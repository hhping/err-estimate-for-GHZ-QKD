`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IBFfiSxs5Cg35h1lIoPCNWYKHZINoNDyuYgep2aunaYg4Gc76mjv5oKLMeoxWbeq
QILkvgTQhWfLmrBDy4exxzr2f9hOCAXoB/WLFz3hDnNhYtm1WRr2kBVHFEwuuP0w
kofqUEQKB9/bWV4ZDRlT8kinX5P6SKcGJMaaclPXpcYkgKwTPNtYuNBe/l/kYCWE
UgzdAzvL3QOUUkQNByHKJoDB47nI3UoLg5EI9nIkM/AUslRQyQsQBuhFBeaoLVVg
deaU2s2UsBCBhkDwYFQLNhG5F57pwNC8K0Vb6A0OPIKe9jiYEt2UHpyjfkvVzR1P
NGydRXUGxGoO2BFNNA2lDEZJuqDl3CWRGotQYR5x1fy0pp5t8/HxbIMKIiDbRLh5
2ONGu8RCVbbzgMC2ofu4fuq0ci/dC2TZWufmmterQtnh8Fn9c72s88Mvql69bw5F
V7m/1FIklZFlUIs0iUzbD+i1Vhg8xjTucLznoUhARi6nTg9SS2o1DjLtXMQwufSM
vMu5ZeVAd/PKwpTefD0X2KD5y+PyuRJrCLaUwxGu9KOLsNusZfQ+Mt5zckt56eHs
suDS3s2I9ZK2H6U7jSiaR7NR0KIZ1AaHtpuHJv+wiS6qNMh7EEYrB1a8LlTBp4Sz
2u80qGDVB02G2S+seIoOjdX3wmDG2n7Hw4z69yg7JHKdNTo1C9wLZTEz9AReYQpB
2ka276ojYhbr/h0y8uPCbREfyomPg5JlWISMJEmbTf/V5BODuAhkeLgxZg1b5Eir
jODq2Oq3UzKulv1l721af16GkhcicCm3Xjkgu+jAXfYGG8IUe0k0O79kq9K4JqR5
9KOzOxn1bXuBelQBjprgYklX09jsKAGWdfqtURLMaQCapatz7gk7MVifZ5G/8Iax
i7ZGMJikAUdb28RaZBHkMRXuk1INv21S6kSs1KERSAa2dEA++ymZcgXyIYahDIuJ
LGqrHxl8g3U9TMr+BlvBlmHAaBiOkHer9eZJgclc/gG/0Od134n+PhnRLTyYlwP9
SaLWHcyJ6BsCzqeTW+4O+HSiKu6uaOZzG/8b0wnspPOIUnZSXlZVzLNbbyvudkx3
NJNs2vzKx6khRgsGUG6i23x4cSFOeP+9Wb0dWKctORjGxFd2TcyAWFNPCXnva9D+
hiXzBPaZ3IBZiYymloslh1YNsaZLa8jPUbV6Xth8Th8=
`protect END_PROTECTED
