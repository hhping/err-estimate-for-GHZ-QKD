`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1qjUTG/o6HGb9s49gU+VsSuxtxwQERg75+s/O9P4MBhZZoLP6/AjHI3QaNPIvjBh
NHhYCOrdRiFqbOUTcZg5l/2F12n6GUBJnHNDnTlwZxs4qYEc3N8E/pi116DHv28z
2FVvQJ/MCyv/pmzIM7W9cCxQfp48fj4qf8o8Q/8sJnJluhbZZVxo8aexZM860nKr
WYqo2Jiy2VRd7IQbXyx6xMFGMEGLktURQm89erwmjKg0zX6hk4Q1I6O23bw88PQE
Vs3uC+umgr62aSBWrIsEBNACPyn3ih3sDP/gKSQPoqraUMPmyeqM1nNu0R9/LO9Z
PwveQv0rgrusWVACRO6O6tRUsNYjaXC6fRONKpqg2wAliR18VyWXPBIXqHBaLU5f
OMJkmKXW0IAIvAZ9aU21vP1gSqxAiwN8aUc6KLksTn4R273ThkjHrjmUTt2slUy4
B9SB8TtkYqap2JLGwgHzeS2hVh9DrZ9A6UquE0x9Zso7MSl9I7e5QmhXXSicAx7P
yU+uaadOnwqeBXKA7oiqUAp3NUkxWPOmcvOjNIxw2nJ7ATbKXHlIXzsovfpYDY+y
OGHKRi10TXXdIeWH2pFS8ZYxHJeveQtpEqFrBNt6nuve36RhLVjYw3tj+7PSxrmA
I6GWvXhnW3j/dmK8/AEV5iJ0W4yehrNPw0pvllA3t0iOTO0lj7xjEjHKYwXuxH0S
VNnuMcB4NYTLm5rHWNmD0EObyqCWUqC1I0VtOqiJ6MJ/3mdtVwBhQzdNd4GMlueL
9G8D3db6QVm63DSmfPQ9MvXFtfe+9ENBJ51kATx8h4/+mYpa3W7B9+9W7nOEZ0TI
1fKXWPxgjAPHil946WJOBY9zGR1O83akwV19aPJPlxyCCIsAGL53WQmLiq5fU3gH
afA+0HncNN2RN20OSBpAMbZtTfJPQ4ObdOgIw5u8inr3ueQQ/0tizaVLzxUG8vyb
jaSSk9aEsF+Zes/dk56RwZKoccpP1gv69WW5SzlNN/nP0FPPyVBZcQjkVg4/938Y
s4NndITNW/HZeWCk7lt7Z+3RAXSDLNHMRz8iH4iRCWHdjUWu43WhFNrLnkPK2r9i
EHx+uBp5JYXPJnCm6g2bmx/tTETjlmprk0Kk9uOJBRa0Nr6UDwfxVd39nKnZYGkE
5V7s9XqiyLDAzwa5XdSqmgIVGdZBBDgyRWwIaQt+nC8KyZy5IduIq2fBkk3M5LMK
kt61PiaxuBbQ8eZEe4GUF07VfFlEW7vfTe7WxXTI0Q3/vdAF9i8m7rZeUj2FEEHO
Yjj2kXuc82sO6gR7i/Qca76/LghdQNyy5hVnpOGvxmJ1GzJ+fiiws6kmSeRvnqXn
OW24TtR8Mu/fRzyszA0tAIM30HrbdYcTCG/bYYRmuHe2JO4qjPRuRSUpM33lH5w4
enq5bTiUKLNv7XtzI/1k3GS/ZftS2+On0lOe3mnfy1M127oVbmZoUKm4vKzpmrTK
diwtZghGLAFLBaUDy3YKAJegHre27USJeAKgKKzyr1jHG5uvue0s2HmBfpTlZGxp
QU2FHMmGIfD8yra3AnVqEl8kQBfIJKJ38+YY+zVxtUU=
`protect END_PROTECTED
