`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4WY3Z2YRxHTnoCdv0VijKilukiwzUHG/0DCS/+OhC/lfylmxrNbGVHxTNbXt3CTL
7AXUXfYoZU/OV6OSUEB8ZFKQq6wVYZJ/3EksnxOxtt/dfxj4BZA6zmw6qGA4wlNF
GEjH1KRWq/Wr13EWN46Rm3J19w3nsbep4eVrpc1Tr7vtYRi6OisO7WX8qxsZ3I46
uCFIGxxnM0UmJA1yZx1gWPToRd5AECnNGMfDjmNDeeDdGrwdvcqWFC68KfuXaaSh
cv6sSR6Ww2J4ZsDDLuecMYicGLo+9PJVrUDxIYzD9V/zzoHf6mXd3/q6Ftn09+5x
/Lbo0Y5Jj2rl4mrgatl9YBZq7OHxNHXQC22YXGaokHdZkVzjEEt12poI2dvt6mcI
Rm016dOEcQsC1GfmwcJK4MbaT+GEDccWDVx+yVPqBrEoHUyAEutvC0egYsMCZ6xc
PjNSSvbVmn/o+1jOSf+teSKvI6WHDR3MvckasDVvsOs9NdlegYolQGmluvy9ALgs
LBu2PSLJAv85Ov30pk133tPnZIGirpIMUy1XuKXHhJopFfAA6tmR9VMydki3IxLV
QGzTMpjqZMU8HerUhR4MLBVvB1hTz7pFoI5TwwvO8+6BghdYWFi98YJfNpWmcEeM
Cgk+hdMk6c623WRhcTDPXmDr/gMdzkAhUkoxr48ygZ1SuznUUU6QnGH8HwF8NaOB
gkB3x0ORzflUiOZnC0B197BeCC3+kEfGRq6BHfMsy55jOLxWLbYm8hIgfJNmiJXo
FUOhyH7l6zXUEe7L/X84qO3GHNnwMRRv//m/9S+/bWEd1v4+g4mH8jKyG1xC3owy
M9nStpL4spm9RG/yC6J5mE6sXU8oqxdCkXlhaL7FIjHdYRGC1QAP0Gm71AKoIdzk
uEeiLjD722tIz6QWd3drqg00kwK3xJEu+xflAMtgsiX23G8JzOhi5BO9jF3XO8+B
Ay7/KSjxeY5bXb1VJLoFwc2584jCqPb43HqteBG5P7VL6Ydql9cHn8xT/0wR/ItO
Fn1smvuZJHzcMCcBgv5CY0oFnnKa1aKGqyDjlOh2o7xAFMWyjCuJxq3I2UffGaIH
oCZlLoeuHm4KDATbnQLLePTYHWQMWIxxlel95CAAxN4mlf5IsEC6nIkK+OBtrvpu
MMFgd211LrSlAVJ9TY6fiGL4fWgvwMDI4PMHyZ38v3eSv38Idb1qPmrg7k+oZmOP
oaeV8XeBBsg9FzKbHi1YZ0w6ipEP57pew+lpg6rkn5leR0JiJ8pnXWvhSk6gv5lX
C2IBgJtgRzq0op/gXwUIzbzSgx97o5aMPXg+qZFNh8rvUUCZY2SA+fjmm05ul8LI
`protect END_PROTECTED
