`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N4NqjNN0IwjCSlkxJ1767YyF+e/rAFFu35D2ceSkFLnOH1yRz0YoAWR0j93fODBK
Hi2MgNOY+4F3yTxQrj4dz16ChtqfFQDQZDHN0IKrE1kVZS19zIw3P/wP1apw4ggy
R5Pdr+/LYK/9nfUo33F1tDE/Xd6Yly+0eDpMS+x4vOJORaMomkweEu1Jz9FzD6hX
LmsTcVVHPyPpcK4aUbnTjTZwmP9sVxedKSyok0N9k9XUnb3soOdrmJQuLLmKWx1/
A1RuDY6cWp0NcM5aCRxi+3iKxgJw4ZXi36H9aDh16Ol/nxTFAt4Kj5DEK3D91O/V
8oLn+o5e67VWLkk1QgxDOF5WMjLUNftIWu/O3nq6L/3RNiVCmDKdyJoTV6Jn/RXR
CSiRw+EdvQ1UenYNZ2VTJBUBd2ZzW7CSXa2OZA52VOrI034UqgzfFgxvaAlwDXVn
+sMAs4aDj7M7+gXLXGaeV6onS54GbQbMcJ6VvqyOODRy8Ej/Lh1l2sAKT3+7w6Gr
1HZHjtRkxNvp6ZJYgkwAEKslgL0jfwtHJzshmzj0MO9qKXCFWa2ZahcoX9VAvOCp
fo/oqV8xsR+y1b2t4whk9IGxKu7xjpD60zhPa9/hZgG1FXG2aAF07nYUf05+lM4t
v9/wRKxlqmPaKpDtYD3l96PEjgjzUM+NXQyU89ijF3rkw7duEaD/fPyYoRyrdR9Z
Io5/GXZ/NdNQpbhJMKxXsChbVsLv9idRypmu0NL2sGDH3ltBW39z8W3XCh9coKO1
ChQtZfCURBDDxggj6hd/EEBLethSOWCnh9vLTwTkDFxV8a5+e5AGaVc1dlIKlRWh
6s4G2ge8vq7QHJMMsG3vHavXsLcX1YrN+gOBenu0ox0841a8qXVWx0u5n/elsGB0
d0yAhn0FLtV18dQC2x70wDHio5Fvc7RPia+SfdQdRaEijqDLrRnBwrWtFdC5nsGi
nKHuF6BRgjpGb8IR4UKnFNUi333FOeRMmet7U1tvFy/huPzvejea/2eS2eQMiEEw
xh7mnkH5/iJ2GJFADBoKpVRbJuqsjpXaqVv6SJwIU0fOywrpbFeOpe45N83mDcpA
yGlLi0s+Hd9/XtR8fh6zyAdholuGrERfSU4SfpPc7uE/RV2jbSm8DEo9+4Re2xUU
R6HGsFOLb/s2cuaQGgbjMdBrZN2SCQY2DWIoF985c1TVhj9Itj5PbR6ZvdFuGEK8
UsaClQIOEaSOZfOH2x39lfynjdXTtfZuWjDfQpitgu0OyldTH+P5pQvekjAZOlVY
qxObPjl7GJYSbe7h2f/NhCmHbRXiFvpy9ibA9u/Qwn0FFkJqiz9n9L8kDr0pK4L9
qiy+MyFQ4sIBt7CK9tLd+EUhfmURIslYLFVTpuhQS4ERhLJ1b3OC54k2v/CiEt9/
rb/Ch9yM+tjeCBfWWGwFqwQwWkdz/2LGDa0YF1NJuT6e4pXMxjrTkBeuWedoX+SU
o0+tWofEXrBscO+k9CmX8ben4Nm9q+UBkLmqDP4X0WZ0zOyuAQYaxTfp4JPy/wFY
SlEl6CjjnnKJZG8HBWIhq/TfW5TDwydPVk3ILrMMjn/VJmu3zXIyex9ZFHaDETB5
TFITGh+Hi7WsNqRVjKSxHQr/EVbNoHNdqGPfHHZN10HiQB/V0Lmz1Qr99twtIbbY
zsphFJJRW1AEm8Sx6UNiT5mFvVP4AC1FnNYGvdCAvmJDYYR9XP/I2N7b2/mhwn1F
jmYu0KFFSnlvIu27sT9vhEKC8o6N7eVFFAPfy/4VaN0I4NKkg+eQn0Y1tHA9rjMm
+JWN2xHFj0PJ2Z++6y0qt9D12qukNGcboSsW4FxVhusgPuBKwvr9gvWmstWljE8X
30DSg6H5Wy30JfhJ6fv0lpwQihdm/HLMeTvERxds9wwXkxJTJrZ09Sfl1otQbi8+
CkZ7rpfGJndOZweOQhAeGzIjMVZ1Yfy8CZzwV4J9cVCJ4JxojERmydOhm9tCpWXn
GhV3jLHt4IIobsuHwhucoNJNtMZwWLijbpdk4BITnjUC4a/cNuI+5btjZpnsxTbw
FLeCuI3WYtAMs2TjvW6eM/bv1ie+u3Hm9LVpQss6SINl40e0I/WdHf/IkRy62K+g
ELf54398iPj5GNS8LwvR9Mp25G43BZNKdeBGUa4rAsVcQcRHCVr6SUrLNyJ7DD3G
UvweOeH47lvAiELavF79CW5fRPPy86dfzRcLifk/8vSAFhBvPbQKs8sKQKAw1EbW
JZCp2lIXZDWS5ikh7RxtnmtLSllKM481moQFdG8MqUD8HTHieenMUZQiMc+WFIjq
Je8gZf/y4aE/kfrLxAv5l+trFixyyMXgKUsiXdI8o7KlVn4mCjAiNJQaVmjnLuL/
VPi7CItRBUIOpoVKwZh3kTIrkSuebViDQjHUJ7Yk/GI5LslM0ie8VBfBpUbir4Rd
Z0NuXfrjo6p5drdm3zTekPoMj1t4PEOpgBW4usU9qoAw38cqfqfQOAGJgzS17JF1
gKDFUaQgByE7UCPGLMgbuLdXyH/4aPAsIYYOzsM++gmIUP8Z/hqX+ussDJk25KSR
Ya0c1YrGWGikKav13HKzbnCIxwL9kU/eq36iZqynUbQUgeRuWxRO83lKOjM9Unmh
5ucnWAN7IvwGgaY/QztMouA48AyAWoKD2/AZgOAiNCovp7HEeKsCfA5IhF2zjb8x
kaHrrFWXZDQxN+tkl8IOAwxRHhclFOmYRHET3G9sYhCfdUxjvvApaYXA3Z0sL9/6
ttWpYr8GfLr4U/w7+YJwchqu91eXN4O61Zp/ZeDJZeJ483dMRxT8wONRrklME9WK
oX5KGceE+XNpCJ4C/0FcbBkhh9Vs1/BFgxfMvhwI9PaRV83PQ5lKK5domYbAAPsa
NnLxNA9j15cbQVU1eAanrV9DBRgIQSpQ01wWmyUv8B/m9MPh1zjzevV3AZqldPx/
QwAEv7eQZRa8A9A+HUyBhA6a1qYxbbcAUDNoWHQrC9cqDmd8xwARes94AeHeeVct
xcZ7Gt48QyxqVTIRHVnW5GCCTRtmEn2kGuaKjAjNcIFguK6Mhnun1pNHO7FywipN
Y3iO6BnAPX05nxAEEz7e/pkdone8cjoanDZGXywgA3jF6bfBfWmoC1qGMyTGjIFa
/C+8Vk+zKUph4CCPXoOyjpOhePgt/GI2LwLIaJSCSRBNe5vEBsJWEtzAmM5sQRbM
X/DNrmWbdHKnD6UsBOuftgylGE+oKhQ3RL7o0aR6m2fFoZMbCZkUGKRdbxaTE5Eh
XKgp10bBa1q6CETEa/1XH+v9hFVUKfkAn64lkxhJ+HNhDJ2KykCVpm7wIgINbmKr
5oacsATpWwzIdZSZKokhp3f8BP2+VzEnuwhghK2NqY75ZOggad++zq8SRL1+7x9/
yBrOiaQmqSFE7loMRT5+lLQvgrW/H5hHe9Lq3Pphzj1GmtnuWaJyk5PcPrL3FU6+
PlobBALuIu/JfYACmLSUEi2vYNrNBb3WR8lkCAQ7fEWql3UaCn5V/LOp68Trm6+M
UHp9iFYsg6/1tTnZJyevbpa0HCRWFcj79+Hnl6cpaS9U4u28xJO8fdoMe9hL6yzW
0i7y66pwLm92XtquQhPLKCjiSo+BupJ6vpKoRoCtd2Kok043ofhd7rcl2JbsE7mj
t2t7IDWsBeuPoLci4oMWsuwom8wV4vH8hNUZlfwQHtWy45O+C+1u5Vik8FsnejSR
MiUEvSJ3F3XLFuoT6crnHsgqtu6psJzR1iDs5RdogI0Q1Jh943jz1v3LIKlNkYzt
CVipE1EjHknoQ+PnPCbFO5gjxxkJeO2ah4HNSFKymfDbhLvayLO3kHK1OqPwwX2Y
xyJwQePtqXcnpz91zM2+vhGi3+1I1zMfndc/FfAc0nb3iVy8eMZ7TI5axef3dJ7X
DUazx4a5BdtA8cVhN0SuFmuS6VcOYDWPiH09zvE9L4EA/j2B/EDK1x0Fwhim/IGo
JcPnUjE5gzZx9TV5SITXhkJr3ks8EHzQo6v/Frrzcy2EXfCIxlcTTZI3ic5sWK/9
+x6z59hvl7kWS1HCGqXReMU2sdrxaZhVzFNT+fWLqmKeo/EVVRcAlVV8QSJ8Q7oF
qGANH94n1mi4z+8E7opr0MwqCumA59gqex/xH7XouwShCe+cKdufks9CP3AVEO36
mB5sgDXH2xKwGU8a0NmVuTpYVWxRNETcrXnX1nwF0aVnOVBUkC0cqW0EDqDdw0hw
k8RcnMxytdoOCsFAbMiDnEf/jY8Oov/ni0rv8XFqA9CQeUa7q9NAUzpW9gPQg6HJ
+/VPjsq3VAOiIyABQ2hz1/jEh3IKukyFjfuubXdKym5X36qQqobBYkOxbDfVk49a
+3iJhc0dH2+diX1TU6p4XD0aDpFi9FcBk40OxyC05iGS4sZRrREro/8UO65oQnCx
Q2IoRMP3bOzHFqWrWaDS6ZjzYrHmDX2V/Bh5lvOlVrYMgbWcxv290MRTEEiQooOD
8ancVHC5cqPDPSrmZc26Sh8MVEt0VsHfC94wCiy3IThfDnO0wJqk1J0CfgKnq6gg
sFZSg8OuLOnweYmcPb4lWj/Gg1MpqrPlrQ5gQcd5hKQNs61CE+W5Sdvvm3MGEyYb
sxDxsbekdkXwuuLguRO0dDbVyUdjfvll50t9p2yG9gORogl/71YOFq27GXgTipu0
V3GHBwc7d0sjw/pR/o++k9u/qlzFdiCkiPt2qFr6uuBKQuw4rZzzMUL3kxujFE6L
PliOy8USQa8HicQvlgONp0zs0k7hT/Puis+gL0JPXZYJwZckPw+PAbuA7lyhk3+7
+HiAGqjKlszP7iWLu1peUvRwFpH6Q9KWDlByGUDurC4t0arjPzZatcR08kct0Cvi
sun99QPzrO4Qp0lSD+9EejaXma3iSpGY5c49mnM6rDE6IxwdxRz0vzwwHmlFd9QM
CN2eCWDXTkmv6xIMEBc73JVVGGFX5Vn8rFKdl5aKlJYr8lgw7vn4QR29QJ+C2n0a
dOCIeQw8Ow5CiW0xPH+BBh5caVxn5Hy/psCTQ2xPNq//FCeZV/9w0ESGd9fJGxvs
32nWeJ17GkdF9NSuHXs7VhCj/J026RvwjmJXqTisJ/WXfAJDFrSF6ZNlD05n+12K
5YgpWwYH3MitG0ZIlwF/jRKUMdbEDIPiJK5wJo2A1ENyadq3WD9nr17/w0/qZSsd
SspeT0HbwpExNIRbUgzNV6ClxWoXdHBnfeBNYctfiwR6ogdv/qLEThHfDLI+0FP9
lLsXYG18c/zTciEbWoRL8rLC75qKkHo0ne9WZW4Wur8SpotYXGyxPWQxhBFNRPoh
LNQt1KGj9P9ldtqnD4IFaDGtDr5AftHDNSDIZ6e1zlr/y62HBKcBC9wFiWpVLRlP
2XOHXSEaravsYe3m8tJcCS/lBOccOmHZVT9v5nnYvNIvgAMSAqsosXnBRM81bToA
Iz2fIYG2EVDa+HULIJBy9L0nAfIv2/C5S/Z0guU/OtlACJCu3tw0ZFCxDCmaXykA
oQerZ+841Mwg3KLvj+EMGidPaoIkU/Krnu94NXKKyhSAoYqzjhi1M9c0WpxcVcBw
yvj/duDSol/eUmu8BqSf+A==
`protect END_PROTECTED
