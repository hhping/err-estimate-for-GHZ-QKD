`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KBZ2JRuKUubJlN3FQrbu09xiTzCP78xiKEzz9OhHsALOmM5c8Wj5pbwVkeAsf+Bx
Z+h8du+YeCBw2dOJu8OZGsx/YyyYU/CjvaTwf8SwbYg1QDkt8ESKqoXxxLaY1X81
XybNf41vryavglGe+jCfZ6tuBiV5UoX+344wHmioGH72it9Xb9iVqpYitQiDhO0R
oLg0XJy1c2zKH2od3R2xaAFua5ChnhP8UGIxR/1I7JX7SnFKsF6L1wQF88/M1ny8
wB+nIKqfPssglSeh+NxLyu3qZH8nyEA3lo2kp3lWLDgR0yTJnv14p0n1HEH8akhl
dM6bxUP1Obo4q2ihvdMN+oP4cv6+kVElqRXcGyh6MYdo2/yDR2kATsnKqlki3L/O
ygTOK0VBqiJkxqWGV+xNcXu9C7hWtQuKbaaPL3YdzAxJ3T+A2kNQzzFN9yA9k+X3
vGWt+gSKgdaqPknhu4mqAO9XQeGWuwhddoIgPAPmAFB1R3rtTvUU1yVhJH/6sn93
HKda3vUfiOFna8lzTHFP3ZSGoF4JKsD+7NtjvSVEiyXeto4V5RXSHJ/g9ynKwDe5
zcuFxSXN0G7xmHZxMgCk8w3bFVlZcG8WwpXxlHUmbF/5BHX6Dho44wRIQQFNcZp8
ErB6bPWKbHdbJChh8trdKQ==
`protect END_PROTECTED
