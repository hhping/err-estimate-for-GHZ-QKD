`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NH/8ahIPWCNU1WAD1/xoD8FWsbDtJuREoY4JgF2PpmUYBL0nVvc4G3nsv2AEQoaR
vtnauhD6L82aAl4DFMM1HG1lOKnn+b3dxNQ+LyySI+0Oh8r466DB/l/C7hYNCdaw
xKkTg8zkkgv/lG3D77xUhGfLuXq5aC44J5RQEJZzpZMlo9b39iuvQa3sBAI0c+Ii
8v9jEhLDWXxeXRRzqXClMwtlPYXRJtO4nF5P4yym3S191ov5b3VuRR666ZBKDK4h
dLZ6adjb2hTXbAVx0PaLyYdasAZFustg3OEnPwWvxh2r98fztixDH+rifU+YUudG
Q5zgVXONrelS8RNjrTzy7g==
`protect END_PROTECTED
