`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
godh4nvFz0Hj2RtdWIRas/F8/8bBgddYD8I6KOgPRX/XDlzXyJRjOuLKWVTchWI9
7kgv+ZlH9UyPxLZ1jAjzTVikRboP4WB0XisMX51oMQvPHsaA+Q4ji9D5jNnKxWq6
nAkSgcNX2NnonWQxxcOX5CSbSIuUEEFaNJWQrCZBxRDlz4/6kxaDdtmt5m4uG7MP
K1y2ZXf8r6Ex4PwAAcpZC/dFxLRGdFLR8C8jVJdbdBfX+E+LMJsTqjJ9HdAedrwX
gnfxirMfcUvmyuJAb9AMIcG6rNAax+d4INbprIiYMkB2pR38FG3oNZNDaxoE40ru
zvaAUg+9VhQwMmORuazFlSeUdMVfmx/wQOk2OahEXM9evDp2DxpEktnEEvezPYrj
bgT+B+Y0RNgdIsI1+PDLUP7dlNRJWAnzNBqc0mpOJnZxLM2wPw4l1vu143E9rX0U
BxtBkmbX8+Pq6LtqBnH3s6ny++f5OWasn6hFKG/FkJ5+z3uiaCRO0pENK5BTO5dt
tFePUlHSLgZ/yCu92ibHodI7PSFJEBMJxI+xhCZOcNctedVe30053nwtgI+D5nYP
lT3AqmQdlA+b3IO2TpJH3bPzF+aP8UwAKNLY+Bp/135QNmH3njy47Q6ReaHgbUMq
cSy0grtPreXzH59naXRStzqd+wsybly/5tcl5ccOU7J9Cus3Ey9ASMu7JRUMx1bB
6M39GAQHrRyVNHs4vR6xH1I89w01s7hOn9sZ5P7ENRWOfNJkNzenSpz7uhgE8Ykn
6nkj9+mvAKehLj1thDKFpaMuhexLHKrQrUEdc+jxfn4diV9mccMWkt8hOpY5QTs2
VNEqmQFBwHvezuwe3FTG6P/eqDUxILeU9raWV8ioej3mbsA4hCPRQ5bakf7wXIRc
EqfJM9t5roXZwU16b8EKN6chx1vTOJBoYHyVIog8g9O+0X0m/oiB3CPLy4rD/XOX
0mwnPJYa2pmKfD0Nxc8oOSolDx9LqA/qTWPi92zpEV4oyTw/P0ymhl/KdY+uMPUJ
PhN9Oddls7izuu1eheawPtjpwHDzV58gKbnEFj1f/awcaq7m/7dbzJI5x1ilyKWD
+2OgTaTa/nx77/4iYcWE8UqLqzkBUp29WWul+BF4m30QjKP19wzGtQKorxTrEyrp
kgA31t8TySvBMUayXZL0GzsvQGXMxaCO4pAERphfFQR4ORtdpuLLMJ8b+Wu6KUxl
ay0IKBANDX2W6uuNL7AcZiRCGYeDW1sDVOIuDLF595g40sYd+voqLi3hUwDPWbGH
cTpxaQiBMmJuf9eCbZ55ds2jm8pVSy5G91u9BAikQ1M=
`protect END_PROTECTED
