`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YP/ZXjfjS9s797gO5TGnZLw4gs/QUYfYAmq6zY43PottVhkh8TOubnKZfmcS4sO3
F4HtIbYh68Rf3oqigXrAAy+Q/ZmqXkFlDzAGCgeBvl9/W3/1BWqSGjkMsPdTb8ql
YEFLTAZ66oQWn+BTe4Ont40Xkw4jhPSM3Vin7S+ND/OLbPHh442Ky5KoNsTFLt7b
jyBcp55JytgsTGnSoHvg4X2ncPbw40OzbygAoFwiY2HKXBHPe0k3pQll7UKQ3DGV
MNu4zk8Yu/kQX5f7SicwcpvAW1+UVZkXQSZDW6LQOstFyKx/oMKJvl4XfwjsiDAw
tNGKjIzBNxZkPZjEWjFUMkaAZ6V+0KygJ72aJPHsxVPfg6xMIAa4LSAdlsC2Von4
247CVd2FvcoGyfX5k9nZ5A==
`protect END_PROTECTED
