`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8oQwheX1AKNnm+fFcBXlw5DgAf7hs1+RI3oQGIjrqVYES6s3kGLYQ17t82HDoOeo
e5KaBs4lRrX9zkMtElTJquLvhTW1tT2VqvhJln55rDidGov3TpAKc1/pBZ4lEj2W
30ECSinjObQjYm/pHMugTa9B93NLruTcWOHVQAxHuLqZqi7hFGWSzfv8c+zva1v4
7g7dnxytvfSoTJT0cZHGREVn4Bgd8wKKax6PtGZe4A6a1R1CbYT2fuRjxsaCkVBp
c6gZfsgNy4r7Csi5kAV8XcYOiLw2V0HKLJQa3SPsRgTX6xPC3TW7etSSqGo/hj6v
lNltaCmmd4GgxShGxQeWTgshLoj8RU9MH/ZKrcsvYTy2s4cVIss0/T09L0exaJ1b
5Owk8j7phdbQNtIILSFXBnq2dmdD5ldI0W3iOBins9FwTHrlkxZpdaRt1txifwt6
5F4KgNrLbZmgv6UHD72aei3ulWW4so4k/4O5YNkA8nmOLB2wmsSJH1v3kL0LLQk+
ox9BJtgqYVhtO8zdRFJB31J9TlQ70BhTiQSb0/1uzGKeR7UWq7/nPZ2h94/AUCpS
zZUhPisPz1L2WtPfVI80knHt7adLVMjODXBNuv9aNUh/0cMsgSQ9Lxz1BPoGpQ5w
IPnqakNPF/10vHGwXJQNOLdckwGwD45a5y/rzTIni+BhOGP9uz+2+pAklGwGXXZe
BbpGRDsgvv3PsKS+yaWym1U0AmYXRNEm4FKvwGRxQswGHX8IbquaWm0O1uohIb9a
9CDmub6QIhgJzq1g7hHfdT2f9P4swvPBCLqQx9UIc0lgV/Btoi5tpDkCFzEni8tm
RAuE7gwkUi3OOZcjO/WChQ1l+BR/EVHET0hhSxlQDhEI9/BEKDMTv6f0whTYltgY
r5gfQ0EsTMxwovvoHiJNWaqY01qqaNT8w1LpmupvJeBeWTESHv4UjWOeKVK0kYrV
dp50xmfrYwd1BkObf2CAL249s+hNcEIwoKNnXUHCgn+/hIwqa6BAFAayc5QleSMw
vkyYhLdTqLXc0U0h+gipzsxqPjSpagqM1gwsYm2u9P9Nnd72DgRR7FPEOYc5B/m1
i9QP+tifYS16zw4RKtnZWyNHjDD9cF1b978o+c131fmyaYuZcr5fwM+iSwGSD1Tk
Q+vSFBmi6oPP/DznsOgpaFZRUwLfg2CcEn02Ws4wH+nVDdtjRuEgZIBjB2TGtRbW
S7L6CVqJrxPTdoPloku8XSLPOFuM2LDSZEapSD5RxLBPhd3BeMLMSguCEcP1SLcS
CUqKdb89wyB1k0wi39bjRuQ+DDjG8M2Fhl7MLlxC3RQsDlSDPzjqzf6VgLeuyp3d
AOx0mo4kJbEmAmCblyGkvvV5CT5++YhXcg7Og8H0vd/uACqfN3Qikk1iVkvBlyTS
hbRSeyHpQcHMpIusX5+3r0pDe0gCQI5GRachSrVGkLvk/RFRWSSXqTSa7hhoSQJ2
iMqqaHLE7NT5SoiFuhC11z9YZewm4a4YSWRFQYdo41lU+ek3kElMHGt4e9rSTBh7
yqiuWbGRwLEFBlvsyA7GwoCicRfac/bn0y0kMT4vEkEMzFr2zT/TGiB+iGWKxTIS
4LGGd9sjvpzdoBMINkmyK02rm5nOlUR73pNXO8db7Ym95H6f/YBq/KnmfjYOX/H9
L6cMcH1P9k5NIeOvtcdqBJ4+WREQ0pKDAkPawNJIWRH+Uu9d1eYfEs/lL96Ictik
rkbfKV7JUKbbaop4dqzhM5vNXAtCpimvWLriEZVFt0lJ+hAmwFh6o0J9LlJklga5
GGPq6Fz3m/b7xtTxzUUDqlCBQiKUCQNqhUx/rk2vdl0x36HpofzYDb49pEIr+gN1
vLLuW+L9kf3QzOg85dhfenM9XwiOY6QHGXv07Kwg6exk6PHfyKI7ZZkVNiw+twTG
wcMvGxDsdPpNdEktOF5qPXy7b8bObQlAhUOMoRZTHIlaeYoHnB31eka7AWj/qAbI
eTXoB+P3F/vr78CxukTzJm+mzuvPPWXN1gb15qb0oBdbqXet2Xz6HGDIHYkVHw5a
sSJwoe/xR5pPar6541m0SD0z+ctlm7q+IUuYpkG8tE4U71gJnH21577mmTlJj5k9
tWhIc+ygUY7GmVeUr56BjoR59xibob+Fs5WKGz+Eyi4Zdlprmr7nRalIo3r8PXd3
E3JRGfJgvxWFvWOn7+TdXERZ1VqTBZFSlEPxUuJQ+5IA1BOA23QzdmXw986thUiM
8T2dS+pfkD4nV3ZSS45FThpN0IyOk+ndwaO7Mft94lbcqg6wUMZXMLDSpXtr8wOp
0xkC+lHHXADtd+m9QpXoXs0KVJoJ1Bf8lC/ol9dMFGl0She3c8wZqoazIkyt0GOz
/DCLMyDvk2g1PI3wv3IAiHHCRKQoHY5n1GQx3Iofj6haXeX25qeXQl003jPC4n4g
3Mhl7jlG0IpOhl1JQfOgFqFZ7wsji00W7dsB8qL7O0vSbigJlZKKRIRAZEu/HhCn
qhr/gDo9p9PO8XUvCiyNUTwhLoNflBddFixktI46YLadlL2NxeHjJuj8YZjZ1mXy
h2WDGxSAwkvpK2nKuln+46+Pud9XOac3kkfisKBZ8qEaeUtbJGAmPGJdwjXZOWIW
HW1ECyXOUE9WkpTsxs+0ngMlJLIxQ2M4Jqa+n+vqqdrO9cZwVsCtsDDek38Juks2
KFtb/dUO+/cFVGmflMSIhqOJ2pd65Q38Mltz7JPZur29m2rFDCh9UaQ5ba/QQKAK
QJvts45wBpkzIQmEusfNboawfuYRxq6xGS9zZyKQlpiKsdHBY+/cV1P8i98D+Cjy
xlCTVnTjXS4wVfX/d9FHCMGeryBQXTdpiIpuFE1/YcfD6vq1NkgioNlAV0x2uysy
EAsw43j+uMhAeX5mczjdNx7MQhDMcQUNwAF8LR0ujr6Y3kH6VQzfM/wKhuGxdFCN
+63chrcz2VgzpbK8sxaBvjA5sB9uHxhi2H9Kqq8f2f6HspCyTAhp2sLfsHql2O5i
Mmq+D7U81ModX9Y/A5m/21H4qixf55ORm/Ehn6kfvYPWwbU9sW4lHipagwg+TGf4
X2I50Af1487fMRCdFy+idmE0zmYn/B9CeiNzU7upApIcQP2I4TFASIQJurxjGkRh
D2O3q0o4+OruLVpdhkcpWVmbiy/TwmEvROoHJYgoXR7MSFmAq0XCRCloDr8dsOs7
yaBGXSJmGrJcznX4edSFnyqpzhgYN/PqWaZNMgwm3xkd245vQupdhy9fflCdaoU1
BYCYPqkc5DSoVuNTfQ6LOfkZOK+JCh5TS0XVm2Opn4Nu28gohlcZBe1AneNg9jf7
PBbhx+rysyK/ehQaSf9UIboQWnIXPC1sKl/9wNlEvyrXyyqF/DYJRpdDncI8Ipd7
D8zDV6/v4gw9seO2vC2/BiconXE8J/X9l9Tpk5GFtB4zl03q7jp/oLDIla+XYuHC
t0598E6j68wukK2/XmuO4bMobqGPWLFxGWrFuHGf27BdoZXxZMQvZL8w8NlYGNcQ
W2PWSYgPKRzUW+N8F0+vBOe2KQp86zhawnaGO7tmZcZxNKH73zNt5PxOcmafcmN6
Y3XzRxDXfK2Ysm0ePsaXI+zDr57QRYNJKzIFCdgeygHTzUJ9ZuZYAFr/pcuBsZ2e
yj2EOgVsaw0sexL9zb5+pPiDOzRVTWKPljbfOgOfXCVCqyfFo88DQCOULBarQCqa
6Zqnwg+Usw1PtmnydzHS1BUUZRYhWeJLDwBjeQmNY90o+E0hBTMvhwEWSrTMZ4Uf
LwUeHgXYO5xKTAdoH/ev/CIkMyeTObZ51hDNpjqOV7V3bu2VkalfkpBgP1crXHyi
PhLf4J9AAmf3spy/oXc0gxyxpXKPqwbflzlHiLkhcCJ5CsJz0X+8/VgoZaX75Tgx
seI+7QSo9oM46iyXNKC7HJMUZhM4/PT51RfAldYGJYns1nz2Gq2XifVuIykBkUi3
mK1L5Xg6a7QYmSKZ64nDQrto/RuDHGEmiM8oyu1ZDfu142APbpFn0dz3e3xsORk5
g7++9YOPclG1foGYlKUFCIbQ/tQ+j8iac6N3UgbM/PfyXDoIuJ/EnV1AsXl0TtB6
uyLNe/JxPaXAj5CH1ufIsoQHYGIDBVJFJ4ubipiuF1b0DnkwKKUAYwJN9yMeNGyF
qk3tFC3oOD/H5lom3VOpZpJxq7f90LU/mdxtAE7v1GdfVS/t6yaXB6oerMZf48+2
N20s0QWJjuNGFmmPO/jD8KaHv81pdcUK5ZlFgNAIVX/kmBS8HWzupf04GIAbimY1
8Rz/sjOqBNbv5e4ArNwotVmcaoq+74P8HLCi6Dt7f8byMwMckl8FIGzpPnHA3fMu
kHeGqhxHbLdp6DLohaDSKn6GSfjb+iL1CMQkvTifk2xyoR+TbSEJM0d2j+IxskiY
ayoq2hQBTr3TwDxoKzgTXxYbMysoGmq3c9WLxZ5dOcKrzvEHqRi/5grEKjJ8qgV3
j9MaVOMY7DJskdUxMqmJAyHg3tCPFPhm0lv/Zg7MdZX3udTCnJAyEcFtdf14ErsT
PfqzMJ0PfzRuLOxO/0M+yQi6DBNeC4919KCBKRViWmUO5MSKvDbfANLJnnPACfSH
L1KlYkGpQa31IMIdMBNbMP/cPtjEJNMKxrswYx+c8Sit7nWznPTUEV4ZsvBHCndW
nNK077mknFZEb1ceSZPc43aPRDtsNsRIZwhdAypsft5V3YikKcpqFwJn3RIddEk1
6nKjRovT5Ix9XP9YXLxrSJ78eUdWyIi46V37GKa1og+waNQhBFv1ruN+46FBESra
2OF/At+JCxzEOfSJnwrZxrjYq1Z618eGRP2F2+ztYOcgfwyvHHyv9WhSgqIIbS2f
2UdnQ9nLiQ3f/oci0fPfC7lVzkgM4KCo/EFKZu8VEC2uUGqTD65NCtKosYa+2FF6
sYQ5BTp0LiJQ7Fa8o2sLZ2Y0nueivJFyVXMlK5GBiKzrXDHTOVQJI+89HUL6Epuu
i/TATwIlD/Mw+Atr6T+4jcBzn3JaerWNQjByU6btbTBk8e7I+ZbPWXn3FoMAQ75u
v1ot3vX/sWIslrpk56LRHLQVQBsO8OTA1CWFmqkFhJsEMShj0SZNNwrSJ3bgpMxF
JvXmyVdxTMfd2YAZweS4/pYImB7RGqbF01xnAPEL01HGXtOJiy210B6baO1kTW79
7PjInLPmhvuZWPy+86a3zgdzKuJctH0OMFrYqvIoWSCJMPfPSZimyfYQY0yIz5+b
LZKDcox1wpp7prC9hbI85T9EVS2No7nZP/nl5MEImHJtJUg0hvWxhPsFQqlEgwM1
YPL9Y404M2yLM/hd3nJe0BDYhymvGQcTS4FXf9A0GGNXdj0721bjnyVqcpXVKAKJ
8R04v6mosoZFcwdJURb1jV1cSvu349uOnQ8SwMHMKAfp7QI4C6AUm9VgzhmELyvJ
xiSecIF8gnQBNODp0b7lcPrj99BlBqipgG268onCaAdbLHYh3ZZPT5k5Rm7q67C5
MfkSlYLql+sbUYi5YwQPpPIYloE6YppjvqItbWI+mMRNtYn9cstRS5jh+MjiEzaR
9/+riFsOeSL4gQVStJf47kqKnyz6f/fYEZjmsysfJIkABKJdrCIflRmPdsBuJ/aH
v/F4G2e4tnrj5B7PrVgx0jugYC1wGp+zJDmt7XPJxTqRdx8TcUbIUWiXSkvelCny
gsw4GHOHFQpBCe/aeunhe9Uz5dBJ7QmikfFAIBPhnN+uymOKAK0PlcwvaPrLWX7d
Tgay1W3xroKcG97TXfo95B6P3YLY8Xj/w73WGngseh1NcBQIBZ204UfN9YEywyWi
TfJMBNZHvS12XqIq1SYKM+Fwir5Or9hpwOIi2Rq3pZ3hk8mLxdZhZj2dyvMxDGVI
dZztriiUxgxjE27mE/7ATXTA9ZGzr5eNdfOG6fvwmOqSnSZPI2KHLbplTpK/GCaN
u/f2R/17UOs2xGbh388D8O83zpqvAOyRThY1Jf9iB/P1vmOi/AQO100t5oC1X1RD
x8MNbH5MR045VaVVZ6O+IpcZsPNvdHehrhIw3n2+R7F0J65YIlBCXAT6cXdjzb6G
LB3Y65c1X/Tb81m4jYeT+UWMynKnZAR09fSgst+ZAFzsMItzYcoKPFcS5pgejpv7
kIfETHyyhm59LkWsMx8b1sfUGBILE1J3oaaMiKV+x4zsHBkrBCeu+V2EgfOQ3N04
OIBPv4wWkGqew7A0RuE3ddEiE7RWpwwys8f4A3EhCX/k6Zwc07TDJ/wyLlA5z6IC
EzdrLelLyAB23bDSyoKNub3D3QCmdAoNInH1cXBNacQAx4Y1495FiL0tTG3AgoVX
KMjvYH7l35b/MpFUu5GU6MdsrYqvsmQ8aMdSz06495+E/eGACpzKvCQYqtWuL6wm
PcriJ73r3g5LZrr0315M/1Zl70pXLc4Vt70IDfWOMpd5yvjYCn101hcXO1vE3ywt
6sZMUWkjauG6bbETdb3QyWjaFw8e2OksWTqs2UtDNuUCblkoaQplGapIy/mYj/GO
hDn55r54Iv56VHfXZPi7qbZ32LOaa4ad8hvcRiLG8z7+eyn+TiFakY+KyFDVpm6W
y4mEbCl2xZSI8wM70dnXKibKwGeNUtHiTiRHURlkCnuKTUMGOEaBJ9fhupW4sC96
jHguLpORUxYSZNAuKqMvZudxTtCKHEGvpHsLpSSxjX3+K5CpqENmJp8Ep4I5VLII
3Q0C3FkuCmfJfUNBVVxSevKywNHUH9BAr4m9e2T7NiNFX3Wnn5ZZ+JpB28QgegXc
RZtkSFOowE2WBqZmtbTb6eXHx9rc7CF70lBLy6XGfxyxdSqL+9Db5rTWVE5qsi/K
MzvDLaiY6O7SEhf6RbNK5lYw/3cvs9z+VCXS3V8v/8SlaQUFIDd8Id23XzazoVAc
WcZfyysm4WBUjXimGK3ygH9btEw6pKT+6A71ip1q1LQ7Gy2i/YGTKoz1/TYsljVT
e+coIIXd2mNueLeKQAkD7z2qslbGcJH417Czv4K5qTGce+1ZwG0mYX60ARGIP0Ac
dzYZsme/fEaTtx6LF4r8Hcd+LijTzXADaxsJNAjyUqiut5QZf5WDOPsnnb/V58co
Wk7RP+3XEUZTNRxk+wMREZFaEjyomw0m2JELh3M6jecTFYATj0tht4Hsvz1xMcz5
8v4YUApdQP9Wsb8vlVTAYIRXI4F8MhLdTEP/vfbe44rHX3A98OpCQ2Rtva6kOm2Z
3TLw0HQvENVFaHT7A9bKJZy6iKgKvskFungwHQJoMePZshapRwYUS7L/Bl9wW6PD
2DYqPIZC3FtwBNlm3xRqidlTMBSYsgDfBtGm4Q+fsadUd2RyWWlpGWcdbSUsXvxo
sRj/xhRDcXlVmpgy+x5hW0HmUlfnM72tkbrvqAHDCLnqIsx5laIBSuF/VITNqBaQ
8HLk+jDEHw6euTJcONJaOvZR2mLxsIgS7cjWBPRL7zK9UbSIG+WNVgIiGFiyn9p5
oTYTZdsIw85GoJmti0Cokoy4HYdIbXKm7BH082kOnEZE0nrM5slVDa0YG9kYOPiN
2dg15Xnii6wxuTPxIxwJFcYmf8goOYgT0/pyuwKmwO252rqaRChZFLbbZaKOGN9a
0YD9jaQu8tt+Nw/ijL5T4hXjCeD+oBgJxxWYrHr4/3kpHerq64B6tWVgl9xsHuC5
eSLGTI9GLKH++ss80yaDQ8CrZxwe3tKEFGNF/YS8BJdCjqra0RrJjWLA5otfe6eX
T8Qi/d9PxXtDuipF4ij69/FdKBChVDQMurxhVYfkcPSYWZ6Amc930UJ23wVRCtrd
LFsRZPvYm4PIaO7pZK2b4TU/YwQ30/OSrmLFcXS/kXnI+K6W4RGkKpHxsqhPqQIV
WQ9QEof0CUhE+FgUGSJ/e/FNV9TuXoy9PTw4HwXjGjCn6L0VZ6mkURIR+hBbr2sZ
lnZSGhYgYfpjpPV5GjF85zdFvn3V0wXMa6uuzaQVmqSM8zRfLIbOOZkyw+si7OsA
bYTSGodGxHyRS6RWGxuJS/5fRzk3t/jEBLQR8tpMp3o4q5HudOVymjZgb1jVJkZn
aL911cSIzabFUCKfF3UWlOryOI2RHuu4D77v8Xfi3oLBCkCufaJCCAe5EQD1OU1T
1sb2YzMyfL/bLM35ev7LQJewaVKOfLly/ESVM9W+pDHqVj18OQLXIjs9rQ4q5EBw
uVC+nKI1lVpRq+wVIE8LW0Sc+tsBAqInBLJUXdXNualtosOWh4tIgT44h47LVPs/
H8dsqTg0uikD8tnjQCnzBCbK+tZHidoPolXwKszZ8JYROeZumtdI3N9P17x3BI+w
sSVADGgnb1PSiAFXZ20Y6gKoedHnQl5dVLDjrOL6hoAYr6k7pF1kBXdOZZDqEY5h
s0N0i7tSwSHu+zjMxBclcAiu/8pDYnjjraY0O8ztqqeq1GpY0n2Y6L4R5rKlKxDe
Jss7YyHwlc4D3ljAWb/TZJqnU+dbw082PXWWiQOR3JdD0S0zKtI6oe5n3u6ai07A
mGN7yNLOX1/PpmyoxLEqQrZiGX+CSWtrVnC/cK6mWOAB6m9w6eYhlyMMaT/nyHzd
U3PWlzCwTGCJQBY+ShUuqTyzE8O8e3a+NziRceNaELlgyGsys3o9ChQ7VDakiMuH
CH+HNiAEL+FjoeF8jEe7VHvbeNdBK5yQw/h6rITQ5rYWza1k5bQQKYq0nLxi+o+T
h5/2dTFoFzW2fKDeft3x+v94TLDdelYNcP9/qallz6njee6eYxQTR0d/xWVBsEff
vRmzMQtfSZEZ6GjlbGhdWtQcuWcaLEFUQV/PxSM3eDu5coc4buA3qudobCn14t+d
VtgWZcws2/FkM4og7akbR44jXHhfpjP9r0Te1VU3BvWOzqid+VQTO+ibniVq71Em
naZMvbMHxaDrCGA+GFJjFqlSea8dtijdZjhgZIk0wuOvy6E2DD7JZkK9P3KhaeU7
VXUAyV9YWc98+p2WoMONWSiklavjMpsr5Xa0RmqNiMA=
`protect END_PROTECTED
