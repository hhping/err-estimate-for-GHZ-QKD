`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wuzLRoMY1Cg/8NyKX0LaDpi4mb8EBtOMBVIcZ9DK3c0uu30glQCf3UDijfGgNK5T
FnlorlJyICvd4cgVJtIjPUUiCep9gVhcijFYUo1yL2lHVjUXYAoCpgIEGkRSqOuR
PH/pSSgTjNDH8jqIeWysFC6KtUlSnR0PRj+FV19H5GQYs8i/4iu3Z6Tu552O1a4x
IIh3m1eGReEwRsfBvw3a8vFFefSVy7gGw7wMScYyeAi7Z+55eiwBLDJYK5G0na3r
XrrKNiFCdulD60+fvuszJJGf/BiGyL1Mddo8ZDkzMyndh2WBy7A+gld431HLC2eF
Mkx5slroe+auP3Hh7uHtuH2jrET9g4j6fqVCtHnyZ/TG3g+hHBwLRG8CeMJAprjo
5GmtLy4CcNvkPIs0Ku5bTT6NYt8CcLdzVgT6rPLZGndnhcpK7/Q7ctLMRg96TZFl
Kg9SvCZqhR+VUXrgFxesLVfnwSUGvOUCYLmTQDjnZSlH/E5O5AkFKSYZI70n7sCO
9vjjaoeD3YzyhBOoastYIa19/Y3xMXtCL11Xn34yx5YX0CstAz8WaH9cJM4p3oNw
G4kPg2wqV0ug4Og57rKh7EZzfe8mlT7bnD7FUwmYK/h5+GUtNKNhCG6tM8IDBuv5
bmxhdryUAdnsFnNhwcXT5xp1SeAXBhZnLWsz0+2eSQLhwF9rfmhJIo0Q5dFkOF90
FEa0pUkBellifQBtoJINv3ngMHEw+/XtmMwNfdNa6Q+DxaTem7PHWFmWsmxavCjq
q7LqUep9iYAKlo6W7zQey63DG24ryxWANGEshJMlnnDY/6MPehAy06JA6yvq5nMm
WCSu6gQnd9JmuXacrO7XOuDIaduXkVpxGNTgFpnIW738AwM942m1RxnxOa2bDUgq
6HzAl8lRSSl2TwNYs9Rry7x2lDVAc1GlfUmXuD+6af3l5iZ05wCAGuSL7gGhv/hx
`protect END_PROTECTED
