`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rd6CLBa9UVWIWsAkhl+Ms2vGKn6z7JhpAXPXYO1QVInzMfNbGZ4ZUux4OJIiX5cY
Iu/MvvkUChImCn/hMwfPl/WkenP1lv3/w9dIbDgv5SsYD1DHdFCDZnD+B2a6itES
0lb2XhhY0QlEMWzKLO/ZDuQr1r0GVU2sBqhV4128hkLeoyevtnFcq2FxgC32Pa3m
c/8yPOGvUKtlOxoBgl3VncFnSZ2TRGpDXkf+vt394xDagKSymbky+R5c5sBqrGdM
BXVVdQu+MgaiF3lTm6+foNbtE0TZGN6RA22X/H2sZZw51G61KqNJmnrHOsviPxkr
Xyv77oDy9LiWsj5ChzmOgKDG/kERhk0spFJuBgXnt9sHor+98Y2Cpai0GxbevpyY
mC4CfztEWgYqu8qrvEIiQ1E+20H0QOM/FoXvKkcr+BkjPn4JGG7syefDKZJdq+Fe
`protect END_PROTECTED
