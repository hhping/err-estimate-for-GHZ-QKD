`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YSgHewe87P/EZp9s1Cp7kWf+eE6NBpnhUOfsdDxbSaKe/7oSCBLwzcyvOWfcAS+4
xZgCKYWZTTL19xgqZDV4RxSoTYV4pXocpPaiwKZ3g3OjJnwM5QTDeap89bNzmcET
mmQr7XoNCWfz2+tRqnvFZQCNdMCfZKBsUJqoEaekP9ntJstkh+WyEg+XySjfFL6Q
7mCLiXLS548d6tj5NDofqZznsd7/6VaMPsQWtYUauXgCWhtv8Lgtp2ipJHZIQAA8
zMu9ttJJvq939r1L3RozGVq8VR2YeNW4DqTOl2BdMrSGA6FO3Dsc2AWRUd+5B0lK
`protect END_PROTECTED
