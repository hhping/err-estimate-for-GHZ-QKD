`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iCo/HU4ahZLAeih6O5cEa7rA1jYSx6BwbNb9j0UrC/tP4gXDQH4AGJapKksv8ozy
wOYL8ghJNHp1L2YZG3xQAX6ZMgGik6NlryHuTkD0SpOe5Rny5fzfdSa0qwcLbfiu
5e0yqHrHBHqHxxuMLPQw6cgwAiSAnJP2uc8+ip2aUirIlXzdlwoZTVWmz36ddaA8
5VRUEQjnl2aCvZhF43RCXCK5Mf8OMp0wBfVldnrJlN8ktxZV7Yi6OWzSvm0oRykM
Bnfrs9EzIg2lN+7B1n9gPRBHgCk10xRYTYo2L+uj4ffKBZMW/l/TFpE4bDRxceT6
v1TmwKLTQnKlk8URRInQ2UU8OiQ94BqjFwJfDjKdQa5uoyRIBelR0f4xe8oxntXe
g6z5UEDEpe7MTv+1NyjA/B13nn97QeTVgbcV8b7V58BPvhEK6FKAzefOr1Xctutf
qoRVfBrC/w+EBgep2DCUBoIoYTEkCB/QJOOcm5WdrM1hfUlM9RNbx2DVY9Qc2pi+
WJxG2ruTNk/xLYHzilKny2mFvm1LI0eYSlSAu2gjQKU9MGZtwssSBSBS7lgrZGv9
Lp3c3Xlv1LujqSo2/oAiqCyMM3ZuI4jE6qpGqMy9VIzfKHK62nBW3ZGHJAAfkaSa
X7XQvqae1/5EGgQiomZ9qQ==
`protect END_PROTECTED
