`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dtFvRR/xoqhf3L5V4FKi2mKxNFVuyV/vXQ15ibLVBnlxdHXOSBEgGTR8sfbIra/U
ncp1tJBfh/ORLfu/I497Ay3QNaM6PTJlaNEFPOQiFl58ib3mU5B/JvpSBhkdjfVO
9CnOK+ta/7PExWj96CBX5F+DGto5fPPTz1b9RQpLhw7E760kcpmJdfUiN0CbLfVx
L9fJqz82WAJozRdCW/Kqs2rPmNjGRy1oa92mv7DzAm21G1AIeo+4MFHiUNJbEyC9
LRLTFN4FlqA7f7jxUiq3a7ZUZKR2yoYRvK+U/ruQFwl5Z8N0JkzGahjNaiIBPhsP
b76fnVaI2yuXdAaKWXgwjsDfBsgcu3Oh2ch+holcizK/bl7iVSxqPkPlRu47rgPK
K9hc8VEUPc9bvnxlTsobW6Lulc3SAnXCHsEcaFOvUN6f8yYQKvEyGgzm6U3GT1YT
Rmc02Pk3YS7qBl5NQH9fYEEfwdzDQGXTyb1nckVahxo7GHWc4HvCJuKnzedEanKR
tM1AvigbfYxX7HcdJpljIfNuDN05b2KXp4ApW0U1Epuv6VT98T4bqje+WvELcB4W
Ugy3om+7mZ4zg0tEy5SFP/xcRR/p9bm0Kjq0ZkSiaVNMnyWj3f8a/LZwsMOS4rEA
5rYyhe9X6VmgoTwYLnfNwaZizvySnGBPTHv4KCJOHoZCXu1y4bDtY3FInLy1ahGl
opZdK0LlsNA/8bo9TuD36UZjhE3DYUosKgDBRiVDHHaq26kLed62GMhhbnUcwTY2
Gslcojxvp2ONrFcQdcwSyOjTixy8Z//p+RGCf8ijlgxiMh8E8YgpBAPgjI7tceSI
w/czpaHab9inr+6aT8F6KJmLS8ZB+8X1ghbSnls7YVg=
`protect END_PROTECTED
