`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3Vf1IlA1+VkRqg9445Ky4GFQ1hTQMbX3u35xCaYMvbclTEIz6STkg+Fty4j12+Cp
aTpmOIA5XPCOlNOQzGPr7RkgTmbRy9LbpWSqGXItvYGouEfLFbmpg2ncK3nmS0V5
W+6tv6EyX1Cz8NCuy5MvIVcNacNU3mztkzyj39lWbR40trEv5EdN1aPqWl7EJllE
XGVCud6oWq0UVf4B44vnWLHTkuWdThbrvQ7r2/VODPXBWkqKZRm3NkEHIXL7k3wB
CaXAjGua+0T9oDDQjDFT6FcnAzk0Yf1cUqcoSla09f+4HQyE18UrqLpBAxdjIfha
Antvr2tfYyO2X7y6hUbXiVAHU7bQmIS3ri9UBzO243aduCDCuva3DwwHTRr/1/Ys
xe1L6hnYhhO/vPMw01HbuolQzNhfX4+4lWt92T9b/btyAMblyzJRZpP+lx6xjXdU
Ffr5GIaeW29SW/wETTbHAZyJojBz9+LguZBwU/pQxHup/fZJFfa4VsPLyryqY4Ct
3F3vNUddz2beZoCWB3vYGFFlJtw380Uc/ZzhW6tIp7DbUAZ1w+D4pIavafmRrLbS
j+iqP957xcBK4RZoAVKdqIyTxSAFfDfcfQBVddL4rTK4CI5Rh8QHp2GqLrxwF2DO
auCfo4+67mJLsEQmA6Yi1dep2PpiurvW6jPT5aMQvkinthiuHIlqI2C+Ii5AAw/B
1dj/Rr8QiOrHe+q0r7tMEolmWKa/GKG0rofrJG6FON6VLOEtOPPCWAx/eI22deIy
0QFurjd2Ix3/k/XR21rYSEiaIHRrH6g72FtrkU4OoAcSoRifDjRWUj2sfmlUYNBz
Zgw9Gbh7L1x6ZAmmut2KrChmvQQeLTCXXRCiqWl7LPuYyHcJ8El82sbZ3QQ6laop
6UOZep/djnnp6axoZ9YyphBsLQ7DZPvTXZtV5/7pIrRfMN4Gc7OBu138GOTPENIR
4c6R0vNyw5/Mk3oDdndJhYgMbviP1t1CNafmlb0nGj3P4MlvjT6yVle+RhC1tTOI
klfijkGqhPyTzSol6VQdzI3Odd0QOP3EqKISDC1pbx4u3xSfNfquORfhRMXgpmWl
UBR8hzI1ev1f0qoq33BJrx/uqJrqEP29zIYagAYuax1kTX/uRSPOkbxK/mG42vry
J1gtE6BhTJw1bedk62odnifRvO3g7Ft3H/78/keNvcD7EBRZLMvc14XP740qewYc
sTfmJF8UiZS08bJcf9wdslsnN5ey3mi7+ra6n54FTOfh9nrmVdZiDmCm+Cl1Su5x
cKpdZUc2dqNs6Q++UoU+pWWeLJ51bx86hHrK43vv+Dx0GUKAt/mLIJIXKwk3jhBM
PbM2oXg+9lhMbdk/zuiCmpJimaC4W9KALjo7/fPvYAyN52dap6MmZ/GSBQnYnhwJ
qMciafJ6SOLkRUQ3NBcS8k+Q8ThaJoHVmWHTE1nJZKykROoi/F+XDFe4MgOYBTJs
OXSg1Pb9SjgvtQaJIAPOeetmBaEXuhM+QQLRRfWL/JBrs3xzzM4TKt4t290dgua7
dVJQAthNVAVZV10JbnBwSVLFVQl7nLkLxtAHLhsfoS67PH7ZdYZNgiQdnrd1Hhw6
TVltrOwnWLwWEEk5kR4gHBF6XcdeRxnqllFD75T7pwsKVdxaszFt5kmoi6/+ahZ/
Akin7ZLuLTqUhnJvAwTsgYSpHNw/UL+kpd2dk6Dv1r4FeO/vyDzGpa2sN+O/Nq+w
BkpgWxQvagyFi6UcApNA7zTlrTykU2Lhg/b4oKf8i2n8TimA83KqXKsTdf7QWnuZ
mPrZscVYQHF7ZqQkRzDeIQXZJIzRzWwMEQqoxxbeRP+TcAIrUhRa3OXbxSvdMUo+
cbswNijLtKvUZtFSZd5wy+h4Mforma329ixoeLj0SU3sdDBgzWQ4o7TW1fzxzCoA
yJOJXhjxhEtfLwS8RM1F3BsB9QjrsOy9iMjAZJCoWvvw+sLI6xgyMaHoTEY2C7Nq
CB8p2NkMdaq+8b+k6B1U8Fx2g8w80RG5f8bU5aylhvSpXQCRCdIuvGpDadYhzDPb
L41bgFBmqAe/PxH3G2Y/zC9Mr+MgKg0uiV5DNonO5me2EL5kK7quABVqKZYFu7vR
2ECzlP9WIFfy5STZ+OpRQWII8122dJNimX5a09H2+RFS+yAmBpcg/qxQWbS5nbxM
MQrH3iVJAjjjgpp4wCUd0IV58RTBxr2GypQKP/1FKt0HDsRWaA8HdMArkV8lVe4s
yKtvilPx0JEAQ9CBzSxqVEMNQo00k1CktQXFGNy9TiiEL5IaO7mVR4efFv7Bxhp6
5kii9jmwu+V6WIjSlbSZALlavp+rQ9uKdTz/W8AEAfn4tlVz06KTF3P+2K2/bN6H
LWAbbkMoI4W0JBcUnrCzjBEl1HVRnyswNlrqZDcuFSlqY+LuEmGg1lNDjlDbmXYv
bKqndk6BdLrpaThylVQQ0dfnhHLWk1fiFQaY4uJ+QKatyJb2u3pxNeAUOGTMEyoi
G0nfpaoCLphpeRnMrUohRjRCPhYRfQYLMKAWV8u4vFMDnMCUzCJDGHd4oO/om+NP
SFpPkJJg63iWjom/aKrJF1pxesxLJtDjKPDpAEzQfaBqZmZTvFHmguohl+3w/Hfq
10cQIpurgf3aNGM6N8hKRJPsna3rjtvDLCwjUwdrQ5LXR6+DOVLQZ+SUPkTT9YHe
lWBLS5G438tRh8ORb6/oXTw2j60cfU2bFhm0McuxX8q3cX0cD2ODKlEgJbINE/hq
5FB6at7nN3XfUgMs6xnurv6+DpJQwgbeR+vcJ+t89aeA4kqqmztCoYyT5bgTcFdo
q8T+FF4zFoUTUpNXRIN2V5T7eCmtnsDz84PaqLz5ast6vEIiGNlxzPgWAp/L6U8u
ioB/VHL/UmiQ0/mUPX/VS8x+pQFIDIHmTxFDSb15EVYgtx+Z5rqeycLtB6tDD5/q
ckj2weixN0YP4dovXvWq7GCmLWyy1y7nDbVXnNclA1BUodEbWgKhqMIpBBq25P1G
P+j2kdvpDUuUTtWW4pj5m+6iogiLufIcT1WbA0aKWVZqMTmUOEwJN5OOkL0ZFNIc
4M+HNy8De9DqHAd23DHQFG8OW7ruCzZbtGrzQLc0E+o=
`protect END_PROTECTED
