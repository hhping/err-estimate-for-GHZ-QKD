`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ppwfiWX3Byw0YlENbIL+asn3eCN0pLRKijKjq8k2zJRM3Tco6hjEypyXPD0+yGdc
Y0v4InFGMg8xO6FLTmEX4aMXy9ogtQPnKYPznx1kM/noWhw+gAEckx2BeZzcFOZK
NxkCYaUKjg3kBoVMSfEf076w0CZiLzdLpAOk0nFL3GwwdQcJeNgqbVesjkZ+T1ps
xyDL38JVjc6W+ENy44cOC4wCAsiOjXEXZQH/wgtbS1SY6P1dlX9cNSHvhRqcPC8n
ptvp6RYazlpPQevWN/H1HnfRxD/uaP7YNxmahYbCvvlubiNCyMDN+dqTpRH/wtH4
3xNHDH+5EIi5WmCYtmzFWViJpcIqIg+5GGihtLDo+12nUtJWsMNWeT2eIzrbniFM
vSNEZBn6ly4eXoemK3C39D6QkdnRqce+UBEbWtXaaiiKsao+0py8yLZja+Dj5E3R
FXAhNFf1LMxpZLhl+PSxF3yMA00EEJj7TH/0hOe2I05JKP8BflipBixBfv2Ir9Bl
jd/us1oqO1kz9lQSwuXEIDqOcXLp15p9lLhSru5/b5EP2tS/knEULJEvuXs+eNx4
axd0agsZnq/6JLR4BSQ6SzcfaxFwPTnYWaVtOUa/kpT0uD7id+nT5JBzzvFNpYTb
GrlFe0c9F13a8ZcA3lW0VGqUt+y+N6iUkBGhIH9VtwF6HvYlHvMVHhPjkeGWvBHr
gaprIFpzzDOi2WxLL1HODZESkV/W6uQDYwscnYrnRXG2S5U7DnLLFf05w9iZ4m/c
NYuLlFJX3sYm6bov7s9+ihChABH9Etp0OW/ZmQPzNZKttOWJ/sL87Y2DOL0kP+zI
+kE0ShqWHQNKRimdxxjLMkUn4BOZgVeWDhiKrGbOasyG+th2Hw/B9i06h7bwy94h
QnndSRDTQ/ZAR2aoU4a3BDD0OReLlMsUQ66mr4d0ds542ONTC3MAjfOa2Y0SHMwg
mO0BLkVi1oWxbQAkwgWHA9udVRoY0hXcIOU7x1l7ek/pIMdfh+zRwqC0newvzC7F
q59+wKGFs/yAISLPxlCd7QCfU3HQ2wyll61f//LRwijB84rWTQzyb/4oLL/ATPHj
++nR0+bGB/Jj47bKopoUnuohJiZJilbHaAeZIjqLyyRZf7GxRBGpWIGG840zwksj
iiHRPZtDubT4+fvjyBWdSJjq6qADEIll2Ipz/IGLASkDDVEcIErHZ3c99w6F5X9b
DZM+gFdGiEFh2B9dqndRG4uw0F7V97W4/tcLsSky9vhdtrrtarKO34srRGbTUwMn
SspSvv0fxaV9TIvQaJS4UiKPkCVUxyg1gi0hGNVdpZWQ0jpk5EP/QQM6mgM5pCjq
JEJwg7WTedLfK7tVXHEyRlDWNoD3nQitXRg3DPOajkz5GNFadMKyygUEJ87ANfYg
UgkhPGg5YY4/+SDtEpBBree87TmKLBghEDMSV2zS4XheJa0Uc/Io+IZsi9imnYB6
ZJzooh6wXB3Qw3MQQJVvbUNwBv/nsWY1B/aolS8oybEecCMyk2lpuZElM8XBDXZd
4rW1fhcDWsD1+SoqUzZ1WW6RqT5IF3CZ+LngNyI5Z/kU4vD1KwOX5oAP/h014ZQc
PL4beC/WKYWBjovnKz9Rrl60xBR9AmsmqMrpCKOkRxGX8/OOqYIgjkkzgkJ7bVmd
D88y4oR2gzwPNN/2nxhVZ5xlB5kcbziD/wlpsTStdElb1l9t8fD69KV8SOl3rXPa
JfafRgPWt2xqH41IVBMSby8W3k1gx5oi2GkwSBQ8CTxYUa973tk7ii12+n+4o3Qx
Bx19n+MCGw1riTEzhFX45MnB+mPBC17x9whVQOXr8ATGFEkVJNORKuxN5pxERkxo
pPY/0/iXTOupvmObYjLtaK7ybPOA7gI0QmbZ45u5kRMJRG2A20S6uuxFcIc4MSOz
Q+w398fVPQlfi9DRtMJMFhSUYOPT5s6IM1jVl9Q2mXmftKaQwahi157mMncwjo8Y
LvtgWbIOyDzeJ8qT75Sxz/w69C/bKVgs+e3C5VohiwONyi6zrRR7v9l60wl1AsLT
5Nav7xrC28d4QM86LTev/aLm3B02TZrLZJCqqyFO6c4hdvv0F2hHsUhti2fvz7yQ
/sE7RIlwZmtZixSp3nx0cwjWsHAcUzDSwlEi4+0hUuOIHwTvjtsQvtu2Xazsqp1N
oZQvetxpNAelryN9fW/BkL+hc2ttnN/aC3FgfnthtaJBl5Cqc8UXoi9QvdXOX3/e
b+HQO+rW10JUq4XLc5QYRuKy6iHTqux9QCXR92kigBJ+NL+Z83LBHxuNS9ArrTOb
kNDiGqnQaHTo8kMVKXbBZs8xWWUXAf9qHlMZLMmSa/UKqX9TiseG6myyBD1CPxvc
SoAxOkHt55z1frBDkI3pyEt2208z/xASkyrPpnMSHZd25Qel31BcCnb5AirRZvEg
MAeRRWn2iTitYqWBAGgqTqsaGnN4TL2ZcHpXqT4ae3kgjXGYyIQZJJzaX0Ec7/0M
yf/raArvfxv1JSH5JtJX78a+WSaJLprAWCcM+t/wmW1vHtE29QtKnbotOf0UF3I/
0JSNaBPfEEid9OxdPbkOygDmv15PklR3he2Rm7HASfJyfGE6fKAiS9VKrfIEa5/6
Q0an9gsubiDaELlITZu9MGhEBrA08NxmEhYU62TWheAlWAOwtjKM0V5njcOZbrEp
Sspigq+Re5ScDu4JmZAHa5+osCJJUsjXJprubyZXWOcqrozd4mSyyJ9+V57oynJe
lrn4eQI2kmV6IV1R8+S4DLTPo4klsY8q05o+9HC1M1UIy9knKOJx/jWW7M/wU3NG
1XNDzy5qpHG5lEGSs/2laM7GRktUkxptLzOH8Rw8x0WQRlM1yTu9+PlEycopkOcT
eZ5AFdbDuFVOzGRTjalUIJLIdGB2gYvqkLNQKyXmp7QddcumSXTId/NdXZb6dwxc
FR6Rrbgy0WaBQdEPpGcdoErapmDSObQ6IyuIJx1yT7k5mWYICsFP4xr0kmwWtPX7
HMj1aRug/19yY7yB/sj4HLj9AwHSgDyCzZkHbQWYaUU8qySasV0+9xilwUycpTik
u2lnNpRzH1ybffjFK8Wwne772xGpdSc08T+ZRM2nVQNXeHMRbyQf1VKg+E/R1nOR
ASsVLA9QLTreKeM4r/vCZRxF8kKpEOqrjMvaQ/ADE4DDZnrwqt4l2w4nnvsw6//L
e2juf+sazpaUCQnG5Hz0m72gmgFF6G1/HzRIMjvy1afW7Ik2y2KFpUN9lX7JYPRS
N1NxfIoW5blJia1EvnpGvgHQF5zsOfOtp4/s/u7Eppjh2gNEvf9sWDiQ8A3TkF+N
iLOns9uQkkPDhStofZAMfLFsqCoEuem45+y/taid8MlLPkacVuDiXCuGM2Tqe17d
V2UrtwzsUFZojBuYdjOy2b7/L4u1Xv8e6r1x/P48Wh4iE3Kiog5GSlhxrx4NltzY
WoDfv1zugG7DPfybyPCWqmswgnbcL1f5cGHdUQYqoOcykp3q0J7QvvR+J6Ot8r6I
JIjjzMisElAQDJd7B2hIALvnxBfny7TG2FzSvmLgusO5bN/ah13fRT/tXMrOh+eV
Pn6eDqrPU5ZDwPA1q8Lt7Liz/DRzcj2EvV9eCdvFwlRZivoVw/sCL1qfkQ6oXcZL
evC5x+BIEIdrVqggbLigMRftjXv/IrxcUx4lsuJzsUylhdBaOqeZ2d1RIyj0AmsH
aGGgs7H7WHy0zFdBMz1tfUS8FMjmWSHHtKjui7ykesu+RuCg0kk7j1dFqDNprQeb
xaqC+K7p3bBCEGhA1JINeyivuSn+574AgBVzeG+VsINkfZRmEq4g1F/FK2eRMSoM
rH3zqq5a+EvrOrExYy9GZlgFm/2Un4NLR98xNrlla04QfIzmlqKQmxIhcEnphJtZ
EgEFS+BX4J/Tx3506rkgCdpH8RRO465P9+rx20buQmkLs5U39DYyLreJLM9zD/Lj
oZz16x4zOYoyHFlvjVDUTXP7Xj734zSm/g5hAfscV7hsCLNZhnpB+H67d4UOnBgl
klVIb4cqYsa2OKU04iadc/66ubEnsfgOKFU59W3pbCjiE8C/C2Rk7EsWTKENLMKq
lWemQ7FxGLvcBYO/W4vN0g==
`protect END_PROTECTED
