`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8XOt+jB7IFZsE+hWhERcltaXxwkis1x1sQtLd1WWhvNXnV5rAxBVJnNenkvzz+w3
01mXiVMb/bPkJ3uCBcY4UJGImMfyKdvrE8WxqFC6Iu87ARJPBg5RkNCFFJMo+Kvr
vNNOtYqubnzTRTPozVb9Zo39RiYJacattdaBtBGHfiL1rk/5P7XDNr0dF0OgI5kJ
/oabsU2unn/B6pMET1x0GvsoxIj7363VhslsShOydSHWGovHLH31dkQ62b/b1ZRB
KkAKvF7o7b0NqtiPYKbjO2aim7xNpCLJ9BVQQ7VO6usoBpe2IZR9QSQ7eylTjJXN
BGLbR/4/MBBniv8GdobnuzlKfp1QGKGFC0BvDiayJgSl8z/ZXuQGg1RIdDsA+Tzg
JTLpuzNoD5lfswGpCfP8UqZUmnoVI+tb1BZD0VAZMd5gPHonJzkIRUhdT6EcFiYX
J/nmkrGC2bMJZtXIbiiyWG0y1mu2UtSZ+x7rdq8hI7Jg4Ry9GFqW3Ps/98KM+jnw
BsPMK0OU2qx2HzDBDHZnzEd/0qxfpQSCCgtwwgqC4I78AHvHDmPZuDpSzZZQq5wq
0AcC7mVuTZ2vVY1AMWHZR3+URccgoa2gAxmCVCJIm848UFegJmIhpPFZCMybByHP
LxcIsl9tmhga1x8oCwWIhBALXqUjGYakF0MYA2M5ISjMfENs0RGqiPJHM2+nVq01
YbVyV7pJuFYN6msKVXaN+gFijF3k5KRZkwv9SUFq8hdtxv+DAgVyxd0lrNTnQw0M
6BRIajxh1lxYIGyunttaPhoGOnf1cYuzbLqB3KE41cjR5KwJ0iY5nNQlmvHzj5uT
`protect END_PROTECTED
