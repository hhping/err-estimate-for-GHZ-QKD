`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F9VpM/0USPpZmR2nLbAukoe3wKLni7lOBg3L00bqZYuu5TkyibUAK7IFeBGfAfLp
mGCLXnNl26O2RPNA2TJvTzez26sBUkEmzWMSrcvQgAAbCvRGG+0uBp+gYeh7cbUL
xFzyJpM3XiD1oWhki9m9EL9XbibR8A2GwvUAjgLwjafp4yxBgUlz1ra2+HeVEirO
/hbfirEUdahTCGMEE+uOfOJHykDy10d8nl+Le8Ht30IfULfViMIRkgtP2GW8ii8M
SVvNn51u0zUg8lTBdyEjHY0F3NuAVG3lqE2iS1F68ReQ42Yko7h+0ygAFAyD4NYe
IlSKxI1q2FfsmtuIY7YHZt8TEardu/ks2QRcBr4Sj38BRXn5rSnVe5+Q5HEX8Hxh
0uQn4Dqbevl29t818/xB1ts6TYTKQU8wer/NFxzg08s=
`protect END_PROTECTED
