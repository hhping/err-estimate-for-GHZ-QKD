`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U0SQL2kxZZbZQEDZ5ifhSVOJutTEq4DRRkR3ESnIonVAZpBkP9luECwmg4cbjGHF
nXHhR3s1Kym7S/i9GaHx4sJoKgef6sX5TwrmLRwJwgB7NNQSUDlpgtnLsWS7j30O
xwC/1lndd07qHzz6hfmR5Mg5SZku4HhVFCZBgVKy2ANyaZ6qTPpmFgStvU0ayRTi
3P3EGa/8lM6NGadTu3Gw+TO44OeLJUYdNsgtiumRL8tgzqWYfZF6AeZXuJlP0gu3
TK1wsJnvxvqT4Uk4ARMzH64X8v7u8NEn6t+TAHl1kTNHeAKEs/7ngAPjkkN2kytx
9EAVZaHmPv1XXPPgw4DWVi2YzetKcKrb0xqWNhRjvWBWPvLW+DtJDtaJMoYmmRsD
K2Y6UcKglzhIF3tAjiu7kJAMDOGiDWGxnDO/ZIftKKW3LQpBp92ocBFLghrUxQWz
eaZ+0Ust5xzbh4kDylKjpJok9B+mkZx6gagTMLDRncQANfzqmsGDoOEz83wWfCfF
MgePRXUENKr583m3J3zGtOreYexu4PEWdIPtsy1hZO+bkeiVzLz7ymko7Wq8y48/
9xGGD5Y/t5btDUTIViyrlA==
`protect END_PROTECTED
