`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tbO8p/yvK+5d3jy39pqRpv8GJpvRKUrZTyLBql/v5l1p2glUwWpkS3qmiVqp/vPB
2Xo3yGYZJ038ldtnYLQQ/fzRkD0O7Ke3VezPtV8uZJl0OaDvAXKtdyPqUIQMroxs
yaZ6UWPc/pVWe8GT3iPOPRmLRviodEUujNoaaPZv81iOAblgUVRBniACZk+oCcdl
q0+DCpX2++Y8fKmhkzyzCDee2AFgtpy97CzUmPfb/12r6E2lVidLpBbFz592QXGC
wA64rh0WM7TGUu4gsF6OhdSH+wtWPZLTMBwy0UVirklnWq63Stp6pGJSDe3oQoPr
+o4Omlhb4L6xEaXyXsNgnAsz6l2ubKnu6Yt8uNclvH6/jyDxLqrtJP+/NMeuwvTg
5Xg1ImmwGx59hm6RdEtWhFRXQgT7InkAE3cSmS9+KKATKt3YrJu3xIKRkXjOkwc5
oN9ms2HCSRp0HP/E2FwJGYgrNggErTJbhYmu1rg92Ku2DL2F6xl6z3ksx4I4wQkG
Innna8I6Qc4ukhA3i38Qcv0Lxv4AM+wu8gYP3xonfLq5Nkk94E2Y7IyVjpiNgUJO
FUCtnvW5zgItEn2yZDb5A+AE66wrs9JEVYo+1LS8bgO7pxovFo8Kp+KITtBDwCEH
pzG3livlD86GQvm/Geyin8fI20ff75AYCXI18bsMH6e6shWkvXHaJjYnA6qnVecF
Hhuz5qqmTpA5Red+QWGUnKoc/3D7YLgA62uRbTqW3GCuWgaV3A1bgUuFwedHq+xs
GV0YLqc7raTyVqiG9o7Jz/5TgERWImXUHXpIvEJsR9f3tlsz/snUkjjgUCExT6yF
w/J68mPdD1FW+RVi6Au9XagotbaFRs/i3JxKJib22p6K5yUWZkiimdzsxsxq+V4D
L6DLWr9sZlND/HCwLCHH0CzROx4IOAme3Tf5DXAfZHpvhmSmvWk3k0bTrtbuEnxv
X3Na199Ck5DpLQj/OnFtnpqx5i5CkeO+ghNqWmgYND9pzC+6frmhDrVbR41F4wZo
Nfl0SmoO2wHxOSgBml4e+SZYPWajRwLoCGqimf+6IOfnGRMV3NUgchRH+STRCvIT
enfZiBLccwuBWJAj5MyWbZTqpJyBPvPHwibwDssv6sjhAFZmTV0gUn+d1jpICAZ+
WqE5UvhKHeS7c1aoLS7ox2BgXGaRQF64aRZEnney481dRfJ26kYiC2+4oPg4jFQY
cyqEw388B+KPZ5DiAxMXCprfyxK3+VqgsV4jGASH2kugmDVtO2aGnZgntYCYHhCh
iEJF/Ldu1dpsxI6/J/eOQsZec3Tl381fmpAR/zOnQgIyE0sQQdqfnoF9USz6fwqZ
RgJYu1ZKc+8nL+fqrNG4A1OyT7s96hN6Hi4kwtiKGwhJXV+yQkJGwN16B9pDX2Pc
50d/J5+KeHY2Juv9aFJwmuwoyRAY6IddExAZ4lT/iCmEBoHbvtdmJKche1ow7r3z
EZrLuOXho//0lM103Utr1apMCVIK+OyXP27omYvd2SXweT82XTZTF66N2FL1LIjw
XGEqCYH1G4jb6vxsuQH6S4NTKc6iWSho0WfBucRraLJqb9YwG9pn/VEnVt97KvhB
XFHcmvECO9770f/CdwzLJHeQIByVvfJvznvAjEORcYKjSHOIOI5y1PDnjdD+FsiR
sS+I1yF9ttZX0DtMZ7AA5DTQVsG8K45hp4lp//5QGwJJ3m9BC1dldsBSy7nLE+2A
iu3piVCw2GNswZz6n/qwdTpM0v02hohUKWHHcm4iTNT/XCjMODFiDVBAqrc7h2Fx
RjvCIHRPtkV5wg22UJ8FosqiuspbA90EfYPjNiMthAMcmNK6KNzF9oFnlXswcgY6
RGJwkYnhMRO6guahrTidVCGspBvSdHV6GJ1+vvUgEEceJf77z5OuXl1RVxjPNKu4
EX2CwjkQO25/7cf56g0zsK+j/aS9XO10gReCrnowHh6b7T9pX10bZnY6ZtpKX15F
djAmdb/UUzpf0/1OzQgn3nBrEhAtG8Q7PM9GWjhik82A8XMJP6tWsvlhdmfKMaOy
BFCVeC2QDkVVxYTtGNHDtswT8JYGxBPePIt2zFkbKd3T5kRZvDcUkenmjj4YDf+b
969/aY2zwWUMaV644fodkWmEQ1ei1Cp6WhJSiv4uPmMqh4/cgc8vgfTk6t1BrrjT
v/8D5AKGMOI6eOeI1Wn79E3DdyY+H76OJFcDUMoESewXAZHAxme09gkMfrT2iTKm
vtSXtyNRuAsw7bBV/c5Al39lGqwsxnbi7OIzJTM7gkDs8Y9l7rSqP8VYtCgUiPu7
pUNeYg62kwyt0f+/x2JkF5mS36l8iSj34nA9uEZou5jGXZjQ0xSaC4Fl4188lT+m
/IOvCjoRoUFDNfYIumhsuHJeSfb0q2vqc3hoX+7cGbsaHnX1iZO4wX0kZv4GdFIM
lXHqx3bELtimuPWNe6Tt9q024CqhQdouYc4hA08WoRRqyaqTo20uU7p8MBiP7DKD
w0zJQ9CJT2Vp/NFC5Mn9UFfx+PvxufYQRlicbcXyf2Rafh1SNuHed1iRAIsbKhkV
oGoGMps2nDgYfxG4shSOD0CckYqft25Q2jdcjsBrZpYnKG5vTJOz+utnMUjk/MKR
WQbfdYJDsh6csNGaOTEMsyK04588FzNMADUom7Y5Elx3OkAMiVwfY/g99o/YmbjY
zAiakjh7A0uTEzb+rdTD+uxbn7wgnzUhPaOYhqjJLOjENlzpTovxKFGXxCLJpIHv
Hwzg0Sy7RWOiLKt9kpJaaFgbgUhStjQopA5dU1vTVFn7WjEBKf+S+ykXGWFBTY6R
PFjv0NnBgwfXJ4yEXn2xqI7pEoWq3WOneXCtMzJ/J0Cdz7JjjtYOqbQvXvzgFWZV
eprkBVDx7zJ7nKpopTy2y6zEPhIMnSlVPJQ1kAeyBvUg41aExUvy2BKBuii3o4TJ
SOSdUkkHeLY/8FzswmFxLabEgQmm5vhOYOZVzWxluaAm5zZs3jv/nYbvdezCI9/4
2CF+KWSg0x2E/FJwk7Wn9qiGhXeYWCKwB0iw9H6lUPOj4fmOHKvFoVSQoiOeAsgk
f3cVq2cR0LVK/4sBPCrx1yYSNpt4pu6lki8FuyP3pBTMkd4H1dBSTNzX124zdjsq
hUotjEVinAYFqaoqBc6HXjh2I1PE156U13mz3eV43aqAxayLCnq9OXW5R8xQjprG
eX0DLzmZE0wCIa+qcbqRCoI9TSjjPcX9sTX4fZL2FHI4xeywrXIhusEox2p8aW8X
1MW9+cc8jg8NUMgY93NJWLIfLwoq5nHLl7CwWVvt5JES3niChnt6ukC+r7oJFx8C
pmW5CijIEcJxq7VySDOJie478lOGywbKmFTLSi+Q+jNcDKqbp2e1co2iq/ZVdIaM
+zHm6wFzcSqe7OWr3k+WHB4PqXsWXdzk+ts7ztgOVOA1GiqPaatTRS5V/jws8jFJ
gXTiNIowDYYj5PZAC/9FCID0ZQLJcc5TuoZzyiTBhdpiI3qyEsPC4bdiM/ok/VJ0
vwngzX62iQzbNO13UJrUljVGmODWG1bvt5gFjU91zV2nu9coNzf5BnlCQ+oP99Ty
fvfMvuZfSw49BPLh5kHjhhmcs6UZLXcuDBTas9U4JXQk8S2LNADBkls0Ft+y3mxr
5tT+bkrouQ2yf6clKm5UWWkoJOj7y6/ent3hrj73NTbq8d9AqGO6uN9sBYg6v8qD
JyiJ0pzsSSw1mcuNPnEl3corYpLwLirkTzojw+ltYVqNyPtSD5NmhJZloXBL0jm0
z6m/pcMqQg0Uk1yzvdH7ZNjwAP7R5EheuM90RGI2LLIl7Ot+RBNQ5u4eexvl4CCg
fngt3a0kiAIonpONX7Vk+LFQg78eCCr8WGcARFqfaMYQrJGO70kJO7jBWJU3h4wE
FmTp4FdKQcVRZEuyLtTTLNJUdr127JnOtXrNv7/rFFHjwoSiQyVWU+v9bDjzJxLY
sBEiWy9RQjUaT5COvHc1FNXUBHsobqSUWxIJiVQRhX1ASSrwmhXldI7ISeLRGpmW
fT5n+YhYSlTwfIqvlx8Tre6yd2FqObA6/jN17ivc5LUnxLJFPHcXLe/MxyKOgrjv
Ef6UfY9qLCy7W/oDAZeT/khYPPkopgN7W0i09ScaEjdCIRfM4SgPXdYIUSnu5Kvw
k+3gJBumRz4xayPD4eD6UywjKQR3nCaRsvMdAoiYo6Kzp3LNw+o+dpovwPQiqAwS
RyIA4Of+d5SlyZd2AO3sJoz1IkFzMlEhPcCcTEgjtFgwWPHc5A/wVRpzZ0t0R0Vw
2LyoWaJTXkVZpm6W9+datT5chh5b7s66MmEWRpCju1mVMmgFX/E39y9HPsQlJOun
U3gYyYON10Zk/KriYkuGR5eT+uV+7JKfPA4gniUufy0PynydOUGHouaMLM6pMVAQ
6wyE1IbHix3njrELZwLK14DYydl+0AYBJFvEZ+VXfpn5qYR209GoENUTiTZeBy0X
nZ142/CgesUu/ue7j4vJiVuG4hVpSxeoxa4qOsqufEHgadX7YiEof/sBSyGuWy7Q
OGJ7i+J2Cb+wJSD/V6rShlzh+Vo/RNfGIZbm3E8iUf5uyGeLQ7saAFxajbKph4J/
nSdAhXGOWz8LBSkckFKhItXbOPhcSW6rYG2jRcfYRsEapb08uv0ByP5aO1HfAXtT
VFAQxE4La9Pz1YaiYGdTs85xAOnkFxcWW5sO3fixHLBmnWcDAjF8ak7ZCQrDTEaB
//ziRZhWUV5Qa6YbKPNZD3wAeanVuvaKto1k/n4ZQLqGJzFOhYMwPLB0u5V7RvF7
f2qEMu7Rkp3WE1HT238d/uf0cs4ZQMcu5gj0uniXGJxLpgm+COMvbfgQ4h4CANj3
NfFVDuUOX/yjOnyF167mbjTjGAcKZ4iktJGPrygXOwCzxC83ZmmV89gzg40QBHRy
GL4vMgrnw4ZbJmGeR278BlLTNRlqrsSHrzlYMMO2ErOkq6EClcgAwyHs1XCAOLA5
UcxP+Dz4Kpe+xVfDKrTe6VY6bdtfKE63ZxDolHRlPf+anxnVfpneStWo5CSJ720x
56VJKGNY7E/xhkqNgC51pA+FS7skyJqhPG1kzrqi/Z0d5Qbbf8J3xfNarqlkCy42
8UuAm6zB+yP7z1XfJtav7pJAlRrK7teyhPusBwT5PCIO1Dc7aEu3EPqSsxU1tCtX
xXLnsr6E0+ZMpkIcGrEKlRksTlUGrT4K9/GF7JwYx0O15EtyiV6yjpEXvj9h+2Y/
mN2sjxv7dofzVXpJ8bDfbOtPBbU4rF28fW9tKrEBgxERAteM9KIc6onIw1UGCYl/
N57xB0r+3HVOiufytC5qaqFsvQg2YGt989HW7hoCoeZLf7Jv/CA+Vw2nJNtzcRN8
e+MSyrxOB8Mm9uCiQSVozIpYFgVNAZhjbELm2aCs0kpgzKMVq3Z27zJQ4tUDiSaY
sTzR9ejKi1RspUChKn85BUypLbQCycuV9CONYefB08ZSsOvuJ9McfFAtyc67S2R6
4tAw8RRvGjUGwhRv5YQSFCoTv72LAU+R0lotgX0W4DY1RHjxzKIoh4o3dmFlHSHj
y5h7783G8q093ETuVo80ewcSnhlnvjyfb0Mrf7ylOJguv+g6DTgU9/TYwfYXwZFQ
ZtWr5zB+grEUp6Z8n7x+auocYSLT5UFQLraTF7aPxEQR3Q6y5v6VMacDHiZgpHJY
E0/gBdBJsxbDrdD719gdsr5RpJ4/JQ4lZxhXhR+mLSyw60fA9+DOG7Wnz9qmtOsK
EvLtHiL273GhvI5M/3mPRY2GSjHdezsDrAgu4TZiubRe84JpWIjJFTZHFBysUAaC
GGzNnHe9Va4glBYs5chQ4GNYIYJrptq1yM+YOSZqNhGOPJ9Sj81TLSSqdPuc1Nzo
vecBYEmoBTaL9ZOCFSV88huVRUYGQdMt0wgeDdcdHVraPO18JEe2gCv0sDA/HL1b
s1JKJ5lOUi1c3wkoXBb84mpCiG8MV7ooZyT05gw0m0pu1wyn4EzEyM4jobB1TJIe
Hj4jbWrgtDdyIrOKTsGkM4h3X1Q+gMjV766buRCNFB6Y4/LtAkgMaffBtOLKjov9
mrbTGhN8ooav8oyMa8jKUn9XaPspF55Uq/+8upXOKKdO9hg3UKZ1CFIirD6PuXCF
fcjirVp6DPocprFG5LpiYhRkkxOfHhBdzj3KPbRNue9jatFBz67i9FqbEkokUtR/
mJtKv5KGbZBeABjuW8JZqlkFCXdB31GfIkle/TUEm0MH0s8b5J2ilnO9YXEvzpUW
8NDYSpMOQMbOYEoeZs+iz161AoQ3lW4O6l+nJT2cH4cpDYtDxUYrMYAvPzXikkIj
At2vttfrZ7BR55sf5tPZIcGT8+YQolRog0x9VJZP7NE4/GnR10rl7qRjuvfnWSOT
L+HhIgxH8e8J+APThTDscjZLte031udWhmoVKQ/iik38tFbDzqmMISXltHlW0TH9
0Pq8FN3Yo0Q13enfx5q+SV+7kLvJnhCFlBqTlNja+zjPV4HACKJ9QTiKeu2s4eQq
eIunwh3/0aC9WHfq3Sp72qZVVYB3sYzjwXJ5GyM/1dVXqZI44idhOEeMM9Vn4t/F
NLRdpCfg+sKsJ3fAIq2LViLeMeY7jaiiGEoGiW/gDgTQLPJ+CtkBU6V8qC1yCBVA
5zntMW8oxidDth1IBjmKyxHL9yW7/wuAmq58bABF0Fl9H8n9tTs+A0nqvKjELw1L
2Oo0hdwSmqUFNlijEmx4wsaoTRJwrrrjDkRoag+E177bKDDm6uFIh/ePSbC/l5xG
MKjErBC6t/aNDgDKaCKIWU+fzdRQNkip42AJyZefWDY1Qiddhob/v7xDPm4kIRsb
m5YTKyPgj9VWInReHXLz3+Q8Dg+wILcBwNjqCa3EJAqYln0Z+sZ+W5MbpnX5P5W9
sb9OeOQaA5/DD21QjeoPqX/i4zjNeBND14FzIl3BUjqxaINPfjTBO0Q6axD5dLWZ
8JZuC7S51U9gXva3t2xXBME/6cpwOsi+GvQgRQ+VZvA8Ew5LMt0LR7UCSqrLdWlM
oo7ffQePYX2gYCJ37y6cNOiUwNKE44SRIiPofWyC8jzuWla6p23vKyqtP8NffyWc
BmK/8t0p5ZzGHhnhGQEwHypc5lAIDu5CZb0+ynkvi9zCvGa9lmb8R2UYKKtljlBU
Y7C0IZMXW9sqcnwho/rzdesggmT05466AzpqlutV2U8AF2Jxxp/kpxUGyu1ixnsv
ucH+zrSp7XYRA7KOMLRRiMbiCUw9Wmzes2AqvEPhXRUV7OTv9m/Wk4Z8IFlJQ0dM
iwOUQmYOFGDsdXshfadMzh9TKI81CizFKcWyMZQjF4GN2lOklQ7esGEqU7L8kFD6
yzMzsHHSf9NCqVNY41wQZJi6UkJYgfFH/z5kHb26bUuKr9xP9DTMYSoL5Folny8p
IUHwn+ZmHGkIHbNpjB38xeQDxlewfnr++dlEbIqMY5nG3Dy5Zise2mpkx9XCwXyy
WLMgkyQIel9CXrl3t0Qgh1T83GgJdJ5ekZ5CZ3Pxu1ATS7m+j5fyXwrM599PW2mS
2Y2l5Ig5QYznuuCmFyX2ZUCgi718I2FoTnWzr2hNit7rt+WILzdLPMGTtZ1A4iCC
GLAvyOLbFgbnVAYXvBjv7DaJJcOx+6AZUi2MdHRTQx+AcYsgOJqNReMChxnUKwaR
Ch/Q6NlDo0F2E5ghu5y0Ei/SFwRGvMyY9BfiN2udZgNCtw6ZP315FZUpdcl2JFDq
0K3cBGnzWzlL+pE2nFm2YzQkM+UHsHY4ER97Mdj9xch+G9bNnjtJWoMRdohpEnAd
p9CX7gWRylHPEgb752kx7MZPT2FhUElFWEx56Ci4VMeaKn8TXvnRyUuP7UEg37yR
LwPrPfEXz9r34nxrftQ5CRqcJCWXDtEx4b28RqmBkmJQk6ZYu0Q/iCXbsnb9G78m
L6KlZJydKt0ao16mV/6y4qdW5dZDdiOHChsrz1Ayf0wwVvGRGL6ZbHJNrbjX4RRr
BpJfEDt7BblVCFdu3mQ1RGBIag3fewnQ0vSKzL4U+jKIF1K7eXm6pbqlgFiPzZxy
2TCqLCCJhKey7T00If8VY9gWa6ahxVtiueNSu+9ie/atStG2fNle2qFr8/MTGoBm
H4emoI1piKsYHBO3UO6x4TukqTeCENy1dvfKMLd9W9XzgrlJDzkrGHb5chDTupzZ
M8fVDJ/bxxA8cr/K2ng1uAnSk9jjbW8u4iT1a7L/u+hkbtiPqg38ZUe+qZNe88QG
qV5BhjztYqN15f/67sKg8o9CoRyuduDCBpi7xxN7Xs6EvwZs2iizzUVYj86x7XfC
fauTTFOAVw537okId/Nwtq+FlqmsfJnrBT3rMS7fPItuWiB3TuTLvLy+whSXxprV
rvfWLggxKGy+81bGg2DXc5Nm1OazNal8BA2gMGJl3sjROhNE1VlkGtdIROgjp6yd
fzUYz/G58tmQkKc5RaoE8OuruqkLCMLSY4ly8JncGXcpkDlkiVQ98YimVDVEJzOh
sl/mi6uryNQmrHSHByH6DX4fu/8vJs8jmf9HynvWcETAj4WkGGz1gfysRT9lhy3A
vVqEHhVFyZ/Ilo/wuIVO2zvmkypSSTINiDrtTOU6xNTv34oULZ/r8cDmtsKw9lbr
ct4p0QAfw5dm8YeRp/5mvDXMNNw/IuloXzGi69+RJZATxdqMSBvtrAdFzn5Tls9e
eBtCDBdkyhW7IhImZSO1+Xhxb+qRGXaKkNiH2I4FCF4q2Y+IxwpsqlkpCYrwjnxG
emstzS/wO1XWR9/3nWwZgaEJz98xVCFa0N/xTZK8MgBq9Z9tnszAdT2bIrs0tSNv
F+fIP0fMxB2n1zOsOT1Vs0aH3tT0HZmA025N2NT6EG99pVVOIoBVDusLGLXQklpE
hCc/XZHrJnSSDQIBbl5bgg6SYqytHUus6N4uDpzhaYXI1rBAEwwwO7DmRwIgnc3C
88DdtykEm8jMe0vbx/PO+U3jno/ZSvj0H1f/poJt/IzP1zc0CgPEDDTnFm4ydRtX
Rln1Hga4S/NMm0KazXBlzLUR6UG9JOGruWpJ1r88gLgZQSXXztv6QbmBHM+2Jq9/
fwy5SNKTPstlnwXLD0r7U38vzIXBhqBnLITRbk+PBj3VRTu/p8l7XHAYhTQRuDEy
1TkVHqb6W+BkhxBJND05hExvUIqJ5TbNeCnb5m0S4CVQhw17jBs2shejgUny4Kya
jQbYXZjNEj1h16QMFvJsjMUW7bodwW+W8yD89zpp0BazcSBXl2K3dmRez/rQWRKD
RziFIVL3jrrnzvexEIQjpJBGpGrffsVQYzi/4EtdLZvlp3R2m3RMEA4g/WI9/xtM
m886pwItq5GZdxa9LrfyhyPRzhUoQHxr1sVm7fkliLHv38R9TtolX6+SpxmZXVHX
5qg+lxWC05KuPc4v0yNRYBvQukAnyxCp3xexoOyN2cEko9jf7m5llOSQETfDLevB
vDMbd7ZgU/KJvtcxzgnHTUwyMamfJeP3r/aY1bZEi4XfxXq87H3Pe97CSuZYx/e/
G5yxbGU4X6Gi9fPu9PEZVMnJ56wkZsQVl48wNfe2Vm+l0Xgr68Q9M/7WpjCIJtm+
b/puPvC8QHt0USbl/QC3VEUMxHZaGEqh/YLEDalzhV5E//8A0pp8j6wHfVjhGqDS
G+jBbmDU0brZlksSEsk1Mg5o8hYLdBYG3dxb80RSwOFlCHm9bftwoO5YGQOsJvf9
xT+5a9ERvFbVYLCNb6tsFIQaf4pd1rnZHgPapz79tuPA8Gjx7z+C5BEyj3YYGNyS
Hm3BTz8YfM2vkP6L+cYtFZt3yXaxHgD0RK3OoJB2nj4TpqOGEMA/r/epZH9APHad
ePto5mADMw5ukQUrYK3RgFAuC/veJPVSjUvvlv+jH8BJYPT+4+/cPmhh3rPrmhFY
Kit6dqWXdFMXcqnfYUP1YMNFobpJl6fdxSLv3+GdaIDKbTDrXPvPCsyS7Zj1yH6y
dwXYxMEg4gLpxNbzsrumI/+yFsrhgBYy5WEpJOj8Pod5XbXIFnR6lWE4JgrWHGVZ
CyNvTBS0JI14rTfC+NcrAT0ft1zsd2B99PP4DfBmpaAtMLkgAhUseWrjczYd/i3j
pd3yhJS9NjI10Ru2RqFEh2ZlBchtELUtrkH4u91AEBpePtuJAjSnMt/nUq7OC7kr
xSn0I9tEZi2jjuLogeYOSgJ8PgiRivudfh38FWcaoX7FK/wblb2wf1XDxsXZu9Mw
T7OFlZ0fy3c7vw11vvxZCOqRVXPkLuSjlft2h0BEsbroF9M6qE2581/XFPuHdrul
Kinn8Pxo9ByiwRmbdDfZATgjSUZUCTMEmCUv9lgfKNPw0PKKzH9WzQXR8FKk0PmM
u5mWBQkyFtag4OS6QNrJ2ZXxrnmtFQ5ohHkZdq2brS4yTR+tVK4ni2vC+cNHL5B9
aPkbkJBxmsG+YRnQQLFYsI2V59bXXrolF2a6eVlL36uL6kNgD7v5BRjvUILgTCYe
OORPlkRM+GIw96a+YjK7XInS5eM2DkErgp4WDNLoz+z6bae03rJNp+X3r71Wvwmg
YTq93qpPase8Oz2uo2I0kTSKcVSBpg4NPDEA9V0mhryac8uhQI/N/7CGtXWedYhj
e6xM9okaDsL4XfLsnwWXX4Ktbj5NpcLYfHP+1a+fa9nDr55XY2SoYSP5FfHjkHsE
IRrj9FEHcdQfLCUkr6Ae0iZ6K091vEnFvLN+FZNp8t+Fek+vA5rprBR/a5upuZm0
8ibBAu3wNMxNQODir1G/GUp35/zWP1h+Vd9/NT9j1rkX4TMgS3YkXMVAypv0n7V6
nQ9BLLHvcQl1SoPr8Z0vB5ljI0gt9fYf5G3Yc8VbpfRCjFE1qrp/cScCIjmu4zqJ
Rk5vRPKNi58YphbwMhTXf/GKtldFedCR9C6Fl7hIjsYpgQQGevc7TWSS8TBJIjA1
LQZ2WD+ygmim49i5dB7epo7tvQ8Pd9Sbs5AdxxCtuejbxJEplO1oUkWg57aXbujb
71/kL24PBlyVf+jxtRfKqQw2jCtkyGOjrp/CpUsLt4tvhSluxlb0bQROHmmPPIO3
+hUpnKSjx5hnwW+zj3lacBNMOPhPBuxbl+RxmNMpLoHAz2Wswm/XuwsMz5vGTlZX
an7L6XFeh/RHtvjxnn35UVaa5ELt4KnA9Q4rpgH/+yuq+8YEioCIlOIPBII6HeTK
LMoGUrArA6SXfOBicsWMcpzzxpPN+JJkwwZ5RJfZO1C/0akHpjtmQpbFRWkRqTef
2o6zJCdBWQVI0pdqTn5vmQHEokLCSJRD2McOG8/ANRE9a++a4gP2ieTNjZ/LOcjA
FCBUwVrDQXVlJjU49bhVa3aCnFWRnIHMfTLaeIcCygB1zk0mBA/569bTIQAfnUDN
RqgKdWdVTOGxhMZz3ZApSR1e622kfV/74B/rg6hjI3BKwjBSiQWKbbn7StJSayok
2Al29yajSfQcS1m3bfvw3sTfEjpvH5FI3/s3/o3Dp7fHj0G0s915C6ZJBRxh2GQd
CXve2u3HmpzxHEjEtnbI93oN1hh5xrMGbiMFaCBzjcXoEKIeMOZgf+qhDZlKOa8h
TjcwGROkCXxf9cIKEN0KEjLulatvC1f4yGxSvLIJwhVB8csGnzdVgY0qAvEX4K//
y4dMqjOqiZqLYXXpTXYyP457W9FVMRfhxBNcuZDiZqbQJIqLutOyWA5XwH4cvy8a
zo3fct0t/dEjQgJDv8pPdM55KfPjXTu3hV2v3LiAyMGOzNBtE9baC01F2vZBRWh3
W/qu5RFSV4qK9wPfS3nFEULP5q7BemDuxBsJMRllSOSCOUmu1MRRy4nloXm0Lcze
wlAGJAkF+vxy8UV/Y4ZQ7kR0UP5UTG305ML2wpuStNQclV1psG0esRZEkY2jMMmU
XAvPK3QeRI2omS65F14OFgxA8EKm9zR03hI0qVROsX2A9EvwXttkgwDIrtF1M/nV
PKt2FyvSWM3AU/ay2Qwf4i20y+k6a2OGi6A7ofoTr9aUF8r6cY3GOxUHUjWVu1Mh
1Ty8hfLRmhcuwCzFTkpt1WMfASRHLp76EjgOMab6GTdzcMFlIETHXPzXGv8QoG1N
NfR9TNKkavYGJ74lJN3Qe6Y5JPVMx98t4TD0a6AlobM3km6skQ7e5OTD9EbPDVGO
rnoMUMegLWUvJY0lxoYESByp1kf+7ytd0sf6mK7w+po96fZHsZdlJzTwNHU45kcl
JhO9d7YcBSg6jM2R+qRAM8DcnhJcyIEasDCBf22JYQqFkGph76E46El+GCNu3vN2
SLTxPC//vEist0rRCfQgBhWJsBBvcVFmsgOKmSVwOkrx9XGZb/xY0xYzJ3yIsEbE
uvcMWeK0fPcpMBibENNGHgsvBJg2uYCbHxRAglWKlJGci7RW3iSVlVHQ1A71zmhR
S+RL+Y3ZSXYBNakmEf/qciu+XUNmjh0vEpSDADWqD6xJBVnAK+eyI2GeZr37uaV2
1WPTSe+nYs4uE/W7G1YS8mpWVpgy0tEcOPGcYJpW6sil8KkFsA/GPsA0LqRCWTpB
RYZtaaGJZgWydZM9yplPZDb+XmTNs9J/nSCvvSL8ctpaly0B5qepPgH2XYjlsRuT
r4dcLMqgqVQDg8NBDp6liiq4bZJ/dnCWUJ8VOK/kj595oiYgE/hGV4uBfeY/gpkG
lXESUk8YtGNfHgs31JCb0rb31fPkaa+vEW37/Nqs84jI2x9qLeRGHC0ptwuCwDiq
8hYOmuyik504uDekJtnicHz1pLEpDj8CHGot5l/2r3Vy/vrFsKn7JDYgny3Y3XTt
u2FwEbbqpOLpCgU0rBzLfRQEFIe0w0n/PHv7PZFenwBLyWjwPrOkLFospleJH6E+
OJB90sUQp7CsBtSnj8AmBpTUN4CsAMMgKcPwYlYrdYG4bZGy89eHBtkUJaRdfNH4
ih4AnSUFweO476cAq7P9zXB9tnxk28uvWXFXfWJi0mo1RB7m+MD2rngMjGSXlKz5
UjEHsBQpgUQYHft8CldKx8+Tal++a8fyhCZn2GaXecwP4RL+9738bfUNM5ME2fxi
xVzRV9/X6iRSr7KyIHKkac2Gv0htYJL21m2vvbivs9PwY+M48YVl0JzRbVdbWRnA
7AnGPoGkP28gADxO1wfiANagjhkjdun2VL//4F9sgklIzAtCI6yQTxp4xI0YwmFO
u7A670yaJ5JgieLPVQSMwj76uKmrrtGkYs2RHGUZdLQqQkC/IM6dTnQfTv7LGuTA
c4+5qO7dd18G8HefO6SrISMCuWYR3c5vPmBWiPWdb+cdxG+ASTVOeX7UktjHQzm7
Io2/P/V7PgIQfOMCQ2eaMcVYxx8tXDjQWxiNY+VBHz/0/S8nmfBKosq0GCvZVCH0
J9eP98ySNXpOGvx0GpVRcBPo8O7g2cntT0ScLykk118Jw6X65DeC3xh0hSPvkfrG
5VE5ufdtBMU6Pezg2viJOT6k8WEMyYMJ0BK64RmgW+hWNxQfRn3erlRn7NVC7EfH
hFIaODsyIzMGsgjguxbGjW9lsGwSrH5pRS6/ks0GMXdv54sgPHTH+TlketFXuaeE
iBQcBjHL/4G/V8kKb+8LuBL9sPOaFT3Dpv6E30IcUc5xJsa46gmUY9SfzhXjsAQ+
3bb4BKNDhnIBtWY8TnQPmZhlOhi20HludBBvlLJiyxWhUSkY8hH03s/UFlVZX55v
0B79gNIaI6ZJGv3EFFuW/HPgGgxVncvbApipz1ngOppueYG07nTz14AQsGwOKZq/
cfUh3Ekb/kVd7tITxtkBg4bXg3X2Njsv6KrEfUdko28yEuERm98Hx7ENhBORYBWE
fsBH+Vdyq7TgtiphYyByBt2uBt6ouQLxNjBPSvLCNMI7tS25RqRT64UgjRNdDJBy
En5hDBia+5XY1SM3Yv52RFd/GNa1DGzoMbtBdV9XXBfLSfLNe+90MMnPZ3bnauIG
JCkQS5Izs5D3zNqHywtZmYGa8D/3Fn7fl2OnoiuIZO/kzBNWyF88EWaIhcqPLv/u
hWjggtn8SZ4Y1Xn2dDq6W6m5HZmtpeUHMEqiDg0siDqhstlXW+dSECjdR/UeQJ3h
yJW+1pGRsz68nwVXRfi4NjNKI4agh9U2zb/6COU3rK8YQiVvgd6tT/ckmoNuPI9a
VUqR1xcdvdoh0QzS6UEu5ARbUz1C+V66waX9J9XC1bmX2vFSqJMd6SyPvAhGU15C
9Feqju39pSbhD3LjjQfVpeGRjaRaE8MgRt6zuLCYHP1L9uuItHubCdSF6CnlNbFL
XtXIj+9NpCut7cGITnZGyl6zaNpeWGdfkBW4kEpQoS4FZisspLOe2OYuK8vqwoXV
ToP0i8J3Bga2zlBDDv2rDMA9D7sklUfxOAGuib4aED1/0NFhTTq2N+6woY/DQ4L6
O/3zZVCyXR+NzWlqQy2ntvz+9ANJtQ7A9UXA49YWFCINcFErkgYdLBi6vPOjGFhd
gTOzD1x/oesIVto0EeIoCQJIdL5Av9BeEg9kv3+jAmbLkIbmbVr+2CmeptLyNUDp
4ocpH35mQMMpncJso5r0Rncl9QvR9kPzAaJcZEJNwxLkebSVTgR9f+opbpHPf95/
8aj6hwhqA2eNYEG8TDFDbQgLy2DP8Qv8pmAKSUHlWNpYN3wh9fuxzcEfjkARp883
gNbp4uHMp0ASKTEkDNdiWueQUNs2zGNa17w/NlDnKSjP/x8i4Ga8KVZ/Kx7hyz1j
2j5UfiwpJ64NzQTT1x9O64X4oZMFcYP7cnlzt3EM2yAVXPCGx9AzkxTQgXfYn++2
fVMuusgMODH+OrkWKnWHNOxtTaXb0Bbqu6J7xsvtQB6x7rEiu9mKn/Tj7esrZKz4
tAAXmvGeh+JBaLQLUKkgrCoGkhywcFchfUwszBuDHte/a04S4IybAmwdbz8IFJQY
r6hwgHlbevBdeGaNi13nZ+5gusF1whJsNFQZ+0UJv7EunxDj6M3oTQHDwv6Bz5LF
zD3Fedq2CvB1aQk88NXMwzZhDmUsSprFaKITojaV5ymC+rtyT8+OaV3OqYK+1fbW
bOBUOmSnkyla1+g/FcpLQr2azUhbpAPkzrozLrLG9wjDvlgF2Tn/tyNB0aVtnCZt
K47FChn3sO6J74kWcVygl7HgsKv3RONZbzLtYZclv51Ml62GCzfi8VHJ2sns/Bgq
V1NHzj9/JVbhu1xAqX+sXG7eJDs+perE/rjEDKfFHX+B8M8qpxbJXfapdGbMZVQp
uAYTKvZ2vyX0qrlaTBbcznd6MObdhGW5B2eEcGy7ZU+gH63hPTo19qpUIIAzr3vf
bEJFEcaBrU3KOzsrSeiBwq6OjQkJXJHIshQEtO+Z+vRDQvWmWMVAr/V+vCF8dfBS
WjsW2riwDkEmwUxAaLbuJajM/pltDc5PchWfRhHAyc5ok9WBvzu8wc7jkuqOjUwV
aQ3Kx+/DhfE4+tBkaPPYcCeuZ70DtS2120Xu6fUFZsSC8xmwD4O2VnP9fDDt/79t
YF4poC+7RpO54qnYtlSkK413WadgJvvg13CFw3qlqaRyOeOibWsUPQz14tj8Bc8H
rAeF2VaoQoBStD0f4AWpO/R+tyDOH9WMMmaSs+VxQ6iVntFMAWhiz+g2G1QEmeYI
qduw65t9AKl+12rWh9pm61pxQqllVCz+XNoHN9wLCPGB1LcBUd9edp2891gqOLWx
/pLgKYP+h7cdm5oXaK/mjJHKGJtS8MoQDeVpNeiQrTKc19+kbEHvPp5jPHiQi42+
yUueTlCBsFGtLB/o6b8OA1eolj8Ogg5cCUPc4fMuLQ9hYPJj++6jPO5chZKj4RNV
LuI14ta/lovXzo6qwASaMKghIOxpt0TUpQ1hClM3eGLzwJAROquqX2pqWoDHjwZO
RpcqCFCqlTqK3mpmJGmIp9WxPf2X0k/s9RrV6QXxaDvS6RgxzCK9fBmvmUondaNL
GPIzL97wjL34+ndLkBpCN4JujQcxtgMwnLvO3TGpdBZf5ab+6dimC6yMqApt9tbS
BvOvVavzVRpkM5z2GskB0oiapLRMWe2jBAu4vTPE7a9LO5wIh0Esbo7s4w+WAx6t
Y9MdxIYMm00BPpGWRvM1DPVme6LaWFG6iCpcVLuB4EEw4i9zR/hM10iCtMTrvUV6
s13gdJVw2qm+zWEx4b9nxveJY2fYFSoJGKIzmalgKqTZ5j+ZAKsPmtydYpqUgzq5
5IuEv6pDlmsLIFNen6qUC9Ffere6qmr9Oi/baRumYFbv0RcxWsSZ/MhaZjdF977x
QZ0X6wtJsfrIxcVisPgI4oM9u8nRyKlPEPe8l6SVa9CeuEgtDBrBnL5pgDnF12Ya
0bBTqhnr4YFoZeWJ7kGs2A7JZ2H/KlRjOi3l1RQWJPgpnlgQs3P5ZvnC91AXxBRC
LSRkC+GhBQVlnP7lvM0Z3FazCoVP6r1OycUOJpzByuGyxNjCiSxqJGZ8YLcD3ET7
2nGJsafFFY6htV6XYwc8p7LZ2KSIokgdPUg6NJO0tnsq3SUY93t6nROCdLma79z+
7Kr6Nc2lf5mE71LpIqKX9A+EXe1s+1TaLkMXzsV+AyK4iKOslWe3dk5PabfNLAID
v7vK0Dy6qvDBp4nzMJ6o8/RX2zyWXZo7bSIeHxG6MMnXH4PTKbxdCn0q5L9cGNR4
G3xEin7pvpHV22OOU/HUpym9EomJVlPC65IWHqbM5NTwfZcKUsGD/kCweMEmr8X7
qdf5Pq0gvEdp0Mnk+DzD3IIDD3ihgSiRwEYhBUWnVJFTIxSzHRKkGRSyq5h2AZtW
xPqABIuEXN4jJacVJO5D5uaere5xO+n6o49xMrWMN7imkNink83zLBHJRHLbTM3h
IfCHoLAACAcJh5YOKa+ELZByFeb9ufJNfa8O8RJ4djpowAVNOrR32V1Trky3YP9Z
SL61QfUz2Q7iF6HyIwMKKArsA3bNTNbRufgQHlqp7ZeRVGIvsAZl/7AnebGjyZjH
YpWDswQnOEj1671YXN7ZtkSvjYEJXxFbpFz2KHTrKcbcxvcI+2bcEmkeORgjATKO
NEykkGrYzTO3lI1wmqssT3G/gPKoRGfH2RuyMmPIFrntDvqIUmIdqBlqRX+wXxXV
/c5kyQDHTht8oduhrQfN0wj4hr21BSUHF56JmdOm63vZsnnaAzwcjaUkwzX7/bFW
uGzta0D4MnS19+ElQb2oQu9m/NgOQBBSl+7k303QicKic2GAW7fLH0uiy85nCq99
VT6RXBImOKUJJJPYWx7xZQXNkB+9UTDBiKf2xYYC4gO7+k5qsflN+YUgSF4qSY3L
EMZvfhy2FMFKgYXR2mYWbqT3tHeRfVJ74HTH0ZvzNgewI1GGelH3YlUU8ffR2Uo1
mCmUOpopO9pFypn54R+iYDdqGAc6glTzxpKG7iEB7o4NjT/7zMcEEFDSoudhNATQ
eS4h83qnJNnmMrzl5hTbjx/h5EqIy9quVg202Ach6l72PQpYMng7hRydakk3+cm5
9nDS7xS6mskWhqQeR1sTkHCicdOgJGcq+nKKV0xliiP/FSKQaVusmA+L82WcRf84
L7wVdc94OxSKzV/ljAjctWf2z/7Jnq7u8PHcuKmQe4IVIxk0Gu7aveuW6/fZ3ke+
2evl4Xn3RYGij5c5GPIuJE0GJ3KxF9TfHajX6P+oBrIyyC1HX81Wci+42WD79KXy
WSbGIamwtC8R1/pNNXGjOGuwQ/bFcV+cGOql0ADwuU/DB6CXNhelBVOSwSt2VrMu
hRElyezbIqmwCCLp07j1paAZ9+Brq4sXk/qBwhGjxUCo/3h28d9fjdIuZqS8XdZR
T3tOEke+4SSK7lzJxpIUKvwz8QfpwtcXXZ5oL2kvtIlKus/LTMWaW6OnaAeBjqwg
5C1GITK8d7O4wFPOePL9bITv+ZOMm7mm+G66rOAgC4PIz2zqU5yRGu1y7ZacE1He
Z0qMPvcUwaznyOqJ1iI4V71BIW/HdBazOyuTW81zRkDOW1BqYphVNsvnkyVnmWDn
45X5Z8GKqYUxjnWZHfItn7o0TpFr4xzSPdBRxPvQDmp75Fwf09yMi8gPk5r8NuHq
cqAALyh/NNCHlyiiGbOp37SqIK14smtSfdNTC46Lb47jQJrd/JLwGd2ULR1C+mvF
H7HqCmGfo0S+wHZ/Kn5oxgiVppHuggeVSrx6jm5/ls3RH7xfR+x52lhk9VlzflNT
17K0Z9kBbWsA9g4rNJT56Q/QHj9zwHMdeRjwENiMG9ONCqp/3nku7JUJJ9S9NlcP
fdEFW3KdTjiuqbaaz7Art1ibSdpszIgvecdRmpn5xD6go37iejR1phKu8gYp3a4e
765K7pdVq8vu4OBmO23KczNlZ1NcVwL/ClFLIx1GovlsV1Spx+P6xUsUCAViaAh+
qSCSS2+6WrwCBaZ+j21q2mMC/lz8AXWzd2vEzdTwb2IvD/MjspQrn/Cr0ViP3R2t
MMQ4zJ3Hsa6NtQjDGW8P3YkLkM2SfeskQ0HTaeBjD+lzPj8F/9bub2ThLjoJacSw
vQ8OJa5F0fZyeXpotYjcN1k/3HoqgHwYPfoIR0z7lKCk5+USxWvfWQzB8azzBvg0
NhMC33IOtbifwhgCPHXoxiry3LaFrDAluv8PIxP6rZNsQ+axDzk9OyKENwAj2r0Q
QspmjjuaaYIXDi82STsp/gyfiovaDANv5lyIaAkqoC+GJqrUqO/HC72YtzCDJUJt
KABsUitp8Ak0AVlaCQRcwhBfRoWdJVkRT++jmm94KWjRPLoVj/aqOXkT2xGOBjKf
3viQK2JjUjcmeOVwtqBBXrwZrwKK16NM10JGHrJ0jT8aRp0KewWwIK20cQff4lEc
lmyW9dX26+bxYdsKaa3khTSRmfi8mkU/pNSYSGyXibCBuKvYpfRPGnNHmDPJdcVG
6HBwmn1HYBEvTpzMswWwO5PM6+oCSA4Asa5SPGSIN0bdntB4pmGV7Y1Rmd8fJ4YU
1JSUClTLlPIb5XWhfrvXIutYFiDOxgILFoqb8xg1nOsaxn1WQwkp7Q78cw2msUie
Bjr/u/M0UEwW/+akC76wtkhsKkqV3V16GXa6CRg3kfRNlag71GljDhMwiCiCmLYo
4IDCC6SQtfZ0gOhx737MJ2c2I4YgBp2I+S1xE/3Owc8nPaQ4bN9qdxyGd9V9IkG2
7cf1Pjcv/IFMbzSJEJuBwzAiCCNmr1sC4VqarUA+uJQ4XSVR8Bs86rPVLdyAmG4q
qzF8cLHdpqG/Aer/p9yYbC9Mq/fbP+mH+FaGRv2ODsnvvAU7+161wpoTm48NrICG
81uWMzadLcLKhdbugP7mVVuFkQ6LoWZu3XwSnWTrBlBsd3TbFv/kwbdeXAIRShEZ
HZTEWpw6+9sMXhGeYK0O7Ptyask7iHC0dBqsf1TcTHgI7tgjMkcif1YMk0nRo1wQ
fNmofH+in8sD1CZmmu/DX6HXsrNzw3b8A0n54llWjwsv2+yM8aW6DX9gCoqIJKp1
yo/Inol1LLz9NljTsp8f3O/ALD8ZuVLYTJe3rAbYZQXrgbGf72RBvozBegHL49Gw
l6c+4bVDkrYL3TsN9ac2ivuexSQuTlPcFDCBHn7xz2cGW+xXww2m7igYuMWtsrjW
RXGnUXfMw85wDQ2CoJTWY1q1h5awfbNAl7wpft8xtUIb45BGmZKIDz0ulcvq72gl
Gh6wu/AuhKtJjZSxPKeNlNZoeXmG+pazdqGz2ywfXkQVa9yd3IajzlvFNAlDV5mZ
28yEX4TBlRSEbhO435eoFjHf1b9EdPOPba+MjhD4xyia2+3dZypiT/tIYFAgGJhC
DD6pK39hnz17X0a6UF8qWYplHHugMPKBx/nsWITzRx0Larxn9FCe1zHzN8ZpkIyV
iyAY6Lf9Ce0RB6ue99DCOrgp4kkW8VPFETlqItRVWFq1kxBlnQ1LiEmRvAfqt9X6
xNV0FFae6O+XcpFSq8wA22TyMsjEJS/agZ/BsTNpSipj5/WlGItwuVbRrenNZ12e
4/txMjAnqpSuSG/W6DTun2kPAvIAM4aIFYhA1HBke+H82Olu4BhpfzRivcERCc2X
2byu1H1Vf3Zy0LmDshD7dF75uQ7XDYtvaN8RS16EKYtS9zuK7UL6VG4RAbP1sYRP
Lf9ootDJ2nisHtaZWYD1KRvmNB1mTl+ZfhInNtPkPtIPMM6+xUjZWIi0IFfKsCPj
INuMstm0C4qnrGz02Qt/3RwrnQ3dGhofmzamBvSYKHZknAS+7WahNnkBvIiWUu3w
xP9il09GGgUvQqTTHf3WKcyhGu2q7sIAwvoS1oMlmqGiFI53NdsytMqSDM1L+mmt
ssyStxXV//O7Ypx79CMmhY7HOA/BCtz6QMMqOydPEPVho0YIZhYwxt0+uE8wUFlJ
0lzL2/X6qMwGPNpMeL1ukkbIb4DcOHp089UPtrU7/IZOB3cL/xVylmdDbHCtMfPg
IBtGWAZBcvMRZDQQdLt32YQPX9T0UmX3Ruyqa8cdXQlLsT+tlxVwsbF6MKHrkX7J
NnQdhM3PaXD7nelymiULgMfrgCI4SAPG324tjfkId7koFPYcIc1YXxD9aefNcJo1
LMp/eOyzQ8dCqfqBCpnnbMPe+Cs4kT2zA8bTo6zR4BN33JS+2wqD2PUf4YtjK/uT
t2Eb4B2K4vCTED+URPXxFMckwRHFkZ8+FEk4WIGBdPpilZ+PqFCelXxzl0HVFcqs
DCuM8+x8GTiENIB7kdxdQ9hMx6gB6pAr6I2xDLiQd5G4O3Zha5UnVkim3A0/ASXq
tlPiOnlIhJVyh5W7jlkykAGdK2zpe72i5M9A/XYiYdJAJ5poF/QiqXo3/IylP3T8
ws9teMD0SYo4s/irKLdscqHjoFClXJmMqpo2lvrZUG/NvJmBTaDr6IVN9RtwuQri
eQyzTUWnyWgVibhAFSRmRctvLQVEDikQVK8wEDETtt0Pxi5vNQ9AAm87YflZrRA6
iLN9cfAioyTX30PBYIBngxTmtcq3SXw5RfCuz5ZwQ+fvPzgpP19asZRolRplX7k+
ukO4e29Sr3DJPt4WS6EAuYmwArRvfmz8arhOxUOaOJNs5fCj0wuUNiHXUDFRPq9+
H2sF9uy6YhR+7GH+7hAyZXV+jz/9bYkky05xsdpZrxjw9gZGpgKl+bR+iXi/s5HH
xcSJvueR7OQR+st0XeRGm3ryig1N6hMREsAFR1NmKdZX/og/9m2E4HxpflhYIaW/
biYdaMwiGcpXv+3iDnJVwJorG52tyBxqFhfDMw6SEJNgjJRo4GU1YP7Siw2eqG70
pqpadaS/38FIIDE2Z2LdxInK4FIyks+HGE6UaqdkacqYLfw9ApH1luDVVVPK2l1q
Oih7bcJ3WQXSSvntLOEVveTIEAd2nyf1ZFfnrf61431rBYWBmRsK72d5Q7P72c/f
xn361l5H+Z/Xq1dS29/XD2xhrX4nLJu4gbpAfIiMkMxDY3Q19qF40H5yuH1U1T+8
2R7TqTcQxN903njg2asWiiRLx12VsC3ItdMaGngWy/xeXgMtNDuh5QwF6DfXNqQv
d7YHy5BP1KeURjzZoMKLQO1ic7caekG7j5MMQ7IfF/hW7a0jsyAjCAkL+s0BAp+k
jZBsLGqSWtM3Yy5akR30Msw8ncNXi8oyunGLAyiMp8YDPLqWqMGAtrljOsag6bjr
L0byAXMOxFcP1Eu6sWPEZedwHGVMa/O86FstoeA44rpHJO6A7BbOqjAF97qpIf2J
LWViD1by4P/nIXKwoorqMQ54IMOkgM1cfsVX0SBPOOGdm3/6brYplVyWX5Wpt4Dl
QiCR7q1aZHSF6DpPviZoITFBSg6508Cg7Z91YAdcoK5E+ZvlmLrW19mJVWM/wvxP
YrC9lBaHBYqOVBwS+I0o0mM0fjtL1Zhe8k2nclKpReFH4YZBnCw6t5Uztaxii2Lr
UBaa20eLjtIaTCdh2FzOPevS1hILdmc19KxrNb2ilZgmzNQI8BH5mDcMX2BVua1J
bAklccqD5f2Z2iBUsIz3WiY9n4kyWgCHTJUHhFFVAb3jslp0dWY+chm9oIuzzCz/
0z9/9XNaV+753pA+hy9nlMbGS36i8N1X+Q58017YnJ6k78Ps+Ca1a1J95HeOH/YW
KNledy0Es/9HJ5dJ8GJCrbbRhGDy0SXkaqCMLyuiSRz5iKHKVVnT35YhgUOicJPt
1ZWdczUqcypousB/VhWecm2hHkVKlpLsW6E7DdN2hPREJmPIMv6vye0ctB5GHxRR
WD+SMPdTg71U/EaYRUm+n+fdRavzI+Jc16MN7S0Mm3RQVcWKrgXA1P9KTuDKlQV1
Vnn9de/bJGDYqe8QLVREXzo7+8oHNoCw6zt969jE4ySkEGgP+P4Ukp6joqIkmoY+
sGrLxE+FUQ/PPkmONimBJBxotb1yDlBt11ibJvPp930jy1v0Xt954KdBMKpEk1X+
mrp9YIMbg+b6cWA2dbWm9SlgwYREC5d1QfYMauUgsqa8PW/bD9rcagdcLwcH+9NC
ZkIYH6BB9gRFMQK0wHKlo9YdNXT9dYoUX+R508ddiG3kdD8wL+o5ipNJ2CcSs0IX
2fhILrQ07k/AaIlO/PZC5Ya97PIk78SCIMzAIcgq4Pg+DjD/LVjpNERt6UuQ1UJ+
mAaTG0g8LUkB01MnSQl1JXR2DiGnvD15EvmmhtQw4rzMeVj5qWVTM4tjQ1JBpZWw
Zt/AT5SmiISVBQbZ9Uws1uRKspp0+QOCwKbHYWxKOOVsi8YvPJndX8v3/HEiQ5QM
hs+2cbWtdp3v0xlAjvINHwdItIuAXfoOoUeUqJtXMe+UsSOu9SG8bjmT2uaHucSq
hgsdetkI46townpaS1GVl0QxbN/AAzvzNVV2/RBKhQOfoC05IuuoX5AZqeRFvRGM
+TiWIzRDOwzYbDY/Der++2aeOv0+bHvw3FeFYTMjuInzyi7dGl7Z0kiqyxRbHeSE
ZJSObvIZu+kwK4pBhC6UIefAmNdv68RCdPPfF+CibisqdLhtk1u2E3po62OZp3Pb
W3WnUuzN8qHFOhSF9/bCxX8ZNCqV9DmrUF1qj4yrLhl6enral2PqlHA/dL3gtMv4
p2bDhCXmfe5BHzHozdtfwJT+JD8ellSJw1nfpeMy+ap2bTdX7LiofqXOlhn8Qses
VvAOmYtqAivKkf3fVkN2rt99x+ifGsmbQzpzqm7agA6y0n8xTfIm36DBTRLWCWcJ
Wortk+ttFodZ7nfJtGLdzMF8O/vbu8zJaxZmeo+tCxh0Pz3WYF6Xw/gBIcPd9kvl
tILNGfM3hTQ6EK7y7FcN8hqn7I1IHIFtQ85Zipo33w/0pZJ9PsdS/aDoCHtqSrOH
q83lsH06y5GQ5ZDJBKCuL7LaJJCCmLpiKnOJOtGK2rCNzSsjXswCbtYXp4tVcai6
zcPUvEWIsQjuVI3UmN3XOMqWjrhtyRzSGRCMx9XS6qE8W3RIyqMM5taO/nK53004
9LJTmpzob7/Ee93Cnu7b4k6GJt44upEjNVgkRZ3l6UMw2EsunGj73LZFmWTrDY6a
R+NWMRQSl08+Ym28fjv7RgFLRxZT6ugzLSoDClz6O+Lk/kdhjiqUlEPnlqNYckqm
cuFguDtuTn66LrMC5A8dIUPrY/45kj95fzYOciEJpPKYW9lUxGtqJKlNEIBQXb2N
Iu04uJrcVp24yY9++HPnuj9CzUIrfa64wmRT4R+5Ehk2Fi8Zwa8sUpZLKXZ76zxC
sYDDwP0JjeQcv7sUBeyYRuhSqWPfRPaPTCdtmOx6uUA7tnWpj846W5RCvC5g67iL
WnpP0mV9/Db/Qf1mAYomQZe504EOZc2x7XNkfTRj+Bf+dRdJJVP77BrwjBmdPQ00
72ORNCQBK70ccZ/F9Zg2V8fg07WX+sl2e85ue4zHw0COU/PsgA+zcrLaKi0BihLH
ak0LfGsMFgXCC6f9JT8dhuN8jYiByNO9Q547cYb8xapky84uEcrnRgIDTz8vQAFr
wqo8XDSj8cJQ5o+qhdo1qhX4teBWHgU6x4YM2vNxdZJYqbYfIyz90AC20nICHN2I
MF7cFkDFY/Ryqsz1mk002VS6pJqZ6D2hqV4oH89sV0CgAlySfpn6GR29zlgo7tia
apdbQmLaEIeF1lQzhVDPlIgKAfHlCohxq2Db9Y9kCMxB1reuVF9lherruZ3LdLJO
Y9Gl8sA6lFrXjw0eMa2ZWJEB+JafCiqPCd0WeYh9nqKM4N2q0Bymy8tXwhoXktgz
kgXefvt2Ad2tuniUibqJGoKwwTcpcqhnc5JoSc4HDkqRtihdnsUA5Qeq1UdKPdrM
98niGM0uM3CoS3PfFV5GXZE/QuPPkYclet+sj30VwdNPqTU0mhIFh9KvsuQ7ZZA1
QGu/lfwO96ATzCoiM+9C6itW8FLDjFoAf71+vpXEEqcCjZLzSmD2lt8rvuYgbrsi
RU4Xga+mLcx/rMlCn9rt2yXwEoKJdLMth2bejlVOlcgwh0amw5f7twTJ32vgGQnH
USfcwsUzlgwELNSgKzpOqBVI5Rqn8IM0lr8X3xx31fm6TYlA4ktdOpm4EOsA96Ue
INhO1xPYj53hf8iy/V/G/oLBIIAB/1paPfz+jqtH01MU8c3zeMv4L1e9GmneziJI
Kl0qFY28JQrk2Bv1OBQz2VY1tn67foEeH+GjCw4ckOqUipz2Q2JSukqjAxEvoE+X
pY/xJi2hykLQ0UcU5pqJcLGbFj4nN0mE/ifuXIO+Gp7/6fjmawyqpRghkz3+Z54U
fR2i+H8sx32eMZcCKT3eMhIoOtDhE+/ehZM4hEyDI7OTGx7Z+HzzVZnZDhC3pU/z
InXH83CezZhy67kyi0glzGiTjfXxwGnrD8HNccp7XdQY1lxSYmWxC0+UhfYeZ4m/
EOQm7ddmkS/Zvc4k1XQdHZnE7uKzNoNNhNyj5cP2EjrgkALeh5mu8Zs+PG5rQ1y/
aKiGRjd+fMFWmoa8JvO5M3xPkZ1OFqd3dFJqVTIJXEhyX2fppzwbK9EENEmpQ3YV
kJAmZCjzoO6ViwVmUYOU4AHfFmfJaeqzer+bS7nStNXWhosb3YwodjFslmRFoJev
OdMBjOsCCDzriAZVEEUqI1XUkdtMFXqX/M+zIo5KmDWEyL2x56Rnjc14HMY9o00X
RyAUKKEshRyFuLSlEOovUbwq9iZyIBSsPQgptiGY5u+G4gpoe7yeyXyyyieAIs9a
kmliPCM4Wiaj2WebC7ZhK3S1zgJ8HEkX8xYmwBLJh3Is04N80kjhYfRiSA2lQzEP
jGxnNAsB5rUu0Co5unFtq6FY2Y0K8n/OWRy/jZZ/L5TjJofRpIQ9BN6d/F8mOREn
IBwOcMOztDqKg3iS8NJ+GFhn4mkYzrmHzm0gVGfhRgoSM7SSO5n2m3/GcLZx+lnh
avsBl29eypVd50u5eyyc/mavtFO9Fc52XDj0U50ZLe06RaG4ywtXCcZsytu92ad2
Gs5sx1O6SeDS8/ZNzz/Gx0UV1LJrZu82k9Lw26zu2XlrzXAv1jvjH2tG0YVHqDQt
H5PcZs7ssDiezTpBJRYj3NwkVJRs94Joa0xB62E3Uewy7wwt+7xj9KXkYoOwM6EB
XN36rz/HjAEMJEyrubaPXdjQ266N52MKDS8rHv9GPS9kpE2knyRMjIcUfF/o7y6I
BcBxDU17a6ZDNWXv248cg9wihTMtT07gzePrIvRJrZwzkZj3nhxGhmLmUqBYJoj5
Va2SkznerIgWs8kMWgQrDDIR2VAGzaFjbszErPKlBsQQZ+oLr08sIQKmqgLUw+k6
M04XQHuaQ6ZX+vZYGfzaZhCv//q7tFCNergo81gh8omhRuirC2CVs2stST2mi/lc
3sgU7Pqq2wXklifTPDRlEoKldMSBxzjMCA8tdVC46bLljnpHnHt1oORnhaGO/LAf
Sh0IpzXrwMDeZvNtuBxcLqr83Bv+6coXMkomdrc5xUcQSgAyYY0c+z0D5fCfkhH9
E+Top6wytlaFE7myJmB/kXf7xYzhqnVIRcoP71AnaswRXiupR9crG47z+SX6VeFD
sXMQZjC4ayLMcvKg/e9oHrdtMEueB3Ar41KPmb0RSTUYhDK2yUMmmBBIgEbDgJH/
TKg4QTXmFkpmRecBQ47NIuxnJOLzY5ozRbk3HKzI7j5LX7m3RH16ji+hrNYqlwH7
0kFnHM0G4Nc1ktkNxsucNu64SotxFb9wkjPUQFaQ7erfX3ilobLpwN5f3TND7hVI
zBpIGmphI3cZ9n19bRuONB7jcfrqO9IFbMR8tBhWdgZcmkzunRzf/FLOJX37fxQ3
udw7SZWFVD35y1cZ35K7uv8VmpdUEVivcLiOXdbuOI4cpYfM/8Cy7GXM+2SF9iXu
6PL/GuWE2zDiqvlCFORH8LUqoC9rZ7mwJrAqN/ReThKYwLc/sAAPQ7uwb35aKum9
UiAEEsWTYUJTiExV1tqQC0vmmQxwvR/VqlrYiSXSdUbMN6d23rBdfVP0x2T7IhPP
3ggPQhhk+j3UsFEAnpceAcq5Atj7AVZ24Aogt6/p0hOqipGRxJ8iFhv/tkKMjEdu
+XXUCJZWr5vJmSDslHC87lRmIrpn8k9ToaJlPJei0cuCFDYg4V8FB3aZY2WyOuNN
svdwy9jlqvnBpWuQB/oNtNGfTfCfrKZqm1ip5sJtQtR7gBSA3l1B39IgrisMpGDm
FAlPwu+BxXF82vhWhrf1/xyD3AwjKfcPTQy1pKZ8JIno7Byeelw20IF0PiBQ65Kp
S8SuN9dkFEPIdI3pqMDlJXB/1XMNqjRWBhXhZ640WlgV3An1c3LFTIN/vrAwvCWx
Tj6LMzes1wnyTBWrq5jZgzBxvsvc+L/tc62cKOVfjGPG55fuf5EwAt3k3OH1Lw+d
q2N/vo0JUH2yHYTA8ceBBOHQqsCEXasDbWWMgPVxBXEM4+N7VYCF03LPvF2BhLAk
APmpCcXOoSpggaQyx2LObX2GbhmQguX4AnecCI56XdgL7YyXfUoGXp3E1+nkqFff
GC7ZO8CKGhExGRWB/SEw62fyUoMigh11u7z4yyOfa8poOneuBN7JaEcIMF2n6EUt
mOCiHxdUvh2I+VSj+9yKgFRb20Kj88nVV+eI5FywCwmIRAOBt4sPsW+9WbDx3IuM
SLY7iU6SmyV+Q0yw96PpndVfijgcqC9I1LMiTO7KxWMCzmAkllFJTHyDVqARNGVC
zJkYeEaF/yx5vfOSmc+7SHPT4lsck+V/B1v4pRj6ZgoOfQgLpzjtsLK4MGIa1fiT
ESezFTuwi8K3KvWU4xB0h7Rr8PNhWQhgts6YzNkB8Mhyv2XSp5PjKxoLUjUPuO27
Rf9Ngj40f0tJU9n9JTInyjivFf+hZhi5KhYRDVzgXDD2s8/5GUU2ogP4TdVOzFcc
fC65kcS7JWkKgTwToZ+nR1aG/KW2PwYPeNsnnxGhGI8m+hsSrIZJ8ofcx0xbeeL5
eOu530KicRwoRF1A8V4+M3buoc1D/cdS68yW1mgzY35uBpBilOt5YDpk1qjysWCN
+qQy4efxsZtMBNlkDm4eAmVFXkmCwxVk5ekkN5VTm+o8wKAVmV589U7o9+ZfgJFg
MO2d6TIX0W1dxIDWwmExeN0HTrieomvombIf+llq1xciL1LkKQopVAFOaFeyPjPo
+FiC68/Fa1bQk4dZEykUPyzIycTUDl8la9VjPrYQPrqHhYQiLO/aKRakjQF55DwX
xtHLXjFCyQWJ55yeak7bJndmM4VNn7x85GUsntH/j9eqoQfXrnf1RyK7rJBCEU3e
EEevzy9qygdnq1odzckLJTGVZ3oZVEtaaG7swyde8Q4YxxfrAJ/2SMpZkeNpuXn3
w7b8NrFDwqCx3X3Twaf+id6sDS+E/ZRvflXyN3DJ61kKxaomNC4C4NUEXZRroysO
yEyrVGbdfxyL2nQYVJpMU++ji0LWUXXlif0k8UsSpBUgA1cCNzqNFRwjTA2gaOk3
LlKXTHJ5Z/o+DFWNci6hcxKEUjlWd0VrucjrWEiYZx0u7icqBTepfHabLqaSF4aV
lfPI7yGBRtRuE6bXSJGXR+o+r6TyTssqJ3aANXFflUn+7qVncRJXM0ex7E8JnRLi
VX+RykfIpApzod56mNuAsRfN7AYGvPn66kSncoYeNY1yFzx8ASln2F3RI7wcGJs+
oNUWCxwIip+tCmiiIsBSNwpy50PPBB2bujfqvv8S+ZKu/I+nKWdQMqnMx+46C2g7
N+i4X1S9Fin3FULjdWnJ+EnGINNgir5wWen6WxY4zsmWJs/HmDVb4EcPwy10g8kt
qfjw2tnWbQX9K5nTNpgqxELwftAOG4dGUMo9MyWyCS8BOVv2lIwsa0Gds5zhLCvw
WyW/7voAHIK/LSR5OM4eRsJyndOFLaQEtakT5toyMwruJ6WSa6KtR3eZHBXuFwdo
pw/ueY0WVe0cpAAiSwONo1Ra6huBhEBR58wy32jIFaBwPSziVg0rRNP41F/C9B5G
vLOXuskcZzGICIan1SiRmzWICYiraWNqQEr1oacnAou+LibI82dwCvpQiQHQLTyb
uJsd42eMIcX2LGtQCrX+rxct0TdIIRs9fuMz28hVL8AGdITuiDklJSqknCYsnORQ
fszBpH8dTejJOAOJmxuA6GmC7YlXGHcpVsaMonoTb9RCm+UTHx1jJ0lrzdaHFOQn
hcZlzpyl9osjmRE7pggG786uHv9HujcIU+ecirXTeKlYMcFHIv05zBK785/ICIA8
6PCmdHa6BosEhut74IMys6LxsZMNuvKHkbnyBET6H78nX8gRV93DPivVAoFEJY3d
S96Fk9A5ano6Z9W+6quGgUzmtq+24UZun0sVkIsUuQzDk7odHuJc2pEjtnq7AGAl
DhdUFAChE3aL4MGkGMBISoR5WrB9sVEjIoYxd7xNjd9WajQX0+kYVKj4MqQsj9x9
MhzNdENgeyq9yAZ75Ri+HbFT6sIjhgE4TU74goB9qPpwN/jl9eXOBM7d2gboUONK
V+Nthr6dNp30vcQyjXmq4zFf0txDopL2uYcpCl/2dF/WrYWCZshQNs/ZM2N71gXV
+bX8JXMUBp+xG+QYpPUauTrizjzHvhk7V366S6lGppLOk1aca8qPXEAvpbIJVjEz
yk0uoBqlN4vJ/G187lot/Nq9T2FkjXQCkN9Wu5/qI5We/b8YGoZkZCM8YA26CR8r
UUNMlXY5bH1s4EVZ2eq+BRuQP3DJ/tkgTa3Rdh02pZMqGrOjygsiBYv4m12rcH6L
Mpt8lUgKkq2xebp59eGA2QJNlG+NArH1TCJ/G3A7diP0tGy93/EzMQt3sL2beowZ
o94GaLoKyD78C2u0kUmBdr98KePHDwq0KTc8nZf44C++JMArfWJH+X0V6ywaPxHT
v8aH07D2H2S2WQU1uCDl8C6LVvS0cf17g5qgVITjYOKIWzc5WOZR4yQMvpTwR8ql
cS7PDCfsfH5bs+mooz1ypFxiMeZ5SdhAQN6RDo1JfmIVoQnqm3JIF9gIGgHl47zb
KPwHrE3XGU87pKefTZ5zqxeJ1zz8u8ST++kOeaRP3dxyVTX3KHgsIEFHaIWHhlsu
DX5ofq0EjkwjgzR6jWO4CEISRvA47M6WOU1HLTj4epsJw3bEdcvI6I8GTrllNPoj
OVS1ufOCP8Z9CoRpALVtQHmgpe8Uo3qpTEA1rQtB2vGeApBuy5YepXqkHk01bkwn
7FiRaWOth4gduSvUTHe2xSjLPyz0xpInE6URxwB6DJv7GS02lDwNobDuVhyaZ9Kg
ollJd+vlACRxmOOC/IHeZX1De1nkvoFlQgkvGX4mT7bBXHPniPs8R7gMD7QXbCke
Qr0nq9MXxjDVqvEyKSw1oWLfqgbMYmo1CeYvxjkcmVfUsE/Cenev3JmZ7bM6m92i
07sG/DLMlG/wx/4SpYATSobQuojd0bX8GPDqoBUhU8c+1YjVFbtsN9BGuMR9LkP0
E6BarsrvOUzcFJaO3M3GOSOsiCLDEXPQXgYR97AA1NB1Ut+0I4xJIpQa6CnkiPDu
CvOTYEBvN4sQTRM2mXpanYwhgpLatjUpPxMfnDsDevZJT2lQYlRV9u1yCtS3rSYd
gS4ZXuo5l20ztRDAtgeBVlArl83pL6uQPLP1+2SwJPvTegemdHPoEfCWFJEX6i4d
eEq4TEp9uKGmuhVCsNTd2BFqE/QEK0MDWfhx1VMWE2b7A9P1rHgxTNf/BAWHPj4C
9VaOl9sRSQ6yAX9uiGmyKlKOwKiZFAsB8+KAQtSKCT9bJ8zhAyNtZCKHOjQaVrnf
cXmdN1UoaVngmyZskR3lOYlVvocPaVq1xvrLbiQ9AKlKAmaKAelu7G9EPS2FgSuw
2PjLn7lwjNibpuJ3iFQ3LNy/LQA/y8R4HplUCGSS9xG3BwPBbSKca/hxLg7ubwkz
cVYDCKteEy4U6BJoHp0xa2HCb/kvtsCCXbXqRmOKfw9eT3vzDhHO0j6U994Ec4y2
NEg//wNlF0O9Tt2ybniUNtylYEwOjdqRPOog4JhozqYFhKTcKRihM3JZrYcdLBRl
EH+sEa6o34M9NZe9XyEbFJO3kK1ZHVJiXtqQk10MXzrElkkc0en2ARGE/uM9Tr+y
I5O7Iat4j3psQBgPzYDKmX1t02kQwkSV57p8VYvroNHlftFeiaXdd5b7/mQliy2o
8YuSttgprhi+XdupvpQKhwzLU8hmD2JvBzf2epINdRkOvc4nRZKZU+WNstHrpgx6
pygsqmoof397k/BIYCHIa/FLc1ShYKlRqs/M5F3SDqV6TWWonKMNv32XD4KvIgjP
UyZlBVruU/43Gcvb34oxJjVsMML6jp0Lli3KceEtsc79qGnw+cA9jCWD2yQfLB+4
PETpfrASoyJnDAm86X+WAFJOPMt5FCbpGtwVITTae1JcJLt+tI9Rhg/6Cxlo3t/b
N0Do+klvPgjfO/t0mAKVu6RySSEj9xnk/bUWiDK5xQ80ocsZggXQr5ECIiXTS/Z2
8Cy5B5n0qRrOHRRee2O/Y6jbTLbGGg8QKFa7Ucx5r3PeHKO2h/jqbwqqxWIUbPij
vGTAuXltslBZzbmQX4/otamrW82lzUwadUEh+Gs/ZKofwuNQbepYI7inmAabyt/O
eXeahKwfgcbY9dosCeeyfXXRjbXWi9ibwuRmYaiwQoD8s5k4+nh5TkkprtW6Uy4/
erIgX4fxJRRJeCl73yX1wEAiG3WOlVjJZCcM/T9vD3SNxqdqx4ziNswwb7LIrJeD
qJ1wx0tfwMqjbYQNT3dKpozMsthyhUcOjFHmzYKpazaDFS7b1MM80ga03WylqSGe
gjCbWetcnPF2vYsEVcLMAofdDeMdrt44/DwphDtt6YzP3fQZfLH3OjSecViXmtwO
olJqnNfWWxdE9TUdLP/u/RCBYmmMNnTtv4mtGvBNgjnZgyQrQ4t6STGR7R3wOy48
u5wkyRolJQyx/DK1cJBjBAR6YanUeL2OnwG1xpE9YyKLLRlADpoctRjkzFgVOapZ
4cZghe/Mz2uBN8jERO6R3CJHOkc63kknMpsdG1D61VlBxQTYygM3QfNuY2roj5zZ
0v8Ib44BqN5GsosoOOpjN0mpFrp3/k5daaq9YjaqQjn5CetiGIvrPXdxPewWiPKN
jqq1t8BF49TwjL09HVYD26k0bn1XOyPmQBw51MiDIsaSJRU558wBX32gtqrZlHEr
EaLf4eEIdNSfMAo0Ajzm7TrAP4efT6rSkPjumxyp5aKq//S+k6Fdfhn+qt+2j7j1
zRvibjrgtRMFpYekVMLtZQwMiUf+q/sisVwpIjtFdS45hnucUw76I5o1jRNYDSSV
mL1utP2tTWklrYXG9YvYzquC5PRIkiBXHPrH9TJ/12Q2qKdsxst1A69Cty9SPy8u
EjBiBMIsIcIrs5cd+aFKHV8PCq6ybXLEkG5CqsHUJoBw/Kqmxu3FxCeFgUvCNfEt
Ucl28zjgFLni4IHBtbyanFwsixVyOg59AAoRYcsvVsAH0tfWpOFlml7nFFbVHhKR
BTkWwudxqHwaquV4FaqjRemFzKCoyUax4ZEzSxWMAQ3GUZZeJUI4bbhmz1CUnC3m
PntdEGpLCWX8tr+Qig8wtUXDGpSkFNvAQk4ps6rXFQQlY0RchldtfjePsMmu0VrC
8hrsb4wOAD6e2tm2pLN76rKwBwwEW2uxC/iszeONOWGB8Or0h8yCFMsxzk5qUP0j
qq2Drp9EjPg8Ugmc/6x22hgcO7OKSyU9bvJ77CgT1vZAI5gqK7I18erJ6EwZliAJ
spWS5WT80l5W/F4OCwmN/HICx267MU0tiWz1ppEPt/p6DFa17gtNxZ3x2SFW4xTw
VIuLCxCrnP4USq6Fyz/kXZjrWMyiFn3vnISYF/PTBTD/LekttQWT5j8t9zGyKett
H4BnfeFHlESjX40AXeonogjDMk3Rkp3s2F9RlwmexzyKFTutdFIt5nTJUicBVloZ
6urRp3BJRkrJSxOEADFnfIQGBQYftC5dcW/Q2VTLlG2UcXM6NPMha5yntHYzfO42
tttOE4l0f7htsNnQ4m6ef4ki+J6WIh5azA8Ue9Ae5od2rA0wViGs7j2KN8kd+T5A
V1wC/VS4S6ToMXUyV9QEjp66oWSaE5sQEfMn61i5twqTxlBEcnPubPmuTq/5SZGP
L/spSF3yP0ibluVey9dX1xvOeic5V876Cj2h365t0hmKcLKj7u812kmXmtaYc+nv
fhwzoCoqDed4u43FBNaaqUn7kDKzRruLeNKCPEGfBc9QSDzav997BK3MMEyqdCnA
2/qT8v5szEB+WfJR1106zPlh0LG0N29+HJF2ZAUauutCkArXc9qkyiJVoDk0eZTc
4yFlnuIBIAJgXMnxsWnMvqMoLicmJ1XlkEuAszs3XD2wwuaoNy0Pq1fNBztORNnt
VDVGcF18UOtmR3G9DPcV/EWVIC411YJzVHRe/3LSO1ZwdaUkLKkjyAc4Mtd2jmdk
st/PyB4OSGN/ovwtOuOZA7zIgY1kScxBF+MUebV/ugSpTYLUJdMnCCaArfZ1dL0s
8rkuQ3URXFVeJnZ5QHyAkxTC3g1vqv2dwiVz6KJrI4wYYM8A6VfFg+z4lhCoQLf7
m4ps6oLfLL37MiZRHrucbjQxOQ1u6GF2u8f2o6EkWzTbdnS2ndQ6DIs+mZq6oDFC
8YBATw6AMzJjZY35ntxqKMl71U5s0lpazf6t/zYJWiSP4NmMUywTJi5XYOQTYsU3
6K7VE9fXV3UKvsxHBPPnk2qHIAq1TYpTx2eiuwB4V+tJmZdzrYDXAISdI8FJTDOB
mpQZZFu6yrSwodjFzaH8THLuZCw0df1HMaM2a38C8MqaSzJPFATaOGLGatKtdDdC
73/vVmg7Ol34S2hDPSYTkMe1hMGedW90l5U40b+bczfl4HcJuTRAOgstXju5aU25
nVNAd1Wf8hWj8v84ZPyZTiHEt7aS16xmktSVE/qVtdfF9+ZnWRg2icQ6sReRuBi6
fogsqYu2t8mAEqIjAyr5vDva3l6SJqH/u+qqS6p3OGNGo1tOOVafgo5jbzPfipbp
RAtTgRLcPkNzidUEkZYT1g5IxjLhXunx9+sQ3f19hA7gqYhr6qXiEffZFyC12am6
GoKYhjRhsQ/lNZlfoOt5IsDYmKYvXeZvLwEqZZrdsW7NSqPHV3v59KS1RYAK5VPL
TNbVstRN4N/S9IO3tsbOQRlcwaVBZ0mM0kEF5qHfvJgd/1ji241i8RHzW2D9Ckd9
0RTUm0jfwCcCaddSMhMd4/Noraxf34ILS9rGPOdw004sBQvk0pgWedtKRUV9zWD9
lkg+n39jezGsGVZ+Sy49/jq0StKiVvJKWb3F5n8RKXACoLD/ov7OiDBsWadnlYUc
+xhej7xNwWrCna62UmyupZYgvrr/RnIcjP+bMoDhaBlCDZ4LcBxKeQpduHAGGShQ
YRsOF39n5FZ1jXtnKTQFiUZW5KSstCfsopJyhIQlloG17/SbfN38uvAUxDgxCQ6D
ogKHYyJUOitZfLXDlKjnce2wn9e6SMtilpxKbrXGpNRgCccS2VlMZpuCJaR2ob/Q
1mQrCa51Jtz8GpRGjbmincvvghJdI37MWquUP1bB/VKGelxNwidwGRtaAyM6KXa4
zORXrB70boRxRq0RhH37C68iHIV/f15PWRTlBt/7BfbzrTnZFlPL+HIw+PK8CrQF
GNzo8hoejzLjFxlWz5paokomDRhEFjk0HSqnnopPSfoLesbv62BCCJ1RJfI7THJw
I86ZziGlZifw1506rhWcxDm5LwL/tlZv8LsLdDkX7nat3jVSOgS/1YCG1R0qlDVR
v1NBAB2DUVVbim8mxe44CvgFnOdU22pTB/Zcnwt07Ym18QVZxXCFNjvA1IEULxMk
XiAWGO5zvM+sOo/e4cKLjkXsT9vY67qfGGB87ublEYMtIkBXmHe4o3pKEHJV6bKB
HRVY5hQPZTKtHPc4c1RZW0yhlJ+cfj4kzEI4aUHKZ713TJbzAAi/gEmpe2mA369x
1yvdyi+QcIXv+UCDz1oZGepRzdFGPCJ+uT0+Str6t2Xokjjj+a88T1553s5B+qhp
o0YsMtZJvmOqJjRkK4q/H4DgbdHFOQUK1nxsIbL0V77KLIhUesUOaZpbC4oOFKWb
Fivp5wS4lwkGsXcuzImKlLqwu+T6nIrle6f7u+0Nf3w5WHX8vWN1qwjuMT0h0iZf
buthTJUbbUNFAiub+ZX79bzBNoSM7zIpgU3nrrEP4+0RWOgjYXye8JmCMBk2Hqq7
p6kYONl6aip38hBszVk2neEWfVfoPDG27zbIvBAY6ENrZgS0VZ6wfx64L1IcwcN0
0E6VTnK1W6TqYIAf2AMNZBMUwkvog5cr3phL0oGLefpGuwUahlKnbPgGzLGpTTsq
4ptFUq9BjdyU7pLe0eZQtR3AYMEKo6wJ7h8Bi5moGZ8AvIAk8lYJ55MnJ6qYjkuv
cdGLNvjJgWXm/DhBRfiDaHKKtr3V26Bd0d0tSQxKTUQKPx9Oq0uw29G4ug3GOICn
PTgx2C9OtEOUgjZEOCyghInfp1WOo7Fs+Ym91r3tHm9eDstw9B5rKyLHC/QYghFK
QnbaHSNJcnLWD3dyP43Vb3KekWp+vEj/ksm9BCYhH3NH5MT+bbcTbGuP/sWm+EAd
lilNca6g8cCTJ/ndGz2bid0PjO6L7rmE8wFINSaMIWQChsV5Ne2TivMVJxUG20nP
C45xDl99YllpU0xsuQTATQjKXBSw9n/BLFMqHf0+yRbwgLuO4aFgxJPHNWeU+Cx2
jPAnvNk/DlngtoRJt3cS4eiydR6z4zrjMIchUrF8p2kIAX+OYejmPxwlfpjLE90F
6YLtMCMb3POa/HQdTtt4iBHhXUy7pIR3+8OEFedKVeC8k8CSKkvyd+KXq8FHn+sc
z7vouszX6k6gzp8OwwZ/ImueptYODUATwCuYGpBINhWtBl4Sbt2+97CazvHbNgYe
kMI3x2YhWzcrxSqR/rY3IATkYkDL4Zr219G/dYvkSJqTs5VeTWnjUzzjCQ8dSdp4
CitrhCxjYVuH/fbJG+qZ7f1DCdxieD1NvH1NEp1nRUvx3DTrX36+GIKKNvku3gb+
XLeETwmJiPeuDxL7JudmlKaYigpGBKzVEpBsxB9/vRPVenSZNmQB2Wg+eyrWX7+X
+RwNDvRGzdE5nYXHNqGf+rtg/tkNZcxoEp0whbpd3KmzkryCHkatiaKCLjj5yaxp
KAbEcpsP/l4LOTcwrL1ug4XcidoL7J4AW/9A4XxYRSGvDM35QVIaYLQvbcVQn1Mi
Ali5OLeRYP1mErLlwi9au/P6b9At6psoraOITLRQWiJhtUWaGA1JtACqcJdvvIic
qwfjDc8Uv0dk4qeJxdAuTkRiFr9RkO4gZvR06Mkmf9sYV3zwyQQ7rOx6D4TkZve3
pDxZjISA9KBvF+1EYt3kMrN3cTuCvX6uQkee/S3sYxvB06Vxk1sF4gSNEFQ3GsUp
QgdZKuvZVcK0B9hD2VHeupKRalGAe1BUx3hjQo/O4MRecd09iqCYOnM0YNkV+vbc
bTPvEeDtjjDAUuHZjk/h837TO9a1jxZ8YceTptj4KMheHhkBGSUboQd5doc6vlYE
p91XvR6W+fj+jMcQxpU8DZMK3oaQnMVBe1N1XgsVKwmyFrgeUzYndwVgMC/UH/Zi
KO+2wLFJ7tUgznfRyP9lSpY9bneajUNbqK90tmIVokch0EGaY/sXfdqb66Pl3ExN
3FNPQ+H2awNhNtkt2HkyZ+JI53ZTYn6+RbgAOM8WxcjlFBdG/gLPh4iR+7+ocHh6
1EKK/P2NlEWRqu2t3BXT0vReOkdNaMln5UtUUD9o7j0cpnOCXE+13yP/lnDZkQuj
5slyxBFHvpYnW7hSQAzHrXvmteUl/EBGh9x0bzPHQOs9BC5Nikffbu0F1EFuc/5p
8brEarZRJ2J87DSX06huZYz5b5r5qaiGIRJvjVPpyGiZHbAST3+C8M/DRV9vu4ub
OANzAW9LOXP4k+nZfLQgW9ivAgCIz8T0dfMdSUGLnHwdeFT7k1xuHshO/fLql1YD
jbNnsnw42Rdby29cuPh5Evst0L3ZVl698/rXaMDILVZI1oLskzM+k7/wTPLNLra5
Ze073TqFgloW7KPFOFrBAetzLaHxjmIK1Daup1eI784Dlk3+c7/Aeb8MEwpyNzlc
lH6bHMNKq9sHMCOrupcDBn4fsxhiaEjufYE7G7PxYFNmMnFdJGz787AF8+8HjqqF
UIPsCY8DIbxeUDhGV73SXC6ZdtcaKQeQPH6Kq3hQz7jMCyLjExpnxP8LOesixJXv
wPF0vErtMduW2kQ05rbE7gtJyUcSXtMUmJ3AsNtN5FhVqi4WjG0WmqP7Q9GLd0OE
ocIouXxN8osC4qPPZYi9O6qjgCLdyPtsmg5/0wkOccG1PtNQMOQqGCAY33VN0o7g
v237jDehli86pOnbfxS0km7pnumhgYHSPn/Sib2/WebDSMKSAVS5bIC1S0e2ElQV
vhvjPkcGvq1qkBBQ4tfK0BtZ5tuF9j4uFVGeAXRLvi4Wr/BTBqZApC/NYJ08tOTl
OfX1Rp+3nKM9Ebp+AiVjzRgOwyPOhTx8cqW0GLxIu7WkSjEoe3I7IjzAAl50DUeh
Mow0GPjVK2GatZZe8zE8Ghu+FFNOBa+nLXZ58xkZhLkwV4Fuap4QLfZ3dJ3d3E7F
kab/DqCCemQx9DqI/jMUL6J5QQWxNNs1xJlFFRRR/j5hqezEty19Azq7XFuyS0Nv
yOQ02lK2w5PLIbpGOgeYcdY/RplvktuCVWhABBWAf3FBulpUWB8FNcBl7in2caE8
9wi67mzdcgtClwIZWrvooXYo2ic2T76reJTnrhYK44nK61fz5QHCJm6CSiEvAcGv
KKaP7IuA2Emf5qbKXZatOje2lB9PQzbyBeHTIhbfEOwdWUOdIbEzSXJGMeUjWzeF
xDa1SjYZ80QVYaZvgYU0sT6sk7Xh1zpZTn+2ey3TldoOAW8QXbbRwPfcHkh7bBIl
NTCNooYlgD68b4hUXOQXej/COwjgWgMVMGWFi9/H2n38wUZZzxQBvgSOErM686bs
eA2eCPER8xf/Eaf62JCLhmTsEuPTj72xrrjnu7XCjfykO7zpEgGXZIJuVUKeiRlm
LkfssH3E2l40ghtUWoJScICUimIJLqRsGM0gKwAbk10JReKJr532q7QbfQ/WzDxU
9MkrPbAdk4N4B6Aqdq7lNTauVAeCNVxigOq+AgW43nqx7ch6QFcNmcLUF9AdtjXu
C9fPWGwGpPQ75ZrQsx4AjpT9JZojFpF3dXc6AmHFSkVgEiJgKhcGONHIzrpJ9FUo
g6vhHAmyk6H1HQrln108ifZ7/Rwd8UmKS5wE3wTssF8ovYRMLBTieZeXiLYIJ9Dk
UTdx+9mHQkhyay7b4wub3e8mJrLvcZ5P80nKiViqkhPB7QYFQAF53A19w8bX8CzK
dxVgEmzM9SphuwpWT7nTWU0DVW34HpQ8NH0ZHwzcnAEdouPW6lbZZUjVlmcyvFW8
agqqwVQlYbCJniugn/SYoqE08pC+/u3PiAV9Gw0VRtL9TI4a+P/ECcg2uFihUJ8I
ikqZct/Au4Q2E3wSiOQtjz9UVbSkBshxxdGoYdPdpohQLHeirrHIGUzIsSsgElzE
SPGVxUTzxRRTudwzK7gIp24RMCTbkER1hfxVXbaABvq6wSy4cDBpqskjze5WzJC+
pZY2gFTW/2yz3YIWIcIFrQHsNTxRXuuO0xC5kOh4tEpUlZL07g4KFnzsG9tyS6tk
MqoKmCFqIslrqAy/pvQNLpIO9dqceDmp8nks0vQPPUUgwHjkFM999Lap0k+gfLw5
Zld6L9y3QDmyUxD6D+eXsYgFgmMaIZE4EuB3sI9fk9HJVqTWCplRCChNket2h//T
4A8t23KFMvjl4Y8jpE63AmYa1iTAuiO7GIWY57BDpGYaQ8jN/KywKVoNKnjd4j2u
0ejNx0L+ZGw44CU1XL416tOarD2lc3nBO+lCzlmlWFJzBrXkzD+3qivrqeJKAPiA
I6N6RAIsrdfNrIsRsAwBt8kJO/jzg6a7Qzs4wDLHDwYmeB1/UrUkMXHWaqM+Xtsh
QMlJArLYzzsV6kyx99e00RFt5KI690EBRMpmEKdm0pY1Hfc87Q/u7wFVjongjCC8
hdwQxagqyjOp/itgoYMNoCwJQGDWDcNs1bA6MKYpq6b7gnKKvsyaL4OUKEUiyil7
edWFUGt7FvDl/xLhqOEVEkPSTb94G66bMXm06PxnswdBlktfaZkqOb9rZtaKwn4I
8BPulmT0PguhCMfT1oFq3mBQrJK1/0BxtGpWCm3G9O5ZgDruhBWGo+U9Sohrc/xs
AgOWHWVolk+qSg7KQDtHrkWAMFMtcCc+g9QUvByAehwmkxm/rrDEqMgN4HddLh+u
8smKiO6EjS99Ms10Q81abWGjAcskstq6EUFLAXPN4Ot/W92BK3/D5ECtCTsYrnN3
cl7apG4kBS+TlAcrYxqKBwAqfnW4MJsSlFt1l55GZ5epEim7bp0EYnj6YXDETIHO
bo9csfhqB0ft55l2wCHDJKLcUUwnOfS6d4WnAtfz7ROz1ZqYjTn7wQgJIo+YocZl
Dk97+RzpxPMDFujF3C7Kr6hlgjuJksLyS1H0fAvjpazEfxctz1dTWer0vvXWsdzJ
NgROi1vBVa9AdUuEyqmXQENq3K0zT/Al/zPKBJYnklzzaTHmWcXTO1VRvqSkyasf
qfJbwHJdCFAcy5FG4rjBSBuaU/07rjQhB7h9p6VKRBJ0D4S9ma1GGBdsV18Zto/p
b0T8nClMkvbvCzIjguBpN9EfsAdEHTgx3Y0rZhkzZn8DS2my0N15I7uMic1G4TTI
qhZnAMw8cxgvhcI9kjzKVoPsIIggi4xPOh1CmF8oYw2HbbzRumn8LRw4uwQ8kby6
T93B8X6zg9SY5cjh7MHyFP3liWHAAB62qEftQYI0kvwdAKI5eef3jAhzZ+ddooXO
rNqWgcmLnsdTUAgbWBi746poEkZri4d6A+WAoEkjfZBiyPwX39AJo4kYlC1XjqPQ
ZWPnvEUdk8pGoVmCw06T5GAlQ5Fx1fHg3olESvvs1/4gI7lI75rq2kDCRJwOWxLA
XgkY1oEt6Xy3i2QQnsXYpnIS4RNbS1gvITC1FGkHsHj1W6FSEzXgj5O83Shxhlcb
VPLL1m5wAutILVZdf0A2paxHiJR8Rg0YSFLsS75kPHOVl0jcK/cmL4Un622Ag6+i
OptSPg8SqIReTm507SWA7WinCsjgWU1C+GM8dzD0ia1PzF4GVkXqHbftmT253W1h
+WGJRSMzL1SLVZ4IXxlMGOb2+z3AVystHCKkM/HZ5SCnOVkU2UD10F+CM//1621z
/Aq1ycQbiu3eGKKqrPN36C0Kpu7bHUmgcmFKeFpSQXyIegQJJSUHxIPflU+YX/Bb
E47Qxuw+FxIVsz/UBSK5Ll03z9RUFgDdvl7ix8PGgYZRggqXsvKGjU9Du3+FMoJF
AxG9TyGQQi8KvUPip3ExEfXnRC/X/jzvNVWpnd5USdQE0IVQchtpYkJ7gc2msSWM
YSbzrNIGWCi6iPzZvCH7zf8HvgQOmhmhIfz5p928ItU4D1wnBOdlAAyOQ1ogFgRT
3myLaRlsFp9Cfgy5oK1dLUxpMRxECK8BDr1bh/9oG/FyDdbofbzeZN5cNZGfn6yE
IlEbRaqcnAxNu3iKGRwexxBD9JvVl6JaMO6pyGa0Q/1lOShdYj//i67xg7vhxBAo
4nUgWXvXnVNTZHdBpbaorv0DOcyNISXERoe8oiFxiWBmsya6am25qOVooyG4dfL2
Ai/+TSh4dcBvP5O4eTgW4RiF0Tep7tm0NGMlCQhOgYWedkmiYdkUpi/JwPUPtA55
NeVCLBRdwy/q1UVFl7SpqA6oFQqHkim4TdUqS4OOGEQPV1sGoRIFu5gWm6HMVV9x
AwH//rTsDNAH8KksOT1CNgVPtjD2stlEhVYrJK340rIEP6NnlwMFiRGY6umM2F5a
7azqZ/zLfeERh7dBxAelRwLEHl4e2LVk/MaIOyEn+kM9oDRPJ8b0ena5tq07NZzB
uMXPTSRkX0zHVakTTbtSjyZ5bKmFo86dmsJNBt3I5ATc90HtBz+D6SogXOelD8m3
7DPTSRB4HvuRgUGOgZyEtV7RY9GxLP6esY4j14gAZMeBO0lcf5kmsd2rBWo5WsGr
FH3fTq4BHmhx4GNWcVocdjV/av8yqpMWo6Kd/BNnjuA1oOuxqECYbYGnAlKOfXl2
2XitOIDGdFVA6eavRyMI9JKfaqX/zHdamkKTtzDf+PAZvoo15csS8Qs0Ci5TStVv
mu1z+n+8UaTd7MBV59xuUTktC8GqDg0VIKhK+UcN2rhJ8+4cdwTBGEB92ll4hmt5
igoGXvjsADxhyCt6SQeIhBPfjAycxCIvtL6T5njf+Qh5FvBcEvQI13cs89ox18XH
ZqJTr1TjzeEW2EmNofSB5979+VCEYz9CfTLSeJKWSkb+k9zVZRqkpKutPIOy6uQo
icjzoL02YYlQa3QVVy3MA0Ksu6P8cqXqxL24ENJtum5BGS8QsFu1rcMnp0l3bjpu
KTl1kwmFXgqk1eO46y9mheAuR7W753sJ1RBzGStoZhFt3kSz+k7uD2rAXqPWDb0P
9v+o744E9jkqBuKr1WpC+CZW8w8VzlhYGT8r8KrFde6IjPvsT2CIFBIa4u6II3Ic
N8abWTw/aVv8rysAYYSr7/719L0EMG0Cd9BfniOsR48hY42CWletFyVNmFph/1vr
fN900i8uQWmFH4CS21LRdc6RcPwWrn8wzGVRpyAK1abChcKhkN/bbVmoErwA9NRZ
92a1DwQVuwJqTRQE3djSU5XpKA0rvVz1xlrKpz8svG03rrzngQdmhU5A//Hp4JtT
wQL62ori6vdwExbwWRe4OWK39myHQahT2M67w2OLf2MFsIfEsNmReVqAVzfNB2UK
iJQieptSG2d4Ux69wfvJvYufVHapeJaZ6P1jN0Z22XQ+4hM1j4qOeDBdgmUIzUhf
58StuF4CpFkUfGHFFdtJCFM0iXmaeAQnmQhv1nrfsQcJW9FtC6NnNf5SIUg/Yypj
Q2BntViLIsgrzDmiq/lNugaoE9I112uQqll8KoMzdqZMxTYGi+obEJxG2L510Xgd
K/tRlKpn88gIu6+3KbIVzNjDT0iltEdd0nyLwelpNu3vgVA0LGXiUbK87bhVLES9
KGV5fMWzCpE+f8euQ0tfT6MLcinahKdbAuTr+S1fsjWuq/lh9IywI6rVKhZtxpgP
LRLqjUBX4DbrrFC/ftelApIGIPF62T+Janqho8x7SiXhNry/O0DA1E7WILQl7TKx
m8SYAs9vg96L1pvEgAd3bp7yaGwb8kYxViXpI0QsV+IphPGjYgSuXPhWCc6uzcjd
AwxTwO+ASqwjCz6yn50DgZvu5/Uus7yY/H3GjoswPWqGbm0wfLZumB/PgGrEU14i
/4pubyZNpPNVCGyS8p8ZA5eaAYlJqQCBtsjHb6yZavGFgBypwGWS5aBqor0LoCxS
b1WRz+rXl/dXTWNP8QBVYiHD1ssCK0lxNdgAFqgvELy/Z8Gjkh+VatPrv0iA2Tk7
VQWsMYETb1+QgsaBPjsMogtDM5DBhJGig7MISqZxga3EC9CT6anRlUqzl7VKReff
3dNTO4yWVAYoGk0FHNqUUtHhRf/F4m/l4Kw+vsijcUi6gMXH6ijcla1zCg9ll2jA
cBKcGhbbzjdZqYbwB7Qa0TGnBWoG11OlrV/czvfklwSsLHMA9RgsHOR2GuGJ+iHr
8Hy6gfmfjlqorPLfXBWpvm2hNRvGtGZQq7ljrukdVAsTgAT3h6IxlxZi6x6a5Olr
vpFD9TeS0Re19VgS9ay8v7RO3elzjwd+mjHsB9ReHsLm0vX9Jb/QxTA9TeJtErp6
MoE+kFc712QBi6FrMd04BJ4AcDlv+5vSMQbLsc6u6pJ+4k3jBCqfCdd9ea1B4WnZ
3uz7dgzn32oIo4uUHxYzE3PFls1/KURUkqmArlBibxgHaYE32Y617bhCwqkUM224
u7i/B49o0feYuUoyRzW5zEyBRUT9Gw5v1Y9kSDOWyBgN8ROBgpRtJ3Towh9gCetQ
RPIrqITODgtCBHmcz8G/622DprJzJk1oJ2koXIL/fgBxbNvwPVTMd/KAUNRMMXdq
4zxOy6bhSwEsigw4KH+8gASDfDU7UKGlQr2E4qFQfMnpZWAIRg3F44eWLpqOkayC
1aGc5eJYVivFU5GhOVehzlTBxYC8KvOyI55Ubv+vnMo64RGnzGzRnbWJh04Qt+yg
KjPCQHzDqULL+qtE2h8NpBvignL1bESNKWVHmJs8YGoA4A478UhriEY1M6WQsiEP
l5pVIxeNQDz7MFICADFXqHRukPnJ9L/izarQoLyxvBUeHB62giccfSkyA0GY9jvI
LKPKYkh56i8BccOHA0sv/EjqKFKhUJ+Nt46bZaloAqR0TbijbUr8GPcbIjQ5kCg3
4bErRehKegYUt6ZW8BM291lJA9sX1d8zsAKZhxRdP1reRxSmLsxU40c0pYGnBJ1e
MIyp85D3ue1f5nxhh4IGXobjTqFdXRwv4Uu26w0hghQGk7IMTd78TAuxJYcSmSLG
NWgLcTyDG7pu8qtYm78e0EMnmCTC0al3tvxSa3Un0SorY9uq1O4rjD9SygFBOArg
Q5B4wdCvsnqsshkwCddvBnnG/if9UdXCdEhA/N5jYX//KI4chL3/4fKcvfsvRKjg
iHlc7Y+ea8fqnVyxkltHsCHpDD1hDzGhwNAzkEuriswX1IVvLRMf4xckcEwcvY+H
/54ZS4GVf14ca18pG+zE5qdW65sFprvYnmQTSvuVhxTSY6PkOrx/EySjgVGUwMz3
1UrRePxsLOCtbrXeaW9/3SfuZ51529XinVKqS4zDYEHkZN4TiQ5aPYU2F5A/oCCh
Y1Tj9wL5SgusKtXcMLLIJhQgl3QX0K2a5Cx2Jt+yfZZB8IsfB64tupzSIQrZ81wN
QoJF4AuS+56sXfv4zCeeEtx61pnhiHn8MsUDDzi+c5xxfaNqWQsEcfF+ChCi7Oal
V9DMdks9nUN6tXYecqYPfEpNKoPDUnwzbgIi1/GeAAQSL31bdjUwAg8iDJ9aZGsC
6jBCGqiql79tWXLJEl2r9e41odmb8mypjzAjhaaX9gIn/zEAYE6zgCj+u616jJEk
L3FrFikXbr64WAbyI1iLTH9mOspJ3vTrnEA3R5k5ZtlNgOftp9Ri5QNMmz0RhRuV
inA0uakLF2lh1kHVJYWVGY5rEC4lZaGbw8fex5iOC5KNS1KnVNXPfesOaZHh8i56
yIHsK/ts16BpPmXP5PYgcZFD8icYiqAE5yhr4m2buK7nve59NhidhgIe6kfjRznK
yylGth8uKd2Pu0MU2WR9kpZCu1YvbdskYLHS+6t7UK+ZzSLflO0aa+ecsjRpnesw
nUKuFj9vpw6YQeOU1+SsRK6x+rnrwohpGDoiMCFY/pneZHQ6drtJTBJVoOSMN/Ij
PVw09ym+EUMUDQy7X1kpI4dZwaRw/cSqwLZLPDgQbKIeNTYQgfZ1+RtDaDFAKLvW
aTCbc0xG7MCRN7JDsd+1ZF0X3Eh2E0Y2ERHyEaOw56J4G+E+z10KKRaNFqo9of9w
BOZzp1B4t+T63aJLBXVDPgEK+WbO7d34W7FQtGFTi0zNOfEQBYJdAn91rgDx3FxO
2B4PMsuCMc26g4RdwsuRDCpWegVWGooN04uiiDw9z5EzzV5LyyYuT6A4JI+VHqA5
TiSjIj8A7H/2537T5GmvQh3j4mHfHunoNWROuwmsDFwEjvZw68S2wYXUO65ijCMF
vhizWkLoDXWU7sPOulewNZSjhXiOEBo3PwzBPzWB0BgqF7HlTL9PQySSrrjfWvAa
rAwPzQ7DdQ/+iK0HArg7KolgasCv/4gWJtJICFf7flpO1A+U//rC2XUoDI+13oqD
sEOMQpNel9jMWtPISVceOHg/fwj1uYWy4IbRUPrlmoELhNRiVI6J71eqb+WOOWzU
ENrD0UeFu5jj1H3bbcT33HttVa/Wd+tS3HvBYKrdptMUjP3gQwXuO4ZfLRMRcNdZ
9TgU/fKSPFOYwloSq5MaFFSG5TYYnpD3l+fiBHbEjv2FnDSUVEU5Qk2v4Qj7NEFB
TIhNaJ40icL/YCK4+APhtvDrRCa101cuAufL8eDU+YXZ+jyr9NKeDiDgkZMI0Vjn
TgcxSMzuR6iER6FvUb3BFgZ1peLrMa7JYJ4yMrLYfPnxFfSgDuSWeDECAsF2YfMk
4KHJIoMD+h79iyhi++RglW5dEntFDp/XJEv00K+kisQeQSEz4pGfR0/kggXnN4Q5
i9xeqfeCW1tT0x9WTQ7Rk/jy0OsM9UxWhieksjfzDnoY7cn2lDpPf7BFNXNjFQFQ
WvNxV0+ENcBJjjdxJFGaH7zjhEL+wrCxwHBp7gotCDioIJWSvTUjjiyOxKHrgFKa
OZWA7Nqm+1mtId+yYqUVL+kwc7+WdWAKRaB6YJkkSDmALPUY2WExzadj1yRghUoy
7gVya3R55d7RkQxCCfC+WNdGQec7h8mDYQqUoKqU48S6jxgYLoFu9Be5fcHnsDkz
CQO4d5HqtxuyKAa1EOrRChxAa4i9GdAxLEILwwAIVLjJqr7wQw9iYU+Lggc9dC2t
pFGPfJRICF15H3WMztuf3VtJ85BPJ9+t82fArmdCJYKXpvdn1dlWvGAnqDXZ3CkM
8er8I41lD4AB0Rc62I3rkMCOFrPMf6m9tHjBVIU9vfQW58Vm5Bc2wLUrCxAxL1Yl
2nFm9mAxg4Q9XFywD+u9T8UOipV/kejiILVtuNelO0CdgxfZGZwFRM/Gykht9rmy
+PgfWZ5i88zotWejeGwuK7AgJDiqx43PR60Ufzp5oxfFIvpDuNhIP495ISU7BKs4
HBd0Cs6Ps2hKyheopCoZvPgNo9dHBdOEaHaxFy4E+lrZvClYCCb3KSV4E/5YIimQ
I+fhMq14c1zAElIs+d6YCWWVg7ej54uz2hkCVJgZK11MXzlN6TGGU4sNexJ9VUxh
77LoTdXUqBctQt/7BvxWelXYPd12nCRVhhqI7Uu5JVxobkayYoWy7KV9f0lccA7Z
z8yRu0aQrdd41e+4NZ2wJfMjv2chKFFovefbEso/KcYasQ8+5NUPjgrhw1Ajk2dk
BQ6sRPQmEaTz7jUm4schk6keUQne7vX28k+Mxsz9zdCMrPySVMCphJmFtzVwgQx5
GoZakNVvi+j+PPjW9fbil3yx9bPBFv806n82YmCYbUT6BS5ahg1C/VIo7zPKGlcE
/SMygOpjblxuexjYoK25Y6b6JNgCG0QWbQObYboVenyYr8yrocYV91Qy9XJcqSe6
xA+pwHKU6UFm65lT+2Eb1R1mVG++BnPa8if9EjQWZq/rzNilaLuhosINy0b5bz5P
bMdGfIoO7M213JpbbDWVfjcC6w0oih96x9ZhOJMvx7ZEU1AKntf05Ef3xEe/qTTa
3KWZoQFCAcTZI2jNDpIeCJ2cmqLVvVHZvxA70xd+RyyIjJJON3AxzyrOFoKiN2Jy
9wCWOx+VOnwWSi/4YqH7/znKcJUCMhixsiJ3hbZrcVE79kN1OAH9t95d4MRlDo21
NTfEOMUBnsLty+7CxT2OyXvW/WFF4xMtEmoL2GZCY63Hmwr+7Sj+Q4KpO+a5EzV5
zjKmyxdVHxEpq9Js3RaFIx75IqpETMrvUL97Hzg9kh1Z3qScBzOjpZ9QNhx6dmI0
The8nkkstAZYFr4DS7nI02a9ord6eWw3PYbTxgHc1peeWktck/5U5n94HG4E4Dph
RO9xyJXJM4qPxAW3wfju8jP+zWC4f7Zk8oO1HyciKA3/YpHwbg46uFgBbLXd1Bnm
lbElL4OMtxDSEkBxb+je6U6K1Flc4ZUkZQ8gN7oxqpTmCMLG3YVHrlyVXSRk3MEz
iNa0FytZ9Zf+NlOfXfUdBW1tWUvGnpHNWeyTOJkBr+wWd/kTVBgGIX5TYdnv4Bxr
rBrAfzAAFjuVryHpyIENIMlPZegs//8c02YA4o2eYcdytwEZ5uGJBjPyrJt9cVSK
3hfzxszCy6bFpEbfrsGLue9R4DSz/mGgqPyS+NUUhwx3sqsWs1IfW2Nzj11YIMSi
fL3hUtA4qujHAreZ+wTMyN9yyt9wcIA2c+0uS1lALfCPrBz0aWf7IqK/t5uA0R+Y
/2t4r7SbTPsSkJ/inECqB2CbTgcF2nmnye1ZduEx3GduEaQxZHsXmWY6mbyqFss9
DOGk2FSccb5NH8bjtZ83LI4eHfxRnJpYohmoczk4xjEGp3HyIL6Zi6VaL0gDd4Y+
NwDAkehC2uexLDjA4/mLBKHhjS1cV3/n14WyjThDaMnc5GgzhyPGe8STsIq9GHKL
h4yjy1ciXtW1fL3JmK7Zi5NqBzKKT9Fw3T5CfnvOwpx9wZBjQIs5Fy7vC43sRa5S
p1OK8QGD3wJuAXX0mL0qGZO0RHpPv92CSmibTLCGMQlSPbz3uVY+2eBR7N12VbKl
n88QsM3Hl94HT1vZM9usYTeB+EFqPFWH7Z01h/hS5ssDGiwUNoWYuwWjHb1pBn3D
wExpAPrUUUHbrLUL1LQanYTl3H0dopLm4A4F3bY7DdxOGK1DrC0uNYJsUU3yoYc5
Oi/XUoaECNSGA+H/Ljh1Xvzrdd6lW0w3sApMXnutLiSKFFx+tdRirsgqr2KMUgLl
Yvd5bGw1KrvffkYzLdULnv148ogtv8byQ7PkDb7b1RWpgcMwuOTchlOW6VBmQM3h
gb+xfGpvT8BdBlpJvtrzQG1vduB/Y6ww7gwxTVsnMGQZdv1SlDzplWIyBD519eWR
YFL8xmuHDRhBE88SijFvWzJMS3Y5H0BFAhbD/Ko7N5gbSt4/9nz2HqVHbXdTFYHu
oCzo/cej/XDCOG485Lt9y9BqoVUQZjFMu+nhlCCuX4cS3zca60Lp32vTB7pY6q4q
rrO6VohnWB/5U7bkjVKNmY6FaeeUDDMqdFGLPrkHZI62tidHGHM7PvG5U9473PlJ
bzAGJasrcTUMMMOvfiJzz2U9a3Ay5eIYimIxpNFGHjvktaWKkojL9JVtED32nq0L
cuv/FDz68//UbRVxBL4yp+VR5cUdPUPUOyeT3OyHEefZVQdPBTT9w9GBvANjQ3XW
raEfYb18Ck2jTRgmvEfpzeRFudFQ6XPloZ8+PART9MdMFGElY24GABBNeXd6h4fc
sFpK29WH2smigvymNYjAMh/EW9f9EzLWNRPCZHI31tgkVbv8vIwRoZLH0K1sx2lP
qJT/alA8MUzPQ5zKe87ByrIRGkeytqi2hus9Ev+GoIYv56N1WEo6hug8ptwYipBM
2iMvWrUoVMqRwfafUxH2/Bghb8WGnVYPeBgZm8dDhtYSTzFGh2Y3SXwUjHetyHWr
IQv33jWtowCWgZCuUfvQB9DjJF0ChV5qaXgWkzAlmKI1tH951LSFRlNQxxTkNPxG
uuClkbk06UMSbiGWqHyzMMDqrbo6uILb8OgsOdyXwJmz+WJir3//XTwV5C5MdDd9
LP1u+TsvWUr3gmwyiIKqabkpyHKZ85+kNgoEUMMMi6sdIhoQ5VIRYTgJGaE1WUQQ
jQLDa+0f5xLKn1oxOLSsA8H4RdtkhGPum7uNj1tghMAbYuITTuviJGaaqTcNocSQ
UcokINF0639iR7DHkOcH4OT4JKypV/F/J3tYOjK5qCpbX21zk/kcF66D2aPQlmaq
lzuEJFeIvSTNS/ui9tdtgyxtWVO+hssCMtgGD4QdNULhtj2fmtjaHdoCNxAuZqEW
ZtiM4MPvH4timqM7mIevt88R/QY483tU1rFJSgNGz/WWM/AYosDHpENYBMvY99re
VlS185tQq4qX52LNywpGJgEQ6QuhotQ5pYm2FvYa4gmY6lz3ZVVS0pkCcOFgmnug
/tNeWISdLQBcR6ZohAsVw+Rr90yshWBc05OJD9Qz61MEVjVATQ441jobDrtkGDkJ
LQz//ZhiiXcP0STuS1Xdf2qyV5Y4hVbAb/uMccDW9LNx94y1qqX01oeMOJ65bTdy
DlUzH/+SrMpxqyvNDwLkxUxEUTNYTm7FGQZAqQXCcedc/Vht9/nw/4RWkCAsAClP
zX4thUrLx3G2gJ8LCKarzGSVheInaqPNXY4YA4q2IigxHvcOMK/VEPFnC/u6+MpQ
Cg4vz5gaBnO/I171mBMFLgcZLwxxajeEctyJqIeb3rDRPGkOD6tHSQ1VraLapUwr
0b0eHCIv49/DIg1+Z2SwcoQOALB20tSqvzHpGySeT7xK5vwxXrPR5vDssrW3KGcx
sHJo35gfbnux6AwBujem8se8mkn45QVh4toFWH5SCc32ik2xwXj82jxyCef8+XID
UkCEdQHftH2atyiX7YG5Q8lo/nlp/l48RXEqTFEcqVD49B4wVjtkkQ+jASLPd6bG
akvi3Ri2+ycWwP+KZqBDv4CjMn85xXklHsvt0paOv6b9/qJFw7DdKpMW7rt8kBA1
vv8SNbzjt20TXggqlNzBdhBA8Dl5UDlXIH6JY9v4kkJYviiy1r4kPXGSLYQoxRJc
euB/hGf6w5Z9Dm/K2QlO/ltybMEKCdBdcDl3SkOCU3ozQewEfufi536pJDT3K3zZ
MUzpBP0aCB+sGTXMxV8r745wd7brRfTQ8J1+F/kmznhrNV2lEAdeufULte6FT2Qz
NhCZF+vDu6BICZYHwUFk9Ly7asW7dreon0ATk0siJ6Og72TeAaz5Me9fIx2nZWrw
QgfJRVnoqUxaOp+SpfoJ6F8445h2BiaUUtXvWd7X05WZWi0seVXGU5ovugUQF7ug
ACu2/hPr1A/zxegytE6lcQ3UGcI9Z94VwK0u0WPk6bkyx/Q/P6FPQlWGZxmeaMa8
iArScnYp65Eavuko2zbyEyBDsVpLMPWSjKxzFfaSb3qLmQuDf6IO5VoPtVpJgaXF
U9ODf22RIV2dlY4kOmwJqgbB1VTefuLV1ue0Xrv5j9MjyLpannKdWGzN8XkokaRA
PDI0VsSkG6L/4jcXu+AYl5on7o6KaFJXydLU4AT8hkgKjxPaGFFy1f/Cl5B4WF1q
h1I4A4KsmauT7xXPVfZXnMK/AS3mJN94e/9OfCbq5rkmpiWtaFkIb7WTitK6EsH8
xgDA+0gxExLhFumj5M3w6JhbpCnvZgQ7ny6nz0CmDrO1DPmwB7ykj8rMNET52B1W
TYVQfaCiYtYgeZwgzYSIxp03b6a3Zh2okBqxhN+GPi4FOBFqgQA8VGzcjnO88miT
o/tEgvAvn4xCg9yNgUkxF7VSVnHwG/8q4bo818sB/z5K40CETNCevZWBKORcreyY
pTu/aBLKcS1Cja6D/Zo9rUXOsK96KbxhKlE5woRxLlcQzpc0uAKGdLeO7sK3FZTs
0RddnYNHg5A8bCB8D691m52jRD+VLBn4NXjjyxq/N+EtioNyELQoYXuYKoAd53d5
rKxi2IcDOpZEO/aCxBP6Gm7xz1Dj6jwnwxnhK1bPdSW9RT1ZC7N+jencRKXF2ur+
45JSlmZHDd76Oggp61t+CheorRUyMAbmJKC3G6lu3pT7X/ms0AtnbWcm19Kq1h8u
A9jweD5rnkZeXoLyYcSNOFDZCb+dawXauZWwG6+oPP9Qe9jY2SDjHiDXOHmyEfHS
vkheAXgRYKr6+05kQqXhTVJ/lipDgIrX+jg0b/yNdfCq18CiPVJrCbS+rfqcKGi8
svB4dHh0rIXvmbX9KYe9qojcbNTWAMJjJmIATyI3gKc2jJ77FND4m4aqANQMToaj
mnd7hSg3c0xNzHe5d8azcEk127hXjG9REDGUD8/llBpI9cjNpoOiQzdloVgTTnj1
NvC1kNwB7pjjpaTTwkQgFhkPItts3hE1ft67s7GBNOoKb+MoL2P6oNM8dTAXPj4v
r6+g5R2EpAIFA6FUQz9BrzQUD9Wu7bmiwVSPpxbVNmzqjAy4GJT2Fps6bA/j90nf
KfHKnmBdPPIF9+W9a7smQu0WZ6a9Yovh3hJIoQRXDNktR8BSnKqBW8tWnkBePCer
5OyP6fF3NFw9G3v7tO1yi+9ZaX3EETVSvO9YZJwr5NOIVLJ0mox+PxcmRTD4D6Jn
eWpaO8zy3CeEvkzSpghf9/RNzMxuREaTkkminCbEFwNcfys8kmfnKc1Xbo+SX7zb
cJDKtwuqSY+kGR73p1lsrpAa3PtHuWd4HwaZlIv+oXywk2vnr+D39g2cZb51b7R8
hH2PbIsjlktg0pf6cfzRna24OIEDp+FdMpADImdqV3E6MOwwImJctvLlepO8jVYT
OdsXheNRWJ1P5WcuvPV8wxnIUAbFV7oXvKwtlffSHR81f+Qxd7eFcZ6n9hkV87Ya
jNn+eoQbEp1dnpZ3wCVFaN3L3hW8EGjCI61Si3Z0OZFfLZ6yWDCWP7PwDvITJ2R4
xsAe6EVr60XxNeDqJ8C0EfCxmZFPV1ZPVJC0d3YaVMoXC+H2wWHx6u6XZJxwDmLz
fvU+ihrPbavj2t05nvEA9wY4A+tQvmy0B6S8BDq8X9JpuIHAGXQJqDBsX6MyubvN
IyNXJbvPQH79xeAwxeSXPXFa50z56llzzDwuB4UC30aF1Ldf3j+uUhqGDWIusW6c
03NF9JHQRSD/4cutB0tHc/IhvtgudWkJTAXgWflGZKP3QzYJohmnpLWf7tnj9RoJ
aH8HI90EKzcg4oplac8/iwufJ8WchJ/CE8IU4MYDv5rVsE2VofcQEUumW4gBLZiS
dU1eojKM3pbmPQY4bjEydoPB3rgSelH7WYAqwvH8S28bNDdrGSJirq7/JroOHmiO
fBmmsyO1WU1rYDeEBqJk7YmvTxnEq8lVQHob7Xb7FhKIc9zz3N8h5Ey1r6HjfL4v
TQBQ4s4sMsSE0pE8dKRp19Kz9L3Dyurasqxdzfyh2DfhnqVb0g3yMl1nbf4qSWUK
GLciSmfte2dVGgoBzTfY1SKWIufi8HokmVRR6GIydZ6TyrVLOD86aYdp9Lr5wm8S
EWH6gKljk5igZsTQKEsnPJEEiIy5odV/OErJnK6pUZn20s9nyYzSSjNuTLP+he7D
AsLV0nNN5QgdWk36GeqkTUe81Kt7wHRhUe4DhkG82BqXaok4/FC5RWu+KNVuf+3O
sOVVFVQ1TzVrzdRcsRhRXjLbeiAIaKtc6xhqPORl086yhEgtQAuBQ5ynu79qRDaL
17M2F39cibHsK8tF3yCrCnYLzkMnjyvwDHFMOYpeyFhOK+HxqOJJya7xY5HjmQFh
KwNqh7+rz5q/FkI8/ZsU95XG4WLZgCFppZP0PNfk5sYVuaEixizlkcmTAp2i6aEV
CEhBD6Y+cAh/79bU85wEAXnl62836GtR0VutKsvLmOm3e9DxgUQjczIqwT8595nP
LQYa6zrvpGwZLn/Fc+mb9iTG3VjYAMI7CtXHSXZSZoV4S1g4IZljjgAAz3DfU299
uN7tcBy2c7xtiH+N6miHJgBoeOVATHvpWYj78dPbSRyv4gK4ZnEYS8YWlG60oR4E
rK5sVDx7PV+wwqU2p1bKCPaFgdxz3mt20D3l+0eEhdUPItnvcY7g3Nnauk/+TP2o
pit8rZfgyi+NqhTDqzZ1s/1+SWgzfuLIULwW1vArLrIoO1xOe5bMBzrRh7r+g6wh
Q4i0AmcURxjnHPIIJhAQIURaN3YxGmci4GB5dTEHjcDMilUvxE8yfG8P6qYzE35F
H9JQkBIKqopaOnf568kJa16KnvH/oOFyecO6c8jhUtvgFFOc3Ge7WjlBsROol9fD
wsP+Uhv68BfolqDapnHsv1HjOB5KQogf/5L+A6Sg6mcSZ7kHKvLZVoZo0/1i8NSN
XUhKTtE+u3dRSXMfyqHzzmKSvd4e6tbO7DfkDVAK/N826k4FNYa94bovqIDz+Nao
CA/lTJHgBfywNe2aH+WM323CRe85RwD39aVXCZeQmYik95A/iS/kAMepoot2RhtL
vCkO84pWsr77yyWezuKymti3vV8dfpA88m9yze+TLW6mO3yF7yrHiIb5ZgJqU5Ve
SMORHTYQ1CfVDgI/5CFPizdXt1gipwjBhlpTpfnQp7yQdLD9SJAQ4sG8m5L8e/Yt
yMP8PxqhBlz9h7I2RDi3lGXOkDrX9M6XA4Pj4epsjDhSHm3H0JciMRyrNqDfBogu
iuWzyeO0UJR4AuV9xKXjHN91NkhvG35dhcBGATOJ+RWTORfw1u8n9porbvk9kLK7
TSN5kQQ0jrxVtjDDP+VggAt/BjoehunGdImVSMGTlgYT6ugQ2W/jeDcH+SreBiu3
F26WjDAOvKIQvSAK5uSIFZAcAWbsuuOkg0CmeKLloukxSiBLetIYmwjW2yuhq5/I
E6J12p4ZSrSWeoImmrO2qoWU/cQAC/BKB6GJoZLVDs0nDFQkaEK2y3rVWNcJxOFs
2Di54/Z+uAnYLQpVoAtJN7zs226aQ9yLMUiW3HWfITIAJN1G8d8PgvANuviN4rwm
wGcaDD3Ap4sbaDHx9h6jDFuykDs9n4IZJUK2Fs5Eb4JxlU6uofcBTvvd6+l5PrQV
SiXRWZfPCSktcj11Wf0tFGHUNRgrJDqHP6xAZsUOUcvChGEGUVb37g1dQmSMHoML
5rVob9j1FM2Vt10NtocKpt/OmzlC+lNM+BIWFRafcLnhBLlgJGTt/H7DmfjWA7Vp
j1ZlQZehSOKorZBlsvqUvEak4fVhyvX+6bVCzJyO8ucfR1XzhOhPFHW9Q8EMBp38
ZQ5o5Jwh2hSym8FXwu2fS6lEAYEvm0bcLdV0FRlEqzON9wW0/HOhANSXw/wBl9oy
1DIkpIIBIERl9WuftdGvhs7RzVVk+vSKgvaHsrFYo4+Y1Kb3bZop/m77CYPZ6Qyr
bYEQBE69wwRJF+tIv9xTeRt9k8YHy4ymiGxytzl5I2svMx2MexoCPDmRbBP+2rz/
G7kzpImKXjJzd/BvDlh/0MDBPgw506n4/oyw17JdZOBR89lRD4zIadLrZ1owKbY1
We9j99t2Ub1uz+tcnFQSK+JWEtBoLHQ3PQv9lsVcY2jw2k5QPlKuC+pt8kYIgkvn
IquJrThhpVsMG+l/7ZYfrWMQgiY+y508NcC3eAlVgnmNNaOx/OFpqyUqI3kGGXmf
YEmcsF7fqMr8ikK5JntcrvrdymZhbU+I+Npr/dkG8vw/YLjOuezvjgitwaQJFyOX
q7HB/FCCEtqw11m1ecBYGkLfD183Cz7PCBroSsEY2UbZbZ0Tvc0qcTt8gCGvdK+t
DAo5MvrQuDHo0Mce521oCgv8Mt5ba0gPC6j/13X8CsKxHB0aXP5LTXrvuSRhkKFm
p77E8Wq8OVFxelMvFa0/5vrcuj0FG5gDExDlfeEdd//G7NnVgu42cGpS43w7DjKd
4oQ8J9UX3xjUlEXeBwy4g6Sko/WXIrnww4RQXhsE8dWmcgZCEV2hzLB88eWvwOON
R7yWIxxCAA2OM4XUQVljC8Ev5DvED8PJOS1Ni5Ry+SrQE/j5LNaYrPnLx6dx/yls
Z1B3rCoSyO/Z683ohx7ze7wWCEhfOcegzgPTufSKhXr/Q7d/QJWF7W8VZnx2VNvo
KOhAa12nlsYh7wZohiNFjJUWo/r6onCBAQ3PiKDsDX2H3Njdvbl4JnWlamFY7GNy
LzM4ySp+qQHhvO8Uuf+i7Y4IN+mfDi6ASJXauPFSmYN58odyLA4wfx7GNKSn6gqv
6eslngn7ZN9UTePPoTv2wLg0pF1A7lzIC/EV8xJ7j2BKnqjXfniPM+ALsWtsefLe
48+k8q0mCSSxiESARCWs/D060wGSFNa1JhP10vNb7Qu4R2aKpCQgbW/ooogfjIS6
bFQIAvjcNS334noqKxyk6JA52L4Rl2crMR6YBPIfP4nIwiWvwPe+Z2ZgxKCdHNIa
VYtlrnWSkS2xECf+s5h67VAe8l2GtqhmYyrA7o/5gUt+8nYktxSDdZFPrysvPshd
sUMd8Y8DntgqNLi0twhTKgTPZ5Tme1XuP8ydskTf7aUoMO3dLDN4PYtmOy8GnX+y
JTqjk3gW60VrxZO5S3IaG4fY4BAtm9QgLq5mjt9AsWvXHb+JwNDFoikIjoCT97Ud
Kmzcz45aUOYJmLeItyzEYcLUgyD/1d9PRxsjLZ3aHz9sD4+E3FCaBvYmCvGgT3gW
ByTUYapU/GtAGSbYWwT2Snaf8Y0YRq3Ufgo2/LBMjIoYA2tSc5ElCukUNiJb7nDX
aN6wD+FfkOnRGjR2YhAYT1As0EfzhYE+wnidiVP0Or+BBuFQTQXI2ViDz5MWJncN
YPzaqwntyBh5WtEmlEhKwyTwLEdyhHqkwRvZIhQwkERqDj7Hm/4WJqGYCnX1uRaA
WqEH2QBBCYQ1MbnI6ui5OlAPrM5HZqBF/EDa1JCLgmXzvKIWjDoi+Y8hcQAWknT6
M7KJxIqmJxyfUDFa1YE3CKRcrYkrBKnp1cD8gOFrn045Mnu48ecTDtkR5fj/kYGG
KNunW7ACMUr4p41a9guulqivGvME+kwj3Q+Cw80ujfTpbnLuh1XPpTl1EbvTaHju
U4DPHtW5mUbnFRA8SukcvZtAoHaWUbtZO0ygJfGcy937lB4lkBuEB33gc1j6TsDn
PBWECq+xIIDioh4dX+pJ553KV0FVVbUVEhqqUGaoAhDk3XkIgQ68Gf9QE21B/oUR
dvLKUjCyuKoHivSxbyM0okMIcuL3kPwjYbCogrmb0NId6VIjyaKry5Ziv58Nke2D
dWXdQcc4vHj6isnMMhv7pcRLbnh/k2ku/WnQevMIVWBACw1AD38u5DBwvSLb3e44
VoZoDCql9hnAiDFhDSJswQrrvpFhUmYg9zgsJOgYucclo/f9/s3PxfaTbev825eG
JMdvqMwJIhyj9EFXIhLIJJCcA2oYfPo+GUOEs+oYZ5goFvM0f31EVXOXsvUJn7Pc
1LBi2SlPT/4J668RDtk+ZiTaI3h/RjFKNYfiZYP9q91zFJ8ToTlNxTMKu5z8D53d
HxIeICqQ9iegu3hllN0B9Sf3lFgrZkpt8yDHFPsezvZQ9VhicKMNSRW9iwncyyzd
ymSc8DAqkW9Hp1vCpGXdYiZkZJGVSPYB7JVzEVQetIigJlAHfzFRbYerOf9T8To/
HKB88s19DffZHTeMsl1rkUTZDfSG3DlyGF10CshlkNgq3L6yuYEiBJV0fJMCW23/
trYrIIgV9suF4ZhNS/J8wRebuX9fZ0TaBiJ3O9XC/BLtKMBIQKO8iAyu5jkTExFD
uyfeJ0FOOZFUbUgVgm0GobVW2uGZaxQo4a2844rzyJR5UOOv/Fwog3RzKo4Ci2Uf
3SoddenavnLKy6TUw+Svl4ngeiEh37JGWfMn/0yOOfxhV2xQjBGbKvYg2bjxEGbm
FonoIXmHg5ZpBOC6WZQD1FlIuTUrD0j5s6fj3s0xMdbdJ1mMB3PIGpwk27jTM/Xr
Kr7jVMuNx7gFIuXbrS9RP3T+BcQOjuEd0iCJyBwwu9IMbsrRJ/cskD+e2pn+RBu/
2b5GF98mwAUAI/XDfoW1xuvVpVClDmW4H6rW/8/fTynYBaJpl9cl6aLnwMPLfsal
icF+SBIB9CEp1PNmhOI7xRdV3gm4B7YFOpHvKk3M41yXoJiBTO0JyKhV4aDbeOzf
9oiZN+NT6RWcz8HSTO4OYM2RKJpPCpxCo6U+kqyAtH0/q0iLJWtfcq02NJwD2hJM
mMvj5g8esZIwPns/OtsTQx7n8Tay47mxi6EwZ8yAl6IWFDsLuapguEkWZ53WU2Ya
X08auFK73XhWvu0m8Y7XeovAGDh6rwJD4amaPk/62uIyVHIedPmDnZTNmRG2NnDm
1JqjkbkiZPuVfrUkUm8txh7Sk+F6r1CflcdrxKH5VBE7HBr8pNEzMi7pN7ZJD5kF
zM+bAGoyrbc8nvLbwtLqxEsxN2Lk1qKAAEBvA5FW4VcpmSuOE8MNMRU8XVGz6Q1F
vUsxzyEWuJ8W2iChSUMK4FzlqsgSofRYMrxf6dQr/8BF26UdvmJ7NpTZpCc2V1tW
WedrUqui6m/RKU/NsoH3yd4mEwThFkV99P6mbJAHhSsKd6de0Md7Gm7tRshCjZMY
vVIbRwnjm8+8RF5oWF1Rv9akPuETMGd7dnmWkEcO6FzIV5jHKd0r0qbhdmQFx66W
j0UMHAjZYQ2xW+xhhLFUgUHAxuJLPoI6fYDT7t5+cFzktrbUSIZX0/Nn9N9VoYno
WEjbOEr4PySNiXrtehmVCsoW0v74WI2lNKR8uhb6d4RqLGsVdA5aqfuJoYWT7TZG
2jOdzTKls0/yKrAEpaXBSPTN7KSh8UUeyrswwThE0OcaUks9oJV4sDxtt5bM07lB
HpNFvYJ5y9LwXelMSIGOyPOSn5h4LcXDwfPkXysBc6sJhseY4ITEdE05/g2/KMWm
DzIgr4s+j7H6L8zuNHHJqQ3VPIeUV3s/9R/0qyIX7PIpMHD52h48/iNy2i8TizHk
6EfulTV2JDNje8MwGAL/bQ7W9oMVgwpHDRKvDUauk5xqQgzVwz4teq+5PIj/cKEH
DGlJT57nLrqNEb3yjSWh8FQu9vYgG3PaxEVyyaurY+E+gryzowVlqrEryDoV880+
yE6/4r5yBjoV4tjm5wlkGFjc6kKZ+0kU9JcBHPWgKVNYvbWKM95p5jFhJOZ6OWIe
TKo4aUJZyh/U1AQIxrgC+zuJ0ssnIFaoypoHFMWlKpDyyPxdV0fdXrqN/rzZqWjv
eDsY02McY1VNxlzHYrawZWx1uQnxgaMyowvnI8Oh2nxaJZsyFLfCsYpTxP8eSX3L
`protect END_PROTECTED
