`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tMbCcqwwqrFz5tOo8sFhpRwGS+bbukgrtz9cjlcNFwtXdIIuaMgk926vBafy3wHe
pmG4dIr5zjJlqzUc+KxhTPJyQTU23w1VlH4YkrXOajnrjqmgLh+ZKTb6NVIityok
IbCn0D7M44xxTVBcOeV2FbQg83Ig7IIett8ExKZGtbA5P0fC8tmP2aR4kZtrz/ix
eBwqbsbFqZbA4WaMJHIJZgfjhCZqY++qLD+o0lWQuZrJbMI4hwGYmZ+avw9Nc9Y9
1s7teLfIryQsLZNibdz7abxvJNWYdbwOOJH6SWzNz6XsZY5jLNeFiDa5lYwEelDA
LJrrsu7eRnJtJNSZVgRiz2yGF4j3TcYl7WY/bTPiRX7PhVLoGnjLuugyC/M+H/tQ
bz85ILPPfHAGCwoGDnozeU7uiE5hxa9+33AAWUMmTtf9IGu4lQKeEphwJfFHYmKy
aABbZgvc0CdpeVEoAfstx86rjDBuEP9aE7O0VBIpYtS5MjFqk1AY1FEIJu6n1MVc
SkYVSrTdybrGrWS1n/yAZdo4JWajwS/60QNR8N8ffPTg2JoC5kg04Z3D/kdHLGc6
MaPtp1OKLBR6jISHou/1snkIZuq8imhAyqps9SmMwCzbOljKpa+KsNHq6JwI6NeT
OAPIwuiZgNL6w3ANwxFjDYwGa6XfnpBNpUJvL4O4ZgyDqqh/yNa7+6Rk5eO6SqOA
uz1dAyAMfA6HgEJInAyovhRzRfMdTyG5Suv8DlVnkT7f5i83UvFSU28EjSiD5cFK
QCDOoMz6r1ONrXKExQzROnGb/muTwHDMGh6VyskZtjjHH4WP5oKij/5lbHskz8ph
zy6yELr7b1EHACMP6Itdbet0oyoAgxWsn4RAVy/77uhJFreYySpc/jW0wZ2jYhc4
CRNwT939BFQQq1jyS2PMD+4RvNgI0NBLGnFUxjbEagPEhYVgVqxJLCtiQ7Cx2CNu
wMXIjdD/hBnWu6C3jptFHlIyFXn04tPU70SKYE0lc6w=
`protect END_PROTECTED
