`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZYX0buQBOvWLW2apRAQTNAWCdnMgSSNCJwLnxT1djX4H/7IHIWlKVjfe7W7d7dp6
5p5ImluFUdZzwoZ4Yy76jAQQIcZuCBsYwPv7YdHUgUKLsaROFoL35LfVLNPDZh7R
8BsQ7Y598gQUnKtNLU+LBKnLJlPidt2Je7TGuOQ8IaG7mUaldKopzs+mmYHcPgwX
x6pUR4UeyIYRvsu7dV/Y59c9B1GFpuEmVrOWn0fNO49nA9LHHVFtEz7pa7PBKvNl
/UJlVGEP5DNXluw/MyU3DMWNqMYQo44anddf4Unv3/TflZMIsgiGemH1uc68b0Qm
rPoJ+luoiw95MDcXaBWgKsWz6cSBT/4pLDeMq3gte0+k//ia+lV3pkQX23jdALg2
Kj2FJfGB/f54hm/6ZCAFy+0FT6lwsK/pjGB9Xxab28QsxaXiwI9Ys4ezhe4mb3Dw
lm82T2Bc8sfQbGEc7QzqrtQGVEN8hWbk1fYan53+CaJ7L7dVvhdzNtmJKBAtgASK
JONkAzgeDUGm50FN/RqHibals8stmGbm9clJV+cIwIBSgwpbZn9tNM27BzWJC0NA
TQ1z4h0K/LrtUv5v1VxBrtOhILmJb0HGWGIVxwn5Cr2VEqxkSNChy1kh1mNH8U9A
K8Fx6kgUzwasdM1KU/8O808eXjdBdSSbSTkx9Kq9EBYfVyPNFp/0WQ1ONFFTvIP0
5CFfk5YWBFBrPfFUygEL5li5tngTHpYMaFeE1FsihGsR9JR7OOLeBSIWQwiYf5jL
7Fs0DiMF8DMc6ugUswPXDPq2v599Qw2mT1X4wayN5H8Vf9OMzHepMFMkB0VdZzMD
ao+xAtZMsd33FQEP89b7MUTS/N7ifGx5JzpGc8DhQ831Cqq2mXPetB5sCPA53fLo
epG6yUOt76fY0dx+/sD+M1qpp/MSvAiixsfaN6kV/SuxUqIUvP4ZRSnDuBUyw85M
HCnBxgpo6K/6pKvF1LbWZE8sGwTj70SZg+4sORAgoytUb7CFZkRe8W67GOMw55MX
BsdP6YCfPdMooHR6+hRtgQ==
`protect END_PROTECTED
