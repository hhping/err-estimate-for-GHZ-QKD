`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w6HB7dk3VAl5t8lGqg1eTdGERlykaXiBsrIcw9Ud1neDOuJ6kYvZLPLmOZqga+bY
1knGBJSZTyAEJpf7Ir+Kyns17Bo5tZ79SeqZWDz/UpmUWS7mnHIjyf1v8BXJLtCp
bfcnc6AGAupZejAo2vc3crE6tkgi+y4BVjlQaPnhqPoGHorwXBXkej9uNOalNLai
DkwjG20z3DmY1j2xoaetuAbx3KCaGSD9koXr6QIPSInPjBtk5CYkAVBe2TRx27Nz
ptsMLw313cJgZebI/5agpjHmdw2TI4CA5gwhi2eI2Pzry1nDn+QFRZ5clbmkIzHx
PGzv0C7K4UOAs9YNIzfQHKi99YflFF4OxqRK3jaf2FfbSDaRqCNyPywagcqeXrXG
UmR0ukGxsn+zfjMdl0VFrCRu5OjLZySnWgvsQ8WRKmWzRx9pqS+X0U5oMuHXmusk
`protect END_PROTECTED
