`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E8pGZ+uYv7DMRbPb0jDq91vjCm9dRjA5hHBCjpASaLYq4skwGEK0JgvrH+bVt1BH
k1RIuegoqxlfqrRNYjO2m1HJq+oSYraDFGnrYg4w/eaBKetJUxY69uQHiOlkzTpV
UQ5dsnYiM8mdMukHDxPgVr5aKVKO5j6he4xi7+47dyIT6SnHuBdoD+yAqjGx+26I
bgKxXHIhFjC6Cn8cZCLI1jXMm6zFhBst49UG/bjHRbHVBJXYbPOcMVKsmolxvvV8
dz4liuNziwLoxL0M3IsAUeyD3nFksPp0PvEQRZUO3dDcyoSfuZslIBZvgrlZmjde
T7ynjmgBJ+G0aRa9kwyY1mW9aGjrWpYTn6KjrxK3cXqPGCPaGj9N0PZp7zjFREsB
d/drYEgVs1EaP5mr5im0TkcEkwwzyuxlfC0HZEcc0BucN0PAMiTamF/+BpKtTLBt
d6JIJ9lAetnXlMTs+vIyII0IFXr5WIlD0j79rEytHUnbRQ1+yUEuD/3LVuxusvNI
fzZlS29PiKlmB3FWyiFlK0krI0pEOYpCvyL2geHf3PwGT+MPIsCZg414VVKgDs7C
lyZBPe+ilE0tjgc79nTvNf/0Dr9RV/H+0ihSsMzUbxehEGD7FQBF/1/gDX9nt6Yc
4pOrBTcKhxdMNBYmnpL5r5ly5XbKFAGm+WSx+V/Zpa1m+d+d8xChP1XIc8NQbgQy
dnExP1iN//00kBVWThXXhPOMQySn1bhB+HyTu83wU8sY3Mypy7YPt1Ju+tHDh0nT
bdgDkwF3wZ4r5neEWZUnPqj1VQZnM3h5vzFmx+KAxR3SG0mm8l7Arbzb3zFStuc5
1St5vwQKdFjUfnAFoeXsm8LgOCoV+X8Lq2y7F91n+KeKZ1vwH8mzAvB059wXYbxV
aLGxl1+9WsZRuWXIkAf7snQuqiP1DCxNwE+MsD7ILABqZj7Le/hAird5OQUFKwWu
6qXe0Snxka+j84DJej3t/owaio5KMLMF8LvaZJhwgZhWooWEwd5JY9fHNSybY31T
mhVlvFuKu5bDQNga0ipbFSqVN9mEA7uT71fsiA/YjHDTxmR7r59YZGoqJwaSBudo
bHTgqzaINS3XMOe1mNHFun9UJP6nJsl8OV2Qrt3Rn7zCLYL0pxi0N5+wIwqrM9g1
8tRWnfst7730Vtr3QecoihA+fydEJ85cns/HJ9xdbLx+uh1M2RFLjw+nVZ3RDHuo
fYgF3Z2sfbM4l+G5C7o8zD9cYdptNG7S3lFL8gJ472LWD/o7Ya4NkzWbnrTO3Z4K
O49NALncCtd/0U+xFMXECOtx6c9/mhedYcn/E9VO64lQ19XMqGiaRWY5PTpLhbfL
U+sgojnOjgUxy/wu0EgHJTAALK/iXdG6had7h0EDakgQOl1arPpvPlwIozrh6FYS
vJcTTZep4zNzyou/j1PucaBgIXnOD/3mCrZQmf+mS+vwJslXKrdMdHh2ylZQP1BJ
sl7r8eIO0tuKZ+eBP+Ae5VFhbEsTD8n9zt4apYZ7bCsycsyQHCLY35OEWkEl2Gea
De0FIyoxsDHI+RQlI5uphdnU0kp9E1dxfA/vmPFA0rGZAT+RBAraevP27XvmNXl0
EeyOFprJ0E5bvquEzD+fFYgKVJbAOAuD3ISRJdUpSOFmah1LL/jAvjTMz1L/w35I
NsASrzga9sa1muYXiN0V0S51HP1qw9bAWJcasFNqkXkTBscAXdqDBTkAJV3Tcfgi
BG4v+tN6sqOpnxaz6mSisJb2ry5Z5y6M4poalvRmFMus/TKqVlpCTm+vlJgyvYxd
lF4VPgt+XxmP55vfRHEwX/TB+uZLZ76BlGy0KkHLBk7tTQGVR2nm5X6v9pQxXe2x
nFIuCTS+IkwqTyfg3MPDAAV8gA4GAVcFr5Hs+8EOkeXdmzs8nqAbKQSoy0r1miqa
dX5r0CuRl22mqCEG5nv4t/1OH3i8TSN8OnGvDYpkfLOCNZ3/q3TOXjY2A8aBpiYY
vjKTWDwkYxUwmvr1UAv03X1Fp25hk/bs61a9a0WCwKyyEhTxpRU2bYaROwR8g49C
+UcgN7H3YTSpdbJCwsdfreqZdGByAK3Bo0AMNHecYm7218zUmkbX58Tp09nCKfXl
aXBvfjRzuTI7DOxb0Pr2Y96V17pW9jxOcvRVeIHP3UbXvEKl9rQoWlnIdhaJELRx
PTGIH4G9MCu+ngNz87/RHsIOqT0NVO6wG3N8zkwAWY/jCRePqL/cLPDU/07B0OGq
OL9oVwS5R9zLJaY4/BMTl3FHgAJl25WohUtYkIpdpRlO2q2figz8ck2yPRkZlzCM
hQVGPwqu7v4KO1fB6JdeauF4X0j8Q+Ipxq/+vTMCEnzq/TYLLNh7eJCHsbzRNQ+8
`protect END_PROTECTED
