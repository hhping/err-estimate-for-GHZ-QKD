`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m0rUo0AegDBTmX9M7vUgIk8xMddj2LCXXwbB4ePEZi1PwGlQ5C16hBlICExdTaco
rA068tK3dzr4jmVrCEBQ0D5EPHchiAyYiJxlElHSv53rsRpfn1l8MKycjdRLjjeH
0obtvux68LwALXwx6xoJT7JCGUxenXOBDvhA2TZrEWP1508PbpEq/b0PB+zHb4KI
lq1nXPpPuR4GTxJjUayZ3p3iOlUgE8PoNhD1CK30DcXaVUtwgElxqtXEZhsRUDQ6
CsgnSrewX8BomFOO38OAomuQhXQTM+NYKHsMlL7DItCwhYgRvC2uexujDsxv2pig
yfGaDVcr0I2CGN+YuVysugPnT+fgQcsOE8a/HW6zaGbj0IjYx+bgAayUOyfps58M
4phZNI2We8jwQAxniuWIrm3dV8EFsgzqfaJrNrqo1XN6z+QRWNHWjIG7Shbg1Clh
AvB/CnS1ronKhqZbkApzOKsTz3QQObXGdKE6SDj5NF23nF76+V4wHHgwa8MPwtbp
XSFymzcWJFeED7izt4BDRvF+KUG+FwSzhGrLWHdIXUBwrikzGq80k0zaBk6RsJLc
39QS0oOfOUJ0aKjKhId7OYXTEaVuZ4Gtl6TmYK5ALzfxpshTGehN8o3ATYUEC9OL
9gTjoGFdkb8NEEW7eO6rE80O+0rsMfsyMG6ANKQsySkf2PyGV9V4HYM4DqnEaqDB
5Fr+0bLe8DP0g8z5CBewzm8CuubkxkF1WzSiLCJFPcKS2T2kLEjUDtJucUPLzh07
/bmmGsswRjqGKajbBSAp07g7Y8Xi52/Q849Ai9322KG0DY3lpT2YrYSBGwUeTqTp
kzzYBu20TGPPgRnxxAa4Fw==
`protect END_PROTECTED
