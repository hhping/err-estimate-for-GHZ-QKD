`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pu4aZhjQGID0z+R/OoOM9mhWgU5345suaLxbuJQVK9TRJSRwHZOh4mut/vC9mZnC
KZ0f6bveNkCXqCXWvj/c9JtrFcZI3ZYBkcYDLCtLKLW4XpldmryChKXqDvyvp9Iq
Hyz+/Cm9X+QWN9DQUyCLjYtmJMSYB0rH3L1pFjfx2wWVy5BG7EPME0SYPJLryeFG
M7Zk8Cos+leSBwAcBGZw+8mnpe0Wtl2LrhHkw/nPzVrppfGsWXQsS+/0f9QzaB9K
G40pMOZPZpYQQERxrLyvkQB673a8dhKoyN3TQIEaxqf/95iZ2vsTEn1Zjl5peZsI
MqY8RVpD0jbd76XC3435dthjU67jtTPZ3MZIu5txRcX3lMD92h5+SF//d7V3I5WI
hIvemfJgCMbYl+uxrm7YjSmIVucg0BsYbUJLViYXdiLmJFWmyNS6AfnoDTeCCZF6
ZrSNIK6ZMelxr5LaVMlE3cnkHEHEWbSHnkofplD3qCgqyWf3y3UH2kbTL4hvM4f5
soFHhRbDAIXy3q0auxLIPTYCfKyaJ+syg1GpQB/obxAyGC+lztMft0NVH084/zc0
PqDOsa0m4yJ/WrBS/qyuoB43Vgub0D3NBx+taeqjypzyWEuntij35Ifppsxux78z
8VLS6za5uTOUHAaL02tK+4FO1Y4hD9uEknCVSbQ40Qc0JmQCe64xZWUyT21F+/h+
AzjWfQqh8LVuPWgQNki5DmE8BEA4HXAprkj5znod4HGnuan0KbsvyGtkaxYvZy+/
qe77ZcVguqc7A+rbotuiQVbxD3pWRUUpXQU6tMIOoG3eV2INHc8uGh9chvrhgoJd
pa4OJ8mKYJkxZnEuFiZtQpEtomS1w6F06SBZA23Hou4bvhJ3UeFYi5HQFe4g7Fvx
RS+E3xgUa9DJ0hD5B1JmbgYAPc5G6feckJRP0OB97bqHf03bSr0Hsdijwl+6gzYn
cEVi/QTNWCLKQAeO2g/kqoL+l9ziSawMc7Y+k9nOTHypDe3JNcZTys8SzPcQhKcG
/N1lMNYBLUYsmKyoTGbIwG8m9/fBQfLHaMhhL0ts7qXZHakHIU1tVb8tZCbUX227
gs1J6VK1jgJ2VPqDAFS7wQef0qV6T8e4HmdKEK8DfeF0Ls8jzh5LsOZnBn9Gg0oe
f2uw8wWSnpOEMWPh3FF5PXgM9UI86lPrheBd6TLF2Z1N/iXs5z5Vo9px9O6zokPJ
`protect END_PROTECTED
