`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sJpFFB0J9VQI5njm/jiqsv5LQnDknLPm+dAx4KWcgRJI0eUQiIPBCPs/xlDyZpJi
RfOcuubFH5kpW5tx2dzEaMV/E2Ms6LFCigDbBmKv3nApya1oPgxcTP8eTIM2dcRX
+Qo+HADGzcZQEknkMzuXqmAQ+1XuMW3sION2ca6zrL0IFefvSNDq5lXAozIGFsmo
jNheJY0jktuuPftvvotBo+JnLcHl/eyXY/MukNb3YoI81A5eOCtWaH1umn5FVykc
qX0V7Nr3Juf/oyrYMZX1CjEQbTOdd7ij3+8JN9JVovdLY8tKGWju7i1Tz6Onh81U
4F8Bf0lSbfW93q7+Ty+cgNghlI6hISlfkGpLWVhcWVMJg2MFFetA49tMw4KmfoOQ
xPsKpoF6yap7v1lnEg3RCQnJK1a1pWj+fkEarOIYGwNYXCz6yYkUG57Iec8EEmKG
0DuD7FaZ5hpTK+ph1oDIi5aXlWHwap3dMmlBwAuz36Z0ZLYfSWiYyAr/fFitRb9B
24hY+sv03iEiXZupzXmlxz/ddR3ZS6cxP3ZzI4YUD+CPfnwDTPSvNoqyGZqR1ceL
`protect END_PROTECTED
