`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9GXtT4Vr9aVkk9xEqC+c72f40/sZEIPBHSCvqs1ZEOZ4KKE1rGTWIfgl4SoyAPQP
dZPp0b31AN5I2gRJe6UK39kW9Mlt3hWg/sxgfelQ7pNc4AU3H6NbBQpc3G7GcL3l
fexerVIFXDfct4JXqBjveV5bKN9u718hLf+qmgFiGO8u0HcgDYK3ecxIKq3bF4aX
5Hm56NSsAK/Iiwp0RqB6b5BXtqM2ll+JJEIQAm2qX0NdYVJkLLB07ITuVDoIY5Gz
EEVagKabFuWGnUK//jRODiEbXti9NDui4ETDLLYfW27vNXKTpwUMiaxuQRj1eh8M
Y3GG0mQAUNhsafJ6WsbKf7pynka2rH53WNoyNv7KmvNhVczM8UYT9RVaA/rvy1yZ
76eHsMgLtOpXCRjSA2VYlV6z/elV7dNFossqd6O1cLZnYyqIqA1AZ/dJcJpJT+wN
HYkYvI+5mhQVFFqArqSnn/H1Ps1xw1bKjiz03sElgGJbmA+GgLt+US2ScfYV8knp
cOuAumA77rZytB7AclZ0btUR0ilrVcX6rpcSBQuQj5U8TVbxIBmzT2RS8HsaTCuR
4VxEQW4Kg55Df9gTrN/Law==
`protect END_PROTECTED
