`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f94q8pDkSXKStdz6des4Ii1TAN9XQREvlbWnq/UmLsvcDk8dI+ep4xOzt6ek6zWZ
ciMIqpvIClasWBgIeeEWTmxBUbjEvvVrViEwY0nArT6TlXgk0QHDAlQA/nWOx4Xz
k4LhAZuW/TmB9CFZ07PHztqWyNa+ZecGi+b0KTtzxIy88ZmfFPqcQpXDOcJret1k
M6opFZcK6wIN4R0GQfcVHcbpnvtM/xchxb4nRflpAXYW+aznp0oTMJljX37EX2FS
xIhVH+AuhmaCakI0XZLGeADQFf3eHJNc8oA4SHdO2eOFHHqLHRRVxfJZoH8Ncm1x
p/0T3wtruLoSol23L3I5WC12cR3SHVHGi76lEmnkyp3ZDPwEyljaH9KoaYh3DkG4
UNTAbK6VHMKB3hhMFnROtXvMtZCdHMKsLFMuwxIgbfJBhssVStnLBcTgPAR0thk/
dwcsk5fxgwVuZaAmqOXB96MkLFRz0d3YsyS3AGWXwaAn7V69kUPR3l8m70+IGEWT
`protect END_PROTECTED
