`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QctSJVqj1m2qg5rbxEKygwxEIlXt6l8TQke8HN6sSGuzyz6r+6V1NmMO/xNVZQpt
A0nqfs9GCUFvEx2a0MG1ji9rQ2VTDJiufwsyPob36S8jwA8MAReEchgfP4wH6z0f
IrNCV5ufJp8wSfKBn8BkBBTLldUCOxX6Jlb8+qZFic4L6zXw1UWs3HJF7XU5YQdx
6qCLIzt8vC+8nsAVSunbYei3Mx8wqOttE7rJq7p/MEJCnXUpVtCt/4+2WDR9Xd5r
AUT4BQnhVDGklgw3O4P3F3aU2807dvPTCXwuVtvcvkU9shX+LQuMvpDID7yluQLJ
uM0z/R3o1sDtgUy7+eX9Yj+76iRxEEJw0U5FUCSfP3Wp/SmXCGTcSLtuJU0D8C5o
U1GfTJQPMpuKFfDouVPL13vlWjbZArJIaoKahNDMP7rgz2jNtFW7/iXDv+NsYW+m
9MmRmKyLumPeZGfN91h0WHJ9rd38Lbb58266OXfJlB/FGuaFcsAt1065uuwNWsaN
EiuwtUvvpD3nbZs4kTIbYdE0NxC5EsUuBXWFFdCfowKdz+4o7MpcjZ1SgjZqru9r
U9CcNXvgig9NrgwOWxP/85OOHYcIJiaeTHBvuuwnlZdZAJj6MjluNZUIfZJSDZBg
/snF7HGgTUzG5f7WuylQMsgAbDzRuuGJIMbEaHKe6CXhy9TWSThZW9cjikqigC9C
7sIoW7smq6gq37LSYfaYYX43LSs/4ssH1bUHdwIA/g/kCNDv4uwYoqur/ykxapaU
p/cGR6mWdi3PrwSWeTO6xqHMTeKvuPPasbcJ8k4E7b3m6NPMKBuRDNsbOQI+a+A7
TcCB9amcd8+UFKzdVypEeiWWLZj/BnLsojvaTzUhwN4C7tr27jW80tGwPeZclZRQ
oBb7n7tCkDKjC+iT3hXyf6s5PjGaH6jAt4IHMh8kKFvs/5CVHvNdnDPjattVOMxt
+NohD4ojkjA0XfUz4IyctLz3Vtz2sgGbOBIp5rS4+70ovTBnJi9p4G6uqxaBVoUE
JTy4FU1Y5H8QjoAbk/IDJ/+X+v5jj0Dv61fl6f9nb88fVDJYPz8EtnIhndp4YluF
wHsqP3Uf0lV16l32ZRoNOoViwjo0EL597FuTVBgtnmpN5Ls0B8KO9BG2DvSl8k+u
aIEB0/MGX2dMsQoKTGZ0IhRxiuWvZ1tycSKOaWJfFDaar2zSOp4FK43FMsufAS3n
+/bTjNVHpwOgbrDltBk5TgQO10OwQrpPHwFiekMUEf+ZXHj2uG1jjbNXN0UWAfkt
2tKYiHrk+ik1w9EBsHzLwyprtgtbmDi7/NG0Clw8cZgtLj2rL20jrS12kkRSjPYj
N24BYk7VVHdh6eqTvyrb7W2N22hAa9H7zDUo3YBraG8B3k/ibGUTACNufN3fxfk/
2e4vZWxb2zyhaB0URigc9n2WOxfaapAkeTHNmoo3ErWkY8U/vV6YLq0B/oNxURo8
vPzHuXu1/PjoMj+HYxLcS2bC4NZ/REJO9omSmEQVbNLIj7BgeDKfiMRqM/InUZJ9
7MTYODeNDIW77mqHri7Ov/FxyjVrDiUr69MaW35Qi9qkalWg0zl5irpKbCh/67Gn
g0hmrGn816LeFwx53TnUXRTsPrSsDoa/GWYC7l9vs6PdpH0Tgawotm/r3z5jUIX0
61ZMo4j/nfIXHmi7GC47BA+qB/cevK86gDHQYSWggpHHytcDqy5YucUbEwpucYsA
dWvr/H0CBavb+f+lEMQKMYz45hvH/P3bofmkrEj5xhBBDyROnlSaH8KqJoHETyyw
BNHHheAhun515aNobPn6zmKZBABu2ksRRDXjiCkPkICRtahxmyMbADA9G+5xvZML
QciX2b4KCfEeYiWVm/a3APCpBFb/5Br/BeGCKxmF8DqFLkiBjRBT6l9iYtsOSsaz
MS8cO4vCTkqXHzr2NnF0vr5HB/t1q38Ge414aCGdef/cfNtLLW2rW3NJK4N3LzIU
8Q1/e1unKXUB0R07nAdAlr9CoKOXiEWbrHnMdJcnAyrLTF/pd5tqPE04S1CyqVQM
1xFZiGms1nB3aF4JSMlS6+kqJZjxbAsbad4l0h7ceNTB0a90A0la39Gne/t9WZoS
fRoDEbW2+RV5f2Plg1ykwNQzfeu4hOh/M1qTlE8CaZo3IYGKEnacJOkqr0BpCC/2
VqMe3jt5xy7eKLg81FDXgOZGDJH8braUm9VMntEbt5vFy28YvMHr1NiigXqdO3n9
Oa38fJBQKHCFPylht2opL2PSqv9a1jcaz2XaWk5g/fb4TgkI0bOkYotO2heI3YYE
XAtCr1KRQpAt1qm4hqVvo0DeWYTQSgKMa8ABvqg+FTXW04e6Nj2lvhT+uO7P8vba
HmgKCmbOArmZDf+MSNompQQR6296r2C65VKL54dGeocq/DZKm8x8uout6J9WgsLT
55Rm8s9pd40+RVCJvuxazUYuj5mNV90ODHX+gEb3XR5z2mEEh2G+qCK5ZafQYIbp
xC9Gh52wdb+iT/7VzQHRzL0dQnIkufTCkZHlS6LsIo3vRhZjFQ0vR51pcgiKavZW
IKHUUa7+nyheqC/ejRxqi8fPY0M+2IG/FjRnwvewx/uEE20UqUpnj3b2tRFVulgV
BJBeFRMt725bw6PyZXDbp0C5kp+lrR/PiAfPdSPJlqMc4DIXZZyGhfgDsVpAwa04
akBAQwpZTwuxo1Aq3nITPwUt+vtDRkNi/gp6t8la2i/eFW95gbPd6hj4YiPws7Pe
AnCg8NvSKHagnkhLiiFvOerNvSE7U5KIasZqBmc2cz1qk4wCaOsGO8HOhNdsPnPr
rEKf4WqpdoPku96ngfLLjG2F/9BZlTNU9Ix4Y2QCYlHUiPcLXZAOJ5H77wf80PSO
ymBgMDibzVJCyZ5E2CBOZKCq9Kb/SkIJO8E3JiCouHlQgPr+rBFp7SLYOo3LZuWI
ZhylBOUtRVaZ9f3ha4Or5wY5Yr5LOTwFF2uS6umj3SkNP/ENM2ZPIsy9iwsV5CLf
M+EgKZ1Kgjv55PukRkTZXHdZScijdYAhP58t1gETsm0rqEaz8bwczA/8o4ryTaAg
7kzhtIUk7B30lybgWp1UdcO65IPiesKj/OTlNtJRrwiGQusWUyqR+0yyCgpGwp8R
nPZPNeARVdUtQt8eORggN86jDgNdG0qUT6e6oUFmkE5lGZpN6R8g/ZNnw1Rhv8ZJ
kEhWQa6cPiNfLlGqIcrG5BVtKDasUOQ7/N2t4RXfQ0c9qCyUnFGutl9zmff/xK5g
X6Oh9sE+s4+iPof+demh6LlWY2v/IOjUQzd4MeThB5iPCk7j04citwSOeDY5fMqr
kPa+Z9TS+6qLFtnBkDnHEvdnc5L4RGVQNSNBRFsMHxBRxKY2qo7Rpac/yfSrguqw
Gldi3UxBhmRyE8+HR4iITkJh2QTJg/v2cQDD/XWkfq4PY6RBVC6e/UUWrDs2fZF1
wO6Ls7gWSjt8Q6FRBA2l0CyDYZ8P92ej4q1ZQQhRzrDmA8QbiJLQW3lR2F9w8jNB
feF5V5cfXbi3tUzm/6SFxx5UOXPOxwWETr5EJA0SZcuBgX3doCaCywUevfXhkdkV
82BjM4elc1zjLJUK3lZsmp7fZ2BTfcc45uFJe5zbwTZnXmm7nlcqxQIUj8uvYHYv
kuqvQRcVWiGSLDHbdWgOC62VkcWtwtMPQ9/VnLiKL1C7felhKMbbw+PxzCYQGE1y
iU+2DvLXzpZrMpE+uP2FlcS0idTlMms7eKuf1+JyD2hPbbBDG7cCLupN+a5PJ8G1
Jk1Zjeo/BokRoGIH98dMZuS5Cyh2SExbnlMFhIg6x9WZRKIJsuK47YQ/3vz7xx/y
Gb8pgMo3J4UZ/oIQRFYa+WPwM7kQp9saWmxA+TBcJbvCx9Nyx1jAYn/uN6vyAzdd
LUuqkIGh86xzOj+EmN68QbI0KEX8PLLeOWC/Y024NTA12AQycbBM0S+cAHkQH29t
DNFw/fPBGidKBxbpqQQNwZmNQ6RHfRkRZxTcmwdQ69vg+Wg9SvCTZ1fY9SgWVpq0
IYDMqv3B/ajl2kV9IKQJfus+bjhnPmQ/Ne57UYphnt5m3iGoBFarUkQDw4JDMAK/
NJOMKHqD+gIE4BEvV3NU6/oVs5qLIXGRy4FGQAzBpjFEVhfwhp9USbvFhcozzGq5
wW9VqDGhjseoxsVBpvYS3WpdT6g0PUbBJ+1gR44II9XOZ4MCUIbouV4W97qQtJoo
m0BwLAd47U3Ezgz4x0wPMCfr5L80fS4HGtBDSCZvQrfJEi+m9+Lb/QUOIJoSr4Qs
VxcziZvqmX9zHKpRUyHp0yBrB+ewBg1jxyrVIBbdsl0i3UZzYwQSZVvLJ3JOuaf7
/3It3Nwn5b6SaKGRd7IE1ogX/VNwbpY98hIPuOvW7m6H60BU5q/80zg4occEbMfM
j/0zuXmdoGyC1d8zM8Zh1YZ5uLsDv462BopxtClaTkwr2WTJjaeztDiF2IsL0N0M
w9IXPFyN/G3kl/yf8Nr2qo4RuEU+4Di0409ylfGVuEWRnaEtMb1Ggs5VyHyZevBg
47bv3suGKtcseY7Z2ViRJrZkTpnLJiWaNO1GfIFUBEf8ouvR0fHcxfqYoDZauPv7
Xhi8FRX8fw0RTjlatvWMP5tQoRaoMlkZX66Vtgp6lKcuPX0OgBOlq+Hts04ASamk
gkCEcx05JcFCsGzuUrqmLWaPqW7ueJCX2lEOdM9JuZgoyj4uFh58GsB+XvcTYq85
6KYvB0E0YoiDHuVqWfhhfoIh9jmFE1Q9HXGN9nX2NQ6FTsgw0fEAajvO4ug1rfB2
4L8l3bZpiwGrkSHIL954LOCioNM3CV6ewsJsX+itFOS/CioueRPdIDBJ/Uq86YuU
T2bbnzyoOwMMBL0V37H8A9Zs5srWZ72YKDNRjcf04MUwAeFFzRh0kTBDtXeiAiV3
gx1dVzXEyQI2BC8VeLbbCWghDZy4/BYcUe6Ck0ge1SoWtipHAVulAmY3E+aJG9jq
GoCUwD0rvZEwdsbqPGrfvWobiSQAejNwbC8IVExkHv7URGyYobUbMaqKwdVf+UOR
b2TgbSi7j06dqYBjOHus19cVVS8Ns5ndXxoYds1juueKKEHJDnpka012CBW8TyIV
xzg9QXtLIy6rjodQXP0Si1YExDFxjDOO03iJGThu+O9ut5Qdgh2ZiqvSteZXL/x5
n4dnRYrnWDpqXOiklfs3pZhI4wi3+yrLYhnHMoB8aA2tJqJhYrt9snW/r4V8sfCl
JE3MNZ9d1gC4uJkTpfMPebDWRbhQwgV+R/KHRBqvWEBFCMul0MyfPWRcn19N936h
WzmMsPS6UOtgMwdvQO5GSzAqjPLuAIFTbtSmFdI+3FvNFSlT2cAZ8oCEU7BHyqWZ
70FJ8xUODyVf6uzNekzePrvIoPV64USqfVsHNu5yw+oOC3ju/LXqSfuHpvqa7EKo
6dV91BVZQhrq6u4OnExDSdLpicDr7LmDVAfb2XWhKr+bkSvv+sm40h3b2GJYcL+y
y8Th1jdi+TTeZOoz82Ag0qLGr69Qm9Ig8yyu+/G3Mx51oLnM/AnlhhyOID+3qyZe
rwFa2DeE1TW6ye0hF01MXFSWGdWX2LAFGL7h+Kf1AW3OrdLmb1nz6ExNqAUwgouG
`protect END_PROTECTED
