`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3m7bCefZtFUePjUheC/PtP9g8kucQvTQN2+IlxKmjJHiU5ptkK0Z2QAr6pJR0Yfn
vAzw8phYCHvA4TKuhBj6cki+F0zkqdttFQgK/ANk54vAPyL+UE+RC5Y8Dakrl6x1
0HsUiKeAC8/wDi95jBAFEyCp5nKx7nwPDQBcAVvtO0A5b9mJO/tP0eTexusf+tfZ
C/Pgx/zX+qpL+lOD8MLnFZB03od6uPiDrRe9oy09iHrHjYXXINb319S1D/XpG9CJ
7peLUwF4s/lbhanavRBxnPFWagfN6HvyNTw6DwVDNCCjYy3KGlt+2rRz0gGeu53Q
JhNluv8Cy5b/OfHumOtce5xsBcV+PxLa2JvxwxVlnpRH0Z7eCWN4MFIcIPLX/a+P
LALpt8grCGdpcyZsSamNohxqy17b+lIewPys5Qi01941aJa97b8q9vtp4v3ic5oN
yZpCu56QTg6BahdYC9NQAqLtoCO+BTgtqyK7PR3+7Fl3rCmpegMRmtsC9aSNjnqA
9eoyMvU3SgisCP4caATC/fK704fuccfQEvGTgXFfmnTfNGWQhdZ/pYledqmfnKBT
S4dY3cuY2grDoyepzlGAxkgB7EPkkF76HXjk8bx4hMqeJ5iKbGNkQRucon+Ru9Th
HGUgXwPeOd/+Dsww1whNhXdKdR5teh84z/vVfylAeCQ0zU+LB82ewo8b9bvVV8SH
T/px9QEGPICSOMiim3hJp5z3i2UptXaO/+ur+8qu7cJZkp26gH78xNdgh25MzH9K
t6U65x089NICuPYmH0K0SmmvSDNDry6nb1lGty9sCW3GotANCUODC2fy3xODR7kI
ysOQrg5GL/m0Mv2LzAB+VUrtwGfh93YrVibuD1DYVDs1ODj1tllink3e2qWF79dY
TZedDbCbJkvdZeEU0FPxl9SZTkmkYTXcJVrNlIP4t2BIOUQlSKHZdA5iyplXGH9/
ZwNT3ivq6D17NsniEp0SCwfLkLsvTd+OT0smfp8dS93h/YsPnlJQAAFUFu17vacq
mSuxcyAzgrb0v7GeWktHFFhYnWUOTGISxBkXRTATivD8vjvj8OqcanX18/Uxm7S/
lELTiyiLlSglx8+iGzCLX9Iz6vL3fEf+9CU0LUkhrOkle1q1J++kwt0w+mbRDtUQ
5Bh5ekxR1jWgTgM8oRJ8lU24mTanbKDcJb1yFQHvzN75MZkILv9QYIjoyrNW+z8S
Z0tcahsBskpzgZ1Mn9xSiJC3Ne9McL6ecwxF3nqxJX7A7GI0s0uzjD8Hjh/4760I
dpaazSL/IwwR0/sj53Ik6yHrqczpQj8aJ2LjXeEwpy/QDJT09lYz9AXldZ/ImL+p
wfNlKgg2ZCTna077J5ThvJaKOEjVR/kKUT13CT6apIw/0mhUL4sOJA/dwRJDW++Q
2bgm9DEDfGrIHsZTFs9EW7Ob/BzD1M2ugLQXVDMio2Kcq8tTy9KSr0i057KjgeJn
VA4GvWZ2M5q5uBxxm5wNbhDIMGv8GMScUFzYfE8riBOr+EUpjGa7KYhUoJk9/3OK
XXjCb7IM9s5zxn55+Z7Y/cJuSqfpz8/Vk2PvV2iRdKdJDTAZFxI0XWMxwCMPnwtY
z0W/JueVIM03Jxp4JSIUSAyYoh4wYHKJSTh5WT2cHZeiIjHhErHSY3KlvwdLbwU5
p50Cxbm+H8vg6d4JZlHpsR+N1bZRxpvEpERtyEi+RNHt1YWZ5H9klBYeIV0gHY80
`protect END_PROTECTED
