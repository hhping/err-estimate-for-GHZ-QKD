`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zAAsbZDRTBJXLqkXtpPFDnR0F1737Jye6v2qRz4YDRSdgoAsrENoGOpuVzzvGG66
Hg9wSrAts6Tx26EYotap5RusD9bdJhuSHyrnxFkpOQxnhPd63WAge8XFczJdx2od
qpl6xVLhBqT/2rIR31LRIE3newqSivUa66esWB7pINuQL+mI/52fuZTxVc19ECz6
eiHDjRYd+8HHr/WsR8BFS3kevAkQBP7JhmG9Z4e8DxnkD3rmQm4IEWAaiiQzV46E
bUP/RW0yEtls/h/ahpPnzoh5JhpdAV2W+NtLRmPfRGdJXnwvkRfZRrHSxQ/h4OTL
EmnGd81EWgD8BciN5itBrTjEbDzmTUSqcC62kiU2jpWA9qGPNtoPXXUajnLlUJ0K
isKek7qFWYOeoyzwB4YcYyVQcJr6q66DysJolKjlIkVJOM/M0xKLh7FNTAOMKTSS
eU7wv+gXthDnT70PCatkgJ58Ymo/zQ2nS4NQKOg9If7YwukXBjMkUkxuILkwUZoS
AJE2egXmELf7q01FsXzLQ3IvRq/3wtIPVglBHD2XPozmG1hrIP5SGbaQiQwALjZJ
5OYk34z1xZuO04GkbdF9kAsKahV9ro+JZblXomlXN0wS6a0TVPCvLdAqdCkLmewX
WRoOPOyqfDz6oo9qFwIut2SyFTGDS4Vl5xPgrNPscNG8WmrWGD6ygLMJGQPd4jbS
4xdCbzP9MsJN8H7tCVNEQ4TBfrM9biPOSX9v5faznPIUFAIWEA3/ymOQGV8Nk8N6
M7Z6M5/oGByxcl3yvXVpHwg69OM/uor7OdJ85XBxrXVt+vqCawMbBWgb+vpLJT7T
5sRz3OoUmOTbZd2ZdeqpYYdduLZcDTEhlH2usPZh+7qky/eFMKsfcnakPVhfijS0
n2/uu2chYeustwgKCd6eL6HQW9osjCTGnDo4JYtl+0Uph+qyUcFSwe1p4YJbYkGc
v0Zw0/zimfI3AmF9hWKjLroa5nmc7FsC1gBflm/ubbaTSgOKTUtyAn3riAILzYDx
qHm9OcSWojPGA5ZQPddI1BBVckA4eIsDvMGnplgZbfdx1IOgDiGwy5KDZGPB3+Pf
4/iTlIb1uGmqZ5ISGV1FtzgxEFqPQ8u+1Re0CzsvSbV8Rci5d7nHARiZF7e0W4G6
3Kp8JlSH3fFn4MRHXT3BXphPoeehw+1nYoArdhPVbQfw1/eGKXpiSXkZJSpl8TmF
hvOmXTxx+GGIwDxd40XWkhdhrN1SzWT7rZ9+39+kfxZHfcriLFKXmdzx3kqgtbAx
VmJ5CA95VA+QV7t8rhjJm1dqC5LZaYMSMs/gtUtaG0r8mfY7fYoCJeXqDDECx8qA
LkoYROoidE+SIAR/wJhHVKgQtC+cYfVN4EAp/QW1oKGfAnk0B86d8bmzYq6tZccz
jP33/x93f94vGXfNWcmeaFVplfMesLmHE72A6RMjqcB4blzwcWoPlMpOSmKBjE22
kLmgqggh3aC+tydN/89p6AsUb7JhTU8j8MDETmhCkGBjD3hqcTUB2he3NxGCza45
bnb8E9GXgpaekq6LojCYyXje0QPqvSrQDTWtaIONGkUPf3pINgEh/pXqZnqPRqE9
+YrBbxpbf/W+gyy7LrKIQ3+1MCmF7OLZvB865ix/74NSXGwzrle6ZXDfutPANgbM
adGFr1SomkftVnCZxENLbcviAwbIumav9FQLLiKCmP7PwqnqdqtpzHttVd2qRSob
dppwVfpefLCXI7ls5/hSgY/myXVPsTgRrFhlmXopzUU21cFm0VoBXsqHY0SIrxyZ
leimLVFy599zZEnhixTm55XTyx2Q33z0WUca+8WhQpWOu6RAZy2KVD9t3aA2/Fiw
lVb6W0e+VKjWAXVp6v+wbnthL/Jpt/hN1JDaraHkfCwpoVOtBjq91sGpCxYCX6f9
avcHQczoQyf5ngy9IamE28NuvrVNw0LDtpEcQ3l/XknEgj++H7vnIAMMBMZS+eMN
oAnX/gtSSOVkMrtb7HuUpQ==
`protect END_PROTECTED
