`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GieazlxEcvISp4JqabaJiff7oOp7CoM0xR/shAGUaa6Bl1Zoe4qJ7w4l5ujpS/Mn
YpzPv8RB64rbNgpmhfQWaxaw46AOnLUxxev6NrE0ckrL332PSXY17vW1dtZxfevw
it3JDOyvESciQ4xo54+jaFEpjQ4N/mDHT14xMvz75WzVUW6teS0Etj2Jt7uA6ixa
bCYpt1QXNGNHz2dyhmnIkzfOT4PX/e4ajR7T+Mo2SV8lXVagcQf4q1Y5xFRVzzpN
qS1pHfqFbkYfYl5jCWEgU5bnbPB1dBEJAgUZQDs5Jspygz+8NojKf+qp6//DRLzE
tFRaNC1WNZiOP2fexpfPKp6QWy9R5eqvQKhBX6Xojf+Cj9f2MlFB37YT24X5J20n
yZl+sGWcSZMi3qe6AlmVidE40m9sl3JMSDLvaGOSFsF9ANt4AdsHvkv/2Qnx5hV+
y87JbIfrhLp0G9/vwZK6qiZ+nvxxN1oDzhAnJAzPxTwsupIayhaDoTccjSZN7DvK
nCckY9ImBAgS7D9jnEFDZALdJCcT5KZI7lYqAfqnn/WxLGLB/LCnXdegu+sTmk0O
mYiGNzlCsPtkgwbIpi8QSqmKrF+HxqmmyQle9TKJTIyvgDxfMg9wghqZ8jLvxEMm
zsDTGi3lHk9Njn+QL+K8xfjT2TrU640zXMNOr4LFhxuiofqort+VnxRmYeQcgUYN
L5+jXnaK50uzbLYv7cgmzYk5wq2VgUtkPpVV4y8Mu+J9RtpKdl1/HJhRZ1XWc3H8
WG1SdmYCqNbqkRMSXfUaErXesd4JyuDqpIXesXzJsq3wDxz9Obb+PMsdm1Bla7RS
ZxUb1/FMjS/+KVmYxhpVgK1h6dexc6ZxCJsZUz0C5NwoNpBymbW8qzSmqOBvNmx9
eoaYVsG26ToebKpOtK3+5hG50Dn5n1ob+4o0VQAxjj9Lgks6RkH75s3iXK+1SjuE
li7S0OaBZBRf8Tbk0hUu95uU0w03/NEBXM6AU5C6nN0RfopzgoeHpV5t8Sq/LN5s
pbBLBmhnG7Nromoh4m3rezpRJ2wHFZ0wUqVAvbWRfmfzzTbaoKQUrngbCGehgt+6
1oGbYGEq3o3dbrROW2GDXOKQXQeeg0MQUaehSGdfRRS+h9U0fFnkTXtNj4Pt6DGX
2S7eD4LhPUK5VMpbTm99haJ8aJ6zr82VKXDhRmD8TQwhXlxyj/bc5aKsdH0DGe1l
Xd7PHJgLCDMoTRcExk1oS5YZSqyBgxmzFXGI46l5DxnL0kb7eberIZqNScDnz9T4
2/dBONbZc2A0mPI7Yo4dINhQEoS1L+Fbyksgb5JVLLYhvudO2kOdofxhAjHiPTI6
YmIyWntU+X4S3gW1jIVkchydl7Yzgo01EdZHypfTw7bg5tzkGx9vlJDEOqbfVmbT
eLmEV84rUKylrSkr5Nk5K9RCxnPm2O05pBStQtfUNesEJQqhJuQBwkj+wLjUK6eU
QML+0qnv/YgcZEzF2YuuWBv4yBghtdy6vscxR4XOPMR72ZWsQvjvcUMfB6l5Xvw7
YCH/zBz8ZuoSADtjMUraqM6IvedXrmp4jvOjwDr4r0uIRvoBBpqV4A+siPYvHnoO
W5/lG+Lsb6mHfMd2ADgzLURwMDXG2Ja6ZaxJEV/hgfe4ta3e5W+pBOFCpxM0vFJL
Qz60XEcTiY6FAqQ1wkYHi8O7NRumsa06y/cPSQvP68+l4irh2g3F0a3wIqPzaLoI
S7nfcWpDBoBM/fzlLfC6xne4Zd9w1oJOdpG1N38sfMS/AYR8GwS5zo8zfNq68MAj
Pa89YgIbT2nvngDXHdoT4VZlFwPJlY5AmAPD/0ZmieMLpdq9piAGgPt7S2nmU7kF
pMbllW/iA15rjvr5eN4h5dyz5NOXiEaI06vqitgp5qBRaKTARV+Evj+rBpMcg30N
Rq052ZKHaDntNIvB/4t3b648DRNKUmrVOuWIWf03EMaM+ebla0H1OZsQ+p68A9p5
a49jBm0T08uawvwRajCmXSA9ZM3xBkgP4uDmuI++2Yfjho0vevwcqOn/xpL/7AoF
mlbPdqYJ3GLpNnh2xUWj74nricEojGyMv4ex4iqt3cMFto9Z49ZgNpQxYgXx+3lN
fZD65DQ08cjvx7kgBjS1fbAdl1D2dgb0/xrAZltPgHHp3/PZS1d5a+le7x36dt7s
gKFFt9uUHJjPkc9/W5VezVb930N3tp+op/EBKz/tdvlCayTCESmB22q5EV18WTap
ROD8kGxTl9RNmqwVsv9ivt15JsceoUqipMybWE5IV/mTNDAAoBgc3ZrR8TewSF5F
kb7b10/vBNWABx80aex9dmqLDrbzi2JxgYYKQjIhAP13pf2RUT7/84pmuRW/2VnS
Gmj1I0lcU/SbkBNVKPTOIgNRi36/1aCjcv45RaBeSZScBXvKO0WTGR0GYKEjF//b
6UPVuy1cnr6M8wj6wdE0xdCUPtzv5mnza+SBvnLDYfezgfktiVMT0Gwgu4EOdDmw
Dy7K08+AyWmsudTo4e67TVf8jbXKxCCnvPPqx9xOnKmozXebXaQ8U9Xdwbsu4VbH
/dhz8f2EsvyHlIpwsb2icQ==
`protect END_PROTECTED
