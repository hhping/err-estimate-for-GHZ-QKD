`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
irgwndKjoSPFN8Ltp5WkyxuV8jrUmpi7ETXb+fkpVcDfPkjsCg7B9McaF22Pwi7x
Ex1QWnqn8Fhl5InhJGcJIp3NtcVLcsK8qP8nTvtlB8GwLY6lTahRfQLfgy0Oo0db
YNqX/ZDGDT2fBsksH5GMnxVxIcq2xMjcDdKteSuhnjUNM8CviO2XM82sRLibZyM7
t2ifJznLGeulFbMth3OTCbPNExennn73PCdPdFSrzIg5N1w7DLYBEbkgLxi45GOU
F0IjqV4dsiAD6Ok7o/HiLFX7A1+S1FoDba2GheL2chY5i2NFAC1AKDxAYXh/0YFQ
Gcy5SmIl6VzIqrmuf23A69qOyCGam7/qlshIzBKMwL9UQZFHc1p3hvsZxY6JzsKU
rFT1g/Wvri39nC1T5v7CmS4quiatMcyJl4eaaukZE/ouZZQaQcGNDmHIEUNeiWQx
oZw+OPWAOb/TbGW2RXi3njU7NbynBUVvRVICzz+vYivrJoiZNVglN1K5TNoPGdvH
W2WfV1UzzzotdjFsMq5Ybtdx3ZWRvASVtwY3iuoE3FhjTaKwSVVF/vPl7ELkF4v8
w3FPohOz5mqipEE4NECayj/kt1S3b0DLLM9i7s1AgaXF9T406RjMejPN5qpYQ4me
/sfX5gdhKn9vJQBTd8hJ/FA0X2KU8yBrPeJV8yXNaURvboPKwDqZxqkqUk/ta6mL
v02Ziaoqf+jqeztpHlzkZ9nHyPj+cAOKr6v/vgyaKZAUbj5jWLcGDRsAETwkgN+j
yrLjrfsNyK9yoRj4x3pYBD/bdQTebCl1FTNA46pUtpjCzfhGUT4U0wx6Y6q+yR6k
4On2vhCnTjsH224yfhahUbJgfnlIixDljbTY3sbMVTlFc8RFn2gLR/3rEfevErur
YD2kfiqv/Urr8e0BJdEJm/GhWWJw0/kF/AVYOjf/kBUSDYkVKXbAQ7YPXYzunfhE
loJXC4Tff7J5MZXNo0qneAUTT8+c2TCQCt17cahAMRv35DbM3844tr/w7ULqkjNJ
YeoWSKdHmAxWie3J+M/WcdoChsKoFOsMb0ffw1kdJjrGUQi1nowB6Ipl2KX5U55v
e1MPALptw2JL6ZKN40+foY0GhW+r2mS4PGYAie5bmoaFUEGk+OX9dkdrgpSCYtb+
YEFV3P5OHEdmubjQP7eIbJIKWv+RSa28DbNlID6ZT2rl4JElE9QW52Trb3nD9Iaf
5dtbuQFUoKAZtHtvySH4SGsGNWhHlBdeoAY1IfRucsssoQu/WUo5ZM+imFxSMj3Q
0Cei4R9UjkkR6EFX8IFUIysiLBlpRAe4wugHPAnEevuCsnmI4ZzsoRdwL2Q/+j1w
CWOGtTcTSOmnS34VMeIYPVhTnYTOKdPrU/v2AqFEqUOQIAC1wzbJugqbIbEkBFmK
NHcqaXYIjiROwDqHSotxDAfakkuIskTIHtK6iGGOg5/r91/xafzr8dBlw5P0++gV
GA4iP28WnN0BXEkudCbA26IPpJ1dyTg1FtWWRC31HPUUSE6jsa+oeePN4zQXlCxd
8CkSPt2NsflpeXiLJ7n7RMqKWg2y3kUFWCJYDFDqdBR7k3PUD0g4BoVxFi1C3qTr
SLbofuNk1qfyR2gVsLK+dvi9aIRqe082eRaN9z/hj64H7aiMgHStGI/Xw7MtBCT6
zXxFNrHw2iCJlDYWQtCM8pVOijdIbEpVmCVkXgr/P3JsbWhz9EiMZSQcfOUGGCNt
B4lhmicWkJRqBDpVo4WdM4WqwqIvW5Z2+XTMSu3X6T+NkUIjqhXnFlB8ZdQAeXqu
HFrg0ai33Q1lWM0lY2wdltlnG8dsBygOUeeJlRU3lOC+w6SnNyYwz4MCpZYeiFtb
Cd9Bff8e89pYn3MCKp1b+8IXxO/mYoIV/kQddHI98oCFSFhVM06NUgjJrtjLs/bh
wYLran8UMKZgzNipfIxepUocMJNKp023slf3IQoUTSrzmzfFdW1BqpXcrGP84WUR
xjTKw2sr99Z+wkaRulBFb0sYx9S6j03Vd+F3vUE1r6QluQuytTqKGeMMsc5e8Zxn
XqHcaCGImCITxb8xEIJFEvChLP8dw6NXYCUhy6UoIW7UeeTPT87bKuKVs0SxO1Ft
Ca/E/4LHe1RLQTBftCiOlw==
`protect END_PROTECTED
