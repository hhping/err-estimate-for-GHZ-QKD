`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QOD+oRK/DsCAc3E01vRIMSzBc+q712dBYxI1yTttW/nneh8uTRuZsp8ATQh18+2d
AIn7xj9VnDc2aTER7Jj2bCC12hyjeOo/j6OBRpr6rPYf9azfj6nHq2Jsc7r+HexX
Dq2CudcQiqIg+OGmT2AYVkqUdSqJQ4u+sO3LicdLM/r2SFLWcmXTb7vqhWXd4o5W
3Qt1515uphu0B0RrzRn9/e3Vh1SQpj+Ow9YO0mfNbnjVDXK55ukB96Z+tJOc/AE+
g55gETlR8v0hSGK5Ok0lF61EJUWyt/q7YJBwuDp7nESaLvZL7hotVkDo3JZ6loP2
DVI6lIiuLcZGcmd5upyPny9mdhivewF7fmW83C+sDXAIi3+4G/wxFGZxHqDNxanx
9+HfvWc8lTwcSYv/DKqHddmhDPZSmZww6JmITso3lV3c7/252/oRtAMcpaVKyIdw
zkqn1zI392KkACmAoirsD1HEOc6uKu2mIJG4ZBlDFvk=
`protect END_PROTECTED
