`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
99wDInNjFxZn7bqcO8DJWXeG9s57bF0x2w+dABMEAKEbwCbaF+4ag+auvEa9KKzs
IvkkCXE1J5Kn/RTlusnA7jGp4O4Dh+Kqp0STYHQAJ37cV2ammA5r8jSSoF7FGLIq
7XoOL05d/HBoMD3pyG2DaNF+til5YAPfCXNQIGE1ZgAOp9UOqqJ0GuEzpntMsnxX
kB5NeILsm/AHAQPwDl0vr9TirB9zeguwlJyksF8CFt7NJJ/NwdlYE0d8wLTqHT2q
je/l7vq90eecvXy16hkVW98ebtxuoft8oFDt3cN5gygpzcC1Jx70Y7szowd4ZpgW
cSDtMcpAfWxdcB6q2u1np+1W61EmYCLsjy+3HLxGXe1EmIbXTrQ/LAx0AQs4gJOQ
qcGc/sEoP4YLXuhoggxFPDJHvJpTyj9PC70IfUhVPqyUJ23lhYV/cy4VIIJh0CJB
iABePtU1Yb8cleyRICQ7+J1fmRcFybawMrY1tCPxeF2IkUS95Da3E1fSwqGjB0Mb
ATvTPFCryXrJNFYWZ2BDNZanp03kbcReYJmQJDxxy9I=
`protect END_PROTECTED
