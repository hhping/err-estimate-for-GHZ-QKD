`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oFav/Qm91jQPNxbVruk1euy6/W3JdYx1Yg/Q+B3zCHaCb3LipwNUAR/wpjaFxMSf
WvPMW1XKcbVgtC0dsI+i7JG7C3rqR5hUs7h1LlS9GPErKlZIDlWi2cliNN5nr0Ff
uG8af06I6f/DLYz5CYjk11JRgUitHfaT23vcvZdJge8NKUQFlk8YQjQeVvkalMwU
UNsBiLQbU0oekyv5Xaa73a1GiuB6DSh4VO+p3DvTyyqjM//rD/I8wkwDW24h/jVk
wlDeE5LihqpJvVP0UpG7s03KJTofu81zYXpyxP0T5Vx7+IPLFHnlbNalluEMa60C
JEU79kwjxKOK8njpBIlBFQ836FfosqoNvxX/jyqjV4WakRFKk3CMkRiXqKdFtsEj
Nmas3r8Y93ym+76Okc7ysnDHeeWaxubCGdbSpxt+wn2vhTZf/+tzQKfGFQDzB+9/
aUULDLHyZbdbMfUkReImiLWHcsqrC2wfjkukVSl8RS0/PDGm7zuZmgthFL1BxqxC
KMMIoqeJfZUkhLdP9O4JuNcbTdjUudf3z7W8ioqYxnCRrOjt/Q6b4ZYiVhs15/ES
HPO8hyqqAw6M3ExJRvG5fZGSNxpR2RSIRAx4nyZGYphLcyP091h6ojRCVp3HH2WL
qL2IORUdCooPYFjmF0FNeROpFOHbSWPyszhrfWGp5kE1Tc5jVoZnGfSA/aRNjbiw
m4wb3vduU5IDoi6ouLNeuactQXPP317WKsmGhRaEha+UlZPwXcTmQexum6Hr09+C
ckqrfmL4dFMxXqwB2gm3JpxgHknVqohq70/xpPUs0oHmkB3dQ3Ovrvs3jQMI76mk
j6neRwTYizVid9sywgerAxAsCDUbDKDi1yXl0sVyWI0SfV0N8MhdBPHqAQ1kHyW2
q4sECZ9ZUcqOSbzdOIGJ/RlbxnuntxQQSDHmTsfT8FuMVvtyjJogfSciTH5qsmm5
hFkIAn1p4Rp876Q3ikP2VEmQWY0bmxYqMhnRCwnJvdnmX0PcIWhwjJaTDLwe1rWc
Vod7iRAzTnQ/VvXFQTMGSz9gfPv6rTaGSXRtyC0nSLx6KLGpZZnow4gg11sgzlNJ
+Jhj293Yq5+3JCoBa8ZZCYCHbXwMwTCI5HsEKjT5baPzOjKuzOUU1gaaC42FVrqb
LUORvrZdCn7PeXLK4LF/G+rz/SgcGFLE/nzTfSTo2Z+fFJtrGsPwr5cLEwBeJ5Oe
pEkj5XBpmQpAa5fy07J+SQ==
`protect END_PROTECTED
