`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KruFjDj3qhT0VaZDLGTDD/K9CPLuxHDGge7mtFg0SqlUFV1b9PNMU1ZQvkXAyqFs
zIrTmzxRE6iN7+quex+DjHJl4HtX04R5cuzQ27fWNT1k47JLVmLFK5j53kd7gXDB
5M66y+nidd/FWA3LXtX8gIb1Bann6I4yXT50z5h6fh3dNkqWxOPl0MLRiw1yAQbD
YQLbTFsUPUOO79bHC97TDuVNECUFjZfW14of8zenv/EQQdCxFgh+QSzURAn2Npir
P01lEoedNW3fCug2S3p4eh15Byc5Sz7k+/6aBLUSEUGUbhoY2tesdSBPX+xZh55Z
ZYhntPlkfXmjjiafJXYTbyi8CQfVgnugw63PIWH5SXcHbofH8Cv6+SP7F6y8reH7
9vaDIzAoFFwefeJR+0bHdXW9nNPxBpAjltx3eSsvpb/tfsl7BL/brB45iPIYnu2P
J+NxPhslYTQUNXAgihX8M95CJb9iryHYHbg7CR1ORm5JH9bnhuL7OEXfzTaHYGqo
HmRpXVJlRHGkKpl6VUvSk0qs5CJBE8lS4UAANfwzLlhLV9AdKQobjQdy529Gz1nw
tq1bPpvoTKJk4iQYtlN+JmgY6A60edd8HPMzgE4K8WbNyLBU+OSw7Mzo+OBC6NhN
g/e5b3jvHBXdxWiuY8K0AxdupYojDeULZ4vE4qPgqLB70rznc67ZXlm49fz9XDPC
Afk1UjBi5iOe2UH6rWd4+E11KbvdyEsYR5fXkr4BxNz7FzIzP2Q4q/ZeI1a8BfU8
cjbqLJnJvNYoVdn6/CFc8k7kbmgaks2PNVViw4cWnTpGf/qybj1K7786l95rzFIC
Gtd/FZX1cOb+laSnHf2WIy+8pOrck5x49ZUzpICGdXzulUjy+Y4Z51mtxgAY8NR1
2xLjEsdhuukGn6DHpB5CFXrPAYPsE55v3Na/atvG0D9VrxJy8Nt1PqbJzdiaoWAI
EdWnkKO9Jx4zPE3GBmfwdOTfq31rc4hDWh3kSzCVtYVibdMAjyJKwgc5aAYDaAsp
iGpIY20H4RaaFA/rZlEsGsxX7C1fKrjV8c/vWsObjXgpKxfws7mwq3OUrqE4S95A
WPX7/UH/5qKUb+vJL0XNbS010DkqAN1LxcNGCTD4OrCYvGMrAjye4yF6epfTQaPs
dcnxwuAxfFGeg3DdXQOZM53kBN3xZHLSA1D83D7QdGyrdRrgKJEitPhgPzbsHC92
yL7hQ6SG4QY+2o2EmMFvlAfj44dcVGPfA+owsJewCaYFco+eReqtQ/NE3N3j9Evc
uHDw3oEYHyLKIJaaTlNuC/NvlGV1mSP4vj8zCaV3wgGugNOGrROXRQJHvYF0KaRt
Dabq9hW3R+NPFQ/5vAIyqcNxYtzziu8MR5OZhPt5xusFJ1D9pOmIfrZmg+sVIAS6
asW2DWe+8UYR/bCY48rkOdDprt7Uc7+DxIesq/0ydLIDl6xMNogp+zg573XdfSwW
TvUOr74d6A9DzSBb8KJpr4S3XTICxEJhNn8y0tLqAx+uavy1BrGwYHhoikuaLQk3
ff/z6zwBZm0DqXwVy7SyCBUt1St4CMrbXUjfbZztU6MHQyBzUBCXhpVsLqBWb0bL
t70GqUGfGtO8LeTnvUrmXq/AmWK1SHlHtxcwZthJsZJzMmUR6q60UZ6w+O7yK3lY
Rhi18YyfNrISrew7pHDzvR92ubTN4x53lq+oNZbAmZYTISKFvzArjTEDXuF5goeJ
ryrhu9KTxuO2BFoe7hcVyGXp+7Aj/1YoSmoMx3va2DM0b6fZpvKiE0pZd+r5J+d0
QRwre/ZnnUGnGJHjroQ3mk+/pBvc9yZAoSYxAMu9K5vH0Nd5Wu/ogIUntasJBsfP
sKfdJ6NfoXwMjvwpireTWCRZpMI25fbZfCJc5aXNZZVnuvseaVrXEZ2iQEUu65lU
mLJwO7KcmcGbYfLTYr5SolCc6dGV4lSM4Dd0U3Jx3vvOMcUkIfy9QztV2GuC5BSa
/Kkv09oEYVyneo+cg25NGfjgXTx4HK5Ben7COF1GFtO1SWv6h2+8b0DdVhqqWshY
NZUyEFY/GG1QZoWljPkxYr26FxogBmw4iLr7s+vrxFN5nh1QlIsCzPMoH/brBM/Y
65FnXAcH6YLkqH8G24CExblhZMhA1RTH8iSdzrDbsWs=
`protect END_PROTECTED
