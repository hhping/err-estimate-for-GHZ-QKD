`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QoNqmnBKkh3OlR/x679sPMJC0JyEs/G3rIbLxNaEU8u04YCkyV/ujFndcjkJXkVU
SVTelrQf8QWEOirlGy6aImAsT6ww4Dy1XQlBIK2pJMWnD/OQP8OSooZsCK6LvhOd
6TvnfHPA2daiwM+R9CECDKtMLvzZgegVmf97SypEfDmlavLMPcRMkJ/sUekRT1X1
qC5Uz4VPedKU5JtKIITaU4ssPNdiGXgDhkHX4ZimNAq0IrAKneG1Ds3qqcftneNV
Boq0uPiWZvaDK6zvFozy6eVbf3p4CrUm+/rL6QL6oA99dikpzLvJmZ89FjKU8Qtj
GntxJHd6prxDixFavux/EskyzsH6dOi+N34VT+VdliqqcKH5tNRsXd6SC97/PfeS
Ozd2y6M/Ji8fe7/YbqaUzjNn3hud1jcd8kkm4f8c+zOVE2ZAtGZmtwij/jkkvJ+E
X8Rr8qIjXOUlD3lKTHul3O0d15u9SQhf9k/l2uGrlE1WnFHp0l6/PkAFipFGl6Yr
4+2h7Duf+7t4LWAAQjj52vBC8flb7jCIgoZjlHctHraUhoNhaqRC5kMVImFOWUs7
twy57OEr5IFlwuFR3TiTNyc40hlkAdoM3ejB1qrNYBQ=
`protect END_PROTECTED
