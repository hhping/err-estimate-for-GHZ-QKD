`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W51lrcCfm0dyAOMXoj7m5GVuMRLDm2pM/IcSw0YwDFaO1xqo4wxtfgSoF07M9pvz
V7XGKYM9XrJ9lEAp1USnnsW43E9+v9eYO01prXcFiZsFiWxS5mVIKcwt1fV93Fhp
p6qAUhDW7k2WU/R+Ix/zCC3OgD8DY+NKZxW2MgyrIf6A4N69JfQEjeScn18RYuSb
iEZeGoZNVeEOuwm8/6W7KGEeLkcwVjM93VHPlF06bq9Fl7P6Z4MrdhKcq8Lv+t4a
taQeGD5q34os7GIbeaXqMMdlojfgkuJppK/kNQRn3hB8ROhqZWVs1Nz73eRe7qGJ
JW1OOK5JlnInsyOlMgaAFAeDXZJ5S8QvTCkhp2omP9VfXER8KS1U8zqJWYIj/uxL
hTqDxpRRv/DJB1IFRgLlF8jUUviPpMuoEUVs0KT/ojm/kvK3BiXCJSdeUQDal1Jl
ZTkAZVwZdiLUerLQdzkfcJFuFdL4iMJ89sBoVVNGUMsOi9ZdlInYeDUXuT7pLmqg
UGr2N1CT9C4oN7ickE6uSWkUhT4XOst5vSC8oIaZPOihJ5Y4XSjPNbiMeqivk05j
UA+pGN3xTEJQKZOxTNgBWzsULEOPOmTiZ6SQ1nr5ejl5RRc9sDWZyOptoxMO5gh1
+TWdmZkqZUFSizSwTbQI0+uQ3KljiVdxE6F8Y8QP5DGUGqpWEMZ/4xePka+/MLgO
uIkBNKurRc66+w6w1TGHkfbAQuyWFMIeJy2h7bPa98KUcReTKxQFth1lq6tKa+9R
qXOntQZ00IApJLHKTA/YnDNq8DeEBiKGejSTe3+vA4elvaj6ELRGV3+xU9J7EPG0
KB+WGoKRwAZd9W7H3i5EFTtmYR+mUycG0Icrw0vg8wmlm2ZczP/i13GSTgImfPIg
zIfKZK1xTfgWFI7aV33W1PM37J0W8/pNsuetmeXqiJTGbmfkcRihNe5iX9qY+3Fd
shHvQPGdeWQvTVprDd9R19k5YcGV2YQeF8/tqj5Z/W72cWF/+xpGGhtSd4hG/0hR
IWCo2fq9XsegCJO1sOtVHXJQqnpJ5uOw9ILkAmPrWm+k0xzmVCr7CPLdkWXHDTuh
U/uDPf8Bf2oTMe0aKjFdBg+Bsh4TsEGLh8wx7RNKJDF415rrXqMWCw3hAyTZd0J3
oiIGHzIyU4Yf4TtWEWvR4642awDtgYLjmrREDwy44Rvr+bJyIThLxi8nPLd2n72F
R1RDbTJVpkR85YNtOgpWYaOeOP4qoKLgB8motntiEmUZ6lfprvlLrpL2VRRnHmvb
6NVYzU2NLKucpszOlL0sNQ==
`protect END_PROTECTED
