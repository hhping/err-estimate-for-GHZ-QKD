library verilog;
use verilog.vl_types.all;
entity twentynm_hssi_krfec_rx_pcs is
    generic(
        enable_debug_info: string  := "true";
        blksync_cor_en  : string  := "detect";
        bypass_gb       : string  := "bypass_dis";
        clr_ctrl        : string  := "both_enabled";
        ctrl_bit_reverse: string  := "ctrl_bit_reverse_dis";
        data_bit_reverse: string  := "data_bit_reverse_dis";
        dv_start        : string  := "with_blklock";
        err_mark_type   : string  := "err_mark_10g";
        error_marking_en: string  := "err_mark_dis";
        low_latency_en  : string  := "disable";
        lpbk_mode       : string  := "lpbk_dis";
        parity_invalid_enum: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        parity_valid_num: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        pipeln_blksync  : string  := "enable";
        pipeln_descrm   : string  := "enable";
        pipeln_errcorrect: string  := "enable";
        pipeln_errtrap_ind: string  := "enable";
        pipeln_errtrap_lfsr: string  := "enable";
        pipeln_errtrap_loc: string  := "enable";
        pipeln_errtrap_pat: string  := "enable";
        pipeln_gearbox  : string  := "enable";
        pipeln_syndrm   : string  := "enable";
        pipeln_trans_dec: string  := "enable";
        prot_mode       : string  := "disable_mode";
        receive_order   : string  := "receive_lsb";
        reconfig_settings: string  := "{}";
        rx_testbus_sel  : string  := "overall";
        signal_ok_en    : string  := "sig_ok_dis";
        silicon_rev     : string  := "20nm5es";
        sup_mode        : string  := "user_mode"
    );
    port(
        avmmaddress     : in     vl_logic_vector(8 downto 0);
        avmmclk         : in     vl_logic;
        avmmread        : in     vl_logic;
        avmmrstn        : in     vl_logic;
        avmmwrite       : in     vl_logic;
        avmmwritedata   : in     vl_logic_vector(7 downto 0);
        rx_clr_counters : in     vl_logic;
        rx_data_in      : in     vl_logic_vector(63 downto 0);
        rx_krfec_clk    : in     vl_logic;
        rx_master_clk   : in     vl_logic;
        rx_master_clk_rst_n: in     vl_logic;
        rx_signal_ok_in : in     vl_logic;
        scan_mode_n     : in     vl_logic;
        scan_rst_n      : in     vl_logic;
        avmmreaddata    : out    vl_logic_vector(7 downto 0);
        blockselect     : out    vl_logic;
        pld_10g_krfec_rx_blk_lock_krfec_reg: out    vl_logic;
        pld_10g_krfec_rx_blk_lock_krfec_txclk_reg: out    vl_logic;
        pld_10g_krfec_rx_diag_data_status_krfec_reg: out    vl_logic;
        pld_10g_krfec_rx_diag_data_status_krfec_txclk_reg: out    vl_logic;
        pld_10g_krfec_rx_frame_krfec_reg: out    vl_logic;
        pld_10g_krfec_rx_frame_krfec_txclk_reg: out    vl_logic;
        rx_block_lock   : out    vl_logic;
        rx_control_out  : out    vl_logic_vector(9 downto 0);
        rx_data_out     : out    vl_logic_vector(63 downto 0);
        rx_data_status  : out    vl_logic_vector(1 downto 0);
        rx_data_valid_out: out    vl_logic;
        rx_frame        : out    vl_logic;
        rx_signal_ok_out: out    vl_logic;
        rx_test_data    : out    vl_logic_vector(19 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of enable_debug_info : constant is 1;
    attribute mti_svvh_generic_type of blksync_cor_en : constant is 1;
    attribute mti_svvh_generic_type of bypass_gb : constant is 1;
    attribute mti_svvh_generic_type of clr_ctrl : constant is 1;
    attribute mti_svvh_generic_type of ctrl_bit_reverse : constant is 1;
    attribute mti_svvh_generic_type of data_bit_reverse : constant is 1;
    attribute mti_svvh_generic_type of dv_start : constant is 1;
    attribute mti_svvh_generic_type of err_mark_type : constant is 1;
    attribute mti_svvh_generic_type of error_marking_en : constant is 1;
    attribute mti_svvh_generic_type of low_latency_en : constant is 1;
    attribute mti_svvh_generic_type of lpbk_mode : constant is 1;
    attribute mti_svvh_generic_type of parity_invalid_enum : constant is 1;
    attribute mti_svvh_generic_type of parity_valid_num : constant is 1;
    attribute mti_svvh_generic_type of pipeln_blksync : constant is 1;
    attribute mti_svvh_generic_type of pipeln_descrm : constant is 1;
    attribute mti_svvh_generic_type of pipeln_errcorrect : constant is 1;
    attribute mti_svvh_generic_type of pipeln_errtrap_ind : constant is 1;
    attribute mti_svvh_generic_type of pipeln_errtrap_lfsr : constant is 1;
    attribute mti_svvh_generic_type of pipeln_errtrap_loc : constant is 1;
    attribute mti_svvh_generic_type of pipeln_errtrap_pat : constant is 1;
    attribute mti_svvh_generic_type of pipeln_gearbox : constant is 1;
    attribute mti_svvh_generic_type of pipeln_syndrm : constant is 1;
    attribute mti_svvh_generic_type of pipeln_trans_dec : constant is 1;
    attribute mti_svvh_generic_type of prot_mode : constant is 1;
    attribute mti_svvh_generic_type of receive_order : constant is 1;
    attribute mti_svvh_generic_type of reconfig_settings : constant is 1;
    attribute mti_svvh_generic_type of rx_testbus_sel : constant is 1;
    attribute mti_svvh_generic_type of signal_ok_en : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
    attribute mti_svvh_generic_type of sup_mode : constant is 1;
end twentynm_hssi_krfec_rx_pcs;
