`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w74igFKzNYL0LwVBgpmZBWintP1RG2Yc717ZstdggaRpKN+KNiL5U32If8zZ1Yga
DokW0LCnvrXZFWvyyuWOVTWG3I9JTvnwNhK1HEmucyBnmQSCs9fjDJN43lDimTDM
PaXa4NqytQ7zp/j8NCMtlN/lhezBBCAi3bPsQEu1P7CB1zxCqBG7HnO6hBVdrLh/
O+11VOhzG/6yrjCMcRwVxLe10popb83R88QbmQzWHbvMBCOYbwbPFVd0dRyDlol5
vFI/KNrWG+LX4AA1xa7IYESPLlZlUMXHU1fnApdTtPR4Dd44P/r/Da/pxXpjwH+r
MzKKMqpu/nCkturDZyzBJRWq4nuvGdmHK3Fp6D8aCHDpFKKjhT0hH25qKbbQ60K9
DTI1HucmiAtsnq5IXo8xrUWmBLujwbU1Y8A0qoJRhu2vy+GLtII9HdX6H2YFplbZ
b8WOmb283KaKKE0OkUlHPyq1UQ9LxrlKC30HiToLlkpMpFrp7xlPBrP/YvJbq+su
jNO3hiLTwHk/fIm+75SV9h72BB1ZZqBpHNQVGf/03EjM2Ud16KgOapvgY7kNFyg1
+4MBRoQ7Z+RzRwAKJI+p/3BP91kPML5aXjH1Ji07Ijo=
`protect END_PROTECTED
