`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iMIkfEPQ9Sis96edNfusvn0XKjBa9D0Kdh49iDEjyWb3z92oRLVR6dTLYvS4Ra3D
USaY72ZObWJCUeBImvSGmUMT+iB4VCCvitLTOsenivnSG7MoGefY0Znih5Q9Q6K9
NEjsQXLkqrkq0maeGl98uhQtRurbmF+A0DItXoFxwbrcN5X6JQpCi1L6t+mmmQ8+
Y3x3m/4IDv5FNE1T7CmiCQVa2Slrgtdr/A2YN0bbuVOUo/DMNAAxMKC3kXtR8HXO
n1/c1f/e5J+4GV+yg17xWBkLopaxaGyznr3oTUXrgz7tbr1Oo1TQ/TvFNYX18JIO
NyjAMVAl+bfKT3UksfrMEkXCkvjrCkaNaVOXrIo80E5I3miHwZ/TJyg9xEaXRQHe
gWKlrweb+Vy9Ty3iCSMm3qoau5ZgPF7Sw7iJK2vpXnQTk97KYHNtuPXE2jueSQbO
09H5U1GmUvEkYLK12v2l274/FaGEunyrzl9rsHkUH79TBM7RdFPGj1hhEslxwTBl
0T8ucKq4DOHx9PI30TkTRw==
`protect END_PROTECTED
