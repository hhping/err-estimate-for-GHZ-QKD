`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WNuoHfb03OBrHl1wYjrU2XbQuXXjpjiM/J9GN41/OfNfjYmpIU6hrCqEHMWl6/kj
+ryRsQ5q3AVs37pr7QrHn036yvsUQUW1BMpFnATXfJcbtF+EPs8o+4AJ4Y1hhnbD
5sKbTg4BQFcMFrVgDi7kCTO+sXCZnY3xmkOyuM09HuF8Cqlvb4EgSC8Z8RCIVcRF
k2TcJUP/Yg95XpJgaVWQ+KEpLeU3mHf2iRFL5lNqH7HXSEMCGVVgUSaGmp98yLJy
LZg+FpLoTlfYpOG0OtHlTzwTxn+QRcTOvsifc7nKSL7KhqWP06FnOrJ1MQ+bXDmj
HzyWoPXKNbzX8ciLZwA36VIkmtmrsEiCn4du4eFZVgNOzRiGfuOgIxMsi9FgK8C6
IuLE7QJnZ6Q4aGHBeWo+blZ8A0KbX2iXmMdM4bSstmV8c8DeMmvpLgPfyTDhiFZR
Us2ELIfedaYO0s0yqppsGDam2Yeh4AcxRXfgW7SYOxrhAb7YS/yZUBNcojpcPm8q
tGg45dlafl5wv4zFKHBlcf4r3+TPghewa6ROINW1nE1pv1jJ61F90ww36sW9k/UC
aVDems0bwPOOOhsvYVMTy1fIQXp6K/jq/mE0QpFl4/Ouok+bqqp5kwH34hV2HsBW
mwgT/C+jXGFGDUGJ7wWZAa5ITCPLHBWqKvTVXc+GIBJOQQ5epQaRLnByrgKBICaW
6KACau1yDjvQ2CasBdrqj4pdEibk3Efd5Qmr+IirNcxKGRLuoWqh4kSLlACN7OKX
Yvv2uwOQM9j/9e3N4HS1hntbNbyl6ApwaWQ/QvkAKAJvvOr+evTWblTCTgFNzBiT
Y3d0h6pAP4oryKvi7p00DxDLTyENe/vB1SUDY9Tlxn19sY5DBI+E4Ct/P+6zAf5t
X/pcbV4FKgRyV/Q3smqWtCKqcY8F3t0HmDsqcGCg11URQ1bTrLZdCH5VlRalPuib
fcQHvVEysMQsTNkV9I32l6O1ocDaUrmAUDkUqzgtsxBDjefxtaWb5CKW/cIxip1X
FpuptFicylTwlfY7IeBB3DGS0SdaDGSUP0neNQ4mFp88AFwbb79oT/PsK7i/z2Ju
rvyLP3TnFpb7c8AOLgocmW0jwDn9vDbaPoFfxGJ4xpdvHNPWTCKisDt2ojyOFE+Y
06H55NT47OF8q3CDnZPsyqN7HJEUG3BJ1WJr71vaO9Ug3OHj4J1XCvT6CaarkeH6
lGmal3ytWHauHDV/9ooA6pMFFHx+KH2C/ICKcVjKoH75+FAyI23BD0yTElO84Oyq
JP96TBUm/XgoBZ4kWXVl9wMxe722KGDMaVEhUDDm5RkD/B6Hsl3Rcbv/rMlPjIXO
T9rQWmFCtrOpIh/2F0vylMuI+CG0BSPGDQGDm2i0Eg65y9MWdJgtHih4nvXG6TMb
zViyYEYz5B5OQG5p59LiRlWrhnPVz24bxUi3ZomPcpu9qbNeyNF9xy9xL3Z2ey0U
dfR+Ais3TTQsQg0pHcutSLY8BmZj55ZF6taHuXpG9s+Bva/RgW5gl+Cy3g6FFWTz
uSLW98EWOaCbkiV5U/2JMUm5q2MbKyv3DPtA6FjRb2Vx5k/ufAJfO0Nesu+STtrp
K8UCv0NkifHnLs5kcCDDsgnGIecdmwncLxg/NDS0x73Xss+orYg+K0HTjkioy6Gx
/S5TxLNILOPzgidHnCiNEVCxKbtojdGB7M5y2Co3kxSO27+EGSp6Yr9QjvFlqrBt
400kUUSb85SD/S+lSWeDgjJj00WswbYIW65PW1vhhqujvfNYul4sDt7BjPj7aCDl
cpHnUz/CgkhwUy/MoNiJlkPddqlKG7+KNC/rWZfLBOkIiwiS80xjogiLHeKAertU
1MDh1ZV3dZsrRpaNHHUQYMiu0p4trswiSmoygkNVo5W7aC1+aV+hE6QGFHOaCxn7
cQKDKpbu0hm9YBrGxcxybyxqHHYnUIpBe5Clp9pj0iDecPBPLG/hQJ5AItapmIvO
90ULutV2QYktXD+jE/qbH7O3ZRgHBcDaT8JfChl5wI0NC+jhxewthbvX2pzNHtK+
Z34f431fGOYW/RxopejfaBCUHRPOFN8Z3bJzA3qmOkliJqvJN9sBOuzqoy2WWkr8
1cbcvqQ9KXnVap4cMd/GWDXabYf6Iwu6UigaHU6sYk1PgWQxCGLrBCIrqhUjiy+X
WxZ9f362Vpx1YJQFZt33yKOkjM6pRKcBXqbLinYz8GZtGxAxtlS7CrMv8dKt4PxR
Udcl2obaTqhrX2p/QyWwzxoEtBTWa4vzZl8q9igQxVPP6gRxc6RLtUkDHaXwydYB
wH+ZsNDR5DecGe5nfErTPdceqsqcwPpDlJyImbfYrEVxqRQj+7M8SaDBOtRUieLN
RiLj7DCgteZk0uSqQbJFTZsoThmNqC4/I+YZRuVATfwNk6tUEhAfy25cUnhYZEjE
A5QEUt8Lpgq/tJI3d0yrO2neU/QMC6DUf2nlxLD8w33/hIFOu45ZQTSedIZn7uSp
7wSi4NKHKJ0PmGXZ+xvEb8+4PqUufR/dPeDDENn4LJ+z1a/H9CWKOAPjXw6C9eja
6UDdd/6VM9ZfWNFlFFrBpWPMk7ffTgigbtnC0ofDNdsHQ0CIs4WfVzgBRepi9ud/
qtFgF9GM0xGx8AAJOUGuxipGcTdx9caRNyZqBgUa/Hi836laf8Jqa1yNt9PkHY3+
ve0MfAGpJVBbNLy50g88FxIbJepiTFZl4nxMmXYuCTFdOog5KCa0dQl2RmqlpALy
Ln6Ukb/xY45Ryf6g3FW4RE9LhVMlB6BoZZ45iY1Z+MFO3dxaWip5f1B4y+MuEJk9
7XpXZQMcpqsji1rv0yT+kz18r5bwIIKnbPBH1qIYQkLaIHeKuYx8myspoTbwQKw9
v7po/emX8eHT3VWJmD49juNMBNf1PMov1Zz05XvfGuNiBhQWM7QnbldLMjp9Rxrr
BtQJI4BbmgYqabuXAuF9SNmdTcSj/HjMVXhLTPUvQb3bOj23NcnWk4COyeN70ZyS
TNynf69L8lVbfIremJDma1ec2iMVDGCfuSW213lNddFLpOrNs2+qUs56bcccpzMp
5sbAzF57oSwhPDVEI5waMZTjdivqcR2HZNHrmeEoEmmDIAaiyNygfjDbJPARzA4r
G3VMZYJOTSE8URFOVRqH5ECxx5vDyajO2cnYCA0muVWxvPqhJZWGE2kO+U10NW5L
zys448z8k7cSA8Ycu8CiTudZZ5nQiNJZpt09eY2w2ImrLNzRt6dQo/TZ1ky/eXcL
L8z2tlW98lIgYw5dQThmxGxNueMwRifcFUreizK5ne2NOWXry2vYH9YY9MC5n8zp
GEAfrqrk280gFDpDA4V6uFS7lZn2tXG8Hi2HjCZggLPryFdAi28jA03uY7TLg0mC
fEYwHZXp6q0tf8DJVFYkIVFVcCiFoJfInBeAdfqApPaOPxhIsk5OalhLS+N52/rs
KIeYizpLx7Iamhy6KZn3wRCzFM25Lf/ChUV3adxbV0h19EuZFqsm0kw6KkZYgJDQ
5zy3XWXDEB/WuZUqV+ZNn4qe+Oo6sHyHLKfX2ldSkYdhevJs7nOOcICoK8P1n56/
HkNLL25CjfPAKVh5AFDD2B4P5wkfT1vjhA6Ix55lRIPCTMZItAcmZN94voSC1gy3
Tzgq2qmCac8le9ukiXfjSK4vJvCIENkXn1qa2jjEocjYPnJP1khndGfuHQa0ByY1
CSZssJ4XN9Ez0UyvKedqsN+eDCPWyFbX4C6QIlv2v8ERsKp5djRhUvBkrumLX6un
koAL1mkM4OSLw7N9StUO0w54JCSqvXGqM2bM90R/mLhms0P35i/XTWxhuw6DXrI7
sTq9tepVXpQzJOF0of5tAvBArdmJciG8oW+HeGSoOnzPmnA/pDPe8FmRJO5XXKjw
YMvgf/0ID0IkgiE482gT+9vCkPGaxLI94GivC5J8P4i9dRv5qDRV+Ccf/wsf24uk
4bA8hDuqxmxRTM3AqAUZqkXi+cKyFXdk4iylBFlmNaYcTLmzwnPBKdRK5c09BFsr
dAA3jzU32u3kkSLPuAXrLTIw+N89RhpRakD4K3G4KT08x2GhuGQe0Fq5GN7wZKr9
S5I5uF4v4Dqwk3IUjfl6O/SYUZp+gMzcwIrDNuiMoqN5jHexJC2/XFY491H353MU
hz+LKurP5oCo2nUH/HvW3Qap7q3rstLMXkXJr7xC5ysfdvC4q2jV7PFVNgbLK7ua
Tn0K3UlltA1EIIN1gV8SqCJzav0c7YploXFWghpPEVXETm3MCMRWlE9g+TCvQ39z
ihuELMHD6cIwbo4kWaFx1Rt3HRcm1gMs9C/s5+O+W/ltKwxJuP6hEYz+pAebwteA
46vvnPGLpMuy5iqLwUzRYlTLoWVOPSFkajSNzlmyNjZa56E2ipiVkmmOJAf/jtKI
cLRn8wjVT1nfrVeRgqfeaE9QW/9VEuUyAHseOTodh0n1S177pu0027omlc/WDg0p
UqjLmlbrWfRRginFaxFdkbagNid1/FzFPdAnsYf2+bmgNLIJy0sKl39qmR7elcv7
+Xbp+X7reLqjsQXIMjbUFcrqwoMrKL/H/lJRkX8e5mOGU3fOLVZ/Z8yXl6Dd2FB+
c+duvAM6MoF2uH2NbJmeBVHDvMT/o+4BAoKUEM7dbqsr3pguPXMMxeoLgyocpD3H
XW3UFSY3rSuKFuHh1/GrvlZT8ddXX8JawXmop6IZNm0Gv4saq+LYysMW7liTwtqQ
cY/3uUpBKTrBnU74KtN4prvS8R12NfYflaEzuo2W9VjKC/jgPQ8tVcNz5yA8Jzig
G9aW+UePjBotU8ezZ8wVRhz8T3MJ1ZXKEHGilghpNHsZht5F6pTFpnSRM0M1AN5U
9tThrQCp/5R9sMtkTu7ribrfkMal4fZthGLuv0WthR0Y8UAR2w1D5ptKBJGsgpaw
/dKWTGO86ymJ/0+3B+eyoY5rxP9wrQZRGh5Vf4cBOO6p/m2RDoTdlImkHPzh3Wlp
HDTA8kPZiollX8axEfcSR3Mu2JYmyOXwIAkQpnd11SDLHlwxPY1qyQqt/TQxGzTM
YEcnmW0PYy01+Mvx6D7wo5N/uYCfeLGC4g5VvZIaGihJJ5N/xOarUkhPS39eOlVd
Qhct2rmBa0z7PPQqVJQKv4HkYBRqY9bQpeSFyYo2LowchoS7vT1g3Goe9Xp8L7iM
iUZxuCxLRbYP69jqQr5uJOJJ2UuT/vR6ROvt2F1q3bMWRcjrKl0bWWB+D3nAFLnf
S6qrDfFMdPmkLKJrp7t/NAlc7/V9VF2CvZBUzrOm1hzRpE3yYiOl6IXyEGrqRkmO
Z+KfQQQS1gR6zRHBmSu8KX1IlWP3YIzK9aysGc7DedYNl6FOOHU9aL52E+D4BMjp
UBcratV7SYYdJiXqFglDx02zFvX2UutSO9OntccQIMgfq6JH/eweWtCzsXk9l0TN
qIgJYhxtQsQiCdzCLncwMe/G2yNG+3vGL9KD8de0aNugHQTEHbYAHGui1RZ63j5B
A+8KHFgN+dZNx3IT4MfPDitb+HB+KjpsPDGV4UOglbyttYl1wEo86zkTjGXRbeHu
7RuBDgOek8/IUS3+OfRz1Y8NYuTCCsWhhk7WMRpO0Qyx/5koj9rsvOhWycDpjyCz
DttQaVMZUpR9EgI7LyKOc1KvA6gxlHjmn3aDsJo02p1zWVIKDfpFIxL2sygUt3kO
d8C/eOtIvEymchvM/tPfff+Dw0u7Q2Va2u+3VIK8UrUDen2pWjWOceRW9wknxlg4
OOj0/8gdcZ8SWYLRC/pJ41oMgjIe4oW/uXVAVxfyz1ax1cwfgQ4saveHObx5c+Q4
tLWg0jEe4xe6K9QQ5LDFAy03ROGN7lZpXVMzuuFY6RrEuxVlvjCPP5mefkFy5qkK
Dd+Hi8wp3+cNkFwzgA6+8Yh6ba0fC5emPUM7DlMVUKhaf+C3R0DuBEHhXxxZRb4M
y+riUDYsyyJiLlFGWEaI5fBje+F0vvGavbSKt6pHZG8a7tA/qyOjuJHey2C92o0Q
VQJcmC8Qsw/kmxVsTvyJCAor1R46cN3xpCaO8RfDSY15niK57OjUjPks9SJlByJw
yMXjow+fzv2QSJ2uIvJygNAMwkvP9FQxZEM3q7kNvoosFDudHi6eDCbee0jwAbzN
eofetXjo24f0uxOY2gmyTyD1DqXgUpGiBOqkBuTa5IXY3NNVLPyZ+rHtNDypubd7
9ZUmJOSDle/8fi30kxX7X2sqh3FEVzJzlm2m2+MJevqtTbWJg4IHvb8XC5Iv0TcV
V76zEpIebeyftO31WWtw7clyl4/HaezavZbVVviOt27bWC0qiyg8eDqEa+719qil
zJo4G07LR01oaZwcMcWGRuFQgUdztViipxxqC5dkikEJ/c2CS1ZWvaIV7DZjnn1X
lZk1EVGq9TmXvz0y/HGyVUD9ZF8UNPERsF15W6yOpw13x/gsYkWb5MXdRFM6xbnI
NWi6UaWAbDQgZuZ2hbnKK//Q3/ySY9pu+BRrCchFGetlCmzLZrcvUAqtq4hCYtNW
4bXCP+B+bhGuhTZi3sYogX6KE+oJF5ZpsxmxlN6wSp+c8glfctiJfkiBRPnQjzxM
RiWnmxcdrZPnEQ+2WYDUSetr34COtHCMIcdLyKiSGg7PqWsoPW//v2PiqKrUtxgr
sZcyf2RnENF6G9OIC1SnZMxrBhwbJylL93BCDOCWFWVdziEQWNTw1qxvcRWTJWkn
YO9wVbm4jxTnmmhRKhoqefBgEXIg81Qdwf3Q4QDWFmyn3zM6mJQUo3AdSFRVLgFz
UfIUBXSbEKbLlHs52iO4aAT7tY3LKeF4sBa0nrkqXqF+JGmtFGwqclwlBdNphR3Q
h8TvAJzv1TONEe8OjWmUg3Wl7DyUqgo01F/h0/hpMxqiiWFifSJ14Zc72eym1llC
SjW8qwBqePiK4HYe3448ukLegYN0uBBxrNnlczlI9VKVjav3UxEaunCmc37vStzA
CTZtl50yU9m+54S+vzgMb7pR4c3XZ4aTNcFEObtcJ9lfiQ6W55R+dSXm9ym935yl
U6+H9KH+TrKvOC9qY9212QCacdEWju7iZXwHcBkU0eZuODYPXEu5099WM1entoH6
dWW98wKXzlQB6jUoR8bktP5X9qASpBzcFF776SsX24vNZnr9sVu9wvzu48n+1rW8
KYa1fLuwLTI14acWueuJOr2lOZ+y2X19AMkh6SCQ22JZplUsqkO38F9FKc9slDx/
DvKrz5Vhdv+0kH9MxWu2wv5fr6N8ul7qmnpTTj1V+KvFRcPes3/B3If4PcaQkln/
/hoykb5f2kgjTLlpZmhiTjuhOj7DTDRNLJ2Iq12BhGpDk6r8CD6Pxr0RVkroe+X5
WNslyFhzdvKBa8dqeQzpTYSke+l/fgSR9BfRrEUpnphfwy1z39AClLMaJ9ytonVO
kL1jla59qCe0DwcHc/pbjhcVF5ge0GFm5WFyX6pvTmkQ0fcvJOR+8UEfxfExPzjE
DVXsj9eGJq1XXCSaDLZ7XTCgXz3cYHqOpRQBelx8XRSRisOttctWhiIFvA5YsiaY
7jmo3Ihnjq/HB/zkiAl8ORlQpiawX259N4DsBHzbczOYSARN9NMC2y/OcTCWD1aQ
YP7p13/mnNz0257bVRIkiqAThzrOjHfmRX/5mqyxet6dkhkSr7GaCT9MfuxCdhPJ
BJsrW9kPDLNfBIpdTbkbybvp+9rFORuC49AMCfH1ZYHcBZfBX6poIt/ejg6kRUs9
odhL+S4RiZFUZOWgAaCnvY8NOzVl6Uonm6jvQ7EdZXGtL8MouuaUVcH27grlPN4Y
LrPatE7dxZTYK6VMuZQMcZBgaZNmgUqo2wJSc3elWxmXkM9kzMzLckh1EOdBIqbq
lX9ibwaNpCi9GEgLwe2u5Ovou3IGclOEJMAwzY8739TUuQSNpL4ubeoRJPMwnw8R
mHDvyY1I80lsolSAu1Z5N6A9VoeBBf1QaKJUjwAd5mNjLFsr0WBl5kLUsuVSff1C
6/4pjI5mZweWWsmdu7LhyCbOMJw6BkVh9vkQUBDpZpLxifC2aY9OfSP1fnwRzgz1
UbZQ5jXqXo5fEQuDQDVU6o1/u1fK0EJaNh9PyYdbv29znrGTpMQCKf7Ci9kE13F/
MCWQEx/PiFdQSFduS/wdS2zegelu5Rgab8xThEBQH3uROMPqXWCY7WI1q2502zbV
VPte3imXOEI/E4xCjAmOdN22vpEJSybp5ps1iOcclMnsPaHSHbpvGbLNg7yhRCKs
FtnkuPsAxg5Yc+pKTnQQ15jEedk75A6j07rVDommYTU2amwn5/4bv8r/UzWni1NB
ThVWjMtm0ROma3Iej78wLJ+cK6UpOxqQcLzlO4X3VlzyQy5A5x0oN7O1RxBp/+zq
LeeQaIA/Qz40/sOlHHY6QHGjSjHh2fWShRSXUFaG0zCNMnf45cz2GpZEmjLUWlZD
xlQpIY0wm4djvDTlHRMLzuOtYUgCUhgjLeuNVP/HG5mrXvrcEkGA6wzdxCWYbLgU
FmQs1E5jmFGtMmRFxT/cGDVkQJVmSLD62WkZoesMu63U2iLpaff7Ph5fwCc3GRDG
ng7wFfFP8qLJuGf1dUJZGzawOVi9LitOHWMc+DKyr+1ZQugBiBX7W80GlpdEQtn8
euaQXh5sVmiQSjIhyyFccrlqGqPo2q9Hiw3DvN3D7q0LAzrZ8zAtpa5/3PVI9/4E
QWRS19SqA85+Mz5TAvd/p29lho4P2B81pHo9W+uWv0PdUcGQY8cYdzhNf0oEKJrL
JQcPIioc2O4qcynxFZXRHELeiClk1IBNXTj2uCqdkxcbDPK1kpQgvMaqSSd9ir1r
KBxVALN0ou4+J1IR/LmPBVn0jChjuUnw2NKtG5TNfqWXohgH9+USaDA297nEYmOX
lFaoc3y0Cow5f3pb72OJaU4s/X9mDmbyddmkkepetD6s69I3FjcSp3LWk89uId97
kZx84J5FpXSmdyBBh6DS4g==
`protect END_PROTECTED
