`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8JVqS987TGCUdEQh3f09bxDxWwAIuV5Fz0X4+EwQVUedHui0ndiOmhL8XhtYsDdR
1M/OYUDW+/n1zV1r3jrJuJ2QZcKo/ipWxyRqv6q53mFaw92w0PBPcz6IAHypPofD
iJtBYfrCcA+p9/5WWLjaemiOutZZPImjYpMLffPCNeMwL/bYlA/qLQ+lIE77jqyU
r3uKsbGirX/sKRTYAwsTjeCpU9GdjRkgacgM1WV2hgBlu8MzoF0S608qPn6K978n
FkhWBnmrBzrI9wnAh0b5oTVj1NTk67omC/VmyOq9ZIuHjTSeLhjhfypH20b8FacV
WfZkZ3YCIbml2A6T11UFQL14spjdwyA2pXf+FWtyz16SM7qYPKciycTi4BrAADoD
39mCUOzk5blyNIsXBHjlyr8EYAhQAVgWkL5vm9fNz0FFeKzcnAJu0sQ3+bqFTuVS
b6uZjMi+0tEd5DIKtS341AP4LKieetHXuAusI9OUKMAIFOIOZPqVv5quW6tjOzb6
w7gczE/xkODVCpRovy353dIpXgV4cAcw1yJ9D4jsZ/el2biV9/asnUBASPpclqj+
zSl01n9Oe2HVyb4E89XmNIrfHojOpwb40o/aBtsZy9qDVXNKEttHq+wWVwFOxme2
iW5NIwiy+ATWz4EDzOGKapyUrg1eBKQ8av/iNBAykjCXCl8llW/nT3hDBGVUvlPk
tjwdAXat41v3KIY8gJipFDK8CruxMq4UJEL55Hlq0jL6YxhmSAJYiE6W9LCSrx0Z
mHRbRT1a4qfdE4B3B1/e/+lrVpb4EZcbUm4xgMK0OVYczAfUMzrS7Q/zWokCzhA/
tDF1NDUWg34kbFB2aLHjFYQIkzD5ZC8rUdPEfqXiTBOGacMUISRXSHaCjPn8+m/P
Gz88HqohuhXeBp9VOzKizFxAdvhDYRqTslJT89e1bLvHN8+7J6PG8Bt6eLVkLbss
9WRVUucReRbBJ4oPs39vDC2x6uPekt6RjcbnbHw8L6w=
`protect END_PROTECTED
