`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6ldo5RXUmWX+E/zPXSRioz0OLCZqixoldO2grGCxOIlsGS8m/DogmkOa3tkz4shf
V0f+lTYlVGG5xXBzSrolEu8lg0AMolLgDoYTSJd6hABexp9Sy1KbWtnbXKnTQUbA
rqfhXCvGf6BzNnFXahI2xRGj9y2JklwelX6PlyzQ9ArHW5uG1jt6GpdLAzvsrL6E
2powKsqEWP5GdIl1PO1AV+sor6MpcclQxDxwYTqIG1Gq5smgMW2/s+KRKOScwHec
PT3yR86cmq1bSTM1wiCr1gVi1SQ106sZaDPpOWl8FSSCYLg0RB5w/6fbj7teLsje
eVyXUqNLVFRmx8IgoeCRuk4LpsHXTIArFmsb5fWOlr0PsN2Z+3hMM9+RYZBSlWkA
SiUw9Pjt7/LM8MCo90hIlNJKQWH8Z/DYYm2a+EVPhcBAy7R8ovxunRVrY5px3eIj
7p6KuplOkphHQPfkAReFcHwZ4Ia6eGx0KOAp5KevlocoJ7+hToXev66IPzsXPeXh
EyW4hIjn38H/NRLgkkIDTiAxHE+0AbqNnJkmLtFhs+mFAd6owRgjoTq3vxD4Ww5s
`protect END_PROTECTED
