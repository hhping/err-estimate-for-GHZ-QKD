`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oaypYOKsttvKeItUTjqoY7WanboAYo8S2qB35hfxb42fDOb/cEaPvZiIaC4zs63W
ufAeasQiXSKzuyxBqGzPtSxR1CV8ROXWnwKorcZPET2FoLDhUyo9ti9gf/Zso4hi
HACNeMfFtcPVKdrWt4dXC4UfTsPG35YrjcxZr7qaYcjAzAewM5IpR7FpAqCXk9Nw
D/WCN0yUNHQk+kF5PLgVWBTbnvZlVUErdQuvuVx7Oa2X6pUBKgOuUM8XsMmyusfI
iaZIEWoQoNdI+0Tpbs/kBc+KL1ZziZ3R9SkbVkAoJuJmz0leeGvqkPCd9gEQMREK
BnQCk+5CGZubgQjINyhsBSwCcwd8H/CDp2VTUpNFgOseAVSiim/7RpFR1QM3rQy0
teYiV4FSQ1eZ0V90jJLkaC/6tzWTy41u50FIDAr/je7i+esqn0/dTmGHszIhnCfW
Ty6PKlHE8LG0j/6d7lvX0Ykk1mMl2GBiuQesGGCdAW6NTlKwvWQbOs0pTjgr18UR
YxW/+y6y7lxH1TZrnsJ5gdfEM3SzuvSBjrwIJ7C+1vMlGBibHIFO/s2r/1DMraEJ
xF3tWUvW0C1Dx5QyopKCrjqQcgNDZzT4gfYPnxLa5nkL2XmpNBp2SH6GXw4Ixt+s
lrpXFYff3WIr5WFfT5iDA3rU/MOrUcECt8oNtH4RsC4qcKVmzjhE3C9aKzM10nmL
YItKaue+jGteDrZ8Z6o4vZE7chK6PTMgfhtVWTbTuEAQKpXShtavABwkRnTZra/F
RkiCQyUjXiuNWklIhuTciu0mBQ08JSxmd0cS+XQv8sffiTUMEmkA3JqqIE6Wfjd1
aYPnP+qchuprbpEp7kNWzfgXxqBoPqKFom2uqIRr8VoiWhuqsPRBUVdpRTQO5xAU
PIX+HNNpDlaC8fRwMYRjszjMBSlSwn4RZ6JCUvDo0GAK6gi8BGJLQIYc8od+VZxb
1I08eW3LtXn5eRscg1jd9i5sichXSVi6bn/64+uqCDCUf4TKEqw0n3L4xTXWThc+
iIy0n3uKqyn/Y92XPgTGzkCj26VN0Fd46kR21x2kAEjccQespC6bjzx2twRRmR6b
GL/WePFLsa6oNwftzm21y0v17Y39dw0CZE0rvWzsfdD1VwQKTxqZYhKFmbELho37
SRN+fELgp3lGiExEccXeP2698qiTGE8pHAtH3zvHnSw3unYYhCPxIo+0ehVtTufa
xxTgTdMlzz+vK9BjZivIURNDud5vxF/sy8TtDWSlUSpBrdUqelN+9UEoaDc6tBU2
i5mtHr2OvB3M5bnlbfjKVv6u5SYc2PzqyXRX3sEiWGY9kF7ATjnf5ZCGMRaD+xJt
HkE42wcDev7RPE14N69bZKOsENWZoZPAUJs1GTcLHQ9X+XZMEWdc5EGEz/QOBKMc
6JNaNmgZDHLH7AXpS7SLF41DPVZ4JfF4ihSRaurO31cbEpj6inGQJyjZleAoeiV9
56jQVdYakodv76iHKMJL8j2TZx6WxNxRlJNCkKATxCu7eD2Fq9ABoin6zlSbYiMr
NeDSgcH4fACnDeZ4Eg4er6s3yh3CUeh+rhU8ke4qxqu0+TJHiJdNnjzsII8ymuRP
qCDDn8Z2vkpoNt9jwPzaqf3HOwo98o3PoQM6PTGD/ZYWo4G3rROdswMwxdduJZmz
zEzARCqrSouLIjVrwKl3LTaAapJPCG40p8TGqw4sqr9+zHcpxlBV10P1VysGWbo5
H4PriA/LYnKrRrqV8HtFBTNn7kjj5iMhQcLeaMpdqBiLgezF7wU57AAX2FWUR9VU
aVFhFp5nacW30SmxBirZan5ofEex4QKjz1EO8/QfNEvYIyhCLAmQFRF9blLb6EtH
ytI3QjDnc92p6RJ9cbqYfj9vwO8tnkWDaYPbBV9OfPMELmNo3rULbUNN03MgAKBS
1A9Pl+kPL3JavztPZLdFklhsKs01Cg65jxDttFpBE6lCqOB8l2ymMLDae5dtYtvC
muVmw7RnbwOPs07T9vedgZSrfCFtzN/ttB4KKSDl5JV/BBDsCdOEYP+ks0XimkjT
wVmhfy9NhAEyNFNQRJ0qhzbrSuYb/p5JM+bcj3zq4+ex7k4E0V89adnOMJsIwRs9
HpAUG54hRb40X7/99T4X07L3k2M1kIb/OskCA1WrT1b3JYsJ2E7RKqGboV+sulLd
kt/9lDU1uhwE4vC11eRqYo22GrDea1XYFyu4RQOiDKODXeKbBGIi/jbGd+FrHv+l
8S548uyg/QCX7eHgKGbx07xmrXQUgc4j43W6DPgwxeojoa+Sq5kDDszOnXTtFqbp
61XfYeos1cn6LnwX5P5sKyuQjuQ1Immrjd1Z/yZth2gmfD1WXBud8tAxpa2E+2od
UIOwXBE3wchWZR69Wv81wij33nnjwwEwNJVTL3yCzRJiIs4D56Y4usQBz2j+KmmF
+1vuiIqgrJ1dHYURNidLfizZMWQdp3EHVCz/M3nou9f7xZg16XFhReJSbtrTz+gS
a2We8U4xWbNOR0rbuOaZVM1IOTdA62qmM81OaWutl4I7w2nAJlRsU4on0M73psDl
UzV0yWgysnzobL657EsqEanS0megaBxdiY/DqntBMN0y+Hg9TY1BZVCATPlacjaw
XynMJ9e052k0lsJPv7NcWh/g4IOpzg2gnDkrGv1ggcEl0hlBbMdvRovD5vutZmrw
XhCfdl16wOwunOgrtdua1z8jBUSWuzGL8+Y9lhptAHQSvCnbF23emv6lCxglCz1M
sgMjg2mAE5CfgwXiVkSC2pGZzjN+kwNU/r8+BkAfzPd7gRazvPWc6uFOaW76x1AS
E/vpqXV+ywkCBi/mjPUPgS8a1FCGql424Bgp5G/uvTFey6nMFQ5n1MWE8RdnD1+P
Di1s1BsusIDXBbWSG5SXtUX4ubRLy+j6DkuYvmPj0YiNaHzqrZ1GTjVIXMnH6jqH
qGww4/v4KXV/ktZLKxpiDpq+AzDGTKhX+DrwX7fw1tuhS6WBhMQjK6zblInL1ms9
0aNz5tGNFwP4C+YnmlGQzki9Mc055VEduXp6/bsBukVUvVptRsKRjU/Kgn7PRA7P
8zxwhIirYwg0jt+2NHz+Ng/SL+WfLZnsIWiMPPvTc5qeWxp8t5JwOTsDmYOj1UaS
6lIAb/PI49Uuox/o7ljQS7FUr7j8jd6XApHPvMOFWffZpjjAIXH2cNnHsFrPzRVI
29DfQ8O3b7kt68TeyP9ioZZgMUkPtmwgxWBAJvfiG3AlpNDBTucfB/6RKF2s71C6
CoPobosmUUrHvOBznFVQNUQIv00+DG7BS6VxvNommKxCTw2wTnvwIU3KIvkqhAfM
AbNxWUbxpj/bSiHsz3ij21iNGp+BQpOPqdLi5AWPNW7gWEneFrM5sD961BtSYiGg
sb/Ob0wOHKkLHeOwcuqhZc7O1DbPBqtF8ZQyythIDdqKRFnBOnO9lgsT/Qacmk2A
99/IAQC5kn+at0G7FqUSMJuYKWu9ML9FjNJ4a6MA/QZh2DVys1XYB1fSzfuJD9r2
cXcLoLMwXKSU4BaiSegWXk45sErfBCjwtjzKFf4ME0q0qOnKXNZY3znkH5Bre7DB
kjW98ArJMy/s6mXXFhh8ji9wVl2qLpnJc6uviIZE5ZoQBIgg92w1FTeeZGu1axv6
T9299+Yx/EKWS0lrKJRgCx789DvaMYiE9HKppQloMsJYdBBItyDDMnWaX+FqEsb2
NEeeNcAlVZD0jh5JLn/oYpDZLJHUteFnoCEo8JupnHI4LzsvFqsnLB49IEft8o3u
JmXzmxOXZUXKWXRc9SySQcawQqfJVG6emvVzE10FJdGh/MGdO7yjj9AcvHsKNNwT
9Za9LdhIEkLRtk0zmP54Bi3DR9vkEAS440Sg1TiGfS78w0HC1h8UTh877tRYSNHZ
o7DK9C0k6OMau+K10E/iot4CFdv+HMYouwNEVGEhhOck323viK6Cxo6HM2gVUTw7
p/JKXU/DaS3o6jCRBXvHe364odAy2xHyaurc4zb1xOogbpl45ru98XPTSdMqqQu8
VcowFln8tIBf1Js/MeamRTzFkvI4nq6VU4OQtYcDGHPeQEYbcQNxG8Diz74udR2u
qa+iMvgzaV13VziooQJHGENs1H75Z/64HvXImPjYnYjkot+xNpnOWj9fWExfm0qN
+wc+Wolkj20VxsvS+606Qx40Za94XbABDm1Mvx9bEy0HCU/KQ+ckxdzYiw6eIegI
dw4iutRCY60246JPQ7UYXTWIpmnzPC14wwRAdfETYyl7Rx1SuGLlXaWA8N7ertJW
qxAeVmZ8+dN+Wm4Bi/dr1ohw3CwiWrA9ifNa0DZ61YJ1i04k+qdLvA0uxgiXCvfK
riUdIbIf3TR5Phi0dxa3osbMAMEVuy4pNmnEzBazHVIrIqSKSg3KW4mxj9ynzai6
Zro5nRXrAC+5jY+/Y92jyvKZsQZFo0uCbHU+ZxWWIPB1LA0dFcs5kZ/GdYcl0FXm
qbSZtrqqSyOoZejwvdimR8KVcmGOv+WSbVZpA/VtditcQVbJPKwsLXAIr7qeLr2y
khB2rt+hFaD30z9gyJBxBUvl6M8SDc3argduWJOnuhv4tQ8IxYjNj5f1YW5aNlLv
+JI7v7YU/ZxAc3RO7GmiD06RB6gx27EubCI07TkTHRIXjColBKWHJpogeHF2t+cB
H+HytEn3x0tLphQKcye9pHHIzA2tZVoBcAR49YUTsJSpfCPL4M3XuLwD5hJRbEwE
310guQKVw1TO5bVo/owYhn+elSqSra+kyiuLPxJfWSccBvCZOzayLxtoudUNmWZO
jwRGaPBcHCEVTmKjvCEKA8cI/IxQjzvfDx1QwHiGCvNYXP1fxu5X7qQ9nO0ng9xO
EnwAi71aEBrHF38BMFxFnc76eGTdCtvBUXyT5i9rq1/EGljIk+nXjocB97UIXmCp
UstLFMd631ItAQgM5v3OVQoL+NC/zPso2ids+knqrhH4JurkR1AIbOJqRMrs9S2R
ZaxveeW5jncQyam8edEevwcf32/5rv8ByMjh1GLkGVJhIb5Ce/L5KHt4HaYh6gsE
gtK88DTp6BoMbvaFIrQ5bJHplyVTEhXI38lwG4AszRffXt3DyfBDb6pXvRw9PVKP
fZkRrC946GI1oYX4QPSxyLwdXbRLGFQa/zzw9MF3oOhu/sA19eWIX1dv5VZENZb8
FQ4+23XAuIvfXtGqn43ycM2jzAPWH74k3cbH+3O6ea0k4XlsEjPHptX58v7HIt7b
7s9BS31MyIB4vCws9vlrK578K6sBpGxBg/hh9v7tya2qm0iiatvPfgNvoaRrQhV9
RTYX2z5gv5zYKEdQKAb8bOBPt7H526SmpwZkUYhvyG3xXe4EIscv7F7AXtNqgksv
kXMzUMmjCfsv+TsPZhFsf7l3v9kzvVfJh9MvYD5aCb6iv2b0Nj2eyWgEYwp2X6K5
He5bw7U5IxoeBumlIW2zL1HDskuXzIFBviST0v2OunWT3Osw4pJ6nFaAFE+oZ6+M
kwb4tOb7VxHRCVdihWWvY+GdoidiF7mGJIgpIHiADWZcoawb5vTpqXW7elwWRDu4
uit8mMh2y9tsEAwD7HmDCFTuhYtD3dS69/andT0HUdYTTzoA/Zc1PbHb4iIbfvHd
C2ot024xw9XC97pC7YW9yfeEri77rClIT/MMU02ptnnDRzCYyZLdtUR9EhJkvpo6
mOXrcLjBJaQaZdie+CPXh24dCZKKHGoewNkyD05u/snvQeyPPI1sR8vH+JZETnvf
Sp5mRQtZGxf7jiAWARKFLzK2wVTX+JDLP/j3M65HXzUMKowpKk/mxzfrdfqKi1zg
CI2Vo1mVqKU6o3nunF/RVaxJGW9gd2TIv/Bjnu6II896mI2vS7Mu2ofd9X1+t7WC
qW1mmqE8VSFHpbMHafAHWE5NVmUFX5ptd70d6e94t9TgbLL3aEGYrQqGjgCs+ygQ
gXm54u6Jrd8JGhkoxTCb0oZqBR8dp2d85g7sgtiAlv/+JsKPsMU/Hqqc397NxiFX
lpBlTA6YpJM+I1d7WT6XacsEH/EMWI4r+TtLs1J0VwIJ2kp/q1zZYWbPwgri9LqK
bsORo4q3IXZHSBCY4AzcvWqRSP5FjuEb7R8fPkVAAdmZdXNvcdlg4SYEMOwmGw51
54h1U3w4Czm6tkNQ3R07DWwiB30V8gXzt2I8TJHEjA4Tg2H4IiutGni/p1PcppTM
paxKGPdaGvGV9DsvxiWqKSwFTTj1H2E4jbWhN1+iFroYU2pwMQW78DMjS2p0GZSs
tqZmhtpZmcC8QVPak/Y14DNA5zQ6WlzUgHcHWVCSK7wx0rc8MfGI4SIgpUEQTx9X
9xxWvXnm5uE/fzexj+5CrP8Fl9lk9HUio0tPgmcTZmzKN3k9uuQg0dPv0kTL3RUs
5R1+kcmS0AoSiFwNn4+eOfeh/qDagsKvBxfnReX0Rp/AufqN6e7i1oRmjzy2Wf+0
aqUdOfuHO/v9UxbAv2+dzjCWCLTvjU7XL4w60OcWGftSlUMSQ7HV4TFAwj2Uz81Z
lehIRZ8Z0rrai2pV+9ibLOnTQvP+WIWqEQgLTZdOjRd4CNqW4wijB4W+RDqSnJO3
guBtikEHEJr3CLwNcxPq73h78GzmFb1b5rzvGKzhj+cZUjkJPf5m5bY8r7ojrGoJ
lAKLtkr/ojcUOFV6VeufQljbTGroo3vlrWnNjc2ABU1PvHavWRH9re7Mj/itOWJ4
BLXcBGGRSwqFqSy/s6oon7l4D/uuBu3itDSxYksA+sv+Cid1V8+mrgaghYMdy+9N
VlsuMUlsk4+vzGYqHEi4oIWGloxhe6eNzpK3/4FQ/XDEmHzHVKYBzwrxO7ABvrr+
asVlcEY4Kayxw2+fVKhZB82OHbckSlToP8zWTGUjCXg+AszCaLm6C96XPFtpT9PV
M6w+wHdbdy6mcb/WV769lS9CqtbbDOjNTk1jM2JZYUyll6I7fxLqVSjpNASWH4pU
kFE1BaqXkKIm2s+gSQcn+xcbouf8F8u7gtvQpofk7Hls7NfpIwhAoj4Tsrwo7PHU
aCOglIF0dTvk1qukhG9VADLBeMwh5UaFGJkUrfUWG4SHPkM3jANCn2mR6Dzc9z3o
aVKyF4wthfqUjYwCwgGQdRWlhEHuIU97tHD3Vt903Fq7beQmIBcL9Yb28ny0ez+t
tq7WRpUArFL411T1ees425h/DgYLY3TeE9RoWw/3F9SFqSXNYJd3s+zYzugSocw2
HT+xxnnO2mlMcSD8m3BrIQbzMn7PWr6xbwaYvfvzIsDXSkvHz0OlX+RWZACsGzk5
qO51vV68VOa+ksd6Wk67H00ORBS2w2hzeVo8HRf3drUDX0QFGpC020fU4bsz7dTR
6Bgz6Nd0cMTTFfISsIOBtuk6rB7/GtrAOHMJBNJ6sMtkASP8UuNPer0F0PO8S0sb
RqD8jzUtgA0vk0qOaumQ18iBueqIGc0fIwqWvYl2OpMalUhtPwqxBnpV3yFnH5ci
X9K5AKqO8cOY6KX7BeRxcp2Rx1Nmk5ihq7yOUzIlvrPb5JseraAWAfdUFstB5yDW
lI2J+ubV5XHGmsRf8zmTSjeA5djiHrkFYkTDxgsL6m0vGBmFYYRmz8B7KRU+rLbK
rUdfcIZaMXT3wDHL6aE1oAFCx4B4YCkBl7DiCxx3F6AlLMOO2iEcrEmKJ+GgEa4T
rUoMAz8MylhnO0OvY2xV/VnYXXKTzYdQ4resWz+Mq8xMwex43E5vCeLquwJP3/Tv
+QT9ALuA7nQsYd8EiMVMUPyeFcH7BVwrQBFaCF6j1fpyMU2UnjcL4XlUAIErNFaN
arlSqcj0c0lEB+LibJ0pzf7guI6oZc4nbxhHzP+x5APyZ8K73pO15kNdAruZqHo3
XAwtalci/LJ9BVu/ZbjZBpN//99ThApt8ViqzpBkzfGKfBlqOuvM8lmLNEn2ykpl
jLxKwsyPSt7UwXUuC2XqcKe4raU7EkLL6cW0maXqndw7JtU1bgl5eTO6O3C2+zQU
AW/d50UZMb5zFNo2WrTESSuOkdb4kUJMBhPbsKlEcAR9CW2DYA3JmMo40UC7KKXw
73J368B0rimU2GiJlBUv5VOmEhPSphkJ7Qq1A4+YOzKgM/D0KlFdaERy7kM3rnaF
hNn/XbbLvCnr+MD6CXHHa8/V1nAoL/Y8mAA8hnhgVHvhtFms21qjkaXwKLmeLafw
eWNRmrlKasZE1JTdvGB8KuvLHJS+Gu/zKemYJA6Z/eznLv18ZEVVSjrmdns0gscF
9qow41DMwNdtd4H/csaEr9B1mgzcHqdfs59ntYkOmHDHhRTyTlxZgczRV85l+vCZ
PmNU3lITXJPcATJlpye30cnv3kVeRVC1o1tDMNooi6VhCsNjwPCWN39w2g9yGBw6
YukOga3u/g7FEbHzTvQdNE9W/YX9L0iVgpapTp1cwN5sdkgdIxUt1rzsumenehim
G9Pvz9tK2ucWpTr5OiXgjKPe55rpB0XT0nHIEpE0xITt/5a45XhG/ucDTo/UT8Ho
ih1ljnhmkvpmQwG2p6rEO8nkapM6Uvlv4MtnDpwMte1+Xmsf7DkeinphLQytW4OE
X3AtnAYOByCuCmgkbZ71UwuuoEqYroVs1KS6+RPrazwE67Mp0TT88aF3PeL6EPtH
DbfCjyiaQ1Q6Z+ogv4nWn9Oibf7XX4StHNnaEeD/l2JfCUYf/A9uqjKl/eFIaY0e
msuJXybkz7dGbMpwyZPSJ8bL9aSFpUKHykmE5qSmd2UjMT1WkidNDaQ9YjoKDv8Q
9NpzVD5/ShL/AyJIqoSlh27NHJNr1KVhvOkFIGtKaOdMvLeFAEZhHAz8gFClg7H0
AIJ/nyhtFD5s0S9ExzFvyUIyfdOVNulWCDOZXUCcmzqmZP9XfYPe6RJL06V09WyW
CObSXCUAEowcMUlBRnyQa7WGV09LqPNkxfH5ExbQeqKszyatFbaXbsNMz20XrK49
DfD3kkNhBIrKkbi6xOsuTOYVKekjQx7j5Y/9sBKbuWYfUQijZDlokR+TiRjsNucX
9/5shNALWBRJt21UWWUE5n95ZGdFEO9TvlD/wYc9Bo/JDOJB4RTch5sjTPqLCwaX
NOuiUO7yYK0iwqxC1kMIjsAUj3hkuUK6MX3b7/WdB64eXklrOPJzMkbFJbfQTYMa
mm8pBDtelS1/EIXxY49xz+q0HwwH3JAIOZUm2Hl9rmENv/Qw6J8vxUlZl2Ym4dnw
c7n8jvutG5EP/g65tTleB4ofX9Y1MZN6cbjdt+nbTy+4qwRzI/5lWiLHx4myi8eP
jGIhGVNyTUfx9026ktTx3kUt+1CkpPKpkJuL78pKa7zaNVrTGxGk1IxElDDBPxCn
5URbiWnCQm3ZsH4QPgYYH3EYLQVg3bdRiSQxJOV4z+0cXbhEU/mZuL4DMSDiZ3zV
Uw+CMyOVQf/GQIXf6eNOskzWXjY8yC2sApjDIlHaV9voZYKe1CETilKaWYmFH0Dt
g7UlS1A7PCp6kcPCNw4hGi+c2ZSR9ShurFcsJ5ROVEzWYrSjxvZmI7wBfr0esFeF
q3mZbDyPFmIs8nhfHmYzsbOVO8+D2r5+c+R0kGi7piGw1gWT3sKkxK3kgjqgxYQT
t5ZTaSG6W4qd9IdMer3pufyWyiWqYJriN8TozLnwyaMCMNmu0u1uGa/2V1BdlpPk
Hk8a6IpzRQLAKItH9Za3AkKm0NUa5LbqsMkWVJZYVoWmFB9XRu6maryeATSJ5loc
Mwxl8kR/P1HbzzjjFcUcEEUdGpotAuiI5tTPYy8Nal+kynlJUFYJZ7TYiOx0GuBR
DYAn+ySriJiTR7J/HrG/hPLzWh1utFlKDp/G68yY8ltdQaXtVhQlm2PRgHw9QU/2
hSJ+Db9xVMHpK677jIZnlukvaffbwzBtXyh5jHzhBOjHB/ODsOa9VUhvxSDu52vD
zhhm+Y0La/VP2/mOlkCF0EEc8PAWn0/EPiOR5wS8nyrr7QBtbf4MsZumC3YMk/6o
31iD/hJtugMYTGc6W2vdKG/4i7yyJYIy9Q2FRseI0SUmImzCiY9ZiQsZY5rEIZp1
vSQQRO4xErC698qw8nK/nc6HDc05WtM8S7k3nEIzBvygBxwh/3YykwaoTj4ApV+H
s79La/sSO4A9/Y9UTZCH2doJEgRJDzsGEADg/DP5vSdTFNb6FFPG3B31GvYUhWr/
RYGeXX1PFzD8a39mCel546EPwtThHJPaY86shri5GVwJxGSSA6l/26hk8aCNKS4y
rb/QENLUhX9HHPxA/fqwbFUpc6WX/5l1oUAS34SZjqQ2kzs2nkHnXaWkYWu+yaEl
D7BdMGNQGOGUjbMYue0WJu4evqBhSlaUrPYVqHmTM4PsxyTet03HnBI48X4cdcQH
V0omob+q9rj5zOtOwyIhlLoByQX6dnPeN4K40g9f0WFfSW6yrOoLoHu/Hldlyx5G
aMxx79sboHkbOWfH2Bbcs+xfbZXGxodYlyd+GyeDjIhEIpdRzvNLp8b5EkPrbaO+
AaO4ZAcSZaXrHHg04dum01btVlR231V5lC4N4phwovsrBQ2wkXLPurPV4MsDeuyp
ORSJZAueTJd+TjihjlUl5iO1AROIVrRLBKLtEFcH4EJ1TuW8J9Jif+XlS+mT3GCD
1+xVxY85lg67ejGurm2DhTnve1yO3xvTEjsfSBVFeYXLBs2D+fe05X8IdVCKD2JP
LDvry1iyLCYD+C3zv3XVJI3uz0KA8bd08w0qQs7fNox/iwk9lfv2Ebl5zjtcMTwe
sp+VRDMBFCWjMxDh5S/tCT0YbZ+hcaC7v9lKosJs38/EmHp+xR26d0hTZwc+Y54o
eXcI0B/KUMF7MupRGu7/F4iyFYd5L5sm7J9wGsR8KorG6g2qATINruaajUVgTgmL
nBvjbIRCXgd4GgrZwkbOZ/IqNeH1OruYHaJ+A55jx+iTHaQuZ1ZRJWNW9J4FG1hJ
vapj6bmOWNyKUhivKHscMz+F9PPw93nvtVIkZvLKM/DG52CWN2Miz5k+cLGMuh+F
5rZT9uDOl/ldqmddbBSBHZ+ShkpwmUINpOr27hqus9Wm8qjkuxYjep+lzOs92o6h
X/0NkAM8RfEKg7fZbbx9hMCxwJ9ieTUKWbrV0G3Zz69P/jRAyckSJGGzGq6SBY91
wxywJKCm+rGO5+rQwv5F5Cb/OzdMLMV/G7I9iBQHp7YetcNDNYPnC8GaDSncR2SP
XLRHHKxxovddfggTCxN9FYh0Smp1fBdL4LMHvp8LwA9/aM1EotgwFFfufLJJFb8Q
tJYy8JcfcFD1DpP9ij/UgRZJGYb7YZ36KSLBM0iiPZ2dahb+UF37TtEajIMfpjJd
SEi9HXUL6+tKQJhZnYvBCoJgNfrGi0KQZyVJRUT7X/tTd1UQHZTYhZqr9H8F2r9P
vL1MBjhkfjp1J5M1bo+NVSNdVuLUf0C3gvE0CjtEdzfKD54R2oQS3XN4+ZL1Chl8
WooaGt2UAuivZExKWaiFTBr3uyTY692LDKsIdR7L2UuZK5Fwti+WCESSAPvBS9IJ
NX35QHLERDMi2PCMEOgrtXSCPxi+KshnlslWKxGR9/KVzz16CBqs3LFPb23WtWB9
2L1JKfqCoEz2HjexOzjyUpj9Ra3lHJkBttW4d18VY1b9786yXyvbh2fHKk+Trzq/
SFaRGiEiGwVOQCjr9ot6nSeGXrr/co/bPoLTuNBDzemHD0uB9L8IVQoZHaLqOmWj
J9LoW8Hof0ZmaZ+KkJQfT5ih+49sB5n3P7tFs214a5GFptuqBi0ZsCPsx8Bz3VjV
xdmF7SXHdKXI/z6CA61ncUyYdEgJZyP5gGsimqwOM1Yt4HMfGdeyWI8xxaPWb89U
LWtMWg3dreFVCkeb/1Q8ke/yoLiIvsL2IpijEFsYX281umEGriQVp+vgUKzE4WAT
Y00gKo5CY4SbY2LhN52kBvXZ4zXHD/WTDhNDv0EG9JHT3vIzRd5Eh0cGztTI2Hmu
IC5RDQe37SQhiPp2PWt71/femIsAhtQHah2GGypIlLfcNU9+1rLYN0p6J/mcnTfW
+HT7KIyE8Tnt/93RGbyLGLUaXZfYpnB/VkeVCMUIPQj7uPlL9ifUq4/CgO1+69td
FDNfJ9v+DsJHy5B2BmL9lv0X5yEPtAfLQPB+aY9zASwd4z5V0cFzWWkf4gntHx9z
+ac2AGoCMvl0lNVIV6cSvzS2CGj4rCvcNZp8+0qi9Bf6+hwbeW6TVxlzP9QkcoxX
ubHbJLPHsXA7Didqi+0luCvDjsEqzCKvMMErZW5Obx0Bsb5E8Bz71dTg7w3uVAov
K05zwhvpm9R4wKYmlwax5rjda6KA8oqJf3qFp0t5X5Q1LNMW4L9ufsgLRIeNip7V
WuXaJ8WGyWHvbUesh/7GapTB2htRGU9oePVw5MmVaheJGm1x5rFJrNJU54Tg7r5U
egQEX8cl7n7jRjhaR2LA67u5ci2y549UZIuTD17ag1HCQRc4E9pWVMAbKt1J2yER
rAAfGyRcMlPhQ+H1lrVxx7UaVdJiq6Oc7j3TsxIYhzMfE0qNPMH/X6Eyq35V3rro
dlVzb6ycKi/rH+glwFCK5ZJ+FE/aQADEBKq3RjCfudZON6/X3KvdBKLEzG0W5F7M
QTy0qC9GANEfWF/pBBx7iam+0Enl46MTkRtaOUG2ojRBlp4PYuc5Tgrwwttluxoi
h+x8udD9Wh4XlfrL6wHF5aF09AmreWoeUlrZeNAcWnbWlbjmkEDNUgz9EibQpnLr
QBbmAadWGld4dgy/mqjjodEeQ7wdvTVjIN3W97BHledztMbqS2SUlGCmX1Snbqbt
GLveIuhn/xIuXnoF10AYNnWukdBeRcfej3Ts76w8arENfE1GaMpICeSt6uOuRb5Q
/yJG4Z/Bwl8nTCYjo/dlXc61p9967kEK/spDo4uIOuqFzX2NBpHuJIREOIdsGqDO
U5kkweC3oAZTIepK8pey7YiI2sIPW94HmMNUiRZ13fNaLCx+kd6f6hOI+YbX5ZYh
O9HL7dqRfVHVbXKbnqL9J7MopSyeJu8ec2CKFRLXhDyxSW9u/Yeoykrx1v5Re7Nm
YA3DiFsr8hflVtbdrXi1G5SYkjKKXTWJaqb8lwFKcSGYc/E7KHRIKf6+3Mfqz0X7
L+jke0fNW78zHcYXpgPEiCllAhV2rW7pkRtMqxjJQOHskVOZn2Fr7IMeIRakTs/F
MeSEsuU8fhNOtZ2pcplkrricdpSRyqdt/eS3m6zv6vARwj+tBLNvIynZzScUjWP7
CbVt4zrYthf5yCxP+bM9dl1BQMNWpNLWVBeRUuEBPTMPPaqiW4trJ0OG33A/n4Ep
by/OsJZYa8T5F7voqoxvZLCL79lwkn3eDwKifJeJBu9O248qTcYS4BylNmvfnMBO
zZW4gJ3kcSYm2ITSUHgKN0HP1JqXOJXZJMzxR1Q/vxW6OAqkqoZ8P7RlUgesljpi
An82d0LlPTX2nUPKvYAIe80ZNI/cYP/Oq8ghQkYtg0LZvTqSXvYBJ/DM6Z/kn3P1
OxuKQ7fYHkaIzbX4ydEjTTFKvZqCqDVnq6LE+zGjb9WyOkBCtxEcntmefeEVmWAb
1yYfYoKBcWL832q/2mDvrz6P3+whS9CCoBCD1paCeQQ6Tm+3CilS8hZU/6V3Ee8d
/lIbW7In1RNKrjGcSoNXQYZaVK6OJybuXkV1IDZtzHr8lpkRkEvLSHhTxvd9kTlG
CLEU5ykXKUTKAzHZCu2DQoKgQP81ZESmbGJ2vG/MI80lbGNd+em0MrfdB/UQTlJH
bZuFJEqn5wZRlEsVTRvcimF93AyNpchnXHmqoqGbp0tu1RGmDjdW94tEoU23SDZg
4eZkurJHZZLyodgg3+SzCwPLRdWbQNGfeZqy1Lkv+Vya7rgPh8z8dQ1R3o4vTMcU
U8NXOmuJ0Qk1ZJbj2vbPbTwKJP1EqKJ4Mt2B/pamrAebZ/m0sIpJjJuotBoHbFDR
vFZYfVjiYreiShkZYSnpU5RyDSBbz4Mi3aCyRuiI5Nx+jNk/t7BhZTrKO8oQe1tk
lSJ0DDxbjpHckuW2J7R2YXVSRx0Nwf0gPcQeoG7+d+KK4OoI/Wd9bt46RNRzixnN
aS1jllC/0CvQCT70eA/+dbEzkN0G/ptnvmvTPY7a6eMEeqdWJD/HENRAsmaBCbSy
6PpENgEKYHDefpz+WfhM1wkHniXH85Xx/YVuze5ny1PNNBXUpeZU5xhUKVQAnd4B
4WS2f6Z3WSQtJ4j23XnbPKQ0MG+V8u0vowwniQjxJfv5a3bD9p29H2Y/pjrL4BIJ
cEKqMjEk0HW5fjRWcV2xJhvoB7E6beUwSsSaANA7UgaFbP7Qu2uKcnLpgt1nH3K7
TtO7Nvt6AtdIdlN65rvTWFWJ5efUiXg4zHJcTRyzKDGnm/oo3IBmepZgiAZtFgef
lftOz1n5TPrRiigYf890aWzge3GMMhh0/ZuJ7qP/zqowOjDyAbMz+YCWFOvjv3Oj
lL3oZOc1fJqt17JXujHRQp031NGJHLEOi54eLe02enoq+UZtIxc3pcgmprvqUg0Y
gMmICvfh3dC60NIfLPGwcvYUU4sPWWmNkCTnUaMzAXpOL0iXYNvwQImYVQ/BSVN1
DEE6hhGzOFKZtkYbVt3X0cF8Tq3sJS0IPQKcY/TkArhAshF2vRevg0O8hQaeh3aQ
49Rx8syrHt7p9aPqdVJxaqeSzlU0cJp2XbqNC7OFoAjJZ0s6tRxDrVtwlIW4E6Zu
o0uIU5R/MycG28TdDltrqfaWH2s1xK9z5JuyEh4DVUiMOPiY5IexDE6Y/omZAmJv
X9OdZfGPtmsJZbRxnNPRm6J/5RLF3Tjbi5aBBlLfAmDaQ2CbOxHKa5lRBqtkue+e
XpiqHRIgJCup96MYqYaGffABZdFW4vMPYkvCnRYyLAMvFBivWgf+ox4+nj5YeIsW
On+/ZrLMatf6qoqPXJbRrULZH99qFhxRekYPR62sylF+1W4w6/8Wp4g21JvR8m0y
vNpyHkaXtHLolMzIljGukUm+0V6DC4p3Ju97Ydq/7i6UswSVBJwzkxJaZh0xYOCM
YxIORBCrP7zw3mx1hX5NYMkEv/8Kx1tFFi4qSOJkdHsW9/2GWKRFOnO7mjq6K4gq
AOPv7H0VA5IoBbPia25L/igsxXu4ZUNHY1vR0qQuFOigOKXIynYPq3eTE2VuFlkU
5FRQw6dkElpcWbXKWy2eJnWejPiIotdbpBZc08VbAn610YA/+9OgAM+h2bOIGLSa
9/Gy6zDyARnzZqxvhSb0rez7dgsv7XqdKXqqozV9YHEIDl4STORwVKNxLFyPKqgR
wdFUnxOnKSowxrqUD6FIK5u/ZFXwU1gM9rJAgT8w9UmbHShIu3wa+CJJN8ulyUH6
TPTxdld7SLuUjJN8R8dIl4OXMaV5xu9IdM6TevqaNZBd+mKvlMDBXuLAlMuB8Pkx
8cZPvCPKfps2e0rpkQLfQ2B0FaHjjbCK9qtSgpEc9kLihAFtf0LNgesWhvpLaAKd
ByzOq1g7aJAutU3pMZ37C8caqgJv6QA1D+Dp7kjRA503+pzYs4aHGh2sPyHl1LgK
2rigNtCwZ67ZWAG+vVrY/QAiiLS8JDSIZVTT7BoiRg3bxm+4nqAGMgK9mg9jN9V8
kxfGKX8lR2wD0gXmkxUao0HyvOmI1rdn1XanrW2swiGCYpFqtSe1U0nGtMKcn+sP
j3cbUdyXm+YYwRxWiuRZp9l4ikWVDiafNFfJvQs8zf/LDjfi0iWX5XfMoSQTk7fD
rVR2WoX4WA8V11PzZKdXy4Bq7FFJPqk1D+QG6Jr+kKyxFha5cYHzzpqgH/FOVbsg
ceK3Extm/pBnyb3OSryqLPm2ejfBtQT0PAE625Jo715Iq/giMfGgx8qZ6kH0Ipp+
grYFqvmHd8ttIaGkhHN4z9dBIWjb3QohtG75amBv4w/YIuleteY5PHQ+VHes4142
2McgDxTpY+xfJom/SsHnqGru3vYzyks5TzvedBmHYDMjbpFhHlPldExls+GmPKqB
83atDW/5nUD6bJfJ2V0m1yTHc1WwLdu79R3pLplfs+9DzF9yFZ62EQehrEA+pOsI
zxOsQ8o9EJuxhd8P81eRxwFqRKrTvUxoKnDyhF/6B0O3iNKPiqQuNIDIZd2MXBjC
jBes+CGsDrTRFumPsn5nSRBbDfqqad0AFjExoc1oiss3maxxWP4hp6TsEVRUI+Gw
l/ZVDhggd5Wvyvnbn2yEUbjHsf4xSpKJEEIWeF9rfbjoP2mn5dPf9nUuM/l7nJ82
TZDzpJjHoLffueqLTQAVP57YtuqqrO8k7AMNvE6YuZPQ64tW8WWcbyE8flLwx49P
JeVx/DI8s8kkFdP0CkrwDna5n26NV1tO7KbYbc/F+id8CQTzkPwh4iME73oixsDp
23luNVIFJUFIJH4wnZT4jwQJ8/OzPjqtcdWsOSpIj4fZpL8ugI5uEsMSyNaH3MyD
oZZPyN6vvl3t9uXrE+gbajC485jbrsIZGyNzwJPkDCy7tgaVyRarJBd4S2aufoSb
GXybbg8b7ncI/UGXyuy6sPVxiA9342zda75cexFqpjTDgo0HpwdJuAt6L2I5FAop
ImaBPXpp8a/WW+zvllc841ZpWuk0O/gJc1JAAcoAv3EUuIMc/QY+IWVWYTTLlS7R
HtSQ6yxRfWOtQkrEL1kCzXD6gBWygbsSFhopmSa/7MUJm2XI9iH8Py7eqr8u8Wii
KJQthJH75U03ljzkBeP/K6wxeiuBpI74rMHUKbF0Xy0u3OpucCteVccKnuW+i9S4
kDBLY/ScdYzZeaT0dxZAucPV7kanPqMqZA4HTHgwteKl8u9g2Q4GVglpReiK52AY
t14lmu/qVpkiSTScTG8SFDx2H1hz1Mp1B3GDoOidUlA0KeeMtOiD7zRQvZVXDQI6
ilgeoykpCsatG45jdZ9GMWpr/rYLQzt5NXZK4Yl2fKTQjpwEPQaLok9FZI8TuVzW
pLKg3J1zZgiOBYDTSz4PI5wIJyvnlRSHn29R25L++c0DAZDCe3p/4YwkuIw0v/3Y
8rkn1P7OfQ+LH1dk+vm14NOHYIQriQ4y5cU3BVJDD8biTUmvtqYySu7HyDdGJfeZ
ymCCVrGiKxaealmI7jsHcz8tOdzNjG81RGU1J8DrKujtY2qQgr6nVDqzOSf37Ass
mlitWnIfkuAEet9zFbtQn6oK1f5OutfxWec8vTMIAHfwJRBhgKVXYRnNwEzGno2V
bb4ZrBVzEc4O8rCtaSmLFJmgohjHPrGYIQ7QphorcUDZn/KYHf7c0NW4TQMGtmNx
CG4nIgIA336Wx3nzsgK8l/AovuaiKF4IMdLOzpStI1sokDyV5SDezfBD3U1vQ/eJ
69K/6YOkMkrhOo6F+QNBqzRhLi+OKxf4rPllIsPwjky6Y88uJQf2zOFxIVM/vQXI
BsQzLfbSV7nWqwpZrThJqdEzq1uGmxhmr7BTgpGyXLytYWaiACEgrn5fOpWV1P4C
dN8fnQN8l+i/nOJ7GIpCGtiHObg/tAuEkqpYtz+g91EEdC6k/a2RRlpgdbJloYlR
RgFKBpfEXIrnB0ln3zZ2YrijesuXJH9toeM+WZ9WwHQODlLo++g8EA8tWBcb6D+k
tkdOYBF+P7h3PFjTGoHS6V0xgweWJ7daiwHqTCxPOQ4hj8z/r1b7KTzakg2z70ZY
7sRNAcwlvTwX2U9zTJ0I4W7MQWLpmnqj3dTExhfUVoqr86sb6S6OcipJUbnnr70b
qe4//P0fUDzzTA7cFU8pMjUIgRKMhxPjQmn6kZgloF0NxNRNADLtEcYlUNMr+ZY8
4axpKMjD/g9PCZ9kD8h04xxLKXx2wzzyraE05P1gxBRx72oEgxcz4xxhtvdsooh9
UwzjYMnfZcvVGba+2Hpk+5ww7f4O8GWRTlUftdXWpzpEN3o0j/kxNmEhqmOzxnkx
Cx/Wa44GgCduqKinQiZZS0hE/cho2zZh14RS9GMRRdWrl6pel19ZtF3w48gH7oZ+
pfq8w/8bqs6qjvnZJeYS4nEX4msx0dPw+7gHcjigL+rLyE60FaR3rabUO4z+s9T7
+rHkglAmMo5ZBee8c1Ss3MYBFnd5k9FCHL5LpS3wyn6HUs7g0X1xlXtcA66nWb24
1qGA7Xtc7wPfYHd5sAUU19EZuJGk/iQelgXpMnVyUhY45TwdNY4ljPGZ5v3O0e4D
uWTHgi5ehurwy5Kev/X22BcizUxcF/eCj1WJ/ZbSzDUh/Vaa7j1UgT7NMmrbSWqb
do/Wa1wUyFGWOvzzjur5W9tmYMzw65/UDqRsOhPpxcyRcE7bKluqcPSSC2JR4p3m
t96ualljByygDEGYJ0eQCV/1Dmu46V0bY4ZMuUbzyOxskSIc+KcdwBi1CSKXGsMq
ItJkW8mAKirSl1fVRuwMynXEhb9jFZowAVhUJoBIoxS5+4QtQIk3LEwiuHKXnQJx
3Np+wNwse6t+xUxgeuxCl4FVrNVcTFaAy4Dh0QBgrW3OONMolfVPJCo8zVcb+ODp
5w3c9EL5cAoqHXQa+YldmHE+MIF6YbfdMwN5RtYRVkTs288Cr2vIoP0oBoyhGpEp
5Ma9DNxsX6ZmKwuX76J/U6KLEnwm8bcJR3BkEBWTc3BgHTs2PHQFy/dBw4kJGr/k
ItolaHkh32dP9Lt4Uk+r3USbpiFcNgLKAhzWCyi7Ll19UWVsyhkcH1VstGeG5An0
dJKaN9tP3tLl/POuXml9eKMUEypbt8stD8GJLbyA8+JPEBecfMTohYbZLlmNKmHO
j0aK+lNn1BFBc+dQVssIOl8nwi8jqZJScBC+Fqn4jQRuoBX1YQZ2iIwqmOQ1OvDj
PKlRGrWIu7pPEZ4pYfNbRdBY9dxdrJe1mczxjtaqG1Sq1WroeLd5Q5OWPisEFRsf
N0U7+bWqfiJniwW5YpiUP/IvFEOIvFPyC9HXHYKCTs6oFtTNAq/0VeZdrW2x4JxG
4+8MgHimN24FsIecz3bcKA1Gg8rhHnLewWrrKC6/8tQF4jkXZYQbVAprFg+lnk80
NyYxEIZAh0YbWhzarSH+Ffb9vzjIGV8p+9S5V63VvlhMPXFo0C94yjpqwJD+G8U6
KxaAgBe6vuB0hTP1K3w3EVza7dju+fcbUuhp84Rxr7qOJqGE4/d9P6hVyNUl2cvc
A62abF20+OL92BdBRz5SKgq3yUx+rNs2RGDyAfIxrrNaAkXezKRcyAnKWx220ts4
rNgBbXP/UADcaclyIvBYDB1x7XOZUlWPyPWFxZQ9fUJCO2lRB2GXhnhOD5z3by0a
+Zo+NJmHbZih//RSu3zaTHORexULsfOXoq6crsh99wTPSI2k3LHcd61+uENqsQbq
8UrV+tdbU5UHpq3TI2K72xW8EV9vP1S5hxOYmlBKynm1IoQlLV3rCy7VG1Nf/omt
AG9jI+AgMAjq4LmCdIS8PePJffiWROpRL7EMprJGyFilWyPnocfLUIc36dQaPZhK
y/NFmYym/9iMKCuH7K8Jt4rHRwQnD2KA1a/cRCpuG27mEmbLgcEsyTtsJvkECsa1
BPZF0lVenZKLtm5tJ7wov0zn2eFOittwYDe55aaCvjJUQ6eZ+wOKf24ISqPv7y16
VI2Dld+7lUH6PM2CMHjxvi6xoU4HFdDdz8Qc11XOm4prWH0iDbBZD/ukuSfZJx7H
44oDejvQ/VgnrJM/1X/GqVduy5GVk+M7Kq3ing5zENjP+fEC05j/MI+87/RHjW6o
Uhpk2Q7PnOs8jNJpd44VHSv0i/S7UlLRwvpa3MOTdkchL0cNN6wlnKfW8h8gzwL2
MooE0nstgobbS54Uz0gkFcbrM6TQGogPFxhTNpCKX1UOhdfeo4L9573wbQlYnJCc
IU89A3Cact91OnwkU8kRAIgQNT5ZDhtKeRCRPPBCk8S8a/h22/cfWpDFVvTRFWsk
vs1WXUdDMDSskfOc0PDpD/fW7cC4f2RbtY2ZHJkKO9kLU9hydNauA7MUnXuRKMdg
F1V26r/iSx08Z2vyH6WgfqMZhgoYgOYKo+sNnKYtLXJO8YSCZuI6+bNEbgsxWKk5
CtQ69BaQh72epCyBpLml21rBAm6tGjiV9GD/wbvbSdAZ9nmskCuvZn4cFj4IzNH4
8R4XmVUrz3/Vh6i0u+1RffjEG0JH5w1SYOP7Kx1jdGosOzqPOm0LqA+1GPmKzRMI
34CUwrfkkuYclrPlkCePYDNvf0RcoohdMusAhf7fu+67qkWWLA1HGSrOBN+ahL+p
8PFQ77H3faTijTmYtVhUSJGkLMl80qPXMVzK4ILLLzK+1cYAtrAOsQPmsSm2/led
U19hkggu+F3yTaIB1a9LQkrRz74j0Arnd92uW5Zl3H5tbFWZMpjvr66w7kudtLSs
LheBMoTlmbPPGMuCeJUGRkH8EfetQTZF0bq6edgmO3nFYZBtxbu4gqG5/dWawhMa
FQlyx4UrL/QbF8Nob7VZ3o3rYskWKKAGVmDau/bdiv15/NX9ODA+GXTdJzGswhcE
8LXVjCiCQw+kehhKsZ27ppyccUi7DD55jtZTvLnV9fDCuFdqWsBPFJ3S8rNexB+m
XwXg3wfqVpL6jTEujKEkEI27GTc796Ho1OcarRV4YeQhS91Z9wsEFTV58CvhjIZ7
O1RIkhkctDCO2lx5uSP+w1hFZNg9tNGAQHX/pzcPtS9UI3RZ+PS9hGNfrw2yGVBd
l4Md0wJ87wwjwG2TJ/BHL4g4pMHZtMgJF7cX7zfpeUIsm3PjP87iIB8tlj+NA3xr
WOCeZkutEDBplyEkWOE5T8Ssi+ehymceWP+4qi5aUAXQjmvey6bqyP9VyVCu76DW
YmMHZjKNTksiRBPsjLh9+aKpUGtO+BEC1wI3+MG3B1wvMpmf9ICrxtyS3UujHDaJ
YOEuU6TGUIeizIBxbYs+R8hKJu0XjnrWxI4zxR9As6creZYe2x5qOHEGgktssXcP
xF7ay1maR4mApZpaGKRbTMcXtszdQn8hzcUAR2pk5+QZcqG1SO+pqOW7HnFel2Pw
cL6N86txg1FesNtJAQ7oXmn+1Kp4795RGld7rS7MzJY6m0Mh5uH63qeiFOIVNZWS
kXU61U28H6D7+F5wOWw/MgMUIapsIipcnZVTtXxT8ca75rADx+xDtokrF04jmsTO
cvQ5NL+v2OAM2JOgHugVn6G3K2Fe0oubJjhMWwJ1U1dmO4+QIoblANpkx1unONtN
rgRZ689VX9H1DY6ZhhY+XDZ8FZtBDBQA5dH8TSN6TOY1B1bbuYG6CJf3VyfHX3fM
P5A0weFlbV5GC+uFMYW9PUwJlJ6Zfghkj0XL1yc0deiqUxP3EjNrnzoMToxq6zFl
czaNIpaXlQ43I18VW+cIH0V7LiOzGEFCkErMdbfy96x8PSIsHoUJ5nG2kmohiSEl
YvbTE0F/yWQ7Gzp/m0f40iLGuaqJ+QtKRDeOiQTGGngvh8K5fzY1YoyU0p5Zhs2E
kO1A7iNSjimcuYg1ZVGVa6CzwqqpXz7GrdPXV1NWg7vrkXaxUDefG4DOrHNAM6UJ
hd691dPS7zBHrvsR+PDokpSBd/hWqPh2u14vrsVsh2OMHMP8pcmysR5v+/+pXXlG
Umj0lD6tbgR7sV0i41Tud/44s4erj5hOhtaE2cE/65ZFIyvcosPfZXJE6ZpQeU6s
ZKU5eL4Yq2eDDuNNP0Qz4T4mJAi/N+bFJbcLmFtbS/Z3otFXOFTKlpjpEB+h2idj
aYyQZ+562kNFVth+kalExMxtwmVxp2JPnSm/wUkkc9VnG0jsv563vAjMbl9RDVYC
j+yn9QETxS3Dg4OJaI1X+0z4yFUFYVR730CIoAs7CWqhKzPv1sErR7OExTRznW8N
6agKzrdNpW9++HnETOu+LUecMIqsBQByQK1OOkfiH4Tw1JPeu0Crre5t6iGf666Z
t8zrmDOGiWkSTvclswMEdQ6tR3mcvVUYj13ZRtJNn6k=
`protect END_PROTECTED
