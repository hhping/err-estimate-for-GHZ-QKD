`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1nGnacO3k/Q2kHSukr7pS1TlFUKKX+UR+8RpyuEcoA03taxxMNG/hoibJaMFYqP3
upkaOE4yQNuRmdZerJlnPmZQn8XxUsTjI0LO4uZkxF9WLt9pMQEImTXW3wnZJ5t3
XE4rYEu9WpDNg+9cRrTxzQKoFzPA0LeHgjd5qfbOTwbc7QXqzTNsbrA6KYscNWGd
PIpzLPVTvBJWbtt1VZSAQDgjLMksnLAxi2gKrdUbsj7p6KiJCMZttn3OpiUThg/z
AaQCL9cnn3nRB//Qv4oSYePwPiQ7wcPToGl20No85h35hnLB3kVS2yCbgdM2Klv5
gDfnbpuq+B64xTbnog/Iz+dTdXeC8RsunYFY1gaSDTb5Vorg/eQciaFH2NEnWsmV
8BT/AuswHVAJz/FONJ5t8Fa0RRqFopYGBNeFQa0PlF9QwOD8tqm5T3EAE6bPuYT9
DL+aB4HGs53mfAhmRM8PJfyd8xFHDQHasCUtsBdhRlZ9jbfbhQG7HsFgWTN7OZlb
lw6f5w4xk0RAd5W2qf1Yc9QRXUj0LRE7in27n/8t3PJJLXVczFr5CPJR5PgvaLHx
nSD+C9dw7cvTFQKdaUccVlGtMDFuJaTPZr/WuHzqu37PxuPPoQKN1kiTpkyrj6Vr
du90Jcn+5kFUu9V+DsRG0H3nnA/+TVGVIY0bvTxCKyULOt2bto/mTmTUjdZcudeR
wL8I64HDPU8hvQdZQ2RzXjf0O/aGR3iWDCeqyQw+Wuk3JU2u1JKLQpwlzNMf0/nR
OlxB/BZQOKFkfgFR1dNtUPDvHUg87zT3QGTL1WSm2kvtrjw7zqkK91/O2k/0dtpt
GqrVtNm6hPtUw5SC14rPxQ0n9/HE1FiiRP26Pe4X5QYE48RaX8yrrXfjxwW5hZ8Y
GRrhKzOBVEJ4c19lPMp76l7vgW8jxtmY47OZzrDwl+aMjZ57+FDjIOrdvRdIhYUr
WKOhHVaDE/bc40fdxKoZJ0b9wdhc3RbAp3+ZsZWg3Pv5k7ZGXaJOZ5U3968diRpq
II03Del3VrAr4tfl93/xNA==
`protect END_PROTECTED
