`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ffHRBBx7vNxlvb7ux8Xc42/rinZ4EAuiC8JIAxg535DETj3Bh5HRHUQAUTvrtdQX
oc7STNti/5w9sfHRlVo2qud0TNEfhNcbvz35NNk2sBptnr6KN42DjeV9LeJKgcPy
Ryuw1PCbLFXXFc8SgD25xi/jfVlNPc14DHoHLOX5yDcr+6PHC7ojhnUk1Q/X5quK
elPJkJAtiv6UEWJLjeeqOCnbSs4ejKtjQrjESFuqGLCRFzr/1swhaUfGX51WFa4p
8T9WTKZJ5LwsUXo4foeE8c5c/gVaeWH+J1PVlyKeCxVSv3sIp7IAPONAO8BuuV6l
YzTzbkbjo8otnDr0LDKd8CNT3dv4pfVL4TyaKN6bf4aqQDdYrWGo60J9QPHDx0Yq
2hTC2S7Mem0L2AcTNHRktjfv1f+ABMAzpVr4nLxvcz8q3uXltAW6pGto2vRRxVtg
`protect END_PROTECTED
