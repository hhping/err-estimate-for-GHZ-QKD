`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
75LGKAlOK5jhuPaMvmqhUgRg0PGRJdPidlm5JuXYLpdO3Gtso+5sxvqbtOuReqh+
O3SzvotmvfIcW4jkKexOhQmsNkPB9mridW32idftY5GDVwTY0Yv7EjHm1zWyecWv
KLuzpOKjY7BaAliSX+gNl4WJd9Lat1GkAQQPzXSpot/3vgdObZW7N4AfbjNRNwsM
s/5NWI/0eK51HhAlbNd9Z2IDX070jhHHmEbbXqW8CNapjXrQ+SLKtFu7zVWd/PAS
VYGBudGBQWsZ1RsWvyNrZVr2tBcKnue5u60uekcHk+c9pnZAJyDJAmBumiiBI+RT
0RPK8vsQ9CQ3qMYW4x7vWyPWt2wiCsJA2d+gJugsuLMFS+UkKFWVJ/Ws/cgFhTFP
ZEkHpqRuMNHyhebigPLGbqSM5EOQLnwL8ZMYeU8rJkpDUIGhID96uJyhHxGzVUPo
KBcsngjtCCL8maKLEzkZRTf9e0JRpNhprBNiRQk6aF9mcIAbq7AL5ZQtB12FpLC1
4ST62t6TqoI0SXeF0vNFoovKkRaxkkVObEruPwGFlTKfZK2F3VZzxrBDjgkBPLTz
rnzftBMEkNHFqWnZqeaO+pHjMbipHxTKJhDTZWdnfRfEWDyx1jgyKCk+4yaQgSOi
LdxjKaOcydy/rpzKZ2xR86Gwa3TTe6Mlrphh9oiK4ZugLuZOQpHEBvXOZ0+hCF7h
m+9yjV3SWTkfzMfHes7NomqMwWu03xv41UFODf/fbwX4hDirg+ANUtY6gEBQBDUa
/NlZyLiVKs1edArYgaFvYVJ04tRkOoX6sO6YXX1ufGo=
`protect END_PROTECTED
