`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fVoeVrM+MQx1PsM8k8Nk9rT9lyqUaKj59QiXPlAdkTBlmnTfSl0DTZ5VZfUU+auN
ybkooUPJ2FN33+LrwjZn65Kupsbq0zoAXWBIfaL1hnNqYtsl4rnawy4qK8tq4j2r
a41ozKWmk8vW7ubbfHpr8VRGx0XLD4sJmRu2sws99CSVdCnNVA022K0QZk5cqtM1
KVWFyCOB9nm3RdrcY/6txYfQrdttZj2AFceX96M3SPmiuWtfgw9456wLWdCxf6sA
VQm6HeckMGAWLqqXvtsHhX9v7NJbci/1GzW+reSKZFA28aZ6v5hKkCmGJUNCAfbO
U+ivGQ0T9Nqt/L0WVpAzx8pg7leQXDLLkJgsGES3MgJ22SQwdI/kROuXAjTNnPA5
lmWOYeFibzL+3lGYADBrdMNVLmFVsPM9s/doIRlS1M4uf+RLBS43eMwSE3E82+eQ
SKhyDdVMm9pEtOmN8mnyaZh873lz2Ppqcr9xnrzql7OSLuzUbGbAy/YEAz/3sgOO
VHr16E349d4s822uTmhUl30utfNn02Pwp4JnqCWelHTS/4Y42NrGdkTS9TBZM+s6
2cbxnpa9jKl2uq2BePbpbkNiPBvVwWQ2GWoPue3DNsstcCH9piXfhTcZk0yUoLCb
4suwDkpBSVsYO/HcQeipayKw+aTlmqXUCQN+q28vg6+4Otvu+lxRIv/Kkr50r9WD
w6l+8HMVADxbYjX3od3sp4zOtdZB5/7cHx6UHU2JhdR1T+eQ1Ahn5mEyDFZDl7YB
8nOum5VL9TVfebhLZJmQvhm9xsudWdF/ry89GqfC7w42OhNHXXuTdB2a7qzYgWT1
hcaNFjGNmgyerfwOQDiR0LWKaK5oez2jfJcvQFuDQgaWTHwJvH5ryWKHmS+1DQIk
TtWvTU9dJUxW98nvgGtkJVhs5NMb6znSEYBdvNQMUwdPSDJXnCeeQ63qvwUInbzx
XRXbnE2KAratHecQbTijPmOl9lwWVCauqdb2wdrNNHordXtajil8xfG9XXOJiODq
iZ5AimF/sXcqJLMBluabjAj9pDnNt/DnuY9dfieO4ZXQiFokoJ33HJG9ORzDRhqw
4FDs1EAiAiDgSjJ3wpd9gaFwvqxuaAnw6Cy0fIHD7ul0qjB5C55twpioY9SFFRNK
Xnh+p37jYTUCdPTIe5BUQ0BlSf51y32PkJqnjOiVS3wF7/K5yFMUByYpIluaNDMA
IopXDS7ClQYtzCv7b9fYh02SNxncevbvZDeGkfl2MV/TFCWo1g2bbPKjDr7HKMXS
iI8wujfbrD8RnHD+0rFxwZGYiOmVeZ3EBaUs8PLdRwhiRpwkjKJB9LUnCoDYnP3O
hcfWk1RFakqxF+V7vHCm4cA9oQAPYeCRpVid+CnfTmXDuHlHWxuT/ZrM1pFihMeT
KyyjchgEIMxBGk933CzadoEl4yDv4xExFzpzWaJpzx9e5zKXmN2h/dQfss2lUxPA
6LafZdD0rWjyKCCVE4v7KhIisVeKLB+Kq/hE/PoqN25Fd3TqCZ0JN2wAAS2uOtog
i+r9SUCffuovLSSSQUC9X6Uv2aMIYLVkqF8n96pglnJ956n16Eh2GiVx76XkmOs2
J3xuFr6zUZXstu8PCsSD6Xf51/AbStMO2+IadWnhRgYUnhaGL/50wEyWtTwX0zuU
YZ5wRe5AMGCGUyMU3qIRE5rI1dQhTL0J2EMVjSVSs6SgiVvHFuBelLkwlakyC9Zr
F09bCTJ2GGYrjWRpY1c7u6Puq3MmwZ3JaQwiGxDXSWt9DIb+/I25RfJ/RwivfYcS
Qh8kBdkB/bHI86rQgX6qY0tqyYRCDVVdbv0tJBn4r4MOsuoWMzUm88iaFLEWwpmB
9T6xMnKYmaF8K0qKgtm6xnCJER3Kca/DkbA/VOmeW96xsXiuFY4sK4ynGqajg4pJ
pPwhDIC7Aas0gILm4WNakIAcjRyVjjbrjA0c8uPkeFBS7oF0gD4yqe03+lcaZA4c
wk13vrUo36A9pjeU0amVqjMU0huKvHQazDSGeEDShRiarWlsmxHSaapADd5JKg6B
GeleBQRcUL/eUcOrPeb3/wkIXCuL0u+kAs3qjmL91S6OflWZaHLZ3LGl/JcoK1pf
tEGId736DYySxpyxaPxPp5k99oqkC3azykM+0521zJPCWH2oxxXQeBi6oZ2y2x5v
ysXqz1+SG7qiryp8LMTtF8Z1tc9EnHQovee0WKK2ptLNVqEyVdUVJiZwbN9ggy7W
4qnh9y1vrw42cfm2saO139P5y9rhmGrGlOGg1kWWpfP3M2Uah1dKwV8S9VOpODjJ
co8RK9VoC9w0Q4awn72cqX1cF6wywPEMYPYLBOGsdQOSXAs2pKatdP0zHWkao42Y
C/5PJLF2fAqCKE+lzM6B0mpVwHuSLwNDcvuYg0AmMBiqWWFsa0Zr66gxzQIEkfD6
1JaDkch5To6/PDkJ/BbD1p/I+C9hREMH94kc3oYZtfAkRrCcHSsrQRCV0EhIZ1xx
O/h60MUw5XWXvohTFAeNyE66nVEoDnRKTEroaT9DfY+Nq9LioY3wOQrHGrCMO8s7
eBz3vVKGvWiAGWUlPYrifSkCsRLQbJ6Qz1c8OqUDWPNpnI145Y2wTPeEyELQ3IRj
GtwBDMk8TRPSn4lG/gV+G/WSSdw+F6psS3lARgeGoIhr+1i48+OS5EnUjJTgHdKn
J2d/OtUhTVVK9yO28VPYaJXmOWf5wK11akJZ2KgBECcY7XGCDmOIgiCu2MJiUqzm
+0comV/A0z9edQMuna11gxhttdgpugSF/O7MCX+zbV6HiEFR8LlJki3YPX8b39cc
RLH0qy86UZPEcAMXbI40H4PfpywdSlyAhl/ySeaC1JvK4p+IgpLNzAhEZW9OrrBG
YbzC6fUAqH6DbxGn+S+qWWDWtRt3ITShN1/9KBRQ586gJtmyhOKBkR1Ycfk/Mos5
jKUDOBxf8OSMAtu+hxMyZC/UHgoSWJXQ79YBI0SvMJilZi2a25YOvy1zFBMkwIkm
aOuFCMwGV980TkK4LZcwTa6+jL8Xn8KdPqBvuHSu3SqYdmrfE8ID2CCfgBSfkyaP
C8zEdmTF96RdCEdRkg0wWIse/OzZ21O2wb3x18l2Rd6AnRjmnYpkXO+mYl93CJ+G
PDtJ57G0bnq4KyPlNC4ExP6vOWcWTWEMohWHHoOWuMbmAg+XKc9TwLRCICgIjj2+
NuKSEl5lfTUJ9RLIedFdH2JbeiXFMDEw2x/Qac5hqRwIWD/HgNkOJVUMNn3vXoCD
OB6fFVtTQXvRilHvf065dWATOBjbwEj2jVK2mR4NM3woK+gpwJYgUHoa8+4ohSqR
3zCOzPPeEMynwRYxvA0ZD5UXDI2aJPc4zNVk9UZgSlWoMpXsX6ZEpkkTP0y3aQXM
IFtTpXQjWROfh/V6+Hpyz1To+4LXAMiuhgkmMMKejk8K7USPhW5zz0APvgHfzSzu
H+y0rjTWXLHyheOVjAw80WoyTLIoRUWxH83UXxYIyJXmJdR89M0tgb+rM/EuDMPs
jPn7iFp8mlfjvbBBpkcXMO0fwBZssYapgp/KmP6cmJUZfv5af0Aza9aNDbwdtOYj
Hr3O3Pb6JbTHWG2MlwgbzUwPswZXvWIb9n438yoRHrwf3TaewxAnw1Gpbqr0ojAn
BiHpsqFc+nEzUunYl/RcthekxMyqvqrcJ7lajR5GkrGyKmbDF09g/sIReZbOnkkm
JuQmakEt/F2r2SwlCeNp66VCn9lcwoZ1Czqa1pbobC3KCDGuLneBaypL5cHpMmVS
WYvKDIfGv0KC84j34FV0ouAZM6EBKwtMk/ktLbicziKUCnDKMvoDb0H+XDc1oHWK
P1jvpW96amiO5dTecCXpwxZ0fMOdOhzX8jjRYMUK2XdDQiAckWRyPWWkrvjHM9pn
oOxC6JbnRFUBfUGEHMLtR+yAi+leec5iPMRFh/Bf+uD+WYURpckq4ECbtluNPAiw
Fhrw89VgTrxnmHtqVayi3J0k4TVTIu6kImKlM1GpmwbPKHwrwiucM3iuKSyM/CHu
I7d06uvpIcmQ8RtfQZoAvLOn4khvV5MQLA1Ti9E6QiUT2Qtyy4sLRfLIkhpBM6cn
yD1Qb7C5HLwM3dXvWAjwHFnb++qw8fd0DZD1nN4JpIPvq4kicYsyNDi7D28Gh+y0
yuXbF8LNdy7OyBv582V+mIx1bH7PHSWk9ENir5FRyyVuiDi51mCpQ0Z0cE3HpOvJ
ICP03dZ83K2UYGPbwCDamdtcVHYTroXjn2ffzcxoOG1arAAi1LvpXBrhLlIRyF+W
pl+8NKkbzbMbPpiqPScxWPXa3TpbGLuYRfdTzgnFmRZMyT+cogE5x8cxiK5PfL2m
g+ICCkKeLL2O0cHLWqYiQpufOWgHpgLNJlF5jlw39SlZY9qdaK30CHl8DxaGUEHC
AKob9cvwDZdJ8QJNLOTgU+u2VM9TJHSEHjAKRMPoQh/Ms3BWtZgcUgTk3W0K2/Ks
Cm1VQojm3q+kynruKaQ74ZXP6uGtz8E2fwE15PedxqDlY7iSgZmI6TPqyNPbsRuX
qVTJKBOHU83NUUkuQ3IbxHfbXw+fym7PDpZQytIgmlKyc4D2x1Eg2wSwMw/cLiGQ
u8KiGH94IAS45fMx7tQdv2f4taa7vpPhgrZtCVhEufumU+pqEYF/MV3bSGhWj2/t
pz9Y4kmnj1aHYVU1ULrAcjtvEXtQ+WU76Aa7ssT+eWIWckWQT7AoqYO4S5QPUUdJ
rDocAVqKdDEtx7WeFQV3y5PUZrKWu7TlMpL19xxNv4ga/1vWZGHqilfmwH4S10Z2
nvPDgoor1GamVu4dsk/UzNcogVes5OZ/oWl4Jt7R/MNJdTo7+QN3ycgC0XV6Pubv
RomPv093MHekxICbMIp5Vcvh2glfhudJGULFxrStRemALjGUVM6DcfzlXCL216se
OkX4dXZddZWmGax0H5pcqx43259TA1tdQGbp3SLRmv0=
`protect END_PROTECTED
