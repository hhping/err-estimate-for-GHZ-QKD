`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x6/U1o5Th5MIgOaTx5H4i8RmRrvREiid0N3vR5KHPdUd9JXWmILzKAgQNALF6P9f
xC4YJlM+aXMf1mYVWw8B+HMpmVVAY2N6ZRf2+rwEYFIZkSMJrhbh1td71BgP2lAu
49gCJjQ8i8NNQNkdD6DuUG+nSHdbWoJL7y7KAVtHADmr0TzUkwC6l70xnU5y+4Vd
+bzhy4F5Hi5BC7CeFoE8FGKPVlWsPQBttpLj8wD9TM/c1alItybTJeAe8cLlELmW
Dl+/byskImJvtavRi6Oet4FxfZND4DyFGn5PpWPUm7lFAXfNdGPPdXc6PdEpUBmA
zp6xyasZOgw5P+oeuSPVtuaayJ/rhopTKy6YfJprB4V8Q5jYMDDGtORr3/gXJVUm
wV9sHukRs2H4tl94WVaM8yOZJqBcPK0rjvHlyjnqbvvQZOqaeTbb3DzJqQUDLXLm
Fxa6NOyImwbr+cf8ibuzrcxwC2en7saruKB5tcsZfKqlRs9PFUO1vr8MdC4z1he3
9YyE/en3AOH03KQvTXGvFHwlTdYg8i5SoAY9BZD5wVIsZ8q2Lt797ozOHeP3TtiU
4vBz5Zd8D4aVqoo/6xIIAdUKW2lbCKnS2aUIKNgREh2m9nikA/HuKTZlEN2tzC+5
M6Xshj18ZWKCasE7evFTYoUsZRNjKCgJWQXQ3c8w/JxbksjeeHdq6uRdR9qDzA6A
WsbCapcorPrV4sgwYJl2zdAZuxMxCAcMs7FLuotJpcM5R5AbDpH5kvo7hLOlPZ8t
6+3ch804g37/KN+FecG4WSBHXK+vIqGIGPuSj5VJi/GsG9satj4LWVjUalLTejlV
B/xvnCDDlpM7ErhaYC6ACMRH6pNiZ0rb10jotUe37v/r2UN5fj9UltC4V47Mr6zU
oODoHm3dgkbEdYVTIAQsZNxHDBpCV/rXO19qyhadUSRcf0yuo0GWu/KOWya+ikG+
7cfsDpSDD1ARWNaSF1ut7CrIYXtaAwziQwYDv0J4JhVs+Sp6kDc5Jpwe4icVJFaj
oh/pXe6IrTlbLrdgeLNPp7O9eHUKfio4s3VAM1emhfEGrsFZ+S99jkxpDTsKUXkz
7dcb8JtpboNuyQ6QmgIrX9td1TbLoUnIa2gzO1iphHVrK1oJOkWfdy5UbUer+jDO
54SnI9El53kU18YJ2mtNeFJb53L/fIdleqCi8Flz+L1I6953DuKyFN7AEI+S/mF3
iT7UnzEeyMbBcvjPvZvfpDcjejpiNqhOrdpHbPDnDBKrIt5AXRTZSrDIAWZ3E5dN
EE0RkSBwgLydytupTIqdHn78Cacnutwomt3KrVFMZZAOfANBrrEl8naLlv/vjfxF
TdDfyKuCgcEVvqIMul+bsi+JtnYy0pMLLfx4uwD+NpwX33LeLcU55mvgY2V4DZyf
H2w+ZahIOTzPqjfTU2fQ7nals4Oka0jsgW4oOkjmaKRELtMDz6liyB7znkPgQ57B
KK/3ktFjXumTOBHHEvPGRAU6UrF9Y4HWKs3Dp2bf7Vjr5e3/GZKrX9p6aSKmyYU8
bRzcpNUXBeHWWjGpZcO5+VR5E7/vrcjwrZKIFgl87BHZKbQ8pOOQbKGBxxDR/2Ud
A/a1wcy+WA0Ef+qeANIEjmxNHh3bfJOBe4GSwxmyeG5ABRXxpKVlopyCHPzVZ9+8
243fDpSY8HK9GC55KlfPcKeoul9rnrg7wuHlyFUA0M77q8ixfiVsTh9byCRN3LoB
aT/b04U78ry4oXW4gzne4s/jGaF6RB+s5Cs3rStpttuWYXEqu41Hlbws+mNIdfZV
dzlTYEY0GANSQ9jDVE2KHuMIIiz/C8xXpcNUQaka+lhdSEPFQVQHSh2laGO6gn6F
OwyYT2tydOvCoyt1yA0mDqFEMrtVSgx9bj063lrHbc6pz1dwZapVER78snvIa0GJ
Rf7lGX+/l1pyvl97ZPQfPhMG74uMnjjmjWaNyGuse+Ido9cxmFEaFg7myhEevy7l
V1ltL6D8K8oRzNusfK9Itu5bwfvbhdFsOdz/p5izrFLNXYHQaDXCd5dfmFDzRiJN
0nZnTgql0znyObtsiZF9fY6jvq4+tnoEX+Buip0j/avvO5gDwSYraPcrljM58i0a
5M5YzRYRdX3JJdOqVwoGhS8q0dRm2uR8aGNxmlD9KApd7TkejCcreqKS74CBImJD
HFpJCsTR7UUfqiDH3g/jfvStUoGQFlWReJABDtmrS03RyW3R0rxHvJNytYTpnPBL
sekUL8KA6tVVEeGOzAcRX5lb7bzdYNSAX21tqpXCWPGHDI8EI8ka/6K0XdfNxRN4
fD8Coa9R4m0mYlAGAMWI0g44S+QROLePm9quKcmVvfm3/FPsLFLVnV1yJp/Df0Z3
LWdcoQRJ477kv9yXkOlSt2hP4w0xvUwPCThQilz2bRS5nmm9y1iS7SQ46pVNa+u2
eIWL0DAPse0GNheBRYJnLSKOYBRQdAr9RmkbTKL2zpG9/PtpvjRtmJ/G4enfp/yT
Dx3oaTLeUyrcgDSXmtCCsTgrI5psQJjBDAcGSfD4eJ5cgRye8Nz3Vrb2G48GeGze
gJ3+cIpbFycSQqx6f3Qa6u69fIlBwA4ONHEiSNnC6StvcVXtxyrHl7IrBruu/GEW
kZVwotG7AS3tijrUYeEhAzxIuyG0B+fQ62rCY+dPZfpc3lc6auDLGP9qfFNphQwF
UOluhyc2z8MY3xNEz6/GRDWtLNsngHO2D4NhxzJTIA6SzufQo0nTaMIMT034uiFM
lK64x5sAI4DsKZYmPm6QqacfcGO/Rht0/ZS6YyJ1w4t+X748Q33VvhA+UJkDFI4X
Do5P6QbWdg7DsjP7eqMqI7qZpHfs6OA2LIO5xP1jRbu+4Fd0XhWxcK8WUYUZnfPt
W7KQl+gvmLkP9IIyproEGUeB2PAK3NNq3kPVcxDnM3p6wnuNJa+7jPTl1Ij4Q8G2
tucNyn+GFnc2C2+sSdUhL3eqemm9ygeqdi8XroBljBuit9BVwqVzatD2NDiYiXWK
c7s1eUaC1KZKUBFpwl/b0L4zLnCDc2xuSt4cHm1vpIpfQ4ycrGdeP0pVswMzuFNS
2UOgvn3v6qVgjLDITkY/XD6AqQPbT0WAYkqzU2xEoTlApSHaC09kfOBjPFG1fIZq
9zbaU/BghlLGkTaQcXxPegwTZ9A03fx+bIzGfI5M+YYt4SjvMqfaPUs91EmAWU07
AXPF4zQs1u5/s5a/s45xbo3qwSAowOaRZNaJhASVsooHx2YxPtVgOg7lgasflAS8
/LqbvKAjAcgo39J+8XZHPTHS9a9xGqz0+MPP5LUA+N1ZS6wYNX/moCEdRTig9Ylo
CVazcKSFnnUrXpKIjYRSUO0xo0VtAL8cagZ8kSrcG2jOpTJQoxEw8TuUyR2aD6ci
3RFtf/r4NoH/LDIPOqQAEgwjwyTr6XiOoWapypJbwzMXm2Fdp6dNFyGN33Rqh2NN
NC8PKSkXGfOWUE5hURUd/NKB+8JwzZhVNyFGO9mkm+Hw93jGbkLzfA2leVEqphjd
yBfPuBHd1wnU+0gCx5W5ThgPwCOH+2wny53+dE5f0HGTAuUqmPfvOJlbwC/R/UKX
TgBQg7K3t20mnXjDEPAaZwXdAQDY98PvJqAT3TztuYzLSWSMxqrjT+bugWfubpVH
a69JJFBEX0vcPPAhrjpSoF29oW1rYmkXhfkATs4HJy1HTflJo8HwzjChVB5YIcBT
JTZwiRLdDvdvwLpeJh005qPiKb7KSF2/VEK+PkYEuK5p85X1sHKe3KqMknNUxGv6
+W0rl7YGnB2k5GESt0Mvx74hawsaYWX2cQgd1zGVq1diIgwTjEWzce8GQLG98/Fx
hqBiySTLle7cebBDQXN3jLxOAwIBPePBOMHQ2oqsPe/RNwRAJfrlYNyyJA5uAru8
AnkBuHd5DzgE4E5nFKEK/xmA2ELt/O7e6di7cBcDhdl1RpRHtu5n1/YWWLXMbw1Z
9Zsu6Wce6hgLZPxw82dcpB6CmiLhUGD4L/xzVn2WQTcAygihfO/OHcJoGO7ob0uT
EoIGMW9+z9Q4we5WB8jDa0QUz7lzaUaX0n3y2DB22LAezNq4J4HwGTphO/d27DpN
kOJY9gHNaiv0ScvYqEkeLysxpiH7HEfJJtD6AocCNtFc7bzZPg55Jkb0MLGhajo5
h4qWYg/w3OILTGlpBYjuLtz2a2ulBWzyhGsamimMAUpPtw/Ka5R5G+2yiK0IU44X
zb1dZnRME9IY+12kS4H4DaqH5R7T5iJ1t9EiRIMnv3AlP1puFbccg10O9ez00EDs
o3kQbU0uZjz6puVlaC7EKH2N/ApQSMUYPE97zFqUXXCCDRd1B/lkpad4aXl21pnH
gP+PtL6ev2XyhlO7sJLA4iKd/kefnDiClvZrALmkPTds4p0wg7LesGTDHl415GC3
KRrkT4a0DRioTJl0uUR7i6mB/KcNH/MCzhJD9J2NuQ2+VjOYOB9SgYUDvCAVCcgf
gE0XNzqq6KswZu8PI4gG60CIxMNMbRj2BGN4IL8/CIg75IyUcFOdsVKn/qOIBDiO
ae0aDg4HJ0rcSwzE5knLnJPHN5nm6Z1DzgRCXQQwKvlPqykyFm2I6Kp/EuHmJjz6
UAz02lSl8D8mMlWCC1VAYVGF3Xr2cRsCcxm+0i7/oglDeVGk2/+Zr/20I0edZ/gj
2DRa3C4It1xI1dnrMh2z4DOc/KrllN9BvmuD9P4IqOcAVFbFo34+dgG6pQmI/+yF
OqPwilNg27r5iKu+QeG9JRxbgUZQcaTGIAyS4o/mk1DbWSB8KZeDbQmAlmjJ0DU1
HWuJpvO/Z9ZCtNrCd4MlJfhg8oSFg389UQn3za0E20SOUTm04cD8gxDTKSos1XrZ
NkEH6b60ke/DX3kREpMqewG2+ihG6kvkLYmC3HgrV73OiFtOU1kAa/Ql4Pznbz6j
QvfpMzcK+PibNupxvnHmGKQi96dvrXEw9zRjCxae3KJl6DKb7pkGm4pmVCI8WjGy
7vMW83lZe+CU2I8oFg5OpZ9ui0PKMLcTdkAbxqgrN1RXb+8+TrQfuXRG1jP6IV83
8pQI447IR6TS9e5xZoYzKxdxrB+8Yka7cxTlI/8a7qm/Mf7O12jVDLdD4SLDtFBm
HKhe+CD1NTwyOJDVBdyLdY95ae8RwebuYTYRgq4g+DmRBcoNNB8mm3wAaBkXU4wk
XznOdyywIArCteOxUHKQHgEaoTReN0n/PS3hYo8E5odXqDhy9QIgSp5XFxzBkfXd
2ZipAfwam3c5R6ZA1AZQFFcxIcTBTLt49fau66V/jOFdGdRbQlso+5AEJCmAPAla
KMX2VKZu2f5dJ9+4Z2HKGTGbx1RfMTzAR+j5ozTl3t4fiGgiRxzk96+TX/WOtI8o
d7R+ED7qcM7qEBHkWTGnl+DgOKColcuHyTF/izg6S+ohTPPvvMfEp6M2rcZo+iYm
K16dbrSPInFrDDex0ncvrZGLXmRSkh2vkU4A4iqFM3195DFMuQuQIfug7wwqlqK2
puB3eYD2dRX/oGnsuME3+1jx0oLdWrxM5lW7eHdH59RjoryYc3svIqjqnZpKJUCa
hBxJUmjsb1o/WMKrDoXjFfOM1gA/xdvIq/WX4hGGiaJOO5z2BgByRBemrGkjRJBn
j1qKm76cSZr/6nejMwZDeKaKxLu126Yr/SRhnVil0w0n1sFmHF2dnqQsjrZYpU7U
bNcyPJZ8zFTGBNsD31Y56UvGAWqAjT3Y6KNPDiDfzWXHQAlOLuFcbz9xMk6jDWGA
fvn9ZI0wvt0264iBPci0KHBeBnB6U2iul5Bkg938/5B5g0oo9lqfDbRA/wcuhkFr
JdQ1Dcu2G0hsCtyWpDXJAprPNwLoiyG6mm9rrjDiydOAiF5HNjPOKMD+8G8jitgg
W9mjxp6RFz5qkhEj6FmlST3UMOZxlgT3+/6R4KIvXRny3ejXIX3sdkq+jtHGXVVS
3Eyql5V/Sy99UUoScyawhBLo0b8pue9otiB4F9NV7q8NIWI/ii5REjHRjyxNEgVe
VosXfRReC2Pxkg6T4mWqG7CbcTW9Pg8PY1IYs9uG43zoBpKHNeILy3nDo2ioF0K+
CLsQO2+vzrWUSuDmrjPVnX9zYP+4v/kR5bjuv8RhIfBj2ipofJYDz94lTcVf67G0
GOEJNj6s68UZ8CtdxajE2g4YT/3OTvID5wpguXtHPBlXv6IR5RrcxUQAIxrzEU+w
T9VIr8ymnq92VYQgFQPlPwEykOIDvmQ257vKVo5OFw3IBLZKSCzm2uicrUPaBquU
765jRuiiZBNxLxjyZX4i0oWC4gTpLWtcLNso/YoL2MQPXDT3a/wxl3TgBrdIIITE
p/FxLJB4cgI39uDxgyGGTHnbdYWbIyu/yq3/4S3Ir2cITt0eTbiHlW7qjqLKOBZb
MzOwdxIDOpV/w4J0/6t7nuArM33zqajQLSJdqfEFVWbQIwuFDgMeP/uvwSDw7OaE
I2/TbGog2Qy8hRRx0FJAleWhq+Kn5tnLOzoPP+Ox4vFF3tSzugRbK26J8J2QeonM
nVKCq+Zs8NgvDets5YdbmSfqs4raqCMHTVD0wnk0imLYxrXO1wUGovrjkc5+2/5E
8Lags6uY2bEUhDaCYNmkuGFfgVQ2Qry4gEy+bAA5Ug4y0ZT6Yhq1BJ33x35JhwlE
9UDHdjOgxnxsshG3fX6OT3nDUwPQjYIclyGSdG7O6Wg55OHppxEw6JalWfV6AwCi
duvrk3v/K40RJKoAtothd1TtSux9G/zLOacQEvseuc5VfapVBzYbrU7TRtZVj6di
bMC6e9b8hW2N0HDawDWQV1ha0DT7oeYuqRb15iYXxHTXz8LRwjYgvC9VEbFcubyQ
/S9yBIGUjhU86jWi9jY8Bo5SEN8EB2RUHuA4h2GmyQfmpVc4h/Uy5JJpLOVFSfyR
hUydfayYOxK4Jmzuu4Fm5LG6lS6i9CHzAH+Lslar6UeiGBg/Smd+pYdNbJ2S7n5p
hjy3pdtRM7ZyoxMXFa0FmTv5wZo0gELpmvgXPxBaUyIunnt5YNnPPHSY6UnUTUP/
yxnEq6N0exNkPu+t3k0Px8/n2zkJhY6qSDiVln3TKIRlgJKjtJeVFjapp7iGZif4
6jfPHss83fOXibydUZ8y5mubIO+doNrORBCtq0Vx9uve3hhUIy0UIORKTmkJL9Nn
z8/usrrFMV+e7nOaVTdFgb0AU98a8ZDt/tWj5v18AyLdcYJQmvvXc45WRGOqs0Hz
QbXGsqtmVQILFSZIxfw8E83h3dRAaiWgjtkZGyqlHenuIKNHsMG3oVipL9gK8AEv
t26FApD24qwBgbIJk6SpM8J+bjqBTPLvaZPrXcQOTgqj/JtFpAJr2Jcd2nlwer7g
+dqqby+y/A1+CLq0ncYIlMbrjKLwdZAorQfeF3EVIyDA8uFPTNTZ2thhTlVmXjB+
XdrrbiVIbK88hPFk7/04E2XBA7FHZc4w6CCOZcVxdBeSOKcR4tlHgFk4qBoSZNv8
h3BE/CP9LeRhHwonaPsAtehyagE5CvUDeFlpu1MBK4NfHV+WUdfhi+FMoe07pKSP
J090nfp39L5TWY4LumMArsXbcOkKJo4I8Xmkr9yQ8qc3rGRxnkIk0msAUuUx1JLv
Bu9U8UrJhtGpleTIrrxUpcoKpKfxxxKTmQ7QxI1wvVufNNrQW7PtXA+3hY5XTTxf
+xr5vMBRt8E1eIHNVS7yhdXwAMb67+q2SN6u79037zOMI34/jwGNQm1sO4B8G/4j
cQb0OWTv/zxe03YWUayCKnIEAJsA2Asa+LsyaxmJmMMSfBjnbD2LOi4fucG3MKRW
HnM4n6qC73x/ohR6fbyjoPAqjkQVrYI2AoidhlDFrggqHWaPezsu5MeLGfga+vSf
PXxMC07kYxXA2LjIjUCpR41ta2X7NttTeeoGkNO9jRy+OdXm3WO3gPzkj8jkbLCR
EeL/s9Xo1cjLeTpLRajgCnG1fOM3ymU72MJBAeJO0AZ/zJ9HsozeD0Leyq14WDnJ
rPb4AIW2afkMMn5cxYT8EYnceerU9bqTgI0y2h6LFhOjkmjoiZUpE6qhUV96zJDU
m/PSrTY7ajOrFuwaHjcCOh6WWLkPz76Jwphge+YtbbZyEFEVJSAws/wzmONS0ibz
cgZDqrQ+sWeNiM7J7VYGnELtHZdyOKlpOquIv1nn5I0hfheuW33Bj31s9f89NaKv
QalsgUatXMbXJiUgEJQR+UFFOWY3QfzIunRKYyIpU5dARJ7Ab/SuuCPcupO+kig5
L+PtYFNdRLTCKPQU2oQloq1McosSEtHpr2h+tc9i0F6uSkUHHfwbuSOdq+rda7to
ebccTxQGd+nTAPdjsGTT1uDjdsvAx/wXU2QR3QxQ6pe4xZlDOoN3gOgmrhubQ9jF
v5JR6bJhkSPvp1N4TtB3xGTo9YFAxUFiZ/MPzrqFTCDjxzGSPrAAFhe8gkMXA/eu
9F46Dgie0sY9iojCzLg6jfj0Hxa3NJnxT7j9fUGhwIt8fPavScD9lby+Y7dxmINu
3QWgaxw6l0Jal7UCQbDKBOmHuo42PA3KYwB1lsYX0VtJFt2kClRx/g81OmQ0s0pa
TpFh2bGXiam3qWBCyur9+qh7ByxaHi0Kh6jb4HrrGJ6IgS9jZTCZSe/rCxtf+Q4O
W7NeFYXPZ+IBWF938Mfux+m/Gapnzek2mZxbDKfDhlk0BE0J8TN4q8Rp8/PQFwTR
o4cQtwq4gwt2dHnwrvPlExxLHSlTptLfv0+KDKBMoLtC4xZ12HE2aKM06g/VIAU3
6Sjn6C7erwAWOqoJxcZWRer0lSnFg8SYdHUPZqOQwHx01j2VQNLQVFyoOZyURNGB
ZOt6X0n2xQeqX60Qcs8PtvCqkDwxACrwGhUbfmHo2zz4hlAzrucn8LMIDwEG4Bt6
IMbDp6f8Qam5mYJdph0e+16NjqsPbn/0/NYoB1P5iiVrii4PALLk0pnGDSc/QD/j
HaN7a8KjMwWNCYamHst+TOlMPnRKKjizbDpO+tEFSY2BCJd3WhbNTscatmIk+M6L
DpcjWcp5TP8V0zqHcbv+4v1H3SkyzNve2aT7HE3f+n3+2tsN+LZb4BCC/4eO98ZL
KAnoS3yvS033QN9r0WuCyY538w9QSypS6/1SvgtVlo5OiRLYaSkvdO9WJUW1MGkV
rKTvdLX7OmQgIZ5kBY9MIR05SKIxgg7PktezUm4Nw+MQsre7oNwXpOGqJZEz1Q7m
d6twa97KCZf8V4k83x+DquWyNC6sMis6J95vh63MSmwxq2kSBg6mZgHZeo7Bn6EP
8IUlrU1nRekb6rR7bVDZHj5aHpSg9WVjELTUTX/MB157yulB7GkRDm5DrZVBbcmZ
1cAU80mpTKskk6zRWlwTxKSR6ui1CxIs32VnOjlyjzRyLicGJqV89RX+MoOYr6YD
ryDp8X6ANn3lT1mPgEo+VQWYypbzOQgXrw963GYwy9JMlTFTx08dMwCh+9Cwypgd
VgLQ29CiirLYG1mJo1CDZJSI3orZ+yAuxMHFuxY6JUOpKuvucgFOec5btshI8YCX
HgO/XtiM6JJYAPUKF00zTkbGqedBsWhlExuvn5h7ilBKMIhCw5P4dRFDnr5Rs8UN
3cTSvY9zQeBHepTNuwqTDrMuH9xVpJSk7C76fLGkkXtreOE4KDVnDF0yz6aYM1GP
UChsI1+e+8U51iMH0lbhTyb15Ti3ZxQhPMjBXUDY9kO3ENX6CaY4njcO3l9+pU8+
nTYuPx+fmuHJ6tHpk4fAmrJ034fc29A0SPGh3zA/hXzP4BcDEoDZwnDJOkd9dJ1L
1HtsE4wsCEnz8BxkRSC7OPQdOAz+7Iz/drcwk5xx4KXoWddH0yTrGThSVKJkYvTH
kdJlBzb6ZN54pqZiQqt3lwrTMcqD9Ssu6UtaKu6jqyA0FQ4aHoPZegXGi36PD+Lk
pE+LJQTiExN6VitZZRKospIvOxhcRYT/WhBwtCIiFBu+wdWGaAcauiwB2NSHjmOM
YMalTTDh8a1mZhZBQsWmqZmqOFcmslGazOfGO7vexy3OQ54gKtt6oFWhIPQC3ksh
/H+mJndKn5L1DYkeP7Xa9frvkksLMIsLdDkk3OA7CSpK3jNbGc+4dZXHPVLr1nPM
i3wFL2SU6u5K4cO+RteAL+qu3lToroGtotyvs38JpbK48Rx9nFEaCx1oqjRl/NMZ
6Mc7AgVVwNLHxJ9QKpdcSG1TmV+hIPI7gKgNsaoPsUFx1m9wbQviFQhMUT1YME87
qCXVEOqOLyrMVIxvbj855BFulW4xkTmyuS+CXGasm5XTDKBhAvEiTWCWdj28sOT9
YQXHpy6f/Df26Tdmigts7AM1pYlv2t+DCD/3feQCwRlNLMWDsgWQbLb6/dJp3/10
wBUyZWfpR1LZjK+E5q3Wzw91l5/Szz9Y7xgsMWLkAzBitDWVC3it3c7+qq8v4xed
dg0xaQjNxRSKTVqHVX2MiVkqR6lBAQFJfMxLFAEwNl9MmXfw1CaP81QJPxa3v6Ob
+B6gwQD9mvgYvhUDirHWEzjkEQgXFinp946ocnV+V0Nc9rZglSo9l4ZrzKv7GSX4
fAaVSuVGlEW5RZ+JM9zCU8uk0+Cac9y4tDBXapMFjelbjJPO7lIRAf6NCAI55Uir
nGNEy+gPweBUNuxwEUoyIZMyc/9JQImJXu4FlWftdZAss1LZCFuXMoD9rhqTqbry
HZO4dNC0/sOmSxn/VTKNpS5WLSCovbqBZ1lW5fLlzMcA2uvLEHmBiHSZrFw1jl5m
q2afpKlCjI0YzltVCBh50jUyns/0Mgoc7p/DLd8wIeH+8Fq5WteVs9irnB0gShei
g2lJ282P0O+/QXMMUOc3rbRbvaTt/lKXlYUGLW7VWHcFSI2DaM2Gf0X2NUn/HFos
39oamQGFoGsefZ4e7YUnNAVRe2ip2DXU1XBrtb2Et7v2eKRnYOz5cTEN1A4aTnW6
zy6SM0OTc+4rEVW877j4GW7lkEJAeOAfvfTiqozkdn/97kVEmWusHDohjMW4wUsP
hkiLsWMeMZoNuGF/Ty3M7CepPxqzunhnbTdFCh4WullbvDAVfq27hiitFdlOJ64E
SuMyiYFoM3gOs/HpNYXhTrISvMNk95GL3F/9q/IsOWW3rVYV5hMTlJSXk7X7fCgZ
yNGOR8Mf9IfEJf34/G3cPKHoFfuvFnjMIIEVxZINLf2ZoGTTbq0pzKV80tw7I7kE
ru8NAXgY/2jBeIZ2B2OlBj3jT1I6z2Gr9n8sVk12wyXv2usiTL3LkqI3V52MTzuP
M7FtstaVEXrvAJjD83NBaotuW1k1yqg+d9et8QJJKK8rUBIRaBb3f8u/tuGPv3Yz
nr7u5iLDe0tIeNM1NgoKsAkvvP6hZKcI4cU58GhLc8Pp2ONEGe037DgYjutsyyDh
d1FdYtJS/2DHwtZOYGDpXRMLxoWC6z2OHzBojHNjtNg3uiGLGUc0efpwjzsQLvy3
yyD++TgIv5Laj4f8988DjJEcVdPd6WZWB+OL21q5PWXsOc/fZMWumZ1ODG7bepM5
IRebPaIJsbYqqV/2+qBgDvpHkZW1ckJQj7MPUVC2s6gtNVR3Rvn4tlPiZ+g2TdzS
PdpNpULLCU9f9ytun1NlPmXLG8UE5iR8MK9DuAPwE0k+F2I8b9MroOUzdlbNb6AR
wIU9zbz5PbS2gAbkI/X/DgL9+Kk56S1z573C7GLou76MznOiaUrfNQNXw9MOF5b2
KEDL2inTldXR0zEYwo6zlGYfG+W5cU3L/ziD4Li2w6KxdkHNjRmSjfxIA82k9mxS
Zgvyk4VacRbexELlGPze8Rj7CsVuPR9phBrVeE1/vTHRTYiliKLD1PN8kNpHD+W2
+qIZzyoui8stgkSIwilwHcH8mJXjsppoSSFp/KnuWuWrTXGkY72Fmf2IMl9I0k0/
+nStw2UMqK2TcFOqSjrRa10liys8frxvmIVLeFQfzQnnnseG1mjvn31/vvNNthJ4
gFrm6InkHtyEbWwCz2aYcUMl63Q1ng2kUMxCyBtY/wCQOpcB+cPLyOE/atYaY4Oj
+X5+siMsFphEkavqnpmkNadS0koaEW+yMi28kqSK6pWMvYupGb1qfHHsZgWLJYqW
P3Go4heJG6fPNaOq2XjO2tswA/1kkVQ6r5mrqCo38RCBx/IyGO9PY6+fTcu8cRkt
56POIzvKNDTmHIEwQmSOnCuQ3CwrsCWXvCVpWS8qwded4AurwXdfbd50+fO+qiYB
KxfWmpQW6PlUVaMxaIp09yu76pllJksyP6lDgzejX1x6vMqds/0pRKxrJ6Y+7xfA
Rtq++uHEi46CfWgsTBA0pyaQAdPcis/ggm6HnsAuHQISUsKYSshljO+xukomU2el
byc8wacn7ZjqR0SKeoBPIwhW03x3FIwulNa/kFH1fXDd0AHd+U8J7++mPzpZ42ol
2PZVnw8guizLfQ0ENDswWMX3Dy/zAHt2c4iE9VdhIpXvujtxHrFE+G27o04DFknh
jvT3D3GhY7N9mYWboxALPK9UAxJizelXFekYyrY6z4m8NL7LPUwdTqtlMJBluHwu
GQkguVsoiN95yoq2wrSpXZPzmntbFwrvJVSJFIJtASSktTrh3uB/kvOFcjOufEyJ
aB5XJYpO95ihVSsHx9Igg8NQpW6p3ekWIgB7G22RCAeqnDSxcsoYy1tB6W3gqldD
HQ9vEu6KsgHOjwoDsQScUC+AKFuy4FeZeuPfAnYVmuCJ8kiA8G7Bp3LNcDGaBdtf
4ipm7gW4S/NnAyHGMoBBkraVxArzgdn6X5xm1BWGVp098HEf1gA4EonNcj/Stl/C
x1SGKOdD7uJmMpp9BRlWjJ1Nr+wqdgWFHwbcbQB1FHFJE7JabA8VZUn8G9s3a6yv
QWzqhtsB9EH1AY/dR1U9AyggNLp6chMt0SrMXIDKZEq8XphVsULaZ3u9QkJj2GeB
nmqH8c7ms33NO/YDieKC8k72LuOswzGKHc5Uyq2NuMBgPVn3/gXn8QXN2zdWjd3Y
MrXmVot1PjO8VeTnOechzIwHymbxSizKHyNUXrCpHPDHMqPAN05C4Q0KG1AbxeMv
GrXEHy/vxc25WtZRi+18yNNQRMuU+nbEC881B1vHquHF913EnSbXPFpbc9Ish/rp
BDzK5c3rjFkhOPi2ErDGevZ9wtdvbg6hXrxlhOBHiLV4+13CdUo4+A7dACE3soph
ygV72lVjg6HN1YqY6keu54Ld5p0UAb095/3f+knlmJh5dERi22dHD8Y62fYn1EYT
CEjXNoN0wi70b0pXUDjvayvlUq64Boc9w9FqDkcglaq5rpB2usml0gTVwCEEjqgM
ndZdWJlaOfcOu3juW/HvllRfS7+hHiOwV1/SuNpJdZjgYKbcPUQDgFZvumXAtcRx
gNOen0LpjtEl2kGRWrMyWN9zDpsT239kTD5On/Kn//+/UMGPLJkaDxGN0DIwM5WJ
w5UACt+u1i9kPRsYhQIZ90rt74msGbVO0wgMuifzh42S5zXtikbP/s2uD3uPqvDi
CqsaDzWG3Px/lrqARU0VSyM+uDqrxP4s+h+3T/MjgeeSNzSrmM4ha7C+TGIzcMXD
y3vnnQwxqsYo96qtRuDk0DinPFAxWP+2fLpSDrOk0BHbiPkdQshXy5gEmZokohVb
W2tj6zRTEXqb4N71A2qz+l/LR227xfvZGNcuzotp4OXxTs4zTUyNk26ou1Fn0AOX
LumSVJmclcDoY+Mdsl/MtQEQBjnAsrA98laDfX0pGG4rmoShpq1oz6tP9F7pugER
84n8FAaQyfwPq9zdykKiL4Ko3Ay8Gb3JVq7u4YAanmsCGClhVSv6LuosF8Zqn2Zn
AMTgvfugQh4Gfx0+BV2v8xhRKtNF3sSotD3AwrzUbRaCQvIARC/IHKy26d2zlGqI
pjb2wpk6Z1XXgeNCTQzlJHnBnrtx12XWt/T6hvch+HbMy+l1aXqlKYuYS/N8DwHB
Rade/Fwbhm2wgPt+WFIvGEFMNnH7o/JLXPQQ0C8nUG4Yb7y/axxwA9Ex195XtO/Y
Q7z4ExaIYpdTDUDyS/RH8xbSDuNY5GgHIXSYxrHTwuQxckwNCc0RxT50lV2EO8lb
tySSoWGIf4TPgPJlTHxY3DWbZuw6nQyGOhu2EpFTLd8JwTGWDXrPi5fUXnk8Xaav
UkTyfxbU0Aq++ttw+UiOsEBfYTdcLUDOTwee4iMSy/Dyk0kxCc0N1NvhGwDTh6+h
gFlIZlbrb+BikRW/sWpRMYuQoqCSMUQrroZVe0zyCwNAdxWcqQcNTP2+IS2b9Lit
ci4mkJhON82+Ub1fL0Vt9tA2EbW4O77VFi10sVw2wK1p0etTee0fxnfDAVPF53em
GBV0iQmOLbSzF358ynz/eTS+BcftlPXLiYWz/kYkELlzvs+pn0Z2w/funnJ2yjdS
e850jQ4yahO6rX/ZP35BAYW9llVhQHCu+P9qEzC/AzFckkvYaLXVTrszXFPKIC0o
oBM+dZinkF4rNpZbt46DpuWdWAsDjtfkd820BDY2eKfHqSWijqyZsqwMlHSef4Oz
xZ8IfxnHZxjjd8bHLXkMDvRfO4QhzEnwIdG4AMM/vwrOr52tY95mwZoeCpdQXCDB
867t2v9FND/cuaaCfnXBhOzEFoErSFZ8VzE/X5R4Jn11vuwdhWL0KBYrQB6LWmTB
P0PtM9zOzNgWT0ASSPcFM5OAavfnr1Zc5ftJB5NeVeFWCHasxXNR9drsjYx5DBz4
zgq9K79zdgcvjBzdijKiqgPJshCHC47mqEJAQeAuiLPsZintS+Jl/o8AIZ32+3zq
jvpBQ5FujFbwlC6a8yTKxvcvVfHcVBImdUdKb6CWKZokH4RrrDISOZSdprCXbIaG
q+KVOeJYJCrFQSPdfC4C6iqRCVNJJ+2d9u9ARHFhzhufSLfoGAKrkut8xLiv/Yaq
lvXIdgsH/Z0qe0lj+rWK5IdcYyZGyRe6kR1iV/K5aKR6s5Orl6iJk+ePHj/MpiYJ
9iOlqnn+AtcbnJUNxj0BpOagQuBLKoUI3ywOp0lQ5ePtpH9Sd9S9siBKcYtIt30q
QjRFTm1NnUSDVg2+CCxUVQhDvv20SSGx/20cMTtv6H5EDeu0j5lwMDytGSch0LZh
EfbKteYrrpzNqu3ukxYpUZvsLzyeqoOH0bJ7QIA5U+XOB7NPor6Yx3BzMMe2iofn
0TtxsTSAqlzK0IjYyDxxNmmY5jxYTpgwt+jU8ElP5HcLDhCa515TZhGt1JDxfvLh
BFEPU0cqoh0UXzhgsuBnRsvCCHUCcVZWmv5K2R5fHFL24rKPz6ZjGP0WzcXGBgIB
jhRsSosscpDy6ouCBvAn+pVRUUbpow6uJYpMSebG0i4GeKxNz1daEktURdqDqf9F
GU5OZsc9n3i4ApIK3sNt7ESWvE9gz1VLPQy9dwxP65MNzQvgG7EyusysEmuPjlI2
VoRvfodWvyGcrGD7GHNp8gid8obRs0uaCf6gLoWnpUCCIqvet9pVjE1oI/VKzucN
z5etStXej6Etc10y8O/QOTJ22PMy/T6ODdUEb3zhdvN7eFdqiIVpg9kt1j1hzgSd
9gOq2XciBxl5FTb1TxFXZM1IfiuuNUii0Kfqnm35//8329mJYnUXoI9ZXyyqYMwp
oUWrG/aKEKo11crpX5FRMgT0fBspBuu4cgU9Asiuxk0nnx/ZF3VLd6mWnCip7FqS
it95malHkUrtsuR7BRpsRNIpmnmyF3CBGopOIujQ2R8ci83ORCLok50IgHpH/e/F
xd4c0Mck/9uEmkoz07hKz9Zm5qS20yuBiZIgHfU6TfOP2xlOOyFqiKA1FI4Og/xq
tTgYO8NTwRMOKMIAfMu0FteHPop1sB2d9RSvDpoXOQ3DqS6UkVrUnKyEEmAQbtr9
ElatClHQyrn4hahYZjffTG4Vh7a5AzUngUtJQ/2RmtDzFSRxPDvl9BaBeZeE2swt
eBHT364P3kbdcxv0ea0RC4RYfAuD5fzDi8bXeo1oSTUddfQ/yWN0/UCeToa6sD9D
cp1hSCQLq+0csL3jBxgnK5Qj5l+tcqgFymR1RhX65Dfbx296odSqPVoEknB90ykj
xtyA0fo71JDIikOTeIKtRzxxVORFlkMvuyq/tqTeFaOXJs4kSKX/v6AySdh+a9SK
awAPJIYx1xR0JF/Lc7plpfUca2S9JGVko8EeJ+lVifQtUQIbG/3LRio4lFYR/f8F
jICHqjRvLMp/NugzKHqBrRHrMJvjsPdfpFLniPFepa7b9AsBGeZfIEMOnGWaL9Yb
IvZMSKctqxr8x19nB9tDpFZZ4N1yNpxhuqO8CaJa3isAHkveivgrITmuVLUbluLs
cj/WylOBu5ZNL7+bwa+JSSMNGk+OLKpSyvmMHlA7xypBF6gFTk3PCTzr5QD3xCLM
IV6qVDSJ8DvWth9tnDz9wX6HYF6O5MdEmQqG5WkHZ4yGI6hl+RlOz6rmOVQhqjdB
d8gGadVh9VwvVWmk67yG6mG/dGGMZ8FLkjA9/E/2G0iEfjIdYyKS+dOoso5wb4Ov
DFZv+glOVmsC6BGR4l9araXmOPBgYxnP8yKftl9WNeuKNPQuJWcl8IpNVetWDN66
3ElJylgj5nY3lN8e8tYJSQFSW7xBNHqbb8HQsBV0GS5Zms225D8sXcAHs06G79ty
EkIWRe/gawN+QBagXAl8DVVzakvspyOF05kVPf3c8BygQP6tF0MrMGGJaJCoMD04
AeXdqJraMW6SHQ/uIhGSJSan52QfLLDUrvN+TsnA6WSWHbk7nV7dx+IXh15eaFXc
pfnv8jsoKh3LzeF3/urWbHPwTZpmE4CC6CYf8mjVcUB5BO5VDn6GPU/DR2/Es0WU
Iu/u6AVJNuqe4XkBTM++dEhgH6dsNJ2AnpWMbXBfdLk5p4NpewF3FvmqxoUsVoWl
DipfSo5yh+qRx90bMMzLyTQnenwW//C/agLcXCcCDYq1/Iglkkbqm6YHCNJEOC57
D9h1mV8xmCtsVQSBPvh6wFgWWBgqcUg2ayR0URgYgnRabRmxSjQEm2cEmOcq0z77
QizUMg9pBF+Tu//fcCAOB/tqz6SW25fvs6iZ8fcUsU/ADrV4tD/W//jpudrEauJK
QBPHbOUHKhmc4aCGd9QguMVSoVWe2YX1yFbbwZTmxgamU4cw5OMYuodedaHw6xrK
xocNX7b1tD8agQJRFrz6mGF3+ILhg1W9ijch6DK73SMTWBeC9AgBDObuesOeVW4Q
b/Eesglq1U12fZFfUbKFi1TY7XC2DTJzR7TV5kG2+Qr6h5xSAaOF1uEcAl/EQwEH
L+8kamV9YqXYV/66O9n9oYpAxJDJAke5e7KbEC50+CgCCuv9C3guRJ3ZRf4Ye+x6
M+O9Acw2LuTYBAIg7+LRjjTt8Di92H9SkPRuvivBdTjAKHyoCHof5DxKIsXj1QG1
o4iIzf73zSjM8wwQiS1Y19P5/18p8eAAtE6ujBtE7mroxzerV7APNl2nKWWYgA1b
0IWXQPbLxOxAdqFg+WlGu9V+5896Zquu+kG/yR+axWWsW0pCNq6MgXXlRT73AbXv
X+LOdn26XcpFRiRilGo9eHGydoLElfiM+1AD20EHVW/VJEWKINJ1NPZ/CJjJ02Fx
hmfwdk3GNiV9RYT84mv8VlMes1P+59W7LLmNz9dw1ThKdktXaRa3msBcTwO5SL2x
1UCYjvtRv6/d/A7EGLh0FWzj1wzm9dKhNpsFK5u/UDUCNGYRHER9xBg7mbIlEyec
cpzmKVd0xViIeABtzF/okR6MML9DIO6VMKB/cIM28+UZEFDMrXZsJSpinRnMaO6e
8BdLTREeF2ttL0Usop7NhzuNiIpwf2ecBUl/GM+yJSXMkvzT5bhZ5bFSgE7tqnt+
Lu6ouqyKz/pkFJJXCiCW2PwRR7DyLKhqDBTyjdCdbLcYZIT5GJ9/MIvwGMrneKj1
xAqMVGui8vnNI3AHOQb4obXlrtzaMeaZyPtC4VAlxgWxW9IvtBgr2ZjW/v4QLJfe
Zpqfzx1fCXF+aotaGtdohQP02ppB9lkCRwIGgsj2YinzTzUm0HB4s6YhoVr0qa4L
7Noy10jqU/3EZZypr/nYnF6gJ7B9i1RBW+1G3FKB6afYUkdwOZI7BqyaPr/HAPmu
1avhkFno0LqWbZ+fX1zTFTZW/3JsVbDs5koEogxEBqp6QSVm9bBnyEQ+n540j8lt
85aBaVGiLmBO9gwmHCOyLb3U0l19SxgA4CqRPT2xEik2AxiciUKlRCC/2FTffB67
rJBcZ6FKlHsgxkdc+KQrzr0TWP/f582EBC2IAIlgar/tLc2IqpAglaK19iP7oZVo
4yIYjRz2VJvNkM9gbodfJEjb/kphurxdZy+Vl7mcPZnsTUfYV3zdlLh6v3zJVCOj
rLvt42FAjGJR/rboFZGzREwaI2S7bVKvbTrQ2hOrCF0ByKi7JjGTQEJ7DwUpjC5q
69QOiFt9/RRF4NsgmMXsp8MiCbMNZvqEEdMHGcvDRiGyDJdS0zh8TP/jNyPrrX/g
9l8wggWEZjV3Q6Fo7uasrxK9EG0MKm9YGIL1Hwa2mWcxQgyOX97kIl6x3Sddntwr
Sg8zE/TUU4u5tDXczF882J5EK8LWD4kWAXp8brxvgk6s30KLVTc6O/r+lufgpqhz
l7kyO9iLJdoA/CUmEYINt4AyPAdMJQTGg9LzzB+0QLS2zZTLCy7hluD01gx26uf9
f7chMLNfcEfURfADjDADifUw1Crr3T3KF4agjyFv1h6Oqmr1phSTafesQeNMy0ib
MNxRGW8K45bpa/n6eOfI6Kxkk8s6TiWAKRSRrEO1AB1vRDhK2CoiLOsHijcI0nUd
Xbqkkr13HpN140Bqb+PIwgNhcjRUA8l7EqJWOoP5VnvwnvYeDCdTlYNiPSeP2aUL
daDos6Z7iPPhfAg0rc3ko3GINFqx17xpIrja/Mo8NdMRFutaoyhM8F5aqRi6abKN
Z8Qfsv210Mq2ZaxZluk0qOqWm3eHSDVd0NVHKR/shIrz1SVjD7FGIEGJ9fDz1lHf
bpmEXrzmgHitSeS1nZFxmkh3KzgtK1ufzPoME2zRWvrvVwt8QyVQ6g6AsjXRmxjZ
JshgbyoGEuSKSEzKlNN0TuO0b1wc58zxNU/g+rvoGy86imzLOfbOYe5Ks6EQwIS7
XWhbYg+wVYqZQzKMt6w3xwCSK68Gg8CF8MeRpzw9LfzSKHzpNmJ6z3sor667q2J0
9p21cOY2pdCdQALroZb2pyffx6TOj41kFLJeTTA3TQy4LNqNjWhWf2iwmgyt9xkL
PhvRcKZ1qskSnMj7yVxDErbGvzqdNQpUZJIMxMxzABktB9uyLn3AkqYOf5JUQ18C
OmDs0q093R3g9g1x4asX7hhTWjHdjp1k4gx2I194GUO0P8f/0jpLbJ+w7cwIg/OM
/WTPAczpFYxNLZ6d3XQPk/M1YDrFYKA+PYvv9RYdGFBxAA0THrs4dy8BQZhm13Kk
snyPjoyj0gWzmol45R+NFYblm9n6emzgDNuzisB6EGg+1jsEuRClLSuTjNTZgEFM
xtq4QhisRk+mL/fxOVfBfzvRK+64IGiThTsDj53gAJ63SWYFyJt3YaiibzSwbvwJ
8cMzT0k3Ht6A40dFLvMNszP3G5hlE3x19cw1yZJvxawnixV4uvmQjdDF+02L0nTj
NHTkNBaf6Yp5Mqgd3UStUE7r/NMFowYP6GQpP/JcucNTMQh5QpmsaQztF/871+TY
bSyJW2OkVD3HEBckwnCYFNrPcV54F9i7ZfooGpefsAGC5fFNewxGhpmvjO5wU5lA
XyYOCG0XGNM8gk2/0QjijDWTOeMZvB+/GaJruJo2s9/WCZogRelL7OrhuGEIrAZu
I5yp3pXGnJR9Hou+XHjQokJ19oJgirxZxOKZY75IEFYvAlsJum1W9MLQjFPIsUk8
C8edqYXwjP76dC/AztOwd7DXUZfrsKGUx88BDQlhS25uGRIO2+l3Px/ulcJFjlTX
T+0XqvWeJO80tQb4Ao3/S5A2LSuOqAFnYOtF/prxX7Bb9heuftz5yPapoue40OgP
ky/8S5JkllsrCNA9XK9on/0IG9zFb0lu/CU+mLOhfh22J2pbOQ5i4YoDM2+9CrCJ
wiOt7QZe8ZplY05KWXmcc4dmm9pDXGJ7xNDrkcTNOx8yjsUUx/0UROMun5+b5gKG
vKEyeuhOSUt6jU/zEjJ8G91FuOkVtSMox4qFMx5k82qmTJ0rYxDp+nlsCVubR+dO
U+Nknr/VcbNzfK5TbAiRIBudRJfNKq+bwo+3KCKZZCAX0igHQTrytTrfdWdBjEwe
t+MfZkMi7U7iMSppcUbpa+LdO5plyVPeGCOO51OWXGU2yPYrnwMUyoWaOXiMwULk
68vrAa67DC8U0FJmSnOFfd1KLlqQkcWxuBvHetKlekYy+a1cwmeHY42BUzuiZkKp
X5oXEF53h3qzLl0/bmpl+/hSG8VX+IfWwo+jSaRh5MHhQiSCZYZEGyWreueuaGWf
aoXPpZcFfK4r5PcS0NdqrJ7oP0tBDJt1bKipLc21ZDEiF1mIG/Jv9NgF1FTmM1jv
Y1rmWTUJWAzt5WndwzxmInoFgqfNd4W5qhRXZxZwKGmpjpk5t9kz6yAsOkay7GVr
GBjpL78VLslPvK7XYQgM3pZlpdTBQpp2l+C5W4eldwykZ1Fb8VAfImJWg3m3aP6Y
JrNttuxHaZwZQSCdK7+z22K6vRFEetbtq7P0oUiMnZUYdsE2W+Vc1ZZwCGOEhrDe
A5TtFp44v7eDPAuR3baHtMkWKvIhPOc6nzb10kRwMfN06ACf1WlbmkQA444koFdz
GGRpFgDOgcEdaAXTZT6V1yy1iwBKkm0k0rWFiZmKe0KA5URYcF4OE5rGvZScZYi5
brRMSdTI1lm6TUsM1JnsqWm52UDoB5oXeNGRwCzIMmtisT8ni/4v8QGhECuRILMO
e05Ezu4g3OOA/yGAzV47ObgjcIo+RfLbSkgygkDnurPd2xLCvcqhS2191Uel3+CH
WcgRs4KA+NpirXqcQjKu9WBzT4zSat//Db1T+karTE3Rx/eR0IjtlKTR7Y+L3nlr
wMLzr5ZMiKFM9W48+xbn/Sl+WNg6Q/4pxQMA+rLhqKiW5nZJe/nENRbc9eEL/c6W
CRkIckEt4RhvjwvhMh4zAvv269ctxaak8BfpLUh+Ym75P9FkaD9wOnc8/NeJ7WVt
wE2ALUvvq3Zd7rglRF/3BaUzTeyTjEY0EgehbOFOs4yUgZshKIzKtMt+dgqRh+eT
7Wj7K5XKOZKvEHrNCttaiGgCoKiL7cEIEfWCl1UkGnc+XwYNEKnCI8n2rh8NCezW
YOoOnSQHf6dYQCa+9OE+4dolQaouAFDrGphs3Rq7EcU0OlcC2J37En/QAdXVmV+j
YIjrcuXiOBnd34+gb2IKkL13Eq26lb9pop8pkkWIvPnARj0UId0RvJ+w8FIwPIU5
+HU4M0PuBYzMn0Ou+68/9yfATQcYJJaZGVl/ZaF9kGMw2O8GzXvNvkUp2Ns7QBIC
E3V/TzufcdVmO9gDbeKBEmEaRr3H1hUZ/yeuGU5EdZNkhEIeOPSCNeKb83/3j6ZX
eCKkaOoKo+hIj4CJ3CFC42v4/XDVGdsx9m958Gwi91HGv+xkvwtLWeW5ub5/biV5
z9Hzo+u7bBwx8PKxa/TP2JngqZ9XWVh6D8a/K1bO3JuYjRfL1dSe8LOsDwu+F9v1
h/AkMVzGqCzDFZrAQGowEZ4u473f8RafzVVhlJ/BhIZudtBXUDryVjdgeaUaFYjz
Fy+Xd/aOl6oHUn3U3ghL0K6p9yOePToKV7cEp6vCM4PNYP5z3qV72TBZg6CLh24n
Z3GVEvCIgxpPl2XHaqdznKj9ABgeZeI/mL/SUVVgN6rv+JrOv1gyf51T+68IHjHL
Z0fQXwhXbp1IkMUa8X2Jc+J07lapLlf4F7woPTsokY+utbxaPpTV0GYqO9ohaBal
18D2VaKixC7VGCyMpwYHBRFjgYdixtsjKiXZ+DMYHEkdXXuptPxZunlS0XzgB/h8
yaFBd8IBYbi8HZ3wfQjZtsXi2psdM5gXw17EjhJ5UV2NsXI62XdZomCwRIMrsF+N
sPVlOLDK/2HC7vq9BGQD1iE9fIW7e+Orfe8246ThQ7Njm5C+jRGikzm+wlTZYdpy
XJwNBQZIZmQUSGugBb6UKhWs12q5hwR8i2oi5bQ6Hm9wX8k36TvfdCCE4IZt1Lzn
5VMyGPl0KMJUR0ZMoV8GWvupLvVp3ZPNvSaXPgu8KSQkHk8LCf1cXadZExxOM5Fo
yLSKgW+sSaHA94A0/Tku2moQy5skFK24mrgg63qXlpObj9HYj9q/pGhp58PGt4j9
ChW03O9Ung4uCAA4Y4+V2NDFkUczKJ1Q6vPinZ70ZQND8MSUZnxHnAYNH/AagJT5
bV2EqB65DTlI5tpsokW+uIfweYOPTZdcILHovmnfZzj33e8v8bq+O8Rl9XBQcWMi
aWPd3WriIBwvjretvZC1UfFaBGJQsR+zI8pJouS4FgatWa1hG3bUTaf1IrkEoIAW
uFgVGmGy3tS+mxX+qCs5R6mqLcfZl6LQr6XjbQLhq795cf+uPBxArBkbgOK2pgQ7
VwFAdley1cRbEQC+jFPvkz4H1YgjfIiNDl+49WWIbPSVGz70BgXcwV7PiossYp/i
XXqexynsA1UDx27H40ZnpGsCM0j46roP9a00KQ2LdZhbpxN/VFjyOoPtQN5lQ06i
+9U8gyfx70MtSeAWTUAAbGuuPMAxJy29d9rH2NEs3S7iOdg/ui0Hpo+QgsKaZlWL
uB+XlEwHC7y2fsj3WBbKkxSjqaK/+OsbFL+fSeI1pJhiO7CwmXEOTp2o0rj+JeD9
e/2+4sHOs0nKJ5PvljI5OKgtJZ+AW7b/Txkzq6BsEp8B8HV5tBeGsN4jndLPVAgx
TvYByR+3iqFq+sG20FTXhQsZwZK2emHv+7i+Ibn9BlwAi7VKmy2gPL8x//6bRMJ1
qRCMNES4szNylUgZpQbst0WKKRGcmeTtYbvKI2lnFQJpa++PoElwmbMzLoxD5VIf
1fg6tYaHuLtrXKlHnFzNxG6ykj+mz+Rkc9+6ebjcjUxyXE/OnSKDPuAlXAeHvJj+
gB+ClEw5tS5Rlp17CEGlm86yvLwxUEbS6BnkcRd0GlHiIZ+XYaBCs0C+B9p99jQx
1vJQm1qcm9vc9A1WqAzvQoJdC+gQ6sg2Ab1vCbz/lswC+yeecXMSXstU/biSQrHH
Ka9bgAcirBVEqJQIToRNEKEQ21wlbbfAZEC5eUz9F9oL8yY1+VPEN9jqVd1c7H80
CvKyZ2xWPOrar5wRDy+UGKbcJH9ePAbLGe4/oZ88L3FeYcMjKkcnykrELEBRJc1y
e1A1BmYAxkgFTcIqq00wsqgYwUhneJ84N/8BAi72DjVP++slsXtVzitLs5/KlIxi
Et292YmvoPdGG9vyfGo4SuuApLwLDzAR/brlWUV2npGe21SprgoPtnenL+hD+S2n
n9pdC/bpUquLlal+OknRt7eDxXIPFBTUu2gqfkq+dOcFO/a2SUdHP0t4UdSjH9ED
dgDYb8In2reFmMHbvSF9Kae/pm00kkfZZ8CIEaentNFC9l2NNxB1FPFzUCI7f+G1
rg9YAMA15g09TyXJZ0lopt+dp9WDP4HWrUMM/J3lmTMOPlXQVDpb4S0Jy387RFt/
6AXg0EFYALuwVLyrVvKQ/tt3JPa3v15/WKALusbz7kbT9k0v/Bfae6ZV/2unBUEP
v0ltzVEiwPX7y5Db4B34e8gKHSaGKigXVOsAb/lGmoNvItaq2rbFD9M6tqdKAjfX
U33M4jbezHtb8/clt5EZLH44ilFBk33lfK7TAU4vIeH6yEoA0qCdGgqbvhVhZyUF
MSI6dnvIfe9ECYGomnbTPk1xn4hHCYUXo7SjODbwM/2dWmcxKT4joMPLYg6G6OO2
GjZPU7XJ59XRW4SxYs7sos9mLDAqu8Nw/30zynzhnJpql/LmUbpQ7YBP0rdL6iZg
AES1eGFUPJ+dQwGaETnQJJwkbSo2x9sb8zhRQ+kiGdG44Gk6GQKIEV5R/RiBk8rc
gDUIviSfo2rWkeI+Jqc8+vtiVQ1AFHDBc6Cx801qlpbBhrnsny9KiM9O2IDJm7e1
mb0IB1UMRA6AFLEJjJAm8NnrpkGjdzR4oRLCklY6n2mmNy/Cu+BU8Ab+zIWa0Hwy
3Ad3hn5dUhVl9SG3e+lBpem6kXZu+z4amYA0b3g4ILWelX7GxkziMcVRbHSwvLNg
bm/akxvTViwuhNzlnMH1lCZARwkQ0vQtGycSKTOgyd7alywDONzn4V5DLZfyyT/Z
jCDbz78wV1rtpMs5NbLjyFLsdaPCadqEBHoniHv57UKoTmxDeKYfrzHZ9aFMra2z
5ETkv4JaEjFliTU74RkBQA4YmZv751z1zcqvmpwmMbX/XnLVEOIWxVHaCcrXhqIb
SI9ttIT5+aVItBNCQWdvW81rXHng7+CgfQQbQk0WO2pzkGtigv53qH4q0+2WPung
ryLAFvxNFnHM3BBm6A3OuK6vIWyDhdqMLtnq4R/WGLF/P6UOuRzieI0gZ0rlwkDY
LHIEy5uZVNRLTevlHTm+ibSbEFExkMdYnfJpm4BLAHZcp/BYHJCpJdWw9jrrC9Xy
LM6OF8oCt1B1kQVWtm34pFkQHSfKFaPlBKwlxH0dqsGFVBq9eUvWmrCS/5gadezv
u7sXhvrQo4DQgUqf1NvZDOIHS1V1PV0VmhJcfaSFu4PBimtMjbyirhY+S4qvUQot
njmbTbHaSihQd22w90RghyW3fL9ogY6wMgjG6ASTgiEAqLRtdIoxRC1ofKOsZsNn
18F22f/cUP+PxzuMMJzy8xtQ5l4Yx8gDlyT685SH1EkfZOQCAXUlS6nYOOVB+Bfu
RSYkNFHvSpaVFuCTMu1Ip8dU3NmFlIKa9HxC8ZUc9/+O9mqRFfYEInOHTN6V1nBL
IAj3q+wWA3+J+iJt+IGU0FsLqo8jk6Ztod8SpgU7bjEF2C738Eb8ChyWSOJxTVGw
My6ADPc8ywIKL1OFy+h4+BLmkzGhT9qFX8PDK0OCPLNPk7zaP7784SfxjobXM99z
aH6bIRwFwqRd3F4vIcN4dO8uo/3vxpNUwS+fa8Av35kq0ZaeOJHHrZw/J6b1UUnU
YfHaIo3dwwQQYEGkhgLyp+vC0SbX9HRa3V4tfa+JQBIhb1ardrZpnJZVTLMTsmUi
8TT0qS0PxAFlCDr24Zrs5Cl40D+Vw950E6n4fLieygwihQ/K3vmDhMgWJvEjzk8X
FzFqfffkBjMG+sAV1p/AyJlZb89TcZHP4lC0rhdgSQXRWaYtjNnQ/VVgwKWraTp8
D+IlNTy42ydMrImHPQokqowyN9vz6QHcrtDRrsE/cCkBbDPHdtUTQ0XQszV0r/mN
BBaqa0W1EQdbI4FRZ5w88txKvyyBbhiHA8paU9wo7K/qsZeeTy7Kxyaw0IDUBRlt
GkY3jEvjKgPiNe3AN72pLzQoNo1wfid9+E0noiYI7m+fwW3vXarGhoeNF0xFj8Go
8j1hLp6tKKcSLXlk/bOzQJ+/9agAoV8oxvXPJwhAPABUfx+Tt48ZyMQPtkqWUTT0
beYNxG2/KAxRQVg6TOPIPGfi5XdYBwkgE3ZCdWzPaL74nrpgLOh8G41krTdwBrlJ
KjXM33Bn85p5vYeb2s/AllHi57DLEsUBLaAWzIes28M1boEA90h9Jyms7G1eHgkZ
vvl2nwStLwC1+0FCeTah5QbuimO8nFOLnuJDgKQ4TB0x5ZTXj82z5wSkMl1YpFVc
mLKeV2CiYPEnHThE3RaLBbg4aV6o/UNZYzmex5RTOcK+iRN7Ge8m/QKsoAERspAl
MgQjXWfLXy57MZa7uFa6kdBiP12Ee6ppigwIm26w4glLXKsjr98Vn9ZiS5lXzjED
ZaN3dAL+mbT5Gk3xiaYlUV6tobv9c5VqDFGU4Kx2w/OpnbD3xH7fjYZO+PW7xhNg
anUOV5xFvlnAf5Nzdd6n92lPjeu/v4u31y4/Emh89GJBOKN8r3ShWrrDFXQOCR6n
/wH81P6oQdkZY7j3k7dXc7MapxX+/gQte3spHuEJ/Od7PGEiN3KUOWrGn+hZFyFX
gnRb47kmGGFxsOkjXfVQbAmvT7gma+/700hWC/r4o8o/wLggh53AASl17hQDP8Gj
ijck7jOVK8IwJ00f/385DcPp1fysxVnMy2K0cIw2RBFiji+DapHz/mnrWZxmnkgy
UzMi/Y4Q99iKPm3/o60Se2mafSZCjitrCzye/VRSegF6KW0KZQih+Z2O7FZJEp3P
BC8MeNDNkOYgYELcTrPMI1rHAqJF9K72g8kkD1zxqkFoWiidoqt37/XYcNQYeSR8
Vr2z9sqpxeuh5j0eSs9yCSyT++GdK2cF+m9I9zO/RhywEhjDQEsm4VFjm9XT8Uyo
uOQdkrVcwKFifsGlLmOEBvtJsQzvhgI7uc9rMJYgnWfzMJtbGeedfeGxwj3X4q7f
kOejmfFdyq+9GF4qgar+kvxuq5hhFtoD/MimC4X7vw9gopzNDxQUuCGJNtkJLBdI
kcTzna4SiwWCRZFwVZ2VrjRnZeV/7qOFpNbJ6uOUgfoj6JUmcLgQiHO8WkUnavFR
T2QZCKvYY1SOL1cFo6xzrP5mdGOJqycCIRqrVdHOaS0A4qP/moRUoYU68zYrUiGP
td/OugSwT+zCqYXvDVD5/r3mYvyz0s+/YJ74gT3+xj7be8SPC2sLm69n/2NlHrVi
5BejtZGG7Vcky7gixZAROvhOcFv8Hpw++6DipI3GP6SSuWXRuG25iULWyBDhozpC
rksc+GwvbTEfTcd1hOZYE6kqaWGsLrRhlUF4Lm/duyfB3yy/i5A88Qcuz11SBxNU
T06rff1QmuxkB8SF/ygo78S1oJKVETtAgYNdjcWFverC1timtFJQ1hspWy21sN3Z
4Sl/Y2oxRAAAfPX3IKATheanlMwYvxfR07JEMM/AK0uf2jF1C3I50FtBbj2DOLPz
O+21RprexgY4mMZsfTox+F4KPV79DYTr8vrc9YuKx6kYuFOQXGpgf4ZtRDRjkSaC
RUckx6xZeObVigE6UG8r+6gMFfnYnXiauR3bfXqm3MtSP25hdci3/xURfA/ZKBDa
EO0Osturth7BsSpJRg5UzUvTGrnV1xFXPKKPyqSde90RT/LuBTw6wTlb6uiIaRKJ
wqvWFPlhpIiJWc0McZNhUA/ljTUglS6h9alThPdJIuUCNh3A2ClKQ0E4FnwSDfdS
hoc2/NdKbi0AsWthobABxyYvye2A6Hv3nk10Tsa16dTz+cy55DcPxEi2gaEuNUsp
+72SWkAQgTABxWuj57yVhhPkX/yTuPy8yaV0RpNhiH9aSGijToq1yQDnUBojTC43
Negk44AAMVkKlU2s0sZPU0khJxv7d64c4Ihdq9yfAdFGw60K/Hz2EBJRTUPeG7dD
ZQN+er02RbtAhYNxtP0cyn3mF5rn629hAfPnG3lMLiQ6EgEW5Xying73bP/nn/W4
Z9I49TI7qOAh0sb9w3t+qOAFSYDzUOw7camdyK1BK/RPSWTBGMdihAmp+aJupHpD
iT5VbE8KKmr1f0B03HGgkJqyFcYqjWMAS1vdUhlZU9Zkjusurs9LWRn39OjyZYB+
DKR1OooK5g+g7TCxZ4EBSc1dev9g8MOuoTeSX74vB1mUgLlLY40aSm6aBvDDjz7k
XsT26JEIwggkq/WF03pNjICjrxzYVxZ6UjJ4iDcmecDraSwjBAB4JXmAsB7o5mE8
tRlf1AxPc+lKo7Ih8G/N/Zc6F/xE+UiQ1MrkKT/W8y/RhsiOceghNiMeX4zDdoeQ
zVrLqHtS2VAWKWED1/e9CsAA0led0REUGvvR1erB6fGghOKSOl4UqeGRCf/BMgyp
uO5un4PYnS72eWypO4zmg5q2aVHLnHM+Xbzjt2bWKZClLgBbCN+tAzu/dxMHiarJ
w0kJziefX8Fv8H6qdyvw6+riXRctVy7e3PznTw9yX5iYwDpPxwqR2bAax/kRusUv
uOHj3bQ9vtfJEUwVosljxAyiGcjaJ1O6USH2zsmYMFKCr8Tmn2qqHpH+R4inJhff
rJlN9AEZV8KYwAuKkVs1FVwDNFrVal1ZusVj5UdppxDp6g35fDuXkzChzU6gaHDZ
azpubiP5BsXfkPv4i4SkEM8aMlIig6hVJcAFdmzejYXAip8Olg9LCnrh7fsNI5lg
EVPf2N30Wkw19AA6Y8oq3fK8TjHcMB3lxULOjGR/JJ69TLh5mA/X24XblpU946kU
IAJyauibPWDSnYSmyKVfTf/mFratRJ9E9M1quMFoSB8COwTKDuGxVLRGGJdi2A9L
PbD/w2G83GKeE9P7gXfEK9tIFzkxoSW8DMaoaqQfskL3LN3zFEOMYmx4LGAvPu26
oVfGmt9oq4MT+1NwX0iO9n6eSulP88NBNZv8wtSI/PhFJVgt946iKyhWgvxis0eQ
vv27Dv8dMbtvrOxo67lvVYlPzzzQs1OLEbSfL66EG1iqM62D0RdnesgvSKW7MHkf
hM7oCZdxmS4/PgAUxROgxYiLGjraZHdyChLqQi3LQ/26gLooPQSbAt9fSXHljsCI
F+t5fZii9AH4p2+9R0GI1s0t3EDV3jvFF9+XN33XV4E7v7UkYIdmc5Azw58fsvU/
EdjfQA6bfVaw4gZcvqkr6eno8wawc17RhFwXljF1aSzFVffy9W5/iMc++NC5e/D0
MIGPlhent8kTH5HmrCdnpj+rfeVnXvFwhelsuazdjCSf2R6JnyYlrlHGStRJMp3z
T4uUr1V0vAUymsZMct6GWRUicF/Y5YLjUfjwQUZ13bXy/Ip7gXXMpUB3CfNO60z1
WJrjdo7ni9pFhDcrzK9vqbZH1acjysU6sGPSsQJnqKLwgnj4xR5a3zKkGVD86lfc
3/B4MvDgOOw1Xqz4RluY0b72D4fN+58N5KoMDZpmemVDUwqLtOnExbbdtM3oi3iK
/p/s6XxFBYnp1oZh1YrkvHPOVykF529rq8n/oqdQBFIw3qb/Iq+wJOPnLjquIHRn
QTDetb8FBEWheuQOnYv3t8EZqBbOuNKR2tzb9aop2+PuAIzhO5bQ2hSFzasFhEnG
zMikE8QZXCo4MJ3LBmp9doV+kFeUNNzrnWmywNQrN5GyB5ud3aiNK9LZvvvV7CW0
kUrvrriW11MTQJioOVar/z8d1OqXOX0t5Lc6lx1IIkIA71qkwcusOvTAkEHj5e/r
hwqvdRCTtEQODCgfOVvT8tlVf3OXtnm/rDf+70B/M66W0jl6e4UL1V76+lBFpF0+
asTjKOIj6r0MtIgTTZm5cUa/vifLxxQhP4UFVFZ7Jsxr+MWSgwALHpEC4YaBUBA+
S5NyD0GuJVWSL2roviZ1HbmIXRoGxEpDoN4fIciCR/aWEErOYh/0eQSaL9y6WA/m
pYuGYXSOWEkUnLZbkzi7HrK/Ig4EQa/qVdznxkl2tRC8tXxihhTZVkDWuETI5XOZ
RDgf0SPMY6QlxYMpygODhNw/SD9mC4s3hyCzqTCkqt8RLWt1OFB7PTMDuTFDiFqt
IF5+ksgWDU1mQ5RPJv5FNJU9zwfjE5eGiwSoAU1iJHMAVMbk4fR+WaP54urHQZlg
Ul1FERk4npJZ2muV1StxuMQMiEZBUTkMhLWJChIZ6CjTBcJ3pUgH8Leucbjp+x5I
wv2K+DWOSM5D3OjCR/OBxxwnoZw6HnQW7sA49ALftwt3FK1RRJyXNZt8ykGouX86
52EXrQyVahKtUAceFtouRJfNECoj4lzsdPyYL/MPaOXhWXJkViqzgZjXUXka9LGH
XocOOTZuYJ09LrQ2+Q8x10WkCtwJoTaWQAKrHS93HvmFLWHVWJMaLUdK/IsSJht9
OkSW3mnl8IYpkGOzx9s2FaTkSDzB6cGJMViTEbz42Nleum3QSaPGaHXFQ/Xlu0wj
xTMxG1erxL/+vocU5wPOA3S66iICioIszEcpRVkTHu85TEX+fdBIVh8XdZ7UdCAJ
DzCYa2UKiARvuf2shWwl7YcxfpPvdZF2rFmrjsX0dTrCNS8uMuRRMjlfHqV0JJjo
MIemo7RIEypb7E7uJcx1VA0MP9XXJ2p8YxzKThOcLz19OAsfNy/OaCuTK3pDEeg9
mgClZXlDtJFd0kUrTtYS+vEYp3CZ06Eas5NI2gNKzbgodE06uvI843GHiqohye72
CHZaLhBOL2GTtpjJ7IvoHGWWk3MvcPR8I9HWMf4UN/5Vv+xPbO42j/o7m+m3e8fD
9UZC4Kc40nkySRC2EhHFisvO7fqvqgE6SM4H3Pmzy40zWWFBhot/LMO48D1rjWSP
f6TloBbyu5Ol4l4wu9YjVAMy5KoIjYMlUGf9tSlFXhzSzvqWJIFG/anDaZKgd6UV
cn9o3xe5fSKs4pG6DUeWH8LDz8cYlXYhEJOyxHJCKUQvF9uXzyZctnPVYIfLhkqK
N2E8sEO/tbF+8aJ7xS+O9dPuvRZ3bAbl6dQJ9pN42zt9Z+uov22+48zxmOE3XGqS
Pf9CbhE+cFYzyUnjhJdhPgC4cUpZNxtGMM4V/xjRHQ6XdE1442T4mvOL/H+SDfQq
CF5vIjQx07K2Zzfv928H+Nit9nrb/bZgDSFAG8RxC/UuAHi6j3WS9t0zSowT71EF
5sy/trr3kVz1Alm5WNoSDffmcykhHVeScPcSCXvZzKhLQ7JVj1hK2/085HwHQB8T
FHeqv7hc1UqYIjFIbBVpfIaZW2URYFdwqIOUvG6p8Dn8UPnFnlem4fBZxP3xfYaT
ABplQjGxrnBKQa/rURZgjavEZC5NqvqJhJ+7+IChUS+iQcc72XxMBQi6CxSbEggs
YsraO8+UWiESBoeaJl9vzrOLPuMkgRMp1M4p8jeqgLJbHGHbmBy4koXodzgnVn+b
gJn9y3Ep0esAT6Yvq02kLcuGbACHPO3xX0PwxeQizzVg4JnOD04Aa2UCS+yBGV1N
Imm8GXHOCTJs1Zi6NWD45rv0TlFscqsVlv/Tf9YPc3VomxIwj4Mc/1GLMUvvuB3f
1uIR5HJxeIVUoKzPDZBwlIIl4QawU3aGGtRrws4rHL7gMKrrPlV0MLExHlK8DAot
jJVVcXzmEHw+a9FYLtaAtdJ28eWcuc4Gd7CPc0tlYfObUCF/9zOA+m1agTQuDVdw
PUnTLwflzXi8sMxreUV4kxqyW3rzWr9rBSsP2NLYkV4Cm8hW+nUIG1/LuIR8StZW
MqnrsXdpd+dlWlaioaQ3zUlyDW06VEDP1IvlX2J2pGGN7bLezRVCTpuk/u2PCOAs
tFpztLH8f00JSHao9+0WJ1k98b4gSgeuSL1tbCiSA5eeXNMfnaCa8q/G3u05AMtJ
IdduUZPUfaYmJos9q2fSB8grB1AQ/XveGBbcvd6+mL+MnK0u5EXiuI++EGRwbH5v
qqccFBSxkPHOrq7yNHSpcxnfNqoa27PAs5las4YRbTnH+RUmog12JqWcOWWzGzgN
MI8ZUkd8OvnUsRAP6AAmi1Hih6CqiBKO59FzHpSBCMiNwcLMI8g5rPXz8Z1a5Ra5
MZgQfSVqN9CMVUs7KRIIUXycSOWZsLsSrlOVhPd93xCgd2nbNvUnUBEKrpt9uPMZ
yLd+cuuyw4VVhdSoyHzbKZfsbZ8m9TnvIZ82+WZB3aPN1Gf7or7RUyO6F91reRfd
/JM45Brf+9inbJkFwAJjknH10cmFHi4Yq/9FhZZI2XOj7mAWK8nlyhdrDDpFmHIS
zUTLCQ2dOev8c0XyDq5H2pKdPgPYWQfSZiy+Yh6zgwh6IxROMOHoccJJpcYNXKcu
r3EI2w7QgCWMKezPxf82o9pL7NTmSevctDQRJXhaHTNKk8uZAjyvhVtaWmeaQE0N
BwNoP/HfK4VfqW44s4QRxXiWHksa+YB5AuODz2n1X07TLj7b6JVgy6snlyi4KSup
HSyvsobx9JFEJctS4eCkbhZ6UmF4aOgWywnkPYotn1ye1eSQOr+HpEXaiqwskbcx
OiQ5ARBTewZ5xEw47A7KWzX3h17/RRTj52cpiXeOBRzBtfYALuPkRgpEhzTLNrGd
dfVF2D00OWhQGJG82m306fSyWLq+SQ09Gp6x8rRK4iOMVe2fOclt3FvW812bzp6e
TJVXGLUThByoWdFv2pk5p1NHU02IIyUAcsrHTj7zF7NgVx0TX0SHYy+31RiZ24Gg
ZKxaTV7ECJVjS+OMH/yWRRBnbHhUGRLAjxvL0oXmk/jYryCd+Eqlty89iD/1zusE
uGCjf0F1wxvScj403uXhtp8Q2FUVCu9elQpAWdhUxFdOam5nw3+XYKIExIKHpc+p
bMmUPI5WFC1/s9qAlM4sqFJfpMsY1m5llHA4CXk9TBKDrwHciVExrpZrXHQDVAOS
NbPC0vGpCajHLoGq1XYxbiXBkXg8Qr6dG7OIHgm/zBvRLBcnYaZfBRAq6c7L7zzs
/nWd1P2TWi4OfKAkMoQcoSY84axNxm6fo8Qd4NuK/BQMxnIbSRg0lej9x2lBFFvV
2Bu75pn/NkAeHIoPZvdqvrL7+6qhixXUfHyzgbYXlQEr+8lyXf+AJljfSZ80lKNg
QaMYOVnppuRJrdZPkY3U7am8epUOdioS33HLLSgzQm9J9EEkLCRkv5JOz1Jw3Ur0
tY9lvqu1w957EGu8jXnDYqrYvJnZ8TnQ8Crd91ztEyzH+mAJDIlLT0EAATcOb7kO
GMne5jEUB9zOOa6q/3tWRHb1hmv8uhLzRdDfQKSdFWAap7nNpha0jitSufyaGrx4
XlXwPNB8WjnqefmghGBgFrgqJzb2pWWqHDruiiCjQtaK5x50efsyL2DcthyQuRkK
N92/IffX4JxzhqWnVWPdCWhn3fgjc8Qin2ZE+QD5BdlckwSSkolCSImKQ44F35Xw
cA3w4AqAP5wZdXEOPaGYxOHmzHUNGX/NaEsDTSMSuKwuD9Ds595a0Q3PNcmbmTFa
YwiQKtcWql/0nMr807j9bhqrBLoJbw6KYfLo3611VNqL8CLt78iv2gRpTOoc1lbd
NiuZp6T//vOO6wp1jGw+AjCFPH/O3+YvdIbf4jlIJBHQVbdniereG/TyWKMrtNNj
ksLYvPQP3I6ywbQufd0kZIhQsic1zvJv0h8lFI5+bWuI5c3xJVs7lddz33GUzq9M
kA+nmCeOUyfD7Hp1B6RKx3T3kCRqU54gowYoRXQz0PDf2waZIk8v4mEY8ZMZvbmW
9UMC4pDYfwFqTNO7dFLaYb/kx5koG45o1yRAsjCFzosDtsdwCGn+jUNMY4hRXyWA
VtZ3RZ93Z5Cs93kW400OqNQtddCv/aOOxUcBKB3/HGkhTpK1e4Zmm6S6x9bMMQcP
fPZb2T1IIhrsLod/WHSKSU9sJU5nl2rmBnP5I64o9diBVoW+9ObIcWmiIwOpiOEQ
l3eOk+LVss1ZhP5RCPFKuaqVuvcjZzEFeR/IOEJFZxj8nZIX7cmQjfNFYrnl6mzM
NbzpVkQ0PMD4bsn5jJjHpdXyK7/0KHpp/mZoDK/yVH6y/+GWtVH2+2EhY1Ewv16l
YiBMIOdY3O0eaTJH8LPDgI9qksrEMh7ErgiHthLAcIKCGFOklAEkPQ4kvvKU4Svi
xENQXJuxBhhmM1NhGiqMrrrmmfaouFw6UVifvdS7bX9SJH1rudDwBEGFBgT5/lz5
Hhorq31E/QcOVmpUuoUjt+Zaa/5mW+baqBY9xinCOE2v3YoZXiH+nSFduv50ezGt
VERR36uL1QpKQ39q4Ks7+XYd58/xsrlPqd8uHbmwu7B+z6U/mry6yKRfcBZP+uzS
IWi2gzHIGsBq/N63ETwgr6DFGGGnRTapHUkWGwNqbkTQJFh9SaBNrdF9P+ZewE/J
nsJ93UiZFXtKi11knF68+lJEzEr2faLKopesr5D+HbameJ8P1LZ9RR/uoBs9JUtg
MzFoJwXsGrfzHYy0h+Y0iefn8IlhwGlZEgYESBHLj2TUuGxL5qBf1d5aTQdg4K9M
oSgM78erCs8gHrjmUGmmvcGb8ARyRkJkqkmDrRGbJnnL/OBwBa1t2B3xPsueEqnJ
O9h2GtRlCrMCQ3YTfavA/MMDdKNhmuVrNkYVEGW2iWGJQdamkO8hsEP2raWyixT1
5AT0KmMOvP91aIOwLi3eC3LdyQGVsFulfnpf/Xi1mFzBfTt271kLXZ7dBzUByEbd
/e67cDoZapaUgFCmj++hxcceJ2R1zgQuqZuAfZvA02LlVt0LmUbapyNrAw3zCbEz
nk3Hx6utJ1baGEuZIvrwHbqsc19vc6yHIrrNpBjignC37kHdeZz6nPc0V0+eTBvd
WJUj4NipclaKdxCNIuVujTYgt+tXz6ckmu8x4FHLBVtyDH9FgjdM/fQoQ6vj30xE
mulV8vExl2vhB81uR4q3NphlxNKyQ5QPJzp4P3YEEiE/VQyV0rsidWx3hw9PLmuI
oYJogZFypOVnDsw1Ix9DmAmdKIw90x6Zk9bSsSVD80fTsF94HmjUiSkN4G7B9Xvo
GZNbYcN4dIjqkvVEe9l8vQVwPP257KbKYPQDdNQz5uAPsEE3cuJw6SETeqQwiWx3
L3m8voTm/ov8F1h08K9n5odZ5+UowHcpkQAKj1R3pe79Rqamf9pql/wqCcB5/neG
8xlWuvUqLMxH0dm3umud/v7BES0EzLy5YOR/3+XWpruC5wAA4YHItRQeuNCzaxPa
Krdm0G5OpMIVjxZg/KlHueueDem1vVSrtUQ15ZcCmppIFXfvXxDC/mG/fsvJb4H6
To+3zW+x10igfVq3HR0zcGsBxiR/385GsjtlsAZF2Sbbmpes2Qq9J1guyfoJ1Ym2
uOxGs+9ofCavg7E0eOmW3O7jlmViMRARaIaOByZCDeEtaOFHaRoKBIdSuA7S4Ngt
PiZ4zljrxTzrnvs9cCInNlriovo6NbDc1dulXLdNcHQLTm66a+f3KVVI/hippCbL
C9evj5MViG/ZzjjVfpPnD4lPfDbkRl18Gv3v+/FWZGUwssj3CiSq6/c4wR8ydUtB
uZYumi2GmSvf/gyPtfgrFO5P/wKYu/wgg3c1gfeaoe6rCN+xC0g0PgJsBKLuW4MN
6JRKYl3uloxW8ELYWMQj/Nigy34j35kQyyORG5VmRuDvPjg9bobl+s8mZ6UiDZWF
P3XlQtJPv6bE9yYI2bK/HNZ43OqpxELcMMI3HdZHbMANtNQIMY9w72LtVn4ay/da
iloIP6kJjus4IpkzXiuPtcsMCcZpwlj2zmeQyxGggz0fw5bl/09lQ4MG5eBKL3xk
ZA82Toh/u9dHntn6IpheKMLqFHCSBv6iRYQmFNK76hLw7wfMxWR6We4sDMrfQIG4
GtLCtawFGadmh5FiNmpGiCNWEWo3rnLoDyjSrrl3thTVffzMeCozkZ0IEiWryHIt
Y+oYXppaKOT/6jI5/dxbfMjerJh0gkINfT5ofBQb7EyAnoOShGSyMmKDKK+eNcWK
HMHtGyP83kFe++M6t1rztwWk+gKmKb3dy7xI19uLanZ6+efLauybcUbnqWUUZc+L
ttiyaGCEx4NHoTo4JSo590KskK3P+7xOLe0w/KcVKvlS4ylN/4/nKVnrTKSOh1SH
7Ano8BOcWUYPsYxRTIjrFnG0k4MwjrYWVQhxo0aF3rcLr4nBDd2Bduqo73zN3C9U
p9B73k5Kuv3DjpfXux6r9n18iGJazE9CrYZdYDVNLjatoAbP7M+fiw7YnJ9k+B6s
M9G5bhM72G+3Em778Tzz0N3IHJfhjY/1nx+0FWROx0MxeOba1e6tKN3+kciJi/vW
PDMVyhsgJCfk+/watLu87gJgAyBh2N+TUGyRBrm6AX8x4YB8XL7xdoHL8NuXnmGE
csRxym4z6GjXOXwrk7OLO4STKDJQgljyKQZGy0ieclTSOzWwgdy8X9MSclJXNOGK
a5KBqupRkkVgK20Lje6VDYOwotewZoFUDqyED9+IZTB1c6qsBN/wQuM1DLB2uGnV
Wgj5Y7/9ctCtIkVR98Sau1JwxiiNAbmrFg5qiyq/1IrSASNa1eAoyVnKCMx8SX9L
O/+Ega0vr2ptK641hI5N0RsGxUyfxsVKn3LnDuVR5SmD7sNSZtfx2cCVVLpTu4/h
azUImEtl7Z2P3AWmkjc9wtNhow2Gv9LTr8fB5FY9IeiIgJdYreCmIXigxt4LA41V
RMQz2l1RAu5CLFpaGOz3M5MQB7VHiw7n1FUh5ncTupq1pB56aQsJm0981Tqt71Aq
Bki7glfu3c+HIspGrw43w3XT6tByN+xJglD1P0ciw9/MoxRmIu/bQEHT5ycEBsYD
LeDzLRAfJlCjjdUxplFyjcQ0Fai1S2C81hp5er4GtUQ6PNHMZLMDJX4qdbD7u6+/
GEe655QREoRNpezZBoKk3wIXlQzfITET4uW7N6XbiZLKDLTHakhgar2l78KH32kL
w3IaL8m4yYmXzXbcQkJBLodidOU5S01CEw4lTo9FKgKovrf+8wvV9H1p//eMldh+
8FlG0JqNsKVxthYfHBIrJY8yXdBb29pze1GH/XpjHs3y7lNEiR0nOm6HZeKp1x8n
bJ9sif0JcGkCN9PTEoFOmq4BjQZOj6mNeYDYL4K+utvoZf4Hi+xMrSKqXVUKRWgV
BWN2X9S9V/i1iUn6Ibnhjzx8hntWInuqMD8NKcWREfzFC/nK5Fp7plRfOoOPzcmV
WhcIUpVhQzJ6xsQFQ3OEmRRwBS9cW17GZJbOAmcbTe3HSIFmcOqvE6PaGvzMkX5U
SXMADb00zA0yyPHkRTI/DbevofyWRVMNass7uD1VollAFG3cyaCGI5OjmRXypjbl
PHzuWvzlNKWNooNp50fG5SLb0dUOXWVBbwp3hAL0Ht6LtBfkV1L6vqtJfVhzA/V/
hX2tKpKm7FHYGYMKW5e8faaOMcxo4zZTGa2HUId4XWATJU11yXYtgP98UW/ZGAA6
V4+4tpryG71ooGiRJ1au7YbQSOLLOEiq8v0j0HnAumYjNVBRInWBxID2DfFikFB0
2E003ad0/hlBwDgvoyrgiNrNqHUT34ZGIMrJUyn6ka8jBuVdiq56JwoRhz6zAR1L
s20MLXKmjXDX4dMf/yfOywUE837riKLaSBDe5ukU9APm0yH40bohuhyBI9UJTzx6
zygFJi+NHrFWqcb4F9FMrn9t7un6O5sjyNRbfeo4ErAJZL7/rpnHfpbqYbEw3IOx
7wDH/1/x/SEJ5Ki1fp+v0gk6b/n67JrIpqq1/d3k8V2AS/YBpiInYSVtREBC3mTi
oefzsUb9FZdepocThvvgg05wRPVDnFSJWVpK4cIQvDgq/GHVVuDYXsX/ulzd7zlI
YT0p1h/Y2NpqDzupIxVDadNiPlKWS+Ku0vcwYEAGQ3eDZpnuCzzENhz5+r5NWaRq
D3WBLBLk4cdptFZ3MQis1Xg23RB4ZByI7VOFkfoyBvQjVkyDJOJEIzwuu68dtwov
pW3U8u5yonyHeASkedU8IKvzaaPj8wdQv+SupI9CdTcQXvpNt7j18E4Pu9KnKXRt
O/TS7S6A93+GjaqcQb73Wvq4TdkIL0lKiEDRoALHl6lbapHMSj3lejAftKyU7gxC
PUkdIAjSD5LwI+Me1XUSW+vfiT9ORe2ha4FNZSUUefC9IfCJhbx8SIMYoqKChsra
dNNO43ORbgCI7DG369hO4G4+csFJpGflueBLuPXbvByKwSWKTUARwpNxczcW+5a1
hGiyfPZ0LRYkEX2Yd4dQiVWTc6snyCEXMzAQMTe6ZWC9+frvpTzMWGuYfwWRX36o
2PswW5nRDtOOex7tJeF6b9hJRgTxn4AEkuUiaB5hJ/DsZltdWnHwudO7m+pRqTJU
F7DrzUUtiBY2KJpS3708d70fLmOn5dIsYGvTdl+0ckzneL8ON8v8sc5rA1LbHm3v
8OwAxnx5LEVZdfx9WIAfbhi05eFIP+jWNO+tLj1+RwWFImESZhBuUpv31PbhneZB
tIxjtSHhraoU0Ca2eof6yWhZZPtrieE+jn0gaD1qKqaZvZrXA8NjnwTkYU3O8PR6
5wkthfQakTiNFdZlBZ+ae+MHI+eL/hkgTyyYow1/BzkLARpk3lqgeutrtZAFQSJu
DHyEA4SbifG9TpXE8eSTUeMfQJ6+77+N+B/n6lPh2nvCIVpD+C84mGA+kbsJbMw6
uvw8hTi6XSoDRt81GFzSbND7Ut/AcagDajPsQX4i53nK71IBSDD3lzPFfJxNqdFM
k0LLZ2suTxzJcSecXq9UuvIOYyIjLTz+v1jJaYO/tr92u9ePnyjpwzXUdDQqOwHs
0zB6vuQKcRxasWSBun1IcbfEDSspjnayfRnPIgMzsXD3/9NCYJvGj89GCkoB0N5w
OvPTY8pTmRPYodeDYoi6YhLsrg7sMtktJrJeiLn0JEkn8+kJJ+vN6R0RhgPrOiSs
wUGExfTxsGbXItVYhcCD+gff9MGNuxrN1FGAX6OpKZd89XXuqrpL2lfVAg+fwyC0
DeKhX+yZiWVHAxNVT3horPaLhxd+byrFJ7my8KMZ9NEZcjDrrX8ByCQ776s94Jqp
8A+4vLYAROLNg6MU8kZdZIOHLkI5Ii71cwpKIB071+OEawi0U/5xw6uDBFmQ1t9M
FUMQbQvlcjKiM0HGxFl36XIrfbUAUzlT3SuOQsZe/1eX9mT/VrxsjMMWsiBWCIu9
dLCf9F1lvU5rGkXHCId+hN7WRlkphp0yZFAuj2KCYF//7SkkprXtM4UvEF8DLvfK
F6hDgTmE1Yjiu+XBqaKArgY2f567kck9/Bj3be5nsHNTkLWMikyXRWJ3sRF3DR2o
X/SJ6K07Gcb5zzJ/Zv3o675j70xsCJzpXCNWQLRqvsAZofzHafeT3B0HKhrcAUhc
7RpQh/2ZdhZiQAqQCsc11OdLnOwxNHFhDsFva4/7YJ70SQ+zBDQtfO4DNbL6kFOk
EZ9oQlCOWjfYWKq/viURiZrmgNIbuAJcBbhO9+cwg4qmilGQ/q0eJH3UZCUxW3rn
aAK1kFkMJ7hJ+ek8auGS4fmDJ5XJo1aGIs14+QDj6nx/O1JjOzK9fAGjSOtE9Fow
8B1iuWH6dUch7sOun/Er7KzKHP0DoX53BLd4zC/yDZ97yDYTB9fN/iEvVjY1Nt20
bSrWGcRDL6/6zHhfadrxJBcDoODY2jLGF6ahBSep5OXx5Wm6ok7hMQ3S/r49zAhY
74eDpm0RLxyRnvJ6th8Ypq96CM1MsQDMwrOtAVwzQD0lsdWJN7c2hjLRkAhxFUgf
elJ7e+G9F4Q+ShRvSN947g8+n0hup45tCBKvxPetfpa9mNjI2Tu/ZrRR2Vy6INIb
epHo4HFG1l9AAWmJtwYoi18qKMs2agv0dAp4SrENOdhb2WlH6ha8YgqkHMYA0SWw
zdGRdzxv7MejGFdqdNmsLnmBL2RkUAFkQoWcEUILDa0S9r6sxpdyvg8oGtgvjZeq
ID7aPISqA4tfmT/h/QFaOiOQ0b4VEkp+KGedw4T3xmJgTxnC6vv4clAw7aV0t0dS
NIfbPNGgfmKXqBh/cUaxxI2edNNkINmZ/9gfhRVsIaRilo0aqig912tcWDUxC+gZ
clzC7TEn/RcmWUcrNLtu8DztpFjGRyAZ0H03iVazSmCxabnZ9ltYauugiMecXwmA
UoMidhXWNiWqTkPoUrKYpGaSY1zmueAf69675ZsQfSOSM3MsrsuygVRcY3RDvChR
WrpKRsHh6TkLpTDevBOBqK7ZiUADuElczTqxV1SlummK2EyvgtcbWrBuQTJ/GpIu
Bgmi/dYF6igMIiDDSWzo5V26jY8wuOPzwov4Pstvl0NRdkMgUmUlXDZyJUGyXjQ0
R4/4rHXA7D591AANfbJ+WPD2TJ8+Tw/fIZ6ddY4FtysigdERDiQzZ8PpDbnPSikq
/zBrZbpXPlqZw4tVugrnKRzlls8v0AiSHHGgOMnZUwxxzy3KgOzzS+L9dne7C+zT
/AskFYSaWFIgK4Ws/U9p6kU8EoDULvHN5t/QilJuDtvjPlFqu5VWyqdTnAB+VxyO
lcfWS8waXIBE2zn+kj5CUuw97e5d8udhsj3EaZG2r4d/fp8EpdRWSS/yqKbbiOLK
ke570fvlLSFmEPGwVsKTw1D7RuWy/JXMyZ7SH+R7AqxlBGaBwtcz6tOxfJicHlUR
CbWbdkgHuZLLCZL7DlFb392uSkriquQ5CyOX2uF7HxzMXAetLJexuL6a9lfdsdAU
d8xJRddpW7HhgAmXZxmw8vy6xc/nTVcqC3gO5PY+K12lraZ7w78cx0nbXiBPTn7T
9FdbtPvegy3RDEcRJUhnnEXaQWZX3bPgoDbr1IzXC2oiD0F6NNdI75jCNp6NZjC2
wzrVadTnm6dRCH4axmMY97cxpVig2le5cZ5/LFGKxpyq4VkL0ICiSmcpv9lo6XEM
UX9pOUhaaEzatqwVWc9+BGyKasyqweFIvXht0S6wwCcWhaY4155likDxXwp5DPXC
9Xl1uVVehD/izpV2ihef3vQ+y2mAuWmgTNHHay14mPo+bHjk3AlDSClA+62oyM2m
OugrxPtARwIcnInWxmzR5bIHychPR5UlMABgzD3uM4iNI6QKzsP7D6S6CDiuSTzQ
eFllzcDgiz1hPYsyEraeFuWrECSTMCLEoiRIAizLyor2AhpdzXpLU0ooS8kYPDRR
kZQL5IpmHEKEh6ia0F+svFRIFJarJTfqJiO1cdZxwY6mmRI2hfD/sHJwsW56gzVU
/tUOjmiab12HSamBCGDuGxDY4fuQeeDhnHp5P7crkA/W+q4a3JKg0uoXmfSGhJRi
9/BDgWcHOVqO+GKIlC+UUEWZ00/STKauDDnFrqsa9omcN9qPqQqKz8L/8pDfM1wM
WoKAA5Hs3TpYUCZyF2P3BL+WGQukcaWaXjK03SQXGSZ0cg9/8iMwSt9is1mPRL1Z
yy9Otaqfz9FEVOroAxY6BtQqrXxmAPq28b/L/c+U8hb9lk2C13HCaLFWl16zD+wH
EpPKI2O7MCYbjMnwSls9oyJ0xHv7EvdErTt6DnMcfzlCM5xbaeWaSJtXMowkeXKo
69T0WvJzg8fLCclXq8tTqxKn8eySdC6CPutksPfnrJFxMwowCLb1LkA7GaM6ISk4
kp1AiR9aWWWE80uCbZLQdnmV360R6O3tMPx4CgDCxcBOcAwyl6GPKPBtj8giyd/o
1bWnyhoYhKM01otir1k52GcNRc64IpQ+bzXG1LAphmdAXrCDwIyE0rm2iiy3uWJA
w3ERXl5shyEh4Wo2p2616ZJCJRnMgljzp9Sv3+7icpOI5PWgs48R1XWrw31Prum/
AqUGhe92aFSBx/WLiCgtX33qzCYyrRls35uYxgOAiddaRVMrw1E1K5CHEUD/Ej3O
SqQmxGPF43eQ0oOGCUrK7CqHOcaLSvbE6hUYqfKN/d02cgi1GPtN3A18BrXpfgS3
i6uB8Z6LTbfijhm8Syi+bDj14gHLxyJiroHqkdnND6P7Dfe68WbBArWmihJMTxrt
Q7675orNdnyKQ09X3YMZmyHuDhAblPTAg3rbfj3jfYV6Ur8w13twUm/0HkoE/PqC
4zxifmpXvuACMPJE4/QoL7aNKd/WB3kx7zVoBAq37IJypSNVlH/3kJ/Ke0RzHPax
pMTLr+4SfeG67oOGUD0MCSrWwBVhugXvMhzrMTI2Ct4oBFeUQ9kne5HLCi6g2ef9
SEPuYIC4UhiIuFYmpML1AucE7qavcfU40U1v/R69+X8Wx6HcPcYB5phGAjZkGox5
gI3ELxhL7CqRWJYpVbmbhyoYmCOO5sjJ0zJtEfuP3OUXMV4voOKZF9xGzKAjWvTG
SIvMN9Pqx0mtGPoo0Z7Onep8qQ7TiJAluXpjYqqL0mx4US8UdgfDnkeDqKoUUqdc
ZYsdKW+sUJDAc21EIHzcuMSs4RF7rGcif1kcXYpQvf1V9fjRt5QxP5KsKB07xA8Y
xn/hP0uvFlmNKQPQvITSyycmk4hyPpbaZbeIzmEGlOWGAcXqOWLG1dcZw6Vv0K8F
hEGyKRl1e7C9N3m+5TlQ63u5VVhph7G+1hdAHSULS5javXkX9l1FUcFM2gM0y71D
rAm/k5OJvwyTvyNkAxVcJJMOYJyS/RUWrDhuwZwR1KNQA/HxrAYwTHaKsTlikP6p
7s8JHWYl6s7RPhLHw7Bf32alpqgHCIq/SbWQduM0ZkNrIAWnBDgzR7tt855kykud
7EhEEb6mX6JzrzcRVuDY5ZsvHoSsffa790qc9LqCGwoGweQwdbT6Zb3BV8Fvn9NS
Qw6gVBLCA5pLh5YA5ReF2EQOuK0A3WgLqOevHTVtqPQ8jXDkhUYsCuS447Yc3pRb
ZpYA3+WFsoeWbRSka4nM4wWy496XtRZT0GtJK6hgWiREj8sVeX/+gJ8zWfT8CPvG
md4S4nt2TMz7L5ea3t/tBzqVeBBcPnlSHBUrCTF289RRXVBLoDedt7h6eaclWCff
d95DwDIbg9/Bep04JEuX0lxaeVlc5GS0PRsOAIslRdiHTSZk7jdkMMPLJlDgL92K
7FQR75pEVxcmh6m+aRjqHBlmzs0O/w87UmENRgyg87INpS2V+jOaf1aExFGbwa3U
cSvjZbuVBlUyaWOlqr7yyEjiYll7f/GMHAXDSjcI+LMAqLg960sAzUMgcguPlZRe
IcdJUygXoX5W4Q0LLOFMJ/wWAt2JqqzCrSXus3KH/jwcl18XKvHDA/j4WEHwxhFQ
x9jYmjS1/IX7eo6BGPfXV8wXoU+TY8oEnnmF2T9egB4d+VyXJ3FqexNR3M4bK9zc
vfP6mA7kXPwMHUNjfHx3SBv0S3+JMchEFQswAKJLsUU6khhshtMYzTlvckUzbW0J
SewvY5q4Ynxr/QHhvyHO89x4JYVoV9/7I77UzouIL2RvMbkwbDmmOlC7iu2pVXJO
6TTB8ZLZdtI9apQJ9jpbNRp6PBnH+8YIrz0XqOejJ91c93aDB0YJOi0qMgieIb/d
QBAi6JrE8KCIGr0QRMfGwnAo+E0HHhSS2dK5o7j2d05He04J8h1ntooamp+hZVbd
UdlIasGvF4f05NF6a3Vi3AT3dK5dhLt2gecDZ/MRNhPVOncbMFAWR0Ho2Z0u6szA
Es/cjP0ODPBORAGxS7ouF9X9hsn8vPgo4+R7+sBMki9XHEgC8IjvUAMXf2xuImx+
72aHfpwF099+c4q8hZOGbeCHWhVBFrETaChaNEDzFb6gEwbkltT+Cjs/pMswYZdT
0/L+kxVc6MEctumfxP2Xez/4aCkqmtvc7H50R9tu1aSI4OCzijmtmzu5DeimXyhy
yDTesB16aHXcKUoq7lpSLsMmuTpwQCg14VS9KAAvNdtwtSOQHg/OptJvWX2ZCe3U
oj3huQ4SrgXFku8egkghqTjEF4lkNcx6SIvWlxppShN6OC9LMMBQME2yhkIsMWke
+3cJnc1aT1GvMlqC/cQmMY4iVNg8GqYlQ98szyOasnTkqbZO4m9/kjuQaO8FoJqS
7eAIIPaFRc+gJMJhRMuHBIFlu7IX87O8AiAP+DhmQ3eM6uHbFuGiR+JeaZknLJ9G
xf5i/Y/qPHRN7aMbW7XmLErYfnTwyrLpTOMfO0U2ZN9eUKB0H+hB2LtRBaRGC1WC
1zLgQ3hQjzorYZxG4L6G8+yin4G/c7P4/5MOTKm1KpoucZu02r9jOqp6i9BKhEIG
V3muGzfC6pOvLvmQsABUgo0J5OdA7qTuni/xQv+RAA58a2Py8I8eBx4LkkHl9bVm
5AtEle3jLLekACXCJ4e9Wl8wv/pa3IbTavox5O2u4jRE85DZPqqXmAopoisljOwQ
F9S1fESQIAav8atDmQxP3CT3LW3M+qxEZd/pLhS4O1cwx8ZMOtTF5UdLrfWKFrYW
P/Qr1RBqM+hTb4S2vwtvYSZdpWOzf8V9MdsQ+4PaOT08JXSoBxtGsFjQ8Cdj6cvB
CzStFVis0ljPS88jTrA723x/3DsQKAu8MPWXOQNOkn8CCAwWEGWECOKGctOuAMAd
eh6+OnnAj6+grWH+yn+VRCT+2tjsCqjOmaUI9B9OPFLpRtF6qsUVvz599tBpOlyu
Cclw5TMyxGUoc77dEpkFF3gSxqddgj9BZOM4umgKQoSyeelwXBgS1N8+cUzZgIx0
qZO5j3+EjO9yGbq08fk0NsVYAXBjupae3kdbBObJMYwfJtE+QUsEX158V22uGYZp
lfzkNAR7dlA0wvOymRW5h7ZvUee/+jolHuhzpnopBmVvqJwAJYUKFJ+3M/+uJYJo
BTX2sgr8JQG776ZpzvdPjP7ohAoXhIWJtJLgSc0m1Giw5RgC2nLw9USjPO+MD7GQ
kXFgNV8lLNQTrkXPrwbJLSg1/H7afHT10dMftAUi/lEInJX9yTyG58aHBnygoloO
ZQMnbMscNlNz1/vq8ITeOydi8W2i4cHnDFefc/63xoEW/RO1z1nxsxSoRJXI2WvN
RzqmxpcZuwZmmDZxRnz0ByGKJuV6YLrmA2KVtY2IG/vCIF7NdzCIc9pQ0xS3pHMm
X8CYIxKLa25MCVOlxtQwdks882IWApN5K+N3n5QCsFCAuU08N3SEgAs7zFnq/1qp
qAenKqJm1Dw2gCVtc+3atanCsFxn90JDYevKmu/vYEZHzqgSthMrAdXoOCaeC19/
9Jf1b6FnheqX0XyQ7qISTx5ZTaUrxL9CfcFzRQX551hJhX044FuKi7FoZUQXoFxj
Dxe8v77gtd5/+CQJmz3YAUmrCTLZAmsQH/FY9ZUqbXN9kary8sXiofYvwxsboWBr
IVq9RL7KKVydsdk7hPGsxxoNMIKa8J6hAI3JXeNxq4vJGdv151uJXzKbv4BX9NNe
Y7lwFYXhvWvlKNJvVW5LiYC/iHLsQ02ASdGvjrXr3MdrrpExNMHUtuwRYk+ElK6o
m/B442TrcBu3OdkchuBJJH54jjC4PIG3TuCKL07aLVV7gX3GxmKdHakWZpBPp1T4
ovhL+4lmuc9S4ioyE1Ybrb12igjnRJarNDU5NJjzCyerbf89Lrw3SOqozUaUqUQP
kfwuE6t3NC+NQ5eY5P3tA524gM+CDwwpiro3/+CgvWM0LGPCS4gKreOxSONWmEly
7+iUWO4sXG6Us1eZyqBUus85eha/g7h83goVrUYVUcz81Q1Lx2IGOEjPeUsTDqHF
3A0h9N5gxFASpnV6wDtt2ZlcqjRgCVH6stlooef6UyMjJM5Go2H6S/U4yKUexVqw
LFNLgJ6etjY0e/vjLKxib8GuPvv97e6D051xJTx+i1b39Zkk2KV7Uqfu3u58BHcC
3t/ABqcsJdijnF4iYfavj9ngShd5C4RcLww66/Bw1X91PVJs51+h76eL+xzzjmrt
uqU1iD7S6Oo+quSqxByTXd5vvFpwy7rvr/U/ofKbHk1ztxc6h7zjvi7sXUAEVLUP
gSPp8rMnIVHIRcrh1TlU6WqZn1BjCY1eNTkeyRseMd9hiKERiIV9vEF9XPVMeMNs
IB0us1bMrmcTZM42515G7WmtZqzU3TtsaWBCMrLjkkhcbWcWfsbVmuyE+83p3oiM
j+FtT6Ig4qFLnkv0V0v4h2WQ4Nt3tT9W5xFyuLHTtfJw6FzhzB9lAsI8R30ftaDG
CvbHbli1L9D3MsnEVicpH49ynWr0+43dGFhVUdSbGG+Dg4Dl7ZuarpoHlYtdILWB
fGSSGdoYFceqm8E7MEfExo5bqxYBVS1bqRjd4cvLQD5QHyAybE5jB7ZX+ezQ0ccL
n91mqVZtQ9DYcj+0fuxeNOATFIJS8KD0uHSsUP6ua1Ts6IyW/k3Zg+sFYAVu/xM8
8/A+rezULI6DlHQui1LS6I0rivWATg0npSi+UP7p/ia3GGY+Q9rkhYE/fkwTpTK9
zhe4RT8jVsa+90D1VTtncsaaUceTWJtE8cakRqj8cjkzsdRNTdND4+ISckEE4iXi
2dYxC2KN9pcKaKuwz0qUO5TSKak46dq5X8Q2XdUvTAD6Ll1g51d+Ur5rIC93YEr8
Vxjhv4QBZKzvFsI9AJ7LF+In/hY2Y11sfcmnBaak/f673AprcQXDfqFp6yqkKjRE
BQ+Q0XMu2kPjzxeeXOQ/LddOnyQixUIAh8ng1QJDLneJdzO+cY2yJykQ6ls6wnyy
v/K6ER0MAZgNXpystjBiHtvjKEywyjUteo+Ky6zcBMZ8bM44icJRdBgQS0Y16lJe
aE+FoXTDN+KD/QFuOYREcRGpzfo9+UlUJJIc73klsGptR+3ZBt9obNy1WdamUXaY
QfII5p07cLNfTvcBx0Ii7WopAc8HRlap+yPLGpXZEqpIsXwZYWd9nXrcCi566T0U
xrxGWgaj7cO1zVxvDHtfw4/bxeBetafj3DuTgbEQz2qQRew5I4/OQkCKWQKPV4M5
2Nn6/INiByxhqPUDX04RPlm0yslUFwA4gqamIIg7XwD1UeEJbCcCeOEPzuMTjw2/
WvDInT+/ZwLXEMYVzI/HKqfrjjw72aX6P/DQqa3m+8UAL9FQ7eNNAWL/el3urY6R
qpIVc156a1v4BVivU/9G41iwnnDllQK6hGFunjmun5IJB7s5KE3WWb404NL6YHrE
Ve0pWDPdZKNmhtxrM7hYCJ/H3pGbSYldbnUIVKz6caf1k4lHcZ0N3ejQoiIp0aZv
9+d1Y5pFADNdP4Q0ykKsBmtaVC2eHwBbZlAKe0/DN9vjMteMXGQJSPWwwrzQ0jtE
+TBo6pomR8QXmF805LqTHcgJlcbLaMyUpytqLRDy7Z46U5xwtTucnQ6vDWDqaimI
b5e8rhpculD8DrtJvMlI/SeW58Kp2OJNBQqx4Ybu0QZR3yetinAPmratW+LqLg6V
wB56KaL3d2b2DIBQ6IYXOGA2Mt4/2ICv7GsClJ4A2j54UYs2TL3bo9H6lmLCHP8V
nQR8bvVf9qMP4ejnx6Zcbw+Wi5OcpMqFOlKyxbN67xIkukK0NH/tutiATnDP21v+
/sYo0t4CLFMH00FjBWVUZ9bRqqySgMIrFoqQjo418Ihfwo2YHBJFPCYU/fLPrSVr
MXQ8T6UDqR2EZwEQDw1RH+5Rub6SiGTpfXnIM21Tz2GpkK4cL6fGTy0ihl9+4luc
tzfxqRoktGapNT7GUtaL1av+Vn1P2pcAuUxYENQ20XUL/q4i0eCJUQX4I64occTF
OyhQtQmXFrPEB8BOEuHVatv0EJFQ61To03bjOCM11E1+F/1N3ouyGZemtgjk3xCK
dflf2Nikek/kCA6qCXU6E0c+6uzFmbiubzLIqIP3XR5j1fs8HmhkulXLHOnoAcX8
e03FluTI3afgKHRhzrIDQVtNOsZojIZa8SutzWQOeYeZB3eRw07cC25foOQZDdOd
S5hDoWjCwA/ttxfTGq3eMclz61jqVEpk++6jXrrVosVp9lHYn7qhjsZJVy05O/Yl
HPWXFLBudI0mnjHV+MMskGtE0lUocRmspDir+JA7kdcn8PiN5FDYh5WufJa9NFAg
31LW26G7lhcgBtoON0WoFXclbSdDrAr3WS2ihqVaiBAnw+iuCe80CRkJTLNwDYB/
5de5EICNPc5K1NgUinwVActpswFW7sF8l/ExEIpyG8chotaMa0Nklbe4THU+V890
MlERelgC035Lz3XH2MyinnTlt5+IQ4wIue/uzJmQcv4m3xRM0ydN3e7oXpWAqInK
n/WtY02w2ZF/+e5fOaVcVCemEI+dSdxOzDxJpAHiJw5HAwdnIbV4kZULYqWm4x6w
D589FCZRfn786uI5gocDroxxuQbvRG180P93XGQJJf7Uj91JA5ViK3R8CdL3iSIB
0ZLZn4hHXCjtL1sfApncT9pzE5Nr+jzphgHyFXQ9vlMpogGAV84jbTFAjT5bSuzU
SCxq6kRvDwv8PEESqkugzufPPw+sD1IzPozQmzKSR6vZBLuClKvEo42myxs+9eDY
TCZUr0bAjefmptgKUIxbeNN0x7LjCjk9OnRKi0xusnt5i0UgmQO3R9DC3P49s7pC
nvRTdvkbPUreVYLd2yQkUE5P1ZhbYA+RDXWLIYhFOgJiE341t8TBWpXPv9BDN9I+
U7/sskZ4AnMqEyc6NzBR8j55X3jQJCpTx3lZpf16JIxfy+v5poN8CQ9xe2vTYCrW
/QDOw4DcydYhjJkGoA3DBOQP+yFHeTQ8c0np3HJGhCui7FNRyHJv46ik3JDqQMq+
DXNyzov58GsXij8DQDkxAOLKx+S63z6F4FAYp+qpRn7qE3mt/yQuD9sziOj1NvAt
2BGeX1Kzy5m1HXYvpqwi/53diIr4FJ+ZQ/OP5cOzaClTJTJvlh9+FSX5pA87oIhX
kv56E98uRHMyFTom9zlWOzH3Tu7a2N1Ucsv8VSDhs0OIJWTbmkwYzmyRRKXpkc2K
iJEn7hdyHe4juc60uTfucidgIkysNhYwGOATs8WNj32Qg4C71Pdblz+Vd3PP4Pny
yDUy8JdLdpA/1nYHAIWztW+giWnJnBraNx67eGQIEQeWH7iVmogFWU65HDIyMIzS
Zyl7ejJxuWfwsBNrqTUpzL2HUXOHaTGgz50WAHMt468mIV+lKr861S3soCqmA4mn
Q792OGQue0daxISNJSK7CAmT5f+GFtgQ2f219zmfBDUanxLCqQtXzk9aA8j7whGM
4feDwqhSrRYonS9zpqLyxLl72XQQmo/o+/KxNQNCGL1tDptruW0gwgNHY5i8Fvxb
xt3okFlRDaNP0CWOt4OF2P/wys5fnew8wdVns56M2VWDeysnogtGvWk/xQp8rJoD
WpDKvzjD7gjhI6ww06H0cky+FztWH7plTERsc1FP6P5aCEa8tP1E6npBsMM6Y+3h
CZPujUdw1dXs7lBJsnO/4IztZn/boevxT5kHoHM60odYW94txlLLafnV1WMuvhfS
ZwsL9fj2oqjgrxdmeJ1Hrex7YxetkN3wHn37Q+uRfxmjj0Xb/Ph04Z6S/gMvN0RW
Tf0IsyrEm/qp67MqWbVmW9N10KxoW79su0lvKoWBdtvCTCBI87rdNXLJzK9ECcBA
hhzsI3cGTM2/HWO98kEnZFq5MzV2JGjpYmJJnlawWiVRyldy3HDDtWbS9xJ2tS9y
tI13QEm956GokozhHx5GfhxFchOQlXLqqnOm3N09r1FxTnzSbysrkpwT0Up1cW/I
LQNlt3gKD8cSlfCT5DMn5hukIoJRpO1NvXKAclrhtyo2A9+C8J+tJbC90npYWLjm
5uG41IubwDlpOAme31kprxkavLLFMeUETuYkIK/ElaolsBct1bsVjenLT4KjpNJs
OIcFYYyQ+5Yn65qhEQbAdz+J5tXztaJTsM5SUEgbS0hDY7Sc6WHzUagebtAuFauW
SkeBdFb7quJj4qXFFFghhneGuBdSRBecq9B0Pf9EhO0ZiuPPHCtZZUKuNxL1e46q
DWA9Dk8jn/bzpmWq/wNx16Uoy9zsdXZcCT1rQV1F2jm88Itet7XhbbHI4ppu3RzO
J9AQKnTtdIIaE5ybI5w03imtxMDElgv24/qCC3clVRZ9wF6BpVJSkRWXLzCR6hYs
GLiLuf1IazcunonmgKX8d3WHDshg87VxVVok+QhVQWRNbwoLOCnjaWZAXLdWoNXq
9dgo/wfsnanmNZRhs7HBKgdIOalXiqZfgmODWp+fK4fgZXWB8g+W1SIFbvCxEsaX
CforH5Jm+icvIx/meNUrGMX8931DRxu0fxMkC0mWF671REy/0jClhOw2Ok8fs50p
MUlpW0VWJqGGKP4ikW9RaR1hhHYkTK2z2dWrdyLQaLfhokSkOcLrS7tosn4jc1R1
odXk2UOPlUEgDKN1DRtoRtgz0l+bJxWc+SZD/D/ax/DrTmohia9TOQoABvA6//UV
HoRakcDFFHaGyLhvaSBEcKEaruBr89Q0bbEkbwcPMbQkeUqplVnzmaEub3XpNBNq
COJuLVejyUhvF8G5n9m3GLBT1DCWSGBTDrtMiMYbfKaJZJiRnnepo8oeduHzBxX1
/W+HQDwpfYLPWQLkYb7V1juv02ecHP0+xAg/Nd5L0eIflYdLxyCo/BF06WeXXl6h
GT/qcj1LxgE8TMruBr562q7lT+xTyJEpFz1OE21K3hgAp70sywnZqN6VaQHqoSnm
KNj9G6w0mKPdauB++r+w6ekb0+A2P8PJiuM4l0Hp2o65gSnXSmvfdQye0o8KOU2H
c1HW59wUFeQxjh3HHB9jthejeg0nYmf5xt4bfeFlnCE+Ewvxz5bB+MpVEjpMhAot
6oe8omfrNWuFzT7jnD02uwtiQYej+h7vfJImgFE6JG8ufTXuXkWZEnUapo2OBQKa
BsNqKnPJnl7pz46IGrn6CP7Tt23TR5UIbdYqK3LzyZ2QJov0DUCNzaXEuhtCNT9r
CAXL1edxng81CqIG6gZrbCwN09t4ukiw6YrG7SLhVI6r5kcq+95uPf95CF0fKcVk
gADprx3SMM/vLIgmA6ZWXVY6Yc1A/fzcfonPj2eP5OHYbjDBdxlELyKJYKlWymc8
UszMuu9y47GtJJX9V6KFi8AkcbIzWzdNMsacqprXTgbUBWNyAWaZQP79+xmxVHEp
v1gNdbOxDQY63pcEV3OLrVQ45OwE7On3/ffnBKnjeBDHNSSKOoLTFFCzs+fIRTrw
HDi2za2Tu56OcCMh8CV1ERejWmtCtd5LWgtjMYKdgmhKXGDCm8PF0zdSRjKQXkiQ
inbOWqmqALk6gjuh+xPG77gK2GZ5UNGfW4W6CcGezB1Xi7vWSFmOPQQgdr16xdEV
3xaYxdQMs0nrCvmbC8kU0zcMKKS9GSemgvvC0dG1oi0ajiR9cz16Td3pwzkR8QGr
vzWscnPtKcSt7xjM3ezIAQxI8K9D/E030YPzXoHxkPZtglCgenjvEhV/xvaegqxP
Te98zCK6EJtkmmQZW8nuMzArXme8EvO79lIKIcL+SV1u0hs6rPaBm/EU48HtKWvH
5hPiAqEXJrYpvm3oAaoNy9TEfO9nTjPN+rBjoxwyAaB0e+maadjtId6MjBn5NXdt
qUvnYwZ5GJRrJk/xYpiWTZh9MRTRL1+2FzpC/+dUuXmFdfaAqMvYwvvkIBWEfPBh
Ja3rn0rMbUKlmHqwI0FSXZhZuIOJL/ZKDQNlXi+M348rkpw+kuUQlPZusBaGZUD5
25JGkddeThLfAKKysyDwPwYgm7ZfKBGchbRb1/3LGhP8Zb9m4nfiSJ/0JH1jbIBl
Gc1V3UHGAMbcRlNOejVIGLXwgOobbCdlwCq/Z6CoHp4SgPTSusjd1ebWcuSFTMBV
tGIfcR26NmvXAflb+tdqV2KRrJSjuWHcNPGuPmD/SQ6NyJQohZv8iUDmNDZDMSfy
6cOwCgdJ/OVKbz2I9ZasVqE7VOM3j5uyOVvOddMHAXaRXhoQDcH7jUBq1oyVLFZK
ET29rrBUWfTzK7lrYhpMnBNx0sOSDRGxK7NhlGVULotyQk9zv6aN9gdkQwUhoSGw
WXR7zV5725qiy40yPnrV+oeunXbPX+hol/q4UlUZ50yD23Ji/b+U5OoZfR1AeaFk
r1Tu55ab3uqVfD8pyk4jPQHHo6rj5pW4vR2oi+MLJjbokiUa9H3R6eXsMR41lVe6
KBPaDj3l6HrEJhZ7T6npHkZ1iX7wc2CB7WfeFUuqkOBrXDhhn1U9MbT3ljqxtsIv
DlZNEsCQJ3AlGEyZU4MSVkeGyz+yU2i9kkrAPufuT39RjyDq7Sl1AOE4s8kTQqUy
VazCUgtWg/yUQsmwux740ORC9xeVtRBesaeyEo4blLAxoip6TFZCXIqZzft2iTjt
3PVTykgunT+/fFX6ggu2aZT1qYvRE5Fhq2kyCPqpnCx3JlXCbuNwLxb+skBHT5DE
hj5r+c4JJ/trd16U1ybVcHgyT3SmoXWQFmj1vPFU2NIxOJdiar4urLZcZ/VHw7HA
r5YJu7vV1DsQmytvbnCCpR/ErsWzfsHDTzDO+mR/KmsFJyKVuWiHjRJLXbomqRre
2yn9zU7Jv1v16V+LtlirTNPJoINaOm4J855XXV4rmvNBemD9EJ+BagsIs50hFaL4
yDO+dAME/SV+BcFwmsf+dWjlK6alwkCsRVPl7jTJOvi1uz5mom5vEhN4T/ej55S9
uPLybjTfShYOXUYKH/v2U522D0oF9W8NdP1RFKHQnu6RqwYcW2ISJuxkm870+Lf6
9n8kCV5YvpMZg6PDl7j8hEYW5CqenZSzDjtvDEGO5ZjWDOgET9XCfntcbSHzkYm5
Wk4bpdZpkaYRevY1fCYp1CDEmpiQR4NcdubtTRa7rOxX2DJ1oRS5XNsJhjCmR82e
r13GfJVWLYnjmyWFR9YBfdx03inYx2HRsdgoDtRlNK0Dx0qJH6/Yaxy7dBrpI7t+
9uNk1zQRF9k1DljazM8KdT/Usz/tk5NqbOS9zhsR/HlTBWIHypo2+Ji6Upq8RbdP
BvFJZcpsSoLyOOjWmmIn3OSfYhjGQ2V5tRUEufRuaQ6B6ibyY4QM9wMH1vzxIluV
Gi/ODfeOEmD0Hfw/UbXzhbKEQlG/gb4xbmvLph44yI2ErhZIXPXumQ2im4nYBJ17
Ej/PmO+mCm/f0QYxC5T9JFor1FvcEatHVD/LyhcTPSkJFE6nQNzKOFhavJ5tDHys
0HkPug0cPqMnSNpJGUHdQvuKK3fPo6oFHXE7njBp2SPWKIwN1hW7FNDxKKmHYuil
62nSpQmkZOv9XTY9EJSr1qZ2246kgWvjG2DEynHGLAf2NBksttnT2R4t8S6PLF39
53GwLBlEV5GBvw58jhushuD6G10rZQPSadK3Ijh2fEwlTuur/UyCewSf6pszHvCd
g2qPQp3vLvCKR0+hwnQupKK5ExESM9M7pl2+PvdkFYdJq2xml3Ef/yCrTFeTzaWl
QOoJ2akYIpcoVbQI2dLGsi2+eypvIDiJOSgIwIjN3PFaZyKNLyNhxuDofomgyC0m
pmRfUeLnyNnsVcuofMUTDIYMC+K9zp+IMcfBz4EUqPyujK+YumE+QRyfykkHlUs+
mTmgI6XI//ZbJqGaeMl7SvCj4z+/VmTVoP0uG5ZT21/Mxif+F28neFl0Fi88Up47
io2TROpKTJOCrzwuH/iDEVZPLyLZ08xSqMNkgf1C/TNp+xe1ANRhP67S+rXBtepv
izHiz4pN0alPHgvp4VJ9kFwPzNr3CuTRaR9QBz88kS8MeJGAu8qxvHNtKpwxooPi
spj1WLL4dbuKbePNxsyZjOC/PYv773zlJZQ/mpOV3DfSphTBn3lp7t6qisKel7V+
CAl0AaGKbB4wWdAsqnD+lEO/XWI5rUHwVb5Mx82QX2p+rPlSumT+nrD4PnAF7IQm
avludVlEM4+BhQ9s7sWfEs6gqZEupt6PVvRuoCy9I+HeOiWk9fiLbjZ+2cNSE1DJ
XNc8rWbh+9B7rlVfWLjBZr0UEnQ7m+wq28vz0UV6bCAtdRFrb/16OsAVtBH3+C6b
gdYHQ0kZgG1dql1thEGjhXDn2GgLcL9ZG/kQDiDIVP3P7oZmxSlU+CSMDZNCpaf/
YJwKatT68SEb7vrAltXrnOFy18nlJagkiRLV1u/3yDA3+/U2NF/7Dtck+Cq9T20c
59d2p5EBkGJZk8FFLUbgxRwSuHYhK7cOLtOZSV6UndMax5+SsrKllAD8wlVyOa/x
CxYQDNd3512HVf+oB2oWhW+W4mSVIu0kk/fWl046BtSoBPJ/TUmGHwB3NJD+76lb
Tz8wPTsFz4AmyVsiV0jL1ePJMx0KWr7mzgBxpeZ1Kn3J+DHXSnGWp9NQ43d48HCt
isrDN0XyLdoYdIjyr6K1WorBEQ5RKwA3fv06YZsHo250mVDjfA+kztQbEVwISNc1
SXP/fRKho/nmO/hXMSv6zu/YY1/sDtGntn8dEn0bKDEMQQLkJBKCzikUs9nZOvhV
u0yZwUzjS/yDuBpoAVJZ758Ob/1MOfbzv0dg7UZvjcgat+JvjpIKG6aJ45CN0ivU
3/WkGQeW7Usp3Xhpjf483s5Y1zhShuD1+1ulONUGH9CUO3kiqqKnnfHBI7eMX8j/
30rCDECx0nMoHAHBEPXr5N1XW6pymfoUOkUNNCOymBInclq7qy5OqXuGFU6aHAX2
+wiFcbk5Q41sjW3V91vQUO1ZWuzpI1h02uHkK68nLzjE6SqIveVaduY5NTx1zgLa
c6wH1moX+NPZQvtjnDjyRBdKhPvkRUsy3SrwOv6qQ7+/3Zrvrragieo+4mXTbVgN
CjA51paGse55w8jbk++q3omyb7JvkNJ10/BCN6xQwW3ujF8PCdYMDVnlUfCHC4BU
uJNsiQeQDR+CsgaBgkI9QRhJUk0G46uQ1qvywVggi7kXtE6SBM+1aLOWWC9GLCrb
X8uo1frbuqWeAPCguLag51ZpjWa3L463904A9oXxOD/lKTm6AtIVMO8+lJRhYOUJ
yRVI6VPA0RhzVEgshsyG7sw0SSiXZ5rduzt4YTAN3WDDRchoj3A6KQiDUhaVXgmO
9RNsHRpCtqPaLFxkz760BFkO/aBUQ6WCnmpfFAPH+x5PC13pzXBrlFTm+3akkqDe
B7SbfdTCcyVSX9dv69NhQ6s5QgEFmO8tQs5uO5D6iSJINPcVq7ON9FE0m8twoHz1
935NFUg9MVnEmFyOI123wgcZL2J7WnWUWJakxisAzT9lJmBqyZi7bia+7/1DTyQg
PcmGGg8rL0CbGcS+iaom1e9MxbzkryMFfi7QXG85kkPbCmiyvi3FcolK6dEBc43U
UpyELeJ9Sp1SnpqJf2V9J8NSkI+YB8ZYETKOelNyMQo8LiCuf7FSWYHTFzCTO+Rd
HRy/WkOkI7u3ScsDXqUQ5ejn+QJUjZWQhV3ncRdsZqTpjwrBu0QSXeEEB+6z0hbU
saO2qHo/LZEbqZdJUdNMChWDqOh6cBXhTr/y9iPmEc9evQDOe5B9CkSAUiPLzZFQ
dIlxAELbvvaeXx2FLI5DrnSpLNCiORDUw5lTzwUvE/Yvm9JHVgQuCgjWBpZgrxbK
R5g0/uBz1wuk9xAFivDecytghveCNbYomY6EL8MuSjDCNSo0cMtQRQ9vhyCdeX2o
5jXIE4GD3XrzDBlCwlfXPxjKiTuEj/lBRr9aIwCmRDbntpkf3W1oY4MlheR7Uu4G
iY/foHto9m/HeE4iWNH0X/qmXCi7XXor9rqOqTULKZDYMC2IgCRRG9LaJUDa9Z5P
x9hIMRw1FMwDEMEtA+mo2O8bQi162MWn4quqndLxq3C+PSXZWLkdqGUe+wdDO68t
PbjrPaPq3Z3ynHRBstjAm62HfZ4Dxkw1VMgalBobyZRqcGnWZ2x+rhrTEQAgva/k
fNGT+abDri0cN8gJk+Dxg0T8BD6Au9ZU2+GtvjgSp47QfJrg7FD4pU/+pxGQdxXy
Wn7/K4Ifcc1k2rIp68XtQ9H3u+b3u4vDoUm3Vy9/atcm/s7IJC2/67/HxMll6vQ2
9rPxPb83FOLh3mld7ES/mdWUnw7ILYHnky0bMJWfUC+jcatXmjJwEwOPVRmtS66E
mYNaMXOBW+WdvN3J5NlgcCGk9v3LcoDNyB1FzhxWxQnFVUoGibi2kNWMySZXSmT3
6K9MvW6boHe1uR3JeNmc0yJ0dDYacKGOcM7TVDQf7Wpp/M/ktfPFwV81eGziqPyB
+TiPhRFRZtBKETav1Kix1mY+gdviHQHjz54TiRy7vIs082mSLt8113zulaEdkZ6S
rY1zxvK1HNiVSR76XYz8sgd7XErg1UjwZ33iR+yO4MxkXNReIiXlTipOopqMb8S/
hMMjZEoT0yWSOGhZWqGpRCOwrsBagVNOP/vO/d+NiFh1TUm7mEMGUfvSyE6wG9aQ
emEsiAp0cJjbUjDywqvyWBbaEn9wyGtHP7u/ay1hvf/R8KSV/Hclf6AYzNhd8SqY
rHpjODVqdTIRmajwfXsAmSSY9s7PIfoWWq3zgPdCJYqa7YxCYGI9siv8FxqYDCh4
NIpGBd+xy3FOta5rZia/UOnktloui9BLwukBY45EkMWdrV2jpfXr3yH0PKQ2C6Py
Z2JCrklRKwd/ym1YDyxpw4ctMe6oLhQYTt7E5nM+Q58meA/Mu+mQwjiS7OFI4sp1
EpHA0tsd/kHXuBlubXg6034eCNCfrfxZP45hns/xmEgD+d0w2+c/a1mTYRwrgsl6
nqe9x8YSt2smJBBNyHvl1YajjamnXzj4hnYookSBPPokR/R0erVhW6oYv7+r8cCU
V3KKkQAzWgcvAAdTGteNRu7hVGZkEbYpDsDXtaoM5jdzdkDXv/w4CCrdbUKCjU8N
oSuCDIkkLkkvYuBOXme05Vj9Sw9Tst0kqDseoBPI0l5Uqpa8uUeNluHmdrEMCLEm
u3RHUR5vtwupDO6Lo524+JE5i/XZ3UwONMYT6fXPQVEEGod6kinV8aCk4ZG6mPKd
q9SG6ddTLHja0/YjSgNUKdavkgVNwwd/3LwfHKXglzmDxbzB5kPjX+9B7LeYb8UX
BU+jS32b9V6JcyiM8kEhsZsBsB/PWJHK9O613MJw76VSdSSIE2Z4l/2rwzCMiB6b
uRn1oPdiMDGvq2J+Jf5SIPMPSNrBUs7FwmrvA9Cyt/qEN1lBMrwDk5swsXbshLtT
OB1jxKtCoX81got6fGhRofvMeNGitXqCR0W1/GKUutR/3evXdW2HuIjOOtCNuckS
bx4whEqAwEaDsKphh87D8OcAizJ2xt9xxiZd6LM1aSCsiHcARSMMH7Xjl2/4l1dK
dYbGcT8KaSInKA32KcvDLMQptO2upemZ7MfxWroz0Dzgfxdgv57Frva5t0oxmcyC
TSXmB8dbFP4it3FES4WIzebZga4I04FjN6IlH2WtPPbW6xhjI9M1YFjuv2NI5BCt
988rmdDDbXVLdisxdALIY1g2nmjcKF0yLtgLNC3EDZnRmeZ+elAQbviUKindyzmY
enW+c1dyCm8La4/BJ101t5fq1dpnp83D0peI9YOqVp7bSdbRnlJeocvN7uc8gxc3
1IGZunVMYeAx35Zec6HSQ/tbm0XwUU4/ZAKwuzC/TE73lfqe5b+rNQ6KGmF7GaiI
8+Q2OLVYcWd7yV/JQpmmlhCBxmgi0aPcNO3uf6Zzq03tE1nFyGmx88Kvh6yOiMv5
mF1lXrGZDfPjqZEa/g4ho5YYilRdgpgKE1J6DQWZ3nwYzhMcgWc65RE4tZpSVDGE
fEARRH6JlCJq9KuQEC6IUrFlYF3el2y2/7N/87Yk9Ma9qJkCO4OYAF+iDjdzL44s
W/RD58gFHL3uGMoBgf6o2mPO5LANG27cxnRvNKvRxwfLLVgEzqakorp3eQ+yfKJr
laafVQv2bXorq2Qg0st+kNZ3Kttzb4B19TVhUh597nnVdmAWTdLcKitOycNBs4/g
SYXV1MbuFCvfl3pKF/S7XFLnj8BRKPm+UdPHaQ8bgXE1sbxxIODM6jIWaJZRhFVF
jaqOWfaDTSZRLMl9qrRvXZ98hm6w/sqX6Vqzy7pI3bSgieIoiZUHGHq4aEssBzas
zzP8sZD8UaDl1yReN2C7M+lTM0f7g6AyjAc1u9TEHIZELDYz/sa9QqnanIoHUvVg
qFvuap344io3f3j5YTPf66hOPhRtMO1bX09mHq40iFBFkZoOGGrO4JVuxjf+ZddO
uUAFCY36DT8jHROEW+ZXHm9byZcTuS9mFhrVsSmU+2NhJi1Z9KimMnOfDWC3INSA
bVEL9LusPbn+EhLmsmmQ6RfFc1/FOb1XbHHW0RVCMYx+9hJulVTbIH2xOtA2xy4K
KVy2P1r8UEdMPh94PGX9ZUI2VViMPGxkKbqjNUun8vE5NWBTRz5uoYP2u93XZMQ5
OEe0zlRxotvTVAFEPMdr6C7AJBWq13ShbPi0BWEQRbxv6SGftTtteCINAAWRBBLG
br3nBQpqQ0x0rSn0mrZhCV5BBsCGlgJ83HxRUfcH478Dox6Vj7g635lbn22quruc
b5jaGphydYfC6Cl9/r39Lqpx67Tp72F64kaMkQjYXeJysopfzn5imGCAxxzWBxe0
yWIkefd9JbMDWCJcpN7l8qRBQ2+nrK6NhTIoJJWIUNh6x5Uiv77uQVTD2UTdshGU
D2U5PsKGMEIMCMt061cq8K7dxH1GRg/pRmHcaW2QRRo1qymTvyWP25lhFmnRi1bJ
HlUmkj1DyiXOek0T+6BBGjV5A5x0vePTNRTDCeLsdy0HDFlxXfsKM0SEQzfDX15D
ptEWyT9makWqWyBv3PdEAcXxXPlow/Rjv8RlhqNhLxXZ+O5xia79TnwVfN0cIzqt
PsS7rVNI2IhaBLeMlzI5cubmOL9gpLtMLnt67cySFhuzlzS5/8GnPI9jUojCPQhB
/sVI+PiWXBhbyp+iZCyDC5xDi/gbXEVa954UOVMBYXSStlUIJfF2X3encr5o6Dhp
EzB7QzHyTV3MgJAt8XiIhDdbSHxUe7srGVq7IEa6QbpMNCyhNtuUB8RTLzYw+ut4
PNgHrEFqHjxmGnm8nheQbGY2iPrhM1kXGXomlrtPqXNreEE+9r2gGaGNRcq5S/Nc
CaOUqaz4o6RUllnISmrxuifFdC0492mySL2uDqL7iFFgb+tsDqdKOrfeYzbuA/bB
kb0ISHzIeQ3AmRu3FsIYgoPnELt+9GiyAL3xDRvNdMvlmbaqOnMXUbw+U+G430He
xyOVCPWBBifnPHt2BZ9n2qcaelrVvIeYw915XDrT2azVmR0Br6CmB1hFioioEBqm
7ytM8Uwv6jVULyssdP7MEGNXS/DhyBpFmWFGyyFF1tJMgBCUx7MelSKU36dQG0Uf
1pEYKgHIPWoTQ4mc8IIHtSrhwZ/gOPihxagxpIWhzwqwBxYbN8K7rqHaOtztQdHj
Z1egbzn8kvgdo8tYc0zKjzt6emTkWrih3c9WkzdBWt6WQypYHIfHN1oRqS1pummB
T1kOQ28F0KL1ADW/P71MFr3B/6bR4p4te7sfEV8eQccpEtC/a3A9n9N8fcKLoBik
ujI/EmG48JRF9qZvgwn5IS1AjN7ETWiK4bTpo0LASGkqTmhKluY2c1bVq7JxIoTt
B58mKAM++9ka4wKvVKkG6B/7c/yYdkYxa5PItmcidiUylwv7rx0hiHToZWcmTT80
TypCegn7nsrX6Pc/QYZa8i3WFoYu/kjNg5QJQc0wMA2Ba6dzzfR5955kjKRzBBKK
9yPAKGAsD8qGMe4pp0dv6oYiHHxMFfYMw0702CNxL+DsqV/0fVLKTq6vpDdPPyhM
UwP2Fe2dEc24ZeN+MsEM14AkCOVMZyp6v5FbKxm0MkF04D7q5Yl2MHScu3gaPwpx
Szb1V93qXIMwcaRzlWv9A7sGYPeMGG7graOcB3v7k6PJ7r6XxZJMw9TUPM8nTW4s
mTok+I3758mM6USq+VLvJT1XHBXSoCENh8F1EXn+w0ncXhV13Ken92OHKXtZ3F+Q
6XssOr2E4QlUZDN+JvKGyEGQq7Ie8OuV/jKKohuvluu42o+SYHo7CvqMThoUTodm
Snf02Cmex13jQeZ/zn1GorIHa4othV8JN3kGHO7U9Km289ZhI0o/Ra2XU0NcWrKc
whdW7wbSbDQM7GszWhoI0gGQZSuY3HG1Jde5yjR2QPnBAHA95H1T7YSWayXcQ5oI
JsMKqrwFW5ehITu71dMyf73P/e+TlFEosSaAMl5wWtNiB2lL4LPAdjRHOHlkUUU+
3e0JC+Pt8JWA6gEAunqXfHNmV5FFmXxbozF8BOr9MaedUNuzQUp+t99+BgRaSCzr
jIZRhFmX0ThW44QVv4Ux1bVYxk74TnbKeZVaKX5RcPVVXx9O4L7DYOwkvhopnDmK
fC4AQNfB1Ru3EyA6V1QQfxPeJennFlYF+4C7LS42qODErwb4jsd6QudaXTinG0bX
WYrM2UYT2IibqcwvswKWAzKCJLLLalvG6HBbInNC5AQrVCgIiIl9rw98NhejUflM
YfgcqFW4QDuQjf3AVy/6jV3b/UHHZYMMT5y6vwV9atW5+4Lj4uvppxZPcHmwDkVU
9UCVpLUgpL5DLVzZGMmV6Wf8j8NjybozgrDhU6Q7EmgElm5PYclHguWhUmMKjUyI
W8Oo+XqTPBtFNhq2+Xgj9GY9vigPWCZqnnC1NekWebuo6w3p2EFGPakKyvCghYH8
j91I0ehf1NbovM+ZxepLCl1kCebrZipwF9XspPHmOwIWnmCrGJJdJwGrkgc2Rx99
VnvVyrbdsk5SbERxR+B84Bd9i1Pg3iFbDSDdFJUHVIdCVB0bE9Q8M16clFneiE6t
pHWnYOlx32sF6p4QGxi2JGiKVh9R3YhgXGCgp9WGmFcoUBhFF4CwgCZ2SBIEVzrC
ETvKuXXONZFV8Ynb6e85CmEbmthwCv/09acGvZBejsLqFLIFwQXdAvuBNn+rP3aI
X9DGBkKP7Mc3twoXo7CwwCCFyenTTivGtZpcAUq/3lP4JK3AR6YdwS8TKzWBbPh1
sZBDPbUR0CUD/bhgIBOjelRCrnMtKEmXgZhGf5W3J2mdVCAELQJ1oqbwj0AC3FpF
Xlu5VsZ7pQ+8/IRvuXN0MdDTmye5nTwyPRt80PEbkFr6ruMLUf8JqjYYPEcwbVai
PCv0asas1exiiAzTE9X8hwSJszY1WMckntM5/HTkTJOPW7CbqLgMQsHlyUrHq+1d
gojTJsuOI+EO7YjJSq3fNeVg2wtK+mCk18fc7bxTyhoiF12p2B619sCjTK/3+iyA
0DxRHCXIPmUV1u6DSLC79G+ezIG7IcsZqd3Ui3bc1MmibIfrDhVLWdXzXcB8XldX
Fitj/v2iasqHooeVbEvyzR6wC+V2bWbVtCXmfSj2NLgGjENznN/LkjNHcBq7n//Q
j4LDNsFyv63zvc3rP/dzH9c5Mo7X0ATO1Xjt8MjJoBqJxRH0UNj7A8QkdoN16Z2V
Z+HWj/5bseAaZ9aMHUctTBsNJoeVfecGWyQhDIuR97DmW99ZRVS11eH0pi3dJKhR
D6Xfcf+9BXJwwsKRcyD7hzxI/UZqNkSp0Os11GoWUxqSa/Nl3c+ai4mZugSu9ElC
L2h29Q588AgWtpWFfmmPahTu3JEp3lsTr2pIKXKuWCbszThcSbotrfMRlK+Ulaq1
kIRt/6STNMAxgSgk1yN+tShtX4FzjA409Urz7sYTdFeFiF4+B/ttCWZ8UsdnkN1l
6OpR+TrdQLthPPynl/rmLn0I9wtIi7URVSPBTWGziWTZLlDCbFfggHIrq/X48LVo
WyFb5EL8NZnN7aEC+rk96IdHElk+vYGgJgB92dwWx3xxxl+nPioEk9hla2lRDD69
huLbjiX/v/alEM/Kjls+I3UpQDKmjl+Qcw9p3uN0eS25UsbACTygG6wYVVaNUYPi
xplkLoXpSmrA8lJ9FvMAhj+LBPP9nJIiaoWoYQHFYQij35BFabi1HIsg07Wl/hGe
Sw3HwBZuQsUZzORf3TimrKItIRD/32f21/QH8IKta8kMetOpbg8SOy8FAdWDRPSr
O7UrUPPgeGFe3K5DtvB47TBatwP+PUA5a8H/UI9bOrm7y0RpnOZ8UCAaA1vTgLjT
eRFuW8/KEhvVC3QAf1BIrxAu7vCf4+GrmbbMqAe3MYCodr80KyaD9XoYPzsnuwT8
ZQ26f+pdNdk2mgWWpSLeyZUnVmPc1WlUf5P6tnP1dFNXYszJM0G0jbdw5mmT6A/Q
8tOkZ30KyQc334jP4jDwWEdBAIfgIcOqIlJa4d8Ja3uDKNf0vk4p4tCOggpvdsuB
FVLbyuRaWQGZ86P1L9w0cvOQ8f4GFV6FgyIq0xw56YHw3iiIWeW9FmwDoLlC7XWc
N67bYBX6fsF17l/1ki6mAod7MQAWqnYPPK8e6asnIu65qwaY3TN45x17aD6VN3k6
ig5KBYUjPe29S+fqZn0VHA==
`protect END_PROTECTED
