`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yqMgRkh9ION4r1nL9qdUkuj0mWAQ5y9ia0ZdLcfDbFBFpgNyU2NREPG/Duetlm3d
cRQNBn29Z0WnXCaZ27OvEMDLcQnMD2JGhauO7Wkxl1o+suX1mteSkGzTQbRoHjXg
8U2uWutv2jv1ZWqo70n7b9+1hxSfL47Tu0ws6pi3szc9KI4iz4vftCCpF200pmaO
3fAzCGGFGQur1MTIh9x2lNQGwrQoR/x3HBDrsECr0CXmyOjzUIZ70DsEdrn6i3L2
MRO6TgC/v4ZajzJsaY+HnAgY4QLwckdIy2nWVNgX3VE/uYBk3HbyK8ddMGIzgb8g
5bLJAsPAJMkZL1JvwTuMdeJv43El5UM+2GMiiPiEXka0se6fD94OWg6A8YtabrNJ
Lr/gzBgdB3jptwQmAzmSsmkrWwj9fhroeltEbF+g60uwuY+Enr/WGOK0Q9uniXiW
Qs109E08eBQL71mP3E0Ufk8IeQk2SH0wuDmuvlgL18K86uOAOKRaPuN9CaAPJupW
TiO6OAm1srEysASJYiG4yPs7DpfLrCthgPXK+HpoI/I1FA17jZFOo8xhyRUDVmcQ
Gp8kj01ouWGIMW4cvBTiseTfFbRm2xzgIggEBBdDWMk=
`protect END_PROTECTED
