`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hAH5++AmbxX8JYPsHqXovOsHNp+WTrbQGkYzHDy2E+SV3tD92LcNgP0PfhC6xs6V
D/kWcxKUKG/8MezRORAEHQIsg4hr0e/p8U9CAkDsS1uAnblVfNCU906bLB1OIxPQ
KovTYNW2auoPyrkTy4LcXvGxm9wAxijtMRxoj4i00V0Rwu6tq2GOLmSeJ5JoWSXN
qn9gZJEpaZ4ffNmDne+iM991bsLBHGckyNJFXDkzueNDIj2UnNGuDI2xFvjfn+c0
oAQ8WFUqc9Yidtqu9ZKxoEY9roI7QP/u0gKfvCIVQU49v1Y/SIIKf1/NEIXJyUzw
zuSsDWneFgcrChdw5d9Q9m9i0QXY1Mw3tz6xhNjx9+1ULd6II2T3/iGJRICDhLrR
sfkFHugtr6FtHlmgfyHwbY+Mstx/y3PKXS8MR+m5Gg0cVdWL5XTjR530gCyGFqkj
TTzcbV4BfdLBnzfAduaQI9xxntU6ExtJe1t4zNFDMciCjUMlrFC+oQaAPe3YmewL
zoP/nffS9lnDL7dP/QVlbmDZtUJy6ssdPwD5hhxUc4x0L2rP4pToxbkJ+5G+28fC
WgS7CLLaflRsVGhuI43Kg3d5dpORZjK4Mxu4/a6EG6C3njQBKH0rDb33D5c7WqEr
l06bfWGfYCfbfrrhcW/44xh4DKeZn3gN4HkevJlf0COxKpu30wD7XOICDtgnzLF1
GeesrN7VPdElJjDHi4ywqIqc+8TnJ80Bf89NjgtYEuh44SdxghS/lkCIiYhHsOvq
XKljkk8CPl6UgaVbu08a8YwXrTz2FpVMXGa0JhW0HneogdpBYsNWo7UL0vls7BCW
YLC3ZsKnYrI2pUXPtissdxytAhlhJZ9d3E2XipwiY2KJeFtb4V2BFjPOJuW5ULMG
CIVvaiqqPwJj97+Wt7/X03C1Nz9EV6NVpAbXAC3G68U8yjT6pJnBsNv4JY7EB50o
QDagIfuXWXBWWiGSz3m6YtxhuOQfwcTiG68qbyO2tc1nTeg6nV8g8s7mi6cgoZek
0KYOH+9Z9VyMJdzgBGGGPWtDrZCYxSi4QgBlcP3Ec7AfkJxj7Z3Y2sm8Fz/hFLrb
bLZ1cqcjAdMUSgf7UScEgiBUjrFX7EIAwlqRtGVEzd/WMbvU7OZhycymyGWFpAZX
UoN5XNYnOsEsUjTFKGh5h42ZcT67AGB8gF7TpGwU0J4XrVcGQ5kRn74MKlDyaS3O
E6o1H5oyYFWCUf4KNkefHPOcXnXXxX9wxX3II2xMZYDbGdD+A3bvvFu48NoBjZdv
QoBguzOWi0FML8C7crFPUy1J+v1jVeOH3F8SwOlioTbZ1VZssuzBsygCkyikj2LJ
U5WC9V6dq6CRLeHQagknhaXyfgZULe5Qq0sFRWikcc1nSb5vnVOfysy1WJ5kBuxK
fV6el2HWcQ+vkagem0QmlVslyZmg6Pusb5mL4FGkdI4RPiNBN99+0c1/25Wq2uxs
pWZn9jWXY07U/I56XrNf80nltjKtkyX/1qScMIGKxtA+twBVzpEOcAI42TR53XH6
hjmVhJhTEfuBdTZSgmiKfxUbvFnYsROvvjPLn97440NSwyZb8NJ932fSttWRTiii
aQaLgfa6kJvx9xs+Z9YTqIPHQ0sFjd53KT7HAlTzvLgFftvFJaTX5gKMQIJVrSKL
i/rQv5RLDAMtMqJBxiydOaEu9MG07X/mzBh4PEDiSJtWPicXw+GD++8WbvNLYhdz
9LrzM4WjC/963mjFpTb+sEPxvgGHaQuhosrY1L8gi3wASFXwt2aXlrTpLTDeCenZ
An39ZHqiAV8EmiOpRLkciI4QT174CLkUIVAkvcFzJKdxBWwwk369ex3020MgFc+v
H1Ip5b8SmJUTCS7/1PqoxtJ+ImmFQklED0DODCigIrl6gdCFqLGF3Z7RimzmXXMK
E8nESpLFeYULth5/rFDfZnUvmKeS/IgcFH1jHiip0x62SB+RUciqlBKfnh8UIJA2
oxC5tK/DnX5s3XDRa7YlqzKHQG7+93EGr/ZsOG/7ayEhFRnElTgHdDT6sQYG2bT9
+WQQMkM3NAV+aqqwKHItGwqQP/okFRLQa1Kuf/aPAaw=
`protect END_PROTECTED
