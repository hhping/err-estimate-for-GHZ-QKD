`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6HFRz+2vV1oTfT20pfimj3DH6muD9ay2NqQegE0B/ue9426511EDO0LxzjSmziB7
7TmKTTaiX+4RPK8jS9KjYhsxeZXGbfPMwTPmkCIttoyp4ar5OmODWd3SB3oNry3g
gGSkUEDVNdv2BLL9eArrSZ2ramQz85x2ivwJgP2Rwt2w4MaJJ13sga0rguVkjqJw
lpzaRWg3Yy4GabZ3IUkGNn7nGLWtjyEcXnlrvBc3frMHiE2X6umEcsIMEGmG8+Mq
vLL5sbh6VpZLalyuTIghWIil6iQnEq308fwQXZ0LPKSFUnp3KELorm31TZnnQlw5
b2XByUE9CCISV4UBZRYQDEYYCG5LWgr2v3hARpiJXIm2QbROJEYlDgJHQfkO4aPR
cESNrHH6cohkApbsIk7nECRy0dsrIBtq3Cv0ywGCUU0QIZO6xnZpHSf6GlYzbfiO
uJNjbdYqhALCumTyu6xb/zlm9anclTMVikaTQlF+EzY8ks/rjs6NKKmJ1KAP0sQw
rTjA3EYxgEEnmZvqYDBMemk0BheHQrNJUFVa7ml+d21bZV3XTMgId4438dMTP4X0
hZptcXwWRsAIwJpOvsdoT2taZkmhwJkcZhx8ck5uOwz5qk98yIMsK2buyZ0RY0sg
eKe46y1V0aUhIBrxndArfKOJ2Uzeg5d8Hte8mz2YaoH1a2h7IlpoUcLZ+alulOxd
CdvfG3fA0hsO7P7f/Bj7NPWskFz4KuB9eWPp5lQz/LJ0eGQhf3a2jbaS5j/oByhB
WjTPTZrO088E/z69aKKtN6retWx8k1EzFlE3xDxjIkTAVaY+RJBQCnJHOUET03fn
jPz+yx7hcyTC7Y74RuF7yzt5Zdm+e7nGLnv0KEbyXNFj/fy67n7MwqXRV2oLAfcy
GgFV/viXmi2PSwGgLZO81IvKe6K4PghDyubnBpADUxVdZmFxVgwwUIMZqc+8pXMp
ZkMHJcgf+311ckGfFAvOc6b7pDXx0VrByonNSMTp57c3GhBd5rrSU8/M7gsN/8PM
BoLS0i06Q9GhDRzB/jkgyBGFxEFf+3bs5lYSeMWO1GkzEyQttkTUAOrPjVpNJjSr
Os7s98GC2l87clOz3KM7V5Q0NOt/0n48Feplo+Na80r6kKsUDJDnulFCLQ4z565s
rKw3uou3LstA+azSQN8Yi5932X6yKozrda6OB/fPTyXsX9ZxVY5AEbSnoFoTMi+6
42j02RvqJIhpioFEMLCGkLEg9rzLroBmBq4FI1O1AwOtuahXK/cgmKYfyQumnz8e
Appxe1SNYbGtfAsjTO5js2SY5ef5ST5Pt4cBrqjEdkkGYMLFpMBzoH9epTkhcMXg
lqGyF9prBcy2sBCdH0S9Z1wZeENDe3IzJruXbrCt27x/OLBvHuFkv8j8FiNpMKl3
/UbLwIKFd48/ZUoggkQXD/S1hh/u+0pbiLaLOupwxSCTOxeTojKLN+x+y3tDASP3
`protect END_PROTECTED
