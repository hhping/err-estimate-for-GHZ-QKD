`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qBaEqJAYbg27QWwhgp4Jk1P4Yo4qh0Z94nPl4lZ/4sN6PVBu79Hkq/edjhp+myUd
K12JAHHDzG3eO81UUHPsMZQG23pRLDwPIXAbxboJ2ooqslzNhZCzK2Xjn1JM2ME2
rTlzAC+vjfJLvH84M1dTGBgnwhizHIu2gGb1hSHu2jzDPj8pZOQTRaROUpcIjSnQ
+U/cNGdz/GlWyT/3dnZd6tJgi6iGPpWCBY4hN/ZEG2kRNRzM2RAo4erZ+z0SKSWi
a8NnxMUWLlC9UhEtz5QpNyRIMYmX4QAGPb44TSIjg2SV11OYsD8C8rjUHoSSHyb9
2E5T5HcvVoM3VaqlW34N1CCwVJswWU2DjbpmKoWzJq1a/2Syz+YcbLQ8owTsYiNI
2dwPkiKRuke6/dnMF4m1T1uSPw99iGDZJ9LaFEd9zNAycBWxbLzSndcZbWV2mEON
4s6IXPR2EWql8fLRBzgfYa27AcUMkEoOUfiAjPUT0NUVVYCKOuBLC+BLi3E5WCQ3
59f1JdfZt155uJ2plop+zIv1E+dcSUorUNi7eJO1A6+ICE9Bscy62vlXrbdbB21t
tPex9x0+NUmWNF2JltMdkNS3Kh2ZZ/xw/Svlto7UDuG016uuw7JSQmnzQHdRHHsG
TDVnaIyzL2dCwdWD9KISGc2W3Dy3MIsYvi5ibrCSLdw/iB1thBveswLO1Mta2nZN
us/D2nuCClzcCfm+3fDgJASWUFwaNCGS706tsH0lyWFLHZWdqabNhFOD7rZWjuhl
y5xeSI4d/np4Z5Urx7tDXyuQVONFP8ERUWS6LgU9uPCRrsZ+UHH3bUYbYdXZ+z+H
WYziLIqI9koRFPA9UjmWWOLJkTPzzGJLajixko9r9TlZkjhuXsxzb9OX58AKI9Qg
KYzZ9OI+HChHidmO7xPvME4pFA8yEdxPF3oTUrTAkN2X9Ba+++Tz2uucKb885kOR
9TNhTTcaQNqkP78AgmxGttK6diuJJw9K7nRuYg5vyiMmsmpV8HMht3uNsocmwu4d
OUqymk3BI6+EaZJevXwAIOHBav2x5ffUVHzbb6E5qms0dNYryaDvLbes5XBuvmF8
mhTX/dCfkwvx7UI49aEW3bdd2xPFfjfLfFdeTfvZTrBzTdm5zJi9jRd7dNBv+c0o
YtIImCBADI5MxNlM1aPVQSB87kHEF0SOWSEnqsdGjvemnE+FJIV9R64euSX6Ww+K
zZxUxwUsZGYjqhic5/SWZLxHTq7n4l3OICVyiUfUM1snFs2Uw033wrqMDo/PsmbY
qO+K6pTU1vtj25T0drq+yH/8KfoVInGFlEPptRPM9ugs0qE+hrglzr3eaup+mXP/
gzY6FPEoN3AgqqCf/0iZh7eFNZXd3aNppMMAlBP7JEKD2o8NiFAUh8sfaIY8VWjm
u1buv91D/8YkI1LnQTN9LdmorURP6vgQGr+LgloJ5+KY2niulhn/H7FvbKAhPc+0
uMtG7kPsrdUUTbDA+UK9qPxo85dNE08kgKQQnfwOj59PMQoZT/JxNvIW4sH2j17t
8Do6dw5kBKqJJUqlwlCAaa8zcb5OjvG7HpQNS7GLArsJCCQvlCe4XBb8Bwfj3NXr
Os65pWTR4QabfxygY89CZuJKZzBGD2v5hfRlTJvPGXvtkz4asI+FQmmrsdpRchUe
3Y7o6eBajIsDGuo5D32abxNkl9ZlyrLnUuj/e7DRa4itLEXjKfXLEDYBMOTyJhjs
kvfbMYTPKyIH8/NzbNU/Lz6kCLpEZB17e9ZbfH5BJPrE1dFB03MtTka/g2pK03qK
SynnaP45mFk31ygp1QoPxvvakMxhv+YVWNvpzamG2FC/iNzmSnx4ZDTlJK6cxk/b
YBJLoWeL44E0MCnqbIsKQXNnPMl3SLB1vrfzUTQhIP1B2lIPsHibmzmb+DyOP8Zo
z0r7pQhWxQZJbZufjdl9jdsJG9xOadmwAFixDHM3FwLcTcUdg8HrEtE+Adkt72AQ
ToTKM7uRwLDNtNuWz8e1mxyyp0Ogk8EIw0m236JSOtiRK87f0P8OvQKU6ElO2WFP
W00vT0OCzddgpHe7LBQj75IoyKqQzWlLfYOgIZWfwK06+Ct5XOqj99Lzfac0c/oZ
B8WFH2/Ak9f68B3tT1JZO7rYkTweP1zAaffDaTdoj1wVIAvV3+qhz+fqobHPJI1u
xen7+u14Me9Gx6KEdcaB5Rd/LpX3y6oLi6x6OtkhT8i2I2CpDMh03HDVwn29kPUV
CyavuiQKE1c0FA6AMEZ3OCKsInpMhonKTC59NZkeBm0JEJpcFb0zg/pue1IkCty3
JBW0B12nycxD0Yn2biFYj/qYov6OG6At8KYSA8HPo4UJQ0yKe3b/ip7WhYP+c8FG
tCGaeC8YyGH/JKM/oqYY7VJvEwFPHAU0eCiN820AM1HzngNFWU00xTk4aKEUhIBX
bV/FxB5UD3FRrb1PCWbgrGUvafiQVzw1TCFjLHEh7EPM/TmU0RR2E6AZCpVITiCc
RbUjT8vxaliEjJUcT3Ayjrjdj0ne8WzggvW27HoxyFE3R61cQS5+Knx6f9CHAxOJ
lI4a2pV3cHGI16ix2BZmTY0QlX9NFxXsN0y41sB7QpGrMih3OXe4y9+JjcZB4/SN
LSOoegZBWQT1G5hWlHm+ljeTXsyDJ4T0c8EePwOex6XCeOfK60mqDZGmqICRERZz
2nIXJI5MxqJGqtHPDK4MBJrihb01rpCm9crZCjCt4FDVzXOoQZp9+ED7BXIywYyQ
dej4sI7G7g+6ykrJM9MUsMUGKCid82x6v5JpIvjEhV4G1HBTpe2lYkE/m6y3u8Nt
Sf1kwFZ7qu9HhrpnDPTHteoCvPp2F2/ZSu7LRmPO8+ssX368ALyeSNkZM4gZOCX4
4NnqStT78dc4r7NcfugUHqqzvivZjQIt+Paet6kUSz6leTaHSyWkMWqz7WCss480
NsXBwrgk2jOGAvSqkO+wc4Gh5gT31YkaOJg6ckihEQaRLhuKkbgP865S0ReFoNzk
J6Rs650e6sEaxRUjTyUtABRIB0rCjL1nLt0p/phOy9sgW5DlyLGkB0ddEsFlOZv1
kGAg1WBjE8PYFigIXGHFcj3YbRhDujyN3oOdT2kEY8/+INhaKSNQPDK/zy50pcaw
p1bd1KAR1kaZEougL532K1OB34JzWlNwy0i9Zr6+vR1yQjChjJPAewobkiZrnk52
rw17xw5yGsVWku1jW6mF1Uih9lBOsvMKBP6Dpr8iqO81CSCgQKk989Fvvgr4PEXh
1gN9BVchKTQeKaFw5ihId5YPeOsq1udJF0MghqJN3RMnAfciEOrHz9mF2yiLsRWD
NM2Ql4uB9UQDjJAQtNbcibBCAV/tzUGewSgKrh2yQyRcVMzPCFvcPxn1Kkp0dH1d
pQ14tyO4G2KZGfVsgOCYVvX+W//uEhNOn/ZDPL3D9MKB2NNvQ60SYhyy8VQN8ksO
pM8RrJga0tQ6T8PRgCMQnpethekPPrOsgCH7rP+SCMJjOwe4zlQZwUGF9pMbJb/p
WR88IGAkM1fxhcINZOkhevLvMaiGr7G8DnwiVKbeM4mCU9rmq1BGBiNE5CvhldHB
0+931lHsWt4A0lPhlxF1nVrnRY2J62OuoUdXiphA+qEirQYPr+YAUHKwOIBjapyc
uZ60J9+csQauOKzzYDdKO5K2QRbNDvIJsXb8zU6gbQ2RaEq7r3TD5vEt4fdTJixA
4RpLJ8wxzAUrKDMl4ZlbiOvWpI7JasY6hByLN48Pz/3bxWFzr6OqwYE5wRIcL9ON
AmgtNYgbs20x57AMjcWBBF1v3jPA3L90AtAbbQOh+QATTBb+1yQdc+jQoGTdYrrf
gLZZPXn/2X3C2d/u0C54iO9scCNV42QvVr7HekInOol150wKlGHnFwnCk9JFyUHU
vYqkIPzeLJE7ZeaFlrbIcZm4PAuv6skfYsTQzgCJ54SC1WlJwTw55NNCJa0PE+O9
CjMTfLoOG49P03J+JojJ814cVYWlMeEXCBa80K1MdQOjAn73PayEkkk4NNYT6Wuo
h7ReiklSZPc0wS+xlHlTxRC8YwWZSL5fRP+VNON8X9ZzH8oQFGw92yUlHy2DhB+3
1oc0R/kdoF3LM0u/cyA/StzOeK15YtI1vWZYAUBoIVn2XxdYW4zGnfoJ1fA9OVBu
b8a1wz1NjKNxlsNKvHLXcE7aG6nSDRcC8lNdGqsB6+m2sfLyF0kGs3e0ThxhD93c
p8/TATa8955CMlwXZZHHL15w7urG6m/TPSLOxFUN+IJEbn+s5MyvlCU9ASbDF4kk
e1xwrC4jjCXoJOz+VqOtZ7tWQnaR7u5YBy9Oy/BKSuDmFpZNg3RJFD+/fGdzuRyT
/BlFu0W895AdvtqllDhd6pACIJaS98L4jWH9uoOlI6VZpe5uKHiuy5VbSOC1M4Sv
xjzgpqzw7BoQNib9X1BRrwYJwNy3kBu44CV8Sko576YtRBO3V+NdmEzBY1q5oOOe
U/df793zODd6W/17v9g+sqWt2aC2tfFykWHkdPd+OBiXeNeJMx/+GqyH7491eMM7
1qm3tXWCgnUVJJoPn5knMTumve22Dsxeu3jFKlvy+AjaHGmAw+soGUlX07AROK4I
dUZTj3NTMSXAtAc/5HEi2VV7HpWrraTELEN7LdBP0ns=
`protect END_PROTECTED
