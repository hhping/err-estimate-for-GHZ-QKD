`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j2D8Big9vmVMIldpj5fGly1llth3rKHtfpgr1YAEQiJu/4Kooh9BcIgB8nBEJ4sT
v/0pCCYFWrrWgaxCfMG5QPemH/fPxtXCL3YmHW29GmSx9AUQZoAjVCgYNyt0N+mN
V/0+Ke5y+8KVKmMsxyzYorAXvckrzmL2Mit8XYodmKmvXxinQXJtZt7185PM0Nv8
Avbx9kX4CNJhw6Msr7P/8lxZxttxrjCtnieGwr15Y/w7453lHM/TJ/eIwtti6aDW
7bAMaSu/6n0LciBBWD6d0oR+D2LxgaU0BILD/zW6pgc8u1u6VQflfGHgymx5rZHZ
JX3rzKFkgBIGdhjBE1l8pIWIsXiK+BMfAzedwZCQy9FyYYpNiVb+I9woT+uCg1Cu
THn561LHA3rkBDgrMq/+2RxorWamQQKVzC05gT2ORdi/37b+hK9rVCPTsTg1PXsY
9z1s8YMLdF1oKZ0i6cSYE/sYrz8UzKdkEa+fBxCa9tXcLxwbUdfiG7kMm/60+gQl
fTeTryFZ5+vTWoKqe9Yi/zw3YP24669O6Lx7v5HZ6a+q+zlhWNjxJmu2wMsytrAk
I+rb5xtJ4I4/5I+sVyocUGUQ3Nr1kD9VkAGEA7Uu38YXi/PlGSIqNn5xMC+noY6W
0b8O9HQEX4ZujeDY1qaCnjgLRTiiRf7bB91BKnmmnazhDoPkGrtkx9BDgUOVzxWg
lJo1kmNqIerRFFrpHeTqQ4ECjRkk0xZrSj1NWvZI3HRsXEbbZPqCOVPsHAlgn5r1
cCzOYvMim+BXdfA7hUr08jq+SNSh2NT2z9tkYRScVXGM9NRBMD2xOe3W+CbKu46d
KPAU2xNp/H98BMvd6VfQI7NRe1zVSH1kN7K+OnCklyYDC4wSeazvRMboiJEqENE7
JGsgXhD+BRnHhsEhE/kQ/4XMQ0J5mKvUBd3tEUi4VL09Zg2x8SIAxxz5uPAV5I3z
By+gyYiQVuajaBYJklVwboYVsZOrJwbq9NWuE226j1/+7xgi4tgDPu7kMkVyK5kF
rPW4AniLiDvsGh4ARPzm6sofBRFMqyYu+h9RP8N751HuUS3JPHoSIiD482YLXSEj
ejTQxG2exZCfdFRfOXq2MghcJQEzS3vgjGp6ObqMnMMmvX/MakVx7+WJeqKk/nME
bzZMKJPl6tkQ2tT7wrRevrx9BR9+qrueCyLIL6JPNu8AoldlLbWEzIUdpkHVvLvA
QXPfZsHFTKx1Tuis1kP279leWDFGAzgOnOL8b0irX+igS4MBiPyOVoHn69BKCR5A
tQPpKMUQfX22Fv14zpvWQi6WDafBc+ab08YxLPk6zZGOdUYOyu/UuqCN4qZhM9M4
ynrSX0u/v9z1FoT0Uc4vlaQ5v1Z9u9xfcctKD2zE1FvoYACJQPQeFyOJvef2esSi
CZSntviFMxhWbBD/1K+AdYIgkWuQJYypUqNPGpQMgBGWaUBXB74xWIOGmD+Vjxrc
ngKBGxleL2VrHRNjg4Jwqcv8FCibsCiJXF1AYeJAC29pxWuFNSAKgk0RLvS8Ac/b
RDv64sFOFt25qnnRdJIRRvrrK12YF4+Gp1G71yFv09Tz0SLA+UEoGp7Re/cjerb0
/RDI1SsjP1BQcWqbglAtg0mq8fkZKvzY8YtvkMk64N1rBbFQ21zDYD3roqvdSdCT
G82tntXfFh7x9NC1eDiGFFuuQMZc8HCK162/DhuV8ol8Dui3j/gJ4Gh3t2W/N7Ul
gD2kJIgYEzaZoQriXkh4FKr1kLa+l3bOAQxwoqlBGJCbCVtSTyY/OLOwft5lKwYI
8IX5lff9mLVP75XhDfEPe9lTcRHBHBGErq0CfGmL4MvCgkP734YAjByVyPjXqd+9
xVove0i9WHI2id8ieIqWyfKbxGqphyBTo5fEXVdcD2podsRAcQmvWtrTFw3VRoVM
QXs09iEK+72bWNd+PfrKiXooqWjCSoH++hx+GM1S1RJj63RRH9/UZnT0OgNWKwNz
DEudPsWKrr8lkQHXBOCVENGqblDRVY9E0R/lJzi9PwOWcK25LXWCiJJMGsT9LTjs
8dtXYuACFZL+pI6inwTMpI8cCfnLdWptNx0PEBkCZQFcpdQDfAGQQSMzLoFm9xvX
eV1PLFCT1Ph4QGR7EBFQc/SOuFPwdzcQYqh6DpCE+44NezlQC9I/XlsorrotGw1l
5Z9y40KhPNXnAfcyAnTe34feUq4FjLXf8BwKev1sX4uS5aSbxJJCcNKkke1YN7Ny
zrzSCnq8MYpVgMPY3LV8DgaBliOr+y4BzriXG0VirMMTb6G6j39ByWz9khKL189O
zBB+gpFRveyWoBtQicJAuvjCpLCv4cXyfkzIlGwwOG6/NQ5kI4KlnnIS+PZHsHjM
tpRZd/fCQe2DMgmJ2AY5oNX7Xyf/+Mw0ejFM8pEWTEue/TlNzgNllWB/cfuJJvb3
eSI5tsjMm9YyYRQcf3YKAMzYcXpRsqdAkqKqXnywZE26VC9351qqmVh5ylUdDEZ1
cXFMKpmCdNPNAXz6HWWVjpCP/vMPyJSU6wGfGkGnBO/jbVTQTglXIQajP1/mO8LL
7oOC92TWzVKLhpqACDGlJMaKCtvukTGGaKYrUbPS+zcIU06LnGqg+LmdS0w00/Tz
scAAJQ0u1dq1aY20LCQh7iD98vw5Lsk+sWwaZOkjN+dcLQX4tSaRHyx0j+Ey8DlE
vmG5q33cNAZz/DOu6glpY1pGkU/xtG13gLDNMNxl70HrsUevzXsA5wTBecfPrqLo
d7YLmpVvjVDklCiKQeIt6mQaMei2lJGt/ZDpdkqWmkvdOFEJtVcM4JnQgYyredP3
pm6YL7CBDUZk8hbHuMLtRo3wzxLLK1TOnDIN8hNpB6UShzwd7pV8thVkHjzwtMrI
uwXccUgPynQVcDkfvIP+PFHjSroov2qmBlxtYMdiNsjfYGV8q3NZX5OBYEcNKbli
s+bEH2rjHP4GDcSq/gQnTm2cBF7vhtqnB4mbEOCA8KOMknZ5QAvRs/x3BmCWS7gW
h3l+3ddfnDsYFlz6daaJsuwW9V60qFnz8VGijT1TLyW1G4uJuvYoCzpBdcCNTWzs
/FKls6QvVXEpBnDqKJVQaRVs8YljgyShq+l5kK4sInD95Xm+6dkgyV+XL1E+fp36
DdnkfAeer/+NO2YjXKwyP357xIl09y5cx1q6LYkp4gwZ1pujhR6i9aCGmWhhs1oe
6xc9epnQJNmcicEVqk4azy9WsAc7Ae/GdLJQj5TMKp50bvP1Y9XMCY2tBRHNZk12
WTxkineOvpH9nskf5QQPEl/UBwut/CpnElJGm31RJc+zt+poRhklDcQKbLWNYO1l
CpIIn+qq4RCOfIU1J5XUeyIQ/gGIUaKE9sMyp6aWkTsXQE1Ok/Bj3cYrNsef1Msq
dQYm2ZW6smchONVCIe3f8/VKF6UHoMgocpwzEYQkhXxfGkB+y/q81DnxBrZfBzO5
+sSKWjxrqigKU577M3y+ktVz2aKYD2NUrPdagzcdTzyQS9mZCihQm+XHZhhyAenn
6W4B3ObgbbyyPuDetyHmPbfenaWhKizcCDxmSZHCwSh71/ymEPj6yLMyAki5Y5vR
iXwqc77QMc543Uo34rFYs639BqbteZRDVLpvIxpu8T6Fm0ppkN/tTeYqMumpYlUA
U2qU9Bz9t2OLloViQANcB3RGxcQPsx+raGQo3sZI8hU7NjxqbM89heXlxheX94RV
ZGufX5D3FXAAQSjv7cP5G8ucs+IkSV/H51Kw7j1mXXz8x3tWsHsA/JghXFr2sE+E
z34Nr0/F8P0wMCvHgixJ8n3hcpbJyXtn0T0urDJBlDnkSaX3Ur94S9U/FP84soHR
112zPGJ7nYGHw7rkpiEnKXV8pj4V6BeF09PKnpnUr7igAqoKf1O3soBa3ejaBm5s
WmasF+Mjj78AMdDE/fscULQL0Tcgr27JOS8Car/ZRprjamk3VIhojgg9vls2BHsE
11xQSXJg8pSvwOH0Eg1rN+tm3pi7RZLThQqqZF/gla6nLECnh28Oh1jaVuhb1vXs
rxaGGQRZtOTEP/1UNsnt9ubndA4B3viaj73nUd56y20eLCX0LNKo+oaivmUbh8sY
YjZdOCBsSk7GGrfoj3F5xvFCynfPGBPzMWiWRoP5ZXGez4o1qWr5uFskQFU676wY
a+9wQo+mdr9U51YZRpByY4lHCnZ1PL7QhvjfyjWnnr23EhKB1/LkbDg9Wcpt6dl0
3U7VfCOa60qU5Iu4EcYr2R6L19CtXKzvN5yU8gSWYtTGJJLp/Q3jIkX0VaMRgSWD
LvzHOpAXKE3X9arpMtMDe/DaJHofkcrcS9fiuUNyEEB3IROC1vigxB54px6ud0HA
/MLg+oPGvHPeJAYeyJ6wKrR7sPwCaIHf4rUqYRQJXl0Uz8r2Dxrw/8LaM0Lrm9cA
ixlBUIpxWtVlP6y9sCxplj/DGxHCrDLiHgjSDxv7RTUyMg42JRd1vxgEySOAdwWp
QveSRar0NPkQTMw9KbCGoeyl5pqh2GcoiOu/463Z9tfPRNCkSJht2f3VxbIWMeej
dA3YT7Gjfz6Ayyn2XzFWdPlXbQ0/TkJQ8C/YzPc/KtKKDjniIOx4DaMvkvEW9Jh+
erkR25fI70NJhPXUH64ACElVNmFnxIhIhjd+cMrT0k0kLbN8kt8qA4qApLMK9jyG
RwxL7OfCVmbBAPug1pbe9iShgceHXcmHyS+pq62GpTCdKZXHvEJDUkGUcj4wEnJo
PWnbo+xwcPKyNuNr2sdF4bKXynfnMxPJrCG75sUsUw/xpxLd/tFgJTHmGOY0iV2B
/d+eTg8aGbDQJi1nGt5aWc57e1fOseclj+OQ9TTT+3HkPL/kEI0HmqRuIRNEG9N2
NA7QwgDDVlpyY+MVOptB1yFRW+qF7Z+MbJY44WftYov0cNw2jyfbXw+w1JPOm37u
N2VXxqt4dkn/56OOjs28oKJLTCltrQqRMLDTV4pwTrv0K13YfOprmQrOttJiqU75
mOCwJg/v9B7+Jj3I6gAZ89G7feEQh9Kq0KfN3/YDR/OhV3W5A4drLJgmKI578EEV
mO9Y0E3RxQ8WRvNwCV13KnNTmKuO49nFK3+t9GgNsog9ocapo6b8suGpL9Eu1uMl
mvCZteXWdko5kZcqzHDKXqLn65w/GfGcomTLzarCRqUjEU1kOXOjodicPpsiQIVN
7r3l4FBLoNDLxHSDSjIVCpUiW/SaSq69CL45/7oSHVMnifc2hr8jMG4991+n/gwr
BSeMhKTrwEKr/V/1XOZyUlYl7v4OyaE8jEpGUvqyyZ19LCV6lcfRp5B3BF74SxjJ
w1JzUz65/iuZJkeIJ+LKwmTMUwbMVwJHEyVkXyZOo2iUY/QL4Gm1HdQe3CMT29M8
pz6yAtkqgIQ94bh1tEpHyYNARsDiFS0QtG7FeFKNE0vtrxTPUs4ItRGi/LYzni1p
Yz5z53eV5IykcE5Q0E6IYija2Y125QFq6FmKSO15I/xY18sikGPQ/SYOaYI+hkiy
0zJbG1ICgUAtWxR1J3+AyTzimAKXh/C6Rk3PfVOtw5eWspBXVDu8LPIzOnFNJAzr
E8msfpfpX8pq813AhXjcZ8vk5uVd/GpwrGVMfoT1YiBan/N+9tCjquttVdHzT5hw
hUsOPZVVMiak91XUYbvHEPy3tfFotNXwkApXBmSnSXX+sL4e68kexkEnLVcZO0zl
29TBdfk+FtVY016jOmc5XtTDn1NJiGVEk4NA0YDllDtU2XlU8Kui5HdoTjzWCJgg
iy1ZXYBmm3NnvnQzWzC/z0ybxcyN5Kpld2OMlxj3xJThmBXqGIxVg2B88mPzZOz9
EhLOf2EkGdMVFoCGRu7dgBr6zip9HhFWNTjlC9GN3qybJvCPWMDborELykXkp5EX
1t8JvdqJribHqsQqPPx5DXQiM+/4PmIGccjggwqE8Vj7gNjQ8nXV3WxfE9pnghtB
Uzxppp/NNVCD7FHkPsQx/AFMoi68chQCFCaP5ox/MELuH2Y1TE5dv4IIqcCCMIBw
MldufLdBTkSMs2v6Mtn4OUzQ91VhBg0WXsFe8yrYhDhWSu1ZOJRDnEn7RVpds4FG
dL4P1pBBrUfiNoGgT2RY2DUXpWxnle9Hs0Wjr7bqNLmEZb7tVZ+G0As/zHCXqpk2
Z+3PBm6gKPBdZSO9Y1BnEXux1tUAqDQ3azueXoizDNf3Ci3Gp5WUDP4T9+AtL9tc
955olS0bJqHkpxn38WxdfZYNrxQtENi9FEWv8P8tKDtdIxRwbi8O2spZqhYPGrc4
nAXP+mYboDbUFmScB6D2hG3pvApbzAcPhhBpgC61EAjHhpdBi0zOJsVkcagC+vYP
ocjtzgcZPkB3qVwZdb6GjkGmtHt8MpZ8k/hwNb4fF+tSz9lFZG8M+/PYEzBTNpdv
/ZZnVvXLbuCUw945qVPkVFfF+MJseeC+lROuJCpkTA9oGy/9pR2jTUjHsQ5uIKUc
4KhQBfPrf8va37g2xcZFmU3r8L2DrR5vpkK4UDBr3SQoGaVGVWoGVGcx/YwZrvjG
7AyiulTikZTR1ddwhGdBcPE0w3ML/TYy/HxgxggZVyq7GPTxM7hqSv7i4sINF+QS
bAcmFOXU2KyjPo8w4cfmgNMFa5PWy0NFSK2iIjroRy/3SQmRuiIlAf9vKLVxlQer
3oTLHZcQTbVngMH/39Gg30GKpXmeYlERfefG7J5fwWhKY+IOcqMpCiatGQu+K7kP
YdJXDfM60NSeVq303qnum+WkhpD1aYwJfQoBtl9p65zvKTlyUDi68zbxiwrLGZjd
JSYvwkFuvI7dmqb16svGigxlW0XYVPIi0CuFcq9tjemmit1gQzy5j9plZjDZ2tWY
tD4x+QSl10xhFRGMifA+1aewLzG45mO71eS+ecb3j6DgEH8MJ7y5TsYznE3ppF3M
3a84aHhWEwsqd0zlfdnH/Nia08eUGdSKZUkfPsstY9fGZf7poePPVBXdFIqKsYGy
eqk1Gs2Wbakpomb8qy187OwzTMPsSmHWSIDCgZCdjQAG0rjxgtXusYfGmOZFoLJ0
7H8v3FTAQtYyAdGNcnh/tBs2fcjEWXiEJlCMJ/guKkG167nKN+u8p1TzvnME5Q81
q7mRV/RqSuhIb9QZQWwX+J+euPOu9whtebr8bv8gqNpb1XZQaIt+u9cgxIT0BG2P
/fGeH1l8vCHoYIsx2fAzU0KuecYXNInIPAZvcHt6qg322JUvijks86Mm0vtLfKF+
W+88lB8f944siH+plyWmoYvp16WfyAc3GoYLya53hSRFsWJ446x2Q25r3n7mPcIS
MdGXZOYKDbDyZQnsZeygigw8Alty52nRqCW6s2tl3zcME2MnUXSE0r/t+Uz7nun4
DPZS3+j2h+N7K/kQsPFSDNuWcWFhIPQqZVmhseSMTABdT31Jg3SXaLQAuIIWC3j8
olYfOcl3Ko+nn/AvQqofDFGU47y12HFMyTV80+Rx/4QcwrVHgXNs8PWjw4UeLffL
uqx4oWhhi+DyTJ0VSqaPaCWmnoo1v73CJv8zeMLtUGRtUflejgdRLPcv6Lz+2c+9
9o0ouVbGvFntGFvq5gzaGC6NPhZRDcZwj1YJ8eWlqDKWsBM7ADLL1xwNws9AX/W0
YqTPt4W5texMcd1Ym2G4LO6ktEhp71NwGUra5mOH4DAo5LMS0T90tvxw0YNrzkvK
yzcrpmXpxCOzWgSHbbz5aOWHhroo7evYdKDOY7fGMp1I5zTMD/ai17GP8gESrlzG
pnOBn+8JiB4ZgcScOMQGmCBL5xumyWwiy49SVBBOfP5Kij+Yj7vo2akBEhy8YmEb
uitMW4jJfasRS3GvuiZJYt9z+MW+cWbf4MHfGURPh7tw3uLOOej2C1umByuODpfw
fLYLk8uYLXzymYdBzHrdaKeGmB5EO8beF7n+Keow7AosAbDWjNixPQrV5vhb8fld
Vka4AVXgxqKeZVdieGslX66N0ZjOSFTbe8zdderD72F6p/k0YWPHnFSMI0cC+NnN
cj/mM1cjxPQHa8JxDnSBQQ9rZ1b4RgDPCSt+EuHvYp5TxcpAkTYRnZU9Dmm0qxro
dRP4JDFAHbIXESWdsnBer/rWRlCD84QT6br6BotmcXDp7tCBCCkxp7/U6lhQIJoO
m5BPF7fRM8v3+vF2bsXQ6o1rPB1r9zX97hl48eh/RI42i4jGUT0NFAEZjW1D227N
Ap0JwHgHLdX+qzKE85Ccp2iox2RzqZ3va10Mgs1VCs5NtNtzx38yOHijqQinm2rA
NI/ZFB0CKoWArMMha1LmvjiOKweTqSAbDQ5kCReQUDw59fGeHQR24MCkKTkXlrPU
zUf3OY2+7x0MrF97SOy4CAjknY+4IErqTK+AQ2fRpHx3xBiyVqGvrGrjVVdqaxsa
NFLl9mBp5Sg9BAX8r1m7/5X3G9B6ut44BE/xAppnEO5VTdjwcWgSi5/PV2IN0u95
juE7V31jPOMpf+8Du5POUosIP9l3C2gg3zPBUQFqQDvYTMrhv+lOtOv4SpxXiniL
PReD8EetnE+vs6msz82oxXuvMcZOTaA7e35ANWY+Wz8VzyJZ/lscalLe87MvKnT+
yYOu1eYdaPr9laf+0cQB2dF4BOSRsQ/8cCLAP8DjKQ6FhjGEOwJqTndEpqr/F0mF
KBziLuWUNY5sys0PZZItn2CDGy+ZTMkgKLagEL0fiynqVZcsyx/eZpVeoEXB5w3V
FvoAZzUPSQ4nj7EI39//OcQtFIjEtfRTLmo08Yz8Wb+3AlFA5dOUpShle2D//7kV
5vAgJULV0q+toemwQmu+DyL7rk3O4C+MbpQSxG67CYWvJIDIODH8kRt8I9IG9eVU
/N90KzshEy6t/g0zuivfCMVZePRiVurHvjM4Uwqhf7qsz1enntmxMsI19SAspvzx
HM5Gvd9IZVX1yiyn+bTsrCxcriMqYgpjwr487zAQcs8DdvgDGbbMuMqTnJflInrN
uSCNNTqubSDWxd0cdDg74/ut39VTyn6y7gLYmwavjTx0wTaiAPTa0g4f9vy2UWvv
l73PbSv/c5QQDpbPRlaHturprQAmeELHK6PfzTPEmWLhO6EyOO9Jq321zcDrZKyV
Chvx5y/zCMCouaAvYO7R9aCjk2BhIXqm3hc5z1QTlwaqa+1ZMDuV/Ydt0cupycBA
BBQUsG0G86z2CJBjEsq8VH7JVyGzj0M0qpIuV38itbW3kJYQAcchuDsV7cHFvjFp
wcUPf02Sb6CCzCKfYj5rFIb7nZkmDAVHMieyJljDxL+hF37QteE8jbrCUqtV4i+V
AofTEr86DwjNzvAxcK7K1C0y+WCFMzu8EEPrBsGZy0KypSOCBEHokBpCTeDQ1L8C
n8Vu5bCBEKT9pSFWTw1bBW0lrJzCWRjEuw0dtOtSkocTo2CoVHmhgSUuN254BCgQ
hDdQStIOnXURTTKK+i5JBnTbNdaInQVT8AlB4ec3A/1iQrP3m+cx/xTYokHKuX+f
ueq/JjU1Bjdyt/02Q50sGP0sTVSUk5X13IEbElqVCvZEUXSRFO49MrJLhNvpMoV8
sgJpbKQe05QCbBQvcAfDQFNxmctsiKFaNmEOVfO/3WLKKLjvsrw4E0iiAjSX0CN9
rO8Y/M2ZMO9X8/nO3OF1ayzdK3e/pNewm0QFwT91bErGBG2T1XvzPWoueA6n0Mxb
yrbOWdgqTE7DQQ8XkvauqxDI3h9uOsCpQj0Awcf+RqDRrtMUo10SmmecpkUTWmiv
iwKRjdHT2Lw/IX1stZwG4Rd4Sb3S4epnhr53TsFxL5CCrEcUkRf9DykAPk4bmEzR
uWF1Qa/NcJ7kj2CmdQCjYf8QLjlKs+K+p9G8e4rMHTNITSq9Cu9Fe2OnEXuLkn//
kBWeVMvBRv/IYSjXHCpNFHx9ymv1iBTAde46HQ5i9QeSpC9aaR7JFq1HWepGubfj
2wHCFsNjEt3bU1s6vFKC5sV/q4WMH//lwMBTh5CxK7UAArVoF5VyiFTBrRNnOkqt
kdZ0AVk7d/nHZXXJnKrLENOGssaaFsra6zQafn9Cn5Vvrg7A6dDTdf9KCcihVzdd
x4lFcOr1QU39jD16WbYVUPf/psTDrEAVm+uIeSQF3fz60idAc5Wv2m8nAJTA98VY
ziu6Hxj/igeqaow6BqfcV10Ag110zj1UK2GnlCzJ5kOYLOCbYDxiLUrRTlQfsNJ4
2cXV28vF5GyboqZV5VXkSviDOY/ezjLbxL9341toEeG8hG7yuER3PpUsz+wj3ybP
nUxlckaCo9RbsNdr9Crz0Sdfn6d5AzJUOuDDd0m8VRDIcGiRiIGWZ8XJj8sAvS1X
jMpfQ0IWCW77U+nb2MnxUG2piU/i9nJG/V+cVwj+nqLcpsSANdzi3/s0apijN2VM
TdXcvALFGan/PezO1JDHp4w/nz4B6K1WicqGHknKEZjLJzGiQSchZzo1KCXeQGLN
bLsQzeRqqdyxzPkP7gu+lgseCCYrmwg19QsyWFXsh0w09sMmlYxV0AcyFgaAIX1V
Ab8r6xHo7yZWC+YY84HSHpPQHAEMEftevybdZM0upGpyrYn9S/B5Fnzg9VpbeZ79
hzEi0memmC2Tj1oUCbAbHolnCzZiw7pJtTuRRKw2MOJdvGe2lria/A5jh6ZGJbYU
tTEMFwqOXI3E15rUxkegOq6PhSLMONTIdM3EvFTzF4Yiid76usTtc53h1s18tDBK
9KpQ2PuS91fioGM08M8lTXzoedlBm/Ak6qm6u8uv0WVzaAelFNeTVu71V/stu+6q
HpqOzk+KLu17rXrZotAXWmGU8xyDYnRKS5ryEEa9MEQnr31pnDHaUSSFKPUpwo2v
2uZOK33PU8kyIJsWHCaLGgYCCNoZvswD1mcRLWoBi+R8o+YjD1HezbdFdZBbgCLX
qMMg012b1Hn91hpL92fyZmpDL3QKHdz4sh6ZWfQ6W+Wd2DTjG6naRMpfeKW+OZfP
sfdX304E1zOVolTZdUodAeCHo+jG/f54fKrCGqJwiByHbWaxmtE5juksVZY/fbcN
Xhk/uzvB4pmgIs+k215LUpPDLchu5quj3oxlFvF58ZGgpKdPGD8/6EXLwsvS28qQ
qBrSUyCZZO6v/qsZSbWHQyUjkQQepcnV+cHTuMDtpWYfyKJ8PydCbQzn3Xy4aFdd
mvVdcwx1QtVDPEEk/idsnYEJjAcoYSj3x8o44ptCkAlIeIPp3vZ+PTgag80bK3ar
fcZN61QDFvPgNDEMBCoWBzwf2ZVXZvWRPj4xZo/l3WGtAtH6pxpgUJ/iCs2zxo5a
fkiYj3M52ePuHkoX7onU1cXQCtm7y5cyGeB93lLAi6Ll6raJV+1yCaJBfjpFDaVG
vtmjT5TEx7KI7JtGTHyabwAeu73Hhz2UHlzYMvP74m/s9S9zplorXk8knMjgt0c5
rhYaitw4byqfILGOLYafNBiv1BRR5RIYZplCTDXyB9xcvlIiMS55G+KQC54T9IDl
8zEhY1PcW04Kkd+HxPVvAfITBNcd7eFKcALVacW8o6rH7K8o9o7tNxi/2w+0o9Yo
oVxV5LuHRlZRWb+VQwzW3MV0ljDO3rTBndNDfAM5KISVhsF2EcYZd0nUE60i0ieZ
IUaOFhjw3e8y3KSMyp3FWeEW3Av6Mwx21LsZXty/ymwqUCLsBwiN0EaPn8jeJPJa
XvAWr6vY80eDSyMHBDs4a1jH6sFj4WGSCAzUGDUcPakLg5z2rEmXZFKptMfGC5pa
tQFtzmzUiuIgI30c6Fs8urj2U/vIVLi2TZE9TktcSziDzeUtduJQYZ1RuTGX3FE+
04w4TZ3tvC3sPUh95oTKOEK9/xMMHky+puIsytWysgz5SwNuALHbeFspgqA+F1/T
zwrtpQUE42uQTRhaJJe7xq6H5QT6DlDnuQNiUIQjEO6r3R52rhFi1PPph9poK3Ke
wVE/iIUpRzymwlBPvMhK7oXzOVZHROFE+tnUyhZP4AUqPtLjGK1eN0bWCvYW4W9Z
5MXcx6a0qiLY2kvBO1VZDAM1L5FDsl8eKqg09yXbAzLrP0kPJEmfzqFnU/G/M/l2
5JJkSY6CvAqi3w2Y0xr+dTOCEWNx6VjvXx5vCo/qfsRGFG7Oi5vjzkBeWJaJXPVr
22nSKI2+5EMk6Qikg26jTnXZNQfoaYoV1SdXzrzAhMgunBnOvPoQ+JVl0bQ48hAY
UJiJms1JODHpt9+b5oQeAER5bV0s037+usdEdON7tN03bKSdQoG8KbmhbHoRbZOJ
1/syqnAarsk5lgpnnA7FUgRwpmDS3UYV/EEgiHOc+UPhL4jysPTWpwvB6lyWONZq
QF+UQIITaUXQ0mY7kHMVm4ga+XOK5wFD4j47yEWum+FVtvuA7fDvm/R4vOFQ1D0g
w7DtRsSakOp6LzM7KIXrI9KEG3iq4dbcEcHtEmLssFIkp+KPHJwHYP0V8qrprsR+
7J0mIR5eI4cQaTIsFkzOLNsygtaNcYNgU/gO21K8hNX/N39VSrvycNqcuoRBQnjK
ukyInoPf16sL1Ky1ylFMS3C74KnRqTtk1VIf7LSYgP5VwAIAy0xh0LK2tErvuCXN
u65FNAt8YduesZGdxFe+u3K1QSzhZvfuT9KY7Lp2777bD8Aty75vbvATCJpsYmMk
TrlhRVuHRBcTDa8Mdp228kjQXoTWGWC++hzqoZJcK55jWspyMxDfDW594pV3e8ID
c4o5Qj6ldE1lCzX1Wsv3vOsSeRoLUzFEil92BFYvvTWuAJMXWl090R5j1LPjuuAN
PK6toHxB84NPNv2giB8Xt/zO1de9A0sZX57mZuQPjDqaMfN8AINteKGr2fLNHiG7
Z4NLyiABv0LY9y/ZJN1+X3YKyzS3vrcFScLkrW5saapFD8Rv+G7FOZoAMuhvsV0p
pn5SRJdnvtoPuX6a1O4I/Y/+GPC6bInrba/AsAAQoqhkVBUxG7VJ/ioF+z6fBSIl
kS9jxNYEHsDMslUOMNRbJ6cQvZJxwu8vt9yek7cItjE251SS+ouO1DjTOA5sQfak
zX2gjIphv2ZRd3fy/EWn3+xJB90hZD1aq9iLNVtj0LYuRb9DDp/wtgI2fw39Asi1
18T/7c/RbX8+O/h3L41UpDPu5qfwgI0TxYNGR0IpzoNhcAtSLD246zzQvDjOXi1c
zbJHlQX2OSunlov6nkEJQJrEij93TBtO5K6fZnY2Y8NgdtekpYjey9eDNuGQfPjl
vXTVJgjSZPQ2QPbSSrph8CstW0tA01vCE5bzaQl2KeBMAsQbhGZQRANP01lNlsmP
V3wgUTbi1uQYA554va3s5szsYzTdOx+2WY7Wa/q/fKfIVuX/HmlAPOVpgjPerzfj
Lm9XTGZ6lPq8tghPHZ4hiqjg7GGnooWJqwza1daVY5+XPiVcWRI1vhjqRIiLCP34
Wv+sPKqqr27g197ghaTAetrG2pYGc54pNiJuar8lhsxR3yeHJMh/5rBkbewaaMf6
Tiv5J8/J2XxOVrLj/z43D8hGP6lXQsVEQcV6jzsEo7IHfOCxih8jC2I/ZkSfVTWK
w1UNnpVGJ9ZfZqCrTqMnKJemIdy1QIIpuktDvy0vzkTFKCSGCxQG/pJJdlJy7nI0
cM75xDu6pJOajE7rkfHtLbhLZUXqvQBEDjpw6RnvfeWfaftDMg63cEUpJrx7S666
velANWi1DccBV5hsaB4L4Mm3BRe3bxEcAfdAD+NMm4JB3ehLtHXAv50O8Lau/c2t
CPoZcNpjgbpgIavLBSV25IqrVG8yVUJRUZVi4XJWKxOfsBymMo8puXLpPTjVOE9W
8F6wLQkakpc7X8iZzEoQulf7kw2odgv8h6z+OWHtFSQmg5obDduFZM78kwW0HamU
b0vPQDS/qblRzqMvym9byGiBQzl5PzK8BP3RUSzDj3H3LOtaj5cFim271CUqmsah
ii4cT7H6mgMQBu80EsVJWlmVDlllkx1wA8C1iVGvY3lksHY5T9pCpLVesZqNnFOE
pHH+mE/CrCEJ6uHk7iwQKN9fYsVdZtdRl4Ly03F6u3jO5nQaPpLarw020jP5TMBO
fAAZxAzNCUy9NlXqQCFhbH1wBNDTDSU7Q2x5aNDHOxQotv29GK+B3VRDA94PZjx1
KTYDB2ZExd310Qsy7uwwmcEzLZ3c7msOmHUJLZm6wW37TjLWRsQbJyE71za3s/AQ
WZ0Xva1CtsKQyrhQGUl3ji+StdS6YvZBpjUGYy28CAagrC5BDMEGH8mE/s7wQOHC
nNx3KzGuDST6XetLAou7lr80MtPrKb6oNCku5KruDpQvmoKP3cPKUzPCuTjWkYT3
o6XOBswcZ+V1MIH9Oq+fZVaUJOoV+pgeuqCE+r9m14TRMLxAKAz867S5A2lHV5WY
s9tvLTq/2Hi209nocjeKhu1Rn0M/jzwTJPSTyNsWvk/4XNH9lVD5T7riHOBTftYp
UiX+iOITW64HOgXidK2YhKBmRwkQXEzbLZC4XZWbU6wlh2axF4d17TmtfHKN/pNg
hFrqd5mTBvlCZJ9qRbE5qmda/jCFM9QV8QhLUcbZGVPbigoJuZ8jZukWUEjvtVIU
PrRLBS6cCq2NIm0GbTrzcVfOym2CD6KiRJaJQqCYDVoAOh5hBpgq5CmMPewgER6T
52uYdnbYGgv3Q8rsBtxgimbDftOq28ydfXaEclglDEBYZcZILICwgzwqOv+HwhUP
aN5dPtyTnXbz0hs4ZnukD5OAFxo/MkbRNKeDrJYRFnidyYnJlHqOKK8iaVlOQKGi
zC1gSwhGBN/NNtnCBf4Fnbe96n4ukZ/Segl5UOIIwVN/evz0uBaJ9HMN1HKeEwgD
Wuq0BlKV2jKSV/AUV0IGLZQK8hiM6Qmt70OH2Mq8Ik1evcAQ2Ke1dBVIPWhwA1vp
7BYDD87k34Mh6CL5iu3o3UkG1hAEM9QOW6drEq+eWmPHhkHcz67t3GqR0vVhXOzs
1Zgpz9I9jc7M/bbDV3ZVdkm7+3ILIa37uJG2uz5pumfSR1O8NM3Vrb1g1FTZTlob
vuygHpheMoLG6D3rxu2Nq/mBg9yC2ejVYjVYjPyW+3ZjpUyG2ZjdtvZJKT7gUCa/
eDtP7excSBv3xKi744SaXCbWmMvdhkQvFZYEnhyrl4Sz7ZhEOHw120Rc7+gv/tGK
Q+Ex68RhDaO7ADiDwI0t6cSh6McVNpPhRfmH0SpBvUR3qsphPdSGwZSY8Uino3X0
v1qHCsFAkIdyn0Uigrfx9eMPukhfHy4CiXyV46WIfrT80nyOZbNwulHsqeYYdb5s
5gZEI+X4bxjw1XT81gi6A6R2a3wTdJ7od/zA9ZsNJm1YbP1bQ9/dxrknTnpbdXVK
hC3x9gxi2Cz3IY1wveiu4sQVY9LjscWVxetq5ARyT+dFCjmg9JEHGN9givr2SSdr
60qVgcsuRIovSxBzIZULls3N6ga2GhVSV8oMH0STLkdL6kilPJWAgXJHY3Y807t6
LRWEWPU1DwlOAPYZrI0Z8YgUW2K7iq8MWOk4YmVEYk26tp4yrsoAbPu69Pn7TBqn
XrfSokk4HduZ4aynUPLEGrl28u6q+CFjWi7uh7TUOAmuRLtlKeduBnTdLfXzdk83
X4BPWiGNeDHwXSifBzvpFmw9xQ0cpNz+Fo+HasICJa6OJB/BAqQaVBCjY07gt3yR
MdPSACkogKYSzlI08/BLlvAx4ANASkqoefneRupCyiJrxC35Pqt1rsiwFGGYMN84
77u71dRSwjkju+QxlxRXSpvUHDNZh9dGnOROm+veth7jaurlEV1ogGPx/CTyCJY3
wyM1Bvdyprl6BvZeNiCSV3IOYfuRrymLkc2NMcmmmykEAJxkRSHzWYldQaZiW7fi
8u09VBL8Rnhu+GbSkEu12xFxsbvrYSzpuyMEL0BnSZfxzQNS3nO3eneo9LJjHUF3
RM4uS5zIFf1dWjtgJ0JTHzAw0aYf124h8p49QtN3aELgNVxVjo7+DOIHa5REYK3q
sWTO0bRutIgig/79IuPCQtMhDT+wlJejpMm646N5GuFJGnO+fZ+A4moYBWOA0a7m
yZESoARB/Z8e+pEaMqQmlq4o4b3zvrpIlvGblf6wdDEIaUFsoDqd+KB0heC2UE0f
28ZzXcCwZHNqiLvwp8hukOYUEh8eFJxbnEiKvqKPqrb/YtTkCJtwMREv7d67TPv6
obIcq0iW4XGKeO3mFeGWglaKHk4XcJz+n3KOZ5MpfsP3a+jyqopOfxywdu+g30R0
9H1Fb90hSmh8arp0Jg8snXy0kfyO6mIN3+j1H+aAoaVNe7bmzfoh4eOU9f8o+i3M
gseosMfRTZE+ufipACAs5fk51CVhUSNzMHz5l2kAtVWj4M31O2wGbkTskM3dFcC2
QP7UHMWnQvvnbw4irfhGVp3PwQ05iybxsGjvRj6xH0grS83kGenTYjq/Y0B2Wkr9
/FL0qSvm38x8Z9MS8vrjhqgEOL6CjqWaOhBQnQfjkuNDrLZtxWpUM+DviKhnJmoa
TpwYxu9LpEmQATP6EUxrd9Y3kx5wBwx4WDUioe+ILHeYnhijKvyfNoLzcK56gepx
m2VNXEcdyee6hMFRXTjhOpOFwvDvLesAWfxyKbQ+xxVTNoyS87Z6Q0pmJmSh7hxs
Hkk1O0L+tz3eUvAJS7fVkBBba1Iz7GoRUAj09LssQ4l6ES/2ejaPWhmMYjhDSxPM
5nfTuCHS1arJymFs3WstU2vderwnBW8Ou9TXyVeQW0WnUJfRR/2jYgzqLEtmGuPP
VNTBsTCa2JQ2u3tsz7SfbTudrLkfbOlNbmjFMlpp1UVZX2RNH4FlyP2743Q3ONrY
yLdPVQAOT5Fa/wOKvfCtO4O2XA1PRIbTU3FU5Q5tgc9s9x5yUOyQb+XPcfpTZ+87
MRpbwSpt50aR9VwWpzrtsjmhjjKhhiFRObzFWTUNAa7QHlWHmWt3hKbELFBrmjF6
rNN4xEJnoEcFqIx5nJuwDrtX00ePFmg2kjocUEzZhe7uE1d34NCCbLo8Nrqxtz6X
thSaQtMe8JVxr/3CkfgyKfpZcabBvgoG5MPQsSXvOAwrDgMKPX67SOR4qYmNFXF6
N84f3ep8x7VMB6wpE6eWmXJZgyeZEGuGsYOtPBZmGa/8/CqTkMES7IFtP1RiUpDR
sJs5PlTDyGZbPSeu7xk7x+UpX6ZO0Eluy4Ds4yd0uYoOmnTBoUVkd5B3irwovw9z
du47051rYQFh3lSLbGhjsk7zJmbs6RwGWHSJtILOQGZrUrlmyUEylSGNmz5+oX+/
OVr/ZxccUJiLwuQ9kczPx9Rv6VkCWDYkC6Nb8ro2FXhd3VCm0ZFOCv/Xnf+nOCVD
pbJoG0rEjFcX31jGbTBmfYg//HWXp8sKO1wd4IDHy+g0YTUflUG3z7VukiSoqdxp
ZQck55h2vzFJJrom9VX7pUrmb7GJDT12K/G/TV7JlzRC+VunnszkXsDdtHQOaI5j
w1zGlP7pRKKoBsMt+oo5kYF/lfAymwbxWBeo7Mx9wt455fn7+YbVVospj4EXkc4r
dqeCtQ8Qr2jP6dSyUshfSfHuh25DjpxqMALq+sxX6FepCKBpg3VNyeM9LuCIjL9Z
HEBg1A++0RlThWo7/dE6Du1fgULbmvULNj/EnogFj25DSWW/uah9bBWVvFyWf2Pn
Gcu2j8dtTLnKvPZHE0DAZp061LM/6DGA7yWDImMmJK04yvwLobqjXR+OMLg0LfgL
RYJbjACqgPdPRrum5afgP36jNEk/FH9hpXFGv2efKMiHlVbRGlXjx2dKiEs06koD
HMZ0nQHEiaJq0rR34HathQU7SUUtm1c/ZS7cyHItp1SSZkSV06Sps87iWLxYUP0z
X/c6Hfd3DZbQb+3Mlh3yOggpacNfgqlJQJOshXooBudE/eW9xG9Imf4Or/lxAZ9U
7kEj0wIVIRfIOWtdaOUcV5OMX6sKb93ksqjjn6JK9AnTa+zART+ozAFHB/eYQTUG
BcUN/8pd8RDuL1sSmm2JXpF3l3WIE2HtUMFnxHQmqhvaQIjf2iluBOPYettcN7ph
cd+dXm3qEnnTHi1fBLWwYZOObFFWKApwp7HEg8gSmUTCCZRkFxpfZT3srX1oIPFT
YOZtaoHhg8Q8TruNq3/5TjqYZlOp7yKLhw4XW1Leh9k2JYX/RgnY0A+4lTaOw0kw
tGUVEHErsdE1B8sF9o0DXZy9JSPkCsSXCDe7eGLBX3ZYODxnUonAtFyImVgfVhzS
pvPvtZVkCvB23icjXr0XNVJAGgF8QcP+YrX74bV/ftoifkwRgvAT8dwiWpwQM5Zk
LD6b822EwiuiC7T/kS5RMYbE4AGTU88eUv8i6TRUirTWVfAGNlxbP4kj0tuM6oBQ
6CDpHs0wFDMr+1aqTy/PgdwK0MDktlbSKa5Q+AL1SiGGQc45DrYpzCMqMRWKnbT0
0njR2jf67dm5QQCOCDQcN1PM1avqRquJWluwNSAmwMkV/pbItc2YKqHYgGLjZ8HV
wpvKBjXQzhI6eTz5ZvkMWvjXTH5JNnQAOSqaf6PGDsgtyG2NiqAh4mCbFow1JTbZ
kDyK/BCJ0onvRU9UK2I2JCObAqdE5PgnOY2kFRqwCUS+nVuYKcHM+OltM4mnAOb1
ICg4Nc0SOcyOKPpyjgcL6JUCR7xZYhLM8qIdbcJ4svMxuEVsKQobH9EIYHwO98FF
vcmvAPfCIAVozOWTGdVwFCjJKMJpvpeaRcFYS2r16FE1a+/oaIzcDAEBUjInk4JR
TQMKjxZfA2swiTOXrXXI+yTFzRbK/wFsb7swZgoWatRAGiYncP43LojhwDK43y4o
iNQhmCI4Ks5Rk3Rf0wlA6iTKcBLl7HYpVsij6+tkfl9n0wVsbK/9erPmIkpnbog7
1I2HnZcJMfVz7jSkM5oFxLHMSgzWU3qJMBLiGZ0tdWNCkcftL58IENOUHA6F8w05
wdESyrrfgP2at3X6WqGW7LFSmIGurpqe9LxmclLVaAuhCGpnLabkjiIJF5ryNi1x
0N+eyUbPsHueuFqM3YQgEEFq7Hycs0DfXHpH9gxo7fCWB7XoKrIVfuzPs4VqHlDU
qVeV7YXtOsh8XOCC2RZH+4Sm8vlV2F9Wl6TnRbIIU3ppTvVdgnZezFgArM57pYbB
be+OtLno6nJe27lF6mth1nE7LB8rwt3AIJt+1oxRRo3YmiM6nE3bd5xN6bH+q3Ll
oZTDp1zkJEqGT2kMnAR8OWem+/DSPwM7Lm4WUeiGwCPDboEzXkFtFW1G476hNJXd
ulbAPglf2CAIe+j4SFqYYh65o7BqSsRcXkxm0cRKPmdJbWa5G8yBH5QSJiLWnvpE
joW9HanPhmBw1MnbUp4sagCcepszNi95vgl4QnACNdEetNNH2DU6s4Pn0KU14YRd
tgzCCcqyFpfVOe4FqFY1p5K3O17ERmf0DqG5YsKY5l46S2dn+uKOxgbBTTmAOLfB
o6WyjZmSt+kr0zI56xdPgSoEcT6iUyZd7a95KhA4zk2qOjnniSH6RSVD9F/5U+bJ
1Bb5VwDN/QPgaFogh9f/8eTEm5LUPcKJJjy9DtrWN6vOrFDa2lWgkEvurKmRM6Iz
XlRJvU5EerLR2leN9hfGOwk/uC8+o0hyY7KOAQL2Qsmc4qipSwsdi0SbCXh55aEX
gvCI5LRho61/Kzh6E2ceAJbPGrTaJ0ozpJpft80UTZUXO98VWNf9b0uHWgSV+dHo
EoKOA5AJXxNBsHXci4Gb1msGUpRqFLomMt8jrocAjARCrRMNQ7+ymxpMWgu6qGZR
ZmOeUv12lcbT4Fcv6jxcrGD8OMD9GbeWLcjEacl7Zw3MUm9nNOIpHOinmGbLxw4W
inrhPisezC6hI/on1PBf7Rm9rachOT7OTd71TN1VkJK18o0kjNREMTApkVRe0kPn
GWMmHsGG4rp8/kR4YkhYJF1eTmdJK+g5MxAUFGoUQEYAESe9bKJ0n80kKBys8Ce5
WT2uYVOxEvjfHY8/Nfs34lKxPYh6noQrYGp5WmKrIAAeBATc/omsJLAQbz44ve+u
fHRXpRDZVtO2QN52wLvXYHg5SwV81Bz1PICpf0xNg0rLsPu0TbhF4ivynFLaW1LX
H8Cy7yrtHZotaVNJ6MW9cMc1eFewuU45uQnzLFzT84rkTlmT8pgaJXK0RbAuSiOV
FO5xB6VWOdGhHBs9FWPfCi1Ec/uqJq+q3HSSETiJzDyApDH0N9ynjEPvLTs4khNx
2XNSOpvRyomFuFDZ6MWhZ/dKIT5H0R/vROnXUaftRYbS///IK1CWCc36y58vGMVf
11an7oPylQ3gqtiuA4E2rUu2gTqa8mL24GmJxioPzqpf/QyXt8JOy6n2Vcw4FYvO
5E+QhLeQ7gNWgMe5JHvVqBCkZ7G6l0qo8LyMWozoi4JxAe6hGT4c5wtzn5BtETsr
mCD9OkwAjVqR00fWA9p929z+pVbyQoq3zPdVCGE0I1KjmukMD5NWS256n0K6DMiK
Y5flekEf0VT2DRlBJp/YEXVBY/V9sEQN0rehdSC84xD6rrdeApwdmRLplwFVdlLE
T/zdx5msSxcK2EibDOWTGUHwJxJ2osDqE7Ted9/DbwoxLA8Egux933tPaM8Q1OG1
0F9gyfVgXbZXfnHMObCQyzV5RjE0q8I1qV80/CboYNq2YfQFdILL7y5l6EcAIQFt
CZlsMGry/UWoamwtbUazVq4dFPOuUwzoQ2pKmjUsEtEk+whJB3aG7qsVdf6xfZc3
g8UA2iiEvT+ZuX6/LEgf3GTtWrwcdPewTR/9AyZlCNA19+P3QHdsA8GRmpO4+ip0
CPHXubVXODDC4KUwX9oMo3hQWmOGhmKo7UfuKxtRphZnmJQ8fbm8yqDfObdTUunX
uDO4TIoT7j/vPLdyPpTlGBQpNLQLLCFwNuI0CeKa09Ghag9oKD4XwEpaWshOVyv/
EHBj4Oy1oiXdb1pmmAKkTNYGjHS0sgL39HAGmtZI8zCeSUMVqNaCn4UuozA3LSKk
16yN0j7BZ1eXsNyX5WLsqv2KJeeCi6diUVdUq7LfPr5W8ttKbZh7d92oACYVxrW8
v+lM8VOrYjZ0H06f2IXH/1uF1dkU13K4dgU2NufyvBl1TMRDV4eUy30R2rqv+gLB
A2j8Vm6Rqwu6z7eNene6/1BKmXQBBC7X07W2hIFLfGB7JpOxtpXHjOb7GxDIU0rK
ZmVb8oxS42xUU+VJfQeenHNUX9PK2Hg2nQgnZ/Dgg/2jivt6wzr0Dn2G7wWq3Zgz
jsNvmX96so0pRAA+z/cXF6CPcBS1Wgta4nlN9t76JFJg/rNUsvUsIk96IHnvnQOp
/yz4mVE55m2qt0PPNojvJXbRWjywc/Wt3GAiunFxEaROc3c/KF60c8IJFeK6cXmr
RwlseLtmdKt4rEYYgrewc4eu6TDpyx80rLZ84x+PIS0+533QR5ggt8QeRG6AHKWU
ywtUBzUOjgzKiy8Uv6sFbXIiZ0TxZGO5pU55IGUhZxwuf8vmllZyrXtlCtJtLjn+
KORjjglwbJbWiSMFJcKEgPa4Kv7lZF/E/jhJAhMJQptXnKN8lO3qKRCcd3li1AcJ
wIbmS6AmBksRCWst40F2NQsM3Imnl6JFFQ/UmNCzMDX02AWU6MJIkst9M9qp/xgL
ueXpGwDGTitUrjo61IsxyCOxCHxa6IjHkkFk6I44jvXvOP6fCsKfZTULoWxUQOs1
J4qfdGrduyHgEUz9gKXbRoPrHO5T4ihR2KJhLY2/YoGN8A2clGX2nUgh4qk3wWqO
BHRzIdfykq3oiGFsdjvSnPsWrctdxePE1cb7F70IPgD2mgEc5qZNi4OJxsBbZO62
Gr4kt5To8rX2lGm6DAbk8Em9Emergl4R/o6ZNv+Aya24O9DUb66YCoBFMt6o4xpO
cAFPoJEJ0DUHk+03UJEXUHvb66ffY+9w2NUP8+Ltf99Im+2RG3sNLoocJR62rK8x
BvWmZGjiMw9JQu4X6UhCh03XiEUNui0o9gvFlFrWsWqWiV8/5nfFMK4N9W4FLxsE
1nX4PCgxPeUTmF9JC1ni+Tj4gBlDhr3CGJH2pm257r2rRAAnIkYwGDNny6HWU59M
us2OFX4+8mEL0YBqLFE0vCSZofEfXexSDwKFJQhhmtcf56NgZlW3clUVaFORytKY
aJU9sO+OhBdL1/jBIOJwe6/saJ9zWJig47FW/FvfiTmtu8B1bgMcyRfwmob72C8o
34KJ92GkcVnO3EhZyThcSfJWAf7vdLppNmsFEFHZHuGl/Ew2+c7SYLEoJbcq+x6/
mi+qL8UHnIbKqlN9wdcBYP7jDIAf3W8ycwl//T8MtoscnyMdhSrIlp9mJsIU7Klt
SBVtTOyd0LweXsBPOasVGJWN1NEluqnFHmuuYsPpxyt0hP+dbmprD400BZu7A7uV
f0kqmxVGrYma8f6qJ+uVL/W5GNUxF53JoZrZIIDKpnLE1ArlTcV+TrFujzEy2sm4
Aj1bpz9pIImf6wQuYj5amYfSNNmVEQR53HuXOWU1PIZet0BqHi+FLmhS+V93x5hj
qnYu9hZDtPIAgqj+32kPS1hxeGJl1672FvE8CNWMC90+YusBThJ8BXlW+JY83LBg
8MpNgjfOg2ML3LJYukWc3C6ZgpWHpwfqWs5NsyBBkPVBPkKtsjnoXNZXK/bw8Al4
XVHC9GLrdAF9+EM9/kt+tdozv3VPk/3GvjM5ya5Lh8cT/JbkoRrd6N2YHlYawyic
JyPtDAFvb2Rynw6qiWMlZN5OWg77lz7sVfZeDCuOuiX5KsuMTgcDbMx585dsk1+a
i4+/iT4bZ+urx3fs1WXtVuNtp63cg2ofV7sk+1wK/0uyPThEtq4r+4jODhdyddJi
SG1i0RXzyM31Y411HmmBrbsD/BJXzpOyaP3W9LJ6M4YDCQoPnzeXDtgUlbT6EE+9
cYMbSibdwSVQ07ygxJuOUKTOQI6v45stJhgGCcMa3L8mDH6IT1dCPe2C2E7P/xTv
RZEZsY2+f4F8J7ZzwpNZysTp70lZ0NbP8UFTkRJBdtE5Cj5PLo/TtLRzHWRhAJ85
mq1yFznl32nPc8DtFpioJFAa+MFVjFGXN7jbYbOl7uSvQBgbbdMqu4YbqbgAkHSK
+hXODreJBNfPgT55ea0Ut7i+TOiFQjjAPjz/8BR4nUWszJZAL39pwCI1nTfp668/
qtqqTciw4l1xMzkVQDH+3ZkRtG567awLH+wswAyaf9azqux4vMXsHO0iGHqiSwse
IR+5T5WyWiQvUUR0V4yeWuoBWUt69YOsybDXcS2UhChclCak+CT/v9baI4M/Es5a
ddvuCoOZEoPZRg7vTn4ZtH1GoL+Z40VD9BcGNO/z9oIEh5HF2LkmIBHUaaitWisJ
R+5w6yZbNfeLms2foKZYutpHzr/CT7C82dvOQamZebPWh6ey4uNyPxO8Vj5R5nHI
ZkfVXIQFO008KsAcTR3R9wAGA2JsPdlbpFiPM2NDYfhrd7/fv6/xl2cpFdbfydt7
r7NZTYhOZ0GpGL0P9gABI6Y6MkE4JIWZQZWGvLGGjF0ekI6+hhNZPahU2jTkZ0vc
slDU0esCvgkKFWh7WLxfOBeiNc1Fhjgxyj9ZbyiOz2LYSEgMqmbkGzWaM7Sq4e3J
RWmdIALJOut3gDOLJQpl9M/xGSmhT7LotcYxbxjpA5yiFvhIFv/EH1kQnqGKGAfG
uJ9SqorQ/ZmZw1tDXVD5DOhCLA8cwhNAOODQsB06szz9iqRQbsu3hPeEVpuH98Qd
UAc9s8skkzdIxz1cUNT3IWwx0NofYNz5oUKfz1z0QDHxLfOAQf1HqDs+njLPh7lU
B7veLlwVgwKbh/gs4z6XE/Qd7tq17z2VU+6uSK8k5RJ/Ktyy1dg4fJZvcN01076h
BfogQuOOUx7dIG7JSGerms89Zr7vJEn3ivVJcmkbGlWpwptbTH9SaA9kit1e9cUQ
ci6OBv3Tr5ohiLtmN4NOocseK50RzdD7F2Uuu/xwZeNdYAGCvhAlBNpJc9DWNdn6
ZUk+nZVgg+VoDwgTItMsgnx0kJ1VMmStfHyka7/cHHYidGtZ5gxSp59YqNywJ5vd
/OEBikiIC2WUnPXEBGkql6SzN7hsbXzI+9ay8c2NX1RNWY3cpLAnstWh6BXiDBoj
DdZTRcocVc0cAHSUuwxaDy0dRiaYddJOjYVcaoY7n7jHNuxYRoy+MgiLMbJl+Qg1
Bprvo290fmVXBkMPnggUWgtO/2lYm2ETgPz86sum6Ttt8SzvDCNOBJcevi8jL4HA
W/JqNomKQIwxvJab3NauX3p99HSnkN4jdtjU7qQvaXjobbpeeUh6fUri0/IQ3UhR
taMad24n98E3vsgEL1WkE6EmWO8vLpdHGK40lFztPZ4kr8tqu1hFucOxC6+/QBnc
EHOcQUMkKA3txnUBDZyrmcElMEHgA0xepy7Cp7hqVzjctS7Fedfo8StBBa3ugSRo
z+juvd6K2js20nnskzqlADe3yro4D+iU1pMEoGAs/bpFCyszN5okmsfM0A1kPQLV
RnulG9pdfo2GOV8SVeLymEJpC4xiYcyWmM5ysi19pzc9SHrLFEOCnEtRZ+m8+Eou
jEvllVfQpuxPoEcuiF1Ha0vDmp0iXYjqnNXYdmuMoN5sp5VFtqDCopoYD0hm0jS1
/B9LMX5fc1/NdX9687bFVxtKYT7qcTcbNzcXKmqL7PgM0B87mmGtXttJ/5/ydb5e
yAwGyb4yQhdMiJRkkWhq4ynURi2sKkYYkV65lkvXapSbHFnV6htf1ao6YUTQ4W9u
WoeoDf+4O7fStzUkiBpV8et+QwQiIFyesAjWNX5vUmWWfIAs3+xDoGjNuGQq8Lfo
PsIfeTTTjlU39jx1gKKf3Y6zps+mifiL9dc/AGfoduh9yws17C/lrhtwsPxQV87N
+FpBMCnyH4p6ScjjnAyag4yI63+t5cy6nM6s61pBScF85AWkvmBzoNaBDzeazMhc
+Jv6G1FJ97wG4l1TC7dIvFyJ+JMNpfWu2jcsvczoUfFEKawj4DPReAs3bLKOPEaM
pn2LxBVU+DMEcY8EfnAda7JXqgDNjq14RSocYK+UsHnVS8adnW0KWJf5SIOjzFg7
qdn77V5f4ObKTmny082YE/84Huy7AfQhpQP/04rSYesCWpLTgZnBoDNxtf+a9XJE
o0ZBA7sc8crW0cbKX6n/73xs7j/4kwvP4n9Ul8d8/nj8yk9AUka4sKlJLkGstSGy
BP625zEp1qK7pi8QuaBycQI6NLWRB649O5B7byGnwkMBbAzvdtNH5cTh+lKro3f1
GV3ViHVPvHBLJV/qpQzZ4866OmZGZIVEqnXWQfOa3dDed6fvbDFGjRswlCyHBNiK
Y9UGiYdeG1rg3ydBHLXm75aK6IuEWcOrDiVfk7Jm6ZA1R2JKrGOQy6pcBOd2zUlP
oH6Pk2O8HbIgCzKozJv8N4ydS8d86IkS+6JLXFRaWzHftnl5BwOaprM2OxGD92C4
dHx9dHVr+aMKclR/OAzMHtTBgdX5LBkzypLlR5Wz9OYn2cb75AH6Xalyd9ro32HY
f3u4mASwYgw9ifnEdHW3VL8W6lRORFo+rNFe02zCXgejPKM6X5bGCgBCWQ09hMHK
8aAIbhbLBMJ9lsdeliVurKy4nShWAelsRxRKCuCz4HkCP9O/CYGiFKG5OrMqamkG
/g3uvPR+dRfLepVrjIw+9WANRiZ4u2os4sKAoLb8Jacg3OvHaRIwgNT671qMnRed
2erfL4ehNnJ3bzWrJK+k/te7yJDwqiIvW8fnuc89WjWwKKNgv3ACIUssqgWAaUhD
PnaEUN85Pai54GZhEwVlykJ6wY2xjzVo4HO/NG9S4/YhlY6sg2BBsW0MiLTlCotD
+EGHOpwR+Kp4BM7fnWiux2pFTp9ywuOKYngfPuuX88GHThs7lHh1d3P7Yp6R8I18
/G1PsejIL/UxTPeZKZr0mrOFjWfuJulMOuXooj42u0JfcmO12jxP6sBHlm1hG/Ic
xmjbd9/r6RzmxJgB/REu49xVW80iu+50s9vnCcZerglb8w8+CdvM2qywaZOnFOUK
xFzjCVFIoCE1XRpxI26OWOtRNaZu6Vp1G+x2q/SK08fVYwKztPHeatYlUMphQW1V
nm8G0c4buhaEkCb1JTYWFdcz2ywZ/ObaWl8CO8iaAEYT1dbSxHwmF/w/ibIo6BSp
aF/DEHUTaQm+/zP2me5aUOQZFUx/WGjFw286QfBieb+CnoeqIN9vLHCBufs/bWTL
UqQTZNzNGE2XckSNW3kFxndBj8zfInwQtD+kBATRATchbU4FGOOZURZEZDsAV167
m9pxa/62FsNxTtgZ/OdOJRK0jM4T8zAqwR1PeCecMbzwOP7DjMDZhI2rCLfK5Tuz
2GifAjwKl87kbsQWoc+aqXEpNrgOReoSfYFfT+cb7lpVR3cgilhJDwSL/E3be+u0
Of8jou2L3Gj39iTLCcQq6apJdryT1wlD2TmN8aTyeTnYGmjNMVhOhaETSkNgOckv
s/IJDBCX2sUA++l9Xx7wU/6IU9HDxhaWeYYBCnqnByS3wAp5DKkvId9du9AR5g7S
rS9Bfwxo7kzXJJ5qFogJnEDWv3G9Ic7nR0qhguuRdvy9uNtnbn+g3xi2AMHB3Ign
SwTgSWMZx5XXJG659ma1tH2p4j2evw5FBxH+tWlZkuz2v8ZRhvBLo51gUrXU+r7m
Y5axg81l9wbCcKmXQMDAKr/v1jBjJSpdBz1tjLRb/Y2g7D797Dy/KOS1AMkx4Rld
0h/YG+6js4NyHkOMsSj0gHtwk0hEBDU4WHFIUyyhdYRZWGzIo6DWksQO/2xgd+vr
3m2cTVAYXNwuankWOAzNLfb3LaeSSdTJwM++Eic91sy+/4BVOYoP9jgRRXCb6BZn
jkJi4Ddc3Dy1HwcfovqdVpA2SjtB/zVDdbYHwdZul4175KSdBY/KyaZ2jOuHgVap
m8C4v+W8AyYT16ljqXFzk+rRqf/1/u+wyb4sS0f722SB2u0VUDc285Jog8LquX+c
8h3RSy+88xkltaNrL7CUJRwbtbHEXZVkdQQB3ODfaSpLoF+kQ8aXK+75UERLwXnC
IBd7ZNNtaT+vtqP9MKtkQmhB4adC4NXJR249VFdy5pNYYXVetjrXLYwBnnrqw8SJ
kl2rT/CQbOkE61n8Xlqnyn1uzFZkUkYa8XzL0DyIiHoqPTJqJQr6SqDwPqQUEXss
gyGZqwFsoKzEMi6BvFa7DiFbhdJ04UgK2zYQXsHZZWpAA8yzo93rB8NVttmpFp2r
QE3xMu4BCOeI0YjwdyHxCmxfn1GCTbomRgUh2dlwTQT6a73yliakTcgmnIOBoctz
2/AGbqOjcCpNKAWCyTxx6YSHeYEihgoHwtdU3k5/dlfaqSmiKtH7WNC0oGOV12BH
hApoLAbKFbk3R5YjMUWn9EjfhU8lW6qEE8Kz9FMCyo7XduwDcGZn6UjOlXijR1y2
pIg/3CUFG4CRLjwpLozJrQMJmtbOmpROLaog3/i0wHloaBkJ30V5BLMzu5mTRBGI
DsOvayatZ6gTI0nW7RUo8bQf4XFzpIMEiC1jw6LiXTHyhWYBg+j8yUtpH5pEwD90
zJwp2eq8IxhM72k8sYwMJ4d9AvsJBUj16aQ8qtI3Gaxppy8Ek0qHrx5CKNvID2B+
H1rEOo8SsIelb+KtlMUkn6z+K+naWWePWG30XIBWlwrNnwy/UZddpNhZ/vpyt8VJ
YHtrznbDbO0CmiqAxP++IytyQ5gaLVGDZTz9n7Y9Dl+jMnScBpIDRzB6qbymE8Sw
fJlSng6zzStzV1NHwL9RFpIK/46VZtvv7OzNVGdNwfZVDDotthSLWumSTEbbVSN7
qiJEaL6MdbMIKzBk9dV+meYACkJLMrsj6eLG6CMVetVLBLp/VMuOeinYPIPdQB4B
30a7QWkuV/a7TGkdfzNWzTjRkKj5kQ3hXnhEehGtTuUQfZHv6oY8nH9oE+7KEkjH
AbgKp2lrt/XKtb5jCoiXjtHpitm4AjeGURCU9RdaD9rTsvRKEMyo030oyqOVrlAu
cavl2oSXhmLsJAlgGJ/139XLTNeCOUYNQDNF4WI+FGFPTM7z2RFBLx+OH/WuxEsM
bLhWxm2JQCSUv7oHWffW1j9eghYFxXFHN2b1HVxw4LHUbiUPZJCBblcKTwVLT6wc
WeNnEb+13QlikyG90vsjY0trTEavqDUiFXwjHmtpK4mf62TSruy2NPfm6sZHjfCf
jvHrEEBePHg59owoMquqR8Niyycl5/QasdD9rtLYeoIhTYl0e6inUGkeTFua0c+k
7E+acNAMgS5ievOXyeFpj0/59dbPkQcjfnp5wRkONu9OCbIhF8Enlw2pl2IjIzCM
Php0Sicxp36bqvMFRxFgYFRhlUsMzgemsa7jBy48IxnETzU4KLXgldRLYny8+exN
rzrGTqV+WDdkwXiBdW96j8rLNS2FaF5mrVWkPhoeQDkQLPS1pTqYjmy2u2PvGWT1
YEHtqFRou+94Nsvmc/QjYJCqG/zkR+3Z3g5jzqDMyc2N8cjVQ5C6CD3l+tjQw71j
UlmHigDhusQL1NE+zRuK3G4yfAlQpu4qZXPUs7ext6OtRn/rpb3LmuVfpHfHygYd
MekFPDQE6NgX6lTlYL7pNXdPhNeL0b2xaAhJvXfNr0fotogQ1jBBRZdJUTNpQkOx
utQvVV+0M+wvW3gMKZHjQajSDUsvDeNbAuUlNehswupZ05XY9x0Yd42sNPjcTLB5
JFc11nR48ixmIPLUdBBYSjU27CtZ0IRteh0RT4peg2py3w5MomSW3DvnPWIQsW0e
LT1SL67YpIXC7kQlIMKTKVNWYeVJDWYV3WWl8SLGYEwT00rurcukQHGoSnKWpPXG
gRfTYgvMbkC1rTY5boo0SiIzQQeBUndR8LP/Bm/sFzLlCro6D7pfh0HyY1+f50Y4
mbC5G9Q35/S7FTITXer6tyNE3qYan7guef5zAQ0ouGuYszjSAHj0MskCwQbfwoMv
V6lup3ozdL82iQnS2Z3qn8x1ZW5rVFoWOrqXXOzdoW1upaLjXmAku0YbtQOqCmzW
xURb8W5dUk+Oqv4UZnw4xnZckkWGvA5J0mzUUcExc3CnYrU6OZxDgKrBxvV189rh
N2hISnpbzBMiwJ+yi6atdqKIuH9rjNELXsKKlV1bVm70lVJRS3coiOKgYa/FZ6RG
AUuWPjaR0j+3HHBQpYAuCMfcg6Gc/esPpdDkS2gBUdW/8VGQwt+dDetD5jcXvIsk
VMUQIeWWNo/qkOZPH0JpLQFlPs3SPh2+LsPuefyMKnUyXv5kMocr7ft3Tz7XcTOT
WlZTQys9M9VARjjBQ7Fip13QmTY0gH57TTHrmeks+cNyh/YvdVGpFIIZ9h7OOBmd
nbWaAR1DIMaIBevse0Ih+OmUO7FDTUSl5fgMrHfSFY39+k5m3+56dk9l34kZp1SQ
z06nTNUg05FoVTMwAkN72daBrlVTlsdKzh2vdvUel42MgQI93YP4Uou+CYzYZLYq
7347Teb8KvTFbFJrxWj97zA0a0ciRHp7HGcEIibGSLxWBvcN8E0NOKfPQb0TTxem
mG99jzM4+qUQZ5iBFdi3OLwDoY0N3V+TYFih9r0GU/peD24s2bgSL1+XeqSC2qZV
t+sDIE+6UIgKXas6JpGo8JQASqORrTLZ9BK29zEIaZB7l2M32mDiZLPdK3xfzM8d
b6DKwBXW6XZ9b5ddmmO2idLiJtzuNoBIWkPkMvSQSKWkHf2h0Y/prCT6rqWqz9Xq
Tjxjz44bde1AOcPHQKqKPIpKu1Tmub9btu3NHj/XNWq5ixhdP074UHt8mvct9moI
hrRNudcJMEDH+reHDil/v+ZYcVRUc3cfZOdKQygw2uP/PQlWJ/atsydqSuwT8c1i
r/j7uqCqwmKIKsJ88SGukV/R/Pp2p5BPPHwwmxIJfANuQX1vHyK8RaIQ7VRqVIXA
TVGL/e73KaO1hFqAKQGHpDDErhKGCukmhuNvNR5vE5WHeoujdNn6N3LfbnGs5lp6
0vLo9JDc+PrfeWDcVGpSNNj+ABfzaXwRnklNJWpEGL0GYcpCq3EB570l28uA2LFE
oGY57Fa7oo5XpkdpiDSKMdKUiN1r4wk+S2Y/PaO38brWvFAuYgmJFDTarrRSZqsW
FaDhZZls6aJo/J21RjO11PomJzEjxcparTdscjM8ucujdERS7dERK1g7Es6O5WJa
trNScNp7sVxm35S02mYwaHXyCohyAVi+qDoZCLzLGaFd5yrWsf0BHKlNB+ZnDKUs
MTohq60AKAJKfiJtjCWKNKtqIteVfVI713vBtLVbUHPsyoGC6hfAK9vQcSLfXXPu
j0+fadIhSMLGMKyqV/0hzHC82c/+Tyt5UxztUdIAl1ZU2VC5rUsRgZjYXDONI5u2
xuurQ13x6Z8uxCzStksZtgf8TNvSE4fS7+R5LvUFKklSP20XVcQZVtaeTATSpeQF
dLfeZCEXTyQe8qzPE2DvoXmQIr1Sm6N3nHq2GO+CDjTW3W7RQLwpBeJlsudN4Fpx
sLd8D7stE1I9WthCLN8cNXn5cuCCjBZlWYUoTlFSF8/RZ2MIUWthtQJmDLlwlDxB
3lUVuGZofAD1u7MfUiOCgsOr5/5LCN1LDc3DNiLKv8BfGaAlykASY2XlBbN000aJ
9OIelbJD3JFsbnqEcKnLC73cdJKZYaCuUqg4JbcM2u/Jm55XMYBuQzmhj0g8tDkX
FQeKx8uvoMamzybNi36UmOeWYU1Iqh9v+TMDzmxQh0WYhYHidYDLWBcojfZmCG71
H2e1ZLjfu3NqlTL8LEn8CsGiGTmvLBAQnBfKfpYe+8MM9YEc/Kp1M5V9LMdQS9FT
OpTyCv5F6FZ0GFX6wa8rjaEqmwzhPh3D5t6YZ6W0v0+B11sW+Z+xf0rq6l0mR6PJ
xMMwfdKOaay4taw2vPyTwe6jjiHEJr0kFL7avqcUCtFmBmEI5NFVd7BX8ClRd/We
6tQafuCIfXnpsCQhypZOfuAfmq16fiwBPglMuqLQUYnoUhJrpBIuGC/zetMnfOzZ
G6tPXcpdjKk+uVeKpm99P+e/J+gP68ZgLUFTNa0POVRhUu2k3Px/FJX2XKO0Eh6P
apvfozQX8vfHGzouDNFw0ixqRGR5ICKtILJ1r5hZ7QDZlWJiHu3VvXxSU9c3xyuk
/0+0NgegIdmeYkRzxr7/z0Mr4t38sGh6zxmJUO/7BIalZPsLSVKwZECx5GHO52Tu
j7jPlN8ZzB6BKZBnzOLB9SCPVXJlJtQsRzb249vbvIosi+V20Fl2GmCykDOhA8Lv
HUQo3jVzN5wgwEU2aKjxnI5x/DYPz60epSiBNn7i/kFJXzXkWxw0U3jp7paYKRWs
0ibEJALh89ratz93lpeiKPYmwX2NkM5KwaU2wdVHhYC9NKWC2JBnw16Gt9iiGVli
iBzTEaMAqBx+3OznkEM1ACIFNRpB9eLFLY/Tkvvdl4YJRRgBoqi1oAUGybkGT7ks
jEOrE8ZuUnN2vvJETcLgFfb5OZx9/MOG2KAQvniYLZbNEsnZiHJfDzWQEmXRHmnI
dtJYITpN3OUXOpZn3eMZpSTuDp/hVvS0MrJWdcvP+KeMwGzMi2Op9cijiQGUZPP9
i/mEvhuHVrFBk7jKuUneitOQ4lw6GjavYjv8C+/ho/KWMflYULbzhB7Icwbqia9A
JvRyLX6gUKGPxTX/h1Sahx04qETNBU8eT87BLIfneQddV/vUhHX+UQu+5Cx/4Wqw
wm2XzpfPCGe+BfUnONZcR9NbZbCeCSFSPizgby0Y7leyowVmjyFbRSOssK7gnuqV
oIscKxaUqFY9qWvNPSOurzH9yzQwLfee8vpQu7rYzNS9GmPOHGAXz5H8MBygLre/
hi0as440ymBvU+Z1b9kUROk97znD8N7/Pv8CJwY7hS6ff3OhwCJzeoUX95HlIkUq
CZfvYvA+TfNM60JZ08OUABjjSxy/1PsL4p3PepUpjzu16+dRqvdzHjJ93wmpyvjZ
tJa/4YPdVS4ADkle6WBI6JI8bij+8JAryOkohYnnffj/JvApaAWLmRvIwxv+V9qo
Vaben4FrQiUFeESWm6SQkA/vMrWMsQHz4Ad9jufUup5ociUuZ+eXNaZ62FtaMq9Q
6dYf/UfWUz28VmH3FQX7dSzCFF5vLxXo6Z446G2K4iUnB3qzNM6kBOzofkIxnQeW
WxjB9b41mfgVmGynmWUVEgE4LCde736pkYlZi15CjUM1ZQ7CvzYz6Mh0uFiFbDT6
MQJoLVAs+ay15TE1oAI5WLoaXL4UvTLouLnnS/eLZ6AyWJ/sU7OTDHVD/Su+7lmT
BDgpud9aOmhKWySxqrZai1OOpuAw3mQ0PkBFl0d7oX7YXd7l87hGuXZmC/k0gQMZ
7bPRuVv+HaumWji7Bv8mKSZO+nAiNnCz/vhRIyQbxgGbkxRcLckgaP9PVjdywXWA
AFO8aDxTMWpd0Haw6OzPMnFzq+JgRwTI6yr91fchsM/TxeWxxdjlaJ9R1F7P1Nos
02Np9tlAIP3jXRBOiXJCcGPiwyRTSVVgnk4Er+jD5ZwrEyyMVfjRA9rKN12jEZXp
lGYU0jTHw9kfN+JBoJT38Pp0SgVXtbq6I20DJ+MqLN/3Dvo1NJ8/Dp0DmGr49i5c
KlHKVbF1BgoCBN5+O+L3lKQS2aCl8U62hZ9py6WEfmM/3TnKAq2iqecwf91vsnYl
nxU6bHvKDmlGELFU8nVpTIgLgHZa0O94Y8hOEtJcO7TCHrHKM6ZZpkCZKx+y5Ndm
6h3e3EofF/vYCcMnhhsilZPN8QybXes6IoRlPGw5ZfWDBEENRim0WsGbECtbZEF7
7hzZbDeCbDTC9zcDoQMPlFm8sBXIfov7zoDKmAiq0qFJ4prT3d4ZBm0QllsqQDSp
W27PMrdP9Mlp32gpz7Uv0HGEevjYBERLFijNJVo2/Tw9bIvOI7+4nd1U4fkk4ySR
hk3Jg+w1OapDAn8wi4KsdBKSlqzbA1wDgrVkNOMhimwAmDHpjBLUf9V01i5W5fpd
6Ome9yr0gVEG+9hVvqLzt5ktV6uOZhVKtW2zG6G90wspDF9nC7FL32VT2pxaGHme
LP2LnrHwH4k+UWOOqHJFVXvcRX/EiDRQ7nyunDTN4D3Q4BSKvytfBZBI0o/HGgsX
L4kJM0x5JlBrvePylXk0eFglAKw/PN0eiKw5UKEmObAmfE42Gn0hCR7ZAQtT0MkN
8sZ7xrUflkSPqGq7mDPX0GHODkIfIb8FDLWh89G8pvr758C4BkmXgulJn3xIusGo
ukxbMYvRHUt9HWgGBw2GtkPFFzlQcPCfGQ5/CHl7N2y+IqhHRMt1Jy6a0+ixUQG+
4SVFdIKZ5AsnxCCXTGECL6kDLFu9sabGqFzGuEmw6w6GG/rk/RGcztp9WgnLon+Z
SLmBUU04alYd7GocVCU4ncx6Bg4HYXmAUZG+pJ/GTGw9jen3jGcPX1yeYrTw3sG5
j/lHs62md8HvZ5qYsy/bGYAtv5jMBcMN2GpWhodCUV14eVoLVOjhR+K4ISIZ0m0Y
4lscbBoyRIR/QQlbqj4+BOvUJD+SK4zqLHwAnpN2A4nf0pUswT3pX9x7HKArTG7a
LW1HsdrPkygmXlCzjo6w+BlnIK5xMJjK/lguyIAJQ+zpyLY52VDTU9HoAoCaEhZM
dQFx93WBeysmt0AOz23U4ax+7mi4r789jAnn9vsZJHxe0Vp+kEA43jw0/sEm5Sdf
WVYqvM6plTEp9QFHbEckVVWT0MZ5yujeGmQ3DlpHid6pAr8g04fXC9vSzeFtEc7e
Y/KrfNWvWQP6WLtfC2GcTd3KDmSmsaXXw/padrbjookevWdX5hoSrw7kmML1maZM
bzujr8iCQWJSvU2+cmOGfqmROQFOpJ8wRGQBY/ojsQmK+OYq1hRpqjOmjMd3VJRa
7gs4mIAH3XcMSgtO0SUQrhlE7PImy+UWpvT3fUrxYmlceczT2IzZxuN2i7/7PRyV
/kXAP+iQXw3vRWnBS/Z09zNaxUIACAcsTC4lSOf11Oe1axfVMfwnXmLGm3qzXz2g
f73KKHYxWoErb0xB/dVAtbSDeL5eOvJDbGrhhpa8I8G2dLBesUZ1Qg4f37qUmnkJ
1uU2jZCi0Ih+gTG+gSBHOtWhuhKjy2Ki847aL7kJpr8rk6z5muYw7fzVxypqCMX1
+SBjiH7ra2gK6avl096QIr6YBmEPybG9KlIXfPxO7360Sya9Wfv4Hu91vc4uRAjO
1V4JH+JR8cBe1/wtCmhGZ+hctYmJXnA8vxiqXRbp1zjwQv9Eq7B2ZMPrfqVh9VUn
TheQOKrT8soYWVuKnxQK1Fk3yQngn9RAz3cQUt8chr+2h748VIxdJ23cjX/8tZ6A
ZW2DAGr0B8Db3BZ7d5w9t5Ok/hC0ytkFEz3lyDfewUGbmBSCunRC/tqogDcIAeci
diG/lKJp49luRNq0q8hkfnJcE2A+qRtgtI7Ijc9DPlOznHUfwVmyF7Gcpka5rUWm
3Q3mvK1nfGpKtZO4xeEAto+fBDGNaIRBB6ub3LxgWFjIQEorAUf9B+NpYqi1DL43
9x09m2ZNOVaK9DXaHmM4S6EF0+xEXcSvXlijPjBTcUvQcvwC4kxPwMeHCJboPpBy
kYddPB3NW8tRuRU2zcH5xQqSGfb8HTDJ3/XmjONYOftlLhjZ/uAON4LKrSSMmePI
Y3MJBBMh8eLcH6J0JPR6j7VmgFaW+Yj3zxXgSIT9d0yzMWR+TLTWPnq+t4eoRGI9
r1kqAvZu52+zcPhvAOXffnas9CGkUAjFJGf4EnByv2yMAshsthyoUMmORXBjFSn/
CqpJl1UA/1/7ifBRyjMwcSU4Yxh1OgADpq5XX680Tdg2kTrN20bQQpub4Tn5cuSX
XNni/Ze1GXG9vPLDBdas0W4ZVnlurlBCCv6rIChWrXPYFLZyVDfqtRwVli9UGYsV
XSu3arESFjZYfzuRlpYxNkvtFweqVobqiVXy34y+n5PIrpaloMdMlr39MEwmPcxx
aZvXhteGvY41txbulbO/J2n4h4VNmSC8+XSvzFjCG/U2lUHfgeqwnOnwvlaTUAck
+cvqgH54mBfTkHgEWUSPEoEr5s6KlzirIN6mPItkdnf8RXm+XXJQsf8VxXdt6FF4
owd9SMdGUU3/mDP4jv+lPnUcWQmp3aaXLzKGu2HKfF7DOLNfnQh7EcRdpP/07opo
vXFoqfT2pXY/j7eZbl51snHm3ae6vMkHmqlx4iXjR1u6rDKEJt6EMX/wUVLCNOCq
BPBftUkr/FooTKsSzLG5g/tOJ6eKnx3hptyttQ//ksnJUJdwY5qW29tIhjvDaUH3
+sicgvtWc4UG8RDP8OEvDEdkEGfl3xqHX4gXSv1PqAbWHNZZc1NTwf0eXQwwNDdq
f6eJFLa7zajyLr5TNVxHBWPoTeTJ7/MJvsqZS2KAWll4JxIA+6LaTuhs9CYiBniO
zyQSiftb+dQn5NaN2V04TwbL/jHafQ03+8XqETu+3a/ZUJM+XLNyhY/H/yQ3Wm/r
3/KE00Axy9xIFEtwJIDco03MquBwVuCrheLZyUrHw6M8iumJg+Ps/1kUKlNLNYrV
SZ1Klo0/jiEP9lZBH+gmqQfWfvkqdTs7KRCN6EUgL2auLpCYCm+7JDFSO0eXInWF
88Kl5Kq2/awbQaPx4cJlMqdTNzifwLWRbI3+Sjzwy9TZ11HeZHOFrweN6i7rXdtX
YZv1JTJfxDAlhvgdnH68cUbKOXZfUoYyP0ETnWZ9Lyoy9jA9FNJFi97RSkdZs/ke
BuQpZRVoL8qOurAhDn3KLDjA957Ut5E1DuIUIj08zMevuynj79/kTO4RCKz/673O
Kz0GW1jWd3iSuqLxVsaX38UNxsaFuJzxnWx+mvFE+mxr4qDWlwQLVz35HkcqP8lg
abPOuh9Hm1kssUMzp5+2JTjh7Ufp4Hvkj9w5n0/d2rfj5xmQOAIoZG3fe0obSHFz
jh1je0Gb7JC/FjvTIn7bq8P0XYgzB2aeh1XwCbPI0gUVf7XC/x0cCXsMnN5ytEts
O4voDmDlBHIUgEEmh4iZ1+C/mhpi/rmvTurOajrp2V34+Ei4kCPuxCyHHOKYCohw
rN6B/sk8havW+tgZVAMNRyWr5rrJio/l4Xz9+gey1mpRCv6xrznwwnVAQMUZHJNy
xXsF3IRojeVBAKPV2sudezLUdWu1fqEjOYakN9Qi7drKScI16VeUjsIpyTlzViKw
CJz51yi89SZhVe2Ig0cmI/UpjMpdqOs0PWBdADdfM5/Fb7enYFbP63qTItUGKU1j
to0xi48y8ew8ZxuCY5wdddddYHAR+VtZI6c5an9is7E8HXjogVwrQpg9CzhteyDE
T8NMQMjJJN14LnA92DCEOEBRvxGXdIAo3AnNvDA3V3GX/JM26yMn3VFA1pxrbOEu
aa2nxihSd28nxdO/zmoXjnApneEX8xqNK1gMsgMS9j1vXMuCmFTIWRlZYm/V19K+
VFM5iNJQKhQdZAom4860cEhox+b7ufwTuOCu76/buE1x0eaYgwE+zcUb5+e9MMIx
XN/xWisi9aZ7SDqczlXSvg+clYlUPqL6qFmWuxPMOFWan5ulHd4gh5WcCTkXv49H
tcp3r5z11pceZ1vl32ssmJXxur3gniXacjRa/DY4WQ3T8upNi/ZfHU+PN7sYP40P
WhbTwV13jG2yvij3XgjLV4273FTJW5O/lYb2Lx3WeGW5Ap3bZZJQdcXJVrRRdOk9
s3cyWa8sJPgNbB4dDOv6MWod0fskGVnVn9OWG70uaw/qbZbixX/RgkzaTzQvrieu
ahaz98LPHiwjRCJNJHapQTjCchHlyTp0tfx2ptlDV3oI05LeMTyVTrykPlIbP1/s
QxqbslV8A6M4wbPhZ0q/+W9pkzrAyKVayA0zaLny3YaQwH0LRvgm2R9uWR3voIAt
IHOq3KT5hE2bwuGOVaRIzfDN6/lEwEAydGQky44ViWkdX/xvvGGgFt+aADb2vYh4
Po8xQJnUCTRnuRJ2hPruThba5aFMRQjOm5e0bI4DeYCEyjKfdcg6XInGayiQmX/V
xNHeTIR+/oj+NcOf2l6maIba9dTZ0F+ddNaXri2lUMO2NT8pEZ4i0TDHKUBx26AG
HUS81ygfdZJEK0X9MzLk2IFvUP0F5LTc3wf90WSudEXCSiC1253m6U3X4YAzQxzZ
Xcyldle0AVDb8dQCAb1pvsohPC9TxPyl1n3XPUgnfFthGGOV+V8B+Z4DxIxUirMT
8rUPATYgbdCkn6vx0FVwkQL0ssVDrLfMdgkIMPFw27ZiZ7zLq0pbHjFWnqtQCe5H
69V79WWcBD94Whv4LzpU+fGX3JWYFRHCXv6bRLAR+flTha/7PYippkj7jc9K0M6o
gWP5x2pP4PEhmhqxlXCMqIskek8fsvFI737vvEEcM3Hrt14by1htUz/xODSNbLF7
623+ad8jYXLcp+3yuJtSDzPJblAuRqkiuA/F+hv5SFDOugI7RprSHyyr/QloeKll
GS2CL7R55rGk3M6dn+qu65uh7ORUo4SxglMdIDtGCmPem0fQ/yWz+HTPg1/i2ibE
4vBQCgli9bMNt07nSLGcvp0y38mhTC82d/OIR1+jQMdGunDpWJeLRj1bpI/GWeAi
zK7lH6J1mTLMyKpSJL9d5MJM2z+2pE3NlkYWZUb5/XGqSDSxj9xvLHv+2rSHyx4n
BkEwmcdIJpdglsfIog27p6JlLQYzOFmrWMrHj8OWgrwqvehicDpaKPqwHL34pUhM
mYQSPygjiqzJniz89m7q7w4IO+3gwR2QVTZGV1M45p83IhM2fo2ZDLlK4ULQSqx8
kBqs7mDXn99C4WlM4mdQ4UcAz8rBU11s4TPqzSypHQMHyRDJT2PF4LoNejaUn4iD
jIcuZ5LBh58wvlls6URdCm3M9SWHZv7SRaw5ayAFaHf+tv6TOOO2QvWSmfnjBZ9p
c35QM09J947L8cH3YiyUnXV0FPwZUSxEWXNxNr4kao3giMZDyw6QpJltWe3t7v3J
aSEDmyCWavt3t5n3YpmKY/h1d29v+LFdOr6Dhktsb1tx56t1fFlwQqSh4/oDOZw2
JwHbQY+lVlj/RBZC85Wx91REHc7zTwLl9IDRVOlfp4muVM3i0BYzwP84foKFYiUk
nui5WKLkEI2IW82PoSqghXWRtd2rsil+LcagpSr3mY2qB6KaswjcBRfdVVwzwE1f
P5+U2OQntlYfnqCGrPQudOstXrkArNC8avB3srqY6RtBvGa3QOSUlqp38Hv5K8sa
PhD8LWiB5rc3OVcRVFOfSf19+EMl5ldn6vcEGDq8C1yXb5Xi7fs/3iHXgtd3uxNv
8NS7aMev+Ini7BHS1ekaaXdpMg4HV2r+RD2G4pcf3aiWAIylrCEgoObPDYBOtzT1
DGjj/yBIXTOomxfgrH8DW2zbE+GcusJeDjbAze/fIaJQtOsXcmy/J2oz9KVFkmNT
aYkXpuFAJe+YGWUfv64r+bKhxdEGbKcaAeJ/oNoSVqR/nf24Urvu3yDQbDDZ7sYr
GU0NyjA7pcH6dq7DSyhczxgfwjxjDmG3jHZPll6b2OliSpr4xZD+KnQjNG9YUpfv
azner1teXnPYP3X7FNm2ZBIIR/g0bXDwOmBXa2KlCLjTsH75bpP93IS0JbSzz4Xc
R5Mw+4wFIxy1zDh9lCxbx32q61kn2TvprQ6+3RtqRUXHrw4H8HsTSxqIB3UQOI2r
qf7VraCIo9JYjnwnoWW/m1M9xeeUMb3G575jiQ0/x/EQAZAaZlqseuR6HFOStHl+
bovQJzgQfQZKS7QZaEEKy6BdMVpBnh4E+JpTNj3X1HqwbA1bmrIYtBOd1iAe8gLg
RYFxljWFvtH2R2c12dKmezfOJ6j1CRn8zY9iWXBM1c64Il3Txa6RJopp5S/thur9
sfDBVFhCoyE/1pMJxDeYJg+TgmC9RT7GaaVIhXAwTlTDNz0Q4zYIRvVyDa/spRvK
9x6YhbEUFy3Hfmn4gcCiCWl4aslFBFtWF6Z6XnPMgakEvjWPPCXvSgxUn0hhhPAW
T/YTj/by9XMyMI7QEGUJII39v9isNn1j3veU/kVyAkqWbYJsViL9bkLE3ANOFJpU
Op+Alc2SBy4FXVFBtM5pRD2zGg6MFbsODnUSYiTknPl9gSuF8vpH0nxYo8lEsod8
1hS+hFbEtLkcle6R9N+xLxZTNpGkw8zlUcSNw2hfW7u1s+VJdNjgJLkacqNxVv6X
5QeafghOOXK98JiUKty0SwvGEbik7sk4GphK4a9l8BNf+mNwWvMxm6mTA98bsDr5
pOnBXILnldK2cPttjC06n5uDH5Ef/78BzsOET3+REPZHLgdn2BnLmQM2ilR+hq83
ShYx10nx1He2nin/ceUK8ImEAW6aWmBLKhplTthv+7ENJo+gwrrDzvyqpTBImJHJ
5lfYq0picH+UTSZ9NO95u3380kgc/hC8bz0C8qNhuGHLY+cbUq2R91fYmv09APuz
WTApY1IQeUyI21YZyE9x6jijrY5977zfwEku5FPHlhm/zJ5UWnuQxwr1jYgi0+QP
zWdvfRUh9TDcrPdKArJrKJ5+VxLo7yy3XrUh6tcC26W6btx7OwDKW5rRhOv8iRZV
MOfXmJuaANxmiWudpEFuRaWFLgfZZv6CAZVVrM7G/M11mnA/dhIVoWNKgZxdABud
6N8ngUsqfCEmOB54spbQx4fYS3/55ygaCRS6tmtxjfpv4pZzPp9nzGkGvFNCK6e8
HEce+VeotoBWYcnrZtQmSnXZAi7LvMovXljujpzlOmXTt+gd33Ep08iFZ3GGCdJ/
rLkujjLmtBTN018cIyas+LcHrkTQw4X81FpbAwbYluTuTaki7W956+2oBbZ94+7J
UpsEDGbpr/s4XDwaZ2IEbbWo5zVI9JQZZ6kzllgiiZSWLioJr2cUm4lhOsoN4iwt
jnvNalIKQtZHEAmCtOCPFfs1d+bHhCmtulq+HMnjrM+3Sv+J/qcbyECuDBNHUPfZ
UHxyjTlLnAab6RBAaBpt4tnHD5bMn9LvPEDRO/HrGxiQk61j99buyJ5kuGFfnbez
fJrqPRUh6+lqpSoH8YcJE5BoEsU4EFP5cfAwlMXBG0YgldAN+IGAu+XIe/5D9GOx
n8y74uW5uY1yh7x9ZxN6lAj/cLvcZoYy6ndX32mA78vK4C5xOy0n1UN8+RrrhhWM
fbiH4/Fxr6qKax7cix4kYurKEhgXkc5cSS/XWedp6I4a2b3Mvud1ciW9FzqWTR0p
Ob55Wuku9WmXMnsGvz59c1GhRcWRnsODw05fGctSFAfCO8Oj475QMYIUNa7z/o/i
MNegTuDsMiP9fpYSvob9JCLCOpEAnidNWzVH5B8XiJZ0FGrvJHZwx9pOxV2xBRNK
FNEp6BMvSuivZNC7wl9dtcvH+Ee2TAyT1vpXdUXj7N5+MypuXcsU3i93FOpn9IHV
V7itg/NF34nX7pEJxeAJkkotJ0DsZqeDYFqMJp3M+JgrZr2tAb0GEkWYGKMdQJqL
tsWFszeGb3WHLcnta1hOCHS4Y6B1r7Un+ac77MnrZdwjG1raHSKzJaJFNUyP0Flc
9xUxNPB96tAGczi0gUzjBoyPd4N95FflvVkncP6CEXV6ZWmbY6zn4wsNJMqbQ59C
QFnNlCQocD76ofq2Q+y+Ge53sMyC1+tlqx0HXqPENinKJEtRUj/v4m+F+Zbh2sCO
a5v8JsXnKzUiZTimmKe6F52o3zqllc4WxlzuMpq91jqzA5M4Jhl33Y0IrYz/FiWR
ug9TLcau6LR4+yPdto03BK1PbA12YxI+3iFuSb2gBh2fMjiDvXh3byzFyB9Fsk1c
+c9owZs34X6dgskEbwOq5RCxyH21Gn1xewNUJuZ0CDPeqRQncYY/tXnS16tU2mSO
pgLPmJqObBUUeDhxeXCgTdXXIX/D5+yKELjEij3fSVix6ZupX1GCVwBxtYOs7ODv
x1/pF6Uo/rpaUMpkXpvOoFT1Kxr//9pzjqYnVhsWMFf1saSuvtvOA3oFkxj10Y8x
fmkeFo1PrqYkndx12z8kJXk8aV9vNM2jHNmwlLVI9U70RErBM1bffdb+E7ymsLeq
agCgfoTgEGcmdmWLvLEebgjWqdZBZwCOoD9/Df/oOg9bg7PXfQmozDIKcc6V6tZo
CJXEfX2ZogjLiSVxqXJaVSs0ItaecqN4t8SV+Or6VSmbAI3QxS/USkoYQtbAzQXF
7hxQEplu89wcvHy/OJK4ecrQvi0hIXST4fTYhPg9qXVOyUtDxHIG4M44sJF1JUAW
KB9+CbZKWZNCqltK3agzsVO/4CH5BH3xjedxJOM3DlfUZ0ZncNbcJV+KrlCPQbTN
PSmMyTRgkA5QJpVY5qHIhJ7AYOSu21RAPl5HhOF1kn7ux0PGIq08fDob7qcbMlUT
67RWe9y+KObvBIudOOdFjiqGfRUB7enyomVcJbHxN1DIIAJQAVbAtW8U32cD7Vvv
X3dBTE9yr02t8WuzLdw7fdnK1Gg2W339Zi75jaEeqrLnwhO43QqTiLAxqRgoS3KW
+nJluisRzeJTwHdSYIk9cce6QIF7tewLpr8SxOl0w8xhcvYhJYPkoUC49nQUnQuD
95aRIpJD0fGIBfXcNQf8+jmdGvsVyw0nZCwYiiOXzPCY4X8OpRpfPqHN0sCNCEYF
dw5AoUDY+hHelgPw63p3wq9e32nZgZDPnPIozot7pmjUED0tTTIlJ50V6XP8GwCL
OhG/L3d//+Ynmu2uiHc4taqQEy01bB7ajg9/+o1d7dG867Fnj3lfC7jSBCxltj5u
jjywkIZM+RuCYtMAComTaM7dmJPEVLTA2AA5j74Q47pVMJTE3n8C7nrxwXvzHX6O
GLxWbuSwEDFOhy4bEfA9JUTm6UyZj4bacgUWaOQHDnDM/GQFT3yqoSvIpwYmXDxM
QQZ9/v8MFtbInOI4Ml/lxVFITmGLKzdUD910uONXDY68pcwRk+Z2CIKPW9YvhFEk
q0VDCGmTVnggEKFS84Xk1gYkALwHH0mBtQpDs02Xf2uNFsUu0vU7hMHsy/ktW1kF
wAp5xugzoSUCC3LTeuuRXXrrUJNIvvBEGwO59Mc6uKynE0RxF93lFx+WDCyXWzqM
g5282fZtP9D68w7cOJpmzsCdMVWSqwjnYXPOyhaE6ljQvm0wNxj2lt7U4lE/6DIi
u2c17gHHfsKjpWVSOREnLUNZtc5uXA5aZZwR0sJR2DS5bYKi9bLYQAsY/mS6meRW
v7a4Tslz88TYoU4WKmlvNore4cF29CZ522lgfMD1DqNGkWdUD7w0Rd65abhj1mx5
1SEUxvrT6l0dbsyXGbLGNwK2v7ifsmVI6KZpGmXDNbTsExvuHKvc5muDxxuumhjw
E7Xla9lsloBsgUAJV8FtN1wdXHmRHOLdzKBhZnni0/1cGsbMlcJcGTnV50TvInw1
PFSKSCsKjLwUOnGsfYUXtm/W70yGwcD05A50N8+MbAddyx/D1Zy57kBMST7EANQq
BPzDqAEhaLd4cf8t047qdp8SJcb2Y0rJCinRP1+ntVonZO1lUiSDOC6vaHtm7Jrc
tjxvPKF4gs4DoptepVxyLpn6HylgazsXjKDG+7aHTo8ZIAM3J+PrUtUa/B47i6B2
YHsnM7eY1Nwn3sH7x7lY2DPWzu+UTJjgIGtEr05mk68TMbxgXHcFtBSh7YQ1mYBH
EtNWBVprGP/GvUJnoXud4WFQplIkQ5rYB+itu4vDFPjecoH1gXF/UiI5D93xo9JL
f/gOM0AzZACLdQBPPoa55fuYOaZCUTcK+grbc4uixfgoG+PGfcmDJmWH3WSvsJsD
5wWcLyKa7LZFMmiBIrOZuxKgcNtQ5AGWux5IDGKIReUkmiR8V5S0yDdXszDvQoT1
Odhsfwsw0mgCss8GBg1MYOABNJkT0lsSmukaWqT2mEBkQeelm2gLBHrLuC9a1wtO
ilwDW4SmSAxqAy9CoJ3fi9iTjxGISYJCsEGSsy0cnvY08KlcExV8YAhWoZmgeRVO
7V5BXoSLr72Dn/b0kMfG2HxRfTg/cuKL0pWfyQVtEBy3jDbhyibiWqLhuhYPP3mD
hMgCbIGSwb2MN4TOBsXJlC1cirU1uzrxJ8JhqnHZUzEgfZ4WDO5DbT3iLk7P1GUJ
Wzw2ZQ7jPIyBxJWuP5XnjJ70FtWTSw4L6YiZJ+avsK+CBv104vaMRfrrI2mQoWgk
e+hmN6+opdi5hcYNmjS4rHQJLZQHLrjFbFGO4ogqKFFrON5x9FqmnhSQtWRhkKly
cIOeKwAOD0eQ1VrUDoUjqPQXUE1DYblfXA9O3JtTZNigPHKMPMlu4B3AR4pG9qg+
OSZ6LZpyNYbLOy9mXocnoKnipz/CxpuYOYhw2b08U3hEJJM+boJEOiBMgtu0Vh8Z
7CU//fPEsyasVCujz8GI2q7dePMF7xNp+ShYln0fY2P/CsSKmvra4bmwWLKzmNYd
/XB52/zIhk/+4Mg55wrMhO4fbOea9g+SrLCfNoaoSqvIi6ayDvmuIy6QyS/J8niE
qYR6HVneIRjWz/gF25nO8IswuvDVPiwHFO70+Ka/okumZLZG5ZbMPWmHOPHc1O9l
uavA9Hwg5E6DQ5MZkIryiMyf20P3IvKMkxonqAcm10C3yLzKG8eGoTids1NRATBF
Bd5GWRVwyy+vA/H3HeNSmuffe7qU9ZzNJj+lusr+lFMc9eXnvLbH4g4RYnIxH9z9
vWeSK3SxrPOf4qDKnOMJZrTZB9V2dtE6tr9f7zywk0lDAvgzulXczEsi1sGerP61
ARCDx9R637pXUX6CU++r4Hjo56WjGUoOJlrYpq7VZYQYWuKgkGfwmtpaW3qklIfO
5pY4biJrSXUQj3ffoq7+H4WRriU80TT77zLWzLFawrVQzVz0eaMzbpBWGlLUXHoS
nVxw/KGOEn4CUa5bb5Ao2c9ZUM01bHAFZZQrPOqdXUTYAgJHhu6Bw79L0Z/9S8so
Rr0sho1EtX/B487HzdfgkI91lkK9GN8XlAQ6Jv/lup6AiA86kpYLeQW9p9s6PWoT
fxNa01AJAjRoQuIogLHGxOBWx1aQb+TBb6befRyZp6IufJ8sDosUMKJss16KK+Yw
cT3xOikwIzg+7q1oKaqCoeef10VKkBmOKFKdEZIDyVp/KSU024jQbl3UerHQKmY4
vRAz/CJZC7HqC+ceAvQ8PRZP4LVL4xQVbtCMESa7ynf1MfftcMB7Acpe3Hr4JFTz
NPSFKkPcCy/NH8Gbr6E0d+vxZvVPnwT639epw8inhBshe2TRbg+0Pvg5/PMWXYsO
3hbOWoMFTGfLc2Nsyfy6bI+CorgskGZwEpXAUZFfxGnunG8Q2+onCKUslxiW9QkM
M0y7SLwIy2Xrwtu+sf+YJQq2JSAt/j3wrRaB4zLNYStYdpm4/PoG3fpou/C0t4yK
gmxB9puMPn2Vdgy8AfdHozZMPUT4OMtEEld/agpMWS5cr3VBSWQ8y2mm0jHCp/41
Yt6DBWsH2HKwAV8UhkhBQPioYwzZzbzISOWdkz0XoCt4gOL25SABz86FDJR2glto
B5pZTEf9zAEVRm4gXsd+wDnHOsDTcgo4v3iu9yR/J6L1kqyha8NVyOMXEPEckcIJ
13JBeghbciy4ObSYmcR7Bkb+LTQapHo3FmUI96aN50i89nDDBasUWKpv4dl6a1RX
dL5Fv9Thox4oZSv4VQE2LtU7XrcaHXttbWCaEnZJR4J2yqRetJWgUfqWYOFklDVm
+PJ+KXmvei54/PnExnHLklljAvrey17WjrgjYA2sAnLbrQmo7hhZiEYQLuUQIoXb
4tNErhNJRWA3Mo+1cFYMgOnOSc8XeCpZ1joERyD0eT8b2paVxsrk+bR+4QXO9RRL
utJevp9b2yYZe0GYcIupDswpj7BL4ER4uZQ7h7jMI4xYv7xyB8xrfqo5txdOThHH
dLbVc4zLV3FNqZpUl9bEergDz4fn6qgtjBGhVtpx55UtZcTER9/xzbq+FaEkT4UF
cAq/0cDxazyEQOnZvc1CMGG2ld45+DjBFWYi0ofw2MBZUW9D35dBdXV/IMCHECbP
nVRScsIzoyXy8rj2PyfzfYqgJpu80D5/j+6Dq8Fku3y1BiA06HQWNlepwlY2tl18
6MvECprJZGKYUb3MDFiwKNAhZb5h2q3i0tei+AXXotGWW464REbI1sX8GomQd7ik
fUg/FmMeO50JgIBpygcQkHTGUCNbRIOUdK/GHG9damQoZXPabCK6NbnwQbuAAJfe
5ISChLyOGPtz57NVnPNdsJIfrDat4zntJIolvpdhL8dr/9JWIMQ2GM5D4LbZ/tOk
LpF4D23c/OuOCiYgUqHoJryR54d9tIp0xCeoC4LsRn6VX7rUozFm4HGk14WlFfD3
MpSZidG8YGkc2Ygk+2TwBilfn/eciCPth5k+dVg1AbjirjVTNXXU6KY91x1+p8PK
zPyEiIRA1FTW4Q/r4MoDbsf101ZF7Nb/VXQgX/olUNUM6cBsYJYh2qHWLFCOQuRA
huGXp2yAEEwK85LebK0Cgucy5+cHVxGepuvdt1IIGbBuYrcszFSNx37e3MYt5Nve
Pm1QIt7HddBq3QMaQm1CGUB0qEUXi7DGchFodrk6g8JuWiuu82r0k9CZNL64xGuu
KI1x1ZKrf2pJ6A248SAXcbw+wfPKUvaKgzwIGd/vLhKCeW+USCehAWuHqGRj+heo
nDztFy53jpu4je6KBAi4nQArhjn8D/fc00LUjiHuPXsjeAYaRLcCRlCx8d2jBd4T
iRaIuj4v2hOKrskABR/h1zFCabgGVM0gbqfTDRBP4THz9iNZTSkuGgLfDOcWSan1
2hDyj4+JNg5SDOqv+DaQjRDaTX2taoP1aa9NII0MaeLwmjYGa4tqN6AET1xwvCfR
r1orRwsipJeB7rkERrHxuJOp3f24LMykkA6MPNVLs2eQSrax7aa9iog6TuvR+707
ADeAdAc50uwlK2WUZQwuFtTqibkv6bdPGfVuT28J+Macjp2gXXtLUAGggE6dPEjl
lzg5GQ+L8+kkj31jXWJrCL/ikHnIQCQ7ooTJEbbDplr+7ZM941D2FgTKQuUmvdgh
7kWdRs54Z+UMjQO4dpt3T/yec7kXwB2ZJwU0ZaNRvB1odc6OG2+X75s2EyAZe5Bv
avFSUyhVSXgMgX5vh7s3t6SIctjs9UxpF2Rhvu0r+Mf8urMNRg3gcHFAdYwG0GZ9
WFbFnmd3AVTuu8omrPHQVi4cI502IFCxLKUOYruWnDLEf9Zi3Ug0jyES6Au6aJOM
W6imfg7uPifOgIvdNAohopQ1pBGkck/NETpCLcDmVaYdQsDghJKC9C9aSpWi6KHy
t5iSKHJ6TURoph8OO1wcK2JI/5CyV4I/s+2C4Pav5j3wO5duDy9WJ9zN6BADB9pU
Xk/sZbVTnuYOv+6MEe4DSEszQikF+p5wlyRA+/xLIHEo7jT0YMiUrFYGOyZDxqkO
QP1Di9dlcSCOmN6TjVdBgnkJw5l2krUIVyRFbv60fszqy775Wr6iPnAhXSbXNRXk
TZDryLTFSJBDaBe956AJ0O9LxIcDDOlckbMBWFPFhFoOB5qF6QI4VM3OBLdUZpXC
7LXAaGIFx4Oi866ItPwKlpSkhbVwZXb/VOjeyUTUnNSYYReQvIq4nG1Zfs6jQ0hD
1sTl6uyH3CYLV8+OPUAi0T8eex7nzIEQh1Mlw3JmOrm3GHBqBOuh7urc22OqZ9zp
EF8pBERQ1a2ICsL2UVg0aM8FYtrDw6rH/zft6k474cDdB9izDQC6lEqAV4O0+ij7
XgGbVWVfl4pJsEZJNCPQUrzEI363pfVvJ6hS4kJZnaEsZr4NqH2IrTbqa2YfuIFE
cw3rrS+GrWW1b7zHhxx8Yxkm/s57A7L1DhOwKUm7T24n0odHUmVUnoZ75CcR6nsm
0+N5w+ua4ZenwSbTIubl/fAHQ689cF6007q8DEvUnDDxIfAUqLCXlYi8LCDh0+Fi
w0P/Sh4aWDDSmEY4qNnOu8JAiCxIgkkBcyn/w+FxS4rFlxKJInz4ZwDG8BVxwpF8
ba9OuAP9otVw78s3mtpgfcoUooJQTp1H1zY5uwKcvxt8CvQ56OaVYkZZ8Y3D74gO
TUtOo+cawTwsZaaHf1OgIJwA/KG/OcDtAu7vo1HelNbyFkTdiuIotCvglnnbl4d6
Uv0KOg+fBw3Uxmc9NDQjStjeoQR/G1Y7jKgnf6VGJl4JwZ/LCwYzq3PhsjXzYtyc
z0Aj3Sy2sLgfUmLoQrLopWQr2yiejX4WFpo5hJ/HfIYq8wLRljHQZgUl78JuRDXd
VSsNKaH/CiaRAqBKG8+TXws+9YoSXXfPb7XeAczWY/nw2XRQ3VisQcjoddKVjfLL
nVIUb9DRa6BhDOJmG+5uVh6SiZUG+tEokhgp77gCmRqxFjO0iSc4Gtn3PWk8Iomg
IHPHN6UhPzK0nDZVT10pGrGCTUnKBWhlbMuqNWdzsw3n2kaFIeQ/v7A9ushLRsbl
Gt9bY0cpQUCdTXfmRXv+8KkDHp6Ho0ZhjqY+kAttIN0mQ+2LV5EG/SbHuAeHFY09
P8/xyp1FC+0iScd3wsLJbUr8UsfHSjVk1J99ToWT1kc4pLrRVM0ABbyhpA2bmGPB
P4rC87wwfMxxSl9uEuUNe4p1GX/0WDWKkyCpRos2e0GnSrefOxuyIjY5vBW61M7V
TUqBYeCjO5y08p83p6re1IHnQ5u67s+SdK2+guzCYseKteTwICv+2IXih3aZOmYj
45Kn+XRqlja7fsbJAo5SMRrkXBVx6IwNi2if/C5BN0ge0MWCfmBVwvDE11icKeN6
DUYJJ6FAHMmd61V+CuFM97SBZnn8AACRowb1Kd7p5qh0jZ187Yn5fO/V6pmwYkdp
EToN8aLxjBFJwp0XL3lNESciaAf3UqOiHupgOkFqjC0opMD99NA34GnFc5uiLw3N
6/A0OldO7eHcGu1iA/BUj/Ze+j8/c2iSXqiH+P0I5dUi3f+/5bd7PHIRC4MTWA8S
etVOZ+CJFr03bPzA9kMDVYz+eRdEYYHco7Y52hVNkwxb7NgKv0oC24ky4/N7Qw24
Qm7T+ymPw+77DoazXkGhyWXtclSYYZjSMuzo9MScaXNyzeCr8+CstVA4/F9RqlS8
yj73kQSafBkB/SyIau/0OSb/FtsierxjZlCzh68zdgkzz5tyKgFT/nXTdDyikmSq
8VLfQsTg5VStcG/2P6wzDR+yHiDYF5oGvWz+pH1YRU1uTg9YyfnBCPeDh05JIYfQ
wNtthsHV/vd8DtIamcYrOgd6XwrzRGq72qzXLiEm6m6tlLeQVp1LTOYxON6isTIi
/2cb3fe/Rs9GTrNV1B448saR5NZP1sSlN/8CUxtZJNufCicg1EVCCtrY7bSj9dIb
GNXTs/e2EdKAP97T+vW+Ks0EWX+/bVFxF/IDI+/64R3WSGzYFgomwCFmr+3MZ7KX
A2jcAVw/tT4IQ5eT6fzpR6yVtX4deB415jGeZyzkxGpEWyyn1P1x+r5OP6oP10/R
tQfAixqPgSaXyKjYRdzpcDInsqk7CBtgfLaXFUzzIpa5TxdqaWAU5UWgBMxPtGMV
YebVtkbZ9IFxeKAArDKhA94EgWP+PYIW9bbtZXRLLjGUYdQjo68OGDd0Ag5J2QyR
TPQuDzKK0C+KJ0/oZZY1CGUmTlXYRxEY68vdPTRoElZQd963oHRSA/qDm5ixnuvN
gIx2dEIaPLeCrJJvy+N72jkixRUD6mulL3Q7QHy42mT+pyFZ9aZWSWaZ/KgjP7QR
78kmhgR7pVtG4+lcx5/urCHr7N3+Rm7rtNxJKfbtlmLKJE1pibxnkXmWKfhQ2Tt7
jJjfMIOdjEadyaKSXcgAnyNTFQWEhs6wONnRFyvcJWmRrjOxS7Z5w4T0YmDMf7tu
+5BE83wrBlN6PzgHevLylx0DJe+yfQ/ZMkDVKYXki7rQ64RF5gnE2giEEp/ELiN5
2TJe8HbB731soXp9WMFlj8aTEeSBlXp2BYpMRMW8Sr5+8InR50W4tiUPeT7tVD5z
jdroK8cxuVzMFYRliegqJCSmYOaK4a+Sn6GoYULLfxRbkW8Nl62AbTMIz4sadk0e
/7v8K4kkJmN3gwNSlQEcFfPHDnHSKnofiNjIyF/TgPh2sIpxY7YQju4DKwnTfmy1
maRSL89JM4pGng2Z2Lnhxs28R2KkFpCZTSVk10lGI/GQ7yyi3Q98Cm8whWGuDt5x
Wb039pA2DSFZY0hVjwWjntcqdFTOySHS+R8+TPlBXk0xl881MXyxP3ixhcWEiyre
6ho7BmToOSBxPgMZU7gYtH26cJea/avxf1KuNt/YAfHdnv8l891N4JZb8mLQz1K1
SI2YHE60diA7U3Om3I9zhUq8pP2h1Y78rOA0AaHw6LDLxHdvl+IP868ZfqkNowKq
J55Mq8/qK/GZXUk1KDh4a2hlarFl1qklCsUqxm2ipzdh8XtY5aYp2pVz5ZmSR42v
faCOmuLuAyASx1oCex/cH7UrHrgIZdy9yd3pB67qJi7xYn07ca4UQk1mhwRt9Ew6
XMSGfvs7FMdyVdde/hik8/ObXp+wf6U3YpZbwtU6dFF6ICDjV7swpHGdgdjU2cgJ
y+JMZs4sXRA658aHEAhgY47zQgy/BnUrikHK1B+sOds3JKnb3wN2TLUtI0fvjX0z
yHRkdG5Ew+UzWJnPIZevocSsMHT4VlxOiIxFAYPGYnbUofCUKHogRtwRT2q26sbI
mNl+l+wwioz1FCYMImBeEzZ6XiRkhLx35DBNN1ssDqDQmZ7nlNCel4CL84JeFFQp
Ub5yW3ufNBf0XB7+IsBr6A/w/dHW0xXn9ngZsQe2njdsM6I/2S9sQXwmgOtEIZd2
B8VieR5dWzXyAjp1w/tmlrCqiurl0pQwa9BurkKEF6SSVvdygDX9xS1CoDTyRdmo
VKPAhrd0Xo/tYh6W3KJHQ62It912ZeQAQP2v2qCAFrbut2CIZpYh8zk9/WTh8gQT
aoOh6vQoEhB9lIog1+4PwOH/Q7goBE/+IFHYUNUru5eMgu6eZN5jXUmVh3Pfqp7j
CtEOvtsJ5CF4tc0DSX48+15CQhOqGeMJc9m9SqyDGEVSij3ec6zkO5OwVAp5WP4/
0W58kNelfpShW2ODd6ovU93GkqUCxXF6DjybFsyCl5BHrsXk4AvaSmFgWod1OG1u
+CO/+3fHdeIzmf3faN1jgaGqeOH4LDiH3gmTlzmIImjXPFnskpv936PZ0EJdqFaR
NhWl/H3nsxG7YYmc4F1iR5Lt8tugSDSg0VfoIdQFhxTsgUdUg6V8kUjVdc3ijda3
NJp+mxgaK2P82crje/rZFtD/bFHecymGIWxCfgICJkhgEBHbQbCxlDqmSFHp59Zo
LqnfYZt5k7ffS3CgTyFS5rDF/55kRhbWaSirzp/TOSU146MtHp5i9ZLsOR2yRU3B
q7yyr/qJ04hecucKXB2oqIWROIck5jks/EAJzqnOYVut1fA4IdfRsCC2EH/CjYgo
wEohH/QinJ5D8j7opBjyo6caOPcI38hv7MVaRNX4OWVqvdaxFK70xIKGjCOkhfVQ
GpHn/XstYS6j/iHG1Toc6G3N0ykOihEsOX6K3znFr4KenNL+Zh9FeGvkPnywh2Q2
xLmXJG5y5XThkeTS5qMKt5XISG5ClMR7NN6igM1MVd94UXL7l4CRANQO58I0ZJud
dA0oADQpz+txRp/PPXCY/VO1KTxlJhEUrlXBiXtsetrvx1AG2cxuIeBu8kqKxFP6
hyDfCdk+vtiYPRZR1HitdLSA5dHtrFFkS4Qd+nAUCEQVK3V/ZwCjwPCx+ulMGS+4
A1vRM6XEzIKA9sJouejd5Piir475PjzzRCWAUXNC1UGa5PU3fBKPv+yppWlU3RX0
RGT4l4MGQG9UhbSLIU0R0wvV66/KWloeLZn5E7r1DSMReElrrwbst7mwnqq43rly
OHZBpGNxvZE5UVKKmzcojZFLrFfxaHPvNoRQrb6dPRZa3czdcuxVo/7tLj7UUbNl
yC2T3un4mZw3pxnkSnGSQ2rxatD1NHIeJAQGGtU5YhDI1wp2bCJUVug9S8/08njN
rrt4xW4cZo2nRrp0zTvKWVmWMluQOv8q1OmfwqCyZeXBkIUiUJhzS6cSWaOISnmN
3TGWBhC8z9hzhPkGfTfaAlNSopVkSIADcUK0VvvrrXc2nrXKdjy2wDk6GjhRqIIS
1yx0snH0abGw69S+6V2d3Vi5DzHdGEy0TlmGmU/QOzFtya4AOcefKtCd5Gm+7hks
V+L10jHXW1mxqKl0DRHsQNPQdVe/R74q2rjN/dynBwcVwSzfMdHm1g7gJCjiJXLM
uCH4fgrSYCuWv8EKrk3jIDi93mcsZuiAQAPxiJG9f1rdmuzNYnrzGpi33oxBIHbl
PDPkxuLcZlzhFMtC2/o1b+LWgKoqwZX7DENYkUp351xal4dIcXmgyAqtefFZVcuG
GgPwE7/p4tG+nCMquPnVbBSqB+l/iksaxaPVtnNhnyz3Pj2iaYgTJod9PU7DKmWG
pUFAKGnwr5TPWxdiOyq8FRc0eCPqd2RzjS/N9R43KZXPyLi7fKEpAcFHWsk4HoLq
m8kRz6PbNQJK3KgmEpEgRm8l3MYcEA7AtNPeSshF9wcyqa2OTq7fiAv8wK8kGB7M
hIDnGK5H7+1+tXK56adzw07+Fw4rVaPQtWUeeUOHogrFd65mmYJWtFkpYQE2c7wF
NW+kCNCmBo0uyhZLGt9berGdV9L0w99kI41VfApr21w3/s4SaR4ImoSOm9fCjhyG
VT4gwhsXxjWUV/NOewmlQ+YM3rDOBj169tq7/bh6yzZPLUenFyXDiOv8HWEFl0He
TZRms7iZsew8gLzVSipN07+ZRoPZBA8ZeLbrYAdEbDv9cNUsSSYEXkrjNn1TNVJb
vz13860RdKnhVfPsjOAkkgu0Bb8yFbC3501uPTSSf8VlOTtLB2p010+6M2vkqOBs
hkj0WlMbeww73sVZ4EZ+Of8npjZfnDMdOZI/f76bQHGwZyz+5K7LyUjU835Nvlh4
ybBv7rmpFUewksFlN+Rfx7Pu8cRBJeiA/dC3fv4oUM5Dd4l8mBNYMmKTcetilThs
KDrwCl+DoaVtkI/B04X3XfaF5yMh0DMuq2RIbBzsiACOklIRwchLMLqoBlPpSdc4
9PdQeSS0GIasH+ZPQP8igMucDnk6DPrYuLIZTzwd+ke0daP/2kQf5CBKyKjKVLHL
5Apc0xCCBvK9CAthCeRvvSz++nKoSJWepSV2ws6F7IzPFNkOP0qldCbUycBRS95y
3jvWqJ0zkMd8N2WVm237DHREWmnLoap922ML/gZbXRQW7eN938Wvb2MU2RgKb5cD
PfrpfaXNkC/wEMmeElwlkD2zfIMhhqKRKf+hQbhDyjl5WtPpG2KrS5cHWqW1YBQ/
yoJFOHdXUt6264hZYeqtSyDRJnPI5hoTG5nPJoOL3+sNzl96pVADoTSyzNlKAAv4
lKOenweeKKmQ5lo0FjYKHgis2ZwrQlPoNwSH7AcYRHrxZ5G0z1AJNLGD/Qh6IbWK
sG5AvKsivwILZ8mbieN4c/UN3F/vGwRfPagnKoOvAffo1inpkKOvhQw3RUlBUGZX
aqLJYx5rF5m/jrSo22VO9A3JLfSDG5l7zXjJA4xo2xA2FAYgcrD38M+fFY5pY6WS
7uEwxYzDzldBSHJAJw3sSz7lAyx+DMVI6V7vP2yG/h0MkRzsrnHkvay9y2MJkww1
eJ5B5+6KI7r9E3OI4TjByiGjhUGWrSHo/f5zafngZceUMTim+pRaPgSwh0jhD8+9
8/rHcWdNn+YdVt4SaXIGaXacEV3z9FU4UB6sWZQQGbT4p+mGluu2ny/R3zUgr48o
2DXVzS0naiXU8XvBOfhEsKbh+8qite5qthhEuNF7LE35RKZObPnGHIzFTlJLMl4y
ZE2jtJ/vEn4zxNAaItkOIydkG71f67d6XUoMBazDDfu6nfECxgu9+JnuZGqI8KVO
smmsgabxkOHFb8NbIiudaHyCPZKELQy+5oKtZJ797X+Xrf//tYk2cIfWanZrvtuU
Oy9dlwh2C1Xn1ht1Dp6lIub4EqwRhLhX22PiGKn/ryCAAbs52cBsi5LxPplDtwJc
h9xfGl+Zi0ZMJL7e5YQ+i5GF5b5fbdo1OT56WZYfqzDyYbNQ8pvg775N0+zRkyU4
Js1CdMWeeegagztPMZm2e6BL4WB5aPCwXg6cqO1zMQKk5Hz3jXLuEBb63Z3ytcM6
wuyKS/SDQsbYWGHNyn7BF8CTv8JLv2hqPxoKuxuy1IIrRXGEdGXDyXPczi2rlzII
2iXsnh/gQ4Spw3ra84M9lc3ZWfLMiFIXMhW9SzZAnohuH1GIjgVaoGv4dAY8BUGv
9E0dRJJOIsf5OobUaJtkZArtwvxYb3Jm0527MU+G/zHT8AanEEksug+2iP6ijqwb
Ivj5nyAuhHdPQZuet9XXNVdDEAjphosk9yFcAEX1DtSEiNa9GKiAjVItzViJcqOP
sAmxoURJ5PJ+xSGZ3z9zaUjXOvK8eeUiJ1/klVyj9ej6lP/o84XCc0Ux2WNAMlVs
88g5Fasd5/pgiR/VgtfpwNQfuMGSV0Nu8/uq00bSfsHQTXoennT8jsdnA7yR6jvb
F9Yz8GW22YbTQCXRebIqwPnNm8xWvRoBwW4MjRPGUi6i26tafJztMyi0mnmxdE4q
djd8ELk8wYRcjJdO8vNKMMALnPsJX0vFTv/8s2Tby4eSKjdt/YNwMnWGyiEEbSOT
0Z4ZjCLvLnPVRUrL/iQ+/eBfiPUy4ppMVR69Hbv2djAC8wT914s7CBzaa5ZqJh4m
ffVDinul2GNKVb0W9zgWzuaWOUudcS9OrVGOfVP9VwyNCVnJJvJ9MEEyZ5NAGpwU
wHKQsPIinnzT1iHxP57a9gw+AKIXZNO2eRMJsEQ8GHRQdabRVJxm45PfPqRzUadx
Dk2ysMdIFE3o2+HZUpGAFxBXxYfEoRiBH33hY1iEHYt4pE9pNWHVU7zt3cHh8wL1
GpVq+XccaByE8G6Tv13aidtH33WBozz++ap+hSMlaUQ99r5p+A91ydWw4W90+T+L
sNn6pix+NWCJOBm/4gRSDPs2IuX8AIXHp66Bv/ihn0i7eagzkn1fLYqw9ouhRLQO
P9ANA7PQzKV2EHW+x7CkaTTdcJQJ4oUJ2TS2AP/PB9J30en/zLSxUmx76YNGqnY6
19KueVVEi/aH0VaDpue+CZsS7MSPC89riz6PE7bZNRHXKAOpixZ/BUmzuuLu4EEn
61BVvfETm376qWZWvyithU6dTFfLqNVlZ/57DQE8bwE5/X1iWT/CedCtxSms/OSy
BsDcarOSeA8rhrgsTQYg9AEYuqoKp6WivrkyGRoNYu/0PesruDxCyOCFTq1c+3ZR
RmjV0CqbyoWGpsDQ4vLawGd0WpOoflj8xDRhYGSeLaWF86CF3NcJ5aKrs628wEV3
rbXXCDN3P4XwC7AvZqpBqmpAnqFv81fTKI11VFbS5OVK3F6PU1FVILVGvq40MlOn
HOz7nfXBytwTkR419IEp464uF7SxJxDLXgeArpYGdBycXqikUtO97p0novKROhFj
iz8q5hyJL1+v43tEnX1wA/VT8mD5wbHYSuXASBmSVwTtwrVnetRvJO+f2Yha+rr3
mpAXLiLGPrtQAaiTzFt4BbiUjRYflijwnB/rXwsoc3/+1GfjuOBm2ON0eWtc7acW
gLHsoQBDEPZT3XMu6Uvktv8iNKqy1RRIKb3WEng2/JZTjygX7txyzATlEoPMA1wE
fFO5fJ7Ox7YAeX2awXf6tc9Oz4VVe/7N/cPUhjUtCWTruX+YZOBQf+R6c8alalUR
CguAg7R6outV7e5Q+YpJLqDi8/QyRJ66xTGoUlbfUJF3eA2c923DIyPwuzsI6/b2
8YO5/BDuGzFVwqJk6GxL42FWGwU38xKCwOPSQuBbYCgoIfZsaGmLVSNr0GZtbQS4
qVdfUoGimNupeqe0zaNfgA9RAPGiohdN2/kN2VAEDL/J5kz18AJGXD79Vp6furOU
0gh2yMeOCbgf/FmJf+jDlVISfzdNkN4jG8jksUZNcGWFSdZ3sitFwx/8LcRXDjph
9pN9g/dYmvg/bTJEMhFq/a+8rSUT7CJrh8TA55w8PGTeRHNG+2dokhixHGrM5QNM
bXOcnvEHUDVZ8eqaIZzU33cFPXohwyTYqUaK/ZYVBimg/Q4VaE7ubQL/Mr+0Mk/B
GYDbVM9w8vX8rTLrsEihMf7VuaGecGLowtsM3MDEdweksMdX1WniFwSIJddGs7ST
jCCoQ+HbmRcAkJQXYf9NDrJRvsZobhh0dMNxQT7uPc8bcpGRH0cFO3Zdbt9UM9bK
NvGRsX7ztXTcM9YVTnN7OzFg8uIgVA7kOXF+Y/6RYYACiFilvo5SLZCa0k/i3f0i
xLNqF6Hr/2DscOno7En9pzGe8JOxC03PqXV+cDk1xwmKpWPsGw8FAS5mQ0X67kIA
JRHgFeB64DM9LWJHK3I4bAWlJln3gYsq56xbikD9fW4uQ2MGhzRFZmcJNUEGYgVQ
Pd5kwgaaHVIIwMDfzXy6RvHlOelLJG8z/j+BXgu6lrI+1zouknV9dADO5nx0vzmc
EVh8JxhZn6+67gR60RqQV02l65KkCAy1yqHZ2jWUW57++WaiK2Pzn9W7HCm68oq4
mAR8BEEGmbrp2tnIGpFRCnfEM8MdgE2TCvy+eA2OF6L3vV7MZSZIzjUY08A8PRnw
JaJ9XQl9mH3ssAM1lXQwX1PxKCNA93kFZNSxcnCR09Mtf1NOanukBZJCSXoTKiAK
sW7BGncLI++4BBPEo1HsiPLFtZ8E3llQuO6EGm0IGj9InOpO+EdECVWH6euvm+Va
w8pPEDAVdNL10HEpyZSpra335Yk2pbZMkcK4/RaKane0gL0nlEvYnSsW57REdV2b
XtehSTKUDKKNz6bjss8txmtfUMScJhD1AuFrN8fTKZQ/7lKoqBEm9/AtS2LApVOi
zqfs/MxbWx55M4pFg+zHpgmFcs4yw6wO+/5Dl53Qitam5K9lBYaQUQHGuKv8UyMe
myW2DUZaQlQsH43X8leHeGjV6OG/mAc5D5zbt4DbR675ufziMsIlGD4N2y6pZPRI
sp88ToThk1voJPNf4FPGyfHW/4fcvwWs4RV1wCaToSj3lKwq3vgZhCaK9pwxWd1m
JTcOBk4EZRo/1xFRGDOn0R7VEIuN3SvPQ3pjCKtpoR/tPYkveMaQ67oojYThkHv9
ztKBVjUAzmAJxtqWCBbQz0QaDWWLlESBm1STjGvohBTCQRUCK+E4odkb/Y7NkpE4
ErT9UYmQws1f1GIuW3SlzqzNOQaTPDcZFDvLVZBT45+zAPZeEw83Ur3//ASFTftV
uN12xepyr3prrdYzAAiF5lRjJjNeFvKXweN6i1bVqZ7dsAZqimcTb7//6ynao4uD
m51Th+uiLz7QladvahkagDlrctSb+1/2Wxijb0xUNBTfILQbGKP0YpMDd1sx9+AK
YZdJuZ8WjnbSe1cPOs4O5JjNA3iLAxYOpQJ3ivWOrR3I3PuUygT/BW/OiOL+A1UU
RA3nUOz/aDr+4ztXZOtqyjJPZ+x+z6WmilwrAfwxGFo6KvKJ3bw+GhZsP1fhOvz4
CBUpASayvEjJIvVPktvDClkrh/aSyEIOas9dydTk1Xg6nfN2sh+QvySIuif3qw5N
mOEOgGwih4LEKaUcmhLzq+NKQS6UgA7SJ/4TCdfgtzAcWrfNJ1Gd7HhKADwdhnzg
3af47APS5CgA+G43DxmdZzmWK2vHcibwbqW3R/mbtcXkAmIUwTO9YDBI7lg9YW/w
64RyJla/DWyrJkWHjRQ2tnMJ4ir8lYIzBsocJ5F5PY4gffuKXD81qm2tWTNZGBV4
a2w4Pl0Q0dvGLO/CA7dDRvc0/cZGCknnfZf0lIFzbaew6q4K57KfMtF9JnvbfuTj
YClMsE85OHFtKAfmlaTT5ez10UXRAAyYDJaVo1t7JPcGxSWaGMbBXJwWf9vwXC43
mc/q5L29ilq2qwvQyRlIi+Xg17HgIIw6GaS3QfRSY10xW3aog6sKc3ZT3zxRgmzH
kfOvXoW1sf5HZAe/yZa2eefTXzY1Y1hsXgSxh58D5OKD7irfAoRLDFXTVUj+3BzX
Vsdp/b8RuVrMiZK4s6nUMHLH+vfLXw51siKKBzTUqAGny5dDwvXH+IUahGrk1ayM
pUScAPleVwZ0KfGyEW0tH+L6txrcL1l4CBWAtxTOklJHHFJ0bZcaDkkPEYs6OuZp
bgqz7npv8dh0NQCQEUo7QdfRx9GXgAV+0qnT6tcRJn9nU03BbLCm0cR2cQe/48D5
xkVCMRjWIssQzsZ0rvZb9ZZEpK3PcBFEpJxVyBBe3c4CpSof1rUeUka3xJeIQeDG
KGNSnNpVltJ43e1KfQF8Q6Iah3AMgugUGwmPOuKVBKTWY4YldrOe8J2ltYPqqzzq
v4LivTISy1s+V/yWu3jFLqWTwG10U9hEsBATnSKc2SyzdGYVUxv1c1GK9ALYxZWB
kmioew6y3BP5WYvxBdJEw0Mdk2YPfTtPo7aewQYb0/A1dL4lwRGNXY+F9Wj65Vs9
VuDhejsnvBTq6RfQ2IqtpkUi5nTUVTqscScuc+2xAD3kgGMF1JRYsep4bl8ybB+J
EQEp2OYPeru781gfMHtW8WbbsG8/NNXqF1JZ8woWvIeDY164YM3q/MISrgbs6b/g
UYeRGKXrB/f9c/vP+gi40ORmjNutU2etrEVOSWAV13/hlDXeoLM6opDuypDF2Zkr
RT7E1Bx6P+IF/dRzP5BFNqITbd04mPmRgiUdfKDABlPt7X1dI8lEkGJOOq2yJ/m0
Xqm+zeV8IJaeWD8BdruZ2Zkxg8yJfaVD3C1kbaiV9LbUmGr/NRF/u6jKO37DNG4L
dNwipPgd/WtmTxX4Sr5If1fJFFfn57BHYa1bWwTtCPIj/ZLT2IqWKgodoA4pYTZJ
7RLpAczUaNfgXAguyA5ZzE4hO0ZSkt6C2RjhXJ8+SUSqyPdvvMVsvGuz+Qo2cd1H
fPn6xIQlwHgH6GiB4qrx5PSxK5df8aIpBwm+VW0jS+d9L07+oaMgVZqOobknTKch
nE39k0r9pfX5y8yGFIvmRS0ueegSXRohfusD1N5T9mrKk7RhoAXsIrUP1h1ycqUP
usHgsULIV+MSluAlZtn4ynDe0ED0cD9kr2htNF02s+YWxVtt3aweJamSeL9RdbIu
6EK+t/ftkUPlqDxY7Uy9UyW1H5+cAPm+aSZ2FvYBGqnjpGd29KsHqeQ4KxOn4nGU
ucuJuFRpWYvnrcLmra1SmjHpQgJqeBpa1tKCtPaTjHzJuT7XYov41+bOt3MgHZmk
YYw5m1ipSwn+eEi5tOe/GlFuJxbyCJ/eDJmI83B6uZSPurZKfx01RHlA3TYHg9Xq
VA33MIbJQM9ndaZNuOiPR4DSI1bCqhMml/Qc27Uqy3GeUDV+HhAW7CrUVb0jSTqs
dCdutMnwDG1VVBJL8nfXlsIgcZ0hpuHuJIJqdjlVcnRTRaOnxHJfRhAiZcfkja+Q
CgGASv3VQm9vsrLegnGq56hf7N8/pKQSIWeathtRwrdlXYhz26UrFPrA9Dw0Ls7p
CEsfLny4VddPDmsAV3dWdN4cA9oUv0lcEa/KZ3ADYnR7GOiD3KyZ9McFbF88hJ4A
qVVhYtQVwNb6oHJ9+O1jLvNTIcrezReONCc1cfzh9W/fGv151TnV8/dpIvtiYoRZ
8WC4me1eczXTUQPKHj6paoNZtNvh02kl2bTCzbPNLhFsU4qehMPgmUg5y/OuRPAG
DkxrxAyPBiLMQVJ2fID+GAWc40cZdblMme3CIaQjJ5bDzllUFwSe9ueNFon2ERsR
2fymNP1jrIZy1T0jOSO1j2NOcHc1WYPRX5Qs2X55YPrlTGmqYBsmpWwY1OswBo6/
CPqHEF1CDQs9yaIt7ymNrvVmpIr3vdnvWLHy5yMUSyUkJDSjh+/5Aj+VXZ4c87bA
LNpfRMNaZxbdCDuy2FR25ipvsukVZYhSEEaVoHyhlfzE4t33CdY5GMHM8AuyeqEE
Rs1IEhINPRnk5RChjvw8IVvWY0ej+WzfXJteaLMIGV72ipywJZaHxI2oE9nlnWMV
MTqUQgo0+UfS0LsW2FNTsYakrpTQtyiQ0acZ2t9h2trogT2zb3L2OCKQ8bmMLX2T
AxWnD8f9HvMKb0kty3CpPJZU6wF1GqXwsJgvqDptu+jWv8fXz2UF+PCcSJUiF10a
LuG+vO1dJrFYvWSTMFwJ3odJMRy/lYv7Kreg7t4X9ua4CMQpcxSe00AyywFE26t7
DD+Jw+C5sDqhGu228pIf6q63FkvrPWsxq+ZO/a2YpVM0wotJoUvbHeq7vkPwq4TK
e5Dwu8U9R+zcZAUf3T1l+GThXqTxk1qC7jkZKNhp37TYZ2zTWtuI8shvmpu27DJm
ZyQc5HPVy88OH4scs/2rL+un9jsZjwMus/LRSKBzCBQ8RAQxztG1XRejWsn9Sbr2
7f5To1ywOl5eQmgkslBFGvN+Lyng0V8rz4vB1mqFIhVm423GLEYzgtLKfssMTBuz
aYwGMmWW4qrVv44CwxX3ak9Q8VMOqXDkSf60mOnqWzc2JA+kr/7zCykBkNuxpIdG
+ujddtjNdBQl7Tnxz8anwZd63YH9/G8aARyB+W8QmTW3eW3GzOKSXonHIKgyqNdp
eh4HJV7qsmW44oA0oPiSTooyC/HIP5zufn6/jcTXpc5et55TOahbwyh6xqfqUlVX
ssUJNXxnc+qjBnN5uG/ZNe1o4iiGrzCwBE9Cj8ixE2mMQXhd85QFeXKYOW4PJl0I
jXf1e0p3n6ndl8mJWHrANcdz9kpyfGTG7/M1n44ZQUknoNwsOszn/uoHQ8au6SHP
Ia53DNavbf5BgI9YTbAmAbY+RlW3JxuHzp6F6bwiECy/FOc2Ol3h66URrae1Q6eE
jSQgZPViGDs5ffHeAe4akiis7RdME5evlxgrh9cS5FHbqJC9shR6QENtZmikF3Ic
Dp0RhDeLIeIrf47xpyWuyETefdrdRs8NFIU3OxSndBcg4Bxx9kvRpmy3jNpUDsNK
pa6gotwUqvrlItbbsgOwSgzqA8yeSfmZixPb2RnUXD1zYMHuguQvgRRErE2BJdu8
e5wfW9UIu9UfJAjTLFaOxSxAk1bVItXtDl/1QlTxIk56dJHwILZZbKVr9mIKN7ES
QYN9BhHMWJgrE6a2RJMvgSeihbjmXOgjsAUDbQIQAbMg4TuAQEDo5MOUjmiECPsE
W1R8wT5Fd0bL9x3BZVQVRHaaXH0+2N45idBJbEg24ZHsGhWCiXJ2n+0rjgBAsayL
NbSzNLj69L/t95F//x5K+BrcjOPLuBeSm2tI0XXt/bvyFlPVG3V4XBhn7vx+PsOs
XZWvUEDFA/jG0rCZcKTYFJ52++N4vipj4ZAude7fEqZ9RLKHqwS3ZMUByEZpBE8C
/4Dxre1xipZkuj+4MVgtQK36lZfiw3zOcL4ujjZwFnCzwae0Wg9mZywYplRGVoJR
veerybOYdcpWASYk1ry3adUuVJtN4v21Gwq1DEs4/USyVOSs3IOIUyvQjjxNmBob
gY9o9VlghMXEJL5sU/7ktc1NtjwIIZPCB8jmsa1nYqJGck4XP96wSTFjRcH/f50W
PafYK5NtwiBqDxQQutFyDG9+ITNOY6EfxIo9vtnIPMGLWRq5WlJxqDb9bp1ld+Vg
WuCOno+z1fqCtIYctIrrFQkFejM/PPvUV66o+udMBt42AgtNL/eVwAq1vWhhPQ7s
NKjc5rNGgjWn4ELoD6V3/QqQdGpqgDyL3r1ntgbRAcJ976eVd7f733Bw9U8mA5pN
iOViTuxfLr8nch40TuB8jKDQNIMAT01bweyPXrWpo1tw31J//0oud61EbhlXXIld
B8fr6ZAhv5sv4FCy+n2foT5ee9ai0p1A4kwMXVAqUUcBcXdmjv3bjhXDx6eEKEX+
Nk6YVkZOqkyNcvluV4JrDXxR3pb5yL2ZomRmM3cuUsHhrMNf50LtaUhcDLYPcfoI
x1MSD8tzNIRCn1l+elS5SXUcxwXLwFXUY801dMrtTQk8zN+XG8hxt5/s6jlZv9g2
7ZmHnM1ebG6izH+gHSQjA4FVaxoYvugv61y8fhAnSBuz+inlOsIKFXlWMnNyQuJ1
02vNHyNyMcgs63LkNX8UA5I+vwdHN3187DHxy2ul8DksBIwXmg/CIE4NnsD9qw88
ysa2mTWHkYJN3Itl3fW6BtDApJH7kZp/61KpIPww8VJLIrH6w1OlURmYzVEqnZRF
ZqddFVrqEjzjK4U+YaDSyrLCRJPw6S+yvHmkk40RV9fscH3+JOSq9dtQzRToUPQW
JEXB1+Ly++R0bLhKGBY7mvOaXAGtJ3Vp/VRThNBiWPH9W0C2RK/+zByES044ByIw
ML0BGi9UZF4+KwkhhZejnYvUbOC1N2BgJkrIjyDbal/bFx6QRDim17WwYRAlVMIm
YHU2Nb/3U3NGGeriu12xaSJ9MXgVhviDosRC3aN9pOm+OQGjb05GoK10+DHo6Efw
bzrYAKIC/Sq67+JZ2ILdOsaunhTglu+BI8yYQLRTdEsprExyywog9qQKQ8emhWSM
98ia/7kcX9iQ2cj8KuacvmfAxG7lZoTlE2UmQp/5+Fy0brngfZz5EugV7d7esGwK
LW9YkVbps6RUOFnzoUP2Pu0/CkJwAlWENpdakQlVdxdsx2sKHE3qPneFLZBe0Qcq
2rH9VtvdVQrOHQMG7Ce7ujz/1UqqQjz6ky+WCUZ4g/TRyKHps6kIlwriALGx4QdR
9xSSd4oYmuSB68UhNoMVzMrEcSHk44hq1v7cMYSVWZ5kkvJc8CQj5fH5OaL7yNgE
4i18BWB0F79ErDG8T0HkTn6+lbTpZ0MiMWWuKwH2AQQJ3lViH9tgL+6iZnD4RSGh
Sz0Ub34UHFcsEnPaR3sY/07uMrnJKRTRCJvd1vhqaePd0vEQOLPWnyf6jrmnhP5t
Xm4wlZ53e0WuO4ZInAUfCR/eOBVGB6CRbzt4seSlhbsRgBd700nVaF+e5yZOV4cT
uGPkQR29P3+9jci5xoSR+mp/nFiyAcFRQsvgam+wygTUCpaNzysdIfEWu6oyXya+
LMC3Yz86TS7ab0u3bJ1q00FiI6URJUpkq+5+61F0tSkFEkSXX8nHV+ceo4JJMlTY
UuHxz5R1u/ybT4hjR0QEmYU/xsSkV1XzABspjNBU1JXdp1KXv53f9BVFFn03IVk4
Vfiyam5U+TDzLCwBBj/8fJccVF3PTDWraUugrzUhgwR1Z1bBc6OneYnTXUK2Hq4f
Q8maGW7X3cGZ2TOD0r9imqG3iH2L653zyLVF8zyT/o1Otkwkb36m6i3HwB+qDkGd
l42Rppa+h7sDfsWfff45nxN22FrcfEsB+gJyR7h+c560l7/nuKyFQ3wf2MU3vH3f
82/UM2gdllVpQ4qE7ZciRu/h5uDvNDyfqDBFxDK0druLl+dwTnPi20Btn+hLizXJ
7RZd5vHhCqYhaAky7wycwE/wpfQfmvnP7CpBWUpeKf/FpKeRcHiwgaZWPcVdPbhR
yKGhT36s9yBNyIaEZwh3S2tSso39F/VofI73Vg0zCIIDQ4cm+xSDIypG53Z7BWq0
6BWm/hlRSW+XcrrOdFJkERpoXmORMW9tVniEEcEYfj/FMea0rMoKRNRD1GtjEMC/
oaxoZkdRjd3fnhOQr6IHKcz3g2+VRntb1Cval45q7Zg8cETok2mWPN5RgvtWBmnS
t4pkqhI1IWJqzZKNcUjVrjnIywWemqnqerh0sogSLCX5whs9qkZ8YrQAUSllDPr1
q+UHI1pTl1Zj5M6mRGsxz+AftsHjfzMbSJNcigVTPGYjPGQuKgl/WNkzdhIfrdxy
QKeDo8iXT4epBZCfN87F9C1ia14UkfDCOV30OnIU/wjSYWuCMqcM8zzCBsXXAVpF
jCSbqMH8WstoI1hq7XD4dhSESjJZhc4vocpblrFyhG9pMvqOAO5Z10F+q/ZhqYyO
fYCtU6pvwU/dDgWu4N/z/WahlBqo3Q94K2We1U8hlkq3utc4Curvkh9LX6Gu9nFn
GRLOlcxJPoG+/ItdABSkMsoULMkvm/bZcoYZ3db33Qcng2cf03A6vGELL9HqxBXi
vMJPr2O3uvY7V8lL3BuibTz67RTnUyj7oH4w4BVPhQ5rhgAOl0Uyw7fRZvs4YCNE
whC7SMEnWdATemChi3TfPwzxZyQ1KoSgU6eXvKoJSonC4JmSJQS7LIYNwgVAcxAt
9CP5oFv+3e/GPgIhgzSzDpFy+Frr2XJy26anEodbXfNuAIye0fsJbBpoxigAPKHM
xUUBUmz5+arEj8lFl0uRYqT/Pnr9wgwL5E1Ix/9FtHE+kPiFJdNdvIojhQdLOZx9
/4f4aaKPgcAO3H4AwAGVLhPQf4yUD9wlK6TYaJUb5Cq1z+OB7qrMYdrfajkrD8GE
ao1MxI9GebNiFpGinPX2BA40E280CT7YeBL4cMNwVKxgRKnCvCLmZrLK/JXhoMO8
ohEP8VopJJxh+uKo/GiO5qCKpxN6MrubN2BDgCySzGNr7mB/0BFz+OkIJ7YghweV
3bIbGbzt2r9Jfzei7sVHUhWB7lvU0KJnUjLEcn7PnDy2Wh9oBSZ266MeVnljYxv3
0BeTHpJFXe5CzvhT1iJO9bYyTPbfW3bpnXEbvymcBRsZQyEyunqJqPz3Nn2XqZlK
A3gBaNwOsRcpGROTHj/p4dBgoEyKr6lS0lJjtmCBXur/wN2L0H/jt6P1zZw8cFHx
iEIENUaB453fBPs+wMqLT5kZ8Q9Pk1EJgLam8JHajrozCg78RiwJguE70rPgU+4I
MKy3yz/CJX4f52CjIPaQgGHtmAZXYWt4KP4pkESd0sK83QHxgdpTPK8IHhNI4uiU
Qwqi148nt4qL3PRhLpzWU3KwZ0ii0a7jLMIr/Vk/2w8nGgdd9JBCnbRRsHmf7cs5
ylgxY/9TRNIvMDt5ap/Zf80R1n/AWO1n5fzxy50GsliCIftekNHwnQa+Bek0Mf6E
btH4X0VZam2iiJJ4gkZ0mi4E2Lo/VgoU9PaAJkN0TG9Z0SwbzsUO4CWAnuY1laMr
7AgL6iM0XdcICzFk+39pKYVb98Ln4mN0VfqbOSgp+zFYMsR7NnNqFnwY5HkQzJHH
AzIGVArEoTolXzRP0OvxtueUGKnj/XSH3TOXutkhL/vKguhH1zuIG5GVIXLOfaq9
rgYycsYRpHOQzLDs5pNhAneLvD5nAtni4Foc6qmGqKzZfXl9bJJwhV2iu2LiMDC+
y7OCv1oWY22Lu0HbcyQuvRmGahrxmu4TlWxcgeDtsMnoD+Wsy8MSAyjdgy1/3KsA
6mxLQLFRHXLiuG/6kOCo0ietVg0BKd7KbgwcOmo2S6U87aqOv3jWcx2k3ZjKazGI
kdNH/0Awi9NoE7NLPit4Yk/l3/4RWDOyYvpacBLsxV2bY+ceieRem+0KoysysTIz
HfvCyHpHCg4e9i+bbKh1RdcFJw9KH2ShXcH4YNTHIY+AHQIXgS/4QqoUEq8DfJp4
M+Udn4S77lvEjrhmo19byOIzF6ervdF/0Jmc8wey85KGUd0OpKRAr2CA5aDiFFwB
7UMHkXNIjRsnov/uJBy+YNiD0J88q26h2xIFBJp5p2yIZuLq1MPE+7XvfXPi3dhn
8dnq038SZSx658JXaI/6IFZNfXWO5LByv15w+ZvgTjM39lPs0XLPcUQbcybeSSNR
5x/AoHoI1Mt1fGb3mmmRnbaE9Uio5nXnxWbsuUxwxyCJOP8ZFHx5P0oN111whE47
yMWAr2nBSEfcDQcBDVcgD/zsDBf3sCOh91VSpcSIxlIC7iRoSp+vUjzJhG3zZiO2
0p+pud44ewPEiR/1shzWenImrEln+j9sL3txtHycU4VKob3V16Eg/sG7BUQQCXxT
HE1yYLTD3GfK0JkwF6rSuevjlSNsc1GNUnYTAd+pqScDPkpZYGu15IZWNPKNYYyZ
3kCx0FpMOjo7hiEjcTrFVw0JrqqCqmN/nzfIrp4efAc/PhFRR+J6BJ0NxL8m9/tK
BikZVTCdWQBxKSa6DkFU1YoFSTOdzEj+P1kCx51TPGG65AE60Tx+xiE41gHRETF8
XhXWU7W6ySF4IxQelcahEzKj1ZxJomR7afQMqZZIHzDNHUBgZZ1+0e9w8DLq/H4V
lG1S+EebNPYRfKYhyY8ZvNbWG+PJfdSLxDARdIejuhyJ2bOGYl+3wKGvYGqMXs1z
YwKedAtL9jQy9MUKI76XhzQjpRuJFn5UCT9FmH8VfMi9MiYz2GvCaFlQfqYxvWi6
Uq76GuNS4Wvr06FOGyxlmiYCd5E6xlk/FQFM4b4+hqFCkEuhpvfzty0fWnsxsdIx
`protect END_PROTECTED
