`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z4QgWb4vyisg8qzpeE+tvahFDa3lF2QJaZs32mxOmNK//vfjkV5otQX+4QI1cfL1
rlg0fBsd95xUp7hqlP9MP5rcpp7r1P0sgJvX1fB+VtdqZAbcMXb69P6RDq+yZax0
C8XX99aAkSLoAKhWt7x7VV5HZAJHUqJsbTHQbgRrE/xGdWtuuItn0SXSHzK1Yv1P
xUaXpxZYX3fTLUTjKEj+vdu+DIFSmdk6S/SiX0N+kUzC93YVD7rqzGDkRJbwtMFk
JTr2sg9btQZmah/fRbU8vJbRY5WHbpX1FhA+YRCoyYDIkMwVo0ZNmgpFDmF2jLai
a3y2jZ9Buz6uldDtI/8JFWCgSSHxzYbLCV2d62KNce3H/3Sr5NxTvjPY/zjPHiUL
HNYSuNv0EZSM47fUMT3fZbQGqvAVfm1lV0xlcSWMY0x6whAa6kJrAju6lsifZvXi
7w7DqKEKzcqGhG2ZKsASO7m4FOx9Sv3v7ZVPIPsWwQEM9Uy0AIxgawqtrkPtsahx
3ycHKlyAN/P+NhLeDMC/skyB7jGIpzcp3zpQwHalWeMyyJnpM7ZmZ3sv+exzS292
HfUe56PUHwvP/tiNMlcKp4czYqcjuS5C+CqXpF7n8W3Bn6cCj5Fmbe6cSY/y62k/
uD92GKKqUPcZXE9VKlPIhbUIqh/C1ByTAVA/b+GzupVT4RBXSdmzYr2IrkQ0rzWl
SXHZLiu4oeHWleeE9h6eZoJCEfxF5LdbgUQ8rbcubsipvoyEJnaeAsh2jwN1HXa+
WjRJAx7+evcyXUirjMRHyCg+mnYWaqPOLEDig1hvqLvEYOhhVhCrO7t+HMRdqAVU
b9yD1TzEVlFMwRKbMzgvoRbEZYJjtsl6tt0HQRplUh0Z3L4FF/ehxwsJengzctVJ
UGvIqzcZb5I+xqL6gVeT2v0AWRF0mIUCp+0arsY4WlpZIXLWi3tZtFs82+zVezCu
L1FMWLG4dqQbjwUxLKf8PpBaGAXAltX3TYurOExYYy892F92+4HkI/yeqROriZrb
Wb+j2+Er2KTiphiZnwsVZ4XyBljAfw14QX4rAwpoNM7xnaI0wLp89u8DTDcVoPuW
zYgyoTkIS8TrwWf7DWICHysadLYhCl/ZLX5/GAV8jZSdeszeb5KJ9hyWkZHI4cez
8gXhb/VLfmG62N2azNiGcwjojPVQ9sUzjdZcnJvvO3IriPiJ5hZzBMISgJrDn0Zi
rqs2abdXs8KOtyOqzIf5IH0g7Y+4WGn1oS/3umKZb2ye4Lfxe7VmoxWMVk2vBfUF
bdpeelmwQhMb4ycIOtNPeCU9lcx6kQpyYjZgRWJ8WHaZ3S4Ri8XKPNE7WLsKrqPN
6AtkUmWk0z1dweP68x06qYEXxGTo7cjI4jrQlLxwGpoN3ttaX6V/YuXXWwf3s1Vt
By/E3eSu2ZMXYD1lybCN1EhHVc44qNQ4/zWHUbvysJdF7VC/BFeZIzXVDoZTjBaL
ExS5pc2QrHI2y+nxjC9Td523z9+dm8yeiokMrW/5vGSZRCsOhXN2YDzgkTx71dgG
VQvSPEh/QQxF2Y5nVoLIrC78l7PTGBcaQhwSWCKFOr59GTF+osxYbI+xF/sxz0C6
8QTAuONYUmkGl5lVrcR4b6QazMSqsVok23sRI3sqcptV8wF7RVut86zTfNFC6Udo
OAlwudcu8lirHlIi7ech4UpDhfbZ5tVgyqrjvIAw/TpFchpneAEFzyhVQ9oQd7jU
popB2TJr+9rNqIZRs9ZIe0RwgMnF6Hp3t+NEzPxsjBJk817PCAxQq/lxCmZKHYvT
F6B4Pwbu6Eim4vq2tZBqKr7TSSaJy+fpdkZ2CvBdV0KLiaHeiSFv2ZlZI3Orv1dm
KUUMScYWf60EleMfb2bIPb2FaKHHGvycIJNpKAqekMC2vlqgMigRPDU19qh0LXlU
cavhAHsymAMGW+y6bh/8ghTbouawOm7NgWV7P+cQeh0klb955Tl1HFtx7FLDav8u
nRBYXUWgdL1NpD91QtVHy+DkVETx3zmArDWSXPWwwNs7JZEaivtQDu49kxci12+L
YOMMfRs/6ZoZfpRBPv04Of+ZGzHQTujagZqJEkdNga4sQKmFHDKC029AFyFydvm7
I23aCsBTrl6qfWtUwgnZ8f1Ei443Q+9zEaaRwltaQaVmTFaNIv2GhcIFTW8Xv6lz
5U5ousFmCJA1+alIOJIhPOycZR9jI4MUfHOg2Q82See5dscTpy8IzHt0M+tHxyml
VAB2tks3a6aihcPUcLwRuPmekGbdHx0H/ZaSEpoW72tnve0OXYFq89duB4by7ocs
`protect END_PROTECTED
