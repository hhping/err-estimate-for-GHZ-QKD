`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dT6WFgPxWsmMnimvfNsznYsTDtq46eeLQ7GatxLddmfi4YWBjhMwqPSFUH7WOZc5
QtwFgfs9jk0gpssry7naYUGX5d45Pu+bcTwwhqbns/dOikaa8ACgYE2/piWpqDMA
7yLS1HINc4TIhguOJlx4j3SML0JvJdP1kPv0Im8aE0u+ZEUCMBiE1z5ArxZ95a0G
CYqrAWgEvimeYGmI4vcLZNVT7HKpr86LQP2W4+dSpMF8hq4Rifkpx5sJRR6/PWhS
ykeTBc9pNkgy9MgS5SCSJjnjiW4mgGvAdkU1c33K3ukdaH1p7fqvbtOSI6XfrAft
QCAA41gzgRM5hYvNTDZDv61HVorO0PWty/S/7S9Gf/OocnGfQgmas3dztqjpcof9
I42YxuVa/Q+Ga/xQ9WJ8vnYhrK+vd0/Jzs88spSLr2QZf6/ibAwPNu/cvzEoxF99
VgrNbXG8Zg9W6d4zMZ6oRn4S9ptnuLBO9vI2LJNk1jVJEA7Fk7j9HEWiASvkFbbR
tEpZ/VI0ixSvJesJz7zJ9TGOS0u0xV0guNvAd3hG7/xWS6ow0xjn2XvGrwWy3kPl
XB8W+jN9b+z8omTmbSh7+w==
`protect END_PROTECTED
