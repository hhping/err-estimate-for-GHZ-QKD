`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5pYEnQ7DsyqiFkFE+jlfHfN+JF0VtyQXDR9T4mfLOxZ/LGvNpnh76HCG5QQCvEoC
RcG9hM5VYeB8WSj1/hYhYBRN9l7k59fd5ftyS0ZBr+Ir/5TxcOkMHEgRsFXXJUSA
scWvnkxAtLTQ4LcrIMXZO7a6E09a7c6jrBzuovuMO8DNGr3+fNgllwyJgL0lkhDL
4t+LUKbjfZdjxgVp7+5LQB7SFFPcfT1UiP1ppqCzVL4eYKQe8wUwLPGMUoDdqiNy
4D+99DOmkMr/yUw082uvLvBS9TyqGktrfJNybA0Ly+7ueUK3t2aMgGXBbIDjR40I
ETaOaVuO21CpOb5LsSS85stctAezBXhYrKcibL/XwFithMQGCnGZ3HWo0+OPmoKI
EvC3L5fYDC3aoHGBvBxwf3RDYWct4l0FR4yYkwHaaTd352KlmC2IADiyuDgXIedn
wrxkAwfI65xLbkr0nTs1RAtnFFuZiK2bKzPKEKkb62aPSgTAOT8TlS1YmLK/aImJ
236rjJ02bHhrkN1jGM/WVOovcCmmScb0VJw6OzbHAjbXXCTe3ONAj9soNUGP67K+
lEDCBbAc3xmVG8CU8WSKq7HGRdqOcIYMWzCL5+ThalCr/dyhHS58eYC8BmrzJTMv
VS3/uejJrwuutJ76maycfv5accLwvg0z7tUFIBmsJp4SjAb665/ks0YT7w8Hf7rF
u0Wi4lfg50d8CpewEU59O+6UXbhWShBumdMEU1/HJPT+8awXDgEHF+yaJZszP+dF
zfXDKx+iEkEelDm4eH0Ee5pojjI5mvzChydCCWyy8LUMTMypN9QS7Url7veDfhLZ
CPURbqPf0H3bi88BlGNiCVWPkFHbo2jKqa3TlqY9zvonRC2mqrIuZk4Cp8Kac8/u
JSZcgQubXnt+UOd9iHOhYwqunahPD+wfxRJ+85kc20wVFHXJ5+q/0qItNM88BD4J
+0eNBY07cplNaWOCQLtKwvu5io5DdJ8vJwcJ7gt7ck+VkzzYybwMi7JQmgHO2lv1
tKoj0i8/V/9QExpZ5I6JQuQHY6xIipXqFw3lFHbX0dDoFV2wR10OfanqIw8Qt344
UDCCPDm9INWEugRK9/nfbddK2mqgDGnAxPRbWxPOs6hakUlghSbuW5ZD2WozkS9q
14L2Dz+4sc1U3z8J3ioVeSOROvJx+QVYB00Fxc+nHrUrG/VCq3OvqpcgLUNLWafY
RibQqUV7byD68AKcIJSH9Bv35w3A7W1w1pHODy6IstxuDe2TY/A+woKZRPAeWpOk
ytIx+M247CRPj9sYlWglUNaHNvVs/bMaelZTZL1L9BHCX3OIAoCSboeujkd1PNXt
affcGwGMhuTSe+0fCVmaK3e5W2FfuxZSWDrP3yRHK1bu/Cj7RObMT6E/I3M2vp/G
wTLC2ySxJe4jlD3LfXkKxA8UvS+aN70ZKLIQ5K8NeeeeMbAbEriILflDMUrMo0MJ
BKtx5MZwIeO0j8RyRNw6+9uAP7Lqr4S1hf+LkE+nQWsXsTq8w0n0ZstGpcg0zM3r
7nQ/NLsGqzIYGmwQ2Zx1Zdj1JbwufBHyE0QxM6cUubet3z0R8B5Ninw/H/J5Qa6O
DKqzE1CXR9+8Km8vXNPd+EakD28HI6o9hAaU639nUrpMvR6wqYTdUmjZW2mYUFvT
6qNc0KoBcJxL3GViKCwnfneUif+z0WvTWKzLUUlYHEI6oiwgZn/w6/+ELgC2D5GA
TXiAvZ0c5jBQQxexnmsHArjDnrkEZpX6z4lgVHsu5Jv+4FKNlglNCcj9jV93R+gc
3h/hLHtlnCB4Qk9qrmoQ7HVTGeb1SyGW8I3myOsdMO9xk/hi6LIkU/A8jfeYed1f
VcNa9THdYQq6LAg13tJmK88TOoItjnwyavGrVMipCABXaqgY977HTqedWuucPkss
LV9K86V/zhAsc5cSo1D93aZnHGVgnPmO+tW+wesMPW8KmQ3AfKVfDqusnSQhO8xI
9F2jgnVdmHpsqAWEhLaTQO7+sytPr00Sm6rb6DTx8ab1MAee7pcrqFnFQy6OtOjm
vm3VTKwIXbZ3Vosu8wJDzwI9rpB6WsFcojwJprRdVDe98CDD8Wm0RkocG1JlO3Mx
ThjTNx0wGcpfdNqihIE2rpZtIjV6cb1M8bv2/6fTD1wDUHMdkuUENvEM8S9wLnVw
TJgYyzN/Q5HrrGMWOrpokF2UhcQ11ygF1LPLVZV7WS4JZQC+boWSNCR0yicinDkU
kwfDTC/8aRkg0tYNELq2kcg0gWc5Hq/vxSeAAzCdB0YmR2Vml1YGM66B/f6Ibjti
MpqcW39VNE5sNKEoqe7zHd8xf+IjnuBnA4ZExJSJiO8dvOEyhGSsCq8AZz1GEQQj
xzjv7pRNxfNNg6cVnI0dWUdmHDce9VOZb49ENF5s2lVVhWI955vJhr6dqa5zt1nK
BG2d/c7v3F625dYO1Fve73uxcd6E7aqQHpjeiJnAOH+lJrkEDYefkrRzBywZWz8B
V9Pg4MoWMumKssXb2JuafqCH6duVihZT2MDy7zvRqgKYQhsiNuOQL6GNZCQLo3kL
CupG3Bl0q59BZ1ZlVXuS0iMjkuofe+Hdaor8pmyebpUaLru+d9LWnPkPTZYC6h06
ZN3jbCMejf1Ccqc1rbOEU+WX9XF7rGMcPzqXT6qV+oRYvyuPmwx6phHmB3t9BY4t
UAz+/XolmODHomoUTBXBEVdAp1oRAhPf6O06AAmvjglhazSup4JXbPOPSO217/Qj
IIW6T8F6adQakP2yGuWnHac14xSCGZ5cex5o2ypdekR7Jxx0elpJ6ixI6szReiSN
FvbzY7OkkZWcHyHgWPSZ8EjArOXGJDFKY6d4Szv2ZH0=
`protect END_PROTECTED
