`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LnCTMWKzfMF3f2WAHBe3YlcXw6dJDv2k7/oFB5JizB62X+PFVc9nMWWfh5WcubJw
hpO55fAnJxPhDHXBDcSjlaBz1PPo/I/Dpz72dO0OoFRqC3R1BjnjK4MIjY0DozvO
kUaWgsj2E4PbGbTEHZ3AIZ1Wm2+BH+bB5uoWkJd61YcZTV7Vc3eiJ+Bs3zk09OuH
qrfvJseE6Q0HtYFfml91dR9pA58HrffYoCRNVTwsPex5TZVZ0WoUMKmro66G91PX
1j+GP3qYEQVBLB4g9YLHQ3AT+3Gng2CglPAc2eEmEgWdcJ0i4jtC6NIeiaF+xDlu
AMOube97EgRresMNWL9kLlx3VoSYe/QE/L1LW7NCLAQP4ECTUMXumQbz7bpxX9Zb
3pfqGytEJAylJmvW1Mdu9Pm9Zj7rIuJPT2gKLWD3jGt2RfVghYaDICs9lDsJJd0J
gXzp+jDHRA3NqMxgcH7udGSki9aAqyTwqdjbovnHXoiHS+J/XSbHwEfACpK5Z46k
O2MT4hHuLyMsIgeIQkQa66n5bMkhlSZSvkw/6aE5vMXp03rDS4/7yhmatjtcPDrI
r6j0sNuvTcUNF2IgZLcjWyIVolFPOJHMzv6ftu5LbnkP7KMzWQFd7wcAXAhLlV8R
OQpdMsW7ESRgoYlDvqmBbotqSqHOeCYpFVmPIcUBi+B6E/4zz3RlEYuEZUkgmPqP
ssLM9s3JT81EcDc760ME+iXj8oqMFkTwr8vkhXTRmOK8Hx/8+Ob06XkISxiPIoSm
TePC6hzStCNUft/u7y/hm780xZxGmwR667nz8WpJ9krNfxab5chtHJeGlg1zsHV9
TIL3gxIWGQivXsIxnEvQQvWz27z6f6zx944Q9QFRcpRjklPx7dyQKx4Jva4ACjIn
txWyi9ZtXYGgXMC1zE50WViLMNahrBezjDkp498xDMwQfRoeq7DsVXOsRO/ZxBVV
WNoJGg+Je+W7Chx4gLz/qcmtl/PYtZmVcoow71fm5aymOgTWl0H3rcx9yReRX+bm
JVeRQ31KLitF0Jw+zjs5Zi+dwyQwAlrxNRTnkjmo+00jHF0N62G0RSxcTYWBAUII
FznMg4QntQGlnyeyipimFBZhzxabpz80bkDjdp9GCIp5BGdu+Af8guqvbng55TBa
e7THp+cW0L+5sTWM5bDOuOthfr2kerXA3XseFhr4DKseVQE9Rw3fnXNGfDVyoO75
/Voogpi8TLX7OkHOl4lkLAtunJvX4ee/pn5zsHO+qDoGonfU0/fPNS3AV0PiCgQP
Ahr0OOeogLSz+QI3gj6Uxzo+1F6GS79/ep7Jd1DNHtJE9sZCETBCklLai11fVP33
JExeuhoMnaJRpa4Oh31SMpcbc4MKM+qin8/45ZDvtyIjlEo3cntkYn2f4Y2uJ7QI
EO+RHogCX8PxAy5Ij1Bley6ySwc1Q3cSlUM+qUt4Tz0knkttDFGUpNmv+z++qZvp
soMdsAj3YJvYt6vBnE4lZowrHFd1OR2LCsqQG8KXKqpV3xDHX578VPtMxKSfdZcz
XiMbAoD+QMpMKvccBQOTFf5ozp6X2fSMwqlTAHSIyZ/AYfDFUC5Lc5lb1OlT3oH0
Jipss81A6bixJAvUwoQ8SWr5MbrbxOy3Nm5oKJNcoHr9iRIyx8iq2V93uhvYLNW5
ab7YeE5iv2/b0kngzui2qSHNnG33weqjCpDz2smHXIqzpcDgo46yvxVeKL3NLh1V
J6fjqv+KtjgLYstlycpFUyEbNZQ0PdYMsLdINT1r2INrAQCJTiL1lYQER0ODiUOA
H44nBziyFAhhjLRrFjG0ws00BDSnz5wpWsto3arome9dRSWxGPvVTOphVhZQE1Zh
P1inlPyysgX8fhmmyG5ywHyzRIsMjCp0sjxT6bh0U4zPNVT2rmbIkTCuzloGnftw
J5mBGFOfoJFVkLG126WOXOfJt0XqMAjdNhcdrnikWAL1Dr7vyv543eC7Su23yMEi
J9r3KKyDBAoWnZ8XdJDHg6OK7yLT60xoo5ptXkrCTHrBz57jQbbYfSqC6IbZ4/k3
+YJ6mYpqOjIDZIuuGCCVKlfTZgaKc19SbLqZMg0w8oMdZsISu3hmutl0g4KXGwwn
upb74A55/b0zanB8P0FRArcf1zIFuV6wTiPzeumEcjrtx37hY+YYicQbXKkIdxQL
ls64ceZYMZrrYelqqehyOvgPqZcHgo9f7WSUGejMKwdAFuMoXURC6RKIyXfAGxrN
d3EvIvaNbiHPpyYkRXuRiw4fpp16VJPR+hISSf26/VEhDz+Sew/KpUETiVchNKrF
YLUSADeSfew/04HNIIS8/+ruRtZuw3pyD8u4VWHXAn0lLMyY4L+1bVkObOghcQ6n
tQauLFaszTFP7o+DtaVRO8X928mmxnrRZR6nTH4dwjoIN9WSjkJmiWkil74/kqfj
EKfk8U2VXJDkWP9KrqHYoYkVE0PVzH+htAXcL0H+qSnwEN3CLcllf+73G39XJBw3
oVGCG42zoQk0pry706Ypdw8WNtAXBY+yqN+y3XIalN2YHQQw3KevE82wwIp55OrY
484W9N7NMhDT7eZyEUdPUTsIT2+MkTiR8nWaK4Es0CScsgSsGrS4q/XHgoyuscKH
frQb/Bjo24CCYsCjnJtZxmB6v/QM9wfCX2IivVeQlfnWZfeTSYgHka2KtN7ciCu8
WS9KJNLNPshVEdNsu/dmsflBHJuDjqhIc+IRDA5DaFy/GTmG/gcFocYZd6aW4Sr5
m4W4+SOXBgq5O4y03F4UJiPJNI0GRVP9t2SA8hbHtjzWPHy5zJTf9tgNGlIJUJaa
8R4goUyD77fgYOK0HZAZ94ofkuEqIAvcKo4SePRkIdNrS3DNZQZqV3MOrXt9cNa+
AshzGXbhD0BZibkSzSYP3kFtbnqlGlLNvw0HisAsuhQPxGErw4HOUWQknYq6KG+b
+hyXBrCrmcxMmazP/MbygtHLBYNGBhMeYqXs4si0LWnZOd38u2/wH6zBuAoBSJg8
7vBcpRzjpu+iovcYQclJmAuZszBkvYVaRi8b6PvRbkbJ2YHS8kAEkPBzfyRlb780
3VloU89papGRO0TuyxuqtC8Rz5XIPivDJh9q7UwrFsAUWTLh9/Z/2CHzfn5JmMtH
FZ4OJfGraWGZoWm58JteTYhv0If1KQHs9KNr5cuJqq8hCRiW0RHEfLTptLjQaqzH
g/GRIGyrxyxWvBZHqFTT+DoiKy4Ai2ZS4KXbQfpC6qnbHALRog81n6gx97maaHQ6
pdxQn51LftqsYcjcwpKEz2l0H4TotN6oPV6pxU147GKCsSdivXFZo9AF3ZKlcR0l
vGKOeHq31Dl5Ssa/dkNOWQ9enrFcLq9XDhd98dhDQUITYboqVMqukkSI4h70DW7B
FlAWUj/UII81QR+kqNy7r80/8pUXWW82OeL8fBMe8Wizgd5DEQDPpRJLMJj0GYm6
TAvM1+zauylTDntU7+F99taLCltJrHLxhwCkrmVTK3W/6OGiQ/7Ldj6wuqyuyGZn
b0/TH5KzDrv4MsuyXrLljMDPoOGNrvXPBoU47wcfqYtqsM42Zm4yzm+waNUGYdRv
lKxPP+o7u3vvX7PO30IkZov411gH5/d8OJkaReq8lc0vi6lxvo64R0zPRmDBh4lR
afMB+tQGtVTtgyRGbnfHtvRFsyqexNjNn5uFObLaEu40J6MO09vV8UBRPD7CvkEQ
MPZUrZuITIq3ZEL7CCzN/zgNzTO1azpPhvKjguTTsT/+ArunTXC1PR6LHdpDSIob
WvE9yD4GFLg7qN/yZmD7SktION3KJb/lhewStvnKB/tS/IYIc8zoX6kttM3DJyDd
EtNWyW/aEwmcQHVYaeR0A7lHoPa9uCflMQ3yDJCqjzLEdyHuj/g5zYlB2ekTxr2Q
UHy/B/C3ZbmVOy1jyLEmNOQLGl6WckMskF1Vb8sK087rnCwCSirSgXrGwQmXQOcx
0x2Yv+XpMpBnM4c7vcTpFJfoDriqw4QgidgZXZbOJjsvMQYg1ZJIVYRYqeUrG1lm
ARwrZRB97wUJKX7tgyXIUs6h3hvqEb3uSjA03ZxCvw/qe6UFR41okDBEx2BRALei
svVFI+xYSDIRyssSXtfuDq0C9hsUW7rbqOrblv0Y9Lyzh9c8Jew1NbbwneJ63GuI
UITmtkf6wxLwqbjG8bbUgqbAXyokKtPeLAtA1+6BaWiz9Z8+tyGi+2VOU0ejkAku
8VRsuMaeHCdnaOmu+0pQ6mmQXFPd62gKZi2XeFDh91YwF6hB98LpAjLxNTRmbRL0
9d/Pk5YRhOFQt4GI0cZdZMK0OzE1IakV0lVgPiLL1vCSJ5Z0b6swXPc4gAAb29Is
lJEelXWWIkwkpMbuQfYC5jEvLnaNxsKXd0eiprqRH8tg+/11R5KcAaMqh73kXIPR
5FoA0DXIz80AmkAFIrLlEH8TAV2s/A32hlpkLBpMi0VwRWcvJQkQXFsKifgyXLvR
p8eN/ZXGi0I/V0hQyHScUJqyPUvci1B3u6ep5tgRewd68YeBsefnIP7x5EuPgRuL
fZyDki+BLkh1fSpB6Ex8FAjKiVsezOkBPXP8i9AjzulXkH8i2v/XyxKNE2DzVk7x
U3tk/EWfbc+m9Sh+Pc/whaa2uzE92FPiNNVzuEEH+T7bMBoXxGOfBXdLd55pIv7o
oSEjIcrztnqO21fS/VHVJUaiMgjKIPLrP/gtfNjNDizBQqJ3nAK270XLXkkFUu8F
H5O2zUQWp7LxqOp6HkKIDPuu0hScotq15tpJ84JMG0mnKFiLfoRuHT2B1Sdz4Vxy
KiEUoQFJnYJcGIa2NcDw7CV7luF1YN/yP5f/wBW0GeK3yzy7DgSp9l2zuRjjYUb0
lBNaEQuCGPqLAuKYnUzh+xcouz6W5l/iiB23i4bqTDEIKUUItizCzdHhBoy5EJ92
d7tForkGE47qf9eIGmD/0Pv7sOHMHBKNzuE8+GkoUmq8r/NsIxAIi1g2XyCD5Gp0
DqSnrKh+4NnCW39n27UE99sygKSoOmaPRTHhS7ANXCFn34QNtQB0WErGPVgFMeH/
4y7h+ofxlc8T0SMW0CWO/OjpnNVWT8DxHlncm5BdFQFVAgrBikaEecaJc7mTc42U
mRkhNNFSeUVhv0liAiHtB3H/s1C+uEA7v0pHGuyyfr1vyRYZpyNIoiLRt7MP8jM+
u0MyvVqIgNt6vBWy8VfPGFII8Ic1Hmlx7QAD2fqxNmISvllOlCzdmLzyCTd5JZKj
L+VbPZ6TmGYrvFOM+iOgrOOLjP++fYW4NTCMs3mam8Scm1A3LYjnXL1jb19J6EDf
jYaMiUa1KuyTUepF+nv0yeUsJ9BQ8q6bM4vChUKyKfDxQ8MQa1FRtPqSM0NJapAR
lysV3z28lUuWKVKxHwKBCziHJPnk3xlJYv6i7u9AS+tyD1K/aSkZ0xnQtO8FtAir
FycYBQK7I467ACHrgi5JMe0bCzWdrWtAjlCiyw0nD26kbUJW1OsLXIXNhorR1mbO
SlWkAxCW4QBaZjZA4tuNQ3nkbBoz50duLNmhLEWXuPAGcYce+erFGoGjvUMKwSZp
MQdKyaDneYNGRVpVR+1iPjhracEu5EWEIdS3i5H7q2Ic+0G1dfcfYekV/pXwgsGT
ytgIdOtJnO2NKUf4yjVPw2Mg30LGqDBfVWUjTXhwnV79DZ71BR3jSbb5wcpeDB+i
UVA/blaaN3ojs1IKdU869U4PGF16H08YzBVhgXd3DTaJCpbDL/iFTXtTpqzPhZfD
08wab0iSJR8/SckodAG0B4WaX+egoi6iiIMVnhC/0pYuQtLJTGmdh6v0s+x9w3wS
Gi8Y3TFvbDdEVZmVI2P/Ug1IjBpuHm775Dob464XLYrDz/iOE5//vHSsCuW1kooB
t1zs2+RhgSLJFgsNkvgw8L1CgiOD6NpfUnIFhbLqUHxTXkMKNsQ2+PyfmKduE8Ou
jkIrLTq7IXZVv5+nILjVPsLLHWxlmcdjHxYtb1p+9qj2GZHXzGbH4MiPnXYGnvwc
xcdmv3bOl2b1Fm+SFVOq2BaLBTMxSnWrWv4IzEs7fsAn7ooOZBMzQaq9R19yasKd
7/OJPGNiYLqolkTgajIWBMI8TWNccQ4dOmRAZivSygciADLM+Gki2eelM1R7NbMl
Oem8mIkerhnu28YYLV1qn7pClQsM/KStXoRzO6QFGz2ZKeo86Ohmz69cOKxNIgzN
/FsmMF29deqf0/E0NbP3NEaFIpbzBSQCpjFMNh9+DXcbPGCiBc/HGOzEzK3v2p0y
hfxPgrZHkYNi/SkEU6Vlqk0lab3qFo1gkkzeK8QJ8XjAczJ+AJ00ciVS3U29WEpz
234fSk1NGxyRpt8W77ZQtOuLRDtflbyfA9A/qY6hlLZEyr6aEiQtjU97TsjbOrSN
PjZstbDCe3HsqAJQ52SmGUFWoYPAHOgwZ5KxJoIs6sWWkyBn9i0dk6vH9YctQwSI
Zux2odHsXokWAzzKSL1HXR85UlKpgA46Z+VdqG51/TXstyRgyWTcyaELm8vhkMWu
ViI3x/DhCq6mXT9PlhF9qsy1S3iyceyjnLLzCNvOY5VK/Hetg/lMRc0N2W9dTBNK
1ldTbzrF+z2FdOxzvU3ZCYwV3vzJjeR9Ms9XUUgBgnb0ZZF1J4CtvQWSkllMCdPc
KvqPGXZrC/+dMlgBwiqLs72pSmnBEMDQixeWnLyJwi6ovT2pa1Z2KcWN2uRrFe4F
qKu4GIczifvILqYrijd67h8vB1Zo5mul5egiLkxzJJKVVdcSMPS/iYlcQy9PpKLt
Yfc+UhRpcELVF8ux7njIVq2beoBbVS4V0TXBbeVi+ak5O/RI9pD4NYeWm7xtzlxv
/A40NrbiSQbR495rz3q3n2DbeFvHZuD0aozfQVZLB6MkWh2xU2bULF6IOVQtTWl7
HLONDTFCsVwoDc5PGqik6DduR8GcX6Rl17alktZK5YXLQjkloMUNbhI2Vx/ejG0d
Ik5tAWT96pbxQa49Fjzbw52yVaYa6wilksOdyCEqn/y2eH+012KI9LKxthb0enr9
//3VimWZUWVDc4v72LuNdxpu8PTSbYoeOjgLzol1ODNn6GIKje+Vu3kt+6K4hXLz
G+E/8cxLv0D7nsrMvAgYsepjkwUclQ+4Svq3cVA82xGXCui5OTarn6ZFdTFBRTxU
1QeTCD2VAku9A1oARoAB5FHO4DaRRmwkXuFhZe97IZkOFh1esFoFqa9R4xEBTngj
6xqTQ9n9scgk0NhlktDX+sigZukUU9mWHLuEz4nBZn7FEMdoLFfLvTBNnAeVp717
34cbRTJiyr0mVCaI+HHosCYjrN60cdkZHpJ45+eVEZEokyOBpaiwGIVzD9KRsWjS
D3VbtnXPixPZW0fP8PTnX0GFwWFfdH7Rq896cHG0PTFeyp3ye+4ny6DakQZ1EqH+
9X+Vq/rZx765FeZZynIXjaKXDVrCmqkLDPNP5bn25AE8DqH0NtI9U07Zbo+3FJdN
yJOMqfFKTSkXFEUBFGI6P/68VSSf8XLnWYy79pbYOcwthaqbWXuVwB7XTJXStMUi
NY0PrOCC9xnyVK8D5fRLpHmviQZMHtn0U1sXPsUgW9OOmrKMrneGVGLkGr+CL3H3
fxBzP4Gfq7qHLEdLa2cU8iiWXrn7+q+DcUYP/42SKt/dLjWsNiCjVsySeVou9FSc
1YRPIA5OMModT7e8HbWAcMd7ELKBQhD6FPd/NLPgmU1aXfSOLAfkOKOLG4USi386
xHXgca5L56pgqFTT6f055HKQO/wXYBhSmRvKTmzMFNdSWffZSUYVYg4z8MK1IQO8
rBw6PItJifC6j9/f9lJtuuKwiiHhkr2+nQ3bwlvUWT4sLHsGQ6ybCS8VDJUC6pR6
Pd8IESdhXXSTG7vsxj6tA9i/iQldgsXAGe3eE5LGbjnJM+fXI4bBNu7Hfeu6Y4f9
h/e2P/8oE5b6Pyc7QN70FNpkaYrZ4kbXnNGPVOty9om9DAZNAjqckBevCROYIDUF
lsnFl+bOAPWbjPsuFZjpjpt5S84Hf4BtCzrE86HOLhBObyhRfOdiES2RIVF/J5OB
uQPiq2OodFzGlsB8YQT5uHUbQVnzWWcwGmM9IXg7U1LbVFu3bGgMA/p98liYoRYz
X4CaUKfWzvtCP5AmJOQ9e4D8iw95cndT3hWt2aT4W2rKcASQzk+li5gUMpWvSbZH
yiOFKxVm4xOb1mpaUbsKBZ8webFJ4xil2CY6XmlEEA+PYSHa7tExf22m/nu6IMf4
95+Gt/tyYm6XDrgJrhzf+Gs+0APuWoE/F4dfx0DkpGUu1AtmMjZ26jEbyN6MYqEG
xkKv1yRW0eJ/XaPhnjrrZotnvVRgdyY5lr+EgXJbwO3FLqppACpKgpUHaL6P473g
JSa9WZYG8liIm8v3Ffn/yb+w7fEKZ3DKSZ6v43vv/DPMLyfv2af/kUF/fxMv0lya
CgEav3OkU5LXnqKyRlKTpUXz+eCOOazz7t/OMDadj/YnPLGrLUwiFrZDcBMOLw8q
skYell37QlQPUl5XEHyODyilsx5gz4cHs3saOY1AdTqXj7zD/t61Q8MAqr09TzFL
djjLTjIF0Mzx4Z1PIR752ZQMl5m3/4Gg4lv8OmRLcf995siTFRcxnSI7siR6rfe4
dPrIRaMinXJBo9zY1Fq1PPRIDmCkYAGLlq8MX/ImZjjyifL7Am2PK0fadjgBZIaH
HCLqUbFaz4bcEBn33twlf46eBsCKOSDJ0gcByo+8n2vDHOc2OmVSMVWV7o8yeBV8
HqnkZ5N/NBrZCBUwfQeMmtq8XaAY9ZYJAOgF31phztcbVcJ6f155GgZ1LnJsUOvZ
TJQ7Zx20aRugwke8EiUNXyGlV8GAqNdpQzda+h0bff1XDfpQ+YdUoFDH/1oLgugb
B/8MuOwbe9ko4wgpzq2OTnMnvZMs3lxoE7NcspBlbFJ6Qlky9J981IX0KB50FG7a
etqcqBwdn5jv9/mivf+Gk2+rUkRJ/Qvf5/2pxoRxwFA3yV4AzgzgP5hOqagEiQCU
qc2jZCRLfpbT2OLpHSeQMwmD/ycg+jADF6PRuhWx82yGjbv4hgPjUyoPt6aGhDfT
LeK72CDOymyVJEEt6yLayc2pDk1oHs8CFRmuynlWYnIuNeadJvYeDV8zOj7jq9Pg
0L49z463bk9Qb2fFvJFcGvMgEa8tnlK4/9v0FKSSfqlCXDhhMUZMvjiIcyOUdBRP
foJdgbcw6QpQ15+SyDdOiBK74TrCk88mSxrVc+/IGXBXpjD3Db1YSTfYsUbz7GXN
jKQA7KjxNwRapbj7v654l23/nRHd+9kuxM6L8FeHcl8LssnqXE/XIY1L9Uuhvw3T
yBdycP0bA+R4URSUF7HrJ2Mq+e6fRRI24JoGgpI5h+yR1iUKr2GdwHQJTfS/AHGs
Qup4eAlsVnh2Sg0M5kGizOw4d/cmBYF7uD4GD8sEEHONs/IssQgEFYpWlpG6o95O
0HkyHp7e2kM6AF2wlqrQnCYH9+FgPYmm1AFhrC8qgbs8hipoIAH5MJtnJbxSxXTe
iMaXbpq7ZynVLZLHYEfOIpWJiyEFYuF0OXJMjPZaNsqW1JZRuDhRlAQtBq/abLe8
3tBhtQPPqZ1Dq05bUD4sZNiz/1FN/xQHtrtTh9ONfhh9owPmJL/skU+DP6WjD1sy
8OZqnPm/l5Js3U53i4XUmQhJxn1sxv2hpvyZEN0ADVrQSLykOWIHjlv9kxB6a+nv
ZM9hf7kfBrtx5WlE1bnXXgewy0KDG0DmY2HPGgKZLb71xSub4iPh9attueLe1MH5
ZGIXxNuRFqGvMtyqRFHDfpZyhtFUP2oabyrEqgtkGz5Pd9k9/DumxPFDHZL7+YSA
QArXsIWB8X5VX3ftmx8Iz6AS0Rdkhyf6qme+6evCZQvRWfigfDSgWoYsQyFksePx
bTw/H6PElc4e0TZY8+7snVVkPkXMvkX1LPQ96ag7yaz9Ijz/GI4YUDr2M1hTCMkd
6bHqG3/c6SFX5JbHSFgxIGx0Af2qgqJZwNidvQwxFoBlsw0QA1Am6BGwN3zosorp
YgsqI/QUtlBUxdobXlQ/Qxz4SlcdIqly1PwGkt8iUpFHzYXUhWA/Ic1G4aCXw12/
R2UwqjbGBOaUx1Uyq9Ja8R+c0sPJFcxrJRqWWESTf7ySj2w3cbIx100iCv6bBT5P
enI3rr1F3zYFeBBxb1oOg3Ae3ZVmypKmYUOs/X4HIVRarW/c6q3HtwD/JauwrZAQ
5hYfIT0bQPU7MApRwgSOKRG1eJ1vqwl1td6C6F+CMIjiRUhFi1k27qQQakbargKH
P7/l1j7HwCundCIpUbK1d7t6JOJwYGUiCttzb5qFBFehN0vRvMRgORSQLi1e5G3F
esTSM+BRYUViTjVDxDY1qygQh6FqVP1ecwjridmP1A6C+Yn/XHeBBztLWX+5To6l
UVpDGbJJXFOkLNZHILeicGlhFJlTb3WZHp8jJMVWxxyv0ePjnfuGuHfF8YabEkrg
2RKZ37kA3JdnI6ad1u3fUsXmcITCUEwGatP2SSWo2hSF0w/DMF2TfY58ur11Ay+A
yzGF+K8eGMFrteJHyFb5x8xTmAKnWiUa+nx25xqVm6JL3/XZTFZN4RJU025aEgH9
wwSXJMfX+r7qkKx3gMEnDrNVPJ02vSf6yVfQbslP4qcbgF/OyE/jiS/M3OwR5hJA
vHKJrCXqVIQZgExmZtyAr3ajSygLeiOckrFgVL3J0zxSWBhiNF+tWbJ86ZCOTdSA
RVsAvPoKCVIFw8LfEQoRHNyJAJ+mSdk2YkOO54WcFbQXXBQlFfR5+623Ax9O9Le2
5CbnxPJTTwLqmTGGIS9LOKXoNYso3es4fEo/NaKBnp2HtK1yo7FWcPnb7dO6paHu
R6Y8OaFbSD9xAVZWz7C7LnKx0H9ldDkaUVZBQ0D5UvqRZk5GpxuQfktJytpIdPai
XWxscwzr2bSU8bFsbA/dSMILJoz6izB87raMlT2EmGQt7jraJiPZ48EY/yPllzpG
wUILR1DjjpWXQYjl4EuNKHGmBMOfeslwXQJdRnPZfCZgZhJelRG19DeFnWPC6RVZ
6lZOTQAxT1+BguRNqLOIc2SufezuMlvT98Yr9eH1AfwMvC2rB8xsm1/CWanZNX/P
roMN0N8Cqt3bLwhw6tZPB0MLXzMo5/qOX/DN8vtrdtXvCGpSTWcPG4XDdhQFKWgV
n0uYqpujEBtdpNrElggN4q2YuOjcRFCeBzktCOU3IeaGo6I+MB0hXj3OYrwbqltQ
Nkozlt4JTxe3/eqMSZLolgaafCQRjGBDtndy8wZTwKt1TtcWWEEgYGh1zBqKCHw5
3ITbYGrCdAp3u+U9YfmGz9ofClqta1MEwjE9Awit9kpySkqCkx7TdUICXTNH8ePv
XBt6PqKE2YpOlkDZhBBNiuFNN/LAw+m8miCLrt0Duk7GReup/O6E7b8jb5oGVmpd
TNZhEhFG4o3fo8nXrb0VaZOvfJeuSgnFVX+PNvo01KJhP1w9uhALW71JEaxkskL7
qm5d3LjrcsVtTBOVH2W9q12bcCFT2MM5IwA8QGvLoQhiWaWNg9ls/LReK2nf8qRB
C4Fs8g2oMHkYqLf61hCzoCEplNPBbJbiA5Paev99wpFB2aKtp7XOmbI3O298ll3L
lyBkIjNy+eBHvsGaQrdjWSYmeW3gLnDuRSE0RsoFzBZa2//GjbPkkaiAl6z4XkGq
Wo3N0SANt8jZ3KEVbJl0rQzSBi8aAa2H7vrrjcS7/zJBa0SzRDygmfQQYE23NLym
Q88m5Ade58vag54lpI0Q7YZFbewtiwsXRtsJRUG1wpNAynsQ81aixkDcFr9NbnPH
scTZ3kxBM1Qi45TgDMiCT5KFyS8ih4GhXIaoi73NhplTprKS2i6t26TzLd9yQtvm
RbVqdoOXX7Hy0ooKm6iJupgOAuBSGAYogZijT+1FkG6ZXyJAqrYUKefMv/5KgF/3
K3fnAPNf5mWp8BHbi2NDgcgjCRvmEQ6aT4N1pUBmR5b94aRewBqsMhAAmKGRIPCQ
XwZjIyQUaZ0ufHYxoxv7vTpt57t77XBR446LfvdEmMpGFSSWNuO3dPP7RvWjxtAw
uSnh3yyFvZuhyVMBPCIKih9SbHS6/lJezO4oVCuZ72RAFUy3Lbv/YhR1YAkTS2c6
BsSXFwFeD5X9/yT1+ADXiZyUexYIk2euTgPnd4PgNCairnrsaM54KQ3pGCw2kFiD
T8Cg8Ym2re1DY0lap7DOye/CvFmKXJehJ0nVFZRoNCdqyHMpe1u0YMNloxF7BSPe
wcLHkuceKnWycLgCl77FpIZ7l6u2RQ5sgNbWYWjWcSKIMiBXnqEQl1dkJt935WJv
SqC87v1oydfifGbd7ozfFZYhxEFzLcjv3TV8uT06hlLJVlkOrQ9fIVKC+WsvejHa
wwoJg5GTStJRHZjpgDy1m6kWBoWFNWMkfqHDc76/aKDcJpAUUhUMxfPv/D/ZGm/S
ZXEdGpZHJaXvJadK4f9Dx95bkirAaNIxJMMEKtfgTMPxqALVyfLCth3riOlw/k+W
vb5dCYGbqSc10MddHZPdIrc4DmfSjIHD+8EHVwYs7ltzGrnREOXXWeC+9baFUGOP
aJ3MX3el7nqJGwdVdha5r/fedE+G9Ft95qr43Y+2zKtaK0wmpvzc9KCfqMuE8Rby
Mcs2vFH0JUd9qdbguKyUjuNsqi8AcewRgHCi3A/NIaYymCqTruONFXxUEGriEltN
qkT9XMpsKXpAaLFRdLOux/kBR5l++ZItcCudkagCIcctn1hKhVUb9HEqjYsJ7/km
NbxiUtotyZ/t49c7HW9T0QPoJmYX4ASVtPD5HxSzpu+yHHaGAfDy9dS8mISt+z/x
yMmfZ0Z9xgekuPCdqHNPko1MLI7zDIUKDAh9U5x8/nuz14KpbUu5Ua72nVyQnbXW
EaFpbBEKBU05OKNSf2sZlzBYUuf7z6p8tUBKjNJNzFBxBkCamoy4Q5N09DHjtZd0
X5yGEer2anYI9eP6Ul5NV3sBo5eM0F7IwSVD5/eRP9oojyAw+D68bKQiAuwM8AgE
M9n5+7qArbFUfb5V1z2StOSb182P13SodIoJRyX/SGmMkEP2yf5oohRTyfqFsASn
4LmQFzm+QzbAz1+sOZ8vCsM8cgI2tLgeVS0KFMRXephzfEKK18rhIT3zNFIBUCHH
/gXAMJNSCOUAI5yM/5vel8ActTGJwWrNWO6qFnj3THyv1wMXnNy/o//HCcgezjvG
peL48aKa5wTL01JOFFemNdlpUYcjp50aaXJLr0m71i7tH0rWKU5Owy/BHeCkWxUd
dSzNkO95Vik0RsHZmMzNUbMgchFWPrCt7I3UQdrHXoN0iZbwD4DQsK2iMcdxjPts
FSqnlke7Ww1l2aDQK+zsZkc2xBxWzp0YgNZHDwJzpMmkL/biagc0RR5wsUTkn4OK
gOUiXl4asJrqAVe6m/h79QSAhmtZ5wbS1ibFB2TG3eh2GagkbMlPXZhaVh2ty6WU
r78F2Hiqfu5+DkqGkW2r4R+1WVJ8zWA+OFcDXH+hdEjO5QNwTrUNFnFUlSHoyTkB
ja0kN7iq4qNj2+gA6chOjn7br8iIgk41TA0U42xxa04OjgfWmCAmiUaE3YixTtXk
jYoenEuo8Ln9vaNGx6cl9iep4NkCLwZfA2VlfmJWVf1cjGd2q2BgfV6RM8eq1K9s
M2C+q6OhgKtzRaiM4DgZpkR9b9wtqIKHF/eTHAakU32P9vAusdKlCzTZIZDd2do0
NP5ak0VlJTU07ybyebJLfvQQOS+faKIscgXmsHWQX5cAdQXVGPtk7FqTBgdaKKIz
U05lCi3zgNdCb+oJoIr/AgV0LZIfUlLDRU1/ddtH6BaMVeGcy2V7JtTfIX2+hkWP
uMPFjiOQKYZKh6vkbpvig9ZR6ab6pr61ozTABCvdkOM1mDkgLre4HOU7A7aicJ6/
jZrcwAHPqcMQCESzj1Rv8n1HI+pz+3aJa/aPsZmgAPySkERjEbi0/5gxYY/T5ZbU
ivJg6zbLq6c3ytvRNLR8SvzviqC0fUUyiBtZdgr/HCqd8DnsyK4DGpA9XrNxFSS1
zXKULEiwCzzBpjbMbtiyRKB+Lo69DJSFrX9tO66P1bUVJCPCnnD7Q82LwncROeaD
DA8twkyn8eANvrEksfQBdHxly4NuQ/UZ+DFFPxtuqPI8mkaXFhw3qPXcPxrhnSHy
89euJxFIN6/6Gj1U/JoOflN89R4a23DUMqRsIOC0b+lk50ZN/kqBbOhpOgTrJ0u2
qB8MmUVQOgtWExsJyp0e9qR5XJ+proKQLzie9aE0rnAUS+dbO+7gldiSo+zVGT/e
LX0UAahZRn9tt3oa0KvHa0Sfg2TddJBTGLzyxdEjhrOZeNwtxVnAgDJ0Z5jGkwzX
CZcqmR/I/ThoSiWjhqfzCs2gGbA9hQfe4HCS+djwfGcGS/L8Am5Cox/n4KvdE87N
TT8LrNgUyBP3zlEC9C1HWjQLXUsLuGrlqqfHG+khwBsDw3v+WIBKQhgzDmSaS9rq
JQ5+PVtripZoP9mmVtte4oAtdLtWZ63aqhqSVtso9fwEe9Qg0xfjbI866glH1jWf
8p+TSLFRjMKt7Zruii09kxcTFLdnRLzaX/ciJJxI+aqWrr4URazRm+Q3NUtZM3ts
h3eK3GD3PqRV1svjLPI3+UqG0Y6GWyMXjg+51WvV8WMoItj+JnUZagGIse93SWnF
uSAtRqTW1wddqypE04bI4BP04aim/CAvoIiIUWkpDPNN6V2gXxJqLff4WrO0u9df
bf/wlsNnRIgA2tuJmC0eWhY0mxyIoIy1qYetdbzxGuc169rhZcU7Z+h6xLDrKO4r
/cQT33dWJOgJZTanN3PtK/9ArZKN5Tx5BLyU6PRqF4CQs2+iVMJ+l+MMjI8h1+SL
qRgCRg7QEZahJ6/CAdiq+zASB7rBoCExpbAGSNEEtW3aDVvoH2nW6clhO+teOLkT
VqNtHb+4GJjtxwqLuN0FaFIJ+0VG7sigrp+CRg/F2rW2/IpSmkF6MsjW11GEq35S
zHpGdvRUgLEAcT775kA8D6F6MLR3P7lQ0eLvDvjPh39H710Hgrq9ZHEJqq24/HMo
mLhZ2C3wVLVsfDXCrY9FxdNf+1TEFqi9+fb3a64/y7YOPpVJdWiRaXNGTW2FIUTL
ylaYzgi5KxoQRw6T/cYUVYH4GYjg9BkkyCwaOZWwykxo6S3SV8m3S9ZsuZZtu23e
cSTK00SvuCsB4uQqHxD3gHr+iy/L7cnBWpxUFDi5aIbSXT33PQJFx7gJrn5BygIV
PDFVa/Wihe+vKvcwDbVB52fTYI2QZ1tl1G9QoKV0x/LUhtoq5xMImG9jtSKZJnSk
Gnl0DL3hN9UlFZ167Y98Lj9eZWjEgvCZ2P9qlv36v1K8ejOuVrjRf4ly0+4lY52a
RHcYOMxnM5SDSAM0SLbX9aXGq+5xhM4xFZlO7MPP7eyNZ5227jq1Tww3pFMRM0YM
72/+wFaaUzzWjiQWLXEGMCNTg1YqhxiHyXdBM8++6wXRqDpjo6dv3J/bs/hRlgAf
W9g48mYJW1jzPftXoUHkQmDfdx5+MIYjN7l5EiV+KTuMymbvTTCWura2Fq4S47ns
+QIC25HW491jkGkB3nt3XkNGQWFtYQOnOs0k7/BY/jf/PjDVo1pByUKH6KcZQTqN
SydtMXEt5qwaTn+AMTP6OAIb+HzCWjsnLlKBEDX5n52UxtzxgmDz0LI23ye70Ycv
lirXc4G4DNqjsiI1GU/y6/owWyZNneUJxTCqOO2jvG4SaCTAaZRCr/g+cyaJnqK/
XXhEP4eAIJwgBmMElC9l/4WoDNfQ5BaH5vP5d80Izo+CqxPtkEWSsNP4KoYVe2fj
dnwTmTtcLGeY2tnVpqgJwOs1kgdivYmtJJshRIaJ+6wmO17EiCr34uCQcDsPhhuS
lwuGgVlkoWdLU3h+PWAvoBnNHHVUlMdGYP6UBfJ5IQRda7zyt3X2hGlscZoL+Hnz
1MrWvwuVwj7rLb/8KqNcRI4HSlGnoqt3kqttpcXo1sg1OBNQxVOFiLPWQVP0RAXC
8dPr2kUZS74t/822qxjFYSLBApAohJhr2tf5cxI+QCQH17AUeVy0hpe6cTPGNBsq
N1n0xJpFFAfyPWgn0UKya2sg84tGl/GaxAsGQBvj79F9rW+ll5BA6hUSFYp375L6
+atgiwJ/PqtMrRsJEv+mxzevGO9p4gMw35kk8XgLfL+ZrDZquGc6QZNiYqkNEzr9
uW6tkqeBh087TvBze2GHVou/ny9Yv3d0fqlq570MFDL5uzugaQw777l3E7jHusli
ZTJs2q/U2kZLIaEegbcG+WCKXfqnzwsGXnBT2SKOd0UE92LH5Rn+R56UptaiFaM1
Rv0c5bbsjixSmNJTQPgZKuBGSRrZ0MyJBBnznR0rYHHl00sAWSGHrso5fxr7Jfyq
1EwT510iUfJ9UhD3IaZotyKTU75YuIX0rGnn8frV+5kX839yC6HF/npdBv/4ITfA
DkY79pF+Q4HYFXNnuWjZby/18XqqYn0bTuV2LigTOlP1rY6gmG0rzOmLgJC3IBtV
/7Ga5vEKr7dnXmFGWcFYLJteceUsrdGBjCeFRwpGeZJ7stFkznuaxBLWgjlfgWo+
iOME2G5rRSspQCCKAoYEHs5n5B3FiC/VeI1K3tXmLhKXHi/JYdxzeGy+E3XCN4zE
9+BuKwnie5ZPY9pu1I75bh05elFUc//psffZ0PvjDi/Bx24cLBW78WH4l9PlcMzI
IxdTot6EyiRrlJFmwNNNJArtieoPSNV2kofSuI+LGebXCXSNrCQkyl7LMqGlvBhK
ET5j8PUcVEMxr5nFCKfNFhdnUdHkOSgh7woB/YQyVYyTEpWSLIU02uGRcU8Ehcbv
FXBpgFxEbJ+2IGzT3YeuY62puPKFL/+UrsLGTIcaw15crsr3HWLhCWqQvQXMmJUY
THiBn/fhVeEtTClUJa44BSNU5tQ186jmYcRAAJkdGwqHyN8GY0xFW0rGT6TYe3Hy
RRSHeoyj5cka6yCDJczEnNSPXnCwuJZxTHroeHYPGBRXsqDrzk3Pwx6qOX9nYDaC
zISzoKreuALh3YDiBJR1qOLh0aK/zG5rCbYxBo5l/KvjdH+VfCLOOqIknd/XYWKc
+mlqiTz47RUBg+harqt26MU8olF0IOMzOADkWgekuCxcQKz6C6k5Dw+CuUOmPskS
lOtn+cWTcnZX4ZIik/dwZsa+jWIt0WMqz7ATRoYCOmWFAISgqZuX9s+yCZykdsdA
6llcBU1xrwkO92YLBR51xtS0FQvMihHQwXxiSbHNrPQR9yAP7SM6x5tXzgLE5XZb
0j0JRyUlKA4di3KUYtrN82JwqWKhUncL9PHuBbEL5GwcaojZNgsUXCKiTvQUvexA
5rT/zZJ5yM9s1V7GzynugIxR5DKIjSe5suNxaJJURWrACH+uX+66n9T2wZGwuJsb
tuDTmfKcp/elNLXojfNGLRlkKd255ANYxXA00HH23Z4AZQNUkIC2zr4w8aef8L62
B7reP90RU/KiTQEbMLIdbk9Mpi/DnetnzlUeNMuQTZ8cujEaa3BSN1VHkUgJr2Or
perqyNmvU/blNEEMlXiME6OA2t01KP15BpWLOxHx6N3PN4sXedPf37qRbiKqSuKR
WALv9QovlYhx3u9WLu1AW57OPcCpKpE+uiPDeG3I8SY1Zn8vo42gshsl5chtPzAa
SighKtA0zcKlVo2fGCUspWWxeSJoDBGmON05iQy3XoLrmjGCPV+xYgaqIA57gnjI
Kr4htG395BDsUHJ/DLhVcKhW61antNxsUIfHOfaLpW5jQmW0UXRflu5leeb2EGOn
E7vFqXilDTp2nK6yANZVCMyrkvfpFM2JpB5SD5pUbrdNATyIAjd6Ryrxn4DfwLJb
ScWs8UgfAJ5/YQjnzXeBC69FHXs3cET586TlSeF9P7mTc3/x9DkD/eQ0rOrqaDyB
4UveYG0pKQoR+v0lP76TCavxpNVhBieFW6JN4/2HGT56VfrQHqAv+cj/ff1r6OxL
jrMwVFAE6QB2aoiVRkTF2uObTJ+QvFZuhACU1SxFQbg6joREwcm3orKxOIlG78ou
QBI9vferRykEBcXEDLzEQ/pVhQ2LnQrGgqukYBwL+MCkANZHSxBtIqi5soo0NuMk
0BH2/vg5R+ZPUa3GacARvUFi4HNkzlqzgWdk5CrekJ/O/vj6jWRB1FdPFQ+9qXY6
m7xUEvHjg1ZPAG7k2ILpYLwSp+1uKknB9t4x23yGDouyaJYSffUmOG+Yd4By+VKV
7TE2VhLL8nPBKcadcJql+6hp3OuG5JC++ugNq0g3tcP92W8QoN3ygI2xiZxF89pz
aILZOJ+2+7fKXlfgmVVpqKWWCe+aJaWIqYCVNl1s5uYeOQO1dIAv/wDMafGop5Ni
UdQVHYifyu5rjiyOX16znofq4cokk+n6JtLMquC7CzpkEje9QpMMJAvaLlWs/Vjr
2M+CyAwTVYR4ia+X8qxwMW7g9dXqlaamB7WigZPfmnaoZkdcfsLcp34HfMQcf+UP
uSBux5akNFlIkATVSQveUEOfyKxygc78zn74KCvSIHIYx977gKazUPTbCZZX13su
TmKJyld8yHgyIkerr8Y3R78/uSEQXarFVe4BLsd0iby1nR10IZXb7uTsG7L9hSnB
h9WM1/qXkxZ9WsWIiEaJJmdl20VG5R27bHkQm4TDYHufP0jQCAQ9n54+2os6o4ko
TMFqlT7x5x3IJN77IiR2bzBk+w22VNwk91BVETLckwfCddje5BdbPIGv+WcMeWTC
S4GD1n2FVht0O5sqJyE5ic2oE4vLPMyVFrRXD2/dHpnokJ+PaPRqSFUfY/RbrS72
Y2nDMARj90wthOBwf+uj4phzC+ORqh7wMZ+7gheL7JTF3U3qfAXc9UJnCVdRsnRp
SvzSbsvWxdgN3smOXjYYTVdvQw41m8EZUrZx3AluLXifciWvceBAbljGDkvTrXln
PU9MCIxeXDC/mFEaNKIrTxA6SLDV7p3sfhNomecRN+X/inF3nh/pj0aiWzxarY17
ieGCNVXWB3dHgh2pErSf2o8shyHEwJHWtJWBPy0Skm/g7ylUQlpYLVUWCVXMj103
SL9WawYlIDs7+KOotLnsKIvgyhjZVLlTeoZNFlpy/PfmegzDlLo3h7TTGMGHXdqd
nO1qIh+1FRp8+iS/4L4pUCtIOLvXVc0BmWeyldBtiHEvgDprovT037ygukTKFfn/
DoPMYL64u7alLyh5j3QFiFHztxNIMWAeeq2gpt74R03rtNnT1ZckvD28uPKzpPAO
bmMC/8BdGqAycpplIIj95OyXHlJQI2Eo1dISjm5bxo/9cBv4/2Uz9/24xGAeclHf
HyD/fFeLPbrzPE8em/ET+QVmy5iJU7jVtIACla4aCsZ1KhP9mTa8gr7mKcnup2GM
0FSwDSwXbJXYt2gDdWh4BXzDexy8Ve1AxID2VVpWPXW6qUg/4nElFK35/ExbWBI0
NzL7s9q3oWFn3Et0rTLEZGRmH9SSkwkfUl9Zf4vDjwT/9ahs/cTApjvNEeGdwLww
k2nyhhaOGyrZW8BhF/KOExr0Mg+Z3z5HTQ9Xt5a0dboYHeoD98kvmhueC2ZXvpAG
WACDFNQzN0vwMDTIH8pBHTHdM7T8eV1CXiQbGTxzSrmwhvH01mYg4ay3D1cWugXE
5CtlRglf7eqV2KxAxifiCgIPYO04/IUAchfF+NCC9DaYEod9Vz+DBr/yvtGy9hiN
+Wh4/2RHRn1l/0qw2m4NjEyI+xiXvVefngSa8wjiX8aIIPa0xUQ6xNKSKECJ0UNv
HfRAWjSQjLVJ2rpsMYp5VPT58Be2eMFDpj7GuuwXWgcbz/r7tjMyBARTp6cT5/BI
yGflxLfCZCSLDVOO78YGcMmqqWqC0dwyAet9A+LCzU6wg4vkif/VS+NeBonYtEoU
BD94vnBKn+GecMkvu+4bO+YaXOuORiruZoe7zji1roSFSGNUFYVoDGqhVpHNfLAc
3pw0nRVe/Vf63phzMpPU6mC5w+iqH5disur3hek9DCOjiU0EfZLDH1kTi9H2gL4M
3ifrb3AYEEG0LSigC9iI3DJJDzx/nUGrGRb5lt+QyTPX0dBmsc28qzzbX2RAx2E+
2onQY3MRcB2oha8vZ8utfKJheYDvRYMviY4QqCwU66ztFaAHambpxa0pDYCu/Oiq
55+As71cUkA0zpCIL7qL94Crie4TAZRQNtm+sGbVxhYiCYTf3IZDo508ytzn7xlI
m563h174x6kOTuOqBOdbUT/aREKSdjim9LqIGa7aGjZjtIUzTQuOOP2ZJBlb4gRJ
GuWdRSbobV9QAPpUhk8AzTclIcd0bVmX6S+SDyD4o9zXU34Xsh1ef3DBov11FDsH
dXa4Lp2UuUV3CbyEiWUFbUwnxPkm/1D0ynFK5ySToH86SZMxJugyCFABl5aB8MI1
Lu0Uf7Hy0ophtdzGkE/znk5Y1paDllehZl7+64OCb3TX10pYzPxXLRdEoaK+4U17
5CEJUGB6esOnkAssiaV1ab+EzQyCvmzymGN7WIXBfihkzOzaNoJAqveoly/QhWFY
Y7SkHyb5LmIT/64hirelj+CQSzwMi1q37AJIgzChwAf4lemUVChflZKw88EVjiEg
zK/CunxfUaqEYuePO4ilZ6IANbNxJ2h+l4QqtANMtPELUTEJwJ/RNhTQWLt8Z7hd
UA0UHFXuUxfF7NHvQGZrizUNh5YKOAUPhZpkgh45X9/wM0gB74nDnizUwMzbXdV9
0lNunR9ePph702/tlnauioFbwcHu+4S8l0kk9Tk2Y9JSmI3+wmt15JsC2Ncj5kG1
8gIyuoSTEIlNqhOGDhMEX93kDWt6cxbRQgyxgcYCPqc4RGscoNY1kw/9OfY9nVQ5
WxgwSusD49We5Jw04eNEyJjDdARLkyJZo3TazPyfWqA89ss5Xov5Zw+sYBALPcZD
s3Qkjug+L/ln3CeGJufhHYQ/i6D2ltCzTsEsNdFXtemaBP/IFk5Chs4OwXEiP3ub
qNQevCjmaoMa6/jT6+Y54Be7ita+zSl7rQvzog0ygei3rLKyWyoi6ZP+wRgkI45B
dgMvttK8255pDdRWelZmvkxw6Ak2nkeNbksn8XVyckSdJwFo/GF93z37lN4Ydogy
EU0EMbpUKBIlyMqxpihL9/CmHpoNKUOKfDdk8+fRYL2/Ii+c4jrdY1MEnS9hij6a
ovJoGOxr0S3olIzNzF8kujqu9IFkdAsGQdN0O77yi/N1el8h2fwFBV3ecCdVpU/o
YfzYYEmqt9UDU5rl57zuLN6Hi27QXsatsnA3hdXsuAei33beDvWBrk179nAi5Rs1
12ocK/1yvSZpZ+ZZnEXJOoct402zKJeIuv8NeW0jex60m+IedNY78FdWUK1Arwsq
HAKmn9FidgZH0cnK7jPx70i58oPS24IJ6N8sh9J05vxaF+236vhFWZ7h1P9lfM35
ZKcrzGI/wbnVlgn1FSYHn//YhvucsMLUBwW/ExcSEnjhcnN0Pbdn098gkuObVWg5
d+hJOwsEcG2SgMhYhIsJdoP247v/VUQpNt53m/k9W3UJxkCFhAMBPfkOHfd+00tK
vm35m8EreCICTN5QxQVr/X5bT838HchfA1+tFAB+z+9pyMsxOBd6bsIXawcRNdDT
V7WL3tCxdMYIZM+aCCoClL8Y7VUfB4iy+E+wqKyKjWcfLz8L7Yft7sUYI+4dLb9x
+8E1ZDQ3oUurM/LYxzkOgyDoCh6m/WAKLRkQZrBgmNMzIfQOHlfN9uCbCNM0imJ3
/wTvqdCLSYZn1mgv7z8+15B6+RFHjIE7bAgVCqsJBhS/GDV4DjDvRdq11fKzHxiO
PVY9D3tnFXFsV+3g8/CA0KmYihYwisMiGvRDwrqtM5s8Y8qaT83Aq3MWFK5/SJP8
904uzUA4xrXihtT6jpO6ws4wiAHNSwz12ZpSX3x9HyYoRXkgmCA2UFrjrLZQnbfj
oqUhKjnHrgoPcX4kM5SXJYjP8Rga5xu8TiqiikIxoPcyDxR++mFNJhvXGrQuNfed
ACHbzjjAd6Jph58Ksvoy7BR/ujFaEPHIF24b9EXJdgZgK/hlSdkjTFjrO6UpSmlu
1XhdT/jORiRLLth3OpLACA1kQzV5+vxqzrZz0tnL1ZrXTsA81ODXkJHvrXnKT/D/
eXFs3QeEGrAxuYmN8kLW6gEzYCHpx/P4NlQ1Nm8iA964mq+ZBFZ7SIuTqGrDTKIy
3er9bIJvmQxwqb0b14wXZvBO1GRmnY38oyArSc1ZT5tC4f5dpwc8gd/lRL0+S4RY
yADSaWtM16EG5bSGyxEQ9xzq8rnZfhtq+4e6ISXd8S7XXIMYig+OjWfhWheTF7mU
BgmpYoppphWx2QivbMRxFvJP8PRA/XheMIWoXBGZy2+onXwUWnfi3xy4znu3TqC1
9pF2uAiNaee5FbICj+S/1l8/8TH3iKPQN121A7/WXiK5XardCrEbSFjlpS07f07m
X/z3sFPA4qF338/t0/+f8pAvHEk8BvGOQwa5AvAp/XkwWl53/CQcdqfQ96qrcCZc
7NjxZVDoJFUNffP1JO8YNtvlgyTDa17T7dcLZVzsW37A9sACHCwmBcAcxKmBvark
ZcquJBzHqJLTItLXmHQYxHS4BY1QSrZNjWskQ8KbzphwbmcEOmKzyxEu+kJChggj
KFFZYJUXFKFXx3BX1nGDCdyjXpyeRoeCtyWNO3+bM50lqlXwXgFFhAvOpOJWhhEr
T3eHVL4e1tbGzIzqyTwxJXDyLCEk8zJSLjTg9RJfeSL+MrE9NRbm7kV56gCbCWgH
FkEIAKf9FxrQeIrTq0L7H9mDGFNAf/u9DOybtB+eaRUuExZdnlSP7pO2I4w4eb60
qvoOMndqB3ktMRQfwcmKou1jWcZdapXLIxNXnfO2gg9zAqca4Sg4D2D0kfplDr4J
+hAFPO/yggxiT8kVoCroiYmQsyVbmDgQnLgBdxyojk/OakqjN1wOXlophF3W1AdW
Dba0DpUlaGwjS3RgTcTW6HcLaJtXEFMI7NhDbbCBjjOC2mD9WakmRpueDANykvy1
M4tzCs1ueuzAp6FsGYJEMVyCwGftLA0ixvKhprKuz6YoFP36PVkgauMSplndLwCa
D6nuQIQngQIhPUdAVLLd5gcgbPCvxkuuUMaXvreAXLuFOpUqI+K8dAiM54v9dNUF
tNamvNcPhtc8A0Tpi+nQCHu5K3mMvTpu7X1VELXAqZRQHgz+YCxSi546bUrFAmSO
LU2cxbGZUa+qU/SQvrQQEoG0w+qu9m9PnUp1GtmcsAaa/DtCKULC50Hjs1v2EDvu
EauAJkpCgEJt8WeixcAhHFRaxO+Ctay6IiPRlgyUOt6+j6HQzmgG0gizJr7BTIbX
jfAZGHyiOUZVrsd/6GTxmCS4ACbUqPElB/1H5yeySCkgT1DHuXFci6LC9Hiw9wkT
7tsUeocQhd72lX5Mj3Cv2iuL4lj1LRagEr8yKNb8Co21Qq/UreIg00W/oEEbLVp7
ZUtoD8KtuLkylzFPT8Gqqj5jKySx23rBJd5sQ4OWoBiBaRejQ1fYZsiBeUL80klM
dEnAiDrWJoY/aAjJsM4pLUkbR/ERoHxj1AKWwTpcMDEMCq5APAECAhnvry+guQFm
GWeaD73B58Q7IkqO1GrMkHCerijEcHZis8gZaj/dSkQzIi197K47CR5RQN4LMPU6
1xJUOILi36pVHoLVr2rxZws+j3Qj90nIoGjq1s8xeucy0CyFdcNrMNS9rqwyL8XE
lDLbMl4R0GS7VdXt4IQWSQ6GNrL9gCn95vlb8OvKW/vHhzcW5Rg1d7mQ6wqxw38N
/a/G1iM+d2yO9ZQ1QMfHCD28Uu3Tu5FVH0aUCYg22exhdmv741zemTU4c8+l+0HJ
QBJU+frMYeKTpcDpmKMQ9tmboGic7iYhtuAN7uZtWbhv3VLsUOO7V1viPBkfXV3K
a9FRD7t3NGyVah4aeZUttIlvaZXS5r5lLv2mgScQsr+QPm5i6nxUJbWhxBjTRWwj
rYOHUt0+AAsQYOQnuXM2cd2/dwkXwPq+gRzquEHRC8obZk80bpb1AFb7KP1nST0G
Ta/6AEKrmaBccqMPl7zY1Os0e0vm8LTOrdNLKp3SpzJYolugLIRgg4OVvJx4z0oH
iG1sJjWzR/UMpND/FSPkSOpOm5H/leU1Co+BqK5291Hr7q4Wgkaztpm6/DqKo8Rn
NBB192oxSL4fhMJhfdnZEUVcH6fWr/2ig8tvdiHLAOms+ArZI/HtkoLAgc96MCoW
bZj2AXIkrK4V6OaXy8eoYQSpRpiH3F2uhclbBS2M8CYRND/89K4Vribl16JFmtPn
rSCp5zfTGANChSKl9m+j+PdhnXSRnmb30l6xw2qo9u7UZ+wo3Kq1FMf/Msgd4Lmj
JiN18cuzrS/YXYAX5xn34WdvnoS2W6DgIZRlmlFsIq/RXDvFxYRUr2JJpUm5e/4M
3cgzPKnfE1tB+hwu/UT9y+VLwhpB12qE8aMmuWo+MJ5ziucmraRlBwmnjDWjuYvP
iHN4c1tdLXzfK4CINtM/KM11HDvROJ93X76urjX5x0Q6IS4XylBL4MEGQq9k3tHL
lDXN24BJDXevD0Hyn6Prahizzi85tei+UHqLjvbX5PdBv39F+YE4Z5H/GxgTBrt0
Yd7vgLBQu8uJ0eyhyXyM1twLFKpgE6PpoxBWHI0xfYeCzBa7StZl15t4+xDALWbL
iNjQOCGHRKTdS/4Nfx1M5EanHpRCjikvw3zlT+f06jH996aXh+ut7dAzB3nNonmt
tzVEPf3rblqte1sRKcJkKQkJ8ngqJ6SJQjivjwEEQDjO8hXsT2WwgjU9V70vlUjl
oqkmEkqYjwFiV7aPFo/LyoiUecBReuohJbI89cJQ6NRlEd1js04iGbfpawcyIPCl
aDp6HamNkQ/L2VC2WEyOsfhRHpLFTJ/CINw/2q/GutlliivTdwgozRsxLw4G39qp
6zntz8siYt/+51fcIll+f6vDzCbJ+nhDeBehnAoISXRbZQeIN109jPgjtKo8pvbB
9UZvtlrqFH4IlBMqFbcLOFpqT13vw2zJ6VCQXsyLxf2HelVrdmvve0gXtb6MCGwG
QHElsFWx7Idn1WiOmLtVz0TyyPPTToE2+0cUKdCkkfvNCBjZqZLTgbOe1lB4ShUM
68ZEUrLL0y14q6Vv/iHKamRcPQUOhV/vPt7XsL7gtI4v7gJX6N2Hb2LEIARQyV7j
RcRiJO/0OlMV1vlO6pIQDFjDMz7bKwy0XIqSN8QUWONC3PglAOLstd/ejWjkPqvk
UUoF8otEMI9jLjlEo5LmXqniZPvNsfFXgye7PZNVWEMWL55gr0ExqALMkc3i7skJ
H0i+mDdbcImA8RyK+kGJMF6HvbQdj0J83DFfZOY+nRB5QtBwJBeouqYigrZmXMGi
Qo0AgYeuDGLD6xywNn4k18bxBBQvNxapQ2XC5dkJtXDwJRuKtpKmjBiT6uXowFer
25YgUs6LC+nWYv2SV+r3sM0KpV+EfXcNC+lO5qUwv+2b8GqSCTirCABUOcLecSDN
6LTJhcpbsY0sYl7A7LGZCCSRZ+ARDph/RkEGxzvyc8aqtK+I7MCtXXC7qvhfDvyV
a6Wijl16Bbs6pLsaavntiQ==
`protect END_PROTECTED
