`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
opEh1oSFmbJOPlazcANhkXNMX1yFLMIlayawVnfR0l1+4cAQRGSWLM8+RWkcVJ0J
2CLKNXLgMHWqC0aVmRfP5oPGtSauNM+m2yjWmm3OLSeCq5ZMfD+pXySPqy2rbEAT
wR+IlENPZpP0o2+8kX0Tq9UsUXbC4lgzu1HyscFP5SfkWUo3CmJxnv6VGUTZ3MLW
8N8xvxsUqt3uJu2pp3Ca5s31b0mfRaV8b12nA4AvVja8lzhb56tE2S0/XJeZ/h27
Jl4PZhlgOFOgckCd3dNMA4vOX0AkzYN7m8jNyhglFI/PQCY27ft9FBmJB5PHucyC
V/VZc8v7Oum1bnOvoa+1T3GQ2yt9kZOoI5rYNxGfnO9MZQpGkssLnt9ouEMRjebI
kCQTTvMnwcIVx63dfFBxWTmnNuMnB8/3T6dYfGrgmEQngZ7fbja60I5a/qS9+q0F
AUb6g6Egnudnz3QANRm7XOwgwf9eHtO8+zfTm6j5yfrRB2ymSdwPJYyqcMxdnu1C
P8kB+PwhRZYpxGNeBmCQ2N18cadMSAdRrLKZXy9bkvrbJDl+qilU4I1WW5XJGw7Q
/7LqtWhBph35VK5gKs+Hn3nMoTGlM8TKj9NQ+c0lCrqYsmxWkSMW0cLZGXg992AB
vHs+8aRxv1XFN6tUxKpYr0zbdpZSGB/hZ8+WrfKK3C15goVZq6WUMOju9r+C7W9I
Iy0lONWeC4c9tgOqkY7ILaSiI2sdp5eUjBYXJ+yjFj4pl0r67n6jbFs0TdR7iCq2
lPqyxBDQ533SfSc0QbMj3VD22LTT2AE8iMsIEdMVhe0=
`protect END_PROTECTED
