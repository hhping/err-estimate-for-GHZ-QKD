`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TzQyI1L3MTBmLuTHg2yjd6hrGySOLchyP16Q5DLaULwK7488KbuUYyhU4sVV1aFB
JvvDRBK5v8MKgRiMlPinTF5Cp1VpYjrID4yYbsco0L+esK0wvHQAYYY+wQF+cPeM
2SlHhphqsM5CRcSRF+RK3Myab2cdo2LPjseIOixvQ0FLFt6VZbXlrXBJJhEbSjvC
FebItUW1qX8MytyGnZ5V+2haAJqsA+zBs0VSQ9ijk3bAkHMSNNVjVqzsEUuBde0t
1Y42okaFU187h2XTr1Pf/WpdgHXQdKa6lrdmT11hpkHZVhQ81fSlxoVACo/3djdT
pLb1qmzLtgvxrSiKf15oBkVro1xGIa+U5OhEIOhcYIHvZENFhKsXz36e0b+7Jbou
1VkbMr2dsWBX2NyTZuE46lq53AaORajzoJ+mnrmEE6ptE++V7fB8BeRlfJTxG7OJ
gV4wLRGywfNHBIyL1EnrzcLr20dFFj8BXGTVFpiGK92WdwEfQ1IXwnL5KVkSZLCO
qQInjk4vW6Ib9NPdQqtKxvz1JXja3N586b4FXjKo1ANkmoEpErFSfRIz1J5jldH8
9sao0wnvBLWHzNvpv5ULirfVJUxUf/eenXlcO+HYsR/P3CVFRRTBVkLVXSp6ivFD
ys30rEhyWhBR/AncdtZWKn5EUjxlw5C4iAE+E/GyPDGlOg0P/AL9wT5rsuUr+L3p
azURuxDvCQ432dc8vRSvJwthSw6G7vay+JKTl4yYExVTh6A2MaPzHuSSYMqkUOpY
YC/0UtEbUVOvEmvGCoC1+m425NivqTYgAJk6eI5qwLRtRw2Q7pDHvYDct+F+pVrE
`protect END_PROTECTED
