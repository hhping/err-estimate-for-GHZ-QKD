`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NlIz0wd911uI5f27R/HPKuLiR3MV/f0BK9G3GX8b/UzvO6KSClcI2kWVbzLJ1PhZ
womEv38xmEsuBkSf9OILm9QEb+4yzKkJ4Bzk6FenxZmeMNW9Nh2t6lS5OnnK3gmF
E7zw7EtLgOilDJvQg439R9Mtgrk1sQLNTZi57q2j1BCFRoiJ23ATI+Z9oI36iGWo
vQRIgOzQrFRh/4qKA1Kfm/Nf+1FOTptgTTkdB2ZMsM37CnVLp60oSxa7EszW6nB8
0KI/iYOcm7fpHOYvLXNhO673Iv+8OBjKzPSqrBVx9eYDS1fr14DUjUU2CPoGC6gt
Me6CDSmci23Jk46/8DCqXzqLf8OhbRNNtD5bmOI8MneIA6NsaYvM6T8i6k5YouvQ
Bcq/wzFUD2jmbiaMICFqjxWSBU6X3M4l6Gh7ut/zUHJkXpnl9qALE/WVTekjefyq
KIGFQFdo0j+zHOACtSZ9NtUbsSb2zevT7bMojuTy4Eqiswrocq1wDlqeCnC3wi2n
CZSHyr9JRDOLmnByPQbOfBqc7nk5uoxWuC13XnLy4i6MyuUq5Kag4mFbyIqNg4mF
kB3uEr+g2zFj4beikKENTYk4hDcg0dyYV+5aB4jXyvAXCn1k0IpsRjNmJweQyWwH
DDWoCP4jQz5dmi1IqLfPSAV8yEGbq3vTrtITZpe1znLmv2WIFeUaxSYRrihAccGR
ohPBs4utBBUIdGxo/7JxDbWMARkdTZbTS/zHuTOaV76mZGjkwXl2PFFGt4WdCOtG
o1WguWtEzrMMle9NTq+8xAfHZvgvIUHIHMaNxPKg0BDkrk4XR4lAkkIbHRhSgkdL
V8CKHQahUR9Z4uVWMq/8q7csqU57lTvEnArLmCk1TciLTn/4kGElP/0WJ7qRx12S
6IRM20M/gMOOZyw3frr3Xo8XvS7TIoUs/tJ6KXR3ulE7D4UkBJ3HsRLcWTsDTga6
YMfNeJ7IV06Z6g3s8DnFote0zBOfq4BsfdITuwmiC4BeCezO5OSGVkQDGBgzfBWT
q3+kJr26HuNwkJiXFTb+NGWFmtBiy+uWHFcVXHsj1CImdkzyy/z1B0Tv9SmrdX3u
2vPiypyhXe2oL8b/gUGSMFTkifeuajSe8B7ikUh//peXcnyQn09oAklax+QIymAf
LqUMBUucc1iN+rmPLbiQ+4GiMW/eEBu+VkKh29Zlym53BdhbPKrpSAcjUn4QeOTr
H1WTQRqz5i+70B4OwWDpUQuUloHW1D0UD2CpdDJ+DGzxmcIGclqeTl1pnvfBlrKX
tQcLEUqRwfTb8DcfW7ixvFJRO/hsMY8X5bKtSc4JUAJJe5aKk/ii2COur5++YygC
uU6HDl1gtkLoeEDcYlAbZBjZLf/RAG2h7Zjs/G8g4Gc2f+d4LVI7yI0TnYyK4O1q
lbY5MG1D4skhxM3DDPqYnU81i6xWh9upOAKehp4KMxkdmW0jJeXKPUHUfzet9UPt
cp6nfOaK3OEdoxDxOOBcmmqhMn8MjAxIG7G4jUtwsvT84xFOIYmUzvfMUfqKgqmB
Gm4hBcQpRDgfa8FbbuhIoibantpOLvcOwhkoe0GNRJUyKssXYNdHKc/0hgyrhJEm
SrcoS9JNsM8qh+vcxqLszU6pYGpjPX2b+T0Uz0JCsFkH/UVd9NPHYql8JUkLW7mc
6McD1nCy03JOP/mZ6wzIBus2zbwoX1BX/avxEo45Z0tsUDj6/dy51KX1iCu8lEcv
1ta0xf8EiU5IFOxVRl7dmW2wEFNPLliD7E2ZLurPB30poHVao3Kqzv6j2E+owSZb
En1rvK0kX8Al5BcIqMW8iCqKEwiR3YwS5PcBOvol/zQH0pjzlRMeHbgGzrpZNmRa
3En5PJbTOtkS8gFTnSK2mq6x3VmRgRuFYEHKnUfFTXVKqkdlfkDWYpAcFN+pyM1U
Z3eXc2F6PQ3Jm22jwL/8C7rvMBxmiNeinynbqHQK7+v/YlXQTT/qQdtT1pKCkniH
o9EfTDB0wKepp8yQPRoNzncLOHQ36XcLwEPA1K9Jayy6afJ8R71vEDSK47/pToOA
61OFSuqIX6IFSm/r1V0E1YzSlbMVjklPcxyCpQorBeEAO+jOEZ0uJsNlh+NU4nu3
EJSrO40IN6uT8pGcRT6sAhbhLe/PGlzmImO7CgD2AwvS+2m9XwPoOiJZDpi06Yhh
WH0USBBSChpUSZTudIXN+7QShmjRMqfx2YJNqBVADvjZFR156Ul9bezIeK8kNs9e
PAvRZy45G9ggLF7ZUkQLUuBQnWYNiF0O2VmonFtctNaAre8c3vmLPDbmXyvvafrS
cU+nMf08dDnx6ZaYzm7ZbRzUISGzEqUD51CNCR/HGnt4p84yEASlahkN2bZQlqYL
c5z1JsVnVVuZL6jwyYaa4nYnR3HPUGm0PHLijtGBS+jIvJ0qrkr2xJUTZ3hYgS+e
C53g43JO46OhBCGTbFmjFxk7q2ViZc7R3NmnIAvSQhMdH/DxeYeqU4qmOibMP+NY
kQnh7JDS+xdREo75dgZtS6t8EqL92Ty3O6ECm5lT592SN7OJb+nXNK0XV5RchieU
+2+PEWQK/wcXXYBKoy4GhLLSxDsB9MKt4OZqrN6gBCH+lIgxTiqMJX7hcjg2CfGB
utKYt/ybbRplV2E8DTgaF/oAgECyoc0KSMPZRTpgiFQRIemhy2sMmHUqKB4vwhXF
T39kF/5OF7y8tWAHsbyJhmcR25gSrGGcKgLNVe8iURBEH5ofJa10htWI0Y0g+9aF
zVqKCfBOPcG1a2IiVhodNDXT9j+RK2TQwvILDQj5BcIqca+7p3LILaPMjfP9rgGA
2yu5BzNaI6VEbKKCc/aKEZePjSTrLF4mciJd3e1in2jri0zWUiphivLFW/Q9LfN2
JdgD+3nyPNUB49rzYqBv5EIm20YQhD6dasCxW90XRlQnQtx7qachGWBGAhZBS9A2
ot9dx0xRwXMDl1KHdSmbXn49LRE5C5BiHZBk+VLq0exLD/Gy7/UjPEAjnOnzlmV3
n/Xup5DVJ6YoL+5NdQtpqmC2k4grfiwDc2lxYr9+eRI0gIxxRcav2CjDTQvdYilg
g03WfyT6wWUddbOtvPAJEidk4PcihgbucrH/ApxRMEXgNRZDHWaXTA9mHe+iRn9y
zJNxNJTdvTnP501jNGLYn4hsFHqFNIRs5R68md7lM3oFqdqfhq/5CKL0kcmFx7Ht
jXgVZPd25XiJzJ6WwXTA94nXsLldSRIMdF/reGoxNKyoxY7QHVw4Nj09HKhIeGVl
NVt7ADN9hzAlF3W/pZBfRarjZVtw4SihaJ96MzTGPt27V9Spn24Q0F4Vv6ffI+dl
6A1dKAeV9r8g6TKXNwSxHU52kwYmc7HtAxth0/4vmYaGqBLd+sms6bZ3jF3IDsbC
jwqJAeVVBBSoLJAY1uZgsQL0e3OQ0rwvFlkWX7sKCHo2LoCzAfGG7OYH+xjAPEPZ
WrZwqnEZ3p8GglyuQwXDvZzXZ1qnM5bON7i8R1vrtFO564ZWrrbTmM6cQxzi6HNt
EzfFLmUnLO6/v17NIPEnXs5ssclfKs290lqzehzV8FrxpXDyDEx2j9deBxbT5T1X
BW4Qb+TW62E/dJNWut+0OtKQRZrVEGB9t2I5UEEYqNe8/OIkfMHaStPKa88gVqKo
W5sDQk57M2/XwE/EccI/t+PaZU6VL0FRS5j1WgjyhB0Bl0W+nw+L6ieeqCNLvR79
RyBd6Iiuv6lIvykk9R/mqTkbgmpIhHLRtsKVUtH2wWGMyeF7ycbFWJo7hVwBWd2H
I+LHAVJcRMZ/H4wTLC55PzQ+14RO0BhowOovIGt7sZGPNU2FxE9w+vpYCxd4fq23
kbFgMSoxQaikdsP6CFI1FoYCWkIRxqsX349qRj9cziBNzs2aQW4FUd0Wyr59AL1G
Xe1UgNM/62jU8Q8EmMldlwPigkQj3gt5Nib5VyjziJog01ns7j4/houoEJj1hy0R
R1i9s1vHti6Xw2b1p7aF8iBrkWUrCEzatfEyH4/NXUI9J+eJzNTSpow7Tvr4rOtc
RArzbXPqvERE0LDSvPoMuZrOmZOxx/mgxI6veWiSxLfp+jR4I6d2A5CNBPAsh3zW
Lr0Mh12d8Q41zKMF9ahqiXcxHM25UDr1ppJU2P4XFo4xOfZbl6UC5b5nSPHDFmUX
wHII3PWjrwteo8LbXR2XLM06iNI6lZ7jOhl7TC/6yiptw7YBDPlAYVabEk5wBxUC
HzVmDr6VaQUZbS8EocDy7MdyJbEBy6CW0zSqMMjB5eg6D06sV2HBW+GQgtDvtto4
VOxll0nvDVH5VqA6NFO33nmmLDAG2srYaasUF+eAhmbox+W51457VLU3Z/ai2Jf/
AW1LF1wXFa2vlYS/RunuW+ad5iqPwrLPW1GI6wzSfCu1nISyXX5dIJExJLJAfJE7
22ZYGr1TWIVp9vPv6CsyNC23Napwovzu+pwJs7QpwTY6qU5DErph84Uo3bPAkwsO
fObK+gU8ozwy2nKued8D/e22ufoK7Q3+ON8mUpLaryALK5tRAQiCQEOyveFFyJRH
8dL7zp+WIDAItmXWRxQY7PhlXRJYOYXnYhRndopgV3qOvN7GES4Hb7Mlek7KexkQ
uvWaSkzGKIUbTUKkGw3K8wHDPqlIg+/hxw/XPMhhbBcOJq7b1ijjIjsMoyDxkUQa
5I7zsih2YWnzxhRzTJNz3MEFgY8gVUwQ4H5wTSHgWFSerhBElqWcg0Izho1kBhxz
OBn+FlbNPEtR38rD/J0KwyNgSGVuBKqX5ik6Cx9/UEbtcQlcmXJ9WS15RhqW1JPK
yU1PmJaYWqZVxhP9K5qqoxbaetoYxIfjTpBfiTH3EDOWmnTOl9OCwCYCXGr1WFeo
4WwdgaQixbBMGEl+38U+EgYr8UFrLtR+hk+HMOy1lXipaKAY8fSVojH85mSZkHQX
mo6bdALeHLGMRKD2tdZtvJ9VUaSoFGMQ00yV8M7acUuqRJUrVlh5+WqkIGiMiNpn
Q3tj3tgEkGEURZao2k2L61LpRdbvyB5lxu6eZ4EOkKPci9/j0GVK80p9UWTbJsQ+
6GpMB2YAcz4fwmRSOZF4e71efckiZYJE4IvSS76o733tmp/qmfM9zURBQ+ItYX7X
pUEABFPSNTGGhbb4yLGmTJHAQNDkLuXM61Sh6T020H4biOArsTcQEkMkbqJFur0z
7zn/PDUeb2zKYm/t0KOdkRhC8LNvO2briHZBAPTzLv4uVEjFlMd0GI7ZfTdRx+pG
3jKepixXXocKZ34rsvWaOrkannhN/ngTaPfhUKiglLWmIUWlUc8I8Lh2bGt/LGyA
a86rQIrlvsb0DCdzKJRKUvBQSIAHKi3VqouFYxzHFnbrQHdBEwjB/8mh6gn1D9x+
l1/ywoiD7SkHfNrmIW8A+NfDkUKG1oHpAzYC5gApQdDkGGYYz8BKtUTtu6CTQsRe
ZEzuYYR/ERHGacb29GEQZKUQxAfg4w0BdXYHTl2j6uspVkFWog3nw0Zbct5s+0qE
Ukh4eAazlkxnSaH8wVJxMZBH7cA+GEP7+lA68mk6uqL/e/ZvNtGmn1Yab8GQ2DSf
yTNszz2d1sc99MrlikCzXzWhb+W9adtVejZt+sOxGqfl7iEAzePVdJkKqd1/oZdZ
ILw9sm3/ZHuDHhwce1rVGBkbcjQPagyvqPdZNueFcJKItM35cHtB6dyT29er3kuh
PDQ/VddNJdesf0N5n5Z79HNGFGmt6U8KT5rJWy9bimO4dzvohp5E3hVaqFM6cm4C
sAoaKgSVyD2YKM7t+eLeMonPP1p7u+hyA3QBdYT8TvV+KPUh69XMrUQFycaj2+ED
9Ena6k/ZuUnTpHuVeXcwMjx8oJr9K29dYMyBcNaXbNVk7gLOHIcZ0Co7nndPwBHh
r6D0+9NgAow34TFpKmhOoJwiwLnnip7Gb2w+lZKO6IEaItD6gfwuEt1EPuB9xDCE
ABG+3ru8jyrUfcMxVT09q3FnF+0FzcZxDjO54O+7kIPffld1/8aH7wbI0N4E0OA6
NQcdob8MvadgIITZHPweiEwMUIMWsnjf6gkm7WCoJZd0oTjcU7/TNo+37ExKpz4K
lkC9hV2/ErXAWwCZp0Vapqg1M9NIu4ne8aftV4gsvPKEbV7AZIul69wwyl4E56lT
PvFFceYc/nhql2w1Y3CDpMsPQP9m8m5iN8z63Xbl/VB6Cx5pO8faJBinncEAco6A
aT2Jp3Y9WtpCSp+RfrpMD5LzL7jgS8e/Fa4KXUV6HA6xrkOZGeE/Yeb5EAUDLkkh
LKIOX4/BZKmE4VhPhTAg0gDzQo9Qs0QmCFhgRYYO4Z7GclD9N89C7GED5QF0CudJ
7MJb+yKZNB2lpmBLl/7ev5xJsYYBdNYrYOhXqYmIBWHVEzl6JfXFMTUwtCRqagMu
oGtQFSVPPMMoVmAh7s52LGRbJd7khXPEDEwAUpDErvOm5uUB8z+D4WzoXzuHq3JR
ldXOkYb0EY+Y9XNsdFs+QnbeFyQ31u2QnzIM9Shr2Tt1jk/GliJOu4SC+BKfCYyY
NxrvdHZCcSTth3UPjSQ6QGbuuOm+VGoeqytiM+ZOhPsnHKN6KE9WBfu7OVD0rBGt
j+b8G9Y9wSeWP2XqwncQOE3+mAbyFsrDc14zcw75qbieQywzJD0W4pSQoIty6NF6
o268OO/OspipciH1H8RbqDKdujAx61TRyDWSTyaGRmZmpAIODQXT/3uvB865hbIM
rZd2RmUj5UjI3T7KH51sBJw7/+Fj9J+42NVEpOBHbaoJu6/RCWvUQvY6EwL49oP5
rJkiRi1Gl0pUdEjHlTU5VGZwfYbxDJD65qSHw9Us2Tvdv/bxElvoM0yaQW4SUKAd
2Lt3tFbd9/eRJ6yHwoqHaAcXT0vAwRUTEa2zU7bLjlB+h/t9sJhPzDeMTSjtusJE
Cjq1PulLLvWUR0Fu1X9SL1U4XDmPOxkg5bLatSteI3HqymH1NIylnVjdek7VHf/y
XQ3Ys73e+dUGez05YMM8pYr8PejBPMARNhnkMJyT3c8p8semukua33YW8UY4rz1g
yg1aoeXdN9mm3dBz7vVXsScnXNalF4ZO4CU9wlWrTd3FW3k9Q2vVwc8RPnTMaybU
iuHBZtcptAx3q/4SwZa7DQRk2TCWPjwubC2sY9Jw9J8H7im7FrwC+XKAtGlnvs0Y
POAMQcjnwMJnJ+NQADkIFz6vfIyyi0NLRhuHysdcX3ujzJRo70TpuyBjlbeYWc2s
gRPFvVs4s1JmVpcMyUZc+3aSXC5faUMcoYb2Ev3LAnqLq8xUvaIrHdsdOiNHU8AH
JY8c83q8YEh7lz0N771cAMhELkKYbLBRPuIcqEqs4y5D0Izk4fr40ZTZ5cp9KDkQ
eBLdIMnka8N4L4D7LJfvxqxieY7DGkx8uaR41j5CWTWeCoigeyVTgy9BsjMk355x
uuDE2QDXsDmYELaYXmEvwxMRvn4a+o29CGFFtbvctkD/KGT1tBTvNw+GDkTlRSYH
z+ml6YX/WAxcuSh+U4iwvjDeUnEY2YBWHHNzfVzkLuTRNNrmqWr6oyH+qfsmOhMR
b233qJT1hjDxrt9xyYyf+RqQQIfwYd3vzA3lHZMf+bg4NSxIaS3vHPeViAHisMZP
4bQ/daOG5KollHD0CFVmATvxTh0jO6qse1TYMhgW5jxoJcBZKunfIEoFX0+TDQvK
D15D1//SCowa278my8epsLJtAnYh2Jy8nG1hrktrTh8I1iI/pabpp/Aohzit+YUv
J/KyMrwvLVB/6zbekRCnjLvOG40Kog45NsPeJp1ActP7QKLAZm61RMj2LibDoX5A
mXBGDdETX+M/CKC9vrJ95Hp3OErI7ED4Luz6Eh5zUKhJu0p3WQgke2759W/8qg0X
9PqGeVsOJAv7AFwTc6Np4J7AKAMxH53n+fphw2k2+rZojKunwYFTzOrdEqa20XLT
TWneJ2+iIyRXUwfQx3/NZY0gXHCh3HoVqwDRX+GXGEE0BUDO9PxJfZJa9oydwoeb
JvrOuZhEqCiSkSOXmspbgqp/56TY93eM3qlJgvu8MBy3Lbl4I1dNX/iFR2i/7ErZ
INKmOhnlo6C3Mf5uxrQs5S031Ckxjz3b82ZNWZXA68vAWPWNte5HB37qJXXTIiv9
XwN1S+I1ZFguWvEGSwOwf05EISYALvHAVHe4vIO0wFHY3t1hcnOMo7DJK1elIwsW
Kbz9SM9G6rV2+ghRK4HlIIG05CEKQEHWQvaeOyBtyZfLN87ez91NbtFg2GWe4zs0
FAHOCIw3nczTEGifKg5mVvamRaaM0YkHBctxok3MehPnl806nDU4hltlSC/ARYH/
cMEAIZj7u7gH9xGDWl7CYGZLMUSaHDuRQOSNelwYKguQEVRMK1IQT57Km5kH38bc
cMR6TGyACVPSussl2UF0QHNgFDenv/c/QPK4hlYvcfQ33O28M24uPCYLEf3PS32x
m/7kN8MCNB2G3hdDgd21Ym7XPNLRrwaAGQiwbsiFWhVZxa1QdRFqUuXrrRvSf0OI
huaWi4Wa0gjpb8G8+61mL1eEm97TxvykrnOeRrItjmQ93jfKrzxBwFKlrBGRyq/n
+2XilqwraKzKRfx439XPajuEk9+LPBoTUtz5a372lT9soljsHesd68E+mSuJqlYn
gbONQ/84OZ3D8pjyDDQ/tkdJTA1WTxhYmrRJ6/G1X/UrEqtwbJMb2Bvci6cKPvtN
WwUKJ0r11H5+wXr8z3/U0EjsD7pE+JeKkbVe9F5GeRSYzSUVFApf+W/XdbaCjF52
c2AqsdeoAqNBOgy6ZQrS3Yzua3K/gLe3zddBbZVqgzG4u1jVxx77S+U1z/58Tkvg
ukqtK+o6uQ8EgUpm1mT1jz4DpSa8GrGr5gF5DaN8X9g3eqScQhA2PEuG8g35glWP
5rYGv5UhhKCgjH882aaNiT1RooFYoy1ZaTZ7oZIb+jFLAm8dlIAlCW/CawBlt2Z1
a3+qdFJAC9U3Um65g8RAA5mWr4aCHVXNf9HOiFxavOTZf27v5HQZlLjYPMPM50iD
CFG3FbV04oXG4Ix8LfaFr4rtOMyf2U5sbyTyA0YQSxuzEPG8+ihXzFrn60mCGgm9
yJYkZmk6lI9rlcUakRm8ItJf6/XifArOD+SqyEEsOLKPB9VYG0IT74sl5lLZ+1Pa
WpfHlXh9GUa75aLifrwW6a7IxmxKjTJmW7iixwFiXiCX0DEhBRejPEuSdzemyfSH
/1qvSUff4q+JtUs2Q3wHNf0qA/C0M+S9CWUILlk1eWLL0zxK0rRndoWCNUVDu6kB
OXSuhYMN1XIrNVTVrTy4UvhiPj9+bWu5hhiFQbrHAOdi4sROv7ckuIgCGVKJQnlF
31zvKzLO9TB92o3BIOHMVxNL8iqAMz60TIzbzuLnHOvznEn9rg3pnHfVHqjlXWZ6
p0XzuOLTMSmf9IZf0u7jUR6Hl3sYimHXohVzleNvfWsGGZ35oOcA+w6LwYFyM/fs
0++QJ9JLgVis9H9DC4HfLarJXqegfL1qvUYF0yJsyuzIEGnDJSpOemmvwnJzz7O6
8fnLrA6TxGyDxJFPmTGMMxCFMQpDjqwyFrIFoNN8gSnBXH64w6ZQoMkSNpRXhOIc
Vp5DnRLu9w516DQqe2JybitqgV/eDaUER8TrSHk792ogbRlZkqlekru5b1uMl/nN
ZP7qn29MnAjrtC6oz7i8tAlBxDHZSan6rrxZvPnHarowf5IIiyUn2lpXui1g5sRj
KSWdwHeDqI13saD0y4rErj+BylANEX8zA77yYKR6YNnXGGBV+OffX7E307Uick4D
gVszLgLzswRue79yJgvCEMi1Yn2nAR0RvvuTf83zizmO7MufGhPu2Q+4eDcE7USN
8y+hL6uSwp5WB9MSsPc/UVZytf8eTraSL5gqyK5kNEmqmSQBE3v7DIDsMq2j0QZC
W1z/2+NC1GFxuYZRyqvdUUKMYx2DgXT3OLVQuNlfnDtXD0r609eZ99ahIEnPPFiR
lT1nM+TO6hRcoYIdoAtD/8Kh5GD8W8L+ZnUCihh8c2NwIsm0V46FWqxsn/fR9hbH
N63zngG8hhvCKlfBJJThO8oIZ5jAZwtXoHYhL2cWvYi+3amUMv41/2eTTGmfuExr
vAw9H9Ng2B2y7Cy20XI6PrYMA2GwGM6a11LPrESlYSlJ4G63097HN1Ezq+TsmG3Y
YepwHaWdlriCH48tn5Dmio7a95Is2fnq4frgYJsrxQUcVaSRWeGXj2oU0X265R6n
jOuNUXG+Mjn8CoTo4dfyAUKwF7aNDRWAn0nFIbnSlz5MZ4Xw9RjUveGRD4nh3p5l
Vp/b/8WeSJS08YCGzHxgSlzuaXp7czC/9Q1jfwtVuOGqMwsnM81HPHcQDjetaURd
nHENdABnPhgHe0yl5mHYxVWOFMF3EYzE+jZNcm2R7J4CmbWhzCPkl9Su+Tm7/xzQ
6r+4LIr28guZCoI3O3GB3YcK60kpMQ++BnK1ZU51BtcGuOsMV0Mqdy4YWZXFFOhc
VUxzbViuX68Kn19Bv9C8hpz2dLH/h4j9oZWjPcWG0ZvURdjqHZ9CKwx1IDDIHOQe
6JmMmnn8h6VZo1IHuocmoS87EAZz5YlE8X3+VWVkKK7Mx3BQUrODXzdq++cExkL9
RqF/42guKLdiQfkuBh8w7d79k3K4iAdNJlI1PmlnwzkPl1XUiYmTsm7JRCDOGmW5
98A5vU5KpIgWS3lPfXERny5vfPGFGs3WKLJmVhg6ZDURoZWGD/w/qhh2TH/1GTzj
A3tmxJBhPRbjDKhFQHefQcqYGk4dEGVv0XWt6zCtu6HxeL5KEJnnNiUTtsVgHsrZ
O2ezeriLk8j4EI3WE+ob6oIU6D29/9ZsOV9Tj+3++npz6dCpL9cj07CHm10Ym389
85h3+u34fUBAathB6TWPabrJTYs3Bclr4qOhujnkLvV6La3ZszksWeSSOR8ov4PU
JlVtPS5Tp2RPSnlBrmV5asCBwzsO2+lmUO+c3H54pG6HKU7BixmjBaUjzsSpAhYr
TnMRSgZO/zmhr+srQUwtfEBl4EEYEtkSw+el/PIDmuNba9IbER2wu98uzMexVCNO
X9p3jiYG0RE8zbhENt+5KkGuE+pZ71XVu0hxPO6GltjRQewetUnaHMl4vGnGcZ01
9NEuzhCvBM6X0vyzlPNcsz6uF1Ut+xssAoNsGp9rqMdVXXW1ZlRA1eSBIDfYWldr
OQr9jOpSrI/Gjs/3BO2QE5ZzGmiF3QT4H60aUI5BKa2NQ7xmIqOgQWz8yb22+eEC
1IYMKPo0OlzT+bB9ADrKl0UGJTB7qAnglU/HfswCXFiSsAn5tuaLZ0lBJHrp734u
BPfTCm11R7JDGvXBJRRnQr6jIMG++3YmoBk0UNXzp/8n2FcA6/U69dXsaklOmczW
4SDOQ9sHvn9dBsWRm+Z54NS8O/X/jVsUQZq3qDxPDNJ9v7IWFL80fNCm27EEhsRz
ICWuCBYP43JFnFsK5X0F2moi9fqLL8EOj9CmDyyd+7HNoNJvsCEGOqvt7owjWMLQ
GaPXJIWtBpUZYZ7gHU8dgnH43FBhV0eVac2b2pd0AF9S6X0SoJg6maiwfJcY3rRl
jyulI7fu6z0V56eJ5YKCeO/zr/Skp8/m1d3NZeazTDzmJjbIlwbATGquoecTDIqE
WYMKSV5mU2IIsL+AsV7b+tE2I2AdDCQAIi86RzHNMaisc0FkbG3KvJK/6MZjBV/Y
798LdoIOC8Y81fdVKfLo2qkSpjDmqbyU1XarrLf+EKxbgmkA3tgdNfazPS+/SUvF
+x9lYm3Dlq+otT9zn4+waBCPIKzV9awt6opnFRdHWGVPZX65X5ld4te1Lppokd5A
X9PUNnW2V4/6h1lv25WrSQFlcjymSPB2VqwxSrg1EI065nMWWu/1OwkeMycD9Vuq
VDR6RoEulKsDUhhml46OXWaHg2KTnYOB+rcDUAvfLK9Baqmml6EJao0bBOZvMZjU
Efp0j4d+/6tre8Now4S5N3mLg3ybOXrA0ksNX7TS3Dnypglg6RO1oR+BsZxsB2tS
f1uWNifIiknwW6s4/CidDcvfEKpTKgISEg3r8PlkOjyKLyoWZRinai8GshgAkpMM
Wi6OEryJ4upbGyD32JS9Odntlfn90NeCaOJ7d03SoHnHe5BuixYSIPxWg9/+ovTk
wf8JKkgQ603OY4pw/gp8nvGjgnU5MqXapCui5HhnfIu1pj70F7XSSULFervWLLAc
xPsOV01fW3DHJJ/fFkdmvzXEGNxJrublL24IbOe5QpcGrZiJMkALCL2lEqqxDSHI
meKk2aBpWXZQ7kGXU/xgrJf3tpgbloueqnqFGZQo6UIWAa/6u5f/Z+RdT1s2T+bG
a5/4UMjvaHPk4gzETsBExOUxsVcJw6ezb5wNlVXNBfvZE6yf3DsFjD0zBPpbyaYB
C0PlcmZgiH3bREcuVHffcCEF6N4bA3Bw6JRLCqAkDUFa6YCoU7vuu0MSQZ6vOY3B
s1ciwH1Gs6Dq6JaspoHGOT8EVouKmY4sMr2tiTA8l+HAeXIzTup+6fwsMSBL9100
AtU0psc4WdFhYWCLhhZCU4ADb3TsdG47PU4Imn1SHkZs8ZILyt/dnWi91QkDtG5G
`protect END_PROTECTED
