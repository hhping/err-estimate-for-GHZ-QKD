`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C00Kn+PLByXxa6AVsxwGkDJA4aU7MrDQkzsy2BhoA011xcOh5PaHkDgRyE/3jyts
EtfseHsq74QMzpKhUIE2OljEoCmSOa4VkRfWj4hZGoZX5MBa/4MaOkRkR33b6DQr
4c4ptyZHv3mSPMJxfjcPbMrmGPqrgOTkoOjRkGic92rO6MMv7hP9CCEG4ataeYXw
buHSULJU6HHyeaeZZtO3HRUBjJa8qfxFMKzHAQnsa5m+CctNanD5y1J9KuxJVCbk
wm7mPiRFHPIK2v9b+ect4NWTXRnE0tGgLubF5PnYPJ+Q/Ka1CwhkRBfXEUfqVWB4
Qbu7uLGxPA/Ed+twZLD9vk/8g6fX2tmzF4R7wQqI6QelJtc/7G5saWJ5DT1UJCsg
uBIivDJ28qLaecNNB/9jVAGrQq2G1UnZf5oS9bfsNP4rQeBwCoS9M3lqhKvApidF
JvGln+UFyyE2CVY9Mm3LD6ruZlUwjKAbY+Pqk1ru38FP94yfu4o4eiP8qZSLl/j6
DZxK41D4IhsdbdHpQho6H+eIGW1knTzXb3tcuHA9oKGS431SJySwStEnttHRWog+
wrX8/jQqb75yeFytuBuT12NoKL/z1ID/e0IZhswejs1qfysx6GgxjPjCpAr1skzN
n0eVSgaAWXQwGrfxrwNbnlmoxTMSJ+3cYoOoru7BoqBYxfAzqA0Zd5IgbG9lWE1N
ixCndoCbB3/MEZsO+drQAoTIjnsPILiY/HSUWM2VT6M=
`protect END_PROTECTED
