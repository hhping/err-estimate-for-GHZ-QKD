`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FlFOzjxV7ltoy52X+c4uJj21WPpUq/BpAXAeCzfZAWSpJBwLokcKUfD+tIEOZ1KT
ABPKLGbIqyQ0WI9qdlfl6TYeEQLK/chJOCze34xNXLYhHgJU/zrE7P+ESt9SYP9O
ggjY18lIPZZuLB9dZMTdSMY4/8LhjyoMOM04hW3LbRYlUjN388DGJkutzJqGmNq1
r9S4eOtxml2SvZwlaGeUbncIOYG5gvyc3Y/kTH5pv/YqFCr5gqylJm2r6ByUPuxw
vdCa0sJxnvBkM8ytkhn4IwpKdwDpa19otuqlm5I/YjrQxx5fOXlgvgoVOsoQiW86
/h4CLF+t0y8g8Jq96w+UfiNSy673OxmWm9MW+vhVq5UcJmVWKMgISOFqJEl18Zwd
bSyBBXed17h3iBWZVN4CGJYy5UdQRb4xkBdrSSb+nyYmcWd/u1J8gDRm7NTKv18d
JqwhZZHAnpSXdOj8UE5ESPkQ7lITFAH5BnoFm6zxnvXusSqnfj2OCymLUbg34U3i
ZpuP7At/K+Y+C6i1rV0nVUFDjnV6t7CUAPXjVBdlrlgWwKuFjXrkKKmXqjgiM/LX
FOpbCfzYNn5+FhOuhbN6Qn/9lG7W9OW0mOCGPPjzRAWZ9WBxdJeVQWAAuY2Xkylm
dudbThq3qpC67EMbFaTH7Na52lZMET7TjM08yk2TAC7F/xPh8dOdvFZHWmbZkyoc
nLVYDmu4nFOwjiIxZOPMGbgVzLa+Hxxw7d9atXHah+mswYE10dMPOTyidHv0FBTG
UsGUhGqAEpXu5w7654XC1XxNb4ShgHsGXoSj7gZkcIEf8pyuOtaQCqxEuZg+BiM6
tcjl5PpzBbCmMLBh2POA6SRj4KHxub+gdTsOn85TDD9kPCxeyAlhXwqVW3Xaj10o
`protect END_PROTECTED
