`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6f5X4KUtWd5yomy2lrGIUbq0mOJMByK8WRjIGZJgWmY1AC/nkv/91zh4B3bDO/XV
xHNYxiu8YgXNQ4Xfpq9dw6t8s784VKc+xamEUcpmIn9Q+lzOcmIp1clqAEpiC6Z4
1mKIVHMMX3G+fSoPZmxau0R6HmI93sOfLcGmyy+o3xhrSA7DtJhnc5BQmEht84QJ
xezIaF+njCJ0/CCF9fSqWlJflbpfkB8ZfJ8fY4qFNnA47DBLvSQ/lXLzlrykZF2P
80cXm3LjGlY2m3pZ6Rd8MBdeQd+dT456xaK9hFhXWqoI9LgsTO6txx3gqwi6aImX
pFomKpgVYWUU+QEe4N1P8xw0fvyKYevMrKL1LhIh25rXr3XGEP7vjttE4Qblj7WN
Brcj/xZyYImVrv5d1fu56P9w13o4+552LtpKwDst07kFpilx7c9r0vqF067n9luI
iEtWbEsYFgg/lJKDqlN3NUIgXbrWBvWsKt254yxtacKbxCitD7j4zIBnQhpUpyv+
m/bYfoK6/T85HAKwGBqi95+O8UFEHP63cOT9Ve5W0gT2+sbYxk36DrObZarque+V
amb9T19tajI972QVOHEs1ytNsCEypb9D/OBrVzRNCjomN95n4AtMIGPoD3ouQXzj
QBqBS0LthvCqOYUtDqfDQkKnw6He5CNRWGLIuIXx5VBBzlGMRvlCLPvIplwWR00G
qOHw31ZF+klC4u4z8NwW42vH1bwRanwbnqAJaNXItdc6R+aUUMEo5cq9xyRKbfpo
VFZTSF9wMCpyx+WMkXC4Q2M6t8f5xy3B430C1ndsLYNtf6mLpIwWbntmeP51/XTA
Bl7Xw2WjyRWZrSGXMe/ikGh5mGmyGSP1681P9CTcmU4WlrYfQKewmTk0F0SzIHif
mzn39mDqFqL4m3aqz0CwGs8WSUkBJiD/FydAEHRan9OPrpZJL0cl0mV/ZlAwqaiU
IoqVUduPWPEhm2PCsd1CdyGPqGFBn1YMMCdl4ErSJmJxjdgBjt62yKCcEr/Y1xfk
mlo+9mq/0C+Lrnfuz7HuUyVpy9J/tywqEz7YyMORVz4YImz9ZKzJE7FDSs0UsdaG
UjtQ1sqZtlQknEIgbWGfiEOriHQRJYGpiynbk9cnoh8/C/Ru5grn4VAabbbtdjpI
eK7xvJjIO8je4haCHJe49nlxN+/7rSOWMRmTEs9TvEeGyaF2T8VqqaKxSeaGapOG
goDUYZ45PbjzyUKVKSC5kRMNlSplt7EFL5uEnofu0WnuJZdQtDNewTHmuXA5xk6d
0/ZDRImH4Zj+os+gdZSaRGfQ55zetSu27fAd2Aum5aYISzRNbyamcTWDtSMJA3Cs
gUCvqf05g3pweMrM/NF7Gc+fE7GyhpjOwJOghZFzskZYXs9HeOFVTlpUx2k2lGhq
Lvy+X0w1bLufBG5enxc1JXznDykpPjcdr1O4NxCoz2VqmFSPhGzRGypddzz0F1n0
0skoo2kz8sa30kX+zZR1DysgjlGyo/B+HyIun+sWo5M9kmzMf5VBjuezskp0Qwfh
nu71E9fzTS1P5TRhwzzfS/ZJXLCsM7zLPI9ZMqnsfErou/1KgmIgrko2gjAIl1jR
ZXzUy3VM8toaWM6r2zo49h43mzrK8gvlm514Iwg+ldEiLVbYIk3xHcgRAmJAKkBN
a4G5drFhB4rmKfjB+zsfgS6V6B4g6GSKAWpPqjIZNYgkEHye82FtscwZwOhjx1mU
7/BBeYr14V60EF/i0+qtHqg3n6bUoRH+EN9N+LneXTA4Vfjr0AJAxF7uduSAsH+h
wQBqp4E3Hz/+gM0em3MlhyOkfKByofiiY9A66108mK8QLRp5QBH/dLecDEZunnGY
zLZgnMocnO26Q3l2I20IMhtrpc65HZfiC8lr1wVISJ6ZZgNT3dqV/GAcPb6DchzY
mhJKUhsgfYd2iVAAIOEu5mTZZkauRJlS4STe8mZgkHwbELAB2AwzEYMT+YMqjd6H
oxfm4u9tz6D8Xr4vZn0UDlI6R4wTbcBwxgmok8vmuA2O++TY37I7V3NgG2TWAakD
1Y/psHavPEztW4Ano+5GhdOailHf9FhlhVHiKuL78sIk4ZNbq5/GRH1+Q7MMTXIf
tf2JIgWKxPafuAvr5HY08wNfk+Ttju4Ec9qnOOnF7HctxqwA+HoyqT2aX6AMkfc3
JzWJzaRLdko8aCMgccwlloPi6T4c2I0o7i9IG+7zhRJZm0LH4FJ6ynEJpKKZeMLs
cPD5Y+2Ckx1lapR0mv+zkOQaDMpo/tfXSmCHxj3WH4nkOaUVgR834/0Q12y4JTr7
kshkWlUsWxYH86AuaRisrELu9EUDos858D1aTxualmsGF0oRaFQz3+oMpjvYIgv/
dCJD0jhyffhFx438Fm3enzop5oK2lop1qExxC1Ctz0p8nbambYZDZSq/Ik7vBcK2
IJdhLc6SWQINY73nDntT/r+8HWS2ZCxpS8cbbmUhTjAROjR2NiflFE6mqghRUH30
ECwA0oUE4QpHdKIjWcrKkbInlzk44HtO2z6FTuHPY1uAcGOmWAiqtKFsn699pLeH
N9dpos+zPpIkQe91JzGwX4daLhWpdPZifT/mF9nWCKBbV6EMGm2Ft9yAvnuoM0Gz
ajOQTw1vVMSfvi2rqeOWL5dl8q3cnN4qHIgvGh1KrKATJGOf6BvT3QR97mieO6jL
J6tDvFJYADyhaHlgu9hbAfxtbMeR6GiDgciq1pi9eonu0w24jGuP2LyD6fI1s51/
59wejZ1gLD5E81FB85oGbm64tUW+uUZ38HXaZUCk3vMJ8FpnhrMlPaOmHriTOTpX
pVBvDNG2WxfChy8Pb+jccnbhfS3plYVqE6fE2ZZq5h9sGM6MwJhKeLq8A8cYRFr4
jARv4bo8DkGx569VHx3YRHNGpu59ehVVDidHaNg1xQEhDJwS6psPtMDNUpcHQUQC
wYw+bGbDSqgbNBTwBgl9Oh4wxvcSBR5A/1K9jsdJsbLhYjmyeqkQYcb9sArOoHNt
QFWEDRqkwA5J1tYk1i8kbZr2uC8p/HtJjNuZqbBjqE8Fjor+Uw/g5UyE5BhBOXCm
NUBTIlRuHh1L5d5oV4lXtaybhYDLRclZgqmPCe9Iv5cFoamCx06C4u1HXXdoANCO
`protect END_PROTECTED
