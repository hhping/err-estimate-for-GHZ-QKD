`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7l+iZquGV2Y9rIG2VAz96neFQc0HGfax+Sh4X1pZvSkCb4PRPXqzwSbTPkBF4T+d
kGI3T0YkWUD/H54NLslqeW0xBmibi8AQnsQ44PJmzTG7dEFjwjxBce/BS5ilaOHg
jjbNs7TQMZi9vzoyG2QwLN/0DJBxAQLb6CX0wDowDcZrLiQXpurZSdx9NpbFqhq4
ET/NX4Hnrkl+F9TBaBeeKdDXm+pDnO+dBvcK3ZsLYezVLGrowWTuI0uMr9oXOmaB
m16UWPm5jBWoTKoMgVaRyEv/q3Pbsgo+sx/UDkHV+HLNIXs9NLu+TXDg9zszh8wE
Q/qZZP7tNFDIpCTJSzdHt+1KfL/M1o7W2qu6I4I+ZZnJDn65arV2xcaXo32XBieC
xfrswPCpQN+1I8lnuznv5mRfnhD1O/VBvB06i6D6+B32AbSry+CDerpnzTONjY20
PjpGsFQ6xI9x8khfY9TivBczH3ZW4MeS6H6ZIcm45pkzOISed4clnYhoZY6vCLg6
sm6VrAZEzWUESo5XPrq0fbh1kNf9ld8xd4fqowN23p8fgxIUJYyZ6aWAEFTwDFwR
OygzkJ7M/W6mumJupU+zNbxuH1FHwjgYb8inw0wV+GKc3kf6W2RFfkp0+lWj+SFa
xVL2bgNkI5MwGzN9lAtw45GYp/teG/EcycyOtebv4iaaKG4d5IMCZiyvLx5NCU/y
N0JZbXPN01jcjYh6+RzJqu2wDgLUqdjkW4nDw8/2Ddx+EJH0lvf9VjnX9f+AsxeO
mw8bZBIm4pMsC56uF9UQhH8qsi11HfrdG0KGzkCiIPwGe2YvPCfMAlyXRLTG+m8S
jLIpLxWqhq1tBSLNerUjGHwkNCN41nxoNW4OMvJHC18=
`protect END_PROTECTED
