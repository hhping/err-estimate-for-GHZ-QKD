`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GdmWlvmf9QoAjd4JBvi+jk6aDqDNInTK0U/4qJBVqANzDYcFBRkr46M+pjNd4SON
REG6gaRHLZ38mWKvc8FDgTis/2utZKsDcmHnNPrewDt76s3SOOk5nkF8hEOuX656
gw6z5YwPtPj9VsvCYVdYzzpuO9vsMb0PQQQyDY6hlnUboTKQcrSbCcmP1NR2Kjv+
pdpHAiFV/L1CElrQxMWs1TvtVKbmBVOu8KtGKS82AfawoZHSD2wilGCJXzUzJgVA
/Q2qmfygDT7NKUhUg8/xsQeJAclaJKgTO9EBIo3PxbICfgeK12LjRfgTgLj4QT3m
DKxqpZW6kRSBMKrYiyC9TTBYN6Mc+2Es25E7aNnG1s9ZxOZikYotL0x7Ph8g6zeI
eqOzt2T5FicaQhJ3nsTdmxU/dWMxc0IWrLJ7p9E0tL4TmDBdMH3mPsRr673Wvt+Y
m+NmdqrrMEFo+LVS16fLSuIWuSROb5/bP0ePyS9ORqhoDFOnj6b7UJx6KnamOIKz
Sbm+UFf18aJgONqTvhpMPsJVpaMM1q46yF6gpmRVfwpckooS/xahUPu01ZiFKn13
+6LdruRTnleHZOLH0F5lVeP71nmTAkRl10rdBMnDB1mwpOfHe0I3shvDuLOudJhU
m0hQbu87gdRn+iWWdvqDVAaX1D0oO7h4tYlUMryfjA4HbcOr9NzEcXyh0Brow6/l
Jms2t38Z4Yy3hZZCVQg1SoYrlfETgHBCLO/xspHxRrLUt3Dsguwcuwj6Wggd7rjr
Cl5qaHlwm6Yc7AoH6trPX6glZvfHOJgdeSLOWFsABbXcAqxTYZGnVrDEjUQcogcm
eZq8O6fHq4LqX6rKIvJl64XG3iuT9PuprKNPLEckTueuywzxEibh6afI6982OQzi
E3y5H8mld6qON7Ov4vjcz/krFlnbbZwIfplNbflnzRBrKKSD2k7UAgJt0Kjdz3SJ
etyO4ulSm5bncJ30TPI7X6sJWU/RQXdcn/VqBSJiEALeS17DRwUvFpuE5+mGNW6L
Xm3nquezssqKIN2F2Fj/DlxnjqgN487bzz94RROUXARiFEGkPgSSdk1fMFa3sRUj
zz4wtVLNcWRmC2e0Tk9OEbjBsqK/bQeWkFIAUXY9CuIeoQP6ptDuDgpgFk2+zzL3
29zcFpjsS6b8JHctSO71Nhn99CXEtwa8PejlOJzn6PVucBbAmDfhh0iR1WrPdH+0
8Minb8qhWhrFrmx59q/JarJTp73RCtHg1Due/3/j0i3jzZZvcbbMJDz3cUWjsBeP
il4k8REg00rxo5Bdu8/P01wsG7DYaQikYpcZUG9xiKgFZM30XXxKLyQu6azaJvPZ
GPY7z0ikd+NNfTKFsqUlFZBCBl4PDRepx1coiB1XUgi1f61Gl+LrkIDqzR3C0GOd
tlltZV7r2JqSEcjhrWApbjBbaOIaszC8Ni6HfwR7vfJPBwPM/H9RYst12cBrbEQf
ejlG46Qg/1QmrKBQQe5+Fu+7qDbBC7hbSWytBXB+C20mUGf+I7hXFRsE5eVIm219
CchXsDtYIBiRUfdyNOTuQP9UV5jO2K1lVL6SzX1Y8vNjEfMQ2BcmMknP3Yp7403B
/603cPffUtNqwumztk1VXIhSWW8rTpwHPwBx5vz4Y37qEi15yArC4FrhkKiCNLpi
mwII15UpP0lNo6SScugmBKma6Ipvnx9PegvRkp7I7D6N5jc6mIWEqeESDXw4XFWi
I4Zc37M6MvEfR2sICvIPS/zujKdXsVmA1CZkbJQXkKXR3UuJJicpzSuKwkDOWxdi
ku3lE5L0Nn2rKE6y+8cO4un0azY5OZP4hMo+VF8RzH2asLFv0sJ4UJbRcKdWyUDE
Y7w+RgnBgHinviWFNFC/LLykv7Fy342sCdu6n/+oywiNNaR5Cj0/F+mAdX9XmSas
s00Ea/mDCT/9ERItpqZSItRjR+Cnje84pBMDlQbkcK6ekZcZ/fDLadGy7FX1APDT
IUKUKXGL5HnIJqBf85j4qWBUsKtNuG1tpl0L6nrW+gm+W0pP/oxBKAYKK+GuNkls
7hRWd5lyQTYlpxnggXfOGCJixDTtQn/0M43L5x2sMBp9KTIfg+phfgh4Qn+/vjeu
aV94FEmjgmpxAGG9q2UEUU0fE/9EeGDlxzKsbSF7UrPFa3b0zz2IA+7ziy8QkT7G
gHk4kz0kPQxJArQmLGaIKn29tTMoWSj4BEKDxZL3X6/qurkpAb4ZG3pwaz/D6V92
MmaHYYNx36rEjTb/+IMPTqeEg2/wKoPpSbo1f8fsyJbZ7aMeQ29uvfT5wl5oCvks
reti660XoZfJS8nxd3hrlb9BxTuqVIO+nZu01JOVIU7Q2HNsjPkZ8C7L2gFmQqIF
P0Zolx0F90IPsbPT2XjWw3o3r0UmTU5X+mo/2TCzvFuoor669SEznb3iGlH68FkG
OrLBoyc2bZt4gRvC8PJqPpRbZ0vhK5mTGId1oWxEIDjU4999RxfcrQET/61cdUhM
tpeoINYjqwo8DOsxUZcOqPNB2om/O3niEf4Er+3Vk+zFgpiD9eu3WS6oR5rwNUDG
secquMp/aiasQk3q+dSurqSHMM7+1RNMFYO7n7a1MJlsZ8f1bVxXL3nJA92K3Wcd
MyD3D+1i72dBI1CoAbffATYb2FaGuv75YZ8dY3ChxJ9l0JvQWQkf3mbZ4/AFxGnj
0HLo1ZvgwRDKpICca+NeFzyOjK4ZVLD70RfeTeHP2/GS2ksM/PTyEzv0F+Dwby2I
iv7LMfLldoZyrnk9tL5HNJTbGkfeXDaGN5SKMUxupemBNfFUVrgv5NbKnTwXMYeb
5OYfCLjnbTT+M1/CGHohdeV+xGh1f6LWqR/H3u3gEg3m3dP9RW7+Uv4Ot3w1IHpq
xsVfMo21Eiq5U1q/mLG2cqpPM0ZraZ8iaEaoD9KukwaWI2I6EpkD/bqz2ym+uXhu
RieVep4gpc1Yfj+/bNOwjY/anMfKOu9LuIGstrGlhbRbyiq9x/cnGDZRLo7V9Bqn
SNsMeH7xaORdeX1CVBtWpttqopFFh/1BGuYPQtSxASHy+YElf8pL8l8lhAtw/GUd
lxX3WQ0dLtZ/bRYJR9hXWZdkJXHIo8yaUOLHhMZqkf4Pq2f4AM+I0EJvSCaW96tA
/nnI3Cftmc90vd+/7d6SaS8QrQiCV76vojBWyHTau8G3zdcQi4/gG4VrIqZL3I8/
3WZTeYjIEBmpu9SYtGJU6JMVFkydZhz41cV0Oyylc34IAEBTVFuEoQTf1kVESNqJ
6FkAVFSC7sRQHl7IZHUVVunC52Vshc2PR1wnM5+UBhf2AjIMlPYyYC+p/xBKu8i/
sQGSBDgdVpfvAh+Hhhaa7BvSPaO4qqp6yujtY9qedpglhGk2Ose+purFeUmmH4dj
+pWGZwa5REfAP5V5KgrteDEXASCOFQyZhSKM+k3dyvqNacMApVBcT8YTFghYhcCe
FUqc+3+2Tk3m767bX8HkAYaDwn1OVeq+4vhgn07+JHqlbwzIzbVgv1OFiYRo46gB
KraG85sLNShIWHCRrdIElJa3VmXsn0Ck+olr2ANEwZpHBIGFrXkBUEe89tUGJbqM
IlXcXzkeuC8oaWCPI85R09ZOKwRU0zDF25cRceObaZX9w6O2ltrJx8gu6NL12kxE
ycnN6RFMpadaHFNtiv53uTzwNueSkN2SJI940tQIoEsp6daMhJ6Zoph4/jFfZDwe
p5Y3oHlwybqZAYXjma2C5PFt4dSIqGhGhy+VKY2Q7Jgg+yHVL8yxYFXedlmAN4PR
cWZJM+DzIuXHbxw3JE8UnqbVk+yajHcdBJoaghfa0pPjctVQ3djRQRVNS0TEVQpY
yuAqSpFxXJ7TcPUk1I2Izl+Mxn6Gr1Gfnp41c0i7guzjUqVVtvNnmutnH8NSvuOT
QUl7rOTvb7Tq3wyrruCQjHzq49OAWq82lpx9jw6pEtxgCrVDb4GwmJRGnaIu1g66
lPc1mNK+VY+sCWG91DREMXCyf2eCw29o7h37kTimok+qN8AhLTMhK1i+G+xc2+WN
ZFLIZfTZGODj1IxlHWTc9NTybuYtRf6gC+OxLVRqdWxhJsnKH7sxutZ0oifSkWeP
4INruGnzxYfFqPZy8tPVvLp37As8QfC8LC1yi0hoZq0W9DM2mhyEh2jB8wXPOFHE
ArHE8lWCqg1N5MZ2CbHGfxm2Mkll1P7+Hva1KkKfR1DeweF9HYVh64EDjwevUUAG
uNmNpO8NS/2jx+cug5EnJpWIviMM7W00ALakk0hg+cncsS4Kl/0VWPmonRzKnMU2
PzRrkqjEecqmHHxXxe2JId/tA5TRwGx7VMICzhnsZGeIoR+41M9FEJjpua0EZq7Y
TdlIkqnuZbPFB0aXn2gjQqozDcA3l31uBHB3pWslf8MXCJsIYatVi/irH8XJPkWR
Qf5fajJYe5nl0ZFPGJeK6AN+6AL/1BAW01ksmNOPK1wziSZwjbAxyj2u5EKmOeNV
XWavwhHTowNaIKo1u7pYH3OhNzeCLw18S04A2MWNNE4=
`protect END_PROTECTED
