`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u07+tyGNWDSceQcqZ5AR5XvSnC0ofB0Qp6aOzsaiOdazBbFHNgSDEbULhgY2tq6k
NGnA1KAXVoan2nNpO4jMc0ALV99aIiRAC7qp37HXjKIkzsiEouar2rc/uAmes6+T
FrM3GCaZ4cpXt6yuHuOPj6zu6MlgSc/ajG8flEy5/molqA/OiADA9AAoleoXnlsr
LtX8NhwbnUk3F3ex6lIh+H1XWSrRP0V8o490kdMy9CEuIM4vutkFfomH4kZ5E1Yy
RHzVHbN7ZF3VRWVtFU/1T9Wy8fq7uE/8CGzJrKbOX8vXYH+o0CnVB6WZcHHubwr8
w2or6P9ZSId0bG8vvB682wu6I+P2Q+Jh+ChInMHAman7mLvtcisd/rdOH1D6bG6m
QAN8lcQKk4t3cXcMRCdvqNd5okwUpaQEpppo7nZxJy2BNvz1bXa4q/6AEVMdX02O
VQU7z1i5qOqncp1ReEkGHRU7epfpVimYRjTIK8+LFGA6NSNBE9xNNi1E0yARBaXM
PYPinVShQRmGQffD0l9Qg5qzWeBnUe8m++0GM/faRCRdHagVDEaKL9EZbDc8TL1n
BNYGQVfpzpWELQSvshzs3A==
`protect END_PROTECTED
