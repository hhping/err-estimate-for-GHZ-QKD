`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zdfvXlc9Fu6HRnxW2EW81BfpYoEFqe1z3tkl+Hxt1g8qmjcU8NfI+NbZIdTfVaUQ
I9ObFJLqv9QPyu/KWPDGV9wBSxiTxyHbWcGqpdh+2HpPMrKYBXJrPKvjxZWU2Oe1
lsyBGts9ArCLs//c8aIicXLH2uWbj+TB6Hl6Lc+3wPXqRRQN3O7LG6BCnJPmlsrs
Be0e6W2liJrILJGf1GtXxNaPaG6BhMXUaggOyBEbnglphgig0Zi/u4pTYY4VRHhq
1YVj3C0yCskE/vQ0si0EfSucDLlyKnnLerIKrPQ7whaHLJ+Y+VwNsr8nYev5CfvO
UYp3gRa90GpVGRtTrYSqmsmjGtqDn2fuYHNhwrI/btFWMgRBpdGWhy3H1+4ti1uP
ouT51ro2dYS/8ZH5GHFNGs3QXdaXDGJMc6wa+IgnYHcPLbgXx63aSp6bw+6Jsvmj
5KPrSI7xvkIBSrNmbIimUFL4WA1GzUVfw4HiYjrfljWvf39l0YMxiBV+8i5D0oye
J8Nf3ZQa+HzvLgs1diwMPpKwYIRpN6ziR8wv+A3BS7nzTCkrSjjxKUbNDwUbbu1H
FqvvAkw+WJZOC/3m3gHm9xLNJr/mVuslaB9xXXIx10pWVvYGp47U5UwS/NLoln0s
QEv1n1nFTHYTaDQrVsu0YfamfvLqCEIfMTNX2g3eRa0GkwvZvh/5bZcn3078JeIO
x6h1bUZdRkCGGgT3QKJgwWR4MDK1gNUQhbni26APrVrqHCfInITluPmoz5yJeObJ
672pfpAlWcOrUKrL5J7Q855DC4fr6DR+nfhN6PAiP6OIuTfbKpSGGp4NWdBpMokp
+f9giGxjSmfcjD7M5SqovKik+GZrOKvoGbrQWrgsmm8=
`protect END_PROTECTED
