`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DGkPuKWOatSCnuZ0AGGVvMMX2UJnUDiHoSdUkB+PkFgt81aTcNcS5Uconwu00SPU
Fxg75+15FxA0lViA8x256Q22fnq7T7F5l6fZ14jOCJKHGXrkkna8lTyZuIfGYHmG
VfqvPAn0PRuF3khhXGGywcP2i6Puzygoy/RF4tj4kvGL7LF3a84ndrAgKxl2Wffx
aorCrxUbG2T7Y5gruoi8z327XzO73oWYwAbYUdY9+ZXc1XnzybQxGFDQz7u6IVox
IjtPmNZdTTnNLtjNCwrlW1Lfr9pSMeF88h+B201WlNEHjZq6wXm9yS9vgBMgM07x
K+p/5QpqRMe1BWoNePdLJ0xtk8aiqm61UbawMDwdHxbTz5oEqYNKbVzlbcMhlfvl
o0V47y5eVtVW8phdJMK8lQ6VKvfcTlciKqYLLW6bvhAQSp0g3JtSwq9UiIHQYZyS
jo1KKBDTKyJZe+qE0UrMIBDfOWJGUqOjFDOeR0pfQO1fYOOwd2Z/o34gmOy995/4
5A0JwTvGgNDuDoCwOo/XXrbPfQTRduVS46st4yTwKbX79HX2vFWV49f4otSVz+n1
s8TWjWALQBHlAXfye2woGv0Tu/L7yTAB6Ug/12QfUAqCCUZ5g6xxzFwab8HPGKYt
Yf66n5aFSeAI+7nPM6VcGGFVVTMt5EsxVOy2WhRURHd5v2frgKbNUBi/4LZM8Yst
2D06chx4Bvx9EUCVN3BD8w3DOg6xYtl8yacW2UN6zEnmJzeqJ5/iVVRs0HVyCM/I
r7mfhAlsMJ9+U058DNCA9f5poAU/Xx+Enjnr2+XLQ/JKtBdieLuiKBKAWr5/lXPL
GDPhPF3xqj7PgTDZFwDpk6CJSWK8VTBM3OYSli6hrxReO18ZMdPVjC6bHyBlBnfv
Xmzcca7VgHqql3YcvDResHN1+uEgf/8+U6xFzUWFPwhoUhhRdcd7pbE714F1VcKK
lFHmVApzsEgh2HKpJrigRUrm6Q/Zy/czY4EMJIa3NvAj0hvEMqz6rd2FDMxegoQC
Zd0InMxB43igPMOjVWzBDvT07FLWTbgekYUYoOU1Ar/vH4Et/fPc3DF+Gdr8ERTE
Br+6L3iLA3tPlo2lMkhTnEPD+Z9Ti0U2k36iaCRQd24kVzT8Bx8qwNjysZyLslvS
O2xMNlfpiwdbR6lai960QvMeCG5DVxMmCgDc745duK4NZm+SmJSRQlPMRJygH1A0
HqqDi5h4lwWrG0f5J6JJh3aj8U1ymfaPYdmz/V4MNXvIbyWyckILs9ELqtUeMhxo
x1r0CXhcTwvV28x/CrDNvPtEdYGTqPrvR/BSyaupriQXEwTiIjAClKfKUW9AGwRV
+yvdONpMWWH6scDiXqwZI2E7+oPqJxusVWilTTqOGk2Qg8WFYpGeFm/uL/onR6Ov
L/W4Lo2Jo6CIKfiemcaFdgzzRCcRlZpMjoRay8fkt51EL7h1o1ScJQyPIboKsuKX
`protect END_PROTECTED
