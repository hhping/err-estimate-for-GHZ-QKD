`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K0z3IOtJ0TBbzuvFzKvpRNDOuwxNotgPvQZNrIDUC/gDVIoLuDnQWmLWyrcWDn6u
pwFJ9TbFUqhCrctSQ7TorYxSU3CBDqB+fPBCKHRyr7LmZ48XgShov10R/dtgk9XT
z80bkd1e6p62RU3yB9RDH2QVtdOXnBxzJT93Gih3Chbd3szaXjnfcnpTumGIqWyx
1tP/UmScIa3aHcYTOMKk3q3JU5zqaVMRaEu1RP0qbLBAb4yIAmcT5JJZFqxUJEHv
QYfbRgDTe2uWeKBtOg3fZHej1SAClxC5QIL/a54XCWijUbIPU62I0l2wa8FjdM1F
N/WLYlOYl1y4pauVdoqPA68lXqAHpvLhHjnsFvaCBEzea1yjNeAmO5s28sObWmes
UyLF9ZxFMbVZq/iO5mwzvlt+kFYcz98OHzGSVsToLHRFHNDs0bPSiLTZmXupHDdT
LMAGSF65IFKkh5FQZ7mFGy5NkFy+ZBhY9gfRN5KQr04EbAN/xZp/NTQIchyWQDjE
1z7BAba2lGlKIWdBOu1HZbzB1wjaDNeP67UFLWzWTRFm5yZUzM1Vbm6CObSIb1gv
L7uoMa48XxmS8Jh00ov6G2welVJRvowJ+bH3szhq9yRn2B0RHbpk6dhVOkve4qy0
5fBARQmmCR6oxQsrIuW1qdfeo+3e1Ht3pXl4eb4Pn9NkaE4V5/90c9uXnbnbxCDE
QHu367pMWtGLWzD2rpjt40Aub4DnEGGDHgSaXdQZLWt6WOIPfdhW3pMuhbW9fBDu
nBSysARAm3+RenY0tNcF5LLcZcHNujacbD0FUp+LcfY=
`protect END_PROTECTED
