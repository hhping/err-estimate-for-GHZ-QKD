`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a9ML/OkIz5TJXke9qkPO+VYcT5g62FVLbAjgsOVpr8FBeBu0cBsYpHOtuehT6qgr
dt0T3CPp9fRrlD5Xmjttlu7NyYi8i+p5klUnw+0upW0i+VhCHt1ipMtSsj7yW96v
3TOd+mBYteOxfngQ4qZTZIPYDWrNwBI1eDoLenhn+B/pekB4FbelI2+SUTYyTK+F
3FAsBrF9K58rRRQhgwuCvMbJcOYmZqJYscFU6k6a0ubChUiBwhzgiAtDPe4czlcX
a0OUtB+cWvzhqevxQBcgiRalnyYBxjp7UIAyt1eHSZgGVw7frSiNkH1XHGW1lOuE
Eo9zIIkzqFifrpdhTPDB/naYLdjK0bJZs2kZshFUtetfDQmhXtc5VCCEeOiJflmm
JWWyUIa4GtNHavBBbN5kutxmq2Vd04aqXgNNSksq0PmxZ1fvjbunnL7HHIDYENJk
1I7Ik/HSKoPTwXNdw/XxOz7SO0njAMt3wcutRmNCu372m9Olk95+jWEWXmSP1iLs
/LZmB6BNAX/6u7gNfSnFX/ovHrMrCbbSYVcMJEjfFqOxBYQUpHVIS7QVREQMzs+m
gPf2ikhNuONIGeUKLhHtEE73Hoprys6NFpHXPwl2GYUtkV2ts8B46T5hDKyk7EeD
n/jZAmzb9XtoZCDQw/P8cxwoa2XZCBvHHO7Ub83M4PJXA1TpcqrtYc/8ELfBfFcd
w1OYmABW9//DE9zneidxm1ZhHzltQ816qXd8ujDuBgEpuLPk4ur7tPwP84MOI33i
Q9CAr5mO7Zxs07YNQjptC7i15ZluJdEqXQ0bVIXH9MTEGjXy96vqA6r5nQHrtmQl
uwXeA+ATMeH4xrS3FXMUCIVtmaHX673oyALlTBN6ZgaDHNXOm2hRQL2ltFEOibIk
`protect END_PROTECTED
