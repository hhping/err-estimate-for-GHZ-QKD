`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8K3gcd+IiTjqT/rIfGv9cwfg34abUGzsAmRy0iAfN+vhXUvfj4xFFEgC5uFv873C
mij4kX2hvap71vkww9Kj6/VMVWL5CqF9NEkY5wYNYd0/zs8p9PK0HK53zMZkMRkS
SV7ywVgs5xM2iqYe6A8KnT+b9klQTRpbQmJUyLAUUwG6Q5PsT58XE1lPqavZws1n
rixl6M0BXaKwoiPcERqW7bdeGSrF3zgSvOtHpIR0uftmuyy5BNvEZAfGXP+x5tZc
rra64OqEH0JuZC1ErN1rn8SqIv75keFNQvVg2clRJSPc7AB0nT79oPtNqL/DW0MY
XAZ1mFyJE59tA3+lL339Lpv4cB6AdhC1AnWWoNKu963vVirNZxmeXRUbPtAkcyMB
Fz5HJXIKDrvEa2X25PObdafCXYtaCWuXjT3WnQQ+EhyIPRMUSfTMLq+itWwpW2S/
C+bGL+zlmg90FVMQDJ+8WZgjFmeWkQUFqRaLsfHnMNfXH/Gh6ilnaqnfTJVHIkL7
WEPJlVT40UfgyH0g4+YPJ+jFugsXO0AwY5NHeRHzC7zW30e98GC2q0fvtOBuPTXX
OFyc4DgXjOt0I3Rrn75ExITY0ActCOW2tRoGRTN5c8ogfSLra6m4/jQyR7np5/fN
hUHottfwV8R2zysB7CN0PCm+J+BUddIUIlCMnbB4HcYLShcsiPXE8RH0g4PL8Oqg
Hs8uj9G9n9NuH6Kx+JFDgsqDB/nMpYN1emhTIQ42Uq5VNTz7vXKAZYnoTGop4hiU
PYFb/wpK+LfG5kDag0zJ4sDspt3KCFIygsRn67YKgLHdKyDkpzAIW3TZXCMh+oam
ai6bq1Zo22VIN7IcUeESEb8NzcuQKdlyhvzJEfq12Ekse3h+IJA5SxHfAHT3EMHj
7HjA/3ZMTFq2yhdCAtfG4+6Bpvyb9UpvZmDwTRkSeMpVPe5ljbavgZKvsC9Sa298
qZVj1VybCJQRvgBvV7yZibU0hRDFda06oVvfeWqHyp3+GBxag9ed51ajMAkeijVv
QFdRsAHn/t4HLuBNOkT9Iu6b/4rccQq4GBSPm9h8/SFXHWjSSnU4Cd+fn25a2cL2
KEqLaEzGjsmBU1HDOCb1znJY2WsdQJkgHm4vw2PWCjQs+HXIoxegQ8m3BFoEDtQq
IxMFcoc9bQjPD+tdGWDq1g4lqQS2szH8XFc7M7O89AWDRmyLXVbP4Hs7qXsAsLIR
NPoAoNwDjw2mDkCbiA0xe9e5bkIDFMS5wsAXC2EM529HFHjaioIOGrLPARuimQwR
XTO8xTAEHvx91akbu89VLMXiGI4M+vJMyyHDOOOb9YQYsPykzIqqW79ec6AJf7TN
9DXMPxQ9mBSAosZKWkJW1viRwmZaFQePgWq3kA+ReWfBQ42VEQRcmwvECOj8a3fO
l7Y0PkGVdrVbP+63y1bHI/1gkhPPLVZyElIpDSnudtSk8HG9w5so1tsP4C6G1HKG
HxTmqbzhUIqrUUMkKmMWR3CmRBAzdXytiKHOf1kCcNGIBBygxOpqVa3JarJrovFx
366mmdAEDqZdJxmS6gTOKpzgXDGC88YuHTaJUaUZdDopaKWVhVKknf9C6ekFNwzO
SQgBxVmXJPXU807yjQ6dJbrLOTZW3cZxaqcGve4/u/o7+FR/P2jASb0lxu6rhlXC
bafB9iBboHo3/24Bf6MXKu01hS/YpkoivBHxyrgrkKK89mHiqxSOBKUJwLOEuk3S
a8JbZSOAAbXHyVtvL/cy//aO/QqxpfhgiLUK0KyaIdLlWS8Bbm1Hct2cfoWmR2gf
wvUGCAnbz82seLJWvrVgNqd9/aWSCMN68Ub6GDZahwO9N5+eXqwDuKcX+JmjmrK0
cJm5vU7sCXQrzbak/oq6Ww7z0KJ+KAHo+JJCbP8bKZYIpMg8g4g9wmZPL/XdyQix
RPTWCr/c/RblZK+tBzHfbIxK8SC8DfFur5U957UyDcvPIhySqgc8PDxDDLAm6PlM
utx6OWLN+5wTmskkjHq39a6EV6gtgY1BcOFR5cIwoN9IQKdfgYjO0lMAJl0XifxJ
efXijxguaZfjIEpMz+4TvI56o5bzefwpSVXK1UADCC7Hr59Cu+xZ1N7Oa07VFPwe
yk3+4JheJjouhSy2n1VzmS6jMN1eAIZLoMsxCsqquSJ0Mv8cAp16rlT56Zhl3eiT
sBLas1+xcWNDAO2F56VJeqoR+kSf3DWCTvhqqDTH2UeJb8jhmVSXGMi8uETM11+y
FQ5TbxS53YX71C2oBLyVKiaiJZ5LPq5jSeK+t7OYihMsnV6LT6j5Ik4qv5sWWeDL
Tge829MUfZQtBT0x3Gf9KNCaooS+8LfRIeFTQtgo0+RYs+jgo44OeQQ1QRXsIqcQ
4cRb4bmG25bx28gjWsC/On59CZ+PVTexuW5XOUaq9K7B+ic7rO12nRDcYVrG0900
rGwKfHDyWsb2ewXnpB/nb5tJitZKnMJPUuqSu8qY9XpAEF5YS6YJIZ9RbN+ElYzq
2UrdywyqhI9+SnLwErWJR2EU8JE4Uy7PPDtdzYJKhpW378OwgwTh8B7jhRS+CCCJ
tDH50EZzIQYq14C8+7Q2NhalmE90NWjrSRB7qMlU2RgRCCqbrupkGhcW3hT45+jo
dFeFFY/aj3qmA2GawSoMQ3cMXBe5h5dNQ1hynLimO6FyjuJOKTkP5vkrr5fbZ2Md
WWKuMtgwVoI8WYVbmFu/f9cacb7HLq9CdlYmt8gwi0I/ndzIGW56Adb3ygB3BNUV
hWYhDGqovQy0MQqFuaLDQO28w3QdhgWYyCedlDO3JkYbR7Z+DBV8LFbUYEYd1YD9
8vtGyKUVmfwX6uklJ80w6Lyx+3h1KJ0qVX5qBRxT0LcHChI0JKs+bsW9jws5Tgff
CQjlOHn1CJj5Sbo16Srk+7RkxMXJ4G0PnRGJUInDeJ5hQVW3BCA/bVK5flGGTxZ5
cCgKp2qYizoHTp/zZZxgZI31a+PG/duAbfYnJfu2s+eGChyw/jIKZe+DHTMgxdaN
DDTTD1Aeklmv6JMOrCq71HTQUU/30CsY1QCkq8bfVgbsKhqJF3xXQDp3IOzZBcJo
0ZIR8zXgOGb4v7M4XmrtIRWzeBOYMosstxn5qilAhwQ1FmUsn6fdNGQp/QWlsJtA
heA99JC4eQt43aBOLLKjfl3kMxuDB6cBfFAPNaHTjkPvQD9UbhuqUPhEGAKgLkRz
jdleScRCTGCer8EI4H23zzUnTAX4xX3gvaUCr6dh094s2tgsaH+FUZx9DFRpFAKI
AOTltxYYuuEyd2xPuv87iiXd5ZeCS4D65wd+CnEyWm4FPxfQHLJWjfeaTdQaE5xH
+07z/vzeTvdYnpmROfN8BD+2RO+YpH2n0O06lth1qJ3T0H9WjG/SfK4jytBTbcNi
YYuyf5VCs/F1MA7f+FLSiGfvEaNbStG/x5swWspL7ne15/v0jcTm1HKqfPk/jE2g
CbDcH5G2iCpRzmroYGLGrkSAlElk8emZgBvRlsfPrANeW9EOYkW1N4U7nIAseppb
ZQDqhI2DE+jKXxJoxKhDNrdpnHZwCg5v8FTQAvdEXx38ZXyFxi10eyy8WAreH50/
YPRExhDiF17LR1dbbCzP65rCzelqcz9gHml8sl1AMn1A7nIX/cZAvEGdggKXm4b6
luVB1JSDBCMQ9NjAb5NPB97yfiAQShFMXy+P97HwXTk+vQQmxpmFguROjK7FOx6h
okA9zgj2RgaWlJMqgr+X+AWn74PpzyEokx+hwTCkxmtxQCiWUNlbdYOYA8IiBD+5
6zrf0JIaTEoK8QghpCec9YgB68uC/0jWHcrsXIekNaIRiijzkpuM3JMLTqR2jVti
W+jWXvHUtwY+s/XIw9GdiWEnl4PG5Sp0T28072L6n+aceh1qtWoBbpF2JTvdft9T
+Oi4PvfFC85E8stIldVCA+VIFQXwGBAQUxUf7orxodcaUx7gIaEip+D/asQxyZbE
0j+LaYzIxHntRScaCP/mxdYTlB/DX2GJSXYKIbLPVj0GFAIZCc+9RRfaHAJOG5z2
INwQ2N7ZnqQPzmAAcbVuPYJguXidraeAqreyDGxd9zTYMOhOfXrrZMwgbRkDSn/i
bR6g3DbjlES/wQUh3ACnAoERQn2hCcKbhxVI8d+XVQwVQABNAIUZepRUEdHDzYMD
TIM3JKPlYnBy65V9eKwZBjdPDqxIw4legflWNANdD+FQl/gbYHd7ofdOr+mZacNK
4dPjVv/HDBgjUS8vJ1+lURa1kllSAXEdpDDxwZGeIEhizrqlYLP/tH0TPiJTKJdv
7/TeujUXcWJRDuBU06vTLFnCodAup7tOlIgDdO1wY5NEtYi1U4velgkCfQcmC5OZ
AirDofzRxA+6/W0q/cjYFIrWGtbFY8fJhb7W7g92SxjHjKaNhh8OqmcNAZxAIyma
4t8SP2PKVT1NZZlhLyZJYCFJEaK/TgR+Irzu0RPK9+4DLvzFtQij4cTbHjvHzSTD
CskyaA40464lYc6gblGIfBnXXkA1DhKu+ILIyDzhxQ7IZi7MKMBW8ipMvkTY6u0i
eXA5is+/qcsWUyFqHeIOlX/35NQM40DfK5NlGIlgXmXtGkrlqLCBpblyG+eiC09S
H7q/FddtBQ22GHxn8/B2Fgi/t8D1C5QOp2B95S/mauFgiEj9YhlO7BKI9B59oAoX
Cihxt/zeBNlNs+9ipMIvnTZmvbgIomgg19N3uRpURUZnVwjI35SL2dkUtq+GsPuJ
7Nq4HlvGYNTa5BpMeHf4HV1FCQlglvrgLeXnzuUA2b1MpaHxZRpsGdrTG4tQgibB
hnx/2Epco7MUFvY86QFMeWKKSVyJgee7gTWjfVgkgXI1JmV0fuwH61YKsUlVCAl3
9062SDv3bo1c1C9Vqb0bDyjDHOfi/sIyU8tAOkKibsOJRVw2re7J0KvlpOlc1uFP
xGsFUs/Ra1NPfs+s0rW+tPwuie11GK6Sc6hjKgXNo6eRh0M6vYmiU+IoWG1CPdhi
uFdhZF21Gnxg4PnTyX26fj10FMlWhr3NjNujBWJ8lOk+gJ4fRa4dY6j1biqur96Y
tM4YfJW2Y2s4UyRqeKAhMRqBVbU/Tw/n3hogvEb8HQvAsmS3o++bmctCqb+g8N3D
xaFcHs3C1OvS8lTQEm8QEuqwKksDGAU6uaRFbhOhhR/tUHTx3DjyZOR4dkk+Yyah
X1/zx+19t+hxHQFL0VpwcWs1G1qbjYVvKbgUI7nST07sDJlJ2t61n3sgSPg9Gnza
TWG9Vp45gI2ePTyHCprsR3Fe5RHY7+BLNsLT6nVkaa5S8chgUJaRvYeHOYUal/+a
4Xhc6hPaAC2e1vEg068566Ns/TNbT8dDepWH3vp6Ca+JI3HUHR3dO6K6583bmjwn
55i1r0Wot6+yLRXZXANIXar5vUuaZjkBV7Rbwn75RgL7ms5UyFAFn/6fGtKeuj1r
oVlMoC91fI1zxoUUHNBst0zg+L2RwWLqVA/KW/r4WHrQUtLY3wUrnslY5kiX8p0L
aJMP8M+V6b4IEzlP1vBNeJNsS3t/wn/RfuZW9cP71S6gNIXKWRY+wNdMbrKu+0y/
/E6fSMUkjF/Om1OwlQQ2K0zH6HmwvMVAsqGye8CT2JCsRvWj77yCc8cWUNtJyjtj
hETLhOLHg1FJGhR1IEgy9gntK59GJv+G1MXd/6dkGX4gu0bizxriAMkzRWAjNcsX
l0hj2LL7nOH/RlNAftkCc1k+aufJpvcLov73norJOdv99N79Ea19tHjN1ufMY1kX
EZmuBGHYxy+l4in3QhVXKmC9cHE9rNrq4dtjR5IvHI8lXFSGDGPsEEOCPNnx8DAf
0kos3z9Rv0bDBgOxTQDVp4mW7pEMJN3XSSYzowiI+SSscDL3QC4CV0O2PjQWaAhy
U5cWHziXWswMkBYZkies+0060S2D6xFlRThs+iCrgPC/Ax7uRyL//1DJnwWt1tTY
NOp+MVsPq54L+fJCgzcRlnzXoE7wXky12HetpbHjr11AXhy3lYO4l2xQ+HpG4moq
qUbT4dP3HgD2g2PJRJzMT3vHl2mY/0EDiqAT+PKrCYthXmMehL6vHGLJM646Gf7R
SeGTdFD+W1siVwzumclww1/ulEYSKERsRfjpjppLfvrCW9GKzLGjatzw3lSeo7PM
DQQNSHzoRp6th+mg7kiehAXXIyzk+xlzW1wccgTCCLN3DvGnVdKMXbLCcrnw+T2x
9Rh3zMa2zVB/i+2Lriu6QBjeCyBIgrRVUxA+SBdLDpyPE86LTiNzb3pFWzm19omp
Ig8jHBB0BVPMY7ahb0YwGw+PYRanzcXMg3LD3+TQlnqutsk8aU4iI0/JDsR7olVM
qdTt3/fjlPc0s+9NjHFEujZu+UfiNfb5hkr+jvAim+6viMYyhEIVqyjRZOPs5eX6
yDighQy27AvCueQdQQE7zXAMegp2CtGhjcArjK8/3vKfpszR+Dh5LqFQFIu35bvf
/y/reDJ4D7WuUex3/oiCdMypi++zt9CCgcJ3sV/qKIGBh9iHEH5zH06r5WgWGe1I
w+52ChS78+9dfGXxvr8CmNLRJPbgQJSRIMLyYCBivOrwr/4eYffKghtg4PDSM1CT
BaoGiBaHG1vqC2pfk/o8qy616oleVRdMuy0oFZpDs/VKKtoqa31mvose6Qt1/HKH
kt8cqj+clzj1FdoaeCLaAvCogRDlcf6ht/U4/65y+jSDKJCzLgbO5tuuH3c+fJwT
WFCuBYxLIf6fgCbz4y1giaItIYiVEh5HtbCghDG+1HtXf3qLNVVLgOZHwQLfTJFC
KTPvVRro46+u4+3Uhwn1mhwHuBCLhM/vhRMgSvTNOZB767fs8lexJFxcBnjXJCFF
z5hkqCQmVVC+lR+2/uEanORJP6F4QMVYRpK25vn3XhSxPo2Fm6m0fInyrce0nCV6
GJkuLAkjt/gURRinHCFXfMuGEhobwLLHa3qH73c43uODjvH3Vc9jp/jGQviAXVR+
HzhP9fH8Osa+xKsZAwDID3p45qH9j0US2JMM3yLX4cwbEnqxSm1Tvjo8+A+IvETn
brf2Pc6xUDRDPm/qhYdIFeEV87eRoMQYI882u6zpI1r61bEgdqehM3tK3vME7sxJ
K6lhzjI5mpRO8E5pBfflkmDyxSwrqufA1o9flDgFi0RPriVZdT94NbhOMCJLg/Ju
BHxHZjSbUcAkS4UFCmW3cZuB7+Pm8Vq7Ip5QrmOnKgWDB9sIWesx8j5beX64Yanl
7Oow0FlsGcMI5yCaGfLUNvbWob2YvjC7JPqpUGRE/ARgY3M/ibmpDvzoA/+9hu6d
YHZE6Po2Qv8jR3+g6PG/Krn1f5PqJAHny0gQU8kKxtdkLyMqMXUin6LGIZzsWNw8
0IAqvswMaUpSysbipq1hwgQZ7Za3VMQ6lN7RH0FxpqDmWsmBjD4f0LQPv4U00Nmb
HKYxj3KpVmOLOnU8ueG/nC74iVtvOvS3mKkAiucvEvayqZ5HCpKVQxKCmMVFfluG
XbdFtyzfxOxeXCcKOuiciMTWI+yA7plRn/BqGeLTXiaHq85zyOKXWmrZET5nACzA
k8qwxM7BhSNSUFWjImyu6l/mPJll4oP3+JzNzLBjwuy63vDSbPg8JylrteZHSmw/
YgnQsCDAbYtH2JUa3PUbJ4pZ5JK3ehbCzTv1IPyCENsTbpVUT+EkpCMTD6C71y4I
ON2OGYXhvfVFCdm/WKaLmUQ4kG4E7SpkV0GF+77zfGkIzDnrDNsrf3TMcwwiCpVR
78ClAID9+Rr+zDYR8XLjGj5DGTLZX5LJCGNpGNdU0cwrxe99jTzZuPprMIq43VA7
iEQnXDPU/u+luAl2udh5kPeWlo7tG5drUXyUhj/VnWO1v5RoZWt6L/UZkX7Og7/d
sX8GYsajC8dTjmGxQMdwfot9zTO0piv2c2AyctZzly7eSm5kkp6i4fYLvgqXXQ+2
sx0BQxCwlZeXNAENVkpl8qW6ww8X1Fg6AKG5FLj4pvuFMkc0rsw7GtEjxgPYAqwV
nULyKDNsjgCxbn3dXNb87S7yMPPXhGYIwETkuNkjeldqAsZgQRtBPC2t/7f2zhJG
EbEXKpAw9OTC6Ro/92q+uwEMJBezkFObI59E7X9dAOq6SAq4MxAUChaSgzLrMim9
p2ulJNduUEKMdGg3kKY6rU1DbcsFhKQKF/6r1NfmjhfuMC9V1Zg4Qtoc1oNRcpwb
3XDCl3tjDAjBvXj6TLV7joUbJ7Wc1++FZnSfrDiLp9LsE3974onbSg0lb0LSLVPT
qPK2PyhjAjv+LzS99d79EkZq+5HgW2j/idGG9Tj8eAZ/QQrjH0rg0bmF5fr/988y
udwe5vj2zrMwwpoYfgKw6Dt+FQNwlvdOOz8yviplSu+PS9Ya0ALCiXknJaZOYj92
ciKOyedqyzM6e3maYGWzlRvrbo/GK29k2A26KYv0qIo=
`protect END_PROTECTED
