`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GNlPXdzewT6eLMk9rYN4u9W3eFnizZVpliTPiJPm5xrzL85NEYFKX4ozgQGIINSP
q0CxYESDYy98mqBVqGNyd52n4tzx70A5K8bL9VV7HG+ct14JPz/WK+iDI2Llcfyy
TtdtXBxIX0IqrbVf1Iy//bQC75ghp0PM3vU92zdVXor3egFuZHSuxr6zlsVE7/YV
I/vFoDUNvWABq1FnDPx7LRj6fwSFHpbThYan//I+k+l/4rjo7B5NYjN/efUfmhng
0sfLte77R4vlYeKvB2Uctz/IZYQ6xGxZCTdAU8TcQ63jKzoi5pl90ITkiOezqqAy
yOJ9aKu3RDKbSl8eWLnodY5I/jqyEUv+1uRy295qh/bN0SvgXGQ2TUWq9LcZUPmW
7TngXiymPXJH0nbyTiu0LiSD6dfkuLDeHYr+0P7vfOk/C78Uyn7AKwOtVEPB2PbJ
ipFcCKygqUBH6I/lpqEZuiHNhuz3kubdeyHQmJLLMdN3OwWS9rUUgop6q2qeYVBK
8yMtDshNabjvGh/JnF6L9wWrEz7CfYvtXeDsKKNKijMPiIaldXe4kCgj3MwiOEZf
YpYtIW10gKzswMuOXAoxJqvUcvsNHaMSYami3uw9uMWdKunDV038BnmJiaNuBcuo
IaTR/411bnSucbF7b/AEmtfsIpZzlPwhgesNwo040yDJuT7NlPUWJ465JJtdrkGG
et533kxiqEjLZycaZLs2kW6U0HfNUn3bCkHngyxHPC+DMfTUld+5xlGzBtjQMLPQ
tFLdtptYg7MBB4XMcJRooxWiAJAdSzzQsoAOzwYsrDoNJwd2nRsoj8l0irjtaicE
hbJWAmz3ufFvlaCKSA+A540B5cz5j1A75GTlX1ImpNhXbvEigMW3jtlkgSFHp/lf
sOzLOFtLUO/KnMhrvMJ7FrNagudh+uMAVu7CY024Oufh3F/WZprio9egENSUh2e2
OS1aeWs+NFxaHDqZwXW3Y++OZS5bU9hKckBO7YAMlxU4M8MNbDCyu/wtIWzrfmKJ
iLSGGSsmWDNaqfVPgdMAjepoujxgOYnzovSCbptEhsSB7nOvJuJ4RDsBQo/7bDNC
S0dkqXQ/ouhihp3QAE5PwNFUTrBjPkmnA3WJnKbhzYtDt++pJdttM8aPzKfuBSiu
FSuLsq5da2oLOjrEQOIT96CmBa+jev8GEdrgxmk93UXwxy56zbJAlw6ZEmYr744N
IwQFETWBC4L6RzcNozSpgwCpxGrYAETogVehfNDmk0tojf9TrN9+cznddGgk9l5h
VD070aTvM55uoOd/UBbvI/XDnAEuGRFDofDAFqsBr/hchLX6/p67+xJSBy2c7SYR
uoUEEhE0GglbkCCnzblgkXlNGz/fYSLPcNXL1EjCG5jbDvJ83gQETl71d/FCmxQz
bkiaPikOLdpumtA61Lcg6RfWsw8HfmQGmb8IPsLTMBbOjvfZWIhescARQO50rgQW
AC2OHEozDSz/GpvT6JlcsyRn1T3nBRohcbfQIj4roXelvvFnPEfoCpGCmHFF1q7x
mVfBQg7SSPtkRUavXAwXnL6KDAtopSoFSg4zwXPt6NojNCAa5QGmslbw2BIK+IUE
9hyi7HSsWTeYvxPR3HgjLDVTjBhr7InWWLDEmtnPWK4Xp1ydhRbD5VKPZpNacnnb
vNUf3TYfINziWO9ja3vZou0IxXwue7TS4m+0qF5AIVL72eHnItBQDm4gZ8NwtPmp
5UVWErSEEkh/HFkRWFFBuxYpTT+B/TQrhJo0xJeK6U5WmNvbTsaZgzXJJ5IA3ntR
5ryonVCtUMeKjLYh8qFRMKtyM7kvV4j2cS/Ozfqht7EYUcDBTegNkoXdqyrkyNvb
1VT3T4ntmu2fLv99discQQ==
`protect END_PROTECTED
