`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NfX+wPNKJxnB9B84zQZuo3gVZqKKso1pYsBfkTK17fxQU/tQXCt8vYo6FcUTACii
TzMOxWeAmh6L+OVj/49QvqkKo5ndnOde8Oa/vH3u12ybKdEv1dKaWVvo8CHLV9mI
I/B7fdmuIrAuFG9w5wmpMW71EhnL4f19JxEfeDIHJneVKOfJ7+lYjNBnuN/MFE4B
/VArPbrOuFIwhk/XLZ0REwQF4kToff1N5X8sq63hfuf4KZmlMRb3UQ4updekBP5g
WF41Whan3bTUF4h7Xw+v1vzBho+buKfW/1grAKeIZm5vUM8pVWNY/iIb+SveGejt
Tk75o+qwjTB+OJBE9FvwebFNn4iriyBwghq38AewE627lF0E6KAb5hvXZKkZR0wD
9z19otrDWat53q1qYZBRfF4Yo5Z9e985WvUlxKkwPI4ApJ9K/i1yOei9QzQdFAgB
OWjMOJLsTSuTRfwHbwBUIwOjfFydI3rzT6GXtk5FPmsLgVqSWDrwOvfP0YAzlHdM
H7OZlS9qP+yaHLwRG2wSUW3HeO49DuTcmyG6PM/plWP5KL09gRubeCzjE4VuOIbw
UkUs+g3oI8pSTQl3x0pSxg7FNoXgUsvUG1IBpT6Lzh97GjqnaZsaU6TW/3a5U3P3
UyccBCbqcTWFuXihNr1P0hFaARyDHojTIZ9pO+bNl1MK2AVo1JjYOS0baHXnOKa2
JEks4GBBO9HnkQroofUdH7mUVINSzvhE5w6XkvJpv4wQ43monykyg+u4bTyu4MGl
rQPJMUXhFP8e/nkINvfnAJafQ34zaSvSq56fWrqJQsNZsD8MkzOFkyrvoZ7zkEUD
dmCe4+RJPxjR+0SD6i2ACcB1SDqIGWZUesjJhYhqNwAZhYU+5WYw3vQNq6RAWELC
O9A+QN23Anx09VAJ6VSBCleGezC9P/0mIr2A9XFiIYlQNmN2gZa5id0tUezTZYDL
AlDhk9KxsY/FY8ts7j8QerKfVU0HDiTj/inYCl6Hp61vqTtfsmSjiSyj6H9sheVk
1BqgmyXbh2WXTBWe8rQEHoM0eUiFTLoJjEyw6xsUkW8A6Buk6BNr8qVYGkpYJpi/
Lve54UGOhtOjLP6UQOG5E/n9Rw0AeqU8CzYH6vchI2T44r0DNmZIjeFugnGaDhTP
MMIyiP3q76ThOmdrIkDBbxHOAI+0i9sG9QNTWv82JKS9zsMXbZQtVBoMRheircxM
9Z/qPJODca1PgCbSTTiuLSXSiKXOwKtcKaT26BddPNZMHMaTnTHruXcjKlOyfyJa
qYYyM47ZmMgC4x8KdiTEk+S2V9FgjBG/gYnqiLzojLB/z9QG3Gjz+GnJwxM56frP
08xzF2tXDokN2Aqzdo1zgEiAIvE9vSNozez95xRFUjc=
`protect END_PROTECTED
