`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ch8TLXAxvyB4ci67HmTHlIj3ZGtdsby3RhNh2UZ5yOV10uhxCMIk+QGfd/XYwBKt
Rfqb3R1rRYlKKNfo2bKCwxnKxV5UtLcsxBj96yq2gNW4Rf/Z+s4h98JmoqilBh9I
+tCSeXdL9hOsuKWDL63Ip2UTa6F7q5XZo3XKclalLEEJ4ReJ4zViFvITG8Ibtz1K
FaXypVLy/zZaPpLaPl6zZDV94HUm3GAn8CuYZ5XpuumaWE88y0cyVOeBSedjYRcq
4ooBbL6KPvhmE2HjCoF4jxGEQJZKBFN27A2cRc213f+Z06YDlo6PkMDCQ1dJhs6+
XUTByC4wabjGLjttfw5pdrjBrMcH1zpL1hdlYfrRFyo8wPAylmcQRH/tD4nVp+9/
PzAUj/I+vT5OE3KYk9WVry80XYlplOEO5KZa2SR/ree6ToaHrJBghBdUHdLH0IP3
wVsGsiimODows1ZAqoYlZtwfQDoamAGu6ItTz1J2iQwbFGFHhyq33FPuigI34YHy
gw7tlpTC3K6dvrZZ6ZbE05kU+dES3MVzZP5QM2+MgSOu7C74zbcNcOavMEKfEar/
c9r8q7I4KIxJklmowBgNVq5+p//yCevVQXbDuCrpUV7l2vABNjtk9Y+J9D0cXk2z
kpShSkWnB9Uun8LUXSg+naFvkZ24FcvaW5gQRgFDDF6t6DZSDb8+qqXYeGuV0sJK
8Q9CVex5+R4S57jDtk1tFgsABHCwabRoPzMpPa/EK0X4gI5SC4WThmrt6UOLIphE
FevCywY8+rtjHQMxIYgLgzfpynZ1cnBgqvnzg3D7G0UIuWXeDbS52F1DFrjgBYc4
kyMpHd0MrLHRdSzkIw0M8+P9MhUuZhAVJBPf8TqcOgK6TN/WpNt3bbQ59QtEMxZ6
drcX3soPeWb8BgypiNkMwDyJr+h3ehHT5mpwcq3hFG/f+9tj64I+3fCawK+bj0K/
XLev7aSW9u3TTg0IqzyTA2TnUvhA6tVG5d+F4dtz6J74YwBEHpzHhq+aKGRmBCC3
3lio+gPIr1T6zZb1YYStZDxLsGAf50xe/4UL03z8oiWSAigKzeFNnTGQdnbcRQXz
Tu4GbsfHBebRbGud4jxea32eVXc8vHNtsQJk+5fnb/zphy4Cl9xfWjcIHW0s7fTo
LlCA0fa8Noc66L0hseKXcQPN2Jqv4r50Ow6qx3J9k+1ecAhXki5Bcgyli0my+mTJ
eis8PodenA44/ea5Rd3NjnCiHXty6w+u0v6Zo/aAzuqqvtzw7ZgywRilcBUM8ruB
E1hl3diM53NoYTw0Gr5nqiX3AS+0ufUs2r45ZjCh3qEsI8WM7eJb1wssfFVMNB2n
Z6ST3YxkXaj9XSRleXbYdE9KdhBw7E+Uvk5ejv3wJC8U/T0vJKw4M0Z1l9pGPbUB
9nnxNKa7jfzqCKoy5lvN6pUFNp9igOPTA9umiJWnPxVnp8OBBEIWrUp4+KtMtLcW
gsV1Dnk1KpS6lc/IMAsIHR9sRugn7sFWahIuS24vGndEmt1a7JiXLVTilbF2lGIu
/+CBtwJ1HXjmZe/167LJ3WROAdJU1Mc/nv+Y6JzA0J+k0wAp8XrD32opNc+jdfnQ
dqhSJNXCxG6BvmsXugVosmaSei4agdeJncg8+/CkEjMP8qOvWjCrJ4T1VTqd5hl2
JrFwTpTlgsz1FoeHXdOzxK61YiVYUmrt6gsdJtFhzIUmeonErwJcmp1VU0R6tty9
RFZJ+oWOMCYyoZYKfcAP7ZJCjVpf2w/yxb7O3xs2Y44pXo64OL1ycXszCJD5lhEl
H8Xs3VapXAVXT0bgQUMu8nYX21DJPBjwxAuiIx1qJ4ZUN3rfkch2aOg+JrLWW13R
qnb+xFHdAxzx0UNjNtog/RgraGfUFJYDmeM3zE68WBu6OM/4o0r9WC1fDIiykiVi
Rz+C9E8Z/QUqLSJb1wVf0Q==
`protect END_PROTECTED
