`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tht0iGSW5eXs/9IL+M8f+Dy9207P1ZalvqPM2IhnhBS2x6nZJORwKl80sIQdDMNo
l1zDXkJiqtQTUrWbgSLkKwBnbXZE5fLGw4w8qtwGwSqsrUE0+YYjqfqJXKYnhxRe
nw68V9lcIMiwoz/VIz05QvGNB1zT9WSBVmYhg+1sO1b6iXfZ0Q/uKOdbuHw84RA3
ddIk6kE/Wsy5MDRE4mWsAEPX3H73ZFyEoXFrcQxhJCsk77fJS9CDAVOHDM4Oqxse
WejT1R4Vn3xTP4zd1eaIDiU0n6riQRkc/Jn6FqyLUsfJOo58dWoENmz8Ivnv6xE4
DyRODNb8z1BXAwVrGY+mbvcgxdVilmQu+U+dcDaNR7/ItWUdDo3s64YnKfXjE4Nc
2tzF5OhHomygQAg6LR1rDQmCiiUjk5epUcjm4rJSoOxIEY82PmtspbK6zla6mcPx
q6hr/ad8huLp9IlEEYo+gch6uKHVwYoYc5Km+ButBwKfA9nlq2Yf8osr5KNgXdYi
UIvQH5elT7G6Ve5ofmmISm/0GZx/kP7ftoP6/tlTXAHRaaJnENfHJ0rErLvZiKiy
Cq5LGIRsZL0YV2TeltH3NvmChkWWH/ZQZq7gkK4zoVY17xnrMkmWHHr12vOVGFNK
Ob4lHaaKCRZ91my/db7tWhJ3ZEiIKF9iotXPZmH0+9YYUyqt5fJecX8dIl3rk9gU
wQHY2aI4fbhGD+jPDY79uQxhWLFvA4+KPoOg7fjgUnIUEyGT1FwuQZxBbIVoVT7Z
tly+qsteYHHq+FZti20zPv6ZLHLL42sUCgvp+5Ri6j2Ud6M0pQsHgXs+VWTDFA5e
kFTLLb5ksG4uJFxy/ajiZWLoPB+p5I5Zn+kdyqTUNtZnkHhAbdv+j2wT6bXtgXnM
8qRoxqM/pDrYxpt9yZe1c4DSNBJE4acOreraW1wKeWsybUKV51BetGAxZks8p0++
1xjsEEn55miuW+YrYZprO0DcjstIeplAxLjJa6oCsMbCJk56nq+futrA1/9bkOwK
SBRa2tnNj3hdWbsUCqB/rp5q4TS47DwZkj0bWGRevPM=
`protect END_PROTECTED
