`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z9ZvDSAS7tQSz5tpjPW+NeAMOzBovQLVfenjGNr2+BDcIIcmARL1I1G+4q50TRKi
i091L2HLT/F9DVRTUSiMMhr4+ka89prXb3Sf1oSmZr7vIhg9ayFXW9wlfgUASdmu
op3hwWpoqnZo57O2qvdLCqutV9E8KZDfpV4JqrVh0C5+Bat+/Z5yHp9uVCLp5WRb
IM8VsybDiC30cfBnmAqkOaai7rJAxxBcCqV+2EiNgBKXplDaFXhmZvik8FQBPDGc
L8Y8aj3W0VclWCR6Ozvp3WNi5A04DehGDOApNLZJNzBBPN8HxoTlkkRLOG1PtIVf
bH4TxXEPBUvrRBsoBB6bfFJ9VD8vDsahKboCfYeIL39685t+MperaC+vP7/Fuau6
ouzoGDag2rez3AenvNQr+0LtX6xmKFXS8qtbDLaNaxnJWB6Z7vT7w/OtaOAdfdWw
3PZilZOIh2iGOdouQezxC+yAWt9urrs+9j3s8L9Tv7lfubIfwfHTnmPdK7cumJny
QCQn93OCiKzYA7xyAFJkh0ZhuvD6S6RYj1Z2wIztOEbP8wV6tmBq9xmrXCQ6givp
VM+x0ShJDv6myKgpAOfF/EiIFZAzb0SWt/hivFzPSAGVOWryWuzR3ULo9AxRreQY
I7gYWyw46RViT+biSDOghVfIIxQGzmnNPAY5ViG2r3Y=
`protect END_PROTECTED
