`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bz/siTRVof45wtStCUCab8SDH0UMymSLTwgV3atp/7XwHvPErKh7APAmJDASRogM
bIx6B5eNbSxib0CYPHpdQLVa/HIda57II699y2xUP7VBxR1LRf/EdR4E+K4WgKPV
yPwtcjT0e8+m0eZoI9cf62Tivz/284XJnRvzRhP5RX2djssO1XiN61/Iq/ZO/c9b
ZUHJfoC25T0v32RgQ5pyNdisdLpsxPitObxDEjNi3k63Mc0F/TMzxDpLCXk5qtVt
XyW0QHdS8cnV8N91/0F1ecrOBb1OKVhzn/ji66ENvcTa78olg/fiuMfPELlW5Xe7
13vbet/fTrqQEPC8rBi/6Xf9JnAYHIVWjQq+/SnZkn0YnbmEQVVs2RBwPZCtz3FH
va3Grn31PYM7l1uk1CyrXe+ttkeeYrUNrOqmKWbvgZ3dlBup/kp/0SZtbOXRQtiO
tRj0r73IVh2xQaT8pId3IFcMdZubsOAfc4YUpD/zlkfiVzqU8+3A9h26bP2DGKHu
`protect END_PROTECTED
