`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hvup6vdQ01YjrWXvBYawjmRpMtXBsqeOhk3NTpWHp2MmPJe1QTvxEmzI1TGhjFtP
3bAvS4MD5QGWCbX3upAFhw0ri5o3XBw5FUoQ89th2vZMWhdAsmQohzCBP8ngxh2X
vCzvav04bOPKdhZL1/qlWoNu6lzBL2es/qEJiu1ZU4kquim3+QQtmoklrauR89la
ZdyjgN8gX96laOegNLHi9G2DBqjlBTuyLTHMamP7Z9V+9C2rUNk3qG+7mVN/vC/p
gy366BHzGhgUBJVINJHzZ3/HybfRXguPQ15OSrf2GjRc6xfEyOVMXfQyvLxVrlDl
Cc5ndicu31MLndTAEvdBvLomr6spSz0u8HL2ZXMSVni65KNUoKFCkj2LT1BRh6mj
I6FDqlVWq8bqwAIzkC3h4u112xX8YVJurcbpv3Wf1x9zJYw6mCHMBpAEW5JsU2H2
cPW2I8BqxmKfSmgduv1sCG1EhvpH6lJw+N684pr7E9m+EKSkQdSobRiVan+E5wAt
3K4rRj46WnjLyM+WnpyimAs6S54k6TQc7X9EIP8P9xPrEFFfZLzZMvgrTaXXYf+V
jZtXZ0p9m7RGQtdHazLNjDG5ncBOIkxpnKn39EJUvzktDaiHhDxn0Vnc7eycOdpN
shoS6CEXbglysWyd84VXwgRLwb8rusYzsLfxElc9NVT+Um11/152bnvHH4UfqRrU
kaufsq5wmysEnagHtozmQ4t1te/PKPrNioSeo73vuqyflu5UvbvTiwRnVjKbexej
v7Pc/vQpWcTVVw43ulZK8RH1mq32sbcnuXPOSz9w7kZbPH+ARST6lQNbY5XDj5qy
nZvuZHDMa5Fb/rpZ+axtAsrBbStcQgHwdNG3+kYyKe7mGa82/gUf3axnYwIaHubc
UQchkq1rEethsJnHgVG7oN6vSSIjC72XbwHxGKPsPOhVBy8xVz+dqCOjPyQa11iH
lBlZJfw1hz1XOi/PlF7rPX43AJTvReNdRlsal/pN6xdprkMRA41N1hosw2rz9ZdK
RqsNOLWpSIeEE0jwLpOTvA==
`protect END_PROTECTED
