`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WvwgD+VtrSclFc8X9gdKAM2FV6C1SJcTUM9SbAxjSwyE8yerEJDpDrMvSZc/dIhF
ZOCENnk1m8ZvI7Yz9tJHCfhIaI70GuIyDergU37mYLe+IvrI1aoRTWRHOgZE3WqF
y4jTXfvKVw7ZwHTltkz2mvtpHniHDsAp4eZqYrCwaI7LBjb8l1pqcBhm9MIvvina
4MCe46sYBEVpt15SyyFFS2k5zgfn1/4ZO8OIpyoaU/3F7x7IRNyR7vNCzGYx1kkq
PfFhOX/LORClTaiBPu3njjIGoFrqByyLWsAOjXiji6xeR6U28Djh1gN5+tbtGRzd
JcFmVnb7JWzGD7J780vxtbuUdGILBO+G5/xfJmuapl9iUTQlkHoDvy70kyeKRulH
AGxnxCUbbjZcHvQ3wkIKtjg9FNqv7s26kYwASglxlN7Jq6iZeCZDmOTXRz4uoSLa
NZsTilpStmpgqtyflZe7DrU+xMz13CrREkiLdXg7LCuyDmbVFhz5Hh0kP4GjY/LC
spQhxppHEYtsWTyL36fuEjdpMasHL+BRfWP4P/f6rb8Ur9PUYNcRCFkwtf/KyhO6
TUOhXDMDwXLd7vZXrGWIx9nio9XU9P2jUd8rdgP21H5eS6WxLU1M8Y5G5QNeqiAU
yUnLimnDDBa3MkK/G45wROJdlRzJIMppR/fcJ5SZnnEHMikl5mZC1F1XuMHLKSaT
rGPHnI7JwTmqK8qEFLBrXgBPfTbxq3M6Far1FEzrpkGZ28X6QCt9KcQmURxwwYDh
qkxGiowDZV1q4yuxCMUEy9IHiP9fIJqpnZqWYtPPE2HhRcKhwGJWDAAQyN3dsNR7
tkbSTu/OciQ0R1n1PIJI3mt8XhpFoAaMO77K1Cp/7IcnfJ5ImIpuRNpa55KmLElo
cKfb+g7H5SY6pjHsu4iCR7/wQ5qIO9Yppi3vn4Fut4QJcdjuRUeEv332Tr28WSML
K+JwVtJFYY7qXOhavNF+lwzkkvOzGnXslbts2cZX6x1IF3I9jTRV5EndQS2ppAcR
UA3yelTa/CAb9ai1qd67XK0e7YHXCgqAME3GnOI0ZEyicx8Qdl+I8RBL3UWvHeRd
gVJlxiPdxoa5usAwcmLrO5qNFFtGm+b1A/bdv19R8TFx6hAu1fwJS41/Qhexl2go
HDIdsC8g3oym15bDKcJDKMBAE819q6jdXyPvcnzbBnbEG46Ut5fautB8vpffps1T
MoheX3tLDLCioh46icXb9HndnQwBfupPYBaVv5UxHQGHqTfpjgSlG/6F6PIGttdv
TUBD0QpA6SqhrxmAwjeTc2YmzqDB7fekgQYqcUVfqpFrBsAvJtwErLjapzx4QZST
OSANSqMjyYY3lnsb3Nl7sFRg21PTXoVDv/saKO7YNjM82qI+mnZzmOAjLyA0pvv0
Nskbsqap5rLriEmIkoNvg7ZIzvkPmB4JHGyyB75PvrjgcM+4oScu+p+PAXBraKJv
ZbbzfehbvY21s7JQGnYy3Ewjv0j9Payq9OZgsff/0p1J0Kk9imvN8vWuyaeCpA7F
YrkNgOeene+Xa4IkwxWtp7RA/VG4pp+36bTcK3xQV82OMdvayOT9IRMpnSJ6w1Ss
x1vj8MVQeGmly+X73bxafIRRngEDRmuxES6qPp03SHKO3sI8rHoziISLCB/afie6
n54iKarnp6wM7wpP8peRm7yTltB1Kj+d/RIenDSKqEHZvq0AyQQxgeCFMneF7jRI
4Uyvjp0gX9f00C+L9i2NOsJiCn7IXFxyrJ8x+cTkq0fNfbIJZl2UXV7SQN0+UsRa
xmEFR1B+FB3qyhirHENGZl+AcQDITRZxY/klqKrg9kkigU4V1l+hnFPt1Iy2ACUR
iysp+ya9eBApqR0TrMeiBZYsOz/8hiinmliiBdEG8etybt0lAqhJLY5WO7ay2d2C
8lWa/s7jtXomze84IttcBw==
`protect END_PROTECTED
