`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HiHePf1AwMyG+HH6zkmqekce493fPI/JTTHxfu76I3jHsC7At0ySnuJCbS5KJHXD
6XZbTMZFocvCAMoTmcX0omLzYuB6lw24Vqc4032bhTrwIy+baRlfD7yOK6yb2vsz
dvadg4VlsvQc/cE48Skt4k2WPmg43auFt9G6/6appz3oYykhJFoXj3q8zrO55jX6
vZjoDmEIuG5DJBfV/zpXVKXEsparm9YHoiPQlnrpZm8R4FOl0RtSHvcn7rmocPKs
J1CPmoAeCmnjo/lmexiBGIVQgC/v7r8Cxmfe3JQ0bsacETuskPmmhcnq6UcYZ0l7
ekWswNcCZhbiFMOGrzjYdE7EWKoxplQC2eaxWwMWLp6sbSrxG9umAhCVUAdOjW3D
/vzNw1MdpECqcq3piid4yNrK2J3zdNlrNBsK5pGzQPemPhJJau3y2LmJZYmY0kqj
36ejmvf9ofNxo9/rlpSN5OsmbF8BrsGbEhyBiZpIbKt5HWi0RKMgihMecchiQTBa
0Z/ts1XVh8i3FeK9tfcCGjJVHxeIKG7hwQ98K2gpnllJd6MylTJbaCiAoiWAQZfu
w89xYPB2pyVFjOJqlbmxDJraeEOuTK8y+E9g31qgciCllIrr+neWFtyn+S+I/3nk
lwSOWHc1J874OaQGBXnOQ2OMfejJKmCY6z+ADzsrZHEcfcQh7SIygaFrRZXRcoNN
CXNVigzA7ZlbLLuaYw1DNb7SJYuAYLYhZZyxGu6yAKvf3dsNfEy5Mfk5/c6ATLzg
`protect END_PROTECTED
