`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sTZUhJ2FEjYPnTOIRqGt+yqdo8JRJyyrldC3MpfCoPbsOm6KYXsKISKXsTCp2GqV
x6ciUXsKMWBAne+0BsGOhjsT98SPu+d74/KWRzH7OZv1Gs1XfajbBJFud9suv1YS
rxdHFKEfBSTuVBhriMCdiPKC/ctaAAGCLhd+UoSw9rKBc5+8sROfgboFJk7MxRZj
uidM3Ds9oNH/34X51WCGlUCEvz8Nk2kjaYs8WS6Vi8pxJK1XCZ12xnXLM3bZaWAy
yOZjFXJ6UVdyn6GgFbyMh/i2onfRf6GT0CxusZKFsIwR8rWOllSlJyrrQgbCfDEo
Gg3uarNA41GAf9i9c2uI1/XldDoGgvcQO65usZiGkHGyP1nRovs8o84baQ4e6s0w
rBGbThBF1jPCtYJf6xiTSSGm/cb9YU+GuFzkxx14KXPktkemfC9gWVTRVYWdNJJ9
W06arW+YcSuRFsy7SiBYgprdQ10rG782mcqkEfZL9BB/ptr+Gj2JBRAHxbBTARIR
lIHoQpBX8AYv9yV+FoJHwr9GT3Df8HveY76/Ix/Eamg0Clw5iAlf0npBc6gdDqU1
yZuntnR5jGbWqsmL7RHEd0M+FF/S42goqye02ouJQ2D2aIVOySCJ/cSlkGHLL/sF
DMeVRwV9qIoyMolrnzCv2wl9zMUpmrQIXxDP5Ru7tkzeehc66a94dNJo0XTko+nU
8dLI9Z3Ri/gXdpkcj5qI8tSNEreY+/Kl8Sw39tWkJfkOxzTay6l/O9G5x+hrs4/S
`protect END_PROTECTED
