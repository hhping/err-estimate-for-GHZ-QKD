`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ihJmtXakPwP7TS5pHbgDqVj90+Vb96rEsk+IEOBMpe5rUShH38CgqqXa5MVnpy+W
FtZ21fJavaTPP4GA1hOQx3/aA6VzIeYmjSmARvxo3qJOgspXfPi9annCERHZ3BjQ
7wmfhWjLOp2oWTCVT3nGo/TBI4YwoTfUaVeibVnQ3DyO2M257OWyvvVd1vHpeBk2
5CzNk39kcsxHMte4VRyT/N9/3awaQE1flqiXHvAER3dSj/Jgwuqmp4JBEqecMRq0
5VHlpHhhaD7cmn6ejj0sAMLKdRt+FT9lIhJMhGmYmMMc9eTdHgvrjPxTp9LKa6GP
pz4F7TxySgB7X76xOiOXTMAaUqtPmCLtl7c2+dFpe4qplx99Mi0LF07rVWgcGPY5
KtTJ/rdpLngQtXBt+xTOJX8FkNQNCedp4oHQ8ZX1u6BQAlCG5ZCXqvIVEMLpJRyH
lf4eM4QlyTApcf7vltzRPgFOOWuRluCcVr4WWcASo802V99zuBjl7Ic+AEvwiJFJ
/qp6AhhG/JYf1SRTloJHoGxqjAq+Z/idVtfw+WuE4VV+TMKp+5ewA8FxPi80w6kr
N/tfMGcooohM705BywxIDg==
`protect END_PROTECTED
