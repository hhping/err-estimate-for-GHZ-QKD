`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EzHQ31NWWH62Ia/l2gnK5u9qTrnD7G9LA7RT2bvbJbItrnHK8ZqKw6gXRo334EoO
o02WjgmK82b2pvqe/E9NCJCp6whjf6eY8p8Med50lpcRY7gaO8i+J6v5d40zS6fl
KzIh4pdl7ByOoupbtcxV/gYTTdsxRygOvhWbVM0Ny1znUi4BGz+dtkgTBeUd+OgF
67LmLh2bg69+bcnze+2SObcuDlQ1IkpUnirzgJT1hbXFsA8tjhHa4qVBTOqcBWlb
+ki0zUHyP8jIL66/odDvmMt9QS+NDTtxPqciWz2zXOJjxgiFlqsZ+HYt7S3uF5wV
2oPHc4kEDThGsDmGJvfceWRrFnSJ5YEJ3sUGFv1JtjHGUzMWQIbyqDer3oLPp2LT
nZPCFw6b0r7fkreTsdNsLOIJp4tV/w6N8n4Fiuss5KFVJ8C7Wdr1vtQQ7hia1Qy3
hcFVu2oLsoUuNbMkFLE1ax8Ry0q3xbxvN4eXFuUTWM0L+nzTU/zbaZig3mGz9CS9
Gk05Ypr41ShjR0/Cz4PugenfLoONeiNMCBu+HuRlFIWdHsEJgTFbgnEB3W4H0zeg
8NigCnfACt06FXtUReigwCQuYAXtWlQ/NZFzAj+qDgpHhuTkCLl6LhIkiquaXqrk
A9KT1a7Ot+x+6/zeoNTNOuzH5LOHgPhw3C1Gw0xywlB5zq8jv9MsNTjtXeHNTJOs
N7xoQWS557NlV+z6DiV8RITI3DBPsOlOm7AWDRq7fxZKFDxfFD9f6H640qZ1iQzy
JdE2xoiql3sxyb9hMkH+cG5a83xqJ9KfAlEwZME99ZzwNc6R0w70B/5V+wct0vND
+lxibvud17wxwd6hzRvGZ3qpkwfIYV9aM6BCEoqNr5TgSoVphCHEy+MddDvy0dUC
PKkk2lcrrnA1htLSw5dJZVJ8Nk1ACVF1UBEyRxObPWy/eV0nb8oKBKYicpOemvnk
n8SWumJ2seEM2+iQ8/RCe5CpXiu79zubecUhGqMm4ytNcPbAcZKnKKSl3ILQ3Xj+
d/xuoOYAznnLJDDe/Q9m5+jscmLlPPub/l3fB6donv+kyELwiOYI00z7FtAsxvrh
lX6wHY0f2O6SUDnMfCs3DwhVywHIGxyBwYaC6adlOE4O4cP4hxbeYo6xnJvEhQAy
Y7yrKC5kLjsVNYwd8fsGInYrh7NKy7QMThqXoiJDF1mCal3ZDU5C6JjBsUzsI+hH
R5pH+23pqL0iOhdjPSHG8eXzbfXQZFBjPcJSWVstqgYTsoMElfQN+MX+B8gfROoU
ZF4X6vHGreEtp9G0Uv8wmxAo5RS1oq4gjRLJIj/Ah/3Lt2qbr+H//+7UAaYhOzHO
Z31i6zvt/S0E4Ymr+jEtkmNTNx/w4g0RGSSsct7oqWRdo5UWBZhtSQ276mywthA0
IFw8+OEqsntuzMofngPiLpfkG8nlKEfxma37vrGfFpP3hOKYr+ujQSbQjU7NZruE
c1Fiw8LueMhj0WgrnA35fbFANFhQCPzySBMUwX5yzYuTNX6rwH/6SSaoyKey8PfG
f+N+2oT0EOWsB23p3kZpaHhJAvF7nBNck0q65C75I4OpJpmEwvAA/C0T8aOebWxB
7D9pWJsQEU5MVsTifjczpJ542bRY0MAYOYjYfWk6kTJgE0uU1FbSVR0H54H+hjYy
3/e8BPoh/VLTk/9TCsP7MORf1UkmRJRIQw52v6tYSWbsFrlnUoHCaG+C+NiycwTJ
TWHBahebmojk0dsHVXKqsuGKqeoDXqrKatkCZCyrS9pz9muSpW+KqqmHEn817dep
SHP2+m12qF4gKjzvWUkwTzqI4uOGPjuiw1xhVtPdJxoWezsuTRwi78KqopTu+r50
+BF4rOajEQqlw29WYKYLOF/F/dVauKlBHflz5j4iy0Z6+nY0SAbYXL/2sa4JaJtt
u8YOwWdTtu21SiOTRxSzN+cFXYW4Q8JPYTRa2F5mgJZR+tR8yo5MIOp5abLUrXx+
ABOlm4MOxAgy/GgKhNoZmOFwUDtIqigR10BncPUJm1WVQV7Yt3bspwOcftGwBm6O
1po0+goYAYRwImQkwML9bHazsgS8BqrRpO3mmMDOJC9EQ9r5XKv8E2ZhbByz+urr
wr09+uZiMs3ErCDTHN9gMah1FYjtssrOPLxJKnFiK8ZJM4fQP8JbMDvyX8sQkGJS
s1hD1kFXbUKeDxREaqsAKRtgMzccROHMYDo0QtFPtmqrTdXU+m9J34G1+KJ0rJuS
wCFhs5NVejbVByzb9AEcTYzSgMUHdXKDrbJp5U/dSM0MmZXOYz8o+C6qR/s/LkRh
jVoIPtGwwgjuhfntFVtMsLUeFikk2dzvytdQwTM4ZF/PJkie91AYFn2YXfilBdhX
NEJdyOQkze7IwpuGxSia7ABEkcT9RdAAnpKAdRw8VomJ7BjAUP5CwUZahHAcxJhX
vN8WkcawS0LKGxBt3XThaWMi79JivZE+6kXDoMA8f+GNTrwM1YB+Kk8PrtgjFL9c
kHxYoXM98LH2mAZxQ++a3Ty/AwlDU41JHmtlZAoBjtHEYHW6JmvMkYsgvTB8azkq
Pb7vZJlyL+D/eLkeRN9u100F68S/oD2++NbUw9ErIF64BzdFrxGfUul4W97wP3WO
PwWsVRMAl34UF8szAyXlZUmNG3fwF2yN15/RvZKTRo8NP/K7SOKOTl93hrtvJCfX
9TuUk9Qy8pS8W8Ru388NUa8emEmWPwbGjNSk7b4+uvS0Ym7gB7mKMWrgFjgqvl0D
MXSpF2mvGwyONxLmPAgPxK+7eRMtMFD3xLY4r0H3ZTXjCXASz8737EfO9b9xTL2L
+zViqEooZKwFaQ5XCKPWWvmUtwqDebONu7dtETPn+V3ZYKplhahMxqu2F3098ApR
QpKGGPxURmeAKBZ06BCqsA8f+e7DlXLUdfwIl0wJWOyaGkxXju5UCemmLh7S13tZ
O1JMbMm3rmGQN1v9Ytn9ugid8yazIrvgJGocS1LP6SbNiqaQBRyhWgy/cuhLCvad
bTlv/Toxf0ejXd8/Z6LRa+Y5tzhxp5mNfqmfPWgNiVmDUFI2nxRUo2hqto4Nvxnj
tkDKY5DfNMjrdVRrqgmX3JZR3f38OkZH+oj4JbN7QGuBeLAT7/xxS9NmCYGP0oS1
txRwxYSNJxKIAz6uR57F2Hk8O5qT+mDA1f+PQrFqhMNfM3LkX5jzbXwvGo8mK1XY
AcznhjlFMp/kLdtQ3uADywkRtXPwZ4lgOMEB7+uF9Ml7FhOZOyi5KzYToMJ5l/HW
ZP2JjWAkcjlyy/6pWN3ZCX9rgLrDezgzSGSzbRsRkiy70ecEaQH8qDvnuGXe8vHT
zlpPTUaXARUEW8hkrxw4ErTiaAKX1EJInoXiUtsDLUocLf/pp5Bff4A4kUlNl2V6
geTyMF5zV8KEJo/zXKaio5xpuv3kAk9m0AgD1+hmLbpGIFVjI7iSEG+ejIfphfNd
Bkt1QqSR+2z9pUDBmmJUML7IIn+vJ1xZILnHJPDEd15y69JBvpw1GW/YqRM9URIg
LA4ThvtT3ZbynpgugwHHtAtnuKr66CCZivl8+j3L4K5HRyn+6B1rj8pACc/624TA
3CgboT9XX+Cw5JbJIPaLFXzAYIZukQCc7SP9PgbHdhVqsuBNiswsswmCUDHMwwFD
dWzSL+kh0k4K5KV8YWyyhq6A7l7GWy5SB4JzZf1A2PxU2o/85dUMkg1NkAwT7c1U
xpVD6lqkC4SXFiWFdWSKXfOTikAmNHs/reEcafK1QSpTHcN/enudo0dK6gzMnjul
leBFqefoO1oWe/Cj1vq0kY3e/HSyg9GU/JIIaVoRqf+fBBZ3UvfYGoIBSduDppKX
iVV+Vx5BiecxmvDGyNPw05ay6id7kDvP9i6TuIsufPlUTJ+9FPmgWsaeH3Jv4Nc8
sEU2Ny/uzVb/eT0nXaJy90ihEmS4GIbLQgwQtIz0xFezOeil67Y1sxEIAlgyJ2RE
dATt60HI92N9eQJ2n+DxKiZZXp7Qb2ygX+GesIwv+/4t8us2k1NA+nPBB8shD61d
bN+EBT316wVtrIk+ZB2XJLCouZZJca26Gm3ENlCvPfSfPLiZ2dfEC9EpUiUBUuUG
HgL+VLn8jVrNuROGnPlMxByo5TNM+VsiKs+USQc4RZgQV2Y7iKBHmukbnvkkw+DD
3Oy/oe3GV4d7oeqwfvQp7n500/BJzKsWn12obyioTWwD4f46l4BE9el0/904z1n2
SZhlr3S1r9z+Rzhu+jKAJNWZqCf3Rr2qR1hxSxgVMtgR6Zm8XcIYHkL2V1lzyhBk
vukBlBadhOUh8exUWPAVN//DiZzLmaSYqszLuhQd7kA=
`protect END_PROTECTED
