`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
psT8jmzOEFIaw2cOOS7kDVSSXRde3MSCPvYMkDMECFA7nYc6gbp+9tcXHAj4IEEc
HTrFc1t1CxqgyYHJDlqulIuP1YfTXQr/wYWGqLaDm10fJYvKy0wHstrc/0aO0OUO
X9XRCMKzImOSk+JdE2puiLo0vHZUUivluLf+F1wobbOmHxiLsP3XSrcLJn4qybas
Dq5qiwPjknKrrujKx5bUTwj/mEg48DmvqDssevwh793l9XFRtx0xkisDkr6pfFKP
smPgVrMFl1BJwCtm9n1F3H9LFLsM1Od8yHbytdjbwtVhhi8q1H5SW4To15KJmI5o
NAbTzmrYeT5PoMBq1QsYQpBuVgb4UjOLEkXodCp1EZXzTBxU7IG0F8o6mqCP0TMv
NWD2d4Y3eMSpfqCClrU6NBo5OvQW0KnphLmCDgKOgzj7TY8wlnK0ACD1/KERDU0s
slrhDzJFTnLKbr7xqcLn14vXBay1Ov5IBkick2IZ7gJ86mNrUc8PApyDuIRN8Poh
p+ImqA5V7cl68LCSqPJKkL9hCayhNyzaBrYcyT9ftQ37UEjb2IGtvhrALGkQy6o8
kAlpBuW3u8Pvo0xoLP4TDd/GbSXcEgkbg//EvfxPl8cSdrkgc15M6CdeAguU+VZk
OLy6A9dAgTqy52wIz0HfcTKL5gQxfGl1TEahWW45z5OFZEqMG2rAGxVtUd6nolTX
rG7q4D5boOmF4Up+hXV4MNbJ2H4NC+lfHq5UC49t43U=
`protect END_PROTECTED
