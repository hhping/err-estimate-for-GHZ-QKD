`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pSBhPfUICslwho2Hn5mr0MiboS+8WXAI2RzCSDMgsqh+VvWy2sSVkqUhvoNvDI0q
sVquPTQdxbdow6rSrF+SpUaQMv8FBrfMr/TA4SSBsN275zPmPQRUCdigsPN87LTQ
lhqMlCIzvtxcuZchdnmFq6FN6jOhG5u+BbIP35aihjtrfm/iifV2IJqWOJNv+vJe
Yv7lZEuDnQbF48LfQj4ZzVdYW5VmPrPtWtQdlZgq+VuH2X5g1zaD36YKFRtUJrMP
EBGZh27sWhxkjdT+eMR3iIwqYhIBt5NY/TF2Ry3ySA4xRUojQw+pMBag4QkyGZLz
yg4vosGx3L8u3JDLAytbj5ycNUcjUWkRjEgpjKAuvGaHbAS8e0OCHXbMG6fjvQwn
Up0R0Yw3KA2i8cOEV73/PcW7G9QvvObWEDSTfLHu0AMX/IOPC/SW4aOTEREMV4OQ
fmDohE+HACgz9e3bjvyjJZq65BEV/ei/WgwPdtH797A6ab0b3lKS6PWZ0lhzsvbY
m8agXbhMJ5xwY7zSnYYHvDEM7vfaXmSVn54yyRbOucOUR121yBThKCEWNYaYCzDf
SYI+Jb4XNkt3IHY/EQgOKaiK2dvWnHfjJUijjSQ5kFNLwoqeQS1lGgF8k9t6pqoy
XWWYkT19BrL5OcFWN2h3UV9W6JArWk9B8KrvhhIQs68yzblq0H7Rm4qZ3OkDDbPo
aCO+0VFgrBFz4YEStp+ZW11j9WqylpWvBZQ7s3StH86wQGt3rUR5FUBxZ22LUjYr
lPyu+e3R6gHPpDI+Bd7UUXcxOlROBgHmE/YuFVvkg/j5VJsSK6tfsHWSrJK1E341
LGjjVxx1JN4/h2LKEquT1fm0MhSUx95fGeO6IhDnK3sqBQpQ1o5PCYVVqpLs9vjX
1EGGEGYTR6TOxMGAzUK3RpjlFnwfUgVFjLVUrAUD7zYPyitnPoeKzUl2w1IT3N+b
uVeVv5gR1DW0jNlngfZPFhiIWZPX+9V6iWbYxlSE+OdUUvv5cT7gfX/OZb1gfnSx
W+pYGeDQUq5v5idB4zVqvA9la0KA/KlNf2Cc3dXHHtOrl5xELw/RfNjNBdozlc46
QjFYO/yOwu2S5vMZG8JiwhbOMYsppYjLK4T1yiHMd9bG/VaRZwyiJa8rUqiq8G6y
XulFQcN4XMGRRTgfodarcWvsG7qR2TUyJ1jaZYTbWT5i+SpxjD0d3OrJUKAc58NR
Vl7FGyaVgOkByJ4LY7Yk5E4lYCN9iEv+padNf1mvNKHgGi/gjHxGpA9QGeJOix8r
BpTognNfXkeUdbf6D6UHHZKAtfqnhf91x+hVjXpa/o2jhzatj7idn0DdmESUZsVr
XTflhqtMYKBeDSfGv02tthVz81KpxA8Nkik1l/NjJ0Zf1kxgX6ymv0Q5uS9D5op2
Sfn2Hgqbxw4JWwlqtScIEz8Eubi0O2pzguQendfFwHoW/KScMQUs9RinRgU5A/+V
EfUq4LWW5CShAIhv+E/BY+mTSuXHY8DffVw5YdSeutlOfkZYXqlqeLsZJutYTxMD
0wdyfRc9J/3zR0eZcepey0WQ311mDyPGPmbmRvVW8zDeEWSwS8h+2mPAfra9rmCI
6YxbcmVyNaF5C3tPP22LnbrI3zqK9wBVg+ImcB8pR06biLuYOQkrgZCnBJmiRyf5
KxEpGUSj3JVftfCkZNGE1N5U7YQtG3DXYSxvLuQp/huAiJZ9AXvj8qHTuYlPHRr1
f1Kay5NzWRyYffWPf3LiNk4WXnXUYeOIK823yXhwBoZ547/1dCzmVqNdAO+Vf+1Q
gWlnkYAbXIqWaUKrNqR1jigbK1QP6wr3yEtsD5HbprlIe0sIpvycwj5f3eWPb2Zf
7kO8Htq0J2OFVH3s55TQdgx/ww4z/e5PGQCvp5ojM0U5NeL0Y75OlNq8gywtF56E
`protect END_PROTECTED
