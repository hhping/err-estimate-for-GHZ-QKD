`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lb0iJ0sWpsMJ21A6tK6BKRqsn+alpbWpNLY2Kj5mGdWiBqzIRkZ/ScCJ0COwVqaU
R4ryJWKh6GkHnxtdYRjp0MQsMH8SeCNwS5GACju7+497/obHc11/x0tQkruFRYTL
nyOFK1v0LlT3/f3G6dwUBgpF0DY2dP96FdHjFiUrvURfG+79FobdMwEABUUOiciB
W+TdGD7Rj5cQcjzMiy33KrA3a7mghYR3bMuj6ffAgrsVnN/dH/NJpBqeV9EXblWJ
GQhm6/DXJ1O+rLoHfik0yKkYZ8Xz4GW1m/cx3rCJ5jpp7fMR5fKCJ2FbI7ku6AQz
GJu6curd2RKEcd23WT1sn+dT8+v4WhegiM1ey1cZxsLnX4jikcRrwpDZP+Ne29/X
ZoD3+ydl/HZzXrt+V7tzyO0eKnWRIGYn3AM8pMf/9wTPMtYNH5FQvUEo8PuWmy4T
v8bPYb884ujrcA07EQvdWZJkAaCeR8IyglZHY38s/2N2k42N/bXRQK0053CikwOc
HSNIXURUUfkgRgAOorqm0GwUxetN3QPN7i6oI1uDY68=
`protect END_PROTECTED
