`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2S6jmr4vInf+dDLb+JgTmtaZ+pJcKggIOPZrcFYVlqDJ5vgvcou+bogx4F/jVL7M
O23NEF+NU9GgN4pg1H/UJrEVZp9HNptY0/ZDWCUQ63X5xULW8WXsdv9O0tCEX6QG
JA645y0joYegzZPHneCFY6eZyGf2d/nYBZ/7BxK3KnyheRTqma1FR71vd9y92o2O
V52s6/fnVQJd5Kw+uVFqHXNEPI8SgDNvAEfhFMYrJ1DMvs0j4o3l0SIlRKCcaW4M
V2P/JPHgd5Hmcnyjga+psDG659q5DqKZrKXVyYZVyRb9EBKnnNehadfmReyHfhy6
/RbMufr5tFEtvb2uVwHJgPXX4aBi7ooeM0KjTA/Ik99TRNyWaV9dk/9h7mDtbOqx
bm6gX1kU5EBxS+vsv/Qgg8+LirJpRRMTIzdOv2202GsYRakqRF6Eqan1odkUo3Ku
Rguc8NH+LXmy1J5vJPSfby5CxdSeHG+lerwT1yX2i52f6FKD7zALVmnoM+drDOyy
qkuZp0Wn1P7Z7w7aRvfsg6pB2TT5RzHsd7TKZxa2NA8lERAAiLMEyBOFa1iv5PQQ
Q+1nqLECFRjXbJJbhMizAnKtRmwLfSG9rA4HFHSFoLA3Tqvlh5p7UoC/aRVtYeSg
zlXqK7p51xsqyVeOERZwMjXjCfEf1fQtP4I1DnkRpGZD+kXeEtWA1Lsh5waq5jO6
SjIhsf6cH9WCwk9gU+p5VpM4ZuKJnRbIEdHN+kLxzhCx1Tj8MgyiWJLW3MwJtsFN
OU00av+gd6L8SC7CYhJuNkntuv+aojwqrQvwSqX7kEEFtQ0XONX2y7ndUzNgxL+s
v/jlTKbIOA085n9hT+ldKh+9v24ihVZp5bahlHjKXfmKIu1gI+1K8OFXRwFkcVOw
Wj2/kMetH+Os2+YzquXNcVEvis4jRgkUJaV+gNsA8ySVygxvCmTgfLBRWKbcxBDV
M2hSBQpwSGoMvYETSSbOtkKuBXT/lxlyvzgFkNUmQ6G/ICFq4oLvArDc/QLYcoD/
yvnbXg8jb0ER59Bo8cyDe/CwBUJCHM6y4GW812qEpgNEFIXUzekkZcO9qr1j9nUP
H7TVXChNgEhAPxE3hGNOyTBV47vbtKSVDsvOaZQMggggmBYj049ZILoW6mX6NIcT
VAODjTCdqUA5wFcJmiZCjIvk2mGHEIqFlu5EVvs2+cG8tJlRmjzRlUMZHwnsjYGb
bnZBd6Z58SR74H3ViEBTzDKgLowh/JSNgs+mV4SY2Z+5hHO4N/+w7OO7WA+5FD8/
iuAuSRM1Pm/0Eb6Te2x5ErJNPdMEKwDQxncJToFZ2cMcIy8E4vIwaIMqIJ5VMJmA
LP+xE2/XGDhY6oEogC85iA==
`protect END_PROTECTED
