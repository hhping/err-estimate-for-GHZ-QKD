`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2QVvWFyzY6Nkk8Dc6FScLjIZMvnqdNilcX4iaHAmiAzJg9LSryIHpEQCrgo4I/mD
BTHcFoaQpC7P13VeRMzczznZmINRM/0xE9jmVWs0s5+XPc8QeDe2v4qL+Lh4pDkp
uLNB3wcgo2+JaH2JfCFk56oMb9C0Qqo0uc/M1jCvTUD9GhopX1xpC9q3HcQcXHfH
9ftn+kXecQitXD4OalM5npGatfvo9GbuYp4KszyivvswAVo+cgTeZcnYaOzGBdea
G5IhtrOhLJuwiLNvwi+x4fnybhuj/Chykk0P/5L98ZbKsU3gnRuiUIgiZIFWtzB3
gOnYcCdwCSZ8bRv25v1d8k7kdkalB99dMtOmdMYVNcTJTFSq7oba/CcUeQ7m4MNy
lxj2OmnXbaMC6YYPGVjYFWofDCEMCXeCyEbcgAg+KmCRm8dJdqN//ZYs5ZosUPEo
fYOEdLAlJ01m5vMXebhKEO6Xy1OJczwIfOgbzNHSu+Qv7As547lrVQIplhW9yAk6
Eqjd5UysW3pjd1Zfs2AUIW44I4YzXWU2LUo11AfS/nldoiDN76HD5usWQc1jczgg
xXNyR+oDMbBq5SUDGDuzNLFOcoJrxk8KFMfddyG/MFoYiNhpj+BQ9wjgiES699Gg
vBDAnVp+/bXX7dHGe/c/G3N14phCjIEyJizqOKRoVgxpsczAZRPzJmzCjeCzdUdZ
5SxBHawg9X0YTDjgt5ntpvx01dNwxoP6dawwLB4mmwN0K/BueTgvu7YU1behOP/r
mLghNY37NP/66ku5tPMVi6V/AYiaUUw79aJ8rVMUKFWIZy3HKEz3ZXuY4U2E6Te0
TFMPNgml7QQOjN/mChju4K5Kxqd0gb+PEsWL/bbAuoezeZrdvQdApoL/Paa9AHSz
a2Tmbwv/EdGrDtyKfC8ks9uSVWizCdH5bUchQ76QLJ/vCb5z3tydQOBCiQa40B+o
SN3kK6QwlkoTHvwFc6Fddl2BXWvA9X0R6PdDDygFKvRy31FuNJIGzfJFQrBCCBN/
/ooPAc4RfLiRNL/VaegAtN5oT/auU0x1WEXJTBIWdsfjUL2bjno74pF0Tr2MBVem
7sJ1RTeifLRjB9LathCNNSJdQd/G8Ll7PBhV6DCU6RE=
`protect END_PROTECTED
