`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
chHgQJ6h0hbJ5jyKQTgbbHTZ430AtzQbsNAtt5iRG35jKMQW1Smyg74XmTAaRzc7
+mw5tTCEAhwdeRLUkmQBuNCpsanNr7/IGPNL4fmrSRk+r9aGhbqEiyRvQn7UlwBP
rU7+DTzhzf8AuWPZx32S3fSAgWW5cVP9xE7oqwrKZWI9t/cJl1sJKoeVGMB8AUiU
UCSOacl7X6Z1G9d2ORw4/L+piCiCHDFWgMUEdIMHgkpp3RMrRlQ+TPW35ESEfYCD
T38n0NtPfD2qwdeFFobXHWcol4c1SweJz/2tJmIub4w71DpiCoIvkYsWbm7UA88Q
H/Ux1eI7ghNAFOijHAB4KIaNTZ1y2fD0HQ4I70HWtkqFwEKBtE4QCb6MsWxYuI8Z
etrCG5/cBV6az0A0W77fdswP1JNvIZUbRgIM9EGhU5q2uBWkpC+XEvXGkQwG6FJK
bARJ7uYL3wWQHavCOeZIa7CSy1beRjoYrdHmt5Klk96eFZthj/SMXEai2rcyzglT
qk0rUycY/zgRDpCNVz9j+6L8wTXbS6awQXeu7LsljOcsDa4aPJkZ/dW36jGYdytC
pvkIXh1hX4paIy2/GhNQaudIw3Ccx6j1KRzwrUJb9h5SbAZW2SRRb2kR/DwPFtIg
QfH2xkc6CWV8RxvRSJIDyMgSQ1mFfaeM9yMlPXT6K1EKeEMDs0AQNHKnZMQxkxX4
YKVKR37jCv2zwBHFAYtCAQ6+T+RFzUA3V4ablpEeA1k=
`protect END_PROTECTED
