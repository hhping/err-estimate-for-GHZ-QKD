`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2vLaKEExuKY2hutXlQoG1YSrllU8VEVBIUmeDINuf+fno6Obftrj2qAtXJ8XHHPm
g7lPRReo49fOPo/d5YXyFpxDrx4I77TcrLpGU0kr89vo+ge39bCXg4hXMFZejCGo
S67YAF6Nx7FyXq6uFuztpy6YeqOiKkAkK88Cv+cyoIJsN1J6opr9X0wuTpw3/100
etYUl84NuCpj8/05TFmp47Qz1mtPCqv5KJbUwvzP6G1dvwEHx8ZYC55ngZ5BI2o1
z960tRCveSCVZoW2mGjMAlFKb8vV7jeLsoGdRfWSBtD9PGdBuFjj562OzLWAS7c7
LsE4CJteCuF5LohOSiZgsmhS2+s1gq5ewyUzRS9rclzcSnOzhz6E68vaTxU3z9cW
M7annRPJVdvkxsTZBAiDIA==
`protect END_PROTECTED
