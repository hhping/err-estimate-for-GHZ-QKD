`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wTKG+cXEeIlXb0nwbj0W5xRH1FfpFc5gYcZtoYsgt6cu4+qed5Dc8KKtfQ9uyx9+
gr8UGoS5aJIVkxdlC+0hYLKAO8dkX3wSqym5MlLdmLHb9w/XkJzdIdgAMrsgJxsR
iUVpJUdMICENMJa7vq9qoCovPlguYJA4Qs2Pq/7yDjqnFrcpjz/oX0jEjyA23pVe
sK4FNY5KxSPGyacxheZK2C1UBJb6vsT5w4nRG9nc8Zio0jybMA6RdwIefVWErxS2
NXtlzZZCR5CMX79hcavs+3DoWXkPDu5fgCcgv9iNOza8HEovaxWbYRuudEMIZ+bO
rD742DDo8GoXd0w/m5MMu5+sLYrYE4scWRchSF2GSVfCF2nj6jT85/gPEO+Y8TAe
CW+frW2Niaa7pzMTFQybPGIhHPZGN9Q7AiodNbV+Et3/Doo36BnoxTXzgUnA5/kd
gzZ1IA+r7/qcwzn5RVOwvgWd0priAGTY6YhbBJHAR25PQv4tYz2I/MkKq8UNmW2t
8CO9i45XuXerPfOuM8GqpQ==
`protect END_PROTECTED
