`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i+/HYIBo/3001apvJ2DbqNGSG0Nsm8jmHmyPg3/aiyDDdRcOdy5RxxhANISGKAhk
EbEJerv9VRGIKLsgcQLxMD/Y7nvifLqKacCN2LNqJMQN3/RRT1qHVO6J2yVjb6ix
7wERubyFIDP7+Jfp1AwqmggbzC+07ghfdjSaSw62s7Ryo7cxVTQOsqUIZ2Sw55dX
6gRDb7O8VjKLUhfMO2qzIvIvqULNrFdQrj9F4DQcCcEwgVSII2SVlskMMKkl99Al
oLwZRk9r6x83+OiWp/uMoDME3jZnq4bFrhw8ZUFFROWkJgdTXQxQVe2Oe3vbTlTh
Y7mbyM0aBkX6IWmn18yJKLDfsf94FGzlxfIZ/v43pUtZh0fl4JUk5voCg/pAG+ve
pvCk6VUDRXBOsO1a7HgmSrhsegQcl413LzN1ng1E6YI=
`protect END_PROTECTED
