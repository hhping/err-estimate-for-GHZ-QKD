`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d3uu91z7vuySOuwOcik+TKhotcaLIUjPA1WAOopLhFny133KxCcevWTDZFjq8hx1
3XbdIYGBNySLPCBtgGd/fpkJXxt6dorBMkfImKnC+wzW18K1FimztnZwnl77JukH
1a70RqQ1CcJdZY0Zw4qh15KbkV0QZhIhL10gmR57+dOTTqzBbjmIND2giB6m4X2Q
gTuhVwwtT1LDsre4O+vXkABKsU9dXN2Clv8GbB67IiDr4+SX8B3R5y38TcvkCevq
lnZFJjwVO6XhX+KJDmK01sxtgwbjdQVHQX+lcGPXlS3T/E6jd3uQCz51Fwam8ukK
zBD1YSt8xsD0H9msKWTwv9oFzKaM+FBJgLvr0ShrM1fI3CIgt/DTVVo0j31nlhYa
iHhXArr2aKpaHo0sQsq7O0Ez981ODK4yYLDnhN7QI/z8zgrZ5fGdHe3tDv/+wP+W
Xld06fuCok1eZMzRx0yku60+wsbWDUc6qbJ/jDBWDYqBxT1O+aQDuI3WDKBpC+eH
qPRllqJIGB++VlcX9xcgQErE/EWsOI+AMpl/en9qzjuXY+wHf0t5pERhOiRoHkfc
lW07D+A/vup3c08F8pKxGzX5CORN8Oz5mRgi5vXQ7fuE3tQ8ihmaCoktif30yjCs
XnDWY6/OgKVPWRZx3N1qlbqZhuQ6bZr/TUW9qopZ6R9Dp5fWLktsVQe5bEdTK/7r
bD4V1vPWW7ZLiAqbWuE2xV+nvOnP4FMvFN1NxMDZsvCcqioeECrwpiq2rhO16YGk
JxdV17JAGQxCOJ764qWkNQ3Sn6stImc93RUxxsh+or6YgYM9Kn+mAa/JyOg4K97u
LnF5AccTBtKU7X0NTjjWH8OezgYL/CiWj6POehapA6rT03bciMTa4weE4bKTyJKd
rDeKTabao4y6Csy5YsbgLJIXCrV/PaYnRwpGlWmH+2Sz81eLYJds58l3lRTZV7tf
5tcpQ7DXTvIZMpotNWniMY4grBKVF8d2TChRFNen/d1ut2NSyIgM76lzJS0T2oSL
AY6KU7/O1MQCiQaxoX0+6aqY2EeXyrTPVf8iIBpsmgogldjC2uMpoolhOND+NF58
/TQkF5gSxQwh8VQg23irDcAJL5JkKbtDacdIbBSstKNN8xnVnqUBEnETuITliM5M
LMSv38hEkPlfzm8usT0h5/HYYzJwW/o6JsXRRHx+tdqWjdoYgaz1RPVATqgiCHGq
1x9LfBjdJe7vA8lpaPcmHbsPY8vTl/Sc2rwNuCkZyvk5mVWpeqvBoBElnHwC/r/g
OF6F0Tg69AHvnOqkwe9qm2H+D2RslMZnHFpewx/0Kxi/QE3wL7R8Du+klKkJlJsM
nwpSFnRVnrlu4rh3hRbPN97bSEWkKTgmOxFvTYdk5VBWuk/FjKFCDndUm3mGL9xF
KhNYCMnkwF2A65GYafbFUSFP1MQMXlMWAxycYjPWYECf7pFbu0xO9AxQpt0txDeb
V4iIPMtz9i74UE7KO8w51IoZ7Jj+igNNqua5+gvdP90FCDxXiv76EFtViMj8O0TI
w9nDxIVDQr2SFntmg9bsEhFJb6I0HSF4eXdK2PvLKvQsBFZmqkt7eMj4JepWMOh+
oLAP+WW6vgLYn9lHVfD7KHE3AqMPqU3P/zlHNETuNb2wFtUbfPe0QFJeoMTgPA4E
lRu8yj/cFSYf3Bfe43NumP+g6go16A6nEQfClMXy9OnzMYMp6vlsYbMexBVeAGf1
O9cm3Y5MwTG0jcyiIf2vBzwzreM8+8zY/6sPRiqKNFYBm3kKMIg4pAbFeMYA96Cx
z6s09tA2BkAqbO7eirtbS8bkM15fIlLZ8ypkfu54Pf2agklRvtRgYdbYiB5dNow1
3nvYfiARz+hXLL3EiCSnlxZfusvW6WNQvayaAtRSOeHUzJH6PyPFDvHymGqE3TtX
A0yU3Hzwvch7MCFuxCHvfFNDh6mqUP4Lfc1lcTjJcgQSLMeOSrqzAH7FR/d4RAir
MxhKoMDuGfVV+8nA5Zc2dTCi1qKRCes0OKqSYO+sath87dYb3dwMktTVAFce2CkN
qaTiM+yhc0vny0PnwtRXuuD/QhXrV7MzlxSnsGFYkLJcVpLQhU9+hwZxMVNiA2zE
dtlRjyaXFYv4da0bvbqVpokRH5A4wshkyq2Jsw07aXwRylTLZZRSaSfyWNikvPbR
7y6DerfuMlp617nvjkXiW+Dak/b/JO7FSe1c7zlc9kfmjVBgACgIeBOW4HVo03jI
8sfvAOwUsvluSAvOQ5XClmxbk8VSz1qbl/+p8soomPPV1dWZrfc19SIj2TlpEZXq
`protect END_PROTECTED
