`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G+5oMIgQJangs78Q41FvNHT3nZ/+vMfLiGQXSF7ZB3A7ObeAz+1tmCaHmTfMhtqR
baQT+348H0qXSImV8E78vnfO/9Y/4qEtnRW7uO1cTIl4Z5dI9BDTjrsh9yFld9dB
dc3fdwwxdKWXtZPFqNCvYcblR3hZK7psQW5jUogGRTou13Bwl2pvarZbX5TrMNZ8
K9kKXsIsuhrrfxgM/oa2J9Dar+qK71ezCtU3kbFXcxn7aGyLzIqliuNOPqi+EQ33
aSV25YxFLdZDgscBl120/gx9mN5VYAafmJLNTgYpdx4dUglctJz0mbbI9JXqQ+Na
nJb+Q1z3iZV/HCe3rmbMA19T8vsqFZPr56n3aGRrdj3uQXEQm32a0Eo2gSK6e3HT
Js4iCvb4Q7FOIQhnXxYqL5T7gddoHqO1beRBJ7L/Mr8L51mn3T7HelttUTeCGLf4
TodAj21zs9ejqZNu3c50WfJHO3nzeZrWrklwiu/wi/PRBmNtHr0dqWBHYw9W7JSi
W0g+dflwQUi4uVwclkGg5+lgm4ru+3iwj2881CZp3vsxw0V1eW4LySV+dDgS8McG
g6hWbsKYCsNHDvrBECuJgwQKoXzTQkd9S+xgm77RPOPs6ma6t5F8wXy2VLCCKkG/
cS71kSP9K+h80rslqJedckTFhRjXmkz59JACs83Csxs=
`protect END_PROTECTED
