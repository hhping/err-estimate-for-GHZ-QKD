`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZAgGj4wCDZAbzrvD7Lyz/kxL+uXTCkv01c6/TzN9yQIvE5wLY/fTSo48SZxgBS/n
t+WFIPda0/zb8mYVvSNp9rWs/F3erxRz97WBBdtHGhft5VuS+Io8Acq5reySTzvp
36SDxbNxZ9fCYf0fUgQozL1mgOE9ioPdhWXf9g9o8JW/7caEopCXuffs932JioVP
6VYBmUga2XxaQRJ/il5/eS/RpyrIZEQyOMexHO0NanFw6hk2HDwNx3/t5BNVT3ht
hLuY6vbxbwZ8oafH/JpTjMi3PZ17JFkOuI21dh+OlhRMjpglOF0NWAeYcjIvdShc
TpewxiMFPSTjQV0Cd26URQGBbF3qYYyw+DSnK3TPkalHeEfYO7rP3/0aSqdUsh40
d6BycnkkHL4T9uh2aFJX/7fcwPz6i2eMz+cTQjmXxMEbS2Z2c0gT2OwtHdzxfW3q
F/tAfCTNWGQkn09MaCqg3Q/o9zBbNDUdPkUlbaOISv5v+mljinZX3S+kiisyGIpX
Zg/fRX5uxY1ZQXQ6Q0ylAgeNREgZZRS1W59bNg4IAA0HE5NsFDuyflb4C47O9vGO
vZ1zz82qGegcTCuWul+vKJbG5vM3smHs6CoaFkFpW2qjitLNnDTg3WCHqoMUoAle
F+UAJPz+08vbriCgbwYD7jf4IWXbv6NRvJoAatsg6G0aJzBGAtNCrOwCEJfLRiIq
MktaIUoBjXMHCsKg85vuUHTvRlX2/borVHBVeg33SPKi9TerL6r9fZn0I2Gfa5jN
vJd09SyeOvyuHSP3grQNePDpzuXu3VhY9E0uL8oeTC6ZS3YwIm3lilKTqwKyGW92
aqkzsyLBvj6WefTM90DCHBSvYOeoLnOSq625nzaEGnJM/tqL/TwJ2s1jVahVaGuv
Me6vgePsSGVat5dqdA4h1Yt6zBhtlYiJ5SO+cH41DmB48i6lHtzc51CSNfidVJLl
axA72k0n6VQpq5O9GYNWGAGXvK2oiT/z1jPBuOExGMsOA4ypMk1bwUzKl1uUDtzh
q288FiKX7KyDzlgcplBEfrDV0n1RNpqxpMX+HJolChxhyd0Q6a39nbSGdxc6oI4L
2n39P0DLBxy60V3xYR+TxGL+1HXTkXqE4hGzwEuo8rymgmUW5ThKKBpefHhJChVI
8DaSGnZlD/NpJFNYWSLS5Dd+vsWvvMqVC3INvJL/MH4=
`protect END_PROTECTED
