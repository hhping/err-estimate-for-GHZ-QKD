`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UQ5k+S8R0520Fyk8oPEqM3kOqPgcXGFkiicQh0j/URtNSKWY+jwovfL3Jfwi6X4Z
P2lcjVCjXi4ktqKA/z/NqOmXGovcDeGkudIIpdY46A7LbTvE4rDNG8wiVfndF4CK
XN06yE3ys3N36yFkPacSDbAnL7H74AfcRxowcBzLH75N9gmW9eV6B4CfZrYQ3/tr
hXpbL8J/beaKEOjpBLAGaOh+i4OqYIjZwcZgwryC8HNuVPkzbNYZcGMeL+CClW0I
4CPnSNwEK+mo/r9AIm6OZ4g3KyZI9GUz0dP1Qti1yQ1sbtMrXgOI4dBNKv5mdDqm
LHUuHDcC3koflKyfJNDMS3+n6PMdhaVUoyJ8FS23/wF5HJqxn3bTzuDB7G/thYRP
U3vx4jgLiYwtZMT4vzi4O3bXKoBIBd6Chwb6SGR5rzJPE9UKZa9szBiyqakbbILg
b0ZN6Urp+UjxQmyt6zo25bjBnD7Jag8YaItKkGUhF0HMFBdIuFNFg+aRwxXQOBYW
FYQpJw91LZ/8kLW43dWqKyAiT3tExBavpBkqjjr8m+cvkM1AtiACZevlmyTk5NMp
R1FB9BEx7np8FnAacnKjjD7Y1RWLxm5bKcArf2DQOCxJfFQqTLuFMuECVAIwiGfR
ITvqwSCrLl8ghb6vzYgUe8+KHVcaQC5Vk4Z5KAfovdWXIgthS3GOK3/4EbExlCtA
1xmBKa6g/KGNGd4KYEjO1iXwSLclUzKqLRrmkvvCN7+yru5EhlS6dDb125En7eOx
ZyiRigG72bSp9LgJraY8YmxrWV4Djd7RdgOf20k5ngWe7K+2NromUUEvw19KcKwD
W7Bs1e5fbIzewjoqI4mVepT6vOSqNShfGMiaVRa4rDWupNandj53oGlIuENXG24r
VTX+M0IGB2JcY2hsL4WVmAIXId0kMztpx8JcZIOwDhVM7TC7Z3gSC7aSaknDLk7c
zI+gra4rhuIQ2VcneIzT2MOhKYJc21CHHw+1gaj/LESfHk1Qgq/RLPApLcz03tqa
yerCPDkB0vk6+vfzPzs/jfeiwFKi7jb900Osd2nuX25iTxrmL1yic3BqB6EpHpKH
AtPZtJiG/j/y2ZTqi36nvMj5vR5ReoijtAbb5jhQlWzZYZat9HPwdV4tEXM47flD
xUty+gmi7OtuZW1xMD63QFuTz0/IXuC1fikJOuKemiYq6AwUAEfi1M2hRF3+kSHE
ZJZvPzC5U4n3whiSA7Zum0bWsj25UTgCdvL1qlK+HASjV1PROSOUf1dgDKlAjDad
JcBzolgUGlqFg8dgnvXkyUg/C1/68SZLmQm8JH6CYZIlODvsHKA6IBhOLco3xbFh
lhqJjhM+7T5LPx3lRP+cfCBNSMeb4+FRdYA0P2hy9m3kPdmkNHbW3f2oeUffaYGU
2/GfsuntAe3/SD5ixGlh71ibk902yDysgZon9VJ+4/CeWRB0S1YLg5c4wAPwxQ+E
mT5HQBlYTrYNnZ672K4Vf1YLuoxibJKOFuwJlWOgVDhjDG7IppacEwmPAXANtmtR
YsB1g6LtvPV2Yp02nirqcA5Rghx+T9VAMRk4ZzEN2V/9JClHz4mVgk8qSG+wxrJM
alxgOzqj+rVpXXhumN8J0s1tUwJxlpJZTp/v3Nu4pTeUGOjjuDc7f2dnbO28jpeO
lpE1FchRoBZ8wcfEGXsXhyqlC4gx5oWtIH7CwNpwRRlu06k6Ex9aP3mDNx87G6Sd
G4MxIkmFvyDzsczU8+ivtVUSXV2dolfc+Mu4+gGfapZqTj9p2K8iV1OSnKkz0ER+
A9rOupwG20BakwOqr+na637BnM9CcLUxgeVPvlCrRBzcXh4OVNqJnhoDUKgmaVka
+2gvxF2AvQ5ajZNHsq61zFmebIt6eDzR7KPMoRH3iwiBP5UtZM3N/WtyYVwKZJ6l
Ekkdm2e9YJnn6tgXNutuXVtKP5jCNWZC1c84Ro1sWnrONtU+GP9k5bzp3hRQXUla
v0DDK8BxbdTbvoWmPAXdLRKcHvuIJ00b7O2uPFlRdy3VdCZIP9CjW9N7m5WJr0Xs
x/UyIPwFTY+hXK5Idsl6tG3oL0NQHhiIRUY2W1gEj/g=
`protect END_PROTECTED
