`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M+eGgsHArRnpkmxjgHOVywLJsWuVuAQVQcomkUJqolP6SheLduqLn5U2h8oo0Sr4
V61TuhgxhDUANu85lOAXymuvzdvHcLqLbWnQ8+dKNn3LvxKafnXXXXkyNeSlQOQ4
BGYVt4kA7Dq8Li9pc5Hrz31HsONwISdvUO/JXHeaKw8bsMsxc0f3DlMkYFdvr8Vi
c3bPAXdruRkD90cXympvd781Eo89G2iDyNFyrKN7wZLt+rIF/QPZJsJFAJTQ8wEB
fJPdXaIkypV8s0Buup71inTd0He/UH0vdaIz76D74uWGUstQqRxpdOM+6krAKR66
tPlspDu1DX96/FhAY69ep7Vr0QTKE5BubnYnHPBpf0ciUg3OCa8oNYmwB6OHhrmh
pq6PVXF77WzG8Mf8ftjhEC4rxV4G+Qga3xv1i5QBrnAm34tmqb+Yat6byHm+huve
MKmoQk87OqjfVrlnoRRMFURjQIxI1+AyLiRE7GghbOnOkFnV6+OK2UU9ozgONy2m
QHbGMGWPaiFgn4d+CRPC20sBsFzPbP1Xsg41EEt8piEOJlw2mtMiWbRNwJPR0lXE
NBnbUb/EzUwAj1XRpoM5sr5sDcEWqe8+pf7rZuLM8IdzMqgRrp/9sy9MfSZGAZKW
pbYx/zzWYPTHf3JCQ/G6IQ==
`protect END_PROTECTED
