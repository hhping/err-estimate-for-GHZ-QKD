`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SXBWOH8jCiGwA69zj5cxbFLF64PuA0B9Fms960Ko+5jLNi+pnQyii5ORvjR49dlN
K/7aGZTDKmUKwDXPNenkDD78pdwxelIXpYqswsHTr7ZN3qBo/XJLx2VBz0PKfOnZ
uGHATyox/uBndN/TAIC3/6ZH8QtaYtoEWQ/l2u4i67n5PS0iO6i9M6ZLGT39wPlq
E8RCBAt61ot5r+rJjQsgucPM58fzQmacYrgQYXpmg0hSt6rqd3TErZTenIU/ImBm
UBBbMIBHkEZWJhyf0y8NxhXN/3RBA3yEZkfKHeAM14IPfjXCQ5Mf+ycP1enEku9W
ijeqCEAL9nDTx/mx8C/2LwsAh/uAEPZ57LmGaj5SRTcTjJ+060Wgcsl82Z96EAyI
QWcbanbr2laEJbxec8sNmiPb4yF2vRb5bspZ9ar+eUjHIzda4bUaIyxanB2sPA/E
Txz+RF912lBIewsQql64r+Vom77OAP9O7LKZR2b2gFBmFSbVb+qmM4ptnh6lUHVP
9SqKVGw0gbNGR/AkzsK2LcfFBSlc6t472NXzSZZSevOBOLyk0m96TRfZFX3QwmNB
pOd2YrUkm/DEzzxv4yRSGmau5RsKfDynO2BMr1QDIt2NnVQB9BREVqUFaTHZfnsy
/1Dc8/clw9LW/fKs2nAXKHrvHn/qMqGNnfnX+NylSRD18H07zCjU73nHL5b+EaYQ
WZ/6kUNmpqYBuVolrx4byUupu7xHSQbZ/Yij5NOHZE5gblFNLndd4TVSLCRt4ioY
A6w1g38H1xjv/kOEojDNt9xzRm9YOZmz9wSeHoq59hD99Zy1IDrTjAuBEnwVRPnS
c5qMiDTgmd+7MWbFoLBqQItG3HFJz5jYVIdYwvDWjj2dgl3hY1gYB5LwfdQnGfBr
TyzXYh0AOXMSMDVY8+NHb9stYicMjfVdAMw7YiEpvKq94A7/6aHDUG4qkUZuzevp
WTJEGgKpSneqFxCIZ+rwLnfm+WkF4putY7Z4irj+WagdoKurPJTu/9nTEOxGiImG
wRzsvb7BMvemF0BshKocAMBjxs+6ei3mmKqv9cOLGOfLs9Z6/SbgE99U1O09PQ/D
EKmnypEbNPerMY6VUVj04g6xOU6nqlEGNno4YD82QufsulbAPSQX4swvpgcmXQJj
1KDVmisED4LhfLanMgvWSoZMfgCjyNux2gMyZB5U3cQoeXys3BRAzSNOuAbZ2h/r
jWlDBCTi6GVFhTf6HToS5dd/Gwn7typw8p/yANOscr7fOMasz7Y6BO/9d+aO4rDW
IT6UjeELYpMRtiZqOupp5jsfNy0CkggLQ/7nurne96FftpQvRjmYdc0R+PouTrxp
t/gobOB/g8LIPybcJScVsde7gNqN79s77ZXmgZG/61l0w6lsC+FqKENjIsmMpYG2
Fg/jDRt8XmMbaN1RxB/xAHKcSo4b42bdo/B7K0RZzCncqVjUywkf0e2pZ5d5LFOR
0LvuPPK/bOgaiQ4nA6pDimOcTzt9IgWL9Cfct46IrFs=
`protect END_PROTECTED
