`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UuN1IhtdbPdLFPCGgIMEThOeoGUrFJdK9H2W8MJ2eBx3w5oaJ2h01p4fO1savrkE
tD6SuGsEKOhaBqvM+maHKkEyO4Xq5ArpoO8E63AG2GVAxQZ0Ah/VWVtjrv/hAqD8
Cwu+TwPQ2SWrZCnXcRWTOTFMOPsXnW0fPkfPzU4RW0jhrcG8CsFDaJ0TVY94/bsx
jsKfxPau4i7Dfi+H1xG3EVwflSrL/muulJwfZOlf9M2fJi6r1ctY/fqd5uVtxdKz
sdRG9t8NeEmVS54WnjUuk7goPSPXXyVB9h0GZU4i7Hbcco5kvZOWhsD7NH0oh0l9
iF3GB2zRAkcUpS7JFd7ZD7Hy/w08HB+iekefNnRPnri+4fHsUXq5LZ2ebc07ZKyS
mYEYIL+aYEog7M4IBbuL2ho1jXrMEgBJPrgCfvG6MM8wTyJcq8xxCyl9vWjLWu0U
YOEvF8+LQrFeD0Z661OIshNia6Xt0CApMhBcrXPSjAze6Ipdgkllbb3ELPc/LNd7
FL7viWN9d8LDW7e6EVbVfB8hNakLKUMAcgEt0c4ZTRc3wo6UA6hmwfi6BIzKGsJA
7z0mILzbMZZz4Z1bFlRxEUgyS+nPTKppe1MPceSMIUX8UwrOzd8DavTb7U/JHqD+
gm5RKtG6JZ8TSbdT4SwZxezTtsjXHiYVt5ml26GLxymDcBSVCbXUaDCD87YPl/YC
Lbbc65KOyHjIaimdrF7mYl1adUljPvQ00HYjutb6TeCqYcL5sDxDNZvcyJrmvNi/
k3IVv0GEHZVUcOZyZLgSBHe85UePQ2O8pVLeCVTXdB6vhrOisToLOAC64ik6bheo
kHbAmqUT48KP8vrtdo7VypvB/ZJc8/Xr/MeMtIeZf/5Kop7pRJmLarZa5TKdR8Qv
GucWuHOwNEVh9i+zQjN3DHKse1N91B/wv41yji1x/tjkKcwHhJFHV0C8ZB8HPtE9
bOgjelCayb7m65nKG1dMODT5uQyW8QbjRDim1GYC6TzyQrDKzJPaju8h/k/jR5XJ
+uVMrdN/NnDTFyCOJjS7yH0rVuF3Ut9y2AizaonGlngGCMIBjUQV5BizoL1Nm8rO
EKSf34M9rBjF9mdRkXwTd49LcoJKlP/b/2LPSbfPKICem62JSzHdbSiOXNW663Ja
gy9G5O7nsiBsHWL77GCnI4zZSKQ+78YFG4Chb/aaWy+jOlP3dOV+J8EvFKWrz5ok
hHvu5lse4zlrtdrpYwVfZTsnlPg4WCsyzttYzzLXHzXbs05S4QGo4iM1nBtTwY1q
vkfADNzNYeDOidFMDUREgLlVAwpl9VpxDMIEzWS5SC+c6vG7Hp1goa6IySABdpBW
b5TIEgb4P8swXIoUgsfinMrmxM6ILSzcImo0X1TJKKdQb15c010faOqoM1pkcH1S
jU9/EPbqGlBKbaWQk1mvcAjQ7yfDHcO/dWmFD6rf/cOMNWZhFJS+/cY/Qos/MeUi
cLEKByVr6yKr5bwTbmD2bn1kB0Vr91++E8IEAzyyCOekXbiLvy8XqhmN2A6OzedA
7FI9bX8MyKNdZaqB6eombexLTJquI/FdFPiEahgUbOR5bLDwZMZKHhCosgif9DG8
lGCjXt0oVkhohq6/ZPz3IIwBEAJKfnYRGOsrdOEaB99N6LCDx3HatZQPhSfzQY3D
1wNTFpcKRyzJSlSC/EEcUeq68UNo0JGGdzBmW2YrRIJxYQB8rWJRtyXs7nUrUFVn
AuB/qLSsTv9mr0bg8413T8isSdEEG6X68M6hIGXSjRJ+To9bPUb2guc/OnrafSaG
DwGS4pa/G0/JkmtRGxl1mwo9mJFoZppgAeW6cHNXcAb4fO4Lo3UQnE9ohE6/4WEz
hmRpXBTABzDvKqyiEXb1zj1VeTcehjmVe7TZI32QANGbPyZEAHypVKkVgP+K9fGA
DkfyDZkmVdpjU9i66uuA6JOm6tHtIeMxxiuobV0v8okNpzRN3pa+J2CMSwgEuzlQ
Hqa5JGEDKvfxkrtvyG0IRysp5rqE0aqhW/enbGgdFUHgmF2l5Tc3O3xjnjwtY7IM
Se4HtK/+wyjmFV8yIkMFbVw0gkAN9cREgxh3f2qPdfrizsMMkSWxTrxt+BGWp9a/
3EZ73wSBeE4+lPSdPTrCVHgL4XJOBTSuhpSHsOtOANGjlaCNEVPW9DDf92MzxN6O
WWccFsLhjEEnTxG9WLXKlrvlLMFJx44lrfqWq+JgCemJkDN2mNIjZYXq8Qcd5BKp
cmY7NzfujFIiXbyE5isVwH7ReRxJBsRmvGT6dc93pr9iGSZwvupWZk66WPg/2dDz
k1g2V1+qeafVAKfE9z3g+nslrh8+zKnYz8NR2lEp/b+qlou+pwBH7oPBY9Iba9vh
NWcnW5LJWkWfbMU4/4ig0+URMMweIeF8UPPl0c/glunNTNkqWQgP/ib5Qfb/Mchi
CRKlYMNQuamXrlLEPfvHzSLToY2VaKs5hQC1Smi32B//dA9lNyEDoYrJey6Nvo8d
X1fBaSgOV2rmgR8iups1LQqA3Il3AN2H5lhltUcV5uwRDuCIAb5W/Z7vXX88GKOt
H8uzjCyIWmmrHJ1SYkMv1AY2844QzTxpnEGe8mCaYjfiftv4XwZfyig7Rv7bn2Ud
UShU6ro/Jez/Gf/HwFUEmlXhXUVMFynG/xdfFmL+yknTkmFuUhdOQR1y44VCrZs3
Jp8U1/BHcvKesPRb6G78qpYMIauHU+UxRHAEOrGwzBLgRQ7XDDiTVqqyO9jTvsZF
qcCyBcWCeqSGOdamFZcO+Dlj4fhtFQKibLeFj7fjp9gV/pxJ+VBszJrtuFmEkTkM
M+8O7p5OuDDWeG6uwtZ+4aa1t/9tbOZ5t0eRADE0Roxi0wrvgJdah1uVKtYE+y2I
ap23vvgQrcJaXG9uMOpeCgP1ZstBPTUvrJ5WqudPR+fHsk1fZD0u0FIYEyLU41IO
jWmiYdBb1m1TMw9Kv081BSLkonTY0CXI966P4OGPE3uUBpirfDftqgKz9jgRwFrp
xUkVMeWcPrWoyqtJ0JW+IqXITkhVu3vzl79psDCGgPYRNfj8KPI6/p5MqyBfBKgv
S4qARnPFlAYGS6/uFWYBpARNTcmzjhJPOILzLfRVOmvDwBaTuTIROZHjsy3fAfWe
irN570/EXJEkU5QVgWX+Efl7iT/Nnu1Z3g7ibBvu/oo8NWcvNsh2nBj71VdvAn2i
L8KgJm30kBFOsi0AnPUktTGqpA14+J3a/qXvhRc8rqFxGUW7qeB0Nx+f5yGbfiZa
uOHKjRqZe7BU+6KmYAK1FA/Tt6P5E2upV5QMfmIG2Nv5A/2ZmxnQckQGp632OXA8
mRxmJUIzdAjCkd4pToKxChdTcpQYamKLumY4P2IVKN+bTrO95TehflsRnl7N173H
2NSfkY8cNdPNJUvjUVGSrHuHoqjbuNZ3ZFjLYPLQbpEAtTtNAoDNg/1hiFJRGJLQ
Vf7fvyMt4Qss9dpQKKddF4sZy/ck/i4mMPmRGSq3zbHJSVIuFbTkgoSkRbHXDrF0
wqWQls87d/HGAe4+9/u5QSMnRy/N5j6pEdjzF0phOUseBH0HwfDl8bDOqz+a5S+d
uA6///l7Kii040Xp5JVCgFBuYq4nVt58CRvY9bwxUlFVn8PcDsDwqv7cWzXxra5V
NV7c3CK5DczSleB1rO31tTmdZeN9xdaI+JRDt2Bu9pX1rHlSleo38Rj2DRhG40OB
uhp1Xd7fl0s13pA1RQgwB9ogjI3Bsgngpfm5MMgQ9wQDihwWtJ9osS12Q926VQx9
T9PiLWoQ1VnS25rDR0oKX9Si86IJGE6PRJYGAgrOWoGxLLyl1C5yAJEpKu+tZwjc
QsPqWVyiUY2BNAjEoYpc3FIOdF+pSmrEVaQqWuJhG79KUVf+2Us6dtzcAuCxBhjC
fz9cMZ81EMoV+cYVRxvV6UyeQcChO2A9u9X6077AdK2gYhVxjeh8YwE8wC/NghQO
x29c7X62Rpl6XVW39K+hS5JLb6awW2BzqjKig3R3T7ttVAHX9lGWqrL3xBKZ3jzj
CXxbPWNzLkcpRyyoLyKV+b0IDKge1r4tSiPn72DyIz9gLxkUk1+p5GBZUMhRHiy2
fvjtIj3VuigzMvSE8MD44LT9k4PlfnI+ZYB/nFr87tXzgJtF0xIgZvgWW0583mhi
DjKMmG8lESDQR5FrxvcU+n7UhDEhoSNEuPURkEm2+F0cWqIF6boWHLSDqNvcTMBl
whV96gSnmpoL03ZP1g4j+JmZe25cLQXygvDWWoUe7BCd4g4mMTYobIClytR4Iaol
JlBoxw2xn4HjLgtQxhdfuM9LKg72mEefGcDZKXWYjDsScoc/eApCv2Fgo7/SlUuj
IKS85W+coQNHJ8mBa2r3YjHoF4hmuR9R1FtB6aeQxFPMU+FIpEXAMSlQ3h/ZSdUE
yf7FdckKgyU4K+zCeJJXyRiQ//5d0YM4nfB8PhEoLoSWU77o2UmK9OvwcT4iusE6
ZH88BKaeMc+JVay/NwPovW/sQqwWXumMFvHD5vf+GJ0HbAb29/0AWrNc/bTNDfhU
ziD11eFkg1eagif9ayF1ONSf19QfmsOerH3gm0GvA5FhX8xuiTDUT0BSw2NCDah3
DBDBpcWuKe2ZYNhbBQMLyvf9c/t6gF7UzwFEDjU+cxEdOoL/2OcNrySs2Gv2Ov3M
b8Su5m2qTM2sCCf5Krgk0pakAC226DWkLvjKTyARocDO9N4hxiszWyNPifrbaZ5y
G/bra3BP1CtdyiafbdKhhVlvgRimeth3nPvt5c2h3yn7EZaXJ8/EfQsARFqNz9Mr
g2z8w+TLOLzSI1GC37ZWatkSnXkBLWhq73iPTkL7z4Y/++W0nQkNjVEPe43wN5Eh
3XeVj7OFgHIsDuEnECVikj+88ma6d5SUt9lssWByoSUiH2Xz+6xSyeUKiHaiZcDg
njB2F0lIgrS7lJGSfPTYamcIO3UswpDg08Cb0RFiyjqVWH5AYpHP1kw9R4pwvCXv
a3F5KPmHJGZ7iS3IdyT9HcGkiBxKRpW7rt2fjvbmolEY54zF9B8Jphlo2G46aAHB
EEfefjXTtsJk/U84jWybHnvVt+XAyfMHpP9XGS9OEe8tZt22y4exKnfeaxetFr6/
WMkEagZI+/T6Ta5Af6UmQTTzBqV5wGAQYIcJbXQtDGkmVUCW1rYBSn96iGRiQkjc
8kg3nHv9wO7crSIgSBH7CrKd6PV6iNCgLPxkHx+zCpr/7BsRzblkuYhSqMOGN5WL
aoAvEijqrqrenpKbQhylyjv9Mh7p3t8/myGxyb/r/9RMADiWcyfcZlugKNYza3CC
Zx+GKVZ0swH4t9WLJmjpcFA35jI5utqbE3+uDYoSf4FQ0zyCdn8rK8d/gmCqnYNj
S5wpoK1orzBCHp7kUCrJ9ik8B/oh0SOaP78LnYIO98rrKCfFLhf1jh7tWjemTwI2
PtsFM6yoz6rr6k/T0SV0Z6ltSlW3lGBFAdQPXmeItnqlASzKfeHYUOuwVJqjSvt3
Upe3i2YvcpQbuC05FgsOgKJ9SQnx+ghzJ22rwTK/keHYqq0j68ZS4MFuhKSAd6Vi
clT6QAvwRATTMyTRgP3gDdSwinNRI6UiZ2jCz24Bh7jKrJ8pG0R/+CTLIi8H31Mt
AOI5Kci9bXZFOWsPy2gSZ+oJ4EHUNijM+pFJZhVb4AJ4yAB9cmZ/AG0mIr6Z5WLj
b5qzjCeyZ6DIkTofTQ4FkV6YFSM/tKIKYOBep0O3SkMEjumXV7d3udRN+F7I5F1N
psnfh84pUITl4XUu+EB14H5F9r5G5et3BQ32oNbRS0QnjOm/cX4zKxB79kvrAuJz
YvmkxMWoom7pyCntIejAzGS6eAbxns8QrDwWfJEezylmoKHRcIUhwVG8+1iLmdYG
v6yx/zMIjZLdlZQCe3GPQHsiSyE1cy/P4u/GtVqD8jpaRoJ1AevamCftgB+W5kmF
82/9mmKY7ttFPR2aQpsR5Gwp42yd2ZZbBgWoHuTad5WJr+RSE61fdeCOV2rq5NpU
hGSEFkhiUBc7ivC3mE3fqua/gDmZt+5x3y1UjG8aaj6hrz2eGHI/y+dJkPFZOb3Q
EaPhNa7E3E+XO6bFhVLPQkgjwoAWvDxQBvCrL+GonISo3lcFU0nvFRcxvbFNCcyz
Wk9YDsIMEqru3Qz9CWlGkctQTIhzA0JWZ6eyq9JPOSenybsQcCbxlH+MRFo2b+mB
TnVDf0sDTdrwOeL/K3EGpCSdMOT3dkafDvJduXNJR0GON3JP4F7ghH89wkSaozDn
hdR4VpFkJ4JXB+RjeBHOTiRMfwMeSf7fdNwUqqnFG/eq4XpY6lfXqZtwOjL+q7XK
tncAVmbHFHDF1q0AeiPEcv8YLhWdvZj40VaaR50INMgwdlV0xeH1+SOMQbppqa+7
STImlvexQoQn5x5bTqwULU3S6Eh5Cr1CTN0J0NyM9NPrY+yDvJ72q/9KkTZQlR36
GRhZ2C/AXbFrUgJOcget/pPdVJ28Hu6Ff2jsz3MM+cd3ESYp5e1SVCWBmWf3nkQD
gmBL3PqbPuZbUcueIYE4voAvZAklAaFnbg9P8+AsH1tqa8B8xiADq1lfKvvivp8J
aPO/M9Hvc9aPlGFPKHj3mYYXfasp5kiGR47CoF4nznML2zjcrl6J3ldAJ2DyLHno
55gvn2e599cs2V0iL6MZ6FWQRsskhE6xBt6HZWqIgZJFaiII+61dX+0ifWrM5F7K
Suw/GQnJx/Ppr293JOqipbJxbu2KTljR3cjV3bFgWkIaYfAwW9hw4TlUFHGRoeMI
7bmEVTd8S6xAPEVblv1iHuFJjc2mfsxVmzMtxQXqzKSYJNhPjSi3xBnHn8icx/cY
B9LMbG4Koczf9aATmD2Tu5kOWkAPGCe9CV6hJ1AkRw4PaznLWT/+K449m97zbhf6
SSU31RBI3IChXGPDPYNocoYjQmqGKgHXCD9Fy2U8JValJUhD3TnBHOhUZT2kUEpy
V1lErkj34nLiqLhkLYLbYYubs5V7vEKjaChM66hDevxytEOP2XfuN2gTtLdBx3Iq
vERKJUq7r+4ed76FN8xm2w9cmhE9CFWMp0HWvz3lbF26/CCNrC+/+wSCvS2tpwqe
pKcZs5v9ZLN+QE4yMCs3Y1XMAFVsmu6BGFmie3Sycv2KHNp1m2xOm90jbNjziECz
R2qu0k0uOQAmx6mMVVKj+eeD6b1k30r++Epa6rEQaXr5GaLlYztQMiITNrPZIRrs
nziPYUEoIwEMhvizFk00gEAcZUNisM29ZPpzKCeJLAwOy/QP5QgftsGxyFPW8SgX
NQrIWcqijZB28cRZoFaqSf03dhiLohIw54hlAziWnG7VVOPzildvtgz6Mw317GfJ
7+18AiQTjxWaWfh8hpWbjlFLPXrpVeefMUIoV6dJjkMEuQOEEdjoeU41tAKzEFUJ
Q0r0hbWeBYlnAEcF/lu9HsvGMH3Hkoj+HpAF3B//cEPMKNIlJFxA50+dak7OzVxY
N6g2udw7LN8epPINzJS2DeHUxPtfqyugMIS2DXYUQEeiMDDuj5SrwmjgNMk8OcOq
b8P8PNo7RtDtNzLZaAqPhiV7duhqeOpkzapD2Unr6qlSmbeEmQX6P2ooo9fIEB8G
Zg7GQSTEZNYawntUaPiCMXHMZeO2oAypoilOtRNkjQYZ7gNc6Sb/gwja3zrrTsG7
1w8XeImn3l2HYMkAiA4b4hfBSmXgaornOx30+LU0hOv937xEWlKc9ZqgPRqI+s5L
djt3ubbmdVrA4tKAc3ntzBCTJQHBYPKsYRuWRZe5TbdI7h9Nh+gp0HhzbW+kugpa
dXEecaGcdXk0xyxwYzIziLZsdPKb3yols3QDhC2ZCMs7brgQc1X8ZqNNgFMyA+dZ
bhGVUq1lsKDIaFJCC8Vp44rKHsaG7bibQeG0pfM/GsXL4eGwwTh/RyoC22Ytgg5o
oZWaY8eXpkbhMr3iiOJuW0WJDFoMhFtu/Gu9CS/2i7Bn5urKb0ARSM7xK5W0nKYM
a43drq5EgnCkTdNL+hvpYLvX3Agdi9C2fKkDkqRvFia8v46as8iw1v/oyYTHlCcr
hotKzKMBvm0YnjoTGy8dxPfAJ7g4TZmKVO/tF58t8kBfnUmK0auIHTR+noOziaCk
O0eUcIID9qg/Ed7B1JyzLcFLGj/QV+8FA0lybps6u0+NhAu6qjHC/34HitfcAZtb
whU/oSjjUW4QPEQ95OhgEV/yq+2Po0iONSO9zQt3fmZF8Saa9fknKBzEO4UaM9KA
WmN+6MaKWKWzuTHb1qWHGycmwF+nm+gMmuJ0r/FMRJcVZ6aOUsggMX4xlYe34R6w
VwcPwJS3Gjdw+PHmOwSYV0lvuSCv33/sWnmS83feL9NLVD/1yB2pEYfzjce4kbez
ZW5SKDys0swDbwM26rPnc8DjB8cloDBdxLFq83riIqzNkVrNDJbxuAz/8fURqmzh
Zrt0DzJQM3VufAUrbsBEoZyPU08yQ9vW1YhODrr9IoUQJsQ4Wd8TkF9X+7AH/5lr
U+TsPVJvYWAmMrfzSGkaLhoKlrwcLL07aaFNe0q6LzrIIHF9QgHQhxOp1TdBovw7
TTeuF3HJLlXiFolhTeBM/nbiwXSijF3zHGsSrxWkHf6hL1xoZouYTAu+JNMMWu8J
BNDBFJh0a9xE2cTaYpCqkPYG5oBJLtAFfz0q+QGNMX9tYGBC6MlCSjk1fjzKmScc
iIB0hwdr+rrnxSkv7Y1g2ugWecnwpv+sk8I3a3GpjF3P9486oia41+9rf83zNIJY
64j2/8LIWGNfg6ZCjrv33sGhlbvFV4F7lQOn0hvDrL9aygp6MHdd6/64sodVjXNw
FG6ECHSKnzUgyHT2/fJjlsTGV1+7uHvx4NINvqnkkBOxA99vhbWYTpbFWLEc01q4
PZb78mWa1Sc+KKpUutuXIfcCxdeKLzzwxez/5Lve7+biznk8SvkgQeJC41ksmcFW
cf9rHwmDnqnJIrc6xbxG+2UyKtF1f3tdsnV3Fs51jSXDfRpvEz07rHT03AnDR6jp
yeSTjn69mPLZkLph07Nec2Qiv0b6ZqeEjW5fioCseD0horfGc9feXO5PlnvvBvh9
KBZXC/x3S+iP8/38v++Znd/WyUIYtdes52ex010tkdk44fA3r6ks+H0ix4R5eJKt
IWxEVVo0qUHzu+9HitNJkdYz383tM9S1uMvnS5y7xxdmuO7r574wajFsDiMwuWX1
b5+A1SR8Qu0kBPwaiJE78PUhWOmQlhsRH2fbzl8s5+cc0s0ORokSKU7LbeRUiz0E
8Pd0jFkDXufWLJS2bHn79VA60ybDardz0Q4rR/CYknlfbxWBSjZug+WphGZdiXwt
hpV6QGv5y3KhOzAT6LXgnk94m5NHu8gFlM5/dfIkV01U8yCHINXZFHNepBbMoSxn
QjkP2oZE9W0rmYpwTGs9PqmSt11SqlOGD0gElcQqFIomgxgsnKRXcJb5WlqrNlX7
e5WpZnESVwclr0zEVHdnxad84Hwy0YQEgijyhHuuSAImMMZE7JxPD7uIPm7P4ehC
MmBZynk3d63W/UN4fZrCF0yf9SlzqJWJu/oo5+Z8vBxBOLpSsVQcuQuyOhsQckV6
aHozk2bRj45vVldlpuOIAgdmyVdd8UjLBloQVvhTlqJtYD5cqrpFe7jWmJBIhrfc
EVVbeViUaEuDMBomHX1VBUvKRKuJDh70fgxKpRBWxS3IrFRU5GVkBGX62RLwJQzm
Nn5Lv8fioR76MNIscDqK1otATtgDPGOiXpCNiooendTMklAHr9b7g0TFwUupr4rb
JvZD6mjRWhPuHu74+5ElLoDKvnhzLUhUk6c1ojoyvBjQAhc1mjd2IO0PBifxnr/g
GQZvjkDjOEAc/YJze2cERN0LOu3hsZOsBBhS0c9v6Uv5o1CgeQBlHD7OiebRA/TH
8dSHj6Ct0836OqCiaopLmUi5iN2YZ6vYCJWg9gKiwZkUXPL51l3cvsOXwXcPWRON
LTmzO5GwaaG2IgyaU9wslPsBpBI0BHTco06C2a51aE3NUlr66TnzmL0ahnWyOgBn
ZuiD/7e3qf+DJziA0FKCzda94J/btujCH4Px6ywjt1nzkDJh6bpTouNsDQeQ7Vgi
JoVBKccVY1wK6S/dm0cHqNCwXIXLDq6hGLo3LQikhbcCwjkvT04KhuHLUny6RY7F
pw+jTZn6R3M3UggXxq0gcViFU88YZ12/vUwBg+AHmnXNh8j5be+rmCfJQhNp+/Ty
XrR+wo9262fcrHj/my7FqKDQdqUr/pvqAgWcDHSULtflA1X1P4L7y7QPej8iL7Ox
Rr4b0X0qVUGqYRtR1kpYePLaFNZQo55mwrJjkPSpaPXp4wCd8KVocqMXhpH0FAgP
Y3OpMdQnDKP3hOczLTIKKxaXN9HZH6fiRPOOcYeiw3SnqIdo8X0BA2kK/bKBIUbN
KxfNnwCZQBSAhpIpEUcelszjCM8vB/2bFAD3FLTU//3608jjPiuuWtoWiLyMB8xZ
yPuzIH7G1/GCAMlqggN/xmcsIl1rii2wAwmkBe1Dq8sk5d4UjVppXdonmSVRUPjS
Rj7Obh5AWRsODnGKfLh1pyCKIb3A7ZHLnSDSOikl2u9xgHb0ah5DXqJUjtI83hF+
4JiUNrk3deD8y/R/eIFyisSnks4rr5D3uN9ycehOBD3lL3F/wCP4CzfLHg6sbiRi
bwgCaaaul+b43/2Q9c6pwtCQv/o5UdnIOrIVoA6CQdWiYF5vLKfJ8TBOC3D59KjA
4VAc5XEybh/fEjesI7OU96r7Ouhc/k3Jrteor1YeffBp7jTErBtcJ3DJGEgQ1gTk
JnnlVOdca89wPx7UzS8BiRz7WDO3gUv2wnzwxrkKXZOWA3mvLwxDB7BKkr+Gto6f
0Rsro98Ryfi3TzZYiaWo8g==
`protect END_PROTECTED
