`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O2VP0v5NNn/JRpd/w+BM2Q8Awl+w62kWIQXwa+1GERTRpXn+txPHaIoN4E1NrZja
ZNd4XsfoSaiiVlJjgvn3bYP0YIb/T5WJSI+ZWdpj9+DpWpF1j/Oji/F1tnoyfGTg
QrNiQtUPgux2rwv+DjsMBsvyRsREENc5aV7XoZqqO9agqsU+UwZ1C3j92CcbqAf1
cLMjGWx/558JUM27+h+hIpecuywJw+zB4UQFdr4a6TcOXarHtgRGg+t403HJnSlu
cr2rbbK1V4lMJHK4280nRTFbLOp2X5Vny/1Xh5jj5PO15StBRtfDFsqn9pthzIvc
/XtUMIZhCgzXEuAiuPFvhxRpohK6EnQ9JHJmA6OQuZtSqb35ybX6x5AC3KezVHNM
/KdglmV6dw3paTPsrlNjZmITrPgimsBlwFk9QrEY9JwdnDVC98mB8yMhDFKEd/8g
g8lRs6ijHXuMj+OnnBEzSrAn4If0gbzI8xCos51ChCSg/JR0BIdSu2q4ZsCHi/TJ
4k+K4eaZ87QScBH6Avb3Ky8a7l1JoC4RZYBRDBzGZqK2t+mMyk2BZwo6oFvWgjDA
e50im04wT7LY/8W36xl/14T7xNDwXNd9/eHO7Gdw1utxI783bpwwptn6UA70YzQM
66p/P6B9JdlbkSJdj/PVGI9gmEckLECwE3PujPikzPCqO8ekDxegqnwQ+oxxZZpH
F2S6eqARlVMuviUUMEeKGFRkixFNTbbxGYK2kXvqBXKefH2DFnl20oerv8IBeGJA
m1t8Z1yayUDCcZ6cA+gvThxI9ydG8DbslZ05TJU0uGaZpcxFuC5gzzUYUIVGndld
a3H7LM8xCCC17YqNA05RNauvEkJ+AMtUwkH+PU9l4aJaqh6Q/NnGzy/sy3rPDhQT
IbbjKPHrNv5T+fjSHci5ZT0sXmkAHsHoaDI2JrY50vxt+9o+bzJCqVB1hRir8UWd
c5qkZ1KHKp9VGvhAy+BMDkVaKu5lVYexMdRWylVbR11mRCN+uChGQjHh/WNJi1aq
VTqa4rulg1FwUwdS1ADl7uog/iWmdTgY0sMK0SGHWoUjR64REL1w1YlrHGf2sbbA
51NOPvLEZu9RHZ4PlTKc5xFcfMCcNnMSqeUo1ewW/zgE2Vknm9GvOMhC3/PS2hm8
9RYe7alA3f6lbkIKueTbfemBNusCENcPxL0Fr6p4xJvF+VOxscWGBDnuJvSyokRp
AfHA7DhfB09WNrO8CDBbZOaBEdv4tjnUWxb1gP4CQXfP3fn6l7H6p97i9iC/IZyl
Hzx/Fe+lhTaWnuaf252Jk+GfkkdzEfdSTNObTTKSHXGQzGY50PuLnujd8XdWKTzI
lGIbmihcD1ZOojG/TslmpQ==
`protect END_PROTECTED
