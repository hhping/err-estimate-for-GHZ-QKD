`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
akIbTl0xX92MP2pxyMfYhVfEFj0jP7mnEU6JBWsCqqHaaLNC2I1ub6W3o1BJ7XPc
bTMvCVpS0OSeRlYqxAoC+PNxoRObM+9SL+d7gL7b5HiRK1I6qMhsKgli0ppS4b6Q
6Fu0c1vfB2oWbJ1yfHpsLNYtbU/1+9mcAteAVKY41dZSHDWmaxuccx1VOf4PP1eM
edghrFNo0HPNvNKFzB6yD6Za1flPY8yew7W/57ve5ftT69MhAoG3yTsSkXAWaSSU
sV84xYQ5o5hTS4u0Z7IYk8VrrcYkuJVxdNx3L7gm85oJIUjQFLkua7tN7HeXYBVg
N/adKRrkOieuuu8JjEbMxlGCQvSj/N1l4cV3ntQUMiwgFA0J+bekgN+lzl3X7RNc
oIpn7lpvEUdfxRTJg4Cz91K3ifaaxPrtBonpqgcWSV1VoNtZtwMVGrWKmnTTmG/9
9S4z7xQjOMjcKZrZN6IT1Utj9z/YpW0ZNhtZgNyRCfk/MjONEtsNQb6mByhK2u/Y
LWxdxW+OZGcaIIkx+6Ri/DO1h5GBrjZX5cCGqsrO+Exj7wJK9y3ImVGPGnIbWDpe
l+/vKpC615HkWf57GRTDsRA/72vMM+Dv39+6ctBmlnVIB1Shz3jt39s5/D1WBMo3
lz9uGMHau0T5PrXgwZCJXWORxNkrMMGuhNk25bt1m9hZUXaiKq9VkyckrhAUDkTO
qKTwwENkBM2UVhRML7TImFrNRyzYaMeAk+OH41GCV0DrR1Xbrc5LkAIx8Sq2ulYv
X0f++VijApnzxzjnJHsbMVZRf4m9qNvR4av2agBnk5sc7Lrt65ovDkUTRZmkBj2R
fyhb6x/wQfx8si/x42Vo3Ysz7aDPUChjiJ9H8lBdAkXHsjQhtP3OKzBSG4/7/w07
bApdWjLWJclx+zpSDj6pEnTygydmpQOkv8R7HPIxB/JtA5QrvDueyrRv8/inZq7C
XoffRBX2eFFIXAv0k10ouXzWfirsdslj4myy3Ot/VG+jfESWTBZs9SqnriD+RkqA
P80zazmex5ciwh1yJ2SWgsqAEAvdHN41M4Jw21T9gfcJfXF+FLjvGgkdbXDO+JZz
RXAWQHlWd7JWGqfJ3FWRit2G3yx1LQ9g6KFMfiQzy2wieirgZLD0lLjW1IIZy2Eu
USzKca1DO83p60ARXQLP200XWtkhvQp/Aom2Kj98NJ0jt/EM26PKCo2MthzrLgIk
D0b8gUps0zwW68MJWbszQs3VfybyFqjJjqytVUCl+iQpxfHN7D39RDdCANDdcMGe
c9JE8GuEaM5HsRpc5gjLW6LNjX3rd2YHfeTml7u5my/pO+zjN+hZGa6g3xFi3j3I
ISOCwiKK+Pdks1OP9zWkEb3qRu36Xl3843GdpGRT9ZuLnVoJVchHtvLhcWa3hmnA
AEi/6Lr2mpwg0bqWUcREdI5FPd2LKf7Eg4JSAjUgznkNbpXpsWf5rsJaOTPwfxUT
GGaX8ko03uqpdZ/oP/+LLdfMNRGXv9bT65wdIE/51gGO0AYIczi6cOPqliyqZLyO
azcuCmdwYfLnZ+PABiczPI4eus2idfHOAjBmEpB9mLUBcP+Xl8ax2WalhBMkK2pc
Wh1oGvELyAavax4pgAhrVoABFMyTeXmS7kahacHkUDSVL9Q2a0iyE5vJE73Dx7nn
dsDgkTs6GzNovoKeGkTjMNi6l8tNTzkogwXym63g/oEJbpwmGGy9CHnI+P9bS80d
LiPvpmy/n84Vl5MYZA4+cXxA+KzTYM0Unb0vHrdnaW2yHaCrkgAJyrV71oEwdQj4
3HxYs2NtlSixCzM/eRYt1n1YteWezxcFNE1HDVsSssFCEiBqrWwcS6/EUIsfoGHN
bnl/iUbf/JZ84v1ukTij/EbC2MaucsjBKEpI7I0UGQ2duFggXF5vvlFzBY5rN0yw
wpb7Qx2OOrWimv6KKE44scGD+NIOsCYoAH1I0OX8yFd6q/7gtoum+dwIMI/R83ys
4Cgo/dNR+nBsTwnR03nvvimSbd72ofPIECvUqfXU/+aoc3BFNMVB6yF6X8mXRZ0Y
RTrw7BxiAgjheGAVLmB9f+UUyx7VWoxNLeYnFjAqd+DPS3TpORhEs46GXhAyEKl+
rS3WpK7dO75yRf0IxwX0YvHVn0vTQxv3LvQN5wgNhe+TAiV7Mm1gTFr63C8dUKMQ
FNlu329SfWYfsiSTMI9qYLUhXSIqN5xkh3D7oYKYyPJipBKitsEVKjwNClHE+9ml
YFpYPdRZUzj8xPerJOJn7wdwwbmEmce7c/3GW3nFptO7gXeXQmjjI8dn7LIUP5yp
uPJ+VCNIV9OGTyhN7/DP1xKUo4JpvQEUWZ1clAA2QFm64lN8RoCLFukipiWD4Zjt
JFUyaO/g70Pq9oiNRWuHWvQJuZ7lNZaDEqn7py6px5Qv4/1YclUoK4qKyxPBkH/K
dV+it3Tvip+Q2ODYPt4u9HpsWf7uIKf3IoelDPT2Ye75/hOrMpeqFEcLJhcC32no
Mnj4B5kqjVh1jaEPaCb88PBnu/KhnZ/gDr6IjafwmUqsQfA1RdI10OMHFCEUxllv
/R2Kn/ckvI4FDPPCfmf9cYHlTp5vlU04Nqc+9CU2Lw0GZntgPhvXgxk608odwmRA
sU7ICGADdDkqlMlN9FPrLw3hdnCxkh1tRLpu6DwxmG/V5R3XD0b6ias6Dj3Npfu9
7OGCgCpdrdK+bHsYJn2lRU63gvmD+56Umc4jCJEQ9CFX3q3FmZxlTJ/nOy8qT9kG
auZiX9jAcX1NBOvhra9PXDNsfGbLMbTOoOM+mixE3l5gFPVb2l8pQ9NZRnvFubHw
SlNIbiN1gwNo+/xoL01W+EljUB3vq30LxEf6btWfZ75DWC8+1du0TtPVZUYOPElX
EzleIobLz9whhsiFRB1bL36wroY1t5wJT1hQY+jPwaoxfXQLioUZ9O8uZBwzQWbd
tizoqPm/f1L4VLdbo9LBprB7J/Z8WMhi7Bd7wjK7lkZ55Eu9F+IPzU1gH+Ytift+
+smmDZGuvJAGSygqjg+oxMeO+8rHlooTuYQsjLJ+A+HDlbdF7OMPbfaRRTuW1gLx
wZEQ/UfU/5kTPQrPsZdZk0VVxEjrtoDjWXDVyZEChliRFU2nDus+91/aHhZjA2Ll
lZwd6Pb0D+DVvOnQvn0ZJrVBAuBrHHVgaJrOW56UnzkRVF+BS7yRszRcw3veMMKD
9a4HN59oz3em+3N9jJiw5Ff6dsCDEpjaqzZsAoIwV0ZdEwT+6QXxL5Gn61smbR77
aWYHhzFVUlajI7YuxNNXLNMSIJx4Vzp0QnTRTHBF8RuZv8L4yE/KDv+UTHFmgsSl
V7fQZ+sudUkssn5qn2T6RYiwkUjWo0UIO3qgBM1J1iB3MS4Oj/+DYCS4MBQWDWLz
tiY/u5pnXqhFFzN6clNQMCDgsKPuGxAcMhDp5guxUCpZR5Xfgv5Egu+mSzGgVORY
lUjNR6Jz5McJCeEfFq3A7IxNicIJvgE1gY0IfS2Ta12uxyzDZ/RhBRpryVhlW/qP
wlXL97oJ3TJAHu+X9WDfxkd8ElKiG3i+usF9Cy3zl9MnxCXVVhswd0N1wMA3cRV0
VngrLjVNpfgFzdQHk9hByWli/tExjK21U0ywxLDel9m2KGBVnZuSCvuZHIdd9Ey4
N14ZGuWpbRWjovVMpl62Jk/i0JKhy6ASY1JfgP+aHx0u3BBX2R7jR9WqaVK62QiH
+Pp86j5MTDnEFazaq1el2NCBj1/y09WfbpF1SBYvqyuRU8kSUE2MfBk537/lAr+Q
aXASvdEY5b9Y1tOd/bVwX9zryeNp+Jv4FcYX004mP+LU20B6oSX7DszdoVQ8CwYx
F8laK+DotFT5owJfRlegskVyECdxpWUb4ceijmGqW/KyH00KFibL3wz2WnZnpc3u
S9z05JBZjcmZ0DvMt1/kVw/uX0yy2pWXvS8AcFol/m3Q6RAgJ/QU2stMElayqsFe
7AxHR/Oy/dELBwQvNm9klBiCmWX8L/K+ZimIuxtJGrdhBED0RlBzxZK8ASMJau8l
0bQoG2nEj93FW0IaOBpfr/A3Rp/PBfiezMYwlio4fvSp9Ts7tim1+yat+Pnqb661
E5IvKmjfjB3sr3f6/OlhJNjqYiF/F4Hs6oXRIBGSaTGEaPazNwS82+JGWaCdKVKE
BbV6j5FezMhqQMqSNS4R4V6RQR63S2dgRCMNl3o5LutR1E1Zg2fPtX/xuL/jrk2I
cfEydjeKbC4e4IyFjLbIuwxLhiiPoheqlTmvn+KzKiNkHFCwI+pR6mXqDSf3Ol0I
dBs3hWtas0yXmDerw4BiBA75LsqNsQ/n6bofqxB0UZx2+6f3Gm1kv1ufNJdt9d6z
Ou6V+rRH06itqrI18evpxDMac3IpUQ1r8RevJ9ZTAH1GNuBZMOI3K22gdmVbHdnG
bJKMuA0y0vHly94BL1o/utX/bKjaBMHwp8IsFLXXumAIWaLz3IfIzwIVH4CFic7g
mK9oukuJyk35PasUn2SiLqB/rlyrRT+wBClWa8DPnKFba0acRHxbT2QFiN5LWsMe
+2N6BVGXBCiaK3OPDinK0yoXfIJSosebgLI+iDIlEl/R/gl9LwLc/4d9R0by9YIB
NQOpmJx5Att6OSVPyKtEs5d3v90QON6NfwMQkq3cz2cGw7f7Da4nHxnIkHqhwczT
h3cT3MYNZ8L2rFK1AMSTaQ==
`protect END_PROTECTED
