`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tDrWAiLQG0gqXCl7i83GkATo7QZmce1vTWBo4aXO8uhK7b9k2ydDnx8zhRPAJxRx
VkHNg3bKa4FisXl3fCYQrcDrwFsaA+WjK6uLCoHk4YLRI2xOXOBVNaCqOMZ3+b8/
nC6mv3B+HIJNG7xDr6a4zLQZ5LcnVxRr+62y6y/qZez8mNkbOXrDJ1/1GEczL/Z+
gEqrH/OTIOovt0gY7Mxl3GQ8y2b0dM2HV5YLLPAANEDwRR2QBBh7Yf69/09x/Gr3
1A+gd1JiX6zBB/MQHx5//Cp28TSYqksu6I1Tx5FhweegsjkvKPo0bSJ0oHzLo4Yh
4k3mhi1OQN/tH68F0HAMItcm2NBWMK/PCH3NJ9Zsp2QODU/m5jAXKjsZmVGZHLu5
SwAIRVeuzFEr039jZ4dLLFFr2o1DTikwv3J3TUbZYAB5WU5ZnjvFD+sQYdLfrA/q
B/2GnqMf21BzOwVSIeSmeCBN9iditE8oMmfnLh22aMDdeoDlfy58JNQGoyae/Pxm
ELlvARRfW1CRroRF8zKGYgAZakfB8YEn3AzY55qzHjrkqn8+OW+IpOL1rS/iiv17
sbSqA2GZwwM2LvbzYfpx2TLguTZKlPTT1w5EoLbAR40=
`protect END_PROTECTED
