`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m325kmb5B31l0aFb7moBWhd0Zg9RLNEujh1DXcPi8ztQsobBrKhoBNh+zg8RwMGG
AFDevYpN6+MtAHHswgUfauqTWSHK+GjByj20fGbJBM1YeXSXzm61cAYSzNjTkiVe
KB8XIOWpCq5NyC/4VKZ6OPfSwd+/85Y6XlxtLZ/mrwvPpsPprbsLILetF378bkqe
fBJGp4ljF4Ke1s4hONILCoqpaVg84qlMHEE6J/hnpAts6dIHUvGhIeiW1SmszU50
kEiSeEhLUWEJ/BZ6/xxjAdf8Yf7OqXC2G4K2TZOrAt/KqsJfXgOuPe6FFLidaiiI
Sqd/1DPlLC1AQM5noG8N6N1qkr38wGQKlCkbE/MQnwZz5oCj/KtXff0OgHEfVW/B
3CWSXB80j2tLapgWMfWwSyVer2BZJ9lV0iWG4ywps6yQ122CApvLwpMc6Tg/yPv/
UD4uLWADw7+N7ebph1metXM8tZm9NbWfP3J7oR/5EnIk/oGht0NrqxyxAsCLSFUs
IJn2xj+4IqrSgJZdGwi47uZtRlDTZlMlPoX86rE9CWX804hMZhKgHMIahVHaA3uV
Tp7kBL8VKwlinj2xIFRh+lTlPow2DBfAdcVFflx2tfQIRrfWTBzMPkWBairzAQED
rFlJzmaVDMWZuEvSpqS0Tz5xZIQc+1OY0rJtJNP62ayuci4dp5BZG6nAZvcWsBni
jzF1mfmI4h1ggggkHKeBEpA+lsHafXyRtUH+/09CVCA=
`protect END_PROTECTED
