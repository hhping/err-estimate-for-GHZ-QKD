`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9cQdmLgYtanMNaWqLpCsbmp7s0COdbmuKf4aMl3NrbhWCfbfV/4pEBdvRcJWYDzb
YO7hsAtAzB3o072vxuAnI2DKtq63dKZC2DWP2zrctdimjfPTp+0e3AHGPRjZjwXp
MRRzgALgUDMkPyfbOy32PbN45UL+vpVjxFkUPQYEp3dXPiwCFfQrYUCyaTu9Ws7M
esgQqGtsKw6yfH7i8p6oHyk7MPfvioSOBf50a0cugWSC502Mrzpn4z3CEq77waPg
knTxwZozb99g/v73cB6SmZA0z6Aprqtzp5+PV1+ROGrnwELRIx0nL3uNXylVLmr9
6SZrR9THn0rjde3mh3TeD0b0TZVM9awWv64Fx28yIlE+eE1pj8awaX5/p8Vfw/3W
KFWrqLkq2u68+qlItdioqRdPlQz7Xjrwv5ZbCzwRKW5nF1HGjo1JgOHyuFvk8die
XWNeOjovR82hGCRVTMJFuXWOBm2iX9mkpSjFKOOehzSMvUKO/wk88BX0g2eim4TM
unVCXmJmHWyaOU43l26eqPTrjOCW7yWhfdBtUNuaOchwhdIqD6qRqHZmqtZEVMHY
Fq4hM3uguw+phFVAnaL/bNvxcuPmCZWjC9XQXi453Cu4KNLs/db+BNPjuhSM2xZZ
`protect END_PROTECTED
