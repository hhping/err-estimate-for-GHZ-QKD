`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EDXVpk5KwM5JdShS1f86F9UuqJJeoIFDo1+7CSjX2AmSl/3zGII9GDoNOPrrdqSV
C9zqPlJ5CILhfHVw/MoQ9gb3RZdV6qjDEV3OprKdWmjjt22wyBg6V6QWk2IA6hb9
34fJLkWiJZ988/66eVtfNmy8IAsgkqVarKx8S6KTq5h4SCdpgCGxvBAw+n/cnzta
AqIHUe4I3ne9GSgy2bOuG9QuCMFiiIFOiYi2cSLxEEQcSO0P8igGv69TBJTjdvrl
7V/O7/o4LrdiHlkQg3d6r1NJ5ICSuGOMesrU8H+KA3JCA2SJk9MxaAFYG7A+Z/tP
ctmGbErDpF9sMESAnxFEu0ABZINUby0SrAoifh9nq7184eL9alpStZDLYsWr7FAZ
BRmy4obd3mO00akYeZDJXchRC5Ki8ZI2JrdV+TTCgeOyMjhqNJICysMtfJLWXnQa
R4Po1kCvwUeIXlpDL7BkDactmGi2Ol3Ykn5bWzXW5gVQatvPp205NMSjl+YxHBFR
kns6g9kJ4S/K8TNrj59L1ZWxWKKq7g7kn3qhEVLH6stLC07G6BC3AJ/ZxJ/dd9Me
4o3PHrj1VMiYZKYISgYv7vJqBN8xVVXhd62M4QVloM0Zb/QRP20BBLS0zd8WpUZX
OUWjKbXXlmPYXofx0w/2IudegULL/XPPArAoo6dKHkbE1KFkezOA55z5qfnm/oRt
fWhnnBSDjAx19g67xyG0Cn0LblehtzIA+4yfXosMeDNRDBVAusp8KTPCWdk6dS1A
eiX+wvjLRCBhjAqZ3j7yW2lkvGusQzWKt3yLecxMQgt0CHvJGdKQU9PDtegGHVsY
U6ip99wHB1CMzCBKlKXE75jIBuSVnEt7mF2fejAD1kGUTVHCqBVPopdocEIqwfwN
uSXkrGvZS0uZIYnmbz8hwKuQ2KCVz2chQDUCylrY4lbyRTAc+QxFqYUo5CPJdg/f
5NJ+ryvy+dtdXiyC3UsnxNsqL4L7VKDRgj8S8DqBdFhMEQ1aVaa7gzE920LvImKo
dq0wP51dDk1U7Xh8VzUl13fmkFkC3io8dQnrJIsQJMmukTQrawa1xuC7ZEaXWds0
n7GbLQi/tNHYyRsVxeVvZPA05w07i3zHLWjNgXb8SMaPMaq4hQZqrTfgk6KbO7XI
zfeG2fQI3cLcUXAmoiKKNUFBn/Im5jYiO21OdIHmZ7zIwdQtqHxbFvklpArrhTYt
UderolGHJpGh+ySLAvq2r1smku1HAyuCAQAc52ayROctcbhIKoOxMPs0+RcYRXYB
uKEbuc17G91wAtieMUjrDFQJRD0JAY0keP56hg1srrsVyY9Ag1OQO1BW3qi9tDx8
qRikvteNa7u05MKWcCqy+iGFg1L3Ufe5gYI/cO8ceW0L2umqAh5xh0gqgnqsHfkm
pAXi25MlhFV7Ub+0HI4HiTq/hqiuIZcWqrYD9rzSayUK29VAGEHzSsnaoWjc65mc
KQu9kNhcJVW5KY5wyWQSk2SovpTEnx6C/jZUV77/akwHNOrP7L05x6dHM+u5pynP
6oO/nB6azFHGwTTOzIBRkXol/LXLtKDCBbkjz5ecYLc=
`protect END_PROTECTED
