`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oYB87iuRJ1kHWb01/r1B8J7NnnY7bm/uOBBG0OeDTCQVFkZu+czyzD+iRKdnuCc/
lynm+E/7sfz1dGqVjsMRbisDr/pqYcgq56OlhAIZnalxSFH+D5j3/3as4AYE5gXG
a/MiIPo0q0BAJ/q/K0Pz4bqnWRmDjZK3pApHejpj3mxmJF4ghULsQdh+vCqWYrk2
XZZv0sYfwRffow8meqOMuVxlDoeKRnxWOpmDzl4Qc4whdyCNfktj9G+lPm30HHrx
x5uOeTZGfI46qqWGpgqlSnIlAc+aqz6eMkDT044MHpuqyHXhZ80DxqVN5v5OAfwX
ns+UjGs+w89oIynA7zlKwu7R9RENiiEFqecUXPx7TSHX1mdm+xQyt6tqjWNwKZK4
p38daZ8yRiwtu/OGKDNM4Ee7CeRZ2tUoUuJrypfKSnROrezIZl3daCNXE4P2Po2i
rwULakbdGS5zYRfjVzv1I9H9QUR5hxZImzZ2YHq9PJKJ1VnzDTHE0IQsVgVO8Rs0
3VZaKnRJCLV6YYu7Wz3/OpcXsqhqN1evt+J25FH35FLInG8Lk2Ovk1qtkTgSLISD
IpcZ5Lsh3b7KG65GipL3JMr5pWLp704FfRzrsq4ZeA1swwh9ppL8o+42YAPiwKo4
`protect END_PROTECTED
