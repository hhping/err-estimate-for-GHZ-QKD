`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PB3cC39OPL2vDoeYlVyCdA1x2eN/kp8tQidrEi3WBlCPA8QbewmwiZruuC4MSk4y
WyaKhBr/rAO04wC/XidXwZrWkFQisHUfQJs/1xkfSniYc5UA1BLv8W5NZbmuDfbj
MG1/t/sE72/blCGUAnXtrnWRBPOHfK9h6ingwbL6uE2Zar7Eu5GPRwgGMWLsC63P
Vnj2uCbKpwXnpYQGqSQAFWTPAvxMYptKufR4IEhtweC0v/T61V9skNrRQTS1LdcQ
GNvL3VnTKHSPLuDlTY4dfUwdvpkJbicmEsIM/3wG0c3eMG5W5/SxsTJN+v4Wssfv
UDZrYBLN1yJJ096m0nGMUrwW/zWy4ggovbiymmEIeg/H6h3PtXCy6EJBaljp94MM
/4NhFTB3OSohFRCCFrp/WLT2m2I+r+HfB0y70ExJM8xTnSYSpdUKL5z9zmPxrpqn
n8sVIc31e9nnVxBWA+jPbO2F+b3XuWLwMFpEeUsiUeMM28G7j9b0m+DJ3qyxi6E/
KaMp5j6+5cJgtSZrN0+c+P2cCOO8QEVtlppduk+mbsQ1E2GCyxKDRnGoi3QuDYNb
Ylm/DRSkOM//JQ2l6WkPUKkjcBN3/6aDm00oXpEoY15uO4i1awKGeyZc22IAAFND
R8RSo8UjxtnaT2eCkOi+g4XHi2UpmBLFC1F/GTns48yC99OxEJmj0wrRQDvqt1qt
G2e8mal/sWWW2OAaHcVGS5IDNifaUe61g3jHyERw+/JlNBQnxaAgINZ73bS8NW23
z9+OR5R5jsUwbSSgVgyEPFf/VCFaM/bB8OSsU1rQV/ylBwKDGIi9ddBl9J4DUfQS
Ep/r6iXrFZo4APJrWEfqxSZVByecJeWTSndREK6mFtQpCXrPCqpZdW4BmWuv9oDi
MxnZcf8dljgrFekYy3OQbMtpbfuaOWJFmXcue+4bR5v1o5mPvWYL+wD3gIUyrIY0
1d23qrEMHqkk2Xfga2lVuLW29q/qfEhMXSzY0LOB94bKCx3p9CNv64LfOc6knGLS
qWBMGSIH4u7JbAuwE6tDq/foyPHFxSAki6o9nAW1SBEE1e8CWOgaXYi7oQIUcZ//
EeXANtTAPphtj+Ks1jlajl1Aidl1xUeAM0AWpxLmqtxjgiDIqi5YFSnu9KVCZaZk
qzjoQAgKvGrKTp218b67B0hnuwywG0dmp4SPTrm46tjrwcSSPgjaQCNEWV93UEqV
ovAjGK1XTtnfF+/QiQ2pVdWLyHSt/2OLG132Cyn/T6s0FTPhMxGBfoTdDbqbjDZy
H1PlCmILYosJcWGbCKck3bUCJtXwM9fDM8exeAs5/PC1WVbuO/LtiegbCvr2vM0k
kGN9SwLDgmWv6aWXmlgck0pEinDUl3L4sykZbX+zQ+HrSdZknM/JNraApzcoQfr1
JgSFbwAGBu1jxdsKoKfFbZnt17edEBm2ZozG6axcv+TSdiqfPq2yFV3ZPHFF2bT8
tMx2+SkvdHe92vRSeuc2eWPDyUifd7OPpiaiIdX8KvBvmyn1zLKS8sjGuzXBTcJm
OW2YCnTSz0MNRdu3dAxwsYVfqRdRALREDrX6nygH+yMsUyPzmcH9EELqwNvpbFfS
WcKZb095ckMc39X+ohq5CYnhCU7v/FbjSYc8xrcuu2p9u3DM5Cg96or6rr4bIM2T
PHMC1mJsnDHEpgylFYN97NwF9TgeaXmFJAyL2gVS0AjlkTw0rbKnudi6xoG//WZd
Z1382o10E6uu+byZ7bmgzdeA8zYhUIIwk4ADHTpg/XDSQpGEg834YqN6hf9nOODF
UeflT/dtycG796jshZnv6slhnp7xGYRrTrOUioVKxAdSCnfVIpEtR2+yBPsUNFJl
iBNA/BLmWrGOYjtqfOESZsC28+PHJyv7VLP/infB6ed1Q0ayGLzEIgcQ9LW+0fJ8
+52eYIVcN/8sVXwfCysu6L0Cqp3JSKaAOTLpzYbfldmAZ5rhS0QwlSQES5P5KvJm
XH71ryXidMcfsMVTahjgmCpLgvtMKE4gvvxP8lMX1Aw=
`protect END_PROTECTED
