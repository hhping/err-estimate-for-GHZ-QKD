`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NOnnPTCmNUVGDUtSGHsPhsMTkahPFEtXEiLtWgzFjKYcLZCZi2qwW1OSomJ/i8sL
C/pgeeDjbu2jq8+uBRQ9bN3Cmaj8VUJzDNvar7b1bkYJQ0taJvE6kkiDcaMIu+TO
0DsQgt06xJPlb9deLx6FTnw9wQMRIvDDzTntCJEwsviy1XTILnmT9iR1FDxr65xJ
sCw/rFxOZojgqv2/7vv+x3S1v7RYZd36hbS8bODrASIeaRumtQdexTjCLEpGbHRj
Jg2Lt3ewpZyCMuKKmljp8FH1BU/GHdu0YijBSUqBVj7HcHEM3mJteYzsktoqzMjq
9uH7F2ahqgAWq+DADrhFMgwkJS+tC3TRvPHNmnZlfytOcMgjKJL+4QCwf4Q//bxk
MIDzrx7bTdvBNT3r8FDt2VKhor6BurQEmhUZXq4Ihks2QQWhjLOiA13BrijWbniq
8Hrebbhf9vISY9Jpt1CqGDnUicU5n40bgALJWQG4zGyJtLevdybVFNnbDVYJmkX6
KDioqann5t4/3Gz0niAQIRBbJ+EEbeXO1hNjn4TT3cWo8V9dP4Q+uloz/1YpI3ND
2hKG2KXshexxexCtOKZA4IdDoKks3VZrvI3vmIWLzN+RuQga/OUpaO75zEfssKeQ
Q6wx/99J6MiZlW7Au3XE3rFaVoRMtB3YbZs8G59IBTxAtLTFeTf31AwulO53sg/o
+z8ToLvDny9PgbV7C+Pseg==
`protect END_PROTECTED
