`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I5PeqANkfGVE4is07yAI5OpwZWKMqNMdfD4ozzT/0UadTt6gqAXkxvGC2YV6OPZS
MWTZpXQUbT43cZvUysznKqFcR2z1GHy1f0PKw7McVGV6MNQY3zvdRO7WA2YHJmfq
cYUv+4vDlkeAN2Jg5VI+g4tuYbwNFQaYK8PBB7LsAse0qnBjg1lmfTQF2u+4gtv9
tXEwt7fLAnnSGAMXqWetzlQYQV2/r7B2jrUIt0AFKD+LrveUdiRvADPfPQKbf+zy
o+UlhcS9ooBL65gUmXTsegFhZ6zj1b5DpLA6hKWoxSjJNWu11Bk0cJtJ3ZkW1m3O
fv5/5LxlsPOFHMe9+9p50R4PD0RLxDDlG+qZMX48HrCypEGfYtzF4KkhCZPeQqey
6r0FQIk0BSmZ/TtFvKtyiiFJeqJ2/27UH2HRDx3tjm5jDr724Otkl6SLnUA+6TaH
D6Hx9fZvTw7fUvlTi+bbNotPjh2hrX+ZrErdG2E7KLG7H7Vmt3x0XVYcDT0X/8Gc
9PUhP/aTRH4ES1otYU8GtUOJJNSuxNxnml13mzeT/KL53mPPUq9B64JPtgkD47pM
RRaSppF9HAhmXx8uEpIzCCwtSzZ4a/a1EjFJsYIO6ZbuBTAqkRdF9QUyBgG4y4Zl
`protect END_PROTECTED
