`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g4WZaD7oAkGmY0F56Rcdp1O7dMu8hrlDTHL9quIb1OiETsAUENYNhgjl9X3Khm1n
a3yZiqT+iW8a/TLPwkK9DJjor7G9fqHPA5N0KlfYpEJF2hEgvyfWY1UBryJwwjNQ
S+xneXt/sjckWOBaJ3/bUY+1QNUsemY1QesbVpdz2Qa0YXm/XJRJLUMSVYMA6jFd
mhZ82FqMLAEbWY8/aQ5dDVivTDF4t8Mj5/ZaYk0h7q0s2cXuvnSw9gv6OilPZ6VL
PYZJpGoV3/GyUWQEEqmO1kNZ4sTF+Hy0Yk8iRdmFL0znmYVNEGE9reuf1dhsp6Ff
Ba62YC1ftt1z27XZyRW5bEMHS2L25TcfA8li45AjiuyEm8O8gJ7Mk2Qm30M3+xcP
HtxQ4XWZ4wRDBIFTpr41Qvy838BoKQSje4q8OVAeqLXqoYLb50JBq1lt5Cak99JM
09iW1hJiOKPz43ogNYFQquCv7mEluJqd3nRNfvdqURqlc8tadsN649cbnWYlD63F
Lm1801KVRu7+atNkDNXBtxa+Nj9rf/sxyTaZ7xKymODYzIFLIJcvAJ8/pUpFuqtT
cs2KJYcPBb2+5kR338UbkYAdp/wibh5lBIL01QCiRE/nYfzbXGSqPrQ5+NtpwSuh
wvZB/zDgV9XJ9zSERy6dF6Mm9/OyHvX9darc7yckGMZVSo7tveA6/D3zoiUi9bQD
fzwrf4xJtDcWpPWshbgEXrrg6MdoKzLRdKYCzkw0OvGgDzLxcFXx7CCXYvlv6ABq
3uDwnuf64NRvqNYr3cm4POSQ/yHl3qnhUnvg/2Hbz9+/wkhI2cA+jStXaOD9lEuR
ZYl+RlouKf9uVQ+UVmQdNHBa1SFqAXHW4CyINkdKXNcQJVM3VtdgNIeZAZASSp/R
m4FHaku03OuSIdgbuqMLK9zi1rwuWXoI41UAiSPSS1EnnSts7Y/jRe+693CcEX3/
KettfeV0/oIHd8xzVT+Hozcol/fHMNXEo4S+W914xNO+jO4fSgkTX6ZElabq4jOb
ZgUtkQeHAHxuOji89veKIIQDhGiThHciQlJGbEdSA/Le7MkEOlm9hWPkZKIyaL7Y
qPnqEUCnpLgiNdqPAdJdvn6rfbqkaAhdkpDXaxXwviYw2BY4WOTlxLzLG+AGRjDq
hh6yOxHrp05/nx9sRSYgLCx+zQ6DEEJVRbvTZigjbaWM+HP/LSm/se0yECaUYmpH
0FE3lgYfWetpW4tezJnIT73aX6xbceUf+PqkR4eMcv57D54ry5L4AhsHsLNlHCfS
uBk5rfMv9O51ZFKY1CkbRiJ4lRjqjfZiYt2FcqFwt4e89K3Pdi/SiP4COzK9T2bq
oHCR2owdS0nFBRes3ZjGxnwa3hQRPlr6+0pSiklzxH3jXuZkB4rPQAHsZ54Lmu4f
i847I3YY9ulqJtrm6lmWGjvselL+snaUV2CXRyyHIMcQlJWzBIN63Kh2t0yqGEmd
hNhM5e9qoMYR5p4BOwcHFx2fCnYoVumjmIFmf1GFp3yipRzfGYC9a7Oy3PR1yu7s
NlpK+BL1x0n0Npibm8YtNfU2XQoNCdJLtm7SVda6x3+SxQhmE0vkVmz9hskHJ3ke
iGIZhCSCFiJ2WBOyLlIfmD1A1bIMfZpsJ0d2aZY6O4t61JiVwM92fmiLDMqPwVUm
RFWmlAHRGLn8iZuOLxXRFJ+ZZ0fUa/IsCuNTNpT3qPWQwQdVIQ5CE+MKV3+9lA+N
d38SJ+2uOSMuqPwwviG5RSezA0BzGf1aqi0tUd2em5hVCAiTodQqB/aIhX+MStX5
djMvFH4TKLI6XNf60xdHg+J44X6MdHFVfxyRVNSBq6+jpNil87hGlkL+cZb1fKot
FhRdXTiUYK2J6U21JNLrAzSResDPsSwhn3E7oPKBk/a5zmwG4a/LpDbCZpcI4tsb
+e9vf12OP7r9ePSKI0cODpqdom8GQVnRSM6JQ39ttLFsIJFgG+8D1gugwK7TPXls
midhs8mWXhZFO/FwsCj4vXTLX75hzZdXfESRlMTDnbWF6LFXvWELlNvTv8vmtT9E
fxcJVKHfuKLG+JkNvniGDeI5jtwQTLTGe4u0AMhmTp3FtHe9HxHsi49Gzs3GiYOD
ZAFXdIpqsHBwgmqwHB6JMZXRRIMlFG8lQ2LquCVgx028bv98NarFuJFk4KGy3uRu
I2IVs0VOv8klOgFqVE8Hh75yoKvr54eCChbu8ecFlDuLvAVgPdI9BtAMimxCRLzP
i8UgpCaSDtcFS8aHb7pGktHtcJ4kCWSzGnuHo/rsFwpEWzXBDFv6OH698CXoLRTC
bxj9lOOQ/GRSuBATk5NQfeuS7UWBo2+JSMFHFsaxSpZDT/QcyIcpYTjYhAHqBdkV
E/jd1HEVIt1ck+MAifllvwbpLWS2gE2Z4/sMb3FqIkhpkRvldzmvxNS7DC85D46v
vs8+CYTvjpiH+Ul/flPHijT8rAyZh5Fa8WgCeNHiM2+QHPOyOcrKpmmPDomkVPNI
KFW20oyAJLdr8TrGnXTpniL1BpLOEUDIntpNpXEdE+iWBYeUfDQzCNC6xrETyloJ
XFnJjukLSmh5Y3S6CCNHKoUf5hAUpeK5UMLHTh9R+UP5b6UlxMohRw0OYSdnNMKg
PJuWFtslMnwuiL9R+UQV51QrFmofcvZRgjccRHk2QRsS+logmrAfMb1VVCwz9dZq
qj52IY4S1aFnxcuQ0BzHIAjgjtt68rkbD5QpB5gBROVh5a1Whi1m2yK+mLkdzdI2
Wd/3eGEKZ59OKH2dnYfPJpaEXHJQ2PwA7ZeUzOAesP6JqkW5D0H4W8CSWEsWLoYl
ywGRB+qb4vkxG15kGLlTtbppofOprF5Ke7p94uEndD9u2DmkN9vo7gYT9iy4B8BX
VXiIAsSw9oZ4IbiuUFxMXHDuT5//OXqNvJwyfG6hSi9nDildHgtZQI1X560b01Oe
UjGCZaxZgadzSVHPTtycZOMvxG00S7qBaxk7L/JTuiadq+ZI90yZCtKB+iiUkZxq
xonulQCBbI728I2Nt5li3WINNZdN0j/JM0Rfvt5MpVkXWUyt2z+UD1XJrPxjVilv
l8pRD/PJENmDcP4DFzByFmAYNdoPuhvdDcPdFZhnMyX8KTd+b691L7mpaKfYtYHw
kBUwAzoqRZw9S1B+H+NA8w4UXr0ujoQLxe78WpTEcjQk4cl8VUFK+VRS7YlvuOxD
644MqylAKOCh7sEQ1QZ0kDJLw8VnZKmTBqq4xs0gkEVTNTE2YL464RmhuLftsKV8
IpT4xce9P4Nh8c1RzZQGR2TGq13H/JglaTOqHxjeNwD5y2C3iTDhX5pAMnbl6WTM
kqji+IZXYDVdrR4R+a1wKDcWAkg2gpRxHWMxQaZ0UIL2LaK1vTsTeyS8o29NKa0z
vj6nP92Juf6L9iySNaBElzTvzqI3Yk63yVppA1lY+tv+2DIkZXUrS3YR2JugcmK6
DBeVH17SxLHzBIpYhuJ5EzGx9IIB4vkUdSvxcL+uj2gBRQGWfW75htIpNZEhY0+a
zlWSck2i3/NHPLyOWWd2tv7c6hz393y0jbWc48aIYTX6WLGP0aklxHjCSh8AaweS
BUrW9AkSiRxCHYERGc0HVCwmhUbhEp5In4KujxwVAv73WlOxKqay98f79YGiyRr5
YuFXvWXRmVGmYjyjw8PkZWfnoLF2CD0HYRK+xb0mAaxB9TvctkjxzKM8XFDywFD3
JixAir0X39FOMvLifafn4/Gbxxk2YQ6ESoN7j4IFvT0jz1+t6gI9QvesHfK+2Nq0
dM89+8+Dp2phnwOdxNpT186Zfix4mifY+A466o/bFphPfnu30IEctFaNmyxgA7ZY
Wylv2nwpf2Un+67GElzGet5Cy507Bxmfew9eflw3sFSiPV5JQILMYHLPhYur6bff
W9qwdkSoBgUTTofGanZs0StL+lnqbrfluvUibAqnx9XrrgdNhneSdqa/Fu5p0ORz
dUUaGTJVahE0yINPdvqKBwHrqC9NWfeb5g14IiUweP19L1nsNXdeiFf+3yNiDQYE
h/5Cj5wz59TH9rtsaKPT9JagsXDaun8io+Oy18T/m0dBGn4kYI+8/4O58mHOX9YC
0GU2qNdVg1Zr7KbX/hXgmqq/j1hCQLuNextD9GhfyivwQ9Rk8TQC01noO7cN7x/b
rVCqOJPhZ6ygVQ/CuthaFdAJbD7DSXOvB3bvk+LZXvyIPq+vgodQO+x6VaD7xvNX
a3VnZ7Yogi7TQ6gtHpbvytlUiJaKZYuyT07KvNtbtYy8GtzLe1en4clkkPNV1jyo
OOhEVH9pdvpBLVp82Eiy5w+lQBN721IG+sca4LZz8HF4lNdSQijK2Ind0S+Zyinp
M10dsJs2h+j77mX/Xi1/qee/kZVsRj4UX0laTW7cmSkySUGPei8/Z7fmhCL1Eifs
IbVNfZpUc4vwniMPlRH10IcdSOgrggfAATetu5VhBqQ9jwpdyxcvqBEvGGfVz85Z
y5AGtFq28kdzv8TlJIPZiHTaJDrY2TuQ6xPCBKEtWbLItWIfFh3K8thtd2LT9n3C
kzehPnzHzAXfXjIcfiNM5W9ooQRt7H3IdtxhgpZMJ6q45MNTpiDV1E3x4xYkGlvm
73n5Te5Ev2vE/AeTYK5gK6Tv04+Lox6hjJQjNRwT5/s8GQet9aVsEXNxnRejH3+V
cFBV1MjgFM+3ceE/Xcr0AMSCmM+eSwK41TuBvKrRPaKP09vcvR6fWnshPNJxlYwN
JodTvuTJ3meXKRcT3oWCzluEWdPUcYTj1jvEZwDDAMT+v857ifREpsxhT08oqby8
az7HQxxOTAZSxdiT7p9lCWkovU2rNbKdGt2twcAxQfXcegugOVbic9D0bh1YTZlR
S8EOhA1WyDBMU37eHg8Ti7NDhqZ7khaUMoF6I3eTuIctH8PA6GzLs1HhCOIHeSFJ
uYR/J6EUC3Kcj18TLlK3W9vPMBAi6CN6UTmkUrd0bsNeAieRbcf4zgesFn6b8O09
P7fapyiqgaQJt1VRZAGQdqpMICz2skgleuZC2B2uYdnh3rdzRj2dYAHJnsmz8Lgo
WCJhMgj6J9B06CIGM3b6618qLnmLgYvtLlvU6MWuGCtuGyhuDJ6Kbh9MLyeIin7B
MEArdLgEc+UaUzDl/vk005ZIms0DTx8EY01Cz7t08TeUoOof1q8w29yN7Y2nuUBr
w3WaBhPnBxp3MG04eShjRDDRCY1X5KlBJGf5PrtYxs9X6JlsvOnU3iLIkUCG5rlr
OkAIAihxctDCu/s8WFD5xOxK7FVG4JtgwcLS69bmH98V3mEKlo7O9VK8XZqFZpqR
STtyvednUAK+y3wat/AOQtZE5/jtUfXDTlwHISZEL0aS9a3JdO++lz58I0NLT/Gu
CFAFjyVs8EMNc4AtvDoaAY4eeGusj2HOqv0spk61I+/HKwjSVSmn6SP7nk2uTlqQ
sAFU1B3k/7sa9l4MGD95av36De29F6nigxMQ/DQgm/D8NmfKPILumiEKXUBm5G5q
PteyoAbN5oP6nsJTtLFw2E/51XbT8QiA5DFeaNcvGu6L64EYFA5oU88m7o5K51i7
dWYVhmI4CIkqMYqvsydSYW4kBp5A/4TcH989JjsDMGYUNxGcWY/02YJQPKia6PzF
Wv+gTLpOAbe53atK5G1pweueVyFECFToVIbMNUsG5MkyxCONzM93wQehULynpIWd
1hg0idptFm+bpZ77+1mWjkB0YsnmF2EKYxh9X8tCwBYj910yptpFabDf6UUOI+Ez
EqjD3cFzxD5sgfmkCm7hrmvvBv0duF/Sm6osGvf4pPx4qtZN9jeyesLDviiJ1Hrb
Ia5DZeruBJCMRXrBTvLlt7/swuprQNVYPKbEo+jA3bzEuJZlFRMs2xf4+yDXxozy
XujiGb345BeKx3g8FxhldVwguyz51/QN8CWFi21AQLY7HnnL7VYGK7lHIyXZvIKw
qh2wnSawGaygj9u+wEORCCTEPR7Lm7WGW5C34X/TwO7rL6lGI/+/hYOKnryaUUUV
GtLpFsbH64K14mnf3xtmgGov8zJri0KZMKUI5IvpO3c10JjPamtwrrmeYn5+JXgk
d0QLlXFZcdBmttYGGS33tXQi5tU0j+8lYy48cNwgOwkLD5XXmCchkfWGYNXQbj8b
TdUK2qFSKvgYug5QvIERRtfw+HzOA8NqvAlctghxJc59Pymq5PtxuCfsnE4+BPcp
9PLkzHxm+FrAG7YU/02aoY//hzQyRBdZo/PIRfsYFEF2z6wY7EFlxjQEaU0m35SL
364o3g1hZEiC3ZljYMA7LOOi3k+9tRvfAmfbsRFnt5fn2OXo8FsEAAgKnVCdHUsi
HS3OovI5CWQHa2gGiIiA/EiU66RDFqGl2XFT3EeuxdEWtT5TehF7hyEjpBtDofei
OpzPp2x61UB8PZqMm6g8WCbQZWsrFx0AkHsAWOQ0L4+z9BHx2/HTTSLlyGG7rxK1
lbHclKFUMqZwRL2zidYaO1aX9gBRjMQB6RTe1Gbcw9GE3N0vjvpyHfwB9YEfZN2v
JbBnir6OiSldY2vieYJPTbOMqoRwC128RSpLKQ4rYatSq8YYSf8DwPujYhLRp8eE
u6N6Zsj0ynhjl/1dVPys2WP4YMF1l37k4wmuesoLrGbz6i4NX7jhgtuO7/zFExQb
FjqgxcMzLc3bnTB2SB00PBXL9cebbPWaIRkZ74BP8yJmPqd9VkwGTWpilNGD278x
OH2ZgrHOxKL0JGpExmtbDf1VqGCHaZgTfNNobTKn4D3VoUfGah6sp4m1/iaLKkN7
zbEuNs4h2v1rXhCY+ykdJzao6N7/+mqbUa5pGPjtJhaTNRvgsNY3pmtnAHKGE/Oq
FJQ9FWVdR+c25is64fDIz4w/NkzDA/1BC4gJRXbpeam1jpnzeE3XeAZkuhVRWGeA
i5DIgTl3W+uJ4R5kvLZEBrGnYG9eW3+5vPn5oSovocDcwujLrhESJ39y9VCvXMbe
+CwHqPxviujdqkeryEKQvLrSHXoeBAqtgUwTARrHpd6+EVxwQl0DvvqaPH3Mkx8R
cE2S6h7l76ZoWKqTekcdwpV2JaHcXTO7P7KGq/3wPoX76PI23XBsqSEUf3wtGVs4
JJevHpVrN+mRE+3kfPiBDLHGOSvTvL62261dEzlkk0PE0msXQgopg5O4CNG0hrB0
TOB4Xgsk10MG6XE8pwexTY0fr8ZjVAGvJO6uEo0E79vvIRB41wIzNZL7MvpW6aWU
m6/yEcdVp3ZeN3u8HW6i/fBvX63MH4el+ylPZQtMdc0R6tBpl5m3bhavI2n1Cwbk
alHwomHXJQG0bm48jtZwSPNFg69MFxDYRPkqo01tBbKQiZzjJWe0+lUlpL9niKha
ghqWwXIj7sO1q6uQKsw1fzD+ZEw47SW4l1KU49cf2N8Ozamt9nHtH+OuGlx+NnJ7
4WlOuab5Vj+49hkVTjG0zHBqO3EAFwmdJIUXZPJ8YQmw/j529p/I6IN1mintc1x+
qkeVnwpizj+09qjdXgeLN7dZYbpKvdE2UoOURiCivvqokVSO/lEg/MY8+eb6DSUM
rFMqK6GoNymc3cHU2HiPG/qUvJ/8D3VRH7pyYj+BNsibm4/EoCeTdfH40R076/RA
EwB6Z7yaKyqga5scwvHhtE0SEq7cr9I4ztlp7KiFhU3zXQuXKr2c0/xDwT6G/mXv
cHoS0Xhjy9bxRu3h+3GAqsvqS6GOaSdgWtuRIfKim2GruBuKsLPDuEOE+TPZ8YXH
O+XvQ/2GwmyvQgpU6aDHoKmjy0rcJGE9KwpCrkUPMqSW/t6rDkWG6siHYOHin2iF
NWLdwxUfAu43H/1qzx48XwjujA1a2KyUWisHin167dTS1aP2NWz7Spykjq1WqGyc
wrSSOfQ9i/cFfYPoJi+p1sU/GBxCcpm3zww6fI0px32Ew25/q0serXMDJVWn23zv
gsn98IY32rn+IBpJup8CPvNxrxskabKl5EHh0kvIb7//EUjoHfWxhJjeuhKagiah
QUADjIpE0fE+t2nANP8yliJLmBsq2+pqQcE+oFBLG4ujmMZC92mM/EVrgnNFjHEP
ixnIPELmUUZ3P0orS9UPCUq3NS8t9ds3Eh4pmYKB4Jz+HL9l+w8OnzZSGG/aI3a8
9qkRbNBPxrkYXxBdOy38RBKbcuuTSIuSVmF9K4taWmcdT8tXOn36WYLzP8Vvxgik
YgbPjRTBezs1jrucJMeDj/Ff5O6JhjwYFW4mXm9LYi5FnBxgleB5/6Gvv6QmBzrZ
qa3jzq2rVs/p6aXr44uw5Yl24bBsQQ5Kb2zgnu2/RzvKMYCfAUvCTeSCwMIjLpym
eJvq5VN8txDZYcWtoegcRtQMWiykCcSCaXDwoEBpOd2gRO9Ym43Okh4U60EWPl4K
vZ1Ncvd7UKAbToJwTu16Cf7cIM3dlxOUuPc4BEL96zJy0WRf8AKo/RtwYI3FNR8d
Xb1E6JjrI9DQmfQevyqOrwv8Wh+0NH3QezPibQHT1g3EbVurmIPKVe4o6wh37Ivt
71QjJK4/Lho7QwZOmAhvS4fkfis664yeCo1DoQ+06VUT4pWB+lZHsOsMAPmlmT62
2HvnUEgLG2+h6NoDaF5ilOQOfCu5Q4dqdTsDffV9hTT4Rf31X11pXv63/NHtxlE+
kSQqRjohHwRay/R7Dy/Gm9lj3HDz0U7pyifwa6my6SRNc0NPmShlRuyizj/1wjj9
En4ZMK8OvjwxfEYHfrMyVS5r5x35AuLmXBetZt2+1XgR+kL4dj5IxFH5HqLIo/jj
/jrRUxYYwTmexQGalH59IsVZYRYm6joIHUFQS60RzWlKD+KJA39zad/pfS03BxYb
SZouesR7EN91DTOIjvyVWwaOmR8KWKzmcVhMofrg6WtqCknRza7r+PtsFkF36Rb8
KhB8ZpCacXy0D/3qFTqtPTQO8B7UrLFvE29Cgrs65feIHG/2ZOzP8nqBPv5dWFKW
ArwAF0pnvO2PHvDERGFu+RXTjxfzTSoDsg9kSlvqgt9ohhKW/YSd0lx/Y6oTiZm4
GQ2hsT7wlg6LogsMhYb76eae2oKrgK24CdGa5fv7ABpJ4pGgEbVLbCMF/u4ToG+a
ExY/m1OO/R9WoCTY2ez3/npyLYGxXB9/uwjJWgK0lWOiz4UywvqUXtP6ZtBbGPws
Ge37Xw1hgF9f49JiC8UBkf+RFaAWzqwpxUezpoTwECmiIptiGX89DB/lsdBpmcjY
9pmfE4/G+dQwopa5IO2C5lueXz9mQUajlLy/tgOlbp9FKVJktZiMNiMUPGySbqbw
tdrPoRthLyi/rSDGOFVIAGBO1E+ItqXke8Ez9scOhzNC2iGsH5BD3IzuFZrYJOFV
mCyEtDl6GtOpDrI7d4uwyMjCOiGwVQkHwcmHlVtrfiFYjixSAvameIyaq5qAMs9m
HeR7jb+1aF0x1IxeynoedvJDI/4gVCH3KhhFuZBq7LKWwvAXO4zeePY1KK3boKhO
lumezUMHJU/b/IMnsQjCxdk0uqh+XoaYCZtSjCr1rREQnHM4OBack2K1oYcLPPr2
bqd+X8dncj0PvkzZ7p2ZxdAMirkRrNVBA0FteSxzf8lR2W3lCh+bsZvb3eTUfDYA
i0Vy8ofoOkurlUMMogDJQukoqxfKDV02/WV4kSly89MP7h6nuAZTEonuR7vXiPuJ
jRm4Gj2bedP6bVK1RgS/61y0l0S8F2q7ykXkY2bCQN6qWebkQ+N9hbU9zX/sIL+r
OGpx1wU/zDBGvN8c/61gUkXSL9cwQKKpSsGEjf1anSUV8/iCdYa1mPtNvehU5CSi
5IJ/UOEQuk3sCrnz4wThi9AVuZ1BpCGU4dbC7XmuVzPb2AyJQDaynlmooDGNbsW8
Od+DXf3Xi+RuJv/8C2RPJhsCay96UWbkMm6NvNTn7JrW0MRQPJ1cAsj0nKucLXjX
jDQcWe3k64V03Rc27OhryLkaSgeHsYSYacT0u8sMrOkEZz+qANZMG1wGDwy2CBXY
IhVL+VzbNCpdn2azks+vSg/INzGbaF9xKl0MBhT2eqGoVSiPqcXSONQb4rCG3Eam
8CQhS4ueZdlCxeXaR2faQBytBGVraetNbYOSfHrEHZOy1UeSwAQF+V/0H1NXUlaq
c0Afe/bIdhi8uwYQU2Jx0rTqpGWPqN7DkkR4g//yVof5bmvT5yb/c3+6YI4x9s/I
mFS3jnVLbnJyhhPD4a5n7zif8RsZIYGdso0VoYplt94pyZXJpJNBdtpLWRyk40bq
a4DIwZtm9C5E6c+JlZ6ne+Gs5aY4WcYVg3GtxAGrmGSbImc4dIIiXIBxUQwwYKvJ
cUSApVcWGvI5UwIAWQ3no0OyXvHwHAV0iBs6aYDQbv5/CPfiA+vfbJMXqOjodb66
VGToagEP+S+hmW/N0RR2+5YY16+V9T7WzfVciXj7wFhSAX3KSiPlnh/mKuwBtESO
HMYpS9euYcVeKwDurQEBkujaP2dKcIaGk3St+MJvChiWYMZruFrYRsOGcTySUstb
OQZylYUORSvC0PzpHPznJNPNpwiX78bjADudWMrZ4y8ACSbljBoUIDF7T4za6elb
zcGH4mRe6sI3rH6AXpOdfbkaZ5/TAsLp0Swnrf2Y8JpIX5xDgjfgJ+YgfelbfUAV
aQT07aC4ZP0twSmE7K/0Vqdu6YHJMO5aLkNfIy6uWGpICD0+M5ALKhI+GvYo6Elj
izknsM8VHne5G/AItCDb8TdnETSLL9ptKM55TCjyQKN/AKPpylj3whULWrWVIaGE
TwyFwy4im1XFUA73KaTrjjspEgt546+IkTL7GppORtqAW2bMw/YySdQc8sc7S0aN
Jbon/oM38K1ozviepkuJg5Nfx5LAlfOPnafl78xYNW3miOg8f3601mlAYUoMTS8j
Jz95PCbnIBh0G/lVuceGFvPWOsiUT/l/oVlNvo766szAbYeUaHA/gALgIuo1WvHs
uoMg31msfju+NTNRHrMRO6PrgVD+xXC/EcryTaz7R1Ky68cOLogQycyLadvOslgU
CnQad/d5ywD3WvIW82ioeKK1PUb1oywYmLPlnnE4cMmJDVtO1RCu02WzuLPZ6pnm
6KAtjdIfUpbSRW2Tvp0Qy4dj/bfY/kU3AAAkPmlSkLu6NOMP8X00ohynp9CcK4j1
lK+RdlkHNedU0bbUQcF7mS7T/vuyee1bY3XdQ6vYm8/4gg+50f/5ZgK/ycfIhwEr
2RXgO+fmLiRgkDYzpLcPJZkmR0AlO0z2m1UuypQwH78Juf9OT0jPogY7EFoEVEko
2ODY/ZQZzLHp5mstT/swq4iEzPmHduivjxlqyS4ZcWcInh4d06XsypRc+yQ6nnZj
3vrXBhdvc2hCGW3m+nt9t9xbb3MOuaF83Jasptv2sW2ruaX7v4n0I14Ojjb4zrUy
Rvq0akC/M1YshTsAIQJaXh4hhVy4I5++I7Y72ZnruapAqzK6dhShWjYa0EWyjS94
2efWj+u66GwtyBPhDFlLStq7yFaceOWjE3W1tVY5J7Q59ZcC3CpTAkH7i5UsEZ0o
XL9B6nmBXhnIKqlubwZThz5XyO4ZibnSAAiaoNv7uhm7IhVqofH8p5LRVugxxYpP
YtUakPnx9woFXge20yjxnGsvulItfMfvYiCkGi6V6F3wYWi1OlPBgUlZ1gPmJ2dP
GF1n4YaUoSK1RhneRp3RvqEl+gotDnVEFa9PJJkw76L/c9FZKM4pCKdkWyGd2Q+J
UKNjPVxj3CnXGmZe4pyr/ZKXOgahgEAtmqqnyoJEWuDaQGndHdtkMuX75sVMAdmh
ZucFc+ZNCN3AcMjkleq0muBti5iZy+uB7FKkR+qMIltyMCuRis+uU/pDCVS/vWzJ
O7ij1+oZ0FA4ja4wT9A2pI6j+NxcUBG8u/sIMyVtiblsFoVHpY8bmwaeYR2pj8s6
fFauFGFfyPVPrqp1dIV1ehO/eahvqIR61TPlKSslbQ/n99YGrnv5EwGxEDZTZayx
d/yLY4KAkE0t5ZsQI8TSE3RYzDanYuib+ckCjpmfumxZWZDsXROAcdi5CwQipzKK
cFAK8Jda7LXQeLH69TA1kRBd2ko57s1B88T3PbA5zSvGDHlaHU3OJnVgS3U0rBgY
1jgBwQG2ndAVOfstD7ahb2Zm5S7ymn9fuQAoQnuiCSh+vtwS7bzT+dRnDUvwgJ/R
7eFFXJ1ZxE0oqI8yKidtUw/upj4ULBiHtPA2rWWS/prnOsq4ivWA3HGU20UgUCiz
2pPMewCgUvaDuhfE7ivNfSGByjGSHMmzgY22P0YXSak0aiLrYFqN8xSsevFKITnt
Z2An/YnwfjWmZLkvkTTUr6Qc7+H31YZ++K57uIfqxwEsnRXufJsTT2ZM1YgrIouf
eNqAh7Yu6ULkkzmIT2WhLFk184fZ+L/xmENj+1JpKK76DjbjZn5oGEgkFLkLWR4R
BiKkUshrdkqOb6Bqib9EZuqHhuLNH73ZL4NI/roBFA6QNyLGqpBh0n1/sbL9Qtql
cJEF0mCk0z2+oI4NEuqr1Cxmyr3tnEmjus63Yh3W6MsPbCXITWnW8+cJNUtqTgn0
DGqc4t+uK3jX8m5Iau35q+llcWazWe/guJpvr6RsbJtrh1Ou6eUb9ya2PplmgVQn
KQMfYQu6Bn9U3DYm6PY52dby6uhpOfEYS63UjeLEFa9FzUTeSfMbqV3KTORe4uQG
wzQr4/btLUHu6PFoBZezgMwVM8KHchYYT++J5fn4MZBhTVcG2xouhs/SEoG9lgk/
DFtdy7XFlFH8M6JmSF6ZGIeT6Gb0AhCbo90zjAvCvB/wFGRaB9WnP8Uox0DHfUUQ
3teqrUvVesJ0qm7P0I3BDGFrRcRBzbQ9KlMhHjVEUy9E5me7ccWk/JXMw7IBJRop
bfDuS5BKrnUc57Dp/QBsv/n78aVo3DMctClIpsAcAFFbSSfAyrVGtbAIzC/qn/+K
T35zYtdb/Gh/0UhNGxPvcogu4yReyVt695DpuQI/bGUr6kb2SK7O+/34ab7H7VrA
WN/B7BXrIstvkxXnfuo/1Bu/GQo51OutnWl1TeEt6dC3fNQA6y2PATAn4UgpylYJ
zSvIxlfESWU1QUkQu77AATN9kvJAEFwR+lj+wbLJpgqW6UYfCs9vJaQxvK9O2T4H
sX6cdHJdc/AP6mw+AEw9n22V1+VWEQoxzEu1f6+1JFn232znc3+zHjMlKNvl5THD
NuBTRmYhsLoYiULEEz/y0IhYwLQOE76ictMKKsi1hXt+JT4WdVwR8J3y4O7B72Sk
gfTcbAWE2eNbc0LRkNrOJIbpd0+5dshH+DKPWQ25HI5N3Nvb5fqId389ViT3Nwmn
moST2/AuvDz/UQPVhE9Jwm4hXrjn9gJ54DehGjlM/amBap/DSFd0YUGZFnC1CMc1
fAGnHYj25qvNWXQa9Km1pHrQ9N6tnCRxqQx4zMPFjvjGDahC6hGTGkZ1tzfG9c9m
46ub5XDt5/04zfpPxQnS4FK4R+n+nDvIH16lpv3DulY7+S9huZs9DiCxlvZX93o8
3OxhvAfaJik2fTilZTZcvR/QThjyjCvU7kKYPuHU2A1vHBEMbq/wSVeSAXLHA7u/
L0pYwgZEG17MDsHYWVIp/5VdUzEx7FJ962L1UQq5kzZOblrytWF6kNtHmbDDYfD9
rn+KP40qoxOo/BIXl5G008Uc+lmVfEbId55zAq7S1BCP012yVe2XJHEXahD27B+P
jn17j9tW2uP7x3RLORm2uV6/QOHzDQMtTAmFRPiZBNJUzsLmQw0KWk/Ngd0HKMhR
nTwKa5OQrXvpzIaw70ZLpUSKsuGRIb2rREc/A0OhLvASizapp8GaM96CSR5cd0T0
SRpfH+Ub5uLJx5vMZp1sgENOAnvt1PIxxy6afrsux/+TH9FraflDU9DM6EKEre75
V+y/47OIrHz+8dIJwzrZUNNCHddNEM+2+WN9ICYf13Jp8nTH5vg/h2eJGUMXplBB
M8P6gyvhHIzpAMP2P6D2ZvbfuWgW0+nLQ1Yg2/9StqPLAcN+kQVE/8XMzIR5vRaG
e3w5/TPA8PaD0mTyZxM4V6ZvdSLY+c87Bdk+/ct3OuW0ksUg2Gf6T9L51dda8Lxg
wKFvoiqLjhb/vq0kBTJXQDIYZw8bat6SNf64/QehlobEevrjM1h1ve7ajyC4FxrO
vemNC9SN+sGzUIfqPsp30I+F6QMhGqk5IKrSHavx8oCWjtnbXichjss2RDpuELmV
ZJvB2d9CDqK49zVJtHnwsSHgqjN8LvYnw1PTtV3XOPSjLCt0XuWVbHq5UdlLN/Yk
SdzDy5M+9O/goO8f5XcyKKG9Tebgy2QvCaUQbBkUN9RTsi2Lqy0iWQiPFwySTUVS
jh3XFS0e605u7u4kzzqd47bR5Kc6908JWfceL3ziQupwEKkGvudiGEPtusnvMhhj
NbttdvEYUOVeZn1faEXx8u89FYDpmMcTOhQ7D70sqrhWg8YGt6BA2fkn6GKVPJbs
X5qvTjnEzqpk7tWI6dFrvhLfnnZ7nEGQc7wnY4dobO2Rtm/xL8Imo/SaVgOIf40k
yGRP0/PAkkaJq/7+OmqxoQZGN/3PyUe9vi2AzMaDwzsBARlxBO7Fa4XtsseWBV9/
c4fFWFPf+UOAqMzcA8AHiooYyOgPOwhmwmYOjzcKDkswdFw6Zi6sjaq7p+rB3Vyf
Y7QQqn7KKNfnoeWTWF9DauIkF9bwLhH8Afjo9c7eH8SBnpeDBGTLOXn1s2OTkwsf
hif/tDhVo2Y4K7ZLPMiNc33fDnuSef23ec5TNH24xJXrbKbc68cTu9J253zhQndH
9ZJ5D4BkeRvkZ9J3I7vkhGfbcC7hQl3eUmJvd+3IFl49HbjnmvuOCuduT74QI0s3
H/lYYeb2HpD3OYJMxjtrIiBh/LDO8ExldVgSGinrkbQV9vVExSQvdfqx3eq6NNkJ
fos/cC306Rl9VHoNvAsiMc3bPa1lkQnicpo1jBbUtX8y9bbwcnkiAMg98b3groVS
eCVYkksFcogML9yBBAW+BE70EypoHcVMex89DK2YGnqg+3tnl8jFag7tmCkTpTSv
Grs8TOda+lTRmo9TO0vbbibAt4FW4Y9NyqejvoJZaRsbJ8bV8T2qfNT1dMfauGUb
Ys8Qr7zVHPGGtQT5aXLGCnRsFMrsdJiKtB9dR1T78R3YJDZWl6Dz13lMNkriVoLm
BANGxblYiOkCl4mddCja8I99DBBPJyplg1RCpDMBTGXcdxXWk6JDu6ZxuvYjw/t3
88llGGgxrRac7JdqwWypnLngf8JKTg0QAfkPQEJFJCt5VqWbVkP3yY4A7J9pyh47
nZ4alCBMGHeZq8T17SPV9uxOK4q0GvX+lr4uwe4+yroOAiGjwrJFw1sDrtZqfqyU
WstDjEPNCb4093kjRw8Plk4+ULZhIv+E2ll18Fy9jChO5f7oxDOT9OcJgy+F/k/e
mq2ov0nkV3IuLnmB6Yew32ZZxae/CFV9FKH+QCetu1EnVEQpqIwK+kt5KPhR+VfY
vmFxSC6IIRwRoDgcOedUfgIUaK4CcqlOFWIkU5T209Mby+OQcwXUcwv2YAcdTJXa
d6Xx/NQzFM4eKrvuOSUbHnb7HbOXJRhFB8/jqjlR+fyUVqOAvy9lGafam42cLksM
XmOeX6uk3D0OMGoA922HFG/PYI4OQY3x8/P6I+mtAklQWix+YA3masDlS3W05z6z
ugGyYR9fGI+tdb08ObF72ETTfWnHhEJBSyl8s8ILiVrJeWWdamUuqpimzaGGKaEX
0Xxy1C/2+t8ofkP37V101P0FnB+Q5SVC+a1o1qhxlMO5LKhSWfgdW7EyIFOKfMyg
ZVyLGiiDAEdFz2ZHkYPEXqtT99TjirM5OaSMmdn16TASuUCD/p314/gp7Pu5kWVN
Ctt/UgUgZpDXnBu4OltT6N6UysYRKifQJv7+r9JWgRUZKrSnX7MJ7nhecB2I2gOv
zRjMzhYDuDFAGYgv98hNN1kqY4pkmgiNvMlztpKnRkUC3+EL/Kl5efjQKYPll1Mr
RtQLSFyzYzcIRonre/ullTzRH8XOkrWMh60aBs+QriEIJ40e6u8dBjnoOr7+OMxP
hPioPzkYkSLZoekaCrm2n4aYiithAn6ImN0Kisq5/r9+qQLkAOZa+Bs/3jf09tUK
K2a6R+3eJiYotywdObZGhTvIFmK7fWooYtWxJPxK4vyw5sT0qR+p1ao5TCc5HJ/c
ij2+3BAOqSglwwhv11i7f/dAxIPPyV3V0q02xf1m+IVUhHSz9pVfifurFOpOUdB2
aLstmPE2UO/sTigPvnp+ukhIzbon7JZ/XhMj2Y3Kd6geW7x4PA3FB7zML+VjF3zU
+wBBBPnXJSXhJupF9nkB2sxwWsEFlRYs+Y3mENR1GENYqU9sAA2r0Pe18VXvG06g
rzhmg+Ams4oS+XxWFxosCX7SPW/4fWUK7Ff2TSC4n4V5Aniu35h3Fy6rEqBbMoHe
izkOPjeeAtHfcfnySvEHP1DZuuH8+lQgytB/X36FeVMqN3/thpkTS2WQxoZ8/bQZ
HeRooqScqhIUmsVTaGvBO+LGE7JM5WVTPNEHLe19FXhgAlOyyl8Zw+9dsO+3m3/z
aMdjNTzS5kYdnD7iGjR+IPYfvHaIWvO1CZ8f1OOYqev1GNlgVKamQXKt6TVMBZIt
gnElGvJCUH8AL+fSwytr8KEhoXbwZFLubAZISXuD4vu+PubgJCxGav3pABWhyqu+
fHRNdG8x8FfuoNa4uD4v1Nubeog2iGIi07tgEoqrdpNt2Gi6uGvfXHhGzCzqiIi9
tsh5gPVOZfXHmcE59EAp2ZIkw5us2VIwjuLAMj85pCBJmYrPkuJsbuYoYEhjblSv
K+MSCV6CifZXkdk6XEfaJaMFWsW8MiS5p1j6V9cxTKLPMXH2gi+nCWKaJID4mCnJ
/asvceQn/A3DOSglVLp7BsL/PR5qaPcCFa7F+fY86c1Biu3hKgtXKai8j8+d1w9m
hZlUP3kT2QXFR4p6sXf9h9XiWn5jpRVVFNWxj7Wdxdy/4idVacA6dbdDhzw76cUt
C35Gu/2s0Pmh2pbIL6yBDOEa2pAle4Q4U6GBtqzTCKotfrIM4lvxFU2Sp7xDQVfc
gb0Qo2m/QgnvLy4nqSQajpD+gLkeRGbuuNjzWw5VWTktROWgb2fyQsa7gErOiYg+
JsTF6MgpPaQCFLkFk4irOQfnzb4kt5K2ArABGpJSArL1cMGeBxQOokqhUXTrlURR
xWeJrnGfSjmLFTqtRrMRUm+7a9V4Qr6Wl6SFPH6CsSDrV5iVwmwXjNAZ7bvXqFBe
sEKa+n3UTNsd05mWoYGWYgTYzjKrVQdcHmX1a4zra7kJi7HmC0LODblW+PBzMTQb
JeK3oGuCr8IKB6OspqdEGkmUSTVq5blvTmdbMly/MN94rPHXXxAfC+DPv/bnCJUB
qyDM7vIqMLQdxMZTfRhKb8OVw8MIooSlKqs+A+iEulfLC33p7ggJFflh5fbTs2yD
cTV4xB4kUi0r17G5W4++8FNaWMlUKrruZjVpu5XyGGAJP/GVxp7yZOPJYREYOnXz
Hs3NyKV9UzLMIjfYYRSXX6n984nz/JzOlhstOSDdmYJolKTN1AceDftHgNjgHAIW
qg8cHng2Ek4dyRUGc25bzUgqkvoUB1uTh0LC8loaBLrEFnIELYPdli9BdOb9UF3Y
aOKOqzLevf+ImaW1H+MRIGsq05M/i8ncNcRxCwpomBHeAHu2ue0jko1HyIeT9SyE
SoQ7mn8nfiLJQlCVXqhpvIXRqqkllIaVxFT+Rvk5Nz7gpL22zGSlYHJDDooCXPaf
YhDCYLmsZ9PsmYEYpszKi0yCCdCROcYz0jDBiiVOJVPgKeixZR48+h7jUMAJyy43
Jxcxl4VymReet4BvvHAi62soQG63gMV5Bd50YXLZ6xHKtzeU1UPJ7bfVKYjepSGf
IXW/wituTezFyb4DgNfNAB9V4f0qFp5hBZUpk+TE2OQIahi2VqbxfZItgWoCf61x
Gvhkmp8d2ZX6NGDr4/BeHiyYBlFxdP3Mzp0F9OdaUUHy3Sh5AZttzbz7gsUmw787
6xdcsmAm/Z0rCMGwsgkt9VUJNu9INZ9uDTgm/M45hJfcG9v7A84CLJEPOAewSEQx
zm2/aMLShYR7Q3nYrl1Mi5YvnUifgw4sgFwaufjJHsOVLSM0MH0F9hou/oQAEWhG
egDD6gct/0nA9rY+vDu9GhDW+DtP1rGE8LaW4M/tqWd9oRR9pFSFbvsIxSNdmF16
yFmD5phKpo7ws/I3w5KCKnOiPNV0RhhKDCfF+jq70f+mRC+CWOTaC/QxpRyeVCxU
ikTPpeET+YBUuD7y73EKkDNzEWI44FyhlNsEk1dEcXyll0bTz2n5n7dR0oRmZBUN
pqrJieVZdKxzPdwqKKsDpAFFLOvRcOA6SPCIlGBfYclCkOAOUR+gdk+TBw4eJ0/e
yCmEqu3x4fHrOAxUFQZVvC7s42z1Uhr/r7RgtIAf94ZJkxqgJTbFENy2ppQhAnvj
XfEyn+FoR2B2ro/ggmpfM4qQjyZLC6y4vMmah3IqUpMBwFV+Ns35TY7Q3c2GoStn
czblUHNYeVt1CvQgHddu3tDbKfQs50+2kQkTczVH1LxCJKzjFkY12ES+VRnkpG5D
AtBu1ZYOd6sL36IjBEa+gYOEdgBb5f+nlJVpTzD43r3za3sMhv0q7ZZmkLKWMwvN
I4+PEogzFMtvsBooXJrfF2wuVNzXa4ao6GfW/Ikd+BmLVw9z2UsTIGUYHTzIB27e
hrMbNcbY1fUFzhChq/NfR27ydC8Ab4Z71+NhOnIUSIRGjrYwFn5F+UkwD6ANnBe0
2q1mc0tGuM3c3tNdCLanxPk6a+oJ1Hgpxiol62vRaK4dl8UGsO2IMTJgEKZjoBk0
UU1aZUBHNjaiDp+XxKGtt7Z1wEukQXAUbSW08gdst4e4AsueDmDCsI/RtSQgfzMe
1nLRVN90yO8WVdRox15S+HeDIsdeXC/pIHZ83lln2Dbk6JU8sPzFdOlQ9uMqtZ62
MWFk1FTZJ+dlzoAUdPmBCu0jM6v3w+OCLBO6lZb2K7twYdL0kchVeq5dtJ1BQ6FZ
fJj0fUKu3rO/2QeXRXlARn0eNw6PfvlJpGEjiStBotsxd0EXSxi5f7+/S8lasouO
sUg6SOach8LA6rZMpKKpnQdGeLa6B6xkAX2fnK2y6Lv+7yPwXw0PCICrTdB2UNAr
Q6H1yD01DVisBMotlHKNbDPJ+LvAYlDQfFWx92/iUfoBQudnBN21QJATgp+gdWPA
dG+tdkqIIicF+FYKNGCxv62E4IVTQrpuEFC4LrKSk7WNk+mCkZ3MDge2ukbZA5l7
40z9d9Pb6KuAXs8CIHhaN3WKEyhAIH9qZTG1/TCLr54rcbYQNuJJ5vX1f256pIFf
1NsCcNgg8i4+McEEekqlcRIH9hjM959S4QBPO9A5Q4cbnqqW6VhHAj7xR3N2inLr
Kkc4GP+w2xouApAap1oSuzfkXmcyBl+Zr62L2noljxFccHzshmo2XDy0RbB7pxWk
AMh4gtAvDTHfu8KmOm2RM66GzFNjp616m66pSrv/T5JA1TmOSeWsLSbJZXf6c+eN
wh5dj933S2b5Qg807u1N82s2lN90fSXyqbHk0c3eMMiOb7VlJF/M+ZPwzFfChnye
zGHO6VrRV2PfgbefAt/jwCpl+7z4VDu1z3xJOIwEQf7dXnbEYMXnkpGy8TbErOIA
dtR3d/383A3H8UZ/hSFw9HEj+LFEW5mAg0i0Ri+Q4ofuJoIxwVy1IrKnK72l6B4U
NDTlpjKg6cvmrHjvUoumrxsYkFyez7WmVWdMn1R86P7Db5v+GEYRoOeKJvKyePyZ
xHmoyojzzQCQhVp3Ir3W0xEs4LGIn5FhB5YxNpg/KbB0FdowC48MdXoecliAGpg1
QiaxhPm0t2opOVDXGaFO29ZMg/AgwyngqlQoDIn9xwPaKlzO+FZoZgaXItEI9cR+
a9HOwoXu1nCZzdanXrszwbKavcSUhzRgIFHWaL50jGG6MIiJNHG28DOXn3Q+/YhZ
mV+0hFlflDJhbsO/XQzPCfIKp+mpbi9/d/p/4YDHxzN+FbHjKnx6KGx2LXIQT91k
jiMn56Az/O3MlwhGEZBgAxmlJy9mpMlB4HABMrgZ4dPUwwmZkeU6Ois2vFJKfocj
pbYrJOF6Kb79itIweQ08jXsvxC4pSWNMTrOYEnQiN920CCBmGZJ/b9n7Pfs/hv54
x3ACgp86PfuaPud9Gb/COo26TzyD+ZcIZ+RgzGMA3ugqLetfBNrZNCgz4EnJV4Vo
lZVXAGofmCLU6L5Hc5q5DcmhVHsrDEwJ4+biHU2uX1c4TpP/A7EgPw3goTgdg5++
C4Qh+B2jXcIc05r6uHcBfYuvRk42jFG1f1nBJElRcxj1/yNAM59EWWaRDsBfxfxg
S6pk7RdLiMDnifKo0fv6EG3j88uV4KuQS4404nrVe7IPjkI7Jaud87ygbhMfySEK
RufI3JrNiH0ZxkTTGF/wZ5AqPobsI0AGu58v9sBssj43AoctVf+ZAB1ak5AlICFC
mMse20kRqRy2X+jW/Z8yCfkqoNaQ1fTO+5pxNuDURru9waNRV8YEeNnYqyQZvjIA
1U9NofDJGbS/R5rSadwi1QdLawt9JSAccZasr0+cNSr4/Qx+SW9TShFQnc1NmSDy
d8A+bBTwV3PPhKc8YFQmdoZD2j86eaIJ7xmu/Z7TdmLp101V9WoOB611yC1rb2UD
l6/d2lpTD5ZjXiXUBmr75pKWfmpQO6sl4xn4qI1Vr/WKbj1JGaB0/W4VI9cc/mes
BHBPaemCQB6YBBzbGDyQn6CzTYI8+quWPZAju0/QIFlHE0YJKRjsuvBtJ4IuoBVw
mFC0Y8QiDnJvHr/1rxAdgPWI6lOvxU4yYEbKKDkmu4Tj8uUA0b03wOOcC5Xt7ezx
tPwNpFEeGdmcc51Luv2UOEfUlWH97V4KlHz1YBeOqwg2rBSlc4T9S61Hl//UYjeC
kCoXut2XVcC5FACq0ewrrlcxf1p7icymvDJqZqMCBeV2b0VDve83PHcjqwgYEanT
+DYzvDD/ty4dy4Q1mzz3pUTtE/vP0rI+KeqFiuqfmL7wj/P8+TkDb0BNcRAnhqN2
Ny+nqLAWTeGvF/2A4MTa7fz1WpHEcLJ5rWxpMp/Gt5c9DZ0LBIB8jn2tfnjQC2pw
BuvuogeTNrOtXujWahIMbJVf33CXr1aDrh5EcXxwsTCAHTJKu6JeocF9qllDY5uE
icsB/BKfGA6MGZHznPwXyuqYoIGaHLVy2qxO8neSX/Ppx0FIYsXsXzHZpcYOO6gF
21TLctcE6KqxrtTFtDzz4TUexQY0O/Sx7kizKInxMzjTNXxlL96/Qst+xZtiBWKE
/Y38CPKeTMFagjZEz+S2J9SHdK6/e2RaZQjPUheL1a5Un5go0ymLzmR1iPEmG6/V
qGUNwlzYu6EDlfyIJTmDP17iQTNj4l41rhZNcHUv/MDBksylWzOotc482etYrBse
8omizmmAMl+w6aVAZHdDqzBt1f02VVAe52tCopOogz/k/AXQXFcCYuw+ttJ61TU7
+FbdGNW2gDe0YXJ//i5I7jt2rUEat4EAub/FCRQwepsXdDFDOo2VfVD5a/vpt9Rq
eymJDg2scu5lAZaG4QRsNbAykPUwgB96WDPcxrcBDRqydxx2tXQBW6P7LBzMaTSl
UmtQXczjq49RiH6U8+LrqyDqKpLc+ZyvObWoGq02vrIyWdFoLJDziKJdIUbFsioA
ctZxiFaSgTR4hLHVa8jhQBXVqZnJByN1qLTE1vthNG3oxKDLb3KNiNLzJOBC1a+q
dioiz7OByI1PXrneEmjdlwbG+hl2kdBFWLYFToTLs/os7z2rMbVEf34aeu9/iba9
aQB1n+nvTuj2cJuO0B5ouUhxa9XqxMFsk6hOETtEZ6S+1xkNTKdBq8aZBGLTp45Z
3Bppj0N6WyjHQWOYuq2mp9s8cXX1a087zj5jG6Tjh+vZqXGS6TZrUrc1aIjSrpc2
07W6Vmpu9geCl3gD7apbDi7CPHWYg+SdLbXQpT6lfA0fdFBQVNxlibhwosqw5s8r
mpUzjeT09NWcNBDB3IaaKir8kzH83ZV82rEzh47gm3m+tMswRzDNvYVGy+nDVBGy
jn36TlsWW4TrX1ImfUKfK1fBaodANXp3voSfNEVxGG104MvKbYMp3xQ6wDXxuN3N
dHG9YnnBv/a4h+4L3RcD7FV1RK16eiKARtD03XdEGN0+b4q911WTs6M7XEKJod9a
URs+gm920C6gVNZ07Q7ptxGrMQ4z/KPXh4lQEWZ5AiAljdjFoNniK5QJ0kQbxx9r
dLNo3kFAMwtohTp1JJ9vMKB7wHT+XfZ+oJlH/DtMteKXeTFwPQENewxqsiyqH/pz
Ww4OMJSApO4lil0agvKd/Qse9gs8ttPjTZobOYyvAluPTjlwjwlV44PzjJEBnvDd
OFlq+EaNoUosNCqiMkUvsUIyuxmkuKH9+a79fugfY6uyNuVaWsNQcDa1Q/EWQPDP
Hu9ddTPI8nY3i3YDacInvzmUvRCt32YfW6285qwwlmzXs7qJtGqVuC9V/aloNn4e
XfQLUTdvd3ZBF77eKk994Qq2Cj6Ggq4PlI+cjT2oTZCxowpxC36UnsmtarHL0pga
+L7dQ18BlMdpc/SJ79SEESFZZj97cdDeiOlpZpmzJEqIejqTx94lJNmyNNQIqsjJ
XejOLrPYP05lIwy2vnVNV3/sf4KJAR5p5AIcNIHsYDM3zKwCgdQPIXXogAkE+r3j
nreZB9f+o8dbnN2H0AzoNQnw0WhjG0rf8TFCFS8Hqvc9B0zWC7MNO7F+lUzMGZ5K
0ICcNHMSMkME7jnUi88q2VQJ0+HnDrqAaxIiJz26ZUkLeqysV4NDcBnjDiTJtHIT
EETQ5Ve7ml/de0/AugsJEkDPVQiVLEmZjhevNjSb6lG1YAkhKy7x+egavhG/jUTW
9V5NQ0+6ON5x1iOuISVTpKlDeY9OzciuDNVZEGMDrA4e9ihZQO2jLSIOStPOmHnQ
fZiPYz39Jfgy2JZVmX1xwR2QIxrYJN9EWqF5OOauiDz0UU6vdxQBX5YZUHAF8CBL
nEMNUjc6QZrUppvyWawRpfL9qJlUEwBVlx2afknIVeA6WnRyP0O5+w70St6FlW0T
r0gPFm6tnW7rj1kkHCESEPz7493D5O7sUw648GXatsFc+UbK69LRo4VcVvS4qLHc
TP1BuDHrgfFs9EbmeR2Phs6YUOSwOq7jNR4AksK3Ryzd1xb17BtB062S0vjcFuxT
2i6tUIdIMX77kALUAASynCB5uolH5X4TA8PPGsVG+xfKtpl8iwa1uJMNOjEpTVW5
YiizI3pJSXCKRLBkjp1rLDgJRzBgt/A+zhyVlH/ix5FUU3ht1P3yUnhGsdz/W1bT
VUzGmTzpwD/ZvEk4+fYeGuWngbUUb5+8mZoTEueHQ/JrsvRcgSXSxviEXATpxGbF
4tdYJgekxK1212nATybI3XCaHdoPflRGx5lovcyT9g9VwvRITKAq2BgzQBzfJ9J3
JeODvMqj1lnD/TxrVJ4E4NUyu9QgqfIP+NbEYtpcxrnSfmwAb4ChiDxXrWlaRQlw
Z8Orq1C3eAM9AOKrBSHvqtDSZ2T0p+5fnOI1z2/taShdqle3ITOjW29ldrrGBOGY
pzx4CmaNSjn6qCQE0R98NTwkL1uHAzofeCGJbuyB2cCtbdsMhtrh5YZBlsJZM+US
1Bkg/ITtF0JE+z+JdeiLumSIkytlhp9VmNSdVGUziXXDrajAmpjNu9rb31GaJ9c8
klm5z76qUvcIh5hnig/IO7oz6Nv6VKIDSS0PifXXssWMCYN7LmwHUychQ2Edk03+
KAs70i8kXJK6eVWcmYf/US9ousiMQKqxF+Te5g2wU9+yRV2/0gAtx05blR6nWg4v
VNuBNttfYM2412y5AXUssNZQQuyutuNjWOLQNucX0BJSVuNIMltNbDHo6U4y7MFz
APGQxmOp1Eja9EYOj5AY/pMTEpjkGJvh7+as+BCqOtt8sEj60Jt5FIz0k/i58Q99
Hhwj9MpOApxxOXD+SFGEBGtIpooVrX56Cn5lTddKzfWglXoqSkuiqbqic02wGuop
+bWjFD1CoNVIBJFheHcMONlJcsBPG4Y6D/T7XRgWKjKf5E0YF7jgMw44Lp0i5ZqK
FAEZF+XmHCN7GsUa4+04HCD1WgOW9S5d7ZSBgGNCU+fG1trxi6pDnvfLTOWZN5ta
FS7XUa7u1Xpyb7PNA5kHeUpoyk/Xs1IDyHAY4t+BqyhII4jlEoxtFyGKvVsvtQSC
f7FrIoEX4X5tcflqajMxdvgOrQ1v5BCjTonm5nbxRFoY4VjLujO4yghPDojuvs46
jIO7+bAzOvEcQC2cR+Nvh4oxoKW3Ud3HhPQ1sKkWhR2RSUV4c8Uoo9IowGUuTtB/
71FY2VDCgL+VQ9fEJ/yvfcpnceiNHEQyvCcsPjPVhKj4X6il/gIUmC1nBGf0ZDw/
yV/2xXLzBVgtCeuWd/aps2AtuA9koonGMVvXjpPHrQksXv1scjt0viAKNvjdjMoz
uVKjwnoY0Cijd5TrXXIAc93zdT3CRbO0KySGTcel+D939LTuzmQ35ydwJEwA8rbM
MJEJ9ejAciBHuHtARnil10YU0nWVk28lNxi7GxzFJMFJedVUoGJB9qGgYiOOuoeb
P1JerJjVhPmZuQ89996PEPNaAWUS0pT68bgX1kh8p42kG6z+KNJdOpSOvVPLs/UZ
n6LOQwdznem+8DjRCQ1W1rRNX6WuXV14A+TuGSr+QI9goBbh62Oe+S63DmijaRW7
FSJCRBlIahkMyibS8+imZWLVR72lCQDAq0VPHfD603YXWLoWBzGq/Qafx4U7sKmV
ZoAF5B813O/1SIZgpMT1bqxXBMlJyMvukBD93VxRsfDBnW7NfGzPJ9dAnLzNw1ld
XBLPnANbr4UNBb7IE9PnhCZivW21cx0/SjIPPn3QQO7NozhoM9xS0oJa4guuebvb
FHoqzXZUxZf9D3Bw1z9R/Ww/NIWN6plnPIoB7tzdo5lmbTFGJfyTp2+9QaBFyNB9
wwJFoniOqjsUA67KURt+f743TzWvPWeLRDkHZD8dA80ELC6KysQtg8qUrlG8OAPG
fTuDb66UawEhDsHIzaP4GngKX49Q0wVH5U9GM18HqZnwxzXNeD1cr9u5ag03X+ZT
lTeoHKZfd8zECUi/sYWbJU57PYtaOS6IQGHchm/9RPQ1ewWQZHSdSgHTAkwGt7T3
hyypr7s4CBnmTbVWaQ12st2ThUutuIf2Gyk8wBEIos905EJyrYXCHSQ7lge+uDF5
w7l+P8nyYEZW10KM8R2O8XKUPVbcWPI2hVX0QvpZMV4e1CLBjCj2dOkZ/4lkd0aR
Ky5icsXIMowVCVU+X8kFtgGTL+pM7hPQ55FjMXSkw//jKFUp8iNqsYJXswifm+4p
njkDunDRxVT4e6JY7KABgd6ksMHki28d7kYjIKRqEzK6UqL4gvR20k3cO3vX4ZTW
2jTlYMsnOC/twIx/IVKuqFSFOlJ5VIKSmy30svMcS67SROql5xSPM79d4qH4txKm
9UTwFmfqX3NcluFg6MG9TQ9TaMd1KH3ZYlcOiKhJbxgy9c/K771PJd1r8knxWD44
BowoAIDZyqwvkCVVkG/hkiLFZek/k+RIorZvvAjzU9KKv2SE0RUBiNbvakzbkc5R
IwulODgydSiL/hiyxiilAvlZUnysuP4yQ2ZJ3e9cIfyDh3xlw1ifTypUhXpbg6E0
CfL8p68dlNysnjvIw3BYN8OkYqAfEr7kp/R5uTKIrMBPzeyIrQXyuH6L7eXK1JCB
QVgM5GTMIH3qSaxS/D0aJV5TbsHFnOig9T/igO7IIEEVbF250+wMz3Rz+FIP/5M0
4mGa/qj5cDkFOL0PaIxKNLEDboVoxer56vZHHSoNvx7UijuAvykDnulc1xtRZ/Cq
N+avjQ2nJsLcrt0wpzM9JhJwnVBr5JXyPS9QzoI7eQs=
`protect END_PROTECTED
