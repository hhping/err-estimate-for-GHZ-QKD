`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cJ8Oudm5GEcYmUEAzI+ypi70mmWwfYBVuSzrG9f3eIosJzH9LhnCsK1Vou9qgTLe
LMBpjTi464IY0AiEzMz1PiREcfxkskOFEXugRcUxIUaLuJbu4zw9U7wPgYOZ+zGe
J4gREOOC61ZsBTn1zDZKTT5vNuku69YwGOsN6qyAnBerBOrus2z/s6ofwdqPEurX
y9EoqUgr9hHjvSFD68jfHFCfZMkhIdgLvFMIJvO3MoRdpCwkqQTtMlzKjIQSl8bY
fGhK6a8P3TLznmzoWoFaBfFI3IYU2szqcDQaMRC/o2l0kynx28GSYe/d6T8Uw1es
Wqo6G08W/HaAHOEcV3noF5rQgHuHwt1bN14LtAjmOB1mEfYOuna12DdDno40RT23
6giUv8Qdb9NRUyTzrWUsYKUlHsS8wDZN/7mXWXd35i3xSOGgkhu3au7IxkZtfmb+
9oNR/TxYsPdZ3zzcB+MImy7qasMDYXzk+JLIKhk5md5t0E5Ee8tqU59wIhWX/+Ls
N88Kj9rtFT1gK0SEJ9tT8xUAogx9kQ1nlna89nl4vQvQY8z/0Xq18Xs+kBhq9BL+
GlbQm4+dPt0bf9TDK7wDgjUyQOchVVse4lp5o4LmTi7R00s1JKu4sSRfjKuJGjTm
Iujhrv3gUs7+FiRLn/zSAS70c3OKpKuEC1C9+p/44geWZL40tz4Wl2qlikj/U8Xb
zRChntstFWypx4BV+b9zW7wrt2zYz9FaN5//28z8iGwAXt+8Nh7OeOFyRQf8F71M
zudM4cqhSwIYWnc9QH9QEAtoYscOOXE6GxiDakcjkjoo8J6PZ5sX3S72JwrXj7NV
MyeKSg72qwBy5l4eusP8XLAI23fGaoZORcb+QIHGpH8dUdZnjajwkCU9AwvOXFfb
Xk0RafL46xOHqmJ4Z/MPeG0DNzdSUItafWmZQ4eus+o5ocH0MqbsGl3YaR8aPVg0
EXsNkfYVFrx2Z8PlCsnJBvktd90O8m0Kqd/wB6nwOXHaeB2JbyKYl4q1Nxwg2iJ1
cOXLqKSMMBWBv9iRX879iCj/nl3H3c0MKZvOK8CkO8s/vI48tKQTT22oTV6Qdo5f
Fdz6DkCp2MQHfcxM6nBJoDwfSHAmXTPe9+RhvA4H/WssryJ5tiqnAF6VTfZ3jNTm
santD30u+Hai8oI7d0ZhyvvzHw9gaLrmjGc0B2hKr2vSEMMWIl6YkJE1dF/GmLSy
jSkp+dF3MPdxjoLLsNcLggf0H8NZE9b1mfA98gbdXFzaVoi6Vs9sOpZOjFYi+iql
MueN69n+3ACIyQzpWhTXRqFuSxpI0m6DxLdFmJGrwK77s04r3h7VLPf6PosPVJd+
c0JOO6OpvwWV/TXgaN+1Lif6e4f3LRirttDwLFKRyfhV4F4Gfa7oXCjLhawybMpl
e0Z/yQxBvmOBvmLbhIr/dtsmAUtndO4Odm4vsvSHDzIRDxAucwBZVvrz9cQlgX9S
qhYbCOKj2aFhFaGfW1VhHB5g8ayqX2N4xtu63P4Z26gRrQHNO95yW+heqD7hh1lT
MgrIiw5G69b4M/wvn5SzsU81Z5pZhXfY1WG7e2L7LjCksTxBu9a5EWpbGK3n5ttq
HNBtFpGIm0dAoCC9IOMI6quKu+9nQu7LBennABZe39RIjM/j3+fL12EZ+ZlN+bCa
Jmqj/DuG6JqbCvgJxbSONoeP/Lg+qU9c29UVdXaCV2AkTY8nTnLvj94KpLhAJ8Vy
UkJnOlus2b0m896MRzURQ6N3t2TCSXb7AEkubqWUru9nJpZ2l81D2H42ftNDOue3
SV5pJAwaOkqUyIiLyQEqaxtyxDp45AVz3FCVODBgvF+vAF1P353wKkWkKoQHR12b
E8xH8AaeJfxiwDyNfI6lG5ustWDGA+IzfXGYjSsJZ/27Z1QQOGc5CeAWz+BoNnRP
ggy4+B1DbesLfUP1F36W2Rb+vPURUlQTAt3/0EgcxScTsCnt4fvaBUnwycAvU9iV
o2QBOoNfOgGSm8dvumKLoC0mwX10zJ3qCpx8PbgzycaXYjPnqChUhR7S0JCZSBcv
NwLrKUkwTCvR+SVijH5SkuCvOCorNR6u+qOHlHAAdd32IQ17W9EP7EoeqYd71T/C
UoRNa3j6S70+E+20HdZRxVp4sqXbTq4lGDtfJz298PdVv8qzRIkgBBexOopx2fJg
7Tit7JLyh4O/L3JjG/Nkxc/VQdss1o3IB+ymRoD8tqtmfBjHuKPDt9qANFzyLiaq
WhB45JgZ0iozxHo5pbskqzNhP5mfqqv2F/fDwXYFAlpUl1KlDF+cQLchlF9YtFen
vrWT0JeGgSUx4u1FES2GkvekX9WPCGhtyr2RiE/tLg/RRfddCocg3/EcHOZUeFHn
07WHeJShieEEmp73IP0v0aTrV7ApH1UUOTyd7VC/3OV91TPs79myZYBp+8B6Ph53
vzj/M780Sl4NhhOQVRWG8pihbMmxyBTPgOf+ZHbYSX30bcH1EB9NOZeipV64Fjp4
vUr1wqfYsVfkYYg7bFKg3g==
`protect END_PROTECTED
