`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3wcyOFJeBMVTSYJIiTWfSKHqWYbLxhpvIF3v2ABspnH6+F6xKAApcJgsJgKRfDeL
35zHuEiBvhoCZAIJWXvj3VLXXj8ZNoodQfH1gYNG9FEmrlxijrRKKeDTrSWojwU+
2dyURW2BvsGs/Hxk4HIVFGA4eWDWUq+ug25KlxZ+G2SnWPapE3nmAdptRFGZ/gYz
INLIf8qoqxusHrygidbFD8aXbBqwJgQm1Zy+ZwT7iA4DYvTuiRwT2PvtIGrKK5ji
jJ9yDiO0VMlAC+jmf7hT69up3OjYvkmbRujV9M0SEzCGLBOy39J93NlP/yleuJ6q
tVF522XL8qc6k6lNX1AlWcZefGU/u/ftJtJdHopoajxuZpYJkeE0aqH0V3J9sqJH
v4xUpZS/AW7jyL9lSwwDNLRO+no1MlBy1Ce0a3x2kh01W9kaFH8XK42dYRlHJx/2
4r+WuuMS+gybfn+SSmUVHmvB+VmYzQVzn8y4JrN5ONjoFGE3+kGU/D+LYhS/3yP8
uQ5QBVWLetzAf6fR3MyIU1VM8x75pXj43HxN+iJftkNT1g9OX5cvX5TcB+2vwbQz
rxyYDPUaOEh8OStULtrjQKVECQqC57mr4wHZS0KAkIs/M3gh+oFsl6N170g+z/kr
KZjC05vUeUPGTnDnKu6/no6qgO15tRWLaxIkuuFJGFnVIaU/h8AOYaelqmxCFIBt
CK6z26Sh0z1qmoL+stc6ASg20Bq6vRWszT8IV2495L+owcLwNCh+SeSZdto08f7e
gYs7il3GaBb2cZyCf6rbLeIGNxJMywfPo4sAx/kSjSSGHn8AMpeDq0rMlb7Iv8OS
T7di/XvVDQlAHgmfBUGH5QpDMUg/9c1r5pwYwMZn8CkNf6IwrqTqh+1S2xqXZOfa
1hjCpKioDjUNmVaXgxQYgrCbqUTb80Wis+RYvxZvRsFmYEAJ348+p7HyeWstBfTf
JNzWZ5kwXWuVjmvevFwSB+i6WcSDQXOi4vqcbhrvAnyC0S+vs44RyigeGWbI35h8
qJEj82GolOZf/V8x8uQfGL+w41eTl6uX/TKXVXa6NwCa9ckKmOTJqIN52t2Zhs/r
MkIRKHGr5C/6kOS/nlloO5//JD4fOEMLjprvJ92iBkFnbyNgdb2r0+lMTbz27RU/
w8gs8SJm7EUcFg9T74znXduYklG46Z2nZ61yBP7Ahr9HzdMzc/TFqQoMbo9OE5sC
kaDvM7Z1Q2ooocnF3oyvrM+pSYZAttS597pnEIFx//VfZP/cNiTnPCyOneMgg9yH
Qpv/NFAnXfeTMEPeypo87jHxL953YvjYR79nzzMIrNcJmMNImWc0Q+8bcM/4Dauv
NyPUE/Am7xh8vRQKy4DD/1476La09CrhJQIc2VpmiCj7W0E0j7xapvVW0ZwlImPh
Fdd0QWpF3eSbAupV3BhWbQgN1yJZQqRLKzFIZRob3mrQHP7L1AhorNrV0wFymMae
XT0NB0mphNKAtSI/NZL02LMLNlW3y1kcNCysidt4rsxCfS/P7CZHlDQ2vErr8uHn
5Rd6d/XFvLM6Xg1EoeixU2/3xwRVSgVy3Ecmy6GJqsn4Us6rxnx0If4arshnVKYw
mxkMEctI5zAUKVqwpiOUdI8hwZazuo8PAiDSvYPRZqOQZk5AkdW18qRVIseklk38
MZevEa0gPgQc/tsSD9AwbekO9lw8ZshodldwXLxk2QbKfNaLTwnDeBLpJHsyeOQ8
HE/8TMMLDGEkr7sukOaZm60Re1bflwdcSM57VNO7ykU0sWnyWB1oHlpoGfePS7Vj
chiFCgnPxXge0WPsSLDn8VbhmAczHgPV8Ev5nI6k/2hGlA2NDvnPXU6QxxRBTFpQ
O9j8VoBHUg83liFhIYwhoq1BBJWWr2ddfQ00F2MjUvobFOWI/WSVvPDbNGHxN1QA
d0pxKwFn8wxctGcz4hHGwxv7C0Gc+gqxDR6hG7eR6p0dS6Oi/91/eHOP0y+UTx0K
AERW4H4QsSOdtfNuUK93KKKkQR6CIv2X/f8SnRxJ8hTRKl3LtG4/hp6wV7Fl0Kfq
KKDqIxT2Kg13SkqXGjL2dNdrVkK/OLdeVqbWacrSXblpZbsNGvJ57j7Nj5PRBqcc
KZP0txHNwNmxM3q/PrXbImSvMCV/IwhFVh1iFKrDAAydZAirnXaPvGJwic3G7W0b
BQfGy5QgaWxG+PkQDgg97icv2jO1ZFhUtYN4g6vOYx6x2zRrcgFizJqIRUWpKk0/
nngKR/JQPC3O+fJZwXaiZLs3DQr7gHVifOSW1qI1wt+d3I/od85FIP1CIipO4AXt
3Xg2oSUFsMnkP1bManDO8KgKtjOuZfzEqkVNRO0J77xuvPk0iYn9eB0f+efL9ueu
nFee0BhaO9DBjR0G9wGFSWss1PAVs2IhB/VHDuCMAU5lBYYC/z1bcDCxjZa9LQLw
Z8+weZIO7ywxnrW+JGiNImd/n2RtphK+JZLtzBtH2rmmMmiogAUtUc//hTKB64sy
Dfb6a3meMASX7J5H0HMiilQrhfl6Soae4p1emBLwowfximDbMzEKEXYG0LFkXr/3
YfUiG4agmb7WPx9lKXiqysHA0LYFo2xrotA+lsRl3FBvF5hXlYBPwZr0nQIi1TVS
V6onlaSB1sLmjz8UQzN/ObZY2Ie/9I+mfQqxTZrm/L7FaWFwMvIr560+RlKTJbfD
IrZKpXoIS4wuSRjjWj8l8527G4BbT9GGEd66LixqPc/hYIKlLphpvWnuTIJ9X0KV
D+3ZmB+2rZP8CoZnCGPWeuKvqDMPoTYeDm98Y2WanJwBGb1Rl4i9M5qybNwoa9v+
0LBXFSn7XU1bM8tWG58Usv6ZcXSeDnrZUHH2zbjT4wB1IIfWEZ4kEVsKzyl4eKMj
6B0DVSFZ4Kfo9Zak3fyBrBekM3SJNn6RxAktpAqFzNztkIR5NPIUEwgcw1ME1cqI
7FOtTA6zwcLeVwDMoZ0V/7mVQ+bq4ftYYAOYlnUhABT1K0LVKzOm+Og/tRS0wv1W
jPt8lmQKt1JMlJD+ThxoBuJAc9kBNI3U95qjLr6LfpNhVIBPtCOapJ07ehQ1OYWp
7GCiDSnTRnB08UgQNqjOjTi7NIOG4sb56Nwxdxr2qpFaUTPod01ThhPPcdUzPCom
JeorHvso6QhEXJwNvIZBDKCnXQH8qQWSL5cYj5rC2XA=
`protect END_PROTECTED
