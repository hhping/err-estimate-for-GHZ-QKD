`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sU8sJxsGY4WnSXo4L4FMmFbsnbtRI2B7J2slDWiAwTWGJbXedXP2UQ5a339Uzh86
puG/oeiYIPNx16915ZSebgc3c0r/Ag/cYa+2xfyU29m46ymDqfz8gwVieJEU1htc
HheshdYfcUA+A+YfRvqsdEHoGRMZPKwZCBpZrstbp+HuB61Ck/9Htll2ejRNZiEK
DNJiuNARF7ZRm8lIrCqqllt7dKaywiOeGhZ7tAIAg9PQtuyJviMcc76SztHpZmPC
HLGVwSxSx8L/MlX2j3OnKlZZH4zSNAUNx0GojOOLv1BbEohJpjKyeE33R2B9DCmF
39g4T11VHRsG7glLraNF+fpsnem1K6yGEcm1lb/fqXJf1NNxwU3xUILlFlJvHvUS
TGuNAmZTcRz8ULYIKeWpZzvOEwCcc1EJ+Se4XE1Q98xy0P40tJhXPKOs0kILB2vQ
q/XbE/sgukgVrQmNx1h6v78B64H9RPX5fQiferzE/sywlZiUdCqkpWjzHYBKfuP9
`protect END_PROTECTED
