`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZXvF52kG4Tblg1fA2oICC5pE0PS3RoPSJbQAzdXcvbbHEYdKUHt+xvRFtTYZ+3xs
4Uo8nOk0Incfb1XaimBDNh6N3ZOPuhgMIsitMwGHcJ3LmnnRzylNeSCePOGYLFTy
7W6eNFo+0FIYYq5eJApzv9MSLG98GzA0kjkd+X8XXGsMfTmzItkDIaGvthy70kbl
1mxsYzcDCJRA3LYIU/lqUlixzQ0FaaV4QP+VI36ZeLdz56IR+2DQh2VT9ED7ghuL
aw8I2AI24pmzkvTiUFwmJ1zmK8+DN3mvweh4WTYQvuJBFn4INnn862abICmOqEr0
+uyX/lfd3LesQMOX2NRlmmhp78zXzzyd4FePhM2NAG1mVhE4HyaeGrDYjmp2Jmrp
kD7plfwKI963K7uZu/SiHX9Bg3rJ7w+0wXsRrB4NVXvPoJq8DTnaQAJCCdWn7LGc
jahmlqtMwhpMLOjzQOcHrlbTdoUrMtBsto9qerbH+ChsTljRsAF9F3sdOZr7zWfr
GBJeftOxyNLFZx7Xt5bbVWM34RW1daentLpUy1SIzvfekWbCvggJKflNhxPE4NFk
HeoNY4t6s9ckKtZ6zbla6N9X/JJcG+A0b7HamQ2kn14oBlt2EpTzN7uj/TON01cW
I97L2HgvccBkgZuqD5Ys5n/eqm04gWy6kLBZGSFUkrkpHcr2Qqq8En8pX9bnRcyj
CZ3sbZDYpmOdobcCPWoWRM/4We8AW0NOgW0hqgAhwYA4WCZMtjB6rDtHzEt4T/HF
z/zeuzelvEtnIt/hBJ7Nkb92oiJoUHJ8Pk6vGiuGEbXksEdsE7Hs/UckXCjdm4er
LjMrGpo9hMu7QjfTJ+hRfYNzudfiNa4MdVX4YOlqDs4+7qRO7hOS7K95PHBgJRur
ct53YMB0FUd/IJIRF6izuX0oPbW6qAggFSrBuXqQ/PCswJS3uX8QeUPFykyX5r0i
FiHX73jyh5KJA+FIvSsApIxZU+54saQUYdIIale4BWcXk2/Uf7F8MYmCuxxJGosR
4i3D+TQOUQFSESBz57+ZizMA9F6uhKJn+upEirT8gqGYDpQpdsF8QuGOaBLTnzNc
p/PVcVu7Wa40/jDAmyElZIzWZbsFiz+8o3v27Z6g30AAbzKeC+n04jfZQRG5Nd89
5T917gDOiFQVpfxU19i3jo9MrEVWPUgkXy1ttU9116M=
`protect END_PROTECTED
