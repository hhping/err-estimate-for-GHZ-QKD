`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ulZY4belswCfwNb7hHp4C85ffwxRrZFysewml8HY6BrLbiYzeryvOyZYSk1/Lohu
5sz+tVY1FBgFPr1yq9cavjjw2Qq8C/qIJ1HfWMUhkKriuWt8pPKI9v3z0ubikPIa
j1G+EigCyBEr+taUIRVGRVWT2x0D575ijGkatywvsDA3r1vqL64yMcMhpSSPM9lW
+6Ysp2hFKWbd8vdXPpHUpnrCporg04YFUHDWYvaCpZBliEItIM+F4jz1C7loqDoA
jBoVIUCUV1hr8MCPoJXQqef21Xq0C5q3DkNmKQ4mKKHh7mazo0ru9FgNAVoMvvQs
HNsw6brKLh8S+ygHJ53BuXlrEX/yAkJPqt4+Y0S9e5E/LRArEGeInaILYa7AR/gh
rg0/lvTF7kAHm6p5L/Nl1X3JlHS6Yko032u458GjBL0DMWVYiKThJ3KAxMSpTYhE
nbt8Lhkss7u4QZ9fCYwJNrfpgl11IcVMqiVw25ZaSIh+YZG4GmJbru+wiam73Aiz
WmzmYEL2fzLHPyh+m0P5woUlgUoYdxb9aAoRT7n1h1SHBvMgkyvyN6kwN/7BHi1h
cFGxeKLvDo30S45UHqK6Wno+wiimztnpvJXlZ+ulzUhBScooPWwgZR0Lx5r4mHux
2PVY1P6spJjrBY47Bphi9JmRejCvQSFYeVF+96Kf52KIC/vv+9wIAZn4mKt9W4MO
mUAuSJIBGrL+5yEW6xWGOoyCx7OvKk1xIoSqTDJJEJqDu88PgWIiwWwDIxgu+5xf
NI4jzX/JXbTIWoFkdrRL3OqbX7j1XcVyBgJi4yQsCQn7/edy0v3RcZ1GwcEQeCiJ
`protect END_PROTECTED
