`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XycvhSnGY0pblN+zFbfTlhLp553DDlkFNYyOUHwS1/gEE+dvbNa8PmEGB3W3oRfN
QpD6oIL+VRuWLOIgzxfp/D99jYryvDNXaGC7hXfT10mBvREabos0X/XqugsfbUVU
A7hgNi70jNtQRq/JZDjMjIuO3uMZCvBN0nh6ARrn1le1/8GfCQtmSvztEsUyhwai
VkmygAHR+Vu3MLkS0OY+xwO+PXuOLUu2144i7AiPsCaRjQVuH+BerdomxH8j4ewz
wjVxpIKlmYf04RaAuIlCDceoaF6OJPVoR5xJEvU/kdAJg4z/07QQw0KKOp1aNLhK
awHmmgBTdTiHkqxCEjYsJ681a/h/6/Lz2zmChYqncMrQWlwjlOxA38b9vIoF4mdn
DJIyyHsx0oEeww9CscCC/lLrrIz5yEdUih3Is56DJMR9VNeThqDPVZS8bsNeE7CY
YIUOJ2QcBVnFdbCfTmhEVF+1xa9+8Bvt6zvbSgVXWBipljQFU3vZAlY8M/IfLYV9
xK2LHqwbUuE/ZxEAQUS4PLXvCW3B7YgyvXmklbmkgdNCHnk0fgoyJuWvzxvjsnso
oQ1umfpFtQStgK/2Ib/Q1Fc3YSEufJklgu0exR35y+nZL3lgc6bw1cyjHxwHdZo/
UuVAVRxjzlh9NCoj9qFyWtRWN+whu7DW+Z/pzQeIMepOVQavIU8+BU+kYThTDvui
2czIJKg0RIdEECeI8wCRzeK2LCAIzJD+m6qZIO9bnxBKU1ti8qtESdZ0xa1IRxiw
aZrQZF1nR0GFpK5sLlEge4DsNTxELWmeGuTNkzpArANXib9MsM2zR5eqjXGZlGKS
y2mJrDxi/3pGhRXUz9HS5aTZsC4mqB7/Ym/ZuO0EdZGJ6wmhkb9ErUsrt5B2w4P9
ceorV8C9X1DkMDkuYIwKN+D1ubD2PhpxpkoT46uxo8573LP+VLm7XP22qiKj4uMA
KDc8iYZE/E0ug9n3lWqLufB0IFvPQHw0MIoiwGk5e/YVWM1Vc22os8kZuCjSq2OR
+lhoiCuQI/Ze3HyRzQjT0o+g24witIVY4RaSKXvfHyGeEcrrFyusGBSpo3qyjmzH
bGnsSdRCnJMQfFYdQObbtsVE43PIJum3JMCX4wuYAFs9x7mTRsAe1lPAIOt2qB2k
xmbZNlTpMe6EKgw6/t1WvyzA6IPQItXJpOnopYd4GckbikgXI0LfwT//4GG9PwM2
2YfYVILrZRwneskWQfUw4k1VkzXRkrEVGGc/W218ceQLx8jVDBfhH3wmpcTY1co1
uqMHUVOhT1YDCxFgas0/E7v3Dg8wXZrEO+iktJzaMSRV8h2jUiedfkCfpq4iSTS8
tdHRtXidjsFRNj/4sFd3C/YK7hnsi7DKdwFKm3vaSFoOL+rGzlWKYgYG0vV3n7oN
okEu58aNEpbibAQLuQnU2YeCPHGGSogNx2skrBcndjRHdh4zy6DCPTd4ZmM2l8mE
EywpLvthcbuZDNWZ0qgp7K2IfXAyjMejAU4SrygEZhmK2e2OO7mUyzN88N8yllxu
n6JcjM97y91eAx1leeGS253bN+ewtLtt6ihBHh7Sf2Lc4J2IX0qK7Y5y6vYaSBZ5
hQGkzx04Sfp2EATGdlWi1K02MsR84t5HsoE8hXMdTVGlSP5Ek/WllNvoYE6bN8Sf
VtsbnLm0fR3GNek32nwFMEzzZ79JspSUfeaMYQ179MDzBAWrFxLclYMleIYZuOp3
NtNJDGrWWCfWQtaWNYZaxiTTMkXQWT4V7Z+PwLAYmZgp7ARE4noL0tWHYMzlGX0Z
hq0TkjXwKYlN5rawR8RzO2Cn7p8XQZlFzxntVbayv26njD1zpH4tLn5NAdvLR4Ba
0H4Ggb3QJRIFgOdmWMlKkBtIq5OyCJ0emVKJ4wRnGM6yGORk6u0JrkGvNxOSVfBO
rcxEb83cpoL3ERwn73eILy8dULRu5l7CAzpXRI68hLyEtaFPaK+9KhOAz2ZJ1OjB
Wvw+OeQPohwFHUB5EerfXcIgZqNHzqPs71xFjIjnyEOCGMf7KWFr62hkmmW2H977
Y8dybC30qg3eDvcYDDWqMRIp3w3dkME04ZLfNBO6jds=
`protect END_PROTECTED
