`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l5Rle3Uq6WPHsQHFIskYVo1scafze3TfVk+BnRnNQCmLvGTncQYSBDQUhPdEeI7e
PYLiMQZQImZCk6MLZZ1HgA6K2xK0aKx2eiFGCgrzFC2aIfoHSayLU8Nbm+FvbqW7
SOgECnTg5AqEhplCe5SBVwUn8XWhZxvruNEFQaCvEGPyW612QFUF9elLKCmg83Da
YJMtLM6i/xObcSFgcjRSkiuM2MnAmCuBjooyozhei3zdEVVTJ0H7cndZfZQJGSIQ
7ShLTWouXDPQweuzuYpf8gx9DIcfjUVPJg9ThAGwYkm3WVP1IZDPDGuObT1Eo0wz
fKt9NXguzxJl7eT6M3Qx1ma+a0y4ngmxAhucsA82KwUtsRSpZwJrFCU62HeWLvKf
GJQRsqwiazRhUMDpe8cU8daM3oucx4nzaGp8FXn8uFexI5nvxYxdY2fWdE2eQTkC
gWFDighpWtGURDk3N3JTrFMljxdQiYI2uuX6H7AMZKBw2Mmv6qT91KwjRiqEyXeu
ofIkG3QpdUIeNDDrZzFxo5ctir+vr6ffZqtxU2xtWWNbEAd+oeb4BQObYdLohSCI
W/GLXQjR9uNOWu+bI/OVE90yvmp1GZu8GmxFSAMlZAjVPqBFexlqwhBbBwzdKyIR
7stpOJK1/7HhiHeynxMZm2wFp+WOMLW6hPYOqEWesTzQrX6DQZbEkYeprxWFh+HL
0AgRtY+TY3/Yx6gwgeZLNamKthtNjgbfEe+uxU6XKhRUnSu/YjrRnWxil3dxh8zb
T0qeAXeNcCHrSMT3qYytIQnjHMZSl4a2Y+RRIkEeCLiVbIXTUjl6cpQXfvTo/5TI
ppl4P1hz3+sy91Csm8elg6VEyzK2CDl3odQT4wouyaw8GrhA8e5SZYbH25NQ4a6O
OODxVr2vCRcJRNAMEh6XKwNNC7RPsKOCP1cbH3Rq6S22bR6PtL1kG5rS6Ob4Cct3
bWSSs1sEce/o66ay3c+OZvRHHiYIcczl2E46cmNnRGgfILWczeOOvbfDR9oWXwkb
ncHdkRh/hcTciS4Pz+dBmmqrZr9nQPM4dT12oZlMLAQcusFyBK9JRwretvgtHrNF
UVFKSHC/VpQ3sgeq0yYbDAFkNjVFvBQheBfRrQtj65jmqwG0dwXOAKIXwHvAtj7e
fuptrTt+2QxvyBIUhpDtVlhKemqHqQyLFmEnNV0xs1Qo/e35e7HcRhJe07eA42g8
M4LRSZn6YKplRq6qjg9R4OJjmzGkgJFbJ2QmogdKBcJP/y9m9DA/Ej4H5YmXPTUj
jFkd2e6TwmIfxM8llxXke0ujK/FNi161tGiszGlbAtNDTMrNjoq+h/gCqOsWLISj
mJAmOkGKuVfm4NMvR8XnXUTrWwUTvSa9kesRqvU9gWG6/zC6eE1HxtLeYSypl56q
yPFo7KXZxHtrizdmmLu4R855MV1f6KUfWVnuBCPfwIjeymbYdEidRxDJW2HYIqFS
dHcs4IY8UDrZUifupIcB0Ofz3vnFHAixxZKnfm3le6WUMaw+Boa6YDsOgm3tIjuv
ZNLRAAE3UQcG3O6SnUHzJNiDhleMYcyiQGF9haF/vMzhC/O759aCbVSBjIUbeEFJ
6IAI9sHOzra9S3Q+vRnp7vnp5kxt5V35Pk3WYh45WpV8gPXVd8YIvrrgUDgTCAGe
kZ0QC+x0Sn122zd/GAMqcgnQx7iS+kb/MzG8SvLf4JNwdKUDmZq+W9R3xSSj7nbd
NxzB2LrAryPl7B+Gz960BqSMNKwayqKiDI3jIA1pTta6AHvxdKK6pQ93NL62vbgU
SdIkb46KWpUax5NfjoxExtShNKKzrlzGlAV9mX4eXF3NNKlLmUcKhuFcdameC1VF
8bfeIGImBCV63nVqbmiw//YcFy+2iziaCHDgRfc/bg/CMpKwLjalnMVmmuHECNU2
u7jEafc/eSxN6pSxFn0hHJ6FJKrjCxnIHBSuWqVB7wp2Vubl/UoqZAQ5uVthLzAg
sqYiXZKSspmsjvuLIVg3D6aBYNw7WXuwL9wvh79HXPTwGdruZ47R8evS92ZA4j1w
zLTgZKMaCI2qphgvXOrmD/S81Is8ifzCmf4+14+N8lfaiFSm/2WmFOxuQDzI+Gs7
0e1cpBhXqJ/lM3iXJTuqYUT59WmHfcpZ9AtNrHH/UvLCNredFzt/WgfG7G+TgncN
qGfQmD8+f3VrRzMlX4S7T9XO3o7FSBHev3iMPCdSjKBEycjYs3fhuxl/B61edDhG
6Qv+crtga2MI+WbHL1iLHL1hNxpPiVWtsUMC1xhQsxdvZXMx8NCm9nEzHNCnCE0Y
g5HNhU+wFVxIawAUSd6+uBSXIonntytWvAif6Zc70A0ziN3Q9YVLe1VmfGrurI55
wB4+cQoKLwZDlsBVi6YUXimurXJxCbHRGyMZjnbjm+pm1LUqUjyxgOjnXJRoNAuQ
yuVn6lGcZCpYHhGqShYjgZrWB7yX543EaMdRPRFDH2/Pu102LtArXFEzypz1jPRQ
6qT+bAPtaaYF3qxZ1vNRNBbzgEjOCgSr5C3AGXy9zqVQKb6SqzqE+msfn8RRJxHA
Bqt5DiNmot/03KGrwTQ0snGxAgxVkkaiVoARIdmytAxru+Pb6UQ2q8H8AGm7LosL
JtpLvFrFIO/Z3fwy7KTLaD9/MQItlO0HX+J7kI5tV8bhqfTbQa+m6l87tjxomi8C
hPOXq6yf3AkH1hN/2nhhr0km+/eWF2X+MjNE9V51h+gDvBrFKmTo0b4ovpGfoKMB
HrQWkaPl1mGISZhTjKGRbEUlfZ2UFwXL9KaBcAG/DB4s7mT5J/OoceEouNCXuAgk
aQN4aTwP7o7dNxrWX1dOOMAnXbmRNb/NrsLHPs0QXGervTO9MicBZh/m+VTy3iIQ
e4IHHsayMHfOMJ7n44LxStDvAywV6UyfHAjmdhO3CutahM6bcZWWhA2iZ/WnU7LM
gaH7PBEfHt/Jjv8VgW4CkRKXhVxGe5RnpIxQTOlDF0plsfdmxxRxVI8iQfobI7NL
ILZVbDLt7qje5H3yVVWGByR47YmsIJl/Irom+m71Ccr/9Ac0isO2CcqtkoZMLNly
mZGS0F2ybsjBdqQaJitd4lG1kWPXgwMgEI/IBJvOJPm1qNziQRA/CRb7ixSxFqus
xLW/O6KL0iG83z1mZS0F28bbvZvMAT8fJ1yIMJFFcOIEAIVMMpYF8w5T373PufPS
3dnz+3aFRiawwuAXlNffMFv3/pj7d/YbLlE7raZcAF57K03tkYL0TbfPFwGkQst5
bN75omfOPbkdz9KJ9SaW5Ws4K3AIQjiF7HZbI3w44gdoZBqr7T/JwajHVl8AhEIw
Z6F5wE1WneR8AjegeWksnBwM9K/9jKKqRrs2eE3U9qhfl6XRyFK41I6yQPJRALm2
6HPsGOYup8RVv2hhxRC5Ddndo+CvzxiujI3nTn/vAXt4ScIuXT8n45TPYfOb6WNO
H04cTVhtiQhqKxE+dQ9JOVirUnq2mTem2gHitv62ttQJjjynduNuF728Rb4fglgw
1l+Eff7c/BZZVnPB+OOV5NIGNvpUKcBaYczIvsqgbXZwju15ecCVV5Q5J1bndxaE
cf7cqmQfJLJaI2tZ/WprzuDAlfsA+7l6jre5s4JyfgQL13pYXtMNE6URZ/VvyOvc
SAn34NOciytEbD7AlvGyUpz+TOyZm5Sjnca6h3E9lZxRC7oGNW3gd+yeSBVSAsm4
WCQHPjV7dk/THnItnEFqJmR8Q9Kxkq2hEyMCMIzE5hDcDAMkvhqPhAF41GpTFNdx
/vE14+dqij1/k+xyM3cy9K/QCLOQvioSBTu3ttZOs2O2icxw1HVDClllZUVkYtia
n0ZAjcmRrdQ3m24NohcXkOcLmoE5BmAT8TnbNN6qB8w7+LTGvKUqMZS9Z5t0kLjp
52rZYGlJJcCPhsaYq2LAIdcv1xAbEZwYxDS4k1If2iPmPn2tnvXA7WBmRKfuZOr5
lxENQz8LJuMsxNMOprrBXYcovLtIaUGI/TffAeGI2StKAJJWgcUrhn4Me5gZYEmM
GXytY44hUjpqUVfxhB84mHlgUeUGcQmLoywzx+YImiBlZbNnihYDfuDsLxLdz8P1
gE0il5O9+36hg/Ibuq9Bd8WXZ8p0SJEep5oWljPdBZOLPEK/LsFudNhYIakF+a0R
W0QPeCFxIJPDkGcGuey4SWMRKNCrQIlia3Cw7EfffxqsSj56ShQvhSH8QEYZVcTJ
ilfURPG43+uOhnKJMkrWjMim5uZioZkGxqLZ/JomNYhXpr/MNDHreDdVXtwfHfUq
8yxfi8kObGfs47fnlBDYtOUTDmDUc04ZZBZHhPSpZHo5QD6U+NGHr4Pi7D4w7HXM
7/fIUDKPd0RymCWoAYdHmQ==
`protect END_PROTECTED
