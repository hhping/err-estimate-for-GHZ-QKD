`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M7CtMhn9bnBcyRLlX+g+V3ITMp90hSNW1YO//x15ioCKW6KbNMaVrlv/3exnZ4Ro
3MtrJsgKktSyDQfDuFPHNjCmDzRt5S+YQ4hDuj+Ir/j3Ap0Pc6jJJhqjhbcwIdPL
L7Ai/ZsHQIz4apXSc/duHOt6VknNfU5iHBo1IMM2P5B2FS9v9+SAgNnZQfYsv9i1
Hec3bGAz75bVH1OHxzo6cJCkENkXIRqDtIHYYZii4FZbx/6XC+CAUMnPnpDhMVFT
ksmkWn3+Vmzz7XQE/nD8OYAhAXCtQ6MvodW4DQGxvqKbk0n4fM+Rh0duAXFAeMbl
AIKSgr32Ai+4rNfzx5c+GKF/8DviyKLNYIKeDMtK+7eTt0AjWAgDTolb741IMVTy
Qa88w8by8CzljFfjiI2g+jhV0H59DkChDA5aqhpXlhEi6T4iZUrG/Cwh3/iaDor3
mdiR/1bD+j/jVccLv98EPizIYQpxgINpDfL6VNBS06AolhezNVpbdtt4Kdmdg/qp
hjG/4fKdrWNNxFVZOjnoEWmFLoBuwsJbeEYfmqPl0VpjweDhDFVSFd3GZFCoPY/N
QBDsJZ5XdhGanQpqN4l4HTZgYByKQnQDOSMAtzjWZdqBICrZMiFnOgBY1j4C+WQN
1yQlE3znus7shRZfK24R7tNixVRMtakFy/+rCLq7nQ5y1Hjyih68OtLvMgTkTBCe
xOKdV2NJCxk9KTzpWjiHOHz0P/Ztz/HiucpOc11IWp0=
`protect END_PROTECTED
