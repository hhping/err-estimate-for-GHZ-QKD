`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HOFjTN8eGFkR2/snoNX7dyioLtXFjw0hZeMGr3NjwlrArp8XW8zMXdEBgC/0Nnnp
q86l/ezxT3vphlUAEymDIMPeIChTGupPTOcGlIkfMfMxHFQYwIPjEfnkTw/xx67X
az3OxEY9qyGM7VyuxY5sY62JIHqfT6FQyGNg3Twhy0A8hFg33NYmh4VKz0srapJo
CrTNaHP0I2KjdoMP2xuNm+sk/sOLeFwHXQq662KSNASLHVQZJUtFc4pHdFKmt8Sw
cyETtFVlKNlnu8db9WMO2pbHh+aaTXPq5brl9yFCS9RGxAU2XEuGAY5W7rvWsP1z
N1dRmi919Sjk3hOkdyDgrLla2QzX2jXJFheUCUgpH5jRNSXRPlIBg1OhPm4o7peT
qntWj8cR/HwO6Sk4n8EY5uvIjLaJSjPGdY8S7GfvBVyaT7C24Jt9lXayau0CQ3hn
l0TLNRcWliUt4pSUFZ9SxtALZcfLByWOe5SVNLCEKDSPEXV0/WG2XTySgnYc8SqG
`protect END_PROTECTED
