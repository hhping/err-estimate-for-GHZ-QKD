`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jIH+xRzqyj+So/onIUHscsPXpR+CVU5tybuIXoio8KJ7MbaABsohs5xZ8jFdkSlt
NHLg5F1/+qKFkEqSAkGd1Lnf2VazgnvGWW4EbMU+WNOwzxWmxJcE9mhPNLa7de3Q
a2tmngi+boxylLZF/x7pmCYZ6E5FRq4CJ6TTkx+BCtSRQN8Gaf1OOBUps8h2V/9V
rYgvGq1UmI9cfy+V2vYnZOwRnYvL3jI64ME5xWL3ZtUITNepOGsiQksiOXyhs69J
hIlYkoGbj1uYWyKG6dHVAhItqkGFNx5Qmflz3oWzeubbdv8L9REZxBazmd5vkpbB
l2tLZfhVDyTAZI4HUiECPtA0bW+hMgc2041+zknPE6GZl9sqn6SbPBrjN7LNFNUK
gVK2MVSu618LRB8b1IsBwtg6R//GcwFTn0cRW+6aatZl/r2MyhW42FhPmj8YZ4cZ
CZoKf/CBFU/aAdMX8euBGdNgbwnA9Cz2LUt6oqgpbFNL7xuuTReJGjecFreDnSvi
8wuV9Dk7jmjppEJT5wWES24AarugHGgjPS4Go+o8LZJ2Dw22dbaGP2h5gPcqBDZe
GxqBdnE7FHFI7a1cYEHFGr+ILKabk8xwrIFsngN7u+eLdJWrhP8qCnLFg1aSbljf
tC9adU7Aud91c/YLnJgfpSFStXzz1VxefpxetWEcs5+ZwZwEtwoOzZAdIvqEBazJ
lS4xS4yDzO5M8a7raWTTH6NWrFZqzNZvD76ruAdi/1Zo6zZtdcTGfxkRGuUAAV7f
t/uMEVOeHvJ6s5gsls5uY4en/F0CCiFXMMh+h6Mj9ASTqSLYZT8xCL4ww+rx5bK5
mfq5wXplJiZMo/s0jQGEyo7AJvvtMAbidWCOFoGmseMzDxlfz1lc9OegWLQnRG49
Fu0tzRPYEt8FspNqmuCN0Q0Fp/qLtrpk3YKyfh6NfGwxAAi1Fqi1GZa/cSpYEFBX
KDs3mB0Iat47qpq8jqlLKNHTe0vQzaXLnkuegMgW5UeWdSBgtjiKgQ9EJUPk9pmG
BYugeswdlWBgfiSU6rFZGcuvp5/CHypwL9qQJZc7mF22hKfmCUuOnfEc44/qtgKn
OZ/BDwnkkXY3W44mmDuONG0P5tmEuudLISnQdqqmDzSSSdQIB+kTa7mFgAyjJ+zc
9RcEvFDeh6mnAhmW4eVjOsG+zFfXJqzMwTNpk7EsU1jh9i0Z3LlXQJLMETGcx9KD
Kj3LwnngG5D9eyJMT8WYuJzBOwcexLvhotObIOLNAg+2b5IUKYWiT4LKstUsfhV/
j3OYH/tgRk+3j1nb3YY98IzNfrHqctr9PELYroLPfX2qf9h4tYlJcjQoLJQyNpOH
n3IUZyEvAMeFEmwWPYOACgL8Pw4+guvQlJR3LqEjZ8Pvk2k/bgnDqZL/HhEuCo/u
OvsRatKetwzdo2tDJaCCJYWj1NYZP46p3nyxTBuxoxj8PmV3vcWQ2kGkWNXUD18p
E4erWDS8K8LAZCugGctNeUYpzU1mI8Q9mFDZpvh4q3dPZwp5JOSnUwjuE/0Jg4wW
5/P/uXY/27xfCT2/QQWwRbnxHIGVM3sfPPP0v8jrhz8X2Vnb2mnrwMBv3Nw2gskY
BUL+RPNY1N+A8fu6v+P4OOwSWaG+Jj9WaC7A+/7Lf1Oishu76IQcqBztkZirN+Ff
claeB42RXAka/obq+MFzkRFjoiLy/MtcFnbzgtiZHpwNztocSpGuI+i3mhEOjvle
qKcfQHNO2MEMOtWZpO5ff3dMJqs2tmSY6udtBwe2glBrOcjFfGqfxRx9MNrSzUbf
9zGp4QA+DBfHmHEh1Dlbb9M+iveA9KLJ9dsUPkatUZ2L51XPQ5hCuM51YSmZ/iiy
CakavFiUqwe5ak36Fg03kikeo26iXjKyi+jvQR8XR+w2LSirD/tX/H5k+6rvCpoM
gu5FvqZWoCOH9ukwozsjxYPt4I73wKoVotGVRXy6nYx941sSc4NeeE8EQhH/l9PK
WyGZud8j9rnjkIgHt35us+Sa4x2u3InUnh8vCX/4wHyeIsTIG5N1O8yYrcs0GUFw
2J6IV2/AC89LcYWhwwQPZ+BG1psWDvvr/pY5Lud5vNmr7esE1jk+15Oevf6LCaFZ
P7vVFcS5XaWK+Ds9ELsG0H41759wsSnrfFTkxVM6Ock9UJnT6KASvOOoidADydlk
0FKzTt6suYvSbPa3N5UoA/Wg/pYn9pbQl4b68VA45mI4QKKK7OIzZx/9hwkyDOG4
zSiEYPQrh9gTKxatf88ymcsrKdZNo7yBLc+0hJJ4fhG6egyVMMp5NSxxhK6eSUeE
vz0ZbAOFhkbpk9reNAPVcLMpt6CxLPOREoWqZ7tkgFb9oROCqIu6Gj/a8lBJu8QQ
teR3eD55S2pSCWs9E+4trAAE6hsPkw5UbkiUx+AhChI7g6SzcJKeJ5RkkcgW0UeF
mlfrjTo2hbO6CTDFuRqUFgFmGqdyDvY2+gzP6MM7nGcIOu3Xcwk1cttDr8ajTjX0
AotR9wclpN0rOjcHYRAl17HxEoOIcGBfPLLIZNeQVlo29ZjubUVa6HxmFXkgfbxL
0GVFmR9dSmve/HM1x1pEqYD4/VcyiYfl7NjBqLCUVfGEjBCdOkodfs7niwPslJ87
xMoNeYHjJnzryrTmIEYjYl1kpPfH6o5tyyDF8s4RG9ppTYMxmIkMWG3/9xu4E+Il
PBAQnuQOVkfpPFmFLildY+dhqH+ZhGmY0Kcb9JEfRn1xs2FKLkQsDh6uU1N1zRim
q3BPKq+ZeGCS+4zKbPslsaLDhTMhdLPW/fm/3gKFxHJ5Z9t/iZi25vFlX95kbmd9
0QaRlR/bypMjjOCk28g+jQJSm0WSSLwF1noUIZ/Zf5vGsu8GVP4zEt99dq4SEGx/
5reyzVLR2rEKTg6laNn/N+DUOUp8mO0A6ly/zGGCqFjYwfYYTaIty/oSD329E7/d
RvKkR3E4x++TlNVU2x4TZgv7AuwpgsR4QJniK5cdw3P1wTZljxObmrATosyLL25K
TnMbq6/2KlKp2t/DWyzm5dAkqQIJmtSsmAJfhGC+82reACYW5K9YUIvjBrOXsfD4
kM6LH//fleokAENF9YUE8xhfhIZqILtxCWF6vnti5WCmhfU9g+C630K3eVRzv9kg
2IZIGa7x9hPhC3DOLyPc9kDzgYz7W+XWY+MBkBetRbexNMfBZZVsOw28ZpeEUVTc
wUcXDqv0SWAyrxxckLsAhpZxniNA+rTtbtMcON/FumnaRV4LC/y3VtPUwG8fK5RU
p/IxHgKyZmk6Buj1BV8moz2XPDuHb0VrvOckSVAE+yC7CczOpxFoAo8Qu85Cv556
z/wOr9R/3nqPdWcdl32UcZ0rWARCdARvrnMsx1x34TdtoNrGai/P/CP/o3dSAWdt
yh7/URHo6FOGFjyrdsaB4TkoYSM0nq+fHO/oPEPze3VFJh0VcU7JZXbjHSluQmP/
pg6T//29ZDVWqJZKpH03ywemtoBLiQ83N5NHnMnn5mr71fTs83UOMZMeIp68y5ZP
10tIrLSBKPUOTud3dv/31owhtRvUFWy+WKeUZz16u87DceYgaDbDPbYkhn4MMj8m
h0Fi7n+YUTqPl1dHiduMZnCfjIc+b16nB5SNdSA03KDHCg3/by7RBQn1R7kicplV
Q8X5SZ5XvQ45OY1V/Ib6q6+rDCFcPDjjLOC22bL9HK5bVCOGlwcxxmipqa3MwwoZ
RPYrnq6r0/FNLQRiCQlRD3Jkx/7SznYXlTdxWyscZzahhLZpDLlp/RrstNhoRf5s
dDXNjlmIZsmrxv8SzgkSGn9jBjtZmIseeHNZjkiQ2hqbTiTc/CgOAx0jiS2cq/rn
EIIFp8CGdx7a7YkaSYMshJmCc+bM8wGY+2+ncsZ9zZ1WDR+pUa+A3/XjNmyfbDiQ
kBhnFQ+E+jD/WYl+H3XSkXKwLf4QwXdnQbdBLnZ1cd+1I5AsJZHfWyqka1x8jQPD
5PiICp1Xp+pFs3I+Pyj1EGZMGCpeK+wDGZDnULyZ7JfLajPhSWPvf0lrOannPxuT
tzmNlz1ngM7kewTFoiYSb+VQCJcxz4Vd4r8Aq/uT3N8DeaWRsRo0QFxVWIRUopcI
TQFfwLZCFDFRT5pzqhxx8yCL0A4CkcEx+5VngtwTFY65+awEF5smm+n4KwfST8xM
OASasBG0eK4GUow+Xx5Fl+hF9LotpzGyXz1roFZESzM0ESzJNT4B2BDAk1YelOv/
AMWPaDxQItkeF27rcuKRznOVZTWgmL15pSpupUuYS9wk6/brGHl7Abeh2xU0/uEj
EPgb8CgRwqygcUUok9GvFrzOZ7vnZD7He/XcJSl+UjqBCJCk17HaEM+9SPXKGZ3a
ULd4qCNjNW9G/3LqhuikQLCSSfyU4Ve2BV9Y7EE2/oiRhZcouEPQRfR1AIXug612
vdVNeKqDBVCe9/AVMXmRmArLrW3MGsySb65BgrxsxJIIclnz75sVUoLVw4W2fTI0
jSMJxHQnLBJgZEbeewYyuZG8HT03EQjQ+5sJP2q1Fccd5SYrflZdHfk2u+jCLaL7
/mQsli43fBGmkqfBPLoH3jvz3qVepN1XTLhOeMmJtZN7VYKnkMfNqycz/WG1TfXr
Qk5AXsxVyy31rd1uiNzzw3hTVIokpWjJyX1TkfYO8sMuQmdRpjv1psq3pQ1qXwhm
BG2g124OnPkwCZZu9n/Kim28IcdcKvIYDWCj2NUN8OAQ9whsRpx3cTu+3CJvAIYT
BAVb/J9sLYEDVqm7mxhfwMQmxHmYdrZ64rSbHOnzo48tKz42OesrHfflZQAruv4m
FS7RYg1oMmC/Gvh9eNl8t9gRWgXfM045XWcXEqWzVOgZynzynDzSqGamY3HwnE44
EfOln4P/r1eO8A/x2tv/XFl7Jsfg/5LKQ8fabPMgYkn7NC/7I2+rMP5CRZ1Q0agh
DMsHTSqRt3TSgLmyJUztGYRZOFeZbyex83Znk6IBIGvI5iyDiwn1Kts3JHj1df+Q
jra79KECQfpJysgvL8qialig5FOuVEqRSagdiwN0Ql2XCZ2XsH4rxV/dXhYWspUK
W0SpbbwuHawj934lShs+d/m/CHyNFFuUh3wEv8lcAiTZwFS4Rw6IMnOADwkzYuwY
c4nnjSYQmD/qf5hH20pOf6AeNtv9pLL8V+LGPMxq2Dr+uysAZQXsPs7ID3okjoIh
5FR93pJ6+y+hqd/Te4DHC45o8jSD/32lmRuqEkjOmcg4sfkl2Ko+IMLD67q4/YR6
hPX977PtO01uAupwBicd4R0g/TXF4mAk8DW9oKjo0hO/3JCWTBUPTki4LErdJFeP
qWLoLvkcc6+VKTLoAddurC/Nrkb/uEdlRQP67ezhB2vjD1yGcyfsEmE3F5CYm5z8
P4gvOEduylDv4YB6wRrawxOtdh/v09dtbDI+HJ0jO+NqFrOg5XZ6ddhDpBpCTXdy
Bh0zJxtSQHbAyy5x7+G40o7rYKCJ6poVc3HHyZyOgJxatKbVyOH/6VZ8KDGEbDrs
gzJjCRLMdKsYMrb9oFSQ/ezPNyrxcaH+Xsc005CEe+Ai4Oud6kGBzjvXzDYHNEf/
tpIwMFZHn/N993JyCtXi2772KfoTvFhQtcHBmwospoQBwp6UK5zcOgoaBdXT/Zv0
NytBxvCXR//vlc8nBL0vGGF7SduqSnZUM47eEBETcn7ydhzxM8X7hhlEZgl8g64M
/M8dg1iH31VUQybaIrDEjyK3ZOpdXN3FnhsuxefDgDaBfDJOlseqMHLuJyaUpb0b
3qhvk+DrU4NGut5S8QphOUyRQQxR400ts8zB/oZ6t1Xh1V+BNk8p7IsO+RPsF7//
NsTZDWGIKKAd+dD0K78KTds41P4KX+6PYZ1nvnolBf3+6LtAwTNVfVQCMgaLulw9
dJjREy3oWThhnDeX21XAgVL/DLrVLmGeK/XBwSKAJQjIUXQO5xDAe+cJ4oh0EBB4
uXhVhXjnCgxTQgZMD1UXt/hQgUvwn/t8aM0T9rard3VPK/w7Os9u3uCOJ1JLLiiX
rFDDLswvftSYknksAkhO4xuNflqRtW6pV14llPPYwZ21gz2OAVVTUl1hGv5n6Xko
vC3CUIsxZnxSSvYCyRbKHUzf7KIPyfGOaPgKNsq5o3A3cn7JUF1ZmNWfhu+pa0rN
nSJStUUgEetc+fLxmRg1HFMv/45AJbw1GqqllkEOiOSz2i7ZlLDZOC9edE5QiXiJ
56m4A1SN+WWUVav90N+83l6nzBVFRGdaNvIpdxmw8XuETuJUHsWzrQewHkU7I0R/
CtZwWdhkTXZJC/zyZXJNv2F2jfzbniQT5Tnjh51QVyRkPw5RMvFQZwxSToLaMQdt
Md4K5nUVDalCx1hrfAFmgL0YL0x3z31f9iOlYx3HcU0Q9cpAy09yUew5rbBLGOx4
PiB1FUas6GLENEEfGFUi6yQKSkFVd9N+GCZVXyYftVonFZ7u/kgK6X2OxeMjdJna
94fOJHXubUD3bbo2NB1lVUNkJn/6vSyaNNUGfyQCSLZFqGtYiomuzhFXQ5yHcumN
bFgFx8t8Cl7jZesg9oeFp2Ya6gys3/ULWMg+fDwfBXiLLVz8uRk0aN/GL0BXuHyQ
k7SO8VU0SP858+2hMTu5DjoSGEaBi7N7rFIlP/dtnYEX/0h8V58hj8CmCMyvl4mU
H4UVdpd/ZVZb7Ow8CpC14VnIY8IYK7iMKYVlcfPTRasJR68x8sX7ueFNxe5JrHiq
eJ4WECwNBZvBzqq6xDYBq/8DYfXLBSod4pS7xvjkUQQV6QzmKjwAzokni7aUiuf2
UqVVP98ZXr1a74wiqikrC7Ss2+riw2kW+1k6u+nUGqcesiAIQuxgBeWxVNgLh0uI
PJREr268BcEBRGvXLoMT3LEw44ZP8oKR4AcJVCVB5kSifwCZBNOasDvKOGAzYI60
VcrIGIHW8iHLabYiQDoZCq6UNVPt+ZPN+8qOinsztv+BVwVmr3rHsRhCmFPhTvWI
QsJ7gFmnBo/ZAASXHpSgmNfIYeS5jSV9ZcpAZmcqQBGDAZE5NqQsnTuNgZiYtq9A
yc15hmcSHhyALME9qDnD9/rtee6LJYpIyUDpJgm6FC9BVGB09OAzdiEcWBDtvQ4K
wIjejW5RFphLxt98mFKovjgKYdUeNNYfhXmbS9vpY4LQ+TVoyeYyvsMdqspWvizK
PpAeyuC6UFoh+LhLs63vf1ehcx3DFYuGXsYd5gsrNlo8i+iNOnv82lxJ2D8G4BXD
0Y5X1ELlaVdc9Qk6Kaix3jvrnls754lp7B3n0TgYX4mPG3wgChbF9rzWXMC8dRGw
rWFDaW8riY4kS8GJKugYVU9aKUlxET5XJLj942tJWCCoNcx4+v8yXN5TBmtX4lLN
j08t+U61cBmvBf7UYHF5BFVrLJtN3vlM7tXh9aP1D1yEGdvK+ZFS0RfCV9gUkrly
cJTabtrJgs+ojx+MJxXXx54tGyyJhyUkZdehDgcCZdtgT/kjAycPZy/uvOLSveHJ
wLo3FK83DGKOltTOWyXmJXfmlQTe5SnWpevzwaO9cKqOWDCKMcdVAIkwPv0F2w19
7I35g0iGZXdoN4mT04JGXZxa5dOhZiOUJ9ZjCid4X2N7iWeAklPU1E7+EBGvGM2X
Zt0GwfQZW8DSKI8ZHh4F4ujFz1plseVAi7dZ0IBaAnV3iw4qKvRntSQyf7QFkog9
`protect END_PROTECTED
