`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XiTQUN8RXG+b07zX/rDVryTfqjiAJ8DO3zTZdsk+Nlqho9sUgd1ytNHRj+AYzg0Q
cFycYoUOPeDBjL6XOqKWcwB6yS37dgQO89a/wHnSZSTGQl0XOoGvv4Q4WDxlm1it
bUnFshfxo0xyhigc/Xe8iUoYNSFHxBHjkT3APbUzNUXRgTzMeqFNyO4zhHHpOQdU
HLeYkzFM9iMtPbwgnAae7B3stFBAD81E/6JJBpYtvOdj5z9SCv6J2sToHDG+JLu/
y7N9MTajt7MZpQ09CuEDHkti+oB6T1r6qkhPMwUqC6ozdLOL+XPoD1/27n8RNjFX
Euv+hJz+l6WCXH+0v6fPOhZYsorJRPays0u0j0UCX7emnK9HbYfAuaj1dS23+0Eh
P+/egcfUTd5QItn/+KGahwYVhjdDQ9p6+AD97SLhptBQSQpoBMW+t3Q72HWZBl9L
msKWNwzp6VgzL1bpaFU2qqbmF30p9+70KIDsapY6x6iYae61xXzEuK3yFX5wx21a
MsUFBOZB/b7lrwfysqM2iA==
`protect END_PROTECTED
