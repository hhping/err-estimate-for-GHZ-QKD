`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D3S3R/lh+FakAjYxfD4gsqjtyw0+PhIWVPq0K2ATP5h5XVDR5APQaV5vLcfEOToN
DQLOcOY60I8ppA2gwiGY6603dtfqdYkCE68Q8a3NIbGc53ognYukimggWuhHXLRj
ib0S937RPXQCtE6/N7rgCCOsvyfuSQRqNAbXJbnioc2WRnUpGjbo2aAerPcHbzV2
Vneb1uPPoHthd0i0CRYj5oCiuOnsXxcNzcx0Y4w3m/rl3yJBuyGr2bkBCqJQB6gQ
zTcmKvX7MK1UuWfexrCG8KMT81pT+uhPONJt/fnC6k96Fpi2UPrURH+FcrWusESf
dz/3II3d00FIiBFY/O0YgGlIiVwXmFwbRzgBBRZ95eMkTqR26nt+iGiEdqWLmVfM
2cNfdKTxlWmklWnqMbT39kNqUgxLJ4i/IuD3azWzQ1EaihGTx4vkDQ7YUE7I3ufV
YENXLcBgvGdaVR1dmXCTG0hUwe+6prxH6vUoliD7m1KPSmOPd8Az5eVP0kuc+7yv
ZkxqUyKKg6bs/LL2EySopUl4mr+cUFPoF0OJ1Alfrf5/OTMaBMRaVUAJicxq6ywR
13z8yP6wqpk/yBODXQUUlxA6z/n+4GRRGLekgiYLmn3SHZWxsNNnN4+LWY9T05CN
Q8A3vVwDsboYlNROh+S8yT/gw2pBnqxXgzvpA74BpR9h9xET6aCX+TGB1RZ7l1gZ
tM/OSuy2j4OQ2h0fwGgeIZXcuvy/K1ZMKtiUgudM5SgPvs5pCvWUtz5Th4+Y9g3W
Ci+9G8ZC2dAALccRqXMtBD4KVwC9cxnN1V5oENx8/pmSyyobaG9rTLkBX57ei9cP
rYvkvWD07V6ICDahlCBu3olviMzmZL5FNJy61wjaDcK9cLL6R9UwJDDAhz5qCVLr
gkH8jjv3Elo9ndE9EQRxbuZM8FD+kLWWVrnd3MrhIfiScM0YuYTVqpg/Kn48LT+e
OEkwI5GqnRtne817Bi9GNvluNV1C/PirsxiUauyvzvGaYkqjNB4ZwlDLIsuWxX0k
FNGHVd6ds5ZECFFt8Fr5AQ/ID1xkVQ0do0G0AEeCq7+XQBaV0lVdlZCD2zwaX2Np
khW7fnCIqTktOqxGL9YlEuYj+o9gfBOi3M5Ggf4ZKcZLsFXZCiFEye/VlVYm3Zt/
tKDB3e9+B15mmwr+8Jhekxslv7ex2pa00beuOLHyw0uyt6WQe5jBc2Dzr295dZrT
fYXeTcUgqcsEVME2j5PfkudWWUwres4xxBAcFCWiytKGEJHraCoCVF4JSEKyYeAB
ZTxvTBZEYBFVKz7kaLjO7UETveaDgIJQ9IeduN7oxuSLHThio/MfMxZ3aGrvW6tm
qDM/+KZvj/7UjJug2NJkmjGmtISz6yLCRfbMYGwYMh0WyhGvOk7NEv2ibzBPh1ay
+wTg66Z/UbTKmRsv+KqtIaOdODCXQphbSMyXkbROdySc89Br2ui2E6xLF9UD/K1y
wYvWlplhRey1FnMVGxdBDcQft8T3moJxMumoPyXgrVCQNl4jHR2EC+ohb9qh9Nc0
/erPwDQEbQCnertdeTtxr0xsmxdweaSKoZv8B1ZAiIHaocqi6vGO1bS4Qj53OU2b
Byh4aMibDrxrpjoWFzmCmdvjuznxiBAMgPrbbDaY2vQgYPG3uRaX37fnk2AHbSoV
ydFreaJ0Bc6NAAdrlR/+XJatDDlRRwSTdLlAJcwi++xvF32tXoctBeyzLdeJxk53
EowfApOLAVGL3v8uKOdAcdOGXRUY/n9C9oLBn2DoXsiNP6xgwWxKtwc3AhFQdFg5
/BRwD37lmnQ9vGOPEthSeLfeSOxhCrDweAT56lLpZsPCT1xoG3jdRIGni+7wzZdB
mgdZDNFcrjNBuaqrMSa5HeWfNXbMQiAVymhg41tTqQ6klOm5MIGiE05bNxoqmvjo
e5VnFsBkAy9iarFFY5kCX/fz9+LR5GVXH25bNtof66hDik2nqXVs6ZCX+yMBgNYx
RofN6RUCSNlj3I5+s0IiVQ==
`protect END_PROTECTED
