`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uIzGovTfME0FZ1ZNrD4/gJn7yYcO/NR9nWiePC+o84rTF6CxEdspR7VoR5y1I9le
6dv6hfOQ+2XynnUhSaf/6kNM2HZdLZ0swTyAEGktuXhdEjlzRIsSNxGIyK0GK2x2
0jta3ozAPqSH6WT+LJfPQk9UtFknPaFYTFEHu4kNVn2X6D78p8rAycNOu4RkeAup
tQ2c/1vXCUdRZaDeEj7+Swurm1CllcorPdr1y2qjqKjHA8PAslVuntPrDB2PkxDS
GSqH5vLmetO9cNeCTPmLsX8XqNyb8uYWh1MTKfwuVls/OXfc67pd7Aada+seUT44
KkONJ4KzNn2cOYrXj/DSZN4Wr2YBLO5R8xUCMddSwayA/yoTYH/dnhRzXFn8WRjj
Jp48/xmuC1DZXs2rUwLnadiqWw4JtmMHnzEOwhoiCHfEfgZuyHmsmOTZ75jPgAaM
pMXLiXrxOKvlmRDkEdzQDGIL4VLfk5jsgI85mWp3z7brvxf2fUfAwXiK7ZPPbWiR
P0PJYu3MXER9AdhaNee4PSiuyhn/h/DFepHKyjV8zMw+HZzpxpkk+ENNIrE7/q1x
hS34ZIadd5EHEr6tTj5TPEi8NrMAAZ4j5IgayXnOFIQZFwMkjUYAlyenRuz7WwU7
Nxm2UECfpdHhGucbYqJd+tGDbx2+QzI+6afVn46kSbZu8yNlvDUmBnLGAzUjd1k2
bBBjvCDOsjXp1FZbvqumKWNxj7pJpfTU4m9bPA2/wihWzbEMqDfoBfftLZycs0bA
lqxza39xb7/oMrhdhRbkRtaZzIreIN7ZCg5+/a/jhC0Zwt6Yt4Q6sDKf1GX4nk8o
tmTyxRIgW4erNbN7vv6eYZxjNbpeComRUaqrzNb66h7P0xDs9g7XTkB10cyTZwen
ZtqK1nEjEBLkXOkD+S1V33/ee8xXKiZuXhYl3mudFyErgmpMO9cvkmtyepSuk8nj
e7A2OMczlkL89EcN3lHmQd2G6Te8YmnjZNhVRmCfhnRalXjlM7snPaesp0enhCnt
o4DtqQB6I3ZgTlwM9Wr/T/TmktuVrtU0HRSVx1HtSazOu5dZE94V6bA4LDUei8tM
mMoQ2Sjj/H6cz5vn5ITVn6kBNgWYsNB7D93yFFRecKVZliG3O1qt0F2vHvIfbDbj
CWtDasJwKEYwi+AGuVxmNi6kPLchrn+0s0YYqM8cCZ/0iboB9gOIvonb6yaMgtUC
ATe8YVBkNQd5DJK2wSyocVVgW5yWLXlyCoqcF59J6EkMfty126FV6JIGVraPg7KM
8njwqxhejzyUbFqWFRSnQa25rfc2nciL8gJPTD3YRj/2FRlbIFCbKtGium6TYmRV
BRW+jryXWfue7bNe0dPFtxi/csbunU6nDcwdICnOKaejQ0H6CkpQLZvVCqd1ZpWu
Rf9UqtN3yYZG+Pjb9lqzDkw3tkRWF6C0mV8rokTyHrkCuT4MxXvXgWnCp+CS3lYO
M8+C012hJikFVvYMcPob0p7zi3iLw45ePQfXW4NVdMXvaWoXXabcjfLlBmOpsqW5
QToSs7O4wBau7CyyWPPN1EeZ7LCtwwatiA2DxQjbDQQ5ckEaOF0Oaxk/fnBHF0Jb
+UniO2c67F9BTGqDfTY0lLvNTmBQkuHIQFYuNmEpG6VvfTpI8FrSw9l5MRfHALCN
CWZochWxvPCcSkzXwuybR65iOs6YPuOACDtkHZQ1p8kmBlI1zZQKcCSwyxwW0eXd
XYIuYTwUkal/dM0mnA+jNzgnSA9SgKhRyc9TWMleDS8g4rI3NTBvSZ3+LabeUdn7
WX/ytp7qvFn2wTkzcaQ2sIZDXkdZxG/V/olhMB48PoBm0xExvlJJwTVpxDLCE5KK
UA+oOGrtTi/BmQeVvam5v02wlCwqDLHrAq7yBItfZwdmRKANhxUTVweoyyyyQxMK
VOSWxDGHTZTuUPaI6F944SGYNk3S1X7oqoXN9YeYkxqkm4ae1u+3UMEHv7FNAq6d
60tgNg8nVt77kzmNwBxw2uAa1UNyHWR+dzdl18f7ai1O/tv3Y/DTDDb3JZKLpPM7
f3E57RbQGPBRMS12gdh/NCIYp4c6Eap/Rb2gxsSsjk8tf5wMDVNmlvsAbVXtpOKw
eAuOoc4HOS+QgaUgLFTcxI1vHyrplWv51Gv9OrCwWTkDITl9oTnSsZFk1WM5GNNR
5goAsu33B4aS9kgVf4pPVgtCJgnR95N9RpVW/jU/hcZUn+4y5xySTdflZXjCO82k
IYDkxBhm3gfyfsz7gQZKR11pTxU5SZv2dXq0CTiN66S5KytRBSVrYQapL2Dc5UtS
X7Ujdr7XeyQ3m5FdDsQBxGBo0yXOg5HjLy2bQKa+sI5lM91+LKsodN5FOVomOnpM
N9El7eZJ2mEhjt/s9LSW0FOw/ql+crhozf26oN//fj236xdpvplvfHYWcqGhaNbz
QzHZwRCtsfLRRJetB59si4lPmqaj14RsfXpB5r3M7DzZANvglYrJ7Rjy1WEbW6TT
b0w/NM2qkNogLNPF8178YLq7sPCDYYRicqlVq85Fd4mAf4FAU6XA6+5YufI2xEvI
wrlWSqte1ktlujVbnt/q+Usi7tq8Zm0ZnUfPa2W2ym+rHff6vPP5o05oDam1E9Wr
lUFfs5hhPlkBaEtbjxZN4lmOtQHeR9PeIGGloVFoMf/RWTCuRMMcl1rEmvvA1Jkt
LP3LsmQinkuqoQT/VNAjbF77lmFtG0q6GA1Wktk1Hd3GWGCiWCB1cRC9C2KCkGSA
J18Sqx+NaRqwvjhijLjf/95ThLUUMq8+OlBLvFbzhGLqlUi0PFILGwUgRT7Caj4V
W+ghUe37OZwfIs578Y25Z3fttuchNDSRXDLkx2jcjAjQUzGPoLUqO5RXOmUyyXOq
tbbKCsf2sAYFhecU5ysPeUjndyy/H5A3mEjGleOVOWoy7n7QRrJYvwi+hjdjCZhS
sTF//cFKpjU5dCDVUSVLnXJMPGJL81rrHa7dVz1kuu687OTJ9Q2lTuJS1jFTmwF5
xNYyhyZO2370ktlhv9F6jg4f64SHmIYPDPjJ8yE19nLWcO2xLsO7ImgV/cJk2YGU
4QEqP0MMvqokHOBGOGdtXjCBwGP5B60kVStNY5Fl3yNUelPf6km6GCrspokn5iP/
e2jHNM+kM6Mwc3lLY1xjwLYiJtaplXQwxU1Hg2BkhUU=
`protect END_PROTECTED
