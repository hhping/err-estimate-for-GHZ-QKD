`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eNCiqdF47X55hhKEIuEu775Bx1FpHPxTt+vt/oka/AHSXMZ87rkFe1r6ZN75S06+
OdVQ5w+9384amdiAxDJswrfJU0NLbKhwAdGq/rkFLcF3C5WcxhVT6F/HnHaIgio5
sjdAqunUOiAwpUctziOuLtIzNOwd23Wl/RQB/fxSj4jYZK/moKySlLIaosWhcfPH
rwt6yO/o0bVl+FdF8T/ZZdgXkb9a94/F66aChFllNtcYE+wo6gzPDkbCLXiLjgr0
/o9CtDyCt4rrvwnRg7zrbcp5HdxBShoejW0dTb5S8r2d2YXmo5kC42x7IYknmWiH
3BtFZmkrb1fEUBSU/y+Cx50bll/Y8EXo7IayYbNzyB4CBDQ543KvAfVZ5A0jgONM
u18GRbfe3uSlcFTrqs+zE5OXWNb4o2abPES+/dFzxBZv6iIqGjzQnBuHUTz/T6YT
k04xXObcTdz0TJNXJ+3vxSSMU+W4zKVceHqZ0cJtaruD/jn9GyT8OMzShmi5fcYm
GdYlZmizef3iPFS8yZS3+OqhSeIomshtYWHdA+pjcm4t+sx7IEu2eYk0itMvq87i
2jpFRCqa2O2BiYe0j+RHLXaQ33WjXXQF8JdYxqoGRg0h7/6jnnJ7RCYOcaVETsFK
cdWdr0LArAwj5ePe8ZA/fQf9l5ZduonzTAxM2OOyJdkfP2V2Rw2QQue9AiHEH4y5
cpgF3vmBX/o1uBZhXXe3CZHPJ/hcd4DxA5GqFqxPJzJmPHlNWvFHPoKtd94pv9Ob
Gg6XIIMqYpaNO/W0qVZDji7d9kUUhDYPrYA2YgZooUI/mg03KMJAInvwVgivSZ9R
zivpuCpxMHE2XQQ0kP1HqCSPmqFPpEpfQrC25OnOErUQ2eLPuQFdRm2zCB/fUGBM
exJwzgde2LgjxSwSreEXeTf5K8welXoytzR1rZBj1IGaiojj5w4WqGPvOF/yKsht
TEItp39uHop6DWS+uqh5ix/fM1k/19Bg6rJMGQ9Bkx3piVYs6g4CpnLdHdaG1rGT
pmZzgLRTwKKJHE4AMtvF4zbQJ2MZQSTQcvMw2bOatwXc+Iu7WnPLW81I1V3kRRkv
E37ja0ETQix7PqRQoMozvptRcDK0I571gTYltfdgTOS0NiS6bEhx0/8zhLIqnEhx
`protect END_PROTECTED
