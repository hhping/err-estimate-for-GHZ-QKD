`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tEvKMGbXkN9Hc0p8/BSdNVC/z43dMPnEbLx8DsTb74aNH72ZR94oVNHGSRMeN0R/
wwl7sCMbfoBOqkHuFija1wITxD85Emphu/z/gdc2c7dgyn+VG1mzdX0AGE6PomhD
qD4c3AyAv9vt3rVkdGXqYPTX8NMA+w8LYvqVB+tXcqeeNYAnM/eqyosNfXcYhnws
yxtXpHi6NwdN2gNCmtgk1iYOLhHypxHykkpGEDb2x21dvx+EaYk4PQxOvOAcp6Di
WBzeQBgcTRmOKmTnjl2T8f3w9N0MilbCECfUmF39iiwycjA3lB7lobraExQg/0DU
`protect END_PROTECTED
