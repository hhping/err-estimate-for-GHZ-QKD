`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
abw8t+/oX/LYIeB85YlnQ2jsaQW9cET5Pniclwd3V0YlcAxqHlwp5usZI0WL8oJs
pjKTWolasM6MAGmaOp01OVNEswgPl85Y94LMrFihTvcU46PLbx8VB2ybB3pqC0ZC
5xOSXmLNpSDyiCKfA1qCAQQ2rW0HZwO9Jx8GVRuXdjlGzOoZvH5q6Tqb6Sj0qzm1
OOGtC5ViniXnkahOhQoyUMol4sSmg9524P/IzNTqv+yapgIiv3WJr6wnAa2MhuDW
bwvuIL6X1aekKU/Pz49DSHhxPD9HL/cc/uWE5lVlk7rJmfCkZgIjJVaLc2AtdaqK
DZOkI6bkmiHJ8bCw7bbgRWmpLVPFHKLnLwe0XSe8ofevYgn6EcjbETGQBLcOgTv0
6mIadzTh+qaBWznr+oDq1eS/FHpHdD4n1NaMCKVgglowYeA/wLLeXbj30izZ8R1/
DJVUe9bgxNbKhY5YNcmdGKZltC+NXA3OXXaxjX6+97ex/R8NH2MdiyGGOo0fZIJW
zqQ80Xp49RJzmchTl1DuUciEK6qj4En0py1QbdBTyFnKd5csrKE0S1HOuXOSjoO6
8JJE9A9tqrM36rGFxXXb/2V3av/I5ZlBIs3zQNEMtGvCrRa4rhzbfFZmU9QNXoU+
q+eMp18aCPQ6I3p7ogVINVPixfEWJJyp+JF5C7ME4nOuIuXWeI//M2N515vg5gm5
xlhBk7s8dFhbj4hEyMburobUJn5kD99e9q5gHxGvBPs6iyNR9Yc9CagJbHtVF05q
uR7YP2HgrD5vJ6DrTdQDx7F6s7ZVRYLoHw90LG2QKw1onYfroVWmG3fNkcI6WN8R
uHM3RWDVoDldkuwQzldsE6RiCmfkw+L2LhYboqrk/zs8e5jUrjOvFBzL2ev6xVzE
2hIxp6glgpvlsOsHHgjgn14Nh07VT08nX2bK1Yhjn+I7jXBjCyW9d9kaW3pRixKE
PesSjelOQzQMjJsk7gPxOHWdLY29Qs9NQsi2Ywiz4SxJmHvOsTGOoQOwJGNRhJ5I
Xv0/YTu8N7sxlj5eCyEmbg==
`protect END_PROTECTED
