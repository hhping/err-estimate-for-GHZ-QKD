`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kU0qrpzNEl6ScF5E4sSjJzCDXcudtEfi+6ySK4+0OrlkkaMrqYRvRdMxq3r4uGkt
7LloVSyWrLjgKBYoMyyRACcUCzv7uuVPyt3cF61/aYshVesft/YnScI47WYoxdYE
FgBKK5dIureDKECRuSXkwQj/2JEuxqOS+LYQt5+Z7SXu3nfC1yykZD7y9N7NnXmS
4oOeZ7XfVvrUvqTjNBzT2gURmNryJDdcA4S3GzrTf3ACGNys0awvf3D6y717TgO/
UzaSQV0YJ2nyFUISWFdafcmitVBClQ1GXaYea9kvGg5U6oxlXt8mIbM7WaUcfBEU
S2S56RvKUvBjfIxlFC2A6PJnzmbwQa43ddSbdUVHmfX2OK/5eh9IyTIS6MHSDfYK
AfIZTQV9s8KpkjAE+lU30H3Bgl/nqBnq1EeD4RHIy7GNTdX5ae4NVbbrMtmAKCOy
kMI52RWUWfXf2XojEU3OmkX0lsdvhv6yA65+zZCaP+0v8wINovVfGn77SQGmd319
nZfrgke7nxM6/iuwrVl+r5L6/ltz5ZCvMEtfRUZxiBJ74jCjCSvX6UJqFUGEM+38
ZI5VfslyUnvCn2LK5G+6Xq4CKy/StAJ5uPaWRwAYMZux5IJl67/m4tzG34u5nN7r
lTjG9m1FpyctVk3QvSNX7t2W7Z6pAoSxdoixHnQHdlgvs/2WSMZxoB1F0CU+fM05
+srhN3ogygTwEVnD094PsyCPeQ7CfBr5LzeGfY3+bs7xp/ZdRWutuInpnaOCcxHT
`protect END_PROTECTED
