`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hwdZaZM4lv0zWQNlHx3v96JO7PwhZUVr/VSnQ/1JGorWvntEuufoUZY8FIrxTsOJ
3jPY9z0XXp8fakvPRaoeKHP/OyAY/fxmsI3M/aMnsUSxGF3YuYaxspBOPKbJz1fv
U4y0oqUDb19XgW5Sr4NLrqLwL0UnTrEz/e6zWz/k3iPmbBmkSFc1tQXhzmJM8lzx
a9tYmhcsW9tRc/sSjPRuUFA2Jd5ptI/n5fGsoq3fNczVSaSSCzUhB0sndyubjKyJ
owq3yDlaRIZPgfe9QX3mZe3P+iZTnzfeF6xZTn3R0mebvvYbvv0bIRVWTNlT6psd
CqKZjBEYRHef7Q5nVmquMIK1m1C6OUTIoj3d64VEvPd5JNE+A5KnWLnu2c6dKpYN
OtT1Z+DrBf5/HG9a6LORe7+wTVvJO8TchaJtZbm+xJdR9ZXkM0VXfIrKmlbllDYU
a4niYBXbXUA7cIn2Ggwcav0zPE4PPy18P+dvgSy+4RfdkHn1i5iqO32XdfkIKKVM
Gz25marnrWX3O1Vs9RvIoLI7yL2i+EyLfaiRPJBBH75ioHVY53uqcCmV4DBsd+ei
KqFvDC8sjF1THtw1Eif0+KKleqbg5wHDrQvBNF6MlJpdhRnKMy1vwlXuswOGKsIv
Q0lKRtXqfwdRY6LmiKIcAO6mEO+WgBUZ+HCKOn6CcgGyvU4PQ1uooiDgPxVBG4d8
uk3cIXeZWxYCaqTbpHiPbU32h5IRR5DRRJrdQif6OnQWgw3gij4cPjj8WUnaLbxk
ypancYxt1AioOy+U7Lg+aHSclja2ktPgYCFeIMzXFhijsuprU9jeYAtqmhF9QHgb
Q9DxMnWGBsUBrZDaNOZfzUL0gtZVMR82kEf4Y9dfvWfMntGreqOL7LZY1cbzz1ok
mQ1LMEhCnEgjwiujMpT/1klhkFnnuQPlaWTdsk6e1SlD+vyHIZ3Tapw+2g/IK9aB
5RjaBh2+FJaaymuRLuMd8l2nV6UmxfhWYqc2IxxvCGQQN4U9/J91IdVyutovF14H
vGG+wVUpdbYnsvHryEI26hwSraT/gBtFIzfN1yxtsL2xvc57z21yD12bt3LbYO+O
E1u8MUjCRvcNVRavUC9QQKVKhR6KujdY4oUL8DGnHDm/O0FPFljom9IOTSWA1MP8
kqzLcqaj7u+sgPPHu5LyzRf8jyiF8iD3oy9qc91lWBNfA3D1xk/rntA8reONWvwu
/xSWbVsNw4CMyioiuIaxkkDlXHOuCTteJ2cA4hSSRZN9srbjGPtr4mxf74g+QKw2
zpTCHMnnUeklT2HV0RV1ljLUP1PIiTu64dIuehOLXMwwBMsuzBiXE4ynFBiQWq1c
cbtXJsvE1UVXaJu+5FgshMB+SzM5tYQRSDXvOjb0YKfeQR6pGRitXW3K1nzMHwBK
JXeY4CtV5RJE0p3/VDDWXPl1MY2qk6MIIPlzYKIFgBmsKHoaWDtw4qdo+wHPiR6y
4OuQKlBWtcgFWszFF78DtM4SKaCFPVYc/fL4b2ouFe9q1i3QvVHgTicyuhEjWLC1
kFu1LVp4W+rzGI0gxLPu9OLWVkz9PAUqOS29nzPF4igLyBj7yQP5WJ3ElKLsm1gf
XLqjOLuyaI4uskzTIaOqt63SBfvCBC3sKw6vWJbPWPyvpR6y5K7G49/wqbkVVfZ7
kyuexgn+CR87cEP6hrH9SidY57imQvyfOf78/u2ti8fhwrIO9rOUFSnU3hJ2NMsU
T58VitaoBAorxdA6omEsTQ==
`protect END_PROTECTED
