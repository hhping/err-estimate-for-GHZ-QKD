`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QxuSkFA4S3TNcQX+QU8vG5XpVmUNc+wH4FSHUNf0r61aoQr3Qju7IsB8cqpxTUzs
p3WTuiK1oM5kCPJIVFUdCEQBtjRjDEeE2OwY1F4m/A6EoAeiMaYeAlkZVjuFADMz
VKKJVrCGtGsI1eHeSnIik/q2VHhjXRIR1k8GHy5+5DkJs6Yg2Ja4fuGqG4kZ60pI
YTt22FKsefidsE5T9Tprm4fgCfsVvbTpPLcjA9PTavXgMx37l7RUhEMn/OKQwWh+
sFI3l/BeUnUTs6Rg751VgNtxuKt9LsV8og8XfUZM7pnUf9mPQyc2GqBWo6CPQbJD
EJMrqhM/zkwEXgz3e/BPGZmwbnch1/KHRlaELwifGroNpDE4mY9XQCjL32lGcJjC
xb446vSCP/Nh+xkNQc+j46Xbi4z++i2lmtI771S3xHKcgP7vNQFM3sF8aT+0aYk9
zXs/qg2tvoM0HSc85Mw+RogHoG2+C2TiDqh4Bj91ts5qe7V+z9FeKstSH035f6Ee
xXQpQ1jksL6nw3u5uWqxdiWFnfr7EmDgGXUKh1BczcPISNPRvFRIEDZMnnXbH2QB
CZ8guT9t1shY4MqvnCqeSw==
`protect END_PROTECTED
