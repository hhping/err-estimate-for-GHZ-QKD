`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j2pao1DLXhgtdi0rYaxTAwuPOGC2mswqiYpyzqQjmXkdc5Uf0S+b5Cvnmr5KpANL
Wy3f4iS8n850jntpGXJlSkBrpg1oAslpGJLc8bKHSCjubqN1Fx/MDS369qP/GhjD
YErcPQXEg1aeR9u80GlLKf8dqu7cg8r9UCso1IYKf6+WNfhxaipPlhTI7Dea12x6
G4R1ls8byAwYlnGWHIFvjWeA0x0L1DGwIzE8u90gOqBcmD1lW+j2RsAory6sjFuE
7F0WIHj+zcU/FHBn9KqwiR3zv6TwqAkTGHItB3g48ow8WbzcRxn22AA9pFGM0AsI
eLbb+O/eMVMcDKmAGmKmjxbwJWKIZiTEv4svu3bpBlBvNRe8fhA98W/j8Sh5XJt+
K9OQFLeHlXJsPJbw4n36UPmb2WI7T8qpuN6XYXOlCugcIYerZNAOgQnEnoNE+ms3
pu8EsAURf3jgVAJwKU1cOWyl60nMcAoVKGB0Sm+oA4msQbmXazAf8/g11nKmUwMx
E7ShBXhHlimTly+cBCLqhJG3zoLqQFsBOILI+7MNLXoXUT00mN88WEe5C7+r5Kq0
1qPIujzoyFy8hXjvHXNYSC+EiKfmBGyhUzbaDPAtpAELI2D24hRa9E3O4mnawcHo
3CWcfaPpULMekcOjCYMNWSlr/AaY7VepHm3JZFK85U32T+CCVa4p18Lc4+PVW7Wo
RWQHph4PBUmsrl5FTnVeT1sqeXXk3VT4ELD3POIsIwsTSSlaQ82Xme6H3hOoRKZL
m+nYPuoogFStPFf74p57MjSLv5EaWefJWCmDtiwgowTmjzaUmMLYyXBESteNkHfg
T94RHjK7r0D8lozIPT1bhX+wYVp29jypRl06J14eImMKwO1pyy2Kpqcr5e0D69MS
7f5qLYggHau7pKy20NoYbRyhAJV1c4SV6Yp+2yFYZlc6bCbFy0TdOTjpsw/2cPs7
ThIUUCkfcuSNP9kQG2dcvWah53dXOApsIscL89qAf/ElLOwX9ZNGRV38UWauwEPe
eICPqqUMx97ELjvGemWY3pELeJnyb/jzdAYX7Fq8/wVxhgAFJsTjD8bqYCmoFGAG
S5CGdJ0KcZ4wW8mhD0kjWja3btqF9uO41DejJDv3euKRXt1mcLcOTE3YOlAxXnnN
+WAJbBLI3nhSgWeUJEOx0g==
`protect END_PROTECTED
