`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5vQ5qEGT3goTHVWgTHpWyrUgucdhgB9zjvG5QC9DoYWMNgrpF148VKQIu2MuFj1m
ZrZ1GYuV+86QLKgCJ2JqK67kstQhACtpd9jkxxMoYX5tm7cuSiF9CDkLpbGXaxZJ
28ISgPjEsqqSV65KxSr58CvYTvfdXlWMHWCu56h/N3YrkH2U8aquiQoq0nuB0bS9
1FPo72PfU1S0b/SSJiZUYaKna5D+LQKDwHOsLxD+d6lP2LL3QAByJG9POM7fh+vy
XFR9mP9MyjyhqHSGAj93KPjth/pFhyy68hrUg/aLWUEQ6sJ+InIwdI0sGmlGYx7o
UkctDsWlWq1JkWIAqNZqw4p+DAsUjrjb4kUwlzVdy4YN3rL6c6IGNFw4/dHn7K+S
py4+htmYXLffVh2qtYo4roC8NyXpEI3CXwfIysdPHTQWrN2OCyE1ZgAD7avDPu5c
7aHpCGHA3jX1v+JTJO6CRu074e7z6J6OzX11zKA+G7vFgdG4oUY/21lYMm54xdCh
0jlqThekaK95AtUkGyEPk7snj6mwM4rh2hcn7h2oYlAP8PBChtMwi6/RKcjlpZKB
GuZjJfj6KOfoiyJIpH+Knu1OogFf2o5hEYAHAlsfRh/QeSc1L+mrfdkopxMxWZEB
xsrti9ghFiW3TBQYLzry43OCHkiPke0hqzEpurriX43Dkih1UHKsVpZhGzFrsvqk
kcesVzz1li5eBezRrj3l7P3+OorSYrywmiBAxw6SntLrlc13Tdkny9jluC2apIJZ
0ip7zb8Qq737a/g69nd36mwY8wLhrezPtxWGRY/Op7m747AKg9hM/mTUDhM4BsDV
tDuF2SrkY2+REIZc9vrIttl5ZoOIi4/eRA2vOgph1tzg7hkFz7kmcxWWUZopvzoC
B1JxXupMvmUxsKCAZL5voCk4fgGRvCTvpnBQHhmeDQC6uZ5Gfd3tbPuyYVRxh+ti
CvXBdV8VM5HKDRyj1lCUc3Ln5bdBjlI5L7dPmBHsBiQ/diqPK+uH+oae9sVPFefU
bghWzwEVpLpL0ZX8r5OP49STy3GPuY5EpFbJ7boLhR/4JVDdiZj82sj2IhRZcyrN
2wimb8DozQ3OCBYT4RBy0Q==
`protect END_PROTECTED
