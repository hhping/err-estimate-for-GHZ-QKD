`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N8ajQP0YCEall6q4ffVXqhagBjnQpjaHl8wjY3HEC5w5h7RVZBInX6TeHZzavqoj
iXg6uvNYiISphimzM8bdTSB6ik2ghO8LQHdAl1e7NG7ghNkFHeX2nHlmeDbr0jE0
ZfCKrivGnzMOYcXk6mz+Tf0lWx0TiGq5fRb0ThyPiXwY66PsUqqaZCc1rfbWPg0P
VFGqHOwzHbeYVQgI1P6W81wnnDJHjSLNf55eQvaEtBX/o/VtDpc4V5OQJKcvR4tL
C8lbg11W5PymMzzivj5GDjv0MxDPJ+lbFjn/0kvRpb9CModKAzoyyhCIZREx87h7
LGm+/rgjjNkMosU42qe14wfrSsW43dPNPWULQcyWofuGhKyuPxjmYOq26e1rfVpW
LWz1inZzQr/v51joDpZek0gveNBC2USYYxzsvhimhw9ykT+dWYzYF9yp0a5LTACo
Owgd5+RQgtYwDyAn9c5sWve38J8QlaGmuFH6oUMJRxk1adUPxo/quXteRmQ+1gNE
Y2HJKQXLn3sbPdGIC8/+YUKA9y1mZ5GC7R1XF+VIVpLk/9cBcXFAqE//omIQHSmN
1yYvxBOU2pnPlKfAbdRxLuPkdw/0wHd5ZMsAdSp4yCPn6ynPgTTSlVCsjFqw4S0M
OQSiPBjFBE4IwFoToE+FofRbxQVkW1hak8pdbe8zOF+iT3e7Nwu91lig3c8KMHsc
+6xuR8IFoxVrMtpfNPXIrBgZ8LFRgyZJuYNKygnIfT64YzrOKCrzMVuRn1PLApgi
F3k3YxJQhmdXrA/jg5/02CVVeudIRfKiLAVzjn/HjP4=
`protect END_PROTECTED
