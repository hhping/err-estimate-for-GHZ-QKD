`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yZALoGDY7QfdjMdBwOG0TyLt0rt2MK7qmBSOo5U0vIIDvyy7JK1TY96XUd/yBkYL
nsYx9Q8iEqa5aJrTX0olaRbygAdCm+g65HXLviUFC5wend/efOeWDuUUQcp8QG08
Arxm9GuQPYzz+Sigzwz0lYSLqP1nm9crKRRXXQi1uBvNkV0bxZW0WaNhU8A9REAq
e9Ot0UZZGeggMcNMSNxucQklwfUi9xVWdLBQXWmEcaQl9YVKF7wTJzqb9NAxVOne
149H8rxjz5LuPvnCpjojnSmdA1PozDTsy8tFcXc2XLe7mwMQ938RfkvVBQESgw0O
1V0EstvvRWIe3hYHDwoHAhN/oQeUW+34kDDrKFvZGQo7L7noA9eSrOYnb+5M2bbM
kFYSQMo6uEy/QSsTFcNarta4qej5PpRCB8pyDJ3WXe0OKyzfQk2a0NSVMpXk4Gce
jNf/eUnJl5yM1bPVxgyxWiMLqXHVOO4AchIsWvQzWRFrsPDk1mmbhJ3mrvrrsIzN
UcYb/OIOio5ob+B7LRadQOLDCAFTmpOWXwgZ1ytPDIK9xh7DD+E40RkTjqkDTDmg
`protect END_PROTECTED
