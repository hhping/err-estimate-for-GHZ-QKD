`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UFTxsWvPjjDFNCWugB7ktTCwJPRewwDnhMB3PdJER4aJhAET6LXKFayfK/m5JD0C
wwnhpSZ8ggLYNdz577GoU7f/gfoTiHq1adSKM6FJB4ssW1j2X2H3Dgiz0b8Cw5du
FEBal149+yW03ntCykuEcWMh25ZXHmSnNGslDfZQJR6W1THxakcgOGAgDvvu1rmf
0fhHnFUTa8iINP9jh34VHh8mLSlliM2elCtMMOELwr34nuVt2FknJoMwRMT87oU6
P/JwS48kBVHZbshQh2D7CPKl/Z4auQ0fDvgwdcynk+EuC8FG0iKQ+9rLY2rv7bXO
NuWj5Gb6PO5clQ97QCbWDg/fIFyeYvMGNU2SQOqYE/c/8thPGk3ixHTH+rhE4ehX
Wz3cQEimjmekhfIrFSx5daJko+6hTFAsVcWmuAZDkCbW3aX9OT8/xG2IgjYbDen6
oWoEaZS6AIKlzyW5VqKWm7Kx+7boFdOQhNBQRczTig5Q4Wt1EazwFuM/tLoaM29A
wjjHc6iUcAYyGoLWrr6vwOfIrAp4AchIm/88aDWoGTE4HwUgqG9bJdsZhfVETZY4
aYXLcX7+uWeNN6A7JKO34DcJdjpOF6R4tJmEERr5sm0M38rtOWWajzuVCIFeZQF/
RTlMwh5KDDS5avqyIGhE0cOyglgziJ/Lb+d7P9HSl/U4cyrGUpiYA0JHu5R0MrFl
ioO1XvDZBwu8Yv5ohtct8ClQvvdSHPaxFa6Ag83q8WSS5TvbbeffPiTKOUhN1mhD
QlqkGo9cRPzmSUrrUIJniDVZyQ1QJQuHLlbWWCqk+7zSitMn90VOV8AEu9Mnreo4
YqMclNAnjDoLjKTl9hCtKrxzj7QivrKWip7pG82q7jEXiGIEw10t35GmBV94KVZq
VoeWeBH8YNRVtZXNtYE4U9z76I1xn9glaGIPV1aszsxR4yxNDZGnB/rVq6gxEp04
2IqwiIqlUJZZCOOvj2JmAkFMGAk2NsikzQ0EyEFbiTpquZo93lBKko10n2oFhgq9
u6v0X2V8Qgx5FuhSCFUqbGm5vjoAft4oWqYWg4bLA7FC+vX+y+hKvXdwffnVQLKv
LbYwIzTPKvLFF+DEsL+34Cf5LKk1RQvAmEdXtSVuCHNqn75Ut1BRnsx0bJRNUfU2
RIMDnZ+FpZ+iQ8rp/RbRpW0XiDbvlqphYLCQa8sx8FdnqBtx1U2PIUwQYnY0j6+a
LboSl3wjZy/BG9nNWQHnWhHATd9PkEYm8gZihyIJZdpB5VsGBmKMzr/ekIgA03HD
`protect END_PROTECTED
