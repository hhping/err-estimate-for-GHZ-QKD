`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CNNKSclWrG3op48YxeZoM+x04ApShI2cnmvQhVyxmAWHONs1YLe1HMjRQ0P/fffy
3K1dkT4A9N0xiapA8Y8krhgKhxjBZeO/fWYM8Zm85xCxIo7IUwEmmjTJ7GNo4E6r
5fOOBad+O2x0nDB0bwp24WsU+Z+myYaaT9d9QykBQnDGTKeUYcioPaV6AKKxLkIr
XO07SAwkOjPveIQkhJE6e8zfvT26aNYWAQXvZhCj6iIEHv4cnvA3zE7mQXgBqPRD
YMeB9VovBOn2rH0pmJ7O3kZ9uua9XKXyJrR8wVGYPGOaKcyfj7KyEr8MK4RiRgje
po6TFDJyEr6oHxfwgkKoDnQYXTMLBAmqeodJLU5LUWF1JsJOGIO7zmTqFf+Xg0GL
rT/Funu9zaQCpsXM8FKgmnb9kYFC4WNYB4f3+zrPfNdjkb3rlX8WwHFzN8LNKP7b
FQtGd3tLDa1Td1LLshcO4tyq+7YD8tuB41dtYqv6hBrmF8lIKE/Ym1nA2A/BG6ir
aA6RN/ELWGJsavUHAA+OXGLhhXhWbcaOPorlaMiRCzIuhL+dZnpCFwz5FoyJHJgd
0/ldHSxtJbEKSaWl6+sOnr7KpWDxzcjbomEobPExGpiq8C0jXode8gQGXeDQ6kmm
WRtAT+G9evKT5tuWX1b02YPht9Xe34dd2WA6jc5OlaA7r6E9mcbsnIxhXowK1iGE
YYbQSl14vVOO+lmGnuNdCyjrh0qxHHjUSQGAfu7ajxqFbkA3LNGeJffB6teIXFDJ
CC9CuBlVKErmxkHXhCg4rUiS6t7AquDfLZiccrBDdh0jAXiVVJQx+fi/LARt9WFL
5IAE4rFMNLuNmJkAUusw9AU4phsBxosjkh6lYNEGb6aBuK5vKcHaVL5vo+ZReiX4
QKUbbPyt2M4BCXq4diH7Heb1z5SmDfAd/rBn30igqT7Or6nZszMbe4Tj27vfRpNN
OGkKG5h5pQyJaEXDdU5RLHDXNu4PDOycKWh2FrvHwCos184uqH22JAncIH9JxByA
XtICZWU0GCd+wabC7o7LNFTpB6q5xXl39FtCu5plzjrjtXPuKFgYIn0vp7bCEWCV
RMPOXpC16HSUdylxugA0F9DjB11hnpYr63sYcoEeRg7G34DAU7GUj1ge3PV+pgqj
hWYVOpyo35ENQVJTSqNkG294lW9StI0yHGYpF37eWybgu1zFEPMm1KqeTPIZMAka
nY4lughj5kbJzHNF5ht1fGpg8p6u+O+EEtKAxqXr1/Gkg6AkXfZg2HMAFGA7vI/v
5C8l1mhQvDK9hkfYCm0nJujOtRmM+Csh15Yehxf86oA4kf18UwW9o77FsbO6qb4T
3I86TeMHiah/5caYo1ts+MDFh878FN9TNcksEdg84FB1Ts9rd5fRopYtRa8h3c7l
Y6IBm/1ctrZ+9x/TBl6ku90HptbOyNnYdTiUwBcCJyYEOAYgogn4bMZhfF/yFPE3
UE3sUShYVrayzf7Nqx1c+Zt08r0gIJymnYSLz5xwjaTEsfvL2G9OM4vYWdXMCftw
t9eCmVkWX0bKuaz3PpLldKWUGrgFuyVi0kNuTaUBqmT2KUw/r2TX+wW6pksJRdUO
wwQnO6f9mSMnKMUzn0w9527UTIqPiCKUwR9f3emxEsOXd4RItroEMvUVapVIClIF
KT0xmuCa3hZIwO4HVg7aASNh9nFXCqZbWKPccmvgNi7KmoVhp9U5PxRQ4R8nZ9r5
pAVAIBoMD/UhpttPh08TTN2UU7zUOf8Lu6uY93N1xo0=
`protect END_PROTECTED
