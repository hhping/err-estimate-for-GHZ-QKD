`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NraYaaGcbdPvDfPtpzLecZdzTjcvq62OgPQdYMW9EVWHPzzbs0JaphvP9E2gQJIW
PU/iKWl8EXvw99n2OAhmoJPzJGPXQZ8APzUFvHpDMpIQ5DDhjUWzv9VObcN4XcCE
Bqdm67oW6DHiBqg+aT6HT42TG3McllttZ9vy4xrnjgi9n7/Xz5IY8TpnW2MGHKQG
dEqo9Jrxf+2V6Qu9DuOiZ+xdM3FFhIA6jZauNNeW4OfrNrvToVfYwLDTJF+wwWSc
cahhe3e/QIl2Zz7Tav5TbBFBXEl2xtjDR2KCxGOwJ/zmlJdG01Tve0ieyMB6Rcie
IptXtukCBNtxwlJqMDHbgbRJfJHu7y4VCCNCCScmhJUWKAEAHjZSedLD+o2by8Aq
6a0qlA4kjN1NpuOlxEh987ZQlLdqTFl/P29gjoNBSQNNbDcAboqSzyswgiPW1jru
/Epvltqpjb10vtUTBOfb00UlKXAIf8miuQ9KxSWIDBjltVr9/48Kd/W29TceTZUJ
vvWPZJw0r4H8BH0GhyvsrJNqmI9G/9bdv0t/NXD/oE3aRLEPY13RPKQQzaQ6vMFR
`protect END_PROTECTED
