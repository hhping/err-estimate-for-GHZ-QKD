`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bSrOJnMIs9aUaa8bY9vKn+tQ+eOwpYCujin0DK64kaJTPyn72b0mqIRVxoqLeH6x
S/XXuocGxgcnHP5bpsqNRwnczxO7CakQk7hMaxc1rVt6yyn82ykAtTN5gY8qa5d1
e7t+dWbq78yoiYItSIOmeP5Uqke4ZFoLGIB1ivULyy8Nsl/qYu6eYmVOCr3Y8P1c
H/DuH9EXUDqP2KEymNlJRtbiYtYLnhdCvrJEt/bjWZRiuygXtVNY33R2F3gt7N3Q
gLCrcvLKizLYps7hP2qko9fD2O+rxW78yvW/4wO737LjnOPAWjf5TJYvRWbsTCg5
k7FPUhmfPLZomqbNFSodefg8hVqEcwlHE27nOgBlTwPHMR8ILEASAxblEbsamwMx
CtgjhQbVJ49qghwKxKUHweI1l306si+qsMy8xmY7SDq47/9iIfUFwerZPqK8IQ+d
ZAmDTpedC8PxdTqPn5s+5p5UIUh3WEAhYt/OhOOfGVfT9d3KcHjNxPV4kP6fHKT/
aC5f+ibJPhkzMfaVQaHLZsOgVOyhI8ntPmdQ4+B7yHg42Vul5cAL5SgMDWYPMQ+6
naWgKRpvgGr9QtoJMb0HFkoh1HusInTAVPjIk4ceZs50nptbBCyYUf98/X9+vQye
/cp6ukdJ2z6IRFjNsfpvGunni6y21yIXrV/9Xtdz6MQXFfUkq8NXNzTG2r6yTm6v
bfOaGuoO/y7M3JItwkm3cYxFO0EfJM0qwhJ4yHmirFWOh+kiLpXeyqPi2F2jY44g
9K2kpMXFzkRME/83EWDsPJyzuZFBNFRL+mcgy5FMgYMQ5C/gjZNaew0XT+7jKCHw
`protect END_PROTECTED
