`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/edxfOfpSrvYgFBqHIuXvbO4A1HxpZXNyN2lHVRmK4RghEBK0bNrykgk5PTyRX5F
jer6rXfZbz0kzR1PEswqzr/KcJUWpOmbIrz7yKEBvjKutOdnrDv8yBliVruMLYJC
7NdvpSkhu27ojTgzBd/QYa/Egoga2ELWYGp1MzeZV61sI6w25otA/6GUsdO7rIeZ
g5s4tDCn5sFiQId7a+ZmKH0TbtY1mSIRAD6hemEILvbD0bN8ljnh2ae+dc7g8xLV
FoDu780zYehQ+gPK9JsO+kqBea2dPmKmINyYYEjNn0uncI8hVASGwpsAIVlk2xcy
xgStzHC000/rM/s3DPWJbWGXWcSfkqbACSYjyXb7hx8igMRIsanbrEzq8bjGQIU3
Js4Tl19owIXgHqRVBmX7eYexgCWMDMcozSGb9qXveVghnKJ2iCCkYHEqKc8UaW+T
e4cPTiPtbKLgXgIJvTel0OJEGpsWmyZktj/vzfe/uceKpZX1K5hRnU8KSp/YHhRW
RfSfxyiPkiHdKDbAqqcaVCtmbiaHuSKkKsCG37XDNUE9+AAJiEDU7chFrn5kUIlw
0ESzbAE1aEHTLJLdHrcvtUqQobW8DRzLKHMzMHLFEkp/8UER0XF2n1TxXgqfvcqH
YKLdazOX6zZt9ueC4fC3oujqklU/B1EpKYv8TmimWKWtwxBNcp/+5dKehxZCfQ3U
XntlTyfE7QTj2Q5CEEMj6Pt1Dok5/W1fYRs3Jzk4rqlUCpKS8CNBoVK1WtpKwdE1
uFREGStovJFt6BUJbkm3NnKIOf1YGpshjOFs+6UtciyiV3a2CV7spv/0lOoAB+37
VHtTTl8cZtSila4MpTisxIHfv0+bZ0a4vdCf1AMriiCtH05tgbaBB2U2M3fMmZ15
vLXiy2DSyDhn0qYSan4TmCKb6i7BYQ99k9VSB0U0NPe7VxYajToSagOKooG7osjn
z/51gW/+yTMA0DVJkcfDVtmPkG+i0CYRWyY1RBix+iOQFKvUpvvgZtNMc6l9T4F9
idsHnUTx6V9UDrm1xT9B1U5SWVtaMbf5sLi3SG/kQ2qYgyTreytWZl3AcAeZIvEX
qpUT8XYcW9PzABJ700P4yu8Gm3q0grguF6qOSvN9L+q9s1e4IQz5CgidvlhLq5pE
iAgiS2h/rutE1C4DNp+/GKmFMLqH0DJnEMXzGO8bAG/s+P5jcZASqqK08/2AF1cg
Q1DblK93UMvjr98d2l9nzAPYhA779x7RwZpYygYWRRm1MwGZ+m0W/7YNQp5T2dDn
K4/r5shWdPp99/O6Bbw1dkAnj8t3WVXJINDz6jBBuapwXIQizWlmKySEsc4QjS6E
fzk/wjL4wByDbVlMN47Ua7zFjXzB4et1mXritPwnFgAqK9+fNbfWRpKCn/nqE35u
llf5yaDw5Z2cTipOQzY55BIa1rlfVy86uW3L6Lp1Q+CrDDrf6Xg4mYA//XsA8X36
TDxFbvYHEGYA/OHwUfsfuxzRPRj0ztyIDL2U/PbkSZ4zhVn2OQK+YXyDEbkSM6oy
2QpH9N1MSJ3yIACtdJL2iqW866QSibvDCCGhI5566XZYd7EPQKmMRoyR2ID6Uhha
xP7DfTUWOa0GjRVEbOyGZ+met/l89OWefz+CIlOkzcmeaTF3RTMx9khdtSo0WXtw
zuI417ktQ9mF7EiFGcFlm8QJvZHYhuT9mOH5WZMY594osg8LG9b5smKNhVtDsIDA
7+DhMRk+xWse1PSqmVyupJIoBRvGWDRnNDE4d/+od1XTwTzRCZuzYh1xmslHdNJ3
jM9iTmsjILLz+cBEYXEci9QtqHYl4p9RA8dKwiI83oL36N6fTxq41kuNdznJ29lS
vrBDI4WrgP5RpVqjMwbM0ar5rxrChzmGtnP0C+OIwBpv9L2OC10ckllzzc35bcmZ
kP+wZL14PfFI1/AfOCuzJ+ZXzHYkcs2nHiJSAZhX12rz51MiVVK9mVD4oFeX3Nrx
iHnAqlGmLOEwRTlIr0f6F3G+hs/E3xMvGVeyy+ex+BhUBntAwi0RsPm0p7ToMnYz
R11zewtRxJFPbGCkmlyOEJNl1yEusIvvUbkJZi9LSVfhJWuub5CxeySkYqfEq2iL
D1tpRE7UIB5wKOQkhqbWihWXyvCuma9TLhUhrZ1Lhqo582SqmG0lT3Zw3IW2J+Jh
JPosXEgB9fqzCXhl/vTIccliuFceqLAfsSjFUMn5oVrDaW2f4QUyWUcp5V6c8KOV
Cp7yXI+W6TLM+53LdT0Vi3Yf1yjlKY1C4xKHZ6J5byNZKDIYvY7OzKKNPaGP2gw7
aFjDv6GR2Km+1NpBGEYDU6D85n1BpN5tWc456avyRmzab/M3uQ/jAeZBiKF8bX7I
C7U14O1nq4B1HwP1MLkq+lzEcGxlaKLwWjK+V2lgF1sHU71jO+KEcPjtaSaGuj4u
/x99ZDRMDkJh1Iaa09o7KX2Hr9TiY4O6d9j0GJRGqMEYrT9u0aDA/VIFvGw6N0CN
M5peKEemhHHZSDZafsikEQ9GlNyZhLaTsmnsAVaY0sljnHAbFxX0QFNxuApjt6EZ
lCatGabx8RfUc5vu40sodxYpz3gY+vgTFli7iaZjnGHwKq9rz0gTcnhhO2EJg679
Hrja9D4674S5wHZKj/DWLdCegLbW3gXojsDQGkhOq8l8RtHpg/aLmqafgekterD0
+CFZULUheO0i300iz88GI12soC8irgKRGjK3a49e0sC2ov//6+NjX1+2Rvkct0BT
752rd0DWny09yQSldKVo0YFdcBMrw73kyTVPw779jBey7cGVsrgJxeHh5hjCBjIT
gSiDCjVqtuxsiouZofPf06xECIG8sRayfW6snhK0UF6xrMi8X9ZL/1lSrhxWs5Kt
z8CGZOiLFj5ePhLHBZMJMQ==
`protect END_PROTECTED
