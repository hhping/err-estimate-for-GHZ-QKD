`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/7z4jCbyIQWrholihHvjegcCtjK8soq8pmKTxPNnDoawm36kBr6Rd61YeMwrorUX
RGfP4AOpjoVgvDttHTuJgZMOvZdqO6lz3AvbJF25Y+hfCLWfC9YPkdkmTM1xqt6i
Bke2gjR0u+dcqrrYmByt6isoXfCmhEn3at6mMj3DVyUH4pAoJvRKRVLwCqvytlyf
EGWE79SoDmwyLRN5U4m7mMFJTyxdo7LiNqqVG4epI9qFRyH+O9yXvwmk+Qk3zWMI
ihlTOGwkQqiMn5lr0C6nPdrWzO32arqkUjejfImRZ2J/cj0OGTKErBx+ZZdNgIJi
n6nSANGO+ec4hBZ3xEXn4TDrOAwfIaPn60leV/SGo9GnanFnvYzZOqdmCrQbcaj0
95+3tbaaBeaKN+pHd6PmcopcOvJn7qtb4FR6xNlZjdrekauPCTvApoiayGj6oV9a
sS5nsTY5phxUHdqXblCLJ9XA43sWc8h7wkPLxJWn4nGrlWS3KtBYFLJSshD2zDjr
lTQNqDdYbF2Aol6RB9E8qTA9sCzSKjBV9OxhQXy5wCrLsftveXslskSz28E9juMn
`protect END_PROTECTED
