`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jDfmVXjhu5185fYE0vFkCg/gGeVcnDqrB1jRDc3FOopwheDrStRXUQdy7uprXyg5
xdlHnXjgy9ge0W8f384TMrdwB2sEX5vLI4ScNOMt5q4rB1EZUhVvZ1D3L5RxCCG7
OJYXxPC0L0v5/cFDpAPnt2IA6mhREw2+vH7p2L50U2kPavyh/mct2jZr7Dr577jU
hwPtPnLI94IHIj3YxYFMMnA1bcx7POprDIVeM/RJZKoPFlb3a5NWmLhpBaA1l8kB
zvZJLMjFsixA/7MJoNkHQQDypJfVzV56v+TbDqD6TJeP5G1rp2pDrvwfaQYx2S1H
ufMGKY+Jv+TwIAl3+R55Bsx4gcWvYoK9l2RFekI7FOEGfjjSaTSwzrjeujYpygEY
eL6WL38LN6dh7n9ErGY8sFUV6SqLPA+uylczugAv5g/V9WnpjNCHnbkHjAONPv1M
za+NCiXrpmhO8bfigq7AXuDiBEjo/2Sk939GkIGEujfvsq/DPz92eywUIjHSqp6W
8PNSG5DYOMkl55HawwDDV2cH4QuUKHUYS7SLYjhhTRQ2SL2s+xjnnSWZFXBq0/L5
BKXWQ4lUSQBfcWv9qXl0uZKtYDqIpfq+8weRmwfpIU51TVThWAttxE6/89cpCkuf
gHDRypuVREAWiazxOVhCmTrXKvkVVmqUrUnb8+ZqcSkxwjizJONg2FE65IKvLseR
EeEBR9x4qxlpUD5/DWJIWRt19E8D2+am8CI6Jhg9pLKUb7H1vcNx7Ky9nQo3SrWA
ruFEYoNzOB/oGs2YlRWwhvjRodvBLOkt4S+Dm1boQcwT9xXM7ZdsmaXBp4l1LOev
j+kJcKdCIMpJUu0kUmYz92+NMfyn7IT0YaShPz/9N6tlRpxooj6Hkpu8qCP3YPg3
alFGxaNOhjupkAOiTiQ809KiyVqot1OhZA1EO1nlu8iJRvMxYoNMatEWUr+9Wo5K
O3rt2Trbnv92i8ZPc7PR8qCXOeJqrzIG849fidSm49Kc3byNYHYzei1fwhzrSKBg
d6D41wfgA1MFaWoAOsZljvZ9Bma3Z+bcuE7GKtH/xwKX5WHueHvN2ZwP7pbIDi97
6XKSVgAYxU9RBNblPA9NR/9YEVjdKp0RRyXBdwR8/oV/LmdTbobe7GKfig/pyIRs
ejxPRa/DhXwtDjmeQoxmGNP1So0RUBu/TaBfJmOSk4RtUywrp4YRXmRqBHgC5POI
W9xqeDHNhp+GljBbIRbKFOQOQu16iu2SCbitnoOAxoSp87tohliGK5gdAYYWU9W1
hFdk7YaGV59SkYNJ2cxZjOkGV5NWJqsz6lhs/VMmBkw=
`protect END_PROTECTED
