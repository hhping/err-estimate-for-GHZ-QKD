`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0i9rAHI0wATy3fZJwZiR0iRNfMlnSECLOB5afD+TQ/41HBjv4fxlN+xUg6N+EAUU
HJYMKc+klJ01+dV89W1q0PWyk6UyPwjVLPICRVjAsKAKBHw0kZryymn8ORpfq2av
Gkz2chZ4KRJ6g8Wiq7qOEkvfLnWRK6CYt78jf4d0lWvI3KSyF3GYI60OZgHSaUCO
8otFQxsH6Yelkn5a7f74GVQY1steCugUNbgqjpv0ecOgTMEOwHmI4Fqo0Lh3Rv8f
wlU8QNTvf2TS8MIwLWBh1RApqPfFrKVOqvk0ZF6r4HYjy1U3yguJpOELPNvedEKk
ReSaABWh8KS7p34CLw++gLj/03IQ487ygypVKnBZizoYdvOTuruWFxGwZ4PJaN+a
ImvfmBqrwBOpv9nnH+qZFhaxK5YkWdH0VrDi3zAV9l8Z5QkHshNSpRmwNag8WRFu
4y14fZKbJunbmIdhP4socZID2Rso1xl2ZrsKNks5ckiHRFAGJs27Xn32v5gLrMCG
LDj1vfSrsxorN3Ub9+K2WacwvdusNNmmlAJLJNp9lKu1Ho6Bk+4wwqqS9yWg9w0r
hNsZ5Pt+oapydLiIe7uMw9u14j+85npCFlZbevouKhBznlPmQfJ1UM0lBtuL8JhS
99HW67peD1wEKcYX2Qg842xHCVRGdjJpgLLNE6p0MAXQRKFdwUKDnc84uczwFkV+
OwSaa5igSnyxeQBlzOdrrPC7oAu++mBac5XW9JeUC1Sbf4rsSm0JPAXOetuAD6LV
EE0XLcN/iEAMX/E0pEebEHtnZGZhThFJDAP0iNlj2Et9PnPtlcxDLGlTLDV52Fqx
IzD49c8W4Faq955BLKweNyeKaIh6jYckQna8zue9cLFWEqmYZeMAAcUD+VRRtiGM
8kjy96IDw/poCKd0s6590cYqOilnsYvBe2sewGprm6rXmqU/v83ZlrCI7aBwMayH
1tePwxiRNM3bG86pD1H4I5UdckyoSAvBuBY7Kevx5ugsXFiqyi/G0BUCf06o11/z
6GHBtW+jYos0HiOYT3zYCbEseDF9b3ySJp1fGiEh/zTLeCLqCh+ipc61vsmvAtHv
Yb8r8kOHZbUStY68qxr2/dU+aIn+fS5k8nye1U6s2KV2D+T8xO1BiCvkCBBZP+FF
OOgJtj0QQ3UB1ynVwW6QwPnVrU0eQSd3E6Mjq2tJEKmp0an8gC12KRkOHAEbKLkg
kefvRdbP83qpm4eDs6s4YTVbKHzTnjx0kiTQgxzLyVJbWA6zLYGOtiDf21dVRAmI
1TNa7YvFRZ3gU42LM8A+AstrcqL/2PptvEIShyeSRKiiuA2Xo9lDw7lVX3d3QG7A
9FaSixzKqx/4nigkIFktefKT2Nl8LLOkgrzlGOxfmFhRjjfyZHgrWUfgUuxJVlxK
60GfC0B4BsPl0XemgWjFWu/+jGLA0SvPlRgSTqYJWo5b/4D1wU2fBPksT1VO5cmD
HEbx3cw9croKiLaMeho3AEmpZP6Myp97i397/Tc68y+nTuUP5jq9lUTwf6+e9Qj7
Gl1YLb5MMsbi6woiRQwgo1Iu52eygNMPTasr9I/YOifHI6j/EPm4vibJJ+cBQLCH
2Z0DaFme49A1P3krK0vkHqGfMjKJHQjIcos6BIfx0n5m8xyNmjUPnY1xEATYMgR4
RyCNfYLDPRsb3+x+gWd1EddOvzK+0fnhThA8HeMqSCPzdcWQ58cQqeMKjGWmICAQ
GWWm3GOuM1dN68PH+aJyIyGsY9FPcVUk/ie7ulnDQA5+XKOmd9MktIrboFsF5V1Z
jcLzyASs8Rmvm8YoEp3OkIK+JpJp7r7qhD7gvGrSj5gNTNcoCm+f+BxWrmysgKmo
HHO571yj84xzFpYGcXoxxEgkX4Aux0pwNa/AAseyIWlbg1gl06gyevcjzMKcON+L
SrNqiZRKLPS+dsdhUdyKH4ptoDwRWgxFFoJ/5KXeBsZyM98CfRNFnadiILqLeMcS
E2DNDHiguX9eiyzeuSbVx3Q6q2FjZ7aAOx/Hy6wL/rwNURuK2a6au8/BJzx82kkt
n8fz/Qurd0r45MZxOhJvFMtxBUnxxeIdAEF8DRYLd87yvXxBwG6jIYUDpMbTFD4J
kq1VMgGjAsW3E9ZzocQ+gnfYS97qiWeZzUStElV3Wpw/1Jbvs+ule7TrEcs5GQCK
WitdhMTFLAbhfGkvb7xCBmWKYauDSP+ORn6XzD7CtdtjLF5ZLPrevv/nNgUjwnJi
`protect END_PROTECTED
