`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KZVBeV5NfkhxKoftqs97H5BeM1WwXIWw9/Ui3f79NeHM3/XeWGwvtNtiic81HaU9
QqZb3UlPLK3/bcp+cdu/7BaGo14IZMknBFUf0T2tob4ZIJ+nvJ3oNyJpM2JN7Aax
mv5NbPgJ2XhtjhJQtt30bFclKRgKPEZJWIHMO/fczlcqAa0xFzkfRR//3MHEnqk0
BuXVdVBf0SP0pM0Y6vxGNERQ2NXiQZBnPoTZtPZKiU1WGZK6Kuuh8NvUV9gr9FWW
OSOYTddRqiFiLSltDttpEqdkZawBV0v8p07rDpWiQc497yDYBO6k9/jbWxj0Us4k
dQAmaSVMpTRzatJz5dFCxzXzdlLPxe6j2+kkcDHr2SBq3WBsRFdm2OMrMey8cSbF
Ys3wYN486s1CVzC/B5+HXgxvUhLcrAt7Y8jwO02GRvyFMQUoU2qwWFKlfi1KWhYF
8z6+0A6NNmtH5SXZjW7xflqyUMjDWFcBpP6JNXfgItIzOKSprLmOpuAaRU1FAX6S
Okyaqy9Ls3DaLBFQn7kehXf8c34GkXlTQ/KA1sYxRfxv2jbKE9yf4k1Eysy0BwjR
7nIj5sh4pxMUuyIYF24lFNqZ3rr4xXhgdEjG84vHWA6MX9NqezS0vjobaGSsGk1F
2cHa6IkRoYIBZjT23O6aejZSMlfCbQwxMwa/2ICNd96GhKscqSrx0tkJCcMb44in
skyhsKsaL6wMypwe2TckD4ZoWa62K2jZ0IlL2uIHdHPnVSzTtN2Dsmvca/SBrQ4k
aZtXLrsZskOu8NBfhcJP6EC+0ox2VM9qPut46Qiun1hXpLMKDigjc2NlLcbpgR30
hBtkpMXkc2LMHIh9ZGLNRNPf+3eDxJ+u7czvts1jcQyTBcit7mr1kZpNzxqqdMAx
kBdHnyHI43icikG0SH0EYwUBZbIk8ng4sQfSfhOcx2DpM1WlZJPYhCYjzkfvhTl6
qAwY1OTVr0ev+OK+CFjjbm6iJ7n8WyJlkrdrUqTccEPOViFiyzbxgqMHoG78Cfio
/IUYL1/LedBh6gb1Mhy5oibjI9j+WVzW3Fa5+xguzEp6HdTO9/ScdpA15+NvXB6G
y8+kH0yM5BnxeWWIrJsuZWaq9dN+ezWw/mkg3WriuSN87BoDrd4/Ft33MPP8K1LB
M4/VpywzBkGTZMJiaWQ6ZFNgFks4GjfCgewWuMs4CEGjlw552PYf/iW0bJG0482c
Z4Pt8VaeQG42yrJEyOTYANtYGUVDn1du5Gc4Oe/BYzDeek7lzVQz/6URTwk4cyCq
+A6cGN379AzzhkJp8Navfh+V+oCusIRmfzEmyjm5Q7PiwrnJ01Ss+KDj2/vJ+a52
Ml7r/Tby51ExKEfOrWUHIps+/WEyDahid6/EeWL3eVZvbWJDaMBrI8Vr6cnr+ZHe
pJWvT3guLrP9ZJW2PXSmit8FJidbaoKLt5NWKeZ/NaP3oxh5cqxfUgHCCTztjJGU
RTmzPADt9FoGNwFet8wl/rTa81y2zpfEBOlg2iuAzzcaO7T8/bMcaY0QU/u5IV9A
d6W2OQTE5975DkwoCNZNVxvtCPpgqjCE86hAnCEzGh2zZStwrdCHPmo6azGub6jT
zpGWykR56Io/QWCq9ouEsU49zdjYVwuVFmJDlurRcIkdnquKSJCeluYrdAe/8/YF
Eh/rEJZgbeUmdHlDsukn4d7u45nNP55SIgaPvtNGfnWPV02zB9TZHCa4gWTZvCJv
pJZf7ECDlSeCZDWClScopNMykt/4ojqtCpMO5lonZ+OaewVgnoxQplx8eLt6TfbJ
4DeXQrNht4aVzD3HSLsmeYf3lbxMhJnYHWBNuQ6Y7nNFsmMFR3nsUFIOvP4siNbV
0jlZohXuWY4hjt6Znaj0Btb6cdke0WMwjJsnih6OCciMSBe92OyW07fHr3nfcqQT
X9lcS48dG2X0AHm2/uRz9w+JBMlwq28VHzPW68XuURE4g9fwJg82EyJHhhpwrz2W
vC8EXskxlRINL/zrcwL4G9V9zrydwJ9Yp9HP1SboRM4F0jPNJH5CnduNDONLoIXe
bPvtZU8gc3sV0pATKMaACDGDCl1MOvELH0iU2FfwlxSoBre93ZFOrLTyJKvHDQXa
zuAB2ynBfkW05t1xCRyAQA==
`protect END_PROTECTED
