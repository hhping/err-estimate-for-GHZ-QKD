`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UOfWKu1B2TKFy/AJbLZenTW8M7GABZklXlmuGCh7Q7EnwyFBNQ69DfTUCNEUz+S2
9D9BFfMIZxlvepuJcpNc8PrL4G8QKtKlsnfb+PA3pS5F0HP3hjPoFzuUhpQNIQQg
fRv5bpT7+Ob87tfAQ/BNtXAPgrfozTaGfW4NUbL+X4ZJ2VXd4aXtf/DoY2yzO3Yc
NulQn4gKYbUM9CXgxWXPmn7CGcvpckXpca1V9bLAZx/yfG9lNeVORAWgobmnwGHY
pqWJo+mkODTmGB+z+I2oAJMrJvbo7NrW9RwsuSIf/oCZS4v349PsV7oPTUm/fczK
DcxrpR2pz74j4eZ18XEuaMDq7vTvwgGlFdiNQFYfP4OWd+nmf5BuA6BOg4Tamwrk
vR2DI3qLkBLOrL9laqXwk3vGzLU1UI71KyqqnMx2L7cHHULwFMCmSFcUwS07pMu7
b9p/iwZ8UKmxeDZ2p4INT9Y3bRQGfWzQnm1BSehoFPSOjAr9t8JFMUHmJ0b3YQIG
aN0V6hvhDtfLZjemTL7thdwShjLEkJv2pG9n/uOKK5fdce+2t2AKF/I49ZBodLSN
mDKv4mZwDaH/9cQyTLAAjIQFwDu7uaPVfmfkkT1Lyk5zZjwyXZwTNPrWWHqGjHJ7
+FL8nFBpKaPUzn9+gLdQA+8sD17+oB7Sp5JMb+E3wXc01LIFTUkyUWaEe1QW434Q
xAF9Dl9KX3Y16fAPfPHO2m7rGDHrFt7Cp8j/21KHFFfxPFOy30ksNSK7T1V7vdxK
rg3VHqnd2qeUZNt/yaFdNZLy9YcsEdfZVfRJlqui+7kjBvEvrKefZcPj1eKcHqmD
jDCs/49RoalPg/5AqS8NVtn+85uGVFHgYawn3+mJErHeH9nkS6pwYJqfl+hRdo7z
G2n/KG3PiLAYIdoyVeiUkPpocTOoUfAHdqqyP7X62Bdm5Z/JvDz8O3OjqCUg1H/Q
/m6U5dvpLpfn6pb+fQ2+LlAieQoGKoVzvmPPwxGLm6hzU0Y2QMA29G7+RD4VVurT
fwb2LkQWSh5Rh9eLf4w02snFBnN5/ZOU/7pXz8XRFwyY0VDPiU37zeWtdYjWd30S
rth3d+o8TGe9qT6QIUM2lRm4zNRTV1B1X+8rfhVSGjq3t9Rh9D2+lruR/10owPEl
OJic9ycMtUmeLq+axYelUewYAvzQfV+nYaGJfX6eVGwVrN71BkXtdU35tyNVIqBf
u++a4SHjMyOzxECoEGsTlPe/X5iK2aRdi/+dk0NPqkKmt8VTwBoMNRxJw0whME5m
CIywE26hZ9/vFiKWJp0Gu6lNAxaz0XpwTTBLatpm1t5CLuuqGN8RHdMyFGGAuhh1
wEI9SeBOgG2pLhvHeG0k7wD5IOilm5GHg4dvjPAAjasj0LFX+CCjM/KikiMCKWU1
2r3mX4uues761/FE9jlL0PQAOTUrhCg9B6NfmCNSvVb0i0kFIEovY5xF3SieOOun
UzDZOA/bYjcUKkTiyek0L8I2KkVlLUb1slobBpKlxxlwEkzWFHPkRQlUSGVqebXH
CfRCVkndUPdwWZMlhQ+Y/DWX9K4GYgNoOYUz57kglXIwpiAxST2w1J6S7gPU993M
06Dfmo8VVxVEI3hP2MvkMsZB6tdVGtMIoFve02d5KNtdTRVbQBtTAvdaHdFG1ZTg
0DlrvK5GTvwuxG4ilETINM5AnuHZic7Dr4dC08kdu8CIOfeT2wKX9yV+Pk1np0qD
qK1yeFFplv9OiYSDmpr/l13uaflMAurB3oGZ0SZ4SXHGstdbfv9bbAoV6w96BHtj
9jvrjaZrUBLAufjGdDQPdvi9scG3F2okd87Z2wA9sewSxRZV7qbUALJXoyVaiA/8
9VH2ieWmVV6SUy0ar6jimyUTwn4sI0xElCoulRmwOPtlX2aDz2fYZ2mtWxpdj8wS
q2xWRwZFAgNfNFBcsF2AEHyjMUZ7U1hpeuWzovudpNHH3s63w1sLFzX0n+sjQRvi
qZLf7eH2RnES548EOEIRJLj3q+fwltEQyndrtUIUU8OmA92csD9VX2nYUk8/OEvM
uzqzUk4vwUUi11XzL4RllYPYepvharwrB67+rpqR3FjLIojR/Grezc09y434/5Js
EmZHwtrujxzvLzUKBhkiUoCOWiEuESMB4WZSAAFS6kSIBTEgI/Q48rPKcV+oKOp/
eeCLNQi+K+/rRxqoRr3iEyMQsq0TQaytp6Bu4zw1Y1ahXfeERd+C41qVbNd8Kv8Z
rjOhMjyD9kEp3dT5Cbpz4dCD35bLZOI+r9djGz2nxseKwbR+joVt41yvauvh9Qxj
0C4fsq8+E7CD08q4LpUK6Vnu9Y7qNyQpjqn7GmqFTSaVs6BqAvNgsPVZBoarYE9r
9TRm6gUmeU2iQ9JOYeHSlbzcKSmQU/kfpvAw+pwWvbXMKV9hayYTCIh7MqxKH8UV
6ffHjwBaY/Q0q8WkjWBueZ5Ka7C3nzkYrE/thUR14dn211QPSG9lhg/u9tUZh5Kq
+VaoIDRH4sPx3NnrLZaBXUKEMULoeuLidXvN5T/R2xZEycUetrHAlGGiFpspIPtu
5e3SVin9LHtGirgW9uD8Sh36IbC2eog1c98FFtHj43U7z/DHK88qZvaq6az1J+6u
Z/263R/2MUSlG2PGVEO0z2DdDau2YRZIWcRqzhrjaWiFyDboomPFcN5f1SMruquv
l+nKbjNpL2IZdcMig4IksiNR/iIRKGxzuisDoKs2rs4TEimHDgf8WYsuAMgbZCMT
HJopJclT/19NcygV6F06KINsOzmJkKjDN15VCiGJBENoRG+Z9wWeMyZF/bGsPkEG
lzekhOO+ahmzP5Y5MRjrAQtQ9WYQ94dFxIij1ROhQdbyftOYEoN492Zwk3GcYs12
ju/nE4AVvd8oZ0qUv0+a6AL1/TZhXMgdoqFtIcGghZLstCOaHfCDzCSXgy24eNlG
qbuTQH1K4og/dsGPiHXSJnaHTVZIWLAG9QE/7439bRF2Z/nzDVJOosmvvngzse/U
Uw8SODj42V1leS/4TMgmTZbVNVpRlESkq7QP8QCX3w7aMM5m/DjT66XD9lW3CNv2
YlHrSpA6P9zpP/KzoDjvUxH3KKEJFI9xJMZ94sEVdzRcpSYQR4ALj2MGdxYYMoQ7
HEFXYtn6P7fblJ2YSl52Y9UApkDDZ5xHL6GoUbaCYsjWw07Fv2OOx1zfz3kAeqn/
VhrK4OikRru2Y4bQuDcVRqqaZ58dah0yii/Y1Ji5dEJPIVKjy+FnhiMkaPW45IiF
QU3bwW4yJD2aNwCGiBKG2tU+fEueFPv5qqROVe53b9HevSx9ZAFAxd6b+e9V7AIw
bHe6T8kxsbG1Z0qDlKTZhLioE2ZE/cXhDTAh070cQRTRcrU6xgSdn4AqSRKsI+q7
CyqnI5x+O0FLNxPD79F+wZXG4tsukTresqg4sZls9P+6cBuZd/JwV6UVBywJpfZq
4vjZWkTN8fFYxSfaZ2iDmv3JwB29h+zG3buxk67UqAOK2lo7JcOIIVeWBYhquf1m
+lLR/ahaSwEkX3OzSTuIfy3igm6UCOt8a5FHgT3ReKXDYF6E/2ncVqh8FTxkXs4Y
rr0vbOC7wUyGinJolQicQIj8GUC2sO7PIETqdQOjHLo50Hx23JTVo54RH3u101hM
TMK6+TcOOin+elmSUP7r33r7R6Kw8Cr8ZA/u01cm8XBUcqcLli1u07Eq+BXZsBUW
rN5fQ0WJh5sWMftjHc6ycxrOtFzI1Tru4xNcuhDAT7m98/F2xbYWRGuf+fbNde2B
hqXdS71qPqI4G4ZoDBlLXvK30u1orUVzO1Cm+kuDfCtwdLpwYz0IhhFZ0vy/ogEa
fGM+VM+UgK6stMI4AvLFK83FxDKeHvGQsxTVVQ9SSR693/8HI8JYF+hcEPYyuMCM
L0AxNECD1nKaNqAPqd1hSWUVrK6KYDxdKZXnOsRTZHRouCqnWrCpR90Hzcr6eBtc
7gTgRVVfxQ97NoXo2/SLkejEdfOI++Xbz0qRRYgTS+tfE2mamYRUf0lcXK0O1hmB
5FfcqJrueIaMrJ/xra8UgCYPUMtid9comhlhhdVgXTdTva5JB+B7b1nAMSgMelLM
FRJq0gpyXJG4nxRpU+crt+DsUBsIEgrvMNrdbaatnJpTCH7JCZldrBNKs8tCH4NY
ID8WdAsxQ84V5FrB4wDbB0Vty/6UT+d4LxZGE21euygICSzcEQqJFJAqv8dI7FKe
2XIaLGwrhPkDphYZVZYDS/+9/378mrGrth7IRpZn5WuHCyVbstuWqN+HkZRaV7q2
Nbrigu/iY7KgqRRA/o2GsjC1/3LGzvDxIHQA/+nP9KMxutTrCEj35VRkhrQ2Q81b
oSDZw0FQLGPPQAxC7tTSRhly6bACW6gqffl/C/jQswNgpDFeg+k+AmzfKZrQMPZq
mhcEVkQWRvDueucqXnLXn2l2ahqewCHCufwHeb1/mRqeGmFp3Gkk14d5iui3+7Nz
1fO9BVE3U1kOp3E7FKzRYJlpwNHd72AT6bTP/ZI3Bci8pV6Uy/NNy30MKR7+fgne
K1mA9eljkKR0xG3B8B2wRsytlijt9zqL/yZvFe74Vk8GPxaNyhcZOl9O83yYNGVk
SINJA0Yea2NRF3ZraXEIqqk9OzlKC5+2trOi0n9BBJeuqD5npCeXmwOuqJEgdzz+
+5HECRQpp5AuYg+7buRvXpzQE7QqzU0M1Z53pQHQqJjtj8/DF2f4HeOSIfULsDy9
gcEZeC+2Z8yFMGm1gwMSrAaAkETRqFKFY4CU8YGwR2syVxm6a3+U44NC/260zFXf
EZJnVdBDNLLqkBoHyW038+XuN2Y6tmjwrVbCcFxqCZfqx6tCEJOQyshjE8ws+Mu9
tv3juHCogO59olETDGZ4tN+mm417mLCTXfEkbvZmfHV8Kz9t9k63tOflpzjkF62l
2ylPtsQerpwTchmV6uA/RxjtduqJdlpd+pYu0IYGVC/TGboN486Y7T6Lanpr7iua
P1fbZcmDqW9bAG/gksmx4p6HEtmRLwtMCk1CWS6zVoEOkt78/3mkkXlJrvozkd3v
cRtTPiXI1AbtUJ3hZuJ3ULy3zGYeu79HZW2YyFt+BOa/Whuae9c4gxwwJbmHz3V8
ZAMkIoV8voKJWmg5QkXQW4O1Stervw6LkKxWMFJX7No3TwKtvYlNB5tc92q4O+gQ
EIv4aXlUTUlpKBToOQA8f/MnFQ8D2Pb6xhzi5raZwCUjUjvEw3SzuCNsaEu3EFm5
ca/kTAIVeUt4ZoBb7m3FpdRRlmKlKtEy0UovUplK5fhATI9PlFuS3MKM1sEDLqIn
1F8Ew5hKXNm6k4YvriVVn1O9t2SJ1fIZ6ZNW936FRoBEFOt5TsYeXLTEiRbD7Bht
ZSZzkteJMyTll8Lbn0FmHhVMztQFpYkbomy3BUCK8EB/k9TIO+RnhF63QXIuLDWS
oD43eEOsLJvCF42vXKGa4K5JKfJCROpCG+6f8V5ycQGAUPR6+YxZNNaGuA7oniHH
YjmbBdPAUOb7VWy90CC+Rl0UzSo5SAIcR0PBrtW7hpM0goWVUwmyIAWQOuR+/cHY
MHtQ6AU1122D3JeoPL+DblSwl0yEEjiO8kWJbYCBacqqeThqBs/3WWz3BXoP03Jb
2fXwSe/FhYL2dMXPDHc/sDv2UQsKXYHRQzasvPAAgd2qwGMCdtkR7MDtGdq/zq88
6Jx4LdUgm8KHLFYK7m7xnkAaARUzxSTk3GPRF9UpCJAxIYZjTt70gmrTU04zRzgJ
6DfRQvI+wlyHoXUK6+i1YUddDItxjut/+wPwHpLr9PMb2xcLCublrB+THMEWSyf+
A5lPVWs3eUHcSetkeX2Mj0IpcwZEQazab3Am6B0LuiwupzPRfbwy+J2LQM3wgH6x
VvFS3LeuDJbuK9EUATCybs8QWxxAx8l5G4Mr7pSScg7ag8tB64SKdjexnyT+Sq2U
eRJNSQka9pXidHbc9XnwD2abhdB1HUQrTuS4RZxiuGvbxxOzGqHTkpR5Ej8lukin
XHk+TpQiu69D3EdRpSIoa41zKaaxRrJKCzJPQh+t+qyatyaKmr4HZ5ngIEaVVK/5
Ea7dUQJu9y7fwMHBEkNY/IK9xy5BsIsWVYDP4rpyPwimH/M3JFqBa+O5n/rkFxFf
X/w3u5ZQOFnI5uRY1czlVR+erIjcrY4ZRPDWETkhM2GoURBaEzLCg887tsAzavp5
JJ0vO/aOmUPIzubmXKippW65h9psEWO4os5Xc9/jF1vPLItx2JSfukOstXf0P+x8
rYIiaGuCa9fZhB2JoeiJ4kggd8VC1H22a2z/2fRJb8mWhEGfbI+T61CbaWDQgPtc
NH5lnWlP4nNNWcfxmf+r2dmBZ1ZroUY/eqhc5e7lx/zydFlGBVxSa1b4G1VyVWwy
z16VLd2tz/PP7N0PjtuS2xwJqkEzd7YxV0xEf/8ECK1txJp504zLn6LF75i84tA5
ybQ4cOErUJcxDJPobGBM992MQV7eMYjFAz840BKuXFsZUqqPKnMBWYtO0MI8lN6Q
2uQQ+GCSay8f0LWSM1Rlxgb5u4/lDVeXRwnqkZjtp4geoUBiLDZMf9580PsYNBcK
k6Iex/fwS/Ddov/qgHR4LoKiDZ65TApcnYP6ZXQHxceveCkxTLVt+qLAA6yzBkVT
SpLIqjjQTx87rSK/o6ZpeVDvbI6YhavhoScBjG/t9KTQVXucKVLd1SuLaCjWeFHA
6aOtGBYP2E/oVtlwHEp5jmBy3BFhaDk43t8yL4H4GVa8SWmPvvnscDwN1cF6clDp
0Br+aSo4S5Lo/AH7igG3sQQFS0bvRLquTlJHtETC8ZtBFFi6rIyQyaTRnBUtAmEl
tDlPfnA8bsTjKCVJZKsDZi3M7+/Cch8wt4/rClaHfemoHRIvJgc5oxLJ6O8I2bBZ
qq9Lk1QV3s3jXSNlc6HovY+q34PrPKPsWxAJj/TzsLGX/4C3BZK+SYlmTXacwVGG
0WEWlv7APCRvs5VpvKrbW5glXHlp6NHZJn3g+gAZC8aA54LXKFpB3tDsaUzo78xn
NVDdBTXJ2ntNYAhfi5zDh4mQ43TsjIN8mrDIm8LiwkX3x4lc3ZrRlLswQQwOryC5
xxt5BmNXxfytKxvFhFhIi/BoEkyXbqmMioVUCSt0MNCxJmSrW7RXei0j3okYO1X/
qUTkRCxn+Ldgfq7QyJNFr49igXT0GsEqdUwhz35eFqLz9v2Xe466tZMDLWsHxcXS
LhjURsSfS/hHfsKh9F3WBlg8FC4V9osnSmXJZ9XHvEQl4Si2j860eBlXLLmBEGsL
YwTh+aAB8VmDqAHJIc6jRhcayca6pRJrzA5xRW3aVdkkOBKvzlaO0S39JFyNLr5L
PvMc7M/L2JhVv4AQPdOyXZ5fXiIDEGHp5P4Y8GVdJGzM4CbDsZUU/zrlVFZ9wTUo
di6sPtZYgWlk6oY5guvsmdLnVvCsayhPvBE9v0QJK/2+YtKk91IVi/GJA43mzwc5
XCVSAE+d+y6cf79NHLAvZO9sdXHqPQE4b4p4bYWHtdEgs6d0HvT6zgmFfdCNBYBz
Zx+d76MfeYgeZ932p49P8DzGr7L6YTREptkcwUbyvtQvRdNv5VQP1zcOih9WBPkU
p3QwlpLHe13CezN2S5ePlVfUyU/FgIFXeZKOpWZ40wIScKdoXaeYahI8ZHrMc8Ce
Gjq9i0x7O9tQvMJubUx1Gt4aE1Si2jvpsjoMkh6212TfC42pVgP6ATM5LuFEJ9I2
ahVEHIDSyG9p57nNVq32+Ia47EQv6/D8gh5x1QaV6D87D6HDrMTE/nD/3phu6Jll
oKac/omibwlbeOX9dw7kdNVJO4G3el0RRn1m+JuwebQqZawxsAh+6HkJA5V+d/nw
U8xGCSSIUQi9liBEFfpzBfVytWwoC6O/wqzJUAfqchCrJMbICCmI8yPdH5Ou51xM
VKBr5/NGvR8AsDWT4EROqVyqp1cXeOi7VKjPj51Qxe7e7KQ2JXsbUnPMnYCpTOYK
HDFDolSJ6g4epWenlLXZ4NtNq6XD3Q0tmW5Glfg/Bvl2w6Yf5KTP3090ze66GWYG
MjETi0JYrciif9q8BaMFV3Z+BHgdlHpkZ7aEfB5/EzlSv9eK4Jgx7JiCke64d5ue
g1k12ZV8FQQHGp4FM7+GhSxlNrb6sqaGY2sa2uJl8Nr0YtiweBLlXtXY/4QsMAjc
hI5HsSiZ0HEzO4f5yvFVv2WqQl9cgUe7/cq9aNkORxccFH7pAIZaPdhZNSHz9tEg
zXbwUoOqkLUT4nvUKrEDZJRqP6QfFMTKhiMap58j5loPo5kgOmZF93YazTJmiN+e
Ff4TMTcpH6CUXKCWjbsvSW13xY/yQLkwNOOCrWTzBSNT+ZEQhGskZoIo3SYKawDQ
8US98uq4F0QMDogm/gqZwX5EHdLrDy8WR5mkUntgyOgUT/J8aAmqrAy2UnVRKXLi
AtY+6R2QgThKRQtRqK5hPzD+1nL2i8RbiLOrFUcZ83PmXSzeDFcjTi4VkMthmcYn
Xo9uOTEUid6lHr3M9vBedPYe7k/CbvgcH3H3fYluJdGCoY+s//58BaWmChb550SW
2sl2pDfv2Nm8GTA8V2Iy+js6JLxYRkGpwC9gl0Y8Vr6DJcttz0USMIR9lRt1aa1c
vhQamm6KfiCrfgWLQPssWwDEk24bKyHs7revQBBn6THAL/PCo9GhIoKwk3ch0EEk
0N9N+wh5apf5ROTvH+a6LB7+cMNks3UIcWFm0CITc5FxFYbQqtZUhw5oi/H2d+Xm
N959+Wp/jalvENyMc1nM12j8iaUvWi+4Ky2/Y4oWMJaXskT9RARoYcbeKFO0vUUU
tyPqVxrxhksUhDnTtsQBv/EIcL2jWidM91qzWjUU8Twg71+HvWhNcNr0lceDSbD0
b4djO3gfpr9YWzfZClo4CyzxNzBNQWV+VX7sO647RZ2/sCaD3cx5rTrLauMjo04B
jbIi5rEyOUDAJIk7OAKNpA==
`protect END_PROTECTED
