`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UdzGVkEqftv59PmRu3LZ28iabQ5zBcKWcNhBENArQkLs+AGIoa0eB9x6851jeu6H
0Qiho4H7CvypzCPS79CLZAKvTuV/kHQ3SftfrP+etHhogboRCbVh4csMgcUEhfLo
mWKqhPAsL1acndlrlsFJZGdgSw/l4JeGI4AssMLmanEOoQMLUox+F4jNobzMXhar
+CWBPiptPmsu4IiGFuPrbWv6DIorUz4GKL766ZO2KsVKBervTH70wf6eIdfbSufw
DTdpbHbu8YLtBc0J/s6szyH/MvcrBkj3lgCfTRc91LFe25B72YS3jR+k8U/l1IsB
5RCaPAgQMMSWjZphGVQQ/UifrER3HnLehtfbev+yza0PN/yopXG0CO1OPGWnkixL
b9I3JYLERsayoPpPZ9IdiCStXxW5KHH0Lfbq77ZVj1AJyN3FEAK9umEhfkXDFv5q
TVC+cb+sfzdx7yfmqJONlDbc/l5gH2tWvmCCMq8g5cQe2jQAmZjawOpFhJyuleSP
WIB5mXGKctJdJS2vmkHCp0R59pLR+44uk8JRloQTaxLcmOvsSEqQMrA6RMeDu5UH
M9kjMr3VVsQMdlC/KserPnlsB126Etff9C45Ex0QT+Anky2q8CcpZvy14+UsTt5m
R+VdfuXstmETyLWPD6CUcJDHysgN56yTJVAnkDQv06D1pE7isO5xrTQVvg6BEpGZ
cchhQ0eSQVR/zUKUey13TOB1O3WnEhp297KCljhpLY9KeiQaTm5drYIl8nmxdqR+
0y3mpjhqyQCSs7Qt5BwiHTtciPeDwGFchSYtIgwMVSWxQrekfzrfGhIMjTR9iIiZ
WCqz6O6WHJkgmUEG27g7jIBxA4fhWmaQdXA7c5C78gnxUWUQyfgm1cdVtonwuTRa
giXLh7gfr/+sb0eo+WJOBeUN8LtCWtL9A0fMZB/c76cor8wbfC7+Hi08zaIjD/wH
T0LUCBs+WDh0ZvIzR91WnTvKirnxBFnOcrZD4K7d94aaP9sFnE48fOzSbAlWzmsx
`protect END_PROTECTED
