`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uGWRow+Rx2KGA1El3MhJIekUTvuqdTJA2syoDZ5L8R0F+l1lUz7g7JvsxnUsK0oK
vjUGSQ5Nsggfu/r6nzawWivfuOADgVifi5Lc5OaPSUL5gbFmzJ9nkPB6LsQw6Nif
cIw0rqeGXmQh+DUezUBpK0GgAPQir6YMpQGFjXsV7u9FskB4wopB9rp8lYyjUI6v
B+fpTsfQZpjkCbTSmu6bX4TmFxao8oFowigpkdiIZ/bYEcT1BxwRtufZDNlUdT6O
TVv6r2cfnxIvvxPzGIYhleji0+UWSAd606TKPxPIbNthpXB/Wg+Ogzls30sK3y9B
0YQox3hOUoHroRztYsbflfOg01234upKEiWH25ppS4ikACyEmDmViHAU4/Hlaf2T
iETukqSLTLCp9RmeuJ/RjuD0tfZUxT/Cm0aHvC50pgZz4EnVenwDGZOzEfpYCLGW
5kwM/JzslWM6zEXEqa0sGe4Ad/clKkciIYgzMfDeJKOyaG/5oOKbtZ5Jwwr2pPZt
UUbq8gXh6VEDmYEr6hM3QdJiMUhl9hm4B+oTAXklVCxoOj8oMdTRlhuSFyS3Tzmn
IpGwaLIxql4tHj0Xb1PgV7bGICG4VMGOvGkDR+ZrFAARp6wzUC4W+taWTWtOr7Cc
3rjV58A+lUmmDzHgD6QLwkKPLfJ+CWGVVbfzjk6UiCYFJKgUpXnHudz5TPzekpgD
bZVQ9w2kzDqPZW0GwhryXUqoh4K0M56z/52XKdgaFxONUcORt0DBIad+4R2KMM5r
hrjUGt6l0otstWxz/l1frYxs3Dx+Upl2XZ/RnZnfA4vsRslSkqyfDgJqp1gLvN+e
oSJlXRaKLhv9NJT7zblrRRTtS032dIFCQ//7wrH7VKZPX2iAD8wdCAdyYK79xThn
BTf2DWrPPnyJMokoa+WsRdGpvsJutGpzdHoAowkHAGecFEAN8i0BVTPDuPR+lyek
ViEgcwi+i3Qefn8O88gCk1skFmS/7akz7oo7pPtDcxcCscGrE+okk3kRFRTC1374
rMZbGVDKFqju0QaE5Y3HsjY5BeP2/h1UnfkurkCqL5+zOOLBxEeGPt0NC9gwA2+F
q450JzP2ZIcsbpe/zeq8mgbBEvy37bnefr0MsawepRCYAWdBWLE2iAPaFITjVEAd
TwUDxPwna7j4fDLoW4Ga3FJwcIESq281FUFxDkTlpLn7CEaB2/xDZzB5MtgLL7gm
TrjomgzbAHyPZP83YA/raEonhOsZQWnlKSD2jR7qQgTvnSE4J+INfPmrIZwYthWQ
FzWcBhvLHJ7lK6uj/w1VN58pFnIYCVWVEbSfLtZiMAB01SRs8ib5AAgXBFpxLKWL
xv9/e1Cwaaryc2s61jm7IK6plXVPhSxcqhTzNayZnsrS/irnHVWCek0u+2KLKTcr
+Ur1bHXSWtA/2mdA6gBbnTjVDcZxGkWTl287RJulpidMLkxvqX+CbGQQD5mjCq2f
FJwm93AzkxiKxw0tU8X5NosNX0Gv8u8pNNImpTlKL7JTXTknFy/ipLHH+WB+NPLU
aMdoyH95bKzAZ1f/cz+61+YrNtemalypxazTWMt1VSlvzFsdIxHN0YSZwdhYB2Lj
hq+f+AqFGMckIjNMTete+DYBcmzV7JUEHGmUy6VS0EqQTF81+iLJ1tvi+M6tz20a
T1/8kZz4KRtRyK7v8WN30FQQw7jd6sqgFMK2r7P7daWlZjTHao5D/NO63ikz30jL
JTPKaAerGNppuemtphr3GcBWB8Lxe07CnDQA1uQRIcQCRzKhawyMOyZAguvcLhe5
0sPO959xm1+XcU7zlfaJdv43pu7Hxztb05UT0H2I5cawHN/MIOWFa41frWzKVj58
6Zq9NTm7l6kFL29hLs9iE5mwTNGPrz7g1v1tqL2JsZTX7ifOw9Dze+TEoIZWerCZ
+HWktuIfRMAFnTHn2EVfNIE0/3g/0hGGKHLOgVTVQ0J1CglaNLfjbqc8J74aJqDk
O3w7+TGYg+aq//iBCh4oyWdQQfNbp1Tv5OAPGVL6X4ecBSdPdvVzmUyWc74kUv3T
LRrtfbCicUFyktHvUAIrzTzYFU/MU12353tcQDBs8IiwkFZbTO58g/1f3YAlHh1d
X7eoMVYExX/ZSy6gmlWquSpZbr9ZHb38EVTTi8QemWZVkYbncOV1yTA95HCQcpvR
f294JJ8TjnloLkcmHwkJXgh4g2o6PFe/MKsc2EcRXkYSuAvKwteVaNgRajLZFEyF
rwg9wp6FfRcLk4Il+JtyfHf9yuIRxNxm66WipGxQgzJG2ZUGbTSk8X+5H/+nJZlY
1SdtdaqiXp4nSqXKa9FJQ2FvnXH4AndMHfo0nX2sqgrs85+g4mzNT8WSMcKvBZzK
1AWr3lo3BfVn/DwrznoDY8owWvHqb+4IPqZtdrFVTuhQX8R2XWC0W+AeYsrA9aO+
p0kxnYIqMTFDXth2owfDx6vjSIFmlMhR9uQImPlADT7U3EslhXOJJsedVrEFDd4z
GgCeFKhUeIxGPaENYxnhPB+OHjrLZAFEdLAhxYcrJ/4X3LH9xAKEv+KLD5Yz2QuP
HcR2mN2ZN3npkbsKT5/7q04QmBp1ZMnnHRc43Q79KvNnDdQVCAw7s1gq83TeK4ri
B/NJ1V1NIbvVnmbGSLGLBdZ92qidRVNnTnrIt/Cu7tSz4fqC8+uPyyvCOxHHMMNd
SvISZI5oPfTN8/gZBZAnZwKjZvGUhJRrbjIaAoCMEeXTJYZ/dZ4fVgsZf66QXSa2
Kehn9GfrHoMljCY/2SamNItZf0lN3z53/Tm5mGryUKSz+5q7um3ot6VqNSj6kjBy
Q70I57SguPHQSgs78tLSxB3lWxM906D9Z5mL9Cw4XjdOgyOgmMXSDpX5S3oN6TN8
6fL7ou4Z2qGswbTHPojpERsn15cIYqml+TTVaKdNjPFqro+sZB/WJ4MYdPOfZDo4
THTtihOfhApSRmwj4f858WzjgR9uMdMEqu/khwhHszVqzYqtu972gasSovZv6SjE
DYuCN3tNVyMwKagxKWRMxIWBpKQkJc2pOaau2fDRv669vmXrC1b4cQCYT8jGGsHa
jtMFIvhCS9Wfe2gOoSPi3Q==
`protect END_PROTECTED
