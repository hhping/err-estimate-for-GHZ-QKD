`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0mtv7omthDARNj0KclfPEvrIJj4foCfZeH+wofSsKBFkBW5iUYFxtX55P0m23yOD
rWXgD7xwm14RrEINJgo/acG6D8YiqsTUKr/vNaFacAgdJ3dtHezGjUwFY6zag4AA
icQTXGkFnoOUufcIST9FS9lm7txvP3AwRaFh48vbzBMQkp+7ry+BE1UtI36GYCUQ
FaKiTTNQmmrSq6sI55VHiPpdDA0FGTVw6shz6uVA3FA/CQThsGun3+TMAveTHxnO
NF3ki25zAel0xci5nlHE/F2vIcih4sd+LMZe4tTaAXPNG7qoi9tLF2DGUJQkDCHC
aO/pHqa6ELnMcef9t/Q2NI5tKO6JzBdO+DFgSL4oqhOmTzXbcnnfHu5aK35Y/hAO
xsdmi4sWkCAgp7OjZ/5wSTDGn7eFx9Hr682Sot/FDpIHBunIzwUQd9rv6ctUsrQN
zyuMY6mdj/JnyAe/8duSZjGDl8aPTCuTzSGLPAM3L6Xi8eRDDLGYe9JKO7gwug9s
UcFwAvEjMjV6hI+IOFEPHj344hiHAxw3slrhpsD4CYRIl1tJjqCnWM3L+SmRkxSq
9jUK25Q4lp35kqDgvG0eo9HMocvUGx6YcmngDzS3t0L4muAdPaqrUpP4HrW6UtWU
NFzmri/1jKBsMuMCF9cJSCskgqGesxCRlkgrpNexShY3gqqqBS81cJMSjgukQ8qD
+5rIq6tUp5g6eK98FM1eCXT8VYL1Lrvsp/tnIfc4S5OKg8spYIgPtQcFpeU5af92
Qm7WL/jYdTLfdWGDabRCA1npFQw9n8xOG+BNx1guZNXkXOhV+/a1z3pV19DWq+0K
7Y0Ca+249NVEBGVOEm8P7UoFmfT8HBot2Vmosncc4ijAeVQoFYt9gcQSNj2prw5m
GTppBTuSGfBBYf5IT/a6c9QGs1Fc77S13RSAFgUm5Bj4Z/qkgfD8AhisW/Q6RkcL
qWcjaccl8vVwPqUfPeUdkHpT8UHDgxUM+hLZLd63cGz0nXufU025qlmsaxBdQ0PP
QqMuwTc25VOd0ajeOGYjExzeBeNpSSIZl+Jm1+jwaxY=
`protect END_PROTECTED
