`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
feu5z4LX5DLuezMhbQDIuV8SKgUV4istRPk9MXuCS5OqazYCWCxRAPxdy6pSGf7r
g0GJQKZ7ifJkCOSejurLQRJ+f2FqY2LLk3v76igwWgbZZ23sp5qMGk/HtL30Je0f
gW5vbkBsVzhTjVnhJDNgSWr4DMb1ejp2ALI5FiU+jYAC5VfjpSE0JZcFit0L5ZOP
yr0BEIegtthl/ls2z3bMTNd6kpnYxIPrQSrlLIC3l4Yiqgigupnu8V+O128Nr+Rt
8fz4coU7MGpRnma6NYLDbMwp62iRT0odqspmolZ99coUzHdM3UunMCMhYa3wH9wI
4yPq0hG5ue1rGEHFeQ5PgD4JBooWo4EKeRVFAMlSzl4BQyxI033iWPsPczC6hSrn
mO/Xm5adlcsg073T8qtgSujRgtdJdcE1odpPaYpwcO9/Z6/i2mugdITon2rG4vCT
eqYreNVz1VurD9ehfgdwLAF7PjGRhfAOhke+sG57XEsYtUHbIYpSX+j8SEHgEc+N
juUcULI3rNSPJrtjiZSdLzCSlexPSJVpG10QMJTxNqyHfU525GZiqzJ5dKNPnY1R
NjfxcrbQHurhWmnAt+C+3C0fdRIeM46tkCtTsDovu6cqF9YnL4rvaaA6/yg5rxMJ
RtjXeVxPsYpKLM8kweRQpYS8uiDnZ00XIrkfWSPW+ZWa5ozJCiv7GISg7tyg2ldg
9N7osTz769d/baXxsXTIiQ==
`protect END_PROTECTED
