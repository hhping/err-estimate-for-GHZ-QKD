`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OPl4yqkDgEdUfM6mM6lsgC6NW1Kkdlrx2beNwmv9gNkVlXSy6So5VwSmTKIdS9en
T0AkDAXLcJVzF0F+yzqLLfefBnR7b8yFv5Gmu6n1BR26SlyqRn6bwXcY8gj1aamd
GIusoz9G1Xzf5Gmr6DUEHvJ6J4CSV7KmVd7anbsuMbhmm4XKpStlqgvzdnqzVVgW
Phsvwju6Z1My5dJhDFZ2dmvXv4iC8C3dVoaZORYlzxvtUIcl0HMERQ0dY09YwtO6
rEo+oHXZy7NrSuMUpowocdZCwmdqlLXhOD+Xzi+MBIM5jnjJDRWJSpLR8Pr1oP0b
6FYFGKwRuQMfojqBdhHQxlMfaRWNP2tWr4muwkU/gOS3/JUUx47ZfHlpDUn7MSFt
KusLHs87aJzOmvKqSpt2neShi3n0LM2xFXPm7Ck94iM3KWom7vGBb8vJFOf0AiCj
yhVbqzWqMzvBdsW0gvhlCIq15W8zvs1MtRDhUNQmDvyl09HjtPrJghdSm5cPOA79
AYC7MBU56vYUgqmzGJ+m/TazVQaj5XjYgek9Dy6FbiuaU2Sjs6ntUV5aAapJbc/r
NSzBlq8x47UVQNQaJgouNVBG/tPv3cQPe8ToMiDlgDbeKbXRYRYBs0wq4TwglH5h
7eW0LUGNgUcLaKQ30IuCI510nN21/meuSV98I8FMWbvMI3TCgGhchGvov/6cQQB9
WgDITzwzPGcNrU2v9OybzGNR7NLTRfqTIaFnMFZGqj7HFpyCqx75pU9/O6H6DV/H
36/7QRCZCy/ewqko2uCd8xQA/mb2f/gHkr/EQJ06xzMD+F71XFuzZIAMmK9cmQMi
vtM+tMRO+GTVyqgUPeI6P+JXvkCkGCbpSO/xXFLzxcgpCUQyyZOTMkhtPNs+/WCw
xqdXnI7bG3ftxkEhAJB2X5uhbNGyf72YP7jGUPMWXzzRNEn+/Amo4B8jjyCbfCO+
TduHhc3BZpmu8fP2YuC7rSpxeeyY7h2L2AGK3VM42tItrcRRp1RHicvf/at86svz
mpkfeFsaY1ymIJUd2HM9LXKoYjDMDByEHPWoVGk7bdXwVTOT90jeT76YsvihHeQY
tgKjQiChp+/Pioqa415cztSxYfkOWzjcqIK1yDzD3eBkxcbgjy2lUPU4uXkcTo2G
KAy0GDJxECSYfvorir2yzGrUw7GUUo8hFfp2sCzlhQGWlV0Wx8fXxZ0sUX82VXxi
IqcqqJtAUZ1eAbI/aPKzgvY5eVCV6aAuKlxLGyNIh92qUTaw1clEFz2Cb/SyrV1w
RvWRjbBJN6Chplj7DgoN1uR37uX4Yahj1YDqWajzQ3OdyAsvmodYXrcg40GFQaTc
+AZh7UKsEeh+/+6rSKTARzc7zzW+BoyUaUZKetEJ1U23fGBZn7Nh1KgGBw8obVW4
guG4a6SLoHvyclwkfr509skUnJy+dfGIMrWScrzpsAaejC6kxTQtPqCKN0ANQKCW
8vtOPV01JeeNhVF5hdnppz8V8CQZZ0cyKO/0zPv6zM+I4tWPMH6osQQD5WoEWckg
2UK1uSDVGn7o/wf6s7au0yL1doxlUm9XMwHEnhM8EP3/2z5nh41Mw/RFLHOVnvo2
92cxpM87HA+txlcQ3JRAAddKdF0Z/qOzINbZ7LbzpdSaO/VSpShKekq0DXL+rINf
5UgWfmnQFIfaVAa12fTXVpC8Y0J5GENeP+E4EpfzpGtGZVXBdP4kvTRFXZ0RBDR2
6Yh85EzGsH0dePrTrCc7xIwGyuiSzszV7mazWvPNFy44VZ2VKdcCupK3I8gmRWIv
LNvu3kLT89ZtOkVoGEwClGiq7YRSt2Q61HIWsanNLdYrgn4vhPsKDL54EwCvKDrh
QgDjaIaOXtI6YsMJvw4mQ7trszUC2YelnooqJsvCeT+vNQ0ypTlKBFu0dK6dnTFa
HQV1cxN0dNx+N64ye7yQSvrHZKkmUMxnTP9nkYu3zNSPZs8nQZs0a2QkvCZ4pvz6
DUU8qnaaWo9q7hwLN5vfJ7QJ5OCOHCvz10yoq8yZN3qBBfN24Uv6fXZRv4vgO0tH
yEJKMlcFxU6sJgeXHlVJXOtrcWRPCrtfYZzoGLYyvwnq9aH3uYLaVtasC04XAVlN
Pue1hvKmwRMZAWfQ1KLpN8jJx5Reg3narsMZzCO4ELZ13aEt+layUxBDbQ1MznZj
zrobe/4gjXdEWSrptPp1unzGwM810lFeFk4EgnAMAKtXUs4z0BEPQb64hCUj1xWY
8PeK/K5Qm35wc0FKzsgUin4rbo5KSIr/NGCqgm1ZuVKGDGz2cjp3hxtnIMWgvCrx
oXfryo4cBeJmxK/XcJWP2UK0G7tn6hZ4oTj97BIe7zP9ECJwdM6dFqQlHe5hdkfE
futg+kjI4TxEZEukpFHtu2OACP+GFEe6AjMac5rTfiCLpt3q4rcL08vXehBPAtsg
2VoyF+Kl6z/Tnox50k4wTJigSniOyJvBLZRSCWl527TE0oS4Tf9myw044GR6OBNR
sbyHNAZm7RiZ9+fMkf9h/ulE+2w3n1sWlOCOYLtZ6ouLAU6xpmT+Bq2PUrDcIOUu
QskQNNpV+iEVBP6a01XSSbHBX4QRVQ3i1TdvsjBEpD2+dABsdhCGrBwD4sOCDwpr
GKitvGY5LLgwe8CDsWr4ZXm0fyx0AJ4YaIijASQGvmtu6vlhUbJaPoPcolCbffrm
Ghflowh4YDB4n2M12EXjvJMInNV/O/G1dyAJNklE5IGPoQ76upV5MpdBe4cLxQIF
Of1AGzAI5nNWnodaevpgX9LR3qQIepEAWTM7/xq0kpzeW1FQAhzqMeQJPWucs9AP
Tv0G5MMD4SWutpBRxVEDi8+lmsXU1zH2EN8g3W+7QlBlstzukl3mxQzve72D7Qrb
UUXsWwdJ0LU1l6aMkjgQkPJmjt4kfNyZs8MTrX/yTRJNFshPvpBSXmImHQUzy6yX
9ljxJRURCsAsyHLC8ikUuEyZNFPxdlLQQQygGdRuH7W40wOL5n4o5OW68KR8wA0D
ysFXJwEiCk91E2xK7zNWnathVPVLyNFZsfW6RQsBb7OyXFKT/B/jhvgszzZxAmel
1wuT7uNll+84qCDtqcLU06FrmNyceQUQ5/EHhy6lALUxBocwzCMudu2/9Nc9T/Me
gs3HAXD/8WbtHTUAsOKpHzCFJOde3YkMet5zY4qqLBpFmW7HJXh46jwhQfueaYMl
bOsuScbgLLLqVqL5EdBmJXTupi+s2E0cPx6zuvNheLquGgf+HHYW+/+zBKUpY1aK
JCXUVg2SupKQORlcd+RePpLPDUyGTxyUKPhzVKiNfotnawykp2l62Caf/m8azYxK
3CukMDR3wHhs5XabC5stHJc8jzuIp2gp2DfrYaxlkROw63L0AYUz09nOEitWxAXu
KYP4mLXUNzNoDrFkTwLUFqIvGi2w0pY9RZnd9OP779Fit3TwZDtYDGwP63QmvhJL
Q4axVA0ABgHdsHp3oIat74bv4Q0swC5TKKiMLxI4G72O6x+JaL7C7XDOxkS2s+H/
QZKEcEKB5EbCQ/27IDMV9IJPjwGBGHOUqL281ZAfRsY53OoWUXc6rSCU5/08CAT8
7zXg4BiQxQDWJVYGqvv4EbFj/s/VMUyrHy72AITN8tboh5w9E4fG7dBiVnUKe1/W
RDcsjjzmLnpAJuSiNqIt7EasbIQ9YUZXRttbYo1K1Y0=
`protect END_PROTECTED
