`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H9QvwEXrVWWsBKCTl5iOdVRPA0j2RkEZQr3F//wldapvnlP8ApB4xujgnNf+oUvQ
kids0WzBgf7UTkjdafEJp1aDjvREls4y1gqNrSI2znmVU+LND0cOhbtWoOstR2Zs
N2/s+2lA/DRuxcyyZoIh54nRzMGqf52VDQLvgo9oSarUmW3B48Fa++sRPJiMYCfs
GJyLjk2FaFBvSPWbSdbZkT5115gqG9k3joEXeDS4ynjhuY5jVHYE3rWBCxl3U38r
SyQT8ARo5+6JYj/JzRypFL6eXs411UX5C59LfzLiDtcLBr1QZGHvVehG4OdBw5Ek
ye3vnU6tvjrnDbrzbLh0rvRBxUPWujpe0r3Qv+DU+GzK6+a8bCtiW/EOcgugWl1g
zNgALRpUc4IiyE7Z0hyurLP6WdqAHTBsdacNY3/1/nVYVjcw1bCGt9OMM0xTwUG5
WZyseOkHg5J9taNN09AXRzqVMfAJLon2cHS6GyVCsKv06Kp6O8+YdqjeN4sUO2Xt
ERh4rqcXxVPVyDQR7CDPi0+JAO8DMhI54C37vyxwotqMa5fh0mQXYTddIrG7QihD
qI0VrkzweQNBRY4gxX2SiiaE+Mhyfm5ozz6/BDQ9dxJLYR7GPXWu8BCjLg+q1/1j
JMit/DqiWdZ0+6fAlPDdcCs441TNM0juFtDpwgy5bKbSW4RlPVq9RkQq2zAlJmBy
q12R3QLu4G+3M0DUda8KjR9LEMgMgsq4mdBjp3j5IE5mYQHiE/k74NorKMarV7De
4sf57oGAFHVraj+7WKCqDb9tanPbfcWWNKzrk+Clr5UEAco3hqn49unXLV4TdBqe
QZKjOdAaTLgHQ7ZFxjtelVrgFCYZb9QnC6TBq7hHwnjNeFkq9LOQckDCCQV6ryQB
QWq3MBbU4oqVDBkq0yYVR8gy+bZEF6dlmNuHIfz+lxCE8+xBe74n3QMCt3Jvw3sP
key4iIReEwMJ+RORB6ztwUy1VLU+E7rkoPUVsK4uug7T5ZJ8AQGAEfRx3YRH0vRi
THUV+8ZRNs1APDa+za8FVWRdpa3/OzBw1UDG8eD3vi23GJQkMFX0gcybXUvyTVF6
fuIrAgykBxZu7dHw+dHaZmmK5pOWn7gjpz0XbLhAUdng6lDfaoBouqisBwoTdVdV
ZyMRS48eMl/Ge9qQ740w0bYp/IHGTkBAViFt8jDxiUZ//wnxTqbh/p1kiyGYwKjy
5nFOS9K89MnJ80Cp0ct/toVnDEjHBLK9YzXml48sY5H4CzvbQsl86FShGO+iHoMX
hCa1TwKWyoiqhl4FvkdjNAhAfHPOvI8BpV2AMXCsmQx3x4GCAVmSWgu+2SmnMmCS
IszbNNZwwzUSO9PePYfmWGbe2giq+adz4cnMsqQofWRLaiamQa93T5F9ux00F4hO
gloWWhkChPjWgO44fM9YR2RcymAPttZfn6+6uRiW/GZU8RrnfhCl3v78LiBHUJh6
spzz+019js6X0+KwdJhqEjKnjgJ3gm0SY9jZ+NyXWxBa+jQ5pPHB8EPAS7N2CjfN
MXl2RrO7enMln10iJ94JGwmU2spAR2l+JBy3NFhrMNMZJYT/cy6tA878e8dhwf1Y
AJMfKZb5qzhidpzJl8z2lfYMR5rjPGPfSvTUO5HJ2bdKUKzYrhWPHhzceoXzw1Jm
JWpBOBK8D/HYjB7LirKpusnntlQGu281n2y6J9IJghturQSIL6/tvbA704QIVHpE
NbWek+Dx8BHSRJsLb+dsIYhEcwsAxEdW91HvmYbxc9jD7PuNRG1jEupeZf6VKa1S
`protect END_PROTECTED
