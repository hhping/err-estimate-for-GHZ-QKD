`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l2JlRSkHUrLN2XLpJF40KCi/gtlhKjhyXHVl3HKZhSizsD7gxoWi/+CFjjLRjIeH
U0WPDHjBiPm5NAmkLoL0MSzYThQbQtM+zGFug31Q3O4IEPdClQTGvW6iHKiOuDMp
EZl7FnjVZ8tJQFBg01f4b62ttY2ATwaC4Qn3DmlYOxuO7T7RllpD2ibtbPlKlHh0
hb0HlYzsXXYPBjAgBE+i+JPViQisKUsoR3eRMKqL6vtCOVOXrItDVYbaLEHMdH8/
TTXWF9nOVUcvnvxYY0Ppu1tuYxh3HK8PGxwENHLin815ZMSmjKhEbE7y7MaHHaRR
jghEpJfgxCbYWOEoBoO3bQ2a4BmL02rEdHZhUw3boaKT2K7RPQ8WuXkoBFNXY017
pm033Ib0LTabWcOMZ5Sl3xEsDFVlDiB339ShZ0jmdNtSrY5ESxULvXF7c0yiyX9n
+hpgXJqdIsZ1VXsc7bZ5e3F1e7B/DLBQJt6wDRj6A8lpnXX/81hYlKE2Z+HNxNrq
KuKANNXYEMv0b87k2MG3wN0D9F/Z8o/bmmalO0JkCZcFLI/SesVH/7FnpyDbs7fj
ihsCijDVzHIRBdpvri1OlAEUOVUJoZhcx+xkKO8JK+BC5ugknosyd/lPKR1gBNZb
eXj+7H/dy+Hss2HU+EI+ta7IyzUslcwAx65vMEBhSZLnaIdV/MByCLXpD65sVqa+
3yyL/v4ssASg5cdtB9FI2j9APdWsVCRyrl3IIYLTKyWP6aLct3bSEZK7bDL6FinI
g1qQNgwpXENxa+r89jmoWX8AQLN+C78Tt01+7SumV+XcjD35W6zMM7dP7NRfzOQn
LA+q03xAL65iE4xi5rGqr+DN4ul8tMx0+XE/rP4l1os+/surYp0ljVuJWACwnJ1b
wSajkFTpqxbfc4HSY0AXKn+34COjR1HhMNVDXGE8EOuYtYfgJumQSXdJdYpLQfsS
ajbmwIoe1QLNmMthCg9TcKn/wbMoIMVNmLc1MgLEx6H/imrFN7eQFWLn86CF/1ko
yLOky0MCd/zFo4BfX0CLD5MdWJmyK+wQb90+vn9sDeh45wOefyYgd4g7xSbaQdPE
wiZNCmKzhLGo+xHpWPsN7JyQs8mB60U/FCrpny3/yAiuxflIZsywQ7/wWXGIoPlC
2qKQLHbgZTYKOcaN7E1c7P94oQRfIXfwlnOynjye1SMtoISM8zEtA6qvdrbQovmG
1B0eHhS5Q37UKKJ36EsWD0CijbAJZTo9AqS06VZS+SCwl7zlMrf5xAkoc4asT099
27B3KwYsCGTnX2tyEtL7RILSETdjqFr1AXPTAWyY6zOxIF/HFb+pe9ikuuXTPq4y
68hY9fG3yE8W5oGwtD16H8nrkjNXEqHr7GSJJua0IrdU02TsJmjsgMj+1MxVXKRp
L0YjsWNOBJwcvRvAaMWA4FRdyj6MH0k1dh53in7Q3j6J6okHCfxWPQ/uTXg4BoWU
2talK0ObOIy5mCUlS17dy7dXCj3RGeMR7OBDq8LmgDE=
`protect END_PROTECTED
