`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w3zyLr/tFSuCUi8F3I/BjY/bEnac5z5PWxEPfO74v1fohYncJ8E/lU4WpBdNFJ6P
f1SwEHCeTEj+NV9ApDLNBoDwL8//4g75kXr++BmIwex4Fu99WbSKdVPzYa98NFsK
B5dJBZwxrsDP9/jB4x3E4ZvNw7DRroLKxt2jDgNoQD2Bw9rkMm5fPXxsei50PhQ3
abMYyJqyMUlUUh8lA3jRZEUgU11w9291gPiUpq5XRX9hgEwD9ie9jEA/YrnNS8c6
KnXmVnvzMeFA6JR06+dOQm2PanIkLn/FksXsW2G/CPS6epzyF5BoLpEOsA57Ez9J
1aQQlMvAWfMCHGVnyWgxeZNMM6TtIhV7zLJIDnpwh7ChVTN37RGCgCwhboKxgurf
1stjHL1zOoUAQT1dq4K7yLAxPF8atCmLXeDYqNHsl9NTSu/zrcFWWNKOEBwd8hRR
W4AvY21jrpxvLCkNSH0qMdGa2cfN+/EgccVC+9RAkTdlIda91OgcrNTsCUjARNwV
KJ7rHooXa17TdGCpa1BHh+bm7QP3R9eufkdRhQ6tm3ndHg3/VXF4BKRjOVJqldPq
3bVq5o6cKsZkCfQk/akpJ/nb/q6qfY4m0bxGirhYeWxuM7vvINqB/rQz5vBX6/UV
OHLTwxIaectDY/fKFMK7mAxsQ2LjZ/l8bVEOGmLVTHgqvFDOwV/zQWac1pNSyR2R
ZBSGzTfFXwyAFvGE1zcf28K3tdytCRvkfJhit4kwn5qLLCOlgdOilWU9EJIgpLVj
EO4MFwlYVhWkeO0yNnl7J/gTRv5ZEQ8BJ1Vhz/1s1Qrab8BSQTtH5oyDufsaQqiK
tL4T+eLlugZi5C+f7r3WRwYCyGwgJQ9wMZ8o/P+mxzSBSNQ5T4LzT+RJI/ZIp3Rt
VWyVNu3OaZdhqiRJFTwMVWpCC8kCwxxlCinuou7T2SmLVESm9e6+Qkh2YXMyYkot
Niem0iFSls2muXh+vj0ZN7+OET1jJhDdo1iAti20Jn+TXRO1ikgW8feg8Zx4wqd8
j5Uoa+lrn1MiSSIAT4tW3ZrSA20UkXpqlvpxGiAnpUtMMw0OVcQ4Kg1eeBWWqFah
ETnrQ1+MkJyX4nA5eomFKe3vy6YIlnhagQi3slq99yAj2vIxkBKshYH39qRLqtP9
8D8chu157Um2jIM7Ap3fZ2V6j1nAP98DPQYox7GFq0GAHTYFysmFS/2u/vYnOqNT
qL8rZccePpryBMjnAEIV5Wpr+mZgAl/mvvGhlPOUhA0K+EwG5cJM3UAhO8Xw+w0U
+mvepspWsxabnvHNjTA83zEQ86DUNiirVEIcO2CsP0Sp9Tls3oMiRT+VHINUHLgY
JKlZl/aTnXekVxDahEb+7IiYNImSCttDemu6wNMdMERVuTa+YfSvyfDwwEGwmcPc
/ottRj7cCV+eilQhfEHGyNCxAvZUezC3RvulMWk3SUPoDuYFUqA3hYWIp5QBnnqr
6l8WtmXkW9gOt9+tTSBOL0bTm698zqJpATU+Em/nuQmHZzj3PONMxr+zto/1P2uq
HYzqbq0TUfYxxumYPXFLxFrssOkaQ4y1lAKwUiw76opAkSHYyMCePcD9N222fgUS
2/gKCxvtmfpef9u9M2Ohj1DRw7iH1MepyAOPB/RbLDS4P+Ri1epP1IkScJAnEFbz
QgnEm0htSbqZZjEJozflqnrfrM6DU7OWpig3pjAS+FKCmgtBmVa4HMqfXVsAIGdP
ZJ5xMYOU1JBIZTzFC63Ncq2Cv8e8qYoHHNMAsWsyRI5cWHPfc7xAupoa/mV3IALZ
veuBH7Nwq7FjnE63LLlBfH5IERwRoSsSkNgmu9LNpBRVqe5oT7ySesy0IxaWRW/K
0BJDR7C47i0vP/v4lt11RJkucTsxzzC7DZrzMD9fpYUyxLLutAvjG2ber1vCoFvB
05Z0tso5zhjIL0K5F7rWElP4j9EOzDde/uVEN/OfEGA0qepEvPiWNa1hslTCGOKc
3eB4ytegiw+nvgYvNbVKn4dy8pNt7FEk8vSKHniY+bAs5ligwe/Equcn0O+AlrQZ
NZ5fFOlsdZ++VdUqrpVa8snPSIA5ebJM+D5quntFU+brwWkHQziaCgheL3d6DMRU
6WS5Fje8Fn40n4Yh3JjBVsgAiZ2TARF7ynCDNE7PMXvJFYx4+KisBpYYa5F4/T0W
7P66lzJrQL4wK4HO1eHva1JZAY1WFfY85d0eDTRcMsPBgkXo5HwLZGrewFzKz9CZ
aZdr9Xxa+Bys6gouIDmE1lkVrn1wzi1iQa1smE1k7eaApUpAg3kljEuwfjuPwCHo
BYDnBAbziunWVlL0z2Grqoh2nziJ/0+K297aSDkIPNTooTEtrYss+83/80fJXviv
bO6KQy3vPVZgAfGZPNzuFA5Rr/xg+51O2ALkzb6fe3Zd8q3O8MnoJZSBEOKFpd/J
ZEV6ledUbPLOotw1Be8RBSDExvUMqKqofz+dT4x4V/clOQhJ2gdOG/VJSD+J0NeD
a4YXBgn2HqMUc+Ya8gyJtEK0mfkWNzNb7BSDMOSiRhxWTqlY2CWYAVHhZhTouTyI
LX6hBGDSHvFkC54SmTjFvDt5GlmLq2MmshN7RmQ5nHdHvvqLV6gOCh5Fh5xGGwed
iKVgwnNzKByPrIO+7hmWJkYqhqBlGzOdt6u0AcRlXQ1N1eG1gEvxIBvh7TrPSdY1
01U62nZUDpI1zfB+gYudOE8fju/dGEdByyGebHFyI7lIHwZl8Ih15ZNA7kMHWHNJ
S+KgOmgryvX5YYyXv0hqmqUVXSclyayVCGa/bmfuUgTyvh51Ie4bYtp68xdbUPCT
CG5e62qvDNXBhhzu4HOWueQbrdUNQbqj/jahyx6p3puD89f28aIZWMq0Aqgr1PpJ
CB4/JbiWdySQjYqEiL3a6la5u3O5OHAcC28KLYE5SXoX68wPvp+WyyewovafVxgj
Bg7EzEPBfmiMgQLOLU1666AG9cXIzaNohlPuWgOV74uva257rCZFN31+ai3Vjflk
OHzvCgBUADVRel9PmyzbXbm/qXWye3vxgk1Wbc+CQIF0o737koR/e7+r9Tb9CGsd
94f1PELFV0ATNkvNuN/0215RFlfmDWskf61gZ3SuMac+dd/Oqco5NDWvmStYSPpA
DeKZC38mDjcpHjMTzNaYn/jZbajwSQhD05c6dvZUhd4=
`protect END_PROTECTED
