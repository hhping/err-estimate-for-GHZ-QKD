`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6L0e9fybA/sK4vd31BoRF+hyztLQWtTFpv/KZXjcajd4+6Ec71Ywul3XzMjFztuY
Pwx6ys15Tmdrkffscgayx3YtUhbxXzRV9DDX02TH0pApHAQtAPOfAmvAyGUrRJrQ
PpkHaElwmeqzb4PD9dCwwSqZtZV9s2jmRUfdvZhGhsS/VIUFdkV9B75sUaqHh2Bx
cm1Z97tJ+DH+PDGh3NYvM63Q87XEoiv6+sc5PZ4vT0xcgOH3QaqFdNgMXmu6aNpB
8/penDw7bUFGNquWCwLOL3YsW60iUdM4A9Z/ZKR8XPXuKDfZhCZCqVi+G6cjQ7yd
gzuuFPv95X8O5dhjJft+eIpbpBAMxvYHZW8bsPUsJzLUsrAkN+8Im+5rIW3pGVWw
R0iwlex5MWTXla6hFbo8sxZwI+bs0dz0VM99xv0UFIoBW5IoC0PWDizltJj4Qa8E
nTo/Fd2SwU8udXL3DTjpwGsTE+sPyIplYj5GKvOmI9iPIdUquhZeS6HZfeMcOOI5
4J4B3Roe+jwo07fJh0cCk3E0fyGzRxfgnGNbQNgfD8CxK7iSChfCq8XTJxK3zv9U
xat/LNlz6EAkfyItcqXcp9A4SONw7291TNETSV1tlc5yvnsHtr6Hlc2uUb2tu+qN
wKmZhJiIErG4DCMnenLJyHYm4LXQT/uBNX51Fhd0aGKelDRQoO4VgLo4pkV5Yj2V
q5wiTJu9zcfGjA43RJ/wu8nxPXXC13DOoEeh4NEF3gYkBPz+LT2xU3gSSy7365ZZ
oQe+zS+KyAyKvLuZN4rGrfoapb6Fy1P9zOCo/6QYlA9kXE2pupu2SNCVrZqoPvxI
//202l09utbvYlvlQkhgYlfd8yvtVnMExmF5uWFPy8B5JONyIltE6EBT9dNBOzTY
L0kfaZ8vUb2f7FiFmrkjCsTvU+0Ga4nqgOa0XGAc+Pm08ARxRe3a/3HjYb0e9dTG
USmjIMdtSV05oJT/XGZO+ystYX+qLPcqHeHSDE0i0TLbXqBF61NfhtIxW7o7F6XO
LnANXnLPaHNg8j7tTS1UuTWBRTWVdgU9mtUUDHtf7URdrf5msrYU9vzs8Vdnan5a
BfgU5OCgNMbDxky74L9wiFLHILLiqDjNwnLGuHKmMu1lC8Cp1c1Bh9d9bjUlBFpt
RA2+O+QgRkTElXdpp1iomRP8fc9ErLnB0uFtVl9DfmqFEnIsHraZN3fYrjR+EePz
aC5Drq18u/d9xmH1+KZh0QYkBuYQM52x8rJBaYGXy5H8MvsVpCuKGMGNPXuDN8CW
OFQ3jeTzn6Hhplc8UHPEDmR6mxHVfG0LkUZJ+apGF9WKcG5CicUZVyawySqyqJhk
ZxGQyY4YOr9JD7rZGaS7B8/HxWH4KNFE5UNJuCSz9Oo6dJ1VRtwEcevJp/i5QAzf
6wTnGp80IE0WGvheA3Ugcx+VB9JkMJs9PReUITw/rmkFmwaYP0xNaKGf3VCJUeGd
GWvc8445FqkJ+zb5oXjI9Yv6BrZR4mq1kQHfKVfNrJSk4Fv6VhrQRLtdkfnRuMcE
HC0vt/b4mLn8zYJV7avqlUhTGnfxr1FvcTatzuw2uIM=
`protect END_PROTECTED
