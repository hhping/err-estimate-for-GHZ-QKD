`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fSyq/k0hawEo/j1WnpykI585LEtVCWLxmcfOr9h13RE36sSt96lssNBsQv6Iav0a
pr8dsQ+sczdH9S7tHbmGcmGQWxQmVR4FHKL5RwOfA2awsC8K6kI3qPHFbPKVlCal
BB4pgkM1CwSKIiECrCaPhjkO+gg4PTdTvXoKDkY85JWCkSBRpvorDlVOCJr5O3JO
j6rpseQVFQsym/LtuM/M5Dt0Uyo47cIU+fs1jFmc5ysMyCMMbL8KlfjeimwIBmVa
u2XdDusLwNFaECDDJX5JQ72zluGnO1WtET838OWRcYU4prFoVYXd+hzKxcIwlXaA
zH8PkdFYP8c88wEmAJ2yl0keyK2QWM04XFNQ8vLuTc+5wGWbvJOwSJebM3dFOy6y
YN5rBAdgkWnBXTTaovHkib8fG05FxpoTkm7hA59OJqn8PW72RR3VxApHW9ehpOf7
HIb/VL9SDLCzU6mKxFv7+oi6Ay3n5iGQt/+KNam3UG+nuhDfB6IlRiFBSCJKGRlJ
3z287+EjvOR/+F6riSJkW9wuY1+I5Hxb9JJh3kW78bmZigHt/NI1kWMvNo0i7Ed1
QsbkgxF5MQviKS7npg/BYVHl954BIIdO4WGacaHi+6lSjS6mqNbRMgMNMnsNnIOW
s1S7+7SbXYOmuxZgksiFvZhxDeZRnCFLaFVrz1tXc4uf+jNj69Ug2lluvmAHBwoF
O6RdgqTclE+7LDNr1b8yUm1bPex0SxhA+n+AjGDX6GxCRf40bmSNwrQz8ZjXr4Vo
5b47gEBHms7B4kv/o6zMavmhbit6sWlwBC8PYtU1T0Q=
`protect END_PROTECTED
