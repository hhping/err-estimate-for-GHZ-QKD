`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8sFKVyNTuM99ofPcWBv/YNYhQSoq/ddXdo2ld7m5XpwPJPGBoHvfLO1mQsBDysnJ
3ZJ0ls8XSHg94AMUW55iHftQKiLq5xRAfeFKGaoC1kcpFCAfbZiE2/aVUTUkWXCh
aFVE697CIzRGkflF+48SeFU7NhxmtcyrXOzkG+KDSD6cZGpi7RL1Wl2GsiOu42nH
nWxBsFzcl4sFfOJZyTwlSb5ul0pl4c8i7ZMxHTEdqRelu6ueXpj6ryk4snPxCpDU
EE9yZ/VQzl8LV5DehavedNVX/pFzEkMWDXXrSMFAYM/7dDqMAPsy3xHfFg4dL+5x
X/IF6FAZ7GFo3pMQY/HgdO9gkVnq/ZdCcjShxPn4k2VBNVQhhqqCqDMCBocACL5v
RU4B4etRN2/3gEZ7JJ6Zt5/SystEqdcejhAY8oDvWA2ZAYOPKh1QD0byu+5mHIGt
mb1bfcLPDfWuekGg/dsWTmzGJWsHpF6MnE0VnU1PcrV9Wb9WQNxHSRd+pCTlmpdU
dFeHEGNIvlSp1qLpFvD0zqW0erl2bXHMSFjjMq6eDjaQrfm4wssRMODe+yoEsLVT
UzyyMXUNhWL5/zB5pzZTSCpAnbmCUaiynYdyrZl9sbPCxPE23/NVibDMm0dkPHQs
+TFOf8/Nbc1XTdevkysoWr2lLZM4ZC9YwgmBpEpwW7CLfrcA2xSXvxmPsVbrfWR2
7VNJfKSaIehtz+o/fqMaGvGdWm8ozw/CZdlIqfFSZ6g=
`protect END_PROTECTED
