`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q2EW8xmKJ6iv7vtkMgge7ofeIj8wNVV7pbYBmUgdGs1g7dqqTN/SBRroRNOmep0p
uwHghBDtYicJzi4dE6QnG+GoUZ8ji0c52BD9EOHR1vIkj84mUun1I85WglqhLCYz
div/nrG7/IDLWJRSyT0wnFGc7abJ29DZkGA4h2GU/cptYkGd13OjbnXAcc4jx+pF
Xx3V0HGpkbu8pQsYjfUjtgXtReOIsm7xncMLyVQlmqnKTx0MizNgU8T4CzrRtq7R
2SjBR0QnYljqMEJxBhVjxdgJWuUsfHfkZwCiFsdOkIXjGNr3MFBc5mWnIud6rJz+
kgDg4naBAv4W8B9n/v7qIXKPqUqC6xKJY6TTZR92a5T3m3EpiLWzETKr2ui75/jf
vI2WFJ9qszPZ4bhjdZvOXE4FVGa+ivLfztZO7HACDnmctVuF5fBI0qWjj/H0GXHY
NcpI5TX3Abl8jqlRXGbG05eX2twHzB1k5eouie8nDtUc/YFPMeAfJGKeEiclc54k
R+YGkeQ3hIXuII4fZvSKmkN4Z1ix4gCyscG/I9t5T1VULPayNzl+B9HV1RAIYzhm
Nm6WsK7gQSqiq+MhSRcWG7N4Vw9WbrgE6PgUM7jYK+QVgEp2gq4HuO/96CvUXu+0
1diWjHKGZc6D+59Pc8qE4vmK15ocR0kCW7j0vNdoccQU40wFrLauLFl10uV1wabh
HR3/gXjt9g8xPQ6ybufwY9a0zpqOYU2MViwa/4uMCJh9TlUGrdX+QRrnG2NhRqpZ
`protect END_PROTECTED
