`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rsFtkM2ApjZknVBTRY9KuaqaXBG3osGPp5GOG+opV2IB5O1Rq8xbFgkpJhWkrRU8
MYQviMpRtDcAytEFdVEDx5IYZAu2pcFfuBW3ByqlHUHL0uyWc/OMJAbzXubl3FB0
BEykBOj3BEmOhScq20RY9191c/B9NOdfMJ2opSoks9AFpP+FNpbYU3u79GFuTGFL
x3rLSCy8ijOEh5rGSqJE7hxr0Ya+qNopPcI4IAS/n8ANWiZnIhHGwxLq+Gf81kJ/
ni/iU1y6CLIAV+K5yUcS/UJjU3QONrJ7jd4P9VkZ6/1iSp1bxlZgPwNxOWMSCZyV
HqiwQGkajcG5MnNnh0o3ULhuf6bJcEBXdLA94nVe854OVtxdbvDYe8q8vY7BrTs8
HRyJWAMxDTp4fNJSZz4svokpPHMTXX6smELHa0J/9nty8jhVmpViyuQxj232kocJ
BwNtV6cDE+lxzJXrL5CicWMn+Y4c0DBatRklc8tuNlzRWOMs+QsosRJ5SR83VwLk
oNHmEuA3DFtxn9lzsEPOFDwy4o8wa1Wlj4lNahD7FH5p6MEPc3mADMde1vp2hDo7
le+ReFgFI2Qp7U6upLo0/jG8uun53xt8gFW3BZ0hFAtQQIVDa7J4AnrgBdBNkIAY
SW5I0PbA4z3Hj+m9sNadJqeX5e/J3zGmbWGgFSKscuKNWPCGdE64+7CCRfG3WOzB
KDS4blkjOHPsjLHCW5nmYddgxHbRulvw3Fb8sOa+2ihLETOBfMA9VTVYEYSbu+uX
vgqkfNjJ2PWvTRHDQKlfhkmhVTnZd1xFQDb0/qyCR5IFKZ0aSLHoZ1INXLgPspbs
VjWOWRt6xZlb+JFJkQT1fyEjDo4AhSnHx7l9gdg3NvulGkRpN0AlyBlcE7CVF1+T
/1R89YsZPUW1mbInY8gTt73AWYmBFKz7DnBs4CUOFkA8ANEUDffZz7JfN/FLq/I7
vENQpV9fh+2hX+9Zmtzy2GvCT7Ugy+uPjzGAWBRPOuv7IldGHID8oWWc1WvDdEce
Nb3c6+X6f0457Q9X5O0Vrwu6X/nsKfh64bpGrDxQy5IMkFmJnHOnts7V+5KXnScB
I+7G2DmOolZHxVgdUmu6mDZ8XeHroF54E626Wv21QfWwgQfF8L+UiSZl3//gTw9S
sgh8ZDmk7FHj2YcDFMOLx/ypI8+HYdgBOSNRNueCAW/wa+eLGEv8uIMP2uow6iKi
dqkaKnYNAYxpDV5OJgRK+TgDWDa7C63Hw85sHoQyAaPu4A0RFoV1eeed1U+jWolJ
cXXrzMa3XbdUQujcbMoyz/MZ9AED5SC2sWI+mX/N4DSTsg1XVz3t/5UjHMJRZpGy
QnncPPLJ0QE7XttNSM6SQ04TnqkpKGg5ylWF6jugcgDjZhmYqWvGD69t76dijgfV
jIorIgQC2GokidSRSi+9aEoQxsnaKWmehnOq1Pg35T8p6aN/i0wsU94t4t3oZSxD
JmVWysLI8V4xjVLoPkhInufiwCjh3KaR4WnhQYtfSF4M0LHBfEdGtiQ1NQ5lujI3
z8bML23CrZQvTz9GoPRQrFJyChilR7CzJeFRBxjoe9fLJzw/ikkxHjG/eWLsUflM
JuQljpcJdS3f14NcSh+LOg+1jFaC4AHYI2qW1G2ZvneVfkAIK6R6CSl7jIiPz8i9
fRKa5MXOiOzX4lb6x6D1jWxHVcRuvYaKU1jvOBhXY5soQt0qUpOPPYvlKRw0DhOg
jbXNJ5UZzog7CQZAZ3//ZdGpL/k5PT5+urT1zb+0mmchB91ZxxLjC7YCMMygmNni
Rev4A/TkJ62C/WICX9WR48eswsjwXcX2iMun3npp+oqmyiygijFr5x6tCzXFPEGY
1ipy/anyLs6P4K5v7eP1RmvxhiJafcISOJpJLAFDosjZpAjMyQ7rZL3DVzeTbJ/F
hzfbJWqsWWP3WHqFy6SgyFkWl7OesBQDHBXuTmjjVu8+M+3s45SEOT1jO1or2oAv
PFjXuh2VYWJjIGht3Nzgi1gnUMB7cW/tBaUl790QZ9/9orwdt7PmX14yCwgwg31K
BJlPFgjJhZDWxGwIZNLXS7x8AjtfnhTMTYCks+CGpUSc1DjBrRMacqpFt4V5nQ3z
E9ct400Qoonnc/Bvptk1cLzeKNKnRqZvaFwKGaRyqyau+rUqiG1Y0MMoMIf+RyZ3
qi4F86IWRMQvI/WpQn3D0TJxaFZxMZzI2hapNB2RPG/xBkCJ76/nRiajUGdTbbTH
K16nlojSNpM9nvOpZy/wGWg+VHlQkYdPyz5u1x3En4fxO6zhiDl48xiGjTGEDodu
p6PhAGJlcuonGycAn7G+1SHLo0PMpypqWkYtl202Q7Gn9gr0eFiXKLioKg2odApH
MFZdG84xe01WSMSVvS7Qh+5tZi8zkm3M8Q8KxyCvaxDb22qStmkJ2I3hAdKxg4wZ
/ym+EGcn5ivZpwAnxYM8/ZIsggkE77W1KSkO9LC8OBNP/SgEBr+pvGShM4z0E805
CAiyhxMSFRISYOR3UexyK8HvF+FOiFzSm87j0rSjhljwQ0OMOjrqRR1YmmLvGyPh
7kEwIWBxLfZM1ds8YTDKMIyCqrd9wegTLtpsOngvhpUCmrm1442ShH8SJAEHEjLg
EPm5rjKjHq0kcFfM+5oaC3b1slcOB1g8WHDXvFiu2OqWhj4B92Sb38FHoXKwGxp9
DBcvFYpJo7l2VAdMBDDCQYQQu2PMMV1B//BGpGkFcUF9UeBAoeSxYGg4+LADdu1A
mFc+MS+89wFz9cBxKM/PMiXHMd076pX3w83xxbjCJwaZNjKZa0XfIqkw6R9MIQCJ
6Tcf5XXCR9vH6GQUArhzD3dUXXJr5iRrBuPYPMg/uDqrGuSuM7UPwwXYoKo5EBxy
SMamAI/ofFFE23j0iWPn+bYJoiQVpQgMLBa+n66BFlZusZYxcovQfGwlXZS/wXt6
lrz10xTWuiMLCvlfonp0QVpG5jlKOj+a0t4RuvgoNpXYv/Hae5bEoG0oMa3EWGNz
i/+rS7tFUL8L5x/l6QfnbG4mwEg5qtEsY9znxZa+Ya62LdXL0WmuiO7xG7kGnigZ
VwhxlEuhZ9IJOUXheIKPjmUppb+qfC1SCgEEDCNkezGj1UE8/o7wdQ3xfimtNDVn
uM4ep4Vehk2VDr0rpbimc/kg58ZOV/rOVW9EuamNEIeyQ8KUQ7MIUKulOX4Yj3lO
v5O3f2pCp0wXaSxsmUSRMGBX4ON6QY9YGzbA/HHj6/hh+2H9jkkYdGd+kNuyHf9q
zrfrCxnjecaRFGDzBvUrrA61nZCrH8xgU+7j+swnBSkBKUpQkmhXe7v5eCG+A/H3
f4oIdakNfuSHVKzPT5kO9uMRlOclrnbgJmhxIn4CqkTJnO18T7OolFr7QQNlGI/2
9Lc4siG/M7WcGaZP2DrAR0h+JnywqVOIXbX1sl/zLLZW3rjo9hcS8bSr2V6/p6XR
41Y/NvgrndPd2N81E4bqfe4ICKbVaizVtpba+rXLMOLlOSV5XmHuRODvHdeNg4NL
uOzZLx3PXspSYYT2RMWfRYvNmDVsWBhDsx+DpI65kOFpWkQXHgPu2UugBogoGNLU
HBC/ISgpRXG+3ziqiFsk2wL0sBbcjI3XjTSifqoOqXO7ckHc5e7TVjTbbRsKGNab
YcfowfWeTPXayR395Nt8VyMTid775QNgc6MjLc6R9HMjHfoEyRgFHKBp+LBArmec
y9oHz/b5ISx19tfvsJr+2bXKcPFqlNr3vSAJe+Fz59ev2aIgX+ZU6whbv+o5YWkq
yOLeBQr7O2y0D9kEj1cwJm1psDMvwMS1RnaX2T/flqul0DdTVfWHPeYYeTU2b733
dG5OVQ0HYfRoraKmJRwS6FfbZBiPXsB2+46Xcr16bvg/IXte9eQ/3mWziQKv8oHO
hzO5smKLCotm7pi8NGzsU5bITG44yOtbbcUZxasXiwNAf94cMT23giv7Xo3mfHDe
la8lboueyTVghv4/bjp9OsVEPE3boUpDId6S3L+/B4RSMIjiYWSRYfA8vAZfqfw8
BVdmbZwJYgwxTis9E8zhLycVJKHsuk7mxllZhYcv1UXRlFUb+OthtcZO+OF74c28
XAUinMsKP42r+AXeS+Xhu1a0LQ+rhtR6RA1f1YYtUmlp9jJ+ZeoSNd1kmYcqDbzc
V4XdI5QnB5zTgk0L+8BiRpiC+d3Bw9s7Xr3UGvP6E+kS4yrdj/uvDjBRmhFeCSL6
sa/PRwMxyn80hEKhUUWSmc4MbVQ3aQDr/60RGJwy0JVH3WfE2bBhWFdPlDEu7ztE
WKafjRB11ZapcbUzVYnMNyaSgNhRXLQYdF9LicI9fpaWFijemCRZZMKfpWqNTO/g
GHEp5leXcIDaP6BwNse3Hmw/Ut+kMRLL2ohN/28UoFEi2otxpkaR1jOGUF/jQCOV
WUIo22EKB/WuhKhobipscsRQtsqL92GlL7ntewWbJPw=
`protect END_PROTECTED
