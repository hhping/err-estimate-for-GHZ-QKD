`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NOz18kewcErdyf7brcl/2HWU2EN5Bb7D4bacMbAog7veHlWbnG6Ra9T1nNtI6rVu
W+z4ADC1mM6CjE4jxivQzrmtXGERXMHl+Mi2NGqgH4VL4h+p7HFi8aokXqRJyBFt
9ZVEvRuSPWzWwDgoOcNmZUDxhyhWHIH0+/tqWhVPmov/4ptF+ov4y+tiH50p4wt+
bz6nNtScHYM6ko7jLwAy0tkWiBg6r0UFClmEbH6USc7I6kYDnvT7531Yn0LNJiMk
Y4KntG4G9mYWJJ5lSc/fLdOIRezRtpTxTCYlQj672NYc0VB9rZv64gi++Xyr6PST
JjklbPecJTG/3gFialp8ybQICgX1T48ltc2DvOILngJWx2v1V2YAHyD2KfQd1P5b
3wdj9vWOcopMDWieCxFZe7v/TS4kzyVR2qJBgKzUpNsHdzJACbQJURawhKHueF5g
6+JDZlGSfktlrI9O57CBctNcIyytJ6KJCzNNhfVefunNfCdNStXiQmlA/4Geq6ps
xaboyxPE3LLkznMs1DZ1zKePy15Nh7uZDzovsSfmS8QHY4I4w5xXaJ68bNUjaNXq
aP3zVJHjN+EfRyXpG4Ila1lf3SuOFeiawNBbwmJjHSS2OJqZuUXJibnbJ3u5Sh26
eP4tfiQ7bAnAspz/LZoV0rfSp3sVMLj3ipMkGQ9zHL8ArBIbn1k2FZ9/SPeSNRfO
vo3AP935Xmp+TV4FiTxlxGTg0PnT1njFU9zc0hJUc7mDLuq9/wbT+BjvUX0xZMLB
5PVjNqHe0H73AitI8XON4hD8GWzwYuoPQ3pape+8LP9aK6+NSufljF3s0vHDl1J/
e/8iBg8C8Pn7sIH/p7vSbCGHRYt3AYrSfiKhHMpc4V21V4XTUftGcVeBDCBwV1BI
xI9Ty2kEof5k/ekA2f7Jvs/1oVIk4I6GmEHDw8CotUFyyzjTYVAX5YOmHSTP7nVY
ujeYEQxWKcWBvjCY6rFj0lachpYhvkfV7JXIA3VUPffqJK89kob8Py8UfDAlHx+H
8ro9fmp+zKLFIiyFDY1aDaHuHHyJa5WnjEfL/hg9iFmL5J4mutuen5THH+cIYxet
raoJ97X+JhajLFscrCeFULcPC0BSju5JxHWxrySlWlSif3befZ6ws7QeeEVVF1Sn
bnCqte0RLoVY0m1Nm9N5kQq7BJI8zW2BCFt97usWQ5bWah84hawZPjQi++3BxIMp
zMAfoElITpVvT4p1ZsimtOCsTVvDlOrTr+YBXwIm0zA=
`protect END_PROTECTED
