`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dAHlkNp/fEmIgraSxKWSMfLc0Hxzqfh3oySaZxRLeA2z6Qnz1stnnx01ATaL9AGH
ZG6tecjtlggZtywRY+rCSX6b0xIqHMwy4E1DtztswE2FMFAuUlmui6wh2R/XdOkn
zYzHs7tn6f/7doVmKSau8D4ICPDIzDvWniO66DPP2O3FXt7i061PsAUTOK19cJ5M
s4GdIOErNRvyBWMYVRTFXTMw++5wGE4NkI4FO+e0lMyxAolR1cr3nnJ7CbfVSdeD
SykD/KfAr/8lAGXyTXGDcFEOf5B9c0TJrx1aagPaLv4V6kz1oxNfEELN69WVqHIw
meW9I674G9V6fc1BH7QKDFVzhFo21jbYU/Be00f/acCbSDFBV52w/nWv+k3RnUEm
zUbt554gkKwe/Nac0X/MSXhoSEVbPO9QSfk0V0EiKdy1NFWD/4JfFP62kUCsjJgV
D2z07xEtQUQp49TGd5HYqqxahIBRKNwD2nLV3OEPbfv38fYfHaThBLgUEZsbk0BM
V+w7Mxd6Mn0hWmF5rBZ3PG+EIePjjWcfRr4vI3yJ5D4ung63h/Jr773zfISy2SX6
si2OkrVaXmq65eDm/oBiE95NA2Y+I1f9EJ4UInb2DfRcvDj6KTH/Nlo3T7vuFeT/
wQeAANWiwYuc/tp+q62ZvCMYI+C8Jn1TMnzhyu7Xj2uQzWM2oVldmWdGciMoXzbJ
nyjmE/TR0MeoUyRXKHhDfQ8V4MytrEB1qZxyXpAa2cbyMAYDpILRaIJRrhlVtWbD
mch4f/4uFKeiAoU0LEPKqxAo11sdKWdcO6aYf8wyOKWPm+yMGdRxI0LM0ihr0+QG
m0oNZfB853ZVDJIgyVJdYOukb6l/STIFtruMTezkqwIFlD+vlmkM1bSRSV8MBcS0
oJ/dYBvIgIElc2i9Ro+nZOxvl+eP8D19Eddot61DZM3qZmcL4pfPPlbJJrwsxTXK
wmKDbGP49G5ylDamjFv0tUqFPkHmoRfKvRVR4vwT6+y9+ccKuPXrfx7rvWxj99Vl
Jfr496xMhvzvVFccZ+/ZW9dHemJ6xQVoVneGVb+QCS3DvpT//NgDL8hWWY7ucP1G
xSIP+RNpyi+uCKyE6y4ah/4GXB3FAxJBNHFBkWsQA/3n+7jUkgRKkzZlqiU7f3gf
8FRquXJCSPzymk+kpxAAaKudVwaTLnjwK5HAzlHioS4fqxOTgUJSKoSo1GmlX/oc
ktj9opMmt3kWY7iavth7KDCNoaI0BgU6Jv7Zdc3tFmVOY4Xak/pr7Gp6w9OvO34G
0+uuf0s0a+s8XegJEcHiA+iBimf9TwJQX1MGAyrWllI2GBO9hbeyLg/7FZ4J76eu
EDqklvlDVQ+/DeqqweYwjfQYK2l8gcD5Oh+NCSa+7ahdcs8okZ48VieR9G7H2ypU
3Z9EMBCGdEfYdq5o2O5QoGupHYbrb+G6EgVONFqi0D79xSOEPkXOftq1oMnBEmBN
/NoHsIV86n7CuCr5sHhBIgw/nxw5Xm6ZhxvyxdBFgSedjVyIDol4aLjsMxtHdrHX
3AXFV7N1bwx+309DwLkrMuE+Lg8xUnm6leWGYYdU6lut3P/XK5WJ807kK11RD7LU
Chpbbp1uPAxURR7j4YauB43LOpVAg10FK6glnUM2JneiwV25rS1p7C/tqLx2x0lK
hUXpkH1BjYUhNnbq0zSxeFfiYx6FDJ7G6VE/309wtQjGg8nCBWIw7RuwKaC6Ms0p
ta8+8jeu5eYfRTHYPz2liwWGoD+EjnfDACLRgBfhaVxzJSNU3QUlPSSMZHN6UEFi
Ofe3UjFLtoWMp1jsVWGoq8mGtoot9w2cCvm10PDC/ijboCUBVKZ4QJOG+d5VUJ4b
SvzrNdOwe4nK0EkX6Qjqi8NyznMnkknd3hA3zWRu+3VWjsOgbldd0VEWLKLDXrD9
AH2RTC3iscHSapnolpCqfoceSXKJUxqx6mAd3AwazigayiswDCMv7L0nf6XgYH9o
8ZmZvBjpxhK52R7XwxP6a081by/xGKFdeJOcaIA7ey4kXQ3L/Oeiefm6XMwFE++A
cnC2H69KlwLm7wlZuJwqWLnMdpo/FTry+0LBCAgmKoqnkkTaHoxZhnHypWhJuz0f
90YaLarNsOA988NW9lLBuhJ2mdN4EDFw+wGyDkuopMXoW6+tuRpXeBVm3PQ0QDbn
iWU0ux/+26mJBqHOsr/tACbplbmFj1AmJ65qWa8UBT7BMuV7+UOVMu40zDE/34ve
KV9PeKpXgIQ28B7oYqN9BaBIf3tGZNVOKgkav4VUP8kRf583ojsVDCKJwoY3Spf1
KJSGRWRo6y2s4uvERugVxno4BQaiiTcOCEHeOqcgpFuwSipJUba/NFbjH4uM1fx8
1y6dL6IBDHaQvV7IqyIcswchm2VmbbOoYATwTcYD1oObMal9anRIxNrFfUFD6jbp
B85cauPogxUwN2sYGtKRSxRxXZQPq2p5DcxZuA5c/hBKW6iUlHuc/zHS879inrYQ
TdMLqxCxP3KVAdNmMs3NGVBxd3Uut9jvCsHhv3KpgvpOAvhPD2JGFKEXKzkT0IBp
MttBCEL9hRdELifPcmHpwi2sPGxqNBYn9HtfdGk+F3CfpvNKm6M2c8aZWg8H7gzs
4m+gieEELrxmz6Y/qav93s/kY/qGeWWW/IeUF7cfrC4dcOONeqTBGZlfB4TOyT0u
FEloIAOWAOdFqkJJR79voK+6xlKYeqAQoRAo30tWeQ7EC4cKF7xiAKqYg9GUw8Mu
/AZdd4RhRF4VtMqJatk+4iWoSvOyc4noSyRRidu+u1qnDN0FDttTpE6S4R1gQv4u
93m3/vesGA8XJmC3C+hhEMAJkGN4wbkVaL6nFb25WSOARZlZQNKipsYLig1ycS69
SmfxtWxRbkioguPOwzJWq+jG7PJB11ClDBMtS0AFPPQrUr1w2cqUIpMQr0ZY66fK
XuKKhLK0I80lgXcwzctnSs5PSIp3Fa9BHggqSx/uWprxs+Uo4SVNG7aXB8y7kvc6
AbXTc+xGKMb7zkZ2I5M4N7EyXUs8m1kXU1aB4/V8lr4nY11NelFJIuArMRhsgZDy
sQqomffs0h9k/NtiSXvnXLBr2pVhJ/nYTl4S9c15Cuz3MyvNX1T/NQydk1rhbIQy
kJpCtuVmFHm2zX11x8V6TaKBh/Vol50TdDJ9ZfI/8YvVu8OpRdU+xnq/4T8Kv1yP
HYKU3QgJacqArbYIX4J9Rp+TlKeODRpta2ZMTzu6IDF6JpcNo1cpOTNq+c17jiZZ
ylnsXaNXKjvbxdgegMheKvd8NEXWExwm85m51gtIo1nSAih9YBpvVb4VyOdcXqFt
5zuwnaagT8jGHEyPk8wCdxHpDaQtDjbxOwRjdwDx3Al4atU7hKOqEG2LKQTjR/bi
CWgwrSGMwZqC4/zPt88e2cd4D5VYYuQ+ETUw5+maupkumVbeuooJxNAMbYnY55gf
xbrP/LteBlzUgXB7zeLWqCIhKdLrp5vUQu+syG5W7+V1TV3LwsGbPJOh+27SXHRX
Mowqd3BST/thyx4C1/P7HaWHMUIe0zpnyEoKp3GMSG0ynCiUSlkrYWD4Z97JbJ/h
sMH8VXvaw/8he5ml7TYfcD9KbCPddyqr01Mfoii1Y5ds9pUAgdAjInWAD8wrnnbm
gSbDHOlo8SpTySm5TB/qVxa55Ke7Sj7OzOqKitXbAZiwP1oJC1RELAyrgSMTHeFo
1V+JN4sLPSZLM0s7VJgTMsvDAU/nb06ymONm6Wqryl8Rytx4fJfzFTLaQ0gGNe9F
h0cl8wKVlJs5pp/Fvj4T3FxOSAx4Ol4DgJcOAmUeDqwu1DiqK/QVJGJ+/V4ZT0fM
GOoO4WyV/AU2dt7FahvnzYmPFRUWft4QJ/V1sQaPfYBWQsXk31k6xQhgKn3/QfqA
xoos/57gtZiBMqPTCKMrQr6OEHUzyrsYWs/HnfCicKf9+KFFRC4uwPb4hT7g+bui
tABud8bOVk1eCNklPUv17M0aKjZB/X6UgziZPFhtopCkjFFlAKOuBEq9lAzlZyTB
+Ozdgs6GB/Gh/OnM998+LhVhEvQO9PQ2h3qZYy9X1jI1TtVu0Xq8/5gCSQXs9oV2
HUv1DVAxQSMipEQt1ssAd7Texxl9L95M2U6VOy4aBb6eku6aKito9jyqSJsoEKXT
Dk1q8JLpS6bU02CCiex1CyjhZxx5s2y+HoinxAQQSWvIqrzTyXutlLL+liqhXrPd
QcCrzenhfDOE31cK8hUuV/+p7whMJlBlKJccz6HqASpL5CM/Cp0aNuSI81CJG2gC
7hV3x1fS0ws8ul8w11hBEYsTFkD86WilNu3PA1UgWAPwz0SmyJ+nL0aW+wVBaYZQ
sg1Ygvd/C4B6BwU+XZBZNabv8hf0C5pRYI2kOjWjFty6xlVHi7kq8DK9JXbWwb6l
0hB3WswwidKliRUOIh5lX5ThB3KB+h5ABftgyt7cxZRLAuEuLJW5kQslY4eS39mj
TBZJOX4zBo9PU65s6qAgEr4CObvhJTK6DOnDNvSgC2sgXex165yxRISkn5y8p1m1
xUPQxBIeAJwpVNxjENx2mjKjbw2SOxj9oF56o6L8CWAXQvwtcPoadoNnISnXlxCB
drmpxgqGXygDx0OwGd+SRHa9Ahrw0U46lwzzZLkLD3P+ydMiOachiOHrvuhljOFG
6p8qgryXnuk3sBKoN9n/MyAyyRMCM9IsjwQrdIylrtBdzBXfLC7oOFOSxePLOwn3
gqiGeuwgcn+KsY6Sf+QQ4f8Nt99Bnf/OSHMNXfKH6FYRPHb7kIBS/FhOLdN1K/dG
oKm4PM5cxjX4AgJytkxauKIOeDdY61LVyTwY8JOK8mqsmzxTkUocWbPcmS+rjnci
gXZQaY+qpLuO4BWwq47SHnfpd6n65QfohP5iurBpy+GWgOIvzV/n4LXgtvAcuqRt
0yi/AuaGXst3oaImbV2kATJpKkRlEQxjGMQ8BtH3U+mWyBNcfcrvwrIAhIOEpkQn
16ly4UBC1T4gHyQpR7qM8LJhyF5/Lj3BROUUMv1FcqDfZ4m32X1Rg+YUQcM8sRgw
H02hjQNTGce2kTthFs3rJlHdqTpxZDoVqIpMMZE8YFOapSYgwpszEDsM6tM6Y9Yk
Fe5A7/Vu9Y2cIJ28bZq2Q8tGrtIoLq1KHi5V8rlTVzXoRy/n2nXySlaJNyY/wFcB
V8k68AS8EE8KUvn/v4Z/y8pM0koXeB9sKIdGYyKPcTiyZY7h8gieby2KZ1TFFDDi
ksBNMKAeXRf0mMPVpPYx++Oxu6Djhnc3Awjii2xBkHDZB8DDzA8zKZGtYIZx17m1
gXshv15fspNvfnijcmgKhTCf8q2E5Q2iu39mF7FMcJAiNIDDkA86VtlQ0Ndl2iO1
XVEeFyitUGuZXh9yNRjIdSDP+WUSE+OZQEgYnQdGfJDbzZl4DkzRu/ONfJaJvFTk
y3fPi/eVS7BTc4HKVsy6itrQNgNGxk46Ava47RMKtccb5S0fx9Ooj1xjRMQT0SY8
jUH6nuzZvKWB6arJDjXonpZR6Dx7ZPUFbXTEwmDq9J2hbSUwTW/SoAbNngh2MXx2
VwWOkUpCWlxBIsVHGYg/0RZJXcMkrngUF4j96L+Zec9E7tqdp9vJ1jec0WGyIrY7
hs+ovTu1/TNcHEgbpCGlxlpce3RMmJU31HaG+2V8kJPbpc+qj/JCrjhAu+duH7Ka
/PVtDeAfQslxQvLgnHn1+KdaGlrAbhjAK6jSnhIUv7ZCzLW9kWLW7wWwKLoEOe9L
ZUBmsrGSIhHJe/K49/LP3OOOaD/GQKqeF0VsuNg1AVZUzWMKbo2MQMrRjLo+YRjI
9Xo1Xw2rdSfSSmj47eFKFNWL2xd30BFVvbKn46Wbb9S31EVEzsJYTLE0dZqW65Zu
1+B5lQZ3RQ2FpH887oyqn2LAXdbJRZigx1vzM1iN5YaBZro65Hfo8djJeoR5dt9e
SP8EXe02rzVsHLMbZtuVoflq+dUicSe1uh+Hu6EQ3y3eMMQ8W0iBUYpIT6NjKFwB
3MrgyQ3CHO1B8wK5A5Hz1y7pT0K+4rdDjh/JpVh+H3SoRt696e061ztcx003RxBu
DEp7pgP0QNSaNJxA7IpYfqDctQfRT3oCWohImNuCVjHEDMNXwZ6z9MYxhvzlPofW
g1K+VwPiXMgOVAlRyLg1HC47SJNBIgR9LQG5XF63zDQvQUBG67m36sBsAKz1x2dx
MvADKJI/Ks1KOWWvU49OcYbGPAmXbgR/E93evwToD9NaClMc5q6N99akbDzhQZRD
58pdiJ3Hjd+nTn+IsZIJCK6M5eRlQxhjY8Pp3Ntht5sawsUcVREXM0ULccJVKxoy
UYSoAjoYUsfrIFvUXHMBby+aEOg/qjWbDh2KQrQS6P2egAqsI4lMcacaVPW+V9h8
fPe36Skbwx++FfW8ouJQWDqnsODNmjJup19b8mpMdbaRsqst6+OEbS8Mq3svc/4f
nblVJ8bLtJJsitqPmcwLdzAZBySWSXVne21T7rTlXWaPZXfwUnBp91usWa0EbDmj
4nFFCT2vItYsPzm81MA3qsIJ5BfQxcc0VT55IKlXCLtFX/4QpH8hTVyvZQe/Wep7
OJIN1y9IAou9MMzRcYBt6zDv7Z17qpoPJap/F/cGAveFefdCFbpgQ8jfq+/oKGaJ
rExWBDN5dPO5sFvrDwVm55aoGqWHfss9Yhw/7CbY6xyFNibeCZ1ZmsoKJ5FpGFbI
ZnfE/wRq8mukoidl2fwhH0O2MQ9aTutZMvoGElRfC6xYEAGrQKWlU3xaMjXTm5VS
MiHSwHGwZaIE5fHd5qAIC+zU+k4gBgXYWNjNKDk9pe/fqXk1k6RRnFldqpNbyiLI
tuAJjKJL+GEVkPqjE4n0hsNbhqG/MOIlp6AZKEKVZaiYgyBOe6n54gTd45Rt2Vzp
BQzffAn8ZIny+f2+dBiuF9kkZGLiQ8Glhyug+dii5zhSaeXZ5fWIVTqr/2tp1Wfg
P1RDx9rTVimkYTZDJZiU1KSNDfEeYlgwIhOraxbaQRt7ZAfJQGAEM3IjpyokErlr
OS1ndVqM3ktDL4y8RPVj8EYKg+KW7NRqlf1bzx+uIrSMmBJF4umrmN2DK/f8r4gZ
Vhx6JOPX3U/Cmzo1g1Xg3CaIXJjc18C3zTfw4SMSEu0VHs7NHX7xS3UXqt9BW8z+
+tWl53cs42JUhcgHnVfpR6P1HwBLHBlGS9dBbf1CSBp3htc+uOG+01W2nMEBX1MQ
ybX6jWYNS5pWeRdWB1FHUWNRxkKeEiND6t6c0ezozLLk6ZD/TCV2qK7gtF1CfX/G
GdzBtL6+JpQYIDm7UPyvswOjXy/LbVnm9KZxsRRKNRBscqacy2gETjwOQ5kXWqY0
wdWU9ZnWDLjKmdTcte44ETc66Tq43Sjdp4OU6uiN75V9YpBX2YgiN/khmZm0tuaJ
o2MZFVuJmi8cAvb5eUEJU4YF2ZFkr8sh2zsPgj8XkrxRxwxbnv08BE23fkMHoJz9
Rfka0kLpvHoe75Ci2vG6t9JPXeM/yQwfOiG5Nfm1fzk8V3pNY+P1QTXcS6Rg9U/h
rNxBHhBY6o5JT0w7oV5JaE3dZNbysQnuoi+n6I5g9EzNl/NIRJWVTxnktEzxpfRw
qhUBrO7NEUYC2UgVVaDXSbH3WHODBLpYt0/4oBm3pypKVyAcpRAW1tYSla0/9n5O
wtTIVBkesFK8MgiADf7RilkwdeLzzX4Rf5zJYlc/g9FeWxbFfDJ3MUhMuLelzddb
2N8HdXvpn6rI9bbSM2sPQTBYGvLQ+VsB5FqktoWtqJ+26j3ow7E/CRxffMNts8SL
vqp5ob6/ICDewFxwfdN1X0iyTf37npgJHddbSwEhNPUi2oEQPOb2XaEnjVGEz5vp
6cnd8lhVli27KFU8X5UGeHOd77w9emfxXokCAiRp8kjKw0xhTcdKnOwXonusQQOP
7y8DBNyuJpyz4pKVpN8PJn4BGgMzi41AQNEqxwvEYaaQi+DKSxs1qGajAIZFGVJV
kMWitHQgOkFYph0KGUy8vNl/LppBbz1veUVXzPYYpRAMon8jao5yOo1oAeDb+qMd
w15B8NWIza009IsgR8b/q12Uz1wdU39uqYQtgVdbm8RR9Dx3qGrAFLjl8FCxS2xx
eOPLer6pBmuqI5BmImZkRohg0bnMVpW45FNeFn0/x9tDjGgXweqwEUBm+MWGdBz8
j3Z5Nfv2bj1XkoGK43lcX1q1jK61eTbnd30QwXLe1c/fyu3ykWa7/QqjEjMaM03e
Go3qll+2c8hndQ+cN9upxq7eXkEB5WjmBoHKOAUWkqMiw1F4Z/uVd1hhsEvvUQ8+
d/rCIiuBryhoIs7GXixWaB1ryZBGoPiihBh+YX3HtjytKM6T6HeTPicVqPxsqkfl
BSdgNa8tjep0ukzIanrr3LPI+f2uwg3P6jlsJ5dJ31fZ+SG7Tnb8jlBEkcx6rS+6
8e/NuBI+qjwl6qojeNNEmyv+vYtiDZeOvCLB8kQi5MyswrGvkefK8wZafjfo597s
9AiHl2ywP4kbF4f0UxyFeSjl5qxfS0GtnNYRxZDDT6F5J0XOSzfKiYw26csGqfLI
vDIUPwfd1KdYfqMse9h3YKUFlRqGmm399obdmdSkzeFo8KDiv328/rJv2M7opnKk
yp5ZUYT5ITYFAbnQzrrxamn5676f4HClGOHKR2I3pqQHCKJcol+pPmxvZvFOiol/
QS3EDRaXNWwFwolSoYKTpOuDeqVLve+T2m8Vt8JdhUgYbjN3FfFAvb2p8esQ23wL
shMAwL0ik5lo2DVKxzbfUTEIM6a7W9UeyGDqNqhn1Jr7H+ROQ6wnRXPzgHzCfB1a
PVj3uW5t9vY6yE9hPUoBJ0A+OpikX8pAei6wB517nJCLXf2schb7AtcUS1lY4okX
Ia2A9Q1AwIreJRRafB3iIQXY6GhZSwDMtNwVbDpWu6ZUvQeZTYLUn1U4/KBCifcV
f8HYD6TD1S+XfjLr6/emq3dFCt7cMEM95i+VDIar1+IX1Wj+JaDa1INVNHHlYEBG
B6001vOrujGISlGsTo55oSMMhw5jOAKmLb/rLJkgA73EkxNm6nzhFPtZ/g2c+zcH
w/hG0YylKQDesAhPJ4u+4HD2DZOaKWZmo4DOQw4UrrmtiDt3228ClV5PemwHKTDc
yIlBrUiTSDAL9XKdoj2GiyMN1y6U27xh+eSvRVCZt99hPTlQJsF3fC7hnEBhtHAR
pkdv2t76J17Zje5PUjc9h0tT0lzXLGFV2qbYS+mxl3SMyzsakCrokn1FYQfA7Jst
QwL6coynxlfErf92dTs4Xt/u3Hmry5iNsnLf92rEQjhqHOv0oqhKE/vLKDmYoqRT
H/yw/nGyYIDzAJcI4TKSC+2HEuFtjqLOPgPKfEF+5BsxCcp13/r21G3HzdMhKrHN
pNtgGpkc83ASrrIEeDObjMJ+ADtbR3C7LUkJEb3C2gSmUcGZwT/v9KxCMxrkB2c4
jPeJkMCV9SrzQ+IKQLo6HpYT8zEgbCkKlzcbun58zWikDgzW6+CSdwQn7k/v34Qb
lMJsD9DPeI2uHIybEv7Gj6hTilQIwpkMTH2/dn2MOLGjIEH1wTyp8yWLchr8nzUx
c/AngS0KyPnKqDFLCbuUC37aY05m1D6srhGNiLIoQUCJARofih4t4CNJqODAy0xJ
0n00gmvHw1c/5jZ6oNShn8ifQpnbVSTujjZUYBIyaESBLTUUYvwRao6tOdIXxBoz
UIDDmlOpm7vHrctjGpVw8554KrYTn8lDedl9kvrrD6LPQIAmTdWcX0sEH19pYqCI
P88SKqx6hbW/ffZJAldA/F9FL/tqkvmODSpQk3OrBG5pe5+k9yOHZY3g2sR+6AcE
zmPT9UQm0VKNiWl/wqoEUdZ1L4vqCZxvt/V8S1JMCayNsaP/xVb7/OPSicEoGpMn
7So7F8f7gKlCfVMmLK96YQZ/QntkF1Ax9A7bD2tHjGGTlbGbZMjoeqekZ3IBfizY
ur7FVnNAQ83BuEA5qbp+QLyrosS9eFK7SaH7ZfDwjuscjCklxhrrQgcmeAFs6EgK
fvKV3Fqd9TLf+zfH/xxySdwYOph93WYwRNkwrwx65XL6YwOa7UxqwmQenlL7o0LB
5jsiYyW9tBWwHeGPTmsDm0qMZtYSelhBVhCToUQmk8pEqBhmaIW7z9RQ4K2YIIEH
eNEtfTlthg32rROqPUWE2yk8UGTWbcRWhPF17zFZ2RjIYyBQIcvT70IcsXVkaCYo
nSgM2DrO5ybzwic8+ck6mHqJQeZ4XlbNG8T3M6mW8rLw3HZcfDg3wis2O8U+b0qQ
yPNO0ONroj91IkdIHxeL9cHcEf89FCtlcchrXtkUyy+zZuztWBMMTB24axoqc615
S4ZAZ7n/U+Ct5sqiTSMDsi5F0GCS1rw7+93AfoXU+8/KiATNniBfaMCNPpOJ3GML
ktl8ZNUkgy6CZ1slnUsT+eAtFmhnXsioOLIlE1R9y12QdPePsNaeEcL22qgZUUnV
v7rt8EudiID6CVKUScFKd+yzO6Nikl77GkIgIUlUa1nY1KgGllAAYLiwssRwas2Y
mFhCxWKN03+39/aUI7cN3+W5x1hWTvnmZrosRvucwFIvODmuBdJ7pP6/+OFPkPwW
vIotSqBEfMdUJeOzUq666gghZs9VRyKDNxIp0jxYDebRhv1hLnIoo1RNV/Q8JYix
+H3CR/iS7EVG2dlNR3AFRkS8qiv29hHkiAudH7yAxupcI//SIMKXJ4rG3V/3FghA
lBjoOsCv/C2itQTsSoCCV3oNpyA+oQEN8pK+9eRxsHXSScmK20MgzIJ61SYm6f/1
zByUL9yGy66Fub95klRRjPOtey4H21TKsq+62DEjGlAiJ7oGcA6Lvns882oP+3ow
7T0SIiExHdU37nx8j29jikaf+kJqazNS/VHPvYQ8IvxujKKN3ObrPO3fzeFpCbRS
AS7JZT0whcuGporXHM2UrY9o2SeEa74ESi6XUcrK0JK8iH7nrrFaUjig5HuB5UrB
kEnmrQWN1uE0AgRVAzXzxZvTIc98+5HxZCcDGe6zy9TRiTd1KiB4tfBVoTLLKjoL
16bt3vNNoijvctENMJ2HS8By4KO/btLze+pBKTMl/35ZlV4JTgZpl8EgQDJ0Bl9D
FZ1Bpi0FX22GXHPlIhBwcWmBtGbuw9BToJYRAGKU/HFgL6aHqHzzl7VB/J3oGGMp
+Qx7sD9zpN2D53y9RC7iQ3vPbn8l+DSyUO3piSaFaqS+EwgV+jNSXHAoejn5lSmQ
Ts1+hiUp2b+ic37vS9h0GdLkcWt+EG/p2LkPFN72Kn3ZAenmn/NNvzq85TVNKKhg
8C+HrVoTMD78lzASETE4wd4zll3O5KtypQIAae9vBnaMsonaXUtPKWcm1zMihuAG
2dEM81lQtFKrPTPxzCtBCcNRfhkZlN07JbdRomT2Pq9EDZtS1S+uQcv/fQGvE2ua
RZoceCc7Mt6/1Sc0XTSVvKKD92hpPj9C3ZKGpwl6isHBDbqnDoyOkKooKKzS8tjd
RQSGerQklA1Ukz1EC6+PJN+28hWQilfqPHJ/v8yUobnK97zvKoIYi7o25UDnr7gK
bTXPy9CfmHKtXTco2IskmBBEzkkBqPFgsNaf3eHTvJ0BPjFZOnB95ylLrT9USeUV
W9xUDNsJU23gGESBcNryyWc9kQumyISsasVmbacprAo7UzRVxJvtlAxpjRoMIp/l
jA0qkT86mfgODPrwJjf2Z++HFbONgEulqEy5sR2DwtG5ep1TU7ywbWY0L+/2wS4J
HJNOuOzI+re/IBw8M4uyiYzg96c6/2FCualm41AD8inq59uhGEBbKwGuwwQrH1PU
wH51E7TxRUOgx+Nyub+2GnWaGQ8KP0rBw29cz7FmzD/Ius8VwTAdFBZzp4R3n4NQ
ISDMx6jiTBdlXZG8zqbpxg3YRGHs2xU5/u/4a0ssu3g7sirOvi9/pDlZoym8ifzb
d7P9RG+xQOnmrP2OYaXNJISv7dBqMncXyWvvE4YgVsE9o0gSJMX/qdGgD9MXLwf0
t6gDjzaFM+DHVMiyImc5yspxPyj9wL2uSxazALXz6hOJv22NQiA7F+ypIEFmbRdB
XtHC5AUDe/N4+wuW8/O3/obRzxjrVKj88b6u/Q66TKIMRJNZwvJqRrWycbj4bYE5
4iSFzW+s0N4C3Ko3bj7gT161apWBPYB9whyEvSfLud/QU1nRkd7fAHOcMuVOS05M
pUmhnok1iGLJd8L9cxnWSpwUgoNxCJtTs6RdS4UcgYbYjlYHoQr8Yp1eAGOVUeB5
LwbECi0NqPpQvILE0S2expAhJ17YGhXihYRKBtIL70GbnXQcXdwGFuYgMsi2DXu+
1PkenIrvoY8gLGb/+dnbT4qScpkGLe0lA6Tc4mpx2f8COtuwrGj8NXR1XMPMeq1l
bk4aHtHFreg5tOqp6lnDrVo0cKAdPNtoM8b1fb4efUl7Pm26OqY4IRX20CRMxM6p
7xgQII1XTQPheLcmDdEknzhjx1kILROQk0INLLpyI5AGXcnd/Ds6sNccHM7c8pNQ
wQz0fkauD+qG376UyhIJY1QOi4B9j82pZqb81Jku7/6AQDfn62qxXIGObcFqaPyF
cEDFROOpk+QoanFH4zBr2vS00qywZhxZ0PFYgn24aI1ju7QD7J7C6jiigZNzLcZL
eMWyRa/BXCMQ4B1KmkFoAMwUIwMatj/zeOwVjTlc05VAZiHSyWtlzCMTLOEYY2cA
IjaL7NrZO/WE9K4IQIHxCg2HUX3OcNZ4pceZlKtStvAYulyWTms6vAndh6XUlAYO
QdjrQOYqGsIRRv1T/q+pz1pSGoTNwAe4Ac1zb72fienoifKhsvkWoSAwMZx3cPjV
nTUoBKY4P+93gbUeGbsVpRuQUZYRDSB7lTz8ltOdWVJ0bljGNk9EyjrFvuBz8iNB
Q+5wRQZprkzdH8bL+gW9KeQHt2tEBlhRA2ejAOBFLsMrV9mrf1bzSZxKk9nBL7/e
3B1GZ93kr4LukwDk75SY/RBCqSLN87aU3f0s01W1tgE78h2EYl9ESRkP90zUbDGR
rhuAcovic+4HDwnewVzEX/fi7sFlLoa5VmGyJduaM1xOnwBOm83XJDz2ejrfbbkx
kt8o3nSIjF5bAYH5Qz6jgtzXbeC34Hc2eK2qZ0UHHVF0cWkTmjdFPQT/ZWRuGmn8
C/R8R+agyb67HFuCI7AuVPAHxGprN5tUO48ccDu4CSwENMO0TAGXDKpNVq+hLeGM
/OEey6iiCl2+GoR/rr0IXTJhs8D3RRP4cbwiZ4FzEP+uzBhZDP9ZcWhTZ8rDb18v
/sPhqMY+VN5dkZPba9McXFJF59XIG5Q+yVDI0dExsPfUzoFk23QQjY/NzLllHFFc
iqZge6D5rCbbxMgx0UlasQSGLQ1mZgJ72Js/AJHb2Nhs657Qo2Iw3LZTZHeD9xlQ
RLPJzr3jnMVp3kdS6uIlUIfCPV0rIJSbdZF8qrHAWJF2Gy9S+2iL5Nr6FCRfGXjD
l3BLOYHSfRPRBR2U1fzLZWG98/tSQAvxMZ0jTHtXzjOZIiSrZX9GN/pkKYVuQ5pW
epwIhAG+CIgISeJMXX1O9XolGhzwcYhACOEpHUMORaLr6RgLYIR0nXSjnT4J8mmw
T3QQe1FEsTnLW5cEOCjRdWs0Wyun2vWUAf/2w2rC2LhIqWSaIBaTRg1vLCMy+Hu1
EvykhanaMeVNFRoTedQiWxtnNsyT0kVzFCuRokStpVrkzRc7JG/kxHoui0DDlXx3
RIEFbLfON7DmDbtwUUWn/ud+UEeuwVwZXihRD6Z5r7Qqkklxum+0brprTirIbQch
Tw13v+KUzyLaa/b3vSIozcMbWVXah07F9GfRM8ZencvXXZQLeAMyrewzzB3rCrfp
SIyiX/v6HMVE5YRgj/AKY8AwV8aJ410pufwrtXPeQqt/sSnQibbHUVgoneHOjhmD
MYftJQyByljfsd0Hdx7tmFD+48F/pideIn/c4GAhhQIcqblpZ5QQxS6BF+J2vn8j
hp9ngATn0EXHqNaoYC+RxBcVP69YWOggiDqUrdsADZ1eqE1e/YS389wcI5pocPRm
rnmcprSg1F9B6OydcLQqnjLLtNh+ey9NY5O9ZDqhNIGJIB44RVUW8/FrHYB0afs4
j1NVohPpHRIlCystcQcx2esAIJoRqvuC7N54fak7y7nFWxsMC5dPvLJ+VhwQKaIT
kv0LG09Xc0a0FJssogd7xi+n3Wk2neShniAc9S5ASdced54AXOpgYr5caU5lCXWy
qSFAHHziRGdNMU6dduYfQ4MH+OEIYx9SNtTka9q2MPPx/Ia7OPpCAXjXW3wr2pH0
v3yKqKVxrGhWIOBGzShWVmXuHiHKSHBpveIT6ODpgLy5eAtiOpuohwXmMXXuv+GW
6x/6FMtnozBhAuvkiYnGUQZmFrwP2jjtLRHuyQNidHemMajV2s+gbPJZm4houNow
hE4keZ4TFRt0OL9qKb+uiOyqkjGsUWpqj/PB97uhKXySrAi82NaFmo99TuN3hYPR
gTW1Qny7k0mn+FJHUEsJ29+kKs4654l3+V4+vPvI4OeuxYr/A0s/appGKih1DDbH
krW8aKWM4mPNuB9qXDn8f7Vi6bFRsGJJte58JFtmTVHtNqNK5RyH9mtW0mPupeXo
2JXPZrXGW+EwNvucFkOVzjziWbRV+0Kz9zHZv9AKPUQnwGwANHOdCQXDSdj9MLNz
xhslZWF0F6sxAr+FLz0ZrMUpYx/uWmGqxcn4tDBKdAOvmBZp7wHWEohdgA2w+LEb
UYK/jRHgS4g0vYc2k4VRPDFKMgBlve4lehpjCRYDB10aJgiw2qtJlDdza0QroPUf
CHWjSPTDQocT2kNDqCtehUVdW823p2eGKXRJbfIEocMYyXWvHdPSxuiWBQcnvLS9
M1YHfbAuHwRoj5PZqEESgD2zxbDmb1jVkwzZxWEjORQ9+vCc3GxdPtiZlbb43Pqt
ZxUZmgTERhD8QV2dcBhbFHAQTVbHKp32FN0pt0p1BvUdjJ7FDqutWgdE7kvJHFgT
p6nKmTpxfYVx1gOgB5Fi+UxPRVswP18ShcgCdhAbj+vVsOQZ07+p2cVOk/UAAkzS
OH0U6kgVH8bsj/bjPDw+twZKeeMhOxr8TYpNisS6RqUV7UcVaQYKU7g0iS+sdCMH
OXd/cAsxtB6F+2VkgLGuu2GTfTalwu20+CI2pk0hdTJiDwFNJhLxuZGDPbwSGa07
GiYM78g7PaGd+GfShgTSKrNDA03WQjXr78/pVoAE1mRHyBZxrZNrtz86fbkPPc6O
IKegisBgl0O7Ijx40RanUPLckimTw6QxXxv7wdnTjPg8oIyAuPwhjJBpvRDJBOJt
winZ5W/w4PhA2GpdQGNbvkplFYdDwBaTESD8MH9OdTA3dMemuxbYOFRnS6oVaFNM
KXtqgmkyXkrFpvInu6IUdcqBFhcM9QqAqZQHfBieRCCypCzBvRVftKJ6TL3jKihF
tQBjd8YL63iMVGz+L8RDRZpTQGXdYifocH74rvBORQksv0NQZnSVM94hq7HcNAjC
XbgpxzgjoUy0tPsXoBQAmRVlPRA5PRWms/MpbCVmAw13Ci8qnLuoqlzYdm/rJrbk
UcAH/Fa0vetom38mMOfJsxU8sZx6xOt7rGYt2TYDZInhMXkk2fI6DCjD2DfRcHZR
4g4x5/Y3W4luR+kOLrEU/eBZ40m7JkECScXFnxY+6nq9hUq23jpV2lZLUnvDdAYd
UCw8lACCKcjTdmVo1E6x6Z2NaDJFhCFZ1vS21xT0SlIP2S9K5XBCK2ShsKx3T7by
l7R2qLjfNGE2RRV+gqLqOPT58Ri4qRvxg2b+8Qgvd7okdZJ2RClPeEWsHATXHen2
oiozax7ALBRKbsZwyvP6ykYCdiAP0ZyoGVmvFL+W+6ziemSqFiNSatIax8oRdrNi
1PteNpsktiB0szgFl+7aN4ZD7Ix2UMsfReb45szWcdz2aJMYcEPHHxhd4XR5zJfW
sL1Zqo484URfdaaNHMb4XnQxD3mUphlgVWLMXup4uA1Ovpn499cpoXJh9QfR1qfx
DYNDaF5CE6rzprD+ZbW+XXHhNVAgnchKfZCyzdC0HW6sJgdCw4KYruQi2miGZPXR
wBT8H627Z9wetyYHbyprJ8NouY/TqLy4JRVJoJZSsyZpqrKSGH5i/jfv9jCm6bgq
ZdedF3v/W1SKFeZ00SFC8co1cy2D9D1YIUMjrUDFMyvogVBtaWMkmH2loUepu33A
aJP9pHtnjHs3W1Adad9TuJ7l8EF/byjGLUifhLD+gpd/4KXbcOyg8eQy52dc+fsm
0N1ATzY5mTiF5yoZk8BsPzJLfYdLGXCu9F9o1rkC6noI00ZwI9dRoihbbH33FRZP
UjedcgS3lfG9arP2QYX/6KUb61UMXO69AVQjchSAVqHSqirC9/hfd4m7dmkv6sP9
nhkYeGK20dFKTBE9G2fuix9q0ghwISpcnGk59kfUTSMPQm8DXlWL0JkqcM7CjWAP
E4kUYbylzvNhqmaMCVaIFG2iM966bZd7okHa0xJzutTirXJB3/6o4JxzuitlcaP3
ddKgivtfjGYLVSHGhDS0xEFgcZSZ7EQQHf4MWvtPYpA1YmDDDHr5R0i6MDhUSMnL
NEdzJeTxBi3x8LzoYg5YZdn5VvoAGN1+iN8KMHd96Iiv0OsxJRcgjIM06xgAsQPN
aODA06wAJfbrBWTplDhCda3kvwm/1ykj2bvtXUO/cIvA8H61adAHuEIZh5wwomVn
kRHY10Szvu1UDm9ofdnp+y9/tW3QpjFRmX0M3JaD0g24PE1mwuhk9pr8Thn6Loqx
CUmQlJPUEGkjjCSvLeLEPX7v/lkzt2DagSm9xNtSn+a4vJ0NDRVcGjSgv58mbs1l
b8+SSxp2ZXKdUm7q1VdmfoZdlIwa+3qKNrFo5IQ/gtSpdezNEx5aeOmBx24JeBlN
AjRihS99IOpnUb+nenVBaHw1fMD/geoExd84o18OBs5GQCEANlpfhkLPvCKuBtD4
f6v3X/pEPjQGvrnWAKTB9nqpS7WFkHdIdMu9vHLE7C3+YC9sBEFWbkcWf3fQoQPh
X60hXmThVPb5eOzu2RL1v/qrwUOsCmtmFqnpjhemqq4PTKMFzCGqf+TyAZJVdP2x
BlC0khZn7c7vuzLBp9BjRu8DeAduKKeCoJN5yewnNy55lQhyzh0CVMFZ2r2FUDC6
S5nQiYdFmCh0jt/TnC0+1U3w/w5AQpIPm+NpkIH34WAIPOxX13fSvQTVugQLybc6
9gSBWfL7gW4gRQFo8g4asnbt2KfWCWV54TFFIH5T2/aKKBiGreD37FKgQt8O5MfZ
8jWTi4+tAU9veEgMPyXjav8vH3xmsBlkh932c6RKOi3PP21OQF85DxAek2oU1LAy
irFOC/mHWOW4NgxrPhqSRu7Ds8/xuNWQoF0vTY7cqfXJZa8QzImQ5r8U3xbMt2LL
lEPlbdqoGgGTkG0+3eufXLacAnvB09+hamiPeSQsdZEh8aSz8YYmTcY+FAjmS/qu
Dt9ckhOVljvH7GbsIWF1PJZV6SxF2qRK2HdEHWlDfsfg0h9HxXYmeKLE3/+LIEph
81woHuDvfwLB49cDTt5NBj7EED30oMxBogh1Y7oCxGhcMSzl0yXVHtAAap4tRB0X
fWFali2nUwBkNcT0oLPe3DlfNMrjZtaipYfNS2IgIFeRQ4jzIs9+kIoO2YDzWZGe
zeRfaKKYxCTiPwiamgjkdLSedFJUpWnGPWYurLVSd4Dfmwv3btrEYPe9DLXF7Vrj
F5OhCeZUy08/Du+sVJlFmor0YFieBCZUH3sGBDTJn62vgzUPOtB75EXWQHUTaYZo
Feg2gbPiME9g96P52sCpoL3hbfHjrzSHsDpQNf7ypL2RyLYCgpTaA0VAp5MMmAi1
FNYG7fIJ3Kmbv5INmayfpayAd+FihKN5nlqX0AcC91Mbktw6FUPR9rMKPIHMnBRM
u9HKkuIO2fKln1F6o0EEOkLmYn1nNxikcC5Q9wj5ZslNZ4cOjcJKfkTFlwkzGJn8
CAfnZXTxWQ1qAN23lUfL8CDmO+qb5wd5eEikAOkXa8bk85g3fHmMYPyQthGD1zR+
YmZKdeBqoE0OdPykbF3yGQ8KEpS6qclizQoloQjfd3GlS35cfOeb6x8YCasdivVu
D3JjdartHPQ1xhXhExkzQH3o2tgcTEfP0DL7QcbDSgHpyx9+8ATpPhl4Y8wYVKQ0
dREdaG8NaNirWF+Y1lC2qi3NWeXiguhU+Nza8MunpswI4G/MX530P6UmAQ+pwzkK
g9ntJ01bobfu3fZToVBp6/0UGO+C/0t/ZKi0tszyeL2oRYGoiUgPnl1E3S9WUUDU
P1+2LCJU5OlyRRLvWnPTcUjJdSJoI7XVht1Mgz/l8u5BHnPgZBqz//UAyZPfN/hR
9MV/K7VuxcEN2xNTDpXHJUhYRvD+0RmTTGFrxBBt12iXrlGpCFrAU3Yh+o/ytMb1
q7c4Xb5pdD9QiqB2YYZoCl+kARUxZQwrA7e6ebQyJgAMYqGCWATSHK0APGQ6VsUV
7CbSxb96LNY1TOhxHLOssfG87ZZzGMTA8Q/1UN9+rZogQR+3WyHIp4Y0Tq8i/QhU
M7ULkiG4iJwMTDPdH3yZ+qRdAJdRn4KXYndBY/f8DpYXYJ0B6fv0rAtqB50GBfP7
4/e9odkriDxrdrxZRB0DNlMDKdravoXv4Kx9crdJPfIqBeJx33FOFFY7LpaKD0TD
QWR26HhMGcWz8Y3L78MmWNfiYzli+i369YpwO8py/i/BogacLMpjpcq651pBS+BH
qpMefVpxJTkeu08v3WJwIeReTQI8jICu9gJMAfWcTR/cPTqnbRy4psgrucPS8aJZ
azQgclr004pV0AtyRJPjo/MhgK6kzrnNLvTMN6Z2ibBNHM1+Tg+o6oHXxokvD9bZ
JRjMC15asIjTmugCTZswttRiNZbl3Rb8KrcV4lQKmdkgxppD96bF+HR92ln38Uj4
slSBCRlatccDuxdZPj0V+iH1BgZTcuTt8cF+XcitlabjLsnyId/WKsdG8ffstNBJ
llPAyHOnd/AbY+lWLKV0PLJQwFcUaACZjMHDiAPwCiqLUtJE5BA3KqgmfqE2fbhK
6AV5o4BlWwBiUQe/wyNYJdRGW4q1vim8ZvNvSXvvQd9yc1gs3/UNnznU10Xf+Yxg
i/ioEKMIdklC2A9FZTi/Ybw6Oych4gByeg3lYm4so/KSlWNxn3JQO9sF89kmVNji
rSil+OL2b5j3srdhs0iMqEeWEzcfbhUhnnswu406Kvahx0wNXpZGXh67ewR06oFI
4yh/lLx1K5jPG26+I6fcXRvCmhUJlURkf6WFGOvqRUzQrASiTLjP74nm8XR3im+r
2jdBygr11qm/NJLYx0LLmFDYVXHbNxv/Ce4KgwnbDLFiMGnCjcIl/v9YPR1cMPBp
vdNNAJvF3sj8Vs8DqfaWf3MZYjC5Hzh4qqgxWX4l3yRqVLapqt/8uLWKHyWwnoiT
v4IDete6zXJoe+8bJtcLQWa0MgTCaL7DOypGskO529oteDGKVKPr6U6mOAdhS0qw
LLZzgZFlnMJqfctOX5Bej4qQ+gKnv/0mxoAnFCSYQnc5Al75KS97h40z3H7dkKWx
3YbPVZ9+rMW8LKLGYhFEQxOvW4OookzSVQTj37bATXNZS9TYDzUsFudrqvSidqr0
jzAUYvvKtTFv/wfqYfNhcejWXPRFjGfAeL1RDqEPd0bUHBCvEEB9G0BmzbAUCAcE
BYS6GkwlZqH3gTQAciNl7ev59exq59p5tQJzNhrDX/iblFiNa9RaY+Akxq/jHE5N
SWi33dteT5kttUfnAGuJGjTPIMZXGo2QS6KoHeCklGh0zXWV7BjP6AEaq2R7OJNq
yibFCV8ia6K4ymWE4LKN6qJuTxfYuD+bt6cOeTw5K2+0bQIzFVjS+AQDPLA9TF+3
mTctfLC7DTrtS0knBTfqd+fbsD5qHRbNg9u4/WoZz5OML7H0MjTN3Jlh6n3V0EX/
wBR9o+NueaDjCfxS/gkFYckHLMvNgMbdjX6GPxf6Rur8vFMLP3AMpbrf5Aw2VZEe
1ib0ytGda/25LuRyGr9AzxZ6tvfdTlqqygIGsrFq2cY/8XWSWQAqfyUy0NytWiHt
/F29T8piKVBx7rG2zAmixI7EFkmpLMNP9HkpSrkMbTgptl5Cg6IlksgXiy2OPpCQ
ZHD9n+PqxbhBjPLISY577ZIuYxbYdfT8b0rH7q2vhERVXSTZCsUOqw/QGV+60QsI
TLL40+XmKUAi58EGdi8Nxw36O8p4OeehGCgDEEhv9q46jvUYhqIQwKVxdTTPjCej
sED3B/EpnesNezN9XvgQ8PwhUeBkWCww4Fz+DwznTxmzbP7lzFwtqyd13WQ+ahQG
LmaT2WxbCECXP/aypPDq8sx/fGIjBlmBVL5JAQIiYae7Yowo/orpoZVcdNvjF+54
k7MfE11JRXzZBC8O9WNMef4NQBg3GrXaajJemluxchL6kRr5ZZFFO3KhRhRQodK4
qDwt/Q50uw8QB79gUJiznk5Cgwa+oBGigi1bqz4TIeWV28SEx2WazIfWR0yFXnkV
K/dflPWf4ULnAYgSLSWfzcK7+8ZnvvvX29jdMjOJhzmuADSrop33mLEyD+wt0Oho
JyrvtuS3OmrAWiJdW443ZI4xvJMQHQqFKacPxLbF+mYAwipFC2hIyHIdHX8dwX6+
d/tbuG1Dihu7K9aHR3NmYHP3J6FDXEYKSj3D4nSkge77RdfU1Cdu8ACtnGiUwj5e
YEMmgqxD6ShVl4URpOg4CeWd0a3imftudyvfux4GSxmsBThhItr2Ug5Kuf+YYAB9
IrhwrKjLcni0KqNPswu33reDUCwKiSNPmLJ7het7GQbNTKQSv/qUyXtju05DYvmz
SOXlMaz+AnFMnGol/zkc2g5GCpeuSPtDsIQYTVo6Dam4+ewDpvmsd+lgpxhpZwhz
9XI3ZIQzyCvF21oDwaM5l8idIM8fQr3IWnxvgGKnGCPr8SYAcwBuFsXydc1rTRxe
znmef0d7np2PATy3o3h3evIEKHwYIkUvHvXBuR8N29ik2+YPPaLlLg4nwJ9Btrkt
FSvc88CK5kd413Goq6w5tFF2juxNhTSKuVqA20jdD0axG+buvVHHg/7uwRYAECTa
pz6CaaLZ8GiZrHFYM5cGuFxPa8YYPgohA2V9H6hbKtYnuY5m10DTQ0iLj8b12wy0
mqQfMVzl2VDXcAueuj1WyzQFikJsn6rXnxpAz48DKSnqxV9eim+YybmOmqtsmhgP
bXSPX/4Po219EV5sQ6DIMvTx14BClhkR8iuFKTCjB8QdD5/Znm+jZEQmIwEnDI6S
ECeVjMiW7gcDCh40WyR6dtuA6j8vLIrhyPOpLakxfs+FyhgyFprosYHSgwSTU5qX
A7WxuSjL1PkZJdTkR4RqQM+rHzz5cH7TNgPdxuePNZ1qoPcQybYbse2vDgAdxvT4
dzXAfSokrnCISkUOylhjYEuaB89VzWjV1xaOH/a/YHlzIuv+veJu4Rlw4f4vJIWT
dGTxuu4gcBI6cQ3pDchQKEXhFMigKIZ0H2h8D7zW9QENIzZ9ECRVuSYltOQ/Eju4
TbQutpfMOQTmFhrIPnGI2t1tdHkEv6gRVZnt5WA51i/EGvDwknJzzJToQtJCXuAM
2j0Ef8wSIS3tD0ltA2t96n4DTf7tksqrNuYhDgd23u3OqqZavuZsYNs0woq0AIX3
suJRw3zSZ20LdllAojWuCB1l4n3qyQsE/35MT9SQQFBd7zghswa/lT/PNoXqeA4+
NyYWPgbZ/bEIvVLTc7xK4jtT+hPB0RbW3iEgymvUM7sBIDF9OFxJi3G7Rw0hGYzG
hB3RHFo++eyMc/ROGci+Z9xwgXX3pex4kiAQsOFNOSh5qPY68cquprz4ocPgx/5I
PX27+hvQdOSchuWaFjJh+Z5x/IF68DUqtdTswriSOCDMjnw8awCnaTUEgcR/QW3d
K5sqwXaweiVRfVgA1nqKQ+4k0LO0NGO9sMH1Fb0jw+ykrRVmP/CCsl9BsxvAqDAu
5FzLmiDCxJDfOgurs0lFYKyeEbHVPZRTAittgzV04Gq8mugMPtl//4ubaPPJltiy
cf4bvarUefm/STxay8bULcKFJz+yd3dijNbGlN1D9zVDfZrMih//onwpFofVijBa
u3MDioXbGQhWswJcVLpaFdDLVNt0tD1oA/fsi4dTLva1qfqzLAz0eOL5AdjZg9Jm
yyIsCBGFLoAMINjxerD6PC/tdef+jzSs0ikJaoow86evt6fSF/5yYFXAQPzo2TtL
D1P+yS04SO+w6UaXVdnykehrkPOlqWiBDRjb3J6wwBJgVdSqJVErOKMxRXrJmCUK
dZJ2GGAp9oOdOlig0GjBGzvh5EOJxJofX9Y21IvlYjX6qorots8ECtQDWypzrJOX
rcXRKWflflCVE1H5RoNVd8KU/UwJn9GDIhXzUWrDYbCkZ+tW6KDXTfcbwz4Y6Phf
PWKvj1UEE7UiKbUDcC1dbvv++SLx6BC7NOQr0M2j23T529sEmd6CkAkiHQipAUpA
T9tz/w7fmRqU6yGEGmz2A8P05ahTETECp8zbSV0kkuu41DmX0fMhoplnAQszsrb6
MYr7eCCs3OfnPaubPANL0EIY7c8ycjda5gKbqp9ibAorf7rqoLtAZ+L4b+Md1LfH
UYzwVtIKnp6lI98zT1csilkN5qS5HMqdMDNqDaH4WpwqlQNwshYe69V4fWdU0f9q
e6ppGoXhP0Yr214R3FMYbqhBOhBA1rJcUtUQkeWoirM7RzN09/SXiV9FZ7xBuISg
EHaFHY1SRQ9TbVTLmKYD9uYmkW0jUnb3Nhw5DnAs5+Hf9ccJCfRkmYmagh25qQwh
db5vA3Mo+u1EUNtCVO3WQas1HFnI1fttRZWAATT0LT1RROYD1NEEARhq57+5DoNb
zisu4or/Tl1ynzkf4eNOls/gtnKprSKsyrmgqmbRgeaLYibJNMb1p0GjuNYD3ayn
UBOPoU95D/L9E80l/hRBip0ZVztt+9UFIk8ARIcqanWJ7scZE8a/qXrRGn+zYmTA
iytOGRJvXiWgM0SvpuRjsE6GwwR4c/ZeuG/YWp+WNV3Ml7aEObA9EC2ZYti5SINU
+6Nw+aPv51x0I06qVADtypfy7y+jWTOBH39Zh6avAum5PvDtx+IvL5cuLGLewyCS
KS2/RpImO9ZR8/iiBuFgkfM4Q54O6C7ct5R1bRH4c1aDd+BJ/WSSr9ThrPYo6nGq
hnIBrOxvqRDMX30ejLhzSoAC8UfZqsbwdOeFFT27ugeOXZfXdFckelpOontlboZD
fs3VHTnH1FsOXM5yN1oKkWO/PD0hqUyo1xvlFpxRZp3C7Ck3UG5JpI2MEnDNVY+B
Xi+cXbDUueTODY4ndHGV87SJYvgh1cCs3WUPwQjhpO7YhXzH3ZZYqDY76D0lfBfv
az/s5d8S3VvztgDnvJ8He1q6k8n3DOmCi97W05aajzP7diZFBZYLCiy8mw/dewjo
0jdd+4susRMfnqWKJA6NMPwpKkcWiZJ9dM4vhCRDB3NnCnzU8qfVD+c44Xvk4V/3
dxcx1UBGztIbbHStKl+BkrWtzLkDpbmDwG7ekNhAGdleJmy0US6TmVzHyotdq0DE
o/lgGEn7uDvXRBFQtHBwQUMrHLP1OGo762G7X9ZYVJ1zcwQzwI80h/4E7M3xiaXU
vGMupN/1GXTPntXz2Iwt7WHqtUbGfFzY3nvWWacMEOAwUcJpYJzEgxEWcYIEcz3t
AQ1fpCURH/5pDGbM5iopZNbxxCgM02mYDbfBajw1IBe+dQJQDN8rbp6XehEJJltE
Egqzoe2wPT8N+bHfujXHnT9Cmv3ApDmAimESPxOzZnFwaHG/1b6fdb1A6PD6eg5z
wD+VXGvj6vkY2lW/s6DUrRfjmVZW2lCFt/hfoGAV9xnhkNvzPMiqp/wGvYj3bT63
/6jQH+E7Ep2UQCcZRWW5VolFRqeEqxbD3LDyKSHTniZ197tS+znCfOVXaYlz5E6v
z/2UmO7+4PFjZTQtmEniAmGVnX3GLecDquTPOc3FnGv3b8h0ztO5oyKufm52QAL3
7QiBSKMM6g2SSTf4ofXOZwbEns0FE9v8q9Z+4whsVdQ/mq4HvELkjuCPWgXyBTQe
fzQrJxUkhochKf1DIP6YZf5ZGH7qAvwnhxqAcdpPPFSClfOR9EiePKAqE8Ixsjvr
ZNYR1p0iQFhnHiFl6HeJvl54sK+6bx5iF9MLCNgIytvaloqjbZyztadQEEQUEFsd
Xan3Mcg3JHyxxysX7q/7xHXg0T5Z5XKVVyc4y0rwzrHTpNGyviLQJZP9G3U0NXa8
BnVLWuVi9HZAoDZz4SI4mrmXyWwXLAYnt2qateShOT7vLYa7DvHlNYa0IS5E9NAg
1Qki7rNACOXAUorBAB14fdPSWxh7NYcGGt5pv12zDnaqg94RBlA3TRuuk6Qox4t5
MJk876OhCdD9sk9BnfUtetGckiatyB+0rpe9iIOX2nspuomkihdJjcZkfvh52H9b
WGYiztE+w6xPErISPA67zU+4VtL7ror9CRZU1jUVBzvDyH+5Uei42ilW99SJPKGg
QmZc5sYwbk2F9SVdU4g48x8O79gtJvf0ese5tBX5FVunYSPMcbSFsnc6LZDX1bTj
KnXq96jbjGusoMBmxV3yFTCA2JnYq+lFT55AuCMhC4YKqCGOitVi8rO9Bk6Hf2lw
ILq8pwCI5Fls8ZEqWD6x2/oNF8Cay7JHTyhqmstQNDoGVK5I6IEdYHAJT50qfrtp
xZb3AVfdOWZoO9rx7ytQSv1GlRGuFFrpAjkC1oENmoAsaZL2VttMdi/UPZKKhdCm
6qcNBMChMEa1Qvrcl1STbYgRSUw1r/cMa+dAHZ32a5k4vnOn/B9A4WKtS4XGSVh0
WztfOzcU7TnR1KgasXkMU2Qb9FSaUYt1PorVzBKw/YUNbU1g0q1qaM/aDmApcSQV
MLO9V7kB3LIhXDG75c6IlleR2LQtXNXuo1BdNgQ+QepZAaoedb3IEYo0Ki0r0fHQ
CrgdPw3hntAU6b26G/VNuJpORzl8+HC0OxG32BOKYRU4uk3N0SEuVSoQ89w1bsse
2vANs49aG5pN1tuaDMJnh811ZuQ8J/fHTjORghxEhNWjGBzmwuj8NgCfykfedIXI
hs3VKX7gOu5nTWYSOhpyO0UKxSpvBADlH7nYbWAL2JzU0JOKGZEHNC58uOcX0c08
8J9SFz9mTHh0EFDC2KEqlRpZ4rvs5240zHebh4nUt3DYZOoa3EIKopzY1mY9V13I
vuyHpHJu+My8+i0tWSo3Elj9zZ1yFBUE7Njqp0U5LLJSpadeslYT56sCtQ8SkIwt
PcTRg1KJJwiACt5P3OcSkj9wW37hDZ8AZ/4WrfoL5LH4ET/+YwglAndBQK6WoWbp
1wSlfXNTyQMbKr6imrZh5W/Qj2K8B+VgwRDBurTcy6yKPxAPcClrGwNNjApCpF5k
2m+D533lyKwrG9DPurC/2mYLFpDOls/R/VM1Yt3iRM53mYpR/TwoTT49qI9/3ZwC
LaCEb32YTSc/oj3+0TN84+9E+njcrHGiMAy+id6djihu+65jx2YNNu1Zb2LYLuet
oj2yDoyIV5WCHe0IzjZLzja5qpk+YIS+NFhgCTxe5ZHjBm/GawyctnVcCacGL3gV
Fvbot2y1RA0wubujCMF+5vzo+7+M2jypLDhC4hvRCCyaYMp1Gd9XiOvV72g0J9Cn
JSJmvFNPdese08kB7L1LEPwuhQOnkC+1zQk+VV/oK65VnfKIq1j2BEF2X0zCjopQ
GONkzOPNYw7plzJv8eRKwGi9DhTSfzfslt33ddTH6M00e/ppaqD99u88ShlnrMQR
dQVSCIs1bUATfMjo5slLBZvc6jv/niECmppLK5pfp5oX3sSCFWNzh+4xl6ZQTiQn
/4yAs5fSCbmHyUwXpand8uvw4+Vh8B2hqFYjkS6Db0BsFnIU8+pUVYhJkoTpUQRd
GqSogvzvmsxueIWfgVpFauMJ2AX2XDBptH5+eF50yWoGOrnAX3iKQzpBhBtWIHRc
LInuH/vmZehLX2nr1JNZxhqCm1DRBzDHncOa9z9T90hi7IYKXqIETmtL2E/8dDo5
+sQMaxRkGhVKkySCRftRtehPW1CA8Y+MCn2kI88hjO/caKpEcXmuc4tvj+RTgVSG
Lz7bodglBaHAkarA8BOQw4eikgymgpTRQUgfqoGdFJX6iW8gfz9ghX37OlszGKGD
yQeVj6MfgCZJyWizKvqaWFyOllPvIaYreGL1eg5daSs=
`protect END_PROTECTED
