`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O7yZmPhfeam50a30YrGZbPvIadEw1+2yuQN9VrAJjqsPcJeq1/6RqpqjM5hH/Jke
40KJiBbOlDLGwVEvRf+1xzxk45Me+pZB5bFL7oWbtEaAFp0gXoYOKldDrjjQqAXh
GrB8uKXRbVI87GvQlcH1kzAyTk3NoRX0WmBwUFe7b9w6CBsRuLx/eHVm2BI2ujQD
gODrPqrLno8tooVrCsJXBKlJE8Tl+cOqvQ9nIbBRVgtYX8l5XcVlw8SAV6S6T0Sq
mkxXgSTGRvxm6H2CEHRpgvQ/ACSHYuR1WIyCc0LeSU/he9NkSD0Z3QZ9QoHxCyTH
7oq9BX8sA/igWpsjdWgTkAHy2/AecisXAmGV4tbzqb6CctSyXNXp+lIu5sY4dwSM
KADcMlOg+cVbxjkEwkbDRaAUCJL8aS8tUIEB5s0Bm2U47NuMZuTAnDm+Sw0YC7yX
USluI6kvCFj36lpqMmRAXwC6aizGREA16Haxq5a3/gPfUfmB8QMatfvOcpC07wr7
IncxB98y9ot7qeVJcBF19PBAmKxO9C/JkaNozoIzNBhuibCMvEc7T+mpMi1J9zIK
kt9kNNKu80ALG2CMLaqpM2XKxbp83ewYuw9FaqrZfadGJLDnmH8bpJdkkn8SFHbc
o7GEITxqe/15vpjgSuDpAvy4DZB6kE9HGJBS9aq/kp459iPj7sLE48EsZTnzTm22
PQnm/K5G73JilZL81jzBDwFn6vocaD8jJu07PMkYV/XNgc04yMSVy7pKAQXaQFmT
FhriG7mWYxTAWkvS0bnjY4h1BDzNYZvkhqMI3sqOj7g3hAxCnDorktqB3Y5jxmh3
D/Dd6gYLui2HNxK6/w26dfkdaq/aiqX77L/aJeMXe+2z/a2DhMmr2lMNWmvf5TT4
`protect END_PROTECTED
