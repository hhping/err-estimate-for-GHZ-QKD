`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qnjCSav6gr2+Ua0XmXZQL5nRm9pGiB/H3y+Rx6CeJ77gmsat9AL/ooKtcIIHSVOE
K4c3Nr7sd/1aIGqPJZ7P9q0wIVF3d/mVvyljIB9pcRMOllaY27wPJrcbvifV/tLl
06r0JhbVhhkgITNDaE5COB71Z4zk+kNj3yUb1fGjuDTXWTDio7YfPfDkr06VyWOW
GxhhpSuCwyLB1x9A9xZIlYh4ImSs0eedsE9i151Qfnr43uzxWH+7vj3+PR5ilAEf
5bFiOOCBPO97dKtUkXKlYo4b/5QnkDh3SVp+LOM0oWd0ugo9C2Wqj/CW40YqW9SR
No3AHdX4D4SPDR950cp9EGhnhPfUk9co+BArAeSBntU2w0xVWd17bQNf3Dpr3O+o
5vCKwjt97w85iqvfz9WQ4nyObjufkiAk5G+75e+Ssb05DmhKhUK38GD//s4Jdav5
Ej9nB9Z4raEpvZlEWm93CaGoJBTFMsciBcHEPao1F5WFtHLIEV/KMJrQD680LGMO
0tX+H0MsGbg/W0eNlZzGBII086wfE4vXUvHOFTx0em07MGY9NSbzLMU+sj3zorc6
lE/QhTNI3X8NrQJeTEQye0z/gkZE4yv5HTVROmLLF7vyc602vGmOwPT14XhZlJ2o
JGGc0DVTb06pHX61G1jCjO8uifqPMjgdn3LDMQqnL5t5i51OulJLmO7xKXwHvJDG
sY/yuWHjyCagOri61JdBZPvdvbG0ZxGHM3ksAOqPxH2LGq5gVN3f1PEccQ2Tmvb0
mxiAQ42vNPZx2Nx9gggSlH85Lci77Bapkm9KCu3JveuQKJmmjXbDokH9kgE/qWz2
7bHUJDUOfVpuBFs/JINyb+lJcOVCxoII3QCzh9lZ8anDdG7PCB1FCh4zzqb9x7Ez
e7FbRIXh6TGT9MwKAsJ3N0KIhfh7lF0hE3yBUc59Ur8Qpd6A5o2cy1xWoAZWJXxh
nFGWrf12K0968WhPaGosMXVKVS/9zcvNHs4L7RNDVc0RcV4bpr5y3FwWseOXYDt6
`protect END_PROTECTED
