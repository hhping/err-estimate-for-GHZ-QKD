`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4UTuIObXnfN9b7Q8N11wJ5AiPSPe8RpvmANtu4WnScLYQ8XE0m8xNlHFg5cL3g3b
t2UrbVWVCq3UJDHTt7GjzgUzb5vp/BvpEYllX/AXT8nl0yByjoFpIMP0hbjGK/ss
AgSiq7d3KCS70kS8mErcphGmD7bTTJFEOvt/asUhnyuAz6xUvpRQ9lIRCABItvir
7fAkQlDnYaitLQA2jS5buKsNX+ceyh3nGvdytX0LpkOvMOQGRxAFIi51ifq2UPqU
fBHFSrs3b4gOddEcEVj4OpFrAYSMHfgMVG6cUQYQzVZUJ5cX8YhDS69QUQvCOP6u
EO2E5ky/+oobCRa8FGphTIk29GYqHbrjrOsVc20zJAwkYvfIxbsgitUyJy+e3KIO
kQ/VOvHGnVDx7RjSxeUgmlakxR73tVFaG1Blrbo4MJmeaWBiuLTORspd+pwwob5G
GvFSwK2UJl+RGjT93JNxE2Lyopwuyi2SnNXEbwkgniXoDhtFLPivDX6tYcZvVbxB
jjxm7LMuZRZOiP2nO3kblBuYp9bBeT2tLOKWDFh/9/Vm7I8RknS+b6MmRcSHAiX0
ykX3fBE5WSkOs/wjwCZv0N+v/LPGGoXUyiKpH6tXUyD1VkHRsuykB3RFrcrC7aql
ZukHCabsEGib/s/x8kPUBLh9CsSqzKoOYJBYE7CAoP76wxb/vOPKvyPCDwYrCd44
hp8a7SD6rhr/T4RSMKQ3ZomZ368V8w1nCXTJT1fydQFtfQgweLVSXUbfxSEbcT94
KmWmbdIFH+g5iyp3vsR2AyGFijpmU7QBS2fTzYbVfEmP6mcexjBEPTTv4Pp95ZwY
YpPi7VmjBjMuO8jn7liNMOomFMUxH1DJ8MxSgfe5oyY/PThoZ5rvHNGZDhj9JFHb
Yg1uixDST4eFC8n9vWAa3U/+xCKH0rwtZ1TUl1xjraYbMKYVa+PZfKCxfUEFfGFa
Rqnvmh6qqeXaT4ja6k2PdS4dcjmsYLr/U/rUClyfr3pWYaoC84m4WKxPzsc6TSGw
3BXCpvajzOxJTAda+Y4/iRiQwvNhADeBiKZilXCeJDtLFZEJNlqURpJkNRd4c8xh
vyQCvmBNAWBdzf6QJcxL+A==
`protect END_PROTECTED
