`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v35j3oWajIF31QUQlasf3E5ZN9BRJDYWoG/XaI6bZtHJtGOKZBPd5iaGJL6YviiK
G1yvNKjAICyyqNBMLVhAtzuNC6LTcOvK8885Xtu2hupT3Di772rv7/E1sfjit32c
Bvs8B2UTFAatjiYr6dEdgiQq6iKb6jBnKMZKpPs9gzO+Q8Gt3GNcv2Teda6z/Msa
ByIdN6jtPxuH+zWKnpU9A1hjMXcCVWVuPzU282WYVgNkhUTlr1ZVziWrFSPLraag
w/iqdXPQoUNwIKfaM2V3s+r84h2YHftONrhavVjWKbXeCiVjV0McxT2n61at5up+
wRgGbaqMncxIWr28PmYOJQa3XCRLtB8Ds32XAzyvf4ndTypyO0982d/sUC1IiHo5
fmwt4o8eKDINQc+zNc7C/RXNg8r9IHi4eo5ZDp0fxoCxkcmptE+AGXs9j6iMu6eQ
gtySCjxRedLPTBMrdL30Hjxj74c0qsKzVFdGudImVtcB3yPGEw8+aJJVqkt3Eg3Y
3jyYy6PmafBtl3a1yUlEmJgOY+h2k2hiPvC3Zk5mAHiQbGMdFES+Q4y+Z6gcLNBl
UC3evuUmwp83qYmusnfLGqNnETpvPJuyKjnykiHCdEuXRFXh59XWsGATD5KLnlsS
xgs6Z3N+I8SRH1oTi0TatRpNBceAo0bi/YLnaJNKJCKYRr/GaymsEGRbJVD9XdAk
EDj8+fdnfmJKoreI6WdA4E7wmvY+OuBJo1Ijrx0pLE/DkpkP0jSFw95bLPa+JjNu
/cViz/ztJa626WKBTL4R3jVQ+yBNcgsLuLQ0R2WGc6AttH1UlMX8YtPhncWAYIKl
I0KPeRuQPPB2bEiYRRpNTWUSDqV1nCwaSj9sD5H+BbuDy/4VDdXEqPDXaiRoLdO2
oj81SJkVQJNeSXMr+0pQ6ehHye1toM9pUxGvx2AzdwsqpwYAHt0uUVabc002RtRU
9wCpCUFAYIOSo0wLllyuFxI+8eofEGUsz7GDF1fZzR3pfEMM862iqKiX9CdqmibJ
knzb9FJOqzVb6eoSt3l9rQ0mPBmsc1FbaZ2Hr2+Xzy5vHLgWx7kI7Z7N05+ztDcI
1y/etXhpm5HK9pIvu6w/lB9Ce7d6uqWz2pykGUIwxTyD41S0wozeffxAkIFdiN2u
VnF9gvsAsy/ZTXmEL3HExT52keqjpRmTqlnnPLVnzqubgnBfqoP9cJQ303GTnn0Z
Izkn/DOnr3slsnhc1npaCDgLxyU/Sx+BROsCHB6PGabN03jbfdsnj9aZbtRJeeBC
6Y2LMyn7nayCGJBTevIJbScD3i1xqCcOyBLkiHnthP9ui9b+brScHz/jGDx+j49w
+HFs9AIXUzJd6dI4i7xJeeV/oCXkqnAO0db3zPV/MGEEGZJtJO+vADMoDSDTVDOQ
A/1O62GHcyahKU4npLklrWn0XMxjrvwMKcoye4YPjVX5Z7gesbvLbim7EIgsxdd0
Rra5iaK6Zk9xNlzJETOsDa83UU/+xS/4SPA717+t4EaEOFjjp1Z+UjLx88fEdKsL
dQXY585WoPA0HKsQQivDO3SpcJ/qkoh2TgHvCABlnrIgXOpHxpnGNKXmqW7ZdnuT
rv715NWbXJUG9WqTam4Q2LN5kOKBfsNJL7gEWWDJ5cL4uieOSr2douLJ5z0qQp2M
cfKExSP+XL0KTwxnPhfcCSfbSbhbl8UJC94vP2EAZ/8mkmDFqG3We6KHTEt+6YVx
jV5JYsYjhLuNd3guVad0IbEhEeVtfVNEea1T3xXyRR9gy9tuL5Nc2MrZ9b6yO0zc
QR+I5ZaM1kJlhSjwoZhAfupPFQyHq+P4GzFRzF6hwAJTyqAiLIoTtNcbrEclxYWR
ZBkJqsNMPqWI7R0jklVt7rskPKuzGqktvRFGcseZSvqBzn7i8tuWzrYDrtRYfNSq
Nh73F28kCgFbTIyXJQ2HWwRpM+I2piYWkP/BsuRpcffQeW6dcttfd8BH9jeQdLwG
OI2MqQPNZeYhq+x7wep5IXgDvwHKplpehrnGkXjfKikY+VsL52EHW2gwXPDL1mlu
mOp2SmGFsaAMFyUmPh4785CmOIXsOkPUDgzaaKlQPUeNUIKU8EuK6EEBPPORgYeb
N2+epZ5JMuQZ5P/42T9nwGyrbD/jugEHrrvqbtO2w6+wHBJ5yK1w0Io+b/wm7gVi
2ZVqIFA1tqt1Us+51hfIul7EZJmOOt4qvJO9I1uHbsnyg68dMTp0ajY7Q600Pg+1
wwoKgB7/8V3RXVzvxkQnJYuNxQcCvqQ9cegd//qMwSnOLlkpk9uwHJPh9ts/ATv/
J1BoILQSycbatSnIYzgXPaLEGPfNrEaOGC1iGUcXhfRqvEB8fJYv2vSH5l6PAyoR
/IfTS5ptB8A4zZNJxu6SHsamAAXwn/aTBLVagx2vholEWF7N0wsrFn7+6Gt0vM5f
JRrabescIpu+LEYbofmXQ2OHhexca1MM982DYmAJaljOjaRdOISqRNtOrDpWskbu
ycglUUU2oGyfJ2Hf+xt+zq4h7HkVOPQ0I4kUsDVXgjbPbUnrqWaNsZWZPYwXzZFh
dOPMh4YMPgqSGn/kc1NNtE1Xm3lRIWYJ1mmDYY8zXST5zNqseQ4Ofr2vplg1G7QC
bkV8LcKmCfAgeYjq9rkk8pOHPAmGtFg/WTrdb/0dtIT12Y8RLz62UQv89VMTSEJq
Qtl85eeciM2Q5HJejYvOqK72hkkEFEOP612ZEfuCffFBtwkU16TMyX1kcuBzvHKi
5TFw/vYWp4q9eceyV8GZLPNooTlG+skuhTIUNYaBtSU=
`protect END_PROTECTED
