`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g0szAE+vodrF5ZnKEb2D3m931bamVQKfRuuy+IEmJPhn6Ncx/dqoOBLTgUs1yIBx
UnZv7I5HeHdxV0siP5HBU94iV/zUA2rTSuTNFAyVPg0/37m+cAF7N5D1qbaa/acR
nS8xcx4AS+dSzJDbSdTe89lSA6quENnpZEbfkNiSlnb9Ig/6VUgrqXlnjkX9h/hL
bsHCTSg5413GhvkcqDXiKtme1CFsqReL9wbsU9YiqCQFSrJ64Iei6fQrWJ0aQnVZ
5qRkomxxup8G1PxnnxUVRWQXaiX7fBjANw8o09QcUjSZ1ERwXfnA7sF1R+EKIITF
UwEe2sThEJOfAErXSZIu+YOVoOaC8rJbMf3DyXACyjGd6Y/YM0HpNQBj0un9uy5C
o5gP31EFus+SwWytLroZgoe0Zz0vy3CJ8lbkDUGhr6qIvcpnqtLrLxSz0xmvLNOj
7uR+nDGSiqL9rhAakAv2quSMLJm09Wm4gfsx1yNpEMnIK3WaLMcer7demdoPMWch
trQy3EKzbrz2HPeZZkhNvdZWRen02COEEqoE05m5bPk0c0TqBQpL1X8nQi0B+onj
K4/XaF0qzT/aOyd6dT6daeauyStELtP3FHrpD3xzItAZO+dcPPpBYewhf1mbTsHX
8ZdImdS75ePcJ3B2kN2iRSKvBedmDLTBa+DXalevzO2CwT8m7Nu/e5Ak+slLtxec
oh4SAMRaEMiQzNSgWF8xgpJCYAEKqo9haLHqfuXgJe2bIWEfqkDFuRaKfc7f2WMk
BaC1z10aaAjar3y65+qjXhwgnsph2n7mR204oUI40GLWfl1SYopG8bKpGhrNilRn
FjevNephTYKXVidHjCbQSsCqqK52ZIeP1Rt1XT+0OxcTTSztqDDVbSVWfDmckhOw
bLlQl6XR+h/UkATxEaPINSy4GJGa8mi5GNMDw9A8qw0mjAscUP10tpRSrLtGIZeC
xNIaptBkZs45CSgNDgaSPg+HwGid9366E9j7/lpK8aT9gYMoItzF1eh9bcAyHG3o
ne94CTcgfEobPstGu16qwHMmZ8fEKSsmb+U7I31xRU1nWtNUEnTXNSiDRQPVVn42
R1Yy9Bq8AYoz/lh1hEiW6RMVVZYkapwvm/nprjRwO/6qtiXmBapFtssrtKIj9t7z
IB+qxkUmWdc//JnLhTQ6lH2TtfD3azLwmM3rBzJ4IE+IVI2yaXkOr2EBPR1H/Xbw
yb+KXe14eKZvKJ0Fjn/8d5gXuUdIefMpe+4zNX1Dvs5FAvNTspUI8UMn3mNAXUeS
p5dGDJQu4CK2Jxfet/dhN9tkWT0suvNKqHAXLYX2JIDEg0JSONqjDsgjOlNTg5qu
Xjw+hS39hYOmSr407rBje5KobX0nm7bllLkq7gjDaUS6xUDKegVsp3qdFHxL8SAy
HcUKX+9v/++1GRulmphr3YS36ycdnbaAOFIL/HDOfoHextDoED5YLFPNn8kjz8Vf
7FViYYlDFRj0SDZdKKGBr8yYXcSHInJOaxdkEkzICGAI3hqKZkzKEib+Y3ckh3/O
x+DLPWqWXRZnP89KU8ncMJrijr1cy5miU8tIvDVlzSDjLwSoFjiJxxDfwKzmslkU
BUlMea9YQaFPdEqf+4aQEsCg2NoAVKi9gjmjSkJqcH3JwPBs1bkkOGXa5o75U7i1
D25bWJtPoKLPZmpbLqLGfmRht0LyXASk5aHcIaZc63x8Oy+2MaNUVtIE27dZ2jot
oE/kHHU/EnPPNs3PwFq/drLZgXi5KgK/ptYTTu22oXh5lcXrOl78FwOKu0GyswVX
`protect END_PROTECTED
