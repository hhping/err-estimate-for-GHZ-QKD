`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cf9wgUGcWA2+Q8/vSTtNPNcJbsGu3e91J82cak4G7g5ZGePIoZRFGf1fhAzYjefQ
AiPD2N7fvtdQG7T01hlUlDLMAI5BhJJL8t09rRuCT58y+PfLE4YaI9BBvI2fOpdY
ZWLccvtz+PCnXuWb5mOqB/2i4HydQ48ipkR2siYYgHsKHdp1b6vee6k1IEvqLbO6
WygmfdU7rYiKUAhnHIq5WTLu8S8qEBbt1HT4N+m0/FZDYCgTKv+z3+/8MPngcOcV
fndslsF2KVqqXypybze55H3AOPlNUth1CmzZGou1QUdPY9x0iv8NuaRKr3JhTwqV
m6vq47CbJeDck8BWZAzK1H8LKAT9XfmWnxfprULmGB7qYRLEN1TLUnoduNwpma2e
SWi8Ti9EBXbqOgVpx/uGPSLn7ZfNCmOX8TRr+D55MkgtyxLMcB0EHuzpEVc2ZpCY
x+YNvjjubNvoGsa/lf1krs3xBK2ztPZd4rsIx/L5XuRk2oQIdJO5VmCcDHEwsMmt
hMMy43CsLK6PEgi2oYqyJthi1WlP3M8lm9MArRzphrEq3FxTko9kTPL3Qql2jlsH
eBgbaI1azf7sMnwk94VrkRI4xzUlToTKVffBY1maaTC9uk5lV9kAnxTqwlJbkcfd
mfLBAZ9sA4VBIEItNLXT/u6UDI3UFGp5v4JFsXTLN2F6mArFccMlpdxLGwyTUtK7
u60gLFnBDYnDtACN+kybIMUbMG5vgpNL+NbDXiHUSetyITyHf2RymxHpZmPLWmFe
N3eNN6T7i2JngmEyAjELrvznFY63kILcSCNODRS/5Z+h2SCeCNk34yT7lOANkA0T
RQLd3lfWAgvdxRWPPLwxbVedYsdQtBXpAV2+bmM3L37/CnuziE1pH94L/ZUpgNjA
qSTvoY5URjmPBRoX7YNZeCK0tE3nWHQFmFfSu+rZlmUU3VkHaT7oUtrhtswYwVoO
+Y4EpaXSEzBePJa4Ac9PEPOdP+BXpN3wAAQmFhh+G0clU6jf07TMLoG+JFavDM6w
R58OOYyZP8dA1hFgEcdhJ1vnfQR7yM7XQfRNQJ9P++AZ4sv3PJTObH6yU4wc6/Fj
vz+CaqKDsbCLfdPVLWvcfj05rRaUsJkmHX9s75arrXkyVo5CT0B00nWKyvahHt6D
WUpKo+2avbFwyGBAjY8zHdSLMIVjTzWHTbYIOdB7Uowq/+c0HKL5JX96FIcRWZyb
YY30WTKed5szc/ISCwipqTnKfFSNJD3rotzZnB6nMYxDmZPc90fLvwbL8h0z/fB1
ASFP3kqqj5yKNLQtSU8BqAIbJF2KIs5h3cBqHdneKabP7K+GqD+bDmPjcXabualg
wIxi8+ebfuIZx+jVLrvVQM8vqtTtVxnbTWsbjeB5g/ypgXjil4gPixbgW9frUH41
tc3Huacr8CJBNHxJkbe/yY9UkRST6f802H8BgHjDk64Pz8WCATSz9vXiVRIIpbF3
BnSMq4+lS/rjTwq/lUImkKoOc+qOAsHuwldTcqXP2MPTVPcaTqUzJk37RcRKlJGD
wq2rmD8rtIpY61ZNjDeWeMZ8F9JYBWAE//3nRH7mgViPhf49e5PZzOdEb4/RKy9A
Hs5p9mboYzrduLp+8ED/4mhy+8bqY96gVycyMUWj9HhkeyluGjXJ9Fb1J4j9VuSa
xgKy2wLDpgvqPaE00YWfLYNaM2Xj3ocmNA08RY8uK4dYmJCm0fDqwd2EhiWjY0HH
xVnjXizDJPjeDqPDJag6wOgZ9md+ZHiZj1Met7KPaggUTcxF80jWjMx+uTbzl6r1
rW5onBURTg7qigIUYOqU+YFk0CmAW/zBYO9ftjrZC+7HZUrzc2gNuKCBId4rsrWl
Ou8WwkmUytW1pCC2qtvo8GfOtL0/2xaD4LARwg9NDx2HUlrkfGqyKdEFV8HmCW77
AVxVeao1y3MJY35110eBMeiDxfp0e5gU/Kh9KDWDS7QW17bz79fvXmZv6QGyedt8
RXDufMsMaAhEUbBfIFMAg9+KPTCQUVd5r11ShPTAPmM2bwlJoRcZ/7bRk5AgBW21
K3lPx9VBbi1M6OvHpBJa93LC8FoAoPnOjiRVs9jgHiwQpn018dV5Thji+sCHsfa3
VIKzWxqRcjfPzoeJbf3y5nRdO7tf9GkxBzHTha+pJg+2Oe2ebLMp3kvbgMhW4PRq
vKl8fjdqipdpEe65fY9mej9g0I0X36crflcT3oNwpR4uCbZPIyh1HVtFRy7aJnMO
YHEgn+C8QdrbxaxEfg9vZdsSiIB3k9HdDTNdAaUTS1Nwa1vhyzZwxe//TqjCMA+0
s8UFtQMddIOPUFM8lq2wZvIOz+NJm2sCiAU86bk8j9P+CxNKiASP3uk2jLYBJ4f8
lojSGoFUVsUumKh3zL3R6vdIozQbcBPKuT5VPo8JoKZYV35v+mZlK3vbIxjcQsYe
4VTq29cjncYVyzFY82xIAcO+X0OB6n/APLGvHfFyTa2fzgzIhNCjhki13OAtfDuz
9L6a3m+X3FOP2rMCYeIXr4staJj0ayQJ6fdMg3FRrY7Jz6E4muJr+Rqq20j/JPhv
e725b7l7ybNwwNHXbm1X9oM1wvFW6IhoVLkwheSfnKoguG8zcwG3633viS3Nc64H
W8JKhE5437qutdWNl6uQiWP63/uTZeJILhJ0zZc35Co/idNs9lf1PT157Nn0osJZ
wtXlLfLLQzuFqTO/goOxD5PEBXMSXLD52QosdPn/4FV+jbmXPE/cJM9io3MBBEVW
BM374Wul2qTxzNw2rQRbAiBeComkDYGFTuZnYOf+hXK0q9saju8Eu7NtwQnnT1Ny
9t7M9cQyusbtPa3c432Iw1u+xNGGJbYvqoTlwBkr5Z0GpxuCK56xDUXWd27M5nQp
y8caFYua/MNOhlOTKs921ede+jUqj9PPqQvNrKHUA0vLH+lcyI+dFDUwzO3ShQq/
5P21BNtGORPKfOEqi2VezejKAjQnHQ6MsM+5spvxpRn3jxqHxOY92/+si5RmS3nA
p71SSRk2SnW9jZTa1hzZkPRQph7ChyPSKwtyT/iRtXmFq/UufwC35ISfBlViFKzC
q6/X94o3VxU6xolehfi2qkaG0oO0yVuGS2R9GuU0JWJhG8+sMl0zC6J5wNRiEqMi
OKMyvMr3Mk7ERhKp/E67lNoURnBgZ0OX0vODHVYBmBbsEDFsuAd4GQpKNwiTu1lz
saosCmXsw3x5bpkESxYg2l9UupZt0K+o6npVQg0d+9ejtZy853SBRvaBTlPLMj3Q
wSI77baDexZLiyx4ihD9tFaBP0NoT8AMIO8CigdE0z+bqPW2Y2hScH9+pCUnKD5k
X1RfQtkrVGo3c+b9cUlCa3toF5oMRV9wLpWInucjyUjUMLqHILqgDryoSqyeG4CJ
D/maP3tC1Owwji30dKDeNw==
`protect END_PROTECTED
