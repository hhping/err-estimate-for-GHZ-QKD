`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hCLgBVsVtDKx7M7GiSWHlEETPcsfBSLyB2jgxhHPRI/+S52TiFAU+AmRgcr41YJL
v8VKyS2kwwr2IiaIpGPkdFEohoRxpCHM0r3h+MyjMaxwdUzIh422yiojCRRWoR49
R6MQuXCNdD+ANXnsOnoCv5JMv6nLHZ6ZT8KKcuI3NePpxLDrNrBtZSyRGfJgg7S7
nVja1m0t7UcKyns06S9ntZ9WO/MpfN77t/Mq3D8L17bKBOpjIBxw+U54N68jio8Q
2yX7PD86JRlT5uHg/2X+sluNPbGVW6LKvo+GnB1l7V13oR5C+wisdoVdWhX779OA
DnDT6ouw24MNFJcAXviFI23gv6FUPGdpxa9gokb5BpzQUUpA0MV2gXTzfmKSvfJW
rSe6Ml444YYJQTDBdYgsUTvXoqMvTIYmwl4z4iP1hJkTL0VsW5fQWN+OHp8QJL9p
MdVoBVcV8r4N1E5zO4qP/2ZM+QM0fOtcGGv9davkhYWSkCwBAly7ajagRYN30E41
H/QkH8Z4q2SzLwYk9UU7fmpPZHDU3Tmz0z7auzgyHqNZohxWMbqaK5M0TWf2VinU
izC756Ux2D21I7Rde5P7zh1qW66+spUw7oF/vIK7rHprmGvKCq1VaKPTQmP96giz
3Bzi1RcDeNFW3Gp8eTtLQDdbtTJNigAh+nqtGNRRVmkN6921EqzxJA8hP01ow4ip
`protect END_PROTECTED
