`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1VQPMffShhWQ6DevJ+pIkNGs5Ha2BYd4kfhduQy7cDJJ1Tl0durbfT2iXXi+zh9a
ftzp6g/3bNa3/BA0/mwJv2DNx9WHNfCidRmoYo11luAbjzyNPuOmH/kaLKJ6qffd
3QDkUX7wz2HisQT/jmZ9EL9tQyDPMe2ffsXbqoCwhoZvGL+CxQgqz2eid3gK17iJ
WRyKnDHKT50cCx+uamemZ9pLCz3OluYLSCRxdZaxI2cLgNqSaPvegFN8YYdOk1wr
2xx9MlojB/CccwSyIOL0pE6FvRxtCR4UBMMEWe4dVakw1/ivhCSFCV8y8XoajCwV
fwqturcIReXO6Eh2wKeYjvspSaQ175l91FxchA1kuSxX3txoMbuFgjU8j+B1DjD0
id0xoJ9PGOJ9hCUOdMH9wdgl8tUFK/JhM1Iij75mFkBBTgokUzBYPEdC9xFMAavb
Ixh3Oo6UNTjMVuZfUlPK8YYlGTcZfhaI7DplDTHiFFv/JZsXZqosT6sizZ3PcYv2
7Qc+ov355a5aKde4Vo+FudhdX4DkMK6h0fxKNLLEQLPmG9wbO0Zy3SFCF8ClARXd
IWs7tiiwkUu3wYBj0nneIOKjoOl9PP/Q7rwWZ/nON3Idx0vZg73nH3VmfAQsQgh4
FygHKtDBGe3XcyI05JZ8S+UvreSbLvrAR2saXIE58CyrDaRPqsSv9CXpgXgb3Yrr
eOjwPt6wWavtcEZFFVUyUozXiozhcQvEUzh5XSh3WnfWgU0cv8IGZhsRYe3DiGnh
Jkh8iPiE7XKEbnEaZcUu6pPpZZClYmhdSWFXnx+ToXkE9jBQKkDDGVcKVuRKhMiQ
ayVmB/s4pnRDAsMtrmse2HMgOjSEeSz4SlyPI2j/8ke31WYOdgPD3Pv0H2D6CH5j
O8nM2fxpugDaziuyqwwyAgIn3gJU+VLJAzZja5aRTQHqGoKy4jC7XOqdezLfOTxL
bM7rqYgDjaQ281jC/wf8Hye90TdMKETTkpU9w65lOFRayC1Mjjafvn1wom8Sn9ID
6PuBEa59I8mY2pMcYw+ZUk8H6wZDy4XU5gapINxhX+AGOU4gkQG/xWHPtIzxE4Fw
3ZVs4PiS8tkSsJFRI1xwNY+/RSk/Eyj1qNJLEhsJtBSHOc1RF+4IqJQ3kLdcz4s3
syKDCiWp8yli4oP7yLspJOXtdwMsw8/zh7t7nTVQo7v1/NsoWoHOUNy2b1kj6Hv2
9QLCb8AQs+KKeoFw7TM32iGfdlIIwFMMW8e6PJZM5Hgmj/2N7OrI1E/M4Gd4ZxrS
x71QeipvVWzkNVHy+fMVMN5sRcREvz7KmOsJx/axmysV1D2sC0tfxo1yaahUDJG3
Aj4X0mWSBwKng5iMrFgQ5sZiD4hrBN6ZXy6hEsnZye87WCCabAkS0xs1pdGf81pJ
ZSOOG77Zy18bMSpDXq+1NQ/aEo9/+yfXj71pqqNruS6nGny5mW1Oc4h01ti4EZM3
cZAdGwm/StigiOJXYZJAIcCNKJKH2hbODJEaUEiQdUXCQ2hd+SBgldhSBJsEIrX1
y9rPPX75dO0vrmhtr7ihceZs2Juawj7xhP/DCoPPJ1h21anyqbtw/hbPhszXk2rQ
eNvGOzohyOQ2xShrtnS2Fol/V5K32/ZU0qrk6HD1zMbY5KXwLbxEPj96CT/uUK1N
nu8xWRpIN6uajT7NIyZJg9RJc+Tl+d9aq5reD+Id8OEGLn9XM6p9tgPeDWxW+/n0
rNVuYraU4EcLGslp5RrXhbnNJwoWrm4UEN4CjoIRXFDZZjC7TdPVTkWSpFjp4CU1
xjgskg/xItQZ1FuW9V4PO2+WWOF0bjOJR0PjbE13DxIH9AOKccFNUEsxvLM5S7sc
i1RLV97DAd9FdCMHEXzuVtfWmQjWctA2iTbpYaP/ns54qirAXGccNzzJhhYOYNS8
wNsrVdQxMfXdGOQCQ7TsXvTpo9/9Xr5s4+LpcQQ1Sj+TLJW9A1uXc2n0NhCOgNQC
2x6kU3dXwIb6DF473TCCt2W8sTNyLgrENSftTA6GgSme6s4M1hIml3t/aS5SMTGF
EXExUL7l9/L1+mems84ace51U+QSELnswb6k5XIqVBXCbLkIrsTk/cTlzk0Ykn5U
Iskwyj2UaeMfOA0+oNDpHf2iNjn5GoszIZP/Ry+/bkXX8ui07Qcl7vmPb/aQZW5p
Mtm2m+oB+9/fVrv71gunPapBnGnZP7Y1E2JW9zWzHYE5b0bEvMpVAeyFyQrZ5aYj
tDqHCJ+1qpUNhmMFbZ4qgHRvCz5gX9FxOk0RmRTqllQmJMTTk2ms7kyfoAzYvwfA
BrVn0X1ktvT1n6/4ul6oUtzbY+WrcwWaSbazTZRT/4GL1MlmQF8U9LR1bg7n/8ou
STgOdEBqThPbwCg1oLIyAEsEKGqkyjS3zHBZP4mtKPLJy2UcbIEBujiIfSAN0PgP
poQBz2gG9/MYueAvZvCAIpYc8Nqv66TWihIdhl5GfZMpvk91LU+eshM4Xcv8CXDm
LPb1McYn+clYm4NqjhS1fZkDDexuPGj80VqbpuTTVayguJMmpoCn78T4IFFSj5U/
b5F1Fs/CBoMbACRZiobe6qhBTfNRdf3CtZXfPQhU1/BUWCwqNVobQah1V9XRyMPK
+DHl2s4bH9/pqTlqwdpGy5i6hc59Jlh7kaSCbzl0eVPMeTJrWW/N74tyWZf8pB30
5/aGDoIm24Wpn+f0H2xssaeddPOAqom82H+98qLjPNFdKjJq9obUDoZT+JKw+c8z
nnKLyi0of6wsMTRmwuDmxAt3hxdorPsK/1mJd2fwZSodZ59O8Aveh/vshZ1nAYvK
g2mi287qsOfxMPIBqRTK+F4jUXgIZaETk4Atp8qRncunsPdgZ7NypBZHitQb7Hyl
ZpMCFFaRsldkQq3PP8inLmQmKFLTItG94pAiNiyD5x1/apMzoBt2A75syV/ghFvJ
0eh2eHYkpecqQak4Gj0WvSj6JibLTjzZLaYKgDRvEPY=
`protect END_PROTECTED
