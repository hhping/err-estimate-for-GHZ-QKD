`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LCDXcpRQqy8fg5fS5UnYPXdYR5saw4U1MN3XubqpdigTxyl/u0ebdCUTW7V80Rp4
KsUa/OnsopMUNkVhgZJyqeoLiinuqGTooLO6ublgb56zF8qPlIvTqUFSNpFBJ9YT
M0Y0uHd73HjPPJj9d0hLEIKqh8WRLDyPeMysBCMFrccSBwgAvoCjSlgS+gTvl3KC
71gmDiqNCc+++EMZt19D63dqmNE+3OrooJsTSZSPlf/Lc0DEQ7WjKbKJGiU1ebm2
mt+NOLzSVVZB1Rn+Mm78EfMSdQx6xiQcHHjyq2s/GmHkgdDuPpFgmAXLZCyss3q5
lilWguAqQ97Yut1qGc/1lz+2Rve1aSeuqrx2Zf4KLgvHb2CYkEETQ+nkphyi59j6
jjcBPfc9g4cNHTztNdFXAaLP1jq1HCR/iuj3veon6s1O6npX7lkMjUMHSuizAOT2
x2H644VwcyFAgNv2qa2I7RtxUbYpgzq3NKnssQNDTrd2HCXoJzSBbifV6QEB5CAq
DgDyXW8JUMIPboA3YVae+cyscjhZIJza5KNHOI8IjFdFrjIYStnl0cwd+P6Z+ljD
JLHp0Zimv/vJMRzMVO0KO6aTxIzyLN9Zi1jKBfFSnPcxwqZGTpCsw8X0g81Hee3I
xuklkA6v4fdC8mqcm/Kwu7ey5Tp5p456bee/9aleGo5oSb/eV94R1WLnAhRwH6tP
RyZsMDFYpm99Vc7ZGiiEwldzFQj0jb5H3vUPgMis+NCZ0MBFpnN/hoY8SwMJfQ+r
z1u/nngru2NGbfMff48px101qg4Kjr1SQVNVHEdloR4mwACF44vk2A8cO26nnTEQ
N0wVP4t6L2Wqw/WB6+CCj885plHRFQX9naq6eOha4pRvV8u7GNGyMUjBhNhtV5nw
Bc0pNzZ8JibKSeGIXGkjPHfdBEWBN3PpbUPekJQBsojbjLEmst8Kd1HWfkPDLYU3
7TwghgpfU3FGWnaEvfietJJpbnzTcZDR06L+WnYHZxUKQE4L7XEOc5gBFJ5pVf9n
GizKfxcGh6y1CxE183P+wco+OlqgbZx/V/y+LrUlN1Vy5fdxJCaDIcmK/298pMtH
7ZsvDkQi/nbgRtDxCO7FjwElOAwv+sGAPCYBlvh9jSmSHWpbxi6+fGunBDjHAxQ9
+quv5LshrYZqM10Jx0YaJMqxN0WeH45bh7E6hl1fqW87E7GqnlaaMZ9v7GSj6buj
eIaK+JFu1QHX85nLVAsAsFCFFUW2I4TUtQEd14uvU2e6/JpiR8jcQeGSA2yykOmA
oc+Td61O0wti+7ka4mpkdYcImiCfMfFZeWoaJgQm+GV5ifIjErTlDYRWnyauSmrL
XyPOOTQFaxfU7KgJcDPAabRukUuLr/lGDsBvrdJlVxjtjpCwQdWu28dWRW0iBd7r
CBUgD6/aI/ERbU1gTXZlMdN9scJ1zdZ8Qj4odypkKZRHBQvjPWRSmlIY+U7OVNAd
lVrrgYyqoOFewi3KCaWwCoIMFIbr+MgWOhwraWkZcrpyUvJgpRBSBeLa5iIDJaKi
5mggcrql5e6C7sEtL67Rr7M0cd/hycB1nhdjiHpcP1fBDrGhCc6kkZGuYChWuvKy
O53vMoHy6755m8uw647krjhio5uMMoJ2OXibVQboyv0tszchOQlQlw2ps75FOkeT
SOLlsUoN99nGLWTj2nMZYITlkgE6Lj3Q6QsJF/oWuLLKAvqy56ljJj5bxpH83/6o
cYA5BHHqII7nfzR5VFfU1IeFbyU5Z3c+Gvu2r7Wr68gI59rDfgpEeAawV4taZTrx
3MPAQwX0LPlUmEeYiM5hlbw6S+W2UBNOqE8LHkn5lmny9J+0qrlDjuXlA8CJwflh
DKgPmAzbKazri4wuP4H/pG8PtEP8MNz9pXlfAL7i05sYiHDQ/8VdS8TlKXhhbIt0
bn1MxkbHDZWSyxhzr9pbCEqH+fvjYtchHwdbqxp0hol/JIlMk2WZTLYHno4b13aJ
Nho/2so+bdMfT76d9c3teKIsdEjD2reW0e/755nf4fzt/VGwQIKAGhCzUkwGBuHZ
5e4HIuOKwSK/PVey4tXy9N6DBbxB96ntb6DtStumqrvT4rfgmxmUhfoOpWjXVBUG
YRmOXcAfKbsuKBc0eY10HE4TKhUG0PA5HXzq2JN7cFy6OOOh2Q2ya1dD/47AgQ69
P/DI393Nh50M6OCN7+M+u++0poIcNrV6Yrm4GRSzne/pitOrlB9VNjPGgjOWOWwP
4vNp9YaAEWgf7aRGGTkoZMfPSYmlzOhcU5WDSDR4XuGQRV45FQ4ZDkWNC03dQ5Fw
PVz5BkvfcZQxg8MdEzpBdWn3q4a6+klzK5ckVP5UPvS+2fKEUU5kExMCyw6GNERk
/X8TwWWn3t+pNH2S+2Iq57VAdW7OZZHsBK13nj3adGNx93sI9OPg8yDcec+DksGz
HzIgqFYWrUb2q548DJxjC7SpATjn4TcWLTri4Pj7VN/OPKobnxGSm+42SRfK0Emw
+0uJTE+bG3AYNeHGWnaqkAyRdMMPQybq7iIwv6THb0LgLuU9RPcOXYWsS7fhIAWJ
1zazCqA0dl2XT4Ps/SDDespXeInz9oeVW8o72pVsoS5I7/M4OthI3SlY1fSk+DvW
VoJdSc7E8BwE7Nq6Yn7gRbhwwnl1W8MutQmSJdYhIszqwzOEko4y5GLUh0EvuTQe
AmDfRdr0eQYckoFryFr6qGQYEfXAZwhkWh1Js/p0M7g0sCiSPMPkhxDDdBO/SYxZ
IJ0+hTRe/W4XvLhnnKsSHg5ghlbcXQRRu2SHsUgAECVf6S4GaMIBwV1Ge1uRp73/
5NKpChO05irOZcdrbL42ZOm71e1lVSDufCVcBA2smALCRr4/sKMRHPJShRlknJVp
WBMHTRfJtgP78iTtn78/+rngfgq6isNzmM6ACf4vImkwtZ/8hvt1BGjiCZQHZ/Ml
LVBM8n4Rz0zbE3j2t5Ey2yeqyU2Z5sSXPuFL6NmyeNF2gcsjOUTloMQ4MZKCz4pk
uf4/UGSNQM4h2HWInYCiq94QSO/T4dnQqI/sTjCIp3M=
`protect END_PROTECTED
