`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gy4G/Dj/0c3CFgOK/212RTTVP9FhVLnc1ENmr7QILRdtUZ0YbRPUNgq7uymUoWpj
gy+aGO1a3Hj4qy4fO1euzjPIBWX+ghN6L896GKoOdD03Zzf0VNdZz1j4F5Qg653/
uRSMDA6OphFg/0hgJWUP196OP0G+eYLTa8TLiCjL2dPRaRno95RkPz3XVgRRMoCR
hhrw/jfk/VjlxepRajc/evBDyfTSFNomaM+GkHDDMvYyTXky1cFzzZyZmRe6QuRC
bqv2Z+yyKYrs4t+poZe+IGYMuENv7+JBA4er+vzK3ksBdljIuAApMpJ0QrmRPkTI
iRZBmZDergGpePn0ynaxaxW7Qizjk94BYWNa+cfFj9NPquDnMKj7KG2mVM3+uPup
tt0ZM/08YHhMiS78GqCoOq14umPp08VI5y4zFfGDkAQazGFLuoZScMSzcp2w7E+3
K95H4uxV0WMWJ/+/dNm18qoMoiMjNlo1apUr/jEd9WJt3tiHGW01R2l7SvG5iBGn
DhdvD5OOpCSXkVbXeUcOwoEscl2En0gZzrh9iRy9fK5FKChAquMVDqvscn+sEWxB
PftVVUSZ4uv1ApXNOLTGIFcocaLsfTnQtV0teQF7aOtgvZdpK9I+Z5yitrlfqpRU
JEWO9IiV5uofHZ4wNrAkxo3vLS8E3rTIZwqheTcZiXIBUYALY97hrXfiEsMU0ndG
SWz7RD6Jp0hPoINYYHjFaUtNYCW0iN6gSVaCVzjFGZCZnMBJvrhS0cb+1jSW3tvr
NheB3ZMGe2h+wmuPj5Zz7a6O04Jajsl+Idfqwg97M5jCKG/4EzyAOWUPxaMmM6j2
4i/gEdm+K/XmHLKBO9xO0tNIXWs44x4A5Jt8TeChf+NHzOEmMANil0t2t+s448fr
cCfBvMHeXMOsZX9uyRBdgT5TBxsJxuWFstUGGnwxegunimUGlS81/MTTVsYUxCov
ttIYpuen1jhC7m7DbDA1iwNeDvP7+6MnbP8EnDV1tyuRMvB4x6ymYHbEgW+vk4C8
uPK1AsqEzdgs/7dtDp4Zr/j3x1bMkfMjqV/UVffTwPSegU9I+rr0NBDDk6Neyaen
K7bG5EXJ0dP2qpX7Yy4zQO9czByAI5TkQJB6WcD6IZWLYw6IlZ1gCPhoGt4cF7wU
vrTBhSQ3IvEQC6qdT9z62xbs4ey8BnKfu+aYrGzpGfP9gIV/umQ41SsCdn69PdUU
BPm6mBrnMQF8pOaNGnf0MfMHUGOl/9BnY6uMdbGUWVbwT0DtEWOxwB9Q1HqTHXvF
8fCqqNz3QN51T/pC02mH0KEK4fRPwdSlYIjmEcUr6uVstOm78ZBwcBYNgyOrqBa4
Dj+VFJu3qsoOAxRaQ0N2m4PGLNJJABNcnY+u0uxVj8NzQMPHV+G7HgFLpSS13Acj
rO7Gorr3M8m49K0ZsPbgA0EN2cZY7lRp6syc5PnjpAA+NU9ZPfQ1HDJsboa+u2X5
8mSDSCmXXr/l0brDD3qkws1ZR9g6MkR7MmikY3g00uzFz3/SkKB3GxXH2RHXgHH5
0MXGBS1eG7N2SXz6iaLCMLQwbCXYyLZe0atim1orMMWNL9ni7gf55ZcGj3uQLvKU
gLz64ioYVcd0C8NasAzR+UcxZwxb+JpyShYHwVPaXVcB9nOTrt7Zc8KmVjLTs1LD
ly2DRMpg9/YRy0+hZ39uNi/wFehCRdgvJsfAeBoSK/eApCnizSbMVZGotj8FcTjP
WbsnlhxuuWmIrzWTEYeOOpsDk/s9cmR8ZBpzYT4LKYiD6bKjmM8uIVox5jCvR5hP
GVDApyKpVFxVoFJF1xNVRoBp/YoXhD9zYhScUQgN3jNCNxabcO39TTsBOyUVUwst
odNHx4q8uioFAYd+bvzrrEtDxrL2p65pYF+69lD8Yz7zSV3BMhXBAS8BbWldVYnd
LZvqbGZtAoW02RU6Ke3/6FjqsizFXAkm/TRR/FAkoiuQZIXPTzHyabF0cA9PRHa/
ezNAhhiHKdKIaUfM+W5lvvJvmWei7iCranNL/sp5w9kopuaDg3xlJtTpqhmT3niR
9afspnyK+PyiSisRvupV7PZz1EGvcOoYqgbtjCYtsF8rdphCV61K1pb9hRXlyoIJ
Gnja4XUtQss/fUti7342tQDhRIukP+gKCJU+bvNQ1HiMv6U4hjhsBwBplIdI6FuP
+QcGchiXdY5hrYlMmjYidPpYlrQpNETYXfbBjlomcI3iaYmQy1EcONXfnmOPuMoU
/zCiFWiyRrYCGcQIZvAv86p4i83IufU1JCpybQz6N5ojAg+lo6MuKxMr7xeRphH/
k+Em1JEDC57n1rVnYTz2PjHzlZ6xCmYNZUMrBbAgnTCK8zPqv/ESHumcyyI17wx8
VOnyADFxDoCrgiUEEIvLky9xoGaigWXy+NoWyeclvZxoO9PedekoTBZrgpL2R3/5
WfpRRjjNAqiF5oPS1+XtJhEFszr51GNSkr9A+2GPh+fOacpi+OIA7XUzGxzITFyB
olBCUb/4cW+pn5YgKflPEWxQ3INyKZOcLaEvzLLzh/+cD8gVc3ZOdFDOf8SmaTB5
XlckYzapRbN7CtgB7V9cqDiIH3zKeYOCOCkeuz9Cq/LNLNBBGrVc4QuNUattSQbj
YMVAu07+H65BMXS7rXB7i51jdTvk7GlBcPuMyk81gRE8VXPJBz8vqHaP7cfprCYk
nVY+/nc2HnwdWXKMJShQn29ItZyC9cePWdRjtHhhS9101FddktECAttMcnAKgC3f
DBTzzB5NQlLDJUaCL1NZXgVMXAsN9M/6k4P8ihp4St9Wpv11vLvpHaJFk6yOkXp+
rNccvesJnUDf6WYtRrYHnLYPJaip6cX/IwOTjE7+fvspr3XEqS54XVTQezt8I9wD
y5jk+7Z0wfoec0ra6+RKoo1h7lmrwAILjn9Ni0FnpRjHYSmoQXtCJEZYKeVcXGAb
gnIxXlEftI6v+4pVQYZyXtVBeWYWK/dmsed15S2ogvaAD1ELQAF6udzWEp7kHEtx
YncsvUts9RtmGEP8gwqNsHWFLRNqiZHller50QMEu7pSoykawcEf5TlrbzniU3cu
z50TZRdrZZKWSfJTMQ4O5CLvW2cbiYiemHi1uV3qqZS0rOhK9b4gfIEnlV+iHPBl
ZSJncQiyXXovRQt+j4VwWycaqN2KSMuSJo/YqvoXM6T399ILtXlKWZp+Ko7Ua3m1
7SqUVLEw+2BZYLHw/IEmZHFIe9oHau7mB1oB43mj3PH3Z+B1qsjC1vJmoEbo3vOB
spRdw1TRG/sUrQ2aBrJaEGgByQxCxJXOzH8fmZzmnQnDZeJK0+inqp60VYF4H1A8
sVKIRcdTOVvAOHlC18rGxcjraXiCvEM4rL1y8FVRlmaJoBMw8WfVSCnIbAB7yeWe
grgrBN97pownu2PX4yXUeMD8YSiM9pZzgeI5kuCiMO5pDwVoX1CKTzuqmNuIbeq6
+ggFyzVgsq22xt69XqqphTQpqvUVWKbGwhP+MoVsQcKHJMFi1CUGZtrQqytT32th
njfB4hcNj7OH5HwvzQT6zXCRkouGTSHTzauUp9G4wk0XXR22IZ5RBiKadAF4iF3+
xWMwMsqxi4l0qeUc21lt3kqH/k4uDPP8GmdZnOG+P6aoncwaZovAbiJVBePYSl9c
QMmuZyL5BYgh+Z1WJgGXK+MRCtBfX/1s5vLq/RuAWmr+NE6AUR39H1RfKSdl5qjQ
Znf2TdQg9CGUTBA15cv3Yqv+q/Bmyv6/87NkWAJdCyCIznGqlPpdFGxTT9VZav6Q
Pbq4rGeNN5SLHJCpuDfa06L0tAiobFDqquNyD/03CRiKLuIeEuRVP+2NddSzW3gV
reMIzwg3VSWXeFiRxU8Zz6uOaHdW+mwcZqxbi89uHP9Y4f7mGgTmQpf6d/HGR+dD
3tdMim7mwbGwo56jEJABducVjepMncwRYsAS7dWIx/Y14GhTCWTuXLUu0X69Gina
SKBbmvySuLaFapYu/6lJWu8690aNVzI6BaURILhZyH6K07PhZhnaDEArXjZhgN0o
USSm9k4ZJbXEH0PPWgzErXIaaY7D4ZRCpwJL0X0XdISQWWitFvmzWOEXLj4Xk51/
LhjqlRZFw+7sbvxSY9hfwejr8OtiXswwU1QO6FH2t07Df6yhubpSH9yhp5P9mcys
3Llt0f6XbfFMhIvY1uQin2bNp8FatyY+rHlWGHnL6nZ5si4P71gPFmDhV0IxmjKF
wkpcg7YXwts4WNC/mE/rX2lPcZ26Y4fWlBNpw/B58Uc9x5DbvP6/xBuegmhR4cbU
f9e9YYvtqhMyBZyXTBIhjW06K4jLujCaiy5TLiXgh6FI9pBcGl9hUzfZqDriI3UQ
zIve139814tnuRFuGVDNYTz7tnaJhZApM4dEj6T03B+S5AEv9Q0kSajdxc2C6lYB
6JEYmEX1mOxaGy2JbyiO5OQHPQuKeRjsqC3gShIZSGTLRxOkJ8YsTGjFnjngzaAy
NFnUJJ+oJW7Zi8BtQicGRPi9ebop8/FTQ/xFxKN+ZfxGQjBACgrbYOcyN8flUrMB
+S9SJqyTuLsojkaEboYDzO6GR6kJ2MHS4EaVZE1WWRSa8C5vfEevNoHdrI0epF9L
Kt/7JVKFpkO5XHdwOGsamTSCE5d1lgrc/eyTYrrayB0VNLtUEEE9f9PMkRrWXw6r
d8ZqpC3NcOZRuNs/Rk9PuQvTwttu341w4dLkAqgKVLa5zO7SDXj46qi1Xv3FfUTT
epFqOxj65niSsxh+CO5y6tjYu9EOGTh4KpvDIGGPgtZB5TZjBKnJIVNWeE7EbMy2
odkX4ToalBooH9HqyCKGwU/Xuk4wPxVchSjRqXVQekL8pOhGmFH8TypksnyVtXOy
s7xMQ3oQfEYazCSIzrE8LOanRgy171Fe0Vl3/uPdlnN3cXiBjqMGLF9gg5FXjsOX
1wM71UYdgFEODFeadXVQQAZcPLY7+yZTVTrXtSdD8n3KjS1DoB5N1KK7klj5zzyS
xdim4QEvQ/iRTkd/PwxKVwFuPnrAoRdQ22UFJAyErTqoET8BP1e4il3B59TTWP4A
Hodv2B1nKdFBQJbnpnil2WmYi86gaOxqT6/yTRYvepGRoeEnqTVn+yzpQV03cU4N
Ak0GLrDnAa3SctMNw8Qj9Z0LCtEomGUCFVJqQZETcS8SYA5a5p0OeB83tcd9lQGZ
3gG803kFIcAQk3oHYZ+g3ETEylEoTmamcYQcEzTEGqep263dFLuPHpyT5uZLHaHN
tcD/llxZUWNpIS588gjkqWuEz31/vONx6Ueexp7m74GamP6Gl5X2sJF/whl9Ovy4
DqcAJpbStEdsxgS6BvBVSInzL70X1vNc3ksOLBPmjmMIIa2oIdS/kvey6CbELk7B
akh8UMi30gh90BAPKd35BE5VLquDthlX7GtYMdrlDSvgPSWfFODALUfmbWqoo7+M
D0t4eoSodPMiGThPBAyVG10MWCAgDh0H8p6yhgXpQrRuJm/aTjxVMKKKlgG8MlxK
LGFkV62e0z3si6C2Ye7OYD0xJ/O+92ptik7MjmGkO9tpEYLfToLLSQRCc1f0e9U+
K3QhNkpa4cT75MUHWXe/zUVkwvpzb5kNW2kv4lC+NxeFOK3MAIAzYXre0H+fxj5h
p7Ms2Eywae5hiZgpuhHsx2DseaISPos0jIWpwhpqqCL63pOEIN4z6vsFoLMRtRrZ
omK4a6kwc3x47vtjenTioi+DA0L6CHZnH3LCxInXUM3+ATcV5b0THj7ason3Piva
YMWWsXOeto/RM+99S7UWyUn3ef8gsAeyPEEeETQfaDCkh58ye//9hL1nU62Z6gKH
g4FEyWW/NB0S7fXT5db/wl8J41r62veSWPXV5H6+vNm7z+/ikoStDXLRjOiZmZaP
ngAGSHF9GvyhDb2sQ7MYL/NdKKh+1/GuwXlluAYfomVkKn36AFbc9XrmZaD8piDX
Z4p3IhMgvmLXl6h5PmU+66dpvYzyP/BIo/XmkZPfpPjXCUREmqz/wQzJgEbhMYGt
qN0F2JFJXEtA9v3mMbbAyixeqJt4TxvqY29xZK5jKb+tecoljsZk1ajbS7bwccnV
GzwhedmBIXeDpSDHD35Lc310InHFFGHrpBkF4NVWOvCMObT0pYZO3rhxBEfArOfI
snv9ybcbzLiqAMh+z0RUL/4cCsri3q9jI96jLIgiTkclor2TULCp6aPTsdcehB7n
htYTXb6ml8Q2jsTJPP0bvXJ0LLYUvIpPNjuPWeRIOlOZXuGtN3kAlq+uTbhdTnll
W9NESsSNx0u0MWBM9zFijnAB7JMX7zAjZiklgy6V7Y65MO90Z6d8YFGaX4EGvaqA
DOxt0fapPMjS+QjRBGHN5/nFCASYmckYZq99duMiCE1VFDT0E4G2yxk4e/EPKu+L
e3TLwnJaSS5/gAu2v8GLE2Ng0etXvjx75wph+QMLGvOlhqYAFQkPDZQ8fpQBKoeE
6YYQeJG+301VpNsR6i+Aa3TCSOZ4/0Fxnx+d6CFl0NCCUBHuxbHB+AnNwGQgfO6k
OOzOSGUwLLl7OKZFr7eUIAXKdbf7rmpH9p0WMO29XXsyM2GNk1fbcDNoAFb4gS3V
aAaoysBTjBVXTf37AqQ+a09H4+X3ExVNzLxL8omImpkjKqjTxrpTTrg4csY6fB2i
T1ayurodZLAf68LyWz1NDpPwszuqm/HOObf25HE1BrTWNOtzFUlUI6S3SCnDoQ6A
d/+yk86Iqg7IYm34zBS9C6PEKUbpBr9e5lyzVJOmat8Pl72o5QOIIZ13GP677dhw
kRN6e1yUyZiDvrTjrM/t3WJcZnPR+/gBSxeUbZWdhS0dMRXgnAPyyXO0NyiWq5DX
XPXw2r2kF63Zievs6hbAqjl7nV2nEdpzjeiKD6F58+an9lEWXDmgYhG2NnEpukcA
SkBjqWUbeZ+rypKqsRqh57PH6izgAv03rzvrFDUFimxzUTjxsSFwSsleMzolTkn9
mhxY/0mh1c6YWcVj52H00kHIh25Bq9n0gV9d87FeGXtPkKj3MPylKEHbXdXHhn1c
Uhz71fv1I85nslQYgBFhYUrFt6YepuunAQVuyJnJ6kLa8W0AyqMwbxtWM1BUmsFd
`protect END_PROTECTED
