`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BwoPHUSJy6TksZ5A+2VL9siEb+lhI50T7kYoTC9rsyYG2t3s5P45928w8jsZ5k26
wvpy2WS4Z8cSJnlTk4X5Cx91N3XSZYMAJ0+p2tVoOiVcQGHJejP+hz38zfmNrfGf
9ZUzMDwcSz7sHQyAnvhmkTtPxcfsIc7UmUfAZZO9Ys02oN2bFiAYyY2tFfOhOAhI
Zf54IBCkbRRWGCCe/U2u36i1lgnXEuSAUzxTSpkakZPphP91IFYSPA1Pjpksg6m+
fmP84ZSJDcKUvp1AnwH/W9laeUXWsEiGZO2yuQSpP4EBnWM00LP+uZlCiw2MtGfI
oPmtjgC/OxykmoW3BETIX4WmuAz/8k41LvfkUcoEsCceaTV7RDbSNxteOvSGsBz3
zbG963BPipKiLOnAe5fj6tG46zST30ErIhUc11icN1mn04qXfObAO5cQezX9qmTA
JceQJ+YRqRPs+K3Ma4KJkEKMcjb8177AHr2/06JY8aQmiCPPrEruDWC/P5SK/10h
AqGJ9+LnpaDfSIQWdjASJ24Y6THgc6rXPvUwsMDCr1QRP4bubbs3Lps6mOAQv4mO
vRRT2+2pbY7IMDQNiSY8tYq2533QzgNT3oC7ii15nkOyLRK/Jr3/m6pYyLLij8eZ
kDznmqmSmq20EnKtnxJFxQ==
`protect END_PROTECTED
