`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4FN/A6em3iHDfwnJjzUGoi8bN2AdpP0BdjsC6UhJgJjP5UdmTOFlkDT539dXwMr4
m0BVSDZ18/tg2TlkEf+N1F4v5nOvsNzDzeApRqiHcMSouKgprr1VbCgTd2TU9sbm
WqH/qlSUfFEP5UeiT75+5rPc6rH5hTEyz4byKBP9kPONvR4DBXq8CJFSA1Vs5BtV
uL9Mi+jV1PFaQJ5W9ouPlpUTfVsP9WyiPMwcfgxZVtxnR2sQuiZBv9hdbetOgy4Z
fUHRbo+v8HzKYliv0uxztz5OMJ+P+/BAOH0LX6GwkvIBVXV6ZnSlGG/ozbM4f54t
IBEwtWdLQcqph37WUD2e9H25Qzxn9KmOuSyjIfp/DG5e0S+wuNkOh9jTcSfog8Xr
J2nItI4+V6KWtRDwdMt9ioU/CLFIIAohQ8yfzhqQj0yycUPBpkxjBZ6HkWQe9cQ6
1vWKgJ7dAraW9yyxsRDPpfiVIItJebT2KFydkC2v/QcFjvsVfSkSDCUfD6OY0tQL
YXKbW5RI++mVHewnmk5gzwVSjzfcB9sMWLOxRZKG8iAosjamzLwu0nwCVTp6fh6c
wcz8XY8odlr3Ml4E6vHDYx0UB3w6E7lxmdSOr9nm3ojMlksWdEDWMguJmx/HX1Ml
edusOdkkcoVpNDgY1dlhtkHeBd+tLYlhozzQ4ZFbvhyHNr4aTJnN+NfGi7Akk46/
2s1iAkfcv8utO0yimcv61fY0ZaNtnsb2dKowQL58lf/ed1JlPVIg6NiwqC+xv86D
H5LumU8tLXot2axi1WvRVEnBdeHp683YlwqVNdmfdfampBLTrjD7HQsHzB3q65Xv
GwbVOQMjt2cmhpDKdmJxk7DzJ2XKLd0L/7m1AYR3iEGaDpH7qnR/oyvxaJhdlQFu
jRtXelmwUkFiumVHcKSX6DTHiPVrnmLB2kwnlR39ATkKHALXO14LxoN/e78CS/EC
sbLm/kI1OYuWKbCFYml+5YqmEcMMRDSaRp6RHXp+Fv3cSGhwtTqwtONRCiGZcK65
+LwAYRY5JzrdkOI6PDk9aNHI7siRwTRvVQ/gimblJvunFJFXTTfXQ5NCqIbdkHe4
sWW4fqpNBC45jXNfeC2gztDvtvK6Ec71nz67Li4rJk/Ey1uYkbkOwfpUPSGULisl
TzPZ0jSDt86hioAN5OxOPsi7HSP85Fh7o9FcxKcBgqCUpERVXjVnRXORAqEfM3LR
3FxD2yaLJ1TrUXCiu1HXglkmu9Nz/1jKc210TjJOpu7y0J3+XWONExtWU+a4Jd+w
+e3TrVwqwhdyL65EeutPgjKCWWBPIf84KtpqliGQmvL/AGRUoyGP6itK1jhWCjPI
PpAVGjc56+OvstxSypA1Mxr5cvF+4MAZNtlM0fxD8pyNGRC5V1l1YLA7tDVqIL9r
ZA76df7xf/0wRCDWlswUM3KSdABl6qz1ZbHNLIghHKdaOXruKEJizAd0FpjumJgf
QbN9r78RM6Qfq4X6TacJ5WeFPjWsdVyMmlQ4QxbNa94=
`protect END_PROTECTED
