`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xcf2PHzwnokgQ8PzHgIgQjJfWGtbioF4Odrx5ki5ssNb94YAX8WNZH+EwB9N6YPP
qjvWmmkzU6K6A6BRI8/xOb+ndcmKuj0ENeZHBP9mfRJAYRR5ggkFkVRUl8LLxDVi
UztRXlqRiJPs15DXosFabTnR9ITQBvie2Hr8jjhCJreejY5xpFkEBt19YPSXdAN0
cKF1qmFrKcPjEtgRsVZUY7/hJ5fW4axZz0blp6W5Fcsjmdd591mB/9s2nyrJ9EB+
nR3GuJfiZ7D0Vjoi3eZ8tKPAcJHvel/re1HRNxfJR+G69mJYX3gNt5ElMVkUmNlB
B4xBFvw3+3jI/sAF+mYk8jWmq4OHCiZtkxHKo8Ti4An3TXfQja6hYRHanJFNgG0d
7T398FEhnLmnMFj35xLTDd1E+tmoLpMy+RdNIEJMv0NAkUq2ElRydLA5slpmCFI9
Zy/G0KeGkY/pwF+7rrRqvAgdG/PGNlJEEZPyjKP9LodbQk3fDJJlnGFig2TCHTiw
aXWJ+s8uEqT47+EfJp7s+eRanr/WkLMFU9GgQAyUwiTPUsIPysnE1cfL2+zLWJJp
h2hreVwRNFkSPs7Id74tcSFyj7k0mHv/YZ6/meFySpQfaT8yBt6cTsolP5dTYICx
2R5vzh8ERtbyrtGB4Dza5GKfZOTAX17gTWUdWzAsd8pnUksTKLlEefBex5cyX2b7
Lz3sQHjkvzalaKKCaeNYipZzXzXNfbpA1NnRdw4pK2onN2E754BHxasVCg5m2BPX
OeH+gMYknpHqRuXz9MBF7ogVKCbWL5sGS1NPoNZJpMB4A/AiTWhA/Vx5JO3ZAq08
8115+pEeeySuZvZFbJ6ZdS/zZzpNJ9YyYHQWFxuuRjr24YTJ5IcPo1jq/9OCjoEn
Fi59/q2JkwIqhxAopHgcgGlf7rTgzvxngDaEuWkWz4bgElaDHvBUE8AM7dkqKe1D
xdSaN2Dc0Sqq2vt/qN8+lgRFKMFeGm/nv8+dq8ak1wJ1yxl1DyWBGNsANOTJ4I6y
cb1IXykZT3fA3bDvlnZUGoCSPqKa10R5kTjqmubcHdR9i5Gzrh1Z96x1BP/jYa8j
2tMaVkAm4PFhQNbsvzIBq07hBFBWYM8QAfaKyazmRyE5172VVSbRuScZu7ZR8V6A
bw1aHWvxru+BQ+dS5JaIkFhY2LxjxMNQN8Ba+3mtKCKclToRixLMaqc5uNuzT6W4
j9PkQOgWpSZuIJ+WxDuDIoQhxgyE5BhZPNmzS+VuY3cdEzraZQ9+xT+XHD5Y1hdm
uHEHJGZ+twwWowQ3gm+VuXb4bOEVWN6hv+Q9OtPgPQqXDvoraGcYeit9y82/JZ9y
Tk1RQKJJXqM5MJhy7ZY3YgGaCJDNmPoS0ZtDioN0DdOcYP9OZCVHDXyuIOQTQ6Mf
dLDu61A54L9NPAL/MZWOZ3g0aC5Yu3/mLqjh22GNRDulvflEoZiLiFzS73xzHO9L
98iOK2FRIywkMO6oGdy/TrxXXtUJcGgGFUWJ3tptyq3NdyO6/BgdujrenkSJO8n/
whFPd5aXXAhtjagJFnEfSqpzapK0Nqd2YPQXv/hjdC2rH8b6Md5flsmvCYXI3W4A
Q3VZpsqahmd9wNpLmmihYac5/uYezs68/wnYgHO/rW5JPbZtRPqNI4gw8jqLlzys
pP8Rg4s2lJWkPkDe5jg27XMI38UBonuTZCZePsw89U0JWwmBb0gQX23bCstJ3J59
XZ2K6GZP9MulIIYll8RK2fJZe7dPrCzhrjc9WcH30hzhf5DWRRgHVR/YvIpSYYWI
j8ecwpEKtZOJfFE01QpM3w==
`protect END_PROTECTED
