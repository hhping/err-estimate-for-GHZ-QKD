`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Alm5tz51eFju8nm5QFzSP5Yqx+LFBbmD8x09bp8kQZMa0eKWk3/QAh/d9CW1x6h2
TrE7qP+DsOYE1pVlNW8Hzir5WPnEXxfrq1HdKjg0aiglMDIEG1y0g3WYhPncg1Nb
4tPNBy9c52MbKdLvQZzFc/YulgxNOYtz41TVOAU8vWLlr7dmdXHHkNUFiYF55Vuj
TFyXP8bTmSTB0jvyeXQRyd9XW4Z7kuKbfym9GQDE/ecM1PiQSwKjYPJ/xGKVtkPk
PlUJg7jXUxZp/PMo/4tOohgRdcVcrXCew79u31kbWwUNUQhGCrqLsSyL/grZSdK0
Lyvvt9sMIsyYTqUGXKXCz0nthZhPcIm1UhLqx9Vigt+7ye2nbJBv3T35r6U2P1yM
fZ8iZ4D0lVLLHLOYSiOmiO7ub/XH963C+upp1M85cmERmNlOTUCGdcfwSABP/aa0
sTqcLT/jjaMm/gIKXtIA79ieLdHUf3PU8N3fcgA7mksd+EpZjq/SwyGLQ1JXoIDL
Rnr3gIYsUwbCxe0oTrqAZQfGrJPNhRanHfRSDApc2s0ZFFNoR3BZMVi3/coVx6Rp
5/fOZOn5wnsSun6/y2bsWAlsc4Pe5UOStXfzjnRLqXb82T1RDhyYNWlqtEi2Mpnb
Z65dPcPncmJhncHvNJD5R5uVSjCIdLOAwBxTAOl2vVoOMQ4AebipmIO1sDHikWPn
UpznOrpGV3sXWep7S4ExIV5KW/eNy56UFzuKFK0Ux0CT+Tq40D+cJbovjXZxcGpe
BJBtp/FVj6nembWHa5yKLM3Ub7A5E4s98vo8jIAks4GQgoZz8+x+3aSe7KMoi3RM
IZPasbrMqqfIgoM8sCsdg6AMrekWy/gykKyfBRz6aNvBcY9suTIkHc5avbA8wi/Z
Z+IN0FqtBr11g1e1+vOdwwVRHuo3seFITxWrZtG1BYc2EXR5UQSgkyuLHras2Xph
K9n2AZHRO/jBKOpERNmveJEXvcyQLFWeK7gHLD3Zp9USe3DOeQVgl5f3lu5Hxs4h
zph2w64VZ2XMkfDFSnaGM3I0uKr+OVp7+d2nEcJEVMNurVJoamp0BTEVodQKNl2m
6g1gcd9C60Xpx0iy3BejNtUJtD6TbzdHHYLridf6geoVBx4mFFfsbIiQGUz9Ad1d
8XsfrYIz9BfNbyYtsvX5CatzC35L5koroMZWGWyPnOv6c/4K3dQ8AZZklxToryYp
7Ik8erVAQny1ZD8FNfi3JQNHQtsMZROi3mYk5SARbBUFbbFBtBp3GjtJvGiTXElM
VwqM/A8Jf2+DOiNIojPdSE0KQgHy5Wq35IhiNBdbgF+QyJJePAT0QaSIOh6joh/9
6twR/KD9Dye82cWxLYF9y/LvtBnCwZM9ZySO+4KhDYry8bpC4848wb+HgOyjFr6a
iW4mQRcj8jKUa/kfqX8KV2S0/73Xa3pDT05tKSmQGEt4QxEYLeOr6nQLTD8VZA3b
1N5MacOOIBMWS5LttBnLzqe/GkFRdDXjIYnIcF3bladScc6e2vxk1XUwti+MWrmN
mbCGMn0Ox3gXqqEpfb3rjH5twX608yoEzL3bnGaKuwr811UwbltA0MSaTLzI0lyR
y6C13LOklfar9clohOdd9FKvd2ci8+00Ob/NAH6zuIp6Mp4DCa7ZtBrWvQ0vVIdL
NxjPBVUzNC7tjXDgb1PfSuprwpNlP5YtsVhBIcMidI9U6lFS2F+Kb5d3TKRuRRGX
2BUX+vyTzCJSte+ANB7Hh7vCb4aGoHRmAeQg5BjnPPggifCPlCSWRomR+9i4kKpD
Rm/7L2jbOG+U4J6p+lFMpIJvRlgUZ4BA5nh32ofrCzbiymtNHwoRMMvgcBqFFrWC
WIxsEowCGOQQ7hyoU9YX5qleoXhxzO+a6GlsXYTVmS/498SSQcXF+MgekRMh1MeT
rled7umNAvcQwQgOEB6Z+t+NWR8PIQdp0SydkhPQ/4xpYIXOO+IDnUa0vj4/5cr7
3nfNnLx4hjXM0pue5trwikkYB5uSWICGBAJ8bXJ1tP7rv27L80VCnVIWnBUdcCMx
Y+jlRzZjLsvIH5fso4+V0AVQd/h/7p/bfgxZKNf/W5IwfBqqe5Wj9Tz2acu0cv8V
+DvZrGbIzCPiPzgRRFYzaW+vtMtakS3150hUoaDXq7dz03NZLNUid5HCP0MzerSH
6h0E1Kt2qNKjUcSrThVXa9u/te8O+23I9ElDA1NAvZ5H4Vct7Q/bzBwMJ3cHAXNi
WZ7XCPty8sIzq3kh9nkcdS+77xrykKVvtFOXNlYG/Xf3k4O/E+0GZoTk2NG2DWwh
O+g/MeoavzzFELtK8AyS3DM5FN+UF/8Pqr54IFU1RacUjv1iAbmDhLUTFcsh3fBL
sC9BrDHRpv/lu/FHWJdKjwbWR6WHWBtpsYMC93QUMwtOJU9tBsR5P+24K5PeYDji
eD4kfgaDajiUIX9zUzdxzeuA+67FLK2yaNxR8cH4PhPsy0zaMCqXSFM01ZnFPkRs
EWgkv9kswn4m076OWcD4kgOwHqLiDJX/XggRN/Gy7vyTcQnmNuLP4AaqeFBePy13
mcpwRjvRaE3OyKHekvfxj/Jiw0m0r4Ylrq6hnfEHUImU7sZdCuntEZNsbgZwhCVl
oAFoGCnjJmQ7FnqV/UUMp8EkogjUrVcmgw4qmFyPSl7PYELkYDPtnqb/Pzm2EM1y
50siGGr04inTXZPzy8SAmTcA3hFcTLBYC8qzpTO1iHqOuO7kIDfko3ucI+RHKFaA
fjgxOy7basZwoiuSJ9Bq6SZNW/rpadJq3eTX91d9YzzZ5utVC+xksfsOOdhCHxz7
sPJPN9Z1pH2yYme41o+g872Fjz1loNbUzUA2zYcoLvtIQp7cHONU0aCXgvwKs4Jt
2Gk4axbGbslub/7uf3IpIxpTs33iIVvlO7L0msBIQ7ol9WWtbiNqKn7iT4lFhZch
IU5b2Q99vxmVbNHZmet6VRwb7CYAoHEkQ8icsaxzgt2WPC+dJ25FUu3RZWcwldFd
bGgQp/VKt1W07Dfj3jIZHFbmJJhtsUBB0IJ32T/H5V+Gk1O9HN/Evno1qNiYtwli
Eg5JpNBnbxjcje80rm2rIJRae7+AinbB6r7OWK6pI+3G93jWICiezSSKMRUTv0HS
VsBWXmuG14BoUam9WQMn4Y9pBRzoQibGtkNCFvYkEO+Q5K0R6329jKHK3/HeipCJ
RWx47LiNjegvTzkf7Lxw3l9dRgCIJOv50I0ClDRFKnw=
`protect END_PROTECTED
