`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gVUb0DEJNPJXSRFicdYGmS47hx5eSZYR8ZKEvUAaedRC50yC8RQ8W9WV70gfMQ4t
NfSHLVPFhQmXamneXfA+pkzdLfgAGE0uMPzKKYPST1P2c7j+Y4PNZaRauElEyal0
hngcqOd1IKIgVEJk+m6YAPhBSWQSriGl5NP7nmHakVudWjuCSBA8aNxJCfOHycxz
w7AJIHZeWxlj9u/z6MGYl6+Ykz9FLfyINsn2r+PmyMSIADU/J1sC2YTehm0wopsh
PKYqeE69njH9YiIyvPAK4IqoKp/DRC6DkzIlvyKhz+aDGPBqIFcBDRA3oB/3uA0o
FDDwLp/n42RV/5aA5bbbb8sQIcU2ByYHsiK7v4tq5YlI8APS9tL8Htq7b2+7T4PX
BPNu3kZ3XKgFwltuL/PPSVJvPKdXn/cA0trJNkVPi7FPUTTAsPIfaD28KXpo87+X
nkpvPbSlgYeRnVmPT2LjWjd0Ir0255Spa1n9o70OuhBis4/vVUYOgrUV4QKR13aI
/gvVH1j8XeRFdgwZ4bDgILQKPU558XcC8yOom+wKcW13w16RyBPam0cJVZdbEWTa
2HEZMhY2EJEW9s2J9U+6Ncc35ZjyLV5nCsTqT9CyTiCHbHgH3Vs6TFbgh1utJNR6
BqQ2YjJE5QaA4q1KqcpIOrHJxiqb9AfsdIbCRxJDdZPXTE2/ss2XmS8wyXQ8cMKt
eS4djKgfMUoxRQ1+ufzqopJYo4sIa/VFWYoll1pFNv3xiWVdUXXRa75y6qdsv2b0
BbtB3D2bWyWj4UGeLOzXRHqUeZj2gsXhU/aMYIPMZ/Uv8gmk9eAWkguXCF10BiLD
RG9lFUNMq8ybO+8EeuYTT250iAEdNBpUfgkLd17cL1t0BEo2phiT+CkNg2QtredY
P66zl4/lltRbe+uIcP7oy+m5Dn+F2+dlK4kUT7IzWvInCoH9h9dibZawvwToNLzE
wJxoWiYeWyJUtCEkDt53TJ7Y8fxr29DgWgEenBzYVZ0Z2NrFxRBsccnik+6pzpFy
STM9FlxxQ0eEVI0gjgvXnUOXYxC5QDh2db+3+CWtUIfPZUnMNP4Ii0oPas+4s1NX
IzULRL93QGAATvv/CsnuFcccuYlNDEITUL32lUFbN2QvJ3R/iHbqobNy2DZQIBlH
kwl6ziRVxeVc/F0Itwkmiv+rHI2je0lB8GItoq5736UF2CbtuC05XxcNJ6mPFddV
GU0HKd9Kd8wRzy+11RzITvtH9WbDT5+4UzcrHOnt+HbSz2sSMCLsYqRdzsslR/If
ZtFwjUFzjcUTb4eOqo7E4AWCbWmd16eezv5u+gz4tu5a35GalRl5i5DZ2azaePvg
EW80geSHod7WNfWhm432mzcAXHnUeW2JuaGOVv2DFRptnalLRJ1uw2wm086FeGuU
z7oGoQgGKwvE/M/OhdBiAnCUfDzXvF+N38hSuLHuZJ57lr5YOq7eHo4E4zAeHLsI
3UBNAlAk+JpLn80SBPDUpf4rPSVZpRNCaYmkwsvs0sT55x+nDkCexnAvNclF2Hrr
vfnHwxaAY5dvNxlHXloZ2aaiGf3bIClBzoDUk7UZKDJHJZNEhO34k9tdECtaLMcR
1XARoI9GSM2NMfpeywxPTmW53U23Fc3w+RhxQGMaYkN2K+TnEr4EMfBL5ML2SPDf
pYdo3fzHo2zN42JZjfMXDADOVgI6Ci4+m4J/0m95N2zDMm3u/PEjUARXPMHBD9s3
Moq2JV3HzNC3cVCzTqdtkg==
`protect END_PROTECTED
