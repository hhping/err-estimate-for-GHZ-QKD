`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
McLqTIpJh/T9pAtJnjXLOfU4r2wBZqnZReGalN8Dg44LUSMQvHXBpLjMweaC9qDU
fkwrEQiJ6QRtbbWcFlbvjOMNfpMVN1KgGJhBe7CfPn4ggZBhvNYpChzUOL03tdiQ
DPzfs3AFQai9kZU75ZiZZzTFnXW7yqJos/bqwTmeIU04RnemCqrJdN+oACCLrOEc
ZVIwabtFs6BaOgpJWNBjpELaf8eBbBhLZoMBz4FOt+/Y1skWbxuviHpJme/vjnlM
+emZQEYG8i8HgqW70npfFMyjuasPd568SZjtGXnFmw4u//5s1qgiqx+Cu+hF17Ob
nffhx6zO5WuSZu3B2AFEtSoPjbbNcekzaTuvMx3mXp8P6IQgP1vtHg4jsJDJCpg8
eyOt8oOBHwicUaMvDcfObnKV27XxbFsqcxFZ63Vpc6CpfvZvaQrr3hDs8IJ5ofS5
cAx9ssb7GhRYKq2FvQMtKwa8RvkAaRb+/SBWQTQ8nA0szq1pIGRwgaIImKznP8/6
/e4gtB5dplvMOgA1tXTZ8nTLtaF6/kHWuItDBspldPSi4YP/KzUTVrqcE821JeIb
Sn60VUUCJM3eeR1XGkfLU2tii5S8EaxQaApGm6U3mRg7j8yI26AFCVW7yl2zv+c5
nFSvNKY8jTmRu0HwR7yTw+JBX/aNZjVKR8X/DGG+n+6IfPt3mqSX1d1q0DaqMvV9
Yz5cB7l+ti+7NhjiEyqzFIQWUsY0ZJPw/hlYXwllsq9wuJaVikV9EfbqH24E0cCj
TM2i+WIlqzRGbK7XqmkbqHHrRAq2pwxUM5ZBqEYRjtfWGXMd4zxvutuOyDtFBcmo
XCYFBVf107WkNaXd35V0mHf84EGs763Szt+F0CvDjMw2fIiLNHX9ret7ghIpy6zH
5TGR8zxl/WyFSMonRLfE2Ce+wVw3sURD0rzda+A0QP1wwlPGpSWJNyCu3N8cXcvP
xEMXeeUn2gMwIuk0MhFhZAPskqFQEoCBCQco6nWl8Iw0UpRnVT0lYOyLGkJPT9KV
2KP2Y3jjYW2/7RRP1aszBArAkinb0fvy6itsa0lBRMAiZK5/VsMMV0/UQWQ50Ayd
CCIc2rPo+sPX0rtx2fzog+y4YlFfzk6G7S9G+XuymO44ZPJzEQZMOkHfP0rIQHXd
yOP6doLjhFlnltoOMWyndVSzV6IX32LIlkx+cfuH6eRq+nS1VW1OLYu12bBbc8Lt
1GaHb5oDOZz68ZBpOFjfiuJM5dhzer1xDmq6cZv57O3/cPdU9sQPAEbAVXgN5TaH
hmaKDYFyQcrbj7UqEzXzA0BpqltEjlkNqnxhAeACrCuf3pysYlGXOz17J+rEyLh5
mFU28wT2Uwy0fh/XPeymf1QyUrm2fG9r5vKVpiXADewm70A8pito3MJomXtFjrCj
n7LOxicNqKVeAzN1SCB6sLk/4AkXBkJOCYT0gu+7BIouoTPEO6y/RSVQhQrIIRdh
A1Y/v/v8KfPFWEIXddvOg9P2ZMPdBnTQQlIGSFPMnBcnwCyun2w2DgXI1kQKsMJ7
QIjfrXdzo2qi88CIFAUOR7Hth3b9gxB+/m2PMPC+vd/3dOkSlinCeC/6DTKi1K0g
PJEPfKeNFNpYk3Y0/LWnJjur2JEwYcY1Lo9zkE1gkq0Jtqg21i21G0Y9A/851Rzr
9BFKzQUgMdlTew+g4Yj/+lztkhECK18pL3nvKUymK/BzMNJ6vCuQBja1u3g+TX1L
33+cIHDK/Pae51y+r8AowjA4HaFP1Uhxp7Zz+g5zTpCJIWezEI8M8qzqJNc32vhb
GG9jxu+yAI6r20h+eyWQEjhMBHX8mz0sUsSahv1KIYVXAbXm7RF9G19CK+RRt1pK
0H/x1ljFh13aqf7PZxnce7o5ReotsKbR2ViLd6USVC2R0zm302xfocrPMDcMfsk6
GBGcyS9kTw2wqzcc0EiVrqLZVR9nzoITrwDPSRRYz9uWVEvm/RFhHAG0cj0J7iOa
LIcMeOYXTE8D764Vbin48Eeuppo/IpXujV4LkSGw+Enht47WVD8yuNXniqHaphAL
FKUEgds2sTM8IIDHvDL7qzaeQtdKU/EzQiCZlWao4UTZttHH9IBIuAhTQth1CS6P
bg1juPF08eIbV2IYutDwobXhoSGjenXli2rf4fk3UrhXGLXPsZI9uvm/HBbeG5Q6
//p0AcTdxx7AJx4llTFBSTh1/+v3Xv78LiC4WZWr9ea1faMDZ6qMwXvC2p14qnPq
ahZkJi3gl2NvwF6gbPIM7nuRsmuP5JH8f6aaRE+EnysQtmpncUP0/FTrJnajOMzX
4JzBYlVVkw5Ia5YtVwHlLfBwh+O5M3TuVniAf9MnSto3o8S6dlpavPsrXp0GSapd
Xt/s6j4Oq8BBgOprUHu2L7sBBYurOi/DAkjO8V/HfDON+a8bClAP48kzkuJj4iQg
VN12g0dZwzIusNHRsyKPt5ZyFfevejzh1+jgtc3vGx5+K4ntjQoCkLV+j0XYX6Jg
BsDT7+jzAxDm0VQsCykQLokVvtIs5T1YZnUargi/LPRzWAZlqwRY2yC67XJhyBXo
AH+prrpTrW1qOZZhI5wLJoX1H/Pouvoksu3Cd4F8S39h0XK5ivKnwBijwHWH2I7w
qDqJfdbF2DqX3+Lh+v1XsnikA3IGUzmVBDVpBlSB4OLcc6fRy6mYGsNJ9Qm1e5WD
ijqYdnzAjg9ylg4n1Cab4rhjkSIg6rLdj7k8cK4ZCFd8Giz8g75zjOSd0rwLAmG5
D66tzVQ2zRVdQ0x30UkqBP+YTvVet+qxACzu20GUyo+TP4o76jgJL9lvM6NshitZ
WhFyzug1YNZ1i9+v4xHFWTjOfY7eqoOE+C7hjnmTBBCwGqYUq5d2+k/HIte2+jh0
Kc0PGrKEzYSGTeD+2B7IN4uLL/jjMCCR5fk6Ii7yK5zAxdunNnFQluCh4jFu5kXp
hMO/QNLR7ykUp4BanRO8KcfTHsUHY6teKr+uxXALPkIoqmEzbet5uiaul+jnZLQi
1UYuMFo5Yyu+7yLwiw0tGBdzrrY+pFRurAV5ISBjHmTxst8psRR4WP20gm+ifXzv
6dlIC0ie3kz8HnLvdPldYAQjPHTn+T6TeOUIHm8LRpM3CZ38ocqwFcl/CIk9rUBO
f3UCERT/IS6fHPBTrNc63R6sCupxo1/X7zVajZzvhX8/2Pftipz24br5mHu1imrh
p5/QsP9eQCC36a6Uv/sXRIO+ON6RIZ8103v8bD+JMo0m3R8clh+Xt5OIuEYtCKgS
Pn1LIRVb7Lebpu5PZ1+5DQL7JJF99a1KyQCDVFNJlvW8dQ2iaYYEEjOK0IgsUCrw
vb4HKgb1yw+nET2v1uR0hzzL24MplIjUhvfUmt35yQY+b09opSn+7W8BDGv25ynQ
A+Uaun99ZgA329lnp8MsShlG3VVmgmxYy1gkGG7S8ocVXA63L8h9n2haBl2qQk2K
U9SyveyrZe9qn2/Gp8kfemDfyw8+sN7tSpk6AQ/n4fWdwH+wdgu/2TLX8JxSVEmj
9+O5TKmkNAAsSvLvv7vmTk22xuIJDtn8JY9JAv7fwNaqGSC7njgjva2BKy7vtbTA
WdTPtdzSmuPi/xh961dfonfIuPgSx/VyhVL5dD0gSjaYUQMzFJE4QdHqj5tRIMTU
5OxDLWunZ4o5wmfJ7amtuff0k+E9RHYgi2hVJiTK9Yhowf7BUFwFjHtVLOVB9y0J
c/4wrDb/aXOSxUqkCIw1ZJwamezkXap69s3KWBtJ+4pKu07yWb/Md5+A/smv0IhD
+mLdjAIDHUN1OVa5QUypiwvMGeyJnQQWmDk5HxbkEc/NTkfTpi53gh8/q9D3k9yp
s3zVcax6fwUnelSzWEGN23kMGDkNr4oG5Iz4/jZ88oQwhNl/yBYQnhw4LwzC8B3e
MHtWBlQtEbXRtTWAI2OkG7gs1ZhPHoUV7kLxrS0Ph84LJelFqzg0tOGB/04Ffjoh
`protect END_PROTECTED
