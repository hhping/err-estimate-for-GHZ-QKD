`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ON9dLfPpR9zoQ88cY/WpIBVJgDRh0Hom0EhQtiDfNV4dS0UVVlRv5bvFVFXeDAsv
uCvoX/iuSrphy8dtIomPCk1IznrDMoy6XwVcLLwji+qJkwExDnv7lqSEk6UrO8AP
LZvAYF6XIcqJq4HAt8E83yiRRIylzMFmNYZRZie6j97q+OI56e+6s6afye/AmkUc
Yg2+/qhCRk5FU2lnN2btBGhSnBA8Q3h+Gcyzg/OvdCHyZZ57aEaMY8jblZ+UL8t7
nsYXI2cWBlhCRsEJE5vMjQxZMz1CCywHYJV0A3+YtGh6AHxyuuLzODiCHqvTiW7X
mbTeT50bRbI4F5QXD5C95ViOFKO8EYPFlddlCBpf8VgWsFu4k1KkyUV58yB30hCi
bhUjCZsy8Zjw9iydP4YAy4jwGhrqdse3+7SWhZaPn+MCsCoIbxnHeLsXkX6Eyc+G
leMw5wUsPUCGb3HcQtdN12V3hu7vv62gtzvUcZR0zzm+Tm1v4uAV/dyVuFVPMG7Y
VX/ndnae6r+mARBqDJ+jZXKDsnc6rs20JnRJ2zqtM4BMsPQDOmYdzgbAtl5FklZ6
lSQs8mGFwxZro44dwnKoxvPwyKxtm8NbfM2H+EtD0/+K/AA2i/V0iB2Xij+CZIfe
QPBeOcyHkyTI8sQixgYBDilmjccEUN3qiYv3cosDkH/KXCY0Ym8yZtsPPzSfDiOM
3yot8c7Tky87m/POEwyraLlfkFdDgszNqqAhxnqp6YQBR7pFJjs60IuwfV177xjZ
u/MFVfN4+1olXs6lDuCCi4DBmjQiC8KZ3vwtuknh1286BJTin57SPvg1C/NShfZa
XO4k2PAkXnbV8IZDBLLE/l/tSqDkszLvbDfV+LNuypaImQSnKY4ycGzF1DUC1QO/
q8r8bXo/4QOoEQ4NAq7frx7Fdsvz5lwmtpxEpPwyAvS40pPO0PsCDCTHb7aVQtwc
Whqeuc/Nm6Bx7M81U5osf26f1YNTkMXfG6r38NRbUcAeCTEtZHNAbZRPGno5NntX
EAkVM+Ac+gWZtjUWmFYfsdIKmSsI7li4TNG93IgzFOx7Gu7AXA9xSv2hH+tESkrD
R0HVxoAiBCOvqxcYHJ4BxhhAv2VVW7dB5JAC9xWRSpzU3ACCu6YdiaMGdqp4pvu8
PxB3EmQtcxUH/e+UN7pVVOm11a/75JO5pIZkVKVvHX6pMjq4qXF1SNyRHsQ/Jcni
/4j9aL95tgX47bpj2xhhpMD66cKg2pmi+2lS0U+JM59jLm1oDsIpYQWiH8t6+XS0
QHAbmjIoc778+usyD4k07bnVToT9eocQaIvqVLbl4A+a06oy2Xo8JUeL/DrStHKT
tdlu5tI1gmlxOr9m5kPeSnt94kKc2onp+ZTqt6Ku0088mgpoRg0EjecqKcIylSZu
uiWPE4thKXwl+SM/SmjTQ1X9v8h5ZJc7k0aFGmsWMur7plANDbrdEHEG5l0VICu8
mNx+6IlaZk6RbdQogvtAXQ4EFopiKPmLic2DNp9IVficbU9JzdWoQbENXbgxyO1T
c6HK+mz4FbFOjXHEo8iEAcF+pxiSkN4v+2sFxIWAJ0QA8rSzELZKHQJFb6foEbKL
89T7hX0VuTIY4KS+A+7ayjqN9T/y9pC9Ii2r5x7EHQ7TiB2tQqI2EDjwMKGHfOwi
SnqkFVJoC1+KgY+Mgx9AyVw359xNC1yeMB4T1Q5nE9DVqwhiv3bRGdFkHxqEyGFz
aB2mUy1zPc9PR/KG3ubB1SGSnJK0GibNm+NQjNjGtGQMEiMvHpH4OHakF//iNfe4
ZPeRoNMzqCv+pLgvUcQ+jkasWmhaht16DeZxeeIbbqZMtR7Cr5PAf7RQKmraXdnC
sBqLlDlmpcwpjvs5f8ScDlG+h09eaZphb6DDGf9oa8VFSC+56/pYGDYqDXSSIqEt
MUYDbvvPPBNshrebVfn1JyvvZMbGJ3StCQTalf5gp80=
`protect END_PROTECTED
