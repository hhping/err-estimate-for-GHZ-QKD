`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HzIdGN6zY6BG7e/Ioj8UCQUV1uOQnUpy4ESPRPqTKcMoLlfcBL8a4wLLo/K9RcQM
KY6aKSxmciRSJPU9SxiRu60oiBSCcQx77R9157DAbWWePoGurCYHgQGJvUQvJkNk
w3S7ZLXeOGQswH7p6L5v81HMzeGudeQyMFF5m2TpmCv0wAWHvzprcGTJcCGsdU4Z
tw7SQPnj3ulF1tWj7DmJjRx6tVSvB5lP3vaGZj9mLpmUj15lV+1MzqhWFNQT3+ih
U6v7yuBDh5CPzDdIVUXHQXxC2co+hMMRFwN9JEpoHTAC0+XnHjyIYvT5UkzEJoXT
foV6lUHwxs6L3VTJDKyAWWO8jnFuCXqWgvDHq8pbVjH05XoV/+dFIqFneNPgK0eo
4an4D6jE6soVvI6baikESg==
`protect END_PROTECTED
