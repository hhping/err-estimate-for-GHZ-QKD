`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5k7sChpU7QRk66XC4lX96YRQEV53nzS03I76dHNSWybV/kNWBhbTK0PMbwCoao8o
LHUJFsX4Tymc0ob1v5cLkuc+n+Lu8IfQD1inDxSxtqZn7n6NqE5V7iPIE8lK1u1S
vODMku+14id8PzjiqsJOBnYY+DvAYUWYBDLhIKlAOWQLHpRZr52UNRe9Sey0AlvZ
Ghyz3Y9JYA/wnrK4sJzhmncazCfGvDRKpsaNv41kGfZF6xfaCz7/Y0SE8PoKJygn
J83ymv25hFEn2rBPFxTw/a/L2UbYshBqu3p/q0JMe2Kd82O9sxFCfw44SXYzUNUj
8KHh5TKbDvPqfhwJCVDoMsbM5HjtuJtXhoyoutFxcpQA5TvU7yCUkdNUpEreDXYh
xY3YHUNa76NDUIouQggbXxiEHL0pQ7nkSYMTto3m6rrh1zMit0n76+GI1QfN4BJV
wj93pHZSJJkWEf36I9Zoy9FNO8q2eKkymaQ+G7zl1iyj0WrOBHlzoRHqSpg6Jroy
/fm14V0spwVzcKnAbAl6E50hRThzSmgC75VgxKj3fPZvPlC7rwjq6iDSbRkQMQXx
EdUVvFZbejp3WXM3tVB9Hw8N9/vDIVB4PCrhFASmLCe8SXDXWNr7rpWpT3P7BBkT
0mS49OBkjWdJ5QqyBbXZXSaPZJXoZfZd5R3bxtVt+weQy24l0KNFz5LxpOJ11/L4
E8sJIfT7tN8w9csZ9quy9gG31tIta7tRM7lPvWnCcitYdIpg/ZxLj8qaBy9n9aMj
+YKCTYNtYwK5GrNTR1ovsWyd7+xZc/U5fJbsWPFsN0UPpvHWgMkSBSxt7KkhSF7U
eSyVocXSgr+9/KBEnuYNvumyLNQtt3pZOnj9hX0hK1X+fMGGnOzw65npmHdOpZnB
LW9ZTMUw2RwTNPVGzllvxRV/nYQo0HaSn3NwiFF0i5EeXGYVvRwPOZoc4oIZzX/2
/NMSo6NYwxzJdyovPN4/rht0SDKINKRfW4JI5S3Ah+JRP3AK//4oHOjF5sw6cg43
mN892c/fLVwWASGzS9MGhsoLbR1mXaVv8yx+kQQbE2aE9+UbEdeBPFZn4v6BQ009
fU3BEccjyC5VYc4gDnp6GQUrDdQmqpftdpVrRLCDCAbgI/FPELs8rQjhSJqgQ5H8
rRPCo2XrvpoVO9JCf8WYvvTLJkz1Lq8qLvfe1orRue49PZkkiqoW2xV9ktzT4GN7
h2vThnc5uaH5eMBSmYK3cl7ErQxFYAbKmExK9siHJ1eX4ZijrlTU2ezDfAUKsS6E
b9RjuPEmlCyVxj8m2vEG3Z5+GOP0WJsrPaz5jup1yutao53J7GLeTeUMxbekT/DK
d1weKOGRhsYgeHMXOR2g4yt81pBR61KEZuTSICYvT2g=
`protect END_PROTECTED
