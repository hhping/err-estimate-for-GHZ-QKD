`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZBNapxYlbknIt9e2plU1Y4NcdN+ex0qYzWif3N9CEgQ45dz1hpS6TtoQaXKbhmeU
HxRqOmhWUwxYOYlrRzQ6a3OHFKErAhjnDTb597ksQpLRNRDnSRwvXZIbbPpIaP0+
Qzffore4eW0Flh8Omfa50/woq5Uh8Vbq6hx6osR5b4ZigJgt+wluEgxxEEYAMilX
ryYLQ3htNg04QE0QeA6+aTkAGLa2NXf/eR8bjiVIeknyte/R7xR5tKvOyqlLj9HJ
WHRJSPfCaD3NpViILYpVIH8MXhj2XyC0mSWKJPK6XGXraQNtPxtq5UCREQUyAFQ1
R2+SBEWIcLEWnpQLVOubMfuwgLiiGZ1Xw1luIMxMZCZjwvSlN6SGOB+NqQ47nJiv
lvfyBGh+LshbYae3Ty1CI+VMrvfdBSHZDNxVTdBm7M7HUiS38DhkxOAz6a8VXDic
1en0k+pQ65CJ8YAE7JMoDKxvM5JxHgT+/l9opGNcawGmp9kBGG9rtzDDhdBz8SSG
Z/AM5vvO0CrrUfaPaHNmNIzyR6JPlS1bq4RIyDH2psSvQb6hzMJ9vdun9Iu+l0pB
/H0m2aBYg75ygq9ORVDAlzFUKZcdNBJVlulEXUBcsQ8gtkD9f3V0zN9MrQ/QhV2o
BGrah8e8Oq9qxVvZYUPDUA==
`protect END_PROTECTED
