`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fmQtP/YyugB8ldybz8KawF+XvV6f3ACCgs81g0OR1MU3b7hDfAKfiP2vCcatoUPG
utPiTIO/RuFZSxOOU7ORHp6+QgVDfS+u1fFoKZtI7yZ/yhoT9CYCFxbbrrPwvpCX
kgq1O6NJiYelqQHXdOvRypl2bVYOniYSCnEEQeJ5+YQp9HfCWgVtmO6vqB9QHkbd
GlOaJHI2Uo9neEYFT3dz0BoJ9Eqv30X09hu8WwlYapsANkRR7nHy/6KfT+0wyAfy
XMwCFi/68pOON9lSJmYDTZIr8mwj9mox2eX00k7ZrguqCfncuURsCwRkPeew7o2K
3+DKg7Af3BQuf+U500D2PvlSti8y7wxilKnpfC+nCS5xhGDt/e/d07Kj03RWZZVP
kDe32x86jEBNC0/W9635VkKkb2aTAhzADtHSLyCXRjCOC0hLdxA3lHJxlNaaao9t
kBM8YF4gOSngJFw86VrqXxQWsq3+ilS0BlxaRyy6ztzKE5lKv3KLgOgX1hrsUNdI
w2jvAj1vSefui+kosKK891BkRMjFcXr1VDKA3fTGUlyG+ZQ6U+r/9RB7Oo8w02PE
sjD70wQneek/XhVu2I4/pDztwHHS9jMaFnnKefVQwOHoIqYG9rA6g1B6kZ7ATQtk
`protect END_PROTECTED
