`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BYoZQ4B+ZIMRiDec9zTjecTcFLqnq92Xcjg4kpPglJJHJUUzdrKH3v/uV6HN1CxK
KilE8ntnk44fHX43SB4UI02rfuyO/9qpIlasjVQCObSFCI+6aN3FjWVUN+pX69Ko
5OPrhIrm6QX8ZySEnMdqO/x5TdD7GmaOsaXV4/eNJ3u+f+uSAoM34ncPf2fPyW1D
CqTcJl/T3RaAgrIyulzqbMH/6lmuPa3ZMs26a3w/Tyiy2kvKP8MEPtodsHrE6LcH
jAmK9cOVoIupO96DGFigcr2e7duaLdJ9dHeJIGFRIUbrLFVOdOQnKy+fbUV0tMKr
KsCweZTu2Akw82LrFS0spSkpWJe1Vo6VzBbKrGPVSLPxUbLSsMTHewf5tqjKRWVS
/C/yVpZhLuUmNb7odu9NSCpQ1Cy9bPG7OJzwqJfQA4JGsM5kMcEBuEGJC1EarodI
oqJoMbm0Fotcusc5zV4M8WAZXZBWeDBDKBmiqn3JOjvz4GTkzT+WOsO3YY0p+ZfC
Gx+iJ0TgGyUez1K/D9Jr8zEgMu20Z5/wUaH2L6ICIi5okv9Eso78l94+1xcvnwn5
zZW9VdpulXi2tLM/y++bzG2yuURZVKSd4S8nsn7R2C3p21nKn/K6+XkDPRERQMzl
ToPKcMyCz84/n44E54fauo9TOkms7snNN8gCGrWn3hb3iZuVcSP61q7P5vbHyx4j
iBzXm/8IOV+yWg6OiJEkfiWcsU7a7T4iIjH6ucQtPT/g3kAwqvrrPnbiCT/jsPoJ
WgkGkNHNmukRdZdCvwFnW77MmxbkneY/5zso1b94Woy3stZaF1avFIGmECgHw0c5
bDFeqxmCP3JC65JGwdSlF1Eo3YzLPavuhTFeO0g26uiRT9D2QJ4e+vZerVO0FlVL
tHsQDZP+GeQ9exgdT7JeABskN6YPzd4e0mUaW79KYsazxa12hMEPx927owH5Ukhm
L0RCjvFRyxSZo/tjkGqBluZWpc4Rbw2WOzzDHhDKk96uFRZIDt5eQVfAThbnutWE
NBbhMXKLP+EjL2wbwDpSDFiPO7Z4w5Q6nd4Jh1AnyKAoFzHvSeupcUNmzFe9IBwL
05wSBr5QCT6EgdrmUEkXmhzWfbaAE6FeSegIvuOqw/YrAYBxJ1CyWg9eFxv/cb/c
miD6n+rB6lzx+2NMUIiRRte70/42KRmXfzoqhGQM0fih231xXOXeA3GOycN4mre5
cye1ri3ATazFDw2E+51jIhFsqQrP5BEXDvulEHI9CfJ47TeWHZommver5rm5LmRi
PTh0l0jU6mbpxn7c9nz2zztMyyvjwzF7bDyac8CmE6aw/tHAfWH3M5hXOtldZxn7
Q3/bKjao9Z4WwrcGPB1y8jddq1fRhhdQB6oZoQwAgK7IklasrvGhsW6iNCZwsvwj
krq5K6thAkcaQBZd93a6SAEAYn57im/AAFrtPQcwE19MFVxFep/SXVhCpCaXVJt7
ekLvvBqdnB1znbomPxadLFWVLME+FnKgjiETl42KN+I=
`protect END_PROTECTED
