`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3LRhnIaW0Davbktcu8gLm9q4OX6YABTCl2qg3Mx2T4M+E+dfoeruL8INydccKWKS
hfg7gI8sf0C/811rYoWpydThwq5JqM3SMntq3fswV/3TFeDLP14RB0ylFlcovhLs
8YNwJ+ZxsJinNHHd9EKhxsKFof7fH+qtShB5iOb/KXQK10ytBC+65oFgqRKc9u9U
Bhk+E9l2inULlJ1J5Ul0aldUTcWpHRgL0Q1E0ZqO1cLGXP1wJepaNFrlU811EgFH
QSyZft7u329k26JVv+nSZC0IjPdhlPhBHEfZDjTPMcuUCaSnEksTDU3IWlPPmpw6
3+Syxa1gMCsyks4Q73SsAZ3xEVZzbnXiqaOk3xEnO8rsAOpmDi+zW3IPo5q+Z/Xg
z6i8kivY6EzOJvtDI7V1LhIW6kP38G/dVrmqS+NvQ+PVBBJu/ytzAz02B4InSLJe
65DkR1tImTazxome5cafK2ZQdBEKy0AdwO85nUyhLetOVNKRrkxjyskogfAFpZ5y
PJFz75UpRQzSGhXNUb7OzAM0OhZItxVYLnDSEhLxHcgXHbXVUULHWQDWkRMIIpdt
Us7eutF200g9w/p1fE70HgP/NTDeE+Oggwn/PhoXgk9roYcb6F3bmGrWXqQCXb93
rJf48IcuqKwgZ+TV3+E7dBZArYi0ei3tJiLAqAYy85qS6UDO0D6dOlJEd4JRqugr
WAsV5dV7yQdBYgO+wsnuBk/4ibjuunCNzdCKmD0fDhn3VVdyl+zXMPv/kYwnM5l+
8/nuX3rX4hybA9Zm6T10VZtD5Wf4DyBcsEajTYUe5nD0JjIv3sbvXRGipb53/529
+YDZ4tMOGafl7KBqod5osg4FHZh2/VJgAQtv3T0moFOTxhc+EpmVd5Qnl+imb8v/
ARv1uX1HCEZkRyyEKa/Ud0qND7kKgvm967ultdr9tV2YuFjKtvN5pd7+H+7CBNJA
VZk0qgA+HxF/FWrr8pNTck89onfva/Ym6MErh8RxZ0WD0Q5+ujBbun/h8xUUIx7o
RYFkVp6ImIj9cVDCpkOcsxDadz1H7mvzWSAEjOTLcUEgWkQnmjwBTcr9SnrSOSHw
vQh8HbHIaex6E1HHfmFE30WCBlRGolYQ5h/cneRTrzKuQBGOLd6R1OEgVDTXhLRX
4eNusz5yEeEUzCPMzkQktQ==
`protect END_PROTECTED
