`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
moxzxEjfAyw6y2U9sNge1ZDqsigfQUmiAk26UJa3PfUHkLZnS0vWewnb8yJh4X1j
AzwnWtay/jUQfbhml5xrGdJ5rxTlN1YgINt/AT4tbNpR8QITRddkf9MC0mBxLpOY
61S5QicCAfUWHlkqe70foCy+++seZb3bcIryvGrr8e7p8TrhUuon7DY+qHxTGM+q
NpJEd3fZQeG2xK360vVwNXURN62Rn1x+PkD/9AfmRM+MMTI5myzaZoeTEnERw42x
zutfUfR+Ayf/u0TzOwsdIGZfLL+J457rJ9+4no+jGFMpyhZG5IaEzQ13tzTBuu+D
oBLTEfnoNBezVD/Ez8R7Tkr/OPajPchxzR3bLBYJ5TRPyLAxKiFBaDsjv2PX9XNi
aNcOF5rynl7VMffk2ZmcXyXclfj7gAJ1JsEm/lnUubiZ4uoknbaHMRIbKJI9IxIh
ZQsyp6WByUuzoGodZYbzILZBUsruTHUj+xFAjyY4lfXjvBMcBoPkrW2z0f+F8fgC
QHguW87HcwOIXa3QCNhXnALkT1AeEFs/GK9FhmHuqntZEL7ekwbX9lL3Tf+Nm1Z/
ip2t1UB+k5KdZMfZ/6JtUzbnnqAKvWWh+mrbaQ8qvodPY4uuFX6eLPK01yspc09y
y49ckNECvcDeOqPfXGKuzE1TdMo/KYPbJs/PX62vHl8=
`protect END_PROTECTED
