`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pomt9KIysnk/zUYmNeZjZT30P3qNj2r83Gp7GU7ytT3k4Uf5F3bjh9IMNhKR/CaL
7VZd3QBzDZMO8ZNgtiL9+8LtYybMKRjxZR7YP1ycVAU3wH6uzu5fMqziO/2nvIiu
jZSTAHrPr9HjSxJTqzr74H0kFqUTHmCJd+QSU+eQIeV+X+ZnqMAkfp1N2DW+kRqf
PZ4StZ52AxGXGW27lk+nczeOzZ8h+AgdqioEZB4CDSfVj6skmpRl/D6qfKKTUlvv
DZDq7sDSj1DwaFAgtDMvz/+rpZk6lStipnxw6Mo6tpYAMosA4zoJ5mM/manHHmh3
y9vyuCcKpcBuhcocvhqhrLgRqzFVYwrugT/psROmm13KvjQraPKoDxeO7wlLrGvg
286UcYJJ81uxq42xhXWVRFmj0dpasxAqVXkWV+Pv1OBOpaMzYU6PcGkScgiM2Clo
2qEqYy0mseeiXsrIhu4Sn43a6UJK6ImLjga4PJ2sogOAjstiueRCkOwFBqGyfzCr
63IbICGYYiaBMbqkOLekIZvdFHwf6dA1gvSYusdVfufTzThbySGFjVUceH5lZTk9
xGPtuUJjEBkn2zvjEpmVteRepD1ekhpJYe64cIu8v7AKfxTmb8Rh7NorOUz2YfAp
d2txpvlN/juNZV2GYv+LGGFlWdxKxonf3mCF7AI6RNKxaskxXI9hA8bhh9ZQ1Okp
zQNaqIQh3zwrIxmce6pFcnPTrDkU72jSicexgE6FuWRCsmLy4XBQVIsr9veUIGJS
daPG1Bd5V66oOyC1E9FM5LBMlx0xrNUQCxm8rCDxVUxv/LMOJOZ4eeHwVKhIOrMo
eClf8IwPak3Bg4JxjROUdhK96pVnfyTrqIEEVM9OABRIgLlKCnU3MZF7SZwTFrJO
YfJ7EkKHhZVBvX5OEv08cgz6VWLOnwGV8nmdJLfdn8f7GxeGHXWbjv03pAuPuuhg
mPn4/vh3mvN+KoI/YT0lA2T6FbihRtXi5ENsWk4ynN6+pacwriejHIZRMrcrYxMk
PfjNb8p2KPNsIQItAIZlH/BiDaLH5zCWlDbF6AcSoG1kiGxhoAHp8rCuqOt7gvh4
F/rGn/xX7fFkhpnj5Ru1MajDMSxH5bn+QalWPti9uMNVgw0vPxRn+0g4R2+cOEoT
fNfwn9nDrM6OH1szmWi0e77e/HWGdLqMhO5ivpOJsaq9C5HhXN+rC/nlZiApxZuj
vk6UZEPJXrM87Cytoj91MncgC/FVLrM99t2gsKwW6F4yymmqVYZKx7qgNrZCyyWb
6BkQVIqlZJR5woCBuMJF8/RpxRl9o3zkd6Gr4RmbP4pHpUpx1mtaPsTfCuqXsHku
OeAmRWItgHGZOnLT6mBqkZJhh/zj6AFXWeW7/OUpg1rStYIoL+UT1hxDtTp0G/hO
ZoDTz/lNSNVnSdS/15oh3/DZUsHar4bcOBdLs1ZcnQOsHA32vCZ4Mqwfs3KlUiC6
+IUZ0EfA35XCRYv0CoeU75WGusEu9i+DMqaTyxVTMMcxJQ8HqpSPjFA0vTlAGX9m
kq1WrKdlqpJ+2OFCfa8mN0jPjOStFHuJ+Wk/vOmLVUVGa1fr5dp7c8HxXdJCv0Hk
wYd3C5FMMmPTucCiTioeLn9I2d06VLgSzUJ9TkEOnBQgLMzzgQig7aIdYEDc/6of
ebNxoAC+9saPChCLqeKeZPZoHW7uMm10OLdNkpfRRXkCUDfrVOoNn/Kk4gJ5GmCZ
K+sMWS4qn9tuadRXF1kZByWG/a2rRIkHBx+XlcqkkeCCXcPw5ZSgdfORRu0UPjvL
MIOXz9AWZ952iDG5tPhTj4d2ZTP5djDMDP1HQTimCGMKddyeHqz17BTcVFJu11bs
Mt85rfqK4gzjrTASyNvBGOfyx4KEef0pSJfIqz7LksO5njJkKEfnApWc1UVBYweJ
gdqkiT0g8z0Nbhs3G388Hi/rhVY7H+RQBhS/GP+2nHG3iPvgVCpgax1yIRd6goTO
/qJ0AEBznpmHz1E4VuA6ZPXXTlEeYrstyMkaD758r0sjnKPvk/f0A3RmJcKSZlEy
5lmfsLlY0LgNFLiOujN0XSpaT3kUDiOtnZSWLnPXnhNuGXnnq6MQ8hru5ELA4Dke
t4e7bNzjiAnKKNwiLhB9X9VYV4TyUt76k8WCUfLivHeiH7N4ggXTTslQcxlO5zdt
uWCOEiLimXZ8ijcHfJyAja7pt2oN6tylvn/qdp5I/ZgsOErIvNoP0jv64x9ViPWI
Hx6HRbEE+yrB3b5bOIqpP/pfgEPb5s8Zizaud38Eo3qX/yIH5qqkCd+zxk0Dq2iB
HBX5pYI8IPBafJIs/VZ0O5k4IGwjWi1dFifWC6axK31hJLyawYH2yK6a6CmoEnSt
GOKDWrxjAhpAZBy/WuJzd4ILowRvauUfwwHUwjE7o8UBL5dBCnAaHTwkdzl8sOii
F23cFSVV78KEJbRPTOv+kzIRo6JA2JYiKVZuSwwVb1ThJdY/uTOAHRWaCKYyIvV0
DdS3u/AnG6roDy8GgeNBBOKKotXNhoXziFwbCmOW4jai+mwIXjoOSjeAfTa/9lgn
F3Ba3V11tbdiSQyNw5NCl09030z1EZnmcyeTbCXoYU3OZZxlMqL2Fkf0gVL2+pk3
5s7+fWXxQiE+wzygzANPtBUjgtRF/onM26lLsA2zVfpJn0+7TWEqp47xyil70OW6
HC9O9eh3LSAvHUkvWKxlCKUIB0nOYoBjp2YL4wCA8jZN8mXmExsk5kDA+//EX8uK
Wmrqm6gXldAh49RI50ldZdNUR6ahPOhGZPTqm/g2TAkpZmxB34aoYm0LyUJXBcPL
l3C0ymgUGL9PFgQEyJcGk8nbOMuRcWoWYFrZLWU5aPwASN1ZslV8o9S0zd+3j5n4
d8znSxMfgH4KbWMAakBJdE/jJsni0Ez/WPzZMTGj8w2+lPktRdB9q0yHVmmoDGhk
wvMcBnXSZ6Be8j+4/PLsi2p6GC5a4/+zzZJqVeDf05Kz5xc+IG+FzOW412y2uwtp
pRCsmKw9a6ZRdmFy+lSu+VqOLTzaReec967sowl89QKqGL1oXJhCTLIWQQg5TZvg
p6xYwcnzhoDLrc3mvFX5/GBNIUoZQsGx3DTlL10P3+ixSH7hCs/hdd985B0tqKai
VH2BiC2TnGQZ7/u7tlAOk50CNj9QAhMuwXjLa+dCgrE+ucLNqjar/9u7K+DfS26x
pxHECxGom8rI5dY0x+SEhlOwDCTZ7jFE/ZLUhDG/Yyg1inlZlAYQbB6oauaUBrIV
TJ7n12EAbPKmEqGi7JUn8yU/wAwY1aMKfqRn2kAgHug=
`protect END_PROTECTED
