`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tf67HDwDRQm0k5ae0Dhf3xD+xpD5B+paglIqeKGrGpM7PYJvMg9Zn4/jHZszfPXf
QFox3kU+C/zcwHGfU7e5kTsYQkSdmiD01JOp2ujajEq2e0aEYVYd1ldXkMsKZphq
IbJd/0oIdWYpKKDUZN2yycnCsbGd9b+eOqUpoKPgB6r8FixK5jFjhfyM5DIydwuI
7AT/8h38s1TRYcabEeocghhEGfWN8cLlcqE5TSJFtvZ4vmxVw9DNOteK9N6mH4J3
/0OonYNi6GxmoNyeSzH5s5XL4Zi+GMKbcCRYEQMWLXC9IYDrrt8AVZlr2XS4AxoR
CSG+agPs5DYXuavnq18HHqitYN1CTOrCS2TAm3/zCw6GbAdzMLnmGtLcox2ixEQY
Br6b8YUWJlsiHpC3AHKAoLvpHNzLjQZK7yACzQ6WJOTOkGcf1XUmwaKQgubc5+2d
4deN5f66ii22A2a4hQzJA0ay6W96DTA9pnzNzFl9m2xM1IhddvBtHkY1TtFT0Oyn
8p9yPH0uwpCcHaFjLm9dFRapXMV8Ps5ucq+8hDR7NXteT4ppDGPIeSibn5Vh8jUr
hkC0PonHetVaMMTVsKC7EDTq/kz4U092ksNhaIxwc5kUxHC8gbIvefWnGa7+ZzHi
2tKb5SftMMnhmoknUlSZHPH0ZwAX59XpoEY0UNZ9kth/IqTBJKV/eVP7uhFWchhh
iblUkhOXDVRYYFiVi+nCqLoF6AzwSTbwiypvW09jJ/i/uRECGihRh30HgUQmCWSW
14HgHZ3MGqRv/irLaaGLXPyo61/q94ItxYYCJRpAiS8OZv39xZu3/iLEkp6zDBbV
4xkF2p0DAOf3Ca655n3svKXeYW/lyqEzqwNrL+NKHdT1jjskKraJFNwrnoQGQtJf
6aPGluizcRCO8Be9b3smv9L6dgubS5kCBzB/AUE/h0Woj/Mpiq3jErRGQSVIo2+s
DPYGUacamY0PHYBkdWfpD7QokFEOi9wUfapGg7BVu+/b3nNQq2WA9OYi7cECTVuR
6KGDdHHoWAjNKvrF9u9Vuy6xCwxSBT1u8xWh1ydT5mv+6I0UTNeRQ1LeKDMmxI57
fvLv9iwNb6ggBr5wxAdCSYjTuHSfoy0d9vpAJ00jryLeXKotmcYW12NPRk1aI6R4
pSXeyoGnhxauuK/6J1PocSJoKVzctWaHw4osIMiisOD9Yz8dNoHFv98i8vvrSXfs
+CtTt7q9ISRB+9sQsPGFJx73VPVuHL5hBN7Q56xpZg9/Lm9JHUw0PoZ9Y2JRpKgl
AqVWR+OW+mfvQoOS7iSJxJ/mOiOnpecP79VTwjDQ/Gh3xvtrcUoYqFQOJVu294o0
RYiHI0/2AdAFFQ055/OcKyxQCS2xVd5Z27uWhY4gxZ+QI7w5An2LDAKAL31dzvR4
M0n2A98cMftnC20mgYgYpZmFVYQNgWNB+KBY9fO+A8buKAD+BNz10DsGSu/s6l/m
FNdlRsTGqVStPLolQi4oKMfffn5IcJRBFvyrdNUG0aExQLv9gMBszqhLcNU8KLWy
SqHfwHXWOTm/cSSrkA/Sk1AHcYNEOvvvLxOIOwhZ6RUdfgRQ4H7sjRI24BKrwAM5
jw+UtaQ2/lp/muWP9Ag1689gEMwi2LWNWEaAlfhQn1jH41zN4NJig9jlQplVw4th
0v80SxtPrkd5bCTduAr3fsvIJ0ZO3b63lf25jWdLwPGAMJv9K1A5avbrK+RCL5ZY
/cSZd+3phPTmuo4OChCEq4WCoBm4CMk1kLu7FlznuhzWwVkciBRKKbb+bn5Rq5cZ
Y1HhKUNWWX3yx72fzl1dzl39PDejL6w4eEdylV6JWqEangk2xM/syo5bot+aKiCC
50ge6VCeETGor/QbBl4RIbG6NECxFoytu3ewaz6I75gQQYhgks2yBzThzurMBp01
eYuujBWkx5ATTwOhpMBj91gwA2L2c6StCLGnxDWfK3BcXXBZ5j/kaSqKOaFsnvfu
2ROA6IL4Ods/kpY2mm+uA8FdJ9ul4tehf7NnSRLIbxxkMIhgk3HPvl6NLlnoE6xu
d0XOSvK17WZIZ4vHOr+ef4dEosB7yJpWsSyESa62rspamKfqQuiJXEg78KJSd2cL
s1UMFvNvoR2CPNWZjmHo1KZlCpCo4p3ldTfwjl6OZs2W+FyunnAJt5jDeAe+Ab5C
yOyUW04CilmNgDg73zrqyK/KLTd8LlLRL9/9vQO1ofTPVVHX3FXhuM0zlg1Zwd1B
1poN+OlsEmAQxWwfW5WPee/2V37k33qWuA0HS+f6geEpkox72Ies9kSDIFROnOHO
lSe5oE7ZjQimniXkY5UFxNVmAGbbMsO8QtNHLcFyuA53gURKmzMMnWWsVejltvIT
70Q8W+VgduXZrfA32effZjCT35pLez1H/yZq9LLk7b7IqPOJ8BhJpUn6X1JeKNFY
xRiOJPf21s6ZgXo6EZce/PIfCcdIw/kS464Mo7Ua0FGvJV0t1LbPHatQ/3OipLzJ
eqDXI1qe6xkXBSmcJEhB++yAiBDHZ63/q3B/nwHT8zHkxzY4anVueVhe62zWJwMJ
hwEHSlG0MlEUg5oxOfA5YbTj4bEKxQyDjxnz784CawZC2t1I63Zz+X8+mEwuyUUT
AnpKe9TO4VVfuKqMoLj/dbVJu7YOU7nPpnLkdzLefh6MZyKlFecQCF5xpGcl9uFb
AaNxpa5LfhLxEkqxiXZALOBxc6k7emrsbisBj7roigRvIkVZMFvXHRnYCXbhrQbF
eoGdUEuP9+tlg4ND8pzyoP98ookwOPzILkOZTAdWevGozwk16PtO3kyZleRgQmFQ
FKgsfM/zFNmKNhCEbLKubuUSoxWN6XyHj6Ct8AfHPhxs7qHlU3MRjH2jhGbwFWP8
6K5T0kiQH0DlN9J0qSS0aJZtCF67lEPBEPCwLLNvYohPGyZTWiu0MPXDPWk4OEmv
b43BR7zNhZoTAEvWgHoD25IqMdWub3UBY6arTvGCjx891F/0aSbLLkRE0AmIT2Ud
CZueK0jBrQmzFYKqKkNwf/sRF+W/HxL9hTHyCW0+IlXafU7kbZVr+rajvAuNDZbh
Jaz2DBCQmaM7aBclysT9avwRu+5un3GimsQuyvt3J+JE1t49Ggy3xMWLveIJrARc
dMCq8P0o7KucCgVzas6WEF0pcNL5osz5qofDBmdf63rA6IPoKvVGV3Y7lRGPAzAa
WOjUpFfy/DETAxeftbUNECRV6f8jyu1UCvtGYLClmHGLjMkpIDhMno+nnj2TIcad
lGN5qR6NPnnXp84Ho1uMPoj8JLKn5iI5hq5d7U+S4Qw=
`protect END_PROTECTED
