`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wsi1SPjWOiysngLuuSLkDs5uQgeFrDM90c6AHSBHEfxgGwd+UsoFPZKPnewwL24k
jgweQSe7BnAAQ9BACWM5yvEwV5b78N0OWnTmqC4TcqxgY4xQ8Xtu9oSwkfto3tK7
Jg6WZz1lc92mpsH7KHbwQDAnSEYVZ0fFTzcUpTpkENs2lVLZkF/18ARlzxojfBMD
GicFPa0YxGU3yr6EQPJ9AJNeOrxGDQDzWM7SDHnDqcvbc+ZxCh7+zEBC2W82ewFp
6gAWfCCRCvRFPmhqpYICkh40rOqT3+yJ7PoXkVHpiS//DN/YRoAFub0vRNeOpOYQ
FQMxC6jgrD4/aFkD4BLdUfO1CnW9bEK0NMZN3CsUOIGzSNmfBO4olXCpvuTVnwj/
l15IJ0KX8V6DbPZqwbHXA6/mpvIaBDmipn5JApWqGS5M+zYc8hJyNK4i/EKU1V9O
P3eePg23JKeeNRkKm5GOXpPElzUN1MGMrSwk1G7SoFLExtoaRcbr48rT/izXUl13
XEfe2fdUY4IKcKFp3zo7p00a195pjbVu7goSa5JXSbsd68yTwfM/hkZx/7qtIZeh
rN2+B8wiyqigldVJHFBgzNt7d/47AUlKQzG4PZ5GtouqFiVkeZM9QAp7CoiG7zlj
dzVzTmPZIpNX1iZxYK5+ub683ZjJwFCdei3Q3CRPUdqIkOtoS1ylg3sNd2smSWKy
r1ZQUSvJBD4lSqOS2N3Rgc1LDdihfTnLqNKDNx3prVoftATW2kApfccTDzFSwKS3
6AGL1h53nm5Uja1f3icEXOgQ7ztnCNDUP0gABjJ2WQGvWjqfGGYvtn/FeQK0FweV
R5/5B5+iR+GoKt4j+5oIdw9bx9TRJoz/CAgdwwX8md2H0Q4e8w4DteR59ad1gIt7
VVnDTlppPGlvPmZwKuIFT9uURx7HalmA8gJtSxFee+vvqQkMxHYCmLuSuCnceih2
L+dmsMxD0TELga1wdMXcokcTVtrrNsI4o6OtW3JEzQTIlN+aoFaV19YnjSnXACtO
OOK9WmkoI+cIIX+D0f2k82zgfbydFXYLSbAakf4TAN8/3SlY+eP+2E5TL8R7SPJZ
jiG1HMASe0tqAQHwcdXSIJ7z4JaaXotaiM4cbmNVA8wHUkrj2dAcgj/1TbAbmpFV
P54allCmMt3L/AHd6cIZ8uA2uGUHpZgxMu5Q/+pRleXCWcEzxYHoVFUcP7pBIlkr
+HmDp+dr93kAmLON/6sO3EGvkcjFC79xPoIKqJ81qLyR5V4O+vIVIw3PWCR+TZUl
biri0aC9SSf4r+UhHnfbhCE4WhkJ5WSwqE9oA64JFqgeMTUh9UH96HSMoYUQvraa
HNXOQCknQhV0/IbpEhWf3h+T4QEHfsff+4xTsE/i77elk0RfaEXOwzSvQeNEVEDg
E0BgPlGvzPtqfy2f1ctCaxdvjAMYac2MAk610ByFmgkgNctnS+afNX0W4GVx4rqs
nrlwjw3sCDmbPkGf8yQqjEysUYisu5vPvJTktHYrKwB+axaVYCB5IZWq068aS82f
wkZ39kCpajJLPpNFAxdjJkdjQwilhVMt06SxNHhYdABOYECa90v8794nKjbhLexT
s2L6VeDUklqeE6TKclXQyeXvfaUG+A07RtKsru/R2ahbiW48mM4FLLkQPiGqghhg
lVeb/6pSDmCSVLPhBYId7yhW5zWCr3JnSo2bkN68H90w3uKGfdf4gPJF4iu+jecs
xmEiapLyKLvICj/IesDA2NpY6YTO2Mj9l8f9loIOLw/OYx6RzHm8Iejc0kQBK0PP
KB/UTOXhUvwLWZTkVheQuyggNGdpN/bhn0BNJjJRf25aOcSNnRuuhr8cyBY2toZB
b2TLtbY8uppJLEXJQ/O6sxQsaZN3JT2TxMCUQuI3t7lIKTwmqoBmlfwacuAazpUw
XQSeVKK3RgncwvMKwIFzbg1I6OfidYubFHXsD7UUXitLtIQZ5hV/row8FizWnNvQ
Zoaa+G/E/OPF8JBvAunDR3q1C/ezVX4thRcSnO26Q9BkWI46lZys8AiIeY11xs5n
0cb8v5r72eWhA9nENvEdkBQNcNrb8MHqYsT2IATA1P+MX3CdEzhMzVGZdIHU4C2F
UsO1dXgaqrNJdjyWqzXd9nsrh2X/pndaYRg0DeKG/csKCqZBkQNqeRStlJB4R+Hh
O1S7G90jZzs2xAT/LHX/QZAR8+W+dP3q2mZGo+FK9D0r1DoPZQE+58oi+hznKxCt
O20zKE99swyBU92zrBxyqVAl49bfqwv+fIMhkW3XKJAqS447WFT9B2RC96rpdNAQ
/BJBrRtQHLeWzXUsuLDMtBiDEzKcnAI4FoBhPrEwN4QvRvBR4oAieGdiADt1b5oT
QWqwHqZ7a6rS2mgAF1bVs94UvrmEg9UrqYMeZnQnq2ob/GJgO06UdjzywVQo1jQK
MyEPuyuLHmKsddGuLsIe1IZ7DiVOHxUPEdZ9LjzScVH2Lbb0nIu77a7DEYrizGaC
AOboq7jPXcpNCQfvOdDHN5G4IEGVZVwS6EZZuPjatcf+/6VF8FB6iDUAbd8pHFnD
nq3LOurqT2uovIub94cCsiP2K5seMrovqfCW5Z6MTvm73p4YZo2JXiKu9ULJjCwR
dOMpvndtlCo33Qk37O9C6jENHql4+1W06U9/o9vN71R+tpmYHmuWPX5iTWGVqON/
MeBUXJDRjqlvZse47id3V1xoEWiEW/WNWWyTWDenaJF2G3kH6nzoJX03q5POiICe
8Nq2StTKLsRsSYDW+tafkMlG1Iri7ZkMMPa+HeYNvHx7RbHnHkNPus6UFlSjjBlj
PYEkHkHhQxR6XXn/TQrx5apMTMyxIl0I2ieOonu3V3pO+mdIKfCBywWWYhg0Uxuk
FKqn4iBNQrLDgAHsV7DyPaMAOaB3ah1Hn0loRw9uu65q4tTCGOn+7rZ3v/7TNXXg
+abTwc+CBKbkVrzWL3Ezirg+j8R6ysA8qzIlYIoE8mVTv9jSQ705/o/rZPIihy/x
WRbcr2HiadUZVAb8w92I/B3xjPdr3caXGMj/gaH0gucthbgoghU6QYScoWIllVWF
IrNKH8yD/UygL+4ViwfjX3yXWqi8QJnNv/IAYfr6D4T2EEJl/kGRgUukfZPbtCTM
LklXr+UsGDGbiQ+mLNiRY5ZlaOqsTZDIaXWLi0BBPYwZU9FfQ1sIFZI+OGKhySru
FwH4VEMnZaMn6TRjDJGgOAGyfeDA46wsg84RVLQvP5lE3ug2rIQ9H+Fd9cCA9IiN
jTEGTtrIKqJ2C/mzHUktaqOpzIs9dgmMAB0Y/g6Q43bq/Ekv0Zp2ukHRQsiFU68e
BJVCEMYREIHnJVlhUDKEmA1Xto+RuTrmfYV6ft7/VqPgYTqP8Gh47eWA0mt+dH1B
PoxkbFRrMa3CYJnJy31vIlBOC8XL8VCaa/mC6LTzFJEl9Ds3Et09drEPa41HHpbj
5sKSHo0oyyMgbXUNrBazwzDD0wfZwbJRBpZe+hNOs7HNYCRJZCGRvtrKPHnRtsQN
bBf2wDpfdrhwNnZdlL9wgfQMpu2+UXRsUPmafcAXr0sVDLbI3f5euomv/HHBA4WR
i7ph2znd6qjBFV0bkbzrV/hWPAb4/6VJWjW+hTYSk7uHWYIDQWLo5MfSVBVPtq4p
/fC8aTOJzVpDEYuzeUMaQYLwmgDONEF3QczcmGwL3+V5afl7RFFfxXb3pAbxBVqw
EBMsws9GwcXOlp2fGwqh6wnIrGcnehGLegE8IgmjsN+5kQ02c7SuL/QZ+Pxjfa2m
gQUWBuElO2z4CAFI+d4lHEkaBK2Tz5viUNoCex3RgqHn8IYGOBiZKB6MF07/NSRr
tvE5Cq9ed6l8Qwx2t+Q86j6+MiprmeMvuzLUL1fpzL2abEUIwUAlgMQ5QWHDqwLi
kVAcOkDcDs+o6Kzt0sZVeURfHzAuQCcPjiioVI/9utHYwzBTSOGS9ZfedX7Gpq8M
2Io/1G+qoSnHIPw2gzoDdpHVTV/QNCE+G4oJgt+5HZpsrwfjBOF6++dR4Dchm3Dn
/oBnqh/Uy95T3Kaly2V/Q0eB7h6hQ+diQCtjmcyACOoh7z/6ecs8K8riuXuSIsmQ
d54OoCuC2ntdOauYd4mSbzw7Xm7jE5NVY+ROlivmmTbrOKZMTkWfzbH4hoBTG+7Y
GEfA71aED16ATOdrSGRx1kfUo+yTxDHG518LeOqdmzLuudUWAy2giLYzTZzWjP5y
t0mjfX34/WboQwySKguaMKDR5RAIqcTTUwLdm3mGdCszr6g45aRVoResSYtXw3F1
PC5vde2fUls2vAFgBYYnbY/xNJ9D6rMRlGpb4SibLXkoM+ismy7K9/RADd27c4Iw
KLW4sjpr0706mgcFJXeAznIgnqKrXT5N3dOfq5eawhxXyi2CmRKQuGDWSv7o8f90
avh/24aQuRBkyZvNM3ykghu2/RmMqGvf98DfCOWhewTzQ4nnElXccoMURJxYKFTt
714xp6CE9x/MPqKij4IVTeY1KtPioB7+JnyAD2+s035TMpHT+q1ApnV4T/+XlGaK
QdPoEM6nkjlQedXCREd5NTqKQhsBlmHDetBev/A4UloRMEsxiqmR1GycbjwvKpn1
UQdoQdgfEpd4j5syDjIe7tjzV4X3w7W2PI/CSG14tfFvhiifDGNtckRNbM6vmES4
ovKaVtTr7+lWw2VSZ6karG9ekLEZ1S3oWoNWIPXN53VSFx9r6W0m35Czvw2TDkim
0hNhkEWwWGSZoX8P7RbOpfoRv2BJzI90CNCEOSRUWgA=
`protect END_PROTECTED
