`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MyWS8/WILYQwEQKvh17KiBzw8Esy8QoZw5KgW9bxgamCPWZKIV8LoeIhcGfPyXIg
d05j+xfedwnMq1Hvi8iuUzfxyJ4Uii+c5mqY9tFTJ2QW2UZB6VyMtebqvRL4M6no
RC27TfeFKlziWXZ/PU5+THmgzqOaLcgteHSVnlzg/+CGSUW2Hh6vfDKKJzWd+JZf
lLBaaESN67ywjg0rI7dxooqbes/QRk6BWWxZTxygtYVJdnagvNSOx6c1Nw0Pp8Q0
vIyroDXkYfIQnQE+xSkImP/EjKPCbvp+BqIWZj2DnxJeITehXkR9q8ozbpa4JTXL
7cU7JOy1JCACTiC3pFa4V56+v9nCkzYs+cYRH5Ta5B/v9LfQUKhjjzQi1TiAqswl
A9QjTgkFx4+ED6Gk6Z5EyKsD5ujGju87w1tMj3Ba9gjuKGhATc9Y/+JK52g6thAp
A9s55kWQu92DDET+FNUFPHxQ6kCBBvo83l0iVOD0LLm8y3e47Nc816P4g1uEjiCy
g5LNgvGSVO6E0qXF844XlUshKi6JRTOC9P+sZ+B2Iea3DGhxfExTNQeWeaZekcgm
085NnwVK3863wEEcchw9hj0jY8KYgnGsnoqZC671FMszgTRrNoZ/PuaQRwp1iTcU
`protect END_PROTECTED
