`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H06eIYi50NKC1SrJnvop0rZq/QTckTcym7DAFDbwr6JRdeqhf5Lch40z2vQTzJ6M
O3Y1mOcg+l6tbrYPDjlOU8lY23MO2ba+BfxXvZr9gSEM82BF0ol/I+ladhLQx7Ln
tm4yhzkU6ud0Kq/ocSmgV6fhYmNawlskv43JU3uEiE53xqTMfPqVyJw2xuQiMVtk
VdLaYDO471Os/kaEPgnuGbXSH8CLoe9P4vjEyrMUSodoWSveYX3+lRx6R4/iBgk6
di4mXrA8fd+mVGIJ5r4+YOvBWqMb2mS+4yn2vDpFUdJaDXRiYGgN2eqysEq2KjjM
iUNmU2IlZV54Ctk7SPMKtdVZZyzTDtAPIXJ378iBU7i2ms1QoWXwte0rmksrU7MW
VyxGI81EwY14J0RztBEPIczEEFs249OpaObTvfQGzgc=
`protect END_PROTECTED
