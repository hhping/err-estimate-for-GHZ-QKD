`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n6/SEguT6E//+eWejptKQp1bITp0cUMcAmwY6HzP+t1Fn9IAk9xNcSCILlXv6Uov
GR+0qQZ4P+Ktd375CcGT5V6BIVRZWlPJejPPoV95L1605igQ7+/0NepiIOQWEDtL
z/rMw5DtJNZVKXYf7ldCz4Kz1xYJgEJfrSw/xXI1SN1ejD5IrdYgCzidDewz2KbV
Dqx7/79Z1GIOqobvilDwSdWCTsV4/CWe6jEW5w/95hqPvkO/Dzb6tm8NdVIQ9DNU
f8UazqGyuAP1f7C6bMGRv13e/sCskxKp45JOH8eI5VS8ACSUvKG+zS7oyfuxpufs
ghfJwhetJFgGseldbUL0WEO4E36TkiQ9XJA4AxOQ/1cYuBDigonPLbz8Fx3EYj7O
F58AedmsiCYiD1JRLpQ1oo1blJCDx7f13DYe0Ble2au1MtYeRe4D+1FsH4XHBVBs
AA/8lwC2vBGqd+8kZdTZvQxOfQvJV7i+IOgGTKDI30dwXRLgp0DKb+8lV0mokBXQ
RBklw39yylIfFCtV+IG67eTxBvNy0oZPYXCqKPAaIsQZGU52nyzfuvrqBd3qxsfq
cZVPvtKTTRDPtSxZiEziRf5OziX5KQ37uP2arqHpg8pCaPBPq2oPnLzVgMbHkUOy
B4QdIU6zB09qICwd38BCqTcgPl/ozBLYL72r5uPRNqkHgAODB5Rvcv/M0Esidxpk
o2LUXaRlgQ8akBF46yfWDkm/EQq9lbTwTm60P09LI+E=
`protect END_PROTECTED
