`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8RDUG9cVXTCu8euIAyh9Zeet6Q1mZT11wXa6CRdshgYMINYAUso4lyyuYecwr9MA
A7DyKhb/qrL6+/NGm9NCmVUhqahrMqH9bSGv/7wwTcN2SXQHD/WuBbLCkHoyImit
/qYN2TfEWtd0RxwnTbD49ZUwa0CftUj6N53nfZucOImxTvFSzAV4xVr/jJ7JU6YH
90EYHe0Ps3V/n/aU2lxEAqC2Tbh+S5tmd6ZdxEXCxNVvGUU1BW2nmRhTU8SpPZnV
+wPaSjorpQ6+T2Ut9Mn7I04AE8DV8QnGdt3+ediui+Z+HTAKOusLyRd8zVlfemCk
txBEgyGxo/OOfUlScEx9wn4921PrCSsnCJoSbDCzTnsydEEBhChkzixi/leYrLkR
elvIHZfiNQlB+TnyBbDZUPComVNuXMcEkUNt+s2uz8Z/f2TBQaygzGtB9HPXGpGO
sHtHBGBDqH1KOmQidgxK5uGd/o7jAQlVZn5fL0Fjd2vnHPv/2gKYIPA1VMpIeec7
aQKqCo7dBtUlzdnjCGIKZYK7klHqPrOIR35448QZ8LS+cJHy9pxOAWoyQpRMEWz+
AH/NJrF5m0TYPYuhoxJjk0iifVIw5m4FbbcPzQ76QXJumfCoSh8mM3waYgTKwruI
5d90RGvDHao5COP42GUdDGq1LmlVDt1e5NTwByw5FEd/2Ds6IQZ/7Qq4gFVRWKTn
EHF1fKXAV9dks4hb++IDEg==
`protect END_PROTECTED
