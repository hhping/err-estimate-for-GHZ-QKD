`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VhIgVT2Fyh31aFCwns0wXgO9m+54x8H1ugg8EqMySMGW+F2OmPyYpAhnq65Ce00n
n92vtwOfhBQsX3S/7AVhMxLKBTuEXhYSyMW44FYrMhCdLtQYnuIWFdNmMFUBvzvo
nh1yM1i9mWiZCoL6sU1DZL5oU7IZoxqd87F6vVlF85OvMCqxzQErfwP36eYc5rte
x30iiIpOKwnOLJWws/OcZHYZ1hGsMMnfEg9owAM0M4RMxQwipNk2shi7jCF7dpQp
nuZZ+OpMR54oItM/dalnl+h6QS9ja0gmoCl+2MQmuEPfR+r+eMinixEvf5G9n77t
Rvkr9mjTnn6SBH+8jx9Fl7IY1bPVwPwNe8RGqfmeslEa+GXuYPZwG1WDchfe/KsV
VXGOdgNRDL8USN6qrQSBH24T/BcJJJq7qYTnKDvePD2Nszb5SNeIUeHS38xw1YX5
1njxS7pYhQO/2hZWils82n+lrGcEqUQtyzqojE8L1xV/rKKxqcLVb0wA9WUlSSEA
VNuGVcShCiN+R16hRnakgq++62VVeeKdX1AdUXL+a/rBgTmH0J8LEFgCL24cSLtL
/b/F+N1M6jGQPi8g49SD8V/FGL5sLxoFf99NxjKe0JUVqKHukQ4usYUxTk0HJ13e
LDGsoIQeqtiQ+pLZ/8iiUiDGUpoRYLvxJwbDxV1eAe2JwSWvV55K1j7BJDSLr3Fx
5iJsyv4GD+T1zUJYKhf8Ev7eWGkdrAILwzIrXIFhlozWMll/IBw+MRszZ4ICHWQj
RX6cMfhVXyV7n2Yg8c8eLg==
`protect END_PROTECTED
