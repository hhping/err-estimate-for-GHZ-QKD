`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RE1HfozeyzGD8Au8FQWhcFMRKKwjZxoPV/46QkpolyO+xzHUEpceIsP4NDzxbJuJ
7dsVZ1L+4KGoIqFW31l0o4EltwJsrD68eGcHZGOM6mdqbf4URLlZ8B17lUpE0s3W
hA/JarH6YQ0+ERqLZ66tx1I7whyHtzXrPnJWHkBO9dFr1MboWtpGXNek0dmWBXPW
U1LNRVzwNSq7tVvqZTs9SjhpmIfWGZlhLyeKe6mkbEtqz4yzdxh5DE7Jneo+J/jb
OOgNPccUAej4iVzadYwpk72c7HE29UgYbQ7aJammzj9ccX5Fx9I5/I2KRdB9/8iH
Y9LUC4x0gupRgeRG+j+RrAfBVAOc+JCZOd87yC4zWIDbwbaUP/R62EbB+vQznVDZ
R3cV0hPF6HxdNPFIb1xp+unY4ytTGJS2uj3wGxtLD48QFgtsLtM68VYc96mv35+1
i+GLhmea9WJeS71ujoHhV3qLSeckYqxnyzvXcjJwUcseGzUwEMUflbjQUnwVXZOy
M55FJjWGA6pnQ5wA2sF7dDxQT89SDMNtqFovOP1YGQ6VUwlvc4hfuo3MKSq1DVD9
F1uaHo1rMCU3L4PGFDss550tn5/Y5Ogv2bLaeKE0+Rqkx6tVxyufg2EnLKeMYqWa
sSxY1qVTOnusvHy0fwKG6TEBn5NAWQr+cVyyknC/brTD+2bTKohLE1H84v0pYCh2
8qBhevAqNtRKGRiP+tNmYJT2Jm4FwqFfku/nNZzbiHmZcpV3MPIqNOBPgV9QqobE
idU94rrSAU6QEEfIHSpQScxYN1DVIHSroFcLTPb2uRjxiW563a1vuA/Bhw+uB0Jf
YNU3OheMyeRhY9qBmPG1eNE5avx3z/9cEOVku4GfQU3y5k2SK7Op2fSzOl8R2Nzv
tuR4C44pnqfZW4zLqI0UyhMDQ6HVofz3kDPIDCT5EK4LGvDqtyWpuALhfLIcVFnW
/ZAdoX3EwXeXoCZhdbcsArHGmImTkuwhnnPE++uWcytt3hlpqs8cM7vBBCc48Ruc
qgMHvgPOWDazKulJXHTbJlaM6239WkPhfuyL+TVBaxMJMiYBwa56wpuuST03sFuf
rcnN3/W8CUvG7qSgVV88yi6AVxHBMumDbREsjYdVv8CbvuYmzO8zBE+Ibml2jlp3
mhngNDIF00I9hfSF8LCrU7KmUXPplFbINU2UHw4st9Ct/ym99worKsR+0qgxK9Ua
EaID7Dj3bU3yFXy2KJtwbYZk53zyBu+zhncqbqIuyfdt87QsowQnykMQB6P6a7ju
NtVJMVNdTee6Z2ZUqhHMey8dY6cJEN/puLXWwNUQ1jIhejmPIFLiyMWmuHb0KaT0
wZ7nP+3p0j/SYXVzerX0jRo6BuFTzComtQjQp7xD74tO1JI9pABrjyYpG17gN7fl
JolOYPdeJpRzgdABUqLxyxvEd521MOpoUXgfCafjIIDkW7mBU6VaVgy53GgJ9q6b
g8P2QO4wWFihJQCGmK8Go/RcJooqlwnbAcWrZ45EDc5jRMEIAAHwvjVk/+AWLe93
R9VS8Q4U1Vzyp8dq//xKilyzyB0d7g7rcthKpFDPxXxY1wYHqP+lpQY345yK01Nm
PMP7qJOdrPGnHkoTu/mj//Zgan8YrDPElHAa2u/Tm3Q3i1do46KH2r6hQ9nxxRJk
Ns2CQar/ImTet2s9RxevcsCQrwK/aK0Bsa+XjDujvKxOOPZndrrHFRUw6LKnQAhW
WXHs3dSXbgXQdzipz1Zcym+5dVH1rGeMEhM+Dxq3EtOC3tAmwCRTkDuNubwtZCY9
4JpiRHl5XgFcxwMWg/2Zczslh4LgGEw8rf/GggjlYlpAoLetDQGA3vLW8/NPjITN
t9Z3VwEvJIIhtvMTrmbqPWK4fWKT6wBrkdkvrawN5A9uwiF4/10VAethjPmK2EQN
frcv/HpdKekq8JXMSP6FBA==
`protect END_PROTECTED
