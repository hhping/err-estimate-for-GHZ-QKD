`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VCqWBTzXyhdcx5ZCjkk5gxfdv7m6giDSl54n81w8GzAy1m+eERGbyiN7vQN/ggYY
Pw6GP/epuQPK3ilQePxGyGmW72qMgYRSuNg5QI/yZgheajrqvLqFrT7OCL1+1vAC
Eq6YWBHrrGkCBvBjR0vPEt6FcGAlNipei12zaduiuPO32FRB4VoDGo4F06vHzLSc
ZYvinExa5KF00yUefRokCUgkia/5p0gQYemveHAv8lL1tQ667L9SqSznZ8mnBM33
camegsTNXVABzHdcqtDMnw7UkzxAXn3phkkK7cpbJBAEHpAMMb2HFozEWtk2KIem
9h3YV7BMpJwHCFA9+evLxANfbizVCsBsNo9dWmTf73qhZAMNtHd6tswd7V/sA3io
Gs6TCohmSZUe6PsFcin19Y/yABWGjsnl5Dj2S2GYIfraIDzB4t1We+NDtdesZ0Oj
6SXdv9tiy/SFIIld7OOzml8ZCWgu8xBMvsEzc95kthPsK2e1W2lq6Y3sNuzun4yO
6dzcJX3kWOjXc3EXM9j1BdpbHIOY9Rr9hE6YdpV4pgCg9JN8tt4wl3yhmqisocLE
1XUW9Uf0q2TFWn8hb6kMPfMWsfjGBSh/X7gzM8mImy4R8KBCixNZlUcy6ohMQPy4
1AazpKNZJttYXHQYHUC1gVumLdG0SZ7k6WsSERoaBEYsusEB0WPjPLjoDwKaakqW
0/c0ZnUKiCkT72HJFyS7pSqEjXZELaVyUkLZwQ/pq+5CAsqagZLnVGN8hnoMtxhH
cJsyHS/hDPDQlu6G1YZicAQfw+jgeLVgxX2vl+nX+mlmbHVl4gUCWGVLppqSK5/H
5iy42PW2zWyGBJ0349dZdy7W5/P+ZRW8iKGaDjMW6yphA0+EJ64pcs0gndd5A+mN
3iAT+lMFbdmInsDbk6PymmpkUjFw9TB7anY62/lblgwCcpCYtwFNMQzmnEw70QRe
iYmuRhTae8OPlzuU8ht1mnsVsiRPEmAMk8YgvJ2aZuPcsxzmKK5kqc3cMPhMS8XV
vNityCr4kqz2kU50Wpub1JXYdkoNp+jUffWL7FbrO8TPH4nNZE/919Y4SXuSb/mf
wjpezll5xf7hfbY43sxR+rCddVQ5sFNSUVVYZxPHmkbNfMEOtYistmlnAU2RBxB2
B9sSjb3Rn1UWcXzwLEdmjRjUuS9dizbZk00jmCqIey547xnpkDMqQa4F/k16ImnE
b845UAtfBkOabdAvFKos7CxA2d2oNM2Q0zzpv3c8vWQ0cGy4y5d3alMa03xWbPXD
G3dZbBshbBrygqTakU+TJ1d42z4pNfRWU/92DB8HXxrn/Ls1NcwEdP6HJyJKaM1B
d7pYluysx+tYOBRCMos9C3hB2qQw8xphRg4DXpHN7Hp7XDunOYb4ekYspSF97gg7
+2kYnIqyUFrangJH/7ZyLJ1lfoaaVC6W22kow+T8j4PxzMjwA2PfGt0gPjRm5617
juKZ3gDOxpLAELjiUawcw49+XfPzQpxyqpSPRDIMKeXQo4Op3hNYkVuY4Q0x8JH4
b0DzVH6AldSZEynRlwhTMsqnEbwc8WfGN3DdoLiz+XjL1Z8Th5z777Ps/rZwhGkW
pyRvBEn/rUIbOJXLok6KulOLeii7WGnQQXZ75P4Q2BmCetuC3PLm2hAtKexkbi4F
PGw78C/wLI4AVh2tY6b6+oKnJIQTnAHazcDPzisizTHW0MlFNwuORu92KW0dobRc
u88VjmwzWa29NLRq79ghK6E9ezESALzFLeSPhhRjN5FVtZDVZh24VDXK9WkLvrDY
CSF1QQIrVqyrdTYbOXPJT90Slzq2J7L3mV+H5f4mqIJGZMIwo+K4pRd1G/TKcmMA
9o7lGITGlLN5LuIM/JT+T/gpv9f/mf5+7a7t9ceyHzi9jCFpxLzZFqHp6zN/ZIB0
78ONdhyQzexkn01LnHyj7TyiH+53RdzMzmxXGANQpLEVo9IZR5dqKtsq1OvT1K7Q
PHeRvJpmHCITpJGn7ktybJwH4UEPwLofpASGDr6v926KO+kgS6X6bhQIGo0omecs
DhSx6SIzzVHM6gItKgXh9Xx8b9+/F4IKzAPavSGDZCjz72uwVnOBqwz1xQjEtF+x
4tluR834iUXpxUYpExsEZKAk7HlfDGlhInUINauHoXoVOSv6yh2qPnt+415/52+M
HCyrFEr+gbcf6hSYsokond9ohZNo3UBzP18sZQYEqelps4FUYv4acPSxKKSYpyLH
rcwUW4C71XVIPRQB1SUhq1+x8wtcFxkOscU/UrE1lD8xsV3n9xp1aLNR8JLXGHOM
NfTb6HvThqFsYTwKNmA9eKWvVl+PqzOj1UpVbWNFcKEaBMLxjtH6048CY8bErvIQ
6V0COzL+36AvxYOPHkpIUzr5c6gqBlv2KH891uZZCIsJvpw+8naDvIDBcORTBwFD
GaF9/dtOt9aKWNgbIM3RqFPVa4YlgcCmnKAxrnzOihWtP/FrIuDQHqujoyCjtb6R
6zA1/QoLEFs0D77lCrHATflyhn8ygedRhaMqlLp5HZFGZ61JgjzwFm5ATZt4yyGt
rqTspnSNxBPRoxUAUlyGhm5gBkO357kRhf5e7yno9M8FLwjpBm45nmzNrBBDkIu5
aQ06+fqcX8hPM0i9p8bfCl7+ZGFn2RZ+732QdtUleCJP0iqtjcj1SGqUUYEY9xdN
G0JFvBViSLViE0rFIXV44L4H1XrMeWIICpskXLCzzqYN5DseZryUTX87X7KdcOnb
OiuBPv7Lqhciftlf8ECmHKUmQiAXfZawEiKPsy/fCbt68yKE93o7nDVRVw47Y+mP
3gBpYfgS1oxJ3w2YHLmjCMRVNtyTAyyuCzajv4E032y8VThvPXE4u0zCKa5e0iVF
CManeRSc42hRzLZfgQaIyvGiAWdkuBUtG/4Dj7FvUu+Um5/4kI2E4U5XzBGYhPKw
ciCZO8Y7R7M+c/bMtHVuVYl5pIO3aJDSvMbRIgFoDbVzH0767Bu5xO/d/IcsHx48
KJhrRY3OGmui97qWxuBHyWc5LhmjahBe9LS1GIeWJ8hbfHmsBdLP41yaTSolknsz
qVSKsgUn6e78S6O5UuENXUkO8MrpSBd5gcDbWJD1zk/+eGKDCDQa6dGD9/otMPx5
0wdoXLZGwChtFbI2SrnT9dzstvxfbWjZFaN0D2rFLp3pZzZUUFr7t8b0Gfg9rIO6
nfJh/fI0B396sq8yZuB52MQ6GchyAc4y4svVpid5gwHdQhOjhGhaM0jpUsjF1biG
oCzIOUVT4DQsCad+qctcxFAAbb66WdjxqugkEACK6VQ2Ox2Ckhhc7Yf1xT1Qpr34
x5/GaOGxkVF1smzv5mJBhXdN1Mz4Z08hRxy0Cc65/9yogXRlyPTZaw3nREXfV0XX
XfxjYINMNv7dXmvbqkq5M0mBePuMcV9et/ZXLcDudqOG12lwZ0hgRPlVXX0gczzS
Ixr6nZPX4ipKbFSZ9oojJMQ7I7MtvGRrEGWEx6VYc9TWaUG/FZH286HVxHYVu1rM
PRrPTuyj1qJ+RNHdS5iwERHsRbvWx8RVYNqhmsG2Xn9WL7uA7WwDzFMbA+hIcB0B
IdLLuvZVg3F0nRAjtkK4tru2SvzAJQhC/Ub20Ah7DZdi2TBJaDmuGjtNhWyyVBIf
c8x3TlFyCfm/9cnzDswZ2+F01XY3PR2R1dl7SXJnmYmJ/ZjmyhUNwdZn5zEy7DxD
3ireeMjWiXJZPHLlbyNwNr/ApMOw7fARChWic1t/RKIL8dfTwoczlnHOhE1d230k
5DDH/l96pIPHifJ9hZ87iFx4rOUzlPkB8d9u9cCK9bCib4JTtD4gxisFCjkVGFiC
RWZbFWC/tqMTwMnNqYziUXulEjvvwGUajV01YOAR3Zk+q7Q7+3miGvqpjwfakUcH
Tb6ao2pU9cV003qxqesz+Tdxs7wHAtr5KmFgtXqpp0/r0owvr9Zl1TqFhKS9rmki
Z9gzM6uka9nC/TXm9VNClbQBylfvAgk4LILSMapo52YiF5oepeLcj99RF7WlGxhK
JLmBi2HnLAfq/ncyny1/jKbl1RV6w4+t7x94bKqot0NfeEVGmUV4IxODzU4WlZuL
InfHL22AD/WNeFCbREHQrrIvQykNqcQzzpVsVbdE0w/jSuDY412B6vdGE41obnqI
P2P+v/T/zPq30qCrqizOuyFgrrKANLF3IJN9nmsvQZN+SAiamIZBPIB+k+9EebaD
Amq0JnjNnodTXixR/e/0Dn0toZAlarbus/X7Oi/0mA1irPZCE4Q5QRBrQdhQsFLr
Qb6jN2tZ9Gwu6ztq1LIQ0uUijTO7ldeEUVaHMDp2y6ZZS9chGcolBwMWdxYh+FEN
EWav1S/GOcSfv6OiNgC4NFADi4Q+7a+LCsIEe5GMnYt3BJ9G1Nqb06RgIqFQi6Dt
bUtawc4jWKWFePKeY5FdW9pP+h/gxv6ssIhQ4/z8YlY1sNHC5Iala6JekYMTBXqz
jP0PjEyQv8BVrD696eSCI1PHz2mkSLGrRtQUizq5/ceodd8kQk+6wWdi/Z09IT2L
YVy8RQ11N9oaOecJz4OFassmwr8m+BjEfxcqILOwnJnYn4igsjb1SdQvXrncaQWJ
8OG8xZbrNxJwPgzMugGsGjzOOa2hjVC4hNhelazK06Di54eT8DlpIltNbY2/6+K8
laI8pkiMzmNQqWEVEZ84F7kOsK0NSspzcc1JzC7AAGBED4VrJwdJuY+439OloXok
coDglKewkxijqz9ltyPgXCnA/wUdVESNsiqx+ar+fMzwiBfNRzb+/RW/nxPqXk9A
jwcdf9y+FmQZRdoIYPxzBuWgV32AAvEKqbPQMGb7oHunjWP5uNDEW2whA6zf6NUw
ZRnzH6ifNTL86Y/zu7T6uqsQiS39uj3TF5z+Z1FJYA3QZLkdDd6/2apc6WdnZv5Y
fN+zGig3LIrcdv/NHqn6Bpt/Z22pDrDFitjwyGGxOurDiY0XOBwopCakEv31BsjB
Hs9SLz2XpFAfpzPd4/HjF83VARkojG9209uW0uT9dPVI0UwjXP5ZYHMuN6ekG5IQ
mqrIKMDQRD9NShfC2Vy0yE6TB20b88QehApZU++cVVZMmaJF0yAXKHzz25wrwPBH
giFmYTjvyUNqEm8L1h+Hf78N24bwWxwKYrodlkaQVqTYqLR5U9MnbQW2TD52U1Yl
irx5jSV9ZFSj5j7PfS8pHdjQ7oxmi8d3aBngDnB3D+n1BrBnhl8hWVzdEA8zaRG9
CSzGM6PBYPijVf7cbIv4+RRT2WCIrOML2OzxEcwPO2A9CiPHl4SvWfzXyovp3Xpl
NhRFOt3qwyUJSNrDo6lyjHhkvPXhOreNXDJbM8SyQWXbIXHNrDxLMEuGMJIFhQCF
/C3mPmZwAemZ4YIEGSsjoIQTMXRT+yT1NZqebQS/Hx7d3IQINlk9jolvSPto9p7i
Qq0u0qq2NCa5NhTGuUEtIM4+0sJNJaawLjaSJRS9wtiI/ZKX9xitJT+es6IOK2lZ
o86qhKs6wc2otUz7QzVLxBv9JUXKhYt7Iu47213qfWtcIjjWHXE2iKLgfgPnBIAi
0VLe9al634VPdbcU787RXTNqNJawRP1D5GNNXU4SMJ9LVCyDCe7Yua/vfL9v3g+7
sMeJpebuGQUi6+UVB4JrfIfsHRDHvN67s4QH+UJH6wGIsIi+VnGg8CeYHb11VvaY
EOzIC0ni+VRNcUhR5/EbJ0YfNfBSfMB8dYOU3nMgkryfF2KW6DuEldvb5+F50oJ7
tldfaY0K7nnxo0P/Cb4Pu52H/3ZvEUqEEMPGlEG8ANuZKmDvuLZm8G1edEe7fhd+
sv0k8NU+6JHVk0+eZnxmBQEeMXTRNSPqzxlIWSRLJAiIhEODnTFRdvpQZ0T/9I68
oytT9nGYLxthBPA7byH6icl5TgExmeMG1sJ+93CcZQEEE7ZxZugRNxCnmmGpNgKS
68/vMkbiZ8pMZnbLBpeXq8+wzmWiWKiZyXybJDRPOea7G358qP4ERAT9+hiXEes7
OtLl3KYhTHJI+rbdC/QBoNDSLnIfo2th2Na5LDPdYE1WjssMuDSo/ibTS+hJ+BHW
jr9TH/4rUzD7Iu3u4UbC6PXbSk16qpfb0VaXC877HKbRYRJCOcKqCrCFxuqZDBsl
FgSoV/48lG/26WVPajNX/U5ANjR+KBBmzhLij5av7l0BvMl1uMFPhvLw2P0djp97
GkdJd2/Yh6409VwWjYxnp1FDtEmS3kgZNMZHpMJDY/0i7LDBnmMBOJ4RtaxyIKWq
oiGNZn0tnO0lOKdrbEtDN2u++B4xq2DThR0n+Pusc3YqdraI3qu/XJo9jk4gyoaR
e2XrS+EJY4Ak+rs0GnujEmzdDnMVxMJ1qLBfBDQ2dgHE/RvDF2zuOMojXWn3NX6O
l2p3IZQsr5mC15WoF+/5lbbB5QtmhkFTkfRVcIPTjkKSXr7P4yel1xd4GB219sR8
d7N7MRnduTjWXLGKRESkYYjwlgMJF1CkL9bmATr2k8uhD/e/6nB6dLoT3ucAEKvJ
4dhVl7lX1czwttKE0aVJrSPUrN9O6Gllspiws7PofX3zm7iPm/CHL/0SU7SI79nt
Pi3XM1hdLqkguZcb21wDwzkkybVh7lXSmSwAVbiYahbLYv5SYaBXx5V+dreYZdip
aPYBe49FHFfU7YCFb4yE/rKIEYMdlhUUpTmSTsY2gJgjKnZxSq+WmzKOkohWNuJy
awfavFFi5FNcjFf7T+uoZewaJgcqUjYj20chV/mFgpF8+qCHQWdDw4s9cn6qkf3+
La0hdD22c3Dz+BCnrQHTUxd4mZUnZBsRYRZJd5s0r7K3XzJ7ZHwTMB6K4cAKiej9
D4vzIVliD67OkpBIFLXS/chYLjnFVB+Asj0fgP5Nrk0NBf+B52JOyLAdsbD87CRJ
pvTjjC8s6ci6PVoaC9PDa+Wry3DZXg2kWFJGtdLmpnGKtJ9Tx7k6jk2YumQ/gBjl
agEW8iovKENRhz2EwJ1SajEgHaMxpQaihYwgEPUxEKFmWwlCmlZa/vXWpEYUWWwv
KpGQ6lbmeKUEKz0epm93/6Ma/7IyoKub4sGNR6CFpn5BlbuZGAdGlXl8VC24Nujq
9i6g5oATMemtuHXpYX8wz2lzZwvXKGu5pANCH/wcdStHBw+D1PVCBAc4GrSjG+Ms
IL1Z8U2Kb1HAfmiaLUXB985grQda95zAOv+57vh/ECVmMIcXEYBA6hVF5s8S+S3B
9+dQ3tgyluTGD/X3qoIm0L0CTffphxLTWl/k/20ptbclvdlBTpGV6EnZbc3cuNLL
GBofCIzkKFv62Dgjg3LU/QehMcxC7GptAQV9RqkGLC85XxLGHuyV57G+RvounJzP
pChDP3erCO8a0guH8c2FXvCTfhpHlfMMOOMD0tVpAEC4Ubck6AuIOMohFLQBpjgC
21Fsw/4WdjDki8r+DQ6wfdgRIpcTBVTqqAxbFrqOfUbvRhDF/3dXepB15d6fE+y8
mT5RCRVGJmY76KY0n4WHLT3nvwxyta1EkIUTXzhDQqyOSTp6Jk6V1RiEHBQbnnq1
pd+/HODqVJ18495to47rOAB6bPYkAsbmVvY/uAdPrEV8Lla02VVrc3bVR8Ww6OJe
jrbrwL4wjxWENFEYtAWtUbmsWiK8agbEy9C9hX5fi0xCDUZqxhVM07nQ6wNb/cRG
e8B1LIkJqAKTqyk9DM9j32ZPyiZY8f1/Lv4GZh/hLRBk/NokO0Kh/p9jcDD70z8D
Pe9Om9Pp2rWjEuuSoT5NDtXmaoQVeFJKBtyA146vH4NkBC4CTviTh0M9EIqjDDnK
cF2mXez8VbCaatcPAL6gu+cXu7iP4nke6TUFYgnBiIANoQtpUmJ3JEb83C4x9ix2
ZFkr+67gQMCUKLYQKuRjempuGrF/4FtW3KAWc3rNVPGZPJpfSx+mQ1/KalPQqca4
2+cKZDEpWh3JCVi6rRvNx5TnLeLfYIWrZ7YLaxBTkZlFulu+cOAQMSciOCPtDPru
6vlFV/CsBhQ3CSTfpvKUT9C2ZJ9Fph1R3OO1hHJT5gmAfrBklWPXaSEkg5uffJhQ
oQNf//NT+m3PYiU986dBFqWwVnxDKM1nr1h0iEQyXbarZwk1zYdGosgREEPvfpiK
7VbUfY0w2EV3HHzahWjhzGnIiHOfU5A3UWmAXOWMZiIcAUswM/bXtG/EDM1Xxsji
vjC9MDiuc9RYos61KBoG8vvXruq1yXJiuTCWSiax983eEyNW7Kipm6qGa8MVKX6L
58vr4eQPvnpsPxUhDdZqqmOD2IVhTmCFO7NRcbnfi1ktOdSU6ISRoyLfnQwoCL6N
35869voRGLi4IPW/xbOaqWn9no43vaZxvUpYOq3lZDD/jJeicq97dA1fE9AETh9W
bV90Q60aCtqUTUpg4UzhkKfVU+hVYpifNF7/uA6eGKfBOT6LOuIFeC4EM/DIuITW
MPW+4OkVgGz7+9VN+JJiTrt2Y1cLlD2/yHLxWOr4u+qWp1qKhEz1407fdRI/licn
K3+tbmYhETn6v8MApTAomLGFBAjNinsjZzVk+zvY/7tgnqkXsLkD9n7z4Oy7jzy8
zYxiuFEWeUn0JVya1LkQN90zh1xoIyWr33X+Hijp//HCH2nm4xG+0uK0V1xFHmKA
JvRbN3s+uE7OH3pivq2fnxOBVWOVAIHxcoi+9t7qBdGLzQLBBSw5hSSACoX4THp9
Ldmk2MwT0dIs8gyEr2tdcPRSYjDSygwMPlxpYA3b8qllJWNIVplrWo6hqS/2h4MY
ju0+NO3pJ7zbsIA6/fQH50dzDuhOZlDoss40QUviL7E3KW8vGiKjZgfyQCd2QLTd
CXeCpWifLMWZkY2A25JwPOuOm1naZqbkb9Qis5RUUyNplsPC1oADmQ3kP4RfsQdI
e2mphrzOX+Z8I/TCxxwC20Og+oiyxePA0SKXk2eZhVHetmqkK01EO+PyhSJYbcp9
63T84qsWGlw4pdRG7Ncxc83uEjo+E1LKtRlJ2BbKbrogWbtyiUxECqjOb+lahOo0
iRP5CRyGOZ4bMn/wro+vRa4gWaKrC1vSAJmn3E7oj1o7/gNCYBcX3kOqRof993Yy
Z8mhmnwEbDp/FVp/gCTI8+Vg9+oRIFwGr1DCX2TkF0fgvL4P0znsaRZZMjk1hXed
nA2LrDDJ8AKqh8ofzsMj98uL/tx2hqEKWWs8UkSntqU1gKq0HkTH8jI0ptBijW9w
iS61jBhnst+KL/zSuYcw05j1tGGzQ5qDhKGHUP9RJgfnOXODDF63irhmFGA3s3hY
uKa3be4nY0nL2yfAHUCJ73LwyzLssvPcjko8V4rdRtFwtfHUpFCSklRNRKKRQ1DQ
hjcssTSnEhhfIyANn9J68yzuFG7H5ovu02ZRpncbITGYxY+UR7DpfyBZM04rY4jk
BYazZDGU4AGqi2BKJJsmARpGMrwnXPPR5dhS5lrGr9KTQaN1IB5r+BUDZ8Xm5T5b
b8wWUy4vVjrwcJzbiK6WYlLib+RyAQUC0BqclJnpbv3/UuZ455XdSj10U+CZRvDI
cdrriN+QN4fB+svx1+dDRqG1IKKnFBsKeTaDu1dNWFqHjvRPjRR8JxHfDCr/GDao
/lqa1ccNsvNwgxF499/oIg0ITMd//Is+gUzHNJQ1NtcngzyACdQE7QXdYctYa77U
XmQcRsxgF93oKNOnRyZsIRkWb63Qf4rIsnb0JrmWHi5CtAHhmJyb4GyFUmB4ywIi
0Lq65rtGDoaASO4gJ97+Ju0nEeD/fiBMZxsg7N0P5ybyE78pbZFakeeLxxQWz2vO
LVn0zcJ7qqleT4mO2YIYn0MdHES2By6JmHpNRAJzG6O2lpR4tRcEvIRGhW41ugth
lzMwp2eAy82fa1PQGfaRz7U6C6nCEzPka6VElp/iP/mtTIcN5JtUdhG1eS4R7QS8
tZFkDbV/7bcUWOGEwqENqGB2rkZ3FjY6KoV8gRQjEpsSDGXrhc/HeMkiQQUP190z
N7Jmd61ovthRgnEWWUriGm+oU/HuI87Kub6Z7uPhrdLRmDGZsEoZrjlcgvFg6YSk
bTzq+6oizh41blEdtRzlY99+EVIyBfhC0ivCVUiqrq4OrnDngTJ7eo/heW5hcI5R
BOxyb72pIE6bb9o4OJfeHsRieYEtSpOjAdvAmVrlDemcJ8i2Yb+gOwFky5SQ03gN
WJn7/MyMRgkA6Zqz5T6XhQ8ULsXckthLRPl/djNwian/w2586fbqpSZBJk9/Jw/6
oeoRa+WXWWOpjGLge8qczdE2xIU0iBn53E3eY82wtqG5sTWV6Ul+phVT8RYkZ599
FM/aYWokE2GOte6TIsy1fZW/E7m8dl/B9zphDigatV2cDrgtZ7FVyckKLACvqL0g
dJv1QtHvkVy7Nx1Nvbst9+sunMYWWUk1wpPilWrnCNoHDorTl6kwuzixZ6EnXwWi
eK9INt4cSwtifRXyIpW+9jI5piaR9b4yaiIu6e90nK9uV1E4LzuFDFRdejMJoDGy
0+plWduS2mTxxrkxEX+jC9uxapfX3SIfIiN9ygocpUM6JdADxCko46JwE62wzWku
MmNFHJK0QKMASwg6NGv0ZxF2FDyJR/8tMvpHJrW3UkQmB+CFp3d4sTKQyb57TQB+
2CLhzkzkSecoppx2GYGl7PqSdmGJ0WB7ZGlBbu3JNQegXhoyYKL/v5JbcSTCyGku
M4hUUpiXgUnDB/7F5j7Os471+qBz7gK761Ujsl2h40mXyD6bzQXfdr5ngHE8SGn2
+tAAuD5HXC4+u9ss2TrIVnOjSmGbCJDbPIWlBE3WLo/NG+2XapbzflD29LBQWyE0
r+fzupkgkWsDBonLj3Y6r38d/WZ6knnehd0JMsQXte3r7z8xKDnSuzZuxxAELh3y
B/Qm1IFJmDB494cHbc0HZ2iWS/weNnX4KxDT0WAt78x1BPHofNXtTsgcZBojVvlC
mcIHff2JAL3xjAZi4qbPlxpp7lquU2zactd+D6ZIKgPiyQ7zLbEnr2QM3x9YcfB6
8JiS58E0lqnhbXzOX5G2zFKrg0nYM1yQuiRHTkBUrg0RqtcjejiictITWQunV5YS
IQNXj7N4UqLbiCFx93o5z1yCDrD1rxvGbgb23LrdqPWSxTKBalvQbuqixcn5tu3L
QqQA+BibMlfbVCyTHVrwiG7aKnxkD7zzVtkQ3vLR2WKuaFAHOJzGFe6WS954PUsD
lPD1hXzCMN+/DZgXOSg6VMzW/IpvHMprZ3JFnmbZlvyJZGVKUkfP+183c/DZM8Du
P+dnBBwPC+/YE3VAPG25HIvQiC7kOYiGbTw2qlZrhYlzEXcR7Dop6jjfTH+XYgdP
0QUzziLZP8s7VrpXBqO/fKWwJR6xR//Z5r44o3hJFCeugyh0+FM50RWWxzuyJ4b7
6iK4lavOPlq4SSCk9gyE4MMN8fC1/RLd+NCy9VltaqLEU/5i+0BgWJt9GVlIRCkG
R1zQlAkmZRmaBqa+b66idS2iXlrBqo6XJhGmiSIEUFt95shvN7CO5ItS/ym6cOYh
pU1WP5QAe2OXF2FAVF6k3XDdS5ujhbj6q37o1JbqbTiNsXrhp0LGmB2IG1AZdGn3
fQE4BW0Vt+vEHU9R0QhYh3GaTnK3u1fYb0RAXOc1K+TRvI3ssEWfXGnwy2E6aGB1
h1LsfPCrG8k6GzmYqA4Vq6w7VXSeNPK8KGPRaoVKMmYeJ18BImlCe7UdpuZRVdyF
mVTJTYEWkLdq725xl9s9A9wbkXf9HpTU/93Q9pmarKkOzRFu2HaBFFv2yr6bDzI0
5cU3cu9oGROjm3LADonPhChvP8998miqnmhiENeJKfS+cxVYjnUUeqDpJMnSyuJk
DeDqp7ahPG3cRAVO4Ir+3Fm5upZcfYY5oICDS049ZMFbSCYThppKshGyQrZJ9zvl
iPgPal4VnDNweg2qFzPaPkiXS126lBi/UHRazTeWPkccabwTrJ8H8YSBLJuTax4N
xr9bohN1vFkrbSNXz3cUWDQVjthtKsxTohWWGxZc/8ky56bAwfuD8hOF8iBIt07z
cq0QPo6UeqGgw3unjatIL8VgJLUhFUwafz9LL+lnrrfp1KdFm8wk9bLgKAnDExmG
nOvS4y94p2t1LcP5IUgHxWdd8Clz8z8mbaefvQKEyw9yMShu8JUAT7jQ6l9oosBW
aAPMsJM9FPzM/Js5XEdIowcfu0R9/pPTr2btOm5w31QtSHdiB0PpwL74SlzP3EAU
JkGs+vR8RXEpS1NWaRPLgP7TbA6gq/RmbKjcT/ZqADK8MoCJyRuX6Ja8JW53GH+T
1h3JBw0cNaYK1vpfcNxBcoLHERozpbXzwJKDfkLpVv1F5B2IkdZ9lzH8JsD6UK+c
cUmjFa+Pw5mKg2JRjoGllbHe3pbDz+v9vn7P31CZrOq19Hd4Zq5VifGGjBhsthSc
339cdrbUueGVDZZ9VWTVKt0aS1sUpMTYAqLmLLe5U8DpVdFi2WpSdENWEUAVzZWi
dMv1JkWKiVg4vGqCXCVhZTeU26RG1d/Hy9UkzFcYJQcpJWj1B6sqcdvMjHtJ89CY
HpTt/s1nOMvXppTLP0/7M53B9nTRjsxfqSq7u9FlMIs3qvC7v8+r8m3CM9zapVbW
JkmTwFfviTonoURhhXUg9uQSmj/wNhXcjLax6Dy8gTq7B+cpxR0Z2jACTaGrHsqz
WVHHX+8GFHtmOTc5MV4hjihGqsdg/pQd6rY6aXduyigOGkmQpfrGd3IW1jGmUwvs
zrk/QUg4jTXSRP01fOw+x8Mg7SqAOYtwQxsjM0KK1DsDSMoXtE+b+JtabemhNo1A
BWTlKHlbe22Obw0EjSTA0rmgXfUHJ9OSIwjxhsamRjlIs2AFuHdyTag5mH7KLoTr
giIMOi7SR780U9H4g1MNrU/whgbDTxcsw/BMQW/GJwlwFAyXHviJAidvAQgEqYrc
06zOp4AM4ubi9gjXjCpdhV5NE84WcVY/o/l+WqMmqNWAyxoau15strQAV0NHcbjO
MRg48YOSkaz3MmBUQ6DvFoD760O5R1O+/s+JXjxakYYYO2ef9/WFT5DXA2f0mbAr
rF0KRvBWkY8zLqM4278M9qzxaHkhovAJGcGq2vdjdWu2G03KQ+LaQcm4kDrl3m6b
ezHoqQHoZ95j9iqxn1uk8ljTOiX8hrYOxOhF5jDiflXtAaHMUFrFMXOf17/bq+ZF
+wqfuQc3TOKsVLzDCAYrZ9nySKbCigYbm3msrwWeN60hnbFQeBQvesobVkrVqS9B
WT0jryTW5WgYDWXURsmvwDlwdPQLkzVA7l62oG0iNpBH5s4l/c02wldZuyyJUJGp
61Z00qkYf/iFEBsTO6TR9+LTf4rRzsR10e7x6LfKesPujRHAo2RP57o9V9qwbZ9q
HjvEstHzKFGudvG9hKoZxGhZuVlkFfdkH+/ddRjo3eqpkcBw5fmezC4t+W7X1YtS
8VMhT6LMTlFL2dQqsu42rivvccZ2djDf/e/JYaKGiyyBCUX9tSO7tmnsG9+wvDFQ
aa/r+TAZ1tcu9JKsBNJRpzSmNWK/w6Pt3lgXrNXU+okLEqf7wcH4EMCT61y2rZjl
LSPkona4N3DinhAUlHrrX+sEljvXELPb/AQWywAB763B9cBupI/oqYKuqJ3bVkam
xMv+jhMN/D24OhkxzOuA86LaA54A0m2kV4oIW/ZpH1ISzsknQq7Akigjk+7ZYmu3
o3zrFvhqKqg066priyfYXscayoYOHFxE3nubaWZiDgCgXCOsarsqYEEdlpYvijUp
0QmQFait7SS4Wbyqa3+/FRoEphufXDblFGVm/AWnuGhPbJ9KAkRJmOvTMAhLR2Ob
ULA572BVtUxM/DCoEY4CKuSkqfnU4VnbPN/4+Uq5zBY9QmVstt72sKiynuNv6MlG
UifoK+NeO/J0vQCn3trN5ZBXqbKNWd8RUaV4r+FkF2UdsyCNleDqzZ0C2wSX5bEc
FIRItXRNs3ukkS9st2zepxZZRsTPuKgER8lj2LYxJbOREGgbLiAwteswDkTG3ZQO
/WPyktY+0Grl7xZeFInndZnzhEP4AxvzGA2kI2etnHp3rd7ZIq9agQQ+rNpT/hWb
A1diB0+2QjI+mQ5pH/1uNObkFZ8bU8oWusFwasLH0Awpy9yBuOWVi59xCndfEa1p
oIET0dq5QVQbKD4/BRXujleCEvcVOqg6gTZqEcg2LZPtZJhhRCyyG+1e8vIOKX61
JvxSpH2DNzgNrEnU+rfOwDxM3zLAflwvbuNhffXLLQAUjpYJVPIezHaQCBU125pZ
HC1BI0spQ5Wen8nVSU644LxfFTriUuCB56nOH1inJTztHgMXRz32tZaQC3Tv2SLi
Rgmfm8Eb6OY1kx44gN6l3nVSV4y+e2miguCOe3wC7mZWutE9thYw90gE7BJl2B2c
wEJF6Hf52KyWjSSZ/Xk0xCvQQ1b5ekoT2piR8SB3xJHQN14a4a7ZaLWaeo2X3JoB
i07VOWhhq1dMWDb4TO8IDnuZUxY1XZe2/1g82232yXOJ0V1082NrhTJHG/HWJq1N
pfU75Eecy0wGmM3shTQWHGeQMDmNgpE1nKIiEO7IJcKUG29HfX2xyAornry49w6/
gYY0skPYq+HEQvRuYRFEE+SWaPZrZtqogpWsrXwHsEjKrWKfTBO5NUv5FcJ01/vg
et/rRcfY/jwY5WqS9lif8EdNd2aiZk0YjVzw0cHJqyTd8XCNcN+Ft8wisGvwPStG
/hXaUIqSeA5/cNhEL+m0kZnLLibq3zeIpLOx8vkgS5eaoRxYuVjnTPR7qpHRTNWr
0IUkwmtHR0SgUT1fqo1guDWzwr13nX9XPq7NB2FQmtZVRrnpAm3j4CMFAYbIvJ1U
O2sXWvDelvQT4zQ/vzNOjSZJu4lPXv+E7Mm19Muu1HE6FImTOniEuGqffgrN5Ctb
dS3AtTzFtj5bBCNyAelk1d296d+nuOL0EGrbxJcPK/qjPQJmVn08BXXR4HWSWgu1
RlGKPDirkrSjVtG/7VHj87pUyxnaZuTTBXubNqquRJPl7mnYCk0fFOE+clXDUcFp
loT1xrJwdWwkptxuxXrdAHwFDQjMclOhIdTMMgG104agJglfpyNxveym6FcaKi8Y
EQhjHZm7owhoyxEWs05s8MAYgNQ9+AHauw3agzojbekiu81FhTYRJgoWsX1n+KT8
vklhv8f5cT84OkdJd6B9KvNwL8Y4br033D7y98V8KeGjSxAwLf9LvVRqqLGeJ2oc
TqMZruL/9koNHcaa0J0OFcvpmITksZEvgpe3tmTQKUFa/8l8G8T6aqdC8FyGndV5
bPQyHxqaHEH5cgpMZPsb/PH8Epj4a1Z6ujk94S691psNdF63uDqiQwHV+dC2YJjq
tp+eDeFM72Ibn/hOf9+9PfKUJ0BDNEi1o5hvQ8z6cu0wgL+9vHG0UXV68M/1e9Z6
f+SeD7mkkRM4kZx0f1wbcHL7XehEg5cigrUhE37dQa0Qq3oWAxgvtU4fUMSFgrxJ
xPdZFa8uD4ccfMli5iIcgL7xtFqZ1UlTWA0z1uy9vNiaXP6iDkiVolC3ilVxELk3
PkkKfA9VqDBt1vstJwYCThTfbp7ErJhjXpbzQViUOESVufmP8+2QW2/FvNuFYLns
GtHSzOTM0o9nB6KZUvBX36AUWoWJQZsP5qcxs5EMq7FMYGzHZRW5g7GeQoCoQY+e
RAQsUZYwZmUgoQKODprWAANZ1Ih4vdoXFcsY5R4g7Xp5nVnz0lvwd57Xa0SYJPIW
ziR1U52WhsaFyyRl+bxojukZS9WLQlrCRKAna2iYVk7FS4CezwE/lPhnH0ir+HeW
nuwwbBGL8JQwzsUW4l02DOs3IDGF2BrV8sZoqZJtrDL630PJSq22dY0rP2PAQDyB
3gSD2h3BGnHwjDetwhumAuZEiDZFH87W0pIR+++sZLg/df29tg/pcKanbMUHHMWU
wzgdYKBVAJVuD6HJ4aVfQgJaVoHHVHs83835vyktTd4306pU9AOl0z4uONeIS32S
n3WdwA/yNv5hfWjJ3rCzMGDDoXBPRFjvVM1jA/s0VBNF//HoaMm/rrbvnLx+Wf7W
SoZU58EeSrOEzAgrqMTnejlKmjlnZg0DFy/noiTECD4cH21jam8nhiiY5EWOay4s
+h/h2pEefqvgzqO3VdUDX4mJ1mWW29sp4QmTQWXCBfmuvuN5pcZHzcE1h1QQVISA
3rzn2zppxQvUXL4LevrXu/EtrtkRy/KTiNAWRBSYMnzX+ldKhLaNCy3UorkCleff
U0PzbnA6SE9eMe5HN4y65F7M1j15hvd4e6Obcz0KjIvZzY6A/o0MUAKbH0IWhqBm
+c8OJHoZ7kilL6XV3rDIFWSxbXE9MMQqIeBRhoI/3LhVtMv3m78SNp0g3CMu1Jm6
vRr2Ey2xWCHPChob+svaQVBoB+APEnCb3BxY4776c4qGTLrp0JHIJruDpvYMj+5M
ved+WWx8NXSCkvsVu5m+OrsEWqs5bB5xqQYmoUhmcopFIbvWbaITT8QVLCoZ0fUS
Y5ZFzNI/zoURoZK78Oxjs2p/O6y9+/Lq5+4pErzOwQoM0rkYrnFLGjMvq88ern5t
xsN1L9ppxxdFZz/KoKC8Ye7rPSj/QZh0YrtbnuIvvPxWcmUq1mcoYLe2qYQ0RxYs
BuqDLFNSE6+OyPgD5elo4XUzw3Z4EgnPSg1UdGMCAQTzC6AIk9kP+BivZmryN46t
5g0ihDltxBnz26G5Xto73N2+xyNjB6NG+m9Iig46a6YrHXeBryJFLZIP8GVUOuGc
LdMblWEFbvaizLtha7vKRYPRcxoYIoQgEp94mqcbn2EvkDRzIWdgdbSdPQYBm08j
3iP7pFlTNgatUlZ1hmzQbIHgTXnwiWZuU1fjxxlq8sDYsc99LFWaGYtwSbUhCKwb
jKt8v2XhWoNlGpluWBsnSRo3iVSQqO7ENDwbokPjfYdSgWCu82in8Ysc6gCwmP6V
lzSIbdxb3H+ubTdMznSPtl3a72rRQnNiX15E38Y9uLnrKgiJOmiG6d/vhsmYDlI5
yry70vqVHhxCmD3XK2gBEnTZfC50z+iUDY/zRqkB00EEy8++9amx7EYx2qulSPLV
8yaOx5wVW1/HCMYWxY3i4E9oDBv6NAHTGEHznCsbtQDc6CttTSH2s+ouvkDJXbBH
pE0QFXMWPBMf5B198kR2jSDmdODHznsbd9oRvz8ihpB7FLmEgc+d0fFayN2bdn2x
+jyE602EGEJtAShqvKWKFBElZusiwxo1r2JBThpAMA3Z7oplYBrFj1XWa7WjnNpk
vl3ny8FFtOhAMkTGhofDStHnmJlrnh2CWTJkpXjUTZghsNkWvMLsNgcbNPntpwrn
b4AWQq0T21tPJWTgBSL1MjHMwa8m7OdYwZShGYv8u3iWCtl5f3CIKjTr4OBOX559
iRTuGpBtnNfDyMQTdt4Or42q2BNGeps23yrkyGKHE/XnUg8yP2qiMhxpALmneBGn
QoqGCMtGJAJP8GG60XzK0XJfCFwr74XxUCMvSPs9yBIlAZKlBaCW7g3o6WKUKdH6
B5Wd7+IIMwzb6gW3yeJ4uvngsOrrX7o5NejV4P/V8IrDUC/VOYYNiC9STTe/kNc5
z5Okl0A73B3+v5OMpjElqwPIuQrNYYYRNvEV2GVUUWjg0Zx47LojBlvZtBtGbnub
7Lkw9PcWt4B4uvRlDtUyK6znHCrBPmI1buiZgNr+zOXNe6TNOcBCsB4LGhJwVEBg
ZLdzq8Q9bpyltPS9X8FfQTC9tEC7eP/7s+WJifpBpSWMZQmM7uU3N28SoPVslZTJ
4T36E5/LGC5/5/cUc6lPKYJnX6Gm7Aw3jt19TYYJkiufu1JwlKGr2trurC0bqRG+
GpsnOzssweKjxAHChGa4+8jQGJrAzlDYmCshgDrAvOA6Y+i0aehovkdVAIZ7O8ol
p7azuiMeXpIiVbEP1f2jEXU5uFz6T7FyLJUFlEEV3cPBwDvnwaTa92JlmrcnVUdI
7ISCocZrSRnWNFHAOIH4UP0pbT09urMoY7MQrc4fD9zqbmhobBOYNE+my1EIzjUY
uvEhdmPdTMw/XtraP6wcefVrSaHlWTkvwKsrFFjwdbY48hEe/oG/BVRVc/x/eVK1
cFZsZLAsFtQYi5Lxr5bmTHUrufwLBKLXa7jNLqzOGkkCT65bo2jLfZ2N0GkycDlS
3qRQV9uU39KMgLycOUDjBclV1HaFEbXzeuMgeZ2yX4eVgtJqT7gVWyJjjb38nXti
BD4I8QbgOTxIerayqNwmuo1lJzOpgu4aPjCOGyGrJzsCUwCNDa6B5OAO+5+xOhDh
JfTEO2TjsHslntXgknkFkBF9HmsysHXPcBgczBMK4zkh5SOWkX5xToECq5QlTxn4
rhwOR05GQtpiT3Yg95EaItQexfOGAMIeOKOvroZoD6xib+N/+tIZRv/F/InUXw3W
BfLHC+6vomiyQtVoYBvgmPhx5JQTPUEuGdQlLY8LkR4Bh9egYSEGsAso50WwL221
dnixV2nZPhZPdsgpO9jVZa9all+fFfaqMZ7m4trtAplV7g/WQFB/dU7kHKoBEANm
5osDAP0HEnmbTQk6T6qeN4MTBoElIKvV7iw8Zd8HCrH+kS3s0KgoGX2ZPJyLQRX3
Zin/SYMyPQuTKASIp7oe3HtFvKGLPDigrP0kvw5N/GI=
`protect END_PROTECTED
