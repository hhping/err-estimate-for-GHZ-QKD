`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l02NMPKrrus14ZTaVM083GCkYutYTKkbTLzTdndDjNvYzzwR1qcKdChfzo2xKnPk
CUkhcha6UNUVsmXClZ0rjIHy1EA3VWI8XUY3PCYmjTrknpejGE8X447L0bVlaLIk
ATTBz+mlxcpND+nmnFWa41i0qQST2ii/xR6uTPKNk59UgvGVo6NTthN0RXxg1/FN
sehBVlDS9Vkgwtju0g27BlIn4cJ5mCxRcyjM4+en3L3cEl30tYZcbk13XBsW3vuJ
APjBEebRxieGbOr4wS2PaZK97CS2waNOv8H4xZ1t4qxUe9IfUej6IFVxuPNiqrIv
gXbx97AA5iLfOCzFMYn+W+5IaGZOJ25dTrVWc3/+0bDZkGW4BrCsOBn2qDMZ8YSZ
hPpDThDgHMxGXSaObUeSpZS+6mqqKm6dTlsLPd19rrazVyJk6x8KBvreqfbd84Em
e0Kq8uEMXwbDKulACaBOV3AdtGwGdt1TstG9in4miWrvUOUtBZcMRg/ko5R9TN7G
Q8PmCEHpD1LOCqCnO7WlePOf0cwcZCfk8LJntO5KFuxRUi9/Nv2EAcb56ShTFG9p
Tu9rkSDHwgqNK0fTm7wP/6Sxq6oEJcEZTBo5hOsU1ghqZ9juMCu1n7s/KKpDCf9/
GjPp0i7TtOIlslFbGqGTOiBoAeoRRAq877ZCvpvVa3Wh/Cb9RXMIQ0LR8jDZTkWF
jmu31fd6NXP7yriUOJzq1OkPTY6xnvDC+1sDiWqGQbq8bGDIlV0mvEOQcB5/nF7R
OBS42PzHq0n5BS8i46EbUoqf/xyKnKoVSfXz2r576Q71MAkX0YIt2LpDpttu6/nk
s7UIJKrALCQrJFvn6LNxaELWH5IXqOos9dS2TPMPxHPnPl7d7qIPlH1pE/4bdSIR
HEGwT2V0vnF7F1Ni1q8sfSPNPTpPu2XK/sXb7ZFU0hrdnW0w/bJN/UKKUu0Or4UA
OIx/MXlkypqeQuGlRbYp4Q1LH4vTxF86mEa1LEL9F8rAodlIPo0cbL5Hx9dJNTY/
KyXRxb8F0pt7OcEURYMwptUp5UDsenScCEn4zT5fVl3qTt1qQg1jstniTbcuVAjH
PV8wQTEWSNxVUiITi6fvpfJYrJmhJoq0juWh8ANgvqT1QI//LOXd75kMAi1RJgw+
1TtSK5z5dZSX96REaEvdg8OLvMHtUDdcWMfhuQIZdYq8feIoLT+vp3TCTZyWVrTo
CWpYOcYy3I8fsyd5FQhyWMwQiyCCmxSs3V2AiVxqh9A4Gax/YEEeF2xbSsmJWrnC
DKyvu3Lledlczk+Zxcp+RMyszZGcj9pWW8hNzkjaduF4wxM7uNBZ8ZtBPg7NFe7R
sTBdupnHBxfuhdH0Dsw1s0fBHijT7nx+fVA/AzPJgD/XKCqeEKBX0TUmmA8apQgu
XpM4uRes7OJDhkSQPopJl2mMUjiMUJYYH3tnZC5vfpkvftH32Z0w+wg2RHMjBS3V
RRAVmM2q1k90ysgBVeU2OdvQ4xwUYc7IkyC2vEnhFbkFZ/AJ/lYAeK8bffH0ZSYJ
FnNuV6kXzj+Z/y2oqtzHv5PYuIwYUEa31aFxtlFK9tsC0jI+zyZxTWEREzvjVLcv
MrKuxwXUot53KwjZ85tg3j5CEFh835f2FQ6RwRRHSsr4DIOtGqVMQSuJPaJ8KG5c
bn7ZaWMheN4MiVIudxwjPxz8T+TzXH09GwlqYNGbccR8AHqPejh10Wq01NI1Icxg
yCQzik3QaxG23c3pgI3z5sDD4EiEgIzGPtQBhrPyMWsGc3zXG0TvSJyxesgnlxa5
tfKxuXh0bLRM/Jn5yPTUbkhOv96OTqwYRbmfj4+mrKpj0KtpCTqCT5HBoF6WbxVH
c6pcFzspBQ0JWrOmenkjTX7NmH0nyN5uC4XKVQzhaqgj496qYOyJ9emvaEPwfTRk
KnGNy/eQQM7avFHQURhMoJc3Uk1gdNl5Y24b7YkTiuL37XLAe++3TBddlhZK64Nf
2rpI3RGsE/Bqr2pFtKZMa50nWjeVf7AIV6cwn6Z3YGHIAZWsKQGEmVvk5ZYsavkK
CCcYU/qPqlKukFnzOxPPmDPrOBhiJXsp4iWF2BzChsxEHqzmcTe2RarCd2dmS1x3
0ywsxk8KJhB0SjM4VsUn3chnjbkk/5PdcWhIDD1OxaRXkT70qSLr83Loyq2L9uFn
3wcFDSk2QB9DdUvqaIR/p8vRnZESk8brG7MdhjHhd/1HW+/g9DpEwS4UTyO8xDzU
9+wt4uwmKVlaGK+HeSOX75aSkWL9hQ6A7Yg8nn7KUwv/Md7fUi3QbMazimcjQsPC
m9n5d66vQzKE9RhcrOMrS29gA1CGFqx4T9PhQUCWPireAJL29mDvgqSQ3/HXWc2X
ZqvLL/FeHIssBDsP9gSLR5Ifpq8kc+W33f7c91T2lUxUGewBgPggwaXlTPqJ16R3
BXgJOnJ5niiRopEMq3C7ZrVX/EyoK9gmUWd1DJP39ej5H3vaQTcDwIo8M6BHF9al
UavQUEcKHwsjL5BcqR2xo/7Xap9WZfhSf86CfFw1nKvjh/bR06cEsdXzCxoTELGo
Ba0W8ZPUkFU5dUnGIRrGhXiMX7no64svOIp6xcu5CsuXHmIhhc65eaiIQdDSnUsk
Mhm+81sWFFj1npRxtF5DIzfjJNBRGicRkA8iZC9HEC6rIga+TYP9MfhGwz1Z7yPX
4AUdMY03K450oFNXLwMpy3JtSB9h8WC6s80zwcEGA5MUwXm/dRdXct8PEkod9c8Q
kgx+tjcp9oO4quSuUO9Gs+rQi1CXxbc4QaLrGodRLFS2q7fexaQ9621Ou2leiOHr
QtXGgWJ3u+klEmjMWwD6QLvjfnguwYb4ZwEOz+2vStWx9ECcR9ZGL6LWJH6+Dsi4
fGGm4GdEx2Lfbm90WBoapNcLjS9Zzn/p2O/EEfQqWvzxdJoYKFom6ybF4Md54Dnb
kkxcjPjWN0cFSEzyD9CuESmYLMWbfeZ0/G7H+MJkvf2DK/yWr3oMWhKUx+7nSFOt
Rrl0f27/0VGYvOc/eOhY+s2ISyBCg3aR1baRWuA0YMi3E6A0sQWycieUOwVefJ6f
bAOTrRgq3ePt41z/JNMsFXRJM1S/0dlhNmM6sHfTfH1kPp4K0/8P7gqgVbIxREii
ToPAxEDGyCOxctWommkvEldYLGj/6jvRwWs1Mfps4yD81dwK25tOq5AFoC5EQMyQ
zzu7OpVmmkLluCTufLCZLn+o0tzuciV6nx3d1avhH8fyw/wQBPmGNv260tMBWOAg
24zlo3lPF5+3+knDdBaO1WBSITXe/SnBc278RTPBWGFuhLt+43o8gdkpVWzacqps
fvb1be+X6uVH6fCJrQKYaESFo9jHx3zTI8O6hfFFo09y1/yco7PmhmXaNuxLGjNO
4tqejAFOak1IX+Q2FrPGtVb1sz6hEXWH3Y5qozEuatq4CrZ65TfVo1pG5+6mPnum
ELmJj6sixmHDaVbZ8RuSnhzLfEE3TA0P/4ZKrTcNAMqIFBQxZlaCbbKfQbEa+xMz
+6AgUgdcKz4L8V2+q/3usLsasPhUZ4GJ/tMhrFHaDc6W85xASapYauS3NEPGfFkw
5nYnsPp1WTT+fS18L28vLiaNlI9nU4mdVbIplryz/cV6XBhA0yvA/n38BwgiLc5S
jJZMycae/x+06ensuwIxy/NYdxKubvMndBB0bvmL5v2XpKtNR4iruj0wpG1cVCE7
Z80iThP8a5wcbJBSctPRyaK+4xZ7/+3uWSUuAM05I864dWd/gR6/4oO9QRUmSPve
2zDiC/HWZXGG10Vo+41cVb9Ayiw98k9T/5HO6AP0dlWDErYe9S+ubrxcWKaJ4Okq
IMk8Yp5myUfiI3h1yPjpDlsXMRIkCgkaHy3SIEq6iILz6e9qdO5gFFdmjXA5wrs+
h5DGAiWnDYdyIxVHT77C5yvhdn1D6ihYeI8yFzii2kNOuLOL6SCWNDl3eiXif4ag
eJGu2x+nU5f5jeGWEWTOkqtKzd9swU6YFQ33zITroFRJQ8kflxfGYpN3gqTrljsv
VC51HnVdA6eoo3Kd5ugh3OjewsmhEyevAthZvTTbSVpx6qb5HUw+gb1qHng9atcu
QbcW2D2mdnS1Htc9fU36P4+A5Kyd1qVlXYixK5PnfDT7IBfYa2BAXO7twX7ZI/sS
ayBTJ74IEkQdh9x6N7CKAZ5PeAjUKVJB7w/Y5LuOfMf4DCST2ePZhb03l5wHZm5E
T17HIB4/D5bu4NLUVZ21gGRm2E8ArkgrhWI1FMYe1UmdF7uBOsnfhKNW0vZ9j8pW
oOjDtn1Gf5JIwXH38FJpyj9Gne8jpA/5s3tS5NuGbYNRhnCcAjgcSKFW+hqTPtrv
mdg7fwj2NseCH4i9E0FW50ocbgP5dDVUhF0hX0D8W8EF0XI7hbqFacWdrLFiGohh
ABnAEIIJzSqxcbs7SbAbJxbzl0nv2CM9Q4G+f7WzQXRKe1VCWwtcmVlx5+Dp4zOO
JSUU+49nyJnIrz/ppHS4Z4qT3dmmeMKjr2lqod0j7/HQQV0FRUxtJgEmyujkIve0
81/irSBV6ujQDV/hojixCDOl1wvY95dNlLJWpD+unxwUmQUIl7gck3NHCStDdsFM
eC7MmSBjMU6reYvjp38e/Nnt2ya/aCGryIftBIcSmyhjZkt/sCb7InKS+viH4NRR
r4E5R6bjlo6jygxqhr5aScUHEarn+9CBkwY2XnZsH8B899Lq9XT0Y9yghOEhFnCO
DU/W2s4cTUTvcvykwZsDqHwID0T39fhQT9yzhtd6/3BZZUfvRX7EgqTNx5BeXSlY
5PcTxdo0pYcc70ugVyN+Sr74hY0+xbQIZ1v2Dg4OtmtcHDrovOpHlmECnnhqxEo4
8i58/Hpmms6/XsXoDOROQ3h2F7a9uP7krr0fZ2N6x576ZF6zE4uuodFhOdpNR8IG
d6BpytP3YG/qMRJF4CLpEhVH7d1MN+N+n4A/GlxGR6mkP+WXKPI6nYURM84f4Kx6
ei2pxcSqwhR13X0mjOw/zGfyM8KisAVYVknJ8fWw0qrO/KQrlnEEnSlZUpWzjU6r
/kgFMmUShDy98HBCaDoSFzwt2Tr28OckTgntKID/LWnlYBMvj52btg7OO6q/Kovu
1xrlHxA9XmVnM6mVZia3/TOWCbJZpUnM8eBMrpBA2YASXERKecuDw+P3CFpHvDCc
89D3ox5qjzy9fJKX0jg5032+EcH9dr+RTa1r5OIxZfiJc2S/Gy2NLE1Qb3ejs9Eu
7Qn4CbrrHykijuhl17t5r53Fnc/Ev8NHTJUzXH8CllFqlPWjUKTG++7az2GpFjND
N+Y3MJXVqqSndfrD5lj5JiQq/3TX4RGmZ+oNByRwzk1f1SNBWAWZydMMtur0iuBE
r6DbUETG9d7odEO28FgJVFQ/A7Tx7uIJU90YrsuGWNzAPJWgBYP2tappmLDkStKp
/IkVYhqAKOihUKiaJ/F76Cp57fUn8nnWvQK3JAX1EOMvVkeFXgGrIKsRN8TJRQFy
/l334RvuNoSi5CH/ruw7QpHeQKLi9YI/cGcX5olepguOOtGfhDGx6pI8PXvhFV8Y
DyKW3IqxcLYXOicd43TjzNSwejCYPyPmTWEXm8A4RauMIsTDyDxIsAUDcdKZi2mu
jM5Ty4Hceo/RPys9BM2Osq/AMw7OwNLyT+dWNqH8Y+q38hVUNa4o2DK9+JSrawJm
Od1vUwG9NM+XsO09KrWzKcXUu0C6dwxVfjSrNruh4vraDCuixtgqVbKRPO+/iIc3
htfZ+sNTekav7nL2B5h6Y2Qi2AA0xYgtHp1WhgurWbVpLQoO04xA3mgPBYU5+GDB
t/z1G1JaVNBOYo7G5ReK2cLlx6C6GbWIEDE579cuWavfqYVRJXx72U1ZFW0vLFaB
kfkGuM2tqnH4f+HdfxkCN3jo5EYuyQSMTAYr0mMPNkm8W/R4AoObdct+0rAYd/R2
xyDUsSjCPgQ21CMqOXbH8bSbDyWyYJY3LHAMKIj0Gdv/3XA1T7EH3W8osZBiP/IB
b64DV2wDJXXiwf+Vadk3adJuHfUaBsVIyglnpiDZtZXdAfXY9FRmcxOOtFoxhUzb
EcGnoTvYP42vLQ9iLRgqgqBGzjOQA+Ump9tggZkRhO3wAk7j1VtmpVnfWAL8HS+F
n4d6sdh8uADvHNZIUr0HiT/6rhyM6nRnOGu6fEzMmj584XU38AOqeei+2fvUcRL6
N/nkyr1qnf4HgaOHmWVLGZCBLKRbOzGHFMhKmCPSWhipfSv2c29PEZvmZzTfqV7H
mBsocjRf6Zhw2ly7UjAh5qUatqJKuqb0YI8uqp7sD9cPvmoFK10919ImfsWlbGPn
qroo4mxvm3VOTEkC5kd6UzU6Ee4NF2PuJJOrDG7dw87e3Cj2Wvq797SW3MTLbUbX
8jrXd/lbo6vqOJIqaRJ2xmKq9MCZdegwlqFGLIePBaOeJtI5Xrl7wVLKkEYS9hsc
/1UGCCb17HIIbWoVUSk37G/UP3dokWPBwrVf6Xk5jooT54Ls6tg0RTKHwpfDxX5l
+gDioYr/wQjIii9yjo+PxlXeUmFmmCCILnn1oA/5nwLPG2gwfgfXIqIdPdBUtnfP
FcileAQhy5C3VAdRcdVmWXfp++Ri4/4PMASvdsqfE2epwdS8sFdKRC3uJjs2pHgf
PNqrspkGXE+MZN5RDuMmUDbFv2yf5SMCMKCwd6l8G++hlR7HSUhGhWGdX7QDPwG1
PumYF+PJ5L8zPvnhjZ2nWPf3aFAOODCJfEmj1ACytCB9WT6AT12O33HhAxVZalQD
oyIs4A1yzBJLuq8as8FiJLN2ybl+NEOLF8fmJdCgzNBndetpE5sWB6TkDGxblZxQ
rL58yoKf4QFUj2w0t2pNwdKG5Wm601VpmsoVRxYZpp+vI3el3FB3Vhn2U2J+h/SI
AD+0ssz3UaDyLwjEvcsJ8UdyJv1UQb9asoqOff3yhlm799TTHju6th4n4zHhekbB
FjYm1gLH0nITxtDoPS8RGq2xGT/7eULHDwyjg5+ZXQnBDvQYHad9XnEoVmPpoyn0
JKGz8udBEpxO5wj5LBshSpzimTtP9LoGw3YPbSvHQ1BpxVLR6nczOoOzgCpY61dA
Gz9CDsR83kzZrn75uwd3pifusy//jL2RI5WGeoWkn2FGh6z0XTZ8CUJETkhM48+x
4OKNBNKYPJsAkHpiYlmZE8mtsodr6xBhcSBClV6qon6G95bgoU3oqqdrWUSoYRlS
v5SnDy6KK7eDf2C00K42zJbzxHNDbtFP5jmu3gzT1lCGQeqzCY08OHUwujUqVBo+
KZ+0nJLmT7R8YiNTt7ijI03u2E0iPTPJOsGWoW6AnABs2A7dEA3HhscDKdLUTFCi
7mfFgxMFRiAxJbJxZW3JsgSyYM/wpv64KyqrCoT7oiDP9AKsZyV0wKOi0/NrfeGc
OIQQqzxGzBluAUxbiDio/If/68NgA8MElMHJPiSx6KXAp9HhJGSgwOGY23GRjyjd
rGfLQiuuhWBxBHySFmIkz3MjmYW4AdMh/8vCjXhEHC2Vr/47UTaV25SzqEGQeu8J
M/9R2ewfArOsX+arxe9xvRwwjaodJua4yfVMbNJ8aMmXb8DH51V1+655Pj8wKP2Z
xmfVrktOyb7XDNXG7qH3VuV6n++HQzW3+vdf+rap4c0WQKlswrDqmDp5j8N+242p
tPEaT8ut4ie0EH79/dQ+Z42/rhrIjrqlHZa+9XC9cBDYouUQTviaT4u+oOZUPZ3q
I8UdpcYjEKXKfp9YBnUWylJDl3oIqFe4EB4gH4vCyE/imChpQobkmkQX4hbS6PPR
dhNIWntxrtcjq8OFr5Ms3otuxVfpsGcRSw5C5aW94AfuUdxa+TGd+vFtZdWmkKEW
rNKnycJLPHFKLlK6swR7kQ0FDHn5pT/ZG1Ep4fKQpZk3AMCOQJ/Ek3zHXD2gfhwe
pMcm/sKLcUgHTsyRRyHah+GzdKYwrUaZXjKGymKqKr68QCyLwdiBkTsIhTDS+vM2
nJ4Po6pVM26uNnBk2dkd0F4L7dgZ9ZI1nu9gbMtUE/3E6Ti/bAB2uf6N/kMDePyJ
J8CevRJCKvZVMzqQXiTLjkbUWD1TpQLxLMdgwXA8Xre4rI0kcFS1C2DwKF9Se4WS
GM3o6MU9e/93s9Dh+0v3sjiVOBcZOvJrkI4rx57ASXATbsEL2KLruQ4qPGenysPz
mb1GT7PlyEZ4XNsPjKV9DoN2X9IIy4rkhI7UJ0uza8W86Xc0J+dqJrz8oDQ8Odzo
cV8QdiFsJqKWXPndCRWTnGlchghlPYQOxNi+/bWtPKtux4iEcQkd8kKT/DcEK1rW
bk88ELkxLk754AA5+RJSarysUCmJo6TJ06BmeFI7ugVF3iTSYPbCC1oE1yzqT7h6
T0buiClitGpJJB5RSVmvDpq1oqTNNzlXQKDeMLaRtNkRxweDRI9tmXDcCvkEt7J4
K92guvDmKrvQ3XI+IKHeb6w3FpN2t6SijMfX8DRANSP2q9dPvBFLlxSxiXsM43p4
WX9wW4MccORsFLRUejfHiu7XqfK24C4YGpabtek383BehvuS52RBu532dWemTmTz
gQPAlL4TxE/rd31kO+M3YOJ1uzi0r+NO0CGpKOJAUeQsgTM6MZS6mQdV6Vzrv8Gr
0WwVHkQoCpdAN6ff88oK0zUCB4nVrQlmqvirat2qsyClI04W5vPZmhecDGKTO2Ey
hs8+TMvWXgbCdlYHv8Axl7/XwoIBw0CFE8OUndDaeOR1kY/cpHvAlOG+LeNrokaM
CHkUb5+PXzb1QuZZO7xiqF3Ovuls2HW3895jRLjnT1ro5latEbTBblkcLNps9906
CLwB2ZsndpnG422xoSYkkyaCPAsAkE1VP7bonx7aVI1lA7zYbvh0vIBzCg/YfiGW
/ju75FeBPvMwNKcuNaD/HqAKASQDw4GvGztnxsOUPkV57+X1YWoUP5SF9mAqaDSR
tpYmkq3HjikSoslSYByHuGzTBfy5/3YG8mGSlQWMqO4nSCGvLtJXwRvbu4bsUvp8
mJu/hOywBsC7hmBDVHWveYFfKlsil288kjTDkonWYKTs0bAPO+efW+kPgNfEztkt
/bgLTBMPTLiu3dbPEbmDOaQv113ta9wrSBXNbanpJX2xuo/WytgKmtZUdfQSTDno
+SUe7cUpvhXV1eoz19R/WS/NEeP/AwKN+g9Vj15/2vUNCamyISzYFIzSpSwUs2f9
s6QDHr4v7dBQm+7NkjkB07SBShL37VXVMX2TThGv+v25DHX4faf3xZe8Nb3bFs2w
4fyuVG6rJjBPJI/AD4PkZvU2RYypC2eItubQGvDTTJDGhB0zfdqLKtUq25HRmBR1
r6qdwJRJRKMJ8XcKNxpv6AB6nWyIXqSq9fe/oU5MYLGTX82OPWSBEpW9jO50/G9B
dkC32IOVftNfGa6aOIT1TpVNCkHF+9ZLwFgRcXA5NyZtYK2FLsWS9785NQ124fPL
3k1i7EHcyCZJaoHya9gJZBY4BsdGn57PvvBiQqYUxooT/30s5ARWMn7HQXG910nh
efm5B27G1tbbg+Gz/XtAKhc4DJ3VLqtiJidhY7CYs6Y/Sf+tlaVV+d9KXDoMLdAb
o44uUeo7ckOsYRbjTZ4yW4JE4eGnuvb/papGLGp5d+U8X2gjOfgp1OxYLcMc5kF4
znkHdU6cALiILkjixkFxkpefiV2Z7rm1xGC5vbJNoKguGEHRU6N4RmuSjDDR/bEk
PgtMkEqbFvER0kxMzuFTM6AnBvJf87B5vJt0iqIwYmhOkbu59QLz6SfO071X85CV
H2e5E04pUECnyYTAajdwLqzllrBnEtVafc/R0cBCLI/+lXfhK8ODY13YUzPhQaN1
LJX6u1f8u3nS3XHdjhhLVklpcokl0oKd9+W6ycZc9AXoew/PxRn1ox1IkhCK3EOQ
Xk2GgUBsRAiHLKkEFmt0VUzfqLBMQCVHnN3mufTZ7dKnwulnih4xmII0pus65jN7
VpdVZ57AYxHk+pfJ/C9iStoEcaaAEm85G1GvF5rjrvfVUtvDoHa0Ec1sA402woXV
yGfsvhDip3bJDKwWZllduZTnLe+5k5sFLgq98xqFuIPXGvpYZbA9Z0b+i28QvAzG
sNVBZF6omLn0N0UdntX4zCMfEfrm7FpzqbRmk7ME97Dxl2SB5hYcjxPbRcIbHqwO
aU0Ej0QB9dj5uBAskNm6a9hJttYd3md5AH1o6KN6UkrvZl6XVhRoAHxCxbEaGXKo
3sweLYU435ZrHOHNuclnHLs9I0yLSwXSZO2h+TG1DpHChntx2J1/U16GAqk9W8Os
nf6Pf3wpuu13Xs2zYleWhRDH0KfYCu1dXwOJ4qyt3cBIOCLpUgq136bczTYxVfTE
gOdXpDHKDpsZkY0HWwkt4t9PT24O8T65WXGwZKYYr81KKEPN+SYezzMfTR/6tvix
PvvaKA/h4s9NfVSFeUPdSHq+LssW6YTga/gdwehPRAJuiHyTNiuSlZCrRkuMMW7K
r9yAFWuqLbxGpWWMsmfY1AwAy4dUDlAUymcAC8OZRmeLHT4jLV4JWEWO4rq1r+Pf
BXIydwpD9Z5nskDslzfxs40riwukadfVLmaEiaJkMn2RzGaeKltwTraKV10XLkAE
tFWhZZ4/+1w2pWDW827CnGSfyr8Ycl9SAT6BvmMMfTzhht155wPhthUpIvLiYTdX
3JxdDjFBPGUclz3Tdkb0rKKBwNViPzR/aYNd7wh2kR9Zm99BCtd2sfQu16P56ekG
0mILzo2u0Q6EH3CmAXOTqJ5JAoZHdFwooYdGdjDhr9hLDtAzlkx4kJdk59YGZQNq
Irx7DVkk1HonZ3GzOvOoajXtArPg4l/8XJygYhGrmBS7yweabR9dwPhd6XwvkrRg
9jO40rlxNk1gMZ10olS5hpRVWr5XEfFY65iR5MsA58UQt2Zg0KF8b7g5SFGm8kZc
bG7uXc50FNssRIRJKMbGXxJq+VLkiynKlJU7IWocD7/mrRH2oDkHg+vbBeG8SF3G
Gi09ccvljPgPEuTQ7qgR7C3g96m8nXKpzq2pFVIlMuAqAMLeIY+8DkfWiiVnavm6
JyOKQYeg8cbApwYIEI/sviOw21amqO6jevoAxEsMdr6rrlWhccqjvI1zlvYnD1Z8
YiNZIUehcPTAhtz/97VbYXN3lD3H9QU/aSrjTMmlRTuqdgbQ++jV+GAcz/sfK/VA
cfFTO67VoVn7K3Fb8nHCX3akqYs9BGyEZ1NN7owuNrQvtILK50JoiV8uTTH9POEI
6i3/QVbaa8tHP81JFfxeH51JG4H9DqTe8nNJowh38USLRmKja24ZzZBdsi+i+sSG
pdHej0vKkv8QZ2RCjaAlG9YYNVSXY5AYa1TmQ4+N/FSmWF9MaHU6qkzSniFcf7Gs
wWYwQZIEW/ekVLh/ggBP5p8fRkNvQPzhV+gp7gK4JHjCD4X6R5uT4KEQ2sLnRpza
/SAvYdFd2o+ADrwvP27b3M069aMzqwkTwR/mf0r5r0zV8hBtqnS1QaPV4Vmw7DIu
LweyDYR15y0o1Ckqk3rDbGtXFQFPgrI4G9eHWz5IdVbltv5zACbgfLDs24gisZhC
+lrzX/FkSAV7rg4cZO+0xtHVXnsSpiLv2w2ZXfXQoUa3OlD9tQzgCzOnSuEsGDuP
2CokTGbeT9ffc3vVE5xLnVMoX4sk6X6C9iH4g7cJkKZvAPH3HmXtNMhwjZxYEhGY
a6w5RVSbuJuV6qVIolnU1Z9DLkdu/pZ7q4vFvep8LJNVahNC7SFvWlzhJnaoBsxT
0PUoKHnd3gHkDukECGCUOSepIExk15SbhbviVHL1snry6pCsYcj2KIOC5X8LrP04
mnDHj1l1h9JAmH3o6xyZFZsR9mvQ9f8wUoC8njM1aIfDLnUIxjClCNDaEbsr1pHD
aIXVtmSS7yzGG9xbEZIhNkB9t4lm3aP6tyv4iTS9jHrTn/bR0hMT6VyNKbyhAlXU
aiiybfp5JBECu8zRDBTPri491zC23Oogh+gpSuWvthoroL20xJfUc3V1VOXYH/mI
GtQijBQT2eq3P/Kut13nzWVMsW3tRdZlQX+pW1iEAFmMb8+husDNPStHIfu2Yoe2
hEBKypVU7jeGJ4OMUXwci86WcstU76XM+bJlhjoKK44un46hvRtu73g5RHXWc8Qk
xwIwQ+lVR9H/Vc2Vf3LHBU4/C7NmBFTCqahGRextNqjKU4aC6+xeo13E7HAt9DWB
Na5rZMC56s+yW3BOtgsPXjLR8tYoto/t4rtMu6P3qy1dlllNYTEptKfcPJHnjkkL
A2S4sWQ3NrO0jJo/mXtRtzeymC/ciXsMlbJVXcZyYlinXf4dLJWcxWps0iG2pYJA
8ADKryulUCzDc2aqgsiHnkeb/eaFmXJUPTi6DQNyZjRgnNkFnCRb+UcYne+gS+4e
JPoaEX/KQqNT5ICjmjGNaIJZrYq8sZDvRYTPiTkQohNdb9rPIB8dPwmlkp02IacX
VJyl+lud/BPgV8rzRK1NCjx23Z9qK3g1A4r18FXbCy/T0gWaueYJP3YIoL0QfCi/
GEsiy7pTxw5MlCTWf8MfELaFRwLgK8K3e31h+XbfeHgGGwGqAdOVHRPxHBdUqAdh
/emht7iUpeaitNj4IPhm6yuTSlnqmLt1FC09bnVodBh925GJuvpaXKhM9XTobzNw
vbFZqqjokG2jHC8DVAImIg2D0WSFHaMGSZglCgGA+2ynjlz2YF/3hs/P1LEpTOOg
cX9F78+iOppbxoHQCsrcm/nipRq23EBukUKJcXXYe1p24eTRhE/QIVIKOe37W6i0
JdBTVotB7XjB0SkSjKcFwCzgsH+L0UQQmZTqphCB9DIKMs+u/uT8BB/EQX2uFFMs
kGq/UFIXPgk82Y2baV+hu3ZsK7ZIph7FgMGRYGIAOAA+FhH3+wX6tTE4I+w03oec
+ng59I0hMFGQg/EIMq1c99e8IReUtwrnGdLOFJtPFcXiYJqtTAnppUQwdq1eowi1
8AwWIB/bZ7ULwwjGi7Y8zfLh5klZf4O2c444wjg0bTexTVqEYX3N6l4UU7uYaKDw
HHOHQ7YKiRUGz/BqMcZwE0TNZF8VFVYAKMjquLgwr5frEx63UDSsxCgBLFdUUZS1
9b7eBEoEIbusFogXjjF4N70svveW/UXq9xU+gFXP4Xp+xrBng5lUcGNPl5M/XPN0
On7SyMXorz2mRBuBXCCfdvi27U/hM9pJYZ+LvAExYEaIzWV6niih9FBMNdxSYySo
lK0b4avVLR3aZaB883C3NdPYwojSNXMIFjGBk2YG/SWGx73djJU76EPhyYNp26av
q3i7fX5RIxoja/0fGfy4fGwWlY/KH7sElfmUZo54bDngO7BjS874i/wgffDwqOmy
KLklWWOVqhWgHPVKiBx5pBMSC7OYb5Y9UIs9C35QgMxWWMoYsx33G7wwrXPBWS+a
Vd7lbHcWKLYzlzxhRqUdb6LhcICS7HCV3SYaW3qzzDjGZTnPz4DVJUEBnbLlJ81J
CE4y5W5TZ/leboDVTEZRCp1kFSbyMvoL4pOtzubM2bvjUdMrMH2Z5wKzMP6PJzl+
LFKpkRaluJ/M0vZFQgiqskvkf1rEjGIBmQh/cXecf4ADkqwdRTv41uXxXM9xJQJQ
TZJ0fJTOICy6ZMy5O2bJ6U44o1PUwfpBd/5SJbjszScuVJaR/GeW7Y3G4SnDs8VY
8WTTUbImab+vUREcA/1qSxwU4VVsHkck/QVLMruRgsmMQ5sDDsDQGW9XF9fJH1DR
drSRzSLPzJgFPHDWW2Il/78GE9YvYeYG3MuJ6iTMkNGeP/C4Sf0ERzfzFLr6JzO8
xLem0obvFqGK1iCRZ2cSpAn32oz7hMqKjOnjIP1Uz6iJY8eqAixtteibZq7OsHNv
UJaSF//lLrOi+Jl+YS+wPiD+/tubZvDi3Qr+cG6VHU/0Pkhj1WuoU2ag02uSiKJ+
4s868J2Mtvw5cMhfwuzD+YM67fAA48P3s972WLMqEUfq8+thpIPOZDu8b8t/IH/p
ODdzta234zCtuPgxxyi5hFfs7mBIWo2F9cGYBkUf2EEK1RCv+sXGonkWzCs/wDGU
RGJgzQ93CSMBCN3NHrSApsVnoY1rSrauP0uW1sAHqvNr12gY1TjGdUyAqD0YPeCY
UI/LVnr+Vx3cBqAra+vXYkGRQLvV9StS9OFYYZ8vtiTBT/B9L51kucwiQn7M62qI
aD9zCgtSx6HINhvk0flhZy676Yk8OASRc//BFixTl9fpk+7GgErr39bQIvIlnJZL
GQATK+OcqMeOHXwkobrPjt3wjdhQalslu3cVDfN2rBGSt0wWnp9j3wB0+YygshFe
ji+BzBf9s2w+BX7gVYQkW6r7atefmNO/B3J0xn/eKZFc3JZol0YmZ1m5NkoSVUjm
01msDq4jFi7wNvLI0qZUh0y2017q67pOH5LgrcXslXxXl90k9/ezuO28lWkIOx6S
+kTeTmxrnPWRxhytZpWb0dPTXJw1m9kVUTC6MsYn+0sunTqLni5LOp5+uMEXl6IG
xxO0W723EzhSC7TLG4V7InWqGTtDS+xlbLQw06BSogERMhF+X1TaVRQcq6wGfTRV
iNLtYl00z1Fc8+ettG2pMN0fVajxvWq6sO5Smv0deyfoxowIzCrzY3I9TZd4Ka1y
kNYFldnnGg42dAfPU2eNdDWlqDf9WLdXEpuFYi3I4CQCcZtSfnNED48+snk6tzg0
t0IaspZkr31AAcef15oNJRZvKyiVMRJIzmaWXxJHztUvkeZwWJho9hIzAxmOqmtd
qAvzfjubfwS3/zYRt91bcb4WV9A0hQpt93SxFnXhkMNUsCnI1By292pDulYjK8gE
Ck3uLwVYq5zh03SchosUThp6DU+pv88ARRDVOpMNDHlyB0qiiNzOHqoPVzmjhroL
kKXL4Mf9oWLL9RAk/zfBhFL8OWu5JBl6GesRS3l6jEyIfKRDSALX1LC5Z08FvmTA
NfD7j4WnkGRuBvaIGL7K8VQfmLqA5/36RTcXaObjGyjwd1pUcTGBXTkeaqYbCha4
Fjvjoc6aH5EF8WY255JvOx06Cqw/XkrrkPvafPOLpqTHmZ6VXXqiHdB1v+wcJaHE
Dwntrq8d2FqVmKxYvI3luHa2xat6aYdRtjkzOgYGOSa2DOj7bTYSVvi9cT8plHWQ
XNjm2MeYWoz+O3l1nSA/OxH1GXXuf8C6sr06iBb3h+AA5o2pFQAN5UdnlMKCgTcP
5eMSwPnDTQSdoguOl9k/w7MsNZjemSSM46ktxgF7vB2MEj2AOLTeWKoNrdoXmYRh
YKY7vkDmul0qkNSyMeAF41eQbcpHF9RTJIULSkNsaYt5RF/xG26bhgIMwf3cByIg
nVDzCLXFxyqw58hhqFbsP87GhPEV+XONudYHQQs6nXzHNhTpPdfA0/ptKg7Mu1sK
DLQreKuNFkSbKRRsaHW1n+V7/EbnBMA8uhkcnOmwZGOTaI2lUURfwLYzLBKF6zXp
HDNTBr7ivtLxbglkenRnIqPH4c6xaybWrRa/4gkYlPkgUE3AXAj7UVJgBOOSecJk
+/Uluaes8jHso7b8L7X/TGVzO+m+IO5KenIUhGF6RSsAnkF2jXDoS/xiZ0gKifCM
uWUYV7yp29rWATh9++DD53XA1+FgjaPRM4861D4P1EQzwo2auR9ZQQx7QLyuBhR7
WorT8Xxl7yO+vHC8Jphs2ivBRGA7Oz5wIa8e2l6bw2Ld4qZm/3BcCdTrEoJaCrX5
8qIgjS+SRykLuGloSCEcm/Y9p11xEL0ktrelGT2p6/F9a2wjTlQDdCh9o2oHTZwA
QQ0p1U4g+xqZxfhkOnrpOMOvSF3sRgSv0RY+oPhckvSULChOVVqbwEqIx0V9xOMd
trEK0nFHQHF1uSA8Q8nsRe1Ut29/XvgvBlswHywfBqJ/Ieh9dXUik1SmYwBXLMJV
t7fMQHmWhxIJHgc9PHWrICHXT2vbHeMdkwFql+iu5qLemU2P/vzt2nps5p5+rp5l
aM0FtFA9W1jPP4bLY7pSPhU3tqE8yyb1t3p/Pu11NeLI5pu4TJwWxsyOdBDQ19I7
D7maECVsQivejbWMlrFk97vFjV5jYxlBJyrk6aN/xuXZZlaCzayO1Xn2B1WQ0w8A
6pDQp7jXrzX+ghqI3XakKI5OrPsv+KyIRuArGmf936Ubk/5efjzmkLnc8mUX5fb5
PnBWSAmEEjeG7gPy+MqbEQPKtOWXLjm2yLp0sLuTXmgkopW1ym6GkgE5H3ZSdUpt
zUQgA9cwxq7ufLPSSinzLqdpyOhNTcqVV8y3JhIclkc2H3N9eufSheiO2R98IoyY
19F8E8DceO5lBrHphB9lBC7i4I1f1hl7XxP5pR/hA8oiPVihTDVMQshajFEYHDDk
rGNMRChX3N+3oN+N9Z7vlTzXTcHu07fsK5p8fV6cFWSgdSPeO64gCDMdWn8dccRB
5WhFSQ1PnKBkdpKFONmwVwSRel/+Vw9GpzYfzsX8oRidvXm+fUs45wnavCX8Pw38
uhe2lR8B0rwm4wtAMai5GdzDQRZdArzxst2ZZS74U6g/vHwevZ5SkjyOqsIgnQ+h
G0RNhjRvpGlCgjpIiDUhm6IYfepcjSFy0qPUa+LqK00D9jjx3K0g/IiknAb5MtCz
c6DoaNZYfQoUfK8i5tiADFRBWojPvMGE/CMGQ8b3YRE8+sb4h9A/MlMzhVzklnAl
8nAx5igvJBI+F3M05gp0KJ2op9TdCKNwbyyYAMA0Nf6aKnZrfj7CXZvXV9mqBnps
DdLj83Ugd8Bf7l5n7WUO30tN+FfKegxM2ieSABoqZrTtpJ43My/fUJX0unIF6R36
+VZJwhy9T8VvCjWEZNu/Dw0LmJYEh8u6jHpuSIOAkJ/+tVENIKk67mZi3hMjzlWu
EEs9ZEQsCY74skC5ae4ScLpkoZ+qDGl3lhEne5nJUnCm7H9DaTz4VvUgssLgkGrE
HdeS740kPRxAaiP2bvIXd/nkNwz22Ua/hKZnso7MMAHpOvpD5yINrc099FRwS0M2
ZjpxenCnWyMSeLuVt0qMAl2LKQU9H6EDbd4AmOdIOyaFd0PwbU+qqxY2oHbeOiA/
16lQ9rIV8nJA/6kjS/XdFbZ1/1cgmWmk9lIH2Og+9m8lBv3nWvb/hfZ0hUus1jQF
PfIiZirUvxEIdUMNfhKCslETgxM0x95N/Y08IcPRsSX8b1mYC3qLxWUouAMgl8dr
31cquXgjdlYtgelOZjfIR9qFkel14QW4Q1a2z+yOcdpL2IBKz+5FdMD2jtrAL7/Z
dJlc+l30j5ydf7TOUx4jzWMLzXluMAMr9AXMvlTkUMk2kFRvLPnyoGVecThensX2
LRE8UZnd5zh9FGrs4hkzJwmGoY7ViyMudbACAunDTR4Ua9a2JkSMfwMmM0cQg2nK
vqHJ/iHkxeCPZ8XNFr5YlojnI2Rc20FlC3NI58HvFm9iv8zsTCJtZA1pg+0CsAsY
ByqnTdsKnaKrchYgc0uFKxYjpH2O9XFU3/4BDxqLjxXex+5GI2nzPweJMKEx4y9a
7slcsXYCaOqUBqqZlI7vBPZjBXzv4zMZq0FYqREJOpwJSU/7ttCdszQT5Q76p3+a
y/A1Hzx+BUSNQ2sxhD4jWplb8Ww3/ejyNMqhHVPMlFeWna4ds9xQ2kYmWsAccdPr
8ACxK+eXekynA290MGcGnuYzD3gXx/tcPqFK5OCBEScGVyG7lRw4E7P49CjW5NNL
lAruE6kqVnUZv6deP9/ZA/O+1KUq2Y4c5q5WRGR6Cnk54K8Px+V+OVOjcKt1lMRB
dpqWA6XBYxqBNKt9LcJwAr6jcX1Le1BtVpPOLprMjenFlJisdVUnNEFJkoF3IF7T
3kJoKRRqzIHegmwNm/7yT/KoUlsJitJjAAtx2g2Wm0UXYCktmvSf/l4iA33r+SvN
lWZAYdnGFiYin254QBYDPCmJh9hOPv41OvLyG7Dx505LkiYN5KNgesvjcjjnGyO4
1B0RXIY2fZsSyDRJiTn1HfcKXoB52buJcbaH8m67f5QxU51GjjnyUFvOzQjVrJD6
2cuBVYuKIlAFF35tp1qTk+yH/yLghbw+5JkNj7uN/Xw7RIqDYHjwkMj/TmR+xIaR
2oCxx+ZwWvelou0r+7Q8yXmCtv5Kj4csicud6l3yOwD7zu6BuxJohbLPAt74mrmo
1LK2k1xTClUHH2fFOqdwCUnh3JxUWwlTtlJJUSAMm268tA9D+R9ZWFje/I/tcHd7
wuvNhT6u7EYc7DDf5v4Wap9iC5fvHL56gKRT1++ta7b+XZtTMRI21Ozyv60Q66x0
9k0bZDqz1hBudp5renTUA0Mt3otUZLmfq5OTiexx0Pdzn9YPnkudHukfkR3XP35e
gyLniimSeYfYCI9omnyVEq5gkmN/9EehtOzMh5Na5bhldqq/wM/SuXrzeVOOxa55
evbU7Pcsn5CDKvR2L2OKBC6ExjIGPdBgej26skroiINnhf+wbvd1lzCthpmhPja9
a8EZudohnoP17MJQ2KAkLM4gRYk9d7746ECH/ynURBSm2IhpqVehzC8RdijjmxQF
Rpqz7xR73zglrT6aZmjIgtN7qjoLubap6ct/uLYxBJHhCUmYsAInDITa+efb/CvB
t+NpSiCba+1Q5p3kwZlj1ZUjJp2vPy+UtVf74L2qY0kJB61YUeXz0VTEzx70a8c1
2n89W7csjNfzJmGjJ9kNlV+zJQZNELNQQhv78TN4me+sr9SN+wfUrDlbgDy9Ot0W
aqlfzukC0DFjL6WU/RGP1RQPgfWTey51QxCGZRQQQfjmUNijMa5Ur7iK7ECdtrs/
FmI6Drs8p7apockaKBQYWl/TdEOBmKfeHno2p0kt6b0XXwjw3NImxk7JB/WYaGJP
6IVKeuYe0G8JxxfGxD5BASBkbL82mLBfAIIMLJErqLKjU+VZFWF6QgHHoL4dWDGZ
K+Qm6TqJZ0yGZ6zVapWFq723HAqJMdxIhQfYv8B1hBnTynV1owbyg6uHOE+yCcup
pRO7CYdEqUSyQY19dAD+5Ik0CyHDm1oM0ZMpqhy2NnNaSD81z/99AEMpCTjTZk1S
gLe4zKjQt43Akv23Dl74XdWBxULdlj9SdKzT2lGqbA38TgZGwWgGF7UQSSnVHqSc
FBRA7q+90j/mvy8JAJfqLi6iAFuPnihFmkRHJU0CxvyAWJzhEKNrX1+jzfCYnnro
kXif66+k/WOSyziwnPtcyI0DRba7SPNc2PCRzRlKNDFHaKAAOK0gm2Qgu+a+iZGg
45KGTNQyWaqLt1LT6ANZn58k8RHgT/PU45lE7uABgsUA26rWBhKqzrCvX7ILRkIx
LqWtoOh+dEMjdA+sgB7W8EFSGRrKczaMr5mF6uTPsM3FuF2tBNnBY5P0U9pTV3dj
8F8N2gsLkQa5yZ3s0ERGx3XFaCq69Qb1RaJMj+lcITUi6yzyCiUuEHsD6jn52Cja
qYHVTHjnCxyviWzpWJ9VXHHu1m4HX1syFnv6bN9yrJBF/j09alYnFExYkQlkJLSP
MzHDBZ0fDtwXt135E+rV/pzfAdMUauRkoAdBnpNlX8UMuG3iQFa/09N+b1XoS962
BMNLMVFnf2hCMOVkEwo520+TyBhgO3CRlHY5AI/X3gdA8KMhpP7EDb5dnNncxpVF
8Zk1RIydynyLij3XCrREZHb/uY3T0hHs3OUTcyjDs03H1R0R2dB5KhoAHNkqL5Ml
GYqpiiN/vhI96Zg0pqpHHoA58ldKfwDhkYqMgQJDAlr/4ZVBlZbMCzXp5NxY32/P
o8OmMJHAdHMJQzaK+5qcjd1YadrU94Q82O9TWDtUjehb7qEu79lLEHcK7z2cAOlb
5OCt1mHzhwbHRhinlzKY9RZwCx9RpdRuiwtatSjTisDcQ3Pja6Mg2wEEqzWht1qY
ozZgvKzQLttj8OXknk70qAP6wkVcdGtsgk8NQqKVV7KijeVcras12nuyle1v+P7+
vOi+N0iz/i9GX0gBu+27mnTBWqiZSAXISDtPxYxY0+krkUWlMDvJ9lvAYyNYMK0k
u5gSrPIohS7f+gvX4ym3WYlXJfTY8ATrdM35cK9P5ilQWy8KV3RWq9myFzd1bRnZ
z1FzDdzCQTmOimaosJMGuJxanA6eSdsQtH22GwNvFtweT+VH5JM1LvTvFIUt3KnB
C5wFv9drjgfqsKVINiC8iot3w8OQ9HJgnaAWW5bSoF+59YgdIfxjWZTv/HsACUZm
/V3qywRLcn0sRh7rMKUx2AHjtJrWUMKkvnrWGE7Am1TtXEjspOy9bx/hh4l1KarA
34R8e113LD8xecvpoxyeHD22AZEb5eNEez2e/ClOvya4PH30r00AhWSlq9tHiwfc
DZlhwW3XGxBcfAa1D7BN9GzjBZFcM3BBHlCygEYG3tvQkq8FdYa1XpRDq6quKQIw
W5kLQgAhG2zvwcB8L3T2g07Do0hEMaV3CwgbRAmY9eEC4YFrjXgzLWRzf7SpiYXN
jgFQcWpPC/vJih4Vpcampv+PZRRWH1Q9M7y/dJPZk/oyf62P/TUNKWLVmYuMAjnR
qIGVEpWRWRAVtZLMKUCt82i1aRFbDgWv1WrAEVGzmntR8grsVWFGjUPaiOxdsoCa
5PXCmA+Fkve7o9Ry1cqUWcxKnFYezl/swa9PQ4yx5VIM7AGib2pTu2uxAllGVA6o
02m0usc/rGQp99DV2FYC1KN1ekUCpN5W+7ER286HbVy9SYbOppC5uQvbHtQmgg2e
xpgHmdCdimImOwwYLw26yOZrTshueNECJaJFIaGfcwXD1M9a/Ga7aJpCCGe+07o/
IDblkmjiDXunCvNCNE/Cpy5oTe8FdIOYA8bGzIFDiAaqjq/X4QKaYpjx917RWN0O
kta0dtH+Qzqy0Je3H1mJnZj5DZpHlrFH3yY8L01JILsbeOIZrTP8o/ncDFAK7BKA
sFmFqXaRC95kO/BEMAG1J4RxhmTH6pdArAL8tA3oDgDE0cf+29dH5/yahTHmE806
pqUsl8hl2FkJMf5/DLQZjYwpq9Tpsq3gCy2JYiYWIjKcLR+lpLfgSUKpHFFAPrC/
DxAOi0oRynMkJtUtu739Cvx+x3YCyql0a4LR1uujljmvX1HakYiDBrXlFspJVQ4B
02+r0ORmUHX1dE1yW8+yrbLE9shD8h8eKzVFCLvpLIh2mqQiB6fXkIWfzcc290XY
Ip9n+ebYPZeUyZL8LeGkFgsqgPNkjuu9upZZ6wkiHSlU4SFdJtrMYXVOmRgwBPcs
GPh+ytDsSXFB6Vn9aMJiRzEMpBVWnQ1dJ5kAhQfSIciD5pOgYxxPmkrtlWDNHVmK
mP98mBLx7tdNPRfQQTzs8UP3CVdgSjlEnkoxb1klV1GyzV1lHzvLejieUlU3Kbb/
TY8nbUzRktQT5O8rD6W/FG+d3hZEJPIcukXI1hkklafF5+AuYYYIq4nD3rZWwU97
3yBsScMqzRvnwVUT+TwpKM3g93x6w4RvW9bOtoDPxTdowdNBfXaZvrVQ0IQ2KeZk
2ZIMpSU9q9fok5OYXXDwJ9Lh6zcKufRXmmtVEbfe/o9wWuypfoCHIeu8bHo66pmH
TeJ1xcrM6NhEmk0CzR4uwG8vqFK4SFCi87G40UuBcezh1TJpNXYsBmEU4L1Nju21
P6CwOnkFJWlvCG4xttOOjwdnFACD3uwLtxNI8S88V3gNkh1yGUhrOY5nd4tMOYFc
RUvhaOvyy91XbFPZun65QYTOBmYsRSuU5EKqSepRzmOMU0DG48FFfog3hKVqvocx
G7lT31yW/wA6mKXAzY34pgG9hXAkyYFK7Vu/c3wMgJTrUSiasTZ70YhA7o0Gmwi+
AJhe2zrGPRpaESxWyaqb69FfdW8pHLCoTVIMZqIIxGGuVAn7iRiLFPfGyMTnZY4A
6+p0gQrIAYyC6nBuMeSfB8UWcjEtyf8+EBhDZoHCoLBp0ANgqrXME11rngWDZ3iB
2OUI0poCXgNWpVE8G08/sJgk4rrCLWMv+rWA9/teeuQ6mkOHqoyNJ8uAV6oGSEvm
Do8TrknZp98V/WlK97gq3/HUQ3FHKPCc7bwFjOAHfdbHm0kP2yDlD7iC2k8ZD1jj
c+jc4DJhZYDHCbTzZxwQ6kV5Z4wJVs24Je+AzSiYO5CdGHrmH6NalErYKWPniz6c
caWpq05rfjuyjcvqB1BWKFQaau+evuMcSz/Fo+sbGZYQhq5xRdASR1ktnr+FrHJY
QYuqL+/4ehHDf3QMUnqpaML4RFA+14yNKiXVf/7UmPOZ+w5kK0I1uPyvIgugiW5R
akPXlfM7OLaLmPg2zmHhb3LsfDir02IA0FDJB26Fo/6F6+aDanKeeAKi9NOuZOv7
XeTEfhKessBS0of5e4eG6hkxGRQJydZDfyyfvCVjrj0VNxlQRXHkPBbmoW+OxbQa
LKGFeKnUSUV9TWsVz+wKx3LvkLxovWuljvpGK2zNDKjGUtsyTORi8jp/eD4dyJDh
zV1ZKz0IU5RHOKTfj6SWhj96IrTjNgFisLHL8rFd9uUdhoMhL3urTEhj+tT9wrfm
mU5CvLsNKAS7fD4Bm0P5X7ajmjPMnzYCaM4E9X2tXpOCzr89Jtos5tve9QmWExqy
BmFGpAMrZxwEZx9yvM5Uodhd6FGxVsq6Ch3fDlvqgRtKl2SMvJDN3VXlXy07jBFD
mEVdljnrZEntjxXsf3/kLj4H1c8ptWNlovQKC8trhWPTj+c4P8bPmPDAwGggvBZh
hdYy7qvCaBx4eX4WpdPQWVhDiMYal2tdIBQOvbmHKW6HWV1ufKzX8on1f28Ax2tl
3oyhRQufm9EQ2VN0HMy6PC6zW2xJJhbD7HHdaE1e/rCtoJhIk6xKZj4UD7+2eKed
F/RzMD5+Kol4rRu09JwLwu9tshopnXhxzx7k2OeGUitu9tn3A29yGOWhnWdAgrpb
/D9y7herxb/reLG911p003XQ3Teypk+ZCJQJoPBAl+yrm3GAq+YeYcQ4ML8WXrhB
gKxzPUcBI4PJpMiF8BUq//FQgsFaV/7nm6FjrH/OFmJX5G3s+7hsb0uWM0hZzelp
+K6/KfeS487xuC63onjSpvJymf8DbVFSqhnGhr4QQG9QGYb9/08gew8Ggrl0yo2m
WjS5myV9G9gN+0x71qvl0BB1d/ONRd3ytbp2OkIt2AGmtwvoISTt3n3b8fx2hDoU
5QjSs/MHbCEak+aLtQYzFihNbcybMn3cNCyLxVwMTk2VvtbQSqp4imXj1QKN+MYz
DYy7tXJ9GuNWFFTByKJjrvSPJo25g6sVRa2c23/qRbeksd6UeAs3K66QBQCaAP7p
qGUBgSXJASUFKsTHW69lN/46KFEsk7rn/51ysjcRjsymfU/R2hvPRn3OhwcUF6NM
Gho30QF2NAdHg8COhT/dW22kfEzVbY8anhAdW2HrzeLjzZEmAYV4qirK4cVBb//n
YEtraQk8vntjXyJwjY1xFPvv8AO/qTaaWgFEVVR7JmxNtdTNly76XWWa8zBeIdA8
/x4Z4GJk10bsDo1Wh6fMUvVDhIlI9SrvzwDPKvyy0Bz3uMBodoh6Tr2HJZiznMyv
6FUm60PFuD3ftBCBz6Jp6xRF8aftyfb5nAWBpg5oKWufVtYgJBj8QvYZtAqbDCfl
Dwhtir+8vueyaIGOu3WW5ae1FD5BbZe1cjn9sEnD5Hn4i8m82GZCA+QT/OorWQUW
DVzbxTmw/Q7CQgT71xYj3aEG5bcoAQd05BN4FY5Y6t3WLUBCSh5qUFSS1wi1LjXK
nZwce+o5aA8Fej1GfkGjx7aoJw6FO35E/Bx+0dw6wVBecpuxt6how7syz9pBPJda
TVAJieQXD6jGI227kjE2qvBAYexP4FCCVR1wQkXuUqVRQWOmVXcOk8KnalXGg6Qe
vuX7IRH73F8a2zykCVv57e1qRmnJTurBZ7n5sLBCckjxUfzb2p/egteCbShCsdFU
djV6X15fRHbT8hTJXwT46f8Ic4VRU+Ap+wvQVBhCAIDZb3ZM+7JPZeGJA9WmZENe
XqjWXxoZiCgDlCJuoSRbY1a9ST8FoqocpERcqZw98boRwQ41RynR9WekHJtJZhMM
cmS68F1A70wCNdVdnUe+eZUiRBaMypLo0YtwL1Uo3NQiW8C+J8ubh00LE98LPeJU
fmHh+hnbdkyiwDwlR7XNhOsT++VHIQ5G7ueT7KyHAY7HvmFGISvyi6wZq0HfHyCc
NhVUXXFqLIeTN02lrokAz2EQST9u+7BeRmGpTBLrlKSSQBV5c7hBqCq4ldUMFUIy
fyHZWtNG6Fg+OB9gPZKRVlyyTDzgG/l7w0W0ptBoWZNFk1kSsYESE4SLyxMXgt4Y
BP3VapxXzrc8sBZXJxytIL9OLby9nRNUF+hUpba58oGwKj7FSBcr4RipEoqJchf9
flxH8f09DsKgVcSOQHgImdKLmfbZa8K18tVP1ah9WNKfuoBhqqZ3o+0qvKuDlw/V
WNl0W5iO3aBlIg6tSq8NaL6Ip35nDNJCKVvEMnaL2eVo0uzCNb2Wju3n/U7we51f
7j+4KC/ek5gzw3WzBRoIXh+oon+XzTCnfWymNVcUmLwMSADirI3IlSTonKDbo95s
Lx+iCdd40LAQVUwENNiLJHrw8/VMhDM+NF4AiF3f0KqqLLyp+tR9LJ/b7Ga2bfgN
Cw5HfmRJm9OX6NiP6navPD8GqF/NrrFeSi4D49ytQheLWeAsQeDRQMRZr5eL4Ysn
1WqTxyaUqfSU3BL75jdCw/Sb1K/7QRus+qQ8TeGnSYcjvbLrAhVKl5gs/lSCmV23
ckTWFnKixna81vBfHSgVZi7xnOoJO0OUYkFN6fMkI2X1bjf9toncVCS2Ro41ZRwv
ejRIObf08fFhy5QlQi3KwuwJ5zy4+j/Da2fr6tNHm3vjnxgDmu5SJIb2S2IlDoza
mM19AFiz1DxcuKV/eXLxMOGrZJpkxiyZLZRi1LQcumRnMr8PU0VADDi488wi82cT
jKCZ9r1S2wmr4KQLshTrlIHWfa92TnluockbePFdflPuJ0899kL9RjhHCWCSG/FX
GsE5K+zie6GOwkLK0Qc5kk/uRbRb8pBaK1SXbqu9rXZoOd76RCdVRSpFe7w04HcZ
PADAu7h+jAaJgQ1+55V4OAwhlxPh1jmuV8dq7invckSsZHL6tBHK6RA0xrh5ph84
+Z3AJz8YRE2mPSRozXryQbeLBuFP1mZNzHQ+WuQFXqvlRsqLwmFBzGU4lgxkqQHO
pE5P0VINjIIPjrpYV0TbqrzO7o0845z3BlKhhsJF7WIVMeGvWutAzFdM1NpI9Gva
ylodG8V0nnI7xS6Vqnf7e9YXXQ/Xj1H2IEpkdAYWoX7pWb/C9kw16jmovnhZ3AOa
ZTryX2pffGiSYiKv+4jKK4BydFyQhbG7eBxyQzr5RYNtWn/ITBkyBB45p7Ppkrb/
ZnLgh5/b7onlAsAheM76fEqZoPuYxiLwB9aIpUp8z+Sn92OtBTaestn6+0YxaFj6
hQ3KZ/mXJT05ZWBQtT1yssSwrfx4zcPuvCm3TX+e6ZIp8aiNStXuTMrFsWsCg+Zb
+G+mmRLsn7xyCqiFDK6EpGJREBht90wBOckTJfwex93yFqLkmnwMvoViiSW0XWHw
Brxo/JLuJNImVNjMFPZpPst3BZJOQxPdt/qMdIJJfjlCB+2+B4GN2pKqs4oDriaX
NON9v3+3gKjsufDX/iSiXftA9RZNS5ybQKda/VexvCAyZDjAHoNVbyHTwchvWziQ
G+a+WH4KktjFYwwvwofWNbxUmFB5j8YCYO9Cm9bkOLgyywoeVCq6FLZ59aSTtQiv
BkCd8Uqo/fWhVHLfPf6fG5yeEa3vyC9xoTEI547pMJDhzlCNB6vhY86uLZGu2oUe
2lK4goT8upWAeBS8502nKK7zeJz0veWFdL2LvyiuelaLOTImIQ245p+GaiEGLqkd
AIQkF71+DYgXvVDOWiuxHqtIrS2/DfZfqDs+qg9JZbEMaqtBbHAbV57DaTjvYgRd
bLcuL/ImH+f/vJGJ98d9UXRwZweZEQAjxkRYW5aj5yH+Ud9n1ta+bQUysTywfEM7
4c5Z1c4WJNr2g3PU0pjC7l9mRR1HqjwK/o0zzOj+2wSutk0g4gxQXDLLa8s7ori1
j/QByJrfJWbPZEEnfiazmUIEJtjrfmdSPv75TkmZu5NNTAuADw1LuwHcwlsrYAS4
7W1Va5uwialuvPyBa7zB+sYGqzrHi2CepezTHLQXN1O9RaM73g34g4rjzJMYNDsB
dDwk41xBs2or/EJXJdpvwFpew7gSiikRvGktOfWNNpnqE+ThYDjtTxpKyvn6Qmt/
Vj7aGwx67cQIe02eS2NhRoDG/QZyEb9+jg4DIdMHIeaWKaIlTq86KkQs9/XMUwRW
XvnZs+b3P0gQ6mhIjMoFhTggJk7qhrmy+dxvsNnS419PCKgTRr0G6uxdqZkVB0wj
BC9nbO3RLu+6laCztyEZ6qQIXnsDsaZM9YH/TPWr6s+MbMbT4EK/hD8878TJzn6z
1h8hYN8+/w1gl6yI2Bak2vC4dNqI8BnJdsBOD+WLSfb74/syrWAV+io1FSmml27O
rsWmpa/xLaO1o/aWw2Uo8vnJZYhaLAMXiP/WOaVKeloocK6SbBPhCafwxsa/TYKA
9t9kBljhuP9SfdTNSXnKsD89aucylijP5wnQ3dvRI2kg3X3AMhyzsmRYwEus/lKO
xZAI5kAnn+gKR5U4afO8T5sFe/eEHq17igX4Xi25t+kSTK3FslaArykMDHG6qQKL
axChv/mV/N2XRPeKbiUNGHhiHzjESZSSeHlSvgAjibzA71bIsVn0MeA+VF0cw+NH
pvRKpeb+TsJuQ3lF67u1jgQM/5rjFqlV9A/lgJoSyp3+GeAiAKG5YqaQ7JxwZzO4
DCfaUupwOOTFfszUBgSDCDUvuGB2QXbzlbhJMx6oVHD2aDuGcWZnlZUOmGRtWF+Z
qdnTriixiA+PoDADsBVQaXIxvEygskw10L8bMx/0tgej1ZPV/oFQnWQMmFZR0y0g
Tw7sx8rTuVg+uUASYqErVakf+vVHsdkQv1zTMLJiTLhLoDCC/ow9ibc9rrF0FA1Y
8iUNsJMMlddIrrjk+IJ92nm0lLG44VBj3S2RQ2nb/MnSWIpmi0rCiIj8vKxV7iIP
PGrQcFSBIV5XkUToaPZbdjb7rNnlHgM7et7Zen3SgisiVThqnhp5our30ePVR/94
bqQFC2+teGzUR87Tz22c1p+KTBpEtxN/D0cY20CUWBnwMQI7uOw92vTVgh9tF9kn
eaEu+UMv+nVPNUp62P7pNf8FnXTI4RzpAjirhBihgMjwzXmlOwZfdTvgA8fjMdGB
QQCiEuSGjzwrbOjUCplPVgnSvpIhevh4P/ieu+Lvh2KC8cZ3sj6/uhb6ziKNuQvM
9UZAr6xf09pypzsRmQXxi0YCqemr82/io1xB6rkXbAE3IjsienJx+RUmLEFmKz6M
2GmuTj64KbzWrIKZG7tpQ4oc1qKHP4G4IolVStEUlKB7+K+vaKha/BgMqg6U7qmO
HcSRVesgh2cFYzM/LlvNaADzHYvAp46SHVZQ9dkMhwHnFT57YGuFXTLb/CARJHY+
Fd/UXcRPIc44zf0gVKixNpHTPqJzZxv8GnfZetgEnF3GwnMKo0X3/5dt8Y2zoBWe
0INmTrtaWIi/8b6dU1aAV/DcU5toXd2V/A44wAF018tAm1P2oe/+cHp2ozaFXB0w
u/dtjBWrzEzmKEQxMjBUxeQ9wenF7p+/Rf0XILFlpr1MR4vB9UQi318+bN/2vjA3
g4AkGefi5rQwq2kpf8aXZGGWGhLmXwj2qC/YPE5iXVHvTGqAo5S/HkTlbuBoWAVf
fkbhS4QOI1IZlGTudthw3XOxiDdoHgI6x4+MQMfSkRTZcPW0OpoDmA7BDbv4p+bP
Dtwm+lcp6HH3aujXvxGgUNF9koAyKiI54jVTkIixbj/+YC5E5xO6kb+9Eo2q1qDP
zyBdQO3U9vau7Tv71qmjqgRjm41mSPKHASCr1v1lzXh5u6OxMEmvEJtXqnMJ42NJ
D/4rc3cUPQFboxbHrmc+Z5lQ6FD61kTjILEU0OUkKT30FMPrph2druEr7II/4Ogg
MGC885d84PXPGQhuzz81gXHKyfyLjZc2laNbBuZ5bCVlyhPIm8mOez788yRpkoVt
OFUwgZBrWZ3a+pzJkG6LlsJYZ+wxk0ct9qitIZ45Jp7owfwyMcVuw81iYH26sEPf
vGcHbXdC0VhDG8yW7zYnBwAOMloOQadBWDYeAuK3xhctNA3gk3covRX6HwgKE3Kc
GLGVUWohbNg430dCsTIC7sulpqCAeEF2eexl1k5GHg/Q0IPi7eCLOpt6phW4GDZ1
UxYbLuj+BhJbeAiqx5yZ5QLwfFGBxVpxy7YMJAcDiqCL/TmDZJtqmjLNkLaTIudg
qeMn5PAbg7n+qI1DLt8rb8rPHLXMgowhLsnYN92xmjXkGIfAH4jA17LsbWsWm7x4
vdLPJQC3vEIQPjvgMO6BKIIp9tWpzT4F6FjD5mtwbGWmGHdxExWEGoFVWYDJ4VZU
TtjrI6azEf8bJeIcJHrGEkwMgPgoK0gy6y0AjbABk5zftiAYvTSNGFehP/7ihJNv
jlwxFax/3hAXBwdFgbFG3hh0okpyhV8bKEVSNsXQCCStCr1/4XqiL4w8mQ5fKYOC
6VkPxVqGCPkBBXOwLwQDUsVRJoQJBS1H4AmuLc4c/PUkXaA3bnNkgbC8XlK8ATLx
0RGwWtlPdte4XjwdDRg5P4rEj83hQch6j7JUPBCXW42TJHQOA+VW3GiURBlSz1uz
bCnRT3Df+1Q3o338AjcWwy7v+8TViHa4aQuETRdjQ9LKYn0PcYMda0gU7g79kbZT
1FK/6qKGJGHHZUDACpO/Y84ssVJdhnxaVf+UdI56tU2B7R3ztUbcBPUAP2QHHi+R
l5Vw1/hEmRdBwY6rs1l+KaOzrEDfis5Y/2EmlojZ8ZKuqBd9XE3OZqdoPr5z6qeq
N6wgQ5o113IyN5dwi47G7n1EmT7mFJJLNPEBww1fb8+JzZMUtH9zsSlErZbBj9Ws
GFGLNOttitewbTf3a/1z42Y0Joyn7IQI2KCOSCAaPDO7RLyXaNSt+c4mgOQgCWO1
WdtsKqQcqJhNWS23NL6FLSw+1AeWQwCyJyObcA7bmt8o2v9mO7JdzptfrVmV0AyF
yjL2BxnQR8orgf7vMakJj29I0H1L28zQDkx8rgnWD4s2wTNu/mKaD+I7mDHRDgap
IRQGs7VBUV6CGrvjyeqFNJFxmcKC4o1POU8rBah6W6neti1mD7WxOBoWtERrqfBc
bGUBIjY+jRoyu+wdduE/yNPOqDb8ZtNZvPhEQOAUj1w0fDUrYoxRTKd7JyVUxsFK
gj8vTu9ENp3SiTMgivJPdb7yEGxH82QJZmhEnQrcFwJ9QNJCIHbls7MCebixdSA+
TQNTDznngyG872R1w4zZJOScgNEQ+1I2PlDs+bn+MIroCPhdsZqdnk6AVDHWdRhD
60gJM3wGn8DV/E/HBieuNMsi4mLnIv4ayT3Gejgp+WuDxVnmtU6kVJ8WYUjhzPLM
Jw1FCgWXJJg/uUZgWDev3uxwQ3Eeg3NTTtifbM5ltxY91NWNvejU0TMCq8fA7KCn
pGJcmmqzNs6uGpT2CvR2CCGFV5Z7j+RDYoZXxy1UEuUlV4ohuUqTwD3nSzcqFURo
9t9K5UKpZP75PwQWqjwBrkgHgD7Izph2szUvBmlM1Lvg/9xQKdEfPxI8KzCq3GvD
NENarafEkDuhxKAn0w/xaPMdEWc2UXv+Luw+TXGx+WeCVxt0sNL9QQCxx7iCPgEm
jOcyL0nMLbLDIiWyO3G2cNAM7uJAki3uKmbcNiZAPKdqvFRUgnzcSMgrRdUmR0PC
PJZC2fnmp7fb30PIKjPxFnUAaWdgcI5A0MQrkaSu8L2VDQvx+Ok3cueECqgtg0dq
5ALxF4d7KDckfwrU5ywJfPou1Y8qoQGHYf6BqCb9o5paq3BCvxHokVgC5kIGKAJ4
/v70sZIViPx+92HoZbwGV6IkaACerlfjQUUmPFJ4x0gGYLlva1jGyPy4BSxCKgR3
IEGSkSSYPQJnVQPpUaZm8/Gv8gU9J2NRa/cnEr12FfsDEjeY3tsAOVW8f3lg9h03
HEzR4WMn/ewqkGCJFxYf3B9XaoYzFKGqs8syQ9zGSsSISvjz4BhhvxxOFEYjVie/
AYi2CSfOcnna8Xdr5KNYHefqE8vdDfx6vlIBrRqnVBqiYO/HSn+bexoIKc2OXpAj
EZXM2Ira8Sp40+cqG8JBaGpkf6nv2zHe+SybTjMyydDrv2QJOtYgPk5Zxc/PNfG7
wP1q9C+ygyq9Fl+rwNNDqn/KP89cX6BEGkK4DyclELx4A7F+GtuQ6xZTiQzao1RT
lEJlHz4qUm67aQ+LIwfv6016S2g/vbmlWZ1BPoj2YM1FC3VyyBr3YdWyVvyGcqol
gpHjWQs09NUJFSQzQZWy9KkYt0wFNia7xOceq93CmqAjyXI4wpPPuyWNi9uz8g0s
fbSj1omENoDJpxDgHGpi+7V+mH+Q+kEme4OEc3CxkJ8Wpf48FZ8bEn61B65s+Kzu
VFdwMn0vPYh5ye0FuzOQCnzmcmWXQbr5OJ1g74irWDwyxe5gM4EggupQTMyTx4yh
ivpinT92vMZZgthroQxbckWG5og/lznx3DfjIn436d0LST/JJHJs/HdFnYNq/T2r
Nz1cuWWWs2KlX3E5hGaFagwPEv+C4GpOcei/pvQQ5Wc0BNv838/ttNMOKtFiYeo0
5O3B7mSFzxdTlxu7TQWoQWlR2FXXIDyL8uhyaG1vmbv/Vu/b5jvTd/2Twf0I3diC
iwO/fTAkSEX7pPAiwK8pRCA/H9d5gw6rr1yiKuzsEcLiJuHwByytMTxHYZj8S/aV
KD36bBL2/qeCEgTudJPhvPebuWKcUZq4qfdBIMHUEFDpdkMGPuf/47vENlemUG1f
T284jSxaJZfC2wHidGkFeG1i4zicM9SAVNM6OGvjYWv/TIQcudpAViutMdtWE1wJ
QzQ8Z2VRk0ZNE6PzN2oqj+NN6Awgtij0A6g9myH3VKN5Zvw6RQY2POhRn1Qsd9i8
TG+jXXFAvOCz6LJAikkohBPOVEMqCo59kNzvExdvSj8tQ3HN+54U6o7quTFs48WP
rlcH+zbo8zbUfQWlgkp0nwa3zjcJo/9qUXdi4CrBQmrBeMAuOO7yU7WKPMwYhZX2
I8VcvHAl2q92kirBV1BkqiVf4/zd6iI6BxcLA76Oyxce3/FYKzFlVezFXHTF02Bd
M1ED75Lyz/bHok7/MRrOXm/yTELiwcVG6RJvTLe4Vas1TCKkvcCBePjrhyP83wCF
1kdA6QgeqGTIwPR5k8yB1lrJVFnc5CGMEF7YE722iHASZ3onIEiIXQyNPSUzguIN
gZmpwl5o5g8tN/R3dLnvjwOHLN2/1SMZYs7lqYUgC+gMyBaftuvzAifU2jhrbh2g
qedmYI8y2BcTlvofGYxeZ4KAdBRqHQZaNLgC1MwjbDZXc6fzQfXVcJGkIS96B/zz
Yope/RamYUw4Ke9wtII9Hbctrkb1vzdeP2EHzPQJqQWJz0WRU8uSyQWmSlIqCfGi
Bj4zEok0YkYogW/gaDTIymyZNghYoOYqm9LBTkQaVngUtoXLgTbgOxoFnQhyOihl
4wlgrYRLXcccU+06jZz+hMRuG5QP4YuLWDG1LWIhDasLFITFk7PxpFdEo6uVAX5G
1lD3XdYjmiJmi7bvDgrjNzyPf9g+ULkUo1rU4bcH7emFB7pl/R4qXJ9XZ2ki7CAV
jzhV9t/o2gZUn2g7t/qXlLZqW102aC1EVAxDGnPQf8sfZkugA7UZ0QGfNHB0/rdu
u/e9H6WcNBHPuYXmEL7Kd8asYD/jttfv2s97XchMzmCKNCZO156Cy8J8rXFcxWAy
OH+K29ZUhjUBAcrmJJy++sW9OUNWfBIxnBU6lCXFiOvj66N39wh6j/PxRm9N8bUw
be/b6gR+ccly8icYYFWIOET6ruj2zYWVDuynDIeiHxxiEgOK+yBCMKBelvL7i0tj
lPeHbcOgNpVsSmLcyAQBn+RqRqk096M/brjMBtPuaPgRWcFXAsduUG68fQ2eZ4zz
VSqMNYjVRovJwNqHSfvk9rea3D59zaIWusyC3OJteFJmSXnYISphoR8o89YUkayS
qoDc0OsRBONrXeXV6tjvT0aQj1Eizi2EWrogyFkltWbVjwXnF+cPy/3T/0DktbZm
43M1ld2hRAl3+XBFSNmcxDxusyZpY2XO+cgUZatO3movkbPfnkPRgIUTzcO6FW+f
B+JtvKhl/mtZRwTg6+6tqS1Gu6HsB9EIJl5X3+N39RfVCUOvpFUV4SnSVusBq6RS
TcGQNby3o7vAg4vtTxy7fdHLQ7H8HHk4a8520uPsSluQYDVsDs94k8pZn4eVUOqh
9zGF2bVakrjfHC12U5T7qevShPrTpnJ5HTeTMDbE+43wo8c8aL2f66qwGXshIo6b
PugFcapvcwdEvDi6Jm8AYwDqlNrdsyv9f9ky3FDqOhu61590PhQwfQoHI4c0GZOX
4/jHa7r5R9UneOwIrioUjrX6Y7wWbxoLNWJ1pdoqzXx8IWvCUgfANV3whWQ5Lmn1
7eROnJ5A6albRYCpzJcR4lQ3de3/uQKeAmYv3TBz+ssSViVKK8lQr8aRvHDDcjGM
MqQK/YJflGh1zzXkT/0SemhCAEx+TPx1j7dubMIt/1rGxu2CRDcK6xTRw9FdJHv5
lS8GMZ9kcLFTNk8fHwQrRIbgx6gM46mF41kRix2svxM6/X1cJ5UO/hkSFXt6bNqS
FKjArIYDeJbJ2p4xLa2JQg1SYygvOMhvyZXDlDk/vYKGxQinMDA6h/0ftOTfsuVc
nkvaCLWBkqLiPzT1Wv5NNDR+hFC04v1YKf/ZHkRZogxQvbQbTiEyZXHpVQY4PtOW
z4tvjK/SOtX6onpxr71Z9eCdOkUuq6qVhcCYZAFQiFMqvV1ve2U92St3pAEJtWYD
xztFZ2Ls5oxn+b/lVp0mVgF9uAwXbMdwXRrW4MTk92Okc7Dbos2/1F1aAI97R3FP
IzxEIq+jYLHaBuwrZsPhcOee/raunVXW+VXACVeBnzrvSKQ0g40nFJZpareEb5Ww
UA3CPQhfdMw09ZFs/p/DxZ3DMJIN7OenR8kV9VobJlpLZWw/kHvp3ZXizG+OUK2Z
dPolA76ya/Kaf3BjSyoIznQUQ4sbeCC44cXZTCpd7rtM7y9P8cE7hBypeNnBjWiT
kLxMmrOcn5240rxCc5tgEWWDu+8bTHnaZ6xPHGoL+xUSED/40ylQHPMTtN5uK8K0
3YkuKzecTBmHPz+hr0CeELWHxBWtYr/LChejwHN1vbeUlQxJDcQVvtLrOsPEfpGH
sACoVV9UQV4ubGjkIH/EhsQOEMy2zFAVvv2+PjnEWap/hD3nt/v/gLB0FASX973E
V1NatOlECtlT382jVXiK4zcOR/frJoUZIZ+LH9N75T8LdN54AMkDl4WJHCQ/Xj3p
e9rmMr18doc44DlXvW9st9/ivammJYN49SVa+/sFKicsLiTS6uUAQvCf4a3GEkHj
2j/NVPiI+llNdTNCrIjXZvcnX73Zc2p12oj87vBc8J4fDHDd8NdcXCQGobmXFYaD
EZCjO9+xcuEAjAZ83PmKkD6Ip8VbeIadMG4HkuUTFurUuvDwDPgLmcjdLYI/htZG
I7FlHFhrnzOA8v6G4Fy39JKosxsspOodbPTBViCDTXHbZ56O/ZpwNxHphh1+c1Gm
TIV+i65WZ5ibTJPWIUYdENweisbkSnpFH0YcFZWFz58MIsOwvhvroa1UnJLq1JLq
O0Kj2PccQczEuhV9BdBqF6SbMNNShe09u4bngzTXESk+sdNhgyzQc6W6e/wq1pD7
V71QP4hVy5McAPxrDWLP7VUCyERYc4dytMZf2vgnhpXDcf/MpLcR/iaQlc4aa6C0
bO/8C0k1qXRip2m2mx/2zbofPBbSmGB19ULoUtH6oyGTFPNKZ3W4TlZ3+K+g1OTk
X2gxFomw9fQhB8xl7n0JMUl37ymw06DfFQT+0L5YHI6wNNXwQtvagTygicRr34VG
O/3gMCgcozZkBrPrt3VrF0i0X13XgdQxgzr5Dz5SHQ67B7GrwPuTfbZEhIOgsnqk
GW/xJERlM+38vv8XiMaAI/NAqcB0UFlpX8OVQTIHU6ltNPyZBTqNYSAMq5l/HK/H
l3LfdaGjuMzxXNfwWSnHR9vzT1RjGOxGDEMHSbNwJgNvuqzSmEWghi7DCH/gRHAd
mc3tDw999WYWTaL18fKwSnwOeH0kBV17ur+MdQbMYEaJztiU6fmwgTP70qC6jmyz
37gjLQmdVOGI1PYGJVgrEVHKKbyZ8HjiA/dWV9v6tj7rEmz357kWL1TxwMkimvOr
Wp5sH4qkQgQ7jNoZOX+HaFqMe3ABjQ69jh5oJpdGU9AEQAXYS0FgtNeQkJVa9Mx4
tM6PWyPQNnMReFT47YNrLIrNRAklwwcVvkaP8qvkCyf4y/WLWFmnxxuRIOU4EjLu
Y6/fXigBRtUoLLC2M4LeoluMZd1HEmTdvBd0RICcRzUWRFR5B4kYO7Rb2B6FiYnr
Fe0+xcOCe2Svk9yOs2y72RB3wmODEW8dM1gbSC5wkLytyKCQleLOX0j8lKVlRSCM
zBXtGQnzCOeqHpdni5eJVS3zCiAVIpijInnCJL2Ggr7gvGmE7BOFO3OxaluYT20B
RaomLfPu7nuJUNaSqb4MkAapddVi7+oKJBOCs0uNjc6XjYqd1dasZE8snav9pfue
/AFR0eiSECHMQOLR4q8vptX3bM0HOv0V4WwVheyrbIr8BTV9NI2QO5RGS2JYRs3Q
++BqvqLkRBUpK/AkDtGR/ANCQZBoKb50CYw85etF89pYjvSp2g6dNR3eHLhPxz/n
JR5+ZlA7JsE888nbSqx6ty2H9K/ysBLYwBtcPUX4+/kkEV43yT3IvpMdfWIo3Ak4
KaXLvojGQ8pLeBL4Toq3wLZnMHD+GAWZ6gCrdwlc3Ab8PnmdJqzqc144zA54QO2s
DYMVcuCQqr5jfBZNSNiyS7XiaO9154vQaOHqoik/VVvyWMjhG9o2fFmnMxPtM21n
+dEUX1LW5gNm9Ki2dtiumS2PxB31MleS9QXsd3QOAOJRTMth5n03ljYX8j+rFop7
KJZgt077+QYjhJP1NsH8aIU6BWXcWamqeRr/9DFNbD1Ef3fvuIEQYsUMGxohLRi9
Imk6sGEOAIl2e0ZKifAAj/WWXVq4Inp/kLTVTaCqIcCN9tIxLNnlG6WH+YSjncZ5
PZoBMOPEYpk1xihp9Zxax+d371BfgesljGZxroCn/Lmzxu6mnuhljajqOKfJZk78
J7HMtbrVNfkOrVp4uP5BqVW+9rHDaSsG9+E7z63kMwo3q7XQmXtE/yqOGrg4IipU
Et0M5PO4drbie52Gl5eqIFAP8AUYJnoud0sADEjQNO4pnjLkGm0z/t2nIsweUNF+
nKzklCQzS8t9hdWbLDVXX2mWe6mBd+iinhgeJh3EeXbTXzi0aO+va06DoET+k/vx
6GntfzuQO7Upl1EyHfFWalGkbiuoGcU0juPcWZPbKF6yzAzFRry2E0GA/Io+0y2C
ZVeRB+7332TClktGbyaNFwtIPjjW4HUrlSp34M3YA1kNWog7qcAqP7RXsi0mqK4j
q2j/J9vUjAuGJwk5nFwKHsHoMbSfLmRAX4dcuoGZ1uKmpe1/P/ni9zi+s4w9ope3
ToCK7MJrNerenptu0OulB1PyAPfkKIH5naIVwxLdIMIXvnr6gebvVDmRZTADkX4A
7tP1IFv+Pava1LPRI6kQiGF5aj6B6Bv18YcnzZBN/dOCGJ0HemS054fLI4KmCkzD
3/kSkTMrozt3reLPFQYJtZnNAsx+EJ6r4c/UK9VshDcogUcshFBeb+P9iS3DaagG
MAomekFFL2hvRzi59gwUXkMjIw1nLfOIyHmoBzWiSDo3IEcL5Qkd3P6V8cODkNtG
XiQYQAjh88w8xur6RFJgOPOOYQPTNaJuO1dFweud/RMDGdzswgnS+DmZrBwWbNNN
WLXvQbIym0FUMcIZAmxVMbc1tpaSKs9PJ38m93q7pcTvDkUmsAuNfUzBlzEDOvE0
H7vWW8LtuOL3Jakw/ZQ3JCbEVasypxUc98ZiJWYqTgGzXX+iA0xjKkN8+XOIMxYA
vYcVpN8TakPt82R3qIezjXS2ou4RdbSEvuXYiZR73j8JnIadN37V695l7JrCSWlN
ODrDdpaGBQmqC7QHTnHfs8KWhnNqu41TA2Dkff9iT6agmzznv4yvS3rhS1GLCf6G
RziXlf3K6qSOnpZyp0WfO/OL1XYgYAelZS9kkftqFrccrfjO8EGc5Xh99x7slolj
V0O7jobIIGoG+yTwfPCw4KPIrPk/DBNI4tyef4e1Riq1MTL1mNghQzdY7oncBmvU
yrN+fLGqQlhTLqWLMCc6CK0YOa6DaqFxtvCNMS9ofVMAaLllUf8StyufU9ozAerv
kYUyzgaQ/b9+wRcNp6FrK6hizuwF4QPDs7pzXK/Q4wj3D7zlcec3d2/WpTwqXSrd
3tEkS2bBulGWvtLtU2Z/q6+0g7xAis1zDReiCmRpY9XdqOskY8900CyXfoexmj0O
obolJ4/X70f49+tqoR0emIZsG3PC02xERWAHKHmXWWrxPr9n9A9a/OAwMT21Iera
ymX8QVY/OPW7k1JDhEIem2pdWziMsHP+2SdMoT+mzM4L7vD3TKTZmNnAuDHFOa/b
lD2PrFm/3oPbf1j0X5rFBZaRj4ZngtMFVStV0+Fnt/9B1Ro+BlilyTmi2E1vrm8r
iakyK5Cjasq6STvfXj5dpQOuBPbovSYyhYen+WRiCBYfO5n3k6ZtfLD57OqVdvSj
790hvzKHhdkArLVQAo8S/dvYGGZF6q6awFzsy/ZMM1TgSRDSz+GnNRlLH59Reb/3
l2vh1OS7TAre0GdW49XS8v7ymwul4/fNH2ogQKcy+nmQ5flELuH6GeZQFy8AoVE0
phEsj/Hefhex3bRq65EQ5hmR/Fk05d/52A6rCI/RmTQQC9k5hnEopeN1SJD5qCym
aE84DNieqeK+xApKBHrvqAb3pxD0flm/7umwVYwVqV943IyG2FWCwHEMvmi9YZYN
gF614bGAJEVO94xHbylfWcYrk/XOxfPJP9daGhVCYV3ZYTYZCKwWUSfPzLa8PeLg
FpSIG0/vKNMMTC36kEQbUlV/+D40lEh6Umrbs697OANB9/CiAD5omm596Z1IYB/R
WxjAAaOIHqq9X4y9YRbW5Ol15h92uLH0bUursiHTff5RNyki+l5YZ7uO3U8xt8W4
Y/vnkAXtQmeH5x9AhAjOg9/JvkZtb0n6AIpCo0mqHruk6dWummzcI+xnPRSToz1T
mFxrZgcU0K3dUfVRXPImmycz8UBEPVlPYNgM/EtAuzGr3mPFahgalpAbcqHE6oGX
k6zrIOGtB3nO8hba2u1wd4t+zcpYajwU4GYHuviM0ozOWSut1fvOOR07oTYvQPFm
z3pAbWVly5XYDc1BF03kD5cRPspWAiuybE1oPtwrzO4iXA5Fos1w91oAmQTZlRrV
es+Zf8zXL5a1adwCLoFqVrHUzr/Hp4qsJbja4gUtvub4EUKU420bSzXz4rl6DT7d
k3n9NB90iiYTBFCJBhmG9CxSNWk3CSPOfTTsTVeNIWhNk1zm/uBOAUG16U2i/nwY
YYNoKJwE0891nrQu/+BxDZknaGdAij1xmoYZB26inzAXZk2EHuMoiKm9y7m9+kNl
b0cjCfIg4QSiOCBA+yvMvNPBDaii0trzZVsr01Xsl4ipAtIIi62OCd7tv2nzvHE4
eXmen1EZkYBf5rrpiqulNp+PkLAeZWmX2i1CUi9esYzUerBm9eJyNjCfN/a35W/G
24GrfDuoVEoRNobC25t+LQsGdtolJ4zEfO52TZpCUUQqBzmtPM/uuiahFtR+FCZk
/bV/BbzcgRwvkOTNedhDNmiD0o04qgYZt4Uz5RvrGgWz0IzWLoFkbQRirNYeJLg1
rYXOcBh+AypXtPVyE2ihpyD/1RDovYiFKKNRZ+TRXa3pWle+W9AAUK2et/ct0mj5
hSfMO9rh9HxuEi7HN6XbIj5liqgBdyZVIxjaeBKOQpIfImnJQ8luL3b1chD5F8da
HavERUI9v/0lAcpQuXW9CnoO1/aTBsoUJ2Z5H7q4eY/rlWFCBkua63tNOW3NRjBJ
jAAlq/ypENunqMgpmOdyc8dqxqGsZpTk/KjBGiVzZWSjzfCnMsG3trTi3iUgHdIj
rgRUhUDtQXKEElO+l6pZ3PwHHCIYhOaFfS2np4al6QSdQL1PSDw/ZqyS2tu6mEMa
T+2J6HC9F7zUg+KO1WBHAiXNrfZXeJZb9Xq9qcFxdPIlqQIKLWViQEjpcIntqxG+
RFArfVMeixsGRGaE5ViTknieVJb0Rywu8/yr6VrPV8vUfigEYxduQ4PA2MkifuOH
XP56dQ+sb99IzEhPTMbNovLYs/TyTTnQ7Mxe3gnhfqW7VyS9nVZj2/qOtxVgUNRM
6ysyMctwM0hvtZjTSsT4BedXyX6z04aHEkMrdADXZt9VAhd+7QXLiVtfzNMF6SpH
3lB9QyBp1Ew5uOgFgvYfYRJ5cHa8vOGWB5rHbxWMX9wmpVrhayvwV4nMYVTjprKn
72pA2ONRhyhZtG840EqcJAA9EunIX/mubwoYWALJ88HCLmPnhcc+PN3jntD8YQMx
x3lIZyCZdwD4a3npVR+ws2bWfLpip2Li2I+oATzB6ukJYS9fH09wLs+sbnMjpTQL
rjeocXq65LT+k5Q2X+PsczW2DpE3IA6n5tOwTqbLbEOK0uX6Pk2zx1JWIYPCY2uR
Sn+1bsJtirLCwuhFdRtpy1gFaUpMMYtcO0m2NwY2IaS7cwGLc377BxaDt/YubAiW
nm//LqCFamtiXNofZQM7588alOED9vqTyt/DQ12eAkOWlu4IG4XGw2Sr4zwF++Sw
DQDYxfYly4h/aSAyvz7uX+aImJb02AHG94fMM7AYIV6J+um+XvmbZ8VIkGz1Ko41
mxx5G52AiaTMOj2izE+UFijvjtZxJOn7l692HzGePq5tNdkGdWyiRPIP+qZlWwM/
Twi+mTm/+6vHriicoatKNC3At97BaIze2y9Foft6d2DaroEb6ZvKgo+Yny1+7W0w
u41lGZ6jzwc8zu8LcpEDje+x1qOlroMgLtss5/e1r0XZ8x90FAzh9KDhmGNSlagn
w+hC1/Ki8ADBknA6v98QlC4BqNA91L+Ky7RzGuFBpt90CZ4a0vb1vgxwpTHARE1C
njWzsmojOZzzE9BidSl7lLch6Ix/48Hn0bM+QsWvUCVDFTbBII9HDkuZpPOeBeXv
ePjXjrzgmtIW7Jcw1s2Lf99CW8xvP5CP13SPCeecMWu7Mqe7N+yEgBnN7ActsDRW
xIomg0QbqMve1AGFRCf0tQsU9IGh/OV1WhpfgZYRtFpXueBUwIl7++5fvzXXE/hk
quTK8617gNhupGlB23tyx593UzrR3j8VKH8TRwiUPKD7zh/ndBFo+7ykuv/VFmzy
tTXSy9VaTHoxK3CWLgTObOg+DREdu7F3/P/T8c5b11QoKK6XJztTnkJmmJ3TmrtI
WuLMZ4qpNQVZQqWc9biidreEWn0ADPKEgoKS95ggahHh/JMF1Z4bPKXB4akL615R
1tA72sWrj5qR7i8kG2anqGfQ/ab+QNa3Io1GD2N62N8gBMKlWtNUUu8BP8hGH0kJ
R7GcZAQpIZVL9bMCoMncjAZtv8UTXDSq0bbyTGq8gC2RqNTN51rTVc/yAJ8i7rq2
2r5IG9ZaIfUQ19bZ8gpQFipsYH4+4d3iD7aOnYeZn7obmqHupQ83W8imbbt82GS/
31OOL/2z/FsXHW3W65qsvSEOoQ9z84KcAPK99c1pYM1T68Ed8op4X0mq1f4FzXku
ujzeFNaLyD6Nkm6WbzF2CThluuCbH+wokcizRkc/r6Ny1NiKV6wnYh/dALGvu1MB
2UQUvMDvvqOAE4uGKZfai7lhMMlRSdeIHblEimP9J58GsWgeKUc+QC2T6OUyM9Iu
bEmYWMvO26aPykBLveC9fyPgyX07rbNxOdYu7EMV0KQJB3OocSJiTRSnm0L7AET+
Fd4P3yAwNFtHMV9VOqN3MpDjc7APX8I91l6AW8vkq0oxl4QWDuVB8xpV7kW8SRXY
iekJi6/HPZjXDVjw9cPjV3yAto0MVjYWNITni1p81oKtMhHM9ArdWhoGL3MRDn9F
o+ez07WTvbg+sAcUM2wmPuEt9Xge4WIwWryTw9K7AttRhLPfcp6cgGq0sKNjkSim
juATlFoqsHb0N5jD9HgxisT3YRfHwKJPhjqaW1DgmKAXNvTP3c7W6LNVeKprBXWZ
r2/9J0MxaE/A+Yn65duitKQfK3ePIL5iFpJ40yfTQr3lgqNKIaEkRnit/xJgEaU7
5pwDMYa/tHx92hyj391DKuTxKO/aekdwNBBX65GzjjKCfKNCJZ8Duc+J3v96Ue3+
CSllruJ0kith09a4VNWcdSejzKIAb0UXTIMVaDij2UkTkgp1xAWJtHLRUcrq6SLf
IQq5h3CkBMtyrcotoAokk+YApNHDPJuj817AqafS1cvYCM7+jhNSZdesdLSOKRWr
rAV+UCwYyDUEq/JsBtHhHceiJ3NbK5+n+eImN/ad+axUtQ0k/PGOmYkWW8AAN8dH
9aYUu5B3Eu9olH8mChTNdvLeq/S15HccH79LsAZRCnfFDepqA1EyMwkZf9UPwFqN
xmz0Pqfr6guZUpMg0arZBJA1lPY5FbUiYfStmDt+hMbZrPZ4VdOU8Q4Gomlw1mMh
iloJDinKke69SC80aXSoVd2BETNgpj6LQYHaNb8qENviOb/cwx2HZ3Wz733OX+VN
frfT9v6rWxIHO0twJEevtpd3b4BNkKM33fja+yNXPPd/KDGNajMsrsqoMTBYdFEN
gh8knIfkupNye+RTIwEurcV1ncnuaSLdxqBEHaKs9pzQP4tv1rR1PY9exx7QJpHC
LadhMpOvcbGpyq1lp+mx8PQdXHzE2Ebe9Ud9UIojGfNFuDbKBw+S35pTjDiJ151q
AiYB3ST1yzne4txWdDmGnwSjCnHUoa4Qo6lXgXrm787AejQ5ODtA9LULPHfOBcyU
aHWjyjOB6yoXF0+viH1OoGG4Q1NPLeJK5OtrvB9DeWlFVmKmQjTx5hECFC79Opaj
gNVgGbt3xA+9NpbgkmDuLmU5BAoH824eJXLVzLb00bdPUeyZ2MAiTHNEO7F5+GzG
IEIxpB64DWO27KmzIG3cxR+syDneb22cDgdLaRNBXtogiSi4KL9d/DPD/PTwmYBr
gw1sMyReLYYmJoOU0L5sVfKDjCGz9QccjTmjkdWlNpxP1f/X/ig4zJHjP8linKOa
mM3w16G/8Dztqg4W7SC2PldRHVEpydgVg1TvjaDmO/vbo8UFLIgQGfYYV0KP8yRI
5H8TcQY8ciMHeXS6G3rvyocQTjeD4i8nbL25vtZIQMLGeYzU7ld8k2cAvbkvgjvK
tTgrNAxcImLkZ7P0DF8S+/pVG+rN9+kL8PVL3vtvpeta6z9wNJl9HzYx5oy8Ho9O
yG09/zdw9ozzrNGqGgnFD390d9bIqnh/xFy/0qJDuFgjaVRhgV7SDJ8mmIxMPfA6
snPo8zTj/zXvHlVAN6H2RdgJwlAKR1hYwUHDdIfsJYmzMcyFfsaXA86HwcfbzBJn
hUihpKyJ6i6OgnSMdzS/9s30eqlxzjWW30mGdH58h/zUplMUZ1SH6yoBL3lybHfc
CGcog+qzLknyJLiMwWmJQiBOppTrO4HxiufrzLOZK076VscOedkuxsUoTFdO6cEk
m1+TuztXk2AbNHaHrH6RDSQqOqs0nhg/jjFFfg3XcDsEZYZHLUmOTdzQXsGwCmLW
CkkbXsL8D+DNtFy4OX8kamXERNcp4P/IceMmtA+n2So0bPPTcY1C9n+tqN3/1i0x
IO1EzT+8tdCGWREt7Fwwra57EfIBb0jfPu2Kq71xoBPbUeJsSxOx7hwIRz+Kwfwm
RsThQA28+3rPq9Aj0bsBykWEvtbsbojqKOCHEvHvVseDpBej1AlQE+34zV1pSAwH
NT3vO0hyh0J+nzPxXAIMfwjJ0PdVFFbXtsvLUqldOTyd6SFof0nySWLZUk1Nbf9o
dd/pL9trSmnu/Fc1uWXdlqYh++rfn5ofLWktw4p7SzApQstRjb3J+Vx7+FzHRv0J
znT4/5csXdRqxa9Mz5lZEWQZLuja/34Yb7U1PuKapK7+ZdEIk48jo2/zGPfkN7PY
f7LPPnJ03i/AN18k3fPnlx5KvacmjrkRXPYz4DA8R/BwvYlWErRpTu3xZ+oVGlbb
xKy/fMat5fCoVEE3+bsfAiaXhyxzgnLpUnz6S+icymUuouzgjZbazWddmS1HWj67
7ltJwoHZw6xKI42LYiwXkYPkHyBNj2atJqJFS9L6WxfLVxz56sE8lhbkk9FmjdPS
Qet7d7gGpKuMAEoJXOqbDYkqU5/zwUBXl7OGiCxTiDmOz7PXR2NAZCfKehT5bzU2
+9uR3zyEIXS3nmfjjyusSymMHmlF72KRfQ15r9AO3ku4HLiewyvJ4xALZ2I3qXcQ
/avJvxT1NB2revLmq4UpMf/9gmRXP4qw+0HSFxDarOfB/eG6Kay+nHJueJ24j5eA
Lfd8w9b5SykMj+vU3y7stn1fQtK/Ipbi0v+Vj2oF1+LXe99MALBOgv70sJPb9CgV
gnY3HeyPwXOMIiAhBVKMHi3r5f40ZVfCTJmVhlkyG/DmoWJnKn82muPggbJ2qsPS
PkFC+uEsjNJvlb7VSkPuYA5JTWfsoBZgY5W9mgqA1VT4PLaiIgXqSAqHsOFiIWNZ
lOc1qJi/c5oVDNLz6+yVYIsNh2R8EvfFZeIo+iYgjMpGnaDlenVXxbkf2zcnuEHB
XaYeynW7XEUvtYDFM3rJ/OCjFMlOwwKltHRolNhZWBrrP/wpQODWLVTjBkeAU6t7
px6MeJa3CyfwqmEYdg2xZaFc/u9hWOZ84UVkgVo+/XRqej295WmwsfmHcNecYr9T
VOxnug3AFxX2RhxHaMQJ41RyVkt25nOv1dVPJtLGiqKXNSBqTO2EozDzXy0BWKmT
Dww43U8ev3dy8J9igYh2bsabHtWTlaDAxAKdrFVA7ZWt2532PbsryAkysXJU/HWN
ZpY/6DjNibLx38ZXcvxSawIYm9LXx8lB1bVgCHwL6KZjSMA9oViZTG8WyvFpCaAM
QrLPUmax/Ovk9cvOksWhmvJlSD0ZdLstdyqzSZH7bNP0WP+6xsVTp2VmBJRUhOTT
lbkor9FPZJApRaF7VuXwlBWXrzPVGOFv3F8V3g7mWmGIt23tRJra5e3yhrIYYyje
7se1r54khhqkgobpw978BvShdaSMR6MShaEQLStZQlGV+ylYVX/EwyfYRRzgin7N
A4NJ3ZiU4hN9glRoll/xgn3L3RmGmhJLkIqT7+skMg1wQRdpWmyfodMJe1xP+RB0
yjF9fi4LzN2zbQiownp2sbQCrCpydlB2YYpWOdktmr8GlE07atipVSs2ePwCijVR
GPdkLwXJLZhShKysEj6ANcON5/+rXssNvwqZG++s9/zd7afZUcANsEG936kbLjAY
TehYMQU1/4G4rEbFZdNe3pcZk6JNM+jf1nm/inQqAerHPtxlPAIK8EMb4tYZ0zi/
vW+qQumKDDr8vOkFAlX6AdHGehI9Hnvt6wVUAZ1PLJoGUXXsC00Hh8/sceBZ7bDO
7JAlKWsDbWOpgoJTDR1rteQ8Dq2RxYiBRXWh8JYMuC8jTkBkkHyHrbF0v+t5ZqR7
UFW4ecuWiGVKUrT2p9Ytoy/kPov3G0QvSMrx/r8wVLeUkgCGVpr1bx7L1d4kXKBW
EqbZsKYtCLeWdPbP8kmUo7R1SuyxKaj0XYmlrHdHB1+QfEmsHs++npXqA7ajgnv2
bqx6ENjtALno8o4sIRe2eA82x8X1nkNH1Go+6fv8IV4fPYqBdlWXGx/OiHBp4oQ3
2WFkKO7N++O9iSSHMQSbW9xOEcsSUcyr1iyqwR1maUitEdhBv3z2ufESe3aRj/hQ
yqesXMHjSL/4iD3nfRuOgoHbUhV4JxQFmcx2PrBj0ox7ZRtsmt5jqjoAg8a/ZZP/
uDoo/tIrH4tc8wZ3ntJyVR+A8qRNu8siz1eU9Vc3hfFZEdcVer1hPeXr67vtjFbG
I3fxZk8Hd6a7iLRi7QTnC2l8acL095Bu5FGu3zTd41O+GwIrEEMwTZrbW4WnUbwg
CHPYx86Y6bYEC9koPxRSRDLVDTlp3tS8+LHIP75M+GjCXTiJiZu+G+5bdnfVXxQG
bVxHY9SgVCGK2sqp+QkjUqnn6iAFYAJw9CxWPnEgjdNtBl5biwoxSPqnVxafOetQ
ymTS2JbRcteG+dpmnqhrGh+DsPIkqtZsoTb8nFK2s40mqtkRHdd/yEPCqA4mgmJW
PJqiDngFT+rgWZYbR3Vc5/BXbyTvnnVyUN/kHcVSmN/4vmhYG7cPY83arJ0huZRu
gtkOzH+fO5kMJf6uTkyqNdWrikjWXv8VIMWzhDmA/0rqM0c7gIyl9hxAxgdAgPbd
iV4pwvMiIGmf9WkmBo4llwaXUs8dj/9z/ubJYm71VmOcxrtPYijVkYAu7tsCzutS
pTnnvJdN9ohOGYg7f6F9ttL+yP1S7rmVfXgZ7GmDgBVTu/77HRBn5PMnE6Tva0nN
K4Enx91uEl+fZShqsTdywRdUyoGl3uu0onHSk0cb+1ugFLZd+Cm/XbvxUm2tgIUh
/Q+11K+bhvT9rcluitdSuzjXSidUZkvWf4rZezkhnxheYxOuXC/TPBHio7naa1rg
LjYjLOzU2SWpA7xHw5R2wKNeMxK4pFlfz5xs30CWMHxEbI54Feid9ZBtDXOdGOH9
0l6wF/kPUbSNH4SzRl7ZHneq0bWqcq+K+daKYh3B2luWcTgPyLRMabm8ccBXBEHm
QEUUzzFFUyy32bJtnxmrta717M8avMTa86K7hzJgMJ+pXQqejdOtF9ZYmyPEAuSl
Y2DPQ3AVehXFT6IC8PDsDh8C9NYGzOdN6Ftx+NlmBDozilk2/1GfO3jz9orP4VXr
JgtFzqf9o4/firzW3m6YEOAvrPsQLMzMS6ib+LoUmRP/ub9y5B5DiCkKfUN4vM4z
x9VbAlxZAQtkP4wFRxwVd8K2JzKHky+boZIJcmszblEixq3zWDY/A/RCiIWowIax
DurETv15lFuvQ4pwg/yqaYHahj0+7REj6oW6KUG9KZe7FFf24B2+3VCVqtvzrgtv
JBWND3TanuezoDgjw3qNoL87C3J0FyDH0Mgp8dEgHnyo1ybNPQaJlUBnzOSlkVCX
EXmWepcwmDTrsSFzg5rQ7DQUNhhVWb8zLIqITfhBQWnxRR4hPQf0hVpMZasQRKHW
6pgyhxLq8zha2SWaGVBTFZxfaiYc4SUXqFGYijuDMSvucRObzXTEa6ZiiZw9kJjX
m4piUPUS7BEIK9pmvx6LbbfMPS8xMBUaFbhk+idhy2lY52Td1QW6E36yYJsl6n2k
bv15F+0wCTQcugR5FtmUTncmWZ0rqwicAvH5kQvn9J9kO4AZwcqeBkIkX46GPnuN
7kx1TI3BVMvJxDsAeGbQJUBmDVn2sBNyuTFwxjhoa8nGY4QyXIc53utlpv3HhAAT
dmRsMzZVuSVU8XCzFUcDe2ebOkUHX/71Mr6R5Cwqj+1/fE/q2x2ztUyB9VoFvist
GsckumK3wbW8FisXZnRtbfluU6kaIVw+/BQBRa2I+9aOn43X0kh48ys1dbC2pL4F
Yt3YjZKYna9z0w2766ATQrAFbk9B89K4XFMuZsraHjFCRkDGUF4lifsGAHNIdWW1
AaNGNvbESKltTO6ridbQcJlXybfRssR6uHezq/ylzxjrsGAOeTb5ObMhrdfrFP0L
rAnhFHBPzea0StB1RCfZl6/r0mhzQ74JmdE+I8IKgs2cbW92P7bjUmxFiDWPM1B2
xmYy2zBi1MdVk6d23vO8dxCjGGR1VFJpGb8RqiydCQlcmQgmsSWPt4stfu8GsnAu
vRbgK7G4Y2U1hBMed8/OzEsY09mjB3wYWjQrELxsX1DAubft4NvNi9mdegi/tGrw
SSH8NRFvCQ6DH1kYFeQWbXyphMkOFSpHZROZz0iK12QlJyGUg9Y1vd7xtbw6+mQW
LhNY8U4oRa5NEpeBQ/wt0qvi0e79FDk3SM54L4kQrl18H78RM6ZRaiVSnecYl/pb
+FQhXspfoj5KXzbjS0u0ELfR685Yv8lZsB3tb18UVvgr84VHX2Sxji50KC7bJ+Ua
YUNIilJeE9pMj3oaF9OWUxqXJsU4hMwbl/W+Ni1BYAo8/3gwRZgMvjkSebTodSTX
VWalWerCTs7DLy61k9jEdes6AZf3vzBNcD2PeL4/cI5qTLU50tHb9I+pQziMIyjq
Q821SIGKHI3/gFUnXdWU0zUiMYD7gW5D8kqlp6H59AA+8uWRa7jXxr/KVCuLZ8Ff
MJJp4r+uIKWBJWkVFdSi5j5vf5UphLrPzJuZYA9uTjED8cZJqAoSwLiKn/OXduPL
fRApjYYgJHMCHIYwAAV+5+4R97Jd02wT5t9iIU+fDBzj1ytXOpmxtPvzudVNWhTg
yYWpu/UzZCVvdD/nG3XCkznVzcykcr8m2wpqR3hgXQuSbRFogok9IEX6lvyuRq12
quIYIm80KyiVahl7A0M8TGLaVJItquDhsjvHeL2r6FrnAd8kk6W2EkXdZOWuIQPg
doOhMRz5GRTXqbMfx0ZfhoCcGzElovO3iWTOGfvSHtv6Up0R5sIDhXKj8LALQwle
OA3SamtUI77uZ4Rfgs1I1s4fvUVksCcyCE9gyLuo5bqSpC03iXf9LDKIPGVtSmL4
UXDnHNDMo8ZaV5OyjW80KhTw96fTATRzX4slGgMcpvIpbisIXPxqxqu6l+vOjGzi
FFRcO7py5HLYbRHpertOng/xx5Tw+Aj38ejNQX6Uw34bR3Q4TofZL6mNWOAtGhJs
T9PzBP9V+f5j3RVHKRf04GyuX8srFFEGUMyQQ2OeamM0AcjzZfxOieuk70ar/lYC
7Y2jUXPSkXpcUOI9Tmghgjs4Vd8TDSDqyuYjVZrUUCPsK1jgU/i9BiRdwwTGyQRU
91+yIhHU0bAP+1oWO0QOinctK3pAHxPIuhK6Qp/IrvG0vubXriTpOqxe6ECqQD55
vRurh0rRsBF8oNpzs3Fb5NDDcLn9bP26o8TvJFzA/TpMRHALo6XRmBwbzs8+hBJJ
jXUho1Xoy6iER4ZPOnLFZ0xm8HEGBII+87inA7Su0BjXt+sXYVeAN3taCeGcgRrz
bdxynpQIqupTyGspFEftcgPwMJvTbBC4bym3jRUMa6/7YLbwQDdbw3OLkfqOfXgZ
uGxyrAjEO1FtLsycfPJ0ObcVkFA17TsF8JcUXR/iDn5WWRnUU0wyYxfOa+czH9Re
u99VBjuXtaM7i4vq4xMgVomFFFVMZIMfftCOolxfQdGPG+bOQhRpswLZbJuSTTU8
CE4tcoVGpqa8RE2VgKPKXiOLvXRdS2y5gwXsNIv9N8trtkF9rSV2IxKnW/u02x3h
DJCEzF5uovJBBTBumupf9DPj9SBQIbNzGvJoJ8V/YiXwDRNJ6qnHAqnnIhNISXEF
pRzXGN+z+E47nCLOo/Mkz1bwkZMyh7LWKFnQEGTeDTGBknrdL8BSlpScoRHj62Bl
Ehs/mc0/179JA8/t9rKhLHnJS6bKmdnnbBMEiW2C23VOv3LMloMrz/6G/H2sbgUH
QPcOWOOLOaNVwx7v/hN+JWympnlgjD/3Ip4W+6UqzuEFrKid6C7mG0geST7eL+je
jqm1h13hgRA0OjE8QBX52/+wfCQH9Y8NKgjp3KLt4RrI9+RficjCQP0aw2Yhat+E
2SlPBA8/5tJft9PFKAUOLlPSpLu693PYPKZfSwhlTije9Tsp19vomDIRNUsu80we
vBAUHztgOMdG+snAAIaG8e1IiREOKN2uVzaWC6/agWt/vCJ4gLjT93JZIdB/U/fZ
LgXcJiS9LPUGamKiy0Yllv2OBAmYmJSutp2MgLWgPO1Di7p6GQWf579HU8PKmzfT
+ojPIx2rTF+AvWAl9uVwsiq6eZfY6s8iJt2pUFtkPCVhlc946vOo6mfbHeswqYs4
fOuoxvHuT0CSngk6lFozknCJMpNWwnoRezlt25q0+srYDIHmyOYTLtuk9WdBdiK6
J/FdiTn0TxAxBiU4XU3p9S3go44DkEGQzzswdy2yg3Com7YaaQ+rKye4yPrMufaj
el12sWCT2bQOOnvQsw3GSQFbnN104kpDOHYLJUG5IiLvffZhrLjQBf05gdA5dF76
j4HIEOrEREBZ1bSA+K6jGKUHy4tjZUj+rEXL/JAC7st5oV+9u46+tA7O9/dbVA5d
Vvp2G/5CS85qHf7ueYr3mO5L26T2/P12H1A7K6kx9XvFB2/4PonYCv+WPSppPp8v
29KrFwmHhTuZ7CavQcdcux7F56pqHydV5F8/5MR01XPhsaOxcAOMSqpxkSdmd9Fb
MbTTlSENu/gIB8hcVjP4j61Cen3GoGS8ckaPI+xY2zUNzKmW9x/HjzW+fO6nqZm2
HyIYqbvNUyAOCuvvgfRJHFj9wE9rKKgEA0yWP/inGf+SigNE/aXV2M2VYicSd3Mg
kv+1or48llo3vYoYLHQALY9hEeTk43u9wz4WIXbS68JdhyqDNO1mJIyQc/hvaBDS
/lDWcxmO88Z5exqU73qCbeu3CDNRnNfGsShh35PZ9xWiPpxNZ1zSkxE9+IW6jmRR
pbUIL3quU1GQ5IzjsUJk1SOCbiSQ2KRsrt0aOhawtSRLCPU3uJ6uGQxVD04QS332
Pft8/70S5BDKzV0RGJaLYo4GTpVNQxp1jjj2s+PaJLIj3A07fuuizeOE8UMW5eVb
x6DtKgz3B2TWv/RM5dgbqXAj/YURekkwUXXe/0PvLWqGPOOxn90XK3jgFRPhjCD0
c1DFrwlOZlmlpXEaBe9bBZhOmd1uRaubGk/j2aGrmANeZjs84WloYpstErI0xc4Z
x7Ta4t1m0zk52uqVdcVQ+81eso7F6fxcJ/SYM/6lbmGOLFzCsyR0edkzbFaU4Sfh
uZt91Ho+zUvKxewaidho/4flccxm0KLHIJafe7cD8eTn/J41KUMWKgBlQIee0yfE
xwi+CKfYhP53tLI8iIU4bzkEB3hbMZEvK+52mAtocd5yVIl2NhxSje3XVXpCHH5F
V2Xl3btD7zlIrqQzAa47T0Wms5S9laC4wphgBL1mq1sRd1AnUB9IPxQAaBHHM4Sv
lmpUSQld/m0XwbNqgKmhFYFC7RATFgWDtaEjOzVSUpbGKNZByOY1iZ7um56AjQVq
joZVLkjB7a2hhAQkWeAmpLE46dMvhpBb9TsiHmInvZJYn6yxuCXOMn2fxyY0DBh6
VJ8Fc0X4+0e7oCJ0YJeO+KWQlUe8sj1ElottrJpeT1HZ0TePKybTBbkBfnGU1N7l
I9m/zk0A3cx6VJvGS8VB2ZjP7ZhqRnsOd74FD7Ff1esUQJsM1eqhnbwfxU8AAyzp
L55P0QbBn307tQj9NnjxYFvx2Ods+Xy40lBEZcwtazL+N26rlne+yY73t3/R9Zu0
1BWEgMLNlOo3O2IiOe4uWL35O0H6oNhgGQRJmQnEzJwTSMRyQiFE0OM+/m2ApBdm
j2B3JahSSb9ptViXnlZ39Y7SoWEIeQqXmCwxgmXj2a8xoiPOjRA7qxNbOOI6jedC
pq3YOIkqfet4HRpv+GyzdZ0dXzyMsEJ3dsoFuwawEYOlMUWKSlH5MXvXzMTBLwAe
zBMeNNeozpHUoqYYhzN1qgSton85S+Cpqix7npD0Ird/LGOBvQ9B5akIhs9L+928
WWuIfGwCjRBWSiaiNpmcpngrogun+PuPh3mZp455Ar9f4XYsChfBXrF1ItfMJ+ro
8rhyh8rjxEbEwvAdErEKU8TPP4EQKD803jIxUKO7uccbRnteq5QKk2Mg7pHDrgiH
N/NCkK5RXjmJhdab5vYesxQJ8z9d2GzghJRICCAVRvovXHbSYlY68261w+EWtYOU
0y5uNi6dz87LCNCSux0bmgbu0kg2YLE/1HMkcz7ydXkuO5ifc3Ps2jhMdkck735U
FiZeZg1Dr2MemkPccfNfvtt5Wn66EAOTx2dqAa2Jd2WltaNjt4BA8/JlGvV5Zm1r
BPk5lP1szlYY0xAGSfoboeIpf+CzLkHOPla7qnqC01nJnWWw99ImsLRKiviuVZIg
WAobu/3JrFjZJ7jNsvPZJ3QfDa51866v3EyI0qWxh6fQR0XQHeTKAq/6EpeZHNgW
seNhfG20GbsuEth3y/zaHQ1rEqCkrQYNITlHjE9T11K1A25b1XqnjBT7YuEeW2xo
xJbtMuFYYR0VG1hz1CWymOTvXXdZO9TJ638yGjW0l6mtMu3kqhdP6dE44q5Foaa5
/kIbrUy3MtWqLbIo7KoM6ubvHLmu4psHg05iZqZWDJkCTt2uES0/HKUAy3AI1Bm8
dmTacjalDAgTGkGidQWbR9VCTUb6WbrTSziR9P8hkZapAo3FX3Bbg4ef4g2BfjI5
yOyNd506SMMkVaE6N8BoPdjYH9YwbEV/Oo01ImZgDMJj5wJ8fPo8YNAWfgW2yH5s
TekLb/5kDEdeeGRgMaAu4ysDevMCBk2p9S2tx2JB262ONLc/T2OgnTCWcSsAWePX
+6f6leZh+ugYZz0mrXABIrwdNTPF4fXJaouaQKfq+Gyx0ue5+qDWi225z+Zr+IU4
qMp16OttqlesJKNHwWURignOahkhvZTlE0l9AfjomcPFgBJUzX9UUMUbhV8+pysH
QXok/TtnzxQL+3W1d+oq6HNxqgUj9X7PFkflKEyBeGFbQm1LnLKpb7XI9XY0CVBf
grUy7AiILV4i/SbJ+BaMYRsGATCWG7ND6o/Pk2/lxeLFw6RQ6ZMLqJcDUDxeB2kI
/GV9XYgu2lXAaTFS+qKCX9CDMqSFesOWjcLpqqZvtg5xow30CA7majYmGZY/IvSA
BBjjI4T2zVO5h2ahOmkUVsl5/Jw72qoSf8PaAreJ3UXt9hVtDlrCLuS7fDWdj3JZ
BPkIx47HvJeZWYzPj3yZKLWimQw8o3pkam9vE8haTy0xvEdELWpDMzSsaWHPMetn
+rjdd0Sqoet4GMy3psbHs4FRnKXhr0VFEWEMmH+6JVPP+4LZucPRzSligG2II578
gOmj3WLbCsL1grh6oMatA44xZFjh/dMtifZb0M1z47bPBHBn3yWP5PbO+QnF21U8
8b/0MnlPyk5A9hh8j0SUWclcUwP6LB+jnQAWZTgEjFlOLQ/cVbdTXLDPtdpLKA7f
SaosEH+ZJ9+xm0exCdIPos4B1Fu7Y3nkvZ07pCXP3E0HRqPC0ejuU7FinQPpFAUz
7QXQ3baPLxhlLmCBaByJZHgGHLCiet/K3b01JrozNP4g6rJ39b+LIqRebEk7er34
HSnjGDEVovn+cidxovpvHJHaaT0Lut2N6E81rl8naS377Dx39eLQP2mpWwrT889r
69lr+E16YVjYG2zNiVYYs6RBal21XniSv3R3pa/c/V6csySdhguPJCAOEI8YIBit
8ZZcAFve9kbbE272PaISdNqx+3M4CaDfs8EbwhZaPAFRfshFY4v0p4lKI8toWJeN
CIPNjiDejtEHI5ytKoGGqAGFqDvrJXTiSqa06vZL3XuACCa/iDQe7761Y6/0ozVc
tRowaP+CPsnDs0xYDh1N9u4RWAEskIPlJzhZ3+Ngfc6ZLiN56o+IDAY068aKRNIB
mCgr9UNRmCBhZNoTAoXq6dpo7ZQhINaO3wr7KbG0GZ13tV+IzrDOzEhzB9qpj1dz
rQQPhXvs+MKXprAcuYVNRXpxSTRqU264Fd8PWz6sYSwmRmFBURJTLTzA0EtFSpQ9
WZQeczJCNVRsNRf9G3byrjZDaFFSKFJ+VK2Zf7oZS6Dem5OKhAszsOFijnKzXu2m
bvzfpSk630mXgMmArVv5JYGXHtGLRoWP9SgdCfXhr+tW7wmAMIBBkQDenR6x11q3
3SufqYeHbQ/aWel7pIsDLYNKD7A7WtmS/NV2oxHdZsoxeYVsz8ZxSGf/rm0+256h
IjeMOkQiQaNCoB/iF8Yk9UswMhQqw8MMatUSHWxcH+ZuwcCw+lNWQfMINuXzHFJi
3ZB+4Wc3Nb7nw/KiQtb60bDyhlJMrlvdJzDwMT/muShiGAvLJFsGeJx0t8jGfjtI
tmNd4KDKLZvk5LHUqJA9r4pHKtcEbJnNSZEP60miYP+Dt8kyy7q7NdZJSVL0TGSQ
9CtdYIBOTzJpByKVF7Y7/nlJujeY2c0XeYbIZqrLTMpmIDEicdSC7lqeul2FYa1I
bcAw1Q8PY5ANVSGiAOdF8YBT5kL5ks6o/GQqJLtxtByz8x3kabcHIBPmPMA+vKaI
Eucy/BRkqrNw8wRbmkVghoeuc/JuCTDAFAGxJdNyLW87xkLk6B1SI8a3oBFGW9xQ
oJMvgLx/CbdsDres/yXZQU7u01qwsmANEKb2nxeKH5y5WqB65ur7/KREytv20oF9
tZJzpPlmApXTMfwqY2+jUUXBqWF2IBAReGrv2EwQvRUBUvuHMgcfb26ux7dow0qU
MIS0P0tB45FtasTCvv5VepsoE+sfB1lr/zn92Hsam+H34k0ZG3o7uvTK8UxqVtDl
JQpx0u6/f+ldtHyJlG5g+pZvlRiJMW6RfirJq8Tw75rKXiwHrX46+WOjc3Xaw7Ua
pW8RRYYGA23d/HmbbbcgD0AW2tQncC0Iy1dKQBYlzNjhGG6M0oHTqohCGA/WI7Rb
2RlAM74/CHcHDmlLml2ZBqyM4l2XLMcONoUu56wT6I3WKwfgmD9JmO8VDbQp/C+B
HHKMTw1/vul+jn2emaor34Tso7M24sA6itiAGQ8A9xI14S7W/1bdDyxEczwIZ0Zw
fZRvUwvT0I4DSlmX5HYeT4cKgU4ptKUIcjlQF+FIYvrneLcL8RCMPTEE1F0BpGDG
k/fgrON72hCE+Vzi5v7LaEdYPDTZZQT7T70eKzdj59OqGqtY5+eqXk/epx7NV8AY
SF4wWBIPMOOllxUgwBeNAVaBrMd7JDa7Inlf2cMRB5TIqpDzDemjiM2hhzJpFrvy
zAyi2bFZBvvVtP4UXmYyGr1O+iiXjKYxEH7gjKEMq9hCuDyI3pptCPfXCcZRkcOc
Ez045bDPZnAyyi+jxwJrYqmlAC0TRRGpG4bwF4hagGdg/5M0CdSDAu1pdBbNTD9b
bf01DDK22vxwxxQTObplL5laL0MR1PTZHXuUB48pWrzP+NctsKdW/yTdpew6BkQm
uJ8ZIC87XMMFvMS2c6I8eUgWo2MpI+oZdMrRkOyqgQ0vcIf/IhmZI8EEENO0Yehc
lbMbGQa/sv2oQileFXTBSxtEJaJMBROG43+P0ATBEAl4Dl/28x1ROtEzQFSh4tX1
SLydi16qgU9OxMU4+N7Y9NV0HHfgsLMfboQVSySd9RSj3tosILEWWXPNcWrItEUX
V8Mh+7StxUzaik4KiOj1qWVyiwmu8oq2Fsa9zAJvkMVjJ/ZuuUxo2NfqDQUSTWTo
wpFd1vsPBSnfhs7Ptn1fzl8HPdYZdPSj0LaHEA4CZCn6ke5kT7Zthv39ynf9yWmi
0YXn1aIEaxHPBA7K5mmppz53Jyfuwvvw6nSzu5hlqaZS9VBWNCoyiaFEnrJfmfMu
N7lT0qgLALengPz2S+CulrG3o1NBTz7/O8YGuGDMKhSrWeKWEuppmmgGtVNtQqqS
hvQs3rVLJP+zZ+0HtHSeneJ6r8sPa/owkc2OgodH3WRfwXxEameUb3VGqW4bw+Kq
BvGTH9bpl3kqJDWLb9K9BuoVgyr7dG5a2PFjgcJKweCs5eGAf4FlD3quxfeLQM45
SfG6WtgWOI0V5HL1CdkqMLL92MZf1Szi1A5VPN8pD9Yq6iqxZ2ruwgSSEKReRwiR
WnoDIR1w2aAlDFfPxuuPME4KCrs24rv6t1Jc5sFf3Z17KJmfV8vxqcYaD12ZBZfP
Btyzbi0YInuBTp4jZAfzBlncPqXPzHnNWWLor8kqQgmi7v6RHPX6SUUq04py38U1
tbc6kshJH0IedO8EwlvSXsiTyeaER0z98LkTOlKeT/nPqpxeIk0qYRV+F3OdVHq5
GadgbrMtwwq7mRFkE1Hi4W/lvxsDBPQ+609anbnPihxofoqmVs1kinAbH4CuyOUr
EThJCmvUGTpXQdrpkhDIszaOImvafSsSUhRlEtCaEmNM2iq14nc0so6KCWDNjEtt
ltQ9AnlGCYyLq4V8qmj6x7SL082fYC1KTKWvMvYZMqlZLTzbeWUR9jcONOq0A9RH
B4U55Q8hOhtZ60toZnIem8iaNzeEXUYsSx5iFGtqjKhXbVIgNRPZZiSj0aW5OrE+
K7+l4ILArql7ipEY91/a6g0jbpzz+G3/kbwjCreW6XgGhBdvHM36mKGA/Izutx3p
HMKST/2/cexPL3IPH9q6hY0drVHZP4V1aemhEwMMX20wzzHtPb6+bEfrInQN01m0
ZHUONPdZvK4ZXTcTi9kSFJQUPAsmVMpZJwmKj4v7rQsyxmCBtdW4Fgz3a62GpVQ4
SkPIWWDqqQzcIKCJBOfv1WdsNDJyx+MZEzUk/KWqWJsuspaJVnij6/kZhAaPknna
dn0v2BK+sGTYcRY+6beqQE7xUrLlsqmWgeuTOBSaexPM3raQUsvRNQJwVq/XlAjI
aR6/m+AhQe5szPMofkdckwvh6M/S0rB2tsNmlnMmoL06hqSu+I49pI+92kTqyoDa
iCVgIcsuan57M+vY00wJ36Dzc6xlDicko302VnYyX6nD4MY42Yp2c5F+Mj72TpXg
Wsuk6F3Rw/nPVjOw7Evh4UvRFskx4+KtNlOrVVbAU3V8RmEwq804zjxJxjqfTiu7
hozGuhjMD7Y4bLiOxliZXeju9Ap0HguiafMGLlqfXPGlsVdpXgQFiIoyW2bAADLy
xxUUqwxIK8KcjN3Xk7OkjrId0NaD4Y/7GFS0U9sCiY2X6ctlouxcHGoJ8YBShv+5
apZhMCQJqmf9hm83iBTeqjtdUxa0i20G76dQcTe1bfrTLKJvGIiNgDDt8SgsIUkS
ZdAHECG7gc4PAMoev6mjVZXsqwFNe18T5xWZIsaUv1F01JZl2A4Zzhq1YkL9bTr7
afpz+/9iH4NpmTx3rXXG8GQuGnNeJQ23AS9X9SYOGUvRgBLP1bMtM9dVsbnoxe/6
KYU++52T05cxhsjqRUBqK3Qi4LhZJb3ljdmxY0DiGqqkygkGfv8WsS/rUcdeBt4+
b2m8vDT6RtUuV4iu9bIMWjCUZUSVwL7fXswPK/Kd2zvNgSt76iQrlJobkqpGtFQ4
MbVwPv7S7loeO+mxUF5+r9fHohSiiABqnqyrg57JCpdFmkF7RomU9I1jyMkMwNei
2jnbSijXzzECxqLqjKl9mLL3IpUmXzdVk373cm2GD05jQgE0HBPD9sTASpF4SU8J
r10ZQ6WM55nhpldqwthjiVtQCdyyKPRzPGsVXRwO4upaHoboN9qQhCzHHklpv9Qm
B61jWMfPLO4UJLyxGTiMyJsEkbtyWfNaIrq2tpq2CeB4TZl4fAEpkBkU9e4/3VxM
Rmg7D5DPdAxygUvmqQ53alJw7hyQct/bVpmvOqj1eWP5AZg6ENG/lWKnznPQkwvv
5Rjr+NiXo4ZJnKh985S+8ixaXmy9zMRKxPmHVbYVLW8pmSqLhk9jO0snF7oImhU0
LnAwEJPMj+VUbM8QFLhb+vfR3criVN5eGb3qhHg/hNVJRWJr/dSoRnXxBWqJacde
EBajohpMjUdaj9rIh76idELO9Ur7i+04SvvDFgWJFAUyQSRL3DP3bMfGkmEHUrEa
7EockX5y/joEppoeyfkzA1TkDvXqBrmqi0RcRONE5TjJP/fWA1ob1NRz9jkw95Tw
pMWMxfyXEAJfVVX3trQGAgYuSqTzXqBhWgwvaTmBhgzbmJrNSTxAfaV5Q1ZX6YhL
Zt3qTxSi6bcY8g4cZBqBhuydljEdZIOPn0TDtvJd/jZ9P9HvH9FmGJcIZS7Gzf2E
6aAmN8FeKOLIOslW866nZ7+pw3i6oWRqPpe04ZbnDFiif4k+tQp/vY0SIsP404W8
uaNWUD9i9plDfYGiTsyyPzHx8lCNOwr9sHHF7D5U/AG8rtXq+n5Lel/4vh/3FTS1
hnqQXy4AD8IgkKUWwIp+Sw6YRYac4BG/0940EtHx4WokgXupQzV53Jgx5Hk5AeSi
zaSeLv0+aWEolTYdVF7ZOLqfprPDr+tSHRBsP6bdFzRi4nbYaUN/+hMwF9WdwCx9
fc0/wbfbLZH3QswaopRDCHSz5VUZGJUYYMdN9NpARhxXY7NU74EWhzDsjcS1P2pY
POxVMds/L3MkJi7usxn7zto4zKjCngexU19lOQljHXdpeMbTn/wnNDetvV3OkAcm
gTdWMMuiPOp8uYsy8LCiqP5NCwx6uY/ezwwVIWVh29YZkatzhSiCoNcooekd13bo
qETTsPTaJdi6llTXxAEDlMURPjo7w/oqUVwN8sM6d6JLoKIF5e9roKlUyaIbiI8d
jIX23xUsXx45ewCfQfX5KBxpFNsEe16TrQdYNmA6qZBd6XDZhEO9ci8mOe2pCJ3g
jWr37OBGhVOKcoRdmsNFu3XaYQGV88N9VHgVrM2hRvzu8H4njO0jnFdr4KY7bBoZ
eI9CrEPA2aZCA2W5bzP+qK/pPQpApiHJJlXTFskmtQFhYE5zdTgzr9NtJ7qSXUQg
QU5981jjSScW+U+oiupZScZTSd6dtdsndKCXvIIjOGSu+uVLMbAePspiRgLLTCYL
XfgB6Hx1ljcgwvq29jczSVccy5p14iLfLjY9a/kR2oA0zg/RGOaSW9ZmfYEPiufQ
11QBQiAVyIoko0YgOBK9prkbiAhrUSwGSGIcmplgKXnmF7DFwDQIu1Uaq3pB5qFj
l/9W15EQ3kEqCcp39Eptec1UI+O/JT09qZdg9rGXM4V4TNM2aYrUxxz6hB2vKdxI
fdpnKe8AVglXvyL1KVPinv/CxNwvovkWee5AbClHMUTP7QtfhnjUSw7DmGMAENjY
8Ppq4kdFuG+/hztJPEGXvk66bjbp9mLvjBkuEjgtUNsjnq/dBvfNVqErrtWkx7Tn
JA1tT5qpkCetI4oGcDM28cqhv2SNmOZVhrJ/b5m2vOd2vsY5MOPYFt0aCdUIAVRs
No4AQckyq1/z+NVg+TciCYdvkH6ZoLiTbxYZtOm6zDmvqfjFzVk8mkcndW36WzXd
6n68+CHU6kpZMXkF64qeej3gxLz546HUXqMVL9qVnWdbWCwkPT1DJS+D69h6X00q
zTlmZ31ujsO13bioCorq8FlxDyqCKUcyvKUBbJgBffgz4ElNp/fvTAP3ksS8WVQc
zBUv9b5OIzlGrlYHT9q3UXcY8pz0/8ZrnmQIQGwrqePDqfp+iVUy2AIOOmrUw59A
yfDBfvq6vpUeJJ8A0a3hM4mHAWMLEuKk1Q2GwiKv8FmQSIWWiFWeowzydTdsQf6e
YVjVFeXGwtNWRtONHOb1eZ/86rTuOZCVdSCx0Oua8UmOCiXFC5AK8Iso0arE0fff
uR8BqUzjSnlDccQZk6SWfV6V+wzWUkbwU1tCDUNV4uieN/CjzMW4BfdPsfuHPZKv
D/FhcWWC5koEYsP/zs6efRZ55PGYnyMBPfoAGYCGY7vVAwNAA3MaiMq1S7tvk20G
z/GlOgEJ9JHv6jpMc9PrETxLY0xVm6LOtk6q+xEGYvEGFCwZ8H4frmNMYPHk67za
mNiNN5jeVBDIJVhX7yAMeaZXUwzYe6ftL38V3vNqHiC1aSHo+uSPL7jT5yVZquPF
7AhQIFL0YohKU44IE/48yPIdmdJ16JXvoGpxmd922XP+HMDIqN4KRIUGLcx497tq
fiBIXF6yVqoxBG60MEAcxygqhBeysCoBjKsQ3IdeJ0dTxizbptPUcHRroI9biFwQ
dRTE5CT5mAE1sGvOUMo91gehuRVkL2ybX1Y11wLyonV7XL/DNXZaWTMaOBmau0Y8
fgeDe24/exnzA8kRLhAU4JlXl2Q0Om4mFPreOSluYzUd9c9IHz7OvitJCXikIBcr
PnL8u30n+/DZRUsqLMMRYD2jfn21rqmETRaKLaJKYZydTBdfJm5EF8UINctW6Viu
QLfO1Miv8MVQroW9Ed2zA2fki4WRtLOmqTWw996OuwmV0mbOFV7MUkGru2vZmWfs
CgyhO7EpUmWyna/UnnoVxlp2MxV+DMGqlzvq4OwFHxCAntKS+m59i55REu747ctI
f8F1UaZB1cck/ulCcTZvz6TBKUH3LRPM14FOjVTL+P8nHneg0RxI5MjDkoYKp9my
v6CvPCsOB2/fSPnw9kEnVAgorFlfu/PZtBotumjm7b1qO3EC5ogzKLQ02W2WoJbU
k0D260plpeudm/Av29ULaOcN+m5JZjApewN9U/sWTRene30k735YWywr9BMML1aE
SD1yUVK29Q2XuwoCXwqiRoXbjrZKn2IbuCDiT+WbaJqOpzBxPP2uoBxwLeqvJ1vY
bz3ZqhQgokC8CtjlhDsrBV0PyihQHNQEwhSrf7rF1p8T7F6jtwIsAatZsWi+NLSg
OWyfczOUBcfTsyNAk3XkCszuPp2+wQ0HKcwiU+8CcsVUhAmXjLmEdbFpur79Q3fR
v3dYvuVMeW6KJMsbg2hkhc5sdRM+ahPFkOmHrgqP02mqbuxPFFh2lNb/s2Kauv4P
DD5OrWOPFqfQdjCNMKLkORGw7by4CnrfyT/z1V57ZEBGpRdavHmfGWjW/3pD4TGO
wqlCS2I+qs/Tce8uh7qzCJRelH1lsXF6sdOJdt8OpzR7DCv0dqP9F8Jelce4eNMt
TKSID1FHK1V1DJd5lTJf4/AA0m2AGse1NgE3Er4ErvCJHNVSrS3IlI/VOidXWY8o
`protect END_PROTECTED
