`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r+YhFxBlhMgKOyxhMsV9pVuO4aZ/uU8Oc4z54yBKK8OlF8FKmCCPXf0CcJ+nbKCz
rPqAm75FQJC4KFzZef9CgqUBQcE2WFEk7j+Tq/kYQt79u30S22rw+jdhTkLVcAIe
Hv7zyo65aDmlHt7y5jjsV3irxpbrVP1HH1RR4fIuoaY2hClclsg4UmLphcRhF1DY
whaqVawmpvsT3Ca9RvIL/GqpRz99LMMt2kopf4t9OOfY4Ht9Z22Tmu2Htn77rDRB
ZfQ72mCLuhbTttxT2C4ijWuydDqIVSvkrmATwgmodeq2p5a4HQClGiguEPJmVCkH
r2YXqpXfNc7cQ+PWnm++axxoI5kB5PAWnEscaPJXN723LqNuKiJDy1PJKcIjTBSE
lIrINZ21dYeY1E/OUu/bFX87lZ77dNYV25pQxDz207xK11MT4Mcz8asK6WkudU7w
ZZRLC7VIHfbMWFgP6gehc3ssKOm3tiFZuL1xngwyfkrMPU9e4iYhobB7UsWhCiXG
OfDeVBaXFAh+Ryc+ocEiWwv3Hcwwujp52mKUrI4xExX7QjAJryY94ij1u789PpMk
cYeLPG0IZ8SC0sAa2E8Y+dEhl4OiKXlRYTBdK+goKqSAbZOkDQiWhi4p/w+YLxG2
Ijg5lyzNUREbXFHehaIJHSgIg+q1Hq0gEULZL8FwhaTosWMA5qf55Ewv2x6RibgI
agEEdNsA8vPccu+/LRsyNNfy1E0KLoAX/Df4ljFpSyEpAVIriFnnOWYWF2B7K8Ma
Osvq3WRNMNnLeONAUgWyMZeAXOCImcGC7foeC+sTkHi7+q451KRSgUgEPLRPsAyL
eO5uuXYZJdnEV0u7DjYUbW3uTObhpBgJooKPy48uqbPUVlaQG6X4go51VhWOzLys
5h2xVeGYU5wZsYMXbqIpOgSNFNQCwT4g8uMmgtScft0Y2ih0dwkkLBTqNZ2uJV0S
uFGf+SPelY3jOnojT+l+T2C9VmDsOKyx9dlRY/uPlpnJLO87thxQGZNLjRrKZ+9H
PBB8h8D084pMGgSAS3NwOTeb/eVZ2VozRhinb0praqVADxMnutRXObWMAQVrynhQ
ij75Y4pC1RKDa7vOIizapykEBe07DDde+6FGo6C+EPv4CSTp6PV7Syy7Ze/BffuK
B3JSal3dlLo8jeBHbHcu3X4MDr6lNeNRwyW6oT1V0fOnHgc34qgWNaflkspocXNg
bs8le7qXKJUI0a7jZnKYt/k6xPRn4dUVihS3rpgRz9b+rOjAXTF7G+n51n1t/00F
0xIsZFpS49ewimPSnTIGxPLMT7weWdz2durKvcs1d99TgEO+4P2aNiZGo4+Xp6MZ
NGuP1qCrFo5Q9r7g7rsdk954rD/ll780jQl+JYjA3sVCsggcEwT6Rzw+T2Yre4+X
I5CRwKe7+O5rj6ocMk/2B+xycYpVndgFX/rkCN93SRwlyeXnyU5iJgs2SGZSp6/W
iZgfGk5YxUh+EkI3MUxLO3aa49Mxf5f+UXi8ximu+kf0JK6JIP7+J3F8ec0rGjL7
/J9YUHrWcx0YCPcJqHf1YoK6oxHkWpzTBCgsEF3eNZzEG5s3RdEgvOgxnfncKh27
6NYN593t/mLIdu6Rd6kE0kOf/1JMBa09L9v649PUKGwENLQLCZmqG8fHk+s2Wt8d
AwY1WYjKPWIyvf4g8HL/he5MzY73T0QXahSlnq2JBLt/R6bvUgwQuZrnFyngrNui
ADZFqhnMpYKMTmJSNi+MkcfaMqECBnbUSoFUykUDp7vPQ9BhWgFQWVUibjWqtdFm
BgcR9hV4MZS5l3qft5cTwpfIokSpqANrQqB4JdybZgylYYdI3CoOm1wXh04zHhPF
`protect END_PROTECTED
