`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+MczfNusMWcY4f/hNQZ5/Vc9CgvD4Y8X6zg3hDfXGxFw/K6U64EM9eGaSskVtGfu
85RURoTdmYKUu8kW7vW8OBn5LoHcehR39UZreQOt73FD6QUK2YwCrJ9UkjmPcOGg
a8lpMR5yVlUJpHttM8c23LbTIwOAHMjr5nyA72efAVIOqjlto8GNCLrLGL9ICGB9
RB0DsRnDXqgNnLzUrT0JL1wdKKWiMqi96TlLsiJaFPaKVCeW5NkNZOGRkmR7zFvo
fCMHQIT3aIs3GYl2WBMictbQiR+BUt7DOQ3u0rtcRQ4vHpi46fPjYBrKN28xQ93i
cM8w1wOs3Zo1fzYrMRW4/wB5ezktALMqvwq7NSu4VEwkDmWRGaTnKqjOWGLSauaf
EgYlefOlOEQXBgqAeEUVeJ1ca8nsJndR9Ze9CeapUFX0hQc1VIc8oY4sNVt3exTE
o+fu4YlqA2ofrB9UO068+pzCLllkze65kb7YpjUvEU+q9awKcLNMzANVZ52K+Seg
y/tvqN40V+YKamE/cR3YEv+D1jG7E75HDoKRDL7Gh6lrpYoJUp1Gz4qdivx9gq4z
1CTlefPng4m8C1VikTkSi6+tXzYdYhJj4/idGGSO9c09z25PmQOI5FowYsviTiqb
Fb8xPyibrOXDZJI6/AAqiupTv65FZh49AqgLPdqfmRo0lQyrnscTJTJTuDQA8pVI
ELFJT4YtDjw/OWG4/Fh3KPZysHCaOHCaXrj2vmcyFQckvE7Nd6vXmLB1kZ9Z7chr
KPMkGdhqG5UkLjYDbwhuOp6aOTAv6CGt/bHgRnlqMOR+qdcjyvrLUHCNgles5+FZ
mYQ01WSGLz4zdzxmOYt+8HuFrLFU6WWeSWt0MafiKdIA4k5dAGUMrQsa2W3e7fz4
HydnppJFcP4zSslc1X27SiMaEZplXMP2r2pJw2Ec08Dv2ONRmRjzJCyLV/0lP/Tm
hwiJLIDizbZ/SiAIK7tZqNNkLaPA8rNL+VV70Mq5t2PtV9/XkC1ZkHvlaihDQnLv
1qKBgb1TAZop8zDoRUBUQ5AFtO1pISKNXNIPa10ArKxXgDWvM21ZnZz3OtMGMOnk
GSllmRtbNxkI4EtCKsPYT/cjCquEJOosN1ikEptsVWerxfycM3JCqlHZn0AE02Z1
RC/2YpayLKRf0a9IZGFtK+zwTiUEcTn2sV2XURGki63eLeRqbHSLyNDHKvMGdmmq
RXjwrHJFtVCyFVbTPhknEo4F2ZNPypPSNeTzyPQlxivHjtHH5SZVRQidNSUTFkxk
0+Zm6KzRY7cJztPCntMz4H1MYjS1KcWy7LMXpoFsOar4w5XElUQmDVDT5kf+qbUQ
Yi7fGr7T1CGB/BrQd3u+eyzhwCZAPeTFBXWcnpbmw/YrZ7GbnVynp4MYCT8Y/WHJ
G9xukHbmDDMhwAGsEylsmy1WzhukL02owFfZMuycPER4w8GVYUL8E8pkAki/ewFY
nhf1dtp/zM63iN2AlwSBzjBjDBFTS9deE7o9d0k1NnFrPrKXd1YdmpCzHR3FtM5+
/4Fa039bpARymOL4GzPcay66acQZrfB/aqXFbiaiu3Dmh9OjMpznLhKEmtdcI6U4
/rmSdF6PFxd/tKA5nvoDoEToomUy6ipwaHts/DKgFMCSTCzpq9velhG7eSktwcZJ
KvEDGvKpuoDLN1Twb/jI8NpFsxnw8ee5W4H0szHI5zVT9VbkE8EraU7cetxx20Rh
d9FLxLEt4fTdYEywcGg+EynLBsqr/+9/FkYsfXncVn/xgc6vwxQxTIQRovTLyG/2
a1tx/j1UMVJdt1NkSCpVkcjX3LEm83oaPTlNCRC2PeUs6dWgssnkaVOeqgYVSOxN
ZvyzXNymumNVMjECSt4a9yiQOC5NXb42PKZlPsF8xzDdtS5Bi5JvdkZeGA401NMy
DTvQOxorPMvIlUVZUcdSUTP3MVCOKhOyjWbODV04fN0=
`protect END_PROTECTED
