`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vgbOWvNFCb8SINFibDX3mkgqYxLXPnibld/mMk4U5NUl0jAeaUo3ADt3xAASkbfH
KQWD+YjOFWZoy1eX24yZ+j+Jzxt3/vHHjPLth/Z5FjOQhDWbA0E+Xt/t1h2Q4GLO
1psgXp4yjIy9Z2RDjzX+6lhaC9YfilA3VStQeQpNxRxqSBGDBHAO4yb1IQtSFrp7
HckOwE5TTSdwFoULsKauWYlcnsET4yXyFeA3gSDWjRqb/ei2KJSYGoRCEBS6Js2E
NCtFpFoyzU13I95/ubhgkOpDcak/R7IDbqXGkdS7ivVLOoNlmeXcjeKzr2TZWYX0
T56L1lgnTuIIeGXBY+KPtm70M2KyJAkhvzpK0H36gImqQsttjmpZSOLn5++rNxkg
Nesh73x8L+RTbK50nkk1J0IIOyyByr2Hr679YfNW4sAAiVIHGfwOtwU+lsgW2Pjv
UJlqmJlHSDLLUhiCp1KpFZSKe15hXaM1/yisPup4+9awluSFewo1cCENMK1b3Zxf
pNdPxLJk3WBjCTH/GVpyaFOzmomfy+fkz2I73xFqQujC/6rPt9HFXjt8xPSCOx4D
eDxsTdhvSb5eym7t35HOpN/h4fu7vs18Q2/eb8TdiFVljsnI66VN/wc7uC+EUseb
SHefdX1apY2cTUVwCRXmx8aG2U27Bp4AKyJBfNq/OIUbfEFFO0mTHUdZSWcFSx8R
Xo0/s/L7yQHviFeIhl3byybQPWvo4QQ5VSlWszatqPrh/NK7ynUqN4A9HzPjWL0i
t8CBxxZDOPGuvNlnQH2OIIeUGlVFu/7EtTHLiO887e+99XU18Iarq+0ng9OWv/Jo
iZQsd1GVKPV7fu8FFZQREGkhopajInAIikTGx7wCUebYrpmejDDGUxdNy0Dy9t+p
HnUsfTwAqtPb/v/fzhZlQcBTe3fWed+RIhELoRzRPFzENqLaUKxmZjPir5m3CIwq
VlEKXdYeu2Ho7Qw+boUea/ViFF+/2DsWS90QNeE0xgiZQkHc153uMyMBeHI5Bz0/
2wUEaJ/9xGrtmwqktw+lUn1oWz+IKhGmct+0NU6cYIYXmUunGfdB2vkWVPQT8vm/
Un2ARw0olfnsEWnwRuVSgrOEMCMFYXHGlUKn8kASrVp0D0HYPLLmzOQkaH5c3erG
nBVl74BpQeuXTwilkMGWS5kNoOJ0X/7Qp7UiqCwDOUYTX41kZf/7HQsrESVLNKlG
1FVcNRn3t2isH08RXxF+7h8GU8WawvHjPpor3kOZbNyFAahATnnZp874le7tR9cX
mo6YSLSt5fC5rq2ra0zjcKvx4jcLH7G5xQvk4In2hRIAgKZmQ7KJv/7TrkKqebG0
rMUnwjCNypvWEy2hspJefB/QjffdZPe7NlF7B09adJ4h8ypjs5rxtBtaVxQqPwDm
DsQjZunFAPlbFuqvVlbNvxBIb7KHQ4mAO5pMiXLdTxTAY/DghX6sWJsrRmqJnY/E
82bSdi5KQTTiImbgOuTBRYjw4lSuIXuAGo5ZJDdjK/11Utcw4WHSmOUkjpr8sPZ3
33H9DcQmdxD5KzGrBUSELpCo75eHkWojW6dHxmeifTrx8E5TDD+MinVw+1zYwMzD
Ji0su/URWENn3bdApQ45rqTXMm2JJBqFMUNE7ktOEMOTe4ofAykk4/w6UItm9HZS
fGb7qvCW5ADbi0BDOSFJ5MKTQ+9+t8JQH6Sb1ZG0saLmZgyCJf2Ay/twhakj6rDX
BGZOhUsn2sAUe+t5zIi9EVM7Ru5+goYWscdrClAa/SiAfQCRGu7806WPQTTIxndS
zPr7NhKXQmhOhBpIRwBUwgB+s1DnqsDps4HKdPUQdOJMIUOdQF1oKivG+bAfO6vw
vwITw0yhs/Do9s35NYfxsj7bLXPW/ZvXo++wkLhseHSx/rcRGC3SjWFx374i3LgI
XrGySTGamTrHXMpxIrEiKIJ474VYadg0X+WdjXCuotMmHf8XP2LYvrAIZDXin8z2
XpQSCORvrbVrOdQO2O9/uqWEYC4r1gEkOTU3N5xTR6x0HhAXF2OSlSyekLCFBH+E
GYoqqa1SOORL7eUPMJfgaiU8qLKEcYVkxVzZGCKsKDJ7dIqmw5hKbZ1luovikCd8
OFeVyD7RD2TGowm+OfUwZvayGz6/agCIhFdpeDeI2P/WNv2I+Fca4p6PwfLxcmcV
rhROQ6kAfdfoPn6Wb5Ckb5Oh4gqflizlDB0fTibHiTctopAwJePe560pnenl/aeX
KmltiPKA3pA+U2D8OW6rMxtFZMqfK87gFTfZ0y0zWItvENSLDsZDPSGHJ0CL/ntJ
m0j1G86FcJblzo5pRWTvp98dL0xcBFf59c7ZpcriuumKoZOMSAhSE5AyzKfONI9y
Kig0g/Vn+LpvbyaCOL8YMlpKqZkrFozJ2qFgKYjJ9jF6n6IeL/lcjV8zasdP1euU
wELz1XBMBfiCbFGjgser4PNO7jOaAjzuPKEfnQmMAiIR/3Mm6JzUSIt65vJRmdql
QB0JA1/SbK3PxNyN643+3zYQoet38v+dwsTqki52jCnN+LjaskHTO6PJ+24m6Ixl
KbxMW3VD1deDeaGfVwBy1Q2IP7nrK4zraRLtqS6/wbvI1BegeeGeQ+oWzlEBEnA2
0jKtdVvQAJ1KoB/IRoQzstKSZ1UlAfktBG2WQ+FtkaM/ag+mUwNY1F+e5d3/JzIR
LJAPjKJE/J4sq+2SZfNTamd1blY+At0bPElvhNylh8G5dG3e7YnxMnpkjTK+kcqJ
3sR1sT0x5RayEdBaolgGMT+f7pW93OLnfqQwYIvXi0oCU9jUUHg9fH3IxmKIi0jN
U95MMtqJPtH2CVCmSj+xhSFN+N/r3tTXsiR6OpChrevUgq2Lkn+Jn9QrlM/axQdp
n2gs8kOaD3lkzvYHO7LLePqArInIkAQrhsc2mynyoFYVdxbm2uFyMyrpZIACJozj
u1UuXyzlH6wH6B/MPW5r691dzK5nkJAFnfu9i90EAOookLL3Pl25A4poHefdEr36
WifL0aG31eV+ItGPqgM7nCNBUjpL5l7HZ+taLN4DVu+LMn6P1aSUnu9++maBgSGN
a5idUoxDfQeQ6Em9IvWKn7NVVrtElIGPik5dZcIlc2ivvKooO7gQBtKioMALgoFu
wOS7q714dev9V84K7U7jPM2KphThurLHLU1wxEP74YSXoJ6HPdC0OX30kBoa6grm
yEcpg3hR7mwb+Fis+dyd1RZIAKHKNJ95u9NmoJn3qArwLHm/TTV9OceNXZ30Cr+1
VjFWVCUgt5ezB+NYPdLjUwz5Dh5A+bjY22V6hPr/ipYy0VJegrarTTIGr1xDTkzG
ZzEdqXYl0MnF6qjO+kmSEJATkei+sNQC4ypJUUT3SLmGse8XuJIf5V8CUX+uHWpI
UX8oo9B++4IykaK17E2ApD6yfqvmRRr7NGFmdlKI/WxH2nmHR4/ddk0igcaJJXWb
7isetpmIotro6+UWGCIZPYQDlDgnDjCyhBYbY7R4Tt4Jte8/TnSpgcn8FgKRAsDW
36oLHUqPLCuMBAsuHkmoE+2NqW4SgcY8nTNskeyN02RAwTBqXJa/2d85iv+gstH4
XIWdAllvcXC2Wu3q7K/gpyHxqoICQJwep7Y7kRbp5LEOrlI9btSyn05a8FMnbT/k
toJGa0vUihjPz0rRIgR6gBeEB9RI+dd68kCtMzxOQlnpKYkkiPEuWATE6YY87a4M
i6SzAc0lQSXBt8PNKJy+Juw4pQjG4c9vlg4VkzOwncBtaV6VohcGSJNTraTwXHY5
nUzHk9qg58zmTSFebL+tOB39VOoKnFe0LpqqY/rjE0D9qT2CVCCUpq0o4n4ojyhV
xX0DnYCKd6gmPQcSi9ceErolhyFr1g6kITibM0Jin2nG6igpOjbEI5ch32b36lmT
sf6fMQ41rQ9byGJUG8bo/BOSYiKw+Ls7a9b2fY/NNzUohJNlyw97pHhaJGWISTYF
NElwYrWYZFur1Po7Jd3EwpuLcgp2qhFalgBfv0m+7Z5K2tafnW7Tvegk7Ydd4aAc
`protect END_PROTECTED
