`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xklbsqAgEOOmTjxdv5+oVUxEgtfGYb/2cLsop1Vh001dSEwmflN1v8NG5Tei7oI0
RuFRm3ImEM3xnHD4GAEQabPmKjnRjydLp3wPvj2oxDKfagzmUBZBgYdgv5Xsb2If
S5wN7VLVYisPbjL3/cPQjVSx0bFYNll/GZsfOXBCBksLe227j9a8DW1/94OC2+/q
l/gF8mBmy7qYprSWoeL/woHs+xSCN43+mnkewoV7rFsjPn96eAzD7ZIOJpyqtIaY
3wfPYLsZr9eGPSqkDUCmzZI5CVenzOcuCT9UiQoJyDv6kSJXjDY/9X80XBqihdI9
KDjRMRpGQLKl/0VemTgdvUzz+VAAWmWwx2KEPkNI/c19GOesRXA+WIBreR4KZj3y
HrEj8+EJgsJ/dOSnSfnNM/traAemu+PC/Uxhn+zWkjKLFT9HjrkpxcJLb9OVAEbf
7iYHQ+axY03sIcN5bzOx6D3uUJ/OidJBNs8AxWYPi2rMPEKDRWJTiCUNNVnIIBDn
E0jQN84Lcz7nX/YRCWVa7Adhjl4b+NXSBsgw+1TKIjJCd81G1ozhZ9sSRvMBc2mx
dCvWKuqoyVozDKaQmvX/nRF5HclnPWopOi2eWcoJE910SWkoPkxNPtYNB9T49H2f
DHLjXTZ3+MO6KPXZ7cFx/yKa7pgW4A6jly8f/qZScbVl3kCBmmcLAdn6v47cKXwx
NdQPUZrwyxJK9MkMC42Quc4I0ubsHV49S6MFnC5ZV5gPcDABoDM0GrWZh6JbzYHj
5DOTZzSdalpxYGpOphlpaaJWWt/JnbPUCj5eR1TrNiv2H/BdNAOcJBlGczgz4DHy
Dpc8CEykT8945roHIuW8YDez+IY5O0ar4sK7Bv4GuVc7cGGH07F0VX02KMVKKgab
1M6f+WYihL2V8S6lwSk17PLd0RmdDWcm+eMukiZNMLnM8huAEeod+2x3wD9PIpjP
xxukFo8sFDcId9p1UWCkBjxCvoZ9wAggZtCYMeu6IXQONYcLXlZ/PCv12Rbol3ka
MP3Ht+bxWyXdgneHTTxT8+GQp5P86m+dknXPSxWwY8GuEiCOwcYAnWepq/+b3kIf
HJjDJKmDU4l4SQMSy910+JOtYnLhS1OIXJhOnWONSJhiJmGYqXuCuxKMeOKCVvxg
RiTjSZ3JQdxAvcCdponsWoa4NwAnu10V2AoVrMSY7xkDQeTlbftpD/iZNy/HMIjV
yz1GCDSOGuZkpmF8whja4aLcJY6PBw3H7tjc19cigxAk5N6uj7KDThvOmSb5/b53
SX1/SS9FWMjlqya6yvFtQbD9mqWv3dfGx5VUuZuxs+h0+Z+a/2QOwexIx1PPUWAY
EXajgEAMhVPpzLGxtePhZsNF7KeI+Y4yve4KmHH1WDaoogXdEBcR7EU2JjiHQf1v
04qRntKCOhY58Sh0aN11+rKwlejr+oZBmclUGRNKnAFBti6zPu44UrzywfPGTbz1
W6iRQ+WWKvxdoe5P2XaQ5SAlaBaSMqiwEOLd8MNg52CTd2ioMk3sc7qaFBNA0bsi
tutPFORsBaSBRIcNth4Ar/5b/ukBd0+RBPBH/jeVjopafgErBTkJV1PE5UJe9h9B
JkAQbJq8Rb94WkP61jYcy7bmscIwm5COS6GSFyZk4IN6ZCT60uOoFKG1xdjtj55U
VI+CTi8eXt0mR8vYvQR4W81ad7kcsZa8lfAzqK6IvKW6q8TD4awzW3Md+afLjr5y
EugCd8DtXbXrCb9FehKl0mPz6CSqnzQjpGuIT+hPCg1Eo6+vC0Na4T7QivKTUz3P
ejrEcvyygurO3j5HGhY/nKTsnNXVRohApbOMuksd5WaaoRccV0S79Rg/Rv6xmUK4
tr/21tzjD371BB7gX3lrDg2I7hodd85iAXVn1S0qC1MlCq5LhMm8ZNKTYy30vVlL
jVukQws9XTq5Q2/HJGhGQ5F3PZE5ZNGs6PZAUn0hedyGG/y8AB4Zb3OWmP7pS3Dw
C521QpDCPYTYN4zTB6iKXG8r6iYx+7dGDk07e5fvEQ8N2fIu1/HX84YQeCm/4o3e
Al1vrnQH4P6t/PrDGsr7QIa4NowNMFOOM9KuTjxfaKkSF8IX8L33GXD0R22coiTc
8xo1YhisxJtRQJ954U9H1zpLkFY2zpbiTX+rRvUM1WFSDeS1ZuNkj4FtW33ofBLk
5aDiB2nhQopsAQsC+/OnVK1A3hhEYY9YPGoAm19fXWM7jar1hbTr4LIm7bLRIqHt
jowTxoALIAUX5sT2auBxVmE71eZ/JN3oNTtGM+doLb9RRUSkdO2+VW+KkW4H197A
L2kiNEKXi9itQC/YRGOFXosXGSYYHm08UskRv2mZa0UBfsx0T162KehPcaMnEfXn
TTR4xPBoEdvbnIN8mGrM5WOuukb84wedkM8ZZcmT57AtumgeqQtMpK0SRWZhZk3g
J+6aXpoPA0m4IGrCs+uEzvwp6QmyKlWp6kafy+xFB9x6+/kNPTlNVQxcDlkbePeI
HaE5KkOJhQbCWpEKjPl+9Z4tFEbzHLHgCV5jtmKRVC4j8Ul6BBMgLL/WVAcvaUjz
IsRRGHafEn4gvN3Cd+zr0ZTMlmt4N0MTpomTtsOlvUgptXHHlwXW47/SwK3FlWM7
KYeK3jnWDNzZnaLkhSQxeYexcMqEXI+R9PeFtatxppNd/35FH9iu/FcJoGhmX+Ut
kcoqc7kKhoRWCdHg7jq2njoYTOKHmZ7Jhg+IyP+fQ0vqlJdq/RU5tPXmGrySSsdY
525Onify+4FvlH9BJGyuoJYCASQPeD1v4gPQWFpqaxGe0ZCo8sqIT27B1uEuhvRX
OmHSjahGrnu1dwIcGc0/hTJVMBWyujr8QueUikihmhtH2ArQth2ZBQiMB0lMG0ct
RhTZQ/TM1ELu616qABFkHeEnBDZgRGKvjHfbE+dnkIKLlZgU9zLQQbC6B2cNjgBp
3K5jwBmuLoIeF2WNKJGdBEQzJMbKk4k91e4GJY3BDkj12dG0xX7CtK8F022wVn8m
24+hG/ncNmWdfm0/dVyztbX3vNiUhwjQqN+82dXAvt0wSwB4Pe8NsBP3FVuDzVo6
xnNlx0VEXsqnAbyfahnAhVxAr4RwSpRnIT/w3yUEOQRwy+xw89sOFGUMgb/Mxjk6
nByFn9b6z4mb+MddqybGoAm+6X4oiPceqX4b4pt52N9CRl/a0XwR+qdbIvgcjAcV
jQA7fdfzB2xTInzfnKWjlvt1niHCefjPEe65LEZNP1wyei0Ts7pOb5miORan8T1P
fXJlc5pTFmxJel3FJhMpecUirAvirrL/K/v5NK95XihSHwiK2VMFGczWGJKguptZ
A3Anya102dcmXWaziErPjny6dHQU7G21pWXr2ZHQ/GNtyLnNtd8k7IAq0suOYlWb
cBvxFwqinjEEGtDOHbvZi0POcJ31N4Ax6yPsnKSBtJVjSx9ML1xilZ143RQzdhq/
RCL18kIMwShsXAdgkqdXMO/d8AwwjYvXp4dSSzTnM6pEelstPinI68msOSd1OX3s
kcMj7+4DjU3aPlYYoZtet9FNAkaiT/LAeBpV0RArG0C41G3bTkKNQRoBnoujV1b3
ynB3XqcQIyv4+wRsRUUHaX0CU3ZFeQFB+GU/+JvAfd5ZgITksRythfXNbY0327wo
TMilQw15S0xag53FDM8cVgop9Jmur1hk9OdFD9svZ+FEm9BV6H/1Dx6rVDlblr3j
Z3fufhNvnG6v/WLz1WfctBbwU5i76vZuzLS7zDHBF5yTwrDGwKChGXFU50hJudbJ
E2P03abvQ9kh8bvP5MvMj1LGeg0aI5KaapqMVRMYOTwtHzIc45N/dv7KtvwKoZ86
G5/7e8TbPGo71QbwqQ7RdgqP/EdUFJppKmy5lVPNfBTIAKINL/jDiHJjw+jRziQ3
YjoSqQi5T4lFMSLaPYe1imw0fDp3657lR7fSynH/Pa8=
`protect END_PROTECTED
