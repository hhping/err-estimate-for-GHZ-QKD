library verilog;
use verilog.vl_types.all;
entity twentynm_hssi_pma_uc is
    generic(
        enable_debug_info: string  := "true";
        a_break_vector_word_addr: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        a_exception_vector_word_addr: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        a_reset_vector_word_addr: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        cal_mode        : string  := "cal_en";
        pm_uc_aux_base_addr: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        pm_uc_cal_clk_div: vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi0, Hi0);
        pm_uc_cal_clk_inv: string  := "disable_inv";
        pm_uc_cal_clk_ph: vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi1, Hi0);
        pm_uc_clkdiv_sel: string  := "div2";
        pm_uc_clksel_core: string  := "disable_core_clk";
        pm_uc_clksel_osc: string  := "cb_clkusr";
        pm_uc_core_jtg_rst_disable: string  := "disable_jtg_rst";
        pm_uc_core_sys_rst_disable: string  := "disable_core_rst";
        pm_uc_ecc_rst_disable: string  := "enable_ecc_rst";
        pm_uc_engg_opt  : string  := "reserved";
        pm_uc_family_device_info: vl_logic_vector(0 to 23) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        pm_uc_hssi_base_addr: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        pm_uc_pcs_dft_out: vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        pm_uc_pcs_dft_sel: string  := "disable_pcs_dft";
        pm_uc_pcs_rd_lat: vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        pm_uc_pcs_slave_count: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        pm_uc_ram       : vl_logic_vector(0 to 37) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        pm_uc_rmw_dis   : string  := "enable_rmw";
        pm_uc_soft_nios : string  := "disable_soft";
        pm_uc_sys_enable: string  := "enable_sys";
        pmu_cal_bin_fname: string  := "nf_hssi_cal_v10.hex'";
        pmu_qparam_fname: string  := "nf_qparam_nf1.hex'";
        powerdown_mode  : string  := "powerdown";
        silicon_rev     : string  := "20nm5es";
        sup_mode        : string  := "user_mode"
    );
    port(
        cb_clkusr       : in     vl_logic;
        cb_intosc       : in     vl_logic;
        core_avl_clk    : in     vl_logic;
        core_avl_readdata: in     vl_logic_vector(31 downto 0);
        core_avl_readdatavalid: in     vl_logic;
        core_avl_rst_n  : in     vl_logic;
        core_avl_waitrequest: in     vl_logic;
        core_interrupt_in: in     vl_logic_vector(7 downto 0);
        core_uc_rst_n   : in     vl_logic;
        dbg_dfx_clk     : in     vl_logic;
        dbg_dfx_sel     : in     vl_logic_vector(3 downto 0);
        dbg_jtg_cdr     : in     vl_logic;
        dbg_jtg_ir_in   : in     vl_logic_vector(1 downto 0);
        dbg_jtg_rti     : in     vl_logic;
        dbg_jtg_sdr     : in     vl_logic;
        dbg_jtg_tck     : in     vl_logic;
        dbg_jtg_tdi     : in     vl_logic;
        dbg_jtg_udr     : in     vl_logic;
        dbg_jtg_uir     : in     vl_logic;
        dft_clk         : in     vl_logic_vector(3 downto 0);
        partial_reconfig: in     vl_logic;
        soft_nios_addr  : in     vl_logic_vector(19 downto 0);
        soft_nios_clk   : in     vl_logic;
        soft_nios_read  : in     vl_logic;
        soft_nios_write : in     vl_logic;
        soft_nios_writedata: in     vl_logic_vector(7 downto 0);
        core_avl_addr   : out    vl_logic_vector(15 downto 0);
        core_avl_burstcount: out    vl_logic;
        core_avl_byteenable: out    vl_logic_vector(3 downto 0);
        core_avl_debugaccess: out    vl_logic;
        core_avl_read   : out    vl_logic;
        core_avl_write  : out    vl_logic;
        core_avl_writedata: out    vl_logic_vector(31 downto 0);
        core_interrupt_out: out    vl_logic_vector(7 downto 0);
        dbg_dfx_out     : out    vl_logic_vector(15 downto 0);
        dbg_jtg_ir_out  : out    vl_logic_vector(1 downto 0);
        dbg_jtg_tdo     : out    vl_logic;
        dft_flag_down   : out    vl_logic;
        dft_flag_up     : out    vl_logic;
        soft_nios_readdata: out    vl_logic_vector(7 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of enable_debug_info : constant is 1;
    attribute mti_svvh_generic_type of a_break_vector_word_addr : constant is 1;
    attribute mti_svvh_generic_type of a_exception_vector_word_addr : constant is 1;
    attribute mti_svvh_generic_type of a_reset_vector_word_addr : constant is 1;
    attribute mti_svvh_generic_type of cal_mode : constant is 1;
    attribute mti_svvh_generic_type of pm_uc_aux_base_addr : constant is 1;
    attribute mti_svvh_generic_type of pm_uc_cal_clk_div : constant is 1;
    attribute mti_svvh_generic_type of pm_uc_cal_clk_inv : constant is 1;
    attribute mti_svvh_generic_type of pm_uc_cal_clk_ph : constant is 1;
    attribute mti_svvh_generic_type of pm_uc_clkdiv_sel : constant is 1;
    attribute mti_svvh_generic_type of pm_uc_clksel_core : constant is 1;
    attribute mti_svvh_generic_type of pm_uc_clksel_osc : constant is 1;
    attribute mti_svvh_generic_type of pm_uc_core_jtg_rst_disable : constant is 1;
    attribute mti_svvh_generic_type of pm_uc_core_sys_rst_disable : constant is 1;
    attribute mti_svvh_generic_type of pm_uc_ecc_rst_disable : constant is 1;
    attribute mti_svvh_generic_type of pm_uc_engg_opt : constant is 1;
    attribute mti_svvh_generic_type of pm_uc_family_device_info : constant is 1;
    attribute mti_svvh_generic_type of pm_uc_hssi_base_addr : constant is 1;
    attribute mti_svvh_generic_type of pm_uc_pcs_dft_out : constant is 1;
    attribute mti_svvh_generic_type of pm_uc_pcs_dft_sel : constant is 1;
    attribute mti_svvh_generic_type of pm_uc_pcs_rd_lat : constant is 1;
    attribute mti_svvh_generic_type of pm_uc_pcs_slave_count : constant is 1;
    attribute mti_svvh_generic_type of pm_uc_ram : constant is 1;
    attribute mti_svvh_generic_type of pm_uc_rmw_dis : constant is 1;
    attribute mti_svvh_generic_type of pm_uc_soft_nios : constant is 1;
    attribute mti_svvh_generic_type of pm_uc_sys_enable : constant is 1;
    attribute mti_svvh_generic_type of pmu_cal_bin_fname : constant is 1;
    attribute mti_svvh_generic_type of pmu_qparam_fname : constant is 1;
    attribute mti_svvh_generic_type of powerdown_mode : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
    attribute mti_svvh_generic_type of sup_mode : constant is 1;
end twentynm_hssi_pma_uc;
