`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fzDKyAIkQ03r3xrvfh2YKo4HEB27NbAoqtnMgKnJ+K+Ym9NfzU5IlhszMaFNZG3L
9xBvGTyuY3Xpo06O3G70End8Pe/LzYbWPFYGvhP22MqvaNlKXzp3ICtgrAcWbVfg
4LAM4a3AUFAPSbaX8/G5xqisb4ksheEXnksNO2R3WbMSOsAZ/SwUohhdn3rc7enO
XasNQkuIC1iRws9CVuSKhpW5cHIMa5VTTJd0mV5TUM4UvhWPtNQAzk3Jcg90gDge
8icCgrx+pq1A9gBdwowoiTlRxWFked8cgvPuofwrR8954HJRjXZY1RI8GxKv8udH
j2E+XS3oQLB6joCnK2w0jO3J4W7FVFTw5/SaroMSdqNPkYMcA1Rh6ITYhuUuez6B
ZrQLVi9ECLaJiAHbBYDrYrj4L5/2qBXOhlPbx2NF26jrv7NW99Djqo+9wao1s3v9
nH/Np350l3XWqbSkTZvtwQyl1BDkWdRkJW7y+XQQCe/tc09hgWFhngvzbnnoMfgE
9oe3+ptxcof02ZDwy5QBFQ==
`protect END_PROTECTED
