`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7HOxPUBcya5ozUfXmZtS2ivI0ykqCNrv4daQJPIq1g6UwAil8OLRxt4dmTseunUp
JtTb5OLAAQq8iuovjtVp3YQrXCRVNHAtk4ikjIIu+NV0oiR8TMV2lk7bcRu36Frb
IVYc2TY6hx+sAQEthhexi75BKSA9BhE9iC3M1lg4oGo3c/XlQRkn5C7H/Tcjic5f
ZTJL1g0qb6OVeT1hTyHIfXLWbevWjCXJZ2e8MtsYCKdEoBfo/rMiW5+jfQ6RJ/VH
tyR/XlFHytPiIxDRRcbTnkaOL2T4foXYhlZ+XWxO1oHNWbdE3bZMYP/r101HAyeL
LnVM27cxoppmJMZHXGCvaCIoNfoJnWt2x9G8Ywb2cD6VZ2EDWh1uFc8+5S3hlKuA
gSXIXoljUc1HbcOhL7bTyu5Zn/Dx1Ujhq+etbDTack2Zm/7xJkOhvpFsYg1RJiz8
WHQh3iQvKlJ39PZ7JQ0HE3e3SiOFiAp363BmK1VUYxcI8PJ9w7V+RDUVkndXSWIS
5+D/kPUWnSG1fJVXu3YYcJiLHj7PTbxmpg4FXYXetA9m1KVRni5QSZLkul5Tpj4a
GBMWxmdxIz1MTJjIp3bour4buvpyE9oXwrWlYwoVPknkkdVfPdcikzxvcMcQiazJ
S/QX/TcSdspP4sc/R57R2YFFmEnl8XoUM3vQPWV+iBfMNrqCXkQ0ICn3/dhu6bDZ
k0pUIcjtWkM/hzo8YA57NF72cokr0Sfa/bvLa3owWYtqbThbmMzjhXfXOPz3zV73
n/A+uOUuZlsnVJME5Tk4zHfmavEvBlzJD/DpFTV2xOyl3gZYrhhJyEpz1eGt/qo8
Pb1pBRU3gHI53BWBVSVYgGpPjH93iqQPdg6kyOiSHPv+KMbaaUZUacJD07O5rQKL
2xTJA0iZ77/FNQFiNOKhqJupQB1fTs8rKe9kvVyBNZEKoj+u86jmBAbCTGQvb4eZ
ISoio984vVSwvjGLiM50Jp9mo+iomi8ofqlOekjjjy42P6CVaZpkdW7k3hGtNAyG
aeA6DLIiUXrSAC6H0j1yjETJuJXzWaBsk5JRigQ1xE6a0gP+G2L3bItldwnQKmBB
525k3mLYpt09Ewv/jCE+PI2xqVr2A68CZQb3hpAL770=
`protect END_PROTECTED
