`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vlhNagMHJIOW/rhk4wU5OOxfSTPiWDYn8wxvA60+Yaeu0p/GGcMFThSPL7MSymMT
52nSSRAkHWFfr0V7uQ1vgaJVq15jsMepyK54asXt2sZ5nHHCvw2mUxxwHIqbd3se
Gt+H2a0NW4R+qRBnx0IMHp0koWuFWQA+VvrVXSnP2qTA7hhvtxKdE9F5kj3AWTZX
pkoWHSYNTcmGu5fD95vI9hEwGh8K3m6FU/X2nq7aU0QY1IiEElPH0Q+ctVhOPgUx
x8R6PkP9JQPe/e/feg/c7WVt3Qyu02cdxddTRG1BzOEIaQbEqYxNdQQa7K4Hpzki
TJO7T0BxNzubamjtWwcxIoJn2AJJd4pdPDxEKH+gcT+z79rJN2uWc+jGyFOHfeBy
S++S/YlbJU1g7qq08WqGf9ErUGRJVpb6dQVkU7T84d6xLnCVbWU2zTK11HPFsjEk
NCsgtj8nJ51MvJC3p+6oT3yFYQ4Qirz8r3t2PekwM0Mxdzlrr2IX5KMqFKh6sDD3
c1u5+ttmF8MDcT0z0ggK47PCaaOW0JYzSoA+LI3lAISXirCNqQL55LpzxkPH8VDB
wzEM0kgXvq8IMdcIX7tdUz3r0JD9hIapAPQiSfZH/HDKRvWWFkUFnz0ug8mKYKOk
E3oCVMdsPibUwPif9Kqc0cctMAuSg40cGwIlCInhrJsyQafa3qr6/VjygQfEsUqf
xInXrjPJuFRchMN/IzPh23pMPBi8uz9S6Oo0AskKjfZ7c+dDNp70+IsfT1RhHjvK
6ON5Jns2YZmXhYezc70az5tXwrmMfmeGt22RRNWu8V77n+4WLQsCUVT0dQo1UHuj
oQrZkSd/IopHnVK/aZRVksF9iYaDb2s+WHwpuUcrVITVVBm22D65PXvYZOWDLT6R
AQVMUixPzeIXtlhuzALfJ98weSn2C4GZlRizZGPG2JSm0ms2tlES4CWSnZmH4tXI
lWvxaioUfv/xYi5ehh+ntne5pQ7U84Soo2Zj9AOKKM/ASOpkcljNPb3dkEqRt0NQ
4EH96nffy8l71b5UtmGXS/wvghtpVtUIDLac0pqO0DsZjWyX0cYn5K8Hb5sQX5h2
tFKOV0oNGO9ufraM+7ykZWM1fwJDlXlw09AMkcfCGmKuf+OCanyZaD2pD0PmoJDR
tQ6TFsWVoh0GRaGj7nj4OrYuzahRfyH5xfEu7e7XQ06ZnB0RiytJB+rXGIMkQuFD
7UQ6SF30tRizSVwpm7khIMMl83TF8K+c0YLx7c5Eyjk4LRHzmMIbLdW4qU2cwNFl
DXZgp2dAuLV6dw2+LL7Mnm+rrgKPSBOBykkG6R4DI6ujc44cAP0zvftCTk+pt0yA
B+I2S5xTuiDybPWz8wjCSAg4SQa8HimDc/BGGtKpuA6k2+dpSKhLYtPRsXCQ1uVI
Nw8kedszWP/KiaWqB7099nwesaLZI43TkK1NsuYVZoNB7nZfQW77UeFhmM/wLoHj
BT30xehmIcF8ntfoCkwlrBVU+IOce7r6QPPWNUENISmstRafeqH82WKqCLWdTsoF
wBOchf4wHzG47BxKaGLTBRUcLUEfDTcHydkv7bWZ6SSVajsxOx6mFlzpc8OIluuG
cKHaNIHviWQRgm91lJVxRSYgIBUyXiEQghNP5OPpBE1MEvvv4cTYpRxYuU9yqiCD
4AhggisMt+uxDVW7kkbvGCj4RskwY5PGUlNsODCnltrTqWd3KLUW4iELQ3He487f
uISHHO9vFFW+/4T2/cInKyXd3MeKPj1GM3kl/mBLsDfs3PvdulJOoRpGOT2SdkxH
HZ6+mPrPBmgy5CKZESNt4tEp/HHfSXbT3B9issUozpcifGMNPjg93MTUc7EF5c4g
wsGgog8Qve3/VO9tnVUUDjGcYmieJi1qNVDHni/kInz8aZ5BJ32IeLycYzco29DJ
MfdCr1+tkSeseHNn92uyLl7KERHD6n0tcWqQ8z+2sWoHktY7g9PKTGxfdOtb7c8W
HSKZ6xvd1+lD76aVpVXwPJPxm/ofKl6NgCWwGtV6+yg9GACC5CwNz5N042cn2PYj
6cDy3HWL93BtrXpsM98jmINYBa6hWfsOKK5gVfv3RBa3mFLMntkLFM7SkTws1XOk
rBz3D7T35Eg0vNH08VKp+uNHMMpBKTHVUoSqP9f06GMUA6jGNjQoBBEtqEcfV/ez
ZT7Zt8wDO39DJH5U/xhNcSJpdWkxIXmRM7jD6FVw1z3myOG2GNuSp37aT1QvdR8K
ck+6trR96Rf9Wd4i/2/gn3ssVuFq356EYV1U4r0Kmbthm7+rO9lxCX4crSoFJhGO
yyE4tBCoCnW19UTb6sGazgkOV2UeQGPIhzU033BcMB057LEKaCNmNlaSpYoq7NPA
xKFnwlh6pwp41qXpThWf5jCADB/40wMa24e5BY/bq8b+NI2z5VFKSbM06pGbQN44
Bv5cm1bC0uKi+7X/BbRc6kNHLrWd7qXo2odn+JqWoZUOlQFXTA5UW5M9seyZUaGC
qXuXySZ9BhZJk2I3KWzrCsS6KuTihRTDTWUUsYn4XiNzSWSNXOG4OJGr0GSRJVFP
KmjUcyPM4+DoX4ortOtECLMNx+5azaw9nIgbRc2g0+Fs0OLoPWRtwUtPRlwyr0Hi
7Wm3t4Jmc8ycQXCdfkii1ABpUw6gXbPyCpDvvjhiovOU1H32jjpa+En4eq1RhURu
OmmEhVuIlT+Zi0Gqxhvw4PH0y2TM9HZJncPBughDr7/3X4fsq1gDamALJE9Cfdn3
ZPknWFmpJCRqgE2fS8NtuzBCQlmjv2gPx9FBmMoKaIAFNzdk1QOyLjijiP21VJqG
TMdQBCPk0r+MusEHnqdYgzmUF/CTvURyt9BCGGlFl/JkNhBOLngPp43BQM1cXnJ3
Je2lflGeUTJNhUTIn9+GkIqOY656OdYqL5a8r66Go65d+EGenKE2D8174o5VNE/H
/NExopErOYl2bMdU0LMM8/ihtw9EpwSHT51YMPakqBs/2cBh5UaeDXf2z7S8up5o
DsaKYuVz79Iq2pqWRX7XBSUmooVLJ0R+96meYULj8I57ulVyzCDfEdjzGysyrvV9
rlil72nGB5GG6DtRpzAJIqhNPfo9ZPKdVxKgoa/mlLBCDSiqs7Avg9EqIJBwCZ1D
V0mtt/eZQ9ZFOBGeTE/ovyWQpMli54s6zvJ0s0WticJs7wdYdRjhLpNpdMeaRSTj
OuUqIdlpSMdQYzRpIU65keAQhRow1wvBEEFBdCnTKkzitt3x7Ic4GVrILnB1//AF
7NU6KhArl4WRFJe6ZsuMBVNOrzfGgTDCoUhTChWb6hkQS3lqmvrO7s671/KJmf2k
7UyOxeEd45idNbuuU3P5kfboJJwfO8Udix0UMHEMxP5/nj/sPcYrp6oD6jueN7I9
uk/fyWOJrrYzHpnclD4wXPr0PeKYz6HyAIQEpktvUTz0QGmsNR4/Fj7xmk5rd/7l
wQXD5CRhmqiWvOmQLZTYgbLhp5Cz/zKGjF6MPZ/weLRaarQtgi9cJxU6zKR4PEQR
/oPM+I+dvOWJKMQKBUFBjY+2EiE862LAWRddPTAq/wabU3WJVclgmq/5XxJLnitc
FsD4/FZ2LQa2eoRhNAyGe6wQFas5YBnmc0qgPbf67pGJ89kSovHYbcTxxJ4TbFVB
XCfixFbWdrnl31vTd+h7AIfUqoel312LxKX8LjWjkc21Fu7ujKyVQCQvwRhO5dF+
3POmQhEoCdrml58olKCp/hQK0tAYHVfbEhDr45/1S0O342KCRSXu1HRcCQEayPWJ
QOKOSot1jDLNfSSrc33J1WwV+7AKijEyoPjvWe9HWaSf1WusOnU1VKX6NsG406U1
GhxSQ6Gxo/rJV9QfjPFmOrxVAlzvzxr2w/583yuu9PcOGQbR/9u2/S8+H7FMr9wd
zAdV/gAOKohCjbiQheU2Hv1r9lnQSWi7Aa1HKgFSKXWvTumYxNZWy1AKERthyHe2
lIzYdXVKUkBIokbqhjHieY5H3+7CSCMEeC+u9kVveGtcg5GuAkIIBcf0t92hllKv
MMW8MqqUSXA6lD9y0kDb270vP+MBzfjt1sA/pBWPmap/sL++1AqwjdEumaeCPPyc
GXE49GJtOOMjHqDXFTqwZcaOfI/FLasI+VMp3axiJrzf6mRpBzlwbafn2xhBFbto
1lFsMWqe8NOS4S1efuM3INyXFy1XZUfXjVZiQtkA/9gSAXnULEAbth/S6ih2igVq
KQ5rTa1V4dgK+FQDp6hH3k7X9yIbJq2tnhwje5vjL1pShPF7aT2pDnntfmeYq3/9
7t+j9ai0BzT9mqhg1qXXZDoI3g0Qx4OjPN2BqhxXuUBkekwkGf28T0QWDGlvItoI
EevH2SFjTNTPQwmOw0Uj0PJzsX7IbvDZ+FmqCeLKbB8NPD8IJnXPk8nfeuf4I1Ws
uaNBPPhewDSDhhRG2ccJ+vJU9l65UL+U/Nxt/hh1ZMHad0MCTLbKzluMKaLgYD4w
SfNcj4pBXBzU5IVlUho4J+8YuvmsKcTSbs2eKNLhyaiZnX1xUVfG54l1IABNXJKG
Kozjob1KC0qbitJUr30VytZIrWz0YnBh2+oQZw1rDLb2PKCaXQfzzUzqrVCMBNUl
TzgFqSn3brGgQrsg8zyLPR6P298rT9IgXNwgsZaVenG/gGjfkLs+/kcfVIqk+ZHt
UFPJ5s2dtXQf69Z5HXmSoP0R47fmRFcjtBkj9LYFw2GomWy85AHvMiFSMBrNY6gq
Ufy8S1MwtkJOX6/SSqUB+lA0WBpzsuGOnhND+RZiNZYgXpzZs0cy2w6YvOy2GF1E
RKs2m6vhP5LVH7cY58f/cWqBjXWBIAdBB5qRAsKof4DzjgMZOJ6GhahHWXbgMWqa
3gcuqvzQ3Gpz7lv+blUJ0AfcDobvcQ7Y+Kkuj6kvZ40QAapnPCDXzbHt9AnVxeE3
/3YpCtwNacCLxYpPal89a1Jbtdut92uCjy4HEaxfhvLT4iIfDnftAnTbVBNKbBpy
RrItv/EH4xIRDMzUBIR555fvI27BXVAlP7Z9tUTEwXAqm9iw3IuUdwjHNIGLHXM2
DhIym5U5oVVZtDvbv70YOayLv1g8tNnLNg6ehjZBDLiknJH/H5mzRYNBxeGZL/AX
74IUIEThWN93Kd2JQZPlx1cWgObBr0hBBfmiTYVF6HZZ4475s5iyNDyxC4wGBPgz
jHQm+FwQXETZSQs7rZv1d7tG151oRPdn3PoyKfhx+ZDEia4HtfqhlOh2x2B0PHF3
85lQHtkIvEpOfcOLfSm0J8RAQKpQb703I5a140pM0SU1asDjNDJ5hLpQlR5xAO2L
kQKvSD61/zgTapmy0E6zs98dBuGiZ1Zk1eTQpc8sfjttaJbYCloiQCqy8IjFUnTY
s9jIcza7dT6rOgNDmdSB5j23sMgI/WX/UwQJvHDj1mFgl6UfZtuTJqQh7T/xfD4g
5SPcqE+VRq1ZzbKnJXbI5scj7/LEiHMiQi2u/a7X/BX2DFbkSFatgOBeNAvkyCYO
N/pQfzTTw/v7ullqSfCr/YxxTMbKBRzNftt9mOhC0GA3TgCsp3eWa6pDcB+yXPMR
p2wh+NaQCWvvnbxDgPI9pKbIE7GyZGYENuMayl5iiRard47vqJ4/yxsL6k33UAqs
PDSmwVGJXP/0r4saWxdcMP3o0njcU+hyouQWFs2J2c4LHNpGv8xZPn9VqWZ8ifIb
l0bnD78So6occPX5OFhQ48B3G6k9btBB9qx0YnFC4ogSUGX9WWv47G23kzFMDtuq
LAkLvDFtQg+dXSs90d69bynPMkQ3D/dbv2JSr6RR6YARh3crXSjY0I2VV5oaA33g
jTqwlyR2fwg8AZ8V7YKsvYqkzvVA1aOg1rUoJ0VMRL2P0K+1WFS8EHRcGDMvU6Gh
fJSiHwKbc3jXkvXFogfysVXVjwSDkCIjiKqjCOvUtL828SJDdvhNwd4mfT3drsW2
5nEjU6hGvDx7AKZj48TBw3/oHJtgnji35iO70syCthEpc+1CHn+xXVWxEYPyfvxo
Eo5TODy7yabMzp4GnvKua4CxSqNG0QnuUyAc+n4f8YNc5ekwtUlut9wL5GcXwwzh
SH0vRfo5RWLLP/FKG2zvp2dV6f3YwreapMzFenOGkSF/YWG6sf32HL06/lHzwYff
QhuhgSf/Y+NP7Chlsun6LC6LjojzbEw28SD6Vg9hCUe9Z8EFaGKOz9Zn8LMKfW/s
nOCb5ih/qIM8LvqZwvXIEzwiYWVoguCBZ4L3Qz70dbULr1wFvWmcMzX4VMluRa/S
OZRVICCnvEVKj86kkwUUWtR2Vo4ySal3UJkM4238gcT4qG9/QyEZvlLhyrtoRyb5
oaUvQHzoAXaXKf8CsrAIj+AorfsOyQWICq7jL514OLtUFCG5ALqn1N2vKP+sg4Jp
FJUPOzDahxVAw4AzlK7lnzJ2dPV/FpbwSXBj2fRD2SxdXGCsu/8ZC++p4/pPzBgH
Gsoo4+hi41pHs7Dy2uJPtlmbBl4fZouBSfieHj/Caoc3fZ17x9snPYROPOmfIegU
0V3Sv39tr5tXtPKgCF3XoN87KSRowC27MjwPi5Q47SYOqg4ed66Z1bZmleJ6DQit
PJ8uL090y71HFf3robcsjDZ2cFgHZa1lkOfasVAMPXmU7Em0Mq3dRn5X+7GFG9gM
8w3tixHkV2xRnE9JRT+tK7nvZCVXJZ7HzfwhRHnc8EiWqXvX9Mu40N9CiNcRyLtq
JbUJmgf1FoLErMV6yWpaSjs0gFUE7WmsnUEQYMbFY8GbxvZrDH0h5VMD/klSacta
5wsP0pkyhTq16dXbGbX0hrfGljPZ1R1CYQd7oSI1Mnw9Ie68ToxzQb4eYmIkvohm
Ciahe4gN9rTTKZs/ln25aPZ2RdIwdKcF8KEOsOwwr/vosrc/CmPHRqy93uXS3j4D
Z3+9gEZab/vQFGRsQQbCzsPHRAroAT4sheXa8ojj1nlSseKzYCdZmMPRL6QGU5xa
Yq316H0YceeeNMMraariZaIV2wKqD49FQXAB8nzQacJyFMpHGwBkL/otPRwo9M/3
7UVhq9JwrTKCCKfFnCWVzqU/sjbwv5LDmLmGPQt3vYLRXuRFka3rkGEKDpscu4of
L3QHaBu/B3XNmyS/f3hMPIR6hUOce3LVjSTB98B1fXYny0Mm8QtoUCZd10Xn6vVa
fUyBrfINonmbW5+2SYwHPKiOJv+Q2okMhuTf+0BQaSPGpTzw4Ajyr4LLyRlG+SEJ
/2k+x46fa4PWGutRKGUKNbtrQXAu1HzKpqY1GqDmwYw8ZfBTvopIZYClGBpc3GNb
YvwDvkzDgjr2giSENiF0Vxt0RzcxkMmr6FtRIfcOBktOTsX9165SqeBjSjToLpD+
RYQz1MQbtM477ap/yxD4tuqHccIVcmyx0akLzCcl+QAGN9HpAZONnnVDp799ARxM
B//2dD2meHWDqyVsHZ3zlQLZw3b3JK1gEwc2sS1y6YXUCHlt6H4dtgcIIC0NlIvj
F4VUGiXvTmUTDI7YBiuQDpgLsKG1L+IvK+3LZg00iy3uYhlTIYA2YWgpXs61Zsxo
+Z1vg5iHz+J9jzruvOfRY4b0pLazAuF6RQNblW/DiD4c903bxyJ7D8YHMkS+UadX
Eej+lvni8MYvaQUDifCtVUR305Mc4epGKWpccAK+Mch+PdDU+T8RaHmmFgkzNRlP
aMy8D0nv72pJDRViXyTJndOt5VI6x4sIHhSrtXFxcBloAYAmzfLjDMuakQDWYrTL
QDTIJ8BWUNYOsqbuB6yA4lg/qBeeIro12+TLnkIWNQ/UooEKnmF4/VJ9Yxz2pmc+
zZofDrajm7Zq0ekMvW6y+DLqKldNASMJEPHap9UAWLQq60hMPJ+ObO0HO/nF9q1F
SXZ1YeIAGhcerb0b1UBbIWKnP8BhIzUdzCoSDjUMD6h1aEpAkdbeDTm/Mul3nXYS
A6lpxkdkmgiTS63G3Vi5k2nnJb5rXXbC0F3gqG8BQ0ksmp7crpyz0xZItQkEQnO5
BzsOTMl05uEuORCLuMdUSQVM5NKpKJQ9zF6BcjrN3qX+GCyT9LNyfkk6Kqa+OkhV
+wo1DPSA2xSS5o7vJnNFvGc2O8+YiX+yqILybR94KvGBCo52WCTHmETGWHdVyEyR
KPKC8W1pzfRqdNeETgKa/QETlJjEbErpHSr70t5Dt+V9F0lyXBw+M6hfB9nc0wfo
l8PUxVftPYPixUTx6dUjVfXky/+jyxvbgNzqjTwYKvfs1Tf5eqd0OUue4jPFgm1Y
b6GRiZaMXgVn44gk2mz//WEimwuDlAy5wGJPz8a6rsN02BM6DksiWEZFJG8End6C
b1KwOnUDZ3GJCihe9qBbtjgNqBhvOkiuQWdv1RLkQqSTCLWXw0QeNQxfZpAOv8+4
0X5vfrdipiTu4yx3JuzqU8xkunFjF59ZOTxanWF7SndoPNCqGGyd63AD4OixY1Un
6K4kUAlEwVOCx0c9Ekdisa7Ip0RuAr4Uw26aLQA0ZXrejnSwk9XXLYSLDs6OJZdC
QUbqsHePtx3ZH0gtAcMlw7Ga1XT5JzVo/ZhjgxeLj4q4O1CQbavceYUIQMpl1V/s
rFuMEGApV+cmmCQjREuI6kQvg93IDkCDlmVKgkBs/zWOY7nC4zcZLiO6LOQF+W/R
103P+61qlmEDubRsfsUjaPNSsw9EbX8fSQpfHd1A8p9rVcsIRWcLCXC+2AnRf99Z
FfJHpzXLBWB1lthWwoIEGoz2fH4hmeOBKxoJHnlHyhBzzYGQnWWwP591IrlEI2cb
l+74zgpK81Ciab2yPwCdt81C6i6gZfVStT5oxfTE0E01tddmYROdTJg/b6R1DjXI
KX5Aeua2AOiSpkvQnvas2IU7tKDt10wwbanjOgSMsvmV4lI77slin2raH1cAIm71
flr1NjkI1X0qG4UoAIkQubyT+cV/1YKq7EbT3kgyFMY12zT0Ra3DvfkiJTxsxaug
sfZk9fzA90ipAgNuUGGVd2RV3BRyDdyMNq3jw39qRMWEnQ7HT1A4OeYeyNx34znV
OKboAZqFYeA4qRN7oLEEkHWkfOOPXCCPU6fdMWiL39K7/iQTGheqoucpIBpUTC/4
0u1PTjX8QhoD1FpS/paLnxSsZTs3UJljG7Sh+C0BJZsUGG1JCZ66b9VRHFlnW3Gw
TSMRPeUA13rleAy7SaozeYuG51I5ziy2fbY5f9rSF5bVv6QidlYQ3Gp5L5jybRab
JqRUy3mj5zR6V+GpZcMI6Pu+CgAp2GRlyoPuq65yOqxGyTgBjM696q7m+gdT75iQ
OK1TtrlS0WNM/CG7x7KfzWD7bBPqQv/5Y8fPKqmzDAzu7IQERhs9sfr4u2Gghsdb
OOmrdn2ty0MNSynfzZkgV/qRQ62VCoLJR6vZ5at+duWRBCUc1v52kATHSn8LRSiE
/hDadI8S9urCDiRNFvvlpfb/6euTbmo+gJxfZMkmjZhN/BQ7En0cATljaj82CazH
BQYiv+R0HhV9ok/ZfH8oZkCriubEHa9l0nRGC6vnVbsVoo6CLBTHd1yqNk8NjxNQ
rUf5FH+7iQEJUNc8e4qv74JHPFw3Z0+4lD+MxGqPF5vmKuTZ4ARlr7Cmd8MR5Qmq
kGstCRmkol71OVh58hLv4+j7Ih4rPNLRDUBnBIRscz7PttxWMGKYaeMTMtCmGsut
7SYSe0NpmnliIre5IAN9m4ERJNgzBSacfpohd4ierKlunBPHAdxU6MREOn1TRarH
WQ6KefU8uCHWvit8j6T4JGq+2aphrXCnO1w0Xz++1SxXBc0H4szCPmS3TD2bR4QK
othqdLAPg1Z81AwVAWfD7sAV0XJw2TTz95dsrVEAAum1g7GlJ142RYDeT9Yf28Jf
k+oY/vw8oiW5nrqG3BWtL4hyRb9rpDPNdMutiNO62pInybedPO/bpe/VsZ7m9m0h
x+Ti6dOm2OrLYLKfmDzV2CXOPtRfnC14LHVTp+Z68gHylaaQbosi08JD3SGrOBmd
F7DHmuGOh51cofSFPEV9Fh+EJ2RCqY6VDqMkarElluJtEHpm7cRUz+IQ99xxncKz
QmpvoEEM8xeRz9TgXSK8RWDBO9nFIgkR9E/d6UOhxfQDfYNJk8LXOnYe+JKCrHoo
DFRq9WckRWJ5HOG6nLspQ9VxtNxHfxym0ZClV3CkDGCjg9ExA0BO1BSN/X8i+CtG
sirKtiiNcuF5TO2i4Fj+EOL6sXVCpnd18RlJT4Hzo+vSEj+0LFU6wXuoWJce44EW
KQjADWwpIFgdibZqdxagPRemdwMiZEz9cg1iTQmlRZxmloQ0fIoOGtX3BMnMtGNv
yKP2o2t5FSIhtCNjY8ULjMrEi/Ou6fY9//xQQk0KdbhI/T3BHFcueDWJNHiC36ZF
4kHxxnwLG7VDF+y3IYxcxVvWgj9hxZcDoBDzgv1b6uh7MPxDzdyPFzMfLxkqo4SL
3AkWKId9S/IhRBTP6yMMBUmpyRbcHhso4BKCa+MeyaRwzDoidwcHnMdUrG3JbG6f
1tyoA0uCyqAu2ptOETqh5tKB7KHqTb45lHRu0tQ/VRLnMRA7bdqjzSKUenciTQKm
+d38x4btsQbmoMfEFZMVc4P0M8iBKDeIrw8mDSOMh+sQ9eWoNW5LzvkKKG99TMHs
dKvcvb9ZFAzr2lxipWhAR0Md+/3HwKowFruXzn+qD8CuHmNMPIVEVQ5NyOarGPWZ
WnmnGa2dFJPD3UccHeVKoN0e24OgEw1FQ61AnfxM0py8S+8c3A0849OYxrLmsXCe
+kIdEDYrj41pH44XXBvFXC2jMFwt6SxN4fwi48S34zQ3RCA3ZECuq9yJ0nEtPfMK
t9ub2CDreczApyQYNMQSFCvz3M+BG43QPDTudANDF7N9X6Gi+hmTZphuIIfl08ng
VHk+FIZTc2RNOOEVQYUiKfo+0D5LDYY0hOC8i0I4d5JDAckSacJCzB8GuJtbowcA
/jAEVIZjGBYQitOZi8TTzVAgYG0O6qyY9+t6n74uXq4ZUD63NKhDTzUqFHucsJIT
0wbhgR8VjthRQu/q0eubD0VULo4pQh7AiYjrnG6JZqwC+RooqMsa0JkjOy5GkkeG
LViPRIdt0F2uCvjRAYs02f4RLtY0uPUA6IqoXXwBp1lmXPJUpKxlE4K2WkdtZ0NC
WDsBYNqyG85UR+eRs6wA4kjYLiNJ9hxt1NGKERRBmtU87b2W223rynzPfxPCGB3w
AQBoBt2E/qJIveIiZuOwK051UDCKuCePzJ7CDHVxu94HOEbOo8Es9PxFS2Qjihj6
uQq7JFxJqLfo03uefVFud1aenZyvAsbapJTtg/VO3v1FQFwzNmhOV+f01eaIQLIH
Wny97h42BNSq8yZiUZL0fFaesNUSE61apa/EVuJbNZmCY0WR56s6BHNeLAJvrS1a
1f0Y3maatCXo6O9HyPzoWO8PZrkc221LYgruvDBhW9aymgmtMm/8H6ydFaHnNi10
A02fKBMYom8jBTyUuTkpcm9tyEvP+pfukmfq6hBdBLpKcJ4ycDQF1zGe1b9XHRbo
ya7SMG9vRqgZPFukIuOS4ICDt6G9o/LbGW94HVx1T5fWly/wjoSkbU4DO/xzOhhT
VfP/soHnEFsTMpKIChUT+xs2hGxfTJ5YAeuyPmd9ZECSJ6bjf2c+LzEA7H20TMwF
GJQU8I+IhHQQ1fqJgr6xqDuAc9GGORkZFa1jJBk31mv/5wh808E/9heRu4aRIMnM
heATs1ElHof0SWLQ9Qm1tN8efa6z8XD3uq2vEtTlzQtRje8t0SuycVVqnqQVeDOp
R3tyNfwLHM9xjqT+9/gbjF8A7v7OGGHd8OhR3u2hR11Pcbcmc1OkpjuM1DI8eyNo
mjYTh0YXBauCQyDpNHfycRaJKS+9E0CerIYcu/WY+blOvGuCFNOTwJaW2ZXGGhgz
GaVk4tGQrQmzq7Nxx7c6Q4b0SW1/gtCy5evxVRg0lO+OHQrNIZGle7iL1hTesTx/
nKvhRfVXLpjmfP4GULU5MegYBrLf5i7q/5Xt8vQTESc4yDbEYXeq0JYtBfu4m+Lh
1oUlaekcv+8RLCk7QKdanAlBBKzvtO1D2JuqaEpM9ds+fLNcVOlwVk7fIAFnqB9z
SLBB9qMcrj6APx266lQZYQh6uhqrvvpAoa0nc47buPePKipyJD2GOlMfSIXpS0DP
wn3qoI8neL0G/3nMbz8RPs+DgbmtXGx7Cs5Avl1AYbK0myfJBwXheZOE9BV9my/J
lsMXiZYxMV7LjxdvPLSv631N1rxPvIXYZOR5sQC6iUojCzJgNwd7nOOrUneSmGXS
UyMSWWwhZItGtoygvMIF4PPGh6hLUgMNfPKk2QhZ+TV7m3yegmm0BVbxQnNwsnM9
Fm/lzadfU4yQDe1cBydW+BuEaGmcJO9s4dnu+g6vwSgRs8ZoJFSLugUaYxjrRJAu
pfUVJt6aGcQ8Bb+9C84vB8CSV2/ZapCQ5kurKVZ7apGBey1l4IaUrK6WnISPBmRH
JAFv+TBgbT9D0bsf/96gHrFtjN9V2ozY7ojwzv2JbQj0REGvOs/4pbRY3ZF3lWKU
n/cjs3gV+tvhJJpDnYAYnJayUhjawlYu/bGazv7ZFrLOLtL4LL+AE45XSMdv3XZ/
m8BKaTGhTwKAexT4exo80DyxDp52gAZQ1XGzI99PJzoRCKLW+sWBuurGDvO4/e8R
xFwhNj5CeEn4I2s/kpUdqUkKc7uU876fwcG9RUvEFoz2qCQTTC/8mcmdGFpOjflv
CWcskdOt71tVebuDprkQFYBDnVOVZubiXm92cLg8/JdoYzXv6PEeimB3l4qJkUUb
gnqR6UyKLIBEtkcULVsTVw+H7mAb3tdZOC+2KIXSx57kcNu98aqnnYcir9dsxWWC
32nuKVkDLbqlVQAm7F9MneMXRdr6bsyknoiYbsJ8ijIZi/oio+4xx0MePzGUvRhX
q2ATyOeTasa7OfsYLCBQ8c0X9pUanE6Pkoi+9Tmp87AiufIt0oSuBCpryIzsYcjh
G3Ru/995MOKpaJRdPO/ijOHixRaTLI/QK7SP2q2ShOgnJbFBMj6CxAELGEbn6KQL
6h1oCxM0i5ilLyBys7/q94lRXZu9AVwnBP7kPYpYomBTTJZxKmqjLgF0y2UJSvGZ
guWDSN/0nEiG76IvYCa2JdK8+hipkTqsk+GLabQFfnVAfEXTBeSInvK/U+I13IpG
98Q/EgsRme1PNDG1/6ua7vSm49HeSj4zxG5YFggYheSVvxeXL+byx3xd4lGBspWw
qsSST609YDULbdjTj2U7bn3dbG4UurbEQPyu8bfqOTnsO136I5ojqANpLdPJZG+k
WS+im5K/jTQgimq/ewyomuENYnxn6E9fabaeRmxXbjikZUKAnK6INwX+HS/Drbmi
C6wkxJNzf5feelwn5vpnqkQFa5t+yNmxD2IFqA0SxGpWmLEpJB2QEPZ0OPFcRtZw
ihPVcyrMPJUhH9AB+3zDdHm2E3Y9KaQCzaJ/hJjY86R1vMMvL6D0fQe1vQX9CYs1
j+oM+Uh5FjB2hGmaz/8xvTu9LBXlU92wzO0+7n0pOAWkl0ePpYgIIQYv7/3RAFlm
+gJ0ox08c65eAI9eYLzNyyPFJiEIC3dhWoorC5OSqsARyB3kWnLO2dAYsJJaGEEE
lngpAIEQtg3VEHg+2+ZaCO7q6SbzoSctN5pk0TRVlbum4t44Qhm97pkA1m1+xlJP
1oROPBVIrS0e1ST6VgUFok0ILu75AIduGDOYg75uTtqMdt43mwVNHs/GUcQLiFUy
z0VDuwgFxlL3zPzeQGUa4jfiowOzuYSl+A3vfPnTCCKQn0Jc9q7lYRaNVpPSIJHL
StJabRvY1TmvU9vA8nQrx7reXgAbmHcutvoheIQR4x2Mpz2S2HORxPSHbXmGdNZF
dAd08ualSN/kn3GmStrBnjGcgSux9rExqqhW2GfLylHIouS+QQr/2vxcvfFRNcaS
jD/daQ792yfHgUlHD8LxsuwAVlndfUgqPEplMG6YLZ8Hay0qn7m2fXAl2O1Yfv2y
LnYGqX09cUPxNBuHJ3DusNNd/8LTkK8TAUNCcOQ8ne1sF9odejNidAqu2J9B71Dx
JzxgJQ4n9My4drqd1j2thj0k9O+9SI0y5w1f+ke+jKhh2hfM2lpW+cmqlBHVP6RC
mWJCJ8qI6cEKYeBQKtDA9KIdW/aSn6Mzf/uhCyHjnl0ahKZwW0W2/m/IrPqIO2pp
0TsUYyyn7bNcRpqRNX5Xrl4rRBFYkBTba2p7wHnxnvmH00ShEhYnxKlJAlpn7MXd
MTsUxo1whY4Kh/QAWK1Nmjx0LO0JzCp4DFN2YFGkNc2CoVzt+gnwUXpLMD44ik4J
KwjOfmuZ7Rbgg66Uq98Shujce/zJ52Pg4Vl7dQYwZcS7lAWp2Nb0mFsUrVm1AfDA
1B0ktl9UkbQqXUFBuHv1U5wmuCHNS98oqOXa3dt0a8F4NstLmTzdL8BCn4/BKYFR
eaueoo4qF0D353khAVlvPesXmszjaz2Y/I4TPu/AKIAHPixDVf4EUyScRSPOveJI
s4djy4UJRRwnMIp3IDgxe9VesRuUzZT2L94H7DUEJ3K7T+eIUz1IDhKnYlKR/CWZ
O9v+SN0df6XZccTQY48aw7LREV5ds8IXhGv0JvJB8O55BVDRRoHfa0yTNO2+paDM
gxqPHAsno4W1LiAu+dl2eHpA2VVE07x2wOFJXdcGz0D3aEOz6t2w1rJ06LrtKFph
ELj7fTPkOyyJWuvTUCkuT8EFrBXpCGtwpsuUZQP8eYJImp73LOdr6bYsyUGDutYh
gIidTAmJQ0armdKD/1FM1H52S/74WCLQImOcUcPGn5+YAPyBxyI0cDUxKyZZJpEi
+p7gTus46MQFVrvms0DWVt+9RVAAeEUjrZyynS4LvJUOIWtZxWAsL0m8juE82mNW
3DoUOUd1xO/fecTiyLnxb4JedUnQexbaRq/3XVvBgqMInJ8sQ/XlxIj4yivw8H3c
S6UM1PiT7BINI24aoVw6Mu6XSFviqLBbSv6MBiC01ECMXuQIcrwSGIWIBuVJf5C3
/ja1H68nG3XgAhd7OwKp8FEkT5Uyyig44GssXPXiZ/Mv+mKET6YCZ10TQQ8EbQne
7posPVdP5XR2ks4rkTbKql3fiSLSz/LnUleOP2ocld0r/JB7fDmaH+hE8n+vZ/8F
NrTCOcv0HVJ8mPPlZqolSDYQ2xn0C4yy5/qwkypxKAoQhPCkj794VJ9UB/gprTul
dNv/v15Z5rOIM5jmMDTbo6dNlAXVleNQPRmfMZBfqaggTkZ+5AdWuWieDp1a2f8C
VKqtXr5tHVSYbC5nRxuHjrbFJn2C0LhDj+5JGp3w69OKc84p5Og1+fxTcAJkmZm/
bwAHOE/n7cu1L6jj+LK7nWCexyWH2+8KNr08egnEkUM9J+RiSsMTQ4x2Pdn1wMg+
0XzpQVu8+TSpZ8QzN7jxW/fYiOF6OZEHm7fUkxxwbn1KBP2s34oRPk3dvMFDyeOB
eO6dGXXVUp8PloLRiWwIr+RGD0KABfOqZ5lmQvEOkcNDonDugLur8vuCIWQf3BrV
cu5yrtRjuE5erAPiKTq2X2uWZB0ZJO6S1romPiMPnlmPNHmthBP72/C89ZgMoAHv
3YsnYIHJATYcZVjpV/VW0AX1eWjxEFZlLIxC4T78/lMwLaloFHsxvhMVz0Oanwau
c7X5dCHs5dg/X85rcyLKFS1KBKDCuuB4DdmtcBeXFWIjJziDt01N5XMyP+YPvUhL
sBkrJInoibTfu/baQQX8ybcJU/n7E6Wp/yJtt/Puz5d/FlCw0NhLPCnk6vBbtm1D
AZH81irwRiXcYv1Gep7bsCJ+EtW4Ly0REyi3efRW+O/e2RsdUEjTRqMrZvpDA80i
ziHa+yYU2qUszWAqPiwdisuNXWXS0wd9RjnrbkBbx6tbPlb3am8BdneeMwWnA3p0
HoYt9/g326c3imcStN6w/pnoqNnQ881bpectsKEFit73iMAguciuiDUMpZH4N2je
DT3iaXrfJaguC+beXFfnFTnoyizlsO9J/1LdCQca3w/AXkVnWVRV9tSFdq6F07RC
KvU1t3Vh+w34wDZrsTSpYzIyUXe60LqculjJ4rjWd/67/KPAaDX6GC7vDpbNC8cv
TUH0Pzaghh2ZF6mer2N+6l3H77zwAGHWET1rEouyjbfAeSx9Mbe1EIIud+mm/ILI
q2CuUEH1/4uZCKWx/f81/EJpaZxzsmsZx2csYzDj6bdQp4u35CzxXtLLyXsmHzFt
QkRYVgUKiJeLifPq3gfi6hgfP5XHMwoAvQMBVMk9k7fqBM8R51mwWKmn0/dkx266
b6Xdu8KK9iiXIuOm3k61WoVtx91er+9c4VIBgedRCSu0DZXvigJI9e6NU2DXP/j3
5hPSZaYDAJcmoY9FiBxVxtd+vsyHywMkyqqp6IDx0Srwetoh23AWfAykAEosMXdX
dQ7Z3kEAkebKVelyVsFUH4/EJmUcF+3f4L9nsom1/GFhxpqQULKP8qIDEQjeze6C
BnjQb7eS+q71u3jWMtl82UgyPZ0zyCyT6n8/gLEZG7bhtmppQ1+pLWprv3jz9AsI
ihEdPZGaWfVqgGfusemoBaEm4gm8Ke/RneSDwApgefQWAwPgp3NFxaTFpPgXjdPn
jC1wUNFfPwpTuG8D7RTeoDKzsrWLpdzllmV1pvcRR3fHbKP2j4WT+RWfRNuVd/WE
RvZa7Jh7gyPgIQdXs1EKANC3ZQHOhNvDd0CqMI5IBA7E17XCueySvsLtZSb3t5FB
0+OK+WCPy4HUpOqk/tIncVcx+GrPW/3phAL8lCTBWlTsJl+02o+HzDGx+8CTrpiE
FniWk+Vx3QDfx2qLxcA2Zxk+k8OBS+RDC8lZMChisLTZvIXZ8q8eakz6tDhh2a6J
xQMubt6Zsy3eUYYz37VmCVPU9detOeHz+kUrOF5F2MoWh8HtHV0oA1/w4Ab4YWPr
nHTRYtAJstlMYKonAEI89Jx5UYGoailJ+QzDRnG5koWlzqGSjOYdWnh+Wd8H44L2
LlB4E2RjmcLOtfbGHq5fg+p4YcEVgzfPm7ZBNS2F+784jJqhfQvKTVTIRpgC1Ni1
ioe4tdV4+qUZaXzybgjL8yt0gP+wkk4JZoVwoJNnCyxHLv/7pSDS2nFnvwR09RjZ
+HsVtG0BkadWxvA6MB4Ll+GRz3gzKJsu9l+EC6UCgwQWEfH/XjF4oSacHeUJmLBd
mZ3pl/VCl39fsLpIDp+8UY5CdQfmd+AG/zhQlV8LzE1dvlzloXAi1yjiT8cJ/5yK
CoVjP+3/bdmaQau4NAadHOoMD36DeH9ZfzAECttRheYAFX8pEAy4luL2QzsNSrP0
1ahvLd6SxJ4izeF5B8eFm+ug6gEEZecfEMrZ47Ix0wYx48rtZTpAXwRsa83ET/Q+
9khdS2mc7P5w2tFnnsiRVsD0td2PWhtp+81qhyS8zDJg6JcNosmSPKMuyQ/0oZik
1KOIpNmLU4iDTC6DesAL/Uvs59qMTUAfvX/5a969DCDVZ53Bukcbq81EVvJI7M+S
VKaOi5upkdNSHS8dCntT/tChXflsQMy2DapOQNXtNWKlXNZZDLAQz81rL95RAoR5
XSuG6jPDfyMbLsiV6Ox7QHIkNCZ4Y2wj9u2YPAFNKj6SSjDacQabHwob5s7pwYc3
CJF7HkCzbNpQsmx5ngf8MAFfwjH39yKOyTmPIZfdiJd3+8+Wk+0EncAnvrYKZLVU
fBkCDeEDPErMmihlCG3KZb5EaNMzUxm/bsUkuPI2F3tQ1c4WL8sipnAH3BTxPE44
MuAbmrcqMbQOsuq3kpkLn5G8l4gbyJ60rNmpEKgX3UAZ9qre0xuM1pOn4JmxYJy4
lyE+U5ebFJ/g6KU0PMlM0PXwU07FXPRv8cuA2yuYVhV7HKBOFVW2uvUl8tS5bpVI
xdHGUtq5zP/BKoC0GREClYOESCqqhvb7vlDx9XDSorOcvp+9cAUwcUdnZr8z2GNA
kY5a7ZZ1kqiKnAFfJM0W5MlM1T52ogO6AfubVbOljVeb42F01PBKZMqIcmBfKRiI
SaGZJikFIXNTlrLr9bbufgi9riW2FNoeJfCRERmVjDXip9xFp111YaHRyZ/gT8fT
g7C6dJUYPw4MrvpLX87kSBUs/uGsJeIdytzV5JkLgX4ujaK6nrD5p1mVGVUiD4xB
hP7WJI0CQQ2ffJ5HxsUaeF56ECk8TFkJ3uiu9m7VGvEQqDTknKUXzIqb5BMzrNge
qBzIGYNaWRyS7NtdmJnhSwoF8MHSXp0suwpdooC7rmaNMg2oP6Xuhhd5ZPq/iFSj
O/37ozvAJnjfAriIBXTM9aMYIxT63YmFMHPO/DAPyWN0n99lCKt+DEmw8gB8hl+M
HM5+xOd9PoEXsg4Q552sKmZOOtX6D7yGLqaXrXpwJdlHivavxJ1DdWaF+PdzCkRP
8e8iY6gGvXGGJYh+WlLIGCY/bRx1BB/v6RHJqTB7WDEqnFL310a5KStFtZNDEGtd
LLSZ0UQuZ9zwM/yO2EdDcIcLQ+/vqk+3ABcKfWgKXLyvUwsn/78M2iYBGVlNU+11
x6Oj7PQULmnnvrEnYyrPeKpn1rJOy8iLp2+C5N8Zzq8bRVXs5vG3mja7WG1aWANH
Y0JxfOepaCr5bAiUkQc60ouWsYxfpGx1hMM51PaLyx2mSYE+8nkfAQM3YAL0BRfV
Xa5HIsuqjMj4S30S+d5QoZ1JYkvMsjmtnyqbDxfcAhO6BOZqd68XqriMKhqyLXHE
affFEwOpkTVbUDATlIBFDkihHB9UFoVee78YB+nnaCP7iCWyXjK8WMChI9dr/BH3
RkIrXwT7v1/VJJWlAtjZqv9Y8Iq1LWiLEIGJk3cjbNwhl0BIxUn+GsYCTJg3Mudj
kPIRCBYKwrGKTiFq4Mklvl+rFMvoqdluEXUpnVfubSkKUEFm2Qf8IzxxFPF7RsOE
QiQJpPL9JRCYMddDN0p22ogP5r/YFSjMBiBaXdkAJjRuCHzeL65Tq2Ia781UkCI6
biGxoVxuUzb7ZkcU9JgsNha4+buJu7wXjTB13F5cPpYn105F1T2cZLTTQ7EShqS+
hJVnTTvSbA7ZR98vqN4RFzTWn54VZtCU1k+9vcW20NLpIXI87DaZ3xGsJMb5WzR5
MtU2mce4dw4odCfFXIOQXMBYiE6Kv5ITpIyRvnIakFQnsHYwH6yRQjRpFEgyOGmA
3mDWC2T/q+U8PorhaPfzNG0RCvaM+KGIkxPzY07WAjW1sg7bw16EVz1m4fYP3YWI
p7M4Wtgmf/99740ax+qeTAzLqfIJGAp8ffA94vOmG0xH8/zb0ozsaVyoYpDDHxmt
Y2q0SsreY9BEWmqMXspJBc5ca3Fbp5Vb9P5ypWew+yf15b5aKQXaq4syk5pIAGcR
D6UHzRHv7qIwWQbWpseq44rXR8rLHbB14GWYfvXMz+BHuMRXP5I7eMxuWbdiD4Mq
TIeye0mQNlo5BWuCCuX+sGtz8ttz+tiTkJtmrzSgWnyPanEfteYqm3iqimPAB1lo
XFhLu9bXVlN8Pg+GxSWtXag+5ijg5q/BY+47781wocT6F8Dty3+gULoWyJHnAvN5
9XNCA3TZMkDzcw2CGx93JVRv9TeBnaMPJkOZ09K4oNLUMa9GfKwneJ7XW3HXRnkP
UtL3WygSuo07JbWlKY7kjq2zFtRLfFD+worSLUVat+cqzPPMxXYL2ILSZc1UkUn1
3RjtSqMYdOl7LMOUCxc0ygtZme38t1BuLnXVKC+1J3qZFk0MIV19DM0onYwONvB3
fuq8sWPxwS6fjkoNbAbdpWA7qGUh99rLAExOh5mib1R/vgKmU7/K+dB7umPc4ESs
SpIb+zXzpJc+EDfNVW27lmXFNMzjB8PZj2KABfxHjO8jnuXRPkcV4H+gOa4b6sJl
jkGG15aKSaIpiBNLBx82ac5ZdjfGe7SG3RstxTpm0++dKKm9iZYUSTWYsVWCFb8F
zlP9Cqczix+87Q9AiwRAbnTPCFlcCTIf13J6izsrzOj1kBjtAQdcp1gmMOpaxrr+
ZcxGyDTIe0ARXsh1V1H+15Z4HjvQwqYzpcdfXcX6qa4U1T7C8V3Rjg9P5Mi6O8co
L16sF4gn3oXfFURmvGh9Lsf0rid9C9uXBhF8s4toCk7FpM6bSzinlYSnQOVBtMD0
7N/1aYaqpzYRtNAQXttVR1vdZHLxTgJEApBMyikXPrPVYGwYTN8g5vdUWiMwE47i
Na+2XgSgK38QfS+QMbr9iqKYtrkvmCFF17XktnzwZIRxqaJmllc6+okPDfw6zSis
YIEkCU8vKZSUYwieIOPu75D3j/3LzdGCNSuubQvTdfgCiemwnHHPYGuzcADnK5JQ
g2yYLmLgahwxG4OuVy5+gVdseiNm3yWmXO3kVc06rlsXxXtcXe01amgX8W3gvPXa
RyHfnKNGgy9K+F4Q62QJFt7v9d8gUHFQGgOL9htSBbDl9GQexqs+CBQ5+S3hMVFv
Z4xqt9+FQxkYH8kZXckYA5toxinaUnunYoz/W+7fdYCa9tNHav3noN3KcEeXF3j7
heqEciSSOCQEolhHpaH0dWdPGjOGTJcM24YfIj1yn3FMp4doaploVl40fo4G5ixD
mhVuGPE4F6tIqhpB+/sd7XizBijuECj1A6bUBHMnCM9XgD+ivp4OeWbAaWRz+raL
OlKSXuWOTjKT+ApUlk6wpwhPU7/sS+5zew4JhTXyXooiX89MlEjgsu7K5p74Geus
qJbsizGnbP8vuVHCivxRXjjfIz6/9rEQXq7aaYEUNXNycazswV2IhV0e4jHrWCFf
seKR1meVSWP7SdpxuqXKOIPM9T7QrpR3ogP6fIvxOVjc6W6RgtSz09a2xCUlX459
BntmrlKf3PCHdG8nKr5C+yf0rRVc9tkGMHBgnZN9B2+tk1g39CV7zHQ+RWmiWR9m
4s+zTGFXGgXKNr8eHXRZWyHg+Q9Mk8P830rkOrmMRH/IDyPDoFPSoWY0ARZ9K7Ra
N2Dg6R32+Ux/4dZgVN+mFbhdnrpCuSXKC+Pff9GDkByMQ1rgN4Vkdwd7dY0fULad
IEBYqDwyVqz3QFA77jX3fokQ/5GrADy12IfcS6jkCNCfwIiu+3BJ8FdQi2kThC44
rslGGfv3B6Qq55Zj9ZfwiENV/7hYsWxn78sQA03BNbJsWOrpQRtDqPHEBmzRTDSf
dpbvSGMOSHO6cTIn6o/V++xCJxHq5UPOlcwQwXqMkPt4LA+VkDiuOprQ9tXaoDYR
kqzLUiEnTNhRePO9Z0HxeCKWJ2fBU5dbWiqaNYkFs2ZKR/cUJhn+HmA863AYcq19
asnzwjSWb3vHsm23MoEeXrBbk7YOATfBQ/5mn1IvEv76Eh8e4UedCxT8bI1hAde2
60tl6J4+7ovhzIIfBhgPspAhk0MJi82KWHQ7b3+uCNq1BNAkU4sL0TsSF8O3E6rj
VuyTMe5OlVOefrv2OOX3wTmkrPsbf9cp/bqQ1hDwxMMsZJO77H7w6g1VzcVRTzn4
BxT1bjowtFyqfpYsOkt9uml7dyLyno+JVRxw+R+wr8w8ctoBbp/XJ/Aee1Ka9iu0
oDKZE62RCtacTsdf6Y/83o+4cbfaJv+8JqMHUjC7fj5sX59IhJUv9aPAyl63qRdg
n60CCvB9i/atJha2PxGYFqJ7uZT90vIIzUmnFJkOsNXXNrqZnN0o1x0Ob6QJb8a+
pd+nHYVB7XmdnzrWYOe8PzBSxS9bjVznd8WzYF+9Y3Yh9/qfuN8gm6tD8ldm3eo3
n4kxx3EEW/OxmwhPMUoMOSoIZY3Ig/8RweGmGA/LSyH4uz7yJvRzUfzuIZG6m1Xx
7kFGaKGKDzdofLHhZKkMTMhbBeLIjd+PdUmb0cKMfrrdDWDvzqWgKKoyJz47KTO/
a5L0n4sSBKNjRZlcWVTHAK0hqluDBtpGdHKMGnUcF6URsgV+ynISNBVxSTOR4ZK9
lElqtPHTAKiT6eACuMizoP/4lCRVHAXY44CixVZGajwoOJB6zqNori75ic5tliP2
4tGmH9XEbrDSPOz4qXoelvL592KaFx0p14ZaS/QCT+9328wBYmMrOJu8RVJ1QAZt
HHdVN9ELU27gqQAAMmS1bKZMUcdhqNQu0Cz4rCNznJD+NUCLbzA86NtDqzQ0S6j1
mObLcGr1ss29UPY78GJjKi45C1WMCv6s7hLCnICffW6KBDG3P1RuW7d8jxNsHc6y
tlJhTVqyNZgbusWp4V4v1b0GEyArojPUxEqLMSgm6U7YJV9vJ4kkCOQr8yWxXmBG
tF/2z+usDfShmQc0SBU7L/E274a2OZototY8xj7W39N7BvgbhjqIOgUepmUUSwCo
AJpaoY6wiCF8vYV6ekjYST+U7lP5uwIJ+VkylhUoTMyP4IY39S/Rqn2ok5AGSZRa
odBe7C0SRdUZo1Xn6TK9SPV4qqO7qW2CT87Ph/Ox/asUZqcX1sv4owa+D8+DJvpp
OaDpjYqZRy7aXRWT2ZuwfTBifQAbW4sFVLKs1KgFzV4TTfYZTxxNKy5txIAGTp2d
Glcfa3KvfcOweFh1bF2+f1ccXY27XMDMwH9d/3gX8KQL4DFOs1T8DgZTp9DM7qSX
25p7CFP7vNzucNdZTPFOcd8sIr+WqSx6ORk3cys82atlZVHahyBz/4l4gHnXppGr
9mydHw96Q26N3hSbCLVbjCGvGTkzmwaXATxJzpOTogJAR2Lkr5uLszy7QU6fLpay
SBArpxIH77HdWm6DHEUTwJ6PC+D516QMVKdvO/c9b8HwumTfAuoIFl7TPv1vVuft
5dyfkf/EsXkUggubeOanFj0d8/sRiis1qp8eUV7I486rVIGy0J8sW0iS8GlZilw6
RSfb/Jr4M3N27Yn9xfmUao83e+jfb3yE8gvFYcb1KKRXbEQcMHzIagE+ZE1U/+KP
fnUz9aTRySqtS0aT5lZbFWmJlz0fkERIiNQKMJ6uTNVlgR7ZZhZJDn6HTLPKq84L
IduacVt3mLZHzeN8/vdOFXGzK/E2R2gPlfqsM9QTvy4zN6wNEO9/CMqZOiA9mgWt
XVUZ4pM9XVW1Fjxc67DR/pD/x8wYSRw6jfUHiJhKvK7Wi2oVqmjgi6pqPLRTB9Qn
kLWpkUpnWS5Wvq1+MCnsU7phqVj0dxpHwqBiZdVcZfx0+jypjxCVh5+kloT8sHiR
Z0qKyizCOJiijFbEExNjKiOR0MqnEyN58Csu6Qx6dKs2OXFoejkvkbiUGKbzYjS+
4LhFwz9CkrkoaXMVXZoH5aMD1ol94YT1g9gB8qnujYeCvwlWWlGqVaauq2fM1feh
ng5vfOt8kqi3zDQ2X7bZIUxDksc+a30a2vjtTwGQXDsCOABvHkgJbqDAqwh0bmRY
hO/ZN+0a+KxQS2rdSBLkZbiMMv5vSEsC4HEUgiO2T+BcNh2jtF8jD7C8jDtLpSP+
NN3bNyNW5/nCw4cumZNwQAmm6gXraYGYrg6NEafXojUTIYnCLMRanNI+w/1xW3Fe
j34eUKmo1Z9I0iNiI5SonwHnIIjAj5BeU0cbYbKLT0FwtbfRqtoqo1QeV8hQbvLL
pGvK0F9xvINJyVjmxMJoYI/+GFVaE2GDIkbYCyItzzrL8M3fos2vwG+WdJIUkT9R
ADSnw27TDCvjoXoFFu3wXJcXdgZQdMfao2r2yxk/9qFt3cWIQ+H4Z3l3XcHZwVdx
eNZo1q449ufB31RJYwsy/1kGkAqMWZFhCs3Sl8mDrdkhzUuthiVPnpI8BPpu46Ed
2kNDul4e6zUDCrQ95oVjL0OC04zy2lNXMKw51sjr4kd60TIDhwZPmBwqWUsqoIG5
UXym0v7deqrVOYbKR7bqcg2pmOnGS0nADaqfpDtUaiCOR0XmsfUAwueYmpnkLec/
IskcLw7BjpZ2lrwJDi4iljPHY+Aa4tGpFHBVQx0iFEicQUOwFlknPUwBr43QhFZg
csSUCQKndT6OZAOUxLECZRlVpmNhZj+CrKglI1YxQcxUAF87kgrIZZKSWrbQN0OE
so/WKRHy0HjxCxqrKS4SV3PV9hNgrBjvL8xyvAzfX/prWjLGtWER6yjx8LMaLLmA
U/3MwncbrMEaZ0v3HIqt71UzPfusyGxP70PgrCfnKJ2KCxtRlW8HHZgxb4ynGo7B
k5deq7EHk1s7XcZ+Ot8X3rh5p7owB3DdWSjTfhYqbYPr2UdQrC/Tdc8YXLeTwFar
TCwdwFJtlQhIkbzPViH5sZ2bCtJ3MveKs8j/oLOCz1sdKTwWFzZ7dc6e5RmA8J5Q
tyyuum5xutLnBO85IxUwFHvmHl0SaNKnFlMOHRMqCVZBxFynXxZeN0BKJ/D84+8k
2iqQWb9lq3H6ySNYaKtZWWSxGkuusNp5fxE1sMQSPFLJ2LwUlDu5LnuSySHObIxO
OfD6SukHASkG4okBCu9mlzR/9lr9R78buvfwmob47w0hPVQLU90QhPLUhR/Qejkm
gHILKvs0M4ut9dPfwLhQ5S3kxSG0x7eZ0jDCelUHbE890Cm9Rt2SNo6QbEh4irPw
It9lArb/5q3jTeGogxlk4VqyVezzBws8k/EW6LIMqd7UbLlkgOspQQGMrCSPwpo9
cRheYxBzK1aS3M/zvJRPXOClS1KQ4aVgEq2XRAIeC8e1V8vCmhQ6ZTO1jXNFr+/Y
Cnwuuh0SBVcNVeU0fiLVu85v8fEHrvEbTGsgnUuRBvR32n57KtOa0ZnOqTa8mYg1
exf+ABqGzqy+RC+PGpt8KxuU5cf0yCNXxpFTz1arkMVYp4SLZwAxoiA+/Wj7fefV
bUnQud9aBKz8wTNFRlLovZ+6w44AFdmbJFqEUu11t2JXGOuDvUWgCZHJHv9g+dzM
VVVD/xxXwxisc1CE9B+0oCowBy3wNlmpEYp447RX5RwN6YDRf0p55nMSZ8nDnVd8
5J8Q/qG214dzhLcq/eaOzswpSrxaoWFXwQhLzvD+v/olkoKkPUYKrvXBlU0hewGO
mkvlmamXH8IkBDCXba6vSp2ror4yKQkdCQ7CRTROWrzZcwi7tON/TBgLZ4aBiUFt
4KleDY0siq8pmH2ETKIT4ZyPuZVN8CBqbHZFDC0uIa5fSX8EU3zm/4KCYLWN4Kj+
KrEm3eZWqByV1Opq+h5ewuQjZKcpwLS5oZz2kDFDqFIAY7eIoMO6cFoCg/dSZpUX
qj2yOFKh26MAw+XdPOv/CGtHnWVBA/sAC4SyEQlmRDg11zm0EyZOXW8oA9/Pe3Lj
MzYnPk1/38GE2zhZB+aOA2GvMB59xaqIA5blxk3RXcQuMTZf0HaNnbm71L2mfALP
r6Wpm9DibKRaLgzR2kSqrq3HSU8g7EeMAoMOm3RNcRl9VAw5mYph+NTE1+59+LNK
zFEa19CrXMjPo3KrGXsXvT/ErEQv5f9UqW1R6/xxz/w9UOZsc5gz/jTiFDqG+hlQ
xhiMirHSOInjTE3GIOJTTGPbm7v3yhQRSqN8BwnpiT7b7/gYuNccmr8HB1lsEVg2
iAnM6qClkNw+aIqJ8t1xVVozuMXyq82q2DbnJ2/GMo/UAQO9amhiklaw265OgPoZ
ncvYwFItXQDb/dzhcUcXzVaD43LnfAgAj9za6QH2Bl4t51bZkc+66aP3kbuxh8kG
p7ryqRdBl/qRq0q2uw85lhDc3+PoUL795dHQiDQRx2LK1kDLlxJ11OaHeOlhyk5X
1/dqSA4xwnnIhULPflBufYDxKscpqeIsUHPVtyVPa+SJLZBEYyt/FpFLm/J+pjcw
3WkLojc1mR4pD6NpSSQdRZ71IF43E9c5DOk+/BepQFZRrsqGZy7B4VuZL/TejQDO
fJNN/jhUyavL7V0bLj68Ffxsgr3KQvEhWEk0m0xE5oI2Lr02iT6CnBTsTLJC+ltA
jo04DXqYrHndh52AwRuNMdXMugQwTPImSKEe2G4IYtVtQfAl/xVGz9oU2g49WX0I
7HBOpQhQDk1Z4agoThR2qMtR79ohRMUxqibFASLsFczXB37VGNId/H/mnrJ+/Gy/
IF3SDjnwGlR9W10kOQsP9ii74L6Uw4Fh1paaoqNpz46JWDSiqDVgMY09MRHCDzg8
6YZOEvAJM1Qs1KqOFrhgIfxhME10sHt+Ow6fSZ4+BYKUBj2XlNRNhOwkjEpiIFzx
YJ4Ubu3XLZUp+8e/2TrouyNdHDAdvoJK5veDYk+kAg7NyX/jxKljXmipJoMO9qGQ
3tadeKOKPaQWWHJOfpYAqykZVzIyrfA0cCiojXmMljEGMzUXMEjpWLZYZkUx+9C7
96J+u7N2a1H8rdSHxq9IWxbUKiTe7Kr7mdgMJXNaiEdqcySQw/8xAOrJhvOZrupF
jiR9rPYeHQMW6F5tFjtx4FJmvU6WcCy0eRCqcNRpIRRfbhw4J/NEi8NC9dAN1bHL
AX7G8KbkMwAXV9SgDlMJT5YKKhWMQoV+BAwL84sRdrZ9S8L00LiCW+wUq18Qy0ZM
6Tyx2Bhil/XVIvTSTEu7swQJ5Xo+1VE869Y75izXbl/B8h5PfGOFMrVD+zfV5NDo
feAUIXOTeUp7ZNk6KckxxafXsTqbuDNw1/yFj8/9KZmZTrdbUuBgrPUGEP19E9k0
ZjZcjODI3JGFvpPKbj+fLsO8otnfHm0DakC31ypNzgxt9TiZs/XO1nrwKrfHDBkM
RZAI/JevwrbhLcIZL9bovuPB6RHiPIfyyRYMfjtU/8Rn/AykwLBtLZH8ehEAdckI
Xq8AGanE0FcZ6Ceu8T1NgY1bv9evoBLKTUFUowk4bTJIGrUimB8uoQ5/PgmY3TQn
Kj08duMja/YQR1Taa/2Js9oT72FeeefKqbJ/qPePculDopfI4y0IIt0tXY7LeDH9
rCBcSTo5ebeXpbWDhY1BE2B6S3CYqLL2CTNh1scyNoPvg24DQ5P3Gv+/4D+k1zCC
UWWLs0wzSladw0S4dsV1sWvgkgMGrITan5CnRGfeNSuc3dksZypZaeTv2msHKdpB
aFz3tRKRQ0dn7lqNpWUYNo4tAEkYDGgFSpTp4yqxG03BxXqe218vVbFwTrijAZCP
kZWUvGDrKrGRmKru9LXoHkDcHQeSqiCMicUamficUkc/7r+WPxy1CbdWDCWp1ANz
C4Dt8RIG6nT4dgttOXJsTzFuSnpfpTntCmTUQ43ZWDz8XAgQdI0I3ZYrmSsPLmAA
q2bjJLm8dBBk4zN8cw6rporoNv9YgbJaIqoWPwhxck3ospBr91ktT+EejiZE0unx
0C4w6inPTJ181YmQf6VeqEz0hrqWlpUiAkCV2bCPmgYPF7hICM3Rh+BFtebAQWqP
64hY9AQimDqhGlUJCxKaLNTLVtUbpyOzEDBZC5w12TehLauRwiVp7zUTvejbH7v4
nIuGucdH4smNk0po0q8kEUFpanvdr7upnpxpoMiO5eGBBGe3Y4ysuQAaISnuF84B
KZLRcmhCd0yqsmdvden+SeIjcezzExeTCILQVa+3YWGyG5V1q9Ktb+T7qABl+IAr
YjMZc3YuA5hY5XCvfuPEanHEf2eXubUIJHxUQ/Ad2ZAWoW7DIRixRuZKeCjhXLeG
LfhefXwmQ5gGhS7wK6+/yrdwoOW9oyFCI57g5WLPfMO+8uXUczPzNaCR23thaKcI
NpA/s7IZm191Ntkh2n8oi6jDlp55dx8nBM3gaCTC1pH6dAFocMerbSVWQRjxuhGJ
UJddQYRaqsR+PmdA0rwdyEDrZB46WJ5icogIvcrHBW75KRbPm7+Y1brzcWm+WIhd
JXsXBXowHe8Fzxt/0ZiF7OX4pnCWPVzUYFHd6woFJ33aQKHnAk8Q531Z6UON+pZd
XSTsFOMMd0l+3hS7y4+B7o9/zSiGSWM/q3w5GYgbxjjgKpbZD6nfFe4QZMIujA8G
l1P9Te6oqnYFLeDQ08flLtqJCn7O21u7EpMwCLlBG5aM/ZFXQlPmyrrXxtFgHoHy
uag9V0ZRZVR9T/nOT3z5CZTFQx9jovOWYH9bbQapNMINImfg3omP/VM2P6tzphpO
yw8VlictJGqMC5dtcBMqmFOTboIZkf79NMbp01vJ7Y21G7MOAF+mVZUEodF47eQ3
RiLbEiapv2kQ61yp+NHkq/HwPrVGbXKtXCHjh1zaF9r0heslTS44uLNjjmo4aok3
S8Kyc8fU8oAoRDR9P/aCLELX3ZPfn8NmIWBR3gFE9sHi7VszV4Abdn1LozIdthoP
Gw6RLaUlSVQBm3VLpsdGCNM71oNeNcMDjMVY7rtQ5sI2cYo2QtP6BmFT6HxJ9fch
oMyDjbHFhpqE0nk1J8FukT9q/7iBXCTINU/rjniYJiTWCN/GWVayBDA1xfABmlFN
fRD7blmWDkZjXpzd6F0TUFSBSf1nt/xyHUmiOHa6og1lKMqcAUJDIj/aCmdX8oxS
2QyPfCLX63sAJc2JHjlxPaHNiWphcOxDpkpqy/2sEmQA11p7KWWacbs+h2D9mm1Q
dVmyQQdE/wrjFRjBNnmNe4KZOqeqmLp4bhBBW6W6FJRUfUbDojSrybug6j0IPV9A
kRdx7nqu44CvGT3Z+jjlVMubG6ubiwqqfyRgZ2Ba8gvk346/99alavwFY9gqidSg
wH1zGCouYEU/H7gcxH77y75d+Cu9gV8H3POTEiKiiLfUES61b16AqZVo1dncQ0WV
SOr7U8snc93a222gALNC3SLmAC0jJfnzKYXhMnmU1NCP3KOzg+X7s53NWFxMAeJm
XT8ku5+XIpBGtvYxEd2Yc/gKQLIsrGXReu0SARso0JnNRKiHVIM7dPUqQED3vR1r
eUV2Gc1DxEHdZnkd2M+biS1JfwleVucm7FBDigCNUAC3bWxQ6zW2fPFPlSW1v48G
ZH9AastjRz79a4FefbeK452COgQ3Ne1HOa0kRjbH1oFuJiWt+ClUulwIRK/+ZnCm
NJx4DNBnY/G31naENrdPcihNKCI5+85edEzWehvSuE9531kD20STgVbpGB6fbLT7
HedqIE5UXjTewqLGoz3SIKQrmKZOwZ3YbA9ALQi+PWDYnbXqxqWEL0AI7iRM1Zxy
EqENHT1FWnICpktepe12a6atIG1PTSefRlHQabaPFdN31qzG70/wLirAa+HlEiw8
cxvmeOwnh1x4r8BtlQe9i2gXr8eLP0Bg3Sh7MfuMMsa6gVoafaeuykd4zlt+adVR
l7mr3VV8aY+u+p5XVsSxwltR7e8SzhCvjzgv6/IoYZb6zgqq5D+XQQPMQeSHbRPW
j8eXlynr/9vjaZ/AlkcOJcLMyFWH4SUdZ2jThfBnQ51/sR4H8y2JrnqR28NjUOK5
1BNm/hZZsMZkXflR4xUi8E4ipgVxLnzeEBY2CqHYxI8kzpcynk21oc0vi2cNmidg
o5psohL3pjdUbpdzs+qPndGyzfE7h76/tMVTffLlC7VYAfHUAAf1D0HQ3JTq5jYP
SKlg/pWaOjFS/ySkaiSfnyae+ov0BFZdTwV4ZAHbndJMSUXa8TM9zI2eLHqdN2tE
nZhbM/nOmU/fbKZ8ILZv4KvDicFGy/FJJiltpqGdO4NDUke+dMPwVZwwVjP0J4yz
Jlf/48K1K7psFR1+y7rRth9FBmEbr/z8jqUOc+WzJraOqp/D9fwd8+usBU8lVGIs
C7bBdHw6jmqW46kEDbJ6pYhG9RHbHOOWncJ38GMEBoV7EODV6GdxEcgATuTKmsBt
WoauA1jAbva/Eu4UKkVwpiFsQufVdzRK/2W2xZiCbF7ACtzWmOiatbRao7oVvemU
hikADeMpLgVq1VarjoROBFBhqAT3/ltnbpzF6dP37hRbtniZC+TxERzbpA9Qzdk7
HU6NyL4ckTYyem7ULmiQV3nrriln7OwR6dx8tUaBFhcpgRq14k+bfENcCWRz0gud
J1NCdlP2IvMqyq0PDHhvqlCBg2l52qInmCsipN2EWuBEKFsZe1c9mZXyZoHYQVuQ
ScfxevOz6yk4XymAWwIdIuT7Qse7cXovn7MK39Vm1IH3CgQo9Nhoet3yjIl1YSQy
3b1ZK1FvSuIXPYTlRY5nHhy9eFQMC22bRBZvIzjIfnkg7Kg34t0fsARjFj90hQ9v
jui+wG4C0x73i3+IraN90Ms97l17ifmZUnNwdLzazHItYt3rIt/R/MV4oWZ0EeoT
Mlkyq6fBVGeOYQiiHfeqCipChIatkfLANZ8rsYVEsY3auJUba+Uv7DsZ6LBzs684
8Nry7TEIJ8gapj3So03cYxffNvHo837D8y36iri+0Vzv8KNSrvgTnruUXA5ehHmP
IdMj5AxEp2xWPt307euFNTYLWPw/6Mg+9mrZ0QTtFi5rGqwokgz+vMZUlkw68OiD
v+wUV7pfnoGUIOTidmovCmuPG+HtQ77FGcx3z59xf4eeK+UbxFliEWa2P7Qbb3IO
qElGB1GLmfCL96R6YbCkcWGZCAUz6o4hSysxceUqh8+USf9tODt0TQsrSvZdkmqV
EJXNyaXd1ooBUM+S6L1U4/f3VkZ8icT5EFl60KXu8dqNyvYcrNgJLQfzg7moDx9c
CA/oY4GBr87KCGbXQKnSUX568WWAKppOk4633kwfyqqPXn6FOu24P2a9sbE3xzZo
U4yi1HST/LpAFqFRs7cPG2MlS8OirJGAZ6UMjTsfXmpD7+l9v12ylcHsEQXN097x
IA3L9HDC79FMhZsyZTenf2kOkrELq8I9HmsAb9cKNQ33Wvd9oTVb0yYUecvihLbV
t/Y2kH5SJ6hhbUi1TnPoTJc/c9CrMm76RQ+9e6DJn1ydFJ09w99FON8FdIF5UHlX
jrW0b8vWLXVciwIQqmBlup655d9nEfpnuT9ZxFTUHyquGXSeg2fUYuvLEqEn36X0
jsvpUnFvnG38aaHFPr/az+apE7Ux/2TwFZYtUdslfl73J20MMIIjmP1W/1pixnqW
MCeNj+hOp8uwWn2/g0yjUnhA9AdX1Uf/64RczwgfiiEA7/dafLnaMLOht+/DFl6l
AARZp4XJBR7o99Fsn3Pi1T04Se92LyvNb5XNjq2ScbrBoUYxcvgiw5CCh7AUe1tb
246PZQcpL9vjvqFGaS8IynZaUyl1aO93V7U2ARhpS4s1Qa8Di7AM7pHv/tlFoa+a
aXmEgQDKgxDo4WkjPLC7kKxtk3aZB+E2kzv/SSZnwXwRPqdfADcVmoEO5RQUQ8jd
FinQxW1n1PsaTq697AfOsiNWSk+buYLjben6OJfDYjxxYb1EocQpw3WJvaLqnReD
bUsMKNKO+xJj8Pv3BKxZrFoOOTG2igeNj2sKVKsoTKBO9rrWOSOOWnAYVgC4A7WT
/paeEBhuazN6KGnGQ1s3cKx8PLk4nj/pH1Q6zgezwUBsDuYSHFEh57rDo+Iw+i/1
uWUeDQ7UwQ93sc4iyvXwsBns/AujZwcN69mNmhfiABkQ+VLgVcavRpNFcOZmXTZT
HqGfGpsV4uZ86PFayJBGiSCnXBsEupM/9U7lSDWb0oSQtMZuSjyM1P66f1UNCfSD
Ahde3AtizdibVOyYIU5hPTbPd1YhNZRT0mICQOJ34R5fK4pfvlNngmC10c69vm0u
mS8cvi1XvVhZfBFJaoa9BywA8N8HqtAUvsswtuKVg1yaAB73c0tejSn6o8QZAgEf
EsHV/xMxvQSxz2y8dpjV4eEJtvWkcMLg9swiVtC08FASsVyi7Lmpat20aVyq01gb
t+mpyRaRXFly0Y9aFLBQspJK3ToPKEAP54vOaE2Jr27P4uCyhVMeOl3lka5H/1qE
wTGj6a+83u1XUMUEEAHWzr8VnQBf9jxB915O1PqYOIV3Bu+RIc6QbTXRWvB4G3H/
4wZC+thCvXl6UiilYXhK/hOyoj1L4kePQOJID9E8k8p/vEqf4cXNU0zzzQmdFZAC
jRZRPdx+66/fzLVye4Mugf0muBzmSYicFR/dsnxPr7gFCmVyVJ1B4D8tpb7Hzc7K
B9j3BF831T6k16XjVpiUF+SbaVMWzXfxRjD9qnQYzqBvz7b/Cirk/auYY9yrUzVM
RmwecG0yN6IgxONgPoVI3ZriGRp8elhGX6qgKlI3TAoIVB2E4F0JzbXjMnOTKsOt
Sq7/at3OLtYL+bkvaBeRgiIMHLkzlX59zq8GHbWlQO5SwB3EIEiH0NPV4TZBM4HU
T3M2vesbPnr7lo+Zgf9NQQgb97ZZlK8G3PsIy0+np7WjEWfrN1Ge3oLWbQAZXtgY
DejYO0R6XuTA0VcX7zn9RxUs+bwsBr+NsUYm7suYDPSCe3WaHNeFWpr0uEwQZI6m
GdQAOq6EiA74PC3LKJ7nmwT3ey0PLA2ejEmxIUktvDwqpJhS6BRffcRz0RMcbnWZ
+G2x70GLGf1WZuxfteCUQnR5H94vmRs1LEANeevFH7G23c7srl/1/dXBcNe5sio4
UAsBRaqMTIhIP4itu26Svn1zN4QqV+ZkuIJB7cw8Afu1pRkPLMQnHjeO/w3rxr1y
mQUWtp0YT/Rhp2D02n+5yqEn61DNkCZIUYkK+vAQDR9xXrMUcgZlN3pB1UbEMy2d
fc8clc5H3CWcSR30xAYe8iGZo3USg8P6750z9uvLDV1SGg8ei3GW4aTJokzmPAUQ
crHXK5+rbhU575W02W4vTHqC0UViuA6aflkyfyxvO8lVO85hMyjoucVrELEIR/qW
J0YKrZsg824uKfW1sHnGWhb8CeNKrXjM44lD4Kz0OhVkFQeOM2xUysxsfvJodIw5
uXwaSsAQb7UQ6BQATyVj+f9bn+30bgSeaxJDN1+f88S1rSDBQgP2w0Db63U2tyTv
mzVcuDuH86z8TZDmW7mc6FXBF+5PG/NAkgLQcn8Ol8+U65UPv/USiUJw1Ax4FaI7
CX8+c4rIsV/2qgxi72FkNV0l7KoUeFVtDY5JulZgmReSiHhP4m7MBDh7U9Mg0For
xfIR0O1Px0T18Tf4499kOG500BpHxFKUAl9Mhy2DoQpGXFWBBwiIOkW/vkNrjidf
38ybcRcgJZtGIFAiJPv+Ft4SiKeaRZoYdz+ObpIUkmwvWwftqGGAn90HuHje+ML9
xm8kmJddEnT3EOb3rQtRcwDvP/9Q9cIPWAuOK7qF8oNsvf5cHiPpOnYY2PsEQsC7
lYUQiMhsMEf3fPcHSjaijGm3SV6sRTd8wXf/xVMofsyd3dZv5yE/JZm7KTsBtfhD
Za9PbwAqP2wJ5mFskmK2IqobgjlbsttGEbeBYH4XuBIv2euCjIRmnF1TbE34/7UZ
rx+ONZclxS/nHRrqLD3Y5J+TjeaK7oPpik4GD75iBflSubjkn9qH1UukvHaH+040
Qgsweo2qcCT2PigDd8mZ+GxE1cKJeEbLTWLle3JxRZPAqy2kHdCThz05NDCxNt+X
JMinBypQEnvYt1PC5e9JdCyj32zF2SHIMSIG8a5CDRocf1RBkAUfupGObKrJjm8P
eXkp9i8go4SxTewIfrWJCIROdMiSF35EYCnNO/JPPys+OJXmmRPey5DZqLG1dcKT
OUWzSLGo0jwh0C9C8uK0rDH31QYiJKiu+XDdidpwX6jr+oldnOLei3iiTaf9GE/t
v6bbrJpAH+mkv2sJFL6EgEoz/EZEs/Y+0wLhqXsCdZBs+yeIdX19xX5JbT9rMGxQ
GvSVTI+mSge1VYS45iHk4BxGz5rtRBV0FBOV3W39KRXDvCpkozQm2it4NBmaNOdr
Q01Fp9upxNTsdd6jt13hBV/uA0+FdSGa8FHhkWEBmfqcdJKcp22vHNlsk2Hf258L
uXlEIrvTGzZ02hOKxgd1iK4UnaR5zwhnJ7mcQTUK0NvFBQNDUbF5uXNpdQgNCVo/
1nYK49IGpmegmJ5JfzIGzO9XczjxT4ozLKVj7nITC1Vbh2hw0Cc7GEi0IX3jAAtA
ZEGqOz6ukuGhSl8vGWiGKXjO7HK125H6DNnUODx6UCLG93IkDTMSQpuZs08DpFSr
HdOexB2kAxYOxTctQJq9t/ZcNUwL78VjLMnDTt0YxHIBurUmsQ/2kl04S7LZEoBl
90LD1UysJXq6IyrHaICh4CCJg0LBe7lE5iC/fy+nX+T2JiOTAU4li7QwYzhE9/ea
unRSMlG/B5UofrvU+3ySkXt/blE7r0G0fbyvmlmVm5raV5+Fy9jN5erh4gKbMWwj
0CkpLBAHijRQXBSdKs46ugPiPxrtuD/OuggPyhS6whFqt7S4bsFux19HymLK38ie
nLcLCr7wR7bBfXg9bA629Hfu8X6x1ChpkvwH9V24c+vUB2XQkAGQ5fr0K/OSpkt3
F/piVD0ITzJKAQyFRKEukHze8snuULzBWDiLPcIjzK+G5JwYhw0oJaqhdJswsh42
PNCfhNSva6x6dU6YJFu3UV2auzWANwcuZb3vTuuOuKr8V3vxe9a75CfeskL/y23r
T0cD5G++1+6UtbxAfab4DPPnYB+BYOob6npcM80s+GdeO2+SY3si3814WgrMINB8
8ZRvYd9hXmDbJN+gOksn8QrcocpqWgjeMN2NU3E1+A9LXx05KMNoROTNCXHHl1nd
ce0LkdW7Y1tE692lSDWgkAax7L6JEapYP9BFXTFT4pLk/T/lkI12BwOWELoG5H7p
D8UUcAu8UuYNSSSPfQkTjnxRwxRZTJlThmp8XakHf/fciH02h6TwteIjWwqzboZ6
ewomb0rHp87eoCIqX6bZ2gO1FmUV8aOZQ+2lBcvR5/qgLfVFpKdnntTKoD4/8Ssd
azDtphzfLYbRHheOg6un959q+GmGsM07biWZTZ4CcfbOQVCq3NxXbL/deHSPlB8C
MQSTWSc2G27XBbKWBGp9duHQo51J5BlB7OeVOQBKWhC81RE6JtUBbqSfyQd8D52F
u2U1IEbtd8CHBlHmtWtc+H/H3XphVTlo9un57OWlcRRhcNuo/bnoJqxxTcn/TKpU
ixbXFWbMb9BLeyN4O2GCLsYf/Q/BFa+VO+oE0yyBSLKSDqNU7YY/BkPkf07ARlh3
1ehkO+cTtjJx/4yHsobYnBxVglWsRRPOXTW6WMRDhhoX1OcliBNm0dNMNCK/StKp
/etMbtBLaW6gDhy4q2ljjnn/Qrm7MBa1f1RmF4qiCdicVH8ELlHtCBzUDTIrpPjq
D/yV9et7QSA25d3kEybghk+1I5hD04p/RT1k4O8LtADMWCdjo6GweSq3gK8BUYv5
6PmV7TnWGvaFTUaUZPWr8Ryp6NDt4+ZG/aY+2upjdp1LtV6x/JRv0EAHJAXbPfbt
Vu92ouI+SBO5DBIPgFIPXyR/wmGvACmnlKVZCtALnFv1AEZrrSRJ27qKYtuyCk5v
vfX8ZbXmOb7LZa9NQSExYOYa/SCqPraAIfD/UWqg9eIGWvammK3OTuI0G3Vo9vbh
kSAK4U46L0JIQEw+JiBF9qM5x7NznX6qyrk66d57cwSHGn+yfV/jnpRMAqe6wg/7
NT02DLg0Y61i6vqdHbrZ8XjgLrARIks8SJCW7k8mKC1Px74an7Vr4DlCyNT21b/j
u3QyozvJndAG0E/14wjoE0u/qpnN5NsLaLTI/S31paC2ZH3u7FW6b7ge93/cPTVP
hcygGpbm2G5np5J+3G/nl+6qlBB6hd30TIGLCIS+WAJNw2pAt7x3tleekbAaKIQP
+3CHvJe6EIVdLVEJCAYAmClfsG+LOWgUXOe3QHYFtOOJWbe/Qdq01FzUenVI6y2+
Lj/qMpyzsI1QLQ6SzKECJZLxu2reHHkpz/Rh8RF2GJKKK7DdDKLZ5rG8aoO0vh3y
nm/YRUx+gZzhhurW2gBGMiroO8OFGZ0UMHKzv3PQ8HTdmGObBsSQBz4IhO1kVYFy
vkFOTtZ5ImtxbLvhOIlPUxtc3IAQNWga+IprZGga7a67wMXZKN3WmzwBUG1znXQR
TaG9Wor+rC/qA8r+RUJXltPecWX4Nae0jg49jwFVccIaE4NfPV5GqbX8zTdJjpKf
iNbohhLHf9miuufmz0jL7ecUBtXcrO3+LMTu/xKxkEypSbykH1tNESDh60w/u2bc
qGvmFOP8riNPJJifceWauKF6AHHutZowPygZmiFgxm7zOQBzBpL+KRLZlHtEQXRl
k3ecFdJzsqRD+iart9BoyUYJ/zqJrviJMQi+vdGtQsd3mbwJtUmLlzh78MxX9yjo
/q1dgU47eUAWKmCKcRpviCYUHWcTEpo/e8Dp1iGFf76X50vURocyv03SvYUpQ7Uz
nZk3j7RmwJOADy5XYEV07QdLcvzn2gS/TONTLvBcTn32zCTbEoUlJHJ2MvGxuhII
Z0wBSeVhNVW35pklf9h5kOPY2UU7mUB+kpv3VGbPxNZ/nFI6elfwqMVMfPQLiNQg
9dv844YdfdLKFgUIGxqldlp/twNCS+1cVKqPJgtQlrQBRnqUFS0LFdsj2EDeYWdl
tLwx8KMDU/pQCvkXqKLyPF1pcrgM5Y3+wzd0zOMFuusV6s1UidUstzIvQy71lvYA
wvMXMOl74HyHxaFImWiksFfdBMLxuijUNQzmdt2HfwgGMZf7R8/gjPdBu6yI6C+d
gcoifHjyzXxIaP8q/1AbGm1iNdLH/jj9d4R+YYssruY+4F6K3+xaDQ+p2Hv6OJ0w
4H5o16FnJknxBosrN7Sl9vdMBj8PgxaWnwTxdLkWIkE06t7HH1/4yp1pTz5pWwwb
usL5/o+M8mWVpBUz1zyxBq4gxucrYTygotAhjIJPT3D6+yFghBPinF1Ec0hL9lnw
cJ7CQqQ/Ems9defKiz+umfPf+lV6zQlmb24uuGLtlym1EROUYMy2Jycgy+/R4IvY
/x1jyAFAFZLkRbR+nn8771AYTChmetO8T5cb+fR7B/yf9rlO3hnysHAJdAOlwT//
s0B8qZA7qy5d5TAF9t+faM3VcsK6sUvGqQQVCN6gvPGfMPRuvR2gx7yG0SdFxHxm
Zh5UiIWuDBVQpzLJVFNxXe6DSivGsxYM9nu6LuPLrqhLr9nINuAOLy4s21hKbw/p
O0lXWIUuXWsfofM+lDRqMjNvpNL3Icd0uJPSMrZL8GO4nuheZD+JMhDr0yxTJtC2
WTdTHzBOd62UjuSgzTLJsJXoBTQPmvY9xBZEQuB7UCRv7hTmZO/cvSAkjWIweVSd
QhqNj5nJK3mu6Zv9xFp1/EPEzPIW6CUzQt/JKewAlbZb0Z+g710nzhu01v6v+tHB
2XHo8d/Nh4jtkdlv8yT+fO2Z29hAN5gZfm625O49Qa1jctuLg5gvflDdvWA/un0N
d1+1BsObXT6fUaRPFZVFU7BLJHkq6Dc3PRx07++HOkIBrMuiLIUowAnxao+FYzu8
AufdrhO7QQPH9AeTVi56dkcQE2YHfylA6VcfmyXqGDl1VTOQT8Uui3osTrRfWzuU
LttSQ2jBFshQhK6fxBYyJelF0szegqeLcRNluQ15SDFCEfjTfSNV4CPiFv8TH5BP
Vg73MX36QkHK/1WI5+KAestL/OMKup2NiabQkB8ikEOTKGmIE+7CRxTH+7rTcXxW
qzAngbkcChqHNuawBSGkom25ksK4j3I+2Ai2lUMaWIXNdnH52kBf6zN7D74Pv9TR
8ZFD2n0gN3ymeUzoYmyTOv1kYGDafXFjXrcBrjlCa3CPEkp6A/+55viRs8lrCzFL
rI2qCk9lHKv+f2yMXMFc9rY6jSizlP/sWO2J3kQsfyUiQz6GG4E0oP5NeGfNA4sj
LAO7Ask+v/3tasne/J4Bsasc/+RHYlzEbarJFAV+LaSA3uFurAbp4oDhE1rS4gbS
f78Pn2H7NikKH23eTL/Y5aVZu5LHkmzio2TPkTXpe76H/5Twa07Y9zGlcp9VzckR
XalpMjPCg63+puBYPX1QBdJkIBrQv6jw/iycpiUUlhZdICRyrwZuFLQILudnmDR/
9k112PDUmWOLCA22Y1psw5/PYnW2IBBHzCSrXKeGu+7h7IJW1B7vjXp0r5/tUMIE
3JmD8Q+6Rl1Gdp/0/Ud+2HorO9EfemAbZ1A1zuC3VOMOIyJwpZz/sVr9HPx/PngL
BStDQYlIHmT0FrSuh8lXIS9iFkQUXo3VsvgZK8NthHrY/1WiNhdTYWycXLG3+lxx
x8aud1W79taiptWP8M5Dblhzv6xPyriX+PzJXrwvqra/Hpns4w4a5vhytb7dcBc7
0cGKQFqejIfwgMXlV16PZIMYOcGRdoiaBGoJ9zZE+3Jjtg6e82j9Vt9iNuI4qKEn
8s1ZUZPL8ZeqsfWo6FSHtq5aC14CO7evIEy2PxOnkc9aJQaRjGQtDCn1RL1CGBEj
zeDc7XKVEIIjogsueJdwT/2Yxq7I5Ir6PbuwIULct0x1FbDsL7cGL2C4lUNoJd3Q
EuT48HaPRoGDey6090t5SoH1g/SB2tjF+GgMA+T8Tzxc+9AqsDHD/sbHCeWm4v0C
nY5zdmVfQLth/nbc8qHHGGBPOWl3cj3YYOLlGVKbFRBIXBfP57exc3p/ux8/fE0Z
6BZKayTff3uF4M+2egxQYkY3wCj3k7GyxGcB31etp6eLrV/ZhCQGF6KhS7vvSXYl
z/ko+/sx+eAC4PSOm7jdb9P7r0XOoIfPrTEH23JEkkjJ0PnbWYmQJ4WUWF0fBxpp
CbiOqRNp++aE1el2eXHiFpn5rBLl4xUJQAQVjsOGQKQprUflJAAzN1dQpDqSm1fw
v/eulzQ512+h1YkI3P7XpHtGGoRWVQMYOZHpT2GOpStQAxkYf1eU2yJkOWx1I/HN
25oPSlRW4MjXBb3eQJrlHMoUYaevdjYfRgAlIrtrMB9FmIUFRyB42N6LcZPS/sWI
rgoiJtLbLtGFJZvIsDORitjv0wEjKPsAVv6c02Nw5K98mbw1ZxPPeaezH8cO7u23
BuhmC8Z+3viv4R/8oUZipvRtg9Py0zLPRZh0WBL/0cdTP5uFw/Vev8JghvednTCD
WDF/QRhBPkq+EdsGGS92hmkb3DWKWSXT8dp0bn9ogV39L3XcxfL8n0h/DV0gl4tg
AEc3Ks9MzjB3DuwG8l/ogxmq6XoPJ3wNpRWEu+lf2VjgVAq2w4z/ynxw1u5Aa8cn
4z+0NQ+/FQNv7OHCBt0gM9D00zW0/O0Wg0MLea8re5eymOu3IPHhDtMYsgmxhiOj
byCoxT2S9a6y2XlxCnsXJ+0Qw13g9YxI1cRo9ztt+s94fnJ+/3S7yEFjZxaOr03Q
IFLmN+F+zk6i1mMla0QlwD4V+KEVmWSkQbvXPiUIkoUDdfHc3vAbrbSFCV+IYFw9
k8wlDZCSy95OthMnRTpR2yZuIJpACdsPWpX7uJaHaqmi0hr2XCyVJy1RXIx4vZFf
GnoV4j1B7pi41vDCa2DHTuoCldaDx27PvyFOWrK6Z/8wh/lwVYW9dujzR85QElrs
CWrss0/zOqsxSdp93QbBjbhWaMJyzJTZIlOHFXINA9BH7HrAmWN6AvhIoKzu+Syu
7xTd3ZxIRxv5eym01wf7TAk6txu/DoodexY/zGqkqmpix5Dj+YcEFWswCzbZE/ZS
W1ScRB6AERA0hjJsqG6e3uI2GVrcXHxCihGhcdrg4XuUNBvAS2TshHR8QU/iSedw
1AywvF8np6fi98mrCN6FPS1Z5+0BxAD6aXBOTc1Gpjpus6zuCsePRNFuwmrWiPyE
kgsRLTsifJ6QTHA2FgxxNVb1h/MsyWmNivqexc+GuIuwfsuRp/Sp/iau1mXJnzpa
DOxwmZ25lgVZgwP1NydJRylh7VBtQaFXs2PMZAHvBdxb6FDSeOwaZd9XkzZ0Ny0e
FKs7tZPCrgC7d0RyZlGmwwIP8IIHG0sfzAr0jdM39Qw+mWA+ttACZWXzbp0WU1Hk
rsMxsOCoHc22kKLKebzOD9cKxeDA+zCPTOsb2ycDM01gK5DvyrQJ6hvsZPkV7coW
QJ8yerBBWjkA3WhRemrO+Cuk77tQqJl9rwcSKbtwrVEPPZtp+oFXOZle7G1DinRF
BDfkW4f2PD9S9f/P0itIvHDnJvsC3sPd2vkt6/7qxxMwSjxo4eo2DGQE/H3QdOtf
MbG8RdSJd56Ordxs4YsHMhI1n+EO+gyLHJwgXakgKcLAtEmkM2PjQPEcB3QyNIMM
e/h7UES2hLOO8/0IhCxZ1OPBjPoSFTr2SPFDKlRoKCfqFhzKq2unGFTQzeZTgUv0
BSWWby3R1BDXfvKkB+SryFAb6e/UUbMgP8kRPYppZ0zaKoeg6BVbkZR81ecBcGbe
kMSwyJmQttVvmlemAt4Bf9qCq1UMSmghqCY9ns+Hja3jiIoapKjX4m3R7K1+m0Jd
ZIMkfv63rAxG8KCXBz1XIa2Fm/yG3freq978JxEC2dYqKIZUiunj+ztNCBJI8PKq
OjpwkkZNRh1wVD14RwrCrXIJNiWYuykaYH6SV50UPyEBu/NVzjZ2B9LypupM9G66
NDAaIU5eVlfhT7AKn1VIhamTyTRZdaSzzstF9zpRGyFgkgN+PQ1m322o5vq0f55A
sX7pRQuIelgP2CXaOxlCl5lCwXDZ/q41InWaMOETgoBy1lmYGFMKIM0AT5As/iWL
pRPtyYJaONpSKWX7nzLUlNHD6FOscRPaj/CeTpDtAnRUfC8k/6MZ1e8alnsl3fL1
5n9Uu75LCMs5er4lCJ+NmqLPTm2V+W0gCCS6ym7l9xhSb2gdQddSbbTKNps/ECZy
BQ0W1l3NLGrILD0paHFJiDnWfkOkS21foIqGFipb9ZqhyrFlkxZTgS0UWykA8orr
czbPzNV1PjT2E4amc9S+tBBGti9DIF2GjyUX8D0KGPU0XKFVDWfXofleLjeCTxAK
qeeSot5q03ekQHPY3ysYwDuusO9oT+MgEHO6mZ/2GJSfmJGWq5QuTr18r9UHbWHB
/Ct+nzBlHjYzKqnsdM47AR4I3Ry64TbmpfBRyKFRdRFw+lL/cklIYeKx0CmQT+Ul
Chn4H2LnHOaPZuM+esVqby8u9gidAqGlAN6kqZFIha4ADlRXUCMs51IMP0eWOaiu
q0DMUYHdUw4gUJ0+99SAPsuHrF89C07uuGnlizQK9WRk+TF1DO1QHiv9k0m3RZhZ
9Q3bPiSwR1RUHL/Cb/gM5gW8B0kuOVVCkQa0bCK+7TTNru4XGTMOBEsWoUC2MHB8
WtJaDZUf4BoYkU9F5nfVCTL5CzLnEZt85xege2VvTCKRGqp4ygulWT/hoVrITc2X
h8M7jJzJ91ORikGmZjp2Ehn17lwxZuAiBGK65xIacOlyjUBt9tcolh04Qv9zFgrK
9h2Kp5YIGrvU0pXwbemqyAGiCYLkNowmnvEvljKW7u6i5yYsPlYkKQexd2baaaWs
UrZ/u+/q9Ti1mFAMUj0ZyCndEWRMu1I2yNMhHzzq6Q4nS07gsYWsxMnRLE606c69
bJm4074dADZq1xm+v70evaafybGiKdPQ4s2nuE/OTXXBL3kIHTJg0GQtGGEu0Zo4
vqJLNx8avX/f1ZfYVA0miIH2CrkL3C2O57miK155y6r1/8U8mOoFH6Qz5TOJ+AJ+
CWVdNU7i7Cau9yqDDXiYIxC/7XS6f0omDnxYgvSwi0nGdT5RMK16oG4Y6R3rrrpo
Ji8btUSRSke1L0I+jAkzQqTH1g85H9jwb7NMc2eQFMjmjw5DqJRf4Aspx7WNF81i
f/Aw/2Y36ZR0fgYECgbaoUHxuFwWimYGi3WcklHStmL/Uk2cMsQ9YvmABTkFZooo
FZWGaPPlmlY8L50+kcT3W3i9/R3qQoqA945vyrB8DnEPiJUbgJ/mQDys6sztgbkp
BZyBtHLDyPEze37vRuV7cm7c2yIT9vTcFJxtEON6WS0cVbnsTkYf/n2fCCpTlxDV
OrzxwZKLuVeu6rBQpW7VM9pClQHlWjvL0vW8mTJ6V2nv82oasTImI6lOTnsKTd82
gIdIXtUuTvYCVEm6wE+V0MtaPl5R+ApGYDt+chq+Ux4XDBqUvpttRlFaGclvXZcm
XCb9dUE8UEQ/2Dp3oeGQPinvaheWnYM7raVJNi7vqRqFLUoon1LQ2p2rfVPNVrBd
FvjzhTwlelBuZJtIQy1oYEHPbcFpPV8w25oMWe4LSincoQpyNKwCW4Ope2MRmMFQ
f2x6trQG+GZHxd0ynjp93xnMt8OFUITOTDUwLsASRI0Yf3KJl1eBZWPJjqENLGez
4JlvWTp8ZObyi5twq2me3FOOU0oyJIEqNHT4TND57CIWpnekwsaOuMWwaud5t1jU
BSzmiThb67/w55E4tDky0oOxXRU8djp5burphSxuAx3DO8IVIfSbRsKxI49utQ/h
uiDkJq35IPgzajpKNZe/ipU+9X0sMJh1cgzjLMpCdggcQtwdHWsKi7lSBG7b1o+R
cmD/bcuAAoeuMd1uMC/aQTibzl3KZrD97R7rTveg0RW4wL4nFQpP5rMeYlv2PUZQ
WtYHwTAw3zsTYi5ScRJNEOp9FR5bnzHLgVo8rf39nJk7d0NZzVPjV8ND9JtRT2XN
n0xKpEOKydEYtI1d8Gb6DjmZyNN4DpFgzVfcqktZwkz11JRhpLAkU7KJoPS8szvn
/SVc9ZwhgDgw8FQ/dg2L5svjQlWw4PX+GKuCht5TquVx/lzcQ1jw3Dhty5DqMM8h
oAcfJcaGjYIMFMGVKmlTX3RUQDAyUOHkWhBLF8uKI9ZAYi23Ey/UzV7X5FwylaHi
ebJYK9GR4ndkQyOnOQPT1YFIWL8vt1fCWeXDnhFA0Ai8srkEqHzhkPLp9zzkrHgL
+IpXNymTSkW32pBI8Ff1X6u0oWC57O/XZW2EY+rDsOvnffkTLNdGm7Jk+uuwlXzs
GGvun5QT4r7k+TldPpfZKdCq75lYT0D0o3Jh/4PQIbKZhbXs83Ewdq/8XwuGBLij
B2bE7Xj9ocfh+CkcNVLNH27t6+uB9bYRtXYiBvIypx555E0/n+cIa/gOshg/pa3x
Gx5zNWDYscvLTjW0br2qidgB88T3vGuok6qnDQgtaHaOIY3RjnpAw1pIVT6HIAkw
lCKVCunqb1ARbY6WgQBohtpdsCMpFwmpCsFvj40Dg4xE/9YJHQVE1WHGoyJend6h
2xulMSXq1LryCQeZo+OPiYHKBDGC4bSeAb+BIvJj2HvL9r8usJANVXXBdTr6C3kF
UyNVsAtWk3q7+u+qZaJUgfC4OxlNzFtl08MIHCn98iaryLuwwKWIlExTWIAl+B6z
1dmJKtCFr2o8h2Ypr7Q/IFLZdHAhFwP9drkMezK8TRzNTtAhPLVOuZFV9OqUPp98
vgu7COz3TCoiFt2FGiS6s1gMxoxhmn69E7/d365JHxrOJIexbsjNsCRrgNf/VkRq
nm6thTyHPX2v+fmnbS4XLVUgvyO3lpio6qXJcf6mxHqqwwwSnGChY7ZiCOFlGjjq
52y88i9yof3i1nHX2Ka+6mwwsblamSW+mnkBurL8YLA4zHTNk5cwCgO/2BIvv+Ac
YOrLBLyAJkG0cS6t4R9rigNyYbTucZrlhws5Xtn2U8VzPvjOR+4HhyTZHxLk1LSB
TVcI2lEGOdjUv3phRJxwJC94z/O4zNedtGQ0QcgUxakI6fAp8nUoJ9YCU3rnMhoj
WOMfE0xWUeyX/3ugRqquNaxrfx63OnXj/3/aTwlBUwZXrhEoOL488XlrPNodClWu
4vQyYtCl6IIzZotawsEN9uuFZk7E8qtn3DXVawjEKBpA3mnQ89g+nMaVGtqwfPDX
vjdKV7ezkcxoV9o2CHQnnLBfBrPwpX/DQJ7lP7XVn3MFLjEvQjK8dkc/thnjdJKm
MAttVq+YQ+oktdOdWwIkAgRBV1W5c2YR2X9M08P/+spWB4nEOA45N59cDAatYtPF
DIlLI4ACuc7M8aWka+pC1qQbnATwFV16Sw9VkdInE/KGRKtk9bCnjn71jA/NGuPT
1aX5FT5WVuS6pRQOEl9WHokysRWx5qu683GM7dBdSecuSMbYlnssr/7dpeW8uIUD
MXkcj9sWXM982ylSHRhaoB4wduZ0LEKQznT8uExYH2nXPdZTf1cwjDl2cKaeVmXG
wRidwRY8zrocOKY6rJRMI9pYl4v2gdIjKMEZDQXNJeJ3sAQHz8havnu0EO2zaopu
c/thVhloL+/tIEQgyBYluuNppMndp6RPOZFEf8qA6HMzseBZQQYS2ThepAC14QBm
RyGZwgRMyCcAetD8F9YhXHD0qERdsNwU/L0PCx7dYynqXBn4dmh9wj4CS/u7fyf8
osJR3V1IKT9Jk/XmZgd6PrbSYSY89nvAv80kchuia2Rwo7tJHGsfZa8ZwJZFXoD+
hR8vOHNooOtZubbee+ry8BbLgboZYO9uEihSz76jQSsGk/OeFJO6JQtS5Isb7LB+
szLwNbyBFe7cFRp9JS0rJiBjfVm69N9dd4l4r0Y8Byfb9AGfqBTgawu5N0O6LAdB
OCEZv/XFhS2tXYRcVfd74pp7aWz3apcEVHHC6GD0Ld70oui1Tg/P8FYusKMWvurZ
oNcPsbW+Q/s00vM+kFWr0oqOZctgR//BNeq8mR6qtbXs7DrevFSwe02zXiPSdZeU
O+R9NQYhMEWNZQg3e4ulOvRLqrCJsrp0PJwKvXPkqtEy5PzLY3SiKPj4u0PKh6qs
eX/YzItF9gNrf0wNVLTa2qBZ/U5SGz7dV++LsC17rHP2Xbgrwju3FQETQS+4CgK/
94k4jUQVGGtXmitdibgNyg/5Cc4nXeVFwLe7SpHzEeKF8k9ar2bSdz7nduJ9TyNu
1LsVnmRfwOMYTWKRgKkQKPgCVOA5c33pzNyWl94gL95gLKdvcpEYChhqZb0aM3lZ
o+Gzo0LefDB7FKE2ShdCHlpQUtavpDSmUyzKQLvJ2xaK/8bArmY/3ucX8jz3moUX
+JHI79B63VtDaZX5yEPAEMyoXR7JNlDvOP27WdreAxGP7xgq1Vqx2b5e0lbufC65
3zDcioCs9uHZPGYtAfV9IDVweJyZPJ6TQTz2umDT6+Bzs/E+vk4pv1UfE5/0DaMV
AS3BsBFitGcFYoBNeKGDmlPJ8R4bFP2c2N01cqCiXqiUDYPFQD/kK1nGZCQcuG0E
S3QlrQPu7fQ3c18yXvGWuolS9GxYreUAJRbz4BEBgeYJtEZISw3w6wHCC4HhFCCh
DtmTaFHAenRhcKljrF2yC0kEWH+BNmhl3qNYwseQ9FJuA5sYcdWVmVMvjZgcRG79
v/1sN9Q7+eCZhHNF1BdTmzxbEk5Q9GhhNoukP4B19XTaVzhqU9mHCL+nyvvEHBJ+
mKAvdD4P6MUQ4UOfmjkhF0GXucSf/1NxCxwy1eluQKxzFT//R2sHqjQJ3KLPhJE4
NVlTDxPZk0jwB4aywIGPyig2/ESSBdduA7CuO3lKW7Oy1kf8hCP07sMBfz+S6kHR
8jZhzlwQX/6D/2X6R2kUJ+5NHjRcpdCBPYZOv1g7FQgdUenIGxqT4hxQeW2hin79
j/I/XG6snOBxKOy/vjk3qRlDNQC6YsoT608XJ0fgqINLqcz9hHjfxWbre3EmuuZ4
itYB1J/7OFFEyptmcsBHi8CoTZUhOoX2dtA3LUgGyWyQWEcxMSpA3OtuCk49EoBb
5yj7N+Du5QQkObqwAAAThnUXaINDcf67h9SgLE8R+7snAeFP5th/rjEaC48viSoV
wLdInZAWyUooj4uNhimpUO6n5wPHkoCqGHmCjBDUYqP2K00T/2cn0Nx3hFXK3/xu
uxxbbn++Cyg3Cx+DDC8b+83HT9RY+lPFe0ZhcmQu+U0mpDNzBiR2BQ/ueO4WefAo
wGFMGzVJCMctmptQyKCLGy47Sk4vax1ZUruwT8C8595sJQQbVXZ43DiYk2oR/gdy
bo/PPHfLWEGjlEroZTR+ZvE5fqYj0gkCwH1NFO4LU4JySh0DAfs0Uhe4wvsqBcQT
v6DZlPD1/tAYOYet+JL9Iy0tpcI/012SzlTcKXgT/lqvxevz6ra+oPsNJAxyDVDA
vQAcxF4RyX+lExy2mp/27iHmWOsrORa+gvjosDm4RR94eFUOXXYy8ISAyxakdEXa
GTezeS4R4UlFBZTCoBZ1A1Nt7ySvHno7j5uqiMj0IBegCYWHqqZk5IhFdWm5tf12
yQNjXsA0u1aTO2pHc07xJPRFS/eRd5t4UhEq1ExO1itVA4zXW/Aqa7psKSbl+fnV
XS6hnP3QyRQgBq+erbBABxZV6coOLZrSuWqcpRXvAlEVeVyqUYgFehQgobaDixOf
7d0y4n/UtwY4XbOSniWUMPFDADoTB9RoOZqIMp0c1BVjTToE+ykSfr2BnlBBMKTa
wg3eBBN7ngemeHYp80UEImUwPzl0iNU6gw3W5yuyHiR8dELJ4A9DkGg3xbZWgMCR
fCMw63kOt4t3LgBgPvgbycjwQ8lAGyQU146PglC3wpJZMZOWOKq7scgz85KzbmYj
GIhKeT/pjV4mYAVx3JIsUXIKWQ9yyb8yhqMSl9PUDK4IUUll0aVVWm09k8Jmy7iW
6WeniWrC1lzCYhDcEiQ52fTM0werk3aOWINMmZxTjYfuHnVn9WBSw1Mpmdml/628
TChAurMZb5eKhfkjYTybQFoc0wt5+DzSGLzzYtAwYKuxwBynOx3L0UocOFtaiaBS
wlBJ5xAziZjew/KHUZbGFYpoBMBReoRtyzoy+NI+9hQpb9De59dCTxHBrV781Mku
HsjgM4fUVP9At8I62Xvf5dEdR9+0Jwb3XlG1OND2MTO+ZUhslXHSCOD/TrEnXPpw
T4TvschIWErUhAxXncJ85P5llUF5XOioO18nwO6X1alSakoFQy6qiBUAiO35QiX7
Vw3Hha0WwiqvVrBDXsRkJ5gY3HC0vUKg0u/fS4s6MzT01sshNYujuS3zyXfM79qe
rsawWqseqoHqZz+1p7hvIZY913kh+AX1tiZRNn3HAPTK1HWjfAHsywJgeE8uZ/Tl
9Cgq/GVemPZsBjQP6UIDIVnr+H3zNrTCupa6RJlyPrN0FZLG27dAOlsLDJJg0+B2
vMVVy25/NH7vrj/EdII5KZwJ+uKLgRz+KMNGYqYDa6eBmNMNIJ64A2tiiiyIEQfy
IsS+Kt3++O9vIoe2KGQmWCXXo/aLEOLZFpbFT6TIGQJ0PXKMXg4OIY7qSETN8wE6
kXCQo3YmUyCnaz1WfnsaQojCzKlaUvk8r31p2i4M/rZao6/fZvYQ3LjDQ6USX+MA
9T01ab6nYsJ7YJUiTtgWAcBw4sJN4MWeAPXUxOjwbYCYxzrk3zbo4RK0rZDeOf0g
FD8Cigh9Rt3HJasS5BO8Nqw+PPIruKwgWuylG4jtctFm2NWjdhxHAxTSHxUUBXDF
LNZKWE5lPMEyqu20mvJiIAMvQl8kG1oGb0f+ATJwEOHi6XuhEVrQm9HdFtfSAEa4
yQLur+hABkUSp5XXnZn9VkWw4FuE2aFta4VreUybDuoYrJmryZBJrmoc+s/+Q5a+
DE6sDXWpTrp4m3A530DsCsAGkWlk1l4RDdVwWOW0pnRoOOIeF39bGvAwmKj5dHWH
+87aHtYT+p1gQs8HmdWPEURppq7N3W2Vdc2HMEI5wS4UqK8GnnHm+TVe/iImzMvH
qkQGVJdKiJkKi4Pdg9COayfnh8qaNc1DJZ9atfdgZJUii1tUSwzdfozlAYgKi2wT
fEoPRtqOMdmyZEmEwKYGcH8SkSSAW2/Y0Murxhkv2VvV7ifW4fjXvMNB7BtVisFP
1JDwYOyv4sjfR7jBUl6vYplbfUFJbLbg4URGbMg7aaIzy55BZ1bc7nA7hidiHLHg
RZ4U9rBjZyBe324BC92+ONIRBl9z/UeeW9ZIcRdKA6xEc5ezRqUAuagTGkfW/Vs2
nFKLa4RBkmMalC0IEZ6DXdTfLdRevjDXLj5eIki0CoJrfztmhoWf16ANo3969yTR
rB90od2N3RlAlWHUGf3fcZVHhCVCdWNPeCUXT6aq/BPPehEWxg1+2NoMnqFg2eXZ
gTozk3hVBXlgDY3aVfMkQYW5jjMf1qmuel5PGVJUArEetW7cAx0A3AkQPUh8GiE1
QhDyQR5u2Maibwr3LKr0bKt0zrbLp+05AewdaeztQe2ZDaH+WCGCL5qn5TuMV/4X
R/q3jsUBAZIvNnxBQgnbd4g3QIR+2AX5w0ARP78VpItZZXR68EshEHXRJFfwskpp
mUkpbpcMzOPElf4l7faC/RaGC2dXxyv2cbdy4LwdIL/eVzMiGPdZa1glsQSPMrd/
V46J6SfTltcZ5MSFlnqDrWgRPJua9y34v0DPBflDBrNXOIt3S6IRhtrXp6U8FBPo
akIgXWnJdAwSpqzUZ99e7AuyY0gdgwN647Bcdha5kEKuOpvKvjrHS38KORxcoS+q
NUPhpJQqFLTePRt1vPxvzVU51Dp0kxNwuOejsUZOO53dtIkr4p4EHlV+EqBbB7iA
/l5g+aUa8R9jKOstwPUjXrAoXmllHyAmA+bd3cihd64OMA3qQIqWUnW7j0Ch/osG
sE0X+XLjw31f5aGLAhaFOUZzST3rZSudRlPjaDb1R37Fd0eJRcV/rnRiT9uea+C+
CA+6tNkaI3bdZp11YHNJLXzRT0KEAugCcexH4TnDYG76sMmkqImkqEmNPaRu44+F
ChKhnZrURfyZ0fjWxzdUr4iKHHR1X4a/KiMBKxdDTY/Yhrx6gxY9ShlRkLK9sLqv
Ls+Y6fgjdeaKzbYkPYXizZHPjnAOMFtYTBad7NfjSskWoezPa/IphIVJ5rSRfILw
um4a35Rw0cvCxISJOVVp0I/cub/4Geq4Rm1KlLNaU9+3DiU/K8JvJ41ZkjZI+Y7k
dOafJ1HAStDG6F87I41gnj9Y0qaEbWwBc+pcJvAKbCpujDP4KwtPkEp9q9Kzsvny
FW5dGPyn1ExlxVllVPDTFolpLmZ68ASEBbhw9DkxEi+GVW+O9uleRCjL+w8b1gqy
U+yfnC8qIApoLx9UGU9blM0dHRv+h3DGVYBj5ke2INMZTsHNbUkpE4giE7vqxzmy
ntx5925mgg8SA+IIY50XQAYZQhL84F43vbjlYhcheS/0M0Ai9OBBwsStZvo/DNSC
5KGvIKpFAS6u42t3ijPSXF0HYVPR/8CD7hH/6je5iyG/nLNQTHtuxds85PjgWoop
nmWzB8DP35ahAHvfcvQWrays6s+j5wA28XhlkGJJP4QqFYlMLhdnc/PDjIjtTyWF
8ZN4LVku23jGa3DywIjRMwoW4bTZdgjYN7/d+W88p+qwGLRYm2FuO5+9giODjYiB
4d9BwvfZUySL/mLzRvN6KfMx6BBPmpvsIUMsa+qjOsFrSB2ONvIi3z/Qds8cqZu6
jdLnQYDkQ7N33+VHYgx50X5oRkv4//tZBOA5M1EkJBOSKPEb/UR8TmFD+Vts0ScH
OEHYx9sGhYNaud5xmyjyRi+APTsncrtBkxQVOggfypqy1WINcg4iwL6Tz2nmN06k
NX9QjBgfYWycQrNxjl3iZJlfi2kcsPqMYrurgmZL0GaXYGcHz1EXd145fhDAdV60
nUey5MELPY2ABZnwP8RQSXNj7wQC8HG7dSIVqiMkVTtK8wDK2zIGloANW0w9N3iR
vgcwlgoXrUEQTTMKavdGgDt7CF2Qsn9FaOA4YT4eXTBot+J5LNEKt2LlM3JH3mZF
gVHmHkqt/dFpGv2zESIGIWCZezLfVnZ1HhP9i/Cnjk5kG/NkMsTNTIRv1VpLPNuv
gcwE3UfUaVsynP5ck0Mc4jDBJtRqljPqZY1bNfvYSIevILRZcjfB87oNGUkIF6Vj
wyb47+gWxj+XXedDxiOxe9u7y+IHHH8RZAxdCj/ZG4xFOQpfiSC/MrqSYMtlmaOH
zsCbaI8lV5KV4X297iMn04Fx/lS0YfrXxj2R1hiYk1ZAuyGh3SQMAFXFpgSnPeMX
GO0uKZqLaAIJn383iVBlURqJzgJPOvJNoJMuTLuEU5hGgmHZ21N8W0vNjPBWuqWj
goYNaXZ+NZ+w2WLyKBcmY36tEgaymwLnvUE5Bo/0zTODiwrmPY+1bLC+TPWpcJuZ
6OzW9ozfqOeeKcpDQ4XAYNMRHWlV0H3d9BcSmbpMG4/ebOFhEFENBl7Dnc9q/eYn
kekGs9IbtJDVJkq9ypndMsaIIhN1MiYJ3+HB9Q7N6qFy9/q3QUPyCBDY+Tl5acVa
NTBvcJDg5QMFgdET1BA+yEZS7EU4J05Q7xwVCXFxnseX9K31VEkL7IQ9KnlIPUgu
8HGqu5vfNcL+p5gxK7Uv3O1x9SjaKdYDWtBtBhTJA2bR6EiXKOas5vh5M33pPbQ8
9/J2ccfO3uEmHv0nHN624+afjkPVt/+bius+m5m0YOdsBuGtADPJNIYYws2clKdl
0+CQfz8hIkf47pLBqAighp2/rKKJOPVq7f7nlJAH0P7rYO3emWhXwFWd+SaDwjvR
A4krtB5iRttL3mwkCNK9LRxewK4KFhkOOiiQsONXy0U/RdZpbjiD2LqXLenjv0ES
014MVXbtDjHZVpV/GdSoBMGkdgq98/003gc8CErnp168kX84grJRSUcUBgUHC+ww
EHWByA0WzI5gieLrjoXuocLSwDW8x5N0LIemfei2mW8L/i4xSsIHXbWFL9ofQhTR
RlW4y2cS730g5p3FlM/zp+OwH34FEafqpOxucEN43T8ySksS+iukdSJTffdjpwAG
3Z9lNmkHYuPm6grQlRgplYzLxvfuBFn0CbmMhoebqsgoCTyetgNIwpPENVF06T4i
TshR+z20j/dnbI2yvTm0YDKIw67hVZkaEvzPP2c5j96SJgqNlGWPS/Yr1bW/txSr
Ehwv2MFimumXdzWwtPDTW8FwWXy9KHb8lVzX5qsOfxqTmylFg5/ODCjIrwHxa/YF
liFlocNh6khuhk/pI/hLqSTUbw2jVlCo+rVIAN1QcYA9LKDdMQv5c4C/vtUu61xI
b0ol6K3QYBaUZoetvMN65sqxOvuI4HNZcDRC4bVBzmRIByu9e44cXgPJqUSlbEwo
CzwkfSy29WXk2K4ymsmgviTSWIWukm/+MsXrlmUXdCv33vkb2TQ3eDB5xA/vhiF4
EpG1SEMWY4HmBMw6MyIHDE9CjE7CMZchXFJizUvtYbfDHPEmX8GMc5toCJJv3Wpl
hCg9z6FcKMmjDyObNtkxXlAtbXABqZTTpYl4cXgqYYOaQK3wkEjRqdXJLUPpfIbz
vD208uxE/RDrVzDL6kVMOeMdHnlAX1a7vJI1z/Q/UomaxChqKMbd/bdyqmF/HxS1
x7gzAhOkk1c1Jex53UM2R0FlDh30QYPSJcOpvqPTADktP6dHnEFNoNi1jUnJbi6h
qoWt0MikVkvtUwg5etl0tfil4rALj5nV9CZ8KG+7EMH0vyb85VFC+mUjq/W5JAdM
GTb2/Pc/8Y0r24xwop2KhCENuksKZuwGI01nq/Wf2IPYL/zdBhROBzB8FsncvVbK
56cAolJDyTPgCXMgFhZpvFf0wpRZ6NA02CQoGot9OWITzAOmONTy7ZF2WObVBiCL
Dla0N+p5rODY7Yo52cCBm5l+cqHX5rUc6XGXu9iKOB8Cg62NIhFRoRbnVqNkMZuk
Q7SryCquwqW508nQDz1HR5PDg6vM9prAHnHnaa7gHXwF2AW0wEq66CqwxqLI9iz0
CWrG+2je98wtdl6bafQPVOoT/yWsFLCuiUub2QKHPiVB0kkoIhz4WWzhvHRMG2oY
kEUa7qvQEfDrvafUP10fC3RX5BlpLCjB0KEIWHKHqQvISJb+jm2wn6y8nDaHl/DY
nGH2/ux00z4FAzkyJf1rmKm/9NtILCv12/ew4/yReMkp2Bvt/4CTVYjYaRMgon/B
5eq+glho86RAPg++4jceshJxmzmqKoh0DOmjJhkr+nwRlG3cuWeHtN6Xb9dHtJzZ
fsk3pSdrQ+Ju7vTVRFx6HIZDbnbLHg/4J4j02PTRUC3o51TgZ1OhIdHlqcgYql5b
g/uKZBwOd2tMgs/zFfXNZU0p7QEjEKHIKzpRDHNDichP73Hond8N2vTK4vbXn/F+
IHmFgukDOXnmfxXh/iAEzcuUstCusOFr6OVGRIhOs36fYSi3mWtrK4HXuLXCLKND
ja2jj8xo/kubtHcpVM7HdTFSfY277/f66+wpRF35qy29vQivbWFH3IkpgU3385CG
yp982rTFnc0G5UqIrsgHePHf5AqKvhKZlWFJzVGxmnlq98Gds82P/h5LK5vAXv70
V7tW272Cs2n7odLKMCSuKMDEnB5oNNQTA5PtYRwLGUJOQ+GXsk11JyTOKj+l/i/D
CssmH2v4wI1C/zSaCUxY6dJ+vDkZj/bjKKlugp/6kfl5wgm6J3yxmPk5mIW7OofV
twChe60YbJP9rOPHEeB1uI6XLomcQcznr4Lew3CcEqCGCSN4Vi6O59ePYWWtqCQ8
2Ixg33h7Ut4muZ5rvik21SQkwLoitveHNaLxxVsNObFctbN+zBz1druToVNyUaBX
lZ0TzI/iN3qUpnLaLaYcUiBecO8oAUjMksiuBmMQFwT/G6E2XKo8CXjY7lfRfwgT
PrxZydAlKQZDnzttdkyiDP8nOvknS0EsKsoIAOn5bcfiiBIdJyaGwF7N6ZSI8nG9
GPdov+vs58UGi577uYrEfrfsvcT+IGaSabYp9tp/ympSzn8G0mnBBq8mAcmQoxpy
z5O5xVllsmJVNpjDJXzjfLDEC7s9+5TzF8DXHc9eV9abbxP3jieEeQi7j0bBoFDf
ovtF5jHXBqzTN/fgMR40TNsRas9qLQHh9BotxO/K/5RUHxBvIcmfabgCN70xt9WG
2UTaA7lZqSZWXOX/cM6xbFnbwC+ZyoWCY7hAcREciWa15nz+2yNz9phcuqOp8MQB
MF8JtDIl0LBl+w6Qc9cNYzqyY9eTLDjfC0zWRLofJM+qwQDHqLXg00JlbdY43l3Q
5nmBo4vNTnUA2zd27dPC0SPqnIs4ovDPDVyBoYnnedQRX1sHIGUyjSoV1uHCv7NX
/xTT21hWdNAEexpkt3rwrMHEet7nBwgiygGQTiOLewFdYNgixzpe5+HIB3uJVKVg
RxaNuvjW3kqa0Cdc2DhgpXreTKi1yVmhNeBoE6ZNQmtpOdDpdNf+cR2Ob29f6Ekw
KSxzDwLhNbaoPY7uTmYClyJ1YODxmuKBRWx9a1lK5+6wT1uR5S82FCuTyUnLFAgo
ViEszUzHcslM26BMzdKMxGt/N02PVI0mdRbw1lpN8ANdrb3fgQje+k4ghfMu5NdA
d8fzqSbfMs0+pDjlDU2urUz+b9mWlbioAVH+vu+fc+w9zZEam/kxKCsXrfhSHv/l
e7ZsXT2y8cM/9IsB2WIRonPej8rg6btpEUFs+FvpqkX7XrbSMO5Nfq3bzQQOqSc0
8MwQFdiXGAag+3287e5cq9LMwsX7+Z8R0Pt2kwLpEm2Ecbf7UGoYnB+gfxiC4Ssf
6w+ZaUgsR63Xo/EaUILQAijJWoT8EPSY/wEF7vRoB9Q9+34Jc6kUhbMNH5RJ5a7M
9ZzYjbKjm/fKN1ovVgStjQxr6fzRW4+6RKrPFPixSoMyZR+eQxVtKzfqIMJKTHmV
kySyKf9eae8v8D6puSJtrA4MdSBYnvEU0/6+lk7pTfIvwy7e9/rAFEvx/Og1dMms
qsKabexdi/REo4P+GG3iDNdjo+huAsppSu8XJ0/Lah6mfeyV5EJumu5S8yO+sOc8
Zw7FI8cMz54eDtOYtPkHyykq1sT5I0roZP8UqDUCiz8F2LTYvMIDpoZMV78K1K4H
GwWu45+IMX0T5LE3UJLoDKCc0AMpNKcY3MUVBkEvRFdGUctaGJw5W70KOZAiPJgY
9jzz0o/UHdOumy9VyYvZdxcam3tfk1/DSJYbNCnRAW/TdTBrcuQ3u5ixNcJIJNoC
vFB+uqaFtEWDMxrMYXGDmvRfdoj2jRb4oA3Q128l9U+vF1DhxCWFwkORbAaHF2o0
dBmallbtmEATjhx16RyxhecF+hmzT87YFsptLQXaunZPq5aSGExdtBw1VyVHKmzU
K9adSMs6OnxBLa/63sWw92RVDekB/ozyMw/p9E9Mzj/HjVpq0Zxfe+kGXCPPrgZi
KOmJC+/TlS0RoG9+PqvlO8yvUbUEDiYGy9nJDDsYBrDubVLQpaz8rs0WRm1VcZvu
K7bB7J3WpIJLWxf/DYdoevnoaQ7DxWZcK5XqDRcIzR3VcN+0lnPzx5SnF4DaoA5J
oLaVW4H/GwZOegKLnQuGJqs27wRgqanRO2/ujggiJthKBTcBlUXhvcUsEF/EDwaP
pfkWguyUdVcERMpP87V9PM4rR1awg0+2L08WJK5KFKCLla8u3RbfxfFZspJB/gA5
4tjYmf/Bcaw47ulRuXT2q+RWm1lQ7J2ksFReykSWg/hDr5Li953y6jf8m0iCx7mF
RenEN62v4bYWKSxum317XA9QRcoUzcY4350YaU5kjjaLMS61UOHq1Gw73lNNfr/M
+MfsVJyuzuNvFOrG41nwp09IosleHEEa/TYpBLeeR++ZHo7WV4faeWmvSaDX7uRR
FczbJuMuPLHBklsWRkzG+vV58sOCkkAKBeZAluYewdwGrDQeKOKNUhmQlhj4y6qr
1UxbyP7SuWLIFyrb1cEQP9LqJL7ExyyPgfizAHYo5dxcdSIcOP/DaIaEVFdt6SLi
LG+dpVIzU4p+2EL+5ElHcUwciQeQIn6oipIf3Zi6msdzxdnYa+mm+vvvacLUI57V
teTXBZDRXUNLW9AgWJf7mTDrFcchYhumtBuCpo0Q/HQFQ9l1cBwawdNFWxqNuTby
u5cH+5O/Q779yjSvzVw9dxvVBNGC4zYxkPsbH+aW7QAjx9sWGNQ9kE0dO9rr/gvz
ab7T2UEc501SK4hrJ9bNiUuGWcLyrhFAFSIcGOzmjldUXa6HO4nPiwr6EFtbd3mV
jezOrFk9RTkvC+WS3dImvE7eHYVOqZxrbmBiwwFc/NAC9mEWX+dDP/VnP4o3/5Ig
E28DBJIGPo2BYeDOEcQy/NHlp7pLITvp0lpP7JG5T8VlYGZp2qnkOTEYK8bZmuLl
/XAG5eI9/NIBfluKTmMu7ffT8FI3ytXgHUasF8LagR5/k6SNTtSYL6fZB0WbHniS
SINXiTTQeTj1ys9rZRqWMlKT+IEANDNoL19I3tsa6KzsTi5W9adaRzAzowhB67dQ
BCLrjXcz57fZaPIgNEvW66B3FRLobhgu/1ziL1m1oM1s8z3H126i+vkuf01aKCWp
LdVdD547UqDZR6TNbtpkucDOEYYas/Ti52FpwroEsIaTfLClULSecT/RlT9tAsD2
mKDvbLKhjC3DQdBMASU9NchVtCxgk/9KlxAwW2LWKVSfVRofkhu4Rn/RNOayl2C7
5o34TsUlM2jtuu0fpvdfpcaRmL9FZ3aJfEVUAlLQtwjV5xdr40MztonH/lEgxhei
UeaifnstVsNBsiq02Rq/Zd8SWDM+lTlRvnjZq6k73iFm48YIMK+0rUOJ2rIH8NQM
xkeU+nOgDYw4GJ9nHCTSlD9T82aKHKBLwPNR56iT53I+cHojQeTZSUkWX/YJjtq0
yjERkJKO8FGIzTJvO4FMx7Lgg9HsenrK4BA+p+Z2UhskmlIOvwWAZ1cCoUzw33Nk
6idhgJko6hO4oC1Dmu/d3us43PokL0sP7LcR4zay8WIzdrEvGMdGQrPnCehEuMmH
UbHF4EwYbaQT9HRycg5xHosLB9PV6w4jnKM3RrhrwcDKr+JSgGBMWctVXGn0mkyJ
iH9lbfXkEvl+CQf6tJ2wRWMXqzGmKGQuua42SbxXV/D+ZLmZuL/81hsrrLHHaGC4
HY8P/zJuiXcXtFXluyuFQpVZn/6Y6rwDoN3fBdqQnDEf8zBHeEtl6cXdDxlWgktq
hNA1DK58RoPDV6vllLZVaUxsrCn0cXOlnPQ+1a88p935C8VnfpHsiYPcWTU+Vmza
Ss6cuz3fFSsV4xEgRX/IVZ+68QUFUDJVGAs8Bg7AEHZGPfqsyA/wPT1fOx0M7SUB
xqwIBfbbeGxNOt15EQJcqDiXqhiPNStqrbjkW1uXvQb8HXMBNdOYWTCNjaKvR5fO
hvSoHN2q3ujqCrZeKHqF7qP1xi1RA17qsmweYj2wvfL1LYLb55dHidC8w/Q+jic4
RSkI8oIxM+THJiMfrTaE07hM0N3i28XzoVberUTTDvxe6bvfU0p4r1UyeYsfuE+5
xKubXyfOaEPigsBsVQUec+DknZ5ZMEWb7vx68fxBke13FtRPP+q7KBKDQCf+nbZH
f5s8XMae15penWB9v8VKxdOydeIbGA8hijNrgQ1RgKPz5bahTCxqvRT/dxwabwrW
fTRvQKT4rt5jPWlpFGIlLSie1fDQwd3Q1EFMcGQnbcTwV8iDVPHTAk53HPpp9Qp6
cHGVuHE7UfxrnT3WSWXaGPHYknbYqUfbDV8PIme9kMD4cnlwasA2gW3DG2SDLKB0
YxEEmd4ZGsaX8DhbPM21nOYUdNouRIQQkg4AnoHXu1wBSrAnM76NCceIhBb2E3ys
dxDAb5r8w9KBmW0lUJs9U/7LOjmIetpje0iOVQf3d4AasYPKN4C7gAg88Fqlcouq
vCQtom7IpYeYDLUAZEjf2jMbDRTL2vsArP6z24lvuMjX2MJyowwFAnKoK2TjBWhc
Eir8HcGNo3FwKnavmKkiSnUDG8jaQsBnLbKmolgaK3WCWqQ1hWNFs29yeQmLBNg/
NJkrzZFrxeGRxx4ZYCIZmqZCw8pZq91tn7wloHJdVn3j1EGZSY+COTiKFefCbtN5
HJWUDFFrpwctq4+owciWlVRxcAWjKfsc7bKCuUPk0QZp/rVhVG9Cy/7FcDTtgFjb
getdJhLdeSSBJwMYG1hC6ZECOyp0FguHK3JbTub3ElWkMwR/eS4wLhPh7ZywpP/w
BwsGKKDqLkuzgQQ5MgDRTtqUG0xt9rLUaINiZ6OGfKmkp5E1ZTQ60BPFqBds2/C9
/Oo9ZD2002WXjPBVYRjPvGzoC6Ae8Xh6acBuqNgCDO8VGt82HZYUQLsPNAZSLJr8
xOfLWg7az0n1WD9DTejqgQQah1A8+c2c+PBQCcXDd3WtuUYkIOe/7ZoVgWgk+Lwk
8Lk9gEMzGTKn4uyHnlQVzH5jv1ZUcbF5iHwSImD1mb6JaPSnw474itXXII3ChB4s
amti3N4AWH8plA/r3m2W73KM2QX3aCjMP0feBBzAkH4S4K2UECCj+dgAx3mWoy2J
pTR+kkLkOGFaEV4m+vAnrdqyWNt2qWF2dtlEwKGiXEEeR/xHTd92HD421YrtjZod
1/ZYtZzc3CrYsiw5VjeAL/yxmVHDsMdJqBlvauJT7Zf+ZRFcqNSsqbX9EXzd76u2
bQlg2u0pmAJ42UyVMSUFuP2mTZ2D5XSGgg9sNbWzoPZnwYQ0jXrFhsIM8UVcl6oN
ZPcp1brdxFhhWWi5biaIox8mc1Ruut04Y0/n7tL0zBS4el3xhmEeT4Y8DEYqBqaL
WjEA/neet9M1VjKtQoT8by+h9p/5/Zho7yRLyKcS4YbhOm1o1dDJdeWxRgPOBhoZ
nw06A8Xd3VKKfyh7Ks8rFhcDs4uJc9w2p54uZeNnWCZ87oWgHZAwlthuuiKwJqol
d3iamDmvVbmYr/xb+QCMLsydA3sYa0kQkrZQsZoMs1wZi6P1p0mx+eJGU537c6Fm
kMEtx8Ium1Z8I1+vJTqOSpg2LsyotiF8cbvaLSDP7Ub2AfA7uRA+zIKdOZ+ElcgN
YlbnP5i5gHHq58yPAtN3vPQDOluQRbeCEVYsP+gHJ+LS/RBovGQZyHkNsPZquUA3
uTtVgqI8xkNFJQl6VAodTqxNsJtrdpyjI1gkFudABXHYVU/PPlTVKKRwyAlrAnJz
OWt1K5DKH9stERtz+kR6VXlAzuYQvFrVYSZ6IvATiYtKhVjWiD6GwJuqdknrquJC
wbUOLl4kb80z4nzp+/MgsjDMBO0hzPK1t1ZbQLt9S8aRtoVXTwl2jvqwyp5gENRx
ebkfqzkOKLm5c7hjOgrpOUM4QycZDZTfBlAGNxlMPc51pSg4KdI9JUyCy9lFFqPs
0Ymngs2gW95WblxmT/AyKBYLARK3jMF2jQqL0WzstHWuQmyc38/2f6M2t8/wscms
b1iMenkR4SY2pOBdfXQfGQQxBsXos+Q/p3gNezQ/o6mdteaxzUoCwFWkF14WXv83
iUOAOlUHG6Bk3vpa7OC0NQeCy0bMNUK1CtcknyYtlwWrH0+ZaZ//FM10DkN4pyU2
JhNe6W1APjfXr+XWw6tu0tYm4tHb4QxKjmRmH95LAMcFMUTmSp3cuzHFFmTCaVd1
9AAuNUswf8gCszCFafkKfisuJwQRz7Dl83NLmv4hQ90Flf4tWEdOMHBAiYvPFawH
wvHE4OGm048B7ODQf4A+GiR27H7teJVHH5zrIryQ7bqivrtPAmVsfBVDMPu4PP7Q
1SuOT4a1eehlKY/Amc+qsBo3qQN9kD0HZXY27fHlkBv+cMDbsFThMMrBe0sNzIa4
Kp01kSnei3SupHji6ZUN5QHfg/OFNsAm7t2Uq8GTzYfFp5iXx99bzcc4wgsmUskT
yX+hIa6NZRKG5fj+JEC/R9iB4Tw7PqS/cGQoQuQWx4umap4036plL8unvrnXh9U1
sPH+IxK8irm9BrL010faXc4L0bsaY09aaHMm2jt4QXoKY8q6I77R0laUm7ivwUiN
HdViVqiqIiaJY6KQW8D75wEKYzWHWFvY2oINQL5G3UlfRyVXv21U8mRvdaJxmMSu
bx9ywb2SGOSE0YizfT8/0ZLbAoa7qNXo9U+tKlpWJ+1a1pgYa2Lj00vsFi7M/6QC
C5WVEGF6DOAWKH5xO27vHFUs1BxdFWyRpZYQ5jz5eChrGyzxD5yHRr6I+kKaANFy
ws5gharD/22P5fOET8DhTecJc/N/YhMv789mLu3wjLawq69wHJ7KOF95pr7FW+5q
gxBLaT7wTH4A0Q9wzH4GmYwWstYw4TSJs8iRqLZyfigozrE1/krEyfSXY9s+kaNG
yFBOh8nNt6RaLI0Qdy4saanJye3NN2j/4rIrJaHaYi4YC/viSjDj039xYn9U/8Rw
rnmfp6h4oekNPAXn3kgvB84K3+C2xjqggZjJx3S+uut77CerKDc0JJ2P9gGVzicE
SUYh/0JvPAz/uIYqEU+buZ5/5oyxgCR6WPdR4g3o3zPj9mxdgynxqHSSUj7qkmKZ
SWS31sJjZOYsjoqrQ201L/HJY0BZ7PmXBi6i0UWiJjSiKFNYr9bcUIuuod+0BNpf
9Cwch4ovaQ5ayczCUisWf8q1OnMCwShgJA1w/cfhoHeUEFiwbIkFqyY6OkJR+yyX
+zWhZPD5gcEVSOE5M2NQFFQcRZq3WX/1AqRrsXhQwdd1tFUIyW/E+LIn4GSnB5QJ
07lVPcuunC2IWomzuacPBm70BI9z+M/suc6pfo+0BhiKrYc5Wr6QBB99jVb6dIYB
d5kCGBes754dnhYaAaQBN7ZfQSVhdwPSP0U0ebWE/dniOV6bziYmCR4nY+KX2Yut
uMcQrqnWYo3JUmCr+a18EQa14+s0I7TNCEHpzFVOnGiskdTm9fwFaAfnBuG4ePKG
0t5z3TUQqDku8uONPCnJG/+jCgBMSrEtfLBUVF+8P4VX//jcPovOcp2Xn1Gv3+1Y
xITz0OAHkehY0/SsSXMeHmFQD/xo8QEMIK9IrchYJwsf+GnH8z8oCuxLWmUCZPcN
0M6Hlv/LmGy325pyzATgy45ZUsOT3tx/Q3/wY6AjIDcPZNYI/6VjTG72oJjYcL/e
FsSbnKpiwkSdY0UMV5JZXdxbvDaT/JYPlg3H6XyzpTsY86CRUomC/JGZZ6NH1UAe
WW6Mu9b/2FxurNwSlZX1uO6DWu5SbIO5ZiFq26zhxCZoj5BLR1N61+pxAA9mvM4+
93KGsqBLI6ihVG2rNATGE+WJU9TiiCEofSRMzLgO6YU8ImKFLpGcjtQmC3rhrP+8
FPNWrSI7Cm4vdH0a1Vf0I8E5SaC9zxg5VGKHTtvZfWktko5dD/u1TSo56arpNUkH
T+By0ChvEke7EfbMwfITMo0IFOFfSE9qKgXD0zgd3bUimLQaxJRVmXNvOqymlwgZ
vI665nMvp+ZY+94x2GzwYQnSRZJjRLDz2PAsTJ6qQXxszM1R9b42VnJeOO6uBRZr
U5OFjqwvDQ0259HqRtAY01NPZlv6UsCcA3YjSNk3LB4mHH+2q/qB6qSoLYO5we4c
Hls3xqPotFE4Qw6uUSN812pbfSsCVcmptdBDvVgvPMrzyt+0byuv/WSOyfS6ISXQ
1VyjXu7cSSFcW7rFpPszz+gYImIJ07HMNSV7o/mjlJh3cGlqw10pRX2jkIDoQhF+
7BZn7CWBDpT6sKrRvBVu5ZCOk37SPsld2pEuBrqn89pj8UUO+Y6p83J/i9FwD42W
u8ea83OF61V6yVD32LLY4yoqO2au60vUWDEGE1wPsklKqUFJKZSZJIo/N/bMW7ip
xKb+qUL5SxxJD3FvYSZkOie7HuUaGdzVoY1LZDLEw1PdEm8MtJIt2XvahRymnEXK
VWOuxnPqgNBJfHAGUc3n98ornysnUJZTLy2/FXpu4R6RwYxsnK2py4Yiht7XFCUq
pnB3nkFQsHNTRBSuN9Pp6m8INyBSLrRv5vJVpAI+SmVm83dJRSCSGTJJ+BQx7Vuc
fdVWFvEnNNnjaREJpDPlClA9O2YcsL7RgYC6goSMUBrPVnKtBg3tdQNnpXBE28el
BmrD0WzHqE+x4FBO1a2vMS3XgOlDNtHhBN+5rJDoWc180IdL1zMBmDb9cNBRsqDO
CdmzrxluzPvaJ6C+Ek+rfgFuUT2NCklI9jAgJh1QI4T468z8yN7Ric1rLdNC8O5B
/PH5ZDVP8buwGp2r7spRUpT2j222FN3Jld/gLZ/D81Wgjez6DFWq6yvwcd8CNuoS
m3lGS7qDYxAU11jH0y9LL2mBc0XddMVUKrLdOOOklzZROxq0rYuC4GxJirpck/EZ
yXsby9qQVgNxhY9wLyqvJT95ZQ9VDBN2jeDjtP+EWyi8TBq9RsuOmiT62nzEXQNw
E9UGDtWv5og2aZuIsQh5FB/dUsNTDsSv9R66XzX9ULCuOtke0cYBJGUtyGlUm1sm
gq5YwoZwb/VCJeEEYg0QCsFEYozA+9lTqDGuhuDjJcAWKCfGlWjSPwVwSGuzTYXc
6WJwZDXmW9bYnP0XpEAp16tpqOBuTknZYwLZp43mcEQk9stfSfaHWUHiTcvuqhUg
pumr2ApiNk4g+tatvhy+oTyRZ+irgbP1vxa+eM4nhIFtOc7vCvChLMjdGw51TeFp
wg5b5/pMpoUwx/YFTYegWZRLb6r7p73BIfiyy1G/EcfrximDyY9T1rPFtgY3R3uq
MGDezfLvSJTsmZ0Aefbma34HxMiArDl0CgfRAx/dRfBAAML2SBGDwe7y8QIc6TbY
FX5BiHYxPmZvbl2Ckxs28T4FnStOj0bgBYqnbIYrkfMjra7v9RLquTCrbQ6juTo8
tp3jGdBuJ1jsB5Z9RUI5IGwa5u/xVImpeQQtU28/sHCaXt1vRZyrwmSKPJbdBye+
cAqvys9mN8rOJ4116ZHW7UkUNuCN3Uul/JAasFt8g8VhEqM05JiXNWk8BqtwvoB7
GnQZDUwB1zbqOZYtok0A8UcG30UaV6ZG5NHdxuoug+3H8+cIWWIlW3twXXtzz8A4
yeZ1mFK0K4VTYlf5lY+pTJIEq4dt2T682VX3QJsHMzQnf8R7kuQOOWiMJYKvQTq9
oBelCLgtVisQ1jFdYmHQFnaixHqG1DdEBLuPzuJ9SXvnemdpYD2+8OgLIKSx6oxO
WPmSXbaskSJavZYW1FR4Hj1D8Cb66RkAePOeQblrXjm7giabdwkLATp1uBU+UdB+
yKcn0fjgN2waXYqKMTVvBoMD3eQ2tuzUX+MFedEkA+sW1W8owc1veuvjJu1eMWIO
xggdqRYTH4R7KLCVvZ01xCSQ9oyLzyhfBm/gPhPEMehuc1sfdJ+p+ZI+UfCKXA56
KLkqy6c80wznCdlva4fCmA==
`protect END_PROTECTED
