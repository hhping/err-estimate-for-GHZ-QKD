`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hzA+rGvoBymsSKpYwsQleXmw3tB627tL2kZFHk6UodMDo6hxPTXw5imW95AtJMFY
a5Zr/kzZi5qMoySf7nae67ZK/J+cYhfLrTFCSLVQVygK1nbCV2ymBNBRJOpMpPDH
ApiY4R4SBCkSb9boK55kyR4nrUXDnnd61KMSgbbk1d5LYAIX7Ixgq5ZJVNl90UEH
mYgCu+SGOW8OsWaubqoL7PHicfwsRu14MtfSeTp9pc75usrNtaXKm8wIHHP9SjKt
dzIufbeR8hQZe2X4QLnpHnZAGPHPDDL1YNzLMANlOr3/UmP4ZwE65v176B0pT9qP
GIAmeW2aQn4CCuuqNXtSQu3hPNLn4inZ5xzIsTlEw6F5q/EPBESWr7SN2OON+9c8
xsrWD757fcXiScGZDMoB3l4YXTEbYo7oS3bFPInpQc+3ue0l5FyuSYxVKKD1urqk
MtLWo07VfuMQ+E6ch3DGLCR2cHqRSG3k4sgoz0JjqYDby4wmlGOBAQ8Ahh/yTsyl
iCWXIj97Kzu8du10lXfaEg==
`protect END_PROTECTED
