`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lcl7SyRaVRGGMR6W96G4rGLnSD66VY37XiTgAPeET3jFeydQaG8IDRYhqyn0UPca
eiAFJiqTMY+FSf1QSRO4kCtk8LSzTFwDZ3tXpaB14WZFchAwxCsq7GF+ddO+RDoK
W024AKzrNzzX+ws0hWR5CN6Dfb0kMpMiT4deWCRTLlahBNyCgrv3svO/qQtegKbl
Vjvgb3wjgz5t58w34v779OeHqbWeC3U/w/NgBYjwbBBNjEBpZ0NuM0FDPKsW3Wys
im8xyx2WLUXfDDLsB5NIFLioAkzAf+dZoTtHCxWNiV7b69LIzEqLJtIPybLJlOY6
+7LGqwZZXrRic8+3y71/JUyrMlacFpxXM4cMyhnJMsIrfqTMNslAcvs9tzUkX+7K
446Bo2tuPSEf+UWBsOfWfQ==
`protect END_PROTECTED
