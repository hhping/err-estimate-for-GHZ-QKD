`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y76eEF//71vtjoVWvvtBkoEpeIHvDP1lBJqZqLz6ZSqXWSozY0XYi34HacBt5IwU
ucUmPe0t5Vm/SfQP7lE1bE3Bl2DogDVCV3Ia/8bYsk79TV2i8Um2xfrtBiTSqPbl
sTUThI7cJ2QX0cwz8tVm+7Nmkl2jIYZEUMHY/LS3jH86iC51T7rnECJkKhsgFd9B
GK1C+wiDXkbfwJlM8GEyGWVom1x07zYsvMBIrvYub1Jn/dhiiafK2he+s8NVlRup
GVBeI2tc2zZAdsSiltO7X7BYwBohpa8UtZiNX1N62JJIeFefwUAtrpdCQhBpUEDb
2WcYesyp54T1Ns2pC3um+JJ6x4IMK1TDUFnYyYqMsQ3dvapbwAZbAQ1/74QEOcrf
UhOoHwxVBB/K8RWMrC6v/NzY6qOD75VfeoJr5HjXQVWilHwGDrwPIb8xyiNONDnD
qViwMBljiDlxTpq8mwQQQNNUIswSIr40IaS63M1IVsaF+2yf7DDPOqOrSzjEiYWM
UST0Ml8mMEZu37leaxQ/6xl5qDnz9BdWpZtWrou3odwdnACpp6EVB1iLXcevaZtE
J8zewZMKHYDorWWkVLug0KCXFfWE1uO9i/JAM61lfCzvLVW87qjE/wtiXeLZe34/
a0ECAvC2QjSgRUU1Ul0wtvrg+jK03qEJxi5YNAMKg8m9JvX6M6NrX/WgyG/sU4Yn
LqQT8io/7sfwXDrwhqyBFCecTYNSoUOCyi2KkJzowrUge3WOSUzXbNju1QdFwNJn
LTqLT4uxQmcU85WI4MwXwucDZHJFxvs87rLJpvoTSizeOwxWA8EGfSCPKFJYOm3t
p6NFm2xyoppBvUElQ60Hov6vSw6CWQmxxEV4sMizcROw+mlzKCDtJWe6icA+19Lo
pLN3pCU4ekgqr3AduV/0vDoqz+HKR2x094Uk/REhnAZeVVnWkei3CR0CWNqSz4bh
0ud9Z7vD+Bxo2phKBkF+4xaiIuI0/OD+U8AFrDaeUeDbzGOJagDLgbvU2FVIAzSW
lgF8ugWNqqMFdnvVg9ifuiMU/xx/4F9sj0GiIB4RPzFiMauqUNJHEDAo6S9fYx6n
5NTeJjSYu0qOWpDsAkdthh+DBn46u1/DBERge5ycB15A+SBtFGwcCm8aqCscmvfn
jvogqtKXVSqQeHImL2wgLAUFyp7oHF0QsBtagPg4NG139xE5KRtnlVNYR3ybxq3Z
/LW0UNaw5S84vPaavAdbq+jkSgX5fkHbeoWEgTa2ad/IvFZSVsUzSvCqxhAwmy1v
Ufaw19mqjpsgumbEHP/6XvYua8lTDAyEq5BmLZXlssmn7hNpGFbB0WrtVDg3/wu+
/esqTvZlFB2PMfpGZHvE4V+i4WDNbkq8SynwWx8OVpHAMMszrIOqHDY3JgaOrbs6
aNvTMS3dMZdZzjgC2BklS43pCjIW9aTS2CaH2cYoeiZMgVSQf2vvTpzHtZE16Yv4
akLbLr8Y8obAYkT4Jsq9fQ4N17YqAuE5nCOwU6Jmpi/FqFDh3SnspWN6nhJrujZD
BflM6M66LcO1QDaaCCqwhlU3BeBokaqzMYrf7puvzcwFFtq5b0cRXdtW6Wt7hCoy
UxusxZP6LRtQC+HAn/GKRU4Pv0zeeshuMd0Bbi5oBhEWKjbCKZmZGaSVwf2eRo4g
/poIWRZCBuX+lnG2XBTLrsq+/C6IyP9yxK3pnT+4WsC6CCEStQPnO0pam+DPfVCb
SKkFkGsnwtkb/fP1s4osCUKvTL/BPCxRNxl5bqnHXeAjeXKgRPZG4EzJpAIdEZrg
tfLEU8QBh4TaD+3HsQyEsEieW0hBepvk6oPOPZ9ohDJ8JlGO3FznkpMLwXOvHoL5
XjEA5xTNmkKLzzP3TOV2rMndd21lS8SXZecvH4ThbdZsk8RI2+M8a8bKj/5w+Er1
ve7I2+UbRzd45hyIfZkvJNiW/K/IJuZ0fOBTSnbMAit4OjAxqHJE9z6KBuR30Iht
0dmyX1OTWKY5UBp8h8htmGnWdabMFs5kwv1oBDdHxKvvJBZlQaDYctwavD1GHdST
xlR9wY1WLtCa5bYIJYpRzFPQTV0XVFydNUtYgAfJQjjk9mB81NWlWEid2zTYXVG0
ndX6gob7GPYCfonEAgfGPUxIaQZf6uOIxfd9FPoJjm6J6NY7q3j/RZ4Stqo4Ob2M
vce0w4dV21ngFFqb6Qm65sK8Lo2lneBx46JBCkhj5+T4QVotv9xD/TFZtDa62IhH
7l9v7nIL5rJqX8W83ZTc6qf6GyHjQJdl9zPVe/UXVrRZn55yge+qZF0+ilCsDAr2
RpAU1krYCa2aitxF2Lj/BWkDIkTmnfr2vk5apX43Io1jx2CV/Dndiy0ljVvT/IWU
7YxAwTcOZcSXdLyzl2FKAX4UVI4nEx0YyujDZM/sBlvtQlTmo/khLZNMQ2vQ8/tQ
CvVWXzJUdk7QGEIfasJnuD6N9n5wVOWrvb16lhy+YR6U+/T0qZPAvDSzw89SiPRx
6Q6cKGjVhb/uz3zezVaMLK0PeQ+IF741nb4MprtHSZKNPTsqk12dhf2bX/W7f+v8
YqXpmFr9zEHLVnSCcC4tva7M3S8XkEUW9zXIKAvyp+iknS81+eBr8NFgPlsnAUhW
SWgvO6eUqBVpszkKFBcj0/PrLOGvnIYRnW6UQZjYJ67YHmmBYSDET2WSNUz472B0
Gccq196VaohowjmWydClE4hfxavOxd7pWPcafFdhx5EA4SMhsDZsFDqkcr38lNgb
HxQNwQwcXCuyhEXrlyt3g/l256ofzlCVVlntdMRbUCOmda8juSJmeiUYUt9vvjgw
qqX/DtTTNV6TWiEoBSYzAC3gvpS4ICrjiSvF90eCTqXkQefurf/WdNkuX2UzrPBj
2DzgDpUCMd/0M63DPqWI2zrpaRGN3TY4GECVs0eJ1Zv2ZTdArvXOSlTHF59kPUnV
hcIgUiM5uf1rSxq8gB7jDIS3sv/o+MUQOufZKltkYKZqqgWIdBNM38jllmc+YHlK
slstJXxxW3ztUdcs8u2qDLyBRlU2z0pgNSAKhXPVJfIonw7hymT0Z0cbgpQz2rBW
jc0JuX3WU7nb6Hr6WrvC5EcIVzkUbMVRTg4HoeVBTsAGqzAme8zBqUVs7d916d8k
B//IPw+ghAhJ8GRXVVfIAF0J9BvFrvpQOtoF9eCgCMRUi0v1+SaxG2E+KysTgC78
W9kvlSI6XPsjM5koTfQ7eb3rUFjtMFKW+HSyuFD6DWaFe/Ht0odjxFNi7zIv/xQ4
I9Y4YchL3+9Aatxb+NYfWU8rlALEivxUJbjQe+8Slq15i31b6LFxDDPg5MtjBTn+
rgTZRJ2U1vJW86+OsGnG1IP8Re6wG7DpQ56yw81UmbZ9CvYMEW9s8oZjUqxt6m2g
7uCPrwuHWvJ1Ptu31H1vKolAC+OMveHzYxrdoyEa7ILD0mppSXS/UaK1ODIijOsk
TMUoNtsumzp8dyhqAlP9Q5HD3ewqng3kiLkW/5C/e9z1TMR52O/lb+bjGny0Vs+y
LJgJc9mCTUfshS+i0KUYzNZEVsiGPjr94V9Papu/0qnjElOWeK2rE55aqelDiw95
DM28wK6i1rrATnWOHxN7pwA3EOCjD7J934ZEdl5fZNFcOTRYL6tq1BYUNYm1upkP
okNPbbwyQwJVfYigwD1qgF7mdWA9+GycK+brqlpd9gOj/VBJXGKuqjRflN6m8c6E
7QD4rWk8Zo5bM9u7Nq+vSQSTskljynPElNmYCcvIfYDRQYkTNhe3SJI+1gvzaH9W
8b/VNr0R9vXc0SkpVy8CruJWlpsZc2rPlqMAK8UGj7FLSYRQKEG4r6hll84aKB2D
vgAIFZYPVlspD+j5w32h5PaGWuLIQlTBwG4O1m1CPqueFImi6SrxzBrvpvXwnqZg
J3NxEEM8eorNhQfazvttn9Uld1h1WoNtAUp8wxDKHFFFW9jvXaP6yGawpVUszy9e
bDLG+eJ2Fsl1OdIUcncIO2/A8JFAYwGSe+/hk4Df3m+lNi6rLYtYO47msrW3KQO+
JmNG/qN4QuLkDTMtlA9n3O95QhJIYEK6hkWv+iDo8BvGFsDLcMrD6vxU1ICOARO6
NuZxyLhrVGZfbySY+XEHOt8ipMkgi+csIxvj+w1VRRxDujdj/GoAvc9aV23ncmLo
1J0WibNPJL1JpfvWqBfNNJWI0Ahjf9VAj0bhvICjfVn0gfzfxQoKiHMX4K9MxOea
f2AOV4gtWEOY7aU++GaLXNOkzBjMP9IyCqfPOW+NunfcHCfNHBB0AFuOH/OyXz62
hFePTN2sSwRKouN+321VJIUgLo4ADlCX9RKkFaH9SGdIar03NiDhuP1dxOfDVHtL
XMpMMSzT1J/RoTTr06Cm5z4MbaXmAD/RFhwiMdW+2DO+3LHJByNy1apzAC2ILR/Y
9I050c4l7EwX5vCKCAhAZROCz05b36W1nwN3TQAEt2h+Uh98Po0/sXz7cORSTayp
Y14yAlVpEUuGbGRPR/k8mnwGs4Q34bGssiZb1M4dUls81C0uiCGNIcoZaeMYPEWW
FTF127KMyMCzwYzmit5A7nGZZomji6zGGdTGV7K4qAvuUES8ieCihfyWi8M25IFa
c9Sgl5+BbcklYGvfDWppK83a4/UGGsP/38N0EQeBZteEWktfUQGrvnBDDBdnnVGC
+F0n2WXqxZHwn1/bzzC5RSGteQ44XPs2EtUHRzBjZtHhrMHmJzBn274S7FrQn8R6
eMuOefn2XmvWTOFrrNwi7X5oGgIpcJnMSwbzUAI5iTxZ78Wcv8OyPGw/o9Z0sAtt
3v3S6idqSCAGu7/pIfPDRFYPYJOXqhf6+aX/WeNapz6Yrk+jeusMfQhyHXGRd2Cu
zdQ2Ga6FiVJHIGzSA/cupd9dDaV5FlauaCrJQkNlJzHc6k3mPsmCM13TvnrW0ygF
0tIWAMX7sKOqeFjVIP1x7VPv+vYWyR1LtGu8NH2S5+8y3DbgTXu2stF0uwALLXJj
pGSwnycmIznj9CVGTuFq3wkoN7okJ51/+mNzswmEdaHY7d+hTT5uQMIrOwFA0tDg
S5KB9Z2iwd3y8Jcwfnb3JIujhPHxajk6Hzt87ijbNB0rh9gKGAtYNSv6A07ZUn/M
kvXjUwKr+wYBeNGaNrE8232PH/AdG9f4nIBzcnJi9ZTGdicUOxhHOzt3Z1DDWm4s
2cr6ggPrA8MfqY34ek6Fjd4lhsKZskKlQid2z3hXAjw+bGGAFI7MWlSGyPWzeO44
tXik3WPNbQPwdi53UdBLaU5mPRfifDEU4wcqbMMFrT2v3LS1Ma6L1/nzHBnvTIF6
i1JWRFM7g1cqPrCCB7nIp9SogxuY/1Jq41qCLjhF0QaGYr6aJbp4avZ6gk39botM
sHvbDrb/HJGHvzYsGqxXJZ94WKsBwIMRSVxnRM5wQyzAX2vXjArh+Gy9fwIQjBk6
0gwnjaQLB1b/FlFcMSnYfglPkizbN+h7zjM1CRIOO+ySHNy7s7QJMxho/XUj0sS3
0z1vCXmmL5aaqLTt/A+G6oHnl6CV7YV4ZX4tX6XNr4U5naMjE18FD9dOv48zQTmf
2zB3xKz/D/72eZNM55GsaTodJuIcM33H7s8uvYt4TDXKn+Sa3/si8rYpnsI/VquF
6iN8MCa/+5/E6iE3pcLiWrGYG/Db3sNxLBl0Y1zcMBgvMvZkDccTeZVjapPHo1I9
RSki4/Ena5WtMBrAqpUrBlurMChJAibrA29453n5UKTBZSOmfGEt5gorOAhzrLp/
89KEK+Hos7bN+EtbtC8CmbnUK0JZzz7+s1DU2PDDg9EfC/6vDpI3a0taXe5pYYdk
1fSEeqbdJHhEIsJifpJccYxG/09KmIbg8HRpNAhge2pM3m/NzICg+1VXNWQVK9SV
HNxYeD6umKaAxdbPHOk89vHocLpk/RHfmZ7TxxDfAcSqfZQQDc+IM7vy6Bab61H/
bvNm9wLQwcMJdSJtwu8RSpokizWYfqqMcbaBljzt+4p44jziKcnBmYYCMrzR4ZiG
r9HQgAkgqszzGrGjVyUcyxY0sSsJ5zqPIxMvG7m4/XJMBZWXygIhhBp2kEqvmHmO
sikG+YZiLMJb0TFmX1D/uMt37xTlWRzwy6s7d/k/lF7iqFZ33QH8Fkwjh3GNmqKR
CvbN6DX2LlF1WNZ/unUMuOD/EUqZCv8R4j1FAbvz6/U7cmFgHCk0yC8z3FJYclNb
3/9uZjkMEdbC1twAMmfhLWFie0i1j+fk/SkxGLtysSSS3sbqYPSjOrIOisKnnkat
KL0DSdB3rNtRTfxpUTDDgDJX0kMw50OElPhpu24KCm1vcw+LhgZIL6qGd7Gv+J4C
dIS7plnppGNhYpSxZ0kY2AC1BCWO7NgAVym7391c2A6v0ITk7RRTj6wpXW6fwtoV
PvYcqtSPevXGxhpmqgzmxfgdTm4KquaIc2YBx0OxRNuanx81JLyBORyjPtKItQKE
wSomCnVQj76zM/yYN2EkyrE+wobdXz0EPSRBy5jSEAQq8Oz7A7LNDpOrO+Q+2BJW
RK9eDNjlOXL/ohBO7c/W4ceXiD+RNI1mbmAisxRn3o8pZnvFgdZSrRHxAM5rCes9
zIRVJza88ZcHfhdu1WHDX2VXCZI711dkukzxF8NmX6wOzuMi5PPRC4zcCRxVlUHy
5anX/MZv7UCdSBcCvtWzcuf+nE5/615H26b+noc4ALyiKlcZnIpEUCDPXXcN4D30
smstsaRgWAionOXdEJSrK3MdCqR9pWmpwWY79zEjWR2aCrsg1qYsZya82TF7ttzS
arsms+O9KHlc8XSTVFzdxuL4e96VLQaMEahecgfjNOhhqKaqSr2sZqY+UUXq30tm
D2rGnRbm3Id2+2lNOP1n7AWdS+nEytiRNFkISIYERZRvfiiHEEUhmABhI+AiHKtB
FclBnaQBXpVxwTkBchkAjhsu8SIH8fwevqcZNUeqqcBpeEAAbWcemMQDIX4YmoA1
cq4fuPEW35GOchOlg/3A80HE357gGrNoXt1ZQtwyq43VYRMfPDZtuff3P3xHuqxn
gA6J4Z58RjK2vRah6QULk/cOUX/XTd+JtAvYvlYNbJqOthqfx9QW/XxHfLjn0WHT
V7OKkt/PMI8ZxyOsRzzuaX03fY0RrRWeTP3Y/sX7OQDQenRqQMOrHPm853BhwxcK
teLM2DzOSctxbNsAPsAygxL9q8TANDABdFAlDwGlTj+I2iI8JLHEdwo8JwoorzQp
QCv/F1FDRVpao8y/JcY6xEUH7V7Y7D40SI/xvZVd5Lznh0TX2NlbMyxeuOUEvjeP
VFS+0sTZXw1y+5Qhce26PS08e+hzNPgniREJlUbsjXlzBVatQEvmREptdF4jrobg
g3nT0htaVRwZdgGaimjxZ7NZ0i6unS5uEkZtLhRYQl3DGmnGUimePA+bJtfoXTcG
lY8SION3yl6rkIbyzFrwBDPQCfoEJMOAe9ahIGDsRCvJaeAECWogu8+wKB90NSoF
g03tfNtW4s803DEJlwCQ6h/ViXHFTPyN8Fxvijw+a4dRnhnlpXVztnmZLNxMQqhr
+COGIEO3LfeBDEPCZ5Hdhs8bzr74bwjU8OKmhMpznhaJD5/ComYb6UIKxme4Crt/
cipBTi4vffq3lVUPkXo6Nt3EqahjGwBkEcPPveFg1CsSvzpeFLO8+yjMa1GYCFVr
FgJ0z78TMustln67YYVCGlivZKHvPebaW37NxVKunB+LO9JZzqzdJCx7wcHNj6lf
Ae7jUJbJl00kEUIEssD+RvmBNB4hzO8IPkup+70q/2BnjFvCvILELO9hpzRTLw2c
5r4hNZPkT+ouqOe07HH06dmqyx7ztV4vrtMo3PPYaB8WsaikcOvF3onepngVo8SG
/tBNKMPoV+PwPTYVZNl4N07vN4+A2MlB3jA25fQgzwTGLzWA14hOX6prmaGLLCkX
l9PFmwEmgfnc6w5CNo6cUGLpzOfvEpe2qcQv1XgCsf644EpNJI3s4uHaKgsgTQGi
zSazi3ewse9CG99A/Ilza6nl7KZM7FdqmKilHml6fWSUwQkjcTKVT2GwGMcCBdok
+tvB7HjCkamLYPH4IPbY1VN96k7BOrhRU1rryYfhOGW8MR2abaXGjcfaaG8KRySG
YpOVumfhMgIL7nkpyvm43y4oXPLTVpMB44oLJXudfbKw/k/IdU3+AQMjntDYgcpS
sOUwRA49z57tWHeGRfyeGRlGf3l7T9TwSD3OeyS1+8crc/K8VH1ZzgkpwazxzygM
jo06oEf9cfyzGG+yuc6datR9lsAxmBUfDf6mk6fd7LxzOiQZb7d8WuNZRtTNPJo3
Amk3A/p3VvFpoiL8o02Z/2fX0vflyB7HN/KvTddJwmWDsoLNBFzaGMXhhXt2IAyL
btfi9+5XbrJk6ZRXHChUvadi2cn40T+WPBIwjuKQg1BvJpPlNAPhP9elxD7SDvp8
NgGeLr+7ok07XAVQibbpiG9UPUwrXM4St4YSVBwLBbKou53KpUR6WTYZayUDHZ6Y
lCFAxywXFAy8K39o758NWKcC5dbvOnWiCdE2qtj+Z/haoKvia1JidyCQPSUYE9FH
TMtpDzNeOrVA/BHB2/NMJjO0Cs+ZsXtPvXVRUgKQq/CEs6thHBOdOqKDpAIPCSlw
N786P2J93Q9Ju1Cz0Sv2+G0d083uKSyP72szvgkIeq/Fw40yvSkTK4UxxrfajN6S
X2rPGDBC+zZKRV8nIOYivCVV9bQNKkGrY9PPBYAhbaOXtOSEbMKjgRGaFiEBbqQi
POo6K18wPVW2XEw7qLmpQfuGk0vP5DpsIA0sAkdMuK8R4NEtw/UvhuYCq5/DMIKX
Ah2eZhSfW8ARdjWuXmXJQatQUvz3VKPcya1vybXV29HAhkFACSfffyLT5biZt+hY
fW+xKkW9FeHE8TSU56MkWCTZAm06vPpKOrddfTErtbpvjCzSnrjj1vlUgOeaQucS
7v/+uBUsNVEHipFQBK9DAVEmgzkgb6k+4P6tZVRfxH/vgf2qGf2WSFXMd7hlJTAh
V8t26jZQ0aKXNb5OOIJ/Eq0n3RL9eSPNQnueQmoDtwze+plQxijucLrUsiYNFfo5
8CKjWc6OHZlRXQJLKfoNsxi47YlFmsCeIaJIfPK+WYn9zSUGbT5yDC3FfDA9ZILY
4jb9a8qfPvroPqejq/GJkUc1bX67Geg75QXila4csL6JYWVHnSpVqOsJd3uRYdO0
COT80iA6pu8HxOqNjtuBOK+fCLpO1/JyVJnQ+vtTDcfX5GqEp8q81gVAZANpDk2K
TLr961NxYwXbIAEd/71PKRLyv3u7aHanNe5JdTRmpPvs3cqCOfxCOB3hee2DUwnf
Zp41wUkIJ5Pf9G4E8Q55tKb/bDRIPaLVCl6R0Zgw+tH0tFII74oBBcoD3egL0Jh3
ncgysGvTD1VmffWC2t5bcxudemsRrlW4rTDZFLNv+nD6yeGuJxP7/3rUxyP2bdP3
0yB4imbnPhl6BdaweUvX8hUl56IkZmzT7UYSW8tLLUfP1LWeashHafdsZ5pP087V
4LXnbrHMZ82J8Q1hksIHHCOlqMWhZnIC6oWJMHX5VXXoP5So8r6bfBlG91U2yFUV
V6n/ZJvPOvilBSYtIMyLJR66x82bMB/0jlhlzmjWSg6tYbpCE8KgcDFBCVNJMlj5
vsBpliKxYvrZeWVF3PFd9PK+/qHpNWt7XYUxhmrtOwNLvWyQQa/LlTmCYHOY7ZBa
X+Nyj3OhOcYdSQUWMAn3eTQnWXB4BeyjREE6vIn2YxkMN7+ld8Pu3dSciY7nUFp4
Bn6xXS39HWyVJLEyWcZIp52Aqjyg6BbYkKiGn/VlB5kVcCnFN6WLxVxeX2jzxpNw
ILTEM++XToK997Auy+H3aP+JWtQSFt9TeI+uF9/T0LWcBuQOe5cljCicVxzP+1mF
6TQmyWx9KFpoNFrsN1B8EwYf8ak9WltnEUy/d6LohI3ahB6cFinUw8dgQs1N48hb
VU8kHgd5o22Q7XVe4jkgCbkQB0nDn0N0zp6ZTpQMasMxm/w6+4RVXEpfrVC+HxYq
L4VK/IJig8A8nBQNk7jRQrlCbMfql0hrUrFbMBr+WXTNmYq+a+R7f1EEFnDhDgQC
PXCIj8+Cb3frW0R61+6tfC/vFShGiGf2kqrMrR7F281ELgIz6VozGk+jPhPNwlyD
vbwLFarFTKbT+GQ57nfS5wu2k1adMJB8xZcw0P71cX7WgYgHlhtC1v52oo6YNia7
9qq76AbFM+CZf48W2Jo+4NzKXDNrwea9gKLx10sNk6LvpI6CaR7wXgRvMQrBUDzD
1YxZzMdx18fDoxjsEZIxXw9bvN2l1H9tytFOfhg2Kw2Z360CsQx6aQ59lkXVBQ3p
ATUe7JMIWSyR1vDnPg4yQSnZ3g47CIeTO8XfOaKd8i510d6nAOJRA5gBL2ZNCbVj
kCKluTmXb6g4DZWcfWQNBJo+EjafequeZRaSXFlh4Iiajn1N5TjK2RTSWWS6mJAB
bkRDzfYvTW7EeKxokuJXgJFTuwvSm6LEtZ+cMBnSpHUGX0s7GSMXyvLPF4DPGzLf
uD4HtcqEMX+QBKhYjGLjBj63QWtiMGBjUEEx8s4mYCzL4q4L7KVSXCAphqwYTJe2
Ju2Zk85r/QXaZ6lViIFhMS2CSN1uy5QG3owVvJAm0IM2pL9GTdw7/sE08sFI7oA/
qyvDSuFvjLqUGouI6JmvgaEyHe9dX4KQxClgPiSX1Fayfznq+yfEDkt90FK9Lu5M
XIpdv4OGpAL+x9F8hX4fIiDjlo+KaYe1FfUyA85hAFcqp/AWkfuvnEdLy/lNjOUi
GNvghtuQixfnhgHNKV0JkmX9i2i+uOWn2r5gEaV1E/acdrQpGRyZhmMZHgVXQ7yV
zl82deNDaKM+4X/c57FSz7dvlCcAQu+udk3WxbyAx1zOOkvRcTCIgZX2Hgo0uYPn
fSlzUuP5XhUfkrYWYwBVP/aLAYNb2kUR4Og7/fLh/P7I2OwE17r8V8a9WVvqrHvY
SwsN+0m+3qVRyxnXUHDAcuDVcdH0hmKuyMaUuzdFZW5Z23IKkNSJWDPkJsFbqnhf
psK7tARfk7Xvp7UmgEriBMPqZ86Zm/79uISWvkRyxhVL4kckbqu8uHlKTHd6QvvD
HKHGRE+8szpTe1/OUvVG/sOOBjq2PP1UaKWSj7KmzSrUPvgDaM1jK6zmuWVIUm+P
nX1u2XGmDdg14acVxtSyKxuQravxUJVk8d5Skz39Wd/nVtTDreTjh8DELyfg/CGu
h4i58MkyX6pDNA3Lokl9qY3S5WcsICmI2I9Vv0R0T73x0slFdE5Awp6p/LQApTH2
TIBfqXrkrQoSw3Vb1PcEqhNMoXojUDRNMm8xsSCgeSFYzBoq17OykvRRkMUoZC1S
l651y+YGbduLwqloUPIcg8ao6l2jkC5gPrQNugO9XKIrV3C9YUrO9J3ociTpZ9Tg
x/EAoJcpXBU+tDGFn8h+1yjDsZvuPm/im2k5jjoZDrcGUEYXoBXElAVEymt14uKP
fTcObN2+7/pHHuOB+humBnQCH9qpEHTJDbkCoCeu5uUZ5FRebKJh/zV2fhHZcUJT
uqBevyvalhHDl/0u1hZpVGN9jUMqrLmzO/fjx5AIes/AjffNbzqasbINBqov49l8
aJcURHNEqpWIpv4TFsM+uLKGeIlKVkhDQAgLnvef0UVuoQ2957CvTjynEJJJEurq
I/s0lsCU12lzXvHPtIkBMwZADA1tRVeVS5RPoTZXb1MGH3DvjKbYhK9g1WBV/79K
inwevgGaHF4oSZos9dLelZQdrCEuK2NU0nRKggT0YScv5fUILFxYxY9+wdgj1gZQ
sNRes5XW5xTQPG5anLN4eqNeuYnizCBqoLm/vZDWr7vo9qitQwitzMFvrOHFchpl
1XnZBr9KdtmP4N4RqJ3B7qSZXMQHHRBhmNaylIChN6VTlpn+fGii9rOJlS0EnMz2
HkA2Imc8XixyKpC3IBPegfJMGD3YobuOQfhebONgqUd1zl9CbLxd1cS3nAN9y+SI
uOG/mPSlnnwiEngMcHUe2sfS2HQ4KiDdsz3n0g1eJ3M84nTfEeAlXWtCaObbKASr
cM4JqtWa+yhKuX2UH4amgPduHwR8/Xl7KGC+o+e+aVbKwoQw0mlc2NjrH8YMEOiS
bGtUfQqZVT9CVdAa+VcBpzV8swy1Hsr1LA+8bk7XlwCCZZQmUa5/ME3D4yjMB/9y
8IoM6kKCbtDk7oL4E0WBpZFyZ9Yt5rdCWo0P2YoPAAdsvqi9SD/Vu4feqHtRvgd3
1Cb5CraBRaBHrt1MyKhC+zJUo+7+ZDK2ywpGluFE9Jof8nQOXZjJlwrzszE2PzwY
U463Ah57+zwYAxNH/W/nzgOhkCdNhZd384NXqbauxJuMV9sUrfMtcsyRUuPDUoMb
OK2nay5CTN82ekySku7qiZ2XzhezlspvabZfJJTwlD1/TMjb9fKW6o2E7ljF61nV
LZxgZrSm62jdJSFeMj7S9RIYQhm8TCja5MYh5/lskTdHLj8FV45a8sN3JbA78C2g
M66ZOJJb7cu9XRWKH+vlTz1CRlDFYGPSsrYg242V848XJo4TaMGasBkbNFLxg2KL
unuP9b0boGdHDn1BtgOVVwjCVv3Abfy8MjvJJvB9JkeO3BjfEGoskvEpD0wO6kLT
kyHuUlO7id3cnbVs/QjLvnLz5+00ST7RBunNu83vYfhpfaiTDFybdkgekCCdm0wW
m/POxbqoDlPkxgqbTBLnxvwnLMx0OMCRZhp9utCWIk+wm7PSbnl9BUZdwQB/Gn/C
YweGV0zXBgV6tUSm9l6lUT3kI1sVYPNUCYiXxfiVO6dDZm9wEXIkWvtb9FPd470n
yA0vCPICv+aG7CKJERphj36r/8+eUewFphVUoDLrxlRVcHvTWPNmyAfp0JZfXgfw
pOWU7svLky2DlZlMSxNFWKf3yIZCsLhIbZZ0FxcthO12ubyYivee/LJXuwed9jfm
Dp/yiFuMa/5QE4kAdAX1EdnkAzSGvqDbvfdRVwoHDwdPENhP4EhvkrPllfhfLLZp
NrooSLmYvUJozSWJ/DV+Kn++eLaySo0Q/Pm1wrwNdpL2US0Zc9Fz74EoIC2IDXf/
XHLTM3OXFcZzmlYcR082WdA9BrfTHUAy+Lkh8hEqNB0AUKfTpJN1E2uznzri2nXY
Vq5PRULPFKzxUINKhCVMASkqtPxsiFQtZ1LX8CEmHKbwYfmuTJxbbM9YXo7pETHa
Il6bfCY5xM/BB4ulr/kz5e15Fk3/nHVTNmbrQi/19GssoW0X+FRd3rFiADmlAAS0
5eWZ0lhgS3v0KKKO8bUGXD3q63YojtYD9Z9+bhNJqoFd4fBz1MzqZ1g+X+nvSDdj
4nOyCGJCPq+yiS47w8oDXVGYaBNX6M8HNw3G1XI32q/pzYAWrHF/0KJEDPr3JVsO
I8TKtYQyWhklU7R/wQpT8PVwiPLaHe7p9sDt9avY7Okn3a2eNPycyWcuuJkcCvIG
SJT1O3EdI3Vj/krMi2tEfBo3u7reWUyVaCoVEF5hb47ibzP9zoIYxJz104/3+5gE
wMkRjL0SGfVVnnPlqFA47VZZFOjOGYkMbZfko/uH2l/VpdN2Au8O1UMIBxhg5pDx
Qa6Zuqjw2SzXGrCX9vMjzUiqqX+IyCXB44sgvnwk2QffdUkJTn2iJaSV6uhto5ib
fo+M5q4VbU2wXjSL4xy5EQrif7cYO7W48MBjN++9tY/dQ9xqTo6Y0hal4sFie65K
qhkShPATdyEYUkbAoObEwAByvzjxxPa72aLqTwxG1MDh1eIUsxICYLn9ShHu7N/P
1uBjGYGR93sP8Y9k/pW0d42sf3dIfsUxN1xKg0uQek3QldJd84Z6cuKsmKlq50gq
Fm/RH/2ewLD+5otBYg4Pt/heQZizR4CbwCkfol6BtP/N8zwdOkoDd5d9l0lDEISX
DHFqAw9ksq3eGEBmekQ4o7P18kq6a3ZLGLYZlLaeTkO/TLDbbXhFfZR9mCPBodIP
8WoIogWl9cUkeSFhaBCWwVasMUaFcSZ2jjtjNjaDrzQ/uyNOOEv/T8UgUt09NNmv
j4PPQy518X9WN8nNVwrnpdj68F+CgkHLeNL9Mvl4WWFy5cm++aFTsyTre4ZDjQNi
YRsoTUBCwFw2Y4DVOdzg/K3ZJjb009lPi9esuue5PB/LGPkAtouYYeUuKqdMXsyu
W9hnKfg6KybvxJnvlmeNhPg5hzfXWveR6USAqrxvyqEueKU7nAST+51wUBU74pQb
iCQ7y5PeaEIYAuR+ARlqXCO1CFiXiuyrGYQl2x6mlaML2FhtEUltwnvGyTP9Vhgs
UlIfgvMf5d55F9yxMw4RPcJ0RT4hJnQpAcXB3ZyisH9isKbLIxYU2FeoTjJ3wbU0
31+FkZJ0hgBatmQRNNadcsf96ledT3xD2rvA+DzoDV0K6uvfDAIYIC+zRKehxjeq
LmpwAKDWmflCuVr1GuBO1KrMlGP+jX4DRlt+eAPOACey8YkSMmyeQczl0VERGtbA
J/MgLrq4Exgj/AHYy4T3x03XnfFbZiT9vKBVDL9V3BQ+UqG2J5M33nnCiuG5Bu67
ZC5QSPp03spMfCy77kU6L7TmJsxYMxi6fcAhhXkMBEVnBnFy872hxzkW0Rcpvyl8
cvM9twja7QnKwnghj85ES++xY5ORub0HS8PEPd38zPnoYEUCqhKDPjb9QYKvLN8F
0nZnSHoVjVAjzsdIxiotKXRb9AL6D9hi6ZGFykd1hiQwltPi9UtnUJUgelflAffY
RtzAFl27eQT0Wd2cV3nk4nvkFXhTCFyY3xhC65MdaUl3SRG3mNyFj+Y08AoRLVZv
6i+Tf14vWt2QxmzH6N4tuE3WNBvSIHQU3xXxLR0Y1wWng0WyrK09fD4oZCUXs86/
T8jPTHHxT2dJnIMSTw93AVICjxk2lrYwZFo5lQwxhnDqzngT1zQfYaogit3K1PGK
ug7kuGO+/qZUasLIFFvmrsPWWrGj2DDUWylkEZLt+c37P0WhGoaxrq3gQvmZY9Ag
1uf4HnBheHw3YehdCkIxSOoBW1qNLAoccEXqIHzDcbPxJW6Cu68QolIddDJsxXET
WBK6LyzDESp/MXzMJdOxfsNpMThjbnEOFjOQfPVHupmwvsd7HB93cklBBNnau6SG
MbJkD1XLs0mbqeY98wV6atC4hkHKwKZtBREJB/xaNJTiy3hgUfsmFEDwGTUCY+qp
bFXYjFgqB8GMpuCrzBlAL+UJxF0Iu//Gd2fkDnA+29Po5ko7pX5Yom/GkLUaIJva
qQe6UEVSCI5lvTpcJpmk9qT3kJTTPa/jwTH6U6ft2p3R/N+6HVgv9vA+qDqez6dg
TcMcxE8C33saNOVHBIdEbeXKCiODpggRD7LY9AxJFfK1P6m1jv/7NKlymdnaw6xQ
8VowOYu+jDRfghNypXiXhc+1nz5poy5VDv/lTPjbe61mZCxR8uzNK4VW4rdqGZjB
5vk9r99CVcM/l0JExyl9zsrdfYyELOeY+FVCTAPcHNsPuQ4rYoulbBV+uGzTqD40
lkBBVo5bs6B74RsC3DfL8Ah4k+Pb6IsOllhIX/wPNIILxBg7T+CiqGoE8+6tOibx
G98P2FhE7suFjeOMLZ543NL3gc+Bpk8i6M8l1lQPnj8tL4Rm4GYyh9KwYCJMf/Qz
cg9tsdxgs2hU+sszliR5X/sulAFVvVHyrh2N0KZCgRdXnliim8kAQNh/Jw6SPZCg
8qLx/8yR8yZOoJCGcMpqEICN/RdCQkjqvlQpUuRy4EhDpBP0RwvFd7lkRrL+CmcU
0FzgfTdrvX3qQ1Yxd1ogDwz0OcgESkUnH3//EnkFFNoOeL+8YFpGdKcOovrwrUxn
MNlq3TnBIgoqnvlH67UhSfpQjfVtEfPAgKE4mflp22OZndHnK757UMrwJbdzdp2R
M/+vU2R+a6TAi1TWdRE0byxa/wcsIQYC6365fW6w3Q9QOZkoLCeRGttYuOYnNEsv
R8n2XAcDhsa4uSk5lMitGQy0D9M31KIwX9UqneY9BmCXl+bBqF99mGaEm7pBZ5fX
1EHzVHbCfm9zYOsSBCpi3NYcYL4KsKWkPDmxe+NGcKGPMF3uQ5Tus2Eax9CD4wnL
OFSy2kv5RxiL4Mm6+SbmBBIdsCGiOl2giq80f0xddpkG3m1wXnRw68cNX85ID8Kx
vdxMjuRgi/C09HHI3Wtlkj1lJPqKkV4Sg8MRmLyvPKsNE+AhH5RfA9IiFeleQu8k
jlo3kP72j+U9iCnv82k1LAjsW3DsZrysW/DtUTiFHJECmG3070X8sqtA43djYxTC
D6Xr5VU7Hoy5hiTv31UBaatpIGoBR83s/fr6o8HxCZN9tWFCz1ErdQqB9MSLBvaf
25PHPmwc7nLWL3xJ7uch91PnpRwtyHEEjXoLOBjIzfTPlDFlpgi0Zxz3tb8mBR2c
BdpaBIIL19E1U3OvNYqa7Tbv2f+FSkOssPE4PPH9NyPcrgs6pMCtKlzZtBnExD5v
wxwCpFVi1rui8da6iTyA21GslapCPLH1zMpC51Eg8YV3nbwUI5S0FjNmMfmLAK/D
dJlZKRqnUJOnzRKe2c7YSs6e0lreEPbgE8WeVrXN1ksq1VMN7jKorF5ksrExYP1k
b8Fh1HdYvvDEm8mtAR7PJh8IN2ZnJhbvbncy0WwQjW8prxmNMdB0LJibFdxGoXSZ
O/dgK5y2CC7MtRZBoA1J84CfSFuJmqAngf7cGariTQUIlzWeuO+l8ll66F7tKw7s
UY8NHMHYJqJQVVfheZ6uxq/bNXUvenEEKuQfs1/0PZuDqTwCEkhQjZYPSsxr1uBI
U/q0z2n3vH3jrEm2ANHf3omkr1QhvXRRolQwyJInz/tbF2Kc1NTKvE5gulB0z95C
Dmt6sHzxmoXADYYGwFNSjg2OwW/Q3HcxnGIu3YWov70tMl1LKrb3zaRy9lomLmNt
2Y8KojZf6QnzohWTW7urH1FA4fsQ70bfN7QFBawsBgraDRt0r/ALjebNOVc7bAzl
aCf4demPj7CDaAOKxdxzS3FWm5YOOgzM7yP9EgqDgGwfFYLqg+Dow4X5Wn72FciL
aSDdh/JyIbaGIUd248lk/biL6Jz6oDfJJ85OyckmCD5qEACx4g0rBPcVOSXaLGSw
4UOtJewDToQzvRvchasDqXRKAbxnsSMnOAIZ4UxNS+r61RkmnHc2iiEBkRhEtlTM
W5Xo55eVa8FwSGd8f7DoV3+70cI4UT9mSEm2v85vtJeNoNJAl+qiJk7Mm36/3jmZ
aJToLqRfhfLsI/2HFjtDbF4pVEUusLj+E2sS7iAFXzCv3cAFnX6dnGmfcdts/t5G
8J+qRNM8Vc9v/wdPX5w2ZP/MLnAtsPHdtsurEJmnEMGCJcAR34J6s/v2tPfbvdox
CTDD0NicpIf2PsiE9VdC58VdOrmR5bytvcNxebus1NqBOdtF+yI3UFCWGw98FzZC
LDH6kNzcJbERuTQoBw8PsuDcdGGe3A7o7oUO75/OFxKuhdI9YeD/9URFfUH+U48b
Gbgg+VViL1Cyv7kWa/kJ6zkekD599ss2r5fb6YfniSTb92F3cYBX1v8gOwQAdE8a
g26Tgvnl61mkvdyLqENI4+dZixevYeG8Gut3BQG5Gg8P/P2/JIaz4P7oe18gDslD
+9BZu4FaejBpIZ7eUyjkD4t4hqxspDs9qEtJ5pfTUa852ZDPR6mxdiMJaVCcroWF
nvGbLHmG1DFdowa1xpgWrzLrlIr4h6iJIcawfBnwi3XpdpBmuAg+pnw3zveHQcEu
351/kS9b8IpdY8fJ60+2IqltLgzOwaDKa4bkdC8+VcgEaIa8Xal64YAdofhZaFZz
juc5/Ks2BfqogGCS5X5GxR/Aq3JrbUoMZQQ2ZhV21cRnpuDlTmTxF8uxF/e5t8Dv
5Qb/LyknZ+JFl9JTv8VBpVbUWnrKqNEb1gooIJBTTAtqvchjOlmnIRuuMATC1Xm2
yVtaoN06IY/7AXmBZgwK8qajlvaGpfCkhlMqVhvG0I2VGvzu3eniCdd0YoWXjmo2
ZWGaSZIVPaJzS+y23jQDrgp4UmY1Aa6lNL1xfBffgzN9P0LKiv+olSfHmlGtIFRD
IjRqui6i5m10rHF/MQbSAiG/o1nnrki5IqnPJYvsdP7MGTZ7GcNyUqGFmT+3vf9X
ML/Z9gdqiU2jRk8JtaO0LVHMoZATNiTkpcLywaoSWkQEv9evwDs20O6K9tnmOu3K
/+VQKJvVMsZ9PDxVJ05gwGwGb5pEoQU9A6YenqWOMhcZCFtNkj3ACGjkOJS/m377
a5xo1m1gZGSbyCl1oUrvdhJKTL5ANKO4chWvdJIH6VG/BbjpVgk5k/nGmy8vldR3
KFNRKB0LnTb/lx01bzeOvJ578LVKY4RU5ES0g/aw2JHjCFReHijpA1nqfzrIuzCq
1lBb6EET35wOuCpu6b4FTDDxf9xkuZJirdwpCgsAxnWtBypSFm8lftt1mJkbxDlQ
E2qAsiYN3jHC5ReSKAoN71LDCvKVw7WbjXKMIvQYV5xpP7F7W19knMCw+i3vcqpy
pG4WzKTSnkB41aOjXom9Akv7C3cv3ccYaLj9wjcvNibqJEX+f2o69KQ4qdahzT4j
AKKD5y0oFLIDjAHnLyqXiA/qhcduvDDEgaGzUcUgoPwTWUpGfxfgX/Sa+IzgEnob
46QInuyvnfFzWRmOYYoGYZjcT9AGH7/kPZ1Cw8cLZNehojkXdieL5ErMhijkhwBR
jSiipi4tdqxl8VWmFsHLl0/PtLdzVKzK0AyPk7cIMkQJHDr/aFyYePCWgTKgji3L
Fscbsnj/XUaefNXGY6evpRea4houFaPfwYdt89Gj+4OgO8xJe7U2aZgkGA5nhrh5
KP9r65HpF4I8QDg8aCzgE/VuxjAmrtKen4w6JfgojR6/dz8muce9IzS2W4wfehU6
OUwYHYjHLHTIYfQjTozt/V6IEu3u7cb/Egm4Cf9YCrP4GoIbYZOKsi7ntFbqjuLv
byxVfk5DFPFpvnZ9yNsDueJL2KGxMJCgNXKeqi/JqM3nH/iG9dABlTxIKQAWNEdl
1ZiJx3sUU1OdJ1zLdx+ahggmAPzgmt4AYs5Q9/EpJdiGtJMHYYXOvMv+dhOih9mR
fLvt8wYhub6LzMim4OTtaXL4Tpp8i2wAkjrT2kqxrFay7C/k8W8jb2NB3VcV47Vf
CgKp44/Wp2hE4rRx0UIe6LbcMQl2yjfq5tbEM0n5PIzK503nWveptXuNgGSJBsvq
K6zWt89zvelvcmC2a6wlGuwYcikwyRqyccnLxPk0Moc1+oltzkOlrTO2RdhowRDQ
QjlWeYTnWq/e+/vD+nJILvMhLlNUhNfEnZ/Ljnq3Tm3UP2FyhB9Skjszwu9ng+tG
v19U5hU9i8MKUx6yQFT+19nyD6VlWu9Pfr47WuLZpwDgxoBz4mzkJJCW9/18bauc
zBLbEk2ZXQ8BF5e7IIQrK+4pcdDIIIGR8aXsYl+qAGsLJOTjZAYbcjVj9uwyUuEe
jk7P3hr2eAfCrsPlU5iR51b+7bhTsxwKU7EzgOmZGQpGAmow15KUJRfOLnOFsaMJ
osVWXrL94mmI2Hp6kBcgrkjw5e16OLiFu+qACPjdISaaxRkEfJsrGT6dYbg4iOMx
ybRLxTUhUD5uy6zLZt7u5yA09/rgHwmgXc4/l3UbANN4DPaWNxh6fFXl9xJIEpCq
ci7QUpk9uRoGxNpBGA06rHdf0/YprB6VfBcrC2zeZ/jr1u63EMXhi9BqsM9cqCU5
jJemN++9YSArcGBN5DZbu/mmfy6lN1dYjIsyVdkia1DyOa3B7qUA4el9AQpCFVMa
xMCyTXn51Zu87X3tC2ReRjOVJSI1RfGnZPCBtgk/kEUqWk6ZfneQMyGDzJ1Ez4Pv
AjFvqVLVwsBYjI2fzvYRzsKx2lZCo27XeIwalzQST12hBF/4cJreqWOBE9W3h8Af
2ADUT03DMsA1Vfd6b3e3lN+yy/g2h2Lq7uZmmjPnff7A1lJJb88hOcOIQ8NmsUE2
xxrYeAYLqE42GM22kx5eil8jc3LVljnBJival/AN4i0Lem/JCjoDJktuJH/MaJSn
EhQGyCaUJCE/USx6Sw6SiC74SBDjrZyS3yDBCW7XarcPW1UqFeDCwvw4XZm6nHlO
VsZTiPsONFBTqP8JHBxycQiTgHcjv8tNZC1YL9he73TZQVOpodxoJAxxq5bemsdP
yc5NzsitAWzwvY2YmsDgPbRn864R30bamx5LbcCWJSWYDay7Dq7fycgiRNs38nnS
5ifLCISGK5TBSGX86cjVLiba2i/ybhDT7QUL8rSIs469pgjcctpEBJsvGn17+FBJ
qlfuaAae6QtquEeowquEMFNW44hHysUQWJQHAcp1/ZVLJacpvb5yQzMihvbGukQV
CvJRwOmQS5cVG8YBQUiOcPJBA8ruhi8HYnnVcc6KBOEJiq8s51TXTjOidoi0OUV3
VGtX3ek10RKhVxXrQe5BhF9NM3v8SM07xuV4HifU5iDJHsR6O608SsTiTbkk5q8G
9sCvr1XJrJ3NyB9sq1ywiYvqcTxEj0tdHFJimzZfUWmD+pwwIlK0M0s/scIajic2
qcC+9iVxfTPkuQwGV8W2uuAnlrDx8djhTx+nYcqOXvXEDGaW/LY1w3jikUcopJjg
njLUQxEIOGFAAE5nd0wPdiIFvVJ4J0BuLxWFsb3oyMcyC1rf7yqQMArk6sF1+DQ0
b2jq+DZn3hugSqXSzbufJJBHgEDIa3kJd9sgorOzQU677DmjaWoKsiZ/K0EI/aVh
CQHBlIj/twX37FdKbDccfk7b8NyPjIbaR6jmLSang3H9tLgvwoXGopjC8YHoZNeG
os9i5UNZG8Q8rUNbES1z79ugO1ISAidzmBYV07mj6Czu3mm143UFGGvQKP52fG2M
DiP3kfqYInavfqhQYuJeID+J/J4/wjCScEHfCYPEHyErYS1kCsiJlObGAhc7K5It
C6hINNTz/tYGjv9tU65MTYY//AypZOJd08dhQ7TJmTPaUBRqd+DqzvD0+t/jHFtn
Azw5HhWdScSetQ0gCZXin+kK30F7w4KhePme+bfW24r8wJQNrCp840nTb4iqoOSB
J3umP2aVRbCq6wUzXGD4Ldk2xRIDuG8LomE9DFYCd7iX2O2ST+eEgPr/4AEILQvp
DY5ixgous4TZfaI2KB0RAPgXJNEpUwz32GWyXO7mToVeKdbXkcNV4ZFgBaRHZig9
TPVD1zrWa1cK+az+G2QkK/98eMz0vcjyDr+gu+/2JhgpZF1pRbONnpyH/MQTr4UQ
Wg5EJe/PusO/Ey5UX4m9+T62MTtWA/D9A3kbQGIPM61UIAA8PEKP7It603qxD9wG
TWMYdUt5awvsVoYii0Pz079SdRVj/2hG4PCm1OihBggdlc3CC9jFl8Pz/5VoHm9q
4N7t4WkGrxWGkHIpuTtRqNdjFZfk0/bg17Skb7vqPUpX8yjoiyilGQQzJkd+izhk
Qul8AQt/2XvMut7mgNbriqvBIJ2UYdAMr2OJFNp+5G+gGUYv22gsSwbz4TrD/q4u
ZNiFxEXMAUabYEURekMeMwlR2JlX65jOGxc9oxz1TC4rA2hcBi9Trr7SnD3UgQ7d
ZPYb87ULty3yDYDVouLRw1VlU8YRq6GOOPseXugLI5xxmjZLXsbXeS9PBcbWPcos
kdwMLr83JOGubIa3wLtiBxpQY+J14hHe+UxyFhlOYnBebltgItvyR3H9pKJv233n
oKeAGUJ4bIEiPEL7dq/a/xL24bll5MUhqk2bN3zLu5WGUKuotDUjAnxYkRNO0IX/
X0xQWAGR5EekQETw2V4hg/D4tasZ7E7/MgBamQRaCxP0BrZEA1K4ejH/HF0y6Yzv
0L6+V8caVVnEuRbJtbea61abm1zbP7jvzxHEy2x/xgGNrc8r4UxwZCTF4/GjiEug
ACyL5e8VQrlai0TZlb7AwEpeUwTZqvBiuSLVnXEsz5GvVksMhSnNB/DB4fT3Z1uN
V4FTpfIni7dW6Qu8gxShu+7WWKcnxnyaR8xM26BtOK/r+gj46se25EoH98pec1Jx
lkE8AvGhlpSrTvGkFZUeLEZuI15Nr7T07Y0LBNKqT0h/2mkSHvWjq5YmoePAEpDl
iBHxGUUTopVHx+zCyX1rZh4iDOvmBTAVyDnX16rPOx4QHCwL+ICq6Hhdt1m/M9yA
X5Amll5gQydwJKgFCUujSO6iPTM2GI3RLWg1ubxSUe7NyZxmjhKV3dks3HLVrLQZ
4qCa05CKnxDS5O4zHEC8gduiTvySit0mbMLZM1+SgfCtDrKL/LTN/zyZmH89TwvU
Nw6JnHx+EdkCuWBGvpCHt8gDkRPB16yp0wxLksfDdXrhNyIZgzYvhiyqOPbzLVrH
P0gr+bof00DIhylp9ZLSmK7tTknZONs2XQ/WkBO8697jDvzQaaG9QxaHHCgHxDHL
czWHLvnMWHlCidGMH04+tfQgUjW4Sz4gv0lz9fSBctubzn47XRDbk4WRyXgIH9nh
ScoYZPD1+iIWwKfpM7zru/Hk9yzj05IC2ktsRRXX0kwEYvGAfxlHoNJWRaYiEDy1
040ArKBBsRReozoQCrzR8mDCEmEaNvZ+uGDRB9XWnz56CgAzjOmjSLauhXGgpZZ8
HHe7hCiiU5zgCuE1qL0xY2AhRHQf7vTDOVzmu9fCerd29Jv5Mewce6Axl+zOANKB
WhIh/x5/w0HjRzuZEXohJhEtF4nE252tCQs8mc6xkQTNYrfrd8ifZ4XQSpCV306E
MQHGQL3pIaJ+5yJ3UmsiOXaRL8pP4OrElinUlR3DLttteH9sXv68MhvfhFZIY3GI
xJd2neWbzqmKsolPlPOxMDBxolfBJTQtjd3or25Yw0Gt/RN7BBILezq1usZrwj8E
QCvw+cFcTXPql28VccDE2KdOiglkpHqFg7AZTHd0zMTXArPFC/DJD3A7uiZ1mcgJ
T6oKAMQq9M3N1lLnulN+OlS95u89M2EMlPaSvm2y8vMPf3VPYvQznkN3hF7NFd73
tkf3GL3PVgc57iYKz27lHmfUlhe/MDrqTMg02vZb6hI7IrxooBoKJZwOyPHE1tA0
HPpRLjihIn/3K9gi8TxeycXqxOmOIqVU7udRxJG4PohxlFGn1CTvW8Y6GHh3wCt0
h/Uyoec58Inx/1oS/tK+8Lr6NPiSHJFUGDNhgtaMcOEFsrsDqgWoXXFv9wutd0mz
UMLdHg9x//TRiHfRCt49KTyRwumRFzcBoNSYdS8fipJ1ki/4gdRWIC9u5rijSJhP
aMG2wy3JXMnpPJmKt9QPg4X/G6RukDroeT+Z8oBYuvHG9ehSTf1x1JSLDS05elEE
l+JGCUO9CVcAmweh42RLRf0ecpFCsJGkM0uLAs6RtLdvzKyg7VRXW/f2rnkBDmvs
sgjFwKmdLqZwAT4WG9Z457PDZW384mJ6qWQfx4TXdFveDQTmvU+mgTGbWMB/sNJ5
dZsPl89oZRaHZ/4NlzmUt8/kuR+p1171qSgKZ03ihUqRqKdiSx4QSZ8bLBRys4Ea
Wg3M1C/djPliC/KKXjUDIhkzZW8mnUTWVq6BMriMFb/snyb3Yw8fPj068Dk9qF3U
PoJanUfoylRn2ts5rXDWrofW7puzbw1Qe4N/KpI+CRCphDDiV1r1u841UjYqRCKB
abT0CDVylSXR8sRgrcYeW6imRw7uTvw/+vIIxo5A82+HsB/ggENXNI2csTrRSJhg
rTb1H1MSmLyiPbezQ9S49q2a3YGrLuvFRHsJxteK6M9dI3+l0CghpAsw12XMFgRM
zAnolWPa2snCf0UGKYWH8UiRfit8hRBgLQe/a8mKJlfLP0j5tmBKr/Y9T6Zj41FW
YcxWTvf14swz9bpSf15CCFrcLQ9XQirydMaOxNWUTG0TP+jfDR+kFM4rWt+T40o4
BJv8wJH+4GITn2eoPBd9sFYE4xeP1LWaVbxce/3ccIpA2FK+8ygBFYkKp91vIJWX
ug52t866q87jkpfzgZtCW2/OrKH9ao5C+hR/0XnmIRcrH8SX+iqUbUuYRL/DV/2f
bhX5Fa9Xjgq1RcWtNAlMawWgNOrZ3z2l2TsIGirgLuuoL3+ES2DgNGm9zbNAYVgR
a/YBtHrnXPS+zrd0BsBeko4XaANCIBwwJRckOjnZ5SFehRkZLt0ej5Ghkyvlp9uL
us0YxVr7Xuj/+mxbTISOpnmee5U9CApbreuEcRSJRZ2VVvlYpvNHub6JXfj6Lnen
LF1etcgPpa0dIZrDiz/gTPk9cBUKL9wOueciqzxOYabfCTBb6YANB3bWyTKv7kHO
j0mDOOEGVZ7mXKML99WRRaBkKSu9LjVSh+8iRZDIItj/JCjfNFMNJSZNliffFU8J
iXJWL0uaJYEC4UbAaFzuvlRmQQOueIcw6ceoKX5z07cuc8TZuoU0AnCXssH3t+W9
FpCXrJJ2B7aaivQjKBmNHATajtyMyEYxGys6ioyLvlevVLBO+ZYeqWjow6z47jQZ
G2efhVKv/XvyC/vb4NcW0+HkOnWNrrJGJdmYGZ2yA+8TX6G+ajoaes5DIfMke3Vl
DwV/Kfj8X1a+6Rv0eLYLJI/nPgL7RXYW7Ok7Bj8nlqS2TWgE8vzEEGldZ5i0b6lR
p+gDsPZipFXMMSdPcKYtUM4/7O4pZjap6wUqKv0Kr/v1ULug0xaDQAtcXmkvIFJX
KkXzKXoyqsqZTPvH1OHnVxRUEXnFfMTlJJ72cbUtZnbEARZXDrDpRI4X4riIiWpC
TnyoIr+czHMLRlWrog6C9zz+08WJg6Njwo9LbIGsqQrTC32cS5rjuCzX5SpOTPPi
UZTRY8IZ4ANCC2MgrvS3EvCOl5YuUwiheR49VsR34V5/LDe1KaEMtAt4K2wKvZWq
a5T1GLZiPo6EiSCxUEbu9DEUlfjxqS34+lpF5CvoRWakcpRxVO+6vhIG1OuhDBGX
RmfrPs87Scj7skBNDQqLGaMRwDwQQCGsrbSu0KqFbZXW25vZ7V48iEwe36yI1T2V
ESpE72xRjnHenJUJsKHU9NpGUWv8oES5g4yhMIbY9aNNfpX1ApCrOoW0VwnfEacq
x09L92HFSA2AFupSu22iYBTdFkRWpr8Bu0TuoDxCfs3GO7Mj4YmEJof7tr2w3Cvj
kn1XhiOzOGiDAx1OLMHcIvE22baVDGmZZs0zl5ohC4F5O7e9xFIkqHERroB3h0lE
5v0IxAHs86fC/QjlqzA2AdL747GB9z3s+oV3Wa0ru6GycSHGkG5LzZJHNT8G7YDi
ZihBmgZkgDrv5Z31ICjcVAzAATlc2p759DNMGOcO0mtvCf+O/hWbnXE6szxPf4JP
sA/+xdeWLJKPSaH//oQAzyVk2UDgmmKoRiohjpBnr5cu7oe3+tNMeQtpfxCRMidz
PCMcRacDATj2LmXMW0i4qPfJyDWvl90iKWrIxK+XwKBulsmKzdRjVDr3WslpOem0
FpCyMT63UGU6KUO1lm5NaZnlbr6Pxq39VoudO65FNKyWFqX0DE9z+BGKvG+WbQMV
PdThTnolGlWxD/J0Fz0JJwniSSbDbDaK5PQ/RnFxm3huNWXf8CmVgccJ7omwLwoE
L8e+n0w7KPFIlbGCE5c+ci/U3q4/IDI97MfDoItvrdki43LLgVR6ZO3h1BKyYJe+
AQKC2zQ9pBtb3GkJKYf06Tkkz662Q9ckMm/jT7Rg5gZOJUns7t3xycq6iWa9OXb1
xlLmzwh4KHQHtfFPXTJWkHCEVlVH8riC6mj6fxml0NP66yntqINmwU4BdMJBDl9C
NyXySabu/KE3TEj1NIfedWKNMT5czGDpDP/FyC9TI9M9xdoS805LXKVcsMgoUpTO
6yciHIfiy78BkxaMEGewZzknuL/cyUw99CovnohoThqRLeZqBU9GKd+FObKEoGTP
Let+TSHzhvxTHk7JmWaQ2ZS3myhBLo/sHL74uj2tlLJCu3/xwjRIZiJK0UV+PvsJ
fKuOhVro/qqd9ZA8l9FqjJr+p3JvDy54YKXv2DWF++3UZJl0PKzYCqwHwpjSXnTp
wbRwk9W3fc4D3iB/8d2tooKlWDwy4KGJ2J1fx0Vk0dxRJUPVO9FMUT8+soSqpfFW
cBLHHEeSHx2yXqhqsoy2APpDNuMiy3tsnhkJTGsSsQj3D7g6togwN15KHTk88KAg
wU5DkDtieXORajc17qrpjlEaiWjR7El7E4YX4g4KVWpvc7wTGnhwgdKDFKzZvAH0
NjDp2NNxWFbQPNAjsH0waIA1C9vVm/ZSXoQfzqTdD2nqM+4RKh2xPsl3uM9Vc2if
tjnWu9RAMz1aF235u4hli0eJ3Gto3bxq1m1UBMxWHUY0qQWWJ6jA7ghGKdt+NGtd
msCQNMQ+lK4m9BEO4eMnn8vlUq3FJaIKuL5Kt0A/dspvfX2dp/YzH/pI6RvSf3F0
RJoDWqqvVlJvZeZBnOBmiB7ZZv1hmg+wnPW0nbJqeR9+psiXjVRIf1Uh268wD5KC
sXMqPyoKoS6nuRNSZGNVgrrgDsimOuouIAUR/JZYSb0QBMkLhfyHOcWK28kYIj/e
MptH2i6tCxfov+R9cUbPFXVcS6nE0QJmu3zV1a11I5h+ytFlzCQ7mnUl3KghMOGV
ThBKTXmsmcSy6lnFkla5bspH236nVM1b00SQY5K6x2T2DFFO3iM7nZ/gECpqDONL
P4zw8fnAWZjSdbCoDiAOFqwutMtxptI6Ur5IZUUzuJmjJBxaCn0nI7CXUCBTaLGe
qyYgcVKMj1ox2uYTmMexEaouhgb8XrjSE/Nn9b2FhxtKStu5N8Hx9ttgEukWMlwt
Qx2mJE2LQfAoJzWfJFS1+/BUzmCV4XrdClvDCkw+y4SW0njxUjQrJSXkfS59DjYZ
2w57EZWJjdwG2c01wfqgZG3RVoPK3dTK2G4kLfLKFT1cP/hM+TqGD+IDCmUW2xH/
nve8LMkJqy2Nh9WJeh0ZnfnEcEJJuXNvvg4h7aM84D4VJUlcSiu8+LCdfRxgTp9f
3gCrxq61/apyAs2xvl7kwr482dbMw84BWnoYC8AZf15kVwPmaTwhKEdRMfsyflIC
8juGrzcF0ro4BSNmr86gRrmIhSm2preodXJ1Lcl+FsWaZ4LgOUkHtWq65bvhHqfN
qcmYgCY7dOihlXBNDYGxJXjbB9BSF3q19GiMb/d1AmesZ4ASDSQVsVQNZfqxXvqa
dsTpV6j79AxZSZWPBmWcYC0+o1mxKVvvwMozxe+PMTf829X4G4MrVcoamDziGM4Q
CJtf7cr+VvwC2m41Qv+gi3YKoIDmi+lwlyywtJf+1qcnr/qiPPHjAV0UQymvYnPZ
7eGJUz5PQSCXmII2aCEPcTTfk0ldDqwcWXHESVzXpyHEUiJpyzbpvZbpPVei7FJL
zmkXi+Axsp4e1tftl5Zlpe4EKt7Kl+a16opp6JUu0oGaNhMgs0SoFVQHlJ8qDayA
gHDYEUS6Oh24/lBNOXSjM9Aym7AyFjYA7SVQbbv4CVvOJCdqaBh48ruocFtXhbJU
oV8QDQG31cy95u7i7Rf5Uj/l3tFh9nYwIDOh4IQzmZXkaRW/zWq4ghIMM6uWfKt5
iJt1zoU73lxwV+yur6BqBtAhGpCE3uRQWLKSgN5W2Elel9eF+FrDfDlkvoEqGtNZ
4xheYVMkIOgYlZ678dn7iC5u+cpUPv3bRYhurTFnsJyVgO0deeI/rtpRG5eAQIka
F8mi46jqqWVwWoEd3Q+QC4PbXKTMW6pX0HP3x0OI6+cRgG5tdQ3tC3cZpRAp8hl7
wMvam6pj7b6UNX+I9duRkHcu/ZPXdgNPxIikFBNgkHKZHgmftVLrm9H5YF93cXYm
zNMn4fckuP+gFz6bPGDUzXny1VXVY8u/kqF+0LmRPBTC/praQJR3Exj1bpMUrhdC
zhyxPcNK341boj83SazPNHSThnz+UbrTlqPNBhknzzIwRsMYC4UgKxpFI1h4Q7q7
Vy61qhTwfKlD/yGvVkfKvDjiEpeLQ498QrJ+KJc6XNComJIA9viYoSVhiBuIiNgP
YsVFoy2iKe3+LcVl0I5cGLni/b2z7XnXjFbmnQtKEhPZWaK6rCrAsYr9EzIJGCxw
xPaUQgY7QdYWbvGd5h5afA8sIp22XjvUAeaE7YqtP65s9UTRqR/8oEpvXdHzOHnR
YgNKgroOgXXbDt9xcLiut+RCXyvB+krKEReCk7jLUWJ9Va1equkrgmp3J4CQN++J
OUoFjwGvIhd5pUjQZct0dPNT2qzJmv6GNMGOXHFqshNjA4L8yOEQ5Re/roVW9TyV
E3jblafiLx1RHD+EMlIA1XnsaxFFxr+MjMEmN62qhR/R3WL54NeWjMvPB+0I+68i
bnh/5kCh1k6g26OGMXSo8zFQa2MTDz9n9ZS/yVujb43lJNXOTxsMzPtttvjwBwxu
MUiBP6ooeQ1uArRaoVlQJNjlxsIOyfLQSvNfbftIVklu1pE2BabEekZ/cmBGqGVI
v22atHkNGieaJRfRC8BrL5jtdnrtM8McoQoZthaXhvkHZm+VnQ8KC17yeEuwlwFt
KvNPKBsQVehtx5GpyrE7Y628isBhvWkkXMy7IVZ7ZAnosBwdWnVxvD7Z18zQecUM
NVLh1v2budvshYPBTl3nuK/HrCVfkJ5MLgIhDMNJLyFOS575UxTbjopOuxdwyNDa
+iTFh1CDdcQPCmyqEnU9x2bOdUrYXKm2MiLdS6Ms+fPFGD+Qx2itQs6RTni+c1l+
WA7LGZDBtC0xA6U+X+PNClWXIBJdFOjcaN3d/9v1+geirxNgd7Y3wjSwu6rliC5G
QR0tVggAt41AGLLOHT2ymSiWtZtiWfF58GjvAHtvUDt9H7etEQi4mVW+QlyW1Dzd
PY3wuB907qrwKrIel+cKr4Gz4zgvJRZL+1vSs0StdeQd8U0gJVWUMx34fSynR6oO
IybPlyOIEutPf2LJYRm79xMqzPp2e0Vt+aEagStGIJEBoIbjYpx70BE5s17ywBxp
Ym/PfEhLbkQkVEZfA8IMpNxFZy9G97zHC6/AYENw31dBP4DXK7Ogbsyo4FRtWYLa
yab6zx2QuiAXxrf9/a20yKm4vWaH6P985H9iNWn87Oljik4Sb7fSVHUCet4k02qI
q9ebppUaGJUSuLbET1Hv9keltUHbLhVXeTdZIXY/LPXMZ6yyFUoH8hTFoINJbKMB
JtLZE7kEUkGegyecO9lueMB99CmpAs9qxzzHFcZMxRUPo6PQLtFm1ccO7b/rxMtw
8l1ggRtyt8Wwhb7dH6kbPLdH2589vPI/IUNZZgYzvPahwSo6GR2JZ6W05p7Eyp1g
9kdvJLCmnR3ySJpwzwPATEl7CD9dtyVU7FF3HnfN4P6RWCAgrEJ81C4H1ELWLzM1
4n8vePYgr5g1uo4/hqsTcRRAh2X8XNn+3iDcJymFJzKlkZOoLDv68mOuWQocD/mI
+nzdzS9W0GY2d7DNoFdVppWrU0cyCrxbaHG3CbLl+qlv2uRTw8ws+iVvt/mDp7XP
0G8WvcBHLWGmYi6vrI2poNyKcFi1RodAnH6gPfbqdyjEZA49NwzakamU9QLoAl0M
LlRDwr2tYfQPEsEXU4k0aYupQSTYufp+Sr3JXJZB+Stys9HFBDleqtZcKvsAk8AE
EHJsHATryavHNVYcuEfMy8i30qH+K/tjKSCiOmven7q86hw5/P3g4jHJJvMkdNsw
BKZoBiFMgaFrZLNNf2IdyPxXnfRarN6nfuzjepDSpfaDoMTGxTaLSbkIFsk8pR9r
cgdwvoC/imWZja19m50s0+d77mtdgaOboBgX3D2WIKsy83pEL0nCB3ZUWuL22S4d
4vXqOZ7LakYtZx+3icYo2DcCg8q8Kcr8kN4nkrA80NmQtmoO5r7HlwRvSGpJYkJK
3Ix4+G0IbzIs3oLEH6TIMx/2aG0AxSN9cz8BQljwcwKdDlZh6wph6XsTYYV8sppS
gOPbjVfPI4MQIoClp4OrNLt8CYdg8tIriF8IrjG7DNXLZVJSy6tVjwLeVonpDBaw
zX4kbJD2KN8D9+oQjsBtvLYJF3oUy1Ad5w61G8e7wlfAKqclnwPGEiqEAOP8jJJV
BFbr1NpEhFxziFvUf1qaqCu9PQvQEb1Y1DkY5SEyk2wXckIgZsdGWooOiKhNPcQJ
L3AzW5c5/WzH4mmDHLR3XBEvE9aGBmK1vzVx/wTsPaVTa4u4Sl+S9Vk2u9Q4aEr/
/vtlNbtrcUeyOPZRrUgf6LObuZke+HF3/uo3M2ozW/6M7KxnpV5NF5x04ZSk/DYy
SSigTedq6+C+8zDj2nkdlGimuiJDE9l+UTF+EmCOXbOM8x6+bUuSbe7DA/s8C814
AEihsQRjhtSbIt/gOsQL//g0vps5IUgHNxg9XMizTvsgBiOSSXFmB3o2Zbi7BLVd
ESzEZM3AP8juy1lTCdNFlhzrzuWXLRsVeKvNKSKP6fiDVw+CcbUPERqsoXvH4uN3
trWOeJihiYKpBh/PGZqNhkDkjj/yoIzCQrX/CGV8DBV/rDWwxBmOQfJcnfo9Xz7B
ME5qEMz7qtbXXGrLBEFW6jFU0dGvXaDN0VL0nhEKCVBeEJ6NIURXVx7iGeUuhsNE
U+63INAlkEyRyvqiavIBdZXps4ntU5yLWYJh4LnfV+nLQ4vPm4fdyZsw9afezeX5
O+GqJHZqhKoKX1+1+gYnkZbek+ElPFtoip416uV718eP4cxn6gi+/o+oFMbecRlZ
lqD6+SypZApaKP+uWowdKPXT/cYUjcB35ozT89eLrBCDtvaZPZwpDIgcHlHh73ci
jh6aGuY5eOL+1gp6xHlr21vRmxkt92LoQuVEg0j29r3TJHeXw5FCmiSAdPV5UbeP
dzAdK+4+hgM8e3QTMPHiYaYnEjJ6GVysSfgafn/Qq4aGc/cwkqxvZhOlhdO5dYfs
iPqnIf0ZI6xYrNBpX2jio4+aYH+EcfkjK7/V+GppzWodvGPabvNXstEncoqsHTW0
M+ifQ5vL5v/+O43p5ULUrklDYwok5Za3P8lnVd5xBbBS/des2eBpRpMDAC1lUh4A
N/FJ9hyU1bPKETyaRnrSJSduEbMBIv/Vy+AfgmGm06ehaWJoAXyOxDlW8YolfWmM
mQwi+MVjMmPthDtZCtiNHNRb1uXzr8gi/kWIm4r6Ked5jgqruRHHX3bLYNC92Ba9
1NjCa5krySyxUqMA8M3Dg60YJLAZC6ekaUDAhl2Q7rfPmlnrlfr70WWWNAeAsyE7
v/0CATHAVSdbi5Vtcofs+c8hxo4GccY6QL6qy2n2N7N6DLLmGOZWKif9Mo5glCS9
pN94NvlGmloVmd7Rcr4vUlN0IU1rX3OiZbCkQr3Xa46aKOpzqU6wbgslzh+n0u+Q
+FCa+b5Nx7tzCz0oYZEtlATj9uDJxToeREur/1as4VbFpQQBmw4FPa+Ab35TJTTX
DMcCRB1QjDTctJjL+sthosPbHUfU3omGaeC3cudQgERKhY1Q2sh/ytLpHEZq5bKd
AXDs50rGV8MQToZ7Sx/XLXHPiKDrgMqOg0r8Po3ZE1VWR0hWkJBixNz8xzhpaK4K
r+2md1VzTc0ibbm/b88dthke9/a8dq/jgi5rgpzkCeSmRIODtYgVZuGTB8pV0zFW
QlC5HEigjHhGMuHDMXA3zN20XSWzET8q9ewpJxYyQRE2iN/JpgxZHcaRC5YhWLDv
/tlALx3v6v78oK74xIg89UzyixOljBc3ihGX+YefZvBHPdkvlVLPu9b1szWIQ2y/
1Bg/2uTYTsv7xqeiVMLqzRdP6EGWH9tDebOwvMbT++S42snVrJ/RKIGCCRHJmHSG
j/LTaU4DkGXd/VHk5WnqABGDhYWqueOjQYIKilFsu/MeiKt9s9K1Y32mlx2VSNT2
h5rvqbNrAi05EKhCRkpZ5sXV5AUhp9itRxVue53WLid7HO75OjBaFn1i6/k4Pgqz
LYV6ZHki+kO3hiPiWFctzeVScHqvDYHo+Tvxl6jqPZ+Naal5WdrXSesp/aJykq5i
uNWQ9bvlxoX+AHmeIsUQ7ib59au18pBy6cFCEaOewW4O0DrdqXbxmbJheIXoXAdm
iIte6oz+TBGTX/gapBy+DpGHvar+HXKUnUm66sDrPZ2BkEFewRcKGnQC0MWQClPA
5lW0rcQp8LZmRbgJBzlUmfLhN7mrWe8o5IZXSIbQ8C1PQnbceUxI2tvd9eXKLd+R
k01FywIBk8Y7Dx1DLaeTDvUed/jcynw3e1iKTqszysywx2MT3Muce/pGVlx4uOIa
FbEkeQdNe2tyxrwnr5yR2Tk9OZg+VdcQ8kWkmp6JcTaV6N0C7HPwgXS+pWF5NNvm
i4IS4OD8JjjsJm0Tle6wfIp3eQHJTxdjhsEgIAaeM7V5rDTfCMsglXN2hEyWofNg
IpqMmckV86Nc5qTVC8aR4Dy7JGXdjMr1A6baFUiZQ2zchMLLD9FR8mb6Lm93PxvF
7iuB8eMIN27jUPWQY1QSyS6wv3z9hbuNOkCP8jS5r87EMTKcwwwz9EJ8aX3Pal+i
rTn/LmmkHd5aXBXMEhd2Mue6wLLOP0ysuLslbQ34FtD+cJuXivJjZ5fYmT0kKrNS
iZwJu1rjhwPRI2pauqAV7UcTZui/vbKyYWSBLamHF3LSY/KMVhfLv2eLAYQhIBml
iAmIWaNOOBDWJviG/RNGRRn5CZNAOQx9+QokEOY5fUJ4HnInZAeL8nuEu7Nli8QI
15ll6UjDmuth00kAcVdm0NanNgCbv6LSITcIAmS9NTFKtPW8KrL4lIRzfVwrHgfU
26iqrNK/YAotQywx7IGffL7VuYTLHCYp8oukZxSlqXmRSuaNtUngHFGWCNlfnhPt
dHAFjn6T0gQSBlFyIPlxfgpb6iMElc9mLj0xUNGSaFfRioJIIti95LeRTMtebnj4
vhIXhnXENlx5N52BN5iq++gNP7EXAJoLyxy7GLUydciI2Hza/zze0OWPWJe0enof
JUp9FqBOltHjkMCN/01X6NB2NYasd5ZUuLJDNWcILlZnV1fihwtgGw/t3MpPWeuB
XSbuQAt6gRemMzCbVistI5hd0FOZIUq3nN2d6ecl4keABS2mKLsx0ppdb4J5ckyp
m7PMWhEW46c/jy52PRJ6bHLNPy5TaLGO8LTVHFs9L8E48pQ5W6JJiliKpIya0ZNn
g9+w3PyjKciBk87r5Cop8cpWw0cdb0MG75Ko0/9mzicx1mN/rb6BfxYpoA1zb5JJ
XGlKvpcxcxzwOkdsD5IeVlZnyMUrBSd41gCCbvUs1LeV9oQHZqlibRh2V7DCTpeh
LCGL5Lby5f90MyIGHpfxos2ZR/B0rMKIjpBLLHn7xVe4lB8wqCOT2NozW3jYR42u
cBiAHT2b2koxisqplRZnZLNlWWAFdRTVon4O9v8lj7QXfrDUxbS2CXcJpvj5IV+T
dpJHxHdRi9vTu9hwqhmOjX5UuKEn9B7hLneRrskRQJSpQcUJrUkivVgLTDqZf0Vl
XAI7WPx2arIQ9trUGFpF15wfVe3Dm44ax0x3RkK+EBIDrsPtFOxNq9Vf/d1pjZ87
XW91Hgaiq0VEkLVPt0+n2GnEgIWEK7LLoiOzo0MSO1zf0tcc8CjnfG0t5osRh6/N
HU7+CQM02P/cm5z0gqZSMOonThgI4C+Szr7pcGJnDrB/snmTREeyU8r45Tcwsfw9
89u0MZLjQCDj7zTOXv2ZTFbki+LMIdDUireHHe19aacdxlnVCqylVDKPUxL5HGuD
GERW79eMirQSnPn8jSI7WQw8hooOaAjzRFup1lz6gn/WQ4a3RcZCnOpkAWP+tVpH
J/yuyDPfz4K9RL65TbvsUP47W/4TQozXE14bR2fmchAeLXOTsolSu82gXBM9YWWJ
Q0/hGeMylcV9eolDMIGqlHr8vLNm5JDvT6pc/Kpo+cuxdyWbjf2TeJ2WEDHp07Lg
MhQtPSXZa7l347VKBQrN8ArU6EW6KfTW9eknyvLSbardDQxPgmOymDSwKFXcQA59
MeLHGfbpx8bVv0PblMwS1qjLx25+YJ+eb+rpl979OVzmIuTlwL5cebSHdVfQA/H/
wpqsEyLH/tiNLbx6VPFFU62SKZoPaKby2jqR9zeEFCaJpJZZPXRDA4LxxGMnpL42
VC+SYA1LIKgw58UHGjzoBiLE5hb7fHOdphnKgna/MkUK1XGjtFaWR5RRHxqUlQDy
t7vZjOCGhqpBdszSbclYMovFpMJaWf4phLDlYCXPIdkXwhFOeYYRz5te1oWLkimw
GFMujPqS79Lppnd6wO9WZjOpCInbc21QjAlLXf3kerLQJjFvcQUEPjFklHaFTK/4
26q+ezjtRgzeSJCYCwSUxJtDA8qZUSivlcnhxs2YrZH6F5+/mAiA0PCOWa8aHm3o
ig5cOQ+7RDxWca+R2/zHLw47N+hOeUy6T5TFd26uE3tc63JfoFjvVcyodEGW0mcY
3lX8s5vh9o24E7wxdUBfvcSGvTPHtC6qyyu4ABzitVQFdfix4PUREXDltR+pvZ8k
KdPzToYYd+d6rtEcoLwJWRkk5qVIN1ELfPG3J1sqoXjnfESJ7FPHp1MHG8453gsD
K2Qw0JPSWvEG4GYpNLerfLGqht5WfTdMu7qqhKV6zF/bC1nqLtByFYp1cr+jEqCg
yvxpTrpogAoTXgz0E9OL/a17OwsRy3NXnPHvmQ5TKg8WqxaDume8+r2OBW93Op3N
JS8lU8kauAlELsGYAPHym0GEYgB8U0IyYFHkezWzfrPcDCiJFoIfuYkrrkWr4C0B
Z5futgVfaVZqzatD29r3fkDtU4ysTLX0jIcVjRvmrk9/mLbJZP+VjtFAjIQZfUTb
GoFd5vhupIFgJj4sgrK790PFhfDrDaV2d9f0a0nO7nAhFUG+W7WeNiaDOn/w+POE
W1ZnnzcYp5Q7bIGHp2J7oojmLP5YUCsgtqQPXN65zkSDtLsXzOqZ2/fKqUjllcKm
Pwr3htVZvoGyjeyxYdm4FhgbykL5Hv8wL5LMV2GxkhdiiW5Rj98wXNt6O8NEI2PO
T4KXk2HF3PYEGNva3cf2SNEiqjX/ohN77/Q4VBkOaBoTm8SAKXZ+xLrZ0FD3pN7I
H2PyZwossm6gVVcdt/3/fniEZbeO0ZBUF0MmTWe/DfmdFFyD4p33wjMpcVUjtjiO
cY43qjnfL79FkdQNfSGPpgRxqYJqlAghyia87hfha9Xj3O3fAFwJaVxtwqAq157I
7sriTzZpjfNuFLXj4Rua1SxL7NczY5uH7ZIU0Vtl7vAYMyny0TV+Eprc1I/qvwUW
oylMxeHUSkyJy+jPYFRYJRs4N125R7I6VaGKKLP1h54JqShDAFLmmMqU7X++88q/
6DQd9HyZQjS3PVK8Flb9b68MiNyTlKCDfUKRZH3lmOAxQx61nZxwG39M3f84fnxc
tD7AzDxZRA82aHM9yEw43b3WJwuJ2mcQDpzxBUbMTDaOVXTDaCWyrpd0tVzb9Ym5
OGYPPuThrc46mICp02LPuNPSU/FPSBlJ56/1rpQ37DBDYaiD4Ejs+lZPJHhDGsLh
gkoI3Zhr73vmfoJHd6rhJK2LTKqfUPgSZOfZ4ygWZBIRwr52Y+ZwKvTWLXPw2bU4
UaPJJOoCZ5PFq1yzRpY9zt0wosR7beaTdzJioapoC3ZnpbigJfmnRVo4APaGWfTE
5hH6ZYqKgwWpzMr81k7vwTc4j+addQPIb+B5Z1fsCmkvQ45INqDDc21nak/fyhcq
jYEwajXOOZP72A4Jzjv+b3vep9e1CZhos6Lp4/AXdMZgXrTcxgbdHFHHcDr0F1oK
JACm8N/+j2LrCje0XjV8Q+F+4jfd0O9DqWo7gZ5ioLaznM7N+ZXdxMzPhFF7fMT7
ZPwY9X8D68R97qxsrv26daqGdEhYhbLPbtpN9IrOCEvb3W9lohhS0intRsms+AJE
BA0NFX2qn0JFVZf5Y0GeOscifcSHj3bPxzm3JNelURFxp1iyOZOZIKiis1S03xj3
F1tjA06Q3lwgfP9D6oKJXf1844gMw7XZlThW3/+wCnOf1uNujANh+UYKCLe4FYzr
/1a83X7FrmEQc3VEhqOhh6a9ew56E5Mn5ZsfZQ0k2k+BmpH4KsprOAZTf0XtCdfv
ome0Is9nH8+RdxWUlsX3NxMGqpf11WHhhpHK+wDjxoRrfPLHJB3JLeoqoBtm+SvW
sBGHfdbA5gnBd4DUEa6WbYcjzR6dQ92LlrDXNdvJ4G+ku9mwFehoxQ0YmXmX7SVA
SXI9ioL5wtlzuSzfMgL4zGNt2NUvWkpxKucePuhEsHRIJBuD4N8sdLbxmHjtJusN
i6fV5OWQ7Fna+U3lOhOkJ0dQbAuGmTTZko1UV316d/Ge8Oposh4drZY/9rm9/NRM
WhAlmV9GTQveio+oxcYs3mvIRGYILcr0Tadw/GjJlLCt0T50LOnkDZFovwW45P8l
GadQYtFY/J3clZtTanG0T4r/vtypqc2ohvezBBU0acX1Mw3oza0DtyNyknrNZx87
zUeWMypmSwLvoVaZHY7NKyMMND1y28q9euMDU6b7QanTyJMB66uK7TcE2bJd9xrM
i9F48lNLlyPKMTY1WlJiTXQHHk77pHtig6+Bm05iHF44Ki+aAEU6ebvJu6vSrkDA
4rx1iNEnQhUlYUH4DZGghKdGChefeVJEVoLL6o6wYLkR6OJau1k9qtOFDYLJ5Vll
MMUeCCjiN3pXdWVWvPpDtDdW7UOlfTKX4GZj6TEzpvj+u8OgsxkdIl73IRlI/5jQ
mAKzBvuJJ3YHcag80D7393T6jGhzjzhFyIUNij3GH0s4wZ0moXfVJdsm9usX8uwe
QC6VDHAXEh+adkkIslm2GITVUsOVpWeqeR0APIFrirLDaQdyZAMNMDwKa+vxsNj0
3fyAgIVAPzv6TWfI4j4pLwfBQ8ajHsuz1m1fDeiY3NvzRpw+E4g00GL7LAgzENnE
uAZ4LsLGBhC7rS8hGEIBTsE0iFLzGXk8KRJcz74I8jOLrplnIk/1//VELRGiloP0
6et3osNjjd6nd1NEQyWesO0exM/Za9TsM4hDii+V3yeM59DnlAKdFLmvl5LxWkc9
S9unIHPAIJFDUGNEbnLLSXLfkgKs9OeZnL/SIgWrIbuUwcb+o9s00yrxZ4zm2Ocu
twf2LqXKrTkrkkpASzM4o9UBwl+kJZ2RhQe5fS7rILla4qNG79HQosEqWo5RjN9O
MoeA3Zhka6icDouiwOhUkBwr9MdL4XeGbTrSh8BGAE7NDrNeMyUYW1z/NR1wQRHn
qyI/EG9gRokR0GZE+ufqGyCZXOlzbAU2PPm4VLa6b7D9rTNJ2GDIY7aFCHhdUJZT
io4tAliDHqS9/yBMdmZucR17vEPqhYx9UYk2aggoDromA/ylYNQAYMIEHTROR1By
haVCVYBfURiUXguKMiGNhTQJ44lmpqJ2msROlzb+72RJqfPFKmaWb1YPCZJimsQA
qD+1C205bBspAqqT5YFPE5GPdoja/os9AjRnk+FJXjnAoFL2iHVEy5Nab4oAXKGY
slIhvoXC8USYSNrToDG6Jb1TLjOPqXyUKA6Fa9k9ri9BWLA6kV9O5S05/5vZ9YdD
jMSRkIFYLA1kmBHbuv3p4k8mNhvz691eGPkRctAj3+Hd5pWe4Gj+ldUAo/xHGHJi
+MUUGHS5kpzc6aHTQ6/53HtlAI6SfHtlf9O4roQBrHw7QMTmEzBZIhxhHnNdDszD
FAxggeZQBudB2fIQu/A6/gmcJVsD3UzvIbO45XJjKkejxfbTcGsA8gUTtQL8vuXs
eI2pUC4AYSdC4FKoV7q62xa+ec2SrFCsmYvrfe7Qp8wsui/UUPv9q4GaVzt0eTFy
asx/RzPhRr6MdGJepyPVEe7oIe23RepD/YIHKOjiS19wCfo/AsSptF2gORt2uu6L
oagzzz5Lpr73ZDpmyaUkCEbLwVMXVdtf1mslNvB33j5YXLRCSorLkh5A5bXjYnTi
by7z4M2sjR9+/nUR+q0QjkM+pyhNd8tgUV2G0lPvrTTIz94hDtZNAJXQtXuWgPPG
S3R2MMtd4O3TuEJ8w7NGYpkzK9ftY0NEE0BEa1SyCBDa+sXoQVahp4WyVdK4u84P
cWGP1mQKajn6F4pYH+pQQ/dLhsTiAfJQOnaq6Uo9H3/JgMksReUep5PGm4PzcV15
CrhhCRQxaX6sQKsBnd+yG5hCe9FXjA5hIYCGSI9delBHy2tkic41+tRTKlHDnW7N
I/orSve0rLgzFZJvd5vFVoMw838VfDmGjh4kYrJ1I++2enN2BL2TIZJWngx4vUfe
h4IeHVItueIpxR66pmrnGu/FAW+IjJqzkhUCHiXgeXkvbH4NAVjQ/DTZJr6md3W6
8YEN25LJ84LycqvVeC2fihcO7Uq2SkuHIeOGT0CI74rc1JszdWB2T+Vr3gyfvX3F
CA/1cENiOOKEqZKyY+LbmJu3SdW6ynPlB2lXKksMDRI7CGRgjKkeEh+A8//1KhRw
HS+Z9K1jQLlcSaj7pb4excRIY4aNhXoqWQeABKZ+HgYWEk95vaK15af3fLPulYAU
mJbDTNTjPwonOAe28PcKrCWM54GQIR7UpKra0nF0Lii5COqw3xRxWInyLCR13chD
N6OV6Duwovh5+Q3J0hctsPTTvsnT6Is2yQjAX0XthSUTMGzAINHtydb5aeyJYcK+
3ywhEhf6wLGe5SYclcG3XeK8ZfhTO++CBew0knNxIOvqpeqva8kP/gTCRj/cKiyz
87rlqgSQFaJvuAXab4S2rTOaQCADTQRPlVqtwfwzTD6PcdAVT0cKQLk7ThtuinYY
AVF5/Ju4xtB/98BRCGf5C40BQITxOJIFD8CGtUIhyIjzNZl6b+CcB4cC+s4mt5ej
eIR9ia98y8TlkfJv7rPMA+JoR02tbYgtc3nRhp6wQ4KuArjIiHknSKSjw/yZTD7N
9s6DhQo89y6dTv4dETT5c13A0c7Q6ymTOEOU7HAWOjHagtpB3q1uq3oZMVQdKn4F
0nv63tEt5ohCIpOc3BeRJCllslmwtS8q/E0y0dEb2Lw/siPMW7V+tSXuFvoSEL1K
tnHjNTSvJAjkQi3Isb5ctoaG4lRaHwf9vuv9N8PwDC4t/caJH/V6CnyS+Gb1gOsR
8wAbeU+a9uOjnQsPIL7xR1WOOX8C5irrx29PVPw8b4UEekT0eIj1N0kAr+kRIxtR
atmzgPEJOUxtAJdfg/9xKgmuYGrbi/00HBBEtnWbX4Y0a+mEnyW61in17UHCHin7
HisrZkHstd10m5v4X7BpRdEVpXYhJemKI1iAKW0JEIhzxAjn5lEyI5qq6hD66cju
y8k6oJUVFpMYwXfncN7YmUGuQmgBulTlnkFqB4P3jjF5be1mGCN/TepODFZgvq9I
mCs9nELDzbvzUC0yLHEnRkTUAWZfVxcwd1kPjUZBJtF6LDxymd0tL2Bc35b0fx/7
ku+5D83iji1EIKwCqfVp2BNURbDZvRBEk/8R44kfOj0/ICTLiWgKOpnE9SX+xhpa
BPcqayJQgWt6p27w3B/f8BND1HESS2KzUog+hWPo3PVC5eaSzU9ntmqiGg84xenH
Qh0Aq24FErG8u08c6dPbLy7ZWVx7vVQi4hE+n8Sy9KDLxoT6DYH37tUK2KCQr3UI
T89yOmP/hfZV4CGLtlsvYptP19OHTav56RxK2N85UxJeKDDYyMEOW2n80PUNlo/X
wNVw8FdhC+tPohGm5umHS7kEKGuV+88sOjCIskrL9emhx1gEn7yWBLfISkbpAbeU
I6ONus62Ko5iPIA8+4NgIxF1n7ySgAb6UFHiIdkJ0NAb2JSdassZNnS2SWFxvmmA
EqXIC24INKT6Wcw0ZtKkR+7Re7/C0VNlYjs20jIQK4kAniGuibK9AD1B/mJdH0du
8u+peJbaihNshz+V8tn+1ilVIyxmjGr7hUUPpX3pHp31iNSaHdi/FYJJtZUU49KM
9C96EumCaBE+KmtD5l555Z8UJXVHM7gZOg30MWAvoL+7Bl4Nu5JHez6raEJphZm4
Zv6iPWQOax3HaPyqHQ37Etr6V6rjhWMzXHjcUw9jxuY7qaZigGevhO+u3Rj8Gv/X
8Hb32p7fwIVY3AWBcUfj+seP4fQt2ey8Vu5Svw5rLvLoH8/isVRovh4/FYN8bbB7
Y+CMMnYmNXMq2rbPmPKBsFAyArlF8eyOFoWYlGPNWkiFchd9t/L7AcNJc7/dshiy
zuyk4s85zVyaMj+gKv+yNa6Oy25hIXwbNj1RiSlu9AZUCYqlHORHnaXjBCbdEV4B
G/g/VSJDnXIhNqWmKuXaUQrzoGajaJzKof59+rGLccWmMFrgsBi47CDJPMw2fFoE
9AkqTSx8iogNajhe3GJ+97InPNzktrrO1gsRVrk2Sa6aEMKUJoJHwBIWsjd7PAZ8
FJ5KiIVatUWCLxwSLWNFosQ5os361VCQ6vbK6OtSdJ/TdWzmLzWZIzyo+RM0ZFmk
z4P0dfGWo+a6YWZZyf9BNSJG9euakhS434R8ezXfcV9SA0Fa8jDDK8yI1R1/6lZV
b1HKSqWu6MQqH4HF/zdb0jsU6/leqFKtP1+gfag9rM2SkebDUmnGToMOMAeQR6H5
UL/uyZ/BcIOekck4kwUt9JGEdFj/iBslCE6rKtYQrYhwV9Mf6L8QNOrW7YXlDP4R
rx1Fauc/U8C7gUpBocR/o3/zhwrI1CnF2J6n4B3wdTErOnNus77ueabmVWrqKLiw
0pccfQHVtAxyVIOc90hsj1d5g5iaydDMI4cSLweg/NrspFV5RFsBfc4WIm7ybEDp
lgKj9IoC8aDdTEb4K4xrp+cLyvn6SH/BV0fNyfb/gk45Peu+plknZciE3CH8OeQT
vJsyRd7yerR0/Jco+/4RlD2MkJ/682EloaCBa8u/qODHdmoD5aZEArvldMeZQ7gT
MeoGLdE58FWABHOCCd7MXSKmsw6fsLltjtnztY1fOmCNWRRJKvXwTqVDw5ZmSb2k
ysXVFyJmiRgcuzRtVsvAsMIyN+5RJgHar3RPY1Zepn/yYei997zi9BY/bXbLlRar
X/4HaDLE1WnqL7K6GinTT/z70rKg9JqD0Dai3fWV+sV9v7aGgReVWo1E8vQv3nEg
5OJqOdjkL3Sk10SaK7fwxZT/TC5mCd/qZNLXLJQ0PvIRbJ4t9ciBxi3WU9nzmQ+1
uqEz8KdAEEUY1ij9HM7jQQJHSAfSDotDk0IAORWcQLQUUqZbMcy7MsVzOyX6ebzK
BqorgqL6i29HLDhlHBBCM6iI9Ev4RdYVbpMtVHr2OrjViYiib+bk3hWZSOBQUNUR
ZFmJ9fNTwenkM2Pn4Didzhjt6dMv165k/RWt85gyfmxZnZWTlWbLuerJDoehyETH
8i74jd8BUynFiQ1Af2LsDwH0ZQrFJn9hcmo4roJJc4QGQ/09GFPgsm3HRGrvxKhF
rsI1B44+xHkFWXflzD/KJYC0f0SMCdpXu7Q77m9qsaO3gByR6niDTMpQ3AGQTzNu
OR0Gsgu65xkqVnu0ctEe0aYyYDrbbfp8Me1lmnG0P+1jkWuH3UqZ1n8qvHwdCkiF
8jgoqYlK9XapkmNtGrPhdcTkWmjbABS6Teeq165jyMVkKg/rff9PPc/O7aGsev/7
kFeadFWepLMuRLjrGqCGwATz4sVJDj1m8pTc1T0RDH/lk0dDajLO8gJeIngVLG1Y
YoYBMX3Ekd8F0IXjICwtYO5aq5E0eji8GlGxE+zJOnhbW9YQRcchWNvnG/OlrUyt
HreBFBr0UZEo5DRCE0jd2UoiUn7EkOM1BG/M2zArw9ZYq7VSWI1bY2UPETc7OWzB
FY+OoR2wPskApktVSnSr9YQgrpaVVuyJU2bD0O2KuK75Kzi5vwo7DSqyjARt4Jwu
qeWwMI++cAnnplLh5KuqatnaASAQfFxIW/BvenhgC22jphbw3ND5V3zZJhQqoa7/
oPIA/DrkHGWYPWEfyDVypEtrKlJlEZilJS2zBw3SqlOfEslCMw4xQtqGUB0wfKn6
oU8dYJpA+ihoMMW0nM+wJB8WDBvz7xqo7VbgdGarf0YU2cPyJmUombHb/0JKntwR
OUAoW04RcM7SJSFLidU3UcMYjlryHJVXg2xal2+qQu0JFP4/UztCrxQPmJwtEhLq
TTLWCvXLjYKxYx6zPzlMUFHuqmnGGSy7Em3Au7WoQG3qLHSF8XKrZLfAUEZ48aMN
fLbai6PFoM4W3sQLZi8Aq7as5+TZ7qGXyinRHRmTM61cYgVUBVXR00qz/ygAogDr
DTiuW4/XN8Sc/9LFLp8h+MwxyRHSJMhKx61OwWkJqi/rfI/wl4/BQsunlBFTDNY0
TC+gA47egfctODIwehqQiFQjm+IgvUjBONo8hNXkbCTFmtTMdSFLICZvaE9mK//w
BoD7EVLTJ8RvBFZ7vpZu2DKuPiadQ+n9njvGxBtACiMjm/2jVJNnOJHvvHhKuxy9
KYa5jYkxccCJqEAb7yfll3mnuEj9WMG7+bbGUPHaf3KS1EWYa1pC3vIi68wrKd4F
75A7ab5UiwXkAXU4c3Z5ODWSSItm/JRZUHc729yqFBzzr8zRZSruAQ1QcV6dfmSW
MwkrYZSc2HonjHapxnMgDXm4hRrtXP0qwbG+2q/yew/E4vv7zVKb/ci9q2GgqCwO
nk6V3hhzxIfDaMkAt0dmXK+SaCz9VaUbEBPkA5XEZ4y0GoJ9kJkKPbFZbYWGMmWm
hmsc02j7D0P5vC6I7eCWcK5IjH1gEszAwyPNiSSwS6FneQ0uSSY+KnaRne1YhAGi
5cn/pH7k//Af8rag+CSzJcbt8WhxFoJSAhmXOzEV6t5g9GiL8A5PYUc/kQ9VP/uS
6noQX+zH5UZQVW6hFvOqgk3QSNMU1euT9o0OlLNGhl1HigQ+W4IVE8rEQxYdfTeV
k4c6n4LY88wg5nGL+0LvLy6kN9YeUbQ+2OgXxeiEab1P0RiY0R67L8VBuey4Kzfw
A5NtbuslCSNsPhw2FXP/ltXWyCemyuAjg+Q3+GdPKK0HBaZDXDmebDcLZG79UUMQ
aLIasNdAcQaEqVUM0QdGV3ifHWcL9HbYfjTYKJqwdtvMCo6E0SxOi60YDpqAnp6O
lXUWfuWfBrNLtU1mu+Q4Gta2qkG74x+/36ha/Q/TPrFkB4NNrVzIJSwF5Zerzb04
YLIm/Y7jHO0EpMc2L7hbcy7zyoV4468L145wpH+IZxYqwPuiW61lc2lvAY5tVoQA
XoYwqCg232d6VCY2xQszKFPDrjrCQ8rRMgAsunrJ8ki8P7CYIuGT0VRucRYE0Rle
6Z5yNdyc/uEzssDc4HQzVmrFbsWDaYGkS9PNqhs0AuQDNCiysXHvd8OF7ydMktYO
QPnm7ZX8KUjzPwSbsNyu7aDqfEp3ynR20IOXDbfMe2DizQfgQ9yjYVEUeOw26d/f
g/kXf0pzUSFLXCG7U6+loO7W3HOA0KyytpwR5IZ17FH9IWsl13t1kjmyoapqEJWm
EtAnTAn9+fCa0MizORo6qqevyBIykpF+NEcN4ZKD/HHd52ZJit1DqSvdddj9JWgZ
BhxltsQLx9khKX2QuKl55mWadol8PcdTc5AqUt4nDpFE16uO9pX6vv9EP/XrLk/o
X6LicMqnF0V9HUen8OAKwnjXlarbxPjHkUiT9L/BgNeHa9oc+d55j/8MK3xNCGw7
oeoGmblj8wa4QKGoo4MRP7aykqUtd68NtrE4TCemRSgbJ7PFddGpfRY/LQYxD0aI
N7r9ihH62Mhh5fFtAtO4aHbcbB3c81sJl68NqBM9wfDVo2brUY+UMqY5rgZW0q4r
u4B3/PLxvNOz9yaK49x4f2vLN/saVotYPUtJE+1lw6HOkGrNnhGo7uhKyALHnw2v
gcGJrv6kxFYkGGMgNyOjli6JUh5oqGAGXb5cI41TR9mR67qqMm+CtTIceQ5YMyKF
ALSdU2PE5uLdrs8Z+D5Z3ddKKLzYob9uHrN8AOfCh5j8cKoo0re1UI5NHH8xlLZl
Je4+HYMPfRmWm40JsQ47BWVhgsUhEhJ89p+xMlYo27A65EILY8wEdgxqL8tA0H9h
kWqJprN4IdFMwxMOwvMPgpkJ4725H2bsl37GbdNTX1Bc8Z3H7Jh0zN4HYItlJ42b
IMt/ZjJVO5lDR9pjh6l7Dy50WlgTkVvv0rnDF3FCJLZIthavOXp9/N5N+GZFZO+d
QwtHpPoJofzxC0+lxch2v424KpVHi0PgWYoGjVeKvZZtJB4wOPndnoyfCyyXzXxU
WfbnZpyCU7kbrzHVX+WwTEv4bMjCYOtON1iZc7zyUBCCLxssIXcMzYBweByVqLfy
fDRwM4U9e6v13iA1yKFO1jn2ADALTjkUsdsgsxes3gTLilHmK1o8sStFsJMoZTPj
7IUueDUCltKjHXFq+ynmPjQZJXpm6FVMhI9ZVszCmgOB127rwDoRS/HI7mdzckCm
Y3BO5qyepKPZzDJyDR8h8cXtB/xBggbbOecnsJ2oEnxas8MEPVCsLT/d/YBzUEvo
IkgsWA3w1FLGQxcdEIUJxssKwn2VyrBeMMa+wWVC0YvpyVpNEQOnt1d8gp25+JnJ
VhA+RYPgyQI121+assQ6k/JsWSuoaQR94LICLiSR1xOXZuGX6lMguMs0H7LHoAZT
ysuedwxswNiacTnQygufDICFTkh4pv3r+3FkCKWL75SxXg2K4f0iQ/qsb/W7jdJs
K6uJDGT54zruei/72JOOgA==
`protect END_PROTECTED
