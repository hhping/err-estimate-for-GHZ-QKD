`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GB8P6RHFPuffLnatD+a94TO9wQJRt/tub1rqOXhivyGzW5rkiJEr+/f7jQicduIO
SyMDWMY8l2GHr6hvWsfucMzfTyWMpdPQRTTPWK/dBnju9qCo3jzmO+5QoC2YUHQa
+IzOB0R7ahI/TjDYDYwPDOQog0Uroih1TZ3WewVxUZXWP9zqd/XitsIm2gitSjci
SUZBsY4ezBgf9M1KPrfffUpq+XUMwibXBw9sfpZFo3WqkdEujTKRyQ0gKgDtbxrx
rqZtwTJv/htvf9Ah0TTrHRF19AUB4GACFKtjPMCGUxHlfXpW+jQ1d4m4D/v8zs9x
1QW3Ph3FhjM7VDwuOCnX3v7YLFvjGSEEtM40q6lH42Uiswv5WGpqXRlefmRYOX+k
qGryRy5v52VDjy9JcF+F7p3XHEIxyYdBBIE4seH/if7tQ5moNLLM5JmYjjUKXie4
n35KgQFLd20kitF365xj3Qt6gH98W91WIhYIW7uQzCsSRSGzR02ZKgez2iXSHnJN
5coNs22lV9pQKTmZhrIywtgjQUmjl0fCG82uOWipOkmgxRMfcIS3Jczr8+HXd3vh
1ENXMFHipZGtt4PDaT9V4ZyvMrqJZLBtrQzHePxal8bQo5VtICBtpYlrHQkX3jXh
Zx8oKpHXjsAUcqWSoJVH5p9CaPKVMA/PuQvgtnmPa1iKB224In2PApux+1p9HOQA
L0250iMzdig1TvXvfYxMW/YfLbOCh3fD1fj20ffkTAUvUfn88X80P3iZs/1zK87Q
m+mBfTK3kD3T6I2rAIeBiVlFhnX3Cyx8hj7MxvnQrLLfo5+1LYNNkhI24hh7cgkz
6vvhc/1zihvz5I1661woA5E1eDslfZRCZ+UaNav7bOxNtIQHyHhKn/8tPeMBYVvi
MHPrDDKc9yTDzPJjBXjv6/NXmMh34fgdZsbSdo2uDLZoUrJHqIPIDb4hyZW1UFCg
j6TxaNg22FLu4Tx0eMqVzAlfYgcfPPVlS1rIXf7S4ORKVB/P2E9KLEa8iWpk1u4z
gBhXzArRan+U++yLf0YJJBqzHTqaOxTLglkqh7nrWkjORk/d2rSI3yKqNSkKJhvu
aHEHN7gq9KbAsD/b988ncVELZ5nYSD0yD2gyfrou9vGitnN6ukMn5irnuOpdfwCd
1asIFkBAAg+6m6KcYZbATQss5CL8s5J3otMtNB9OR7MkKiaxdcM4XwA8NX6kftG4
+eutv2HJoPs3a7bDW9I+i4aBOO8I1i/G0ZWy4fMvgp5Yt6AXixQFDaoT6Fzi2g8J
uF+qCLrusxjryWvhQyIR8O1sdvP/YyQSjE3DV1MasZTrp8KnDsNSka3vfDD6xVzG
aTWPbSXLSeOZS007nPrYw6C6cztlSrQ+JKlPtOMT2dyL6U+FW+yaZ8cb3JLQYxOU
IyEn37LHhVcEmMijHjWtGZnOGojh42Cl7k9uHJAnoMNupVzn40zQV0bokg6Zh88S
wdQSf6xSvAb2XkW540dGaTO1aZN+HiI8XObigNe2XFlyK1eZpQPk48uS4Ghth0aC
YQa7v8uyfrzAKrBmdUvh3t/SapyQpK+VzZmSdIGPF7V4YTyeWrlKa4JJKQ73ocRC
RThbMbt43UT6ULna/7QNTWf0IBVJSFz3SOeil5Q3eIdZYh9qVzcUAx3Iaet21dmH
DuMVJMwY81t38/KbVXFUi6YJC6bZOp4syWtzxWZP2Ouqeq9ArDsQ5QjvfCm+QFXA
0bqxSjqDyaoGKhT2Kl+m71UpYUZyGUcN7xrRXS2gyF7gM5e/OFjCTEP2egY8+JMh
w+I/OPCLjlZmSRZCE50sABteoacSz/fBLvc4DP7IgnJYQQYlamKGBWrTp8Jbu9PA
a+uDQO7vuV5PM1ALTXQFV2n2EcFqTCDWI579NQsWzNJhVwJhCbhamNYMZ2xntxRj
YGI1z3u3v9bwsCMgcewsoOr12UVFrAx6vVMQM2jc8BDVEhnyOjAm/OoI3MNRArdi
/YctjfnUtzd48Bz/zj76GVXt/rZIQfSdoWv24XpZPtQK7o5rFA9GPgqYh1w7SCX6
6FcoV0u7mtH0/rGBohVNEMpNM4Mmzp776SU1s124pVTQJZcryRNi6TKZolEVNJc1
+DsUsb0PO8t9U362HTKYiRzaby/M0qrpuJT6jHwjdaH/FMQkn94TFc5FQt0RosCn
+3/98tL0TTwW+NPqrJ1xZwxx30bF6rGwKPxrQzeNFB4CBdYVqJrA42usY9EnDO8B
nk/QKmbnAtBD8l4X5SC6KbQ5DNNkl7Jr7E26p3H1SKkdgsqRYGiSltN1lVu0FW2V
nnfeRV/1o4aYy1wrVt+PnxMTf6u/FkaBLsAnBCZxtCKEO0Fe3AwL37Bw6vvrFxwd
dtgZiyOrsOAEMfyPjkCgZ12jkxNZIDP6KOTsibR4sZ2s73lRZlh5wfTKx9KPnk5Y
gF7GHBmhCc3CqXGH0KUr0/uhirloE1cgWLJOvThBBGLgeqfn6KsDIuCiAufXV82O
1ojLO5EoHWwnwSS/mLhzynVnZMLj6EFyIJjkGNsDvyeN77GsyInLAOfF2R+wSYg3
ZAHP4xuQscmMbeFHpyNXO1e88byWUvIi1kL3Rb7d6w3MwkcDF9d76U5TgXZ+LLn1
8PwhnUw3m0kskxZoyQoCjcsuBye1MritUFnKk1AgVy1FmU1+TNbqtfLq/Pbf6zqe
GM5t52B3oWbkHhhJkFPtFW2l+r4UCaCF2tjDTEidR84WK1e1y+MyjgZhSw7kf/Fv
H3PhSZjYHfptTQ3UASdfm/RXzx2LNnJlnG4MR6hAw3Rx2o1zwUkWhvfuzGwq12Sq
y4Wq26/8HGeR/Ep44IRa3JC3Bc8RCDpBfwlbpTLDP+qScJdEXQWXei0rnJ2CtKrV
edFDdTkCYIxUcgw6zZ212NwogdD3hqtfgtOMAY0AxZwREpq069d2JsNoKYYNKm1e
FDjUtng0EGS/xxV5XBX6fHkqo6TTP8fQBeF4jQ9a91psDtAn0AjCt4528wC6HBEz
tIec46ue7dSU+rYPmd29rB1Ypna0LytbF60CGdwx62taOmn8YWf2CpUMDDB7m4+a
Qi2izRBFb7zCjfjuNbdl82mh3GNm8iCCXknSIXzP8RXPUiS/8wLBBG2rB5qQKQX+
Cz/Xmov84MI4fTb+PU23WEKxXJqQXNg02vC3meBiVJMp0OWlfgkqtQyB+mcm9DYi
vcfHOWrRgcbv9n23AZE4xK1x/kqldYLmrWuNtXAfPlUcG96a3bgwsNuLBC7x/MUp
BXaIp0IjLd+xdiqYPb76mjEGfYceZFFJAfU6B3Hhl1S8XfDV//N7MhkagYXzpR5h
fPku9a1lwbRiMLHFwggDXoRdQlSQH9ZFP/Lzoqnf6zc=
`protect END_PROTECTED
