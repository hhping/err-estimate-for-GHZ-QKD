`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XQrcOB1EAbl13LpF1BVnkkGKCxB7rnjIO8sA64waignGO3+ydZv1iTzTbopAcL9Y
FFnnEkYDL3zwgN4LqM8j6XwSyMQxhXIRZvdG/wcp/d7rTb8natwngh3XvSpGtFxm
j2RY6y7HUA1IT5HX+qJweoVkvtP6QDbuhwx6XXiDgWbHR+RQnC0NjrH9kRAHh0h8
fhbF+mjX3LzgF+EZUMrnZQ8/TudewndBr7qfE6aipzFHidtcidS2HggewSdeRmlc
1sU7HqhHdTtFcJ7zzlFVqCu8O4SrKgmUmIMzlorTgrELnEG6G3krSxrHFlqIYedG
hC29RPTpsP8FcmYH/NH5Y/vcOiUdhDcF11h9WFw0EXcb2+ugIRAaxOYexWcg8tXx
c5txTZzR4GD9ci5NVyTwXOsNLH61fSjMUHjpjM8+GufvZxsU6rN6lMyfccylsWrx
MmBpqSOrDVRAK6MAQ68W9BKApl62DYYJtQjVlLCai06Agf/PzI/dKvLUMGn+w58P
A/lOvyp9AR6pM/GJXQ9ANtKHO+eRfB7TqE6GHq3VU8NhewRfOrUsGqOQA3DHO6Fj
4Nr1chkzE/MX9OpCL4x9oeAi82ajn6vYHW0NYGz0M/yh+GAqQ1bpZ18rhZw1BfJf
8T7NNdCfaTj6OXkZKTj8GjUuFBS2cgvChLqTXbAj3xo/Skye4k/eFHGEDu8zirvH
Z0l72sN0xxkrc5LCMvjIhx9XzBACfwd9k8C61KLg8Y0eSLKuQCetv63FsOiVVVfw
QOPEGWdx611rLUKWG4dgFfLwz7Y8iVFleLtNs4zBX9ILrk3MVe1bB5rKQhpGB9Wg
1giiezp6wlaTKfyZUCdvWOPxKV7hBunVYpKwrT0NTa1YPCqDQRNqARoK1Q90bUJX
YJpVAdvYdOz9r96oyFyTem3QK6sipx9V7OzPJgcFiHRSDNx0onAG80jwPAFlWR+A
bWPA54QiNhPkfxPat59Fmc4f+5yJpZjgzf8n1tMk6wb/ZFbkiPishPIdgqrbepDd
zf7XUCJscGvV+hrcl8dAQKEAmEWRdZGYt4c7yTv1Pya4B1rsqD4T8Csjdpb3qnvD
GzHMumNLzxRVWptfkR63czKIFlt+V5dWaapxO5myVuJem4fZ+50SmXAnGFVm1/bb
7kJ5uRfuVvUaMF3wbkHw8NzDyfZCjLVCARzmacsGU1ol6u5DHuRr6lazONr2QAlx
4100+fvryBBnTksJNsko36dyh6i536J3jJ8HKb+KJp0xKXjAzqMlKr6VSb6tq8ZJ
Osh2EggZ0leLY24wfjqGddy6/h4kRrC8vhZeM5i5nSLRZvrOwr1T2Jgax2JwT+NJ
208+Wvl+7zWdGnVaX4Ih6dtPw1tvtRESGQfSR4W2//q1/wGQsDlNDj1wOr170baJ
G8pMPbPgBm/JQApFIkvgF98bwlqHqCvcM4vxOGghtj2VLsemmwiKuCmlqCAsNlYI
RYk6XfRjES0BR4OO3lNdjufjkZ7USKeM7qCRzRnj712/kkjmi6BRVqndVJ15iQ+M
qag95Br0yK8CbwudBIdAuethYin7HO8qfvgsnjT4CPat9WiGozAOd9P+ShTVwiBW
R6oRi+a4oX141G8o1XhaQj8FoMbN4ZybElc1ecWcWMpPMEKa1ZPyhHzBr74Sa9fp
`protect END_PROTECTED
