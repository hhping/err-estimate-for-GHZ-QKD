`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xs5pggu0X9xouHdQmD9pjZg/6L4DlnLQ0bZwkTlGUpniUwZYI64UiXm2fEVo0p61
e5SyUdd/s1TiAxa7BOO9CGRZGfrIaTgh77pgc7osfl/Tv9daqTpyDrNp8J0HIFC7
CvdTyEr8wgxGBEc7e+9JdkjPUeWhQRk3Ix4RR8HBjpczNfdV+msDWvDV30J06v5E
exWlh2oUBjYHNG8HJTHb1Cp7E9q8otvgkjK4eUmqGO5z+u56kWyd/Bja8KqfbiEt
txXkIUKZOWupDbzjA3vrFrwwTx8v5vZOnQ+/EXM0+hqEaGAzDSYvllATmlY0ecys
VSMPu1De1JG+YEs4VnGntofbS7tTcTmpvGcmmR75u1HoV4UGFLt3nvUx+ui739Lm
FqWnyyF8s4dg25x2/GZzXimTRF4emhudhUfp3gM3eVCGZIvb3t3cI5kWoykIMFPO
Zd8cgHSmfsJ8XMHHNFUvK3nGXFWTAC0xfl84sd1nvjIMgxnf9K/O2ExZwfFPXMQS
6H84ZWg5bHpH9M8JqxPtZj/tCHC6/qb6tRH9oCo8G7FTbikC6HmQU22Eh2G5LT1+
j+kssfOVidXA8RBGizVBiNfbPE46Bal7qDZ3ausXkgiQwkGfRes0SwrJfLlZ+L0k
HV7SdLwHElq2YFUPjvIJB+ADHqMQhN8u09GXfrAu03gaZH5UXQJCEyZ/lseXxmEV
sQBw4LzzUMIVzykzKy2SsHdMRzcxFEI1hNKwN4HIq8I=
`protect END_PROTECTED
