`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8EnK49xTugPNlIoUHcVRISgVQkeUbUU1g3xcq0sUbgJIhMpwATu08g828QNj3+QB
KJSYn1EQKJppB42oTLeVa+bc/YmIU54pRuDt+OlD1uK72K7f2i+JUUh9FbMphoT1
SmFBc6YzX2D4Fb3b+hfv6bcAoWE7OEIB/Fp7vLVb7129ZNkGxZMQPFMzkS1dGEdG
Gkpl7aB2rfu3TMz0iQI8Q5BWldz+AKXJZmMn5xCwMHIh8tb59ML0n+47or3OBKtB
i6sVVH4vCVhM0dAqOtmsZ9f8vNO0QQ720WOk4NPJcm3vEd5KpzvNO2CM6Y//HGkJ
6ThkpTaOLTbNvBQCQIPkx1Tyeq1n6p1YicSkz4hAAcCVPLVr/eAng2NXG4h68o+7
hXQ8t6TvNefokV5g/x26pLZ5/64iV9bS7VcjyxIcwz9MZGi/iPYn9fVe81TFiOzV
k5IHZ1fVFL2bqBDeIkmzMtmnYlyyA2A/ePhKkobbgCMGHjbCWPE7HZblSpU4nVz7
v1JmwJVl9q2Vb1I00AsPF4UkWnHnx1NWCG9/G/3EKAcUu+H1ctyi3LKhYIeKCYex
KKC2WIXekJrtWjgunoCDPFG3LSQeXKlT1ehGL1SJzyq00MDNs1Sh1mTIVfQuSU9u
2BBpXYf4xaRRxhOVy8yz/U6MlZ2Aq2wR1pW8QxfUflgN7sErtViVORQNL/IVLFXD
557xP32GZFw17L4/KxJG+Mx+dPAkWseXoWy9o5+ZdXxop2qFZBVV78g/Be1NVAev
OzI5xh5uOpQQkm6KkVweAAFJ/EHO0OsgrPh82BYaI9DBGqlF+wYUn4zy1UDE6b+B
vDEtuAtds0gLlR7IcNezBB+qxsuuiJnpQFrGSMUCLl0H0YG2v7FqMS069aJMweOK
khq7ZmPsjwb8bYim+PjPmL6QDRmJ/8Ol8RVmeGHiD9XHaO3A3CqdAVoLihaalQT0
2P18poF0ODfGelPdhYMomnFZ9jN3RNC2MoRKvgBHXZe51FxjU5TZ1X9D0kNgDsum
mZUzSH9D7Kclhq4H+wvzLmPSYrkGTCcj6OIVqXYxHvgxB4n6cuUSSHUkzUjOrlEe
v64QPYsxPavjMNWslvHa7SBs3k8KuzmbJ99+obGasWYnH5BpSrUqPlcP7dD2PrYg
YbEa0/0hQO2g/CW3LPeCjPS6Qj3PfSmKBx9eI4SX8B5agf/OuRA9p49ScPXxxeKA
EfTvDnXScKafZUgsPOMxbM3foutP+Wlr0Eksj6alpLKHoTQ3nqhNB3crPTqcG2vA
zlXhq6egJ1g98Rralb5+2mMMY1cARfa9eHNU6aeRXPHRRHlKW0fq9g82a67Jb7sU
Z+5M33rxOXh3OrX4uHBunnBYOW6ku4wqfG22wfhyXZT5q1ekjJoRF6hmoXnRz1bW
En8gh8Hjv1jjOT6OCw7vJrYdDkJfQcF4CxYJTRe4m8E/CZFNQuiyiXbVL/eP34f4
oSxzZu3b08A4f4i4jUQeRAwRlusBU3ylCsQlpWgB7vSGaaxZ/ngTJuyCw2uZzo/B
xh66wxRX24vu2hpH9CSoElqe/SnBHMtSA9oq/VGx/B94RhYo/EjX1/qqygRTNS57
jIXMDQvZLizQV+ZbifJr6QdArfs9UtqWlDpsUThIOUCn7XnjqtfA/oPU6c7w7gI1
wv/SF77HGdb/fUfhadDffyMiyRbGHLTUTLv2MAvajZpEXE7hS5W/3b2CfDjv055e
yYlP0qzIH5rY/2BtvSX+FTOXB9ZVVI8qHZXIAXnER5xKBCoMGQxuPkWfjrGItzNb
i3QKGWr1FbtlK0R+RCxQ2omkvs5NX+QXT05PQb4gxePNkO7huMP7w/4O1nu4EjX0
yFH4skAGAwijkApSggyhKuzitfMghNhHYtWtlrib2ndzQvapa8RO2K0W8pUTY95e
poD9Kkql3z63bVS+Kr7NHlV4pfhDrJEv3nELy3cYmT2BeMEitFn2Ub1vgXxOyfC3
Bryr2FwTlvDNba1wi+ZMJZwUHSbpsfVNC594uBTBeO2NcCBEHI+hOiStND+p9G2b
0zPPqxUHhmJXjEOklmgluuMHaMdqoMg11W6hO/ulBpi5SELLKSHwwqzhJwKhevYj
ElFo8JTWmoutsORwqJMUIAi6Z8KhaHHtnNTES5ZHmrXuPFVM1hqq4KjvsurOpiss
Xf6zi8WDujibB95H4yZdoWzGoqoXYC4jOPzVLKRLtYgGh3UffWqz+8GfN2a8KQzI
vkU48ekXhFSLDsIjauwmiHH9rLC+HX42psBudsxj9xazSPwJl3+Cbx33cBvHNePB
1dyGdZo5TvScjfgpHan8aNq7AXj82kJum4MvbvDGQdnd3nvLcAb/VgxecUwAybf4
mkoFip98nNrGkGqb2s5YpZSgZzU0s4sRpYxUpRI5ycG4gTYi7iNTjabbWCzSyQ0e
hWkPHVGhOPTsMfMIjr87pu8wbIr3T8BnWT0wi1oRSN2OgpKnWt+7NmQIV4aoYcVp
nmpyBp8x1yqx9QWK8Kw+WY3QieQhLFjCp5/jf6MmUqWXL/EXSC2QzL8QQnFuwy80
Y4Snb8kU7t0r0ivQdqncoSKZxlJ0gHUz7T3fNCf0d8VDBp2HBakueJmgZ7nulH1w
uwL1HcRyt67HsPrh0YGaQiI02M5iJ1ZHX79Vdl2K1aCt0dhEW7JWiAc0nx7uf9Il
K+tm8mXyXLJRCLZqQ+gZe2WjsSbfiTInKEDfrx4IcAqBYnAvSdmp5nWjLnge/TaS
udUChVVAqPQjRQIaCtSgFoBuODBE1ylcqcDj65Se1vNeeqalBwriXxSEGbji71pR
HqrAtxbD0fS+vS9GD6Z/2Ey5m6haDRk1yTtD7Z+FHcyqLRfQakkc/Ky1vFoforpk
sF/mHZ5fcbPycl/Fm9HmctvVu+CAwDWB3Aqev1HO+NAU5xDWeBELUpDINbmdubxz
t/V46UDqxNjEStOlNX9bQvJxngeGQ5Y8XSyxOLdYDuOk+X1S7WkKA5rEAnz/dEzL
ygEP9525UZX6vX8XUL1ECVjB57KF3EFEp400in8EjWEh5l8PMGISORUTfEtc85il
+/8Ca88QHjMhUUCOHbgHaxiHKza6obKZd6lZI2wUkynFzParA2yXx/OgGTTic75F
1bl6tn3NmAknDBcRVJd5yCV+twtMXbfH4lkCZjYZuKgToMTfZluOVqVBDcwwxycX
3rZsw/dlS3sziyp4VfneFYe6EP5DYAjCCdGey1BW5JNNk943J1G2KZxJ+czboR8W
SIPE3QiQksNdJS95aJjjUmuGKf8grhO+AAE62p375mstb9U8FDUkoAoD33FUgQLY
InxpiN3Oa5ojIs1LA5IZmqQTyfcBppFO/JwSQD6AKF+Ta1BRhg0NGdz1JDKpVSFC
A/gYGJvXRXlXtpbMVXoy20PEe0kRgFItSU3Bc3lGjMly3cUuymkjoJbdjWmhulDx
mO/UV91rG9AtlHFrcFi49LsuCMaBAjEyMUxRMcnxau6QJcOpnvv6dO1lGEG7/U1p
OeoaybhzYD1VGTDw5EkhDV15t2/cjTG2pP93ibCVZ46GwbJlufVxX9YXDZCLVkEw
mRXNcEFkl/QgygqKr16ZwB4ylZ1uVq7RRNjAoRROV9LvzQzXN99FiCbstntISsTB
Ar1AkRXCSIBGAo/9uD+YjpefZ16NkQivzCZ9ErILdtCoXc465ZnAm1qotPQtGkvi
GF/RRyoqQctCMcjS+6OgykTZF7cfKmBoqI3QcUkFPFYGhG/4LbD7Kz6EFETKurwC
m3BgjZnwari8nBPCheJC+W1KSxus9nsyQ4bFBqLNdhIdc1XvqjM3QJejlcFDVcrm
BsXoG1pFR5HH7zzZby5thOzTzEwUiZgRVMsfpDp4Hki6Rf4Y8i97uLNqHHjRZqNU
AeTv7tvYcNQGbwvWbus9jxBgWhd0U02mpcIAwx+VDnr1Jwr4+XC+lt971w6L7Sho
A90wGcnzxU6HBM298y5Dm3mkMk1azdsNxQPHdjbIPtadTA1DHd2DZ+rIjhCUj+A8
KoAAjsb3cjBKNg8zcOSkBzAC2AZxN1WJUZBOOBhlbuBcvJ0i/5gC/0WzO9K2c2MU
5XibgBpu93kE8uYfJ7V2Q6kcAwaD2nSBERVyZoP1hs9uyD+VghY3FHsRxOReqFwq
GcSW/CB5qss2MYjaQ+QoLFMdZlis80EOkwaNb9XEkOpxYx4amtc+zTMfwKIVyNaZ
Dp8NXzHFx+lIPPONot6thFbq9AQ7dDf2iLUToI7UEpYZ66Fw2Th+ywzCno7Ua+9k
CzqaLA82dr5N1Mhdlj6H2C6P86sGiVH9gQOxpCKOavhygmFFpS3w44ta4F+CdTQm
3ej8lMr5HVQb1K5GWRTxTeSvrZ8LKLHHc87hf1ftS5jYXxIloTHv+kzqgc2xki5v
lH9knjuBIjDCjT8PWrMWs/6rp8HSNcz7XLzFcsTm1xMAUlGmgpbRmjmV/mWSqkAQ
x7mmcLHizSNX3FBrI1yn2r7uhgThzxP6TDLX+pF3PnfQI7xLtxQ5wRMlN7TKwylA
7BF1wEDGkefWCAeow1EzCLOh47ZIO6gY1M//MK/OLoa1P+sWcDamw1A6jbKthv6V
3S0gwQTN/wVoMIhbk/mOUOai+fC1FmRHV89nrxVJSZifFBX+707EYRj5TXaGcAlU
ZdJUbRWacEa67Kho763oINxzHF3VKOyWiK7fVGu5pM5IYsGi/7t/3p4Zk/AUc/Lw
0WG4zJZtp6JbMMiazT/60XwL7LkJ/uqIqC5pNvcrv9vCtYNtXWVR54XC/OWohZjy
yio40HEacnC485YIrHtX1bM/NtJ2GpOHVJU4yejiA26ZkmGjoBKVc/xuO/h2ZFqu
797jd0YJNoxw4RKZblIc8kuPT9eMjjOOaw0WCJig6Sjzes9dX/6mHphpv3tn4UyV
/OA7XpZGdwTmuufy58TYoy1bgc1vVgUCR885pV7ei+126SYrnxvqQ2FqxrFRq+Zi
cLDxvE/3DZHt3Dqwvh7/qV4t1bfqIXSRdV0iP58puwPh+acT2+sE5WiZUbZv8Ggt
m9kCLfSeCqwyhTEzfe01ZHyD8uqIOrToTOKTqnP+5+jDmkZeRpX+LIYzJs/x8BZz
f4QJW8jbhjeamBn079LD+5zPdiV26pm9jIrZg7t9d5xD9B4oxtYajotushxiarsD
cxQVuZS3s3df+MN4zKzkwodBTimmS4T8X5s/iYc+bGVB6bowIDULxvr7ReK6b8W/
klutfXfuRNCb2mOP8CROnPP9APzK4wsTsaxN1LTwJIsQMLqDPItKQNNRBMOY+uso
iJGJKUMRBcmGgJJhWPzvLYhzMV41kqYbWGwHg+pS0TRrit1bkn+0gyl1gZ/F3+BO
XP/0/eOjzX7ZnsnwSoPRO6Bx+22wMEPDfOtqz+4Mf1cWbMygVOp3x7ZuvGXzpGXY
iEMrit7tntpuYflBOf3WyaBPMkW+s00BRfMvYOyHheLHZEnV4lJ95NCa/sY2reiT
wRxovZbBcd5OKQjOaUcIIKoNCd0HLjWzPvz3tC4lFfsS+YaIZOLpuA5BWgLHu87m
gv20VQUzI15szp9tJ9pSfpilc2KeeWYojQm/KB0hJ8kEDzNEBq/xhAb+0VaaAfz0
7Imbibc79+gmgGEx/L0nvwh/DxVpDLflX2PbVJ6NnWe/FgKWikCihVMZCAjJ0lnC
nxAPznlAIPQTenT8gnaIi73uAf4t+dK1qu7FDH/6D4UkYC3Dn8V7y9zaj9/xtWUq
KFFKWmM2lK7+NO9SiDRh1IWV4dQ4P/0K88/q+Zeo0g+NjWT5+DKUD8gni5hL222u
ds03hM/MuL+XfaQnvFxaXUay8/3WuNoY9+VKbA3Syhcz0RttCIIFCMduf37plZ/w
XFRUkrZY/EDRQnCc9DnepzeCDBjGyBJN3rTQl8mgeKSW34ruuQuzRCJHncEAWfHm
O+jsFxpkCuJqLIB85ADvcTUmsswE0wGwW33b43ZxuLqYh7Yd+N0ZmvUvJ8QaAioP
Alo5eGQ2k4StR42WmZ8WfgDxW5YJ/FFs/XSeQP1pcVNKOhaKPa+36sLjM1mMQCwo
9ayqXgWpDT6G0Ie7ufewrf1XQjoEU9BZDli27yAxXNlqH5Pb1zavQ5C0bJ2n40hd
WbjGmG1IKPvB7HU2PyWzZILtJqIgBC84FGswg0ENMuBE9Y4tsTg7LDZLR6nT/1r4
1goh50stdOOkrFq9aijPHMWN4aeeCBKZ8lkFmGQQknD0S6soKSrnr7S9wDTRIsul
WLL/3KNrT+hzqui+pAJ/4sL+Cnl+0SgGS5Y8iiVouVxodlfggCk0T7DK4QFf1kVu
1p85NxUvU6Mcrv7pD7MFGDspz0qkDIB5kz0jmsMobqz1n3JhZgUMNEOkke3D800R
yggf3eZa1s25rVGI077ctBcAUTKc0x8afMqVEY1A/oRdRVCYvbmVBVAP3DJAmzK+
8dulwaXMvSD6xGtLGva6xr3pfpwcTJuLmvYAk/QLCT/Tvhu/+Fwi3kEVFVK+Sj0i
BCOI/fmhOosuxCWaCACJV6Cuyxz9tlKNPeLG5rcXr62YIZw6JwNXskttbSJYGUPM
EhvEhhbkK2CZYzpJnCbY5X+INpMx9ao0/0E/Jmry2xnF4tz6KhfTj9RlSmCiD4q+
mSVZjadg5VDGyH2vR4DYe+TrNBF3n6DxwBPTlp6FvFm6P+1uBeA2CvAJJSZKINsF
RTiljSC2gaOK0Mu4IyvzqW7+3aVRRovnYwJW49pBvslxI2bSnzHjoDkA+iNdc2eh
uHpJ2PvNLZAdfHDQA5HH85tNUcpSRLnCUP/+1ah7GzK4EsE8FmevRCe0U0+WRHEd
WJkVbeIw7mN34w+QB3yX2wD3/pcQUdpbpQACQfw1qSZCbiTA63HSkgAQxr/GudD7
KTVvB/NDbUgGsceSEAIIiz1TBg3Qo/8DtfXTvLXoqDZ1OxMj2JF4SEs+BhUuQBzP
fG1G4eU2RxQa/ipEHKACAe3fN06VAbMtSfKQJROW8Flb7IY7UVDhOUTXY2bjhs9q
2g+duSj5yeBKQKZh/yR76+MhenT1T3hRKQwwPZ53GDP66gtIAgXmvd+jHQ+QisrC
uV4/Su/sU+85SXncuinST+RPK7Qy0yhcKhvlKKJozXT0BEU/cfANlqSJry8dU+s8
o+FMHEcxb4zxzmGq+Q6ICTaovhhCgiZug7yJ6dtkKLf91eyAljzwUfC92+lDUkQu
N5oS09h5C99J23JenihGSlXXBba7nyGqO3YqLCHzxOzh0tfmyDZM/kbAVmtxJwFa
gwss11TwILqwhULTbU3yl1eoynQ6iE/hyogoPnGriXJvP28add6HM5XjI/UNz7yv
WTZSuMCZ7p2WmzMpstb6XuTYCY7BxCNYljNAtX37mlXAvvtRfvnhFqwCBGkikIIp
gKp3NqTBTZrv7doxYS/WHFjpbDtcDA3pe5vr2M0TJPiljhD8mNTKR6lU087Lg9Ky
u66WG00AjcoMU3tbd4qAKgDSLTRklxmZgOLyPTvObERwBsdfDvhthhTSNdX/6oKk
QFFegOZqJgsGmtTftIOWSn2/eOW5Fb1r19SxOEmUsmfcmowq+Kk4YHxoiBtIfhiW
rqLesU/+4xYaL8z7fOxP18PBY4f/NTWk5RjaFnLmzjapwByEotvPcYb9hCtdVhOh
KDo+MB4LzFToRLhek0RxzWjJqBxToHedNVLFWN+5CVxk3aRHkvJVuCGntdcEl2gG
kNtd/xP2T9Y8+OTDP7llrm+DHiQmBSrev5fDF5eqNrqeckrdJ9OUwJ5PDWB26FIA
r7A81KKfYB+LWysvsKIAZlUvF0MJ/I3Luuhq9Q+V4Rwojhtk3SSj5D0PyiB3horT
wsk+01eP7/mGXp+QxNjlFeSxASulPCEowvFf8ckgjHaDU3Ap2dCO5Cr/2oZHyWsA
hcoOs8TdJFvoZEbCwf+jM0mimdStwxpYn1IlhantW18TXF1R8nuXm5njlzYAaXkS
vNcc7kE4ub5qQEFBZEN3/3qPnEcQRK52XhjDSSO38hnS3yuojksoRQ/cF/9q/aZm
m346Ku608/MK7XYo6Pyi1QKtpcvv4fDzrWtprAGoYS3XovTm2BsxPhkbawQ+Eq5B
LTBOqMNnpC/ZFwDH5HulISYEwSD5spAwGyU0tZ1ak0zl+rv+emg3IfQBGimbrZhP
kf/WAAvZNi/lRoXzMaNLUZP0pLs3IDpdaBEHvgWXl2sFC8bToK0U9s85B6MGEasC
/zODQptIjFxO3akvSGuyK2Ka+e/vx4owiYKQ5wzyS24ku5Z6ongtDg1AAO11Uhy5
Ji6UA09E99o15M3EeH+3GAM1dQbANCkZO4iflphLRNcIs4A57wCkdPiXQPJlwswg
WQOuvI2qJTVMIcuSM5Ay00ONwRnmUHxMN6egAz9kCg5BZNir4wlcHw1/PatoUyFo
6lzUwlSw0xw+cnX9oOmgkXl/QxeBdfxY81zKX56L7yKcv0Zgqg5OluIGIJnrgD4s
AslO7a24lM4dWKB+PiSpzKvr2PwNJD6+6tTLKFiueq1H737aEpyBEhfn6dvaF6Z9
IQZc3QC5ZJA3FEqtNjOOdlgfU/iJ6bMlN170UpZGLUx5Frqcw7OWs+sWmHmgYcLg
nAeYZkfeR0Pej+dKre/1OkfMJJoDjzyaQbCAH6EPi1lON8IylGlCgeCyFlaxNfkQ
W18F24ptfK/OsIwZey8lAHCQ+Ca7i5PdFfwkcUntwXHV0Uq2QJLhh/dCClqWZwGp
n0qTLLKYlDZKJqcj+5JedWkK0u1vn+wnzFVi0NOF7H/vrHIgkQeF4FrI50MuCWop
11vT/zc7/AeGxjfjMJruMbeJB7dD3v+vshfjxATu2AN/Wh8Z2luAi2UpDyT+Mu6f
t5saHBQRSQt6MHAPM9vk0a93Vv2e8t9LibAiQfvww0wOhIXgGnlZYonYOFEvN4Jl
CN8hkxCboQrgk4e9q8cWphODs0Po98sK35jFx6lRuJd5NK6wfg/TMcydkatgNjun
CrrPh6ovwXLFn3EEdHpNE2GVQJvKnp0/ssw1fU7DLVEAwNj3EUFbwbvFLWW2pbdi
j89F4nZX+MB+mqx7d6nA+CR7/srydEDFpUqRNX598qGV4A9xNcESN1TntjYQIIas
8XGbqrlPH/0veaAUPeSHoiKnvja6YBsHdijMsvJnVC6gCc5n2udXKVmXF8rvUqem
57S34SgCcACgfLnPuN0wNWxGz0qA18SvpafluDywwVupx4Y4vkjM0CbhXIw23Wsr
PxXEMBZ31837VABfq3YMwl/eCZzzQZjyYrww0oU6YC0Id13wQpb8mcnBEZUiQMSt
iliZwNhAY2JeC3V4yAi9yCjj4cfqeXMtam+ou2RWJykTYnm+PE/vRU9rEZJHQ68k
2OeGU9KkgYda6wl+7O3zuamwXlsHz8R/vbfPEYou3f5lcOpz4AvZMHqis+UB278p
ZDigo4idAmPlo3Nwv3oGKgVtV3LfMgwZxhZO5JDwqqyyA2u1VVNckdyBZHh1lXqX
mdj3P2KsW3iNhSNkQezaRKhcq0cbTzXXg/T1kiiWBdI5bOafjqKi1uSkuyG3Onqg
w0s6VmcG/78BDKJdQgPh/cVch00DaJuR3m8Y/kK4K1CQVrn5mu4icYLa+aTe6kuD
1WMIo+cP9ZVCx7o+p8Ovge6uwDUsNGcJCOjVTzOvN7x/Lcd7ucGKunxPoE1Hq8nO
3m9U0SF2nL/M1A4504DAoLpLkstbEUNdq51/d/hPnj5dvSDt8TxO2zxLt1jRdQ/h
bvgxpgBM4hWbnFjjca2DoPc31bsHWXf4sreJbbQD0b1Y33WzH8a27jxLaJsHCLj6
957lMIfkbjcZSCg7NVmqAbs+fIx4tty0AcpkBYkCQzNJ5V4S1/G2afn66kdvEPil
9r3FzJ8qWIMGsfNisdY8hODCOxI1NN8mzuTS2D5U0PonTkJVEVuBUxJDXuz8DpKe
V/OdQdSwEW/thSNFG+FqY8qFrZPbA7yDbMGimDHWZhgDXXiHfoCqMGlpKHyIvJDR
qk4TXdCGg6+YhqGg7wVyx16AiBcPbhHNvRbSJxshUv99W7ADwxhHXWhnSQLTJC5w
jta4kZGgxp9CqqIWTCoQeFt2NWURRrM305Ul5WtSulJweAwD1MuNG1CB6MXBN1Js
saS9ANFNRUirQqi7WOHf0seGZaIzH2hHDQIHWS7LH5kh+Nyowul5Q9DALAZTdtxg
3xDMJLAEIjfF8d/zGmXxatyb4W1DDzuzfuiimAM4DQtAb0bkrUKmAuCHPKyXY4IJ
fhTlDrJSKIgcVHUy+uhKWbdpkZrjK1jMIk7/1KHUEfpb9NuxphwPxutW2F+AJc1N
Ej0GJkyZDbRb4Muv3S8hGy6orX6Yl2Fxc7E9GY7eCVpnIlmdGae0lwNjXJS4MvoV
V7hp43OMO8KdcLxFlzts4gu9dPp1lMGI9GFttOogxDNjtnPNyYVEiQ/ceTV/c8Di
14KrXkH5r86Paz3+8R9ALUkgzb22zjZpmzL81CxToWvJ6gIrRg9PKUuHLNBFtqbF
qSoLcFYVylcsHL9zCO6TOjeURh0hvw6rx9U6auHjJutG5vuHrDQRsI/p8jxTT/XD
7uwwusY6IXaPyD/8jrHBSDqy2LjXeCaxMnZzuW14AnA89FqOrEalK7+QosePBco3
ZFui16quEu8awo0Uzj3Ek7Ew7xR7Dnn8ajY2IC5+SPZZzML/sTXHussEWyHW6UOv
toKU2/mfmStyOTFMqyFFSgh1byxHrY1PUr+IbTzbbkurOrZ0AdtlUZ0wyHqXrjtU
J49v2xZwt5lmUdbSUnT1TxZL87Fg2OR4ecqkzl43GyoAxWx98k8AI96isCayE2X3
UY49Aa8XJd4UbQaBz418b3sybY8ndny5dHoY7W0nMdLWKOsNFiEpAUjo/YiEcLQc
8aGaS/mbBaFxY3R8DThik/u8CEOzrm3vtTUxvvCl75xrk7POY0oyguGBargXpfUc
/HEWXPwZS7j0P6DxkFleA57oVzPuiYxy/RmZSLPHiPXQEm0wGNVdWDg+MI0tJ+pr
ma+TtG9sC374sYN7m/yZNvN0U2VoOclnRNoBR8Kt+SIsbzKVEvO9miXJ8bSwXxVB
tY683Nh3xtaOaVNvHcT7wMj4dFwGznVG0UIgu9/BBY03YIqmcCIVvzC4yykK12kS
LB5BsB7S109bso2vgK5O/Np/YEjEN5/t6y6zNMKhuW6Eacke7++AucjIAB4rbT4I
M5eHIXX7hbW7BLq+nkhs0KJIk0XKKQD1hu3tHX8I4u2Vzq0XSIux7N2efg5Pk4Zo
btjK99ZPOF3PLyxOYW+wRVTHmEujTxd7qm+OuUy5QxnY9Ujp/ua9rWKJyVfrWLiY
ETMmfrBs97/I9bjYzvICe4D4zHT0+n7FyHM+Wj3IKPeh/fmhmWsT+a0mDFqAqPpb
uV7fVSF5ATfQWPX6Yc9z6CVv9X3Qmz5ZfK4XTrhqqToIttN9Dq3wQoVs7dRaAEgP
B4Jp2U6tio4zoMYU2WeimqaJAypOFEkFiJm4JOeUuspNdI2iq9zNckLP2xJL4u6w
vSGPXc/Nceivwkio12xmFmD+2rTuWi7pBDTTAbOzzX70mTs1/U67I43oOl5cRZJn
JLaL84JpNPJWf0dzbCA+MBIvf5EUSAN2sQbj5oVJM8tHJKghXignJiZ8upIZoUnN
kCXh6AZblChYicVcHPSthml65INVHzkRwGVVPEysUbnYGxyF+SCrkEEvpde8U04k
NY/n/HCB3Gh+RvXHURo+kWaSLBHPkh6PFSpeRkXBEw9kBg5etMO9h4FaRvbup2b1
RdnKnKegfKF/6S5urcw4wRgolcuZcap9+wJ9ylJHFCEOrLA7buSZ0jloGJCKKk15
m+I05ucB4RkuZrkMZ+JKDaLJmY0WYmjHuHnhkhnzI5zVuAUjngM29eDoBYsJ1AW2
r/2ea0vWn/UzRijm7AkJmh0i4v5/CSdf5xuiSDnf6/eb5tE0atekcdSI/i02Y7aA
pyClldmntxKJZBrMQC8MNI9VX6x9zfbi7rdFX/Dl/jMYJ7NAmHxtf6kVxEfLJL1j
1NB2UKpgsP7qvmI8uceFeikA0oblYvBfaopHTQj0XVpLUvj/EqMHt/9tkN4i8wWL
6Vz9ZjyRSZBCbwSwoNYVe92lEyMYB9EmfzEqw85NQND/ceSv8hvj/YCKEiYh6lTq
4YNfNt625mctieasz5bZWRPRHnIwjhi1PB+cIUZdTmYPNttdGwujA3m+aSWdHfKk
BdsTbeEyRKSADKBWJjmpvN6cwgkWbJgTjeIClu8zz9nyt9RJL+O65JJ1Up9CGgaC
nZh4HBK+KC4w7mLtYYckKg3wGeOvi7k7xbMpI9rC9VdAlwQUBdAMUfWUgU9rqHEN
WcwTE67M5Q2t4iiC72nhl1NcaHALW6+MI9Nt/iw7xMwwpKyb3lEUS3+QzlwKSqbf
8yiAFb5MiEwciMbN2YVeZUChIAyOqbOLPvyFCyzrILohUPBCCR0jbyLiB4YSeSpf
CvDeVYdc+hxWlEaK0kP9KCkWhxFC/gy9Y0EIPgqEemEo75YIgQWNBYYq9T6Yp2pI
bBgF4CFtKc8jtypV226OMzeaD4/Ml5dSuOA4RP55vUPZfott1L6IE1YJyxIwxJAA
x0+PEEbr5skhl+jdCfkYJuZ2ranK6z1Wx4SzkMYHUbBdYNf/TjUBs1DlPfN/Po3R
mETUE3COb3r/oQYlTtQhXZTStbY2Sb37IBQgF1Rc9oBqDQHnoX1DOQW6Up16DIt5
RSgWR7drarRFSth/arUaf6Lo2ri77rUUAAkkQJux+EWvW61P7ZHjXOrlX4ameZt6
zjtGSHuH0jABN4rLq2VInUbZkqX8FwDhWu+7UtSf9V1ZK3xQ86w9goS/A1Z+8ltC
kS71+nPCKFGHmpUKE7zbuC2wDVrQCN73uKzF1ceB8yqYNjyJDXkXMwuPGvcXYYoP
JtAsyYtsrKtZfwVhgHYCPkhDeJxR08dqYn/0cy1lYwhNuJu75k7OTGZ7L/dqjI9Z
WZUUTDimXqqcA3kdJh+D9zhEPKDrZHpILjX+pufDD6YN+S5DfLDYiJYMGXTRuy5W
bQifhoT89ARAWMnJoxX0AWSJ0mt28daETc0bzXk321ANjDoTSA479HK19mf+zVQV
zSnOGe10XLBPFCU8Nqhayw6ztaJBAEFK7ZhXRQZxlgeMFazkNAwLR45rJxRCbDuU
UdtObJmSs+WVicMgrKLihdnBKavrkm6pgdY4lm1ueRbCuCzC9vS8f7j+RaeQQTLn
1aJnwMTi1Kwwq17Ei+pi0MSWotXPbGxnwq4AL/ju2qYWVhAXQBp2MiXg5HdcBnCg
o6nOOvfW3yKAsHO0MYgNWITT6xtQOAw9cULcHlv/xLFr0Bo6tEzA7C/aaPiFuk+9
4Ld1QhfdAKsYEyonWxadBbCNSolTedx8VCqD8JDQi6X31DOeVl8Ow+9P7EPUeInx
4ajQ1ZRxnoSeJ9eLxToHbBAD6di71xtdPHoOGkO54VTKii1F2nGi2nEqEI9R/78k
YmaXyYgJCmzJXjjM2nuRo9alwaBNNDc+nboQuXaskodw8e4MOFpjXal59bMJFBUz
NxF0YFVWBGJdHDoo+xsmcgNPZ8Sq7KkVLglJ/ck4T0RAVUlBek7uIb64HCfsenBt
lTRpNrG+Qd19g0TVGc0BflxsFax6Motr7ETVSF4kdYi7+KxfdRI44bvbrw+nFcL3
pztlk+svaUstL5F3DC26Xoa91c15pZN8BFaSBSFASgZDVXqBgA1aVzx6yQ+utzN/
kHfIOIKUDuN+yy7BtUxQ0zuS37GpkJfiQPUAoE5FQsaylpIQMn6nk+cwJvkOGlvS
nlN/3n8FhHUbvewWvDpuBmrTro8Kfl0cx/0BUREHGuQdHS7s0QUpF3hKKOizrRuy
NYPyZPP++0pDYfUyTiStlDTqP41Zf1cmtLDBP+rVYqM95APhWHddBhLgiJA+aNBm
5LavdlfCLiIoyY3h/IrrzIq8IsmtB6BHfSXrvTNAJE+FSLfxAyBjIjlgJ8pZJTxc
SfoA/rSfbIpiQ3HKIJnZSlDhRJ684WljSN3D14yVcx7qQCEi3vPu7xpzk73IO740
39Nesckg8/0v/29MFxhmQDdYxePHCoiSV/c7lU6rYFX4pnAT2Zu3O8DwAqpiSMEi
XquA+p59e0unuJ2gG4x22Sqhw8aUHsWq3PEhN6UsNYyO8B/zRXZmAPobGzJo7Ylh
Zzpqcf3srWlsy0N0iN1HW4d2QS4dsh+eUPQ8oisztJ0eDBT+cMoZ5wY15JsxQ5xf
xBA7lPsrFY8pvpmDKXxbcNMdW0f3Yf495BLIZsoGMznTdtACD2LA/In/w46epn8t
BJd0qcrX9NYnp2Lp/1dnySv0STN91D12bZakspEyVbNPy55P/kZWJ2klKuOuA3Ru
lE48x6xrf1V04oBnDkWjM1NH0zQ8d8+g9z9wXL0OIaETAvp+bF75Q9TYq3BnLjX1
kLbIlxIoH+mwYUR4lLpF8LpGgIWog/eRh/v5qRH/p+BI2EmXrXXAyEuECPW5K/NL
bBlz5KMvNr0mJI4lHtK7DJLXF0t0YymDj4Mq3WjVmGwMEOE/Xr3XwQ9Be3mV9kPy
lLYs5IBRLkxKtKn7odXGzaMihohokuD6YhMCuF6Umswfy1470VU10Wzu1C8ySI3O
5NFybpu9mykmzKmakZuhCZL/17U8ElkOFOduLuHnkl8xo4LIEGyutLvJ5wjC34YL
+3tYP4F8CDa+7ZqqVaX34ZR2D1hnpQGz6x0ZS70pEQT8zimNKxT1lzzilmTPCj8v
SP9dQJm3QZNUgOcEFiatBTIjBcZswL9MRTsZpwZ7xCFGiv5a0qLK9bLTUa87AK5l
wpf+aixTNGrdhiP2hB5ncrIjrFK5rZ8XEyikATKIMlRZpS2dhnEu5iv+5YPkkY4v
ohSoy7HCs4IIdBOGALMXA3y/PbR22EkwXKJ/9kBcKvVw6c47qUr2Nt9Xu5dFek/j
hWxzxG9bwL2jF+kO9hEsKWvZA+YJ4+6+OM/weP5Lw0rWuYhO55TRb0iFZDoZaskK
psWz8TqYp+6xdtgnu0N/23EhvB+YLekzhh+1u0Tp6Uh0QPv85PIBICOM/KlfSbFx
EyzFb6Oaewgmj1T47oJ3sQ8utceLcDfdtXVhKxE3n4ctdLynm2fsQnYD9eETuivg
T3F4eyhmvNkb+Rwulh0jLV3RSDXb4kIOStpfO4Ecf0W6d1/eiht5pRiiMzzBl7Rx
/EJ1B5R1aNkRR2fBMpuocFAP4NsIkp9B9nA2hBjvQ10gBvWmgmc2J4Q8mnxJxLlz
MwwFLfOR6Tb+7tZyaNYvWLscNtoTFIaYE9eGGX39nQfjf+kTnK4XNWp25AcUyT66
F0YHNIyc+JBq0Jfk/UTGT9lG1GARPvta78vWJ/pSUKe5iwYeC5GeqJyhA9v0KBPO
zqmqI7dCJviKhLmxssxu9FwVghubrWIUZWjtkyRTd9CEgj9VUnw4/nhqG5qYvLtu
mZwqcBH6Au4D9z9gi7iXYaJ3IG705xqwz8klhnYi+GeD8cA5355Tm2RwRgasrbqn
xVa0x8JY1nWvn2e6/+MjLpmGleQMGmB9vEAISOvGmezyOMvI4J/Wc66QA7Zlt75g
Q14LBQh/xKcw0kxhdmmsRvWFkFfGSdE4XUYO5/KJx4aCh+RlypD9HjDpJZlXvRNI
auOd6NTDDuENi5dgyERIzj3ZVLCoa0iHV7EbvFBFqnehpSU0AYGthOYb6rwWcHPE
Lke6vmbmvfGg5T4IB4bXIrgMiZ0UVyEetp113DB2AUguMxf5CTgN4tn0Cov9EnDz
jJy4ohIoFE33C0GjzhHrexJW/2zHHXovIQbQeRdWCBpgonhmsVipCQsCmTGRMI7P
Ja06LWUmkH2+/nbX6ATiYCkX8r7UgQJXN6ilkSfwUGCpaoRqJEGMR0dAAB/hy4Dd
4Ktspki2ZRYKfR0UWSU21HBz+r3y/v8aK+MYhLmFAZQKTqYfC45cHrxBksBB71aP
LBXy4UMX5r4XAYT91Kxeu0XiiIz6wtKRgSoae5t5oUTX72kwpOwoPOpmmgeFPZRy
qaIa0yJ0UrCUvEaLwskow3lsEQs+tVmMCojA9XC+jqeKnKrHcnVNDInaZlwEoydE
lgwIcIyouEnIQtHwrPZkl1yn6wD6zy1I9qI3czdyvYF94TiOusjGWefe+zZ1b/dt
o8AhVnjM9/GFQrA1/SKSIuGno590Rbhr6PnLRBYoSBhx0UDW1fOTSwWLzlSWQ17O
okdr2wZQnUqUxTHam/a6xINXvfwE3cJadC3QZl3JYc7pt7ER2U5E1UDas/1JIu/0
rA1Hn8nPI1ncxwvE7UzYPo4ZoMsV2X46AShtJczXtkSljpBUX8w6xLlXxxLxONY9
6Zbfem7Jga2nwLTPKuB3AU2uI3PWMA4yJVLC8UR7IjqkFQm7GTKxApjQPwXxrHTa
JNpoaBKsweOMBs/L44G/R1mg9umdMHguTphirrXzxqbh242da/LfJKjhr2O2DRut
uiwdGdMc0K0DkUTQoheZKtkfWQI2hc5ewTazPQISstYVuHO4ZN2dUtrT5z5HIFo9
g0ZFQZhO4cteWn7FT83rQEsKtJaD3YBo1B3g7FnZCAVLJKH4rf+VCOgvz52hVl60
sOzCFuanHCECXwnLBHtpCoFdQmPQhIFsMdlBwrUlhy+BlU5DoqhHvCkMY/02q1HH
fGNyWsgYG4+MRd74f5CTmOt9dvR2uSDAykUcvJ99cMe4Ae9ZHjNyLuOEiuzUDgLq
kqL5EtOm6LpkbK162M9GLy4o+wP6AklqIiyByN6qwEBBxwwZH07wfK8ENHjJ093U
XyXtlTfqGTjOCeVd3JEFqVhNjCUvjmN3FOOqrh1Sndbamsr+DY8Sj1yCzEzuj3xi
/1fAooVtFdi0GQARcDmUPhuYJWeyQzU8BfloY/HANxo8cuZMveV32vT0ap3vYUBN
dEf7zGFh19QK+aUpXqKw4y/CrqPjjQFx3DH2a2V96YJKvPcvdLntpYn1nzvN9e8K
ps7xeKt2RJotDllFf0jRh13G3egaDhfkHP2U3H5ORqBvhdM1OkL9sfEiP9q2DP2f
zsWDcPUdqSvpJ8og8b26XQVqL3kfJ2OKXaH9NBGBpKwoRzrtb6PZvQpcKSZFIekQ
MYYmN9xKQjlWhbJrMpf87JWkTKJbR/UvvEncXokbrgqf2CuNCMVtBr/8zxepwGPM
Hagb4AvGseomoMUsjULOwo++JNd3b68Za0mu8PgJ7Wfvdctu3TWr6WRnE3yOnS4I
nx7VkP9T3fmJ05dA9eXOOdRIw2n6cgUqypO+AyiB6z6cAFj7SF+tyZ1hxN1d1cau
T3oMAt2ET7MS7buDMscRCgqDHa2SriW58gkAR/1WeCgnjHpISyuX/va068b1C/Kg
ddIHW1ZpH2uDw4Ye1M7vC+Iyd/fNJNdcCBkXR/btPFXeKuUwp52Ut+VmTkvkoUpv
zGh0Vy+Bt6rVqcdDIx/8j0dMrwN9RKpH7/tNAbosvo99kYBdYpCF1EJd4iwTKByX
dZcStqw2K1+4Ya4U30zgkUpJylC1yATVown7Cv+79c2errk5WNcTNAATBB52PZNu
ZXXiwroiFW4spATDwAAAttOagLoRK53jx6FL0Uir+7Dy+paYVBnIu1crJZhM6Bvs
6nt02QOX/1IzxK/UmeIZZ6UEDjf0Z7fcVAfZNe+8YrXwrIg7zpFAqUvT4AQSQBAc
RHGWjQ9sNtJmClUCmZoM9vOPzIyLZsrseyfse3qTTqK2y1AMLZLp7QhjLGfxFrV1
ET4yEctD53He/2YZFZDYuDZAvf7Aib9sokayw4ZDvdZgSF762r0EDsigFNJGITI9
iBY+oDG4lx5p4Qr1XK31+PnqJ/3/OCe+C4UBrQuXO4T0oLeV9t9sRQZ53ltorzsr
eOc5WHFoLtFim4400GjfHQqvUxE/cKSztfQ8xX+2CyxWMc8bYN8lsO1J96l26zb2
NagpOqSCeEdQ/ac9dnZWtuuaO9zUlbw175FNSRx2SDLao+SuJe3LGKLwd5kOJ9eb
pd/H9WHWFG3/d2yTAPCQBL0xhSFlFPGV+bGseeUDlR0wpvxC9KOmUC329DcCl3Q5
JUdpiUvGtN4Z+d+lxvfx/lBJiRmu5uT53/5bMH0gNwdAlfwgJ85pKrrcwysEK+1u
yZFY975BF7e/yZeH1kHdOFsimk8RJ3WI+nTE44RiDVIx1I7N0h84RQPyauboNwTd
+7+B9WMhYT03rLEEvMBj2JGDo01E96zeg/HG7oq4JwfIN6LbdKIWnwg57NPl7MB/
4wlQAWAP0A6jT0yDQpa/6BYhXtymR8K3XFqCdUnsYchfBNuzhBLsvg596LEN/sEw
np+w0Mr0A65iCUdF18N6BES/Zj1dVqkQKSppzU3ZlqPGECly3oSnZQYskspA2rke
NWdWYyzJ/VIz0RxvJX9qYCcgXqHM+PKAjgllLB1NuzX5/j019giDsscNqG9AgPZ7
m0ilOUbBtoo5AxzXUVWLOsH0W9zVztXCtPeCsxSPTIO0YrV3Z8We0ctaElaMVf1N
jTp9wanodIfKkH0fRQJ0O8JdTtZn8BZksxL+gwqPBkyw/K10wV4bgdE7Itv0yJEd
AQzmd9KAimW0QkoudHBpWw8Fadf3HNou2HbaCNx1w/UcLFrdyr5JFiJUyVFEhfzs
NuUSPsuE6eukwtlHEedLMH9CUFSPw3a7Gsi2Tcz5fvgmpNBcvvH1nZbgJ1RWCJ3I
EnmcjLkxhAmWT0S1dhqnH04Y3uQZU4C0fcdx7QUPgA+3qfaeI0ADoRX7G0+OwNik
RZbdi9W8MX6IaT95M0s8kO1xybxDVXPSyeK3vQIpS4Db4SF/HHt+udQ7c+ROiknu
+iLvEwy1EDEbdQ5k55K7QQ3ysQY0p6qhcZL0m+mKKjKQABaRB7Ly0N60ywIq6bqj
vn/UqCZgH/FiwnBdqhl8durp/0Ae1gAV8SW49GzA51bGFKoqN8z3AXqkNR6GDVeb
cOR+E72SFnCH9fhfvssYgD6+zA/gVl6cc0d06mWM1g8n26/Aq2rOVWcqtI2lWIIX
v3vdHU9mnIDiflCL8XtSaZu1udTPV6pTaSS9pJCTbIFMTzLs1szgjWkPVxeQNf/M
Z0iK7aDV7wwuwi5xiWekzB8opGMX2yjuZg0fjdkbSHgf19IclwELrZ1eKI5BfzIb
OykP3xc2Ne0ONrox6MhDiZLlv3K2tYDFaxYrLU6hGj5JLRfaR15TFGvXIOiWA+Tj
vHDVYiPRDCcHUA4yCqOsnuIo56dG1yFVfTLIUUsLBA7hTtk5/1qjQzxM+Y9/9x6N
Zv0BA4JJwOnT2dTB1KZX7zMEV7SPRuEuuT2XZvbv9pbzG+2jDtEmXhHKWrznzYD4
5w1LyaNXWqpxcGiYIEd/B6MDjVeo6yWQGY7oaq+4MOEiJ3VFJMk1cHvrUAU2weSR
Ih/ybGFvbotumlKIcHHjJJs3BMFS5ZTseiBZ+u7cv908l8//bQ6K2cmPw07jVhl/
0NTvGKsMiqSnT1/DKZkTKCeCqs8GfctSHD1g0orzmdM/Mrm+sy43o+2Ra8bhERx9
MbALHwxQxBCkK9+amiENi0SYcK+h3SOhlO98T3WOmSwF8hurPvdMzkWOLIR+4NDj
kAf2DIa06deupyeMydAXeW7MTfBqAfkeMKssvZ6BIQJzzySPTz5J8KgO+aFN+s0B
NYPMN/Yrs9y1rYaui45cJL10Pqq6tJjoTeWPCzsLYnBMjKRIDRrcPPTsxMts4reg
jYcntuteQVzztxN3FqPfHYFA79yql19AfgaO98JEzWnJHx9Rr8SiT5MZZf7AmDU6
kl6cX8T+3+cFT6RasmN9xPes1Zrcku4gW+icwQfMjbYtD7oYtndhDKbCOHmd3ZQJ
BMU1/j8XL9McIViFk+9iakNCOUhB4kJpHdskXsl4HstkqLKPBalc6L6piSvtCij/
aFaiIgzouwpi3lo/j2oJJcbvMBvZ3y3Pwvxgskkt9Bp+yXEP9I6oIqDyHKGtJAqh
JMwphgbQC9ZAfBfHYWjUVRDnU/h0K3y2+YqcDVFfY6IOmbjZjKAgds1DdqU646+6
cofNQx02p5Q6weafpXlAAUm0Sm334M2Ipqb8er+JvaySo5QBEqoCTwe044opk8uA
LFSF9tCaK4Jm+q8ko1Leyg0QldYG7X1pby2NQhcwnUl+06PnqOOviQOPldum3dzs
RiBDVRYYGswHnnWwW+a8NfOmpphHPHG3t8uAFazWi/wYXoo8jJEyxQBTWvjcGGMy
QAwOH0QGfJ31BvI/P82HefKBCbiBu9k19dZI3LiaAjZoeh5b8gKvmlwH53I4vvbI
UOuZ4/JXFRvcnSnPx/C8bEUuXQZxoM8jDQveWCZmVD9p6mtK7LiVNXwIlhv05to0
k1cpF2rLezAFadXKLt+Q0Vp+upGlFcK4LgqJxieu8/lz0+O6qtKUlZ1TcfIIyASO
cVf+diWfqLFaAdWqLnf1W4TgtBP82JyOTCirlPBlTz1wlnXFaWS8oqIDMvNE6tJs
Zt+F/9CFBni21LUas32ZWFRndLcB9+9Ks8nhsnkUCtlPzXOGBuN3FLXdP0sR+EU4
o57KfV5jv4L7nZVeikkB5ELEuMmFWmR5Cdfb85TQsOrG9b6apDEHRiq+jQ1ftoqd
cQwVr/q/QPPUcjux8c3YDoya+WiriDQV7lp3WpT8HJHVuxfsJe9An1i8SFmCvGiQ
avVvvIvglOq4EnwEOAFtxwA5yrnOwdNnyksg6nbt7eXh7nEaPDJk5pl1ZjvpJ1xi
3V4Gcqt5PcrAqFYNIq7FXJ+LQFBQRCledVi4NfC0JpVRvNsPuXE/zSxqaRz5sEtd
mwkGa2GemGdLRwEe6ivYfGbVcUC9i9qOcZdsGRRGDDySTRxcb9bGlDx4KcSp3YeK
qd+HaSeuYbwkqc/roMPNVdOHg7ugmecwi2IJjzVS9tryl39v3syLR4toGdm5mbpm
XCVylLbHtmA316Y/aVh9bBHJeuIg2iWIanB3oH38MfvIDGI0Hncciv6bwTuJ2ErC
0P5syFhuvcnGmY7cq69SZ5CxuTd/M3AC+4cFB+AQChjyOHBM6/oa/XNZKLqr2vJJ
mcilYWmAVvxtdy9fLVQF3y+EnaU8n4VVhOi+VGd7GWVkz03Oy/DeaYyiLXZzvo2/
RmxXcrfkmRAOGkrS5syrJXGaNyi7OGXjFU1Ewk5e8ykeV+8HnT8Twl12M5T1u4a1
9ifev+52ngzEMbWwZ6UjNFgmy+CWMcLXe6yLGL+5RUJrnx+daliI6eMBTW0j8QLH
DZoX1UR0pc6emFLBSwWcfVmJCP2UJ7pJNCsIQd3G6uNOfc3bSL4Al1vSzduSBbCX
gI/b/l+Y39mvy8RAlyWUSYqJLIi+aA9baGwa3+kxpijy6PuiSUrc9OMtI14AoefW
eEZqG/78m8+n8Vb00hSPD4woKmd7fajUErdEFctWDbNTEBRTl3GgX6DY+M/GMGOF
5VuA4IL/oVvuDaLcish6EPIMD5INw2avsYT8xsI1d27Sru+Y8ih0Jc68+1s8vJ1e
pioROYctPp2GsGtx0RY20xhHUsXg3VQL8Hoc6dJqaIC6PCvoXMZbi5EjuhR+isX3
HJ403Y2DhnNwz9tJkPYc9dK++LC8ZtbEc+FCwJpWkPUj4j73khVWh4vVx0fo4RXo
W/pWwrl23KtnbNrsObKwezfxQFTTdnJWwfHp11kCevR1HJBVs2RW5BCOvqnkgGhW
770/S6EZiWezYpJpsFwNIFdD4Gb+QQQEaHjLfa5o4VhZX2+ufjSdTBj6IRRfKrta
kimIQqrmYkOZwvUrDsMAGzXY5kNvC6X9BY2eIQ6qy8vLYfhFRhn7ehsVBAczNNBH
hR+D01HilbpSh+BnA0RXA7mF0vuNiOEVK+TL3DVL0ZXHCaL1Dbc/PLKXcm0W07/Y
x+lT5iv/ogwS3WE2jJWWXR01dinrsXlBBG7/wrygqcC7tV4jwBxGoKsV4mOjwVa/
hs3NoYBUQKC7shJQwrLzIcZU1jCLrmG7rk8jIo59sWWjux4YRFlW01zDb6sDrHvO
U3EP6vVESDAd9JKuhgiiMSiF2NUeQXxOp5hDgh2ftHyL0Md6CKs43Lf65WPaUnmK
CThkaFfF/bC2bTm6m7L8IsdRitawoJdkR1pxr3LWXmPlnFOTcJqyKSPpBcxAmvTo
FIkn1+C+MNvVMKmKVnMwAnVDOTBscfkeqC6wQMpMgZg0oS/Sij0B94gm91NQjt9v
iHpy5oF2Hcg0lWOnuiwSG0JwbBeH0z9MaTPF/2eH6jgJYfwID9I/M0gBzbvtOeG5
LaDLlMp6OtttN66KLc/r3VRE58DlkfzEEA4POmzWF2CKtKYJS9YQjZx1L2PoGa3/
ve3b5xrHaNmtDgC+BlHb6A2ZQloKN2CnQI7i0Vg79wyiZYrLj6blZdTFXULxulOV
mTJ57Wr+TSSfzv78JJK0V4+Zzspo0cNAlBb1wnWZ5s2t+9futdKZx1ywvLlLjG8h
j4rPpDaCk3KVYFnZecdrTgeH0ikTJ4+byBlWfAKj9m1QcTuWoP9dSUha2oGe2x8/
hxdJqDkMHJlTr25qrE87ai4ZmO26OA0NeGKO9a46dxXZRHutX8DhrxvSiq033ilL
cVnRhOkcxFF+HZHPIp04Zbu+oWFL7WAjkGDXLwfsEKRn6KEpNVflMa+2YvpaQTQu
SgAytwxVqoKSff9dCJVYlnSlTzjM9RUEht7TGQaQrEKuQuz9/64k9vgNTfOvbiVU
m9YK1eZccyFcV1JNzPcuan5QwXMXKCe99/wc8asdAG7YjqvLwwuqXuzCNFDmMcus
6Z0R2C5tFdVhMHXc9jooksOUp6pSg8iYX+B05R9qazeGIANcB+XIAWyGagNczCBV
HXIyDQ9MEUoWRNV9TmeVdRAq5MZ1NNPtq+jl3Hvuunop1rpGUjXz4yyPoHOtM2uj
2zAMkFm7NsrqPxvirv3tBydlFNtCaTqWHJrkF53pMvijjiHk4m6ROJpN7HeYcfZp
9GZB+K7/zIjVPZko+CfgMn/pVzy/6DKNxx08kkFgO0ciKu/JM+SECfB1qBLrJ3w3
6Hh4SWd9nDD5+qCicjdPL//JjKEGk8Y8i50Svcdmz7ubldBbG2SLyaFcmZ3npprO
f5katMRIW+GRWoXjykaRNJb6hY4t+oOqPzJ9OZJ6qp1wu+dUnT0PAclnjTiuSvHU
iAAxod8d9WIg71usM0W8aV4TS6bqYpoWfZ8cuRAvGCMuMIjPKi9PPya7dHnX0hwP
C2YfG4Gy5lkmT/lSUG89YfoRnQ3LM2vfStv3J79NzzzUulQLCLMge4k9cIV7RBMe
hzYYfuXUHwxB1b4408o36/Bt0WaWxZrV894zGcOS3lw3TnS1oxllVl/h/ZSmkrwP
hcJJff28GD0JcTMlUODG3tMt4JQxNcd2uA0mwpINQhlyGcZuhCMcnNATtuteiC1q
JBfiK4P52qr07MH1MjdgxRt40epg8om8eyctFdKItAOEzsAkLuXOhRflI1qN4av+
Swf2EtNBt0Wg3S5cMavmxWxUNwlKr6Cd8HhFTHJggrhI2Cj96F529eoER8eULZl3
he4FyQdobavrkIrWep1HpVFGKJ/B4fSaDy3u1soDMDgdt8x5wo3aYnXgUNYPb5PB
taaWAdCt6e8t99MO+WOxWiShztYAmRzgo5xwPJmtIO6OGXucMfCHjF0IxZRlXv2S
8fchYoXqv5LODDif46zxVhKL5vTY6iezptqpamSa8S6rqhi0UfyfrPIt01YckNQ5
Ps8V03eEG1FqvnMEGk1ylWkKDMOR9q/e/UfTCBzwwXasSJntNEMt3iMIGwUHU1tl
tk5mK3MpYTFrLAdmcvYx6FriCOP8Ds/vLq+k8M6vXr0o/S9c/ZWeGyRQ/1/Dq1mS
OsBsmoMdtCnY8HyUbU7+oMQLHqq+y99KpuTrhV51BwYohkUp6CgL/Nr1rTkSIeyD
pYNUy1O7L17FDCAmYrvuqwBSzFXND0plZDX72Xajfe0TFGzy1hYuazNaEqiqRWYQ
SgElE1MPVgPZzTtwYX/e4oKVxcgmoc5RLwSFHr+4DuzBnh6NF43AUukiunTwVeZk
TlQx8Gb6ecz9fe37EyAiZ/5oXP3o+46nwVpBwd7lgR3r36tA3GKlXsos3fIG5fsT
VO9/xJ+LafI0pfNrfwcLQdzSHgjfSqj8xPPxUfBJMNjEbW2hZXfLmKE6Yu55WuZE
VYtVq9sBbFT3+Tl/KGJO2Zwcn+YcJYPvnv+NZlvEentysCy5zDSNeZrJc0HweFSP
Fc6BQXd22XmGhcnQ6k+k8gEgXSV+r32Yb9CNQt5FHMZYdpLYpwPpQnU05IEwJR+4
mm0PkNDxk/7PVgXKnJJL4yBWOlT0297RWr3BFAuthzu77sY7ew4CNm15eW1IDKtm
TOOiDuSs1Ouu0YesBixo2KTtyoJmUeGACxzktUwNWn3Nt8yJ3peCFwAce95Oqod7
AP5EXzcMcqjgaPszUIEKCRKOGiMcQwWrXq+exrl4HHIP97lKUipzzLhBYoMBg22F
WYWDpvowm5NS1YhOh3OA6HOal+q+zjMLWTsnh48bi4/0EmG1kO4aSOBiAsbtIm+P
UUUyJKX3x1Sfp2N309yQIId0xOOju9YXTuN8a1yiPbSLptcAcQTHzYWSX5vd4re8
DQTkMJUtCfFXhT7Z95IiaalLmdnVONPrnm/xa1Mx8tVBarM2kKdZJTeQFWAsqfPo
tGwRuCb93pigMjKUloN4xf3DmNswxJJzak4eUwEYPT8UfxDoDYfcEiZy44YFDO8g
3dAqvIz/Q5af5alzZy/cBZTODXj//5pTP+gyq1uUcZZX5w12OTBlEsbf0yOV4f5l
4oCk6ikGaPzJxIYjM0I6SwQ7UtEMYBRsemu/jSi1z2NPLtu2QsFJkhvpGHr8BEGO
jgVgFUy/D/0K8rtsUSAjKdGppy6MBfBPqUMaun2e1XuD5Kvgd+5rzrH84Vv/TrZq
SxyVcUxzrlxycZTjPxAFIHaL6i8J75Vju+ebNx1lFFn5Hoss4ROIqWj5p2bdLr3A
k5pi1HBiqsIWVqefsngpKhs6dvfbQ9v/ZG7cHE0PczQEfOPi2O4OGA2mXuQJrqaR
tRuvqdnvbw2fWjhJCIXkVPj2gkzWRtGDbez36/5Vq61c1kr96ebzQwqtN/H019TZ
m1BBEXPXljhH6gaclpIrgtOH0FGM140D8Ct+KQjkjlbmBr8d38c0k22QPw5tV6Cn
RpamqiSnXHw8zWoOnFzuod0NGCmurNVYUxRrVrbPe7FB3d+xFfCbrHntK0/G8Dua
Ve6Ja7Y3gWeoGCkdzbcSwgab9P7wlPbSP/H9uYTO0KyE3X+fvBFNs8WKyYGNhmeq
oYly2nrK60WVK4MIbIfeNqRh7DY9Q077baT4Qnoqg3U59VTd77gkgqdaz0RExJUY
nrZ9DCq0ramFGDxvcG2qGRoZmPux9HJKAgMFh8BJCoDcZfxelY3x1WaQjNA3H20c
6eFng2p2V3rIk8hu6y04OC5UwwFRrt4GgTM0O4IOvxxxURJxx6g2RgekCeHPDYnU
S/1/aP7ANpiKCHscT5npDRYiLzFiGb8HP8A9Og0kILwh6/shiyomjSp0dh1mb7jt
nC49rXZiT6K22WUGDyEAEozwlBrO3C6nBdzoFkWsDQpl4tMtk+g3nLy48eosBXAf
KZh/XsDdd3jpPdsUB55D81vovBB2Vb/OYYtw3Ig2LdOvHmul6aCHTnhMzN7X8ha6
+9XDsIxrJtNiJkdiehrMjcNr3uep7hX8y8xFI4108eZcy4FRPPY4DghwdRElewFn
yua4vxLQ7fvgY6EevmxKQ0j+0hR5H2TlfHL0Nc/7GHmu87Zstys7OAm//A6LBpjB
oNSnRPETxvddYgH2kWHuB3jEOCnKSrjvbHJ5xaA5DVnn4Rx1ZRrHsdv0LA3iw8a7
j9dZzA6CABZaR/8YxhPZs02qi1wPLQeO/q3BVDub8kYl8OyKPUClNhUT2C0Eco+G
kuXAaAyj0xWfgbs9JpP2roho048CgsXc5MYCTfUsgzq7R89xLykXN5xYsvJrk1JY
Nnuqtebqc5NvgFU/z7eZk7Yn04UTbjDHNYkGQOdQbc19NzerL/GJqNdL/AYGfqOb
tA3ZjDkTkxEK7E0nal/P+vQM1ByNRqXgy5XIeHHoYd1iS44PK9kN8gGQ8nmmm7Rg
nZTMKStZ+alxMZ9MHi+oaYPe3amE5vHn7BwO2rzC+X/CT2Rsbydxvnru1fu5q+jD
5mW4khTyOclesTFu2vS37IA51u8/Vtj+eRTs98YiFe3RowXpsuOxAXNv2rnHJfXZ
HHxFuP1yD7RSDmdB/U0lWlUGYX7wFlW1teHRG672/qLhOYzyAMO8CZBZ8TuEhiQ1
wXLhHjEu8DFyZVOaPTrwHW75mGe/b7EXKaXDX1TTIFDRKixcgGDOMktwi5vk4TP7
CmzRn8Zz2WGRffEWgUyuNnWLHxPlbZBFsA3VxES6NsnZVqfLCnWfOb6O+auMCoVE
mucGlfKGbDoppGcbE1ZrTYy3ODDSwuuhkd7/9S6VKHEPtQqGy14ZvKh9hZUq3SJe
vI2P1QVoSkXEOPnEmjOgbizcxCSX3HFJNwBreet/ybbmA7HpDCM1s2rB7PErz+rh
+HqmKaSmVSVwvNwefbSDnpBadf+u7FdXunLUeGH1tTw6QPYXoiI0tGUZThiqSrAz
H83ATagVnGDIoSCRWoMOX+E/ea05b9AgZqkZilAUajOXuPaCZwou1r6H2HfwrCe0
4rN6zt7wNJMMhoOdayyq13Rn2q2faSwkn26kVBzqDxepCObCFKU0EP3Yq4GRp90T
eJzG20hEnyOoDXdjFny9iOJriuwQVRSIen/L+r1mf8T9HuK6iGSeRHQJ9jLxPEML
JBYBT9tN/LGESxGRz4DRE7fPUWROfbzJeGe94Uqf5rY1YyH8EHiMCsyRQWs3sNsE
v+TQrsh5wwRRprG5pkpgFBvuXuKNWr6QQrJVd5XcOcCwsT0CtSliNoYMcqySKMDx
HNlwPuITEYj5JHiHV7zWawf1X8jsuehTwF+nTvGeFVnWKm6S3lM4tZUcnQD1C3GL
lC00N9PDr3b4Dk5ZgL0rkHzjDwBZuXtgx/mVZVjs7+fdw3+jpqZ8JE2P7Jww4IO1
R8V6LIHO7wQM35qA04PZZd6Yrc8o54p8LUaqSgneyAyF7ZVLEuCVlPZLkVG6k3Kr
Rdj39oJK1EYCyY6e0JXDkus+ddubTaGvAm2FiSalpPKO73qg+gYlHsvevJPQy5QW
l8U1kRD0SvJxvId9O4GhIVYrjtShCdTRzI1+Ynpcq7SSvej2GcdjD6La3z5u++TX
+gNEi4CWIQ/kZvBrYrzjkPLSUjZPzrQ/fhQ9u8DD3founDVlf72YHg+ymNxCnr46
A/zIEfYRXsXYIcfw8pygVMA8HHyTzGvfYiI3f6wxUsTvio7ro1GFd4ShjH+g8wGV
ielM3M4jdNX6ZoNWpErzreQvYtk5/YS/MsRKRTSowd3nGlXK8qIIWgPv2YCBik8r
HTJUJpugkmKDHBL4Xv9ohg7DsuoVmV5VlxlublfgPqaBE8dA2DkUWb60BFACIKsE
xKxLlllJAJUPC9vobMA4RSE4sbVvzJy5DUwhS7FfdR3CDysZ/oZarcEa5+QPmI9C
invvna2HZVQfhWs51clO8j+/BPDNsI01XOyJHijkLaboxUYnk7gHtaZtCQmzRwf5
ZFBYQVoG1J3+tjA992xNe3+0SPwGj3QHe5tMjuipqhYOQ/GsfFwZ5T91f5Ekifzl
Jc7ItE5r12P+6bOeKtbcLS77IJ8uR2z2J8wvpe0o6MT+cUUqH/XKQ/M1AxLsYhco
Dez3qnJQPA+mjn6BHB7qTbPVOf0soDttDRhk/xlVCT+M5DoGJi8fHAovvz97ZfBB
ZJo37Z3UT3pzgZklYHZk9m315AKkZ8tLtjmCdJH4Jx13fZ1yXlusPpTYT/NTYAmj
NDPlsKzR2M0+DoSUVpMmBJ6h1xJ0wIK7NQmrrdIw38QVqYIAEpfBZuyYCZFTb/at
UUDe19lZPH83C8GYfU1kbDAdVf4isYuMaPMUXieVWH83HGuKy6MlgI3rYMBoxtqr
SIPn4Z8VSl4LvyR1TpM0M3lRTrJ/2RlFqQQO+gWU12l1eMN4nKYy/Jidd39xxNBR
jKxHN9WGS27L3xxa3c/tKi+j45CJv1SyI5oe+GOclEcwPSTogLqy7HmKxpGQX4bS
OlHUiNlhUP/jD/ffyz7LCTMFXZ2vWh3yN0pPB8lVGh5kKdi+vnHuSL+gV2BplYIa
bA/pvW24FRP0uTgQr7OOl7HgiLP7VHxWdMjqG6ZdWRpIZjzrGy7DEa4SLaX4sQxX
jndShDWpk0+wHbiCrMekG8wAxJWlr7T5QtcAYgfNvUwhUNmSENd5F4jjkG3MTZPd
34nrEv4/1TL7GiDdrliQDPZt2siD56bxFlViFCRMZCeiEU0vYH+e3PxGf4H6I33i
9Ei1j5C527w/zO83fiTNuezTXl2663tsUYnnhFN5rSq5GHHmKtyp/nHATWQ+GcHA
OuTmCIBFj3acyqJ7qR1lre5u7I+R+nQcXDGM9bb8rknMgFsXBdhNx+Vy/If89PtM
U+TmVmYGKYPg2ZyRiTRPaoI+qLZGhSq6nDMvayT5Jf68f8BKKDxc8sqovJsG0WtO
AdBsiUHUaC0R5DYzRZftKX22C4rxqVGGrKazmGnh1OCo+BQNm2u8zslO68qaV7AF
Oo8qy0jo0pvoDx6dzDjycPuhK29x+lpoAV848UxzkI9nDWPl2HuayzR1sjXvPDFb
6OdaMmM3z8OVHhemMB+CqiqWmazUUuqMoDx2B0LTlrpNESnGSHB/GHzlTf0N31/R
AKP1mdsQKRGCwwv05HGxzhaIiJIj4FOGMfJ1TRpXWVhBR4bqva/E/B8NDWe8aRql
ONRqFDhVGkFaaa1dy7siBtfXW8XMGjjCsgy+Ji98du9lmSFfwyYYnwHfHPpfp/3n
BEhnnOJbd1V5TkluigUkaIkeQTFt/Hid7A2KnoPlH18Q3AGbIJNWSFljRA1wCyxU
EhqF+mvelrc/Tky2GVDH1P8m6Kzj3rQfGWvvJ21oaj4S9mWRm6xjzBld2UHlRISs
9yyIlqO6TC8q3yscbcDvgBmEhtn5pEEcj5G31eTGpk6ef9K4LQXDXUUiEay4saYX
ke4V9weZHk/e2Xf1cDkYtQTPA0hp0MU2UwnCDDStps+Ex2ZmcjWef/2v/VQvnAz4
WSnjJkjD2UOYQQfD/m6pwYhx+14qYiXoCkVilJ4HQV/SDVRSeHeFi1XcT6Tuyfc4
GUVAprK+GaB9GAGHvoLwLaXp+oZffGf9UXb4K8IAE65aM3wJjMbQ5q6SbfatlmAk
Y/cEX1HBQVYl0AWeILiJ1mvbC9XSdOTgm5SwY0r5lLKjhf32ym24OrIXYKARC2sF
9F/b5kR+m3F5Ncxwlos71F7r+e+IgsAHuSHNcPdACEf+c1HIsr6+GMXgaOt93bj4
ULHl/boje5qaiZBGI8OGz0jSK25LCpCYxjvq8ta7MSceyF+HuldUaLeDPpQeyq2X
uzpMIOk1N3zGyE2x0Yy+rlIgNohzDVPluhzAjRzbIeFEgwHkU36FZ5JldgRDgFRy
6bgKP2QfBKf7ARN3qVGdUb94+l8tv3sDhG04FwhJz9AmZLWJqOwd9YqMpTbf/cIy
nq69OPwQmNZHwvZw2DPILF0GbsM66Lhn2ejGx+xHExdF+yTazEBo/OLHMltlSxrL
370Qp3t6fn5aO056WMvC0VY6iz7FGeioxZLXEmwkJUU1XxdNn2I/T8sYpKMYCsbm
xlWUazi1aETcwp+PxR6VikhYMLdOE4vIbSrc3yABOh0OYFKwMuTpuV3+clsDnqFA
022bVRtJi8XjlzCGMFfNE7CE7Y3VHuvUaf5FngDBJj9rQ6/pWNBCWbhfr6obd/92
eujkPSY738f9h3YA8Qs6YwFaCMpspUsZOQ6qZOrFLQaEmp2UxkGFyVoNWcwD5t8n
QZc8Ef9FobEIWiCaOg/k3NmxEjoc324cBhvx3tzJLXopKWIdtjvOic9CKhPcOpqc
mh0TrASlJ8M1soiPqS8WI7FqM8lNgRsolFh3Fl1w1F9GnMfrKVZGBUGunf0dhAZV
VCOxDQXx1OKNMG14DoGNJ2tn3Z4YRWhYx26AfbA4aVzhULd13hojkP3TO+1+Aca+
XmYKL2Ee+AikC8gZMEkFfpphrb/0N8vo0iPRhtlfAs/omJZriH2oq9m5kZmqHxmI
fFd8kA2UjmXVjxevYoBvn8+abNcwdVEH1g9wbqHq63Cj3du2vgYfbz50r3/BL68g
WNIWxi+SqCaKQZf8+9KgRnw2F8prEDa3M7ZCl89Y77OIF2l2tyldf755x0fkFgWR
H+JF8iYLWoQsgd9kdOu/j0BOpUBMAltZOuhOsGM3dGJTcF0iwHV95stquIWypANS
/K9CYm+WE63RmvMh5W9axA20P8arZHMjxvZvddaVc7TlUzuijG36f70SYhqAosRK
nCIfjLZaxs/39KCaL5igx8IfW0dcNuG/f3V6nFpJB4K0yBNeQpdb4nUxBejT8Mt/
TjT7bwsc6WC5fsfY3yMPsgCh/76V0JpOroL9SSK7KegkZHnrV9PwjTW7r0S7OR1x
dGTx8yirl6ih7HKXISFTbHsdvhV5tnhW0uLbgr2EQ3/Q1wudklR18H5SPU6UgmLr
oMXDjdMxxZs0t4ORmY6Qu+ZVvKjScvgJkSBro1WPPDkLmSlVEQDku35VMKPmuBql
XQBn8pM70ARPMvBK8Y8UA8RIOsqvEpz9iXgHdGje2GZfsqoUhvPOeTjuuxXSPfUf
vvbDDryQw+df09/tlqr/35bQnfNWZ1b4rzC9bbrXCYAFwJhv1y3QN9SKcriTYvD7
V28HN/t26Kaxg4yZkmtpiSCwr0LthH58jG4RJrhUfjI/Hte7vqGz1X6U7aJRO5p1
vRK4qJGStcL7C5dSBcA/LHa4mucHD+SQyj3CWRqwHHY/D4OgEsf5tirtOO5vRdTv
wmiyTcd1mXHr84uGUojhuu7gt58XMtHVGcsSd4kXEv5Awemx6hJ23r6C9jy/qTRL
9EkUT4MAq+VqgO8Z2/7cgqbmcUlmS0gPt/viWKguP7Ny1+K4uYUAjCOsLErluwSM
X7Y+8EuJInnV2ejB03nvfkosTedZ3+mMxPGi99MTcjiDwV7vdoj2pyY7LehSbo4c
DYzf6miJwZEE+Z6T4O+ZPajLnx2qdDRHfeAQRbJSb3hHDpVA2zUUkFzdVUbMc9js
eKqWJ0Q7rq+cECCTQhdhfBZRxJrMWbgfGARFQQBZbdxNzaEmLY34C18p+VMqI5x5
SN7ODQ4yMdPhW14gPPywFUl1jPIPLfcYzzVNyS0U5MRIHrEtmFYSEg/SDm2ymmM7
PRDWq0kxOsOeMYnoeymF2skdHdg58t3ZdIQqma6nsZ/Wp08ns88zpjrB6+3M/BZY
6+bzgJX4f3zIFXILDAz+FBXblV3ZbtZf2T1qWzZFKvv3as1Vlc5oVK7/DMm+sT8V
ANxLP9i6W/MhO4BaDB7VrDopyYYrlE9lrGF8An9YzbYJ7JTSN+kQ/9Zf+kMkbqWE
w2JE4GzJ0YalUPQBAaJ4czn23yZMHGSD2BSzxb3agZt3B7+SQDB3z/Beq9S3garK
9tFv91MRAHRJIvVsc7fWdeUPd1OEZcXl3ZWhHHdXLk2EDyEick+zHWtxZKM1+Lid
rJ5SYKPy7O5MV0YqqKGvoOCkqa+JwNSezxLbrPPXpsXPZgMHWkPEDEHrn2nh8tLe
dtK2stvo4u+Sl03f7mVHFw/QL9dbfs2OI8urYU7Ucq9GrHoeXwW9+n7C8e1fp/o/
Fv0X2Y7gqSjzpkQ0LmP/nDeS7Tp4msXHr1MS+P9COk9kVbGQ+yAskml2KpMQfVSs
HxYinKMHKCIQunJKZWK0I2w0CCEGDj3zeQmq5YIjOJLqUQiHPHBpwseuTqycHfNZ
hW73OV+PVG+SyVrvMXOqYGf4dBSRLxJMvF4miMrjMW1+GHmTeL/4W4BcnhXSlQQz
107wkZwyM1f/uURt5kNxbNvSCTyCDm8B89O6DrXZjqY5eihN9PuXUFSFR86a+9oP
YV7opt88QfYV7MZf4qclBKAGmzOfIW4qk8K/E79fsq3E+QFuQf4EEXLBasca0L1k
En0ldbaYIXUBbzaT6wYWj32pC1hFGbsXDBSfe5aL+X3zLvyRqjsglfEIfmbv1DdU
vOFyK+OIcwEwrWbVQPD2p8sZbt4oCozew6gOhlMFYo5cKi84iU2sOLvk/LVA9aJt
bTGfw8Kdgq6Mk8ChMFAgrNsYqcmBTfEaFoTylKBj0Jz58D8Lr4sqsROgZwGo1b3s
7iHzUX7MPUvIT3NbgS68ROGQzDTPIeIKUA5EZ38yVM0rXsQ8kLPB8o1kKRwV1FxP
qS5PtXqxQbHvJugoV2gqn/GViJsUbCqNqGCO/2IXk0bp6o+NfIYdZ9MWNkb9xGNr
VloiR9S3QbGyaF/zxATUw0aLnjt9vh7u3OrnacK7r46Pcq8kx8Q1KzLrXRdmeW3o
af28gjue5opbfEfgF7ieFU2sy3xtphJiZ01TUk8jzUVBvmyN7SxCSoRKwokb810y
jD3dQPlcrpEVsCXhzRtkAO4G7GTl2ob7GZzpXqBe5CLVci5qB3fw4owYDgYum8mt
aOdJM4tIwK0yFWFVis17VKTRk1CaAaCil3izYz91QuhB1Qil4LtTLakranprEdeF
H8CTOy3kVWbgZw+8u6l9txTwxikizPjF07oecGI/pfwRn+VDBZ+vSjrirjMigdNJ
+bb4bVruvSL4B9uvNOiQ1beA/BWQiWKgAyzVypaxrVmgSPfEHPkTy8bI15TFF04m
dMrfq35j2qFe4v19EvZPr7HAdhEGpl6pFUlpTb2KpPjIVD4XvChS6Fm3m9skafF+
tYVRqCwmUO4QuPaKRQWsJ/8t2knxUrSH70jl63tNfLW7Xp/pFH1+/+gu0A97LiV4
RwsdRCgMV5KpinZVkhVfWCSbhKpLE2rGjccVRdM5nBs6/UnQWFloZ0LCIdMYcTMA
SbMwHskxN0LTp72rr3+f5YvHforYD6MfyKTWXV/55eF5BDBV84mBWnAGXYjMb00j
OIRep7zWGr+2mgjrBr8N7f5gR8stEMofLl3LDiatada8ccTut7aPXQHhrUVepxch
8ScurMxmTa6a7kUDmQSZaU7ioz426kORnteo5/IhqY4PD3Ih7qE4heV0zMbjinrs
go6V8FV1swVK8/1nLrpiKtUseQFpBhGHW1jswmNDEqIpR8gP3WROALJnmLfM1pkl
07yYgVVPoJJuO/yifMXmKOsxIb8gCaDyaben+v4qV9k5nM4GSUQgUbyVw2dobaYn
CBxlWVvX1O+6PMFTnO19AQh2rRJ/ovRcr/8lLybIjuotPMBG8aRfN2zuilsK+bNv
8bB2gbB6KREjdDcD3p40B99HDMtwMbA5PQzmZ1QJGUyg9+HaopvJi4U3xqdst7ft
SiAllOjo72WendA80wP1Ei7wuKwquVLKTXcYyfnUgJoodtRdSTD8rEhAvSy+o+DT
GSlZq5d9mOaYY8QcwZLOnQtDDg2o55Cvee0tkgaJhlvrQuPnnbK1GXnDY7ZOG7L4
6nZIJLyIADVN8h1Hr6tlfBRwCpgikZfUXAswQTjJ3AFD8+00ywqRefoobQmVXo5s
3cmGhGMdgfDDzErAkDh2v7ROSD0QF3c5x424FmEzCLd0xzWPMtsLwQS3ndfhqsRs
SI4BQJsjYjmJysKZnt4eZiMkN8NqdrUAqFTrzqWbzqcFsdeiQMRxEX1RfnM0Zr9e
T6N8eTVHQWq/G98E/eOweoDMX0VEJYHq4j4iJhomR9T3IuzuMM7nhOW698KouGVS
ajehqKxUyMkxm+Z6IwSLCMkyLmpCYHdGvlsw0vQ+xC/584fXSWKel0bWNo2Tinys
69VAGFxIMHPrYEVCBku4/FV54/KVgigev8oILU5EIGi/rzGPFHSD7M3j5VbxPPaI
AbVZP5qRU1LN5qA9/muS9MB7a12wh5IBjlMoYa6xvKYqk+JqN4bWTcPpeZW76CNW
L8guUD1MSuo8XHU8SzUOpiL0Mry6NXEF+stGjrwf3ZBa/Nw6K1A57RiRrv2L2A+j
KnF+LziTzAj4x60FGSKTKsdXAVDeldDaMjIS67a7ikKLWI4E8zKjtQH63bqwiUbw
Imj8HQv438CwKyd+DY59iS09pI0eDUrsLj2gJ/hVKGE6JwrDV4Zs0DNacZc8kOLZ
HzKuJBwgPKsabYUeW9JTXQlXyuTeCXyCxnAf5bUrFYmInrcXiL8l9QbOp331i85f
L9TbXb1rVZkjvewIDeKX1FGuHc2de4jnnlYQmbd1LC3dabyAs003gSZilUJbiOUy
alo3zuV2PvzJdnKOsBCw+3EulxGwk/yaaRZJ1gGaXQ9/dFXn/6r2NTjt2Be3tszu
Dc9M/K3eDkOD4Ay4ZYk9L8zRwiLb+HSlRIIG7Q+5XoGKBB/+pi68ohrE9o38BYfJ
uIWTmfghtpPKrugNyiI3sfNx1YxGANhXqCInH1ObAwfQQBlGjT9l8KF4YlN2pYRG
PYjLzdx8XLdQEZDIYLXRTp/0a8bPKEPyRwOHu1OjWV+S8mH53FiwTyNY0fgKveus
+iOT3j8//ScYrQ4Bmt3alkFOqbLDZ69OgUDVca31QRZF0uQ57/trhaN0OjM2dy9x
RVB27dR1xRR9z8Yif6kyVF4V6Ixu2M/Yhw5tAcLmu2lpdqs6TjfyCBmFvaoNsXXG
f2AW4mqdG57p7H2KYHxTPF+HQUSUZ2KorOCpp1So890Cg7XW6XIs5zb4P7bsdtxC
l/SozebkI1cBXu6RDmpLgOgYlcYkpLPQgDeyWrJkZ94w36SuRX7+bApqw7vPYPgF
06hTmA4ehpD/SBJxGpi9CQmQf0Swb9YGASHzNR+6FbEpfkAh2IdHAMv9Ve+8wzoV
IFm9LTkWcQ9ktEa5TbumoXOoBDixM8gtkVsegbUZZS18wuzG+DQZhCf98NzdhynK
2hcnvtbV3sQUmurlzKWF4pMMJXAE3jrZfsVFLfjQQ/FtJyMP5wHl3xl0LOgjWVS1
Z1dLkf56gV0cIt1I1f1w0/ypvbDwlP/ODkOx3ESZAAKviIoypKvlRj39tsrKZ4sR
15ysyCqNpaBHHuYuOyDk3FjcgjmmyjsDthL5ZrpNsSamuRyca+cTVfE75/HvVf31
LNrK8lDQLnOJ0Fi4y2usO0Z2b3QbvgAsro9x7Upep/vaBDhlo9PGORxRQy97dpVp
oOxU+csf8K0LBWfvpXRcWlLP522BaQj6i3hCbawa3cZkb5B2B/nkdZfJKPzu3vdH
Ze4WBVwhGXBR5unIPcqyStFqVh0ve0/cxHrKCC4+beCSfGig6AZPD7qFTtJAU3TA
a5iFJdsDyFbEYv/2KEQGOXG/bDda77Z+fC4Tlipv8a28qvgwsU7IrS/VunXX9sT+
kBYV9EkpKQLNHJI+eQr+5wqhrk3SpPTEB7HVgnP0ejDyz84XbWNQYq2S+n8NUsum
X4uKzvsvp1PVMH5qxOngVE29KDJXfm96QLOssTV0fbSKwnN5vjxqTp6zUu6w/TF8
8A5oELZh3Oe8cp7eEd4kEahmxmk4nz0A0JZb2V0UFXZi6xN9V7KkrQe+MT7g1Xeb
Sxjh38tjlmbnQQfKmgGT+9qPtAv9xaV1XI5ZrwDppp9AL2vnpQ742EIGfzkyMFNE
RhVfljC6mqXBjFSpWBdT5osNBbrS2axsiZTJJFSc7y8D+zUsTUwGRnJ7xbZTe57Y
xZ8Fr6fjCmPqpj8JDvCH2Vmu2Wx7cGsNwRtCudor/wySYV8JBCDObwHk2BjiN+pN
SYWrE6naMLGRoGyHoVf2uDE+JiLS55HIl+vJArRxJq5M6vGBt/GyMqYTsHHefl5E
TlPTgETwOw3chlgZptmczVo+2Lwv19Iae507gpyPA2JcQSYyNI383aQGzsZsYeOr
6eRSWL7cMUh7ja++uMLTXKWN9GxCZYF1aP7OdF8F3Jmah6I12GHTTNcfhMImi6Ec
sTgt/ApMjYa+GRGBWl/lkwavKdy6NXSZK1wPU1Ir1YvIarGF0W7DC+djsC5zRFnJ
GdZgHxIXs5QGdyrKdjY7TyPST5AUxyUjvhM/oOtes8VNsG0cJBn/2M/1+oM3kFUU
MmwAmeR4tgp6CpDZKp78itCmu4v5Nkmow4ZRPqw2fqmQ3s33GZOWN0vmuD+3m9bL
ME+bBf3nXreUp+tSgBdp95ZIc4PaaZbl/SnwoBcyGA8K8Gnrxvc3eLbxXnuld+6J
9NpUNLDY4Sk2NTr14AoLOyG47Y+5n3t9sFXLbJxJ9dOqI4O1yr6Fq8s/Pddn/Qgl
7jaf68Jpi5u+jXGJ7riRwtPNQ6E9ndJ06gBlw3R2uLREC1wJz9JnUDS8QKMisuZj
KzQ+xoARHzx0Oq7Makw2q3Y2HckrdBRsbXtxPW5eIz7Yygj7mE7ash1OOFYQGaD1
Ocubq+2g0T3LX9U8x/wlG3ubSW9axu8Pnea0IzNHOhKxZGMpO80cAYWXaevY4csY
Z4dHFuNKw9lHF17LnEG55yO1mlrIV8hxqGGZKL0kVJc6twBMyUezI9PofAFVyZBE
IfNkRq9ufoL1VMAOXTNMKrFxytaexQcaf4Y7hClc3n4Zku2u/ILOSb2V5aA4o2qr
CCn6f3mARfVn9r8Zg4UG+UOXw0zsR1edb/iNTANMSW2arYrGZY78SeqlaRs86Z7F
yfIbBe/6WYMZ1DLcqo1zlo1+d1Ozmrc5d+QMbzJxFZH6DPDkyD1Y1Iqy+kxlUimj
5/ABsU1++CzWhRwq8go1GbmQfODJWV8w+rqcI6AXFcI1L33ZlzJmoRe/fTASZ9SJ
USeL1JyFxpVz+2z/RqjhR6TnYpRGVgcrxcRJoQr0fsEDb+wYKkHPMX9dROD4J5RE
44qdaMk2J0PFGvW/T0qqRbH0EhRbwyTOB2zusqMdvV8fNB10xevPfrKzmYa2EWeb
bCB3f5hEmGWVAwnGJfUS624NdcbrhRpDQHKyhMGuPdlhhQWre1AzsDLl3//rpqgL
P+2xFjq2hixUV/ycuo0HBm/rIN0S82vbRz/mfAaZVh8bb5QUAbpxxhRGDSqWZRqC
jEDAoMcTz+0eDnBpSjdcbafYoVJeEm5+PwCzotSflZYhjNJnk3pRmOW4Cqp1XhS0
K/VyEsl1MpmnEeiVu8ZXll2XCYQLZxJDJqg4tA3ttA5kWBseKbwY3IgG5TfOrpTg
7LOw5AIm8vAkATjTzioq92g9Dtl9HciEp986X3MQhNHm44GwIAB/eZ/YIcyuJepI
k31yX6SXl8EoUJKZgisKZwZ9j/MNysNSma5tmbq29R61g7C06EMZ6uBbW012SNMu
SdulJGts7wav3LBbDazmiRttrRqYiLP+DgBI7mhN9XkmidUDiXnLPZHjOX1zSJXS
oVe+oY0YLdDnsnsixR6c2btsSpmQHpTK5aJIuxlLPVlNt4vZo4ql7XewpbysclT2
9rC/XXZjgFIA9cJW+zt0amLbCznm0DLrxZMVKC8QQ3tMagCB9PyQWQ5OZPnbiTWL
9EIgPzqEKXTW5WfwMyVlz/FYWCDulhkKB+2MFGmDQexxMS6RzGnAPtE8YtBA1p5i
mEYAt8w/+eH+x8YizWkOcsYCh/iAh3rnV/A2XiVRX9CxMKdKAHS2MlO9UcOTylJ1
dv1MBjZLZeafOgPR3d/GtineGnw9fWbIQT+UA2NSPRxvmvsgbyvjOENECOuZ7FZs
JyiY5adQa2N/rKOP3yWKNIuNe+bPEnI5Dcd951QlSu7fL34BuqQ+Y8buVu9T7kEP
Rhwjqe7ejHsd49/kWwMkvIGY5XruYurQi59Rz1HlM2i72HM9/vCN3Rrf0Qj+Et0k
IZCk+d5FPLiuxdKxTdry6C7Jl+1N2hjO8u3Hy2lb1cfHMKAUi/6juqYzqerthFef
D8u6Nq4oHjkkKVCWBgwed+AaRPZ0zl0rIo07hEtbZghGgQ6Z1cns/cBfnNvWcXTY
P3FXMdt3qOmiEY8lHhZ/iESYTp4bQu0MNckVsNhN97KloHUgymLmwTzzWOWYIYu+
/aGBO1Vd/G0ibVlQRcCnGYY4cYY0IPHpc80Sn33ppmVPzkgN1CnR5usj1QxRSJ9e
I2AJPXa7rYx3Hs/EgamauleiR9EmwM6hj/YSbxPpt5aVIcc2YlLW8ZGXhptmrcwE
7lJg5B8gSbYhXFPE96PH0iPJdoPlJnKg59sNH88TQ0v4auCLJW/c3g4urCE6pRmk
5een20xEMxr9FeOyAN6u14VtDcQwFVLyRuQM1gn6Leucai2Xqe4Iu7besEqWQZrn
SL0mYf1G8sVpyYuHSy5lNAcXTV2I8uAPoltbAb/z+Nz9UL8c1ncN+Xbyl+jleta7
EKXaIHaeA1ZU4U8qUvfOQ94V8rk385DUdGCE0SyTNbEm/I2cjgdICTykrD1T21JN
x0yc+hy9fkKMrHMHNmI4YEPg+sS1mRmlbvmoqK1CE2WEfKe8URzWHMVwFaBqaw92
DMKEituMuPFerdogEuUV8xVcXcQ+qJjLDv3fwnZpBlSjp1I2cuGn3imEliO308Bk
jsUWIQ9ivKc5pwsH/tGAF6y/fTq9/c/02AK05RcNF2V+qGahG82JkKHF4etQdDOT
rayOifpe8jqs0IImXu1zHwn+7ygTk5zrK85S3b2G40dzQWLw+AL+rPx4uFPIyf+Z
ViO/Gh7nl3PP2kIA50snVpI6lQBVeg3h6Ct5nykxRGUe9MmVAch4qIpcDydRT3TK
cYbqxszfUL3xSgDCnR0jJVbaiSwwAH6lvm0rG0Ej5PKrmvmMLeVt7nTUl3dom+Ev
1KW4y+VcYJjJri5tupCKCHyxTUZjLfqt1wXxAHmUyKh3CJR+S08E6iXTMeIq625B
FagVRvX3RK1FNgmzXC/Ese9Ny0qVBh02ZQzgO7HMSY0tPEOkaAAJxI+eL0BYYcuu
SNdZtANeE0mn5/oY3LfGUPn5yOUAiFXkZ9QBHv6H2BxZePYwqI0dOM+3wqw+Fohy
0aWM05Yk/rpAL5lASsVewAekbmKU6qlrjd1vjvt3CRVrfiBSXXl0pAzCEImMRrCb
siFMcOWvj/uvv0HU5yQk24FXlKOxgTgs1qcp75RtzGG1gAPweUbnHX4dhxhrZPAr
ujg5yE9C4AokHc+xE6ehCfDhgeSP8omHNIs6yt++MU2dsUFuKV2YBr468WQlM2WD
LW05kFnXK6uAjOXTe+iAqCre/OkGYMwuezJjeRB+NOO53/2GnqRgJLQO+gP6C5sU
GI/UYzinBu/PEvupsxoixYc+CBfqZFrgsCo5bT0PrP+vtqZyduTkKHMYKQ7dDazw
BVNr+zPCgiI6xZhZ+JM1nf6C0JwM28Twc3Dtoo29eVuiaPlkJctQKT2/1i/jUBxU
k9tXwbzvXEFye5113VPoIzVCGzgkQkuSAi6gO3GiL4lsZRn/pIdmc1luvImm4WfX
evKMwXAE6np8cXmq7O8MHshER4aAKsYvPW2IRX3P/LeXM9i+zrFC0cOHGWQDksRL
NzNBTiizaSjSxe54YTcjwCclPZ/5R/vddSTj0kJw9KZSs/AYKxFySXCZYcUCVNZs
Yc0KEECI8CVgodf2FUl4JYqN9bAiq8VrcRqf/Jh0fySVoUCb8MT8zgzx1RmFfrQV
orepaaSeQ+ncA/BTq2EefMLQjEKiEP2dCfnfkG6Z/r15QuyAVC/H/rpTyZIKwR2m
btYXaDcv2+kC1gyoMPkK6RLIvaVIcK3VEWhEBpdI7t63JlMl1z3AVkRM1soZYEvf
zpoZ/bg2EKNRXw8ENCwIwWSafqGf6IJqPW/sxrXVvRA5R9qhBpU7EOMYTQzb/BZW
COaT/KoK+ZYY0DT5QO2xCHJf/XQwIcl7jfbItELYkf6PHWn5FmX3BuYd81xb4vPz
+z7ygX8l0BVZfBEsKge6KUEcbSb5/QJ0ApnvARgy0VU7wmR8o+Pl4j0cHI8bl/Ac
PkwTxTB2SBdzQ9ENd5mN3n0W/nwnOcz7CnfSR7Q9RmZlYjYWwCi7wRMBUuJIIuyq
VEcFI3XMaFVdNqU/527YCJgYl6dfmLWAxOc2871IEOmi8oZTrDg2cyNTTX16PMB+
TIzFv9QZEMBbcPm0xfGBQ6z85vdLi4jFenhDnamj04TETKKUasheBrEGlt2623qY
akc9eiaAVuD265YCHNtw199531cA+vC/AMsmcTgap82qDyOws9PSuY1VjbbITgfq
FeCH+456dvOYoYSJAdUI3n7kir3GbVOwzk8W+CTbv4uFNS/WnEu1WiEzIEfq2mxG
/SVHSAwsKWJUFcL1hpnVCs/JIWHwKaH988qdxyw6GssEwso+YC7CLvPHQGcs5AW6
Qf3b+glO4PA8Qwy0L2s9Vq6WVa8BUxJlDmTwZKWlDCJaJf9Qrhm3TiSynQSsjUPk
7KBSS1JzvLr/VsG/fztO5FdvdElXkzSE5uhWj9QsCxa2A3BqINdFnhSV707ONn8a
nz+y1Xo+LOsxgnkYFrI60u+ZLinqbILg74iM/YznxDCSvhg7QlinwwqB62gloNkk
Rx0Lo6Anzr5h1fCKm/ST7i/pzTtg0n7wpB7lPCrdUAmOro3ppsaRDVFyd1kcZt4r
zxpvb92QA9Ul2hMXwiWh/c5lvi04H/n2Hxwl8LLa9/+RXGAcky7BGtQYfqNQtfDg
N6vcCbDnXHLLwQ8MA5PNmMOJedgFFhBPIvO5ONGy1UTtSGDk4DHp51m7vn8H73fQ
5qbbO55Wljqg8nVyYrhaRjRCLwmBBODGB91+QrHbHyb/wCam6LVZ9R7OrPJiUN3b
Rl5LwYXaWHniuwo4DtqdKorDprlNSTMshFlCZULM2BFLQw7/uTjvUuH8jbz5RdWJ
f3IFQGkKUOkNHwXG7lQqlLHZ1vbV5OV0t4etD6hL5/F9yH2SZRJ72GcvDhBVG3bI
UEAM+tvPPDJgOk4mhnYMnDXDJuUmJfO8afW00HTc7/58zCJYvMP3Rg0xcS/yQp6+
NFn4ewGnzeKMD3eduTha4v5DTjUNaSh8TIYvJLK+qKfn8oUVEZWZC8t49xp72aif
6zMph8IeFjeZChwv9nwDUP3qjV6QIq7r/ioCkVioiegXmcXWf7qtyowg/+WrTeBe
ubn/FJnTSPnKwucfBMsUQFshnTqdk9DW41oshQ4qNlkYju5FWO+iuNW74qvrQ0Lj
Z0gsy4pjvmHAliRCG15c2Iyqj5mFc87LzhlFNjEvrse1r6vThP+at9R/c08ZD1fl
90HswtqnRMGenqonVvAwphXU+4BqhZXDFkiZbU63WSpOnCB4GTRmIPoWeHo9Lbap
EBcZn50CphHtrF8u71ql+uEEErly6sHZHybDqd1K3BFT9H5btspopR7W4EgsbpX1
GHsiDoDoC3ANQnu4SCI3uzffxynJWy8Ewmj2d/sxs8n/3Z2QMs+7nIVHyuRVuHwI
G4HiwwZmdX1H5tOPY3ak8egLXFGGozwgUW6pg8GTeuBDBPm8mkg9F7UpyLHwvRYN
t/3hJ+Z7kAZr5CahyCcL6ZpdJ2YuCmgd4mMnhGosUlV+DGBOkCY3mPgDqBqn1iaB
JyGMlatTtwG8m/sIYMChj10VG4+ZveehcJQEiFfTB9tpBQr5bkyycNWFWRQt5Il1
BBFmGU1q2ulZ6/1Beg79rk1Q7jwA0JrGSrNcDog/woD4yMv1ey/IiKv48Qz18BiD
dmNzYt4uzwGiixdNhh1IJiadHoSHgv0MneG2V4NqVxbU2MJzCBb78csOMpys/Ccy
/K4IcU75qObPO7XZKJnZXMl1nEyliCAeRE06HcMQK+OHTl5ETe36NpbrSuqL7Msk
2Kb15Ln4VsCg4wBZuM+GU3CAjnY46PhF956ehVuG9lHzqWLHx7dBAQK60ejoVaQR
F4WduymF+fjyahGx79Magp6fzqYzh14K0cEMrV0g5wsdZUHxqCEvJCtI6djVocYu
gB3sO9O78WETNmVOYIx47Myl6RkuRU5XaG9vTq28zEBnAvVWt+P7r4YbkGo5kySY
+0cdc3++P2B3FcCHBuyjHwY0XCpQSu90ze4SMzBSU8cyu3BEqhNrAohV1lECrVWT
bLIam1Fxfoi/tuniP6CqbBbvc9jo9EY20NhzZCfIYTJS8MdQsyJG0r0hNy2zw5cW
Rjk6N/0hj6440pgZMeEy0qSw0B3MZPrjMDHRw28jkhh0FiO95e305OM/68WqpyQF
jv9PGwqzKEFA14XGCnLMtHekjlgnABFjksGzWRWGPk9FRlZt2CA0cEKB6Wmy2uSl
9hHfynbg6TF15Eizo+WFX4Up8VnTQSCxE4s9JeHFwdEWAGJnMiTmSYkuZ5P8gyY8
RLtnpGmItXlsG/aB6jQWIUuL9aGegl9vaqMNuJiqQ3p6BdPe93C/HAmzz0CiZ4eB
506o1u0SH8B46vThYj0gshTYVPloLcKnicDtU2GwprocrSjsFufTl+z7QJD/mNaP
tztpegh/FdsKCAkfn9xtxaOQKTcXvVLBLDjETaFFM2BXKsRKio/uqLf8Kza/axlx
79HcsGPQRX25K2jU9C/KaPnrS3cq+yojs196jmg6rEX1qFkL4/6syzDMYxFtq2uL
qu7IECLXkyO4v9jm8TJ8C8q0iIxegVqqFmYM1uLYGR+wUYpDjgjU7lgU100eU55J
9zucehgFW1wmZoxM/HMMbQHftJcTv+serkDp+w9Vqn8EDT+fhGk2JLsdVu0a4/Mn
toROFL2dcuMsJAzvaNcRw0/JFvSnAuaZ1eI15nrwdgv97JRvqEsXWEhcM09rcbS5
B5iaLKR7k0Rcozl2Sx5Czhkwp+YHIuNEAPKSoIR2e9TWu4WH9/D4wuCApTHWWsnh
EpoYwk4yaITKsaLZWFe/2JYOUZRTc3DgEfiFVsJYaTkYGmttM7QtyFIa14amDAow
xO35GEeB/kkoI9axWQwyvvNFfXVVltQJSTItuJewfE73A9EqRhWOFZU10j6G9q5Z
6FHRWooyWcJt3Xq/d9hYkL50ksKk7u4bcEQ0qNrNu7hzUVe13+XlSNciSqgEkd3/
28+VU3PpXtXAd2fQP2YHgo1ya+U7vNPmkg9s6BNf6gQGn6W2DKSbJRCxfV27mkHs
TefJQZvlE9oovZSVd8i2+CHd2J60TjTFP8dTCaB6avrX+3xi0IZBdy47UnhN6LCD
YiwY3HRafY4EaB9EwPno6YQVJJPfBfCxNI2UaTLGegE1lmTZgHByKhf3yKsnTIbS
f9P/idzRFZ9eaCx9bRsEb2Ccawvn14k3cRU39DGi1Qnd1qEQpnn5K0WBC0DXtJHF
gP/ngI4ZFlY/N/yXL1G9MJfU9V7HaPUZwL7yG3BUF0qelcpYyphFNTny4/HCoEI2
wSZ/w4lA+P6d3Ed6oi1vbFCzmvDqVkmvUC6TiYw42hzDyhTMeNOepIqA/nHhE88r
Fua0SbLfEGZ39eiLHJsekcSTwpdI/BE1XwjZnVGNBjTMIFgX5s03ijVIH1QySAs5
tKFbrT/7hcxwq2GmLRGmPUT9HwzyUvJDsva7WVEmh8PyqCGuJFggyRFL2rlFwTMX
cS0un3OHCiQ34AZ84GWBsHLpMAVdD1kNIwL3caLKEOf3AIJMmdCDf2YfRBevuQM/
khYGfDt/7/Y+YLLrrFgj4H5fbbMzueEdnir6mZwu1DbJfdycyhedhJLheMglemkY
GQ8F4Glksq1l00f7yvjtyW79ubRstlGUIg9o9TGcdkqRzIBQI/OL1rZrhicuIhQQ
K+03IVpYGefQ/+C7DMWddfhkd3umnBf46naToUHVOmgKns4dDLgzsl4mJU2Y6BH/
0bHxyJgr52r+6wD4eF9kaAPx48Jj84DGgZM6HJ9b0++B95EJ2scaZOKsWCfx1GOm
6qjoGeYuVV6yZ3Dk04efkoZgNSQ+1znek/eCX3VgkWNQdl3S+KjqEpe7zD/9Yye8
6C5iEHk6gwGZ6unCzzfTXM+w7YpmmtoTwKZd+mWk/1M/0NqgnZx1iCluiFCi6T0r
pzedeDiFn8okCXy5bw+M9gWtfsRqq6E1hQDIdbOGu0YpMV4Vurns6my+M1en+vbd
5SFDORpJcS2ox1XAsvHF87aGzjX362pPSikQwe+hiKGBEWUQQe9kFtdYMknkDAri
XB1o4p13qSZaaz9WgzwNiHkpK0LooHUknh2q1pj9nbIp4cnNyaRVnDXq/ICMmUAj
JHtMD1YfitbLDWIRdpHYcCZC/mdsmRhZSzbPBPylSm/VKlyeeQC691SeIEthoyF+
nVcSSMn73iVKErIqmFdlIwECVREV5C6i4+bGv6tFqFUVwZtxqK0oY51RjPfVGv+C
gMynQlAv0Xlnc2BHO0XfoZxsRpVcxuUocRCt1OGsDn5pi4e5V2KUqc1eM2DFW+aI
Y1/nmYJWRqfzi0xQoeQonKIEnK9lRyxayKclxCj2Xo7T8CeLCfcwArPMGa80h6mJ
Crx5OcMCV2xJ2t5eWs3eMo9GPQQvjqFfrMR4AHZ10qo5Iv5DU8n7T3HBir1POCeo
JZBXwkl0UC1/qya+Ou2HIEDufrZIz+7KiFrcy6wQW5k85a7P8cBKQkzVig6NyPdB
efLU00hq2lh70O6fMr9oj1Kx1st3riN9MUGrmKl/3nwfkzlhVzfBkNzbeWVoWLeP
+94QeSJqfuajGc3y7iXit+Ivkvwvq8W4qV3GCLTv/57pJ7RVsCd+8lpgM9p6mpb2
ljj99Zb0eUKkPI8QYaHU0OddRfq1wVHBCUFZHRfKF+9bp6dVRAVAeYuqI5kmMi2O
BKc6GMGX3z6hMgLao5ekV/WFyv+AOnyeZLEWqlsiAWkmwDK2wnnt21CME8dANKzQ
bjYfjei1p5dVFNJg2Q9lN0tKT8UFCN+AFPRnLJbdqOx9MIsej7ezc9ZkCg49T0bP
c8SXNhPV3HKrQrBJHANn+nHspEGLA68iA+E1vqoPhKVyNfPFvd2XveVzY8QtPaFU
GiGn0tW7o3NSJFoluKtajKJBlAAXcg0qrn31veQECvEl4ozcOGEBAAw4FGRPtuRA
wb60NyFkN6k5ja7ucD+du4yRtRPRPez4BQuy3bPf4VNX83fnWTP4tH/IN7kapKBg
CX5bqEWbyChAjusm2cJ3TjkCKNG4PMMJUMx2R8GWUcXPD3ydnupsQb9r1AofYkh6
5K/l5/LOznZ8n0tVE8O+JrnNGP+VgFZV1Hr86adU2M4djBItU+h7QGpAOnYCdNv6
CEQsBVNESTrZvF9EshGX/T/V3GYliwQpcl9xV4Orx1fRIr83OxzQLWvFF+zw414S
1zEl1n3DEPuyfMGoyej5JVrksTo7IiwMQLlUXo0f9BayUNuF657R1uUaNn5fAEVN
8bWsXHgGhXgyqIfVcqtHpVvuAUF0kfPDkHtsyive1tQq2rYj086Yv1nzTfKPbT6k
92rvnZN2uQoUAWx03JHkqyVd72Utn/UCJTyN3flYmvOtoAslrIG3qYiQ0/SJ3z/T
nHrZW4Q8i5E5v6/3Smnp8PMwhxJn1Drb4qRcIhOzrlgFf7ty1Uvq69JCSnObSOiJ
tgS6g11JR8Psjra0Yva6MvXN2x+HZcxpQf1WY4wD1V/o3jw9sO9gll5374uPjIAh
+HEnMn2K8sttOpgtNFjA9l6XvhSiQlraboH0iSgPbHztug+tbhRVv3TjG4qvtrPZ
FOqibWh/5hQzFc9TqzeE4U1kUk8IU6kO4zApSktXnUMxXOtxVdGMjgpb4HfyIXUm
9ynl4odMfJuspfSkjwV4GrObct0Odfgt3m+INkvEWYBf3iV64C1T4Z8j8KcJYvAO
abJzIUjhf6XJidqCzbtmIKyMQD9mfpnusnCs5ov+T88JZDAh6BMPyV130T9ZAuKx
xskdftXZXty26mRIH1/h1dKeXGo9m71+XOLuwmjSFXSNjTTcgba2r9zqbxTAmJoK
5bTpWHBqy+EVpvRZaSs/R+77NHigZQDlrvjw3c9E3TeFxwjJjY+o+UxtK6hpc4+b
fx4J6KCcp0CCGN9g5L9eACuxfrbikc0cK8c4wcfT2n0TlxsX+PZSKvaB9GzsdDTQ
dOcT1KGVMURzUyqzwwlq4+CFgVwfhHw6iP2uoiba3LqpGMktXC0ZyHstYWz+xa6/
k+WDy7GQ+itGKaBYHbu8PM9vRQ/oVauxd2ZfnoMQaM4ofPDdXc0cB0YT0lXElR0e
u49O3Dpffkt1uevZP5CPoh2tbWUHO7/+ZoV06/JIN6scu4BeGvlY7iTkgykgxT0T
hwNG/TCYQaEgf1JmqfI6KKHPUXAcHqfg8ETDV3fxH4lNu8KvUPhzA2Yyrksee781
Y0zuLyHw+pLvzpVLDKixjixcTcvKT6rgfi7VhPccGdBc5vQVTjGtqqp9l48mRwhx
yV5dwgqzTkLeKCQaiDSG624vmoWNnZOSyRUNP0PI4x3BsbI+0TgZ8TrEwicIouH6
iMgnEEqQvIvotRV7hLqrotgRkpzSiGAuplwmzeiJE+WRpogtq7pvH8ENzGdYt66x
F0K+fK1xXIFCAyxtcYML5NnS3sjth1BpPeJpqmdY47OhopewGvW2rZ5azU231eHk
j/aCQ29gIv8FPsNbR+MOK1bQQbEbcm/NEkEPtReLCarrw4OaAC1d8msnNYgrTpBE
zyMb6RPNrQLT/BidXzJ1cswXqNCcbLCq0mzKe+lGYR6B6oUmpe490jyrVrUEvy5s
IDywEYkvOsff4DjrVX8wt19CKl3BTzptcqvlVZigclAdN2zaYuOqzgSAOgDT29pE
4SZEMj/otJIGyaRGE7cVVXQiOahGIJnvMdeJS7gZF7kLeasQWb31J5PmycmZxe2P
WbrPDtpQchrCV3gWDwX5awr/XnoF8sYkSBq4d9vqesO+SQkZCu1un2ojGripwnlL
51ccpYYh9bL8twecSVuqqdnBXhvpZAWiNZ2VGCjAqr1pXwlMARr26JaDPwfrK53S
LpMkH8M/WX79pcmjRqHxxGjTNRnIgIc0z6rcH3tfMzO5o92L4Xgcb/JDxhgF9R60
t8QH6qwZRyxgy0PCSrvPLL3qKAI5RtAYZ4QV/4DRw81vafgW5pxunE0/5RVozSWE
LOAvoQTLJ6sxFddd7a6zB9DzaggxFwRxmGbumV78HHXkF28rLtFfMO2lgZPX8OtE
jI17z+nly4JYGOTdVZAWQIPNMf0QWi6TF+5PJfArFJPl/NQSK8+U/QfswMVak4hH
2HMoTGl7/mVuwEM/hXWrWupZK/ioeNIYEdeDBrfmUpJV9migdQ8wutQcVmaXxiF3
7uNbw/VHfzVGvxjVD/JtSF/zv9UQRnw7a9AcYLrPRtzZAfTq6B67bVAjRXeriek3
HVYUGRgVUkbuVMdl3F6BVm/i22cO5u23wZWsBbz9CxV7RdcrGzncnkTXOmBFE7Zf
4a0TroDZQdB7dz7blahGe5hI6Mmxp8i9Xly5W1j6ePST3hdCwY3pnXdlVfeKnfSI
0EEX7Jetk6LOKyg+MDApN6MZEtqubH5XdPXEYSP9ED5+5Xzc0OMoRa+QNSJLb97j
kSyZX9M9NP7XYctZS5GNNWMuR6+ygrEbbtxixqu4kkTzeyIEwwd1dAI/4rE+mUEX
rQZIzBFQAOJcazejifXp7JJDDu+5a/b5wqgr1864l1f/GgSEMUhQRuLXXCd4fPPE
RvLGjjvVnFsjmQihCMvf7McE01SKGOIxiq1Djvuz6vREfdlESwI1taBNXoYVsyVP
lMbZN3LK7IT/xBxt7vagIyydt5E0MBloaLV8oMlV0sgZB4uwfba5LCdnFKWPmQG7
Pjon7Bupa9OSITtU1WiUB2lWyCtNMnLjeiOGMkG6DjOg+OcyumjXAmgKLdzMmCVJ
LA0CUxvPC9PO0PCf40N2SYTPEkIcc+LL4ecoIjgjnccn+9HFbYTnrfqNrGqjGU9+
+VHL2KNEvuOVD56m+hAbVMs2/DthUY/a59cVbOibGbrSCM30TadjbAqaRh4cSLrI
qut+bv9ndV4H6d1OLM5sC1/GhZQAsfyblJa8jsounKnb9+3DYb6kOAHHgaXVM5zf
bCEOoCEI6GPRhAhy7WLpSPlbzHZUruCxHcV+I8apBmYBNWNYOnWZjsqEJLPq5t5t
dXtA7KJkrdjv7CbCU1NVzUjOHQsTBTg/hDhdOfW8jdAJfPaWPxdPDpy1bMgUVpXY
SB/P//Ux3srUts+X6MDeeSBh2/1z1DCRiho9u0jmW+qJKRyHjeSF01HoYyM5EhEe
dIeIRO1BygGv9cv0Z1sbl5dLNN/Bn2+KVeZS2RNglOYrkJzXBAGzfl1RJ4h4qtfy
h1u7TO1O0FsIqi+etS1zHsMShF6kP0kgrawrF9kA+EuiNhpOox+4+0qHK18EFwKC
OwoGZX5QRuVXDkmVmJeqoS4gG4xUKo7xV5rP1uYbBxhTFm0NoddPPN5wJwm1j8Or
QYwtdM+HQT8wVJ6wJ/OSHanYDRUU94xkgvOeya9dnA2EdVUlhMt7CqtF0pndcNys
Tc9ZITWFpyL5tPtz2s5pBXbcUTCT2JIg8C8mk20OJckMrLRE0rlh1tnsfMy2BEBC
kW1QxwAzjqjoHaBEnw2Lhsqw2FdX7QRhCBF5aV695/EU4NSbJ3KMGXCYTiBvOvz3
slY9W9rBdtIplQxGnJIw/nYpe5unbx8I2UCeu2xE0azfd1+cMFXJ4DXQ5DnGMYvo
+9PhIWEMoFBgkSazcDy7cVSu2QmWNc9yxC+OWl3gsL4O+8BQj66HMz8o3HtQxNUt
EHZodWAU+g1I/syKcBkBZhRHx6fin2TdOUsZE4juzvDyFBiP8bc3/5Cc4yZ6Fhm0
vXNHCI855kBdrUBpf05aIVBOpyTvflJ2QQKuZgA/ojLO0moB+WBEIrZf/20DkybS
VHbVUAN2jsH+3rzEPS+V0mv4YnVcl2J4aXQi9nD7Fop3oKX86K95umJ6IGioMUsF
xJlMM7eCR0kn8YimuWytJt4R2UW7D+XML1HHd3284Xeffs8Htm/o2hW2CpMQIxZX
2kCofw2u6mJkwEteBenolOAmiWrZ9aT4UtuIiVRY86GM3xdYW+UHGAtevO0aUSF2
O+aYjXsYr7S1eTJemaHCbAdKiC0BNRppoWq0yaGexorbZ8v00GGn1IfMx58E5Mio
mDu7boLKcC8zTtXV0HoslfX+WBQVFIdsnhA5McoBaUJWZBn9+JP2ZpeX+s53ydb9
ZYSnY8KpME/foCcsZ8n6MCs+UX6h1yAh8nJ2CxrnU4ZUj9n+MA8y8ZtFtda6nzFn
JVPGVVH245u4FK7W9X2BTkJpPI+7U6E0eXA6FKooup5wSEET6bpO+Q7PskISHTU4
cIqMKi+VIhaOtAFqeGgn5eT7AL+c7TZ6jn1XtURAk9BC5G+2W04AyV9eFhfV/kA2
r70rQkN19OXn5Fs92R6hOahZUERVLfNZWIVjtbntpE/PyL184msR+hJtltPuOELC
AH3RymsMBDoOsj93um6IBP8vU/GcWuN/EGZf65xXIVJtj+UyaHRYttyzeRKSfPXa
S/xydotQ6KTY7wIjWndqqG3Iy8ZtX8LA9uVj3B8TQ3zPx7cs9vGE8xoYM/Exz0ul
NcSlUCc0bM9iihHONb/K8j0iW7Bf3PhXzYRifCXG1MFjmcLYpR+Pi48zynPojorz
DCfDZDCouup891js/HXpvp2GTwLeiOcwJ1agMwEKnXXltPifnzeMLbPZPI1qKop+
84or2nhMAApg/i/fGCZqao4KZhR9sxTauFE4tgsanNQnANiBKtIowlVGB8lmxiNW
qWUNBrMnhD/4AwpkM4XbZ2vuAFthrbtxarAfFG8hGuHNyN0C062FgsihZnuTpj50
1K/zZsVn5F8GB77cUHcPnxuCTQLUD8xrlRYdBJA6Ugm6OMFnOFw5uoKz+E89Nniy
Oil64cWaOc/aqjk63ZyBOZmhdTVzZtVLRejiUwWelGARHkw8e9tEcTOWYa01+M4k
vvdeoF0vlU9nElEukeQQfD4ZDHO2EHOU3ms4lh60FJBl+1uil2alCEx9y4cYQyh2
CFLqLXoR2A/9ov6WB2beF73jy4dh2B/zuOynEwdLSeEkEwAavmm05TK0qiCVN5u5
1/Y9bTUoOiAYYRBXJqS8nabdUAFbLfmQybCxJs05F59X8rpGj+UiOjyYvjOv1Hmi
Che3ExC92EP7E7GP8Io22Yhne9IwluvXzQJ1baUUXdwkmlFDcUCkI1zoyShMlM3F
yq2LSbAW0edxZv8LQYHiURCoZBzbLQlNND1gkGvhf8DRBjiR2dfylTNVbv5XUsC6
MzAUFG7AIAbn/+IFJ8zx6vKeLC39zurSdeYAZobI/b5yPg9qKH3vm5oyQVDEOrLw
8ldhRxIlrGCMvlN6473tdg7X8TZMBrjW43zN3KKuhwBozv+APVPlcQiZ1br61YO4
jemIMsADf786Pqp17Gg/Y2T1RZcngLu9CuZaFR0VK+KJwsBV7F5XAwwn250ydUoJ
t8UHyZeR9IvaR6cUps2juXKFxUvga53Lrp7K12/gh2K1ncDH0dYOa5VXxYeKgJt2
7V3b8GF2oi/OBANRFl+Y6d6URY+5aLGQvxAyaVVu2RhRp+uN02rPC2o3Urt7j256
tJLtvj8DF7U2YWLM+yPEcNpTjQCmpHktedF3sNKco7hnhLN+vvjIbIjKyBWAb/4u
FjT5LpBS/DIuuLdgepzWXnlVRfqDeWV6jOwP3St/68hd0esFjadg1P5hVKhPTe8T
U/ao9AQdD7WoC7JApuyiYZjMC5nTLIeRkrkEgJbYLGnGxHM5aBtw5lG00sWFal5z
YqZqDulFg31UIqAMKl1KhWAxHqzyAEbqfnXaHKeYAjzZIau6nwPuN9eWv3V/UOOo
Zl316u4gYkGjHeKqR/vUHCx1Z2pvCrmTd0FNrIamcyS5LR6E93U51dXg/7EDaNBI
XBrisfjdaJ6kXwICdR3RKg08Qz9a5IP4A8T1d2NOmtckooWJHpSUWDeeOsNzHmGj
sHo5tmh5OLg7SMROYllrWWkXw6bi65D8U9n6oc1BcrbYC/tzXl8Svph4XK3VKJqZ
dsPzIONMLktib1HSRaVjhBg3XHpIxQfvTaWe0lTFHCEua72yae/ImcbhgG1/5WHZ
pX/DLpU4LSfis6+NdyBPvjtj6f5OTiIAPlbaIZ26FeWc6++l3mriVtIY1mbuzPLX
L5G8+Zvf/XqI3OfbBNaR2Ue0nCiKeDdBj+A5/7z5nDhWD4XuUAWSX0i4nIAHjkVo
pnSVt1J3NBBIvfWqm4uBT7lJwNLsaHm+Tu0UkZQ7yK4ai97LbwSiUThIbsq0G8sv
SRudzmNd1PNC3ylwcmdy96Zemuy0AaDoZT0/a7COwtMl5AJO9hjoScz0NbC6hOux
97B85Y9Y4HCqV0Ge2qnhtHEWWBOcls3t82fixUZJvGkFjNF7dO1UXtjQKxkb1ZhG
Sj0Y6vwfd59nPAHlKuWVBvIeoj8J89iwfrUkb8JnVxbWKbStrPLJMHMZkgPPFvLE
o8K5MEWLlJZn7s5/Di5UREhzOt35gDpyFfcHGfZ1Tu8RfoG4UEsyuZ94NFYVL63W
fEXozv9NxaDQl6vRCsDklHiElvYN708+mSoFBQrUxQrPnL6mGgpDobkbKhlOiDjP
Z3rwjdOxb6zhUxejqI7GR2LCxsg0dJNH5iPpsA94YYywQ8SaDC177zMALQb/ccdw
bZ/RaGPqHFFOMV6Xr6RuMz+Y5bpRl2LUv9dKY5hS/yiOiouGozj96jI1lIKergrF
vdPRnXkOBEIPUOswskWKy0oSuFt7i+BtkuZj2sfc8vDRrXroGF2z71HVnTN1CATW
scs3L/6mcGgn9YZBtbS/WUyY1LLuTG1LsLGb+6PUAPjuT2bLrTRpDOOS1OLabblQ
7EiWF957CiAPi+XDmQASAIFASB2Kvv3k7agJMTWcmTp1wUrhW5V1brc8MPd1ETMA
dj4glj0AblWzshPyLXGAVaKYoxqoOYXs6oD7uOeRyMP2+eEo/QFpEoz/F7wt/DAB
rE/Tg+TvWWlqN/ExF0X6p7M10jahL7gng4d1yMWMSQlyYrvPx1TL7OHoNlsDQlFS
LLEPrpdR/scuyLJwg53RfyZjB2Nk3V4kZWXC6c63EAAn24SHo8rm18yyZWc58fOE
rtJL9IoeNDhHXU13jjpUoc1Wtg54zQUpy+/KxuabY2DTpf3jd+Sa3vQevW0Ejd1d
yst8DblGtpsUZ766yMfCLDGsniHsjMQ+meZBkSwXPRXXPJ9oSgNr6bbr4sdJCEKl
rZb/gn3ZYyGylDFOxaqDE6ct1KPPjlAD9Ga18+qgQWsv1R60sEM+6Mwa1rRhM01V
CJOk9hTnWKS46sMlNgCSlJ2nvxJQmMExYYBa+ZTmld+9PEJM3mgswqv9/0oVD4oe
jcpHsoTOp8kJQ7KCmGm7zlNsmoppGjumzwcJVXzRlaN1JTtiLJXiOgxUq7hlCwYc
3mqdN8iPGFY+u2j3Fz4wxGbIBl9BbgabO/9EZ1NM4cgt65Iyv5TkmXrL/pVQ4UkJ
zpzkMLCrmBwhNnP0JcMOcA7DMFjHccN2YfT7wdo175wK8wnjaWRc3VjfYZsfaZ9f
xjKuGouW+FhCkPLR1bXE3qbUGuQkO2PD01cPZx3HSsHoC4CoyVFDDmKhEguFkOGL
fcobIlJQqqY7z0aNQafogwUI6nQXYvDfeWy7OaNGEqQKcRYOpeTL+S9JEZMu2nuE
RrZFsRiij2bPmK7H9o8BDGWq/5iklC9j6G3ZH/FxhGpzBp4/X8hXlzZgKzcZryBx
T1FRuHpi2lFvD5ZF4Loqu4Xb3q6iW2ULv1mDEljs2zZUWqEu3DvLFJKP2tHfYK9K
cn+ziDAv9PITblm2nUT0PewhJFYzeeapUI+Hqezu8LVIRK7HJCRo6C8r6gOnQnu7
DeQJvdS4oHfMDlq70xGihfRrN2Rht6sapb5LwaYCEb4NQ5NorycTgZ/+59efZ3ZR
C/RkwTPCvoAp3+xd3GpdpW3apNpqKkHosgSmYZxHLDtZAKw4Ii6EGgupVpQoK2HO
gGZBOAPzdMnL3sXlPQ5kUr/Z7ChnnX8hQASaEqC5NW1c2rnC89xD5YWzltmNAgv+
eLhIDXMBmxckB6HBY4X/VKfHCSBswUm6Te9TCjqjQR3VdobpVpDzup0J3uMTfFqK
g2s4mpyncMz7hbLVkcpJpvbGkfu9yA5bZJcAszNYCzTPU6Y2rWjP5laa83QITN41
B/1b0fK1ayrAyXl+R0qRlUrUpZAJX30iUYSvojoQ4sQLxQkO4PHkliEFlNShafhA
umxIcB//sihtELfsqbMR6skXHHpuwLuq/ANfud/PYblnIkczw/HRlczjXfQ6A6yP
3fvvMu9nnufl8McdI6ZoKF+h1Yj2yYOxd9V6+I+KHxBsbB8DyjupkuF7aUjBGM6f
Jc+0z3Jp6gWP94VCzU5pvLUvTiL3M17gUvtrLFW68e++mMJZsDWGfo/yeRq05E+S
k+JP1mSrR96B7pEeOLpoDg7OU7YTSufzT+d7+XRBzziwqhdv54lLy4HdHKrPHyiS
58fw/ddr4PH9GpXnSeu0ssyM00SNKewhDUgaw1VgzJcxnH600lx0PGSfFm4L1mmm
gK2kLRNxZMUzimKM7twxYtnTUTjxXO5kXomCHX/dXL2QMt256oaTstkmSCJ6WYPM
8IBOSZ9AY7CqWbl7OVOI7soQvsmlsdWRj/xUhMyLMEV9avMIisrQKSyRi5hfDZjp
wTjIeMVm4+xfY4zUTbDagzsmY0QyiHb5ISXxsg2al1F1sXW/LkrFpZTyfxSMbJkz
xyq1zH7NbzqabaTDgLGy1+WDWC5EgsMxQ4R2+nKcFg+VDaBTZv3ki8ZHXMfjs9Vj
C+v3nY9c+KVSjnnlwOeBNOs7wDaxnypJyIOUMY2HsLbS7qtwHxJXzc6aQxklQ2ds
+0JvLWv3Hl7eztWkD5ohXqbz1XAZJQnpY7S6AB5Xe1tWwd7FjkzD96lWS3leph9d
Y4i4sg+PyFumj8k/UhiGyyz77Nl59kDPaD5gGnkg/2+v68bDNwPnXzordq18z/Zr
VXVho5PdcVcJoIw0/kDpibVf8Al+ez98LC95rKOHiiVY5ymndgA5dsx7rAHtuhdW
7jCYF6GdniyeDp9kMfkx3qdlAM85cVkZFoyKrlr27RqeBGz4hIsfa9aqqTrv8Dpv
xoWYHk4wxece0qNH9VDghGHp9WnnKoCQ0TifVeUdiNG4qJUwdqyQSgXxXh6EhFgk
1Gwc597L/51DCT8ILCmakUctkhv+aHM1wE5Qu/Tb4AkrRdEZYiA9FFfet5mgPDXo
9LvoxNcgSoaSEagpLejI+2oBfPMAIoHYnw/oUz13mi7NAZNFgWtdqGLJgXtnAXro
8Td7ukA6Wl1zpbqNQILkb1ICDsIPUPEPRMxUIIex4xuFTZkP64m+bkqZ3ljkEqbv
fG4DaemfLeBhQrr+Fy3+ZALXDmZ23Ox7A+hyiId8TdUDO+nnkubaNRrLD0N+sJwG
E+j8iWPtyaUafhI1uSx0g2z5g5uCppVny2UffCnifwqV3i1fobVN7y6l6RjQqK7G
CuBIaO2HZGVJnFD6x0o18tq0JF4cglMmNUbEv++C1VJjxt2O8wx7TD2CTAdOjoGi
NIaXZ4HThqfB/0TORl1x3coF6iB1+C4Fq+SSOn0O//eri2CTJsrS2FSNmg719nyd
jVbrruucXVtjRwphyX4Quw5ZG5wftVtTzb9YKIII1E+t2kUo+CzW8dEt4veNVtif
QK+Tq9lwqDEq3g2b445Sj6T7KeD2IddA1i5+unPL7nWhTnpPgPidaGLoQ073b38V
ZO8Pf2ZthZ7oZB4EN+L2qTVXikFdgUkU1xyTHzu3JRfaKrKvP+jurrOc7l+sQ0UN
GhhcUW9HNjbJ4ukwGGNHn2+cpoGzlxmCBMdCIy3fzqZaQC0Qrl5kVN85H83pwejh
+jG/uCcq2ihVy2vN9EJaDBFGGr3CO/RbQ2xcSxnEXFcSZOrLuSH/X8YEyLpYOjFG
5aj2tPM/WBxRcipw2+m79WW3LO3+a8jn7/cjsWUsq/hdHSFE1WktRIWy/SKsgT0J
3KDIuJPM6naKIN/C7t+yNPYysByW2MUy7J7zGCxnmJBhua3zdulRDgXTdBd2FNxI
99FAoBYg5v6YvO2JjHFurqv1NMD3KmNiCtrlHYoDK74jdaUo6dpCNZw1U9pHO4ye
i9QXpNA5C6j3A24S0s1KwP1sLYflrTWGK44+gQ9ZiFFbu3FNXQvwjcqVcYfOQeZF
sTcx1+4/4kaJhFCpc5zilXLQYyQu2POpGRkWR89YD94L5pcOxTdtZj2iZNiCPczf
ospkf9CKI79bgRut8hdmZ9Ok50qu8+ck9qsEND8Otdb675wTA/3AOI2N/VbsPo5g
2UxmR3BgjltWnK/zd/QpSRO8bX2yrpAnnjCoDQDRwzQnHysSb8JYs+o0zl5YgmoW
WBIuW9K231rquk0TEXUzjpLFzwwYpb2HCiRa2ocwpCihvKsydEpSmtA8YiZ1mfw+
vXlU4HURAXZXx9Mv7j38GJW8cMYbzvCWx0lwrAIBAMqA6Ei3kp64GxqC5vYAVrMg
eII0jt9JfCpRGazDc/PH+ngMDcjFPuiBluvvroLu8NwJKDYkroIRyVmpT6iKJTYq
o7HgMraYuzcoqM3GlcIZTMaBGJz3I1TGE4KpZKZbFXUIrX1TQ/Ge7707AoqMo029
a75SScVGYeIRlwY7sxECGcUmJCDwMklg59r8aqHNs7Fe9iG2xU9fOMH1Trs0geWQ
wMfjLwi3IcmsqzMpdQa4a6feE6b2XU0GfMrJPZfQzO0RPK4uLuE2a7v0dHdBMdim
zsdH6o7K8f+vHOQ0ro+N10pHyaQe4/VoX/RbwN9/C5fqRWDszXbeXIsCgsSG7xeE
VR4kAjxAyAjdoZBYV4dvv2BiLNLj3k3+r5VSdCt2DyrIgR1yCo5EM9m28ylfFGCV
xqyNgxyblLSi+0N9ZYIzIr/JYAeTqvCwtbpJN5nmWcg1aYBdlJm5VaeLIy6F1/NP
HFzkadvcgC19pUL+czO61Oe4BKLYOacLFMsEG5L8EM+/Qbk/GYR+UMFlH9A6hOtI
vE3QosY+TjrjJqdmzjirHLiaj4SL10Gf4FerGX42Y8EzAM32hdnLL3BUrMaJriXp
jdV3RaB4teghskVTySE3o3j2PodxNRhUMfEyNmxumFvsT10DRRJ3M6AkHnbvb5pI
byqyfs/I5f1lkBskhZ0XEvMy4HC+CcUBYYYB0DPtpueL8LgIWM4RYxFjFvrD1lqa
M6goxZyAHiIgdxa9qJy7XZ2u1DdofxA0jOMrPVe+MObWaYXPzN8ebSmKrhUSGkzv
YeiQAZnT63ejvu6Ene5IwkmNnSS0UHTpTqb+RBZyi5z+CyKm5QvWU3/LcHV7pq1o
KGy08ljAZQqMBNvDvOKSvfxYbS7z9baArc2AMJ1sIMVULREFM41l8nmpLFNIm+TT
LZG+c5xNmrxU69reKr4e+hwb4qscakFSk/ztb8KPx6uhV1ON5j5VWd5qcapgWIqI
yrHF4HTWOWHdU0hPIiIuBWM5vjy41qS3hQZPhaUwA4nBPiVtnCGm3WqbOdCEfcU4
cijcBv9wI6vuwE/AImI5tJcn+68CYNoPcow4dEeGlkKcsuVAaQK9LR7/P99/UGD0
CYN5LctsxcOo0OdfXePaTFudpjPr5NJeQ5miIMgsIZIgnaZZYwUpkg1EBcD11kBp
iZKnilc0BlCIw9g6ZIT5U5W4DzLwRYwteIgW7bxunGPeeiTNWhQ0c7sFlBDBcnl+
5gaq2lAcR86rCas2jIP9MJNkNYTbTXBU/WB54dAxSZG98wuK4n/v4mKwNTwtmLQo
aWV+MEwiN2omFDm4S9f+Ze3NOxW++GjYJTzUVXgiN9n6UHqpGHlryC7lT1kvjs59
a21WN1aY96E0oGL59kX1TnnGhQCUXGhLe4/mSaPqswCIE4iLRGzs4ZJsKSg2konA
7PMOGBNyCfg7roalZ+NywqmNTOtukiVmuqe/tdVvEhsQIdpTGUacNdktcn6JlP/J
xUng57Sdjn7OmdY5H9F4/xd7cSsObEO9cgvwHlOzwzyA48TZnLY9h6z/wdrERbJq
ro8BwMkZ21AwJ7iLoaqckkFaHeABX1nFCJ9JxZCWQ/kErpfNF+KIP/I/RTlFkNxH
4Sw+3Ymrmz/mF9t3o3LU5F/J+DcEx+oxYHgqwyqj0SfVIL1rZg8kenQAA4B/RvfZ
`protect END_PROTECTED
