`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U4rU3IOp12fIniodNGouzA8eSKmqT4uzASgZBNUkGQu9APmzFfm8kL7AScmJIyMG
3ZHvUvfl306FYIg+6PSkLvL4u/ho7g+k4GkDLKEMEGpUZydqNgrQr+dnTJ1Ii4Et
uDbnHmTt8sMpUime+lywMKa4dusso0whdtN3H6sRO2QFTIzxsrfG4c2HXzG7TlLO
6tbhBbox5f1iUjWCmwlpNrDBGm38x5+tEeHqDSyc5SvH5iPieIKaWt1PtB3lFP4J
5euzzhcLdbqsC/eIbANG0WNP6ySqHvJ1w1bZ/zhE9EPI9drXu+wBZAO77/HPm7vG
Hx2zjpAZqTO613EZBvXhP28hVytRQqN2BSpYnzzOHtF73Oj+h0VK747nfh12RbcQ
mqPE+NwoLcuPKP55zFRVu3TYYNieWkUICO78BWfSjWcHLQEXcRP+q+RBKisUltw/
09chJsUI2RXbrcVBtnLcvu4snjRkRGLzMjFO69dNC9bZyC10hWq3aMZRVuVWdkv1
/R2G3vtrOGFHExsz/mi8T5D3GKPU9an0PDoC6sLBnWwzLASbxU5Oktc7z6pzDqL8
9AkolX5J+vUteRwhFM5hcBr0nuRMWNdnYSi3m1jtUp7WATZt70EoaraTU5qlHo5G
PFsf9hkHaLQmr9HJ5Dje+d5Llt1yFHcmiPVRHEuWUJ7vQDGROueJf8suWJCVZ9EB
eq3KVdZiYuMLQI+dgMXzqFZJmUmGlNugyFbuCs9Ku34YuIkeM4DGvmC6yYAG7tU8
2lnE0KdVYCOtZADzXqUkoEfesAflvDOzlIO9AURk4mucKiUP/DffbpzsSEPOxyN7
`protect END_PROTECTED
