`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UX+4f5nuNQe2gL9UjK+Ua6/IpechpjTTVXJvK9NcLlPMGsfc+Oxe9u/aHklo9j3n
/tWF30/1gPJVl0QHhMR0XdsQG/7aZo9z+PPxgBJ+35plBirQN7HYIZZJd6eJMoiy
2k3JwNwvJ+mesvllREyX1MEjmSrU6byS+OOTQuvrqAtHpl//9W4gTxqJswWRbESC
+O3JzEsPBdllWSBRUCt6vIYyp5wiAmfVLVeqmP5QO4Jxs3wvbuee+b6jNweoQ8ew
GN4YInLxMKksMWr+0ok5ypPD84JU+2Y+c+pidwPkw9GbpuqIitvSBI10f05knOoV
bG/YNes37ropxQkovuq+yuGPttWtcstoMnHf+4J9apBiE07RWAp2TObzx5851Xyo
oXoFPPOmWrjc0RZpehdvjEyfIktuVJ3ZGwSK4mi/jFjYi2ySrydDfyNfGfiteGW6
b0vAuBO38t9PMVD/B9RaCwR01fsvEDoHtCTkhN+6LGnA+julUyhmCzEWVyyZjH32
KDNrs7qQ033YLDN0B3L8d1/QfRkdedruD/fznMIG7Y+xJdlQh3GGMAmmV1kYLnHn
gpwq3YVZiYNj+ZHogzNdKTwoFDZgkz8T0A3KcQl+BHEl5D2rOzHUaEwJlfzt7HLe
QjyRNmqqCtHH3c8kRxVDyUsg8zaAqeI0e8c9kSgNlYqO2ImtK5qtSmc/jPg3A5io
+dvv27wnfL7JPX25SXMpbR9CTjoF/OkiPEf93BWsUnK4MnuHwt2VJUYg73zOR6ph
qY28dWuv/Dju3wmaoggAZh9ZF1nXeZrQUjoQol2HODxQGb08empC43EpCK2cNxvq
rMqGKriS+a/QD80ruBF02BqTe/IoF6icE+ZDksB9u60PskUWbtwHIDRnnKAiUf9f
eiWEjslYa5nnF8xfA03szDRQs02XYN/JBPnnfLUzOkQa8/LSAUjpV5GK/WGNF8yy
DjxzpWuzfh+6jNn46VuWSmUr3lIqp7+PUo+DBzl6YtLDso5TJBtTtJxLUZ0fi5zZ
8AMj4bA4FzIZP9DPPxmA7FrsTjC81N3vAZraml6uws7qF+jyT5Z7QC5j1XNcsAU0
XXbdgzyN8nV/OWgmH/22gEx99amEtKWU0K8g08MmNwSYLuTMpGMaKnHHwWB6Noq4
hEliIZ1dTiKZjIdleIPStDXXipxY++LY/Y+XlzOxGZHw5Xl49yQoFIcCcSqwiQFj
OdtHaz8FRwmkSVaRzUgfvuLHZHKHqy1KGk6ZtcWk64fNDmKvlWdb1d9LscfKM1qK
tg5wG0QMnPqfZz+7jQ1/vE8ouXqjV5wxT3kXtMc99K0mLlRfKaLc5EVtBEASX9t/
dOADd9qJj2EYJlSA5TEb58NWIiD8ZaROauoDKyAgnRQrwFwCC4rfALHyfx8zxaRE
GS0e9nY1Wyom45Ui9Vh8LpKxnihUQN9J7tUZxLRNznSGHIzsEcL2++2MMqJjbOxJ
Y/HLgfn0nocPXztT36+YeQMnricXTC4o6bWoq9l9GPZb1cAaCkIjOETCqPF6ZYmv
sy2CgZ4G+lvQj+g1Uq0+2JHGew4WKuBiqQmEUXPGWIvdUv3M5PlMYiiuTNxCkpjK
OdHPWcg13FO5kE4o4LhEq94lwTIFF8pt1MzeI711NCR2f93yG1k8swfFm+S4BuCm
kt7jsCsCF7xpmTOY8louDvhzB1raSdMBzgqy0Bgo5PSA7m9aEWsFWaZNniH3dIYu
OqwAzSsZlCFkmEMJMgxPuly69w71NkpNsbdp07hG/XGqhfs3/Vv8SzxE8M17T+gW
N5eKwGc7seaT+o2Yvc98u/EcULC5RFvkODRL5L8B8u4cxH9dKBLHSoZ2Sr+SfjND
04WRyT71UbNVVPNl8k1PoKQgOTcUlV6u2DNCsICrj6t+Trr5Yu3mqdux4aAtw/w7
eKVrjRZxjJMMTw6CQdMowe5aVKoNjcy6KoTn3SC6tVO0dlCsiGbJPbcV/SIoEJVY
ZYPn+ZuBhGn3k3abLcammk7hhSpUk5pVXsW2blK3J/dGcg+4+N+ujmcH8rZwHoyh
h/zqV7UvSdlP62minDmF6YzkNynAbkkcmL6djv++VASh1FIgOACiLMmD0+VCpRa2
x1eYa0zPMs03M+BeCFSzAc25LQ6Zakd2ibEeMzSFH+yOTWVXA7ZgJ6cXkBsoYL++
cnQVp1Hj+Shl4a5VcsIsQKLka8M4AawK6xWJ8audzMrAkeIVFnRtQo8NPlk4xBYu
o+CSUHTkE+OCVICxp/JU/Zo2CBkdmSZPP7EGFb61OEeAsfNCqANYCTMoioqcoJDg
9lneXdb4L6OTlbDMFdW+WmWs3B0B6jMNOL0xdchrLlndyldPYWs5f9oTEK61A0XX
P9jU/CtZA9aI07Gq6bfaVuXy0ZEYuH6fmZSdd6sGhLsnIpEMTnXLyoi+31ou+sEg
PBFSXCpkSkuNNS1+Ai4CKrcf3GxKmGwHUvqrGQlpXnCd5QWnluvB/alle8iGEs8X
nr7isoUH2MIJo+vSlRYxyFVe6QeVLKn56t7O/DToesDIZk+XNCBeliG8sG7inAIE
3LNy0ZUQyo1fcjauUNi0EQ15TXXhPTlV2CBqtXvMMC+oflKs6V4YPMvB9zbW26Yy
aEvYngHnNyvV+/50Mj0VUKKDC0hwiQeuPuo4FRc0rzodMFYUcW3D6gkraXP46gfX
ofLnAkzmIkSexYeLfrptgonX0k0G/0hosclmW03d4ggzBTiKJNSho6ibr6dAjO5f
+PV3NQvLvFCjxPFiHsEqQOAEeMKrc/HxjLMcg5+Jc1qN68/vWqEFEdULE1Yw37OL
zl9aiF7YkE2oxivbvUwWgsKT+8FpbtVGT0BZSUw6jEtkpLE00alYcl37w104c+Hc
ueSCnHiN1VS0Qo0DSSeVyAREU5gBqJiGYqkTpHTVy5NnkLe5IVRize6SHZCKEidz
nXoNIDHTNW3/aK/lFJ+L5KqVMw9jVWQeH3RdyGDtBWcFILYXizZ9PbIuRFzNxWhx
VIdUKa/+QgbIPH9S3QBKKrqzFgm8Se0GuZP8/gQ5sglDBPg/um2iC/H1WLsw5IV+
1+xh6L0H1H0F87AxxpfE43UVwvHKGXuKayfBs/eKk/7BScxoMvohT+NVNr9KMm7n
+ECwvIL2nnhRG9onPEwXSIZqEc/ktrUWrXb4VxjooN0=
`protect END_PROTECTED
