`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p2w0wq6k16HHaq+nhUWbRgh2OcdnfLNVEf5TZJAfxQb5n6KiSZDlknW41n2I6xCd
7n0HYsOuimwMnrUowyYtzB6o/DvGrd9ZUJrHgi7ny1tcj0WZKni2pbmqoB3lmpvD
ofBRJXZDf6YcxjCHxblIIdqLJxMLdyjR2QRyLxLTJt6aFFsKTBWSrE26kiw1CjTh
EWPFFBMZ91yHEP8FUN0LkECFPNaitc45EjpKKyRXcJJWzkpdcdjtugT7Xy9/R2dm
ETT+vLbw18DvHfwLFEBHkFm6yQbrRrZ3w0qMBYdYWJEJN1jIOoiQfBQMnNGsIgMX
v/JvpPHaFhMHdHy+rJcNyItoScnr7BTVXlPzR3EItW5HaMKSEFHriFNeMUyyW0NK
kQpKO4klcxAkVWqScvf/BkOLMxSVcItmgElFrjjnMfzoO/wiFSGxabouDojFqH4+
5BW0XCciXlLn01/nmpfiQhfkmsxWLC4a5EqVDVImmx7CY9/1r1v1aqyyo/nuSIqW
KRV2zkaUSlnAMvsZGfIpoigr9U1vuKdQRhWujUhD8/tmyVjus08v4Fp6taXj/wDH
x4Fx4s0TleWybmQGOwp+k9dp2loA9B8KJ9TY2/7wlRomL29V2p3jI1Rogo3F01Gc
aBicSZ8bWYfAe6pGVO7dMhOoVmJv7z/xgUVoO3qqeIeNWFJpRqXSwWmOvmnzw3TA
UlTPBeX7DwtbODJc5oHUlGRVzaeuO2BgfGF8tzaRSc6BM7ZxPffbjyEQJlIBXKWz
jci2lv4U9UVxx5+RaaWf1mdXtwtQraMqCtpOjLSuPMyQm/JfpFtJFkddWCzoBLT7
wStGa6PjdqEOgIne1jDo/RlHa+GAf1QA0ky4t4MxRDBoyOn7nJbkRHeKIvVZiaf2
W742QFwASnlw7vWn1cd1NnYOmXnxPDD1VW8te/WrnkwMuuxCdK3CQqqSpUSYIEm3
kIe4zl0qZ734yATF/6pcuA==
`protect END_PROTECTED
