`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v5r2hoVktJnddZkrm45aj+2YHH0o1OTMfxGm+ObrQh+EZc2bz0vKvMwX0s58krp9
ZyqodKg8yUg6KVparpTTTUq9uYcBK/lOJxfSpQMDUvAWgd1ATd9kpM5dhXXv6b0d
6ABH19lvYtlVR0Im9ZUAYFklIVSgLSb5PVKmSY/Zcf0azLNYbUcJ5540OLLmnocH
iOHy6G6vsO5cjv9mN4m6vNugVGUKeT8miGj2wACOATHsRDpu2TSWhtc73bAT990j
plEDexYlzDK+KJ9ybUB9iuhILKnc59hi2eBO/66WxHIdOc89i8XGwg4scyb7bQuH
sRyRA+FGz0dppe172eCKmvmnXBBLSB56Xd0UegBJjJf/sy5muz/t/UCdyn9EzF0F
elYPrXY8qCzY+FZPN8EXnZYY7qqJg+gbHv/tGusM3ss+8brg0ImBlc9YbN7T3X5U
pOhXQ9IGrOQWu7udK89n1beGhvv4t4bu5bpoEMtaKorbbQMN9CuRR8LNHD1/xen1
3R/HQjh3b8Cn5Wme+279QdeEKmNs/40wkGgHCZ77PJjU15mNIqohMf59QeKpB2CT
vFoOtw6WmFddEQhiXwBdHlpciWb0K3qMBCVFnM8Os+4fcF9dBBEiqmfYCdL6O9t7
bB9LMiXqEKSvdYmD0ZWIYGJETr17a/3a8s0hfEXQ2S249GM5bvgZMuP3B3m3ENZY
643WXHySmMZN7mh/6k+x6bHYKGKeGk1QZiYdmS4RVLIKYc471sJ7+Z6OCDgrOVW3
uo+1nMmsiNkHxqElHiRcZY99j2ydalAC/MIy6Ldv1jm5D8EwtftRoA76T5Dn5HIW
9lSmeeHylgAMO6BSCqvkVJO3RyHUfzehG8CzTYsuWlfzadOn3/zz5DSEFZxmH1kz
gx5DS/F/FcNebRh9M3Le1G8chbcOrOUWWp6aDgh/ajHfL+vstXRiLrOS4lBge57k
yb4SDnxwtbV4sSTq1bJil/pwAIGAGWqt9TEagmJ6VoqeFj09UEabVbzNghcm6Nhs
6tV/Vt/G6RlVLjswUJTeSawHqqjCKBqQMeDciEWa0ee517/3t8gXvpX/v9P+Q3Zx
ENDigvrwlXRKaBV/9IrhkwqwldIPy0/ByfCkqeMVPBHpNt/ueGB3+1ONcPcLYMtP
cF1ML9AwbNwAT1KHfpBsJdRGH832xAjIuhOTceaLtr4T1/RWWziP8H4h3wOXHGBC
XQPl2GoYIDQDiYvRk1poDtlX2w/OOrAg56fn69MYYkiwkSLLfL9FQJZM+lI76/hv
vcP0g3+TSVf4Mm5Yrc4K/mUrlO8KBWIk6bYFxpRurOUQFCCecmpl+ucTB3pnsNhC
R1gKkqUiKJVFrWYY0LtYO/G70l3iX//Wa0gEs8ge/TJkyr7nCd56+dP9Bb5+q2PI
qNdFR7UFomRoMDnKIdv0pBnFbiP9I8fjVeVngzqpAKzQb6W1JRi5fcBCYluBP8UQ
Ip1ZDLw21smXB6fX1SWbzFRAJ0SJJsSyBmBOjyVMLTiB9XSR60hkDsNtA3hC8RLb
UuF/wG9ygFBVtWRa8oe4ue67vBAVA9z8vUZF/KwiXVXL1hHQK5wJ2GAqp2qV3WqK
h3Geiag4xnJB5kMXs8mIN+u6dWNJm+SdhX0OpX7iXezBQyVAsdZzjHBVqsL8IQ3l
8ViLELLFMGr+MgDB9eDN94QHmJOmrQDSn5U0m3SNpfsS0PTQCEX/UPPDE207JJCD
PRhSd566O7SkBNRMZfJwoc9KwbyveTecN/5rgbFJy0rovcm/MREPn1qQbXI1LJwq
q1QI9d58zJv/KKxaZq24PdjPgrKMgC3Hv3nEvORsqwi27pOiPJs8nqB8H22aXxiX
JnZjTu1J45jfwmhnXEJtlXmRRrCe9xdG7UZCb3QnCnZcuh48MT8t1+G3O9hYDEgw
ZUMraMYpa7+FVVZZIW8HWnEeVlOQ+ji1X8ZKK4dmS/tXdZQL048fOcLVZWGKyKKi
EvK6LJ8iDITMjHi/xb30rMkBmvj5O29Ixf9NFp8FOiW/ZuDkgD0mu26sjHD3N1N9
uimA8odejHY1l/v4HajyOHXeEAS/RERbUIwR0GemSnfUda2LL8R319TdIbwPXXPo
JRF5ryDxVl3rQBgv/qzl+a4yCiej3zd1BWGqMMHdxvNZOqqGrEGcRb0LcFi257eD
NFJahpgHWMVHMDwhTxfFYPpeS7TaWhvJnlcQlmBITKF0khAS3MKm26HqCVow1eAT
c9KGguW8pviFm3DtG/c5y8c3KmYCxY14p2HOMQOQ2FztXwPhhoINrqgAzYl1X4S4
QeiGkHbcuxiKDCtEnyoT1jBkXbGPMMX0c3zwsijrYuk+bNouDIuw7K+fHwdOXb4u
47uFkNr8go/oxRgw2m4OJi4/IFlEWIzuxKY/Nhsaxrn291ETzmqQJ+DMdj/Z6OAV
Uax1CZIU3tFt1NpAKDWK1b+aTWZgS1b7Ey3KSRdIDSaEhPjO6dvmqXpzBYbwhiwy
Rhz4BgIMkTDO1eJW8yI28SYC9+K3TXT2+YiI4/NjzV8meeU9l7rOe1nZue5i9Ey8
TRdt0aMVgvaTySI3jHDivZU0gBmfERJk1lrTLnBXcMMEtbcMmErOGqDDRudZ5hou
oX3CafGRZriXWpcL6b54UWws4T9wJAPXrXgG5RTLaNgW/pc9sVT2FOZ9/RBfi2gq
iwJT6xhnx7MAsxGuZUtUDzeEfPIBFM1/7EKAOIbh6tmQUh4BxXJM3Kc4jwLlfTUW
NILEjzpCGROkZ7NE5JGdMaADE6mMBl/ix29sSfyiJhTq0NGJn4TyhYxBA63G0SAU
da9AOuEd0fnMkUq9hRqmqc356yxDj9Gfc3G3VsDhi3yCc1im2GQag+Xza3iOhu20
SRGr3qzYodA23i2Dcp8uC+9HPNmw18YZhtTmYL2a6p3zW/4qjBZ9OV6SwK13RYbv
usz0fkzjsPoE2BVKEOBkdvyr1rcgFNVpCx95dSNS5so=
`protect END_PROTECTED
