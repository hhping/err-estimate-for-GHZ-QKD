`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jlVJF6TSN6L0ID8GZ5vKLeWDTFIVfyJzCA87PpYRTcQdo2zw71ribvrqXRdNwsnn
9JvakHyi8jeebTVNiXw+Oafjr+GCovsjaWyh5HY5KUuL6hlGh6lE7iTf6xzbGDdp
v+Vlv6An8/WnY2pAOY9ihbN+sL9tyuy56groQnTEkJZFOrXbaP2ptQSQ9yUFn9bm
BhAHy1JyQLF5O6OA0YAu+5Jh86yH7xArISmEx/oCgMnPettxQ0va5KSBYyvpIysK
c/HxP8eXVJcJ+m/wADGiJgWuW5IDiXYm8g9eO9ioCFlpg4HXZbn/Bs60OO1F96Nr
nN+dQBQzbUazK9LPJUVunICMvshLQzW1Vv+CtdKGSTWTE7l9Q5tDng3jowa/6Mxp
mlJxq10g7OpVLbvP41cajkaIzkf9k6YnqublSvCyY7sGPGrRQhLGiwKlvM8YV8EC
hhlv4fE6n4mXYkL0C4VEIx8G4PZqjlCyrTe883yx0SZq8fpgTpv1rctRzjlRZPbh
BmiInFvtKkT1RHkURiU0ZG5upMfmrtMBfOaauxx50TVK8MHPEUswXQfxCj2e9Vpj
/AfmnXaoXBVc4g0KqVhTZWPJr8x0Q2ccq3TQmv8SmaOTP9MHSuZJL/lkAJbbvk/r
xeGVuG7MkP4fsdZm5xFwt10FG9GfKdK8wYTAtKnOs+10rJf/hSMDMztltUWrFUCM
lwT8q7WLMlGZK9AGwb7fMf3xFfKmcGs76szcpjZpSoMEFcuh86Ve5hhrmUXMymyy
3Beiu01ODx/HrTr817h6G+uuVY/4V634i/YW8S8cKXhrEhmSfsezQNwe0uZZtkKM
dwhpZsRS7iF3zpmHFMyYWDwIsUfYcCOsyQsbaO/55QgLmr/Hl34ILnWyxrrySOOa
my1BfSi5B07WfA2NDIWwOSvh3GHralIDl5n3CvBHgZveq9kP8G/gijpXrp1c2LWC
VtfOGPN8XsYBDwE59BcbImcAM1BU1Fi7gjy+my8l6scZ1aRS5OGbscrvQmQ6mYl6
sNf2iZyQG3rYrIeaKP7KJs8zsVaQEjgA+wi8LSThA7swIuiehCRQXgTvaGDl/o+U
PY6SpYFXiRPSbDbYHaeIiruVwbtwHxxW1VF1cCIFhpLWWjrvyEsr6l3vJB3ITRb7
ITemdxa3WjdztUYFq8fpXjz935MeZfopvGZt8zwip8g=
`protect END_PROTECTED
