`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w4kbkEv21RFCpIPmAT/ousMduM+ZRbCNuV6SdlON9Y32E/YCughg6Y2pS4SQvqF+
gHiSzax/Mja30W1gzGMgiQws/0T9WHQlXvWvZSlIdB4xPNHirvopeMGo0oMAOpP0
DAaXlfONB8qgteM98hqAw3gUKcwge8jEwBsAozOyc+C++278ICv4fPVUAXy3KsSq
TjKHWGKNgEnf80nEGKrstNA6j5PCO2yGoS1qtGcJSUgmiEdfttOVZ1dsqtf0OMOv
H3ARqeOWbF9SJEAi5c0xKLCE4U9wIq8MiZhsjASp6dBuYQGHgZsV7cNLHlTkzMhF
v8xs+9e+MOtBAny2jXv6bFfHG7M5j8VMKbQtusiB32o3akRVKO0ghDPTximJiMmU
sqJR1RG3vt/OjFzMS4pr5p5hQWhmKOCfHpBS2hBSmTVvX7qgyLV7dkOfJVC+8Qqy
zf+8Yz675bzaMOAq5XxBgW8st0NW13ITsD8EKBVgh8vKLX5GEGKmWgqMgIfV+T4b
69/tkoj8+7ZCH2zBwKIGRWPowe48VrGWDaUuvA1suwt2G9kJncpKA58hO7kWJIJF
7FRB5XvpLxJxpoIlpDrD4sARJUoKsbM8z0Oo8+qvkMiTN1Hf3aNI6gR0cPatPhO3
ggAye0TIYp7Vk7UMNiE7g2Vimm8R3A4kzQe58phVHUujbE18RspQqP+cTXQF4FoR
vxd4WymCUP2OVVLiUk8JCrwqbd9+cV+qG6es+8X7kgcqPWQWOaVC2jm58RVs6WNc
+gke6qto/iNjagOF9PLkbKKxrtcpYobR4/yPNdh8XrnEh46fA/D7wCm1tPWFrjiP
QpWG52Pm3l5aO1r2Rziaxsp9WXjtRCYIHQmeeCBGaBC6cSueuzupHYuPxY5VR4aD
ETOrsxBRG1/NpA83YO30mqeAwirbCL8NFc3EMGohI8ido8zD8SG5ME1W6p2JMbUC
fuc5Fnxl/qZHhJhBmG9ZlEGL/oBf/Xbufc3JUs+VjTC7W+oVjyUvi30ltT4YL3s1
5n9pnL4oyEh7imPyYaJd0Y5RaaROPiOopP8X+9as0IlQrOoZWMZo4qWxNwOk1NLs
8jLCnZ0KCgegpa9qFkQtsaEqlGSIao5QN2CubVQ0mSSB6QgcUTdrT5TpA3ov4R9O
X4IysPpIjLD0JrBPM67CXNMOA8YEp2Ec3jIjsMmVDJYSvoZZri4aY8qPXsX6zgAZ
5Uj4mrGEsF3ozbH4XMvQedQfg/tBCMUC6hCGpTzehJ1ro8ZEHMc6ewhXhT0XjEK7
C5bXoKgIMoy6duEzd1QdPry2jfE1ZUDud7BXE0OvEzS848fccPhyuSLJssHB6DzS
WzBD1Q8OEiO8aEsnp6z+TEPDOu7Q8+JqUqMjByk8uEu0gTvW+l0GyL+Y0KVC/cBP
EktVYKTfxqwksKiiGnV3ztsVXB3hopqfx8WdnX4+TbLYQZDhSh/nkgVVSeTfHxqc
AIaT02qEfmlIyuq7QCKysMzY9HOtYPwgazFz9yNzb3iOnqZieNnRnp/7unmO28A3
bSTi2v3IHQmqdyooMCsPKiNHVi5hemAG4h7VjKJt/ZsCOat9uoqeJxIBk/uXhvhD
+e+9ZgamMPWgeDKJT34kIy05pE+I11LTyNVwjEuPiRIABTFhKQd9XD97XjgVlK9g
UmxcySC6MR/MCkJhsgIeoP36ZMQ8Fq9WAFQT5qMYjLUGVGhojcKg6MeGgDHTdCta
U6MxjO128yncwWide/nbsZal9h6YjugMoCj9P3O2rEx2SLKZHVQgFZAF8u8a1pgD
KMT/7RASPpqPDV2+UKA1lCnDM+sGoPvs8CxhEelgM2qxvkzgXdwX11k5pRGZwDVJ
uYPOXoUouFOelNl3Wq0jJtN/FELpngXu9p8um6VIGmTVfOO8w/gQM/mnTRgkpcL3
zTQLk9kJrOvrOdLXaHg5+5d5nLCND9F3QjNbp0FQCKIIEGPj1Ws8rkkIkXbBKdf6
Gj4E1LnKVsDo+bYZOkPJs020HGlN4brR+QyHM16dfeNgKomjr5kBVg7vuruG5tPB
xR1cwP7yCFHLec+qrVwUe8gk0ZjP2Hj35UxcT+Xcuf7b7+NsOKWwyJ82J0o5mHH0
SpBcVE/FEN0w2o6btltaOoGv1wFp158vHKMeliVQWiozqSTshux7310vq9uBhxVk
xPfX5Bt82U4VhcSaJTldYeIiazBDU2LcQPL+OP/RxTrrYcg207QtD8Fd8I1C2H1X
wfbLUC9kv1QpSB1LVzfuud1H57NEiOOPWS0tW6EpHyekhaXN15oOyOqbjbCacsCl
xJFzTX07Yywx84pVXOLB0skBtxh+toipBlSPQW4pfE2GuH+UGlAavoS0yp0aGAWW
WoVsqu6Ufsr3olZmID+cdvdwHWVt3Y1p3CUGcry8v2ok992e3JaiJH01yMc+8ykR
+9lR3meQC6HwA0tv5lQsXmCbjvEKak9S8ulS5j1GjT7R8fiNDuIlyANeAR9Kqcq2
qF+HgX9PZE9eAh7VQpyZf1KlcZwUKOU+JKjOoJNrXKzd4XTQA+ynBb0/1QXQszim
9W8spQlycH+0gy9gjTC+VKnwEd4odatD7M6l+WuaSy+naA0LsiL3eQXrioDYn/eS
8bnj5xRON2Do25Jw+HP5xnAyGyAiq3aVV+j1Vy1pLiKmQwvtme1Z1DGxggrgVBOx
acvPgyzXkFS9FLqflq3voTtqqGaMaxnUvVOUkO9hLf+Is366TPqR67+byOmRsbXm
xfbNUqoQ3ADX9hHF8TwlrvXRyLrZ/GgGa+F/cW2U6KtMLZqZJBM+Yx44YH9YAiL5
dUHGRrvcDZjCc8SM0nk1Vpv+gx0KdPpc67ehHIkoHyWhMW1SJ0NSM+GxRqKBHD3c
RQdJAQ0547sq2XYOqPZKweX+rBZwxAfC5irrg4QMqiEZo6iEisnjTYX+nXQiik2i
7V28e8PnOm1+9IstcuXISuZsZCL7VSjNrPV3l9Qn7nre5OCBCuwbMq59uwqBRpXm
FQQDvKkLPdFNqyocA3W/+E6agB5nmObMWhI0LABpUxjvpkbOFfVLc/+SLOisqYhY
ayBwbvDl7gy8SALa0wSYQRQVycQ7llnt1lG6IZtydPSSSl5tXk66VR0G/jXM37R1
5dftkEhZ1CHS748e8W0sgiLk/HndixWnXUe2F9n9ebm3HOSFy5NynmY5+yheiP3r
28iMtfdUFK0T7KBVhalUnjOeBnIGTFZ9YialMCRNePAGizm4fnSQpjQAVwW4rebi
M2NZ+YgQMTZLmdPvs3DOWX/wzDq+hxuiJxuZcJOFVdqEaHv85+pteAEycIUnuvCT
yhUuj3ozxppvQBl0yvUDguVZgiKDeokKt7qgJqiU8qw8rioKTJ9DmZ9KH54LWvjR
9fe/qtTNNuu8iDw372vTBd7XQ5N1V1tj9FcS/zBo8CccF7wLoYrBnlc3rODqlDxA
hbfCdBgBin9bGo8TpxOceoq99/l9JEnDBLVEywHAB8fHyULdPZJMXGiVmuDbCva3
n5GyYrPllOW24epWgmEWmGuOXQ9q9HHwaqrFSsjb78p7zHVxfIbijJYa21JtDfJL
VDVxF9oUThukhWKyB/b3l6byBPxpibcBYHrZEp8tDJ2FwfYU8KMr6BcVY0Mf5eCJ
E/w9OiwRvFHHWc8ypI8MNRFA6ERyL0e8LeiRPeuCS1tTxf0UmD9xoLio36EwhjFa
afO2pUbg89lFuHslK1LpkygLbD/nqSSaM0N2kDGuvlWItdNjyD7JFeObh3C767FR
/wQtDpmwzE9yJCU+lfQLRWKpgKTTj3sbuYoHB4R3BW5OvPZ4Q2C4zsnBgUcXIvIF
kZOYIpH2tevNEMX1IdNPMWLJsVP9NRSEGj4Bj3uZdvtlikKIw5BqMHAsfZtjN1/M
TH2JYW3EqKX/eMBqWWec0CNokGsxFA6EBhsnhPF4mjfNYfe5ThdzQZJsCQ5rXziQ
kGhkVVnlsm3Px1glf1p8t3r87z58076ZqXtpULHp3ADAU7ttJprroJsyAyFsEy6H
Kbmlc+tA2kJIKeKEtuGMw0JlLHfZxEj0A8cT2RAE8s+85WJIg1rtZsp6puNmxBzW
pGosB/Jrphqufh4LDOsS4geKAXjQRKB7jqLUfv5zQSEeagHk2jVZZAuWsCb7LjzQ
ih4w7C9Ty3v67rJhRgKkMDL0LCk2fDE02TvV3j5URyCXoUnQyJHNvgR0Zon3JrW6
uyUKjpxuUnLFSZwjcAujt+/cE3sIosi5YPRUwALKls4ScPq4eQxOdPHVg8VuOtAh
b1dDlqFMdFBmNz4l8hu61YjTzEATKksecQdwqUF51uk3ArmypqvRGF0pe875fZWW
V5J2F88fLHS1RgrQ7oaO1Wy4SmftR7OYfESEsQXc9QFs2HHjcXB/jj2mQTEZ8ONb
KvxQEd4kuMM6Sr4uwrdWkCpaBlsG6kPj0WyCM2/ksBS5VuRMvMWifWwE8QUr+BMt
EFNs+jlIbzfWjF18EzuMRaWyLz1nMx/LMiD4eoHCB81+nMFkZOmQ1y8yiblQfSG8
cK7Wja5OwZtvNF0bHbzB8/FPPPN4BmeMuL8ctf8OhDfnO0IuDWiCSGMYd+5+AVkY
tRMmsMnW2Wu491ThGFBhHftTeAtlgHGtQSW0rr/+mWbnb+3VXyvxxZhbO24C13Ft
wo76uQiKeqKSoX70/Kx8YSwGnopQgvLcgzx72anKNWQfBKr9bL4xy0FjxPfTUJnW
DX2D85pHxPNEfCn02B4C6cCezO/4ggFuWkZLaMYGrtxaT8FO+vk1/2gjzg93+njK
KQcuToLcpD8ALrzdpBR3zzWItz7hFAz48bTKQrecFpFtFliP9J+kLlfUMfmCT7VG
98MJuV4tn0UuqymxIYAlkM2M9/Bcl9qh37X93gTRGnAzs9x+Hb5VdmXe1mBcREmW
yzoggQ9cf1TTi1N3NUjAqEXiDkbcKsh0bZh2os+FH57LzVnRH+mwa7SfmQdki8RC
5i140F6T41rKz+ytO8f0D8qFU2/cYgAywQfJdAYF1V9DuQ1uOri7DY4tT4TzGrfH
rvFynNbbecUIrrVUseJGp+kgsIbTGMPyvux9kKtc5G/KseB0FMa4nSrMmvHe2XP4
Qyzz6yPVOEBKVegYzYj4ROP4hw3X8Gx5lGdZ0E+R2qvNGMnIoVcZKzFKouenEyen
jAuZrbFaWS+snA22CxkMDwkFT8Wg3b8OryUdVqdwxlD5i3vzrTGnGYu6iaVFAV+a
2LzjbNzkYC07kzSxMo4GwRRIa6l/s7S2VVsITnOq6SIg5u9QQ/+0C7UlprYazOop
VypLobZf1TjNIiSaJPESwe6bW91/6E3kFFk646npQ2DkCuJPeXnR6Fv8x1XXTZRu
HHlq0ltBbUNznKo3eo7RdEFnmy20pZa0v9/5oQKxeNfitTKRDdSbvY5skiws43wZ
8dJKMIGbfHypz9dEfiQjZjWug5epv3gRpJGOjgXi3/LiOiH5rGN//d43ncuMEPNu
a82Mj7bH2of/w6gK/cwMJuAHf9atl+31q5fLex0rmeU9oR0NePNSEpZVwPCPUC1l
BXLjT3uwXnBDeBeIVvX1hacWfM15ylxT51gMya92UvN3i2F0uK5CY4TvLUAVcYmm
OVd2mNwOfNVV1w/P2Wcs0A3Kdso7KinZZYd2lbPjeM1QMxfGt/AhBUYP2+9zdNig
p0bVC2HndQTnlEMdg+ERFq4J2WsL152eGz6I/oStBll2D2E+7sEK82OebyQvNv/x
mERliPFV5CTZgD/3jOF9budXtHuJdjpPMUdRXnYfB2FAeorAwErzwK/qwbUClxrK
EHR1J62LedwrzAYbG2kB943f6Rq2sYz45wKHKUIIjGWEZw8uiUd393OTZa1gUBU/
VS+Chw7F00YKftCZTYKUGAHXZSooQ6ADzHDFQZhrXNRd5/URNMfKwxdGhTs5UPEa
+zGGzfKpZVJXCo341uy4h1yY8uVNz8fIUf+eaT4744pQW21ne8kwsM8DNhCneR4S
nfEgtMd103NzP8fcV7AN87YyRurjUyG/HuD4S27ronxf0Jx/yFEefdpWRgIm0agy
AyxCPVRFMQO0A2XmEFsnL7L9J7bBkgBYqHxik0bS/tGceQbBoggR1Dp3O92LxDZ4
eU3/1ONNdE6oV+wdQGTuhno/i8V29d+K/AddZ9k2sWnMNh1IP5kntBC9GVoCs/33
Lq/nkgml6umd5fIrZ3UHpIhC3gcB+/MED9+ZShI61zGvgKJu2fiNrGTdzjSssqFO
J/IkZRQpsC59Db2bvCDOpMyZwvKR9g+3jaxM3OvkvzUnVfs5aAKvfuE2W1OYLI8o
GQkRctnvAbg1o9NqUH5hhUmoOeWQGzL3sbZLQqlXoP95iLmlNXzo2O348WhcAvY5
1IgBGZSp0gWfJz6U1w3RB8zAwcRo9pT/xBaR+B4FF2KNRe424tZRJvC7tdaVcY/n
FapFlXjRE0TVzhdzDTvg2EV3rxHMT9rwDDoRP5jIslWQ4XZyKKJmfipYv/nAdvbk
BxGJQsmL5K4K1Z0mwhlQknk74GQbmKc2P/DSfCvOQI9Zqjs0Z7Ue1+EorEc5Va+Y
luRxZUk/dR+scv7Qyfj70i4uFn4Q9/gtH3LqKXQrJ8ZF3VkSCFw4qFHQ7BF77o1k
YncwC5lPOXBzrb0NAxmegR8QxVAynqYM1ZiVmyIHO2KgEs+KuIb9sQTXQCyLbrmG
IOxaZLo6LAH3b29Qi1XsL+UnMxgSHoVvdJHo2dO9tgCsbX7s5PJPqyT9mZNtjjey
P9wGo0qZxiLHNDFcs9njt6KcqohQEMUw2jTUWSSBrGElUhBNZOWEn4CVxjkafxRL
v4UHylluprIdGVB8bOjw++ta+/iwGQYtvkCrbTeOzGv48W6pdgz3p8Am8oXwxLNl
FRz0u4DY9JwdP+K8mvd7clctqg7RCBT47Mmmh+R2VihBOdPAWLK8QzpXDsim01dT
M+51XfHWz8JgKVReNHQKraShYnC5vHf/JRe8GSBDwsu/Ttdq9cWVUvUeDrNwEqMj
L/9QGiGO+b7BGsixFlTz5B26iAqNYwAnrQD9c52F/m62w2Xb2V85mGOS+ZrWbeiv
TteNpblmxLd5IB9o9qxA6U6YKNIuORn3DakL/Kr+S7TX1hpNkGHuP+Z47ktqZQg6
Dfxm33+MnfjFBQj7lYYlWk2w9dnkPEQWqPGDT/WXhZodXsM6LqRrJCZEWAiLqgdY
AzlqaMTzG8JchuCXXrRr9eyUZVpxcw9ogSfiRTSomC1la4qMG15sLDB3sRSAtIiB
Tgjh03JzCVn8jeGdjzGk+8+75DVYdFGNLbwDnmsy5jYQlbz/nusMjFqvXalJoE+/
Y9+1cubPh0rzzvoe2ptq65f93PrjNKnpOiEL6I6u2UzYIwwPyYihTN7ZXMgQYEC8
1Yc03YJkAeFqODk2wY7rtqmcxis5IN1Wms3sMyyUp7TwjwOF52bP/5J7QPVSQCr3
bbyfZ1uN0gVE7W1sJDvpJ2eSZcDYyN4T//ZeUeU8szeboGplScrOzdfnLma/Wp/6
u4li3F4uDHEVmju6lwozi2Mx27js7Dbzzcrn3M653IhOIQaSGGqhucBtyD3TNYV5
50NuAvN96ghKKXibLuzOK0liD2T/3YSkBevKiHPpWav+uAMt5IQ59uJhGufu8BpQ
a3iJ5LVNcWXWXI6rRNVz9Zu24OcSUrFoWZbXBXQquRFnO4hk+tHbuCfSnL8YU2Dv
sS7jDbGWuc8PoGsllcnEk2F9nsHZ7rPDO9u3efKvbf2fqudnaxIzoWgkGXCHiwnx
VFSF2L9O/CbYViHDdzAVMOGxr9CFcik/6JKHemLdarQruzyo45yOtwffWvE22LgC
2wGtHF1vKk8aI5/um3KisJqcJaA9a1gN/809yq9zGWZ1Rv9Cm3BD0Kzkng2hsKf8
w13oA9PaCNF8iKfEcO+PY6Jyg2u+lNOoiJOJhZniPt4KgGgPD+sWVziEAzsa9j6v
0r9h6GF+IKXLxVbx15xKWhlGx1az4+2VRKSupWfAELGu9Ntfnl5SjVYUzJZ9PQ+/
x37aphMjF4ynQn3gKncNGbg48rH/P5OWv1/pI50/jqRVjDJcntJXgWMNv5pdDQ1a
j0FHMX7HBTH+BuJxd90cXB3WRaxuDp8855RM33Gz9txjomIlyvWBmeKdNuQYdwKL
uMAAtynvEc2h7CiYtMc+S9TBfMcl9UlGoeo4m2DyDCOsSVaukJsjmQSnU/z6HmPB
3XUxQN8ruuKTPZMSQfqdzxQiCuOiMHDpMgg9Uq2E6jk7TS4kh82dFElbvPJ8LsnJ
p5Uyx6My4zc/TeKZvUHpg4qZbWld+vj5Tiu0k9fo+8QR0ArKCM3eUxdYDoCwp6II
7aTTcNiObNvOnIQ9MwQBubOX0H9nTSfBV6kJCgAl4MUpVo77TyYP3UXMLFeylVmE
U9RM5dq/hguZ3C5r2Yn3i0GD16OSPsXMIYdLfbVpelrpQcTt7k4KGW2KthmoOdSJ
q1wTxGUAr3caNdma1n2AuIjtLNB9eLG1NZ7atBYPfu1qJcJJVTreswccVjeBg/lr
DnjJqZiF2mxruSzfEWEAs0eXCiGgEONb6MscyYe3V2fQmG90m8LT/yCcjmgpGE17
7MNB1ig7WvW6pfLns4ABVIDIY4uAFY3aniFMKAkd7p5y77XXkTAYX6TzWO7Qscqc
z3USgLGCeSjQ3pQCxRjwccmHVwwFlmuaPXPLcfNTKBNx6hd/b/UiNaUOeKlEhThy
f8coWpQDBw6QQaqc8yn+cHTWm+za/2Ht78SKLBQyBkmaQ8HVuz7Db1SUihVzOPj0
FLwF/8197Uy7H7eseRWgfN8yvclrl958VzKuyj2Sa0pFLdPkDV9AzNzo8Ojjqwer
gu8+0b1dznwgXV7bh0D3OzqUMizLSVrx+V1LH53jElFSpXRmqjK3FG0+YKGeBEVc
a9MATdMMN9rTl5k42kdP6WmaXjOg34/VKUZkW+P5bYO1mP9sQAoIH6VIQegS5H24
lMNnEPQlTXXoV9HrGkD/soswFfdMCzqB0IWWe97Qk4WiwpyfO1wWKETXm7K4d5LZ
m4cTT3CRAjtQXqecweR3UvqRKVf077MfLC/0apUDH0GtRLeIXxxdn6rOQ3n7sPsV
1PYADzanEh48teN5bJKyqjFVoQIzbdnQ45Ey5Ya72MzSlUpY96GHAD8ACGdfbqlw
d0etUogIv3F8UAolWI50XTjfZppPgbLn6JdmMsIAANDxrFAMwFyzpkjvy572mYRB
DO8Rz72VRy9lDjUeBKCQzSbYO8X25I8fYfGHdQOZFm3ysrQqf9E3zjO79ZZAUdl+
2c+3lqGWyuM0406NGe7BlIYjmkLsIXgwOjUhYgCC4KWG8+DeeYupq8ZpS0kG1rhx
IR5xKrN1pWDHEGsQksbJgxEZKuu29QzhB62TsT6QTo68vcuHkM57tpt5/vg+HqZv
AHaFj6qAAjs8L/Nwf1ZJctL1yVl6wQpA4YE0TtNxLmwswi3OxxDiQudI58+XmHM5
wABp25pyurTh6Gt/k29h+EhYttKf1Tn2+nPPNBV9YNiBEADZccqA0Zv6+3oNQRsQ
f9ZuszJ6s/ezS1op0gnKKsDLtur+Ndtr8TlNEEaVFqnXpVif1TaoDRyxfCGMpxGw
TxtCJ4pbcU/y3lzkWDYldyv+3sAcalf/fPu6gJRywc5RjJKI1RzQHgg7Ce+MmXJI
OVz2KrYj/+zHKVKAiXS6onu6xpxfXRGApEAs693z5O8ZYJUUjNe5Lqw/aA0tEwGS
ssNqKetlCKTPN7Jg1f59CkCI3w1D4Ovwr4yZIS6UM+ZZc6qewrVyiHIsid50ekFv
bbYHCfvEsmIozbeuVl7h1xgRoWw2UcHgSwgbYdgjkZdWX4BZtHztK0ZFEpeQz6QY
M8YroABjkDTL+/1io662vEgItGD3ZAp2LPJDGQT/TMdf3LYVS59Lf+eTjW7vc/wV
Izc+R6XGt2Z1gb/8xROHVNeku+dNFeRVtUa9zts/H11I2C7rz7GZU1IKKfFPAhj1
0a/kKvj6nuamBNYu/n8QJF6b2vVcUNd+dtfxYWkW8y45c/QXD00vsJb7R6FlBRLj
1larUnPvsQMVZLLgIXTTKP57/ANYbof2W/HNElEkQNsjCab1d4bgPSgy3PPuOgf/
s4H51mZvW/oWpk3KHUk9/+ggEmh2dy41iJlHwtj/eB0Vt5F27LwjJr2/xm0Blc96
R5KItIfYGmi4uCY0nVX+IC9xWppVdw3AcCnNpyERQxBIZFoV+CMtOcPamWkYomg8
cryEgT/C2rVhBAqCDd07qwhUgac7cp5Lb7ytYhpAZRlNQtqGM0FgZ/cTdY3ZETqR
xwYheNDqHhqudGJC/V+hpNHSVJ0hFzqV1b56QRSOpjElrkyOeAG+4wnNxA68WnD0
x1YLw5dK9Q981ZtJ+8gkLvY+G0F3DI6OvMPHNj+Az+6/qMdT7ms/sePJRmXz9gtA
9U7iFZtq4uPFEcHuPrxCCax/4vVX2hVRFpuydVjbZGSCFQpABduRcG6EilIMV4lw
HhjAs3LTd7jafQc5EMlxTeozEz6KkngglsPpZTd0If+1HoZaynQaJfuWjVhLTWsr
PYe9t7v5YGwZTH0Ye7peVJ29CKhE3WvLORMKMYt8CBSGXIbY1owbw9BPzkqLWDqC
jxhGhjdx4gMspMfNqGk6Ojtk1pgLxavaIs1bpHOGyxjl82CTcDy060ESNId8UegA
qHl/qmzKukXwnpCTlxEtOxVnjUk0skbYASMu02xdkB+u79H6BQSbLrlwTeI23igV
fDtpPDyAvIPbkZksgRxcVHR8eTHcUJCwPrGXzjSvh+NiKyKJbN9cbgVZXfVo7dOq
TrjrHmlvcP5lcnKjAuYueJFEaerZbuSPzMaXhUi5ylZptSf4MLyrReh9crd1YxzJ
zFFi0QDmHVXWDVjDcQyYr2q7zIOTGXeYQjmYwLwIwSVmBAMWlIqn/pHmlU3tpEP8
zDpbWsrtJqVYJMjRvqLFj85tnQipgAJE0SpFP6yqN1fATys2hIZstytOI2hiNWuY
Yx3afFfZ5RDNSn4W7xmi5hoNmOijdox3ThjDKbqeqR/WjsuwthfM4/Xmmjk0ofEC
OroTVwX1Vm9Btg+gJr9oO4e87ZH/Y1RHOYJcZL5OZEgyubmThXQ+th8PYFoPFIaF
G/AQQBnBRx5o/V4mPNZzTE9KlnxcUIIcOQvyXmuBqhjPyHqu+lKRt2fOnznOG3zC
NHXWzgOAzT1NZlaAm+OhwSdvKJFblECbMkuWp/9sANLRNJZ0BRlTEwDAwE9XRC2f
UqExEptZ8GdaesFRS3fpKLU6e6wEVULN+x2mWkK8lP6kCtzE0cfvKdYizuFYHppt
rV1vNhiEEfnajD8KBZ+FNJLiQkUUkXRUVPIv4eG6PpBX/hGfvTTW9YifkS+c+082
PsN43VU16QZGLkAlT2lqGpP4m8W+MYttIvYCZbQ3Qm0E3w1nMgS0NQH5o2pLGWj5
QB3+sniO2jyme6zlzdPWzTnLKw3g8JV/5jHDEIKjyF5vI2umYHW2cktZs1rp+3tJ
+VU9vRm6gk+pL5QJhP4t3j08JbB8TMf4fjZnfb3chdS2w+LWNtdmP4+N3G7oMt6L
5l23C1NOuKmGStAouPpnMlnw4D9dMWxyWhHJlc9557sCXcIHzgyO+xgU2NjazsGz
5DI2BwbQWD6jWRn1Qm+4or7Y+GrmZDp9kj+XVbXTo7zK0JvqkoyxdTOBDzgeyTbn
8e7hszdvcWEEg3uvsfDsjExUaJSWThMkglEKmagGHKv0soiMTZQFi/y6xt2p8GQb
nPfbBoiGAF5LeiqaIorxdIaGkfGxdaoc3NZ+2tAR62lC/KKqpWFnavB2/LiitmLb
eQb9tDdQ5tqBu1/XFvI9gNwTeMXRUNPAz+BzlIQeDIhGAAnV0tHmcTy+bStBUZ4P
zL3y/01Z0v39UdDCeTN4hHp+FEvqOpujZ6OhHWS4WngPh6alxmpfA2e9D/a4SIaX
43B2lMeq2rKtSvBKDpE9UZudeoWypg78Kql+LQoHGsllpcPrUkOz3fDFHvFlQyV1
2PZmR04ocYsBlsr8uUz3TnLU634R4uVzDkxjlp3CLIXa8t0Wud3K7uBey+O6FXYN
zqKGLSH3Y1v5BDUNsIJ8z46H+Rp4536cdq/x4iTxSM3EA6s+0Bl8NscI9yaSeTe9
lnFRXt0jvv+hesRfFM8Mb2E2KOYW3lpYtjXcaB17LmTNfcJoaapb8PZDxxY0fza5
T9WCxSV5/AE4amqbo5Pd01Pzwja2FQgxGoGLH8oL+5v+3azR+GZERE4SrIGL4gOw
ZOhhm6zMcWjO90LhcR3F/gy2sZc+Z8xnVRqF/udVl0dyy3g9o8nk9POAqjFB2cnQ
ggG4NvCo0f+SL9b5uK5BCb6flReETNZacQQNYHqVR+HApP0YMalR6h2sPHCxBDJX
6JPVQCy0RdmUODH3Sx2sn5aHTUTzogtxtgEij2b5WYyD+92flJAQ+jbzwISXfmIB
zAz24P5rKeS9RrDNJ4uDL9z/LKmLS3MFRCLqVt/+7vEmjbEnSfhfsYdj1rwojxQD
xernN394AUKefWvIUzmPJIuR8ivpI5V1myPavZikSUbb3gVz/F5KnDvtgJAhXvGl
5F5Uq3B+gvepIkOPH7mRdovlkiTJeKLNlUumf5o48SABV+GZbz+fpRIWa7Z7157x
Z60HEVhzOOFr0Qf+FoWL5rgLUScoFvapoLonXXFogYgIT+gr4EzpgFjlC2EH6Un6
dfMjrJ5PyB85FxGIYnPZ8HcEaG9o3mtwW94+UukK0A5i/9T9dnXXRoI5LSEGvjac
p8xTcLKoNNnf9mRxOtszHRxX4q45orMToiyt7nQJ7jQTrCdkaoatM2VxugVbhfZp
GklbrJ/mIpzCYILFoe4uC0/z137eUNisxdBOjiH0kMEAYVd74sW2qfg87+m/fDbk
XZVKLiVbDOEjA1LZ3asZ7x0iAgnACVlFS1mKFvDuXIpgdK3oZaFouPd1sJOVQPMH
+AJlI4AeL6qA9wt4G7SnWpSOy5xWcjzt/A+1Q5BC4nIrMZS8tCPT6E4ZPJupw6Ps
WUhBmuQ2zux5CGSdXttV0QE5W1bjupoHG/CN1oZGtZdNrm9OEx2kEpvhSigZBgtQ
X46fKKzn8sQGIPTpSaHy4lcFHueXNZmVhtHfLV5Am+zALlJNjDMcV7Bmp45Iihct
kaYJICjaqkuk86De3WGmsUrpwKTECy8ToFcm2lDOa94Y3d3k2IIC3ui/FGWFuESf
Pi0CnyuUrakmbNCgEXKWVmpRsmxcKLgRIboFKe3YVxSN0bvMHh4GzwiIhpI18Jap
7sKwzNtVgm2p3kAA693t/jbG0D3UXvUs0JZFuTlW6rAuOvbnuHJdPhBRmO5IwPak
z8V2qxRm1rq6xteFWibfRMk2gZdIyBY62eosjvPscDHKsdvfas+EVPqPyaxdUohq
1dnRHEdFybDMFhQGmy0cQb3dguJxArY9kVbUXPm+h+R0wuewE467zBHff3oujhm4
a54vu8iSe0c9EYbXiR3DbFz7u7C9HDsZRcdK6FOmCtYYxWHzNsm3pnf74y+HW7nO
zmZd8XTiUwdRRlpSeT1RbV1w8vpRHyKbIMIRdpxBhSdMsd3n2DvfofgXhL07nAMJ
euRx9jFp3UDIUv4CpkCY9H2JIgZju8CjA5zoUhXhgxWD9kqJtC5A3xHteCrrNpSW
bbcMEw3hhvP8Lt5i2/CJFoSYKfnSczjXI4+1bxC4J7l/xpAeE2XiCOoV7gnY3jpA
BzEkE2x7zEbO/32SCWRlBufpMY9Vfk6vsH5GLqx6OwpiuwElASlprTkzwk1v06Ut
Ij+VtD+VaZt0Ncx2qTebDrrL2WU/k9n05VcRpizDwofbt+fwrvlN33UwFGhhXVgd
G83YOzIqdWR5ek8Dxv5SsH+0TAnrerRPvv3mrNKzJKEpjgDt1LWPWqHm+ewMceA+
5hGtJeTIPlUCtNhaVlcwp1yInRTOM415rWfbAWoyM9T+dNcyVr9ZI6lssGbB2kBS
x2PbfnG2TrvG10Bt1WxJJTJcZkLOvMGKAJ3VKrvvrtyM0gGz172TrWPB5Bj5XKfu
Wd0jb0JfgGUps8G88dSvk1qoSXEYjMVQ9csxw32H6FyZaIvkDmU48aXK9gH5Isy8
faAm60GZRrOafJd9XZb2gvkruGa8I+sq3IErafi8ptQQHxSVRjh0Nan2OW+lDOFv
SeE0UU+fIjDW3UuY2ls03GuPeKsQqny+xfLHAlzVMduZAvZv2Tv6xPSXmKi/AYSa
32BX2pHvIQE4mLbgwH1mjWayMGS8LsysWWu7wlvkmAR4vUHcErZHenp9HVaKz4gB
eGIKsPSLB2KzV2tZHrYD1AKpyg+Co2IlI7Q76hP25XB39JmJjBoKjttAbYoZWPxk
rc7AKZZNr4X3f9y/D19QaRXkrC9RV/9ChzHm+5nHTz/rtwk8XssL0gzzxYo5FOyT
gYgFKdxz7sgNI07owbGuZLYOlDIjYYpUPohYS2TXU37p7eAPBkCR5XuqwFTWpXSk
+yJvDCiUyETE1LBOJdxv1xXYb63WaE+aztuswa39jVMVboce5tAMq5N8eXZIjbd1
vgx9vFXnOrFDVPWdev03QkvYei+x07/e25ew/OnOo0dWdBRjUa8E7/0y1h11MkiD
z2lWrSQPSGJw/XuxlXLKyeW+toVQQ7Z/kFzZDCm33XBjcG0LHW9KYw4hQYUuiysK
UD/JVkfhm0kpIQe8BJ8pnK/7XhJKZGWLsbOocMj7Gl5EOWzAU1rXtEceJjoOsdZe
Gluun4Wkxxc1VxVL3qJ1GNPmCFKeILYiKZeBKYlEidHSikUtIQqa1H1lOdb4cdcy
kSvii/VMqmwfTkcArj2POSXDejWhuca7qfhzbFMVsp1nfvbk77bJR3DXtSka0ebA
JTJuMZgYQEt+adNzi/1NmV/+VupfuR4s4LQuuC6GI1S5wcw/zkRyQIaTjJs5w45Y
o/M/2Z6Jye3BsGljcKt40IQ6P0F1+fBEkSaLZYOgcN6wOld8iE3a0rK8xkpKIo/b
4cKudAxfwE2PLVuL27TPxAcBbx9tgmpfcqKoV+o27+BVKvl0M7cdwnDC38tnIUAz
vWJsbYtDFVLP7SbbRK2cltzPkKz53c74lYHLXUo9uuLkJTuql3vyoajahAIogn61
wspfXgKbi10908HtyDwc+f2X7hHnssfUcXAWkL6SAwObdy2CQNueX646dQR/2Ggx
IxnRDH0fkkCkTsIGdsHZYirHVx1+gLYUUv5+8xHi32dv3VB6bC9la/IJqBR0Humm
aqz/fuD9cCvD7hNx7ajPCLy6NFPV8iuWLehpE1EvVb9ZOwqwRJZTqi3mALQgR77r
9nfZP1MgX0pGm9TNoH2/GVpxVmp+nxVrB204VTPa4RHGZP3yCmY3JorePM39C7sY
5HuM/evBVJ+MqOK9OYOp8ReQu5ji1tyysIogT/rMnD+hH81L4Rfmn9Gotp+lEY6o
68bBXhVCdCiIvkFwelYZvtXcCStaLgFsFEuucsyWl6++4qqmpbn8wpbF2Vv7I9sg
E3QBmnYrC4HIT7wH1qQdXXtJX3TNuV4GwIu5m2jppxZuQaLnwZre5ghkFdx1bLzM
LyeO+Ar9IbdezxpCJDXjuPe3v8fouINKmntRAYMLstGu6M1QsMw8SNcfHcNjfc+0
NUEdJLUylJGFFPOTLxs+xbReb5wlRxWqfpfqB/sTovqeyMWzY84z7TYAGcHZm5MX
BLBgs7Yt4zRq+2BnhB/aSXzRNP0Zcpuy8nCSymIsL9F34WlD27j0rcjp0hJvOj/T
KaAVPcliiT0Zn3kS85HevQ3boVqGwDEud1YvyrB30maUJ8q5TQLqAqSmdMp4d/Pt
O4PyISzZp/Bn0jb7nOjBmuPrlQ3HArMR9TQM1BXXKLdTpz1hmq0S8Rl4qOhauJc1
2j7/H/47hRWX6wM5azW8ea+0ELklks39BcyeNkOLdU7HENAvH3K8wpDZtQdqs57z
paXO5C48w4Rytu1o0G12c4/Zl5YL+xEISDh2kwa4b2VKBZoR/Wn6yev4e2L+h0ok
zN+Uo3WCO/itv2dPUJs4an+KLRVLOwAZxVXMNagbF6eYhMNBqXje11qatxWgIgyX
0fAMJDOzu8YJXoyHCYqRVnSDtXfXDOyxu9Gb+QilTocvNGr4lF7UDhOpELsDxkse
Bchc+E7qEd6f0bWSNrtygTZpcUIhQmXuXYz1k2/VJEZR2kYerVPg9lNCNIjA02nT
MJRF9V7naVMDKL4knHwO58pQdDCxniW3MXsw5U1cPttAkxJDsn7+8Cn6mISZDyWe
Wl1eVX5xfN8GaL+iVaOzm8ao9XhUNPbSvHoYKIHP9azSMXEONBCzF7EJ2q18sSSr
p1T/Bp2nBIKIQw8gzK5nnTr76w4uPCtewmMtFO/wxslMaFuGJj03n2N79vqejFj8
zLAh2jy+brCxA1kK1YVf3SE6XEZFSw0PnvaZywiBRCoPUIiim59DkuDYD1pCiBjG
o5fFzNTgnRgED+SLfbjpAr2jP4eF6XHKul4CXXQwWXaQFGiw4t7qkXdefROsadC5
cCI7bXiblfFkNZPD9wd1NNU5p+LqPxfR0RuoN7IcARCTPRURusyWji3VtCZnf3SD
GxtO/5rw2l5R/vLy5ie5ZZDXPbVxgO9le+Y9CkmHqG0ey74U2F5WTIvsoyqapP4j
mUkVPXOCz0i2df3xXhfoLUBbHVYV+FHDEwwuusRknr8azcl8qOmRTqrTUzz59yIE
dx+9h69S7DpxvVsiR4aDaiaAlN2ZvFF5WAXq+eQsh1oQby81rQTqZJxSliDP47sj
RA8lB9HTvZtrjev2+B3rP1xrhEM/7vuEJRIZIlHrUO5yDai0qxUlNUlCgthVoiLs
FMd7klOVaViGtmwDnftzeKpTzAi6F7jdzdiqvqvMNujXJHmO7+vtHW4ceS3tJjRK
PTGtsHJyKpn23FQTLADJ4nM/5m7hFjMLSf1Yv7zPXxziFmHxzWF7fT7r1HozM9FY
qCTgnEZAK1iwOkexWxrHnherGAfQAhky6TVk6c2o44LEpaM+5g40ZxUB0o6pCBsI
niIf9EKPElBFWRlSLELkfuh3W0kwUEa3AiODpe6noaHPhjej0Fu8bH5VKF/Sc349
jbM8W9MMELpsJIiW6Ra/56l7yRpsRw08zXbux3O/PSMj1uaoZ83c8vVy8+ya4SAv
GfHTsPYgbQtZNX58FII+Bu0P+G1O8AE5fOko6Ai0q8ErsfVe9lv0nulSytKGVPM2
tE+3pizRUldXu4gyAO3d1YSL/ADGlf68eFHqB6/VvNWq8Cwz8Ud9Tu2+1s8SDOb7
PmA+/Yt87007ibRTOM5XJkkKQo3o17qWgVDpR+YjBB3ugYmZ6R57YGR8+nUQFOto
NsfdEAl/EntPhmewVsTQDIUtUmDrRHu/976xmQigsQ4gxw+jouK7iJDzr2GhBrvK
IaSp+O17ztA/mrOHe/rxPV6BO/QWrMQQzZfX+Rd9+UR0l96X6Kf2B675Kfe2MXr6
FA3m0ZaABU3rJY/aDjVIth2dcm3mA3Gyc00ifx4mzA5d1YyGVhKewgPB/unzOSMR
SbsVkV7c3OJqzfAkJ6oN2fCMWSH8yu9resJy6gBq51P/WWoKO99LmLuLHCAtQTOE
do/JIdW1EFdH/Us9gLrPA8jkP+TeCY4+GNW07dsSNH5KXh4orQOfaPdA4ogQtyDe
aVFFVka6aZZEdlXNOcyLQbAdEcuI6q+OK0qYRvYzP1VEDDwhm3M7Um5N65NLcfJh
zW+cOg7EDHJ2UJWa4fDJFZlnPRzqfI3QO12hms3gmhl/DGWBe0Wql7pKZf7v4CsB
ZeLkv6N8U3iZJtha4i7lvIW+hyQ0AB1yCz6Ew66OjLCPo6si7K3+EzWVhyd2jNq+
TS90hC7fT4YuArFoDkmj0qUS9/vuaYphZIRU9RijC2V4yemTBgbzSlM4BAxswpOD
crRqZ8+hkMUrFR5MatE2WfbprVRpoqryli4410xCYlRXP91YXZI88DI3WER5+Yg/
RbrpdpD+lWXICdq5IQvWpgTHu4XgpztSORdxWPsJTJmTgeSTAivzLahxxJOUaAts
qd+F0GEWkiYIQ14pSjT2VnrWYS/RggCbsY/JKa2QUHjzrUwRajU3ztI1UXPTPVtg
+sjVIAdd87oh+T+u8Mas8yfFPURoNHaHVZm/5/aEpOlBrTCtW3JemsDdSdnfXnjX
klWnJ9j9b1UQGCXwaAQAYyN9yd7z+9MxBtvIls1+6KiDTFuRJwdMpqDQKfcx+748
wvVSfPZyQgvIfz2k2Pkdu5g3ZEherHON0EWeD6mCbxqjFKy/8SkEt6I1/LNJTKPt
5WUdprDqMMs7MqMoaE16w/mOmCL/rj/g90jpLicTo2EB5wYCon1ImzUbL7yYXoPP
RcjfErJ4FXfH87Tmv8TOXPfEKE9twB2OXLHsAzifGSlDt+TIixts0xU+wPFdtlF3
l8Rlc0+3eD27S2gYMr12qg2UmmK0LXeaW+p9Rl63rQpgTpwbCjixb1EFshH3DvcL
rUrl/haBMKWjI8ikUomJ3oYI92ShSYUf4FO8IAtmlfBhc+Zf6HGuf2ZmnLHWxEQ0
G9wVteMayBcyA8l9F8S71TvdwkahJFdqg5QVwXPkHTcv0aEac0kR8fnAnRYs+NOO
XY3StUkpTsBOdZEopRwrqq/F8qCxwUVPmioH6mEOb55ju2W2EVsobuxI1FRiTBBt
0M3Cri6js97PjnOR4uxYPJa7GONo5RoDJeRL04UaiGQaDwqeYO/YkfziRpvKZNFF
KwG2nULLqGWBakFbNDhiNpgzlcPC0hYv/KrTX/hXMQ5zMsaEcDpp+v6J9C/fZ/eY
tAAlkyydJ1DPpOFLcKqf4wjV6dX9GcfSTlI5PfwmFCGsjeYic1rQ48KdQRiHZcnS
CemGsTOo9YD2J3WP33hP5gNCo0yyt4iZG4+UMhGcNaU9iwmELtF3fgLrdMQT3KOq
vI5H1URDwsy93rPrafISny5jI5sZbZwS7haSUu+LVWa191ZbLds2qcnAGomQ0Y4R
N0wqwDyn8EaQ4aRdUX/as68bb8sz+MBRLexd06X2oD+zGJC9jDxd5muFHFQ/ayOK
TGPQMEHT07KyQkhlXMZ1X9sNXrowUKbh3bzPta1tl8Vy/708JSK8u67Ijkftgawo
F54tGOsdDBlbk6PCXetEw2CnoS0K29gNDRQhXY6UwOD5A/AXGW/WLOb+9L8gMsaA
GlvRQKsPINsTUNvSXZIIHRCM37UD7TDQy/Y0DcOvhQaRVSpRsgYvoXYSUAgQkfcp
DON8yEv0bHEEI3wHKldv5gJxTb6EDUSbthK8dI9lhmxd/4sg8EijwXdtH0ShKVf1
lF69ZAFsNbqoCyeqSyAKLCXbuA/Z82M8s/oY4uKuAB/YYN6ttxvRlr4y/cnPBEij
28QYf7nWy5GNnOASi0Du309xxkRoABU4SQwOsG3JZVbnsTIs0oaD4otSkOciz9pP
51pkjtfhuGY933CLOlutzfwbvjmOJNEFmRI4b+7gDjy/unTYhUsQadeRWGSXpKsx
OO5zHM/QJuWeQbcmHTa5mnqgWZtNYFBhdoBqV3Ub6eJu9ffK4jD4JSWRiXoUoXuN
EQ9L4slhb1Juc7BopkJ10LW25afxFXZXt57KFmSFwYOG5u8kFXvZrmojxXuH6k/b
jSqN41NMCW7iI+ch5ICK9FDKK5Cc+QNJxLPvrzUS6xLLxLYOgKkmFyTsxEX+PhV9
SA/e6z+cVxZvW87iTufpFBwcEHkiXs5SwM9N2QcIh3jSejkGWKWbD8fiy3zBL1dv
RZrMGxVHSujcY+njoV5h/wq9NUp7WtYGLcuHNo+oBuZqriyxXjCKs0p+ry+ublGW
uyjDAIWEP88JDtAXhStDJWjIvo3PlK+CJUE81uSTfZXSrpYs35bAkIrMtA3qcYJ9
2qi78kmWFSMi/eH7BXEwFX42fdN4Lu3+H0mBEUHMPyc5qFvuStg9PJoPqH/2PuCA
+FukwK0AuYEQ3dYImQoDDD6eC9WPTlGkqdf1QiRF3XKmHiuJlSLc4GVkem181bTF
i8NaP89AHfoUvivsx00rDJwLdlmipy4uYJyF4rlKMlMbVNws3EMVGU0R4Seo1hzP
s0fTj3xb0qAQORPPOoNRzTKyGlASQPxXtj5WteiyQm1/JESB3CL5TYHnMr5YQNrZ
Buj2Ti7VbhIrL06ozulWTkGw+7EWv5YvLidsEv07EmX9xhIrYL7IYxht62ve9S+u
Ki7pJ7k1QUA0VEFDI00Ln9N9ep457HiUq/fctd/YMbJPyfh3YcHZ41W6nWqSHf0Z
2gmC5PnfJtHudiwvv60z62DXpgaJXQpo6xqgTNIf1CIKQC8i8UaAIFQlmBI4m3Vm
C0X70rxEV1ucIPAxdVxgihiBDdw6qyvR2KLh3a7JHG9qKeo/DChrGyFFFbvr8o+n
VqQS50WeQa17Hz0XyGZvf99rKbfBco5/mHnibhs0wCO82zUzrap4s+VNeOQ0BWBV
cGanIDrdCn3reae+oxACWXPxN9mHi2QgCAXDJV/1ao0JuZwrE7lgOPHiwei1IgRB
naFL3e5vAzetPlupMS9jSUuo7AEvBNLUzPFWKiuDNqU9VtfYLlBrMjeob/kxTJtQ
0vsQjX7E2ywK92Gxl6a+2bEfIIBPZPTax5Y5O/cxQASl7Lzo9HFnYW7D0pGlDNHW
e/NX+znvtNR+fh41FBcgpSskfKsedgnzZEYZh2HW2jI2ZHR8Pn6+/vxIstEnv29Z
95SnApr2NFzPTckVLdo6f9c1Z4qy52dGu1/5ImBGYqykfzNZUiR3vxoUeXYBeNRO
WDqKDt5NNraq86Sva40JdK6h4aemjW/YYqOp5YUi2agwzRSVzMp4gFuDGY9TI1gR
XeeGJSUbeLBNglJN7C8M/YwHwQ9yVfgu/8zONkQfMIimOli9Ns1wH+Co2BFU7sH6
6O4hb9E7bexJGfuksmSkh/bzcAgmB0IB+aw+70mhUp+l5o8zPoHGJSPskuIepoDn
mavxdW+oZOP2AZhNbZxKDMHoKMWQbMRDaNWWL/r9AWwOe8rMDoHRfrGFygHMbAAF
gTi51M+buHWkXF5DXilqRAJcJqXSooWPLATAZf4yRCJx7xjZEsIUI2uDhSqgOD7G
a5Qp/fQQAgVc0WX63Vxz5psrxG5HYL6CcsCSIiLUO5ZxYH6/QO/KeATJhpkWmyvb
K3Xot7N4xtqygdt2+tjVmRhm+rUj0RKJc8sY6X031HUSpZyhEWfmRwpfo8V990bE
OY904Jg3BvEGI6FgLYmnXGcVcvUyYHdGOgQLR95RRWuAS8Zn6+rRUj11CH3s9U4J
r4rpJGFR/zcBeDzksJrQTBUNuJUa4xC3goDJBFDuIsOtXR0V7petQxu3ze3oH7E8
yJy262ZLXY1OuWN42r196GwMt1tFWZjxPCo61ZuPDbL7VFRZnNKF8OSRm6l0n+8C
6NLXPtb4QEp+yoQHw3Fr4dTXf3QNLEPbjbz0b8miJu2jiLi1GwEjqKk+Xd+XboBh
OnrRTwIfUi7C0hYX9TVRJ1ffsZkTe9xACcFNUmvmu03Wca8F7PzDc18126caAXQG
EmulkeI2nn84dInGeNwl2nEb2QZJoH1WPFTg0M3ctzNqDOuo/p9MKSYVpRcJdOlD
8RZOpUm2Zju80Ay3OMJ4Ah8SBmyPRCNc/YqbxGM6o2KrhsXXNzgBGI0yAUd/yVd8
RwQ8Wi8Gcr0WfYnMwi61ktlKX9Kc8lCmVkGnZanZibudah2CBdxvXObzZDS18l1x
EI/NVYe0AD1U8gBENNz7Z56ZkNbcQlySnIu29xxdv5t2bjmQVP7y7s4+NGXTpbWB
pGgTxAW6OggxIP7FqlUQvYCR8GGBYJ0crTi4GZveuEW+xjaqfkO6/Nkj7cbHbMNX
GixCho+fIFWjBLD2hTzg8JuHCPKZ5zFkqMD5FdRrv5gu1teLH6dWpVLLqTP21g3/
LLt13UrQTLzVSPHe1S+2GvwFciqiv3eIT3Y6JwR2Ry4KWs28fyn/h9erV9E4XX6n
ywtmujod74SyOw/Jvnowu4JBCDZodwOFiBVhURV39nSbfSGRwT2233rGofWhEhsK
BfBE+nYtVDLStel17p56Bd3m7E7lsCVB553yp6v55v+MLJZcm0IP6PVAFrEHSCkS
85bZ28UY3LbaHu7SCuznTQL65Vfamj9w/2cnJWshM16Nw9cUKgR6IJTFpezpwZ32
d7X7nWllpAApcCT/PipirGgv7cEFJiD589dTRNa2cZonj7O0Kdrhb8vrIKDIcp68
KSbRaP3JaxyjEUdfbWZ0Qn2k+JkIddC25wVl6aP+wQ4BuzGH3JRBH+pTWTN8n81W
Ek1wLT4OIs6xC730MEpjwkpsZUrrVXhL/fcxA05S4FdeHz1aByMp2mG8XlyJ+dmt
TjhwkGRe2N6HDTiuC530R71ij5V+Ng+qAp0Ki7NU0hNei1aMbjY8VwCUIbH+HfP7
ol76oG+R05MLRkjtve5z/j6GPEYNOuvAE3GZRjUMcySEcunxU9b/antSU12XPdlM
wWMAqoHmPTPu/gsd86eam+G0gRLrGpFmgffkBwebZmsXsqhF2bZbdbNpB7Y6TMNP
FZuEIvAg7yFPX4t0yWEv4ytViTl5YSHS7Eh4qcNGWzs1nAoiyB7kVbeQ50DKgEDc
7msoi2tNK5uULofK9WLtirQmGUUy1cfKarWBWhtdj5517gsXPmdf5fMJ1YXWT6Vq
Rp6CxquGywsYvyS7b/KcpaT3XHv+GDCMBK8UflMnn0LpdCNYLNB+NyQXefMpOPVg
8Hu0zyD7rFWpg/8uXf0+evUoxQhXgtNR9hY2mFnMYJRX3vc/P4Z7Oc78sbVIzFMp
U9pjY6dsWth6YN0TMy/L/2EXvzMWBzMBgEvkZ4eIU9spS8Z6uD/bEwNxvAX2Ajgt
m97Imcxmsf/Oe2Qb/bmflvjsSwbo5byDTrrWTzBDJQ6d+/b3iLZMDGThhdmKI3Ia
SROhV7kCP2DmNC0CBg/QA5bQSDDRLC3gXTxZxftvBJL4KHHiNOsps6cdD2878eav
hD5tz8kciR+N1xLVABhmj3Rys8zDac+Erkq2ifQsM5NbUf0H9I2v6Iovhwyh9bTR
YWHrfAw1+Ba1OVTc1ERXlYjXUfRM+DwnY8vIyCe5kJuQGwaPoiKFyH4BAeyH4UIR
8NEBOhEeqEO4AdggLwLHkMV8faqZgsDPJCcZe0qKJ288y2dBsnpcKqdf3ZmlQ7gf
Pnfrh7puhywhf6v/HUZU9f5njC2gawIX13d0+NFyAXPBnvwUir1P1TTdrYraDqfs
VD5ezeulGAVZFitnryn3GNuTjydOOM1Uwwvyt9/XQ3xSMaCdj5sQjOUQinfBMgCg
n4KsrJrHEqLl8h5bLEmGB5tTNG1d1lC4s1dKCxGdbm1buyvYeVjnliTeVB6vejiG
oJa0NlS/5VMpothkrj4OPMXAfMBwtm0oQdUpk2Q2Np8fRIT4r7qdnZ27ENi/A9b1
feF9xRUKcGvvZmYzhzfNhX0oWYO8MhBby4qMYMBxyKEgqKLJ5jS3aI6Kbrk1Daea
KR3KxptQ3FzcwmlS45Fzz9hJHp/vidDQjOqpGjtTvkbeZeLiwr3tDTCjkLSaz75A
XXKUZIowyObeYZi3Fkw5xi2yKW2/dhjKWpopXjMxeYMGZQjvvrRNUF3xQNv9n4Ho
ZHUmOQocapZR6o5rV24vzrCaZQma7T5q0gAjYCO5FVL8gjIB1vFCmH9ME2ZD+mLr
RPllLONAaDokLRz1WlH+DEyttzprrGYjltFxCtRlY7TTGXWBE2gL4NJSX3sW7O5g
QPlWFf4L6R8Xatz7L+F9IcIS1p3SjZ6ZEswICzNZ5PxbsRLp2JV31z4QPbNzZkMI
pkpytsHo5xIdbzfNABAcZOe7b+GROHx58nqo9X0YwnGo+zHUEbbewk3/HjfunDTB
vNvB1++dgMBWazXYdPdY39PbH+Iv9HPf5zuNcENqw3o1CWS8OTDYpo4RGhB4FgW4
OP4q/pcDaG4VBS90U87gWgg0WycQh53G6YRAuxDs3kCZmQgY6R4XTML2/1MDPrfU
HUUakbYHox4DAdTqEKlU+r5eE/7QitTTOWe+Lgfru/3nSWnQMQuslCiwWHyJyYtL
jvttPbX5qu4aL3pm+3UwM3cxc+x8PSimn89yYRHcDxPzPNWFNJAZjMFM2lJ01jx9
ygSlUA/mgVHEsyvX55Cl3E+kyFXHHm0fpr05/jnpkuq5yihJw+lgrAe+x97TrDHS
saoMsAAo3zxBF4DtaUzxD02tj60lgiDifrfg/oZoIGcWCJtaaQi/w3sjMHsdyutC
PSy25WXbbVmHZjmwvUe8+drtLvfCsgzAjOO0Stkr8ICTTwjv79GMKFMY9q35HLvW
aexP3CoopSTUsLSJOuwkDlFrZMcWtk9ftCYbs0N3l2cMq/eN4MUV/3+RU4Ihrg4B
JEdffLSxlxfVBXQwE/DhgBHFncZqFcoMdJIw/rGKHsx4M2PLmv3xgnRMK/w53Fyk
EzfTYFgVrX2dqYTDvQ7CCfU1t3HcJbt7vOc0UDQXno8i2DfgfCziS0/+jVg/suxj
mmRGMzy3ZcIuP8WOHJIxDhs24q56BrGDh7yOrQUBlsXiU4e3NC7Sfx5ZEogNAFax
aswbl4D2FwFfaQSnuYvibdCZXpZP18EOulOoJlB0Izu77c5VWr6otYFB1Yoc43JM
Y+7L13z16jPQE6t4HK2yeZIdNoXS6ajXLY5SxAGEGho0CU7smzscUNe+Dex0U0+/
a43U5HkdE8gDAHGvKOn4/wBlQI8LG5ytRx1zrroFqUh7sV1/694LH9hfRRNCuppA
5aPi11ZukrjEv/7u3uEX18rD1Ny/X6/vTJzOAmNKc5v+nWMusdc3TteUedcFES8Q
MioCkon87/FAOO/pfANHd06Te4wgmzNiVbMv3ORn58jpB3KINz9fSQdM95+Hcmli
2OUovy7Ee8Pjx1lYNYdO2zifyfVgDFZ+fqomq6JDgD1DWlSV8ltCl+06YT3al3F2
Ai933GYHfDk5YyEWazb5dG6pkKev2O5s5CNd3nCd4tSBhnGMaphg7eOW/T0SrRWL
7/a/Y0p17XGJ+ZSz03BOpEIFtKyliw141WHxF00E6b3kDc5TmC4Lewb4nMAhk/4i
DMd1KAVMvUGAoOqR8l2AEkBuHaI9n3x1cSdxX5Kvb2NcBYZuD0qfTsOjotJD8gRM
b2bGjrH+atUw96mqxsqjiuLgbdSwFATimnnWC4J/b1cbMO/Kth1vaP5neW+6seYf
ae2F0oDBfL84kY0VIdIWRxBjMUyazd7UrHeRsFkrLyfjW23M4FLAMwLaiHv703A/
xZYyuW6EFLvFlaOOr6N1/v4Qv3B9szhDebZjl81T8qaq8RclpspzWxRtCPQtxw8D
3/XwEZtPZ7z776rdQ0LGZB3oD9D9eelR3QnFKu6NcLSp//wnlzdJoO6NXYe6AjOZ
ddSwvrLmVzXZMqpchAa7Cv2VkaK6YB5Ox3bmf5xQ8OwxFX36C1ojH1IwvuKumqW4
fuMPs9cxGZktvVVwx1Nh4ZYBom5+kJzNlnHz5jCSIRhtKZok2folX+76C6ZXwTDX
9ZEfpl5l4ueRz4GkMnbTCTtJOZFH48+XqQCXpmxSfcEUcLH63SbO6HhOJ3P2kvVc
YjpYjpaZPWswpkalgFNAiBHJwQ92a9Vi2+/vB9OvUl1Dxoci5oiidbGecnVppNB7
FaE5PaSpkOV8XK6qzMzac0H2fnFbw3Hx7sCoPYAFiy28sjctfnLTuq7j7HfXu5iX
APUTHW4uLBt3hNtVUpA8VxxSa+Wc/qEQKQbD0Kd+IjXPBTeA8XxR5u0UIhNvmMxO
HctqmTLsbYg4v0OLE/pPKkhQ3q53lTg7w7+mjjcEXVLeezdZSzHGBz4Lv9TvBRqh
tiOdN/3HHqbor/VPAH34MSPm+xk/f5214RvK7a5Ja5t1Cq5P1Y06E9CN9ZaZyUA0
AOGLkZRJ1r46e8gzEXgNahnYqkUcGOUuJFGMzkzmTdaEH6jLvOIvV+/vlf95FZRu
3lxWiWNOWymoax/7LAO2cmZmB8AP/Sf5+I6gw6ZXJyD1T++DD434FC5i6bR6a/Vs
LoATXE32APr9AMnMH25JLKuznJiWFNVVz7yuLizcmdCPVnyS/66Jcxs6EP71qiBM
rjLtZ/H/0avF9ZGtt+1/lqiQnJ76DJjyO3ivWrNtOC/am8g8j7Zo0FgnGQEMkSJm
0sVoG2VaTsHiZ+tADaP046WMzkEEpf1mg/WmXlPuoYVm+xire7uW2XrfDSfXin2e
2LgQBC9zQ0sPRJ16mGErXLWGO3wQcgdzP6OBCbOcyB+JhcYJc8ldDT9ObKNoUVBg
cifm+r7lamOlUj/miyrm2B61Qo8ZmWweU1xy5FofTWQe4qn8WbeqC7ZxEHe1Id5I
Tt3jTGArQF5ZMhz3elF9A2In6unl90pQUzmFhRN/ZwI7r5JsL8q+IZUT3JI3se+E
uxJkt6hUwD1FTbakC/3QAHiKRMptuW+ZVWXwLD4kN/ze5/ZXvEOvc+KkmtYV6jcN
mSerf4g+SXEKvwM17WV+2Nl0K/dLIcqsTFt9CxIZeRsEh/dEVwp/+0JHL0D1Wqx6
b1zwqqfRWAou+rEc2j/4eEht4ed/WsepUdeQMBBWStSsIM452sU/60Ttx+lsyMfj
OxUHPoEy/tneJr2mpdP2fwbtqpRdjwgd0eNfqTcymCI2ptJ0P057y/WgQvQ24EAT
PNHHV7VO/0QI0I3tzH7ERLY+YcT/PopsuYpXC/KOIjqWmzZcvOV7apxtrkD3BMXb
VbgvNuDDjkQdvD7L7DxPGKEJMvE6p42q8vnZJwFq27kZ4jnzGup0JciDpV7pJG8O
zlkQ+r/PR0nv0mUKbkOs1nx55lYrB7/0/TjRfSheR3gT0zFBLNepd7iJXS8y/vtO
9/DN6YWmN5CmrHzq+ZC+IT05yjlAMEE4VXEyzbOlFSA+68WGhGqfsfC2qpqEiAbh
y/X66eV55yjY64MUov44rOyYrXCnDt1sWn1l1Dgk9ATLKQkvhrEWhsBPxtcQ7F5x
6hXZNHv6TU7SgtiarPxNqa4hRfu849B8aiG56bxIwGID0Rnps16oFIvj/mYP8wAW
vx+AQ/CVjuqnQbqwnSubyPPoKjq/CnI4PxWX+1ZfDeC5mkyaZeLQJ1YTg5vVSBpp
VQFNu8RQm0CSWannV053X0uEvfLGZrzn1K6QC2LlK0lYgHRql30iK/Kmje7OuMo9
p1OZbPPCuRvg8CcTgAL6Nqu0uXCfTAzWlSzCkctO0Oiq6SoRYj/RUNW3j3tyYSLO
ElRo/805/FdKe/DtVCmYEC1zkPpy1xi3fA2GsJfo3q6k5eBPRBraYQkuQ1IJf8EV
1ZKGahKhrT72hYKtForohdJ6ezmjWcF++WWwXYpJUfeCGhIesIh9ywYpmuTadKdu
jVjpppR587HMuTrPja04rX/FWhYR+NLeB+wVelBaH2WeKWl/luEzvRNIz9TOVXx4
mc1Uq49HSzBZZRRr+ki4WtkF/jM3Ff4gcKsVzN/eZof9ycK9AIDrr4pIPmmp0OyH
enGc+lF8u1RXB9OBBODs1XCyDp/YI8cQydpkli9jfYsNJ7AaKlgcWXjDI4kg2D5X
Or+U/+LjF0YzNU8+YNbUt1SHGlB/nbnFXES9C0xUyvbbXaW0Uf16taVeSeMqNmIU
rwu6ak2OWTqH9+27/0wlDa5LUdWQwfgUxTR6B4No1w5fGpbU5UtXEB24tQq7RfOw
RBL/b0M5Nop86IstzeTXkysYsc+JpMfIYEo3vq7LUkmjM2fzx5KJG6Z56n1G0t0S
4/+yo/imF1HUKrGaeewS6xMOPB+RnEtICFxJVI+Ti1ys3mcOI/Vboy4iF3WjDE5X
KQERgNNKi6Xb8r4Au19/lB29jVndObgwm42jcFElQ/Z48Tz4qccIuBH+YJe9tGJd
ASJWfEPjOdQabf555KQgsOz9TCOPjUj8Pwx6KkVwcdJ3W0ONWWEppWWjlvzKzLVd
DOFrzBoI7Ulb5JGNEJHtyY7J8b0USJucSabisAbfzwuM8h+/4zWU7HHvWVS6MNAn
xyj3Go7MeG5K2u63AbeXyuPYSRVvOXH1fkhAcV7bsjXPCMsZQ1w7Z6D/oY3RiMJT
6npOG0ZuKrTeidVpx4khIm3HW1oGOnY4f+wBA12Yvbqi8/EgHxZ2/nMXpSiVPyJr
k3dYOzWjyEneNe4mva/wlPeb1i49BSXwfJ9ZmIApDL6yIUMuFLb4yb0ZOtxuK23S
mfODcSc2Uvc7DuQEJhJhdzsuYZKkWixZLo3VAHYS7Lj7fPLpgpGtT+wCMzI3/5ko
+Bvr+mbATL03XgdYGNpBiDkk8nAdbBEpmjweIgG1eoIWrKnosJAfkw5ioHhgVuvI
qCFFiJBBoh6ui6GIVIEIEIjMeJRLwTz7Is9J0TwcV67chww/YLhnewjABaqN3cSi
1gEd7zBScIlwm5Ld2DJz/E+LDt5ARukzPDB5bi3z7ugDUrSBOEm49Khr9qE4N5Sm
i0hK/XgrNMWkQMIqMjueD+QXTUy4TVXLKvhLXwqGaqLLhGEa/cNj26WO7CfRZcxx
xsjGl8+qSVaJRI8PAKua0C5rvz/6MEdzEjjFLS4TnKfPwy4WIr3Rf5S5iETipNVn
+q6uqPiGZRZQJdIoif7Dj388uE/TPU+1CTsW29dcSqndo1h9PNPLsEYzeE/yun01
Ns6HNo1Wh/+ufuZLNkD48N2AIplREVpGTebgqD3HEGTWfFljlg+wQJUwH/phJcFY
KgAun5q8KzLGNwtG7D0DP+yNGv3LQkN6ZTollTPD4MrYLScED9AqNp4c6MtlcpAc
qhM1Rc4tcg051OQe20MHq34ADoSpR82EMnZ4SV2H2uaXuMibW416pkD4fkwqEtV5
+82ecodG++N9gKjLEWiA/wXDsMg07kAoKpOPj8ygPLbglo/bi2ZVa637g0I+GwDf
5n/OjQYT8wqOKq/ud9XxMNHFKkyJeIUSoq4m/xK5eTCndVni4OjjnS5xlEda2dI5
/mjtDDmQfcuMWhFsxPJBaEq3Jxn4W0sYcPqdi7GWK/FfgThXeCb6bn7KsVg/DKy/
7R8hNyZNNU+v2fUJgSPM3s0GKoP8+kpRFmunDDm4dn3wSuLPRnZIuV52e0hQDpu3
14AIqYuSpKOlVMdwDAcFG+CIdNm/00fUjI9XZ+6mzb8jtTqC7fXyakDAU/Bkt9tW
5Yxr+iwHDAAFGG2JfFX9QVT/7y8bz28wynRw5KRnND7Ln9XA+tCFAQTxQd78LN5G
gEikQyTc2KAUoJ9u324IaVIW4mimP4egA9mhi8U7OaIQNmpP0FZXkyc9TSvv7GM3
f+f+RCNJRhX8h1fWszszk3lkniRJH2i11XJUWnnpNqckqhgNHUF3r4nef1KLiXwr
l39uXkLXH6QEPOVWDEk7mKscXOOivTeTmLhEWjmCyEh5sdjAO7GF5OS88My65Gcz
n2CNNkpzaQZqZ+SnrzFRCb3VYtYDOfiJ+1xeMfLTBJp8e7KeqM6jx+GsjX19v0bP
nMksuh/b/VmJtNMhWGsZkSZRhUsrBliG527l7oeCx/7j7AoL4QEQdiaZg9VosUZm
ygJC68759q6ASmvSihD8WxR7kO28Z+2uS4akoA8HAooQlFCB4wBO5OqSJIHiXDWC
ulx4uYARvAZexDLCtbUlYhVdrCCxKz6PNmJYSMOd49d6NwSQNnf38xE7sJlwNJ1Z
NOe9gg9qSXlBtYtIJ59bPAVlWcJV4s/NENpH2v0hSdiNE+XMXivGD4pUufz82czX
4cC0t8kF0D5+KjMkr19LnmMUG3+fY56yNC+N6Kqh5lZYS1T0rzdKVQd5D5ENSea9
h+UgSJC3bad3E2dq7ljIfdtEEw2PMbWyBrX9Z3kQwduvcAhNfWBKwDbThygZ9c7k
mFVBOk95yAl5krj8GuKb8Bp3hUpoX/xsOShip92VKYJkrcbeI6cj08XqRnGJ/yyV
qe6vvJmcJLzpx+dbKvYp43bwX479PcMtkKQ6774t4mjvchL3NPrFg2pzdhx4YtiV
eKPoDJ6PiX4rxkyZCwLqgJEBC0jKYtQqC48wKwe/y06Nhu9SsUuRXHs9Sp5UM5ps
cb8cGgKwIpxR4MYoyVB7yaKfy15NfVsS/1To9VibsSYRovqSEn4yBNSN73FdUbU6
e0fhU4xBKg0FDfw/qRYRGwQ0+YAyTnNIqdywehnEWJXgP9uf+PPK2Qo4EixLFkGQ
VdTXEDt3Ytcpg+hR8lhWjfrMj6r7sOHiAaZB7YYVhJZEmW0D0rlt2HsqtTbUz0j5
UN4cZdfEY2a5TnFcOSarVHKDn5iEvbOL8wOdB7canRbMOdVrzeIJnCv/7Lr9hVDa
sV4IW96WnheMNNNxedjgCwS3ID+kRSdVkHER90rzVrZkj1zIqRUKEwMzsNaDKIMb
l0GED+6GLJhWDwJSFGhDKNgLcYO9rfpgp84alRN9mvlDcr/i6d0mgsZyfj8HQqKf
eGeRDmZ7EM3dViq0+opiEngFNmxdZOj+4GuDX2f7JsaPhZKrGExj+1c82jkfDE0l
rCFF0lZxkbB0OTsatITlsyZ8TEa3gipFuxAANtaEQJ8aLsbFMcRZkjX9qaAcU06q
1xBTHuhX/6E1h2O/obDEkL7tIgiDHD7/+2Nv6jQ59kWSSHaBunm4OEeigeerypp8
PsJ3z8RoerV2o/q4n+/lJqlVi+I1HyiP8IpgXKFCkSKbjHmMpg0vgtXs6PwWlkuD
2EyK+URE2auk6kb9C4MPPhsOkwllvDuDR3qTHJW+pQO0ww6ULLvRBcQ7VVdmP1oz
CZwKdwWZSP3yvtKEgyYLC7YEVZvffQMsuQ49koJXfj07Xu5KnoJN0nagdOK5Xx/L
AI77K8LGasCeZ9wA56EyTDHd8NBYZsTvxH1zoOBDKUQ6nKQrmDnQfzapz9e1FtQR
cOmUAICTVvqV2x7MXhXCTKrS1w0ZeCphj5tEyUHPOutHZdhzhbzsvdtO03Mx7to1
umZWrKrhBcmsj1K7Eded/WbkTzhCN3834iTQbYGWht7kACZAtzohz+1PhrvXNypw
p5f9tKMyx0UCB9GsYKaP3aIOeo8+tMGeQ7Auqu3IiYvKY6o/F6NwwxOXFUFrU7F7
jEtPI8630dg9Ai7SHg8cIR0h1pW0INlBkzU+FeeMo3kLmByDlfwrPpSfxlBay1QO
+wAIp8KT9zhlWUU9fScsIOvRpnaHrDIvXuiN3CvkDZT6s6gZSIP+qaWnrWsWEirZ
HSAQc2jELUZ0pp8yEAjXpLZXXpRofS18uwwo6IAjibH5AMqUHjKrq3GWGDpmNg/N
w2H5ThbyLm5vJtq1dKu+EBh+dSmIHToIVOt5vMMpFl4R2wSRKhzudsbGSAnyG1pI
wvdeQd04BwM75dMP4NUTBakr8cJozXQGnyDJbm8N9CF5jam6W1TIN/Xh1LS1+ZNi
G6eOdkCgc6ZRNY303TEgTF/7Gy7M58zznknXQ4/oF2ixMEei/kmByJzlUNTFLYYu
eQWaJsbpv/LF+x4Tar9YXiInrHwsMY86jsOwOotOAKdc3iye2Z0OeMtxFBIhC4AL
TuYkpHSjpZ21oyFWSR9+eWVgBaYHp0b24IC/Rxmgh7zvPggvMQihbltfRbYB5ofd
laDpJevccyIvh7AidR+d5zU+n/pawJeIjiCl+1iiGTwfEWbmQfttlYgFuiQFrUvi
fGaQHWjkk+bqjbEMjufGAApmKCm6VoW2NWIdMV53+HxfkW3zVNSLVgdDLLDPhdde
Qpowdq0wcZmlOdS6wYpC4fEecbbVuj3YnxOU5wyJFbza1i55DhfPXYaOZrTjBFs3
NONgwe+sg74Dpwl1QmDM1P9KlGtXUv9VZrovRmoTlzptLpb+f8NlGJ7XVQGiOSUa
Ih84iYXA8p01xyhGYPvH7lFfgg6PdKZmkiWVo8aCjnvDOuDL1zyDsFpnqyhUELfa
JnolR854+GL1ioHfbauGSaNMwIArYAmnY6Y9umYSKuafpgHGcV6+IDDaiQ2jG8yb
6FI5OEQfoHRtpTFb+W77BQ0+5QRYVztB0UlFvYBsbvtAW5Ho0x8n9mq1tJ/rc7M1
32VQRm9ISLkLbWid1HWPrCyCwReghIQExaC7US4N3+OdgjVD2ALAq/t3z2kMyzDe
qI8T+8Es9RUvSppJNkQWcc0TpocLQW7sKRL2hcBZ5hQ/ckaWQ8UACWwecHuUMmQv
KbtOijpaKrQM/YiRib4wpkzrWCwRJKpDSokCt7KFMCqnAi+u3WDM3yLSLRyjzDvl
ds54ElzMDF4Rj3++cBBZj/m2ruBMkvcKWAB0k52v4e/+AXLE3jc2SzTUC5r+K4Hg
LGnDLNkZgC0AO/NOv6lfsb4B7/9rf6TQQIRpyRoUYAi6R4RqRiTSjlm04WOmTyNl
tUUzVArIC7PUgpDsa/LZur2lL3aZ8zJMPW3hSlueGzxIF7groNB6UO92aOE8HlFq
TkG+sC1QeOoh5IaPkbhujCc3uBe6c8mTw4WLc/ccZlHKsBBKi609tEhrte3z86vu
OjnASzljrxb5LQV9NnCpil3yFgVWwWrdHfpSF+KJlrljtOXuMM4Ptux53G4fHngU
DQgz9eIms0OI5WqHg3Pi0TIlwaVcWk3gzN45yRrHBLl58SFnhwvqUCspUOUTfyrY
xIqKeWKGdAr6+ssF73EG1HWUGFHfjGxbEXzpsihHSsZs1yOMXRQASA6XcNpDtIV0
kplrTxw3+NTD/1J/+n2BmAc0huWtNRpc8ET4ZG9px2/uwiiNpPcy4X8JXc9Ybf1K
hYmRlkzY1iEEP3oJIApv7STdNcZRIyGmlSvL4gRm4DdkTZIBZZWi5/KKESQQFnWb
/cxOUT9E0Vxs8Wa2JERbeTNL158fHekU6WLsCHDzvy2nXPkT9ckQZsqgVbfDufWE
cyXmcj1+amwvjs3YefxpwonFaknxfJ6vtpIg34NZvk1PwyRNm2AIStvE8OhYTtYe
xWaxZW6Ade0D7dbzLE67DqfgV6tP9BUQlGilia+opS91XiJ6QTeXOrLQ4sk+FeW/
BOYoERXZ1aDMMmoVZMwFpZw6PKsQ047uUx2SabKjFWobuBcNp4f1eJumrvLyHUya
xQNZFpoYredl9JB1FWgeLm+0x3o3+w9+1iaArV3nQJYkWOP0X4/xVz/Is8+wG85S
htDwUB/1Orn0mcrAbsKHC8CJfmUtCMGbRMlxn3z0APrrArg3M2v6Pt8vT3exdpbp
+AdMy7woYXTCfJ73L1DcecjZhbfKKpL2Imirr9gRqilIO6+VNaR01TdbKcI6iLkW
htq95mR5rj+GWnLdNDmv4NPbw8JvpVRMUhxFSbCGyelJesV89WWIdaH+WbUoX9yy
uhnGOKIfgnogRUfmNeWN035quIkI9AvABpSxQorfWDw8kmeTFN7/D4YrH4YOxlix
qCkpUSm+ExFzMGpB59erixJrL62+vBleTnpTd7ZFBOsBWATzJ+o5WvIYmXm7DgTY
Rc54S4ba3iXG6UygmTb/tsOIi3+LrSeutCoYdoDLV0lus2zLCV2901QFoOw5Ponq
HKQ2ietb7Eto5f1w/cwqC3I2ixrzms/9X34ENDWhPX6P6vX5DzzLpw+sQNHJC0Np
dMfB6DSzFXCg6awqnvdrjuhRtBOHBCCJ9icgX3PVfJxqcBoIJBxps60b0PbFOhtm
P+Xy0Rl1+5oON30JCP5xU9Ga50ZvzkIita0JM86r3t8I+QM6KBD3y+FJlP3tSoHN
+XMdqRBhqGHzZZGj3kJn+60GE9pn3L1CN5vjmfCLVwwdrJ6ay55lyfY3EdLlKN69
KtGQu/ArkhJyFFeXvzywcs7icUlMaEZ8T7pmzKoqYsG6wxWQmtvU0AzFm27dbUDj
xR4eKf6/esN6hvc8FcsiYXnsNfMHZjMkbxz6Rt9tVw7bb4rXG5XvGPsjsBAE8bju
khJzgcaoLvAAgJL0WbjJQ6ssxb5ZVTtYbgnPjldaAsTq4xAi+M0QvknR52EfjggF
txLyXPXVgQsec5A/pxlzek563qFgcG66BiBiREjyXniDQkjLkSVvqOSRukX77P4N
vP+BTlDNdJtDYxbSfXdGkyosQHIFGceiUZaMeS6tRWb4aoZSTe9O+x1VBU89OS1t
cppDmGGPznPR+eoahFtG7YWJHAKOqq3+d8Y904+7ZZdtOvz6c6zQKJQpRiMswGjM
0flFsWdI7sFsXVswpDohwzak5e2uBYNcpuxR6tFs65K3FnqY7W9n5GWyBBhS+o2W
OQfdHt4WjOXXDVyAK0dn+cmImF+4KZ+AXeAGToX8UrfokvwHNoaqtMN5Toa98hIE
bt2PpPcn1OqLsw97zH6lDgK8/dy+EalGMpiF1jv+ZrxfADQqyCWXx1C4886KjX0A
yaWqKWt1MqVw0FxTdLPihuPCB59NQ+biFha+nGLX6ieUlWd0Oau5T+K6L8Bay9DC
3DTtOuTGe36wdI4Pvx39D8gKxjA9IJ4PIyi6AKh9NBtUkU3ZAFW/j/7rEtzKEX6C
TI5jXGFG6Yuu5ZByZvE2B7nmEF7jABZeYGHl6x9N7m8Os+k4KsUe1qV6+4s48wmw
+KG3oekXaFJ98iQFk6DalY3pomYoa1smr7Mli7JOO+ak9NCruEyQf+43KDHwFvmo
rBBTlDP5nf5mOx55D/FIiFqkhv9wiZ6i5bvFanXqjxd3sZjft/MWyps2NfRXCJor
EMaV09jBZdYsHoMeB/VnluhADaGGtI3BvfrG/Da1E08GevzR3ximyMcD51/M+Lus
le71ZbHxiTDkY89ORmC3RDO4+vj0YlB5+XYfOoEo7Qxlpvrrcd4eRUL3h7T4jXV0
dJVm0iGiFLR5oKYQDcPhLppPHwvZr0swfJi8N7e+YbwUDru/3an581omq8mDNzgi
K6cgDVU0NUuBLie14FmmFZNS4pao4+gqYZbzOyRmZT5Gdh+TYKIAI5qasJaEQ9ES
EGt1bugkd93VxqHUYIsRV60oGeWyWbiHEJMLkg3CrEMrNiPNzKHcFIG3Oi6Y2BrB
F3iE3zzpETnFF6b6Q87BksjGMUdMys20i83zjaqt5Z9rSHX//Cbln1PYbnER/Gkx
yzn1KzyDAnw5OOBa7RfkiCRKFw7RH4OO0oPKvqepTDG2joK2u2wKX+ls5ruaLxMQ
gk8j6GB6+2ZlaCMBToIkUG9KWZOt9YCj4HmC2bmXjy4jdC14uB0U3DXCiqSIP/3n
E6s/EsMshbhqsP0/Vby49v8zWPeozxQgU2mgLjKWmOzjKNbM2WkLuCrXfS+6ZT3m
YOCc8fnOFEDdfp+gVEaQMTTtqT4QwcNfdWJ+z4zxM2xClBnX/19ZdluysEqh91vL
q1R/a272RwwSjjgYdp5yv9oNyDkT9QfNcO0W8VR2sxBzDZ5rgnqJiNDTotH3b1CG
611UScE9cXsEFk9fbvFxNqEHx8UQGzHh0JLfVWfWmKl59DNkDSe9HcohAoHAoqHy
Rfd8lsJ+7o5Cw9qFlN3xJHcZ5Fu6LcB2ZRhevaG8hnfTq385IBSGMBD8y3lLWp72
l0yglEmKl049P2ta22XiGio5YIdPnq/QhIN1FCfBFRGF/nf8Xi1zmM1uMXHnYAOC
UtPXp2A58H2f4jpCHORmi2MfxS2owM/g0OWtbYps74IAh/ZA5LJKmHyovINLbzAX
5wt0VxqysAJd2Fa6Y2IVVhUkYtELX99myffbxcdZQdD7P+myrtwKY9lnQbrPYgvg
bipr6rORjI26A71sK+vlIWTeOcZMAkkQcm2uK893jU1FJ73P+afakcYSwydBGP1e
naJ2jxI2xyNJ7gaKi4f6ejX27Jivof0sNuNzU9SiXa59SotwEcCRlV4t5D3zvArU
PwxKzZeEH11y4bHBag3ELz8zTrsZuT6w0UGLsM4QinLhhCXksyhUcqVH+SeKbeio
6UWUwMjrQ560YUSfkM5xT9SJK+918JHjmnCik2F1hszYQzjTQRAamLCM/v2vMomJ
qe9bJHYw/ewh8Y/rA/ADY8op23Pg5fQDC0a6EQbhWaRMSJwB7g3tR+uppUXHjmwT
2JMQiBxoZvLe9GkMPUTTBCRGwMVyLJTwQoYUc10hVN5TO0pMvwp5Zohor6o5KrjH
HB2jYwVGJS8kPTiLSY8mf2MhAG+7e9goHeC4SwGGVR47Ojwuo+ObD71EwrKUBpnT
BGuWknM6JKkE4WUBIVuw+t3jSVFBt1wToG6VGRfYcnB6IGrleIwcKxLaJANRFVPV
nMNOiLBNqA7L97vNLlAont15qZ7zeeUxlqn7Isn+eCFnSzn06DwS/uktysy5E5A7
tT231LwNrACrrCyTp2vtOo1UabqI9J+GgGe9S6OAILgd5g2v/+LkjPi0c57cOi/U
q+o55KbwqX7XBBpImITMUHua8+nDXvvC7U9Yw3+WIHnvS3rhfn/2fkq8dFXbfIdK
iHieyNtpvzh5tyPtP/T0KhlnTr5sNJpoPXgmLPdSrbdMznej4r8pZADbM9/WAJjB
Qdn1GpBFuwbbynvRNsHSfAK7ZrZ9N6PMo4oK5Bbfauq1jTJlbyWthzdL8Ozw/iSi
ypqCK6MmB9Kj4MuOPzDfj5a/Vp8xFyXY/Jejfo/d7HWYV7a5QM29io2Z/A0aCeJd
PJrcNDr4Qo/k2ysDJPYUO1Ce3ig4+0pRaBINcvc1m5qQ03EjTu+tJPHzpACUgTOE
OnOJiDyGgZIYlbo1xIGbS3Uyj2DqrylGiBK73sstZoBypzfFY7u8+wXJTsXFNK0G
V7vk8H5zOFgp/RLlYOf1ldaXvTrWBmS0KVHmcMsMbGBvTEjAKvIbHdLnizZZBXqs
O/LwWgsby6bjSb7wIXz5zTcs46o8czqGykDNtdboBkncJ5Su8qk5IbXF/4RqoOOc
IK5nme7vA3tDZha5lZpHbqMyr7DZzADOEl66sKkxXgktxxaLXdfN15walR1y8T/U
NrKWrcmYbVLsyLwDBLzvGzMFJusBy/EdK2sTwT26zXLSAvwgn4wHW1Eu4X0x/p6p
SfTLhLT/yd9HBKGSay18hb0JZQMOtzj0/U4/NLzPCBlSXBkubxtxBxEnbMEv/EYl
ODnVk1u2si8LIukfwHTaMW5fvoCQn1vU3EI9TDrgqk9KbmzubHLi1oYblORIHrDR
V0Zp5idvsnPytLYAslu8ssm/8tdR4LOB9CuPpAWTEuLx9xQ8yNb3PGPt5+KNuOj6
kGNZ6V4DAa0BV/Ff/b3MTIthPcUfir23V/6mlOU/yOSCA5MJiQq/ty7wCiBnPpQr
CPfvd9FBJVg81rm7c7jAqwKvTHSrImlomhmVhsckIoa01ZqZ2bL3IGZccJmfYxac
X+njNJmqtlqrqTGTde7fU53zaqKGtHMg4tSsBnG8v8YBReWZXoSTk5cx8ZqerCQ+
xBKGFNQZ1j/2nrFERSFOF6graY4YhsnTMBFKSLzidSB4Hi8ueL/TC5EBOCOpKaoC
mfH83zXrrM2Mmo5FtbHkvnBT6q8Ieh6Qs6w/JCPUeEvU/sPYtrpAzm6XwJp+REm0
WB6s8xTAPoMbiyvOWrU3mVgw+6TqbNbdlwJSTHVP2UAjVfgtpkYR9qLxS5uIz7p8
rAewIoy5hdMQU18sBK3+CZuVjtZw92o/svv/WlLB8WluGxtQH08XKlLjz82XG8EM
/mAKMlTiZ4nHkwyiISybvPUDs5f/KzAH0tcp+UtjC/DqXv0kjyx5MgAZwNtZX2Nm
9dxlIDxVny4MNuUfNfgQSrPX30impdmTVSjQ1x8Vc10HsyRQiUUKEMxfoVKBvxqN
DCLB0k4MG0XBgLBIL2D6JB3lK0+88whjXIygva/ZILRtkUZJ7oboYKGq/S9il7rb
y71EkHXriFKyAq8GQoOTP3zL83SIZiC6CPb7FY+b/sompBKX9PS3mP3Lhe3srK4j
IWargYI/qr1T1+extcyEOPWxO3FXLcZhU1hRedBrXN516iP1RrFvRs+brPLPQ3hN
Idkq7dXJuYIdCd7WHN8htd1CJv/UYC/pFbCSEGOcTH835Yr0fcTn3SYvrYU34Egl
EBHhpHg0FU+50MDz0Q4YJjwubh6u4rNbOsMim527fmFNd+oWu/wvMYtMxN1nm2QM
/tyHPKfbbgEqT5FftlPSBtk9PmCbKT1nFurcEXLedIpmP2c0LLuGPQhtOkqHJljC
PTVQW19Js4Q93js/7bU7j6jq9qd8R1SCjmeK8aftVnNxdsS1hHktdOkXGbIZZoOb
kU6FNw486t/Pex6+sgaj7OfarKRIhEUW8JTN4eUa9Yubm3eBuaiA3XcBDcQGuNyn
0wF/tv+pmK4PelDXp3zO4p0ZJWOsX72PdrhkubmGmNszWGfzLbrQMhcne2vk8MBM
5rxYk/QnrrYqfkZgxbWC7mpQJ8U7bpIeLS1M6BQFB/zPh2ifdWf8wz5MW2Nxevz+
x8eoCQWZgbdNnS6TaEU3Mlf9ZG8kfmjuhTXO4a2FaT514ExqaJ911cpcKSMWcbnA
PmBM+PqVMGuwBqlTZGIIoEA9s4ifcHGTwAPCkM4pT+wkS7puWWfWpD7pGLIoRGt4
4dsdZDVapel1hVmEiXyTm3fLylepVCWxDLJS4Bm+XIK/8sFFIgAufO7ysuCCQi/I
DgF2/DuKDdZgK0nZ+7tY7pdzm3GjKn4LsBdf3Pnw1LgnHsBTe6oTRDucsMyZljLX
4d2A1d8GQx1fmEWkeihKpjcM46riWxinmEaBqmN3H7HqkurTxl1mDhS1wXR3OI29
OmLlGQbw1CjOF5Od3Oz6LI69GqGR8X78BmxUJTAv9otFVkKbkcBT93NhfKQplnEd
oXbY0H2867lz+A+xC+0LnTBTSDk8uqglMfz7fHoC1ONzoNYiIdYlco5Ar3jM39CX
vaFTPnkWIK0bg2JrzmvT6IAaHvIvvJtg4XW0nDHwizyLmzLDfgIOYXmuWZQ6nuav
qx05oshcRdLa8yrQmFvby5dASsOc4/ZtVBknH7YSP+gtrM8OwXpP/719QvfF42CO
nv9ZumApVQ6Ou1beaV2aEtT20pCLT1nGuulNa0sSl4XnBX14Bw5wL8r7CfNmsT7K
b9uLHu7/d8rTqIHLXhhSAuT8z8P5SCopDDWkzsTkp2FMYxKXhxZneDfacN/MXtnb
73xDqqXHIdDHjW63QGRAW1YlZskztyJhm2v7SLeOT1h+AAwNek2g6q2rkzf0cQzr
CayanBjnNAtkXV04J05aroKH5Njt2XG+c47wJPq1+E1/1KgqXG3xDs0FdFIoy9is
GCYJ0+zoBVrFI/vPzkm6yPA7/GSvIRmq8ED+/3rmVIrS2duHnZRRqCkRjnTlMQrU
HDXTbQHpX2SRMo3UBgmt/k7mNJPBD3S5FZaajXQTD1BOnr1NwJLbaRLIqt6NrEzJ
iwTjALxhGbPCaA/gHjg49DYYDczP6aPMANWzLsXzvfublBBxhhKlj1iyQ1wIEP54
znfU4vUsSUJ2+AwB+Vn+onpPNRRx9V+Hd+yzSbPDHExLyiiHffxQppcea2PtXHjt
E/c4refRmE1aHRbzIozxJzg7DdppD+lOTnB5MCHd/Xj/2/ACmxqstutes7UrOq8T
LIXUe5Jhz7OsFB6oERYonp6b4fevqY0BVRjWc0cj5Npb4hR14SUVzIyMm3fJstF/
+CC1d/qYuFJ48m7K6JnVXGS1cgbhEVUpTxBqRJlVz2OFgEAFeElEcS4lDHpblAtU
KpP3Xw1CKNZDt2K2ewwFEbFPIlU2RbH0PvCb/0UvZfCzXA1i0eM+EA4ssyvPFxG7
0lfACiNLK1uki2MrqKqba6K96d6AH9cL6yZOGTn76oJiWCRpkO18bzN0Du8QxqBV
/ctVF6ieSpSIV6ofOdURiJxkaHUq+ZxPZR0WdlzJ51YzXhe4mdV9n+yVKZE71Kyy
F5icloC99UTR2Lc0lEZD3yUwbnK+kwlg4ZT9K21QNwT3tHqFYjUtvapFuhFcJLDj
Bd81LsQjoIMC59nyJoArzMJgOkI1y4l4UcnY6mdTY1iE21MX7Q1hNpO6WoUwm7Gt
tdgQPiyRZy5MhLePPpgd4qC0RoZ9eBnSlVcUdivGgAjVsu7eqC9kEPzLZf6ACxLr
4Fzbms0fg+L2luMw1IBstJjl8ghB4TznK6mAb5DxR+7EreX71izITBFUtMYQ79Tj
ZS+CNxJS9bqcn2vz9iVsHkvj6eYVph9laaCNPX/fC3GrIPYoCfJvoEZ+MygqaC07
UUQAIA9m4Oik61SglNSW3yjj+nX9ykP7eUPI5D+nTjmc6s+V0Sj5IausApbmGpcj
BntWhc8sK32fjRxwHhb2tFFh+0RqvRrefgoHI+W0eyaIUJf0eGWn1vJM3pe7SHYc
EoQEHOvRlf3bbU/10ej5lpLupKt1JpHj5FIOOmbs57wE1T/mibP21V0R/Re5ah7F
iFICez1M53BD84bRI83kk512GrSQwi38+ZUyZV89xFb9QtL+MaSNp4PgWG7L92gB
ZRhW3INhtHS6PdjKfQrEV3dJGIL2VGTHi+vSg6NjkBE3cJaCD/6jqAmL2LZjKPyi
baHwt/kPKJEfMG6RFsCu4O/iVY46joEATbKzEdKdhiF9CWk7l2cri6i8tantlF8O
CAV16+n1hwk5uSqq1RrimuTurpwopGMgNpAj+271nUc5MV/PgIob7vK1AVokwp7L
MDGRUlVIN9qM0K20Nl9JDveE0PT+2FQpKleiM+JXrYBUU+KH4fKOV62TjpyDtrJK
tE+e5PQ0TkOvgwETtVRSI9eRHtnrFRVPhjwxxTHdmem50rhpQJuqaTHSHl+BiaN8
K3JlHhqfOoXAEHTP8wh9LErRadRBvLidKiOSv3sp48iV01lh1J2geCsal3B77WKp
+TVBmdZLFX7/Jbh31y/4bDTTfd3k6+dwl/0rIDYqfPzvRUP0tqpncYoYq4S+Dn4g
m9b7FFY1RZN0nfMFE++OfPZ5uY6dTSXPFcgh6oPwaRIIubdS8Hd3bZP8qLSJSruB
Adhy0CPY/hdfkioeWlEiwiHqNU+tWPNMcrsDl7nr6LZ2wOc08iWUGdwrp1o0lyXm
9PIfQvVUzNDGuOfnEJVV0YS8Y+3n/naUxEGkyfvAEbNQFtZBPz5yhCI4ecBJERcK
ZI7HsCij4U9/o5TXIlEkcwBmcKLsEdZxUHVWAN8Qw8FfvTl9fhKZ30OxQDgoi9gi
VUL3WJokkKTf/7irUdTLHE2UH2mAX+F3bmPPscyKc1Fs45ijbcYPNAzdX8HuroGB
1aJ81YsVvCbG6G6Ib6FbfxmYCs+y9V/nrMFIDdQNw2uEQoeZ/hhF2+g8fxX5kCFX
W32wMpuXODhBJvnHW5sD29pByzQplm1IL8rAtxlMXS1q9Kz3jRoTT64T4pV5ASPJ
mNQ2TTH0DK1J4P94u//MqSQELpsEIuXQogjAihEOK5Y2ffxeDSUf4Fz6O/IK/VXP
b0GSARlAL9cmGlTOWIArcjpEsaXIHKO8o7xJPL4gNoHyqDdv+1HcSNSSiB04r9VT
M7TmrshNhjsTQ9nr5F32BXO3D+yw66IbuPdOz6GL67/8bMqMogGjFDZxxzClyVAN
D7G5/lp81v4jzNtyEiYtSDVsUr2PvzxA3bMS624RFBJFlZcPpaCxPXUrnhUjnJfu
sp5/PnuWGSq3KP8t119Ro4CMHdnj7HfwyptBZXlXh/5gl9XgnxFDcedDMcCFVD2R
XXMy/FTKKaCksSDHpre+PyNTD1j73ot12YRHnIWNdcJVUDbJpNYU8vGlWFAv+zeU
+P2tiVItiGshgCrHQuD//27qt6Ag4RCx1wIpN6MJm1GazVBFvb1pXltk3tVeO+zr
vLMQWfuheiMs0JFpgkTm4jqNgXOt4MRZngDhafbJ4ZkFgoGLabGsUWmjZMEh/5Vj
M1QqdWL4270FPDXlM3an4r0HToNjDByT+WSg/2yU6hd4afRQk/iXqCyPby0T57E9
llbeD5VmO2gfNX9gmUdjvgaZMovHUKerUiAScaRbFiH5C1Z7HrckSjrSayERn7qQ
qpixhL4G5guKlZBs7YHNItY0nzaBHmqzSL46f87Nrs2BG8YrthoatuWMQT0T3Ill
1U15SYD6Zh2nx6Ez3CProORA8zCfr38OKOIFgLOZLXGttg55LhdcBgIUXlIjBpni
uL/CkSHidEBcXBgaIGsfmpHmxjvYiBtZjs+1ya3Q6eNxYllENvteZZcZGjYQL1Jc
0ayjP08lo0ko5hRduBeGXPhfGPXHHAv7eMDVx/D5lp/m+8gih1+NEozLnFiXbonL
vbAndU0iD9lv1mUV2+7E6mqZhBDEP0Nrn3DpgPLsqXnCs+4c5Cs4t10brnNpuxOw
U2A3VGocsTz04vIfUVI1NFiu5MiigToTEDWhvymsZCxOUdIYCEOOfBzaS4wn1Wtn
3JkzzMnrfsrYDGEOgKGEUZeAlP898IINSf03HMLwcHwrON4vlfoF5ciEBKg/GVQe
rYzYKixtUdopjxSlE2P1LfxRBOiKDeoQFQdqVKPohumGgeGK4wpNOEUC44hdMemH
c1TxWvjHG4lwcV9jXtH1vDD88hxgUQFkDqNQE5gkEPlaKb8zzyyaDBphnftzvGCi
ZRDw/+gMTXKZOyqeXa0Iw+Fz9awJuPYmi3y/XMmgc+31jJH0svt5alr2/KCPL/U3
+/8mQyexpkVSU4XFGeUioILdHFuVSYTpktSoV+N8To7xW+WOYqEOJbkp9+T6pfE3
Coj1QDqKayaow8CtQMv2iXtpV6tlvtOCALKQdmZdIwNYebe6WAccKS+ytKtISgG3
Lcwi1jJHJgUHpzFScK+NDjHaPJ60oLuw46tJuLmTD5Hyx45plLvk6V5SR9uWauzz
0lkAoyh+Kqor23JZ240VYFXFihNXCdVlopYMMbkfniI+dhyvd09+p5noideyuoa9
EGWCPIutirhzYFuaHPWm0RBtBp5MrAXqqgqZWtjKLq9XA3FO6ein1mKcpnF8ME3g
nvI7ei1VBhTrmE0AarE005bnvYYHDgTeKsa2FcOJeC6mBh5LIdpcO2sdqdhnzCV3
TAmgFJ6x/UfDjP/PLBfIGvpoOlcYYeLMQR3UTPgyWoBZQXIOTl8dh9ItFY169YO4
v4xbB13Dzl4TP7HU/QsFnHBDwmBgSJ7+ExuE+bkjO7xuJDIYU5r4Xx2kaMa1Fgb1
/d1vx5nkHBb0CbRrnYlgVB3xOkrsK5dndvxbe2JBpg1DCz15ME+xCyL/6bsm9vF3
qCnjWFDM55IofV9THJgEA91bru2o0+dqbGo0pXyKivRrOj10e1Q4+QIQkJo4GULs
YsRAk/uL4jIXNVMfO9xHO6nSYobX61V1K3D45s+1fWaiD6xqys5q3Zq34QUom80L
753x63/vAXlAIlEEY5o0acXNBSf0odjtNKYIoownnncTau6nXgAlxQ8LKuqqXi3f
7esMYvt2jH8DgClXZlJpcWJkAvwtCPvpkSpHEhy1JbYvxDowECOG2tbbWZW7zJL9
pFWW/Y78QJr3XOoqXGlrEcDXCOheSnYeEguh5GBFEbN6/NgU7fJrYw2gSLle++a1
rPD8w3Az4+VxZAG75Z52HHo/t5q8OOZmpffsuWZUOrjC3WsxavA7TueVvhaaiQyD
bEm/hdNwBFYJXzFX4uq37TrOXFPjAc78br3bWgTfi+SogDwINHubraea+ATR7JQD
PScJQp8lN43OUIUnOHPsuQCcwHq3Rq3EdTr83UJA/3j54JV4HHYg6aFjYw5hVy+T
Yuc8nPW4RBIYZHnW3TtCN6teKJ5NImxbI7J0p1yEb5g1EYxrX4um+8EadCSt3Dnr
QgYIk29K6YMCgndKbzuQC3M+U40EpDSi/5Q0/KQTG/85jrVrALswFOB81Tk9ews+
RVvTaw5U2nVpoezpIHhuKJGjLvEMaZTa8jolmZdE38Hw3RKnX6FlR+hmMjFsqBVX
xrBe3Ggoh7pZgpYaKiGXNA4vjHQI+AoAchx/ohb+kR6uLO6iux5xgFqBe58MU5zI
mHCR7jiEGgN9Rsz6wXtQs3GzMAkGgPSoQE355wYTWGR0jPk31kiechK/XUPRrfym
LEyvtnBs8K6+t7Qa876jz+/VLlYp9WYwDNJeJxytWOVpvOW1CcZbVOJvOVD0SoDF
B2+meWzTIJnNJCLqQDM87geyNp/BCt3Pgky3OUJdcHDKdA5UZN+13xNbp4zs73iX
j4wwrnpR92TsBRgr6snWpn4gbprOeUNbNel5xOeV/0INaum6eyhH5ExSIGq5HVSC
E4XqCOc8OFUK/nQuphcnIKsBvZjULD3i5G2Tq7m5jcDcAkdjPO24ZIsv2qBYa0SX
Exr+MejV/9w0T1JonEuQC/Tbw4NVEQGoiaQDIhgwFWbo3iaPHdCITjb5U7wXJVtt
v6TZyKOZhFt2wFOYU3Qe2wfWqzE/iOqKkcW6f6Itv/Uy4xbJwKwPcPCtRu3eh6Tw
HIT0vqQm+h0gZiU4KZyYu56yJMTCbVdTej6vuXa6DqLh0pRymcSaH6fxvD+znX6Z
DFD9g8r7HgzVX01Z4snFH+BuftJX3OBbWuQdpqBfRwUzACIoCKDEyxfuIw1NK2HI
I4p4sOxsYVd2sZn0GgFEzq6jgsxYjD0iBylqhpRiWp21vWYtSHeQ9x2UG+r451l8
t0eEijkEjEMRuDNVxua9h5lcWjdGBv29t6Mp/nqGmPWitpaW6eWWDTLGNwin8/HD
uoJQFl2tw70ht/HoPIOu00hildRYp5aAo1+Q/3AQvmChmaq4GxfD2PtxTU8bh0uT
XW4kAloSAwpXdEkDO9/rgjEfyFvTI7Rmb30Z+SaCUqRM/CzI8MY+ES1ro8aUedBz
h0KkB2PFcotFStM/NEzzqIJ9YcU4A0sxjAl/IiM1EeXuZXKW+IQT8qfhbXcgUZ+Y
HXV8nxkSYu0jRWKF8Thlhmq1Jfl6HtLQDXQZkcfHERZZmT8O3/+7lfSLmO38DQbZ
sodpFkOSpOEehBa5O1bAixySZDYn9B3FO9IKefMothEMDttzy7A0FcJOjE0Hn7O+
kycgkg1BGfpOEFuZMgsfTt39mEAh3GFG4frdncEdizRX68csLPFVAjGtHjAZo5+H
TYvMlV17oSe3cT7wx6Zx7XTtABICbnUI7LHHEkYJ1AS44O6FCnEQpO0Z7oAnjpLz
KgHQ/74g2Uu9eqvPX9kDFW5TUj0N0tdiDLNJ9dSnsrtNm1dt7Yh0qmWhICyTxRQ3
OelwlPfQ+wpwzIO6sYl74+eA6x+QZhiKark8Tfnys6BzS1aumcBzgq0lzJ3x1tYd
zojECRJnlVQH0g45VkeKh7OkoMkYPsP876zwwecHgt1F4cUNC/L75GNAgOQoDxv3
NXB4GhhnjVbDs5JSuSoYWZHB7/nKkudfN+WddeKlKEDtFLs6dgtjt2FX/Q6AhSi7
rxbgia7Zeke40LAr32Zb5RuEOJaWp84ll9asbtuOXTWU4/4YI4sExCWLdKuudr9M
8cf40EKCpLo9wIChxh7RiFWfBVmk2abk6V6UnBdjy5tYi14XcnId1XzMFW7EMbv+
SvWnY3++kGLZotog3MnE+tNKtYnD+4VVmh3Fwx+DG965yD/3rd5cK3VxCUZcjIgG
JL/CBD7UAQbDo5mkN0DJPSkfDdYZ6+C3q5zQFGjiC6U/mtAMa1VqQ+5OSoQM+ibh
SgebCzGDsv7pgKO+BKxrO3NTBownK0B4Jkp3SSXHgIOiUdT8hOBTQclSJq5bLgw2
HOWIep80tf4njuYN/Ln6tqLOZhS8jAcAKojEF8xYenKpPdd5ime6ONlHSySxlXeV
XuUAvhB7WB0X7bIa18tM19QYh+IIu4wBTgI4QEKdKqmCmj5n6C6uwZhUKxNaj1y2
mRn07oh+em4BZtJiKWQnM1OKeku22pJdblo8+tMdP7+hZ2REFd8S4yqf+Cf3Kb6w
5QD/9XwQdd073TlDcVyy62PSwcFTXrGCI+2f8qBqObSR5qx3bGLEfUaxYG6ValOE
gRnaxiVlfdU4inkbmrLC5tU2gYi9ltHZa9ldA2ZPT1i8jJFRhb2vTgvzoiIC7J/i
plMD0xhF/5MnBYEOu4WYpHgYncmr0zL3r9equtkZWmwLPv8TkgKyDbJ339yjSDm4
Xzy/bvHw/zNJOyay90WBjLv+r2ILtWWkDEDxbPUUPG39GkZ16flxCU5vaW5JutGz
3HkPpiwWwwOAZzZp+yR7iIsLEJpEgvygiAST9fdKRTG8L22gdRjM+6/ZskrqdwJE
Lkbc3lNEmvH7tagjN+2jKSN8uSgPCvhtK6kvAIv3ZCOQNqrWoC+VshBSa7uwPR6r
v9tgOtf5DOpYRco1w5LBB5YgcW4x9D0Ervu5LYxh4UCcJ/eIucwGpNMgQr9pY/Gc
a2lLDPPnFfu4A0576ceF3rbF4ImPpL89ZLXaOGLpbFKXNBu5C4q0/RNOH2uEl7pD
ruOH+OAHEIVoShOjhS/fXunfJ8wdZV0f8PeVs1EeA9ctvY0mE+Ld3HITPAY9wCYH
wylJfGWqz/DSOchFLU7QHIfbkOlsf+icS3WiINJOU2y5aKBEowQuTbVLFX6a43hg
vZkrftdxRlZEWM0It3jtQnSemw/CqodnRen91qoVclbKONloo9YTKMIIyIXB+Dpj
tMNA7fPDxkPWde4cpR8ZQhLkwn1mQ5BVFEFuE7GlCDT50s62BP80BxrRRCwyT49k
ChT2JkoBtTyVMlV/4TGlwQNiDNzImKpL3M3iPPlUBXrzWxq80+HZ/pjcSPbNHZus
v4KVD0Y6AY/b96oLnxwNMZWqQ+6HbU40dvbtmGtQ7HPK3/K6nj2Nam7IuJYnmMLo
asBYECKkObXAu/1vFvtZDezDucclrh/OJsap8X6vMKcPmzKsCfYlYvM197xhWisB
WgvTa7kNxjHyDgUgsll8hbH0+GuHIbdc2XFHuQekgK3695xdao20sqSFSlpJ3ZTK
Ma2e7+JbxAq62L+F+k1xUMiiFOnjBLWDeuoZ75Q/aXR4tb9zMt7/YhaJPCzNlPYP
mrZnbx2vIzrBrv/bAcjkXiqnjEFoku7MT8bgLtLUOo8Ljiy2hctzsiL7Pa7A814y
c59al5EE9RLsWxTRspZOhvk2pVZSZQynoCxtymj9h3pFR9w/naEF9f9XteXb7zIp
lGcL5+/L+4GHI+z6JWbSq3MCwhIardVMi8uTYhKpvxs/a+nK9ITXJl0cHiXXXO5d
kCM0jEX42v92VpgBzgYVCGrf+2KTL77bv+PjI4oxlHjarKoDI1/bMNXz0SREqbi3
Tlk0hCPdO67WS/TlOEenYIDvyI4/4ZcPbjaWexGIBu4nsafEmTZjNdZqtgZgSthJ
vEyJq1luMqJl8sizsS4CDPlo9ZxpAAWUxTakv+aaeqRI7/EczB0U3IOtmouamRGO
fUF4t6qWRITRIvFk+xhFWfL3voVhMcTVytrwNNxdoA72pFS9G1mmsFe6z4I2MuVY
9hWBnVGlzgoAdVJpbGarxq84hCH3fhgjLgsttYOe4KlsTk03Uz9mX2nyw8LY20km
g7Pr7kJYXJuTysx3akOKiezay4Z/Hbb9xawzMVxesDt55JQbPLP/+n7WsV1BeeNG
umtSQsFGd5zVwLED8/Kc+x1+CN5o8TMkCUZMD4oqQpAeyGP+nrRbZIM/RjwhCFUW
k9QlhIB+1MCfDacz45yxTVpQ5q75LSlsKmXeQ+70XKeZ9cnzkkAtieSkSe4GUfO8
g7MFvEBztbLuZ5bE4WYSPr/7Req/AbIzqrMGlHZZKWFocjpY8GpHcfSt0HKFZ25P
hVoKIXjqLgSGQWvub7qephs462pLTn+48efrDXE8LzYGr+kqySJLMJII5Gt6i1bh
kl4O0JLPC8URk/JhTqsfoH58kBzUURytDx4If8UOmizvue5WASr4l+gNgrSXpqDG
RjGCgZ1BDP9B9jPUf6PpOfIpYvmqQNtmRcwiEwsWUzUSjZz/1VtPh2I6gRDOW9Wu
7dNOUMQufz3e5ESNaAL7Imm3xv+i4HKsBZS/xcy/KYXpf7Su/BJfJKwhZygIaXXc
4N0f74NKS4X62jPwtBvBFpe04GqiBShbGdJc8wjuiEa7t6aFx61uV0Us+QTnRMjG
orDHF0bZUupmpFKMGS58o2miK/05zTFYC3lefpE/1EtzUQOuMrvqe8SCnOs2Cp/v
MQ/V4ugNv/k+ugO58oK5DsBCglsWhrbmw3DcGruYSKR1mH8g0SbbVXbGaaQ/YAMj
NHOThMPNLpyE5uPUHRU9E8mRNnDYck2uf1uSgXUbJLWWit6yRpliWUkzexZZsfwS
zuBST2npRxxMxJCcrMa0lMGcxHfmJGRHJC7zMSFy9vOv8p8EjB+4IMubtzuXoE7G
RvY8wTS+6GmaIkvRlVk6qa3SfIiZWQIBil42Qr5LLOq56ylO+cRQd553CULBU1v2
QDQ6oLEoOaFdtRSFzWRO6szbZefMtAyOKDcndvG62CjqISp3Ez6NlLSOX1j/76Nm
cQCD9ngQZqqEuAa7cl/L6JFE92XqBEVHjNpS/TU3liw47emzf3pwOUQ3t1u+ENLn
ENz15vnFQYcgEfC676cj10rNYvd13xjUlxV+h5wo7A4i3PkY6Fv+D+AhIOFY9hUs
D6V3yxZ6/3NQmeiVNAm0iEw4kb0Fp6JtgXdP5pMgApG4LshLuVUa/NSc/FfvjE4Q
W0G5Mg3VC/ow0RmHFYUubFCABZNUkUSnVXnDc2z25z1AwdlsSBFXo9B+eZhD7VZE
DDDhQz69Hc8CN5LTX2cP72mXbexT9OIdAmGt7LJIXnAIoyp2Hc3/zeykuwKElw3C
anMAFxUQQfr/wnqYoPzZXwEIRhE/6+cABEHCPPMXaoRP4+m4UYRTbdLiiwU/jfrL
INc30kj2loI3iOAorpqCAQ8F6b0vKsCcF2aIqFM8gIrwsESlKkBuldmoALFY/NNJ
KbQQKUOdHCrXizFbAX8BX2ml7C7F3ND0p86SLk2IQepCNK0aXX0N8y3qIkoeV6zC
95fjblVZdW+cy7RBRpxnRcePGzlOhiBANfavmyOdUZG8CoCpVA854iO3xo9FyDJm
R9QS+YycJOSiFjCWAPedzA2fTdX/zE0la4Y24OfmhZLwjqIMbR+ETlwRlg8uQKy4
y17bX85QqNU7Q4pBkv4Wwa/+D5E8B1UAOaZXpkuc4QdiEAnfng5KbpPxwvRhN9t9
vl2SydjpgJR2Xg8C+2aD+cVa1RotNL/Ug+OugnFmyHijXCDieaJ3MRE7tgiqpaTK
O9eWYP+AuKqenjca2jDd0o2lM8CEBH5sGQ5lfv3xZdY9ALwGd/7PUG3Wg5FhopJX
bF5uC0GgHN9slzZB7GThKNiz8iX1Wrasuhbfp/ZNNCWSuOF0pjDN6s1wJBt00Ijt
63Ohzehet9++xVHssXQWF/M5ZeS1vsJ8xPUS+4rihKRhTO5KubScPutiLhqlflvm
xZslK+te5xKIH4+JwdTLs5QsRodUBMZht6cyhMka5P3qAD/QJeZJ51l76bEtvl3t
dSpMwi+Wsir8v3fGLsSmEGTCYHc+n6ilLdv8NTnjGoBWZq7+Dlb9cOugyx7lRG/R
AK5/v6c45qxIQnzPc1aMXST1S1ieDIFJoC8WFWJsH+5TDzWl8YqCfGc/eD7tNpO5
eAVbGHPlRHMpnA4IK9nm2G9DlEIYpVTklxQWeEMerTZG3vu9Rx5Qd9oIbALM/QIr
mjgr7iXY3XOhMvbgx8fH9giSfFXzwJQN+RBw2ky2/BTNFcEsFjbokhc3BoZwcLMk
/rYOYZ6doDIf3miaWWHJpdB60CE6hOqCzh5ItZderM88kGZGRr5S207W8iunCOGk
YUc5enxYiS4etG2Z3azLOp1Faf2rhVBXP9AEmMVT4vOWz1X/SyOV1AmrzgL3OHkj
wQc4LL2khARDt7BNG2htsSRZ6a/kdZRWr4CZLTj1HbA9dSzLU16dSryS+GB0NE4M
Yk2z7tcodVlCCUKc0UVSHSuP7r89QtRKRDLgGt51ioEYuRb/5tW0j6o3CIqp8k0Y
+2iXN4EfSbjScHJ9flIpBZOee8gnHGUJBaqT3VSoINwkC1KbpA5ZAOqMsWVT3JRu
L9USBvbiHvtxPWV6NBxweBTKTdBGslkm5Miqhb0UUz4BgtyczxaZM0lkYfT+qAoo
09t1+gEvZvl/ywe6HIOdTIyJ6w1pljXs6Hhr8foVV9KAic7HzK4ydPF92sP18R5c
WJCl0zXpJikF5HdO0G5L/1VFLMLG6NGyo9CNYblHjTtMMISKnaNzEecNzRZ6ydpS
XoSWVRTvOEdBOl0XpVgASASCLgMABoZQ/V2widrUX0wqAINF96nohh+KfI0KWsir
qioYI6juYWuZlftG1WZeDGHIA2hKBgLb7evmKJIeL0UV7IcjrAEHbvoE5zDK1Q5u
/IfidQwPD2+pCBMR2sGt3rY60mQy91tUJI9Kzt8HKyO3DXtsAQPzcfLOOP5pjw7E
L/Ohu8X1A+xnK/j2ZPYtU6MStTcPvj7Y9RR23E5koN2lFG459yIaU0xFtjxe0YlK
VmtOcx0ZxTRK4alogA9U21tqrhj4yhiNoQy8EbgnsyzDYNg1tbSsEK2f6nOgl7ON
RRsmwcEPxz2RSn7VgGP7mnhLLNtR83UVGKtYyDDRDuNsn4l+Z8TCYB8HI0b7Vjs1
1wrCNaqdnOC+3TAGyv594mHQL44ukPdrzHkS+6MLObiUm4bOzWJHW2F4ToxUZvQi
vwaOakeco4cc2ganiCEj16Mb+3ywzqeTLxm+z+L/0pix9SaEXsRaDyP9HuiPnieD
x3TATB9ZqKEPfaN7BaPuXxPyOmgQEB6BcCMr+qA9XOifcZIDCkufXdMi+rwytK3P
TOqSefi3NAUwo/n0nruc6WRBgrOfbIgaEq8rGHoMIVQaU67QvvBo8Sy/laOsSH2p
WHFCVeSUA7FqrmslSixd+nTTfRtXUz/GDbnPgziXfra8AhCjtMyUudg2aPJfNIEB
sPXklvhjJ4HUD6lu02/+9lWFhqQ5Ec1PDE5pZZ/7yOHG/qUkUJLasJ8VJ6ouUdc4
yUnYq8v9jnAHmDrNHRkMtHB3/zPOHdDv8/JYsMg2zv9A9fWt1gVRJXZET2Rif1L8
5lWSKSz44KdKhW1/TAqTW6W3X+ueqnALRJNfRAfqINjU5ltit46mC9KVmVvAi3Bz
Ugn6iJUMueyeG+hSv1Q5ho2M+3lyp0IdxTFqsMoHJyywK3fUhPyvZHv7ZybiaaIS
v6+uqPbZVGQZJGkg+jChyKpMd4X3MqcO+UPFFmBz9Y7bYparEZvJrVgSpgHhsV3M
lOI5CWP4h8FeRNpT/xD5v/QG2SbYYeDGcwG+VT7L+xh67t8+LevpB3Wd2mJjcfP4
WhkKgX7jT9L6grDXxaapQ/zbuZHzFkXskxVoeFtMHJ547Bhtl8PfhEa/4tQ3F7Ir
I6RU2jqz11TdfHyqvjg0OHVOmhopg2v0V3xiEH7fLndXxsIIrz6TpdwTyDHFRRV5
zNOBb6g2q4FFIPsgq4vK+Fyl7WBwlom1EBNsZ6i0KgsKG1PSg7iLxaZPUGv55cT5
TdU+JfvtUDP6z2YFvMiqHs9tiKied+8lnXxhR2Bk8pCYXNmGSrnAoKnA/DSPr56h
EbG0uEjVbLk/1XV/axBxLSFRj4B7oIEt1lsVzh08HMraA/ta/zVi3/YmOzvzaoGp
PSFonjUTJ4zh0e52hTHjyPifFQN1sNv1Jfp37vW9e57eyR/iLUVi4JDZvnDxLZEb
77zDbwMkclQXalc8juzZ13rINfSngyB+sSwr3VKBO9RfhFUH5D7l+OT4wo2MScHP
9Dk934Fn19Dc2CK19MGMB/l0ggXsRRlhixOHp/fX2UIXS8EyXiJLrMGqXdrlAMcO
pUTAZzdJADuqoFeXo97GfhcDqt5pjV/+7vfWi5hSTGY8+aps/JBlWECATHnenP3m
f+F2uNKxsyiVRo6wCgcYKcP1huPw7IGmuXaZ7wSGOPX+sdTm2AzQI4owmerkCb/Y
+qX29KEPV7sUnhkdjhJxn7T9JdaX7FBBQxYNApZzNqoP0axajuqe9ajsMa1IRiwK
VoQSJEogBWybBE7jFerAqEGGPFQzknUFDfIUzBd7Azxwm0solx+lpv8dpOLktixU
rXtP88ug7E0znVXm96VeZY2WNy5WtjeAfpXHXRrAlz2a4xdaNxYsJA3nwHRvM/83
vpF25mcEqXpomWbitkfcOCbHHPKm0Yb2hwuCfgvF5QIso/8gfGxYSFtydTavQ5uX
Rat3o0gYkYOSSj0WCrDFdYvBX22iDM4y7ao597haUfBHwwTcLxLC0wAe1VDSDKi/
2UN0/ys6imLzo3fToVUuBDsG060TYFeZ0Ev0QavTYD6w5Rpv2l7cTzb2OPaS0ICk
Dzh4CBJYbzbuZbd4gpNBQvo3gzOM1D6FuPSC1DlLMFoT9jX7vgdm3UKYCqWJ2ePs
Y6goJy/v+WCaR+frK3tS6frXVkEqnyyvg5+qneGl7tJ62i8Izq6wPC6twSAkfBxX
VCHGqcTs8XPwq8FY0BuQFeLWEibRmktK+nh8cWD6Ibsx5gsj91+1tK5csbxVNzg4
ejJaBiQpEhXB2jiWlZ1AD6GEZt0NINwba9F8v+8qsGuHcGHADclVKz6V182bIxPV
ZAQZDtGD7ysWFBYSNWJdUEmsXPhLgG2MK3byTJnA35WJ59PEV9WAgd9nKYdfV75c
NjPEBbU5+CNF4msOCw9vSHAwzMj0aSaipejhc8FABzk2wEv87R6YCE8o0ofoOp7L
epcgPqI4NhrWvblDkcDFZwQOy1GkCgeZfdOP5tjhP2JUnmx+n1GVjkrIB46t2C0e
KFmoOuD1Nl7vi8+IsBIa+iwlWF40KywjmCfHMg5hNWO6bfbWigu8856tMOTHoB4Y
8EmavIh51zEANChI/B3K7nXlf9wF6GCaoLGIxLdrmD1daay5eqwLas0xa6O1opKe
ZXItSORsR/94EWlQmsxUe+kwuNwELvfjbTbAyVt6TV9xjoET3XP7HJqzLVrc0i2F
/xZK4sjHdBO5eqo3S78EyDvTzk2yBm6lHGXzMb+v3dLiz4rr/wz1MZHGpyN/9e5L
KUaGo/jGdoMiaON2KVRymbN5tNmX+lKTI8rnnTNTD4IftUOX/ZnN4rGKvYoJdJTN
kZX2hvk7EJERupyfVgHwxngbe6VbPkaSHWb9nhBOcFf4h4wNjpAl9u60u9xMpBUN
7eru4eTMD80StCO2w0A0FrQnAYVrs7LLnEyK+waoHWYHT4p1rvb3DYaB0oSArv+K
fxFtqn8qr0iM5P01IO0Mp/n/QIuU/SArtpn5qjto/Dff7+T4aKTh7+D/w84yq7vy
GSGgmA5oilRtxbfsrtk4fuZpWafiCz4UTNO8BI1P21V1PNHEqVpa9Vea5bkzA+e2
47zYrQ+DEohQhx9DkMP3L6wGob4X/BXqO+t3kwyD5UB+j9YeP43QFXqe4WWruqYM
OYyH4X47SKSDydHHie7VZ6exz7T0lipuK5FZlh1G5qUuBFGTYKEnygTmWirDdRlw
TC3gWEUxiOjR4BTpqUUtxMDui6W/62DEniqOJVMgwpSJvZh+kgBKMW569652/b5d
Ua4L6fLUZPINVcZK1d/FWPI/ouv1y3t25QOfbTt+fdsagnMdYnT7h88RyS1zg7+X
ZAJTNLt2UPYjklugEq8sb9b4M5fOpetLhLamUAiK+96QlydiuuTLZICTYKsXYqbD
tPD+Vlruji2WIAsOIABXvaSY6QZkYXlmLYTW33IJa17eZ8iWlSWcctPR7jfC4rVY
fVEqthEj3+cTPg6VjXTHcdZWbyXGi0jGgtp7Wjfjqdkx1FtmgqeRihUyeoT4VAI6
UaDYqwcHCUHqRmJoDSsaX5KuKWoJCoZGmBvNGJb8be1ucTqNxjv2PdJspGE2KYy8
IPnXboMUKKUFKVPO0ezHNbUZ9qoPCVccivutNHAPH971sgJxas+TAsih5YJsSUCz
Yu1jQfk/cclBf52vWxccIsnxBJmwFmnyFSfUWa+AiRxYlI7eCYCjqUXrej7XaBPZ
ef5/5DImm7E6XGaciWF5+GLqxJ0F0ZWOWmzS+lZNQoHPX27X3mXILnEdK4bQOI2t
RzfPMIELL/PA5HhxBiytBsI9sj34jVY+F1hZt6Qb3eItV9eWrz2/o3Nvkyyo4/vX
erioGGDahtS9noF9oZSn4rSQCKwfnBN+LkDwBtGZNLxtXyqCCxCWT2Nw8dlsW2bG
9HjYEUhkyCIGxJO5dnddOzxoMrC++/SRV8L3mnm+cTeW5IguhpNX6zhh2eq/RUxv
XfVhiNVK0TcaiQnvSzSJ3+4SQ5t9JN17FlmlfxiKhPVKREwmDQeo/1vtFx05ApIq
8B7HyK+WSa7Fy9UiNFJhI+1SZteHL9EYQa5ks99tylBH4zlo5hlY6lBzr/2LBRRe
Vjuu3LAHWOGl+goJwSEq2ZfmPlDVelr0F+IOzYMUD64e2W//FkBsSnCLdV+O00aT
uiHb+6pLsDeJsJzxuuzdbClCN/OwhOMA90BbBhn3AbQLneUhu8R5wn+S4eoqjnoS
sE0sEP8hLNxsJQWi8oFyQyDYOhX16eFWenx2DTpJxPTJxiz2oE0kPe5IkO4o0IvS
Z2PBchLCWFUbKaVH8aOUaUVfgj6EbhNbqNjwwsSUbDe5w6Lw4yFkYoHgAL8ggcoz
ZNYzhr18/os8IGGMkXp/47mlUnfmqxhtXzKyvfKXj4tIbT2Yz9IHkJTZJp9/lmUd
cjKWHEPPH00H9ck0VKqu7pBT5UmwCTOr1ht8zmkQLgEC1pqpDFAU8DxkBPx1fm1B
qsXUjLvugk6y9SbNgBq0s+usgkwTZpXJDKhF2qCR7qwUm6N31GUpBYIQfyGc1keP
Jdlx38AN/fhRU7oCOGovN4iNJW4eraQc51m8cqXKD+XEQZ1VsU/BRa1nQpA9Eaxs
WfySAhNUZnBYmnzfpVLRdd+gr8eiIVvAvui3+VnmLtG9Is+NfGdhmziYeCa8G2l2
HAlklvk9br9EJitkVZFuecmRqOE5n5cSowFwhuqPWMOiVRO/9nVMBW3ptZxhBRsj
6SiqN7jCjFztNJ1+kkUm46wgUqDdvsCG6lY/ZPPA8i8ITOZIFfY5D3zw+mn+1MWF
GcNtmTAaUlHr2eLcoiaSgIc6mQx6Yk3HX4c32vrHDEhZNADNO7gdFIRRYa3mimOR
MJ6l1YkzZsklZBqrqnS3Tj95zMV3bJEXvAvwrOpFGqSZ5HnoPzwekyUozVCfTVEq
LMAHOX4KeJgPixBRZWnxTNCUWmDCRx5EQqKLE14Q3ztkgE9O+h6bkj0GU37JXBFF
JWeMseOKIZVJrUemD4z628vKXaDRpTAjNuVyQRJmSnuENOHf7YADNXIiIi0h3S4F
pwjoSIi6L6QsfcxlS/HRdAZ7+6hegvkTchn0VFeuRnX3ODY17L6XXPi/mjxa6RaE
xXTvcwv0SaHZlvt1ecSS0FoOY0Lr1OTr4njz1RIuCH5emeIxJvuMqL79mwr3JL6Y
1iuJmkAIiG1Ty2ChqAoMdnxp5QzSpE+jDC+DuQIVnBEbyG1BYKOtCmfR0/SqGYVQ
DDJcVQd0knS1yIeNMyDFjOHqMU9ZykQSCR83t5ClNMFKMiFn/Jo9+lF278T5FCcd
0TWnJGrT1b48++NfQlLP68859LfeiG3ArGImhNL3g9RPsfeJIfks5SCSI6CeuJYL
tJwkqO0BN3ZFbQY057omExFqTBrrv5tIttPzw36TJgWwnBOcEPq5MLxRUsKvvfQc
rAiRmNIMVjeND0X6JiOHwqEpBaijfrcCqDaGnlEZ72fWjmenB+rHYNP7jHKbaqDB
WuWD0KEVW7vpYTjG8VHN9blAEdZ3Xd1IRcmd1aqaokeiGdh/44q0DubxGcIbaM9E
pDkNNME0h1gswxmDFtnlkcUupgdzq6P0cf8NLJOI3CLGNRS5cOS+EGfCJxY/OoEU
j6DpleIVLdOWriAa+rcpNi94s9kqY6MLhRqqMF2Z+wIDu8kLRTny2mfuptrwcIIw
ju2WrMsrhUuOA6p68FKMFBqER1djwjwHvKAsZ3Yfnz9/duNtMn85DVJZaXvervLB
aZ3ehvC+8zWQUCCdT4vHdLEdoxTqBK7YO1ex2uKa9E40wqYMxIKanxZtKe2x5yfT
4NsuzC7wRyrotym3s+MS0Oe4zKHTvQ6oKsMbp/+ohGNZlX6Rw0+Z0FPex1kBnGGa
Ft0rcg+j4IV7/ZBr0zgtMMBhC1wHNyIjvEKZn7qJ2xHs14oEDJyR7z8DjgHtWbD4
WUoIbmbYHV7/vfMWRda1udZ297gG6jcfBeGm6nmfY77ETZ1LOyisr/rnbIjE43Nf
KIYzOWOyLgcYY8EoYFuZUSseCcrnjn9SjjScCsELtJPFwE3bdcW87IRkT6DxsEZ3
H8gIS2XtutWcRXEUE53zMr2A/zAbBXUGY6xmDcWB+R2MCmhHFNqf8ENE7Ry2fmed
1UNonkFN08sekX7mxhDXAIi0bzlx4yLlRSSnxB9IWbo4qInatRiuDYvkK3GY/O81
OYnGOawSUquS4ILawkS39QM3OkcHgUVSG67g+ydDbsxLhfXyBu2ilOj30MPFSSY1
V5s02OZH6rWxnHyvXi6AbFZT1Z+K6LJFX8GZ6LCZNo1ERCsXSgTofk5Sb/nC0Cyi
DBvB9H2KR49a/e9/ZvmdhiSCnmkYr8cqK72lNt7ZG0io82d0DOMNDcDsVIUcVANV
ysogkfgAxhI/9Fl95fxRjWzsH5gQLf5BwmtTBFphb3xhHMzszizEQB0ox5G5tCqi
/142lqa3JwUaq3F2zuPXa2RdJVCjoJAHW4UlIzszK7V4tqAdoutfuyFP71BokaDy
8vxE0wG6eburMSXc/72pHuEYjEOdMA8b5dcCqN8SIruVzp8wsf/xSZtNk7iTIXbd
drmvxR92GsyL3xd2C7p82Aut5njnZ/aEzH3rxhRd/13tXtNXE2uNS38+5/O4udAu
p1D+JLhMa14DKFqYH7AnfpKsMy3op5l7pUivVCYPOuLdiFNL4BEh3/qTl1RgRZa/
Ic0ZTwAP1xtxDuNogmuhyPJXWTR3opVDHBf44ya6MC2hDYUeVJGpvt+O1fBY2NbO
N61wiIZ+bvBT/ZR8WRJ811s/CkrlZL9/h8tOi1KRQ9+zRhUJmB36A2kuOPvgXDjG
H6gSqzvRoc5KAK7FI83LzKrpvPUlsUK8cA0qv3wSOEwnSivGXUqqYXIFo7fztEOM
8I/ppyigIRVT78vnUNOUKs+vIUq7hnUPt0G4vDoyH+JGeeJ+Li+LaZIk2fuj/248
1ifkG6Ouy2rvpGH+I0ClYjTTJFnKlAZ0ttyECcNsTzSs8iwIt8auLPHmDURGsEXZ
hD6t1dHuC2kn1CUGSnhcvGy//nxdz5sp8J8mj0yTXpMuaPkAyo/NLeBF0Zc98WPx
Hy+qYyQBNbdTJLuhHsIxDSyy5RZOxkb/4iSx7WQQINRkHgFzYhsLGXBw97gB6B3a
PN/t2W24gyfLjfYXuA2b7B/jd84FyMYmZ+VJhvjuSeU+9XBU31/rGtOW6kC9Eif/
Twpba8A1wdpUQXaOFZLFi53+wm2k4AO54voKCAOVYWFxG1PdT6Km3BDWX5vVzM19
QywZ1oQD6LOWXiSr3V9hoLJd+9fBKaS7yjin8pwwXJDNm6tialYrkK25MqBNXm3e
EIVIHzHs73RGXSCoHtxM4EhS/blsKdb84MQZnWWc1B6s45znHb3LCIhfkkBpIG5F
v3Ozj2aBdJYKYi5r+rrsGy2H3JTsvG6pb/gWPuQwjwCHNO3vWCw3mKCJxW5Xn9pZ
CvMAHiC0na3PF2I0uK9KAXYqvGuVJtnXipvw/Yu3KaIQmpmv1B05iXJNQ0uzFCQ0
37bVTgrjYWIn/i21ntDZztlaqD20T36amuqJ4Ff/dHS2zHcRYywWEdqt5jQXF41o
hv/1bXPutHCnVZ3XR7VEidfN/tN7akNjvKqmtIHPMPHlGqMoxj3wv0bEaUyWpfJD
e3pM6+N+D7Hb7CNzY/cyJTz46X1eILm4oOw7R0hKU0CmOJ3EHSMiMXEqXBKscYW6
QCUlhetvhhypUlyXWSeDjOGbHLP/fEkQcIkckV7Br7bF1YPxTcEdVkxFmbcq8zKx
Mhgd7GLYjOCqlJjIPks2swV4B0oc8NLG49uV4FYQ7RwceDZc61tJAAU6mXGcS0kI
OK1U+g/00yFovtv4+9a9CKwKXwo4iKIg05hdnfm1B0BOp8Zt3GG3ygFXv7IFQH02
FL/xEoHSEDUa50nbEUWSHzED0FPaVRbQWqWhiPlr3vyg+lXKyjmku2DbHV/LTo9E
GpRr8st3dQ/265XcNVpJELk0U78XZWg8aTUTDxSLdBCeqfwC5PB44J9LrwR1G+FA
CIl4Hio+BTIT8anYEKhFqTxRZV7R6wTJggBEyuJnFeZv2z4ZQ5Deh2cM9sJWyZ7G
crO4namUOgmTm9mUiSO7rCqlAWAY3M8jPBnvDoH473lqYc9ZpWX1PbdLEpvrkqre
eGALxoWWAhd9ef7iFehMyNXMObk01eaxMB/Np8EGU5se2B16cpjN0q8bzHlOC3R0
KRjXaCKt6ME+uL63feW8qP3VaIR0ClVfuU4/fnxKzy/YkmYDmROflQtgpwtVDFVX
UOU042D/OApuJOQtbMfVvgpEqvofMn/eIkYt8tURo3EVDWoXYI6yvOwobA0MAC9U
noCG/hX0kbLDoYVkrTHjwA3XfrdbjlEhHgzIG9zPVdkS1TNbt7bMk+nC1Ag/86MO
uIwmh5fz10EDUeKN98Dn1yNxI7rO4gwSB6dgvQHddy1Uku+jKvXIGp5n/Xq8wfgz
CKVDnajVfJQP3nseevsakiRkzjsdT1lCHBU2XNU/veD7aaVtAXxHlONyaGIc5t0P
YimNCQgpjuAoluLe14T5JnCve7qqT1MmSoD7PBFEJfjIjKE9R7ifbndGUlexthwd
JFMv6TogEnUhjyzdEXvLM3BbRjxrc0Vn3AEy+KCVoD6NCDC6VYSx+qLMpia3zUj2
S/9cLe6JNh+zSdIwVtDiEHRZ1tytoAcSnlfr9qxRJbGvaOaTp/5cfjiDfoDKfC0d
+lpnVWmVVVeChWErWNjiUYMogAWoX4x/j0ZrItBuio915Y7oTPzJPZa/cPptspD5
/s80dNmsq5DasvfPMFdRdkHM8GyQDBdos8ZoWwqAIguap7bW5/IB9hflVZiYVMbf
f/T93EraqV0h7v/VlzYbXTAAXosprDSiFn6pfkxHQm2Baygt8NyKGmVo0JieApbd
j5ioqgAUKeP2cZX8Qrc3UNZ5CgDND9pnQ5UUFm2z4grILZUY7q2BRQYaM5pPTRSK
00srEC1gPSfljvw5G7z+3jUTVql0nXJ1/5vdX+LGoDk4NRlRfklu/HoyWPBGVdl6
BcQMqmPLymuJHoj9++uLePAZgcrd8KHLV9yWqKjUzYublrZIIJacLliMegp9FTxt
j54kEdHCJlP62l5bW0PZkv8YZEcBW8ahI07W1minEr2EmellHN2jmh4Puk34tpq8
zJIpZCNXhz6dIX9ALpl2dV73dhseqIZcoCOqDP+NkgtXtZL5IGyaoPtA8U71yrUA
wHzp5PqIMXvK/xIWnYUaetbYAQIZHb7SDohrnBBFx4tRp7ZF24CZPk+YFDrCiimv
i4AxI0L9l2nx6sX0VFQWX/OYlYSaM71wZ5uEcmAJkpo3d/OsgFGg/XLLqn0RDV/J
5namdbQGCUwZLAVsHURH3HMFrZxShNpFk65Tpr+xUdPh6zY8bYJEvX8PwP2RxAg/
rufJGxxHAxYTLbQ7Pk6BCk7C99sR4XLkSIW/g6ltkJ51rWIJ2e3tsm7oHqm4qPk4
7FtH37ngZ90EEHtlStTM2J2cwm3CINkretqzmPfPOHNQK678kNFFsZi0c3qxsUa6
OzpDr/JbAEcOyxFwQoAwwX1n5Mxn7HtRd4XwabM3Pi/zRj8bkW/RoNPgRMlX+/Kx
Ncm7JBeIW/m7a8zCwPH+q03Pi87faq9+Ni7LycZi0f2m4WxJhz+NUhjqjRuc2vrl
xNOgdUMszAIC3Q/4IQv29DaUDyoNAUDfIMbgmuQ1yEstrEzvqrdw7fRyE2glOAwR
WxdLW4Vw7rC9fjGGziPJ1vJ21bqsUiIEpDORnE3u0SHvTBQb2SZ2Px0Bkh6rqB7N
oRs5zkmReP4+dX7f0mUZx0+HTjNMGO0ftdrqoIwirZh6H5MQnoQrcaP0FVTeGlMP
AYg9nfOzyyIqgYXe/K73lY/quBnoMT37aAOqDuCtm4JXPU+fgXsXctE8GIuFSaj1
pYV7cboRU+lHToq23K2wOKNoIoTaa8tWik1CntJhgFcwRBtUEEDcD/NRtlklb2rj
Ib0zHdxmxPDvJe+j5qM7+qqjqOQtu36WU7OTUaA5827vGPrbTEYWsydkAMzGggJ2
dK3nl19jchc4wWd38QEsGgY7gNblhYmRjyCurlzYLlrGnk8qefqnFVlhgU24u9JK
ifomr0NbKqvplachKU62AtzhYvyyzaQvyXevxn3qumVBDem0CKcW9ZDTIOdc/Znz
`protect END_PROTECTED
