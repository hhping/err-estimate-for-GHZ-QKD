`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yiGOkXaI4ykLv7vhSIgxYXZLowTI2ll9syrx9fpQVtfvbqE47RK0oB/1Fkjkql6q
/aKcXRBhPoXo68SAL6fM3dkgxLBApyE+pPTmoguHvYctOBgBdJeL4thpBhGDDj6i
z6m/ywVBcCyClwMcWuB+vpRdNZrm/FdM7Ivx4o6ct7R7q+sXbuUU342bqCcUyHU2
26ZHSUzyVFQIdl51+c8D7EXhXb5ZJWCyWs0od6BOwVDTSJ91DVPF3yAeVz0jWh9J
k6SphacQ0YXvwSlRlIHjBOfmKvQ2B5I5yITvF7KM45IHxkrcP6aUC50XtBuN6u3M
X9pauL80dXKtDvdrjVousp7bXjYGVP5io7DSXEgyfkMKHhVE08UZ+6wV47/F/Zuv
Ng/4pwSyAPyF4GRzD8z3+mRVmUeQe92kYhKnDFzMLnBqLj3jyC+60uKO2AZ/pUYi
2K1l157YT9m7F2RWYo9EAwoR6B+7+j5w5741JS4gNY9afIoYS6dKtvszQA2TkxnS
`protect END_PROTECTED
