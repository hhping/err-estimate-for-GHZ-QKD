`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
78e2wlSVCdydukCGofoNXhiAZF0y7Kxf50ICxRK1rbEUmk75EVusg7Xd24M4f5kj
hETyRbLNf6COJdCwFmQkxNbAIpizKoJcjDkaEjJr746DPiNKSyyBBWfmDk4bY19y
H+LVFBlNuuAGTY+iOVy7O/dUgwB3uUmi4DmjB9BRbr+UWqBPumtKAYVdRpW/SZ4u
b4IbpenqmcctHPwxPR8j90O9Vv0XFEeaJWgJ4sgsxOoli8+Vw5KHKcU2cVJdJQKB
hnqCAnvFcoAeuyk8ssXvXudissJd/Y/m9g/h+Ykff+x/o7xXl5otyV/mIwCjnrw9
Wx8D7sCJ5sJpM+m7cjGAqJno87VHCFps3UmB4FA1W8QW5nBuA1tYf1cmIRVVCUvS
jnKr4v9FNU3Wg4XxUwBvyMHzFwRcTr3z7C5JWVnU42Ktqjr2m0VFN1DNYjJH7Wq/
NvWOiafgPsSTnLkl++h7NJ3/yA8oP8riFogrMxMXGuCoAXxZJkRQIkYCG/08hcOz
039EDporL3a8lFLWu3fIB1rL2StC74BWbWXpGetZ8i3C5pPs2zKJmqPKoA59Nz7x
vnFnBl8DD+hFP6wFNwrAKpefmQmeMBAh5BT8UflVtjlXUV80DW4uD2jTBMsrFjeU
zQoe0MI1tyMlZ1NK6cvzyC3wcoj460XWITO0R41nOxE1ApehC4sx9zXbMQSyxnxM
JzmSOZa4KxzqtHYcA3iX+sAWBTY+wJ0ypCQT6XH4Z/0UmJTH59XywtUoLwKN7pAH
mQyW9PtRDIIne4Wf2VzmSJur0H/vCG3LwJOGcPpwtAAib86sChfyLinEInNRzTB/
8CRZ/69FzGWlI1ohAqGk53+FyW/deS3rTG1M4FAhMXgGyfO4nnHNNuX94soa+9gP
dID6LSUwDMfgiPuYq0AL9qndePLT4cpIyiUbax/mwGtgcYi7A7wUSASKwXwNwAuH
Q2XxGBYbDTJqYmb67IdOOiiaXoUDIMH1QRWq2YUPYQN1R3aSSEN9z4d4rpyCd7mt
ooK1f70UnF9Cz9NDaTw4XFczU/oq5Fy4L3StUrGqAcO2n4YicCi6QZh62lzJwFLW
oGVSyNMHpGtPk0M3m3Ck2dyPOgZOYFZXP8IuGpzYBlYP25mhmjh0vhm8j/SZ6eCJ
FPZCk5RwtcolodnpJDKOsF8qDcao3fDdyUiraEjHu493GkuOCYLipVIhOYcmoK0P
6hZ2MyFNjq9iVbbv9z09cgY9r9IjATQV6gVA3+s+6d49Hfvn7FSJXTbkQLmL9JO8
/xo3RFiVR3g5h1PNwK0NqTcCdPSKP4dZb+Ujr1Rv6RN2Ybz3yOZY3wmShF9iOv/H
7j47TlF9BJ1Lkx3Vgn+1/qcq5mfbSSMwQWgFFJJrMhAl1N5/ZZ9eGyd9V2Vi+2Gt
N8UyzbvVE3CMFK61jDCMyjbsC1Ue76ET5P1RD40K39mYxwhb60bnpCuI5WldD32c
hhb/kskwfuxZH8DvXx+1WXIqzX0KhD088MLGxVy7k7BMKANGS/x41+XEnKhrc40I
fDtf0fOz0+qwawoXYsuHV1sfZm1JmTgSbqFiG/RCREdHJZQQMXRKE/D2mb0UcsCm
OsEZSaf07xAl6rneNBv6JHZRczeWnkNFMe3A2rgXyFA7C2EPt6PGoJgFRo562bLU
ZHB9CwjxaZdUh1zupnJ2d5yH6VXo2M4jDNeN6tHLkvvsh4Vwe8a17GXWfepzRJiH
nfKEEiqxKW8y7wYd6w+daetW/nHNRNix1cE8mxEvIyGOc/hyy8qIdIoMdGuqyvcs
/ukOtmGAv3fBS6aTrITZJ4AtpF68XMekUdShf7y9simPB3TB3xAMuNRJ6KBd+W6v
2fD9xHrI2QZlqu4MRTKB3pOwUF1LECnKDDRNPb4YBquZ4djozMD78C3US4SG+FGR
OlG6UuL1fLLNyJj/+QUC9kPM2O3XWP/e1EMTJEh0LCEanbEWNAGujKn36E5opRse
LI0F6dn15Wm7V/kWO46mLCqNG7r5by1BSEV6UUs+ok4TAlTtgKi2hGwpbmC2sT7f
BguPKUPatxcUodyIOSDEg8kT4x8QBVKlFuUmIQl3J3zevxP50rgjLDn4iCqRfEZb
ogwjPZBkwrUwKAmVB52f96HY2PdofWFyZkDbfHrYAJSBFEUg9npkoDqD3prcoyoJ
J4rzOu6EsVyo8vIiQVdRb+2bF4zRhIFiEvJD9esfzx6JV+Ar0VdXG70LmQD88YAN
bkV9/kdv9eTUJhV/zm9wSPXgeiDRiwVhTzZLLUjgnjtOFZQWhiei5uZb4FdxDwGw
jng7PWo+N4xU480Ddk64Z9bhtSQ05dg7rP5KhRHivGTsnUH99IeraktKkbCAvCdd
dkVFZifEAyQjdKu5piJQ0hRXEtd6r+uNpUviDLXxKPcnEHOW5S2e16XzwM9xCBQR
Zjn8TaiH6T4V8k6U1anjV36vbfS2rpGRw/Mn3ZIzujbZctgUNTK4yixi5lDXjxZ0
cUfn05tYxa07gZbHMIwN8qeLV7jfoyKaIdTZOjAJ/r++fUd7oyi/DPEQGjRK6wmb
3G9geHrdoxM3NXT6DwoqChMyzVaNCFEusJl9sXnf3wNcPTmq9LNauSyVxS8Y3ZVZ
UEwm7i0rzJRVq3G1ANYhProWa0UiGsTsszjlefXPQ77QlQ1SjrMTSuWUTcYyC0eT
meR/kDMA9Qt7biufQqcHvPO+Xchdwz1Mzv8R9Y3cmyRN3MZbA8TmCH8GY0DXtUJX
KOOBX2lmRETp6ftcR++naTxmvLeeWVOvLiw6xXhbwaXTY0LRWYa9BRm2m3LEfSvb
OsYt9oCURIRzDU0GiRDGLpcroN+v1D01+mYPCiEtA3rPruYC/AUwgzCYH2vpjZa/
ETaGcogv/I8blb0Sz8mk2SUKNVX1w9lerhQJYhV9mLOqCt2xFv30ALbLfJsPlvOj
ZsRhLn8y07DSEF5FpyZ35aVa6TAx6fscxNShjWAN75hZPZDTao5RcYlhsah8Gi9U
m0clbunmmOK/qvmU8F8tKNC5aa0DEOlzEHDUXgecdaYm5y1WaHBqBo+maERaK+pD
nFLicV4PIXP9FF6kQ4IQouCPgt1w3HR6Q3/jaFwrNeyZm8bNVbztkMOOFKhJctwu
EObjWvDnMCMoZ/4XubJ2nqIbJzk4ELPo7miehvm1WlKEOKVY5aOCOX9e9hiwvaJC
SRJIT2fBY/iTONRir2pdWJrC3oL6AeAlzdGybaeFCwecPsX3MTg9yxWFzHM4gcJk
aWSrPftuFies1EM171hG+huqMtZHGmLIHrFiodJJwpSEE3qco1Qa8mFS2G1cwxLq
NEkswaxGgue1FOXqTKJQg46RI67C9mv8RCGQif5m4hJA9VarMaMO7xnpWp9cTca0
0whtE5nees6dz+liLjuWKQs+vypPxf/veXhulFz5ZgMYdJYAbKw5HT27kyp8sYzE
YlrckzlIDKGQkevz028+7pnvYvoXVflUd6CgisdiJac0HOg3wkEFzJWJKSlCkyJg
tbplgsVLVwZuajJRJuA6LiPBCagR/Dgb7JifLWblp5nLoc+vdzgKzeDSrwTqQjwd
XCrMa9fzcdLAHuEV7gEdOMvPU2QNXpV8IVcjf1ZnT1YuZUNEaJKT9I9Ny/RNMzeh
KR9qU+qhmI71Q4Umx6tlzwhzbmxYI7hQisNZIqDIx2QsHHXU0SjrdGLyrJgaU/uz
uTUZ2mWS8BBlQWAdjlc+EInz0aF+D6E44otXeBFdNx7LFcZ9ibQT3ks/vChZoUvO
mC29lJpba6G95YdDbllhIz1nbClP9MeK6gOAYxSTmDyqQEVIj7nTjtiO6SnMdgl7
Ph1TyHUDZMYavAmuuuCqBU9JbhvBevvDPidbI0d7IdUxvA7/ZdAeCaAKPt+nRkth
gxBUqyXtoTeu8M0cKAyqBKVYuu4O8JMLrzvEbvkgg67V23cxg4dsxj9tRRPIQaYz
jrqFRl13wQ4h73+8WQ36L/vhgpKUzfWpcs6Pwpk9r7Hfz2mPEOCPSN15QXAprLay
9J13yeqN+kRO6F2If8caPXcdwDOnOncwy+WMonAkyz9IEqK0AE08b8nWbjwyBHq1
OTaffajuKa+bnC0HZiVrKz9VxNxBqvYTEy38alynSqKmT4bXx/Wm9gpNr9W1y8Te
eXKXc/8Nb+6Zqab8xXAvunC0F0oLpR9qiZ/tbtM4NvaPemAWpCfyVoOEta+ovQsz
doWhQWcdlKjWBmngwqcNOr3Zjn2xNLromX9pyyez8AKNy9XQLuBTfM6IxiUvboG1
weMAlf2mXSmSeN0eAx4ohYfHOppNz9KwZ9/EQdwdo91WNY53EYx9b1y4mdk9X4iG
BSBR7cpfLt1Bv8rs292O5iu7Fq8FAlxkeN1Ed1OrDyKoHqsr9bLtgEBulUYiD6Hr
z9tyy4j1yg6pnwrhRIX2vw5ZjhQ57iAxcy/1P3DJ5UZT/jMediT5UafQE5dO7Y7M
Ryc/tLWUkTH7oidubbJsEVIwssZ75OFOI+8u65/mmRw7wwfMdx9xjm1uBf5+YxtV
24H1KheP6YEEqgY2OmK2YmFSXeziN9LPC+2AtCtGLin7+DXGVoSn9jM0/RV00CyO
xksjPwVyn7Ry5P/2JqAW5hETKektETax3XrQ+jqPAS9uwXsIu58niRzBfmERka66
eHCxjfZJrldVSiIXvNN57+y13jMxzoevk0fFMXIyJTzIH6e1OUQwjQRwbbNqxwIn
zkqUGZDmXtaWiNHiAKgYtGSnO7uSIZv9N/7VozLm0Hfrf+5Q4S62xjS8z9/C5tXu
Nf+/5IE0/lF31YIvajajwaplneeF/BvNzpnshoZL3RI1Kcb146Kb/1ZKaIW3H+vR
8j6gy2VOg/38b28Of57MclbkYJWFctBlYFAtkifwUYpq3stNLNwYq0IuQMOEO1JF
k9FZbqqX3BNAyftVAlVfUICfEJVLouvJ3fsE6l+3uoebTK/FJ8iDoGkNrqnUy5qQ
phLCXlOqlkU4l22eBKCoo/llEO/BzMsDxF8iKkRiQRktPDb2WaP1N8RhM53ZMx76
OAVVm3qU3kERJG+HdYHOpRGBhfsdoXw6NhB7PRzbwnU1Uqm/OZnf1eLd3/Z913Iv
FV1hnA1b9boCDk6A9FedKEvppXzygxl8fESrzjS5FyG26r0IRrjqrBXjkZY0PfRv
pgeBs09KZmt9YeB7ZkRmA/S0lxnzNgIrAw5djISBmhIDLs4Do66pr6YP3o0cv6a1
MEjUJ9qg442gUoaYvHYjRclfniUXwKdCBLabqROCh4MZBg5fSkP4uD5+DGqxpxph
qfOC2GeAL+0k19EQtWhy/xNiULQjFAxs+CJATp6tmNKvsQF7kSObuHlsmTk7ekDE
DFxb4Ed/BcpF9BE2dlX1XrlTi6QJrEXL99HVlqw+bU3NRPw7WqZv4kDe7Dv9HdUg
TgAmm46dlNt5PExYAyuJF1eEBye+S1J9uMOCMH2cyeTYaKBbdb3DwHlhjbLksb6w
xDykA0gb63KqL1KEyz6bq9v/C9xud4Xh8aRDDl4Z7HZFY4rWVdw2y/pcpuKWbDsg
4lKuFI1k5SQoMzgUQ8ZheM0BsnkWSw805kS3Hx9bf2nK/YpufYMSqa3dF4hPyzyF
oyeH+4Fj+RJiYkquZP4fj9DYQew1XXVHFMG2Bq66t6Y0edpWFG2L8jsZjUZWmyVb
J0zbQYmHjyNMXj5SA2HLlgE03Wq6ekKisZqERthgXuadtkwTSUHpi6EjBNPljzvG
EHhPGKDe3sCQY6cbiekGHQ==
`protect END_PROTECTED
