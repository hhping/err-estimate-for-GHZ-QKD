`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bvei6JHt1ANPi+y0n+JLcfZzzunMO0zIlJ/iQrv+J6DUv0zdMYyB33zv410IpQFz
EFBm0EbLnNHR2chInaaGTh6iDgxtBPd5UPunkFt/iXrWjyvDEp144IuU8cAEC0t5
xdWA8+wZa1/wLXk4V6IpUOO2NcvE3KsuY7CXveEQGh3DU4MV/lufJaWomLcuavKx
viXUsWBVjWaFgxK4hdtFc4fU+sTd8HT4Zt/MALmT84OldLTk26KjUQId5F8NAo0V
vNLB/5gyVaDZQehDJj7RSUtbAxJ3kESdfVBRUCbOgEt/nwxoQwnu8T6ZylqwARds
wMRIopkhZrNL9cUXU9qV6yIMvW3jLTGmmTj+F6OYvo7EYsKtvrHufMed1hTJ8vz3
O5wUW622L0h2A3vGWhu2sFHvV3fLtGUgMr9/gFIxQpD0PebTsycUXbLlzQWJgCvX
BXLiRC+IY4ndlS43smZE6VJMQSu3RcYKi3S+TeGSD7YptCCsVftsOQJJKKSOGBf8
rHCIEMwdxsrosDZcVHtQHhpsgPyUUE6J/t65xfvWSKQTqGgT3TLa0Hg7QcsmAO49
wT2rOG5ID1bVGRu/K+Sv8GcT8+uFkRMRKu0SzfDeU8nHMC/ZwVjhWOJ54RIvIZ47
9WdgmRlef0lxj6dhUpkeMTwLjfseJXAYqT+2q5Alp4PyLTFGzrNqVJ1ScWtWV8EQ
6aOzXPooh7STmA7TaxokLsxtX4WHUyg+cSQVjGe9y8NE56XZKSFbamzr+64DEl+A
3VGu7Hfv7MPjPL/YedtqAnl2HBDlocQgoHGXTCjIa0g1YC8eNEf6RCPQD+5oqJSx
PSxo0UMYqc3Kz0Jj+us/BErPJeTZL7slHsSxKSLFU1MW3ibdegvjHAl2U1ipEh67
iKD9XZdUwPj1jGXgc0ohel4pS603Wk5TRSWvAkUk7N1Mq4hDM59XtZODhjV+hzol
tesQUR5siE1/Iozang7TkGIyofrs6IGG/Dc5rlDXUmyZfHqeZT3mwngIu09itTOb
QerQQ6mONC+rP7h3RnZlqY1QcIROdfXnFnKmBAY7EMKlJkKFiYsPKbB6nOHwmU4F
sL45XFTqzkKpiEyLZYM8uzvA/SLg75TAOG5ry3ZWt7lESN8y9+PMrrxetuUmQPW/
nruR+NGys50gxh4tRxFWJr23dkjDYqMXmmqlAWHMIz7hxZPGoWrLNWeYVMuz21rp
JzL8RckaZ01MyARWvy7yejgN+L3LoRMVWZyQqQ/5K7N549aXo1QxYLHV4BC+yOnA
KXxjkj/gqZFZx14FEG6podVwGYiD7OB9iy82rXM6pHw=
`protect END_PROTECTED
