`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T9z/KEYpfGobcVE88SoGfH8vhjV+Z8v2qqDiy4lymJTPX+yBUNdfA0kj/ZuZtNrb
FWkLReN1B0W9Ns8ITnZqVNPD23Lw+j0rbqlynBrnV8ztsa7WqU+OX6b9ig6WyjKa
s6d/uk7t1/3YiX0q7pXKQUbKL8vt3ZX0t5YznG34lCbiElauULde1aVwaPnSRxqg
17vDJeJlfvYeQhteje5PEAVn4LxhXSKJRWV8e2Cjnz68wLXZN76DZrcYY1T+qL7x
nLiYmGs98kjAcFJRRfabqNazKPsSHEXW3RFh7cEe5p+hiYr3SEDfm/m1ALKlAbBk
K+7dtBwXk3NDMm7abW22EJZdm9gVeMey3S+tfi2oX9sElXZfo+2F/v+FgU8En0jw
5pbZAng/EQvBZ6xs86xO5JFZULXY48a+ytgD/w6C0AnOXLNhhAXYwU43wbyz4p83
OL+5NAxLT/K185MbsxnxS9UtOlEwG/H/oUnhN7UELa0P2cO6dgyIHIuxBmEPTPDS
/7N1QvACC6az5IzriPRiD5lj5rXVCYxMZZI4tX05DGVYCM6ee/a+EUNxEmwL0Vnc
772CgyEYcACpFnP3qpZzzG2r86QiVHDJ8gSGubCHiP+Tkev5ywszJNbWsWDgpjKi
q4uE9Zzde/Ctjo+RJ/D1S7/LmIFvI2iR26/REQakqYsAhvzCTgS0vPazgo2mGJeO
Tgo4GIyq+wBpjw2M14XmzRa/ytK66VQ0Jf7cqzkmNDfMQSVTIwpHviTwOOnG1/Tz
vEnqwt47FGrw7hDeAU875ufPvGKonxaz0H4aER1EgvI=
`protect END_PROTECTED
