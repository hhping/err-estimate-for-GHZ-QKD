`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RDzLzZGnRQFo9eOdkMkgQRNauZqswIw7l5OUG6RZqQr0ZbwzJKPwlt8CrzAPWj++
cwctx9VYapIoIn+0wB9dCSyd8X4CIY8i8EPWo63nEN0zXOazUNld0QvqhTV3dDa8
tZeC+L+lPnnv1EVD+PY2zHPobQWROTMo9WBcylKZRQ+wk/bMKQuFeEacSf+bt8++
XV5jJuVvmKERuENnnoSYmRY/rjFAq7TPPBs77fiKEREwA6YV9pQjW/VESEu1ys9Q
VVwfaILOhiaXmHyppjJog+k7pVbP5DjMjFCIjC9wyG131puRPJb6loXZsZSQ9ePx
mFybvs0rTAflyenPMPvBKeKf1mYOegA0ltvTwTuoomXW0zHF20Hv+Z6cbn8Jyfqv
VAeNqXHyam+RPBoQM9yhFbGQFOQKcLx20W5bLiv3w/oM4KTSjzNosBeIyZvgx4V/
Fm6nxQFpPoJi5TxS1GsPmt3ftjY//AZmf3grv4smSQZ+a00dtSkqQTabULGvpB5u
TJI8a+z8NogPm7VSlXde1re1/VqKYWxiKVvdiyiDuiniOBbWGXlWZezQMEStbPUJ
U29xoAzy1WosjkShEflvctq47ks2Qt6ZGcyqowOhLmsneYS10ftytdP2raiJKOVr
JyI4lORl1TFggN2OsekYeodBanNS8IRHB7Lcw9IEEczNCpNDdwkLiRNRQvW51v22
fkBGyFng8ZQTX4U2tRt85Tru35xNgMolzYWSvkiN70QWqoXnYi9KPbjxyoQKioIB
yTh49Q37Pwgo2nwimiN24yD7NLT6LeXfARHuEJX8G22DGGQnX3qvCcw/JzvS5xSw
UNsQcMBUg/fIaI39YDRzn6IezhjwFA1gLSNwHHEjitanHbnYBY4Qp9PC8Rs3umXF
MS6QgRNtxs9W1VzziIVnxL906kMbwsXoh/yDskEIYCXCCF4rQvyifczOzV2DwpD9
sN6z1oWYyN5RDcoTX51tnpR5tl99HquNisIUse4RuVoXuIO6FI7Gkv4jTfLSQKH0
muhlMlUM42qvai92P6tl7BALDKvrv60cZtbMn1VZAyL6lLH9JeeaYhoK3CujUIZW
TUU8UXoJCCTX0OSzxzQXnl4oIxF/TLDK3A6tkblCYz43kKvGDkNQ+yUtUXOlpxYM
32MVfzHdvf5oDM5cswsSc+plJe5wLoZ/mRdNn2OLUzU55KxkxEzEv4je6I9/xyBq
MccoA3zWl8QKYIGY9p490Hk9EMHRKPj6gjXW02QQUhxwlHUjYwgZJvk+G08jU8VR
LyxUoC3fWrMLb3HYeXVK2VS9wtyHgCn8jBb/BRYBXc5fUfWiOyTROvGxkXO495d3
Mk8dNVgEbXmq3bDZp7ShJssMJujxVzgb3OuB4TS3IOsJG1CG2AF1Uq/ZdtalG+JR
ICMiXrRqZFi27Wx1CH9MO9DmA0S8rd5UjbN46rfwHj1AkzqbhTJbNP6BcQt2uBU8
R0HM0XxkeqXjHF1cZvrCMIuRB0namtlifZBsLPT1U9OJrWSW0COh4UXIgyjGkRhX
bHweBXlG+QJYlLTfi60kGpSKsZXQOOJgMtHAU+Zxv2yaXpm+AuTEKVeOj50N8rjy
NvzcOPLZ1+tZVOM52wt5Z8urtJCp8QEmJmC8Ujmf96/b/LYYQMyo1d92y5tNyUVK
oWW8oRGdYZw3aFrqN0dPygpkmhU7F+SbJvzfBLYf1GOVvMeoefkpLh0v5xFPMdeC
w8cGn3OXgPKWwCmwO9qiz7a0a0EMGE8UUhhjYSErVbtqSu5wJW8nz5D0v6mZjbeX
aY638AURAzdWzvgfR3VAuA/20VcOTreCCj9JFk7w2ie9YvSVvvhjal5ESxEUyd+9
aHeQgikTR/Oj/0QgUt6EduzOySiRINh1oL6cjXQ4zFIJjnEVFUlCqVqlR7+ujnfy
rs5MbGz8/Elkd/31NKyyyJwcRDnpdHoTV5BvQcO430qN9lmTmYWsm2/mv+wnd6/Q
ejjnsxxRCZGZqbKsKxuJLRsLQeFg1pFu78gxjs/XeGjUlHlKm6e4v/M93R8nAetO
hvJ8/xh6h69XMiwQbh9QJ8L6bTe1CZ2Wn1oDkfhutEbOxdBPMzANty5dFQsdOTjM
UVBrbXR7wGZyjzRQ/xeI+yx1KqiGnWZumOVo7DpkNVOujSrAWPitFUhaBnk0WXDY
HTJnPI5bUMShew3YgGKDT/jw9EqZguxcAqYKo+h7ar1Vymw1aGo+CblBNOz4Lmg/
5ApyuyFLFFEhaXcmwSIQIiUv1eON/lTxSB52i+fjY4dIpZfyjlmO55siB8e9THSn
+DcQQEfHxkOhGsNdGXdq+vrCvd0rcLElDpk9lvg1AvdqvyeHjieIva3wmJ3GnE40
Q6qT9J+y/hEeuz5+hfQJBrKgUelBmowC+hALXQpN2l4+9R5ZRqL3fBeKDzd4KORS
lj9+O9x/LjnUfHKRiSJ2lNpT84vAdEmsTKLAbRWUQr94wZvQmGwOBRYiVjqS0Zbj
2EezO5vhDnYCn+djlE2LtxC+Wvzn6Z94YPhbwLelJUQbEzfvVHWA0JgP8D/kgqAY
cZMhEAkDE/IlhPK0GItGztJwlmvXSXp3P+jl4ZMdB5Inc7jdIr/vRbO53THvJZ4o
/xVx79fP1hYb6ewUVzxHqIUaXtr9KenlDL89uvS/LPqzQbsRITvdOOFJRP1ucvcB
qQwCrVzmq/z+7DWpeU4GHZ7r11upiGn+U1fw85+MC2Apj3qSMhLhjo7ey1wCqiw+
AATnW1vMfG0uvl3fI7izvFnh6o2ElS/mhBd3cAUSsGrRk+pdz4IcOD1L6U/LxORd
amIziv+BdMxAQb3Mbz1BVP1kVtnZSciWNtmKUQoDmRQL1Cca0qv2sm7HlBZwZRwX
oyOvKKtGJ194S6I6upDbiavl0eS403uMgNVLPccmDdFPzwxflUp9LelGV8FJQP3v
Mzy/kMLoC8jTy3oPk/tqJoWUsL2DCXPpgxSNWM6/zug4d4c++N/DQIF53/d2WW/v
4NPd2o4uBInA6mT8ESbz6gsQOKnTNAmu83tIaSBYHTzOgZF2UDrr7TJM/DC1mlS3
0J3LgU4y8nJQ38C5LIJPj+5k55hUlQ1/t9bII8C034T/ME+qFFAJDXs+M8Qd6v0I
opa+qoG1lc1B6L4VYP/Dyj31sXfYci7O/FzYKG/HwKZnCkKuOwWq986nvfBxZ7cs
hXAIZ7lYIHq4bHKMQt5OzA==
`protect END_PROTECTED
