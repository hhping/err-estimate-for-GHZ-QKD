`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
svlHe1ECnyqvkTW/vQ+t5xOzTIwbqODCLBEeBuKeR6Tr7k+xCux4Rz/z+bs0sXkK
gRioubBFprZUACuvPg5APt/uz8ec0ZMpQYsrnQF77osdclRvEt/T58zA9kjMPJQC
oaQa0EPboqX7LaTXj/FcUA0vV+qPt460QQ595yYX7tChfFKrh4Fb23GJYTNUGwqh
PSvaQ87y3udzb1cHnfI4Qnxa4uKbom/LLcdsgr1cnNMQC3fltXGO0gODCpfg+zsq
qC0hLpaGoPFZ7KUeYXNCqxh9Cm6RobLuUx4gYmqK2z4bXBdGAl07FW7LY8aF+3fB
98vW/2yzhFLV8OfjALE+PdstFXZxtDggIor/kE5klktldQ01scyU8aEXBcG+DEnp
yoQDQ3xAyW0pdJowG7yJLdMYxm96ir/WWrDpNkZLuJPLAifb7wl1KeEZiEwRiGS1
1qPiUrvQM82UUDjsEQflzX/8X2eKGZ0X9jXSjgveHTvuBqUkaZjZYgLIeXg9f80T
gtPaEKWP9oY/FMN6cYbARgYa/XO4wmytkRH0aubNNSRXAIzer7o41EXgg0n4BEpN
A4dR+sKgte2n2/laWQba+uQJT3WhXddjvIHKlIet8ruwV0O9jtnjph8xNk73nRRT
EPiQWQiuihM5afFfguW+tCpZrnLu+D0OoSTNWT50d961GrjZfUrznw/PCgzmR6Gc
M/MZ668nWspGcbRH35pf15g3TQKr24HaIEroXdylnZs/x2GOdd/bxFMpulglPMjw
x8YeMSSIPNNGFMxp8ymLtQ==
`protect END_PROTECTED
