`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HsspNbz5Rbrml6fLWqV9gOVE3hWU9Z4h0piRhIVxupJD85eXYRbuWrjo7qGHM4Dc
vrtj6r9XeRFdQa/Z6woi+XB/wA8BJJdoGxjij1Cfnhy0U7XzVk447345LxywjPUs
4TuVj2FFcJhL//Olel0bBI0cpQQDrmia4qTxY5XnsIWNgd5Ii/qyeOC8YTZxEnyZ
0KtEqheYcnjYbqTB6Iseoq3l6xcj0KspvGurrH6OewoRV/+CsgPZEpKtuIe7+RzU
kmNvs5T3lruisnVtXvmCythdu72/ze8qOeW4cVH/SPynMDRgQuYUO+ZcfAFmdn6Y
ZcAEfBJM8chE25lHiWzlqNdBY2hX4icbhRp2Tqp66UudBT7lUctngHyKdcXJg0Wt
XOnkOr1N79p/jOSEp88P7OotCAOxNTWaYVKC+oerWxBMRpsEAfQBvoCEbwVw/zaV
u0sKIrWlTsmq0AiJfU/LZ3aZ+Ews6qQw81tQJobx2VDVXlWLHcfzC/Be4pfjBU1v
b1eY2mnl+r2n3A0btQuaJaggEgiCl/NeY1XADXU2zzCFngkFhMiakZ3cmdEa3AzW
01+soeqQiyVoBicfQiJeQHj1HxWYcXKc2bJ0YgYXy6ExjktQxW14vFF0W8u8Z5qc
MANsoKo3jZX5A5jrvntz6WlA7kEizKhSGbdT8ts2MLlbOUnanF0YH6aUrDbcdfL2
Nqig6tRWHZpxftI8ZXkBZ84AABpkR0Oj+heE2cWP6AWBaTJb53jsEqxIQBeFOeYO
3y8/9QbRVgQhPSrAOM9V2VqYxpUsZDJ6+6T3IBWhsX5rMKq9ytqRB8eY4n7MWdPx
32TNFkgt3ymulO9z5TdMZ5nJ3V4vpXv6w4w7En81U9rK5fnbPhXjpk6k7G3Q2TQF
IQgTbogWK5b2H6M7IctEJTAMUZCmRkN3M+LKi9HS2mwqZZaG/Tc5sQh8tV/hBySb
dXA1DATgBR6zCzjQIIjCYyAjg21vSV9hVn51CJrrexdDulv2uUFnXnfeeoyLxXgU
8NiMpoV8Ztx7xIT2g/ldIblBEFTH8AQUXRAkXlk7pN7Oqvh5D++bsE/IMRYUSZ7l
DkQiuX4uPpLxQumrt46fmYUfyBNWWVYC8idRC/EQtTOh4FJ+MIkTsk4RQ/P4GbRZ
2+8CIHN7PDJP7hD4eAqNxkSvau1ln49nd8uML4XhuAkr/WVzBGpWZyWNWkNPj5eJ
HbVgw1zVnZfKVrTOrATU0Q==
`protect END_PROTECTED
