`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wJNphZiH6HbHUCkksdC94UzahOi1S49aWzp6URHyrQ02YpYZfluZoZ2YcOoSfYd1
uFZUuBYvA7bYEeTjIr/LG+mUPm96z7oaweIegXgrm953XYCNQYC3cg7vmDhFzexm
oz5jahRDecME5tSpMX+eVYBIhzlMmblR1aoqKySNAXoFd7sABf6+nmQSy0Y+/9E6
ypDx6SsXjGR+YKBlrMaiflV6QT/J5hHWn1JjKj9IsY9nzNu3fMskxCMPVTdiEyNo
rWzh6fFLfSRralRyAcLorcs47vWNz9eMuaVg1GyjP4eeC0rxdG66Kc4aQ9P46EK8
Wgb2rwuQfjNAvd/ZcpIcN8EPRZVg49ouXcfS6HHH9aUktSWj5hhE6mK6U0eaahvH
3UydzyrbhsZOFUoiFE2S6eTm69msWCPrRlfYWtx8aYCmmNzPjmLwjEjTS5bBMwp2
0qQIUOKJAdYQdpiLlB7kUzWOlXKJzkE6bRFBEqi043Pa6TtLzlJVEL7OzVCsYkqb
vf0O3+hhwSmz8yRILQ59IWN9Ki1902w64InM1CULdvjoM9Ihl93ge/czuTWsKIEa
eUNVILrrHoc5UpL8u/RBiezsa1A311mMAz/M1FtqIhtEhOOLDDaHMQkoMF/owsXi
D+Ao29erIyxpD1byU1z1Gai54Czga/jfqd+7ywfwVSsfjkFo1SPsyb8nQQJspBYg
jkEKw74KtzqQWxB+uOI6eEOWbQwklDK5DcPMNwQ35bo2Eyu/DlIyJ2PTGLucsV/+
l8hsEPWXPSfkJHF7YXUdUdNEf5IZoTSqbMIa5OBPZrze+fUVjRMPwFZi9hBOtDng
1OezrG04UT81pRfTHc+Ky6tKyyvhbfEsbwFZNbYGeplLWRv7yQJxOhmPLhS5AtGN
eLKZgsctPI/qjP5je7xULRk2aW/Q/VXi3FqBeIE/M10=
`protect END_PROTECTED
