`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6pc4yCsps4F6zfQAUcYq3x+GiqathtXpalDbiQeyYEget3DVsf1bsgnFuLSllr/3
w+H5Zw2RNc/bV7TrrdTcdGR66NU+Djqo5Pz8lQ4qaO+LFlPwLaHjqMjUchG57QJp
vG+OZGSYepJdLH/1qzF8d6/Y6xJwq7JXHJ21XAWoECUjTEBmO7MMASff7grj/ysk
FIkLwkjdfwxZS29Mr/07QOB4mctRWzLuPUcbU76t5WoRXZLVWiXTZ+BXbqE7pJTE
VQboAaHtVcVmvepQ9X4+ADy/eJORJVF5XGfCidfvIDAkjDbkqCN156z+MDUxGDvM
P+UAk10epARcHG494t91T8EuGkxdROxZb/aPImKh/2G8V32V5x67ezN9Y/RYTtIm
Cd1kezSqhMymWJAzm5+M0u7YopNPZIHmC6KvTdXQ/fYdpVTTg7qBp4GpabulkVAl
oog2wKIum+cWnRW6cONmIoHaCI5zqVpvGEHKpdY+3EGsaUpYI5tAz2Uk7mJgtt9P
2QmiI+SgQNvVvhkoTBk7u5jiWPcTiKJpaCQV6UA9oBya1E3cqt63uBbTJq/6PbyE
otyG1X51spwtkB9hiLimYt3G5yxwf/6be9aIPowNYCo1hGBw1wnOiAZ7drY/Erts
wCSedGio3mQwPlQ7Ui068RRIkA2qsyDVXxNd6yipqroD9mU/gD3T2XNRGdpvTnTM
b83AAzEs0MjnI45aF3BqmEcQyUgQBRIQUbx6I2Z+jdQo7vOOORRsb+zPYVqeWsvn
ieQAGo8lWpFvd2IGsfQx2cu7BsiKdH62lmZ4Y3ll5x14bLzheAthMN2pGdKxh4I3
bmskWp8V69sL6taWHCqWMBW2bbfUWzMIe3XQ0JD2Jsn5ObJqTYAslq81RXeIA2F/
gL256yHC3WFZbMkoPxRfN7Wwgefjrxe1d2ezSSq7hGbzc/Z061GXvviowDvs+IVH
WY48MmchVBwaJ+xc2zlYyILaAVT2yLsbW9EIagE39sXGhkWrE5Z55kWe6HSHEHG1
ok9XfEtcHUxbhxOQcbqYLTgaEH3Q9J2JSlUr7wbCH8c5H+4CvtODLuoj11vJnTg3
SPyuImawxrzTSmQp/Vw2Y5EGA9c1x5eyaPNhrGxcvJ3+Ib+HUsUrwUitCpQFDRd4
3UbDjoDt9fZOln56LvKHoX0cuLKSPECmhC6Wo8GCw7YiIN3GDv7nRV4eCsCsUAnw
cx8kiCmE+/bkjPir256ZIZJXLzj68lp4Ubo93CNqLvC8pZ6DgpMbk0WGhLVpx8FP
Ht1TNaktVe2mhvCxzmiNv3ZUaEtBAv8LQnMs3e7+PXg4k4r6yqygB4dhHT/mKCvc
vgdRj2pzz6OMF0zjc4sO7qj+8fOhaU0kJPaYVEdSQxwR6hx5nuuRspSQPRH5Bjgw
d89F4Ml5HUy4cftDe95hM6leyyGv5yJzIx6+aum4lvM6VBD97HYP1bNF//9vFeYU
RWZBvu14vl8t0DKWYMbWGkhGuPy98DC6bQiLWgBODyO7pu2oozPA9vPcsvefwu/g
QN6f6qR6zkA3GMGAQ5mv21xbJj24suya1FeAVmj0mI5IpqoCP8sSu3czKmnodJj6
OOcajmr7lFKoXG/8+uDtBUEVgjfl6qZ3DjE8chccBQEsw1LLOWd80RHH9czUECm7
CBzrZv7XGdEp6u6cYPZMNhYBOJN+ZRFvp6jqno8+1jsDbj0f+4gGUk56h6fT15lG
nt3t42H23a20F3Qsv/mlCKso+5WM/o27qGW/kFr3TXujl3/tCLLOyGMoDc/D6SBs
sflKLdbrFNiO5zonkF39UQ0cOwBhuVZcaBSLphCBkkL3TUvDyCYqom9vkJRfV+5O
0r7ludkRJdnU6jw6k0dE6rLBUsF5ZqNNv5cNO6+CX9m0XxIzSmJ1XJ5gVFhxwAGd
h7XSdnseM7o+OHXjkM9Zhokay3ucCHq056F2hi2vt1FAXA4kGWfgOJOSNTw6lTKC
HPHYkSNcSFZsxya5ycQv9Mv0IkuF45QTkjtsbAgKyVgyhG9vMJ2a2q0I5e0hARiP
tbF0ytpGLOXXfQYoVF8/CAPeoIzM0CteX/Ig9L8mX3l2flPqJamuKOn2K3RtYBbY
OOQ8txEMeq51owXzZtoBcuuQ1q4c9vY3Vgv49CEfaQn9lXkyoTKbuIaVK3gDwLZN
rcHemtyvO+kVGYgsAQhhLf/t15jfaBg5hPjVq4lt26uK64EjYCod8VhWmXTF8zeK
SyTa5ALr9IERFU6Z5dd6OLlK0xjHC/Auh2KDWft4oiPosoOlhnFZBEBvB0PDNTQ4
`protect END_PROTECTED
