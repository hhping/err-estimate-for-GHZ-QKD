`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NMC7EIZpjrxsx4HOqNzSONW1H8zji2hmUyxtqX0wf4axjPQ8hVVHVF6WkTnSbwkv
0cQpqI43RD/7QlAUAS9nHO+3DlwtVBwW3mnAStEdfp9qo08uxIfW+mGdqLr+VBQH
UgwuRdMKJrItlmRBF2DcRS13ClPt+UIzFG1HSr2f7jzoxkWyL0OinI/EF016rq2q
B43GPEpfsXuI4aSbjdCjiLRMy3mx707xraxziBjmzBDKajoFe18XWHiRa9wb4D+M
+Z81VJoNhM+K5XqL97yidy6x6pcWhnxkwPZQFmoqbqKLyNjkZycV61H7MA8GfTjq
AxIxUjalO4JNNxAvJD0MmTOLXVUUkWYX+aBN9Sc0FadNz/OwPGTYbPDB8Re/qFtk
hJgkXLjHIwQLzaBh/Jmmd90526eiExmOXTI9bm32vEb8Dl5/qKgI9C30Dei1E1ZQ
c/y/U9ZbLSq5d85+SZrfYtUtNXWONySfp0zngpPkZCVOndp9d0goJ80Nu3cf62pC
iSRcRGFx8Cn08I3xkBIGL3eDljBKdBnjh7V+H1+3kyA9zi80VeO0/YwN+EKf4uoH
XDLT1KSC/ZrRFiv30wPOvJ/9CUhFM5CwAj6FBhPUbTOBG8SSBl1gassUl8G64bWY
owxo2e5HEn4A1JB4e2S+w9npROclCkRpDKHBQo/f0v+uS3Tr8sXLOhhomNfr+JNf
A1VK8448F9m4a4AFO7AiufAl+KI4VelTLSMxf2i7GsZysE0RIOw3b+4dIsiWmQNM
YUaVoAKIq4KHURjWYgETvTnkxHk5JwaYjUmvbFBnit0Mv+2bpxA+3eUjA1HZRj6W
dORSFpb7/gkzS5FNgFvqr1rxMioc1EIbFAr4w4WimNuUPmyfEeeZV8skMTwAkA39
8zhAQpMNmgoMrFIYg9GBxOHkcgGRnpUCZqNo8aT2ZXbg93m+Kvz6CImmtudh+U1N
TskYWLb84+Qnqz3hiqK+KtQrHnnrTpAATNZlfrNiWLfd3HK0KtNGf9hb5iD/GI79
OyNhX25AlDt3KVs3zu11eQ0AwQJ07cmWW7tHPeflEEoM+ZxX+G/5aSafH1gIoe6X
VYzJeKHLGMhzW61QGe3s8MpDSWmXlb30mOgpd1TVr01dmMFlwyBWfwncWd4V+LQT
/JtYDZDltDHbVI+1BM4fzj7WLWx04XvTrN/4+XSYjTPZ0sQz44s91/K3eAmu/sEn
diXumbDIyZ85gNgGw+qKSw95IpbgystWEN/g20JlDPcBBTPGuh/TAkjMaPlOY5Fn
rMTUmpfFDraYhzTJoEdEXNSRcdMvfX4Iuz7OWpjWh4xZdE2S0b6NtocM1UJQG20V
6kr1O5Jta4OXNtKUnTtEgC4ql1PYV/ysfNalbL/W43Qt4Gxf0RX9Nr6dQJA69FC6
RIBfMcijucFc8aUCwExYW2BApX+7YEXLwcud9lCl514uRHOxr1faOHAeuKO8Zxql
`protect END_PROTECTED
