`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z+AMseJ7zIK7wG3EtkXTLFJ0KYKvx2u86Rnk2Iq2BvG1OtqSRElwUxFdHvmbjAPZ
+Upwgq83/E//AqCilqOMIZos6QTvv8S9k9qgFBlGGB2QodD5HsdCMs7bbbSmFB28
bWDvEkw9h8eaakR3Q8LiQ3UWQTlXYzaIbGU5Sbf+jNNJoJdgpiMo4jeTe3mx9CSj
mpZU9XLY1AAHjLXfZcqRXZ0O6XhiQP7HtF4fgNDkuUujqRTYWTkojSI6J9HFRVDu
kUPdyYidLfobX72jk71YluYomt0YKvxgNS3ZfWM+rL+4hFfeS8xtSb5/Xk27L1ag
qx/Ur1Kde08rM/Q3S4G4uQyUbKqZnETPt1LVRPHdAaVPeengC6+tVisOCtmvYtLC
FnsbFlzvsHsXt0EtqxRkDIVgICYJ5/Ey70jES7jsUQ+ocxC4GC/QB75m0c9CNzXk
iHUikp7Yjng8dPEAXDYRHBeqXjzn6PF8GDc0s6y9VgZ2SlRdYgezK7BZcwGCKW3m
uUbOtsA99WQH5EtQLQKXp78rOeIwFm+Zmp/IKP3tqL9ZwYtub0ehidYLxMdKH8Zg
0Amc/C6ijJYaOwyPlw0eM4HMw/WM2cY6ih57Fy6NVGLbkPJa643OOaMY0AiTCIoo
kVogVAMNioqbqLjse2TJF848cGXXq7ZBM6FVWg/yfe+gPc3JRqyN7qSEbfn9FBrg
HiY1j1pBLtmEmaqhGoLRoY03AEgg5O65eG0E3vdflC1KQqLIa7ydhEwD2/k9K2Gs
kAj2VA9dCb/ZWzhIPVitNL5b5q8NJwVwABqP9eIXgcrXqErle+UeWHhY7QUHYkpR
OAVl95R5KsMl7ipCLcuUlAriiMPrTTUJ+Kk3qg60ifzkW4N+P46RZBpBaZ5NnCkD
PZ5o9tSa/fIXlUGAyRdHa+cDqCT7IyTuCOo0uS5STQOQ8Ip9ETCuQnYS9A4YLm2S
Nv2pimU5rfYFXu1cvRhB9alwIlS02eSXnklgpK4E8SqsC7t2ST5FToMN4GFLfcBZ
ngDKuzcwNSMu4lt1zsLMPEsEgXpnI/QIOaQSW/eJRXt6nrKI3qZWaN5SnTlcvJHJ
FosPWCyXOVXYVfixVjHQoLwnD9bKZRnmzfwbxp3hGhIvUOPEirTr0bn1Sc316y8B
kpS/Vf53JxjJp0lnBTO5jSP6ajBVF2Uj6oGIBv8CCkd+ApgczEoL9zpZFBf3wOZN
1djCvsPyrdaDRMULw54uo+5Y28A7U49mFZ6I00JZqATcuzhJJlNi3+a8QmEfMW1a
XN0oQKbJaKjVilmQFDTTMBqtLMMJGtNLOR26mMr5L+8RjnPQm4wnxsKloVWtpujp
2tUGWxeKnYIBc7wWkaytis0a43l4VUdoVpTTO7CQZpm/ZWGS30trZfp/iMLDQunh
Ya87iudBK//DJj0FD9yoQ7SoU/nd+rEdJhKJ0SF8dAYmKvBfvhsqbL9uht6D4Ujq
Wx2NJx4R9BCj3rX8NeFx4lZpR0U8+3wjbbsCZGcuda/pYYpczlZzSuwJxr/DswCQ
OfiHN/z/49n3Xx2vuzpVTScSG3t9yBTMCAGBLbO5RFH/HGa9WaTpmxfvlysLNNzi
9aniDAigMGvviUBoRnLqECa72TZVxJt0X1MwX/3vPAlSNALo+PS5aiEkc83O6RTq
Fiuzmf1XZu4321fQAoTv0CwDOwxw4YdUoaCGdTv6LogRHSYMXH3xa80VAXg1LHsa
tQ/oJLMuICsyFfG6EWuACjCZhFjTOn3YMBpyJ0ZStCAqWovg0nzJfbriSq1eF3JD
BmVn+8UJq8N+WkLdomsHnAIYJFLWnA26UqsVt8D/ZzVi8ThSsIvnvXXCJ7y0YGUp
q3l2Dm/nQv5K8lPXZruY3nGrW5ypBTErOBdI/aOb0N0RG8qQf6TfmMGc32I4UyLp
fcJDRjibmkyhyt1cmGF6CAae6A+x8MVXkF0X5cKvHDBHMf18Z+f3EhNadJFAre3M
0Q/hOdqJ+bg/k9eKrnEpnrAJtbkMbk2955JlBzT5WUAhn4X1tPqe6FtmqujIOpk9
kMySdiCU+X5BoqmjmySUlYhWVfN0zJIvJy9ZHfFJC3BlxR38Ynjw3I+rxnQP+vvH
fFc08tD1nfruK19hxAjwFO2Ph+NPhKm5jMCtM+IsHIuJPCC2cW4D351nV4luzl6Z
FHw7QW5L+9s+R15sXz7Lcf7iQkS6kMlDYmyVX5xw4muO3gWIlf4dJrrapSMgEctj
UBIL0ZU8VWgf9jFVtpeyYtZzm/+b3KTsEl1jTJXvivfH/8UjYEMJbgIeaG0hB6Ws
jVy1h7KcRX+GzmWH/MMI938mDQoe+Ze1+NWVd9Mo0Yo=
`protect END_PROTECTED
