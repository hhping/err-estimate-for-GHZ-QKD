`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XmKkecYUPx7wY4K1FEiPOub3t2Ovd0E2+Fso3EScplrdWt30/wWOkDSZR7e2xQpV
qCYsJi9dGS9s/D/TUs5ofuarEv028gSJnfVUfYTtwL/ZM9rbIpM0Soj7Etnfjjoj
dAeuei37jv0vh6y0dPxngI2x0zBQO3Sdc0pnOJrNl8kJFE2fDdulfOG6wfUwVKIf
dF5nZKMUo+IyJotqba3EYustiGni2Zb/Sepqezf2ljJUdV/hG34byPWR4d0h+rbg
3c12mAhsNQWplPscD2kJVeI/WuLxzXOGUL4Wr+syiP2fA3FYFehp7iXbiJ2YPETs
/EgqAppOVNG5y532pjb5NUh2V3g0wAdC1mMg0Efs6HjXbP3n2oO5DGUDxSshMQ9a
OXhqmgOeSZ85lBXQH07o59i7+zghqKRVeoKsfWn0Gewb3Ab+6dt7vdXjP+oz1v5U
herF6bhytxu+6x3w6k0AxCkfxjaMqMnFx6gKxLKIoLVZvF+YIzn8j4jwbQibhcqM
JulL9Li0wm9jactdFHe9WbATm3lFLm04mvzdaWan2gFb8XzuIt79J58g7KkHkt9q
Qc4MzzXEjI8dfwrgo2rjS9Osfqv5/2TQFzpLiCREUAeUjk3zicIqu2XJcyYyDOPd
QQU+WFI65pZxAhzf406Jp26rGD61P1de8a2XDckYsZVA1NkeW73kS3HyWMg9NxcC
vVr5FfygJDvGgLpvR8smiAIDwcJeXpZsImjBEsNjW+kwrxh/x91nyWGqfivCNkL9
h4svbHilm7ZEbuSb3fexakQPQeZXGdAFjO1W9g4SbdN3SyQ3MNpgdSGAdYVS5Hyc
`protect END_PROTECTED
