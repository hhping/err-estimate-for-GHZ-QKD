`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IBLlhLMKST/dTxyaH9UkEq8zmMTLonMr3cFZmxS3xwWMdFwp6OXyxHHjdzDHcakx
J1f1RPkOPjrq16mYtNL5jEdXHUXLqAVgStOB1DMs30/f4UV5mu2kVZ8d5A0MeH6d
QOxrAKh6AV48Ww815J7ajVDyi0CM9Md0K4hZjuZ3IoKnoaN+tG1TYZbq1tGRjsf9
aVZ491nwhWlufLvIMVoHimPwlNtMqSI5YkrqDnzRB4SoQDU4hT3iTLHkPLFqMQB0
D8nxzalfr3xfEmzqfIRxVYd8iwymIn3z3DzmUDCribFb7JMMP54cghUZsCN1lE6b
QuMFkw71h9bkXMUlb9M8DhMLdbXJm6OEavaNcJnkg3H+igLa3QTKuRerv/e6ft8m
uR0Yw5bRTyNz6f4tYq2np++th5Jv1Km5ayKRTBJRlfrXMEwuvCuuZzT3y2Y8tsrG
MxDkYupjl4JglI4wB45XLugOQdsqLur5xgDltZBswcTb4/gEhYiUDmn8tvOOIeUd
gPVGtTNFRLkXf9DQKYduvtUBe+o80tBjYOANYq3v4JRo3MxUUA6O1HrDIa0hYMHX
lKBpHW9ymr1o4mnsyXd+EA8qNk/3RjBmITMkVFoPYpNem3j/vgHrt3smmfPnpm17
Mf3LiRGBk/PrH+x+bImBt6fV4/J63AcGI/0B790+KhxMQKsmWPGP/vW6Mki+QEIU
`protect END_PROTECTED
