`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v7wgV/WwQWn27FgzRonD/BPlUxGeRnnzj9mWTb9QDymiTSeLqryHd8zI2qzRfthg
tsjKtCo++zzTVVpO4BK5ghEJzA9kLu1iNPA6pImqnYdatASBSRE/xxQDIHvotxRL
iJ8KK89/0tCpN5sch3XaEilctBVefm45b+tVGPwNeycKvPjnKBiHz7w589zq2hW1
QGnuMYOVTzxZftH+doUXz+amqTJ1ff3Im0Nfaikyr7Vg7ssOQ8SKCPyDcCye7c01
TRGESqTzdxEbxfWa0HtR2YQ9dGOrn3TTLhO9v/i9vVuriA578EWrldx+TzQyAzve
S7/aUm8lPn8LkL7KNMtxMS5NBoYNxBrzDr393nPgmElEjfU5sOxLSZHFt28uT8LF
aI888B3cslD+PRS1Xxb3n/7S569VyxJXqHXyHkJdbU7hHaozIEFjP8Vgqwdqndj4
z3GjwJz21BFlsH/72mcIpZre4+HrQkkDuXdgo68bj9ziV1oEs5d1+1Po2oFxovbo
Ay5drGXoKsMtHn9x5BAKTPcJSEVmijvoRiK1anJ3dJ8sw5pF431YrgC0mNXArw4n
jW1lTRVtI0tQ8kX64KoS1vdMZ9cHa1R9gFlt43nSM0Yr5YLpJcWCYLZv5btxAqam
0gwxaHWt2gKnZ/l5kh1y7970rjkBG8Vxbh7nYzp6782LiYAXpoij2WH9EXduvQr9
IPyEVyPnsqWSeAR7qSHBv8ZMIjfA4DjSfzhPITkd6MkIo9ebkLJF9rlSkYZYRBea
Olh8uAn6j6nQoy3RRJRwGpwMyzSaYCJKLrCGJNkdvTOz2cQHbWBD1dEuKiXynuZV
aLbmPSW620fBv3Z34/oCKBg8x6f/pZ76nUHicNQ1C/M=
`protect END_PROTECTED
