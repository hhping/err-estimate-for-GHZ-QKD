`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dn1Qxb7HjLLAwElr7AUa0yxb6s7xLOi1tNrv31tIzwjngPShxSavdT2yG1rAqz8u
hjZbBBvyN+b4DXGfT4pRZ2n4c6JMNyeoUS8mHW3H72MwpE2y0IfJapRyZk6MMloE
bAGHJRkAiW5ocQPDp7C3XVqRyw+HB8APve84+Ed/4Q30A/T3GcOJWwshvPOGnAYZ
Pd7H6TuKpIjYH7RtemsmTkEXEyMLhr5p42YiLqUlzNcfSCzVlJ6QUkFS30WwAawF
u0PsESeAX4o3Gkq2oJbwSxL+qKixGvbYr7nvOcsfMWpkszz3+ssJDO5bjbNJ60tI
guxpBQ8GmiZ95E3IrSHrrrqdpFEs8BTpPE5Dcv8u7krMxjEHCq0RBU1TwuGO6jgI
Jza4g3MzcGpoaQ8H0iNsz10P0R1eGJLopzesTDjkHn3uqIgOxeqyJqpwydgMt8Ud
N32zXeuBUzZ9yJ82flFS3+UxnPUqmgDf5OXESaFn1oTgO54Nn5nf80aQfxvfBYVH
JwQL2TkGhySk3PZSOmN4zTnjAuhQDH1muVjb3S+kjSZAOxmlZFOmKpbKddcknpuJ
PDUElbtaXm+/sPdYxeLdO8vbijZWzfr42qXbZ+B+lC96+lZVKvlavxkT1vhGskQn
kmBDIRe3owGo8vkk93y49yzyQtu1+qYUQJWKtQS8W6K3gnri+hEl7zyQODQitMOg
lNeATyfghOqacBJysP6sRbKq+c+vlIBgE7TRfn1gk2b842mIwakiow4nnqiP1rP6
n2zE4rsiCdcgLtnxGAUsQDiSTt8/idS8W2qa5RnDxIHi6eLissV1BxO2LmRNCj/S
HIIoZDLr7RusHrRQYAAujeFMW5IfvZX9r9kafvo4nGTC7r2Lv4XLISBQqnfUubBL
UVisaf+jgDibUi/8WCaAUeENAHC9APzxL+IZ3ZFqAfVD9W8g71GYBaxyP6t7KmHE
chtCgbxurmqpJFBSeAdw4BG+XUPIPfdNvw0GGRKUHX5PAyMQAtqk+03DbhcD7moP
sPKLGPAOp9BEQ2VXqx4I6NryfjHj/YAUyghmGTekU6SoUl92RHVVpVvL+EqvNPT4
YorfgV7sgXnVjYw4Dyu+RpR1N/HQpfVWQ+2kEj5CChifSDi4ajI5wRqEYf9lg8m3
DONl+MWQruOK0AEtMiJHdA8lTKtuV47WkJAIYKxAvh1n/SlILGOSA992hULvUBi7
HCqwTdFgjmryvLNSPsUXA8irYGyjm5gFvWFSjGtuCxyag44w+AOUVO60cqzFY4TM
TQ/eoK9G0I0SE/bwz+maiolQcuP0Jofbubg2AM8Ht08=
`protect END_PROTECTED
