`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SMl5g4T/S4wJ/v/Yfh7tjnEDHTFmc6Ex25r5bSWWdPs+qV5X50eY8ehC8Gg8EOwh
DLwa7+Qr2Qps+LWLjN1r2vpfnC401AtCqHlJ6nirmA0RvxHp4WDUDXH1GMLcCUG/
1gydfnA+KGG7eAX/9MUwu60cBy55JAipdhntoom08V9Kxn2Hmg8SpmLoAYUEOf67
/lQGBhYHjaRSu88ad4HqbCCmJ4XFz7OwyQrY9k0IWB3hzE8OzOxM3Zke1E+dhwqi
Of2mzJPCxwLacnQldvc4iOAuziZZprOCa5i2TYAEbBvdt1GNM0ZxoF1iZSZuWHKn
OLhy+WZNAAaivTBrDz50D7nuL87KaCC5wZTASfSSmUWWl99rorvoEmuszXQHVuOo
jLES/XM/hp93ufpp19+nPKT6SJByklyXh0t7faC96FGNo5/EAv5R8C/9cuILeNc/
ro86VW+9UFuqEKrsB0iR1+rhkVOOBfXJDK94+zC5MLqDjYPo4RMdtsDtOkjgmKrh
qNZ4Kz22C8JDOGm84giEEcI/408WLdVs6upqVVZpxTZ8Vin0BX21UDxIjlXYvwGX
wk2FjSlf8lMyVW0ZlJsivw2gvggawKNCu0aijVHsmNNpzs8pQ3/vo/suKezhN+yV
QOJtVZCtAlKLx+onUtf2v8otccE38uhXXLv5Gx+ena0Qs7eXSiy4hgS14f8WTRWK
bYxYJlttI0fvKousuDcuj1T16peD6u0W1jv+VoPI/HKP1AzHSo+mxMBgZCDVHgIX
P6A7IWDt+kXYiSj8/aBFsGDgV3PuqCvAfTJT+DEfyThu8X9XPDZvT9Wsop1uQB0H
+T7uGuQUS8dcZYfVkjMQuUS65zGilSJYlvl7C+0nAD5C4r69VWYDn+CSbYx3baUJ
VrmeM2l/8PP5bLUkRW3h58k+UtAfb+vMwRYuuzGiX6SlZZF9UDYqu0Mf3XroNK5F
`protect END_PROTECTED
