`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hvS5viYvnF5CDjvD0JceIpQ9F6ZjhoO35cmFqEM60+zyfhWCIuzfJcOqaKdbSV1D
BT6iFyPaYFsxdg/OZ0lKqgRZk0yZCwef3drSa8Oif4cFZxUyBb7GOtCB4AbnWFzo
Pk1Lkc5L3E8gEcTqIpnc9D7IJYio5XBsRXtH9KNuXnLDNWSLVu7zmZj8LhpGP1mS
f4vNwbAP8cYy5qF699Lw1Jb14vcumZQJ5r3/VqEj9Fu3rEyNx07hO2Q4xkrwHZq6
vYp27bwelfxdmJofBdEkOvTi+2H07fowj06tHUkC3HijKwbWzPbZLKSS4A44SbgG
FO/Xp/imLOcwgd7n5Na6zpz4A6wK7LGg2FV49DlPPCVENGbKY0j/QrNMWWre7qnW
vrSmzN/qj93PJGEZ2UT6GjV3mEI2/gZwAKF7ndRWo6SgNfMZcjKSUALdgZGUBDq5
dQSUzLvslyLeUXvvD94iFI6TwZ9ZXZxVLEZhF2skaMg2DzHebLIWl4Fx5opnyx5Z
sHIJiRDeE6Ddp8Y1bfPpbd8Gta8MoIfJvEioQNwnSTUq9HB/2mAm7kc66jn4EbHj
pVQBqTpSc2VEcnXxHoTCp9hqeHfaK+VC12FwjbyT3muB6Kf5ve/B/qRfTDYQzLTt
VySTmWEvX+gIsxIUrJe/bqwRdJs8Y95f33dNlKKes3hdYQXeXRKMEl5GWNDNQjer
8gEqs+PI7g4a6kI2CKsVbF34H9vXkRchMUejo1erDUBBIi+PfDPKG+Kqh8YlO2Um
LD4Nj6e82wSGW3dM8q3qxrH/rzYNWhsUlJpLBdLDkeOki5TOisYPfphVSp1PBEKE
9PBhSlnWPy0JbHivn6nccgugSbtqn787vgHwinR1aa8+OWpHw5xui121kjhISHNR
Y7kQ5dqmqEEufAA8zdqt6xTyeGrveMy6ECcAfwMrvz9IfuS8tUS9HT0lj/GIPn8F
Y4zhllySDFivzBoYXqqbrAid3RPvrRXsl4h1FeJQOsrAzSzJpRFFe/8Jzhziier2
OHndSxJWn9rqRlqRp37JNaya3jb6Qt5t2WwWHIsdq0Ex0zzAtCxAnPaa9S7cIile
EkR3BWUIdTbageV4ce1SdvK6BKCLgpKQL+d5lXsUDl1S5POk/zzG4xMZ0P01W6ig
Kj0xwFg/YBeixI1vofizZC0gg97hBpqYLcf25o3oxrQ6CnWOBQlQke5Nk3kVm1SW
VnKIEfIR1uuvJXOsdDmuKLz6FxSJQ/TExB3/i+3AlrNQmL57x2JsdvMjqomcG3fI
iUD4573rA/9sOdXk4GLeREMC5EEmagbepwRTsqeHJWe9nk6FLFM5C7IUnPFz7Tgu
m+Zd7LsoKrEdsB0ugg1/ZxIRcut7NSsubDMdG4n7Sbi3TE0iO9tOvQe0j4LDjGgx
WPPA/ioe00MbSlCiIpGVAAmr9CHQhjt65sQsiNgOZn14ka/1QzcCcyKrES3l1ugv
MHaxDk4MiFCBZ4W0DuM2pg==
`protect END_PROTECTED
