`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BWjlXocmtXww8Gpp30d12ofKJsTl2rQ23+KOP6gCnJvnvRb1H491ren0Pym3psie
RRxyKkLRovWhyRayjKJttdKXawetcs+sxY11+iLpwSGCmks71JVLvzK0oiLURQ9g
3eo77fmRQ01aNWAho1iKrynKzrAZvVFB+4EsPiRRes2bmg1lzv51cel4IzteIo4V
QDBdKKW3K9dzdYF21Tu9I7+Cm4OQDZTJwj8lD5dONfeLIOR+EqyGtld70it216fw
Dfn3wyYOHz/KKT+Zbylosu+FxMWombzGqtZ/mZLxAcFsGUZBI4sb1LopFKMxyUZp
Uvq/5G+iBtzlgRj0dCwmc7zmXr0SXP3aRrCytSrpAHJVjuxPwmw2rlQD1JlnyhoV
aXYEIqkKIQx6OL5WWMDczuFzVewwgI9QyjY4X60npvLo1tdrs89pBD/TtOri5C3T
jT03AnacNP6PHFkSBFTqXq92vOQgX2tuQ7us3E58pg01MDKc2J8FXzxYXSX5qGx5
6k4AjWwG9lOhylML6NeOSrNHYywpY0/UzyYI5zpy2Gr0so3mysbeipe32GaMPbZn
kNLypoBQvSBp3ru0OfsUblkspes4x/Z+eJ97NHCyI+KU4tlcEEYA1WRLxQeJAN1n
ZXguIVkXKgA2tnFBwG/uiqr6Cg3gLbpS+AETEW1dZcn+m83E37xA8Is9IoM2QOcQ
YYBuUVlNAjhkK9g9gLAChEyO/44L3IVAKM9HdyJc51ojBfL23rKiJcfdnm7HGrbZ
3HxtqhfNipcSbnwD0AfYakKdj8QBpFpp0JfU29sY4KEG0Klv14a86udyamsk9PVG
ouFX3GBHAiTu8imws9bgtZywFc4IGv3fTzOmE+mZNP4yBbe7yh/bKb/gZOcYaPeg
o/NXhPPVoVjpAIkbaFvocl8xtF6MTFrPbItF6xOW4pHHVwkYh5Ya2KsZFgM0ivQy
0xrP5r11yZnJauQLkiGlBTNaJjSG0KNCrm3kmNlLB1VrYpmI5Zal/HWIYh9PQlIg
T/uiUW0o0l/nVYx0mDcJNK92NfD1UdSYXokjM6z8BTIkPUvYPUmvjrvBSxuGxzmg
rS8gHQhGRs/fYswBiu0G3XaviBO91VS7ErA6mgO8/Dwqld2ntdq/zUhFT+CIZl67
dfbaFL9DvKFnrx1eWPsUBa+GZW3+3MriHWZJW3WS+EouotcjfIklVnECG6SLP77s
dUDClyMPgztDphZls5LP25g0zYmmjcHTYXRgK9h59ePTe6xrMKVdvB8gl0UUvpR1
3JgEeMZNFu082ut3WF6U0qm99kUBij9gOFHtQWom+b8okmXDFrE9XgOYWQESLxt5
zc/DALmsaYq7tHt2kovdyrdLDY2tHfXoyni0CHfIQXURoTzZVbmX2OX+fzKQEUTw
NXRmJ0NdDiavZ2UjaYbr8LVGhHZGQN6XNYQ6NFkWlZSrMlD0sPJvAZXc5SEQqBZE
sYjPpn0xJk2dhEWQz6xMtITGVtbUsfcRRrFKomR08s6Bu9sp2Gjwoj2ZZ0JbYYPh
jx3O8oLyIp6TKvUMoC0gTpREEFfnRKPWx3fhgcTrDVjOUodNKHFnNxtYVXPlfi4o
cqafHxHty8CXTR6sxF6cyu5QK/skffHD8b2AvYqBR7V0fxuwwzeG1Ewj0gnb8MOK
l5WwTb6BNq4VaoBh+h8mzL/MEk+or/z0/CVmNxdoAQVmnu3ZPsupEkU9YvEJ16TP
TmwSf0yFHYbfJSQL5DQSTXkvD/7m/CBYzTPf9Rd3CSptONDPz1SFhHO1BtevK14+
6HmQTZxilsEx0TF/DiWarpjejKWEZhhr5JQWe1pC/GFCPFlRztBEp8lbaUbjoOSo
Wn5zQPVBqcJXXR/3bjSRwJsiL6p3qvyl/PgFp7UhQdhhInkJrQ2zhgcrhwnUz1l1
YhVTaNTzeof3fCukKDL9+rN+jbvYe7jGIDYG9dFsEjjDbfJ4BRJe0je+vSJpLRpI
JjsMzTEMJ2+jiNOaxKlNN5CksgwYTgziaMj8FXROjBQv7v7kT5eRYbRA2sxaWpXo
9ZKcWnDt9zyROqswnR6vxxiXy9XCCfdIegsc+mU4TgrbUNYumL0cIH//hBqQW/Jp
cha3JunN/egl0XQcjvcGa4bZSWpYsSP2f6biKGPZnfDY1hVRImxK6Go59nIlsON4
n0jDlTlPTP6/S1xBWsWPi2k4Fw/ZHHOEwFNy9YNjxCgpOCH+jMtvF2fdGlWDr0zI
Y82zw1dHWso9cRqxchyRIpGhV8nMjA/v28Y6ZLLnoUjz9tHRGAbKc+kwZ9j5205x
ORPenlu+OGu3L/ywJ0363wsIsrAQvmbP4Q9qZpJ9oReNTvGmvtgU25b5E/54sZ01
8FzA/4/XiHtB8g5gXlZGuZj224Jc6MhFbJ8Z9/fOKGV0f5mVyZpzLxSKZjJ3/aBB
LZhfnZdD4MTFdQjxgZyVJgJiZQeTIRKkVeRZzUy4A0bIDWG92DXMZzPMYhzli4va
PghMASUEErTMwL8ruI0zOVHKpHj7LOQ3x03ZExEkRNhjrc+F5te5uaALU7qhb6F4
qM7KH5iqJ8o+NwIBXr25str1D5vIM81uodKTel4e8OyX0FIj4SlRxhMuiudE2qhl
n9FsSylHki62sn+9mbX0KO2tOKeYX9OwUwYEIJeNynuJR/OE9n6WSDVCwzDkY9Y4
FUYGn5kz+tdVHhroaf2RVe69pgyAkZ7uPDWr3DjL8s6pgNQ4gaTCiIdj9WeXh/Gq
yC2DetOYzEmTOWiL4N3n0LsKMc0utrA7E4o3qRWr7sFjj7lu3vc3Qdb1FpSlrPJw
sdnsYEcmzq6GmqEuOg6LqxILq8ckJYoAvsUaeq1kJEUAqikQfzSQVr/fgFDnTlRg
hh9GO19vxyPN/knw668Jmu7C9pTQJfyBEiwSBjDeIy24Jv3n7g7BiMCN+8nq75Fe
cF5o7jecAk0e6IsbtaBRqfahN7QI7kAVtb/C46LqWJk=
`protect END_PROTECTED
