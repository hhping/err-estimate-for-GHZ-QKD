`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xmF8H21rShSbTZU9kcE46b0j8HQSZeZfLfOxSo7Ldc3hDQLSymzpTYCAuod7R33x
FiP+Ap/Ygfwxvv3BWQTAcDqeRyzMKFerHCj3ZPv7Cs7YP8bv8heHokrAPH4hTHci
vdGh+aCZaBkscLMmObY7LPgTO0lbW6QBQ3nnSLIhJGdSLwQvBzL+bFuxRcaBXxY5
KPQJMfDCTuOly8FKFpdnrYMiF4YYSDg7onOPbzPZJIIdc7sRjnrRM2W9h+HnGi8n
lCUB7UI+OpbE9FAyavXe7EnCeWT/mFFu0+GJJ1D1bXksEDrSIqPtziZ8EHCXtSb0
FeY/Oow/JFtQ6ufBwnUY4je9HUL/3kDK1PveH0o/ySZitTEXq4x+bfAj6FslWp+/
NL38A1vjnLndNYo4FBGYGcRgMs3Uck6e/0U9PRnKoMjk3rsZsKyPyWN6QrwuFdBt
j5pG+8fo1lxcy/UpfoyHJhqdUS1hAIAti+QXAgG6vdhrmFD3o6W8UaN72WvrcjZ/
8Hupg9LEk9Ma9eLygb0MZx2iMcuQXdrmP+MaZf4Us6b0ZlnmRoHQrbiP92vqxfqN
//9mT/nSxBwtG1rnvCYCwiTaqmV590K+utqg872WK0qxdA8yDeW1ifHwzsT5xlcj
wptcn7UTkn4h6E1B+aebgCpak5H4Ai1ypsfVaqpIihD4wkHOGSRJBJck981rmkqz
2Sy/vWBN7oiX3lDwkGDaJ6M84+iFArEK/XGxfGQBrIGjWGVCd7Umo4TFVNhc5T0p
Zo0Lv8T2algIOa39Sle/v6lTMiNu4t2+6HEiwrndSY3c4v+9/hH1ku9fqVG0/5ZU
Z5AdSluMGg1QFlipFu73pm27LJPxuyVQhUJ3PBPJEc52tCzg65euVXuFr+KrB5Yv
adAXPjCIRNyxTu6wCGxwQmAbVfdvNxmFz/tHG1Ji3o/CrAW+/zw+h7G0SJK4yqbt
9Sj22SjkrPdGV3y3tipneY4CawxKuP//CU4ecSHf2sren6Eqv/tfe7NFA1Fdbfvn
4LftmDsYvY2oi+5z2sdEGuxzXlGW1oiV2CgtL1FbTu9mFZrql6TRMlU80NrkY/J3
UfuhpLZXeFy5+jyxoFMn7L7zUJfd/L8npDCUV2m+70EEij+NNwT6BRK3zNZnPPN2
E5JQMxSM0FMC46TO4l7M2J9wt4WwuvQhB6qT/1JQdpRyh6ih6p+0SQ0WSm/R62H/
loll2M2zdw5Lgcwkf9s4MnljAs0oQ4d2nLZL2QUPUu2U3iHpgecimnDMH1z1x/YG
MHWmBKZm/fVVyIM5kbXsl/hTlp3ZW0QrZDXuoPcG+7SJSGlViaLx+b2xJrMfwiz6
fAlevWZ6Nuevfy4sIyZWA16y/w8nZQQYWqRx463dL6yQ7dkZkZikgdjHDVM1nKMX
4pJZBdlZlosI1dzcNEF+L5BTFiqd08we50WHekc72pfkIiic7yESsfEoUUc3F9cn
o0DUGaOliQROGNj73cpnR1sBWNVr1JCkRUCXeRdgQjsHcL8VLAky0mxdlLGGRJSr
MVnpfC5AEknilqgSPyd+wspYpu6bUOklCOzOg/nakwB5wx76MpcBv1PNix/4y4Rc
Now2xwZBV89Y02034H6EOlzF9wDQjC/Ft3Z49XJd1GzHjfs/Yu2h6Vy2koQE0JA8
6kOtAPUhi8R99dIkUvHpyurLetfbdHy1vnCPmcI6NSdb+IiqylqmGGfN1YqWuyV7
90m3Pm/CB485/FFgueR39ISyO+3XGGrUYDt2GojL2IvcINeqR84nvY/bVYyEls17
2l3DnCcwkTxAO9Xv+rJYNUlxiUX/uW07oM57WUMfe7YXoHhvZGMXwHUQ09citKg9
5mZZh1lLcitXtTx7eIsV2yNQX6STKCM6T3I8Mg+1pNs=
`protect END_PROTECTED
