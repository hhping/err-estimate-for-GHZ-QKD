`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a5ogGtChnxsIy1HPus3EXEnJami9lxVMP8hU0ztKe0JE2cUmrv74aKwgxGTxuQjj
/dxXkG2ECUw16g4AhnKBmDkN3F4PUaYWboZOrAHpvl98yMamXTuBjv1Of+x2tIOf
yFKq2PfLK+fGIdRNxe8MrxH6a00QtKHJiG7qaEBDO9sx8Bclf/WBEWmB/DaE36Uc
xV2OgPbJc+Y7jgVL9lm5hqyB023wubPXAaGuviKlEJTWZlFuEn0tEbi6yGsUR1DG
akuGK5Hpqy5Icjqq7L9Wvyo7eQGEuf69W7LDxLhfI8NnXM4m44biO0adaxQTcRo+
Zjq4pLJLXFyj+eqkWAOINQS2IAFCDazWPCrQHii3YDibVp1sRytEFVVDFy9aOApu
b6pLyJ5zWJNI15OJ/C3ErXYIHlcGgUmwG1FJaRH322W2dSci0TpN1ulz3TeRz+44
H56Zk11jvWXDd+4C9sp9EA6NfzbhMgphZ15EzTElO23Yu1Q6laJQibbsqv7KvsxL
SU0DIenJdpn7nQVBwcIbCgT8hWcMFkGYVKY8lKab4NhbE3bCjM6P9OyRFeWEta7v
SXEhmxFRl/lCICBwO6eovelVXtmYa1UT4JV5+cAn20OiBVs8Ye9okkQQJ1OA43o/
80t371w519GmNO7OwwXRzdgTcMVqEFEXdt80CvefbjURBL2EvJ2OrKFj1MgRv3pK
VomyRqZf4lQ0dXnckr/pY1WSY+c3KfSuNpXDiztQl1hK2BzsU7TzUcBWYlXLpeoO
I2ZxBvixolTebWwA8GXN/UbIGBRHoBwi2gGrM6/yyda0idoHC7rqwnCxIpOSRsM2
0zUuouNQEHx6aMbOiqHaYJ6E8Y1rpI89XOk3/HK70TouvJCEx//ELXWlBmZ0tT5a
IFDeMgrHChc8VgK1SUCIJgYSYjL1/72ZGN6Qst0SWQ1bne1e/uDrTsZH2Mutwj5v
r87N8A25QeVCP4O98bOc2R4zVzvS5I3sGj99DmO3OKq29XQ66wtvimXRvQl+7iak
kCgj2MSnrpKFGosM5wOE+1DpcyY/VB11x8TTHipYpBo3JjGY1CdI7PeCYKK4nMVZ
lcHbov334mbsVHhwjyJYPnC6IAI6906a5bPrBXACCx2+1IkwV+VpUtN4lumUK4ZI
cgXOFSetm/TJrn8P/PkO0KeER2V22xBGXXN0d9uGBvwYPy9ShexYzmZHvlLdiyHX
BjHUrF8kjFPZpUesj5oG+nnvJcL7wL8kfIBRZ6PNRb6Z8CY/07whfXBfd6vVu0Bt
12uOV4I7WJesyMbokhHt0zZgO+NipMQ/wm7rZ7hubZ4T1SSpw+g/rOfQ7zu9lGTC
ivLijUd0vUbWWwZ35zreoSFX7qL+AA1t9HY3DlxE/299+5zTsyi8o6lOebVEg5Eo
X/i9LDw4/yXcWO2S9n2BUppck2XtEZN4E7KM48jklBHspA7SB+zqlwJlvaE0QNuv
qYjSGUs5PSMSIXjkbaKiRl7k4ZzLP882OVa+UhRXydSJ2XjVJhfmAKJODboIqFxC
6jj+Wk3r2CfL3P2q9ioR+M5R7x4h7J9Oaz9bv4ohYInhMXx89hVwG9zJoXVKqnAB
KDQmpgz3JYte5bsW7qY9AE91B+LOK8w/p/lp++rk+dTDX9EnS3VQpq3r/DJ12wBT
tG9KTjSrGlSQtuxb4vg3lylJqAI8WmybUhZl6bybwU4/UwtABb9u9rHxlqQfoBMA
EaoXy1psCquUXl7mSLLNPrPwIl4rQDFypiZ0Hb/ucY+4rJ5PBCCmQt8N9GO4m8YX
dqOIe4mQox/iMT6LunooiDuOpYYezEyv63ZzW7CyqLBU/WVKIsZ5mTpM/l/yFjp9
5gZc2M7oWZBTeLFr6wFdLGCVvKTGToaXjK0FG8u4futqxKQBaJrfz18PN9Rdz1m/
s7hDV5nOykqBcu2ovS7wr7y4HfEB9kXJJfFfvpBECwS+P3FyK6e6GqX5afsFbdGx
CDe3Ox5FbCvr+Xcl0DrllMaOQE70IutS1hcUxjyK8Pt4IPHMUcr5519HCMfl5Kqg
n4N69IsVcnI/cG5NfNBPRoNnTWwN383sJk68SqAuij/OdU22cTPEG6thEeXO/7Tr
rHR9VmI9Ny2NRvUEeg62LrOuCAuPD9OeoxbkpBMI5Eswownm46DYNlTiwXBpVb1a
KKYRFo1y07fonxOd9TD90jl8LWBrSn5KVB3/rSfPmj+GYf+XFd9XlMwo2Jn94zI/
yyaPfDRzdjuTHS61EhQYrirzvjOAdl9OpvUsugrtmCL47CurH3wQ5iRZO2Mxa5oT
Yle9aBkkxjRiWkyprkFKHZmIRCHUZaPOnSU5jbOpjnYWF6cCaCGSVGeTQhKRoKhz
RH7lK5NSkHDozi+ZJVa6ShdiQkb54vAzSUqSfstzETf7lU+Qv5o01JOzCArAMLb9
e3qxwX4iS9Fyp2V3rBL5qTUPpbieAhussk1nUKFAna6+Uft65jf2Isg2d+si05bs
uEt1cggyX0jENIbYX2ugX+eWEaxjTXeEvOH2H4GOXqw=
`protect END_PROTECTED
