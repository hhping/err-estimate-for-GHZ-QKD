`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GhFoYIPqMXOqyLa6jEredfGtb17lZoqkCgrQKd6nDZVEImrQGpj2HHI3lpbi2JQj
PxBuvSoBgRqkvrO6F03WPAFibwHNfLRWRRiT4JTto4geZ5QCp9zaFcvgADHlnQOU
hgVBoR/HrTPqLLc7U8xO6NJ+bMVdY5NJQQp169tTsXedAl3WshRsL20SbY6bGS+j
wwhrBh6XtGg0kkHjMe2RIhAWv/zM56YjcNbYsUu1bscxw33iqytbIDERiInkXYBe
Q2E+yuXjXy9qX7NOPacEgq49Vp7iW0Rs/I9vZkdRF8rc5gGuPdw2nokKe6Z2okiC
LTAAI4eOJAmq9KxWPxk+eAkZJJeB87STmHA5K+BiOiDKfVy0LNslXnxWxjy/6Pqn
QX8IYvY7TbhGloK7D/5QeNIdjZ+7UASk03GncfTd0qQquG+h031To7xIoIjfJuNn
j/10EliVqXnXkT/ozw8SsvKsZHKt2s8oeTXGNEvI8SPpwhiauCrZp7f5J/4665jY
8bW0Nie8i8hK4haSpiBUqhntb+lxHyRbdRSKQTGo1PuzFQWEx8CoJhONClHiQi5q
bXZJRC5plmIqpTCFTp15aeUwhHPBgvLf0b/aNxRhGu8E8n6YMFh3QizX9HH7tD0o
R1zGPTUeXY8OqQQWDBQZvmXL0uppXg3DOpODko+z409v2LEg7Hn5F569FPhV5uH7
IVXLvQwDtA500RSl8Vi6ICVjACW2xc+hFNfjhhJqzuHsLUBlE2XFQj2cCloA1+ac
rJ5pmYY8XL8qPyexYHsNxA==
`protect END_PROTECTED
