`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6a2uiBxor4cbFCzfEbB7QjCUrJ/1vfBh9vUccB5rQGJbb2PazuR+3GGUG+qZjh6A
LQqiPXwDCBGjySMkMfroq0iKa8z4v/9QOABY7X1zyKVobSe6jhAPjr/wqy1XIp5D
kLMptbpC1Ig7bzkcp8hPW9hTYJPsKZfGvbmTUncmtv9iYUznyzxqsII9O+9LxDsz
YE/eDlmAaEyGdJWycf5NC8riCNNUoJQfImnc5371NpZNUPaRJSzUazPwo48ulKND
J5uaTASj/dH9975R1Tb30EG05okRm+uQ+AQqrj6Ys21/69/FqfpKEBQPRxj5UuXE
yQbuYttnZLGQoqr5TnE8kvLayyR0q/Wf/5k84XBn8CYdGTapJupcfs2RCjLWRISE
uZggNCawVsqY5UqYfeKHaD/pif1zxAQpMaYDh23N+gIApEBtwcO6RS1tIEVbTmVa
04Hb5nOgNCItE4UZ9EFj09rs+3dSbVAc6/pc5UYAeyuJcc5I92Anl7u+X1W46KCh
p7UQwLpH+eMjq2FVfVauUgwZYIU0GfOtD1HlWouEQ0cS2SRHefgRExVWYhvgmtyr
8F/Cv3rdkUNn0DPWLOe99+wUz4v6hiaEeMpE2/7+49XeEg0fxZSImM4Y/Gim0c6z
atNle6ufJqLus0ZaTuZ/cQ==
`protect END_PROTECTED
