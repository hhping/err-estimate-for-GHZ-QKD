`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mvnimEAF5bAo2gK4tlFj5+DxK0GPurDjpq1PV12He5htS1zVv64XjL7vuZw5HYGe
kL2nlvmaWFiLnA4CbqkoMce2MZW58C7KE+cthe1UwFYTHSjZkAEmlLPxpoBN5+X0
35JVeM5J6BCkjD2lmmY8WjLkHn69gCsqmPbdPNkHyOW2AJcsoPQ0jFIQVPAvcQr8
emj1Qocp2Wv8h9LoapdDR1Jm2FqAGbcZioWaogTj4W4knocFFTrkU2JMoC4sA2bv
to935/wfO5179QGk4AJgkDsJPVliKsrlRrRJPePOv1abkHXaCfk/k3ZDxNYe8j+o
8KULz6sWAc4tNB0arKlVPYX1Cjjc39MwBx5IS4g7S3eJXXSxOlshmnnHfXcBjik1
gsI1p3977MarJtYauWZFImn6Hek0UQHRomRvGhZ+Vp4dee2Fqfbkdkqg8wgryROK
9BokUtg6/L7ZMGYfbtrg8Y2lGNJpoZeRpUQaDtjEjHPXYEzjX2ipJg9KimXFFuyc
yrXvNnhpxnUumigGzg+xOOcxoFGkmHIEkzFV6t5Uso/rgNE4oamjWzs3zWrCejOv
tGIQTggqEwaEFhPvxGW+IbPXIKUfiNOLQpuCkLxaRqhuu9p6iG2IFVhqqBC6KYUU
abWvoXqB40nTKQKh0M018g78qxEbDACuDCxgmvdjdzupEWAuOUcHxsi9ImqmvBgF
Oq3LK8eA1yPDZjxjlZLqJFMTkOlaP2nBk4ds/wBZaEiUNgL/GdlDz74nVVKn5bs4
cYyPHFUEPhZOxnXyFcap1nwoM+/bN/N1Mm8qtWroMJmFyFqm/e4K9rGf6TkxlmkE
TKF/E0xLZjnRe4jqz2GNhkEKF9Gp3J1lVqLSlKU4Z/KnbKEeaBhwSQh8GTVrjJuJ
wFhKXt6dKdDw5TDoM+iUjBtct2WxajYzs39988nKLuGlPgIDHJsOA+cxUTnkQoaJ
t/MklfUODbYqfNwchFDMZ5jbFZCONcyi5kPJLZyO66ARtE4ZNgszfPBhGELTZ7xJ
c57ZQjtzKqGJDtoKpf3GTd2X5HJV0q3J1ryU3wEaChdCoPcXgwoEst1xItChFbme
1kj59TBExwz9Qq82GKgYvLeV3WY4tHUN/a2jLZuz+Zzrrjj/yziNpzNNErzqZeRY
XdDjoXiJ/0mylwps1/SxVt1biQ3iVYnaePUVknSIelCYJsXT2/Dx7YcauQH2O65t
du7N+wJg4HPDWFvY2suh26uSUxfbtMV3zIu2TTYsg4X784NCuzvNRO1Ura3nbUhM
D7no7245JWNEYdCGApGq/Losopaez8Grf8Yxth6lT4TAhsHz/BmZKmUeuBWBjeEs
79Oc3LI7R/NpmnBES9YaHtndBinIXQC5bd9LZMDl0bKOWwjc6OBeN8J5d8vl9PHx
dr7sM6Pk3lFSgoB54dV9AtNxscXrsn7ULMrMetu3E/WfrqNxCZsSbCQ2M55QXGnT
LhaQ/PRC+rBRizlIdmPqsBNPmMSpDFUG+QCYT2QJtM8JD6Z1iPA5SfleeGUoY3e5
Sfs1pGhU2FZUn+W2sz724EnyIC0kQreDICCX79s73mWg+AuU/4rytnNYxXPZLHVY
jtkiPDeu8XInjE/3inSiEIWGgo7FkHW35axz9KxJYpK7bGjW7RawFktD96qEJbMI
zirUncK5nBRFPSP+sm8hn1qlSb+AV7JBcNx1RBW7rnY2osnO4HDvEwlfLZE1cpRa
`protect END_PROTECTED
