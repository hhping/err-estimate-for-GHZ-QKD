`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
keST85J2fFYGOWdYqLLMSAs3ENpi9RmLCDhYY0UCByg1mco0cw+yl4izdXxCZozp
34qdni9A1KvL5GA4pf7N/EgfruSw9yWpbyFNw4A4wvbrLUv9TAlsqkx0ojcWBufz
VzJgkzHKIvmmQmfyc2yPTjgBEwvOxpVw070P6RRctH/G27Gz8IL8zMvRpqDpT1ue
IVILeL1xDXPJggmeNZCANxxfL8VFjXU3c+nzihYv51VPK2AncZBoVFfd4yY+Tvvh
tJIWNQPOHCpqfL5bRmDpQBEWsVOWi9J7NMw9n/fSGpsWgoKtJzBBik23sxzbYpoN
q5Mz+uWEVdO2v9hauN5WOVQVdVctxI8WjgNqycvzBV8l9SJhzwwMfp2V6APsa7tE
SED313NYueoMz2tGPZAagNETC4aBroOWoFN5J+eP+/2/Igsil7NQ08p+7YN9Y9uR
Y6hv9P1YgjQSOAT5kgTcUDRwapAIMa1DPMunnEGyHS55JrJC+FdfsHdLNdHabdAt
W2CFJQ+lKaelwWWNToE6iMpbgeouWJk1A+chKX5l2ERYQGofOXsWMcp2duC7Tlq8
yvlDyumcicyAZiWr9ZQIC+1YHcR7f97UWPu7vLOBayMti6zldnGo3qPW+05d6OU1
PL1qfNbOYJpW30YqEYge083G/dMz7/cY1CoQx0qiaonimS7JmLmSN/f03aFDP2YQ
QmnCsiF3JYKiquP5YwtxKUuAaK8t/rsbarbCQv33jAuJA++bcBdkedIdAKzpnwP3
`protect END_PROTECTED
