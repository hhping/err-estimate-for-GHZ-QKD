`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oVsVFOCb9m1lnEaURA0PchlK/SN/XpjRzqlM8KUE2nY/pHzK0KBUCMBiK9+DRcZF
Di8Rxdsd+PRIeG9Ebf5OsIknfC6cls0v+TjkUGxmESa+E/tgdXl8ZFNs2SE29nYP
IPQMTcBX6I7JD1GfVJCi0rPEew5PY0dz5+rvYo8OAyDDjg8icG+oBQNbv3SVgoer
KH0pxftJYWuBaAAqXC/Psrf81RBrVeOF/EkQpEkwf/0RMBhHEbbalMk7uOXBblhG
uxK1Va3t2ikuazAtU3NSX04o9zX6+XYGzKbAcqR9DEVunB7306auLYS76xup4TLU
j7f34C5n0erNt8mku0RCWhc0Dio0yjN840J87yWCNd7DL8iDcjElxjPtcL89mnGZ
fZFU/F0X9e2F1plOZgPIt1rRGONg5s29ckwZSei5TSoaWs5duTamPlBCDxmRnPlQ
b+iVeQi8ZjB2Sgf1rQPqvnvATshOkGAN1F6penRXpzRtWM1KYN8Fgbuj2lbiGwC2
SFHqUrksfXK8ZIPxHUccPP9r01QsI/N4kuacyFh8Znq1RJSy0jXt0mxaFdRXZm9x
Ptvd71Lcxk8xBFE70FlqJVUCEZQiwhBQdNfk2/N+Wk8txPHJCG/S8mR/K1hg01qj
tBuJ/bpo18h2/7saX7LNNcnBlWZBzTUUXtImJQ4XaGpKcu7+jNWdwfPM/hVyR7Wa
`protect END_PROTECTED
