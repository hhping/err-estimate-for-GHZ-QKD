`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dx62xRQ6+Y5KEoeehfNA0HGldSfivcxOVeqd/u2mU8d+XMHFATZGI/JI4fGgD6Y7
xetzMcW0DSulk15Vz+tK+E0uQBoprjuHeHfH6FGWI+ZqSFChnryFRIUin7mem1mB
mTTZy+Cag6g2Vww8dzIPE7m60tBRMYn8nnu9XHPspBtMxtNwy6j+yKmGVGhD4i1M
hdD88FP6Cytfb1YqmZp16JWMo5LYanDqM4yRb2J3+EXqnM+Q4Pb90uejlVzCUCb7
3OaW1YEQjEvDxq6zQol4DQdl0wo981S4iH2+Uty75v3adqtq2RaWS5ICt3wGNtkx
R7wUMernKC1FKAHsR9hkd5izTqGl2s23tuGU64yMihSCkhE4pQWM4xgO7lopJc+W
4P2mHfomrGdLp96KiZDzLbd7dqlkprUWkpQgE7yRb5kKIlBX77MEFWtgBYuNp/GY
7xlDnZnENqJI7/u8o6e0Zw65W07u34Fj8/ssBi3hx/I=
`protect END_PROTECTED
