`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nM/F0Q96VDF9j9dxcfFwO1ZPmjAR0bqUNfulLiJ4HMbr88AjZDjP1LWGScyaqtr3
Z2ebKkfr6pqIpO+DHRKmxSae6QIWlROCtenX0cjs9G2jc2q8dG7C0Hmps3iNPSS2
+v79XQsbLEpvMeq5i9BelUrGzBzHO5cFLeKooWSA9tlBZl7dFupJVmp06CqwOaKr
mkwoz4rx/t2h++/dwtFYjzGbodxElfIbgzoYfrgTSd2Kc52Qb1Dk+x3zpJTR03t+
q0BPyOCoCCDWXMI9Iv99l82pOJ0DnvqSzsfDfLj7uadNH+IQG/8mR7vRwDcMnjab
u152qV+AlDZ489rL10ABwEJWDzvYsq/+pRTE1pDl0e1X15YVOD7mxN61VA0ZfiME
CFaZuCVxSyEF2qsBHowpOvLtgyh/yR0/DANwAJAwQTomC5R3u9OlioVq1wk8NoAR
WavhiAbgW6Vlq4TbCDDm8GM4VIkPac/u8ChegN58+xb7mEikDAvorOb9J1y/F/10
A9sZA7FNABlKJKWPhKdO/aVNMMrmLRRlYDCw+RJvSAoqveeAb34hFbh6MvK02giV
u6dk+2vEKgZ+eArkzkPnEwNjWE15zOIuLAQVQmcVe8cPNLTYGDKayu6SYX72GQJd
1f1e/dx17IBA1+spn2aZZSZFuV3+3JmddxiC3hfpqZeANqWBdKBg7ihR8/CdnafS
HEKZAxMZYFwwm2ardyPwa6Nkz0YiQAC0cXwaX1wUQIDQIUVpUFhwsJtPKyJz0i6j
pGRAayHPxRpYsLmm6yStRKzs2on0cTxQnb/Z1aV1tCRe4lZDAurGReWvgJpVv+7d
3x6rMDpCo0HJsSSSFpcCfzg3AGMIFqLkVeamEGEsn/EtEEtG/WE6WyDxG+SOqElL
7UILqy5d52NK57SsSDgPpyT+gWmVeArNePJQHLiP27WYZjvJL8velz8KHSCeH0rK
8h2SDl5wvTstOWV167VR2+zj7aNzVYB1qtT9bOO9ZDSDw4lQ0xDPInuoix0nmMT7
LblUgR/SgkLpyAc4AbEa0wkVh4eGMwzCcGkoNhZTO8yE/aXd/w+8zJSXeFooo2bo
WmQE+d+lLbIabRXx3VV1pWi1GuNHfaWYa5BzII6WZNt/zhMA9HN4I5haZu5NJ3oD
6A2RkjXKid8vP6XN28Izs/fGlKHqgc8FDz9ETVlWtZoN7Dyco/6bZ/33B2XJNTMb
o+or8EERNtN0aDP/ICXKnCyfkXst+g8vmKqQoAoABKAFC6nZlLfXmUq9IqjFyupL
KxI/qT5hMpLxaqKD7Ukvpt8MpFlggFQny2OMNhRfSkEuWSxLaipfLc0D2EHpwrfc
UuXqARiHMirCx3J5+KKix+NQFdHDpCKzPZMWK6Qwe4Sd+SwIwjk/ckSq9iCTzlsM
23inhg1UqwlBAYF8aGxFTJoxKX/v90lN2HPAfFK0scVS8FJnwrpjYs1dY4cmq3XE
Zzzqcxd9o6cGYwZ2VPgCGM6IX9Vvrzr4nBozSi2AutWEIWfb0uJL3JiUgmXUckTX
ZPvjLSzuWdXEGLfr1tIxK9IzmH7EySRo0t10zEbJIs89rDxIUpoNHB+8JwKF3Seo
ivQv5cDdNiUkPrGARig8rOKsZHECHqD4L4KIOcXYbwQcP9dgeC2skSr4qWiPBJAu
T3waqa3oSFzkOAqXPMZAbW7MkxNd0JMBJzZu6pXxa+oSdnf7VekcNjCxWtyYDrim
B34ewfnMndMTDaSl8QPc948rII0GeMH+nSKXRxyIckOQfC/3rFaqhRnwz7dGMtFp
ObfEyBXIurFC1givLI6KC6ue9+UaWr/4PV8NRE8MxCW3RFQlZ5HlphCW9vuEzcBW
FP3Vs2Q00/L2M/bDYttoztb6t/EQt9IdfpsDGtGIN40H6+vGvEHzLJfFHJrDxcnA
sdVrhkQRy2Aa5iKA0efBayodWbqPvFVDGsYpkBjidiVxwAdePunRrV5vfmfG+iW+
HFag28rug/+ah2LGTIr99A3WGuumpmQNP08Qr8RZRYaZ0wnMsE+cDdpXUoIM9Fxu
3nKZ71p1iot233SuWvEc6xvSt/Sa0TCCLA+6xohboGNJV1jbU0CdbtnuJ2I4XHGK
q5O6WWrMEoeEYfl5AWa5f6ULtjyOTwmHb/8qYxN5ql/conV8k2UsGgquh5XGn1FC
lqFMsl8vXvSL3SUR12SaNCvbfGrlBb9l166FU3GWwFWatH/+RGUJIJfergNOmzom
px4KDFNFlg292EeS15PJJhgFq89Rh9w6+iW6iqxXlaLr1c3orRZHFKCuEYjK6j04
olbZf8UksENbHa2XNQ6prOq1u7+lVk43YjUSIW/iaCD7qIepsJDP2S+JktDOwSXg
DEWVBd/qM6wTPuLvkzeITcrGpy1GB9Q88DDv2Z2AiVgSn8VlcJ6+z9tflw+efz9g
SgOGJQBc7LDAj0doldZ7WlD+yHWECERdjmzo8+xpg+tbX4AwhnVfaQ1KCu1kGy1l
NyvBwTTnWWMSEWh2F633iFWr38UNO0ELrAqd+1RQe0JzZ/tlxhmF1gTi5NK83jJV
Bm3PVsjAVXXEP7Ey0yPu92IrFZNS+EhO7sMUseN37ggVgFr342OABbyZtkog3xRv
JK7DD/V6uLxF5RDyoXxKjCILtZYjsa+sFOrOMNnp8VvGrVjbxuk1Gqa62ebCwcu8
OmRW3MKbxaLoGC0gKHtd7qCI/UxaMl6shPDsRJQEmvokyF/pYioFkrTQnRlv0Ofy
Kjcjrp/PtbsttqyaX4pGYF1lq3iH3KfDwI1GibGPqc9lI0YGCyd3nnDbCSRxbNyF
AdwLBUPF3ycvt5HromkOVJ+nTzcLjvYZAG/BuY/gdPO+hk4NbPDqIEp5mfqrfMO4
L8iDJisWBdsH29Cp0wdXEO08HZYhPAF9MHXO6T2KDrJBBEIFO8+kWb+Dg7xNHAPO
odsqMHF5EykgphetwoE9mH2mhJ7NRbtFVSpiTujR3p8cjal86T2aOlaTEVbFTTLQ
qlTRTece5G+pTIOdgjqU5zmeYVbAqXJetLPyKgl7hT6HlPzp2Xo20pDnLjmue6bA
G8/QBFn6pKNs98P3Dlh/An7CixN0E1CELsu3kwqFL9YHrlqsucnlTtMpgAfNwDRE
4h9ddlNrwH1mYBRP3rB80HmK38gbuMSkTk9VqBttXtBFKiHuL1G+eWpAh2jkyrSe
K7T9V5LIQMztbqaKjKpCezFaalJdHrgoZqDbJN32txl/AAlLMEE/XpxKSndpJHeB
dod9SitPQr65S1Grph+L90fwZGMyb88CNXoeKRG1/ylTggwAyQ31+Dbp7vUDB127
jQV3QYnxLYMUGkxEjwX1JpJQjwzhKJiepxJURHseV6l7l3JmFxYkYPMCuP+zit9z
gxzyHIjYzUi3OrRjaZjPi1DMf0ejGSpQD+alG/GFWBhb/yCXEcz3FMcX6zQp5s+i
9RVlUTilNYYzcaByPkqAKq62T8zvSNBESN6cjvzWQz9TpS4/3CAfQJjJQqSWfX5k
VcZu0X8TZZPCmizVaVfCRUVQvFK6gYYqthMzl/OcL9c7TqPKdp+DVKzj+5DW+xtW
6BeW9ZwoXjzmVBesQt6B5DPaQjJGxSFuyT6xXdUVKebbHrzJCEE12AoIQx7fn3FL
8sTJCFq15U0Kk/weq3jBCHF+Z1siTMBD4iohj8EmEKZnF+Nziq3xRO/9be1bWzu8
HWKZm8RBvDd5opY2FIA8LXmRN5u7QMzpQY++7k1YLdyRF/B6HabLbHR8NXq5DYlI
zLnZt6nGeT3Lsv6lk7XRE+IjhRqqy22rlLWMcS5fRzz0yEvrmKnJTAnlH98ZQIUa
51gm8CA5yeazmkBXdhzra1i4MpTxifkxSvt/EfgqRbf+8otZZsy3hHDRToB8Q/Yg
Ugc7uQNCADSj7B5OOyAR0z7B/mJnbYjSMIL+q87Qh4d5TzdvhmJpnfDbWLjDKOL4
Q50edsSCsFI2IXlOTRP2GncRBUF8znkfNr8+20ElMKExuadSfTLJzHX2UjaopElb
gKsxNQUqK1sAh/BCFzIISItsLT8GwkrI3XR2f30BZbLV7zGBZFxK5cJqv4kDP9vs
xGeb1Yzk9jREg3XOGjOTx21GYYQapcqBi1RDbXjNxt2uSCATLoLmHMGeEv3OuJkj
uLNaO9GCidtEuF82jGVt2+HzWePR6fOnOIHaZvQZ8elHMGTmajUFNsmllf97rIhL
`protect END_PROTECTED
