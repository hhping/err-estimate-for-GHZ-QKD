`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
99WnFNahHOmqmG0HQ0xw07Otk/zR7B9Ma7/KHiJSWTW/TIAtLDiWmJIAqNYPunBc
isPY7iLglwT+VpC6gnO1xEogKf2uwW/1hKBlRCEAVFmWmsiYtDcQ/puE75J4Jl7A
av5MvuP+Za3NEJzO9bfeCgInvhaIhsEpoe6boHYLNsZdiTY/Qv9x1LhwLGgRQN4N
pw+CzjXj8XlNJMXg247NPOceGQJZ+sfRm6CGOuvT6jr73lJIszk80bVYanR1vaSt
TCUBzhoOxOvy2MBAPi2a4jzzwITOblRXdX8bxh0eYEAzalCsvaGzaAFv2i06ChLG
1kVYbtbBLJ2LHlM0SdkEToWmVKitggfkwUOhwpoAUN4xrOeWp2XtEdn4zqNFymTL
TzrCv/0pyje/o+UPRnFfV4FYEOioMCvKy0G+f4HE6CYBiFWkEVOwSTitceEk8gvT
eKnnDM/9AETOjRNVJ+Sgf58llAbCiSSSqqEzJ5LhBwEFLo8BRyU110eqpwy68wJL
vP3VlLyoSPMfuz2pjkeOOSBA/qxWqquJu4WDeRfSkNH4MR0filIF5q4M26jDzymm
gT2g+fglcJTk7BD1DlZPuCBM0U369IRjS0NkyRMcCtIPGn8OzTiCVeAPKbuMLSJr
EXVdi1ZS21u2idePuvXpqluCTFSX1525tQ15Pwk+zsXKEYJC74ZT67aoMwk+fhwf
ZOJtbCuJnfbmd2BmK5Nbttwoq5g9zskSAsibkgfnTOPTdYxDeCw6WMk9JLGwJvSt
zIEC22spV/BmvyC5mo0q+uPTcj5zrtnjkZeTeWImOWo=
`protect END_PROTECTED
