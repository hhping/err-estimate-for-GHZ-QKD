`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JjhMZQo0sexxpi9XAtTiNsllaln5X1f801y6DT7swPQqvhBQPNTzjfmeBlXXEQFw
JVvvQmrp1guUdiX3QY/Dwf/IJAAaX/9EABe1G7jIYZ05HbtTJrfkQz4d+dpNW622
pLfNcxEN9WEmSpdYnIrEeTRMkyMrW61K6hncyy4ndDNlfugXyz4PgxNB5W8U+MyJ
nrZPKjF2CdcNS/HtbXdeUs1m8I5FXqqAO6pWd4aBPi7ZrcFXDq/i0GtXxbwvMaQF
5rQSc6IybSW0MmtjeT+Y7jH9TZSP6qSOnsd9OPYxN6NVqL1nClnjXSe1cFfTo+cQ
naQirBhqNyMmDX2AQYkJMdU2hP8UjXnso57EHJPKEvAZnHMiAujfX18fQ/yDzbtR
UR2G/GN0rY+RoWA0+4sF+w13fY9rJ6eFJ4bqdmvzFwPMpeyPt5sj+c8k1+PGejsP
F6mKrcmdvtn5ytDaiJtpeDNv99suhHNScXAb+53cKiZPKBLMmGroL07gGhXaaKSa
MRoVbW8SllcbHY/0Hu0D6zw+bH3npDiaRBCXx34MO6cbBmoWh6qwz7zx0E2lDGlz
KfCbKQ4AnFcjlH4AWuU9067dbgQTa1xHxFo0EooKHUXbzJiIgOyBiRzrzeHcC2Ml
Yk9SS4XGDybN0M3VgMBDlFVK2Qal6znyn4BhFAZRnJWP2aSFX8liDxuDM93muDwv
LKaMMGYuycmoRzKtqMyYQw19Ce4Fwe50X7mGf2E023GzzuLXq1Tb7ObYWKqZGyZe
jlASdzsvzuDOyKiR+0jhhvHxIb9Xd2y2IFPZZ7NbhiN1sPsWpBJavwi3ZlEP6KGR
igsNOkenObHnc5RJgDYtXq7KhUM0oJ8GImSLhr2wLJKydQcfLuLXCgAo/B6Oa7b5
UFVmx750ABwLFnNWEp5JI2o7FyeaKhGm6EXZckEgrjp10xvjWmGDVpYeDVvxV3CO
jBY166zd3CUePFedwPTKzGSpJkxpEwYl7ZSeZ+AiLn2Wu0+sn7uoYycEWAm8Oaj7
tVbM5Gg5pZJ+yi9g1ICV3chmoLKENEj6WN4Ff7dSHM6HOm2g4Tt5EdfXOPy3phR5
RyvTLWpOsimEIhayDPZgP533POX6m5cKLVkmAmIxux+Q6CGW2bluoObyMDZytCvf
jiH6e6JoZqwoaXveTXp+PtljC5/ZGSltfpV9reIZkyOdVuODut92Wb9JHZ6WvWqh
2YFGZjOjQvXdl/Z1GUm9XfaEZdP4RKTihpNW30ww6D7FslBkSfAutkkv9v/oWT+u
KM+9ZsHhWFKW9euq3v9OGR+IaIHKAbihoDqoqkYeT/31mjUDEpq/6H5CBt6TSyl5
CL1p6ibUwBv6J6fATZpXdbHUaKWPrMH/dGvyZ3L+DTg4tIarAnzniVLmrEWnqHY5
4PfErC/cYowEgFruwURJycj7VKrlR5opOytm5TLnf/ZXnwlEKglMYOc5IPdQ+doY
Ufg+6jrzOxiFfrSuaWOacH8qkDhHYaYmz6nByZKoebkzYVZ7IgtNx081ejH+vR6F
b5UH5Rry/SDHA3GoL7rXGp9zZO3edcTRIcr/NI1SR5lBBJaTYeKs/XnYb8CRK+nB
LmDA+2g29jhb+2X6b7kZFZm1yaA3WZjWGodVp3077Eu1xdAgSxJ8DBMIUL0O90FB
Xi3VdJMwGQ+stCAmVs6kLvx4v36XxoXFvoNQPlVc+B6i5EIQgs8jmLHznWQcxua2
8B4QC2FPXapSyqP9ed5cXOmZ0YjKUQMk+KwP/5ukzW13HwSnI/AczsKEz20MAFGu
d/46sYUG84a6slUdYb/v8tF1UkLaEzin95Vd/qyXmDHe9x9dbFQqRL7fdn0ZV2Ne
2kTE3ZZgDCGkuqWyZ6/46YklUbvjxFpnNgfGuAN4m/oTTHbrpVqQG3JmYfTYZsFD
VxDPFqY8lrv2dQHehQauxCm62181Kf7OJiUM0Q3w8CKf46iuRzSWKXT/lA/ycmrP
aLOoN/S/03cLUwIjmKckGIjeHp+Lly1wmFBVCyaKGZwiuOwjhY6TGy3cTHhlTQ9D
sYtTNS1FHAxa9icOFyOt7CcgBduYxaAkovrYpj0vnqm7siMXkaSHww0dnGZw3SZb
oK3JTKXhKWPgavQoczQqerv2b2lIn+zbV41Yyhb4v/w=
`protect END_PROTECTED
