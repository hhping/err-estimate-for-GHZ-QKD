`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A2G7N2bmaerLxstL3UCsMDVDqY8o2JtO8lbXB3ZHInXuFPVvI2WaZoluHYBbOtrv
MFFO+elM8eKANNRdAPLGHbYUrkRj0GnkhFU/KPjc4GHCFRmnDxNG0gwMx/GD1LNW
4rQgfWT1VdXE+d1sMolwjzX7khjXfj8nt25ivUwyt6ivTW3/903WtQk2v4KOL531
6AUg69zKLBAG4QBR45hb5KdB31MqoBkdFerkGgtrpCZ6kaygLMAuyp5gmw2yoCn2
I5RxRhwTuEbyVadn/VF9Y1vWNkLIIJhOey+ZlXekyRBT+K/VTfJ8gYK+mppOJhod
Z0PvCxYDVvNwYydmvXz7Sz0CbtdXMEVL9ylHMGHznLxDLNQAkx272pED4yEGYq+7
jFbc9nw+8p9P9Y7BA3Gk626rlFckt6gaWmoltIf3LQdL36HzhMVRADcUa2A6Xo21
iP8AVgrI8mWspyqgpfozV4IZZjox2ZJGk3zKYDP87nUvfGdlHTaRs+s5z4DhWfQg
PrDeVbOOKLe5/syfJAxVKDywnnL46Rf35BFIbsqIRHETgRaX2NmCxhhjVH0oJJFB
CvdIHgCD7ptIW7iem9BcNoao69Qj/KI5YfHNSY0WozA4hjm6TNPTTrTacfywrNP1
XP+eCrpUTesSczlvsNZScrh20VfCp1X0rwOkMrs94Vb+w6bBKXmh7D8jZGirxUZQ
Bk+zjkODrikuZFRdLixmlYip7TjAJUTaeDeOMihjFrG4E2fi7EskqgYAmf/lcH6Z
R13NzJa4GxNPeDsLPAVtokHfgOeUITDShTCgFuJDy+YLQegeyrGpi4CGdk8UYfV7
KwgVRUH4+5WlfCmumm+SnGl6hbISUW+NB+km6jE6zBmVMLoczyOsJGS127rjE6Oy
ZAnWq6IQYmv/X7Ij4/E9nxa65wIAzrj9rRwZvIP3OawxC/0hSGj8jJdfTuMuqBHR
kfigCoImLReV++yOOXzZAE2mPDuuLcLB/QIYJYUBBqGHFr/yngC5XUaWDULe2n0G
T7YeIK8/4Z/or1b/AR0IvDGx/86aV6OqIRR32XZ5qP9Yg6/ZFXuWL6HMKab/xgU6
T/qSUwX5VE7caWoHwifg9uFJ8x3fyjJGKbrkSP0GXRdy+XYkcdyFVf4NYGvVO9K6
VAI79c43tB6N1JbPxURdA1/PnOR8cjyMSp6EMoc97Y1D43HICg6FPll4t/eD0VaF
p+WTCwa4aOAMly7W2pxvlTR/NhDJR96YmlsVqff5bBuyyxo/IpvEDiGDzaaC3A4J
QkG76yAFrdkorZdRwaQwq5cqvh1vfZUofsjDxv258WqWJYzLYHeFBXhL9YlRCnUr
zxMHTmAK4BLLiS0GbB2PqHDIiIjMhtwgnEfEFTNSRRjq6ey9xYlW6u6jz7HXj/ae
T0PUVjetZxKIq/TRz1vwmonLeV8V7SNDPGjREBLSTURYA4+UZ9FQ9nBxuY6Ua0ZF
e8Tpr3V1S+ddKH0vXpzH4uqSR0lO0czbk8LJ9m+L+tC44+vQACHwjYw3UdFSxYnA
7pkQ8sfBYNAuM18U/fVNEuxBBXTuq9Vo710jRtAaJAkryUSZf8YHvHFX4EJYkwJM
I59bG3cDH4OKtH9XnkCJle03rLBOiepFfxAKaQxborQIUJ4lQy6uhEeYBY+7Wt71
UOWe3sXJ3jvs5bJFNWi3W+9N3sgNQHiCbMgPie9emvtLmfc+dYviySAg/1gwR6DE
RCzSy94JIFMYIUy/ASL0+cNUdGAPqC446tKlY9Y7rShQJTy29btZARvZXzxHG1/y
t6dZeYBzcn/c1LUMUXM/s4U5dVxF4KaxjCKIv97dplQ4+cbLCgs0OOuJXfL2gDY8
Ca+UGCfhnknQUz/NdNroPELSaXxDghWfVhFdYcU75Doz9ACI4i3ZezyevGU4x6Fu
k87Q8ylg5/3C07u2vUorJAB1eleDylN7Z35KFP3QLr4XKHQxGrvZ7CvE7/0Y6DON
wRQAjSim9PfUpYiQd8KRJ4ypS8eMV02KR0kRcHhOH91OLyg1vKHi4TyeO362Fjs9
o9YV6Or+VqmV3vKDS407Vn4gGa8saNVWQ6GzJ73iD53P14TLVbhNBH+oWscsK2VZ
XLmhcOUFO8KtGJddmbueIxLEa7ftVhFpLbo608nRsser1XpwlE6zDNw8pwjCjI9l
pea54AJUtItwKmK50LfplgBM5Jvqf5iPYLEV3q7j4V9NNME8N4WZQuzqvV9zUl/V
Lgj8cmP3ZahvFg9HLbRPonTtOQqeghGAmE0SuMxrRDK8R4zVsaP4/0Lr1S/y/K2W
JXZBdqNptXQE8D9uwgkQAj9V7+1HnFHSve0VX/riqgfGyniy9f+E6n769E+hwn6v
LUovbexElDp01pXL4VL8G7n+R7DXdBAgFT4hkmWbSNaY2CHsHV8EfggGGt4SRDZb
cauMtb53S7T2vZWfY2Pxy2ZQmn7HcR+Lq1rVVQOq0hx2Edl+sCs/oe44W7dO8lF3
pD+OtO+VkDBPS5kZR1dsvVuFsc/pYwq2/OHeGUQMNFQtxmCnlkytWV4MbqmgOgdP
cr2TkWV3CfzwEIG5ALadg4FkSnPj3RdBCsNDcp9HLnwjBZULZh5jyXMAse4irTyW
snBLsCBd6ChuX/jcTXoua0sCKDHaDNQCtlbj9N4KHKuU+tzuBy4eIJeLrc1HYCy4
iCkgDkyN9YsPI3hTDdxyilGUYmNrL/2UyXtz7I/XEGdDYkyAQD5bQVS1g6S9YoAU
R6Ixh2PqGjNcS4rLvsqOOdtQutE2RuNWde5xDC7+scKmedvTcUGmOiE3A4QHRIWZ
4nlAeFcFFyyy19LN2n8qH651zXPddMAIyTVXaRrVr3V/dBmmZct8dNdZyufGx8SO
hC3c0wMXb8BJ89Ye4HODjFKzw00rjUzwQMq9sJ98NPRA7qQYdhL+lBgpZ9t+FpIW
HKjWdEmzHx9nBfaJA4nyGvCiVeAHeNCXU2SHMBj6nWtuxJb8pDUD5i8jb+YuN1Bg
P6UYYKIMQ23n6nDggSucaoQ4T+LzVYVit3mewgdBXaOTiYIE0NvVZo/72HmHe6B+
7fcYLWuqSKS6/hJwV80KmZnikg2ZX1BYJDJKi5JMEb0S10MBIHBPne/KfU2u0C0l
y5QV98gsOI90CmLLUSaTzu4tcR/6jqb7nqXfXEyGM3Y/D7V46ry9OilT/TfrD1wn
rzWWI9EDxEeT6yIUxpuXHFvjtz/MvVUR6/mxb+DvCwC8aGv71dRp/SJluznS4SOa
OrGknbE9nDLs20nNkfelAwBusLD6wU4J9cHoM8ln0H9itctEwzYu7n/qns47mChH
d9GCP/6W+oXIALwLwvIqiehirszf8T6rn4zO0P+Z7UNwU4WbFDkFnclO8v2g/Kei
rbGk48Utu5hqojud2PPmFK1xPHxha5ROGAQ8cYU82e9ZDCA71GC7lZgxelBfOKJh
wKodTQyUEwLisXUz1jCDkWXTkl8MTVLLft8ICLmU4+9H5QxCiEwNNQAGynAg1zdR
S12TwFQrzY2YGtGl5SQ9OHKqgo1EfmyJBtMGM1CpLR/C8+VO5w1y13cTZ1IDkHZ3
QF6nUR/O7ApqvTtyuJ7CDD7ZoRlsb0oP+7jU/DfZZd/CpYV/p/1J5m6dJs8cwLxS
WM5QjksYxJMGHxMUgGo0HNwEiqqMnX2TRXOoZIjyWbZ+Oi5vRmoiDiBUhLvzMTFj
ucjxgNv5ClRRSkWBc3mFz+iFyOQTA6plkRt89kStAyDJTStl4tiqqQDGh1iaP9/y
AQxE8aT34LA8PCptj53vQfeRapyvQ3PfQY9K8hcdsMQkAYNy+33GxmLNLKVguG0J
1RZ7H1q1+J60+wxJ28BFCITQKn5e6LlqQwDK2BKUHyO8iEAfSL5v1bIZb//eo1sj
F+99fKZdPFEe7aRo9NrfLfSzAlCUYcn+GeJzYvpeu/Ulj4iBQH5hxgtkA+X0n8e2
HYH9SgElU5Fvyguf3u41u4L0wHhde9sw8Fep/MwGvfuCCsKQMKne/zr8URZzexVG
pDD7EiaXa3QmjIyq0eMaVcOIHeeqkXyMfrSTikRVDPa2I+y+l6fYu2R6SS6vFUBd
d1aVkk3QkdvJWJw2HdTrhB7ZEl3goU5z5q+thE2AxqtbqCExChkpYp3wcBwlgNgS
yCoB6VGOWEpGoobpi7B6GkLsu16xuLiG1OvKFWUo8kYD9c8FWWLNnZrdb4nTInDO
PHaw69B6G5b8nm1hfuf7bkDfux8RzgSnVZX4gg7fy2MQkoKG1klb9kgt+/wWO70d
HMOQ02fcrg2d9skGfl78jJqQCHgoFki5t7eSE+Y7JxhvL5OQCuxJBFwwv5TCF/Pm
+ZWWxzvzRndthpOQQvSTqS1JZXS/00fVMFPNpCyFCwXimh26OfhgzKORYoubYHJt
xH1vjRRzuiRHzJiwLS+7buv3bVYG0M06/odX1rCNlgc2pxeEfEDtRYRWXvXmdT7w
eoDoJmPyVCwEbpmAcvhCuIlNxgTkJUiUoXEpb8zqqWRfSmhRUpcdm+su4NUEj5Y/
IeNoYy4HamHAXV3CGOxEv1LZHVJBwfBhaNlPR+Yltbn/fW7r8sWsYAfV85dDOq4U
edjd4O4aWb3dHRlaI04I4XvuBuh8HaXBPa/r01y9OBBC5EnDLRcv8+pRjTiqG+gN
YvTCl/ZMT6Zm/AJuaBv/lmtQn9TzcHfwFKaPMKDkMta2pf3/t0riq7LdMaTggv4j
e2AsePJWwOpDwQ3mur5W631jwcTfvEaVpWNfNM+Ia3nsECEGyXydC9cWfL/lzdj2
GJWanlakAidI+gp4WvvrgnZMUidAIp7+fdAelwkkwWipCe3tp2ldzQrTvGi9OZfR
LYlhsUrOmJS3cckLDz3VGppFVwAmyYO+1t5UXMqpW5h9oQ3FilS/5JtMo2Q2fplA
BmMVgx02yd17Sd4baql6iAuW/3JcOg0XJ9bHiVjyR2ZLJCXCKEkh475UaYoma1nt
uBded2fOJ1nPWKehrf+9M1RslM6utm9yN89+Iw4/TqoR4ZNsBwARngMCfgPqFLPv
5teL0W6cbB6YpiicMNGyuwXxRRDu/YVsUtSjb8CbtjRhGnrHCVULnwkjgTrGPe8p
BgAKhLFPt5XtrMdwp9KYVw==
`protect END_PROTECTED
