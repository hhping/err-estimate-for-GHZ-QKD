`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PDdy+oMSfh4QjJ6S/kfMtgDQ7Xzhi2tK+jSAaFeUq9/35DvahpyTmbosEVcDB9Ph
BuizoAhRrywgvwpwOVIioXqF+q0PS0fwlwjSrtJs5o/TevOoEeymYhD4X/5pF3r5
dBNXGBpSa+TaWAthWx4q3lKmGNlY2wPzkl+uvwsyFx0amqW21NlOcA/nT+S30/rS
rQTMAHa3RIkrlhjpiPrsQC2eWpXBEO/6BVINE/fnAr6xTqC4Uu3DAVX8TbGocSrZ
O9E5Fkw/z+lO78MCdKWVHie07oIH6ACA5dx7ji286sl3mZos8/4U6PpWgEqTKZt8
sBBTU0eh/EQFjVdIPKSETKxDxF8q/ku8WHB8Gsm2zo5cS+8g6K/cYx/2bdIHqkSj
DAk4sr2cdWBFY5070ZR78w==
`protect END_PROTECTED
