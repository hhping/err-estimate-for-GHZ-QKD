`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NRKVO32AWlXerffaDdy1MDvlBEbCzC2oDKAJDuYE1PP9//ntLeQ6vRJigKToutBf
zQPnO8yfRoButMjPfQ07C8wzHfbgcuaaZztQS3CdO4VYC3cLHSsJ44KBg45LtVFY
FSsi/gFAUlEu4hYSlaWIMvFS3P/wXp8KVdoMUjhBTMnGyR55j+Gz2dzc6f16b10C
wTGJVaMMAOku6g98NimkzN1xOtGso6lkEb/txx8BWY1NXoJn0FPzyZA8ipAulksp
IWXzKzzobNHUiPwbK+evx3yptbRLkApX/sKfx3J878fQSXkEeI/MWsQKNktWiEJ0
IgannfNX+clXEKFy2J1wEmH1cPx3PqwPxcOXUhVHCSEipiLq1LIG2saEjVNL4QdH
Hu6tkxvBJEmt9eBRRxX1fZCW+A+RGeDLZYhksNhF/5hKtVv6Smu+CNd9zCrIZf+Q
fSnrsXrjIPhAKh7uHwPNl6Ia/XWitFhjls9JtzV+o2qudm7rLDY6f7/ABQmb+Byp
JpTlwggi4qY1IbBifY4ViH1diZX6VFW3zH6+ZRfLYC03sspGd9W9WYN1dkoBtZnA
0uc6EM1pbqa5XAAYOnPhGj9cBnFKKy+mUMudKZmzM8q2k+Kx1RU0Mw11Iz88nuT7
5794ip4ACMuLEFas3UyspOX9rw950TSD/hlfCVNl3lVtsUokyXA7NywpkBKwhzg9
9AEmJ0B+ZFxJD8PqPZSdrkIY3T62eydL9m6gbpn1r6tqiIf3i/vFTjHyFmk9v/Ln
N6O6wBHfdNjl7bqWqbqEqMR5tpa2oM+fTGZtkX+nYJ7AMAKpqva0/8K57YpCyhpU
l13s+AAlFyiGPCCYXwn9y/O2JV9nY638Ii/beUi63XVdvXHHMrz1CECY86kx8Reo
lWZeagJnVTY+szocN0+XjsJLg9eKA+9INWsNGsdj1AzSvKRy8jp6T5gogz7RswCg
qSaeL9LvFCafnfHcmRcSluYMZjrF2/6mXqwu0OgESDdiJFtvK52FIcC116NpcJpm
xSrpHlNktm9kl50PPy4SDw==
`protect END_PROTECTED
