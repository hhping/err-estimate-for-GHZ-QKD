`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1XGt7MQR0DzxNiRJOFhB0xjL3bJO586/uX6UsOut+oD/Or4t9nIC7f6c5AUwe7Jj
9MuRND+PaMkPJBedqAEyzNgqH6L8070AkMCjICqmM/cljOM5S9KmirQp1RJ668H7
aO8fT9Xetlyn6x42fuB9ume/R+UYXgm5XMcv1L0wKN+0X7vNYH9AIYLnqh9aOSSJ
0E3kdClspkQTzt4RjqswKmCSNGzWvYF5PDecqw+Y+uOJ7SPctLWV5zGkRKZJbLEx
AVib4tgrOx1snssDmlfJUiXydVYGm6sWUNT2jCMezwo6pO+Y6m4DR/KZXxkCXJUi
C6mLLR0ip1u3xEN3Mzja3IK1v5WXE+PPrVyq1gxIGO/xMx5uciC5efPTh+4S+4Z5
MFy6wTtmj4wxV5pNCTcM60LLnTnyH9YlA7r8JTo8EJL6+8TYmduNteR5Fsnck2MP
g77MYUWWpVFNoglu4ChEjCXzAKwYddDJn9brcd+O6chtlVmdkgEjQnLdobdZXGdG
bD14A14zqPV9fr1AEq0+ocPrXPnPiiqyJpZVLpLc5vO9Y2lmjsPK2kfaXomnfo4c
bptT0b5QXwT1Q5DTA9tj/tdERtJHgMhb5ceHyda6JqYxclvdgZuGWTCyUFO/xeyA
4dkgIUkCnadRA4DTszdh8wivwWV+FS1+VoytL2QAX9FxOm+UlrJjVl3/jh3Dp4Rh
yI3wrm5rDWqdqF0dU6R45ZxDzF+O5ys4JvcufBWJ5NxunJ/jtcuXb13e0D64BJUh
G4Up+bO0cyLHvOHSzdtTp0fbgfAhRRSqE82hHk4DiVL5/PkIZPMASpdkWsNwyCeC
08vwGCIdDer3T+8Gz+18Uo6JYQXXOcKhSh7kPNighb8T7qhC26t4R7cSIDNQMdki
kX5hZCD/RlXovPcJzsaTGKkkXY9kvXbxByA7uM3szulKp2SyrXi/MkXEa5fZ1Wqn
cnAGSibaHYF7C70dc8ohiA96IrC25NH9WH+WHd5n7JIGOhfn5+zN8gWB/IfBWR15
oyZ4E8EV7MeLbSSnZb2hXbsX665zOHfRLsB4Z9MZrUnEnVNee2udDE8/odROy/rj
ZTNhs4uWOPzV8m2KcT5uh3LDAO81CVt1gl5UQRLzIrBT6JlOsK3nHwD5UmSqKFFJ
0akqBBc7N7PPmUKMFSEy4jIpP6QE+FPfncUC73ghxDL5XyQQ/odQ4TAPXZ9et+NN
D4ljvTae66KZYzQPRRiiY4fec7jjduyXV91UCsU1shc=
`protect END_PROTECTED
