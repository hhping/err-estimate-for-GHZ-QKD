`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
buK/AHpiCSoHlRRobC7o0EPChhCTuadG2fnHqXOdcK3RdIcU+p+s1v2OFtvCEEtJ
q88PYifrLCERRadsLCBh9T/Dd7YYpHk6i/a/qN/E3tZlaxpdIu/UaRkeXCx82Vte
Nw5p6QKK0kEpHGjUyOc8mNhLf3VV8bMUME859bqYQPW4hGc0B7AOtaptYDJjqBbq
QcAl281EL/GD8vyguXmoxLUJ95B1zkNdnJpb4pZ7IIsGNDb69HoNAT28DubpSieK
V5KOdX2i90Whx9TbRL+IZ4qwdo6TR2vYUM02miVlYFijxY4254XuKbEhSpv1gVK4
M9DZ1WUs2Od1qwhh0QxtZps2HkiTilICTKL518YI4FFxELYOAp7e4/bC2dFDFY3+
Q0rqJBFRT5Z9DP0RJn2nTWkF7ACrLpekogqvw1GNoVJ5oSqd9l0DAT9Rx7bOErKr
qkcDNpAICyHowvJO+hNYtjlebFB/ioEQHadM+1+3y6C757D9mMN5r30YwhBJuHj6
c/AoviWhhDI0enuj04Glw680mI7hfqNJ/QcrsZG44X0U7m5X49eLkVs/mlD9FlrZ
TER5VL5IFw4dr7+/OWJ27+WAfZ1Mri/L2Uq5hR+jzri/+hjOXK0h0F6rwi6CpaZ2
C3jwI4s00PJmbY758aMbDxU6+Oel32HXj2WX9xyQwD/Cds5rT++qvJgY7phkdTyv
ZiDsgV4o8zxi3nDLV/TuM66DUIjbCvBogAYoCeFEjA4GQY4VsQi70cu9cYoNz0kX
df7pW6YiANiJHz4rMq26JRzgXjaecYHQZenR6lxlSAYMgDw2bcljB6s3/9d/6PX6
RDGWrP/4dVsqx7VGJVSjL6Ny6Qw7Cf5/lMXoUDdp+e1zKhOKCM8cwG4lFyPNB1KE
ZdrL45wFP3wwFTKVZ2J+dzxsDSWdX/Nxse742CyQm+dX23teUy20xRMEi179zBdd
XZdOz8QVH9ZNYdGIDeXEJsDnjdUrGMco65kRsATZqsQWUOE5E9ro8XYe0RapsAoG
Z7MaWo8CtoCKWSEDMZDmbWfzhcTXBkGtx+DgYHRQBBWzvGKUBjJbGe3fqoTgbycw
7KYvMmGEUacSZt5D+n5D38VXNki5lED47CxskONo4qsA7hSHJamQGXVvC5ZXz8tw
oSE79D9OJA9+7zP4JarMbcF1p9uj/TjnPjrnZDi+75Jkjx7SY9Hs9Ug7kQe0xi9a
zGqlmZWlY7lUTyX+tInepNx9qdZxIl2l4eqmVXEgY9SkRyL/Y+RUjjfOJvTfMEOU
Dl9Lw6cshoAk9lsROgW4GOCrYGJF1bESpgKy30i/2vR4ydxjy2qrpDRfUEGZBIt6
`protect END_PROTECTED
