`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Gp3QRr0vqOHZnwyfkaY18wYRhtoVs7sNu2LQj4hakTWu473DxOR3gGmZgmTTSSR
VTyqhbCdPlM6JonYQmDF0DSFXAALq8lF5Qmyid8G0ClSsbzEJM+D6ew+gy6t/qVl
U2FxJZotRYld5h0dkPs6/nQFdK1zgf6gpxll2wfpVoAn6xUa833N+gdhiQeRxLN5
HkJBexo8KOa8NBMXHO7zLg7szM7tuu8l2ATJ8MseOo3SEHVc/dvntAHJckBasd5y
UkTNXau44X/4mz1yE7MC3mSQt41hQ3mdTVaC27kSSRqIp5kkhZK7MrMieMqKZ83L
KckAmRB0kf7QBwhvb+WuM05mujNQhNgi/ckqVU9hTuEaBtRqO1wNLL+cZrpCHsM0
Ez9MfFRys3BiISeUG5g3UjLIdXfbfssnv9pPFjdjabSzWHhFxLa8HnO6cutcg9dn
uQVvUYjz3dl++mv3uZlbLUU77eQ/N0biIX/jnMwPxsqDvmJ7N5EirHFR3TaIJ1LV
NlK4hAB9mtje8tz+AIOliDAfcJN8cDtWT6PXq7Ag1JktKk2qFiX0Yt/li7PTe8cF
GIK4m73FwZUufMR/U6OssUSa371cCfFGZnfnoD50GArchLjwiTk2gmrDHM8Ewjx1
`protect END_PROTECTED
