`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E6wmIayDCPj/i+w8uMyK1yD7ONlcJs+dZ0YBrui7xE1k78UhjzpjlyBiUXk2kmuZ
8lkqj5vd2MoI7203Qnmf0jXdDOaZUJx0Nq2/n7a3llYbwL1C6USembGZaG7VHxvY
hGYNRmDFmy3BowTdxktOLDXPa2a1Z20GCIoESXtoD5lO8NCdb0F3Jjlx+cqy2cDH
a97doxxJoJ6o5nEXlpg0cr/X2LeFl70Xti9Ogo/zFruWjAysYKsVnGIz8hZPtmJ7
JAIvqlJfy64OAHzOEUh9ryrB4UX+PFjLt1n739AE38Y1UhoDRP/7moqktkA6Z80Y
jwMO55U1opSJHn1tE6I3CxDZ5qxT7eoDZ0f5YyvdzgHJlFvv6hzHii3/olBJTBA6
C+wRk+igfZFFAPIhiEzTdSLB/NpQjLw0xDgbLBy6M7KMinw1iX+jbJx2oa0jV+Jg
TJ0CplGwANI2XbFzCu/kmyAt6PCGv0jjh9DikjBWOULdWO1oVDEHITM6AP7+pZnl
Npmio+dY/0oKyc+P8aIZWGAMhlZ36tX8uYIcJ6RAMPjH5y0SoVCIcHEqH4mrjbuK
JIvHaRWbABHAgdo3T975qV7OUBg7h5tnaeVWmxx4RDcfiov9h91bF/H6CFB929ZV
VE6sCWdiOw+vwI1OnAS5nnOR4u5ATLNp1EEsdHFTel3Pg6glKZUqqDfq+9TM+MUE
+FTjx1WLxJDPfzDrHveRaAn1m0nENahbXJkvrpOHATMnEw4rPjclUV/+QTTlwtiJ
2NDHbR7zi64lpEHlvOyqwECR86ZolQHHs/V0ngNVDuRrClBXwDVHp/unSxmKSx3l
rspjDbhJu22Ov8v5IpTJdufGHvziMwZNXnKOSU0pNuNcvzMRqtAcrzpskmgcxIkn
/HRviGbnh8frCscpMpmeTzZQwqGmTeRqXsrinIRuPgkzTc77Sns1/EbVtgwFj/Oc
rsuz4w0TUAjVI1vGTPmwiEoaaKZbnRVbexgdHUchg/DxXlO1CD4pq5y7JsZIoGBb
vhcj+Y8kA6E5pCidlOePz4yQIFNfrm7xBy4yopkrtRi6908iF6n2OStSkKLFbIi7
nbStwZcGp6qzfyxaLfUDOVb28zGaD0qBH0xfvs/E5aN1eH8KwKAZQWkD6WveHaZo
D7GjV1OjA/oLBx9/jblcgwc7PNdRPVCIWTIblLMiXWOzVwjj0d7Wn4CLvYINoUGd
DCRm5M6mepKlX4ms2qvVQ+p8DR5LWwpN9Lx05fgYLtNJShIlHEbOqapoJnHqouLR
mbY49eKU1SHa0PIDNIRfH9w06jzn5q5Egf0p3GSz1oNfixPJCAPMXTnsWv23vRvd
`protect END_PROTECTED
