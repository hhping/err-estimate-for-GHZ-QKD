`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mEW6o+l8tGUlPDTRM0Jtn/8y3T/TSMmfP7qPkr7cYYn75AT68FyeDSR9spPsufIp
MACq2caLFjbSOfMkOGbt8srdEbcikKG2zmoed7eAoaxviGCuHZzNtzvivsXUPiQC
FcZ7MT2guMQXw4TE098xvHyUxpIJ6IjBHJXgjhiDI9vQkxx09x2GE0wCHNpcdc42
7zZ3b/41Tv9N048ZPjIwZntn+wGnR7IAsvA1Ob2efrsE3CL4yyRbOuY+GksC7W6i
/kTx1JJ/OUUj8xQVc4gEbSPrwHoCpgPMk87ZU4zxSkkxdcdMfQeutGyrrSEAIkyD
JkA0t0IlVmcv1LxntYaTn54F7nSsy1QGHNxXLucuVVdCZefYwFlYW+y3+0i9toIs
brP02aVOl0vf8fMFyU73wKrGoAASTP7oLdFeuLoZzpfXnND22eKHhtUNjN8774jj
fBWmNDV/IEtmDLq/YRxXI1tubjFT95WlZ4hGJcKLYK+FAm/948p2/tkerK3w3i9n
zfSveq7VEWRhmzfeGbwVpygifBqpglzMHrlkFB9+xbLKZ5oODuV9jULkHpmvTkuK
CFttcDGn/HZqzrEymzh4n4g/sIgd+Lbf4/xgynCDaa55+jD4O14V+NQq+GcoZ4lE
F1kyHv2RsnFAJYkyrs6ipUbHohNDH3gS6dNOL+4M1fZJ3pmNPMaVMnqBII4+Sln+
tijSxOqD2cEF6oSVqDaeyIVt1+YetieCHnkz95L/kkcOiKpz3SEB5DeoltuOBJaf
ulIPPla6vfSgVrLBNeGvA6N8K1ObOCjQY0RI+NCn4wg=
`protect END_PROTECTED
