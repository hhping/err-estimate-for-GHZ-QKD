`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jBfDEFTgP7wolUM7telFXeCbMPqKDx47aMmSxn7Xg4DCkaGbl5onpya20FXwrSXO
5iMexuWCA9/rStvXPWB34WoghbNxkootaVl3dVfO9ONT+8tCDSxVH7Nib7jMXBxT
rGAD5jtAt5i0oCwMhAwZ2JRSaG2drrFMU1O2WK/GYVkYgtZ7V6gcbCvKiT4RSPZT
xZ6AYmvXpxNVKq5w9aIdgnjRjuOWHNX2shD29IqVLOSteX6vVOwi/iY35mj5q0aR
yufQtpxe9L5mPqedR67PfrPwSRsquU+9u0diY44IMdMBXYH8GJLm+IOFXWfPKukU
UXGp7wJo0UTQjz0vPQ4AkTLlUD2ZvJyzYtASywiSWfdDSP+8YypNHNAcYmSms2fk
5uPelAPPwOjBfANljuxp8ZM9DEfwNdspxK2HUcermvMkFuojzrTYCz1Ke/oUiS5w
8wN4RlyDdiAnona5hcNxM29LyJcxScDkdkBk+ayTvO01f3vLQGgqR7MuQ/cNRVxS
zqA+t5bmYHsl+kGb8N9S1S6xhmk7zUWtVD/HXDKNYsi1C94COFRKnE2YiresPryu
6ko6Br8sbTgdP86XgJAfkvsJbiaXebvXp4BvSo6R1bQEkV08H7Wcknc4QFcUm/H2
lSKcQzHCqsmYlXHNajZyeVQ7rFgyvrwQ0PaQiRLrSpylWPOG/NHaNjaklpLP6nyh
vwhi+Cl68yk3189vCcAX8zkl9hyzRkVMp+AsiXoRZgoSvAHB8Wtx0vldBOlxlpp5
Y7EN3qAEigCYYo+RkX+9z8zadSb8ugOk0y/F741aX0I601Sy7sMGBJjmJKNiK3H8
bXD+2XAfaVKFKQXwhkb8/f6k6yySsu4blxZKtTvZOc5aV9zmnr5PxjLsjNCGyjQ0
7kt56rkGQNm+xAK9ISYojPUyuY4bnI3aiqTfXfv+9/uxDm/kp7VhXvjICbhORvJU
KB7OggLH3iRnX0n+04PQjaaNh9ZXFjce83OChUdFkv66ntsZYPbl63pthVkfPtYQ
4DVX/+XbPSjkl46i0CSMPYJO40TF12pusZZIunCMSjgtxCXT7VckRVaFjF1yvafo
QV+BxdWt8gN3Akxnbr90DR00PFISHBmyCbUoEY8wGjjI+z0FrxPNiZTizwtnx4Mb
gf10p/EN5Qm4CzF9yWYsfIUntPgaHskXQh4qrKTGu97BmAfWfj60o+v6JmZyP0AO
jC0c9v2KHEGSqjiSR+3q2cL6tYmJsubtV6Ffte4r1pTN28NohfHhtNRXzXvnp4mw
SKO3/02hgdY7bGhlLep7UOSqMUE3lqne4kCPqPfy512tVi1QuIAquDSjFJ8fT9tF
yZXBI6lv9SENkulwYUo7uNRfj1tYMGRVUJeydkr635DCH+oIzBYnsvmA2acm2tbG
ERZrDZPdIwVJU8JriKm7KRcKnAErFRqShOYAkG/U14HUPc33euhuzmg+wG2tNiDm
EkWiqiHjD1TnwY5vCBqnoclcSarJpxhPnQ8nr2shIzXPmZNKSAVMm1jbBbSLIBor
M9KBZcTPOPJRJ3iJI3WiIA==
`protect END_PROTECTED
