`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sZpFBuTAsTT9WJGANQ/XeYuuCUc7l2sjSZK6sAsM/LFtM5mg3gF/XxzOLHY/x1T4
VsVfaxx3C8t2EaibYoUuGH2EFelKZ4fWVz/thHdm7/H700BZHVZzemjeGBwXoVKC
ggxou/Ty+vU4Rt0oNq7yGXgK4pkgav5kgyyAv5M9kX6He1ztxJc6MvQTexAMptua
BxRzZ/SKipUPEUI+7MxK4GbQ1aad/RTRIEZ81fLnfpbC+rou6N/daGxaS/fGVF8I
/sCX3+o/QQ4eKoYJ88eha847K0sDlPWveeLHFRiP5ds=
`protect END_PROTECTED
