`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J5eslr1+rBKpwMRIdoaGOaqRPzbYL6XHJ4rHoNne4gIMkcNg750vC5wsJTpL3d5Y
l0N4XThb4YNxTshpIuXPMpdJr72QSuABi2KIdSICxDrdC/Cht1ADPEHLEBI4VJzS
fxpndMWvhHwJtGR5o52HXBiSf8IbjvYwox1UJZhwHa5A4AWN8RjhI49VuJ7M7Wg+
xAzhc6ks3oKn1/9jM2Mw7A1202q7n7iDYzxE1Cv2KYbCJBSMxReV7/QB1OWIyNcD
bQsLNP410+4sXZakBQWdxqkLYNNm5AVQ71xqFo1qQwUQ58ABUm4RPzyIsDuQlCTV
FUn3y3T4d5ZkoLboYmOT4N70d3s7et0vO1ELFWok7NQTPn+HV0SBDnKGIUDabb4q
/qGSB29/8HUTCjlcP4CSZAkkNiWA2QTqE/xzK1OdKnpjDZokwapC7KBL32RLAUKt
v/pl5VW6k0u3gNO5oOZwrfVb3LQokGGiEj/fzsWUKmseG9jvQUUh21FbpnU7qzmH
FLIZcUuM4pitpyrFCjUpCh+Jpl8FlR1gXFI62B5pKHTwzscctgPQoqlHcmIU24nN
t9J+og/0WdqY6fK2A9ryeG49SkWAveGU4S7sKXwqplpocIEhLVD0VvSEOhblvNpA
Q1JY7OulVIo5E8BN/szfDDD5kh4ML/AhUes5gEW2kSVIVSStXQdWuMmX5JVfsFYj
FWHC0jaM3Cf/GTA16CZ2h8P/qfXW/UGGnmF+r+zCXJdOqo9RM+PbXyKCyUi+0n7Q
TX7gv/NLDU/4MnWstsTyeQ==
`protect END_PROTECTED
