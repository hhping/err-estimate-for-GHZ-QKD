`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qm3UFVTkgVBpkhp1RrMEtF7IrSNvi84qqvbo1L9h8890ki+8kLnZ9HUn8TBwKqq1
f7EoWv6iE2MzPeKX1M6mJv/wB47pOxmNd28FK7PPNw6cEdSg0BuCaDoG7sJCE01k
a1deKLq/lSe47y4CPV91wl+hoQoP3xauT0gRoswj+z9ikAvhZa4SmQF34KkqE6BK
bGNllYaN1fVoMIOk8+PVoGU/66zRzM/NkHKPE8ki2OjBW7rCRagvEF6IY7+lk7jI
fC1GuGsN9W6YooThByDzgi1vZt7z9XILhPAqUVF98Zkdeqn+Yb/Fy3ueHq5AUl6C
rMrpoIAMzPxrJPoS5OwUBoDD9b1gjrbjc6Qp3tz0cFNjj3VQgapmJrOrU0u4ZvtC
+gr2y8c9ppvQhIj2YMR1DASOOMNJjb7Vkjz76pfbbvP+QDntdDgvgYTh3bRUjmb/
uR2uXP1n3+2ny2F3Gosym/YeRwfGxzrzBYVsJUFuU2cJaL8M3tlllyO1LuU0osqP
UhIeT4Eu4ca1HrZ9j6ABhRQutRuvtIWWwBLJQTCH7nR/3AEXa+Yt57bEzi3lvMa1
+AmD2v/nbJPt8e30Q9wXtu1uqImRJkc+azvfHZBFTKMNYlegla5GB17bcaIusf+l
ptyssX+ICQ4MmkMqc0aRe58mWyKGvIYtvtgb1X7GO2hQb/OgrhBox2kc5wZOinHP
93UONIrwiTeSZCyuUTYSqzLkMXkEvRDGo1axgqOnREybPdOmkVHsSR/TesnImmfD
yx3J2KBmN7jjlFqyqpi6GxDkzMREmrbjkVANlMUaRsp7YdB4JkM95qppHYLQ7iQo
IQCSdthp5sUbQwNGkuxzMOrkokJJao5iBn37NviyDgw3Hw/hHNnMZYimxNevbAYX
Z+OW4tdeoIwb3OKXrXSnQQhFK64epXRDR+wUlcvzZBSsZ6UHfzO5sgIhBQTiG4Sm
riJn0clx/apGeJ8xl5WQm+0WSr3al7+xkk++TBaV+8AtHUaLcYp9J4HaXQug6uak
lkQKlJRXVfxD/c63azABhs/fvLK7KgQg0xT5KoBvDsuq3rlXvzbL0LujoDfiV73T
GYeveEBe6rzbbKbgh5pKHQ==
`protect END_PROTECTED
