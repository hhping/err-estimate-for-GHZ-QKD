`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mXsImlRmeXCwJhTTPeZAFnALpiXh1iQvOCvV2c7SndNGr8ZK8i/SKZ2sG/b9sSLk
YTewSQDUgL4uUe91VwYMCN1Q/HX/5Otk1p/2mlKi87lVUfpYJWwUL7RgesJIQc8b
iwNhGkAQ0mgXdKmQqGXFLir3XlUQ5YJnY9A4MKMGhSzWVN9/vbhYj+hpKO+cvfuy
gPnbLpz8DjtXKx7LUv9bXVC+yQTwJs8xlu5Rj5csv6d9iC3MUs64+Bfyq7hD7yno
AaDeh/bGO9FBBYIu/YS9ZD+IgN6OroJiaMVgz2SrTUG3ztL8QThCfl+rNrnzqZWP
0Tg3zIsG/b3Fpp/LeBnhS4xKAziUq6wg/QJ3VFxiEeeY8SwX1MYdrzH2qfPBth0D
G9fRM2bFqeTUxt0mR+4gMmcusen2zIZc3lxxtbjHX/8ei2jA1PhXwlsTw9sQYARU
vimoNfq6EctkFt1F+Wxzl6cZWPp3ybUHReNklkhkfl218s6uXulZhs2z7c3TVGYv
RLGrTpts01F4QJ5TwD3j1b4EEBk8NHObNFuREJ2Hdp5ObTDUt0YgSeB4Q3DVo6Fj
LTyn7YKgUK6ZOJpbjsma7VLqh9VXd9WYGTg1NOCuIVvTuetkk6Mi1TSftj7sTCpd
Ayxmp9hNHUll4OSu+PwvfkF7lLQCzvLrAeFqczK/Q3qjI7c2IKD7NhaEougHLPSj
HuhUVF5esmAg0coLAaN4/3B1nWF2Fmurx+LsyS1q2X+M8A0I0vkM1jb0CStK1TrI
ZNPFZRLdK3C4kpKavBLl8Aei0Ih0lBTf29Gp8O4RfWhFn0ZTUVtrLFUwnBQyhDEt
qwLVGbDoMwVFysRAvbHmmQJs4jiWqDQfffW6vEuUAtq2bh2Ik6zVM83GMxTp//Ql
jUkNGDgh0bcSRi941B7ebEgMC8O9v/ZeUVQX1TtA8W2WS/HLrO+lrKvhV7ExyYoO
5P87JecmutokgYfNjSo6UXeKLLu4U8Riy3dJk15VWmE29CmWV7mDacI86Uu7aeGU
W9jw0nEodC8PiGVwrayNjgHf/TTVdiuPsscweJC5Oe/snyzVnqB9FIcf4ttApE6l
agSb3MEP6uKRvXYUl9pB6WTxBGgYn1wAxQLyUmk+7WetbsWRCqEaDG46bUgOgheo
W5gA6ksjpsSaRsJHh/EHdJJowkmjywGDu5P6PkiJoBgQ3L27B9faUGw+I2jYNIh1
zRo3+SlWVcwAZ5MRxfxK8xvwGQEjWjxrc29ujxV1FYy48H4RFDUL81DBOheMqxAl
shXeHa9OsclHDQemus9xyosX6pK2DVmYsnXt08Jshi9GpdjLUZnZtCrTiBRhGd0B
GpMEhvQmGBwFJg1Pf5Gq8ga1TBULrvSLtsmqnd23+40WUGWcHRAjVKX8t1vBYyEb
WcS7qtrclQ9yVk6bTvsnEN55hcuOgOPYVYEv+YbbjVOvGKI3RU7kMia3O2F/TUG3
`protect END_PROTECTED
