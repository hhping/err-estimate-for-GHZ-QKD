`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LFZP4pRv0xYBML9w2dYAzqZWbHCAexbWBI9x6E/I/2iAJJ7sC5hircJxGBAna/9h
jBU8NwLvEjC4TZ9XBMfIx/ZGmsNZzMUCPK33miqqrsXGju4rX+BaqvGeOgfLWOMV
8wx2oszi6uCOZjxHCG96WS3q3yFwnEUfZUC/UV6QKOsNwdHPDrWk8lbvngg3Fr35
7UPFi69Tc7W/cqz7QfzJ3toVP/tUdO64tKSWrbLkpA3U1cYIhcIn337p6qMLEhLl
Bko8dVnYw1pGUan1M6VInCQZvGdF2ttrqbW6VeINhS+Jt+sBd5BxS60RUexWIDcW
2rY73+1zstjAoLDO9V/o5jr+jIdLJqh4/G/MJESgt1mbcEnU8NWGMupe7dQakC87
Eu7cTKUbbX6M/BRBRt2n6uI8o5H97kTu7Y5CnilfbJzr54+CA9C2nx1H6HfpAmlf
WeaHWiX1uEr8cmCdDtDqZoRSSoQNN7McgWQj7HR4PpV2EEscMDBYGWZJuTKLtGQF
7usEZL6rBt/BeyB4ilK0HZ7NrPy3vyLh77orQBrBlqP/JHJFBzXVKM3etCItkXDz
tBsyNhdwZc9c/8t8uwy1JxS0U3pztUEXLVwvJGfwpaD/4GcrGfrsUQaDROFM4VW/
fwywMDV3zP75XFo4OLhGxYYftzU55qkK8vD/NMh7w3IhbyPkoce89+N87a7MUfQ/
pIAWDuAJcKBb6hqrZSVFf9rB/PagbgWEksm0buOWsdajfNq6IS+euCei+7F+1U7i
QZT2tiWKhx+mJmhepU5w7dmgynWo0On0eJLxfwC6Rv5amGn5WJeDT9XH0foBaNF2
vO5UEy68O5xIZWL4nnLXGhfR7eWm40Ur83iH60/KHyuthe5Qh6R007TZI3wQxJ2Q
N3tqzqXzwMCQWEVsp8ac+mW5igUY3dIUFj4vW/LTeiynMLmALntgIlFXECfsnNv+
bGayXmBAl0WycjIqOqUxEomschoUeA/Gn1Twi0MBoF4=
`protect END_PROTECTED
