`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xu30cBmc8nZ+Au22MhyRMhrAhaZPr6KSK7ho/WfIKAsiA5K7ZsCO2H6Pv6fb0GdC
LAExiUj0ZW0H8US8jsourYhqP+IRmJ71u5NRiqaLP4uJpx2mhRMXfibk+cGBJoO2
RxzAejeM9zoLFV1y7l/cQyZVDA0gEsdzjehYImVLXLR5s7XvpLxZ+HQbN922TVcp
RN+qIRm5nkqRGng7BJ9CdGKcdVv9jT1t/E4oKgWAnMRS44jj3m2CbUv2OSfru3aI
u+pRt2mG59GEB6J6n0tskxL4TZ/jGbETg4Nu9echWtNoL5F0Sp1kVx5o6y8S1Igl
Fp7q8sQdek1VuJsy/mkiQWGuF3oOkYC3/Qxs9pKN4m4AkGTbOJdo5830rGl1p7zj
jJPoDpWGV+AFCj3kQezi3ugX5NqfN6kpK3Sl2muNN7SVadYOqDOQNJHpn7gng3xa
KDLaf0K2L3XocD7iE26XJ0ngJayr6H4WZM7JsHzKyB5MmsD6Ek2EhmaKnby2BSiD
we5on/2qhfO2SiMYReWFpd0WutNcVoPhCv82k/sy3LGbx+gM0d71NeP4cE8xiA8z
lg+4ySacoF+B7EWXJlsfew8JeqHTMkyJOz8AfEhkUridwsLrHzYBm80MWzFbvu/X
4AMPqDTbncnve9mXXK+HBiwTQQ4hoO1kMrpfZBu9+aoDyrRY9mhvA1zTn8pQsDn/
Jhds5iiDlTfYxiF9S+l8+lw4tSLfH13g71kQf4EvdVFKloHU3V1r0HYrQnn8mT9P
Fu6mcpBTrUo9vkCIDsL8inFx70zVGBgIGlAmsfpshGDEX44hxCz43zHWfquDp+kr
9CUNw00KIWEstJZh+0JEPjGiDoSKDLCuVipE6K0lLIAPhBrhAYCsGHQB15Iz0CVa
MpfxpvicR216midA17Y48BElzYAiFNOlstZ09a6U0RfOpOx5DVyXOqwc0a4ccQxd
Je/YcObq8WJlkAXFTOEqXgfVTZb+Eg61ovZL8S1kibMdDtjI6tBGeQpDg+CK8NZp
9UkoG1V49Mkqr603e4x68UcQJxCdFeN0hL3jYHCV88iokIUln49xhAEdKxt3eFr1
j4yySzwKyz/EXzja5bXhAO4bssRtqngRf7mXh8eZdmWEGJ0Ak/OoTBci6XFWx45y
yUXSm+HQW7VVK+NsDSTZvp+PIJWIfODOfWr+kuopfVPJujkOJjS2sPpFeDQVFNvt
qfcjP5kOXbPdtcgs2dAKryRIumZPmeXXtUF5pcE3Cy6koXeSBh3euoYInRucXPmf
oDs1BHlNxRQAy2XSssSXsNy2yAd/X1w9rbt1SK3zvqPsN5qvdEM9nUCVAmVLDBtd
8hPRaJIuyMKLhFMGtKNvQG18ftuL08ONg+aqyrHVhWNeFhVZxE2NS5T9tSUPueb8
7zHiG0AMyT+896D7XrOrU135nBuJpZeZFLXT8HcvjDgNGPN0ZBd/dThIBjkws1k4
kQl8rpm5Bo80z3FAHynQ70ZZ7j+k+k+PUMW+IKqroAqtjdVrnQepRCYPAEIQNoiD
1WLqfZiAEvF7IB7Pl1BV5H937QVRSXkGeFCCwHxlrTquH/T8qCbTH9xp0HYhi17i
2d+XO8wJ4pTlV3NU1AcpIJPg3fKMAyF/VQLya0TRzkNEhrDCpzxGg2cJhcV0eek4
4fkz7D+hyT7Z2LQulnqXl9BqqTjtEbWbqI+W9oBHJvDGrdKVvvy53J1F9RhlE5HD
h7xJ/wGGuGHcfQvV0tzotEjVk/52+Wk3TsYmItEK5U3/8vRSEOK3LfzF23+iDw0Z
7C9xI9Rv1s4aSwPI5aZybDNlEsWrBpUnygnZIcxNMOuS3O17FV8wkOrwhlVUiMG5
W7WYxymH0R+UVTEgOjA4MLknhwDeyfMQ+XH1ftl3VFMDAJOVzsybOLm7B8cKn5XB
Nhy56w9Z6zCJf2lkMTeOjooD9fwkrNcvjIOlFVhOHA2Gt89b+ACmZ966js2+JJJ8
OZ6ci9isym/HPh51C4UgMWlkOg/WKiGM5+OcuqHHGtCu/KBThpLFfMKya8lVtBwo
SYPFcu2xcMfEaEMB7nfQjjvYwvOdbSNhF7xhBeb1tpGO4z0xZFvPAC9786ky48N6
i4v+8PLXTNSqR88kLRFX0WnVsC1NWOGHPp9UKARtkLphkV8JiebHls3T6iCn+g2Z
4HJHAOClzmX1Pw0dyBaZcJ/JOHqdnewdK4P2Ma18wBNc6AsAaD62NMXNRhBSw2dd
LZRNz1c1JztBstYLnSS+Ro2s+qjeTHsnMXeJ6L2jq8sMRP0ibqLyQ+d3c63rPhHE
8gRKhpt4iU/E+vC7liESCSMg/00RobRCyR16shVEMkdgVBF5PstgNPNjJbac/duL
Y7xPv5egxah4KwIZ/sfkfxMDXIKyrAAgek0Pz+kWuld64PR9ZTB5wJXBSswaV4jf
5IL0k73+ouNdAlJR12JDElRMVvCmI8nSBXWHDSN+ToHGKH+ruNzE1p0w4W/PHBhK
5jIiFdYWdDQnd5cjqZoixWSAWLOa0gFCdM2Xkevluqkd+3iYP7+cLDx16U9DVFTW
GMvzhb5D1ChRgpMpEsuq0Nnpb66Yiw4n76d+VLoUvEQGt1pMnXT2eKUXMg/NLEPn
LH14v8a0uJCIzycj2Wiqdwo+fJhmgAki6bn8wyStAJgel/NjwCgiy+GbiNF+5u09
7zw7zPnNBef0m/RRq1hmA22tpNgqknJw1uSdc9p7tk0WVZsG5I4357NUa2K64xRa
ro/9Y/thFRX7k0oSKipaw+3f8EEHBMYwaGbSjMK9hS0YMLG9YwYwkfZ4VIYMzUO1
UoWfCYIgVKm5iq4Gs02f7AN0u7cVpjxJ31lQH79pLYEz3tZhOZmQlff3IJzBitPo
4gFUtjHqi1r04s9BCASoE8pixjpgJ05uQBxMjgPOtWLLegyOr+Md8WU/T+FRgSuJ
x+5iRvIcJNdh7xDh6lTc3imx1vDyFlZZO93A4bKinFGa0u1dZ7Z3xJdCCKCP0v+8
+Bu5v+tlki+0kOBWxZRUTHy9ImfRgEKx0xYpjfBlSm9GVsf3qb2wIip9V8E8zCBl
ZTE3smaMCRtfj7Wabz5k8eVMrf/tMWG3ryI/EKvuy+BMtUNtQPeo29h7K/q1dkSc
q003Dv/dapgcB8w/Bp4posx/WQD9Z6OeDwN4MNnr5dJ6oexeGtXdNYVzuoTCxEKq
UU85nIe68tREINRDqQzRNQwuUyLzL+21/X2QNALqbdMoQUwNXhkNyjU8FJS5kw8V
YdCfMGNJEzRhpTmO48NjvEphqZiQ7ko7dCnBXEL8ucRu8LH47az+OW8piocKoU6I
VFdy2LaICLOmmCrRdeVXwDusD+UWIe4NcrGfyCBWVz3ztNsItKtHSvwpyXrm5+un
k+bJ0LGnuqymDTQPe3wsx1c+bhqRFoVwUz78XZIMPj0sUz/Ib6M77fUo7tJNKLMD
RrnoE7Kah8hhA/DmjAxVe7GzpLmYokrdz7O18RhrfbWHpBE5y+zjFRF/lVrAN2dH
IFioPKwMsERZQO4cfQCJwDbPF6dDrXsCqgfjuJvSJ2mJqrsUD0p9zW37U7WpJVB7
o7mMbjOS/V2f8FN498N2BA==
`protect END_PROTECTED
