`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
94CcMWHY91iBF3pOXpIgqo5ZblQotTiBFINo6XNBVAzeEA1i/1d1/vyV5YKx1ojZ
kpmOHBXZD7Vh4xUZuZ41wiYmCHeFl7E/r683JfxmgDnvRbGDj5M5HF5Sg1q57Xlt
uhNWf3EGv9jFfazvic3SD08Ew/PsQNZ6TYBLm1qmbFgK4zrtKHLg+3tWejk94Bsk
kKn4Tnlkp2rfxu0FEg+gkEKAR+zC0q6ZuPZGbsa66TpwjuWWv7PxS9dGyJ/ina5o
aezf/xtl+IvZqI+V08bYjAgMJ6hDF7RIKejJbA00O4QcEx9r7pE5qZ4RzQu3BPai
qjAO3saSjRA1DOudviIy0G+wM2CUX52jyWLqFecAczk4GXKHCiobML50AZTHyDNp
mMx+hHV8ozPNC6SSd3sL/g7eibk9FylW+4ItQVml7aSz0dHXSrMk+9VBuS1s9mUu
xNE8ezRVYA/gLqYAeKSeoLsBHFa4oLfKwN3nlv+KrF/2ht61DKe+46XYVndW8NF2
gjOxhCIQLl4DOq6AwVMapblaWfTHfpUolygkcy4QMFL/yfQklxUSnesREIQOjKqi
ljojCEM4F4Dtq4jgy2YXgRCbjcc7qxEP3nFh/yiamY0qVO5BBRj4PO+UMh7tnT/w
3aQkK9Jh5CRXT8/dspivHvfGxKk6CeH/9/kx7sX0pcl4o6vvFJbq5YEOJvn/ozHl
B5iUesqWTZGQvzhS4qIlJ1Ccjqu81MFk90RPKSa9/P4wGkiXhv/ozDg/fi2n74ZI
HNitPS7vB9W5xJn3anj3GmR+MO1LI3VacQEOZIOQIo46qquGiRM0+IDCV5DwZDl1
xXpz64QB187t+HfXx0bRHVwz+i1cnm3fMujrsr/Nj0M9KaaBmJl/iq09Wx/1xFXJ
4SEdQAdqOtapgq2WvLYWdmqJU3GIR5xKbmMSNx3s7V31zlsBikMZbSZi9VGhPOeH
JBwbcCJKlQ4yBDcqtUSxQdeMGTttKI0Uk0wa/kO3PsfnR8tp4mXnT5WeTg26Ycjb
`protect END_PROTECTED
