`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OYA07GbdiTDwHClYHwjxXXNQtGPKxnJ2yYmMvcTOTXyRbIc4KhTHMdFyiyTcljEs
o/dsduL633d3dXr3KcpdvVOdjs51WYyQkfBQgrbf30YAwBcuuImlvwqs/qUOAPUd
sPFBO2NYfDD9nezzibCbEjVs05SQrV+GUGHiCXXmje3pYWh+9thJ4cI0dqP6DkrE
cJz8y7QwgVpDAhM46cfd3qXyjkuhtpoeWa+T+OztgU/6B9qayEtGQ3z9R3REHgFo
T2Hb1tVsqkWFQW8EBK6AIWq3Q27/jMELkkciwleJ/lY7vmM3eztcLh9VDkd0XR/l
gfIbC7Uzw6hzbcZylAY4uSFf6Hdu2hRpIB3vThgMKUF+M7xzLAbBB5+3wEiGEvUB
zuIZQq6egEqyeCKcDjR2GpqHoReVPUSDJplpksvHitGt+BarIW18EMBlcMpO54+F
75UDRajx+xUiAmkYFcn1CEndQgvld29vslSK8M5dJ3YYsorkCzMqWSkT6whCYRMi
yYvFjXXR5h+FcLNWaCzipF4jMShfOj7Ho9hwk5DMkv385WpTe2G5BhILaghTijP8
pV9zpKpU3hWRci71wnYcE3DEP4q/nEMNaj6MBFzbzPb6f0IbYpFogaEo4bLtJeTu
`protect END_PROTECTED
