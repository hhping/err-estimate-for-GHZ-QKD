`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W8xjORzWQ0Qmf399G94V572d64Nr41GMMYJqoDlt9WWqBcEEAYR6YU6k8iIE2AMd
ZXMMwUhioK69IDuA3RGpz8NXAheEZD1Cz0NcXWoYk8/SlZCZntRhix8hZ/EcQa3P
sMpMN0OXAN5Z5n+LSU0VHPOduu4//NKzdwYEnl1oT+tw9aOvr0oOYiEbU6AOp2Gq
eKhd/RSA6bzkKrkkhhCgzOHsIcRnrss962H66OA86kzgqB98nsdns2AEuOTWgG2i
ZrMrSRbjYscVAWcW9dhWBeXSjofbsF7hOyvRr423dfjE8HK4RGl78nisGpwLPpx8
5vPrtB24e794tLxh7BJOSt+loxl0PmjngUfyVss/E/QgonKx33H1GZ72HWFphZew
JVrJuQfrp7Whd1JuDIGrsaILJWvcQv9uwRbiRXRpOwUjR2R/D0FFwZZaRd1Wql3O
U7OqrNCCpU2vQ4Fxct14VCbYkTqJE+Y0ARon8iSVPmC282Tl3XVBAXLS/jkouhv4
wPDbEVFMvlqta+aAqRpsCyLJ6vC73dCeNDutbhnOAKC5ey0gctqAFWb3sfQRh+qN
yJkKmOcaajvICh6h/xE1y+UoerB8HWQB4XPdOAqZbET3xPmbfqxUWybNvWGW19RR
qBqGn2y3UF86vstwmKCa0e26zOMBuKv1kTCZN0uKiAKtIgBmuUuyYSrCIbGjhpvd
M6b7mQC7MIlk/vdedIN3JmmGTbWV/cDPQA2nXDcRhBDraj2IlCSs0hdprens6B1P
tm9pQsgrmWY5sueeSAkUfPKMDuNxs2QrZUVyuCuvab8+05xAgroyXAdzQtWwbhd8
lBUqw3MvlHlsJvXaP++mPNvgMA6p5XFsFWtPYsDVCZDbe8U5xEjQOFaSvjHlkLpb
QLpuIFbLDlXVU8o82xLbHlELCoPX1w+oLp2i8Gzl/U2vInlYEehlwF8lqFXnBiI9
h+wjlTt86aO0mOZhKFCSM6/s4qbzhVW9p1RPvIYcP5JmJOeC3fVjZoo9uH1O1r3z
wzFREEiwd6+PfNjwY6UiNmpUxd8NzrbiQOOZJdRP7lrBLez9xnAS32lcl/I7zG89
haJLWOH6B7/ItnVPMYBQ55Jx16SuXTzTE9X2MkzFy03FHu7bQP5owUZZ+vWkT1/2
UqC/yYCPoVkA8ekRI9AlgLcc1iSybh3aLN3InUl2021X+GE6klsJh+XGmg1UaYEZ
ed5V6+GI3aIfnYREi1gvlObDhCWUijLourox9/VzI3ztuxuBAF/wEZxxCqOz6ADJ
+7Pn2soX5CBltD5CfRmfKlkTORCpHPT7q1BVun7pedvZT6gWNDzWQTImjdhWSe6o
6Mc676Ig4FOAbd1o+LqXE+iET7y9vcYyMGkTT+P9WISu+TWP8NfQmAPLL6lAQAII
/WOmtgWNZI2JsHMmon8iwP157XKcJUlBibDT3UMCc/ssYhuaQFhWxFkW7sTAHKT1
a0CBp7KC6Hp7tpaGd3yZBmKr0PMTjpw7MVUy92R5guMvsgbdTV5FFFUTLlfkvp3t
rvFRzdNSeDyeu/ZygfJ0LG9fklxwiOeYPg/ai+fj6tWTU9mlXJ/thhxPCY9JdIm5
qwM5sL9bOnqnAZEanLbFllLGIHiWxjrCwarisOlUOo9evDBqOqyEOPIGFS2hC5H6
qgUtLEoueyEBLgvK6x+rB2C/HvJ597+AMjPSlug0VNlMqkMtK6v+mNUr3dWyKjO/
U8LCm/qgRAHRDM8m0jtkR55YHkRgu8MvXb2tsVlfGe1cJQtcmqxbsWi5rZ0unKi1
JJjB2VzSPnX9tp0L070DfcnLn+WIqvnErmWzmlH4YQ1b0gCEqwb8KEG6TxSlH/rI
UEKJ5ZjGkD36mIQYoe4ERln6hK5VJiDL4wUlggoZv7+uAUqBrZvilzMZWQ2B2dgs
rwgRbg+cDFNAx3lS04fA7z2rTMtO6BsQROKuYyjIvutHBboXa1HDgEt0mSa1X7GC
nmOZYNVvTgNgItHy3N5qL3kWvLMXDwVHYXyPZrJ5lv8/uj9KN+TWuBXy/KYgs+cv
laBvR8e1sAGGWh90WKbR00sGeBSthRWLKdvbEAFTFy5pgHoRmKZcaUjyuLojsXsv
NU+/v6Yqxbif4NNodBtoftOnom2Lu6Oq06rxJXZfZzA497hhD9OKSuV0fXu3tglM
N5LaqFB+SThFHpr9fJ6o3j89a79bKb+bLWVAIrq8F6uzH2j8DR62BkU7BBdX79aJ
19ddh8HlEO7p1/AF8T79tirEFrl7gXPp02PvBFXLIDKqvpZB4WqMtucKgpDKlWyY
DdNiED3AMtS4GnIgahfpJnZuI2VGbFDG82V4FcweGDe8WUIJzALqVLU8T0fPTtuy
3mKEliCMZuuqYI5f7/5V+rQpTJ7tVhwTVM461a2EsGxfSeYwbOfPlNWVaPR1AIoa
u8cMlortb4y5vBqh5n3MuZrmEshSg4kyoMQZeY8xLg5ealOLmS/OeqystV2NffuH
hY8QdVF49YNJyazySXnSEgsIluAegm6KTwJh9qefvJc3jSEwvXMpYgaROM0dKjOq
+lQbrUL0ivR7auZ8yD5pV0vCpMIFbHO/l2heOZca7mssPPA70u9EFghm/ZleoQ3+
RlrlihQ9+iT6vqqZA9cBKhHo5ZaR4vr35BAS88EaRUID60XM7Gf99uo8DguE8AEb
4rR+fjdFKDqp+7IVoQ04vYsSkz7fzAaWxZNHkugKwtcY1RQLwsN1lUBlI/3GEpf0
o/6oWwCh4WBDEYMeTHeXCiqOt75e/ee+UZFtpe2ojHTz2XuHmNbT6m4eLvbFkyIz
mmMTLjJ1jyj6X6q+n7/gNOLSrcwfmpBZzd47lDbOYX8wIEl+hRriTk/bkry2udmV
xm4KfIY3Zrd3Ydk5Yhc8uNSz2bd8UuHm15tiNQkY5Ldl17CNCMZnOwkJ2HVhX2sM
NhjldIqloPwz4KViiYSedw1uXIym7dBJtZb9yyjuwS2ifXQm42tWY42faaZLeFh3
kXl0NB8PtL8nCCqpFqc4O/xqzckb8y+k/vmURpQTXQEXT1x0iA7ownMFfM8HzHO8
JUzfgypOytxHoZ16PuqOIWNrNDaYle2NtE1NwXa44mwwjIb3BvmD9m6BlCg6uJks
L995Ej9ePZMloN/8cGqmr3smxVR9AuFFCts3T56psN9SsguO9tuQqhPxpI1SZAiI
bwQe5JR1qPqazV4Q4O6fyxDFpu0e7+lwLarw8hYMabLZVMY+V20r5x4zH7/yw9E5
UxSDp7Rb31dnH+9lmnYqzAI2Ew6bfZLVsjBUHOt6bYdcVcWlkD95Y5Y4PQ9Sw1jd
JOSrC+ZK70yQNTS/c2KMK9B5nYgF5sHbEyTxnJo7n6gSNhsMu9JCXv7MUGtYEjvN
UD4qCFPVsVrAxuPEb7cTTtxGa15VY/bAg4bzRkAfX918UCrYTiL2lRlBONej3BSU
WuKHaWaEdR8e40xjPw3zuWDoJDyaeS/y44cnKUhaPxMsqIFZR+/tVDAOZhrpYEMN
PwAZ/lOlvNi9l+2D9wXHOtsXR/sJxQL2Su53PF+eycKaHusSxDsF+zk+JS73kdVg
gQyel7k49HHosuhD8r0nIYYnv3vqk4afm4b1kZOeFJ+4EOUm3fi3FTiBKFhMwRAd
xPPCBKkpbZ8DxSzewW5IYH9QQCnOvQUdjIRIOuKhCOnjkeGuSuvfLvSml5QEyNlD
B3ZtKMT/Dy69VzfCPvjKKLh8CPYyOwKMaV92eNUKFYdeGyr2vhL5pbLXXWbW+ZcE
jJVgCApTAhq7jJg2wBJvnbhV98/nfPH7+o/BgPIr7Iepi5oN6/l9MxpRROd7bV7q
TgmKdk9QdjaSFoxzw6AIYUxsc4wiR4H9nnmnY9wssHXNCyuXx0hlP1GHq7lrGAq4
ebhEbuu73MPK/OPIlVbr6sh4EymZmCZfbTKn9rZ9jLW31HFEspv4Oe1NqSVwDQiw
SE0S90xwiL41i5nYz+ExA/9HolSki0Qq7L+3sXVdHFy/WDBa1a05ONOXUGp9zGr7
pZAMnSDLNEQGfu9cXiTWexb7S6ubDQ4NEVR5D+7mZRcDObyOy7z2OBvaJJZzOp6h
H1ryh+s6k8UGU3jQnOlZpCZgK2WUYk0p6GQeIurONzCQ37CPWiElfZ1TZcT+ST6P
gTy1/sc9j3wXzm4kl+XLYH6VpXqAZZ8KW277uEe9yXQWTtOwzg89Qv2l2Jr5HS6a
iSDPmbl2Z5eXi64Lm2CAotq1vofMXyWlLNMklHpDF+NbIeaw8p5w9a4LrKoAKqiU
eagex5Q8mGG64ka9mrRV+X/PZJFUVm8wa90OFrI3aNya+Y4rekyVIBFj1CDFjd/Z
alVKj3tXQkKgLfwAR53TKpWnNvryO7d1ive+Fs9dxJORwva7Miv5M3X6/Vb2E3Bo
Se+Q07j6qeehYBNenEsmq2/rE7ttns8Jwu5ELUqCLcX2DsfTd44ZLw5PA4gKeWVx
TzTq6SFVGHYg4RJpohDnpPsuUCYhU0ZD4N0zbOTZoQ2xhHhxKSQjpFsZKIvD9Qmd
7cHa9cmjXTJjn0niRIrTabnxXZ1IXaF22RNK6xyMh7hQ667FPQ828+u0FNrz4RCP
c4zo7wo7unHifEnG1OfSreo2HS1kU9Vu7zrMjx2CqbKKBXV5ryzkFX4G4sFiwehg
0YCElBPYcw/RLneQCemr+ac89l3B2eNPAEATzSTyCQ6I4X/aZYS3IHEEPTaaYmKZ
WpabaljBfYHHozLA76aR1IN6a1/UikZ4bwHgbLx9ZS+v8jAgTcP+W2MKzKkceXbC
rjxZrlKmRt032SWtm/ZxTJ1a/NE0Xbs2WRSbmu+R23+XlUMvriVJ2ULqi7KpU4fu
K94u49Iqugx74tHs7wxp7C260Tp8ok5q81m16vmrU+s9p4SWdFW9Z7x/pDa0p9a8
cP4bJLbSKDDfM8GdFWP7B7EBiGokNGur+jlBZBcclFzJwHAaIAlxjNeFcbW0MZjZ
1JcuxX2t7DyWvzx+jbuz7AqOt9iZPJ97Thrn+tRFr1u+KI2mNTYkOI0XTE+vkJTI
sqOTJp79k/4um+rXxNcskNveqtycNY2QPbAbW7raVcliNqqTG9/T/hq3JEvCIFAA
f0+0vHX62DfEy1gH7HGfaeJAJ77NU3NK1WXebw/7d9np6jQ02LLXBYWUuG9vRt2e
zd/vyZ3mNaXS3ZLpwfVL+lkoaWanykmsD6djVdnyvif4jXcBCZcVmSth4QcskO1t
+QE+ovI/5LEvhzIRycVGLZ3yzYjPq69FAlxq6ukkAETkSqWYuEjN7N32C/u8K7US
v7sQbCrJSo9hZ5+Im0oaEMiS2eLzqByEfQtM0K/28PbI5wegOYsACJQD4JDWNpRL
cEp51YZcpQI+765IVSswwcYt3NgjUureGJGDD1WZniuacPgFZ44ejZJHi8Y/VK+5
+jvGptIP1WxQvil1QEIZOk5Dh/WIsXxGqYGJ8khpuBwwZltgT+n0MVYmef1FCetM
yl+yAViWnwH+bIN61wlzjNpuLVMzX49/UaDqnQh/LM5Wj8tNetC5Yvh9g13g7Xa6
ycSMmz8AOpMCKpgiBMiKkcjVQjtt5GzM1alCkKlVrwPFgmkQARDwhdL+A0R+OTQK
TMqJac02RRgNDR9Z0vGu3c+0h47DBkFF2wvgMzWLd6QCukDKYIA0ylYBgL2+zlpj
2EIHaUHpadeopSJ57H5o78A32he894IKW5ei2S29DbP9AMrmnmvw4mbnsxg57i5r
35/R/IdhQgBqdWWwDEbFFY03hhN4cQfxRCxvL97tyoQCg4/vPf2gIQQfNog1PUMV
J/dV15cLCq8NO2haHTMyC8yXhtnZE7CrAg5pOCzDAKTRsy29CnixeYl68QWKlyhu
G5ry08VmMoCSqQ0sLy3owN2MKE5f13INvy5RpJLFJPqOtrm/smlHvMnEpoGTyIbZ
KRHEedzIo0UnQ33qmaMagXjgivL+wzeZK7N/OZssiY+L1vV/F7du3vr9n2lU7Nc5
fdWC5NJypVTzRmwHl7Rndy2+wY/PCjANCDcSGJBV+bidoeQHY0oqtE5Sik+tqVRm
rGfApELax69So13Og4EVRZCpBokdUZwkGUHOJqrBG7UFXL+91IimZdj2xy89yZ4r
/4576P/jVJYKtzqnS7xpOoh33x2+nst8i4ip00HRrRY+mG/FgRA3KWevmzCm20YN
HmLeVjjiF0BH10eAxxXRsGeC5Le2NwdBVDzWvQjxMUv7ji0XmEWyd/mH3X8+F1RN
go2EthSll17Fid9uOS4eoxByX74EYKGYIiDMxOVqDYkbgFyOxcPpSdckrcHrLvzv
GCjNpIMiADRchXtak90Rflj3C7xhuXmEGb94E379DKC3MK66l30wxZ2zw0Ja9lsK
0tvvd8DV6r7ABsGkYe0t23LP37IvlVxYfErq9QOvBTn4rdcRhem3eoy1mNkqUaVP
FKhaLwVsaTaklliAyJ4Nbv6HbzFSsvdclKJvzu3cZM/SwhuAhADG8DA+3irYBYTo
iACFK/aLz5Y+2qrELwAyfCnqGws0njMYLw0JotbhxHSmqsEm3/EdoSfM7EBtIeGg
zQASYW2BGoZWqO9EvGoY9fcEZ3ehHIloiR49DeNr9HFr/uQeuYNuyOEK+fOCEHvp
zQah8t0M9lrYWWOtATaDp7MoNSVUg0k3YCzXzCosDcbvmxhtThKYGL7+EoeX3J6+
rCeE/nbxdhhCBVSkWzN7UoQnFPN638kb80ZYI6MimjG0UuxSFZzap1H8DFPfSIqc
O4uLcseX9uCuGXNxzj/8gRRwTHwf63a8pIJOSJ+NqNWSeJqTr9LpfjhQWeV+PJLw
h4UT+NMy0Igv6idFmeBsPk/tGh9K4qDIBKU+5+6bvUWbWnsWHPT1Zdm+jw5H91xA
GpyKdI0J1b85WqzKndQoGbe0yS/VCWdX0QPv/nt/2srKCZsFfEkXzXaEFYXIlELg
rW8KLEVdaKVbhRzE++QpCsL2P2NN8xYdipqhiR8IX1x0Mspcb6LgmmiUQGtGZp3u
HovG5mh6ExrH9FnvsIquA1aK3FSVAykEUJT3l9c0NUQFUWztwr+m6ufHlkmQMNws
R1ZDUT+eUj8nKbJvxPbkSU8hAfr18+f3uNusAU2U0JoNO+xjKHDzC+R6fXsW+EU+
9is/EJkgm93rhhIdyWhjZOz0akZDYywUoho1GxB1UkLuy7MKK8Zm+VsfHGw7t5we
cXWnJUJrHw5JtwWg1w6SaunX/4/sUgpc8WA61EcFjQuVAXuYFPNoRZjgU6xHDmSW
NizipFRkfmfR8N8ECAdWaoWRQ/YOt6Z6p5UN+mL8DuiVpBJmmXhzTuglB7GWHQZf
MtN5OX2UiNVRTFIxC0zPRnD0k8XjkFaMJgC9srkxQJ8oe5Ui4kjx94UTlg3rmLPC
XfF5tT6GnXuuj3HgOM3NdntozIZ1+FpQWnY4QXqPq7bn72QkNpsd5U/oLoJbIe8C
WP2IOadqxiRklLxLgRAXZM+iOPaSJsTDH4lcZ4alWLb1yuNkohgtF3kqbkGXkyC+
Ahn81X07iFwOrFjhgVWI+K1AvNkz/Tqd4Ho2mStS6dGdZV/PCu1R+4skhkucTfnE
/2MiaN7/QTMxTaLrZcxPrNVF2gS5UHSd71mXExw0GUTMqLwO2u4QO7cpS+kfGEz0
FWxF/l1eswS0jqOZu8nwPsC4426fAmXq0LUghEphwY0Wy+G3gBuBEHroPq1hHPFC
LcpWgm8ZN/kH0qmnIT6zcHJ/Os8pFE0yzF3Cc2wGiR9xeG3+ngPnzuByxpCTWU6Z
E4OAabhDeZqJPfZrTRFyTIBnUwtrEAu3kko+XpNPQmM4F0jhP74G93e9QvqEGdqC
j0G1wXN06Dvob5ck9xHGabnNUlTZs6kUG2LWBi9ZNC90PkstCuuXCjaA/Txw+IK+
BrV8il8UiZMueJ+6xn0PH27RnROCXL6X2u2YhWvKVBAgmRzpuID/Gek3EyBGgDqt
yzzYqjBenFsM7z7aPex8yL7QSVRF19srGavb8alDlp0TacyaJMr1XO6OwJrUyRKe
g12BjNyq/t1NynT9DVO1L/soRfnhnOXyyxcnM7I5guo2eUN4aFI62xGkPQ0LYL15
psbpJbeEW/Z71qyPRRyr0R9vJMCtWaWYpDzHti6JlfVkuuht1x8U+oKZIaB278kw
YkV/CdFU3LFSpUr5YZtUQJ0GxJ3wcLqRTlYH0SUI2yqbiHpdw9Dj2EiOZKVi+2jS
7pGig1cOjZG+vBqdhuzlJNOo1VHWtgXExns6gIHYsvy77EwrCRZEBxSG6mf+mgkF
ifqgAiIb6J8/6tikGDl1evrIZq0Uqzl0kg3LrZxqTpSU7X3CW5J6gfP84HvrtaQk
tm3Tw2CPiEC1bWLt5I3fM60OH4WHCGCj0HAlcxNPP76zYKsNAvwtI7QaxZglWwFf
z+n0hrOAVSuzRfdqmafy8YgnulbK3/0idKTui2m2UDhngef0Qc6lbtA+umjMXfl8
1F78z3AuhcyCJlrlHSBvPm/GGN1ePUDFDjm+gBflhVFqPmVb0iEbBxmTS5oOEu/F
swKb/LQbaW9dP5ckATQpk/SYGsmSKEa36n3TbZmNpZWe3QxMhGNuyXIPzvI7MYGS
KgkMI5/GLX1tiodFwOyh0YfFFZlwhm0Tzf8dSeXfe0ikM06apppbTPe96BmA6/2v
vcqcaXfzgP7+t9p8LES3L8eFODkjo7miPIIew8wxuMQHW8RJdf7noeE0atEJdrJL
dSo/iYE7OU238OpmDC1l/uRCc+9+9tpPlzAB+W7y54XShQz0XqsQjLHyr1qrkFYH
LsF6J5Whm4gQQar1aVZYSDZBOdkzW9jZW+QpxxuB2p0PSg/a3jbX8xedB5dxgNkJ
s5zPvPftciWb7L3EIvhQTevoKee4UmxMzFVc8qVLzat/RVcNztzQ7mdAEcYuquLg
PeTn8IDFMl/ulqriWigrjo6uaxOIJY1dLe3zdZl8sLj1xWbIOESAEnybW7+6OGti
27xWGgLLv4GCqaZsXwD4Fj3YqEFY134qGPlbR+3pVlsPnmbr3RMDspDa1rVb4/3C
jJce6YQqUryowkxY9LxT1Tl9mBc/jLXZl/qGHCGStlWS7qgkivNPPXWUmkEEjUlt
+X3khwE991lXLWYx59gYiNp+efvyKK0mZcHp8FQQSrMAWgioS9nzNVv3CYggGXJa
SfYb8EtD7QGZQHWLyqB4uhrH3fZ6TF0KqLm7RgAeSt3REoV5w6lqRmy4hoxBrevB
nAEblXn9Ws3hkWVFQsQyx8uY3eF78+90zHIqBkDeemkCtxFz8f2K5PUHEM5kK3E7
P4YNFYFik5te4OKsnWmLTaxVy4VcBrIJpn4Ci8sQQkOlHx4C1rUB4x8hKDQ7siVS
ZCxr79+txYTEmAThSm/eqYDfB1Dyg0cF2zYZJ+GEGD2aVoED2BMShPCfyh/dDnoQ
0TkjgM6omUEq9KR3I1iJr2VMT9VIqzhcxSqTZD+gff+8/Ti+IPrhSJ/RwwDpWUIB
1SbWwCpWvpg9DOI6j+Jk8JSSHb45xpv0I8GamtoEX9G2FS7BTA9OlSECDudqY8Ea
lmgKLrk4rYThSrvA0pMHB5q/sjTcn1eAB+uP3NOn7SiRGHzZGkseSpEU78R53DDg
LKzSDTmdTciDeae21e9Tutuy8Bb1q3dkFEez8QIiZK1opYzYpuSRRctz7JVvJozY
u5iZvbM/L5Z5Cy8cvDeRaFz3Nh3ViC1GF4TLrZmbXV08BWap2BnXI4eaCrWCdULU
ssI6irIRboFtkC0z3nYiHZmrvmuIGFSHmMtcg7dTah5DGlJSdYS5pt5HbgPSk1+X
grYPp8m9d8DzkRGU6tpaGR6hf2d9bDIrJTY88FTuNgjWjkFXEluew1Pkp1MUReaF
mfuwbVV00S2HKXcOstXskX44rkHPhCJUNKCqLgK2RgNEW93hzWoMu+ghgu1FkCPN
/S5QaxfVcEkvDijbepFRH5cqRLUItWMEndGvIi2aIJt+Gf/QXzA3NY6YK5cufZuB
clYuvzH1fZmu+M88rK/mOh9+S5jL43WqQDfv4CGR+hkss+j5MWcGH3aI0bKJTtA/
4GRMTkaXbpl1KPfkLiyMdY/Qv7FLYJ9cp+fY91ZQlJuX8r4e5ObFwVP7Cp6Pndjq
NLyjrkNhH4UO6+xC9ln3BhKZ2bYvfPlTXbzR8n9VI3Cl33m30GBw8Rg7nifNPOPA
BzERxCd8IVgLWIBn8i5K5XVJLLVW8nXwpUcllQC3AtUw0cDy0zkML3x5JGzAoZ5/
YZB5XLLHdsk8j8fPo0cikpkCmqZKutIlw7SmqMhMfxZ6MkN//mhotFfGZ85dbZqx
P82oAw4wVYPTYOrWZ5xzilZ11noa6zHeqTJ0Aimo+QOryyt/Oc2Lf7Hpn4z5BSsN
e4tUyveyFMB74ef89zVaeIEBHSF03iz4urX1DzuxkffuMmiQja2bmt2L3Q4y06fc
2IS4UUcL8Mruy3SbCZrOYfT6pNMJMFPSHL/Msw0+L03vTi876rNn0Yro8DHHE8Bw
WZ/cB6mXzgEOTqd3ZPP7rOMSXmiQ4lcT3weysU0SPM7F1wcA/twgmlyNHXGff08/
VUivn8rkwuPGSNgMcFnYlrJo+wQmIi524OwvqcAJ3XXGestWXbaZIq7zH7+oH57j
3jg3tOcBysNuHX1agY1X6SdjYj9XrrQGFGBY1jgI/QrccC2H4PkzX3JS8DaK9DJR
PPxoLQum+V7O103ZpwxtXJNRvFvruxA3M8k9v+IQgLKp+B6DrXTmSJyc5VIHza2I
YXLcnWKcG7nXZb5dFd+U/3m5vuz7TWJq/cSB4KT4UL8M/Zqd4lqckv+3FGwKV2fu
6WryhIvkHpj6I8yNfPhDJETOSmQC30RiXRv6dYZ+1klcKhwmeMXFosIlRbdtlIJj
ueSOI3BdF5cG3jMl+Ch0/n5DPuQ8fOCcoGViHeHWR0hwfTs3JS8AMENhH9DJLhMj
oLP3VME4xC5iy9Qvx5aW5nW92GRPQMFKa+Bib5RxUhhYLenZtnlUdsPNQsc/lBNf
tQSE3eL2D6R/c9z/KTVqco5mhEWcM23xsCoFLWb8tmIffMa3M9oayptoZecgtoQ6
GW1F8BKuwjPANg06DxNGHT2azHgKCGW02E0lMLqhGlNBlt4LvoB0D+l+n01GNBdW
aUPu7nC6h/ioUkqKv5FQGNCYweKQnsxlr3vzGT0tmuKFEMz3J3w9+vT+MLwpfvqB
93lrf6QQItc1DpxghZfK8DIZRf8IUepTLbQwmfUdYBfA71WA6Id6Jz+MgG+XEEJY
gWra9BG4jpMv2jKNSySZgTkQpl64fxdSSO4Mqae07KT21gtt3wbFQcMzcNAo2sc8
Cau9AmixL1/6Shj6YnQ4Ir4jbaG/EFrJ5DC0w5/pSPXqaE3AYnlqx65PC+U8jikt
rGiZEis0O60G3bIolMxFnjBVpQIeJYNYWc7lIQdaY2NXH4Ry+clPJxmH276IfHQk
L1AnDQxCh6/4bSOE778MGXydAPaS/5XQJA5GP+lOGvQLWwd5h8ACuZ5BmhD0Yfap
mGySzMHONhNMi0J1ORCO9cJO+LSKSROpppaGzZc0Y5VFERjwk0B1E4e7yh19OeqM
liyTi8yAs5FfR9Z1T2jDe0FxoPdA/1z57vweNNaKIMXUDpmiiF8g72H1ShgyzUXG
VuqEK4TuRU98OxXDB/dnvc+QOUIexlgRW+afQknSksg5G1lTzEi1I1FBQ25OqiOT
5KbsumbqxOemYvJoZru6URk3GHoykCFlH4QLUVYl0MjW7upYjf5wMz0iFry9ToX7
r6fkRcXEO1A+8e4r1pyBb2AJb9tsiZMBJ8H39op7uaFgKb6VDHQ+e+lsEo39gvF6
XyteIeqa4DaSyuvfMzlbicz03HyFpMdCHnWQ9VH3FydsSlZsYFWEK3dp6xO6AiC1
l+h+WfzU8aj8TGAXy9T0K4IQNL0VphUWBRR/gtn2YUmnjo/ld9ExdaC/nN4tiwjS
E21BIviSjV5qwKmpziWXgPgLeWp5qi2CW+WMBhWJ7kY9/n1SNZzU95EfdBmnfbdT
7RT2rKVbB+0Bdi+R6Pik4DEI7VJ4TMCzrzKAdQ88p4aNmUTKtAvSBOVeLWb570E3
M46mg9icT4aqnXs7DEwaSLNNaskJIiMM2E7BSU5fgTvaOXwcMQghN3biF8lp3CXq
BBZGmGTZHmZjJVq6Uo8bvkde/2YN8UD/miF/dz3U9jKwwKi/CchBcImGLLPduQEi
KlvVyKySVGS5faXcs6ryWgTV4jm1fE+Z/6aEsgwIlzLLGIaIlzFhU4cIjhyE7qGf
B++AfrsqvT2AaK/KgG4rzmBqdspJzdM3BG1yx14YiPkwQjgRh7x2kh3WWac/gGU0
QSY2P5R6I84bZp2JcL1aZHheFHLgGInTJRDyoO8ENGx2fOPnj3mffXWonMGGGExS
MykWQCPTAhxeylAgvpEvZryqGQG+6LTAtHYrbGjWo6ksnwyjFZ3+7vlgH3iEZley
vkgMwX0r0SrhEvR/YlXlnfIxjfJQcSclGxwkCG5c3qZ89VHYsCvt1OztjE3N+Dzv
ZEFBD7Ng89pnfBp5QdmgAnSroOIKSNSXPOjnsrK80d4HmItiq/07PxauBTFENNNo
7Rremh8J3xNEWyWmNjCy8Bwcy0z/aVtqVkfv9gFO7u6hDlvwq9QU+3A0BqJdFYsL
Ogy3bzPdU6PX0tcyQAxJ545Gp1ZfrsayUjRaYiRWfbsXW/GCsQy+QGES6jbBdtnL
bDJra+6a5cvdiK5wg8D3gSgCTUIXwGwqNvODYiqmmJW5sKB07i0/mI7DkL4qo5WC
w+ETkAXw2wdPoHEPC/3as7eHQus5e8PkCsroqaG89JoFbgCNbTQ3AOESS8zror5n
zndwFHJolleksSTMuhdNmWf7OjwigTCTfXRdE7ltb43kRCYeittchnRZ3YHrO/8w
65JeExmWMkn7Z2nuIihaZey/H54jV1JcvjmL+ulG/ZLM0kdK4AXFGlkpmZRfqKJX
ueRGT0INYVd+b0ZsgZKNfxMlPYuWF4hflhVIFjPNy8SWVfY2OVCe1/5gyL1U8KHh
Z/b/Qf9v19oJUdu5glffy2R0wWE2L1ptASjuZIpEyuF1Ir8Sif63na3JjxfTaOUI
AbZ0lFpmIVE4ficqHX+nsPaCPSgDS4j5mqr4ubXQAShOkNjZXbbJCHad7jfHS3xH
QaOYS9crfCxA6pFDFYgrQqVMTWDF3qCY2b9xz3Y/mTy8NqKRW3OXI+yZlo4FHNli
VdH+bS62bDBUpGfl/OpjtKyspWb3CMEL9+fGWmuL0VKh9XhwO1PUv1yQvYiSq0F/
SVBo4IxtU31bH04v139+yVUyvJTiSn+ttuAD6D2HYPU7rRksDHF0phuYdmrCpcHp
C6Rrv2yVgRQiuuP74C94VRJ5Yf0kq2hyWoV+KzENuRIjSSPT1r5di5o47QiAfjkk
BFuuv6jp2A7/WCDtjE8CMIBQJpUIHBgGi98lt1ebbbdr+ETV21nqNBEzsfhZq5bQ
hG6uuC4huJvp5vwXru0gm9QOafrEI/HJ9dVJgz0e6en8QMmSfL5sk0LcvcVj86EX
v62dY2y9LjizF84OR2FtudvkelMKvp6MlDD1rPZitol8F7btSaG6jMyWTIzU/GBy
As4qiLisNiL0g33sAHs4XM2eYht88aQwwT0jzFc0LZHcoVdVSCp/2K2S6uiWbLJc
cKi6rWmON2fa9MDMk1sYIpqCWgOPPLGBtXcheDfnKZ+OCCkmhkhB96p7ap0CsmYi
C2PiMZtJVvX3O1Dr126SI+3y3VlWlstP+hTwvfmjHUBfgDeyO9NSKqKeIbhSlfSa
cPncQlm+pxfoBoXcYUieK53Rv3Y1b/fbV9UmU2yK/qhjOQhMNfkQUOQ2l5Z+eeFS
o+g95fqOXfsZUZq/ZbWZR7zjdiy3M5nNXhHnpzUz223ahuK8WSRC6n551Ux10o6E
y21NqdzZUxMc0kX8dcqmrJYVt83nj9VecZZgqD0aMUQ3YmUN4ipXarPulGOLkHz3
YFNWILONXfUAyYqr8ox4O1N+1k2Z2kMrlsBLlfTNyJUIKp6yfknVgoAKRHC/Zzkq
XE+f4vJ0mW+GWoS3rKH5oSorOgIVGcCnz9Co5IkRLtcaigQxbuuyw2d/h7xJWRtR
Urvlnh15Y1I3KdEVM/RvMdePbX7ZiJFxH+BMRsBsqnwGdeXbmCdKCVLJ23VWhkuy
nD4R5M1oNdsR5dEwU5J9v0aw0DyllED6wuznQQouUC/sqr4DGnkDr8lNwFjXWdlT
4Jcbv/WhUpTD9GiwToDVI1E0HoM5iU6peK+BaVXY7GqmzLRC4HF3dC7WIwd6bVxz
45ealHaDzDJAsS5WscQLITMhbDqnkry35kWCYvyrEOq2BIVI9b18VsHzDGluLp6b
vj8+b4bdi5QQzccv8gqA3TbgE+qAID2DcA23XbO15nSjJ8LQbGrSbHDlnXhPgftf
K1F3BPyKvwDaiCQR3fd5pjIywhM/AT5TaoQWAZQZ8EgXzNc1247X8vhoYwonRB1T
A1dTZ62vBc/mq/jrwHJBLZesjwYLMjoQAZkMXbzXAaay6bJ5TeEMenagU60rVC0J
A98VP0kzFzd8YBcMnQpSAstFofo86T71eMbRLsl35ME7igLWuM1NbwFqEkCYe41N
MZEmLIA4cKy5jqYORGLMapMdInn6tvU5pAzF6NC0RBNO4f6D9CQHeEjjKzDNoivu
H+XqwLYDbJBmd1o7hu2uzMUr1LCoemnQzAsHBs4lA9taCJXuNbvKyqiKBYpjoXOs
UO0z+rKY8uJByAd/+4jcE6M4qEJlT6aBr2HxMP0yNiaw89g+8MVZqoJEjcz4Vkih
JbpcBSQXRmTQ0auAMXc1EdcQzfdmyIglJEUpLZufO6fA3ff2EyWB2RgmE9coS2cG
PLOoKVQsQcc5k25KLtyzmCxQ/L49YCMmyUJGsS7Oocm6LHWMbhDvgKSebAEtQXY5
Dm6XzbVoAQ2x4frYYaP/pMvlHbKTmbx7gxC6Bk5Zg+kkcTB680L/ZzJCvtriCJRN
XGBclETyTrt4cr+vmdL7F6bNARrA402YV53Swvalcmx90mjdegztECfUmnIT3Yo3
XSrx6BMLFP8fOJvt39G9UUlQcFsXOuBVk1FsxPc9fXiJ733WRv0mtlOUhy4GLq/5
/ixTDb2ogg4Qemqn/9acivWczeH8+6yHlZyDvnxVD2TmOBIhFPvnoYNFIcHWSwEY
BSfE2mEQg5/Nt5Qt7gBYUizV1JSNUkOnDWx7rX2G21m9qZpxFISqvn7QPZSvu5Xy
0tSW1hU3zUSs5zm7l/AL7BrFABTEWp0qNb9cTDf5/ihPSddQYF2r2dKKQyBIWjFU
JQvKPgHrKyFEXfpkZ4osaTw1mFvzHbxlbCDei3A1agOK0PaKpBMlrDowpMvN9fwV
6NThlTIn6CyslX0ZgRgXNvC3kaLK3WdeQOO7AqN+RZijxg5CrBdzunccLFZGoXRM
AqVTeTwDQDRJBxaktDGinAt1fJAcmtWyyYyhgmn4MwJWaWAW350R0xvrGD+69O/C
k+opgq0h/CWBfEBjeyxCDQJaxFtO7X5CkDmj1TPUJE5Z3LmeGyTkHrbGrhkVD5IW
eM6TcHoaaSAfIh3h4ai1r7hT1TNWCM8e5AeQ7EuFv4DALR2w48L2a930C5XC7zqI
XjKh/yEVpP/V7/c6EN4JXPLHyISEs6nwXhgK+u0hCeLVjE2IhItw4jQ+V5gVke9l
OF8Anme8cGb73c3cKzn2etTzx2RMAQ5lS314u4Dy2hajQMJYOGg7Ew/6f9V7dA0u
LA78zCq9S7DH33hbrXXT/vIySzPSpLpVAPCpq7W9M0l6U+Qe829xC440Iy0RUJad
vA9Qinq1kJRvB8BcEULbnEF59pecAcJy3imY+cv75LWEYXx5kO4Oi1NWwE84c/H6
cAJqM6Gaqg4MFmcSbGWKssn2cQnTOBt5oS8k5UasthPgvHZRjwOZ0O6jX8Ekh9eJ
Y4i4QPdTcQcXUsTzqsxsYWEjRXccJj3u05v4B0AzrDuQqOdCGf/+Ko9Fw51/Pg/h
KKvPqwW5Z3Aqu1yy9t0zfD+sD2GrwRqjJq6/mk/2yIyGmpJg0Ua6oMBL2yVGhKAX
g2l+RGQ6B6S4gvicbw18VhN7jL0KeLImsnO1r7YjyWcheVSMGfvbl6fLbO5uV/VQ
j7ZfNmNxqjO9gESBCTohcGtAUFkDANXs4qtXp3+R0JwiYK6Rq21oln3eyn04jcHj
rsPXnGlkdSrQ+I1PFCJmkR6PpFaSi2Q99X4TM4aWg8cXuTS9RNvaBR4jo85vvTKP
7cR8vHYSrR4O+mih7rAyI6QMSWS0GMoGpSB80ioINtbNTaC39BVsiV1xyNzRh154
JPKdna80qAyo7KmVxoD9bdUFZEssOoqNvN7xMfL12rlQ5DPiW/W9/kJIAWWU8qVU
p48c1RbthNkUvGp+KnXT4u4L3awm6xpmn5zwyiubAxhlrq/KAWpsoI6MOQCVUZBJ
XYfmZfeh7YLlMwgxSQOnOcx0TUjTYD0Z0GCwkupjOdFYmicqxrOfFlXlGRDLRhQB
8s2VsaBL6FnSm0b+JtCKvFa8HbVkQ0dUPeejRUnoXgPLN613Fr2lvp0u4FvDGhja
m+TZ21MnUb+qlI+R4rSCIVzEXSbkWhl5uv/I787QPkhwYLNIYvW7CP8lvVgUT/MK
uap7QdhmtVytjLVR7Jj3U4u9UeK+LDLORl3VLS7O/KJWFXee8ltdslyCAkNsH1SP
aGlyLuxNm8OZNpju3i/2ddeLaPI9Slie5CuR3jbLRa+IOflYZL3LlLIq+EwNoB1m
5Yl/8zDXxOD8W3E0g37dvyt99Ek0iXXQuqEwR9VFG0vTKxYmHR+n4uLVFwGt9Sxj
Es7tly2vMBflKgHgbTEFazo+wHsvpSRSggtGx/EDWvEd4S0w54EPbgZbc2peqzCE
AGQn9oGVw1ujMGnhdOV4zZMtQkcBqDWawFdJMhZ02lwNHgf1dVdRtYaod1kCyQxc
uF7Mx+74XOI5tCQT61Od+lJNQ3CAu97WTcS1u7AgQiwQTCy320CTTTXPpcnEoq3L
zI62XKGc/3kZMr/p87+6d/rPO33MD9v0hNuDQSt7h7FhujRZbC6klo2AsB149KCa
6sNXXkv8F1jflQoJMGPd8n2VUFHF5dHp8mCQ41da1kRaCQoYb2FTCdJ4m05vsjKM
n/yDu0MvjnxPihuLSSyRhthw4L0+okcK3Rkcbe4a/GnV/fIwW32eKqDDuAKBpKyA
Ct9Vgew4/tVlMpN2zalulO/YYNFbOYHD3Rm6XFGpOExwLoWWMaw78/0vt8m99QuG
mHjx8z4bBEwj95QYUtYONkhs9udlNkX1i1Tki6u9nbG0LAnDauoImxvdEzk2ykXx
seERCIn3FkiHUe/y2UmEMqSE6e+E9cLJjpEh9kQwDv2mpBtIy6ghdKXaIf0FtsXH
I7pCviCPm9LS1HnB+SGFrE9+7FVB0+1KGGzEH5zgaRX1v6oPxuomwTB1BuT4Vlxd
6PPgTAjkG+OE6O5zL1QrvuoDfixcQy2nm6ng8d9PdU1peKI1DE/PavJxqA5d3fIo
NtixYtZY0TdvDhRw5+uC+j9sbVTH0WUstCQoxjG6f15Ac2iOic8y3B3gkxGEZIKc
RTHz0r7jIZda56GzInbeSnbIpysLJaOo2D2hYNxQxR2+kHXshATK5BIzvw+pAezP
rNgd5ulPpb90oCfHF9lNLD3dsyHureJJfhbj/ZKoEaMEmRtLDD2WUQogys+lF8gm
6baszO2RxnOt5l6lMpJLffXrKJN9R9uKx3mlZcgOD2TWdP62wKxHgw7GI8LiX8TH
LO3v/l/V01EdtvVEySoJc+nDsDZrht2fVlqAROg0JQS0BRsHcdV1YSEG/aJ7r4Yu
VgKYM/FoRc7NXvITCXXkmc0SibmFpKx7Ck/Baoyxic7C+qbKVtDoJzLXSMTrplpT
RiH9RsI3JOF23s5Ko/bf+f7V4ZvCmFSNCgHx39ZfNfNLM6q54pkdkAreiDClTe1c
vwAxl44GYZIl5ztne2BoBWoYlm6jG4Km6tTT03SqWXurdK2+qjrP0ltcd3N8hCX2
k5bxKPT8SU/UJ0PPNlpYV5WQtV6nDfYoDhw5GLSW3eQ/rogwfzFmhJfO6am7NxGH
NtPLlAHhE9dhsMxJslFS7zyceKvnepHztpP7Lcu4PJmEXZx/KWxExAqopAUKxUXx
gN9iUro97p0P948+5KIyREBMruTZmcKYrb/7gpFsPU56fX0IccQKNyA91BZphe4f
aFJ1GEi3cyfuYDFWgzbZZUyCEhwpXzxiecCooqWEZpGjdYpO1INTKDqtCdoDXDT0
GGIdSQpKZsUAwTI3HFFy7v9TSc28PeUfxm46S0lYYWtXHmTSdvwayOxt+6KC7H7B
yaGmZ6fp8DFxmKVfyt/cxoH0zaajKTjtT4Quk+ZhaLnyQD6VqI7kjAhVnjPc0h0L
b4GueyyUD2DImMyhPOKfQ2fYItgmE15yg9QQmZ1aw2+B2RSDxAInD6SC/GTpjG5t
JP+3Ib0Ii/cXyo9hZkZ6gD+E5tee1DsrXeFjgX7fuua9tfqeGDDdlE5vStTMJWc6
sJA/MS9GIS9Qcop3nVre3BN3fURN4mnP5s9e8aj5m5yszrlZqDORS3VYSRlKqbju
d4kpxtxukyxAy5uSSyM/0bGVn70oBFP+oliKj4/IeAdLQ0yyJF0MsQ6xkBhf0YZD
2ki01rvmornaPFzR7L+PoSgpLoN6jTQOF3lP7JlbJqfB2Bmx/p8WkIcTmEBWL7Os
Q8o1wI9xBmi50JethlloFySUkxORyE32cmQ9/z6OimDBhLpnvn1LHmICjKuJATQe
N1TvhIrofCS+IexeC2zRls+GeCNh3Ed10AYaIMxNngHcJoQcwJQFkNYxMH5GRpi8
0jJNWrFSd6IYh35Yf95/pGi6dNxvt5hxU9cfneX25dT7irm9QsThSWUyvM/M7lnY
YJn6Hn/sJ04mamiJOUA9ichogT7mGQ51CXBoJwVo8ZwduPeJQ4XqyDH+g1DoW3j6
SEzhq/z4gf7yXEN2Ds4Na8Q7hXCGJk9mWIgFDWQ9tF6IZyMjxz1KXddjot04sRKN
swDmkQZg5eG2yENhr2fYE0/VkJreiKJoaZNwiN96rBvnjRcyN2pqmZsJlPhI/5Jb
fmXqKhd1Z30OUuEAuGwzK+1UDvn1U06d9pYQhK8ZhY0elM34w+6ZFtfbdvhx87s8
390U6ijv6wno4LydP6QcfdgxVlzjTO1SSRAW6w9YWRRx048KtONGsCxA/klscDV0
1xikglVAzJowNNyhzPW3ManLsxkaU/m69qte19lffC/+PozgVZNbr+CHc+MQK5p+
WBWHit6Ogbe/0Lt1tI2jRTlYRrG40G7/OOP8+QD+GGCuKWAe6AmlPCny8laa+SWD
OICYYKSqtRr0UVM5wiCb8CA44SUldy1QqLRfk9HBO+DLvaZZspWyFbcub2+hnZmS
dezePpEQGyM+exlD37AfmoGtqL5lksNB3U0J7SrhhQffhZ99lI5j1uYgeoYXoOW6
y2ICeo5qUn6XwGaJ1htrxFkrnWskr1X2ChBHWC7qWydgtQSn+D25CKUJpn7TcKzN
De8lMolYzlL5q0ykaD8EObWfoC9/D0WbppCGPzMdHmdgF7bSrLqB99rdofehNpf9
GCIcjmKhlIyQegZGcMbTSQJNDEDhZaqpL3m0a3GexGfEroayhr0E6mGGADnS3gNd
wtaXmg+5LcIgLZPqfSKgc5g80D5kg72uA+Qi6cEOQ0SARuOPiggINRskel9qLlFe
uI6f9gBKgN2ZPLatVTweAmUpqEEOjKMNOoDmMC//wG/uj4Jq2y2+s5ZjAK4N1PQl
GpT18cMVeL2jwo84hwGbgaYHWqKpEvPASpqk9LqN6JMFUT/3x9rKszRyhGxG4BdO
IF+A5jAy3R11BdShhMQE76MWqMGroEzSRzUFOc2bBBnCWC5DGti1Y3vE1bS8WhW4
xENjXURoid0HOc8cEJH5NU9BK217wxO8liBsDpfqFIB6OEFHz+5nIucZq3K5QfOZ
GrRB8LSRRhEk9194WqPl4h1VlGuj9lsr6EzFQuZLe4/3q8aV/gZa5QHhj7k7Ut9e
7PG2LWmPh00amstTa9ug4b3fKou2k79qLcv+VEaTRIHC+IHxDZlqh8scSwQAquUl
x+mLRKq+rb2UZwVRS9CeETIRiC0TPqN2J/XuhTlwg3oAxyGCBkTnsqFng6Gl/4Oy
ePIG3cdzaxSR+KQm/qZgh9mjB04wFhhIOu1TYlAF7FJ4TUNlZtg870NzaR6DMCgr
l56wJzU47xrT9nb5dF27tagVjKRdmDAj/NZJnPy2j9fUavgQKWMmCI81rSR/yYGG
RSolITU+i2Yeg80CqUNAQRi25g39M/skZ5oHBR3WjwiciIMlrV8XXQeluUj0clEZ
ii6EI7oBqt2Pai4UIcGJApk5GMjblN/ozxOvcfbIQxaNnWWBx2x8X1LVyQXdC6yw
BkWu284LE+69+VGwCfPlT3XmTP88kchQA/6DtohyhgWLGOXUicPkBMwTJ88N60ny
PGz2WCFXTLdjkwKiFbHT8LyjCqu+5siwFvCvZnIN/oVx4GrfIBwUrHyq9xCYRiMZ
58KOqDr1GO4AylUmNZEEKTlXpIF7IePh96+fjjp1jIsEGVyeK6GSo+cHhCDqJ2Cd
5EuSGmk1toyLahmocwYPLqexu4Sb9TjLW5n4orv3P0Lcz6gqJbJ4KxwJ+LQEgGG1
c69i+0SqddhfuRvVWBte0d5SnKCBh09pjH3oXnOV9Bvmd0esstbZiKTiz1VOM/t8
BRUGoSDHl9jnwRyTR4QrHJUPmdZGMQHvgnXpxz81MLrZS892BCyCosaNC9b1VWAi
2dKCzbi/3n16mUUD09sc2EOwMd8bj4PWkeSYHwySplakys9r5O4SklL2mz40mJAP
nUsN+z1wOcNCzuoPST/9VZWOXmeoHq+Wr++CFcuUDM4c8E//i69jWu6BsrUvhD5a
nX2Gl/4rwtBA24UEtHx62Gc2JVBBnOrzSi7I5Ve9+PfzhxATZO0e+GMLCfGGbuYp
6zw8VQex/76AaWNmRSFcXh5aqHOa9X+RrxoZCt0oJwMjKFBWyyTAYz3pGHQdM1M7
En9X7iPbaJJ9BETUMdZsi+02qERMTUfio0QuuAkI6TmUX3siXX69vALT1RB5zPTV
GWlSakqLzFzcbYjHqZPzhjgPJnknXZTIyCtb7AYLBcZWN2fpaE872O+ctAl+26aR
Pk4YIYcOzdcTVEXdN9lDRa7d53UIdvh58W+gDNUtkuAHou3EP4aQY8VJk33jQeLs
HJizow/NJ8de4g1b5THnEuAvkv9LNx6iThFpgOzfy9kdgNwg2tXJsOaUy3OoQC+P
zYoPAEmViLEqzWnbZLY11T6h9/zlRYNYnNaMYRrACB7BmZ04/6MY8C42uJsKQAsZ
d+/5pWvO312cz+I7Yok/nRx3A0ki2wKmOJz4fS5CdzDAgfTGG34sZolHi9TpoJIY
6ScsNr3Qd74IPVB17AjPtWKXcr3qXOY/AhRS0uqWd05GFBMHmfOFnWMFw4n8Xl4U
Ykxh0eXooJmoM4qL8il9n2BUHw4zuVb/naDgUZO0xGzqvBQJURZ/QQ3K0ZAndbTd
zyDK/1Ssx/PzBJBer2Xy+Sn0gxkqvjjgOs8tjhu1LZ6sl/Uk5YZcPrmj15yNuk3b
WEq5rUVdG7Yeg605b1NotUaQMga0xzj12PIZRkEw1HCVp5+t2URkh48zTsI9g0zx
Ixu0/Tl79nlSL160KG6Qgsz4e8SOmnbRry+m6wWp2X8poxn2OpJ/3nXzKRbIpuUG
L5dMQKPJe/SoVAOdnK1P2vt2EqF+uI+7HCxmDD0xCSsGD6S06AyqYSQsmHiAcsUy
M0N+knUj0sez5gcT7cLFzr28UijeqBiBUVJkTHsMYCPZrz6ozZ4/YalfsV1ZfPFh
Seke81JAIRi7wGKALlntHlMOntfUrV0yWiX3J4OaZAQyj0vhjuLjhdTkHWug7wVW
7JVUz4TP0sguUUYfmrNpfo9/O+IdfgT4cRLdqrz4Ml1nQzmA7bALdzrPATv11Ewe
JZkMiOSQI5GsnzU+2ShammjB+Gw7A3b0oz0h6K7ub4CGO3yPxihgoIzWYJShfSgG
D7qQR0te4ZdYFpXY7Yb+ywzXE6xQsqtsg1GttgZ1rC1LLM7VJEPhMIkGzXaZXib0
4aPXGRgbsBawOPHsfh8fJE6hCufO1SbZid/vtvpMcIytykWeOYdyXEXM9MSWG3np
kSMk04e+bttYaiqZ8ACn5Iq1m88WCwT6IjIlQdfQL2DJcWfsuB4BUuEo0ktienIS
7gqZw455P0XNXWiEkkM6ts4l/dK9M0pq5JgVfESLdvsvrSbPkJPUipEOtxERmszD
i4+qOtvTzGPd9TE3gOyp7wstvA5uEpCmRUEai0cZ9nI/jezzVaas157mN5vqhqnW
2c8YZ0AMzymh/kLueCaR13oX037b9wcTswS7zbeDR9NzGE4gHqXyk0dsHaEy49lZ
pQJBq3TMvDph5zAUDA6P/n2E9NTQ8Ki013rnQMAeRJm0pcwAZ5QLfMsQDbghbzue
c+7pJetmK5HUZ6MVmYinebWhVzufQGWbsA5DlQ8bPEAiE3t9sYxlNlaNewXDQNgP
EZANfZytxMwkzMyKp8/kMLBkJ6GExdttSLFdjfafh4u8h0Oq1pN4/FlqpIxQzPqU
zeQEffGDoG0oYpdogPWdbV/fVA/GNNkxsnddrp5RSY7k7cMyx6jAwmt8ACwfiLHX
p0CAhey6HuG5tCKcRw4jrg2priJ/8CdG16QKiHfqLHf9xhVCngNVnuV27otXMoYA
QygtCCfgs4xf57j3wiz08dwjLo1lICFRKEbvX/3wHq33Sys2S9KRpPBAi4RUt1V9
KU4gBnMP5OR67dr6bHnbG4iteCCYWGIm7DgRPN6f/pBgd7MWSykZGzc/HKTTwaDL
isNEiuMeh2T1WQ4jxvShzRMf50ebn3ODiyPMPmv7epMJ49l+dJDVmQQIdJ8CvTMt
L/Y+IOOAgtx8BvLB96AfRwy8oZFyP2OqAnDJHsjSC6/+H1BFp/Gvm429uL67ieoW
YsDLuAxmcWjF2UcTM5rZfPHHlq8j6nXmSK5QnBZVxbVmr5Bx49F+V/EOsxTRBDRc
H0stXLv3xVKIcQfCX0lNBHzKF6upa5DJNGDzS6Z1rLr07NBdIdUFC4lHJP9ABccf
v72ItFx6hYuWLitUPYjH7uVE7L0MlTJLavaLGGdpPUd9/9Lu7JJGj/PJZQ/awpAq
+NVPSC6+0ZtKXpv5mGVIXln4hzCg3CYLCMHUkLOKsl58/WHBaVK/knpL9YMpxqWk
zRY2UKZ8gEyQia7Isp8oUwvHwFz9s4fUysItIZc70YyUFt5toSc44McEr7935fUu
h+C1gcjiKjnf3zgzxGoS2aE2O2s8i4rqOGpL6BfDX16ZsoGwVu0LS8g8V2OYq2ll
nuImZPolM6ogtfKXfg+6ENURqkFIjBC2wc3TN98TCi03dGKWhi6rAoDAZRaIIL3u
tOAp31GTzOT1kRyVnVxdxxXEqNUj19nE9gRmTK3BPhArdmXTNX3vSlfOBWDKfrFb
naFpmZTv1MFDtAB0QHuUshyf/w36/kQOcXD+0w23yzEhxOfx1DxWePJ22Rk2c57T
aH1P9efU1KcQnQoqIwDHtqPsoEvCzc/bguXRvZChMyKayIikzMO9mopoULQXlMe3
FpqSvGk1ZP4YJfZi/2zaloYNmMzM6J1orj7tmsf8JxrcSH54+s0Nmj2OBlaUvOeC
SzVboZZu6SfXMk4DIVqgYQSI1d0iCXbn4KjLZOgk1RHtpYtFSvj3gLIhQU5XB4OY
WRCrAH33d+YklYUGcrymT8/pYtQFK2VVYVhL1d4zMlCxZb23/mEttnPtDkuuNFML
BFQ2Ppa32k0bLwONvPXqJr3SdAfyLhGA2RbxqcrXEjy8fOR9MjOjHZX8U1BKwjVA
A05tGZvSoHLqt6IexSp+GYm4Vf8Axls+puxqCVXCq3vhhKVt/NP2poyAk2gA+LE+
UEix4dO1OgoPBe8XRBDOq8WsU4mcEgxz6GpLR5u767QkiblaLci9no1LkbIUL6CA
nguRiXtyuZT8e1IJsX2s4XAFVQVoCnDHULWctwsx3CqolrIigis8unynsdqssNi7
Z7VJdjBKT+PPprdoOCEsi3MKqLDlKcUAgWUuAI/YnYpQNcMKu1YAfsozCpuFTVyc
sE3b+DEzD8olJ2SFK6HAtW7A2dWY1F42x2AAOEbMhtpsk+o6FmKMtpNfiAZLbYzj
/+WQh3w7m+bEUtpvdKsZrg3TsyHMdeAxh6H8FsrRjsdJdSmaHR/1C4OcIA8yJCMW
dNvmRmSy0n2ticNZ/Xf+ud+W9TB6Z+GqtAyGBn+a/FnPlWdDONbAUHjODU3hCMxS
BhfgIsOT9VHEWfhoLbBoRGgYX9oJ7LTLU8ADaKhg/AuhJDnc6YfXRrXp9Hcc5tQP
ztoot4mC74iDdo8Z7uwtki/MyzViQ2tQnLC8o4j0W4ZTLiXmRIax2THC/QrWMdjz
8g9jLvZPpsMSZl1IVFncQ79L0CUuC9UHwBcCJ8+xieCOgLiGCNovRCggRbRd+3kL
fjkzHDus+tUf8A09s4BwhX6/L/Pt8RMmPWFU3I9mFPKceBt4Fa0n+wOdwHeFeVq4
ZfXJQeswHWnVV0wsc4/9Lkby3ruPiBv7lTjYNmP2lRp+QjA8QbAR64Lztnc7dAhq
Ez+DP+YEVC/NT4I86+6tn9Waec7W+iThDUuUqNK639FA+EUWZc9DgAVWOugrjt6P
/hOloem2CgCB6FVZyfDE69BtRFGQ7E6pnOJ4iE7v62G4OAPPHAuzeV62RHsD4RvC
l5vwM6/HiC4EE4xwaMft9nEiljjBwtN1mlTclQi2doVMWYadhh3MeorrkpY4IDJP
raFyZSE2PSp/WQzj6nPDDqh2xz7TsUxCz+/HZf2HFds4fEFonvKub4SclmnV1pNU
4X1BGzRjR5WDJlhCPkUs75Om7OwBhFXVybvz5GqRAQUzjV8ETOZpr4rLW0gelFfa
kkOtb9+Yz6aKBd47zJaKysiCz0Y4YXg1Xs9p9fghndmfv45X118HWIeo8HxWSKe6
imKz1R52zgOXtoywxA6qatPcPbmmW9IkAmyc4Lmu8YfsB4OgIo2WuoLkhDyslwCH
h2YNT+DrhF2YMs1SNJxMnFOdD+9yCQk0jlYtylz+VM75OdD5624TjzA2HEpthccL
WZUfsvWB2ZzdLkebwPv0y4DUGCP3SF2S+tL1OhH+YYmiA8zBlzv6+wGTHYh9W6CH
5ww42PHQsQuPz4By7aBBT8+rGyRbB0VVYRP1okmb+XLgKpHDEhtEWKV9KSQF3mx7
hD1qq8F28M53AcqXr0ZfNXmvOhsP0KZcJZXrzeA1J66bvdxNh4L/Z0Uelcg0v1Dx
25l4KzoX7HHD5GBjWttGGBSQpq1xqAFqPcc9kvnakj1OcRiDSjJC3h4zZyCUsjaG
024eB2gPkrZSfBSBErdmko0VZrKaszaBOdrY3y+FIhLDQguhh30GVocd3Bew0LnL
fQgAEJ7nCh4nWucZ0ANCMn5RGGF78WWYcZu6rlkdpHEreiaPmrBvSqCAGZWvDuRT
v6/b2pBzZjIt5DvsRBln+YRF25q8Hex+LqU54v+JN6/fn6GW7k7vCt9gX5Ml91hQ
/rMK8lV/N6hItrwXsmArbIVESrMJzKuR3ngSPzSNVqjvpb2AqmCCxjOROhbJbtuI
kZpGDDJbju+qHn4DZtQ97poycMkwtc2iC5H8fqm6pf8oQrGHw02YsN3fm2PPyTr2
jDReVdI48jUvDj9ZHzG1RWIype8kLYn4UI7CaXnOC4ttvPmpRidyeEFT/s2xG2bT
LEKUWxY6Wjxx31PcNilQF03Ivqt5yF/QP3pzNcmw/RMvdl97bENSXChr6sox1IRz
hCHNSdkpYHQeoKKE+PdprVqXcGn45SshcY4UJA35GatuwWr/LZOTu3Ax6gF/hMUP
wDD/0UdP3XT85NeczcGDV5XBhl/Wq+FQcTg5HzHMl5it9+6q6OMeGgMH36gLou4y
wTDfvLq/iLYHbge0YVfeMZBAJjLnl7gNMYaGnF1rbfaTyZ69K3W0rTfn2cez/gXz
Q/51JBaJ2RMkX0ZE/eXQhDjVV+4Zg/GEIHCViimMsmCg1dtxYnUDPF4gJlmzem+B
Ky3WNcYUepK8iMu4ztIClizcATd4IDuCjuHj0zSuK/+6SUsMMnZ1UWzwScL1o6mZ
lHkH3OeJR7DB6OklTBQi6f+98ypviZjxPEt/DCihP7dnSfvacIXj4gYoDpFlFESt
3ccovKTspJJ3LlkpJFul/Ds/ejGTqoVBKN4/2JMyYvbnKusz8blOQ3fLVWO3yfq6
PnvKKKLalKHFVG+e6ey4V6gjqajmTc8dprSf6HZmrpR7ZRvvVlHjoC9ibDb4eDkY
j9zI/7e2OplKmxS4Csgy7qpKBns0qT8keuQCOrnBjZGwWNQKbZp9iapFf7IbfhUq
yZ62/+ou1P4QlrPk3qWMqCwjOed6j9nPUyyOn6Y12Wnw8Z/du5nMn8XkIt1coUUl
JpW84RY7IFN7i8CmjwxrpJr4JovY6EfuTBT5r70Hryw9qMGKWJK0DhfmWiif5Whb
0U44EbySkKo52VuMAjoVhK6mYqlNAhwGYVR2q/29ZGHsMd7JqfRbCghGL9Mt4wI6
UjcuHJOVp/Z1R0HON8gdeEuYA4dRP0J5nc39Ucm7lkybuFj+yPuuek7dnFt5EbTK
BzDRcDxUs35gNS63c8C3pZT3KG/F3NdKRq6MfykOZPCkg7p48j9zHEQy/g6LP+vG
Zigh4jRm+qabzBuxxkVJnLeAkQoELgvc32/IShoY+KDgXx+bKhWxPnjLUJFrhZ0N
1xkSNh4edThigadrFP9mNyIoxdE7arLgQ0e1gRV6tQaYoRc+9tivUHBw0YulA2fA
MZdY7nxKFhFXPsTwEJqwf+hHQFHb4y9nyFDklqeWZxi0T/jXy1OiC/EzGDvlkPlG
Lvovusm8nz7m88+cadONG+VT4vcMqfnCiUnkYjChuhK+7BRXF5LTB9WC9+WpQASS
eoZZcsVxTHQMTOw5hWv8MRcktxIaS4Bf1p/DiIhtGm32ZS3eNMM6rSLY9ebhp+Bj
7fpF9/SHIYUPM4FGSRmLhKb4HR1qx1LJiNIgZd2oGz32wCCCrKgUg2rrqerb9wjK
MsxVqoc6fupfRz11GOeS8njBShsIcBCdx3z0coOZph9SJrLYVyLCRdpmXEEF7DPd
luMvNGnhCMkGCF53WfDUdjpgeTytPPENg+bNfsp2XeF0ZvBRZnnefhUUIYwxz1o0
5iT3S/NXjmn2l+dxcPnO0MsWrxNNbqH5u8rxIzWgcCWZNZ6PHuQ6aw7ddY0Qeshy
TtxQrAkkMyDvveG1+rhpVBblzXtgIR10ZDSLhXKJb32hU5Rc6kz8O6bb9e2K/GUY
s/ToyoC47fZ33JZ+/tApyo1qULQz/5qUW532RqB/FM83dHJgfxVNM5veXogMNJha
uDWS/bpYNkg/iKkWkWcRNjYOuasKLg8/4rqU3bYrsfLHuYyjVrV9keDldHp6r3CF
qSrqCbkcS91HoZBftZ0cyLUkCJaxYdKGpiYrn6cH/eRRyemYMGzG76HDwBammYKE
WNrc7PaXosZ/E0obfyKtbIcBBLPZBwl04BojtPcp2zsS6yf4LzYk6FV4V/5wTGnC
NLOhSgN+kSQNfPFqKKkw2IEhCYJgAvCe1M9mEz3REJ9FxkRgSMEgctkZou51EnaT
IVPQiR8sF8P/CQiSl1CFYvuB+AE3EYygtejREL2tNFto01UQ2lXf3rkJg8Q389CV
NgbGdGfcm24TyBB6MPU330+z29Uc4roQ+Rul+WoDa9/5OXV2l4wOdbbC4OyEBIaC
77p2A9bLAxmWtEZ/Vzq5hg98U0+b3WC0ipuUAzvrbnR4Iv0VV9x1eQgGQ+TJc+R1
RLrgZv9hQkqjE+5bDc43n5iL1VwFVSdE2SMMR4rim9wBJDR5D6tuPVx9PH14Pou9
mLKmK0V66lIy5vqqzF2w6A2R02wUMB/rDXw2Dvx75+KRxjIwRyA4Y29lra+iYQ3f
QpY3tKacOJNHP/idtQWLz8zCMlq1OMhfEEPe7DoEiy0tpTowoikcCyiWTLfrAZVL
auQ7GDaoWTa+cW2dCZso52+Edb/VwLVSPthhw/b7ZqvARQm6paxbOnqbZ1aaDDio
/aZt+cPJOnkis4ND82fzDjQhYWC4B+zMlf4XJTRAa1qBv5fvqYGgliejjxkgbbpO
s3ImgnH0N3/gLy7DifTJc03FmH2YKedq1/je49ilX3baPGBPHYYvXD1AzBTMpJ40
2IMOMb9ILWxrJQcBcuoIyAFSy+Hy6gUFBCLJYO5m6Its4pn7PSHjQanNGEbluYlx
Jhx4vyAzstctz1LhSXxTz/eTu2wBhTKVTTFXF45kaY1TtebpxPQtKtFiJY/wckmR
i5q4guujuk1UqBf+klw4awHRhBw2uKu+NG+PV2604wgd9Tq1uxCWh5Zxp6U8AKsj
CV4QT66ttaft7Gc5Rf8U3wDq3dUBdHGfgSmiaXusCo1btslFlnABbaGYGEh0hN/g
Fc8Y7p2Ac9PKVnygzIz89IZfKKG51qEIkIBqkKvN1NobD9tQDLQG9ViimxSzFhbE
eeFqJcDhOcud//yobLexYK4CLCwJfsUe95nlclhywFuLvDtMZqJivwFvsuX2xLRK
lHiWNWEP+Pfw7fRRag4DnV+FueNe3uM5FD77yNVBc/URDfPU9ViagtIeSijAgf3Q
bdJ0lU1nkqeWczCcQIiTGW76TZ6Y4Y/0JaQ2cZ0VayrB7lhPkCwBjJDPc73pnVYf
FgzkiuMQsTgY08aK3ARgw2iRvaXfNRGJuIQOplvIjhrwebnviKUc85nyvlprkmEG
ccaV7JvY3UDck/LB74Gy8YBntk97kH4qyejfRPBuKfyXYp02rau1T166P/zPGp59
KGEdXoEOpUxAKe7/zMHh35ZaDsOt+5p0IAc9fnBC+s76/hzkmUi8zmjIu/FC0mFE
g5Mk0dEQaXvw6+/TMXaYw0DdWybuZNoi/kt975uygozJ+JHoiAEHX+ii/l6OifLU
qfF6VKWTjeC6cmOJ9cfAfdAsEK5GVsYc51XloGJcqq7n+3WNHAHqAnb8l3v7edDm
bPXFLHoXuI/ZxpsFiyDPISWgWyu4ZF0itaykZoh0udC0OzQy2z+AzAaaDaXVpURr
YHLPvc/Ok/O4whdFE01iegU715XWhGibOwUSF0ge0e9SaDDH+Xod2qI/1cYJF77M
aEK7N/yZ52kCepnqvzKRAaw0/rSqsUrwzzCdzdY0Qv02SQK3gFIEkNSoyYX2GB0z
m6e6wnBrgsnit5GYso9x5o7VCCnxyAI/MFgJ/v8STMFdoSxISV/CIvTxUI3BsCpD
TWdkCGpjCmJeAEeBTzCstwpUwWS/k3fSgd4qlMyyiwMX+C47TDQgrJ9ND6quHoQx
hLlsF+KyPOJ+vtg+iGsrWj9kutnYCJ/NUlpiGkmXtmUKXiWZInFalA5Qbdp5hCC/
Mi0wzhKBHdq9yF1MdC1NP5U27/dBkiFv8isY05y44fHAT0aYA2SizlhstkL/idkk
dHfIvQEhMOSjWPBheKp3MZ3UxIrD6desK5w/8qyhKwTmscypmGe3QTREBm5+Xac7
505YybJCBgTMRaaK/oRwt3Eavr4iFOPLAJXf8jy7CuTN/MKHP9TfceaJNgqPciFh
g9YG+Y3zuFweH0ZwFUMPrqSPNwRwH1739mo+V7SrOo51b2GCnVENZKR+aNQ/6zp+
N58QfZRwUD4+ZZhHDfBzQH6xCLMB/Lf0WqwNghSv0kBY6RmFxrQU7mhI+hhvq7R3
Ml6SsE7hg1wWVvLkCenBkKxckE47PJchWm3me/5MoaSldF5wJMcDYZUnwlPQiAKe
3OWlMvRqyAdZwGe0CJlDrMOZxk8r92vC3ZgDyiKFOy6HxAesupV34tkJrGQ7Y4fm
uje/yCVe01At7L+1ykWh5OH7unBMCHKkYO/UBbD9HESdoAPfoy1HQ35VuIQGqsbi
TkIrTabuOpzHuYE7O00Mo/Tkg70qcvcSgXQ63PHLqbqddYmN4FSV2b9kR0+EPMd4
+D3FKQgNg2hZmQ42sMesKN2UWS7+cHGp/bxCf46ICkvcb7HKI2BFELZE7LV0A7c0
OsQbf4nggIfTeR3uJr2Fd4LUZELpT7Ycz5VnV1yAldtHVVPvztSLjB2Iseuc2ZNq
L0upfKlWx7oHqfLaCJtdVe5VTgY+buu0hCJqHvJAvYC17nHdHLSGxiA11yOBHs6v
GvG3NNVrbie3jej6Bk8CzrjYqM8z6DthO8cb6RXb6xV9utmHVuJ+Qq2oshp0ak0a
CqXEFhqk3z9j9QmLTA9U6J0C9LfwAaefmo7Rb4ymIAvRmkUuF8MPZsN1uDxVQJzf
bh6A42P42p8pzKLY+BokgAHFnFDBVIvV2nwaUAHQCNodYEgT4CYBfkI4r/2M+kV7
SuxU8JLVE1lAlcLQGCIKN8iLMxR3pQt5N3ROX9XTZqKfJCpf96ymICpjhElyeyw7
eDRT4MZ7l7Iprhfw85x6Yr0PLz8yIKFNc7dbMQn177IQvs7RPJ1dDp5iu8FqHSWO
WyTqILtvO7SYRqHHbLBzJf1CZBClXt/1SLxr6cLKH6FTelZ6eDMgmt5UOYeWUdze
psrzhquyfs+LOFzDjrNvDYSQoT3PdOaiu7kYbSN/v1dgGrje0fzHAdP7q845iFD+
Lnq8NuTKn9AKlgF33nB1gAvh7HFV5KpEai8gy27JwFK3p0UB+Zd03qwHE1WeMhAx
XNXkT8oLnU4olNHHcYTkCF7/PolxIeuTxqfZYb7e1bpYX1Fepw4QOQK/CnAi3YUz
MQZtiJDxkV/C7zqtGzmnqnE9Fz6QJV55jeLueYCn7WWx+/b6C+0TWMUXhE6fn+Sa
dGrh3QfcR3X190T9QhuVlLQ9i/mCxLeeV/LpoE10I7vD+LgjUchMlNCZuP5gG9JU
Km6K4uFTf+vZyvbRC3TEULcpm66n+X3+hbqSuV5Anr2G90pTnPodPfWEuOIAe2WL
AXSWVJyVPEAoPazHRwd5nchi/sSJ4fMJ+BvJmLBmXpjfO6jMs3OiqsxWP3YcaZx9
FsxE82og3KnTV6u93DPVloQF0WV8hgabSIew+ZMutnALQBRht4eL6fha3UXwy/4M
w6yUlRUyctHsr2O5+nhE5DeoiC3ASqYovSdYKlImVcYaPEnz41iE7m7q5u654NSE
SSyNzzuIZztIWbiydeYkRJYAsMAwDqLLqsdhXrftSA8Vsce6yEDYV4/RaDlp985P
6+ztR51kA76Wpkgu5CAttabCNp6Pfw1kVDSPMJrtbDgiCJJwGwi8MqfI9bgBRGWN
uRJlzcouP/f0fncbHW7vm+HshcAAVYo4p+Jg2GURkDpuvY/p/g3ES6pUB9KxUflX
tS846Q3NPMi6dskL/tGJrSCwyrYL+OHhXmqKpE/yEd/nb3a54SB625XGBXxBiddp
M2hogny8lzlNjW/1WQ2tNoJDFK46bhJ+E8Z2xL3oZbAVn2o4lKx/oOrKzJ9HChXq
3rU8FN5DMeFidcgMCUXxA2K6zYCBEVwfh/snQ7Y6HlgQaqh7vHkPNAk+JnFjMne9
b45ga2F407FSl1zByTJxdpiLvahilljWqlRxf5jFXJCL2f06tkatU/p09BH/a53M
vVs8F8EEKUiso2CB7JN3drBkhU7Axt3Bmgcl6KsaRVpngFHdwf3v+OzUSEgzTzFb
X5lSdcuj2EILKYeYSth5N7/vRJ3I3eyYY0Zfpy8dqMlRlln/nEmkunfAmuF5MXRG
42wh7CA/2GlB6xORTChIrntc/Bc/xQGSc602oYbDxWm9jeoqyJ68E2YNJIN7r3wq
7XnmZ4eY5dgmax/xTzWxThvy+TOHdhXJXGa8Uc0lgPbU9Sj9LtLG7RI2eOro/0u4
XSTHHpzsDw9oE4+aptuA+22vNKPgYQEh4+RdWX3W24VfIPTGr2bhNaupkSnPVR6d
uQZXOpe7INvzexetBx+ZG1WW4a0+Qe+c8ZlgufR7HJQryklf6qLNVpdBdTKuQlsV
4COrtGFa8P5zz+fVvCptLcmzWG7RQiAjPjZk5e44XEIBZ6KiFiFaynwznlS9Sxro
aGUbXrKe1N9qLYzhIOtEwi/rljcrrmCN3qZeJVRg28rXPPjSRIFwnYuANItAjsqS
4yunR7jdebwnpM3HO+HhjK8yACdIAY0LFRPIBKr06xlsuTQkXyZyAjA4obORjMui
TcdOC2ROJ1yE6dPqEiV7fWfwrF4BRGDsquCBP8km6cdsnFDSwIIV0+eQyrKKxXGa
sG/zfUfMmS1SlRbptPxmM/WMSd5QwJFpp05zzoCberQCUDQOnfbHQP040TwJ7GbY
z3WzBbvgMpUGoYNtoRHLMADP2d0HSHazpICqKMT5la6PtvDhE6qO6QCpUG4hNFTX
Gum/TNM6qCc5gCYJJAepEvZ9E7Sf2169ethlj/qo2xSHvmWj1Tze/CcSsDpP0qJT
8vwlKdRHna/k5PzJAtbUNbvw7CgVMyhfn8/so3jJvkylEjdW0Yb3G//pEOf8OYw8
tROSo4Bv/vAm21Gpj5f70Hgn228RNEJQDInpDVZDxvmLQj0Iegcu2GsD9kAHJgF5
+ktcerLtCA5g35eXQjF8t9MfYH0nZz2MbHcvGPcOYw38ezhk32GL7AXIAXL8xpuZ
Xs1zNsy2OL2atQx62hcUK8pLjYYg27ycF3FMnyyiE0D0RMlck4PnfptkOYIbBNkV
LNO1YxBZKalUseNH5djFbp4o+l1wmouz9fEWYVTumgfNUHiG+QPTVzBymXCmgCiG
gQwqyvv+3j+ZmJFsyIrRGgbDf97nugqEIchCUfPNiRf1OhYhoqSSlBzaofGbRWaL
VKP11F01yl0M2coVbucjKfitMZD6XQzeDjSi9ZhXfR7WrF4qamg6E+1wyIhT2ucu
nCrAE7RLjcvSyXGqeB3ohA++Ht5OzwtlYM7D8qydr08hdVXEUS/eyfU5wbvjux+M
UT9nhmQBeZreWrapFpJ8R2s9YOFFsI/FMB88xSFe4aVWExAIkRlJA+GGQezjJZEe
08Oxtrr8k/MxPqD4d80Xjp5ntS68qMf5zqZqVqETU8uGtIKIJmHa/38pcTj3aJLj
5cUb68tonWmeP7fvKzlwLjFe/cvScVF5dbIO/NIxbrNssTeATMbTesga0xeZ6HXZ
6ey+QZmahRqwcbFtsQsWjKNsrT1wLoECiE5cDqLwOaWDi6OpSZYdUzjVfvYjBWnA
kUUQkUHLQ/g7VUz5yuiAY+6W+nN/sGUAA18BfRseSbrKYs5s5QyqVvku3QWV/GWT
sYQfVVSD1IxfggO2Nxv4yqlRkZHf+CCPTrKr14Qm1R9mnly63psyX4BJGqZrYHPC
fSE9hj6RQAKUkKMbAF65F+D60OwSt5g2iDNn9hRv0tFjUHHipVHHFrydQVBnQ7s0
I/5fdGW9LbCJjNAkL0I2SFlbXsZCqIvx9C3mhm2gewdZSNce3qiebE4jJ6apWnKG
LI4yksKjocmkFNPZjk+1jdsj31qdmP3MzLH0d2BUkok4aSPJQIZX1nWjQspmwk7E
FUV6OHCW+JwHgAdVeX9nTYrADGN5yOV5oNGJCnHzqQFM+xFV+zXgzpB59U4kH/vC
QT7j4iBuuqkpGfugDSqxEfdUyWWLqI3XvZ2bQ1pDNlGVryY59CxyApXBpMqusxPC
YlZLpZJ86zg/V5DaUi+hTjnvQmeBJT135SQJIP4q/ZjTSry5wn33gZNH9RFVHZXv
qY3y2fXdhFiSxYUreMSk6NjgAA9WY+wUdVELExhJa2H5RzwauB424BlxkM0dryJq
2WFD8+uG8mCCdP4xvsm+grdm8lPuUlbxkwRj2/8pYf1S7JY2vZwFXPGmDZSBBGa4
V0GuZ3KR6izR8Crv0/LX5snKYMR2wrn/Sg7Jx0W8TWMPJ7xjEnI7SHVARcrjzv0K
Gbd4x50x0/nNIuZx1t/wvr8mNIyUFiMiMrVzVI6Q5dSapNEd7uIdIWQPjkXxq6YW
Y0sOJRSfCqY4ZBQW3iMLtUQwsoUXA4+qSbExnHbx1OyhEnHvoGxnRdMmmB0gz5MG
gvMrQ9JgeK2DZNZ4Bea2y2TKoDi8/nslZBETWUugSUWzbz/LroIBHJ3QGO2fHu/d
9NARA8A75If/diBtyMrwucadTPoPi5FlB9PSrzxZVdYpIAaDasLA1UdEJHkSCP8v
TM9QP51+53RYc1b/PEeh1vAy6CoNuO4YH0ExrmzkNOzxxPKaHfcM3Et+qNp/vOuD
cmicIJ2V4HKnTGn3WYeOAVzMz0W9eO9i0XPcLNZN4r3k406wLJgouphVYBmukAB8
8a/gj3DNpMNbHbiuET4dlK9UNitiuUM2csP5CzeeQOGRejjq5Fjquu59TErUYxp+
b+zZ/xbSlfyT7vCiiGD1hUlngeVhoTk6RSvPGOvjQtmLmFX1Yjt5IVqsx7eOazP1
YtBZo02KQpC9yLkRQiyOU2AAXVdMK/cCajh+C66Ho9G8BDxDGc6RwC9x5CPklOjx
Z2b9Q37ombX13w+AwxLWVLLbYpNnssuMPGMoTna0jAAMAEEBL0lUcnP80bnvP10B
kaAFZneoJSj7s8JRL8JC3QAFI/WVLMf8kcq86+52tjYElFV4B6a7KE0PEz05/Beo
dO96XzCXfc4f2Kk3+0L3tAHcMI0TQhpmYX6xBms1qlC0/85ZMl6LW19fDTN0Dqxt
qoXQPBTf4V7mREd50kJ/XBgEYXnogBqITx9aYmuL5xUqy7bjV6E7INnvqOJ7nGdQ
mH63XItXBY2df641y5DwuqoqUbbfD9BjDmoWcy1ZovvPHqPdUacMtMMhyJV+9NIM
N3/g9Xtjp0Irmw5f1QrPwlaNmvhitxq5PgeDOFpQoJsyi5IPcDznDLBg4duF3yCO
3+VSU7azJvlz26TyzeKx66d3BFJnQkV+sexmnV7T/QEToIcadIaulhFixpn2AFyZ
siRsRsiQV/qLbvb6bK+ZV0PBJuCBdO5DDkNaeQUQModTRBZS3mupZToKsSdjhOw4
kc9fGZ5PQ2eSjPIz901RgPi87FHxosZsP+I+GFn18p2zEKqxTJ514cF2lzj7cb6m
QIyrQiGxrAuYl5ZaIwnSTmo3fFf4yM2CILg7lRTXj/cW+xP7TqO6G3F7EVn71Fqu
EDk7VIVJd5bNHFtbwhME2a3QjjkLX1BK6wYT5uc8swqEXmPYl5vdzaqzE9Y23s2B
UlL3nr1qnXeFewNo+Z2WP22Efi35wIFxbVSd0eSUf7UpdQyMN/V+LjLeenc85cra
KDzyEgCust2AkZ1OR+vxMYn8LhKstLBpAnyORmdS4mniwBIBEqGgqvZCQIwxKOze
EkXcBkRWt8wGXmbgtYU6Z5DH0EeSkVZtijN12Tt7M/FRnZogE6d26UXZzH3YjVeu
1MmwdXSSvpeZi+qdlPLNeRHTqTfbnqr9YviLz3Upbpij4EU8M/SkD0qiijS6MJcs
dKsyblAx+nVbqWkCBu/9w4zXIwauEQ+2+WTySjWdm9NpIeJT/x5JA9M6hGVzHYE0
2KLe9Nda9uKxw9gtJYQsqf5BhPe0PG216q7RTmYtxBUJI07kvqVKguxRm4FSApt+
j6txerfpAJ+NBkflWN32cGmrNvKdMwszXzJ/gQydfnTYGnw4vL0M5tSqZxP19jo8
wMa5V52Ayh7gaZ/yZ89JNH6h3kRoTZCfeNep+wY+qfNwQ1x4/ICjEGHoilkr489X
AS+tSUtTcopmTD6V+wquSWTsv++Rfmc9tXBRqt4znTrZKUZj0vQ0xHjzfyptak6h
gGzNaJYYcyWG1mPZR5IgCjFZGSpg5H4VueL4nJNX9ll9LFU/ELegaF9cJLvcClx8
R3/XVBUwR6jwPzyRmDwvtK/4tZR9Aq5d8VtXkodmVSFWDCBXC6uLX4IyjWRmTbJv
5Z3OLKTbV4jbSNeVKDwvjncG4/Cx3Kr7G06Xhx7dO49qiNxrXUKjPOh95qyqsX84
vWsTNL5B+JVF2oTE3WFn7EGYcSehjrWcTB4R02ZtvVhmkNkwGlK+1OO0uw/5CkmQ
51OgxXQIoipqccS/ALkPABEIA21PAIMuKJKWiq0cGAm4w/CwD0HSAA3XvpzqNnd/
TDAjhyYnd9Uis/DWFsE+i0g8X4EOxZbFvFZOTgrw7eP8Fv7RC7Fd9kCHrmIeZv7O
bABjNLSqm+OjaDOwshMQKJh5pOX1MttEcf2fNnulzaePibJW5YOpfcBssKXK5ftL
ROtM7hTzCXY6jkWEjGFWXbxSabw9331DuF4cmUTmWWGN08Heqre+Yiv7GQla0yhG
ExeY3NXZKSvqrdvsZilAnCl8dOkq2TmCwjrQ0z4k0bteYusCmENjtQjDJSHG3f78
ZbsXYhncKujSOWA7szr6xMYcEjyyKynL8TMyzWUSFDwvYwjF+7QIyFUmXz5kU2vD
WeYovYEusgeElHuCPalPsgQt/o9UTBcwViSya0Id50p6Wa8d7XxZTREe+qkESZ6v
E1D+IQxomM34bmfJbqBcVml/PjYhuH1hYx8yLJra9DfZ9MEiHr3dfDFmILAX4gAX
hySaMTDD4bJKwycBjtc7OgneugD6ebNGV0QzKVNJ86rwIzty5SoLx7eI+qM8hRFH
QiQtzEa02vimD7pSmunc4jr1kJ8g956gwbJEQw7iGIpzr+Vz1Y+nnkk07ocjURsB
rZScsesD0cwOcbF/IpYDEOvZsmTm8q79jv3AOu+GG5czg6FZXzjgBGengyj/NSIz
W0csCMaweZ35YMLlUjq+UjR2KD9Qlve2PIHGw8gVDvM3cXgffTVprdXMDxb5VFTt
V+bxuViDbp/AFQJ8Hc86+s6YWi/9sFZSvOAD8W7BnMKcOyiDDij3p31dshgX55tz
+Wy/O5ZqttvudrZNohrIyAd0NNAoUJKD87V+34ELZS3dW4+q9DwNTuK5f6pFBTYe
R/WXtLRX9XwLS6HpcVbL3jO08WgjioISVLXYwNB/A/rxlLw7VXKxHJYTDtpBKFI2
BXPokKdhm6CkLwuBrJrFTTG3AI/ItLGl9kOPHKdWNhKao2bPeXSL13eV+VssZ1VJ
KeI5vRUrQrdCsLavrycmT61SCqEknwERfezzizPoydGwqKyPNnXWojIjXhjDfsjw
QdDzADMfwVf98ELsXsWMInGVbIyu1nDN+gB9MUsqHkXRx0Tfk9k8qqQ/LBZoXLbt
iy3Ugha7sEjymcz8JtgRzNIXyNUYJurO5iFwUFUDZbpzc/1ODKZr5lek5P2SPA6B
C06fanKOS/Jy/sCcb9zAAi805Cuq2rloWh8yh4Gu/CJdAKUFfOp/In5HZtUptrtJ
z4yNqaOZTMoYdDxth37N0JELffETP+T2CFU9sEDhVssij453c9QpOPLsmIwbCfYK
SFqzo3WhgUYzEJihCCXXUiSdL44NhXmm4sMjBhh2qFi+I0rb4SOXkqvzLDVRmfCt
zKPLLVHXA+UrwSAwiCCqNvBD6THGCr6gZoFCD/tEdFflnBJb4TK7XptKjubwcGrJ
ss+ur3qk6YXT+N/Mssmw45HwWb2xJwJAVsMFXA7ct6kk7SdmCM7jROiqOznLHm3M
8iJWWKLytbfOKXCfrxOH5QUUy7is/gihq67pDZaxnph2wHOK+5igC5qntmzICLPI
AtOtFoJzwlAPKxP4vqe9+L30Fa6E7/0eJCmyK9Pm5WKsGDugdD5tgYVZ1A4dJIoa
xOxUwFCaPS752F8pLlPrXW/uod9FmSE4kzrhZKr+NQEMPVwwypJHwl1MwqD977lP
H/Kbcah7E4dXcZBqjsO9vYScaH43KPwqyu4wjB99dobyVkaEMKizPAnnELFk+RB9
doPALHjHlspH5hUep0iUlspTkZTDtBLnJeuJCN25A0UR825oh8LkYrHxmyxJjuGS
RE8xXm365LE4kzu0+yWhKgpVxisaanU6CujTA89DtR8d6VedanZhzzDF6Jw+7UWV
NrZE0K9/ItL0Qj2o5Jbz36X0Xi5OpeqM1ly6449WE3N1COzVgtbcyT4RfB1MFqvm
kW9PaHGiiSzxj55iKC1/6H00BeXtBQ1jGog4TUQ5CmGgoAJYrQteRGQzYCNG5NXi
bbJOHWzYbnZ9wFwWju/FUTiLzVG+CuxWFG9C2d2cUyRbCb8uW13KR6PO+GsHfhxq
PrN7bTlM3XqeKt9iIrDk4g19XY/0vJwmM+EmdZutjCGPOBk0UVb4HwoSb5H6jIHj
97frSklDlN9F0n1jUE8CUnmoHJiTNtxLKUk0YPVGt5CcdkTeDD0rY0yMcxQ1rqo6
+6FlLro0eovMCKUlKb+KQVKpP2Y5eiHLeIMP2iil5RsKTUt1GwfvEYDd+TfifOoe
LahZKFqii9e0R8b9s1muQ2jfl31RqQE7OzGNqXJC3LVzbYEx+D4JeQIxhX7BtxOn
hy7eagKWuc2EcOv/Ql7wTMQO8ACZak1f0KTNnA+aSHakypLFgQGsm9gHwyIdxctD
j6xyZ4Yu4/u8Y9uh1qRNqdCb6bAu3nptN8JE7DHIutV3QXnpK6rnMAY7K6e70nMR
6NSk+GjkpQhCeDR/5T7enElzAS1knD6K5hrQpHhSmzzUUWoozSeiyi7meNa9hb86
zo6JKxhpVFUHLZgDUXBmVQK7jNs9+bjpSPHt0HX5dNWEqN2/Czaq2Andu7GiV+Rb
ljyASTxgo+1Hlmqnk0iP9/HCnE4SFqJmbwXOGYMiNzqpejVn0gRDpb3OQdvVUhjj
+chStbKaeawoscU4f6ls/1EEIXka91n2Mq+vc4PQbo3IVHc3jVe0yn0foueZCXu9
otekKmD0LbO25ssRdeLa//60ajnKzsQbPeRyxkiSx3QwPrHTPLodsV8XCGU0sltw
k6iR0pbre9ZgFErWcIgfGbI3OsO55h7sHrGOxUDHJH2NWR8siTL/y+UjUJga/v3Y
eXeyh2W1MaKE5YJ15UvcLz80mPAa6McXhOIsKFQL/uwiSSQz8/Jb3lQ7bcwGITfh
mbIkgqoiH2NmxDpKIn2BvEMLkts0nZnnpO+YHPGG2MgKmlH7eeL7gaH9FP5TglV8
k2erYROkFQS044uJhHKpENRjZVVUnytF79pLarLGmw6gZR30ExFxFv0TYD6Xm01w
S/nU9bPi2nlC5ZE6nVIdCX+twldIQuiEeNI0RIwSKNNenIRk+QYGW2rjiVGi9sGa
kxs3LkoCkcw76FqCP0tgBirYWagj7U34Q84yEMt/zoJxvsJlytjQJhAmksoAe2iJ
r8kjRO/uBxC5gZPzNKKSvTOeea0+Z/Z2ZBGwCB1JLJ5Pv9Z79P6s8UsHNwJ4egci
OFDxgXAmg5xg2tltpXvmqZHA22O/IO6qNwNBgCK/VZS3R9eHfKKK/vsTT8BSL7Jg
skaCXKDV5zNDPt0DM06U05zJr1+7KxIlB+9sEqBv3MYT/3ncYE++tUxem9WFs2QS
XXhVGsEELQNMFXQGrzNV2AoTTe8SJPh5YLs1Ds+2bT8DF8Z15OP0dVKVr9zCa2jn
+k86yGzZ9krRNvzT+Gnt/CrP0Wy4rn4ehymBErTEhziG9C4mA/2DZ/tAK9O2ADH4
NYaHp46z8Wvvbaz2JPVjYbwmg+UicYPmvPDxobf1D7cONDBTvGQ2Kv8bxWcvbA1/
SMhaIjev5c8sWKxJ9dL6pboRcBx2TpA6GpClKPS1lx0tWJyJJLmUpJJKDAACMzb9
zYzmNowTgCfAu/9P3/ujSjFrblMU/waQ7+vNsstV6h8dN8teYVfZZIyVV40+YdSJ
RutF6Hi5a3FZZ+qSRyOvipvWUuYAHchN7Z0VWvQ2byqy+nBE+bTRZYEHBJqgvy3L
pO9VV1wNsfgqyk1VuxiEyfM9DSPkLICs0e/GvNuafnN9Q0JR36NCdPpKro3J0qQZ
mWy8cuNqpbxQ1cWoCjzfovuUqP68Utds5QgXTRirYoUJrfAlh7o70BAId3PZBPfP
fK1nKqOSw47KuDhV12Hj+5gVu8MS6SDmH41W6FmnAE5ygynlpLwCX5LvhkCbjvdJ
Ib3IpYRICH6VBjlD+vVKaHpp22vsJhe6gONunUjte2JkaAVDwG7w1AOxXDwhgq82
TLwaeWKQ4o8RdGLlITfmELQalCI0quoM1N76o7QROSrxCm/MjJHELReQTfa+74rL
qJIkP84zoN5eOWZw8p3mGuy8IUNYr3dgu26flbJOQeWIwdEfP8eFeeJO/pWGpvqm
L2RUnWIsqjx17FEu6pxjv/U9K9icqIajTsY5D0K1YIxpZG/x94qyq24QEMy8wm/F
t32See5adSX/+vLeIPiQO4Z/Ia0DgOfeYXDEVdkSIRpDZTUpt498zlSiaue2DBVp
rtQOTRynCZ3VajLfqXOThftPbgMlpvwqwYU4ELv8YYV/IqckBOYeTads46W1g6pZ
FyEyoW0YBxQyVqY20RTbLGt+K51RtV1PSjKGEv3DWSf7hgen0z78WRl+ddZK5IKs
bo9FU2kxrJ14UuAa6UG0sESX59F+XUJQd2Yah/ly+lEm4EtVi8h2Q7RvPHfxoyev
iN2N7E0TjTVi9r+0QuEZstvdphhJ1KpFJhL2TWNav+EHLP3GMgU2nptZ43MwEoYE
CKxJNnSzjqf+ReJDDsTIeGfN8Som0bplXi/uNqNU3GjYYXTqUP5juaTbPi2Q7v60
wd+8vfFxf4fV+Om0y3SO+MBQQp/mCl/RsW73NYjmWHCxSrGEBv0tckHoPory4oZw
JZ83qY3e/MD4iPiEU8pEnoW+5gonX6WXEfssV+MPKA3CFIu5ELTyS/S6lBf1csHL
bS9JBJ2xRWvOSJCiAICLHLPf0OxIrAqybYdh+soCgj6ABgvDJdBs1BuZG4hfgMlk
0fKAPdrGIPmOqxdEDFd5XxP4icg5lk3m05qpFg/6w6F2aHk9YYJECJWZeFGpC5Ri
v5DNmpmKAbmV25w7dFR5r+KEpz737uvYkgSJYdN48bCPEeQbKK6o4xitv/s+aZc5
pE/BWEESOR5H2E1EwcNfGdj/VeegeYMq+U53eBBzjDSBk3H9m8a0QR2CvzK/yD52
R8pTYNnm9Q6qA2XbnCaVhhU4PFNvFXjoENEqOtX8oa9bYl1YRgyclT6Olt8HGNjd
rvngd+veMRfQZz7WjyKy6khjBeRcq6MdYs5HFIEtVQ9SRvoH1zbXCLAfOSyHUor+
1bKO+1tsupaDtzX8q+J8OXYf1n6S4e7AXByf/nPKOcwipu2LiMGXaMW9r5G7IznH
vgBCZ7wgC8UJNkvHEkV9MDDGu/wKSgAxs8QkZ/217IoDH5XCHhTAXvdbAcd4l/ME
zPGd+Mln1Twqgo3WK7HxpMsRBwqlKXDvgqzLcNCZlMJANMYY9R99OPz9z5uOXzOs
xrOtsmrAAXkelbNUTcCwh1kpc8jolrIWyB1CCCUozTQf+a28TJzAMg4/KkNJv233
YA837TVZeanW5jNvPLKG+yOWc4UzPqaqxt7/NTZA+/l9R8Zf+ES7ZplEbvidEwsd
nplA1HJ71MGcY50HWcdnHroBA3qhKPqJ+P6GyP68c1auoewHURuchv4Nbp9EZDpT
3zIJLM4m4Zneu0S/WhtSILd8wpQCM6j4Oh1YbA74YYUgZA1Grgf0FVqwPJCXpNb5
60ou/6m+KLWsxZ2fV4NBw1z6Ud/J+Dt5mqaKZCfdVPKtYi/2z8CQBw98Yx6gBDUD
6zYWCUiAXDjkYuf97cN1krnjCJ0JDf7qZlQs4pVNZKvZs5IuAjQaInGpLcvtmccG
bPXUkzgtI+AEWFAxQPphHG9R5f2mAE7HyeeFbATbh2CTETY1AfRl0KtqJ5BkE5T4
xdNKuY4BEpelZRk05y5NzSOH1gR5LCCPDODeLS7PcOjRiko6P8uW/gnT+xFr89Lf
IGwrroDH5GhJYN7attEPDRbE31Q8Vy5Wx6vQMZPbB/Jcu2fTsdwxCzjwRNveGpYU
U4I0FT7u1B2bG33Rjl0yp1gUKIH5VOxQyIoHtw2elLEorAmcEQaMckGgD3Wmbw8U
0mQTfRZxYMADiIn7b1n2QSNmolxyabz4q7LsBEn7yievMLl3BJfQQggpUFmKWVOn
AbAql2eBlJurJm0/eVmbTPoq6lqELeZPQp9oepkewInM7Q0W4rX2LhWnOmry5zlA
/oLrEkytjZtweLLCI3SnohyzisKio3IfBk548E6TrcY/k2ZJCLVsxmSVc/TTyhjX
IrOJnfx+UGUaP4KpdKsey+tt/9/k35tIOTwKYqtzF0lCt81M1O06/p9cwC0E6Hb3
L2LBrn+dTR6tEMF0tc07K1IOvoSY0vI5UijkR2s+RGxNsWcw7vlqc5OMxCsV3dM+
fYQA0IWwWo88kJ1SOGKrVs4Z59WrUy0Vy3V0GIevsTsGnKNmjNE/WYZVkwpZy7Gi
5CynbjYdYss+9g4MOcVwGX800ijanoDU+V4bRvsohOJLIE8W149UCSRWDVUxh6xz
H4Zz8wsOsiKvyHIDXE4rlEoMncbaRravFaJy+xalW3ebrOPQfEX7tUF32wouJ/Pp
q+AcxwFTnZHjgORTDXLfAKt9hpg4s5/7cS8R7SKDAAxg7qfPVtMlHcNzniy+T7/A
7pnKlqSmxTuRqeAKWqdr0OCKqyZt9YLx0B9qNM1Tv9H6Vk7kgpjC7cDVX0sih9d3
Z0i5HiIco5b9c6W39Ezsa6flyrg3hXMs40qDLjDtDmzvosqjwLPC9iR6He1QmUPt
wfrQwQHikTq7UWbo41/Y+bctpNtCoyfjLOFjCpV3bFqKo7jb/hX3sDoIZkMQbx0Z
ZGRv4lMDJEb1P7wOo555tGjJ0Ed8fiPJejbqfp3nPP2fEk6MvZHKlzx/Je07MpF4
oFhdtjvjaf6yjApBf3RpA66LCuw8XL7oWrA7GKmr4zJ1x/SBe8pKLmkL3cg951iX
HOHXhnnvsOOy+2vXqjSD5CwG6FYcKXMnZkEsxn8MhuUKwpvAD2ZlNMZdDnw9CdVz
gYWryCNudUD3f7UbzmiScEI0VZPH7lmpT6rdZ/UTc/GnEh3bcCFnRwpEZekJfGcl
NNE4SyJ8XbVwcYL5LVrmJyr9J3g7kZh0JAaWEFQ/rjXyrNziJqZI9THyIt2jpn4K
+fMtIUX4dPPjRtbzHFmkQa3ie5I0w3248UgH81BUrod+F6D4kpzuot/lysMliAf7
IdQglaWAHT6epbzsXxw8+TyMLjWublHv9BBhEd/tU2VqzPnltnapPWMCNTIz5X2p
CTt5hZzmjrCbJO5fOj+IPzT/KVuAj+pnaVlIkDedSalLzyWa6Ym4ZHN+FPkOgLvC
KNeQV3Bo7nGE8vCyvDUZm+I0Z8z7EcpillpIq4JAO+G1sra1k4AaQTOLv1mTLsOg
yOOejFpNczLGkdhfRR0iQknQAhgk6HqMaTiwfk/x8OuHEIuU468LRUYgEEKG3j95
PQ0rnomCQM5On0d5knX9q8XnJB322O2jakXJ1J7Z7OeNjJuMWJm3wtxdB+ChUDyt
HLEwvsp4l+ktcjMa7oncIkFJZbLd1aaGirfy01N6Mu8nXZedE4OpPc/wbOqhzW7L
ISsxaa2OIi2aHohVv6+vB+HocFXGkzhUM+hfIW/qBwmt6sZi4nm4SeK+M4AgvZyp
95ZQ6tcQlD4Ylu3ok4ARKb6A8Wx68IdRunryBEsAtBeY7npJ3mCZw/Hmj/VL3Coi
Aw2ReW7KhrKrroDY0qrEj3bey7pY+KzvXHpqjiteuzfatP+0qG0X+ZTVq0eer/+7
hckA006zCdSyrBPpG25zQaoWSbTB2L65astS0OEhYxZG/B86TVq+sk+ZbSTKDYjQ
zxG60u583Guo+hYONgrHZsiEmPfBj7HpLTx5OzxIivnB8ygyLggCAxKE9CmGnpAJ
Zx4p+tXuRkuxtKKR0pIWKyHuQIwssuQUOSlsFTCkTfSq3OCM9uqy6K6HD8vDNVNc
DNuaCd18jlNVIoLOC2KED4KDI88XHDiBTYaOxj8/0O8d/87dlp/MrRou9UUsOCuL
htrWYFTt1xCamRdD+eNmT5MSRK1ciPkGcagiZk6v3hdg8BT+OmIkxQKubFBbjuA+
6VLMxFwotqjWZfKjpUemKzOTpLQiPlwrBZu/f+z2jfZ5V55+d9WdgLrg3FSSeOBm
wkRZRVwt/jpix8m48fytIpKFvBVm3/gmqDnsXE+6Frux6l+yqQWfll76c2aW+UmT
0qW8bCJj6GzqAnFAeW4r1L0kQkWkF+zxWSeuhYO7ARVVYd1JgrohJJdGrv1dnjxQ
5DfpWL7Z9y+2aiiGkeCZMwZuf3xlYs6mWPIvNvDBEEF1PNED5qTZeERueyZkdLCQ
Qo32DC4KcrUnVglSDo1kIw3tFzFAimpJCTp9NFme/l4xqqhVEWEJ9jMipdLRykfy
BWurWOsWfrK+B6Vo6ZEktg7kdmOcYJekWUwmkzKD0PgWZZxP7/wT+HStM2AOPdKD
t2+JXLRtOlUpOFwdnozp6BBvwtH8UNCWiyi6BcdEBbUKWgiZjlqd7WDMvxOXhQTh
xN6NY+yISQtF8K/e+Ey0AIXOC1vFnlQKI2vDThKriEfZpUpIW46s0hCEC1bzVRzL
48R5obk4Us/256nPxatXfrGrRX8xpTXaWci+JAuWCiNS8EpZH8kLnXu9d/iJl5sd
F4Gp/UmluHyTro/puS7q2Khmit9QOnQb4S6ut701Ai4v8ePaR3Ik5yl8A+cJVHIB
LwAA1gGO85Wrp1ZPT4MVxQFEAfUXH4qPdXGo+FFesGA4IV8i1tyBWLYoj7GP/D1o
dPi6TPDUZVygNXQBmufg6ecLH2zUg8LVaw22i5zHi8yLgZiL7d4fRhzTTO7IEuyf
D7LsGuFCUGVH/UhaVy80PebMj5EDa7bHg5+dwo72dU8APbcMsSsoEuqhgYR6Wq0n
TZJy8/gCX9Q8N3AEJ5e464GcZxfhb/0O/ERabK6HOnp+8f7qhJNyKxokfZSEQY7p
8N1vz+frEpyw3e1E9hof9TQuzaC4Ei+SWYz0OhstY/qIF+kYvjShjgNxcJiWt4U0
VFYKuDFb75exgXVxFTMAAcHXAoHpR35hTPma3Ha2WLeqPvl+eA3f349bqJ0NIVWu
07PEoohnAvuLGxC8Z1JyMQ6gEYRI13GIWk/6E+oZ8RPxReSdvt3gzxVq5CKuLqZq
QASNe87bxZTJbyk0Jr+guey1jftGnaHMXa4fC8xvY1uaXwM3tIv5aJD4ctFSnJgm
m+KpookoK/OIOGEr871ntI9Etf1pa8XsZMS8b0f9zzYn0V0EnIDJHNAwKtJN3osC
P2G94RjdwEIPTslSjBuEmJn0oUVf4vsGMJ1hPNjmxLS5M1llxuSuMdEYSOdwZ+Er
CNBan/xhNGh10cyf7fqkq9KQb2U9HyV+4lJepUpQ0kLXR6m855C4vpP7dgehyCcc
rNKkMYqwk/O/ujW0D+KaG+TOICS/OV5kKw4oCzhO0ldPTri8X3Qj/uUBvE1cqSzC
ADP+LRXLg4gzjf8ZEtdMMs4xWSlb47gh7Lr1wQXQyaqbmRhsD0356tl2QA/SWhAb
YJwsyBe7aiQ5FCBPWJpn3y1+D4NcrMrQdJ7JPikNiXDV27qYml+4fKazlL5o+pYa
LwMyWHGGkGx36c7SCttoHPsiuCVF+ZsC2QpwraXbDuRqTGF1CSoQX2wNoOV6phkV
fEMY7yypx7O7b8f35xZPWpB5yBHbK7tSYbtEV9T8RnVg133r9IUNxPn3oeO0Bz15
K+xfw8XQYptB7czEaIhXlb6cuGmQItl/TM1LC/GV1+3OZa5Lg/IRBg/uzN8N5tO9
dBf9RB46a02kbZhtKx7612rQX4Gvwe1SV6PU6TuDConmOHNmqtoCY6BZKEB2exq2
1dpn6sZXRZiokZM0FI+I8LHIAaLwZwCXykmO1//EeF8fn/7n/1zmLbqxt5V+X+Zj
E736sjUp3oE1OMm/f0PZkDsHHezoAA8sFT8f8Ozvwl9Uo5FvVZd3oMfTOSxY9Opa
LCYe3mYRZvFnpbK5spuSxXNaauA1htrHXjslVRUcAdEO5WygwPfzR8wfM4EcNFgW
ZH7ICsRSv5TtVttAcfe0Pd003RLyupkiMcLVR2aw5XXkfcOqvQR8+y9ucEraEh7G
lWSYbgGAWxS/+XbDkaKwYRfVQOdhXjnLzLZJklWqhqxm+VEdIjo89c4z78wdQkzU
+7f0S4ZtWA31yLxWlZPm4nhJ4GxN+t4mZO7LpDPglwpmlbHpFplE2Coktuv69+vz
pyEqBQxGTdcTTkA7s02w6G4m89TcMm6D9V00U2DYy1D9VEEe+81s67xfA6JvBxaM
5IgbcGr2yEHl8pxOmmovSg9F5A8PzlZTU3Rvzj/O5rP1SdrktxAYMXEL1+mWwL1u
smqtz2DZKLrbTWLiIU6xcWamW343yak910H3R1XYIEJJVDM7tkF0egAT1H/t54ix
IlVScSNxQSFBzsohI11awyEfI7g4md+CQe/vpM/k4w9fRJLmVuSOagWN/CpjnI16
U6jJmmWoguXVaUHs247Uh3Hz5+5JjDbRNJlboJj+cwqJwCH4XdxsMOdmbo2U7L2V
LjESWWHLt/6S9Jsz8GETmlu1YjJPJ3mNbRVm/xLTdFRlkzwB620DFBj+Pkc6yk9I
C9VPBURE5YjY+DxeFdWp8DjAZlFG11Ie+SaWOAZPfx6eLlZX/6L53pahZTqXRz4t
P936H0FWHtR0aBssf2LfzWPlgi+DPAFPL1PUxfo/4peqR3DOLMzeYz307FuHvlRz
6K1a6ro+Gmny076wn9OhchbXY+eHDWGI9u9B2uzsdCBsOgsxKe7kQ3714d64lfno
KnOtKBiF14scVpwg/mtpoJv3j/D9AvyOfBEciq4slXj5lza/oGH6u1zx2eRTkmDe
FjjhuTn2E/V2qTHi5Ob8z77DWmUGWXeHmKoSH1sY4OKddp0uN+KLV3SPG2Qq9tYI
DWXMvk0D81fperyQYFDtsTIUxJum3XjPCDJVcA0I5/Lfhy1cJjqtkXhzqwbn4DW8
8kbwdHxekxcHKzyPQpf053K6R6n6VYZlzU4iTV1u86gFp+Yavf/3H6yD7PC9BYpL
JVz5e6KFPXc5c1VtIyN21NT4LiViq0VMDrlseloIGrHpOGRftx1vnQm1sazVjNy0
GgCTroURZ5HcdNscz3MlQhZH06Q7kYeC0LoAhnN/q8W5PjABmlCgQkHdbHYf/JBr
seEpXGmEuRiRd4fjSaxIN0W8ZkceAVFvHeUB3BfqgOf8bGRvM73pgqliIOpn90gM
1QtAIEMuouE29/Hj5/dEyloPgqAxSw3h+qpPrwLS4bV2EDof672eeNsBGCL5Ikxm
hBZ1xnMX+745ZIIGhrtoh3lKXUTZJ+DNny25BIQ99iyvb/jCD6ZrhFoZG/y9A9Ou
z8y58Hvng1KygLgBQz76XjEUAGa/iWcXAnHCFITvOf1gTVU4Tr86RwVLhIt7fVAV
vZ0vEwrK1lyHX2r4m2fIJpPZLRKhn/YRJceaNW/8f7vG+6k1e+BctUahew/5SGni
TFOw1mxL95/Zh+CS3TLe8FsrpsshMUkcrB/i2tB2E06eRp47JTf2u+l/VFpN2HHH
CLuC1InkZv+b7O7a1vvoJZzPncZtAqCbuMgh0+fX/yBbVJ9dSD1gvQRUo37rX7yl
qOU3qtgpCuKzZ7Aro5sOGyMbr0sD1JOLDCDbNp4IjBHvw+cVO9FtjsNkPIB4v/30
Nh/bIHP9JZHSwxAUUm01ONTaWnAoJmz3lESifrNaYuBB7Sg6Bk2yUMYdCLqsxBO1
BWKin7Sv+PeDOGSO+5LakeVGISew+be5JfQjtIM3PNroUVNdG300MUdSCXEZy+fA
GckXEkRdPsKlN0i9HWZv6eIB2YEkvrU84+2DaQjmSpSrBi6VHJB3i7giE6KgUcUE
708vUVd2DY9ynPLp/BHK52hoRrCoWz65WFEsMtDhz2Jznoq0J+wpwB0xvqieLo8b
W/k0BZt35odq4AWVHQvn6nRZb7aOb3gRINPfROzBq14jCiRaD/ZqhK4iVbowuLqF
8cikABdysJLDYUHQrQlO55JqMOd2jMTzqTSMLrfdY1+HsaXprki+ETKU0M2pTwtE
Pka6lJyLGn7t5sksSsgtUGJtWbMyr2f9HMdRvDUdD60xwRtrOfz0j1GveqxmhOUY
LcljGqF1XtSrWcVXHvohySXpSmTFFkKuPkpsI5UqKtLhZ06YMUz0O1YofzG7uuMM
AYajCsI1CbUlInn/LNLz9e7TeoUNx6bDUUGATZV9gPDidvE98CCbCsGPJrqsEctx
dzJnrad1XsA5i6ArLHbSiBOjtNCLPyiZH22Smdo+ck/azzwabuSIiF0o0xDKCki0
GyURseS+QZapGnN0Y79zpIf6wWv6ksC5o6IWOSLgb6XoUZLdNNaac4/5QD7ts4EB
nyCxvWRctE3K8LdiOZLXBja+MEZVBpI/XeKAdNnvfMGupFszBXHQxQjogeVEeddu
EdFnLrT3fLnVgzcSGMC+X0mcgSgYdGFdTQVoR3sX/n4zrpG6BSjdJLHUeb1CIBBk
sNKUudOEE+oluVt3m+sKsgL+Qbd52NUYB2SPOsPj5LBzPaVd2YyEhfEUlIko6gjc
ltKiw+3WhFFUZA4PwnqiNb9lFso93JqV5msT+iw0M6+/6aW3ZWECefnH85cZ2goV
YY0zwh5GJlMiv1BftSnv5AguBT95pdH95XLdOD0a4RD0R9kpbJ+Wr/sHrTa5WAtC
PanHbLoRc7mskAeL5WrZkd3MwPkv5ZXrn2yD++2LsmfMmFiyPSvkO9mUei9wlZ74
0uOxNWBoScOWJbVfxMZ2pPe+XJ/dopxUOc3hpmWglzumQen8kd9KM5o1PSRvfOk5
hf7/fRIwSYquCXLERKnoRJXQWuWqae/EXAF5DGfiRwxnPVve37QveYPKwaHfY7RQ
Ko/u+weDqwsBtvIehYSlcfw5SZZ7ROznA0Rc3t7eSKyOp84o+bnO1of71cNgeZvH
+vrUIP4yWsFxSjGObj32oW01R0kVOSG5Caq6pygzYEiO+3Dl7eEsOBmNjX6edjzW
Z93PSBwPdN84rzRY4ikE3hSj6FWOnFFKg4WOMDcTeRwvYvycdFI2lXizMN3LI8Cc
FCTQmSDHJeq6Hs+0Gm5LwCmPA+z+WQon+tmPbOhp/smZC/u02ZCIajBbcTu/mwkP
7AnRODO7OYvQmcGa1hT8RVVqFHqaBsqDmM1ux25i2gnTr0FZ4yHe25l6AYFWtjjN
4ziOzWWw3XJD52oN+a6hq/BWh4FGGT+fPlYUb4fCdpaIqu4ZvfTWbGZVSlShCUYz
8hiwqstqs/phBhMCuJ2PXTki3EuwLGYBjd4m3O8nFvOIA+epRgLcFwgSQD30pWok
DZ23Lwu6lMshnAzZlq8YwqD3i9Zsrmy/FdivAkyvfMc3JTZYLdgy5hyfFIrqh23e
2HH1OHMi3A6i5IyWwOOKDXMSBOeEP3mrfAkWlQG+TXVnRqU5LdlZj4qACiibsp1+
sZFJCzxsYYdxCxoMgo6DP4ysU4JhLqvMAsDAb2oUSIbMBUpOFfsY8btoIWO7VFOT
L+2bFEP0nUCbEniBtBC8Cz7Vju+SUl5YvXwnsVrZeiBKZrlpo7jZ3bQ8/hptRZei
InFwK4EZW1oysTgtFrFC1k4YE+kxBnBWcY0SIZ00WKrZCHZTp77PpnOVwGfnbcxY
HXkaIKesUfPsIoICIf06hnIBe90fRp9IxeJJc7TnzUjCZsLMmQAQ2m58ZQi2rcHt
o2TlwRvXEM+fGqPraHdS6AxvRdbrnxGVNPZAF1qPgaFQZeW8T348AJKEGWB3mtg6
SjCW+dsqsg7mC6FnQTvTv0aqQqyMk7ZOAjTzLtPNIrjB/L7WKqNVaVDDDBqzJgpd
qHALLAqobTjJ/+xZrZSejyo38EotHKcyTE916x9wgRbRC4Q4OscfLCilHFJdxMDZ
L4efls8OjDZgzsJ5jDPIS5ICrTeTz2/bAKjQQwQbd8Z9MoeE/r68iDm99UChV9K/
F79hy37dHvAjfOburpsG1xpeik1eJILnb+EFg+N//VXUHvIiVqFcsrriCvfy0OtX
wHGiUABzPd6tYyeJPiK2EraJvm3nqW2RvIT420MA52OOVAPVeMlQF1DeTvZRFPeT
JqB4HY8bc7RLhronIV0YWkdXCRZ2LM/yUgcgMigSS3HtPyebftVUBoFhsj8Aiahl
YhLlvF6eg65dciR6wI2bVWZLcqYH/n59Gw2QBEY3fm2Q25Krdl9Nfeh4ya4b3N0W
TVySqBr5L+98p3JDKtZnCYw4QfI5QRmP7HP7ksw3TSeToKB1cVojmk/MrpevHROZ
vJP35bet/h6hPlxC6mCmNQj+0fkHUIhC1spOsJzFWjbCTBrz68Gvtp2ZkhAYKDQ9
wKkwi6Yy5cfSqZrKZPZqaB8SjTtsht0RG7GBYgyfJjcJAaL4P/+PmQwNFiHxzm8D
JkHKHRGvF4XNpTp60HnEjrPi0yQNntBtSUhLp3AQhBOjFDJwqMXLlqXQA2P7LuaO
WSuWaeqfrsKScrgq+fYn9nClm7/NE+Q54uVlXm/7v3beLH3vb8VbZGTz0CPyYU72
SWu5lHdBUByizdwBnakfiwfISExgUCuwPb+kPzoqU/kZh3XLit4vQHuGW29McUza
PoYZk4kSWyNIq4sEnx4jJhnZ1Z/+g3YCOWdUR26m+1RA54UgEBBWaEshYcp7ak1P
foVE8ntgtXZ4pk7q84KWETLK9bcWD8h84P1yRkwNa4AInaAfpyRVSn3J42uv2UkU
/9kC99p6vPl3WZ5ZJ2ZE5+13G4gXCs0MwDHxsNlNHqeCyx5h4+q8QlSdXLO8/887
wzuntStuPErfiLJUkhvd+3Uvd7GHmAQxSV7Qe4F9NJ3ppB+qW3pMqaA/+biLJDMd
sfYWznTKL9r5FCSKcsBG9VCp514YSJRozixO/aAq/9gSSl8/65nsVAXJeFrwuQE3
FLLR9aRoYFdgABn4sGGH9wlR0YZeA8PKWwkidLhMkIR6zzghGyeV1i/vnHhOiDRm
F1NWiWC+8wY2j7FE+bBKcM065g0TRtts7UsJYPftWSCZc3RXnIUpbx4czlv4+1i4
DEKjEVn3Fp0ZdrN2FP+tEnmSl5K9IzQlv2AKll4A274edeaU6g2tWHH4K5jm3mkl
fD3/tQCK8YBLEnvnMauLRHU0amv4382o5yticPtSLg+tY5CmPW2lOmA3serpvIpc
rgjZYSl3QfIrr3S142FbQAvX7DdGJwGGPcXQklfJUxAY+uYIDacYJ4/arJSMqA2l
fykPFkY6WvPZvC0Y0kg2kPTCdiAdzf6WVwm2PlMLysUl70L9C3h08W0zCVr7G6U2
s5qrqnBN806cHBk6aOarKijJB5pr0veBwoh/WrqntjeMoSD6IQt63RIHn+cpt35o
AopHesLnhZrEH/D3lAaJMisiaRnhHHjIJPyHNhkZfT1lqKm0mS+bDUfmWIrlqj6/
ehZsJsqhwuwxNJoQajpjBw7Q2a/Rn+SEg5mpKFQFUQg9yVAotYDhq88TjVjOhbNa
TKcCSZ3wsAYdEInY4ouWi6obNBIz2G/dof6TEy15wWXe69tM91EwzDOnCdSevSZ6
j05dwp+oHT2ElsVN97IBQICbECtlqx0elc6HuCtG+NruAI9OIbx1hFFO/lsNFI43
bRcoEyMNAmZd464FYE+uLBypT/VvhkYA6TYlsAjOW0TjLa+gNpaZ8B9KT6s08YKP
JJA+WCNNvx0qt3TJDiP6nM8p2NRNRaCUVuJqx7VLiEz5sYaRQgG+KV1cV2I0xSRv
EWpueYQBBi2mOjd7jxxysnYaFQJLnv8uRKSo4Dxn/i5U6FIIJluJ3t10qYyWy25H
MglehZqYqphYw5aeLueZYzhEos0TBgevVtysf1wh+r1szc0Dk+0l1c8Sb24JMtJ5
SWtxfTHTopjwg7skaNlx5Kn7CpP9l5LiMLgEwVIPX/j4sql8+S5w308sUJWANUuJ
TG4b5JwD26KWcwtr+17lnBTyOQAd4zU6ZgDeFRNeJULUJ2D2GteT8HIJey5g76N3
sWgLcNAm1AJTCHGB0FYJBLb9dvzuvP45BNxKQf0+6Zu0yGMui7agDr1pG/nkezNQ
1xi8BKgN5v18CBZD4mN31dEbNt62//SIEOjKK0m9vwUDeLh+Bx0pyCSDq1Cixd7i
LFz80qgtcneswtHK7DHNI3oWjaMb4lIZkgBJHCbzggWuKR5VovrkGaiAUtb8GJXW
OFl0t14+UKvfmslhulBhse3HNzvwy0BF5khSMFmKf25DvsLa+mLSESWuAYm1v4rh
bJAWyCvJcrTCs0qKPz1ZcvXvhs+mTCOIKD4VSz3MCoNTHCB/JV3buLE08kj0YMgj
5VPbAnGTmCFDNwa6W08NAGJtsKFEmKmzTRWtOLD8Be2vV1B8VSDmZ8ZxJ2DoZDKk
x25TbvVOVTriwNsV/U/67wplPfgi+vY38dAbFksHboC6HOyERIfGFA2GNwfMW0Ql
25a3Nsip0yJ77ZzSnldq2dWP5aYuuHcBZ+OUD70R2DIEuv1GBCunSxLXb+T01BM6
lT8jy5LL9qHk38zwANTNKX113FQU6wL9G/mI6N6HEYTxjFf0T/C0C3ZzVObsiqc3
3UPccVZER10/mApZf3zMbXpaISUlRqL9jDhazntTLGBSTDqyqh1FI2rlVs2fTFhr
CNRzMCOUgSfB9HMHPfKGB4BBibIhrt1Fw3mfN6x1DitKudi/opqx0I0wMdsqblpP
Upox3k5hKuZZDPSRGhpk59Jc42O6fUXuU5FdpFGSRax/p5es8dKLIbSB8/pqXSmt
84cqCFxTQ5241dHim4d4i7vyAEY9+d13wSQ+vQZjI/7LEjvrVbxqF1QSytc6ablq
S8F7WQRhjC/YwA6CmwSVdx8kgcfaavbj3TGqNHA0zUJNdJyazk9KTO2u1yxiFnEF
Bdj99QwRiIq3Qdc7hdEiY5ptnlY+sJkpWqexOhwm91r9p6fiUKlQBIPrYmVCRINo
ccdE+q4DE1JbDWcOAJNg/mbp3csiwb2bZ/dl86d0Gzv/agyHTEZtkc7oIGagoqF1
vriHFVsb17K5e1uQxsV8lWgOy9buduWZ/DIegY9OLamMGUOp+nuk73NYZxxxHY1v
EQoo+8tLhTjna5MZO6tn85rx90hrQIhYPlBnPSJ2F+Nj4D3nqR6yqizIqQevBi5Z
2qORegaZqTHOKinwNKKQdN7xs7bNwHfQwRw8kxo63vNKhJUDzSARXQbt7ZZso/DE
pxHF7Mjl4vtjyqhFeRFSuGgJRq/Q7nipOMOOAPx40tZ5uALwMaoepFBW0Yc1NCaF
JAw5bHMWDXw352MUBZbbHMjGpZ/EgVgQrM/Ju0FAxxUbcwTNgPg9eiDXElpuKDRA
debGTdPQVcr68nyjjXwydpRvRS4u00Ie+CqM2Ze4U1AYcCh44nc/uAMU0UuEKdLF
Cqb6JpQ4mwfqyVkxynSE68BTak/2WYTAiXMSv1d2+5eIMijM+KvJT5K8JSBF1KiT
AYcuUnN/JWiqGd0L1u4LQz8LtQHNiO6+FwJ6Ko9K2H8Hbi2bzrO+4JaFqA2Ka72Z
bUuPYQgfa2o2K5wEBGDZNPyRFtib0GXH9xXc1/LejJ0ERFLyLLTPIj77/TNCnDdG
3eTOqxboBo04YHvlfjw8vji88ODuxQAHPbvH2Y0wKsnoX8eg+6IZeizY/VF6TM4+
EPohR9N+QY1QbAM3p4DVj7fnFVkWMmMGEizmkDWWCqGOsCwtKQMOc9Zz+VDT8nto
uJ7khrDEeDjfSXjwUfIEv1DqMMYZJ76T8yFewfs3V6UXYdZmrd2U/9Myq1CIZa3j
+IJ0GZOi2eLunBMq9ytq+b06Zw7Y4zRSSFm8gpfk/1Ht5TXSUGAI/PioKA0ESNNv
u2Znl4lLRM5B3zewd9S+HhNmwsjsgB0yBzaH/2HxGOrkNi4hHk/IlV1KWRqRbfFG
zLdRSbmBGlDR5RPJNL8+uoIDwApQvwRMhYoKYhKTh0FvW8vMrKu1DrdG46iupE1c
vh/Y+B3spMDK9xq82EiqMTnqTqCOjqUIr6DyUO2VZavlWRQfXMN1rxh1Bly5WhNT
G1phb4wSICDIaToIjDRRU8B8DKQdw4yKc2IFMxjSybo+dOPKOH1HuZ2bIiCDy56A
BIiSb26F78dApDxsOSr19xsSRkAFMXCFfOcb0UE+Jp0pRJV1AkjtIexeOhZcturH
in5l4lBsSsSwJADMnUTeRwX7fRo6sJYD3da9Mlj3Zud1+OHhTrYdEJWT82fAlWmT
a3xA5i9fp+Wnlo7J2NcEjhgNt3+shYXh5buTrdNiaTXvUjMyBfiYgTEzLFnrtA9j
jgV9yyA4hd7eGMJ/b/NqRqiipE/u5Af/xiDcjeRTByrE8UeH8u+jMZGm6CIVKeM0
qgCBvL3TSSISnwdUm8MJKEP/ue+u4/lHRym31zxGKbN+09VwDLTlx944f5Z6t+lD
5PxvvVqOwWm0lS+BjK0KeMqkdps45n6owTOB5RdwMT7vlrRUqApnKRJfZp//M14K
W9iHgZ1erG/9BkCAnVnsQqIXYFueHvJaYgIJKrZEF9Q0WIEMwWnrWfm7lcQaJOy8
l5M7wSDBZRLm+I8znB/t//r02+TAMga/oe6lW8yjp9o2aaNMv9aO+a0WMVXPEjya
Mu33Tz1a7HA7lqZdp6KuSqZowFrQULRqRSh5FEIHBemuR9MGuQCR0qsZqbBAZY7l
kjg79AeGFmLXB1je2640FYpgBFQNvMhDKJsTLiZYuX1y4WETa/EkTq3FqTBSnBwV
2E8SwyYW/iwZrOJg/RQIJIEysHA7PX1exS8MK97AnJXGebL5xjKFD1IIqYOOFOyC
ju6Eh7U7CqKaxw3hBUDVnupW9WUf8GhZjHma6VHC81tqH9+1p6Y5ynKQ9y4sJ5IL
oOR0Ybw70TwacQUV7UHqy0gGQ0yq2WxRJMuNFWrGAWr5HOqZpOwrc1WzJG9H0zU1
tB5ZI+Xo8QurZKPQLHMH07DL9fi1ZYzyoVEGHJgoWB9se1kF7VRhEgd7SlpP2NPY
OhkZ1RhsZIMSzkBrz9ypaIVTvNK1xwhNVFmKKDDlRfeeUJq7KSjyMmw6o9/ZuvzZ
4WHWwvQCJkAXmD876bJgahtYJP7E95qYksu2Z7P71q4ym4P1FW1eOoFbc2fkuwZk
v8VFPJWdIOCjn7NBuHu/pHUWVoSsMHwuPrqMZGAp0nVnAQw4OBYRVOA5I3srf6xQ
c4FKCtwCC/yBae1fpVF+elC1taPYrjqaIZ5Sqx82cmb8JY4ZvShr8oJs419pKcnF
7BIP7wy7RliVhvjX/EBXJeb5oKnQfnuYMntWk02t3eRliyJtH0y/KmkIH2iT9rGS
c9EoGgs8LhY136lOB95g2Y5pQV3krdNxMoLERRcd+G4SvHOrgWdgQ4O0zI9XFdO9
bl1/oilrVpVvOyZI+3W9JiMtBQaQi60tUfYmyUhlVI6UEgEGg/NrRavIw0a4KHH9
ub/vET3oBprob82a9DMr29/VmC9FNgd1exJFlZSSmB0D+a7/Rb22wqtcmDVd+usp
mkemhL5zzl3/uO8rcpYqLU+p//I9ZzkkFnh1eRAyhT8wM9Rr2+nxwGxGFL28u9Gp
f6wyPRFT69v8FUBwBmoXptbiwEgawBr8hYq9jqp/vqSli+gY+VrDyBY7VHIcBPyf
woH7dEp5oWIzVI8zv8rbtowLPvqsEwPocLI4j0L5UnSkp2+/YYZKS7TqUzdrj+RQ
yOD70LafP13TmPIUzSuaMMysQJ/xC7sgb2/y2kFUgWsPZ2UKziMVe7yKOW7uSb0R
Y8kOGTX9SE50VMbQPv9su8TsYVxHJ0nkSc9pCH8lwuq1Ei7DVyCJYSJst1xnbl6z
xLHiL2m4H2g5OSaQK2JW7ANm4wwRz7dtDVOmOMhMM66G2XaBuNf47CQUDNL+yrzg
2sSHm0hueXHuWDbFrC7f76H7JXydJZUx15hvOKWDYCwqGKPVqvyNnGQM4sS9xeH0
OqVLK9fpiMTcurq6JXBDuYu2TqAnxTvg35dtl/YyD21Oukao2D/5uMmAcnJZlRXf
TEm/LdE8wQF7SmHkoAOBLJ6Lm0Dcycuavw4sYzJPQBV/woV86fb4Z5RhCAIyL6xi
DHJYW28ACoPjPaYvbtiZkyYr+pgnCyEeS4K7A6T1DgE46P2Vf0fn54JvNX+2RA/h
vvccoDFfFq2gufmd5pChluDH5ygahs9bWMBmIm3cet5xlcz4JLMzd6IlK8E8QZwg
nA2DDIJMJmx0whp24LhEGCexZ/GEY8RPBWNOCpv6FTrPuZhyoFmc0E/X0bD+sHIx
V4pdjG/jsbVkfSQqBdFqvrloHMCzhUPEwc6Q+Ir5+NpZRaYDQ8KPW/vkL5j6V5mT
TuPVKzVhlp/E/Gk/VFOK3CvYsaJaihEnDb68ZU1yiGadCi/lSSqYQdgMhYxA227L
SSvnFTC488ZHmyrlYL1Ia3hRzbl7CT3yVncEgslvihwVeuN2MoX6CoHPfdcmzTuD
YszFcx31k9W/WjCEFdY+GQGHqAag07nzbnkFkoWsf2hPthCdc7j8KK1hJzUy7lEG
D/LkdblX8S6CX40mcY+thNyYrcwG9OI2nYymORxT7rTSnKB+wY5fm98lWyNe9FTF
gwSpCaCvP/B02UaSdukNUfPcrjsBZHukItqoKAdF30ka0e6q0WjwDVb28NiOZ2/+
3MJLcZdNGKjUteYsmeRauEtncAHS9Vr1aPqFnvDz6FQlKXy+W1C/a7OtY3AN+MlZ
03E+rJmInqccDPrqHpi3siX1btnSIRB9JaFQa2Yf0q/ag5qxF4s8S7HDCOJhnXfR
Jf4FIzS1jSH9Jmh8wxP+qR6TrTEwmU96h8RWb5aLjAicncKwt4+duvSsRb+F5svG
+CmGgTBmN3sWQm6lMoEfBicIB+Gd71dsVtp6FgxpkQAgx+fpIilBg1CfTRtbVhNO
HN3QA0zxwjXIY/vK5UF+tErjnqh2MQQYXLAhhu6oeQUPQRdAyXsXB5xbyAmDdsXr
+VKcqClTDOFVWpQSwpLS/fYg7BZmWlr4rtRq9AwLcjunjMIGrw4m8VJo4+/aLyGy
1FLXAwxQSzD6b+jk1jHpEmW+vB2n1a18GTNGUlwkiItWCc+Fd7E8DQzOqNTxqZK0
MBAlsJyxzPRzNxyiaU8wc00KfIB8O7+yAu6/MNTAgr6IOTNvxS4MDXoxuIgllirG
TpKekq0gVu1nviIfvhQsNukOjdILVQzhkPJqsMN06LATjYtfcGmVvK8m9XnymSIk
4oQAlyZimDqhgCsUZ1BSEmbKdzOkusgqdKTyEObcbQPkfatEuDVwenTAWKS9it53
gm8CD3RvuZKYfBFDXQvIWSk9hIj+8qRJltN0RwZ6oHrwYQqlKxNBXkhwMjjwpb1t
JeIf4Wb70UPySU5Oy9oJyzWNEG5ptymI9SgqizMFEQKjcYHWnrwdannnEajOM0Z0
DF51nzihlak0xhnxa2zOhNaaaNA1YBX4WKq3JKY8kOMX1uN/BEPSAhyd2ywNBvaW
t3sM7XHZFE556UReoiB0V6rpuAfO9nfp5brFATqIaRccVbY3kykBZZyoPv8iDtFl
VUZF+l2aZdnT0e7cn9X3XYHHSlyXTIKBfFP80TSiBHeAV2ehNev17ynd3hmRXlyU
oqaju3gOXT7m5lqaHYV/U3wjxBVgBPq8XnMRzlNNU+PgX5+FGffcyeNvXDuDpUHI
OH5x3vUVwJFLHJGIh7+NqsM4HvmUfN30dUf3x1F4uQMk15tx6fVBKPgM9vV5//IV
7rWPnCLVr0g5iE5APPr6UBcCEW3g2slubp8WCo9iKxrV64HJsmpnlVMdY9e9m2xV
usXtH+/1KlpwJ3YE0X1etcEJ0Xqkdtp6xgliSAoS1vuLDuPFSCCa+UU+2e6wqSrk
KtZjOxrOjgxOJ5gGQ/aUmCtyU2J8ux6852mGO52dmOOZ8XTsF0o/bI5ECiPZQu0w
qdTX4uk1TPTANEWfsdSTWk8eZhl+sdENoOwJg6z/zKm8pPbL3J8JLAhHq9ErchUn
p29T+BlqLdMv6OPmBgkaEXGLn5gtYLfajSFdfgtKfY43VMKDLmECz5qlKKz9heYO
eZiHwvmAwMmBFy8ktPcLim4c7GXfw7+1QdorpT1zxe0=
`protect END_PROTECTED
