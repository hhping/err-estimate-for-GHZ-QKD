`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DkE7EcjbjYT/o+1zLsbQigD66u/EtIpuPALoTCaqYps2tr3T4JBURlNh1nkH+1vD
ous7HLW92f3J+ifSapQIAS4x8y5F7Fqi+f9YaWfjIBQwO4QBKdWZRzgxk9caQKAD
yX7hulHgYlKJQFBqQeIRi49XoCx8jLIOe6ZbmAWYfwi3/GXuPsR/SMKU/uohLIGQ
sNgO4i7MZuUeKPd1pmiuBigsvKZ7fOsMgBRxrhslsh9SLuuT2vDyl0gccY5Z64y5
zfypjD8tDuYXEmkz7zXGVtbbuv6rrF/bWk5B8agUPM7qbQp+FsMcqx5/oD3ZpYgC
SUXhpODqF8XlUlnO/SaAAwRLjBxJyL1eofnQ3hBxLsLUF4oRZ9KEvc4Lz+DoTULT
OA+KjaBtpwxAHsqp8HjGavl91Ge8DGL6DZ4yzAXCMojMXYsMemOKzgtHcPPyVhJ3
PhGsa5r4DMquVKU56lnQdg0ST1iTH5IMKmJdkLen86nykG+9ndy8ohk6jtCB/B2p
hb8fekMJ/2DzSFc9f6yh2Pgpam7eSSKzdQ+01Hye4V1a1ACOqYbjGUsFxqKxDUNR
VGZ2BHlzS0GNGc1u+JV8smxQpdRyxXneWdUq58nj1i9rWcorqoTWzESU2MPHZV+j
FKhaV1QPSbFaaxIWgXoN+zZsjkZ8NXM2jotdz/1XHgZosnfErJEmw9X2xcuazuoZ
hMez58lqW3CYWZb6FJYftT/2qL2SXwwHQW21TzaoD93Ji5H4tVTZ4VgCkotXeYxM
YRtJPZDTZx5cdJes5o/rIbV7JKltT7lFGu4NfZ4TKUuygfN0TFjPSEbK2lHhHVjC
tx0QId+MxX/o2u424DH97/fVTuIyx9Kb75GrbaYpNxlSjydHiab5n8DrYq2zbVVi
zSI5i12RNPpYxWkuX9/Yo9NllmXIW7rQTp5cEMoDKuu0A6N2oChZyguvHf7NRsrA
+lu47Vizp4ZCP96OGVBHUbvZZF8rrjOuKcrKhc7TFZ6Lpufy1u1k6wfnrUGooqwL
gc45QkxrRr6omSG7yzOj6BFHhwzaYV9V6g76QA5uBsDqPHVS0JvhAxBhxBdlEzHK
fFGbPYUbveSeYXb5gPu7bIOreBRR120lw7IMWG+1iw4z9zfIyb+RSOPpaK77wmcr
b5g0a2kjgBnXFPqFOT+S1C10yizRk4FQua2SlPvU3dm1BpuBsRlL8kR29u+lqR6K
abgM4uAXib1Uqw0LlwWFZHpBhcTA41SIVHVVEhbFHITQjSICCHjh0Y0DCNmLe5SP
saD8llSQmM7Avsag6lbckDMJwfz57q+V5OXedBsduB9iVMg+vKVDLHaG9qcfsZmh
EnynsUsLME/xtzHzSC+mILYs0mvKUhxhH9RJA4G7Biqxe7o3n3orBTW60q0Ssnzd
vVFtSSvCiqBtl9m/oxEOYxkprAtdOMZYFbVsea8pohq/bN2C5s35yCfUqPD40OJ1
WtrZoqtdl0Ci0wL+EzmnayT7dG3IAXSD5bf3pQPqLNLn+zuCDEdU1HzSON34nkFu
hZDwQkoxGT1wcDdOUq8Km9qQZoFsg9ZFRveWPsu9eu6JWB9iHI0npMFlt1jG1a/C
WjlsdLVysfh2tWxmtYb1RLUO8CLGtZUXPAK/IDpBTi8jHHP7y88XWjokHw3nr71f
wTQHPuQ/WNXrGwKEeviwND2ZukIomGNA8/0vhaHOTEERH4C7XavKOSMJgsBGmuxq
BgEEsv/xet46hwDaa53bpSm8Oax4C6eOEq5+b8olSmS65Yv7NVsJdXqWiusZvpG6
FQkRF/Nv9pC+q69EltFpYCkW0Thq/6UiUVfznTjGCIeUKoaFcWQhVzJk6NjlH2YV
BEnKXOhqSQwxyAIKPDNT3Fxn2rICe3p+ftqLQzp47tu0jH1Iw2A++c9ljOt7ZeGa
/WUdPH3hl/MSgYqCTFz8K8tELgG1fkXfyX9DdhwakIdZtwGS77WldLzKDWiRJkLF
3W3dGXi2RLQzuQZCP+6arrHHMoCG0f7Drzg1nFsEoUNj4BRFk+HkW3wifMYV/QA4
nL98cn/QF6duueXTYoAKgQHpd7Jvg7m8x4wBUjOKZdRfLM5ftWH6sgVH2O7rjdD2
/v1SbvFu5hw4QKYIxco6ZYDmgQDQpKWgJ2s5sb6tUacCMKv54F7wgli/eq35YDQl
7BLl2ybsZVlpjJK7vees05Wt9N5jm8SwFmSzU0ZWI254RppGGW9UwbAmLJEuU9fV
tL1C/VEyJLI/2/DBrY7ukkm1SPME7IEvQ34BrTymZ6AGWrV0Ko4ew357AXYept5O
U/fiKhbLbfgJJucZfa2gq2UMB5OtM2pRJ0N8Blufe5SI4cuQ330WeUFt/9PCykAd
Dcfc+zCWBrvAYTRDpicI3K5ieKr8ihQUr/P6PNULaLAqf/QMD8SmPynDlj2y68lB
WCpkn12Wd9RBe3T6/1qFHcoaMrsTNRtNBTHRn5KkzlIi7uUYr4jBCDwnpglrqEAM
1T0ao+rc/Sb3AMGe9MRBB0VF+GNxA+pKh1m21esa2Mdf6FrlnHIOvx9j3EqXdAzM
duTKeq71733bIdF8t7Vkws0vXXk9CqygYOIy15WXbAobh0vTrpEXxsXm2UNk7YlG
Md5CXEzumpMFqHDCwAm2tnpQQJraMGoCqjXQB1F6ko8k9R/1BV534pm5bfNlwKRV
c6THIYGlc3R5jJVShDFxvaKfSXfnjNsSfN8XyT5DUFlKLna46uLYiMeZF3lCO/zl
Zsad90RKNZiwmT1uPCd2QZRMbT+EARe0BnQ41YdPp70laF1k1Y46C5eyewOIX5+4
d180ht7OoriisLJOHf7t5jhEQVyOlZWNF4Vpj9IYTE7h3ImfQ8od36ar+4QqMlVu
z/G54mIoAY7zObDnPnfr48nPMLru4qJc4Evc+4QHmR1Ig4h8L0ng2h9OS3i8hYpy
d18PuVLv/xAUJu+vqVvN/FReubNur+wyaqAv38ulndhTtcMD8Uy00Y8Jwo7kZuhZ
VYLeWVdol/yyFxzRxQtm1L4TEK5lrqb8tNcRuHktcfrvuJsP2DkphrF2kEjHlCOq
E9gB8xPzWFlAmzS5LUFn3JBC1N5cg4woXBicg1g/mp3eDx4YDmW5R0Z6w7nD0F+7
A12ps4vA519SEtiteMwzAGF5HPoJAti+h9U+xLv9WtEECOV6ZH7lwPGK844wCKRe
Jsueqdg0ufpvMSWUA1rcAQRTLWwKleo5cLqc59BWga0P59Oy1U701uiuMs8Hrzgd
DuagdxmM2adtif4dJjscevpVRbxLcnEDyOmXqysCKeutrl0VmgwyrG7t85kaZsAd
7tOcoLRbOEhdncnQfJvSft/H7YDRCrzaloXz21S2ge4LcMmGs3oTxj2j3F26sLQP
GfdlY1Issf38WSAsdmU5ej12JvfOf56e9lGbDlMARhaylsuhd5RBLumuCdPi7Gyd
qUHpmPnN1/kb39UJQmhtxIsnsGe0h/08aoynRGNjJvYg/C2u/6mMD5ach8u92MHB
+6JzDR0lRM9fYfR+ZyJ0XLQh42pKYbRGwOubqCNvbC4MaO1UGklYPFNXYIJhUa2W
V4bK31mKalhcUyPaaZPjWCEP85a320GVgdys3mVJAjS0vf/Q/MRjHzt4tLv+hrFb
rX7DBVeSYxeVZN6VcKLZRFkQe6aq2tsjD81/G6VzXZsOlipjwTPejLvRWAvUBmHH
xkia8GtU9RPblvrBd2E2RNiJOhdytQMVxy7a5JIQAK5Ydmsi4mUAnsUp9hsDB1ht
061Q15TFo3DAyyuSe0eYdOn9uEqfOtDXCxaKihwJompe+KD+8ZXvOE0sMdtdHuuQ
MF5tVvIeKvQFA8cwQNCLvXI2leIZADUtpkCWwZKBKHF9tOZZMQCpXzTISeBEKMwO
+X2ub6US2C+Jm7+td+AEuu1UW8oYWpiN27OntPixGORpXBSfKOVCgdHPcMDSo9Ht
nvQ5bPtXKmEBPJAf4K2RoFcaHUPX2l9fwKW97Vavuj5qMHcdQ0KXCUoWfwmgokb1
QvXyR3ny4/JWFpVK1UA58dzcy9Q0lTbKve9gtL3BG5CCrzncrePeHUMJQdazpN8s
2B3vOalzoc7WH2sYJB4KO2oSvHSfByc8RrlzDH6uS8vXFdJMXypVZZMU7nkfs/DK
f01DgzOfNDW1vvzdRzpryMFSEscuFbVBfTDbHZc2k4MiJCZF7MRjNI3OIdnYc6Em
NHpuke5DutkIpDyXdCq84wO3J6qfDyPYRRkoLet5pAnGtQ17wGqT9vLu30wk2U3q
58BkAiIprPDUX0WyJseApf8WXGhNIZN4d0I1raTNLXLi9exNqc0QauUHbe8me/uE
HX0TCdUe0cHe2UMJbYqG+GDs1dO05HhgUoxORPDwwNuxS9pIeNY9ylbcm/pzKpYh
6Myk4dIrRFbWemhK+9rPbzNgQrXe8zpnezT9TxKlln50XP9YIKKc4yIuzhKCZXZL
h4KmR6+TmgZXnHVvTxYKyuPC9GyZmXq+4o3dPhrXWQCSWU/GJkAgf41Z/ggeMBTx
KPc02O13XtO8nsk5ZCQLsOKr/fbGmTjWlL0enFge1NOpejY2VqjeJi0xp6KhTKAh
2GC5R9gHqpAmhwsAUNUFeTKdLDhuuXRGZuHCYHGHyTkRVzt2vP5D9jcHfWoBXrnj
G0dR8PKLnU9+6A7miRasVBj5xmELvgJTlM4dfrzKaA0/wPZ8GAJCNyoFbc8Z66wr
8AY0kplL51/RmLOSeNLDN8gl/28b+xg7eiizNccm5jBmHg6pen7uJA+l48trLnsr
6wbse0WoVURuHaawtuvqUSU8u0+iUCZJoKeYI3o48PADshQ/Kx21BLmBr0GVOuex
vO1C3nYKZsrHE29sodopN2cdRK8gEsRaqDMbnFYDtfDqYC89P9lvR8oQMr3PUjoe
gAfvEd6cvsvhfln4QI2gBY/dax6KJoMw3cxu6noowvw+EiwFywIPm5BDDEMrY74v
zUJ47aLkAvnQmsh7qOnItlK77quDnXA3s0QqkG3AYHlQXOv8IB/ss5mP881gQVb2
GTsQA0tVIPIMIBL9aTuA40olqPiFg4SJ1Ixcm9JlOFk+lTC5oaMLr3lD9uEXCids
LXOrkX3uE9XSv0VZB/nE1vGysMHjfrtSsTMJJOcWyYx9Z7P7r/T8BuslBf4T+J7p
k1KkoipxX7CNM45+IQXA6a4iaPwxEpXT1KLxp9myAwylpF2Xkv7RWtpdvfZBdcj+
meiog6CInOHMMUStSzUp8MRxdwiHjR2zyZA68hi7wRQccRJELwtXv2BFgsKYtTWE
Oqc3D6iNTrptT266X7vaQ6cNCogEHY8ErfVUpNqOe6eFaINTI1+WZ8cmqWBxDv/6
t9rhkaqanaO2IZhbZfxutXnqelzLR4nWhICMKdP1ArnXgwntsG/DFrf3aDFYc1VJ
M4ySDJC/qYAUO3cBmbDs1E7SbHV+TpHGL0PmbAExaCOJH2JeLNHsh3D7YoGH1Kct
WQ42TW1E6/6vKkdyy1nBJq8giPbzhP9JaCAhGBraQcAaoOeucCuPVVtDKRpOxpkY
HIJfU0V2qAXKCTn2VE/jgR9XqQY+hZaZUgbDKDFn6F+L1q1bkFT0iyaJegZykiA0
ApI3Bo3YFu5bytnyqK/e+STjEoaNEWwusr5UT2Y9FGFwDXFPDlV/MPRN7idBKZCW
qLo3zWkBYTZYUv/1JiK2C2VGSCN0T5oHwWYM2pOg8+16XAhh1MSOBK8m6p8gRb45
qXmU8ZT9ALu7MiNckaFDvd4XKNGEPv5VTgx+Lp0Panjly1pkFTCnRZYaQrN/LyZ/
Ig7x0A3yihldbk7uEWPf0bUgQRjWJEfouGzerTDXTLG5ZAAQOqWIb8XH0TU5xNu0
XykxJnvRUoC7Xan42G4wcW3msls90to0+Y8L1+HOi7nJZa9dpCBzaNA/Dn54CHrV
4QZJNezqFMWzRgEEjsJpai7L/dFRg10Q0gVeDiW2U4GZRhP8Gn9yNaJe+gYuVCK2
4qykNB0HJnajT3/3qgejOiZCC+1usl/+WuM8l7AEG1XLR8KqBMk0/mhjibZ3RN+K
Z0K6PZLBeHzi3RgK9Va9eOcho572BlSGgZyQhfCV2MwZ/IpYJydFwLPIQ73zwjt6
bLUMpo5PvNbMyiChGA0tRaAa6BxU3pCHHdoAae4WW3NlnWxmln0tYfTmzLgNYdxY
rJDAYwFVVW9KllGyEWT1WT6Gws4PYGHt83gm8sIsaFts6/ektXDBYs9FbACK1ICs
QqPPByn1lblqWuqYQHg9lAGdDootIHKCJlcJ/kOqfyVOYGzd3MhbMXkfxlnavjXy
8UTmrENfWH2Tr2ZfHkVSpHNUWzwqqbqvLoQKu5m32++pEXUuaBzBo8cONHYHrpSY
GY2knQ/GbYOyYqEn1VJY0M+eycXZfWabhjd3epOrUscTfDqjRxkGlOW/jDJOMinb
ik9aJAnCzP3s0vW0wIFftDLh+hKui1bEP4zkBNQT0oU8TD4nn4bDrMa0YXsIwKDJ
lUEI9go76Azzl5rPxfA5U2vbEw6oioIpS/VQqTAtoG09WO/luJ8vZRO2Xedgzqbn
Vbc/9Ee9E7kVOFN0rC4ES3bHKgNsSVRHhbKjj0cv27DFRRcl8izIgk49Q2utdxK6
qwz9CX6M4E+hUJUKYqcz+D71xM15iJkiljnBGCYnDCu7llryWY2BoX6mCCcX1mSX
A2PIugr4/w7KnVpEYeeuKuyhSwQwUoSwr7YZ2vvx7OWjShhX1F/XIdmvh1U68pDW
7KEDZS77evKKYR7gMDTF3cSazveGsu45Btj+NtgdnkpgcOB+xdle7LkA7FDnZipx
j+NFSJonqCY2+G7BjXGCGI3JLQES1nnJryB5VpBb/ogWZnoxhpnygwIxQ2uuXEyD
ZBinhKN0vnfO0YlvK7nILyI1ixfsQrstd/ZWdjaCDPhVoogXeBPAoNb3Q1UpuIqM
GSngU3j+RxdxHRmYXMn0Hf7/ZeOJ7tnJdz4tDGKREfIRXmV3dDgmLOdqV+YXHtkm
MuOhTBYpjwsZSiY/M6aLZQs2sb1VKk3JoAHViNKLCG8VfLfOIpyIcqkb2bqpG6D1
mcfkAyzgmU9PuC47m/j7yOX8LVap+idUqPTmFWQw+quB9NBHHceB72ND3MGCuavR
MGOTwbsS86RjHAXFpungGChlxjgro2l7Bx637+hAsyA4WW3yepr0uR2SRkVIZOvw
wmOIbPnb71neFxldF4oZLuIl+2XS3TSWvH/iUHBLZWzoVWjvT0nI2wj7T/5incvJ
FdkEc+6iCjWERGRAutCtZUc/hbQPFiC5uZ+Nk3V2y6ORJgPtGWJ7J3IT9iVWAuFw
vPqIcyox5xjpg7I3yDRTNXo8vIslkyBWURdRhpBUOYy+Ej2HHA2ygEhjBTfHjt0b
+oD0GJ9ryFc4dkMObenO/5LRtWM5TqOMMzNr3dWUJm9XIsYBgr9wS+yDkKBtD86t
tvX/Ms3k4TSeqft+lbfOcK2cRuMamx0TYga+tx5bUsGAqUwks0fQVFuBvviEv3kh
L1ThuX6+kCrjzS34khrRULBUT6AIXc/BMX1Qgru9OBOwBc7HeaTEEvh/j1Wdep9O
JMK0cj4aeWkfuxMOiWE2w5PrMkiPsShy9Db5MQg0TLzjhk8wFRsVhRUsESp/3ojH
HDMTR64vNB7h2oVFUOnOyLzes9DUwgFCuGCb8tvrNJE/Wc13O773/1nL4GUmmXuL
N+MWnp1m8VruFU0T1Hdd8RdE3VuQjvtR+yJI9XHu7B2oVS+MqgcbLVV9FStLAQ+s
sKC+FXfgbrYytQ8Tn6RoWCRn8fB7ZLrXyh0DDqSqCc2mw218sx7vGauwMmqI1p6F
Gz5HeVjnFMXopWKn1dRuipPJiDvUGJgewsVuBYDLlGHa667ah47xpTDi4bIyxRfe
Y6qsF5gv6yVOpiUBrv0T3f/KGALWywNA9BMmiTOVwh92HWadcbmYrWScFDFDjJfG
5X0/z3s5KZwgVhbqloTa5yRL1hGXBhbjeGbjVR1YrrG8d7HygZY8rp+mpjr76A68
bNL9HyC28AN1cD+wHWIt2ybxC+d3yva3ZYtixdM18CzzJ6ySMjOR9VfgVUE6umdF
/CDj0jS+PuiiQ3ETgwsm+yUHIe759CoHGpEluK7IkKIr1OgePWwVlETi3Zcnwjbe
d8AzsfLWSh9mcNqlKf5ycxgK91DC4Gj1fFmzKsnLy+odlxT/w33zj3esvNvpCY65
/QHKCfpwd3UawLns78et77UGOwCNorVMLZ49XfD8kwPzzOCnjvZqLn8UPRKC20uv
VrQjSE783KoYW5kUBzFzjku1bXBQyf21yNXD8q6nmbjSDtZyNAM0s519EabVj+UU
Fby8M4e37+0IaKO0y1PVOen+ocAqBA86A2buPRFIK7AWEH45WYO1Q67MJrA+7S0R
T8DSfke/Fras3gLZckDQ7PwsuOMa3lHLk02gLLCwcSVrfAY7PHxBpDFiJc+C1Bjl
hYXeKbJfTKihzBZF1i0PiwTQtVjxRJILySnuEIj/aMekONWWWGNNpK5JEVg4gIjh
xoPw1xmVvS1e9LADYxJ+xMCZWmmVL5XBVqMJJrAv9uuAqyV/IK07KcvbIsb+LTNm
z8SS6dhO8A6EJLACS47oyIPY6GxKuQOS/02ULAy8lWK0VEc+Q7z9DtS80dsCQfr0
aeYe5aXxKVuvc0Rdwjx5i8vYu0lCDLXUJD00RBE3f0czmJf9r6OqYVwfHz4dAYxM
7WCsQMTcVkQ0faR0D8aC75BDuGNM8vk2qCr+5C3c+KEw9Wk9KYG8THy9q2+CkkQx
sT6Mm7lX6kxqFVgYI4daGaxx186ul2jcSIiTRtyXbjDLzRELJE5KrvoWKKKRtH3c
KMl0eL7knoIHw5sq4ilzjgZu5Cw8S1twY/yLmqZI5EGW+asD6ODJTiGtLKxDg6fo
SheiV2E7uvCeEyqDLXi9qDe8T7G3nGirGbd2U2Fom+RBZza5RJ0mSlMIYb1XFLxC
xh0MOdiSjqgGFRipUwdaFw1o9u5Ak+KHjmzXP6j8iMu586pIQC7BrRu2tfBonstN
gFxWRDZarP5Kn5/pTL0+6XFgpc5jyqSpJB5C8GqMQcA+Ud/QrrXyhkrkUdw8Rsxm
VD91rViFWBZsDKk4da99Ur8nEKWdRorvbUfIv+PvKdPc5Ig5Gi7pmriBMIR76NcM
z0Jmjur5LHIXzki60UVucIYYLK5LaScZiQAtcIJqryf6ewxCpYOc7fznvg+eOlZh
zsw9kU/wELTv5X2RnWybEViQWCEC5canlTF0IbE54FH9rxaLtOlMM9rlYMi7hy41
Z2Q4bbFpmFO3D5+CuNzAVgsUT73OYm7CQ5rPW2NON2iJlvboS2k5RRD1PzHwEja4
LqT0JwKH3AukR5uyaD6r5Ou31pQJzeVKf3rFb6gMEYYkU4feBbvLfcGbewvWNqX+
ZRDO77/VlrXv/Cr3JIIbg/8uz+94W2IK4WgsSOycD03LCw9GoUs3hDkZ3YHyEv8W
kaQGRXvfDwMe8iV2t0D/nkx9iaSr69N+LRJ/FLmv/LAfuPVqyl5SSnAbh/1j0n7T
vBR+Jc8Wn5hoJn3gp3Jv1Jg+eRoh+HzPXjE9L6rLdEkDDELPOeFxGgPyjNv39BwZ
TwQ1bgaGgxnVrH0XbHnGcGYtTi0QJqwehTXi0ln2o7K5OQgY2730HozzdTH4zb+L
fXWpwBo161OcE/waGkBe52fqp2aYOL2tdGGHrW2/KcGb4QV70+JkSSSv9TqGpJdl
+Lwgwtgeha7xL47oCXkIiMvpTP5q7TbPEOJqdSqFS40GQJjeasWzvlmg04FSbTic
1ZZPV2F5jV1cbjjNU87qMrfWJzAeIxBATpjWEbQZJNGgB/l4yZempHDc8s0jAdxg
CE9a2ZxmjrDXeKasoOzOloDjHB/1S0OkpETLUbzVRCSUuhbL0boPRDhHxKKBYtLK
1rEqTR8dcMt24GAW+4exeW69IuTjXQYuUvMxGW8jKgsbio7yu2Y5q0zrxdTI+mzF
9G7boLugT5QSrJfPFWtivyiENL+x7Fy7SvnUWt6SAj4PtlbBA6ZrdaQm0C4Wlmca
+DCPQ3Rtu1lACGhCiGtQA1KrRM9mS1Ixb8XOYUjj51UOMqbItU7l7w2QuPdDfHhL
8DW+FpADk/YoxQPMYon5aN0FlTP0FCIwWoQCOjqBeqpaI0mQJUTs9gs5Aas4W4Fh
nlztjaCq/ZaQWQlOAr+YfZ8o6q7JgUV68vQQc3S/0UZZA8xFPnWm6j+KmXi6IlGy
qKUL9lIGJYhfLykONg5UFJ1L7ltwuXogyTS0m8HbZZC+GpGXGPuCOWs61gyPgWbK
0DhOR0ikdEzNIrQfrIIlvnkNHhFsLG6Vt/LNK8TPUAIUIsaHxCPduwTwDlJnQ6sU
/MA9CSKJ7lvSZAD2UV+XxcQEc3CtBGpQIn/txHLUUKugYbbbkuuVcWsaxlFH7yA2
PuW8cK31O+adJ/s6/0tDJaAp1DzirXo7l56WiuN5T0iY67JuLpV3IdF+HGqqoneU
JSaN1e7Cru+OOGMhx17EkyCOYD0kN8GNVFuKP6y3uYIpwLNbVs+0sBA2L+5YANSL
765YzCq0XTyDk4j+R679YZCBmJ/yZFW7RAFgu51g2Zyikm1QzJuWJNXQbADrgoMg
Kz7a2wdKiggsW4HkMahW10nigYBwKgrLZOqd+DxVlIGAWJsGjKAio7pOEanSkbjQ
QALnUM/dvxN9p1u4jS2+aTQ/m9NJaTmNh8tEHc1eSnkGnp2Db/CaNWBuB8sMzAtN
N7c5w2iOThr+CxWKbCh6ihw5oTjJii8VJMMBboSJYCtvvZ5D/Ngyv9j6W8hdztMl
vh5LoQMccmLw6E8HY2nCx89nLnVFEGS2cfsJHpOeGfQ37nIZV2PnAcrHhPtSqpIr
yr+lyf9t7hF/tU8SqvY1rFBxnbsPoZrXYYpzqEuuwGDOmAel815pFa5s+k9JARGo
bt8xAZ/uM0YbIHQLpxNxSR/YBjbNxuDkG9EJpVvwYC7EBuTx7UW29DZOShHCdpwa
tm4J/hVxx0blg0+YX8+3JINU6AOAWS6UaKkAwk2oFIDVBziOND0yoaLIC5LaWJq+
BCof5E5U22Bz3G1Jd5ahrEPolYLQC2/mVUwnO58zkiJIYXDI4iDXN5QJIYA9RMff
GbAqiE1waykoOU6/vNgjq92Q3Nlm1aeIP3t6VHKXCrLfciP+OhfwDujEpd8g90YX
Fma26Zq1aVRPUTZy6mquw9SKitTQgDzOkwKzYvj7KlwPYagSl2YKojTw685HL91+
oRkkfuQd5D9mnart9Njs38F6YD+nnNrKErO4vTH72vQAVln4dlbVbFzj9h+albVF
uQJaNjc492XFQaGCPADzw2epi3kIfBh8xuakFp6Wk/LdT/W4RVYh+cMp/yh4tWar
Cb2jY/2UVyg3fApjnPZyLYVisfx0VQ9R+zudIbW3ZW5yihqktwy5G7xp+uxpkdjq
ADN4I6a6ztfyOMtUPwoLxKmrS59l0pmi2jkL4fwXXPKvIRGixrso9S9ajE2vV8xM
eFqNukZhbMWx08hWNwT/j0fMzqvt5DQmxuvPhXyGIzZXnUps/1NV/+F6tisTvRxw
3CeSy6oj02LZ+jtBi2/+0oeUPkXr6Llo5UCvRN0yNvNwMexxjPEl8x8eTg2SksNs
tuzPFg0kcCVN9VbM/MqlzuHmbfGtrdv7iG47/PGc+WUb7tlNjt8SX6TnTKFiA6sw
ByTzqOJcLIxIacy/ZYFbsKKCq8EtAYSgLZIJEwZcvIa4pN19Px11G7NZyA7EdakL
9eyEdSstFOD/6CwrhCrkwj586T8jmfHpdiu8LuvvfakO2T/P4ZYTzCWE24gM4gUX
fVg58gpgNtnPuEp84G8v9uMhPU5SBagxVNGePULREvseJobHQ/52v7H7NopHz/9n
/SLPd/5Cbq4w+0yIUn3B7nahvod8p+nO+EpCks7LGm+KZv12SAnyGqwwt+dkQzkR
ASOWM1vTv23Zot7JaYOhBF6f9b7FBoDqFpFrXcgE5DRprlPZkqUC5VLFrRqJL2Uc
5h7hmMcVukZuis2onRxqhbOn1djRWwmOkhX5rGnvMU7DUoVdSTOG/jEj3enyuy0q
O4YWo6CGE12upu56irum6GD9jX6KlsMY9IPNyWkuH5koJLD8D4PRolHT5kKQYoee
8+nlbiF3fRPCwwtxF86VIB8wdoUSpVPhdLue09Cxz/+GehkR5LOMsg5nT1dNfpEu
sbQtqs44a0oZETKHH0eMrBRzqbnFCcJfTTuzWAclZIYbRJ2xpv4TAVxmxj0qWjXa
lobIhL2arEY+uoy546HdxQF48rOgpvO6Qb/QSg3O/l7Jl4k8uWV0TreCWUHH3iAV
lWJxh72lErKORa+akql50vIQpi0R8HQDTaaq55wx2qMDDRZFjsIT3D/VDDqK2sJW
CEAgTjdCMW5tOP3FAJVzJUvq7n0+zzmeefv8H8I0qOc3qB1cK/fa5oCFra/JVokP
T3KVhYCEi/uxFeuwazcco/bIvTZbz1XvJYqjmsVchpMbBdNJafv8HLQnINKf1LJ0
j9FxMheNtDsa3rKUuhBZKIKWJQHPVn/0inR8yORYC98EDYcAMLBNrupUoofGPWph
q0pK58T2pcQdw77SanIPvllWcmzUoHs9Eonx0U06OAZ4RIyAyyBmoR/c1Udc9M53
drn6vTpqP7lAAuz8UursHDIa58Bt7/H6+OlXGG6nL37AKn6zc7Wgcaf2b48fX3iJ
wqF3ki8yjA8WaEl9b6/HuIj4f0rGlQCxq35Jg/YlkahwCDJsrG9xgB4PWkZII+G0
NQLqrYyr95BiBQ31xHgSgBxEih8l3ayaSczsc4sVQUJzKP6EhOQ87pHCcr5q2jUV
AMsrL9RB6oBMqBT0yAyNDC79MR++2OgLGHMiteuVPMlm36ahtgDlbWL+Q4njQdOa
4ogUdz5qe9r8xDdrVfwCOovOahRXWnjJ+fNohGY8zqB0yzSPpHKooKu/K4/sgQ2i
KTk6qE1HZ2UCcNQgSKYE8Y4lWMQiUqvsllWl5b00ozVgit7G8f0PGE1E4/4fXV8b
Lzh5yF/sMgBSPsGdE577kFRV3WVrEanq+F3d1CYCcWm2jctkl5cDc0+Igvu6djFg
4Zq7toN0P90I5dYD2h1RJu75UapSVqf80h5C6403aYCHFqDSHXdFLj70znMtX20j
d2abMWiUVy4MArvdASsDaPEAP6C0DnbWrfTkwRPgcmXgXWe1NhH1oksyEv7re7Tm
CCle2oqt2DFxTEiDYSQJ6JH3UY0TTED91VRxyDwz0s51sdkzG5hUs4DHgeXoKuek
Ue8rjy/qoZWSsTp5ko9yumWa8bS/9sF5S0AUz1Qv8XkZz2HEKE21emSSOkMeIm9P
VYpSBW+xX4mK2uA1Tkyt86l9s5V08zDeX6BNlp8AHI6nDvPOzrmhOclk4eZNe2hV
FBrhzWhfXDEGsRNZg5I9Bfrs3tqopyKS6rFeC95KiF6lRzv7yrkcCx87p+ZC8QLs
oLIO7tqPT8hQiSP4QgayuwKcf+ORRNxlGtTj+ZutH+oPS22ifqQgp0q6Sg5NZcIc
EC92w4ars7VjDSiVxoPBjiU+qeZVQJso575V+jZoc1Bh2PLQxogSGUBaFuawZkTz
9VfhYdxtAvOehxqJfnh3l0JM2u2tQKhuX2GA24WW5lxa215zXLqpsNAQOdlMnqS8
xfdCF+4sX6Kx22IwRcmvsGb1iEr+GOl8mPZSfstkWPmm/2ajVhTEYoM12HgD98OK
TGy62JMhoqDmijjk2bNCdU8XaWZO3mS9XlPXSKgJ/UDG0ghClR00Rj6BZsLEB+t3
o9V05dT0buDHww1wGFNUfTvC4AXwkczwP90IoW5KjmsUOMc8Yu+vr3w2JDGDJgC9
cJbicgeYzFmfJ7uKf+Od+CcsLvc+8uItlN5Cr7AqeO2E2aH33u8X2Rf7QXqrG3QH
u3XXfpOt0ynmTlfrTUMyYxFnFxnG6pMPcn5RelX5or/GCFfV9gVdZcVbuaiXFiPS
KIGa6MzUJ/lck1SehnnLqSgh4djal9ml3qh20FHZQb46lTZmSr690I7j8eyXFV4U
bm2GSOydQMA5stGx/nllneWWkjkAge6kCjrs/E118fgoT33k610gZZS858LULRkJ
o7DXI9GX6WGmMNvjAwJ/L2fsGPfAk3l2/gaUJJMBObuTPuswSwIoCgLBzPLCJD6r
fieJUSobIQpZAw0dhcAFnifHyOVJ18GTwa9ZO3zBURew9+NtHYc/FS6DXrr8jHpL
7QR5M67Hgxr4lMYFjAwOA5Lu6oYESdqAfoTEFRNO/ehe22JHolomMS86NGBfA1a9
YoEJJ+5sfz0yCm9xXT5aWt7tOJIvdDeJSd5KVA6TTwVIsrS0hu6a+5PJcYjicJX0
/mJFBBNwcYqdQd3HFKMwqNXEjl3EnH2vm8lXjLapy26a3bdoPfZHser8M7l9n2PS
5QTQOwQdgmDTak4LoksLOi8n1QalHWiCPV9GcQJr1WohHooI1hhcZsSThWPt3xZ+
dX7vL7Ey4CxALa28sGgdpd/WiGm1eta+9DEZ9cEk+CIA/LHYEX4BzooByhxttl9F
Ch7EyxbV2me+cX0+m4xLxSls8Rrxi5dIMBtXYbBqiJMkIlv/7Fnr+QbSkrxT2aPu
FwfX/OlUvfA1DLzQ9owq7xvXfYldVxPA5rLcu8CGxiVdZbyqX/WDCNTkzf+aa1E7
5sXSumBrCBGbliY254l4hpDEtgBYdndQttL3O3zwdci2CGKxhONjtTOfD2UAtB6S
9u4w+zujzyKJKbeyNGs8TkdyVRQiwJL5HzalF4gWa4f23Yqu9Exuu0KJ4MvVGMEP
xEh7A4ZScaG/q26ys5f/P4iWauRrHp9LAecAOg2rl37U1rOVqvHzaPQNaN5KLpsP
Ej+b0FanrJp1vfWDsCtPqzfYyMh6A3E4INKR7wUJoqjZBlA379vjbGQrgtkFgfq/
gMy7KBYum3dqMSsJFTlNG3S9XCPPpw2TE2lxcEsTXfBsm4NiipvK8/aUSs+VQ6Xc
2Z7r7D+W04XypBido34ZSf0ML+iNyYNbSJ7UJqZPIzzd8mKQADxx050ZzPGKPgBc
Q/OvoC6n3NCKjwonDYlym1cYr3RmxY6/vEiaNvX2GffSr3tqHpfi+3gtU6rzsp3a
EwD0yTzjUcb/mKZ4TBoo8dJHeZnG59dv2kVlHjNxbX8kDBoSAIBUbStYJHiG+Dkw
FKYVT07n6RXWA/dqgKCCSGDdtcShq4kqsyqwOuUVFprRRcOGk4zqg6xuQyBjg3zc
DQ0cz0lft8B0VVgFpMU+5eriGYSE7cq886LnVfOuA911SfeWFIQHx7756emjzPeJ
wM1okwBZhpCeh2w+PAjZFXYqTadnjIpBjGv36sE+yoAsun+WojlSRIEhmou26ZCL
6e2cAjB0ZKWYMa3YoK15dy64XkRPD8fUqiJmpR+4b28q6hOeUBDsOM1wDBhj55D3
9FTUn7kUd5rZuUW4p8iFTXcgXiRKJ8i0dxS81Z+PObGID5auJtFvRqJfU8BYkced
V1ZnZVE+wDgH+7alE4NbYgHtpUc/pKkLjGi3Ry2ryqPi6ro5INNtMt7uTo6B7Kvm
qB71uKPcQubCXbUEwQuUm78FoVa+YcOGpnyqDawkAmk3/sLvDIaMziHazvlgD/eY
X+FGMyFaF+YuLW2naNLqsGBQLOU1za7f9XjKqj2nawgvFeFDOlW2NibitU7TERxq
ggWCbJ2rCDRnTMNeir3vzghzfZn1GRbgvR74qNhGgcoQ1hS1jTUPNXNtXWwhaM+c
yrzBpqgLSIkxA0+9eGKgbgkk7X9yVTjH8kQXSMVE0gBVMOr0RvhzOEDuYxCK8kG+
qhc/ve2k4M8aOg9axoO1fapTlkeCLricVL7sjXW8JYnNfr4xiQ7ilNuz5/TSOGhP
RHg5ieH9UZntA3Q54M3YziAQ2FZ6JMpaUx5nme06KFEFGgxb9vgkcPj9aPU36FgI
aQ8EK/bp1kUxYqBYnkK508z/IaWKE3tRkzG4vJoxzQkDfH1BmjRA0+h+VY5X+f0b
H/0EkNXHqZ11omYnLOfW+mR23g5j++uWIMlA+j9QKNSCqOopS9Rwal6PX/buS1di
CFezDHFscrE6KZX6b91edXvSL+KS0H646glMr35m0RgRttU2ugBtjjsCOp+/qUvP
bnF7+dixM8g00wEXNiYEuNzqNpZ2ye8aksqzY1P6k9kCkL7tI28MvtKO16lmUOzJ
SE4spuuitHUoNBIiUchktSYFtrFuoiOVWNh4CEOZRUkjYxaVru7PslwbeGnPIS8m
of/mlV88URQXyto7ysoNxTxKHCIiL62fPCwfmnHpXfg6Q0R9+PCAznnpWP4zA95s
YCNe2WKjLTSVqRBathbdy7GeCE06AVimOowrVvteMIWTk+lyvaCsxRbf8cMdrAzu
6BM5KMbRJa3kkI7xr981EaoKxtOyO1hEjNEufchXIXaZKLZK36KN6I8Tsk2PWnI4
R2q0AqPCp1c7NL0ZqCCa9wrltv2L6kVEsnZFdiCOb1+BnPA5Swd4HsQGD0PP/EFh
1+YT5SV2kZ4yCnYJwxphNwAVRKkYoD9arD1fKI7xgjOx1yol7pFiLrK9u7SoL5Op
58oEIJTuvlmoRqgLrVhwCFK4h9TzhYNKgLraVI9peFDtmqi4ckprQfypAtnctNWd
jrF5v3zae9HTbWg7IWT0K7f9xxmL+qeSu3x2+uDR153Q9DhTonc/IfH4vdb6ka0U
3VHhDQQufeF5e98FgXi3j/2tfE+I/ZNrCo6v0Ll19Wed8tguIZOsQ9BKLMTPRCcc
Kvmmt4owsmm9aIdI9OdryObykNUBMYITNb9/vSg3m7vzIfbr8K/NI8dzj5Sc7oRg
chV0zle25D/oy8EpqPP3ATSFz29uSCwE3UHg6S6jyrpnindn6br6JQHMrmwyWEqp
VBe/6ufr7WFiRTRvk3ESvBRnNTVoretWGr7/aXLXd+edsnOksLF4pIai4xkoDbuY
KNdnli3qg1pZ5vRhBt2bY9L4XVft6ac+t11UMPU4S5VCqx3jZt9A18/x/SRa07N0
yJ3zVGQwSSIG4k7mutLo8MlGw9CPVHh1fJ0qbXfEQkl178pbABh6q/Gpks2WWv5V
2wTEjDgWA+rh0Kwt2CS7tmprwyUVPa0JIePkBNy4cIA4Ys3P3dGUtiU94nWfw9Ek
ZT9dyfcx5Qz232d2S6eRbisGgu7lPZwBU2IFppVMMS7F+B66VvSQAlzasiJ15OBc
Yq/ftRX/Hzqi/m7hC84y3P8mAeyxS/J5QpIspQMGLnYF0dTJLnPs73xjhaSFeGFv
M0BfYAwHbtdjHqvsSqeEZRwpgOaYu3QRL6pTcMNpz6/ctQabRWut0LkXjaNBic6r
CmrLadca8mXMndbZoYXap6Y4QFKGhKBviy/IJvY4xiI4bv7g1wWxCoxJ4IGNxxnl
FoBFM2Hb8K3BV/uIcgnEXGSrmiIWE22pGJPrICSWWE4MnOfrHvDzJtifQMHDREU5
0jXHN37miTw5HQ+7sdonH7E3oExw+HLZIA2uHVueN4gizNQDGbDd38W/GXpddRpc
kudiT6qlQWN3v/fzkfaZOD44f1Z0zghfzOzFuRRESJwKREF48AdFk4TspsiAXuhu
AbVtLSrijVUfNHbSBSLDErxHB2b/m/iJl+j65ca2EoNzEWY63qpiVQtjKJBBxI4/
Nll6xvVACvkdcRsFqYYB0HAWy2RqqNwHG/ks4cgCGkbCnX5/BiWYY+Gv7ty9vuwF
8zyWHxh/p9qSgnC9vSDuWbJharnkDo4VlS5NohWHqBWvGDopz7vMGUrm2Hc0kmgU
siM2kD1AI5APAZP+e8CaF74+e4y23mQMWKEfI1/Vth9lSzNS2lINCT0QUmDQIHT9
ETcg5gz0ttQXuhc8FE/kHWIYb/qVMP/8E1Y6QNsyTPkqxBjZdyzhZ2621CCWKhMP
G+LIwvqbgaWJJiWYHAkAmmTkbAUvD0EDEn7Ab4Arsdcl7DrDoJR9skwWKs24DlGe
pBPQIOhhy/GL5JxPrtjMU7yOc9hQi6udoyecbZg3HCCMxbG2Wv86jMJDTat8wZ8i
0hfAeMLpLWdKhwxlc9nZXeLus/MR4osJ12cP8aollRu1QcJ8lVW/OKEtpPVdtQiO
gAUnKdukAlf9EcsGSTAjtj20TgHXhkUBCVRJUCgGSUE3v7wqNzP+QGMbtT1fE6/F
dacn7d+Q2iTAYj5FXzz1WoCmS84O7jC/yjs/j4E+jNgoZSDZ70D4qi3FDY4EhSQO
n2kgnJCl6SwzrAuQecodbhfeRqVsViffCHXsitrOL7lMXdiwZz3AqdV9Ma8AVUOf
yLRoBJ5h40TfazcA/0lUzDyf0/Qg+b4E1B1UXufeC2YCctM4OQ/qyqh5YiAaa5cW
yNYnpfJQa+73X18DuYprpGVwuq+439FzO9flQecH1qUVW5zOdSpUVOzpQ825wZq8
k9YXnOutgJpfztYQ+0ByvzsyNtaHS1+XrFa0dC3JxwPH4WPAEKqZDSrdF8zcay97
nvkcNlJLzP3hHY/vCKIJ6qd+tyesY3YNmJ/PyquKD0SBoou6S13BDy7KKSYwUB7o
KCZeg+jNOslUjpMhX26eEdXhR7IJZgkvPAnQlkxaU500iqJxz2ioILLwNJtCVyuW
G3timbBDzN0QIKBp6MlwFe8EjhPNRslQb1MTRsiXekg37xivIKIFISYTGxPEr4Bf
eetOudfRAkJWpeQGRI1ZCHdc8aTSdONxb0diWSQNwBRmGYtwFXbmXGlAqeXbq5F4
TCgrP6FpacO/SG98evyNr0iVh2hJb9oG5vUS+dKlF3n9Mr1qj2696wGWCj9UaapV
T23DrDIxRQodwInZw9LAxQzwQskv9SpTl4jwB5CIEWPX/YHiNkXOyr9mlIJS+qy5
GCLvyfOabcCcvckhIFM038p6b/VvPNFK/t3ghaNPbQsxnADRIIOk6U0XSsx7JNm8
R8XKQL4m5JKhdxs5Rd7bMS7ZUKuEvZ3uDjK4Mrv3Rnx4PboZc7tGFiNukRW3JrNW
QwHXZzz/Dj18S/0K9WeEs6L5gB7rZ3P1tfM/lxadXKAuzT/klqdQVEyJ9+fAyFBA
s9jsxWxCxuVmy1J+FBcO8BtQ+SpkOKyVivDrMcQ499ikfnpOnJRbGWGD2uuGBYlU
cgRhE4kI6q+ElXLr7zwkIRDCbrlTLRZCIobTaTWKNbKtQcb+1fTbu1mwfx+CNJhL
9OYN5J6M/SdD7gwJ+7GrJCaVUVMVekBIzFCR+vrjStKOtxoQkRmTxNrrgo2T0/pq
SNze0aeHlxv+C3d8lljjUaLlGdILmD3DyJFK9PJ6JEaK+K6IOQ2M6zO2y4lYJQkY
dobwZaWb66cCL/HNMon0kRKb+pS7gHmAiK51lFOku4UOJXMJibOgEUdCv0K6oAb+
jmbV/K2syRC578U68yQ1zULM+EjtZTJEmKmN1s87F14klgpRfc/kNsxm3svzL/zo
XP6Hx2R+99R8MAT0z1zrkROiyk1vCzNp+xJ/BEtd1afUJK1kbt3inIx+soscBBWm
3qYxqXx9n7jbXCm/EPaGONMbA+XMYDTQTlIbcBZIb53eH3zOCaRsJj79cs9effvs
6VaBifvgL7w7cOADmAMQy7AsHp3c8bIVd7fblZPajaWkq89QA6VFBNej2oaP2J5D
ofC457jZozvXLyVxgkZSZmSFnKLlj8GShmVNmDYAoWQXinBuDuAzandIEwwCPnU9
BZw77hsI8Jyct9jBWPy1I7zYwdNgKokTzRhM/nQjwwxQ9Y8SNlhh7/HTHKgUme8R
H2cJpJJaRpjf7McSNvmr49LhGyNBrFEpdiRiKmxX2V4EkJeTfmus6KdUzsZXXTrJ
oqiQbv3FFrXFwkxkk0y1AEx/3TKQbtZJxUyf9SJL47AVqpKh5QBKci0ZM2uriotB
TrdLCj/KmCwSIrM4euzlljzpJEzFPKxPv53JWEX6a89BYioM6BIYmH3lslzgeqBN
kyH3fUZ5zPbIYZp4fawk8JEFWeqNFOC//858ja/RM/ztxnd9SEWB71qF9LAD9cos
EcuwzvXkhG4u00/ozJaMAJXqBF38an1WkKkW6hn6TlLqAEM/MtCg9ggO1ZOsHQKT
o2IvWnUhF91aFFyT5InYB6wYWN6aJhihkwvxIb3tnWDi4cuF3cIcwhL+4RN+l8Uq
11iWpl+f2MSkwhHJuo/EFhiPgoFIi/HrWztiJSdyR4OIB0ch2eJtZu+ld4mDykPE
5ZlLlZjL8a8DbPlrgBRFdwQ8KBekrcgEsFQzKYznHMLNoiVtU1b0+go0CtE5tA7Z
8hBG4L90VcjA6veIcGPrEORWRNScYWzvwhYDf5JGXYzp+VrU73FMqrprBjTlV2yA
jvyLcA4Av6Vf+zmXIB9b/JP1fTF+XhmIYG5ef1b2LTKzDn8jbizRmj/cLvXSrnM7
iUVf/B4eVYuFjRXi7g9OGSsXnlEC2MMf58GEcih/QbNi3RLKxP0C1tNLOW7RHuNY
+c3tNnwSyPzKaPQu6rHW60a2CTl50sdY3e2KMoMZvL0x4wp54gY9dPxGaoL0jG5/
5+6xNMr/A7Kdx2/7MVaoDTIPHQ9YTD3po7pN3tAA2SyC/vFJvohwGBaJtnV1f9mi
OqzNYA9g9GN2ula5QoiAZqP/BbxomzWYKe7k2YGDqXrydysAJYvwbG9cnP337v/S
0xCyiCO65X+VrdQeLPhnmQ3+iRZfHecuIj9V/UcL89LFbRBvh5AJt9qulNxLCl44
N9jxQegGZ9c3nZgMu3RFkizoEqVZDMQAOvnYPneMjRqaA7QuOcKsV41+KT5BrNBX
hHMPUS4aPWgbDSk6gQWa/7ZqYVN2X9aEEnbvnfqb9+0zitsy6hbGD7oiomQVe1a5
ip2Y8piRrQGcyD819Pm7AsGpO0AXBdo62p+QWJS1Wmk4vNHCLM3TFb8LfsWR2yoc
52XHrVvGSZTf3DZi4LI2NuOHo0T1A4dNo/rsDmlziRH/gaUukPk3dFjh272ubdd6
iKT9wiCnvYLH+WBmNj8wXvaf6DcLeMZbgwLYkFdLIElvkeQlc43oMNXV3/ogt9/b
3K5tByXf991wKIRtw/RuBa9JH0gU8rL0TdFiGoVnhVdQk3e4NlstISRq7A9XOXkv
0VDryH5SmF9uGIu6zI8lWIC0uaigWKTIARfmaMrZH9lwIVzshzz3oTlADnosNtKk
4nH6ld3XLE5qwO1loOMmTqZhUmRTt5/eO1FvKjt3Mi0/Ie0+IeqnU3/CwsoI+p68
2yorDNbXK/feCiGZQppcRnpn/WbWXDnkK56htNYwENUtddo0coF2ZsGyToUmnLAe
Z1RL7nu1cLMzGnAfghSL0Oxqty4HbaHeqSurERFbBuHBgWEXJJETuHUFdddxnXa2
ZXL6ca10YUcvfkc9Rx4mZniuYekYp9EKQE0MKex7Xhz3azEAzFFdZ4celItqlsZP
RkOURFOpwj0J6aaQFoDI3+UetqPYW6hZMFVmsdSlMXuniHYyODfYohjiT3SgTZfR
g5vOkBdNv20NBtbhZZZdhLtB1pan6Q41gfezuFlbchbnOIgsDxeJmfphgpjShAzP
TOpNQZtjkzUBlAuf5e7tDUaM+lm+agA6THFM+soI/s1c3ppKnmu5qqz+kfXG9paW
DCV9N/JR7FZ/mCNVqlwifori5j4Sjg3237rBWNk0IExufQQusbOIm8NONXzGlWoq
HNVc086CkHiBjo0YgwzaKzntPFcFOKC0Um0PRhB4VHGky+Z+OMfRDLgJf+qSOSWA
YCOui3dk39v6SVlLqnInDza0u0rsfBmiSalyd0IQvl6LmqktSdjwURNGjdHOViYT
TUC2nSwTVapB+RC3H/eenvX1fO36DoBEwDDRAnUJG3zRpftcJNfPuDSep+XFwBDL
7FvdvCF7GlyDLwEFbHSh4adGjolaJZdyWr4RZe92PWa3CIIb06tuYDuC7v8kMVSy
S/hFSItV4+cXIq2UChhzbQRCUSdNZdK0QWKd0kAKZ46FirriMv52DdG17PkV+89T
EVehx5XpeeAQnz1TZ84r32rIHAdaKZuOqG8AICyDo6Npjm7CoPw71HlAYTy5k1iv
aI3ya9eobx2KCKAv3PHA9Rlo3sUJIx4Dlm4uwczW/BraN0K/Aepl59saPnGBxeBZ
4/om74QQby/3wyH64MpuOmW2pV17r/mO4zu9XSHFIQRyWeCHvbb86Z84OKPLVlSg
BLtI+noY28b9jYSrtA0iouZdB7ZQYz6J3m21zde3piP0YRXw9wuVnNY1GP2KSYud
ccQqhqi+whL2iTnP72BswMzVPDawY9k+rBFyt6KUYAE/oEQsOFIFX6QF02HeOYLg
7Gi0y1BBsCoYqH4C54qYygzWq5EWY8MQe/dGkWZZ9TmSaPEiAjbcG0ekhCWCgZaw
ExnU7//gfTif8wBHBtsW4eDc2bTl8UnIB1k0LPxK/zqe3+dqf0uiXPVzf8HaP3G0
cfRTCATRBWwu/vgWBDHyC+LPwEMo+jX5mmpn2zhK1UB6Kvx15SGiZW3/3v0NAcPK
i7haCna+M47YyTX8YICrw6+TeI5+7nVXn2hwX+C3IZF9yJKAXh9DX+p9NXCBZllK
yo4Fsp/DWdeplLZFhJa5Zj9E5csQ3gU80fa+ErZ0ShfpZHaPYb4KMVNcE2RKUWyd
T0YLVOl9GbfMkrvpuQitlq1JqPlrgt2yimsDW9Z2+CvzhJ/MKcxql0XRTRYdMNjz
A+QtfM6nFnwN8wUcZX6xPhi4PfloavekJ7N3DKMaUujc3ENeeEyj87nzcbpE9fW7
tEvHtlbmTRmIMGtJsrL8hWynwtEchPCQDMeH4DLd7lKLYt36rlvQIWGQ0IahPaJk
KZwnu4cwI7ra1SsinVj50jR95JaShniSikdA6jqWcnuTk6jqTiL9nWsqPxhCupTe
HsTAmG8oR7O5tcgGYF2Dr23+PoVkxc96VKOhgeoRWPqX1eA/fuWexB9ACEEuoRY0
0YrTC5DcYQNPmCAS9X9+8V/gTi3BQ8iRwwAF3fEM5vsqN2EUlGb1cWD4X42eg6fo
rUkdAqOBTaougiCu0Qkdfz6vIQpXNPoENAw380H1bG7wBLEU6SzMPjh/kNrj1PCb
vEt6OEgo2FE7LeSbS2NBH9CU5TWUF9nbDtoblJnF9dh1+iu2QMiN34G7G18J+0ic
h2WcdPDBO1FJ9Fmrh8DyZOrnsBlxe9fowY9lTwZ4M4SRPc0e69ULioeB0tp6oxh0
eCJcbZFMD+8wavc95YCc5qedJrUUuWJ+9IPM3QEukU+Q/uHp/13QWGwCuGcyq9Js
jct0zNfZIWjHOIYCsQMj2txOF6IfQ1gIqbwg9rCNUg4DF9vhW0mHe8u9mmBxvL6A
dKxNa1Im+UR0VmADQWa6wscOPC7SiSO7Xckx+XE06Dkm9VDoq4tv0NvDM53TIRJb
aTTufQhWiINkJtY8yrISk3v3V51W3xbscYRy5yzuv2/DLamyCwBMMR4YD7aOtjnE
EEXfgY9y1WPJ+KlFoiruAELWwqIRP7YdOpPsZVPCvLaFNj2mmrpJ/YKsK/aQioPr
dSjB+Vzc1pm6LRhcjtQt0vqLnInVMt/CnKSMIGmi5UNY79SOkcYJFM16hLCEwCop
LBY9OG0vFxtxBD8QyGfOHfGEAh1xWZDLIeuh+pvWVJplhfa4TThhGu09CjPzg6lH
nikMPH8jwWtgL5RfyjDR/7N/bLpbC5giTyb6Mv0wjpTtk5tzonaHHzN8JkqgzLGS
V/3IJyumPH5iydgdqe88C4SVZvRpLnDttz1WobDMOOTZb282oPUF34JgBXfQzwgj
Y/OeZmpMTVIrrW+Sf8LQCSTwU5HviTBV03doQcdKBY/qdqsLOxrWg6ASZHEtIkPO
kjWxywcP3xs4uqpIfHE72QefKcy6pHBu1/FIjBWQmXbnAr/xJ67T5Tyb4nlUfJpn
yGZ+kog1RExTWq91Qv3IqHSpFO6pYXwQbMpYhfYZ5NTRlYbNA4cvAJBa4xkUEhFM
MS9gdlZzx0iJN8xDQIu/HJ3U9aVACU21LSqCIFqXGOY03yqI6UAEQ0wiCp8mfsxy
kFTyLT8MOxda88QUy+d8X+JRHn32M5yKBGas5Gup/8fmdnBz6HTHAYmPAx3Huaiz
L1/jHHCQWWSDnmazqoIGjJB47qmIn9Cu7NDArdwXIZ0bf3V3pSWhlBdhu/Vc2x4M
n7xZfczZ97TXh/9N+tIA1d1MU7yUCyH2SSsQQJ3U14vXQ/QnK4v/TWIZ904xHZo6
sV+BZaKlO1npXLReNVjqEmo60r2fkN735X+2ujrD9ZHIObQM5uDdpFN05tHHAWRY
g8CCD0ENq7E4iKb4z06hUpBJOZyr8G8iW/QWaZ0RMk2cS0wKf10OLL6sSASTBH5b
y7hsZMAxV8lSOvYMdZC17cpYwHkaRaWLPCP26LVq0Wacy9BTu0w05JcRYZIosA/e
MWhtWTvtsiWsPzVt8cfvR1Q/2xafpe+Y8CvvQ08R6wyyf8h8tcG0FYw9Y7V/v/zG
VLpGRWCkcbIXR4bk+SyFgRhlLSIWsdGGFUw8uHkZwAtCzNn+2P8+aHoeAwQZzvj2
7C8VUAnSsVLz+DJtd1Ye6qdM/7ARQOUQ+L9AlLTToCvKln+jAdxXNjKLC8xho8Ei
pfNa5spe0Oe72DILCC619hyU6uDciEKovNtuFPD9cUusXj59A0roM+3/lz1rOSOf
NGmZrxLOPJ5HQWEZjyi5HYp0bR2TsFdjJmvXQ4pMXeVkKPkCmYfWPlf1qdoVJOVD
240cJ2177+ILrRnGiBwCf3wR8W3o/U9w2dZTZ3zsLs9DYni8nKBHhHOFPXNRj/dN
qmykh8RUb3GMFPBRdAKISEVHa8B5ZoJzOnxdQRmR835ufE9uPYphJr1VPnzzHWDI
aYm61z9x7xVetNYL3Uj8paEuBtyVakH7k8PWyAUwjs9rU+s1Q4p0+ysM6MoYJDdj
IxV05KLroloNfxDa41qlzQIWjjSWlhJeBzfXMGgCHzKSRUGr8U++D2dyYPJpymxV
64ma2frGMuChdsv8sGDnlkeUUcb3BsTJA9UZpLZD4ENnNxY7ES7udtmX5+GeB6+3
Xlc/V8EqUyuL9GTyei692enHBnA1uVYvtXJ8TtoYQYzsIvv5PWLohUxIUry563mw
nx8Q/V7qk67T6SJcxTgRRZv4ZxvcL7wNs8jVQX2N35+WrdvqdMR/gm6gICR31MZL
VtyqdMPd6UrHkcUd5qjG1ZpDeLKGgfME32mwPHRsGa5E1qfmLKIr9M36ZXTpyInf
EkLBpAVTCRo5QapOzjldQEzQAC01UE0jEgQSRXo6EPKdCphKFff2d0DNmrmBLZqV
ew8E9fuRASLwC1yh0fW/MrpTBkPTvsMYHf2EazW8PdOPmxxRtjX4ipATUIpcqkxl
WRcofk3ZUuq9GB+ltVmBqC5F8uON/cbZmTe0iyk80RRBa5yPZYPiijX/9sBKxHLk
dBMI1uorGVzqNK8B4fIEWaPv+QT03Ctg73qxSy2ztSSUs3Y5lCGu9HxiTUwo3WDr
pJjnOB2gGoFjFhO7KM9Zu/EPreD5K4fWw0jyBKBdXfJ5uDqqXFwr5uoRy14NeiIt
kE89tnb3ET/7qhSaOa32DOBpji+Trcyz4oo8rTbarc1k+s4/zi38QgMq+u/2tpSW
lBoemiaLEUwYswww9Xp94dVD6PGs9Iy3gSl06oohOrmkFqRQHcILqKPVMHjupVI/
YVx3KFEGk0t7kt2QDMupnIUR1XC9CHLKS7RF2DX3SEO7/tenBAutTyhB5gHT76hX
AsanDG5+1E3afoMuehewW30gPkTca3/LwCtgx8MpEDYvfFKnGSrXF+wnsWkK4ekR
gR/URTs9JDBPqvSWhg/bEn9jSfzGzGDvVb/2C0tGkHwAHIPTXoswZCPJMOdq4Psb
xgpbUSr0kX0aKIYj9gKQ3U/vS8gl2riKdMHqWf1gYC8inBLS241FsBG+Nyy/3OuZ
NCOwBZFFWr9EspYST64mXu7TstId3tSBm1Cu0Otw3eRkMPB2CK7y9tYUqVrsrzOx
gXUAXxZHODFRR62FFcn4+CEvaCpKXFcQ3R2+sEUjFoyvG9+Xd9JK0gRI7mQvhzwt
jxLi+5q2KdKQMyIngx05hXa3xdt3FsXcDcxD64ynX3iIjLE3TlHTKyA9T0G9POe6
zu5rmJGaMf6+5Xj4DiRebpkN8unUwuETcugrsZFePWm1Mn61aAHRTDIfiH8Opt7U
i3yScTSjP3v3JTxrQ6kvyaSxbYoc5wF4EyP1nR9CGUGKn190gaR/wqJs06ic9SYW
CtQT7JD/GIb549H3+PCtETmhBBMS0Fv6v58c7VK/A4KU489GJH372Nmjb14TM3CP
3sIbDb7MMlqboSLFt16chEEUkJWLOtZT+4aKejAhIpI9q0NCIgKnqyfmztZjkrve
7V5LY7fUpQPyZ8AheMDXVTaB59RbZu3id5kGbak3d7MK0tPIpGs86x21uMB3qETG
/XxN7UvGosexeoH5XB5q/id5gPiEcZ1duWi9xW2wxRyB0aLorgOkQsdBlXussB9T
r8Eyvx+OBcjZgHLDsVt952CABBVSBHdRgFn+PZXTxajWvEZnOffTQ/xEX0O7yXSG
9/uA5MvQiTCXF6GjBebgqnT89jt4I9tk/yZ7JMhNPOaGSeqlHHPuPOaq2nFs6M0E
GQHv5x90eKde9dQwaz7WAIpEYYzhPw639UmLY4AO9Etj/DoJV9V86H61o9IE0OTG
Npz8pQ3sAMuDLayTxgWzUd6IGB1IbpG/dwqNe/Mi3qSoY9HXnKQGu1sk5BoXLIf7
lih+v+vbH5tRJhH6Pf6nVEW3gXwW2GCoy0232cbIhunD8thUxQ0ZG0WsP0kKa5oy
8RbymTccggfi9b3O6j2L/TfnO8zBoY/uXWc+9QSU8b6dPaJ5WPphQmvbnhPEWH58
FXb3RXpOtO1mONuR4tKr2li7s8pWEq/s7Ps+7u99ahp8RQKklTgCdKTf3viSn20R
+Wpyysg2cHvTTvyDC46AgovZ3hMx65IFOYNNC+dI10SnDjC+i/0wy73HXDy96d1p
0blDEPMgnXD6vOkeuHn8+oNC8CjA9KmWg0F5FYzEoL/pIrnrN6UyW85BhId9vWE7
YUXY21lRT/AG/asTwjscUFl27K2oKY0ocOXVA587EgO/LvL63TPudLQrR/nCsp0L
8n4yyOgAQlNPO5xhXEgzZYwoZtAgVbi2WqRJ6G/C3MlD26O4m/xBCuEgAnaZvwUx
WGOUk6TFQPB69kYN2Ppx10Sr1cMxCirtE8Mqxf72G2Ftv/0VlkBQI9PB9ZQpP+wG
AeHARqM8cmkHFtHsaB0N+qh3rISUxmGYgkgANF1HLtzQDxFAm3CsmBkBAzzXFGL+
6fuXs9gK8FYEhflcYmGnuHw0cXFtJYOR53LPA/Og+iomdgGs4Olgbx4aK8gujMJF
dTiLOXx5/ZR4F2ifNmARbn4YrAGcArmI5hHwMcaIaYOsGmjxIlKKKLSLbdn6AMpK
TFgKraC4gTd3IJGqPrW8CEYkRNmsjCd/vrA2M1FvP2J31IZcd3j7wPDtxJp1lRBF
Ze7Ar/xJKShV+UlvvAKKkergXO0l8su39QaF9p4wI8ULCj+0AimrGMkhZihPmT6X
FlaYybR/ZxA0pQyVyS+yQw1IO5XIRGEfu4GT3dozyTS6a8flCSydFbs4v+fhygS1
O5Ur4WexQHh+xEt1l5ClSLxZMOsUcC28en1fWTF3INbNXkdC0SvM1MRP6Hpn4Rke
LIjL0wFQtWeR6ziCk36g3Zm0Tcw/TnaeXuzjYL6CP/54/Evvd4Hd1x2gBvnAj7/C
lrjtVsEnKM9YhnPd+cFDogHnyK6Hz7szh4VqDuzz1eATpgi7g3ZlGWYk9drghAyU
lI6RQo5+vaX+cotj67CwnoYqH396glxuyIGQiXMP1lAjEMYNesJp4QNbOQ0PCxkH
t5cLUvTosqeUcePUDc1/5+CGvQQXG7CGkBtQhQ17lAiHCOHsnM1AE1G0z9xmhdVk
OAXCEWNUXQP2Niz0Z6dAgmPkv2P+vcQoK4rMe5eGQ5JIuRwIXoXqruZNlVeXlV/k
oQG8O+4wjL+jV5lgOXTWf/zcrTGts76wUwWzktpKd52KngCoDQlISh+KgO1cuhum
Z7raNRTDfvA0gdEKCojRUNC74Dhfzr+smcjJKxS1Rl8BxjZ8FRhyFICzUws9N6Gi
ZcnHmJ63juCJo77ihZArQqUFSdDmWRDHnXAmOokLVr0fqiyBNJ8VJlFkgeFAhz9d
fS/nMW+/xSC1IpdU7MEKxeROBevJHGV2eKtBUvVxq783rJpvuWMN4Hqw0uGpW1bq
OR0vmQDgZpfLvyFrWaKV6Wg/JXBB5CJUKrFVCj2fDwRWOCvoE4fJxyLETeHxHx/R
PavkhMspC8lZOTQnttDVQEqq9xw2at0HcSq2FaIYNHh8Vd8ocDRX/y1JfkTyi2ZY
9c7cA+Pkj9Hqtr8KE2H7gkPD5pkN5MYRWliax4NOSr8/oOR0LHHBFpmXYR3p4NnD
BpEq+iQRYUyEnN+CS2mE1SzeSuDu3pB135y51d26zRpB7Y5pIa6I2Mz4Gw+rNs0Q
g3ZHLxg+UoZsy8cVNIWj+1gK2s3R/Xi2GTv/vC0gZyREyTzNpEdcQgv272aOe8ka
439K4pdmcH1QQZ12cu9aN3lPADEUs+MAhCtWYQ6D56gJn8srXdjwDiuynnlT/ZaU
B2Hc8H2yIrnIcYpQHxnmf0bqNC4RrXLAxrKBkCOxc2G/RJI2Nfi2WcfjsEAT5qwS
vsZ1ZgfJ2CAqdOIRC/hjAhT/AqY/KK6P7dBWVobFzKQE+wsoYkS3GxW7WDc4OcDf
F6Xg+0Vgfs8G3XDlBt+9La16MRPM/sUT76XkoIDcEAQiZ5C0gBnBUHfM4imspVMP
Qp1urnTyteypxrOr3swrsZLm/2AguCR/pamay6evPHsntnPW8rU1rdkP6X7bSmgU
lG/B3O9sQ2LpefJ17i7rEShiDKFcZ+mcBZtXPwmUTNhC/o2+nh4txbAQeoqwTXeP
pN5I6RCGDxwqfwxdZLVd/PHyg7fxBxJ2GfXIzxdsH2wDCcsurC5MfKKJrpEqwW9Q
zIyVul+ismQHjsyASqxcDloV/7mxVUog6Idb9MCkDjwjJ3RR9PEdENl237e2cZP1
tBm953TCNRw0HYLFz0vwAoAFBW5RkqIeOTLvbUWP0sQdcpZ1TqC94ZPDQhd5X3uX
5rJht0w1kU5OQ7isJviY9nkiiYjHWaUTask6zrORCp1CJO/S8VwbnY9wnI0Gyifw
wt7j3/vTFPvPimE2mOjZbr/z1dd6NbQJXI5j5NXsrltnU+7lNGTxBAQqFdK6o4Vw
sZr5gYIfd/3XZ25LHntvtOL/b8Uo3sCKlTLGfT36H3Mpn3J3HpnHERUGGsUbN6oY
GoZvdDMZV0fGgoi1XAfox7jcc87M4miTsiDtnh3zk36Gn/4f7pexWgQgsbJheu4+
bhRlWvHja4sZwsYeL3h2BLoyJE+pO3cRFlaBEJiJFLp3X8h9sb3ZxOb8kS6uV4s0
v7plgQpW4SqNYUYDnStndhqEHKSgs0suPdb/y9A4J+iI0iNTIpwDoEuVbwlveAWr
H/ySIIamF2YTz486kgNUmr2clBjPqFDcLL4/V8WounH8EbVixlrrAEe6qYU2tZ8K
scbKwdSwVwJcMFowIxUe/joH47tgSLUaS61NlEPoawHAklI9DuNJlhQ/qM+hideB
013jqfPQu4ubEzw/is6bEM75/r1xvwP1wDbYDXzvKh1kYi3nrmyCyC7wtIylejNc
1xqE+D/vmx7ZQ4Up387WkQLNpfq0gEFmWwlKVfOmTNB8jnH7lRg0U1ZhFzcadmPi
/fpeKCE1Sdz2bwv4E80K0e9N/FsZ7ntSQE1TbW/8bt0nkPRzQrs3hLxlw9nNNQE1
uQ1WY8AVFa5qNOCE6wQUaTw4bCICWopGeCRtC7Y8z/nfz4K4at7kgYz2PV10oLuX
PHJSCnZyEvUIIc5IL7PNADTaN/mINUH/xW2s0BO9I4uY0xWlVyTOzPyIGVbxZ/+G
nMyVtVP6ZBQ7B/xiXW8yCtLgfg4A70JaJSl6gj4+dYoF0g5RsOVoxOoNls/wpKgX
tKpuLRJ4dRq+nprY4YbUThzwfrjIcZAQy5inglalrV2oigaFXRGZmrFMTMR5DSIg
3ncV4gBWa0+d9zU6xGzX4QfwIaomYg3u1IOTqTpa1CTSDi0xPgXkvVsgOea3mfx5
JrbOqcuaFFptXfn3NwvSGnLXAvtiEmxNXqgukzfo0wuYxEx0IY0JQjeg4R0D8vIN
V7u0xUihESElaI69mGUSjiNGBkS30VWrLXuHbmXQIcRSTD+yT5DFdmcajVoBbQyD
t9Ae3pm8JLT2kxhhr4M0N2fuEQt9hy8vZnqn2346ol3hITL2U3vbKfNxsEx/ZEOH
Q8xBrwIe2aunBIPFC1vEWOFGB39C1qOhK/N1DIR394Ka1tNEyENc19a9SVAD2tNp
LuYbI6BOj9cz70fI1p2Hyi7VV2SwQT6Wp9e7GKhN2WviIkHCd78WdIIVcnr7sgCR
zJcFTZl94sc+14agFT7DlN2F/pNR4FuRM0u+q6cEHXsprBKrBH+SAfcGIcZ3EEZM
xNxXSaAoW3muAaV0ok9VRtw96RN24cyzfepusPRphEHBtPStsHkv6jp8Gh4+BVvl
jKUABy+le/HZNV+cxDNdSylbPLPYpyxrR/xH0ceCTe5k9ASBsX3wvha/Q8ISGCgU
Hy+gSUPDJ9/MbtD9eOsH/zb0DET7OsfGDSArt+zSy74KgLPylcPZ6B83cWRBTqcS
ug9MtEh547GWrxu1ElDKUKC+SsO6EhwiPEJSMuhCRQfMmqvG1ffLnEgjVVpI8Lo3
OsLT+EZPthCkpJYyzrLFEMibr+Kyr80RWL2HE9xNlp5lmBq0XbWndXep5O5qUwco
Vnk/o9bdGBnA95L53o90t4lPTLAs7W7PORvsjIYYcot6m1ysdBAbM6n7AVvNyrTJ
uRAH5Qt7wtzeUzyX6vrBH6AaOQyU3LXLydCkEd9kOlPHo67HN1FV7iJleH/XDklW
iUTewsXRETDejW3QBXPPu+e+1hptWcFXuYFXWOVM9dm/4qEc4vAuWVw9gSSfnGhh
ihF6e5g4DAxMfUJgcCNLagYchlM/qZ1E8Yj0kIygrXNY3XCKMzVeOFWeJVrw1mcz
Wf5BOVGPL4SvUJldUXIGigssIvsBfnMtRy98gB6iH5JWVo2+l9DFYxR6CR/PYW/s
kHKhJm1tMurZgrei6QM+7jJC2P4kqvx5Ip+95XkGpqT1MA3tgHmr4PqhdN9a1Cfc
v6/w7tb5zHbIHM1pONpI7hlxtFAy1q8839CPZMAKyFgS9y3WOKDotoDOVN9ZvVmF
SnyiNoqajaiuQmqtr6ytJvvCEaj8iQsBvBWjitasYItv+ozR2eQsCo2GMOE8wrOb
hP9mh98rM7J8WiiC7yXFOcLRf6NdY39Zl5wLlvEr29OCTXPzDXAdUVTL4iwOem9J
DoGbNHGcZEIkxRNMc9F47U22tHDpGKhgCC8ok5TnrXeP7zQAN3maQuNCJTQZCbzY
U1D5L3fHrZcBH6GkcrLWHyHIS253CWWDwKfs17NZ8N2k0MXpuMTqgj2QB2hmLAB2
PC8Mw4ML0c6xVcACSbdO8TeG0kBgMjONLApLIGrL44pK8OWg9Kw0cHBvlfQNm8W8
A81cVUSTt0LlXL5HQDV2AEh+CaJ25VXae/76JpX96VV3eKGf5egnz+C0u7B/Ce6B
NlFu29BZGGtmhjWn+b28PYgxqMwArQnrbAUyzYy4Z3ctPncqCjGNE8TjgwcrQeZz
T3rAzgjXFVEUxacMEhB/fRJBmDh2h40UHF6Yanj4/EzMo3hGQkE5OHcLUwPnxb/F
vtoJA4oLSf2eWKO9geHP02zDezETAgH/ya3pXKYHoTWSZ5Le5u2b1k4YQZPE7An9
419CgZk/d0cOwh/VN45cjGHYBAcyydkgh7CvfVlZYa9SpQ6Mksk66gW+uslb7QWs
Dx6fxm5KFGzEhjTsSHIHbzSa360G26SGGD5n90ZzqQ9TD1EOHqzO4iQ14Rl01OAd
SK1bvHCvQ9QAA/PHiA10IQ8HWpkH0SKyU/s5QcBv/ghEv1G7XKHdNQkUHD8lc68E
nLtImZ6Vn3jdxVu0+c308SN3rul8ayfFlVR/4yPgN/GttqRpQuh4kqnKgan0s8cz
kbHJH7F8aqnoli1wr3Q1Yd85C6FJEDpN82Hjkbx89SlLSPkyZF6sq1EuTvq3BTMT
GE+k7mkQt8T1MAeYdtdEX5rbNgSWWw4DMdwOMdGF9PhruAPijTDORVJLtPI7CNlg
utR812V3wXOZ+4+DxmRramkMVScb9gqJLhTzWw4jx0y7QtBoBEQepXUT6Kihvik5
EYX0b43uWco7hn5X2v4LXlArssq5HS43bepBRsarM9goaLQjU8A1P45tbwMZRoUc
JK9UG3ckSYd4+X858eGi6thCefJ5e8Yjh8z7lwcLNA9P8KDG+hOWbHNy5dt4ts5b
7Px0/0HJlH0kSuFpAhVNBUPsMYKMJ+vOj3xmhq8r+DFAj1/7Wto81kDzXoPuyLy0
jRu901ylgxVvsNTovp9Hv7psMRXsS/iKC9S/bYMvUcXXqfb4YOFMLtEsVg10x8u6
mLszjzKvKNzpYClNODa9fkzru2wAvlxQUZgKWSL+gKqMuOzTvhVnQ3bIbV1mSVpl
o7qTt4NASfB3IQywgNKKV19ZDFdaeUzTPvm5R9DpTZ39eLEmrhRWs2iCEDf7BK3I
EzvYWCIj4NojjrvKMDHvTKZD8y/Q3ijSOktdpQRIwZC/+7u1sreFtu8FB4ZSLAFg
JXkBJ+yZXadQ9kkkEH7YuP139IKXPPxWYgxFmgx+uPNzqiiJYYqYHvqaYxRBfdPv
BnKSHe5B1wrNXGwt+y44mp5D2W3iPrxjBJLGW17IXqxONrmkKOC9PaFQgCQKEZDp
qrQhFmReVmLMuKrupz3A+KRy8YaBXsWdyNy+mfyoKrQ/GqrTU8ENDZmgtSabhV3N
e2SXA02LHPuiqwvI/tSDfjLitc+23iTWfTHvfRfon0te6yW68UvTxaErxtiho5qu
qNICc/53WF6z7L++4vWDM02yxJqlm6REBkisDL4X5yrEcrKIriAkRZHZbvHIRIQ2
ddfOTmNo6z3X9jT1IHiWE10Ur/FiDtXuJmPJWe6JCcPqZ2G0DsucVwc133OS81ZC
y98RwLnM3WMu6dGC5bnrweJCosjJDN7uEJtBF87TqmbZPOH8V6c6vYxFgrA9KlQ8
hSko4i5I5yD3xNGapGRKRPexaFgmiwNVz4oJS+rtwR16kFuQEiRpqg2OZwEoAoWn
NZdHDFPw91avpfB8mqoVcLRjmzY/uFaO16OLDNtOSylptj25VM4wWyM906LVNoVk
77ewZ4cUSVpDME1L4FvvOv3seP8Ys83qgPRiII0MHzegUPCdda4tRfZyGCHIuuEW
Kw8JkRcclCTwG+ZvF5eTJSl0kN8ObmH3eOOLJIAtl/tW7H8Q9F8IhLKIvJ5awMRb
DeE/2j/bk6fPGMMsCiLSj97lsQ9o5vi4utHPVRLCRX4+t5LqBs+FHjaEiGZv/ska
4y+xaHcpdzJZrOD4C6H2g7t7Z5N5Sz4b8OKu6AbYOaCewPk3o6DpwK8CtLSTxKZr
EmH5/9d7kZ2Fy022rnOwyqS4luRgEEOQL1lCJjJpbnlR4kEryqWorrgTu3doQMjc
NqQcC/qVF4wqz3hXKMcXz0hC/U72SsZPc2l8M3PrplpCbwm28i+PG9MMVK+nx4f+
wmc2OXJyc73nZ7zeFt5C+ZT7eC8Mc2D20Wi0fcffdH3mwi5r9jQlK1OJFPn0DjdK
IQCSyRHJz/oRKqvTvjDd0pLwdGCkQyeyDZDVRaanv9EavNmbwcKYaZ7xE11G3o4Y
mqSlIE2SH1UJKOkI6+ntkJ3pfJ6UNct9dXNxNSgrPEJcLkONIIW8eonTRhD+E+z8
9R8T5Yc4RkSRkGyK4oIxIQDoQovRjqHpZk399v77o5huQyZXkl+EJP2t1lbGp1YS
UxISTPFEk5dZqTYMbu08ElFDWPRNtY3r+upWvNr6UFA+slMvsplzstkSY2EvdjN2
yVssp3Ozbe9d8AxmUE9DoCwz+wZH4PSWyUAf6UfMnJMDcRCReFu9rMzTHPpl5z1L
E/T/Ea3bXDVda9bVXZzGjDR6g7+AmXtu546cmd5UbzrVTyZ6fkVUYlDzd9K8NOsA
tgyLHE3y2eo+OeJ3JGk8sBOmg8fzKRyQsr+ueRqHLLCuPZ3dgrXoJmlxPfoGT9PN
DlkTIp1zknz5Ll6AUtr70TTd/y3TDsUXm+xpLlqV8AWaSjEaHRsTRZU5uQqdpWPE
+2thntrqLJInoo1EksvmM2L4rIq8Q10F8z8+6NOAaZUHNkg8wdH68/+Ypd2VOUqt
Yqvs35V0QU8+0u4KRhdrSGlh576LY6EyCZQMNILlDIEsOYTJyeyizFVUh+r3mRNY
+4UDfdKuOVFjORI8UgDiu0Nu5QUP/hnBSl9ZBQrSoWWbbRTPEv/Bzy0iaRrSa2bl
2g5QThk93ZqtTsElJNus0G04zwhYvtP7sk3SNzQA1lhmbnqZQhXTJ1Drntp7F2ev
7Kg2YpR2xJQ0YCnpbjcTBu1/h44tUNnCMqpZmIEaGE14ywpTKpnMbOfTE1C4SozI
wlScZdT+73/hDl0weUflbCMjb1EZCE9BDRlSI1H5j0U5t5o3hC72+Mx8jg2sJSpd
/0E3MwRYcUJrbZNfx9H2olLzlDwjm2X5dhaEg/2ZyifI5pDQGIDlkQ69VJv273A3
t/VIqJJm5PaFl4V278x0ObC6f8pYszAQ1FLTHj2b6aZgweRXu3lH+5uJtHAlyWPN
rJCu5kluch83l2fAw0mLgs5NLSzICJaxZRg/v5g9rwm+uEiaMkQRWTu19qVd47Td
ivV/AugdTrjKs6/gQDF3bgW3U1TQ4/UctWKktnKcCbeF0iCKdK44SYorpziimYGt
YoDi2GkasetRaI2yWahhqRccTdh0NIpqqKGSeOOiqJxE1R1GWp+SLK1BRwnPoS6s
K/bk5xfhPm11YWSul5XtH4BYuYM6ZOSTDQUwlNpAo+qQYaN++frMJwmcMxinqHDs
I5MYP9BLyV3Y7kl+h2WmK0FreZEPJskiMQZnQsOfPAsE8lAnn2aQ6uAPFSiJY9TF
rJPNWypbjy25wyNn3lgnJQZ7rWShVGDHJ9dXjvMHTYaApi9PfBG3dVjomSDLKn3F
0+CMftgspyAkrBEa2oSkf/w8jFb7hmct+kyIX8H3ZyEFUiuvy3zj83pKPJcJbr50
Id+MAN+0GsQ7+1BpYuxhL8VkOebd9sNp3IkxIXiBa8qvF5Qsq8Idnw6NcgjEwM5D
iaPHP2zmfl1hanyN2bi5NuG4nJemyIW87Kd9H3mRojeCPuRDQLRk6GJFd9IFvSHi
t9G3jD27tdvClvAeOrl5g8YMyMsWaDADjAWwVR1yNw7wSjG+mi639uawYrAtS4xu
pwHi60ZX0zgcfi5J49VBRu52evbs7DPwGdUet1ss32wdqw7hxe9j2zHlvi+t4kN7
EQGAnAArJZi7RmJTNBfHBBOfusR5grqxNYwsNQV4Ys1c8Cp72harLukeCtYXVW4V
gJqpN0VP7yeENYum644xG0MkKGlKfZmurmm2AD7Djxsq6Wp6Hk6uf++FkC0a90rY
/zqlCw0zckMb5zxTtDbX3SRYp8KZADQbZtKK6dDth/G58Aj1nJVlgXl/MvoMyE7F
ZDppbQFDhUF9fIcX4kcHV77Wn15ll31oiBfl8p7GAJg5C4MZB9MYYR1oyf8B1kTL
WXu05Y15qggznm3isCkvbAi4T0n7GEiQuOGSJ9fwSJAPLnEB+fAiOsXuBWyG3XO3
3qEeTbpRqAbnms7S7YeqXdlHlUXLmJhQLtHVETF1zIaOfDtqHLDgMHZhQYoRxOKq
AR76AGQ3OISXXw7PSoivSC5eWNbs/9ch/siGsjsLxaC+1ksfaCQD0r8vk8QW7JEu
nc6B4DZFo5LED6vcO8HYG9nShDHDDXcUg3S2sN3UroxB9G1rjwZcRxrttFlmUMsC
PaYzyP3EHh+uTlRO4sbcsCAZpgoHuVVoYOCLxoiTBe47EYMG3c0U+ASxJerz1vs5
Bk/QVtBiXAWymc3aDzCrKjuEtaqyjyokuZJHIrtC9AEeoh+i/zch57YGu2Xv5k+r
9u7EIaWHfv6/qgIXcRUxwf0FGON0jwUzLiFXR6JsVuktLSB7S6lS3yBCa9xCR7rJ
imx0gxUJVlPahaA+dotxyrHp1ALoEyEPto/EfUd0V3fANgL3NTi5bb6JiQigV328
c+Up72hh/Tu1YZWOjai41aN4sU9D7DRYANExXDz0ROAG7xOn+vESrZIzV1gKKi2q
QYAD2lCika4TIFnfkb8at8T1NtIxqFRtMd+TURTygkZ0rNv9/+JlSIdetIRemaFR
dgb8OvVqTFnssETAOQbuZQUof67OlsvuPE/4j4EnF/gpaDUKgR4P65nw8+KlmcmG
zZCxAh9KV/iUd/YJ6WXVnAu2U6FMYT3Z57fIr6EURjmSU6yj5tmIAXeT/o3Wa86j
2SqQLwKE4SLlZiCXl90aQFIfuX987BQzrANbX0kvzqpuqv9Hn47AGW5WLUGyntKy
z6HSj9cUufrYMrPxW2NYEHl5y2nn27U7h5I6+D8HCOcu/PPPAtTB1u3UPhAU81yC
Kpva5sOYb8kfD43FHkCN7SHEaNignPg+ltHNomo2LT/i3NK65hz5i/FXFfzNXwPW
PWT/iKDBNdKFJ2obWzAMRACsNK/MWqoHS7oZ0uFvW0/BF03Gv+0hca+6BbTy7gSK
ptEnXG7YIktDHBMs5c3se5jbQJxQ4pTOVjsExG7Amsku04EL8+7B0UCoFwboMuPB
qFvLtF45HB6SR9jL1uS8TNp+LVZY4WL1LYmJBTqKjwGrm2RNSEZKf8u4z1o5zJu4
nvRrXWbIxL5eyOsMYhpcR/meu5JrZ8Iy6XCHyLelNXMBQYGfrS2WNTjnX+kc3bMR
f3OwdIwnc8dlDdaY41lLpnUofrBtYYr/oFETaepBW4f+wkoqNhVkV4dij/ZJ3yIn
2FNBzMs9RjF/56lVFwmi+GeNkuWF08PqeGy55PZwn9MP6cMlpHqHkUddoR79yMLF
8R+ndQrD6GCQ/I1nN9moAorpTqs2eg/HyDEn/ZEuFGs48K7yJTumWjmV9bYpw2JL
FMrgrMT76h3SPkYFHmMx4hS330asFhTdSJGPpQ+dZB24lVP/TJ8VaInaf3PNNVBW
qIsbubAQue4s9ALEkDKzCAu1I8gQFyQTDCTQntOGqeVDFwXPlm3wYKOLoC7UbCBC
DrG6NwgBgySKCsP1i46G3AINyxTK6r6V0IjK3KdDx6iE7JQffUb+2b+IaDwuKSEF
QKM+UwEVvyfb8WyPAqpjk2hooP60gJKLKecRBXizFynNVelGfkiMrckhkcv8w8pV
t2O51FWhPI/2KksQ4Dp318hqqRtPNNIZj6eoDXbWSykGUnxeqtYw0TE1keJWK6Dr
pV1C621yLVhNG3pO4byZbry+RRr2NVCdihoRTFqxr0mTEJrkiUFgKpdi7Vf1EHRb
feznwQw/6AqIbOoD+jT3tPTwNLiPdQ5UU7tSbV4ghY67f8FGDQ0+N2JxwUSYMJfu
1HngBdFRl6PFYZVADiJPEgDX765orTWEc2XdSByoNHrhDBuKbJ13tY9k0+biwVXe
coF+gxsSbux6QM6Zu6bK2gRp3SU8f/Onc/bWheXwtXs01IfJIBEYmikMLp69gZ5R
9lK3KDymf7cIVh1dz0d8PjsQoE16RkjiRogXgddIA6t2zxApRKOkvXbuLZVxF2Vr
KjSokDNMITN2x9U0PxJZK4O3pTYQV5qDPPjGxKm7o7mPCpzQKNFHFxVXuC91vp4m
n5bBCc6VWAJSIzEbhOBzyHIF0wCWqBxKrN3Xu9dp4P2ZEpUe1EFEvJq4s/s1l/Y8
NWTvDemqIKwvNYUQSZ34cKQN3UqReSfxF5+LrMrlfhhz/7JeMtpUnSvcHr03v+dN
OByeC/0ddcTPgT3WxW7g7BSVxNxMM/JkyGW5XnGqkVtiqdaZQ86Pvm975csDnrMK
f94GV41+EvJo6sdITCL7j1X+nWAhxthAFKWZvWcwoQrONL+NRXc1Gz31x9x0BEke
AGzMkHGccfgs6g8UJ8qnJHbFaJZHO/y96J2s75D8BsqOiZAru/Ny8hFb9sdaIUO7
oDmHPs7TIOOulX4jJ/ssHDfPhUK8zGXx8HW3MZ3bpMRtu92AHfr9eAYfYSZDS7Cv
XbJ/tmvGpdKPYQZ9rlGT2N31+PiALLZDnZdTlF0TydYsMb2mCqRzwoiG+r76WeTj
iDMys6mKYrWgbqXk8tK/QTcbQnXJLR5DvFmvpBM2XThEeWy4N7jWK8ntySpkK7MX
bMfm9brgl+Z+i+J2DyUPaNIoUXY7XpNfSj58lGEPbR4tylv1TKe7sgmyLKnyaq6U
iEJyVELutJPGuYt7b9FyFPeKi3pwk3dB+AyQcywZfXk7KGK/UZKYrzE9g6i747Ms
vwZ4WmRR7zDUVz7znXQTSiFt+XSrvPMtv0/C6va3w718Bnj6Xpq7QgnEKLalrkrk
hO0IaIinpQJetQ/jD2VROyZv38XA5hjyexfHKIPiKt7GyTTV8OObgI7I3oNw9tNm
1+voWmjPlZvin6qftHXVigZPwoYbyS00EiqjpPm7ZovTFsQrTZMATnmaMtLXS4ax
E0+mS0ZSigAOCEWVKVFAGV0kmj40TuImHZSTy1UeNamSYEWMGN9B8xrtwMrDWNPb
gK1FTzPJtvrxo7mHN4iQ2ukUAwmQLAOe4fQ8+3L4ROOQ5peeN4NT2Xla41JJwUve
LIzbyqlC0zQvZlxhRwNDHAjbnq3zIqobuh/Wmb8qBXBmxCjixnVUh8KWwZO8Mhhe
//QBYMSYWIGTfW5jBHeKtCFWm3cVtRAIcfosp4Z+GDcoMR+3tLKbEh6pUZ7r3G3e
HijWo+UvXKadcrvrcetvGzQwghQ7QvuZindQCpnJiF4+ksMULNqN9GycI3qXeXaX
vqOpYbBsGW9plunElTZ9bm7/AvQTjIqmCDazPSDjB6fqpvlwJmm8atsdXN6LDEQ5
+idKKZpyZkjHgSYPw/+x/zps+MTir6CbqmyBryoQRo6hB6EDY61wEzW6baAeaCfV
JlgoAOvsutVVUOMCP1axldyWZJp1bqCkWNG6tuSbBAS1B9I2YpietuPwq2dkkDav
bM8kYNMEkIJ27zrydPwdAnQYAuuLyFwjK6ex4Pyawc30OyoySEMhutXDAf55hGVv
TBq7nA2BBix/TulpgHyTpVU9GrLv85SCGrEanDUmfV6+0MX7nt+GXeD0onRALQQ+
Xux5jFFa2Yw61JHFpKyJDsTEwuI2V9L4uBDnjTK0hJcraxFtn975HKzkGyu3yGgu
aVxa8wHuKOlsmRStkpNZxwF6cLO7oVw51xHC2JrPWwfwPI47zL+N3beeHIrtTvFg
qsB28sC+1q8o8d5fjKTQIzf9V6hWY3fsjWOF/t4ZqgoLzXBRpAWlEdvw8pErCGp+
+dh0jsoevx814jpG8OjDeSoIjwJc95AgqKf6iLx0oxRlqMwi131vc6szN5slsSgn
gJrp7FTlGd2VUKSa8EDmGwXr0/lnp4mBlX1dAF5yuoEwPVV9wTw4W1fO359iT82h
7wLxzeHngTHX4pEc6QN7j3Ib1XyahF3e1BIVxV5n0030uZQk2TbK44V8m3LhIE3K
zZhWADQGni+C/8Mh0+O51NhZwpr7ZO2FIkAH0+C93M4ng9Z4AKtf/eKWr2gm9ZKT
ZlVB3FiFMiEFsvvh76ZsFWVq80fQ7fadbfS0AynB7qBQft9BxbSgdctora9Tj6js
Qfce2dST+8vNnbfHDaarydSVC6za78YleatscI14YijkvSOdjpcBeZbMQ8Ci70bw
hlKXO3b/IJnI4KML4lMkY47v8ogJpgCAvYmVQ7nhqDaWlsgld2TuQT2s10N+MFTF
wlsO3bYA/5vda9O3dP/uPFmdryGrYTTNhtrUlkqyXDyL5KuWRAFRlgMwl083+xdV
HB4uBirX6JSC69Peo3kcoNPyQjbjTp9Xz3dvr6EENroKRyTw2GvB9Eb1FdiJSz5u
8ocnF9mBQ7vp4O/LKfaMCeJjLTTbePS/BCUKla72qP8Ep27avBt9Yn2iUZV4x4fu
5OMbPL6qdte/GJ35BwD27Qo6vV7w9V4DP3RhgXO7Ay0JJTQSwwLGVubSaVj050Yc
PHaWRrujxDKPliKRW1NBFlih787XMfK3DMTtTqrpQqHnonVVwiiFbBzYxcsr4mfp
58tLm1TO7BbOcQg18pJN3XIbWf1eUlEfCNZSwlCCgGq0qMKmlNrVkwJP9A4uMEXo
erbrgNumU/8kRtHQyviKJd6zJQWHPrktps+evftkgdPRTJgwrIoywd/SlkNoYO4n
tO4yyrol6b6kygdgIkHld/PfF3q5zhbcpnz/dg4NIkD/yiPIltj530lB7i6sVghe
NB7wnTRP1UvdPIXzS6g8pMTz9uOg8DXbC0qahPDISt1flKco7tKqY2rA5KpZu5Bj
qh2smG4Is4aOPhE5QIDe5OrTaWircz7NoNdow1xYUlUG94BPVh3UrKq1vcY32iqJ
8UhEkj/pXpBnTwtTDvdoVZAwjzjNZ0aMtcmpZdgzpo4m/DRmyfZzcl41EuOradNX
64v8lKU92yivgoSWnAH5fFA+KrYSA1iEi07nx7xk7cNVo1y0rwvS8BsLkA54HHkD
o5JCtDSnBcykhSsAXOPMheICAG6LHo8feKkyPx7umbs549wd+S7JoH196EEld+yh
qAIPkNiluyxGqvbmZpLfGDqEH+jcwaLwrBvs7Y3C/38YbF6WXNMua77H5KRRyGJ8
4fxY0OAN7NdOcYd+8R8p2SSqXAptJE/OQpNWqXaTtLeahx1jcJYWs+KLqhy+4aqF
IfvAVtKJtkiECWLqoNVK0voEseRRSmuT3rp2oAzvB3BUV/SaBwOePNspavxhWjUQ
fG3kFgC/N8UetQR6qc44JMFVsF/9SLj+2mxhWDhogoe3h7ZG+N15iZyQJcgw8eTV
F+GotpQPAnwT/hj/kA7nVT2WArCkFtE0fcLEaDtbPwUjTdrHeIBdhAoYdc++uzvL
uRGM5soKE7zgwxSFOyic1wzHe12+GSThDxmZdXjn9nC2/+BhlwbvoACdHnjsyiMu
I1LbEYiAIHnWPVYH6O8+iY7A8iteC4GbCy9bYh4y/Q+Rb+YMyBXtLcmuGnVI50NL
KhVCo5r4Dux7Nd648wtMV/TViJk0AByA2Dn2Q+1mGk37Vorpv7whPQkg37+zPb5v
H7blQI+qFIgKJ/V1LLKWQ/UEMIY3d+yMd/qroa0XQHSawTRFYP60dzJ05Z6DK4Ts
TEnmjyF2A4NC9U5ZCF5NjVv9F1j4E9N8nJaWDX7Szir02Hf3jTALTtqq1duWnXpq
CY8TvmPkgJqAEWkRSq5fO97zAr6GS39D+qvdVejfgmbJ7HDJwqJkZ/n2HuN0wDnH
xO4SGktkhAC2lG2GrD4JN1N+q8gZRYfZ4gayw34Ef+Dd9EouTCgkl3fM1jmdZjiO
I/ZhAinrWFckTEOtW3kE9TEydidurbN/1SgnlvgQgmOChJpOIhDfFRkkDQcTW/Et
V75XRwbyeoUV1fR/u9BiSwUYEjJw11e8sjyoEDWCk/8I3A9/eydJJuRjwkzS4zWg
vQDf4yWnkeTNBj2o/JNA/xbJFAt5tfsh+SNU2sdvnqY9TlHNnpHIfPkLPlsFhw45
cjlU09yEy3sjy7owDISMXsXrlf2EAodw4WsUzergpuQE8l6fE5vVlrJlAimnE1uv
kPBGGGagmsB7fiWS0WJTFhp9O734OSiWlnMlMl30bkYfLlmt922NygaVimUY+8AP
yWhiRSj20/f6rs/Kjd+ovHiwPqGySR2kPHrCShmIt4lEK6ynlY+06B81xlbuVv6P
0kdruzy1b9ivmWkklPvMSVNA5rvwaR4m+AH0NhNeb0N/zBzbq4SSbnpCKRbjVN7E
UF2pI2s0msq5zqO2QWbi//+Bdm+9cjDnAHr7E8A0xuc+dIHlIQM6KYoNSmSxVyYK
QpkUYR1Ryr/ypDdRPvn3xWigFgrt7Nf4QVaMIO3dc8BtKehs/gt2Ht8dw4ykadEQ
jmhwZF65tiHPvCnAHcDurWgim+ICRfKthuDFSR7YGGaFWL1rwX3w653O/iW/3GR5
/RqIKyOvV5iYzUb5naqO9lb8HDJy+r5DLAJVFa0WW5YimU+PXTqcn2HC1pPmMfYr
LoamauksMm9qOUJbbBIzci0nJRTvWyzHmsq7Z1Es4IKKl93DD1IkhRZc2DBjubKm
Qd034aBb04ZYfRWbhngUqI/0PUMDKTWBab8HB9t9Q+/a21LofIw6uk/xK1RA/RIs
5myIAR0fcELxpBbK1BjTMyIt/Q3HJPi51VTRpaMft2MMh2zo0YG3iCcfAtpT8K0T
oGGlubjH6vs9ubbx7rdOikAAUvsClZpp8c47l2ty0ejisYdUs6IMK4io1aiqBR4N
wHfORNHVEqIPSz8cWpdELmnVIlKt86NdQujmWPjYwRMqPHU5rm4YSIaKt279WmZN
2nzOLvoIsFuVxspnbAqZDLSg9cH6iU8N+UWR8OdGXcocYzMrCy+MpCPbgiivum8g
od329Zsdc8Q5LHHH2nS9gv/M7M10WSjWe8g5AQiH73r222WiKYNl+Bp9mNf1lb1v
dksULgaqstcFAmIPpnNAo9UwOkCMI0rrM2rNJEeSpyOPBAa7ien350KC/OUKqFnR
8dEge+Auwc399KH3LS5vy43iY6KQocrJODC1O3Ri2N+ZeTbw34YNphBZAsjSKuw9
2gsyjh4Gah2u4VCbNexuWwjhxrhACFtKb+x07Lbh0WlK7np61IliZOBrn7BHJftu
5RXLdf/eccY6jXjBjlNl0OVpYVe6S2eC1ItGhETwZAxg36ZYr9FRCjelUlOk0gxR
AVyTm67HTAucJ9U7rBLwvgnU0u73UekN1MQeNl3aQr0XO+Z/DUrXHwPPM/Ogs6Ji
a+8+06VOX8R/a8ybVusG2R7MStvMvDADBxmnUhboNiTI2xxYopIMnSdozNJuitiC
Z5jzqdaaZpI/WfviMPQqpF3NIxdSefCPk2GQcjWqwKlZKUAmBzr+pPOcaOkrgbNf
CkgKYfEXZ8IET2HjJnk12vLgqxXdRdg41Q6w49BSUp81ma9P/PsteklOBTy0sbVV
5BBPPxhWhnTSiWOlSRFDr5qtrZrKjyH6Nabh/PuUNf0TSIIzmJ9gGqYJlWKJLtTY
Nxy4ZxcPPrCbMQpjw0ZEUVIU6l55yF3l88WVt8gS90YKa/PNdMFaLo36NAnO/ZMs
7cjFIMCgkwImdSuIIZ4/8Uu3Zx3mmDntSvJXTyFn/EkeBrmUjf4kDYBypGOisLr2
De7YrMXrabwtKhK/bazn+wUq2rft6XotwaWrxIA5R6LpWQwrg0+cwwTnGYn63VJ0
SLEhIUXrAe1WGNjlzrd64xhl3WVrLqImlXgUj5x7I6Lzv5CbDB6anj8345uOKyID
FLs2TVchD/SgapGB4Mr8dJZ3LlG+9Ye3+gcSBeTWX6sHMn4eZq64fYdtQjM/rl8s
bzqoLRSH7MJdpD3d5B1fvEjgYg8eJNF8ZraOrGZ2qqajEdovFakE9ZKD6kSGnt1D
svAohm0jEhM1R/cLPdm4aBW3T21LuGpoknAk42wxOfS9wqkIOkYc8EHy+nNAz6jr
JMaHoV1oPEtRzjirSU873duF+eStwuGSs5NObn0QoUkMFpQi0AL10uIXCWCArrnr
Wt11j+fq45xsVcH6dzQvJs5/Q6Z1micGDrDaszH23NQ4bXs5I15wwZ4TD7vqkROO
6fNExQyIi6y7KyG0C3vSIRUJ2/ONLKZ2bEcBLlR2Ws9HQXMYWVwYLyYHrNdedE76
wzzdyfcvByDgVoghBgZgcdq+e7rXysNsU5s2bqHM/FhLHDHsOpmofHI3Jd++owRk
82ut4Vs+gJmLVnHpN+fE3sS5Wdpa6GgeJJufZVaz6qg5inyi8ftEYG+1nMbISRSD
/cKGuky74WBWVHLUHXqeBmkBTIfluhtEQi77mAZSmIexPd9ggJHilykGq9FjX3Uz
2Z8++d+r4cn53X0pYDbl/dsmQ6eYrdLuoFCWfUWBGuYUBI/7IX3Amyoqxb+x86LN
6ssvJVBNQPkfSLE+WowLyqsZMcXE5DxDiSvS6L9ohuSM/SpqOoYxkT2HMvJm4Rax
eCgp/RurpiVasMhUAEyC91PWxEHncGRCbWMm+hw9IarY1WNJABxbPV02WbhyFOJ3
wslUTgMIdGiBN1y5hNzYl6Gulxekag6FJv2lbAGLUGe4bZTJIBQ3JVHSsfNfwjEA
8rt1lv/jyC3u6Em2Itqe5jVGgfsxfUyEJtSxIo+pfFA7Bj6fdwzjAwrTaMfsRW3E
x/RyvDL8QuYT4s0dJRD99JZ8WDe+3LOSZ5lVZZJUuE69L3hZtGt1V7SaGNrFWAfI
XLtSsB/dFWhj7Ol0PUHjMYCwFj3911WI/KW1yON0ltCNd09JDlyMx3iV0bJiqZq0
kGAlNoOTkMBLndEBLTCsyyN2UjTkT5GDHzB/189Odt6AuLnC2KjenKRvaIlNOvda
7F2IpCvOJUg9OLNfw7BK0W0cwXZNRv6KeWYXPSIm8dp9/u/FlDordh1WACzSKzeP
CcPNn5TevP14fENkgIRFH8szgSZW2aGXZz+Jecoa/F01StsEiE/JkH7Lrlt1Rd5Z
CWoKzHYqlnZ338p8Lqnbyz4cSRaaRa0LKDgLbQshUL0Tke8RJXrHhQ0ciMbgRO7t
LTOrOn0gHNHA87buBha5bx2JGkYbbIOaM27miS7NsqP6AtPzH7jH+Zj1KFQ5oruz
3ANH+UmWYzPNHao6QdWMnZur+wJVU+OoC1fL6L414xOZlgIz7LMiSJASLbPWbQIm
t9L1Sqqy1N17fwhgKAYGJP+ffBLh//5Dq12dPw4odJzKE5ARqgAFL/YCXY18m0sd
45kCrKmcmCHSTxk898ALu4Fl1vnMcBWipWNlM2fSQL0ZOKmDgkTLDE5JX9xgEhTx
KPwV8PCJqEryRi4Tgq4Mv7ZaSAh1F5nZY5oqLHMxQDQxJa5NAwOznLc6Ehc7N++E
SdIsmmwwoSW/Zm11t/Ul/8m7HqUfFLflPvoVH4AhD9F4S3Y54rQeJ2ZD5U+aVzBJ
6vrloOcy+xYUO01kNgSnAWm1w3tJgZK5B0WRNz3qwpR5Fm1tRlD27hLe7mEKj6vp
gj/Q2Q+4UndUyr1V1JZ8ZkqtxCciLDVpkSIs5vzm9jiZI032Q0T38qoyoNVYhWZM
/LejNABnJIaTs8LcPtLLMlbh0yxWmwrSzCqAdMtaaxruzk5P7vsNJila1upDSw0g
OqTy1ANjQpatD7CQNe/H99YvKPhPufvKuSGuLpbB5gnYBk4EAkN48IGP2juaCKT7
It0yYFU1+SeXNWl3jwCpghSJmcL2vmUr686aer+/q9lIHC6JJqHkpeOXASDrmhy6
yPqtkb0TViRuo02PoBMf2i+WymiIZVjLFggYllwJd4yC9vYB6DMqtGu1+zkBW5bd
8d2fs/dcy+XT7SJUmmHkcIArqbPwMiY7rTrGxTcUfqUOywfFZDgEcMkAFxvYQTkE
duaIKSizp9vHCfkaig/VdC5OnaFlEK1t5l2fnjfEhp7ZrqD+GUf2VWunWZmOnOBn
DHrNZNLH9daGXaeQE94lyurlpbTYxadfI0UYqXm8aBUUR7AwVo/SOWhQBq3J/0BD
1HCeyPqVF7GCdL8r4AzOrNQmuFXG84yRzVmZ0n/SEsdXjKTmjz1Pm8WV4u9EtPzM
Jr9vBUkKahgisn3HtQEs0VfniIPlDtiLwic0JiU4JdMilI0rfKK77teM1DjJ1Jg9
vUVXEOf31bhWJUKi8iKZ/NZFMDzkdw9oJ5UEcTegvYm8ZZhsdjUEk52ymEWjbhAx
hq2u0Jd4pkNT0aoDD/MNgZx3rYNtpeV5RFhsrh9R6RJbu6s60ggq/DRfbr9Wp2CI
WBPyuNuoO3Uz9oTdS4XQUptHhc8jE3ibSVHHS2RfTlgZNfvy62P6VRsxRNdG4/8Q
X2eWrieFguqFdpngDkXEcm3aIBujdqPq9cqUK8yZGb/UJvrHqL5dJymVzkk/A6n/
GezYuz8rIk3tacKBG9UDVELLbO0S0fascyPW+vLpkOQ3Ymnd1Y2+Wbuncn65H0wn
lAc/uNTBUzdHdvcWwygqd/bcmcaKokRQrKn1H7JEid8hUaYmvYfqZC2zuLeASpDG
1flS5dcbtCS/12poWkR2pLNfa1yrAvAu+0DkK0qscZ6OtxTAU5bkeAOtrew597mb
DQRA8LQv9g3YRRh1W9byb27sbff8P1y+ZpebeIzrRrf1xZbBkvefjmKOU/fkQIIS
BHOdCjbo7YcFVA2x/mAXfj5HyYExZxwjdHKUoyfIBzzcmUSzQsA8ig0+Lit/H0Dk
9/GW4Q6VBgDTs+sC3VxE24iU69w516pit6UlfPO7FmvIMmLltNM3XWcrWTdLs2cm
HDM9VyUW3RjD48gR6w3/6oT6R1NmvWIpue4AdFKajCIXUj4j99DwE26JzJVnbcIN
LqNB6vjioSVvWwLpcJqWWG/H++8pHIWWZ2W6W5D8mAaNjm3/yy4laslc2xXEDj7h
WqN4NVYbDJpQqF0+OAnP0iqkVU+8gd0+h0BR+Z6uo59JKdbJbzwWwykQ/DlWykTM
sMrnvW+ilDvB+47mQwrsZKWFhAmxXNsEohhAMXQsMJ4l+lclZO3i/rilHYC+6IYX
T9qdHtdRm+j7IGNsK8+CPpM9zpfhSMaqBGHIZrRGOZllPmYHQdr5dehM9VdGAWxZ
wH6KHj+3YDms1c6OLjexW7vSv9O5zlynoyaDkD8KA7DkM4Tv2HY6zyx5eYJQ3yah
kf6BrnGpZtl+Sr3KLC/vHIjMgtmqxUFy6ulxli/Jbeez166t6HqQrD2XdDPBHxRZ
P2SCAs4AKcP6hx2j3E0cxesUa2CTEVO8qFj7EMybc+VRdyPy2vvPtzU51ksP4WVR
RCjoETFDqYj33KOuxHM5TCAwWq8FRYT5U2XDNfHLKK302c6tGEgJJhG2U1rZFpTP
AEsZ6VC9rTIGbI4/FF/fgLI1b/JNngEi3F6wCA8U2q5OpJG3i+2h2syxPlfnu/s4
w9v3E5DBsSYIBm1vuxvI36Lgz0JeqqlFNsbn4vNwi/FWNnVdqG2SnAfY4lOjP0f2
0hKnruOSHVjO2e4ITWsgAQp08Oei4LGjpU4i5hBz78BnwlKTpYA20u49YJz4x4zG
hu5Ckp++jvO+Hv3JwCw0s4IzdI1j/CLwbRF0lagYMpYiPJCwSgI38GZvtMYCOyf2
J7yUC+PdtL7kPOGlaFYGKLbhjuuue8pKC2nez64zFteLT6h6k5glNnUp8Xd3mfwZ
onTKlEJUKDLvqGTL+ohDOFhpGJ0RmElDZMLx6YZ9heupuxVZLz00pwMAFaE2sJco
utW+NjTX6Z7Zyx5RgMZr4QiDbg/HvqvFswZzrQ4hPw2ny1MGHToykWQzlTuj+Qpo
qpvPzRMVo4I7Tf3Bwu/nfTtCEzMhba+NF4CbcGkAoqldKBuQqozcnYjjyVy4nZRq
6r+/Gfgr3Qwy4vRZHtVRleeAZQgnyxa1FXQ36rLD4yILReQTPSAYFDVZ2YmtIO58
AsF2ITmqce1UrhucgKE39NoZlQ0H5PVZ5cRtc7ojyh4/yhg/PR1C9pcJ/krehXwI
8otYuNUoeHdajHh6lPnW50kgz2Tu+iFH8TEr/AXA0FA9ETtjBli4kBmAPK8CoTmJ
QbWWVrVjGYPJuUGIg9RlFeNGYAEz2o306RkpVNCnVo/da83cbpZa0j53LAp2izIQ
3kYn0FRcCILPkjxOUTgaYP14EJMMt/yn7SlxeLom2O2egAC8lRdqlzBj//Byc/K1
tDW8JYMavx+f4PQ3Ld+QaEic302MOXz03aBuT6rxaeuMime9IjC2HnVjzdK+DjZt
ztvywriczhe09AsUMX9frsLNdz1DldVJ3LlNgLUPLAZetMPy+qSmnMkWwm+rheWq
/lJ1D8ebLaJncKoGdP0RToMKnBX5yHU0/xfQL0Mq6IgHqwBveO2VQjo4Y43lLQBv
c9+97FNta9SKzZ385boS/+ZCjgIoLe0q3rnHisiKmMJObg9qXctv+8dfw+vq50Uo
lRSUNp+S+dx+d3gB2+WNHL4wCOPJzl1tD30m97h9GG98s67dkS+6v2LRPDvbsrgh
ABAhdTDcj4XX1YBEV/lYJOwgD8x9dJP9x33V/z7FaaU46NAY6F/ORkBEnxQ/bZSf
9XOTQCpkVKU8r9am6pfzf9M8kkyc1gIL2VLYcmSUnIGnPXdDC/yLQ4RrGt/897pk
zmWrOyeCiTvLrfO8tOijwqugIUGhhW13rIaVAeU6ahotxx4iYjGd91WKvdPb2rbG
GvyHZLwdQO/BdhE6hqYq6GblvuJBmrKUWPs+QR/8kJMQPxMXdnmUxbFfvDFiz4Rx
8nUHC1Ek3bYP92e0UW3S+59RoYDYdS5mstsF7gvcZjGPMglw8w+crejtUiHeQ37B
UXYmB3VazemkqwKvuCp980k7MxTBvY+lfcgrXCm3rviiNzQGHyeJnAyOUFu6pF6S
eC0DLwaTQU3IdgV0303h5bYZ2lQZ4kqQH6trYpXBr7PiiTPuGVlWL/V5P6t4wkfp
TEV+xyuS4Z8WjgsHJEW8sMaBTppEf4WnYiilhspYn6OFqCZKz38/a9DU941Uuz51
0EiVDqtbysiCoslsDL1Qpd6tltQxfSRzo26MvebZA57qdJ5ZdlpHRUZCUeLUSbP+
hiaroJGgqipzrZhA9LVrD/lB/+n3Crm0yGV39AMyu0jXN2fV6vfOXJjDtesMaMyv
W4S9vpkWaASNAlwVNF1Y1aJIxVvQpnPoZGfNt8gWpdu6OmvkWywGrsj1sIPi98BO
Ptn8PSMksI6JUCjkuSz6PYImwmMmPLk/sD8zU96BOT/OaNCLYxxbcXrQTcexHBOU
FIwa6RGGAj5I1rSSPvHrJ6haUc5vKrOW//biYtqUVoqz47zxLNjD0pUAjQkIKsuT
FvdxfXRaBrILDm7qzan3YHFVyL78Ffmqrvzay4HJKkHF8hvwpO0F0jtSA6k4P94B
06uqe2Mpgkddq+2+JKHwPPaNwuW+GLU3SxCTttGF1ApFp1VfpjlB7nXNwYQDxAmJ
ANDlhc9r23bzz9JuMKPO0lWxyb91mXunD9wKTLfbXk0A7mWRw0RyXz9Oipn3pN6B
+Vq8ttw3Vt/BwiJ18/ruF99PfgoLCTb5Rl/JNEasqiR1C93jHB6d8RgGJBMYikd7
SgNJdxyOPj21dx+EwhADuksv2hewPjyTzIdRqzx+ief8liY2mscvJ57FblX3XoYs
d1f8vXLT2G7j1e5s0RupvDX/q4b8ABrnZrjVCOksEy+UusMwxY8Z10nK2n+B6sMF
TOpHTzLMaOC/1X7WY8QCkeweOOgy+gljRCjHNCe95kb3wNO2T3myK88M/fyfXjO1
AQMfJAxfQGHZVsldORe/gvSJM8qClqfE0EWnUiDlyUu/++AOwcrlhXOwMQiKfu1B
yi3BPctY0XRLoqvTTJZTGE0a3azwaB3qOJSIDXxHkfmSd//8Rmxin4dks3QiO/EW
4Zvsvgn1MkvzVJix1bNhz1henofpojXSXoSI3rR+8W63vNDE7Y430hZQEPga8G4E
OwwMb7u558/MteML9xvOhqT3l/lcHr8m5tszKwuo0rGfVsOlVAFC263+4Niuy1yq
NtHjfSUb1CZwD9MhHilFWvdpG4VqRdWXpkzz0K3qjANUfiGJH7S2gxrWD7TBUr8o
nQMcRYcwb87JH0aSDsKXiKSrtgTgiFj5nLSMWwMucfYvdgJl01axGVFaNT3CZJNv
Xoecjoza8TJ6Harh2oP/mORy7/nWXIbQl5WlEjtfJJ6Gyf/mHSYLdsGxXyKx9bR4
AqWGmxDrGtHkASBn9xifp5lEVw+F5aHk3MfMWJydjfGsyow5xIWsGmU93qsn4p6t
iehSzXcfgY6OCK2kW0ErmtRRmpvjvygLCi/s+T1YqaWq7d7xcplfjbnSlMmOOf+3
ONnJabYkxBv/Yp4ax8wkH18udolmwxUBPWpUewMjkMeqXf6MxPlm9NFixo6pmUY8
4VJ0fNAOCdYGk+dCpRPMD1U7+addsyS0H5gQo90uOD9F8nJwdzEsDu2zZVRXGIUl
pyPOyvuhlXcZILrssAvmG0y9P9tKbapFlNXIJ1Kdk7o0vnzyjcg3aDc0aLq2VGaK
4aYrVMOMNZtkAXHDu7lIIFRXLJMPdxLmF7BghFDY+A4RUnC01//vJXrvXBXDYMBv
+V+XRYM1sGsd1rHw3+EGUENJij0fi3yicpvoDgLu5H9QK/Tg3xx5a8UqSJADnyx0
oV9bqfiZPE4fsgCETiREhvZ77MvLbq6KXTRo+qChgQRG5xg9UOc8XQhfFTtJhRVd
b5pjv9wQzdGpSTVIeDJLnG/H6PkxkOubkyDj6cXPuxYE0zvfWgAtidBM9vbPO/yH
oSYNpIy1C7CCVwnNn9anW9pPqvPgP3+O45o8wdwTUcVHsyM6ovpFpoL1fvdUOup8
BBmthDiyHN+kDzGps9ZbsWzSOtzIjOjmsWsNquVB83G90/FJe5I2pOEFtB8hgOTE
i+NmV8EHGMhcIA6wDN1wSLF14cDl3rManKU4dgk7ypKaeI3wLY62NG9x5/z6wjNb
KvlMtFw/YFpFI2g9hbbb394vaRH5R1Qg9lrnmhm85JSK8dAp9o9J5OkPPjfnrlAX
HCMkVWdwF5i8ko9u+rAtt0fJ3ZyWWZ6zELIJP45g3vJAMfuNcpzw7QpGTLpobxdZ
zOaXOPvERWzENJgG8WQ3my3o2fgUKeD5B4M84i8oqrEQUdu6BcmlaJmqXvLkrUqn
sHbCHKjO/jlvnIBgsu4OLjeXESvtFlZBDpU/TgC5e4vM7ZEJQqzEBA/fTQsf5RgH
1HGqaqe7HEKCTo0lUCJwliHbEN7K7H681sudXUKzVvPB4TEaJImj80M8/08Qu4CN
vWyu/JE/jGTjkwXZ9I9wXpvIH2weGCNfj0Vw+UC5LIdl6a17pBxASjFSyL56TtaA
OI8x0twjeEXgFC7+p9E+ksFSvAf7Suk1yEQ0ORktm4nLiUkR3xJCP6aUwqyXbHTx
fE9A3ZGduVPRjBmUZ5/RA2KJaesu2Zm3QuJbDMk8dhzFo3rZtlHgmOcroTXOxNNY
iXFBeP9rJznGq4jTm5uT1Vd+moYzl7QCdDxQIXsfx6ttxt3yXPIc/aEgSHlEUDSE
0opW+G5owhqcTKP8mk5njnMijMHHBV8CvYi8/BY9Epir5QVGVVsAGDABwR/RQNlQ
3AUd6yCyM5UqaWeSXmBoV6F7WsxYWURnU+6D0ePqIu5y1pZQ90h61XYI0G0hcCcr
MEstR6B4SU6u8p+CGBBBTMNOaozZPgoOVpbG4UHArU56cJGPCNiunlMaZm+Vse8a
d8dQgO42mZT86k+QX72s8BKxPyMMUBgoG4tHCmkKdJc4aDVRwV0XAPkxSPKS4XoX
onbAmTuLpyL/4TYr7tB2yjyu0ATI1jZk5Oqc+NISNV4ggsZoVqDoQ7Y9XN0Gvv24
FAKG8Xl6lvML3myV/lIUDyuEy9M5VGgt3YwQYJtCesGj+XfHSiSwj/Nb9p5f/zHm
O0tukgoTZsVeywp+gae4gPkT1LrEFKlGVQQ4wPNyhkU07HzhPfSP06B71KFyAeqi
i33fIfzsoKAsueY6tzhbtUDAPJqGMBMss8+yM5Gsj4ZOewj5G6Y+B2xjpuRc6v5j
rOVDTzZgymek438pBrVkoxjSL+DoKNWyjubTELExW4mg51S/3IFTtjjtLq2YMzqi
v5Idp7rnu9JPaV+QM3aP3uEIcjm2N5TAyjs1dC583xVQpoMw5ZU+jti4j9cyJdoC
tfkopGuFPZ5ATL/9Vjz8GFoft2lcWEVlklYZ2xhOczz/ctcWZV+/1ouEKEir9aDm
8lzrIdZpMMDGxfxt/4iWyBcp4rtbG+Q5doXuGlmEkVAzMYlOhYSI3rwIzkEiKKKR
SfFrRDZ6CJ2j8tAe1ddhxJE+cAUvzarA3zX9gSU0dUSFO47yQ0yzVcLQqaV3sbpE
W2tzwPRRYyAbvXG31XdYrqv7pMFuddTMzKeWO//0wE7l7awh0GUeJr/Uczx/b+dG
3J6ehYfAO9DJHmRySK9FmL5lAJ4H0kyFxWQtfyv3cy50l4h0spaFfZr5r89DxoFM
0R+Y8KINFg2OaEyJj/89vOhkQOBME2GSuQN1ymkU8f3t1VoIboytvyCHVE3+NWsj
WRe7mWY2AFidpsEHFUmXLlv5aRvdRuo3stQa1A2vEZIwS8C0kriEbf3DVx5lnTX6
ZzzMA+x1qXGHPJ3UQKV5sbyFXPfvzeMD9LfICeMeJbCNZwZJlxeq1gpGkwhSj7di
vHpRyBXSekInqm3xDUWHgZDPo4KGWQVKe6PJhKADvYz/aKWuEX5Pu1F45fJuLHsY
jAlvdg4FjcJCVvY+rOvDy5uD4zoNco9gV5A1cl84vugjsmRAlSK1Po9slA5A3M7J
2p7z/HK6qRh1A/jWLjfaGuLjPrldmiednv9bsDE3zlL+xLFD/4Ka79jMnJ+6LahT
Q7F4Ay9kBOqnHU/J82+cldoGmfpAOku+EmGh5OifF8TfmCNQTCpqfSvz8QSLBs75
FEmIvtYPny0ZTICTz7hG9GdecBiFLexcVFCGWPgLXmyMv5EZuBlEnQSkVVp/yW/d
IjmYqPcwGuTZevBWz0DP2VwNuI1fIWpH6imBHVbcuZAFHuVaJgkKh9fgG9DAWrHA
TMWPqLijzooH0f5j4J4k6vQF9ZHJPwEvLJFpdXB6UcMPxTo5/4bh/kDcXiTEamtT
PO+5vAMX80k/fbeihXfCMY9d/8pf7iJz24BySqgZJVxHiEsvoaBidFc/B0agmI5l
4rxHqPs6jJVJo59Zl3P8NzwP2ZhS9nYz4z0v1ey2WGq7oV9WW1Kn1RiVsSyXsQZw
vTGXi55zt5Cg6X+syBGxa6wL7ELNdhobbHvzkNKrsDjad/aBzFSb0G0/p+c3HHNs
uDfPaxXyD5NZKvpSPr3imjEhn5i023xpOb7PW2ldbPoQ2s89luy+iUpCe+v6LLyu
rQRQW+OhweMkIsO8UB6EEEZKsnS7X0K9Yw5VS/8ifM8AYeG1+XVeSfuFvdHxPX62
78UBLW6a8U3qK4/4EWD4Ae1TDGiFV0afzUBcnno2XC9sheYWtGVsHwzRZtoJD0cY
8OcYOiq+qm3LSULYYbV3NKsuMQ9ySQ7/6Xdi+BdN1WhMXJjKbeyeO4XTfvmsGFho
y6pGup+XDdfvqrjjwZqtBWj8DJAAzWhnycJ2q4ztBT0HG+Wk4xecBlm87I6Jbwxo
OpFWs77racjkxTOVAg0tuMWdirbz/DcyN6z0+6W2zyfMX1kEgRdlBt9eiyzG9NZU
PTgPfKe732xXy5ZuiT0IR5ge2ObZd7t7y60l9rFWJ4yweqV7EZzudrB+IeTGRYSa
KImWtU4Ey6kkIRausFlCRkphbxyYjUsmLYxKjKxFCHJP6ngV37oVr+GwDiRZAN/0
pS3u/3bnut3Pv/hh46BzaZfIyfO3ikc1Jpj5ErPG+YJQ4It5XVglprnPHILZV5iX
6ZFh2WZ4hcG2Q6JYaM0xNhtdEe5vmQ8ydyi8wOE/zoOfWTs+Db726BIrqoD/BU4R
n3dsI284LqezlnRx92PWp/oioNnUZ+7rwMUD4gXTXwykQgjtfHwI4lzLR3OiV2BX
JaeqpB5KzjM6ljpLXCAbrRIy2dUxemKludkhzGkiD95OF8fMD4GYGJkTPZDVTdXX
d1+hHH1N0hXqI6LlpSOwn61ZRU4HOn98RXxRaCyg8LqinZRqbuSfzApsIKaKL5o3
zozK+Ij8s8Nyqswphcdjc2MIu7zfW0tgR98DjPIuzRY8MSZN1U+RqNaQx7EnWdCu
JzX2Veg8zlyZ6FQysOOT40BpYnIqEim06WY+ASa30Dkh3G9jwfu5IivxlM811ehw
BdkSz3MiBltIl95X2MPKWHTJ08ocpQ9SmC2nOmKwe7gDGGZstOF5ZNsxlfQPIqdw
Y35BTpdF7oskPFKZQU9RWKCX9rvNH4vPfSDpcRwFagjl0JxhoID1Db1QvpWg12II
AgXD4oCOZxsnFIojN1ND1DmpchvEiWF3xZqjxRCWReb73dinJd6dru1bKfAsWeL9
ViCoJz0Cqdgi4HJ49LTqMAY8pqNYsm0GBK+KPW+gcusqmMcNdDp8QC8aZFsnpjGr
eMK5dd0nshPLqEN0UqJa/XPazDPMmmGlVXdX83PAhIlKIndNJD5i4sn1xPrjw7NU
DZ9awkDyvltfVbdugEQpJh9EdHHHpLZQBBW6DhI7WcbyZR/tAAJOH+mlYCfbfjNQ
V/GbnGJa2kBUC045EHsugawLu03IX1rKWKP9aTjeGTGptd0X+MNWU86DE+kAGDDd
63SV2Zx5LzvA6qHb8NOwqxG8Rh/SRdqTxaFTzSrKMbYMYzXkZ31Fh/rNtZxlDllD
MTDbvr6ukSnO4nE/X4bx7m8qk7II/ya8j5KR72Lth+yd9gJ3VSyNjI3K9YV8J+Bq
LasvsgyG8HjDZSuxWeStDIu4HH4NY9gHBS7GpMcuA+75ozInutSr6fb6aN0RhRCr
yahVl2KeNCj43lg3b1KWP8yk5Y50X7aZlhi1zNPkOI0H66ehrcJsoqZkVBxSuSc0
DS3DaMFvbQJS+LflaP9d/JXvoeUIjQHX1poMbZSgzI0FEUpCPCq9o4Ppay2aQSWF
tsiN1gFRDS0n+XaNpuKZTotDHFtI4KWPwTeBbDelTuVB9RSKgk+lve5vayRRaFJY
APIq7yHg4EpCvjx22KzitxNF8OPer1Ys9WLD/NoKKWHgO55kjc9O7wQaCHC3DLDb
Oq4ILo17pHg0VyuKfteC7Y513vX2ozyRO6VAuHp7n/t72/G5aRq1tOhHKGF4eI+/
mqN9h+VVTNx5+AvP8A5x8sKPqCJTSfeHMTWLWPjxe2njb6TVi8c0wL8Ux9iGwW3l
UbetvJbZw5SRP8UflQ05gledJVIXKd0WukxmlaZiTAKm8Rye2Ho7iY/0Rd+1XQY/
2+KLSGXKzJv5iAkAxd20ULBT9KqxyVNfcQlsa6xaYhTERUph4hkP5wd4X82bauCu
uU9tuANe3XhCJ2mtqT5vk+arEqu9IElRoL27HTr+XRQx1zPLG9zv8tLirS0Jlasx
1guQ3+RJLo1OQIFTKhzKDaovDH6ZZw4zCODmw47rwPKTgC6uCUMasIVClCT+C3Ja
k656ye8I7TbHSH4vlg6ZZlmhWYTkau9mrNxRw9kQd4yECLmJREgo4vNrPF2gTatx
3WVKr//LXpCzzhO5Ff6PHb1SKrNZwOxeGRF7+MPa8hS/Ba+Ij7Xqk3k/yvsmF+4r
f0iIXY9skpa2B9ASVFSDIBvZATAq7RuMhn404aWn+uS7FvVbxL26SBxOURu0g+CF
NAU2Q7v18PvwgPq+HKG2yEQN3qxB/HnY5lQhzNWuj79qKz3eRL09EVmXXk5xk0xj
2OGA5Bx4lRe/4WdwGH8VEEzpKxSI/SXwSG3IyOK6ZrSaz9j5oRomJ+ZORlvbJqmH
QGsH2GEZ7mgXretR9p9hxhhHczOgJleaMRMfpQyK13R2pzAR8H7KQ9wRSgKLStKp
YuBWr91n701H0NWJSYAp4nfvxQx78OjGd4XC4wY/9f0m4ohCVk8qRKowVpAx4AuQ
H8yDs62+MY1d373NYbFeleeEKHm+MCTHUSOwXptrSAyQFL8FP/Fayo0heel7IFko
HC7/SktTTRrktCJa0fmgDHQW/5kbucu8sqv/0tfuFr2SealQAAJp8NWkNnDUrEXT
vbInRy4ipi203y+rTgKtkcE97ko3j2wEXjjzfxz5poS9PzgoWDcSDl0SkcUHx/cg
+PC6gKpfg4N6FI1Yp9x6+thmnbHQqaWe6Htgm2PIl+diO8TZgjIE1uA7G5g0FZ3N
+yctoM+eid04XQ6kFpqp0UBe/rBtyqIdPzZn14sVi5HRD8c6WqaB4fj04bNWVXgf
PPUEXehL/CrEYsheVAJY2G4/nWkFy6TfRm491Br8i01aUXnJdcyBOHEH2MmcGijX
AM2x5CqnbR40N/SVW5ER6FYlUmfoohWNlaKmPC5FAI2sjIXBb3kjz6TkBmw3+MOw
HdreoGGMvbNL0RlQ+l+5xiEGtcGt5/a/oswIaxP7p+Cu634bi2YukR4g1NfY/2BM
9L+DmBF7uA+oqzJ8CP1DCgWXhfKtup1RvpddPxEcmgbtxBIn98Xy4wCKteDdWBp9
GjS0myIu0jSzkoxN1yloJynqof1W9HuQK9AJbXJwBx3i9kGJ2XvW6lymToJzMJYU
qLvRmpu4kl6u9BJVMtCviMLqoKZn0WeT0UOrEgSEuSYcuEprrzsrZurdHQQs9xci
u01zNEMWoJMstrobr4IHxcYRmJEQimzLz1ykSRBfsZ/1cWsZZTGhDhvgCcOoyo20
H/VRnhgX61WGeTK1gt8ieoWrdk3fflgu1egGyIiLn2s78AZh0PRtXWvduMZmWt+J
5pVCr8eeEusn9LDiUTmlloxQj6PuleB0XBBI9SREHe6eHEW62OKyBVYVnnv/dk0G
ze6K91m520Fl8CaqWeEEZuy4G88VOlMhKvfPAVYzCXrOOozVeRG58UGFhzjF2bmI
hEUrFjwMBZ0lo8xV7Khu7u0z2oy2ZCSr6L5PBqVnGmvd9A6R9XCeyKqH4fwsn5kG
BHRIgnUbmFJvDOHvh4R/aDsE9+9iFFfIisyv4gIQ5+/JETnN1sUBiC7GfBNDFJQ0
TUVi4ZoNtOIpeaAIt7ZVbPRNyes4PJjm9wkZHILGJx36MbGkeU8zKpHKE0Jn4qAY
4sIPNOl8sBz5uZ2DYEvcl97ZQgERG2FMskNJhYPJYRmn6LS5M5mO3kMaT4Oe7iiW
KQzrebkCDzb7CR1dEuWYua6WXdDBpuM3NEiqnOAbJAPwdXOdz5I/wQVMNTuDH9yu
Hk6kvjmU2IkMOCBjKBf0ub9Z5aTj4G54eE+Ms9jQFWc11HeBag+z9HIg1kTbqfEB
EslNx+Y79x6fN/RzpnzTkdhG8yRlcdkLlyuaGw3iNCPBWZhvb1sJgZSRzelrB0Fh
uWiOc95WsveRKTi3uhYkal2BrkP+MGf/7rzeCinWjkopRPbhZZfXlOrNAf8WOvUN
QTRjuJLbjHY6A1d+BWVbooANDpaPyLudq1lK4uNt7npH8o3qeqStvXi9sf63jrng
ZcV3NvbSFmm07vRfGHNAJ30OT0C1fCr9qxOi795cKFEPqf3miaUB96zyrp4Pz6pM
s063+3L6XQ+gDpQe0mfGcLfk0+Snu59hnGzCijDpvDZ7+8j/YfYUQqSnQ1BkrmKk
slaalEKX7oXcdn3mH+fBPMnM32tTY06nH493xzbc+jylw8VKNgu3N/y7rRi/Nkbz
1ywH+6Lze0i5yrWEPLmV6JlMKwdk7E8JJgkzqqgH56aMdS7i43pxHgXC38Ig87h0
OkBJ5uvSrCwXTBf9yih8GlT6he30LueS+iri+Vyp92AsZt7goKoa4SoWnNvehXrZ
Ss4EF404kQ3GiDp0rn+RxfOMcYUbadIvT/WYnzptoQgSXiFEtfdnlpFBCkc0gwjb
SWU2eUQlEFctuEhcqVwmxe0Ra4BLkG/tzbffZHKBM4BWMF+GnWxiufu1I5VypR/F
PqOmQQGYTSD/MjlrV8ozYQDfD5kiiGFAKQ6bmGR9llrENR+NQuhvCRHnDRbgzPJR
cW7NXYaO8tAzRgEvUJ2ecZ+KRjPvZTlXajp+7wAWvVh/RNAjcJEIJCi8ctr8MU49
V4uMfGk5uTmK9MSY3ru0EpzBI6uM9fFpkSrtroDxPFCEN1qGNwnUgsi7ZUY2rbnk
5kEz942X6ZahnzFlA9fUEYdy43OzPlrZu7bVjsUH8zFMqzOPDuVCl/c++FRk2kJw
amE7QwELwDJf/azHxhXTeXfOi7JKDSidxQMxzLlxkcDkWNtw0W8BF29lNZnHzTaj
8TnyD7hQA6moJLI3hTSfyi4VI0AEYsGwgMn+putRXZ4ja4exylhYEIAdxR7AXHrB
GvALtGpjm9CI/rLGZdqmHRpU8ipBr4BCeqSCOPv/5+zD35ZpnXFIpFsEfPkkuuSS
0blAlAcIKnbZjLK2/K8+Tx4f7w4w268GQlOSuBh5arNfXzAiXLeywPqi53vxKPR8
vTG5QO0BTamkWiuAfsbOMyrgjiNN/vxeCIDjMUXNtKiSRQSaRUNwA49ETKn9CfyR
xeY1S2WFxIOEeHjAruUkqJSXjrsvpgMCmXkYrzpm8dIe+2ulk8/sA9FXnTxRZ3o0
oI7cTHR3QCqIYTrYaqJdxFYlKJ+2N4FF5uumbkSZWw51T6rr6pvBFssDQ+9WzKF6
3tCVCKvwS3ub9lNHI/JRmmkJLnPeQfq1tAX9Ik7O3F8ihkbJqQiQmFZH1GZ6OVNN
xOAEG5vVe23r30lLPw3ojy0/NM1aeWJSkb/KAi5CxTDvyw7jBS4dt84zZRM+WNV6
o6aJ1tdjrh6CC21vX9opo39ztuiUS3bslmjugysprTrC5N6gJYCIVL5hwC+2Ynu4
osnOl6ZuLK1cwLUx/kJXCqcG7wT1ujs5W+SAgqj069vYqIdzxlqZRcK8kuPNO1NC
SvCaVRW0KP8+6ZjzzqT8sl7zrM0oLS6R89R7HhMPso5Jy5cEHQM3yymdGh8TmY1y
BDfftLtqamJyqaXz1szWFdO9Kr9P8WLEnE/FhGosYWBwxcTbUbrVd8XVbGA7sM5I
QwcXKo3CVQSnDPwgz3PBwn5PY/0mpoUfXP4LwM4yEcTLCqzOT5NzNentFT0DeitA
h9qbEtEhOXLAkLOBqfr3xO/7eOKHbyQBuGDLptuSjyYf1+BmrwBCyGOrDNVIfztZ
6k6rdgY8HzQYO3bzGT0tbNL1i6OK+zuUlqV/c/VCbbUhE7u9gHrN5Rqc6HM4R7Zx
ET7sbQCGrzvpVpGdaDgFbZsoBDp0IUqB5verYiSLhEvRnFKQ7Ga9gMvrXPALtrFi
yegSMLw2NWGbw4TT4LiWqfSLPFtJ+5lWPDSzu3FoZ+0G/Q38+sTFPHm5l5UtXuVn
9m3U2mzo5SyWOYffCKA8K+2YB6rqgsOK47SmEkbhOhkLu2b3xymK4NP5hmift3bg
AOfUeQmPjto7QIqI1ixMcrzP+ksXj2bm1Sgwr+nAxMy9bWPGIvgNCPsB8JOw0H0C
1j7TnvUwYEz1rUxVk5HaQvVEjgOAE4H8LDu8QTERXf/LRyRY9LX0tFHnLModSpHf
sdN94mnEgi7/12Aep5qjF8zp1Tb/x4DGvarU0OpJhXx3STCjAsXSIC8+tjiHvUPd
j6ELDz8SGun1GpJ9NYlSjP0yTJ1zayJhJ+/0Ba1UcZUFDaCr1BX3EvJrkd6F47lu
gnpFMxLnp/wkBprQS/xpFtdVyPvC6I9Yi41To/JUtuHXF7HWemY1JyLid/xQEAyJ
37cjn0/RrBBMFdQTEPXX61Md1E4SqBlHkElIacSqtC15+4p0v9En6ajJiR6Mv1Db
UM1QCX7/YsJLTB1a5UgihZequR7xyVRs2jUjgZF5PwrzUCsF9FYeCMmmXaIxkY5w
j4YwM3KbbXyGz3wCC351VKeS6ZqSeNDAXW/Ase7yaxI+SKWfpHIHJ2Sjpiinlsur
ooDwMMo22zK0AbPX9xiSEzV/Bq8IPkr8maRQUSEwxifimv1gCYlXVrWjvLmr5Hle
LjmQ7zGdJ58tJ0AFYPnKnOf1hNUQaDJvNkPFPjDfBGO0w0OFQuJ/d8tmEN/Nj++l
hx9Gi00I3lw6+guz6U1tFVQ340oWae9Gk1ywCQRZ+fGhiALtQ0j6TXPDXI7YUWCk
qnWft/JJuRTLyMPhMhYwRFL1YLbCJRd6hI+HXVTak2V8vooQlno2n/LeryS09kLW
My9G10lHKw2dy9M7pVu/wZKFTnBA/+zZlJrcNhExKBHhZjaGbdmuiX4TeODjhOOj
hMhRpGcCDb91Bmf/N+lG9aEa4+iPLIQafJLGWK8VI2E1ogzn8h8ZqUtTIW8mYap7
CGYF/xZXCMe5crIB2YYtS7KIR2JeOPyfnQ0xj6Vlwm9pGKLuEYXip+gTgbao6Mba
VjLjdRW0PIqOLLNgvmqptXE/OIKOCoT1finOzjxbO5Jq4gVTNVqmdR4QARoRwUMd
ilcy4Vl4aHaXN97/CenYP+K3TuZTMx0gJJ7u4pe0Te5bL8bO1mNPJ7KcAgJUwsKS
J3iFze9E6rB9AEUqZuNmm2THyTlhxWsd96cs3Qoin7q0uw2kcpQd15PdYXhhNI9Z
iFPKI+2XD36K9iNTRQxLBJi0t2dUApc3WHOcN3T+hcumuX1KBpGz2us3u8uR5n10
lvJouNQkn2Gchi6tIxwaOBIMz1Hh2S2Nco77jYAKK9U8eJ21Fnoe15EU0KZwnoWE
6R3+7wooPvjo8F5NngzPKorASzXlP9Isckt/IouhEInFdWuGTQA2TS9ab2CAlijH
u2OMfEOX+s2jikI7ffdgc7NjqfmYZPNFzr+UTjy2+1eAM+iYkubMGGZrHfmt1tcv
iuKlF3iLkXO+Llbf+fngtt6JDylaVHzA39zA6bxuuDec7WcnCqBHBRrjHQb+umcH
E1+R5yxJtqbTiBcwgBLObCHWI4H4Ny0qYRTgJgR44usz6xf0oDlXgCc20NPMWH+u
+6grobC3RqRKQVT87bSNEzHj3Yuwe70sRQO4YjVlJg0dAA4Wn9IscqaZUwrBJLnj
df1n2C0u4uyn9Dgr1yQAT45/crsGlRqMZ7pBVJYKTnR2UUjP7eZ5nGBfoK1+RZtn
oD0n1uyCMiDUQ5oa1wBQ3Ws7Trk4cjY+lUkE+3bnHvwsPFH3r/QRlfYVTCyAf/Te
sUVSh6+I/tMTmPiAvgj1PEK+VWzaXJUL1sYBaj2hyn90PZ9Q0uGXdyRDVa3EqtCR
WvPFWAkViITPkGYX63DdCy4+wMr5jKQid8GmepN1dwQPbDnLbj3clDjb00IyqSE4
AiinVajddHIEQLiOXKskqlWk26+/kRGRE5qgR50euL97+nJS2eTL/sh2nGTfkJWf
AdafVzLAK3HRY8nLAL3JO8Pk1c+Hgq068KIDLNgjMfHPB2XiTo+N7CSoWuyLNd0C
lC7W+B8cUun3Re8RPy+xZJKgvIMelcW3c4qDVHwLM6SHXB9KhUleGJgKyNBWQ6T/
0XaA7wC+JoQylJ2UtNkX3vKLhJZtp4Ln1xX24rZPrR4La1DkUf2IOGRs4Jf6C6md
7h6FiG32gj4RsRBVNLmtJ3cUkvOGbYJJxGMBGcmVhWNRgK8TQTDtRDavHnAHKTI5
62DbQZr8nNaWsdztB5FAk1AbD9eo0suLhW6ZcADgdinf5pY0iPatRz6BJAN+zJKA
w1GlPZo4q2Mw/stOHb2n5pxLUxemruf0SF//rITY15aJlJ87d4csgY2VpFfuBA+p
7XMnb3XPn1YpHI43LDfCq7Dra3K9Qn53H/fIrCFrcg8zUCSaUgL38+9EM2LBWiwE
JrIvXE2iUED59ajX7hXP0UXeezxZqy0OYgIv5tn3rKQRRPfIAD9XAY6vsWWfdyXb
PD7Wvxgf24w4ioSRkfHM+zbFVBWvY/flpGjsqsnIkmPOhuT2XGGyxV8nkMn5k9H1
0XQGp4Jkg6o6ldrSlDM3RXdyu8457CKc3fDZh+eIsmAz0o3k9NnrWvaI14tJPJDo
eYP6gAW1etI0p6wDcBOE77bEQTFXN4H9emAaZyp06PcXK0NbGgJ7oBbBQLXT4e8D
eL50cLaYIB6UcHfka+o07ksWJDye+6zBzZEUkloiB6HK3GycQE69XiI9isuBijkd
dBCFmVat5W39N8YPaczVZiF+3ygzUnW4g6WTTfWX1puKrEuNAzVcZYZKbJnIuukv
UB1M56sWY26D6TPG2KtQHPWkt+kPM0gKoPjZ3AWsja2+xbMn7NlqH0ARfH+9NzSa
1ieWOHQAbqaeq6La4oNYCKRvSS63Oms+N40prg19FgidCVw0HISVuVNOBubSaUH+
UFUriMmA/Zg+0FaJ1ckW4/034YFXc1/6vcZvy5ZM6ByNAbCnviIqR+Yx9zcLxXzE
AHjyEnai9gndia1gK69uF/tmIb/Dctqe/sViDFFjYAW2MPPzkNX5dwPaoX7+dTqG
a7pMlZdkxS+kdqOvw2brV9+j0djso4fJ78MAbhFdbsbjXgHJWhcYOi7ddsFj75tj
u2LaJUSkEIIDPAEOX3rhfrakYBfXm+yIIAFh/NqnuREB2xQKpvsHbd0/CGdUr0nk
foYlQatoMtIEznUzbEeW1XoblA9kQ6dYAxTRjP5LcRls560WOf017UmMYQzBDc+G
ElJFHMqq1hTKG/jt7pjE8WP18LtPSMtok0uUo1dD1RxtJ/UyS7q7ZjxVgApRE2Q/
OspVY+c2SHxDUJxKeKmhz3uC9xUr5wnh8TslK+/zcZc9O9qMhzt+upqzp4EEBQ0E
FPv0BHzgxrUaoWUpkNkf7NxOK/YGLPWi5kboXrGtTlkP8lh/uWvgBam7IqgajAKH
uDzkTXFiG8F0MPFVs4NjcHVZQX0C4G5RumecGqGTDd7Jn+PusKej67ykheHJnBGd
TSI3wZ17XBK7PWYFInrGrM6ienxhGWRATy56sdyO9bH9JjoxajL9WtVWwQGuU5dz
qtJFUxneH7Mg9oOpRWaeka+9kM7iEYbdFsvWObe712BqrlzcL/zok95Y20NKhOtv
vb3T5nYfqaiYyTKH4Lxnb/ZpVIo+Vf8/Y7GH5IFDLWYMg2Q/XI2EG8iU/HLZ6Euo
t+VxYXKsQOP/usfrhhp/IFxXOH9bLjkWMXZPS42MB7MWMyxCViHflCcAupHlvbWC
xeb0J20EWWhDHVHN1ZZlq8usn/s8ycu+bugDXVwuUbmyUuDgyrSDGLNwpzMC5xlV
vr/aVZNJz//oJzd0CLTpSE8bRKXi3B7e44mYjKrmofHv5T52bJhYwIfvsO6lfZoJ
6Eb6uSmzE/ZgsCD/sHVn+GQqLl0I4q/F+JYdmKAzJrOfstb7BI/W/3YcTHuxxZfR
2NHj9ItaEnEqjCN3rEFZBPCe/g2xG6wopdFporDtD+yf4PAnguTFQ4gARdrkEcVr
xmIhboKEg8JHhZ4/77cp7j5Cunm2jxqNvIgZivpYFvx69q4r84pZREH5yfdcvgig
VHwpmELpF44M1F+YftKaBnFzqxogulZF5McanyYQ0/vGqdiT2BeSCf3UFh/RKo9C
wqiCTz3DDzYFWMdKb1PAUINKxM6hp1zJSh2xR8VNdKAw5ZXimUDgZZdCIjQl/lZt
MJyC4KQ5GpTHVDnX/Fw4CZ2xldUZCB8aM71PzCcabIJyass/4MaRfZXjyeXTpaDb
f3c40S2wv3yOLxieuSPl/tm0PMTJGIU5Lt8qR9F2MOLbFlfO5Io5jZw08qM2BNH5
Vo/q2ExKyp3NZm+glC4g2y9eC7h1VQ1+7F/GDZhCILxMXZ7Xr4ko67aA9A1Mcj0P
kwKxMKZGQO7Q+bKLt8SQBjGVCzMl6U1S4EWpkXozOYIjrIEKl/OqCX9x4QqwJeOs
iDpY70c7nWweafcFdRL7onpt1YrylkQcU02W0gUTU9s7eqi4HJLVNXF8egrYYdgj
RmVVILFpUj8dLQakPghkJuebzyBnEwl2dQDN2PiNB1bG0/YhRj2jw1/vR1k0c9UX
XnV7tZjB4T3GDvRRQDPSdESHaxfUzlWESTeIzghDjtQmtR1IRAKKy08SibBnYsFW
2j+CmTpmAWid1krT3MRwofjd0ZUZpSibmyfTupzCPQtuhCAPDYz8zyIstnIL+01V
hH83LgjTbbVBXVYGOUrnjmzZTrW/OKCNpwTIPi/wb4/gpgSHi0jC6UN6Ur80IdEz
vJgMeKaRCOJ6eLZNhn/uD4TR+FZrJGD/q9Y0DINplhSTGT4aXcRK3Z7u0Lqzykix
+2XBTSDXHktcx+q+gMXB/mURyjcsECia4YxQ7ZI2yYtLaGMZZpwbq79WAXLLKRTz
I6RJnr+TrqbiaU+CdULrZzN37SGpsaGchER2ONl+LGJO+mDNluIu3gWxWKfQwLO/
laevx3bgG870WDJPiMTPo3DWUeOMQcRB9q5QulDuoCKp4w5Huy6iMqYyGw4oeJmZ
lv/Xn0bQv+7LkjUNlAgV/s5iGYDrRxwxsbXiUATnmQ9qXJHueC+kWz2CvL3C9K4D
PWK0dvH1eStYJxWa+VLtuDkLfxOC8UwHDsFSeqXeV2nXkkK//g4vTseDrQd3Tp88
15xN2SK6XhumGO3OhVB9AuSiw+Vuq6+roWg7jvvLB4k+9bfYDJympAhvFtdh9TNa
dqw5ne/j2XGd+7BAe5FTQQFBW77n0cHgrkPymFDUfQWceLilTt3uKvBCG/b9SqcG
uFpJFB0mKio34CrqFHMjQ0BzCyMMlqdvFApkV/bOkCVvJMhAZyZ3p+Pqc+rSMLYV
Cjb664pkeHkWzDQ4K3eE6xqNr7QX9ViSwknZrgz3asTqU4tgC043XyWUuj9tH0nr
yjH5sLwAoDNzWWQRo9Vtb+ykstuQ0B6RRArOD3NwvRzR0RvEswhWaDX6i/hSQTv6
ekmQvOG5XE6NksqBDHVQUNdv+UkwNQuMDBLXWqIOJruI6vW/U1s1dtnr93uZSRQX
Td7HNOGIwuh7j8HSd2+m78evNP8LdIsXePnrWAc41GyIm/YEnBGaNFRqCuEcj2tv
5j3jb7edeuD8xW/fnuULssVA4yaAX2m5+WqFkUda2LGQHrLAvlv5iJAplcA3QnUs
fVW5AXTIpGC4ws1bbVnD99Bbr08q0xtdFxY3pWcCs+fzcFPibV2yYH21Ognh4cQK
yLQARy4lK9st6SoqFiPFfEb4VRKPPBwrVwFCmIecnvc+OJKxIW6C/2j5LIylBy4q
p+zcxuh+SbzElCTbDrDqT4IWFwHd4PbRE2FUxu03n8leqtDkjH0lItRmpHUZwSh5
eOkKPImlHNaTpM4M9Jfh5Hn9nWs+grnCH9LS8lwbpnkaAZjIqfrlVN48vXuitePm
3vxy4xLVCdSheJN+jTQ128h651R4Dau8UwynPPHPpI3uDyiQ9sVezbYWlcstRfXO
meSbr/pnT1hTHVLrGEJukfh9LB4D6YMekBBCYCivYsFTFgE3aWwgbgOyyMcNee6b
Z+vfmp4ymV98y87GdhMDqr8vScPqZqDAy2B5cbBJrDaa8+oQ1B5pQWmQ3cZjAgTx
0V2U4GK4i1ToVdaBbfliy2OloHZIicc7D79KnO8SXIYavh+OnjUPYsTEgEX0r033
bxcACBTcrLF6fM/yPJzvubLLqIy28FAPlDnJQ/BKm9OpnSl8a4n3dscowJ1kZJhe
jqUIzFm73WrtANDPIJ/RwDBlh7PAyOiIjetIWmNsChrLyHbTqn9OwJND2StNve57
QN4SZjL3ooOglNwUMxLALEsV07LnExKm+wiALxzZdA/b0EUsZn1NpTNAlIGQu77Y
0C0iGAZYPqLIyvfUYQAmYajKpATwWPdvBFIdQb8+e/YYg8FEF0pis6bBUDYyU1kG
Jnb1i8uQzELUj0t6ptdio7OtQtVZSmDTurGPxhj1KtHmNwqMwNzMaxRjrc3dFmQk
OoMEwySWYuzbsra0PnMjCSH8ArA+cDkeAFExY5xyv6JTtyRJnIqN+bOn+L620cFU
9rofE94wnKqKUPT5kAriL7u8E4LMs3sLDbTOH4AQtx5WjzAZdDfntQ+Oj6jX9YIH
zKJu7lA/AXb9jYJlOrjDDOZSKRq6Ucum3RGiPqzz4SWkUndD9domvOR2CzchSWMM
rto9bfnfTcwl6Bb9GJMt9A9ddH3GoMsoSMqa5V1NWPaqnlzfzX66pspcesVK+RgQ
blO3OB8B9X3n9uYUjfm9tJ3D2T+9cHuYh49rWxbaDHOpHj+lulgKc3uyMTFgfg/3
ghTsQ2t954ppydiW+S8XYXwfVXav2IsCs+3DSVSwe3Wr+g6rKdRryUbShCx8iizK
DfG4U8kxqNM7j1PnYhL9e0BEIQn6UU5VjFsZcnDSCxVc/2gDGLiUHUAom0Ub8Me4
2mjGtQlCnQDFVAGbaAkl2E61Qc9d+YIZJcwUJyYcGjj1A/uWNm5ZPJjpD8/PUPHZ
Gm2Gms7fR+pGsTRD0GQpqWbp57ZRRXskA/8NZzJJBQozj1xvlUlCb8eJsVt2orzv
/+AEv+BLdTWDspqINsbtUrnJuQlt7KE5Oi3zLouY9n66eaDmymLrFxCYsRItOE9G
nWUN2VhzmN1lNI/gMPtw/HxaR5Lmb+ls4VlgbZMVINi7MXegqy85L/aqgW6UY93S
1I6vWL0C+3Eb4Ln0cd552tFjq+gKPqeJiByQSBvq1Er0wuQ20vb2MMtm/QESAOYa
jVVPo8OFdWkMo47C41cKKHP61o0xJ1nzKh/2IIH5APRvrTMHa200TWzQAWXmCV6h
16YBmcgsEw5yVkhfZWp4SKBN6KHDyjkkNh+Cy5jqjDo6uHbZlKzAVvcjeFuxdLIF
tkfXezzDZvuRIhp/Z8n4lcS6HMbwuDXJqBKUZVBaFahQvJ2nKafq7n57qiPCu8qA
kFJcx/nvZJEtdWjFqxx2YrQAKaF8XMbLs2T9a4jBqCHlRs4fIBuwPJjVzpLdfUtU
YF7x9Lr77q2VV9WNhaFj3ZIQk0lyiu5dDhZ0riSb6jYOGpBlBp1Sz5asPtlol1Tx
Bd4w2+keqE0xSxrb6ikcFn4Nzdqldn7TJIqPtsV9SvTDrppvs365eqnLloxs14hb
Qu4vhjBLRe8iiVS7Y328efiz1t5tuhBxLMrqBU7A1/Eeo3fnxxZ9fcntLFWtDdTg
pUdvc16TuEDQsm9H/TdMR5ynCdDDqsYpIq+Kvbta4PXLYMRykrRipXNrScL0Ork1
k17aktaqzOWE1Qz5BiZ4Y1khkr5l+yYPaak5/6+v6LXc8zrN+NmjIZjtMmL/koNx
WbDtysMddkPA1AIYeu8w3JRZiMA+iuPQ9u9IWQRhCM7AZ/FIpx4DjfVjAlUciJcI
`protect END_PROTECTED
