`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NiqgRAALeL1epfnYH0h/UXH0ZYAZuA+obB08zBOW01FXiqJvT0trmyjmGJydaeb5
LZcc7tHA+lcdJ7pgVco3aY8Q/7P9vTn468q4lBd2kD0kZILXU61kwiDIHvWPfCTb
IObX/Yz23vhb2EXKdNEEI6y25abUj9TiFQmAaqQCXuTddMmFnOEaeLdi/JM3BlLV
nPmWKPU0QaQLHDK3+7d9aMidbWuhZw5f+ecs7s6vVIvGnE4LV4F/m8YiZNx3XEx2
OzH7iNAKFKzBQH+PWMkmP4LEDldbzjSUnlVZ1TY+HxRuZZZ5v4fBM8tmYP+FZH3c
20iUVKQyvbAErth5m9mCFtC2DJfwpAav8wOkSUjBD8ZhW4yk/3+Ct4/ceQLQtt6u
JBEBlZ/31r4LYNc49aDF818M1v8LfiF86IcsirncGJMrF0ax2/X7wMe5lg/p7PH/
So43Dym8BHHK47CE7AezyCSSSTQlNBTsa9640VcqyHI7n1kFYx/yoY4LR6whZ0AS
nGfDQ2tuGzoppgx8tiGjad9a5CEnd1HjJT26dcUbaqNjoj9vM5Y6+J8amV+D0LeI
5J8Gsow7fjpsA5jt/rMucp0VxM+qgvg3SNiW89uYjWrflPGVl2adnup3X87KI1ne
BsMyMfUwMUNTz+CIdOx7tKNgyX8hqBmGrAtzlaDGmRZGFdUxmC/13g1dvaR7xgbk
35zac1yjOoAbORPqYdoM2ifOM/jvA2qkM8rDhOuisyetf7t471Nf/P0WWPtRrwrx
rdbEgCZBxx9S5AndL6XMgfht0XKI/RRV9AJu1+PJkCrSuwYFIteaI0Cjw4PcZqhs
k4fvapDmu6c4uN4WnoW9WsGatUAWZythRb+nplq8W+rfr2CnIXhMRbNhIYeT3P5c
eUmREcTa5PMPNwXTeu70jSlecyuYYGa3MbcBoYSeMv5svtNlqCeT24Y5ri4/l6zB
McvMTV38P6gVzgipSB35l1nlmKWFSjoOyo3CX+/xEmfU9H3iKpZaIJmoLGVxbG/Q
s6HAWhDJs/0Q5CtuSlk3w4OnfriOY1FaPlV1L9MLu/a4Qji0rq4B4EsEHHi3ZSeb
vS2zmoK9CyiZM0VLrTb+bybkGvIwAxcaAy0vmao7sHy+vWQ3goVyJEAvPvwedzYG
v3HV4dxnd6YYVKbLG8g2SBV6WWvRO07H7wXfDrexV1VWc7iTJXcKaNqyDf6gHn2X
Z9iFqKFrb4Jr54O4K2hU/MAL5ZiAQMfOSD1f9PIY3YyoGOOMPhPAaPk4vdOh7AOu
7GwbsJ/deTnEANhWtiVuX8XiSARUD61qGpDC5639KuECnm3uxA0+8uCDBxlcS/aq
XDiOb/W55JBRWHsJpJFFkw6hge0vEZP43NAoLcf2bEok4QblViusku667uTxupbC
cAlJo8RqAyn4E5Fs9gqOyQr0KDg5eQ+EoGlOB1mT+AlFykoWnT3QjhQSY38jAE3C
Z8TKcC8YdLBQkomSvx3uGPzJNf9IkhmspvmIwDfOuKiudmhrgR/ILZMjEgTLG2Fj
so4Db9uSuHmTZU8fwDUyMMliqQBSmOIsdfHUTqId8S4+tsBC3LkCq4cgntb6Nm9D
10yeulrnkgzDwGe47CuXJqu5THVtesw4T/HDyRRGBK9dbI27Zj3HJ/voS+RPDd2m
VMAGjKChQ48cttAnUTMdhXrbfYYZAITv1YQg/e5lzbpZ6M5RIqmnZ/xCQQf3+pxW
M5X89beEhHxFZgUQsdiwG27+hCx2j69L42cibDmYf8AOmmvc8yvvfi6AZH2tA18j
Sd0x3/KjYPH4Z9y6FsKbOdVNWFLEbSscfejIkCDlGkCFhaUGtcwT7iovgX6LOG38
L+TnJQGJ4Jd4AP/+gug7KhT7YFYiJcZxYTGwdOq/qbTkLvr5p7NllqwD83RcY1/J
osvxX0f+aj57nAwnRaBqSGgAH05UGMBy2HAMUtWb7K17hoRTLQywj8vVIFfIDsBb
aHSFsE9N7cnTNFxs9CAYZogKzHflJjdrJIlp84FnpJNestDscJ66+xsXXAg3/I77
at+ZcRbafiyiTzbtBAeBZXYWV1T0rHIWpC8AlujG9mFfdeu0O6M22VPXYuPmNaoS
lgH2VONcfh4xY/7pIJ9GvAi8SiwhNBlBspjK0ArSGXnSgSTQeOioPARGf3bqbcEK
dIYrwi80XaI7MEteXtkpUsh5zErhQtCXzcc52iKZ7wR8SE3rENmZEkApd+UyAUU9
qzziYiyD2vCuFrwBo7VC6VAQxEGejOIB7F4R6Gl4KOXVzb4DiKary4YM581JTxqg
qTyozLs8kxBb4NPEZkx/Qn7sOn1nYasekjCZwDfMIVD7NN2OgS5EfwYYbz28VlPX
566XIK54qT4VSvDNccaLPraNDwTkxumSG+RxaZKkj0tzVy/fRy1K2YdGA9o7YIlV
NYj5vPnmZU3yaRs9FFntpTRIYxZ1HOFRfB/s4jsTRdeOp62n/gI0UhsufMfP81Sr
VSRiHClOeG8RUyPZ3hCy9QcmG4aP/Ty0hl0KmBPVdpTe7im37GGxgUqBYJUVlUuD
XvKNi9mg14IOeu9igaLy6GK14QYnSa825dbJrUKb4QZr6QLHMILDnHIbY/SHU3Re
xxbsu4ajDwf/laSmJsvgSnHCLRAZ5A8b8ukW0IAquvioDtFspCaW2QGhMNlEu1sk
i6rrQWwHm1O9HkQIHN6HOF12Blx2uKaDfuShSiCb6LnTsEld7/Wc3EfucWEpqPhT
aLQlRBL6YtlTvhXkanrkMbJN9yk8ieuSjE+8BydD8WJz1O4iITruxHJcUBud8464
r4FWx4Si/9v/TB6EDCDQNnhFRmplVKx6kFT8Av0AdUqoG00hgS+cIwlQMN11+HIY
BBYCBQ+KDX/kZI9Qg4b76G80a0y7TEoBfvqEfO6Zd7GPAFSC5TIEJVSCl2eD+yt4
FrfcMqOJrS4CD8yEVGS7muveQhqNZVaSL4ZxWJY6fsxjy0oeeA9bYG+s06P4NY98
hw02ReGvvFW6c4UWiCTH93WRM3fRM7d8JYLWFHwPvDtBzGwx6oEaog828vdnVWy3
+1jSIEDJjclgSD72tG7FeLawthvqxvX99QetPQscgDjehekH0zlc8pB92kXk48Uc
xCmlrnh8a4lJzt23ppVaezBJ6uJfsX7zkav125F4zci2KXM2LHzAZYKS1W4hW9V5
FkRGtCkP3h+5sG9rU2V8lrndmh4isqbqxnWKsvGGiJ0RC4S0QUjnt92uFn01ADG7
Ve9sRNg5/+kYtmj0/IUrQ3Nl5XtcLcGM43LVIYGxmTa5pb29GoalYaUBgxXoc+dx
Bo/8P45p+dIeIzuDgKfdpnwNSY5FIsXFDb0rXJ9VhueP2LB+hRTckHB+8d/qYaVy
/wZLH4xY1ixRcWQ+8d4gOaoVbjyvNttPkqP8UYD5bKaCe2azfDuHjgaaULwvI3Il
HUYQbbDkx1apRbc0M/Gke9Y87uG/yqUcZee4xIrH+fKcHb9du2Gzbobc8QEi5+9r
PoX/N48kRmfHzRbsBPWtbZKt04EplOF5ryko/G4+tOOkFs3YTJgviciroBdf2DjP
WWqNrgMDQ5XpjED41DgTER1sT+9OKkUTm6OAXCYzpY/sQ9HXYxc1zsCVOkG/Ftcu
LYnM9hfKDvlezItvQwZOE9I8q7Rp6uVtDmg9I5Aa87rEKj555Op4JdpU+hTEZPCF
k1pNCoZPJpglijBeJNdcK28TZzoSL/aRBrb9Z/o26S1U5bjUz+JUkcQxiqpP9CjF
dgqS7vxaGg21IgGlKuS2hGqO2JgvqdVGSNG/PONw3MWBEnzQ9Eh62U45B7fuNkAX
xia+ShIEvwc9UaY7AzNlVGgQHz+J/acLSg1bzMnVvwlajKJMa/05ahamEKSossyC
FnakQV7FQYygqmOyo+DKovyqfaH5g29zu2Cb3YBvJwwUbcDdlIiwXE9VLYAcHX3u
jihJL4dfYVKvq11RhyPbvY+0P8churbBkBqJTwo3MLXRdwFe/JLRH2wTImFmRfHx
/aAy+87WWDl9ja6vbBPDRUDc8/odE7ep0B+Hid5AtQaImRbWS06ABVtV3CM4TkuC
Se/NUhidqMdBbTd32nSjwLowAHYjMc8tO8iWzJZ+eXLJcYvgC76wFWojgG1oV2D/
gdGEJvPExX0AtudwbHXXaz1zJi3iaMz4rtoKBr5KKg7OE06DY5rTc+wUCR8RNWXO
QaQ634irw3qs3Fe1ffKCjcoo6gyR9L8rzmbDXls0DEX40pvrscZO+E5d+QOsnaE/
/pL34GyQQBGnPoPkWTMCsdcoH1JHJtassqjXWcB4+C38fwPCbUkcX3m/jKk224fY
SZWWCBgMomJ7SkbB5h34I+X7TYLlOoz9Ds2h94TD7m/I712P2fCrn1BGXwvSEqSU
dsJHGIEYV5D2HhKVcSOtkrzSI9qKr4XKY4imb4pRvKDOVVYkGsKXfWEX/yo6mE5R
togD+RINSA6EeUPVB+XKsxO6qptuhVl/mi4MoaDMWX5Se6JoUe4BRDZo7zgysWCz
ChBm4kwjEWKBQowGRxDJACoDYcVYVJbuduP+3A8ojgd1XUlXdVfkhri52hUIeOHG
GFzZepOAVF0ASfLHdCR30cI82G7Z8343cgNRzQriZLdls3Jyw6nYgQXDCLCKkAyD
TF2AZz7YXEHPJ5oa6AiaIbxBy2tikBjdgYDYcT0ELigyOpPZqH49JjfubQOvQUFI
HtxTtJbPRpSOtky5HDHPBEIc5d3KFjTpPzBqMHuV1O+2z/1UTFOI1nD5Y/NwfeFP
Ve0YOivnOkS/e6ZRJE+AV5kMpI1n7o9/QvDGrMwcj0lf9533JuryNULcNT8Z5pRz
poar8n+49beabYr5xthDFYOmfIJBZieBaWvlmfw9M65ce9mXpuXWRfyE1QHaShSg
si6tAAks2O76QdnabgVnz48oSmbjQX326hwn4sc3hFktq0m0AofZRVzdSyjXrWhX
PPaWDbpPuwEDSPBbBWw9Wy1v0O/Y/WTIPdmztgvR/B/27uzoq6wdSEY4GhtVlTvV
SBSoA46S1ZzJ8MkFl1St0Ad5w+/8wj/sfMpyNSRAcYGbm15jjEok0XkJcSqCqATW
ItWIzJeP0FFKVFGuOqMamlXK83BY7ldO8T9OFrds1A2k8kjywuy57xl7hdZSSi2S
ZBH40SOZm11+1Q/43gsSMcj4Exy/l/m0a++PkrG2w32gjyDmKJyal5zpdkjKRpmC
DCUMIYWUSpeA4eeADnEnwZfxt2uH2Yc8606UsGo9MdTo+MYit5+pBK9TqlmWCXj3
6ke7JZlZZzgLZLx7LVR61nmIE8wF45MBxBWsdVZce+ELjEoRvBhe1n4PtKNJQPD5
JtI+hKqUIvmlf2RMShiaOjjiVxlDjnNmxbNTY9VaVq7H8qX+4twKTa4P5DfuluM6
lbZlaTJssDZTriNX2FC2H4+uJX4hPHIuwxnBVAGi41n9nfyBuvzd94m6QNzGY8tL
ihbQKfox+T0M/Z/YCYqxCZPtAeHSfk1KYv6oAt/MD5goCGLkZuLtDwLlqRL4gTDK
dUtvTAKUR2EcL9oOLLHfMU5UrNuU9z4p4W6oTyACQStx8apEVxJVCROwYjbaGUCh
vgBRpFg3c57GKBuZkNKeP6MdTkxQbwqO30kZB9mfsaA2Oz71w9gtAqOWwg1twYn2
kj5uT6OlGo7KvE3laJ+ViVi+93wjberQABi4dfCt4yFniq1hrmJ1fVtaIN02vieB
IjJaArbpDW72Ah4QfcVsdgn9/MHLAyQY4Otke5P3JN+HPjeAxOYSxftZAzILAa9N
pw6f+O8TmPXT5JFXEWEnITn+iOJiQsAxA+xgHTZuNf3rNfB+8j9QSWDb1EMjivs0
vAe5ke+DmiBm/NkT0qgGuBdGtW+KE4fz12i7rcroc4dyy3689QwzEYmOlfiTv1aS
FZb1ds+N8qRyVdu6mUVVabPr4d2pXdQc7cvwN3SEXXoOVQkRLmuYdichjAuQRoDL
WnVfgFgrYXtaOu9Kl7zPMtn9ASp94Uk1eWkdjCr2gVxg0buzQIrB6dVmqHAzlYW4
ZJtE9X2pTgaMfx+Onz4OpD0z2b2WvyymKNRbFpMGJ2elDPEGkEv7bq6DTXUtvwV/
P7/HfZmhf6zc3Lv4U2dxhSlIgETTYQR5SBIvyoPoizr82vQYjmk/QI1a6eyXke/5
txIcy660mLK4UEROmkU/okTBL1iofZEDFJAArUSnnFV72KSJlLLecvisYszPltn/
/f1Wq0azW1oBMcN4xBqmKYSk1H9KfNHoOdiiVrB5Q8sS68GwRb2BbDr5s13qE7IR
8dOILxaqMn07b3gqRpUK2/NRRuimgEOybeev21wW+qzzU2lby7G11cJ6jm/bZKV4
QP1zegsv9tluEY0qSAg7fL7bSU/tJLc4j9UBiWs8w2OGGF8A9GMOE8ekowL8m9XL
ydhuJiDxhDgXiMLY/SfKPD8k/LdZ9ya4yrPmoi1YJm0s9IMCaGSYOCIGxH4cKXtS
yTOBW1uUSTpPi8W7H0HjWuPZzI+OLTU56XDDhrAZGMJad8L1VnMW07HvuNhQdQ4x
VuFWtaMtsZ/mMosamI+Pplw1xyRxEt/4pRGHTQ/kOF7we6UH3vlIyFokP42FbtGI
MFxRj273ndrN9Kp2qBZysZjKcvBU/WMXJP5eqMnfQdRRhv0JdAmLM5e8pWc9fkz1
Sh30/TF4INRJTqQY/l384LJIVbzYBKU+QdMAChjxg/R7cD1SMXKC2RaiijkxlBlP
x3WvO/kjGN1fzSGKxVMylESgPPrUTk9sR1zsn9DFt9uHiiCNSAeQMpRSs09fNcBf
/TojmTLUSQnJwSs5KvCrL1GhmoaoxFqqK6VLrLGqmFVI5At3wIRpmigDmVFdcTRe
luiEKSPslePPkRoCsSOp0OEmyjwaytHhrpAs/qVUJz+bYTrwjqEdA1YgEvb62fBj
M70p3+C55yNqblbx43CMgUJ+tPlfk5H4F1yLf7T8ow4FOjiZzOxv2SPoN/kjhLkW
L2sMfXHklXRl/1IfL8maQvbtVeLE/LVE5salmmRrsT+ebJ85w8Nhf870Zwm/tr9V
My+8o/UBf7DLP5xqT6AFSgAubZimKTB3Xb4W3uE5lEuTsDgVMbD7U6N9Gq4aq1N6
stu8+KnzTcZ0dH9LCOzEEW6wo6+4zKkrsv8tyzWLJSQAlPVueJ2SzQnNhKTNsoOZ
b8mSddDYp0227Uu7vzM+jX3dsduJyd/nraHGZgxS1HYsB5WFB8Y62glldIMmTEUE
wADTxZ1cgZBwB8RynvLsZgKNCyJL0qCKYlg6Q4MqU0GMFJqDdbTQ3YPYMhtV+W9m
4sIqREO3IA1zyO9rVCw2UiEpw3gzqsiD1v5co+q7sXeUeqlvupUW2QIZAhOu1V/E
L5+4KmiNn0s5HzkGSMKO4LAoS7ynpvZhOfl8eVq7AKrczhwfc7vfBbfsmkyWbAxE
BaDRV3e5ng/QDWDVoSuOsqMq+Kj3QI/DY3J7o6bAYTZK/oykaf5s7QKAPZb/PGDH
MYKzR1EMliTkD6zvR3IwQ6Nhv0wgYgFtXcTs2Sgovip2hXoE5F5LPOwyWS47r6yA
Bty5rNJWZWKuCJoCX6EA91AoFwZeVGPHPxZE7eqiFr8izcxY7+NnBThGX13TjBlR
1GYI0tZBqtRiBVTJu4OIKCQg9ncalaRSFrEKswyxx+qcEvLl7sxQTHHMBttdCiep
m6U+Xe3NFMyoI9ongvEtiG6R2jZ5+gzfpjZAyOH7p/V6SzLZjSq7kddDCEYiWv4s
8mx496f4brAb7Mjqel/uoow/Y/pxXFMnVpH6frDKz7yTBEblbXXl092FcuK6fGHR
aYh6Lt5ApKDTY4K6EHfhygYrIR0+Lffamc9dCpEFe7OCViMVyDb8+3Bqb6HQ1KJf
7+DAOJfZyj828DVwTsjjyyU0gZu+i/8nPNUg4K01ZU9pz8KoAuq1CpqY+YP6hln+
dHeDJDFBzbf2zaqZzsA7SI/RsObTWXLrdRoLMY7WlrTZToT0Ra7TYOy2VDQyEqqw
jVoBlQaFwpwjlik0/bBTUD/f5Ap3p2c/oYdJOQ5B7UWStSfuinhkH8eUhbng7M/u
+b6fJCl6IE9riQmToAlXqHn9Yas2CBX62xvhFU784Br6Gcr3Yhi4IYIODGI4bJzi
MKZRxQSW3cI6GWoxgIls6Dr2XhR/WGnxITs9tEOn3rqes3uOJytMcwAt3LjCFJ0r
FHWLyXudH1b6GjDuWezBUZMu4B4hFtob8RiS2In2KeLxf3eQmD8jmCeBu2Buhl4r
cdTi09bGo8fKGwrzoyz3lzL/j/R0iN5Z73v0mWiUraGceSpKU9Yvfiou2xvdn5jV
C6d9dUhJzMFPRBzKPEJtvLIvTgM96tCF2jAyN1hPNbLxKu+kqw3uTbzPoOeDt2e3
7zx/NGdIxZVWPyS64DwkTtMmwXzgJIwoS4H/L1+u28ly4zUMl0z5i1loIYGyendd
yJTWXye6mg6jFMxUpHTyQxEtmpiR5DyGmLMbzkNAvVRFfVQYccZCRfBtmBtS1mPM
jioQ6vHmfAVEtuRNXX1SCMnYpyrbueWymcq7Fsy94ka7NPzGI5hiRJ82koM8rp//
oveVxkvfN+ZokmuPnmvAPCektbxabd6w5fm3OROu3Drfw2LWcAp3zmXW/FS8cXOv
fEZ7P2FdUh27EAI08JRWmQ7OnI4KgEk8tcTaYdVjKH4gq7X2rcurVAZLnEkcp+Xm
U0TBC5joCmoq+PM4fYcIjTFlJmzU449sHh9i/B2rspEC4obT/FNRElBAzzAzOj3X
0vluuO1+zCRbyz5eABgnBpF01ItCV3ACxsrcN0vFcXE69wk4ADmuFSUYg0z5F4Aj
ebYD3SArEKR/e9GioTul83sXRpxuAktMjk8FvxTu0GzWX8tfH6tQtIuxUh77vwid
30AMGrPlH74CtNghKT7XjOeqPinAJHVZniN4wMLH1x3PzWoEaFWV7daMY9nuUDUW
6CSRx3BXIaXwONGx0E2LVDpDSsxGLlCtt5t5mNXFvhxoee/hzs5svMbOn12/38yT
RkrCs4qq1Hk1h2xNd5RHVa7JugVNIw/FPwYrRxB1Lj5jIrQSE+bepyzVcBLr4KTJ
Xm9XBOmjeiyq+zu0yRsjMNqGXRN2y729fm/kC33yAMbth1vzuqkTKC8VlFhs3Zd7
ZJX0+ChKg3xkOzVec/ZqJrFpU0AULUijgvyYIm/lHOsqRw0M8Opim/oUmGYdCF7R
yB6HUDEXfTgk56j7xTh+pZIQn2IKVo30x68yarwccY2zI3taMdsDlkzGcQWYIn+P
yaauK2NARsDnVdLnxQjIRfnUxDAwVmlWxa+pYdTMZdlQj5gpVh4Yrems5Z4VfuEO
U9WApUGfMNitTVrQEbdzY+UIDSSHU1+z06ImefoVKjf7EcP7R87ZYBwk8I22Ms80
WhK/BSAr6o9zKyP1g+F9roiytXVsY7PquHkQgCYIZus68F4eQey4/Dhq7MFc+DZV
NF0HSxWJEPKaCzPDF9OFyRgWiAQftVArrMtKbjfM5ZnFrQtWGxaC1DxIUxRanvSX
Zz3CPalEdi10XFSL6EYXgmeVmOWIehDLH31kh/eCYN+voVtkR6C75LUZFQOoOvc5
Q/jCzhxxSWOhSBervNOOZYXOeUX59O24HQFqHwVxaNHy5aIGvTVuFfcFAD5QMXAM
URXXWDV/IVoBGsDiyN/CIYhsFvrPcG3Tv1pLDzNFX5bkco/ShgWrI0y1ChymvGa0
m0suu9502TdihEJrwTOvVnKpBiRRq+lj9vVZxgSGPyeEoLXuME9y05mU6Z1I4sj/
GNybn8fzAQDM2GgTGTvXG7Y5R0aVECXCHfoJ8zxn8mRgfWREIgLmewc2cCmguSrM
dXxviSHywaQvxxbEMnn2aEQIH6VNBAujmqucwb9jSufpcyyXp+ErbZ3zpJb43pvp
UU8U6qeII//GKasL2UjGRtxapER0QSVKqUm0UZ0yPK9rbz6Kz4IQV7c3tgYC92gn
qnuNyPJ9bpXqDGiiTAACj5HCUhtA40om7LTyO0QflZfTDA9EkbqQlM2vddCVspUR
cMaVA1RD25IljGw0rN3R/tT7JdwvuSWOEpPM1xuKUyou+XKd4TZ2AU6H+JONLR9Z
QEPasT/hcEu/6ngR6pCqP2IYD2LPMD0Z4r96250/5sSeZpRV9Sb7x8yhOAFsnAnm
D8L8Is1k4Isrf4upuovGHqksG9Ev6rTHwuiDZESZCEiKpmRGDo9WaK7q+50GEY7K
GZCx4kOFFzoFQOBWG8rjIhiys4dHk8eBYPvEO7EOGYU0OW4OwUE7S/OwfqbzE8WZ
wv6oumq2jBFbZpREn6tywtl6wiH9DzCCfiaw9WDq6P3dDsOWiZ2IythqtKI/yLs1
gP2l56hOv9JKUx+7eyxTFkvCoDRV/u2UK0XVhP2Sgh96n+K7JK1/55ExtFWyksWg
vna+yQbVqKlh5Wy6J97XD0gJt1wcJJ7GTAJJkYTD3mu3tvaxMEAEu59T4EyMtdGE
gj3a0X2UZEWybW58ZhcuxskhWGsNLyH/fLpXOem3BGHZm+5RMITzewzOcL4v6uJT
ykPafaeoVG5V2GRb+akIGdcbnCsPEY7/GXQr2iWVAjvzjSXlmkl5lqQsZze9F1Gc
yz6NJ+/b4oHOq+1HOEWtPoqzzQWd3lmNdWVIvfnBtofeXnJGHnEj/v3TVBIkvITr
jqRTRgIIIPh8KF/rTKcC1gE0HC/POaGYoEQ1XL4BKyskZWE+BY8VbiqteuwBv1oI
M+j/xw98z/wEpdnCIAFWzCCo4TJd7b8T4fhvlFBm2VPbZvl/o5Ssn7jgXjg6hTjE
r3UPmMt9DYnPB9p4GDp33PN6paP2b16qza1v/LWmQCZb7ccyFTfmBEnMkLqMKQvr
l0a/31t7BrNF5SkuLWh4pCuATRbAWlCaVRiRq+Nw3XV3AeewKyws4T+3xdYH8whw
UXwLagWz52+F1CUXfbpHhQtzcdLoGa8NFgbaeWVWNW/TrPqXEWFqyCNZ66eEpbHC
0hlpziG52V3KoXAnHGmSA4uBxNBh4CUINnOs63LQzJEkTMKdwgEfqNe4ys8Iw6DU
TgkU2f1Xbmy076BAtilJGOemmJ52roPaRaJup6avL0jRM32duf1yGOoHmlMyAN4a
2C3MR3oRnjHghKPpAiFO2WBwdBXFPLtpuMtavx4pcJZ53jVHHdQdHhYwo2YQfW6f
dUtXk4PVFOpFqyTtSeNIi+ahOt1d+ELAF5d6L5c2QjyjUXQPRFtwz/wZaYeZOpe/
Ia4VWXaPEIsxoMnzOWjas33nIhk71JgooTFWbiFPoNU/eSC/aQLhQrRYvwZk9dmM
oZYr1a3M/83jdYCCPr2i59kbNlSpq+XSUR293HpfeqKjAeBstVt7NFeHLHFXpj59
l+c4wVDzgTedp7qPLo3HJKlPeZlbDvGGx6twIdw5o07eK1ApYLDzGRUUtN0lnb8R
cgUyF97PJCC4g06ufmbpkCUVEzwPai6q3ToXXe4B2qSyNpgKqkuoAbE+VSfz8Arj
3x1SQJViBusKQ7+F9/oBWd+mf2Hu1AApKdo+oLJgjtG3n59gvk0sy0wRsgogVpbm
2jhPXOOPpm+/hEGiWzOJnciPEm4bIUs1lTOaBtF840kmEprfWZCJLudAw3DGocwz
ztC4PqjPaEzrS//aUQwhDxmADj7MXtwgVy1af1Bv71mgmNy7IGq0AIEURgBQ7Xq3
TkXFlwIweKh95h8SPEUtn0Ihc4iEePd1RAlICGhUr2rHFrh7hAbQHBedzY/L0Di6
m1LPfsd7H9LJbouZQ6bbakULK3yWsQ3wjOvB4O/mKhFGnsQ1w9SEOFeQVQWCvVvu
3fzfgsCCfkOM+6IWgBIN/kjZxafhS8idg/vtoyRPzn6mwxu8NCFfnpXo38ccoFk7
js5Q3o+HMbP4EVc+T8I5LOmEcPgE2T6bAv+3SsuJBRyGRio5Zwh1fW/LL4injNCT
CwYGDp6Je+OdBIG887uw1D+P761I2wLkPiQYzgwvM4AcUUCm0tO6uTi4VwnwOYZ7
EBSSW/vCXs741waknfVql/wYJI9X/Dy8xpbMPc6upNqxu4xO4ZltuLeX1kjjVJSs
RwJPUOjQkR0sC0DfbrgEHfnyHoIVYdoUSSZ90Tf/LAMqrTZ2ckHdGPfFrM3vGt6O
lgMIUIk0ERAsp7z8osY/YNvgneKX1CBQ06ps/Y9l96gsL5avamHQz0HO0EHZHOu9
O/tSWx2ZtOntjk1vcVPTuHYf9hNpdRura9WnPTN/LXDb7xdACAlRtYmnRBFGyxuc
jXHVGELH2deGD58dW0RWODzonDvNhbFXJcWrFwX5yt63d90gq5wXiqi0gLFcyB5I
ceDSNlwlFlCzIJsKuv+esky7m8zz30X18Kx1nMcIW4bT4qeYosRpAopRMwuJn6P5
zpEFeHpdI6fK2QUQiVyDurodx2UVQllu8ksryLJrfT9o8/0Uu7iZO0G2nDSCI0dr
jJwE80jntSaegqGuuILCUqxc3ew+n1qjnl+HHHlj+ufyuhSXa8OISU9mXVQXo3YW
WP5iz508JcQiF+5yCQMBD0cgnzZXeyWb12eItCFS0LSr6oGU9gUKXgDHQCrDzEvM
QXYJmQF4yUafrQepW1hB3uIEFm7EP4t0fXAyJ+v2tPcbGsw6YC8L0hy8ftEuOsrb
2WJPcx3SFd1bCM24p/Qujp4jwXxzwdLrB6iIrIZMUuinSUinoVvrgeDCqs5oQcEX
vjNTqQVfPKji8ilr6XWKBO3jvj+MbcBQi/NLOe0f1oKv6uY7JOjUlqv88ncBzm+c
xmxXaF77CoRciC1C+8LMBp9VFRGLlBDW0aYxkofRlLtpDPxB7UrVlJK1QGxId9HZ
Ywu4hC366FM2JeGuDphmj/ZQY7vLHPHHICAkNHTugmTg4HKbhQvJyd1moz6HKjDe
K8uFdwuTgIq15gMuoKThR1SnL9ax1QyhGVk/92lZQTI310Ix/Z7JbQhBvlZ+YxcO
WEZpwj3Nn1DApSORSzLOi9U7j1i0Mi95KEdyjgioKaRxUj0pyWrGBlEciEby5zM4
U3o6i8UU7eYij2zT8C/I4umHnOFqoREYb2rqIBdr475XN66iw6yrgObqIr9SllBV
M2g/+JzTmCWttBoLYz4H2U+r7KU+fhDt+DdIxAG8cf4H9J8NwzApFIS6g48EHJC1
sDR4XerqKvD7wLg1JLi8I4QhLZTSub99/JWoJvNH5BeXLfZqnUeHz2Y0bAUKwX/0
+twqaWvVPqgWrCTIj6iSPRC9rgidnjjvB+SGeMZqnTTrWbQkzexs/xym0j2sjDR6
XnyGVM09HbG62R/RcvXlrSHm/3uMGT4RqgGkYHQ6g+aPKhdZjGpqk5gBwhcUilNW
O13MaqSBqAa6sxFjWm1WPwsHo6gLIe/xSDOKmPSIkEoLQ7mhhIahtL/obytsuZW0
QL7lx85ti+jXOhw2AqrCrZWpSC+Si2Ajv3bf7nxN1tNs7F7Q5We1u0Cun40Bmpbq
1UOn0jDXsUeRSll1M+ld68YyxfNP7nsk0sTCAK/pVCNA3wP4YJFCs5pCt43B+IHh
ACCm4NRtJu2sG8VJB49xKDFKMNiD+REr47YNKn4dCPSaS0X0F7l9TMCswilyuZZ5
qfZjiaUOgZ2ZUkGG5WEp4+/XHkqHW3z+jND0SMGMlb24m8TUNZIpP91ncpzDj+wK
w07a9By5I+U+CwlHtL+2WeOKl3Qnk7bzLpC4IPX1dUxTGyILmwkUMj66epMg/xMt
WjoA5TJI1FJ8BIr7pHkyigsZIU1YORMAhTW3V8dSvIwaA3XkLxE5jO8gePRC1+sh
be4eMLTFyeb/6+JYUPiwWau+zpEp2Zh1qq6cA2lEJy1/GRIXHLo+/nWmZfLcMrHm
5I7nxOpESa6ct/diLymtrdcZw0IkhLmZDU6dLObBAowttjmHdXsC3f3pcV/JyjGq
iRCMmrMh7/uLLbiWF+5L9D1L76T/eksAJj0QklbPpcGDt4pLc359SHtH8fjsOQvd
QDeiY5hMI/uv89FNSCAc1Bp6RmdSPN89GT1DNNdAaofFn8UzN55UOTWQhd5ZpMPT
k4rGeh5sbZERvQo+NJzxvdvypYoA4VD6Wyj7EfW+r/ng5hGY8kf/3jmUunIq5vWo
RiY3navpCMfVLLU3EjsS7LFTBmoTM5vyg2ysKS9Kr0h9xC4itiNJ5J9RZMtl7kny
Cdw2xSfl9sJiH1XCcopkCbDK8cSr4gQlL55MOovshcRenQh30cJh6OniHA3JB4pC
zd4ow6CY3fU4wEpgQrmqtmSDKCe7ZdczT63MlJSw+mrjIJNm4XWq5rICI7/wLEWs
Cl8WT367vimcJ7lBr6gDFgKmXj+ikCPv/V8vmA/9V3vS8/F8ZiK0mpsHBwO1OK9j
3S59db3C1CYNN3WyXfTqkRoa/u10BXSVNdPnoxaNGbul5k/EIf9PhZqH4fwKVpJs
TXa7O8mhYE/687vzXDj5pfNEkSup+Y06Z5zhIY6+gANsDGoLU69S3Yabtki5i/y8
dOaHf+PYW46UCs/fuUOWLOeZkLTDKXj5PE1DybNZz14k/ztQN7tgUd9JySa6KdAl
gPZDyT4tgmJajUdFRq5+oOqvMYGKALNyiMguQH4qA3JVxFu66p2dIu81CQPMMbOy
7hFyFvzltF4IakBjxiu2u1plfrqnpMD2j8ZF2ZC5GDaNaxchE8pjbkVbzWk14w62
fXFt5yDeMttYAOu0KqUj64D9G9ZkYUWSASPr3XN5d2O38Am/2V8JMt+bfd9R55uo
DWnvSfJpngFl+ZQuyvBguZLS/t3DXjh6HyzzW4XdlHkzMmIzwh3W/BAzhI9LQLxu
8c7S0pG0ovJXOpa9oo+uGbHJtvFCB7IY1gmTdf56VeLYtDX+RINaweLWIob3Z9JK
5LgpSVjDD4C0dOGhIxIbpZaEFCt8e5b1IdMAqPBkzH0s3dfNZMSo+pPebLyHxFFY
eVBLtg3CKhzYdFma34sm84vzY1cKYcN8EIZXNTMnSQDH6c0/h5fGc/hjfJdfcvOV
5NJhdrO7dIukp0RdFT+VT22xTsCklwtBo6FZ2KCwRw3xwJHBG9fL9ShzNKB+/hwf
JPk7c845U5CLbYGEM5Wnvwp6iFAitego0YmEs0uwp91WJTClqOqcNmfyAJ4aeKQH
+QNds/glCvy50FF6Ql5VzFiJRqQyBdPuelHxGNBEA6G8y1fuAeIL3YQN+thGBgxi
t+w8J3p3OB9uPyUmhvJTb52K4ayxNECTWO475ZjeQvC/kQdtfnM69Ej4++stLDHV
T1HeSay81QXgwvJdN+vczRnvwYe4LzCAyOOZGjD9Jp8zFwFPhxRgNBmwiY5uB8+i
NDDf+syw+EsvqeA04/rNtdWdxdmN9DfJLqJa2wWQqNUtkFd9uhbsNaJMy6NnE3TQ
4tTxqyCTkclfjCEbI+gcpe8DAs2hC6R0ER4d7zzQw7pFC1ibssva745bJSQcGwL1
uzWRQs2b3J92AJbkpmGKHE42fuZTNSu7fhJo8JhKsFitm+9LO1gTNLgVlleGuSIi
X+4sv9N0g9hg7VrUh0bKG6T6alNAdPx+VBupr8y0vjv65UQ46AM5vmFYdBiCuc9d
TqBd3jSoQecfuWPq5WbWuhCIGz6c/1W8CDbUUkQhX3xqEB7Ptp9lQDy/3ZB+hgIA
RhQej+QoLuzua88AOvFQVB6nOT2agc2+xIzpRFMOD7UGQUijW3cdgsJAKy8NckJW
wz4JDHnePOEIFl6PGi3SHxzdL5Zzvc5H8/kaGVHzDQhOmnh16+ws5Yj/kIcbiSSO
MutFNikdS+CQ9R18oFRvkgNvGu2PzdUztwJjB5huzPC9zPuZ5gf1zsuzGN2/yqCq
xv6vt5I563VmhZ/fOjJ69CfMI1mGnmNTYs0IY1witY1Z2gRd2WTo3Uzd9mpNRUcZ
zeQrAHcXSkKZ05ztSsHtWZvHOygh+w90X2UJAmAwo8FqYVNM2PHVzH62+b6QP2or
SEKoXoZk4+ZeCCphQ75OuMyog6pDg3ZU/xpHHpPqIyiIhTZs5d9SZjzuVeSEQprN
vZS4aaL/kZgdBzNUbtNArPbmHBenJJOw4iwcyFYTS2Wn86V5l8v9+FRrJQVjp0tI
MIN/KtzaU846WyuRXHgoTPsNOKJHb4onQfnYMeCmTj0fOyoTcV1YWmeG9btaFUdn
bKb+l+Sxr4Ue0G6jg0lRQDKE8Cb8d10THkZoE/rJ1muLa91bn226+Y+VjDI9Ja8s
n6iUr1jWpjnjmj2dgjcnd16I3hYuWCkv+06oBZI6LNNWafU45FZF5Wknu8dWvWYA
cMKTHWXuEyoeDBlOZT8xHfc5hX8Qmo9OT/02nTSisFHRe2EsSI3PWtpyJDuv/lfN
TMu7Zvep4DsW+yaj8Rd8LZNViJuGFRLhz//jHo+vWuSUddo1zvt3yTax3chn+IJe
RSOO/CPSpP7GgGaObEwK2NMzwFVDC/lNEJ0fuJpxvwJLKjMuBPqiHLD4kWj9iHDB
rSKqxr2MvMmfM+vEoltSYEVHvFdyVqQMrQfUBQliwjlD89egZvT7x14zT1DDc5ax
+KhJccCE1S9KSuFRwBwjqXSgwGYY6V0wGNXsmSEycP1Sc+2eflG6j7WatidZooEb
vNClMXEhWKZ/380+QyMpEG1vEHPRV91IX0xYeWCgUh0n+MBjbamY1mL4o5lzoPP5
g0BV9ue6xy0sFnxTTLiArzxtJHPf1bIEHTeqixbCfG95wwiVKueBiDJJW1ShmtdR
EeCFNaw45wohOhNEsOPfuBlxSJsHNtP35TAwyVuTmUHw5yKahlbynXbOtz2HDllM
lgAZI8txHAMla0knTMJmZ3AuCaynjlMF9ZtqgdI9Ur/yiEeHkCes36mt+cnp/xUi
e8hmbrF/s9Pf192BK3fLVwMr5ZlI8Mlht+ue2NeyHOkSsBubTS+AV7IVlDcOe1z/
UQxy6mnYxXr4W6pLQr07EPV6ZoIa+ixVcVrt8b9R9Si7ypa58vJJZxBPD4JFZtu7
GQDfeFWRkrekA1SYMmeAhMo5pXIeJT8BJiXnEOdaFENBheSBiVmboV/aX6TaJYhO
Mn5KrjiZ6fzhQW/bkP8oKqiJn3zFvETM5G73QhB31yOd+bRE+CDrAzd84dmFr/nV
imPg/6moT370xXwX5PxkYIB+J5Y3IDA7kX0biVCaaQFmtLm5F4HlyrzPOW+Nm+eO
hXeQgG1VZ0+OnYTZ60wWLZela3EvQpurL73l+5MdKkm9AOXLqu7AcfTUDuYEtrMc
kxnV5v4tuq6mgg0QOmVk/yDKqkrrECrwDd+Yu7hclwmhHU0f+V3Cr6h2hBkniQLo
BdXthYf35u/GAFUlcRBG1El+0GYYTOk16Xu8KpXuDlHh/UE0ZqzRvRyB4bijrOnh
uiNpdpUQlDLRdX1xi8ivj5omejcevql6h0jKyxNB2Z4wkqsdYuLTPJj0UAiLoQU0
tBPvHrjCHufeLyJqpUnNDxbRh/fp9Bck/KH34KmXj8xcuO0yBXn1lFYarQGJgqaB
HrYe5CnoZQd61pAbDU4lWVC97P9OoA9Lu6RjI6pCGsDV4/HGmGy4LehkJCqDSDQg
RXesm2wEps8OV64WBjMm9y/uwGlHK+vULWpk3/9GOovStadpza62gRr3+KPBFv4S
O0j9nXKdb6ZjriKV4cmTC40bLnxvmIMCJw0dh8T8/COqpt52FWNYMtOX/IuPju/Q
7tORDXYF+s2MtFukLO0NjuMRvKd+n8QuZfHi+A5aNTZL+P9ym7pG0+hIqbNgco85
jfo2yhifpAioN2TOIMlyDCyydSn5LeyYT5ZldsEVt7odqB/QNoM1iRbRsQzm+5sm
u0fYIRVWy9KmDsL2KvWkm6b6deaHISVzOx9UmnphI0cLBFh/RA4nwHrPlaAPHJo3
gaHqkLiW//NnkG5z+6BryHvDiYzyuY1edhfcmbRQvOvXeVrocNp+WQfg5A30Xaty
N0roWEB12ED5jZHBHIgAxrP0eT8r8qHwe+/6wLZ1tp7eMpIsF6L9A5MBFWanjcHE
zXucAtGEoXUP7l2w0WRkyEhET2okUcRct4XaAij9e3lQ+1K2t3SWtrQCu6IqHCgZ
kBdgkzunKpqBlcyitB7InwX1CE5eFlOShgKLRMQukRPXRlYGFQVgleSjX9ftuvcX
A3tsBcmt2hI8fLRkDknU4NhOFKclCnZK6KbtxMlPlFJO5pW2108ZZNjpv9ki0tzs
YPqLFCgC8+WmxMvxOWQw5V03MIZLlowkAZpGH0qd9ugoKa2fqvIyMoOjNPxK5Lbp
E7tGUFSCFOX7QNk15J0QEGZiX0hKsY1Epbi8ELpF7sMW07TY3bqI/7yvCVlwu8AS
K+ZG1TDlhJ8T1nwGelNXyyHFp9BU18slFlwvhP/87AJnQMQ2XoU9ItbN+D4TsPij
kWxuTs+cgoNhN6EyFhNuPhlY9Mmz3B76v/WDxlhkZLrWnHvwcaAzFt9RYq5NpgBU
rjMcls7l66q4rFKbeMMArcTBzXuocggcyt1C4hRA1rerZc5/JMAGp0zWaEqKKA/d
P3wEuN5BdlcNYd2MyQ8PCCDAadACKmB6kNtvVhBzUXhIoZtw77wYRzAHZI8Mahwi
CEEeUO3rbpihfnIC2etuU3mQ3lIvCxkV8PiW7svcOe7NinEvlndk3zMfyMEMR7ZP
vI3ZQHPWhNISv5iFvAT6UyQjkfwZCPT19Ju5rxTHX30im324kyRUZZrYQWoZ3XkT
EtSRdBmnRhqv2aMJALvMr+wnYy8HhHX0HF3QlFO2cRqsLRdho9RBZyiqfWKuBazo
z3gFIWAmmNEifBLoNDbMcCj6Z6YzZG12H5JJYTfyZwssUPKQ/D/VP5S3KhzfM8s8
hyGcmijbO1WhJJsBIKIR3XQHjbYI5/SgsMMUIYm1A7jWz8129TC+0A5z1WNO/wsz
VLi6q65abHFBL/J0Ft6kCPLAK0fjX9HmKBdCFpUyAXHhhv0njDB2XoI+fu3QP6Qg
9Lvy1ljoSa0h4wEe8HzI+BkuehhS13prkaAtNRyKn1/r8Knp3JHnB2hyRitClx6+
pQ8dU2fnGSqjCP2T/4CTeBpgHVT6SPyPRUvB60jP/OSCf5WM/Byik7Se4t2Ib1ha
7L9WXijLVWqYOGmTRwggUeb+avYpFYWjJQ87aEg7qPdAvOPFSR7lgHwILgWhni8c
tZcLb95vVcckAVJH9RKI+nVQVlfFo9/zSDrokRm+7l0tRG+EUXY1a/yiZisvYNtp
d0Kq36uCi1+JaZ8cuTZbhAPFaWqDMPoPGqIXnFgHkeJOevO67r0qHgTgKpCx9G0c
JyKligSHqnCJc2K9XSi9Pe1Lhds6qxxYtfF33Ui7gKbwLTo35r7gDbUxhiZHjkAj
+mW1Mi3NT/7wD1D1SDz8tZ1tQVEmIj/5XgTcB0EmSKKeqRx7iUgotIf/ljTwsjM5
grtf4OFEEe8QH7NO+6QZr+gbdgFQxmluTam0qRa+eAtBLVnDkJpM/kobR8l2ORIK
7moj0IoAZlEVo1nnC3ydRwSgzlLl2owwHLhjZ9JuKYrkMVPNnKciyvqnMVay5M+/
YC4tIWkNf4+nw0T4HVv6498OReuUuP+s1kAZ0dyzCBId4hdG4uP0hIieFMLtNaph
un1JeZ4mQT9t585kiez/MLAau0ls7Y525xsMRPv9ff/EkR5MNLLQvL85lkqrkk0p
tu2N0g0L0K/31sTLwFF8v5qPCeyCkjJnfK5COCJoExAJnQ1MbfG4XhThGq7+ieNP
ALtM1luqXEh6+3QnwszPd0E7xuHzpe6PIBVchRRKnp9fMBIFaSRGTEs00Nrln6yL
wB78tm2GaBBNpu9VraV5DWMONGX9IpU3gaMVVwBsJfToi8CmGpmwxZ4mfSJCbXu8
jSIxJkk3eDeHQRF7Bk4AbJ6f7F2U2B+P/mmxsHgjjxTpuucdvlgA51UuazaiQeO7
wTMi31OttlDTU9EiO/Hcack/nkTTk7JE4q9rci7MS0LHo3V943ahprn0KD4AFEiT
xoWIbQQ+YQK2bcupSi73t+FMafwtX34k7AJghpcvwv19cpO3r6K5gshuNkVDnrYm
TG/IHNP36Qco6DE2Fs0AlmhyoTKsQ85omNribqmBXYE+CcGbSGZORebMgydJ2zle
dwjjKsEXv7w6C1egGIj6zd3kV752KkXE6jYpnhl08RQCDGhgdUlBefQkjtEuWfBB
3NXm8Ph92BGVTwfrW2R5/9hDoWiETwJ6vgz8gJyjJuFDH8N5/2d0ozNMN6/A7DP/
1QAJAv+4oNG3MaOM4x2lmWYAj0KV4TwvKz0/JaPZBaHG90BNxthKICkEkzUMl2/D
k7QdeyPH+ojfrJFTkvGwCQIqb38lNh42IsPCX1imOKcm5U0hrtGsQkaWD7lyoOjJ
0aATkIPKey6ElKrYr18YMSDBjg796YKEhBwcdeUjIzbhBs/a8xZzfeNQSyG/JeYa
YrJ8XwF6etK1cKwEQPNzJ4C//fWLupro9hHQ5kpbDrI1xGjcn4g4GGoU5DNezbgt
FCbOuZUPrdPxig1esy5266pGxkIbcsUSOtigSlky3fLnGArM8eLqBR3q8EKbtuTl
O6SVY8idLwYjJC16X2UdsUGUakM8UxYRH0dUCJ8mkF/wZvNqm2sE6mDEhdW23GxH
KsqBI2d4LPg+PAQF4I2xQWRs9eS8VNlIBifrbJlCIBUBY/CNGsicJiZQjhqxJwxD
OfBTQrl8N2kHv5cGwO0uziy4g3ET3uwqcBEQ7XVJG35Hzbf9DbrKJ8Bz6Sal1U3S
yAvnYapgApkiMAcs8kHp7w96JxjY6yv/vC8h4HfedHRWe3hvfHdOHUOp2xOiPrkw
BtAzEr2XTSRdoT+nyxkUe84yYCGLUy7i3F8PW8UDl9R+qKFLb0H9tpORvu8qKrLK
0K6IIe4VNQ1Gh/2J/UCL1G1R44h5tsJOnAOdtY4xW3Ij5JJEnbLhjcts2Jt6R5LX
KMQ/stmGm9g32QXqNrYNfNsdDlpdRzqL9iSW11o8/7p0F3k+cYc/7NddFj6fhqUE
nUdytb3A1AwTm+LFVZzjp4iC72KWcNQ7+yAyCDP3r28/YkLkDA2WtBr8aVpHhp2z
JHSRHoRHu6NPXlOOynhpGCmEgbzdcfROsN2KoM0nE8o3BTUI49Gzh7Kqs3oWcGcN
2b7OR/TBwNdkl1om7azNnF+3ppBFxhCkyae/Ir8bZeY/OCPCanz54Qw1Lf+YKcnr
I9O6Cb8FohG+v1QTveQuIQuRpw8TlPt0mafW/hvnkff1nadxqgR8extbfZQmOSfl
R0S4KskAYclJs0kS2auR7yYdLtWagorB+zMPMUbbCgAdMyURfu6RfyLD8gCxLTJS
TbhP3ZwmCHi+VGnLMl0oLzftUW4gvxQVDvQp0igCdFYCFMuRxJ80Hh+TkmO4ce+v
kSMQA71tPy1PmMVbpKwe9x8mJnaYp5DwRKyi1SSo8Xxk9N0vBHvrBuxUaNknZAm+
kW9MSJ/JABAzv5lCq3m9isSAY0wOznORJ2wqzvNEW/rworogHHwH4vz7wZ7S9H3f
fveijeC68lrS7MH3un+W/vZYKevKkMrinruoDtnCugeYABric5kViBrcfB5bBD7y
85eViw3J3Hc2veoscvxNJApQgc2nAy4ZsJgeEh+MImq3hsEkt/FzMNXaU6U3sPnt
fGBR2wgRdBeL+yZMTaI7a7v+gDumMYXShLI6ZNeBR1hUjufjc65TS5+Zl3VhDEVX
4kZEnCvo7Y//VJZPcfmm4ZgQ4YsarMpWFqqTy41v5JZmlzJBD/aeN8BU0CCBlHVB
PgVoKBBttjxVnFOQd2kqOiWc+oVJ2A4+Wdkw2n9sCQQAm0EH4aQ68K5XgkbP1NO8
sdyV9EyqSXWEbi7X4oTaJBxeFJJvUjDgxN81ULw3VGxvxmzl+dM/PmFQCKwPq9IJ
SpxKLk6rGOm1QpjX27GqXtdghYVIfl3tl2b6VgHcsOtVOCxrqEG4+mtdjFJrvKtn
ImFLjW/ElyDnINZ5z/3DCkpIEBeyWKuVx//a4BjAHonZUroyCIZwQabwWJbzNBSA
K+R7qXjFTSR6r6rqIbK2wrRoMJtwmgdttqJhEB/uWnkesHRoDu2JDwOYypKr8X0r
3JY7AbDrVdRwd3DtoCROUbTi0IbyLl39LEqq7mNmJc8mXjpvaWGPy1uiGamVU/3R
uNB0NXWT8yRqD863aaR2y7ftEGRtmobaS8Ia5TqsPKHVGFAHMZaGCq3oxgsSBJrS
FansbTNW3+S2BSuGIw7xJXgaAOND2cJ/YpiyOVpg7+kERFujySyeYo0NtlK49ZRi
U76txfP/XB5vkCTM3o8xNykxDcnL4odnaEoJwDRPai0JK3rFjKnWVSLSYXF87/xV
uxeB4ac6+Ps/0cFFsZz9wQWtIa+JlxFAsDHyTzKzSsaB/cSvBVjUZEvURvtddtR1
vSlrf9jLZ1lX+RYbASqVgvdvjuweX/7EtQhkT75k9Q4x35KUEftN9YXqED8CFhB0
F6XD/7N+YNnaZTtmn5R5Mmd9s8nVXxNPlHRl5ZrkZr2YfPsaUyzhB3Ntn0o90LBV
WawSprJVTfamjZLfdqRwkdi7nlHFqCjXk9jhTFdoR6UVRSijqKgwOwe1WzMAEPo1
z7YY8SGhtbsqZGWFownordyJNqUmpEBv7vx0VeWl9VZCRCwmRzSg31iHrJV/pZ/a
AnI7F+a4VGKqJMuLMzOGj1nHeWqurvMgfPWs4LosPFm0FB6W6biltbSHsdvokX6E
sPftBnRSCgpJLW0xJdBumstcTBKwsp5Dgo/rWjr4VLrrx38jI57qAwNPun/go+yU
6SfgSL6RWqi/8MWgU+zqLwpwxzLJurVpb4yYLTTTuW2X8k0aLPBbcWNZfRcetBRs
RdmLBJr6oZ40sDpAB3S863IhZ+YMdGhGjaeLW3G79gZ9mVKRdd41M1WY7gGSe7tB
joEpQ05nFwBe3ykq20lNltBlnz3K7DGR36zBRQj3GppiVSJYOnX8gaBLeNPiKYPP
aDyF4MKRqvcbkVXyluR6I3t8e6ixNDGyk415R0yK/7TJDSHLTgfeTFBnJ2umt5iq
mQNzqYOEXfdllIcQERjZygO5rVz9T8IJx4xY5FAptlNgEdMlbIJ29hNpYzJGSBU0
+PBUBLEpehPdccToBngiaW4yhunGApbojfEmG9K7V3HWcb+1ZaGWXwMDQdYeRioJ
sZwl7FKpqmli5XDOvHcuUJTpbIwBMifcTn/LJw5tole90bAHJqA4rHRoGIJHlgBf
GWInnemrU98LTCvYxY1+hl0inSDbvtAsgX/3xqkOeh0p6zQbcSSLaYlwP1RhBKCh
PvuPYNPHCDwOxow2uGMNHLyz2wW23EUfI38kCqT4cd6E98v2Ll+X6REKa1PL+XFz
8OUagWuPw+0x8Pz0R5ymf/ILQ2XsOrgOjTviUINh4CjSN4tJ2QPppao9T98mUxe6
AfD1sKQIz/JG9RT1lCu5TuhZMUhRe5Lcvmd7/vjGd8Ky9d5FdIRAkkbxccYy5pLJ
vr4DcJbVP3/iseyDU5PZfyLdtBz3I4MREhASXnq9TIfnaD/8kj2neBmdSjFO/NDl
8JecR2SmQfxquNfz4x+aixi5hwqPsKks+ZmjG5MU77PM+x7mvZtUObQND5j8o0M+
7T86WT5joyiosF1dtOS95EBnldCTo6CMsHgYXyJ63YRQT3KcxikansEwwlgx43KZ
QNoH2MVNg2d4uFu2lzKq0KT6VTncLzhE0cenq8ifnyvIva26Vd7ZCiPHc/2wUwF8
m97o1pPf5rTLkbwzp9+w4maYYDNz7CDkwadLHkpgzTXtlMS1f9q1mAEs48PuhZ/u
Y5GND9aEhm3jAHJsvd4jB4Llx+jaGl/iBoZgHkgFb2k8AWz3cSdZXXkEn8Iibxob
tM8lEfps55904a1TXKxT8E0iJ2vfUhra7m8rcHCdp2nJTbY2lHFHLn8uaegAMe/2
ZsbTvoj3OleZX+uwSkTqpnig0QPLZi8VFUDU9D0jg51dR68/qdNkL7GBEvtjDD5i
sdekcVK5pKwqQqZrSWl5hKc6ZDv6CinMQuKHnny/uoF2wuhYd6jHhQCdbXNF7oYr
wsKPo1vYApAB2bjTmSOjPQqW8BqbOGbQFDY48tDz06K7WfYHefrj0k4YRFRVZcXl
84QHVJnUbdhXOJ+wKt+k7fq1nWe8YuoA8OEa0YCVbDS/ZDiVfWiZ8Ls9ZBnuxFL1
A9zbY6hStuTMHqcyaCPk4zsZXdpNdL6sIyry8se8F2m6ITrQl2fF65R/lpCLa8T0
vx6sGxKNnZd5pOS3oK4zgM4TVnTXVGp+uIITnh8zTY4uenH0sHBDgv/A5nMUoMvr
8UeSs5LbyvoZoQy+QospJHbv5eJcsltB1Q8OYyStryF/TmCm20dhwChfJizpZxzM
KXW0fb9/8IfuyFl2hi0LS5TkDPa8CT1KkrmmypmmrSZjIZAcX0VMT7wfvQjC+jLU
7+MUTvEw6andSoSScn1huOQCCS+GMbHsfNODnnOq+/KyfA77tD5gRgKX6azq6ccy
cFyoDASV8nBNpTKmUpAO6uY25i+wO5c8uRSbaoJKvtDsa1bIB3agd9WHMyBm+El3
1PfDUBodgTPrS2TX/AzM9SOE/ksf/riGI8K5PRNG/GLkFkBOn5zQn6GkxCEaCAtR
h7Rycrr/YVMl5wUIgVKsSjFFk9qALu6nsaqdEeMilxEAgSS0hA18wMbraxU1W+/k
wdnvsT/DQS2REztioquCx7xDCXpANEY/G+HQWmPswDzeiBOsnLiMRcYLeIAQmk8b
L/W6+r363K7ZC9wKEYGBzWSCUABR/SVoR+68rR6AhBgLj9Uj/eOGns1P7eg6PXp/
QEssmGGqHlEq4xVYoo4ssk5cHLTeyHp4+657BTmUp1JbjvLLLzxYIFnc0KnCyBdA
Xs8csBUGx4if27xOiSO2bm8JzLeyXipbA8TqhVGnSZo7/wLFBWiRveGwwOgq2a1L
JZhzQjjTBmakZhMnkaaxSxexRFCvtAr2kU3mCaBmcagWwI5OqPuy5/UDCPgMYC3X
ceV6AhtfNXrg46Kbsm09jR2a+tj0Kd7PlKnXC1e/HzW5Mf3Qaok1XxLGjWmed3kX
nsS2G/dimpevNSXfWMMakOSaM7Dz4PWJqxP8DXsT3ouvSv24XdLy/RQ3sBKOZmbw
dLWsnXZX/BGAa2RXiH8stprh5psxJXB7iVm+GYqEF+QZeNCI/FmgFOX1bLkS9CmW
JHrbT2aua6ndeu1xgnqc6+YqMykvUJFdF3qnK0klo01lvb87q1dERaD0cemgG7+Y
H/ec3Ak8zzYu6k7XepT6dptcGHTl30xe+qQGvMIyN4+KF/K3iIA7UTI1cJEbgkvo
r128a5bT+fb4xiCnCCM4+5+788mLnk9QSQOWnuUfJF07cBT648/7S5dxsuuJB+Ca
rRACmEnJqUhmGZSceDW8HS2oAV0TfI6nP7feSK/ZM3zNGrMhhJlTD8enEXi5YXg0
WB7Njl94Vdrq7YF4nzhP4+Bq6ofDgHUx5PRHxYnI7xMiWdqzRw0NcaZ0qsvI5Cbq
Tx5Doby6X45VvUBDhHE1EbVQURiXruF8llqVqdSZAZJNjTIzGKT92KRtnKFEqmet
erKzbdABRq4lYFQ1WjdRAApyIZiShVmiT5AWm7ecBeFUWPQKRPeVIQU5Ig2INhxq
bA0b9L8oyign02Eb9IutEc0yptEb5bWDU9Wn14dMjqXZu3qCCeaxlIyY9GoCydTs
VFz/AF62EnPE4GT5qq1FrdzQ3uRSH7o//Iys9zs+iloifILkefmDpwkpPmNjWYvL
QUpowWESfjA2y/nFXhbczapuXmbnihBLHfxiMxc2y5mip1Xw7WehJIUA0VISAnYC
P9aD64wmMxh0/uRegZQ92Ep/ddaam2Ot3ewPPXpZEuje1kJfeAUNP3Na+PrfFKa3
m2piUJ63tbXydlTYxTaMbOYY9SM+CAN6YlRY3SI6ws+AEOkItUU0r7v5vK55v7Yp
MhP/D3J2IBvZA+vci+nfjhkjXqb4j/UtbIMCk/FDORQSAM8+fiAxjpQWK4/mKQ4P
RF/720w84Jej2JNekiFgNhm6tWXfxNnbzY1Jn6b4oopKCLy8+LySOJW34x8yecYp
vFVujw9LOBu5G0VbLBjmd+yHLF3sBY5FNBhmNKG7TZetawI+MflcRHe9Kjq7tC+o
gLGQ+/jFZB+KMSKO/tLy4o60w22QeGWHN2tchqsMfRFGB7C9nWNK9nFvWvIgAhbQ
P5a7h+hw84fkJIKzYLZ5SxEGZobJADy+N9mIVTdf5dtazS5DSx47cMSl5VHUjl4a
1psB8yAq34Z7zq8HQ1R3T/r/2FBpQopfTTcbmknflPDX2aro48U3jObQAuW0A+x1
LFR544/hHIQ9Oktht5QTlAlWQIvGwvI0SMbu4eJaZET1fOBNdt44YXGUiM+OA8Lw
VwV6qPVZP3Hsf9CWM9gcOU8mZ8SH7LgsMLipiiw5vh/zAxEkXRe87XpT53WSjtK2
fhg5OXdcyh3Fwa4IGW4aovSkmpRJMGsxJFrwdRR20QWb5Xfd8RFTWxnQp+ac7Zax
5+l9oXB62O85Z8tEOgnxTcpiQv9/mKAdaInI9gPLG3lh3PP6weXAbUnSzzv3VVTu
E6ngl5kLCdLdQibcjoAM6CXbRyQd8vLB+V3bOqQIbBaKBTKrWhQQAHiVsluZxsZK
/lRO4IuRqNApLvIHc4M+LGQWvlkEAXFsN9IrbnxYxCTK45VKtumf4Jpiivybbwx/
2D15bgxMKsYMU3qflJAivqWVUTvyxVTpsIGNg4BVd6tDkb6kdhenx7Chugxdvfwq
k1lhJLhVRzi3xbo/8mPcOzN1cvf8IhGVw7j7s2/qCLogV4bRxBaYq2+qhVcxCsT2
fpiDVMo3GcrhXwC3MNGNvegE18UdGNoychkcwlKGIKU+8I8gnjJA5eHnp0otSh/T
EXHU3ypllkiRzzRvdFgj7Gbv8wR4dmDRyaUNhvTKQ8jPjTbccZPgtBDhPXVhTZO7
x+tWyKFMPBT1yLxjw62EiB33CyAsD1N+wPcIwyJaQQfXfVc7PDH1PVnP7E+CIFUB
kFRR02+YPZ1PF8cEvP2e3gsgTsawun3a+skaKtCDWcVKcAD5f8tliGFcNI9U/fSt
Byhs0bblF5aJVsjR1PT/jXxhXTmQqs7AFgtMO7XSdM3uLN2gdJ62U11buU31PzC0
tizKdk0w/JjjcNNtMsoSocK08seAAvMYqD3Bpc/liirRlJOJ8BEbCrp052OheKTU
Ot07v8PW+9lflv7WBaP4eDpkMCo9IVfbIFd9DWyGUpJJvxPUxYijxqgrg6nOh7hn
s1GBv19ayzQHefOGtI0//sTjFgUzK1UJwKAl67us8WrT4wxB5+nY06+qXQn/p5MR
zXLtTlLqSNQ19vk4fFS44Vzbj3DKptK8G1sulId+PZ0d1WibxPhL7R1J6dv89cfI
eUGESE0X7tX/5YD8Uj4NwRubD76S7hOXsYaf9M+BT98c8Z60bN8NAlq6TspcDpL9
KaFyoSs7HIdwwmEJsPS27lDzgBfIuVlgjdTvbkV55FY8dph6l+dOT7mFPf3Yf6Lo
ZdlxmmWKQhV8YzcRJqd4VOAlSH4cyb76fxhzDlf6VPQyRkky9Kk4vFv2bte7muR4
1Xoj5yg6OPrlQ5/8AV9bquKVKJu00raP4G0UlAngPojoToCNy4BMHMz4XO59lVqw
D2UixSJ8E1WMZHzFXt84/vEMg527E7gd7GtksB8IbzCNS8IdyCTNEjh523Fp1wpB
bjyW539XxSiS0iXTrIqOK6ZeCLaiX8BztNVPb3ZV7/El/aSuVW+6Ohw6k2pJX9ef
qFWGmrR24q+EafI/p6yDc+QNNpylTeZc7pl1D3WcROXJRIxKg6A4i4HiokQkqQZo
lgCB+/lBW8Vm1ffU0TTZ3Ec/g8PqRhXkm8YMK1iyNY93wHAmjzjU9ZJ5QE5eDPTQ
zIeYS3Zjow0/fnPYIYtAh0qfzzpk+GHEUVJ5JoiqfuZntfsBpfPRmk3aEOEF8wMd
vVyL+pwIVZs5L450lzfxtZQZvTdWiqQwkZMuDu3vhFjd5Gj1xn07gZU/Lk7Aw8FP
6w4cdWjU8el+qUwlF+4oVXTspUvC34G6WIMFeSaLBdhQDnAMoMbIwbSrIqqKpE1a
QmbVOOY/LLCMifrKxFO88Ivc+B63yeICR9q02lFN2fw/IcK0eNcBOsXHjOJATzik
YUoTOdG6jBwzEBIhkXCRz4pwdAMzxfoGJmqI2rFhuDjpHpY2aIM4JlKaf8xBTmwQ
rCIUisq4TGcECj4dqV4B69wL7CxJnOZMazUBSdK2MAjvL5QzQa88VlIicJy+kxji
c9tAD5EkaBOoTJWVV5TWPQWZ0tEtJ2q4kDcaiF5EhGQWca0dDQMN/MJAwDaKbUe3
wpiuXYC5Gf7Y4YWF1lJj9OIBEEbFE0N8ra4wC6Ahwb6TLPOnvM1fiN9dncEjoKPg
zw8P1QeTgilxRTznmo6OZhfwJPC6ZXfgNKe6KR0MnQpvhmO4TNtGu0/e7CnfOWFh
0bv+JOU26rkYEUGCjWAbt0V4hqPK6oTiBX8BDanrn6uFk5jVhc6yAMVGfXiw075H
y7P7Qh8vaS1Ej2hvWp6uGqvgS1BBgBXYCY5yCNAShiqcPrkGUY1VfPD1n7oJ9wx3
gGWgJYwqwjIvu9hzLlYkE1DJmP90QuLSqprgMtbulPjmxhFPUomzD3w47i0fGa5w
Hf+skKfvTL9oNdqt0KWfZ5FIU6XTgRA0BtQryjJ40V9+QOO40RwNrY4ktdH1rtH/
v3Bb83VUZAxl2Ks8te+McczLWReTIAKJy5eIUR0zbheRVnP9amNKM0Y+5eIxW8yY
6BSp8Icwwwm2rsB1zDFAQAnHk7bDFo2SfVlYQAlmt/LBWtjIfNrNgidFMV4isVA1
Xn8ziAMGjl6iaE2Yi9iMOD9PTt5twYIm+KtjjJ79S4wTvBiNt0ygij5AphMWoQJx
4ODp++0Qvcj5Mwft6p03XYGJURH+QA/mFtUyMYVnM8RxT7JZ1SrZaOjEtHae7STA
RT5nClEyQq3JPgKpXW2+AqTZkYHxr8I3UZ3v6QXG+j3sSq1UjvAenV5bRkw/Y99c
EetcBI5iIyOl9hk4sPK9wGe7ryYWIy5O9OCK3WOzunEeawg+fJUVT/oJYwqWnYfb
ajUjwCiGLKwPT4kNrfqCs7OlVov+8F4NsMUW4Klh1OMFI8yFIx4tK1hZC/PRGUlk
lERnBRMF2Ho8i4WHw9dw1vjsuhkpgdgCPJluOfK6sDcBiU99d8WZ4D0KKylLh6db
qcTsEhq9fwwGFKg4OgmfGuLvyp8PY9jCsUpp/4tL1v3Zrw2oFmJ/+KpjBsITEhFW
otOxoJcMhgLMiegaK+hgTZ4/z2ppMdiy89TuNBOIOFA0Zqeuxy3gFlRh6ki7EEOT
wq9n9tnXqHOHJJ2Bl3r+7UMazSiTRVvpD8VY5RPtKH11mse5J9Lw0n91vskaW/+D
vMzuFJTF9GQSiS9Yha64A3jtHcfeTjkMYJOdEw7+Lh8vGAEhz5vJMMXCZmGBWY12
4+PDAHPRVTsknKB93eqUcsjxt7o3AHX2IzETsy63wm6KQy+h7gTCQyhuJDRgJbla
9LoZUeXjRJJe2rUrnSsRHJ5HdOU0a81Zibctxw0Ala434wUnvRjMpOgmbSPTUWnf
r7PSO9wIs3oFlM+QSvBo9wTnln13C1q66v4ces3Sc9HCqMzWlP9/A7zZxBV+ovP6
UOk5kzBimJzCdPEtWhENW2pXqu14mrrWSviRGHbh0DZqAypASnfYi+srPdIx/3fv
KRJ/Sb7545LapBEadtOr6tADi2i9cIh48FfBtCBqWRmmKApLU+gw0NWEDEaIHVG3
UYt80sfTgPPH1gpzkJHjEfFDKmNuH+KlvKI1+yUNbcM7DlVuFZJg4sN7NoRJhHek
0f+jDBisGavxmlFuDldNgfaxTIMG6XZzjamFAuOb1MBEp4rdG3v5Sf0ftHVGRb6Q
36dlBeWfitS5cQg++9Ntki8eN7EfUluat0b6Pa0kUut91FQff9laoy4rAPzs3lrB
jSolr+2Ybc8t+DZYGlkxa/0jn6LJG/eLxu8+urxv11E9an/zXOQzZckA+wZWDOB0
U5G8e/leP3tBLPAoVW6kz1vIN4KxtFc7rQiGfO5LwgHXUEVlk/y9Gtb1S1RJT0fa
PKpIuEAyPZy3egx46d/aTAOjweDR17Spm95TEnPZfCkXRR4m5pAOSsTxmS9GII7M
Z+UVb+6pgZTWx0q8BI0CSDLFkTcldPGlRHqDyyTss+1n+EF1WUrUePCDmVTXMdxJ
2c6YQ0msnHW752DwqxLZA2Zi20gpa+ENTo6zrXaArQ9vZqi++AUGXjj8cldEuUrp
R5iRYgIYEVFncE4yzgYSieC8ANj9CHG+EA54al1mFYrEJOadJkoVy7Dhvf2zyGpr
IUebivDiQx1oNa+tf6ASyj3Y/yIOH9Vis0SPby1jnolm+xh5bRudcvEpYnzt/jju
+epzULpRIlWmGbkAX1HDcCVX34wisT8KqvWppRpvCaRsE1xya1PqwsQhYOtNJoiH
cbMMsmLD1qA5OKhRlJheRWksR1oEunfwEa1Pg52qy+G5bf1pQFWwW8WfTsLkCYRH
tnwN/r4x99RpoH6gH27bOxwO46WfrdGYZkYF17TsynANxRJ1l0dfRqV59OGf44XR
RPVdxQ56i6RkUrFwUy0sHj/r3SOX+hyVPIU3qVC94Ui2kYXbbtS2LMmdC2mdgGCy
oKxEm5tcWLDf8+hayL5rjG9VlGJN0Q4SaFyDNz0BSPF8HsQ2JH9uhTfszwSoTZCP
pztU8Qf33c6MYIBnzNqrzpJvVApkQkVGkfTOdCsmHYJsfUJWm3CXQYJlGxVmISez
drAb+Bl04rhGpaHRNNqFXmFgiIkNigiMSD8c8/F6pR+utPnNRO5bNWysPn3WboW2
3D/XLuj73M8knu+MY/UYTSdWK4pbfZdyRs11IKKk/ClGVBIj0QrZ3XKCg7uFshJ4
aZz6OI0zrIFIUgmeHsesdvcNqlFXuPIuDwZahvX0dJxT0kq7ukcoDQkYTBirv4aW
yxAjp/U/hpOpQNXsgoPD8FNSB4Ef3b5PV1bF631VNpA+3LVha2viSKvsdnPMFdW0
zoM5m7oUq9AmM6i0Yx624tD/rJabrExY+LdREF+aFfZRDEIo+mUnORLumbXp4yW3
VZFhQ6Tkc3poJqAf53vI7Oi0mXX8LBbGxL05LBwivGtgqDd2BzyDvwYM6iae0S/U
STuJv2hkJpdROcvWzGG7ZhJD070bXe0sFQlxQ9OOWLikVTWTBQM4MmB73WaNwkPu
YXpeQQBcn6OzWdpMzGib/YUpeLtk2eFqrOjdZv3v6pIZZb0TR/mJcVJsS9Vr3Y0t
relNItGN94M2h/B8QeZVF6zM+1AxE8+qge3rZU5nxpPHnbDpgY5Df0fbGDKvLq/I
9uK6MWA8dNf19LZJ/mhHI8GSlgDDUFMlQvkUphNMi5CGvem5Nh88ogRyt5s2qW/H
pP8sA/MAEgHUJMhTi6QaULBOPPlynFZyMxWztRXqyzgE9BlGdTht/RxzLk7rvTzc
W/Qi4N9US9CHHD3BDIZeqahoTzJCys4ZgugyMM6GWCWci3U8VRNEv3ZvxxGUaEyP
hNfClpylgwnV3IVK/trXDIk3kzEtDp4IOgM8sPN1/GahriwixZ1CG4TAUcjJeHBP
16eBiMLPuxlWDIiMZ1sZANCECLjeJJOdplMhpuyqFxQHpGJ1YjNq8kkPWAtX5r/Q
Ne99LKZq9b/LnLwaIrOIMPdh87VHbr2t4bhOMSiDoHOng7ekyu0WSsPDl3N54UBm
oUrstAWsuL1BO7OUhnAKgpE3OUOo+T0xuyK9jSDF9Ny2fW52ELlVEDzNNdzTEHfd
Fp2ol3iBZNShh1Upv0MRT7AoLlv+/r33UaH8dtxXdVb6QC4nem0xVWLuc9JqjIkC
QtStQOY7W996zG15/AjNwSn/k+897dhCIWwbtPSzhFmOwOOvPv2HUpgbbBHqy5dF
ycZ2ChNBuH3htL2S6/m+BQbK6tA+tVUqTHegn1i9wPANeR24t8jvklkRjfXXeq7z
WsytTgpIdioMdw6onGyzlD0Fl9b0ZimceixSwlCJmOy1kO+OMyyAQmX8ovkzpjZF
oZMmPv8ipX3zgl8HhbIH3eLyGhh12bvqW1fWhM/gn7tiTXzrIgJzktw2Gle+6UtN
3GBPFXO1BVOh/jfpHVhV4SQEDZMKF4w9NDFH7eZrZHRlzCLgLFnK2CqilN3bahn6
EwRnHfAjAxtHNMgg8npf77dhYsEn1a7ULcIq2AYV17GtpPyqPfSIbCT8PvJBR6Qh
XmD6rRvNY8D04sLphBT2pZRo8ADZghx8AV24tM0uUpDr+7j2yEBLy0w5zqaCnWC+
eSCHBMZUc7T4KTIkl+q6T/iXhw/VSnL9edR39uDe7suj0cizNfS62S1Vp6QMtrsG
XW3zaUODzxyNJSuVMvYbDMotALkWCSRdeRiMNikcMwJ7+1LvPCBKhxPUowAMiVj4
ib3Rqe/Coj0JRU9kJpuTzmQoD3XLEcG+HkT3lMkIc8LVBX/ob6SQWKsvfv0jZlMG
VrNw61ENEWCBc+USVj7KfRgN9qCE8GRjmV/1R+ZEIazmWixlq8US9xmfxVUdyFJB
HcKcOaJEP0F/0s/7q6T7uMzLKe5tFgyaI3mUUt+kvOGLZVV6cNqXhvkGmjZ+F7lc
ULhFYp9IKVdjVfeJ/ezuQ+LqG27TfL4Pk31lbWOebSnsAfJtLASJjQpdHIZuRCoj
RT0sG9PXit/48Pb7Ta8Twszu9zQD3ZB85iecVDLd56Nuvgw8H4dl+tlLFpfmf1T9
adVu9LQHQrMWGQF24bI6/y2B63c6vqkU/6MflTAkXBS3NIyzMxxLJfBYjNDkjta5
LvTtyW9RMhMbVQqxbPsRfGDwWC1T5ZxVR6vaOmH+Uzi59XbN7kvq588V6zV9a/cP
PZ7FX9i2nxukH1XN78FVzVvL2sBoYbvJetx5qUxkkTjWk1A772q+kxuKMpn3MMfB
IHfzcn30frHycb+50Gvy0dXNiBj5rHNlfEqUgtVAjddiZ89nzNl3c/avgx71FnSq
5gDLBkoIg6/HMPXjevWARlxGa6DbyDpvP8+iQvoFptkCaE0R+meLQwrsB3lnf+iL
RmTEt1JJJK5mrbjEbv4hNumGZfsyCbKC8Xt7BmImxGZB1196LzqSczVA0bdWaST0
gr2WJ/WfBKeRakQKcJql812t3hlptyXSbR7ewa/4ltOb0KoDlgB2KzjqCA4C5HG+
8EfeYhS69BBkIP4oxZHX292f9N/O43sB78v26EfG4vrqJ3kV/8/l0p9cHij5sT5q
seKpnCzNrCwgNJStwJOPWycW2Bu1tfJ1N7tWv/GZP4Vjtk6z5AIHzsLTVW0U0+5J
TebDV0ADjatzVIS7AKZIcmmOQk/LQTrbmvj9TXWAZRhRxmY9gNttsns+g+kFwlhp
IozgmjNM+rffJM3FF4Tqr6wgSeeqTzTBxRC2CqFE+F62PV75OE/096LoQWajXViL
6qtXKDnMPL9Z1bIuoQCKt9ZRxKgHEbiOtRGEUAp58s3HrWD6tz3ERwCmhpIUY1Nq
5vK7/gEfjmo5Af2r34zG1p+rlBSsCRAY8ySQTqfNDS4Z/SrMN9pvl0df6a4RUYGT
HujYYRKOXfA7QYN4dHnFFYpYojpWB2wW6kYANUKmbp/ElBI9KMNhrhz9/Pmrc+C/
1V9biekvIEZIhaem1LnnhHXjvEnzSqEZ5BG1/QRdKdXjxDVXdomzNNcj3/U3E8do
7ciiZa+M3ghGZx5183t+7i9fY+bkJ4SrfTIvr4XSdhzcvm+IVDgcWHw2aoREuUrY
ZJXyW/XTd4vs6+X/I/Q2KxZvIimeytWtQqpabbmfnGGWUjujf2OFMoLttM18nLA1
7ml34RfOXQaQIBwKhgw1rbd4TbUE3ChlKUUMuyqmiS9R/C291JQNgZ8PVjygFw9o
9Xj5zQPyB2zuHasWbQAFwP4qpasBwDAibbpZjD25dij/c/cd9Oqowuf3sr/rS9jH
eJ1wth/nvcuKaYrGlsEzpbeCTckAWRe7HpxN7gcK2/0qJ6H4sx51Zb0+nNl6FDxF
SY+riqQyOY4oBupq7rgJOH7pgwZ5ikYyrJu32pwEMAqxdVekgL04BWQ+YABi4xkc
+ZFynbnLloIezdbZ8G1Ifs+jg3lKV6PLf98yAqlr7ZNzm2yKnCou5RTgabwtv6hN
5Dee07Np8C1uWiLkdfPmhJWzVLwZVP9Dg9hrcS+cswCyihLFly8mpT7yaYORGODq
0yC/d/VYTDOmYDtamjZzH+VBda/5mLEHHero+onj2iyEHAiO+MAkD19CV/PGAmzJ
U1K96zknOblodiWHGSy//u/QCaLzDq0vsrKqMe9lEYL9cOTygMEp/MQraxLqX3vE
gyKzzEifAWpdlWtkd2CL1jrJP8BT5W9dUfe2CY10yJY15wINoMpJ92imWCotXENe
VTRFFRyBJk4X5Cqyod72xSgmxAIW9R3B1XQAonCoalj+tGtW0QRU8d656bpfNDMe
m6jcinmmGEY2EQGvBg/Dn47YNAMMm6d5uUzGUjYPzzBE2ObsyL1yzS7+wHH5N3Sj
Ebs9i4ROeST0B/gpvGut2anTKiQh55/f4+D5mQckZmXhu39y+PlOoHcHIisUFdYs
G5gf4p3SM/paif3SwiyYt6BZ/sSj4cimrlqLu1iEZIFMbQFchsOWbgIkFwAqkibO
GnpwUHUki9diFUw9LidaSZJ0KZzrcbHAy6UQnKlOAIGjKAExlcvPFrA+QV/vaGOQ
/zY/LJiZ9x54C1+dGTdTg2iQx6E7KD9mkHn+p0B44mik07HwxoYW8jle0Rqs50Km
n9fOJMY5KiDM6Fu3oVU+UGwYXUhzlLQIyZPGZPtI8JLIqlLUUYVX0MzJrLDcNOtq
NxXLEA42Cc/dKLNuWqL0wbfDJbzwOqDC+0gln6zQfV86wcD+DgXnY9W1lQAxeOyU
Y1YMiOQcPV58hsPIEHQyyR7iv4QjfgAkdZJtfE2x9nTDZnST6wrJZt9WzQeO3KAS
owvNgoZlfWMgtq0yaOe3noihAeqIa5ai9QEzT2IKZjpDx2W0I+rO0OXHjxEk8EjZ
9TFyHi/uqhkEatuFfLAciUBGDz21VbwAHJ2bwUd79ecUyQABP4vepIxRw6gAgEAv
JQ2tiYdlslA0ZsV1ifVnYKWGuPD0M84J1pBDrUSaQRgmE6n4M1/SVNmgrLZnrbLX
RrcutvEsBu9p9OOgvIJWRNXKd/crcHCBPb4maQcmRMd8LczgJ64+VzbEjL1ohix+
g614VSzDxGoWr7D0Ph9WsthhBpki7pyMOYelzlPhYRHnwtpcXb/tb0PLnEGxPVuZ
5kN3h5gRoxmB22GBQZDgNEJ+hZ5JSTJ3ux36Qo55r4Ah3KsS8qhMtURV9di6xpFU
nO2ZNLp/OeUCQLYePd9bgOosL2sJOu8rROqJ6Hj2zzk7GkezWnqS6sUa+jiACgW4
JyFX4UHCdIKxBEjwnVmuEhKhp4ZJswH7cBmCCt7an8ziZeF1/5z5BIv5zSnKTDCt
XisH2rZFPPG6/GfSYVEiN08iKi1+BNkaSMDSLNrSxdAH6iS9Olj06niQuF08Zx5a
MLAybED0wHqpspgZtTZtzBbcDtYPiFgrw9/O4fCcW4KwRn9Dg2dOx0OJTwUtrVJL
yfS9HsixBjoDidd6hN8pCjU+kuXB77SXB7VsTzpG1yA1uzThNi/loGk/E6Yc3spN
xTXH2NwUHEjFIo473xPA/KBjbhRfDBL3ja9z3MyEWiPuIZhIv5EaBfBWZdxNv21O
6xX0O013ZuOH2NuEDJ5LDmxLB8p/AnnEVg20/ORfQaFPmkX0QO59/hX3TP+A3VE+
KtxhLLNYCOc3ufIN7iUAsyHq6fcmY2ROXUCit8eKrDLxaem59gY2RRFrADpmIyxl
3bpI7bMe/jig+VE92sEHuGakS2vg0F8B2TSaPjhlJR0pFEhQzHq+znrS6LmMfvmc
UTOpaAheYxQ2tNiqo+ZIHe4IxN9qUYeJnvoqh4a2LhmYKVeHKi33QJQxzkZ7Ujce
Pp4ZlY2/PwonQ/DKX/Vpsxdh21cCBmt9jz+8CdyWjTlIWv8X62KrXUt9SkUNkbhL
i6rW0wi0qzSsKTMjMv8V1Y8ArkmffXbFyA4ekt5mG0rBVVZb/1+ChqNXmBYtDYsO
J4s0of62i0WFuMYZU9jXJbuGpAQ3Vh8dB32wpBeSuJoS6UhuHr+XFZicj2WBvoTA
aJTQFpmxd1dmu+U18iIFh6ByWS8q0sd53SwfFo5OqhJFByu6gCNy93d2HHsm52uJ
fIwlif9twpK31A3WThFxx5GoZ2aYdpkYK43rrwcQipwCiIrgoyjPWRg+sUn+km58
v1/f/0YUNFlGGA3ZD83Uk6eoqPM/9mO2E/ExD6acoaQ3NVOY8z3Pcm9O7UC8CmJk
bKks9rmoFliyIOYt5IPHZYic4GynvukrG6wz+dcVjZGSBGbR4UZQIlE0pbuAAYPf
1ooVJg5sweDTnF2cjdExFET+p1PCtLaN8sLj54xc9t//kXpTHwwquFQSxPec0x5y
qflmeWL1qPtZ1XlgzmPDPJmCYi96WQFFnBDq8b3MP4ntW2JlEBSYe7Wu9vLqqZEe
xerWoM1Gp5z1VgQI9yfWdIR584hO22RIaASWhcJQJa3rc6SJo7ADJ9Px+WOw1EZ8
e03TgtVYTay57RiTK5E0J7RZ2YO6JhONQ4bd6RRBtFbuD2/yt20tXmHuge6AysyA
HXvkLRnkAQDaGn6e40xvOCwDUjJ078qT6fquNse+lYVjr7oLHVkUZaDTFE94SM80
xSDCSEWQxYUlQrDddy3eDn08YMKDg/q8rALDPQR4/+958DCmezpwEIDzwq1jdZxH
x195NsBaktltUXApBKiCiDngpg4CawaZM/WYCGVtbHZu50W7mfbiEx/NPMKqza69
soUDCaEd3a9/y3Yi6URFjClWnMROODlNWSSu3Ogv1aQg/0wiOHUL/gjbQLbI7AYw
E49bXeDddfrpJAe6BFWenWHxueNbCyPJMJxpo+vrzxsBiudItcQdjDezuAmnNicE
c8PvV0KqnlDlDymNFnUINaqv3Flka2YxUn69NLTHT/gbmbYRDCT0T5obp1/b9ACE
1TKfc6RROAdr5snflj/ahzsgWtCtp3n9bdSXfVD1wrvl9TCKICHwr/8HnPFk6Mm2
t8z5nOpDQnCKZXbRAaGOGUzFQc3NJ6mIPleTrcR1akBH3VpBBeaa2/+tj9rlUg29
0CExQfBvo7+IiTfZuBlwwi/nDDpH/oKXs4Ih+p7hFHuFt7oym9CF9qUMQUKCaiij
2B92Tx0Bi0BCkU5mPxcY0ilayiTccoYiyv9SyVZe+CuvQp5zJpRsiZkOcpuzUBpi
iWnvwXOjri3VIPPNLHmIMy1e+gWrWMZi8cmjTfy8sXc0PFf1NQMZMMopoxbrmUm6
onwQ9TDF/pZjQaCpebs/OxMqk1pODH2IMN3mS4rbovCtrvehZy1fvI9F7pwLmvpR
4rV3HDyA7X/aPvwngpzbyo+oTjksFtH0RSUwmwLAUXrD4+YktLiC6WEUq11hii5k
bUt/z5DJQSknx1LZzyNo+JypcMsp/kEyH3lNm8HTw+uPOLVkh99juUqLtMXoIpIp
Hxiv2V+Rqw7uKoNY/1oyQHMTsllPJXEhTikRtClDBTx6mKU4hpm3R/ca8xoyK7uE
vW6DMhK15X9RWVTJyr8tKoRR6RB9lAvQSsMj0rcoViv6ZJmvaEDUp63FTedjXZ4E
kU/45E9qQcD5obuuBsKHbwfvVh5v8tEWPLHD1d5YKSBtKfv3Hf7BBpo4BlFnPUmY
e4e4Z27MG9omSDIGR1v17RjA545tQUruYiP28XRck2rTvGEaAigyykntHPMg0cnE
kgr8gTh4GIJolERoP+vM5mR3pvma7/eCzDAldkjb4GD1gvjkhEcfeZBWmXkJ4HPT
foZa95Iov23UKmttuVKPO7T9XXfP5geseZ/dVIS0CuzzcYgXc/rNZRUgYG50bgbD
tlbcMNkhJll9I8QznSAXbiqRH4pu4Yjm3GKHnmxLgRFkkPXVYCcGKE0v4XFMvXts
atGHNG+TbGbYvFXoL0WnLrqbaQEJS7NY6W9UTo8lrsXRwC8yv93jBfz+TDC+9gvi
h5SIacQ8HuxyZjs07zjeQ6Sfo6upZZkqyJ2/GjIih1YoO93NrT6buijYVfa0amq7
nQAOrTAe5zLdyFGNLaZeAUDN9ZceiHlSZABQ1FVYyM3DAet0hTtZPKBMHv3fk11p
/k9K4ug0GCDJklSntayQS7GdILSFuGKHx9OdoQ3j07RxPWxPYIhxId88rAxfhYG4
P3J8TtrPo2AEomp3XyxPqnlgGdUuwzHj4Er+rLwX25gwDeZpQ34kBbgzaL8XAK7h
F2mpTWC1me07ygblbTfVCX75IdzZKOIZyjsDWKcnwXrV9OXKgi7ez3ysEidXFAOe
ffOtpCmaHM+DbdYYC1xNPBfO/173NOpNLzVTYTVbsSxSVglKEslkl141oXX0qMZT
JWRcIqXzqOCBubGS0bKP0iJdbjiZSEEF+Wneua4Ap1thnlbJ6Cxipl58yX5YHoug
ghFMANm1/dKjpOG3i1asWdmJdeW/+3E9kaDN03jHjl5aqRIgUqAnOY7d3XFEVMq5
S99dKecKfKj68kKnZWIQVh8Y6VE+R1MCdU5Z9hzXtVzgsrPmjc7JUQm2+N4C3D97
DkUwdEm9IM6ru02d7bRzQa6v7Vsh+wsw0bisVGIeums8kerV+Zx9i/KsxbPdGVyy
vzFPktGyEP7iWdwGcF1tHTNg20ixpWD2p+uL9W4yAnai+RIpzQIyb1v8X2oK64DX
4yr3SECaOzwADyyWMaxcIH4c+rgdJh4x3Gv1XJ5DV8/3hcWMOff5Ta+cSdzC9gYO
E273y55H0vvaDMtS0DPNQ6pRGigYvdvfMWwW7ySsQ/syaEpr2kTMjzaJTHCdIFSw
RGoJ7ALuSSp6/wvpPM5+JoUBW1n8nqqjnDxqCTGXMOhsbXRXvaDZFj9aR2wRdVPQ
3J5srNiaVj/begDc5Bo9OMS5/6Ihh/BFBE8PMune1rcaJpAE/3znFb+LLEw1DMLb
bMU8ydL/mi/sxJC7OT3cqY3TSf8WxVablq8C7xJP6212hkHtLDXuihBoJYNjDb21
OzW+g3WfEjlakju5ygxCtUV8hTxc4oFEjFfd5hUzs6edenB/yCF+KgkddDsMFkHv
M/ga6ANwHIyHt07YEYhOeq3VKHL5R5Mlm8EGzQ6ZXauYHaFwyh0/ksl1HxsIeEsL
lh240HG3Gjt2/CvZb8bVtcMYm9A84oP3Z9ABD+7gLbsxsU+u2VWkCRRZvG9+9dDN
5rFt4uBk0a7Dr25Q6XRObHFUEeBcbcEZ+cAlYc7/TaqbJzAbsfsQgM+gin4MX3CQ
qUTWnGBdGGoGvplPnXthdjfvFDgYDzlEP50VuAY8F114l6i0gtblZvHb7lHi0UK/
hBx0iAGhEAJUsSMD5/526ljgyaZNBZNb5bpzmjweCnhYagIiouSRKgntKFiajrRd
5ZAIzpfXbKaJrUxOumkOXr1mT2Gjpywo5M5KuI2m3yn9eGvteocYFXBHMwwgPxuo
dR+ZwBALsu3U8FP6I5fzWEei8CvR6Ay0+TmmsuNUa4ddQ/CZ2GJ2hrbq5Pk5eTpN
57X/beD9jfjjKDNfvbAwE4e3fG5vklZOCxGjFKz9cLcdTY+hogYRwczQ2xrUzsbi
m6JYrDIylmxFUpgfNA18wNFL/nhp4Bkb0yoZFBSXtDA2LJZGpM6M7WFmbrMngcOh
sBjvb3squG8mauRWQepgHmQ5micx1TpRfSbtN92tMGKOV8bKdx9RSGIeuw2MQFf6
Zv2av4XjHRApCX0FhH1vY16CBLV8+XVoRBOc96itDM52nsAh6E/aIwX63dxYvdrd
Kzft917w+Vkna2L5xJ8ny6aq6a9+25Jg/TSWHwXOlYiGsmOZCVI2HdeHr0ozH/mc
+tw2XZOCy7L0ZjiSiPjdAvEGUAp52k8xeDB8GtlZaLrxHum7O68deYtU5Y7gCw2t
K+DPOkfVnGdH3xVm7bmLS6+PJJ/W0pO6Q1xKDu6UB13M2c+yq/gXilrGiiVTSBvr
RBhe9lbFHj1cT+O/K7+OuB+aBez+Xf29pXhNi88Fli0nBsHP8aFnVgnbAQYnPhEl
+FiJ5kEnvUb/oCaYRu/yOSZUib1HDqkzPEkdGQK/BOIp5/oRqirC10jlFT45hN1O
1bf+BPP/n6VrNxqI8w/f6bdJ4pCQp3mWWq/OTT826ioCUryOF4aMcbXLWjTEZVge
4sBhS2zwXcTdNfxU6FUOPK0WuTJI/tQ4tupENnBS8dmxOu9SMa7mQpzR4tpRtzak
2sPVP4lDV3pv5e52I9Nzs2+OILXRArWFwFIV8DllIZLethUFACMxhnE8WPcABrBz
rnZFToTRSuvFBeNw5sTmJcX7Iq/InzqaV+CUgPD1Ere3jnFLYTUuF/ok/wBUyneR
hGlZVnYn3dk8F5NeD06jwPf4AAY467hmDMLgexEDyEa1c6RvassUIu9tOByvI48d
Xy4qOEX/KH39XAhlAo9nbKq3N8Y1Ji2mbHSvJBkUWTx5py8ojgfH7wf9+zj+OG6I
vnLSGrQ5P7b9nnY3KZMfQ4dtC99SVoyzeLRczJngmocJJe+4pzkyuISqkY9y0BfR
RO1DJSSuls+esEnAlO4UZYKIHIvFHQGpnKrg+n7UwwzukZppkSB+k80S63vDTQXh
jCMA0JQa01dyka20MHKMVfUcVHWzTX7LfRY36kKERRmXRY0rEeR1nfOwG1cv9L/4
b91vwfLArWEu8x6jRMPNMXnmWaSz3vNfbYVJZAF7k+MaGkelKXLl9ILOhZ13c6Pe
KBGSr1IF7iVdXZIYB8eRQj70mSw8x4+z8M6/XkjWerIgbhLosHz7NzpysDApqsgP
dEHa20acqp+MM9M+cASFdYI4lgca4B3K86HQDJDNTQCmj/WwoQP9Q4TEqbr9/61k
jZbYcH9KHh3lG9QZ/PxmnQqopySgIYlJUqOSbluFpKNYJeGT4sJEpYCdPBNKkYIF
g2BSyW9x3RDTEI2Um0fI0vdb83Vkc9BgxdMUf28xp+ZXGoll8z++HoHwFE7n52D2
naZ75E3zAiw05maW/hWi9PnmHIwv88rDMxnv2zw959Vk8kl+/MESSmW8wuE3UAJT
8k+qd4igl8oP7hMjNzuVbr4xmnASUX8AB2q7noibgV4TINw3YmOGuc23H4/P2toh
+vDepwLXlx7jVnFQktJK/2l9Et3nQcohf0teOceY6PbULk2xytgXqGTc1REISYYr
3BwDb1A92HmjvtCL9IK7B9jDnZ8LFJ4rte6/Jvkz5uo6JDETsNYTbbWcYKKOpS5U
r8LiM28TR5Uuo2rfh1y3+wQICAsj2IC5kO1cLvQgy/bSU7BmCSxbi1J1TSqN/0do
zfucbz8W6+0OG5j2Zgd2Dyv6J/v3EiTTbSMs1j8H0FFjlOM4hnXSRIhzXNR7ZIts
a74pFZASEesrpxceeCCa4hUn3UebeaF8LnnMMJfLAiEV/1czhVNkPhUTT+7tICoR
SxcD+9m+NBqbDH9mgaZRNHhD+keFYZsvqNkW3BNlaylB/NHJG3PQBo0RDXUdfwsT
H31k1pdKdDUSg60DJV+4Cyv1VV22Xr5dnj/gBRn7xq69rbzHgqh+ST3Bi6UFgixb
wc1ArNypHjPSXvjPk7z9bT/1XvzI9Ij6ESNW/Ax5z524Tl78d5rBApkuX4XdOTJO
zE0hqkr1++VWR27NudccY1zXN4EgY6wbTxswCMeXLmgFnHyVXPlaHlHX4a7VMH8K
ydtLAOsvlaY9nNdsVCDWUm5ncn4LeDlk9vWrx9n6dl7W9YmfoT4nJjEWl45PSkSD
ygEXlRLZ2qOfmcB48Km3qw22QkPRatbluuC+a8sZOd4ltzH2k4vvbA0xm349vUbI
PMZZl3f3rTpEIHe8L2X6lz/noie9czKaKgleDGH6JQxnCJmxVDY4GvZfP9pr+KeS
HmTM4h501tAdxvAXFzyxW+uJKDBSf5TPQFk4OTgaBGTiIILvzI01rQir9AeqeCZU
TphRXVTLHVLVVEqA5TpmGJTDkfhpuluj18tBh2dETI8YUXehga9Oj0yCXpti4SjQ
6rEVBFVFE9T726YRtnA/OirOs3pII8et15Zpj5t8BcTBSj4gm93scu9ycCbTTtpE
t5GOlibftjcoIlq+UIL98J2d52OQ6/RoYLmVmScRxMFsoMYOT6PAIS/NLUH5/dhx
a6wzty8usXy2srtXqsqoymuzj5Cw2HKd33vMjO0NBmzO+jHof6KBxQBu83Hd/eqI
g1k4fiVu7YZl8GQ1mTt8KH9LCmmMQ0H8BkFJ0VNXwnECSI09QgZypzLR3m8875uP
9GHm9eCrK72TYxvXdQ/rs31/kDj6pujrVf3V4Ra1Vy5KFI0oa3JhaLplfAxqjs8T
1CoKc1v0Tyv5WHOmkdqlf/KFvGsmFzyKcU8L/SGSPvAGYMjGmVS5zUZki7QKwSEi
SZ8rN01+3UQ9EvUYUw+Vr6Kd1msOj+teAZY3V7IMkC9n32k/itO0QZa5k0Tb8kiS
1qJdql9hgSb4Ugco9XnHYyfuUQ/Btcj43qvcI49Sa85p6xpoRln2j2m/8VT23rzm
M6diWK1c+kU57JRwmXOYNwnukCuckQWXXPAl4UvRXtCF0kr6umoBpHRqngZR3dRx
J0GBwekCsVgouH8sp0fedKidMhqtPN7lw7dkEemsamNZgD/+KLV67g8aqAqWfzdC
BpDjzY2jF+PiPvXzKCnCdj+pVL/ZxhMMZlAK7TXv0FBgZszqWkaYYLokGWQ/Mt+m
FuQExZiidYAuBnfyebe5wMe6KXxT1VqpCu1rYTTErHQmvRSt5asUr3jHIVDBzNgW
mezwcWDjASII+FXCtjggnc9Q31fyO8z+Xhv522ZShg3z7aUf1WxFrr9t7/74sFkp
NhScGqMoIzsYEZiZ0UJKXzl3M/RKuHjGQ+NoJ/vc38YDY8+HGG9sCAR6N3miehNc
o4o37bJ/LjueI1qrThr2iXKGJMXRo4UnYP1f56zI6dI+A1IIjZmP2NlN+xDT//kO
GijtV8icgToGNx54CIpbxMqli3iEWgcnl2deknqBxpU3iIrbKvPyAd1Z3dLkhGJa
mM2EY60pNo0m5L5l7Gn6TpmO6tCHIUDtQz8Jv2jApQcQFC8kaT/dfoATA/tyzkMY
hcFs+KMF90rD2XA0DVBks07HNuMx8W8534ewqeZP1eC9C6LtuXET2qU1BpSThjqp
F47+t8CFznRaJpM6guZgE77gkEklwvPrzQFwNXCXQc1BWuvSPj3bSI/ZW1D9o0XG
XdYdJd7q1C5fqc6A+SMdeHk7xR1WV2hqOVuqRmzd80bJGsiBDSO9utuetUcFQDkK
TUOndDXvncMcf+Oq3mtBGSO9tjERZd+MmbVur0UhaBVMuuLTnjM70OfSO4TByQwo
tDaxaxgDnkW0VDxebs5005cItJ1VTCnxkHlxRphJ3JMgAi8KR06jp8mjOW4tlgZp
hR/hOhZWFBXYySao9xVoSV7/iJG9UaLETTtXviJH17eCziKaHxfobMLpXOs+CESW
bgLFr/4orA2x3UeSr5zddkfRX2u5dPRbcbbdwh8ggJz5O+5ZW0VlqvlsLswee26a
Ok+79TI5EoJ1ytMZ69tKttwBu66+/mcVqQq/56JsYM7rz/osdRuL98VCOqdK+X4l
S60UI6d21Qh2DFrYkuGG0WTZxdHt6aLoeMSxmOZcP1FpijWpBysLZDIPC1ZZNReq
ZWHtFd3Q/5zTvzs5lLrsnHXRzrUacohKx/udum37vGSK807gLdFznoj7Ielp9BNb
vtlrPwE+59toF+I5M1mpJQyL2P0Lkp8IQds4Z6/sBwWBTE7ABb/AfyN76UxOiNUP
DcgheYvPeszSBG1RLI+s4y1MU+hjvtp3/TDwJZwFxtgkWIPV9taj4s6aohZiqflG
lJ0qVEQPMelXoNzou4wVV/8oyFDACCd0aa1ougAgD5Q1EGmPYWmAWKy6wwKtg/R+
cM1G5gK6KkFiZx7Cs+y4uvW84/9g6lKV6PmVAbxkAuRoPw03fwWkAvMAObM6k2z2
aMf392ql/XSVHLgoDMqgfDorLSZM3xNKDMd6HE6hnQec/SmPjQgtnDUpZio2CA/t
Bcb3KbcL1Qwm8L1u53oFQYwyXx3FXUGBEuaQ+0QBWOUY3mYsSyAvV/OsHha1XWfa
CiuZvMUDTiGtPo0GWjqu+Z3kxDWrcnFNenuS06Uy/tR4fpFr5XLdBLuzd8V4uLg8
XyYwkTciGmmngJodLzBpmcm0WVuGTLrVEEGoBsmRQyAAACNghjArqc3DCvqvznAY
dn/aJ03kkm0OC3ngrcM7ofRtPoUvRHXt7tjt8YCLnI9JPZjaALBWRExB9Lrlytoy
3Rwy8BckloFwScsH9M5QjTSqTAiNRY0PXwuWWOyo4dWoKWDOhwX1AHmS/7MJJ0FT
srO7KYgsexBa6RpgisdzCx0xwgqxg1b/9tJcYrF4C9dUza8XZHd0lq3L3NePcna7
I5YXdyDvymblhnCXk4XS7Tk5cmRUvxWq7TckMxHjNPKoEX7kZ5qd8KQL22stGgx1
Put1E+yYKhteciyJpvyC5+Gan/iyNvQUhEY6TqNfSgpGrIXou1I2KND8PqyukJnl
XBMEWPdf0veH8ZAs7Lxe5KdKxd4so0Db0zIOtyiZJ3bir2rwJKErN6lSnFh+m8Io
zfO7cMJqKXwbGF6BV4eWXOHV0npJkmdM9l8j9lyOOL8ZB6EZBGoyh3k4w00xBIN6
4B3HFM9bCP3hkFsZ/LTFSkpLEG2vVIloaLIQQuIOPuzurb+DrWBpcP6zjf91lr/I
FFDToNQJCfr/VGbDHZngRmO93nEs16iyNJ7jz1SCPLz0yE0V0Yphnvz4bN2Nbs/H
RbYM/j1qS60HRUQlpsNYolryBJ4P15TWC/KtGJh7bJXf1/Wx3ILFUkNqN5r1Sp8I
eGUz1e5DLJDE+u/S+djFXVM7Tm0wsuJ/JCqnbjmY0yXaO1iBIiYlfAu50DaQksmS
Qnf2CSaMzozbg7jDNTiLk9yrh8ZQIs3rsW3MEKrkBss3QlA56O9kke+cf/YFcXep
6tfk+iNsEO7pRfYuTRSTwmlku6H7e20vLNBl2LetYU2GV6uhnCGDiDrW3BUSWZtu
igcgGMG17mGft67OXcR0CstyGSHZ5dYXzG8e4jfB3pjqttBv/VQw71bd/XWW4AHX
H86sNF67KQgFfRUsc+wzwO5ZxIE+AXE3ZmjPu1u13nSofea9C6wHYbx9tNha8HnI
dlOuP6zw77zTOWxhyNdk2K3XFct6B4We5HjvvRfbBbGn90MeGWxsVw+X+LQwCh9X
T5QKm7vh6IjxXvF2aPiWuWNlrXH5EH1mQiv8xJQZxmzz/LeiZiNo+z0hxlzBt90+
lEB4FX18gBHKGB21MriZkSjchCewX04eJCR0+TJ170WFLiZfs4w9KZQmnYZPZNS/
7G196fzOwNWtlM8gtKOiQxRoIKMTFmH0DCoUliauQgX5hHj4nwKiAOAmbB3zhGam
9w52HKZRyw7a7w26OJF6O9BwwwEeqIJFD/7UTat7HlNUulNiDWy2xYoQABTP/rkq
l4mzeMG/NnkHRK0daQeRntcngMODacVX+95u/KLN+2Fsj5oASQu9SEcz4bf1r+71
dQAg5Y5odC1kHoL0zq6vM1pblyAX3RUQc9OFzTCLRMV6En5gV508h7KBN86hSA+P
2GiqUvGyg51vmmqVFFfVGmACnAbfPjSAyzkTwsF9atvAQkPWjpQ+ZoWdJg1NthP9
DgAlOx0JYk6cEeKRM+md+Kmic7D2ng0mbvR1BjqkB6sfmkPS2SiD2NQ9mD8JAps8
FraBZPDkG8P0HARclIoiBRDWO9D4FIkwoKGJr56CtpYy602Dfyp8iiBxC75ekWU+
XEhCjiR1Fvvycz8xuP5hoVG4+aNSrJU188OGyLzAeGiIZ2wyiBtqiOCVHoOt36hD
Q/6v2aAwICDg3bAQIz5i5knxf8UfX7IYN1bMdTwvIbQA1Y8QEUDA822UuERKKttk
3zo9aQWsinYOg0PDg+sCPZcHCQp5y/j1iU2HfBYYQYjq0Yp0MlD79MsWXmJzOTi4
ip2fu4ZpUyqP663BP+wdPTQhDmBJuxk4urSzfkTSqYXdCIeC230j6GgoCZsyf0Xp
KoP+ZfPx95ZVsCmue+sdp6DLexxGruFfW3Ke5c+C8FlfRsHD5+GiGUt0CNKuSDnv
xDjr+52Rl08oJXG8ayz1X27xD0R4cbBgxqA6LU1KcGkW7Uwlj6u/8Ifp07fGXd/I
t19I516pnC+k+BwsDmYA4qFfD/pcp8EThDN8cFRptyfDMQEWtUfSijGJPN2GHu4/
QjlswNT+cdeiJkrkksO9mLeCG5WR3+gmyyffy2s4vWZxwQCV7J4KDPdb8LY4+SDZ
FYrUL2VlvLsjnsHfPCkiSz2o+P/j6N3njVXZozAZ+rRDH6Jpf3jHrh0wBCKmPb6k
fiGrmIr6mAjsO/Np16TpQjezOHzyW5VYBZBHYso7x+DDno+torGJqeZ/xJ5ccOYy
GQHoaJY9k5YscteBQK0liDCFjccq4KKUO3uWtobfqSgS7jwTUwYKYLrXedu7oWAg
pc/xF4qYs6CdYktaYDbsRZaZSDB+Pzsw1u/vRWuJLqQ1ZFVatF804VuqG8bwK9i0
XMsNfx8yw7n0jgM2Mo8Rjt2w70726FR1twUxZ67QUqqBy9z+5K1udzAmmrqX8QkG
RhWo+mQ9ZeQd/WpjTlNknLfoAs75WKy/PhP4aoyTqAxDPeNKuLeI1rzNhyQJVRRE
Wf0Oq+3SDSu9VkjOydLZT/gJMOEmTbx+PlUhpKMBMGA20FliNv2VuHn3sy9Qstt+
9fGU+G0evsQHUa7iIu4DfB+fSByQWXGM+t85IUwHE3jdzD3sySYqhJ4MfwR9AhPX
0Xsp6SbNGL4/Mz7Nyi9VT7zuKailAwpJ5ri8SsrLPL4FHxGLprtiPBmr9/4mwETp
9Bt/LoKusdAs+VIIK/2HM8Qzs1cPXrp89NJx/nJ4SfxAxy9BFXR0Ja/rzv567qnN
9jNiCUhWcFXM07+wrACcn7yxd6pzwYurSSqP3l/eEWOsdRdLFrZVvA989AJz7QdB
qjCWVZc/5wORBinfV+Q5qbI0Ix2FLvU2Jc0AG0jl7Wsh7a0S77HjlVLHNn2IuR0A
Y06Mj7UDgCrhHVyF6WbVCxHiPqFYA+1gtuMmhFw9ak9mTa25hndfNcKQnlr5hyXi
5McUEucPm19OrYtNijB/IWrwfcyWbG6kEg0sl9iJ98S71NRO/iv3txytxq+ZsXUK
gX8bWzcH+abHU2JRS6uI1/jHpPWjrzOp/EU2dTQm58cLmvEWFMDAwRFGfrb3sl44
aKGPSI+u7uEyzeKo0mU7zQ1PKuIwSSjJtbS9tGALf+L4X5ZmTIeN5rqNTbex0YrE
h1mcqhELGPLcf2Gm26ByDF35eNouxs9mfj9Sw9SgT4d2kIw6pXjJnS8UdQzxMs5C
AaQ4u2BRBmgzhRoBF+TUTLeYLPcXxpmuak3mWXSxOk3DtT0xTYuNLJVm405AdsZB
LtGkkCROeFwOHBVqZu1o2c1AyIMMc1hltJoLrecmvq/S27AHYc2e2xlu6U4TM2Of
eBqgNozjlBg18WrYv8eeLxLuIau3FxvDoj7+A46x5dgMyKjNWDWgfTerfthmBCAK
xVS2k09ol3wDApaAY9cVHpAfc8a6+xyAam4+wBynl0uOKh28XR8CiAX/VJNHiRDV
270QY5mKUR4vhRIOKa4i3KhirO1plY0UJuWwulqO+E7IHkM19YQPiXLeW9PlO/Ad
I1a97eQ1dF7Chr1aT3jQ7g+pF+z9yGeY6hQWFdHmk8Rsgl2VYTU4Iv/YFZn9r8/L
jhJlXGczpoUtwFvqAG7m+rZOF4uqKI+w5xnuaXSvY8fXkZoPpMVeW4s5WP2L5DwM
tyPkQy7Vu0zUU6IigwPn52ECj4xRvOJvS/busOKVShOQbcR7zE3TK6NXQ357VqHE
g4UMBd11ZY39NBeX6O6B7pncAtmERIQOvKhVGupL0i3RaconDRbXWV2tJtL7KfKZ
8XKNCofv6KBi68tkhP+4qCsG+bPBi5VGqdCdE++mP/BgiZ+nIWs28LIhT+UcnkAa
s2bXeut3YAXBTRtGHj0Ds+FNGnmAZYOL5yFSfw4SpBcyMxG3227rG9c9rEmoSbsI
sIvQy1d17Vepv799JyMzz4ov59geUdDsOFe908eYPFppbifR2p2SmgPi9+cCkYVL
342nZfasLAD+vY/keW19heiLUSLGgoTBM9RKiX4hKJpVTY6NrHZWV03kHJ5lE29i
X3GCL2WTK/ipzoXpRwqgbFZ7Ekl8JtV5OFZPHvXmDRbZDscKP60dRHUvwrGLubNC
eYHMOJ+dX6RnOjE5IEc8IYbVDCKfnrEoeW/aOiJJWpGkHqho6+Tg0jVrAvYasH0b
46jbCVg7IMUk1bToVamb14B7wnFmLrYCsj1IG4mpvd0zCUcUElDvqC53ag/kXCNV
TCiMgX3LpyyHVER41J5AVvVIk83yQLxdDN6ESCUGmhycjiFYrJMJydOpsGvn0whg
v8LAyIUZ9AUMPlmPVFrtrPd+Tt3qWaRkzD5iizxVW1hVlhIViqLJS3OTQ/c1+qgL
PlJ6O1/dPnTH0yW5vj0oB4W7CQbi9WrJOwUW1K/mvwFUt+8w8pMYLY9x717IC0AM
SyS5qI3neQqJJ+Wce/qampkhRFSYuDlnx2ngYUhhyxDZVD4SO4P4WZHrlwJiZU80
NYclQOjVtVbWkm/tXJcPregZfOYDpfstTrupVfTr51moglyq3iNFUJTjcrocn55s
FzZaiA/s6On3KGvmwbdCu+6xamn/AyvDkGRBV8oT9K4aE+tD5fbfuZdjWiSYYaOH
M9Vx2Ey8fqqz103MC2SsU3Ds34iKHXuNi8cHYx9oQ0Zz2SIYRYCbt8yWUPApWYk4
UPM3lxNYW5ZES335/cq0NHiVlwpry0hPhAkTAOdZDbdwgnctuW2Hx53I/KgqDSg1
JVJ06E/866iJ13lNSZ1z5eWoag6jRbRl3WNHrWjPEtHTwRucHpjxcSjEB00eHZbB
+/J2cuWyuwoYkIVePv3s2XRiImPKpTE2M8p3glUvz6A1YkiYaSY8nFVwqL4a6VqC
0FqRJF63ECGcpxVMHSGRzpey4xTowZZ6VIpc8gYyLR7b31R9NCPi27Mx3p3NR68N
f+BbNp0v/h6pTYaCYk3YQXcg8W9bh04P3CQVRveZ1rYBOeQYztL+ph3yrhgsh+YX
ED0zLcJplA74skfMEf0VV4psJkdubrhdpuurzppZ58bkK95z6la64mvb9oLC3dq/
t/YKYu/tQByJ55pEQu7MV90aEZtqNQ8NO+3IuFhTQ06qLjnIcW653s37oLqLizbH
NCdrDGWbGmK0pjwzSCJMGPhp+MrQ0xHeEg+UZUFtw8WFwyjYankrpS47kdYXaoyN
BgXEb08V1/vQjytRcOOaqSRth/v8Lwff/0tWrlmfdvLvcJAj1oLOjw/yWWn71FZ3
HQFYraZBKKXJi1dL35j0fY8rqSFFmKj0Azs93ssGyXY7aNfiXn1FN9C2fDVWjsze
wGpvniaN1EnahUsOgYEK9rHz9qbKOb1OLoUawAPXUBBN1xnfyyRo9xRNkrYctsHo
rff2qqqHvoNR6WPSW8FNhJs7YEH3JypQ/GU4t/er2zOrtt5I2ynqcibTBYhzTzJj
9aqZCeJtzHHXYAuHg6jiHXovRBO5PcCbEUuziZvTfPjdgDkCbgJ2fB2op5JVpc1J
SgSlOk91ohEoG0zy1JAgbTgGBJGa2pFQFe5OGHbB36W8u9mSI0wwO9iPtlfRzQo3
PIDftbJourrpNFJ171oxe7v6Zv+sOzt784X9l25rVpBIQFd6wU7MWTlaYRkbMLfs
YbXB8LGpR2Mc2rS5f0aK68rhOP/hRRnDeh8nmD8wKdQneUOMgg9BHgwa9j5yeLfH
gmeAcDVqoWwH9RGKM04TVlv9U+EWa7WuaZOg2uhxT5E87O7GTSb3FuyG8cT+FJlG
8K+ttRG0+efvdIlc64ohX9g0yLLzOD1l+XrJ2cOr7qoJerOYprKSO/aEQtkVBmhZ
FRvELWPJ7v8vmL1n2Ly41h8k1MwjbbCkJ2FxbPuvBKX8h5NqwjbgcjBY9ll1KcGN
O2k52HNxXuQj6ER5CFGXrq02auD+Z8F4aJeDHluSNY7wWUnjksb7AOrkAm2Ui4PE
JRe7J4I2theN2TVrxb1WLssSNa7B0qgcb94pR4+2M/eblmNtN3s5wj8B/9XKS5Vn
7owqesIHAcvaedfj92OdIaqUkgEZIpSOgs7Cg6Kz6EHIC2FjGrBlqwlTX3bCruLO
bEbMzGKdQQzHrn1FGnpSdPmRQu1slogPObWtEtkiq0Y6dDEH0pmzxluJ0DI2/u45
jXdhq6MAZFy53A8QUMByld6DxPTsZe1sZDrY2iAdxwzRzMS9lRdb17vgAdvaIkHt
MmJy+poP0jDVqOpM/KvBR8VFvDYB1MITlkSOKQw8pcZ2NK2T578N2SyZaCB40aJz
5eZd77kG2XwAnJzTDx/SDDM+6TLBkYSivPjrXXyvNNYO2Xly+aqovbm1NLB6Rh+u
8hx8DCOTLfRbVO7o6X5e3DHeuVSFGChrh2pGMXzoIn8nEVSvImEcCCn2LEvmhfCC
xOhf6M5VTUxgPe7/UmqdGfuco7HDHQWPqWnW5X/fvz5j7leyx2dkxzPoBdF90gh6
YPyeZUOGNFQAXkMvYq6woyzRkY9pVnEiXUkF9DOp0kJijtfKyzoIecVLZCLIf0mb
/wuLha08sz96MMCntZmwBFHOuEt9dA8BbHHswKgU6Ezxgoihdftr/gywPhKA+FNH
Js2BdCY3Pswt+cdC+/85VHZOVZp/SL1iqmWkCOC50v75mAEyJxqxphi+ALd5GXUT
kzeVYr0g54Cy75iMt1I+w2J+5oRiqVKWBUZUJAAW/0xMNI5BIqkLJGM/f1Cep/bv
438Quv28HSaIe7k4Ej9lfKd+5eofF+r63gj8rdaiewdF7TWmQeNPalwh+04aPjW7
GvSeVkSIPclPJjt7CX3jFZeW+bvmiHj3va8NQReAI8+kT6nN9c6TYzTXrDST/XXy
iUA4dffEZKLDMQWkWMyNbwwbGZqoVy0djFU/3YSmntLnh8TDL2jhkOxowLy61J+D
6ntf9ULP2z52yCZ6CWW172TXZdrSyoelTqZp8M1Q873izjCMCtfOlKm86XvQoS6n
9XPMohnVBNNlTGBPxfu7S/2B/TuNMuBOOw+2fOqGtQf/Iqt1Hrb0pcPfgfIUN3yZ
HARQrdbuYkL8UBI0+WQ+9y/LBaqhPNe+mFBVHEVpA6dQKhmzJAlTudOOtHSJ3Zea
XgkVbeWn0EAtXJAb/SSIQwhqXJ9su1wJwvqI0vpkI5QOO8nqbaFf3EVZmI6aeftZ
/aWxtMihYCSLkazoF7YT+DiUXI6PDEasZXbJQBT3HUZM2IlU9iUaeqQFE8jI6Wug
VlyC7UixYLzqOanoZ1msTpYiUT6K9m2Le0wzOtQtyF23abF7XtBS2D1LBIXsaiab
DGytW79nPOs5UFLTKLG2v+TmoG30lpbblmz4Lhfabl2kA+OQ69M40rDCahKChGzZ
uBqIi8FkyA9cy2ENo2Yeux7v11oH4hAZmz9mkfj8bIRHjalwyZK0gDpsqC1FgzNz
o1dcOgsKBXygUDl2QFM82Rp/IM0Fsqzh0JtMVt0LcrT+w6g4twr7jQQQ7FwBlmtd
KQicavJKEqhnmxKd3rP944fd4DXdVgUiwFghf7KJRWQxIqme2gl+OMZMNdRzkrAB
DLbA+w+LOJOoUyPKRojkTsogmoAAPv04IGy3NIH1x/h7fsDRbJYFxqGZhlzDFoXA
0EjDed8eK+Nyv722rCjrhsT//ZAjMmZX5m1fcRlaxVVGEhMf6YeOR4FxyUBdzqNQ
qSjTaheXxwFHmXad1FJ4h6zm0lBfdVEXj9T94Q5jD/rGt6v2X3SOhqPytMYUqrio
A/7veD2sR2IUdZVRkDtqhVGxvtMs6VY0roCBH7DmtbYGaKhqQ090IKxkW27gwBlT
SpU8nfrjWYyD11K4UBz5yVXjcyvirCZ28DT5Hn5QSJ70DIqAK2/CXgQ9ENa0Ycux
5NtLo9VYNS88LIUs5kI//OlbI837T4h8UzcRnr6Be9ezObgu7613aliUV55wV/mp
EI5sqgMeNvKj0ejFK98QKF6znzKS8myJoR6yYcZmosU1NG4TWobsQK+XHZJ8ygCA
5ahahiAox9P55/BvpNUyUU/Kqa+BSm7o3mnoNWXU73x6uiylSvQpuvFIq337S2wV
lurpt9jcPW9/0dbCnXM+8+oOhVK+KKWLWhuTw4ieTJFo3mNTW+8WeTP3NYWUPrM2
FSmo4ympJP9/4TvOo74vh9jKWR+lSVYbDc7q8O2CtZ1V2tYl4qwSTwgxEAFw1K0Q
+pgn275khE3/j5V3x1HgxOnjUqYXj5AGhAKXljuYfyx76qw4cMWKx6CACu6bcHdO
rKTWSA77TRap3+swRQe2bJhfnQj7SeuJPB6Xzk/jdSu6+2VowDoouDS0BrUgIug7
PZm1BnnY92Nb3cWPtZXcLOdXdKckt4R5HmnycWEohR6shcxLi0ajKzdVtUSs4wfv
PaLedBdFJ+K3HAeYIpDG2ooi7ZEJ5jKjNZc5/rZ+xqJ1RHoI61StT/wHoRhvEPen
MuvevqUr2GBOX+AuO4+szdoZAmE+d3+PGENU0uP+ntpgWVs2Bccy5BraAsJcU6hp
PWo4AXFXOk7EzztNUvPMyuKf4hbHRHDCTGVVg+pu8MFSzeKj5GAT9f7oS1kU8a1P
FNXbhacIJU3vLE29xs8tyw3RyVTRwsan3ZUHQzZHQ5FOkSfMYdrRHc9ILpuztRo8
29e7nHmg0Xd5c7TOdm69fIwVnGqk2ucYWXPWbuJo2sqLVTR0saDCVkvUT1Sqa0Uw
nfImGJY/DUBnz1zHTCz4eMxWLy2xYR4Nrw13AGRl5zEE999WArI4iEXTCi7zy2U7
jMU28LFzxYrSi7axwmU+ZEc4zs8shYbq6wcjxfqhQL6iV2fTqX4myGXfUznOdiKO
6z8Z/gYyHuroqPpdrabH/y3y5/S0k970wOVcZqwN7YI6ubghDF/PZ1prg+6wNfQK
Q0rpaHRQ0ixcSFrKxOEJr4Hr81IQpN8IJUbeAcC66ZWbD3n8C1R2dsKaTNixT/pU
zJsGz1PYGnKOsMOF2eNIAtkO4jaC+oFZG11Rv8giy8zJQZmz2CTiMKd1/1nxGzhC
bDRii8dzAy5owF/89g9k0sAeNy2uEbDPCpiD6eyXc2M/jY3oMIoVTIqjI3uwpMef
XEbiXhk1XpENCyKsjoI+GVFqPlrBdhlk4Ho0uH1IOec154/+nkRJRFM2BxWVyas6
AZ8mxLL3MOiH1PPhTyFifn6Q2LDmwfW8h2eggMGu5souGZB/eySwbMzf8xR2oM07
rBNYAJc9mGAPkA4xnwQkA4A8cUz6Wa3PF0evArjevuwW6FDIGQ8lvNNmB1csdUoU
WV6doqURmf7WtVcp/+bKMs67qbI1xOLCV/NtioPQymuq45CjPeAPTuhmsFKU9uEG
EB7rTuPVliQz3BDvf5qEKsfGbI7gOPLTtCKb1u04JkAjFwuZgA8wL6729aqOP223
YK3tGwPx0ktnTtUK0dL+RnuwZk7FO+CeGptlVl/plOFwZJAsCezMbKzgEBaULyTw
3DNky3oGLSvTJ149jTrRGuU7+1bRhoU6dl8U4dyeQ9WEJy510vp90mBW5hRBSxKh
7+K9rJbps5b+UgEgUOjKre0iqpA/TI6imzpnHBvk38+gpQFZ/lIMpgMHSpGE0l+M
JYqX+vUK47cLEGY4wrdJmbSaDOCQIroT3uqz1sB77e4YoyNxO+eEL43EdBSZwXQg
4JKkQmiJvet0K7jcdfnZHbOoET3ynOz+ZwfYPloXFqX/lYAf2QWsBAKEhRMh3KZE
H4vuHavgdodzYHQoyU6J9C/0FBUfg1WrcVXs1wrYqaK54wa9KLhtKk19Sm69HI9k
tlczM+4RfydyfjnmzX1cNjiSQsExpZJjgEz0dqQLMUFsTX3wN5tjtzFdqg1qQ+m6
gsSRphl0BoG4po9V/oaY0bYL66y46pQ/ZV0okeAv2188i7rOcphBQBUIl8n+i5yp
RvcHkTizUYzytfU+lSDGcAc2qh+fhEHpHlHVZYoEONKWxqZARtHL7/UOmnnyRnnv
ZtmG2yz2mdWswfcSJN/JWpCpyMBTLNjvRRqgpjbYI0Fdo7oiYDkb27sLEvnvJS2l
vugHCBOLndYMZkRSFFT6s2wIq14Sidahtx/yKu/AsU9rld5lHRPRtoU90gIeVl3c
G8YvVU3mn502eaVmRlf4h02EWKOcTSmpR8+iVgogFqWhXnV3hP5ISF6G84TNgMsM
vXF1vU8vooYGFeDESu+t2WOp0KSlY42n4MIn74+OQMcbpiYaEKRi9gXU/BzORWcd
qsP/ZvUhsQCD9fz5cpa0xK8SPa52GrspZ3q1QKVZP6sofCNHJKpz1mWvn2bPE6mY
9gIFfcuL9PAQRh1WJC9Gf6Bg4FeUgg8sZC3+LYdn+9shVAup08bg842Jmbw7oGJj
89dptpUw1j3/5u9a1t2twb49J+t+oMG5xC2v7z0PBGGD+i9MXZwjpDbyWuRc+I80
y2t/fbMJ72cM8C810aMckOIi+htvaWIwFnnXbf9e1P2lOwu9P12PvC9AOVIPyf6f
850C/kqZ8HzSlsaEeBIaIEN9ZMpVs6Ajygvuf5ZyMPGKmIUZMFiJvmhzwK8ZvQIj
npCrTVwxMGPxLGlhyHLvM6UAfmX3P0fQJ9u6SWuLXccj8WWw9pNQo2rZaTaEau0x
n2BEv0bckVqXslGUDxHAN5SB7t+3wIXcNYPSarfJDREogiFnCDQCk71QwSJDtp33
mf3EBiA3m/sNwGEN4fMFPubvToTDe5uvV+hYRJP/SMt39un+iS8aWFy5/ZPOFRbW
IT7EeWtodtPnQZsccAY5ms9z72gS8a1tfHEfc6p1Nujo2NTl4XjNhTwUUnkvH8Ik
o8Mbk58cL2XcOkp8I/7ZML7mJ80mBDwERdi35MrXoGPQTDy4HP4BJ06ndDoZxAOh
3AhTiKK/PZr6wKM8LtMpD++0cKwwE1QU78ZjyHh04ICagRVIWgYx6iS+Fdss6gtD
yRxHsz/VtSq9x87VQX9xYK9JQpK0Z7xPmrjStUAeH13GJIJTxNJeMnn5fUwYa0My
FWGxbCiz0RTdB+TAXzh8wFy08swHf5069sRWCOzRIpjAX5viSJgZ7cU2YJ7GI+do
24JHsQvJGJb3pE6QeMfAdxSKmM4uEIM8gzHz/5utQErNiHcbGJEvfknSDrekM2Oy
IYpk7K/XX3bQKQiB3SNTohORyPYbbJqOxgryH8duU/ZjdtiPlUpVTr9+UxkhOnrw
GXvPpTFpzKSLcvOSfUZXE4iD8gxDVXiwYkdHCksBKm8CXAnGyiEdtBAIUBOqPIAN
bV5fKVHSkRSQ/27jXH8ATsLVlXPyGTy+awV+9Ag6kbATHheBrOccrRz8KC45Sdl/
uy+WeVYJ+uLsQ3YqIA2vgaWznHs/QuZfAFfA/gC7QQk4i1k5MFa2GFMXHJHEIl6D
eJULRhNJaPDv9LLT1JUuxocKPIdb2ingOTEwjWQ4Q17TrRv07zhKg7vCMrh/+yzV
Zzg4iAJxmtnO4LrNRtO7O1/9t4+UsPrEjnmAjSCWxbyrdfmmKY0G6MFYEj3RBgmz
YaL5X1H4fZ7t+VXKmu77Fc2sSGAMy5b9KK5BNUoSGL2bobaFswpLNpBhsrOy8Pws
W/J7BdZzqLwcji5OdQ5OrLqZrpaZFD8ReEHApQVAUAuJ0VvsI4kn3vctpA9c8ehx
9nBIniFT72ywoV3jyi8bgeZ8B6UQCsMR4oqIVA4oq2dRPlg5ZETtIOi3wfLvOQfy
YXZEGmUP0S6YiWzj3DvJacYOtiDKW8vGZqT5mibChlNxnBQt6sNBduvVkt0SbSCf
m++2fX+ERj2QOATGNkB3bK2O2qJaqP3pvHO/UHPm4rpzEdREixbfk+YypIW0p+R3
CdDGu2xB2vVU6UyN5UjArsc56rkAjxz0DzfBxlGyqc710ItGUqHMZWiZftKq7hVU
u24AFyoZ4kRLnE1I6/AL1dPjjyrFtbXktTXoPpoVLGyXJSvHdYEkFi3F3n1gWNLW
JrD8lLb2O8A28eyoZstIkMJsKxfXpDUEK3GXz+UR8XHXKz4C65Zxk125NN0K3Cp9
PIVMd6MUps5oUznCO3cJ/IkyIN3VQV4oBpHeoqzxvqGLcBgLzkrjKUkm3/UdsklB
H/Vbmua5UVAyR4+cavM0mxrpmsjp2BpL29/kViQWR0VWKDSqlQ3T9peDfUD3wr81
r+8XTt6o59MnXHKK84oJr9CCIwaKBNkhLIhIqJyyX7WYifUoJGn10ynLDseX4MhA
9jfTMAK1U1ciR44reNwPQHcxbEGJxEjS5SlN55zX9Z408SV2v1md8mnwy1pIrdE/
2dao6D26vvDeIseTPPb6CgJofphyQdmXDDPmHgSDCq+vZvDrUkm5ho8lOQkzvvaM
u1Q20e5jnjZJYJWHLP4OKnBfQ59fNwyWWDw0mBLk6iaKu3+wvekgW5T7dM7pO/8e
dVvtKMfF5kslDGHkiWsNsrwvFcLHBYYRGZAxA5MkrRnrKAg3QZB2qWP7Rzz7DH9Z
VO5oUOB1s5Yi6v6aq4wrhN8LBnlXvoBKp8YhQHra2FcCvOuAS1ZM3D8ZTXT8fKY3
ekYslRjQtbBOCRALp+STO7KKV8eg112yyt1Hj8rzOTVkJJK6QcElSJK0LMuI0ZVT
ZCBvuo14SVRDd/Lvo/CsYYcs1EH6lKWIo4ucwsZ/Gm9hD91PqIUMox/bbtlQYaXK
pSvfrMEAgVid1TFMJ8yP6YXlrNZpzhJhgBbeJi5KglXXPJ6JKA+vlGLD7y3V7Nqr
2XsItBgS1fCtcimxEv7dzst3OMeOsRaJXnY9C2Fk2CxEem1Ru33CCEDua5CUHAxt
hCXWzAfCv9b1w9RR3aI1CT0AQyDoyZLCtZmE09o2195UfGXUQkCWO92HhXV9zPch
GaG6GmjqWcKT4wIiyW/q0mk00w4claReXXXBGse9j7oQty8fCp6L3cFZey3DTyP1
Kw/V1KhGFfPIw9Y7cNQhtH8/KYnkGY09EhKIW2OonvVuL9wT8t9q+P1DVAHOUOD8
8iUqlyjfrxio9hkg5JPE+5CLfzGMAQ2lnd3XRZwsTvqdIDztFJyiXooWovBkEtWN
dlniTdopRLX6hmNlAIOAr4yuUwJpE3Ix4/OIFk7f5hyCqi60I/Ay8nMsKxvDBRxy
vlER1UOEZEPWMSAuXAGq6xHswhoRyFBIL4H26Q1lNBOlhx49PzjYOizRpkZk291O
AeufGFAvho2RbWX4nT9kMlK3LyNC4CTDpTZZCJsNMVFLSEVeNj0UslDhH7w2NeO+
rrh53BaBB6n06Z9oY/4O3Ehg9+UD58gKJDlArb5LtVR7EzUYZNggyVXV9YAsLhkm
it1K+vKrLiIzvsQNkS1XczmJoGJ9TbBnfVnB24WvF4R4N/pEnIgO/L6XCD+llfFn
AFnOMzZXYdS5k8eT8xIhRT9RTxmf5KgYg1wIHzPJYKG7dKg/LCp40XXXFbJXlZji
ygo9rB7BUe2R/A4kQF729hXyTa8Y97pidCacFR0peNGVG7Da7jat9UFpbGxLqeXl
CKkMZcRTtk4PCenejEaMHj6i0tP6mAn+Fj2QpnAGZ3anZSxQEj/42hmc8TxfNWaV
sA89oP7qa+ffFsw7M82yhcTH9ZRFW6DLAl4aPJrzRd+0NTbnQ2666fFn7c/LkCfk
FzIb45mokjzle25tBVC5nNgbLN6tCafLKWcfyi8nfXWbOB9Z73rX095fyEblu8Bs
MMyTg8csVM12Rqhr7GyoqcjNLATcRCf2BoHaZbefcFNp7zwZOynd+HjpkPGYh9VY
dtuTmrSEJ920HMcqMyrzpmR7qCA132zX8c6hhp/Cm//Ta74u54evDg917Zi+n9jC
fONrL7YJ+YyUfojIIm31kDBsV+GD4zgU53PI6cTrQYyIm5bBJZ3vfV691U9I2NUp
ADxJ1EXfaUt8ohSmEc6D0fU2Tua4i50NEwTzPawczcD0cFnSdyvF7rGzGnKjY2PF
y3GFaV/9IsFsDlB7JV8dCt71y/VLsEmZ6KSyH86Bs8dNEtVDCu3mAukFU2WtFprh
isJErXAcwtVSJKyeMF6UgcsfzswT1ff/qBRiM/QHgkGJzmwczDlq6eNDz5NMXniT
0UIdvnpk3tdbkciTxtXl2Fscf+SCXCt1X63h1TRdppcAtuDjJ35siBXvuhe0r+8Z
6uYoYA3Jap55JjBvGh2Vxd8QHIc1DvPzCQS3vDnL1JVxyxaik+Z84zmdDsNSjHgB
o2qNsaABTd2wCu7bghRdTPbho2PX5uVl+X1GhE1lNNzsMIEYi4p6k4YjAX4o5oaB
8pHrTQA5qUdFZYAG3HPde+tV4jdm1qwKnOPPIRsWtZ9/Y+Iaszw++Yfb902jtwms
vzQnimVu3YXNR4k8D1WEL/LFh6w1l+qYoZIZJ6xq06D4V1Gn8koyXfZaW4NN+nch
qegpyKl80MWnbHvlpgzMSR36h+Ngty98cMshFqPsxrMqQcCReP89QiKiaU9tqMTz
80xXGmbnBmoXC824xvDJAJzudp4549wVhbgDfNly6JS5WAxn45L9XzQZ08o9SRbK
6PBNTiZJp+T53DsH9HDnC5+U8lUpf6dE3ANZmrcwRXz5miyjzQXhXtF7q+VcZ539
K0eqkn2Yu6/kpZMYB8AmDrzGTqo5oJ8+HPWiEQgRppGpFZAmtClVAZDoD9KvtYFt
iuGjkTTnyYEcViOHctjE+PFBxaWofToyGcgRe5F4+AWb/eyvi+7fwRjWxixzN1d9
nqelZVUVaMBm8qgGDFNmDTRV9a9tf4FZ9GNF97fOy7KDGThofKZd4ngV69g1iJED
ZZGelwPI5elFd+M6EH1ucKYYxoFmvBb25UxfmCnux0tp325f6Dg3rMu2B7v4b7y6
D0GOhN6t6jWrr6i8PkI787+1pUyXSMSih5X1SoJpKl/WZpQYUrus5U0qhnSu4edR
dmf0PbosOp8VeYjXAl1icwAr5XHrh3Ez3j1nB+iJnnEDcJnAsA2G7AnYcencbW98
PtzfKNzpBHIVnDQKKS7+4qbTTS5DtgbMs2tNMJXosTBD70oyU8KypWMrYVvQziCv
WgXR87c1cG9vTi9XEbUHb+kduIB7l83JL4+a7/moxnKJgsVLhXb+MfN7Kayf25FB
5SkvSyJQcwT+l31smtUXOhRZjKhl3iLvB0RzAeLN8fHSTUEENuKM3x0Dnwoqh2x6
VU3tcpkEBfl/CM2EycNxADZTfhatrHkL43h/8qbRBGFjdQE8lltDKfFDN3HTce8Y
2PLSRgj3rfjHjYMNQ7yM7Eu07eLOueJGCmslP4TUDxM9gL6n/LwlsmUXmn5M4Qri
bJJaoUCudTciTSm7DVD5lvrDU56FcGXTqnOWdiEGi31lyzzK7q/OBK2YH25VuAs1
3HYVeqliVfh2HCL5Qa0UKLFOshBYAOJy6gWD5hRlHKZzcM79UAetTkyJkQ2uuBXG
3vLTRWwhtk7oBnXyy4c0nuac10BZEIVWaQB3lR5jtaAq2Net5wk1OckmDZtrUyY5
doWO1gE7lfSx9q8w2nUqCJg/ssxAbFL5w+MHjxG5lQCwDqSRYDaN6bQa3uz5pX+8
iR/Eb3JE8z0dXuNRc463jM033kaYdktFPv3dH1zLs9ntga1ndaggPXKcErSN7bS1
HS7AWe6O6oJbNktFTqNifg/6ZRMyJo6aE+/TZQ7cdagZZpxxrc3K+jmePgjZflJw
z/QJB6/zRlh5g3/bFJxSF3Pys71pjwPTvfNiv+eXFunPnDASSngL+Z2Si5eZfOSI
9AytzMjIncpEhCoZedtcJEtemxeyOjoBnrXHLDh+gnDfLCTcNq8hxcs2mAHML0vq
7CuZHSbszHAZ3YqiOGqN8WZDVLA4WfdWJoWhID/YJ9UaFIcAEx/gan654TUJ5JwR
pczk7Fk8bEqtCkG3aR6Z7tUP/91GCbIDdWYLVVcQ52Yxs3U9QxxBhdTWwCjL/IBq
uMWCe7mHYQmiI+awOgIr9+6R07+mPsh9WoKs+WAP+u9FtRDFJWMuhOoLIM+LFvSk
YHMuAEufjS50supVeGB2nZSX/e9K8Ng8CbYFUX3NOyR0kf2HiQdmHulMPyUMZu+m
eY+Q9IE76IeFp4fRqUkGr3vMi9xz6m16bR5V6vRrfEuR+OhxYSwDe7RNwjgCDGRv
Hl7Eq8Mn8RKo0Vy//VHwYf0/NIp0nHkko5u89JWcM+308fBz2A+zfsVJgiexGcnB
SSX+0gzAQl12lLFYwj+chl3b1t3QJf7Ye7gx9Ghzd9WnMOxuc4+a7u0eXEC29P2S
O55XJsi9O16Usf4MwtLvKs4fq0qfEwDTUS1qZ4zd7T/ihy504zlmtzCaOduGtJLy
C1a8hOLOCXgGW3P/4dTgUD5GRO6zkfr7qpme6YdMO3mI3g9Z4a+sazcK0wGV2IC6
zqdbAhQuCxMzRZN1A1SS04S9IVQkFv6S/V4i0xbvcWT8o/JCeHxB+7Q3a96oDs43
VCyexzHkIOEGOf/7ZVH6N7NCKRQTBWzTuk3cEMt7qhT7zDiceQzwRSb8iM/Aw4KR
0e3Tn90XE3aNPfz/79EGyCvGJ2sYqT41lp3uxsfB4zKPxgBsWLqoaVTweN/saFNe
fhEYZOn2mG2WQb1KdGh2+j5VJZwDtpIXp1jM9mf2j3g2TSU0osgFqNr6eJE4Qs0F
zMVeBeVAQwU8zu+1uAqbVGqCRxdOKaKGvl95eg8yOV4n6hBqPch5VSCvF9A17cgy
8rob0Z1Smbb8pIRzmHjrGxAiY05QwANNoaTNdz25LGZSoBx/VlGk9dQfSWzZiatw
oyeu7b2gLxuYqTHlrQUVyt+s4p6GW9tuLg7lDhi0rZCesXwR97cVkhDwHVTgG3/G
26m583DsciUa1LR/QOd0tFYZ/e/QtEKRawVLeeP9mcrK0We2Ni6eXJ6RPbrVfUCX
q6AZU2Jih802ZevoXbWq4Zt9sPaCfgMYlFIqB3muBLKBz5NVFlAXuyZQgIRy5mF3
s1pm1GgAACIq9LTTDvdm/uC9MCYaTmvCgZ+62kO6A1/+IN0Vew7FTc4f/tjXVroQ
ictgf9fwPluUSTfLzG8wyau2mgjlKq7TVxc8Ig57PrL1a5kHdGyXRuhGTRPI/940
bpV/Ns/mCB7WjPE6Go032V1c/DXX0cuJGsd6k1ceorElpPVPIp2JweKcL4C0Ojt7
u09Z7NqZv26a+DbYbbzNThciUhcs+fTVCCx5un7VKQq8m1cDjg/ckDybFJeOglSu
JQHDNzJ2YkGx2yR+k+ZaOXZuIT6Abq67ynJm4sRpTGn8m1K/v4Q12ckzZnMLy0FU
kda+4XoEuCtvXjS/otHzWLrD8f1GIyxQRKtDl700OTJ0xgVQFEGYgDucfaREd4qe
LzT9wJhWU38D5jrA/YtFNiXQbTrSwXPotojKZfCLjdiwdeC22KLa0vLqnWuglxDe
ask1lmUJBKdvsumfuFzPHnbBUxdNyJ7aqYmBn/aSFxoovYMcDGeIM16wB5l3QFvP
co2apD2nrDAXF10RUMUjYUGz8cyzZ2fgoSgs9oLacBFITGNetoX9ePmFeGy0Wktg
Su9x9usU5Q9PnqOIpypTHlvDeRXiJ5S0jojrDT84ttzm7kmH5UJs7BeWmKRLa64B
UaSnrPFw384IBrgGoT/pJw==
`protect END_PROTECTED
