`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h9ZE2jTgTjOakeKZqMVg0r5Lyy/+5TReAbJ5K6ALrAF9OEkFStxiGZYWZyABSf1D
X8DlQ0txTfzw3Lo0DZNq4xbPOHrKxUEbFxrAQIfELlt0pt8P3gtY5FE1u/x2R+DJ
1mYR1DNwZY5JxXX5G/pufVir2TAJaf2ZsA6Wq5Gf7J51Dttw6LwwqCkL+345Aq5H
L4dUwTs+kizL0+XVPlu3btppnyY3//EZ5dxgFsYUDo7ja8qErbFrM6oIEfj9/+HH
7hrM4TvOXhuKrswU2fXL14eAyklFoFx763pzYPdJLlil1q8hfVILO0gAmrzwDIXB
I1mfnLPFg9pVa6CC88hvp7M9uQKm2viqtHd1RgfX+5O50eajB7LgMHQISz1TUu0u
8KG5Jk4M3fclYgeozZpR/OhMNgS1n5XM2sW4F4dEjh3ytsgbsYI1mieDE6bUGgVD
taRuCa6R+hekiLBoLBM0zZCAzuuLH7r3eRvHlJdJwXsHhKdUWAnpaLJXuDq3XKu7
Qz7TZM9ghJ/0rf4HfemsnzbA7L61sZqPV0uJ9Kd8ZSLhuC8EMyQAOzPTbtESmSZX
gaN6+pGi1WEpty9ebn8QzHAzC1Rc4ybrFzHNDRYT1HLdR7bFWYViP7FAlcwA3+mu
kVBoXFozC5QOi6Z1DIvsBlwVenE0yPUt4EmqVs3Y54K+1lUA6eQ5kFYTkPt3O7Mr
Rlon2pH2oSm2b0Phmw5j0SBxFQmi06AzQGCFMcMTK131mWa9/k+R+FOZ9GUWDm8E
GVoa/9hoDHTCwFtngNETvQjG2WZGklqLzPkhG83SDIlesM+YLNVCk16hMlUl6Pc0
ZCMENH+nzPdOdFoYev5ppnAKeQ7c5k3ZifV0V6vIx7lcmvR+XCH/P4EngypvTr1D
RtljsAz1Hi3DnrzVuDFd6BMy/4YsMkoOYneyPCXglCeVXpo+dlber3VY7qlcXet9
JwksCg6KD6boe2Z3H0Y2KF8erunxzSjYMQWOSaFcu5jWHAhtViQ8AypT15hBMVKi
RB7CenSry5ey3ZnVAy7S9Zog3pN3DMtRgoM9AhEzMw940XsbMnz7CdYkHjgweIyw
0CJ6B9zg+mO69H9J2p/BlAs4EFmFHAnNYP/JNoKkpbYh+bISMt/JYdhfk5IElE7o
CvKW9KHb7j/oW6vqWa3d86FCNfh1ZxCkrqb0vSSg0Mm3knlhf0vrhK8BWIaDcEVc
iiOlPlduGC7MitHVPHab+/wp/WcEOhHxvgnJV5ZFtBsHcpVL4QThXFz1htM87AHu
rzjFj26A3Ld30ETBAmwY0idBi/aKgGoOjiqLflJqKFSQN4AO3yDNhFwSl/YHAxWX
MCvMT8C38mPJg12USitL3xUU/tEa793mBP+vmSt4x4o1lruQc2wDHSkFzyQZ/Ajw
76TWgDBwDHHwrY81g28fMYKLf8x6f/An1PXtp9bkgB7TpRaG52e42Kk8bf304bEL
3KQMeFO1wKUBtczVk+NJs97dhSP4pz6/76DmE8Xz4gt8B8K2MpRicZGDZnbwjPWF
JpkxckZDBqxqWvUbXQhxIyHNBlfxGDOpMUM3R05nLBSsz8OW3gOa8Qlg5wLFgDKy
QMHqiGiRU27SZNfVu/HCOP12bjxqqf+TyBS5inNeCk6NlbKA2a4JfAjdgUuKqQls
JMZJBfRxEoi9hjEheTSZj/I5Hg0MPSy89FDr3ivX7nXL1s2EEKTMLJiiXhYm/fm+
8UmtZonLlJwCPrCTeRXr+Ii7ObiafDntp7b3hwYbqnpRGgxu2YGUTsv0Qhm4c0PP
JCUQTamystCjz9YMLVTzHM4A3M3uC6oXBTthE17zCwjZe0RphxBRsvfS+BNaVGik
SwnN5My3wBfal9BCZ4Jrt0xbn/LahQbTxMN011kNo/alZ97g1vAcvnamMOocqOC4
`protect END_PROTECTED
