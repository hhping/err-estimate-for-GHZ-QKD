`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IbFLqNmN0hg0H7osFq+qEDw1JfIMtJpBgnUmm/FQqR23qJkEpMjk2CFLe9C5xJdc
LgMGpIlcG+0G3dTiG+uIOtXs0qeKcAtt8uk7OZ1ZZHKyZo7zMV8SrnN5uX6To2uG
Ft8F6YD0XuJ6rfsGhpO8ERE2P/7z7SKJ/Ff3chK2Yviokt9DjXG4NTX+vCYzXUxc
aHz4HV0ArFv4vsKfGZBdTJeRysewYDfCwYtEwOaoz6fWHZzLQvJd+95TsSpInPLx
QaLOVdSslKAnSFTlzspkPhGRiTNOH6s5be7DmaGwuYfRYmEH2NeYSJSQRk4nd2at
RQLIZpRRH8GYhKTa9/VAw8Gk4fiKaotiFdNPrsHAsDAFwl7PAswjcyNBVFNQGiAg
vErbRHAVIwu/mFBTrWesnjSazhTlkn0DIB4/5Fqgk+fFuZfYYU1dCynXmcdoB+cd
Hpgt4zlwmSBnyvUHtXFi/KmucE6kDheCSC2BhFe/UDaa3As9ne2Wx4U7PYyQ8SLl
f2c1SI/sXSjbcPv3r/SidUxmfP2cOTrOZc17vQ1e3FMtsU6p8Vef6+Jfs5nwI3I/
0uzDrxqmgiCXw6FNecPabfrfGd0lgh94c9h3zLnVDZJ76zyN5eadkQU/O9YcgNU8
afwsGCm7lio6XYOSCLRwNE78BNxCgaIRX+nyDroU+1Pcp0+Nb0u3FkyMNaAuse0X
TGDL9H8HPYpYSU8c65DlJ2BiMBjpq1RfQQtQNMDuPZ+oczqydURAvr7XvmyuLlQi
cJ5bzO/ThmPN54SMDMoJYZ+ICbGDjdFoiZqhmF9WBMwl0XR5PGh6E60rHRZkXW2i
E8Zia2K+HscElf1O7w3qXmrfiJDrrjKb6NblgIykpmosWeOZuO4FO2ge0MoV9U1y
oN2uojPOzz3ZbZyJ0Ud4E1DH1vnzM0KU+1/pkhxuMk8KzjTSPuNEJnFQRRiLIfgM
IhKULsHFxlYiGiiJgvoh1zdIasxcgGiLotKBygBNpKj+0IDUb283VuXmXrJUkQt/
aHtlwcgTz7o+CaV3OWpDWvvMik1nyIpImw1KMIJiinFpFlz7Kq8FeoZ6Yxr0fXpW
kDXDZJYDwrlhsS0g6AiEWRaq2weio5KM1WeH4EJdkOtf1+lI6B8BbFR6gyz3TbqA
36hn8X0ji1IEFlY2flD/+JhigmwkepfqvySj6C04SmLJ179pL3ZF70ePYOTp68Cl
6lJabjuCFqbFE5TAGAJMJ/9ms05ezU634dmD86kTELM21MeOzXmLx7D9cRDM4TPM
qwXhB9moFoe7JJcmqr6ByZ/rmiT+xoIGqinWPpTHBr5NfcQElczMDFPQvDSOOtOB
5qPz47PxXu1Z/PWMViqkXJymTutStglp1qjKn+OdNqF2Xpxx66NhIr1TkaH/y4f4
2B6VgoAQJUXJU9oSuSIq9aUipfj3J7jmLxVzuSwPt7oYQ5DfEJ5K5uhq7yhQgooo
lbKq3aamAkitpvyeVdQD/Z7lj2PnGfwJvE/L3CbtDI8YFv9cIgvDIpJOiH7dhQYl
DVq/OOsFDpFIab8FTAZ5FKlcDLsxR2VHefdaJyVBpls90oCd7a0DtncwLwkLA90p
z5RVq/8yaBJFCBaDsO8Ce0ieRxSmoaRoFFufjwZUIh71DF8OoRO615dD3ssVG2MJ
6LQZy5vv971PDW0ulSdNXpUV/tRGJ00V8+f7nboRdkubgx4Fobuh3ddZx6XaIGWl
xv69I/KxAusUosr5Q0qclEs6NMZuDOMd4n0HmMArwdaVVwehVDqZXCJ9QdUiwpVX
/CEJa7xdqpVH+SKBa9cBXvwHWoux6DgieWeRLXOosinBTldma0Qbf9xe+jcOgKmu
sDYEwbvNFCkCSes/0zvaYYQ/KOHn/D2J5zBMmlQesbREGlOQM4A46LNCmpE1B5b5
G1JBq8o9Jn705XtC95g5C8ObdrOAsdLDb8thKzSVlE4Ucz+gHQDE2PXg4vKYXWqp
yVN0pvmSgjZ2HfvYmeAEIl6EzyHPDB6jSBmvJN+HEY8yDjxISeo08NS1Ips4j0cc
wi5jlSRC6W644V9f82eJn3Lvg76pNxKhRjVSVvZIi4mI5/S4oTK8scHROrEpxSWE
ZlQ549cwcbc1qwOPCTvvCAI51v7icdlvX0xWrmXwyU2E3xGjPn44ojuGanLbjQAs
LkfAoE9WCsjyHjk9KBXGpG98uGI2nOj7ogdcLLH2zaEsb+8NjQz8dGmK8Opl4cRN
1PjwhaHOWmdf97rPkp3yYyVQaDZ+hZ3AXEtls1hFi0WRtQJvCw/nquDLrtpW/cQt
jYYUZ+1NOOppHYYfIX0wWgqqW/KTJnPHHtTbQ6keu867d5FU/IYvqvUyEvIODRo2
or37m2s4VywIzlCOjCl4hZy9gaHm5YVIoBSK9xnfj9HixnFvxS4aJ7FF9zgvGW0f
CaDweIdQwxv0qEv9P2FNsHHWGDtFIQDxLiffnnR4tWkMXa1w63hF3y6iAlAp1DAL
Gn42LkvQmj8qjc8ieHP6+cNV7q7Xv2aQsWNT5lZ2s+zXupR111MJCXLZ6ygxeihs
FTGss/fSMz/YZkfdVfIJdFf5/KvBk/KFNVujxb6GOa3XrjbPnaSxmf0dKUe4RFq5
GyBmGsboSCvgEuu14ceROD+ATeei0H8UDchBfS+laoHi27Nsc5vmq2tQeqQ7Fw/6
yIHHADgasY/c9aH1m/MDzVb11btkzbog0j0FSlWs4ClK76MDwIARhNYJa9Eyodfb
7U1x0sGAmV5hg0JcFCBobp2SnaYRTRQvUTj+OnNMaUYanKcp1PFk9HeBDpvMAvVR
kMDMDwvb6l5ArTC+fSB68T3uNfwq9Jm6qwiGWnFCyRDE9AtbH1QrbGdlNkNC77ok
QIeGyOgVPefT0oYw8sinMu7tBhQesG9YH6cW6hxwJ8JKAPq7xFzqAOMD4X41rOeY
gmGJKNBaSa2PjnxGsCVIl0EeEruk+G9R5k+R5+EmvJCURcOCF21asxVdmr/L+iy3
bqUL3mmzp4wiEuaCPrAMCrh/iJsNC99ab6OI/c1Al8CtwEE9Oqlna9SrjjPtGlvg
euyqkeSK6gcsacyqqkiHExIXD+9nk5bgtiILsawh6ESBZi27G0+9zl6ZfpUAZ/c7
6sjcKYMdKMtO1c95VmZF7luWBqon9NvYJONQZj5Is58FIrngg2mqml+6QkKb5xOr
dVvTT1du8yvmTqbeQakCFTjFRglUA12ieja9/jLNZPHA2DcNxy9SRqtE+RdIC9sT
0qs3oIqxZE4WAfAD/VtV3PwpJedNimkzxajRRE23zFhm9hEJ5UtzdOnj9sNX6+vv
N8DoYeIEDfGMddvOBoTDEtQvkhbbdexZgGCVAEiSoasUQjILciJWompNTpLrrIkQ
FV6QRjeSA15c2MrnG63Y0It/Hbx2MVclcU5tpy9OSJKyF1D+Q7EZgF9gmjoJ/lo+
8dStWV0X9G3Bpaub4TcC29c4pvbLyHLYMmi55+UJGNmyT90l+1T4y3UmpP76oWT3
8fmoMTS0+Fv9bFsQTNxYNNffQzzGKDV+nMGWR5/HNFQ27buGdDInT7aFRhAgGMha
Tijoeh+7OWoom3SkAlyc+Ssh9UYP/MsBAl6TD+CJR0K817FwOFztIF3tCb6m9Xmw
G9xjC4vcGCIEo05O9+HiQ/JNCpx+khsQd1ANu/hm0MRRCucYHf898KbZnyMPYz4n
J3zRMjInL6OPoQCCFvPiirCeZKcsq/lF50Ep+dhErIq2kjKnFqSI/crzCigR/dyf
e7guP2h0Y6e2QsUxLLc9GVnlPBwBH6qbLsOD+h1q3P2lX/Dse+LxN/6RppXByl13
83zhqS5tusiqevcNZ1dauRigQFfxdU0jVG3Rx8A6wAbRehujFMCFrKkyRC8WBGKU
xODQ/dY/bZSsCnqiSOu+W80Gu0BVSU1N0aozcIxJC559yIB1IvbLcsYeD0qvIX1d
1MRZcGeRJVezwjqQH/W5gaQc6KfxBVYkc0Inr4Nu378uI5hVIv0bp/49YDHka2WU
Lelj/0TrNb8b2V/qUBSS5BdhaabpvlfDOw6CqoYzVzjG5aclujXqZ6XVULS1Zv6H
pQQpBOuv05ODXDdFLTv+MM5tYc+tHGcyjS2JmDT3AMn0UaeeP7bfiqtk1flWNVCw
8otvdJiMMdnn+HxAE81hfLMSH2wsKj32BENc6hWJgzsYWYysCHzQGtKH0lmZWF9f
3TwEk7HU/6xffqo0g1q6Tdyk6YyaGEEc/EQrPKVQiJqsmjiVwEq302XA4bNSx73I
FksiYB8fCA9PU50aEAzbgzcLftqESTxqQ1e3UfSg/TcQWnr6OJ4OKsq34T+5USKL
keas9VoevEdh2p8Q0v5NCIFzUPQybuqFUUA4yborBhaMrNJOd2XGe/xCCNpNzvdr
fLpYUGLF15jWaE5i881anh1nflrRsa+7MH55Ft6wfrwI8P8ZMzf1vi/KpKzbqCrv
OIIpoFgW/eIJMVMUC9mxH206lKrQheoggupo9ihZu8WoCOG4800LUouKeX50Vqse
DSb239BI+D54udbGj/yhsFSUT6gCzSb7BW8sfJ966Ue9tlGYWWCRWaYz/4DTZq2k
UBUBKMHmYNkIZBHvrkI82n+b8Oa7HF3mTEoYixDbFMF+pcDBgB/GTVgKpIDCk+v+
EOrjlk+Y2Q6leuT4R2mJNe/VJnXro0VmHVnvKgDncqU08XrJEjg0/Z8dn7vdInLj
f1iB6L4/6nGfy0hkfSb+PlPw6oswgRVb8AfybEkAw+SUL9ND958VZVsTyBJN/ucn
WJe/HxvJpAE3cIl6B5IKn9obdAhPaQKJkw9Scx91+tzThLL7+l1rF8f3H94vXSbi
ynohPsaEPiMaDw1VIR2TxOl2982yWWFcJyg0XWrVrd50kiJyTEuOnoMdJOzy5II2
cXqsMST3y/hOP4xkhv55UkM6TBMbih6ev8l7OK8eIijeUxC0reDU44ZK1KN5/36C
eOIAAK3FUsQjiMXEZEFq1/ZcWLwIwRU1eC4AaOeHPl+vOPk21HObCGg5rDhfJwTe
5AWr4ITvJZjE51hOrfrFwBwdLfvWJPoVqI+lUdhQRdmFxc0wXC8QmICM7pdOjO9V
cKyf44Yw13U/OpPHnMcrq2tTQmixWsBwxDudCdQAPMJZFbzsqC9UcupycEuos2GK
/vUVX5N27S4XJeQJRLpGkqVx4EW9MvcKCLnfqzdKFBVgvijELQsxH5cWYe6NnsmG
6QZELVqNxYtV1aJwu3N1v7t6QZhElPbjtSAer4LJ0LIgj7WQNDHdN/YNXTGFQ8oa
ji6p3To2pMhTJ+TZq38VY93I67oeGWOpSrr6RbnayrptvAh7pLJzxY0rrqbKa/OU
jT5pZxM44yJMpf4gXPLgn0SR5quCOGu7XMZ8Q1p5pMbtmcnE+JD5pzPbYos67W2o
nAOZCmCv2+GPMDgn57xzI6U9XMpqMEstWRwSsnrFlCI8bna+Pw5wi6rft1ijo+xA
ZZLB1z0eTitVTS5nDwZQyj/vSvjNNMiX4wYL8NgI2zopBq3Z8Ti3V5K3iTOO9Qku
xL6TqDibBYl2A6WmH5h0p++pkCt0TFgQzrFSFP23M349+B9SaXDRiZOtiXXJgloS
+A/OcFaq+OM6yCVoic3PiO0XPvrnTo2JNNkjxtXWwn2C7q9nq/QaH2nGeKO5E1J7
rHJfw1OYRF/UL6A8ueBw+KYiA0fwM9TxZTay12KzTQuSTtc/RYRMCugr+ehP02J9
e7Q5VQUPbCJ0tbWxVz/Nx8OaPIFgGrN77tELcqA4JfgD9GwsC8q2osE0U4xcA96L
6cG6Ow3dlIfN/hfNqgIS7Rqoqp2LKE7SOcR3v0gIScZyGPX6+6qsrBd97yOC27Z9
pyF5rzrHDIfYGiqY5nfrz12Bm8rtXeqbgFm5/YlO9AU31+ThZMKSJtz2o7HTpFyn
q1zPmMOKALpIGbdY6KVKSKFV5ztmGNxAysRIg0GiIARLnmlu47xD0/6ah8SnD9oI
7p3Z9a1eF/9kdGOybkHPfRBA2uPfiZjvtcLRvi7SbxRi0dcZaTCTI9PRaJZzw2h5
eoxET01XVCF8ZUwgin4Gm6yHMmcOGvYJyW0lUduU7L7ieLGkYINe5d2GPfBmfgE9
RUk+3vDfsh5qbGvTj/n/Fv/qSoQtBK2LyTzjoMZmN/nhov8wsoUeTQc+dueAoVXa
KFiTacEjXZ2cShfGYeY/NOQzAEtawAhAvnj2DbDD5goPPkQqDM7dj8jwinK9vBUv
qdrs8gXsPev/pUDLIk/bx/IXQSljMX7ni68wbTupbj210W3HjaW6YOoMb9zhZ63c
WcTqq5jq6po/1frGqjwor3yHJeMhq+ngdx8LU8OV6OQe2VZP32FCN3YBOtKlyZPu
btFLjD1KSDEcG4/yJv5GGsm6N/IkXDhz19zFoMrgqFjD317cnpM936JCfUXnOCgR
LUJZ8nVbapzMYxNEzrQmZIfvY7ecPN+bLNSR6TmiNaMJgbi0II4yxbXcWCObosBC
FnwGRb9Brhl2AQ+xgSgtI4wqZiJQSXXDcjvGhc7FDZNzmqsgB9mXFZMpABSWZrc6
LVo4wi2rR9x3TqYFCRDpSRpI9eANjuX4/OZ6zdhFM675LICJEVbC+3Q3Lkbi7ext
SMRHrquYtvK0RuY/PM4y7eakAf3Pv47Tv30oAk67jVAFkBPGWxTqczflzoLcRs7k
EAxARJetEVt9lLli9wAzNLKiiBRol4xSbDQzGkwLWf/II6co3BwYPYaqPgQxINLr
6WgWrAh5n+b4XLBKsvkBl1sB431Q1V+MwmT8bbBYmo54JexX3kZu/NcUm5L7UWi5
5ofg/AcPsw6JILgjjhTYJgXmcDPrNo0JwY0/omMBDAs3CGVEFkdXUYX/rHDQOWzS
zH06/iYNaj7SruhbE4kulxdbR98ZwBDkXy72flqHSCkCR9CJ36we6PInj8H/NdJK
hKcpa11fJ32cvcHqitGE0P+Nrx9hzlfgBOwIxM5yrGSJQ7tzqCqj5UOY7xnxSbYE
0w3GhJebbqBu+E0+zSavT3J4l9TeaI/T1HOroJXOgeLFuLus/zCXGLN/knYMulPh
1Qb/UGP1NE9qnyua1NFDdYPrQXCp2PwO18ZkKLr6KhRfMmsRXrGqmuTRh+wx98HZ
ILIqq3V13orX+jnbxehXrNIGASdF1iO4C+AGp6pgfAHKtTbLmD+driRjMakg8gWG
aVlqSp9rrzwsP2b/PzoC0UTAOO0/4tFMGgbd4O6DPpjjCwSjEfYXSKXop2KVn5sS
7rwQI/eEIkYTrKgDUEcRqnb9VA0sgiwI5u6q9G7p9CmzATdaxqHQ7drdMfMSRIjk
e0L05JiFPoLYoQyQUJsD9mUxITzVw0SpLzIZojf8pEggtfNk80z1OqVgxLV4E7iB
geeVsMEvlmHtvSzpSG9r3vXJiGB3dQBINUyqjqaN4HNnqPLtdjU//r/3OMIUURNf
FpuCMIUzbrGLnVWN8ffgdeN4DtlHqZ1/XfKUmYnlnNV1QzuLt7IULAYTusF33AzJ
hVNDAo+4cYHyN1QXL1GIZLtK8Tds/v6P9FTLbWKpwW7G93zaY7yDPCsB2klOM+IW
FWSADJsvUrDNb/9EXaELx+FW5giiXvdHoxCg3r0Du7mHdC49P55Aq3v5VKiQKL1d
eBgO/gGb7IAJDzyGkhM7tewKRVEfCpQ5j6ycij/rWBhLaX1rpW2tH5bSgrDrhpRJ
nldC5IxD3v37rwbG1MG17jQnhGbHlyWahXZGG8TTe7wUvNoTLr03VPEYkFSmnHs7
IRvqZnfUJILYB3c3eJirF4IXOc4DRoC+r6z38UGQ2iYQy0wCObqhe0ZUbtgQeCE+
Qsk0euVyWA5TvtpTv4ZOFfW02phZ6H/vEytEUdtGhDUWdWjD1WGuN8fPGaPealOq
t7RRrTKrkOViGEh8RcQhfnCg0KNQ4jlHontKl/wMZYZYR3HvPIzTVAyPs5rclLPm
P1CjYe+pIY0W2ubPupeNaWva3SoX95VLbWSZ9ZGIpCDd1zKC1fNxSWMVvxztsGTQ
21z9ZECOKonpjEdQUGT6SHjT8kZu6QNo+2hDsJxz8d1/CBNbdqLKlRJiODfHEYpk
rGm1sq9UC4Q8vsms+mU/JeaJhR1ywR9ikrLYiLaTW0u7EpD2XZ5PipRbthERzjHf
mXbI0ufA0TfZXv/4XmaNjq9Tos84M/HmwY59hq1r8Pn5L7sf3H86e0orP5Hbpze0
LnXWU4+qwlVzaJnaOoZJKj72HIrKKO7zcfDgmFvIjgKvF6q7mTvR1dxiAndA2Gt3
rPYaKvSstYd2vftAQgoKZAGyzxPKclWPbD+uaHYBYTkogdDzHv1XnO6xBVbFeCM/
ACGoFZdzbS4KIXkZfVwSuza8j5lqBA0MU5UfHE0Bz4YmXfVEFR0JuXLr3lB1Mm7A
B0/8qN5q7SoSM1KP8gfvMC/LqCEMaIjwSWqJE2Aymb6Ut2JnoLiSPcGuS4ISdd9A
QLun2CVZuA2GXJuR8MGn99oxge0TOBkvB+rcFD7voIbDbcaIIkOv0WhLKNR4GiX3
KJNicaz6T087HlcF37joh9w5U7GtRWt36RP62eVSsdMKS+NdI0kcNzHqJlXcJ2zu
zK4SED/y1zu9rTZFVTi810mtKDKtEuK3le0Q2+YN2s5zj74SMoRPIMzKfpSv0mjA
BBKsOh102qasrVAlXsJrGzeKmwMIbQ8yGIG8nT24WTOMqGEc18Jl04JaEHFNO5Od
0WCnsBCTdg1xvtM6152eqR4P+iabyxL8JIaAo/e/A/Lb8jPMPGiAmJCXKI6332+b
fqYzg7NIE2stdGcGWVk1ObzP+7gBG09txOwGhwDyCVA65nmSy7OUTjQ+p+Rp7XD3
ztzAXEumU1wqnJ9vn3g9iw0V2wwzKKYcoY1ZkT1DFJzAoKEOgHngM3cdEovp3nyY
CAbwq/2uBjdisCz5oMhjTuZTbbqL7IlMZZkKwimpVnPSQjDA+2wSCrlQw6s9ukv9
jsBikBqaAY86LFS654W35ijsRKVxAFyvfdooGncIZaPi5xsetU/foiJP/YStrmlW
GI4aFDLmewTBX/sXHoVVjFrski7OXFT1nIkaaBO5ZKNmsxcBsWlra54ICGOPJNFP
RfpaDBH+5mMc+N3I8p45lwG2ZCGUFOEptkHm29XVmfc68fS8oUhXGOkmfieGXekV
mmti4QkHw2mxsImJslfVfsYDs+5Vjx7MymqRSELjmtREDTWdUGyiKtsB1tzvy57Y
1+k2TjHx1RDjjxMZEtAdLUkztVMKDKKYa+UplGvQWcpPXAGtQb/oICNp0ZD2ft/E
syLQP+uSCfaxUtH2MlQ9KDm7HvURiY+yvnQmYAYtRLw7PhaRKNzbdSMha7y88AkU
eIvwaAwtFOIYHvUG5M7MtXeU2hM7Fx/RRKjV+XD3Vsp0ZW2xH+j0HziF8rDdhpmv
xbVwG+HdHHt13c+ZgpKY0yE3SUOk6jmu2jkPTAyblv7AIx3puJhovtCUIzT7p3WZ
h+hbPLxUvczlwZ+X0F/pvCJ0TOoeWYJAozMMuFdy5fmLSIKrfB0cjENFX74gkTCQ
q/JXn/+qsvS20/pRotQX4PfijmMwyNyT0M064Dr9mk01d0e2oeoSbhKvPCIvSbVU
M1xpsm4DdBSHxhp5EUS/rK5xEfxt5/I8Emkm81Sjp72jdb6C/cImLPRaSgf1LvNw
oNIKrytHtU+FjAmb7YP+64DzyfLRRdeorsyt7zdDQC8bpjNPdTPDonOxZkLfpAGf
IN66uGe1OU+cVgYEJ7N6hunqePNylFPCXEQP+1FspfRzUmbp+RfJj+7x7Xt1OlnP
o6QIslfYc+LIVbFcjSj50T7tq3wRmH3ao38tJtabvhtABZETpAuUageKm6a6/+xm
4W9K1/etiEwFXLdrXV7IKdYQn63LtWjAF4tZcz/5aoe39LplSug9ZpaT34sfRSsw
InfZp6fDVCXiyy+UEI6bpwnP4k/eOxeoY+oOtB3I5etBvQ+GqspJQUIkCTAQ8BwX
7L36GZXLz3+jnbDHC097E/IZ/wlonkyDMDYeY5KA8BbtQiV2acwW/U9ZtKGpl/oa
+2tf/dUSij8/Ts7XHAmaRH++xrStatRrK7/Sjyutvx4hHGbyHTQ0jwx1RWxA2nXX
SVmKu/MKplyHFNqscHT3aPX1Wbj3aGveHh45/G/pgY0guV6eRnLsbUEKYwpmmZWo
7uieZrws2DA2NiRG9kIaB2uMv0ZHXfkLlGhxCKB/UgyoO6XWdB1H6S44+dSKp0hC
LtO4fXUWtDqVUAvV0ivNh23i+MmHDL5ZZUKQ0O72I1FuUM0JMaTiwWqVhTP1Wyio
M8UnzMBVnP98FIaMF/R0QbqSUkJdJa0/pohFGOgiAVS3/G99/zNN0A+/aERDuX9y
2vFE4HscqiUnpaFOcPPsjZ+9N4W0JEr1MLygMi/H04u9/zK41WBcknMIlE96RJQ4
3xs6a+HxP9m9hy5PQS7OhGjSvvxfzU+kM9VHQNq+49KdV8A527cc0jegpeDrDS1L
AR5dK79oskPOUwpA16Yqyi0l3gXJi+qKGl87StFynbt7sf+HtxrcKj84pNlDpvan
GA2Sj4wx67N3yYWNwSF6lXkEItPDP7KrJT1dax9r/6t4WYUn8gQMaMqmDGMnDQpS
UO9tUfB4RdlCopr0QcqZ2cL6gF/qWq0dkP7vnlLUACU6ITIjaS5P1EXMu6VgwiRe
WDdUJFL8y8r6WbVJw2TNFgI8JHNj4qJNMzLaQW8xE7Z1iroYnUYCJjnQzg2WXUAh
2KpLnzA9PIeKvCl1mVWZZiHozXbU6IkHxciP89X/oh2KbTmoVFpoaCljMqgXAVQp
oNrTEaMPqb0e2KX3nd9161NDZhUWGH0qyBdlXNCGIlabdry2ixkVaGeVXDZb+6gg
JpANpDpWDMP+6WrRpUD/fNbRSQQxcWJVbOZ2vmDquYW+8vaoArip1iGEiBZ7mcRa
KKn14sX7zPAxYR7H0xcyPQzvq935fDyAOKasFwf+F6AprSeHlrfQx20gY54ELwiE
ewkeJhRBi4l8Mg9VA5yA5eBJBLZgSPefQWXO1OOm/QTDf2pbqVkc156RLHY+YZ0d
b+zs+cEMsMSbhFaj+jWC0cgVu3ISA5Zt5FN2KcxKRwXc6pJ+45v0iaBQ9z8+1Z8V
jGObg8qy5igRgP6xXOyp05jc2tO2GHUPz38GsL1zft1/I7K0qwzL0upP1yB/NwbM
MKRhY83W5cUOKihSf+dEBoGDeY2gJjhvdxOMoXmGjv2SGzv+TxuaFrsGP0gnJ1UO
wLJOC8TAs6d2JrRiXrsI+Wdv4xxbqPF7wxR/TksWCwq8NRg3E5A0BSYIcidxGSw8
JX1r3hvxos8HNNc85q9yjKHtg2I9vJmt3RIruKcE45hSkdczN7LFNwdUBnbDeh3H
5HqW/J0wbxkhwNAQ4Csoq3Ss/KHzahcUtwguLPn1bAY8Wo1fRCizNspXgx+2rgJJ
SApTB9B1MNZSrVDsg5HWM107KVvxC57AV9jdYAUwDc2mtqyuIJSesVAN08Sc2nua
z0Sel7QWkuDz6ObbFm5jj87+Hdak8Sbg8Q0Spu//hfDLf0QKi7CdS6ufzhsEtcBj
fFIRo/3PfMNBDeOb6dgm6EODSD7A2koAwIBuD2Bbk/T+ejMQ44t3L0yE/ilyw57c
1Ek009AC8aBO8JNx+5YXROMEXs/L1+jU/bXqu6JRvM2vPdIAMAgHtR1dACjQVXN9
tPz8ykMuzam9hKFQOr42qWJswaRGiipr3f+JkLWGp4+F7UUO/SYOKhrTWLxr25N8
1A6Nri+xCRNFe5aSybYkGtV71ghF4vOwQkYWpwOqnxXDSjPMxPGFJNjMaViWZe4i
aURqUbQ04nP4zvVKobeGvaoYf+QPOjwkbgbHKh/TwLI6skVcdVB/OoZeoF2xEBy9
3sOy5csUrZt70LNjadjJoQyQsVE6VO1lNqWd5VvMe1O8n+mBxfUMCDKXjgfR0cmn
8FRqC/2GKXgL8mdzFzBIQraqJRV/nxMC5GSSwHWCmMnzrLc63gI9Va2wW3snB0HP
P6xHxhIyNQG8VUt2VvL+2R9GcnPViWn6v40SndOGk+C4KzkMvXSdWDUa1Fwt7wK+
+zrW6N+IrYe8aipjwTv9YtQ1YAAaZMAe/dwXCBe3p55tzt/1VXtYOcYNe2+VbAsW
213NonBl9tFfqYRV/5K5nJrNzYh/tJT5DJKQswipwlRl9/T6LOHMnRWIg6mCAEXa
qP4NN55scjxbgy0/KujGupTEkDVuIUQrWHu+jHq6HN14xEp8/irdWmY89AynERa7
rKkHKK7nP4FncqHiaIIH8kWWM0ScbDhR3tlrDRi6zBngylutr0oZvax44DJ1y8Qs
q19atg0fTiCN1pHll0scQ9HhggkJxaB8s7VpKQGfOBdffwdSAr3euTe33wWo3cr6
jAtY/tK8oHBShssuHwpk8Mcs4lTqJH/48y2hn8Io9edpXzG32I0knT8ssybkqEQV
auTXw51YbscbTnZL1CqH8aUQbvAHu+xwuZv4HaV4o9o0PogMYkFeka2rGSMXr75g
x71sXuL+36sZuZAYVy8zlwH0sUYvNXT8gdOTi93AlN7miSuRdFkZSEvS/4FnxWo4
BEproPZKbnShqv2vR+RvlTy3G+DRH76ru/cTbS3kxyYiz3gc7Kl23dgcf/gKkV9/
Fv1P6VBSBC+JP/PkzhMDgvxXZE0vEu8AJx/kGg7F/gy3xkW3gRC/Lm2hUKCFCpGL
HOmkFtufLkucMNa5gZoNCLcrJjmXysiNzw07nVUbfN1aStPa9/LBbmpzOmQnjY8/
8J2B7SbRZapTCEl9F1nZhtraFsLK7HDcEguA5I+dfIU70mzW9gcMGYR1Rpr/SZCo
XmaCJW/EYVBscVU/Au2uThPCOO2G6oxS7gy/k8HXVPET4rvJzSbElxNoNk5wi68A
M/KELOCrrIPG5TMHO4txgCJ9/HgGHLJgJ72x1Wq5wzQkDgZGOO5IVUAUnQTjPHoQ
SUMvWsFn4BVMLm8kJ3h2Meca1/BiqVsPmd60Izk3anrxIuxZGLZaLmeQzj3Fw38P
WGgJohKPAeeMPIOGBU9L45ngm/KXCIerO4R+he3mpcKnttxE3VPSlUKtICPOzSIJ
lkx9CMDJM4NWtWr7KjJeuY3OuFwo3d6du3hTiA6yb1KkcVyCNyQV4UFrNhFul3So
n9J5IcWfE7bXyFoznTU20HKZqLbaM328k3FFUTG5VGRiLC4LU1L+8Zsc0wfe/wR+
QwBQtHvw9AoGI1oW5t/7eNaUn707a7Iw+9KSxwugwyLQuZ4x4+enB+kOzk0UH6Ha
4/yVw1K4eebBR2R81PY4NcIIEk8lpCFmMWmVjFtxU7HrJv8Iwv1cw5YCy3WGUSvz
Xb+YRq7jAR/A4zJIBx2Nb4qvODBz3dFJdTZzEto7VOJekA1pCkmVbuXrhRPsGoe5
EhcM8tJzyNRJwtVQLTmabKLwr4S4lZI57Uz4fY2jl7eFXSGyqY1qbvlZ9OEHzFeK
E4sjVcxCbtgv6bhRuigsEQYHg6VoNMTwp8uLtn+HfUHKtmO0a7hlRsKKq9ku52v0
4CTQRtnuf4VFKc6f+jTYp3GEq7JcThnI6gilyQVEfONc1Wpds5LYYQdzZR5hfEAu
1aet7DbLOh/vn6k0X+wW9O8hD77PaxrMeWaMzqtkGue1+qVfZIoEe7BfaHCWr9tK
YeH+izcoC7LspKm3Ezlli6M1Aqgzc3vEeUU33bbsORee60kuFsnU5jQhq0K5bWZD
15U5e/l3Ov8IZsfeCU0iWGD3QmCNX+qxdW2a9qb3+CtXiXzWUuAl4nkoMe/fgHgT
kzNKdRLHtlsUnVx5olo78Z+yBWi8nzWyk9IAu0kNBtrAAFBh7fq1hCd0V5yhn+WP
Sg6PoyIxIz4VbN5puX05MGa4lDpM5yvPIA4xtz20wYePza5STmFlFonzzHZMBWOp
hqJxyv6VS27XpLOz0HzstjqgX4r11WCM9uktRHjs+jFu+2f6D26DlVFsORyb3WdV
POwouOVmzt0MFD/4/jNHXp1EiW4r3xE0EttYH1YQuEa17Yp62MHq/WBf4QAl5ZoY
F4dDuE/nILcFNR1XMGMowstty0XLJQcLFynlnAXiS2J60ZAA/p+8oFxZUzaDJGHV
czm4wzH7EqYr/vmOcvinpUVv8OZedXeERIUOJL9c/rU3cOEwWhbEZ+/Vv7QqaiaL
OLhQlQdqAIcYuUrCAGBL38b6VX+6saIYYFErFix4Q41qFzKopQSI1XNxJc1QfRfT
seZuJ6oTset6y4V59BMAzVp0l67xiM++NiJRY/lK9p463zOKHY4ZoGxeZEwtlQZ4
kKvBGR/aKx5d21V0gz+03VcOSARPzArg4DTQuAXlH5nyCto5MKD1CJpQ224GQQcr
ayGV4PvsLEekiSMRzdZ+gS1nLtWWQ1kw3QfySKaAnpKX3DZ7WujcXH2e3mLNqEze
sBqHVkb0AP81/VhAnPNvx5O7ByM8MgDEzbd39mdtsa/7wDRrLophDijaT1sivqLk
NCtPKJSxVbEYI9WQTCtmi54s0Gh3Bd5JBCRFgbpEkuAWgUTR9QZxXwjN38v04kPb
+brYwGpKHKIqjP92yorcAkfFwIzlfvPXC5soskowbTsn6qKl5WoGoM27eqkpNDbp
JJnjK/IkhfIVWPehAIGcN+LZ2GISm75LsbNcdSXXdx2u6QLMjsTJ94q9gsXZQ5rd
vdQBLsnhwFBZXvb0v43MiAZxdU6ueG3EoGTkE5roMbk5BvZoHaaaQqbZEgktcW3j
82UC9kk5Z23sgQus1P0AZ635C8mD9ubloJWUIjaWyWT8EwsM8YzMLF2a+yM+arnU
rl825JYCjuDfGWpq352ZWk77XUZRIbfkdUC9Z+f29S9tmkSMBeW1h3x/FSf6aKZg
hS6bGsNoHSxxvByg7eIdJBwu3g2No/0mvG6theaQboxWSBr9rFzJxIMFZL9nT4iV
oxw6eZnVA+6CoEFNAoEwQZ52siog/zshbYMW6e6JApFeUEfddPiSfyAKNu7VK/Hk
7NkfNGhWFzk9lh6ZaaiOPVmPr+Z4B0wfTr0N38b+FPqr4iJL8+GNwsLfnnYa+t9y
RLNa/h8EWx9BypF9Gp6vAn88Vcv5sna4GSBuTs7mE2mo87qyXIbJpTwJiwfpPUKV
nWsLIU1rP3CYNGEouIdHASyezEiWwgqIbIF3BE57qRf0TPEbrytFLe9RAZllhbMu
CfNvcuk43IfehC0cF8vT5MVg1fjabQivoy8gMURsLN7fV0p6gsRJnuwN8zzVDagj
B+Ac0lEIr7XilEC1n8iW7YZZ/GtTZxMJN0FfKIFDHAtNiilDzeFQR62Iab5uvtRo
5ggbURgJul2X/+xpYvptVtFpxIAOpciuFdXEhAgtj/vuEPxT8RvheKflDAX3mwSy
8gJUOMdP3J62PWcWtAJ9hual9ZI03FY23aMfDiWq7xDbdh4HFa4Nhw6YAgjOUk/U
EShiHNJTyUulfiY3zzc5qsll/Gs0oTp3M06XA0KSMDYiQN/1b+tXRKgBIA8+a/Ws
P+sthUMKuqhm+r5Ko8ExmKPhI29Tlec4txLruCJ7DamB4d3FiIdMCfwUuaONwVQE
JbGhFBdsjG4XluOh8rv4fL4YbMWGEF9kvdUJPC67twY9RaLv85sSGkj0T9Q4rWaw
nKtQTtKZ4h9NMD/Eb3Sh/XcGRVWZGNWEmrjxUJtSO1OzISi42L+QWdzEeOnMct9y
akRKaMr4UY+TlGbAwqxkidV7w78pWcOd0b2EGv1FKnkKA0oZNWSi6RpO+Dxg8Cot
kmwt6EyVfqbHpFDNKm5s3PZVV+o5fhxaSVXZhVJ6uN29aQ3W6mzggd2BL9T0OZq/
I4iq2Fu57tponLwxTNRE+c3+6k257cpay1nuH20ZP3AyOpRg27LIOqbGONcKRwQW
9On33yMXM4EBy2jxnm4FjtrmoJaTaouKyerv+Pjq7qZrmgY0TEECPoIvvaNUE00a
SvPdTcEd6+62WJsBfOABU1CvRg230YVe3OgoagJ1tDLzakXMkLjdaDSYpzM5oC+X
b36Mavwv6yuxx0/WDigFNOMfgtNWKYkoNxdIhrM+Xh3jxLC9COGOgnyh0iU/OEhm
sQDPedKi5m8oSwcBRQKCd6Ft8+hdHf11cvXcJBGJMtJjPmTbN0EPqlFmDdUDtdCV
T1c8iTSWSkaYzRQYszB7kiru8aWKRncABP5OHaQVZsWbPovuz816JAsEAEYeiZlG
ingGiH+sjQnwRUea0TvKigZzvHHVEjhueaScQutvtV4VzoSkb/vzgun19q0oee38
LRYww9pPeR/XVe2XOTvBf61HJazocf22A0m/GwYTYUB8SLHVNLrOVCuCQs+1fPru
zg9EiAk+posCKL3RgYONMgRyy7TxtEGaWAJAwMqzlTKMCOMgM87wX3H3Z2pR+3Ex
2+EbvTicF98O+LpqDJGqfehbUlGDpbUDFnHUJitlvGQPlmDhB8juCiSG8znr9M3u
IK3UxLe99XMHFLslRLRNx5x81U6BlphpNpEw6JAPOvljByayF1qLs5cwPVGrzwJp
lBXKg2fUI4+lsVSgjtmUUfxO0or+pYunBEC4SeHSRp2+yw6oJ3FYa7XbZyeBLGre
Co0SFIyexAft4GNUwWAthPmTh7FfzAQgr1qrr7/S8bnvW5yQWxcoQ17yF/KcDTQz
6ywLwynNMosATZmiqdMEiecHCdY/r5Ruu/qDcFgOLhILJMW2cRKOztsYGoAUIBBl
zfnILADQel/LgYb0z008X9SG12yvfGchx85o87N2OIfseFcoSC80RB5WgM2qj3AZ
+EYizhIlrJl+nDdnqn4UdyOUsNV64c2bvXttikbWOS2m/HP8zLJlp76xDiFNykEH
/vV9MljJJpJcw1jqjuUOAk3bsUoFKdOj6XoY5ceDhapyyjQ2JSRoT5sqYRnYwrRG
4x5WMKZCRzRA9kFVUzkTvAGV1RqlBijEUi0x2MWl858zsrdbgccpCursE3EAhPkE
TyXgtlSwbxRCPdGWkctSLWiTdkJuEdx7AmkP9/6h3C89XUpLBbUqHKvUXreahbJn
XiyHjvXfrkiuPBZJwWMbYp2r/AiA2nAKfLYjZ87RCx1opLvwPdT1+WxF61Ch8x4f
UN6PWkMlN/BBQpYDQ58VT9rDXTv50j73UoKCqBb3igp0s8KONsX0qg6b4yUPWrGv
mwe4MeDCoQs7dsehOB9DNRXZ/oriRYRXpb7HSACL1dfP6fEd/uyoi9844u76Zscg
VZm/OfkT43fq/72ybNGtxx0Up0Z9n0IhwIuSulJU1FhJdiRcpvUmhi/9obixz2fM
pXKsI4ZpH32aGXcaCdVaFRhy+szUTJAhk6jxser7H2IBkSGJJZxNRX+2sHyxWyEW
P+gLe7K4p9wLzYR2v+qspQer+gvDgzZUV4zEQ2+UhVA6rvpYMXyz8dbBhbfjnmLh
ut7Ki65QuYrK1bgu0fzKZYRX3Szo1HBhiS5meN2WS+HePLZroBaJwXeVRis0EETa
yPlcR4LgcRjVYFi9zgbxXXkb1dRSCSOEjAFJFBhi6YAZ/HmmCAuzcBGiqSODy1ql
/AfHPGM/PRj45f3HGqmuHuwI2Q5crdrxNizAbOAMd2Dqv6uMpUFc0vjZYP5faNOn
kL7wFqwEsF4lHQdv/XSKOY5qx9gkS+qdpjD0zO0FMGOE75KoYXB80529XQ1SjnYE
vq2I/7ArqgSJaTKe1pC9SbMJSaKG7rW4Sa6tsF44FaZyOaSTtGhvg5tQZMMp6iKY
N3Tekq+cj6/6/TQ2kc7l3jtPlcH3BiPUebHu1UcM2fiF1aQb9dJErUCfYsOdjkC8
KyKPkW3T5f29i1NmjBW92trGUE/bQc1Vc9C3WaBgoz+QUq5hY4XA6iUn0ktEOZEz
dgM7MXtO4Nms1vgvdMuPyGsFt8qL6GIBmaqtuu+Uq46UIoR/fmdXNbDGSrM2yt5t
AR6NUM3seHeAW64/lOxfz29sSNaAJbiVMMp6/c3wPE6X4151f0Ii/AOCq4xazFgU
eSJdbVra/Ov8sD2GzMhSILgo3todCHzpR9suoKVzVjI6tkidtTd1Zh+zJy8/U6WF
03gJDkKQ0Hgymg+B6SunLWiCIvPYHTuztYffDBT8i2lFHhe3FmTUM2FaIhbYsZOF
uPosSn28tRRR6TERqVdUSM+/oKhFgqLvOkfNhWXuHsEagXJ9RNhDVzNSvnYENMaZ
xgYRYTFtol4ctJrCwyOSA4Ny+Zt/lclhAkd6Ag212wmJHqiLyo295oE4bcAgBB3A
0etZrBN0YiOp0Sh+2zQrHuoldonLl2FyZxpHUN/8ifeYoAHfYzhBGtMXRnjZkN4X
TFRg4+ug7Tky5AG7emqhPQaH/VCShbf8BXzv8BQb5JpcrafR9RAx8PXOGJEBc5Wy
Ooqw/G59Wqxw+KbfJDyWx49YalYoXdZ888nA9LdX+r9FC6hdN+mi3ZNrRl8oIClu
GU190919iofsgXKe12SkvpZh8EvtClyZF0BcxKDbfYXnGq0x37h3hwJOTHWsLH3X
bQj1G8ZrbZzpKTdqtlzfqtHfhhGJLBFrxf/njjHpLvQ+BtUcLOZ+wLnE6OS+2/Nb
RjfXMxfAoqYGOkKU5tXLLUyT7/6fa6iHr50nqoZTaA1tvwnnZ5XPw6bLzfeqoP7J
1Nc7VQywTSsNtTvdjE7oXi4O9r9B5an7YatVtciNMHm1AvaoDNdrLM7MUwLJDIX9
i+kT7J1i76DfitMt0by8n+YyNWHJ+IYqnKs8oE/HkfqdnA8Y22v1HQ/l6VGGuuyu
uIHgnhGnMdtW6oLwlDet/4PoSLFKAywW+UKbuTEYP+fpUkT/SSzl3+zKZIfc6Rze
kspWCD8DlbxDDFxlFSmZwXfDv3cF+JjFiYB6nB5LgjBBm0n5Rwr+ptzWCZL0VwL/
mWNQzEZmsVSN4189TnBfx1oBMUJDwG76W1J88+ABrxgRNRPjty5t+C9Alzg8pN70
oy5J+Jz9vPuTa7uaJa06dXoK5IAz2+I8CEmCeKO/QwCZ51QOCDk1GTbH5CDRvjmF
sO5u+ek7h5AeE/HmC5UZ/AYiRZPZ5jl4UkpidmQ7lpdG18TZgO2V4ofLDspSzqWQ
KcOP0VbHC7GCtXJy/1ScbAWKkvQmAsLvQOVDJF07wzQRYdPVaUEovDkVjR4hZwP8
/lje4N65inq624F7ucoYhGNKFNLVZ0W6i8mD76C6TeTNhgKLeMUwOGVQVsw+fg5Q
iNFEIpP50pMqm0lZFbLbMcwjO3S4pkGxN4+BzKcPFvofEeGkr+Dk3v5mZx8MxsH0
xPq07rWGVgF29Qug3rmnICYutpNsRvxKu9ZWS71wceR1mE+Wzh6ZGRIVEvk2aaLt
uHYdrxMlw4zTft+R1g3JcBN/vsdrNIgu27eHptd+CAT7/PJNiy6x4yIDSGg36p9K
9IuHGRbcn3nW0WNDYiW4Ykhkst2uDskfeb4nbgd3k8QDx+frefoFiRMJM/RVC+q2
f0a+eAN9Y6oWVmeGoWJSYMcdUX5fFqsFX6wOGnbeCCfNM3+WmuUp+ySV6bHOoE65
kdfhAt2G96Afba+ZrvhSX8sQGk8RlACJIFMIuLfdZme9iucNB9A2ciGesX5zDi89
qsG4gnVOyuEiCZlLUdvqCiSAtHaIOMcrYVsEW4HwIsfbsTQw646EsxotiUWNOhWx
fBauyaV3U6B9fBz/0b3ZtXop8fFMZElFZkM4gNL0aitB8cAme5vRRkSkGmWFe70q
JgsonndGknYhtSCop/fYP+uM6TiSawqnnhd+pQUA6oqMGBvROxrHTNi4esMq5ggf
XNj+w+oDT0UW9Q43U4kgvtwrSbW+ku3fGsLxY8uq6AsFvHa0X8cn8kRxqZL7VTaE
i4/juXDthjKzUStY5Gbi8+7xww0Cy++gaVJGZK0hvUDyU2rmBmKu+GveeDY5SbNv
2MKyeKScEIP/jRhAQEF+Q/HratqzMALC2V3nr7lcnMMr/agTc2bPLUiRhZFiBAyF
XwSnUjSLrojMQ1z5wAd0etKSh+Ou9TjY3fBS+Z3q1HHyX1EIz/w4gMX94J818Z7H
iSYhb508z3gKnLie5s18UUBAMGYnWlbABNHctVkBdW/MgGtINFRaycEAW9YEo5Bj
TeqBjIT/qELe154SlZ6jyHb8xtzCHZjDLk1wawHSQA4MH1l8aK2vpMvKESqLjWvp
5Tdra89lOmPlfxesLT+cDkCkA9HZQo7+d73nk9ITpvfPzXS3zTLywFgc47SwOwfp
p7ooUhoy/CYGXTqmgQNyggBJui5/NgkZsndJjemTU6jTwovwkt86rVX8SZfOE4IU
HG/nsYZD2BSjQz70No6+OqR5yFoyEJxoezNIS0vIaZEoAPoGX5I54eBifA4YIz0b
bg4NpEDTq02PRRLoYjCdqMdJRsRQS7/iSyZi6e8cS6P8ykZhYJ5D3pfarM3FQT2D
a18dQeSHWata59TqSdW3ADtGypKjN5k8KrvomNWNe3lQHyoZiIbQjokEK2YFTgFV
gb+bdB4+ALgNUTp7MeUD7a9etYtYGqMrVcyGZCdjnOt36QTfXtb3Pht/Nqx1IWXN
D4/tjgsGpSDkZL1L2T7zEYHgnKK/LedK2FwAilLmWREvz1E0urpgz4ri8BewmsCR
cp/kZDgPrL+YA3RLD418IiHi2FrWHEFexEu9+99FvtraaRXop6nRHrLOdTC9ZhOv
+Ax1TYIAWSk+FttP9SiqmyFsyzmd2o2+iOaZGyB9KZMccPdmWh0oXzyeqfNXNKh3
5PkoSxSkoEdNPoyZUaeuq2pmjq0R5JQhK/mP+CO0gY6p2NOQ0gnT2XGDalfryk5o
nG2aruTbVnKZf9u8/kOWChTI3zdA5u3wFqN/5SF/r+4AYi8caQmjmDdnA209DD3a
DEF4dzglF1naqfMLGyqRk+EyhyIP8KuoAKq+GYLc8RO1kiD5QUzCEYBPNQeK7UIy
Qt4ZqFK+NbSCUGQefogxVz3B0+vvznhIXzcJMAoEipOaEczRWclaB7q8JoE7aUpr
kJXRT5EQnI3ugRiKsqzbK/c7nM3FhjyS5aB17GigugVBrR2GfJ41TiX/9QG2h2DY
2Kgp3LtZMBusABD7SqUSCrjTLAcerzB5ZoaHQnbDyQc/4I7fNu9YrUwUzL6Cwzjg
bYbtyYfw1bPxgzvuqA2L/G06T28YPeNonN1BoaxsPLZwlphN3bE3/Jz2pGS2S3t2
eYBVQl5g63L/SZsI/ia9NHP399PGf3wBjyJ67ClgFoibUHC8dxMjVzHudlsVutqD
cAossDIxck4X8Zf0oNZlmvvWM7iP61xjukZpX8M0cUVeJw2LpslSnammXqxtU5D5
qtUDajTr56gefYuMlBkVMJOGHWna1fEICoRB0cLav+9C0nL4Nk81ZeHmNZfcpj1T
5cIGNK0ffEVgtVYgeph28izdM+61//OGNVTvvwJaJVDfoF2SfuCPwY0DWckBwoPp
xsu0+nF2mf8DvkO9dIGLvOg7J0ypjenMdGfFLL9xm6FQocXNTR7kgYQbCPIB2v8i
ycbMnW3IHqSe+jVZNj6Hu3Vpa2F70Lt3d/5/YizRzyrPqLDM4kP3uFW7+AHa2OvJ
lpe5tBsdpSI5aEzCCyLl27blQUeFkYDjbFY06jXmBUsU/tlqoTxXjahf+SBjwHtS
eG6/uSnPbe2xXwR9MG9D4y6FG8uopkXZO5ffuVyz/zK+PWDS9Axu1HKEd7BYSMnT
cJSECHDHhvP//rd84nhfCY5tymTljYr/fOu5EY78iSm4fYm+PYlureSSBivY3dWc
RwFb/OLTdDnn2DMr1m/83E8Ej60HKy2p1dIKVFPkt6+hZGuTqJRmtzF89Hfs89sE
Iw7AWtzDMRB3RH4qZnzaVRAxXPs77KqfzUlQ8J07UX0dfCoFtHnwRUFBl3t1j08j
IBZlu1oKc7FGdDPqwetGedW4NYCk3Y2WVfF+PK7RuP9PMY3QeQoHzw1IfJKPm0Ix
8V1bD4xV/IpKlQY94E025UCdQ7UWF+Wr5Rcieq/S5K8sfKpLzmmrr4FLtc2Va2Yb
sAESY9knw/sY4O9wKL8Jk3RkYMH9zQrHHNCnkZPU4yPl1YdmJ0AsVFDQfL6wExMC
RBuu6aPemR0lR32MrtvDbfDOZhtX9cL2JryYM9mTMB83pPvdiv3p6FeLP3bE+pE+
SobdM5awgczu48hzqYoCSUPNYSAdoVetfPDJkq0EKDoTroHLuPEPqCu3lY7+pfpV
xdBfeT3A86qZW9ukj/j9oAWxMJxjukXLHn5PvG9ctWB9hMa3JhVVYLjsoa2GeDHm
Br6QorFYUqOnIsRbcHlyO8m08Ip8rZyPYaoQcr8bTJK+h3Ew1aDmK8Hhz27AzGqi
uOzpugGR/jEY4xtrYITIgvGcr7eR9Nh3oc1/iHIFsGfqFPyjBEdY0aSPJ9b5tFFJ
NW4zUmmgsHWJkbnnIl/STH8c0+OdEJQMb+klE/ee/9iRHCCnWv/E42eSldD/R8LV
ijbl0eiiXxpGS7cJdTD3Ck9jX62F4HjunO3gnzVnB15QL5qlfkhLXlnahE1NGOQ6
54heuKvmfN/EsaqoIhYmMT5c/JVOPIXRXeRCst6p1BvlbYSFdI2k9KU66SDGHEVN
4OxyeQNAypLJplZwmSyi/H8EwUf7EqlrveJh2/6scuCIUTLGbdDrpIe5oC0x1qHt
KXi1ENe+xZBw7iUOl9tMytFucf5KZt5oXF1deSRhHbWASLqxXR0chJOSwyYb64OC
7Rma3zO3iFN/NJ4L37IQXvCIy6utBsA6MSyaORzSPNnT0CfA8RqX2UmJNLmwpVT4
dJmsTqjlhzM+aQTMqu8CaBflIvhgPWpb0fqHP6lAgKjvU2rRh9GcnOTpPWfKXnzz
HY1rBYgd8uV7tTThjI6HoNJZAKqJX7wIRnv37H1wqcqjfmTXfPCQEqX8lgdbLvuQ
JsPgbD6RvU7Uo86oi7Tuq+qBYAJyB2wzTS2+vFyDtgYpLfNhRCJNYKqO34ES8iz4
8doF+FCnoPHxYXMsamHicdfL5v71vg/9hncdOcm+4y58ecbZahY8JnCG4Zv+1gVQ
ZEgtnDdsPle+iaPgvQhhE9amVtKt2vgsCd7mR/F/BNjxuC3p/pLWCUJ2B3I8ptKm
0I8KlA9qIF0LlcECdFG3iSCtNCbEff0ixbuh9F5kamxjkihkD+qzhj/7tQhVnpEy
39W0jgvHSl4zQGCja+rBDUqX5YBcm6IizV2kzEe7lb8/Xp3NT7mMDzYvflzEeNpn
20mFcezq+eEPYghXZ+yXQOUmJyCnKPJ7N4+5Mq70ZOV685MmKKEIY41us/n7zVl2
VRhrn/H3aD1lyK+uV0J4pmwIxNLThH0D0rUYQgy22W+Suy/mr8YYVikLm+YOD/Nr
GIJ+pKYCgjkzDOawTLO017Z0CVNlN9pmqtP2cOdNrnjRrwMi1+IOBJae0IHR9rXX
KfMJ4XGl7gQffLdn7/6VBdBmjTDwdkFUf2HinsfRlsIIswfgN9ADBrMuLY6Km0q+
8JSN1MnspBMik8Ug4ToVJaCZIR3wJ/Q7HONSl0Bsvr/ly+lJ3fman3Y7Z25o7QCZ
KwmvfEb/UjVMPxW3rW/+YaRAJ1aYFa1tOd7LwMsKNxEn5IWqR1CCGeCof/o1B0FR
n2YqqPVcOTw1mdvsGm3RAitaYE82V1Jxznm/KrOCnnC0hiwHKQketlfKg/ekPUuO
EiLYa7JCFSkFfZ3SpTUTcuUuSlouvgjuywz9H89nmo0HmUqLwfHPEWbYUzWy9jBL
KvAL6+Cxo+6vtlm9o8KnTIKf+1JyenbQC6Q0egNIGTt5k1/vTIujc99GgcANMjkf
eqVgj/pTBxKFZ4eFAY40yhfgH+6/0FE0OBahJMz3K3BmABWaXzbn8xlrpgEHOWX3
wbW5H7SczdC5MpHEHiSUAKqSPHdSKlJ5C3wkuZIF+ZTaSWBVd2Mc1LsLd5DABOQi
LnPPQ8mjTBOUUqO94yLJXqwDTan/nTo5x1qfstb40z4ZVfTr1rre8nf9kLY14bTc
UuZC8bmy0UwTi1pEeOwkDY04IsYZoEptGEFiWg6hVKyPA2R11L/y5G11b3ovXzfV
7BsTKxCipa+I2WMIXZSxGLwwTIcnhF8NiBv2YbDjQCbjZdxjULVokd1olF2uMLg2
Sl1apFaJa42j1s7crOvPEB8C5QOkfO7KXhxQ1+abXuzCcl4n8uWdwj29pkZdOm1w
O6avXYclHIYfN71DCjphNmljCcOk3eSVtyX/2WTUFaRY4LoPnhW/5ja0vh74Ohwz
xlsYEn5nNhLUTMsqCNDH1ckt55H28VQiA0Y5HgCnzfkaCObJpK4XYZ0CAC7wB7tT
A0fXZUe+ZrFhGvoz8UN/ORo2qnYDbC4PVH2Nf7FotRbfTUzB+jCfCLJq8fEvdmAx
Q94PXyh2TjVP+UhDSSXAmDDDQzWx0jLiNxJPnrj3sYGN+EsaX8Kl31uBDITNP27X
ene7hX2CILylOuOudWnuUOTI9FdUpBVDuiylhcacf2xjhIODEO4Ko8BznXoxBLNo
W7yAaMQtvqzMVIfrULoMvvMuE5kRDPmXD6Q/+02ltPSj0tziXiLkkzCC6PfyY39B
Dcf8uwGG2GKrXzF4UDki3BarXLBso7uV7UHbFQn13PPnc88GRFcdfMMGmuehGBkI
Uo2RPpNBfAFisUX0eFNkgJDQEyhaxT7SKJyX1nWspT5Ki3Ka15QicUL7N2kQlx6j
hwLtiOYH9R91q2Pg8gXTT/t8EAK2GY7IK6xbd2TZir5lwn63d9BEPLghfe/WQ735
Xhu1RVOZGy/l5dID8QyY5Axd6rtXPh0jXLap5Q4krfxuo6o/KrNhACXWC4841l6R
8TAOtYdqJWOF+3Rk+d8lI6ity5MTCmB2Tbgc8I2ZkDt1b109/VGFhwM+3e13cClU
zBX79VpkiM016SWHgY5xUO2qU0cLfxmkGijZ3jSc8D+LhMREhl8BTvytltoFSha2
FXZRZHEACW2+leb38AHo2bsMkOQpMwo9jUhF/yydvIgUoN0G7QXR+4DL6DxNe1Sj
33ybemxUSPtdr5J2B11USFy125YJsPLQ4/UyM9cFq5g3hrzLOqUXUUeu8J+i/UIn
Ki8HcH3ipkZ8LCwQMXtq5i9V8bNp0bLgU00yx1LeAOjJOHnJMAsQ3Z7ZcLrDGERf
8H1a8+nsyU+zriFIOYue/TsBMFyOA/N1GZvo1BZaAnJCWhxll+6ot/wCNBUBVmaS
RBrjOVe1m6LxGgZyTe3BWjyykCCgviiND3HBvzu1DU8CvzhWFV4BN5LsmM08oTXI
ZGbBvkuW8SdqTPcKAPiaaWbjF3WfJgIZiPCIVgeteIEKquApJ3OUKUDq3SPj4PuT
Dc77JgZi7t+D9xB6zFfGxFii7w1vMhxB8JVA/dm9U5ajQUg2Mqb4WTjgoSPgxWKL
1es6WbZ0wULJ1eBDM30rbeslsizAxxijOv7zdQRv/mRYoUNOYzEhFXqY4anR0lpd
EmJGx5hpRCrE5vSgYgOx6xTbXVrPDEuThTqLaOd4tcAFN4oCUyLRoQat4Oug4RrI
NN9wr+pwKqhnxecqdhzhIgRr0O+H7awfo09Fl9qdsl6eDSBmKLpwPvi+7r7ygBwB
mmqYGjxkxGLuvmUWWCU1oJ5R8HlNLBn0ZED8kGJ9uWU60WhRHLE+kTqSZtMau+hc
jqQJY64mm3GnTMYOU0yvkQLgXChtSMALHE1V0PevaQUA62nZ1a08yGaxoTswW5Qh
/GjDtML0cSXRvtL46tSGOtMgyKub/A4h50KcY6kmFcBQFZ9Jsoo7gfBKWwH8Y8E/
GdXvgLgDCMCPQaYuvxEcQF6Uxj0lHKbc1Ye+kQFkNuPbyHSf93miozRD+lOaDeM6
EdeX3wk9bdex6wqchW9x9pKgRiJ6X3EXuHjOo0pBxsfZBPKK6X1SheWZFSEhv0ar
4st/LsM0BY/WOH3H3M4Y1KflC0IcynBS19UEzfv+5UExs1YZFD/QFstsS098DbyN
gSzwyOnS5sHYJSjHCY4Zn4WLr0W5CTvIMa1+FwMqYNldLjjC5hUFUakcNp8I8FiW
cLjUs7Yt/n1ooSJNQjbH1GpmQkrv0J47utGpIIpmncBCWnDlnH+9IbUb8z2zP7OF
IpPDIHhxbv4JsTwlgCxZjJ6Pw3jyVd+Y5AJoQgIgUYqopjWEr0NuGjm8iKzsbKRi
XYdGqZ1BflKOXICXhgmCvXVv5HQjJKWeytWKtqb2VT4LB0OyWbn3lrEtAb8X0ixH
c5m0fpRdaiOQV7m6QCztfmOJdg0QpyQekk1l9k7jLf7W4noS2SqKpMzHu649k3wm
H4ytKSI+MUe8VV8l+DypYL9Bb++NSKeL6wVQZBMxkSi1yk0Y+Bfm28xx/lsw2n31
Isc54gIvvJzodgLSVPAld5081ThqDib7Ur1vmejZFJ6KCk1uGpSHqjMA4PqzGnWS
3O4hK5osTJk0frE91N/Ev5CH1rK7x+HVPAbwK7ccITB97mceR8RxFvF5bLDD8gbx
TITU/QqjZiBuMPqMJ747VYufzsI/wmVCwoSdafKghYz/8KFHekwlMJrCu1pvJ4bi
gyyCCkX9FKmCaUqJphB8jbLobUorUiTRK1z/wifijVMNY/sJ9ICkIqL7+RWRUsWw
PEiSlKCNS+cyTdsX8Xl8e9tWMLjxEoA1zzyq4n7RYA+jhgRa0Rv+wNMlWMLEopn9
775Kt3aIaZPG0iYe+DCV6y7M7GTQatMkGUYSpk9RR4NeiTAlFt6VxbrYyaw/SZsS
AMdTdT1DjZd9XvZFMQQnTwFOZWuS/8sywEo6UXzH+C9AgmVtjv6HdS8BySNyWu7z
2IPUArbPNo+56iXpUbXB2lk0gmiSg4LXFST4S+GLhPVchpk/8GHwWoBhiFNJO0pD
10OQNW8NaqcOk7HMJl1SP81BOj/d4jV1h4oDKwMYRwVLjeuKaq3v/9UIvlFAP1kl
dAul7eJkK+BisP3SHdCpIgZPrJoVX08hbMxRJubav8hx3Pcu1u7Dietg3rfKKBCM
XxkzW9DZ3cnxwY6mGzrGhUz7bMRh3ycVU9jiWfVgHavMR4VI4FAFvgvgkauTNy0U
UCtymgLobke70RcVXh/ya0fZf/pQyuZnKcNZXmN9RB0kjSxqwucc8sQ+8fZibcPO
Bqe3RzixVEuuf+GkOwnKavrQTqEUgJqwX9kxFfwzFDOPveB9ev6lP+uD98pznLZb
B5d/vJ7/LCaQX1NzspC/6FHiBwPI3hwUaFQLLAuuX6uj1FRnB5Fh9X7vXOh+1GJb
Rvo7G02hWRXejNFi4PFZ6B6EDliG1MmPbvFWSTtf10KO8ZoOA5c1bxtnlHwPLhzy
r1WXt7yiaZjj5W3+4Q6Wy3FzEFh61lqEo8nnsPncCMP22DaDnWxXvWf5DOS0eZd4
1qAliyq6iSWrTcQF0B70+62kHpgX0MiLtNhGdBzDlCbeV2jmRAWR2SFlc7RCBiAt
zeN6D/mAx7WXClVkrW+rxZtmI9OyULDuTOUV4e1eKHutaTWxCsdaC6kC5dKWCCts
WTroZMb+tPcrdvvTIAdDwoyuJYG2kfLOfj5CDOmJ8njQuiOCvQI6albDFQBJuA60
9DmR9bHpH4tFVvZPWAIc8gFINGW1Etipnuq3ZPlAlhW2qEvM93086xS0/CJXL7LA
mjfw7vp5ro200KMCHQb8nOj1ahs0oDPJKsajpCLDOhLT66h9uIBsJNtWuSnRgrsH
whdwBxnWhmBmgGKQaF3PbJjBRT8qg+tNrf2XUR5p8TFLGPX41ZLKCdWBLye2n6bw
+jEHEmkqViehM7ZcgQfsVplKuaiBvFhsJJkdSilYF4f7dLhj17EHckaCL42tlI/X
TKELRWijBHU1IcUglVIKKCqC7z4MhAEHLoMKG/uMnUcWD44oTXB1m2QMtm8P7BeV
jM1nyPPlxLRdFsqzX9KdFCNF2ecBX5uwfIqbTLT2Fi8tGl+PjDKI7WiMe+/w0uB+
kyYETW0v7rG8eteck1tDvOpbwsPsiMt68481G00JcvUsAK3HrmNjkn4Kdv5IjcNR
X9BR6a56lOc/05FauQFVzU7VMgjhZEcXbMlPxl7rsPt0ZupuKzDe4ilBxvKPlU6a
I0bPjp3RB8QquRqftyez800ipWls+Qehanr8a2+uOKeDa2w/dkCzv0xXxIgJz7/v
PdeR5k6S2rgDL5WZr2wexpe7AM4thUGDOqLfbx2/Y/UW0cC0KN1vIiMpqXEjy3F5
VbTg3J/4rIyMKMhu6nsTziAkKuUjW5i0yhG/PVArSS5jgl0/drIsftMChCmxEKFU
mZUL3eSaisJyTTsDpZZNF/V4/bUYOYKfuQ00SKSovkodHVlbs1nAOU0PFupqCIfD
QuGydwYNu4IbNRFavifLAPVaGf2Rwh8Tn+5EwudNqQOnMIrv6vOkChXGick16+9L
01r8zisfie2MDtVmUAkfpnrK9u80GKp/LFO4Gv7Afp3HSVJQFanhkYothuI0yzEQ
FQZEMfxzZz4t6QXRNUb9oXvNt9Hf4NN4cRYf8fQbnpjNPXeXmE5JL2DmrHBqK3Zw
3xZGoXmZaWKPmMbxFZeECkxWD2Gynm8z1XHuheWqDEmUqlCQyP5aeJWnn/z8RmY/
Eh72jA1KYK0VOIS6IVLcDy7ylSc/zelOHeJFDhXy++Cw39W1a4sxoNdolpd+Myh/
zECIfqmmQ8af/pTQOLUslEhRTAOjAhvpbdagtQ5xdEG2GPvKTHsxVXV0ZTZDQYSi
oyqPaPxDezNr11SV22/mS7WF56HPvAmf9T4t+0/5Q3pt8QHh3ymc6pG0Y1MYa4O/
F6GZbVC9QS1yXF3Bp2tepipQ2L5xWAfz8mZAy6/ejljBKOGExHUspceK6aVfS4xe
5TN2/orSYnu26trOK6zZAwmTVfjUs8C0xQNW40nMj+1ezcozD7pw6UEIoz0u2Sqm
tl8U6pWaoGg75QoNtz5Y5rub2uu2IVf+yfTCFhsWoZgMm2nKbYkLetcFSJg3j2w1
0unYaRJ6vUIpQmgPey+ZG/SQhRuRhew1X8gTaidyxT1j/kDO+q99iHEMU55yoyqX
8G+/UOvRZ59tKLJPuq98YLVsOUDrQSEALvg0qUy8HH1oHxjtQVbQrGrkPTfzbE4n
tQ6DXHqden+IRYEW02Y8fm0/MCuGWs6l8cuez2yfgSuVQKvGKPewSMojDqtuQ51r
Cg9e+4NEpgTON5Tg7Fdx2aUDJzQvZCGYB8rEVxpTas6bD13UYvrbr0oLqKn8ny5q
JG8zM75ds/h8iXcvJUnxzpUJKpViQXUyJdYjlTzKO0rx9PE7XWWSmNexTJmHxTq4
MvC9uO4RH2qvarPFrDGUPWHwgGh5QGBZ5E/tcDgDBvhaNyBS/e+kRoIoN+s8bN0c
ixclLa7gFjqXp4d4gULdVn+QfZEK+813Daz8INNZK+CELNnkEQzV1QDGfr7KpSF4
6HZHPsCSan7rUkimyVcuzgqEDjWRgli3KNDsJnK6QLXhIiZD8tXIG460wzbDTkcq
jt5sfQlPap0chsxCPtT8ebRwBVxzWqDVypb/tWBuWxXfaU5E/L42R+crpplZhK24
2J1Zn7s20dt+/UMIFrnHByNjTris2Y5wXl0JUQc/YoAZybEV+spUrGU2JZqewFpE
6hOrTeBvwQ/+Zv07I4p/lq/5X0HUa1iIse9pqWdS1uI7lrSguAJezQHdGKqz6BiD
/bbA8g6Q82KVTPxbhW81P3uaPcwBOFt7zs3Mqikq7Jc+d1sosGEyx8uL4OukRzsU
W+MU/uglnUJU1qMqUREAqlF2gtl0ujOI21ac9wUpNVT1dvR6kFKRG6oSLdPga3HD
NpmT7TPNRsRHFxLf/jk5QjUr3s6qZz4bX8HG2sjU2UYPsOan5UQVVBMZoEvzfhy2
EWhFOrsljiCplAKYrBgzERhKT6Jcpf+N9EMtZFDx59GtBe6D+zwB5StznzLjlvqN
O2+RwuGr+Y+mQVuJ9et0AThP5QMKOQTlqclhb2hJqj8mpAizo0VxpxJVTJIKcbIY
RzCMaoJoB4fXYyuFvcrtq+0rERc5YoIkuKBe9twOofL2zYVqZ6aWBlW83XkR2gzV
MmKileDd/nA0ptm7tczVsEuh8UKRzMY1HQ5OJbLZT6V+9PxSflBv9PVFhjx/kNdu
xbLcd4kl75SwozqE5tLIJ+urYQM3Vbi7gtNQpFO/xoSlgHH8Y+ObWSNCgdjbUdCR
BwA5B+HOaxNnbpRYH+B3eoUX2X06alUmXy7Gv4p75cAi7nFkiL6P4MJDEos+npCN
uK6E9a9hNPGQIrSttJajJDHzJ11ECE7f3f9dxJ+sssfvZQ5LBGgjGqOhOnOYCCFL
eh+A6KNTwlfHqyF8paAotySkP7AP9ZNpbY+7Yaj04fdNm08E61JdzfTIMHyiqb94
7wC+vxU7L/bEyUBP17mC9UjTDAhPDBJrWG77Fm+kAK29o78cJqGfFONROnFXRM7/
kfMzCBfCoEHwP1qkBhEcreHct1mWLDoewCG+RvH1CxIn1t3NXHi1RdX4uwJW+dh9
CHXxRqTEgb3BhK81DCIUHzkKaZ6rLu3LG2XswHclQxU2USjflIijPXLsc/dnf4Iy
OqUi4HFlQS24DkxeQurvmrk7BKMnpig78LmPpRFkJTsLnHOxKjhjMYLOG+8W/nxz
6cnIOaY2szYb3fw92RvMjsY8kUW/P+ojm9I27wGTAkm2Qp+AnLu/yTTP0N3f1Dvn
NQtOjz4Ex5tPC/f1OEkLMvhdAiFu/PYXSZRYhJCy5+kSiAGNhqmqq/ZBN9AsL8Wp
ZqPO/zMX8dgKHoJ9ym9axhTHzw10FvXiIH4esYkzy5+aGYnB5W+auC7/mQx+Ith+
HwEWAlreIw2RH9xTFF9tXgqJ35RjDasqV63MmeTwqMXd8C3+kIV+G2h1AVG5GgY7
nkO1qi566HsVu8ZGQ7FN3tB9Qzgc+L7HMt6b7d6ZcO0FvPFWy+SfmepXGI1yfKnv
YhuemAxkYno5FolvEIOD8gExY42xjKoT3m6Md9/xZpEnsRDOKAR9mW+UZZOC00xP
1rVq9EdEWJyWYtpiVYxhvAH7sXQmPrIQv3OYgU4MzcX1KykQisSAmpomAcW9Tqu9
F2vhuJZesAmD66POvJ7tY+LOSpFUIK8QBpoXf3+nHZF61ZZV9ZrKetd/nwbo00Gj
BlJihJTna3o8OSp3p4n2/N2IGoEgW8C/UK/xdoyHv/v1IbcfdkTv3VLzRy6yZzui
n/ee70B33r1AgAbHOxRAusgksiObwBc4UnsONhmkU8e9tkJu0/l6re2EgYEjpGb/
bzeuJCN1mUNCM2/ipnoc8GajanpFlIXWGKYX9cdojNlFhq+BeP5675R8A6T0A4xK
YUW8YfEbDBPFVBoOtrY6TagMs4MATkrUYFWn01vXHbglSmqAAbGFUV9gLnQi1Lna
+LQ9rl50n28GFqpyyJ6BUanVIiOjDnPlbATybIYtgo1pq0ciT1Y1qpNH7wybz7dy
ZC+iM6wSjsnhq/QOpoZjQnGXGrj9bDwhEaFt7EM9DZNlEw4Y757gC93Q8JgLx0l0
aiuMX0fZJr8n1xKjBEOYqFE/UDQGUPneOECol4Qhiee4xGDq9xKw0BHjZnOQkqm2
MXowNhxlwpLKtpBvCVnO1aI08Pk5/LO7GgTmA3jni0gx9pQFIF7uEaKqD2VgZv7h
RXNorE/tJ0nId9jpPcg389YBQVP+pxE/+9GkkAvcTWWh6IIxucrQ2JVg2XNnymTH
s+h/44kpwHYMp7f4Hn4VLfxQiUHf1ImFLUt32QHCE3cS/UD10yGSAj+afD3Bp294
a0SkROX3PMx+i41IbteMFiGVFDmKYYXVkoEhNrumdy7M9JX+IaNznQ1Sr6STqN8G
aKIFUFyCFV2MbI0f317Pj74O3IXwFkDlg0LtOswzqBQo1zbr2PaxD2DxcX8Ah0/J
dUBBN0v/O7OGJ3k83ir9cRsjiLmcSInkceOwLuDb75C6hNtRTxdVn6pFc3i3WfZU
dmUREgFxjWRhyMDT7sbJJMmUFyS5mzTDcAQ/aSHAuxa2kNFzjvtFJ/2X5ODIf0gR
8Ln/KYMgh67MRJDM15o98l7dYSGp5AQitmThik2h/XyAD+83X7x4rvbuQPhh4mrA
Xk4eDI+WF0scLkg4SpfK0HkQq6cmsU9Fa6iuAa7KaiSfhNPtL3D0DhFrTJB/8R+t
uyydyDWlN3WJe2AJA/Eaa4aDA97tFzKBpNS8Xv8/KKF6RTnUj3Z4e9zDbBSj3/dP
zhplNME/wnPNJBKD9PAzYGrAWkc0xtvOnHGNngme7Q3Bjr7UTt6kahezjTfXY+Bd
dvEHHcpmEVtWgfeUwBOOVC4cTo7u7O0qJgMjEFQFbRzDUpjdSw9I8dhf49gqAahG
mDcNzGdezLM+fzawOdZAyZk7ZxqCKyDVwwBdsuI4PQa83z48t5VVSq7rBvP84Qfn
0PaqAWv2ZztA4FuBxWCYrkwuFSvViglFAJrKm58vuZQut/kaSo6A+yfD68Sb4kbs
GNL0aPLcMFCMb4j3KrMfzTeJv6tbX4Pd7iNvkGdwo3w5QTuEWCgiJB9twDK3P1rV
rbJfPY3hGi6+6NkzpMPmq3dFgZdVxnkiSGaXb156owE72WhdaLHUQYFu4CW6DEPa
5qy6xR1qg6obZQu2ak0hTuzC+XvXOkkPq0cNPe5s8cMYGtMhAH5oDn0rTJS7Noiy
WLYQYXN2FTM0muSI72h7zsyRzQ4JwV9ZSkhPTbnpceFeadZ46Apj7ViaWRPrJ1OK
5BmwA5sOHPzizZbB6IKH+hW58qi23A3f6QhDDUEWyF/BKsapVwA9hYzemSNWw/N/
Y+FzN7Hv22+kCDiF6BCWsj6tDaYKen52cqMPCcNwqopRg3Gy3ADDaJFcOM67X8X+
Y/ytH5smHWEA1PAarkJtQdhF2tLgFgoZCFPibdruXJSIaFwEiXkQnyZoCWX99yu+
mTtYExiPKXvTTp3uNj9dtOvYPbr2LQgyKc1rSgFXBUuNNZ7uwgApRCHa1Gd2Dljn
4wvA0NLhNQbCyOhmHTiyQ+wGA2X1d+yPI99dA48PFEQCDbCHAiCpo2FriyrvwVvy
zixmDOg6gLUr0CZ3HVri8YLjybQx1hdppCeOOuA55Buh1Y4XRg43hHTtqdgIYOc4
JPuxMd401eRaQDtDGmMl6oF+8n4wy9ffu/Cfh/RVGwwb3lz+xfTPAzEjJL4aDEEu
Qk5m/qFaBbwenS+VcHGkGuF1/mpnpRlJUz367soht5c5RBdrqjIK2GMaRqzf3ijz
dz5Fyj+OaeNyKeTZUbQ9px/WJVSQZeizv7+04MBH3dxiM3oMTRL8GaJjOUyKNAIv
e67G1CBGZPAYfqHKiEHSheg7gfOGlY8dEMzJDcvoiM4LqC1uMdupTLUhPDuqSmI+
DrIpURkpif4BiRxtwxd7vrULrUWElAk9hvVsDvKl2dL3+0EhTCyWchxuYjd/r+4d
wHZ7+MVtrLC+8GUh8/A5flWIz1ZYCYm3h8UhSVPmPmBZW6Bk9J+t3zPeLhdgfQlS
5/WQkJq48NYj05Zz6bqdxJgM30kO/hz4yq4KkbS8zX5zMYZgMaL+nQbrevDaEPni
HmeW/G95VCRLft80Ka05jbzn9kAYNtDpcZGY3J1QppJIN/4nPedoUNP7YD+gCmIm
a4egbDd98cW7h+POSIrAjpFhEb32zWyuTcP/ZCE1qFxPhChzxTsQKIrxz/fztKtl
rf6z54LMorCH49dgfAEgMj6W8n4SLC5C4NwSJUCaU8dNwMWlACdTvziKNttZY4hU
g+kYbiuH5dpgaaeYISBlf4COrjAAAJbghO+bTgzxetsMgfDeHw8JjDsVCre176Ar
NJokKD48bgOX3PisJ/AteL/9BEKA3vbfoMQG5a9gXAPbR+8g4NR1gH0BPLQR1uYf
K1xzFOK6cf0jxGSzDVdpvgZyBqlYIhRhJbkicSLdzSgDc9YesG5RQPQajlyqpKUX
2I1CwVIk63JvVOHKgP7A774fuzdcw/Aywd942VzYNX9h2ma8Y4RQnoFfy0vcpt3J
b4BXvVAN90UKFvxgYzezdjIuK/rKzKCRqcu8zVqtxfW4K0XS4VT4p88MzzEb+Jn/
sINNN6TthhdwAn20w7hFcpTK3aKnLJdHcVR3M7nPhnuncTMExUZjIdQSBQAcu/bL
3JG/K6oqEogsf9DOxer2U4/QfY/kdzGRN+nWIzl4ihM8K2uzDpJMiFz0RuHBsXGQ
DkM7DaFoo18FJLekh/NlVVsCYbNi2BYaYPUMCeTh9SsnwT4uT3kWvGxbPPqhNdtx
wP5oJiVXLPgMWSn28EVOezIjaJsdEeRp5nBxEzW4dkRIXqLVWE5hMUiG2rC3D1TL
y/ySP91D3vzLqEDE1cBhWykcvl8c4FjhN28mONFXqhf575kapvNkGQVAgJAzDrsI
wyNjCsia/WFn9S0mjGp8X0EyaGvIoHX7Y5MpYFXrhCnj5NrWjXm4r2COKJy9OZ5o
AZ7ciBmL0uA2cuGb7+9fv+V8KA+vTh6mwZ6uFTJW6vK3pj+EqgJ1yFMHI6viAku8
Wv7xDQRm1fHEmTqkmiqfSzy227TXwGkqHfEA2k9VfG4WROMmX5wdS4lZ502JwdEP
DL8XZUZKAzC/igZr382zOAtjn7svMqaiZ8O0efzk/+95eZoE4NLq14Xd2qHmKYwF
26B2PKHRDE9rHvJKSJfD6q4QC4k988VSIuzOsFCpoEliVMe2yg0sTNnPiqvgueC0
1hEA9EMbx5SDCIdyZYD2rBVBCGIUaf/Kz0YUkLItws+pJIUOVAtMH87S807dupfM
I3vBEzphloVz55KU8hbn1ICEAj0nXZcGCCherjMG6M20ss+/jutkazaZInJWY5S0
kHq3b+FW7VS0JU0e70ylisxNLfeHhBdj5leEqmVnHBaeYW0CKBL5HPvbjf0ZFOKQ
x61VURKzff0cmeHQnwWHhp71LXqp9Yy4AhGMnk87PcunBtYeVtcELUASpPqSP0zG
Ls9dKobrNhhylSEtE9W94RbOhLo+EFMbL7q81SrcG5ck6bNck7BhzhSwCxmKJlFQ
TF0IhNZx9bnOnebPzNUePfpeBGSgsC+8U+nPdRQMhC4VfyETBbqAxmJ3sFtazyx6
DuA9IqTvuNJSqkgkRTKV9yT+VyN019VXycIcb3SxAF9VykTtrBL6TuPW93NJUdmK
IINEbEzL8ZCr0Ws8c9EqK/t+9PXYTDHSxy4L4J2JaksEFcXxRmzoKyMxhX6LuR4I
naFiJfdD6ZPUzy7O/z6O0DF7yhbZqsBRXUMe32Tl2uvQT+UDUvSaU42iqR7Fq93r
6IrPas9Ov6KuiK/B1QKiNVZJdHejJB73QnAtTix5m2zGanXIMzf9nA58hlfOjpOW
WV9fI3owvHGq6GMwLwRjKBKZIHbhlGTaZZnaDSm+9eEuU1LIwCvCVwX3mbKgzTJb
x1kl5VR9VM2EaFdWsgG5N9Rhp55vRu3uj2o5fBbh30nslxMU50/hj2d9fn3UJ7Cc
FHW6cOGyibZrFgp4STRhKoH2aLQmmRJ5891zCHkRTk120faXyJuvn/rY8/YPdzw/
eOUL+7bzrSMlgH3bGgmyTXrPxHrQcz3OrsmitAHe6MvbwPDRanQsmpvrYIbK0Kts
DwCvRwCNZDzzFfN3aHYsdZP3tTmch/h0x8PyNOOeq+t1jEwytJLiYWNuDlmaEXxh
ySyP7A7LTrtD7Tq5eUUrM7W0irfN32iH0TsCM0fPd5+IWr5vE9oKUyxzg2hQJEX5
WYg8/sUfNsJQr2sUH0athoJ+gzoedmlaB5x3F+kxjn2yaGS2PMJYbx/p1lqH70+d
ZCrWC4f2qliWWG1IVryr5EpAExP0jErRZ+GxT9YYsHnVKeywXsFogpbLnGirBvbF
PnSmEOc84C28K6jOkENueNoqgLLfgS0us+6FZpu8fA12jINqLtDYLWMBpSJjl1oh
vgWRpPfjNaMFCf8kEv9w49vrAfRCxoORQwiHkp/CckZFUeV2cxgV4jZE7vqXORhX
jcGym5Fv2zvmUE17VojmJL8hCW37lENZ+XQZRH4/VRdj1RJK5qoD+o3k8UDewD8a
6PZGhw9rp0Jm1agMfvfaNhIlOc1/ivhjqbPdP80DARM5+abfTgeaHBHItV0wc1fE
59QQtIWNuhaiw4Ksmjc243xhAW8KuCRVLC9P0NrJnzeJrei1iYeG3EJi5CZg8xC3
qO1+YARuFiWV/0qGUeJZJNKbNQYKop82vhBX5vHio5qdeYcNN4duKdOtqzek6JOq
25J8vn60xviPHE7eK9S/DuX8OexywGxx3A1afZx8zuUroRsk6IojtY5FGr83TW/+
ZIogRg+st/CAuzGutU36mxuNnAuEYZW+jizuEYT8NFz3Eb/0Asd+HO9As4mzgcIe
UolwJlCYflRptZBJjvjXhIjnvGwpcpYo4H4d5bGvrv9GB8H5OnsRME2N5zNuhzM3
rkiNUYp4Xq0N0O98hiMI7ksHKGTjh+lEpm18jOIC+Al82RoipuV63rM5rW+ujsKb
xTpt5Y3hIgQi3K++hLMWAisa43ReMHZehybNmxsmcv4BiQtJARMme4HkZfxE8uIl
5XtMpxOBFQzrb0YSDnwU4j5kR8Q11HkNE8reu4Abk1CG1b81dIcT7DRP8iVUQhxl
Fyyc0iTk7XJs5x6eDoQoYKq4IpyHEQ+LD4O9am+Nsr2iUXAkCIgNKoGrh8UuNuJ5
On1AGdGMePxfhby7J/KT0zD0v3e/Q2WffZRkOWJEAshhG4juN3ITyaaOynsPfxRT
VvkdccHeSTEHqBrdm5fqRMaRG4fjWwpF+NPvJxhfRc2djyC6ESPjeHQjt4XBvLtF
nzk/Gj8DACtPd+qrUfdJ4xalywqDp6hdJJ3ZCNN/nthdMPZPufXVJMtLEEv26IoW
dadSBAl8ZIOYxcAxEn0Fcnbn8iTkHabafRZM/x5j5+/dMzn+Jlmf7GuRNSU8JcFQ
wEmpnATT9JFIB0Z9rzICNIISgYMNlNTQI898UeiOHmdMxrQ8Smh2KWw0WDG7Qfri
Z2HNlny2bdNdoNWU8oAxO13sn7wcDULbO49c+hDYWZNIKtUlyrAMBXBONQUNXR/b
FQT3VQUvfMm/FrnarUmrQKl5y3wCkVHPuMOCoFLZtU057QhNHQuuTAqjltbNerFg
MWCP9NGza3joxm/Q+67bBf1IB7Y4NrtcO88grMMKNOAO5VyuY0oPL2LMgFA9wj3u
1nF5IX5kf2LeeHnwvB5gnQ1kY2K1FiQUDRHf/Lcss3YBaUWRV/7zfPLyJ416d1sU
FBRbQDiACKbQxPv6++nTG4esPAZ1JmcR39roY6HoRL66rn2tCnC9STyVLpBlMVsm
3fMo/mTpmcy5sHNCmZzHNB41jdyJMkflA9jvU+2XZd/hjW5k1khnLSMDWWK1HbKL
bRBepXNs4K72LBhltqY4RAfbUXLccNxUMm/3us5ruPAlvQNWYoOOpCB1GTKsCPGy
UhmqPDahMQvZWoL5aGeNVAnq/G3tTIh0ovw5FKY03M3l6oflS4pNkh01EUInN9mv
GqFwjdSRfQ7/tBQRO3/swW5H+TVdh9xZwfEW0VYny3mJFRmyvQXk1E2LhvlEKJw4
nta5MmoN5WwZkCBA3RgN3wDN6SgqLvGikhG3tDa1ZOaXw4DR9Ifui2FfnjfLDhP6
oB8p3uqKSmt8w2jznjR2ov0MrCUwcF3aEkvvIjnOSCKnc4jiwcq7GfGZpnlq9J9E
y+kJ4yYHjYEBILfoF5Di0+73G5iaJekytYiDnbO60Fs2fsSEPFjMokt4N2rFY2lY
2fSqYPulzOtW6eWo1qBz2Vz5nfPgnZXpjmXUAy+8yLs8VgyhCFpatdbI2YxhhXv/
IrQtYAFfGYbCyZ85VbBPZbYs/67xWuM4/ggGyjbhG9/dD8zj+Po+wG6fAB9Mty2s
CEtx3nW9kNYvOJ12r/1dWc52MGT4ZWTVXGX9oXSp1CGWuSjgygLwVvPXYkXLmUQk
Lo9lDUqKYOye/7DX8hHQ9AWVQiAuADQp/N7GoCdE1r2SEOUlyVrKQSd65qC48QKe
ueEqdBu/mEBYAhE3rZ4MIrhQnTjd3A2STHmbplMFXzwJ5RMLLALptXwFxfKvzXME
SwmQ4xD2548KKhuBVHWoFCCP1IPGmOe7q0FO0VMqQVGmjIEU5y1cyt+Ww7Vd1k90
nGhPWAbDkm3RPtdYYbuuoBgm6D2BqfxvxUCd1u1Bj/v5Yyysh2w13AqxRYAuRX/u
fMwn0ZEyPzjDXOWP8LLw04xB+3IBcr02gugL+vVIIReEEjAlGaJImJy8gin70Mw+
Tg5hmihDkDY8tOLml4pcmaGrcM/sG4zVYqmI4wFTYlwDNaGj2Ef3kaxYFhJPM7O5
LCPKdZHw+nE63fcaTl5tL1b2dAR2ddSjFdSotqF/85wAlgtzQ1bpEAJdR/Lc2l3w
j5HnZcY50HU05QyEviDvd/Qm0wUgFZgw1fJOGxOAubg1ToNOLjSK4+sdxnh7snKG
Ea7upnDS1nSH5HxayvYcSjjslExmHk9UMuCbRaukzMyY6OZxkgFu6we6I5yeKVnZ
0z/JWo6q/I01eYzY4P1E3Zxr8gWzQQpYazKvS/IgvDSvfm4mnUUsTh6MbHr2BFNm
D1ca7R/fVcIOxXMMzyiQ3y/Xhk3XAxDGUwKIo8674l6auQPft6O5FyK5w/c0ociA
NiB7Bfp2GIy50+XD31se0ZumHXJn8GEvHDgt3n87YlU5zvciTvbFya3r5/FETTbw
uK0wmSuRfFBZogatI8cNYh1kf2v+qTs/vPqTQwSrxVqld2haiM4/3nU0MRypEbEH
YXlrniQ1dhKDWOcm2cotDl/UkVhEZQHAag0P5JgAGVDoMeHamZP26kg+fNdfWkuU
ZbhdSDjiPBHVcZ8/sf6mLTKEt797RtNdvC6NKuG5FNXgKsIU95UiSVaWSApw0oX8
kddt/0wZgW0vAwhwtGC36OkEprqCPqQLExe8xxvKqRx22Seavdy1tdTf/bEThxRK
//lIFMDud/Ux4wYOTkieicOODwad61UkpcQRtGPJeiKHg+ehBLVehVgqF4L4ceQD
AbCyEnYtvVd0z1yAzy/FrlzFAMMHMqT+LBDLkyjJqdq0R/M159Tm2IWadB9dSOu4
9/PTaM+xt0g+qlrdsALGRntQtCeN5fuE/ijT4iFL+RzO9lpi46FZJGwmz9zmREJT
NImdbvrQJ1lJUQWn32k9ieSEQfz0Ty1tPJhWnCibyHcZUG0ys1Bj7zqjGsX5gOGh
ybJLP7XN2xFF/E8tJcdPjL+bcRooAiI96kdQFZQgClc66TTWsfmFr7fR+i0c9Jma
nl+V9mNVTXKmAcAam0BjGGwenbPj1xoPp2sFfvELfX2aw85OuuFWP835Q+wkMd45
7eb1tc9KSbTMKDKzWUdIO1ev3YLmMUV5PTNvTE0VC6C8qoegsrb+Zl22NjX+6JHm
tU5/xveT30K0ZDaVcfIyUhVOj9GJAAsxfznQhAYKQFqr/uvxiGFQesjRnO4Fr5JJ
vI3yLYavaPmeFX/Ezfcyt0WZDSOYKYqfgqhXzHUspXp8Zrh+ctOfZyeW9xTDKOlx
4MdVxX22kqA5hjp/0v8WEwnTz9xfLzlHJ65I6sBL06Wiv/zwzg0xRAaCPZjqOgnM
d5PC1T9+BPI6RPNYcx6AWnc9MDy0+ySzj3eSk2ocYMc+wJdzzGwf8t027IvwbcjM
+kjPwM7D6IZI7r5FY5bYno4crdGhTENH6vtkZs6wWDWdOV11iUrye0zBmQCBHKXT
KzE0Az4YnUWA14281AMAc4rIjScuyTc4USW8k1EfE8MripYtBIWhmtUHI1mf8zy+
bvB5vDBTEJb988015KZ7qu00MSApzINI4Sy5v6vHXjuFBhm4kmfcvF6McsUlbdQR
bgWLS2TP/Q9UiHbIela/lSmFxpYZ0EXdrTJs1sZH5Sk+oHss459SyLTgSkYX2LzT
rhoolr7gh18hQcWdkT2mxIZOFBZjpqpcY2vDNUj2LwKDR6wmJwiRCiQl15YJ6cJO
XM6NBHvumk9tMpJMdW3nECaGu/0OKfBmyjONyIJRlLX0y3N88xghX7+vvnx/HsDS
UQJDOV3iW2UtJZJs5genx80hJ3oWKrd78Tm9LLnYqs7PSMLJIuFmCe+7N+wFodAJ
7BI5Zky++xNOHUUyLxcJCERJ6z/v7LsvpOjhbFXhQAfsYxxpcHis1FxytxCYkuor
YSe6Jir/cNIFsL7XHEuIy/M/npdiu+kOTFS1l7V3/Ce0mkQWD3tt5HEZsEe2a6KR
HkhU66H08gSk4vgD/IRXlsjqEGPdXc5tgZf2jdmnsA4BiHR9PaP7t8R1V+sQNS+5
AuRBCPfjCRhC4mJ0dYWz87I+lDXHFsAXnCE3zQMp6LX58JasTFMj/1zfkvHO8XN9
/IiDdM2FKH8w3d7hGwlW5GxIs7Tew2hykP7zxBlfRGOxfEeptqvIzTZ7LoeqrKDW
2uEl3InfWR+YPRrnrEudb4w/0ayqtUGTnqiLpk/ByOitxMR7v33o5wc2eyokx4v1
/dV8j7kT1JHZUvONY+RQMIPgdKBJV7jr57X4dA+YujNIPcN+lrmIQqoAMXzfp+tw
FcLaBkuohN6LDNbS4jSqVi/1UVOFThRwRFT6AHm3eYK85CQF4Wc9TbxCuyjqYHe3
sv+NA8s2iQZwzAGpjhmUL44/jvXM4qrc2yTaFdddfN6gfYYCL0WqMXQWlX7nNUJr
qIr5dUz6ay6ksv2EwxYvlwSoPN8l1Ax9L36DHbv6Ty2DTEMJO2K/zhjrBlUpV2iQ
tH7H1LfgG7vpubT3R0P31NwsJ8JbY1ydNt75IXREK4bOtDFVxlfnDpXCIPriJCnL
oWVTBLMUc9l92HP6WIK8vOCi+rjwUIgjUNIKRD/CVnqOoCj5h5sbCKdXR9It3vir
GT4by/NXSoahr59XX8HvSoS977y1XwNeId+iBYF6wqBpqdngQhiYGDvno3MClLTi
sVVl3N8xcyOM82PtZnT076j6TdG0Di0Cg2EgtZlb57quwWY+WIWSpAcfV66+LIBJ
tNHg9Y3mUJm5BZ7rGuKn1k4Rtgkcf0KfBm97ivm9qbAxL9Jvk3jAvyapYjB+lfBx
2vC3ZQEY5FfKD01C0/ZzBVnYV80/GQSMbIFydTmjqdlffRcCjyRcRVy6z80te56g
gtfWE8dqVUTKDCSvkCFAxTEfPF/cYcgLUw8+/ctLIA1lrpy/MloGwrsLXJJYQJj6
DYPdP3mPDyw3lNtasH9MoZzTyBkxf6Jn/8Qz3vYICQ6zOA2r/ubaoEFFzrWJGWFA
bOw0CGDPWJAXpOJPSvqE3OrDbN9vPuEqe2XPyzcy23xkR5mdxINgi/CF201L+3Af
HSMaf+rKr/ntDSyVohMn4A64VosyoQoLMAGmlg27n8Ip5jxGCq4yVgzldQAlCzW5
LoUbM4WPv303k5QarHJDPbVIhnQVr9bkjJlpWN8wyKiHRarUdaj8uKZJM9TL/FJZ
q2wBrNalLkez/FfRoZqhnxgM47BhFhzwLrRniATdgmW8mkP5JCvgtsLM9tJwpum7
SQf3Vpnt6iBfp3ha/1LxirlsyEOazKCQL6ZuVGC8BjZLDYnohaP45+9BsviNaP9B
N99HAx7WUdeRb83hSw6/wVy0ExiYsz5AY1ke48mK+2iCpeQ2+7wPT4GnC9bmQxE7
kjme4fDE6rAuFOA6bC4S826GZ8ftSulcuT+RcX26rAGlbrqyUYBCy/kzCf8ld6PK
xZQlSDYeFb1H1HLd4s+5nlnn0yP2RnJ52mcMlPRKl5kxXVA2Oa7BZhZUJ4+fP7AS
TJmJuaTJLrFUq379K71Nf867BwZYNCexGwqH1Uaq4LJ8xw7qXl8ridAL4/xVbcpF
QzeWBIg7xy+d0d5C3/FT0Q6v0rzfVswDkGs/3NbS75Ph94Vcr00cXbJynIp07oGR
uvKhG3YwlD6ZkQbztIDvSAR1v94DBJ8Uk+jbrTImK4bWPZj0m7kK2pkbXqdFCo4g
gtVDlxrhjwygUj3cbL7LA7P3/utFpyG91fktIoy4OOaN4+JZFLl0NKTIlGF/hB2N
fTvLPz3uXUk+YF6wKXHEVLpP0C4fNOako88UQODPFR2inejreiJ6ds4amc+D/6hh
9DmKdtDUQIL17kFLVNPy4wtm5fEU/k7S0/64z6XZDt8Y6Ld/OzLqTr5b+ZzCx+js
P1nUn4hZJkQvPgfGMQTFyVmzRkWy1hRQ779B5cuv7CcTxCFiABl2qVRvtIhVJQU9
NxZc9HuQsOeTal08G9COtqm+n2F1DnrHJaZWgFuY+x8TvW0TVcYJMK4Vh91h3CKJ
Js+bmwy9vZgi3WfKHAYhQkrOijMPE4jM1g6QedRfWrSWURKutHNmakD+sPXMMIZa
rL3eofeSUFuJB7GsjnoHJTDGXcos24CIJhZ+0rzjAhjMEC59toJaBNDM08JJRzIJ
J6148Mr/tw/z+TM4fIST51AwA772Irwfb7JNbez+FyhFEU/Kh8FvuiYCoz0PZMna
TdfKmCOXfZmsXKctSwE3dkFlboXnO/jeR6+tFsB2nlJC37vIKde7mmTiHJ/NEg/h
xA6I8BVFnjlCrOZgJt/yE2ortcQjaF7YZFiSbl4PpQNS5VCJRBNBj6jhPaP3q90Z
Du18OFK4erN9Ogi/LB35WPkid8qb34Ls3Joock7U3hcgzhi2ssiZZPD3dRa8qFaQ
A4sFd3MYVYk3ziuBkVZpSNN206FypNMEGe6P5ZN+kAmYwPK/zXHrAQBd8vNk9IAy
NbYatmxH9XCXpRee3c0NUZPUjLMgGnzh+7gW+moXz+xF+/vuyzGK17aO0IVE6Vsp
vQUDD5NeBsi0e3xLwOrzbTIEEC/rEHzzz7Jqok/MeKnUnVyNbyu2Wte7nbliVb0/
hHWDDo7eZfn1RnS3YR08NcEcn5NKjMa6SUOcMFg0QvAq2x5yhrUOo6HE/hhG5V90
v685iW/4KuQxxAUUMA6wJbrmetw/Z/fFuBaNpKT4ba1UC+L8z8XPKcy3wDwbZ9TM
qDSVbZSEhHJ870MnZv0W97M+moqgc75+LbNGPRyQcqGRDiY1Nl//tsh5lZJn02Et
FaV00O0Z7R7ShYPuQUkyiB3IyiDjIGSLijs5VmyB0ABDrUyruroG/A1Ae4XvZ6sN
l5Gtab6d6cSy2kOAnTAKiA2b/fvYR1pR1zFwvqRayLJ4M9xdLnJsiNRrwjDJznQT
dMW74dT083QUuI+1kTCJ5fO+5yGE+NmZTseEJzybnRbh61RuefE4UBSOmv2+NUlS
Tw8gqPELivx3GUp93YgQ1/b1VkMB7apHjSK6jV2PIjmlMX27HOzdF8ki9XFoKNMx
L9UISglfP/fNwmNeszULkzRcD2LXBjxm52oHorfYWdeENFP+MXZemh5RbSBKIcZr
2Sta8rzSad4/8bqKfsF4PAJpeboXCkMl8nBcEJ7dpssXct62vu1HBK/BJBu1Lr9C
9fIn5i9usA8390MLGU/gKEJEWjrK/vhnxAgOvPCALt+D/T4vN7t6dZt5L20RiyjR
gFuVs93dgv/k+gFWtydaQBwwdHoZtjn8OL2DRQY/sK48DoPekvx2xGJcRW4YMa7a
PSZiv64bRsl6v4Rn8WGnLt99tKGbviS+wSw+loQt6WMS9qdzFC1WYDhExxOMM01Z
IKbyjftbQbs48JYLCFEwcWFseJQL2u80IYMYeUjMb7KF/Yux8GFTl3Wf1/2P8itR
SB2DcMpp2v2REOewFm9aufZn1VDsjRiOuWDOF607jdtXsiCSlaSpQIJttIoG+Z6o
N1uJ5Ye0LmSiqPgSUTnYuEQfIOz67FBWy+tIwvDLGVKR8u9Bp5U+kMUcw5l53g64
zSyNLBhJ9z+c6dU4aoBMXDMTukcaoFHUXQfSvlmshto/t6PfWBNCYuUtWMltxeeW
095dYHHzBR+N6vC+VwsgvqJhoalrJV9zJEUAKHAQo9jXygHsPFB2MTzBbpEnJq6k
JhcsbyRR8YyuKaW4Vu/n+7HFeepe80y6YptVtJllDfj4eDlObFd8akPWqRs5X7wJ
KQImwQhOkjh/9NM9hTFeq8orcnY6aZ3ZI+fC7HIZAiB2vleWDMxvC1BFwH7MXaAE
c6w05vOE663+gpBRc/Neh6W+sI1pfXcBbUHTW+o51a70+0A8UvskQIUUslkaZC0a
qGWZHt6a6RZOFNUj/5FerW/Uny6VAVIt/02XVx1D4Ec0qie9ZKJHw1u+zqbcoIfa
gHVscnuVl8Iva3G3aunhtZ6x57zu/okLRry4JYKcewvYCuWFn8WiPhtAMVzUDP2M
fTvO30X0Dfs5NfRXKnjerRoil6DWMN3Msv52V8HywJNXFnn75YIuPDbnoFgNb+uT
Hn99Yn9ptN/V2gdVkUvXGXzLNxb9G6PF33hLBFXJJ74yavJ6LMgydi+H9mqZaM8E
S2DFJzj3q99M+PvcSuWFmPCGOv9g+0i2d6MonRkYq5gGZx1YGYNPSQXKckp8V1gR
FQfGrvzuuXXh9fk97J4mqa8hYf8+VbcsSF1YDe6/8WUntJDuF5wvtStXZTouyhc6
2gThAYjXrt5fG/P67ZLgriv7Sv2zCZwC7JF2YQgqI7wSkHgzqo9fybAXOG5Bc0vM
dabUvAAohErqPsO0eltgR2SYQmry8cqwHQ2v0DUO81Je8YvjmWGnXSMlgY+GV3Qj
fsqaYUIDOfQkDb6i2/RsCrqH/klEXR9H0ZVDEjy9JScJ3BdBjPJsHQbMVjnBPGi/
Nz4L5F7PXpp5ULynwhH8mHVHsVdS8NpkKb4hfwWbAnMRW2pssOMvUis++RtHHX8F
WcjlxhRzxFtzBwJEHVZBeAZN1LuSXR36AR0hmYA3VSY/ZaKY6WuEECOH3cYV0PkN
SNat5/fwyv+jONm0OmFYdKz2Z/LrFKjm+40Os6MmZBuyih6puidyRjNyRbYMlyS7
v7qKo9tzjn6qSv8YWPw28+sMcBTzGgFEPCjPMIuWXHG2jOhqxE4vtn0XR8/ZWALY
XvJpLE2yZyX3bj41085dOsgYNPWFByYopSKxOKLpo45W/RpzQYBooSiHyj9xj5MV
M28k4q+Y1FXRrfxgT95McL4eCk/pWOYhNxZsPA6RuFZhQ3wI2gJbuHpCajjbRSD1
UdXX0g12pAJzfkXf73mEcLMgg6czAKctPOvDjUKw3l97VEBsuL3zCtsZ72ufbJrH
95l8d3xPZ5UvkyZ2gaXUXWi2bId3VamzHJh/ZbbXWfasg0d7QEcrCC7RvUlsKECt
OpsJpHkdXSKOUKlbUE7QuT9nDAVqvcTBIqmUPn5eIFVkdT7KQNeDRr/dM0KRxX92
MArx+LvbUPNHhOVjbry1V4jUohehNO1zUhqSnwoxkdfMdH7TXkfRhfgz7rTN7kC1
EcI6s/GVK98oea9pDDQ0m/x6XuxxmmurT6/cjsHPRjm5hQNTvPQ10mCSAcHFPt7E
j61OlaSTaXWx8uMGWsb6ita3X+wGf0x6DfrfpQMCq4s8HaSZQZ8mwe473OVuGtT+
9dt0ycMd90vznHdciozChL0Ov5s1Kj+J9Oh2/gcU+hKJGkeqsCffySU/ccBEL1jg
7wfgYG+WFK1chCdAQl+A59u/496t0ukv1ZAX9hE7O/84TWkYYrI9COWm8buFj0Fr
IuskU6H7drJDluQN/8USSfsKhyTS6MPLHX3qryLZaefJ7WgfnhBnFfF/T/N0xQdc
S9oocumAqqHiuBk4Pik6i3ynK75JQTajQw+M1uevt2Z++8gFMNHlLJZ1UPNTwX/v
gRwEqaFrO+MH4d8kzEA0RguWvHCkne9m9G2iFTwfE2e4GdOswzuBV3toFk94vf5i
xA/+t2hzeNS6IIAHP/gBfijYV1O20tBZm1wBxGSJpGOqMDqE5Yw4ZRVQFGF5ISyI
Bym2H+5UkQnzhHr3TiFmZf7y0cDN+byiPAwz6ALbj9gXYuOI3VegCxGEv81oLOsj
72t6ln3rjZ+AwOXNSZ2CR2HV+jh4rrXxY8EtGQSJLckXK9XfsGLZi3K+3fGrxrhN
z5pIrLB4BTqFuKW8KCEQIqFgIE1eax7fr0LlFspPFMfekGrki+2k7zaoArKuz0vd
s6X342fxE8+9RFjnYG92xxZgHyl24OEmGpNd4AkmL6eS7plOo3c8u6rSmidncwvf
/vG657qis/QCOHWRSaRwbDwGDIhkiF7gjL2lRN7xgZJZkKrk5lxN1z6wv22kSXnD
3Koch/tBbIESKZgqRwNuPG2HzZfbpQPiHL56xEqfWAyLaPnFqhQpl+djm/qELvPf
4hA04xq/qpRAd1QIRyLRcrWFLOy5F5h4Wiu5FnxGPRQy4GZnBkJpPSVYAlAmbj1I
ZFousZFt+Rxx2oEq6lucMo2uRUntBRiE7q3BcKR5JFxPzebUAvR5e2aWpCW4o2kD
VvXeoFif5Xm0QQeYuDUukhAeLmbGCd0SE5fezKQr3BPEYJQ9crgivq4zqUpFnqHv
dKMcUnETRg9pPNopkddncMVLmeUHS4E6rf5ymghni3mOk+dcbQic6KGMsPVlpN65
+Zf1Nlg9jO6Kal9Tqc1RW9Q6O34EC/3vT37HxxwV6US2CH0v1UCvMqkmcR4FwSBI
/Za9nGK85Q3Rpw7TVKqLCB9fgdxphRF4DRyfS0yGz/ofEk3iBDyC/+6c31aOibw2
N2zN8ij9dTC+rEvMyd9TDb5GFg28rmq/HSrFNS6hi8EgyRa+uEgpJzQ+3AtYhS+G
/Yg55qKN0E61wHsKyEUFzDjMGX6iUGeqm/0g/k0dJQDh5eDVBWra/RJgH/2THcGf
uLKMUFNpwTYJ4W276KUda8xUNOdri7TJncOr8NMCEJ+lLN0g0mcouBajMNjJxfgj
Z//c69meDT5hfJ+hGksepUhlfVDeG7bpuzcV7/9oZzTKTEoIEpTxIY6OIOnCCknI
vbFNIzFhBPYQNYYZ3Om/zRtG6sAmB15zIZ6KYcgOiBV5I4Lhxl+kFjFfAWsr4l7/
0ZHm3Yq1I01dr5I9fIJmKdMCUCpTECCQRFlZw4j76AQV+ISCJ/6UcVc0PbmBqdvX
8Gq6ngBoK1ZkU5z6nkvXLTBXpXMr3gRY92Ypr5mTuxDN/2BwYr4DeQ6ydxNQs0LW
FDgLix0WHwon/eJbhA1oNbhQ21vCRls30nf+8+EERmyl+GcSvelafDfs/2s9RhGc
bgIkwouHztULLk6MORk2f1gyGyLdT/knLD87LGAPHTt//niZAXuDrW33cgyYp5iJ
OfKv0aTYPrPhdiThgCyoBf68Sl9IUsfetoJZu7IS9MeFmG5wCLbiWvS144ny1fZO
c97GwVCtcrj/cxxZxDf7kgBiyHGofKpVz2A4lvugFGCreFvVX9IcXNN3UX1QZ5jp
2Satrqy20VSkepopB1Kk5QmSve0NKflYhrm8plRJSZCyio+58e1JlN5Gn9slOhj6
xp+PAD0XSu/kaHsVDLIY+BkQOqFKqp9bossXZTJ4DqzYZpuTpX4Ea1hu2RF6ilqQ
IO05rWoanxs/kGNmhp12OrC4IQ9VhMoFIRykEP0pdfxABqOWUmi5pVGjxcLb7k0U
KQ2mIotKrtbSpKiDyjJ3SDe+Gl+FKgxKoH/+uvhiXxrDMdqSbV8EAATT3EtgkBlG
nDpqRfMD5XF04pYer3P7edEQya3iWCwNxihCrCnsMdRxh8jpVPCUay6AJ9YRtcAV
LiR/QE8SoClKtVqzjgYGWnEyvq1kezmpY9TQMR4VqXjkBjK+jvT7Gv3P2FH1wYDr
E3zHIWRikKshR4JQ6Fnzk7I8btEfDrHmJNFiWvzpBpPbWU+/xHiVVVqTanxhtjJY
WFGYE6Mvto7sbBDnXsEvMvg73wrcmPpnYoMObK/zqorW3daNHxxtPe7N3XKHSea1
BdjmDFrB0zm5I/6Y4TeSydyqQP7gUT6EzfdODsMlFLjUSwY5JbAawmQEaCSPKyzO
OsqgK95o3gRjGYtM8YfZoi6aUBDzYKPsrV8/x0AG1G8/YXAaHpw7zpyMGqYsGH5z
zeXsn1P24uFzjHKjMKEdIFuSVaM/KjUiU+ha2NzVhFOTpLL0pv/kVKsFV73c3fw7
1XscP4lZ+TWQtQ3YXAuljvgTWG28jqhjmIyoeXYAa6Xohiej11wAS6hFdLq/dDr/
MPlMV+eypNeONe/B4CRFPjw9EJVRmFITmBZFj5CvNhZFn2/bWK/HNsoimeCoUPvA
9aKX2kGqYxYYWr96UlFUT4IWVPDZxeUYzQ8b/QCtXgd7IPuDJBcKxW+ea3aeWcgS
i4pzdd6UfGmvDrc70Y4mzTQbI8n3Z4ma1TyIML3NlYq4eJkesYxSWBKRzOT2zydF
8iULkrDlfV9+aBKLxEOtk784Fu4BrsR7ocZ8sW0X7LiLHCVfwTHBKw0jog9fbpF9
nn1eJDSRO446iZQuVKslIP3Dhfty1h0um4R4KvG/XdLgthNGYSeU5qv7cu6t26qU
gLti2kBf+UsMH8ad8Hv0PVe/4JtFDNDDCl2Vl+tI+fvN3LpgU6MI752JjDqHRX6z
mRpajibzZMU1hZ/IzTEV/dh5y66dQKkLMElqgd0yvba9ofXTJ78oLq4gkP9PlWhJ
6j9eVs54nZsSojxrqbpCQdkhcQDJliV4ZAArg8oLKnOkDLd0WG9NEZHKBN5cLfL+
ht260IldASeo6s48+C3BBTnOJMGbFRblG2/SAI1OwbyXH9YjD/JN/Ao9f1G7Kfq8
sVxPDCYKksyAuqbIB/o3QCbh+7KXdV2goGqCdqHlbYh6FNAVRWW77+yxI9xPRFjq
kgy3YWM9KzdkmgsfIdlJdcoIG6x7GIGx18xsEgEmxDi0Rd/pasfc3k9dn4WPz5wk
s1IJNBNBdQPaBk4CmmYoRqX/+V6OaTIiS7FtdXqZ9LJC1norVKc+5YS7OTLMU/UZ
DDaJ9BngaQdouT37Klbv85PBTWAx2t7gmc/qbai33/EUFQj/iF/4SyXlRdyq1jtR
gzcm/kQ9HyCTrVbYI/mxqG+YL6UNNdFC9Xd9cEicns8oEBfOIep1ACl4omiKtFFU
nYX6vsVZ2TjExzqvp0GrUYZNELwBX0GuB5oBRqqwUBUXaIotbiRcoT+zLxVf/eWz
nQ9/Y5c1HPBxu0AU5Oh40p+Kac92p/sESZV5D3L49SsZ3E8VGHIt3VPxnngE3eTc
0/0nz9KxKHggrROIikXbOOsN8osY9SNGX0HjeO1OT5ePiK9to3VhDJOQUQ7DiWV3
9RqRf87leJMoD12VwQmsQoZu6wPZXVfunSqk/ADRXbYqzemLvoDs2ivNVIl4u6el
SEnjVdew2UcZPgvF8+b7AwplAMOQkUbkMCCkJZHaqkHqD0MYrfTSAP6Ei1ABAj00
4KwEz9XHI2GNvQTBDHdfCNV3Jjv99n+1gpLk+Fz1Axe7QB6XoabxS2j1VbuTHGe4
Hyv7Jt2JklvkPGF3NTyJV56P+HFsS4L85mv8Xap2Uw5YRhCcNiwL7abhHpXIC50P
Kq9sDXGl8wYFUlUlsSfy5am3IY7AyNigNELCR2xYQ5NbXTbjbWr2O7QCd2tQJ2DT
okHAOtXqmMaTr7icB9pFTW2UlAUMUf8oJifAhxczMNzmuxzPAha21JRJNStphf5f
x++vFH5LC3HB0KnaHqkOBkusslBSKa5+QP77EfOfU+Ql8MCj6Ov1IokReqMTj1TG
wa/z1ZMDyW9KVkwbK4A+8KPHh/qNKIf1QgqXa/shoUOvP2kNzoCgDU04REsrqolL
60UGMjvCqX0F1ydO0Wh8Be3wtTjc9LFUO+QSOmG73soxVPurlt8nsjsVzMh44VZg
z99+ClnmhZUBbRPPKbX2ZEj0ytXRYMGIoMa3NPlO6zJZ919BLjN5wtcIUBk+StSF
qPWihap47ASB1tzNpf5NqhRNdBFmP0f7FI/xaZQsa1J3QcW3dHk9ZmClKzWr1Xk5
R9NEHs8z5wTO0pjre71CyPU4IMFvjPDVrytCtO4EJEFW3P78igAGMgewIkgmDSvy
44O9I6BicoOWDheQcRB1opBp6mDeEeKQbh8v4M13QGXtzZKIMsbpIAQ+qPjOqkFJ
uCwc+/bpQY+pvieqJo2pJ2r5/eGtjAfw64BMY5jFfhmtfn3IO6EkrbQQSw1ivNaz
y7UwSQu4t2/8DrPSyr0Eqd3X0HXyVDmsT1Z6gZcp3/Xbz1wLHxnv9JsL0CK4ui69
/GGmubjAis54KjrpObTWRioBFSbJ5mnk2XlNTDPsFIBUbux/6nwGm6SoSgEKNDy2
QBjvt+OJ7EZds15JsPXnwG/peeSnoaxATZFJUbD5zoyJSXDYokyn2ORiqjyDNT6d
1hvgijKSlbrBVM2+NWmyMb+8IU2jl76QCzleob+e8L2nNxK5CMra76bJCJxp1Tt9
UnD/Sp8Xhel+HJZvnsEvJIC64fQmZT+Lc+trDpwmNRfyV8ognk9Vr/YapRqk0mLm
q9ZYom016CBMkOJ+RZJAtV4WhyHKQTvZ01CEumHyd52wFk4yh81Ou095i6OZGSyN
BidfB8K1X/8RTRTR1IaLEmvApBUP6+D2p5H/u+KcBhjMjyB6SSo5GkHyv7f8meRd
eyIog7HqHr8xoCoxPOxUCNcXfBrYjrTZunjtuD+Ou0LoyWiksDW3Bdn39/J7jPSK
IT8flvRMHPzcrsk5PtPtiQnizjVaZy71QsKetEFCrSIG14LOSAIepjiCK2DiE7FV
MQcpHSnITYAY6gMqYpTTx0U9TgUpTxTF/HGMDeISUOLoyakGipwr3nMIxYunYLFD
khfcLmp7pUsu7275NTu3mOJL1S5aqN3oSCu4p8/lP29XPTt+e6NhU22DEvH79jvy
OJS5g4Ri60ExGU4JPROWdluQDW2DVnf+ZUF4Xv1Drzje514BehYT9Bet5fFgXm3i
OWDbPGYw0Bc4pXTJWm7qhHC8OydGmPsDSvWGLKablBIhMXwfi3ilTjgwWL9VY/Rr
zUvWt8OvVpJN+AAFc3vsJfax8KmyzRw8ULaHFbqYDAqaDnGppfa9pguXrwzz/j2g
si8BeXcQjO0vjK8m/WtUnN5dBGWi7pIrpa5qSmwsbMRTwZ/5AK/jeZI/YgJ03L+F
RDnNQPVjJYSse3/5oLs/Jou6HjB0UYi+NC3t6XbsdMr4t9xedwZO5ENFq+4+VFIs
bN5jV7rmGd51ZvsOXAhgntVCjD0uQKSGdzwFaZAlwDmSXjXJBLywTDm+ReoESSt/
M6Tok9o0o0UDNrGFDfdgguaVQyx9BsG6ctyJzJgAXtPlMxoGgtCJKjBZ+84ub2v9
C/BFD2CLEO+JfI6hvxZXfuEQM/CP6El89vQj2BjvQAJiw3+U9xuMR8eVYrAfg1FK
TZXFEFhxLAqZ/+3cGbh5WIZeH3uNGxAq6hY8X2KNUCdauaxbhhJTq4Zd18xrEkP+
L3XMgDUx2v066Xqmff2x/ce0pZF5wBLUK+MxgjOZvxkq6TFWvqKGV+AU3/0c2vV6
14CAE1jUYAls0QUuksHCNMfL8llHmprg1vLFsxTYk037uD4R0YbY4TxH5llxpXRB
bDo8migHx3ObIqPxMsLfukFTFSZrJnMUvEThlBXDGRm0Dg1FrXGc1PqjV+tTWqKV
m3IXD10uSOx6dcvBJfoWSoelLSGqRRFPkSzpEKmYSf3JYSS3xq0AXTv7jIiksC46
4YLZnl8vuvqSS4mWATddME7twopgX0vA7pa/jhJ3dJq5QZHuyHdYp2b2MYuQkSo5
4DHHB9PPRDpzErhOxOmAtdzP0LmDoboYbEo6rQ2OY4x0vdJzLouoizwiBx0jtSUB
zEOehgt4eCj/QQP0vX1m9Bkbch8ir/t86S86luib3jkggzT12x38vC3/DQJgzZQl
I4ezry2QQvA8PbAkiLN9nauAYNx/movotAbE2KkyhAd+zZTxOFv6h/lK5goyabIO
JCaFG7WEPdVX/klK8jDuIFtqii+O4dVOzjFdBpKDZ8uochG3oldIPiJi+8z8Fl8Q
BbI9x8eP9ki/lIfRb+0ywvHm/cLv3wr26t/xO/82N04kEoveTNG8piBZMIWY+rsa
VTqKbavfldEortU7pUON5g8i+e5b0DzSeOnc6ifbW9vFE7RDlzjXITD9eSIOapOJ
BmbNd3lIxqnbVXik9ce99ZzCC47DIQjWbCkQvoJfFDxzBYgeApXqlqMKVYwUh4Ru
ty+s4vANtEXFS3OXrG8MU0rCvu5697bUKEI1/CkaBwbFQRhJ/Q7AM1zz9VbLmZdM
i0aYuZ9QlX9VhZmiVplmD8FijclHGGmSScI2anCXP6tHnRBKm9cVXbMHKD13+M8g
iQsgiP4WYh2TsQxCwefzu2TUes9BTGUcftHa+vnH090+PH/8JdNg3dJieL2lGFod
KeBtHTkgFimdwPPJWsMb+vn5snjShQcDwirlJO5rjZifptvh+pHKrSwThhBXi8N5
tkwXwwci/0Q+1PB3OsfkA3TSkMyov/8d+cWEwSTgIJC7B+UkuYQpbXaJLGtIT6/c
C+QiMdSmL0q7lXqTC6zE4LpDjptU12uyxZFdYTn3pXMpBr26YM1Byx+/6krRf4Ae
tDBQ5qerz5fR46ihR0OSe45ky+H8ZdFIWZhzksaAdR24+htD8ZiLmdcXTN2BJRcO
sTA9B4G7q8eaxaOSxWkxYYpIS/8w/6dK8xNQxNsMU0s+c73MdXfkjk4v7nBruv/E
19e+MI3QsuHkd1wodGgNPxg/dyrxp+i9gsPZdE1nFVVxHSjybVqwyoOUMe4jvvCr
xgyyOsR/wRTMjglMOO5nUtDXZFgb62dbVHxy1HYcT8/e+8Ya//pkFgT5Vqyky8ld
aD62uL1upqspNbVCIXA333UIUejVA60ldqSmU+Hm40PCinNpq1sG+cQCKkmCh9aY
fhHisF/S27g6qStQHStOYMFt/0fdZshJ4aUO+f/9rMrEuMrCuKmh1O+MJhX7dDHA
+jRQ+8+AL76IYucAcvZTD8Q4zR1mb6JH+k8VGVpAccM3/c9AI3YjcrqR/51fKk4v
jwfJo7MbbGOrSkjXzJ5xGZvqeFBwI8RIT2R6lfeQa1bGvjxKt7iAD5P1gqsv/brc
Y38WNheD7lSP0d/0OhrRJSVkQw5Lb0fqSn/pIIjua3Oh+mmXcuzXa10RjEm/1eqx
z/ZyPhWs49GPGYQTJ0/Yn3U8PCXXmcaDpvT8zIBbbHAdHBtaF4Xk6gEtjqU3Dy+v
FPt3bpiJ6iiJfXDP8B3Xqf0shDQkNSHlQqh+IYNNwTyGEtavAG59N+nnKR+0R1gA
vY7B8JbzFLRCj6MuillWo7/BEiKumGwoFXA3sRyUjGAV4YCvLsISMfJM4P6uuT1c
O9aW+kwsR++w2Q4H9gt7Biou8+IY2FTzaLYAGz+21aGBVArXk5ufaOIqyxWntk1W
NrTUXg1S6HirRtUdE5DJjSvCmPTu+acLSNU42eINkeC9P1w4QNh5tFOLi+yimku+
1Rg059l8jdnTXof8r6FSv5vZjTSjL5OtSglUw+6fiCKDMGxgKhD7/CNMDBaXBumB
junspR8bIG2hzC07WgQ1gfiuaCrbycLW/A7r20CugUpwHmAGHnTyg1ELK2yQzU0t
qGzU7BjKezvnt41ZJkb3WQ5aaEADEmaoT669ysUJWxjAVHPdrvH8XBQ8j3Y1Cv4Y
xuXpXBQuBrHKmPpVvGEFQmJwuXlt7QVD2dQLDPdAzfGYKimr9LQ/Kr3JF1Tb3tKt
EAzZ7J+Z5gieitMtzolhqG/AMdFL5hmZWPlmTKdA0UJKtvoeLtg55ugL3lUxW9Zo
OOJbcDpqkDQ3wqpQXM0Wjq38hDON+WVo/HqkhoMwUsZM8MSYW9uA605FpOAfEUsx
3qF5z5wZdECFxweojnR6D5UCZLQKV/2us6b7bTAQdmZIGDrhYmKxP76GrC+/BpvI
Nd3QVYfBQ4tSMGWcxXBH9J+C74QstGMZvJ4/24FCrN87Yuwp7+2TwmnR/rDmHmQH
w6D5LTPHbQPHlJLp1WiITknLOC+Aj97yDlmSf2G/R818ThQDJK52ufm5gqsRMQCe
4S6Qy9w5ZOYhEprpgmRuGPgna6nGFJtckUZRgVp/eQy6143EdTX3ZMyT7NlT1MGE
/ZFSQ7etYtpSTqLcegKSza7Zmvwf2q7UIBvL4YUkpM6AFI5ZPsHXXbuRQMSxHIq5
6i2HFbFGI5jX6AeoA4Qz84Wrs9Vk7fjF5i1+WgpeXkq1eWJav2RqOu13iBMLlhiM
0MalWXv5tmIJvWyKy9ql2TWsMIsDlKniyhVfqLI7PFAFm7segLkg8DSobytGCA+a
/b7DW3SQ3frfOR91gVTqlmM0+9MF2PIdGZC+EnNOwXnUlJa8YMQSYcbwluwL/zgh
cMKNxrpyRLzw3jDvSBx1LDxKnNv8rUXGEqQug2AU8xtWiJqw1pR+myGL8YdgDb8O
CiPnE247eMyQ4gGt2SvAAY9t9f18JnSNh/h57QKYYZ9xPYdn5WMCJUrCvouDbL6b
X/j2fT09IVo6k2e/hRrkvM8PVvQDNS6zDbIIStg/LVy13N/JK+cSTjaLiQ24/x4g
4vqiE4TpnnZ2sbvw+S4HLXmra8IEf7zlXLD1tzxECr/7OX0M+iYrMoVQDAXeDD8U
JZBPhrFWYQROx2W2AZVTdV8wOuVt53gc9TbCN9pwYP3juacV+DPvrUeBsEaCvGWO
ezBWL09T/I+KASOatYMr8BAugVin4GCfk24+69C2McIC00t01qPl3UBJKKhSo8EP
tPasq3d8ZaGGDC6IenzTEFEW4Mg7afeVLF+cABjrlMOVEnDWJDH61m69T/+HmPoF
7dfvt9ffpkNVbu1UBcDrWkSPNE3Avi8In4mcH8ROFlYrZmadse5H7BkyBFAhdhGB
WAJpTLteKGB0v16RNsvYQ0X0bClK8pA4hNpS4Z0Og3gCiEcIqaFeTNRKipkS8TMV
RU09/sMxODs3AMKwDIemv7NaIckQzpc8ztzDHWn+gvwoHhq7DAakTseN4YDYtL8V
S0d04P/oAL4R6nZUGcrTuCs1HoDkGPr3w966js0BcbR2j4+VBhIUHSRCmWnL9Q+S
11E5aYoy3tiS530IbauNNEUZ2VYaGy/eyKyMIJg1wF978dP3b1fWaY/dip8l68K4
qutyQVGZYOLRUgq0NvqB8VfjEwwMjrUxqmMPzp0grCrHykdT/l+nrHc4PpPe3dIM
GlIFkyfz+ev4EPQF7biwNg8KheTiCX9Cdf3QSxX9OPOGSnzZf0X7Ma1NlKklZgsh
xPFDyEPrxNEXRV6eVf2kXz8zFHkEmSIZkKfKgw3zoHuOb9PdxEtUz1XRHLSMbRPp
EhBcWWHcuGg8o427g6IAHLqPufXTJs91O5Kp1BFudk8Tb+EXILINaYepQU5msATb
s6PsedMGbruxg4ZlY+R6zWhvcdVJxjA9inTfZxIdIkJqvH82Ri42JqK5GVWIAlKO
Ph/iRnjBbmBdT+Bk4y2QVgCKn4L293syLQTeywfdfrHu4DctfbcVSJmYKgvG7Nwu
wGjuyFNPNvT7ne7LOuXxnw6A/bRogt+OS1IBlpyKPD4ERFwg/hP7d6St3tOo2znX
IS7l5g1CxKghcQJ2ywmTVj6GTVZUCjo1vSrkxwk1cuXOW2ODBrfyjnrLDm9Hh9MU
ziAjoymOIhUaynV/077hXLCLProysx63rwUZpj+BYhBs1KhxphnZoWko3pCUH5CH
PfhAo5oxjfuSgGAcjnp7cVFKn4GMQyKk0K0BI6521hfg27gbO6E1eIKSFnJiyv+X
enN0Px5/xEMGKjH6TeBVO0SFxn4P8Z7Or5gWbraKiQRNnhmQvDO37R9kznXArFYC
Rjk2wm45cXBYagZddR+CfiGmFEKMQpOn7+E6rvObs4/cMmaVo7aaVD8LEqbMuiuF
94vY8j0xA69+WeGUNZJ7WMgJjIslyPS2F++lbru8pMc7Y/za4ScllfHgOSjc+QbH
CKQ5ZsN5yDuaw4i87ZpTq2ULktpCQly3mP3ui8qMMUzVVLbnkbgFBv3EylBhI4x6
C6LhR1bZFCYQxFT1/dRZnSrJhbXEbQDV1gpE+N3KXqL7tm8ztOhf1N26dY+OH7De
tGXzckPD4KmUmH+hzQ3O8uo1sWJzvJZ6RQZ9jvFgz2Vuuo9RH5ff/URvk5TnuUXh
fyT6sMtqiC5lX/socr9ictqqKEzAtOzm4bOVxnQr4QZbZLlLpgD5R1nUFAZjMGzv
tILJ43OdGNGHZldZqOIw/e9m2YiMzLgKaDuM1hmkrKcMPw1LGn0JYalpslr5H1G+
/S5uKDxB4lrMFhTDVkozuH1JJL9U+B42xup0xRe7F7LbyE+FcmzA/2MSGGGW4/1U
0pxectfSPD5uTb1gIJmWT05NfL/CaLhtvn7novi2ssZiGBjg62zvZSRcIZuXjrPQ
2pcFb23ZVXnR0Dnq/FRWmGndO9DbwWaPiBEPgm7y2sMRw1Fx2msdIwoMek48MbMR
VoJPEg1e/OBJiEcq/BrxCuzt28B2sSj9t6y0sMcC3iT6WUR+4rzEAjPuT24x/KBc
b1KJ2vIrXnH4vv2nSEq92D3GxJKmvBrts8nqbwJv3SOaHe2T933xjvO7mXxiyUSf
dVuEC42pj/Adhhd+Ze8e2LdsoF2Zyx/e3a3hlPbZeeqZLKiWds7y/PSs6ZWKWakv
nOJ4z/IhUMal9Hg2QxRqicPfvaYJInjdeu1ymB2frZaWdejFQwyA2ieKH2Ga3r3Z
S2xxq4tcbWX90QcLXsquavb0LvUXg0/mJeZ6HiBQPDfknaYFrOg9hSX+7V3PRsjT
Kud6lS5nMZVITZOzm7pDQ/wy1ip6k+N9T3xTYciNQYGWFFTVFU5IT6Nu+3begiXk
gWlIu9Gxdo0rsSO12Zm1rDFzti0aTiB+m2WSUPQueoy9P1vdy43o8EqNy1wjcjqd
fANyshABcmgh0A8deWtg8HzjdXtw4ZzNqwb8WxfZJz5Nqe96OZgLj0/Y47yfh8Lx
HZ9K7W9JM0Qd1ZCUSCWM7zv7nSJFM2gmAhvxyTIkbwuPaT+LcRqi0IHFiEJlE+lf
mgqkOVRzdykrpt0+m0YAbhY6cQzAnT4keYdfAii58oMo0O3q+BUQvQUFqSMV1C3o
qNYjrSLluNCs0PNAl0gyveM/uL7azlo3ogqAaMxkdUZfinTokpdhYjhFf8nPDws0
qZUhiw5XorObftjaVg5qjnFhRwLg4HRLlvpGT/H7/ByFyg6wIEnzYL58BtDwwDa4
P6uKsFJ3+hwP4KxXGrndvv1GCtOhjQfgQFFMYN01ccvZ2+ueLz572+Mm2PVE+rzt
eaaTkEBGHFLaEAHLaWZBb/PqQaoxBk9nN22kCKLAkaWqtEPnIlvk4Ubb6b3kU4ZP
O8ZhKO4atnb3aLxWR+FM24T89+mE1JBUlmvR5aXFIdkXyhvFCBTnNSqPKRJDD08v
v+X5dGSgiaXOeLw1R60nFVvDF+AAKItwGKQFlPDB++fXVjpAt4nWnucmD3Yn3DL0
dUjoJvnl00PCfmqdfV4Fog48zpmtOXxriZIEduFrvFSo+MwN3wHYeG23nJNlAKdu
ArN4tN5ANCL/J4Feh4/JI50zo7Ved9eo6NvLL09DpMm2Guf5R6u4GeN705hXyCsh
HH8mjbFTviY3x5seT66D5GjYpvlKoYGFuGlnSZT55TkrWF/Nb/RJbfQiXcMyJ0/u
xTogvkNVOIm9xYUpS/6XgJ+YS7ynyERDohDmM1q9hMYy94a2hgbyAOF8phIfjiH3
SR1u6JKOzWy9bKIROFwiiqAdqt8etqZfyGKt9/VgRHPb0Hr7F17kl1w1QyNTJY6o
YZbVIvuVC2uSv9dHjz7Wj3+O2d/iuvVA69U/YDYb2vczysHb5Ss9RxjA8EKONtRK
gciq1pd4mCbLtICLOtPSXzjQyT2aE4kc6+sFq675D6YO6iyb94X/OPdHADzGdmdP
5AdWNxQG2GinbDEsVxOuHl0fyGJb+SIj/AhKEMm9/fO0FNRTqygjNHnpjtQ/gxX8
85v+LiwyotV08aq4T7QEa8r4QQVSpukwv1NN8WYVfYi03J3JgPUc+Wh12/Oj3UOC
v2VkmYmwXgMxH6cQb7sDRuIDiaZ52PeXWTcCH5fjb6hUyG9K8vIHhYU+fSLoyFIg
Ld3r4zf18XLsItiZ74r+3pTonahcpma9B63s/9UhzGBjtqoWJyNn1ZxMTFY29562
Q/9w0Km1CT+SnFEYY6qHM8AvefDHfe8vuVDRY6KNPrx6fYHBN8FKQBnSiMj4o73X
Ji1eLWS97RZRgbDv9SZQW29Flpks2qzXz9ewq1en6Y/kUA4JP0kdrwtHiaj+7aYs
4b/G1fPs3omkZtnC6g56guBcsL7PqYk5paRU+pVHOwxjxB9JD3eRhNJZCza8gvE4
UWhDjs5B/lX6Mt4iNRno09r2H+nC33wUJRLY2EpvNU/vZGasitZEV+Ngz716co3w
YhTrKKCpfjjxKui1YXOeQm0tLkblxbrcMM2GpY5/TdzvJicru8koJBRfJpzAhLgz
LqZqibZu0CJUg6nMbTOXuFfTzXwzmK0vtgUtXoLAhG9au7fgPG/38R8LdNx2utE+
EEuoDM/mlaXaMKZDDioy5H0Jcard/o2oPOZrXMeyMRAIdJGDj4RXDGqkvBUrJbWS
9PzjrBiEYcB+A1OgG3T+GRW3Meh5+BXteVsvBQz0ufuTA+Vkd0g8JTXtcJ7YSNMa
p5dQJpa5TU3Jjn0EqNd9rWWF5LQ2Jfobvj/fNXoOHdh55Ilu0ix4WObq3NH6mxqj
z3WPdhcnOVKiuwzWFlaVONIyX/MEf95ld630Kdc2IS5CCSb2Pje0XUdbBlaODyDm
u3iYJZ0eNldCgUzn6eNxYVxlRJbPf9R1awM5mqwslMlur5zKxLvD7Aq6ISQdoPxW
4ta+eoRfXGmz9AbmHeshHjVURosdu1hLo9PwoYgL/vU0jvUrJtQbTP4ngszDwzjk
DXEm5dryGYVD3jcm6F/hZ1UQp7oo563ySSO4dpF4HuqAHUwmJLqmuUIHYzYDLZqE
bF3QE/pJhhZKw5s6yN4bHAtSQaqDzEM/JF66Qz4zm6dQpHPn7WpCR/hj8TUzVX6y
J34o3zbuGdPCWSuK7nlon0CMuX15XZQMGob+ijdQ/59gcljJdb/ZJVCWIAUaMuwU
POwMH3M0Dx8z0l9FjLCGxPXa5q0QXKHKHPJjX32YySKvzvyvZLwM8NCfU3/1p7cM
HWZP4HJI5/3bmAUahqCR6qbcuEjbEeC212J1dI8xbsoG2dxFbce6l0SHaPTLinhN
bLOq+crWpsEvALhOqFoiN1aPWM9xxUR/+t0J/XplSnkx3EjLRWBO88x4SJNyK6y7
Fnem5NYr8frWHTOTT1ZsjqvOFn4Yfnq2LuEy2X8QaWpM9dVaY15ZrnxvtegHGcPZ
TrR+3H5GUAO3vMHkzVsjI5HA/VVR6BYmVoNj69cYHljz6cTupmmY/meTgqsRS0by
rhSLGevOXa5VNdnnRU7TqYXhiv5d9HjwBPUDMT2HHG1OSyP96Ryq71pzInR+/HAJ
owSk0ujDRpEur4D+sSXJEP2ThtXLjo50rFvq6NuT6HY4bb82cjofkzOdtjLpifAr
SXfPfe4dQSh7oJBgF87HqitiIT2ikFYAr++C8JbKa8/lLmbUwHdJFFAEx1Od7zW2
2rkCKXoty+u217XXVyGgJy/h8iOHXi1kGuuPg54isic05hkrX120VuCbdBWhZLJI
Z5IKfW7BpkyCYSAZ5tp56nTLEYTIrKO1YJbMIT7s7LQSC3EpNdd8GrfFF89S+mwf
Th0Miv2A+jiwmmP147x9bOA0YXCDXeiq3Nfgg3GwsyhXMdjl8+r3wCTahac6wFqf
JAer7icdHMpCRvo5+RLZ4Nyf+JkAkNevalnQaH7GwpvWMXPnylGE1SrLWeW7dKwM
qLwbfP9x8crhelcnXP1CwtGYeEr1LpApW9o5bi2qzSw=
`protect END_PROTECTED
