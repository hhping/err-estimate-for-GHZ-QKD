`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M/gLyJXDQsmCkqRkFlCteDfpPT2lv/vgTRaVLiPC2I69Q69q9tKbH9cvTX0iQFnb
4EIVuZ2S0FPTrc01a3csOvpyFHhdq5iq7l/OywIRZjEnqu8Wwkbrnu7RgKJdgfXN
jURzE5TkxfTBas0saJxaWRulzez/H52Csh2eU/l1/tFztoif5SAK8EPm06AYwOPs
B2SzO1ykPPTZUbYKdXf+j2072x3MAZ7WpG7hLLWl+HGJkWnuAEpsMEyDyRQUWbGX
0IPLmNOXhD1X5eD/cj3K/35vIMbbUvhBL7W32EuP92g94HUUWIlrwR1FMcFSDg+n
04zxImYnv9VHQxLfEvyeSeU+WNdF+wbXx9svxI8svum8itLIBPjKskhGRT9LytBQ
LcDFKlbYIzMUVQMUPymEJsr2HyI2xi085/nPrt2zezsiDeEn1qcNDbGBoYo9tgpv
xtneNBBthlVN1coz3nHm4ro1R3qGzAvDWJO47rQ/495xJFArCPnLY2cDQvTFOJVt
qF8BdptBQWtVxeZI01CinYEDCAD91z/hOiEQFiRVtJxjRc6DbLCpNUi5kgkQdbnW
Ok0R93Q9Ma0pRjmvNRFqwaiwA7iWWOXKv2adhnt7rlXvpM72t/rAy+9dmySqmEEF
fsnw+4qK0fChTs6GJyxiGOeFk1fRUsLABFSpKJWvwbt13TAsJqTEBLK6/kMjqwrs
R9MAlxV2exz16mXszZYvE7mc6hdrU846UYeF3154RLI/AWb4nAMhRgFWdWgQs+XC
ZV2DwtMSXuNyHJqWy2aLMIe72vh/iblM3uvgJtYkaJ4mkPswMwRcD8pPnJnZREF8
TAQbB7minbxu/ahgVQX94Tt1I99vrKfzqTx33LW8hOZ38Lhlb/ocRlyvnwOTl0hQ
vaqAKjSfaBGP8O9WqbEMPFEiy/kDx7etzEET3JiB4pOe+GgRyEz0YXt2huR5QNil
8KnLtQXKyal7JsrjLYT47+//yHCtKI30Nj2UnExCPt/T2TJkYn382aa7qFsLK43T
iBjS9aNWWFvF4WG5fxYfpP9jft/YW8PEwbE+yuAZQazqDZ2QOqZlwIj62CXyRiYj
gvfGGVN/XZF+7zxNpQ/q8YOP/p246rAj6QtDouU2BX4i0NXh+FOaPsDszYUAGemo
uKie0sH+eBsVoN5LpEHtNPoGDP4S8ZnmWQMDQ35CI8tTRDXCsux3ulhsv2CVWWVl
nKdzWnthzDD7D6TjYbjkejbEf3P+WyiJGipMvQzoUath1N9vL4BwAV/nIP7dHeEa
nktUAkUbQPrk2pqXyV3RUOzNBxjxLcMCs6s83k+bfUJN9qmHW3G37v9KsXe6anf/
3IYyPTpQJPqQfYQkgjw1oslO77qlape/X0v1w9scqv3Bdc1byqCV0vQhQoBbtgAI
VY85q1d4C/MERCXd1UozIAnZTgtH48C2CCSedh4ou1hnCb9uZw5JScQNYWZBGcVx
lxrWzzD3xGXlvjtkV59g4/R336aZejWNV9heFrLMnz7Mhx5O6Dz0VO1xFmYk3FBV
C+Ou2fuL6jkGBXELV+bRPHM054zgnee11OuG/guq/pdRoLagh/PP2cDgZBMmFXrP
fIFB2PV7xY+KtDrQD0zNBkmXDM4eQbBLbkSUZQTtbOFJEy82rnBdKM6BcHgdTbXD
P4Kx6RxRbgZXtLgHcKLo5GablcwBODDwqioPwAX6b6fAeNFnMMVBVyxcRnpK0inW
YHIFCYOMgZsbRCYyoYWoIj21Kg4erD286N6CTs1aodkY+7OPBMoGOwQD7ep4Yfl9
tvjCmSO01wWc1k/EWYYzFGuaJzZGNgqvWrMB0CniuIuvPHQo8L0t1lmczHnXNYwK
rA3KWkEVNYorDW7HqRUg6h7TcZmhmjzXGX7fUIFZ1hUJz0pKaoFPWjnrPILXQc5u
S+R4w0zoHKt5QcjzVVDuWvh7stbb1MfXFI/6U13zNww3OXf2hE8uxdHHVOs/Hzig
KrIXrKMrUKSkqjhKhB1RrX53RaKpVPs7RrNkRX5DD0e4G0RlL+44HN+wkJT75Kfr
SdxHUmU+Oq5OGokz9BTWVJHrQChcp7OMgY179FbChGCT6QsRn5cK5Ujidho4tC8U
9G3iCucR/W9EvnwMxrhaUyje/f+wpXlEEC6jVzaFCwEyrVwfFG6A2rbpNhTLFCyB
buTXSUwYyHk9QIVVnP7+S/nliZkIFOhSg1kXia5qaj6y3zib7JxkEoFvq6W9HIt0
gfZVDmK40CT+OesPzEVY7sXrxeLV+T+m56rtYvwKQmjtoacji/xwaPGnZrchyen/
1ZqLMysxn2K5M0USxPdByIqQloGV/AfXyPm8cQ4Cbx7YbOP0QkfzC67vs9Y9ZjwD
JBx2amqn1vFWEc4KDdFP9TkNmaCBSBIWsCcyMA6a5E5Xr50YVh0es8xT9l3Dtxhm
4DRi8Taacj0GcVOOqzPpcdXiq2sREVvDAV1YTsXhJs1mfbDxmSXFR2ZxwsmuAayq
d6IV42B/NU2E1LAZkS4TFuPipEI/4sp/npqUGoMnx2zx/Z2VoUQXaOTD7yFXlkKl
GLgj/+fELVa4hgKLSXtByPlpQLyorqOJIkAMWicc58e8Gsx8N7YJYAf1T9cDYaMn
LXmwR5ZU4UGcT8Ko5ZIWfCae+8rkDD2r2goBnzOkLOHon/IX6+Ld2PnuRB5tClK0
uvFwXUONs5gyPWHKHV9yirtDjj+wqXgpOgJE2w3o6sEn8G+NETtuW2yhdq2HrmmX
PeexfUpDm55yR1wFYFf5sT/bVEsxlpiDVK1JePNeDpe7G9sXOKCdbsYmQnh1s0yt
lF+Ed+FMKpvdpljQ42sHytWQ3HTLTexEH+WPl0jKkoEveRRhdVcfRVWR0nIlWfCo
EB6no9UY45J3raYsl5iUVuYG2kjDEuTcCmYUuX20URG8cVawqt1TcCfPuh06nMz+
/Dg9YlqYCkpgHdoJfSDuQS6t+gcQagvmH33QbWjRLZEeP8czyoIhVID2MUiKXnCK
9Q1pgwktgO8Lh3PdCeiMEPB/aHLAGyQ1j83LA/cvx/tf2ShEbfJetSolahKP0H65
9k2kITTWOSaXf21kXYnn5LxR3EDs9qM/E79nVLn4BBrH48kYevSqG6hiSAJwNYQs
luNu6Wv4skfkW/2uRDnIB+GYqmSYcQX8vBZRHPANkefOjCVvrQYrMPAC/DleuqKk
47ba8RLqgVBNk8JW9sglxYeyJDTdQW7Mg/1550eMZrkzNavGG5JV6YF5nLAKhB92
N0raqIq3NwIOeHoF6j0k9wYZIVnDndVf8P5urDVj7Uc0VHmxQHBkZmNoxJYrfJ+x
X9ldn9k75XdzWGR9tZcJCxjzaPxBvDGYf7dsarM7SLl0vJD3bDd/GvxdkuC8tYev
1AAdXA6doKoxy6wL++ny3ADkiPA+HOjcVwWsGbpeidbMcdWf1eOmSapDm/ihl9MX
98Kcj3fAJB4KW1vgytFhy/JiFsKveweztMYZIsuwycgVHsg17mD6IUcnzRbwCCQU
2SfGWjAnyV2dgAmHTYufldj8lBraLrEeKh4hrUvNiVMRt1fD1OXjeMgtFfKQ9x0D
zHn+sX8WdtlOvz1GfHBa3WXfELzlwkfmZ0RXHr08xcnpibvEn0NfqhK6QELzU57r
zJBrpjZ1zZez2H+d8qYL41oJOMGnhFEkXD2GU3SpIpT0GE3cQL8fpEj/wVGcfFI6
W87yD/zSe1BqfhVWQpRX3CaPcgpAWu9tIUFU/HnetRZxHM/lsAmmmhbSH/UF0ovI
tw1dspCE1GXiSmV3XQaZjg5GmTbrsRdrD8ANc/KdeSOZn5VDl/KVSQL7D6MXaw6z
241uC4mVWBOzNjY7gNmRIgDxluKgFRZaeLPjHAdxKlim5E41qlV3xBb+fyY1iLt8
Q1WusToJIAVbeR5qyLYlgpJDFqPYHv5eREPC5xysgqsq71jucMXJtjy/qWttRvUA
wOx8lY0RSkKyDFdz68RuIohUNrlRb5C7BCopcrhqBPOBUf+15rhu8VYAFS6vYmUC
6hRzBrhdsM2R1pphJdTweTRKzqawdu4D+5WHk5kDtBXfzLPLZhUSgc0Ri/xaHXi5
0QPQrybN7+Dmdt9hptEQAW5AxEXSLz8GOvjAEua/hKpGLAvlIZUnulHS1BjuJMr0
lzOCsFtgbNwxlJutvu1KuLZDrGyYhKuNsO2YNDZHJ9Q+QTBkAF8FFYNwZFGLNBvf
zVd5gupWtkx1YClVV/vVOi38ueKQN/HPbMjEH1d1ABHhkSOWKPGtYKUzO5Dq6lMq
lWj9h0hK5PTD/sGjkuGjnIcje6zJ4G4wUdLbM4r0fsu4BeESjdwDYKwN9gkdUirM
KqgsXQ7VkGW9UISPdPbqPCvMVs/rtV/lvcXTvzyfsk/he/tiPB3eAuotp2hC9mlU
u++ORVt+ZzcFE75ro9NSnq48jYPKrCW8LQUMaN3OtmqLg4Kyf+3jL2G+viRRgaYv
+iI7/LC7t98XSIjvv6oYqygpVO1gORMyuayb1TvQMqHiefd2kKj6re75EJ/NRO1W
E/IAP+HV6VyBSxtXlA0tofmgawNR2bJqb5GnIHOOGkXpQZWoEpaF1ZPErv9f7iys
4xQt8upW3tM9qhuGg929lZEcz1xIfJPLNnjeAGjPFJ+9nX/zpcu/Li1TtztT6v6a
i6WA2PEaAQXdWkT/Uotdy4ldszUSa2MB153byxc7b2JG3jx3nmTxo9JzaHdayiQq
f9nzQrG/D/sgvWeMUzcK6CrX/Td9D8dorohhZPr5SABTO8NGTXAvF4OCuzoubnno
N1j2BKeCbbJ4PK1Ehhp0AaMm3dRNRUSzVFxxlhRi/LAONaNkDYUNfzHIJr3iB5a1
JOqjyb+XflpymKOT4TjbXQxa1FTzUz7Hts/Z98x/LurzNr+5jSAr+dKpFpiMYtt+
Qo7C3R3LinyDHwYaDIAGF8ARuKG6cvzeEaU8+Xom3VQiqqFi2kTVtziFaM7/9EQJ
A93/SueNBNZhx4pqkbkkq6BY2KiQWGyQSWEtPg6zJWnk94hNY1IqnmUp4U7LxnOi
90NeZDZvDRX3oBdXf8aJWh8GMR4sMjHlOIj0BLsnAb72tUYjxE3556YPvZTMj1en
dvXxlTYS8qaYZHZKen74F9FQnGR9HWreGbNgJ48jUVFkDXqEnfuWYbAOEiKihCv8
RdlyxI8SraUm9lTiXK1VmRiywPHTOw1nbqePuns3hKpEGY+uFA4j4cH6yx5bgj9H
+9njTP3sZ2dNYEsSt6drghWFP3uzKpWrZCAuRjfYpYmfz0fccw3vgWLYg2reP70a
JnLfZ63QsPuLWstqc+Y9rsbU9Hu6R5fxXdFMnz+thPVhVFT8bzMwE1aRWWV7wDxi
P4U0WbdTa4GfUHWVhk79+GcbZSiVi8PxN4uKKiJAUSY9RYJIUr1jBK48QKSEGHto
ulsX1MtTIvjk+D2rbzHRoKisXaaunXv/4NgGgIc6iBHT1gYZZc5q9NpNkB8FhaGw
owtWIIn3w00wfTDLm6SKjKzkE1h2kLWXeTcygMnpeiV/O9OjOKdNfYffJQv4C+HO
MiKQQldXT0UZ79EWEZx7PyC8cwR2JtBRIsa2IjG4TwRn11bOHRrwO/HYpxEFITMf
15rxX7b6RXp/rudG2P2zF1twpsENqfCBqFtaEuZjIMv8IBlxzk+YxRnGEp5iTd5+
nFmHbyp37a/IrQnha4psk1qWPqGCaC7+U9EmVMxq63c14NoseDaRBDy6ZIauyw9B
P9k3GIghmi48GJBs7VQ35vNvtDxlpVvFkBCVchRB/GuSL3YYVSI1ELmnlyoscCma
KijxjLBSTWLPqc6/R8z45uFh1MoL59GInDFJJv+WRQ/RKDKulD4O36Z/ttA3qNLk
LciJkNrFASozQ9/iBE1fT7/vX32Z3O4Fqob5vxaugEWSv0FtNRC3Yms7oc0ht8BS
jc1NORLyNxU/lrx4t+ahVkODutyupqdWd3IUtLI9m8s5f5UNiKlzoO0KUGEA4b8R
2iz6vgG5d/5q4Y6JvjiQxSpTNizfg/kHGnyR2SVL7W54gUw02r2FobMnfpWBCRQN
ksTixyNCx5GidFtjPROWg+e18iyviXkn21EL14U6PGAjn3OjOukz6owr1HJmRhVY
TM6y8KZhfvBaBbdIiDViA7yhD8RlsARpKWN8qqb8u424mNtYbqCaOu5zWTdnLpYC
uN/FTeDiuq2WZ/e9jruiuPNuNrCtMqJy0yKOMS7JBCsNyuJizE6z4M2th0+XWxf1
n61o+jMdvkw0yJ158OJi52XPmCtt4vt570XPy24BdLFR6rix5ON0JQVuMNQm2J46
Pyb/PECelB6vxXP0C/jwnmUPXdVo6B5yT8Oj4dKCnZrpyGoHj3xLpz1VB9mhpHaG
Ml0QWvKUl6xy+sgDGxhsGHzjKfTfqeRxZOwKG9BsrqTxpkCdcF8aRaDTOl1XiJgn
u0ORttMR1g6aPTTREr8KTATQid8h6Mze57hzM94K1l58S650MAa+1CClBpUOgjx+
QOPkVsh7QJqeXP6xqT1mZvwFlVMf5HdLP59cxZEFJbVk327KeZgclvqMwyRyI0ns
SghKaBRrDsYR5cbMsxkf4w12svlzqCgdC97wtpAMV6WiddjygvQeiPxhDx4FDa4D
dyoNdBHK6Lae/R/TboRQ54vfAGfcd3/Lb7+84Ipv38Y+jXl48ErF7QdNUeiGUoP6
4QzSFwJkuzfB9/6/ltV5ZwYQOga2PJLA/XPctCk0PhkpVE6nNIQAUv9IlsRZbacL
EM5lgwNHPGwedqYcilPwHX1XnFzzUzZOa/2aA2/Ei6uOJvBBWbnd/y25bjJZZ0Rz
Su4q/NT68xcZ+nsYIpz8FVx2c3FPcAokPuICMUTBjGVQdpa3RDH98Le/MdQcb+2i
ucvB2Z65tzMQ5VjyEM3MJF6FIxQrF+GyTAAVN49vXGeboJeW0ZzTE3bMOSWa8ntn
MdeirkoMfBtjNfKGzonj5XY4KwLedni1wmrEsj4dKPqSnbUJRuCoETxGh92mTQIf
5NcRiqs69ac5931jFteilVEizRqLmwbceR0EHmWesB2O+aUvAhS4jDh0eZicXdBB
sNht0IPO+7kxCEPWnetdirM9p23a8SBDmCjutv2A8VRxPmDQr2W9zM7gbko0KHMh
Eby9aBVBNuhrGRi6aUNnz+3YW4wBjYf4qcNM+gM0K+nTChL28sqy5lNegc+MB7wS
hyNVJi86bmNhkhR3qdpNpKwbjkqzrDaS7jAUmf7P6ZCf1jjlPbSxUjBVdLkgUjLm
MyZT2lcJ225udSTf7bMpJACNeSmYMf7wMpM1o3ceXDgqT90bW+OnozmMstt/Fyh/
v5jhNNlntRl/09zoU8SxWXYuRyftZGuQJUo8JCdYcog76JQRcdDsnVRFkGgll5+j
ZGEQRE3NttwjQjk8F3cFlBI1Cd5w41cxsQXrrveINqo2XLjgYAVn0Y+uuzkjn1KP
FpTebalotSFEtNcv8c5qKWyB7jP9+ZBXTl9p/rSyj2XU/yZbYoZcTciRaHiZsLYS
8TB4aKN53/to1Nq2MO23cKT2Tp1wYVKFTvHajhBuYOYw75ybUI5qfmS0K270mtRH
AOkJU0Wb3h+UvLOeFay0xxktgS4OhJ86VpgXvL5DfynwjoJXjlfFthicEX+FRvAD
jXZAmz31Tp0YRqaC12vqxmIbsMp6unANEywjbUcN4by4eWIYFCmyFy0x26J51W9C
7RbAcxsbgBjQ4Vs2ONmAx3kvnih+DfolRCFWbFuZvGmTvdbNKrc0sgjpNTdzdXRm
5G87fygzab1IeB2mvB3A92EHbLjdsnLnc6yp0Y/HVFqmQn9FUHG4ljo6p2K43yjX
PppOQEDw7gIHr5KxRqiRvCOf3dGDfcFzRIQedUembJW06UTozN/ThKlCgZfZI9S0
irqU9Amu4elei629LoqnZzIcNrMm3vbKs+A9keIZxirfZjVAjIFc9+VNEkhUR0R6
5vGM3yotSdy23OJD8avr20O6TZLFTWWGEqg5sAPAmyemR8gHP4cMA2X2hINR0tTw
FmW8xQxRAVjYVeuM6UPZjz9fUWCWzF0lcP1/tKrzkIl82mtHoh3U1uNXR4wsTSHR
eGUvOMB4swmu6refj5q7TqRH+X8vQ95IGs3BSCJav7g/1YC+YMg9pDQ6bg9ohAOu
qfNnJXZ3NtP5ytI/vYVm22y4PoeNsI3U7tmuQTZun7Icv2WuHx321J1DMETzryGz
E/VynZGR1YzVWQ9yUuf8Nm+RVPm2s1d7p2/KQ3XoWd5p7IEn57I1PUlZEzYYgjuy
HKBMWbJclVMHKxlI7vq/o3DK/mS5zm9lJUMVrzjK1hHOqtQggdcq/BdnKO0neQ3o
q55BKZGyBHaei78Rq0rU4YcwTj7W2Do5H2XIOU9bLXkUVZQC7IQ6ExN5Gvbr9OAZ
LRwY/w0GwjKuPMMuR+o8hnuuJ8PbmaqE0FmO9+BkA5eDyPhvMbcJwFgyNHZ+5S4r
iMTeV/cB0IVQ8hwO3CKjH604nYMbeld38/ACF7HCet0PtjWpodp2IEOXnd6430wa
mWjD2l9xVW/AeYg85//HZbd0KgKSRdNYOB690nbOy7plHLwnPHG4wI+Z42S+GNjZ
rDXU/6RbrYCw0XWD+LayK7r/cG8QTWwVhyt8QJvD91hHxRHY6taVD5sPJophivrP
Q3ynKv5NrHnC2H7cH+dQOSn+7c3MmQKxRaThIPeK+bU/v5UoV6/jrBP01AnP06/E
YaBsRZaDetxr2IXRYwb6vKmLYfDazDPi6i3M/f39LOC9RccHyNm2P+lUsGHxXiTo
qA48Nd0edXzmCDQRvxcH2GkS7hAXbbwpM6D3mD/rUxeTlNRNk+fheKWJASO8uiNH
qxEl4LBOjLC48QNK4GU+ky5hbz24qZ2P4/h4HTQ/552geXeBTz3NCfIV/WxXBS4V
2gspVsiQXHWmei/KVWmDNjQEU4Z48ms/faXjdVRBWO/iqS6iujrBFOc2g+Ko03SH
kqBtLeHM7CagG0EIwoe2qFwqpjG0rnqf8xef/6oYLvQ1wAf+qFFC+mFgv44E2g9X
ql5SRpRbdP5FiDVeGWyP6ioQYORagVCVPmkievHJzmbQZidQwrJx36ZYYFoECTTu
WtRrz/rpEQqBNBBgGlj6qyKia8K9YPJSDOMlm8HrMOIGKaI5Y2et4G2nS5HO/7Wy
u8EK3CB5XgIdXOpTuZKUzrWF834YJlOP7ux0s9XRW3lAnGGS+AaF+9cnTELEildZ
OpQMMAMID3UEBVUbnT/80lj4gbEhxmWEHtfdaSOXGLfySOqeBkNDhsM906vayRUP
7+yxIl7UpVP6s25nQEAVt+X+RwG3Uxg10Zc543818ZCtKzcHO7amu2eymKaYZXHX
pe5XI/G1iOsx9XdlJ0GrA2Df+QK+bSZ9vh2Ix0lR3dB8r3bRAPrBHONzVCLWMoyj
tgUOascB3HxFHOMN7A0uIi/udJ/nMo/Kp7qgZwx5siStqi41Myf/0CemlOahKHKQ
/3T36yFniPpuPHKAOaLdle7tFFrUAeFz0U0FJJlOhSZ+fqLGRLbiZ8gVozD69yOA
bgHY5h7NOeMGdA47TqlRfHZf3wX3zqyS9coK+woS2AwEQYmWQhQNev0ORk9igjnU
ts4qj/BnTXPJIvIdbf5Yhi48Aothcbd/ELxMJ7SLAlG7Pow0H/tEjsSrr0tC53Us
rXFiDmskyyGnk+Vm4XjfTTyZ0Q2710rK5VuAusD0d7srJlNNGq9jHvA7Jbw2W0MV
19Yemj6Z+Ikj1NHueiq2x2sTyLTEnqRH4fLoyirsSXGjTEyVdsq9iFepWdhrlABT
Bcfd1nPrLAIQsfAEQVs7Qh9WDHAg1IXr6cMJ14kNY+yAr6W1oZHwvvMWxnVZGI2a
553KC7GqxN603V5zwr3oB1O9vSLzualFHLxaM6WyKmAjUHNHev6EWKFuvckoniMz
psQzKGHRkyOgkAX7w85LbayzH+O8c5HczxskU68BMUWHDFtT4Kjb93RbGXHx+TUT
g4DPIkq3EZJ502Lfsq8GRbX7Xh8Plxrgovj1hLcRFVB/rM6cXO6Ct96c+1Bnp7+S
Os00ulZNrIgSJnkXOKfScXbRqnjcYYNOxtUPjAn7sHgCpE/xV4ysY9ktahxHsrPk
oOfaA8EAUItxdZ4RtAzd5Jcmm2SDG7nMDQulzFR/CONucXwlEpIyDV29erfkQBLN
qQdK4ZfjIx6xGFmfdnF+mbbxzB8vkCt9vXJhwXCPLEua6aD/pNzTgTqveWgAxo0V
WNV6BDxslWjV3HxF2JLQTwhbgYuIgsn4fcUZK8GThTH94c5iiIBA60DS5tKiHmiN
8vduYEFk6u9erlx7SY86Of+NVWeu+ZL8C2xuhgzMMObMpxda+lVI32GjOzkvFfd2
C84z55J5zi7O4RU/aAXaQbb15WEFz/9rcPDOZMw4pia4IeY+5o/clCEKpv8rOaMO
Vg1k8heMM4MINxuyanSA5taqpJwGFPB7FR0NN6g2HUICNXmG3VarRvGAkLLjzcPs
qNrU3VREQWitKbDlFWIdyvVqsP8SlYVcoFHtfBusA0WK9fK2ZbXrZDjca6j1CO8s
gqrX4E2T7sHwP4nMQN8rqyh0dmAl4XSE2mPoxr4CabqoTA+ySuuSS2BbGhyYsbvy
eU9XhmfJozUFds35TD4e78hJwZJcRf5v5twiBdhjhir//l1AYevt3aXqCa2ls0n8
ZFzOHw2wamzTFZsFQD8V3gZfSoOY/VC/dz3Rr3yU0R5FAUezTSF0Bxq1NBDoLzgO
9tgYhj0YgZREVztWarC0WA6Elt3qM9TfluhiZiareWRsw4W3fyUgrz/e368ryDP2
Jqk0R/7wLvyW3svqW4RZGBXbn2v1CuZMKoSSMZF124DIzteqOir1r6graKpu4n2T
r6ZfkkHUlh9U0HNQYWYcX9/JB0jzHPvHRg3XL5v9BndQsRUOSyaJhNr/bjZ84i6D
CN97aNTvyuL5l3UbFG0vdFK2e+SfvbcS3fLPws9AllPNkAt3+Ak3npCTS2v/0P47
epEJuLhi25unldvFPB6HTAToW7nHYdRZWPhP0Fp7ltRZD07sZSJMFtN55ViHwIOr
Q7e20Z8pvG5DJqP8i7JYwxisKY8rGf8LeQQbWEShx06IqLgVv0XMNJ7JM9Y1xotu
pO8BISoC1Skke0awMB0VbJzpByyHMMdvyc1QzKchmLDq8hWHVK2VhVb+vQOgMlR3
CP+fHEAaPZAi0w9S1owAjPoOmCUo3iCdGC+NrSyTqcbj+SrWMYvbwkH5WkzRpIfN
KzdS0lvlRoMf2OXySFNNjRKoW1IHswfGDZj8aFPxE3AVA6H+d2tSakBrjbjJ1loq
KGZdCuUsvu6YBT/11EWpTB5SOiS9MMCHUo/vxwBPN/MXvqJsXSEhHAaDYGLxZr3T
54hT/b9PaTbUBZruuwqaWcDh2/Nfp/MW0h8FXCJA3zDBYA7+oaoQy/Wm+PKhSPrh
Wdu2OubXfy50GifmqHAj9cd4PWOB6v3MlQ24QRu3jzxORf27iuohTc8nk8xF0rmL
Pd2e1S/9aCgGk13ESH8l4Tw7KZU/3b/LavHrPMweS18dzniT29FTd5fR3yOJVDm+
UF5fOBaeVHrfd9JBiNMfyhw5TW4kEVuxnQN+EWlEQ9AHzRZs/Eyh3GUvAr6idHPD
T7P7xHmmAzkbNvKApmlSTX3yeh6rmlx4bYPpn+shGQutyaiac3/pA1Nw/Nf/MUCi
HamR8K6E/lrOlgzy/3dNV6nKNdPJB99elXWLUBsAca90xCsadUW0ucMk41G+0jl+
KK7h9Cl1N9DcY7BzY4xhHDIqg29Xktx1Ov5bfSBQ0xV1vyTrhVEC/NLyR/88lncJ
X+uOSuuAz3MhFtX0rFnphRHgACGBJkjVJw17SmQlxFOwHaKrUI/PxSGRaQKq8T8r
pDQ3Mqd5RV9ANQM+nYJvWbzQternckGVg/Ez1PJSvyDynghS5xIg1RCldiTxzknw
yLhwG9f49x+wIBD3OG9VHJgb8sVQHuNWdMSp5YbWRTXLlFQZWMTRgxVp9lg9eXQX
M1+Uy16M1qwq/9PHzlgY3Cl6nbIDz0yQkCcct0HEYEALleOZbOsaVNPKas0O275y
m/qVsb2J/uWoEteBKZL+6pHZud6x87jYUA6B5uYpIRkip8hFPpuowtPGIpQtXkhi
9I2QLT+ILVwy6Q/7G18Pes5HUE/vI1nF9eU4fw5pWBvnnI+fbfi4K/K1iRGPkjWL
irJ8XNynZxerh2pIn1sTs1m/48DRX6biEgeuEQPaTiAIqGxnUWZF0+MUj4QuzpSt
4PFjnKB7kT3neIU+/xwlhVcViwmKWdELcIRy7RQroJK6KOSO/dkLjG7jdB6sYE60
fKY8kDnHfU36VbjXWmZKCWzso2kxvS22xJz8N0nXl47298y85uH9VuV4UAcmPPFu
FRKFi0NXy3FLFZJBMC4LjE3Y+gxDlPjYKj2u8MK5c7FEFFfSety0LdXg7+VSRKo6
GSQ1Ar9AaYBasLR/uDbl+RZi+9tlgeJ6hqQhRC6tmh5njh9e+SSZHpFY4D1kk7g1
inVeIIdl3jMmymrzfXk7s2bybeMOw7enfNljFlt4KsF8eYL/9VWRk7jX51D+auwt
2eTKapgHr9EoLIxsZXEppVt1dmbsS3uNtmdeK7luYyffChYKPG/LRdXFSv489ayf
RCuxD+EnYZcyHaYkLwKFihCVS+jgGKZeIMH0Vh7DuBZqO3aMAAEDlVY0qc/Wd5lr
0U2dHHhKNC/KG/o6t/+LLEYSjaix1Q+awplg751Co6efsp55egk1iDGDhvy69dvv
OHEtygCU//WZJtNVTQooHr8cJueHNQC6ZW1cnyUfXEe0hU+I6W0FbXM1lgI2cgSS
KwH6QJNVUKRLHeDTWy9kLR+vvnFUFiUDU1RWVrDL338DfixKkk3btB3feSzYrNNU
J0jEaLIrYUZz8UtVCJ1aMWFZnVLrgSWxrYt+o0vTGC0YK9+IsfDGVe3tTzoezQL2
M4HqQQx+t+DqqqApETlriDD/AqkrZIvYz6NgBdT4mPdWiQkm/s5cvTN0Wb4p0+dt
aDURKSYbdcgJWsNCCpHUrEAXqcapQBu9Cbi10pKzqgrMBnDkuDgPyOYokfZCiSHF
JTWxBZTzELS5+3v6CFSrAoocXBcN00Is7goLqYKnd6cXZMWfVz4BG+Jt7gHHD5GO
k2Z5IdAkebhhfrCeR1CrsuE5ZNop6KOBRtZ5sFmzt2wVFzPTsF6ugBQTV/0EmOcG
Uc8ChOObRg+OQRhHt1q3HIQy00YNh0HDR45X99CUt7kwPdsxyLl0uo2fowcDEzH8
yZ4EUQDxond5j2PLEzovKKunawisP5XaGvuLb4NLHEUy7uav5Ip/m5um/pP2GL1X
AZ1taI8dKsg7JZVZaS5fnxe8ThpnBC+B0GlT0uXTPm9jz/NHoovzqQVprujcp/UK
M2svYrl36PMACvX5BbA7GlJ1phCyULIRXLATJ+KXVsOHijE5FZlCejrOh7GaPVei
jcM9EYJTUn50QL6xg01P6BC2UZbRKAJ3tWCH5kDUD1u0QlKvlK6ZrXfi5iTV5YUX
ZE2ggKYEmyLBScB3sJQVRoVVJ4FSiRATNnyDfVahI8wX/flv8T67zqZyhHW6U7yU
gfu/37tWBeGuHsDmjutvkG2MwDb6HYbsMlDAtb9AJAcaSHPIxUwqGfZxo845ctuY
KCSgmwBejqAv4f2nDyDTR6Pc037kaPSvMBk13Xeuqh0A+vAHmm0MOptpeRrsY53P
LsLa3yheVUPo1t9LtVmd0vb7t+F8aLN6dPM6dLdmwu8LdnrKo+MVbJ0aSZhlUeyj
I1tESCzzORvFyqPcNSRB0ncs7QcIoDxXW9wecB0gP5lEn1Y+Cdz7Kq0sPgZw1LO9
++tHnEpQU22ZuUeD64XyYXP9L1NyVazbeE5k810UiIoNcuJPqHX4bpeMeTtUT9Bd
LcqPIAHSb4tyEL1nThnx3WaaMs1VHUPo2sQyrPGQ3BfPT0rKMaXDkoHMm2+r6PeL
VuNgOzfmrtUqBXm7o23Tsbcp1l0NSv2J0L2tZfy5IonRXPC8jSM4Nc19not1gYg7
gW7JP2RDpHgznapFVdOOIc4JxZC2iJV7Qd6cViBfvQ0Peo2ufYTX4at/s58aCX4u
xpq+cNPglLHiOpASI+Fr9mcZcA190JL2N/9oe2JlaF2Z/KERHk5++kk0zLapbr6M
Eha81WaPWA+nOuDjWzpP9cOknHt5EJVHxmZWgmkH39WpPOMmj4x9Ncpwwwh1ujEa
RWp+8vn16K3tvjoC9nfd8TRNlLFpoWuYEWW/rSq5eNT9TRF4pT7p4OCcm+VY/ABr
bJjVAFRrmEVUNoY3yKHtjR0WAUNG1KJiphPJCeYF3f7QsCbZiwf5mYqCcF6ggAqD
NGZA+2VoRMZxZEQAjV8PhsyRTNtyjXrzB7RvlFACd635+IaoGeRN2HXNAxkmxKKe
QgfECzuerIgMTpcvWtM++BxoJJxXsMTKtPRhrHriaTrK9d4s5bg815AyKwscH1JA
e2dELFhsakzCh06tGJYWi2rVDRqCj4ZnOBeRf081NbVrd/hnAvIBio4FYsz5UCCX
s+vpvJC3lci6ANLMWqEU7dD4vuQD6nWZnyFqnvlxjGm4Bd64FPYi5cWbyFzUdYD2
Ciya7sE4NyKDWpIgqztKVzCLNOTg7o8/LgpPsic4+G2O95kROKNoiUWUFyFCC5We
yjDipQ7RtIFl7MMqYS6PPt8mhmNC2h9IxQpczLPgYsh2mGk6c44qZjRy7GyOUtk3
Tw0eW0XMGua8kWEkiHh13SlKrpXhiyR6DfFNyEoud8eWO3mH/7oNMFd40l6wZSnN
3u/Df3ZGSMZX9MzpCbeKCvmCaSpO0rRNCZU16pZXDliWBX5SVtDPJ2FUrnowujM/
hWwdottCRh9Sk2dfLYdIxUcSK1hJRX/xTZteMVGthQHGI+jGgrIWU3cS1M6jxa0K
eJt2w3dEE/HHRet6FIGZ2m0XH0A0JepW2QPRapDn/x6zFIou1K6/nClyfdchopuP
IGplAyP6qPIn2j8rjBScfgL2YgDZs7f2ouVk4r34EoyJVRfk7xU4Y18EFvEXgToy
h9b3ksrZveHaUUAW9QcVSOZ4u1aMwiZUFK7BkkP41+TyxlKaCAAV3ax77ZvNjla/
hBunUeTy4jdLxBIRc33DTCjzJraDiTi7iRSN0mPTwP1eqXUry4IctYoHUSLFt5Yh
UBp+6WOm60buobBfyjjuNGoqeqBbVWN+xND5RQkhxl1971U9Bmvd3x8nDHpHMqfD
6iy4toLHDoioZ5Xz3cmgWPZ+5W8NOZ7/BrOuqZwuAwC/SAldTBjjIIb7xgH87ol3
RSeTEZ4Jfs97W+UhskhU4Xrb1CmK9gx0vhsoAh/8CdPuNl3g/WEc2OWUjvQc4jaa
U6rGLTKRJBta26iYMqg1hi9XTbmRyeTM4CUlcfPTHR6TOfK1r7E40aXdYxEJA4Ql
mm3VYeBl5SPx7HXhGtfOqFcGFr9N/627myJI4iEnTjWJ14mdyAwg5Ypod5ewjA1d
ospYaGgBgrpHKdhaXK+zSqicK3vrQARDyJIbdwpVuJIj3VzBTPitzEJmlSmOZ1jg
6PM/RdJTBbSCqRlKRLuTCcKoL6NXBVsZCL3pvY+Yw1GklWPn8LhybtRW2FSp8Nek
AUZ0eaiAEyyv8YiReDgw9nz5u5A1uy3shGEviMz+QDS5MzBQqkScC6rdDi6XUOE5
Q/D1EDyUUfChBLGzZsyjdrZbwACUXx34J36S4IBbi/O+rNIxbEQJPWsZPKU8p/GY
X3kwBVoWvvmtX3v4trmJLnKSv61lhGgYBuFHao8Nucn5DobmKDrDBDjVr8TyE7uH
uFN9hLsW+X5OZ7qKq/XamFVH5DwuirT9rMkWgxPEpErmmhnAiCGDL9M0Ema8+53u
TxuNoPm5RhcXNe/E4JZ2p0uhboxQncHZTRBOJIlfH90HkT5kbD1abytPSIzgOGwZ
rBkwnQOdmbaAXXcROjs+E/53kdoVGe/si7B8mPgmI0sA7M2Y05/SIp6hWVMf48PD
EPMFrnsDAb7WFYq9H2Bleevw/mEgrlAhcxDnLaOzoIeOtgeneiYdOYNpkUgbNk/t
DKhynRU+mnjUtOyP5jY3ANV2PW4bYmpztIe6Js8Zfl9jsF/gGwcgi+tCuQfRZZYd
qvQ6vGcLD2VsgYvySS6CXjG34SBbx1GEEJ4CSkTret8KdiMTkGQI00PL2wUbPMpH
tH5iCEwTNaZOj7jZWB2fCY+aZlhRPqOAlzFlyBVpiE1wxT8tT8up2A7Af/Dw/CpM
xnygAQo1lsd0k6+t5N0O4Euc1oaT4UWweChqWNM3ro4jC0lt1w10EKO8LT3f1qZR
qQLuVHCGWQ9w0x8V/vSLJRCuks+jT5rOCTe2xjJr0HA9CY13wRXIL3RFhleyBOzv
zCUVITwNjFo7XVZ7stlfflJe5ZjYBJD+AEY2IVWOVXyU2gGDKoJYeTU6z+x2UV38
POicZmH9qU3PnXXhNAW5wX6eNa2oTjKlJOtf5UQ+2902x+a19y7/pLx7UZJt5knB
yNPprqumUpOGwLCkrR82AeJ1bZqilba07YPj3BmrbYc9Zcqpt/eDUV5g2V3Y9hTT
d9iqzVdTzKXCesluJnwDHGrWARMjO8hDbK1dCiUe8kAezbyW+hZZwOpiPZ6qLDdW
sXmGj0ecnbI1omDdgPE29OFQ7x0ywlBmThuqsLY+fkX4Mos75ALEgp05j0CCYFIt
F4TByn7u8W38OKcxZnKcalpFEYl7xs1Sn83KQoThtqKkP1KQ4+sQ5aaIorB0C1DV
WT26m00LUJhfGBWQDxElxNg3eVhi/81ZuzTXpiQ6PImm2GkoU5Q1EHDG+9O5eI0A
cOcs4oFTQqlRnze03Cqjod2C0NUKfc1KKHT9hEm1UOtEwcqyo9zzh6eoUG4y+NqG
Ed61WYp+Of1aQAf2gzHH2QcIDp50FYMOwGP0ViL6dyQwg3+JDG7nGuEh3C8JOrco
b7rOTMTfZTBXamEFMBs07iAd93E/EizjrD5erjlO9YuMhOSSO0R3Dh6Ymkcx5d4p
l5r2CIcbDJpdIZpiZHdSqDqro8r2lCQjaelSL6m4vNRe5MabjsGKMrirkUep85pC
a1GnesIkxyIhmVQy1UNBOzuoTxzoUubEnAGy+JqUhaOHWzKaQXVuSND0nHWz/NdE
3Qg5DphxqWcfHUFY3vxdWUFIpzyB2JTN56LvpsnNcCHz7aEexr0XUCRslT5SPc87
FE8HscjYlyP84tOlhJkjINYONqNblO2cMw2PK8J+7IFhBPgnleUz8jHF0Kj8pcrn
fNh/mPC9bseM+I4t6xhsDtKazhs0gnfYYUw9E+03apM/tTZiQiKyigxmUQzYSbgf
KxVzsH2BbJN60wZ8mJjzzWUuO0zq12DwYwLreu+0tTf3hF5nQpoCUys/OKrsMW8W
7LovXpH5+NJ4snzGOe0mAAktTZq8GCdh9vREPdUiVCMIdjesvb1KDlkZzRvpCA7G
zJuY17jkfB2c3P4UoTYVAZWPVKkrLWxtHsO27f2HMueHdeXNVeKfUFt6kXyv7FTn
REUVPs++ymYXAyPuP5UPuMyoa42bnz3OySpoQtSljINJ4QmVUxd81VI+u+At4hpa
6mpgaEz65Azyq0l+vNK6IbdsbLlxsMH9kloyZk0fnl/IqPMfCHdoXUMLpy/fJBEC
D1wbkrOHe/XqHIbb7P31IoLz48yr9U5pypBV7XDKc9WLcjKOy2qKOal6km0Zcb2M
+ISM50tc8qSERJ05c/GC5FJT2U7712Qwl0tQHuU+tipZixtjJ5NaNLXH7XD8YClG
pe93bOXrODXzj5M2CvIB2vghFu74sEnVi+feCYJs+rUC/ff3n38lR45hev5OcE7v
f0oaS3FvMq8lOvfHAuIa60hcN2Za8xF6/P8Tnv6av8KrO9fPWMFINnW6XwmKvnqY
wCaxSE1AzFPSsh8aCwUShKsfVEUFRIKwM8/BOhIIDofL3SbNyWs51ON2BauXC1E4
TvSrUAcgr8cZYVBK/XN+41cLBmhOzjEGXEPpCkEhAZspcBCP8wcCD2Gs+hK9Uux8
41bTYUNF7dIzirHn1C7yR/el6wPnx+eOZxFpDbHWb0T3zISP6ys81inFSOHyj3J7
DZhC6tACMLyac4Fo1w64p4v66h85Fs9YsrSSSxeWJZURvEOhqE7UCLs26Ukekrym
WwPH0P7ttERqoByUFmmBAp5HrJyqJiZOB9dleOD6dGBs4b0opZiLgB4sExEEqCku
oAAjhyr6H3GExdYmhl0huQRJ/VkrjHSpcJTGa/HI/FwNiOo+3eFqpXVsb6OUoPVC
k2vZLwFmjjkqOJmfNBUHqHx/hiV+kQIkjhCPdi2wSDLnQK/n+f9vxNMM9qtOlJwV
Tceqqyh4L98nUU5VxBWo0fGvdaeP1AZ/hh3OISquePhBDTl3X7kfUUMokRxxv+sO
4IXUrqX/Y0J2DaY3tQC/vPKiSeOHUUDw3foBzVFu2R3EYE2NRjR7lm8J5nXVDZhK
GNe1ZLfkqXbqGMp5KVQLtJ302NSDkx3mutq6ZFDz7qnwwKQakW4RPqzbfN2PtwDs
dvHT3IT99aFry9OunCnHZjChwoQzz5vmLx/yLQDlKB2uB1h2HurdKuEzewoD7EbR
EtkbQbhG/ifkgS3zyPOywnHF/RQssAbFI/POn7hSvV1a7raHTrxVmy8Y2v9Yv2ht
k1FPMoqS7tnv4vLEFstOogxbHpofHNM0a3S3jn5WWb2/lOL404oSwIaYJ4A71l5T
pH8tNNRBpuTdP/ZUDsqSHrNlR2YhF2FXT0klwwTsERZfB/uXqXq7MfVJ7nZpA39x
YWN3XpglaOftN4ZUbcr/e5AyIDMha4w4B059AqkJdJyOWo1ga1KMPIo2Uf9UH/Vu
cXvk6LfOHvJSySr/FrFLOVlXaTPdVtravY/02+mUr7U5hxhT/UJMy+K1scxtwafK
4Bqll8fuNEvy/a2sJw3rgv/fIjR+oHtyUufXPMXRA1UCMAodNA7sWqaCvbw+m76u
WyOipCErXkJDKXbsJJb06M4d3WTiewl2sdzOuA8pX1RW7gHopvv1Ixm6fy81pnq8
VKg5TT5ZP5RCO9A3dtRy6T09Q/u5kFGFeiJ6GrLYTyHE5M4lSodC3LyAK9qaBy+I
DkugkKYOkFZ/iQdPoE6mMmV/A/HO4Jfz/30MTd6MtkGzSTuwuw/mX6rvg/qU7PBs
7aJpveRPWE6WIAcJTq7hFoPslIT8UVbY7EzdFcnT5iicNmUK0yzHO6S1GR2Nagco
Ew4jswqO50KAVpxFVLFLGTlTDMEhyotcoz8DPtmsW2nOU7dvqBIQcaw03j+Yphmp
w9/2g1TJtbMZzd3koNkqEDRlF06dpsA5g6D19mInaQ05pOzmPzcVpLGCzYZj33JG
RBOV058U6VMBoGPkJmtZs7gmKSiA801CvaTUZC0LfRgLuZmByswrD/2vMtotbl/y
5J2XXXBaT/Xplu/AqRIQ0Qx8UkwK3q2jUf04sTMj7U/EBR/T33F9NDgeJXRUfm0N
9+7U9YU72EK2CGWNnseygGGno0yzuoi3VWEyAOtYoXlCqWMZLkR8r3/9waDVPyMC
lPXaj+4I1Tew1TEhRFar308eefzLf9KW6KMJyztPFvXhvii3WlrolEPNV2uNRXjS
/cvIO4tg93Y70bHa/CN1ExQah7ugYtPS7i0KwlfD4YAsr/cp3ZAjqznu+ut8Xn/K
4ldz5ZWCNt2O+vRQ++PhTfGCFdWBQFSM4hRk834BBl8Ta7xeem46V5Qgp7Pv+O93
dmByj1SZnc2sgu0HcpkuCRlQIt0HWjXYzpH3AHXAVntzAi8ktcjZOa7nGlfPDamy
NWnaGIkfZwFgfm59cqoqsunylwtTPU/6xzu44UhGkT38em84t8tAWGyHugHbkQaE
Nc1s1KUdCJVej7DT2OLEGylRbcZgAZohUFby/4TCg061W6GyrccJHbkVuD0LiakR
hQ8pIuR+T/k3Pvo3iIZm1gt96gr8PDMeL6+7JcWXqX9QXi6FVuQU41c27dWxt3WF
YrVBTzZ3d3zFHS1QM8c2EVW4uzc+EmjIj/S0Ep3nEySjLuSH59+X4aEWrKDAMIA/
cilxNDuA+GlMFFKcyRncSqev8sbKt7d8AVvSN25GCHHJ8yUVBJUZiUIzk5TvO87y
KS3XYb4zHztidt3+swUWFmsiiN5MqWGoHTvViNq588kZomFNHLuDQRERtD8DW/Ns
ksVLMSMk6AUui2qonlKU88EMzETE4niYHxQrRCnS5bPUZjfqElpjl45/DCycXOLU
KgtRDr0S5xpXn8CRnzoEqRLs0RCfEfOzZL/4I8iFGf8+J652WI1XaQwBS0LgEl0g
Afa2Z84mY1A0ohY9cVgsUiKAHl68LE6gKLy9PoPfeYDwwGl0J0nzJFF+VYO/umxH
cMrFlVv9oy8wnWG4g4PeICY0b47X3Hg74NgDjTJGkRSkzWS8b+dbHr0g4YtatGPs
sxyYGvdegVTLKVY3mQuyNFK8u9v+tOAbgwZy9xyLZAiB8WW60hSnMkyd6/BKPilC
JiO/lCtIzR8y3TO7oV/FmfPzzi0YeagopwOz5GKByezkcOl2ywkcrQqMvlz4eUs3
4DdehPsgtQO4oU5ljp3aHi9QlczoHUuIenMozBYJYACiYOh0kNk0n++jQ7tjFRoc
RFYfN4l+ZlDk87VPbpAHZZXG08u7kA4tD06L39i2TN52DHi/OYL2c1tJO4+phQ0V
G2L0OsAWGT0h1lCosX0Gz62JDwMP3oCLs7ucKn5LOIDzk3KQC2lk9M3crrw45uz4
XyWaEs/cpWeMaPdD6nxUquTWPTT3H+3vh/nJAvTbJajD3WruhWsarAyb5vBxjGcO
RTCUHmJKCCF/Qza/1A2TZoPwxM+3PVMyNG9k9uRlxRYK12AKW+8WIedvb733b3g9
OH7yZtpqEHb/5iXvxET7gbEgvIsCi2+g/3woQhFuTDHqUBbBr69ALHajnSGo7mWJ
iXkC5J4XXeXWiyUxMTWmUXq5NlzGK2pisBaVE6IgyR9Zai4U+qetbavZo+UdDdi0
KfqTNsPrBIdpPwzF4acbxTmhwUR+xKNYIepza1iRGCy5QEgBwwi0SwzohW8wVeL6
T2z+tgIBavZpMn72Xcyt7HHB3r6sb5DggIbobyGh3p3qpvdaAbpWl8N2fjSUHm4V
gEyAQ+S9O6imFcNT7ZfaAIWe+F8z1m2cp5mnpM8Cqy4G38/4mo4XLRFYCZ9EiN9a
a5f9yDZD6NjwFNRP2fvy2CqMmwyjTwq++GHGBJ5hYD+OdRUHKGadAJ//Rv5S/8gP
sZHIcqq6hbKDKhkDPt0yUSktcXKNna6IrmWWx5uAs2XmqDefHvbdVx/m/TZO+55o
Dz/TJ01H0TWx3R5SdFKKA1E7Sg3kRvYnNYYszn+Daf27B74V+OydDhg6H+CtD/Ss
RGe0CxVWlhf2Wu8KWfIFhubWT7vkwSKQA4bI2YEWZ2oamesIB/mTCZVi7yiS1onX
uSqgo4Ya5Yuz42cYODlu76d8zegKjrjUX33B/3oWY4X+cK7fG9+H616z9E3RpYLf
tooeFH+h7CjJoYZjiAZGUDMyiKZd4kjRyd0dUoDTiT/iDRJdPHIWV/8HeDqNXNWg
WEiIsjWoqsvqbwqWFv7R+QahcVlaRJ6InhrtgW1qJr5RQcIkvaCdQZRK0uAqGa8g
nN4f2pEBW/wZqjFVa568sEFj2wgaGJyq/hrqnQsXYffP1QJp9IJyChgwZSRubt6Y
Kri2Kh8tStZqvklr+PrQPs4eiIXFyg794KhlEVxNBxAuUJ5sMzPwnaIXu42Pr0RT
sYbs2iijWP9CHMU3+cOxpzQv96uINyqADPniWox6ohaT4zrkgXBgP4p4h5rwx9+N
IZj+dQxfBv3eUTlFwEENgZokfsydtLGylfYfSOpxLK3QW8mDkuDSdjriNk04NZzE
y7sEn/p/jNAYV7aUZL2Ijcjzvj5y1tmCKyhpGL/6QUfrdgsQip5y/3Od0ceOPh3y
z+Qm6lwrF5gsidbhbgOUsl53DCxChZuBbvl3zKCooBHCba/pljqkJEDt+LplVPgo
GVkJ8qsS2ZMc+Y1Ub09i9wQepYLwCSG0nBZKGMKuaP2G0xu5x4cmraOqJbQOQFX5
n0VGP2whNpYHkX85ZfXn0kSIVgfiak4KNrFkbTm0M4nTHlKaLluISou/EZEC0Yr6
jnp+8uoBaqPXPdn6Fd5a6gmij3OKy9rz40Mq1WXGhtwyqoknfB33Y0pckYzNcVzf
t1y9/UH/bLUQD4akchWorc7G8MwZIJ8lEQcRaBYwYvQRlWbtorEayrH2kr1raLib
xfsEwDDuowA9gIwl3ZuLzndlJyD5B0NM6OqDX9SoFDt7EYTOzZ0/rYNGtfNcVf+h
W+9YqFYM7R5O8ihj1GiRAZwvQq1x9JMz4OBihA7q8V8+7dxsmKwcqj1hsGWiBiJM
CxLmu9RxkwEJ0sfMNHur9cLjkRq+qpMYiEu8oYExkDcencHO979O3y4KaSPcK6cF
oRGFpQZ/5r7rFZm/1CO6CnXDkEPUn+BUyCUeaZ7h+VSFZA9zAIoYoLeVdphIq1uQ
I7atliUqFOcSBIbgk1D5o1DucROaHot1KPsY7xOoUevk83IP3LdrMdkKqiwnTV/D
N9VEigIu40NmXlbweQSyNMwcvXusM2qjPWgbo9DgzjGiWa3YlXym+JA5Sq1IXT0S
3qSHrJYpuVRBSWd7Nre+ea24nhh8/y/t2zfr+OeBqGXKHqzvdcl7UDUDf1TGCxoY
+buhy6I+nGXqsmHuSfubYJudI2AdLkHhBgui5nk/dQQpqIQfBio5jid5iWvEshIg
tec66mKBmfIF0zZmBSLe+lq89rSIoVhxg5VnuKZwbmTc9f2WKvz6YMPYhDAwdgW0
eMr7ao5mFHtpnL4iI1l6JPJV4hUEUcm0BIfBd3+sTTAVLtXAeb/gegI2GtOKrB4q
aZYSAdZJR5borGRodrpdZjjNEUd0MPlPGReFTNd0b2YtZO4FYbRH5q1LNdwzR3qk
T3ytU1dzWWnEZIY0vfX/7zdYlPpabJ+fgcVDnmxJkVs3Uf7/IYbs5YYBDUZP/cAa
lUHRndEGkkOYbY4WkbLvdR8csNF2TRAW/HTfvQ2FokoxmemVIccImSbz3CTpszDk
qtDYQviPoNxagr+7VTm6x75EUOMkZTZwM9XApwm/opORqwbB2gJunTI/QtYLH0nR
kY4V++/Oj4qUISzkAqP6RNU1n/sWKF7kOQfHbqkKWmuKL6nB2v77I7X2toXVY61y
35vWk2WfIJrIBT6bh69epm6694pDzzb4f3I98Ylyajb1tjIHlLecokCumwzieoOO
4527GAc0+zftxLkONqTfZBa5DuTupCcKPX9b3LQOHuYjnbYg2gL1zZxVC9GemxIg
CU6SEJcX9G/zA2cWthla1gLsapWzabKtO9yrTofU0zBKFCMeRbY0iWmuMUQ3I7PY
wHOLu8wTWNuM/iNhFhmQ8XUfAZWs6AVD6jI9c8r+SVoD9AGs03bNxITJgL1XtSxV
3XpAyhVsjE2ftTM2jCvNJmn0iyz9u4/dHwC/IuAPCXACcMJYAowU9Tx+hdR5QfGx
r3+yA2yqNs0GYbfqDdIiERoDzuVAW7P/BkWfO/QOpBbSxaA+Ds8ijd4XQtSv/W2k
Lt/dT7I4Bfzmgxcf6UYgeeNcGI5IqycpzM1LV4q59LWI3hV6/3Blf6J5JnjbKd34
tu6VpPLPjgKjxX/UaQdNz5w37I0EgElpohZcoIfVr2LUKOcK0VJtoGbW+UMqyXwA
L9HN31j7gwwzPq4b0jYJuKRwHPCsR5LuxONUYiEE6S5vIbDMJSctZeBnvpE68JSa
qZ6cFOa7TdCpj2VSaqN74sRgsSxFsd81VgHBP4CJt4wmXbtUL/+oJsqguvl5OzCX
pCGPbOZfK1AYYw8vHPV3aU5gR66O4Pamu3GFQDM7IiO2VgY3uIznOqb9YjJMJArN
Ggbcj1JLfhLUJRG5PWmNIONh2tV2oL+kccoSnb4tNx3g9heBtMeTPJwY22MEQJhd
4XASqXtfOo+VbRlYBd0/qBdhSe1HcYt/vghZgrbGXH/LwGzW6UST4thFkmsUJI0s
ba6WTwxa/EcErAhTQ0y+aDz+5C84wvfO/vrWSsgVnQsg7w747Bha3OwX4KEJsjdf
Lj+lf1zqQ44ANc5mSE9WzEEP9m2sfbxcEFhG0vpSprjmSaOszN64rPOPTHus7i/G
UTmlJN3HF4QeVlw6fnENs4diYArmRKi4MEG0g5f4K1IoHmZ6B1UsOrcPoX0S67q4
Y95Uxuv/9Ly6Un+mgiDUEIkJ8rusWi1bhnXJt0PYAaPpoB3lKIdUVuumyflgzoUP
6X8usgO8Vh3rTZkg+5zEBm1ZQLWM35CyW/g6w/xWeClBf84Cplf45OeDLDnGgHbW
vblBZX0nCsZms3COhvkQAjbPn/am5/YYBFZ7D6pxC+16HurzzRIrylNMxyA5x2jy
uKoD4qSmC3Y5CGciLYxlGkKpVBfVt+c7LcdG7k+ofyDWcOO7iMLSG8IAZWRSh1UM
RFmfqF1rnnMq+mtEaGlMg8cgTWD9fVo7dSzHdbwyNeFZwvX1Nm6jUFhQrMME4Jk5
oW7JKYxDgJYXMRpFDoGwM0leEDD9AIdXPgsQ2+cblVYX+Plx7hxp5NPHBxiTBKHH
pki92NabXwYT3xB7+8pZbWQJjFm3Iky2LB9UB3ctpnxz328ZSHcSv3t/hONUOmkt
X8581xaKDgXT4K1wbQ5YOoLhd7xgWXMcsOetWLRsQi/jGUo0muZo7DJiFnMfABwz
Rrr9u4L2u5P0VRWfPlxJgwa1Kw88VdR0t0/Q9SulXotoufPzZu3vAqw/sVuOhXNq
yQNXJCvs8iINgoM/s4PSCX8mVN81n7rZW2vbf8fBuq+jsPrC5ImkOmxc5CIspu2b
DdC7Xwrb9zPDZkpDac45RPFb4PM5uwCIorhyvjHGGjEFIT9J+yF9MKpYDgYvcqcH
wAmPsnZbzgntmz77M/9VE/m7WcDwnGrtZlm/D1sdn6FgFWnX2Z+hZ3p5im3DVY0J
6fCG1Imb23KK5Ubkaqn5oo2sHbET+FCJrHkUAjI73kAPCTCgLlgFnjMtJUSzYcSe
8iIbcfPd4GihE85wbBwrCu2dwt3XTyUXQ+bObOLhmgViyqooHlKE/YsgOo5shLq1
f37BlS31LY+r0ZXIh1Dorg3Ub1MP6muy6bqbgJgpRjymwDmjsQpjWvsXFEd5Ip8l
QCjOF7WtLH/6JgfT6EiBOb0PE2V0mU5hIbTRWXuGhXk/XQhF8db4w19eDgdLnoRg
JhfLQNV4WWGgLV+2vILCWj+kHX8zg4WH4zRWRoURUagXQXaChrrzYmGPwhnB7WjQ
ylFxS+k62yOXUxaovKVGkGb1eF8tF/5EtrYGO2+/pBbjA2FRNuzT7TURu1QNNGB/
iF1Tx8CyBfqV6d9bcocx4bYbA4VSaUzEmJF5wpz0f9ko03pDjHLMh4k8KW5OBnUZ
I6kSZPNzgWw1g94x2CIfqVtffnRNM3kasJ0C6YvvMKXSkmxlXRYp37DJ2UuGnnsD
Cmg26K8wJ8L9Ji8m5jEQrXuexZ329qXwMCaYPiLZuR8Qe9+REi8pXzPlUxzX2Zbf
u1A6kQ5fHXW/u7eLy30Zb81087oasIa3zxrI0RDmy+uS9uCavaCrvDHKN+HsO8wh
08k5+AYI3K+HVxWK8DJgEkAwmxdwosxh78RAwq/OVhK+qKsKevK1yQll5iwH1mzy
uq3N8E/jaGBd80xmOtP7aRWBMMHN6QXUCIIvWHFe6AsoHu9NbJx+TRriF/q1z9ym
8l7S2N9nf29B13U7z9UsF9N2Et8GX4i3zbdttnT+/ir2r6GKI3S35T8UQciLclUN
o4E/WtFswpzD8ASriB43jMegwE2PUGdap9ppwp7/t0q9kHmJI6Pz/msld51B8eKf
yO2aKjpTWF6BeFtQgIOVQu7dRP2awIJ/PEdW0aZlDgfYMlpO/v+j01N1K6A3gc1I
NSgCeZ9Lx+jsCZpOb8Zm8gmURG4p1B51C3KVpyOhkwNkub+zopxrsVbONnXtAKAd
fQG7JMGWsJY8hPQC+LGu7IxqKXZpaDq8QJQegPQLDRYEJsN1JxkRqT8ZQHfhJFcR
u4LysWjjVSTKei/MePV6ZdK0JlNpRjZ4UiiPEmusz1q3tbAbW5u6ip7jQo2zYbxq
16gICD8o5CrRGmFaF4UNTiQR69rGBmjgFsIJy3eflOaIixv/kjOJwa3HA/Lvdkj1
CkLuPnALG+1QQ2lk4YzQ+kriS+vKCbLW2fGFvlxLy0YQ2xo8sBD3EcurNbZpaoVE
0JZbxN3EN4p1CEuV1nhCUwP2JRTsoGsOLS8Y27uttvyW7+xnF+rYuKCD8ytj5zQ7
EP9x5s0OyPzVV16XRtqHO6dRym5iKNVTuCQY3PUl2A7opRxloF8FvQwRbqss0PJA
LPbVSKbwsOyCRWgr3F6x12FcNIS9UZbUrWBMqrqCCDR7qKO2n4WwPXqfrxmhZNUn
kUNe3RZ+Ne21FF/1ZejcGIEZdGzdDFL1tcWv7WPFwrNmdMUaCr1IMx+HO8rEp9dq
nVCqNLtmddcpaIVyghWoZZXqomm5PoefKhnsobmrj4o5+MGek+F/QsaYbaUK6aQw
7HdXbwZBawEKHG1I+XtJzjjBFEgJA/hONuD4jkkcFBDap8ROqMnUgjL6w5SUsIwT
iR/UnLZfphe0u6lLl6AGn/IHZC8f6eG61YAMz2+kYDsb+5GZKFUYDY+Osr+cxSrO
WtignFMjz34jf802jw4f4w6uZKDLEEIpKKzwIgSrd/l+VU4yha6NqxyqXQqBMOHu
sqhES5KuNocFC3b/B0a8vERYUzQL+KOtod0+qDfenyD+GQv3z+9w2FMeIhF/HKql
pJQUItQ52Kd7FaxiTi0zLehuMSzEJMSDUTYDl7Ou1Ks/28e1Qw4Qg4JahpqPrb+w
Bpn+i5vervVmjb+RaiI7XYOQNq+OSgD59EFYUi2pEUYDXI1DBTx8OPIrWD53y4Oe
7QycXX51ZKabwOnzS2fongrW6263ndCrg2eOrxwQGwSQW6In1DOM2OtHsTdJKjW2
e7RB5UeUSdKvhNpHVqMvWEMfAEWZYqSqT0gwyY/0Z0Ua8zqFh4rWV4lPXZNSn+th
mRgdFHR9FsCHZj7neOkeOFwxine1lu/zVPT7lgYFiFTAbHdxtRSgLoRpY7ZECvFj
T1cs1RvYj/CrGU5tnV64HvXW0f2r35NbZkrejyrlRFXKKxrhTu/7T4zkCzwfDdnZ
h6cW3ORs2ENvR+3jVawn/6vg4dn96cD8jzxYzhw1HKKLxavRrPg3ScfDReALxixM
IJ64TMiee+OhZj02eaZpDHTjcgZVcWDo7+wQdDwtPVIqrFjBd0otmPgpVYmxi7rA
b8YFFW3TaMavuEzLEC6QCcy0my6xK1J0htKHbwUrTUNKiJ5rZ1/EwwFW4+eLFqg0
oG3FUCw8gurNi98hug7wddjPbLP+50ltRHJYJnLKwu2d8JWq/vWrtB630khYAy3h
SdsA66sZxQVqiRGeykKw+pfYlsyz+U8zagJwCr3ofvs8huDgnnH2Gf2k6v2SuO3S
GhIiQEo5pymqtCov0PNrDhnOfQSbNhQxyEyDv/bwChgV8qh3mydp24AY4FkNwcFO
1iw1XpvWKsw5UuEhJrxSsiGAsMXmPWXrixmi1XFib1lBiLAQbx5Zrx6UutH1gx3f
4MS8JyabLGUKu2R++fHUffAzflDZo4G4bKz+6SyDOoslceutWspviF9+x5GGz2Hi
/j4tCeye6vAjU+EuGF1hAo3FyZB/4QNX5JJTt80jWJGOkc1mBPdRmpTFXATmzhgh
57PkUxLmLF7oxjyQbLeXSJpcGeIqXRSqG2bR4q8GPPzcD0Stq8ZiMavb/kxr1ij+
Ho1hg5uLs4bFf2OGUw8C7xCPX6NuxHXY4JIsOYloiO3qXY4apEZ2M3iMtPrSwAhE
leGKVSS2hv7MLRxe8LnYnf8W59l1PQ/CQuM1z6c51bfgCx/kfRURKWdCnyWDOJh0
p9jswblsG1PT4bz56G737kNzKjIwmZs5XTJXZgtDU/8Xj5OPNgYpZyUyEcyOA7TD
UtDz2Rx2B1Z6OhzwpM+rop4JdSAZeN24HmDyCXW/I2eL7uibn5tiHBHYY/6CMCTJ
qx6nZpwCMTCQR+pVQ/4+t8nTarpjLZQTr/W+tMEM6obP3mBEakZlhTdRz1Yl8cnl
tKdqTeZGracLe+wQ2rG8l1xHTmwJ9hAxCIjRWB/qsEorQL1Ugw51/+mGHaIag+GB
Ob56PCMw1feOrbuDupQH+4B2Vb9BpH7+g2XOnbaIbQIn9B2RJoLEq3HRnkCDhEc4
Am1tQtq0cKq6T842XPXUraN2+DSePawrW9ss2accQX6SeaMk3YpIwubrox6vKRxJ
lQbTYmt71JEOU+BxRD7JLXRC5BIFHz6CApYuJkqPjw5qXeWz0hHW8oXD8vq3j/D3
u6rXmsaC3QFM0RgBMZ79m8AhISNw9CTPsz5smG0Tq+Kf1nBLPRD++bAqUFV1Vgw/
nMwSN1HTcIfljO4SZQYtTeYfy+Nb8JUnrFMp+cwKr1X0GcYytF2j04LESK/lLXgl
ZFfW5NXeVvrEdSSNkBWhGVRxYd8r1p58FHNOdOu69WHNhKlZfUHM9gT4DMPR1fEB
qgrNIGzMpZjIXO+6PbutXfMGGFbYNbjJV4E539bnf1a+4Gp2ioZg5z1R9M3XiQGi
SqzYsUuNlIREzPDr3YjKy2DJ3U+unvEnwnvEfTtMwoUeDgn+R4qJ3DTWJJsxdBJv
AVDHByt+y68G6vl3HFsuXnSL+tetFKt6eJUctq8U5zUw8zThjOsdavrxR1Wd3iG2
1QI0MDsJCMlAZmCcQEdC1RZ0tWRcYjKWOJD6/Y+4AGfte3Pc5C8EDSpZzbqFWxm1
ngI9JVoMdV0RjcYWdI5OQPJSXsGQ4uz77TWAEWKZv3ViOCQRceYxHSN9uIAH1LGv
s33L26mvYp6xc0hMauohahsMrSIO/Ii3225762V0pYgubrn5/qJ/N1tIZ67GsUO2
4YvN5t9kHVeRACkhCpcC4Mv2hMqelCnOyOZTHJ5Mvmvx1Ynnye0JsAWKpBCT7+jq
fcCrV3xoJ018d23Hf7CKQvk6ZGoVy+4WvOt8uJm2Mcdv7QKtKeCotGUuRCsSzWnm
Gc3nndtjs9MfQ5EAXdarvF8ekLdbTxxRKgfG2/WF11VTBWhOhLrF8XuixS6qXWoq
CmHb42lo1gZ3rTEFJIRa1mT29/DXGUrLWuSC2kSUV0DvMoteFlYxgJS+itN9kAyB
Kt04t76qCa6Icxg5h4/6V8RgIOTNGr4H7Tibom+HB78fIX25DmGQuXKiWZfKuSJZ
hDOrcHGlyYEThWGhhnOK+PLu14dkDmlNO5PTu8DvrfY8RQVrENGqxYKyoNhw+frF
S4v6GsRtX8k+FFup4f3cHP3OxVCWTDgT4ZF8niwMjrAz7lhek4hbtR1otcdTak5N
6BSMtNvwTJGkp03Y0Z5WJfw3KGb6cedzak+Y0mcjrrWWo3RZkcriaIm+t1jgzRIO
+QoHjaW/+5+3ipbsFfJwTiSrEKmZci8aMoxIFNW+JHSDWtBtPoUvvAIYeAg3E0XM
Y9/fEJ5oRK0psYqxxOjt5fE3IBbWIDmoRGLjSCVoMsHm8LFOgEcGscTjN4yG6z9k
0HYdNqpbWl76tmL6GHUS7f0QY+sxbO5hdE1nHsNXRC1BZP0GMIWbunXMHymkgBmV
nVnU2ZWCpaTcbiM8grfsjE6am8SL21xRZVuXHYVdgtiJrVhZi2p3jJUzqC7+S9zA
XgAd5IYb29NznQnsN5azg8mta3tjCsiVn5SJhf74nvEuxhUfe8oBD326ymqfuTH7
bfq48XkMGc0WpT9tRJEV16BRzl/f2MogqVDq3KSitg9jFp1rPic7g7GadRyoQTtJ
m5UUPgIWbgxfuhSBzqs5l28kflLJpSvngweFyuanG5UBS7yMpc2QjAIWvK0iUJDg
xwDAVKTq8kfj9YuYrxdty+o7eNZLY4f7ODVy/n21sorS3StqZY16qiepuSV87ofl
NwYvVLEtRA349AF82+EYGlihDvoFTJvO7j7hQILsiYl0uHDpqb9XcIDWekANf2+w
EdjOlNSBHqqMargrqK23jAhgmahkbD6WHqWmHFHtlDyW40mS2goh1ManuZr4rcnX
2nhydVL54ItUaFHLLg/XMiwwg90Nvk89n/Dna2Am0ZBq/f15+CjkTdQ7RFSlN0/9
OMHcY7PmmcOAE+1wQnFqFb12AF3cJi/fC+qrL95wLWo8Cv9bSYMRzzFMtTdm3dyO
SNoFFmErnxBmPLU6fmwaN1cUNfpwvoF25I/BtahkojpNL842S6VpFJ/Zp1j6iLvC
0S2h4ratmQ2SYVlhAkpBDqJvBybGeYj++KhwvjO4IRCxcF7SBwgcdaqd9I5UoYlz
cHqk8f9kDSTfj2HBIwXrBND5bkpwlU7wWOTZZSrhMZi49glmx8eVS739APgKnnGp
EW4Va3ZI6eXfRNvoEVBz6z2GMFQO3/znYCKGbI5nTC1eiT6R6KQ4jN3Nzc8wYXw8
l70H6szdiL2CUSYshb3rOFUp0TqvmOFa0zgRTNK/4rBc3qvXz4yoCTvhxY4XhXqV
ke6HnWceMZE/VIM/v/vnO9S2OOpfBgSTq5TOOrr7n9iiGcvG/52dVeJwuFfFh3Wx
HTcDWOcHvKkIbEgWeAx3btzEQ2xmSOTuFJz4fjXBS7QOlfeGKhePP7STZlnodl9Y
kapIS11j8dDMJ7SY9XEafKnurEPd2UELN1J+V1joBinI/A5bzASa0QeDhafApRdE
817Wex8VoxXgvhZifBj5RKm2Q1JguiZPD8DCeME9TuAMlAZDszOmB13Ah6/pck6y
kFlnhwxDiY9hx9MRqLqgH14YNqxV5DaL+L/bR/JQ8F4eKzmNrQqU3AMqTWUQ64CW
5PFN6q32qwf7jTGE/0tfDZgXrEe0I1b6yiGD+a3Fon8JhW1pHAzKaOyOq8ABYG/Q
pqVfVcY4KUlsUen42vqe6uuAN97tkBNCdLG7dYSuAbWaDcH3jxaaiLGbJCGBTBXW
bHrJ+g0XeTMnmwqGw5ijJY2roJYQSrkOz61sTm2uAazVFxV3bIrTims8V/QVrytt
x7kPNr8swc12KOmM7HPH++8beZT27SDO3htQVdx5Poi1BDaIydxJYSAENS07swfR
UgFUU+fmKZh/0veo4TG6ZtiJTAQk5Nanb7j9q89BhzVaUaZGhs7bQhdyMB6p50kQ
pasgWcgbndWE2xjFfSRtVnan+Flwg1hRH9rN2L9CR0/A2ucjVmOWjoc1IUj3oIqA
xChNHs+YHC4r0rHxsFLpKHB5AWJ01MVOqBjhz7DchtsJ9JjlmLoqy/N9RHG8OtwD
zgr6eauCMGXRetn2w/t7c/dowfpUle3uF9twImyZzBC5RD16nFZ4KHAXGa9bNkYE
sC/nkxsHoamHbES10qwjy1YK3PjBuA+bxqt0O87u3MCTK2Vk9/zKG/LWNdtLMPLq
OBr5ruKFjNRfLr4NyZjG9y+NC3l2Z9JlIsdq7mEO6Lj4F3Qwj/tQTd6c3xPvefZH
j4/aiW9T6s8xZTzrnSYhwegk7Ozj5xIzWvQZUjteEKCUCttPFIlOiBWLbG2TxKlb
5fN349VRWRwfOL8MKLYrxx6APtnaAKXFCH6gB0CgutfPl2udMtC/FCLbp2AWmFfO
WCjPT0ncSmCuNcpmNe0h0EhSC1G2LOB/MwL58DSUzzjfkgY6e6p87ewn1MaaM+pQ
oguwKY598yS+U2fZPIPl2w8HjuCkN1gIQ4qgrejMcxEIRkrxE/MqH4qIqAXc+J4p
VAx5vwjSFo+nmctnvKKVNfPiGcoLoOt1WRuAq/IhDCWv5PvmwEVjeNiRAHAof7px
l1pmKc9RWa8kPqXUGAqcZTaxaZo+hNwjudmbY7P/+PxigD++M30FOBaj17yIqOkL
iaMs/Gl8fxOUVy5phGzUTQ+1MgLdGnEV6gjvKrBDf3T2UHG6l/FIy3Gh5QlPPrVh
UFTYM3+17z4CZIuQKkfkNzM7b448k4U6pQw9qqKpnoJ7KTgVJCGkg9Q4m3+71Gwj
TQhHNKYFsQJA+s/Rrl1Rj95hKNcEoZyzuVWVzS/gpTP3LxOkexjPN8NhMzJOG3ib
r1lQnQpri4BjfTF5Hs4l1o0P+fAopnZMQALly+WeQKMq9HhpVmkni8aPK4agY0q5
Pti0O0ug3cSFaCfqFjBFZF+mrMBElcRM1TCOYR/sSqIouFgiVHrprB7Y05rF8gst
q0DlDrVu4GrvPNtUjo6bB5inTnRbk6ip014Lim2O2t8WwocGSVeLV3tZtDdioVOS
k/Pb/PKbc0O55pjDOTzk+xgPxQilSvD2Z576TnYvRGEfOZpej49gYazAMJ38F9Iy
5LzqbnHvBUvcV3TcI9zw91KsW5g1Z/7MrLKdVuiI1UHv8KCAcbEdMGO21yNpG3HP
De7DJSu6hmS9SpE4Ts+I51lxZNnSnNS7cj/dz2+m/pQ5CxuC9kS5GQK+oeCp99PZ
9OwjETbAILn0dqH3E0Cdg04rlrk40RfJbNRNoC7/W50JP0IjdqSAVrbSA5ZvgNG6
KybjeNRMFrmCTFU5xJjRHYZ4xxYqJQFw2KhJsPbyHnINBkolpQzP1GkZVRq4nAUp
KntsdxMM8/T0TLpytShgkU2gPgebkDTYh7vljJWs3jpieC7Y4hzZlx9QESeefxk1
9yWl/5TM94209Z02r9CVicqXr2fkiq6/uz+3GJYmPybaZ1l9+Pyt/A57uDbLsj+Z
Me/Bw1buj4kTBaddLoQ2+HV/7EQpxVtp2TMdxytw0NewcC9ZD3n/kN//CCnTCADY
ertVIvPaaDwpSf8scxHjBgYQKDk+90cFUg2OzY+bLGDEPaXAcw08Qzwfbzr8LHQm
BSENvCMhsBzAFWPK6QvrxVn/gMlog8jzd+s7RpQ2DY50pAioHvbMVVlPFWqzec2R
9Xz+f3Ah/n6WYOY1U36EegWazc6GG1foAnm5RzS4ckfoWfO/6aX5qBlgLcugQiMV
u/BFezBXgbI8PB6YUJEkXwGJlYnIKp9nO0FPeIZg9nlQib3Q1V3L5DW6PH1DsTiK
bbMbHl1i2Ok/5c+dhSHZoE1sbcwErDOGx9peWDN9dyLNKt+YZUfIIJm65NgB98w2
jS2/FPxB3FYTePcYDHXETtjGcD8gpblSSKqT7C4WWECf1rQzLtRrd3uCMYNby+7U
xmWJRFaaLM0g3aeVQ39qVOyhSsDYJ4pTL2h3fpLKvrA0z+OHJbZ1GM6EquJ60uck
UuChxxEklQFoOEzVPDV5kQ6rUU+nv1OSfuy5ApihUtIJ4r4q4JARkpuNPVu63NDD
nPewrcxNSeV83zT5gt5NlF/QiPPWOq+ToZ7kp+acrAt9dpi21yH5uUCLV3tiGgnr
CTxLR9CAlyPXafoVZ+b7JK1NXVe+cHQcXp42/B0rAXXwo12FMb1dTTuC7cnRAttK
XTUWwoaFjVLbJhaXcMwZ63LY0gTRq08NmIij+juRg+kalVguRMQEJQvpm/KQflGj
6I2Ddq0VeehjzOGVPZJIyzrFgL3SfrqAuZAPjFKGbt39wzFtFqtf9nDNSTcQY9LA
7tmdYSsHi7FeECPud9WT89e5fEaZWcV9aHq0cLP8DMYRkr4utLP1aRSO3O0JNaMb
274v/I8XvQsgCKJCB//845xekJJY264o4QBa58WyvGTkNh7tSVYN4enoa8AqvKYl
PWfmULuwc4zcfqp6y26j6p7529r61VK21K4zmKCGemfxRjR0FA9GzDZjEjHMrrZW
XL0ZauXeIbVar1G/ECBGf7NSGLkzpoThUS8h/mqOhtVi6TTOhaYJuKNG5CubPUTD
QbjD2K8mELOJZcmsuPxzp2dyn0vNaFNzf/3Jr3SvnSzfLqBP+a1/Pca4qjcyryU3
I+PLPtYTtIvH/b47lKcXBB4CALSJUaZ7xwXKeiLOnRITnajrumY26Rst8AlcRdcd
dT0dD4ZMoMKAM7PzXLDaxR1NCbTc6iDXlGWBuYs++kYdUKOkbREjxhtuok4mb5fh
JmvPVsLF4Qa1pjfgm8vGBfksL2WHzyzT5vMyUWCaxW0GDbvLb3Lv7ucJvHYzFeE7
9UGxyWCfDTUFIT8rTzijLM0XkaSKwBF9DsyeHRCivPFsoPGYj5DDspbWk1MqIzgR
OJ9ZFdgxKEzPgnxxKCmSjysWOrrUrzI1Vhir+dcsymD7pkWx8om1SdMl9YeXWrP7
Y0Yfntnyi7bWSIx42rHB5UtkAEV6Kbf/UWwypqfIQqbhYKPXnLRjYBoOEz8Qp6im
twO0AxsDRoS0o5numHh+gGSGmBw9zG3Yvt8130qWyu53rR/opwcUqoclHC30asrA
PxRmAknO2p6ZQ+k8eu6CdOZ9vQYryWkXHDXYd5iM0/sDWyvOSI36oh2hELh46sq7
jpR9vbSvKjNow2FQxfqEYPhIHgGnw79QVL30RG2t4PJQl8MxHki/XrPsDrWsGW/4
gX1vkh3Q1Y6X8PpyVQZnpzxPwrfWDwHGVxIbnvq+5udTV73tyaRfdbO0rptTeLeN
fhkYKPjqRRqc49WwohJ9FXdg+aFDVP3JtU+iE/QkjbOdIPV7Na4ErSEtirLZYw2G
L9aMbJQucOh0onxVnjPCFZonEK4IpCVaRsZxArPWPFwehjDm7Bem6++6dZPbF59S
we0eT3gfhL4bHbcP3wr6KGFA+XMAIaQOcn5Pn/6cg5rJ8yn3MKHtxuI2BIAAKFIs
5bN2n6H2ccB45Ue7zM+9QoJ+SMk0lPx23qIzIvkzxsTcqfBwifq/+pKrlrpZxl/4
NIkATqsScLKM5SbxXIotMW7aqi99wY5bosHseHGlZuLdcCZ3uGmnvMDgqRbuHD8D
lvSXKmoQHTk9CnYuYFcFVClrdizpjc94lIvCATtVCmdB7ZZZEUEM6LHmQUw1zQi8
C3buS8zGcd3/qNSweOCtwH/mY904FiYKbXaiK6VLD+BbeQJne6cg72cbPkMEVbab
PLf1l9T2ADfGPJvclSwDS1wvMNI0RJzFrKReSlf8iNk00d8Ewyk9nr7tcBC3EpZY
XzYjxvpHiT7qnDJTpTCnNU8WhVJp7RPlnVp7Zjd2rz97ZWLcSeOm3RO0Mx3LGhN1
iDQxYGg85NQiLcKnduC0badxXY0QU04BtaiIZr5Q0804QPR7aIlZymyGB45PeMgz
1dBqcu9DS6iPqotxqydg0QAs7yh0IvA4/Gy3YBxi8AU3/nlbKL060IPn3ZhGZIFZ
k0WuLveAYtVP6nCUYFamuSoigN68Hnm3cKnquTSavVQS0+bY9uah/9+UwKmP+9vd
LkDO80lGWwYfRyT8fldAHKeBpZNA9GiqqrmX2bVasMa5Tc7SaagZ2u86K3S8N/vB
q3mhr1Kt1YwctHY7AW888VZ2tnqIhUJ/GFUrjLJmR9S8NrMRZNvMoq5ZDw3IAriz
mu1agcAIKqwWwilxcNJiW+lu1JLOdUwyVJQd4/OIjURpmAU+h9h9Rudl5A+GfAMv
zMtp8XVSeE50sKOM61JcwuxRjnCBKK+qPS1CiykmTzJn0Qa+/bUec/VlxSmJfe9e
kdZwr9iffHEqrbkO0p39Su0ZntZ7cQJ1OFV79LyF15TnihVj53ZfQbJIvkkKjDbn
8cVWvx951PJim0NnzOyENIVUV5SgOrhmaYa0YRfRQANkJxMPz5nA1LNn9x0a1JRx
j20R7SeKIIKhD+DTDK9t3jR0IVZydF7m7kfKxbHZlz0v6eZzXpUWnOAQPS/f5Rvl
s9qX3m7B3FRxEzCkfg9eNhnfz3vreUPLv8K8cOmu1MNHX8x3+5b6Q5UJghIr4nR8
o3YRLG0jtnVxVZuzW1rG1Af1Yo1uenJ/gGH9TNXvl1ALBb2v9Pc3kC5jmgX+JxsE
feaQbzw7O23WAvyJY5S+BiOv6AyI84V5LW1qqfsh0gg4aXavDHJaeAI+x6mFAgZe
xGGgEooCneXtVWraNWiV62IqfrrZ/CcxIn+rZ9UYEeGguNHTDCEuUaWPvqyZixUd
u8Ssct7obhjc9SVzAx7x7ioKJfsgvsJaehbtPNfX3LOd5eQDT/qg4tIIeApuG0Pa
Kaws8TlN75HWFBYOplIa4XyCufpKXZs2bNBtRHACRlfOgIa+FsUzYwIXag5tesp+
jgxgR8MgnZIHgKtfwob4lsDc0o0G3renZA7+2fSFmYpwKm7f7rPxLO3GR3to+ujS
h0MG9CzjcfURZ99YAMhHl+jCQn2mrFbBeITZIpJMSM+phDgvhDKXSi2nZqMcUYfu
mM4/oa2SUZI4UZZDAca/SxKt+Ofx1CwU0P182k5OLOh5dXGV1y/8DyL1dsKow+8N
r5IIGqTnUXYZ3VFzK3IrT1Itsbu0NEvPQ4/Ejux/dZigifRnH213hfZZi/HF67QZ
fmvBJX6j/kj6kSp3U+iHDoIMY+FDMgy9+/uHpJfa0nHRokhYyxUbZlMyslsDRM6p
MnzAZaVgEeTUUDPVDwvm3m2eUfRNqzyTEV8OzWX36CRr44uh5kTrqF0Cw0v1Qqdu
0taT7swK4MtUh4aJR7pheI7fEvxcg/6aW+cimSDVT6mYrFf+p9Uf+vrKCJrj1dKp
pBEKTYziOT2ZXWsKodE++PAQXakRW10OaB9J99poPcq1AYiCGpqohRk3S8DnfFJt
whhI0Yvct0DPu5+5HNvdTLRnLYpky3H0QyWR+ZYaWh6eaG+VmyU+4vLRMfqvyO1x
EfnM1Uusz+0/9IqqlwkG1mT2LmSRTf3C75BOjQrjgP8iRyXNus/c5DQP5tvEFlWk
/2N3VXRxn7STube0etrSyJ5qJlgV22H5a9Lu7biJIl8zB3oKlPlAWQDNGBr0S6Oc
2JyZs2qHfPE3e7vCsbpNsV3eKXPFSI64vOEP+SH3ghPcHYlSav7iL+QJdimywfIQ
Tf1DnJQwu69ozVXOsJ4Je7tRlJyJSz7X0UqvIA1Fzw0Zsq236JaBgSVexGaoERkq
jmpLx7a+agVGiVmW4Xfdhpd5+k0jna1wUu+zchgefM9YH3MLQ+YcrXsNT17cJE0j
naB7VhufP5QwabuKkiNzD+8oWOdlGSErtamJRk6Y5+Q4kIdlm9G40or2/SrKxolB
dDmuMNA6YWz70kR9Y2bzirvcvm9ljw6D5PYFaMEwBlwSS97cCDJkJvSw78RRuc0v
/Su9XgzCiYprSQ6nMkYYqB5Cf8iHOkHO9LXiMHmwwMCi4VLQYsrfWJffIjJTlAXL
BzS8l3X8oAUSPJQiRsecdG/rmna/+vyAdn50FDhhKteWOVNKF1gPxTKxDstLs0Xo
KypHlwLs1No54eJxu4jcWkQhouKTqwxyoHEIiPh+M0+ITNJtMxNBPHx06jAYtZVw
zUrxjTCz3atPSy/HKYeGdMRltAOpZ7dIa8jS7ttQS9LOvPSSasifQOcPNre60KCv
1VWVogH7svfFDiSeYccn0NQg0yqNyQaKGNjH8xVxq0j8zWTd/QpNS604ih8jSAhy
l/vkNVOUJZnYbwinQEadimMypRUyYN3OQAgzYtSVyX+rHnN8QHzj1LjMeBU/B1tk
mtqIUFvvcBCfZAW4c0bJhGcjIP047hdYNSyxD95vKWbXmhqGSHLkWJvKoKnBJXUO
AULmhuH5SU1LprSAUSav8qClnhdRlV3opCUGw9Ez9PLwkRCL9+aZRHzR3IOsZHmY
jSBc9WUGjJHkxmm5WsnA6favSIXJyBbtYv57WPuEh5RQwaW1rtoHZuK4TmeH7UvH
G3WQqmvWsYNuqiDDNUpJcOLD6XoivBLtWkXqXWPUE4cmoaVfwKBjfRNNIDfnH0LI
N41pv16X1uc7YTIer4AzW4/Ho/TrGXfUIsULk+qiJALLlyk0DJl9lWd1t86gSkg1
37R0QEHReSYp0OHyDfRYAOqMgAYWYDnL23qMdscXjJcgWZT3kZH/lSD6hvEUlYcA
qAyU38Ukeap3+FIMDzNsnk0If5bkXmbdXlVBI6HXPF9OPa/isH4E/BAmPkKHN5cN
j/5IkOyIT+YnY0ie1NfKR+0riuPi1hBoZBDVt3wm6UjNhrBKko1/FEW9Pn77UsfX
shL696TaBtVjfEY4wfvMpTGeFYYihFlLkBdiTaXrwYpgNueSKJuv7n6kdWOdMfgm
cDMLzzD+sWZdGUXLZPZ2EOjMYlDogtT98CfZtsta/LZzVA9OnEpG110XFL174Jx3
4045Q/8A27FzYjECpVPZP3n1QGB97+Q66P9xh6fXEIWLfARbi81n8/OkdLM+PPzH
X4/eH/kzLoaAYiymP/wpSMCQJa6Mz/1ASd2TRi99VIXYSx+NyfkY8luns4c+QJg9
QedPyWp0bJf8jVh/RWXQojQxbs6ROpLGTVPuAgQOssrPdUM2gg3H+IZdaicrmNMA
nu4Xj/Iyzpr9W0uFlnbVl3qca0NbRvHOZv5E2Z0uY2ilVqyNmviqzc/TwMp7sRva
tRJd3vn64K6mQG8Hz2neh8+7/yioU8Zxrc/IBG4gIcB/eHix4h6dKI7FS4dDxNoJ
jhsKG91lnoatLSSVn3hOy8DUSj67YPVPCKG8BbkVo436OW71bq6T3J+0JboGzEAF
99E3WmoNAt3w0YVlTlwuSfDpJOM97DFUdaKFEvq/PUey2/ZtPatSN9QpFe4CTh9K
xkSwdhoMITe+v9yhl+JaBL5smqxleE3NvxHMlDhh8Bow6yNKtnqFHd1OzJzH+LBf
FhRx99RouMSf23PvE5nyfjO5K8DqlVmaNTn278aGTuuFijnOQZnmwXNZ0ZKo1iy/
4orKtw/MMOK3krqyrnm/WalUB6IoNBOpPFciSHQCCFniUSHg21z8x5npALknCXLK
qohxUlGDHtWDDog3lzPjFyFMdWVFMzHB4yYxQEc6I9DnL99Yw+H2LtzJDCxRhPCI
DPFfP8mrOKmtbgf9LxvFrlxtcH5er15Bscs+fhLf10Nm/ZxzLjI8RvANi4K7JVKA
auWghpYAxbfeDP54xWdHvm2UoXlqXXOejiajigqffmfpOW43xKq+Z8JILRG/2jdf
cssWKlBXWFqJVCUYSSgjsj+k8kH7BTy+dQWFWl8h4Gm2suekbkQ0qer045/2ySfl
6JW5YHmeSweELotgXkmT6rM+JOComH/YboVCdIv1QFVxzWrflzSpag8IkegwA7WW
uA0LTnCrwB/JslzCYTK17Xg9Y+bDlhCeCxI3zdWxAM5fYXESa5YmWp7qTPBJU/Kz
1IavPZ1yumSEXFr8O1m1QwJwNXjwfy0yxSuf7Nkb2iyrzYEZ7Iqh8jkVnYxxjiRl
K3/P9DnB/TNET9gPl+s+YnXpyrcbaPHnyi0I4fyPFdyzQlvSpXWGR4HPNcRs6I+L
JtvrEpxjOPY9dGxSB6TCMQPaNuzkqyuC3NF+XdZG6oPkzU+wxkvLwPUbedIZltFD
UB70s7CKTKSip4qOphQcY31CMb//QK1/54PU2A4T+EItY9iI7P8Nk9T7/r8wG1Jy
qaIS3BrxopZ63Bmj3dAhZOFzKEKW/S7CQ7YgGJPK+lioulnZfVWSit0IuS6m1up1
O3OaOCkZiUxxnI20Fif+z54KD0AbfxqNPhQfmfgT8qkjgNfBVLjOMzZIAi7TfXJS
vsgA1tzEmlZSsG8isTzcXhbx7TcEnacPCdElR4Y0LOYDRD83Jgz/LqzXYohJNEJd
zP3/ko399cAz/BZkU5dlGxM0hYVV3UxJVBL8I3W2GEP1Vx83HEJFVPvr/27X4UQF
QcEJVKUScxClWNk816i6R6zgavM7CtHxoa/GaU/Zlwauk83DcAfmyI61EDB5jo2a
WbWnGhk0NG9qF6SlZ2vVqOa6wJMj6oUm0uMBOQ6979y7v68Pf1oa5eEjWR3AChDj
Vw2wwI74lxOrpzdmsZmJqy/hyq4aN0cKjEPksTnz/U4z85mli464eypZZ9Rrzak8
4OJMBqIapSgLVORnwgwAgU41mSSMSahRDU7sGwY5+pvaeCVh43/XxFmSXgBRfzT1
wQLFu0h3CLFiejnkisRU6MtKAVDoqYz7KBNUHKZgFM6NuasmZMCkP+ljXgg8Sfvs
1XPmpflXbjeUfCQCAs4P6FmQtX22LVEQxmeLelM8K1K95kMQbB/JMok5pzgPqkwu
NzjntLR9UI0SUX3lSiQASu7F+URN4/GvzgWqIqltzAiDg7G5R4k1nxme0yKU9pKt
HSZ+ZvXAEoW5F4nSE33Cm0Fi5cv8vtPOvffHeIeQ1hJnZTwwJGjm9JDtsO+bQtxI
KyWoldm0jn0m1ECaixZIgkSc7xz/B7T7qD4gDTvvK2ViM008X8mdsJXsNIOW2NVm
snsLFeVvQZ6AHBnK1CWre3LDHuIigTeQu4E/9vklnM3dZBnZBB7wJcfhMXS5sFDy
Dobju/cLLJNMmikls38KPSPgxjZChr3AqoA58wHjEgLFeP9Ry5lvqFmO9tv0gYLB
h4AyHeYZn4o29EgOa5i/qbt2QnaR+yjS8XDj4hGJ49Oi141cEGF0servlsSu5SZp
+eyv43g5VKw91rPdQz2P/HDM+oApVUo9DUiqPaSISEbpJvqFQCspWkKZ6wv2bSR0
sbi7IV7xBC32G723Sw/voS6drjg1hZDxxz0KVlvbGh9NX++3hWNNl91PY6NjIMjx
HayBY6ZFuGZEemd+q7GENW87skwBfV0JwuyJFO98HyfdwM+Wkh6ae0sYZ3+o1qOi
NeJ1lArNc8wKgvo4tHv8Xnkky6vXKBDkhaYibSO7uuvY2WL3HLkTNSLgxTN2a/ew
FKXR3sKGlXZiyOVJqMy510Re9nY5zuksO3C3YyTNQkw4I4ws5q5SuLrcq4XwV/3q
VLSqTb0KeZxSAJX7F0YkWXvgvykHr55IDLQ/OqwVB8IAANdiialMMtEM7/kCSFkn
r4XM5RWwdtQ7SxInqFH6fXP+Mbo3vRc6pyaFaneT/hyq6GrSGAY9wnInKEy4sGUP
AC1XGVOHQsD4sSiv0iAJTcxFN2TmjWbG1zsN3w1SIJ8ocmgJdEYQYZNv3E9jrRvY
wY1dGi82NUp9dc4nANN3lFwFlgrIkowzdarCSI2JNz+A2HZlWuGJjfOmpN5rQ8wq
Hs2/IXdczNDGq64UuCqj3g7RDFle4uM6iRjbUrtU0fbw0UenbCmfOJ54/chCdNSR
dnV2i6SUuGxarc6yFfk2fGTVGcHKZgF1SDOOi3r1yQC72FUc16SzZf2PjsF5AKMh
qfZXI+X8217UfRsuHT4ZHbRqR8M2Kw48Ngo3VTqaTW/e1Z9awe00qMl3ctUl93hf
eP1D8jQhSlmqrc0XhKfwwPEw2XzcGPgGeLJMI0a6j6r3ojxQJP7PJ6JXF2QYlCWm
Tnt9zbotFDgSGPj3LiegcoFXNequVQ1yrq62AkKsMPtfRCShbASDhbJgpiBr3LUl
RpW5YmkbCfj+zPSFR0mkFHYKPQlmBNbumpmuMvV1zSbQgmhIt8CNEq3kBmaKY0yy
l409GQRXiIlsnvIgWYkEatG8ha6n1g0s4yB24SWUYtQxvVVHVxVvPJ1yaaaEqouN
fhbz+dQemYnaJb04KxF4Rr3cpuyJedGSOM6nBYjy188mzAzQznf5a6MgrRqFatpG
vqajMnrd3vu118qiZ6Mr9H8Q4+t+hZws+20MPTSeDOPmAmBQTvkeA2H72mud613/
fXIxMsn8W43/Favg/wmWGzZMK8ODrTBIkj9xpCKCvuWveIHny+CZ2U+lpmzkxgqM
YoYk8qTgapPMr/FI//mMZ1OJdiQmA6rZJekII5IUyOAo9n6quIgvBTb4OtnzCGgP
HrxlUygQgJYWS3lu6ecclg2POEvbIi6kwIhrK8hw578f+J/ZknYMg0SKko/r8Wmo
CXVkPNRzd6st2/VlzRcbIgP0uFTPCQWYg3z0yWMxur0m8lF4KsEsh7iBkvPyU+CG
EhU14XZsaY8EB/6RIp/5+hch1b9FxU1G50Dz9Rf1Tiz27NF0fI1G08y0TXuH6zZO
ziIEwCluBRD48slR4vt7a+OHHD/GgFBGK0wdB5Yc+pCP67r1uLrZeigXSx9/ZBxr
4S0S4RcoE+IfrrJKRpsazYPFZf0dYvfzI0s2IYsKycAtJyerREXisInK1Zp+HfYN
V8JfXl3PeM9ORGo4nVTwu/wU+TVemvj4WBymqpFCfaQOm9dsI0mVa+4yY0oubE9D
9749b8CwlpE45rKqFQj/JCLLLbA+x5j67eI+iLqOc3PgzpZYWNDWGrXGWbzE/5N6
DvmeqxpLrqhXUoVyhzYQvjI0zRJLDqIDafn+JT1FfXeUxS/a9fvX9b3c89Ds5AFW
U4JtpD+fS2TbNdJ00MQYJzmBX+EwvDI8N9YPhcsTvEgUJfUWQX8XS0MYA3o8QVOg
DQhAPIZZws3kpqy2vbMeU3CnmkWIe8eNnXu5DpvIh4YWSkUMM85GbGo/AnRrWQdI
rnqD2Yaq4GqZYFPyqMfSo6UxszNU5MHSnSvkbcLhy/ZcZbKMJB9qxhONfyB+SwDm
FJ9GiDzJIWI1y2NREFDfTxXleYIVx6GOEm6RBaWVf5tom7zZVTZXy3ZVzN2+77wt
6JGoR9E1Gam4S5TpG09L1EOwPeN1DvVlg3GCPJkl48AVzpqORb/eUH9oxVpY+PXA
a5HhOFOKX/FpzQEAU9u1+S1K0FzMSGR3xHANtPiHGaD2k11HxhUs4i3FcK1wtu1i
OKEDA/yPiWiNF/9T5i0oUtJo9b/CFPPu9G1Lf8naBT12sD0IfURvEL53zXQX0Ywx
+4kujimu0Slui08I0qNYby3WZ6aOt7WRQwALBUwhnpQrqRR6zYDK2ygS1TtTO/Ar
zMhLt98DhKEEevy9vTljjJBDmnrni/basFwWOWqnt8LbLj6QLA44K+lv4kfcCG4e
nbO1QvyWqk80e5Uw8m+Ze9MRRQ3RKaM3THlDLZdfnwlrb/7h1LZQbBuZK1iTUj4s
IA+wDiS2sqp3saj6aTX/7bFU7yUAACERJoZduIWlKpwTdUqX2cdBPNLd782GOXes
H1N3NYED9RxBz2DTsj8DVtHjMgim3aOkuAlyUPt/oBO5+2MYflA9FJMleBPFv2cm
aSTpw7+RaBq2qTktuDv9dD8V37GIOu1Uj4wNzEL0gUJIOelduPB2FXRDrQfMreaB
xwVwyha1XFyDKo/21M/bmO5QXkx6fKUtJGH95e4TCv4d4NVKwFf+alCXQmpgljjK
qAnCvYEP/MT9kgJigLWQXGOtj6SxsKQ3eukqadfRclMm3BBy2DPZDNggS8ZBNY1+
UQaUZC+6goaKhbZY4isXr44qIKbMqosIQC6uei+h4e04JS2YgvnLrzB3HHCYMyUv
rHr3QhqrrMmwv4Tkb4xDXCL9leadT+6k3LEaSoODp+RwB/3DR/8s7yCn2at3nY+C
OYJ3iN6RF4/OuhimFxw119h1/kqYBO5PC3K8PgGqxcaR/QJeCjIbie0ZEY4/luIx
eFU0YCRbaIUAeQNKWbDMj/S6zrkVfyz8KxCDJez0hf0NKbmf9a3moChTXHkwmmxU
oQlozRhh99UrB57V3H3lorX4bxzexGFCDfaa7WRDGCMJiZELPDTusQIpOX/+uYtd
HEav2fhrfoNA6ui2N5cnE6CBiXXvmgJnF41fioOgIa07jC0TWYdEpgfjiyHo/NKW
P2sTb0aFmhrAqnt56Ej05FUIwMEIVDIP8yx/83DEy6hOedqGj4LfJALbW7WmNTEL
ZVk2A4dXr63Oi4y5IjqiaJtn7hfHjmNJ7zbHLctIv9+mKPM0Iej8iBk9lwHcApUB
CaJmkBxqlFPoVMKXw5YggrMKh0C1zMvmy4EmWrcidehYOiT4nEFYxrsJFbvSglTZ
+Mmi00Kp6hXWdNtwqezW5Xd97ZVe8o3jkERxs7ts1N48H6r9U12K044iaQYWsHvm
U8+6rxRRfScfD0C87UpiZnhxD2/XA7EjrRxLAQYMDDRlMyvDFX0u8VIRclx+tbwm
O83trGU9PWi/Jn4xvkwb6crQblOc/1IpgEp/0yZhzO02iMX3TSq3P4FfsnWJdUj1
i+JWCLha/I3y731lKaLd0yBOKtX5x7YS6U7+E4NQ916gSocSyyslxe2Zw4ZMRY94
l9fN1lsAcV1TpJzxWFlC22Etdni21/lqmbrj7Hi8kEjDna6oBw6xVKqqc1Ylnh9S
jNyt3ule7yC+zGHzpjc92AtBmBUnno5ArJ2J3yuRIrTz0z6N2L8jxM/cEzGiZrwy
Ei5h3kvE3bfpkLAhsjmSOri8X1QB6mgMGN35nTbPr93R3YhQju2hEhPiwdNFMH1I
A3obRz+APpEOjwC9EvSn5kc422LMpI9LH3upUrI3Hj6KgaetRz92E7Fgfm4b0Xob
KZYMRjnE5+AhbQOBSIcIsbqC0cahfn6x6CHuDThsQQFMRJPYX2qABqzEfFAGC3px
L1lasn+iitxH96/yRx9kosVJs+1JejSyYtIR485xPz7I49rDyTO238IoE5aFkXLN
EUvrhvrqtO5H4yqUe4EW492js+IshZ0bAoKy5fFIm2FbeQiiM4AhxHrwduFFRO2z
Ra4AwMNR8Z52BiAFtBeTwy+UQSJDAQ0L/Vd2rxA8EoudGV7UeDCNnNDn/XGMaOrX
PgltBgndain4q4bA5igS92IzQBUW5ZZhT66nP9db0UFSEVhbXOPN4CP0SpuC+qMr
p6YsTTOrDgkzYwQFRJFMc9n56snaUdjR740MRGcJKPuCi2lK8gexrLHw7BYrwXix
h7aiaNQxJk8/hejaZUin895K75GMJ53SQFjMVQ1Vwx0pZWigD8+ss/xr99oVMQHB
o3vfoSCv33ExYy5rH2gxOUlcwY6tOHmht9QsK5WBOWAn2Z7U4wDX5jRzDRAByQyt
hMs/Dzc5dk4C8gTB7zGTBllGNJUQRPIR1F1GGdk0u0v6G77mYcpdS0SwmwqSKoz6
SPJ2Ni/8aLsStdE+WrAUUXONWzMrlQdEd2dptlj5Uvp2rTTETZRCazzAUbE+V7RP
6tE584A9uLXpHYthlP2a1asHC832of20BmKaqM1fvI7lp9idSOHOTFp4mBLTMi8h
eRqLfa0O4crVeof8SBCS2vxUPSIdkr1oiceDmWLQF8PcaCA6Cu40S+7+AXOSN93c
OXdD25Qm3aHPbl15bnFvJCHebcmFcxW6aDttG4fDbbFrMedEFSiBqQys+QrR49pS
AmJObQj7gEfwW2w/GXiaTxU3kR4NLQVXh7B2Kd6e3PBfDmJvM6fOMGqS8pBmUbyM
rp+goBJqzZyk7ED8XhS4tLiYyccWhM/p8cRtYt5SZMsHGuYeqKXzS4YOCQIySnHD
sDPwGbOw9Av9cJTj2ryV2wzLSOjHfBbmT/lcZrarQZ5QIo4WQHaiKGUSAR0Of7Of
N1s4smq14H66eqPGW8ZigpIM1TOH5HJf01UfMARNyL1/vBEcNLzp5MHwJnkjkeFv
RmijxvWNrZbUsvo3927QNhQKw/ClyxUKj3jRwQZgacK5HbmazKRgCBTJhjZpO9Ik
Ux99KNsL0AIkFcaLuUVeFFm8bsYSOGO5xrwQ6WaPXyMeXKbq1heeqhRusQSRXhQg
cwNZnAAGlwoyN84sPnP4EfPy5jN20jWI/zTb87MTqQWpBdN4f8UH+VcTEb6fmoey
dDJhh1mpvuAqyEc+uOti2nqoXNYYQUVrNZDozWylwq19x9uQqwEHKYlMnQtcsaBJ
aNF0qXmqehkDtiu7AAcvThjCf24XIai9OT+msgqDv39TAiZj2tbqeDM4eglJGrGC
7Brio6KQ4hETd2Wf5V2oZZauB+63f5oWTegKc8rJaJun2G39snHdG+y5f7KLqYQD
5j0m8ysFp4rwzPTzaX9A8NY6CJgatRRsMWGhTngfpFfU2TDg7jM0gdmyLvkHZDju
ZjzpHU3y8do6PfI4CCVSwWG+PSWEN14NdbO5R4mKUHAEF8KjHt5Y3aGjhRp2Ih1w
iL5jP3MNZK3cWN64ipzhoPy/ch5gOahDSNzvUYyyPWRTxKKm+AgPCQr9EpisqLt6
qdXsn+tfNpABujjd92Dr2g3sFdqfnkLKLdeztvuVgyRDG6X3WsxXfUbzPOrMafrz
e8tRLd9TpxV7VaLNEF00cCoYenPRYMkxwHsGfcsZF3LdlIi25rZr/RkfPktLkyi/
gzFlof+nGbMSajQPSwb07WWXQJt93iXfCgJgkH8bbDHtj99JbHMCM8GXNXbJBpVI
mlf87NU5FSErWdJV7JzW6MLmcrfrM2XIjHrfvmdNmFqaws/WLpzs8+H+Z86BU5yh
QcCC4SHw4nr2d0uhXUSI8rnK885Vy1ftHOSGBcTYEHoL4Gp6ZpsVRe6KgA2EEZ/Z
XETlslPiaP/Xrxqdpi3MROvOQqp3nX3wpMphYcJNhaORfZvlsugm1K3XPG/igZVg
F6W5NtOZS1CLIop1yo42I6iEB309RZQAoh4IKCjr35LFd92J3SHnGrtvQr7RZAbQ
nhDpW6YTRDMNntdD5fNshHQf0XK9mAPTQZxlnWxh2NwhPh+6LjR42PPeL1wa/+8t
Cg5GHVBY2UkcUSMczI5B+jcD6hbbqCKNCtrPMZnCby47NbgkAi1Csk94aeYahz2b
v4oN2xCK2+VsSI6pHG7ub0DG+CGXwpMk7NkZ2j/KmWXCSJwPCzeT/OyaS4q+pgAP
I+jjVYdWSPy7SH332QDVZAXsMKYwlRa6hiremAmhRaz0U0Y9jefM58qIy7NOwXFP
2lt6jIJ/kVdgpX9jnQJsaPiEWNFqzvb4zo4rqk9mL4vkNM33iE9y9O0yjC2NS+sZ
kpomU3fjO6JwPpPA8IZK+d65PVDdfACloKOg7Fd5YjrvC/f0SAESZZg89xnFPHin
4NbjVBj4J3H5S7bitCFVGprfgEfupeoQmtasQZNdvmUbk8mRMYxqvQ4Ns9Ol7rtt
4ESNOiAKxX+ybNRIMN+YMci9jbNQZkJ1gdWm5TJT+hDKkGAH0oem6XGUQTxT9kf7
Co4j8CyQp+VVENNouqb+U8lB3L6zRuKM1TeMz/PIifwoq7/APJtwHpNKKQEU9qV9
ZTOVeYfk5iEA7I1cnUTfSWPf+vkGcIad9/HeCK6w8eq09GpVdXUS4tiBApsRK+r5
gEZyAZQO9s7qA5eOt2HCs/yGd/y83aSGCFxyxto/gtHcYuL8LjXyKnaJ2hn8QN1X
Lu67le3rLy5HlAiIso7OMtVBHiwcWc6blxsmOrMYRLkCTel85SNK2VTzfQAAGutO
zN4lyQcai7AEx59IfQQkCkrsEHQURutUWqQ5YfAzl7fbB1PAOeV1PDUuuyIde6jY
7NiCmfIiKdmkjclrmEn4epgCQ7axUg7eGlogHie7KzcI51SQvgnPNZuywDF5ZiMo
hd8d4JSy3PIe7h9FZoXgPvFubFIwFp/0iQ6SIHK4WHGEpE62qmSBK+5IjPouvDma
8hxdqHCbBICfa2C5PHzxnsXQA3ctEsIqyUoWN61ewvHfKxWuGxpyAH9+NVY2i2ll
rhPefFaarMvcHNdOjFwy2C2Lm2JLSMtqhhsCGO7/9w24TtKMkH1RlUukboPzadvi
4J1gx8hcqPDUi8xOb787XqlBfeeQWSBYOn1R3vFSYI6mw1PbSrWoc6fkydCQkwbg
pCSmJtu1qffh/DhYKukaMgixCc+EJpnDRFPnh4+CA8TiRu1ChB//vjIkO2VU8So0
3MnZWWu9ucYimTamfVMc9inMoOqOqpJL4nem4Vhd9LSjTmHEUc9MKtpDA8KpAc0V
AwBtrTwdQ+Pxb71naAEi61Y3AhBLPGALFpnD/3XoxaX7gz39JHEIkMqN99DGbySa
eVDnQC5uGvkt+YR9pRES313oOH0xJ3uxRuieEqOIZ14Jcus/MWo2a7vYS3gl1crK
XQqwTGRXty/wUYB7uUwpeBB6pWPEUmviN+X+ZjkQN6siwPk1RPzVfinQa+DiW4G1
ZkkEFUYf7RWlV/Oer4/YBp7VHcq5rWCgGtDGRCwO4E85QsFnvhjAeBH+TjT/aGgL
RmX/J7cybc2XcONd4exVpNpce3j19BRM8KWC+fgOLFtnOjVJijcVicZzyRJ2azfo
PoL1mvcByjErxan2ErnSLryPTtrsavHosUbxo+dDWLlwvpkt8vRX8eeposxcaPm2
VUahGMnOnrco940vHaCbD6/dY5zRfD8n66376Dqr9eZAMSXDJ688hZhxGovW5Zla
MEmkLpKpUOZnr7a340ibk0l7dztB5PKJQdlnjn5+LCy5h/ukCZExYM/69EBR9gDH
pOMzP+1VAoaLskxRXFHdbFcfg63dic9kiyeoiUuxjGB4nMJ7pfL/61vJ+JHEDrkB
sgX0cnS0DK4NLJWjtE+m4AbhBpRNg54jaSQqG5vk1HMPq4tcexx80s+jrwHnm15g
ub125I11EQBUywseq9W++o3tLS8Hog+ITDzVuUE8Ikg2grTec5dXdViyDHnGqeWi
qCQu2TpL4/hJCQxhuX62d+mJRxt4IxTZ/ezbN+KhkyHgighQftiSmSF88tmHmAmH
cs76ifPsE5QmDasov8ksknjLx18bkmsQi1xcSwZnNJST77JUc9abj+ZZTFMoj045
zR/uhVT1qpiAZuDsQIiqVE6OafFKxyvcb4Di2ua190AR0lHMZUPm4XcOqFaHAfDh
QNfktJidazbZBWA45YeH/IboVq5qELn9Q2/CvXJCKGj2Xw5rdu1VAay9HdfoI/a/
e7EPGxzpLJGW2mkc1oxBkvkF8wjmERoL+7p4wCcW2vVChhK6TLtrE3o06KXpX9Me
UwpWQGAxDgKonusTlrAJrZS2xef+gwaJdFOLqvYhhv4Hho1n5gX+S1r9UTNcepbC
KY3UmnLI1xel0UxmuWi7eGoUssrSNzgEREuPngrwlfMr6TjRJU4r61lpc/MqhgiA
cv8cc+KyPH9SGbOpYXvgyJ3numLxs+ISKVbwJLoA2QV+U8wmfnxht3gC5wlva/CD
ngoExBD6vQHLx0soyDG6oXfqUcfDK3ElIJlJ+e0Exk9bK5oPGzvTaX5a/Bn7COhf
7B+uTDgDilxCOcp/4eGU7ivFhTur+EPmR4q9h4lVNSC+4+CMRsTpWg88NbB4KSjl
zz5yrmQFRs4L1GJ0/pnxIgl5JnMttnMKtbUZoOnQadpS+foj4Tn3B+86f+dfuO/O
LhOQT8FbeKsYRiJzfzfy77PBrtEhe7R5VMffJaeLjmf2w4FsBqIKmUMCGE8afR33
p/GCApQ46RkTYh5jHNg8EBpkH1rpTG0XXg7zMQ7ULzTNs5ll/Sg6lLqFkOBQ1Ad+
Wd1Hto1AhFdOSA68wWUfKDN8Ad1EQ3ikBFhX9HLgMVW8DFDRPjDXWq9ljIXTi6kr
HsdNGqKGmfoQ0xPLO7nvktCdaucZEZVy6tAcLhSYz++VKKDLaFI4esoeaS7fbxJ9
MW6Z2L0JcBJNDLTZd+VKhXNkwojuAWGFgDfzjUrRGc1cQHogmVg2S+51vZcGyvEo
rUAODT5rVXYLUCstat4wJgQEQzN1/I1/GFZDGa+NrTiM5vwpeuibXf/TaOw1gxGv
Mt4FMwehRT6nDpS0G1h6xSZZIIwFputzew+uYT70PK0FEWb8IpS4LllZgPUend+A
41J6l846WKA17mJoiZIGHcEUXIpMZnCdrHPWrUo0X6tRMPPIJgmtSlr7+Jar/qpA
t8VKODI7CFU+9V7Xh1FCY91wxJnIki+BoBAD45OjzT/N6fttrhvK1XuFGzj2kEmW
UXc+UZT7m0c9H0fY996Y15up229zKq1dCL3FMaH1YgqXKaWN3A7f07MBCg9Kuo6Q
wdgyDmDFg+zxfKsdYqWaPwOnJa4KLNvchS9s1u1htGdRGOBAvXvpS6xkJQPM9d44
d2i6cdxl+Oz9BVtpLngBPWmxTYAU+NKutEHithZmujCfmqYPNsSfxeg+tNzO9j96
XA26l8gJnXAkCLh9lXoxcexs2hlA6kNjdq6/dhcQ8w841/JsPUAIoDBtLyaIUEku
tUp5j94fnA4v2J7ByMS0x3foF5IFmCrQ+bBU6z2HvZWkA7wRUhf04IoFvmwyfNnV
bu8b9REZzaPjL9WoFod3it9B+TKr0BzmuOioUPLVDuQ9sdGmIR9VShhVnPLBaz5z
PSx/odtzrvaweVn+SciRXW38sBYEp/a25HLu45Gp1/L1VQZl7UpuR40ClAQfCwo1
8kJ9iNcj0dvm1R+zjuvbZdT33Oie9MYOXB0YnqHElt7LihkTPoi4ZCE3vMB2CeoT
Cqt8Ybfr+ik8J7a1x3Hz27BPAbzrmqcHrzwMkLKO3hyKA3V9XusanUokmrurrB0n
CWzyAAB1/YiYIDM3oLsz/ViF9hc4XTlU3oRAxiFlBp51+nah1ehbEwRTz4T7bdtB
8lFdcA02vl1c+JIHjB4/t9wZdLY5LiPOE+imdAW1n20071rusAZASW/tA1/scnKT
p3tpi2d4NJTJofjklaLedXZ5ICde7DXsda8hUlpBKN5mKHgVYg/IvphBxjoCEFKc
FNJZINyKzbtr3bRReEUgg0hK1TI6tbNyxRpQMAubzTc9j5ToszKNzWPKT+szgH2f
X/1Lf05QNHX9i9cmT5tcd00JwNVBbyf7jcEd82DGUeQUWkEkMedI8nQvr5Yx0sU4
1EK0NmrBAK/D6CslgCA7ruOqpcp0CCI/9dVdB+amCxlZeLqo4DnoEVGkmL1gScrB
/+0yoXh/kwt6MTy9r373oxd08bAqyI+9LSB4znd8bZo4UMnEvEbRMMTpxLZMdzI7
ISwFOVouNZDZHpHhXkOj8cC1n4lLHS9fTeqxZtZvmESlc6y+Sh2oCPTbrdxqZeXg
jYBT0AYR+BKwjqh+pzl5994E0X4z2vRrHCq/wGMOP8YH0YRuDVFhx02oBChrGVGn
E6nnZqc7PfYacgOS/DQhFLtjUromK0KA6Fs8UhecIAbA/KQm1s7N2YENpyzWFzci
942SPQp0CeR8JIB25IfzN2TnvM0HLZ29vopdC16NTS3eiggE0dbenTL8kXzRJU+u
ut7480waDGacqtb3Pc3G/+VqNUWkILiMVjdYbnEwdwHsHTBrqKQxMuv7ew/OLtpm
H5hK4OsYT5zYSxEnTq41AIyAFwOmLxjEOkxj8Z6ZnuK5Ac6iIMHZKQ7HU1SicajC
heffpb79KHqTbHH4tozeTfsJabvvlNLRkvCZY00xqWr+laMOEnu/YGcvgg7dPJj8
nkgLBtoyPFqVb3uJRSgADaxSaudLSiAdaOba3kVU705y2hp1eWJLcbC+lUg/tdQJ
S95mV/uAmUrIbhOj6L36ZfnaYoXUoIyMzk4dQ5vTnYv4Vi2FWUvMoz9zViBcjpou
zWIuEmy4kR4ozs8wo1GOKbDs/GDW9pCBRNgqzscjcAWKJ4naPRtfuRgrMpCMcVEL
N6QKztKVTOyPK2smmqt7mSVE2K3aMi+jSvXpPjksWFINQR0bNAeXilxOz2C8bqhY
IV0hDqFMve8fZwmB7ngwPGwAFNWN59pLcx0KuOT/fA/iCDrWUFFo62nGq98wuROh
yz9MHMe/vp2P8zRxPsWvW47aohM5Oi7GqIAOSqD7HoC2wsbEWbQUL3mvNha59adK
RqUT20gi+jDYdqIY8kGqHfTiKzOV2Cki7azHFRrUzF4crPO2l8d/gN5b9Dxn84+N
SL/G9yMH5Ev0iapHL+dNI0TCg3qFMPLcCt6mJf2TyiqNflJ1NefuYlqD4IzA56uD
j3FuPd/txdp8rVmv7cEzN04F5eShPtwtmKNIV1g759XSHMB4Xm3aQDrbj7n0uhKo
xPToYf7kmyi4l4SzHd9d3AyYgx0XxSUi+CgQyReanoYmChHAo1Aol+wbPbkqturI
2cQrcf9Kd6WEIPsZEGFtAKbE71PjXcieTVBWkMdGHQOEw64aZCjwPr3/r5hGk87e
rSOB2sHkQ36tInc+eSiMvTInTTzI10d7ChaUuEPNLgTy94mGC1xOotJSZOQ2G2di
WX7VNFsKMk3CMJ7X3tVoQg6C4HL+6waVfqYLcGPI27BfElyGaWFpL2jvNxDI7QIT
aLQE9HH0BBb2BVy0WgK8hha2Svau0gxqbDqspjxYau9bq2Y+jWuah6jHxq9Sd+YF
YGeKfDugpjuMRiE86UaA/uhQbIYgOJfBTLwXCkbps4MLtILtg4uOzbXyquMRKlaQ
r1OOqTWmnwcSJIMIhJ9Up7spGhn4EMo0eLzvh21oU46hVyAao+M73SO07HUqXRK2
3YsvPGzumAmzTC0FAW9uYrZyYyc59/V35C1GvUHu2WSi6gn9F+mw0ybQKtkMbKdP
4NZB6Nygf+Ptlgud9rNzvzL496ko32raKg5q5ZAt859OMrq8CvG3Y/OSk1OBYwg5
WMxobq/uUnPzBSEPcZ+jc/75NgPMpE2XWQkI/Fz/U3E8gGUU732pIQDn/U3L7QkF
M6kFFNqby+qsOWaDKDy69pBYDNc4/5+zlEwy1Tk4q2swkf3S+xj08LIZB/124F0w
EDizcbvVN5A6u6eNc5gkqIg2C7SO7U/MRqnpCECCD+iRJh+Fh7Jnc62JTM9oFv8C
NaRjrWo0SLqta3gYvLucqMokgJTU+0X8jUxxyISVpaOcaiBY0j0cH7nM1mzPC4nS
hggyeQKU1SqYnLdIIE+uNYEHPmdvn6XTiMcaw2V4CWoafpz+HkOgcR4nhcoPpNN6
HXbm3++7QpukV5Qhz8KO0P+NJPFuP+uvNYnhbL34/RYzzqRBY0XlMLNmBdBob1o8
crvo8JKDefUhRCyecSiKnoVRooI7oTCFDa32ZRD3uCJvFIh+ZKOd7j6i1aFAJWSQ
yW7ZuJghJbY5x2eMs/0Cm+xgJhxaqTAVv9j8RoFO6jnlEQ5+kvYCLfpItGEqby3a
PCKirn3dkve5ONAL6Xn+IIGMcYjyIhJyX5VDI8ggWNCIOSWGHYK+TJbN8Ja7AMHg
gsq9hLPMKG6F1g4Zv6B3pvzhDWo4u8VgeZ+zletSiYHhwY4X552NrdQr5Y9b7XDX
xsZDzIitwkby5bL0iErxkL2D2oBRjnVMq9VO5wtTKNZ1DGgFuv6ai1r4qAlSJuFG
OgGM2d+cYM9nrVgZtWB7yyoLtmDVTbFJ5+z6eI0gOlmOG08BB5I4ruvxtaq3iR9t
3UJyHVe1naOBQWMMEdj1nOSgqcYUx1PmWdOFcpQwIDeam7gAaElrwvXAmq10p4Ww
KU1xzf5yyOFWvBk/cXXdSKq7nopf2nAbDtPPz2prihB3BSNlcF5Ge6j3xuMudE82
Qou8CzmpYZqoTIOJ/SPkVlqqWZmynrxoBXtr1F7AkUJaarotiwBLEI4CEpJIUYUm
a6XI3kjIzICM0LmdoHXilQ4JC400xrc+xVUIgBKAIfxEMLOINLugI5B9/7F/B12b
sT5Uz6UtYXqStK04YqsFEEy+PgVkUZDWMVF0AfO0zEnCqQ3UqDFInXeaJXwLJOZC
TPDq3yLcjYq7zUeh5okl59BsOYyzOlAJuGMJaf/ReiYQ6wRY0Fa7J6rllROR8WdP
YNoOK/BVR74DTFbYUlY2M+aXxThKUIBl1U7Cl8I5BoKKtLpKLiSqT4HhQKFs1vsE
uETXXiFnSdGOj1Ym+E1HXbp38hQyPXlsuWHxTzxO0+cvEvGFtkYerw1GfBl+MYDk
Wp+mW8O68xJwMkXoORmRG/CyeHPrrGCgsZJPxwIJfobpyyXLMMi7eAsK2BbYR566
tb7iz3+4hcueGGdcMFl/qVOCSFkHdNHrnLuJtMazAmTpFTSYzwXaOrPK+7KPjrZ5
YSmGNi9tcsA139OjneCrTRPGtJVTOWENvM/8ugFW4dt8vxoTbX0PURMCJzg6GVs0
zN58O5vuVB43etRi1DAT3Ab5DHftZNOC0d21bs6AWgCF9AzTGNSkuP+kfZ/g4Wsc
xNaxKYLVlJvmCjmGyt37DNofTq5uqBSm3xb50tWGPfLuFe7xSLpLQfo5a2xsSTZc
mPfIYYkTPnRa4u9nro+svzZEIP7QH3K1WvSy0wwll+ZXdHw5VCkFniA03u6AoclC
+MyY4UctVoj87rkVSOzKt+k0knit1Zqx1bdEYchA1epoLapPPFWidscIyffFfd8y
ske+DTh2FhK9tiLkR71K9w+KuTnnxGt2dT6zJdg3hoYzajiv5eHD3QWi2fY60br2
hWgL4ELf32PzvrpLqQMMYD1zqUwsZpYpOldwdvw/kfzItG9B7tXGgXhsKmhPnzYf
hSyM/acUoiZg24SMxwCIpEkip00ERkORhCFs2wi8oHixofftW1ZjH8Nruw39aKgP
7eX7WWHeDXsHKIhgHtrZeYoGsk98K98mJY3ZL9LWlnrcRNl5XolEwgP6BGCSJMCb
eKtKa+wNVit+nPaO8K4rEbtFMamfz6A0PYk+4x1WeiUK2txvhMyqoHSLOvtSSgwK
SQ01gu7bikyroKtyRwtkt9KGi0dBqQ2ERX9LEai9Lv+QbwOl4TJ9gojPaV1eOUmc
KB5ypWz2sZA/mMpGW3bCYaO5gZz9WUCNY/AHjZjCedo5eAtx/w+NFrbwj2wPRJxz
WYuzRHjtp5DUTzNkezSuxYCiqlZFvCA6FcR0A0HMv9vg25EndB6tz3LCXtjCIkXM
rGyNBYn8+eSPYCxD0cHtdtJYO7KWntWddUAGQPuHD4r8Sv5jgJpE+YrU1B61a3RM
luDhoBptcQXp6HELs+SqztZRTVs3ehxTEOiEE+jHtRFQHYZHfsK1f4zanXzTpdch
KH1RKamI63GVxNDQtwwBNXuqwIpcX1O0vkq+jx8eG6GPzuKNwtZiQoS1jJCgl7Ya
74vaquszpSR277nLW9o9mTQ3xIsnQ1vmjUCkMYeglakJerbv6rX5rZOFP2XHUu5M
cfoSGviKmCeFybXsJUzSsrPEDtoMDq9u3CfKS0vGreVrKFu2WT24XXbG9pqjjQ/H
OajQ7hYpBd/mX9A2jLcxOnyTWwfOb4dNINyHMljYyoitplhQTQ5AIOhOD4wXePvj
kFzg1+g9A9fAfaR656Uk38KyeA1uuuTjaTe6pDkgU1EaxWGn62oeS5K0DGUAvyHk
y6L2uxlK/2rIvCHUAPFS4x7cTjByvsUoT4FTeD5P1cdGkQPlzRwiRfFfaBLVkDIk
19ttQXYZkVnY0bHgZM1/jQ1hGPTmIU/vMh1q7431Sdbnjh0BUg6whc7/dtGL7o+8
JxMC6rHzQXEbJOX4rGZ0y3ryNAs08I6D5t7ykLJevd/PVsqOYDt0fj/zxhEaP/qk
RwO/6CgyaGbLTgl+jr4ioZwGF5oLiE2joc3VtNnMy5rtbzBSmZiBwFtA6wBmZdst
eEtq6nDeB+B8josIJgBU3A9aE+nIXw6xCgVHNgIvrs1TWfD8aYX/afB0CvLHMH5W
nnkQvzE3k35/2ExgXmj3mkKLOQbahtxI20zkB44W3ejigRSBPTVWhagPeKZgndhm
cKV8JtdnYN/W03KMABgrrJx1rxwJlQqYE7TPZ6tp9fpGP8J+d6mBGWahnak0zAWn
Npg79FNj00/GCHvk8BekT/QtY6m3qdMNRGvQ0fsk9WCVkxVEEPb8tUsWHard8qjR
w0rdEMCXF9qb5fy+uTqydH7RYK39wNy1x9IWHY/lo0uB5Ca/VpKod/x2J/KL9rv1
JtRcQWebiGdL0uHXhWFeRiTiQEfFZHKcf+0V1ce3WRm8jADPqemq5hUAtKMH8YpL
SSHnFl6p6Xjqh1uIK/37NlC7wPH8Ox3ufdW6kMyf3yCrv+6yFiNZM1IMGFbE/ACB
KryEbzcO/GENe/ovnxun6QQzEMDvkFlqHcBirk3XwhsidczY70VHG/flMepbfRGJ
3KTVVjDWnsiu4n409U4GPYMx92tn0GzjEJzM+8YCPk23m/nN/BGcU7pV6jN0ik3T
CVGc5TkX+Y4pRYpS+Oh/NvnweOf9vPV4XB2lpf+BZeGML5QVRSvS9eUtK6sMmpuI
EW/JOoOnAZuApwniGtsfWVZdHQpXURZZafjq83vKP2NL4yxuiYW8CEk4aEhDp/Ry
afrsTrx38a//aDKeXHAdSfHCD6sYsgJI3qbFSxLBDLJiGhQXfOfxAhOGvxbBYoYD
cHBwHYQ8b8K6p2EGDRVCUdXGPTs/ziE5dJvB0s7oqql+n8NRJzbnMQJWmnh5lzKq
hSsTWDUyf7fvsr1fUFNIDCYb8LYPrPtZyFE0kCTEvhpOEaKCunuLmWzbl+LAauYP
41RMq2UwMtXb4T6xS7jP53mS1qEBsaivSgBMLaCr5+oKhxVOVPxQloxhLYu6dkNX
IZ17v/6tC1HqmU/b69UXxHvEFp7L1K181YlZEYQtKZ2juJUV8rJx3P7E21RfR/X9
62JinLNxti5LhZqqZDxmN4WsSjIJVK1SAx06DbCaG7eiJdYjfsgPDYqv5tkW+USF
/RCuYMAzVGwPuyP0luuDMSYzPO8n5b4pEwoT5M0FPYGlLm5Zpp0wbU+3bZCeH+nJ
CsPoTJGHsmUpZy+CPy6npLGBmZfAlmLZ6bLKZaIbLmDeyPGULOFRBSVXFKRz9L+j
5iJ+7FiDI2g46fyVwAHxOueyw6sVcMwRH3QDHuB6OonLEvRuLtlGR0ikVwxQgrXk
rGdPYRyPU9LBDjefOG3QLygQPz4aFn6k9CuhkoLc0HdWvpYWsO3mmlITmRjLmgmH
dFmpTarYK7wIRyrOybYsSw1txjXm8yeRjHkweJcZ2RbCkn2nE+z2K09Qu6lt7dZG
00a6zyKjBKB08KXN5vrbtUkcili/xpJhP1yXCd7HPaMI0DQIZmxojDTUh0wKyFCY
wMg1l9tgkb7kgjSvXrVWpOOY/1LLpLxieCM3YRsH2KsesXsUBYy0727aX8Y4vGY4
YqB8Xi0CyO0Qk/EXqWRD4BreThK1+oXjXkniWWGWvW6ly8dSau1lsu4KR36C29Dc
iA/e6a/U7fGFMJ2DDdzoDjJrfaBA5+dPUQTAc31gT/WCMJvLWd2H3nSCeROjbxQH
qSlp41i0D7E75EBlZKqAHay92cjFmVZYc+aRJOZSHd7bZrggnQU1gFnG9l31x9PZ
ZpNcscNSZe1OFnAH6EHWGj3hW6b67YXsTEqgSRn/bx0FKgqxKM29qsKd6q3ErE0/
WBgp1D/tERFaCY2PsgNx8A7CAahGsFoLqK2YK71h6imUeL3mA6bV87Sd2KUFswpP
D1v2c2pIbQcI5tzT9uwekRgW/FXC8PsNQFIKv7Q73QJZtVBRxATnXACxU27mAkmT
4keiqDzz9b+01NR4dCO69IeIgs4zp3N3GacOtSh2Rv/v4s5H8P9xIVEaiZMHcgcx
jUEOciwabA+F19RTIj4ihHgjI6ToO6aWBuHDcw+CnqEPm8Eg0eVJM0expJn41e2r
luVUnLViAWy4Ps8u8Q3hrw/vCmuQCk6JLvd9+CXTnBOLyMXEisknblBfgHcBWRhH
5bgbv+UOeXS5iMapqAdpnYcvlxE54mN4Tfk+OSJGEHa8SfGaRvhQU2PJqumNCYPO
7yeAPOOVh5uAR6jr1pnDj4jKKUi7GD91mGwME3hVUcvOTDyFoyDfgKz+CcRSoBL7
Q7Ho/pCwaZFAzVSNq3BRd5PW7wAf0jVKBqsffv/yaC0qrQz5NTWFRXjRNlJy0Ehx
Z67zTD+lQ4ycz1ZOLxhV/REMs4uhwJYl880q/dCLNFAXN5LFDLRoi8S79ko9wv8C
HBXxmpaTUvqs4TbjUN3+dihCDEMo8ZEIvwpfUNNYTAGMGojOqtcvL35mf8Vq0b+A
HT+4BFJ5IES3jZECZui49VHU7GLfXoFHTWMw5EK5rHTDSoTgwUNt6GIn4iwYQd88
gAeOcsaTvv29yXAo5+U6VxaxKopmtsMAdd3kJ2jsj03RGzReVMmXqWbNV58cdJgP
iVsLNy7/5XG5PvJvBRqrgy+CZfZ7f1TxGLbWuxEZQwcGYB63sijRALAmOrDWWXGi
tkw/HAhldxOEAmhsWKKBuFbZPXYQK7St2E2I20FI7LITI8shkCPLUcOaVzkqIHcM
kvJ2SeaAdCMl98+kyiZQ1qDa4gfoa2/fWUcJKMw+fGkMTJ9tVpHRuDs9qcMMeoGB
/UDF0r3kcUUAYZoajsbTJWRf4TwgUJjWH7qPk9JWJ9395GrTmW17x366VURzmRjD
Y0eRyosx78v163j4oHsgRqDGzbqNN3hLqvCjl1LpkSWO8m0v14wI4+UMcbljz3L3
E/P0BSoRJ8y9/ApQwsdk2ZP384oU0PyBKfWPdvjpEtYNhfjYulG9GYTWTItL5cKq
pua7npfcst8colVWv1L5hLnm8S5DwyTIP9jmygNHhkIQ45+MS8WoePVKo9JrSU19
Pu94tOP0k1LhZZKzOKFYIXVRJ4BkXDbBZmqo2ugkkQENd/5/zfdMZ7fRFwWiFMuA
l9UDcnX1vAdmM4EWTTY78QRZ1IDJyCtmTMyRtW/qbQlORMYuLusnQhUVaRtdLc+O
AwkzsJGpan21UIsx4omadij818/Ex+fhEqAgZ92SQQdV5MBUINmPrtyeiD3XtZ8g
qTZQvPUZ749Z66cG8hPzAGs9+jNlXoj+59kyu9McXNsvrtEUf01Tg27/IHyn65EZ
QpCVQinqhLa3taNF6P/fgL7s6ItEoKVi3JFxNWym28MbVDtDbl4IFKIJ42gQ7we5
Cz9s1rp6dk8+x9AjEmW9lhBaNzPiafTZV89oyX1SVedy80hAVus+WAewrrjNuUBy
KN9YJMNOxbIaKF0nnLQJrjfRfjFSvYQiRpFpz1WSlSP1GUVhW1+DywcJJk5C1K2U
1/iPbR7hyv0CyGKftZxu0h82a3fJBDxdXzFPKHfmAHyOZzXLaBgJUwPASsIqN1Lw
1C/lAITm0e4eaOA2ehKDHm52AS+gtTfXQc4QOj3k0DiQ4buiLt2tmLdIJy6sIxgJ
TQnQM/FWNpowCo6uy8NFXPJVDZBq2NOrdYJBW0badyl+YER3EMl58bLwAeEhWKXB
9TBpHwGyQcWc1uXUyWu5Dxy9uhP3I/xVUm+FRYf9i/e+AeYNZ8Gv6uTAAkTM6WFY
7s9TerdRm2Qbb7LLQEZK3eMDH+LHdtWp7FEqmjo9V59JBXjGa9dObpjr5xRU8t1g
fEbe5YtPleHKZUokhaGlG/EPD8lTHkdpFBCyqZGeaFY4xLRwyW+QsQ/88GAoRLPM
JyX7gVyPwYZIVVhOrRFGAvH43C+uaser6JNYChzEwhJEutKEXiGIhjYExD2lJvG8
8AQELVb0jgp8cRrcwY2HRMXw4dFvpqn8FLsi5DM4lfYL5/K1YNBVCksAvqFuj4Ay
fKYQb3PJ+J4rCC69tI4YWlOIsk1zL9Yno4cObhldlvc9c5jsgg5b4sV8eS/K9M65
NSCM/V2SkvZPveUIP1pFPxQ95wES715SKDVcVUQ8LptNiuM/dL5EaPav/URZnXxP
WIu09DcJQSe3hordLtVHeHh1MFGBi05y8XjRq3y4onuLQwc1XUkis2aoFIH8cS3q
13uQji8EdJ5QCYnnnwpHJ+IvqUGI9KXtNxXVyerJNwibmzUVDRx6gvCDmwy3U0FI
zXeshMShYDCxvpMeeBNT9NhVi4kcbEmavR7e+fd77ipChgcK5ZN5xpxMH1xpNgfp
wQgF+Vr1YNeaYzlIsJNd9O3GincTIMSKCTrfASVpSu03f0Sc7iZWmVX271bPb9oE
bvZ5n5HIdbJnS3V9d1PY/TK7Q5pqTnrw+LsMTCIC91RMKFQfBYv4D1BwqILFszSW
SZgf37BcYeIoifFGjWTZ5cTiFs6w+35fAEmQwlvKml1tY+V8v+Y7RJLKmgNVHsSP
0/YnyCpabPzsoBPB1srB8Sp+1dHWt5PvN9WzP816EZkGdMJnPeADRyF5m6AUPr5/
Z5k/56g5o8ROQHY1/A/sfEObdRbeUPv/ZMruK+hyyO8DkbNQ8PlCPnnyggugiXMI
r1F8DrN/D/Du6a/FwR1hHDEVwbKZMl0EaPLndO3SFtpYvIJTDBJRWhDFnJXTzb1k
jhupv55gK6d8gQNtlayHHaedzlPUHNlUM/I7dQ3Q2NBwHnvWzwhxvS5LCRMxlYyg
8vrjGtuttyGqk7QYV3ZZj2YQMQUwMPvlEfvg2SqsfS2c3jkhOlcFLHKOKIGCQrlT
tnzZuz7Gn5HvvO99l/n1GcwpKzmW8ir5XXuitEbKcSJOM0XepzGZ4iN7VWuXEFj2
0g0GR3d3oBFzdUfGIAwnqO76b56/n1kCSjPimgP+sEAN8kcjmJ1zCM3A+bfBNzJ8
wM/+/R9cyerKBbQiPMTCOFC1zrKU1UhzWf1WJximKO7aMBFGwEG1yiNVfGxhI0jJ
FQr6tOTocgLYFhusTKCEuiyphKGxY3fSEp9X6WKf0M87XHNsjSTj00fcVKVpQuk6
5rPBpgtK3K7rdtGTn1xuvxaGBKAWXslfnRBGOVEaZqNEn1qag32yRSKY99kAVUdy
z2pt1Pi83s/kBqPTVm9NfID4UcCW4hQ4yWCIxTclxO1e0RIyO+iR7F7Of4QXME5G
JapiU/L2IqX/fwhp1RNobZy2/eccXC9yOzCorh73z+K4v43fPpkj9pdSgV81eHWC
CbEtkDNg89E1sEIvEARtYgNMUMDpAFnkmBn9MZVRDZ6vGm1tHc2mFd0l2L7fLch6
E8NvhFQTC0QSEnmFhMS9j2I431peHuPRrzLxnH/VSLnQ+KVIr0uxcqgvnDAezT2o
JxetTXsLUH7mFQckT/1CtpmJKdnWV8tZpmhkrlsD5Il/17S40ztUElQJpXV/ebIS
ngqwrtMu6pqQgXLLid3cIv2ySRkTeO5B7pX1aHxr7jLHQMWrjREFJ0a1DTE7vB/H
D5EcGUjE9sdjgRXscUxO4/9bFPuN0C7MdnevIytrnUEboqpZrpwIi9jAi86JcQMq
RAlJ1XQmT30iI0ioJGqk0BNjjOsrlJCr4HQTs9jEcbFxlvriC3SbbHZ2uiEU9u80
uqMVSTyQm2kiIlW444TDvNWMFKyG+6or8IFJQHYO5CkxH2xtNg1HCkc3G9QVvHpv
yyU+Zm+PheAF8Xzq1Fe2gC/EFuWj0nAqS/XHHGAE6O6P4HXO6jPhu1pdD+i42Ej9
cNW/AWxqYSt+MnvrQddBsjRjb74iAZZIvGUvQdw0Lx+4mM2Xd1w449EOCUJH7EAx
dwbPVo4WEIRDd8Qwsl7dE/CuVbHcsf6CanemtVpWQdWz4o7s0/JfgQcUZYHliRCR
d2ISH7UZNeOrZ9p/0/JHWN/sg8AeL1Q/w5CQqw/tNgJdoJUplFhtpBXg2LxtNVuB
t9nOLf1b8ypxBZ+6pZ808vqvw7Mupt3zFIPYGdLLpSSYLEjVNyqJOHHZS3ZmoPYc
ouLniQMebBQsjicrXS/74csp74c03JNYFnChX9fYj7u3wTuCRg1bqEJrMJCsnNOA
7unS8Vd2tzu7h6yKNwhMUNiz5yrELSPYHrVBcJGK/nv3/90R2CI6dm8+9zdW0n/8
QAq5poQxi2B881HmfQrHsI3IgeUMshLAvrZr9gH4yvDV6MSElKtcMdMGyzqU6MaO
BfZj1ymu4+Gz1Ix+milDw6q9gYAXmKOoQNRdXf6IbZIWb2Y3D6eKlELW73K4+Xsy
d853MVA4C1L+uEPuJrXO4GtIcptix8Mq1yKa1QHxlkFoZw4jydaqkPW3N6+cCSJk
t3ZzNJf46H1gp/5PNHyak1EhpegjPmR0BKA5m6sibIxkc1TdHxXCz/EYbj+TfhdB
Y8Z+Emo85FewUiJmU7SlMrY0qcY/kn7KcFxGMTVZXGMoJdEhY6NJz75cU20DmsWF
VRBSjEoGdx0TiPsG3lT2f7TPAkHvXBYzuS7U14x1wYyInkt34g1XDxYPsHHsry1h
jRpijrIMVbGOSwG9sx6Gmq1D7y/M1YakrkIJwMEVqCOq+Bacz1HYWuVwTIl+EvsG
lozXi9+ENuo32jkmM7xtpr2HGm14XJ6nRPiB16TSnyn7eOa9vsfykymVBJpEqhsk
h+KcArQ0Ot0wkNglsn0eKQ2T2+ryA9pySAlJWGVEmh9xwQM41Rz4u33cE0gbmSH+
J91rUgm3bRicxfSUQzEmDg==
`protect END_PROTECTED
