`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hrXuMusR3mmco8134amgOdhFs+/8gixSP2OscQivHaj5KkR7FtjGVubBGcHriPB1
09rkuGoPrx6wAnHVi7ZyQi4mflKqygCluIwsxUMe3LZpj2WxkMAL3lRMD54az87t
T+z/maVDRPLdKm+f295qLfadyRXtOvtRQhRa3Fy1aSp0tou+1NFfFR7TDDSlhtwD
NWOzaDCH9KF0Fe+C8h3hZ1XUcxhUNr4ZjTGFg4MR5xsajacfbMxZAOz2OqUY/OtF
dG+Ss5uWq2F0EK2hxz/77qWatx9CndrmiSbuU4LTZV6f1Sg2LDCX/cfB4Pf8JA6w
Fllo/dZBjjeUy5yqMWURqTjc7uiwt2rVqOFWoed7nojJZ4YKRicPM2l6kfKbAYQo
gc+95fO6eJtzTNMnd1Yz5i0nhoSWmqhO12haGBJl/PkiUe2xSDKlWKK3PUQROhwd
4v2G/YYvA4WK4cg+/dtCed/AyrGlYGrwScXt0ppHN6T07v2barhGKblhAuMWM/2e
R6bEmmIvFk0saBF+OPJQtNHOx4rsX++BgozRMxznPmN13lftwrVViLbsVY+4PtKT
3vbM30Hlw6WZvRtBT2kLpiP2nivKB3lzmXtsqHWmoryX9+HRky1Z7G419KkBerOc
yWrShCtwIDvC+FesRJ+kEoZJGR1qEdzgBo4GoNmSeC2DgNKjSrVLfGIgS1Hf0mIx
C2bNDZay3Mus9zaGCaoU4NSyPCtOlDaSrlHq9Ga9M2hReu92jxCCpFJ2YuOGBejc
aLboGol+1iIbEGQVktg+rezkXj6vDU2Mo0tTRNcNx8Yv3FXt90wmvwidSy8mySwC
lAVHjQo3rhvAWNFIpzINDdBfxHdMOk6Iglm8BaUKlcbmqnBbRzqKzv3MPotsYrdn
czelDO6ykjS8xlpOkS6j8PEOxYIB0orELPlE5fxv4HoDWzZd56diI2V6c2kapXNK
+Q/JaH/5Opsh8/AWO0tzjsRcdSS9bXqEHD51HM3jH7KT7SLEC94kVOtdXQ1GZ7so
nQvlpj5Js8tmQPG+WDMzc4LeZZTPUrCjDGy3vZgtFiD+cnPr/z+n/SnS8hh5cGU7
JX0bmHBjVCj9IPl9W/gccpeGQ9DA5XMKeghj7TDp7F0GmI5T102XcEaP5UR5e5zn
zjWbDADF0tzrzT986MaHliGnhEUC6Abq6WL6ntu57QjsN7DS1/3gx5i2oonOic+2
TtGHyWe2YrB2nUKCquC7Mtz15Pv/0fdKWYz7MeiuY8f75dIv9ofxdslrdYMPnnLQ
kKot91fb0I8jSJ9QMqx060lrGPuyn4M59MKkwdZAW9gtLCvGae68vQX26P9JW6h9
2FjdBQd6SAHfBjffAN4JRQ==
`protect END_PROTECTED
