`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cwkmWx+F0DUwv2irwZ0BnJj05KzaxFTmaGbiPehJoNMcF0A/v7/CpQ/Bh9RkWdPZ
Yq1ROnn0KViiWDCA2bB8NSubjUafDSfZ/EzexJvMdwucO39sjJdHo7hnIERkT+Qe
7VHOtvZpLOOq2pzYvCAPQ14cjGaQYdK2vVDt5JBi0S5F3n/w90D2yUWiRPQXmuRQ
NDxvmoZ04mXUriQuWpbXE6+KMxIOtOxzdmV4S6MKyMcdYBE0g99674aZfD/HSL5M
jwx9b/b2NkowQJIafUiML4qiyUZ1guCf3HngDmpePV7puQTXMWeV547nSHiuZ2OO
hueH2/Ujx5ighzWVNsWhI07yYKiYkrO+paf+h6s6ELmX9y+QLUX6sBqkk1AwR1m8
kiLROGpGhC3Z+CMtj7TPKmBb9NZD+3jCipGvaTj0tFnHdOz6uNMvbHITcV6/4aAu
qx2YXWSP8qp/AyDFsyaE964qVKf21hC31vSyThEU7jWNtVhDgjgJC59PKAlZKwPf
iTPwT8bdGJb8VK7dJFLmHMrLlSYcBagVsCiNdld26rF4U/pcNP15rHUeoGSbol25
HGGAH30sWNvLvE7dpsODO66GwX6MCd+yHXWe5+B8KpUvbhGAHH39+RumNe+fmagK
A7jDY7+j9aXLJ6rsfZhz4yGjzIUfJRqZBptSIM+/fz1xx9yo0g2ru3Kf177T+FDZ
AjrHq7GJYuzFPulV2Mlu8KjtSR/fRD6J3pgDndlVWKUdvjrWkrqu+BhMpnrkP0Gr
+jBmXXJe/ifQe7UWpQ458O/i1KV0p977lHxeTYWiXZl3qpCKsuXfEjclyoqKSF6l
vTfSRAMyMRmuTxLjt+Ukt297nCtJ+krnPS1UEcF+j9iDsvj9pP/EpTLt1afLNrcW
rW5maV+jFs5/1cjEiHAg4IPuzfGsqvNCi3Uz7ILuuNc+IlXtG7VVUkEOOcF2OlAW
/xljPuTqfLxub/yNDKV4mceMxiZbf1BtLKLZVYFxJ5ia9LttQ+HM8jxyQF0ULf8Y
xCHOGD8vJNPt4Wpz9wsW8O3fXDl8r8TuC0w411hlZPehmoK3XUiFo5Peuwg3c829
NHHU03L4OozsPCl+aIKaopDrNMtHRXU+UCfxqQQCzGN4d40SNSbWBMAIH8FVZJlk
XwDFgtCmVB24YoeCHMq5UaFmZ1jMtBmSOVnIpZ/+xELX6r0xtcx8jjp+3MD9sMbe
0QoEh5BNfHeIF/NY8RkXlVC+jNZ2LqUKbCiacILH+w0Yty/oavQ5bkndTfuLPvyb
Q7ty5/96U9AgVwVKi2pF5VMYiWplDYqV+Jtai2fOCrV7lYwsl4yeTzfDe+XLyUOr
vdl02sU6L2F8tRS61iVb0e+97RtvXdys7PQEGcAw3tbL4gyr10f8mTWZBcoITQc2
91rplpNeCJmx4MWc7xHcK+ll1J4xACIKNsBB5z6SHT+hvVbLn1Zj6e3nwDiExq/2
JWP856rDdYbDN2EbNzI2OG3mrzn11n84UyyLU74IJxmG22elefZVSiNXCh6WGnUZ
GUAnvk519LJEvYcnmEhJVRHAybFNgRzecrNezin5kKpQt8aXUs6GxJAGNKiAsyg3
6r/OhsI6CND0Y20g/7skSoDjcVw1Czz0/66whEUdTDapksbTDxCOAqKcSp85iwHh
6HC4f68qiA/8+jVXB9BAIwmxT2trpf3MWL8H+tXRJt89/pBRAbP9K5dL31JCv2KM
Dr3WmqFRX+A9DXgaS06Y4vXoR8V2GG5iG42W5Z6JwoELndN+KALO6RKMdt3C5YKz
utncLQwQqAtdpzkm5+R2pWxzjseFAfLGPM31B3JkCBW7BCnOh/1ZmlWDXQZ8xHac
vOxVY//GzGNE9XR43C90VKZ3tgtKZjJfL4g+m5hozfozMAonY5dOCm56zAq7C61T
tQLfgZpf6sYlKZpM054jhYcSyh/6XYHXUz3OAVK6mouOW06+pk9RryQWCdkC9q8J
QvGTUazh+APlG7gQ5SKS8ZNU9J7baujLiM4BdF7Jg+WW4q573pP3XCcg94PBITVh
xktFbAB24O98jvAWe5D1L3xA+wjHQMaBYoFdXY2Z9q0lMPdsDnvRVln3XzW/2n24
M7bj/chAlTxiUKsb6ebrWVcz7hadC08ww68Tpz6d0bTwxk7Wmcd9erzcDRKNWuSR
J6wKUZmvUUhlCh+agCZAi1gSQmbutuGT3GFlKHKsVC0nAr8Rpv8p9K+Xf/rwOHXN
tJ6JwIG2BzQLk1leOWwswR1OxZ9AY+OnMym7PjT98A+eVhc0smBYTXNSHNwC6lTZ
Qq04wVCJ66VPpwl+H4OOdzym0xPGNkszKvnRv1DBj2ev65rf1jlSeeZ1cu3WWgcE
Rw5sDn9N4u4BUK85AsXkDCm93R5s/ilPqhWAZ+UJAFRPV9m3Uqfvq9B0jXexX+qn
XDq7KgttA/WBMog8CsquxPgMs/9f5zHa7TH3FxaQU/v6skBy9g1S3sKSvybuvzY5
EylRPVhwU+ZW0BRA1iM9zjsUTBNsML7iMsExjwmTGjTQBrY9WPLjZ4yvN1MhmJ0Y
Co395BgXWrkJ0ZCJhi5zfX0QBX1WCZov2toEyIlxPqZDODU2UZ1xNMx0tlqIbDgY
QMREXpF93A5qDGuUPxkbQ4W03gjpu9FQ6WxfCVa55iAlVpyQ77qI78RrWSpOTULH
q9MbPF9wNTHtRX1dl5Le1Go1URx9rUjbxwrqasQOTevS1asHSVwTj5PQlh8GoVv1
zgP2nlWLOmABGzOp7PgsIpW1l1oARCkl1rSGp/+8y6nKZSO4h7tIwbkm1BZvhQme
/wv1FdOfoCSPFqwB1EN72IsLCRAhrs1ID9TTjsT++xma2D0BWbj51uRej4AzVwhA
mhgiI0STJ1zPLDqjXxrvL7xPQZ3Etss82A7svOTirRwtv9HMlV2kNF+sfWjvHoe1
DTZkeeYxEBbqxR3lswd4QUg8ndT4/LMX0DLb03MMArrkWSmSH7aFNDo7d4cnmnpv
YnkM9YxGHLCGwprr/oHE/FpdmFStkXTqdZ7akcSIZsVcNJTxMwR9XL3NJt5oFf9T
lv6R0RlM3BVOrpFbx0dgdo0pb06zlvFmebs3dqbxOSjvN+w7KGCNp7Ssnq1FZAig
uRL6Tn66or3dsw725KbLAmbQ3QhNR0KM/FM9b0vENDrA6V96p7QtT2Wu2pnCPmtr
RA64ktCDe3IVoMcSTynyAw==
`protect END_PROTECTED
