`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AgOpEZ2cD2arlXsrCVV0Ei3gN8r+zY1imZWFbhwQNh8TO5Hl/b43Wk6txCButu+6
QKS6U8Lv8aIGlbkIu3MMH1ZHhntE/kv/KTGfFUn5/dQj5lGkxZpn/Wtn7iGaR+FM
4aBrPm2OrfqGNgaArm1B+S/vyFAPRRphj7+IVIFM6Di15vw+SqFMtUxiKHQaLrYV
LIV5IIk36EvnJcJGso0TX84O8yPDPXpd4aL5JtX8t4D+fp+FZ8r29AptnfC1OO6i
WNxyysCAB5bnSSz0yxvfSd+8T4xZe8hhFN4uEkDxFt/adxp91rCim+9YF3QezuZQ
BlspWTUjZmP+Ztx/8izHrQOUO6LCgG5ZBo4dypmkNBxBKH+C5dce+hEbJcNeJyvW
gFdtu2EcMxVO849aM/G15wP9iiUXo6m6ebjvoF1R1iW3bQqFJfKXw+UjNE50Kp9+
PSDVzab932LWCnupzuruyosLSJlClSQO1JFBH0XJRsPDT48dHJErJd5W3k6OVg56
xEdL+A+6YUyiawoig6kyzxmZYBndOxyRDkqOYNZReDSfgI4BuasQSLKPFdmpzTDR
KN4xb7x0sCEUWBV9+oYZUox/ed7MsI1j/WXWU4OHHYUlCmQZAk/dLu7h5Prv4Fq/
xIU+Q7ug7U8dD3KOqOv8ok0XwpfOx6i2djazXNkpb2cF0gMMEfpT23uVV9AktIsq
bW4B2pa9HJhiy1YpXmro6DIs69dcIHhymjPNcvVObvwX8uQXvEJuK9ATnjpdtlft
qAemDLO3+F8fLp5P51eOfpzPzxy49lgiPvcAf8+uw9UNu4dkwYQHrBBaL3d+tPYo
hqD58KhMYHwdfXH2A9KpoNYUCXjWK4pRU/fKsJt8xuEZgPrjGAI5Vw1A0I6NZLc2
L5l3H56MPiufEn2zaWR7o5eA2+N2UDvgjRZ9kp1rm1k=
`protect END_PROTECTED
