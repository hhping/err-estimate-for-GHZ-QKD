`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oVwVLsLlWMQTTp8aGggo6WELuQwezSOaFAaPf65eZZ8Y6TBE9RprIVvZ61sPj2x/
zR48WVbQkSgeYgJD3qYzUOGCkvxvCPReJ3Kt0tAkRKgElwmBnJSuHfEgvJgCBo19
Dk4qQCXCISWXBUr8PkzjWnRyFEqbjPUSw+POi11EtijOnvaVgb19Jwv7c4UcYPZm
DRxWfttt9PPgczWFLm+Y58uuHKImQ/zl6liHcJkQh5lbtRdgtTyZrq+vL3DgpJ2I
uwo71QtkqtDASDXCfCrHCvHey7n5z+q98/G3B0CC2adF3SR/Udzpzz1WjsfpoPbk
6BgPdf7Sen4FWx9kpT/ckuCWP2sccFgB+VPZD+VHInH2a4nZdCafkuxia+sAOWSl
w5XIb8dpEDHSzjIqIDM60gkQRInD2J1LLK2/SXijRYhC/JpX83XSf5eKLKnn3UlG
EGcw6panG3d+0ICjFNE8774LtitWpoeqTD/TkKY1/iQzLfpar7VKESHddoESsU2n
hIHZ2VhdTR8KMmGkwU6jeNtjj420qgRiG1dWrNUwRRp+AodgEyYa5QpNvOIpwGMA
NSs5oHB9OLcFibepEFWdf7HNyNUEcbGX16hkrT6AuMkIiRjxhNiGiTpl+JW/jTto
FMFE8JS9oudA0JFxbHE+oPY2YhPJvycxD1m6PF+zsviU6yor1GW2Z3hX6gHreEWn
vm0Jln9RUhvHoM1RS3lT80SFbS0QdGQymwwURwIXrNE3/bJwc/cHea0vV1rzuon1
2+0qboUhdliv2JVHT1PELQkyR9052QJuOsoPc1UahsN6CwKlUvJME7oWPi3RWBoq
+8FPegiYAgNkns80ODEVdhMrN+WrVjufcSMZV7ppTq0kQElRedhx+zko4KP32UxY
XPj3WtwiYfLumrylcYFfV+xWGah/95FBaSLH35uNjxnIfeuQ8eWfR8uSntJEDzbd
KCw8lGuuH2YN93mbRqcOGVepi5Kqurzbx3cr5f64ujWD7QDPnevrIZUvHRoEW4hI
6p5xuNfBo3zo4pkmfqX5OhCwZ5noiqPJFHznGCf3EriPRJ0AJbq0hlUclPQCijB0
nRoBrQq2YqBzilUcrPvslPR57056BEaTXKalR3wgI3ffxSokw/k8A2QsiV7CBF6L
b2Lp96ZUkbWTM8djKlBFsnnGwxG6NoIPMkaNGOoEs+kEPzVsUEKWVkpxie6hRcxs
KXcG5oEa/xOdWx7pS5qM4BOs80JzjZFou194nHLMHL/rYrpVQx/XR0gypFOCtpii
yzT5JRbg6BWQIX4Yl2+JaP0fVA+hTSFoJ1Uuru6akMK89m3hxq06s+s1UuV0wJp2
a2Jt0osNTQATwv51EAiPxRU3rS7eZoagLY8qDfOPC0WLvrnO8APL1fyYBLfJBN6C
dte3QDLHFzhUQIYyomaTs3T9v17YqkRt0UTtj2VZRUyTkt4CY+CP752/DIQP911x
SyfiBS9DtNcrOHgA5CVVyhTVPY+SuHjBNUpdsSrQ/k84/5g/Yudij4Kh7EBnO1JK
KGCJnrRBB/tBp0qcWbsCA4qVf+B8wjoeZzMxC7Dfl7msNeE9UiWE3iMPIXt+U+nM
2UBSENH21FbGSESFL4brRAlqE6haavD4TKE6LimKCPZqbA/T0aiYPSvp3NXibaeN
s06tpwNvuN3klRgwdK25ndyf9kN87DTl7sxytP8A6cTrCsvmjx38SsnaBuwWO2Pp
/XQIABeJFs5nMwQ5zam916p4Jak0xfzVAeTwWUfxzRTQKizJY/YQXZSN2RYpG/Vh
r/s+mbuGriJSXwA2LAeZ70KLFK8SgXZXWvXyOZYTvmVTBEK5QQr/m5ESk1SZReC0
OHzrfHk4SAPgld1Ic88ye3M4RT9CcqQqEPh3fHXFXiB9jaXnCZytufzGc1tD5h41
774DB2SpttbtlQwxvYnwfJwAfg6+C8v+UAwwQtuQIwDhcGJTagiEAaX15mJF4rKf
eOu5QFVoRBe1RhTIhLLNCI+mMWTwsGLbnpHnrr7dmKcOdmutz8wul/BqizSkIcQg
N79Mynl35LEdFzkbD/bG+sWkBzd4ujawJl+CdKAZxbDIhNgeK3butgKmJL7MyRGK
xsrH4I0w1NgjNGv7HZaWVaCSzKCF06V4guPG6XUTcfWElPZKK+jvDV/7OHBH1h2M
yMkJo8AdJw7DveEyXEr5LRaBZt7TRFVr140UgZ+1Lglegoc5jWnwCDXyI1sqCqeI
mJHyYtsWeE1nOScsz8GbUmKyttPNpuDy3oOppdCd5YElzUtmBnrWi6zMcMAoLo/M
18zO5lRQ4aYYz32QUe7tzSZ2crHq8317b2nFVnOc7WKEKO/5VjiHHQo5pcky+Ti9
ivPwF6etVqoA+bTvDF9BGEBYitM9ZU2+mLJ54pKFo1kw0ei9A0Qf2FQtdqeag2F7
GlGiYS6aouSPVJ0WMFJ9mGIv3irYWxZW1nGTL7r+/6YlsHn/2NNAvXYITMjcjMsL
pjqhaKF0DrY3u+PKGzMzdHqbCX0ptiHnqYsH4KPk7d0WIKxmyOZm1MPMCD6PSz7W
B+l+DG0lPMq33TJW/WfF6Z3nJF/Do8ykP3tbGjmDQsYqjCVo0F8dYIbulfU7eZgk
MaGSlSG1E6ck9d8uYAYBLxPqqZO/VP24XNWuAULujetXzlBYOTcu1Lp32+PZa5Nw
XJbNvyjC4/rKaffCnaxkFQ5bJ0hGAMGlZS2RQifg/URWI5HhBFEtHiO3Vleb4sB1
WE7dXg4TAcFaQ+F3+R0bCJgOYoEPh4Q9S78I8O3DGBS7uqilKrpMbNeG3q2LLMOm
8d27pPF0vj6xMBJHHHqCkFbPsGS2iDxchevhc17ID7GayeG3nUWL1c7ZY9GobbqB
lfLVjcWf1YU+ivzyx3H8k2uCXF9UpkSdT7dAA09TPs7hIQ7HUUcKr4WhdyEg62n1
vXc3ZQlLxvrNlf2u+/iOklioCxBzZKY4JJnm4CRrH/rAV4gnYchoVseihFRsnas4
X2JODKhLtDqf85sdk/eZlU9LtbbyEIzVW+gX7SN0BNAJ1y7yaovzyr8LMGOSaCrh
HsKX+XGpZgL+SOm7yDTBIkUDwqx5xklEMPFMRyZwDAUSVyZ+OLmuAbQorgghI2bC
2leD29ni4eQlJEghH+btjUvIzHg2OCY6fkC5VCoQkizKvTYb7OLwTCOxoY7E3FvN
kk+XH9s61kA8zZwL9sDEWO/hasXTzLIRXzyyU/EzfH7uoahhCFGpVN/3jJ0LnHdR
rffj8vT2m6280xM3GxmTQoNLUAjTEC2qWf59SgOf0KTu4CArxOLS4bsRR82Y2edJ
c7cp1EJBRVMDeoXpbURa9GahSyfX3LDwAnNuf2F0kx6vgqOfCxF+c/06C9Iggj0T
BSIe0kpXdTuZgAblA5klPfj0cdT9GSGjhXuvF9Gs2GLuSCG68lFyLBinAH8uYYcx
GxTeAR3xAEScF2FvBMRPl1f8t7sw4stPLRFqp3ViDUXxLbPAA7DRRGkLy0lNa6Wz
nNRjlehakuWQQfnGrZRrjhC+xjysbEJxaNj+Ifj2ZWE+lqZbZrqG2wXj7j7Fy3pl
IUOTxE8nLEmaEJdfPsGnAfIOwV+cAua5BS5ElefZkmXRVzXi8pPUOlg7gJu6QVgL
cfw6SiwoA/sHRjP/XVX1tcJHd0DxhfmVru80+cY5rHnhJMqTULrfz/pe0Tzxkn9k
rmMqj358Iix1rqvReT0vzQtMZXLZmilA//TS/0jj9EKzsaOvW3N3WVnafJJCF/zP
72H1bEJYwhN7mIbA1cIKK3q8tnfBBPJUS3xJbtks/bbPwWG7mHonxOYnGF+bnieH
jpnomhyjcTn97LmxuMapuOQVWMiChjI69r/pzd73yyUgTM+M31Dg8qBu+H9BIhZl
Z31Omx1EPqFzM9sX/vf7PyKQcjyhknBK0UsPBhx5WrslxjwkDRC1DWMtKlxVfrLR
kmpMtUfnVb+6Eevo/YNGOjnyrr1PgPpm/w/fHOwiZKwiONipKHg1HBq7NcZqe/id
DfygpIpsottxOyIl8T1hT/FQcRwr+CCloVJex53x94irevVzQPhkmgbrayM038Gi
z+Cpdcl63mymS9X8vqYTD70WgcUty1W7rae/WwU93NQp6Aa2MbOfFjBR9rUHZiu2
bJQDckfRNAwLKn5hb+MUDz4dzWay0vWhRy344/g9GKJqpe68f4FJGFEtPrc1FVdm
Yn+P/lUQ4/IgLHqHHdKEYJBXjCCEd1Z2fZ/ypMh+JutlxxKROBDmjwFrOsJlmT2p
GBsXEAUksOjvSRoZvxWmUBgLSED21RZC2bTu5Ss8eCkCx4Pi/bceFOT/SpIa0J4o
jWSvWOF6zL4ijuvauoaOXVCaHXCfsOMxWa0+B+8N330NnBp4Us3rWiCSBf+IAllT
gb86jQoif3mFt/94lJHMbbR+IhEr8Bb1Yjc7ImzzZ9nfn+5rGbP3y/L+p8+Oer7k
mh+dD4p38xR6dNhpaJ/D7EMiGvTiaovgSw9EkAzPGjgbAX1Cnwmao0t2VG/MkxTh
Ry0es73YmMax/DXKFd8BonNFQKfMoSpx+yIKJP4ehdVsPj74rktdizzpj6KjJWMg
jenLqu/RIvA6jLxzL8H5mg/ex/+GGk1gAWXaPdDFDypVn6UHy2NIbEFf0TAqLRRq
Ziy3Pzjn8/jRalmYeGnKOEzNIetY71bfxu6btO+xgGUKGiNLuBlKzrQGiRf3orVw
1EN5Quv523wnqsjn65boH2U5VJPZgzuAGrM0IGxCVIcN0fKXYZn3r+SjK91qdh4+
gO/WYzyubC45j7z8roQFHAeARQ/41uq0E0R/HqJMMbGVh4U8hSezGbfUs4StMajx
2JkcJGHi9PgmFvVpJggFZbYNGXWGHjDfHjUOI+OQKi5EhiIsFiqOw4w3jEc/jat2
DNRaq5JL4vAFFiQ7CRcw5S6nigpE7UIZju2GFEOxLDHHLLFScVmOK+h4/Nb4vep/
8ZlfHwZtEAqA1drJRvGKjy0rznRudQsGft1HGAFYsWtl5VXZcFyJRFjxrtqc/SiU
FZzNW1IBkuRVWLms9AhImA9M2LLK2N44YaGS+x336iUOxMFoUisqDN6M0U2M2fsb
JTgjZlxTlhlhZVUZ01RhD9cgz+nmFJDXMblIgyi0PCu4z41Hsucu/jnwERL9euhf
gmBcAeMEmfzowUFFoAzccGZ1GfmGTfkbfiRUvu2jzao9Dgx4YWpEtWKSrIG2h9qF
E9ASOM6uOxfrFnsdqo9qmKFlfmjFZoOD3UlUazqPKjLCLCZtNC3cW78c/cx6N9Uo
NUmfHzKx1vUcmyMSdmZ1MMpVpHktyE4LoWyEURuV7H3SVsPpbW7wLMLOPkXH3bSN
n1X+I0bxDkusRORwp0wlzvcwzZmQRAa4K5SonhKoxMIrsIWtJnfPUnLuiaXq17K7
2S9exjOWXR7PIvc8WeTuf3PzXhfQB0+l60AxF5cnUN4FaQh15/8ZBBvvsCBnAi/W
GV6k8pGrtueW+2SYO2hkUBXn3xNkCDm/s63dZMojqz9KLzRV0YAhQpHpUgj36X86
LKbgFSYdf1wZhEpniJBfd/eOlVM2Hu+Ug9cpfDYnDH+OFJwyoFC5QDZpb0Jo55xT
zG4Ki2RdYRuHCJTbUUTe2S0sUt25Bi7t9om7dl/LCU6cQakngVSzlUYEAkl2xPMk
0yLZ623j1gyUXB5YNxe8vjDYDw8oX/50J5HFE7Mc1hY56/Xf1PVgElD3ERYwJ2XE
4q3u4UYFDTykXjqSR93YNjgfm2oSrON5Udnh7QIWbfReMHdgUCTpfoT801YbSeMt
bIA4bg9lGngfVNDlnREoB+r8VZr3yPiygcDKIW+J+BYRcSy484iuY0ZS9XK9zjJW
Q7LX254yV04HkBy6trh2+sSbu7MHmrt4BcjBNORlwyEzfQU7dKxkzHC4ZO8fV76N
uecXYrSeEu/D5pqyD3rT7eAE5EXtFzOODVtQ5tysARv6K3MC9civEsNh0pCsg/Vc
T1B2qO7ai64ODXT1Y85X19nBeJDC6OgTVK/oKaiJCZy7AOC3KdgnNQYJwMbnZQ/d
PFe6OapRxWqV2HRwGufJrq4XVNfQmXLW3xImWmMbgy+8//vujM5gErmn6sXluLRh
g43PMdP4hig6QbFyatacuwszlx3b2iBPo7xg8M/khGY7XjqfhUnakXhuLFRb8ph1
KrjbNwzW6X68CVk2pKaP7lGFHShSPJS/OuARtRMuzM83urgEbTao1XmNvEHY75li
bCr4zsi1L/Q5LleXudN1YPxlQsNvGcxyUTo3dyYrgUjl98XGKRKFJafxxr9UJrcR
oN2SKp/y+x3PA9HaH8OwoJMxSNRhRmutyrFFeRDUkce71V87UFzBR1LXYtL1/HHy
qUOYqnLQwihwWH04ifL/1xGyQlsdqX9rU3ijMiFZRhdgamusv3SCpGmF2RyOiDtd
W0zi10TwPgfNNyEsIE8ZsCLLtWA2SgObrgvqhL1gOSxxBXlz2yQ5cHagYryyeboD
pV2Mdz2UlU2Mqd1w37qSK14i8ob9uuP/NkkploWvgFs3OTO+lxdfAZoYohDRu/Zv
UdltXUdCcFlfqrbAXxgRULdHIzuHpJGK9wnvUJnrF/uXRhqAAs/a03o4TSsx26G6
6zYZeZJXEZ3LFuUrtXvP9CLYErBAEPfw0OyjvP4+P9ND8wL/t9I/BHDWfNMVzyMO
MYy4XQjUtZith8Ub7iP6x0UTKXh/Mtfgo0TJui4jf5TCnWH5Ieu6SJAnxBnUkgY2
e9Yb7yOf36wM+RP7f5pAPmIYC4oLyQNqK6pbSFJrmvuGUWqm5VCuoSICpPwe0id8
2cz4kfQmo/FKQzrJ8meEUp9zfH8AvOIY/9+zhpHGmBtUyPy823c+EE0BZ3jRYzmS
+55tTDcTEBA199m1AFWT5uBoNQp8g/tueb29UrXwbj+N22ORcY+Sw/q4yOki0uTW
RyMXF+dYE+ogP8K/T4Tqs7Fgwe3Z7HjFe4Cjks4dCg7epw2lOWbTW+bGQX23xDFC
FvVBSZVq7HMGOk7nkKAP+AFv0DF7caywXIfGHljxzx1V13HyYDUVjUx6PBzOgLyG
KRZ08R4RmbZjMzCRY+U/6T/e91M6j0KWty83BHa+Z2g4BZETkHeFBgRJAS7L3Q9Y
6epW+yxqGsjwuQq3pqEze1Y+8s/AQBoYhJ/tBKk0+Mos0ndSz1p0FBlREr4EfMQ/
YVUakPZBKpczN17o7IBeanCDZKtYAu5nsz0QqPhZsUNHThZwXI7KNVruzVG/Sk3a
5/iLcxAq5pIYhOsE5sBYosedsJjjALLAiA2fYsQb8ta7Hv7sBUtb6bJfev6Us6h4
cJLksG9ZixHz7ix5vR/Mq7OBQ/NYPofmpQ6FyhII8ljyAm+9va89P1QxtYoFh7Q+
NI+ZRQXK4bJWMhXPhylbW9HKaEGPuBFRkrcXXn3+omAgJ7oEyRt/FtEJZgBWR/oA
8RWAWI3+8RXluafFJWkeZ5NlOp9iTSw1XCmMBXsb4CsblqbTdm5fN8P7yZ2TXuMq
w8Z1mE3rZBhxko5e3vNoTfzJAa5SHZ4rF5K2bIpu5P/lFKjek0FyR1kPKvxoSo35
btUw5U2GpALZAOtjbBeZa66HGNBOOMNWe+vkT6eQmOixp3cnTvuM3u6+dMP050yb
HI+SGRIcGnkU1XDv6AMQu7RTJK1RnBSFAJg8wI3LDQpfbP02P06xxnh7ubSuVUwy
EDzPJ0cPj4JYPB/1JFeX6qieoxLyAwIjEg9Q9BYWGqXFHUJqWlTGYkcgfXWkJ2ba
B/HMuC2jSGdduu+Lwrgl5NQO1h7w7MMFHGezbZxXGK3kjrcCCY6LqIsYufTN4qAL
1N8BvBeJZRj9rokq13YB3xBXHurr3gNRm6MQB47IObqTmOdVJ8jnTQfMVbYdqybZ
atrXhjENSPipa3sUWTMjgvvD0U3E2s7Sx6C6aUXkvLbbw9ebCwbBFAtwjSaPWoRt
iOACPHa3O5KE1sNGIVHq8+LePvpqurxoeiE6UrJXkdx0QB223Zs7uaa5wT0HgSBG
HbVtKpBhaO/sck6dlfce9Y3G3AyUr5DSHEsLnkV64yIQ5sisPgX05R9q3B+R/9Oc
8KKhj0jKhuSUt4n2+G7cw0pgcfu+ndOb9FBGu7W4DD+V7jc5Tz9h0kU38rmZ0uPZ
yjqn239bmvUHueXCeQJExq+3od2JjWteg41wjMnL3obi+387lcq/RUyFmjivJjf9
qggvWjOW/R8liHIz4Sa+zNr1WxmK5FYKgI4oSOP0y1IKYX6hT79spddC+fOxkU+S
3Aysz1U2JS4/aov1p7BRLFIq7dtyaQ37Xo/JAEhm5uh8/03D4x7DYyKUdA9hEKBP
icq2SGhHKL1jHr3u5Kws5u2oRt5b/SEQCD1PiZn6b2XPtsHw7DN/qBPw/3TZWfHy
iU/m6cG9dp+WTHtX+AigFnc4fCOKKWc5mxByK1pnopROTx6EOX5XyerTxdDaIGmO
pva7v4AJcwQlYUoz139hn/VV0cYRi4Y6h4OIFdpXmDIhSnD3s0/F04Jd/JDedcPC
g6VYm1OEBJAseqsWMqKJS4GW9bLVT30jYA7Q+V0j3hV4j6BrMx5v8T5aNoXuFgD7
Q0XkOiU9j7GXVFDg4ojNQJoW8hmG3iKlU+G8w2n5npmJV2we+SrGQaW0rrtLl0AE
JBWxTFlh07BljNTEsU6Goy1DALUs+H8ntmfWJRhJnllVeY+P361IIAzKK/sV4CRW
Y8MV84qfQtG5buugSbC2N6yBsLuS+kFqnxJxNGj2HOsXokvIzbpaYoJFeIGChn3n
F5gxDJ7LwLqxiSSNPnHCHAuDilCWoI98XtwOaU8DQ8rQIjT8iL1qi+s2GYGq7s7P
siO8+noQWf7mxPzIPel3FUuZs+MPhOt0Uil/jFijZPwHXLpABg7MWVtWdsuX/6I8
z+pLQeQy4y96E4FRDsGXp5WIp++LU75pA6/LxplkHRsQWbYJjxoHR+ZsSvpwbYSn
UMzZ5on83/lhjt2EVGuquI8OMqNw7v8RP2MdD3hBwpk+f5xsT6GKxopuqFJCWlxN
dMqPTSkDp6oNQd/TQFx1F8tbPJViVEjuVlSe4xhb61+WkWEJR5sSfxbV5dFu+m3P
BcL/XsRQUKSbybKBq0z48EyVVbWv6KDnw31OtZytTh0MeDQbf2YOGO/Glvj0fdOV
SZXFDwIVOyBO5f0NoPAZGXoeKXZrnMFVxDjeX1wEz7qYRtQKKsrf14i8oZvBqZiW
iZ9UiiHw+Zs9lt9VAJJa5sSNn3fG3xBjXQgLe+oNgUvlTyVW4L4Oh+6bsdcXprUW
e1OlRjRsQIBK5S6fVxyKWdMBEHWSJHXH0642C0Z6XnCYbeHNHOQCHkSJz8qGA7Wi
Qe2ffm+GyT1KsVnFywvbVxa0E8oKPkIIc8x027hnc62qwBa67WFw9W9k9W6MDcLI
p7jSfavo2jfQAsERdYzXq5INZ2aUttTVrj9Grrrh6ffR7raJpqtp5GXlfewiCcZT
tqgxwaN4nmJmbDp6vSBHBw/cD2dKANz7HLluAiL8X8rXrTCdwAn/gWBq7tEhWoUy
sTTrRJWARd3WvD8x0wBK2zzCXKLXqcGeFzGOnnoKIXN0fAi59qLJAeApLO3CBewm
+pF7q1ZnmpLyIp9Y9DES/bs/zVBjyRXccrjJ4FR5UlPoWKmhovH0aiIlFHwnekwS
wVqNKvgSRyLnLID1Tc+JXaxJkDTgOMGY2c8RRwgy6+t1ywcjkUq8iA/GsoGRRYqD
FCrVQddR2KpDFoV1dQyCyIPKjY7MPkAdvt6IXy+U7T6Emr+fmGDSgAOReclguMoX
nt5Hv79GXu9ewQ8xpl8X/MgQTBbvku0erZ0c9Z0AWmWXxuHBzL349245G5znXlI7
C0234NwRxvWIT/Y8Ubk28oFVwJKmuuMiMuNisS/yDRAh0J0lO8mStoQWvzD+SuU8
L8CwkQxCT2hBVUGQHox6OGt3MCeuDSrv13AA8jLFFctnosN/67tWRjkqxj4xoT9F
bud6KO0qCcIn8o2mgXOUqlTwH56Z8iXS0E5FKXb/BeVxxq+3w9f055DutWo0DmGb
qGAgm+q/8r3Dv+wffyIO3s2bVv1+/k64SptSjNzTom+a0iJn4uxi+Ae7QWyrstiM
b48crXhJr1JH1giv3wv7meOBUbaEsSMVMJQ1A3+7DAxj8qjEl/SrploVpaCfq44X
xgp1qtaw2dTbd6Aq+q1aCYjti1HL7HDSTEyfPMZLZy1r6+LEb8h21K5isc4Zdcqx
1oyD99MdNbuTQ2SPDtijaCR9Zx7KNvBvvoCQgQHGH0dMvTDzgsO96Ex1pfOyfcpQ
cZqAbKevoxrD2mHrsTDq06hF4a9M+InA+aLo2ZdQ7bfxQ7qrx2sx9tHbqD4YUyIQ
3PgMNNnmQHQCcCjy8DaLOgIdux37pMpDM4X//Mv+ooGzO6r9Lf/S9ybw6XyCq9Bo
Td9nzCMtk8uHvutTaowjE0NWMpVlKPkkRk5g+0QcVGpBXOkVPuxMKpR1xbCU/mVH
knTsVvmRcKvz1Lao6x5n3Sevq2v06VcykyLWTe3Tv0ANj1PPNlC5vdzeCy8opJ9o
J1At6STudzyHZYFD9xSdbYhaGpUMWgXVZh5ravqHvJAdU4ChwrOE/DeWxRMnXv/C
dmrnYYXeQaDApevbKC4jv4ukZR1ha0Yvw05q+bxWOk7G6Lilql1pQ4E3HvIBM8Rn
PtYSjx54/ojp/dNodrBS5VDiEvArBbeKh9w9zipHC+TXisSHQQZHEzIjzgB77YA9
FLGBG81U1v0EUDzH8ynfCH/lEv9/kC/qX9UW5U2SLkruF2j1sxKNqLl89v49TiSd
ztQk5vhRgEyh8uB6dIhSKA7dKrpU5HyHyYpGuMVLyl23IBOFNduqW9xYvzDML066
/HZZEIL8VO7cDuYoP09ryHxwpjdoYkgpnI0lKvu2zL8T+fgWv5f5QOkhqO7BYZFZ
hLMZKoKDXksks0+RCYFGkfuJTQxcy8NlNj5+y9jhzCAvIoAQRUDZ2irUzVKbI4xI
EkTuC6wuwL5hmcxAuLrsLMX1Rzi/Oy6CApHNDwqIARL5RR6R3Z8A0QRxh7vnEx+W
S1G6feBNDYE+kYMEO3Pv78UtzeaDwBBIvZ4WjlYtWMytTIcMTjvAKv1EjucIAkCm
c9ZOdrwU83LhFRCJNeyF6Uy0/4moakkuaa7XNBFdckTqZbXADKuiMAFumKBF8mbK
YBcrHJnbUpKmpq+GmODZoOhM7HqhJjWS3U8PEskiTmNfUmLPF3P1SlSxQZVh5RRj
2hdFrZDPiR9OWYqJY4uRK2SWzK3Jo1sVrt9PqG3r/Rj7dO41cOI1O7V7p8lg192q
587q1jzc5FWA4ny2SjddgXq8SIJtKGP9h5QwH4c5Szs4JznYMggbER8Nq0IcoMM6
7sBJVp7eTqkiJMk3u3Gh61FbuHrHnLtc8a7OAvfxLMhsyjOgmXAQ0xs9hPFvxHUF
RSoMQ2q744z4C9qEUKr7NBQY9Kds1+iLqQ94jjqhlYf4HHx7sfzZiDNz119XVUqF
FjOq0OGGOL7j4rHqOEdSYdSrHVONr8mX/hph4KxKir1Jcdkw8ZeMqTTPyqhYi4LJ
M9pc7UhTDOWNHOjqZPjRJ9vLK9+VLhaBInBn2A/9BiYcseXG8J91fFj1Y4uk0AzC
haPrAAcyGH1ZcHU7Bx+0g6I8zcYhECY9ZGQiyXqLXo/58Jcr45UXx62+ZW2+6Tqb
bbbcHbA1hAlnyqwCsOJlaPjF/01pYZOVhincce/mY9IaWVTEuzx+epW9axZXouUt
BZnLWAucsuAHE3XPYVsWWhxjDk+1Il+7SdvPOTjHD6mc4qYvn5mrPxH8zJIn4p9S
PQMC0DMttwuRv4asDIQudGcdsVVAzyqa/IZpMId8mtFmf0bh6sboVfNGwC1zxV62
RYvRDSud+89RQKAHbM83pQcjuavJMBuhXE6qPmnX/w36hvxGZC9Phk5LqAVozZQI
MOTXOa2t6Y4c2DEY8LIykNQJrhqxoLv2O4nJKMRTXslgmgukv+4mNy6v1vEywEEJ
7vKc1e8rzi+FdAMHBA32VaC883pkoKu5eSRBve2g1ooh2qnqy8ZQ13HSa/3n1ciN
UQy5vkB1yxvCS05YJ7ESy0xw7TIVytFw9J0ozqd5Wb2FUg9w5I+HXHHf5BzOIUks
/PyBWMsllDEcsU5vfSQns+ilb3x2G8w13AcGchL0StjGpeNud9aABlBYuuYPlera
BH4FRWyimZnIu3gDNirQhRQ+MpOiYZ8jbQVKLrWcKgCpy1dDp9TStVn+ga4pv8rb
GuPhBM+l2sklEj6mw2iRt5tO3orvpo4wWKXt7K3HeNn/+8d3HKo6fH/CQEaK2HIG
ARSld9nMTYGEx1lHGqEn9JtzkQ0ZoLrEjw9t2L0Gk+21mUbwwNLEfkNOwALDgSd8
VukUROGIZqmMBDsUekMHN197GZRwcwNl4rHSJo690sGNiIWWzwZ3pdlWwG1748zN
wPlQx9GBzSvEMSkQe5VKlq+W9fCnC3hgPg4LIQLWN9pS5i0fSLcdvwUalURyABQZ
qiXghW5kU2j8ksrv2fT0h/neXrfyebsYh6roX2w/0BELCl7Iw/xfklXcgn/wRWjr
60vsd5K0TvEEn3t0SCKqjaFAco98uPaoW3XgA9UY+LlrWLf+3qEqaOIfyeEtlnuo
zIgbThTAix7iYbMLejp2+JVW0HS73z3XpXhwqJUsTeu0FtSnL1D1Q5nNNUZsqNny
BoFHqOc58qB5s31iTCcepKOz2lhyawSeWRvoOvCG6/wIW0CfT+FocpQpTJSX4u8l
uQQat+GKhCxmBeCD12e3DXun/I8jAiJmXSFcqlnoBpUZ2iaY+MsWPYAohJwqFAEf
/HJOp1UvyTlYIBGjkUtyz5KHgdQFMmWmGJO44jbMPi0h1lju6L+sEXIoqrh5Pr1J
NlL4LNct/3GpB6K43j2A+/jIFhSG8ozVXsmjKzqpLvtPH2e1MvkfpKyu+OFyQP/X
tNhOjn30JThgmbe6QNL3ihdDqcubRqT19PVh0XZPo6bFJsm/XZoGrFNbRupHjNGW
RxbTfScbZxPYA030oqKODQjY78ewOBSeFXBDFL3VDnrZwLCCW7a/2vARPT9CLYqd
KmjwTS275/T4WBL9YqMSoABIgvG6Kr+0ZIss4eFXJbWqbF1RQ+z8aEsLtty8N74e
a2Z/pKlzs/h7BtnuIgT/QCM40yXxGn3bxmQZ1iCtojtdQhAJZSFwTXKTFssz/SQw
Sfcgv9dfRX3vDj356Ti8zr51XFSmH0QJs55px5eRFTgslCtl3lCf/niJKqt+E2/O
KkRpMCVzwDdip3WEuLavZnh5+ntLzKYdIHKXC26STBCs+t9ATuH6Ww/YkxvVKn+Y
e6+c9q/7LvI/zeeYDonHYGEmAg40rz5sgvDfG98A6AJWq3EiKTObm81edP4yItNk
SxbzGNUyL8BbXPvr3XtWAOh8lSVa2hALFb/vl0po6+CbBmSLB+ubSn2hjaOZ0wja
Ar29XTaEN64ov6D/tJuw9756EM5o86oC+On450i+DkCYa1bPOoFMGMdmtX8XsnnX
PIie96N5bJzPTRVdT1Qb5WNXH6Kbg/IaHNp46zZMYUQ1rYxtrkKnadNH+N+eQg2+
c0rrLFPDLX4lDmZ6gU6Tnm9IBNPAmoFqBlMUZACC9tAEDx/u1OoUJ1lG7Z/TMdGc
uyXg17f2zYLep69UUi6vH9Gv+f1WTXjGYOomfA9qpfmyNhpygRdsc7XyxY3RsTGt
A0k4js6kJPhKueCqy4ZTCaH9hFyhgzgHZb1ltytdazaol2iZtzvUPRa6W/csRmRC
UXOMVvn2fRxmtE+Gpkpc49coClpIbHna2rkFYpRmTaPuv0YZ3MVTHOCmTmBl+/ta
PdwjRHMlfsIJltqZYR1KgGCRj2rTcVo2nu6OO3Fxz4RMyXoowhOHJRva81GDMRL3
gX8EbaaFFNdcGvK1pc/cnB05/jHm/LgzO9uml3dXWYuSzsyAon+jiy/+BTLC/yQt
zYLwDsZPclQTdUMmN/8JlP0MFAypNqrEbAofQAV1FbEmxKbPMg0sO3DdOYC0bcEk
GDETiCXgxrhY116Z+J6ngC0ibroFGn6TeABsjS1+MxqqeY5tNYoI6GlxolaLGQHz
BtiT0pss4lLxaATxCaRp26APXGuiPI3M/rBo0tWW7c3hqXrA4t6yq0raDZ/Kw1ZO
EeGPxvuvAMhuAirUXVxKa1EuFB0EJGiuWzrP1C8KILWyrNLwUg/6aAGrCovuqARd
rE8U1nYVpw4C5AmfSTGY6Da7emqfRNJOIYJA6fV8r5FYgpFjqZUrEgAawPodWsoL
QxKtNIUBtXpo/4v/LByuPfeNhHagu70+eLJCsSj7F9HYdvCzKnGiuZThw0i8xBGP
6UWUDD8p0lP2I0BzliDLtmdbJFqUFS4FyMGGHgoW+XWM42gL7ls01zLQ0ya2qhZg
p0brfQx8dYrGi1DUeA/OHBJNF7IVx92p5RMbKsGh9TY2coMq0Z4PSBKU7WWSGRN2
7iQpTLvY/Ck948bs7H02m3eVHy5heyMDWqUeG0llxvofdJrSnXICtCWhC64z/S9Y
GvPmCgbXu6NLqn8sQGb1/V4d2ptS39Wkt/LVkchOp/6OPa82CybhNThsIKm4YfrI
TAaUZt5k4PxMgpjamWLQ9QJ/R8u+8fjIh6Q2FO/Qe57XuQzNSIHvy1VTmCHAW7wq
LODHw3P4yt/UOQPqHKgpKSSTxcqRwqiZhYLlTY5Ge29vE5qwmgJAknD5dvXEZIDF
K+VsTZupw2GSqNFA3gRavwJAdVLLgnqH6tAF2fBB8CGG2C8D1ppGK/BTnKEPbgq3
80hQtM3m/d58nyydb+iM15bXkdXJE3pNqjkQC1Zdn5eoBlYGFsNRkhfBMqUqViqt
5y7Pl6KM9JHyqnkTiOhc5WWPyQx1wsrkrhuHce4ov/VOsM29DFQtRW1ipcslAF4B
Kmh0DZcvAVXscojFZtCEhCJNGAdUlHn/XQfpdV2DLQ2FahgOcCEcW6MFbOGRpnco
Gvd/nFcyfEWHmCyFhas4yhE/1cy9Wn29dqYYiZzNA8S1BMGBL4TaHLKLLRqr/cCQ
LPOGHFO5VX4mcDmlBaByQccdVUIwvATzvnQCC2O3IgjaJoLkpk5lqm8UCzBIQk1z
wpmEgKZ8KGZrUE0c1wo6M022YrOyN3B5jOVEJ5il4Cg9Jz3WLen9Txn0OR1qBmXx
N85yrTsl5iPrinr+OfkIdE7SBbK/YClSmoZ0CKwBS3lB3lIotWr8hnxabojZXlGb
O+LUSW4ADOxn4TlslT5IIDNqt3mkvBD1vQHyS/SWdqOg0+pdK/uvPRUG/i3vk8jl
vwew3ceqvP/JQg5YU/K3UHfrWIYxM1VAkLMKyoX4zyhgRHmQjQbGO6a7Lx6247u2
1ExVIPbWbENs2GqkF4FlJf/4dMAnBDw5W0FlqH3MIqea+DF45XwWqh6RalIHYJ4V
ALrfENY2w2pOkDtxsQQMCspRu7G8Hw0EmYs6uaopZ8VXZZIkezVgsNQ2vdnsfABK
fJwlFfRPwG3PsjrjKdeMzsP6JlN1dPuuW3PKGlWq+y6IdaREMpNCwqlu9EL6QHhq
PEyZlF6csBRnymLQPgL8/22owkMEMFgA44EvJrCx/PEpe8sCgGPOTh0xCyDpUX4T
LX78+PkUeL2U2MUEG+4Fe4HhhGRJ1uyP8q+ZP3BpafUYXxtwEtBpY5Ph46bpeNLr
xCEd+XSpkZGGcEH3BYk6Kf8k4XoPbNOEJkoqEO0A5U3SISS96thJQxu/qStoDTdt
1XYXCTtf66TLjrbSP3VLtja+LeHJ+TOa6wlccoYStgVcf/2cg2kX96c+a8vwNj9e
RqdSo2uIY7tM6ligr51hK9dckbptfBMPpFpnBBtsY71SDXbXFa6wy2g2K/0MdEdz
FouHmmdrfQahxJzNHjGWOKe5VeAY1hCF3p34Y+H1st/iekDA61OwoiR6vNEk3Rrz
0ZMv1In1I5GMtBGDWuhsW94hzDF18J6GfQNsW6Q8VIegKj3eV1axBZJa2g3jKR0N
mbiNLw8plehNBHexIkUPAk0PR03kqTcD/oFzdIuVN/ZkD4ryuvHsgtQgXJ21zz2q
aYF9iXHl6elcttX0GM7kWr9xWkOR//AkaLAAjP4taXsClqAjmk3yGl/okT32niAI
Ogt/xNYkNj6F7TqEDmj+e8NJCOwgb2t3I7zeDUT6yh9jNERwaEBawZEyJQamBXoM
X0YCJRQDf2c7X8ik7P2v8EiE+rohKZU1qFNI5JH+ReioWMlzd8QarKq5jfzHUU9X
NX6I1sGtdSZps7PvmFHIFCR1cNt4SrefFZphVENjf+XoV1G6/TOBBJcLXYlyXH+U
4oty5oC8J0Z++Tv5oM2xezZqEMlhKOwSqavvsDqXWtY5rGjxlhQluZ0NT11pZKUO
4oNUKZhGZPEYX0cb7Ad9ziTIwW3WzthlQTN9wP/7/BrfBFW4IZ17kNuBqiXy8WiH
dJ6OOX07UF1wxPfYcHbNPxNAmboh2WvoMZa7MUEfgf/Zw4qhR3STdG0yAvFBIqlf
yjCf4YWCJ7nZLtSDabHv3ZLbnCG5WsGz1P7tJN/PdODLCHrVJLY/XdOwiWI3bEej
quVc5EuJXWrFtOzfGG+UQAPEL1uhbONrHtx1h+8uFzHS/ZQhojS2Cu6Bl2X7G9zD
T08YJtRlS+FbcmfD0Zi6Ad9Eaphm++9hSTUsb1dHqwysp6zXixZLqh0ISiSzXnUv
N7K2RWsjyy164OYg4QpnhSuCHsA9MlrRtNF32FXm+xmoFJHJn3iz5+lIrIYRx3+P
Tf981f3b445ToCNE8Nq6+BaAyDaJo1f3gVUaZVJJAYcMKfPt95G+YwBetTdI6ea5
+KPJltU04BOIkUa/aI1OEYD2SKEeZF8uthPIuv5vtmZOCYOadRt4pF4ZfwcsbKKs
7+4PjkOkgFsCZ/GsUmgmY/D/IM8mXYUrgk3BC1q8EkUFXj78Hb5/D1Om1p10e4NJ
SI5/oHLXJWWXZBjruvTBQOdwiCQ1gOIO/ECsQOzO82E63MyksApMEPUQFJgNHjkO
/J2kIJfTF3D/pCxET/VKekeCo2qu4nYewVik4D+ELsf5HvUGAU3folHQwLYXgsuc
2HTgAePYqx/nGC3bBtk5xXFIi4Dmnt9Rw7OQqiqpra5zEhcmQ8IgEmg+g0y/GiL8
nFc1xhpxGI30Z5EStHsGU5vT2z+3BRMBdprbJutheOkIerE2CrdjmpkuD+pcpdZ1
FMCPZTA0D6UFaMDNbDbwqW9NzceoyD7GSZiGG5VRl7zdiMz6W1HNovNeYVKUqBDE
g509xqcMg4SDbfafh+xnTM0BcNSup8sQQmBB0fQX65EEQOWJrIBl8CCg/7nw+wWS
FS/7Ot82w6aB+eK7hFjYHRZ4EeYCME4PN2KHyZZq/C+KG4QovBi/91+zTiUQQoFH
AIEkaj4fiDgAm7WTDgXdVqo2w2GRvbPp8uxDA8xNmk45KUCtlBmS9E08g7sv3cP2
i1c3IqsKiQY99paJXK7a66hwDhPMSFaMZ+Qfho1GSdzVntkdJS6GDX1dpoNGFtnv
tpozy+iCjgCHPK2itFwobHQJ6pw9zhenllXRmZjxZ5pOR3M+ev2KnKDHaMWDH0EL
uxw+xm/ZsqF9hJNSgJd1RS/ZK22s8KzUrH8++WJHWCwcmZnsvofCyk3/oc7EXfDd
TY+iQRfodkx43NKjlEPVUYMKUh2ZfIq7mlD1mBcsUDE=
`protect END_PROTECTED
