`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ayrn+At73OZIxCTbvweFNvw8cXUnaz4zL3DMZLZ9GPp3u+KQgeE22jcQuZuHYmQB
TcE4h44vj+eF58+mLQjwn+9cAFSwWU2/supbXFYsmPCDrjVYe21xUF1cq2IpZiwO
9DvV/QoiFZO0RUHlG4iJvTuahA3ElyGamDZZK8+Bifn2sZETpXD+0wJKtKKE5dEA
JUKTLQZhJ29ZsSSneJzqMGa+O83aPkEH9xXa/9F6e56M/RyBCSOjIPhHehz/BO2S
Z8PExY6PJLAnbBbM/tZdYsVLXBzGRTwwsP0vwkN/xaNfU67HjPk2kqFdOUVSN1pP
JvnvznJYOVQMUP7UTKLDNviXVKzY8XAC6O0DLo66Gx4rzZia6oF+nnyaHR++xtxb
aavgPxS3qvAHcEFJdlFFikN5Rb6oi/ZYj0MNRYoQD+yy0hyXsR9Prun9z1WmTZeb
9BdHq00LJliBKRq/+678xlzRA3k99moz8SkbYKXwFDt2sNKNfcsMbnFGyaQwOekn
rNgBZlEnsEBhYUN+TB2QGRULaQi3eeBmxY117y40mla+BGP4v5KRo0H1eIgjXWTo
9oO3kgg9kKQAeOwUFUJjMfetPd3XyliwetQgHNIWraXpW/1MWgRm2CyHiu4s1Wg2
kTy98OFlQQ5oxcxrhcVLQdt8BpkkWvNEL17vPOywOQFhIGYiWxkvn2iJb6eXYe4k
jFndudwxLWLn/o5iRIvlsD686owrq9h1J0f2AcNaHsuicHbu2I2GKWhqZIjhUgXE
WeTAYLmfaeceBZXju1ID+N3QbfIlYKMevdpM7d1wqjkGqT9whWTaHMXIYJ4JoZ3S
xt01c1WCCGEul07wZ1YqjKM2PJxnIw7wKS3a9Fg5qwUR52BojBTEEqdenXWoxVSk
yRf91OVoFMHyACqoJsMQQjxqvgksNiHms2+6lrcHsLKucun+O5Pi8agOZbIIy/ws
6HiYA5M/wwS9LuRlrRNWBxcq0vAiN+ykP87Nn8maZXJSgRrYKqOeZXc5XAU2/Oa6
xig68VfRlVbAD6NifHUzj4L/BaKNwK2MadB7mcA6ZHIfo7iqtuEYMqCtVnslaVXh
c4ooNLt+Ui/st/flUNJcQ/C9Arvp7CPYB5Z6PAfqJmNf5Ifa3jnpxzqtdCANQESH
mH9fWJz+lIwA4otf586ffInCcCZ4BRPGPYw68in+c1v/KZuCyWm3m3yUE1qLomZw
IwyK2CJvmiS5WFptX8tlfR1uQRH+gNXAbv081M1XpW650jPTLsyH1cvAi7lY2iNy
F6osCE3ceW6swMScAMaFVcfi+JcMIchMfGtJ1BWmyWCMZXv/uXlnCZGNyLrjHOx2
AzKkL/88ZnHIUuj8pL6322/AySirFvuLf2Dqzs3a8W88W4Bpk6234pdRrMAFa5A7
nxAos4sz54Kq+Z0/7SOiJgs3jp+QnvRAWsavUmRsCF/AOV61pQ59MXRjUFmz6U0C
u5BDiEu61sUX1BeZ7H88DJ1ACqnPRDmwygowfsr/+nuFALqDwUynEPYgbSBCTTzS
GoKzcFf5Bw6AglYoGlFLSgIJEBTAebswjKKxmJEyN6XRq3Y+fA0n3Z5kVjmAjcbW
uyvCEQlRT6H9qzaBizcI3HOFlkQSy1Xscb24XRrf9V2LPHBbpYjo4wklYbwcJTeR
t3ZuSkwlSFji+XmEPNWt5A0gGi+Jy+HqaJZ8uBxGQMg1Vrxj4pPBNnp1pBCqaLuu
gjaUhw6eBnLqhrrWhvyCB4aFKsjFTQgPkxxIGQ3msCSx2/pis1zfWMGz2zR2vp7E
cquyMk34FAYdaaujxXUMsWCIEMI9fK0+kbxaRoL1hQ7sNheaCHQrib27SFb6LT6a
7BhpCQc0M3nJB3Fc/7wDJcMQ6p7DDvt4mGgeTQiLOrKaB7knL3omCsfEzhUPqMyy
ohiFmayL2eoFMXC+j7Uc/a+frGytdClHQ2r+BxG2XHSiskKKDjHv0D1rySiY854f
qWDwcE+SmCrz55MgmtGoO7Cj5tI7RwtiL1ZA9NHKCrc1hKSVCEmIamE47aqZ7uGe
npfEcW0NoGth4i9CdLtIduiqmmUVLM/qkj0Ae3qJMe2cfjxTjdpsjZnZi/7MmI5J
8i7DZQUwfaCIdATNqh29vg==
`protect END_PROTECTED
