`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f2g1nKO5orZiyFUEbc85HXT0klVM5/0v2F45apoEluYs9jULCbcuqrU3KWph5bhO
UB2ZOPkiB3sZ648aNfMK7eqKsGm/s5dOxALLo5S92qgMz8b2srcwtYcEEY0GXvLP
VfTEH9YL96GEydiWoZl1QudRYFs6zt9vIE/QtypWTmG90o3NmjBUPXMSjBZTbSMn
n+kc2r9vhHlY+NoYhUwAuG0ACnCl3JlRz7lGQPjzzrf5OkefcWWR2yvSYZ8Txgz6
Vr05fo+zJHgHT+PgD79RehEbUWA0RCWoONqNe0MyuV6AS6Ra2uK+bXoV1b5/H9h4
AbOPZIoPYOqbKMGYMAMylp/aA3cBzHj09AGOu1rU/mTsY8tIwane1OV7tMljEEHq
eqTXPX6VsDECXy1V7nPzJ4CnB+QCELAoNT6ydW990FLf6SyTFG6evsz0Xa+LCYmn
qKPQhswnxOvcodndPxC0Sxg26TFnDu5d6OSezV62beCF37EPsvXNTnoBfFHc76K2
A9X5UFrtp6arsNFiTez/flOgzMwTOy+Y/Sc1wdYIeGsxOA0iWIsOTHQsjRfIt5ye
q0ahguAA7Ld6C8GFF0J0Tu2YZpqB1pGMNi9VjZBi0o8pAqdQy5sD2fRTPZMcgpx6
HaEgcRDBMI4J06GFaZ35Eq8gp6t5TDaie+Y1a+MSmDr9iHuEmTcvXjC1a4hCvRhY
1yfeJX7/dhmNeZyCO653I8OFmcEKDIJiPmChnWEOlxZkw2jrPh0xNv3TM0iZz0Ek
6pTv7LsucgHrwVdSEcl6sltBwcjBvAbl24maVLXn5/J7kyxVKieKoRGfiFuc0blZ
z653pYJXIMRMjxcYzxdlTgS70fZWK8ToQkT+EF701Dgbnr+a8nUYfC0dUHs17I6A
OVZsI1KA8QLI4/Nrw4TVvwIL3Nbd5/LSqounxrpqPBbTSY45ci5zobCzuv28S2yE
WHEblxjTRJtdMLq4Tg6BFN7VpQduW2ttrEMH3TjMa+EHsUAIZiub8TYQ6FePNCO9
2QbdP1422CYf2lZrHZC3BxORLJXg6u1g1WJHVsa1GB3aiRTd0GsSBHWgiPCUkQqB
yCIYxYM8Vt5A3JBHZ8qYZRZHiyrrLSkrOorx7UOJkoVYCF5VjiO1NewK+/8sDzNi
/pwF7rqJw1PlKorU9+EQYriVsQ7LZRToeNh+tXijgtyb/KiYj2fn1Q+IyL+pCPMG
278N1ghJ5FbbetIgKmI9BW0p87mO/XicQju+xgqPIBjIIUjfvzAkyEqFyDlBh0jm
O7yC0j6fG0zdOb7Bg8wwxerralOIEqOMfN0yfEiwpPGxD0Z9fOxXOQ6klUmFNgxJ
PA38sIg32PFHrsdniYJcvxDLdi3NKQEEAVC48+kn9CendGeHSO2o1eRJmxq0/4rd
3sAcoeTkJVHrzZSb7nA2vIE6ZpvTkBwa1v+Z51QYDl+zTaNBpAh7MY/A/haBWYRT
ITvm1yajW2jJHpJqXL1qzYARPEfjNvsVYvxkThRbSDf7xGSTSATlj/UkEo/uaJiq
txmihPAnn5nXOTXQx3aM1S9N5dsNhHu4rqMmToo3S6KSMETxcBJEI+DnM4dhfoCH
2yrORS1ZZXdlYX5p+/GRHB19BD1C3ZjgHAEfaS7XvcVCCQt+tSAwuyn+tB/m/T7x
m0CRdIWjPb2FUpLwofzEMwrx3GR9wPrLW5FDuMQ7ccXVG5887hwI/bCoUcRsxgDI
o5E49KEATFWaiECgDcC3FvBZw3s6rZYgJPTRh5IN3zPUb5VWN0KS8clJFy0xRS/b
TRYCX5h9nDXS1J4z8/zL6klPlAtAdTOEXfQDTLKVEZLjSzFcC8/A0lCSWdiHka5X
RBnaD2AAwtkHGTqi6xxexiqoHrl153NXsjVZK2OFOPFjbj+pIO1zuI63AS0WAYLa
r+JBHLmzlQEh5rJ9UgPUB+SGIefjyHt2pWFgA5JoEXMf5XhJHrT81tWjcgMdyDkg
YwV5A27/cZQeZOZr+NxaszV2fTwyO4ZfDEiChsFH6ygvFpo7HKHwGhKyu3iMWnEc
Xs6WkaxI+MwITb6MvQOPS3mdcGbu9uemU7yqtlCGC29yvsj9NpclY+Eg1pgxxC+x
JW5Gr5mBWHSZkAkbQFhsE60gqZhREg758bW1oPW6Otf5N0YLgUvO3odNKYmjo5Dd
dhiYqUbHQcpQ1G46PJ8jAV2tMpNl8a3syBgIOOzWpzlhBlKpH//rn9vrq+KVeVBa
oCDPU72yjrDhNsBQjpm7w+1AOIqh2b5TVAk4ms+qe4g8XXq28gLGnxU/+2F3otga
UBhQBDUIuAJhMNfqJBcTRFnkkyWXPWURsG6/20F44vB8XXeeYSnG/Os2uuo9ZMso
Qxh53iAvgram1L3svBDzW2rnQh27scFUOHGlKMf3U5xiiSwKeM+rutN58DMvF4Tx
8dsVhKVkpN4V9E+hzv80SO9iTTuuuAsUCJ9va79TsoZSVHV2QpiKht5+lanFTAgl
1DrwjlpSinHF0y4IV+gQT/P87zBw88btkp5Wtz0QvYiNFmXMoPKfk3/kOxGxameA
+5oAIXWvdyF6iqIgxcNvRSSBRYBOmzL05yn9HNvIRyiG/5okyRo2KJEZuHyWCV0m
UJ3xJvZwaJhXw96V04K+99CgO3u1Q7cs+IVQP7LMK140VcP9A02b+fwOUvWlV1CI
tbLpyyOCN0g5rsEN1J/5nA==
`protect END_PROTECTED
