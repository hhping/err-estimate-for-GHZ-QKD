`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0cnFKhAz+JwzlsqadtBuW2sOKvTMr6oAwVbdvH3fodt39dlYKQUFbrsn4fjbrG04
20EgsYQmcaqyuQN2uPkPOzrF7M0hpqaTA2/tDqoZ0xtRT1d1Q146GH36+nvPh9sY
f1j6Ixm+/0qtchQnEJbYm2z+mXDnHUxszwwWGggwN9zhfAtPT5ULJ636bz8EcqSq
AGpX9hJPezueD0cVZViORfvAChP+lOjaKj/9Rjj5+rD4lj/pOQRmcbVdfGJVFn0x
fwz2PDjNORi8xCX8/FaFEBZ0ywk77u/ntG5ByLfM5DgaW/C5tjbIGlYD+bfy40oQ
QPHNbDX/p4Naa4W6lJkATG5ZGR8rSYFb4+40I45AoFMCEoUqGwPfShKdwUIgXu7u
f3jVvK2KyOwMbeoqcz+Vb/3ohU0Mg95f7jUhSvr5C12TCGkzdk96uvumX9wWhQi+
/YwscITTqizv8kltf5IL0N/qmxkslN2muQYsnWVoEnF36fAczpsdzvUoQhNjKL31
bfzbJtoG7zUtbk0WRDL9RbUNfDzCJ9vo+JWYmJZGD8MW5I0cKwY3u7TI+spDZ1ea
z3R/31kNIkoEN8ZGr5GTTrWymHvMiGi15LljCDVs3XZyAyQqfuM0kvEVcUIex4G/
+kkgxuhD3zaEDm5ZCnFGKLmwXh1G/SRTWTJdhwuoV4FcZoPejWz7nfyEWXkLUlbV
poXqmgPbdNwtsqYsTsCDsuux0g/8QswJl2rpaR1jkK1XEGPtldtDiwgOgYYaKuw7
0gCo/DEbnhgG8WqSwgdRb6RBOam12KXSlQC1bcXpbv8ellGZAm8pAFNuVcQEzUoN
OlDtz7mK0HVpmncA5K/pS3fhJlDkUrdxoR1ROGMXsgQ3CcV3g9mVCwaEs3XHFAko
piJU3YLFQ69f17hvFhoex/bNapdxHVGzSLaDdQiYgtY=
`protect END_PROTECTED
