`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zOutvamJbKhFYVeYtSVbDdA0Pqwg9GVvEFZkndjrgIk1cU4f4DTfkpz1CtZgVNLz
tCOexj8QVZdX/VJy7E7iw0SEcmQDkfdWjt1XTfOmews/D8WDRw9UmEpryVj3IVDW
YUUt6pePWcmwT5MXnU1GAmkD2/+fGUtrwWzoqrRKPomk5edRWTXBRiaImgttiX8u
/2oMyBPFkT3wjiJ6kpTKD+EdNIUD3V45tdnanfrS2ZYO0S1Tdq6Ahds+GC72Ib9v
3sa8Qkx0FkVdLZf2Ekng20ksTzcquI/0ilez0H5OBVfTWT9it6nwRVUzz74jGpt2
zU1H5VN/7JSU9jjcJSyeVfv9zpY0JQvQAJTYaW4NGlgsiQUF3jlHdGKHipvkiNe7
zgvwYLg2xhy/PsMZ8T6KBCRoKDfKRFfU1LhMY66J/uD8JoiMi6BxkenUizfAn0Sz
RJPrL/PfqaJ7G4yNrMLKc2mpswNTSnsFPbppS4curwqHmIu+Plkot7rL/YgejAYL
0R7evdFTZV+bKQSpKsf3M3Ee7SwoYPvN3ig1So2hQlSMGqJoheOspDyzgM5EKjwj
XB9fO8PAE5SUpbJN3Op0JIhY7MRuCDHQcbZgYcLBu91TqEvm1Qy0Sooh76oRad0Z
PqBUATnY5aD3s+Whv0f7iiLnugaJMW/zt2UYLQHPmP097ByF4WoTOC6sycRADr0x
S46e5sus9/UU9qbvUKDPGw==
`protect END_PROTECTED
