`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZTPYS+HuKNH+EOS4jac8VyYugqT+v56tUTAklmAJzJAhiPA9TLwMnnx1rd4vRD/U
VX4k92zda+oZQ5atkExl8IpBYaufNzxmObIo3jfgUAfg8ZohILo01KCgRkapCHjj
8imohlXJqz3kzrBL2DFori9lvx4kC8feA6D4ui9JR6Fq01rWW7yFE0ifTUNX98BP
iD6Ghm0kj4PhHnSoTRL8Uh0Ij7H9WGJRsQpjOtW/d+eJlUm4QKbpwTirYoW19rqn
TX2WG5lEjixTEHjwglsTfxjrH9oZJq1xG5NC64fmnJjfp9vhwiub/mBGoJOxYXHs
cbUsSvpH0z1mi47vo+0g/8qIM6wRVDsLft2563VsgQ+l1bzI7+wrVsJYom79hAlB
nOJzWMJgzOZA+Bme4ITbtaRRUFNoKQdEqrewlLmQXPfom1LlwqManAAdBVVv83pF
HW+dSRng4rbmLnNRtbsMv5ildxa/AnO3w/TQEShXtV2UPrOsbZBTO2tVWXYybCr1
zwjSeA34LXU+fxfSW5hvAnGVsvkcErzLzXDozeipZ3U8pmExuz3cXsKIsonFVf5B
fi3YsOhINb61O8U2ju3Yx1Ub2cwSxS+R+ZdFhmEHsrAYKOPGUrICaHfK67iKgO89
cwuZzNFh33XzVWpPr7aU7ygPHQ6COHwOPaxPXS/6cz1Z3KxnaqCVz48Ma5jniRkO
jNLJBiNL0L2Pp+EIyvkdKCRj3ou7ASNvBg3tQXlbtJjH7R1N2Dp4tVzfUS8bgORY
ZEzHvBb4KQgr7+Frqjdrg5iF8DMZn1C6BX4Qml5Vz2OVloubC3h9BuSLiBK8fLTh
TiTqNnztvlaTPwCKdeU+x6KOoXCwNIdn8rEapie8c0hpBePaXn0S1M7wmrgqsYuU
u1HHiWg5Vf3n8PjGAGx3DABaRlIwnHNLsrLJRK5yQ+m3awPWIYxg3j7Xl8q63qUM
AsabUW0U2LMm0jfUdojmis//c6SC1c95wPwK2u/9ji8/g5ZmfZzu0j0mBKRmwkmU
efDryQV3JcRijjoPv8RM2mNGDdh7/HathJH3OG9K8X6RxqP6DsbbL9GrT74fj2hN
lnRMeaXQrm86OSddJVPQ1FNoQ3J7Prlugc4RewHAsfPIMAx9/2Y17lXyCI10ejju
qnMVzv5uwdN69sTsXkQbkCFqcRHEznZFsOcYKYPqgEId60hD9puWfxGqKmUeesxA
I+LUQbsVO2L4/0BEX2fyx/+evD/p9DHBQ0xaK7j0VmL8B4OUCWP+eHi00lFJq9aQ
0P7fGgfYHpKMLAyHPOB5ox9DBzmPz4kYRYZjnNm/ZUYg8n8PAps3zr68c5v9REwb
nBmlfQ9Ek2jj+pEVH3rPy9m5MGp36OPG5fFc75K8vV0LNEYFk5UY0RFrmwDPFOV7
vgLJA/75d7gxI1DgJsmFKDbi3LK0ZUC/Sy5P7ojZnvETEbeD4OF0fjLhmd/OwPgU
2ASd+N+t3s1XYQcY2N422g/4lPJpq0x6SimExBjKV3hjy2QIXoEG6xCoEybu94iQ
f2XZXZbv/g+modzI1Wd+Bn1idRiklRobr2ho3PY7bySq3x8QINe7Z1CgbWKRMaKz
6NNrTOWMM2LbNIXzJh4Fu3vxwUw+ppRnCRdqz+vBCe64VA/VfhbCH8nRPg/Z2ZD1
It7XJtycTi0H810BhWF9859idbTS/QFw+jImB0yBSgEeGgLXRbK12W7NjrVwdow/
jDYOh3u5qa61Clm4Os1wQO1ldFyfLi3GGbRdDRQfvLB4GLaG6nNXNLdFjTAd2xD4
VXS5OusNUngguWzHqSLne7OM78vsrP3opDhUynMpwubir3TtRn5aMXlt7sYl5xde
Q+0H4MJBVmF7JJFF4Qm/kMveiJYeSLis+z2iXTwASXTvSdnJ0jn3xsMW60UJluVv
HkHRT1Rnuqq3zwDDqXMguq90xCyO7usqDd7kOhfeoBZh+UYvo969qhuvVbEGJkNY
CxUDYa5Ufn8TQBzwngrvq+r8g0c4BB0fMMc4QxXoMHduCcqLEJ7vpIrYlmT1m/+F
9bXkn4ExDlwB8aoQGMRWmlwYcbBi6IRWnPx4I0FiKAvYn13TzwPJl8MXXWA3p9+l
TEA3bJOIFzcYUKJcD9qbhO+Lf6uN/Edn0LaAwIdNlKN7akALbkXCU3DZzpUZNRB1
c8sIcgEoufxaIbnGaJN5ZmP4g9mSOIMkwDd9YFGlPLudxndxq3uL230EpLZ80o0m
O3XGavPDb/3S09HpKofOgEe3IYpDRPv2Q5lQisHwZcsxRFaaHGKNgVV+pqK0ifvI
6hbh2iuyyYAyTgBFk/3O1M/7k47v1C/YO8GJSz6z1PCwkEzi89zdMcpd6UGeTnVX
qE1UwYIuE4uOvGZilEV0uctaIbv4iQCTbg9YKzKOuBBqOtcE8ahH46fWCJifFHg6
Y93McOqB1plUHURmpdGcQGDWNJDrafYJK/AJGW+4MQnh5bQjWHYVupZl0nnaFT/N
cDvnjlXdMGIbKtXEpjrv3L6HQoohnUpn1BIBWeNhhQeMmpCyazGkVAVyRowRcL+y
rLA5X6W/XnZM2OYvQUfjE/gGXre606N31NzW28xDRnsMPMGFrAbvIWGzUnN5wdpy
5RiZYtwbTh/DFhP2ljHXC7leglFfQKQA9b0BeLms9jGJdMWHYZyC7yUIv4EbjVbS
2OQCEa7YACmMMM/fvdsof5t4aw1/XZAiWY4Q7HttwwdlDfzuOayfXcFsjp2p8WhX
cFPEVy7HLUe1fGjX3Hp7NzMygyO2x56u79QUfIE8bXafYVFp1zu/xZDLkrCuKmTQ
Lu/M1GxSEnUa6LrazfoW6iJEdqsn53faXH4MN3yS+RQOrA77bj63PTsoKMFWty9h
yxelWTvNEW4Ifq+TRwud1jDNaRbGb9EOK+7nVUoysdu1AlrBoVWt3MR6DvNd+QVQ
EgaqFSBFtnE8zUjwG9w3l4y88sm3hyBz6tY4ls8NHkaQuKTdu+U0kJynm/m7Jg3U
OL2AJqET3YE4by8Q4L2SbQsZ3rCnk5AlmPDgMH6FQwtivroSsqzCmszTIrzAw6tP
BzJKgOtW/Yov55IhV6Z7lssgjEUfNJ/CkRgqyl4bdaUiYUmkFjG6/m/EUL78W7Ig
3kNOmYMaLYHlQkep/j4dRbwB6e6YkTFr+DQub5D2aOVjLCpMuu+Rp/OUAmqbvffr
e5kxnJjUG0a8JdaTfu2A4jolL/oSrGpgsBuCp4dsY+mteeDlUf1S6yWFFcXjfRev
6hYJGsu+9AB/G4CpBTwa6ZuIdQPP2ifr3Y2ZGWUu2TTXGx6vVB4unVBfu8VACDQ5
F7XbLvM0n+axdGSAytwqRGjJTgIC20AZY5MC+8+75uLZdwsPIAKUee0j0fDB9qTb
aGuM36XrDtDdhEAGVprYWZWPSFps0fWOYrACyDd5V2Wnf267yo3zW3jMCc9O/3Y8
mrMlPgsATe5ePI6n180ZacVoq7bm/PGg7KRG2OFAUrIZFYLy4eeEyfmm09T7CoLx
yo2bQ+EKR4WiUYASG4mg2pwaRhnbpitr996H5xrKDuRUTZbg5KSHjOLyzWsnfbZj
L/cctMiWUiZ4YKcL5RPw9jNmYr+E90otAu5L/VFp4sgp0z6stPwGZKoUCS30P9L+
MYo6qTIlfYcY19Wxq1fKPw7zgrNaClKXnnUKptepLZ/g2E3mTt5MDwnyenRkg8N3
o9ALxoaQImUozTzbqprey5sVsQYkC6B4eA3W2o/psxnW+Wim9eg6HdrsSfG7O9Qy
TUbimo9kNCLSyrTrDfX9X9ZE3wecA9K5b3eonUysTGhSBr4hkbn7E3nkQLHlmnlF
Z/jLtpJc3Uq0EH5c6n8iw8WZrRylCmAnFiG8bBILQZzG4edFZfOhfXDU7l3ge2xD
DFUAv3lI87oRR29wEVFZ6GG2GPolWZwj+Q7WRr8fuUl8jnex7Qjd+9LijQAqC1HF
XtTasqZ2PiG0tj23kyOvqPLAolWthZjuoZ5B7hQX9glxcy9ZPBONIFSFKuMlRxNw
CwUKSOgZe3oHIZ2ZuE1oZSeiUv3PC83Eu2XZzABy+vM/hrKKihRhHDhMO86hqVyW
6iFXwhnO0wtJV5wunCdyYROTbwMczZ7F3NnduIYB0ULldYHrPF7iCu8BKK5CC3Ui
noZEEM1Aw74BiBQFqe4vIIfl3CTkbaAyCpBgwGwM9ZaabcUDtPDYckOqVQHJ3uJh
jn2BxP47xJhzwTsdE2Yz/pvue+PZWZmVw8v54LeiPuEe/khn6p8HizHfn62GF00f
h5GXDC6wfJ5meA7kbz47zUlPKmYhui+EflEcDQuWEQW/tJpAC/Nz7my4A94/sy2s
qxujBG+bD2Gn4S4A06PK91hFw701XHhSWxh8IyAAIgaZN98uVTw5lZLkwODY3wVw
N4ZztdWzta3x9AK/zLVA9O//rm6oHy1fVZf0SD1FmlVLfWl64K9kXiYkGaryg2XU
4yAr+v72t1PIlkUb9oQKk65MHT8Nqas1sCB3dZMfAtQ19fHul3tL0IxEdzEZkPay
JzVWXniUIogb03yYmW3APkRsUHwBEqOvCdLY+eMgQIRmzuByN7uliJIKOYsJE0HT
XXU5bPIZ6oFnPZN1iFCaOg1GUrtLihc9YknObEOmhn073G+TrQdUm/oABQvIXWAk
EE+yNB1UfFIhPtFujabg5yZehdyh9R2eW96chvLIkdhT9O0Eer5Js9hG6AOg4Zhg
ddIxMBfQ9OZ3QPBodNYif5Ef212qAuTUAtl4S3QiKxTm7N5sCopHqsTjFHCUFK9X
gBBsjAswszGP3T3lkfIhKc3h6wv3LVtHs1psONA1U0RkSrAwxfKiKJr/bGPMM4j3
y1Nzhge7C7OXAzuyTQ8bVOloefsubt/UGHQt1fbYsptEn1Ya7/Wwx9UbZjg4qd1y
mt7JIl0bLQzfCIFY4cdqC9x11/ZFPQZ95nbJ0LeKPY0HiLCRgVHlGD3HLJDTHk01
L45YFQGofAVjg/39gXknBJNI2D0R1fDN3bsX5Q9X+fEdU9X5q+jxt6j4f1tl7H7E
IHvev7sAS1qT83eTkCWZidsaENP60Jm3VrexcpAC7Fk0VZ+lejTlVQk6wFUFTovT
k7qRFab6VnKjdTSJkDCtkuOXwWZfnAvqSBWMF4ZEyyBVC+HI59rwwsT2enX7yzWV
m49WD0/aftAUv1tambpnqmgEfVtNXGbGK9cqoQi5G0C/K6G0pNWwS0JXhEcNhK/Y
2Owlr2EhLRPZCU8Z4MoSnvjpsPGb5Uo1De8raQo3qkMK6zn+SQqQGwCzUxP0KHHy
Y5v0ZsklNAS8SlwCn+QZ/X57X5Ojd5ay8oxLLKDpyu7cUDHe8rnNiAU9Ps/+iKge
JPdX7ZFOMiaOAIXM3hBY/2EoSOIdTYt37j2Z0u+jtAnLY7LKCKNVkyNrRGwsvBM0
YRcysOdUPXdkVj62PNnrQkR3sf0/SLr4Hgcb4xpatA3Kg7IKn0gxQUqITD6xzs2a
HkcenhvbInlBh1AZ4BkjJfSjytfSUeFtTLGcZX2QRaGJ02h61pkaY+tFpr5E2QD0
iSTix1AvbQTXBTxeNF95ISFG13pCuCPFzXuifT1OulCOMVEWrR6SyKzepr1P26Rj
f1NjKB+JS2rGIuGQMEdPmXFHPuigaJwuDPvoY4R8sMBqjYymWzsDXjLQBkYYCWKH
BYFWyIXaGHcIAiaCm/r/cXZ+JkcMm4I90iIAfqWupB6xr0SOodj5yhcsep9eEMOR
qcut4iCcbmuEVBYa24+8bRqD2Acpc2Z4PbPMX+Sowf1LHgmqb6nTDVW+qp0LhCdH
kzkRQJpJmNbjxz0mwIP+WIAO+oVtBJ20ngUcbXH9g8pG9zP3rrsy2DqMFBUyVZsO
Xp4WdhWobqtr6pG1AU0jpWlebnWmlhXVR6nLqxoKRqPFiIVYXaaesATbT2gGPJsi
dF2C0K0ObWnthpk2JZHblw3sYWdMzE9HvzJRhYxxRkNoRy5wRh59+eTNqkKmaUTs
bjCGUR/CyIBvAP19RjB+70RlGfl2LvPfJqRjbs2e8eqv8Uv/633b09VivDZHTfAp
vCVckGjjjL5xawOV6m8bfP+UiazyGekX/UP/UU9yPRUkMEnu17DMxa2vpky0POAk
Z3GH6scZP/vorFJvviwp9ZP5MFeB90SFei40rtzX+ZRl/9m4aPyCLr3aYHgQGosC
UQafsTuxE/yXeZiCPZV8ZyIAV56pXU/3rnbFuSuWAuXz35SQycFo2eevlndt+wlQ
PjYj4TzKJzBlF3I7YODb/0K7uLiYSpJQpwAl3gNQGdxFADdZ/WB655jRiDRoxOE0
ahQ6rBLdNLz4WOjmH30Qo4so3HksS/zcJG3+c/zdaNv2vRJCX0USLgqqQvLRrQGQ
/ky4AQvYQckdD3nP2DyqZg2n9+kS/1FATCHS6xLBsv2p5BYNwC21tcPEWt380ThC
V9in1phhw0LcPoFqiIzKYvfNG5dmAx/2zM3w//O9uywIcCbzaduIrOobkL+V/7FY
kVSqreRQLHYmwG0g8PdFj9ozU7FjSBIuNFejfzdEd4lvSnnBkD8qvmIwoPRoB5L0
E0/OaFMejmMEzw54OKsRr104O1HOu0NaYPEn5i0GETnI+bhDJJddZ5BkDn3isJLt
VTzRiqRlHHD1nfYEIalCcwWOJDf0cdnHN5wn3dqQKRmkYVMf64jVUd7UhHOGq/7T
z/w0gCM9ko9CVPOIwRL2l219rzdpmhEJWeGAM7vOkD3ON1SZPUY4e6riZ9o/29RU
R2hVZAY3lrHqpPfXzig73hZHKjS9MAJV/T5qXwA9YXVXQaZ4te7tN6plD7eWRN9i
0+03pgmNZ0siBSc3r+DTIRCbwr0USgtkUM5RgZLxlXg7d8ORP7tiWqnYmaXg5uwr
/1y1KTaN2i3JIN6e/w6BAIIjVcABti2ZuS0JJ8J2LAiul98XalvDYEMURV3uVBW9
lrk4GEzSYF4/dQQ2oOgKjyhHrXmRsFTmnfGiKt8V7ZDBvgpR2AIJbIwTJMNk3ZH1
9e5mCReO6hzTaZOxigD7Kc7OBQ9OXR0ydYKbr7GlHex3HVS5Paw51Su3/wvOj6Aa
kzb5feXxmUhrR1y6eoRJpkgEQ8f4ub0KF36zupGbcuQq44XiFisDVnJ8dt1OTwoP
dvuxwMSYtT64JM/Uhs7gnPkz3gVolJaC1fEUZ32jO3d9C6FqVgIsrwNQwez9ffnJ
SVE1gSGzK9sIaUhBzlLuA+1tMp8QUqde9sFt6kCJvTalCZYGz8taelcc7EVnmDo9
Ju91yH4BmClMFxM7R03rZMpK+G9SYG8fdLQ3bi2EwqmMmKIB8mH9cj/R1MY75IOM
kWmgm4ZK8NFSUq+pw1YaW9KQKNgtAggOZcUIEn10LZKoui5rO4acyvtmBsPCLhfq
1WuDrPMaxAOqPIb0CTBLrJ95RAMSMvd3mYN9gpF6akGXfdFR7Me30pYl90h/7h6z
N51bpDk8+XdLEOVesXq8sXjx6SqUm/OACvITkiH3AH6/WvQKOx4nKSjEU34OMqir
uDcU7OyEW2qG2UGisC+OAln/GxCoZ22QcOVlme1KltmqgepYZTQ1R5SE8BXUbChb
BYh7XW37tfrzibNSXnwgcDBS0S2o6w6Qe9pBN6VprJpESWWwabGrQk+D7cvE5uOk
2hCQaGl0utjWxo4qvM3uI1oIS7RJTp8mj6vOpYuphnRg4ngYFFABfYfjsvvVyr9E
MGLQzM5k1/yH37a5C5ASGxbCyaaQR8aDXCtlQNjaU8nJkGtcIz2cYjUjWPaExleh
/erSqbFRhuinfDDZFivcwJTX5abzk8goJ7anR+xvRDLcJx2JPI2uiGXgXbrhP93h
Td19KuFbFRcw14BjytTDiriWQly5BphOJXWgVJavr8xoRtk5tN4tfn/blC2wkD4k
/IRbDEsDZpaqEHZ90m2BF/6wuxbL89vVUzHtydLIYU5R93dMBhgoWA7snsKE7aS1
ZpppjiH8Pxm8ufwTdgJ6V4HTPRfMTs8P4EvEJDKtMyRAey6CQrr3Mcr6qxqRapI0
nvQlhgtdpGfDn+SnguNI5hiSo9M3Ce3dFmfdqazjKpBoHvSIkD21LWsjj4wmhHSY
MmO/I3nyWcpkWZFqZsPv4eq8fuqVLfJ6aIp3OpWJe7NmtD+d75NegVXeQYuoWRuJ
ieJdaWK9Uwly5qrv+IJXmX0n3Et33XHej6rE3WaztN/IUw0Fut2raSSFOx47Gmix
GwT4hPuGWaWhvKtYJbIWpznKleYophJjJJHZWHwIdtpQwWz5x9rttNZWjyxBvgjI
3wLFZt1KAB00l91y9clEa2jPhbvIG3xBDsztw+54rz0w+MrRy8fClNJM09YDmJ89
PowGXxes0bgo7/BfzG8DZRM9Z/yq/1yJN5n+cLWjYZ66R1sF5cDUVnKrkLogd0yo
QXqO3r/ER+VAZ9rLyNORMGvObecVvB+sVqQbIWQxCIr/xV7jqKF/7P1NHFRe0HgB
h/j/ncEybmYpseJUnUOFMCfbxmSQrrbreh45gA0t/X5+Ec5IbqL32GhqEs1qypem
QWn9VuYwiXHGUTR0VLuA40L4Bb8T4O+yP8MkXx2b2R62IyKa/CcEIjcUXWILSd2j
cH7qVMaahG0ONcGCXVk2TsslAhSYEDRZj+ceXoB1dF7Lfd3/Fb9bxgye8YL38OGf
T0OIlMKIUVd4JjJ/pHkpioPo4k43zQ8AZ/DsH2Tap5rKukJ9W025gmgkk1dTNX6E
Kntui7QmaQm49GCATEjSdL4UlH/skOUTdnAZh1aZATrF6XcYCCrzgEwP70AtoZfa
fPE3q6CWJND2qVGOXnCKsCsDffdsuDG/7KWC3av1JRzZ8ynU5JelqvBRWMOcxvcB
wyKqu6z2fPSBEIcXnHy0/UzHjaPPDHEvQLtaGlueVqn5pAvJ0bGRvbW7O6jDMP0l
QEwIMLufXeV1yqWgroeaDmopVcDsRcXLbn1ZQu73c5pPBG3TkJKd9ugkO4XnbcFf
0YP0dFFt4C8xiwaSMubqPJsitOWrgF7ZFHq5/kmtPedbTyN2TxJVmu01OGVa84Ve
gCGeO3Q449QcSxi4Ekzh2RYRcBmV88QE9WGHev09ggYCg1AKFv0/l4b7nyYV1nLr
O1uAQh12QhuGfxSx2xsBwcWIcwd1gJ8q4RpFB/TDb7CtDJLWwflth+mexXE4CiEP
TTMIFkgLxZGNLUugLPVX7eW9ayoyEoCz5+WP1ZeLE67sOhLMpQO3A2bib0XayMzl
EW7KJhm+FxvIitb1Rx5wkMVFhCzhS14cbieVAV2ncsmNTHOpfpfLXq7EFynK7nSl
9TJyNmWsHbRb0G3rMCUFnlPoWgqvZCFBU9YiBYrDI/xmXNOh+JBxIHf5CuPoeVSa
wkvAnCbTOc2vEswWldbCjPE7mNHK7j67xU4N4GZd/VR3dBl8kJMdd8V0ySZCH+eA
E+82i8dbP2038f0XKYB/8Mi2m4D9pkbPkMV0Wt0Wp6IzejDvjwKl2ULUXd9pjZMp
Sn33exxO28tmB8Y2Epn2LqnfjfhQ8q34D1/Bw8hc2WeAKPpyz/HvBOze8t7kepy8
vd9vvC9ffYxHo8bXwtgZFhGy4zI/fkmtp7NU9ymBdbLEcj3cLtC9UkJmaUq8lb6/
tAR95AjxxqX6hBiAI/JqTjNOyaj8rJPyrwofxa28KgYt2L1k7sebSdRhiDgfJUUs
8PG+Cmg69GqhCfURAIMTUzstlrJI+U9+elz9lmLX08wFPVuoT6if1xzo8w28g2xJ
dMocBkC6gdsdsq+pdZdz/LRPhmmF8feIw4ksukag+dhXFPLGCTqmx0HVyYiJWhbv
iEsFF8UG71+vkEpjW4sSecH5/mNNJqOjZleLnnp6uXlV99GLusXfHYMa8tU0CLfb
LbnF7M6exZjf+WDlnDy5vRp/udXbI9FpaauqVXG8oUA79yDyrYBpPH7PFBoafIix
Putvc5ZveAn1esDbqBR2+/hwHrBGHH5n8YgrVWHBDftZ6xzGJg/w2KCD91c3gLoq
64EUxay+aQG87wmQ6T0C7ZyfTBuck7d2J3lMDp+Ji6+9tyaN1TBXPq4PWrCLhLzL
/MelskLYud9Zo/43nRbJ/x0zFEb1B7ZBItZJVEWEnJsdMEk/aOAF8tuoMhQ9zh5o
WbuvYi1cpGPS3ioLO9Dzs3iqEOVTFvRIvx0QnCrix4KtElq1mkg6sKfu6ie3KaYw
L+1ULh4VeHR9EpTT3B1sfzRIog/GbEY94vpvmP4bKjT5v6TDpp0xc+K5lrwuxieQ
oyLGse1Zrk2bNebD1PkjTyxmwjb8spmaJ1/fz1hpA8qoAZLGGtGpuXOEIKLumjjO
2Pt4WozlVCmr28+ZUPeYE5lt94lZcaBQj8XTtH4xIjs3wWdE0FCPkSymNs9Rrsqq
TnVpF7xGwMuBEcIfJTxbe3YnWsQbXOxwn/FjbnJdKYqgBynURPt0pumtwS+5z4mT
NLIVefNie9J2/azi1P8JK/VXY04bFASk/rNfrpoFLLW46cROQ45/Wj+FuxyzpuYT
zBvXttMfg3/CnqQJth+2eJb4gLuvJ7eGEXKVtlijsFxn4oRqqMbvGOf67SFZG43F
WNdx+SvWQ6IhHlwAtyGWlL2/Bnh5V2tZFgYJeW9xhIE7zDHI9FRZUeFPkNzUsUyz
nmXkVlt60/jlhq3/ku91Lyzf/ShbaFo/so2yImQkTvVG/pS32CYJ6hSYjIR40/r+
vlR6oURP77aRduaaA+o/dnqqL9IMqH5QF+Cv3Ds46C7/OL3cZdXT7WobcfgS6Fe2
uWFlMJ6M9l5bdfzvq1I75P4JedxtlKcud/M7opPToqzO0wzEqyHR2Vp7pnGBIoka
Cwh2AajZ6c4uYfl6GO0QPuPc52BDL9pPyfWEpFTQh91QSSCDe7G9VLbXSzaVQRKD
oCY2RC0CXUuIXNnXz2izR4TZmw/PvV93FMGJQA+8r0Jhg9PkxWHLgLM+xiUCBnj/
q7/QxTAOfCHFpybwyHnw2jEVWIU3v1ALz8XJhLcRfc/p22Mev3Ic1czvW35MMJko
Kl6ChXAwfYFeYY9UcOGDxnXgcAeQnrXCb3Zfk2nmFM7OnRIdTfBj5EuRa5P9VYft
9Muev7Tcod3fgwdeZozwgTNDET8lBfW6iEkc6cuhKjwjuucRjbGWrv3S+V/X5WVm
FszvyvRqQgg6rHQLDYAueYasBmYS1Cry6Fza3cRgsK3Unrk8Wdg0KACSeIF+X+54
CMG0DXCcD5rRIG7PqbrZmc8POMcflOT57kwgdOPFpSdIh8xPq+q4zqjedor3LaFB
YzCTbaNhyKv0tUz3RQpZJ08A+4QkJp5ITMz4g8bgr/2e/KfjjeH4qfEjsFhHcgH5
rdfUK6cMv9vewl3s0reLZ/9zt6YLYOqAzOS15UP091TxXbgRfux5AEiSZsB6BRPu
llpiUTWYCKOnV7QQ2BNXeHefaJgpzS8B3ckkDLbXakq/44RvSdWqMz5ljogh0EoF
CxyFTZ41xsIr1+97hmwHKFqAsyUmMLj7FdfluxBXl/VxA3Q8ZpbKyljK9NF1TWGK
9WSzJu8W9522Y4w6xLN+rWrJ6V371norYBOGniZtkgDT657/MgQINgWq+rLLYJsc
L3A68crcz6dc6mXLu3kqMSBfdStbqnzptXNJOeQpyLDEvAwwK63W61TSg7DWHkhz
oCRQRBYMDII1KpKjTf3EMI0EESbi6/FcgrwH5BpVc7AdJxh/1qIg+8t1S+I/7mMo
7nFOt6uxWFQIIgu5IixjOttT63WCwCtwrFhmTvZGSEIw3BY7mvkE4LkSZjdNI5By
4zFepql+ejPqIpZTk3J4DLjm7o9glSmXZ/p+ofAp4laKBUD4U0jEmZiZqLAont4a
bmyH41eCrRXRI7pX9Vw9wJKDfnAC1Fw27LMwGm9p0/KRl4JXWkxUmVvl6oyCDZT1
vW2Oy7VUXJ1s5JDiF2yO8A5L73geLFYehmJjOqx1v6bHNsCdJN/9iqT/cDqEZX7Z
1HVSg4zscV18k3H8KxOHkr22+QgIeY58gIYHRJ3TR68FmLJ3kBaQ8QTgSG1dIFt5
6xQ8/RAivG9hpg31KKo4hGK2i+jbbm5PxvQ10sSGY9t3IkAOYFqxwoL7IcHpCdCQ
8yVsaJHju95/rqzR9kuALcp1uySKaXVnSXRNqLgv8IsaewbQz9dpKEw3dXp78Cf4
qijT9rBiPsm1hnw97Jpd9Y6hjrH1biVrespG491tldxxlWIJcwhSTAjNBxmlsau6
CadtRUN74QlkSHO3+znGrSi52I/FL23F9nWb/MIRd/fEt0PgiRmafcT1Jhp1SaZc
uO+cOPke/GMgFqCUHwzAza1AoZpfCIzMlM6gBPkH8KHHiR4WoSBUMTlwTh3s/cjv
8VXuQHpM7ZSWNsRR7iiEWERTKJ748Itd1wVA3k2TIkPEB0gavavMdsov//CaFgSy
Mvyyv6Ukg3VfJQ2o84GhxCtSllTasZoAjZjpnN3+KL/79jariL8/+BZObnReo86G
Fdqbe6ilFcnZUEJfG+eZi5Dso0uy0Q0JoKpt1h4dB0VmWBUOtJeSwN4kPxkTiqgZ
c3unBzScwSFwYVfXnaWUndNo1WDR5BJqqk0Jd2FfpSymXvfcFK0K2CQlogW6JzJ6
CLdg8VcJ7X2WrIeKcD6eX7komw8cUB3c98fD465EiiWgYOX1dUWLIIvjIzPAUBFL
mCpUs17oQ3zh3lkaCvpooczRguI+JM6pHrvFzUUa512HBrrKvBCPHuDYq4QlW48s
Th8ysTHep5IRnbB9lXLo1TKzmvp6mAzEuCbKktBgA3DKS8DZazrjvI25NhtCaRwK
iirzP4gqndQ5WOpwQuJc+ZgYqgNay1RH+hwW6IQhqN+DL5PCM+5NomDENuHgsIOe
Utwu3yhAtyr595Vrm2NwdGSysvmq3H3mNKGCBinJVuLUGVzW2wJu6wQdkao7E286
jVQeql8OESE8RJjuqdDcY80jA9WCgcl4E4t5W1UaW3Vx+xItgau7Bqk0d7Mbbg6T
2Vfv/X8+/Ogdgwxdp+c95A0lC0pZbK0O3ABy4JC184eq9WRZUFak9hJXaLZnNsOb
o59F8GGMZVKkVOdb+6cgy8Ha9nYmA0pXBFtXzV6FbC1t3JZXFPhdNLvC2DD2Vg1p
A5ZmX2CenNgWirhedBDzl14NROmP4HPKyLite3Y6HQLo2yG+7aCtt/JPpQElrEtt
Ghlg3Iso82mEzCn5PN/IofscKmXx2u0c3g2YFivtY3QynXGzSfnSZ/jQul6w5dzh
dyinCLZUV8mRbgk7nwhGtQ==
`protect END_PROTECTED
