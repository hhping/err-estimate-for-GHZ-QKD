`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w+ALxAsIT8wmrARrJ4pvuUGURNT2P+JPAf98HlEWq7AB0eXvR6OXGdDAiYFONCRf
BkFbVevXU/iYZ/E1CSBljgMKvXzpGfq49C6OlW0G/1ZHrm9ZETWy4aowGUUpbsyE
ZVnfNEho7PUCNcCIw5urLkqlbaIr6ioL8rN/U7+vdXqYy0i6ijqqu6//wdN/gOZV
WC0TdGasZPKuFSvNwU/LLxKVtIr6qSEj+BYpeqnjV7mRNoGHamIp/oIBZuMNVDc4
AQnK3uIU5nD9nCzh+5fvjRYY7RAmBi2wXuZOsZo2DHZF/sRZUdV1VSC20mZHI1bh
EUjXXNQ4NUO6dnSxx5gBjpyg2f2NQXRJs8aTYM7i8TrYh29AqlQ2fRX1uBGlrXSb
9t4+DhNpANBQUTpDj4wai8UhivRCI9h6+0UP/u48w/eftpba3RvDE7GeE4L4vaLD
kz4b3/F6kvPIz0grXMBQIkCHeHdfAQcCEcOvZcw2Gl5v+ESnQVfZQhsrbO6SnJeA
9P8FGNySJ7gJr6i/d6xqL3iZkzeAmJrGVDgql9B5CoxjMECc4jPPg7GKZ1lEt2Jv
5GHryqG5s6uQIpLsmQHKEHKUrq3W1A4ojZJSlSs/eruAj1yhYgt9CYHepzU7x5Zv
TTXZDaqaZ67svV9TBicDiifnQC3zYpgXrTlZETN0Ijne3UZ1T8K0fku/zojC7iQ/
3aAx9PsGHwhP1fBZDZuEyK++nfNMAK91bTJi1qfyUu/C42IVtGFn2+iJCUpBJhp/
J4XZuqkG5/1SvaO9ypc/u9qk9JzUHSycDQeEVBFseWwaLqDKTnb2OXyvizgBP36O
qhxwC3JXbIgUr16noLu7xGDJq4pF87ixZ9rqbaMPsk9ySzacJ7HQPIa9RcDVtdCF
iWlMTooIykrqz5c6qZ4pjself1BRcxXQywe1EHegPGAd/JCeLbW5SWYLYYXq6Slq
cEh+/u2uq+VMZ6z8vURmYYGL6BUnF2wtCaCc2K53hkVtr27R3sd8FrLlYYlTMTF8
gdxzo6CRkoClYYbHsaRnq9Pq1ZdQAT14SobKpK2bbo+htbgypeZYJmb6Nd818PzR
ZouOZEfezp5DBWhrIZ2AmrMPtdroEY2GfRDDPJXTXftCs1wB3U/pzjY8VrfTbBpQ
g9/CE0cWf7JghZ6QXyUAswtaK08a6t7KIhpRAR0vJ6zzlMrJolBLLsokYxk5350H
Ppz/SXawm8yKV6jKrTjLiH/7h5fGJTOoOBq2STDlC1+1QI1VMCJKF1Jj3cKIR+X6
eogW+UHGjbBHocH9n+XIfZpUiiEiQgEAITdy3z87k8rZ8/WZiOXML7JKbpjfnXwA
SY2IrWSp9qKhq2vLYyp/VYWcgUNn58KKL/KwlaHCzruOtQStpjJ24WoEnwUnS55m
iXGfHxgXtM7bDGydSEbGoCGGB6RBCxBWlpGGzz7W0qVFrQaBZgFzNNQKZQa7U5KU
PdewLHRL+e2rXbqxsyRSpt8HPW7M3ZjkB4xKkFfUp9aa2tSKztjgYdPVriInVnWc
2ktvqXG21w/5GyF2aq0TRnPx+8RVlHLdJk0fm7bi63Fij9JRGumQzTPZ96Fawjs0
bzXgORU9ex7AsmX5UiCHgD1OM5vDh1nEyCJ0FobYiNzQ3f40omB0o+OCqQCxfxa1
8FX5iZN8rvYTPDcrQIJVe23ocwB3uyR74l/aQoATS/l6UNvi9RGqh7XQhC1SSGb2
Plh5CJvbVmtfd5jJlJmiGZRV/6Mr5NwCNS9NcyB9VZ0CoXjsAmbnfkrPtkXoDOPr
wuYOyn2HtnlNZTd1lchC4ZcsmJ+peazbGN8T6rQyIIEp3S2OiHSDpsZbI9SYMmPH
Nl8ZkALICZhbwc+7b5o6PosBfb8mCNcREcBObA5rT8kfb5S3snUeEr/mQWdGKQ5U
MzXz88ty9W0qHTzMpXsxGpqy2WuukjUE6IXt2o21YzmNwkeT4HzEHK29nfmi51OZ
5SrXNm0Hdl6ayD3cvtQpmgyASQ5FVzMzS1Piqj+i1aWxfK/JY4ksHpJp18wmV9tc
HcuByBHbVw1+ALGAmT4gwol+5RjfIXPpOvAbfkK3nbvGE0FlHX9fRkTfvDacM+Ha
d3jrP95wny6jaipGloIcthsIBpv2ss1kbYJr6pg086PJkimiFrwEV4PqLcNhyQlB
4IY0nEfRK00yzMhKdlRBPKJbOlnq7hZImuc0iM5SId6eutmJLuYtZ/eevK/es0K9
F/YobFUjfxZaH/t+dVVrtNqd4wJCv5lfXknj3LssQ471zN0yzOJw04K29dThyOg/
oHKrCwX0cx0DW9U2i5lTBmD1KPCHrVK0AN/3qs1I+wP3eR7OYz07Lh56HGaCFcaP
aqe9jlMS0qtJoaOgcIzPXXOK/uJRr2PTyU4q9Sn37Eb0PIpu6mb54hMR6EHEUzZf
jS3qwjcO1gz/dUTrwfzkG0q0wvu75BQ4JmxjMjW76RXzwQn9rWl1t4v7p/KQehhv
J/LqJRg5tULevvPxLsmC4MO1sO5O4prlDsOiBCxPs5L8jyjAIAs/xDk3CyFtdATc
7kCxf2W93O5HIZQyrm9y2nj6r5HUGl4YelcyGB2HTeYm2kV/MZYSxc3kaOHUmltS
nw56ByMNtXrT0RL8bTsxUHp3k5enTwt0QwUO1lNw+uSuqG08L5AYtjFi+CGI8sBE
exkgr+y/BU8TyMyalRH2/jjofAkgDs7yT1Ee3hCjnM8PhPsOykGBlv4hgtuMsNz2
990BwIh7C9XChGndtcRZcR55O3GDixXfNSd1c13bhYjYJv++8wT7IaVkbfk/hBUu
ZmrTDN7MiOWeFVT1ZQYDDV5N2tOK4NDckGNxElZtAoFdHJ9bR3LRwml+f4VfFJNX
Dz+EN7wase1JmF3ml58skg==
`protect END_PROTECTED
