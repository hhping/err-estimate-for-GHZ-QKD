`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s8zLK9FHPdOS+aVDPIr/PiL3/AmDr9EnBPKNa1fONuJsHZcldbV9ulQ1e5QsV7dZ
eeqDlKCmVvGRjbZyjvND+Hk8p6B/HzdPJUvMDx+e6voYPjHc0Hq9rYK2DdxGqiQM
hFz4bo02+i6v/i8FBtrJbJDDzyXg4wQEnlhayCHj1ozi3k4NP413xpQtno482jlW
3r3CQwwQW6pBwyUQahlpUeLNQ9CLquTWMrIpJ5zu3WWD2Ts8EZMV6s8zme7QTT3/
4XN4wd2QVQRy9QZp+zEEQZcayKRFzVNy6h2FmqKcq4sgBYxkDL0wJsUC7Tmp98bd
Yc5p7eaqJDyuP5gAgQpknRO1GCbD8DfMwAWm814d9rpT4MFzwZ3+FPJtbTB2r3xE
N8dpi7MWVbiiV3eUfoR5it87wV9dyV8S/PoowBuhMTfEOKKILHeA6a8lanYOz7sp
b2LyP7/UhPYUA1Y4Ucb8kNu2Wo8CWsDx/UPBUf0C2bul1uKnDRL4g57Uwvdw4uL1
ZaVBRFNU9huocEMWtOTDfK4Xkq/q5OIDO/i3bpL3NTXKcMVR3QCok8ytdhKqNiZJ
HUNFYndy6YcoA0N/+Gbo51esNq/HHeeMLq5Wk3C4n2qvgZ4zdv2jtgP0f8tWfT7i
A1qHxysYsO90FQna5/AR8IEREJaP5/VB+eaOZZH1w9BhixjDvSdb5YkleNiGM2Jb
0KtRXQPXM6cAixo/5QQXXYNNTK5NnkPepnNIbmsTtZLTIGGf+dwzn0hrAdJis+fR
r6Hq6uGoXnJshJKVWZYbaLcmPrqsirXPTllJzq7jscvyjKOIM2BPsQZuQ1Dfko8i
c8Zs+LsWr1vFVi0k2b0G98rUAfqf5qIYWqaIqicsKnd0sFrmXs5X/codvJk++AIV
RYaN1jcq8N1T5qlxGjr0qeHYMJ8Gr6TQsCvRpmzeaSQaRq5m1j2CBfqCYgm3VG4o
KMoGs54DUp4edlOeDe3+Go/JBdnhYc3kMas9e1T2EWP8kFGTxZEAUsjlPdcrcZOS
H0oHqip9cSdx0UBqvbeu/lN+QUEcelgYIHtfRzQfyhu89pwaTP8+DEvZllfjRSKO
`protect END_PROTECTED
