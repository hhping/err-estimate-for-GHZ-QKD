`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TqsfUKGWLRwfHv+hvfDBRpvYGjOOy+Hm+f0hvExfBkn6LTdckhO8y4XDYqgmqgjB
7d4PlDnn3/uZQBDBj+Q969fpUlhVsUohcywRw9OzIfnoy2v+PiINdcvNre8mDbIk
z7KXX/qyx44m4Gogjvp4BlDMfpwtb0gdHNzCVAXljZRk+7D49uMbCdJDbbM7Iy2V
SlKiZA8fNWxbYplop3JIPiR5mxVT6oAN0mFkALd511cpmZz6V0s3wjXcB3gYbN6E
X1OoJ7qxD3cSWlT6Hw19xKgomwkWNwRXge9sFPD/FvOWjXO0EKVRJi4FVU/pyTXA
G7tXvIsGBAFA0FmzUbkEXjdCAwck1b9RsgHmbDCekBIKm4D9mi5ipqwFdpbAgDqK
AFA9N7r6NanTO7a7D1g+nrY856vVblUU4dQhgApBCjJoIgBmMt3RWwZNanc3Urje
L5G1Rl0q+68F1UjJQeRKs3UaXfqxqSJm+LnI99GigRAJGlu5KhW+4Ba4K2EXYKnP
ayXANIVUuIRtApD9LBSe1Vt564scGSiQNbr/HtW2OtYK5DjEFdDar0oZPlzlJDQC
nK8C33Q5Ob1Fp4amz2rbwbnil3DS+NGrRQB0AKhi9mY9j8JCpaHUpODiQWq4G5dw
Ku80RGfHjPMUMClochEknq2V8emUe5pwU2x1FAIfl9ynKduG/HVfKI7Jq/TCvNBn
162jIa0pKNloPOkm5PopE4vYLkqRl2NzAaCOz6xBpx60nvjTk3IRkPnNi8AgFA/H
Spfi7Bpl1p/lGsoBSVWpL4fJl07rGG5XP3G27vHu3NWTad/iqK7Q1I6opDWXH+6M
ZcIa8qbGY7fFJ/sIv0/bxmyGmyz0Xcxja3sm9ohAUXY=
`protect END_PROTECTED
