`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
icKtqNmeZERBX68LOMGw2WW1MhhplWxTiMrnBwBIoF2wQ2OAaHkNQYphvUuJHZWJ
uN5E/fivwth9yiyvbAc7WjKIgDMqrDiWf0QxmEAs3kpTezwP+nDKuhL4LiJZaM8B
7YmK4n92FEq3iTuDGbNUM7hlkpbrGhzLLIyOEENYCYXYn+Z98i4v5dZd3f68KWU8
QvjguE/tp79xoQBuNkgEcqvwHxaCv773mDE+rJmkyL9C5DHjOUISmIkDv+X8nKoq
XarLZx+MfKgENIb7QfkpKMx85EREfpCaxv6pzX6WeXXkMNB9BHg+5jYG8VScnQr9
dhARiGRg3KyJ2CsuGe8n7XYESJieDlKAtjjztgnZYVE7UylTQO2hedk7wdZCMZHM
pE3Ky7L52ULzj19dfAk7LZV6ELrA59uh6QKWx+o8NdGLwrhtXuiR6P85OSCD39nH
6iX9kzl3/bqr1JcfsuhXSCedQqhO+kdYAYFYXjCtCMknn5CJwmW2YlMbtKq1tmHA
b9VavmZ9+qP435EnQSNID2THR8aJp3wBkjLx5To6PQUSAW2t7KueEzYLwFJTYDf0
Rnru2/P2ebr4UXgE0ns/GikliCZpDibzDn2KfgtXkrivEExXl2TfohNR00ae6njp
nsDko+9igQGuOys3FmF7ur9iGT71uxOqhZnygSjpwf0g/UKGFeYYgzMfaa4e0ug7
QXlqihW06T9jM2tJLkvUhgGRzxtZj3ug8Np0Wvvzf7ch8R/UtyYHpbljzx5FnQnv
80UWqLgPAFIfRCDq9JlOGmTIaX8oXfeqFp2BbKhhcaShsWsBbjtaMqdKLTmeewUS
kioJvbHVS+Ckum5Y6t95nzB1Yh5jMc2yMe8xlpDm+IoeguiQldNEiNvb8KL/4a+J
f6WUQTPzzGpHJEVybSUm8wwez0BhdFEWC6uo/dv1DtixP6aw6Mm1Fzj1ikTFtKxw
wpp2WjnSZt/+TY5AOnAtkgVwuVkb/u6/21oTnLZ6unWYN8V5x56QbunM6N8edpr8
fau3XsHM1WbLMkc1yuvtq+RL9so0ZwVMgwIqsdUJYyGI9sW+/9ZFEDBFx4iWZ3hS
gyTl3YvFe79RxAmbiMcTAD1w0HDakcyh2AP5fAuGKin07qGmgJsQg7hjjczB35bY
86UIV2MHC+FMqSmwqDJjwAeuHx7889F4FAYYKNTeimKHlPTHkeBC24JxqDlvrFBs
lSJPUgcQwGayL5JNAEurESNTZN9PkrcGBcznLQshjh7spyElqSQws+Juzmsxp4bv
7Uz60cLlXIT523p8InnnfJm1ikgFRlFbbgEKA6A8e4J7/8JU3jcKE2zmdesIB5A1
FDwGVy42CxjuemjQEUQUJWVrCsGeb/C1qYlVzpAZrqiYLO+9u1Wu1Ccm1uPkfAs/
BWE/M9HcZCmblU37w8CWZp66DiKYFWXdsjn2tXJWt+db6Zn5RDYVg4PIDQmPukXF
I1osMjtnz7/+zFHK0Bn8NGmbwmCzkzUo4BwGMhdTC0gjXqj7Qoe4rWYtzK8FOpUM
LvSnfOX6T19WAw/ZPiKXaYVg9ElviYK5m1M3oocs5F6zhrtaE8WxFKagEKi5nTWP
Yc2+FuTXpSFdDXKZmj/tcT5PqE2xKWf/Hn+PNAJl4E8C/Dm6FCpKbX3Sj8SZmmiD
yeHeRFEPSnfAckeALwJTjXbjBqtpQP7xUnhpmWBtPg3HNWdZlY7BSnKjwC6pP2BS
bLDdpHNI/5Xc6LnG1QdY2uuP7ERgNrfqj9m5otgh9lTwDL+7r6XsQ/M1Tun6rWg1
iUW3Lv0NREl7qLjbeHk6S90Nh0uWJFXakAh6IDbnJS2CIkeT5mVbVOWr4B3Q5IpO
E/OMaGx3nKfbE5zzXKgdF7uBG17e+JaKIeMKiPu+LKLaVuvmI2u488zBQqnDSQz8
8zL+3XQpC2Ve9iNt+NyT68AEZyspzL+HyX3fVrzd5jhvihaIvhjTKGK4U4GQrhNU
cHzcotcrwUwPDOdvsl1jTSQfJOLpKYEy10XU6pptKBivGochgBvoX82RiYjpXacC
MvaINh0r3zeXzahUKvDlA65Ekrrk1lxTaiqWSjVGIJp9pXsgda7Bc8IRnTJM/d2w
3S63+CEGCERACuHOOFyAEv91GRHyBrmR5PIbM86LCXp+sAiFBCNXAHolPkgsYYMx
SbmUyD6rCWtNnhO1pon72MtCsTblloPyHAAD4VVy1iy+IHJl/6EN8NadFKYEI6Po
zLfP183B+vbY1qF4UUc3IQnHquW1BxNN+vIpv/lsKOOdXxRm4FdzT9pymGE7SkZl
9fb8nRaL6g40GvuOSZhWBdNYKuujkLe2tnkIZx4dwN38GILXk72LGKQZaPGU4UMv
DVrBHhk0/dUI5irthYsBj7mcC4YHCqxPNGbgz7hyf4bA4CWTNAKUokZqkIoTBiJ3
w88u2FBpGLuJpyx7WkNWWnLFm13wFofzOOUW72bltrjMR2QVXZUc/ldWUFf7iWi0
XKkMCstVoOMGnvJjcK3QqNEwS99FzXMBkPyFl7vqWBUv7DUWWoH6Lgfldomu1mJ1
Gc0VDSAMvfRs+LMEkEwy/8rLhZAG2veqLAN/yzPBVUknRZ0axmuKBlkz7sKqLFYg
JgYXE2+Dp1N17J1sKuDP7/I21PkAsfWiko30WIl4DrB+ghiY70TbzMFkH5ZkssKP
6XYwBdBFJlEXqGU1FxHhxBcAEoXcNKdVkKSJ442O712Tda6KRU89cpkLL+1Sf9hs
iou9tfRXNrtNhw0yixvl+9mihZznuVr1CUDBVLG0LKdhaHZMoFXqyU8XX6x+w4E0
7PTDkG3KPnzy1VOA0nUGmorjaveywkZ5sAE22P8o50BRrYHw9N6+mWhhHk6dMBq9
guJ/9q2gakLQZT8jGV2B2Y0xvm1x3OBYis34O52yQrwWvzFndjgaMA53+f1wyHJr
SiplAZ8RvSyII1fVSb/IBPjeXOtoXfmAZQodVMCd7HF95BszgyF4iZQTMNDUz8oJ
5zZAAecYXCF+QHegnZWMnskgFHWuzGGq0QIRv4Ph34iLiCulAYp/BEtD6Oob+GS+
GFHtcePhRy3kdgFS106RxbUtf8jHWUgFV/fvE6noYPkVJJ2SpNJ/v34fisF+0Idk
G4DW/DTV6EjO1MkWHhfg2/Ai/mCKmHn07R+/56RvzUjn7nHNfulS7sZCLRwhm+hi
UpjDjozV+/4Ag31VwEmsAyWgzcj0RpEXsAJLnZPnouCY9Qzic7AVMt6v5/0kKXSP
I6l2ZllokbPDJ+5rmf5SyY+u4SSHmJzps2wW9333vqfxMTs/WjlIIppRhdBJZrQ9
IJ7UmrtTkiZTtfVtQtemNq5vS239xQLpJVMAfS3rKYiQTI7PgEAAHI4cM99LsTd1
DcgWwZn2Fp+LBfqQg4ZTWG3+f67ht0Igm4O8MK2TRVMmQRR4h3Jbmn5MvnwAO1N/
oeXvIDKg/H4mDUi6HutNWi07RnvnAyZsif3QmHXSEBafocU+MsukmdbpwBcRwt2i
WSLUZVd2Xt+Rmz6iGcU246vsjHKgJevPbizlL87Lm5NxLebJQco5Tj+L/+i8zYrt
0KMLZokb4jp6hrSwNu82BwO1IGuXN+TvHnx6DA6aoV2wwYey4d3r7fG0CPehYeSO
FY5ZFn76kx4WvR7xijRGOzJ3tMdkk2iEkKeS/90M0SVMpqk+78yp5WIKprP1sbam
iRywqZTOUP6X9j778Sm0+bkubjNX7Oyljf+cyPHmSkS7iN3ldOwN4jGYlMFcANay
1Ej02t9Yv7oxC2F07HhBJrF1EJq3x/6z1F+zYDxzkByxUPPMzfe8YuSz/ed0dSnZ
V3rk0DKFnt7/llagsQxuvEq0Ih6BuGQCpzeqbhzIeR8y0u1pnK5Kn2M3cEy5ehOf
AREc15yWvEFF2Za3B/LWFDHeFyYj2ygyLThaI2hgJMoq5FCR9s6abcS1qqVQuDzI
8rEzAN4rAuqf7QdIiZQSOve4lqBXiKk/Euczt5ZHQ5/SkW+7VLFO2LNn8TZod341
5j62BhKqgnolDGVuLbI+sozoAspwSomCEwrV1hzbBVuJKNWkzdJk62E9Mfp5nj1g
hbaQo9fwQWSiWw9hea+SfZrVUzb16Cyiav+5ZhL9fZMRY39cyp3I+SO7PcjkmgrS
x9LmVngp5fTpAcvYJwyzFrH/7uWGk+QdzMYKFcXnWSaiMGJBWZJ9tOZzUEzbSVmI
vliZrkcBi8J/Bluvv0EtIpgzgPveTCk2d7O3axFx/SCX2fDwbKWEzrwccaVXM0kS
SHE7Bszyi/uCkoYuZSWLUqH68U8CLv8J8QiT73PXS+UAIsLA6Jv6c6Mo+IQ5krEA
oP+WHHfhlGFegIpfET7Tpjg6XLjOpYzV+a8ykgv7ljMht9sYvrvmWjqWl3kTz5TR
2dsE8wdGemrwE0xw6tdMoMuWhDWQ4sSvamjeHIn3ueG5XrvkIpG3nYUgYCxy8Avt
o6unNHFkxKI1Z2CZFfYRRoN5d55olqeOcrcxNk/vHsC9a6oTivFjLhCZVdTA6C+0
sdnaBnYphU6/lxq7f0e3umtElS20bfpq8/9dR26gamSe4EtWvETlVc3c+aT/lW2n
8oQvEOFMbrFF8uU+dKEowmF1OzN0frmAYYzydpdZFJdP5ZgKnm9iHaC6lBRIV1X5
JEWS6rsl0iw4fB3oUVw8+xp+zsMDOYvOUqBwoNb8DOnxkMxo9pgO0vz+mLelGgE1
x2BizVzJn4TnVaibi3sVqjXTp/5aX+chQCZ9nCDnKWmmxCFRIllnmOuMYPBtPZvX
An2SJqDfhPE2aC8m2ZH8CYlaDwKXlQTT1/3wVTePzZJljD5io+k4mA0t4WnoWU5d
fJtzETaXPLOmXAmOkdRgQ8WDAe1HWAaM1Ab58UuMxzzYZGHbgcbtN3pB37f/CCxQ
EfqlISTTsEnEdWOXJqz//mtS17DTeWgD0bFxS4UPJfrQ7tQ5L8XzqfQHNd/r0e6X
xT58CEggvXb76IrQoJdunPHK0Py3iZVsRYdq7/NAvQQmz0KlBCXXnVbH5qBuAXHh
pCg44uIikah45KwV8fSMQ/7YlCm5NK/YuA3a3oCMG5+wjOsLIW83noUisrir6NSf
m7z1GOFAaWurMc2M8nqCOoGfClBXtT3fn/5pFl7Cx7DL8kCCU/NuarksDRJdFTXi
//bz7J2mOv66+xl42yYPDtOl+UUPVkL0bAo7mNe4EbTexQPzjJM2fLBYz+WW0GsT
dQtkf4I8lEkeoKK9Zvr2JCafzfVf5B8FO89QKct9YgkgPfh5yxAT2gcBB8WatClu
IaPJ5p6EAcFpTDmnWs2aOuHm3lD+PcAixz4EDPtRVwelFPGVXdPav7mYRoms4LLS
mP4xKaMeTr4/Z8aDs5a2kUyz4vne5sbP4mIPeJZ14Fi1JYJdGf+P0mxXDbOd75ac
PUVYd2+Sji0ykrcwH/ilSjxH+JXbXV2n3vCb6aohx0fNLyX5SgYX69kE3FBCU0jU
g2tuqM+QxjO+E6k0jk14h3IOwN1XvG2GRLDW5k86YvvcBGU/R7uUlCiqVn7OPvGI
uThvrB2C1+0fUYl/CmOnpvqGdQdmpc0jpBw/r70ULLLH4xrN4ooIFAC7KH4SGND5
KfnK3Kfb5srzHTl2xBL2EylLbTT1PbjDQ5OaHBBHG7vVOuisY5nU2qg3LgUFv11+
HoXRWFa/0/aZhcWY5C0jNXI7Ff2bQBr8sWxQsbhTsPcF3fie7y22Cnj2k6d8EKV5
vErHHmjAIkgNB9YPkH0EMwUWJNN5w7vpJ1t2n2IkTj1yfvFzZFqUCg4dQQVvHnW5
2BEFL735JkZYzQKU7UrycCFQ7WZiUwUAHHngfgDPWcgrVVML5fpf/5ghYO68JrxI
YkpES10wwZXntu/08iyBqs2zNpT+HvUR3QBuAY/yfR/6/2mxR58AkpcfdLN5OmCz
hUh8xPUi11llHCSzaiucSShCfAl/VF/GAILfEXWFm8jHlqGzTpMN1MiVKyzhu9ng
sRurrwIj7szgEbwVAogdzXmv2hDYeFZ58UpiTm9GtzEylppl6ZuDoyZoXSdx4lnV
+E5HWygjDTL/Ed74DQZpGevCanaw+EKSRghKeTPL/DAI3dxDbPTuLTD4mpdH1aKt
nwgq9cHUDD55SurpffYxON9Qd5rhXz9pPcbRkHLcA96qimB/eM2+iPUFFP6nhoiv
TB6SzvdeOc3vZe7hVBb/Pr87/CPe0aTR41erfZGrqCcQ1OdQHzOdeqwUMyz63z5c
umwr1heaFyLVsva1FDk+pUUP8ODbbQf2v9T537H/KKZ35nEt1xYypZhLusWB42R7
7ViDxJ4PJ0V9a0feDUZBo1ijXqwKWc3okEP7hneNtA0SpgEBDy9ygpMBcNKsB/yz
WncEXiiSGoipIR3+vMiL+1L9yLebeCznwKIo8uTrNhrj1nCAdcWEj9pupshCJWni
Z0JInUSj7T90xiuir0Nwrevja4eBv3vCij417Bw0aYCdMTc9FYxRZUqU7xAZXeyW
GDB53kyYrvkUuCjVXLH1BDa1fpep7HVdl57TuwegqsB69lD+iPWp9+f4HSVGIlxg
SN1YGeUN2SIH4IZO8jUK8xWX75YiurFPOS/9+4mw/8XM3V3sKm2o1MPjhhXN40Lq
+K+gbChsSrAZuB5u0WIw3ahDLKMccL2Iik4KUA7qQskXmsTtXDSjNFwVkGJ7KNCG
8qFJNl1lw0poPfxp2aCMZKsbi4gtCfaafyNcdU+bkgbh9Gy0wddyoQlHOzt4sac4
crZes2cd+sum5Z6DgEJUeg+lqt65R1B+xUMtOhVdlD9PumcANoOF7c6URs0yCDOR
+0n8ihqjRQnoVWOrn/1nVC7PQa6zgQ3R7R9G/qkX8fW20XlQvJQBDcd6Ys+dxd2B
Ytyfuo9teu0rLXxYyHcz6ax9661/ZM1XyLdGwbiYdD6pSaqQx4bqxr6B6sY+j51L
AGgNnCCPYduVuR6fKPRS2WlHzGCC8j+cbIOB245YAG1aVjG5r/VDIABJ2vBpk8GJ
PVqef1B6fiVAcna1iVkFR0nXoJAaYbhSLGfDet7SFc9/zqUzXkQsC0RofVjzRh0V
TI1M6vx9pD6nruisrsRuA2EqxXPSrCl3piRY1FhGVFPK9S+IqKqtvt2xm34k50pk
eQSeuUEn6yFXeDSgVNzJ25SR95cK7Z4iOxsSUQnfnHl8+ZWyx0vqTHwHZfEWNX23
RlkduHW5FIIv/FN1S2o/03SeOjLeR0WB174kp4dMsdZ7lk4G3pgpsPzbRaMw6Els
2D6bAJJfMN3fGoUtmzq4rI9nt5dipkWKlWcNI7MQ4rykaDnV8KPesr3kHosEpyrd
WE0/1qBZn+i+2RbJUc2PdcYIPcqWIKar2cjn3Z6d/mtWH+WVW1jHygb8g6a0ZLFq
xehiQtGhOFAtM3NMUHYcZy05+gOrWqkR5cQ7cVhd/VsKcvhjlJHj23kf4iZUS5af
7I386E7xJOGKklzgzlQLh1XWmiTiTIT2KjM5fZPyuEUyuyCzOJ83wgVIAcjj4HET
w595nZlL/KHSAu7MlOOSyFFASZ6glOQfq3qJbI+ZW4ScQDoP9Do+hODXkMDzI5lB
nPqGLDX4tQ205q0nlLOGIn9kCsm0ZPMfG/zhPjOu7lS2rocXufbos4/NCVbSxanZ
MD38eu2LkyKtlxG1lvF1BVl6LluakQZ0HQsjZZRApG9xItE/E+oKMswQ3RFuTnEY
JsQFS9JiIGlTp92e1e6XaXNcgQafS3lnK/E1RGL36DOYh7vvT6L4DDYdugf9LbN6
ggk7pM6iaEW1t5x3j4y+q2uQnk35hPjpcYt1syjL5h7ra9RQu9fJojYdKQc+/R4M
hThjYwzMvNbl01o85ehkIIotxtjbNunMOOjTU+oUS9nZfYxubyCba7qVLuCJLftk
J5eKnmadrvxJoIWsRgQmDMeGv5GIE4ygZ0zR+wGB5TgLv+jA4c6fBSlP/X4Gccfn
NXpR77O5FLRIcSHf6/JXSJeXif9q8GcBBW3EkxiEMtvwbAry3fbVAoRaBn/9xj37
jlhB0qt68DUxk7WzqS0wy5Q8HQzU2BakEypWaDO/koP4mLYvaG885o4IFv01cie1
lmRqaWXniVSp/nWoB1HggQyF0mefEfnYrz5TUtWrRL/zN0mx0e5FhJ0E9OIAGn+Q
cwM51oAkhs++wlQt6mUKelg68HD51r29gMb788UI4Q/TZzOWNXDCcXz2dy9ITA0j
Vbl/N2NqaDHaEtwZcx7G0ZM5yR4G+bSvIySJY6ZlxsFZw+opZq+Ute9PJt9+zXBY
P6cSzK/uJ5Yb1fC0JxuecvuibF+CMYvtsLv5nUtq0hpk9Ch/xroqi70YO84DJHGg
fLIgMdcNsir17Gcfwbc9hIYfD5V78rPz4ntowsjNua+WXAhIMExJC38GzhiG7lpn
cn5GEWunoshSlkXOrmEVm1XBDLIPYKZqPAGOafatvguyoPXUzpwrUSOpRhwRDOhB
LdMzSpiEBdOhK9K9CG8Kh8flj39ik/fi/4/of4oBkabeFSuKDJfJ933B8H8925CH
3VQhgCmEksrA2v8JD4gXf9GX41v2Dl6+BwnA2eXD0kbMlJiu5oP9f00ehpL59AD7
9vC2j6r4lwMztM1iJ1b1rweLFTZKW8cHR9A5jO/DLWiI9yTXAvOTdI0DH3l6aRnO
rp9c3dw2CZS4u4xphy17QPspVGqCgHwV6afsgBGTagaliMEONK138GA/2yWuP7NF
AVlUYusesFd2v2B8E8LC4shwlvZWIyRHJABajNFSL+ZsjzGmMmA778MmOaFIJclN
dljxv4xkawGEZTf7o7Uvo1+de2BZQ4oprXs6ODd1BWP6CLPd6gi3gJQjdhdplFMx
aGuUmwZwWsmpnPD9XOMh4GWzSJ8RD3oqkwTBwuLX1UGBTZIcFCx4TwzJDTmU+my3
vaKqcBmdRAr3hEVSmtTo0brXVxRzgxS/g0xBK2c7QM4T2kYoV3NurUXRyoN4N+gO
goWtomEfYW0bXX0RImjRc47fSdNWC5B4XiYhz1gIJXCvhBSKJSvSECItYtRfzdVH
TYThF2ee2cLk7GGoVkGDIs7422IQVVlo952xxSZy+1RdfxXqzkV4NfI1WyMKHQaq
zz03sojRBvOLhMDV8lhT8uv7Jyo1IaQ9YwyWrsSoY5a3kQP+bH20s8+ZSCpQXSH3
k56eQdiPjsowQ7tlCcNo7kaB5GkjjB5CWfHnQfE/U8Gjo11vcuTAkAWE8cQwCbLQ
Yr4u9Gr+pSCWQ5sooSle0iVBTytvlgUAVVFUhvxh9qNJ7iJBBlwkuisfIFgv5oZe
JuwWUOdSH2x/WscjMXL2YV4xyzU2eC+WFaUSoWuxqitsqwzJrqL+dQm0Ozf2KBJl
6TVV6kERn89hRhIUyfdp+h1HiQx7C2oKLQK+p8v7G1G/htX9SrFXS5Ulql2IgaD5
vkVaJF/gRXmo/cyAivkJczjhLqjuri7DYgIIKXNqq57elIZ+yzfRf1uwLD4Re3oe
panOOykyOOYaXD45q5ghPP+au8ILQWlP8IMOIxVGU4nDCtT9qRtslndgSbnJiM98
6qCfx5aCZhUcHumW8kivlibymVWSjEh4m9i/FP7onlWzZH3sDrEFsqttH52sAhFG
MXuy7d7O+oQhpasE2DQr3lA8IkhX04iM5KnwwYjPgxb2Gv9SbZ9+39xtJGS7ZOiU
8hM7ihf9M+mW8KWCluJFZw8aU4L2fEl2IAqRksB34MugQhbTN7UBilb0RHBn9o7P
OnZug8C/W/MUP06wef6WxoHJ9+d3C0ciWOjk7lF7VPYyFiXGAacfPrefAgruXhiz
VKMrPdfsD/NlJ6sl5YnY7TAhbxInbSdqM53AmOxFShldPgN6URUNZIEgf6XJFuUh
gyWVWRaBWqmWtEmJsaKsjhNwMtMG1A+c8f9ROG6UlIhbFB86p7q3wnj38KQO8szH
NHbeCCURkAsrW93lU9j5PKoY/CMhjST/RJMUQT1lzXKjyE0bQJaO/HTOmvo1js41
IIiWT4qs5hkBaLvBUUjHsZ3o6rKdir8y4DRS33d35gE3uThmfhLn6MuELhfkCkFx
B7N3pg988nodoDKUuSATDk/Slyb3rl6L+uk65Qbwpp6VOOMlmknIDdM3fFkZ+auw
xIMa1qiNRAdCbQ1NzvntWlTTUd+HWhqPrwXaSwEf/EgfYYBwGW9S3u6oFJRc2c9q
KuKW3w/Oc8MmK+ILN6NfYXXQJpLzGzf4s4IF5oDvkgGca9apbMkXXATnHTQQiMy0
dli/QNkbQTTY98b1PAzlszkQWoMIKF/9UX7tqxoE3/rRvk0m0cxlm4RH6E+XMwt4
1zo0QAgn0+S7gHkTwPr6xr3B/ysEEcolj1hwaCCcO5TN1KSHh9Z561TWPAD2u4XL
zTs3iAElqpRpERkDYZevb7isLcP5wa+fM39iydFmqVZ55x6ENe2U71ts2OmyDkBJ
NbrmQi25Lq9SpgkCY207nL+q+RFSP0pUMfcfXFU69oYWeNFKCALSuwTfkFyQ+dXv
LTBNoeAU60S+8saWOeS1me/c6hKZ6W8YXFhEDuATEWS9h8KGodwLoEmWGVtTMjYl
hWlYwVMYg5L4VhwlRIcVnFEGVC0YqVx12mFNuXqtSdNjGjDtNx4X/7qTaMvmeJNP
3P6Itjk4Q9CoEvgk5/5/2Iu1EqeQRV47XEi9bCd3zT7ESzgUCEBHhf0dz3LgIaTd
hwLaoGiYUUz7hymxhPZg5Y7NeV4k+LsCYjLcb9CHt50+MWQruLqpGDWIBYyKxfqG
71idgpPheJibGi4mAswx00iqR4H0KF+XiXEozolDVwED3zsQXNBHDJ98ogYd3MOu
RXXRe+vNSBXiTrXGQetJPQ4/9gu3I0cZPTpSMkGq1Fl4r+DnF1lbFlyz4MArsGoj
WwHy1SexhXo+6GuFPCMHrbImi//ykN+lV+WFmSPQ7TMRB+kvCuqZz3xQRbwJMnNm
9agrh6oy6pggn1BfQNkEt3Z2WlIqLq5xqb2aLbOQC76rOx9jky4Yp7ap+59J2LLv
kdK+lRpKSP0jaQ3UN+FSRMuXe1lo2zf/SnkCp/ArV0TQOzwz251M0D7Uqld+0mQw
doYedvorwudRKCo//IlutAp49GyeapdWRwqUVXW4d9Gzx9cqtZQxxM3JVpbacKBg
5Z5drhPAB2EgGYbkH0JrIbSRI/ny1qNSCzRHAzWyO2z52IDH7GJ5BHhpBAbt1iCP
xXTw+kUEOWQe1zzAUaxPt6iUBOld3zWDFwaPvhh2ixc3BOLwihe41eqEYJfnWShN
NOm9TgTm7ayg8W4U0q1GvLSbzIEe334zQ1Nx6iGz4yco7mOYp2xL7PMvb2vwJDBS
uOMAJ98MfiFra9ujkOJ6Fqmn6tHGtRsaiIm5CLYN1gMmAhKlMPq6/wn7QvU/mTTy
6fwJNaRWVc1uUwYpx4CFkvn894oD/7gHvWKTN6tAcVHAMI5n3P0QNDxKjVgpdR5y
CCOMjOtwZydSj2L20R4lY4TYVq1KCGX5qV6622Kz4/47c2jESCHnZma0uAW+2DSc
QyMCzrnwlyvDDqYTqd4Unw2pIU5VtP1+aoXQiqlFFsELV7Vet8JRoGhJgJH73XAE
533Z3DLN5aoaMQXdolPE4u6kdUnczKyhYdjo8auYbk3fhBN+BVHoei08K2hYkPor
xRnAwzcVmCX0CSwa3F6bVilqGXWzj/9VcbE4/URU+C7TZ6ptR5maEmZeLjMXKHcQ
TxhG9aogU/B10r9mKecsra3LK3oWGS8yPv5xd9HVCioyEl3lt40dyHjzNgS6JI04
TdMM7ZbDBBuOfsyepBcAb9vQnV8buo8maJymKYG7zxac9YkEGTB2ijJZPQpE5hSF
FME4lqfvNkTIKFQMXCcYIleQfcwtFoMpuNzn+7D5Tjxezp/XNXjRfvhZ0+QbzGGw
vIzqLuMfhaA5pCO4izIMm1hJTOR9p6rWI+w30TOxbnEDy8kVERwfRBRMwhcHBsUg
MtGCP3IuQN5+gc3CzLydtrLS4bqvef2rBtYy4MzkfROUIxVrLgTCrc1AGmtMep/p
uM+Mc/WnDOIsiZsA92UZTBdYi09ChGtSLy/U5qOPf2sCmdeTmvPPJs06V4selzGM
r/PZVrP/qTUNOIs+gRWWIe5Vz+36UaknXfZQVfh4bJGkMEhK/FXxAVOd41et1G+Z
WUdRp/62rYd3SYz7yFTiBhEM/WDOrvjOmkkpUCxfh2vI0MOjVi/j38XoPIJqZJez
8VnHXYFh3VHHg2/jGp809Bxco5WKDDzbykOSp8xP4ejrJi/9cJxs5H5W7CvwKr8Q
NsQG6oXnK6fxdOoV1OZVbD1XJa9g9gpAGIaXfV6PdTv6kHmPyHlwjEUPHzXjAchk
ekfp7o5nA9Tf6xrMhd3nJf+U9oy4BZtgFDD17p8yv/VNS8i6yw+n8m5XgnKWdv4T
xXcDlaGmxejadx4LycPDQhSRx9+Rf5ZIMqj1ffjjNldItPA48ciQXEQ3ULsf7ZSq
bZAORxgbIW49+z2lxGa8i0Ddhkjxel3vZc5y9i3P1uiU5YxsA7M9XnCioZknZwzz
+ytzxqLbJ2oVEG+2Wwtdc+g2Pg1auBkXYqAabFtGbNyJ06kXR+jNTym6RDfb0uY3
LLVyKTfMci5fNBkbSwqiMgbKiqTEvF2dUZqf5Vf8gxjCK7J5ciilxUjMomeyHlCb
TkbLPSwo9mC/R3ghLkjVrHRFkTmAP2vm6Q99D/8GUckiUT2ulVbSUGxqtjGztpGP
hCT479TLkIwHkPdJYOYGfGvx40B7it/6/7cG4SsvTFZOpSIYRFzYRixBtapkcpT+
piiw+Qsbqd9I1ZeYd/NrS5NgM+aNi1mCbC/e/OAqK8+EcdyeJTowcL6YgZJq4jTA
Qx58utkLJi/OXWLsyXyZiVMCAUsyrFYSJ1V8g6RCqNcmDYlBXoezpPXetit6yZG6
Q2iwzqU8eIbrcBhjFLcCS/WvQYbfhocapozs9kJPN5YY56SMHrYLaPAckwAW+mCI
+DvQHNAdEvu2pf5Kijx7DuaUpu7ECmQTMBdVUt38FBgqPOSanhDreDTQfm2jJp/j
qTx4u9YEnNZopnM+gAFN+Jw0syYW2knkyuphyS6XpT09sBEulIUBEF6vdtApGZH/
U6L9Ai8qy65z6EeQ48Q4KYoxVgBileSSpUVm9PWEBFAJQit0QZInsSm9grxWz452
QLu2oncCQJX/26vc7vUMfhPvAFzs40Xby1nN8nI+0MIzrCiEFifg9GVLfg+oSuyD
Gb6h7yb2mIgwyqNxrhhwvN2+VmswNYYC0IjvGkHISIceqXhxmywecFly12pEcggM
JF3R3eHj3wKwL+iYNOGndNuduyEk0WwWsl8LhTM823WXYRU6WlAXj/IsWEcek7dY
keMyiHvC+0ailnk8Ze4DBTiwnGKnpjXjgFjrW1/+44+ooYR2Z2imvbvRkl7xxWH3
rZdGLHCER+S7i9pVZwbGPLH4jA8btlRi/pKI33teBt0hYdDTAPHAunA00m+xMAvw
uaaPKeH21sbQ6orWD3Oi5uLFyOoDczpnQvoQHK0yIMijn5rNdJHEAJ89SJfKlroo
9+pE43v1dH0E3fRyVUCFg8SId+sgmZw7HiuCr5dhB0KkHBRLGqM/EyNU4y8M9KG6
OK+kjNysVTYg4VI83+ZMx4nmXQ+Fb0iS30r6BqQLGz3+li85spu72lUu2PR6GLfK
oQIiGBIRUGBNEYsYH+ay9z29qmpaJgkfbI5S8+D+9xYGVAKYiw/VwVw4P9IPsJ89
XfvVnQ74v0UCoZvdNDC8k///lYHjP8mvR21GsT4z8pU+cz0869QHD+gtb/wc3WgG
Sb1XFJNnkcg7OZgGxd0MSCLhVqXg+x1qwO30u0acJ92ycQNt1tIPYojOV19C/ytR
yPm/gIxh48452k3XRK+ief4Bt4aRr64QMTJFQ3bE+/trmGq4Gd6NH7VaDEvo1NXN
P2dg/+ilSbplWvNwpNzGoW35Ve5jgnPQtqA0g3oK2yNg2YFgeyu7EZlYhugnXW6m
1B+JdddsKpNy/iqQBra4VLFFdpcR3hIE/Q58i8GRPohrfL7sQ4O7mnzPfZ4Qxj0F
jM8sl2Dj1SqDsqsT5Q8Xs+bMwGxVkcHJtRsn44JuVgPuyWCMbM4O4gXS+aDPBJit
60hZFqMehzyhKqLf/4UhtBucmdUBzvUPI+75STJUD2yPiwCBRlWSV9Ei5zFG3ieD
CSA6eGeTdDkPRvnuCIGbqvGvzHX75Ac1y/oImO04xLXSbmVRiJFclJ0T1OfnI1NO
9z41tmmLpPyNtHaMpnYmPtg4thKsidkl8W3d6ljFo1RKXyoeHJGZStRPRi9+uvTm
wv1obICw8S8kbFMYg3YZScBVLouiHwzCP8B/Yit16OPCDyqOgzt1OxuwXZKN7zAD
Yhs4f7orW5e5d0GYQtPrEshBOvZGW9OJ1QiNY16GR7l+FM7x1XQhRu7G8akVqoXx
6YrI71jEoeh3Nscolo+aBo0F0scBwvSexwbG7cgX10dRrEsBSc7AS2Ha+BZMy2Dn
lPEkK/GMlI46ecfbD0o0ZJpAWAIiKk4yRL6qJTyfAlxDBYRsRxAAt80Z3UAbx0b6
sSWuO3hbAgtYQ5MCBTGvnrEd4DAev31A4k2DYbbrStErMWJ2Nc1IL2E6KjVNY1q5
pKgC0B+DTo3iADGMA+KM0txgG6DbqJNIE4ocZX8fXFpt/JHcgp2CiuOuEPZi8Nps
hAMwW+9bfOzSe4w+vOe+EG5Qizw7o2ySk9/RQhWDfIUu9DT96aaoXAw08yTQt0F1
YXQfQQXcReZcIQ0PgG0pepLgcrD3YP5Ih1LumMpQJOrdoC8r9XtE2unE2IeSoEsH
/5n6xMpx6wvWBJwRPoWdKAW65GwpCPBUWXqdXzehQzDiXqbWKiddP0OwiFCN+uhX
7Rwoyxif2TYlB5R8+DgQO8/ov01YILyas+ah4wtQtDxM2OQcIyHbkp0eaG8j/Rrw
lHqe65zQ/Kq82KJn/Troe/A/aLFYlotFrL2RQkRcmbSpHbRw9BU3celtGIuctS8X
5IyaI/OFtNzh/l3DssEau5LNR23ogP+XRJVanMw+2Eggpe7Ot8plMrLkk823gzxk
pD4sEMYv4gD2sC3isiFLQzSKaYcwvsult6nxqUZ1L00eZrAnC04xe2tVxuo766C6
RhQda6xaE7EG/rRarrPDzEflU5Xd7cox8u2V67YjKlpmSJT749i7cGvksGN8g3+8
F2aSwKyitweWKEzqcfBWWo4mzwytGyuj7GPOf8w0eqcP7pz/OBIQs3UMz75CoXqh
Ss9+0DCjcJzTqer8OenvLpkCxezJ473oKQw4CxqlkSUApzRv0HRVg+Sz8nSJul0q
nalJ1/OmX7gprgtrEXjqEgaT/eiLlImbxmQ5dtXi0VOzetguxc1KMwkKOqdi70kK
tFktkTHaARkHBL4eOsfmaJ8CessxhOzWtIG8EO9ZahS/HWhKbDlcUElQfbOkf2am
WfTxB2d+0IPIdvMkfGqLjyD96NdmZm7KaWpaqN9nAVZK04RydedI1Pf+2ldvh1z8
dfRwpRkjXMtVojnBQW/Be8PXBZ5L0DgCbGDYEnMdSh5aptX7wI4AfR4ZDRCmM3ph
tuFbpsl0v4U70vp3pKL8IWTJA/wXpYSlRV693rAxCF9o49EgFRjZa6u9tsdEBAOQ
A4lBxP1UBLvsEWVJiEjWYoTEBniap9bYQq46WFvUg3wlZB9sL1h1VdVW+urxkNlc
l8lYZ5DTxy9enbtebfMt3t8XSHQ6VwOShCjwS0vqDuJg5W58JsnecYjxoTSKS4LZ
cmaXLMxdRwkMGDwMl96rHgFEplLAw9uzVI/dnhlDMdiqQX153de9dgHVpsL5vf1y
JvHMGH6c8tghmQo5gE7aKgHg7xHGhThtpxljT3ho7UWTKoIcikBbP9dH5TgEJCRw
rOL1ENP2T866+DE9+7XCTXOy16FnkdoxZyvi15Zu8med2a0gEHHAUDeboKUmtMlH
vndZlsSUvxj5Rls6unKA+2CtPjUL7tC/mbwk9IEOegbPk2v1pne820+xOp2F/vfR
dysIBw7h3ZmGskObLbKbPOjt1cxNQG1xvOZ0gfQL4iEW+S7XWook6kYdCySFIROg
ZMfKytqbAKI8Cz/nYsrU68vqaOEGbT4uoyNHiWI/NZdf8TTHziBpXDMBMVdmd0Du
ppN8gZXZ6ZwELnI58N9/TqAiOvJO3osAzTtE5qHRSJkAAQDbKs/mRu1leKvk/jvZ
v2OcjLgfGKAj7YNe2euFokPynDa3gzjb8lrQK33q8d1gJSd7ELnl2VbL4OxIUcF8
3Te+ispkwW7K98ag8OfLP1ph6dEcV8+OP/Mk9OGu/AcSeyo3SAnVFkJrRmYK/3pM
jmPb3z6uJ0+HH/i7qWgJO2q4Myf/ructWRftWit7FSpU4xsFVwZ2A9fejcIi0zgG
fDfeQ+Df88oZygP3LMRvnUNwvAsIcZwoMxXOYf3G54Nn0lihWvclRtxRcQky/GyS
xceb+EJfF9//dwjUDzuwvl5V/D5GznIMzhMm3yGazTvV+aoXLSaISE10xDI7yU+E
X6UUGNl8dHBxqaKr3AlC+degraOhObWzhZonAqg0zhr4TYwhjM/D5EUoSKcX30y5
OC6vY7pcHJWfKcm1AaLXEt2s5+ghhywqNgU66882ORv8DdUdZZ8pG3Ht9aER6vpA
AaA0Kt9HdkGS9reMllfWWyEjb0eatT6X9dF/UHPu8g7GDYOC/SovkmLa7/GlO7cZ
hvd2j8MzVxHoGfoMwa4VQVZvCiGwBLHQOO1Tx1IOgVCXecrs6TGSXhDzR1eblsRR
yZa3PlHZyNRYF+tAPhcBjdUA/lP3UUQ4YqwpApwdAtE0eRmNo+mGG9wrhrWdW9P9
o2xds9L6sEuLL2MZcu0N54J703Ffy8TWeR4Jv2gs1SbZZZ+cD9guNRRSjgROv8ap
7uR0YUx/nrebnBmgjsrQDk094Wr136Z2pcSLTO+Gj+GZbqPvBHOaQXFye9F9VFFH
G7W0HFwlUTVJHygXWTv7PSYrtxmCR94n1F/XNEENDzJ/Y1Dlck7UVH1iw5H0B/LR
HjY0j0M7IwiiX3jce7SEtifwjHCBkutnlyVSsuFt8dXVuD0sKtBuVO9DdHZvquHj
QvTeMNQAQolwn5ZfLoq25IWm5NYvC9dPktjoR0h2pZJihQ+d7+lAnHkjdwDPbQS/
3G7CVl8NW5+GmsiT/HUg0chosfGI5l+zRg4II5D2mK3Bcr8qZiDhgYGYIGegvv/2
OZf/+MoXKZmNP2RlCIHhYyFyyQb5vJC6QesgjeXiw2Z3ECg6yYLzNLF3CjeFI2dD
5xTd/ig/bbaSG8n9iUHdo2kHSZuF3LQhK9PHvodvn1Pl8r+Yy1efVgi3Xpf8SfsZ
KfDNZOlld7/gtuskXjCancAWhRbq5tn6irppr+zTgEGmfA8h3SlictFgzvBMfxBP
KOxOj3p2uC9a03efX7RhmEDLKy5ZYx0Z8trToF7p9DzaxCbO4C8fbe9z4IzCzWfj
jje/z8JTgcpHEXsdOJ+tHNYgWw+463mWjHdQ9OcuMvP8QfgRrDhz1ljBPg9XZbKB
HOFuQUF6H9DxN0gU1czQ01cX2xraGxD3sjc7AocJg6rV4CTFeQmQX1gBb/jhfaq1
jgxNp8CNeHtbpv3X0nFP38bQ+lD77zKo21tQp76BdEuK4ODoiRVDPWPXWRNLQ39a
xb4KpKo/G/Vw/D5zD8vHq48ZVX0Iy0TR/cKjaJ9NpqXQyLYk1CWZRNjhgdlIzF0N
c1CVjaN8hsPzzKfsmlRkZ3fzLSC+Goj3WUBZk7ysgro5zaOAEfMivFmUHsjSDjq5
Xn7wD7wy3XCqsF1Y7/H+xf9XC0d7J4PmpFNchpubF1b1gpPVwcobKYREOw3FdheN
QuME3xY6KtsRTMF+b+sIQsWYgRudu0FguLh40VY8ZXPbAzUGSxvqLpr+YQSAgzO5
dUttGckG6ruDKdpMistIK8DttGnhYfVG395vocImxjBr+kE++K9vQwP79PsrqMjb
l9nOtyJSxt0DAaAi0hNzd6Wnlc+vrMIy2lg5XqpmK1TxAQpK7aIjUSe5CIddy4WO
ioCmizX58H0cfwRY1kEmBuZINIekgBcKjN2/bLp5ZhVYtz0vTtuI9mCJsxVVyDow
wk+msxgvLZg71jyqpxp1MrPUNhzgSoQOszqdeb4ATfS23YlTjzwVfqGNF46gdIxC
znH44qf42zRocPJT86bUEXIPlok90IKosf/YdEU7tYEJk8L7Kj4KJuLVgOpZJSSD
HusRngM6PtIgVIAAUbEH+f4ZE8RlU//ao+w1S4/6vdsq5OE9uArFq5zboILToisg
OnOgQY1kuP6bW5M6wP+od8oYEXVRmIHfSQPQZ5DweAwT/PBc0Y3r1JTXP0s277h5
fXecUEBS3ciH8H+VG75Hz/YaUDNhfejh9BmWi5E1nfkqiJXaGFjua0IQ5AHdE9Vw
5lpv7lJ+U5uNpJqsO1uP6+wN/G4obq2A3fu8wpByPj84/Oryu9LRH6sR3SVQzaD0
yuDltxYU+v+KVSsyvoCNY2L+z4uyFsTZX+lHAn6O0bsCMxpd1WI5QO884EHI7lpV
I/wqNNTukvzY1m/wTgNkQv8Nmc18kgq6CJa6F/bodlwF42Q596TsnVd+FIq8kVU0
gZ34tLIlJoGIrfRM4cGbG4vCXgV63n0DtGG9g6yMMreSPPhfD3VK9yiXdl05/8lx
BxSBsKizLIytLYeok1JeYFbgSqW/LFo0vXMimQRznI6/GP4AYHiZHSaHAWQTqfQO
hEZpcU+3MgNEwJHY5ZR2TyFc71XjQ2RankkL5nFS82K8NR/Ya+4FbzP8Zj1CUh/J
jwb1oShzE3G5EihVNBtiXvna6buZk3Vn9LL9qhzxU97g4DsIzcgi7dOHK11M4JYj
zAf2IcoZPq5z/wz7w4kVaSQn3W4vrxzrthPBxGH7nYMXvC8yE/2RFptvEfahXPzs
QEj2JXyZGXwnXILcrDzxizeQC/ld00U3g2ws8jjw4PCacdjoaEFlyN6DOOxymPXM
JL+GELkGxzVVgClHHlJH/aR2Lh1hw+MDzL5rn+UOffdOpmR8DW/tX77fYWXyYbmW
b1yQPJeZIfVK3lW7R+QZS51AejR2nzIkftBe6dJwBBfg9qp0mWUb8mngOnwfW9J3
SWKg0M9wd/Brqzgj/ksPKPSRI7ZU3kydP1jJ84BYKx9G22tzGs9qfHd649hwTi8G
ggBYUxDK3vkz+GIzdyl8B10QD3ohZrFA3BOJeAuZGq6r32p3u4pveu3FqhLfwhlQ
zx7qDnkPTt55QQWFsWseR7EczCo5bEdkeFLpshP8EMYSmIdFNWdrhh47S0X/c5fh
ypliCbqJBR/XzT2ixiVEpoVPwtzoxnXf/qqrNiVUWhZG8jOW1wYy0+myH5njuDHm
iilu/M9PyuMNLpipkIxduViNuO36oLEB2p+PJUD0zk8686ngDl8rYB7XlXOJ75Rr
S7kDulF7NevopioDQYvK4UIrawNp/ec2JXE33IuWrtO1PVIXynLP6Iy0U94L2jVz
gNEZOZNjfbzEVAxmSJKQalRBxAZZvQdqHrIPiLJKauT7cTxDydAHcx7IuQ7uCxJL
nnt6/3va3absbsidJhIJgRlK4jsm09qHVmq/c/Ka5qiUEULSW+O1C/9AwGCZxoJT
M2Adzqz8bEnjEfVcnXwNLs4szL61AUx96GjQ4Yvnoi2s4dfXlepUWARw8V3uD1jh
EvR6jhTBcOqKuiHbr81azk968eKc5Lek895l/w5jIGAhZMJeGDHMQwNqIpPnbdps
dEBz+9AKlt+gP1VJ1oPWZ5a6MLkMrvSMb4tLiF/cJQpyKtumRqMSoh499fgBRbl/
eV5XWF1MUwsoxZIZi8ElEq0ipIj+Fpc3rAaNFvQ6xYReMtiYJLEZXF5M4w9l3r3N
i6UUM/RdM5IijoF7tu1NEwNlcmL4qJQA9nRU5Bwh0/89N0uxVR2OJE3Lb2h5ak4I
p8IAS0xtKb327MFojlFNv/q3zk5PVcP4NLQ1mzQ1b2Y+S59TcW+xS6RMm/MSSPkG
rQfSf0h+GqQ8EBpGPfS62NAjJMZMjFPRtoLoLMS2+Z0xS2vV7AMuFVB6ydl6aOoF
wYaMcSzCLUNrt/IZAumjNTiDyhzoz1fTitFWoRXRJLXRnN5CL4AOqQXfcxIcPave
cnkNxC0SkRk1rWf0tBPOalNGVvyOO5nmXWPUfAIEWKbhxjEJE0fzuFEBM4jC43JR
5e+OOtUfVf0fxz+JsYBtBEPX+OrdB40LaHHsJXbBoojgtGCVQRC0e5cONjQTPmfl
4E+aCD+p58qmXRUn9/9VfirR87dNHl9TmH4R5a/E0sG9Cg7RWPNYrH4A3U3MZPAb
y+ADSiHXN7eVspEVG4jMFaWYzG1hsV5FpOdi8CuywUeGY68QOwgzh9Sdlhwr7LsD
AMXTYa1qDGfVRb3oAcjrAQiBEF5LuTIsiD93GU+ji81o5NhhbC7cmzGptIpMjfyX
FOrB861Kl6k/SEU9YUmZOwgWioZ9jwEANWiI+640Avrm+UH7+gUdgGCAn/2ebdwn
5gqKEPkMv61ndiY4JHr3uaudgYheay7A4Vtd3v5bU0T6NCSqXt2Py6JpUpegUxFJ
Z+9BWtK1FAEK+rfbYorCXBQsuou63AouvX1wy9z8WrrZN4OSdB3UsdGljQmFU7ss
X7H+xiMLVs71qLvwBzAoL6E1pFDzBbxb87cR7ns6ts5o21RJ7YfHPM2B/t3SyOp1
5P/8rSN9u1J51HhniGy9gyc9xc93z6Q/tGdeV6v2EGciryexCYta5o6mT7MrsyAh
oy4NouphIXts0om9oK8sVHK7uImpNeZObuEgu5gnvcprhGTttrk/H6YIIicE6yH5
GO2tke82QAvM8WmAzW5i/UiCYbHVjRp98f+qm25dFxmaUkpUTS6pndvZi/trvwBS
ej4qnh+Ddfjn0aPC/iAOQcDuAJ2p3gSsqL9ElvJT5QyMd3E5CKewIm3LMAgn84z3
E+fa63DeGtVBrbSwzTzQrbouKXxU/AMHa3M+il8aq23Cy/sXpmnrF93hqnw8yXPT
BV4MbYGZ2IM5P3O259IdoVuRcp8QWh1/Y7TcXRrRdVDuc0t9mcHV/1KrTzk7KRgU
M7xl4oqBLF3vSi6V7/6Xagd0NfcLUiPQIcsStpFe57a1SfI8LoRWT4gbApUjfhDi
160xrELWkIdHssDfbEaE3IaY2XlXAx0X6+TWpoHPe9kxDqIKszGRt1zizi+1iCT5
a+WVARzUbwswwQQSkJGpkK629Me3e8aSlircMtmoED52VykgcGkFKj7diafK/kVe
4ipG8tyqrdsIgtsLowvnwNKd4PUxt2N9cZYgS3r2pgfOvKJYIVi+HXCgpLrB3btN
I1lGP73P914nmHLtyDabzLeuE+BRVS0pKNyDjl7jsfklFSPntAScwmAiQ3UYNXN4
waL8+N3hWiqAFjEHeUVRfORlQGi2QgZFfbugD2EYPQIXDM02nFUQgpye1QUB3f+z
XfG7sNsA4eJpnpMd6ZNybc+8x9rDBNPxQ/5xbwm3PGx3sa91XbYSLjODcSNTS8Bq
fctHIUS6NL1oSQiBLabkM0Jt8h2YMTixUu0pTfDMhhEg8GxipVtmrwLIdHhdvLQV
bYadw9TPM+PkVz0fKNtSTELg024qMJ8PPMD7GZSfRMAqFRolo9vOlGRMrZIWcQYP
SR9wOpd/zIthWhrvb6r9JFjT3SiSjanQKxKvnaZzPLefm8js1I7wmSMQ4VjT5d9g
rh4yonaJjZPMr02IjJ42xj1hs63vzHNQFRGqDoPbpjtlR2gdzDZWWQFr71n7s4wu
CjVjsdb1PI6unXepau81fMFsQoQa8uy7eoaRwmmY9VdyeSZqwKohFqhaqgwKox0J
1nSHQrL7XsVpU5z4kSdo7DdLjQc7isDPkOClul6vAnxriSn2fiU4zirwj0AHS0Vv
hltmNq3E4cTD0V+j8khdHXcvrJzdLO6kpDnVBS0+mfqZlHL0xiUNyBpf67Y4A5Kz
00akZiniHNYuUANwkdeYSQ+1bM4XHh9aPODBfY1iHMFrTaU6aUT9hThCwZYtZ8Me
JGBo2SUBOD53iTN00bQW4emJ4FYCuIW/UL8vueaMv4SgkfBuhVeETjBtLnLDiG2u
b/kJ6ELd+17Pt3hmV9Rnh31t5OUAj5UiQqNbYW4+t5LxqjGQi+Z67abTqzYJl/md
Op2ZwmDEj372A4/lx/iUzBIeYS2899hAIrj80sZO7f8bZEuEQ8AhCep5JR35M388
HMoP2rnHWU6f8qyLZ41/J+Mu8NyFDIbKZ16v4A6ylFQ3dFCzkFBS6Vt9yPEa4d/V
dBYtek1fJMhOmKBn5jBL7CTTyC2NFIlJdmTGbEN8pJi4iM6MOJmb89ggA1eI5HDD
sxkoIbOz0EelbMEipCfcrnPppWaB2t7QzHQozoYpFeh/0m3vSRcV7jON0FmGGxoQ
+snU2fPUTcXhAWQPvHLhr2NlRbtNo0fHF6hkJxqkdTL5QGT4/iVG1+P5likxk9S4
v5OvlgbdqNAz16BUWTj/BOvMWV0Pg0dwRaq1Dyf8UEbGCX3NpJNUDVvuQRprrxrS
C8w+Dx2G/yuAqBwPTj2l6MRoTW/NuS+fpWiUKiwvAwBq3WbJjckGhl4e6kqy8GtT
wtlXaO/B0zkIDzdwLrqo3wju5EBHKaAU4UKYG8ewrxYhco4BYL6H3RSRi0+MHdbR
ZvQGKNL5jcmd4TcJG6fl9AmlmAAfyxL5ppOCLknwtwgRIGEpqH5WZd+G621KqBKk
VJTihomXkP6MjFjo4o9ifsZSysejwXDTndpACG82UyRoybg11baAHPoCu47HUZQA
XekC6rf+HVjcik8p5pjEOjdin6PoIreZlkI/F6ywqLbU96fzr+WXG33NGWRwutO9
Qj4NMaC550vxAaFCD+hU1WXzwdOVmJdi5p2xCVXYHnPLIe+s9/anZ55MlzhpfHsP
w72oByD1BcqKa9Q5jcmb7f8gFAfLnqRjQ3jJeP409GrrHe96iFaKO5cnw351ucBh
3iGwHPSjilQ9BnaTyuZZhXQ7J+YlYbuiQe1i769YhVysrWRAcOoi4EasDm0iYbDp
kWJ3nvBr9Bq/m3t2Yfx0iBfWcvITIsf4ZTHVsdD8yY/GJATmPiUavE6ePxcF+AmD
cZAgs4c4sowIEVA/LSxmu39ZW2hCDnPj9X7++SO6MmUAltU1N+OI+/ruBKfjUgC3
7zltxyh1YB67tgLurZC8QJpQliJPfc3WZLmrvfzf/pqKnPG4WOQu8EKJ3tFk+e/s
0EX5VgehYuVydiR69/EuqOM2tuA3Y1HDUsP4eRFPFbTXFIoJgs8l7EB/J1hE1u02
6gWsdnyH4sJV+QytEn4oTl9nLMGz/wfCSInPPP7vsystW0hV/s0juFJ92vqnF2Gd
z5zLKwMYeIWACGuZLa90I7/wlMdG1UDxUl6hp5l2o+US8k2OSJmUrXLCk18R8asd
WaEBydT043Nezz2LSSbSUbfCu203fMjfz2+tgIuQIzg1DURoXpy4OgZy4FOjKe81
hmafkysDs+C2W3FozcsfD1phj6qa8c9tCeZ2hgQwhyhSyDwlXOsxy4xISwxKOBgR
2rWWbbW5vp68TA/OH0ZLDiZX/xQSoq1jEpChDKQk9Rgs/xR90rH8/4iKx1eQo2OF
hR+KMDEcNI9DFw4HDPE9gPrZshsNHGK/JCwrfXxV2FMSRypQJnLvfyXQhvnKAR6+
yyG/Vg938EC57X9XaSaK3CsqCsH00mVKROsN0oevxtMD71JhUc7i1x//zEzqRqCg
c16qxIcxFPf9y3Nro6D72f8mEmlHXdpgUOFxTl6N6Sy+EzbzpPlFgfWsg5wySl+q
O0BFuvtl6aKEF4QBPi7KER/iwmwgVwH61AIqbcfeSsqhZQD8rY+NXAtIQjy5a8aY
53sBhn63B+iDMVdXxSUY5b4tf7SfsqBLXR6mmvmjN2+P8PwSaJ0fiNrdiP/sgSWt
+KY2BE8wXNYsXh0TpCpJtHvenZTZgVtU0Y3vByQLdzpk0RZZ+A9YsVtOv/s4Cifi
Rt/sPCH90naUj7svr4HQaT7dg+VoLgu/uEEVJdhHE3iVgZa90ti3A8FpVB58J/4D
iPeLD0t2Kx5Fbkz6ldTlsN0vepfE2vOoZt7RAK13Za+DgZDjllLpkYlzKFxqW9OT
iBfRB5VPcyxodDK0r+jvkYt9uk+zzyLjWQGhHp+O0wlxuVBb3vuqQeKFKcDRG7fV
3R7BZG1DzUQgz9aNnwHsSOJVXDYnerMgbFs2E/0wLxW2kTndhXDy/I5sZjEldoPL
ZUE1Hocc5XY4vCTo5XABOTv12RmltvS8eT3V7peHx5rRB1ThJRW0kv7RpxGfUoOu
oNMUi/GaJCaug4KeJydtMSNuY3tPALmTzZOGwI9uijs5wViWX729fw/PDlCvmv/r
lS+67z4q43CxmZVyGyO12lNkYnzwI7HveScfTXNhr1gdAAyORsSQrIzaKSOuv+2A
coNcdHTC3zZKZw37Z3i4c9EbMu5jzuyTKupAm4BcdYOx5kQTf+TvZ3SN+q88iDyw
axU8lRb9r9dklVEx54z5B2BU5Z9WgQ0/fdL2rNxAW1tOjL+WejAFNIgATnNR3qUS
8ttyiCjuwVpKQqGv/QO20/WpeKFELjJ6bkXM+hL81CzLiBJPQcEiMumcYVAXH2gS
wMzqpLzYaQKO/9mPM7MSaYEXcgtl1QpMUg/lSZqEONTRTNhdQk4JPdThpz/yDoiS
eWHXGuhCblPt8YFRoI2TZU5EAIyni3UAkytPKfqQqFD7ZqgtdrVAScL/12WdkWpc
dp9wt+Ng+se9ZstSqgTFUwL9MYMt6iiI1GKGyh3KkyF1MuDxDacljL6esQHBcilN
RRm5iiTlv+5vhkmOoW/ejxvZV339nnYHOsFmE3xTPcJu1bJGGctoHM5LC9unVQiw
qHG2XU4xw3rCfGk2URiABA3t8lwkPEn7ytJqK1Nqu++arTos/s+Uo+r0O/FVlqvJ
Bskq6T1fCox1M6/bD/e4w00IGbJyw6B5XqyGNffNtBM2ccu77jGXNUVRl9/mBvOG
6e0V8npFe+E7jGw9qDysY6HuxMqLsRuglbjiF1vyXFfWGYf0EAFVkOAc+6Cy6ZMv
6owMm3muLap4dRp9rjhXNn64yPA4RUgqBQw6BANQdKcWJwwQdsJndcq1F/sRx4eS
kLvIpysSr3fLDXJ6Fw2GjzM/gM7EqJDw9MH2YFjy4lbLhqn1CkdU6Z3GoGtvyGSu
srPvipbprLPEdwyGxMcTc2Y2LyvF+8vZ36AYwt+9ksFTXD4Ycrl10iHnGSonrCQs
lTyokWOoJfSnwF7wOnq6tuKwtfYP7IZ4TRgOiNWnPIGnKgBQAH8g8XHAiThOJ5xV
akPsk+9oMOMqCD+DZQejOT0dTiXzieyyRulD1o1lwiSOOB26yph2IBJwTv0x2Iqe
YYEIqEMq7jg1wN24C7gskh8eZUlTY9jOhNCOSpeEWc/8bUJdH9/yppK4ZyykA24/
j34k0+6dgQprz8dyCrtnGKTy+AsBBLwmIy2s6eYTC6oWq0wrIXakm4kiY4C1cbor
iLXf1DBGjStxU4g1gjN/Io4jecBokeaMQjNvZih1C1/4iMtG9YwC47dGXSHRt8+Z
mg3/z/AHPl4wdcJJLagvD7Adk2Bwl28Zkp2ICaQGC8lotppRElUUsjD+t7UqGxMn
yEDyZOlnXAPx8JvzEzf6SrxPqbsQ6dBHGjjtYD6vjD1DUJ7hRKBHFpbz5NDuNHy7
akBoluEgSygKMb/tu5n65Zwj9gKe+GC4j8rUsCZSUgZHH8n5Zr9cxA+utiwUUCIW
vCLslXsx9Y8bag4qkaFtkQlZMfnHNXvN+qUYDN5kW2cU7pe5ttIXpQGz9SUlSCFJ
rR/tsSGm8k7n7dtp0OUZmp2Y0QoIXg/ljM6vS9Ow0Dfiru6SzvhuDQMTL1tO0SRR
jh8//+stAR9zE4WjWE6tUll/ssxG8TxQGUk1SEp205RnQiA+IBD3tJCXv3KtJEVE
Iyd33ZAgV06f8oPnXkcD//y7IdG8BFJ9GhOmaepU5+U97jrKydu+prCXU+d3JGMh
83qK1kSxZmSRtZeYU1N/HNE5EKTf/+kGT+Da3LkPltalklo33xcm7pmrDLDXOYU4
4+XiaUq0QP3EfG8nyKKDNytU/jPWzXp6N9BncnCGwO4NiZZHF82hyUYZjgRrtu3C
i7WIdZ0URdEhLR3pCDjeG+oAGxm23HODxez4Ikr5R39GPz0+bhZqVo8j1cUObxP7
ipjqHjRoLrklTYcWZ6JbUybnFfSE7vrRdcyWww6LMcG5jZna8ySfQ5cD89F+utMC
UUHIM+VG0tGFS02KFnP3hnUlJEvWcFSKgVrCgK7pvZYa+yglxGzoztN5unL9Qhrb
M7j0vKLEbgw+Ec/PxTTyyeOoVpqml20DS/vlT7gOWg8qC42vjka6sflT4E2/CJVB
4Qov9dD30Gay3ez38G3UzbMoS0K0kn9NDzbxiZgoL9kQDC9o8FmXzfzz4F+12AJz
Gf1uSX8RPa/N1oUtrnnNmIGF+BZpgK9lPzydRPdSTkFTC/e7VhaOKMAeaZqe9HDc
J1mwOWC3MmfwyL/tHd3OEikaH+3lIvZI9OL5A9S3gF2SUaiuUNISg22JM4Lj2fUk
Zf+Rst6W5hACXsSxseMG+S+9xDOvdwPsfM61LcCbHvqYbV2KcWWPgoYQEHYowCMo
ULWK1le3K99LVNvSVC3k/yMcm1vivVYdaiAV1VRX4OvAAfYfaTPtox6dQlfHMztg
bv9TRHZsowoeHlxI17GJTIrrp10RkvoCCUmZ8zWlzZ9yDRXMcp5TiAceS9xtufiC
YSMOOmVZQFQlX/y/ZJUT2LpA+1ciFus4llGS5E1uIdIv+nNnIjmUFQCkpbiNRgps
K4teJqYA6vzyPBhTZuM6LFSQjqKNOXrucYX+bFB5koat9mOP0EhYwFRJm8Nf74Ht
ZHAY1q+qcPofBYezMvlosXvR6UBdagRIZnDvErZsHfk+sGZcUxu5pd0PYzpkvusq
S3AqAA46YSH7GieyR6BXQY6GVK2O9psHv78Er6jFJEW++zx4zsr2vqJxMRKj3iJy
b2sdXZ1sb0PkG7r7MY3PlK619A35OGYuZL7MoMITG9cwmsUR9mPJu/OdCpPdnKh2
XTqLOpaTpSPJUQMNgvhzAC/rwUrbuwl/6jVLhsunvfNDAS6pFep4g3ppD9YbbHwD
S3x+U9Qw7frowul6IYZtALI5HGjVODZNG4E3LBAGFuyx2XniVkSxyCdbRql4SGJc
0MRJi99cW6LqnNeNd6QB2+/mJaT+2EE+RD+Um7sHRqTHPeTXi/d8P2H+yW8EelxJ
8FUM1sb8Q7NeGPE6Ebb2D24B97YDo+Z1aY0hHXxHm7qD7HvDjm2Dj0aTc59feLKE
J2OPsu6sLmTX0KxfHK0JFT68UcFnoikKHR4KyOr4pd17dPqsMyurH6VT/I4cib3a
hh7k6FijK4WMOTd6LbI3wjtV+QsMsljd8S0dpIsv49SXeQfOZzEd94A1b0o9DFfP
bngFekOFPV9/fXhoI3y449OXBZwSQjtEm9CRLGpErFVxiYbB3fK6llWHfYnkEDuW
ZutwJfYHpDUie1MMmWm/uAbHhdkQjSr5v3zCMRQ9Xvs1lqisLmXfBwFmoBWUUt6a
krBfCtE2xjy/a9kCmcw3htBSV3DTUtZwGdElI+n4sUeBin85By9X3VWUlGKWTq67
N2sBOUnz3oSpKClw2pB0M4rvPSVlJI/VPDgUI0+pWHxvm8wmTPN8S4s3VH2fDaFn
XLP6cekUTLqa2mme6trr02wZhi7QRp1UHd+d2vzKuCsYX5HjTuyt4CZ/fmTVl34n
DoiRxZhY6MS5SiEC8g4iE2kaawXpNCQ/3d1xwtY/1Xoh+wYKinq6S6+gs/TQa+L7
6w1sF/R/ddx4sBRCu4zMGMA6Plk5rWp1m9OfmlGHuMB9GU0mxYQiCxT/qHk7hJVh
GqzesdEpc/uF0ra9eNMrFi+6skIhIXnx87udoMus8/PGA93nKqWifms5qDY9XpGJ
OEmf4Ua9lRZkJVDBF1RlQ/v/1h+Ujb5id9on8i8ZtLO9BFanZtfHxAmyx6/16BxF
uV6/jNofZcBf+47HL/qxJdonYH0ZhY6pNYPpo/v4Elu5K7dKhx2TrtvwcDGm82Hf
x4582L+8iO7X2ocwQZdYCVXyaBrPgh+pEDyQ7DvRdp7maBjtpA7lzwWnIj9dW8ms
kMuicUuvMHc9pzGNcyW0fE+24t198x8n/p9Fx29iQaLxs3kDMeb+99qUIFRC2hjg
BSNhSbQWOubyXwPk6ZgNHY8wpyxzhqN1CnRP5/A/HzQJDbZmnRXz+nypfe9cdM9Z
F/kBEWFZTgp1hjx5lYv6h7dZDGUpADFMn12s+UyPb7NwLhBRw98YIu7bWfdeMbXm
P7N9KXlaeyqSWMdW4+ba5P33x01EKsFYdLOF7DbKWm6KgjF0YS0qerNY3n8k9VNR
um4J4nPg8ENZ5O+Zns/YsSscg+60zGkZmZxiYtFbI8ai5kEUBQwvJy9nJVyw9MuG
0Jo+0yueP/t5Lq3CeTL9cU2bK8h6sx9CIxeqaGpICW1BG78Z5QdcsMJnJMEulL8x
tAR+o3GICB476VqtCR8hw2cHM3ofZwYBVxt0uVA57zaEgnqRwIxKhHMF/xLqJbwp
lzlJ2fO+De3Fy5EHpDAowHj3BrhV3cwZCShLF2wLtK/sROoygSogCetCg1ZmWlFx
2upjODVxDVGwu2FLp267X6WsNU/Cq9yQa3LYmblQqaFE682wTuRWQufsqvxxMlPI
0tH8YkPk7+iIW7+vCzG4KEn8vIePgZnvIkT4cmauJp7ewLmwUeNWsFQmchx46Oh6
rsJW6y/Jfq60VAsCb5ty2tvdEcAth0wLEzK/qYHAy0Ifp4dkDxpF48jopDqHCF04
fRQWx5EdE+sV7LKUIKIFmry7VVYQds/YEFXPgI6xRQazQ1ui9CWzp1XrNW7u8cnH
u/WufSOtop+lECefSF4e4aLKmFeeFtnmCsJRUxS6EVne0T07Ti3PnGXSrXJY19Hd
/AXju+FaeVflw2QzWL87yqfD/Zxky/aPNorXs+d6dV6H3QuHy2s+q7XbFUvFetR8
HhmmC+hW/bapIoy8NAq/I46qrevKi65fwDR0y5/fRrm7XFNnJ8RS2uXh2CYCzriu
op+5j6qA8tmgjJi4KINzBlMb8mgcsCBpi76TzHzoPFBV16gdu147O2E5RYLtDmfd
GpZm2jZ1PUrsJRXXvS9VFhn8A7XqocDbL8DSaBO/Ehur+VjZ7aWYmtZUyBr34/Pr
w9DbAvdGp94Hl1ODrILrPYFQWe0iYZR8q0oYrqj6OI/PnCTGu0dTzyQesn8rpH4A
KrUCTI+zo7zLT2NmBKRMHuGC5jMz3OcRyuuktnCbCtnfSuWrE1Yjs2QuY7sT5iJ2
tEgP1qK2V3Xbaxbgg+hMsbvgNrFP9dA+8Dwx0zJL+/1dAjQ1DdOTPfnQ7q7CmU0S
JSmzf3/ZERlaYXYwxK8v9FoZQpfIsF4xH3vxTEcuDcCaoJrBKfDMqJQWUeXaw4yb
De+lSNvGjEQ2N0ZNjIdZV+GbL3Cz4dth9OLHIT+OhXYStsAJiSTLmPSgHIngbdsB
eEOcPqM+H76Kz5V8ZFzyJrzeLSbXPo1+cui5QlZKtdDMP4ean/HHLCfuX5A4UeXy
70f1DUszDKJY/Kchfwv4I2uTy0OQml+XhTZ/CI0R78x6euJXC2w636WFZ7evjuVK
fY48IHwbban4NAiIE0KsqwhBkGP4YMxmqeweWJeB+il2aw8R9croX4rhrL4M3KkE
2H0/ODeq8Ie+WwO2wN1k5qwa2Qjw+StYaiRHTby2PDYpWy0Qfkw8ujwkSa08THcF
XA5Fny5I14Y+36TRMDD6ApNOXJ5CnMIE+jWF0Iv07CvG+GIXa57W6aAdusZZx7Km
ssldBB1i4ezU7uh7M+4W2kqHrKAPlxoind9BtAq9JMV0keXx0E7W4gtS306hW0K1
lU51soK51vctLYCSdg0oD3DRfSSbUvMFGyxDnVV1HPAeR43mEO04Cw69EkC8Mkln
Uv9cSmCRApS6x3A4SLCfF3E3hbzmQPq78EebbfjEZsu9AZbhE+WQS9M21AKPY5mH
SMcXK+QYUkVZ7vTnBU9sXCg/jzrfbS33IVOnoi16th9bPejTs9gmVQjDCfOJvjBL
ZgaDzE8yT2B8w/THLZ3ufcyNAvfUqKfndNS4X7l5m+p4ehC7rRjDHeTaiDb1e+B6
qV3vBlz3FKAt63rPDz7Q7IrWBcTRbOG1k44mNCUzgam7vWAqMcYC87jHzF+8ygsC
LkXqwSX85ZC3C7qp7qRkdjehOLr0aBDPsOoifAGOGJWKDQZpGLCoHeYpEAmA8LOe
RaAmNjqeBK4qJhTx8Gd/Whqnb1FTjoRK7Dr3PwefENXaooR8RNhbWxxsxMD35qnU
XJPrUG8jAOn2691tBRlHZI52jrUPC4Zio49jM7cK6I6apIzwccUYsAsiBIaNonja
TcO7f+q+NEh3mtH9OBArras9Z5gq+n5UcVOc3LJRFSOYau8FH0lFKddQq47tZQ5b
C1Akv8RfsNmDqLIrGO09bk3tVxZa0qKn5YjAObTwlmybgcKn0+jQwYlaMbXXROOw
Ei/5mgfi6D6jxrVH7eq2s5pTBMackjPAbuac1wtqcwLIIPTbkx/oQtbgcNVwd4N9
omWlBvbcY+3srBzkD26DSqnDX1NGwSfsEY5eINU0ul7Yemu3QdiQqPDklWPVB86L
Mmsw6Bdi0X9Pww9IZf5RFUZIqpNCGbFN7rXhPPlmLt284bIgY0p/0Bkdd3fWtBRE
7iuNLH/DNpSKVZrjX/Xk0/bO3TN6/1FZYqmE7AqWniKgTtEnkN9Sm4+X721mgVNR
hvnzcxZW8Ub/aQ0Jgt0Rx5q9yUGR5cUcmrzAweN9uNpL6SS5van4VOqUTQnroWS7
Yq68FUH339P17d/rZjBcHgXHRgdCfaSZjyPlZA6u96BbtTm1DOhKua7hCtqE//Ph
DnhKE3dCNpkJk3XgdwETGTY/qqJwPuf477x5ky49iGJnr7tCNOIvESRxj1tJ7G3Z
zxMtmD6TsSXXVGez0jvHotluabBKNSUJy0orWioX53kL0dwKoEDDMp8o90st/FKz
YSbPo7bkkKiIwewyBoVpanTZtBeMPg9SDIr+jiTcapwMXTHHGzwICzRphXMh6pOS
6Mnx3FLURTSYZmrlM8azscoww+FpM/QmQU9vDvpBisnq7TI8Zc28tke9S7frU/rc
CBEuhaD6lO1qD7o13mXzMkuA/laI7oA2KRL8pWI3Yk6hCfxoXv2ok6IIC14ckvuP
Up+6HhAlwNdQhrwz9jeNYoe4CyjjaXmtD5rGxFD9tHc1oqAO2kg8xnt968JZMiDx
OTz639/hdkOwdQJ6bhzNY+vyQRJIWn6ojdoubcvFpFQTXZXTSfz8IPio7EQPrDyw
V+rHHelnw63v9EipNnvvEBTC3TdWR7KNuGn5iu9LKUfW3LHanf4ylI7i4XkO0hgC
E3T5hzu6DIIpXb8boVVNhe0PKXzEA8Q3ESN2zZw6NcKHHRFqvCmD68ZvbfwY/+7n
Ue10ad+I+TwLIFxcSshVmWI9NzxfKxaJCo/zi7fJlBRJbjV8dmb8k0wBX83oOZua
JLwBp50YWYhWT/4TBgpXlSPXVecyCcltywKfBLu1ttDZKfwsrxMDqwaORWoqTslA
I7qMxtUI1z/lrm95t9ZwvXR79ZXvu4p0L1Gx/zP1EE2peJ6C1dcI13G7JKpN0ctW
M63lLEAKiZcaWnrVCWExFYgHJ0NCWDzBn6DSoUVJaSS9AsF9V/5Mw96tUTSu8jKS
zELJxaL7HC9p0ZAZIgQgnuoMfOcAZcSKZjxvEo+9R2tWeZdTWqn33ztrENYtXaNH
pfuVixzR5RBRczTR0foxBP4IgeaHRUIAomNnMNRIC1UgjDprLVCpkY6B4DI307cI
TExcL5UFua36xzjMhAsBNWsPDq1sGu/+egB0fibGeBRhFrFSvX+ZAxjXdnFAxpeV
qkIKldeqiH+FV4KTuUB9ycaBP2OnJkU5Dl+IPJpAM+kA2mhUHOkywNtOGbtO/od8
kLFgv8EaGRIEyGaM2WEcmTXHbAhvI8edbTX1t1toSZGeLZEz5teRbSLULkCSxJlX
GxeApoLxBu1WdKqHz2HsTfC1H1aCRazDvZP42lNQygfxmf+5vRN0v3hyXLuROTHp
MCc57VpZgfcbX2K3MjtpjpljNiPiC0dhZIhkcAgWRS3SYlmYBPm2FbKY6H2XaMTv
fspeM87pPVCZTBOE3C5bE8R6184SuGyp3MM16h9SlLBQStP/XOoylGlar8yHdkWj
ARzqE+/O0l36Q4wH0G32xWgi7qXYwhKpoKnH9kQW5BsfHg2PganGMXZ9a+LmPYZM
n6e7OXSxwXuf3dLGvqCgOrEea1pu3/fCaR7gsTM2VDVrQt0cr0zNYi7zfB6HIfSs
DVtfxG3lEtoxKF+YHoWlykmHiw++diz6BcWx/Yb1kh0gtBeqJGWbP+7rR2oXHIcJ
2igSQZBVoTEF0zHRa16KqrsTDoaNmXxB7mThkgCP3Hq0FCI/Ny4AEA3TYfJu+NN3
MbKr1vZiKCZmSbGFkN6IBIpCDG+pVNVMYF4O3mTZ7vnNm+otFD6TfZj9vmROwisC
DZhubn6VTDiugUauJFO5PQP8A5ZzAKDgpXHUiYGmCmk/q7O2vf//jXipMowYh1w1
o5f7GOQi6MCfLEnwVWgjxMDKOY+BRgYTff017iFUn5WxfEgXWIcZlPkXkPcyYMP9
BycSMMqq7w72pbf9CWi70Jj5OL84Sj5kTapgl89+2HCBIwdb0LP92BTfIXHNSILl
gumQSCRNfok6wgxW5doRzezakgSa5Ljw6NnI+xQbUuL+JGNj4zCDqQSFeb9nZlAW
3sEYhUZw2trm457GA/ZViWGkk3EZFed93MqVaqaPhzYfokDJNS3d7pMrU7VovNyW
5qJn/ObcG4VgB36cDcR1fCRs0KANFBID+UVowyiXUyUV9aN4hkyzN1mAuliRyRpU
tNv6hD476JZ5AJQBeAZk78NKsNpJAWjOE7gzSGL8wKsFo08yGdWc3RK5f6OSjkfj
/mgqEQrbtp0LXGo6vYDSOMCFrevm/SVgKuzK3s8IMdJWTCz16i5vSaV9EBgxLmxP
k3yhpbBU0ydFVgRpe18DnQAwopMV7kN8kZE41I81sh+IKjZnwwuKE6ppqJTtJOhs
hGf+QXP9+eolXP5BpESYolfbgfUY9lOmdVOXIugX8rn+oPd10Uf4/WiGF6wXt9PL
syksBoFPhV0l4dJwBP9pZTIB1lJcYz3XXB8Rum/173tifW8NQ7LmLusbvBZso+c4
5UAlidHVROQchFoi4eHa2IdLvvuDn0hJ83+4PNVE0JTGEwVZKUrXi/Ighp6VhPdj
/bjTFzv/T47Umtv5ayPGnys9fGoZPzyuuczYBeGGiqaRvF9QB+IbVm+GL4toWNzX
/R+84ZVq+UnkvJ9gMqWLmSCUMRhJGNK5QQn9S9zwVfT2w2p0ghTZAPmLFqXMkUGQ
91Msvv1puBQgrfuP4HxC81EN9WA5tn8CzDcU51fEgoILO4Zs8q4UYs3A6w5gdQ4g
+ahCecnpMb/zNDOlfTdfHs74YM3RXN0FXy19xmx3wclDb4mhuoPzdIpDOhPUFUI8
bHYXk4rW+wU8VpVbvM1AV7wD1wC3XZ+Sqrf67Vdi/8/AkmAtwvUVMRAhLUTJyquw
J1lAyvKUk52t3LsWYYvr1wkm9CqFdijBjfhu1rK8vZKB3v/Pd+3wPuILJsIG4SP/
5aNk5lIhfDF28rQ4NHWt89lDCTO3ytFGyxjbOf248dllJtBsoBgJfhzjgGVrSYlB
TDBpK+1Mknb8eaD/lr5OrY5Df796yiBOEWje6blgoUrr/jymjJSxAmZ5ibwlVE9+
9t5GQ3PT4EQSUEdoAuTEHMN19MMX5Pij85c41vW17UC4IlAfmKCF00p55sYhHzAy
8pzNE4LCIF/O9C4E0Y1iyywXO7icdWPiN5VCMVoSrdCYKVaS976iOZ4wY6Po48kP
UW1Rak2Slb7DLW+IMOK1N6fj6cWRR2uPioBH+HRw8i0Q9jlJclvGP2kj/d2oGqPW
Y4ML32frRFPXW+5adUeJkwsahwXjpKWLbtGtv9geq3iqXkIZ5XO/goV07Mnj1iKS
GohitNXK5J5317/YoD7BCLj+YIlJgo36UYH53aFPV7lmSoJ+gFUBPgzR1CNzE8bx
6Nsh4hYMqz8n+2ftsR0zwZlj6vibMxvcVYkwWtrKrenYvRcIYbr52i6nUNmbn9vI
iYFFaOxEkgc/tNcqdg6dJpuiUFrqKEF0iHB7CkouAE+mSopOlHReYqwbce2Wp0wk
LlL5Hd6dGRrZ6AiyOlKT7w0w+QoWMx+/WmlnYyqfPVgYUEcHOyHMfeCPixM99Yrf
saA3HEwDk3SmMViS9OHB1/ULyhDcaFlJhkCv+3EZR9sGXPWjmM4lVWrlXpiAh26P
7taNDefBXmM/ntEhTR2Niw9/DqHLmuTo6Z1eIp+Eo6YnmmM3D8JEHezMQRHuLdyc
Uc+/FiGmQR3SICVWm8ZA9DJU2wsab4v/5CsG4TegYQFCIws88+3v76LG6D9ipdOa
wRMZtynmKgcTa+MFKlorAZ3irbyDjGE6ns1am4jfAF42FwEdIqvJmrShfJkTPVeo
RyPOtxk9WxRs9EnX3y5r0ORpOttFOgMIJMdr+IZjpNpQQsJrqBuTTFprdm6hgYaF
e4tzS0eEBjJ9Kt/X2kioZaUn3d0TjmAsyolShcxME9f3AsWuS7ZRyQQ9CbOcSETp
w9Rbel9G9gf4nvwOsKPdZsJVxRgAR449N2Ja7FSJcpzvJHFNjclTV4+dDgj2xg+Y
fE3kEUAlgMvMo3ne1kQMdt9YFo9n1bg8kmGQrfUEF/2xPJ/XHB2Y6jgyfQ5INyLb
XNm3p2bpp9X4uBN2ryVf7Yjk+jQTCX8J7HfEfEHU0GV3HfJ8lRCKnSSHai+Ms/ed
/PscxO/IjplUM4s9H9cbOVE6fcvThaLXor8IqOsdqHE5wSiyTfbSETIpCQZIiz1t
Q9RKC6aEjG98eQ5TC/47WVTcD8b7YcpawPYGT78KJq5yq2gcHxtSCvpsYkFcnpcj
DIGusiI2ppcKYrOSCCwIZMM/m5ubV8nfa46yglHI0UHY0HLM1T7gCbTw2UcxzPzn
8KU/xG3Kxt8tr7zHZ7ZNlhMx8xpp4OSV89hzxvcz24Z3+bo8TsFByvARvivlnM1i
fuOvCEcN+e5fvUL8whZ8knK4EuOQlr1Q+e6FkWAzig1vM/z0Y51UCA1XXNn8X/6b
EZrrKnzqd0TzClCxyV9uiG+asmTBzFdlbGubrXcXKIFD2g//5JDP0dSYikGlKV+0
bhTUwzzMI74PNH7KPB1C1OWbNML39JQW/Jqvg4V2IkBVqU7bkguuRY3GqLjPOzbB
KLl1mCM71Qi14OraZEkUCoRL2bBxnOGaoZPpg1gbbi0lOpCeG/wBwod4jyaDXOma
s+aXlBhDxa99qd+UoVwdv93nj4MhXQxJLN/Cp/f7s7j7Z4J7V+ckiJWQ8I0EX7ZG
4eB7Tvvft1aSA8sMAiUr/3n/RJC6/9whsc9mLEHDpCfGT6XapV/VmlwCdY4NgtV+
j4LfbCBj5dzsJHRcNJZXyBjoFbLH3FomHf1syzjBvAi2vDARM0S4BxQblMSFTClm
6TlkcinZISaT9Dw0qTG0CeJYHt4Ni01lj7Lhk8TWOnHjo9u+tQPKUi2CHMnKglIH
hkDoo3ZCnGYFlvgAnbMtkVda9EWmddQi+4r2Q1p8m0iDUn3eRqY3BREy55GTpD8w
S2Oe5/ZR1lGAJBhy2Ppg9fapWyvIOllJYckcdPsCzXP0Yp4xcBTZ94gGMD7Fp657
Bdd5yQYPv9JtEaNqdXU/QQeLQstd0f3bNRjBgGE+ML3cJU8lqBBH7ipTAieznb7F
8QA/hOxmRXWqb/XdAoxeKmOSVC7+9L8jw/XrnE0FE1NbWslT7pytmFd+b9RusOmI
IgmbqKNHGMixvj2laggyiro/vHdb9kU/cUtUDm1zifdjSKXlcmZ4DW3sTsg/gPt/
mbA8JeIrGsBRn9/H0xyrXlCHWSto84yNtH13P6O0AtFNhIjIFF/n2zk51DHeDNnJ
UlozDbb6T24iQbnZwmLetpLJYhbOOjZs9P728YTAO9XOnOnatRuBCuMroAI5V1Lk
uW9vHGMFkwN3mvox1v3op/bWWnBD3eUnWbjWuUaNfryqd62wV33bsHWqE61ZHb7z
hVnUQClBjJPxE+SebkXiIXyrIya+VVEWRsaqhBEHU3/5vKVyXV2roNPO5GXeZTvF
uf43nr2Fp3sisfnYvgIkaNHQDIqVKA7SKjHkmc2r4l3cI/UG1FDuybbGR4RY+3li
OcHCxL2R8/y+4GV+5DsF7HiYJAhETKU5mKzQTaDWRFVON4uQNGw3Iu6UMCfgspMI
QkYZmsr5bsLrkORkhjGlpOx2beCcrbsc2+wCdP14rMIuEU1iv9wnkkz2Qm/bA3zO
MmKCJDMiFfR47TQ4+h7IagPMZkcCKVKatU8eqJWFd6O10Y3dbp4DOg0X8zJ4CO2W
PD236K/QMgtFlMbJ79u3ugZE3rt4n4q2PkkEcOyagOpo58qECJRrxtLrUKbqxaKr
vl9rYJpRALRNidbguJ+UCosmCAERe/ZbSn/XtkqQR9dLsDc+HLNPFNvV+XKmPEsB
APWjSAkG6r9WAhIyuFnEDgit6VKupcqf6YjQY4lYVQExWeQ5q53RJO+S6+llWXRf
S7gVdg24NsO5RxbZsgYbnIpMhHMfLSO451cFc+Y6QOyzRhS3VEUbN5exQRjAirKZ
p3sx18y8VEQbSuJqTw/ONegbnJRxxHP0k9Fcjhx/sqgJU7i0Y823ohrhWB9Tj/nw
aWIRMnf5tEPwasmlMIIIrlnuFGAPt+xGclLzh+EpQsJ6FEPIwP/R74EfBLoEFuEX
kk2C49ObgQZNnw5KDk/G7H+/kS1M38yXuOU+hh09NGBy+tHdaTuMfRNkFi0/skWI
+1W7NpABQLhQL4fnX1Q2fGjVu0lsIlp9eJCxDw2xP4ceE6m054Ae9vk/ZIdp07mT
nq+Pp928Qmtv5l5n274zqp4VgaWe8Hn5fiCEmPKJuMe33sVCLYVkbA+prIua23fq
ivmvNuKbTD300RxpOBWFhRTwYw68pS+4vstbC2r9A7j7xo7CoSJ7sXhti0EjkFJb
boqd6PwOABkM8+XMiVMHHvcWYgreQhw6y8O8Ayf5n2V1t/E/I/JsgOshZZ9dZ67x
57uXtSVvLTZxGUA07tu7uSj+UWAvU2va5quBDkJhWAn1drYUKADUfg6Qq+sHxJhZ
aLGzBdzvQZjDdAArNj4T7ar+uoavpwLHngPUCs2wcSDH4bmqDzKfpG/ozaLlhcdU
InAsNvkwYtIi2VUKBi9AABhY0WWj8OdKPoeqCsk748arpSpoxlhyyAjM26gf7w7P
4E3NKESzWhkPs+KOTa80daLEEuSwdtDQEjaH2I/5l1AyUI+07y7zP96/cjdxob+O
wKFXFnldbU2zRe/VpJ1nhOmhMIup2RIEvtMH1Je8ZthCG4Dfuu1dPdkRmccXDUPx
VTmLqALp/NanmH9OWRIci6zbN4EI0SGCW2mhg4+AjLaxmlq2yGPZsumIUOfulMaT
Ra5oEeardmBiX97HMS0zRgIudoF3IIMX15h5HU0S7EFKaZYXP2xjaqnSjWZih+ya
uZ5P5UgCxJgpazliVMeD84xZyUsM4BOrM2wKcrCGqUMN2vOd1pc6gQmrDwXPsSeV
rKhTO/nE6SJYkSoELA4Ez9pHP0gcv0AQ/tc2qFxpkowCqxZtxPUAutltMYEmkI5A
iR3fTOQoudB1oMM2n8wzYeHqiYB8ljylkxSwPwW0X30sFjCruKADQYOFbKEVu0pW
c9BR6x8q0W6d0NNGicEsINp8qbnSD79wtATn7dW085+UhxyH6bE95lBf+N44IgTR
IhY7p2xUMh++55Gdznq+PWtB1XjHiO19XbWuhHmcdzM6hY3/lPBFOJTxScaDMIR8
/PpwhRr1qUoBOgFPDfBkL2jNm/3wRo2BmfiWNv/UpvZeZyErEW4hCM6F1GGTHxAh
hUcYv1u2337HlTeq8PFBSUQY+EwVdchypgZ8A/hkYnE1BtA6skidFz70Y4kC6zPp
wMvfX++jwuwveEUnntGFRAsuPIP08I7DeTM9/tgnO+VBJ7/u/Bz0YFDSx1+r646a
vZ9HJBfZaYA/FweKAMmpeA1spryMh99oEDFjeKXZ3dl+mEdnJDFYAetDF795FSLE
2vvPTpGl76S2glhdwr0ve7JEWDR0sImOOLv9uu4I8+Yh41arlznCYNwGuYz8VO5I
RaIcZTgt+OipQxn16BmZXsvMOQRTuyhr0nwb5XPUuDK6e/1jxYjJX9Dt/zGS8q4B
oRxlwREUcxsgIbqhlx7gkyDVgjWBBluENaB8HmuxJpNdVV6wFgicusowFFaKVkZw
XVRwcwkdO5FDr7RsoCIQuogiA0pBC1yHjatlBmyVfjj84E2sJ9rjoWpUeTfttDBv
qeD8t7ymN08t/TG8NT1P6lJlbEbrN95w3gbeoh4U/nh/oPILT7Lgkr+XFBpk9DfC
HQh0hiVUlkMTNhx/9IPCp/naToMmTemXqgdZCOTVBrTRkD0jqs34gSKMPkowtKfx
p9YcylPmwjgdik9tR6+uksGyoW8uw6SVY9DZMg3VhWH26giG/h8QxPelAShO2vHW
HVQFGu3+prqeBX3JkFHlQyL5j0O+iJGVBVd3tAuedh3wm/J7WhCpktfF9iR+Yqj8
vRrAot1O8aVqRVcjjLwgy642DvSwEudlNWa9C/69Ty948IkCpPpFyP0VY7lCdGxc
Y2JXNoe1iyO5VjshCemnLY0I+q6C0mdZnvl6mlfCesgcQPD82F3CREojm3LXzFK0
SxdnBIRJVBuhULO2hqI3qA6Ob+R6awwMdD2hnl1aGDGm8zMYb4puVKnuVoDo63y9
LZx7uWDONowS4K4J7a0VsYCf1WS1Ro9oz2/5P7sfuS3mSf3ctH+WF3smDoRMko+i
0cM6Lm8Ij1/PXNOWQgr26j2juPt+ksN9VU4La+gJuJ3uUr7nBMdNsTQbGyZwlO4Y
VgnPhbga3v1l+XRI4NlHlQdsYG2BK0/zmsCEZM1xZ2n2BpU574iBn2+vTdEtHCuG
yC9p41vt2EfBDxXrkkCenGfXgqMcOVRCNlDKKrPiUsb85uKn3ThiyuN5zIvWYnp7
ebJ4psfLNtu0VdWPUTJdrzhI3VSalmWGuBE0SU4fenjLtVPgnrWLczOm/LJBkbfg
fkVNIDWN5e4TxLCEQ/WNrnyxBdy+mLWsBmq00YMKyCwK0EYXvhGUH9+50lcJJEGD
cxbkAZ1IThBaeFVJ/nMSL1Y6qLxBPx/A+3hJyvxVkIf70hGQr+pM9wClBiwibldP
wCkufK9E1ZabqJNhsCl0Vno2C2OjjQCnScyJkMAglBxYQO+CJDGlml0Mt1Z2pqA2
ry1+CKXFvLnqUs++LbbhkLaVc2OmhuUWEt/H7Cgym86mZnhtQ9z44eFU63/0/sty
Eu8G4ugTY/V6xlCi6qQjwIa7GVnjyIsQOoSilxYmkTUiUxU3+dlGBs+J3ZRlMwdT
2u7WzvaLO3OM9HlUhCNFKzoCdc/aw92+EycTtt2n8200ppGPpuxyVXFvxUISt1qE
Mx59vPM9T0PXiG14USGxDbjogrRJHmR4Jemjb2ujJbn3Tn443yBzJph0WEMXZjK5
jcs3VAai7GbQdBAElP25k4vU5XK0zevakcAjcOfAjS4dA8bKEHL5Scx2fqbN2gLL
611sGpj+7ON81+GsBYzFsYj+GYAkaCK5H97D7dqREn4tw/u6jNc+ly0xfMVqHDue
b6872rpEq5MxTBY7t9G7vAovd+UFv2jpZSAMfDzRIzlCQ1Ocgg//t0uytii8+YH7
5r/DHWX+Bk2qyKNtiLZNVNt2GEkDTEKD9tmSki5x584+sh/iViDebLao1/2k8sVW
XKg+C5g8GG5pIq9hBSEZw1HvFY7pHbfJq01vD9/x3sW2gOusE8S90wmJcG0cAw+8
GNiATPXYSopUSkBWSOsTje3jhcT5UQQiGV595qWyqZq1N7wYyM4s9dgNYfVJUL/B
zw7HwhdS3V8axGd3I6aNQNZNOGtv5SK3Y5nL4zbCrjS6YRftIxTxS51atrHarAcv
BozJorOo5dypcy8oRPf1zrnLo6hX0Zte1RrKNJ53x6jJxFz4b6oPBASy8TSGTS//
7pC6q1/gdXpG9Iur1GM6p5Fe3WGLC23VV6lyEfjkmQScMATcAqK6Z7G3a1X4aac8
9YCWQBLAkD9EqZUNZah5DOLe8qhjygG2lyG5s+CqsecO5+DtcZfhhzzKybm0a+nc
KkPeE7briEQ/d/O+RCGU7ilpnc5exTdqyM0tODA5AzoRY1J+ws/oAEbOapyX9QNx
hpAPOhov78whYPyKo0DsNpz+r3HTj3nXSR/QQUguXj0qVYyDSAlHb3jTaFIAnqKs
OmCqUoEz9o39LnD+j5XMkH589suh5v+OSIG9IM1H4qH59oYZr5EQsDfImSPKQ6nu
hboyUVamA4mmIjXY3LPPmuj4ycxKn0h6hvtb/qbaf+MMZiKuwU0yQ0vJykzZuJ8M
YgVLGD98ep5FnpxiVSQy5Tn9epJO89W6HKe0xQ5ln2g8d9VUTsBuZVq/zVQzPEWX
D03TNO77l5aNyshbkfXzqqPNO4/mmt4eW1ELm8Df0yOdnEZRm88HK1YNmSigCLmH
gdtKw9y2+RzDFsbT5FG4MpYcT1Z77xZ1/atchlv6WLnbYd7SfBDlN6eDUhRiRF4R
Oug9tqZX+OLgBKiQT6t8lPdByKK/3uPyVIrD7kP9WjreXoApf7phbsjtQp0nGjN1
ILsfXTaT0Gy0HGM33/G7/ZK7VcQzPES6WrxbqOiw7EVl5LhhyLpuzM7ohDgcqicK
MvN/dzcKbz+LXHBYiMxPIWh4vlWTZSXLcvW8CfVLgvy69NJmvY3IwNWZ+eRyQgJb
Z1OvWOXH/l6tuw1L1IFNLZ7WHALmjbsCAnZDR1xPMUUL0odS6jEaGyVnsSSNoVTX
nN/pNBu79FWmuV3ZyJ+Qv7szI4KyoPm1ncgA8h54Iu/X/YOpsnO4MtNcQ+wKrl+j
0n3YVNRteHVoBOHwCesxIgGCYrYZnjkmu8lXI3IlCZX9vvOeHEE/ejtCr9Lgseaq
HRQwoQgc8Ftt9+4Qacr8u41o9AQStXXy5XH9Lo+MHW76TpyqZ5LH4g1p4SFxO/6j
/qrEGQZOzgknNKC5Hyvu5eF+rsQnptORo/2S7SwBzq33Tmt9X6+flA84kAo3m9I6
skeQZQ29N3KyO54OyrWXlmQSJULOYVhSsvXz+GS295vDc5GnLwVA3tIvNQMvfAXo
5+bLYIgGhq1BSIgI5GQV+3dAFWyvvFi0UlLFY2jm+HX81vKPSe4oSNJXNdJtSYAb
i48m779veQ0IGkgdskyB6G3XdxYz7/a+3AEeTuoKjCh/U8uuBQRzHIewldOQlMmX
Wps3ys2YT/hCpBryqShM0h8xM3//8CJNvj1rYMlUiiR1L3doNtBOEHAxi34T9IFJ
eQsxaeLZPGJgyxQd3V0iNWm5gKjpruegFBIeKLrxnonXUiORqhmMoS4beRcgPegd
6ooJKl10EgKaE+qiwbyRTNYTF5gQPz463TqfMpQ8N+NJ1RfBR+80EhWzmvw5urlh
FrBS00y1xGLXnSzYsDIz27lvxSzanYW4e3EVWHRO5fu5vj8WtcSJ/LnV1RM6AyFL
ISWhdhOFNckJRBUQ5hrGnXjADx40PDq3aXvF4ACH8GUlExb7OS49/mWM7F8Kc8Ab
CSzNlG2qP43dRz1NnX71T2dmPPKqZOUAGE3anv4/XGW+G+rkft0yDhFeBzRwuJa3
OIYSlNpcScLNOqEw+EMHyedEYra1u/Hdzo19XgEcPB8F9yO2+xSnMFH4RFjJyAoe
0c29wqOiOXHbtzsvWtFfRrBElcR5x52n72lFEQmPO45SSnE81etKMbV5kSis46mT
clPfg5YJk/OFEOyaNtCKKU0PO1DxPiMIiwt8NEz64HLYykqaUTGJiMRlJz4DLh3U
P7D28zfn1yVvC1hzdsKADkMiecl4G5orDRaxC1VRbtLCSj2TPA+GREWZ0JbHE3tS
9RVF5ElAczFbKXAiKE6b7c+qyQdIVPr2bbp/N6Q4B089TkUtA/0+JAexwHMm7JJJ
sf4UGxfsKCaQ/+81ve7Ykip1DwPTc6lpqYCb+5kSv+t/7MBQpRu2TaVwJYls4vAg
iUIW8uwvt4Fj7IT0mhnlGux45TIhIKcnMnpx814klGwAR+syMhwENkogCEUMEVXW
cIRmVPKwmRG3BC4l/LoJf0R9mbJpZ5EWFHyaKDFUWisGfDOswEkm7ad5cryYJjWM
JQk+qpAq2K+b7NzkMk5BPI0+za1V0tceyLEaIaLM+n9buC7NjCLGP5RxnNQykTGu
rEXXu+SWQCMx19JWh1ZqE2Q1ipiSLs2s9QfFBp/Ia/NPzOnO3Biwq3FcicY1+aPa
FriuyvQjoF0JNeWKwHLcomRauwNO2WWdVgRgtXKgZ4jivpm5+FTwK2Wh5cCJOpq1
3el8k9e+e/OMRz+UJoRR2J1FdEy5W/HSGimZJFtBl1Xhn44W9FsiH/XSzyt3NPI3
/HeoeSrHpJlmB0TLfIUgLVrIGY1tpComRMkXMTgfLSLLb6aLxBqUCjUZ86QoOmjI
QzB5uWqPMsNhWksu7WGl9fpmunOp86/Y9RX+DQvBHcVX9A6udjp87UxFvDzQyy3/
v8xz25jq6GGNqOU1sTeDSNlpRBRkp2t+C7x3KRWuumNJ/IzNtz5ExKXvPZUPvpMB
zQJfG71mARhm9ZmcrDPXPJq1c751RGYxbPHjmlqN9553mJ76Yay7Xer3bilM3x7s
jSsTwyYJPzSOjegnWjb1cEHH0grjMVPU84FMDDYfRuiF2zJfyil0HxJbGg9KExkd
IEcDbDTbuidOkamZ8jYyLyJyBA9Ck0vt/lHvhwkhZYzBVZsra4oqjL2X5b2JgMCx
zwfVodB/MKtupSpGl9Fy739NCvo/kfSy5VTaSofCq1AOKxAGq67hytLLR2XHpqFl
xv9a516CfMzP6lloq706k8qroBR7mM4BHp2g1cixVb+Lsbc+aao3OILuqK/KcFKR
FLrnwYFEE13+YOR+ZTejjlJedYE6P37UFua4/eVq2S/ulmI1Q/I3H5noieHAUclg
4c5jBEwPxsQYpSagRXtWJU+iJTrK8oXy/SbD3UxFbSZH0S9RBV85E4sauofg8TI0
ItSzbuOf/R/fK4vKgvwuxjDpP1ijW1m3DMGNQ6qU3PzQ0N/Y7OzLjurHCHhlAYv9
fOUZBLLbI39iOUQsGNH5q9/R66TDLbjuCNFNL5ktUKdpsNEiqfPOfgDbLBxM0eCH
a84MRgQGVI0shDgBLZsnwQSVH135jaqg1BCLmEihcww729XJG6FAdabq2RZjdzdk
K0DZuOPFkg0JAAHLCAzWrD6ZtONcniU7w6KxQfqhZAlqBib9r5eCcJ4zEfrfipqi
AZxqp6mC0obUrAgTLNxNw9OViHWGfMA7SZm4ByrHnrO3Bn/vdn6aVSkUhim+XnNE
tZSj1Je69lIUBoiFCOFh5UW25BCs+6hxl7FKkVVNMN9Dn9ivQBTVp0ecehunQTAj
KVdTr61euh+o3fICJgnuz/0+PBLWRcfjxy+b2ELPg71bYyUIkUWbPMrIU2pZZ6OP
CuXMTKDmKb+zOXe0MaVwH+Sd8c0txdLpLSLlvLyuxw4pShmfPsYITD+axQOU5Izy
lh9BUb+YjOmZBONmXjZEVuyhRFJQUCJPTw3ZSG0x+FKbhI1hG405rPbZ2qPF9iOW
wGtVyG/2af18wYRQLWThNQPYDPZHh/0ky1npeM0BHzKzjNwKomXr8rrbjYxuCaMq
NXoWTbKjTT2aSvyVsjIldz9JkB9j4r8l5qSE60OvZWhzYGrRzzYiULcDA/N5HJIP
9fqqsmOMYzX1PQwdMKY9JTuC21KBbrZDAIFmQ0uXlOfGeV0ebS/kvIDyYk8f5ddz
iHS/Rler5P5bwbvhJjgxUzeJXlqAZ1mY//K1ffli0u114RDOhUKitJk3UY46cO+7
fOf6PZ8UBrPTPi+W1rQyptEuhcyIA9uyYn8JmeLUNfwIRvpBr4gg6OrZTYmYtGyN
I8rGRweal4/QEslnjGY4CNXba/+YJObrd8iyhI/BLt0Ma2U7uiI+OF7yCt3hNNWW
hix+KMt3SkFHrQYygG4v2xJVaytqEo8PwoMr91bxyvMkHgUklPHMxSfWvDcTyyh4
j3/B4an9JwEZJuc9RHq1YHN5f8EpoF6BI3B5v6W/0/v9i09kktAPELoXjHWdNOMd
p5vfZhqTfR4Zmq4z5fcKhi+lRaJpV+HOae4nPy9iUA+auMwkGuDB+dtIm5kegwrW
K1XS4Y1L4KWDViIgkTEAr+jgBg+Ymrx6j95PhBDP1UmcKkkqyr8gVMrezEEWUHqZ
IMdEJtG3jN70GKgKx0PaRdbx5I9tZWys0vr6U6ghGrFSXJNDhRzzc9c4UZ1+rZrn
F1W8ud9jgdnzJHkijWExA0VdSIHlEb5++Kg0EIN42TALn0mZrb/ZyfEfla0SZrL/
YZWaFDVPe+2Hq+jjmp4Rnc0KVOz+Ik8csA8nS95FatgHe345b4PgyKywLUsXnprW
dChahFlG/vjibc7kLCefXwfVNaZtI7Fj9Knc/DaNsXjGJiWFVuerPbRUA1MvHTkw
zhto/JsELGlPZV/nKezljcNLbSXY2c1s6d5WO10pSJhWoyD+rwXp9AnLllS5b/OC
V4QUUZ+DcbJCVJ8L6p13B2s2gQCb0yJ97FuXoPZTZMme413xlxBCwaCreRtmN1Xu
mJX9NCcyuaLBuopREGfoERABKwtN9X+EXDp1WFjjOo6hFpiyeqe3STSboc4GKGRz
1EJUbQhYTHzMlCuHEXaI+yLZ6lhgroGt0LUp5/z3RtrMU7ew8jA9tpl/I1+gtxZv
8vxlMs0vg6GxGrQM0ZAeMIXEBiBhm6Hs+unmjumQMqiWud0mLGHUPnP9cra8EzDk
Era5ol82ekNLztE+esjFg5ZfC5mndHhB8e7e8l2VNfsHlhZBT3m5NaimrCFA2vcQ
2TdJTagjcz3lCxxZYZdYHBKg8dJ2heFhGD4/nXJ93NwN5rLsY52nkaeisCxUhyM8
HQIXO0L/y4bqjyxp8/HdnVeDGPyHUXiqTZ7G/+I7f8UhyXtLeYyGzSKED9JQ2Qbl
vWSJw/niKG+atAbwTUwi9E/tS37Tqeh8hgQkk7nw6pmW/o/h9HfKxylhN4QZsGud
XoLrbEKcGX7dGzL67tuWXgKRVllkr/HLJCFBsTMilX43/DJZ3Hq/hmVK37jnc1ZZ
tmWjC0gnDlt0D5I41sYsktXQbOmW9SZvVM//qKEOjJagV5mF+bfw9VuO4T9H2h/v
kbzvUWnzsce9myG7cIOwsvCkpOzDWNK2Lyw+Udn8mfJc2pAH+zDOLcNNc2Kun/YV
bXmKVdlUNgD59OcWh/c1aUMK/0/dV6DtAp8aAerlm07lIp9OgBHxMi37srLz0puF
y5sv7tmTfzJ7rGbCf+FXxCaYYKMSA+WPIAsQsFzK+S36iMR8ES6rCBbuedTYeXlc
kiDTYhRnFo6XOzuWXPqadn4YSeLOgcCnsHxFY/wgKHxX7B1XdtUpM/xGNE+NbFOF
ZLWblO+MsrkEHi7LTamWg9Yi0NLmQ5gmqZblT/xB2LRr2J1dA/eJrXhFLmFCDt1J
uj3RqnZFNXxsx9UKkZtFG6pTr7oUirMOnmBLuwyWynSbqdMTYx87t9ffCr9bwS4C
HHkCC+iSpccB16F44mC8AOFfrCGIfM9ST1eBiOe+x3GaW4l+Pdc5zkQhGrE0hIkj
z5worDWo4T0lvuALSgwhmHX/HM14Jjl7SA+2Gfq/kpFiTOYhXkVs8SzIQD71eFeD
80IsUPNm7gb3T+ZrI8nG3RYosk9t3TVG6dOHP0x4jNcxCrGhivYNX0ddLbffJir3
foc9zwAFzNPmYSM2CvRTmnkY4vD5w29l/301eTJmSybLqnX9flgUlkVx4ai6QFEN
NKg1ffoYuDEf3LIvqkCPGegi/YYo42Oa4lmkFVIIqSAVMGri0DzGHWr1vpTuVGd0
4FY03QjtooocwZ+jGcdMmJ1yAXQbseXUp+rxSnSy8fLRjGl3SN80fMPVQeaO5Xus
AaDtZSgJi1miD5IPWJcBoX7nIenMqdCGODcBpXHotqb1XLwv5X1ECSkVDPc9x26c
/p4XcoRqUppvkqBqyu4KIXAfniOuGdwUXlYfaCluI2Uieu7nkcfgroMy9plm06LK
KDtdyYSJQFOxOcnoyVas155NGvVEyVo51SrPw8nmOmDP7bvax0FfVhjxh0l2XFRM
uG4SlIOC177O15lvMoAHShq/UEPDzTAIJo+ZNUFlGGjIuEhE+eB7qLMABWCzXAs5
kul9FYQE3EVFnUqn3q8qycTP39gidjukosTe+rQhJHDcaAGuK1Iy13eHDyefpUuw
ah51b32j/lDAjKuLgslzACxaYeXXYLtp91yB7ZQ4EZaTI4uZCEAmYnpGMewI7Ft9
xZiZS6v74OFb7iGQaOsBN78+2mMmCdij4nfrTUV5eAeFB9qGF1kS52P93ERLWr6k
FDo007d59f48d+pY3zNfzDs7vaNgxSEv8R0M6GsMNS0HXDQhUslXL1JNTn10aEEN
PN/7ECC4391AClEXML0SJoqtDa01FS5RrS9IjB06K5/rMd8CsUPMulozQmdN3rEo
Yvw0lg6VajFO9xXZ8F0sLpPpUgvPIEoRNexMmLlIk6pj8qJ3yhW5JJuFn0Ps9MGH
ZykzUigPvjepEYV+NHYPqFxvlCs/P1x1wEToSyXlrKJvfccNiPsEVjkTi5WVM5io
kJkHDh8BwuvpKRxwuUmq5/y6Dtdmqca13wLPtM4kSWytYVIlF9Tw4tHTl9b+EfNr
xUAzqUVRzK9v1ySzzwv3cjFUJ+m9ONSCVJbIvQJJdlrtGCL4+oF2Kp39qgJRTF5F
w77FWIrdpjsKO0ShbQqsdu/6EWZSBTvl/qHmS66+iETMVo0PFBkLHna8YIDVYxx3
8TDhX0w+J6SWQi8TfxbEvFJBVAdpm5YwHJoIq322fCOa6AkFM4VXiP4a7w9fvAL4
bvrG6fevqMtVa/TQQ1Tglxefx2CJMzjg57I+I2vQi0SLNRIYMJa9OhDqaDtqcFOE
e3l0tcVF6SKFEpx0iBfA1TnD1kf4CgT5eqX92VsfN7Jw8KHWMGph4y2ZowKjPLf3
mDafgagWVlerUFlbtKcGCyzqPlsa48Z03b7OPVrPvz635FHZTPcGYJWQ7FaKZZB1
JpF/EJcK2wv90bfXMGRKjpuxqb3YY7YfwUEaq7iYjqRPpBNDT8PeK1OxbrR76KxC
fO/tsre0QCcZtbc1SDZP0HiHhvgdpzGfm8yhftHjvI1ug0FLGdnGX/iBKgU7xTvG
0JHEBuA5C/enzqNyaT5BRS6mC2dUGv8EcilodidOllv3SxEJ5C8Aj4/QUlXfSe0U
73PNlolOtTQdQnA2/A6ocK07dv4Yb9kO4GVqn1qkxTjJuCughixJwhPNxgSow0bP
D52X/N5/CA+HYsloFPRcdpSg0kv6vCubtqs5VWujIgYyXawJEBm7RSlol0Ufinid
4+7dJHRZLw9Qgj3MS4ioHspCXw+WYi5Say+Za5OLeSjDRqk99lN3vfPqZLqP1Xew
ZzGRlTIIU45ItFOnYKM1YTUbdZqo79bu2/ZhAhEwNRXNrtSwstnVSC/ITDOFAdC0
apDrOfSnDJ2IteXdy/jqTFnXD7ih2uGxjZ0tb/f24wKqnk/W7fCFInliPX6sJlmS
7xvryBimpYRDnoVRGXg/9SdxH/HHvYlU0vsGmnqQ32KxqpnWZ8sqi+TjDGCmLIVf
CQ7fQRxW44skH2JTby6VOeONuGF7XYI8hmiLrlx1nSD00GhIBonYY3GE5dRHsS33
r/MJmvuc7Bb+DOGdFn3nAZ5i2gMY5I/CbmjfOHc53SlUb3/AivNap3H7FVo6iyxs
fvlsM8RaQ73S5/cUUH+1UuT7u5suLCco50bbDsyE33LZX5OoFQUgonyzLyVYp74B
lkPSr/FJ1g0dwXkNdEmAxKo6988/o/F7Ek5IGa15kUlpPKTe0q9uKfamVqM31pOt
jzMMEYMqJJp0DkgXuhVIDXVeSZxArctIXdVgpNsZX8DbT/YfM8gjnM8WMVbnhvQC
NKjbg0JySaQQ82EJpHF+792As3RtZZKNCT3OYaoitQLC21dN+J26GkQYqrK+ZD0P
LWIUv1B+/liN5wKE7rVFQCNAwD0QBzg6wMDhvsd/xAMvyXqtglMtUDVwAbg/RWRg
F+ve5WGSy1ADHtN8RZIK1kBbITy2DpwTF2Y7vN8TxW84XwHuM9s3kj07SS+Y2L9/
FeC6ZuBwU+STxwqyiV5QxaGXNXZhazc7nVWzsj8NfqQxQFS4bL1PtHU3BDkMuTN6
rXVXbBwQqeAB4wg9HxwaKqJRbVV79B4kJuDZS60+EaUQXhzIWmP+43qxOV++tSO6
e9Rkh7IWhZNHmQSSB9tzBe5mNoUws2qWMnj2H0hOoibPcu5O7ceNx/I0NrOq1ygj
WmnilrfH0kIdFm71cCPOy/aHHy5/EBmRjulg7/SDAaY4Inmn7HIlckH+7GVr9/Su
UUeNF6RdeU0+eqCADRdoWs3LnGRUGzWYu+e+czsyp+Io9kjDDEXi+rrJEoC7jZlW
C4/UjbXKlbNIpgzNyvK3uCcAgnb2DWs16YgwVVzwJkMKO4ho7dm0ExFGoB1u/kvM
inV5oGqz979UG4+E3ANKJms77Ac+8aNUy7aU8eYgz8DkCRv7C4orVLJUBvn/CG4N
lgV7v+8aQNF8PonBN4aCD+qo/XvZ9VUQ2NfVXpfyxVw0ak5qHJHMjUMD95tXVCB7
2KfDFAUNzVwkze+29+yLmgZGiJu02pZ15LGVp4PsrqbAbQLNGrNk5uF7HlP5/sjF
YZ0Q0uyQHmpmCfUMWGUH96lAz3k5DE0Qp/jP+77wxQbhRuu6pi8l6hanKlQhnry3
eFWK5cV8nXVmwDwPc4iBTTrYfRjrCDgIKSnoXEq6NHp4a3DCNWSEcuLTXFJ3ZFyT
zy9P6d5fmfsd5dP6JnAgYtshhYevvRQQSctdWG2jMiPTcEi/JcWkxl5i7CtIFutA
3J0Rv1qAZgcwFkIAnmYsc6+o0RgFYKfVuxUHkZpDANxpW6HXtEqg5wtNlzvk4e2n
Gd8V6utS6FHQNDJAawVyO5gLRNdhdGM/dXS33Bd1JXJmSQ+qIWV/sstmL5W43Pc/
SoE0RKw5s0lRL8VkUz0NAW5VZ73ZPQdCzV6cBCWNUeP5sBupuFvruG3+XrOyz9jB
vetjaLunOVM24RgquikHfs7zYF+chw2OqZk/6AxsgJtStBv88M7p377zX2BMvAkV
j2Bm+VWYHaIVbrsZV+PuxZuWxAtfYEOvGZj1INgw4QDTC8h2k+krBMcWQMY+QuVs
jLAR8uMvPhlII3ukqOdfhIVHoP2QN89MrUbCH3542drYrIDjcv7AsTk39ojSmB8o
cyzvB9XIftIUx3htI2pSSH95ivA/5ujQIVOeQdU2BKnUwPGgGg+OvG532OLzRln1
YGP+dxAAodg91hIs/vSYTFVdza/Df84XTXFhVH/N/vc9CHXfUKEqAMBH3I0h+4Wu
0TuEf7X6cm7oWmzikj8QZItqIcLG0cCCNKFJPSIVZf53OjRg/mi4LZgHpkvATVOc
pqvhMJ7yfxu9LZjrx/QE6zbYdzZ60QaPimTxi7WlbmpXmJQy4UQ4DO/udz7Shoue
7WuKtQU/l7JWyTgzYxxK9cttXoV+uEBNkcrexnBjXvaH7KHJLTYGSbQHd5U5yv+r
HEzeYR6wCegUNxNO4vqkT/F4TfsgsHMSzJB4phtXkY5GtCOX31HxCG8+BYsvHr2V
6sS5b82J6OCZswPFXmqRH2wh9PFJ3vLjPkou6jttTpsOtJQq0QhV2xloMJRBq9Ze
zNd96/W5mP3MjK3J82IhkFATFa/uP44mlCDWwdy0Nh6evqyCOOZ01w2BHKn00QVc
T2x5S3ZRtvTcoxAyTMLCo08p2Od0AB9tKgLwp+6qTgITp6USv6Rx/XXIBEWSPtMF
ZVbSAW7VylVIC678U6jzi2aj9KsdQQU96zffBYzojKdqG4JV7AJvYdNRDPXV6Q7A
SctY5dfhC1V/1INoKVZj3TPYMGF8wPFfke3bjEP8u5xYzLpZEj4sRgr+9alm/az1
2mZCit39V1xJe0iB/nSaJEjLoEegCktGR9v4bvN7PpsxHqUytD/G21Od8yf8qAf8
VQo/h3VdQ7BP7JuHwD22q+bqeEOBN7rjh6vPzhJlAHCw2VmOCGexobMIBrRfoi93
jKJunYSZxpD6IqyToCwD48gp0Sjv+16RyuPFv0KEGGw1qIg3ZVg8P0z3QeHL9e00
d2AHS4O7uL+j+LUwdANZXtCyc9uffUm6GqsbS/Sh63hOzIiGTG4byXne/IyTM9W/
aubswCuXLqAAuxCdQ9rqxA/5CxAQTK38cDG0V12w8FNjBntYdiaq2aGY18kuaLUh
yRO1yOXdlHv1opgCGlxrheVIapdF54B2rr3rXuyza+QkYc37CItczVZau+YvZBFq
9JvwL8QO70qm+3H1PTyXpBKQSABUgMtw2gTgX8OmsWOoWxRvvSQWPhxGCuvrKPO4
2ndiQjpjBh4UsL6n95ayjjgGBvChd6hPIBQWdxF+N8jySWJyp4azOsxnpf5z/Qf9
sxzsZHp0DEgB+KNCLmvT3n5WsUz7yVVKtJVWOFfxTTWEAWRrpMG38/Q+qBPEQwD1
UoAwMpebSWzX26c5NeZIADQDRnoJ8HJXlF+nQFwWygkV71IipHNDgGpObrhwQz/h
ebQRgbQoFyaxV/wJNh+R2s8K71AYg1P2U9s3YPUOqYDJ3VHYhjFGiwv/NUK0CJCB
pfHKm292BfAJl2vZ5sseBcrmZZIOP7JGQeJtox6dBcNS9o7Jvz65XJyHMyn6rJ+f
7LKepOC5ckqt2s7A/0EyX68ox5OpfyG5ktgHmzy3BrCvKOcVYOi5vfBlcMW0w7KQ
w3B09uzCQuxZ6yftGKQsqasX/5/S5H/AwRvUEU/rims/mkHWlXEu5Rvtz4FSSumd
B/Udo3jN4euh0KPQqV4QzWBw9KVxiqHerhRTP/YP3PatzbILn8CMBaIYRKLoPy2F
4fRVIOSkumO71HDYxbLqFqnxJBOOAfEgYuLsSHpXD2Cm+4B0DYZXhiP4ak43gBse
/S2/pg4KicG9EYou0LN6VlFHm2r9Cn9NsPHt/BJFAceqqxKut5zA33KpjteiB7HB
4i9C0SveoZpABDfolPdxZoPuHZknSiAz8vXNJGf57XzoEAulq6umQYav9utR1KXD
RTl+gvp1Dcf51fQNFxKUXErPLpwE6i2XZMdgv18/k9nJFdtX0u8LnB60KTtv0UQd
59Go16s5kyJeloBSis7J+tOOaVMaepVF3TTPB+xI9tha3Axt+tziECPSKRvR3tAg
nfFMiJy8achoni6zfdNh7uDzmrheoC2SEbKySXm2q6wFjhkKJ2Pbc1EfTN+/yusw
/pTXKRBMi58k4KnpDA2KMhBzk4iVn6dUQORJoDP2dbCUTo8eqjx4x29Nv9zW9DzW
0r++Yql4A87aWbHHxogJepdRQGatGidbkrgvWa9MlumjGSVeD6aDP1PLTMMqk1Ub
5Q7NZw2GI8/X6rmicGZX35ggkK6as4wgpOXxvk4QLKUs6eBe37JvnU7cYBVFllIL
S5InN8ctPOGFf8PWgI2dZefx4By220ccn5H0WV69XcUrqFCUBZtKDIldKnICRGsy
mM8bGN04Qs/VtabTWRhSc8AVbx5V506HiAJCrDYdRLHDoTYK11rZS3zE3r7bGCHg
uM5/e/+ieeR5+Rv7V4BnXJRSGToqf9WgGTQxe+ExT53Dm2xlvbVyrfSbCNDV71gz
OUd9BpXj8+5qeoH898ddCdGHdoVOgwVH84ZJg8DJgUoT9RQwYv4XX45hCNyI7HdG
cKH6NxDZ8+ApwU68eh5XXs0ykc+Xm+CQmNhHfTrOZg+3/6BQ/klFcx9L4H1mZYBK
4zUchPh10gmYDN12WjbIo+uCqXvyCtLJRm7R1dRRl6buNZSYFWopjeUC5z+TV4N6
/BICi5dJjdazuohV2FrsiOwvbxYuBx7HyDti8+iL87eTUP9yBqLgEUjGS/QYzsba
vPvFFYZ2lYe3cGTNSOR7e+PoJ35MAz9wU6OcEE/rcYZonlwf5h89ARagJ872+YCk
gSHpFinjKILMFzOmaGYp5UF1H/Pzv/5Xu42wj+6i2MSocYYecoQgWH18PEYB9Y2z
c5JAa3v7qPcFsu5HIlSF5ykySPay+Wc/vHhfKP4DVP7oBVDPV/ngRIh2MyjhIu3Q
JyBEMCivL6FJ67QDk9DkXScEjfT3J+CGjwCCPfxPO0fov58AvFhS9VQ9dM0PSyjU
4GE4WToGFekl5E6W/x2uedAaD9/RowlCCi3VkBeBFcKoQz7XIU5EAVeiBesCH2T7
AX/M9V2NX/lJYrF4UqyWEmrZJae4FnXs9lOPYLH4tdj0cYX3Rylg7i0a7v6zWUhs
Bu/hmZhtxzj1OW41BkgjgcCUNNA5BDAf/Ou3dz6DeAkEgEa1nos54vHIGyuQZsQZ
VMtoTlEb+t5OBK7jnpS4hxMVisSBtiFjVnSuZB9cuPKcOBWzOrdRJf7+xA6eePmv
V3B+4Z72ZWWk0/u7skEjJQDI4uExxwEt7jrichtKMN4Q81LMrXyDWHPA/C73wgE7
voI9NLGj87RiWTIvKDkFuDUwpG+ZrZ196S0Dvav1WSqm8yy5RRGp/bhH2EAb3FxS
oqaYZFSoONFvrniD+MvWlh1cnfFtE3NZQZ18QmNZ7oJe3arRExATkCyq3g+jXw8E
+AnyOB5VDNhXtRkIvD+YMbLo6IAPccm3CtlcZNtoGyVH/LfszU2ZazCmGiO9CKi8
GYBzwf4IPznY4JIuGSDMGWm5w13xqOn5Z/GBoMJ8wjdGSNv5jQ0hmFR9comH1vxo
PqpRkb1xtr6veWEperD8dexCgOCmVF8+u21lgMtvZ1SmKtOtSeqfXQ3c7azok77b
h4JOTXjXmJsQ6qRpXpCS27HMqk7Cj9vcsY4szlImzaRO/ratiIE5KRg8hEAHEoYN
IfHf5FYNLxWnMKyDYQW8JZ7PJRDd/cav8wCoOKG45JHsdDv4hPkSGIF9IZfIOVhl
bQMvwA/m+k75bXTJa9Gz+BrVg2hivzlh+GU/9B0yUnnsR3etzgQRw2HhKM4QJkNG
BstLopCp97UuOpSTiu6kqWpS6Gl633gKf5oYOssCKEDTA64IwDkzeIQVRs+1vrht
H6whwxBYam5MXsPrEupaMSI/ebahH7Nxk1ZP5+NGWzL9oz+N0rzri6wjbb4928aK
EijPg4pam1+JZTDAWm3vSgcIpMEcp/4kmxeQ09IeUeLydrXccwY7aours1O1D1XB
76NzCmx822g4S/waEAGUUWDyHfIOv/4BXgbJXzhktaLJcSJBZv7K0c0GSoffosc3
qG0Lg3UPWl52ewKa+Fn/09WrwCHHXpAC9V7h+ervWOfqS2vPZmfNuDLZifC7RW28
r77kSR/5YnJdOy7AQlP1LadVpv3hHRqr6dTWCYa22XUMvKyJk+AH1cwWS9DD5wFL
nVScJThMDv5LxRvZBmyafvR4vgX926Gj6o1h7midfkkIH9xR2VU2GgzbAYUNyB4M
a+oT1jUj2cZWe5ZqeJ7m4diPG4Scb8WbCSGUtSXwohrh8n81WpzLjRFO8zm5tOwm
Gctnl9C6DA2MmlRZwFePpW3oKLDrqEJNm5Ds22uPUeUfdga1wnAO0v5uVYgTLXbx
uTWhPnWMlawWvqUIDz+xAj2t5lR/qtAJAM6E7Dq+5pCkmUZgxmEe99xGPJuc5spw
MmFQGKtEJgxLaFpbN3dRUjaAEnWPEmWYJl4UVEMyP4pauX4Y+VJ83uuVILpvAtIm
DBN18afJTw27ezs0HPW576YLwhjbFG3/wHBvy8eWUR5wekHZ6JrWIktjkfx1yeMX
QA6uLdFiyeJtDSOHaoxYpYWI18J/aosaH1JaFu4iLv0b21Er6ms5cMKruHqWxmUE
4Oof0mFxQi7KmnoU/AN4WUSOKXiUU0NZT7wJZVcgxZ7x4BuRkX3kZx2ZcxZ7qQFG
4XujAtNmOqxfQiB15mgIJv/V4ML7OYkWbCRHvWVk3ESvHV0dxOfO72LFSNrXYS1p
xMi7C7cqDQZ9Gn6peBDgp3viWTHF0oVmBbaSoK5ztS+tQdhfW4+hEBZyGsSEIwqX
pal+aIbZrYhXtwd+3rStnz61HPZHZk9BD+mghEzMX6FjH/xl0pZ1K8R6Gp4IpUxt
4JcXqvYDb/V4A5DsUx/ZIUCADjt683wUu+aimBD8wGyJoq35x0qBGBbZoxcCXPqb
yeonXsegI+yxUNVa3BeL20uBkPasHEEHES7wiuNgJrbp/AqhTud1DBJKfNHjBAki
nLDViyIF0LJTZ6oqOPZkYryPVbAIAcXNmZAI5DOEEBKLoPFNBaLJaiZ76SDgmAXF
V0jWC5QpsdjZM2Tv1k9DWnmq3ePu5uvz2j7TREZqE64q87enUP6sPwag31Slt3cb
5+MQ5FuBt7sOfU3fDyEz5MZTfZPN75kS85yxauvVAMt9sfPIPtjwOYtf1HXKHvCn
N+Qcp28U0ObXz4HDNYhPKsm88KHww3x6F5f2OyVIFrKhdPA0T7F9R2+ZqLX/ghZ+
CepeEYmO4GOJYdzvQQKJNTKRdRS0fpBDe2lTPi8OC0Q1rtSnoJNrVrAIEoR7BrpE
XlwNsa7ya7MGPYtP0/9zdn/xUTPlOsi0T0VFP5bDeUPKhKYvjyPl46V1+TbZvdB0
ilT1TPGngljIs6AChV4Fn/x8H4SorkOrTrOeUwPwFXJXeEc0rvpcN5kv+XNBCLj9
mrBoQYLlPsCg1cTgC/qEPlumDTYv+mMKh1U3AeCzdcpshfsuNlKpz/McNk/d6CBG
guUquOjibFocUQoXZHVxQnKQo3vPhYcK2tnweYoJtwWlRO2w1b/09vWJBhfwwHaY
sBAIgPQGzokpiW59mT3Krg7yL4s843VDus2m/tMsyYSlE3uyFRMKf0+GApaacUxT
W71kpH/ShZ1keqV3M7uymPCXKGVegIqo4YRw8W7+ETuJRlxQ2vm3arcBfqYSZay2
tk7E6cZfjKe0QOHfqZF+ori5NldL9PPuazfjQkzMaiveA4JFTPefy5f34gdVNggi
jbrlvFt7wNpjYhwl7b+OK3g8iRd85hWPWZxJQuAof3g1tgup6pOnNBjrVuU21fco
7dJW2VAQjyWr66ZXg0gv24UzNawCO/pVAPu9yuIisr5eQXPMoAg9WVj2eGsqBxpv
RqIhwKQ2wtbudEo8Mfe1crmrKKQzENIL9te1isa6vCflQguu6Vzuh/rTNSd5Eu0N
YKLJ2kqmrQqDCymtb9czV+92tSAh8b1jbnaBBZq9THVPGaND5Z6jJUEQOgqMIgEW
4M9utyBDB7Dm5kyrU0XGQsGmoWtKWGTIZVmjtvtfgUfjc2tjVkc0Fl4QUot/aKz7
RCCnXMyZmzxeX8ZpCwwkxMP880qYJmXUd8F17lddsC0Ko6hbM0zp1FxNbnMsilj1
NwHl++KDTSmpxMFGlSVAn8zHgRJsk9uaeSlYoR+FzZD/XG+rkEDfkLp7aFmnzE7F
VvUw1bLvML+MIEtf4wUWSHdeT/jWCt//vfPi25+zeitmZx3ZUGIHLQFVJ+/ToMik
tEIWoh88vWjDR61oHBCUEiLiKy8tXM/Y6rc5dlIuESO/dkRn+15z/jMtiZq5+/6N
Yhqeo3Z+H+q0+1mmqQ0+m1abNNtWJVVcnDjFNHlxYBvzwrPOKWMPA+Vts/5wFfLb
S8SaUh9DOXT3OFNsIIALcNFx10v6u2O/9iALhyfmkI5jUD8Y3WbrrvUaOlhAI8Wn
l1/41c00qMGDv40TJuYCFxPJIDkWPvj1rL8nq0e9qYKT0b/Z/Bsu/7uKPqvBhK+Y
TF/Ze97zR7EASIXUg/NFj2VTohzRG53L2luKOM4mSvgsF+IO+Rd5t78WTCR77mH2
H6vV0FwrTgBLUhBcJ+77OAdeEYjtsHjhHGKkathskEjE+62YQFIWt0ZGnxOyHzn+
2mCbetLZLOl4EtMarhMfhnvL8J649BiTqqhfXg+m/0sDEHR+R3CBHujcvwoSI24j
iJSPPF3JHmXdLEcL1BA6hX5Z6PxXmiBFt2csGqMxZIRo9Z9gBK2IgkC04k1r1s8Z
GJkQZeP5YPvo/dNEEGSKBFpo35uWQLRtzdrPsn74DFz0mmdgf9A1y/hxUAvMs0YU
ZLzpHd6rnM+kJEHNUdSaR+9tq+lsMWoYVu/I26TKIxC7qYnyi1iYBeyDX1vDyPkX
HVp7rd/hIDh4nEEQ/JmCne5qtWJnbCw11eZBrJtl2qFoX5mre5HGHJXy4diOJ/qw
TtYDRMbZC8uQc3C2ddF3UCzDJmypMBSqc5morU8YYng28YchraBSnrLk9tIVYo8T
gV69DAvXoTu+5qPaS+9wnHOykScgCXbUPgsgyPDAgWPbl+I03hWifJ7kh5QDtXlY
VE1lTJxAU+XWQdvO/bRoD4kx+gRx8fUz+WG56mYJL3uz0iwef1Sjwa9ThIhP0Gxr
DTJ4cwWwdfSdaDRPj+2u0prHkUixEt99wp3VeWNF0hbX0VwjjwhTCdwtz4uuduH3
wDb9z89LAhpDUhDH9bOz0H0oXW/XbwyBlWMxBgMGVmZ8IFTzc/xmsEL5YsGs+s80
IIuPCeoWZz366kauqrj4MN32xcOED0US+8tNItEnwriodE64RFC3FOg8ylDjuVBh
tywVWxg0a0VCgn/7fPZGhiviB5tPGPtGrrqOyyAOAaPyeQvvytiKMCihQgSXKnQq
jXLvsTuScjj6M/jGuO+K88KNF8L2kFVk1TH7sR9zjs2DyJ++yk488fxBt+Ea9nxw
EJw9VBP8FD86dtzjABMX8HJQw07zYMHNgrd/bMW4IcZJh/iHjyIMVUu30E7M3MIr
XmAwPU7mj1HaJ9tA1Dodfp7TaZYDZR1lF4PE42LJu202VB0FkaEQ48vqtOXuinEY
zlIBMlOOvsdRB9RArJ6MY1pkLlgNBw7QbfdMC4tqMSB57B5j1ZMFMmY8a/2XaZMX
jjvmckHbvfJcOKO0HNQ4ZOT0r6r437ei16G4haB1LL8dNZdvct7jC6uMIZ36fXHp
d4CjK4IspDEeehGk07kOVuE/QHcVEIIqe/lLmVz9M658J0siHErWSbrcdxnOXWEg
tRAJwQMdUQWdHIQcKM3+Rk+TVHJtHVRgZ0T3SL0ThP6RbtO0WWjAZFzugQ+1x+z4
Vxw8JLZLwPIA4Y/dGjZQiD6xV0yfuebSRlb8ojK58zE/cPFTKZtBBdPBoOrHTs9k
cLxiO7Fdf14hrf3oA5HOpLQitfJ9kWgEEBkPE+yam7YnjYkIzG3Xk/3nr7AyBqOK
FCjr+BENNNjMpdgWYbk8cC5mWVdF0CzbxC7m2retnIZUtAGSaFtZuyXaT7cF1s95
ci0rV34ViMlNkQs+/eVPaKcGf06EXySoduLDToEyZ5O3/sKNuyMbBN2Wj8+MjMXI
CIoD4UrMFoiJEqvxcYM6WXmUVZO3wQP6W4jS9YEzA4U5bwkNf4zPN7a/+85oQAMx
HodzO0s1dk7Zc7Qj4d8Ay6Jb5bkr1neix5BvCU4OWrbpiXhXBWuC2xwjV/KHeLmJ
Xy6F0VDa0BUPE4/ZPEvZO9PFTA+qJgUwz6I8T+bZgy3RCULbUZm8XTZUysvJ6KQJ
XQqocvP3Q37JgRzj1LQJiBrQ3G9mSpQKuaVYmXeF18S+t46c0WC5Pd/gi2pbEQ2h
Fa/wiTQgEL9AaBqti/a9cfljhR2quTHhLyNrvXHLNUr3IkEaaNeD2CZWW071xVma
I5Q+ogvw3LPYq1Adm1OJYucTVQMooBj1/LVvIMR4itjqzE/yIn6jzbOzm9YyL9Cy
eN+BFq1QYsyuX/gKeuOWvg3lJmaRQ8jLkhS7RnumTZtH0UFBOYx/9I35tRTdBk4G
u1Z0jy4JIN02nKKjECUNw5kKxTEBAfScIWpjCHCLI5zqmr8b4MG0hGNFlpO/9s62
SO68X9Sq9kWc1lIzVxQW6tYAaLQOGtjVLaSBHMzgeodNABprxGdF2YlC+L/nhN7U
ue1CpaRwTifVcFYv6sWHfmYn2KE2DP2K4MDa6qUD/zE6SBWfej2AVnM+NHMedIhJ
Arrykmebr0a0gxPMGi5hJ76Ei+1gnw74/OnXlGBvyDR2DMYGkxXtA7fpFMmEMw6H
3W2+zkk/5xJQmqK3Jwk5RMPWttlgfJgmKNF+L1Rf9bPfzbZeGtbrsGC9YFIa4Uih
DlT9IF50n1T7bvmTryacDni7qL31zAa504bmN6Fzk9jif0S3XSRTqC8hl9l5VeuS
tcm/YptFmGLwa/woOV0ytGz8D0FtQ66fJu0CvyF+3e3wYRg6Tc9iFM32bzwBWh7K
ZSQuJkgooCDl24uMH4COAeCLe9qC5PUetnOaRYaI9/gruPD41sYJyaUDRI612K8w
jzOOq3+IEtslOK9tF1NkOuWsmAdqnTCUNnSXn88QnN1C/ST5dnkD/0Wwoz0Glkte
ofRVX7t0QmSIBEZjX2nFLFUz048Mojes8XgIvBDxMKQWqMjLEIwYDvkTh9z6l9Rz
S6WKN7TTy4Bs/nPbDBXYvInABXl7XnfYBLhM/d1ANkn1ljGRxXBD4EWJt/jZ6VYq
mI19RVEjOCmK8GO/2k77FG9WBK1L42SLkNuUEyhrMzQhG/HYNMMBktXseJ9MjRwS
iWepMKbGIqSUd1WiaDeiDu2nER3Gq5yEbnkoDEXbTb+heTn03HLPUpw5lOfBUwir
rXl8lEdqAXluKfq1SnKhB8BN7ErI8cg3rcoqK9mi3b4wVoYDFfSx86qWRhZucnTH
R6JTAlWrrPoyuiUZjJiRXF7ut6uxaeSZuES10VTr6rPot+1/2gZP36rzt3wItgRa
5peZpZQosSd81b8lYf7oVtu6h64atPsdTuGVrOy10aBd0+WZVOBUoDa+eqSf7GB4
si3uEMJcwyCmxzawTbG5JKc8TOGycnKWXIgXCZfW0aBz2u6K6bEZcLtnPqeQglpq
IxL6ibk22NT8JOBEcP/XnEUDKYZvhkuFUVqMVliHm2TWVYz9h40AypZxZhNUYjv7
XfQPSkux7qs/vGeaBi/YsEXRs4/0DgCofYcdCWM2LsRTMqFpIYHkLD1sYPZRkVII
Uydx7hy3SUDgu/8jr7fCyoWRXJ05VUli5VwCMN8iSO8wqg8EU0aUhJ4l0hFSVFca
nYyb4yAjqT4K2Rbmmnj4DEeJfFNvVB2oCB/EJTfkcixUVhrv+O5VpTDJyQnws2G3
WfDeWS36Q/mkSFfM5sRVBNzvHWtzqomAuFmPkI0O3QBK5hSYT5Q9QKdIbHxXTtt2
hNvrN1lOEV8ON8n+RPjyQH1LDgnOYHZ0G7pHVT6reAKMH0ZbyC6aF437KoTTcBeW
PP74Vs+jyyfm39XrtKWgENkLiN7PQNHvPR/7pS6BjdAenBsjVyhhFD6yEn1v2p5/
jRi00deDN8gVrCnZgEcdY5hoL1tpDVqdxIHeSo3f2z2XnTvDEJZ3KUPkxKoZ7m3B
NLJp6cda9ipGLOIz6SJx323eHc5gJiwiVNyr5ke/dhdkb9jvIaSXPNgh+IojWoAZ
8v9ixwxUnkaaNvX+HpCYy9U1FIJgIG/3jfMqNJsgiQG8Id4Jk5ZsuY7pyUV2CTLH
HCj5c9KuxFP0c74cGxS/XSAI+AJpGnLasxovomvzBNIArbfby5JXdil/ozIYfB4P
D+hcNinukdvh1mORqAy2xs5UrLiPnsNjMi5UUHZvG/bh522jJmpoh4V5ypmSUNkX
FZ+QlJ6EGYjPNZ+f+8s1g/4q1CuDKruu7djWnFHGA5pBU51OqtiF85dswaadoPMH
k8TERPh0tyIUAEx4wdkEqB8ov5DqSalzaK3ZCzR5FR7qXzXw2+9JPG/TgHCl7ShB
BV3Nc/1X8A0wIqjcfKYslQtrdJ7wcIVnog++EsEolczMacnjhnpkLGIbLhAr2D4J
VeLL5BbzJ5YqQTBIU0wVoyMIC+7NKmaV8BLtAcXl5dd3esrr8Dk9l7pwJOru7czM
4Sci6/HnJpnh55+kQhFdCMrVxMvbgxablj5LaPmA4dVgkxZCyP8RrMJpTnjaQX+I
54/vBLUjxs6y5JJUVNwvIZ/BAAqNT1EJE8CZ0O+VcNDDNWp3naZQEj2tUkc4BfNu
SKapB96ZO95xI8tQc7JDuIOttXpLkVl6vm7vjOkzpIswuFQxRG4LNszfNhYPXspc
oqdwkDtMi2mWRGI5VMi8vPvN5cO2sTJF3WlpZpcPGLedBr+s+W8jP5WPB9IkjeVd
K1ePr2mWCW7nmDoMC7XrS5vyTELS8CNbG1lwglvPI0gT9DQcwyOfGq15oqv+vA/g
irSP5GeKGZLMA7EJiLfq/aCjZSDNEjBlmDZHuuCwhumVXrvzKDWFi7le87K0THND
GiSEKFhII3x/5sO4syDZ2FWITkq2lOUrMbup0tvruGB5nDjZneTkMI3ONGTSYBoq
fzkSOLW0Eeap+kmPZfH2br4RukW4W0QkoM03b/4SUBxT5hYP+mkqsDWkbtk7koV4
H9tzP6aeInUmlk7BetXjqhrkntUJfr74lFfuarlX/pzoJnS1I/yRtVRNAgvy0AEQ
y3H/ZI58lHuin8iNtJuk5+wq4DtsHVomfJvisigVosDLHtgvmuSWY5a99LOR217y
0e5YQ2YQ4mWgaqBXIp4b+0cC8fKQeNVxyY/ow1wIaGv1Q5z5bvSgLP8OB434tm/v
tg3bzhMaGsKlSpFq2V21UAIqw53AJRrcIPWcFjaHX62m7qY62X0y6sq/uAs6Sfi8
Y6g301Zgpg/jSUZCxvrjp3jjSFCDNyXX4wnmuDQBgbPJFnFQqzD8f1tRjQB117z+
CTEZNBtoNFTYiB7c84bIfDGdgf7TdVWILhRpgFZe6GgG4Of9BP5eT/nbPsodnUdt
ZVOLJkF8zoLtDE6YSlcTX4aYQOJp1rNtW7GILozD8Ge1UWmym3t3or2hKtuNRbtV
HA6e2oQ0l+3vXpO+qeDyemCTKnTALZFQ2RQlMRHRkxiu/Rak6Fx0HlHlTKJ+s6GO
b1x6G5A6kss3vL27Ob8/7SDq2HMOIKzAaV5y/m7q6AZ4FdMJ3VzWmRqgzhmLI5C+
sDm5fclqI9npJjF5EvuDtOqTTf4P/Z1HZtjldaH4hKm5EV/1GrCpODbDLbqWFIQp
l3c/zUIU+HKBnbXfH3dOOnSSUe4/kC+ASDWUTKGrYbNeJxfxumh+NPaMwwhncWKM
OMw+Q/stwnI+PFZzkmRJeP3veqllky+smLPs2329pCiA8OqveW8qzCFRWjQvQZDh
nETHQ3UWq1X/8fKHix5zMtVeh42t5bYeRg0TrXru0yilZHcQA9b57n2U2EjImSOt
zJjIVNF5SRsY9Lf+KGWTJ0p7elEJAlbPngLGEiJxPGGLP1IZ362upEYs3eIL3+Vc
IroZp0l1kFems1fLJYZ19geBYRXDgzXe+lm8jzWnao0/JkugCwDP+gSsdNX1h2qq
fJ24WJFyNi43eGk3f/GKH9PfLsOSpPjR0R3HW2w+1a+Njt04zuhECGN3C/IZaiwD
ZA1M6fzPPIHW3Ej19CB86x3Ern5h0eH3B/vcq5deeZigmeztyoBH0EXlLhaIFCwF
wca6eMwJrUc0GCgfG5xffp2Oye7EKRSkygGGoHccLAoDjgxoOosRfDRyMVblR5+n
KW6RHgYHL7GvgtwGUckuXH3UvFvtb50G+2X4t52dyHoEqeW8cAyvW6ajTBTAHDIq
Rv49wbBTonqGj7x5q3RLme1tOiSHcuapCvP83Q9gexSlUcduYoT2n3ASRLhv8Lpw
7I3uLKbVV/Ckr/RZjMGHJ+Sb4NR/Y50YUITW2UHgDAsZiv0nP9Mob9dZP+M2B7NG
PXnPAq+1GtWawMWCyBw2InoyqWenWNYwT9C/B5YmRmKJo9yRKoqaImwGRC2JeWef
oFt/yYyq1kPXrWt+wSSURzhrHLiGs2gSXLHWCZqAjvaV7bwLQJnLC9ESnZaKTMNg
kYOcby24tHYOS4AGVEaJWdyU2EWhwALIoAOz+5ZjFMWQ5ZXgRZikg6M9KvVPAh8L
X2arNdyBaW11SkgzFwU8qsslzr0fp56IxJPXpGi0exk=
`protect END_PROTECTED
