`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hD16av00i0xT8G/oCuj7k+frwwmXme0b1DY1pXFQmSs+yoKOEHpQAWLJ2zb8DO1q
bXuOwZWRjpob5abxJ3u0hcEuP/qQ/fvJgTh+CzNtd1O2+MIqJmdGXPhWQ1lvVogr
tqkSCKeMlTHv8SZZ06lpVJgTTh4a5lPJYG+FS+Py4wvIrGKgLd6tCKDLGbvPZE85
lJ5n/l5Ke12BbAS+Snuuj1RGFfN8exVoLtet4KLFVndUQI8KOO8W0H7mjB7fOaVH
8eFqdgyI7SURpyB7wKXGZIBeazqf2DObz27yfjQaZsLRDVbLLXyOtKFoel6+Ql8c
0sw5L8AaiGyoZXTGentVMAOzGrVhK5KHvJzM5E6AG8gzUQVHjrtlDawPMOli065I
5pReTPw3SrLjrtYBAWRQ6vABYwaEg2D54s+qrolHgZpovXKQCrE9QzFS1tE7rpBh
Y64LLKD5h8koE6ZXoxw7cpEYYZAa5WZoz4gkSXNYBlFo1yZA1C+jvxuNUVmZuHe4
756UnljPQUoxrAtvFf0OfDGcJbTQFWmUqqewUzA3rtd5AWiI8TSDj6jHNP0RNwDB
h22vNL7L96vhSxgxRuvL6VPxV6t6U7NPdHuk6/Sp57WxhuDzu9SxkUXRz4LSySyE
wjL6f5fXSE9KuMS0ssdnRIOV5Ceav2gpuYw/KnYZyL3Q+ORQS5jJgDRUdh1ar+9j
OOVNPGLfrvlQRKyLpuhGjpS//3gpNTCI2sYu8NdHFVy6nWmwbOk1zKPHe6kOdR60
HADsFtljwCIsxO9GHv++GqLjJtXqFGrwrBPRf+A8cYyuv/VvbXulXrAndl3SkkjR
eA1r4vcAQb5XEt5U89eoSA==
`protect END_PROTECTED
