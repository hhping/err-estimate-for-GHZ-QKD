`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bNtWlaKnpTKbjUB1QoXZJbZ0FcBij46JOqrI9YpoGfTdbsPhohG9hhM7Yl6nVCtK
tpCuS+4LDyTdtUM+7soO961qbQP42QF8w2GOQTsu531egOZrEqqRF3c4OjSddVCb
RH6pH8BLNq0GmnuGJMmzzW3d1UosabAlYzAi7LgDmIy8x8GSfwuESkxfmsG3f3jm
luuWqsc8Dp7CX7ljqyR5zdc+95zJOGDDzmfcrU4FKmW7GHUqD/Ag0Noo6EFFjiY9
CHsri3y8QvVCj124Ark6GJ5hgAMnRRlOlgQhQHK0WPIbZpRAHBAPyQ8y09Sa2LM9
es6mUagKWzxXNQnF3MV8EvhF4YFtvLgDwwPfG5xgRNEAZUwQFsjxmbvlAqRYNoUr
JtvG7wC2cmhfC+4S8IXQko5D6luNxCq2yIj7GC66ULPyihUneFd/38TKTSFLvZKm
sFkSfCR4GfOHSZ9hg1eaO9LvzZkkzVqHq2noP86H6MIeKmQ0IjIIfVpvt1YUAmTV
llJkbOB9QT6F88chdV4M6c48ran9GBWlx7Q+WuUYs2yHUzwTeMZlEvh+Dk6FuKw/
PTjClmYnEyjB2RrJYS2s1quBRlEMnBN8tcNzF5qEdhFTYQhjJCKAYUkGxksImREl
gxygp1QXlVOjV6yNQKmLVZu9cO/v5HFe0tGAfCyZzX2W16V9ZkmRiUonpMawKzsy
z6Bq0Bb8c7IqueF/n3W/JYukOkpyn1m8ppt5zt/NmyA21NBHUZLlKSUcsyFAierj
l0KOmagbfXDHENYkdMKSFnNKZGIY9dPJ/HcYOvFctt+/7zDYofebCDTFU4+EHF1E
eB7jYBNacOuh5t9OMYsdO6d82+HrvNQToRlKFFaoEAUzDDJU3B+cu/CCoOxey+1y
l5F6LVEbjikxYosb9VHhjU2cMUZm0a3C9rukI+POdIShkIzbq+zHr3XS3yrf4tLS
5W32pwnVTpNmGH87fWtpJHmToiQB97frZVCKpUUcdPIGaKsYaS3jvj52o8G2pqUE
veMJb+1ZlAwjs0nhJW/90nmIDkeOJsD9wxcfyQMm0OqvNmD5IsDcZdAkF8IN57SI
8j6qnxSy/oLjobYrr7DdHb6+uVwhUXSR67v21t4ax4eNpO0jRr0+JzKxUHIssP/i
HkuePKtviWmXyV/tb0/TOxqXOHOpGlgDqkl6zOBQ0w8xwYlfF/OVljk4UclLCC6T
g5im8TE3sHIwXBji7gY+fHlZB2pDJRdTyMZdjYx+TJum6XDfPYGVe3VU5UgL85FT
bwICo32verS3LbCoQ/lR8GOdSMHCArLVYgxyvbLMgcnmAROVSbEUGJMIqVJBooHx
aDkt+1aY6BWCV6a75PHRGW4cYHfSNDrOuM/gfqvbOyf7M7yStFXX1GwR/hG04hYi
viz8KIFVaQLWSVbycqtlNKpI/vBBVB95lLaO0PRSEtiE5YUhM+wNcYbnIHwMKZoa
HnqDUDdX6Zqd/fsckAiSssso/CEh5DyUTqjUyDMcmdZTept+f9+i/yeOmy6A+/39
KmYKWJ5qJddFh3YiGh0i6W98Aw4cjrLEBU7oEbcTUdveDjDgPNcjGwc/VDF5TCI2
4C4qg5Kd36zWs9DRxVDE5YZICphbkBZ8mEKN0LetIwPgqrmTbip/BdpgIcu6o9ek
OXclfhCOTCmK+xSXTJsTbfKXkQDLNjKahOA15KbRYC14TjD0iYZ2dNT+0GtuQuMO
FHiKI/qxB6+9jBUcRd1NwwuCAUjY8z57mKPp5+497hPyst5SlaxybvXJIrUAByyO
1h2aUeMZSSbybbRDq4P+OF6K8BTZfdFxG0meZT2AiS9A9DTRRV1v6wBb8lbUhV3E
K4wRr0UWEs3Qzb+KwkBzcEln2P8iTbLoTROyyPaOOp9qMdoMb5LaC0v3dMccM7Ol
JZk8K18r2NZSfI5bExm2QqwtRHWeenABlF+7Mp+7OCsNIG1SU5WEXT3uyard3v1a
Ve5W9o6nQThLnQGJs141cBTM2f/8ztO0Sj5d3Y5qHRo5mkDSVD3YLE7Ko3N71Do7
ZuACYdIZr/t6jcgqceNpFeuHY9TDaS1oDgAJexFvjUx1iZYFY4e2FO6rk/NPlbJH
g3u1j8I1CJJMrgLU+yIN0QTmJ7vF6YgvcoMKcmcZT6EYPjKJ1EdQtSDZf05xrhaR
KVIZjFDWIKJtAez16+voLMZi1czVjCI5CKQzJq6uI1pA9o3KXem2atv/bZh0q/Su
gBQFpRKqr95Qtf07Y0W2pca7Dn3mGVDo7BTQO2XNQgljhPq8zBANNDlWnTjKdNdt
lsoiXWLCo0NqN6C0hrBUQJjdDO86J5cu1kkrUe7/BogWQW4Bg7cYYidOpD+3hqG8
OocDZiwdQ7tZL8HqhbOH065IAhOGWnOTukqt2b9FVuhN96htoy0XHiD/OrVDYTHa
d4Cifr5szw40e9VfIo7O04jmDm/HCKVZG1wHjCVCMtymodrcOaLQsWLBdtYmBoS1
xj9Bs3vi2tufFPbZ8flO6af374Zfm3EOGBZksg0KXsos9B9IjqoLm3K9UOSgwKnz
sAB8F+IsrW6PnBQq7wRqxugXfvigefYGjbaKs4CqftSnJ1838ziOUZk0BRpZMjae
QXf9sBg6/qg8YeRBsgAXEIhah59YgtwvwnvhoDzh3mnGpmvdZT3pEgzyytEkgDVe
VZUBoNxrpIVQTNtFU9lNebr1aZroOwYpF9wfjotVkKBu2HoDaC1+4RfP166o4wDH
qW35XnAz+L6ep034j5XHSrpD9wafG6rxvhFPlo3UhLrULUeeBYZUvE/GNOaYhcD4
cdV7vmDEf4fB45suLQBnnYLbpJ38EiM40PlTvIflhQz27g6tOCmcBsMOOBAUfGNc
J6cqegD3EFZwXubXO7sUpsAj7wKUZV7esAr/n4rdV4W6f9sYkglRE4k52Df5f3fe
QScxVqasm2TL3EfKXjQubhZGCdJ3rc+gaAkSe2ylgNO+a/5ZqARQgAhggPijO5a2
my87AGZHUO9tNo6n2XZCvgC/88DGLDahUsTAJI6cknnQIRWny8hogGgTRX3mYy5V
ZfwNWA9jsW6q5XaJSmwMzS/7rlK5cToxXeYvEyq9BzEQXhQsBmk2mlSkwiSBNPeq
EYbYRpYh9H+fMZrMcwTnW0ZX5poIMKOIpn18MgAE7YCwLkNbilPMrkf5F1w7LkO7
x3l8JrcWBC/pF4jMRG5DCUDnD+r6VHhHEiox/AP8WvrJnAf45F6Jbd4A4u4arzSj
CrEmpX9sVgTdlmejynHmjRFI3y+s/0n4iN+S3FgwcJLCjRtzv9azkN/v8DtInU9l
0jtyZ5OKWsOEonrfExU4RUSvQ73WZkV+27oTAhbQFuxNq6X3kjk1ohJzgJ3sUlSN
gOdxig9sZkLbfZ67VJQDi5sZRjs+xmxNZRswILn6T9qtVelISuW/ahhDNaQMzDjR
xXirUl5PPEflnP76CNdmm7EpiT3rwFFLfKA18K5MSXY2B4P4u4WsYg1ATqaObB8r
PMwhDQCXFTd4sifiGWdOSjn66qcIr9jZDlwK+YRNuglXmEJKsP6o2MqgEkvmwQ/y
1LcZrXVld+eO6m/Ot7cXRIwk4S9CLvCeFCwdnOXInYKV646ixcL1DZDjoyjFUPTS
3g26dDl+w/Bvjmmh5W5A3I2WhQboLVwBxCTxbXaiqfOWU87ENalY0J2MvlAPBto2
7PnzmxenQtdL10Gt5Um2Vy7j1fyx/HgGnreFqqaSYtymWm4Ohei8sDokO7E7EpCf
npTOD0mjGzzhlDBKeC/5C9dMuBeohzRakgqb23IFiFQ50ELArw7bGm2hv9Q0rZvO
Mt1oLKgnygJ4lJXUvQo+dJTcluQE0MKncYj9au4ddbINzWt5u6EWyniVxfMAyvjs
PAAJQxNzTH81UrkXKdsTq2FdT3CBwh4djXfvUaJ5fFAMRWUgwAPkznCBhb29oyIi
YXTiwaUfeWOvIf4xvm0zj6JpwrSxRZD6Rf3fmw43eTfB6d+b3YiOylvW/0ZtPOd4
GYc8nuAfmv69CLLLvxgOXe+8XPPRBt3m4VlD6QaG1D1jMYC3NNCGbqZWM08cI+f9
e8v3/A9Mn8Bm/GmRgL83Y0laFg9U7ao6YJG9y53wMPbDTgz0IYbyST8m3Mzys4LZ
wKm8toIWaCr0pMuzeCGwwrr32CszgYHrfth+dqV2PV0ii/waWWaoaAE25OhISdB2
E3Juol4Vu4cvE25bc3EuvPhBB3ZCTpldGeEhrQuUQUW2Qli+DfW9vK5WHgi54cVU
vb/HMYNRH2XjHkzlHbJodhpTi5iqozc7YmdOosAY0yPFf4OeTCSmvqx4CD5YY/Vt
uuxiSKlgBBE55nAeeRLEE1+SN6eQrntUiRAmSVVYJLMwuvgxA/HW9o5agiJeGtk/
r/G42HcbZdFKdUIMGWGKUC9XHrLPM2w8RPyg4iDEyrIzF/G5N6HM6+Z/1LddFyom
ixnnu905+n75nQUxyb7szKCN4pT/zP1nlvS34VOYVeJdZTN1tOYukOKS/wLsBvk3
22mpj5lyvjzRSCNWbfkl2pe+y4rhqYC0S1EGL0g1qE18gSUFVO6axgiJhfEHuuMS
O5utAnzCZIvhUlX6eZNO4cCEzP3Py2sWOGth7yDJL0EALQo/T3spVPr4HaROAMcG
LdXZOTMnxFU4UF7ZCCiWkGSyzIDEXuwgSxynqbZhcIinFjZnRrRXMGynKTDAloFq
0UpNxIecicRkmL3ihH7I6XsSXe4fZwE6WVrE1qHRiK4EeC9+tEAttQwilyqHGec5
iAEaQdO6OOosg4fYVLOtQUHXKsbi2IVsxG1WI/tSJ0dCTsEsfR1QOnXVh8FpqHyJ
4bxKfEF7E7henDId+fv6+kfWe8rrs1XP1iRYQnEcy5x/RWFYHVbSZTWsdbSbgU/2
7KxZ4jmRPtbjPslk/5Iy2EM3WmVHFpsHvsygbddr13dYcpYP7lR/mennVpVJs31Y
ZIbr9k/vnjcqsm7l7OkW4J5iiqUh7yP2NT8MaWqBy8uKoVIfVyY0Xjd2tNCusuKb
mPUYBeef/8C6fKDRdHLc1jTRNz0a79LIO9MChUdeeVyctmtYiQoip8Rxz9QhxKP7
FBvJPfP+u3+/lenUOhunoLmpzDwAsC888ArXXhwlBsWUDS2yb3MUbSyQyR/pH1EQ
MLNUYBUNQ/inGdCA+b4AfYzx3wMVdjbTF6tECT7h53JFALAY3BiPgPNd5kqtOjdN
0arNe8ZSM1OOwJiviNGCzwNLfusR5tsyNg9jeexy8b7MJpJ1bN1GmOdMlMTlOvdX
Sld+oOE73LMgS7iAX/SAYcA2s8hohQssvbR7hHUhNnNUmAGrezGDb4Ors+SErwN8
nn6/aAPGAFKADDA3srn0tLTT3x89B6wS+Q6sllBYpI7zsqhC72GU5h1+KcadE9sG
22QqsVp8629tUWoBza8brYhQUzOEFgpP8dysbeJunU67vqlCTOfE+1k5JnJtJZSo
S153oqZgTXlQ7imChrZsodtnUzKJoEiCZwOY9TSlhj6rnd4Iw78/FQZpZUOcxH7f
T1o+JJYjORVRRB/17Q6nD8BonY8vKvGcF4UzDZ5SvxdQ0m3LiHE91nSOTNqbCXVe
zFb1BpnnKIMvifY58l5Vdi3LldD7Sz37v5MW013ZPPQi8fwPmc5yb/tGRsGP+AXU
YTODrDDzXZceZjrlGIlz6/x+K3lsG2iT9bdDU6FcG+mzN7UrTwsS/359/q7P14sZ
JvSIb+adF6qKF/X6nYgJlCmUNulsN9wDZgYuB/Bc4LmeFDkY3Kumun5rE8a2GCjT
SgSocy0fE+hyNkKoQfxG4sec6bxxZN+YqPjJixEKfGrL1wTpr/k5yEFbLkAv4nCG
/0qcc9mVn/zbJ2lYl4ophW4G5AQD9mq6Q7/muiimbQ/BswZySwLCns/fqk54VBiR
hxhDsjz/irbuzPJIEBC8aGhQVjAaNFdjUrbY0QM6wWowMUyhE5Yb8YcQEHpoNDNn
/LSdtxfe475lOHco/T7y4Oao5bHF/sLv9PxweRMLbrnBU+tcB1qC/wS7MwPjh5YQ
z1KvWFgqsa71kWVFLQ3NiebjCGRI0gWZlFg/wK9sb1/PJBsFEXTz322mIcZ+rMqT
G+0IF7KfXc75bL3nYVIDoZuYUr1j2DlZRrpDQ/BII7BG4CCVwk99Dnw7FOaJ8vsk
1FgigwnmW5FqFBcdGyn5M0g1ZpQKApvRTIkGoj92C3nFACExwR6A38ywbu8Ls7FE
y7cvMPaqjvqTsNoE6qDbZx0V98Iu0MSqlAOahd0XbN8NES9l1fHXB4/V/0852YP0
+npZ6voY1Y3c5c6awfVs4O0nkO6y2UZ2baMxRFFwwvs8k2/DmWfLujCBTLLzLuWo
FCSzhTCFaJieqnS5t0DQEHbWfSnhk3pjkjXxZ74FjxM+3wO5LnWIA4PMrahqWeqV
Qhl/A2B7BQeWaSeLWu/FDswSui4CyWQp5KLgL/Gxok81pskAN+YLM+WwyoLZ1BVX
NpdHXFtD6gkWo4h84XsdtvN9py1D6LEoJbk7Lgg/GV0R+OirayOGFKx4ckzUDnfD
lLniPxTlmpmhB62HKQvlsLyPtPJh2lVmX3pLbDuL6wt4gvre0vjdZGIlLMyPB0ye
pMHVmF6KNiJsvzDKAbE5eZN45CJYVaEXwi7243NXiZtJc+t8qLGw0qu9n0TCoUsA
Li9EAppv2+hYiMqgSJxQ0h3ZO8j5V+nfBX+xGFMR36ZLAKOakJ2cBmyoJ3H6hCPB
6cX4zCqLv6Z9NcllbI4odziIjm2IlI7IU1mue/xfdHRCItK2nvZkLDZieICC0BkJ
18cteJ9pLaM4P/cJ5uZwqr2B1Hy7+5Lr7se4CoAAbNeOaejayD66q0pC7YNB0S6P
zE5jfJHjZ3169apsrU6Cu0HEMvHera+ikow9kXr+c9qqZGabRTGjczung7v6gXie
mpj99BFdLdML0YppRkAzVOaWedI0ThRc5cJFrT3/kfFxTcYb1Yow7DHWcA6tJz7C
NkZ5F3E4p1E5DfXSTslQstHBZycxNMTDezOK4mv3nHmDAdT9y0vi8J55nmCTI5eC
Q5eqGsEq0zcwq+AKsJgliIHaFagOvmO5bDWPWaFRp5UHtHrRNE6nZwc46zZrlBqC
zCLGuDxeP/9oKVtpLu/dIs5v2vPXQaCQb3dDcTLjUSOvNyJ5CusGjXVi5MGD3bVD
Ru3LyntZ/tHil8Gk003gxSLyPeVhhK3TAGrEgyncq/DUvfAGe113foyOWg7RN8aE
/4EcuZ/XgsmOzZ3/VTWHKzVFFHqsbXm5bDZYONPzTeA/oTWKKkKoalV4eohnQouJ
mnHmKY9bhKAHtU97QTK2oVmVaGxPd65vNPizVlEakBEqAX0Kg/8MSh0x/QTalj5t
hRgNahnQgVExgAMt1rCjthpgZthbSDrf4HfZBwFc/a9lGxcEwW9t8WXwtI9EnRPm
eG6+rwx2oQeXdnW869STjmKHFOM5wzJ9UUwO2thl+4M5AX7S0Cuq6oJAAYjE3cc8
46Gskr6YdahlVCE5pg9P5o0dwUPSSri+/rpCkz836ExHHZGV7nwky6yJGd8nb/MC
VmZAZQacUmRX928k32pVMzkCHPxRB02WRrGJWGZC5DWVLuH0XJktUFJM6/ojSwR5
o1dW8l0P+ivTtbBWfZmqi4rRwmjl1VxWaMzIIec+YQtObO2OgVXptbdzDDaM+GKG
g67DK877WgM4NfdBIaIjIEQWKFoXdD2jHybDGgyWXIHYyNCUagQDyGj8spG714AY
9lMF9aGi6XZzu0RQuReY4RMqqip40OMHokIWKJL1k5RvIczBL6Khgo/q1ylCPBYG
jGxWGV7MwCp2W5pkvJIi180sdqE1dhArqatgkpXAFoPFyWNBBoqSaSUt6zSe/nHR
9K+V+5gbFf7dqKcAXSZ8GLlEziykjH9oa1s+Gp8ptsmT9pBC8YIXnJ2iBnoh+Htj
mHlwMOyAnxd9WCjHsbvA3OoQKbpUNzgjixr7HbJb8hVWarM21ClW8TbUSBfRc3Yt
13n3BCTh3iAQRpKWqVuXXJbMR4HwPJ2lfmuwxi4dpZTSeJorQU82JfCuY7Zs9lV+
ZSx+cg2x8FY5/KA01wLnIRasweuSKRkc0pr5O/yhWcgxWpcQI0tgV90IBcMlY5nY
WexLgxWO29xvv64xLfQQojDgnKr27r5ohM/1S9E1XjJSbEHx0Fy1u+fSuqZQpK1k
yXQc7vFS3DvEuNIjpuK2KoGeBz+gStdKNU7rBlB+Xho1lxEOehH+5nhEdU0bNw3P
hgOWK+ukJXR7piiD5PYoL2kugcxIfEUAi/E6W6RxQTN7X+3nYjzDk6PZ3hQZ55qX
82RmnYDWXlx3F2PfHxCEc0L+5M3HfYfq1xaHaPjkP773N9rpetGYHJ8yXH5hfN4w
v8LqOWGfiZsu4JQhAFGfDUZhZBFrnwQ+2bzXLdVkB97fLERIBy6RjkwWReCYSZGy
onZ4XTXCj9/zRjlyzkJcfVAjm2MrEshfd9ktg8oIUm7FWuXU2bxUBif+xuMIScA3
X05dXKApK7OTx9ElihZjoq9k87m632AvpsuO9QSnOudQJJPMS/ELnjobXdXe+ouL
RLYce1n27RbdsZeq5xpGUruCARBgldseJWDeY85YFX/BcVbxaciHJv8TxwgY7V9C
oO/h2mmNoXXUfd9VBtrH12GvW43BSmRnT/V/S4HrFJbUV6iMH+BzMZyMFi9aVqsm
W1HXmflKNFGaKBOw51EgRyclv8W1QWMChQhojh6aqHdHVbW+RIu2PTFXWAyyDGkm
SP5ceO4kR98SugpyQsd7JzBLsH/gxhFi9NqQlUHEEeB8R6unswzZXw53mKa5P8F1
KWBMhQ6fNsQMDFMKV5uN6/yauaZK7J51tRLvp7Bo0gs6hC5iXsJhymD3qQ66hTYL
BkCm1njRDDqomRv7I6xsX6TeEp7hyIBDRmE1KFWi+V1DgP6phL66B4b7zNZKrE17
fd93snFKiDiTHGgfeUQFAyVljMz1GmiyYucqKBbVsRA4oR7jgH5qr57eBHXxWyaV
rDtLcr3e6KVh7uMHaf80a6pdTTApUAgsuMVEd5EYCsmmFc6eoDAV5LKwAWQSNV8U
uV0+XizM/IoLipheJHX/P92EPWnDGED9hi7uqoQxf4yuwCee3CU5ltuwIgPnSqE3
unvjugLzVB1avDJ+wxIutCBLqKc6KvVqwzIYOcJEXu1svlYukr8LAE+guO15vcnX
5j+fUY8bx9XNwhlzvZWZxoRfc4vk5XPRtaGLOO5Nu6/OdmQWFvVZoFXVpLJAKtRB
pXehiitwUz3ZUMrUHSQW73Wfgrwqt7WdCY7yeE8HMyHF1veehF59bzgkQdrliHKc
aIYx+XXlhTg9T3gKhkR7dj3IE14AOKnvtA2gEfq4cKFynsSm6eUldpmsdNnudB6b
z9gGU7/vV1+olbfvfH2MTVgtRfleDh1eXQOMM28aAhi2V6STBCtRZSuidK1AIin4
uZuj9df1vegHaztIizIrjYLgKh9s33biyEYveszyZj3N5Yzf8CSvvuPUF4EJiU3K
vjXjfJBEjEpNFboF2c1Ac/y3NAwpMcP/X05IOska36CL2Gm6Es0djqxVdwxTn5jM
dn8TqojjnsePuA0n9Qn4NxlJO0H5hUEAE9ZNMVg/DnfIjV3+k9rE0iAMLAKzpGcS
kHZ399LKT/xeSM8ABV45solkOmAjRreLWTwhvIQBI8pFJRfxJr3KPEddnFKyW1o3
1AqaTPajWZI49wsY8gWov8dheAeJUc+XsLmiV+3Me9wNNnh+66JBgAk0G+lvVawH
i1fE0iCNeb9BKXixA+kd3ZLhJZ8idaV/W0ppRcxhrYZ2yDdBLQj2zAl5Fj6Rb1TW
iEGptrJi2AwRg6zYPthWZhpPv1EhbSZvu5z2nEWEQdp6ARaN49t7yyNW1T/HVkcT
5Q42w0aCS7dO9Q4XGreoS9aQIEuLraKe4UuZbs0YlK+G35eqdG9yai0wNxufte8G
LMoOQLSPxzIlAuQxmg6RxIx5HbjTE2yzZgqQjBJEHLN4ygi/Em+lJDk1zR2FkCjQ
97Y2OAxlc8e5VxhPcbTl41w9ztTxGrzsn5FmaTX9dmJhM+WV8PAXAAzF0OEGkLkT
EGIbO69us5K3dK0klQ1WKblyLgeYiQVlug7meSVLg/pJXv65+iHrl2xnJ2kV/vkz
zhpEam2Igyt9fN6pAc+rCHZhbI34tFrCbqDEj+xiCokbsXhA0MWsFRNulvOA05+y
d7Hb7eZSvKFQw+uXpOj1+g1O1sjjcIVbX0r+JSm8vtyENtjzqYXyIbo4z/m7Fj9u
MotsXhUZ5II/QdMdjwFWP9AWnh8Pq26b/bF6ezQw0CJGsTN/9V2QUjLnwvxOaqp5
UT2Ff7dq+TnAIYq/9uTp3/Oj3KeCTcvUytOH1OgyXE4cfVTiGrsulk12LelRhOUy
GaCMFs5IlbCmq8OhmDXjwsiFIja6V85Ai+g596/MnKQgjbnbdJBwLOD2NCYyBQ4I
xtSap2FDBVVE2QvwUbHXO7vk0BtiNikxxeCcegcUJ1JSDEM40zY0v3/+Pr1AcpCX
YKdVP0VS1o5tv7hydr12i6C6jflm8dkX0TMh7K3CY8F6WejmUoirpboucrUYLSEw
W6RVnoeIubJv43ykG5ygslZx+90vf5wH0XuUm9qxO4wxdlbXRzkHgHtErjm8+DGE
MdAv+gDPeGT8hlTMJ2hO+q6bFxyQHSVXLey73idU/TIi5bL9gJ2dDg5FhUim4Bvd
C1GYKRmEvhBOTFdNjZptbc/lm8237idm2pNl/LqYDbv7EAmHYede2uba8slFqk+I
nwF2P/Rpe5HMJiky4cJZo90PR3F+yZ5OZIpR7r+Clm49t68ga5fI7Gm6wHIpqyRQ
39H0ujbKgXMRylI/8W03H/oR56gzpsRGL3Qw34ymPViJ3hCpGCWqOxISJaZuJD2x
QizoccxTQWAQ25DK+PKe6zi3ex6P5dlkn/UMgFLOkGTqYCjzlrILhyb0VFThWJgk
gZTwB0Zqk6pM90KX15hin0EMeRjALdoy1IeNqtLxuxfIyMgK4TpH5Fdd5r/Sl3MS
5Q23huvjPVHmhgSBVrP+kyiRLK6/vjz0vQ8W9TI5DwPGK/3H9gh8r2ZTmwIj+Lel
AdzRq6zGVPKONEIT60psbIqh919ImEnGFZYaZD4cwsM4dhoVo6PBCvlq1KJ4Zvh/
1pzBZ6v8j+Kdxhfj1BocmvCLj5xlmH+W8k5VKedGpsj81ARsrWYiQE8Ui+l085PZ
Oqf9NGjTolR9A7ByTyNTgCZNMNEd2MT4OqmYgIsq97DxTrVcMmI5vcjmCXIU0/ki
XI3D9XOXb9MDj77+FT89j1LIXj+qVka1OiXAgMbikFiA5vZE0DmpmwS80ZdcEKN1
ccntvd9ng6lQgJyjBAUFzn3t3tRsiV7rvRmqRYm7xWbQODlNT/ChQ85Sm6CIb6fV
8XBwHj3hufSbH50yo3OoXPqErYjN/rFuttcUyuU51NmfqMLLKFqC9K3W9gOftAmK
8fdcyulKU+1dXs1M6nLXIjLCb+NYRL0p9fw6lGCIwTT+njSN+th9MUyTBf7OfN2w
0U72MFOlJa+Pfxrgqc+Ce1A4EQk/KuoitsSccTO7DsAQPfgU3Cwd/i6FqNheG0UL
+oDVWfQIQN9OWJiIz2U11404JmmHWWXLUc7KmDWRIIrxjOWewSVfH4IPfPF3auxu
oITO77pRbrPymwumOAmWvuSDJpW0kGolORJ9p51hyq3AXS1sbyE+owblC4enIMdl
ohcRI9kn45vr3o/cWFLKsrAeg4yf9ZhVQk+b8ijvW9bIyuUBAJr9S63QqsgIwzJQ
49P9AP+8CUyOosuQms4+YxvlwrV19te8dixiQuewK4FGSUIdgT2pCkQ41D22xlEo
aE27Vm0pWBeKnIG8bDdUgXxQvmry6atKO2KnUw1iBcyRw7MAYAL/iM+cCBiT/CFd
ZzSpATG5u+N+I34xZ5XTqyplBEq3euaG1w9JHGYaoLByYEJsBVsaQJ/siSh+2Fpl
hAMQIXnVpcO4Dwz133FGfkoTk786csQZ1xl2uN9CYcZxmSw3Dk8nY9mupSIz9FB+
X4owK+D6WEtsBlHKQYOtjW5IJUPIXkeHQnBKR37vAiONkTWNSqVorRj+K77HVp+7
uRYC6I/bOmKK+FaGJIxUaKomIt8/1qVSqcgfW3xO7+xcbPfTIi0yF5QRsXebrijc
mf4Eg93/LW2LHp/TkE+lDlCWWknJJ0+1E26lPZVTNlP3Mr3kU0nuyMlC0z7ki2q3
tJIF383VdlAYoScs6HPRcCZ7ALWWET9xPX6kKIS82yEudSwy/bpzuN1nMOU8lGju
6OAr4a8FwFQenICvHqKsA3lT2KGFshxmcdc5DQAZwmVaeNibLL2Sg0NYGTpXLR0f
bq536+23OSSG1rkrH2907BKVOmvUVqFWiJKIBLyEW9B+sn6ff1nncQcuMhS6wm27
QqJkeHTKo9nnjrAj2olpshSej1qwK1IRo2U/8FwNIpKQKLexCbmpiJ4PNQnvmB/7
pu3t7+2xqagJITEFlZE7oj5x122+J5mMdo95+1D8O0lsnovoflObT1aA6DGF9qkO
otF+E/I3zB92buT0cTiehd2N2akt7WCJhaDGym/77r021U3i5FzkDDywvqbJaybc
mPRkBcnGUyaRATnj5+pudmkheLL+RAWV39su709wIqZ/V72Bg0olRw91v679+NNM
bM98u5E97/IGNMeN9Uhj9AwLI/kuXd70P3psUr4GI9UTTEGyfO4GHt7UV1oVu2L0
Ev7bYCKofnlqPTvUstLJz8LjboFIyXefGaWby8K1U+FFTuPsT7WB7neI+9qMdUnA
txigUICXCZAjVZ2gqyq7soRv6akLi9/xAoqzp0SZrKuGGO1xb2NUnpz8DcIbNm9W
0unNjEDt/RvyLvZzZa3/FARpiumNkA8vthp/t1hB06mSKvkoy9UvGb7BuBRZqwjV
ltR8jR2tCsY3YLtH5ju7pBqsiWh1G8M0AdRpF52AlWWkOmgelKsok8GdabqA78K0
3f8C8VpRO+1qus4zAcZAf0IvKxHWjWC+wXlLoYMLkT/qauTcjyTH/tef16KfeI/2
NKBgzA9cxxl7U/2DGE/pn+aGKDuNM0VnWQh01Ufr9ACTf/RbEa7Rp1AzwxTAaJ90
Q0wtZTps2IxNy2Mz64N8g29a17pYUIekPkn4fuXSpWepZslKvdxa8GLLPeD3ZcYp
MEkKi+Kr/oaOReM0VRnLiG89FRNX9NL2XW2Q9v9GZ8dblCbNN/VnpC3JpOiv+1vA
MTq0T5RGiPHvYIcoJGyMGzn+HeyW3MQ5W0RnVODP9iXFRQATH7J/OwAkvXcOL9Do
ZyyzlRZ7ZY1189pWiqUXJ34i3H+ePrchytzlVSpr7Qb4o83p++kdTT8oAIEXXgWm
7bWGSR6y++Txg8dzX8CsbqRqSY6q8KFqvO+20qqgimzrR3gFZfbP/4QIGT6rWwDW
Zg4DMIMnICk0Q58NuL42XYBrzEnrReTnrVaRRw/BukOaD1Lw+mu8v6sCPpF6NH3I
EU8SIkXWFJoE2vCRnlf7muOYkY3TKfo5dXbMWdouYScCIEEDAxPqS3cBTJDqnGAR
OefMhy9uiDMyVpIaJ+MGAyS+t+6nEemudrKUjjvMorb3qspyYuoPj+abwYYzOwLJ
GIa2V3j0p2xn8pJHemFJ9IMz+7VkReL3vnsl4lXymvYMsjjhKw23sBe96AiZF359
jcF+78k77/Lj7L9cwrwJ6silTexaxKzuqtHVgLLryUHRRdvjR17vd1hxBP5RXK6P
wmvt1kJK1GimzS2yKzSCkLhY/MQhCghMafggqvJmTR2bsGRsdtTdSmvIb/XwXgsp
fZ8nGJUw+Z3PoypUG+7Gx2GQGiaCm5YCE92NWEiGKlcni3SkWvUx5nmwAS97oQjy
awkhDQEMwpHmeL3I/kUoampD/Qxlc2sMer3YF05ektEpz2JU8j/dMCRAtiTo9H4M
6PPGahAgSkj4CWAMhEuK2ZhzKQvKXEqVKnrcVDa0DX6KIHoP0zqWWMUmoxy4Qaee
Ar8tNdZQtOJV4dnEfGM9xpcJ/2kKg22IDsPKHBThOVZezAPx2F8as21iPo02rx+Z
H5mTfoHT1mAXIgdXX3qlD1RxYzvPXvPR93yFMFy0Qc0rkv7W2TefnHkzLErZxDZx
hKO88n2wbwIpO8pk0vf8oSyJEeyScQ5Y+IKmlhaTin6bKM0ipPU/bi/afVwC/2gK
FRaNqt29nR/HJkIXmbEz2ognirwcTLbpCbf2r3vm/eIK/2dPQ6IspQNfc+fyJ6lD
S1IBIJILpbmcJz7mSxfR4QeoTwjePhSyDIDcQjeTGtte/8CkM4L85yXfnO9yKI/e
P1g5DaDU3Ri0YVVU0XAaU2ssVagN8NXIDFhZKSCcxJs6oZmpW9DWSyga/xjrZld7
W0d0GMG/g4H5rhZXEBMG0b0fgUf11jSxOfZmV2zo4sqOcRS9CE7tIHPJqSljE1TV
P1z3BwsArUD12MWQ5Ud+Z9VUgdo+HN+V7AEs9t7gMOHlkfUjTr5cLaNnKxBmgvzT
PaZevD1EiByIFsWsCuGfKlkZPPAa2ysJufjelXlb8GoHGsjps9m+BFBjXiwnwVKN
GUgMJlAHPd6mHrHajJZ6mVyetDMLAIg1gX66Egw8jk4XZq/DSe/WEwJWYqdMAGSq
017seyJoeTTyha09FAmn0MxoJ3REIstkaV0fjxBJacAZNwoeKn6FdcHGBQJJaP5T
Ty/YxDhoaAtr2OD1LoNML7N6QkNqrccFVYO50gZzmXWFZ0b5gcUNZoGypZ5CIaGp
/bE8d1Eri8gfxrym0sbIDKDizrgL1X6xGFxvuILh2i3FYkw9HEcnz0DwJkFyxbyi
TIWX76miQIaw2hbIRa0kK3KV0u1fDXRlr1iaE4zY8zpKUyTRXauiZYrJYy/eZCfM
A3Z7+NOG2twP7mu16vZvQJ/X4jIU2a+4WlHBkWI6tb4ii872crxwb5WX4uI+2/dV
AFXTzb966iRzU1B5yJ+CnCJ4/XPqRzvwxlUucdEboSVn6xuHuXliiIddYmScg47S
9MjSS7f0AGiD8N5u+OrTiS28jaNGH+Cmets7fkYZkT+3be6M8PZJQZogJvpktb0k
wFG38xqZUvooJS1Fa65DXamEQZYPAov/jiP6A1yFHBQAGv4n8QW174LebMo/lTiO
YBhAER5UEzRNp9sOyKyzqhOfEIwFtNCagFZBT40B7165aQIVfbD+QObtjWpfd2UC
OaoD5qHmIdNflHHSuSYOeBFEQoI+whuFwN3BXDEqmYHsXjG0BjGk0kulJB5wzW08
uIBft0QLjAAk4/zlS24ldDNz4/TW/UG6czlhmTT87dNGHLEKsrjJQhqQLW4NWRAu
NI5ZAtD2mCbRX7z625Yo35jHxrxRW4XxegxSXHb95/CADYN+rNMyYAewcpJS90hz
rmPs9VThyOUBfDIa9XFJcufS77E1eqEy54r/O6fzHQeSAuyUuk4h3w/O5AVw6IYQ
+RmhP/EHDaDKofM8SLWmD61QYtD79sxwvKxjnvMIMHMHLDC7SPyvXKxnZMWRlxEM
xppWnGcKGg4crrLW+K1BaY+Iy5Yc0G1KYaMjgrSBzY/Mr6sXbEP7cqJoJr9/bD+4
AH5HIsvw57ZkmZjzdU4+TWlJqXllQmVMgNNeeX2BaR+zn7ECTFXNJWjB6utwJ4Hx
16vn2T3N5wyzwnljZhhcOMMxDQikDqTr2pjydY3+0V2L8pQj/Yuj8Wb6n7bDjRzs
2uUD0QfK1AEvFVDQg1ElUSmPewgXCIChyRDxxWGZx7i3towreghyv83BNjfBQcDr
Tn2cbHX4AB0wHKkMANJCfGpUTQCooDgbBA13/dJgc+F6CJgJr4LozftS5DZTFdMX
+zqOwfSE31btqxrfstV2wdAye/mrmNEMnQvIE9YSNQUOYtA+Qlw7X3MMvRp/vPvI
11WCnatXWfulzysr9IAoa5ZiBkOGBWCkjtqYPqmfsQ5VXiBhT1IzcdIW/gLxy7EJ
YWKzOelBejouw6hfkuBuArPE8xaB3NJEtTaIJkZvCHdaQ7OV9Igp5zrFygeJobv9
yX1M8Hmk88VSuMupdxuF7WbRc7DELQNu2d3eFkZ9vJ2MWmCkfUlqijzzwHJOgmTm
Lp60YUQZs0XAbpebMjGbvvGfdT/pcTeT0asG7HkUOgDNPbjKIxmjYoZAYr/Tztc1
DTyhwpBCQz7d5kFnYjVkPXWViY3CFhVMDIHQ6qeKJbM7sqHvH2Y5VN0fmvbkzbp+
QFqL3ByRXSEky9JayEe2LQmwXEWu5MjrgrNjhrxeKzl4KWd9Ue5qaq1ikanidrBp
6lrIWWLa69p7lJbZ0FUaT0X36H8Z8tvT3UO4RxHecrCqZdjE3InFgi9fn78S3GHa
mUe69hERsjMZPIKXkJiekkbEBfamPOehBRyNwEKFDOXyP4w3PzAnoOR9k0Me0Z6F
q3PnzIXM4duV1z9MZo3Q+nexex8Z983GiDG2Ow8eyQhqAQqTu3WzyugH7dxYxTC7
5swD+aTP11pJ/yeV8wFp9mIvVBDKSK0oEO7YDiGu8T4A8wgHtSONinPfn9Krc8ku
4m48YlTXiEuDziRAyA5cbT53obJXIRe4L/V9CnVZ31ddSSaHXdMbdoH1ahm1Zw9G
1l+/lcioiXxs2FPHIJSiicCLAaB1CVeO3yULE0FZEK2y52L9UeBP/cipNGSnCZk9
iUKh90G15dKGa893Nf2WB/M+4K5NRgvzkOOXSiiDm/DrRq2csTLNFcwnAiyhMlyP
RVHm23y36iYKRP3lPSPTk3HnG4eP0zdW6t/aDZvEqa13OhF11wnxUr1efmKmh6y1
U9f3AQeA3G5QX9FJIKIUvu57LycmRvfRO3zL4iB9TfWqq8hD4jjQZEMKYUd0N2rJ
IRuBNkmz44fQZwIYMuNB+utM8t/g/yoRFbI551JxMjfZvibdV4BIb6nQ9OVvmDg3
Za1gGHO73PZ7BCQzVG7DJR8ycAWrL9Fr8CnLX5Ccc9thYpZaXmSd6E3YDj3COVPg
rRuZKSWecH3koiw8/UZy7xS2Q/VjAV3XRP285wwlS0aEWwXz5bdBeWvr6cRACWzn
VcEo0i60fRngZL/X0r4VyAK/UFHLAYkqV5OqtHbLA2KmlLLcnq3X9iXnFttqo19P
TFChdPYKagm7ahtu2m98YApElY/1d/DZdG9hXYil//aFQylr+9l4OA1XxgbooTh3
yMHZvMykKag1GygSAf9LQoYVjIEgNbtWDgKNecCR4b9pVU9XTd0IRpYAfFZP5AS2
5iYjxH9R9z0ftXWfVth6L0qMV3sAoilg5VA2WzpsZl2OLwGGWG6q6HJD49KOIIFD
VGrq0Sj0Iwu3+j5vofvRTzjyUoOn7U+1THE34Sv33GiZCOmFIcxZzvraATm6BekM
RRM8baYOQPuthMDZBlDGe2sSBzqlfmfot2g56pA9v8XCi24A//BlltJINkhDfTSD
xwrw1xQm47ZZSKTE7jEc9lvKTIGJ5VZjJOpvpwRKbiYfu5PrAOoUMUNCDq/XhskF
QSMfkT+8ZH8KFN1rgnbgnoNqe2b9N1n/kqe1hxEv1cTdi9sbjCM0oVNRADU423nI
Mweu04dzKumDgYCgHMUGIlFP2YGjOYwthCw9sBRlsntgeDN5JWA3MnbecA3qybKY
lv+htpwsbhSFrPjzRL62/ULNPKezcTnt+WP/6a0ztRoo1tI/dtzJqh67jzvHKANN
3gZDF2piLMdn7Z485xDZKzQveTs5FCsw6h/u5pPtfKJLObOuJZbmxtErfjm/V9ry
Z9Xl0mvcM+hBuSPbfmnT+2p1NzQBjxhXeop9zLyEJfMjvSpUZx/8/kHN+7d/DSZO
ybPfSH9H/nFYDNbjqxZooosQHpVXOJmEmVr3NX7VeYpnSMNMopDS1r8EBuf3pKk7
8+jn26uEg5Kq8J8iiw/FgClbrRvLWVN4SHR077KcykOhW/buzUYfPUM3kbFKr4oR
/Yctf5ELWfvhKkTiZh7R6O7KPOwW7Vhr2LmrEnxEsKqV30TTK8RfngLyTEXZBYAY
cAQ02eMSKyhedStWypGVcZ6v+FO6+vlbdkPDSJVFBHFYgS4LBIHbDnKKMrLlwZ4g
3Aoj7Uh09NSM5L+RPvu6V2P6e8iPpcWm+0PbqnK1q1orNdywNeuxRLwXu65XlpBh
rfONsTH8OAjCXsMgGwg2ZMdnkdwAz24AsXr3Ok1bynNbtDyCiwEqvpIvhS4vBwl8
49Zf8AAj07rPybVC95cgBe935To/9Ufdg6s0s//yrfZzZzrvVWENn+8KfQJ4iZXF
qzdp9yvMVk8/Y4I09943fwTMnCIHXeE7zZoHI9pZ04u1VR7iYizwzRLGUtMsSjaM
ffDZ0C9BHkSoNqYPiRPYAFbA4yz6kUosxKnCMjVUilctaBNZkZb0v0tmUanwMZmB
6rFBZDFh8KWz5RAXDlR9fvFFCD/xAInEG6tFZQC3L7nWpfYEuf/dF67wuK+N0gTz
N5+Uw5pTZVMSIY/Yv/D0DppdCx+b5IugEvpJ1qGICti8IuBweosNGnlp1+lVdJ+B
0YEAkH4aRRd3SeqJqG6QfsDuRp6seGpI+TJUaIYKRHHO78D0CJ4pO9M/8OdSm/HN
eBqLdwYrRTqCYZtk8QgdX+Q4NfX6g6BQbZBuldKcOntBRqtkmVjEgEBdQGHXoohr
YfuE9QYBNIeG9Pv7czloB9Jk3zpaPJQrgymnHE2GsM2KX5cuHxx9b3V0xVjUCdek
/xuEUfykB6uHwFvKwhRJpkH3QdCxoJf+spZA040hD3cvKQx7VxGKtmLFwYxySx53
mT08Mfkp5QTHNwZ8que8lmW7Kf9vRceogTUf09mGAVBkNi0GVmOUkBRlV30gGf4o
1sNw174Aqq/H4sMz3sCy4PRrLM3Oev2Uy1S+RIz9EGK4sGUvglKpTSPbs7sSJkNr
E1/UKEtHhgCjxQWhDvxchbV4fUeOMI0cyLVxO4A2I7dZFVDAmBm/bSQwlxaz1DhR
y6KpnlMNX7FA5vgXTwOexpsU+hI4l1aaKRTQ4y7SOXs7NbNeuS7XkGWy6Zx3UXI4
4p/hgnPqH3kednpkg+eJpkul7/OLpZIKwryMjS47wMQ3DUlQnG44MXt6Z3ug2yQv
g2x2lgysWg6YodwYIMh00V850z2rFk0/8bW1do1ZTv2hYBT9BXkx/EQOaI3/dJ1b
qL24Wv4vl6n36JyvY5k9iOnwQFcgcAA2IQNaT4cgSR3Re4iNTkgwde7hwdVbtnQS
k8aAsF7ZxLNKIbi5hENwiJxzXwS/TLyogOVEht13q2d/yrSGH5mQynj0NwuKk8Lh
QqFLhqfC0Dii808Tx4buEZavL15TG7gMnZQl1iqxiVmgOKPTb4Y0keWSMmx3/Pd4
iGvOBjb9xp9wmfQs4um3U5KlnfLILk6ahUfMLktCHNjuDc+W0NTx8vpbM8nGAR2A
z575p05BdzjKyVsnR3ze0ltvK2vANn188SEyRpiRBf/kg4afVSR8M/jrjrK/bi/a
4irmKD28YY/PLa6Fe+b23RiN5F4Sv61myu4c7/454eE1BSYKKRzh+Eqdsop5Cmoj
SD7v34zxslxsQsPtsdoVylUVQjgJng891Onc5bb28zEjn0P7Mbid1xa7gGsTWIMe
MthBVFeYdbuj1lmBFkJtlKVoFCtBjQqR2G+j9X1dOrRlSPcXIS9v4wFMqVcbMVgM
9g1a6U/OT/hrgngrocaEDOG1FXfwHAkowbz5+rVReETzqSJblDasUsffp7B/VYRN
JONRp3nSvbd6Sl9EOAkwg7CzJpy5cP0uAlHCmzj3ApBFrg63u3H52RBu6VNJcPHQ
epiMearfdH/if0Uwm10qOZxp9oqbOWWeEoYr6R6h4bjXpe05Pv0g9luleDp5vgI4
UgVDDDQuzRwXmiQcxGFjLAf1q69MZ7z1R7JKYpuYAOrR6vEepkOpBp9Oem51HjSn
Gf0Gbx2pIQpiNy7B93el00rWuFHgiHKug2UzIpgsOgxjKCzKrDoH46siGW8h/MJU
DGi4pNBguPbn9qRDnBigcnI8mjGOoraG4WhQYHhcFD7YLBr9Sb38GPc9RFV8JMms
R2B6QDBLOzt+5gwb6tVVVGshAIo8uUS/F/ljgOw71LqnbWl9kPuA1853BQCdo/2G
/1Hd/EGmMUV1LbHGJrxI5U5zKIhZs38i7TXD3+EEwLV5YgppaWGonWc1qhnTWTlp
TF/SN411IrgjgcvVmtCCmqA9erEtq91S2WKZnuytVZBVfsr5hGmPEcAJnSGdONOQ
iz7i4lV4dkYuMK/AvDVlZIfpzuzJxE1ybA/SNX//nrQcnAyiVDG9Ph9sxYfxpxMX
Cgn8RbTEnnfsbsaaq0KXUGa5H1MqmlQMbwx56tvbYtmhYBpvOZ/yjV47SF26B6RB
nywXTlO/6HaD0zXKP0CQ/bwTUxInSlngyb+IihtSSXBY/4luNB6ji3mzTy2tbbd0
XjxANRy72LIxsgLzC5Xr6/fB7JjZ7/ApFgLvOkLP8MjkK+VK3as7tzCpBcqv8qc1
gd0olzjXY4gO9DltxGeK2Ad1Csbj3UozESedDxeNEnjs4Lt9drs5qKpKiUv3Xli4
763/QuURsyhr+28ui19zyaY0mtCB1VtqkMYOT2WVUaAdJg09xbOlnvOfvoLf3xNR
g5e3OgbCQ8OZlQOHBytQA8OqUnKLYxw7snc1H2XztSqRb01V0in683HrnHRT1HL6
B7ymvJ5Q6lD4pWDkssMJZaG+XKT95bGKlC9TVptnkjeGmQB7XqiMb//9mKbCCZtG
I7mCVOu8JdRTKdKW+0ckOhTcqWtBQPjora4xMioJKsrdgCxYk7+ln4bl9KPl7WtK
NuH09tDIziLTQIQ1QKjJJ2k+Hq+7XNymmP0f5R9SEcJsU4CYlS7k6Gw/lKjQN2Tc
QSb4sXc9R5Dc53BR4Vlal0294p80NYJHTDAITGEMZyl6JYdY6k++j4nl3QfdZ5+p
p/DDkKxiuxmyq4GKQMn5LUOmxRLcRswdtm6fkeI+s3ajzLUVreeCRcxDs0uGbdT5
dRl2FXkcmDZdXq6ml+qhiCULYdmPJNc0RZFhcgzqBuHEG6GbEs6MMC1szpABBFk+
tyi3b2TMGO6PlKvbTvXnwfRxgJCafzigFmjrSiYdFJWUQuHlp4LhRfxUM5dDJGge
/K/WEfpZ/cnWM7yxhMJteijUYP0t0TVSl9JpUIPz5eLrHKuhhI/it2PaJzCrsTde
SeteC1GDc2Y8QXEIMQ6D75ZKppPUOzwtZCtd2Id0yeOwYno+Scjl9HMPUTIOi+NR
D0cv0JxelJ8nlN4Fwp8vlxIRoU3Y9twu8HNv+7nlTIr/hY1bY7okw2DcHXsAV+qM
/wkVKF9F6AuLFd4sE9VVmWH7Z4Qjd2dvi2LZmci0cTSGrIj9yocnCyyTAwbQOTMN
977bmjaJ/tivuiTEfaI27ZzqSXzThKbeVXf0ibf7u/WZs3C/94dQ2XbIy+dZPgYz
5No13G+1WjNlSyJIpzA/7L5xFDI9huDD24SpYon3AI3LaRY6tuoycpn3Gm1NgnEF
uUVTDOoC6Yees3mN+j8qL2ZBeWIrJGyrWCs7btXXfSnFZ1dthA16ufjNXAUWcoyO
75S5StQODD5CDJibZoEmQW20dOBZGiXVfJ7CUMCE7DVa3fCbTrZTVGJzWwt3uVH7
VINnTWcSgz5i98dvJGq2wflK0jBBLeGc3rvMLYUwQBN+i/eLS0+FpGxPq4sSPur5
9TI3eBr/yjScq7E9zucgN7crcI+DKiLLMXSl4mmXXL/7NEV+/8HcGdW7RtdLkKA+
Tc961L8ECUTPRaMU6YDbuPcQI+ITOAVcWpLqyPbL0/EBj/mMaFZ3ZmzgQbUZkVzZ
yPNOykx1MvUoEdlttIwBvBqrR+gzryoTWRNrmH3iy8fwg1gb0RADydVarovZqhqL
sdEHhGAmLqdjq9BYRjo8yJrjLiz/IC/b6Xk3H17FBQezoxhUX7XS2+LsfQf9j7zb
FJFryNGRYkxc0fopmzJ6C6Fgf1jmHFsP57akIzON81bfldYEIIF65rLImo2waus3
Kv0Ue4sNm2Qpzdyc6NY+SXRSUKhlBqOidLueTIQs3+WZeGUFwhfJtgI4c89OkY6A
pXBMKPIu0erynp6vBszL92KMZ3QQ2SuFdYWlwvGbuqEkCjajXeSGiFkB/ktavXgg
68L5RsYrwmDJwKsGzzJvJTBjkww5m+lPdCaQnZdLTPG7druCq3H+nUVITVxwK8M1
mtvqaNoWlJjsFJwvX90OtK1YYMmZmbMG7ts14v55cLqfLZ5eK1bi2qVx+p+CPSsb
0mhu1hSbL9KIbLzSmNtSPyx+kp5OoJc9INggHqnojgZ0jvYy6EM5yu4ertNtuFuE
1sx3NH0kR5AWp9pSH9VfquzaYyis3K+w5rdxcZagpjjtWL16YM428dfzmdXuruzh
10ONcFq51PVaRWFllefDjarvQWf9nbANorq2S7MjCNDouru+enJXkH5eKIhK1bLV
1OJdbqrlruF8dGhJPc65jBkb0wvWdKuIZwifXMOqIhyeBxhDQQGxXljcIJtPEjab
BGPqa9zrJ5fDcSscaMTDvy4VIIz/vc2FpW98L3mVvCAYtRbNrK3AFgitv4yzgI+y
R08X5CQ+eoUDgnj571+sUe8iEiDw416IGXBpz4OkYlqrrMtT2lDS4vIJyXMfCFeo
udnA2sT8kk9AS4LKjSUo6mDf4/Dd/xkgnbipdoMIb0AdREo04skdVNbJlUWYSYrv
KDiXMM2lFPSRnR5iQyZwRib5w2DT771k3rkWDcs5cq5SLYqIvYsniuVP9xdGX/KP
gBNt6uWGHcVOdOWrzoGUlZuQDSMGmr8xgvoraz/dXQwvp2QayqvHbJrjcjVxEsNi
vTZwJmlX9qd0ZrVAdcquXI3w7Vtf1HYh0k9VPtba93k6EUJ6bqO1pT7vQ/fwqUT8
q4jG6rWTbaushGJfLlE8HGT2z1sc4c23YQuBrj8Csu6/ii3O7lTf6tO1PGJPJQwX
p419/Rr28sPEgbHf7xpvNwnGV3Vg+WgKJOTioklgJcYr23CxCq17W0vQxjsKPyDB
wOlEL5ah/ETmTTXoZUAjuDembwY0NQPh0JJp6IOSa+Gw3PqGP5w8jkBz7PKZpmk0
O3OS6GlMTmEERFO82VDmHix/RwZRa6e76W5K0rPXfMSGyLnAUHgSzyBfLaAWm/0f
jhEVi4psn3fxnEx8zCA2Wjjp4FNEwJMDNUbbJOXV8L333L9frz8UeevnlhbCU9Kz
F+oaWRTYHx/KLyQv3k4e8gyOsATDlaOZRrSIb1qF1YSmevLuX0go7PtHMjDgCKR9
6xziH9yrlgk+DUgRgV3RbXInGp2EdNfmvAgywqLdBWms8dOtlPJ0xaTOWV4Cd3AG
AqS6RWsP3ULkDxUHn1jbxsBH46H3tcKr9j0dr6uiTQLW7KYt+BMm2EnCMaVtd7m1
4jk9oWX62qmHRPlcXERfAgJm0o4dLwzAPMwEi9uLigpf69JoAeCUcdkpXHR+Kg3U
GSllzHI3yvkzXO+pUauo+lzQxU+m0lDIdwC8mgKpgVsBgjhsyFZAMEOaAjfYY8V5
n9iJolExovONeA/q91Smv2ZCsNDq6Q/FT/dQ1h/tmS1TzpNLw+b4vSk227Pj4UHG
BenmgorlcXQCvraAsO3DfwPJ3TdCty4M5u/gFZPvcpICMqdPNsJwhz6LKDOUv2nA
VdcFrcWNLKIXnIoxgOXI548GqRpCISSjtZhQOpaDX/GBvTOIbOlwpa2pJQbpbAp0
7piIyvdKcboIMvsYD9ZyhcqWCvRN2Y277g2a32fK1BInMbwFcMSDB9Afe2SAZ1Tz
9csTSSG4p42H5N2nbwmm85CYB9K1SgBIdDBZa3eSc3M0CORTaTCeuiyt71bonjXB
23fpnsSpQuNge8ux6oWH1QnVblKM82cp9kTLPSeqW16NGPq1GOZ7jTbNa0AL9OrR
wLwMD3+aoXBtsQtzT74ZfFDRzIxhKgG23BRVg7rZA6WTmEFV9kvJAWWyh42Sm6M3
8V07ADXkfPkEMuTDwb8q5VXoAmB9YUeAFuwv5Zo27PfmA5avcquj7QN0L4DzX8/M
KvMG8iPYEKtnjBGEPSYCGfcduptYrrDs8881Cm3jXM7RBTKPp9JVddqh5gSFYq7R
0kFp++4Fp7H+/ga1MTMfP4bzEXs1lUqUpVvMuG5sCeWj3WBBZyraQRxHO8fBU1Y8
6rUeSFQkjGfzwxoHgGBg0CCEiS5VRb+cwJwIglOGiIdsD+HhzCe6H6NfNhIdz1Wg
a03wYUBXKncms9HXFMyF5ZFQcFWREbCL8l8DbQHkT8ZPdS3yUak+JkAKgrcD8/n3
ECCoKXetRVU9A8Bq4IabgTKgNeOnWigETZDdnSi6g85UaMyh0CuEOHa2LI8LAmTs
ocZvn4JWePuJBtFQM7WJnXA9HmozTQStQK64t90bZGvwihwq5mpvlFBbVW9x83sj
1TWpYjrn65tJss8Yg0zm+z0NC1GEhwxNQgfU0sF7VnE+3/trZjuMXdOvVAXmtvDX
1vzYtBSfzfPJFH/uYv2a8ZZ2Y5WXs709cXv9435wqmyjIyeFpUtZtEshuCSKMaFc
0+pKkVS3okzr/qkaBDbq6w97gn35X3ZMgG2giO5P+ZBMTtqAnQqmUpZOh1Qcopg+
dT7hutt2qfmaHOYAbAXrlz7i0wvcl3S2GczWwz8ni0z/4hBtXVv39mmNwe75ssx5
T/7NFXc7Cr5krmPkMzgCQKB59DeBIWIvW3K2/PYGtlD1G4UKW+OgAYhYgMqfttdG
21sQgeV464Y/4FtrvXrnRbIBZSDk1J/iy6vIMopK9YYavRYpRyZN+3xSkbxNDv8V
OqYJlkTzc9b5PQN3QlFQ5a8lRxUp5+K0D72BsSek4cNRuNEDRVfOfimhhnvR6dsH
LKpYydKTd3d1ccIDmF+tGf35rjF/2GXtvO3UZT24Kn1EMt6zKBzgjnH08g/fbTTI
9TkHIX2vpMlwJCGT+fOftEDBqzaPAjHPfLdTTaQjrApbrpqQS+3k00uOZ1z/VKNH
sjIBJriDb0TBXuK6OASRThRVbIb7bYRRL1FIE9G+yzOU/DuPgv08zI0NUnrgt8bL
N1MpXCyvWJBqKG69nuStGLRG8WrO7gPrpV0qvBloeHq0ZFzW/IDKKihW12A+Sa+k
9RipC/LoR6e0Zw1Aa5FF+kHuyLSHNj3wf/rRNkhvqZ0m8g8DqDIF+hE+T2eNMj0W
BzSB0Qsqa6PSNbsqDOhRJL/LlidiWnZtREFGkPQOSUgsPE+qVxBwc4zLKpJD/egs
CXYoFgWGW+RMouPzJZcJyhb0+EgoXE/7s4kJli8L26wlcAYU9mqhr/O1qe2LpDJ4
GNMpwb+yG9INWCZNL7pJHdoOXY3MCdILDHpKbn9KeHbSeyS+AzLaibLRe2/syAon
2aBDUC/pe/qltV/62Ca1etkGm5G63FItZ72v5dMt9l3rz/mKX6MPXvK6Kb0k20ZC
hRBtC2vP3yYFpW6w94xIxYu3zwU7i+HCDFnz38RJcKN60jJJFOXcCSmbofXX11Gg
jcqXAjNenQf7Eimz7Y4vU5KyKkNv7Jrfvq4g81aPHjxeI6vRfqzHA3yNJp2oYhao
U4dDQNeA3jSJF2BBbZUYBxqldXGXs7CBoKQCSCtnXfcslfdOkd6D6N9ztioPpGjX
LVyespgkm6WIw/fx29wrRP/A2ZHZz3sTleRYU/e1+fGUjb85x4xwPqrmtbk0mOHe
abvkjLpkF2H26nTuingoT7X5L7vk7t+30RUgc6q+znNWYcJ9n+aeInLptwQf7YT7
v0Iym9QwJe1M2bLungTk3Ih+KRWgU59OAIpQIAr/4AFPWVxwCn8Xgx0gbXN9zDID
c8uDEUFsLYGPpyark7Siu4sYOPGmXJTDzwLXQ7EptEjET6TsfeVsVhheDuXLIECY
D9ne1teF8fyqnl9iL1JODrIi7Rw4cJfD6JcqFDU+3zQcbARO5WmcFj+QERlA3WnH
jjkrFO/49xNBMDqwBx0zjWOnnSRUJ92VjUNXAvpI2wrfr38o9eUgMdVJBCz7D0uN
ihXn83PjMUY8m3XNFglqMzeqQB4RayuGKDbioe44W+t8si8IC3VBx6RMS5c7ELmB
5sGsLDx/A7ijzitF2+++d6EXyigbyNsFWih/TDoqtN4uBfMr93rrrW+we1vd3lQJ
9THpcHsNMkyKFRPaOW/xbVcrQmwxEckF1mEoDl0LQ1ln/SYQBx9csVgwMMDXMyjI
V4lESOIgd7PKzIhC2LnpeJDuz0NhgbxyuE/lx3DW3+ArVsD5LHIMNHIX9exNnf5h
R3uXlXlmzogQPOvgMWMG0kQsn5ekwCqhI5F0vv/ZVoxCv2TnD1fVv4ikE+TC4/QT
rI0/54QsQGPZOc7I/D2UFd4ylAa46FYml1yWNfwG7ptvlwjchVu8Yi6Xm2VnER5n
BCNCw056672PDWIdQTea8Aa0zA9j4PQOZtPmcPTY3WWPvNAQ0qmpk7Kp4/bacZFg
DM/EwHSpCWDC7DwncPcp5sFxZtPXHpBdaFIrTK8Q9tlLLmRLTED2ADBoYasbUdRD
use1ZIdtFnNt9UEArCZVe2irV+6uLyuWen3XCuYCARQOYUvE3q7MKcKhxcehQLWt
UCACrLj6/iyctLd/+qfVIhxXFAQhbDTeilHlk5e5XAlMdFWyiatUAuqg089UjooI
IOXIpQIKDX8LZx870J9J3E526CoapBg6J9W9d3xgVtA1TCk0nZjEeBY+javvFJ6p
ZjjWQi+eShbejaJ3pzkpPN+KMYo98f856cLMJiOrhtCuBhKDbwle0O11hAZ1iSzz
iPiH4RuhpD+H8RC8yyigY1ATRhuoHsmpb7vPJ44SYsq/sdx8TrQzrJ8YBmuMP328
pCYAQMdn+bO7UoDyGahL34SufU+hE47/rDMkMlDJoE/hPDe+KOriSVrd4YX56cy8
7+BpDVMsCGYlx+1HSSpwg1dolmiRRQt4yd1yHzEzSdr3ZKHGv5/u3mHJOBQMfMrj
RQe5s2pv5pXgxBr6XJzV4yNSXLWTcKnyzSRWBPR380bcAzFsR4w5SMijvEc4aXqU
eZkvT9Gy/hg3YF+BWJIf2rp9kCvfLmI4vF9eJl1ZYq0bao/M6a6PUV7pnfzG5Ncs
Q7QG4nMUBEKqpkIfdvyvA5rUxXYkQFFM+VUkOtf5oapvFQlpk11+p8WuW9q7OUl9
Tc9lnCLsn3dPen3KsHkCMKrGbBLGnCiw9miQf+w23RDy1mZDMHi1BCHLREdnzi4f
ZrCebMqpkdySAaSZUQ6Ld9lduqXxxCldiMAlbz5F2tmW+K92ZU173AuTTEZ4Pnw3
majGTJ0z8sNxPbw22LJAAe+M81TDQSG5HeFHRBBOj5g/g8/AM4Sv8l2vtQbqS0fo
B16i2/UVlvGae2B47P2QudorGHRacCeLCd4AKhdlZ203MfW+Ti7CwTf8OzuNRkGc
VH8/sU3YPHvompiZDjFgrkO7mfimbcUpv1//HAwBmSCpL30IGSHPxMqbcC1RK4Ng
lu2w2Rx83JiLtTJ8+r6NVA+9lvsTIgZ0/G8QjAJofeNv9lPqkh7Ad6pZUrahijcs
Zv9iOhBoltJYeJN1h8n3PdrYA1j0L60cT0ZYkh8KJl3vVg0i2Fg9pbF0HQZibri5
+tljaCat8Bz6MY37u+9GMkkQiUnuETNzOUHv8J181GvnRNasFHC01ZkYlsLiwmg7
5hS8pVtKAMv0A9x2cnp2HxHgv3D0lAYWaC6enixXfNRVCOyXTXQaRFh7wlAeckBi
Cx+elnpUrfkvDMpYAYqrIEX5eEo8Y8H7u8oi41UaIcUbIpLdxsNa064tCt1uFBR7
BN32i10Q1o4naqiNK45KUrnH3k/pMQMwkanbgXxOUGoc+v6DSSNmoLEiDixN9p9F
3Iz/BLC3r7HPp9zSiBKbDR9/F7xjrQFJ4tJknK7SNkU/zltOTWZ/+CSVl79KY87g
Ao1FftrWi41znkPM5flQkg0MF2cK62UCdDXhkP/vDL3W9woe5+cPWIQ/s5cqbYWT
vTjXTko2Gz9WPMcfz6TdvrztQYoiJggSAb2JSo8MR9fRLbqUSUoyeOVN7BZSsglR
2jXMYInC0BJ3MQ6r8cpBxle1n0TG4DK3DWLfuhWple48h2MaH9aNTXOLtM30ndLU
u0F6whCAcgNa8HIz0EDFVUoqfjOFTm17SUTQ2a1PM20SuHCrzWQszWFEtde+kmoC
H8EjNxegGpI7oTtE4PMsw14D5b8iL+nmlhnHbJAAfJlo3Kf3NXCh6Eh/uDOrFAPP
9yHqL593zl0woOUr+V7p8KTPCOWwGnndnbf/ueNwOXFaD6Ab0qizJJd57AMEikbl
ng7BIDVFWoExepdY2HWFFx7F/VQ3CvLV3DNJqba79wyAOcvaPhs8en1UacP2EKVD
4lbzOFkd9tLiPgt4dlISGGlDJ+Y5xV+ijyZg3jXWFhWkF6HoJNnGBn3hLaLMdf7m
cJqO7alfXErltjkx95SQL51e/WgRv1lpYawFmD0RsoVQJ3eMK/5tHAxtUv/1uFzq
Vva50GQJGWpE/KWRmoxHLBWhlgT7IkTDDtF2sjATBs+DuleqdLKbE9jCN3HiZK2h
OeGoQojYByskEn2/xljbCEwQvLGIktlsOmhZuSFcZvLVB6bafEdAAGjtpv8FMoJ8
avKnDFSQoG4cnO1Zxh4knMVl6CpqidKP9iV+T5Djb+I4PWWvDVeVhmjp+ViPy8Kb
r3h+c6nJ8WZMCJjELnw+6alzalpXmcXeM76PthvXmsSdfZfxyBKsu0RzadurpfQV
TVEzn6hQ3Px6GhwRzFGmHSbImjNdMdodEitrXoxzejtkAWN8u9pznTxbCcSib2mG
YbUOkm/8EoLS0wxMdtDHI3YZMvxQEo3VU5eE31GiuORTuIqqBv3lp0IuA4mY2Bsq
B+sCxW82tSPgOi9WEw/Zg2A76AwfXNA9luLU2Sm8dxZAyKlNQ5UqdYkHz7fqBbwi
GyZoLj4PiNb/YI6d2MTwqIpNkgQsrWI9+Mr4OvwHUoOxOrkTebPYv6zijxosi+GL
/+7j0ItZyaUKfwdJw2wTAXyJd7pSGuBPMOaxOu8nF94iWq6uHO4lGQtlVOHX5F/M
Y2HTHDwMur/BblWz1nT3/3V5NvYkYfjbb4FM/dMZwP0l/3VCp5DoP1WOyNT9wWXm
xHpRrwSLtoxY7aM3SxL44TPKosGs1Qq9i1KhJIwctIYGhdkcMFFuh2MWAR35LDx4
ZwB71/KD1OZRAEqOha1rMKe6uKrzd34r9am5uGVZ9S9B0vOZaIKTzTKqJagoVRkJ
H/H3yvWKEoYSx1fTwL15Ut8uhdF2iOsuQ+/fTsLnjroKOPYnhNFp5MBZj3cjtHyS
dXbab0AH67hL+Q8aPDPw5B46vJItVakglRrrbnfs2kHwOb82RbNkw+n4E3sGUS79
pIfUB10HmOi5WF4m13QbawvQ/qtwoG6lCQOTdXXIl9ZKJ3E2TIohnxxsDuOrVcmy
pSTKoiN4fr8nXo8Ygfonz4ficNPOBVGAG+3btEedfcMOoACi5hyVbObqaPRaWenm
1cocCxKutpsIYFTAVFUv0su73IOJM4js3fRBeZv0RwRxve41mwYyM6l/TnsSIzfL
T7o4jwm7OerOJNZTeFMhzJz8AnfjDR6deEED9dtVi2YX9vBoqf6ZCBM3uxIGW+Ep
Gf1IRQ37oF2z4MvU3wmt78h/NwtDm0x9bv8+dFxzVhgNSO1yxHGtHXmbFNWk2Ic9
TWUsP3Y+1vb2E9xPhUkdgq410mqht41kflFbKRHbtNpDlA3cV1wbY+sKUbGIzlhR
jZQ9CRyorrFhekodaZq8yhCoeXiiLs7QCD7t5HLZfstcjPOfYgy2KXUAtfRPed6p
xy1O8Mk7MCkkQe/fGfvQGPEttY+59yGmnBTZkF/S/FNRv71evq1Dybj82zi6lgPm
8rBFEgSweAZ8m64a5Mr7aQNd2A9uM0EutkgGjj/rzaheTw8LzhIys9h9UQuAiGO6
nwzAfGY4bbgm2TdB3KopJyYZIozHbpbpUntWwdDk4HkbCkzZfSgb6tAChDRERraJ
6EbMl+sNHhyaFeKZHc/URjA85UUPxPZOA8CHfv55/qxT7BFuNlBHL2EIvaYUmU9Q
cY2MSnPvH6aG0NiWnQC/WvaObJxhGLpBCnKXRbhhBXTSgNlrJ1ACzpZwjIilIhCv
WxZbLU1x8g173jhHHydpWWOjintmm4XdtN6noh5gbZ9UtawEKZpBpZbzCnZOrDSI
Y6lrbwEWS6OsX8XHfu9KYS0ITEJCkR46Sdemg99u2fHTapqz8j2oCM4HQ3ytNVdP
hNARymvkTV3js4fk3lUHZeuwoUT1ITr/razBdhgFsVdD+KXtXRb4S36JewHVV3iO
5r17sEClAA8v3/LN202pX7tYmugSLf1sIdtXCdL77BIlGVHICsMmN/v8mzGF/4zH
ry+rArZgN3bu2aA+YbQTQnzhTZYBJihm7lsVruERtmKHwyaR5KUR0dya9PV1uBoX
EHMq0Gd0MSAFqPEDlvn793V/CjKrNrl4S9uxsyHupMcc7Ul8HjmhfnBwUC7XkqBx
Z36BD8gu7MQY8lXOiQgpp5eiZtLPJVRgrsy09m2ugx5GP878blWsL9VDaPKJsep1
+o6xoBMPAwLQDIgcQ9VvR9Gbqf3acGRHoYz7ZfKtrKH8eEY8xGPkV38shiytlxnX
gLOLSoP68BFFVS73+MYw7VG7ny5P9qfiRPBfWUGkGqA6/fKoEP+Q5ukLhcF+niAb
m7jXNTPiE9bydXxFAJ412/uwLLfYl580LGeWoXEeog+lsPudwMnDXRp9CNvRxglG
8mQ9N1tbmmYywvtFbAZEl/TDTPav8NDYXdp3AkwQ0Wpgj7Vr5813nx/YxWIxbNn2
Ezz01x/cDkB41a/jZUDJ4c/6C/ziXOt9VvvlB5pzSxCUAfPglR0SxpFoOULbLuuk
JQz9R+Jq6zcwBd2GlVNsBpM8WIUaS79RMh3QrPs3gtJYicQxkH6Pmr5mCsqm/YO9
P4zq2+Q8Lr8xekzyE8zMsafT5aHBKM/SacLLHGyHPWFjkNu3oZ6K14jefTBw1MO3
1eazmoBphl5o0DEJh0NL6nV8wakVVqnqTOLyjm6MtcFHTq2kWxXGq9a6QjIfkTP0
NFKKVc/DksFbupTJGt3Uf6ZEZvgdIV4O1bC2yLRqqNFQ+AH8KYecxY4HM2xCkTeF
fHAfwBBhoq0zRa5XfNqjuBJ0ur3zxYGa+/kQWyiPlT4nDWm8yJYfHhbx2M3MiTsS
yz6h/tGFCm1poKp0vq/+UT2A8QYOshH6n2C83JkFHLNHYGM8GcBp1SkisTJNuvgz
INJq6reIRdytF2fXpZ1sWlpVCb7bALzR2qn/10Ase357meshPF2KOZgyrSujAlxn
m52SCrwWKoj0N4yHXT8vUZ0IzYEbHe0XSh5K4gi8WbrH3BG7U/ZEo1koBQuYH0YW
kuK/MFBPJqLgM6COjNSFadOoCEL0hW9mA9CcOCy+Fl4kPGtlsWEOAfD7VmKu9vBj
bUvjiPrkhC5PuVjscDX7X6iFCh+vqFANIfHJPZIuR1UR/EtT5O3gmuFaAyquRZFQ
jAzN9yAkoKimEWPOE0sz6J4AWbn5VnRUPyT5jFPsRdm76str1TxhMwsJ9XhPSlVa
Qj+Fu4QcztsqfQ1HndQPSHIBgZQSZGHaSapfsC6z1nvMA7z8+zZSRtNQulz3ErwY
6AdmkL0+p4UJUpOCbZFnsv/a3lR9Nh8u+K9svkGjH+4WxNPabcMrIZyla75fISO5
vWa1530CSm+48mcHsnJtUFSgtqiuKIF2dU3U70kke5DVzezIMjI/GeUtrZZeEAAe
rSEfkIadb/yTTIMie5zAI99HyqXSh9sFw+Jio21EGuYmlSHgktWusEdDlY7vAOXO
ypRXOv+o5l3qId5fuZ90n0YvkLZ9TmvdTkAGrzml+TEgryoQ1ekgrnDn34Nq2ioD
Icgz4z40xr4VXH/+eEh/RfR5ynnIV56NHlyY4+uECasKH+yGnd9bxMMRLhYiziuR
dQb/XH8+saiieD/nEhRdokUgKw8nxhd7X3Gji1jNNZK6cP3zcsHAf0R7FqmXiCzy
h9NZ8Td2b1jg4/66CPGijCqVvQcDdxO9XwDe3d6jNmGyhvwptKEAv5VEBu1vyrgI
NTXByvsWSLM3Xw+uLRuYV1p34ntnGRomG0krocP3i/dh9n/yqJSIH3jYGNcR1ihh
Qnkwv/J1qEjNPJLfUs0CV4jXGnO40ejGBOJtyt4ecnG19JbtpYMwy2PySddQJ6fU
Cq+Hz4ps/QdUbYLb1RkRW1A9WL8LQrY/in24Jot+TW7wc11uH8K0hHdwpW671Jvo
uCKZNT1KefU7OMzvVXxsvFr+pwhQ3aEZ6DyjduUTFTQdz12iA8Nf+LZaXjNuqs1Q
YFMQYja0A+CQCtvkRXJoWIson9R1EWgxHPrmLid6doGMvxztvlPCN691KPVeQ5FZ
WprcxfMOxaiDqjfEjXcwY56b8rseNoH1uZ2im+kWq7dT/GfyPs3hjTvo9eoVfBX0
LkkhoCSBoc/x5kMzdX05aocX7jeDhOTDH0px5i7SHt5RHZ2P6MG89fNKxbp4shlu
YnqpeAOAnMNatMiX7Mg3MB8mE0/IanZTHxoMWK86DO8zv6CI7ekha9jCHwo/i17r
vDexKDKpCkp2r62WLm9g1hGHNIJxXpWp8hQviNm8uL9Y/MyoLCnDHH9EOlQ6IoUt
OAhSWrwLbwdQl+/NYhOr3gkXxY6ntc2jy9uTwl3Ei9IjPnhbdfPnfFrW21yXAOA/
lDl72TKOrRekV3ep/LHFri///wp+0Ol5tBZkx0ssF20jEnXuCrkmCi8Ytng23QSD
+uG9ivg9vV61gDsalFLuOtmwceNcrWbJxdP7cB4uQkWqAPxYaPbhjFQInGm6tNZd
uuGi7cwP3pB4/75Bhe1W7jpJLZ0/KWKsUsvd7o1I6NVE8zrptLcM8cByEJE6Hf+B
rT8hv3WrGkQgINHEjqQrmKI58btykujVV8WfYF/hxws4Rt6VF0f3pxz3Qxgvri4j
04/pKZQyhfsbZ8KblHki3o2nADYqrzP4sex02I2CSndFKVpsTI/jWT6IT7L3Evb6
bKZ2MlPN3Wpj6inT8AqB8S2HDHaW/lzhjdfBArq6lyzVLqlOc8AesM6cU2pHkS1o
Asn2PP2gPnsZLG6GIe/g50IR78mPD65pqV5ky0lfLhjxueAAzSorLRPsFeHxC09Q
qaZ2EK5Zwz12glqI7zE+Oi7trL521UAWI91GbTxml5sMqBlVrFVS/4PcS5R4GywB
S9dtFmy+E4uAa2mkDketKmgCVXmXVw2uKdexJSeKEwz3rrOBH8hcP/GEnNuGsT6L
T2zPw8zLPPgz/qv26ZSVgzBCw4qgGT8PCOIwe4HfeH5s4YCmf9Vb2RnYbclxYLmA
g8hijPiB72MyfdMTgeFmNREdn0m4U1Yn1yzp3VlpjZigM0Yd03YxqojIvoNwXgdA
GJd9Z0XICEkG9qTUz0gMQQ4ie5vNDQ5NHSvA5+78j7VS84yWDeyd0iSq801OoEUx
G6FAbyydoHXSJ5S1OH7zb8C66uDN7p3HOFrikWD0BuP9RGopvW9MQWzdn755lBRg
nOVMfCSUbkqHoiyuj/kb8u0N6+Aywkgb6AzBg0FQsTE6z51mOGt/1Oj6EOI3wpAD
O7CTSWIZ9ohsekyBJSAO90LFQrZuU4SelH1kPzARnb5MojGxIrxtVcmU0Yxv5ebG
OMbP2F04278bo2/tT6fq3LgW4tgnStdYw9PVrJ9pGOY6GUGfS04+8wKQ7LIEREeu
9o3fvJbzsdBS1zy2RiHIEKE6/02Z5Gy0uJwBZVne0VC19rInXdcyS5FHykJ6139R
H2Y4c1YTk5P2ICzwMuUnL2+H651P2Gb6vMj+1tRjUUxysGd73XYCBuASfLxKG31t
Y31wCzT21PTdICq8dMaurcftKA+Ib9Nmj5qoti4tm3+xGkapsK5N7vIfoAbVEwlR
vTAsBSAwXKAInKSL5onIoFxYAWaO0cEUz6xkBilZaPEnTL/0U7arQ8qzOiQOgYLC
VJvYBv7KeTe+UPWXbNXfuArJVUnZ2fUpXWR2wwS49YDsuSqnp6DpeXzHHtDRwcSN
VDf26lJWe+JoX2ps+l7hz7W6bZ0DODpF8TTk8izPdKSNBLYWTS5KORy60ASSIz+M
oI6WJq6wfmIDTlrnd8mal6dbWlvDNgVcXji6UCfbrfo1B9VindEs4G7W0V13gkef
V53XmP10eNpTPeXbKuifNMpVOs9v36MggkHcQBvhOpBsW0qtgrhrwK2/Yk8KGAsP
oS2+b9YLwR8UTsGEtFKpMpDk35OpfXKeBiqt2kFJTqgwvwZdF/DVhHH9rU9qqCVp
g+9K/wr0KF20GVqAyhR14B7I4UgHxPZO37a+jO7s9gPkb0T6fMAHlTO0kzKH7shX
ARVQVvh/2JsoF7aQJ/89R6vBc7IA6llRNcgDSQ1OMNhRhzXdIOiE+fnQGhb6J+IX
OTSttFdqR2ZHzrRHmKNP6kptVkxfVEXgO3JLpLTGYQysYS7GZvGbDIKLefr0muLC
6GErH3vW3HaYCHzyo8kfSPX1D1GImRffR05VprnzuT11G8PVfHJstXUNmpwP3jva
oeAkPPqPEbz+R+KBPZ3IxyasD7Z/5c9WIvsiIsFcJa0e8nwat9Tgt1e/Ehoc9wn+
DaW2zkZr3+re22e+m1a93/B3mcL12f7owY2j2lnO9UBdZk3wXRHJupdqS7hhMiFO
2DiSmsYENxrHddjiBHg9jswV8833E3FjSexzQBCWEfUkYr/4csvtZa/ZLjMYYu69
2ASt0n47vMxj8wbisbYJjZqFC2E4bZ8ldEN+iG5A+z7XhILLvejCpmhcz1l9j5Dn
pYdr3q77kVN38qxGzzpiMxuA0LKekaSDCEHMVaPLeMpa8ZNR+onoRWZWSDptpXeq
tZukVWZQmHMjsuK8KJEHGECw9hAcNTuOPPu+fuVrjtqKDqdY2U6xBewmYOfpRdSa
N2P3jEUtk2r3MOmZOk8d3Uw3lbiV5DIsVIAFB5+eWuNxGFUJ1yuF+fNOaHQJO0cD
hdQGJLVvJmBIneQ3LSu6UgAWh6ICN9Yq7H5LjsJEk/Ld+r/trhcbvEoJj1MUGt00
kZ/xsCxNZFk6DA5nINkr6ysxeSkdniCtuScVQksIzx/IE02sFJ6H8+CoyvwHp7uc
pwN+Zgn76v3Y1PxNYR7ubuLMTMZw3pZL+4/+H0kx+m9PWpEda7X8Wlg15Isr7cr/
GmHmW4aDmd332qFU+cvzfEzY6sgc9jaf57BvUCXqI/KlXrBXM5eB96vf4JRp8aEU
f4pqN4cYNizaYYWh1DxE6cjCsCo9hWY+GV4Drk003Y63Km5D+w1ZyjhgnJKkaROs
gJzNOdP8Yvlu22iPf+eLs7FLOkPKOvRY7OjYxdNq8VhGQ1VUUEDp8WIydnP+y48/
wbfHyKsvZ4vw7mTHDT6+LeXmNX4qhZDdZKTnwfhNUYSNuP8J/8rtqkcPnKCTkbSj
a+GsDWVrEtUWQlc4HncpaoxPbY7cVntaATCnOVz7+eoDQ6VW/pJKimypHnbJI+zY
IJCBNA6WS9ddQuJkPiB7Zuhnnd/MObBBpG/MglenWCItNaNe8CO73AjLZNQ7zjix
Ev1QUfIvgPkNhEU602lYOq/UUpo/p78X0zp+UbZx+7f0lk8SJBBfVekPUBxZJ5h9
M6L+pJMWHjaYZrLRxOkTeOXFva4F6BzMyjZHyLfNPuVMguiN+J4DnZL84rnk8ozA
GQAXcaB0WoA2OHtklnPNVKEzRp89c6J0jPuAXyBkpMnfl+HzYyv+RWpipZxZPh9I
jXwHlPGZJENt8PUFvWOcKaU4xDEvongzrXOHbXNcNS9AJa705nm3Sr48c0lygvmK
O5ar+ZBVfRpirC49LVoCViNTpwIAZtnU9vi9hcMBXAaXECp30YvEWYK5rsKBLDPD
zleuDvT+Q/3Nez3JsvdUfCCDWgJ2T3Lnf0uvCS8DY0blFpiz5H6+Sbi84QPgDNqq
QKBZdOLVuKSgtoK21dew/TG8hanvXKhFsAzmfY7F1QC6uBDEMLr1RSct1anPzV1w
SdbrBVWBbC1INq9cHpa4P9lXqVFvkHjKvZVA2zm5YUBixvchiy/9sFs2HAGwpJTE
/UchVvOK3pgWk/sWJj8z/5ulSfvUAtGpQChRaOS5Z6B4cY1TAC5nj7w1lKIlrHuy
FufUMBHKrJIdKc1LqIsdRG7RMpmEBNHg+9Wh3CzOv/8Vgaw/50b2QEIhuZPCrkOd
lPBMfnk3Dinh7L87BplG2wdKzg2GHXUIFp9alqR/qyj3cbKbyZzTnu0iFD5bEqFd
yqu61HSt19NYACjr6pnzZ8S7wL04ABfNI64V8anhxIap9RLJlqbJVUo4kwla+WJb
cMH7Y/SB/oVtXYJter2p1habYQTuGeRf/2in4ReiYJ3xF3lmZJhYevjIuD/ACZOm
MkqaE+ZbUrOu/5rS8ij5Sttfx/QeZwZofxL1Mh69kHReI4Mbr0ie5YKTX4uWp7vu
5LMCCcN4N1LNAtxYdpoSX2DSSpC/On+SX6M/BCFAWoDlpzI5XFnTlB+tQkSSzruF
9PJxMx7EzwWY8IuKocIkthYdtJAzOBXT7m8dEn39PYA+0Vv9NJngG8IseeVaEzCB
JpZXOIMASIAkXEWCT+6hRO+4jpkBYk49rMU7F+4SRjubj3kPcVMZh2TsXMLm9sHw
tc7rLQVg7DdDEFptN1yQNznvTShkJ8mpDhofZm0a2zdoi6sd+6NN71lrm5gIkEcj
9NDYjqpLFGPGf2ZbeWKzkhbux0MK5smhGR4EV6UL3TWVVzy5Vf7UMos5U++h9Fzc
WllZUXbGN9j0rLxUrSNeSEFYI0DggmQII0jvIYSuGvIZwkO8IVS2zUaMzt/9690j
+SXttAxXtqg1pVI3uhfTvl98nZySgMLZjzaknTAV+y7cfSLiA3tJ/Okc4ypRMwhF
tpSp4pDfrm1EinQpTnUnfm6mZSefqOg6zuxEsuRq8dKmX+1QxiO0bUGL6YxrDZ9E
ZJr6hUdwpPomaRsEyrev+bEf6+rz3BXcJ4qA3XHVnjgX6X7FC8df3Cf/b0KyQO+1
MZDGZiXFXR85qZuYtaO4ElUWDaJAypE0bxs7fSHlj+zgeTG2byT9xAe4yRiOwZ+Q
gx5ydodEAZIO06o7JDrld22j7hAfbbwNRR7oI3UqfsTaMIfQaO271gNHCTZcccVR
qbHVRrUTSuhwEomhC0m2L9BjG29L3IeIZB93ufHrmjqTAxNCL2cMeqoiGFQ08WQX
SqN82SMuuq8o4gcxDWZSEqyHaWFeIbNwYnVbBaB8+xHU4hNxPQvwjYsrLm3eRRot
8qEBiRKY+rmBXLNOi2UE56QKt7GCiq0LimAjkeIPqmfMlYj/hW4GRu2gFGvJVY5u
bGQMui89HuLznmPteQwbKR8G4Tg1Vo8hUCeFMnTntvjIbEYkp+422Vi+bDgMqq1Y
IX0rWp7T2aWWbfn8pwKG+OvNrHwJfr/dutMLpGK5l4x0iDKI7VJPBB///fBrpjHx
VaFyCxF/teiOdJKFlyI1IKPh36oFeR1fDiR7h5LJtXleXUxDFc8KG+wwvqXoZzee
XEIaVCPD7d6vXg2tpmKWEzO7dng2DzTfArJWuwzAV2mF8c1g8bqF7iN2p5giB+cw
zOCWejr+BY8ftvD8kep17CCGlPwdBpknk1qHMFOjKLFW8Hjh3ZAO79Wt2m/cWxzc
lCFQaHos4Au2hHJBYtdAy0i/yBEAWDcdu51peV84sLvawudctVm1bbiy01DoIy5d
vcQy0OKRoAhFevRzV7DjVsuBJof43SVwguhUSPJBCcewCDBcvhodsBGf55I3b4M0
32b6ibvHHbWukah1fE/SgK1cF3sTd09MEYNj318u97uXiIbzpzC0tOYebSeDRXD8
82TDnRrRlgw3JvYNiGEB+Col0ZD0KwPriFGO2zaICSqxpsg/ASeNHdvVYr21M7UG
qcJABqEO0fttevZjEWfuw8+7cUb5drlCSH/FgIIEE56UtUSP6IT98QwyBqd/MLRd
bHVeRGI/Rd8xCAFZxSzpW0wNBD0aRM1uWCffhsL7OMFhU/VsLLaxVEd1/oYuMTKT
LQlypSm2j7wPOIieJAsOoMljIgbO+11xoeK5GBacoXxZ49icvRXPT0OnDEr9ftJf
nSh5pULN9K54msBebGlW752aLNxxEFL9J6paNHUqvdx0MT/k+1Phib5TpmsF+ezp
bYe5jvu961p5+fpUhnDeNz6BkpDFZzSwsMutsPVCU5BR0Dw8d5x4q8M4xvbMeO1j
ZjemUQ5+g4APxdhekGhV0BF8fM9nqf0HLWkaSb/x8kAOvKgCbPtzuFNLHNNAc0HY
Mh5J9e17+VA4znvGmMwbkZ0TEA1J6TZIhYgY9GlNi3vq4QhSYKDixPWEYUalb/tP
dqFavntgvkOicw6mNk4toP0hC4N2rfA0DGb7J+ybckkTYkly95g5GET3s+zVaAnr
cxldRY/fagRaT3eTdTtHSs+6gn/IajxhoftsIkVecaiwQIXCJJPcO7NoCLg2b4Lf
0xxoWrSOUiXnyBWN7cgb79LG+YM7JmATVDykKs1ETesXXO0yT2NFlSxN01+EMsWZ
FG8qUT7NBDE6GGLL/z0TFynzvM5gJGhkRAIU7o7mDKY4VXUtfhFsX0QbWPMP/bvb
KjofxgxreTtKijjkXNFuK6WLaUQmhIEjq9AFpohV8+WHT2k4KzcMIaF9q9ZLfzLW
CicaFSkE/7cFszLmGQ0VbCjOwY4dhyQMcAWU/UtIEdhfQf/P0dpdboS/x+nEQX1Q
+RSrh7fglD8mAlVmDqbyt0khsFD97u3OVTKYirIsaa0iZ3dCU04mwFjFGbnA0UbB
pXWy0yDh66T6SVhBdLiQIDoJusrkQYLMcc+SzGsnD+rNb7OC1TjvzYJA/KjkQ86Y
0kC2wg/sDOg0QE41XllsrJleFl0W119387A8gglnMCEfBlCWjgGCLIw8j09MG3gk
7JJXC3FGsDYXVdf5anSwu4LI8mm8ydVmDk7BmDvZAFmXwnfMC9XSwGjIZMkZi1NT
53pw+1Q28e42QMNQtTnPySY4LqVcBk7tvmS4InmfNnTnTpSOdNLbttHoO5FRVobA
oOubrwyQHMOAorUr5+Uhl80NCBPQMnhCwI605I8pWv+gV33X1Q5ls69M3mKeONup
yzxojVDN9EjG3DWm4YnV4TqnQel3R0MVk0Kf17w2evdPPyQzdZInHvc6RwQbdIMP
3pvX4S1z1IeblGrAjMdPUgek1ZBdVGrCcnTKLdBtcbrB6dgMAlYzgP2V8L5Hlj2u
Vly+vJjdDN/16Uv/gFywYYy96XfvKWdRavsuMkr52nNLLRb6iQaJu8u2Ixulmn8M
mfo2OGLhoCJeL6nAhBz4+MNagOx4MOfLkub0MzwJgtUaUBEbF5e3lx57FoVnXyyZ
KvwkPmdAvoWmsGnPYc3mSoxfNVS9Ce8Ja0WV4GCwEgA0Z9hQ/vIaf1boITp7QwxC
vv74lk29l/c1J7js4SR3WJSRJ8nJPR7UYPYuoQahUuCyHr+05dd6VxiOpoFhYzL0
nIgSgpQGVsx1PjEL4W3JunOYLlWWA/jhRQ1ynMXf4naObphwAdn7xSSOUn1Ms28K
X6p1BSsMk/oW70t4IqE3kzG9OrrzF3MyX3XvlINItEBFTGZnSLaITZYoMelBkAib
tLo2YXBTAz+fYrPlqV/1LdOs3U4YMFjF7xF+lyusfggw/YE5DKIb/2i667f7KV1x
qfS5n+GunESSRQeMVYShXRUNF8WKyYGkOUyOdh+z6aVdrq8cVih5ccqfBanpJ/UJ
LskRTKwWD/nJtgBd183CgZgWsuI8hNhHN0tlW46eW9oiRyUlwpJrfFMwu0P1HYti
QDyPJOZrtPZF1yfTMfMDFj8DBUi5WBy+M4/8PFEMT13QNsgKcWbXTBl+8MoT3NVd
TXCAIDQ7MztF9wwwFdDhImIBHl3IOAY0NTrmXMhcluT5kJ7LPP7LOIYq6DqwblvS
hslx48vE80jTgMVHUnT9rCxKuCqUybM7oepic2ruPdIUs2+nwMxAJw/K6LGyH3wW
PhE65ugUnz1NSn/7oSC5aXKhWzdnlHxSZrf3DYtHZMlyDjujpEncsQYKNWSnkaNm
eHEj/5NeQpNMgJX2s6lJ0axz9yxiBcbX8KpFapG8ABMqz2yj2eZ1HOz4KYydUIvz
wt6IwoUVmagJyD6nsrZ4PkxtIwliCu5VzjNPFxiLA8Ra+/NZfeDyEBpT4XNZx0ZN
qRT2lvY3HOeHdUw9wjUHUaWeFFLmT6WTrjNDbEYEDOjW4Y/u3GMRSoeA+C9ZI1kK
UGeNshlZQjuBsqNQlZH8ekaMt1frMqH/bO1ayTInYnv51lczhopUIqgB4yEnzjxr
7C76IKuqFfORpRXM9mNw3dtYtIzftKsMo1s5Vnptmq1zaw66SjJKNnZ4GErkSTZK
PgMnrkYHHGs+Wu9ohK+TAOI3eeEDVH6+xDhCKJwop+3lBp7LcgsYoyWClfqxRRvk
PaHJkUodY+plppQmWcHdzQTpGJfqbQbl4CV+KF+fgLawnjehfmApmpwhZ32htau0
LMACN7P7LvFc338nTdGbnl9isk/IZjYPN3IlXGCnLTRE4P+jWPhNsHtr+/OvAR2r
7KIwYhXTU28wBquY4OWT+wxtf8+RRIKZ1aJQqNTCuugWS/S/T7agBX3oRI1XnS1H
hnOuog17riY4FDvJ9dZue50SycdCIMtyKaD8KfryAWN795/w67daYeg+4pRV0cpg
/7Ab7sq7swcTYmLvVKx9OB0/nti/VizrQyRtVceSmzMRYHbDspjrodqYn//ErbtR
CpYVZqYQ6RmTVl1/W3eC8HsWY7Zl2NO8RjEM9Z3FtNrPfh8ILcgrHxN7qKu1G7Nz
leYELZvBOIyWTVf6aLJOCTeq/8ziV92sq8xroat4GXNUmtYRkT2qbM2QGw7uVrci
iE8CAvYoIEoMHbMBXhVL69wCQ9TZwD5plXvB86NmRgSRI8itx5iAwXlKJqM29SqM
N4DxjriRo7+RDQ9MT1ulmM0AHooSzqdS3zuPs8Jk2FaoLd4KYHVyiocJX0GRcqti
SVDT3n5pjb0OcsG557CSWFf1VZxBTB2ZVXCuvV1B9RXAg4il/fslGFQymGsH9O75
dNk7h2Nfv2TgIVpULgbTU1CkOznyuEWd+k1EeQQDIF8G+1XF0/bMpdr6Z3NITvsL
bOFaM0AZKNRRe2OdJ5I5Rb+p1KX468FH7RIfRzuoglaCwtHKwJNVUvzjifJ7166Y
kCrw7dHvCQG8bo+hF2h88njw706l62zvoBWDe+44khfYtM+LAiG4m68Oel4KHIgT
R8L9nHRLliTd6RkEyvKpQVAYGcbslo8wSQ3kRXXi7xlm/ihyR/C2F+ah1xAWu3U6
StxP0Cz+j8f5Jrcpq4G0kUKWpt1iOIPS57jiTrXYdmi8B50CuCm5xeyRY/kxHvb4
nIb+Ej/rW1dUaG3wMeS8OjwAIG4RBkwkEuGA8EI8YUUM7v7Wgwv1Kk3n6nQeI7Cp
u3u0ZXLSfpQQF2O+TUGO+lecq7PZNXrCUAQk3FYdI1Ny8kYk8xZwAjXIatOQXvbs
TT+rFBByrJwux2d+Biw0zwxycZCYLOCcjGPjLl7KqPBJg/6IzG9Y4sSEeTOhdaZo
XbMB+2nKjkjip+BpfI639CbQbjh+cVargn2SGvSCXY+VgzPCbuUkTESHQMQ8gJqE
69dOHULUIKIExqjJVN/CC42CCLX1TTM7WX5WLqtgnla+KWZyULLHvF9KZC5FETtb
eEjiUNlNYasyAB/9uO5KPJQFGe9zDBd5UwlX18GGYpRVj5yPBQPj9fA+MQ8tGvnV
hLmphgJnMbVJKA+m3X67jAQDSsaOOMs4gOXVVgKs6zoezUXACK8OdL8rWNTiMRPp
diQG0fOn75bCt+uGPaA21nfrbdF4T4bYEuT4X3y1VB0gPgWmFV8Ou5j+0HPlPe/R
WEU+vBcSsE6UpFh5iZMIcYaXQAXipk4PEfLDYjfICdvZ2zAa/bsiQ6nr9ixWK3hm
ZS8GIBzHbK/gOJ+jVsiOu5tsQ69RcRmPwvAvuGapzuNotvGaK3REaCW/a0+XClNK
Gcf17HG0Q4vpzDgZGDZUZSovZ/BKxDyezTKYp6HJwNEv2tcBOZ5iGhHOIOwSn/yx
WiRzlgkIidYddo86besff8YPCU2Rd3Wc928AYt/1cuOpWrOEn/V6ylXXY6ZM+Xlm
nBY5563KzZFiCva5HAmdzmh89yQ4wk5IRLw7vdo50CdrfjU7yOGWCzXaDtM9YNcu
AHLeFnpH5SVDuaJIpHXd/rGlVlkNkClvyZt2ew3JFa1DZm76u8lCOzsEby58vnuN
/NBmHV4qYgSGHb6qKhMT8oNMEbTHxFFDmudIW859fAgG2P52xNu9GH2dJnUtRS58
kpuAkYy8BZTrHE/u/VLV6ua6BFIFNeu7lrcXcYO7GYpSMidlhWSUkeZI/ZzjC88o
RHg/vuC+HEneJ/AtM1b0RarCy2Gv9OW2aUtEwp6p+B0eX+qIO0Plw612WFHsw1/h
to5J89mUQj7b5fz/65WD1ReFL+mIkRIsGlKauZ04j1wMefnOi8wwfNnnYY7Kf8Wp
7S06jAd4PnDsZrhZlqn7lmbMYQ5rnWzs41pBW/1E8761s+CAsDb3A05Aj2VmuqFl
TDKqlkKZTs4B+ZAfcTg89W0Z+d3w8RPX/w/n/SEDK+1dW63u7sVmpIwXRTFaMZlT
mKkYLVTW0HPE2IlA3Y8j0ynIV0ScKOrBuQjmirWXQ5pyrVI+loGxvGgwwpUO+yjv
jZ3YiIjxwhiZmdrXKggyDiMQct77PuDwqHQzrAXNTBOnkmZWTh3bWwv7efVDT5xk
autSSsVCt3uxTkHHo75VJLVgyXC0tzhhXdzBEtYi/uzHUNcQLyVfjJxW2v1W4ezq
G4Bs6JbR4rIoVeD0cc+u1pnUmSzP9i3S8A1ztZRg9WhcGYxbspkVaqaBa2Qv1KV7
AC/w2X4a552/D0sZf+QOuqncTUUW7giAerSGQg7gvhA8vxvFizQGvBeKql5V8EZw
gVUNCFwySGNs4vmj7R+kJ8TNo9DD885djAARu4rrlnuODmsV9kyChYXVnY2rYJnb
I/2DoXpWdEdhGiD7SWMF7BTvvtRUJZYkUR2oCAW+jqiqtES7fkLfHxuq7k5yUMk3
tfKip6N9ZwlUYco5Oxs9MCI0Xi5Z8qk8kQHN6k0rDkeLb8J80/mxfzZOliSMC/0b
6qom5tVHqO9pn8puKU2FJh9Txvh5JjTk+ztWsEphIBTjIvStprwp/0TvQHQUextg
O0GyhmVKOFfW6CMXd+imSANu2viGzsy9jXyaqI8S3C+nzoRrXo943SJgsM9G0RHO
6OlvrZEZcQ2TNWG1AImAgUxfC10TypiTSgfqhVcpK39RsGfcA2sChniAt4vd5qrX
W1qPrsiRnNP/ZS1fjrKQLE1p3MQMLcRwwE82E7ynQ1vFaKEEnI0R6YaYTngxrNDW
+T3kIw4L2uMiH7144VJAnZYT880U+v5kCHJ3DtwFvoHBYMGgZRXzBQK5wgUEKRpN
CRClY84fktNUTlAuOsuMTwifzUxs0IbGvCnbdq/rJiscNpeNPmr0npHJy++JNIqR
jInEnQ1h4nQrj4DAbYE5C6rc3fByCO2/R8eLRWBXCC8N+QVnW6K7ghm+s6pVN94S
8VaBoOXHSLT0mudO4GIKc8aVo+c8tAGVDwz0Zq+fFr+aBGUeCCx6UlO8NMBuohsM
LuGgqzk1O4pdnzY2iwn2VUiYJ+80fweDQbGfhXo/WCPkrfhhcEuKSf+NL5M+CUOa
xaQRsUEzzwlNxfOHuWQ0c/HnJk1yELXrvsizq2+BYhxAdnRwwe/vipm4lGOrRxfV
BBzovWkyEXsAnEVZ+Fidf6rTE+QA6jF4nx1B5hGT7GcF1+jrJlAKDka05iPe7F3L
ak7UQa84f34jKda0nnSGz5Xh076JBFtoSZ+Qyf7PzCWwsQmhRNDGz1XGPfO2AY0X
LblYFExLSXsEDWGoPbCLzAZeXSrk3k0kqsAucGxdF2CGnfV5nFdahs9zILNKqtjh
EHWi+X/XO/txZDs/taU+8XVWFgg7HqrszJkZ/GuOjoZiVs013Qg8ypXk/j9Ixbon
PM58mrMWBS46lVp2zL8zAivmxyYuiJdihJ5qx9LmjtHq69iS7pqRph1Ql/IguZEq
qGQY/wIpEtanDQlpGw7sVZHs/jEaqzUP5giJjNfv21XwfX29iDEDb6JdgBkPC931
GpshnIcI4nguw1HRetrMEwUlyX1LzxazftVlraYDfWEv/yOkV9sxPG+fZKFVkNzn
SMZfQX1x7Qnx90hAdICbJBIx2aX7NsJAYo6aF8xjQzMNT1wy75kDltDBR76j0XYZ
wcbcxop/VOjeNvNCI9mF+npmmiVSl/3aUoBS6SiZXHvQ3GBtHlDlipM1aBpXFF3T
IMj0aBRKupGhocoduEgwLK9nz1QUUTdeQiCxTesK5AMdpMsKVofBXRDAfHOKAAPU
0GFNx5A++/c7zJk7xFt5E1sR2Wa9XmWHjd8Zm18sM4fQ0Vd13B07EIDyheEi4HGJ
HM/5AwrgB5/dBNLV71u2J6VQB15elYPdBI8pivoQe7N2gaNqsnPFDrSeN7KR5Usn
AmcyI1kkV3YQqLaaFlrEjwiYBHsCySSs2OxbUwME68RJ326MGN+gvbBOAYT4yD5o
bVBoo6wyObN+/LxoljlSh2R9MZ+lKdLbXxVe4s368tThK8Jc9EKYN9HTCqAZu+qq
tuQ31I6BpowBnlwMrrQ8w4fX/FcfhQA2z53wCh5Y5M9DWYUyGziOqQI5ARsl51tu
6eSltqH5WoCtDc6v1lHwD0xStq20kYbsw+ZN8ZdGQv2p/3Cfl72mkV4SYcNHuSHc
iyGw6dQQNdbK0YVs8wJn3ymtxOEv24rWaQ+eRCjEn+zvIh4IbTA1LfdBotGfMvWa
CiqzvtTEpfpX1/L6hI2UMUeRQoRntKADGUWfvzOBWmz5GFkGy1nEPC6sM/HbXa1m
mmynA+arm6ct/B3+eItNfHUS5fxSOpkF+h/PXoXmEiTdQzKwIGRTWiKakVNqIL5Z
QTwbsK25jjBe85pkHk3SQ9NplltHIBzMlEAA60BewY0oC9O3v3njMp5EZo3Rx4g2
+XzULPMr8Quqq0vVAQAFfWuK3gOkYkQqlVIsB+5RESSEs1tpYbxxWH2FkTtOZUrE
EzE/JERtTN3mdA7s7qlA56XjViXNTIKAZSKzv8YahaNXy0jbLi50dm31AyDNCvMN
62kQpmYsNN9XatSFuJU21Q5HyqggFigU8DRCyjKkqPxEuaO6Ep6WhJYYEgbfnIXg
iTh341j5F5QMPWLWNIFCKe0HRWa4Omo+kRO/Rj9PdO/+jm3layXoGOJRgbdHaTlV
hW/NyQr5KLDw5jWCz7Dx9hrNXHDq1bxeybDLQfzqxn96cpXxPBHnTmkrcu6uHqTP
wChYbNsLGDytYK+xqjpre3uCi+R38kcwx7WAMA0ZpbRO/tTSajPKerI6qeedI/z5
OCfg4mJszw9mgOOO2cCyPBp86dPqpeMvysDjiGd9Yw2gp2MksGcfB8JKmbIGjrSe
E39RToDkauYNFCn7+wgJIg6nnIdAUn/HYVGY48qLt/27ZXiHNJ0wprGGhfQjiBFP
LJ4NUeYZR3tVIYAb6XEWZMZJCUNRcfSS4j8e/SkmyRDTnoO7hLJB3XOKKuB4pxMr
tjvIHEla2jxQ71uZuaczRNcASUSX6g+qTaIHIrzhR2HVkEquTK7GC764kxtquUIP
DBQjiR6TVV72jiRTdXOwpuBAdbDd4QYEb3Ff2pqSu4nEzOsV0lfHcYGhaV4yVNY0
A+vi010FKwCaQDMp1nK2KTmPkZFEDcrSNp3o1BXaAVVuCjk8LP84mVxg/0CnBO1X
YrJF44ByL4PIAaAWE+tsXV5mIXhat/QKoCq370dx/CxtLsvB24N2xqn2h88iZwx+
TwMnlpK7I/NPbolg12IE9T6st7PfmbmwAdRBuRJ5cYtTDLAjlWNH2pcvzbpVDir/
iIuheZjvNCvhkARTuiWK3xQYEvPXwNiDUmAIEAGf05d7F+BVWSXRr3no+YfaPzNn
fZh0tvdtL2ab+qxAmPGSnykNllLcczFbhENNyKcY7ZN6By7nkctKbqU7aLx90uXF
E1knPwuNJ1y0t1PDRqJm6M3+jWAv/ADNylWGRdFqR2BWu8zOlNBRvNoAzWtPidg6
nNfmD+Wti8WjOnYofkklg9vc3Oc7ZFU1JSPlSXpJPzQ9sKC08u9BZRuQFztBObCV
lvJqZZiSSFvZUGWXxE0rSGLMFo85EpUmWZvE4yTt3QbVNgbT9J0jAHk+d83HvUbJ
mxWcvmzTzruPNGx4kHDL7J3WYfJ98DAsjrOwN5tndnijAvsNYU0+PgL13hNh57TP
0vi2b/B+/y4Y9qi1DjNrXRD22+HyRXPUNJQmj/lWjcnEq7e7g2/igX4pZ7YFQ3wY
IB3EBpj11VFjAIxEAIhJU39G1SUOK7a9McPatt6C7iLibLL54rCIzYF8xjuGzW+a
bMrAoKy9vOl6zhS/8GpDOshcMX4x90mdPFAu+Bx+11TJcMJkvrkCmzSg5m5BJIbL
ePvz7CTfWkaT7EtgxjqwSyC2KtgifNFhtCz7tvNywoR07+EHuat3zN5GujnMGGRI
1JBncPE/+xBZC4rJID/xH+BgYQfLUe9e0rAd/1DGPpBCV/kT06OCVv3JU7wsPBrX
3GuNOlOQxsn+MGy0TqAhnI1FLFxYIpdBhDrAu3MnAT454HvhkEX0unDuTXdoTViV
DlXpdlK76qa+fFTPJRupDTSm5/0AW2rTbrMNreudKiTu+yplDatedji/ulcEIpY/
7R3sHQ+lXmSK+sQvsWM3YuAude4URPWYkFAviUEqeoc/kE9ejgJOHEniBtEMwg04
jwRTodoMxN471uTEcjCcJ/5t/Y2MjJhLYRBLGcmQydVIqG/PKHZ4WuAUT6JqoDfN
J+p3i3y+WCXLxC4axUAxOX2ePrTFe0jpzHUpdhpsnMLvDu6tYAKq2G9NX3hmL5Dk
Oaz7gvPTwglZv9nZFU40Ao2xXOg6UyziX7W07zKt6v6LZIHBnpA5xmurMQziPwYk
sPSsrqeZjjiygbc0M+2hy/KbSCJa4TyyT/BF919IytHE1LjtNQkJ8EfhCG/hZHzd
cc8K91HNp/hpRCmQxNEMikByaobwi4RC0qlOn5axlAU0BF5w1U4syqS16Ye5LvZu
XZCol2DGnfDI7sFY2Mj9gr7rVnqeJbBoabBRFrf8OfU4uoGgLXXvv5FxMpRN1hAj
srfmSRHvQ9aqp4AG/iWnV9qjRrHGyLBzqznjx1EuW73NUqPVnHkxA+6/dXNVpYvx
y6QTGL+XUFmraNASNgHiEiyYJspcPwsISefD111vqdBWppzdxNyO1yQR83XKYAm9
3fW/qHwhtNb21dC/glNQ6aNS283xXhyJDGlyWvbyVeZNDSKBosaF4Na00Pmvqspk
ZW2MysP/29TW+V5MSIELRTJR5fFLuSpFoJkVjRadUSt8p5MQwTjqyldMsCVXWY/I
XxGvzQ/ljHOGvWT2WZsmqCDvKT/vocl3vfJuT5sXwXf3lmpSZna1vOnqka/WY0wA
welJSq4gkfQPIFhFZ3SKBkjLcAKKAfoN5YqaObM1ED2X8wJIDc+0dhOr1lMllxc1
OJwsjewyqKEnXvqWYF7i8wz3h/sR2adiVsVZiR21BI1Kbjtb6gkulMLEw7waNRo3
fmEOVV6t69N2DYO4udIDBiXoaPMjeojMsUjgl21j7VeJW7EIpkwReKWt9LBld5im
q4Ien44RBrMFuxtPLcmScLiIhUcjr5C4FYbKlAWGblIiupPBnuXSstmBF1hvbxq6
NgLfGGqy5YKZevgneobBVFt0mkC4f2TSuHhIkHxApyKYu36jt5zzB5LjIpfJusgV
9wudi0o4JYzwRaFqCNmM7l+hL+WO92ZrdLeWj4ECrxPaxkMJygRk3/Z+eivhJv1E
98MPc7D2D6iXTwj5A7tuRqZnoYNa58h2rspFnGr/FWeiB9affjt73Bpo1Yikz8hn
K2xSty42cJLMdNu3tW/82/Ezp7zIPyNAlrlewsjv5G3i1HWX7AkhcjXLcD5yM7VX
YXxYuhT4wGoms6ZPs2J18Y/DnQ8ugSIfgez0AG5eVVgfpkeVgZmYSk0tBP7ezUZf
JtfWwbKjrq8RI9yO1tTMFVVKGXE0zLrv0uTrkiOyT0BNgbYXEYPh37zAREtMLHBv
VAdrPTe4DUBM4vJqqG18YVexY2G2u/obZmwobKRA3QfAK0UqhbRYRhSOfJbDd7xK
e23giG/GR9uSwo5HYVFycMgVlCkIFEO47y7EUbDUFvaj+PtGRFrIbbiJSAfFwai2
X3eZIl4Ats9dJmePoatuMAysvnB0LU6YZKa2+hoM0/6Ase1zb/w6iWEpaWAbzeZD
sSeaGdQxoj8HXNghBfd5qfyOxTHvC0F1fTnhpt2K5bd4cuzGdZV65Gghiie+LySH
LpXghPIs82B1h05SgCSnnY9HOq+I0WYQuvYQaBHYXMBUVV9HOlo3oBACOZ9lrBxL
ppUXThLfaC0bLpk1KGCmmFp5uEQpeFVFY0Qmzla0NPRUl1CqXB+tm/8yYJPrteFu
jq9nvlD04Ix7lyPFyP9qxK5WN3/Fqw57mr3OyOp7WQsFVtKlCRP+Ddt1pVbveXFC
sKNVO9EFFd0+WlBztR2ymx+urEYtIJhW1pZH4M51LLZrEwG1efOuYo5NLAity9hE
D4lVGTX+vyyKjPObz9YBF1ztgETWYT5CKF9TIQzBkn4uXu05WuZeuj9cpwU3vmoC
KBxUnFhG/NYqQiatCEjh28pUE2MMANCLsJNHAZalToS4+hJDMiKRYlTzzSdEbcyz
+Ij+UXopShOEv8zLx7tKGQ5sZ8/zhDpRa0bPRB5+EddcJQDnX58ppMLTrCb87TVW
AP2wI4vsrbkfE4x4EvBxf/qlEPvvPSAh0mkBj4pV4lgwtydBNQr8RMCe84x0yZuj
Mqwb6FX+ReFxAtHTdpRAVCElNVWl1rqG4PanwXj3+4bkaEougiLx7LgRs9AyEbix
GRQJSnvTno0ivNya2UALsMRJZ/hHrwrw8si1DDgwSxaSxnvYQTgDXtZ81cHK2Y0u
OGyTf+4jeJk5oHsmjSwTzEuiSNsxX7hIvleWbPAl7i4SZtFZ9M+GStQ0agY5qbyc
dKuOgGngV6jBpE5nC/eCtvZFHfkM7kMfuLZJ9srDEw5JFH8dDkUrY0EvCGi2buJR
sU2zIDy23VzuXWmYJ8roDMRmS0+As2bKfwYqOSk5HvXCOC2zqHKbQhSPaE7QMvDi
wHETTziyzIk25t5d0OU0TScHpW1HNLWQ1sCO6leYxJSgx3PvAzbi+3LKKJX4j3sB
20y2h4rnJI9n+5quhQpOKaVP4M71OVwfnRT3ttyOqsy0o6sdphwk/jdIYKS/K/iV
iEmruBXNvuk5CeE/7XNAODBl5Fq+ftn3mgC94QW8A2yxbI8CCye6sFnM3OqITxXg
f52Oe44T8b1Ku441cQ8Rf8RnJIbg2fUoT6WW8UPhCyPE3ck6FYWMmQCxNZ4IzhBP
xZrZTubhAaGQlExT0CsTA/aD3iX2HQnRbkysUTrneqxtW5c1eSwH1bby9mNz0vaD
r0q2K/ydh6ebWAR5W+DHDLNBHGctgLzYdRhGwxGmbK8XHiTIvqYwx+jZhtWhcqFD
04+GlYJAm+70Zu1iTO826EHBqensDkfUOpohwHdJIS/4KXONSX4t+UsBGCGHxwir
p5k3+HFHLuiiUvliKr0j/uvKg6twYjdYhqKJg1ruVj6+zDlKqDFNlHU0Zd5Opms+
Of4gdjBpdV0KI9dVKFZoxBGFjzq9yyXZn2NLU+QMAuIEQ14DBKnm4x8XKkxjog59
ARj93qNkx7NUzeWmdcFUDpgsq84+3sWqsJ2DfpA3XRGW2VX3is93PLUDlj5gryto
NSCmlduFaNIcOF7DZHbDl7VhcMFekRVsMkEW/nVP1sKY7ciIuxfKG8caQ8agDxxR
Jwtt6/BSmKaOs2/Jr3kDoV9dJUyUK0TkHjpJbbMbRr9GMKnDbX+Sg93+Tu+DQjIo
YyKMGCKAYTPMdB81xovEwz3GjeizzXPaD620QqfG+nL2BoKKhL+fRGFSGPdw81ER
q/wsY8bknyz+6Zm2eL88buH4x1MUOwkf6rrVfwtW74qt/bQ9B0YzdKmij6LFK5hO
4Er5bV+OtqJWO2FEN/7e73pm1rMqPWJprrI/tTUNgWk8fopbF+Tt8zCevWoOG7Ae
lK/yxZh4oGvywy1pbY6AN2osjNLMbUr5qRhmT3kZC+EN08gU+A0ale6i39sSgAGZ
a6nTkUpumzDghbdQE0twuPKXYP+bIyN+HPujWP6+yMpW9qZI4fHFQx/bnaNrhDGB
MTI+Jdv3wFFyF8ObQJheGpiXvdWEs58CdZSa3ANyRbHFbNSBrr8hwBClvyTimi+G
w0o9AYjRD4OpAXNVUwySuSlkXjOopF+MXmzkC0ik/TqrhofQJDbPEAUf2wIkaTmz
bxPseRsmIf6XotYE/3pq6BHIvTYWQTLz6vyKLJu9abaPL8iW8+K41RUOeg8rKaqV
Xh8G+LQCSMEVjMbUtYwJBpESNssEgiJ6lO1ZDTvY8VK4HJ7O4QCz23OlqtY6HinY
88zhv2F6rdFGT9ms0F0Ti+YzUndO3KjmfM8kGviRAByTUffgQp65/RT6gyXj1cH8
a4sHVIDthkNKHoHOM3ImPdMZyPkHqE8vHpY3Q2XoHP9RttUEfboSWb5Ar0IPSuXK
vYakKOLzLCmstowHf1/5CLZHTXiDdRguMNQx0iDOqX2p35vtX6btDrTcOhbNMR6C
41MeRBQq5wIjE1EYM1cd/g+686M860xXKNWppy5i+u4YKpoQp778HzH8Za3BbBJ4
dYDeXU77DjnhZQB0WPs2xJrOdDlrVW5Uokvq6RrZfX0TiVNx4mPXp4vL5C0rxIDW
GW8b5sMP60oCNCV2klC7APmUnNTYBhLMKmaQyGCRdb+ccsXKAaP/USqPiLDErj5Y
wf+lEHeZ+y8fVd4vloDLWjPI6Cn2ixrmz33hrswUJwy2a0nfjPQJVQBzXOwrp/0g
Y9BVL2D9hYXzOc+GYIH+Sw3lcVVN5mAGIrl3meKNpvtMgUy4KH2KIwFRxDhQa6vR
eiNnnm4FAFK+9ofNXlb7LQFVEtqIsVdGP03n2kRt7GvuIihJwW9BZDVsIklr8bpg
SCX3TO6vOM9S7uLSdhCbj+vpvmL+3C3fW87vRCZFF7hwlfplrvfePgf/zocNUilW
wGZIqlN8v/6D4DP4hHUgOfaB3zxcSDiqTn6ucoAWh+hq8G0TYRDcEOthk03U8Dmb
u2UQ4zTNiyoQb5IEOT4IDK/odSdzSAbyhpquaSGliaN2O1GOT18w11Kt5XCZCaqe
m4cNlX/riUDXoX6vJ6tjp8Q1Uh0ue6/5Skcww4Uq0Qt3fJI21KwKuhHOrpR+L0yq
PjbPK8qySORyaDn51RdBuyxusMKI8JyVrlGTdfr/AZD3Knk6EoELSFIvxuvPrik7
0aU6RH/MiHqwhYlsptGYFm/WFH6zRum4UXxnMegAKuEYT0KH6H31nNcYPSwpdBOr
QZrMRDxr/EyJfWmDqlsv1qfo5Iu8Mn1AAlWSwhvxvZzAYMAdKr1B8bnxppRLM6tG
/tF/uP785rLx+Q6C2+NdaoHbCVa+Dd/vXdaxQ/eTgbDCBsoaHdbM2b/mVLSR2agW
ZSG8owDI8LK5uxqJc5SPKKgV9mO/gOEORfdVjlUJLerAUE3UT83wHiArurcUPr34
fM9MlO4998Rum5MsTksOnyHga95q+u8UtZNBNhcxcEMIVNU/8puUezFsZ8D5VtPt
OROPe1raegrjNxl5WaMc4+ymsvAwMUFlbx3/tf0NqY3gdcfgJ7SmUYVqHOwqcgxN
BE+0BplaKFt9RmJfaZYilaxD5KLvoYVnOjv7PU2tzN7NOhArAqoQxISyEsVnEK3U
OFhYPT2RzFzmfS9amr1t+YBfdVPll+ZvbaVE90J9cZ4sSAHcSioxFvyHVBg9LUVs
BBNBr1wFrfAKXYZaboBO5wrNurz3DuAhF3xPMpIR0QZ/jN51fdYKAlYly6coX1we
uD5cstKbMhNqMX8c6gE7GH//IizKeNlK1LcPfhZcAE6y9dGQk7v5qj/CUy4rplA+
iiT1YE5pkfeP3R9XlhXVk5Feyu4repHr5tKLwqQ7KfJo8/RdAVoJbw+mwSeJyQOm
a1hUF3bdA3PWLdHi4+i1ftt0prPIqtE+PAh9wtUQo7gatWUxe8d7QEwTiwAdADWe
loKubjpY5CAL1f3PZZf1ars7eQT2bX4kBQ/xkLr3EQ8fmZP/xJILnMHF+ZIyH39f
zTFsuurlAlmevBvD9TFK8WL/pnDaritVuv5jW4yM3I3gn9OxVI3TGTlfZ8BOQY7G
ZxRlwPdhjSY5tWRbJhqm4ri6gRpcyZSP+H0ydZ9Qnv7b3KWFxlE8PjrRjAXt+IvX
jFPJmuEerCJbDCnj85llljMYegvUjAC+Ku0qqXUKa0Pq8sA1KhIUQjokGKAE7ga3
76phWe8DvN0wywTIeClR4nVfBPavhMjbZFhrKx1pjL8X9rZGp0yR6m6D9Xt+kvdA
UYtrqd9cB2Pks1DERKYugbYqYQJ506UZygtu1KGnGiFX2pCJaSnsNNrLFTc4xiKn
JWHXBUFhWKKIvGvi04EStqaN4CnAs6069KH0PqvXjrXuMvVoDfkOwmXATXtg2nIo
Pt1Y2RNGJ5xRLVUo/5tu5VIVIIxocXL29s8SHl7qNZEyOrRJPXLkKVGs+xoiVs+t
QWWY5QOv3bYU3ybBf51A9Ii3JM6xO4S+uRjagYFbl1A7V4EmlcQOca73MoR1Y8Jd
Yin9Wo0YthM7SXK5YpX0KYXV2s9sULqIS5WFPtFE7DWYYO29R3way9vRstr3R2Mr
ifeaxe5b4mMlE+0NfNjNb+NjBkPa1/ltIPezeVG1wuTenW3TsD2d3gv1KCya44dO
gbqNyDr2uq+RVTbN+nE8TclzvZ5dSg4/OCG61b8lUWnM/L743jHrN+e9/b354r7S
9AGYc3acPbUpN2SpoVcfaES6Hlc3X+JnutTKtvnFDqY4wi/dvAxpnO2G7DrYdpmv
BNQpww3jk8NKcsz7LGwwZyqM3vMmdvm0vt6DgkjG5GZ4X7W0gWSoUyAGnD71/hIt
vQd7wqacBqlVFKn3b2kIakFxm3Jm8f3ElWSXWM9iflC0x/sGI6D4hAy1jR7yqgxt
EHODre34CuinuDm26u9vIAk6gFK01f9h1a6aLvbplOfotY9bF9qR1pia7PR72KSb
o0wZRw11eupTg+BjJNiLSf9zLsm2vyD/lmMPRQLG/d2dtgcbDUzUS+zBY2+rrBAm
Vmb55GXngkHcY7nZzNCNzYuoNlUIVCxH3feVYhVltyHMf7ZtqW8Uxz0hOqxzRP1P
8JzXzoOcYCUNFppqT6Y9GdXyj5E9qmg2+I62A+QntRvcDU7YON5F4lMwbQ1GWdeq
8SajaF2ymvRALNdOQlOeA+fOdCZl0+U2w241kjvqEWkSPsUONhCAC67GQzyUBuTb
kjt30zIwLkJjEp6XC6jGIb1sOxGfq9ShvQL/Nx6X/l/r16/+9i0k+I3i67Ts3rus
tbqsvc3hCf07NUWcLI8/2faB1wjTm/jb32yL+mCq5yZyPUUb78ojxXClmIqU0Bu3
AlhBjZgwfagY00S0uo9eId4bVAnrRrKmx4Ja1yxeUtTjRIais5iDv1ABKpdqNkWy
GJ/Aj64IRxTG9n90fOq3j/IZWjEXZspm9xaIujhK9vFAzwHKq6VCsXQ3DarXKyw5
wiWbXdjtT9nVcxqFLnTbcx1PlBNXrslzd0lTpHB7A5YMnAKudG9h60ukfVZLw7p5
AAT8yxzbs6eo3FAy4TLAQJr7VVFEii3M+h0+u3ZnU7NjRl9Q7+nnxBxgoZ+AG7Cz
/rBA36qywShVOKl7Z79R6kinJ04v1k+1fhNSCx0JoGzfP59TOJ+veRQMOBZ671BW
dJbQwCMFm2mbI7sesO4+PO2Va1BrxgqNiuKdcHpzfhrxlMSCAlzi3IHWjdEpE/df
uGDhEwdJzSGNCq3/FzoUoz5iiz92ovyet3NvLkyaGrRyKh/j9TOOdecop3j9WU67
WQ2T4973j0ijoZ3U4wCR+LTvvQl5LAWIfR0PVj+SNipRQrrCuZAaipQm3kZBmznm
F0GH4kFLtRtCLdlThszQP+3SqLNWzsPvS8S+3sCXvqdGZj07ky9RixxMN+/1WFwG
Nz/4QL19nhiPsHnZKXdNnKQU40QJE3U3bAPyxbFjh8P3fZmbt1TuFJoidgeoVgGF
DkDZA57VJBNXuGC7qjaJtvQ6vgz0kkwinslcD/hafeKaraqMlHLvM//A7W1cKgZZ
n0x8wVetqT48vprmOtzsCxG0wdrX/mN9TDxDV97fqIKA8/i3UsDyWDsIAcLkAVT5
1DXAoYlRTFqjcbXMlw+qB4nfuaUMR+wPUYDkqtGIrMgJW2JDeKeFcSZltqRCzIKC
MZZ34K7sA8imb4CijKwq7l6Z0EeN61HOAI9Pmy2HWyn9XCMslxpklcCYPlNBKGfu
0RCx7qGDXPVztItKZTytSh9RJnhFnya7PquUAwbtrna6cDoZ3uzFlaLOdanKUh0t
ie+sHeheY3+u7quJhWsfDw8bX8to5QtZ8okVCkz8ka2Bo5KhqYAibNWY5Q8AaqyB
5lendZ501ITK2AVMT0OpJUwUKIqH4ZHhR6hOOIFFqU+YRWEkhLf67pcrpk+WYvry
U9ens6XGjcwcCNPBcHY2/RfLxjR5ULeAzPT18aS+M0O+X/cnMhMeODdzByyUojOZ
yW2ZiWxRY3CETYd0MkH1B95/W0AaFejZ2Azb9MytIlVBKGHB7dRupHS3RIsu+BIN
pS6mKM4fYDWBcSEA0JzpoU8qUuzr7AIqbJQ5Zv4a95obXV2yKkzrU6fersI2aMpT
3rSumH31OMegllsud0qmlyIqoRhnygWoA+JxOa6MRi1N8aXynHDrafJ1jcOhVkLa
1Bxkzan4NypbTVhZfgPZDycpKZCiC5OUSE5MTXPSfIBS3lYNcNFaFetvZ4r6D6V4
C7LNDgC90cYvXHDLJm+dsTcVYISJ+5znWVY+ijT6Hj1FEYVgq9O3Cf7VUci+25Xj
1nbtbUhgMZNmz7lBprbhqrxBvQOsb+QH69Z40WhmDoqGPV5fdgiYv82Dx2A0nvBE
rKRcmSP2G9NmiZQEEr9QlJk1tDqPCR0Mp6LSLlYLFgMiYxDSr/ZNI1dNdRWag2sQ
xvBD/ynTWqCZ1pM+RPvxawfFppXPGtf4Boo8KN6BCrkLjl6bq+FWBnMr928H6MMs
u64IOQgsHNPYotoEWHi3Lr8fSwcwOkcwm8sE/cgVf8Mf7lQhAQjlKav4RGnCpycy
eUQ8PSdyMeD4jPp+N4TQGBC4AbSChIghP3U5xg8gj0Ursuu3IeoiFBnDsLlZ2CbG
uv/rf8ytcWa0z1hK2kzS6f9+r04BnXY5iSqGrVxvLyPxvUesIEROeIOb6oHkBzKt
qLmTUvqUnKHrIulIBJCht8dhtusIfVal4XXI/3WtM9EZxXpsAJA+dPCt5W2yz2Bb
sC2zJ/MgvxfmeWO93WMmNYQVuYwI9Lq6LN5PbqwXG81xtedzdFit8B6s9b1Xe3XH
xggdUlnR1Ra8lJS8ECkIM0kRkkvdD/bTLxwu8hXgBhP3LMMrK2xbc54E9S+ZuFHI
g93qyM3f1JfK5SV0CekZ3KsDNiNbM5JJR8WMTgdN/4MHl1hpc1AxqlJxCj0hL+f6
FHJk8FPgX2PnloUOac1BzV+WkH6zTWkVSRmsqFAeryl2Z7Er0axGmaJhpH64jUZM
Psrkm0En1ImwErY6F89eeK05rnWLMHPx8aIg+LiFhFLZpw70/T3K4Mlkrd7w7hZj
JDy/Yac94RA7eG/cN3/OZ7sjVuBvRPP0ac4wGMIWrQ+GjR31sd9e8dtXHBykt/Y5
XlvPhRHlWlJTIwZe31vfm0kS7S7hj8fViMLLnkvOjwl9CxzjOnmTJkr6BHReSZww
hBS6OO3g7BbJK28humcG0oFCSVSELvHOMWc9F4EDLiudkA2GdI5mscKS7OuMVqNS
3l5vaaorjcA0zdxt9MMSU+81sC0OQBT7psAUUYwz2sSNt5qWDpHkBTT2U7ciYyYo
qV91WlaYfoLVjZ2VEV1XXGVHiNqi6qybfpR6I+zCnNBnZGojhDua/8gvQ0AfUYDE
1rQBicZeVZy+yXia2wkYfS+nVVzKQBWrpXOtZmJH9Pno3E3qFMvoscebDu8pSpD8
EMVi8xjV4f2QcKrrA1xn54qSy4pkmWEGo5sVwQgSPS2BzPN7TyxYfqokWabGuimZ
x2az5DGsnh1vaSR9VRsuZmpE/1dnMnDfw7bg2bRL9CPXBAoS32r0uGDbCnJMU39s
hcZntXySDf5IHAqsK9KmydyN6XhAkFG0bcr+saL3chR25UTmOz+j6G1wEFn+iS7p
VZ5BIhCVwrt97Uv2kkcJKA8WKx8UTqxgiCK5aRt04BvegyHR+Do6+zgFppDMgO97
m4wswlBuD0laSxBcRBYNvgzukptAI3VcuP9SgOYK7uTjTAo2yYASru0apXg9VHTP
uHYBV4kFrAgJwr9KEK6eRscrIL2MZuSmAYyY+8/KIia3fJG3cXV6z2+VTsgIUfVE
p46AIafgtqs8f28/jb1skJ39I8vfgD9+WNb2RrqA7+Ur0AAB2Yyc1wDKGKiHlg1h
LTVPGTbuVM9dJPR6A4G/frWoipMEYQsRMwetFDab3x+xTFY6Bl3yk5FsEWWvWW2p
diUtn5mbsyAe6FUWo8dLrgtoY2eaMdhpJtzar/o5/P6Pjkqd5H+zfYs2KgFA4T7b
IxCMiwDniWrF/OzBezquF+jw54rg3IAvzsYe1eKVBIU3PsgPFrtGjKy+liw1Cw5q
2QIRFpz0Kka10Gx/7hGpqUpVAt9uAFNM1xOZmHNAmp2e3qumnIgglvB+lmNUKZLs
tiCknH6k9l4SsNbJQWk4HPOgJTeY9INox+Hzik1RST0UZqQy1NPM3sFJmyUIOLFQ
OuRu6HPxTyK7K/irUJfh+3VaoiaDbP/TTXTLJxodTU+UB6jeg+Iu4rwW33nCq4yb
LFt+qKbh+lA9p2W3Ja1XKBMp+4QMdYa4AG4FHMMzjA/3CYMULxbBlh/2sxoi9EZb
7lOuXpyVxyRo6E0/xB6jaz/z6YyG+NIY8VkFPHmVGwYNcu8BinSlQyEQHUsdGBSa
7WQOu+RELXJkUzNDpx5YoJfTd3MtWhIGguSBk+dT3GaEr5G0vpXUTRQ+iulZNAP9
cyaSagMBF06+I/lcnvcITlYUw1edHxtqFoh1jjlLjIPbX+ow/822kbp9fFEMLsWG
h2MEzUnj5EdYZZXGhF9GS5I1tgKLr7nqJ7Sw5mOlGqkXK9qRbcjcrBJM0A0R0vP6
5C++korgxXQQ2GgmA8ERtuXlr9Z42WMsQDxEIojylnHgKa7xzfZcG6R3vendokHl
zWRs9kqsIxLp//bS/Jci0lMKp9LopBqhulIGxPxwsvtRn/BkYRQFDBSOyqAoKjZf
ma/7ThIYK/z8pibxpJik6QhvYU87AeDccKrSI5783ztV70uc3LtIMZU6ZB/RMuaU
H8FB8mH33H9RCdjLeyTzb+DY6q/l3ngZaxtSOZdSDn/UBTfmUSiuhijVWWNbJmoF
Ke/nuep89atfP1QLGtkBuxzGx8iAH0aJZCAsMwxcsEbggldsorQrcX7jynWR78Vf
JmpwJM7zy8dQGXpznxdmd8wwXmrjwvhkxmurFutZjYe61s1lu5InEk13WbWVgBce
65tjbAUrj2QXEeWp8DGdkEBHDl4DGRK3ZJ42W42cFQwHXxDsJQXuhBTu7SLZdSaZ
D+OAPEQq1lz91V3P+bSXY/aWm7aFQ1r9VYTc3hqF6m/U97xZ9uETjDQDDCA4gwtv
TyzHsqldFDbZhYN91vNfDCtd0cLMa8UQmKS0dTKuMZjlIx+DB+Wf3NWgJHTnHkfF
zPsBPPWpdJra0+g8rYNq4Q7qZJugJ6JcWvenwD4tRzsyOJI5FiBEefcBP4ELLAzu
l2GgVMtPOqn/s74FAqZwdBU80SZK7EtKVVccRoDaVxTHUmWZ4XmA1jAogqlKN/hu
aM7ulvkbx6FhvJK6UEWV5b+kgeLvfcOhl0e45xL4vWM5BwvI028H92J3UyUOcDeI
bK6K3XDPs1UugblZLQVf5avX0MOpPhgHsp4I3Wv4X0I7lmQ5S9G+SrTMV7JgxcM+
vJmoElvVhM6/8PKwassLSt6px9F2/jlpVvts0n9fz5HdD36hYyVBq+qwDQXkwGAQ
XLa4LcqnwdcWtSKO8K2xNJp46H8liUf9MYTkoCKWkuXl6sIau7Fhjlf6KLWjzocj
O/LGwa8pHfVSEf2z+rAL14ezXgNSWkq/7vv3M2S3PssrbXFHxiFywD1MQuNrIG4M
58VkElHApx33u4jgGqXqvLdoh7wFjztBJ9Rj5hL0VkY6FKvwc3esWWopr1NGo2Yz
2Czk/Fh/qg556KgeGTapwGSw4sn4vgXwxAsiQylfwRrF27j/5KfVHChhSsLTJLAQ
OBLRRJShNfDPLFFfv/ksme+b1yi+G/YvwOWdWaTewIXFRLYn8/P0VkmhokvU7cIa
X1A5Pcs4f4SvZbyVY5VO6bFXBHxdgcFhsAG5PlH/RUtgY+e6lEB+ecFvzGQsqLLs
l1rMRXhpxw33TUuIKuxSr4zHgbdVB6oXlWHZllYOPgclWBJZUtcLsDG0jrNewEZY
RgX8rCyiri0+0HtxZd7o9/km/Rv/0T8zMchR7yhsJiNZy/i8rjQxF5glO/DDHLwg
c/vaAhzP1t4Um8v76CN6uuu1zcW+VR5rB6pMQUtXhDRTCZT9MjgPs2dSwUF9InL0
hsp3DR9fQyKxhWl9l7V7Cbs+28oSYc4FDL8+FyIcFMyOK5mIE41QSIMCW0lTXYrS
wLqK4kIdxPpP144UBaSp4W78bhFHGq9Oqc3tA2HDG3ZDeEi7YIBHXMsZ2qYgSFsX
op5nuKaqCuLP3Z8nXeXMYSNpVPygySVhLUZu/arrL7nAQ39u0cSUqEddFXKUvlxW
4syk7Mpz6pSKWw3PnpkhUf9FVJ4J80x16GOsaG+LoWnvOVUa0fPJwI3KDQB8QqFa
lU7LgmYppa5ilFylNo9AmmsTX95sB1SHcMP8+iahLYnCwzcanvAirps1nCWzpWoU
v7A7rMrKfsoggxxS7vgAbyr4X6+mkSHV7HvuFxF/3CdefmIq47LtADLUmW1e0Th4
pUNNZUtezy8x92Gc5D2v8WLX3nl0j2Ogxlw4yNATuFJ83cGwTLqCFYFs5w9dU4CX
Md/eaV+1Sq3vSKBCgwAdiCQiNV/EIgLvhJE7YyeZg0icX6ufn0OfanqRCkY7LBpc
u/B7rMIC9bMuj8BzW4Kp3hDhSrKgf7BvNjvfQfN0lE85BAG89wgARJR/5bPkGTJU
/wkuIeigxfmDre5ioHTF0Fe3COfbD3ISJQ4MDzKDmcdNbGGFfUOT34KhKY2TF1VU
kyjo6l6uwlfi+eRstyrCG3JVzpLz5keIFH88Iru+zNhfH0LjmXr+9Zp++M7YX+ro
dnNJ2AXhvCxTV6yE/6czyf9Pn20Ru2ja2e2/LanoGeYvbalUx4WjYzwqcW7uJHHW
mUY5fvYf2dD3bMBSGXUs4iuSr3OKoajh5JYI0CpmV6iYRJ/RW2H3KC7FAoLyuBr+
J5Ysa3YU0aE84eOeIh6lZtl7/yRgzXEndvpRuzikABVZmG9ZAC8xLU0graE/Ik4u
6IMnDHNhZiMe8f803ICfkPvAJdBQEiGde1SHQyFO2GlP3R7R8rdAToFiK2c3PL51
NGv2vjH2FU6gsj6HZPcLZ17dDvPhA1r6THj+d9DZRc0GVZpb/NoP2fqYUbPQ1ubA
RNe0pa4cYiNyzvObasNadA13VFeVj9SuVR0eSlkDYlP0f5xvL91jNxFGCQuR2ukd
MKvJTCS7D0k8G8YMauyRNFCPrE4oGnH/xIXaFs02esm+9Hf36Md0Q0sxwfa078w3
tCsnyBIwqqmm81McwJz0Sj/8QJQWZj7VRvcfD55U4Ug+XMpJ/TrBvgbVWNz/KLiw
7F8oEMkxRa8IAZjTplK3DM0IM0soVa95irmxfOG/dn3UuV1OD+8zxkGG0I3fXGiW
QHy7/nKnJ96Yn81XEMlmAyPx40QSOvpP5ZkWiloulj3tfG5BwTvTukPBRBiFeibd
XwKqRg9NssyLuaqR1wt3fkf+F54756wufeu1pybb5bvhPBQkFVFJhkmb6U8NVTqk
ChMyYNtTPS+2zfyUQtvFOMexIZRoAyNzG6C5h33KE/k00QWgE7I3RG39oAVLi5jq
mfvKw1/rrnMqAPoDWQ9Z3b8f3OrjRvLJxvVmYymiFkLuWNRMFj+4Gdw9lt6vpUeX
yZRZ4wKOUCUDrI/uqk8U0Yoid6YKhldnGP5jsOa0SLdBRcOLBgsPoLPA/aBPa7oZ
t/yS89oWZygF9rHnxJy7QBwHeYlRpJFasiBFSCpkMavPKgXq3v8m4eNC8UBBA8sx
acvVqnyghWpw+2lSYyRmEHk3aBKudzTsLW0XxJMqXj1n4hsPH/wxgbj54x/yeqnP
spqUayYhDz7f9HFcNy1uzBZ4YP8s11xHsbnsRqIR6koIMw+6BT3LQV//Pd77SO6n
Plf+aqjr3KaCkMCeAcaghZGZYUwi6hB1Sm6h5RveOjS799ySvlNIAC2aMKukIsS9
yurYXELBH5cLc264ewZjV33duI3B3kQtOioQoCoVhMggm09YCLBEANk1uBAnWqPs
cw3JM9ZIw1QY+uT1Cbeyu/fwf5VUpE5I/nm1fHe7I62ntR2oifFudcTeWoE9hcgO
OoDOxmVb11xOnBdJo6dr83sd04dVSMdBhZ3kVhaWepV0uBDmZwLfxe00AbrJz6Xc
kwogLJYO6oHTnGqYdxEDIg5cAVGvP8o88eB9Hc+Y/wbtwmaHB9HfJT99jd8MU14A
Y+ixJRx2DbUd/lEwhVih4/HSE+yOc56N4s85QfixPuv5DwHbU+RdHAEvvPBs2kIp
hyE+keh145dgMckTldsrGOhr41sFJNu0/y0LBZ9h8ckkwzFlkd6sG0yZxrNO241v
d/gMBXp4IpMKEj+vWizX9B9GKJZzdTvOnOa1YF3OZMP1DefhwBvEVJHMewB97t+e
ontkJvLVKUrpnlCWhl3eJg1ZYs6lcYDUyCHAAtWEQYDc+5cF2S1kFL5J1wzIKqld
/gsnZxL2nYw1w6asfLcDbWt6EM6L/XOkR86alfrTaIKbDYgHA+yxxteVBnsDa9BL
QQtHMeV3KDgz3BKRxa525QdY2gW8hYPhdGy8qQADE7eU7Rmfb8wSdlU3cpnRPzpR
hlJPBKiafkuBKc6AXN2gxDxN0tiANi9JLuHs7MIlpxKCr3F9WbrElJE/Fn8Qo3/E
TsrePXxvmoMLLX51dfLKGUnU/oJpJHYeaOYmufEvHLJ7AXVMVY0AzTNe/RSYZlAp
4r7nF+xSHyNaGiA7hvPhAHRzDBJYJBeANhcYvFSuhlkXODerLSiOGSdzTrKyNDZk
J4s2EbCtjA4Nk+Vx6QmvJ1XBxk2EAIShojn18pIN7oy0bUZmJjsXKxJzF+AdfCw8
rYrcs+M2aWcNSwv6clq35GOLSDUbJ3Xv5Bx+/+262m7o6nonDyO/hsZWITpadlFA
kabpU3+yUT3lSc7mjXYrOk88co5+DCwwu9AOHMNzX/IBnSyXNh+Q79KKETm82J5U
gb5Nsbq5+/eHDpObwyBSM2ZCWA0fYUSAA+Z/wCMZTL7z6/MR1ZhNUtA2BKp/MVAj
bYXfVZ4Wov57TGQ9ubF5iutxj60bpO3qOp7LaxO5b3e7zrZCMvMvPn8xxLEsDM5a
kWshMvpfiP0ppMHyfdys58cNmW0bPlPPxM4Z/AagRBziydZmNYiQBenxJyC8s5EM
euRaaugyZjQ2xRGYSJRsLO+VAf0sMWa6jCkb7kgiJDl4HncEGQ2T5QVg09Z58RRW
CtQYwYwjFciobGOvjXeGki+w8m0WrBBT2AkVNFrf1CTvmjGijcFeEyuxmlLnfh6Z
zExpZIoaKvcS2BD7wyfw+bK4OaSrxBj67dyISBhlfpTOMZIWcAvSrZgfBdtuqoOD
/UCjbY9siG2dBvHTxEV6GVgaRsqxC7wocEUjkHdCZQvY8tEZlL+ePgjEzifJf3JH
c2uwEPvZW4F91Q8LvrSgFdPF/2A4Bxqz+1FNgIIRhifQ859nIfiThmwIFsf7x/1k
zyhY8LcRZIatc1lzXe51mSX5cORJ5Rwa4c2miTiwbCdDQJNWowrGycujf53hua1c
snAMp4hv9fYvlM9tVbrenrPJ43cUx4BtNZ87Iv3SQXTbzlyeyCgBpIvH7Iqix2R+
K4g45iNprcgL/xmWbKfd1NzbF5D79PPvrPX5ibX+iTui3hFSPgFUC4BDzazBX6RM
LRVOwRMD4OReqOgEVUfijoBhKIe07DtslmdNGWHQQm1P6b4Kf+fulY+9LF7ylb7T
LDbXALlEDDmkrWk4Xkf4ssqpgFXwHkyT9n7VJ1DbUhi7SC3bkbQCOY7xo+UoGDyN
EMAFmZWnMlSlR8Q6bTYBzlUxtodTzMBlHLHwAJKyXA5STxBYXzELCq11YpPTZKw2
kNFKnXMEcCfeswXRBPUXxpfmrF3fqJxef59XlavWvEPDcL1dn/Rv4b2oSWgmhief
AXIxza8so16FJ1IUI7MdI0qltBfc7Zfj3WxyR3N8On/ZAv2HcGW9MUMl0lQcgDK0
Hiau9OcxxZoXLFLVUx7Th/DDCEFr9oKkecaL6I6Sj3nMIQFwLmRhvjO6SIc68Yv6
Ht2sIXbj85ZSrjlyTmtsOhf8gB/3pbNp5im1B/nHsgzTQiyx/CRAZF+eXVYOiXYD
hj4rIV+wsOHU/PqA/FSG9y6r/K2iTPbPS3aAGKHcDSBYB8x8sfLZvdw7blN/h3jJ
J0fGpPYDw3L68sns/wz54ZzveJ5P3xDv08nw+T+0wuWjDJ3iwPPR4/ftesgVO7Mj
BaCiSMrCKLw3EQWA31GeiRiV+8tXBsUoykWPq24+38maZvaqYFYXKgvUQTbaGw4i
H5nOizkqDCs1sWwHstbvd+vlZZfmuFf4voKCVYmovn0IZtQ31hnERXtRyfexc6BE
G6F2rJXdh0y3ryDaqGBmyhUIcLvTzMPr+9YKRHVSYWHOF256B8Qplwuh2b9LdUeH
xgcWH6/wdbXkQ+/jZ/K1nlpC9V8c8+HZfOdQp31GkLOCUHHca6Ok8wzL5t8EvEhW
9EFqYSiDsxQFM3JpT/uW169Uc9kvxkGWgAQUOlmqN6qwoW/sHKSkhxVUX1rPbXCn
ugxDXilncxz2u0+Ci/lUbEM3spr7ncguNtOZl5Z1LIoRUXwYE1XPsPjQA5GYiz9l
O70Fs5lktgZBH/d48MxKiKzsNMKHJv6R53hNf4Vfr7tJvSmqzXiSLluA9EJ3ttbk
Eys5T44YbKeolRZg2wNPElNWWRRAQA3R/mVDPEhK9oohRs7a153hlNykYDCLkEga
ri3ASDoB8UABLh8ZIpH+gHouzS3JbUDFO6sB89U9iDuPuAEiFdqr5v+tI3kXO3cR
I7rRxX95MW3QVWah6u6F0B3yMvBITxtlcF1qpakndPJ/n53HOFUd7ECUYauosrlK
Ben6xktjLt0mBR56HyR/uzZDnnRWf7qCgF+iTG0V5kRnYSZ6kVMbJeLo6QR343BR
9wBE8zpam5qecwioimIshk5Gin4hF19rhVdBHFoDNPiOrMMRbOVnT61vfz43Io8P
NXdsN20tL9hj/a5NoRUFhOlHCn4ydP4Q1lPi3xxMeGliTx25u1XJG3+9lgbNhOw7
6R/fgoKymjBok8BZQNBEho4DL430VieybvAj4enCbaHxqqO1+LMmx/8iZdCBtCQu
iF+7z3fjKm2gA/5i45P0q2nmdFZo1BwZ07iH42aCNDQZSpSTTKyhzOYivnqxKp8Q
d+U8HIIbEAhQ1uGpKJts6Ft6iD3PC35wEVRr6h0pAbzRAteLsVGSbKZ0fQf8QwUF
jSq333yjU6n5zyK0qkwVD6W5jg5DOp0UJa5EkmgFk+DK9GByM19gzURYi7IZvjvn
Vhu+WaxRquQfFVtDF8gPnLoy4XGcmu3nLGEr3X9edT8RQIvnqy/1BqaRyhvg6+sh
zx0amxhTaQkboVCQJUMO1qL9PWO6PomaqVMThzHWWU7PJrl5dxW0vcpg3EbP2q0Q
oweUObSTMswB+ClWfKArIQwRFoJO+433NSdrydtgTZVIs4NFYz2fALEFjJYil0GS
6x42ljUkBdDbsmjeO85CO2Z+9bofKm6etGD9cB+ohH5GulIrdgBkfhAIbh/ENVKC
9Ef/dEuIdegPv+Y6GbiSWa+IL+B6/6ndKGQdC6QPls8q6s/5OLxYWsBgRPLJpDtz
NgMGuTn+kgWYRD+yEzGtpx+T5yfiieUEnAITwxQppzwKF2v+5/isHfBL2PWintMj
9e7xHZviajPQx6zQmLj6cFtY4JvOSjIgDx0c1nJNq50MD3VPrd/+WZrJA5b9Eg4o
/eQL2Gw7VWr7pipP3VxZiy7n6EFcFs6fIdU0R7QfMmNhWpTnKAxno6mgVpVN/zeg
Pz49tCk1ja4FdZgNrNS1iCBR1naWJuqkG17UKgaX1iE1pPtJjnN8kep2Ira+4lys
O8oj/MoRnZFxYpcU0nS7M0wvpiWD2MBfUfBTHoysTIjOPlFX5FLxioKWiPBC/Ut4
NEIS90nv50PfkmQzxvBIpxZkYmignR3w8tz+nDHqX78RJbvFJznAektnw0/YOaKU
OkezihObMFlT3A6dXa+MUTRydGiHSsvGN1KFphVisgLIVGXG0aOro8W230xbRMGh
7cPprdAMp9G6ktPmzFn8vhKJvhaZKBD2fWXKtHIiaMukauTmF5ih+dD0twgNT52a
V3eAX3i+Q7XG1dq5MO6KiHFZMjwq+dxZgcqHXqF6XixqkBdTCeubYKgtCOlO82N3
JA5odvQXgV4c0MM0c5qdhi6lme0kbNhJ4g79f9zOrwnRRxTscvRcz+QAsZgM484u
OfsBAMCy2wFEVrWSUOhSFMK9kUv+royC5QFYQVo5tzUEYAY/Lze3C3rpviq4VNBa
/ZhrqP3dUDckZ+Oopej4GOS+Nc5uhxu+c7LMht8Whz6OXyfNjaQEUeivuYsjlHgB
35+m3aj7x1DnYngHaKzMMk16vazCogCNcNgKmu2oLfdoMWnujAGoQNp1zqz21IGd
9po57vNAwWKyjVrAda3S5CsLMhHTJWup/IsSBdQBsXXngLUPIsfuSc5rRxwCnWM8
0YG/1he8V2gp7/ZJa5QLOSN+stcV1/BPq2LdGneJRq9xl+fC7cxraSXAH2rQRG/V
oWBv0kh2anNnXoRWdL2s0OawVPAMQhBzlEepTjw9ySAYRjh2nybPsicHncfTyLzG
DL0vEsStVtzFHgyBpCDIPeplSqiHlJUqh9GpZF6+wdHj51J9s6hpEkRn6a9FyQDT
sVary2FzqXa3eQU/v8RszKbt83pZvPsAL24YblLy50WSyl94chF8TEZwBPESQrro
5rP2wlkgEK+2gxtIftm/YX3psLw4LWdwNwUowD5h2ZevrLOygUUd9xijyeaFNMCz
3TMHWTX4ObSk2hhPkmaTHQHzXljfOW2sBBKhBAuilSFUSahJ8krHSbPf6y/KKbr2
7oFcsNuC3mLAYuCPOzXyG4VMbLU5CCeScDfbKR6I/mgP3LEX3UeoFeVfHWgikJuI
mGHx4ryk4T4XSLgIErKlbgxg5+4dUcbszC6/z0jfZ4z7taM3IFZ9agqna3fuuNCT
b4Hnd0coVybB/eXVr4AxSCm8ozPcXiI0qAKnkGzBPhzkxtvbtriNbd+h01D1iO6i
9/IWA7W7zzd79GGn9R+mLLSxalHAQ3e/+PDxsyml60U8Z2H8haBgKwNfKs4KRGlB
GqlOTsKmj4Fy2vSxVXwXESkIPsp6QUwqI08PD+BoAvENu4IWlVFzkwMJQBpgW75a
EGAseFELL6VYiHdHT6XRqVh7DH62OnlsHFNkhFG+R6AWCIPo/mDdFFIwToLizmIC
4+2AhhXLteJNqLz4Cuf2p2unBMYhqbE06Vlvf9ibZYn9TS9+yRzd2kWlWG07g/j4
+nsjWVQecvMfu8QirBeK7u1QJZdze54kWBFPoZDv8BZR7cVBdzcNBBMW3DCLVpdI
YO7m8Lr/31vC1F9b9nc3lz22i8TSCjVwHTNTjYoUGazsKX0Z/XFsr5gdkl+J9amI
ywn44BndezgBZeDMhaEHYWchToJf2CHxqcjP2sa4eUqBu2p5BNxuxBo1fUPIGDwt
1Vg0wEpOWgRQQzibR4ryOyZsXuaI7QqFqw4JdBrw7s3aEw1fEXUSnQsYqzruSMW+
A1rHeFo6xkH7XhnI7tShMaNN7k0NYYZtLJTQAZRS/sj6CK0ngVGV3c+Zs7xDHNLe
TBUhDGt6tyxp1gHJ26VtHw4rI0ErKfZUDu2JcNuUq6fOkZJEinujiQH53Y76jxQD
IMuaDXg+78qUO6BTVtECH7T/1itcRDk9OS9srj8hJvxq/xFWqfRP3iVmhdxknDE1
kdF5Sq+jYuHSj2RrfkGSHsiDr8RYYs5UmzYkPf96bUijRZoi9NV1xY3sCImVUP6y
MRQHpZQJJUxEdEJnwAd1FCBozQtoLFhIXWfivQIn4L2k6f336muiJLC55MXg6ciN
zYvuzFzNHR5w7VujcYK+TJYwsFVyWQVkxSQLsEJ56WxeU+F0nu7vFHOLjGhQrFQM
O53aJh5r3fGIcCUCOvk1Il3zuNlTgM9aFo1SCiy7MhJ7YxHzkIopLNNCLHl91zSv
o4yba1MfcqMuiIDaRa/7htK4f2UI2yVJXkKTmrGJZ8jW4Rjl+qiWz7E9tlxMpvaa
s1MUGcp+TJQ2vsYnkD+72vgdOF8z28haBXcUaHHseE+1jopWrGwLQ3PqEG/Z3T7Y
lUcEnH/EzkKpVbwx2631WcUpec+kJ8LhuFqQGrW+iyPGXXFE/eb5Je2O08ywe44j
+WTqY+ZIx+5JqY+dX9vWjMJu1icETYXxwejArGrYLKU=
`protect END_PROTECTED
