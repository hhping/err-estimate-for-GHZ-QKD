`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ErPKFcKNmOqT7YUzKAKsjWPwAYFk7NOkNwIjr/5a/w/u4nJ/375i7mbc81wYgYdi
n3fJ5YddnFmjX0GYjynh8VyS3SEu3XMhhxg09Tv5+Aw8ptSRpG6U9kQx3DtQWocG
YtWcmdTjINGb4BjSV3SaRO/nkBb71ocLYlPvN9Tdx/mC7gD6Sg1VfP5Elv0S2WaB
Wf+zSzYoHEuix/RAprTZsauXrlrEpn8mcp6eVnQ7E0mnJ9VKjSjnWEw+sT0IPpgO
IYLT53qrNBi2ZlKF5fmWdQ9RpReCA5M4Fsp31Z+tLEXuMcPbEmFWz0BnQdS9eqhk
Iueqin8DNSOtOj1qTybjvll44OMHJy5hK696zcNvnDe7eB+Ha8fqqvMH+/I3vuvl
E9iqa/JSAexEl0ffHMoF+m2//xjmk6Tq6IeLYoLvIx3T12NN+JKeWg5vH5h2BkBX
csGQeh5DRVy2vgnOKRG0rqyrFhn2QAyBr3SaUBwd2vneKhJWOD5TV2P4Fa8s0g5A
9PWh3akJPQsvsbfoQJ8VZAalWVUTrhwfec7QmmsTrerz1rcnTqrhozD2uqU+HnfK
0imMYXh+saZC3rdtc5XpA6QuZhKYZFdVyECtSm587lpE2NSrt4B3YFqWgEilML90
tfK0hKOcwDe/HVLEu1bfaSW5ksftMNIJKAVXt3bJ6HyJnJKKJEiGcBCGTCAcQM6j
FxUPkb5EKVRODf/9Fcen47IcB2fbKOnOa7BWoNsg6ao3tqNESeLr3Z504ZDqIuWZ
M151WWLfpqeJrLCn/EPuMlLN+pz70MGkA5rbKMke7z9mf0l6mb8iCAyB4qmGToeg
iGqNrmRLEADYBaretoPtFQ6pUq7YsC8Q0zP75gOl+1VhyoDa36an1/RK2TGxSor4
PFE/ejO5wAbp01h1WKTqgCpr232fddnc3KrrFPWFaHVgSX/EewKGjqMinEIeMRXe
YevaWt2KDSaAEKG0YMZo12+LEE16wQTpUNJq2Ghh344wDL68SyFdaLFCLY7v5K5f
qtVVIgAFBAXYRX2luhrz62TI4cwu7nDuPSyvGBObZqb+UBT5tTynFEwqetuDM+Ff
Gz+TaIKZqJuMm5aBy0dgOs76kuP9YctZWdzhMLtGKE5nH1nIn/0StmAATzaB0R7b
paobJH7XFKc+grNwARKKWbQR6bZKdb6+MzPwDtzLzhJaY9fbNxK3USnXzSZQTGde
HXTc1uxK6DplcfnxzXbvT+UyspTI8mhzg5GOSTZsoQ7009BEZ1QUorEV0BXwMRdM
JZJlSe9Dbo8+LLsX3zUpg60x7njintCK1frtG0G4Ipbot/X3v0SDb+HCmV7LqwlD
2kpeDc1zYlMQNqnFJ+GP7H+DjdORafGwcnEdQ5P+iBUsgbu3QkNZGjzibFn6nf3z
5O7Sub1DfY82aBJ9z2LWmsU9mXu7QBFnywPFWuSYU3WkOAWnMgBkD9mHHwaOy2/T
ahZOS4RonHq98JeVvfVQ0zMXYHJhLFrs4+4VUJwzHE+t/2yCVWmiIgkM0N+dOYB/
sB5vJ+UuwPNT+0lJk28CIr3QPRDMBOf4835oEdGb+kaE8+Q+5fRak16bmQQJ0QJn
x2q+d06K0K8vjmjcw2DvzIWF/bnMSK+zjHnIlYUWoUkhVlDhUP2EWc4Yq+XVDBDD
GPntoeuDzxeDSbnQGd2lJ+fq2m/3B0aN7TVxQpZoFlCmOn09F9etj3Q3sLJ2jHdN
oVNPJnWczY9j/RNLiXptCixXMjUseP00w5RpJxwAkJdf+vvxZIs/5/C+Tcd2BwUN
09OhPmwN7q9Dnsq8qaoX20+SDDS33mx3qOe+WhyC9br2AGSm/mvqsOVMqrYT+Y10
bOKThoYoKkmRDkumX3drJNc+EmvorMtZZ2UQ+F9coLQCY2DVxSWsJ+FfLSSbrK98
kIiqoUmPB8dxjzJr+9KeWwUv7AA9jaaJJQsbR4JoZ21PBRda+yiWD0lQZNy91O5F
iTeZN8pJMlYSbhWvuEV/mneUSUDlT6ZrVoo0gmuhq4nIR7XOqcsGw+P6HBTj9mj1
HF8R4LGeL1WYMNkka1ziln6JG0tEOKeII0PvZaklBFdBhvM5CEdOZahSGcl519ry
DxH9+HsC8vQ+y6zVqT4ixa12XTxy9SyBUOPOo3Vc5T19NEFfPt23IYR1FVzyXWvI
To7TiO6t9T5ONZakNgqmdPCBi1CIkvMLvsF5mkfuIfrLVIUgrxWNX4wn72qQ7wcp
+wSPENQt1q1wrrLnJzTJfUJKBRlG9LSUz7jh5bRrlyEvW3sQBJAQif/ZYxEGKuKO
Mqcu5rwM23lThmWTT0roIn7j3gSCvPfApfipFebO31123MjMepCdYc/J7HUyheL3
NzTvxkTGAgJxEyxP6qRhF00Qovk33Z7ygCxRMo9s2Ew00JyOr5/noYbQn/JSsYy7
vuXVjAmB9UODu4VKbsez/jQERc6KkVbTV3bO6sCD4AiV6iE/1CQnRz+qQSLuO2jD
sauWrZObF14yNzGohkv/wPyulzgzHMvr1r6ed79JCscrNzHTuwOJr3XjG8O1mI/n
gbrgnPrpq7JzB+nibtrJgFoSyBJ4HuyFVpdle79niCxtXYe4HgpY9cxkUul2ZVdZ
s6xQHB2yeqVTvBVHx4rLFM82p+UMU4XyunOx+SUtB7QRHW2gqKoIZTVMqLz/jRbS
MBTr14naejEXIP2YgwxgtJscBjAQNA+nGaR6P1mWyPxyYAZ1WxIysltRbyOyZevt
NkBzaE0MY3j+Z1RRoONLrTppKF4phvteuZGWlt2DAfK85u82BMIof/z1EjjKq+rK
ve1ZfRGlPwHf1X+dfw75GKogciv6dzHTzX23486qEF7xoRsKvXL9bTkZSiWbUWrW
xKaCMtijDkzUQAHLKwYo05kwNpInFXhZ8jYLG2XBchaQ9g5s95hVUuPoiR9duiox
PoGWsRiAAhnX2dRc4qLITn8JaSAawT3ahrc38W3xloKEILUc7DIlgcUrf336IobH
VpK6inuPoSuX1QU0xzwCcxHp+qKAX7oNpHm2IYwAyDJNSr6VU2eLRo6jUyRkeeIB
3xJNSgErS07JnZh+qPayfbAed+2amiymanPpNK1qT5QLUaHae1LgCoqXcvLZDQQD
Y0SR9ctd9jztJYp4dt7aGWpBRkDGsaatYRpCxV6du1RFjbu/t1zC1GJwGatIH1oS
YOamaWdw1u0pxm9RgiaR6slW/zFYYR/ay8ZMSPbmkNPvC0ERkxLGSf/ZOiWK34OC
vLZyRRwTbyUw5LDN7qYEv9M4Nr0XX/as+MJ/rhhzRhlI+P4v66Py/kcjciEKLA+J
YWlBgnBFNjT6r9ERgkdowcObVBgS2HNgGY9aJGScjJSgnyDduKoH8xA+k2xBeVue
2Y8o1j2FK77O8TeOAk3c41q3kwJnBfcsgfUw7CyAVphCAfb6Nu/R9UjJMvNNRq2g
wm296pmxuxMykJIr4ulToj3Vma8nq2Mo6KACGiN22EUpWlVJ9Gbe8ZeUKDSPE09+
rF7c4d6dYD51qgkINj8Wrusjs9Xd5+geJY1CAIkgq+JNPkAutkSzqbnS3OzrWABE
GHX2xIJCHYBCjQfPzzZq2C496all/aJboSP/1FOaHewHCaQpYi/d2hAP+af3gJJF
RsS45O9lmZjX1Qh1eApI4iJMYgXG9UsHMUvAn+dZ2XULwBEieZgvZbYQswrAQXxo
9NxCXmhfmNSM1wsOPny60IgJOfwvR29CnO/KmUc01OEczWrZRlUNmUPQ/DZ7cdIM
U09Qdq7sazxzZxVWnycUPzm8HnWAM/ZfqE1wNeqbXv6SLM//FyK6UyDwn0FrW4mj
ZskjPSTWk2Ur8KufYA7Q7rdhGrIGXeDNSg93uvAsLv8Hsj9FwLxRB0AGg6skwa1m
Hw2Y3VHMkBJbRXtUquaNVFCkR1lMf474GikcibER+WHJKh7HQ+Iv+jym+p2ogsDj
bCxBHDmp4k36dPHLNo/o1DY7pyAzWl5U+aFbg7L699jMCyuFybJAJxJCHUYBtTol
vGEvFSgMh8Dn2FkmhlG8GK8B6pdLrKguePPSN244DxGl+mQYdkvwHicK33GHVdfa
HCjZG6RMpC/seYzKmQ62CPhI+XunQV9VlBt5+v1YJY1I8yDOspDjHU2ktt3qS+Jy
nZ5t2fBxUO+rrCudatlvTlm2Wi8GysQwNX4NaKPc8tYWfrGocuK7DiXgfVLOCzxT
sc+pK9a4WZElbZjJ+gK797dKwrQZI9sYxxbgVSRlsntYHgbzzCMptqHCCm5T6Jt1
DXizrsOY0pPFOArFfUBA8liROCkWwHE4c9t8m+9gNK5KZ3QzMlZWTi2iSAMEKc66
Haj/qmBw9xfEqQHccPIWFrjxEhgz+kONpPcDHFgbrDUmITEUsFVEECRmiyXuRPip
T7WrBMMXAbLznNsEt6UFX3W7iEM3HmYwfvrBqiLyPXuugRrLgkjQIYoLDOMWcL55
9rf7fJ8y/CriMek/5jztqKGnUwCy2Mu0q+20Dr5vaQK2WadCmW3zYTRrpXL9XpcF
JtVQ8Ynzh4kBpqCR2HeXRgpshXa+BMx3ExEsLfuc8b/cAgnnEfmG+0Q+gxzT6mQj
RyxQNjl1hv6ZWJxviAVghtcjoXDVMzJoNbRxahN58d7fu+6DR0Fh94gIfI7l3xWU
f/JRKbpKeV+Y8PM/+Dp4198T9dYUfFm35uxF0uWDo6wOHXgr2qfolDN9AIHHNv6r
qncqSOd0Iw8rVbd3fU8Dy77sXWpjD6i96r3YtKyoMI0KcVBLE90WWXMKMRolGNeX
rSAhkXVtCvpm9drSh9+xKtunqD1HwqE7nxlAFa5JqhdtZs2DNk7OMkLHoKbqWH3J
fEI1Xal+9JoFPUEDhCE7krOTD+PNnJtkFpDN8poOzY6xPZa4GNNndk72Etcty5LF
uVHyLOLonXr2flZrUjNkL9eaX5DneNK+BjQ5IJEAj6soUy35WaEQ9Z0662PndFRm
YvIq24WC0MzO7DR1gwTVOO5XMYDzJN7oGRP4OfxeUwcNHsxeWmHTwZRIjDMt4U4y
Md3rEyUd6VpTT+M7hsbIngoTPFGMqAanpXVPO9EjX7B5KB1dKtUCosTvUFPS8TWB
7qfXbdaXYdmMRYbEx4vZGGz4f9l3dQEcZTmeRAEdnIO6193Zy9eJmFFxbrUUG8JG
P1e2eUqgtEaxtTCMjQF2fL8sI+nVD4GHJzoyUEPF0lTj1LGqi0rcY/5qxwVV8yII
1kThdUZ+8h9UICUasGz6JZPIWMxUenmzhFojgIYro0ucPZe2f6sPPfzJaGhYeQAs
MkLb+JXF0lvtc8IFuLeeRVrpiia5dncgBA/AZJBRa6J7dyys9zIpycXETCGxr8w1
dMNZchJCu2Pv0cQOwmZZQblwG435k8QovYGwuhhJVqHRu2OqPT1MiYz9Dk55A2qT
7z+BQLTN/Vx5k/IJwgOODspb7rFRg+8AKRx1/8Y7k3EAcKgA+BpekjO/U3Z9mi36
AVjOqEkN8H7kDWSbIqM1UK1/LaYaTcZYD+H8P+f5ji8Xbfy7PdCe1F1NV0gl8kKd
mL/KtOqDiV6gVklPqT9GdrXsNyZs+1pZT1GEkigz5/U+2Ab/ETdC3EQzhJ1f5WFS
Mcm8syAzo9zoDFTH1xlhQFcB2I3d522ZJI+ovKmF9mQf5lODusDb8y+Jwqu6OzdC
GE9ah7sEfmoXfkckSx/4Hqx9WYoglMytiu3i4maUSnhULFBYDGTFXdWrxkSB16G6
ECl+6HFYw/My8Dmq2U1Z4jMDmNr3JQ+onGotiTVqiLEc3eO/e5Z9Ie3nWkxBfh7G
+TqbS1OPV2jcvw+CU7L3eqRJ6QJWyvlgamqHFfIUgMiBExPnst+wKibMb836nr6R
qRuSm7+wUvKYXnGf3lVqSKztu/3Fjvcx8jAelFBqT5JZMiLD8YtJUtp2dj10Pe77
DCfcwgOUb/2noxkzdwu4j0DH4ctDdkjijmMMBD60sgCDqtFmKd+MP7cUyKRI27Ce
cT8Xzm4UOhOdrGSwdS+XdyCbmd/IYiIkaRtoN2iEPbxZd/SarH+m1axQTYyOvmhl
5InlBcnpaUIJFIkFIdzje0w9C78PNgBmSACKHBWbf6QEA7ITkiJ1IIaY3LlUs0IZ
9H2y98B3azOslRM8R8nPwBaK48l27V/Lyp5Xv1QUpvS8ouzJSdDhVRM7EfR2gVn4
Bz0iexyLM08CZpiSkjmwyrjJTJTQ+3oCca6YvrOg5g0eBaGdup3m+nI5V6ICXWMs
IMKf4wX4V5VqHk3AMpdpdefFlfVG5cgWLqpn2/l04amaGRJqM74pTP4QY2yjucZP
jKlsiKagcnCSU6iIJQM2uPgKQEMvjywGPoiVHx6JoCEYshZJBORjcxxTf57xfFis
hudV+PW4bhurguagflMknaGKoYKMTfLgM8CshxCy/LEWGJ4ki8gCSPTKY8GNTkGa
nHyOkvGGGzRoZZJEZBqELrmhYKEgv3OnwZK79lumhoC7kkoyZCJ/IPpEzKXQIG3J
Db9dBlKRPUWzkmGMEnz2Pg0ttrndr9tSQ7BNEXZJUfH2nyvtmu/Vj62Eq12W2H/9
tiSfGX0qgSODBL50xP5K0hP8QRabKnjTlJIhi6F8xjfGVQxLAHVL2ts0OADd7kYA
ny7FAHWM1J/JssIgOC7jvY/yExbZM3wrNKAI77V6fcdYDkX4DQ3Utf/QCdALJOQ3
LEfSWS/7e2QvwY+TqBrrD2eGpn23lBiyTQpc9D3tlZeSIp3H3HVeJJjneXNJZBZa
6P9DhpPe0SrRJp6VC1VNG9BPtDHIJTvp7KHLj7X/h1ZRTHmWQKfoaDfmuGjmHYtM
lq0nMIkp6sMhnegSLhpCuf+nAl2v8TcMdruxh37KP1j++sRGq7M9hbjQAZFKp48y
RhsjVKpaf8vzHm9POs1AN2zFpVDFxk3FnVJAnilfKbDSnGiueLtWdgz+Z599+uk/
D46UhmLZiyBXvLR59r5puz9TGrwGJrgq0GMnQLKnRCYEt60PiCqUTLdIJzYMsBzo
ZHuAr4UTG6k2ErRjFgtb46vq1Xki4HyyDbOIjHANP2LCnzN0KWQsvCblPSShnV1/
sTzSl4jhHETZD2CG7gKAuB1p+78thBJ3UbtV13674RZklEo37Rk+drERFni/PqWX
zyjWhQRK3X3xbe6CulNoRhdZdgLl7lyPC9ff4zC6WjvHF53hSMO6z3arNgRSww29
SSJKjlv3KiFLvd1c7Ojne6tLlgD3d2ye+BsHidfM0uR4Gdn6u8yzAX4KFq7/glzf
wUz2sqv49tykCw8wg+Cyz5uHYnFkjkvLkcmsuSms0pvLoQS4M453OUcJTq0GwrVS
CliLFkqtuoesLWx0VS3j4ko4PYn0gHC9T3aC7RyTdAAniOkVsEYxGujbBNZrleMA
C99SmIyWZVGFHq8pmJn2hEvyt/QWnJJ2c3HHbi0eIYWtJFvuATdwEcZzn7dNKj4N
tbk/BaTh3qyvtefE01CgdPsMSeXC6bsrPIihDM8MuG1eeqg55GQeinvCU3csdWQC
0U8AgxroicZRpg4wkJeUyVmo9I//wqxS5hZxOhRXlnJz55Xk5prmiOEwP8mMjVmC
ZuGWDiyPRtS4hf4WibF1ZgF7UFFm1FnAECFwbh242V9Aj3tq0foo/CRaO9dpo2dR
1jMs/0ftPBBWnmGbe4+puTA6Gc+Lb9Xeadcmd+5OfBI5EOd/hIrQZhl2WeieQsaC
r6xYCb4vDjoROopz2pPGSC1ekh9ErhZzbEKblkwMVtrW6FmJqkikhsJBKSRlmyzX
2iTesf3ilzsXyodHuVnSbRJf84f5Mxus9RMmmgV3dynnepjsKpDHFIxioQyEpQFD
8LtFsjZiGvTXmK6iesye6P07XI7BzzP6+txaha6NUP6F58HFxg1ztXhggqo7KAuW
RKboipu31M3IsXY0VNb1QnOCRPrGfYpeE0NZq/FspzS4YL/JB+AI/d27ydLspbab
exMkNc3KfAi8ast31V5cnE4z7mma2VluAacyQLG3kY1E062VnEQrc2lw1gi5xS2N
LzZPalpE8QfG70vZUhUr51hfoasVygyghUhFDOe4rQufeY+JNnwadlcr8l8TyiaO
hY9eN64buraRySctXp5mygmJjjo2BcgXxQaGP/fPXwf8q1cQO+2nJy1juJOmocGL
NQYLtPctzHYmDF7wRvu2Jt5Pha5RTJkAzS/gEgfIO6raN9TLqebpmiV2avpov/DT
0LF5Iaq/dPr6Zm1QSNm/wkeDOQUUy5aI7SBfCXL6tLelQ9JL7KKLlhcRYoNOQT72
pIgrV0CrjMzAZFFKgZIHrlNW+uVHz9GoT/Ngc60VSNifWVGyUIfJpgAEnivotc3s
Iq5IG+Cfa32WnWnT6fR6mu1kz++VclR1r6JzIUM+sMRoZAfPOiHxkNJGqCLfgN5V
E3M7KoWxfkYoyUCHCwHFc9bIgBb5G1n5I/ys/ObnJd9nLrZcwynU6K9vjUmCkyvC
SuVw8zSaKeYUT4s7oVDilPRexqKTDlT56D3B3jB8Om64bCSdZgbvRPFKHsDTpaxD
v8Ox3xnDJtDsl07Rz4HVGFPQe/1qA/YcdkS5iFw3XzNnJrUjP/gYTyMD2YBNwcbs
DH0YFFXdVglC9oI300Wqvo3FFCKjjO8pKu66ZriKI10NP6Um523xQie/oQMojCxR
AMHxOuYP/UvbBhhHchoNbyxwLeK48KX2TAsIpxj8sVkzXQnOyp5djBNxQDglHgbR
yNI/sdKpAPF8vE2FqN00Ifyfpc0IbgIT2+ofC9Mscqnck36S0iQfCXji2KXU/NqR
jyGZrNh22r532DqSX3yTa63ER1SlDVvdlZPiIOXAAx186q510my11le/Mt4EqrdL
Ef4DXGFxVg62HXfq8dR9HsQulk5D3ilztnbFpw+oY4trxE6dFkGCYqA44sEBe7MQ
zOAsYJC3hsRvl+IUvrb4xCeHW2h7nuoGt/Z8Ov1ikZrk+EI1bXhDk76euSZkaTzW
Ulu0LvARzjCztfWmsv1YzF6TBvONfr4vsw+sAo47sfV3XyFoupD90vNAZNugMk1/
1HVOYlyJHW4R/LWjP/jyv+8fnkgFhMKsAClbR+dvmvRlvz4P6FFRnZH3ihbAL1CR
9baEDdP2QJ/eiif6e08sUkhzVtWqwDe/EhO+n7+H4Z9C/xgGXh8OngEYLNKhqqIB
w3EUHwxeg5sAoe5Sv4yFegtkGK2mwnjZ7at4QQN5cYooXmILenclCvttQowR6OZG
20JWwL3moW8AjgalcVsdkCK6iHS733OQYySHkrhdlN3MvOtJNOOuATwRyuUIUrmE
ii3JCV2OssefErLAtXCY0qdWKoj+DpagLfVWez14y73Gmzjf3ODppXD05hglelyT
/WTcG4jA3aepR8hs4m/vvqrLPf/RpKCpLbLQTe8K5tfmWBm7QCDsqUeSHIYBo1Jm
VbVrpbmv9MU+mxu+oDmZJKjZS7mGrfQj9QOAIWHqEdvhc2/Q4Flor17oJwHaWEFx
0Ii3q+cFhX2KStqkZYO1XLT+ORVgIDNTZCl0aTT7y4tuww7sgO4ViUdMyBFaYWYH
p865NSkAHFJgY2KJNcsmWzidvuJiHoWR8hMiXZ37YA0xLi+8IAp7rWdOb+KYhd7y
dt5/sXUElg74YPMlelQEzuNc431yEDVE0ua6vdkh1ZxpgrJqO1gcv8NGprGYA2rs
mdaVJcxd3G3KT+UAgaUsd1ZUeLJ6jDV8ZRyGikqQCvbcbGWF1m9WWHIerJHlCbbn
nxa8hQUZ4hIHKypwxkgPzKuAhRccCZarWj/M3yFgz0vk8RGmeZEJ7KU63ZFsdi6J
kxq7f1A96cJpVGPDaDVUixSi9eaGBybreZcfGhadvrhGV/Vu4qSbPbWBZs54cqy9
Uig8nripCst3rSCD2uszdtZHy3ak+vs1DJNJIN6dh0fbsr0Qvx92nQisLf7sxehj
9pPZY0Samtr8a3EAfteWy3DWVfcRQvOHChZHPGkqZCOhKZiTrW6/80Mbns4y6xg8
O5yRVDrpw/eIlGl2mcVIqP6h5PbDEVeXNPhyjkK1YcP7S+3RYtjKr/0K1aoko5Ui
Rujit6Xos2U6J1zxWQDShiNgvQPxOtaK5YTspw8cZ6nJjjsAHnZPB9thrcSGsYjH
lj++eX3sD+JTCrIETmpWK9sNqiLbfKn5C3u9x0d6d3K0gXXt5UlB6dYZU/tAlPE6
6potbacrA7NQizviakNKe1WEYGMOBPKhPUlFBuspwrE4HuPNLTjOFH6mC7uzrdZl
I6QIyKxuLjSof/U945ICSJbmP6I5O4/KjnbjMNJWyaIT2xgv7HDQZDaLjsni4B4G
+S+G0kFWA6Sct8qwcKLpqqY4I0fmPykRlabrnefLYfU6gc8oUaspFtXbr0xHtkzB
+KGc4V9wDkA+6idYvxyZlM6prvQ2UmLxI7T+2A1J0kCgsOyyUnaxnWvRf/0bS9yF
cjvxNYWe7XQnGLY4W7GNYlOlMxHmR9ST0pTXrCSDaf41S66y5eci+YST3RmwP5B6
QzzlQJXQj5VbsM+ObxQfA8KvzYgwp66wXncPwHUQY2//CIOZQdfhIuCIsOfKW6/D
0k8/hm7gYskQTF82AN8Uqoqg5AHAL/ARaACCmHBCG1LZPtgLENiIE3jztPtHoXfU
CPEb8jNz5b/S/W3bF6eb1GItssqU+wCMAciN3mWUbZaTJadej/QBBERlWfUag9/H
eKXx4zZZwIj0NVItE7Lvv7aDBafpvbwizpOOBJz70QOJD63zFYAqCMhl2hzKU/Xv
HRIbRlM9Lfoq85UzciIyG3UHegMEMwRLjxBOeDqWyZDOls5dpNnrsINOnGrUi/NL
kPAAIFIbUT8x+xxuUsa+I7pHomQjcCJ9NXXQTEsu+bq6mrpvKMogwwpyj0J7jj4R
UsEfYq6+cnYYpWwKLGMD0gZ54BbW0qzkb56Fj6FHKUg3Za2b2GVtTw+/9PaZryyt
B8J1fpiK58X9eG+QOXrobIwLyeIU9Nc6TqjTsUsf1JFoyhr2OnEJav8qEk5s5zaI
X/Dgk26kS1gArbEXwj6TelNv/IfxNvi3CSf31tJTEWxRZ4FT0VAWEkMHQ+hTHyZR
FZZ2LkondMAfxBr3B2tWweFz6k89uAHhLuE2Yrkgh2MtwY4ogfOO2I7WQIbkOWOj
9IiaeqcWx4EF295E99mCunuKgse7AiKQ1SHrp2NyVMpAYmbALmMH2+D/61kaVBwC
ElhE1wFw12J4+MU+LpVAEkkcP3AAT1UWwVU23Z44m78noaq6kly+GQ4wHYWs+3wp
0yVJDsChPgvNW/eDc6mrn4RYsTyyDW7A9zeEJ/izRhU9o8xjE4L1SsUh9JPCRg8A
scnzWTCoLm6mDUXFs1wmiXTG8RxShv8IasDDoE9Is24DTpfghUsONyG1GuqypunD
r2tzrgBaroo3a4RA3XLvL6xtGShM39qfreeqllR3d7/ensx9QeBhUY5xJP2DLBHK
8ZO9E8WraYIeZn/p3Nq/KNS80lCC8qJ59K687gQQS2Y6JfQGWjgAbzaBxvfNwPdq
mjnkx4K6XvFPnKW2BavhihShaOX7sbaldIZ+oLlnL1t4Ejjoq7wArzkxhcdjb6oX
wB4QbbXAOA+feuIYZQVUQRgcKn3wzVVBG0fWVlQGUADYR8ARyVthn5bvCy51wspz
d7TnvmsFJQ6gkB1mdlRqIHILluh18LIRyJ26LKpgoOB6A4iXhuOdQkx65ptA3xVj
xfmGr7oNLTJf3t9CX4M56CMdwbuD7jBbGQN0HbBYdw2Lu4mN/kbVLepRXoCO0XnH
pLOJAOuLrabeOWKc/zzB+4H8zt1p/G3rh8B0kpSLJxvQ2XFj5p2tB1HqAsPWxDi5
2g7+VOSAypF0OAl2u7CZApzT5smn+xLg6C4aA1OAEwZm8RmMyYsxXNiTIvtTkPKJ
Gkk0lpUFsJCAyDnsdfj00LGe08O3Rzk0xtzalRLhd6iPFqFrav7RDI4r9kC39yY/
T+XqX9/hl7X6aCID8OSae37miCvWMi2Oy2cRMfhBcF7quVm9sx5lyVTDMT05DzEZ
/IULLuYyKNPyw7+GZIFPo5aQRAwWewdyLgcoervS39b65zYZthZT2SDLxT3iG1l8
iqHMHYLySVFTEMHAC05BjhQyAlKL1VQocu5Kpx5rg7dcVG/TdLp/me4a1YnPNH9Q
611eT3SFgroEg/HnURRs6BT68v6mx0JevSv0iiOpPbyKO3NEUgaOcFduda13tfqu
OeifpL/8B7IEoy8chNzLkLLzBg0IdnAj/2dyJAak33FX7JQSZS3EkZWzg9fvhgcV
LYFRhYhPTMAa20favbHivRnTIYmb8ZPpE6lnN1uE/t0zd12dvzw+e0leV11kYnNs
xw109SZjgKtq7f4R2mHCsn6Kf3+nzh0Cr9EyjYAHC6MEhFbOKkNf6P5mHhqJAo+w
fU94dZ5vnu3Y7z/+PUNjdg20QyUBdyk1lEpBgfy/vvXLwArctDeThDRitKIFWVU/
GKYPpnsvBiBZHy9f/xB2GURPWxU2MffqcpMfWgzjAH2QJnG7vp8lPh72HJizeBMG
TzN6/uLnVvAhW/KYSDVRgKot1zk1uB4A3wTYBWx8yZL3/6f8AwgoRnz/hM65BYNX
GmGrs+O7h71VbiuM+Zh6KVk+jfBD9EqBUYDcKswncie5ly0n1B0wi68KvQT4aWDt
81HKr2qWwAdReNKkGxrM6UeEz4U4atVxugaAZ9tvK4vSjCOxGH4az4D7ZdhPZnOG
lcIXOqe+Im5rvzNxxgm3PdsogYZDiJ/sHTi6tUqXU4TalHgPpkfOKIQBZjJ8mhUN
yp3dwjuxEqy5sL/O3FTIMp/9LwUrSjblh6F0XL2SDY4GHd1o6olpvl0XMBa80LsT
e4FoVrc+PQA2bqPaGPRrThpWmcetEEKCk7dXliHIa/Eekpj/IMA5Nf9j/fvW0ZB2
NN+OpdnSf3CJSB7X1J3wZtN6Ib51P29D4Gyw3v2G9XIdCecCE9rX3p6r15OzHb7z
rdeMW461nNNr3X7e1BmO0PSKRP7cuppiDc7x8qAgGBYy4DsmX9Y7rL0G6OiSCMbC
ujLkY+56fokejDSX0YOOue1VZWlAaurkwE9cSnDT2dpsilnVo5WrbGASO3DkKOxt
5h+rqckAXzfu4ORT5g2jd1vcTkIL7AMe301PtX4A5E1HLSCYfNI+X+0m87/qlkqQ
SRDPtQ+V4EnclhIaz1ppSVnmG6ZUWW32tKlBb8w+4PWfzAghpDftbcLYvaEHBVhb
eF6s/05BM2Aa0SYWaaGQZ3L8l4wcFzTiJKxJfgvn/E+UQrNj12lu8TpwrOzxl5Wa
c8iNdkpIGy2vFEIH18qczDxq09QTa78jHpYzLtbI+pC83NiJJ31WrfuneENDb0XQ
xjUPgO9bwt6bdr2ibgPWAqGOqn/3tlekeun9gnpGKdxA1eFRudo23K4jZPyYUSdz
hW4bBA9zWDgF7E5ooal1sBD3UpBsvkDadp3fzmuILb671m+hRTgwevULd7VzPlnX
nE1K+FVP53Yx4d00wb8ylZQZY3RfmL0XAipfX9zl5/wf1IFRRXweqoIRp7t9AK0F
V8PZMfVVdyePYtYKw8kw+vZT5gqB6zGL/fnD/XRQDJIb2X9xJ1ne5GYtr33JRACj
x/heWPLBWL17wlUH8k6WUoofWz74pcHycrZ8CCVsFb7Xoiw31Wtlp9l9AYpkt01C
EhKi5YlMecQ/zno80dKSTDBySrjbifQXGImFVbs0ggr7AuyqqknEnnClQJMoya4V
OvlX5dJmM+HvmjLq/RH5DEscfOVBkpjIhZ3q4NkiE6R2f+cN0go7hWE7vsOWt6DZ
pUCMxgI5HhZUMgxGMi/qAvgxI8kxwXJQTAB/Jtz/aPLpOWLGL0E1hQ2Nzrk64qpR
Y+9HFt/Paz8wbmqFiRLt4KmnLNmNAPW9DlsmkH7PMsxVMIt/rr7Tj69IPlR9AUgq
oa4RiDTBSBttt/ToBQ6UHIjmYtbNgxJ9Khh+NvCIUJ1FepH72439pDPtWGI0n1LX
ZXDLsvLjioZ1NzUGw5+MRK3dLbsJTgpV63KWNmt6x2MqpW4Xg+4pz92y3mM8+Bhu
MbRUhUd/2maRFaad9D1IZ6JEIg+vFl7JdNN2MUyQyAv4qZrUA2AXZsvV8h1Zfkt+
e9rruosCDj8wfad8s4uTlhbX4QwU3rjuYOWrPVChOq3t1J50NNlY5Of1b3E4g+Qw
rHVpe9Yb4/9nFbZfBYbbmg8MBK5+9TEPtKKUxEcAluHTAE4h1cxhqBsT8vbphy9W
HL2TD0QrGac9DPzRRoPrZ/hSy0HHdaFdhAboGU/me/gbxxKU7Xa6KUw6kUTz7081
xIEP8LGaIIWTS4zjm1DF9EOwKwPhJEItHzSG4eMd1iCpsM6MCXEO0o/vH0M3Cq/t
yPv8A9a3A8isD1QuD8Im3TrPt1qmll8SXSQAwox3cN4FEWSTRszDfdnHScxduAc3
ODvhjUcJZ7ZNbgDWSNL/VJnQwhWmurv7UdI9E97HOzIPTaPVKUTFTYBBkZH4VcM3
E3tuKb1y1ozoiUvGSuVq8LJg+Miamo8uMuKmGpuxMexpWFjd1N4pKqYk9MhKADzd
lQXxzzr2j5BZXrAJac6ntvyGHTxgE5dUPp0h6N1ZINpjC1/2A+jM5GzkuWOgCjl3
nIdU+otBLexyrJmxQXXdcFc/HwehL3E79tC+8wGV+lTL4vMjKJ9GQ0CeDEp1D6Sg
yrPGYJkTrqa/nOHFwB92lkeYguliJD16/AXVIunU3jWhd4wuymC0+3jqJF46EtHR
EMttJBlsTl5L9w5nH4UyvsR/bEd8qkKLiAmt+QzxcZJo5AQXGhw+BzA16GbfEXmm
DE+B1dz0nF/QiKRpAzUOZ8goMcikl+4SxoLag9r/GUw24xjbxBHvEPN3dAqsbmHC
oz16mjKR9vLR5/8qb9c5fj+/wm8u+yjbdQgdY8JHKuft3u7EoLZ03KDWpMcs+VCv
My69lUSkE75e2l77Y2m8izHdqOq1Ct3UorFO/+DbSf9XyZHN4ytIXEKO2PzT7dx3
wwegukhnoYkoi/RC9ob+raZi9xCK8R0IhQ6JMXOzaQOCsZOOsTWYY3FvXyaVp+1z
Xs4d0RL4+UnsRbYzLTAttWI/h9GeXKGvDR0NL9IF9GwSILlcLKyY4ShueRoXCo1C
Dq+/EHvGXbtCN61wHk07CScLnL7QRZeq2Beshb9EwuK9+5ztREkQLCGbTL5q8Owe
A4/yCmhafUU2OK+KEd9FSdZja9e39lIrl1GqvCo4MrHc7FA2dDY3u6Ol9Oc6yckO
Y4lLpRatKB7RyG8hfxqfntJRnlRE7VNN0wDZShs+RVyDxiT+CODR4dBhRpEFBR5E
y2EWyh+8MbhRpH23hB1jvJgi2+39lgoxIglLjPKdYk5X3qhjTxM9TVSJcEGzcVQC
mBiDhHi9KV+hQdaqF4FIYIjk7U/HJ4Jl4wV4Ci+hd79xwynFycLfFrBbJSX1DTg2
3Ypqh+seXrkRjcNJB26vObImaEDphlBO/oPSBOU8DZZ24qrQ8ATJ8q4PgG8Cmofa
Dxsk7ARof+F/b+T780bhHhocwRlLsX2UWABFRa+FJZEcbga+Yt8RmagV1/V0PYKN
zn/K3VRdjChN6SDXgaTylPcBcxoruOEEy0P3a2eF2/FyladxQI0I5E5orZffY9sm
QQ+asDPGPucL42FryxIittFTcYD3gPPwLdX2rnpVLTgx5HJR4evr74hm5+jJETsi
+9D8yNJPSFt9oGNeWPeLnVxEtRiOB2fc/WKpBfmeYJY1toInvVGR44JR1HO2KDyw
EnTC3I98eeojXvKliPa+XCIg1gLC8aRP25fm0Ax6lHJhNRktNU2Gd/QiXMUr/A63
wC8EDvHPV9hzTgVJBEeoF85zlg+ZwywPeHIJWNPSacajTsREXbMYvwqDfCJEBHBR
I9/JnqwGY41pmRJlJcOsNlvTSmEN8mKHKG63S28aXemucv8alMEDvdNVz+yJ6O1s
soggOXsetIiMeVSpp9eLbyl79xugLrrvaCx7/nh7PGOOvXcUPJvkv9f9o+mdkxfY
PlZQcvUqkdPKX0rYA58bZbm6M1/YocfnUaXWehsBBKatiXoI9azoFa50RtCxA4M3
GVLv8ybQGgAQYYuJ/AWlSwXfvFb44QLs892J4tWbLnTgm9RPucQ5TnBC/gi270VW
ALPxpeA74DiSVPpLf1es/ryXYjZw39eibSGbucwklnKhYeyFyXd3R6l1CwUBX3vZ
BVqwqsYcDYvQFSyqjCMjVFMUOfSc76YKhfZuGMbwLDSR8Su6sYwr/gQpOOqMCoRI
yzzbouh+VZezGnhcJSNvGMerWEjNwAQrssk4BJ4M2U7GJ4TmBOnBm54KG/y5zWaL
YQE5CYQoAcxk+X/I4SO/3DtcrGIhI8L24e2v+1bReZdBeJyE25GduWupbc3jqaGp
noS7J868kbMslaTj0aADFzSv0l1A8WA7zQ+K86L2YyCNafBDOjJ5rNQ+WU1l1TxM
zEWjaOT091D/Xue3japTCiDNLTDUqbRT2j8OSOmMO3A/tsNkus3/pT9klDKIxaju
fkxJScF4I85gU4Z8BKkyPSh84QYJ/h5MeHtvp+FNNZBTu8eCoJ4xGQviAq2tnIX9
OQRS6q5yeETf7iJ+Yxd8zPByvWqdCYX0+Lk10Mbp1R29xYZMUsQxh6CXxM7ye70E
Qtyy7aQ//Sut5AAvVIq0KRFgGaLgbT2Uov4ajttTdk5vTQV4BsMg1xrU3eIjy8B7
9VghNHCNrFN9zBFG0xVpX+ddAZ1jy8ENbPFzGJcpZTsVrSaDij7UB5RV8l/7/jUp
guKZcCMAhsdwFZADffX9GHgYlRyB+Maa48LYLm4opnUeBwOVWfXfLf7PKXetnDzp
q2DkpqrvzB7FUi4Pcyj+3L55FBPZW3Hs1Vn2vXBplAykzIowBW6lr7+oL2uDJxis
CjnW/fCnILIJ5KIhjATDTBDg1IUL2QiNmIFFTVIzhDrJC/DFFCnjAA1o/mCW1Sf6
I2cpW5xK9hlWCABs6IuhUG3sdkLEtV0Gwf8eoA/kwpi+LDnelCCgSPVoqrO7wx86
2c7D4tLvbZ8dcsYzk5Wme8onDCDA0t2zz//DvDj3+riSzvy8B4ZlOXkxEXd7WhP9
wg/CyIl37VxRqXNGnNmSotVd6UN2J2Ky5hkSe0B8FLjOQ7WWD71HPR4p2MSLULZN
wFl5BLOF5PuSBCyZ1R0L5hsCexUmeoxgk8HciPhwzVm9EotQpe0O7BDm6/F8lj96
sVMcmxOt9NZ07EgeKaO8ssKn4vStXvx6r4TIX/ZGznTBxuO8PMh/eQy6STLVfYc6
uNwKAAh1KQ5ZAdjeh3gPqngB2HSIKJFHGrIJbgs9xy9WcjgsUZm4k6pPYPFbJtLY
lOZz9yoLYHN0Ztx0+gyqkHSTNBwUg5NhRLD30QfHXWF/BkOLx44v9gVwnF/O03I+
ozb6yqndz0f9sk9TW3kvVt+C0ZwHLiw5iAnnTkXgmKxNHtjddnWjgFHS5is/igxI
3PlUtbTnDHdE4cF2wLyTyRgJhE+UGeVEev3hGzgJy87MhwCNdfOK22qYoaz42kJ/
UrkRSmyeP5Qo3LP4bb1ScW+TcFHjHij6dbnY9sNFp/N+7kxK1iUimVHMuMv6CY1h
V7vF92FyzXNHVWIs362cxVRa0Rp56VFf5Dc7O0XYJcvDVz3FGoCAb5Gipc5VNlGt
IWOpRCfUnbTao6hn8+LbHBkgCOw+jsu4BU0EBrj02x9NMKvO09uABMDZP7cyu+Qp
CY5tilSRv4Dc6XdlTbaprqIeDKv0zwr01JPt3PRm2QgvJcJf+RC1j1bRyptWZ05+
XNtWZs10k41ouaekD3zmrP9VysRbZbt7UVIED9ES1EIin87/hWtDBI6dTFbZ4/Hu
/p5d3abSpqqr46fsg/iaklrKNiGi6Mf138r442PRTPjog8gBkiw+m/U2RuGDG0L0
DCvPCd2w76Jfka7tloO4j5yrRZOJADg7WIj+M5pHnKnOpSEVqK/o7Eeo3aRoVerZ
x0nbSfaB0LI/5dQAGZ4ooXxRrB5l3KKNBMOHoZzGR+UhnU9+0X9BYhVzlkAwDsrE
LNY+kfp/6bUCbn9LWntazXau6XPGQ5L0lfliGsINzOCBs2XNoaMVnc2+sJnKst8z
3vO9C6QoA56zhsUqRBWpTkHi7HJxW5QfBPMH5WGBq9BiZLYof9988EJG07jmNyfb
tHcNFR94su8u32rGFnSodol28MVUXPuIE3aGQwtRuQMa05PAvbT7rBBrPDcu6bqf
RYRRimNtYKNoYd/odl9pqp3zrrUbkLkuwlVbwwddoWtJkFORg7Akpop6UjepW0XS
oyT/v3Bmq7g2Mm6OM47/OeGHO40Hu2UZxK5JyL6zoJKu/xBcgH9Pez2jLg02ts8/
TLNaNQ6zxbmJbTONUnjggMkuRvXGfJDzRWJ1YGSGCj6+0qfjZZpsRyrZBC8QUI8M
eWtwHxdvvoGmSwiGVdiw+QnWXkVzji2+GbUViYw04Mr7rkSoKosOSsRUw5z4kQUH
t1PDM7m0hpEK8xuX7mJvofenzliWv9bz4+0OAbJAGEwPY8e+8Dsy7r33whYGwin0
/Ck6UHtT6ZhZIOMn6ILld8ZJUFhWsh1/vmUN86ODFEV+tfmv/FGy7WC3g/V8XP8O
3lBcGTzA7uHgrd6tcBKyV14H9uQ+V4WmgrQDXPgIvWqDhtDa95wlebOCAIF2E7AS
S+SJjo2PjtPot3xyo3raqkhKqfBFjEGI+ZH0avIgW56rP0nl3ZIxG9q/iw1ZifXt
dQHYtTgH4fqymGow0VGt5zfwzb2YC0bSHFULldqNiLWmr9czdOrXJ0/IA5SaaiEh
2jN18c6WW1hUt+Ngtv/iDvYOkHQOD4g2LmjKvqRKDuzETjYEX7Zs+jTLVuG54D0l
uzby/SNFFfvlZf7bc8cuvMr1SmJq0VgWqabNGO8ePX00XtSmpqYNdgMsXTmhSAF4
QB9S6no4qM1eZ4xcsaW3brR9NgwnVFJenHepPuHXN+JCo2V78J9v2EjXRleMJMOU
TlYyGE1DZtL0UzXX6LiV5GEo33KDlXIoNAv4yJabJvXK25UeZjC95tRrNg+YJi9h
cfnSotP3VAQeKb90kd23GibvbF+kYNU+3L5TgLzdohS88cR8YjUa0nL2C4usnRTi
kpcp0Gz/miXKINJhb4Lt1Q3cLqmeKHIntR+pXP3pyXHMxIGvFglxJdpYaw2FQGUM
H0JNYo6CufvGGUGiEUm72rccxyb1riPD8olNAfnG5oCNeLtI+uXMGGfQV6QCLAjq
5g+Ok7P4Zi9vbHBQltiJY/OJEmwApkrUADemxAIs1I8a0JlIT0wqQjLG/vIFYbP4
LGaISsVXXavywtHjttdN8H+c4j4qbqJqjRK284ibVjOmqtVuR3J7Tsri8BzCOlF3
G4e/gqSSCaYXHv6oAAlNw25R7jiR0n4UUm7Vckh3B60l9VWL76vIuucRhWvPSwoi
jcxhW0FTWVOmAnoFRLX6EgX7HiIOqQg/ZybuubL3dBWbtKVXYhXm++DDVyulkxMs
i09Xc1c7tQIjtbFHjyYK+cfLkInG+/TVxKxvKqTuP25CNp040kd6CWscUCn5HMwc
q/Kt4ngDRLSttiLjG5Fu7dzn8NWlR/WajEanQBB+0Nn+j0hGKVrr9RzokpM+c6Kn
cElWVhwJdIBbKCMuU9fkZA81OX7j/K5fB1CAI2lnHz+CpSNNYfGTxekgz1jEp5/4
b6Zn21DBeH44T+YkNSUjCGSMVpnFKnmTn1xQMApaEMoAo3pck/7gITafO2chYOsL
tFT/bUtRPPgDBVLlcyxbomuXmrZnbxIeva3oq5FMvqDkS+s8MMytLyVKBgY5Ohip
9ppH7KRHPy+0xe5WHFlUgYn4bZymDxlQiEXxtrK5MhyhwrA78BdISbr+Lnz4+H/I
QGTd63wEaBpDP0FRGZ2Oqr3jYmNDHFdMbBuVWDKukwNmhndK7fiV3uOMq5Wacs4v
cl5WByddHK7MQ10nA9JoOpRJlHK26W3dpg16M/9guBRxCFGLTQ4OLAkwZzeBhvmR
DYR6uVOaBALL7XTKA0quDG5oVlINx4GbNG4MWWYcn0Phrzfe6I7XM2/4mYuOeVut
4JMY8+W+dwanTBTJBfTTH42hP2bel+p7vDk/ynqFWjYYWWhvoBI5ZU3pag1pusT1
wz0LGVn0KVoQOcxSxuFiC0s19sjudp5p4yLnYcUnTmUzn15GzD+mPrZeuGYxEpEF
KwAZd/p/EQTWqEmUb3LZ8oMWdK++nAUybCAvu6ayO45P79xh++1c/4Q/SH/vY7gH
kdNvycCyS0gZ2ZpYJ4K20241jrPTLcJSE3tR3G8grCGoB2+pccrUN3IuqxwZxI9G
PO9T5gmNY5VS06inmPlbd9JZRGhsSc/FkdafBdu1aXYGD06t24H6e79RQchqaRj8
w9VQARbk1I3FxPP2DnGdVQGRA+3VnNQu915cAP+ZCgvSssvpSm15ZzKiHajWu63q
1jGcSjtu83q19YBN9hgtPgGInhBZGRi9CwEfOXE1CB6Vcc5hnLWRTHsSASAvdJSo
qB+ftI0GeV3oIC0qFtmhCGWfETfmNZV6FoVjJxTzYXA9fREYccWzqdkLb5luhnSY
LNqdgmHpEa+Zt7g7l07aR9pG18nkqqH3vPUtRH4vFAwZupjzcZ50IPgi/p3nUbaW
rDYR7i+SyJFZnQh1fExsFQEFz3GbCqJCSBXFY+R51q4bltJxfUolufFTEiC/i+W+
UYfyo1VfpIg/LGe21mog9J4gBQnUB6sgwtU7HqZAQGKFL8jtKCXX3IaqNZMIcl4O
DnIo6O0qA4Tce2VbhseAzAWRJU7pCFikANV5bDZmN369RlkNXfKxqa9ffvNt2xEz
pW+gPrrzrX+5b06857yncM7pZ5OAG2/GXC+z635E/omIuDWS9R8SXEngYK0RqyVz
vhagcsx6mosrOaHELcXiFBJSlszK8CY8W4Pr7eiq7CMrMcE4OlcsEg/Xf0krd4V0
pAuJneD4BucYYEHLerZaFJMhuPSaJFTyj+m8wQOMwsF9FFj1C4AJ/RJbVj/+V7SL
BQs4lfiUdl3DIFmvrwocgVPzSPozKvpEzKs6VlqOsXwKJvMYmo7nKukSe5PL3uKG
LJJ4gQqh5uAGaGj58xBQjiaoeYUDjqnCp4jC8CXeh62y24c7cv1FxxOcRg6E1HRR
+LYG/2zCCkx0xArWWENDOIB0Wld8CdxcwgOX3KMx7Y7Po1utJEp2l/+aCPy+HRcI
HqtbtEM/WavKd5Esg5018AjGsaRwv9W4PnF/61O8WcmJ4NmCENNK/bOAEr3s0so2
yf8YUuHDbUJWLLjKTraJlOJrbp8hRHIRDnaKE1JK1/ub1zXPGoHZrSJL76/EAlRm
pHACg1i+6QxjATJrnGiuSu6hKz32s0Agi1xEi61RjXeIMuqaMqt8a/h+r2lrZJKx
fRmjCl5FzUVv398KTwwtmUegbRVvaLbMrU6H+jERoqh3LU49DoTEMnG1E981csta
7PYlVxoQXInLCldHkHdUf2e4qsijULTRfZIaUcLcTwCqQ+zqWhaZPlNP+A//zYJk
DKBs3mlQIARh1LT3go2MDeGPum5Go0DqqZcIUqhheOeyZNmylOHX2d3FgnxKO4BK
L4kiNQL/gpr/18T2Ld7eOFDNqde7yA/YvP5AA2ukN6zkGhFfmKLT0R7BVc74eBqC
tAQfCGYQJ7zPPXhyfNlNouqC8SfkbafXhfuTiq1sXbaOupeCdyncD6Ne0ZUBW5ER
g+EuGOY6sfz3F92S9OTmFPhHhjiGNphmIDKFd79Upu+qk4IOPwTQCXY4flP3E5UW
aTU+WD1MSGCVPfLETYgPNWNsn965Dwh/GrzsW/JqYpYlyJfIjD+zT+baGl2fNRBs
Uvt8giZPZyUA5OJAFCJqXC2g0UGX/v+p7ey8HMQRUjwMvO4wfYnFVCrEvOJsGwet
R04hTx0ybzxS7GD+sf3PTi9DVtszGkZnBKuDGIJM6lVSDpnCFMAKKZ25ulc0m+1q
H8BXJEFMiY4GvmGtBVz258Z6V8zVuMGRYgG08WS0TJKBXvxemD3O2YCHgRB0bDHS
6MZTgAFEQQ1P4Ws/csPhhFOk90l37Jzi0I1GxTgYK+bhwMhHpeibDZwpDQulH57z
YmyWsuUie/1T0VrtsrlZjID59qIyWo2Inw0QoG/Oz6II2uO7+lGSxJebU+NEjVRQ
XSI6ekNYb8Lo1q6WfprjlB4z32MABGhErUelGL7VM3CCtmZEFwcZDsZMuHIyWzKX
30QGPCVWoTNZmooh/h8yQslJzwqDu73fsmMHWQW3qkWqd9fCXUJC6B7lRDCG9onb
WESWIcFzIv7KWmfXUihjQw4tbpM2yJmQe5GugdnDqE/55H6/xnO2RX3xr0H9Edbw
/ZPskV270XNx6XcO785UYuucKZmE3hnncSVkpudtkOe2v5E/GBwIr37WsLjUOEfg
H30RlK0LFG9gDVtj9c0yiaYyXtx6xZGKGyEjVlQyfwtA1YZ24JQbRV3q7biANUqM
yTooLMxL63H3oxTK/gB7CnTh97cQbK99waYLeIzRHHa98eAD294IiFaiIwbXearA
gM6q46lr38WX5q/0u9ALwJcqPfoJcnfyQwTIExy0SSOVqyF2si/fi+qkJhea5aXp
UPWbHHX/2pyYNISMBnqXbFpcNQM1ywlwTtQlx7/evzYHZATARwJ+tvGhN6UKLX8V
fi//PFSM4PWbPhU1WRP4XWriAN6d0dWPJwG6v5vn7lJwUViAiSmo+dg1QP8XAa6s
6jCzM2mhG1XH1UK86EQ11ao/0jsjvKhiPhV9b2ii8nS/6Ekj6U0qlFZBrYpD8dLI
3a0Sm2XgQNSY7oaSOAh8Cdl6eUf7MKInJIiUWbXx2SBmD4PengSdfWK6A7zRnmpV
xhCn6A8UkH5YVtcQqzfi61cKspXoe9dwYhKFH90jDp1rr3noR68/JRDydR509WV4
f203sycu4iC/LvL7CWQZdXLStJ5d6+j9RETfGc1CPmHHDkD8B0FbC1LDNvC21y/b
M/8NSLHoxcJdBih01jwhRmL+dh/aJZ9MyxN+5qFm+7yDzU9E/LUPbn+pMoQ4B/Bd
opWTaAFiXWh1HkqIiADxlcfyxtHiwc6BaF3NASsLB4pQCrgF0dEir2BbFCMPZ/HG
Ni1viadSOyq6eZqcBlMAbvS9r9MmepESxC2p+2c4asWTvwEAPrWZCiYPDzvCFbA0
VsVP4lF9d7ABjKoIgrRrzv2p9XQMyMb6M4MPJ/7zTZ5Aan4ujjkTOPm0AzwOtgvA
Et1Ay7Dk7NIqBZ6uC09j7OYgCdpLHvntU6pDm6Qf/abaO3VaHJzn3lB9KCRBPzep
+suH7Oot4wSsDS/+45u7jFk2Qz22rq+JBrIebozdhNNbGrHREy/DqeNbZlsraEE0
bBwAtAHo/Mv4T44XvY4KsrpGNU80Ty9+Rs5Ci4Bo/x9x9/CNMrrsYb8vt+vAWEUh
SbeWMnYDqhVFYUx7GfmfqvF3YgL25OO5rEcrzsu5dkRNC+vvT/hD8SkN3rxm1dmP
3yxJhyP2AVNCecRvyNqTaCNiQY9ccMQEWOs0k7CjZyhoI7wjFgiwd5lIVxVqrZz8
wk9QcrBxeAJyJccZ3aqfzJNUXDh9fKm/euMSKQMbJnBga8+Pd5olQppWZOdot7qd
ScxqNfD7DwgOBfs9BWT4592VCqGtq15Ryj1nxCH2DT9wBsbmw4yqpndzrLBzAtUw
7eeBPilhdFRCzl7seuoya+diRKvkNrhOFokc2DXFGYsCDIVbkfluDOqOF1uzmA1Z
Yi6RM076ThPX9XkYQ7yilOkcK9ftWKw+HufkZSU5MaPlhCTyUVxs4jJyDwRZlBRl
XmeQ4OifKfLacUpSXafaKs2vOU2J/JdQ3zLW1VfQ6GNYpM+/AxnwDYrmQbFFq5ra
fMRIqCVvXTM9TH4x3ByxKSnSXETb12cUAQc+G6Gg6K8TWhmgTRa76wsZb3cJL7U/
ykYJfXcJDmBNPJAN0xdX/6yxLRe7o0JaWBOVn9QXhms5htUgxX3xT9KVpfsPfzR0
ik9161Pt3K4uxtYYIGOEPNPpXnfek/WOMWtaVD1RyTh6awACDdYHg/xwK+YmkL+3
1WwRD8FeBEGY31CyCy6Q2Rdgb7EH+9fJrr4lkfozZTqEcsev4AtKJYBLcg9J92f4
1Nkwnd18myG91pvlhr9TrxxItKYmsTQlK1b9qj3h/RWSoTfGNfBPyjxk2lc4iXiD
aAyiSF7eRssOO6hLBJkUyudmYMDlqCtKKd9fFhQgMKmqLco5F5Syjyk/FV8jfB2W
BzMAlj+o/ezi8t3avADGDN+aR2PAH5ioJixZ4FMCCphU0QoFl+5U19o880tz5pkn
XhsUSyy/Aa7GMTPVRoBAf72LHgx+tY8yxeVECHjTtBjsauTNq2sr9Lhz31PY1MoO
0UDQpTSvCaKqfil13PqlhC6MqlQ+b+7fKwGmEL8Z3nE6trxaffSGyVK6VixdW3Om
/iPS2QhSS/llJVUURVKkBMcypSSjx3aQAc5EulbvL5004iWezYO/LrXfRMURKOj/
doX5W+6T1el5SPQNke56NjZCDd5wKZ3EQB/vKTN4Zkb/dv1FfcgtpevEzVQo3phM
HuWMA3htAl31SwG0PJNAYKRPZKjFfAir3md3E8vW2Sk3c32gBJ2Qj5/fg2oDbyUM
nSiBGD8y/s/vtSbRnsyEVlnIJSFemRbBni75eIZQqqossZgLNDLH1qgpHlT1SeKD
g8A49XLgjGLFf3DuiXzXIvEF8eYCGUdj1YmRFTccOrjoJ2Y9bmngSx5qcrVoyQqh
i0FnSA1LnFfKU/xHLa9sLOZKAJYOESQaJCeNUkH0Eq9QuQXg9IqbumQ65hwlR8Hz
xOu0hxS9HRYu2BvntSfQP0maBOY27BELc0+ATEMdR8HsZkC3b4af+rjfRvv7r8sX
fXwxZCPw9BD6k9KK5+KqmLDQu/imeLHJRtLtFZHMPESsz+bzxVHW4J0HAiRDrSlY
cnZmgXt5Kz8sZ2tR8anULU+fIxM61WEaBiosAVj4OSFfEZG1gfmNIncVkjQgJ/Vv
qUeU6bHH4oUIqBpGh1VKLddaacRVbfXgcbmF9Jg2Aqz7P/mdJFMalLKkp5OHepI5
kQ4SPuR7CWIUnskK1N52KUSxvqBTQoAoAdk8++DOjY4/e+FiNFMQ0XJaoay5rKgj
JqFyOuFBPUlamvCk7w6BE4//wNaPJeFGFA8YNhJ+84nmxUIZdGt1SABm/9x5RLA3
mIa9ulVM1PfHek9cz10O4V6H+gdCK8boz+XwS7wT4d87RewwkhmNUW0mDrRKnxHf
YPnRnF10XDZCFk87pUQ4jVjWEGhXpgQgYjpkycp5B/nW5tEsIja4d8N0DHS16Vqk
RtdoBlbeOmtTL17OL3i1MQkOHKiMwB1TpYm2PaJFXHQxYqSm/0oWY6sZvZ+t5eL0
XluPGPQtuqvEQgQxOlVCuzUFZ+xUYooS7+CFAhDB3Lu/z08M/55MWTYp1nSoBaPX
cVWZUi9ZaBaT98B755nKbQNQNNe/VAyB+Y2a1CKMfP+F4Gu+49qyJYBXGlwtToC2
dg4EEGbQvzwE9wC4rttlNIHTN672xMprfV+Ehtk9OSbuado8uUNWoGKED5trwHBa
B57Q6myr58eQDgVkrVNpGINxgElHCMyPQu1VHvKncOnl0WwDHRDshCrA7qJ4A2oD
fxzc+3JZ58hHYh2P0y+60JYnaq2sN5VwSv4X5Tu6IcAm3fTvU0CaMhUoCyUihJFc
Vfh8ccdm/5M5yUx4+pJxrztOBE9y023yLPt/Qa+YIWjTjFyRcmHvyX7RfKnQIHEM
DFw1vIQRyZYZHs70KwGZe2Yo/dby9mJSSmsZ3iyZE/7+ydRB5231hDMOGoDLmFkU
nOi1Fg4Ckq9CQIq99E0ylMjyv4NCrRtCpfkzdFyvdlSPILmy4rkue563jOais5n5
iw1W601EAd0C3n01pF4HQTv9VQt0l67YBGMhDgWnmsmeT9pFVOn76SoU2vasWsmd
5tA40Z8n71YZlzVyzMhaRBVppzRoJjvLk2Gzl34BxYK7KombZcU/Rdf1KEMWwhPm
nmJZb0ucKre60IMwfywSQ6sOOljUXpn+QQHaGXvt9bwQfpLmEVebttPdh/PkI9Hf
5KZupCjwjxb/1TPyw2WwMUUJ/3kid4InFGIZiA0IjKv2jOlhoOQz8pU9C3aYvHoF
UiC/SC6YKn4GJSB1BkvsMAhj2dcpQwbH+JFQJYs84N8Wp9cY6Rij9cw1RPIVXjyY
rspcLYsmtKdnQF6bNdoBuR0hDD4tqivbG3WJ/FL2l5+1usxbVkzxhO9CH+okc3Hn
J8fXNxai6KKt6wGsPA3DM4u0kDmg6KP7b9wxivb9/I2bAw+Y3HvRS9kidxKZZ+FD
IaBgIbhOtgBlTjU+K/sMf8WszB+N1g7Cs4aeuZr/fhaCQmgRitfjLsguWhWltw00
xWPufKMOFDWejUL+0w7siMKLCAPP0EKkyNBMfQ5OxSxIAKjU/rK6lO+Zlz5g4On6
3dL2o6NvokFe/PPosjvQgBeC2vzr1Jq40WG20hgZaHFLAKC7BkaWDtEblY67zmJ6
bw3jCsB6OD68ipwrMvAER8WYkhJ6FfKSBYAz1a5ZYEYkhSrUFHQLPj7PRSykieI+
Qf5bnBCGbkd87+g//zEUZpSJdqLxLyMDH/G05URKEpwxjKXliwAmji3SPS8AZ84x
aBE6zEcj9I0BkE5D3IjsPUAZfEB6xaiDHzxYbKJ0DHMutm7Ht8qWZsaiPIvu0gI9
C1p3Y0Egbbssb5QD9b2h/cQfXrT2LBGP3qLjKxNrLUdQczIybWmmj5ZMIEOTTRmV
yVLhsiyasir/EEgiE+O/Kg/jsVjGXA8BqHbzb1E+5KtSL9TWHH9yjChPiOt7cDAN
fTj01iEO7I1FfCPVbqETuakfV939JG44rMKRkzIv95pdF3MLAo5RpRWMyxQLmAri
o2CjFYslvuArfzujluUoFWOFyvK/m21aGEg2Orf6xe2lPLr69FNz/S8rDUiEY74+
hFjVtbEI6niha0eIlWEEKPnzYnsdz6msyVhCUayc9w5uSfJqsGN+uGn7oFOkyl9v
TMtORraK3YnEKbSZGVAJ4PVyp5em3+4mi6FOPKYRQsJLWS+S7cpV/GSSpSBca1Th
s+9g5goYuxgf8XeUjEo2zMedoUQ5GqTLDnVDgpbt9+h3cIotQSw98//QfbO+5tbx
uSi92Uu5NUhEzJvvmZ9beQyuWxqPdOUoY3vi9PdSEtsU2zROVgj2nc9igCO8zd0O
SF/pgCHFKXQrMDx5RSFzQeGS7pHiU0pmqRf6eoDgoixyB5FcUgzxh+Vx46lTngwS
JRUI+yclwLUzQ5VuLReguNslEu880XtcJTsU8n0f5stjdYLjYMqAZOt6hEiqyRF4
cM3jP/GMzpYg2BumR2qxvUOKM8Wg7aADRd8BW2elRT1GSoJWKEXRIaSOGqokZMA/
+Jqhmed/2nRyKpox99m6wjZuzZa3Yk+qIFfznf4iEQfA5rVDQLgxycsoworBTJ9b
ZtCV/Z+xaeMkxHhMvUVGKCDjRmw6Wju33OsyCxUnrGDwXqEmOhR2niyGnjlxld8T
jOkL5fmjnfbO+i0YsW3FejBHCeyrJA6Si2I4YuJidpxejezIJdaK4P4JMsGZoSE0
9VjZ7/Yuca73Pcu3sEitBd/i6eR6hKADaw5N+HsJZv1gd04bTQUHYDZwfFiV5wog
MjOZ6JqAl4rVZS9uZD1kGgXWn1QhwboTMrUA0sQnJVS+0NopYssPeRWnJe3DAqcP
cl5JfKVmFKZv9LE2DsKE4GYJPKSSGrnGvXdIQlHxMTvb38pAtAvmHw3HAZxSKj6p
mJyNUI4lB1zcyUkMN/K/z6IP5D/D4c/Qzb/ABQ3Y4p7RYvG7JpBkzZZ9jKWYRqZv
DXagdXLKGn/xWGO9Vy3wuUXFrrRaDjVEGJi1mdI8h7K8VdGgtPmKWpLLafu2+bTB
VCI0Z2oMnELiOdZZ0V5YkRiVuIuf/WNd0W/vO9Pcc44Z4xc9RtIRx2/kMAr26m64
FYXrORYE8qzL4bCSH4qpyBXCJlAalolbnYZtOSI4CKHXkhFSKFkAlDgZtNDJ8p7H
ceOM7NijeXKepvAPuDqTlginb2w53+d39IMfE7JclWAODuQw6asnr3Vgihr07IeM
Dn3aV32f63vd37DZyY174DsNMhsLcFMwDkXAMdADoEOpcguOpcrmkqTaeAt6XgUi
tX6DIhEeF8YbJaPkYhTYTqN8yFfTZ+mNlRKqzLI7CXjrd9cuWsyV+DSLHecJo1Ts
P2LRmGQH9eOxhZekZN0sUN4Pm4VRLZzX5d//sCtcwG09WZKRfBC51iRmDTrRVaXQ
LjT89Pv/iiXg1GH/y9LJf8FCctrGEwJhTPmH6vgIzlcpdJwR+2jCdwEvWjpgDDX+
aGrR3JE0/1LrW+YqAdV0AmXL5HDTMtzIEhwEk5qWovHhX1U36VvkZdcCJ2ElN3vz
zqQPRCaZbXsIcEJC2AjUC+vaqPPm1CEbEzpE9+XUpVqVxmfRmN3CQtmaC5Jfvlzi
WEBzu+Thr5Iouh0U2tWut3Z63cy8P/scTPf7odWlT+/w5nAAn2iTusMlG+C0d9j6
rBVi1cuzDis0HRkkoVrpLKnlHBGynd3AH3gXrs+g2nBlRpQ0d89zTy5q+rTDOkKI
cy7ebUrWp82gxkmKU5WCQrID0dg8RtLN4igVuBJ5sOSbxjyfQPecdppy7Oiu0vt0
hirfsCtNwrpQh0fykiRCfG9U9sa1ZXF7BWpjBU8Wdvk9JeOvO8q/sysMm0n1nAO0
YBkVyUJhGUfW6+ufjsLkd1kdeYpJ7rqiyYRoZMZeALbl22LsTDq/CtjrDyEzUkRk
MpKMTCJvAgAU5Qku8+YoKOHmmmV4I/ckPkX0favkMYoTg3OaTyWsMJbPu7ZRZ0Ez
9gQ3O/s28Eb/qOE7QkLXcYNRe4vINg1IJgQ8HaEMdy+WuSSogjQlOouIkgwC/c/G
TfUJ5a2yUetvuLEIc7T0+Grn1CIkByiVdMthK9s4XvCT5+ySGgQ0VfmUvnuMKYbo
9by6KY/GiJZeQ6v+sg9OSfxLS3p7fzMsi+IBxmqbYsAzsAfnhwA7zN+vDPbUkC97
4uUVf2pb8RpEHF1WN71LKkjvljMsskZUi/Bp2nRTx02xd51JseRhF3hR1dTG2dYi
njov9XdA6NnJi9FzYMkruzioG88K9k42TTfnPXMtNFeRE951MRE0BuBUTKEy3QzW
Y+L6nrtmIoDQNk6Xi9eqQBQfxjKxaS1sYtBJqHMcjxKpNKCjjieZW4UvjBLFO6E1
E7c/Tr2/+gzH1SJfcxVQPxObwIBE0n//oMR+vwxqfK9cWLS7e+NaYK89BIUwIr3k
+cpJoyD5100GRU+nN15RogiPUpeHGvnTPq1Yz459eEVChzqnrPDWxjFOTnwRWr90
DnIe1npjn3fD6RoyQxGr6VuLK62BXpz+f0u7ZFTN2HlWnWkzBtQFkMV+1uJbT5zs
j6/W2GtlvjJDWypBSuG2lhudNNem3hyodgaAqcLdj2qt2l5/FPqFFbs0yPrrDBm7
/cMSCmFHeIqx1w62IR2M20yxpy3L8fyfCoCmRo1xlURgtSxzjsYpk+5pQyN8n6rM
npcsLtGZ10vOq95iH7EFqWQPPZCLzwuuxUFDiAGUm4aCLXcCUvqutpkxOu4h/PlX
nmCPAn5sxOUc86JmKgWksDEvtHvob4eiEU/bgatLas3EOG4Y4kMJNMQFSk+btpBb
W1olPYRNDleZ/qivpoJuXvnU5/DWOlsQycyh87HAnZ0jhayQbltRajmAKx1v69fT
jg/aBqIlFrftdhGeVTw517iEiKrTPj2vek0qz0ayy6vnXkeTloEJ8WV9rSREC2f7
kFupzBXi4Kc28Yy9ndGKib9d0cXG72gZnOw7tYD5UVSJ64mXV0NF21AQjHcmZFP4
jwLgynA1rl89vwqHbDC0nFnqIanncmlwkur/MrQIKsEt4les74vqiLm4Kneg/Tqu
UADB5jOLq8CsmIh+voDzKeLIfU85jvGHRsbAh6PZnfrTYWaxNvFTVB3acIK2bZcu
YJ56mnD/0JcoFKtGWrGne1labCcRVAILnDAXnkipDQNR2XXzcNNuTeqAqfES2ILF
PgVkY8I19pdVW2BvhOkBJWAxJUpa/DRCoy7FcXqozWdBJM1ozNBOu0zuaWkIAke8
bApgt6mFuDb33nPeHrimbsF8VHhaDEua03NnSBvp5mZQ+aQtH+UT6l2xpzm6oSEJ
XgbJY+x8frWfySvoaFOi8JsVqWagD9c/K/MrH5qiUPe9ArGDR462qmL3tDVIhcX7
vz9W1+sgpM5exOxY+LL8cRtC7o4fCxV9T4yzs4ldicuebJBvOoWYKs55nOnQBAn/
RFnzoUmeBaS4baXqY/DyItxgdmsQ1GEZH6OTcg2FUhP8t+o1hSRF4OCtNcQ+GJMr
BCca+3wi6P2LH1pLf1GZMvcGxrW+ambd81iAcbapTYEZYPPF5stJme/0MhqcGWFr
uCBCUTr25+DlbqFJLr9rqkZkuaAwrx1TrTaAgzE2D3Hd7x66kCX2t1k0aqnKhigj
XOAXlWcv/e0lO06d2GeQJ/8e1sH6P+EerX4ffY0eCwPKkufoltIoeH5FWsVDWrEg
p72inI0VKurQkrbNVRc4nJGxDWT2p9FgO/or9QRMvfauPJYyFIKiqKxNoJLqSX9S
QwS1DZ4CtgVUFXm6mgrhD2fuNMC06afehFT7I51CZvc00SPaDQIUKRdB0U0Awsm5
toDwMC8CWUGVgkpN5CdSYC06y0jd4Wdh6gW7tPYIQChBKNPTBRbivP38NCYquC1l
uLPr07HBxVQyqQPbGP+ND5KLS+V5vVhJNbLSAdYj4zaY7bQRrMJhqt0Nl8CF4Dh+
bnmKxHinwdrLlemPU5UWjZRVINjXoGwE19kC7/OTkZlGqQogci+3uDlJlgOi8Zpa
pglreeSuonlv0NRMvm9dWanHMIaesrS9WmaPYBo7sJLKT2kOdvxZwzM4ytyQK3pk
fg9R/XX//WU8Aim6XsaZAs2w+yxrGVKoYVCZxr44nOmILl1bDQ95t0RCWnGktXQA
YTDnue5ZTc5im9RQ4H4YnV5IHIcUry7tYFi09bV+P4R8qSbA90GQRNcfrI183IpL
tuoaB7LVHFjqm7A7RDVmI+rg4D2lqgpns0P+s8uRmFDF2t0CB/5DSMXyb2RvMlkT
K10C+WM5mRs/tm5nzVYsNThprstuyBtwPsx2Y7yreZXS7reEGJisIsXJ82fbMkw4
9zpYoE9CAL3JXuUMU3eiT/mSEuKqYbFDcaaWdBXVnv0Z2IMqI7y0cbaM45Oc0MJ1
BVbTETozLPPTVm2KxoOiwB061JnDk/Csh/7xYaC0D0uVbAwz6ZDUh+egDMfCFTUC
QtzMEZWj+KRjgMXF8eF+DOCGzB7UYNchKC1SyzpFTncIqOIEIt6e7ZoK+2koQ0m5
7tnIirYzXFgYDAD2gDzPGyJLa83uQio20n72Ouh8a0H+kA9WUy7BL+HRaiq0GPf/
Atr1H6SMHOF/UuGMzGcHYsM4pwTowRjnH3NKym3PHdEYXBmo84x7W+uTMSMJ5h/c
jxMs/GD9vlLXl9Deh+TK7dHiPLTImpOApyAElWeFmfgmTFofwQzljUBt0nkhDRel
6uPykBMzmIv1VELN3C1dDXOSBuRMxGmLuHV+/Fkd5TfGI8A2Bkw1RabcgpIRq9e5
0241FFN3XgmsrV/4QtFnZ71NQJU+w6sSHIOlONVvUFUJ8FejBzKTkaoMjPjyusiE
jqygwQQgVYusG3U+h//5wwHSkyFIwgklRKtBnktDxcbfzKsNHEci3QFA2zGDNT3H
UTj3tbHlrWHrtAo2zeaxxXQSrCaEdfNkTz2D6S+ZzHYYdGAsookL3S200kiiHbGr
lquFGnNK1kbq/d7hPV+oQbFfqgW9l3bRds/5y9sGzwJMotgATf8DWBWTXcgoTuvg
T1r8oZU5rwKBdAGvgnlPupLZnYk/VWMH9r8918Rg/L7lpOpuWJqfQyGl+iExougg
Ua8mfctzQnhbmk5Pno0VHx+kd+fMnkoWXPRKt8tLH45TXIT4Ei9O/ZbHdK6NnpQo
/pCUa+ekft9qymTKpiJwaKa1sGsyS6VS/XHPT+yPy9fdbjZ1/c5hobiCLFiGE/+s
SiW0jGXgOAZMBtTYbd2sdeJG7bTNZY22lTWCac+NZCNJBQmXDRoBWbhVoYriYCcD
BqvAe4XMNtk4oh29TmEWTb5OmGfOKkEVZgrQTdYQ5N2MUNsWBFJtv2DMIsBIg0DE
bbaFRriqjQSyc6U88mMELsbbPBIApJ1F3uiZDxivzSKst6mldLIZLUyYKVu8eGyR
6DLOvBuxTPVIkSHUD8x9dzGyicBLbczHwZmPbzgLQkNwemG+3v7tOSvqfXj/csbU
IYeUYqZNmiE6QMtC1ohN53oV6OoRLoxgAoG5vb8juHz3bGfxTw+CTfoV8HDcq52P
OWA7xQcNWLJ5CGYWPdqES+4gfRfCJ9pSyvk6p7ImFSwcwBUJBWTdut4yyjREJTME
5Be73rvzkPXfMSY1CYfYZsSSYsADpLYLvuPeeSXPuR7HlwjK+JZeWP1x+wAKhiVN
6eL9NiJ/YhEGFBVpE2iErYKUPw7yyUBHhZWrYOTszKMqgyprq6j+o2t6E2H6plzH
fkf8dMyYapeyOsnF6cIzLH+nLsi8T7IcZnTVUxmRRsS2FA7kPsFUnauwJZJb6LBh
t07kxZ6nYW5H+UnToWgVrTJ1tITE0bM2PfK42ypT8pE1fuaLDAK2nmtK/jv+j+YW
4hV+CP8Uf+i6UkfCY4HFjOmWqbC0MY3L2yLicO323Gs5AAUWfnVcXv9vr0Qqt3sm
q4UqUkLrvKcCf/JHmhDLzYiodU16w0dRGrVg7j+k3FU+/eYhbSM5oNXkLmJMgN5l
DmPu57qG8kDCHjJawL/Qk7qDTMhJEhvmK1Ug0DSP5CwS9agR9z1LZWdaVy6SJObV
nYiw0c2Lk2ZhpEi/e9pykVvR9d/p0IH+/K6b4O1wa6JFwKSjSmAzZdRKTniRPUsJ
gL55idvcrr1l4SwY8xjxfiU/p6fifVmbEjOONAJ5uhGvZ/ytad793tYGBNpVtIgT
gRNwZEGTdcnZrbc5BKgr+j2m8MaV4iAMaZEoB2ghfEu0YSUndKqghsZewFckQ3rp
8WFpBLwzcG/i9D47yjR3GLQCIqYoF6VqHBR1QYtPKwl1B5//jgmHiK8Bfqv7K1DU
nz0t06Vuv+fc5SEWCF0y4VoJqkTKQawfkHrXoEt02uIeZ6wbNa7clShtf3MVgkuB
aB8azld8wFcglEGZ9HoDz9Un1aS7Rh90qHdubhn4bgnVzHiWYGtzE1g0DtbsoMhr
5TeWMtl0AubnbC1iS1oH+FAEKCrA6ZeNyC9DU5CGr5fNS32LB0fZ+G/txuoX1m3R
ue6eJwGO1moxCiiuWU/5hNwJiIvVh7WdeA8+DdzB/J01uOl6bJDsvu+u+u4+zAu7
QZKOvyDaEj3hha/31WpRaj3N3J6s7Px+0JIQ9pHkFOZA9nCwS1ZtkgBPXZEmjtZC
QEreL/7kqg+8sbAN9sa3iP2wGcpttl5zJlgge24ODMQqqs7N2KvOHsqMxATRaayc
hKw5sAsTYi6LZnkDO+3KxwB1oQA5qkSsy+XZ9bTdDYY2eldZ/YMeMCF1/7F2OpAe
FxAlD9+heJILmKWVOWBn4OuzDJG+1XQ5givJTVR5mJnyUjpEQSv+P3HFd+KXzkU+
z6q1hqXaOvfixsKktAVuE9HbhnTK8LgXCxYv0JXRJiiiomvWsCqQdrEwLVrGBpdh
Ks6k42RXo5tUOSb58CXWjKOhVYQvzFh/h+JETf6xwIE5NOQGKKDiNdmptjJ3Tv78
folxE9dAfS2UMtMIMMbxPue/Ax++kSKkCwWeThToQY8FNueieN446temKWD7qpDO
9r95e2Muy76u0RKK0SeqQs+4HsG1UXD3MI9RQh4HEHYuup9lzz+fjjxoQhWIToZm
mH49vLfPNCtrCIvthWygfyxBJU9bG7SLLiVfaN9i5FLTOhQoppGguoGl0lQeDPJc
OhFGk/oYF6yXw9XdpWlnHfv5XzLv9yyFP9tGKqtD9hdrL9f8S+UArqI722iTulB0
1KPE2BaAmXw4P56811hpzoYs5J8DFmUR5RLBAqM/H+VD0Z+PHJjzewKP4DSO3avl
u6yA3/Al0bI3A5F0Lk9s+C10oOIw/iaU8Q/J6WcCVMHYbGQxGKOu48zvC3qkZBuR
zCn1lp+QAicLB/2xwQV2Nt3B/kE+FWa9s0R7FMe5jWvXctt/F1XnTLtFvnjn11yA
nsioDltnw46OYvftj+UPQZDm05RFHByPnJyVIkHcisHtJEJ4/ZxxDhWBmQluf0AE
kvRpoKHG1AfZmqlgMVJvDZHbdf0PHHQ+/OitAKS9He+a0LWmuiZUSmmteu2zin6B
iopcTouMaSl/BjXKpUtKCx8deNGrF9TuM/h9zZLPbkcHOkChVNdFKXCjBhnjzxbz
7NKJ6kPjgLdB4HYkor+ZOQoUogltVqAruE2aDVd+ITUqwOvL1b02rT5lVrRkYHJE
9IPdEoMiDUD17swcH/L7SRcuX+Nu6SiUJ2gyBTqqwIk0zvZYnCxqQwcG6kMNwZwJ
hRhyh4iE8ULf5fWCozYok3OA4JkbCiGC6dnJliw/ANdyB+rsTcKJmVqQnPOLEfbp
4aYvxccG61b5n6qpAUEwH2wAbGW4BCwz/Qfhch/jFF7imKAAUyBHOYEKS2dSgKx2
p1zGzatl0wu31/NDhr+a0vq4dCAoILcgYsLpcFwpiDDcAHy4CiraFHj4r94O8e/7
QJ4ju5epTJGKPM0rWlbqKf3NUc9qyN8P+G7NeD1Lu4mShfFpxQXDPuXl69M8NEHB
xucxuiA4Hga9kYUrslFZlFBz+tcyJDT/XD/kbc78g+IaeZNy4H2Y9X8dwmEthiOQ
qwPmNAFOB6F/lfOxv058zwbXmj/iMKUF9YTm2Dm+8+Tt7M4MwDQa0aUebrOHd86x
0dg200dlAJp+XUewhhzjRZQKmZbjGX7qZpe8C7dLqLO+tohMGj7J3mnM4Jxn6NuR
dl4GZMrO6PRw6m4w4LTrwOZzaqbkvKX3k98YSXxAFhbXStwhJPmlRWcQYpNs2YMs
jBXx7Dr0wXDaIrDznGz1Dpi6hEdilFbrwW+j7gmNMTX9jLLR2Td87y1vohQ02PEv
jLMqDrqhgGGKLlYszmJdI4jiSJ1NWrD4xajQmkjClrkIJuTel4i03RawZ4YD3JEa
0Q7frzmMMgDQTbcK3H2m8Yj0i/bkJHcyRJJlfqIno5w2kdOXnUIdRZCL0soGDTD5
GsG0lJlOAiyMrGAXygIIgVwUWlkN1C4HHhD1aq5KfsrfOA7Yu80RiReOsxc3H+mh
0bFDw3TKfJVyGTJqqAeKj9mMkN1RyYAQH+oSWlIk2F/vD3/aqfYZwGGOcE7MAXUw
tFS/yH5XxqILtXEvPzVS/kNsF+UEIrxmMPpZ6qyA7EM8PITg5nIL/oY/8JWbxhvm
Fhafz0suTCjTt8X0Fx63uo6KvkuoiqRzZ5Uyk7kYe2veK3d4gjcZmbHS14ZBkgg5
QYdiktiO2WfMhPA7oCUNbeNAASSDAuq2gb2uphz5RKrbDB4HQz3Eu/2rnF2is8BG
UKaOGbCiiuNUO6yUKDJR7BrQALVPDGO+ez9ESUrla8zlrZn3FRn4ZbnMbG37Tfl2
DN4Pu44OaJRoQaXn4FPZhzP4h/Ll93lBbbfT3V7HXj+NWsw8sVecz7ADVlyWCGOV
1Dxj+rwwdEDbcn1sf96+VEu/s3m9KpTx34KyohUhFpsLuwYAMRrrWpKXt7eAwG9A
XV5GiguII3t7hkin/0KMHXuwGHU778wY+3FRh7dGIh5DvCclMcpKVVhLKl05aJym
DZq7roY13ACvg9Cak8C0+f664Nf4zS2loMyrp9PRcnpOjTJmv8etFvJij5cQSmhC
6yiZB50sOL4Voxj5HgV14k3haPL6D0lQHHL3jnX4iUUbTf7mLZ6KwnWEJIiR8s6J
QjCY3qYMfavLAp9q/59Mya5jESM8C90JF1KRuDQfRykshbPtfXn5OaEJXGcV6UIB
e5Bpuo4bEpSTfIE4dJfy3Jrwh1lCjYd2UnEvMCR0+rm3/XKY4rVpABG0Fo+6uW6o
TJ3pAg9vNdZiSWl70Kmf1y5wI4RSTQ9CH8I84WZtX+Eg+ctlQtIa9VcGQ8UHTCJG
oRDO3IR1OnQW/1vsQLkRQas3w3g8Kf1aFhlvD9CGfZ8W+uQSdpjokAiiJz9ybPCd
nL9xUUTKS3LTWllgM1GpJRAPMYVlN3VGeYg19xEbpZZPWDdNcpgzHhyad321jUck
u6/50Lx1Xokn2a87QW/TYdpZS/ATfBThavqWSoSxjC7s9CL4ga490JilB+TcV35A
YvXsqO12YWARrtd+j3hOXO0wIEy3Tk7i2y/3IGSX/TAbdq2GB6E4qhf759xHUqlV
Ge4a2KytBTQsWdU0MpChSe9EHjKZF7jJUyHNh8qHuUgUa6ycWLiZhGvo+kBfQhCe
GJMXfdGEadwXpgDOYNFMOzecaQzKqK7z4F11k34gMtHcKRucvy8A1AbIH6Xiw8+H
Uz5YOJPAu5BuWR0d2ALSFqovyoEcozKmujiohGPK4SaQ5H0p/arWnp4S/sGR8O+i
y8cMMQZ8/L+dcdm3kscNs1XsoMT2mqEUK3Zsl/twXZm0oq/5BN3y/V4YVcji969o
bQCFlDRRo6ptg1kaQFK90LAcwyMGpZTnCHCOu064h4SrvcvVl8PUF4LhTfCE6lbJ
szPFhjoe3DUEDA5vtYfe2+49edmBAIW3TZm9sYeNc1H8F7MTxMkxF7w5LuD8z1eU
ykFUlypzJdLCQR30ZV/03Mq8udak+Ayb2mVzXuTt2xEiXI3q5CEaFTnyCG3xJna5
MOHGZb8eDOHELQJyLuVUnpak1NlQHTCbs4BTt3wdfO3wSlQqcJuOFnIblQ+Q7Erw
dQZjdv0yK7RV9ZTmSD8uFnnho9vkV6S+7wyE64wweY0N5gGPI0aWf/UpYMGG9K/r
QSHsqqaL/5uVkG2jThJ3vsGrPeydMuvUQCaSaiS3/PCqYE91+TfsIKVdKYbVvw09
LiWtF8XihIv1+Cnc8aGiRjXxmyK+8J0r3uEEfglGxzx4tPf+NUnD+wzecnpc7FQj
1yBzpNIvx3yPh7UBubgwYv+dnUyeLkG68SGRdYKdhvKYLSzoY4P8V1IlDL7kPq8C
6pcZXeR/zpLZWJrCwuF+jfpzpLv6mj2t6f6rJBHbUxcBMKjbFbHg4nmv2s91OOel
q2cxYEotT/Ux8otwuupq2rOkgc4GpYWlRZ8M3LSLVP/xG8vXAeTL4lPoUOqYaj2a
yQgyLlGqLjl/3o/8foEFXNHO1Jq9a0hBCv4fB3+rnvBQsSDveaWhfad1bD/AmucI
eMgzQlF/pvMAYLakfGk0MOACSx2t53s1M0KbWw+XYGtYGAS+nRZie3HOy5JKNq/R
QwWJZsLD7cjBf1vYOs+BkpPf87tJbZi3gKDfT0E1XsEl1msde2GvNK2kjyNXSmL2
u2lE+RnaLrG4WhbSFgeHOYsix7BOSqvkG63i2E7kPXOGyAuznOXpomq7uOm85bS7
TVKglwGfo8C4yhOEtaJ+hSvpMcxRdfs5FTEsj8fbbIGvDLMXwkU8e+ZAqH8mkWll
gjohKF2E1O2LzzddGmmpGaujcM9oDTTXXZ/9FWmlVqEZZbY54o297HswYj+V147G
Saqw4CYSpd8ITmdGBU7bXLIrmS0G5gssn+oTrsLOKpShY2Yb7nZqbNHi2PIImY1c
vQ6Apv2DxUBQ60+gz6UboDmHPb2jx6qYtdHju7KLIB0a0sLPJnm6NMwHJ4LcGb90
SjMN4fh5IDwxfBa9C9Ji/cddRT3buFBWJ/LP6UOr7a29j9keba1wSyC/7H35xH0v
ko0NdzBuRTf5YzmL93QDPbTxPdcsyF9cEBM/QsK42msmmqPlGf30wZcfE60tPn62
Ug3rT86gitWQG6ys3uvwANfpSWIWC9lEJzTLnBH0Mywi7ia8lSk/BFwozZftZF4q
abOT1GzVC/JGZrEI3XmZjjUnBkqN6KWxLi0nYGdzhlklyTdMWPBdBhLJtnsbT11E
1R1kMb3wddHIZdN5KC0N06kX3Qt6WMJhDtBIZ4mlNxs4xsUtIeyE3/UcUnyYnr1M
HPdgp0LRyjZFKs8kdVKJHo6LFPrBmov1KACg87jkq0YdLOZhYk1ztEC2ib0Vf8t3
jWjx5B3XKguu9lAxCckQrxHil0apTl1G9m3GJqCQ36KqjmqKuvNNd4KCnXcuiIuu
Qg2tB7h7urfGdlnnLY3eQMrALuuJ//p4MueqDYYDlcnr1vl3VTA8mqZ+xnRPWeMQ
2JogyZASesy3p+on7flKMx31Gh5rrbjkReOM/VeoRH1PB6yRASo42Qbrjr6RN5wn
lRNdR31/zBkltLN0Y85+7ZL+ie7AG/slk3ZJI0EJvvTAz1hUxGSSbnIJSocUGTcH
aOxNJOZTLiOUJ5B78HHp6nIxcXNMLSS6nADhNrBYpLOVpXbWaFBYn41MIgaI0gZp
1ziWr0lz99Bt6Y/6HD2Fl+AcpSAsn636gQlG6WoSrMjBnUOSX/EEE44j1E3neqgt
Nry7ww+YtLr+7vWQ0m5RWNR9JmLmmegYt5GewuoFVkk/DppqJOqryJZsH88TuCHy
xEcBNXBXGMHinrIhQHmzOphBSp2UUrm0kU5xl/410Urx+Ohv1+yYdFfoNVX5frPv
Elvoi66CNiJCfkoXrOCw0nNXQPkOGmCeifsngLzCEhMUt6SsoRRzUTulg7ueHtxP
sxuK7AWXV2DvzigTZ9T+9wBJRh6oYCDIyhABZ8Viui3LG9T5zQ7TqrVmPW/X+2s2
KX37Q+6jLIFyEoCtQHt/oc2Al9iCQo0SBvzc/9FSESutrORvY6YBRAzTcLNQGRot
73tel301RBE0fjh/efeHXmnaj//IS5rpfw/aFemVv/AkZPOzAEr3TCqd8I1vWgfE
wruenbMYd0kj0+kxMnGRxZi82Of0PexFrUXyjO6PSZ83t9LGIRuNY38fZ1P+2p6u
rGJ+qU/bZ32jfzSZdBBQIcEfQMKJ9AabidwcO7rC0fcqWlSmi3/Yl9mwdISF73rQ
RrOzzfzWRRtvsEr5mHfgLYmbUWTDKgWV8IcuRUclzdDM+Ucjcpde2/wmQdR9vsHy
l29yqtUA0EnhF3UWGJLS2zjm3mLuze3ALyp0mety0vV/JS9VFkT+hKfyz6684bV9
sLd76FUt4bnDDP9iknChP5mF0w7mV9eXw2O0cNKty1BQJU0Qfk1qY4NRaqiFyT1Z
EWKh3+nYXBKBiEwAdDA0GJSoA2uKWZbDIzV/SHewY0/kAj8UE/BjPtTitiQBEp15
lCHhvDtrEN2yGJmUsLgItb6tUOT7BPjGKMxEzHiWKN6D6LyV1eyDpQPQ3ko12LMH
ATTv/H7qDsobB/WPqVo4hVxKllNIDzGapY9Od0FecDo8xFBjE4Sx8MmgO76ij3UP
NPs8fR2lQzXmVyYnEbAUUfjSMDzec7VeNOEJkS4hE2piHuSTMplFm+Fo9DgF/dGV
JXZNMkw5eyvQZNzwvluTFKKWrNhgvtrQSZkkpSZA6/YtRn4pPsjVQxTGJTKbooKZ
wNPSa0Kn6Bam33oI6k/MXCheOWKH+wSiEp6atQrASN2EVxzE67byifAaBE2UGDUK
mNNcS5pQHDIVhvRG1CvzvXURkIQzYTf9RQQUFWxTqMQrzOHb4Tfczegw+vGZ+MyU
hfvT02EhKvwNVOGgMsqXmyo2rXQIOKhvdINR/OwwRsBYcU0yfe8vH2zDBkTELDIW
nwP1k2CbUDe3cloWib6lh94DWQAR4IDED6AXMUSjtLj/4F+KfYB8lCylsMvlGe3q
st1vL/WFogV9JV0zPO657jjnADB5fy7yz9+s1jwU355MeWJR1xegc6jwkYTN1lKy
Pcc5xcm2FwbmRbtvMGi84cAoVqQ8n2PpP9xpvphTiQ4mVMPgSn+n18yFLgYWrsNz
OvAkW31QfQt1TOha5WrQU9b9HPzbaUTWDf9xerscK+FRcOqEmZ7zoUwOljp76Qk5
9rSkG28vMiyJGkF5rkrkygY4NorDfbcJ/uWaNeEq4Nb+p6pbrPIuP4UcC1+fA/5Q
GnR1tMMBUmh6rPiY4deTB4g8kOare3lbXFVsedykH/LSDrUc4ie4SexqgkP4WWzo
ikSAJOqjF7FLsimZ0nGu67dsH9VF26v/a5NBnPYpSAXsA+5KQi5ARGALsVFg1/Ji
cGqzi2HnEeWClB7si/FrjWcGgoJJjlep49Pj+aopfs8o8HkLSO19qOr7XGqDx2GH
XbMBBwJvOSogwPVzT8QWvTI2TUJX3+D+6iarpZKupRj9jFEp/e0+H/mm4xqlJGQd
Gob1goMbNnGmd6kQKq2We8TXwAPuTKxOKXO4ixG0hWCUgTA9JzW9vE5RFBHiiVXc
HxcbP+pvGoNqVp2tUQvDGq07RF3rv1tAUtEz9H6kT8xyVLXvrTcJgYG/cj9dAOHe
OeJigWkuLa6YzYU8JnqOGZy0lm8jrqOHzYz10Mno8RwY64Fu+Ap16tWbNB0oFjL9
A1hTDs7WH2QbxwjLAoAG5gWz5b+lvldq0jZo/m0Y3/F2GP6YwDD5K6TtRbRlnDTA
OR5gYqllWqHrHYsReuqPpjPuQAj1cgZfUTdEx2aayIrHuB+/GBdx0qQZ5YaIHao3
x38Mo7u14tnKbD5Ih7EhFQwzY9j0uWgeM+Y2Y6jRB5qzTpta+zHQ3v6knDne8uxl
MTBTN3D1r76uON6zFjyEY9DFQDz3LOqWPSCgg00UKQbuyCjToFN/FlrRe/s6de5x
7LS4dWSwfZ4tQxTb7CTgm73eX4e4+dCa90dtV9o4qqOPXZvkQbXziAl8hreAxXuB
QJyYF+zjLRvHkrG4C3WocbQnnaVPVHBn2Wahb05spbukPqq/4gGw28PjDZ7FGEpq
gJyiJcYhnIqGZeHpdKumITlgLJJL6NjW4ZJlZQlSVlZCxd8a9ukPn9jWNFxemLiY
OonDfpUEOpVD0xrPpkJQnp5qoPWSBqDig0I35rMk2+LBMQCFKug8R2hzl0IPbFXS
eud5T2TcjcZ6lrtSH39Vnw+2mKf0b+YRdVCDIHm8RBtg/1uI2eZWiFWiszFxClTI
bRMfH5FuPmqJ5IbQJ1GZpKF7IsFsL1KdJ3yJa6wuC8wSUslY9KS3k2ppcY2OB4/d
IFCmW+FtaGVYy6csNN7zBdkwzfqcUewNPyHZVOMelMNtfJKD2+XILuvZnLccFiWU
EmfldSFe3Al9H5KExm8bzCv/ogLgIpWCMwo6Y1bgDp73QsOa8ZUir3N9dJYmudPn
MVfbduT4IJGNLlSh9N6gfZlWDjY6ZLD8Fsg30iNJ7TK5NdXqS/d6IBYj7zeFtUgk
Z4QCkC5GwYDmqb+IDR6lmpEmyBUS8Cm5cHV37xZ6ZmXzWzOY/ggnsICUeGaVsnNt
530c+Oxh7e44+S0FhiYEWA/MprO86SLjzBia7sgekxa7f3Nyr8sg4JrKZ+CV1kLL
1oIo8e/n/0DxWKVYCUrm6KmRdHWTZiBYTZsDchqtGk7DbR+w91q+gxIOXYtyhe+P
GjZEVLLXimCudFd1D6jfcqjecS893CQH/4VOYKkL6RTuSdr+VdBzHFvSolWvP5Tc
Iv2UUAxmOxP66SJMd0prL2nBRrx0EcM9JDxr3e3+O0D77GjZCmtMPJ9tKsTp3nBu
7LkLMHLs6ZnMp+vcjIqhV/jP4NTsfuDRCgpZLf9LY0lz4lF2AzhxqNuQBrHZAiP1
CM+tCR1zimFpPjbegEMaYcnje5J6GDum0G8r0ugA7O2314gHIS+IrKfd/IaT1OGJ
CtiqvF3PpN9NVgej0WXFCsqm+RKgKmKLEF79mDihLbG5ETpzMJeI8FDR8FEIlJBx
LiHlq+B+6wtq32/kuTMP5CobI5dNwh4ezetqBaQ3BNvXi4hRMsnYKxd5P9GHWv+I
cE2Utqh/bSengJlNedtqtJ/273tMPGe10g1LkqpOeCqCwXkEqV4NN8na9FHXcGqZ
hKE5UtgAtXg29g7PNOMxgvJdZNoITO6lFzXkD+E9RKuEDolos8i0XKXBaGRTTYGg
MPOpi4bZC6dXPsUc1KubHiPlL/dw05sagCOfqBpR1cEEXqA7cA2eP4UKpXxdS7wa
HQurokgoypdGHSOOrX6MHgenGe3M/sFJZjkWkh82z8gqMfKFpClDLEb5CbyJcWbm
8N0muc/gudExvCRJBDkh0ImnmEW6W/JXfeHsOAsxXn9+gLyMrAm8e0EDqLxDUP+q
+Qxrs0nBDgfhO5G04vQJLo8cCBbzvHMH5+Sn5jWsacLHCchjws06041RWlblAZ1/
86hVs1lvQ2O0E/eLnVp8Dg+JIufDUnLiC/tCLAhGiYY86eLRY+gU0QtHVWP4jSlx
EWWHs8Qm3lraTDhezInSj6nHZQ+N9Dv44ihA9dnicsmiQjm1MYsba6W9Y25ye7ks
yg2kWdxvPz/ZyFNIxdUNASsaaRMHrkTnEEz8EDuHXSZZV6VjOZMFAhuI9Ek+tcAj
2lkg3lFuj717t6Hpmhk7u43L6MtOVcjS3ze/6dYoPCzD3a+4Rw7Odx7QD4ZXeSCZ
mfFUiSjJEhz/0rC7eZj0VyCSVFswPbH/Gdx6uRbU97p2RoqTBVvMh2XUEhAnDFx4
+Ou9hz/PIcBvHoYhFiuJAqbb0+5ZpicheEqQN/h4K/6Zh74dZT3E3G+zTIfVscSE
tfKSkUb1oIQTD0TY2TXGMSiH9Rm8kRpYhdXlIBj2+rNYhFGV/CypQwB5l3XLGOns
MvTCLjcWckc45XaBRTE7SdIwfodMzUfDRr/Uya2YwcBQYQJJeAtN3n74focEHTGg
JxQAEznoDmEsLaYM0baCrvU7/mwbIjub1LRALUbcYi1cCxu1G+SFMg1m+WmRkyl9
78DLsN+wYxyS/M2+EiKRX4izli+5bgLY2PPtqMEALYnFStJ4VFzwcuzIlxxst5ss
pmJwEuuk6gE2aqLFI9TbdGxaKaT6zCzge91+KjOCGjfE4PnTsapUgf+8hdgrlA2A
DZSrFLRbUjKbx8GHJD9M64fQPjvvKqnp/p7skKSxcyQy5xRael+dX/BnN8LPnyMN
DLUfj3dyjEPJ9K0PGk3gnCT3GR3ML+GcsjlRdde2TKrfSB1qUrD8PEwzYeYbxGim
D0+UXfmJ+VxDJ/hMPEMIKxS/buwM3LQIiWht0rLwEzF3N8XW4M0UEtmUpJr9BHOS
lYMbEZMpGKwNemmN10QT87SySy8tRDvskIF5xjN297AJiDpV2txY2yb3pi4DbmF6
7qaGjj0t9OUNJRVPxNDk5QnlBcdL1O2/oz8jfmqrl7g7RunhtEtXn4jQZg3q/sIB
JGU6g5UAEhPeO2l5gpr3X29xsLeOGhmnvZqxRvW8KNNx1klKAKzT5xj0p9gKuaeG
hvjx7Gx2gTddKgTKnOWPRx+rZWLwNzoXO3IcxU77ZsLcq9ZpX3NHFtU8NsL5L3WV
yZ18oty/o4lGb6zbmmTPFNch41dRJnz+hb7nQKFiFxOLcCPF9+/Tw4xSEpsJW1zk
mszAZohCcbburAibUxf8EWtb/9LGjgvZRXh9esBdfkR8Nh5jJiuTCXLI8KB0gKlE
NFMLsb4WzOmxGEFMj3a7KcmTs1iUIOMQnxEtPtXg7QNYC6kwDkJfzPbKZiew0wdp
ndYHwGL8P+3BEt4614baR7dIbNSEuqdd49VqGaG+whzKwa50aCrRhm3FqSbjzrUt
2V7be6ZYserBhkn6511xP4CJQFYk4UHAZDcIcuH9HgZComhS8DWCu1o4T11sQWjz
6nySpU0F/17VEnuB/o3t7odX9jIdJ7gqcYBoeP8ofKyQeY34feoU5Xu5MkOrLi/O
/R05chAYnRXnP8HAInTcDJrzE8DUo9JDxQ23R2ZplVBc/RPezKb+7X1COxAqLp2Y
Dh13RRyICPkiON9VSnZXsBQYX+UM44pnqE6wB9l99EClXw2j3edbKDR/VHHHCm51
18hjncz1KsAjqCvBe/GhMU+XYeh/YyAPzlDdMFxngEPdlN7mDamkrPSI1wSYbtGV
w41zTEnUzMi9ty3ai09lmiMagLek1du075yAtlP9q97FllxCfa1hcBEsOUJXfB26
nZSl7ytTtDkqRhtMynNHDOb4JfYx/ESkrfB5H5d0roJLj/4Vz4LZg8o69fKIOyTg
aJBrU9gzZcTBaPAPzd5dCrbeFyfW6VfvAUD6YCUx2AT/e7Q/i3eVoo/6R0WVsA8H
5XsSJ2zs7/ESwDC/Y8t1ubBskxM0iuxmEh445yNwU4nr0iSpRD1HoK8MeR/CEm9a
DBqwK+WBSsJwdtFKHH+M64LVGabss+wJ5OxcStJwUBMgizj4uazZSwq+iGecWHJb
VOtG8rlgL/YLAPWPSfATOCxnCSYMT1D7/Ihx87Ur9zIb+5F1OyVII8tNdHQbfNFK
gP4VJibPIHpJFNgUGacv8xxMvssVkOJZRyWlN4DVcJhW6S1xYYC542a0+CbiXzbZ
Spf+Ecgvok1wgb1meCJBZg2rAtMxNgZcvBxckVgRJ20+w9FWlB9FKvnsh9fr5TqE
jcgcqBJFQDtNcxHRqFv43u1cZcDaIdKKJt6DJ7mb2s8AytH4G9iCltthmcA58WlH
O2r9m8hcoNjc4hZGgMc0h+JYNwWL752lEIYsjF4PUSua/d1D+xDTXol7Rbep7qOf
o65Vi7YBiCnCN2LE7TKLfuYPTnxOdYZneikuL6ec11fIus+4VglNeaCag/cLV0ld
5EV7tykOSCz5aECIku5J92TFDSq7mxM8VHKY86l8mYXf/Ea1c9P01DkBLYh0MCkd
BDcGD1VToelh3GxuZ/x3MjC0aQMxtTEgldJGHhGh55NDobrUj4X/svfcBXlDpuv+
pEWB6WhVKPLP8SYY2uXvnrlKm11YLgwGTmgrfHW3BOCOMw1xn8Lwihs4B89B4hrm
E//KtEBmQBkHSzfUXGVIlhvUO+8plvLBfTjHIqIDjRvh/k1RwXAXIpFwq+L6654b
iv6NCzYtbuTDZoAKO7ktYmy3/Bo+9Fkp883Xtt26uyP0duxWiz5tEYQAM5SC/QVS
jT80a6jJPxwHtk+Qmp+8JF7HtdhabOSaIMqhP5cXNAqiMW/TknlDIdGENL8jby0L
XZr78nCcLUfKODTQvOwAjIpTOZVoYmuc1/02G7yoTjVJ0QGP15s5KKhhd1mIl+cG
Ee52V4G01+oilYkNx29qiQKNpYmpCEne3updw321xRlRE0N0GBp7PPrDiLYBx/11
MxREszoyjpCLtqkxCljpPFx1atSiWDvkU0BrrNkcsrooYk57ZSlB8Ve4dHfu1MzL
mmKzu6CkDzwiaxooD58unApH4i6lKS7j9zU90u+dTaZI+55OAA2OMOaX4/RMWNRo
b1TVwosvMCG7Q0lkQKoEFR5i//jTkiWHO0j5QaUWzEnzif97Xk4c5vCY5QhHXNRG
XIXHWMKtDPUyYQv9MtN3c8g1DCfSVooYs0hAczzF37OQT+l2jZ/wPqA61vFdSNdQ
76yKXOJquZ1V/ln83KhyeHMHMaBW9lIxy9n1+dKYRJg2+DX6SDEoVG9Ct/H6Jigl
8scj3nNpem2VR1xzeX/fOskfdXXz4VG0fBbgHSexMKoawt4bicre4Gl/E26/UmXT
OI9wERiI5MBJhsYSnTuqBQHniXW0AoDdiK90FHrU2oX6FWnFuLUsJE6SdSclQJpJ
Vk+00DKQDrGE2pk31COilGofZPkogK5B9qKo68994rDB5KXPxAG7kDsWBzwYL7st
D57aVUtIlV01OfSNhf1sWacvyQkXduHuzWiPPpRuA64T/CiAcrYJsAXd3TmCxQJO
F6SAH9Dg3wlavW36JvjPaKfDqb1ExoD3diwrCQW9PAtwcmq0zJYOc9uzJowvaJtv
ZP9+fPA3JmlBEzKrOuslNGvaD12J1hUWXfUAJ2L4j4ALcuudpmOU48E8lJeXoawK
FI5bWKKfp62zpW+OQmwL0COqq8GBclvgVr+toQXJ4jTRHSqywByeSHskPoaotsqv
YvcCxnY0DSP8NGGKMPxL8jMvYLYfAjHRs7JR37jgryvVl5M37il/t/udJmCalP2/
Y5orNe9JiTBsVmd3t5ofW8LcGyA3LrwQZXNqaSTKvILbQ9eTYE8vXADPJdcy2Xn1
4JGrjERqisUW0i1ly0PwKoWigNFBuyd7J0ISqc9aQ4p0M8RDHrqVVT6H6g8hMOs6
6vNiV+d5R/HvSqzJ/wEBZziEXiQg97gp5qL0cRdYgbski5rSnwbiVYNiVuDsB+YU
82K6zbxsG+5wwskEpidwqZuJc+/ruZyVZlIFBiyKikXqDSJvz0E1gO4G+NmkwDGv
ZyjmZ9oIegBlP2JIAKobD2bpLG8NfENa4465UlkreDcBr8/VTfNQzjM5CI/RXhSY
HRu7l8J4ho1LmlbjAyjYX3gB8e6zxvCE8ggprDbRURzFQKlIg08K97tq/naDARG4
x4/rQ3n+vpS+7qnmpasRwqAvRqzN9MGq9sqgeuL0PLbF0YtlRaEHvye5i2IjJvXd
DMlUwc/YOd7zURnlluJb1I9qYBkK2gvSnrA33+SlJJkME3fDcEW06sceZadXej7G
7Y5S02k9OyqdcClwA3zsGcXJgs2zVyldtXSoONPCQJxs91pr3v3wECbtz07B2tgk
OV1MkPngHnPx/CB5pDkaLPKSZdKuMMQ9mbmi79tbab89EMbnvNhKKODNNsDiWBTt
7tO/moClptsLLDn+hHD9jHB1883mnjPnr+64pBvjvDQKlf6t4K4EQLopABLI2Y5y
oiqvgHYe8YPJTbXzL4CB4ZT5DU6rqHqtgNWzZTPdeUgfNg4LtsWd6qV4flkh2agp
3d+WoPfvAAxM7xtgaX+TgAxHqAvtktUd722at6gxn+dZJ3mStJsVD65xLu+wqLa2
aTC3W5jSqfSG8uKHQXLHl0VlqmwMXVwKZt2vewUm5LnrzF/Evrm4lyinQuYrAclQ
IsFGFWPJCRJEZnas1f/oItdt+/YTSzR9CJLsuKbk2VVnpf/w7o+2M7dNtZX+vbeV
o0UcmqGXqU0HjBdpCcm1Ev6wuvJeXfCFqIxHplC/vXHtvegORsUnsw7poABoZdfV
o2fEZgDfafRiL7OxWse2s5pYsggGOtNa7SnoIEPoNPLGbAfwYsyeF2hi+5pMJitY
eEzrBcgcxE2FWZI8Emf5BRbH2s1sdZdIpD+Mc9FU/bKOufnj4pTMjdzivce6BW25
Oe2Ace4ZdxVYGlafjMK5K1TiNlRpZw0W52aHofvKxq8oOYTpRnIiwBWHaOzk1iuE
D3/f56QMZYh3+CCL99TOvnRC8w+NvtboVxUJhQWVIQ0KSIINCaARbyM4fuGzIIAK
KfhRfMXAdvRom5gpu53OKsQ0G3HW6pxCNwx9terNLJYzSuezCmBWBzweIzA4Vzts
V5cxpXcEe/nkuqvgwqMOkaPLv7YLJihskuRw87z2g9TwLfs0dz7pGqA6m0eksOcr
8buh24e4e4+q3ewtzxLYpcEfumY9BqdScarDmWEQZ/aObTznf9DzHpAuKC+Aq4/A
X0kYP63FYTk5iSu6MsVh4lbllZM1WR2BOueyNMn3XDYUnqezoW0Nht9YFTNQJkUU
b+5Hzh8RW3nmXTfva+7pCB6X3fZuJeX6GG+1HWAw+6amVu2ROoeN+WaMgD1R6s9a
8l5Sx4Zypt/Hi4d+FRPmt96Tk4bjpyNbBLoUtUbNhgl2rAV4VNymZ2YbeSd+eE2T
SpqS4Exzu/0OIMkiVMwE6riJXrBYPnqd+SkhRRX8ocJx/TvZtOa44ayMEWP2nFdZ
fl2E06y0ACaBrh0i/BgoRKwRC8NkLL+iaV24v0C2SmjNUp+7UI9VKHF7kAU2HcSH
8q9i+3zCcQEL6wPAglre6DiKCVhOfxxhLFLk7Hse+URTt7CYkmtDGIN5/dSsXAae
2jW+JOFAgd/naiVOBv3YjqWrH8mmHt3La4Rfj2Svp7X1UyFqpTk3z1rKyTj5hWtO
wewLd5wktYxP2c2RMy5H3goyjSWRsTt44fFdQ6BDyZpggjZXdNR9TUqd6km5ugjm
athJidzcldtJpC7WQvAP0dhbv7Pa8+scyu54stEVoy4GNgi3OmNH+/k58+Z0D5Wo
Ae/h01j0IEuJ1AiUShrblxC9oyZOo9cJR+IgceVktNkfpwK6A5GkENwpFCXh7zwM
elee4DGgjB355k2LQKxETTcW6gycOL4iBx5kQ5DkhdXHV/Un/MsIDy2T2eZw66rh
4ldnwdlYwvkLXy7sH+m6LgtuyhNXSrJCSPGziaIlZb4l6OdbeynxgOmeECOi1N37
QAz5DnixtyXQc8KXvdWwvmaQPOZv7W+WMagPDqstp7Nsd/3+ML0a7P8RvR4vgTMl
H9+4XlNRlWFJ5+9Me0wzd2YkjpfEK15PxrFRcyiZ3FSGThEbOGrqGuQW9lOgZN5l
lG2vZ4keAQWiwu5iAOGMHgAd9qDvtB/Uw+Hkyxu1kkVPC4h7xVvMkyoHVY1awGqg
SqZNlS9Lxit9YPr3zODI/1En7eUfNz7VcCtMLPzHl3UPEkBB+UJdDgTthDSJnLO9
Eo4w9vH7/hNn5DIVaGprJMvps5bUFiVkNq9Sh8WeNR4OFYqpG5JDAcnUQmo9Lv0g
Z5bnurWZGNy4waK5p6LK7aDKw5wnV5WYF4UmICtvsLrKRRuAznB6YZbOOUJeRMIn
97QWFWUwH+4vxGr+y5Ojac0XTof/VzfZZjbIHKCjLfHI405ITlgSCe37sJN3XfqO
jIjne2o9HJ7AKMrwrcOoeXmC6NAKqDYqEI1clF3kchNdJI9k1eyEPp1lMTgsRGnJ
/2FyIZZMPmEL+JRbYSkOr4411c085vHggdg6QsHDPxaCAD/wQm3mLeZ7xwUA/fRQ
tACFcxcf39AAgo0MzO4kHvPI5cDQHDy+KX474bSkIcuBt/viViA1m74wvHn7kwyL
9cUgBjfaz8WV6Lh0nOcV59jgohrUzGWv1XdDaVmfU+/SAZYs/+KdgbtK91H5wIik
Ug/rfhUqtp33Th4Ux5WmDFZwKKqD6KEHg4rzIffDwEqo1aNkdA6N+oR0LCiclt0I
FYwOSMu/nWdMlPZelIk66W9MRDdFJZs5mui5QIpuuh6X88QjMUrMPCNE3mCLBNxz
Hkw97K2tRaa5uEBTdRY/kUQtTDZ9OAygy/OpPjXYnLn0guKUNV1PN7FM7nWGNrxP
wm2UfBvtwBNIGpTRPOD8unKy02tn8CyJyv+K+Q7Jnc1U1VEjrPFto0edznV8L94J
78QaiuA88ie3SBMAYtMvdY9q2zwHoS4QRqwWo8iXqJpS5kebP9cv15xtfzAGfunV
FuH5EDN7eBSX85QFjULMTwmnmz4GualvjqySZqV8xKVNBoOBnIxP4XCcIFUUt68k
ocrCSy6Cdsin2plNtmW8eeqVnUtY7cIP2TF9r1KgY4BOPrDq9+Ryh0OWdGAoIvY/
gLMaEmvA5qSTFxf57l9EzfUtqdzVd20m6XjxcuYU2vEQ3eoA53z365j6i/KtOsPn
QTpSSXt88rvAsi+XIaTn65BPE8Gq4JmjNa9BsJNDCkT8O5x+dUJno2XQip92mlhc
3urHCuK28T9SYbKU9+uzvDglk7WWnhvKYaS6a7IV+X36KWDYMMnsmHqTqE9msnn9
uhBmOZoIB7Ue9yMr127nVzs7ceqGh6JtZ5aDzMxR3RGGFX/cJpRz18PKlkB/0Rje
nqCsjrKQtGMroCkTMcTSFs7VrLHOGAnRwrMkPDlpMv4KUyXK6n/tgOOcFZyeNFGC
PjEYBO3EWIS2EW3nr5PH7E1yYJovQiDbKlpGWWTrwybrqozU+gINc7O6NvzKR9kR
DLisZgsczMV9lhKM0C4OSiuIL5JI7UMEsNgglCfETICr3CxdjbNvwUMo0Ki3Vr5f
OqD8gCDZbIU4eO5t/4lak8iPRJDQmNgyN1/0aREETo6YcSqP808CKQkt7s7um0v4
UCrN1a1NRD8K6dl+T5UcTFTaGARjupa8yQuDVR+IFI5JteuU0ELLJ2c2DEqC4/R4
xFXOAr30lPdMU0YSLgeuhXNMs7irfUTIhXPYzzhABVIN4iVKBoSyVCKqEiNWlaFA
ZjQNWbWV/XvLmNd6J5BY/mtkUdpWLms1PqtRpbk26Bsa/MaOW69IkKqPysKqLh7v
2Kx7xRQgFP6QVgD6+gPXcQgKs0rjX5zeSJmpNIr9bTLaozM3kv9tQoZkSTah/evl
mKhWwSIBVjHbVL+Ut5Clb6D+DJwwz6xNJCRS8htUAKJMZGKaWB2ZzS54m1mFOfvx
sPx9olwsSmIlrSN0SRzA0OuN7GkY1g4FSR9nrDEuh6hhrHllrhRZv+gmY4h1Af19
gfKcEO90kAsryGR336f5B2fnNdPhoo+WEjpD48r6/CDw/eZ/tTyWDDD7L0gniJNC
dK1EEwuaROd24eBhIa2Lqrcu5cGDfUH5OukEScYKaoHAHSh0jBlK/6bBE7gBochM
OPktqxEy8rvo00xlzE0PnDti+0C/2pyhgDTBh+2tde/s1H3uOnit3UugHyrkMPfO
npwctn0LT7V8hDj2fmVrF6JxJIIz/fh7g6jMawPbKDzdzC/rPXljhG1ydjq4uZKy
WeSuEmFumQtc6WlRXL0NMPDDfoWKMRkMWrsCLDXqsq9t0lc3ukrIqhW636c5YSte
t71d4/JOpCMfNl2O4StLItwKjgNz9W6aC9B97OucaGq4mXi7uwnzkq5SSU3Eb42r
m/jDhiItjruABHLazCw3BrrAZzvZPZyKc08Bk05a/7bbXIyh2rEjJc0ZnFLSJTXx
7RSQ/CCOlHR3swju3B6rHH9a7Tszcp6EMGjbHuz5Im0uRcxEv2gG/q4LudxB5OS6
K7wcVzD6pJ2UxcYm84fa2Aue3E6rMXYWA0gKpSO824ha0DDzy5S6EKjB8qTdyMwv
0Bde3L9TJHp81hz2OaCXsqo3L9MHWr6ayxLaMHJvq3boGwORGhpfMX2HcrnijSdD
RQTont/L2DtKMYf14HVP6HpP+SKnYAOO6QT4vwq0zRLpEtXt3eXvvlsShtLVGHbY
dX0B8zjwc8bQiZqqJfnH67V+ZjnoFC+KzwZxeClhEPGMF8Rp6NfyqR0W5T12G0tA
dlDSrwrCUFueHgtIVLvUpkOVT+soiSEYRLVS8SszDeVF22hh8nuToX2+oa7gIvNm
94sB7OL+/1KOsW95VM3IrZ9k/cb1WLO5zg+9x1w3ZYA1y7LzaMOEgLKyx8YtT/iF
SW0Q93rsimRK7O3r7OGL5adMgGxvmFwfvFzyWsegQp/T3Fq8CSWNgyy9dCYpv/dR
h4+D/s29j/8lkDA8a+g5F6MY66EGCXysyMVCAU9ipKHNZrdvJ4xMX7KmHbEBh+QK
Fy0Wy2p4D+imAKRSrkCjT20jwQLtk1qhAa3QMDPpzvTrS3W22J0obOZpHqgTeW34
Fg0FM/wttZr8xRMLZukB6bX3cyJC1vGP+D3c9+mD/3rnMB+s7kCOakHDcUjzZTpz
XzTNi/GE6aowptKPS9JFl+hpxBBbtkU1YcUuGAE2qQwSGSeZ0h3FRleL8ej2N4qi
kaX+nDN6VIUaBMLn0u490YU6+/R1vpgUWsw+umyBnDILfzaz2V4MAWXv4V+iiLEB
KCc43XuNPWXwlsaHwKQ62pk/efzyDXlwZn0qFuJwIZEIyiOPShcBN4XMpfM48CaF
5wXzeQSKqs7px/6f3U5dJzdvUq6IvfE+tG2wU4HWdDN2sPU3wNeLbqz5MYTpFD++
fZSPr7dnWhZRZWjA+ushru69oIpJ0SRGslFE2QMaZjs8I+MTa+b5f2hllQzefl3i
Xd8PaRtqAXmwap+tpxW5oWVT1uq/R9iyWhQxGu6S8OrFgVQhEH/s5X9UcsopgE6F
WMORabPVTrL1PP6LvAPqlrlCc8uvMah/DDJk+Q+h5epI6XXyaa7CcfI8LAU0KdEN
Pki6P4ZoG8VLj31QqAqv8oNfSHIhfIBZUyALU2UxC1sj4KagwX0lHQQ4jWYKohds
dkyTDKbbfYB5R03pNI8VDeVbZv8Zi/GqioqW7/zJq46HhbWZBhKp8uPWL6dHxZFp
dUITt7OXzVGY4F5QYYT8D9az+Kn4yneXUphkGjwpy6N7ow4pESj1PRjBHTA0bKYb
UqeqV/CUCFpiUpFLxWNFZVhBy5/DW+VqFk+Svorcvo2h6TTigEAFOMjXI0TatHkX
R/Pl/IzNpvld9VGDJ+jRRC9PMzzniPG5EP+iS9m7sJ7SeOhlhxxztEJhvKvumepT
wnp/jM1eC+X47KRz6G4UaxrhU8TKmxHoo5L5e8iNbg21N4nHiLYWXfIftmu2mWaV
0TP6kLePb0dzsLgo4Q7jEzM4xSoedEyxWKIWn/ID3qXkSqNNWvrb8XQdJKUunWT7
xLZVf7DjUe49BIY2zrtMVdxscOiUAPPOyJIPxizjczG4jbhTpU3wQAXgJW27gLJi
HonwevRzhPl511DGQIQswNtfTA/o9jnkSd0l1JMPFhlqZqlPjtR2nikcMQZBz4WS
0LteHv6oQUSeHME17XSgRLmYEgUtkqpNYNBwcgikPLNjyiFNbxzLgq5eJSl+yZrZ
yZ0iIfgMgC8IoOqqkmFmNftOuwZ3JGRVhg5bn9oPa6Rqvz3Z7Hgbcg2RWlw02SFh
klP6xClC0sEBn+8NbHLqnbeWjPianS6KDskYGQUlQ2Q2794LdGX731KupKmt1WZ3
q0SuCovR+qDanPKWX9megoD5/HTyinbQ/+tNHAjcGighVpyZStRKi0mA0mVjbkO5
w+eIzx1Y10B3bhWj2+10Op8H7ZVl05URRGfbRyfOViQYULkSYIVaj3zTCswWvxqh
SqpCTecZje0apOytoClY9fdBp5nbD6O/lRRn7K8XkZpCqFf+z88CSaVx7p77cdl5
bMX/KYXJtX1Z+UOregBenRt3G5FPNti6d2w1gpMzDPylcxwppZvf4vVvV3ge7f4o
HK+yb55YBAQ9dd98qEFrOE3Xg/dP6mV9qQsE31hn/J1eOk1NkneQeiFj2KR3yqpE
2oAUHz2xpnod94QFO/pvYZGy9txBKBR4armo/u6vwTGDfkd/IJb3O1XhUcB6WuxZ
umgGkJGjRbSJN2jkDySbcZnyw9QLDKd35AiCoy37eO/YWpVwTg0BmckEbzeLugoI
ZQcv9G5uOIHiz5ySOacj3HT6btcUasLuUMtESS43lJGyv3nS86zvg8AxVKt1ieKs
3IF5rIcAHnMskRe1BvhMnYEqHZtrfeJ93wSEGPki2HJQiGtrQIQhmOzZZw8ve3yt
+BEMD+qgtqevtXd6g0dFUJ2wQlUrdP6tKUC77Z20pyDz+qmk4PuCJN4YEJukqsLC
uHsMuOKwqA3msMQ9azt0Dez+oqfEVLr4U8USR2jDA/Oqxo6jiVU2g9t3jPvq002R
TORYeQ9FWUULcX+2zT4qkKRzN7bypPk+fnqqMezogvvib+XoX/Ny/IP/OJH2srG7
I72N8RlegAcnCObZ0NjkkvN4gn7ztZMwoBVGfShK2u3mKWK83D/WtDmHPCNMCE3C
O7dyGrq5Uxluz0ojHyTL4WE3/jXFeNX79tshpyhEqeNFS3HeL7AEkADxSRjBZYOS
ocKjP8tSDg3FFNkXfxKHlzFCXcFZKCgC6iz/5JX1Aw33rx+LE6h8BVlF0bm/YzVj
Zeq2O8PcDGicPHh0b1Q//lS6hmvW8zQ3Ag/ECjPi8Q5fiMRX/ax+nxvYByQICRFG
brkObZYPxJvI5hRi768o9reA3FzmqApyKyv3nd5gZfDGJORrYKk1Y9uK6j9LLkkM
7NFIVgHotiOeUVIHh7yuxLOGBQs9dGjYceTPphOE2tfPyjz+P93d2irNI+qStoHv
+Mjh1AeeBPoXcoC31F4je+2D7KCN6UgtmUc5r0jhVYIuFzKs8Wl9XW9ka5JY4JUv
/9XAP2swvCdyuB+vOpQTi4dY1wgCIPGiCnfhnUPPJJS+OT0Ty5Wx60tfiJ6wmtt5
oCOYhYsYK/Z/oo/TvAbrKeNMwnqUruAVnGQjRIny6nPgBOQW42rTX6qnYKuGHAiP
5mecwD8+L3GlVIqzucAaP0CcR7KwyF/WZNhTQK89TtBYV7ZtmFYsHdWiYJiiMDRP
HmDo5r31jaUcnQf1RbemmKYlTxI+QjEoRADFLsUrAcfJRnJQGGLZ1+3R7Djo6vlW
Am5rJgma86VEBPAw660nbfft35zi2H1VbfFhfbBuTaOwOpvrJV0d+CtbQOZKjB5O
1L752chJ2NSwvYG/aLhIAgcaoM2/9XOFZ+ALkNlSHBFeSU0A0A17t6ozMzx9jQlo
1yQT9YTagMIBghLCwITGhuzRj2eJntKXqfSPZVgxtqAtG/Pc4P5Pw+bo8BgZFckz
mfcAGv2kk+dnPJirVjiflKOuCNah5USjR5Rv3PklFKhQ5cZUxg1+kHJLJFb7yKwE
EBdB8l1HTw147bNYfxPmbI14c3gAknhniJNqzftjzKTXlsmGjWoUkfXFoUPsGFWY
j1pdMga2KLaqmzM4XqxCD5kiX3HqH92ChG9Ii1oYHZiUfIiUNMEk5tElgF0ZA2Mo
hyVp9Xk7MdN885HT/BbgHRUiWputjXNv/uUrmrKTCiWa6wic3A9iuYLtMWt7lXFB
ZR6EAzuVRJbrQu0pB9dEpR1DwZ03ymV3wnsXf7E2J+MN7PHz9TnjDuCCg4PGjJzK
arzdB04pdKJMJOIozRuD4puQYP8thcXj8haMSSjIdgX+Y7//nqlX2ah2IKB9lfB6
+sQQy3UPMj/EG2mBKzaAPFe/aqLIc6LGjfzsPS5tn9v2eOP0lEdxUpR/QJnf2MUb
7VjAOG7bnfleH2avTynwesNmdpQn/NU5t7n9OQtJOR8Lf2/IFHw5Su5fo+ms+e1k
maDeuKr1vd6pIbLmqO3meAOHrww+c5EgchVn60bsPrK5kTLQKq/Wcw+LGR2we8HN
F1VU0p+0TG9y3LR632yz0X3PliD+ivcQnMmqos184po4JppsTCIQ5zQ/zJxHCEp6
0hUMtKkRmt+yvKTBacI3p2olGw7ZGJ2uQeCJKc0eh91kUfO42xJAAW9+aNHRpyCn
kCIBmvmbW+JJMoWy6lHnStr18PX6ounMxeWwSlCf8juM5ZEws0sMedTdjyWRouiu
pNjITtCWQ9jTKf+HOp88Aul/OnwwdpSRVRbYzYyXBaRN2k/PM2EK1zAtuv6+9evv
l31h2nLjt4wxh5ZD8527ZCC2+WSS4yhDtUI5t6rUQ/E25NUfkt/VYPiULWIoepkY
qd2cB1AG65JdZ8qFsarZ4iR0rXwTs7jTdQ3pkpd2GCl+kXplum24gmg9kKybSuS6
jGaj7G8kvbgxIQnukyGN9B9liOxR72CwlPABd8IrtppN2ebShcI+joYJcYkmO6rS
uoqVGXwk1M5Mx7wXE4ngEBuVhvzOYl3A1FdEOeZifF/4N5t0FC+XD7QfzfSkbgQ2
kXt/GEwcnI3+oVHhHnVF6DbYGHN+RhfD6DTsnwZe7ig+d1BmJZmaJKeV/aFZ9W/C
HIrRIpcaf4kFGKg8ZCdNK02EgcVC2FgtdwCpyLFotM/EazKbEJgSTyUCNeKGojNB
lPCikF8cTenUZrbPZkZ8uihQvAvfWA6drqSo+/UOnFa9HnKTAi231G3z3u07u+Vr
rnSmL//O0NbcDYbAl/KBuJGGXvvW2aVNsxOJ1fi/rD9r1E9gmxEhrvqcix3rAZDg
3MYFtrTEouFxM+qKSkwcMZJRclEOl29xA95eswUg39G9JKcABTs1uA2m63kReVh9
z+cuzTbLxULdtmJUZblYIOI7z6JgqRZLLo+fQdJGd+UQWsY1hURTgle04LT9bSt9
vZfUPArrjW3b7kEfAb57pWF56mxKCwJcVax8mUsH3tafWN0l+5Jm+aIIQ7e5a+Ko
V8Qb/AOm26t2thjGF4VH3D2U0hOUBPjWf3Y5I+EuZR1cWZAi20bX7Zfe18Rpz7zJ
vBpMrzV/0k4Y/PUpe8zluS40x7ZpX/Ni713KicWvLPlYvIvkdRE/8MzWIhd3rowh
xFy1g/9Mwi+yGDQN3GUwV675n4qR92xxY9ioGC9445RUjtMg7nvePp0aCUwA0CiU
BXtmQMGcYaVAXDaVUh2a2TtqzItEV5mly/UTIabOkThmmDmj1vbEDn0EVCIzrFTx
2jeTbhxnAO6Ux8neVZt1fIbEGSnx/C/qSsxvrhcqQpPGoPW+vhrpQO9ZnYK4E9br
iLI5srNjfycu+OygZJne5C6b4jc64Rr5/ExHcl//WqAumykG93LUF9Tx94fqOUOe
5ZdKIi1rYg1k8EfrDQJSwomlkH/MZhM4tO0Lzic3F1JI8vzkzSGydhs1yiDYf8y6
rQgVHX5FHwBZ0ysXuoHr8fSWAKGtTyZ4eIDbR9C/GJkp8UA3z5oej/45RYhbYqwu
Z9j0kWi1Qlr6D10T3mo5zWOU6lRFYpcUPCuuTYA1X6gyvWWp6OFodV27lpaNaTLR
SkYBv28QRJg87V3b0zF2fTTnHO5ZQEfds48tKcAHSkQBMMj2e6kbHyLnnG8YyisQ
GBhkPU5Qwp/QLyWeVFbB4/c6mI+CgRsvLlU2Xdeuo+ZzlJ1oeA/xSo1xVYayHTuj
zaRpM/A4dQK6H1HyJvCfE/0rI4TdyMoOMBwfLbK0NsJ60yBiGnkr9j4cZM6xg0rH
QqfhgZKzFoydpVC+hd7WhSoRt0Vq5lxnuhlwuFSHMoIpcKYoRJCgiOB59yuJ+swv
DiA+heOknaHdcMu6NSRv2mvDw8IxQWSMriU1a0wgnjlO1LaCo7jlwBn2RHrz5Zr5
+sRkIXEzEfIq5WAVkN0lRD7YPLuJOZLVRLU5GLTd8OBw9PW0xp5hO30osB5W3NL1
CJtK20plVTKP8ZaHj0FbD9EnxkBXwq5+MrmE+cMnaG5JUY0dyBSFN6sZQxymlM1B
F+i8hAXLA1mIyzbJLa/+s6WyDOO5b3wTbAJRh9y8LKJB6NutLvPjQ3msWjUkMRO7
tpEINRoTG21nlZ2xsUmFUVCenBgoI8L2M++NUxgkolM=
`protect END_PROTECTED
