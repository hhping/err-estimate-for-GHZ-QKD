`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V6eJUAteRCBdfC2MTEb0suNLamCXPg0T/lNLxK/Qm6hpaBZ1M+nQBWEc/FnOV/cJ
Yuh9sPAYCGCEYKuQb5AqC+Xmt+I6n9g0hIo2YBTGa/9Jzp9e6Mnq+5Y0hax2ZRlD
d8+msQ1lnyphgLa83jVCZZ1P8ewnMiESY945besO9ULVrpNzeLK+s8xAnhqllTbP
QCo3iefXHuVxiYSENyCPSGCzEUouzffZuRdJTzBbkhrmP414yXwwQVedKwlUDB7m
s7kKMGNa7LVs3ILUMAUbAaebof0ps6NJbflDSZ95jRDa2tANBEDm5ozF5VG3FrC2
9qLju1ADaxrydWcv/Fes5JOFPcHeBGQQ6sIhmg+3fhmDYSpoLBvVLzXhjpe+FcuS
mFFvYFjZCLjzFTZR7pJHjzCMnLIM9JMzKkRdG2A4XfPNLNXLUAGzKDX6IOchGrXj
Rgcfuc8pHRrrK74FBtjah07pWEY5IOyAluPLHrVrP1bYQdPKlU/bGMlLjpb1boej
`protect END_PROTECTED
