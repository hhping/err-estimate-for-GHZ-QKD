`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bBdZrfcNxbTAf6K8kL7adZ7wH9/yKZyCqU125bWhZmuMJNxz09s67CEmYAXM1u8z
l5/HaQhtAuMo9QknpTX1Bi5lBLhG1ra5NNHwTJKKF47ltTK0de+6MyhYVG31Q/or
CZfFCN9Q6Qs6OsLnzcZ7bCZUbQ7DeEpY65nGDl6D0lKxH2IDWUQDqdv+v8ghpQXp
W0brcQjxMqFCrfge7Ws/7j+EUX6mbyutAnSkyTWUEpccMwb8Fa9y4mfEmIWLyPLS
Ew2c/QsaSH9BaolczuYzafe6PGkuTLRC6JCqFwYhnDtm5yR8a1Dr8PnA/NVHWIiK
g9VA+6234A+52k2T84TPdhhh9FWEoO34sJOg3rF03KiUMyzl2Y0HCM5gxl/n7Rtb
`protect END_PROTECTED
