`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MPPBcirEkIzWs16IYmmqC9YaozrMOcbTS1zAtnJWwpJ73WizdSHuS33dN8bQd6gs
KVJRGgwiVLXsw3f12QC6ES0FuwbYITpitpzN/B19+w4BPySoB44C7MwD+a76VWXZ
3R/kz6DMCdlqqSe6x80lawOjLoMPtJrL3CRyFXsRXwCPyjCKQIcrtDj2j01QYPlz
pVTUbGVucxdn+R2cIDDKGsJIqDuDCNfFgtrfbnnjGi7+SsGOYSffBoD0HWuNK/4l
mp07xrt2fePhNUqirPhwf8d41ar5cnWftnJHR0jpHpRnaFOS4RH+NTSy14yUQvSP
fbUTkINX/n1yB1nTLV0xJWluUG3IeOjfE0A4Vn/2EfhIZj8ewtMu6UtUIA6WYZn+
WlyuwWlIVLgYpnFqh/YEO4REk0fIV/3Lv0FqT/ebQ92EahDhiC66RMUsnVAoPWYl
FXqdx6Wr/9oTTHgeKK8yv36yoUt4ncEssoEw9fohC2GXKdkSja5mzJXTX+hBRhSO
i4K96+jMYCFSabvXAGYmbmTUGiu/t5jHgkyq0tqQqL3KVOMdSkVzhK/7ZQ5CDjMT
9zne0w7qYptS2U91jXIR1qcU8IS2VZDKeCfsU5qJUTrlPnljNkGbP1bPocIwvRtG
z7ITN8TlUQYWk/jXy1+/RG3H+Yj+jp6VzqQOOueH+TVKN8ap21XdIeb3s3UcaXKJ
g5n/8bB8+tIu7+rlmjPV/xO+LEMTLJMeTHUN9orQgiR2CADSTVO3kqgnE7FZ+Zvg
0Ysst/jvk5GtUlJCsGH12ym9xR7fSI7i8iHLwiZHIjA0ycgLSM1KbMy4i75x0A9a
HV2f9o4BlemteBNbMfKfwFpRvTt/COKNemhwEW6zJ4IJyGkhs8Dxuu4m0QBC1FIh
KfZHvz2byMcOjD073alGAV4+ZUrPI9zdAaYcstzH65xUM9RKVyAVbdH8fzEH9P6X
Xs/GcOQNoVNfd2DJLST8qawYXu9TMKqebuvdhXd9nHBUf/6PySl8kUGSmjL6PTE8
Mt7WRlSEVJL6dXbavcAweStYPmMolI2NFLDbqV+dkz4bosRdfkYbFMhbye/uOXNK
IneB60rFBkjHM20ugM1wwkfz49xYIVK7G9QcMZHo6/B912xLH3H2sC/JGYWl3MB7
O+vtALqdEh2kvFKHxZ99bN6PKjF/CJYSmxd07RWtQUpisyTqkq29N0nbdx0GAJvZ
+lbP+97X1s/gEd2asLMODzNtfz/w50m8RGAn3kDDVNrWOxzmLEgg7ow6pf9W/pl4
`protect END_PROTECTED
