`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KIxQGstSlVOqaCGsctbXf3Nr84KCcyjhJZ8WJcZXIDDK2EnAPSuNNG1ijuyL8w7P
mJJGaaWkYJUXKsw5BHgZAJXyNaJAA24CWLGXmoM0gFxZrsYasm0994cm0ihih6ZR
VaLvQbE3OQGsEUaj7m2SXvbU0lP/9TUvKKxibm2sMSqYZDlGe26AdY9xyf7LIkkc
P/o44ht4xuHjFaEe1t7GBoFQi42sS80xiqgRlCGU0UKvalmWCsq0CUp9yyahps4E
fxHuSXJ4MPMbKf5VFb7L669HLuoNEChWdWzSr5XgHiA/cBseQCISYH9xkop9TUML
VeDBvyYt2cykOrrk8qy4YuBycRVQzjYoGRVPIhce+gemACzGDrBn7fzocyCMDnrV
PoL4GBUDFkq1vH0S7B5AxonlTKT7GLYtWLFaOCe0YoHKoP+fPXjAoS1FNKdI3CvV
2s3cw0QJZHP5goBRe1WhYU2WX9/UAtF6X6iWPjbqxYD7jQD4lFPkFNIdXNYSinI/
+TG9V8zqwhFm6UbI9Ogx1sV6LzsjRvp5CXh187oxljdaFQfJJ86yqYUnsX2ImkqT
wTewxi84VyMMfo18rO1EE97VTlw3ggTo+6P5ZZ2PBVFaab5+38zzyqOE8G9ahEx1
O+L3o7gjixS3RlWXyee0emnZGY2ybsE02bt3OMwpzNRYecVnl4MQBRrjv/yXz2WV
tVByIo9ZkGAMQ6yYgbIiJw==
`protect END_PROTECTED
