`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GBTLr6PbtQLPfrxLm70u7V7a4cC2kI2CeqJwY2fbSCrrWlkbJiZpdKQ0Rf2Zqm5f
gkuf34w44d8NNujQd0piFElIhgN9x+3pXHJGwbKuvK/MYQ+I3xq/C1aS93ZS5f+v
ICesx7gHL7XBWCUhUKSilPW0XFdAFYBLhymUc6+X27YC09dp0s114q9Obow/KA3E
h56y13TfH17UoN2KYjsvo+ebjRPw8zgRD6obJxsLKYzUTEEeC2l+9bUMJlTp620C
J7y2QYfJLg/asSc20RfS3xVyrpctefdSArgXH+hMARmwCjMnftMATtScoBYMIJlx
bQEI8b9A24DP6CGjaLwgUoyMDEJXMxzMamngIc9Gwx20nUYPJVuH/3JCX2pc68b8
9KsgyS2zWWoMYqrwrETKRtc4NGhxStJuZBDCbACexFBcvVWWKW71QFLRysafC0Rk
ThpB0208WF3I+0JGH+au624b6uU81oSCBEzt4hJhVB32Mu84ar+swaH5japuZPYo
siJV1nOZraCstkEFG4gNCq/YhoqFS3VSddD/XLnecKbGmvH5jzY9zCxsdY3baHc8
Taw/IB7WBIrXePYZBWbi+RIWHKZheTTJhXBGr9J3aUYBxzuLos4qfh7yuceXODRU
cwg1LP3AQYzJuRBbessXo/bNJr6usIHbOEcTFU6f/lwDIqyGNAthgETXyI4Y93oR
zi1A0Zpar2Bo/lpU8ZWwbbSQSElWZS5rkJSdwKZZcjws3pYVbXGexLfGHBbGv2OS
In8OnG+dYrpb4PCQsv51svMIpUHLFbhw0xirfPSAmsrn4vB0OuXnE57a+rVCHkwD
FKiH2P3ivwr5crsM7DrOKWb/77+L8SJxHrB5HYrN/SCWq1AAP9PGj5h2nXy22W8Z
AHx9tkoGz168uwUjtFHPUBdv9xcv9QY2ZM+eYYFQWtJCvoUNKk7f2guZ70z7diWP
hGwhzo9FKMGTgKkEiIrqIg1Kiv07D74n/26I2uLepY0=
`protect END_PROTECTED
