`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G5yOZ6QTmitww9Aov1utoGAMy2Il8SGPQ/ritdjcNIxOTY2t/ScCi+Uo+L/d4mMe
dPD1ZczfIkIEKMjcS65wCRyabyczEumghK790xGqMdRq2ptS/yqHkwSOtBCwLR8z
GAnz1xbYC8XPgsX5euioe6WfQFyLtfaJTz1zWtaRd74oiROX43oUBHhUBg47ey40
WPh0tPLpW3KmsgnvvExRozXFN/q/zeKyHlV7HXM7Lw6n5BtWn/iZKBeoaPr3oSVw
PHZ7PBUl27Lyeil2hU2gQmpVKaRZqC8olel43afLHtPvImo9pG6yEe/ZRhzFaseE
5pu0sM4bHqC7PKDhI358ktRcW5KS8ToOnpvv4jiAnsDoL9iBnAEaPgfSd6HCAUKc
Xkc4ZPHP2m8E//LwKsnl/0SEJFQJfPu8DWGIAh8cvhCciBw/bef42dWY4UR5F+b5
/a09xxZL4P0w/fSbKu20KS1xzXbpU+2crqkDkAFo9TsKd34sZJI1hYVQYVbn0Bal
`protect END_PROTECTED
