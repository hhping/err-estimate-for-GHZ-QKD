`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JVJmsEt2eOKdyqClXDkQ7EXEk4D2HyTg5EUxuWcQopcNOfwKNgxLvf6GwpFWYUTq
82gHu2BZIKdUqYneKEzeDHy3tC6UVddntVD3Wg3IVhpoG04HyZBtiNVlrEy2vb5j
6YOxRRLDZvZxa1ixQIF4UYVUmSZs/BgFvtiMU6YkdQhA0SFDu8PjeWiIDkhKvtbr
pmpDanWJJE1dLknw2WIT4bnVA7Xpoj2V7p1C0BPklsLIoFEIPcJNxSZsWkwxHIfn
fXeLjsRcl7MF3gXOyzaZWzTgOLH2yYY/ynLuH77HHSbgSLj9f3zaHfRgukIK6EFc
yYbIo22JHtSlFWcepT8o85UCWOCGygHEpKYmW5bnXpu4CkYudNpx3QnzBIoDNYyK
84Pg8SF1DDyEn9lTIr+xAS26kEyuBeAN84bTBcTpRGU7HFuE1z/h8KPs886KLbgZ
i7Qh5b5CbiqShAZ1e9swcoKfxxQ0xb54Qo1PQgetITDsyBFGzywP1ZV0R4h4VYnF
YWeBRbqjcuYk0sInZi/Rn6eMSgJEfdHbW8qpSovPQ5c12MKHoIg3XFlSyi4BrXex
9wdApq1zsGLF6JhtnXZPGtRZe7iMHLrEdxb0svDM4llNyrRe6j6rAjwZk7Xp4xrv
oGcU8aJb8D1LejuBukETQmnFvzyohB5mWvUWG5tB0PbNNnLiskgHa8qX4pWFo7IA
3/QhrDb7KMvItQIzdO+4ZstZcHNRy4bixf3yE1VzaIIs6zsgoscWhlgpadC8tId/
SpzSCynA+i25yajs6LcjbisaFMmaENR4j+sZyXysb6IgN5wagI6vLEtCk67J47MP
5nejL5TDJ4Cw4qaA0QiN2oKDFwVzZyjJf/z8j8TZf0m1bGaTnQda5HtfLo3+dDYf
3Y42NUJnGDsYvuyxxM58meBb3vFBvLt8KUQouega/HJ2aau3Ndo6rtz018wRutX+
pgLDESA2MCHZq3epsKzQBT9tgZMlEVqEFo6sG6fRCiMMnHSaI+eYav8B/4Y0wZdM
8jKq7ay8ZAps+r1kAx1jTrhKaP6H+E4zq5iXQw7rAh1mirOF33eZoj0JNIWScs7f
BVnrBQDQTm+FZMCTKqD3Wc9eWDxkiZGHzEnE+ixJn42+04v8crnYqGi6vRziRXrV
YOmQ7deBa7DevnLbGiTzAoksLXZL5sjphLHeOgfrdc8qR3wYzYC2l+Taohfm9lQ1
mmxzNfUAtocnMbm+gca9UkGm12dTSveK7u3HvNl7OeTVFw79rb+bwOP23aS9klNp
hC84R2e9ihHluIZc+kins/sFCztxXjQ75REL/Or+usuWm7rZ+j9c2UVQE2AarTRX
Rhp9BuD8yEjtDmFsaOJ5PI+1bRekH78beHwcIdAeHhl3HxWCDJTTVByl21VLhsLp
cfe+bVAS1CYdr7kZ3TunJu26PgkdSZ9bNly1vBRmDwZpeewULMKSWKAEj1rAT+Cy
nE9Olm9OfILDb6EAibYQUkrIZR1eJBgWIJbWB5L8XlL/6ISW20+irK4qGrXOP9el
ShBsvpfnQPActX+F6ekgvm6T0L83SwDTqqTE/ZpsgzN5xxs6Fkb39srZcCILDU1S
bfh5t8d06VC9sU5PS3CXYjXp5y/ls6XORLoRzRP21BziJINH7OfjI1oihtTNmrb+
RcdOFrH2ZHbTlUafxRetId4cCl3ESqmtKK9soq0U8C57cXLTC/DbbZPxmLlGJkpK
8zkHqx6STt3RWdqGxsr508hvY0Rn1eVRLXtctrltQmKp+coSE9wPr80EVJ8xjOyF
8odi9y1IJJfPRxCa3SwYnxJb9ByRpuqBN87qKs86EfIvPqNJRz+Gnd9md1r5H+Si
DPyOi+o3RC72ZUWUTAzyOhUF3tsqq9niUybOxcsC8PfmzbqlZNpI+ygNmPIAh8Oy
vWDKNol0akOZU3l/eBy/jgEBKxHfZGp1rsP+BtT6KuDoSbLEEsIJHaTFrupIB2ff
VnUwsZf42x9RmIfV2aVpaZDTtSUoYL2iyZfD5wk6gpYHeKmvGT1NOgV2crv6fy30
/4NpXuImYpTAkRxrcyottf6ahQg1SgL91jPXm6m9Zsy3jX/nsQcbVZWHwRXCdXIn
tAKRqJ4ZBPXmNAW7B7h1Kubg0kmU6qudiLqyMoBtAqQdN9unNmIC2XqWHYL/SjmO
hZM7nm4KMcUhRFaNykplltJhtEa47yS0CJNi5rcA/yBj/a2i267nCFgFLEgbkpMq
ycBa7PxN1WYTLhljWcx3PYJcOy11LzCWYIPj/d9+x1nW/s8vCxswZ+zT2n+pTpMW
i8tBuIH9WaoyC2TZMzh3IHzyqG5n+V5dARtQh7bRrtRJQrzY21uoYoPsyBk3wp9Y
tjTir+IKPbDjQPDguw99BEdBWlSrmgjgpOj5wk5k/mhgjdagAFOpZ42J9AjnUQJi
homx7EcGqZvu/ZwXY7MNogVmQJ8rcbnzKUdScEZwi+W8l+WJXy2eOwLRj08gTHHz
9XLt/rquxHUj0uVuYFQ1I58M9T4Bg2XhWKDagsscDVjxGpiKkm1iEMRr/790Puju
bM3qwVK4ckp95h6ldLVzQnEe4zjOPdr70Q9MDhePjjQ0STWFZYFtBao/4yegZ3oF
iFfJ6vw5lVAxlaB3WcKsetpQs1kKO7xGIux5csQNBAfCLxFgE4m/uVI2QOpUV8uS
hzQ7Pmp2t5LiGJg6cTT/BSqynLMy9gwHF12/rC/5F9PNLsH022vJ9jm/0pMFiWT7
rU9gpNh3rmFI02PZ+EWzsp5JMcIVIJbxMcKyxPumUktFLeW93qZgQ3WaetJsFqk6
LZ1yHH8YlmtPLauAnezXMcqB7FN6CSrnzoPyRmmVQYHzk7BM/BMi1DT0IMstKJw5
7NgPCxKhOIkoBDrme/lp/rV+ZVFtPslUL5IuMAEx0p5i0V3juAg/YHjOqfqPv91x
q+/nRYrBtHqXVUAuoT46H3zTc25N57/bYWJ8ZhFNf6Co/Hs4i9Uco285KKtBcdYw
EnxTtX+vnzGgTH24l25Lm/fCnNnjAR907MP2zE6nWk5D0GYUnVVz19ihGvlLazHR
z+QBo8g8Oa8TCHxXHlBB81f9KM8HwzRt+yzGXRo8yAEmc4mCXu9ZwupGkjyI8xIb
KQY0iykuosENYHtQGCPPjDHOq+N1qw/E/t4Gepp7gvZX/zQFq3Gru3jUliDnozIS
w1szxo/iNBRmfFQEOfnzryBirRjcruMj9lbF9ERbYg8Exoqz0MXrLKP0ewSUMCrA
XN5yn2fk1rzoaCC1TPB1e4/dpxpU2fDdfWWD8VKEgdVhd1UcOS/Ija+eph05piwr
OG6SRnLEqwPHlkPhFQU9X7Nt6xJ39DaV8kZURQ6gI0QgW4OX5dc146hjE9PM6ktJ
VzMTav95UkyuMU+3G3I0wWfWtOVBKdQl3nKF6lTkyrK3H3r8TAYFugFVH3KF5I/X
jIAKP37qteo0TsRbfd+WPtEVzH9kzKFYm/f2kZ9UAuXywo8MBRNDK34zAWFgSKsA
iuHZdPKY0DzSWVr8nTrq+yi0nANrDNm4QgVvM+9Z4aVym0iPpYxcQLCxinOpno/w
mGh+/MK/xeVpNash/AN+xrvoUDethq1GMwvgoYlyq1iXeFXLAYYsm7R1F7k/Zjhi
xjMUS0BcrEWwheew42ZAiUtWS6WhWNJV0t7m9OI4zTlIWg1R9O8+TkaDrcgru/Sj
MIS4xHGcPQR01+zhlBvacc1Fwf4Bp5fJwT4mRe9bccSPuZukJk9GJGTOPwrVgylc
deGQ7HcEJvqHUQymVK9ToaszDn9dgoK57wEaNnDxdLPMH+hNi7a/8qQOCn/sUHW2
y7FbZWRYUazGGwQugl5SXZxYKl13xUd+VCpZNFFm+FHQWcHRYwFRpejMwwCF2Yxh
f51B7nvV8SIVi4fWzq1JB6RTi46k6VFO9Webx7xSCrOypzJ/WchzcCxkCLyXUhMv
B80BlrkM5/Q71kwQB0BsonAN9i2QJeHnEFlr7OI2pAkwF25gtBnymLUqxBzdntXO
ssOiBK54lNrYlghF3N/mkrn6xxJrm9+GwdHENsMINhQPPV6bYEV5KyowfM7ATWwq
hI50C6K6Kfw+byM5MawWYvJfS83liB9b1THuZ3mvKPCjS7h27hyaEgRcL9T8Q2pv
jtHbQzeCs5zMgZqVhjzeyWq9u/aqRkp+hjbjXF3oJ+RMaZz7WQTx/yw7wTumzCWg
43f/ITTNc/c+5dAAhuolD/XiJSQ7fJdYp7r3DmGynK6+RPnLcW7Gcp/VN0t8sj1F
`protect END_PROTECTED
