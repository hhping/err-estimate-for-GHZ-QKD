`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ytgpSI2NiA0g2AP5F+PhdY8zUXhIqpKrkstIn915ZVrPx5qumT31d0KMrqesMnvr
7sQLt4KQOmQOHhoa+/Ytmg5b+6ccrlP0nCJ3xghYtoUa09AZHNcShn2/1uzHGcWy
oXQHYxmQSwrUTJamSxnhgFY9LjTLQ2urbxSdL3v5G8cb+JFDMIzGrsmsWKLlgftz
CHcm5vqeMwXqu9gYp1Cfue1wkwG/JIFnU5wDcS23o+yTtb3HQ81NEAkKhAoCZX0S
/41mEKhy4UFAlC8eTtgaNgMB1hNup2XD45jaoC+1yA8N+GlVq79K1yJDmzCt/6c4
LdefmZxh4FT/uVrHTRF3borFcIjVUKW+hb8p0cXWZT+6kDYWci3huEQQPuHHDg3b
nGnVxiqbIdKHky1dpNdNRAhid0/xLefaeVSZIiLZFz1PKzz1TwYqVw4YXd8HXMkC
A09jzHIIlgry4fX56nkbCOPXNRxSZAgR28BqvIwtBwHB9LQT82e9wvOB/3g+v97P
3QnDfy9RKvhiytwuLxYgOoBXgK9OCm/L/H3C4NM/5YGi/4nPuLugno6IPVUTwBaf
bRBf5snQzziOWnvDggWRq94yv+e+n65v927u3kDeCPi2XGF26Qwlb2u6pcGjsGTM
fjAtAhe5uApkR+Th5B/8M5jcxDkIBRkE9oVcP5c1g3Qw644X3FAqe8pEOOL3/1oK
NJk4yKt7c7BJ/vObkNsRDYrkbUk3Mc3GIs+FEYquLDovx1TBaNfUFYhKGwBgvJWa
TCSihcdRTqLMHhDhy3LbjHhgVY1aEJjx2bQrmzoPndPrTx7rqCzv/4uZxg5akZXR
8Pmkw+GQeXH8tBI+wQDBj4CeLTKYuahlljnlWK4DiOJDgFEk3Y8SlGMPmhNRzqlJ
rkCzhrmjqer4EJaeAKkfzzi6N1Lobam1ume9DvUIGLvZTQR+Y61ZboMkC7qEg7u3
DUSHQIizm3zfNan7iP0oih64Jf3Pm+ntijKw2DQr4wkSJ/Fe4Rvkocs50hhj78wu
Lz5eOJCxBK/7pQxbwdSkbp/Jz3rtDc5pK/cHMV3PPC6wdxp0Swtf4/FywSBlvzl0
I0mWGnJFMeSkkSY8PJM1MXDVj4adj3cALXOZn+qmrkWe47xn8Y+HkUjj683ZTS7Z
sFKgNTU8T7bj2QhyyNiAiCXZKpX+Ogt4sfo5WZKQzMJevhFQOzv6ZAjY83kszBUS
HLB+5cDmkxquL2YFoyvsoe2hnl/+rFG5umdQApSrzLrxY9ZmHAx4crb2XCpKViPR
tBVYk4it84ZHVoSz+yu5Eidq2U2BQCYMEga59qhLN4BybopZ/6iOJzVswML4rct3
lujnn1Y37pUMENocx983/IyPTuAHqljOzjzdn/jl/66/lWdEb7fBx9oDiZH00dlO
apYjDW9c//gP3pZY44OTKq3QrKK3tY8+ahqkB3jwynVXl0/mvf5osGG24Pu3T2ii
nrw7PwaTYGhw2hiSxhR35qZne28YJejB6J607Qe5olJxoK3iwY1zNKCZ3jmpwbLE
Vu6pmpyNt1CloJxKR0jmkaTpocQg33LBc7m3DlrMQkNvZxJPFX6FiSKH/MSx8ZXz
67XFRjOcW5owmTQZnmzvuBZ/vJnKxtFIEBd8RyYorFYvxnv1953CJ6YmQMny+erz
VKwoHSq/n8AY5hi3Z2K90IHjC9FvXgkAN/rf0JAyH5xLj0Bz2X7unPHY9OJU43oX
npwG8I3P5sdvtlZjKwRmN4+YoaKqrzFnlyz2boeIHu5txY+KPZsih8Qr/1TgTMyR
aCabKwrqGVPDjMg1vGdvKylCsyEKhYxy1ZLHhHtxuL+BG63w0MM+zROSUFjP1fHg
MeJ79wumiXst5qxw/Og2XggabuN2ZYQZWQHlykToW9JhEeXDRw2A0/gDGa4QCswj
/8MXo0OZCoecQPYZ2WqPB8/aeBb2eVkfgSR3TozbsKYDa8H/gLf9kF6v7tfPKU1i
ow4PnC91L+uSIWux01Jlo9wO+Bom4yXYXUmVQ8+RDeHSjllNvOGWUrP+xNX3/gS0
a7FXzi1+phSYG7JGKUVKbbPX6cgbndTPfnoK/SoWvmURjFL1OM4O7k71D8KoU6/9
jT9jhZI6Xurhd7J8SvmcClehwXd/QPNfGPdl57TJY7QGo7J+yMF66LtutciVN9ux
NNbBJeGou70igbhjFygA5lBFxOa6DXeTf4+eWPeNnc2nwMEWMrHSjTKjhwXVLlDc
LPcwUwLXSKirBwE0S+FJ3Sm5WfIJCojd715mRBSwQNX4y+O4cRN6fAKQyDrmDrJ1
vToJNq9sKHBAtY4IugBnoPHD0Dg9HOWe09f/9uK3NAaQ7DYRNKk6zuOciupbOz7a
LEwR2u0DemkQtY01wRq45KXTVjzXTra1v9sebJvcJwfZgEessx9SB67AoLHrtg/D
JVU2Fuf6qnsvDH23dO+nTmubkueUcGfW4LwQ+QN7OYKatlZ9FPJqJd5lhyIp22EU
4DUWWzDH0JhUgt7DzxQaJCmhZTe2YaEwpTrrO8erEHPuidAwWIa+tjVaYSVR+l0H
X6h0GFDGqcg0a2WgyunZX1PKb5MdnQRuG/CYhyqufwcpqCOKgWxECMTBMBLqzAjB
QGViSb3Zbdive/GOW85DUROnm3+py6zc35vARilMY7pTiLhmZ3lZzypUPl7B1X9J
QLmYkSh78qzftZ1zU6fVAHXaM4CnJzPST6kwvJeWVbELLdfsNVgVF/m6Bg5YZRe6
PjjzdPIaBpib3pBAvy0Wj1PeI/qbAeTiuMhTfLC1B5ntsLxJ+EXhEbjU6VJedmaC
`protect END_PROTECTED
