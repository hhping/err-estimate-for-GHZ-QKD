`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jehxjggFfaThKk9owVKWo11tOo/PjSxrAONXmYHqs/xUsKlh12J+4CUG7tLbGk8p
Nu1qMhFf61vNdga3f/TYp7A0T1X4H1RTHSzALlYvhTnjGStzKRn1azOh+5FJ1ibu
bvXoYN6vEKxyRhAqtp2lq4bIdVmA9SUNQBLr77nq2Ee/rMvta2utCOJiRfOvKs1b
GwtssiFLaG8o3ixko0Fb2ooQzYlhWY/k6hSGezBdVkwCZfZzNN4CZ3yGSfIGlNwD
QUk2LVAI3yTxhP1moS/Z2zwjgpvEA8CNpx2cT6juMvUlumFv52qvb+5hbUBH9wKK
ltoZl/qib4uhIHXch7Dz3J9cbhPuoepOzuGg8Ai+6ytJlgvQqQpf9fjajocgvGT8
j95B/pKi7kP7xQ2wV1JvTA==
`protect END_PROTECTED
