`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D2fOV42ZiMAwxVfTze+aupyQOEq5XbVExt8lgID1nSJXSZOSjX+PM9YqG8H2jNNZ
k+SwE3/BrJ/aOKdEM9HIQ4fzRek2yrWEMNffaIXFkQljf74a8vdp/3kIbV9Vs4tg
TkGaakEGNA1tVTdZ/eMqayFmapnJpXPH0TfiW5zMhkSyXpNTRExCLhgv+7XNIx24
CgrrsKNPSQAwIgKZ1CoK3i3oEV1NmMWkjiXcI70cQqncixs+bL1Kh5tYEWWV0NYw
/3nl9Xn5G8vQ6zD/a1uQOq/V9EpuyZ3tPQR8bMWGR5H8dRZxnubQwzc04GlkXJun
133gCImla3ISeLNU+Qkhq4xUu6LiRojsTTbgdxh0OgctTCQi9CdupZZhWlBTiTUV
9vSzBwcmZpKXQ1dsYfXCfzS4LG2IvMji33oAKRUGPDM=
`protect END_PROTECTED
