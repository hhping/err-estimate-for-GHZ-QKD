`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GFiZOkzprZFG/K1DFyC5anH3QPHNSbu5Ouhd0hqiV1J39XnXWuF3fY5AkPUULohe
2hiEL2nTDhJtN8efuVoY4k/ydfVAmapao1XsppyEifft25gfSzOl5MA6Caya0jXn
1D5UqKStMxbcZQ8ppGOzK0bUaSIFn5Zniy18hA2D1vmBObDW2zR1n5D3J23awedU
tEgmppSO304STGE9b/eR+U0mafSIEvHPrZID1S8y1wSGN1lY6bYq7SMGWKBrRw3g
mtAC7//t5ZsMHGNXoYjOxQobWOeVCn9Qm0MuGb10/bXuQbF2LzL1cGdC7MyZfmxL
pwB3wF1n9hEtktkElvTkW58UKFd82SSxh7rNHJS7nazrPoL/TjbSlxYmrpvDiOd8
T2fF9VKcGm97iNTGLzpXiAtHg/krnmle2YJ3aB75dJEZBB1R/MRw+hsC3VbQ+K5b
Riu7bs9QGDbccsa+ebXnNYsIMTX3/1AveMEQUznuJZZZIQx6V57TK8g3O0McdNpp
m7W/63R8PLCq1wFFI6Isv/5wRcU4EAY4lhIE5C8S+5pdXDZauRCGyK/cRJlyFIGq
j/Z+Xh5wOCmhjdpao6wcdZI5JyvwLFV3+UKo+/d4nAlg3616rJsTj8Au/1vjGxse
AV7t7SvJS+317WlzFYSiwBoOYWblwExU1yZWcKOHjFzDMEtV8GJlZz4jRugx9Uoj
NP1u6aaoSbhSKVkJDLRpdssFaeYzlOmRJT7Eih4SrsCkAy05AWRsXpTESHEn4phk
HVmFlLBEagRVGjbJEFyPsGWncr0Rm+JR7DgGumyI0rdMhqNs/qH8Wnh/yywFas47
rlM441WtCyhPpwUn6rS3KInqAy4ZZUDZ8oKutIlkAuBiJdQ32wJCntMQqXkhgjiG
CKYc9c3MskuILUaCKOZPA1csOq+U67d1swspuDzj+bRFxOBA7dLa7EfSwpWubWuY
FzmpOkco7LUCYOdh58xZC9FsQAk84JTniTzHwchrU2elc7LhmUnisBe5q6WkLQgs
I3Wnesnq8v8/w0we2EunNXEsQCv2nXncO/SVb5GJTES0k2rpMsvzF9T629wertSE
YAzEV8OzreHfE9GrIoU1PxnIJXzxsUSDMBbBpSBgZ1DGSWWcidsGH/UdB075CtZE
2w/b09wdSkwK9Sxq4oH+7IpQvZKKnWV865AW4tLH20ZupTNMxoT9/lUUvcOX9Gh0
A/hiVt+J2/W1T13YYtm0V//sWW2wJrAtcVVVzxNEqli4IIZX5P+SJD6KV2vyxDg6
qnPBsY+v6fYDKx5k5WYjG365PZ3Fb8kMXshyBcL0BY2t6h0qEAx36XTn9vhkUhVZ
v8kYLH5B38yHSXTUxejtqnQsSdo3YOFx/MIPjOM1Feo56fo6FFcYWmtvWR9BtIOC
NonYSVRXXIvlNRot2k2tTGuJj7NB9aJVH7xDWvldu6VB6OBorm2AwXMdJeKH+uDb
VqzdSGUWaiHRn3og7tMpobApOSNF1qZoguzTOAyEQ9H/QdQwnINrRX3KP6Ops79F
NOTOWbt5/wdYr6UrF15UQ3z1MFzfTNPmpbf9pEsS/W4D9YfBYD5Ebpqt2TtGdAQ4
C5lz2NVG+fSMSLsoQuIN9WEqM7tUNkSYk4PIqgmvbsy9lunbEoz8rZ3KTLlc1dLj
t8u7xIfMS7sJOxOt3BBLGHWwSUfk7xuA+dSxFadXyWvPikKiF19hTdwGUhqs+Aqj
iNiyLpEH0n/GJBIgDh/v2HsEy4U0q4CqcNdjse2JvX668xKWSxWlW7US9n/OUPiE
S9w9RqNwrdQ2HK9XJeXCGGeD53osnob0c/2FJthyX8Pr5RnHI1WsBpb0Tyv/7GKR
bcitfAoL2cz+lta2dMPw1rqC3dFPsP6UjyC33rybwEgQO7dk6ZOA5iU737oEFzGn
aosQUnD5rugolcPIL032rgI4lWpJu3Xv89Hj+RwpSXXkHFjVJoAV5YbYPGlvXpk3
2+WHVvAt5ebN3AR4S2MPX+7FjHISOPzlmlTQx3RC98v5l/JAdKw3QuigmZXW1jmD
roYMQ2PseFlVjOx/+jW4mH3QYvXoJN9KZ2aDnT9Sd45W0mjH5HCyHTr7JwMtwvDX
lR+zfeSJ4ZTJUq67WaX+hHFgcQP3JKz+CcG5xD5enNEiuTxreYA0mAiJvXS9wm62
00BgWYpSQV5i6q8NuzE2YjV4ToOx3/y6DugLMQeRhqSGgu1I5j+qofPIJVXMhMxy
ubsoA68a58Vm7EcikQaTWCFdJflAV7/9W0Qd0qilYTBVbZvKTt+wF2ptlkBck37M
ENcNtdjURJBfC5SzFkmeCi3lqmLOUrG4k1mAEzbFpVb14wMR2sVTUVVXN7wwiKCW
XuhyIad/8hIhGczwGN1rq7e8KhW4M0hxj+svcDOOCvGxeCnkKc2ON2F47sQWFLJ5
IywtPe8oorwJy16D78M8BvTE9S7b5fb8MjGEJvixSyqQnWXH22zz6ZOLu534L7MW
XnLzjMJOYma7k9wavMBGue2IEzpUWpWF/gUMZb2q23XfOUIZVy/KC+fpC0HMF4y+
4j1kezH0BcV3FAZJlTz1300MaYcK0OFk/g3nAFJC22bScbChY8CoRycznCgsbNRC
HQw96xTr+iiA8JDzQg/CxjsJzcl7PtWdqLigGIch+3Y3n1tN+TL0feFnpk0SNeCl
jA32fY7JE/kPByitRCjYl9HPO/fSqbT94tBhwvSmk83n7pwD12Fj5w3OZEFsFFIP
QLnslgB4121vY/EXiJahL5Jmu98zOKRnwJefsBSTbpg2WopbwgZPHeGbfmjQ+AU4
WOT8Tnb5ZyhVDKsmwco2HK+2mTse/VTyOT3YjPNIGYJ6sNOtbtvMOGWwY/7evG74
HOXFpVC+M4rEeAT7wMSYpqXHCnvfw3TGXG5Iw/gjrotRflvccMNeyP/uQrwz+1eZ
hqDTUUqUHFtkzX0RYIikHHuV0cLb2lUbyPwVdUaXVAqx6c1sAUJm7yKy57KkuoPL
KmbyQIVuCHDC9SkmcGt69C/XRc13tdxXqBQbFxXPY12CXpvf4ZEW2VbCCGEIfCWm
8gpBQzadLCk9BpxYqlv5JBTVWJa/a0CRm1kJIZOXPXPvkKY8jIgfgQZJHh4qTB5H
G2DG3Vzly1Jzs01HLRlzm7PqA1Mr3HtCHC8LieFHxS4Mpo+Ixi1RIwF9on3A8zD2
0/IJMXBTshwnJJw3PTv0OA==
`protect END_PROTECTED
