`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v1jkl+WBy6+mgSjtyM6de2ZBR03kTfn5o3B38S7FeiqjZQ5MbC2GZoUTh0591579
56itkQ86Z6M94PeA9Yb2nXA86cfxKgXqCFh/iVN9G7plloMaS7+BzgW3zZGm2pi9
EAm3QdwePBRBNcbKZcHitl8lH5p7joZ3VhXNZObQwB8J7HP3MXJgiAi8m/HKooR8
emK6sGFzeN4wsNMqe+3vrBwX6o7+6LhS1rcXZ7+NNqcuvluj4J4NksOCvtmNwi07
tFBDngWOS2YrMzIKGkQc6V4jUQOPEs2ykjyuGhxQGvJFd0fa1G/NQsi4JLBaghfY
IszlUgwESyNBQJT6Vr+oDtf1JUvfVRuwWfPWzbNVDETwxWLauRfN1wsnoaSDMaLl
P0hIVhjteh3HT7Ng3KhSYkcaUkF+apH33q6EfdqbCVywptyTmHdM72cP6Foqn1hN
uANq9YNyx3pXe23VEQ1pdCF1LgSBuTZmXnJq6t9jXmAO8WaDFb4eXaksSu4V5MjG
222X3rhaYyWjkcs7TCad7CRV0uLsrvoLcW2DYTvbVDrYgUMBdErC4bA/dcypp+0Q
2ZJZijOqW7/MmJC+NE21+R2Ihanfb61vRwGk5C39YWpRtJIamw71C72dHJs5SxMY
4D7dejHmTFyBcGfkhl7oJItOk3ugeBqThfMZ3ol45ScfrHmsgZkhj4pMZMTKHDwX
eQ+mRv4VVhWyo99torJg9GPvH+XWIbloroIAqbdjzBYtR4u+jGoq/7omHomXZo/Z
YksthorBPAYDuvvU1knvQcqCAjQM525TTLG0kEkwRxCTi4bEvnbTVYys0+7AOtPk
BSiLlUt5EQhr2LXa175fPHlMjZdzoNVTGgYxE/H39V8n8cgpmiuWjomO4pT8Bv1S
g/fggme1vU6B7zH9dIAElNkkTRAebJFQ0UH8IgT/h9RiASslzIqqYdXbZP9Xtoyy
IsgxjvTGDiMM2ZqUn1u8B1IF61PTPvhVJi7qC4h/vjrcDW2C9Saa5Wdz8D8BwbWQ
B+9F3xIibMsLeHmwpPS/yDtqJ8Sdsmh89dXoYAIoID5Jj7QzMpeTCuAdWerhvxPk
iNBBlNJjJqAnXQxvVY1WaxXX+ZK5pgHJhTyKqRq8GwWKrruc/318pVruCHjlc5lw
VIpx7IYcjkI4o3k9WjjKQjVZeIKGenZIhQfxqXBIu2ZjEhQ44D2u0ot7TAEU3t3F
voSUL6tZZ89I/fWnkMEPlh+JKn1XL2CJC+rfr+V77VkQ3T3XlVANzOKRYRRf/mGL
yYEujgeLTjy7iYPPnGcDHgkcjvTlXAwcRiUm4730rdlghNwNR8KbpxQzqPe7HHQD
ykw7Q+221nHGrTMJv7q1oL5CTRvb/y80zVaKowXLHRdUvmE+sVxglpGzBgVD2iio
fuMPiGWLSAXGmqvmOh1rWzYMLUSUgb2dPCxo8YV1bCDODgUfMem25hZ2yoNEwFks
qsERpusKQndxFoTzXyzb8+0GeXkFfUyB14VxaWJuUn9gZm58MkfornQvzyaUz+LC
rROs/VHRL+XU4PNlKt5+m5VOW1gvOrhAFz77sDFE+Wlvck/l9Pq98ZzU4Owy5TTt
H+5WE7FcYJYZ+VEcl8BmN2bTbXF54BHje/0MTgK0jxCRcaVLKbYt1iTM/yI5F0sB
umt/IqjudYhreA1Xd3yBHQc6jLcAIlypOhMdBMwwwYaxGoqT+qPLOAZQbWlk7JR4
pcJTLROsieAb9Nkq4LIoVBu+zl2rMfDhZlrpw7M1rpbsYDcVoz+ip8xYEabGI71C
5dL0GB9F8fmUT2XivY5LZH1a9GHtXiZTBQrOCqhkOwLrUiUZV3TrACJtPJTzrstE
rAiPXepXKF/KpgAwVJ4y8e/A298qta+kUC23bHAb5ldE+FX2zwQYIF/KHOUyVK/+
6ofyHDmMceOxzER2vqxTWdajZk/qI8jR5oSw3ZwSK+h02SIqGwR6AzDwO8K+qn77
jKU4rwLhWs5fnznhsmPb2t17d6Au5bu8QQAHvNYSEHt6+2Cj4SVjJDxJvrUVihnA
oxMi0GOH75ZquNsJhvqpS5THUe1LdiYnruvLnAarDnFVhCouVssYvIOLzmTsM3xS
4Y+vZXGWHucxkUkrsoZ79jjI1jsc4eQaKliIKol6BYFN9uB6eL8bms+efECM1nwC
Igf0eWjdh0N6BtqYlud3HhT8nBCJU69ImdXmFIpZQBXXFjJa4gc4qn8XHWYPAPUN
2nTjdDi/sOVaBljKXvFBUmH72dVgXPlQMP2DUO+KZCSg4ym9XnwidunGsqxV+NhY
kIhTrAXm2Zu5beKOky4YvRNI7Uw6UzFIpWOtlgCbnNheL0Y4MIaumA9itplrxtZx
uha6jU8n8PT7zo6HH2RZjKDJpxckwbGJJt/lJ8s4zUB9gtIm3scApoM1euqd1E0U
wKmGuC2QHcDkhfvd831G5Xn9oYp1SaNkAkRpRe3BSD5K+z7wCaRCciuw+AzMocQ5
U6HnssQwO51y0OFrKOVacR/yYlZgdYSxVQUHWNQHdtWiL+u2pis47s8vAOKK3zrB
oHL3oV+quFze54rN1PdoIMXH9M0a2uE5VPs2VX/0ERN+7eMDTVSvADT5M6ZdkNuI
ppOuhFsgyocqdLs1ULgewYNi/9/iQJCzsZkBePAXoWjqeI0VK8L9waz31lVsEa7H
RasPASVkZHqV2vuKBu2anBTNM8inBcF9I3sh7hIhpKt5zKlZz+yJmonQkDFO0pcC
O1N893It8bB0ymPZzfrO1cMddW4vo6ZxVflH/X8VY7RZxa1D6LdvWDt2jAbAKj0n
iDL3p4uRKKlMNY26nzGsW2b8ra/oE4SrDFOpr6m56GsEOJKGCwcPsINCkfu/29SC
WONqrd6Hj41itouFDWs/J2byTUhJErZVfqmbwT5vH1wEb8tQKAARwCAKGbtfzvK6
X5l1H+onqPp/qu+pnloSlOjWaXhXx29tNP9b+MhkGQOn//QiXKHI44bVXNZl8Ix6
n6+j1FMG5APHhrovStiVi2k9hvkL7O76LkSM70d5RNabDJABiYwQQR+vQTajPKFt
8jWfnqhtb7MltBdqtlVk3V8UN0sVWGpGC4Spx4bGj9NY+JO8Y4eC1UmVHLMhbgNx
zdoupxjwthArUjgXEbE71N/KiW4TxTEE15BIBYTcudMX+AebD7ky5m/hrWYF1PUH
d9Vvgc0sQVq4cnbBV1IQqVJLga3ROdZiiLnTIyR+bpqu6MYYODahwKl+rTI2NfAl
aj6RbEy2ld39vOvs8qULQLoiuFjNgmvx7Re7WiFteOuUjZciiUFnQGmZb+SVzJ5R
3phdoEzM7hZaCawACFc4WUlMag3586090Yg+uCrq0ateVGcVn9W24f0BPf8IJfad
/PS4zE0WS6vPVYY1XbhjZvgLUWGNaVNuS95WMriPNY+j8nGXcbe6ekqYVVB4UGPk
2govwqQFLpznqrp5a4xjnP8Ai3c7LKOhzim38N9G/CrLinzO/9yOCiZRJaKw5R1p
k0hwK5Qu/UrsUjpF/ee0UboelY9jtnljwagbEnaGtEHAsWafWsAoWHObBWHyYHCa
zZVeW0POWKN6bDeyJ3S9VLOa5RoSPFnSetDbWnxHTOpzt5t21NNf5nfsprV5SYDd
xYVAASDlpVcUTy1VZFJa069/4xP2bagGgTDYn7jCQSeQO1+crNJSYtEKn8IBwgRy
8zYwvNciAikmEcnp/jb19WXQw8wRNhj1Idnrb9fXk5wVtBO4ig18Kffi26g9yQto
28tKvYdIkTJtUIs/QTqvHxNLCGPl4U7AOL2QO00tK2SlHcZ7iS7H1dyx7zat0A+j
7EpgbEU67+D7mKTEybm+AYENyVhABmKMeJFM5h5EvNwNT1Nz5ZrfK+WlfuAH/c29
65qlV1PhYVQY+lsnJ9c+QOCqRK9Paw/dydP4H/A/pArJM/QYfr8iN1YtMuiRTm6n
QprV6b+LIn6OjdcSRRUnrmBDmYVLGXsfNfd549ifH9Z8KiYP8ojKU+xkaGJtyUeY
kJ/EysTv0ST6qNAJJIFb4bYt71maDWz1GcDIDvaOYfJZSIklrvS+GR3rufWTXP/j
LzriKPhgo+Y9x5tC69jPjNop05NWF+XPpu+aQlkyIsoPAVOci7GAZvVMkp42/FXn
1DL7y0Cq5+l9+nplnhc+3sn/m1b3gRxHFpswd0OXN9kV6cQ27oSfYyxDpUjUefFV
MmBWVjR5cKzn1RtEyKcHKCA1RSQp1ppImwWjFoFqhGbUFPTyALIIKCvPXL8mT6zM
bPgtol6SUY7EllHD6BxE7jwslQAxjOcN3q7b2Yv6KBmKHOfN+dnBknv+U+StPuLN
DQrPoGLljIntf/YbyV7Fqt6KN0DiX17MpJgXw2p7AmWFLG1Fxvqnd8byuuaMZxn5
gDe3Gum7PtaWaM8FNN/9/KtUpAmRFxPK5yFvWQM8PtCVEpeRLDOnaejDGDkuO/lV
YUbkNunq+Pc0KEzDqJW97PwuruvQuJmlCvdaPAgzlkVI3vHqVmyqZ1WoSCnvdl08
lkJrL29COPPHXzs6xCYGLCVaDouefq/28eo4BB277ovcJIMaeEuyvTvVG69Ispho
EzITgUya3CiW1b0Ofq/xkxWdN9mxt7ln0k3qMdS364Yn52SkmNphFYwpNnqTR36G
p4jdFE2TEBDRV9vXf8ZzGfUIcJzw6/QNmMe2KID4k3jMw8rMc/yiSdJGYqN/mft/
joJhCH6sA052K5bkFyzGXgpXpNhBRjuGIBRKCcfqcmdb3k74q4miRPZ+QSfZRW4B
j8MdrTjXE7AICCMcJMPOmWgLe/w71gyGaRZC55kbwdH5A92Eap8WoP6uJCBAKSN2
INcAAH3nOU9U9EDsEhN5qq7Ggkddb5XBEla+MyGSh6jF8TbNUv2K9S/vMi8x9/kt
/COBzcYlf/jhmh2o0BcTp1i14KG+x/0MHrKzPCwQcMv7TZcG055DyGXsffq8e3J/
0dplOR3otPA4HRaxDKfoy/wHFSJ+DLIBEbE48yo5FIKLUNOkCq9Zg4N81EkYt7ei
K9QLniIbL6A7UrBKV9bqgisuxE6hnJngBC6Le1hWkyWDokQZqXdYcwdVY/rhxCvY
jv/o5l6IhzlItwDBhluvLeoX6/ODxqsfW0L1ob+eTmYiZOGNh4q9Sr71oiLQzMk8
+MtbCZRq7R43jSxQCII/yHgfCeZWjV72PegN8kKPHeZDQl/RtY1OvjUXmHwUAwrw
q441Nj0wimu3kfLI/Xfjim3EKIrpWGog+xD1F9MWNtrHwKV09uE7FlEMC5+mkdJe
Ntb4CR0OE9b/bUiSpFuDrooz4+x6uLh0m4wc5t5nmt2YrWryJb3fJwLtdUsU3xgV
q16xj5kClg3syDL1NhXZPRRt3h6QY2RNPn7MzdTy7LhS0ZO1G4/6cqXBUOm31e9z
AUmx4Jg08h0gllVtOT0R0kjX78P53rt5awXaLR0oJwXJSKT8zHt/DntnfXoIytM7
eeTyA8g/2RQCV7pOi1Kt3mxHBLsTKIDdV2OfbPHcdL7lL9EowAYgGgoMFPJvBJLR
qp8Cr38WJzNs5R3HU+m5X34AxwqyQumCSuQMOOyS2XhaCQoQVgL86GKsgkt8MfY8
Z+C8lm1+Qvci/uq8bc3BMlM8Z1QJ9aHZSSK74Rx7YzuppXjBAINqRsz69aeFB1Af
XYPb8moyYHGRh8M1nM9lBJnQeaWkguQ82EejRGZEX1m6asp7UyuIa05magpSW/Rf
ZLYUrZKKw/z+m8UAB7Hof8emOamZUHPVjc2CId1brSiGe+BBFp/qpEfz8cbabwr/
zezpLaAHqpKlfNXyd7rAOVNIxoFxtBVPb5uTWAENSFJIacXle68yi5boZ/OCtd7k
gUkOkryyyuX7iqWQiYwd7A==
`protect END_PROTECTED
