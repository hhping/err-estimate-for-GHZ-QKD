`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qHYz4CZFb9uUiYFzZI+E/vJM6MOUH9dZetol/3znBfk20GlGCS5iFSWYanDTS1h1
vXu/Z/Luu3XR6ETpUT8+NEWzH8JaV03/ZE2zaoaB4ji5Hs9sXK9f9OQEESg8h22z
u+e5McXxRwxmg3I3qHM84EbjrU3kVpWJConkJ5erPg2si3PpKDMnFizQ/DFfsg3L
q1Fp7z/rkGYKS34jv1OOONiB86u0OYsQanvK2XhSlOs+ErO/h5pLns0pqH+hwQ8s
Nk/uySHaG0whSEwiUx9sj0Zl0cFMBnwtnoK25SCEsrVxJfseC/O5kAikq2Vr6I3c
HAjrkmYXyBEua0zv2Ws+qPmusq9o0tQAargWdePSxckkG4YtzNeh5csECkC/E77/
0PdHmt0wzPxH1DY4Lw6wLDOMPRluHAWpcPqeZtrdpVW9Okj79pegkHPPW3ZaSMTT
6BTMkXMkm9TsPWrrS/RUqRuEnO+OR/hVB69uovPxo099jal9qspVjEPX0c7evKaX
NAa3Vadj2ct6sndvetD2lvNMDMIzHCX07QRf91PEbJr4JuTDbnq+h+e6fvP9rbMz
+Tz5QLjGXX5P70xlmqjkr+BpH8qRZ+R2C4UJxOen5zRJtAJ5YkYgKUPFSDmJF3hQ
3j4boCXTcmbzobvBpwtsz+vGHBCpnSK1ktRHmyYcoNsUKA8i04qPWfwsWaqkuHw/
Jb7SHhR04qOVlbaPdRyR1BElgFAjnZ3r96CxwrfOPpOytvC7cE3LIlg5UmQy9San
z78quTAIhoF3lzQQvgEWlFbDatEp41PjCOY91uA19TX2SZ0yaR3KFYMrIy5SoMS7
YGMRXoXAyr3a+ejinLV1gmRPveofnBk83iAmc9HbY3xoUrmXNTDqNXWnEsV5dSKw
2uMDH/KCGaZK3P/jeBwoIN0HEOL/c/PKoiluLhChdGuUCSjimVyibXeTH9dLC+92
wKSWVEIDb5xlkz4YQlJ/S9PpecrHTiJmfxzitQLxcQIERiV0Ov0NzgEzvz2AcrDD
IIgiOiGyxvvL7/LW0D3qah+juB1Z/+O9vc56TKwuNrL+y7M/51JVI7JmVn8tbnx/
`protect END_PROTECTED
