`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UZM39+Up6jZUkvwZtA4oDLokLh02hiw1fNtaPViaVqYs8VMGKPZ8m2gCOx8Id0Zg
8S+faKS6DcNy253/KV8MJ9eVAkYIoEqmlXOTkr8ZYNM9dqkOtzTlDMnmGjKN5Yi1
jZUdaWdn5ueuZpGnL4IiTk7mwrcKpEKrmuEbSdm+Fge/5SjzAVwXzJfnxQIVxjWq
MCRg9Vb+mVo/F0PCvQ0EU11qePoWfFp1WD5NfnfT/3kFeDBLwQ17+fmlJuTdnXpc
4QG5GWujPpsIpWiah4W9C305cRy0abn7xpeCv4VLnDRHm4EtxONwQlsvRZTxPm95
zX/D7zhdd/CGbqujuIeVQ8YELuFYeA6fTnUjbIAsUgiPBgoH0lAo93NaDqg5NOqF
BJ/0yDa33S0JodHNN/jz+iYUy2zJ60bkhmj9lXjQrAaGv7XwrVCXUm2uv+s/bwdI
p13Gz0IYfDPyT18t7nIs9/tm8RJLOL+6ihPQ6yJbhYgxLJoLIQ2BcXPMKbi6YRRD
`protect END_PROTECTED
