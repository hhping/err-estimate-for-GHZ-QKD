`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iceLAPELUrOiko8RpodU5qh7dXSgZ7Flkss3hMSeRW86/o2mPRvf+cm6H8dWbaPl
IyrvmhmXWCRyzeKJJXDX9+2dXazvqN3KR8WiaTcwzyVBUEmdEXNt6YKsfuKAXaC8
r09pJiK5MV0KlYt4B9KIRa+mLUDdZB3XfCmPZzWAewT3Txn6VdA2RuMNCA2Env2Q
dflYKu10/gT7LqW3yDIq7mz7UxAuZ1c8G6B9VaQKA9HxLwaG5UxfQZEWgnO6jqh7
w/LheqtJ339++R/SBHfZeRRNkN9FNeH5h54IrFVpnnQvyH5JKkQFrwWFOv7Zig3n
nk9hmgWo3fs3IhZWpSNRpqN1tI88rvUcKODyjxey8N2CaKQfS4wyc32EGVX/tHNP
heWHRwXgz/2X3rRCUuEhc8cxdzvtDTbNM2YaWSrQw1v5u4KooT9GSZpsogyhs9p+
s/4haxbqTLJtclM+Hr+7PS+bbLMJ0Fb0KPnSEfrG5SQD4GoM80GPvYRxLYgxSZil
lgMwFLfRMLdXYiuwTt1jwg8HUXFM53L5AWaKzJqfGTmuqBVDVXKrqGt0IXshWgF1
BP8sPIIkExan/Up1HelnDmu2YGn9bNiKyxJtyqcpDY3uXOA5WCfXGnNHXNVYGf//
dWNBixnIoD08Rp7ET8JW/GOlQ9y7swRhfQ5/8/FDVTFmqE6Lnqt4ejck+QX3eHfG
heYNizL98lCVD35S994Lt/6Ufe+rdff/OLErvjWHozSxOk3FlJyK2VQHbWgZNJRO
uX2wrekIvolpfwG3gPvouA==
`protect END_PROTECTED
