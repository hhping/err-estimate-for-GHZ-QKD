`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Us4t83RjK2olSflhT8Ma9LmqRy8Cd/7gDcwdWhl6qpGPiwEs70Hn3xkeDrZ6gPAz
lbESHB4LvHHD+FBNFIrbYlQLvBiM6GBErbqH0+FDEJ67z1tlm/yUO3G5hquWErb3
3kXU9/Wm3EdR3M6BSHTVdsTluCQCrN4tDaI4TJQMBYVplO0iEokXPDY6F5JgFOxI
4E2Jp+UJHrfUXH88d78QQott0oZl4njN66fybBFkN9u+KUN1zq9c4d9OhCaiqN2w
m8cTHZhdz77UAe24Yslpb/WCCiIKgoKkgB2+7QbxGvSH/btkxAY4zNNdOdqpWsjQ
IWORXzDUnb6Bl9Pjt6Ty4LE2U/J+ARZakehe6pB8ZOAGr3rLP+nCGh6E8SuOhssx
H9WcNp4Ow1czXXYJZvt9AYKhP6LgQ/9qtjMKiBsYlJAG1Q8BZ3Y1ojiYq5OaSMXr
iFcBvPkfRsUbzo4kpgT+UHgFhWPYjilo7G8f6FqRiFE2Kiag24+7vbr2r6tEt1yT
iyaF7aEQGv0mqGdWlfankWxGcXUsbjyA89T18KYDPHGdq/7STXhUlklbHKhKjE8q
8R9vtU826JVhS3AXMF9DKFtlU7nfRJH4i087qfZpCKl+LPpLb+KuJfxfWpJKIQpl
kv7wWGkHwdglUj+nqMWI/EDqrdZYwVU5n4Fv30Vfh/NgtjlmqJbQqxP3GIvux+yU
Ekrh5ofSdvMbt3iBJUJMl/2wVSmhJfILOIgXxC8+hSG2EmfRmKU0REfi1H0VgeDy
66djwHfD+Wp2EabzxPb249/i9I2a/M81hyperk6OqqrejAeF8kaIKaAZbOOfDyVv
mGcoOScnCx6vvn3+DPeOe3Xxje7afqrGUnKAxYme7TldfKRCtHP2Fe51sxk977tP
Px8PGBxNJ+Jsgzm2HXqegYiA+8XHlB17txWT4Z5FE02EC+Eb35xFEG1Gpc7BiwN+
25dkuHtUXsj8hPXycOJsJPxNUe2+7IosQYrokRIv46Lv5PYi7l4BAVI7JIZMecI8
dK+e6Dh158jW193qvnYxkvonUYj6+pQZD1TVEMZzNbreuICg5bX6/UzTwB29yHIj
OV6XW7+xrdUXqC3E3Gyk4uj5YGFvG6nIJmAb+sQYXpqfO3ztLeF0VMfedkMVYCel
2/f6+FgZUl8Lu/K0Zw/v6ITuI3A5L7EHy82fmhHwAE+9YxNPyQTb6N7M/StKj0hO
w6WUS0jwCNzPGFMKZeai/z9iTqooLAvSJ/N+OLciMN6Yhi+EO5mtD4BF4vhsqeFc
de7G52duxG5L/ANJWNvP6SSQTJ6+ANsYh5q0T4Gixrlz327MZlNd+vBmd903Uu/U
`protect END_PROTECTED
