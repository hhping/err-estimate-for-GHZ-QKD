`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BIT9LYchKePaR9akpsVayh+QZEhI7hRR/fmfxTFJseMaJzLpvSvU+FXKfzkJViS6
ozIgskPJNnGLOxCXV6PTGMff6pK0JcdxM4fbW0KzlRayTQQll5svqTV84y251jyz
/36BzfzKMczBzHk542U/yiOvqASAiUPrXnKm+G+QRUM6yK7oOPMf/iyG46UrP/Fn
DID77pwsXG80agZRvhNa7fvdBoK+jX5sVOOPL6yE2mW8GlgOXSCQlVyTq+yXjVEZ
/rASJjwyvchrt+LZTbvvgvZppiiU9LEVMNw1PTPuusrTxQuEpZGJPOAK9GkNI5SG
mCG8mnKwU2ZqCk3wvQbZT6cjqcAhJ/AHAIYz0Cv53m6oYtIXPqaxajgB1g7MdQFR
nnbz4tJlFGUrpNKsvVlNAkdUD9cClBlk1ILOxt4VsT7bGc7DYSqS19Vln/mqsHVn
OkZ25oGMUfysfucf5Vg3C9Q50XTNEfIhKDYJEPquiTmj1pCLkkMKzOgp4ZzvaTvF
Ob/PSnJ+/ulfamDD771UlAMtEZH/k9WV8TEWn6yp4Cpr6XD6VwLCGyZlqL/rmTwL
mYo4EGRKkmwycfws5NLA4e6DbzDwC8dYFgJZk5Wpe6B6LfLY8D4Qm1vS0pU7zlo4
ytELEkB/3Qt3BelsEeiTWAJclEErGiS1Hsk0vGteeXWDJVylUNvZvT2okm5VtwzN
T0lI6tpAb/7nCTdB00Aa6aynmmKemJT1vB/4h1pZBx3Q2onouulZsQxpgVy5s/0w
SXeXkP5z5BqeVRvYMyemxBerxmBNY0bORm0NRLCU6Qz+FuQ3VIeZpxm3LFfPgQsG
xDsnOqTNWhhj6UgLAHfBuI+S82RpanYKalauXrhNLWDg/rJJIHQh8BRxqG8EaFiU
jD+EvXP8ehSmyLQ7rHHfQtAqRXGpd9OmWQe0QHkNFdX/ezaY4nw0iNsKVdcwzm4V
8bE9jxhnDcEEhIV0N7hWqcRl4W63g5wDli1RXfP2/mxp0XJuSBFjjkZHS7EbCV4O
P3KgGL5Nf9+tlVlvHYEPvZmcoZ5Ma1n0f3hSnW6ge4hZX3wqdwiwq6bSSNIEwCQY
WiLH5U8rGsmvGYOPQ5XUagD1GRU9RkziZ8pxQboLU4PPMHkYC6+c+/i0RWL6ZBit
XJymczGvLriWp1vMfGqG2owBKKnG4KnJ2mWy9KqNAmOZSbC02E1n5KOSoTnajEfL
q84ZleX9Car2A9X2cVA1pOL4bWp/W8Jkg2TkJw2OtuSeDCLFdrBIiUr1I+BZr0uV
Ve2433cLLqjJ6LqyOzsWN5qpzj5wBt0rHWmhrU70xdy2D2tDVFN2cuXehC8DAtjJ
d16GtCO0B2aGTxVCsvnS1QxdCrDilHPAvE6Upul5dbpfqRv+x0av4Tp0m4LEoaTq
UecXhqyah/0iehuh6mOVjJ+pbiZq9RjAjm9qeJPTIsk=
`protect END_PROTECTED
