`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nr/2MT+Vu6TKM8J6MGhh9Iynmuhz2A23eNDzSWolFugfNKxFqSw9jxjGJyisv0ny
olE/RAvpITeiHqtg34KfGErLNE8W9dvEI63hmGVpEAArFEeo6uWEViAVQHOjML0A
dk979AdZXM7uAVLj1yw7asZ7Sy/quA13wvok5K5nw0N0n52mkKB4hZeesXpsilkK
Thp1axEF1DsPJ8VNaea5gEFA0qUg6OZNOvYdCMd8tFnNu5yYDhgVi0lcRDQDjt1T
TgYBFILC63vSw/wpUo9t0DgU9JAhI6JfVD+0G7HxHEo04ffSCCfnSvIHjEWn1gkG
Ow76W7XM8HWGilE+QQ9/XQi2MXDfHSDwhUbowpg5GXJqzofIyY3dq4esVn2Sp+1w
OHe3tL/GqEdikpc3i5D1vqg5dB67yMPeJCqwBpQK3iY0dawYvlqgLiICwOEoKwKx
raHRfckC3VA38Yg3MROnL8FGRvH4hOzRn7DqDoGSzWZl/evRWNShamO+cCbcV2kk
Gu5KC22o4xrBEZ6pJxB6Q9aOnyppeOF2V+WVHOhn7i0kjws62uBwjZWdgoyaU0z/
fvrcRzU16cXCjIPDcL6I2xBDIHWhfhe/YClvUeATaOe3XC5ZMU+lJJz5tZTr5BEG
G03Ri70nG3Io6GSLtX1YRrLH/ZlNJNNmM0cmyRUnOiRTVrrEMJNtce7QdSXhdjwv
xLN1MhAjLkKXzMYH68+5gd5mV/12SZ7k80f7Oe0Nzv4/dd5So2IDO1pzCDMZEaVw
zakT/lW6M7X3Z1lFtI0GmUTLcNEL4am+0iikZCSBiBramWxe7qWLq5kefm6RfJMF
6oMo0ZlXSX9zKSMx103WN3fEZaAz8tKb4aotkQ6DCNoau6mr1KTBtbuvS1+yW3uN
kJZfCruN5IKGpq0CjQbA3MLnS1C2AzMN9A7lSSGs4OYUz76H29OnR1+z/1BIOzH2
bTUsCQcNDjHuhOBQhJliVs1SGYDXKuTa+Qkj8mQ8/AG9T5g2blOMxMJ01hmDFM6a
FkNcFmEv8wzUEMMt9Diw3/3Cm9YQBq3YJkoY4gj0KvpeFlyDbBcCY+nJH39WlKzB
yqYvEe6y1bUAFWxDbJD1kSOcNeOQefzyw9lkgUzH8joGGg9yl+ChZqTZm0cTuEEW
L3mwldFLZpYM//LU1/6rCrzaRg+5XCqhLqU/gPJoV7D51OOiV4dyaVFGf59msAyA
+O1Ih6omgUpSiB2+BLQRdM3QM8bTQ36/p2m6ftDZGevSUK6YRFlj6MiolJeNcT0m
HjjM9ilCGTfznnxjbKtguyrGLX+A0cNmAzJgQTMMHLhCIRf/6AyPhiIfOLkvf3uS
VuHeXkVT4dxdzextriiINWfibcRRfZK3xbHmoI/jo8dnKKSLObQcYixhnaMIl+h2
jDKVmbEBjjY+SzLUTY3c2R3ewFCU9VEnQxOIB670A2u4QDaWw7p3uSUoHDp0Ctx1
I4AkeCtYHSOztPCreZIe1qoLXAWOJq0/COCrgFsgfgKPr2V79BQyQAFh88sj731E
/y/D7m7bVDd2T4Acyxf5MTruN+ypcVvG6TA+XBfEXciXG5DUp/tP6PGwnzEdHhK8
t2agn8Iv+Jz/oandlGFgh7mAvhi8SWE3NMkuigCIL0NOGcZIF3Otn80Yi9JKTKgm
B/jagv87pjqC3DPOj+a1uDW2v6X/Z/IBmMC2Y/ABo+2n/zcrY0mq/RIYBYrOnGtE
ZgUcCFzCqIegIiCKrbHrQEicATliFvu7VAr0PtssCG05BfI3Ewg7HrN5BX3cQNCb
oII0F5PZCdRhSa34/TxZXfzcPP+MY0ZxAKN3Q1WWSxCAO7HNRwnJIlcDT/Y2CW7a
sISBxMI2KaiR7XyUOnh8YAK+Mjt0qaS4d7nG+Y37GhfFbDYtmk/9aTy/jGvqwItO
okOSp0ybhvAUqFPgbomJlchJLW9x6EGvxaY4EqRHvCSXl70YME7YgiNqtX4DLqmL
xMmJXjh6yhCmnO/ScdMyCe7LjBXcbz8mA2oFRHLx+sygkk8Z1vSW5VrjwmpxZiCS
g5jLkC1NVu7LLeejEywnbizvFbrNqgqfy6ajPsQVY6QV5yCctpAnzr3/POzRdo69
0E3C723rBbLixRQKRxWotuHofMAjco7B7pP6P3oTlJnkPy5I4bkIBsZ1shII1EgA
Gsv8mygdHt6cLUdQKle8mrh6beq1mn3Hzy1cE0H3vjCF8vH9n1la0hx5TxV5w0+Q
9ffRsD63aIBtNqjOK5XhaiUbmjH+nSxqTodtDhtVksKR+rvHLYupVrWgzLC131kY
fwdzBHC3sxDaLS0gNBkhRG40ViiQ/Q6WJChm9eSVRbiQp47M+bxXtpaoxi2HuwSQ
ylfm3m07oZi3obdZWeRHRx0Gi9y4ZsCv7usxAhdBocRYvx6u1vojhDKLAbFNMkU8
`protect END_PROTECTED
