`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y6tfTrd9psYX0VtneF0rEOHKcuRclyw75ZX1w5L46XeWoM7XV0E00xQo17PBEUqK
tzInGJe0wAE5JbI/16BNRlpc7ffWU5PdwU7a1vMBhae8OWOL3wgJDj4C6cBd3D7H
MFVL/m/RbeGTzTPYN6n5t/OSrNPPznURy7gPtyjsAT565rnh5Zv/irwGXYgfU+wx
mvvvCqlpUPF9Lg4vqrD9CYipFZw3obrl2er5XdwXrUy24f+XivVmgGyUX046hW1R
P+AQNyd6JX2nriHL66rhxLWTqiOE7Qgu5vBSvhKfta2J3u1GSNwfx9Zz555kAfSB
JkxyoncroJZgsIWZS86oBWkWFBoysa7nPALxBKL16ZW3c4p81YN4KfBZXgFQY2Ql
1azZHCQe65RthFK7IEtfkO7LZq/mQYRklJ/JhIXikon9TpKlKtuMYDEoFTJX4Ipv
3s7Q4bSHUFYab4805n0lKlP4J58At1I941sjk+HDvu5I77a5kN4+kWgZ1/fQ51hv
4NCtZubeA2QZSrFknG6UKVguTXg0NPb8R5Y5pIn/ba7dfrhyYbNswyA3Dhb0xwQx
ICWMhXYjxRaH87k38mnHF6RunciiXgr3pY2G6TVl0uNj4I/MObUfCl4HNtekQpIy
yjK3ojwZLTAro1lQ3ZqRlEBEQc17G9R5QeZR6ALLu1fJIy5j4h3kVQDMrCkh8kPp
BVHaUrnadFxiRICs7eD0kAD/dVOdacXYWi/kH+Ji3cptH+wOyTIVN1HfJ9uD3uXY
K/uVr2H5F0TiuhkCmHkSzTazJbbd7TJxjKA1+Q1p8k91ojVZgfIHoBcPtC0xmAmB
Ofjnoe4aeLXI0jX5jCJKe/sS8JzL7PCOBlSAQJm8FEOBQ+mMtTe7cYcNDM5DYBse
XV1H6PRf7pfb4NQMTHjhD0BwOp5BIMma3s4EOruftYEn0izPYNqlBIIfqZezy7V+
7RW7+5f2TE7BmwAP1OVnvE91laptVu7XpJXpmf4QJn+ZLnVP7JPs9TzbKjCuualO
fCZ/HrnIdDX/2bE1ilOieJxpRzdg+g/elT0MbJ9r9VYYXAOmPsdrsP6BSXnlA6Yd
NOaB2JKhjD81V53Ay/1Wf3KX8lJo1wSeBc/67EwyBsooPVJ4cGMKzo8CPot47emO
Vpo16HC+xRd6mWi7ibMxR4kzyPpT3KEwItVTxqgcT7L9QO7rb/Y3uRnF4HyF3rP7
CzUkDJfVabgJFa3ZO3rb7BCf1Ewd0bzzasgzSJ5cjF/zm+Hah9NM7ijt8Ho4OIs4
u5xQvQz22PYagR2uO3KI+fmeTui58LGPHbOPBT3tCoF/XOqBq9mgvzndK29vWn4X
OBi2KKlhaTrLO75P6ds9WGJ9QB7+5UcCv6/e8CTJpspVLG2WKnHxplQxdlw8n2nM
VTYj9ZDcHQYNL4xMKYlCY5gFzOhhY9DInyyObw07E+aIc8IsBodaM8D0TpSqaCb3
Yamp5fQJCT4WFeygVeC/0DeyilELto0ycgfmyfZ1wIt8duWqozlcQ2uenEL/siIw
p69SqyWnVuncMB9TgGYuWsYeY3OBRsGGygCHOvKSiFiBpusnXktAvD/VPh9SK4ug
ajJTi09fKy1b5Jaapwu2xoFy8kfk1SV0hmhJoYhNy5EXhrEmwgc8iNixn7Y5DJXG
T2hS/XEVBbQJgtS0862WPrjxhs2f7nb39p4EAC0jYp/gTsW7CpNLFrzSxrYfidRk
BkNNtdTmAp994WQw9hRkfzlrKGk/1tNB1YGxmgBUBDCc5V5fya3hlQHU/yKOZkJZ
YqhLkgIUDdIirM3kfeKG0CoVZszlnizDr0njz3AIhA5IZ2Q+Kc5k7byxmZmnjusU
u2sZ12niLe62mFmNj43i95GsvooxUXm0ZfbslClFz4WxZvUHn//O71lrIvp76/OZ
GZJQkdRtRbx/u74evAa4KHLj5qBgPqOktGF0ULYmM2vYLdJHyfLm30b1Ujfu9q0C
3U3bPxRwk8Ys/2j7KHapBcQxhHhConuy/1TdOVLzdb9nn1OQg2yxd49ZxaqtWTRd
s5hoRQg8cfLq2t4pnyX05Uz0r2aGyCPPPvVNxPVzMcmu/IisN2MMIHYqdhljy1bV
jAfXQUOP81Zvhl6m71yMHJdS9zbkg1hIAuhMnHUrfOmpVBuaBdlN4suVFQqQ6/MK
h6ZSVytXK7KX5yezIAAd8nU0AR3ruQYYhuzgYg0MjsfanL4rAwFGQ1AzzxO7jOUe
/NF6pbm+mDZFESL+p6t5J/B8xl6f4wQD0KGCWIwUmPzgqIi3Wu/tIu9m6bp9VXX9
FLAjmdxuHX2xsjxqgPZpE5tCdB5uDZRZHH/CZL7xRtBttmkrOUbPZY2b3mncm3IN
y3qRNNja1Qm7GFaU02VQAzOXbq8xTvMWbKbBgFXVH19uBUmEcAikUd7RhgWSR5il
+k6YNQ2OYpApbVP/jtpPVgSDYLOqNvZxAKfjrJxQAuz5ssETEe1Gl4peqfE2AwqI
UwBCycjfCXWIy+Br5UmGP39+zqfi9C8wHwBb1ycK6KwJRqIYvYAipxB5pci60rZe
NlLS8CAJwFPLEbOxfOZ/Uswk3kk2RTDRz8U4EkLJDfmUNWYoGdo4StRMDkQZcBsv
sd+Ler9QKJtQyxBnKUZIkoITh9BINuDXJzuYVOqn0v1xHg2+JvpC0bhf4nMxgH6q
kmxWKz0K7QoG7xW9YwZhrR65DFnYn1revcaTDg7FzuTzmTsGoUs8geg+qIyKeHoQ
470R5D9OdmnRwUMvV0HK3eMXQODKQgjxZPtQ70k4yHtpdo50mjiW0vCxWF3EXnHF
sSGuO0d193w5Xp2aAW/8wWY9vvl4rMKHedy5UCxoQlmkQuR3Jo6JN7cxKfhS2q/W
49lZaFvmgIYywJDRgXnWKRvnijXq2jSMB87Fl9241SqCWN0jufbnaiDGmFXjcHor
mjCCAWHCh6oXOPK6vVj+njvwYe6rkAbESXsQHBTEe8gPEbzbtVRNQny6lpZGUpJr
jJw/f2cfT6yEB0QRWQsTmju1p+OFFpDkmn5DKKqDTcHrh0HecBE4ScgHkuB0RIya
vTfCXncrIjPG8Ri0w5+ZSP14FJyEcxABG+DDLAKkW/BTQlzP78IrEjxD71SvlmNj
OpZt5oi0cQmBPpvBZOPAde8v3hjHxhOnHmcBwJEIh6tbUkGQi6EOqab0nb+hSsxc
c33dj9jSs+jI0kzTfDbYHeLYIKITzK+0yQi8VfZLU+FPA3en3xT48N7z9W1r5ZfJ
eWQworQEcSeMcgQCLUvzWwMDM+8YEcXXwNFaL6TmNib3PDqYlril6KdyeCPflyfs
OD+rnME1wcPUE4H28M7Oeh4C3j3EcKE3BL4kjaTJZYjiN+b0DIUWrU/9MNsn3cVW
6gS5j4Dv+CbWBjLfzR13aAki+J8zkTiKR+98khLmd7QWe1QVnwvszKNUMxc7+3Io
70ccH9nHYvL4tK0J8s6copJ1zdCQQ5KjKzac1/rvbxZTEvMAR6f90zzwNcGIn2AU
E2xhr27SA+nKsLpS5r3Eaq7+YPYXyd1OT+ZbJ9j5B3ayfWxGFZM1pvSKrFvY5XWS
vW5AXeqRbp+PxT+tKqDeckeXRiREC28vjYE32Wd/aDRt8wLBrwEfX3iHu2xBzSwA
ry2Btk10MlQJcEeMPyn1rSdG1VbTxwL9Tj/D6blHjikpwwYB7L00s8/HMRw5oN4z
OqeqnP0NSxB3z6o/sNf4KUjQPDW0eDA3knt7kOn7JGADbUBscD0r9uO5hDCIXKLk
gM8ijfBSAJrdfEuMU0dRtOkPr46IO1ZHm3fg4iZe+RmZCBDCcBXye+Ac9Iu/Ql4/
r0mX9k11DI1k0XpF+59/nEDpTpoQyFNB0ClNKNqwfW2aw8elDkWVqh25vaTHJyNv
ElmzdhZ62HM/s8lEqWAIpS4Uxyvw+dRpjGX4r2/mcufBrmFA6/i2Yxds5aKeZlLV
JKh75178qkbBrI5hiiEuVgX8jj4m1gF/4SFh39MgBdJTTtCry2abuY7StN2ZNdO+
iQKTTONH+n17PjKg/+E0punJVtEItdoa8t6esNa019hQr+koTwYccbHiD0K5RF7l
W6Vjh5uc0KgBmZI18m7+dXDGpnCDbu0Y+skYoYLt/unTwM5M4yNVNZZnFYHxkAl+
NOv/+ccPLMrh8t+rlLgquKzwNhQrul9XlnC9l32mflT1zKFBaJDA6VzXJRASjEMX
jag4RcdleG1UqCBn0CIfPHPKy0vIhxw14v3lNBkiH52ckdPkOi8Pu40Z1TkShnwS
3PFTMxn1zEkw+do52mznD0Ko5FiABWZs2pVMonR0KOU76P1ViuGKWINJ84jStR8N
6NHwYytMoa4QJSha2359d72HW6rQLrxvZF1APAxsG9OtPGKY/B1IVnQzpaK45QV6
T6a7LE1YM8vtmaPlOkvqwmERJQHnYQGsP6kjtEO4xCb5aeZC2j5zPRgATeM+W020
UNiMhA2em9xQ6EZzfy+/JzDtyL69eioqzGLwW+Nw/QNkVTmT8TM5555WLCuIZo9C
lyo6WgysVL4ND8/Xivad4fsw6AWIi0pZx6YctuIV2eQo1swrI8H7nHLwij3gSBAZ
riuV4onAE0hdMMN0NvPYOBjQtqkjzLMl2fmfZtEVlUp/qS5xnxUI9hSHn364H7vM
l61h6z5504z4mHBWe3MleEatIhLDBwY+nMYh1IgaWfB9TwxfB3yMHl/OSRKjdR5f
pEyzh2PxFKiArvOGSzpNISdak80Qxx1dkvSMCCOKJHepsIMp4krDip6kas7xPnvV
2G17nJDOcQ1F+UIsNVuzmf8zt7/i1D7A9clqYEbYnvxl2h7W0OqmGqN3aPWre7Zg
pmpctabr2PFp15aXSQSEGhQoNGon4N2apBr5re6YrH8yksIkfcDVBbGw3MuCRUIf
47pMmbYtNPYdenekjDMpHTMrwyrcwEBZDQbR8GIAW2TGeGv8h8CfOZ4d/K/Vt8A/
cFqh8PYwv0f+ilqXqgptWCZL9/Y3c/8vKgsTO52j/Y0abFbmViHEcwd8J/mCGD+D
rJifPYJVDCdoe/WdXSQ7a0KkCCWGnp/X0zvr7Le4mUVy9E7vRHO3eQznFc+8t4ly
/qtOzxn53GEqqVQ/yDCBSkjbnAGcG66TJP3V/o52m8/kOFDP1sY8uSueLYj898oM
lsb3jhVu1r5fwHmHt1NYb4sdI3ta7c2eIqcY/w58oR+/Vs/ivx+oLxmNFKjZyqfO
0S7dLpDNpx2EM0uaesgLN1uXi0WKzhUj04ric0vYmJCT/NvjzXLSdGmXNuNnimP+
X1X9uu+CzDyokhza+vvTOOPDq7VkVZdXkqT1OU7dMRSJCgUqOQNeAGW9KHa5Jrwz
Ql4WiZTJinsGHTy8TIr/tUDqUH8wcfr4K9cfiU2I0aaZNBodLfNHJSt+HHHhnlXV
7I68zl9+RZzRVeGwPbamQWl2CmukCVrUWwt7YUCTvzhPcSilZo06IYAxpYfE/d/4
oLAWxxhc6Qm+WUk9Xrd3HrS3YjQJ33488/GK2TganEpmFbf8zDVvhpi37mWp5sj4
Id3ligTJM7INGd+rJvZfqOnOkbyz7vepjzIFDCZ88vi2+SbnBeoDjTnfIA0Cogh/
DxRHDrGQ32MiNYnz7Hew9Pd2QHx5D9yU2VyW7eEApUFvaGePP4Kx3zmQM90aPnnz
eMdhWn+mqR9IVurKoBL8rHaFJhji1ZhvXLoOEfzAxqJS7S8mQq9BYzvWXoC72ndf
LaIprjZCcHjtwhPRWdeuDRt8Sj8Vvb9l1RQ2QILpxuB6SNX7cpEA4FBYAyMVNIGX
jn+1kREsD8v4plpxdYB6tNtlfX1A8wo0TWrzgXo2D3i2qJsryhXPZYosZpCNXryS
Opo5GSlh12JsaCZXbeO5TK3q42ys0i7nCRCRdLEX+j+gjRoWORCpwfdFpAysC9w8
pW9PbfpmaMD0dADhm2xZRw4f2T2HYg51OF1I0vKepr4=
`protect END_PROTECTED
