`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YtkI9/GbbtIlFS+RwiSIbPhgnPpbp9HkPbUyeqVYp/j8H96m5dVSbpU4rJuQADhW
qJeGodfnJmvsD9EVgEHmnVVPTTAqjR8CjLsQSqpBEeqGZVm0SMPQMoJv8x9UFZWJ
rBHpjzG/3SPnGVNmBEsr9ISKJtt7WJEEGB6lRRq38ur/Qg85TcGvpSALgpYrh9t6
hZS5we60OBOQDJiJCvDLj/GV62/UL08UqMzTnmQTIPCQQ48fCkTy+r+xvlvs3lo7
6j+YxajfEDkjQZnd7uuG84Ct5vw0WY+jLm9/nfKlXH027/AFa8oTTh/QCLuQKSJI
wCca5W0n0KKwXWso3MdtvgWnNJH/hyvdSrptEIPllxMxeiQV8bafx/BFKNVQ4670
a26TKMPtcf31YrPXlT7j7RDwj/MJqftxgzjZZ15GNWMh/U/BuT1P8uK+CYS0+B0o
UrePWgJXYEzO4Pf8mCF3glh977CBM3OpUAYScir4baq0eUTcne9hOcZd/dWl99dt
XqVgpyGf76eQpVcT/fCS59C/TKvz0FqLv/j6Pvx+qyyKkZnL1dKy61YIwJlXl4WE
IjUlrN4umlaB95nHl7m8UrB/sO+Lj4YQ4gf9DD16w4fVw9St4KAqMgEiYw24CuL1
BhKA5FJG7upcALHQq0S+yxdk+/dguQqVMMaRMAvq30GoY2A96P7fmUQQBRcJ7k3v
YApaJcqlZucyDUG6/FlkmZ+Uc65N1jvAu6jNUDqT5nA4bShNhdHTBkxQpUdAS1Ll
+6MVciZC71R+S6AntQhFD50/I/4BklCqBtWi3xJB7Lr0yhiWFm/jBgKqCY3n4der
WyzklsQ4rjE3S2Mr/5pa7k2XLfoT9OLPE/h8TEQfpJAQEc72S85SVdjS/wp+5dNy
HtLQNZs0KHM1LpsVxOH3F6Gx6qoYEdgt/Ok+Qf/yiIXIEKm2pWm2M2V4uUp3KICq
RMy1kJo9ONiJJ8F5xybjW8yyKddTF7cqrJHDLicO9BiIahstLan0Ypi1xxE1maMq
K1DCllfjdWgQnITf/94pFYbZ78q1T7K8K0FLzAt0vLWDQru6dIu/pyuKEZeEWZv7
WaGtXGKV5iTx/wXA8tCqgVE9RlfxvT1I/8yi9m4fI5anqASXpNcaZXir/CCLOnyk
lzC/h7RSFMi8PiKPU1Js/h8uyxSLh8Mp146FTBHJK9HdaFGA0g6mWZEX5SUp0BiG
gZsYQjfIl11640mTQz74yQ/NhNbz9GvdUpjdw+KWnT0D702+MNxL/MlwfdLdhk+8
7igyicWeidGkUYhjn2Ga3dTYPauZI9zO14kGkq42ZpvRreadBPD6KojY8isvZ84v
8l3h9J3YBcI6IUXebcqgOGwMrISPPWldsIjJzosXxkRiWFvYPrT1zQrgoSZ34iG8
f3DLd2eabs3ptBn1bZJ3Kqo4PBd4vNVRVcOu3BkzJa/KT1YGfGO1ScmStnDIqgUE
g8aZUGvEyTCtbSefv8p0XINqH2pXC1sH52E2x/uU4T+PwUd9QkOl9V+6YfOqeDSd
ZIlXYTrm2vLi8QKo7xYSQMpDaOwU/54aX/Kgh/DBxzdDrhV1onKTXBOlvPb0DI9a
GHBohMZ9PFRdbmpHRcFl0xTb3BX8Brn9y7czUYBb29l0JNwjdAyrZXT6sFKJUs4f
GDvOYTF7A30lJNB4f3VGKyu1c8NDFu+/pFS8Wns3rMEKqMr/oG49GKnEnhE9vc8l
L39UK3pTjS0XTDeZ+9ubQ5kCQG/uJ+0qg8/Q5OE9krboHbc1q51BT5XHbz57BosL
wTU9FRjcmtAh4Q2UEIGoURet5Ozq9bHXcEEg9OjRlfUQaLSy8StNJwsSw1Y4XMnI
n5fsXAJHIIMpLRZc3WQFvKvkAR2Z4K345wseOrHmoLWsFgZUz93Jrl1m3mJR745N
uKytRlDqHuT70ZzJmHoAxeOj6Kc5KJZakFb2YbU1dzSNHGPX2xLMgRl8nov4fstV
PwApBo0CeC1b0I9Ng/bzThRUNwvnu3hjOxJ2s7HrSIXPXGwosL9M+E4/weBY+MW5
KUE/5UfucgfwGj6T2XDL5zHxGvMPusyLK34dXCNHQ8WjPCVmiDd4YeNLKAMzMMKm
`protect END_PROTECTED
