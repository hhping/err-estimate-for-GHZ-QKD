`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T++rsWVOW3sizpgnf+ma75rDBpX/BkWLAfUK6rgnTUYUr6Wgp6Oba2z55lYOK8XK
rbSfbg384beHZc++7RbWilYspGxF1M4q7g+mugBrXnvl1YqhQOazU9Gnutx/JYNm
aPzRbQrPTmjpoZnF2co9ficxJFTqexdiUB8gKwhGiPaAtmnXY4UfigjVOu3wrH+D
qXu9jPWmNB7/FzftCuQX2W4J07HJkH/xMqdrYAZfI4ZEXKRRgwJfzBfQDpvTfMWO
eY2vU3zaFY63V0+2vMjbl5Y6YjN1AC6inFml8woMfXRxyJgkVfb1cr1jtCYEwixG
dWgJgvC1pR9MNkF/DOV5YwMof+nD1pVmgcjvrMag358svDBRwvDibmdUe8JhwiVe
n6jr+Osyj/hzG3pMVstagCMq9eTKA8yGL6sQjSTJnqvC/2K9eXlmmtRXRxXjfZ2g
l4kMqZ0qa9gV95W6avgGkyloW2oRsu6o1AY7s+kkFCa3NozJ/2xTYu2pzNZ31gnb
o4i03b0IWXH35eycPWWlpGTzNQfycG+a42eyMaM9QMqKzRIzfHJi708J+DxECYic
euMJSo5NExwIrdMtJTC351biIw10dPEhn+cm9CK7JDIAD2NgbgIjsfFPCVbrjfFM
SP1aAfJmXBQ0yMxaV4J/AufYg9igvFfxEF/GHbo53dFlXbFkHsk8LUjJ3rn7eu63
UZBo0nyNLduvOR089dl4s1dh/umjoZ4K8cCq7Qi2zC9VGTxiHXXDUqzBiw9WrytU
w/gUy4TXkJwaKiRtZzZmBQ1b8bmjWS9HST9LM+PutJaKkRtjExvwDniHJ0bROzlx
6nq3NKBOxc8NdLs36c1gxybZ9BmR2br2e+YtcIMXPjQ=
`protect END_PROTECTED
