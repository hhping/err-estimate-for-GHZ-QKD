`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gMD84kccv31BAyl6swmJ8LFcK1G0qEnNRoDtbvYAhsfm0gWSntPWdXIyYPgiMpKS
S05DCZqXja54Xz92jhJNSb5KptBSul4qIEf4z7eF4rItN2vPrAcNAbZ9+o2s/TAM
Tp8arZL6bRUl6MdfSnD8OUTNsactMohj1hwpHUF6Rhi+gCfPHf5dMbusaYsff8xH
VMBpDGJurcLwEVy81TJIMDVjjv7HGU15qu3WCB0BCodXsB1f6PkgQR/eMAW+K9yo
Zg142lUGE4C/3J/STWHV/JQzUq269FfpDESHtxZgVAngvVGR1fNutLpvyYjS4KQX
LvyXAu84wAB2JB/MNHgMkvE/O0QfGdfdn9v0ACGWil95a/ssf0Dp8soME35WyHqY
cHKR3NFHVmS3N3NrErfulDozjarLr4GNcwzjwZuOfHMfW0iUl8yE1q0fhA6LNW7i
f5sP3DiyPgIb7zPiKv1tqQ==
`protect END_PROTECTED
