`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QUPZ1Dk1QCiCRq5jUJe8zRYBl7ym5RrgfXSyrwd/BYJqeXncuk3DediYLahWDaUN
j8upRzfpTrvx6UosqFheYiaemxnuYu1C3HtfIbRaRAlk+D2RSQQdyMoQ7LuOysCZ
9iPqfvAZfr68kxFxPdfZtvJZfpTwb3jO/uI1LY6Jasiz4b9GaM871QgbQUeirFff
I8CwXPxFuT8yF4n58qqM9vQXH3Aw2in56c2W6Yt8scTRxL/LHnZ0tiAzBrpjvJDa
aQRAy+S6UE2A792OVcK/szb2cDyDYujz+ZBMRcYazJ4zxuiZK9+99LE6rycml+lN
GO4iGus3auTVN/x0dD78Eav2svPgIaGLbS4+fAJd8uIyTsN8KfrNn4419gI8bvtt
VuB302E4L+RefkKP1UbEb2DkMyrM6tsEvm2XPXKhjSRei2ZXiHKNtdS3si/8xM+a
HUvu/afKnALuX9gSO5xhFaNimx/gX4xaZqwOp4Adg+rnRz3H3bO+h06OJaht/9Cq
4Yo6a8WAF0bVW2oWcvZiQHiKbLuelItlSmgOEBVzZtTGBO7nX71800jXtpFS5Lbm
RcQ4pOt2t7c+8BQbqWBit+CmoE31rVVZyiioNE4njm81ZJEPzyK/6K1OaLicYiAN
mPevsSJg9/b2iG/lIle72U7P5EM5N9Iz+GvtKNzYOEiTlxnezgZOMO5+Q03xpeeA
weR75vELjZgXKQsWMokXHOCuM3sHCi5Es6t2ceMvL1usuyQr6c2eMGUi89qKVhdK
3B7GFTVHNGdCH1ZRJH0/dSt1pOB2lCwUP8lkHaQDAWaO2yDAvxfM2ImTSwUQaNic
puxRr46cPDOdExTHxXaDo52GdnWSdN2j5SJKPLXPxooxFZqkcQmeoTrhQjhR7LT3
ZkZ545GQ+wMt22/2L7XqMP9/JNyhy09iYpFokVTCf2Y3wq6OxB8vy4vQtgIOnjpZ
fLrMtx+qs4HHePL/9WXq7sQ7FIgQm2bcIbYEmxKYddnXqa8Jyudwt+AtRXyRBPq4
0kMfGuQIFECKw9epvR+7okcjswc+GufNsvbVXBUsWT3M0Kjo3GD5wl4Y3gDa9XCp
/KKKHtOwztK+j40pEFWUlWMCJwSyh21ui92C6QUgodsPDTOlTZUwLj36xKqisyWV
UATHAvFnqkjoz7gX+wG/sTLUzyrdgml/AcgDYwUymI8T5L2htNovMiLA24JbdwbB
m+p3fb4k0/5yqyGdd5MImns7vvVvCia6qEsHQjcPE2xB29ZkrHVLx+75mnp8DUeZ
nFYcADvwJzTASgpSb1ByKJoQDkNiLMMRv5wRQziB7ICF73G4+2QS60e/YLLzNE7v
0bmJJtXKQysqvxlufbtVhzB/FWRGwWqDYeiw+TH4nSPnS6yQ+y59aiRGjps2c1mJ
ML9VoGP8JgtEe3CDgRZkLtHh2Pm+c13fsAwZOlB0ccNQRP3sjOGvqBwtgTsPRUjh
`protect END_PROTECTED
