`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s+uloY2+K1nwg/32VZtUA+/aM+CXNXfGGPAonbOV5zP3OR4QmJ/IYtI+V+TacUru
rOi5mikr3dZTb/dxeM1XlIlh5fM91Rqi3+d+bxBpSIVcX6nnEN41JDqIWpquwNJS
eSZV3F6UVcEoYP9D26P6Be2cWwwuuNHYg1gVCruhzsiwBbUbE2tnInQE+NjS9k2B
XjCJ+KleT73iZ/FkjExpWu/hvxcvnqpe5m5bkjhFGs9PHApu3yyHJWjJZVAhtpnN
N0t2OYLV16HWsSxCvNFhpyycShvEXxfi/7JZCa7YwVQVNpDCXNaGv9dKJ4ZvUM5N
CTwGHdaIsIajRVFZnCDh6D6UtMurRg90OH/pxh7gux+lEDKefgHeFOtGzJtTavwO
Eqr6D8Zveeng0J2HXp7ujCBvI6Csd9KaEDh8xE61p3wjrSd4cYhy4KmKx/8EWMy/
WhlRLfdbUQeKEx66PJA31ZlD+2MTY395cdIxEBZvn4kI1I8CkuNVJDQbLUbm8HxU
PSM4YMUm5Uzs6kqcIc1dZlGzorR84S8b7evS+a/H1v5bki0kG33cXFcE4CpB0FPg
YWdik7wQdkGI66mcEmIZQraLf//rgEInQx78BwIKfvLCMIEHCciD26hL6xuRmGI/
rIEXJvbWbtTksuvbXisOmTGElMvyMLgDrcACmJ3yfjF40x9VBSSkI7HysjTJl2ZK
kpTJmoefMpKqPhEmoSTD3pkhP6U8f0ogXJpU7LEglhEQNgiv3LP09iamr2gDaD4C
BJBg52SBM/OSQ82IIPcCVylYejhvYcKfBKFMNvCgeR1POVTa5tn4YfiD+f+ozjzc
QkqfE+v4Tk8e1seoI3BrZY9HeTJIQBgIU58LAKF4qNEY7FdTVOMfNkmb6L+oWoDU
Cab2Xiaau9H1kNZj3csQZuR7btzR6DSItw1J8dK/710YeYPIHP8Q6FFRwZRUDlJ/
gnwY0OPm19if8av3J6FnWPLts5oGkjM89yzK0aP9L/ZwX0HDmmyjTu9ZHPz1AVoq
GUebJb/toUlMTLk71btMimH8QrNZxTWJvNLcyTgU+yn5hOleZB7vbvL3miI2+w6B
WC9N3YSv9s5Zgc9DWnXkqN/0fIoIQmnZ9qACKguy+VsMMr7vPriBch6Q7e+4hMyn
ULLDzU6rDCVHZjjtfKt87tKAV36L7n1Lbyu2psmZF5evCtVTCX2fYMw2JOuKeA00
sl81MM+RiiqvtqhbZsaLzgOgT/ZlobVhrThiUr9GGiq3A7DWI9SbqHoX1TpB9+LK
/am8Wft25tp0AGBcnshtMMKhlpUtfKtJg5I1RmIAuiVbpTpULXKSjT+C64QqIaQh
zu21Cte4BkLYmsLHY8z5bQ==
`protect END_PROTECTED
