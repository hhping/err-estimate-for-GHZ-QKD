`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pozkqLJTaK8nKv036n63JkP5XRklI2e0zXHNd1k02pleSCgQmbrv6PXzyP+oymxV
E93AmoWDqt0LZPIs0xyb1aNh8YTJ2xCgztVXiS4YX0KTqx/pRkM4FpP7WM9OhXOS
fAJzqjosrdxhjwtw8hjyM9gZ6C++B3ONKTm6jjlgZEX8uMm1mu9VSDSo32kmSsaf
k4hVmbjiszxgyR14yk7Ob4mSoolDszr5CAvI8LOFfg8CsjHgHY54wLxly2CISH9c
WAUk0kyXT6cesK/uDnl4zqbSUEiELYnAa1jtWYbnjOsYiVXV4m9nmZyxw6c/Bp9Y
XHD8v8dymFY87x4kqKsYcG9YPt2olJPGrTm6+5qnUkvLrmpGTQZboIZgsi21wt43
lmfsdgsBceyx7u2oYdUeMXV+2MvAsTcBz6YvDZuQog9R6z56pkUuk8XJHRmXf10n
wHhtbUbpCMDCBexsv0CJasH5Zytfj1FKRaY+c5D1BX60tmckhucIPCjga5IHoUmv
Qu5uMAntdj0LF+tISGrxXPLc1/JxwSm7K7K2jl4nvYpz3pU8KFDOB+7+HxeEHwM4
iBZVp/dQBakKxrEMJgFthbxgHVg5Gq9vgLhH4dbTWR2hjkwIGa4aFKPnmD9LRgpW
599tmkh88+g9MPdVORGuQN+ei1auOx5qN3DHqTRqOWhE4EvDCwIg+FLhhC5Lsdwm
Cbd+cFhCsKzBRXGU7+nA9IP90qUMZvNajAPraJmL/2D6Xt805TbM5bvCYzhMJwl0
XT7UD+3SpGJVWFEyqfI73WT43FP2q9kSABQmpkPmKCNW/HHKEF8zI+B7QiniqJr/
hX29YKBhkl+Iad1W/7XaxnFhOZrTjKhhIQ97yzjnUuq4ciMwp05bb9Q9C81uScJQ
qRIWH//DJroAuX8Z/5O/uILTnhZrPFav//lWQx0bIQVmqiHjGAafc9+O6ZQ9OjnS
kjrPYJdeEdthCzJQhO3oFHFH3wo8a4eQ6+rWaQ2vFXo4tN5Nm/8tLJv1Y+rUpa4f
dHNM6zjzb6UcwyhKonBbwyl+TXIXT4cle4umKZ5TxjTFPmPaYD0hmSnHMJ79Laoc
JD4glCGrPDhonWggpVTdD9pUquR2IdMcx8eFKmn1cv68m2rc5FYNGuwGty6wsMk7
RyUNuB5x/18mHIs8kuPe2C6jH1zwW2zKTsROPI+EMc21vWu+WClwM137LsKJ0Ry1
52wYg36I5HiBeTI97O1BVgZQuKd/qkr8sMVl22cpRNU=
`protect END_PROTECTED
