`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dH9+8h9bNHKeAYvYBC+n+sr2tf92IsFU/d1gOyUPcYNdebyW+UbN5phABLzZnDM8
dvX3UoeNFWSAjVztrgpqW8j5PvL3+Wa+Mr0m1k/JLXWkQbLFMorvWlnjsiyWHrr9
tK5QePS/S48rt84L+JSpVMX2CAa0JIhZBypWBavmhbiJ0UYqHx60VO9Y+50qmiDQ
xQEl+TuBciCD1Uqxt89BM0RqJ7HS1MDwEuYWTvkvK37qnz2t7utR/EMBT6w+rNM4
ldN1AslKjR2XvacwynLLRPJUIoMDLa7uB23SzcWnV5NPFC4UcMGRwMKZehfosaVa
QqJIb3aQ6xLAWuAO8mlj+7wAhRYg5Hh/bUPdhprsWAqwWKkl2ljNNZGq4PKNQJqI
IAnCbaoVcwrd4Yovp5Y7IgZMdjUnSA0jrGAygCyPsS8wOqoPxNBfJ5B0xcv6sMHw
uBl9x0nXxcA+ozO4U7MURmMq1h8ChRGIxIJ4BXT2HJbZl2mVPScxUzU+uuMTcTyl
8do81uWZ22Iy1HafxfOHQCBaPIhXrIu+L7ISkOLVRzkLFGp/8MdAIrHiFvDVTPAH
IMcj5nUmtPC3mFyeiwkL3ry0ny8hbxuNQReGDBpj9Na9huNqIsVDwlDMxZ/njut4
oRwIOB8WqS5ehssi0J4PKOvOltUkxA4z79evwlmbETMOO4o7v+H1/V2nCugMDKkq
kK+98Fk1UhFdQ5GFVKyqrtAtF02mUKBKZuwprxUsy8BtodVzTstlKasP1dCA9dBx
+es8QjwQCCTGRKyGuHrFAiD/F374OhaLuLR2JhobU7XsfuBKPjSl7D0i19jOW8a+
YJ4RJhgaX89JoBkPdFRPAvuXED67RSEsfwEHc3u/S5VGOh3hvaxIZTiS6i0MTqai
gtgAgRdMkrgvQ0VTVzvdsoIovZ0TfxZRdSrZSHTiOu7Tyjrxdki1PrW+eUY3mfjb
s6O5oNiQh/93YTWN+M2h72HyNnL8tIx05eruawUvHkAyGDbioq8MfYw2ZpYjNCiX
Mrm6lZ0H5kcMsOdf3XED4HVv/FgW4oFJhoTAjvh59y1IkyU+Bq/9af6j7AWv6XPW
J8a+/55y4ece0EgfNlLpehwPb5W/0O+HMa/1VnkYZQqkVKu8dZ2tM5TR9tmSZOaZ
Y5CHl6xXxwQfFum0CEOMjgBYMXpYZy9d2lBQ2hxyRLdS+Go7abUBXUVf2mEN1krC
lZQysQ2oDwoSEs3HDM0yGxEkgICUZJtmZxKjP6ZWGORhPKLxk2GAVX9VPEvZhDcZ
OQRF5KTdS9Wcl4k16NCxkdMucUC062dTLR7s+jWA+3cDC4/zjxS/onkqtVxPaUdd
5Zb7FKujqo6l6CJQARQfgOHdrj0uiBKoNnoL2EwjpjY5vLK7IG0jEP/WMYh4CibO
0moT1gH8kC+JwvGnZxDWNLA61M6oCgZMbo52RPUm6CrHIrwkfy7iMd2klBjyb4sS
yZesfdq1hWD6FsK7U1mwDpVQX5eQjwglyvRhgBYk4cr9hsZDMuwrhWZa6rQPZdkK
04I4q2p4GYDAr4rDYsU5X3FCGL6DpB/SZz/zwmnTHz8koYswqys20ysPWVeGccJS
TGIqBx7XrqdHVOfqaPs4DJ0wn6Hrqqi038rgT/EhirM=
`protect END_PROTECTED
