`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EXbsugdGzihEZ08F+ewk4+8NQBk4P3bc5qo3GIgrH+990Gvmle3UfyW4zNZ5O80j
AvhdIjIx7vNzx1iqqAo2pnCBYkI2/2PZ6U6G7F8n3ds0R3U3IJO729RatsN7cGoP
TZffwok3FKaEuDEdQk8jttpUKi+v3ETre60XpHMoMZQr3xs715KA44/U4cH5L5C3
MJisVnUvSdaCu6QB9/ATexJcs9HpVheWE154aFnVp0K0WSEqhLrWn5SJlfrXugsx
1BikTrzAolE85sXQVRscYziR2wm59On9blKthR7E3zqcdVHYXn3QTJp7pt6zIsS5
hb4amJA/8JJQdTL6/2dWoJ08MeJ6wdYebDSRj2r94KvZ+XMlK98k4qRM9cMH8bE+
+CNleReuu2mc6W0RznJcrX0C47FBtG9zYHPdETfFG89PdXQFLrJko8mq3GYhpXcM
uDGgMPRF8kz4smcD8OBM0UVch58I6kAQT4vfLWAAjFwHzyj4dn6TGb7hBdzF8riG
qHVd37BodVsF+HhoP1VIl6wgemkeQ9MBjyg1P3g0bTuFIJOVogiqr+BniuxBB7GY
iCKNtO8XT25NwzsWj/P608ZXH3KS4F2vsSH8wcNovGhJVA2epGpIu11j3g5AeNzc
kfdNgAJsWQ+GMTSBVTeBNydxJdaeAux5R6hsVcemUgLdEaZ6vcyoD+Q5BGJQ2ljq
//ZeFe3FwVRZwj46mzQKBrki7fdx7RUQ+XuE/k1PlN63UrCKPajr7r/1aqqHa4Jx
G9A24WX6sqxlVytLuASnzQ1Gf1P9BystIR18osbKbxJtzrwGEPRybrZJNi3Z9PUG
3iCOa7bD+j2ZVjWgvz/lKE122TqmMYUq/px8gsZSwQhn8t3PjBVlXMzI+HotSCtE
L2d5nwRQlxPqdfEF84ihjjJ6wz3IW69bR2+QRvNT/F5HAe9/91ERtVOptaKc54Uh
ZTHxhE0Y4nuCFcFCF7xwEbAEaaxSU1F3K4d5H2MktUGKfg7VYTrkafn+eFOT0L7Q
xreZU5aRNhk1gDxFf0TyR2RMBsa52OWcQUA7WjQIhskHFxMiOb/SxBT5WFg2+Rsb
M2NW8g/ytpX/MZ1WIvQDWB4q6vYV5N1mRgNPz+8NBtA5ZC6dXKxKE0PTi06HsBFW
dQ4fL8QMCliQgVaY7N4UgHcCDlmKLmPZ2P6tuYL3VnVfb+JVCwpK7C+l1Or7EgVI
4R0YxOvmGWOfC6C9VylXEh+IL3ougVjPJEeVfdHPgBaeeLIKa6tqqDsncP0CoEp9
An/6fLqUgyHQ6FbKcp6vpz9WLvYIOOrASCDxoGlG6Whl0NTrmKD38YmvQfkByjvg
XBge9fK9n1TOb2/XXMgR35Mh0ob7IxEDaqL0tBM9kK0BkJPWiMm3ikCexmof30t5
MDz5V5J1sHXihpidN2AucTrBELGlDnf2ZzBSmMCukmK5AXHleBmiYxrVOdjB5Rei
ti6FXOYRZvg/Sw32Zk62vkUUY51mbw/D1Mdim+CAOt+e7J863YRblk6SCNp7Zipr
1jNrkrHUWe67n1Y6Pn6X1VRxHxWcZwVMKszz6nmOoUiQhx7PT0rdAMIP9fTsiKT2
MkngITTb98P9YRgXcPPYlMc3/xzsqTX5buHFl17txmc0DkAzrNCrS1vQaY6h9b6E
KBbzgUYr8lQOe7alt2qyD8B0lGda0Qd52G0JR130eR/MNWPE6ieSLBCZnd1iJIdH
odDQ2Zn8pM9e4ZkF8XGIb3Q6UB+xUFvkvIkRjxncGprymWe0CDs/4MiFqPPQhB2D
XqcIGND6fqPS8JHnv4flIBbyvVQZHFqXphrWSMwUrSzp6UpaBqV949Sjzz+JzaUx
7TSEyCJPeTwgaI2VhYB+YFD55JaH5fx/3fJESr5HLvqZMjXY7HwfRQ0OnL2HOTO9
q/BcOlvWzBvxRp0IrHOXZHuZAAQKlEaE9kAQ9/As4DOX8lmlYM+GJXs4VDzqI7MH
tG+aMn5VXQ+mKiq8+Xsr4ZuGMMHUH7ueVXse70uQueqqU31QHgUZ+3d926Lu9+lX
kafuNRT9fkS8WDO9u7joBCVm9r+rHyA6HGe8vSdOXmxqJJ5wmPaClg/HqDD50xiZ
nRvik2913XXe05NPH8glip9GlkrzIc0ze4qo+JNTfSEc8yOoFCtCebHH1iv2dAps
cdlKX89QDuSZllsgpaOrv3ZUe8lx7qQggEZl/Q9nd1BWhWnDtH0q1Czs/9GzA+Gg
iX6pPGtYdN9RhDh0uwsuyYdOL73HAyINf3pd0Kpooc9hn7yKTp8gW8yRd6+9HrGK
f8Y4+Qyt/KGqN6Jux8uylagySV/1AklqKFGgbqTEgLSFBeCAlAejc3nTcKX+jAEv
UJ88eccm6cXo96wJMYZHmcez0g0wOnFy8COpPSa51NJedZvMqFQ5NwcYz18IOZgN
Lm1Gorlxrtmsnc6+17p9fOCiaywtWcCsh3+NwJwih7XmfA1HluBCMavAfXf9GSmH
urVQ5NzoFn7ohNoV8nCbJJPEFz23jubkbGGBAq7RoYFdZ62sE56N5o4329KFrXQ6
x0al+efA3fTe8XTFgAmmH57JzU99rm4S4/P3icz6TQQoLdCUfIRG4yTKeM8Lftdx
UUWY77gJhV9bFGMLd0ID7bnULguVmfEAcPpoaYi+3Co6j8q8lFGYFA65HgCma/3v
tpx9m7HH/a6n6kNvIFmNqoLO5iFZ0iq4G4PIXWQvdXZE10YUd9wzXCDL+CA/89ai
LmS3PA6BApq+tdP387HSQyHIlEaQ2LtWTKsHHExOEM8FLABWun5AGrOvPqLRFX3m
vq9YOsJrjd3l9eK+1tT4P6xS4/0eTqppQjJeYowZQKXtpd80ULGAoZzyjc8bNead
WmYV8e0dwRTO+WWX1nxogrpf5H7i4EQA4zFLL8+TIDfc6XfaF4gCAIbh1zgStqy3
UwVfIsMkK1aorwXWIStJUCVPTBcgU0N12+6/KaRNWQxEVr4A4hm/LR5qqm0yZ15t
wvG8mAvu9FGcs6xumBASCfMJySTA41ZC8JVL+OouyNWZhh4Wp33BDEAwu4lkMwbA
w9dx5irHPnfJndXyZas0Cze+Q5FloNin7Ppx+fg2P55cCsb4Oz22hlMPKGwBDwbk
PmR0Z0GOsm2sJHN3XyOXk21xIEhA9cxPyeP/tf3nI5XK1mMtPXj8zGSHkDKRiSL1
AiBDmwygHJyZKmD6T2HcKtQqLGyrEMSABhWx+tVLMqfRBjtaLJ5oAiR0qXqWgIZE
KLRfBvmA64nGtyK7KYa+kHySdq/E6BNXiQGH/XONsVIJMYHD+QGJ90gH09pK8A8o
MAFPXX47GT3dVDWYWXbyn2ZQNBfU9QuzEZ8Gjo1UxZyJLWvRIcdE2FgQqwF/2jpN
f/8grmcA4SGxEmvS+sVu0eq7Mbz5cIED4gyekCmjPMlzyswkP1iuomlnntaQTNOQ
RjpH6GYougAu3fH+yFDSXXmRnZFiLEPU3FITmrMGfAvJiu9+S2DnoXeJzug1+Xma
NZpomkh1hBE9eJJ+27inRRUrtxkAY8sKOqweIE4iB6jheC3O1bC4CTEMuBGK4Eix
yybmij2WiWdDzpAUAx213DNpPhTgSOKqCo+42epgYydzY/btxK1XsYoSgcxCQnDf
7TK/cKX+nBWKNXFQjAe/kRLlQaVZ0CdDsKmce9DRt/Xi3KFC4+7vZaaaHCIGUQ+k
Dd9OirqwIJASS5CAFP0k8u6uAc7Et9f1b+cwEYacY5Ud3Px8m+TqbundL6pb3Jdn
j7XGql+NFdlnQ4RIZy46Lf2M2+15unZFm6/yynEfQ1PJHdAOEgktfbCGLBo9Ii0k
CyN/Fe5OXKB1sw6WJDt5lS2um1QgcEkMzYQcWLNgWfcp20pGHremZ9LIacYYKMde
YU+o+LqW5PW2Yf5bsGdcCOZdvO0DBkBjXxnZneSAdlHZxwHaPyLzdVxi6o0U64Yc
13VLg4iwv0twVglRrsO4+nNBcw4u6v3NS4AG+psOKZIPsd0GjLB6o7lKo5b3Ck3C
Bj8RR6bsOFGRDz8C3zgNHN6I2CmHxec5vNEpTsooJTFGK/f4AlFwVDGJbhRCBNHq
HABi15c4XIjT5dcPIduss7vYZkJo9blpr97vgOVwgXoDr/KGfkQASQoX19zef/5l
Tv4Dw65rDADsXR0i4VxwqODX8d+ExnsKd+pJK+brcOHKbomI+KBtjSJJblDf3lGk
MSr/Z3ktNm/vMmGI4fsDnmbExqeIThfrLtkPtwtrwGXIc8itH0eDaFGONLZrfg/j
3sIEcT0qYts8tGYx3pmrSWa3GQ7ZviNMp36bl//WFRRPgaxmhubPE6NNHt26wesA
3gp1Z/j35osgW7mXHRl0etYgmpTlVetXfdaHu5ASwGQVJ9IImEkrhU0gYqJE85Yu
ReWUVs79f8bOccMa+rM046LnYJezCVM1B0tYgn1nmYblx6dasbPW2EFI2nchFXFt
iDc/uRL9OaCZKHt3HdaJctQHJWkUUg/3zt22+C2D1ZFH/yPLOoB6HFUjUMkfrzH4
p/ITk/s1vEpBMC1l7nAQWs3NMDdW9goLzYRvc15hyiJVvlv9A0jmpV8ZKoTHeKsf
g8qbLo+fES3LIBoKDk7csMo9jL7bYVXJ6bjgX4oEKYrKwWeWHmjk/Jk41VSlxqUg
XhBK68nHk/a+fP5XXmd4IApVdG2ZuYQRipPwJHmDfjdr2fNQcQ4zqGrjfCWRDIW6
a+1iJjrOk44J7AAt1qKpmZGb4xaDOPh2P2rAV8S2RzltiD1NiXkXelLfpxAIzFBM
9I6GD5D9lqF07tLDAbmMavNfPRvTh0LSmucpryDE/0id8U/Sg0LPERyytbiBzX+4
JoyilRt6fDLuJR8gsNHIO44F7etPw6oyqsgQhgSUwJPLCcreYGZLkZ7ntScvj3gz
ee4oNrCnKRE+0K17ibRq0ZXRdCvMrm7Xc5WLL7a3keeSvADReoEzuSiEXwaBLg85
0WMpoUpe164FAokjax6au2UVOd8HRx6R3SKzT20orqaOV8Z61cDyzByiUjAHQd3U
xE8r/U768md8z3jcWgOPD8v6EDG4WbRa5nvBpmTZR8kCzUdfA8rcHBqdH7irNPYM
vWR0zAVODMG+e8LHKHTy1GoPoFF9wBO73nbCYp/hwLy3y8JwvvnRYo246b5ZFwVJ
n76rAQ72soWOwtvBoywGANJiJN2ilDMIHrCQtrYvEZ3+0iy9kvZ3VHWIReBrKUjV
tKCORr3/NynazqzRxJuPE3EAVYegmxKGhXLaE8spiKIlj7bPUjDUy44Bv6Zb1BCZ
DCTF9+KJQT+/v/gW1oNhGXM+kB8KASjKvVMRTvbOw5AnTdwqJZvT8lpsX5XfpF7x
VHAaCQZt3SI1wh3BhdSCMIFWpeao2WJ0knp4/kBJX4giR+1cNjtLnkhkT2g7SbWH
uKEjvXCGEK55OSx+bFuft3+ZazrfOhy4gSEAu6iTApWB7AOBz6z91PxaX5Y6zbJC
jfTqXgpKzAxluDuTPxlfBcjLRuY/mqed99niBLbBFzzHlPLskfoDIJnA2unz5+Ya
dk87LV3aaRyJNWh33hN04W/SZdzVDHnIExP9FSjaPvMQoIfzRK5Pj6eXaBfGaXXc
jV2wJ9jHqTnmhox9DuvfgmS15lLG5w6Z5sjubbc7CE4HTBw+OYfOO43dtQ67s9Fy
+NP0eB6f+tY3Gzlgq5PT091jqVC4lFuI+5flO6KHCe/eXhHW9Yc1Blrzze4EFIpS
//7+uq+GsLts5h0kdl3mgXXjNKIMu7G7F5BPRRXsDq/sn2LD3qI97DHCvj3gbhRt
2R1iVh7sWiBEw1uHki9rHnNbogBm+mMyX2RNj9MJmzRUKlk8nR/rwsMSna3SYTDI
nUikhJ9WMCEIWg7XMs/OPcuIBmGerJg1qPAolxIpJrhy5MuHaWJWLMl1Nn4MkPme
udREMt+IERn8ObYTXI2sscX7p4d5pUrrDRpG8zX1pU94Hv+tgxY1Tjfy3cz/oNhM
DXENlrKCIbX7PrgurtgQE+STC9PpjCPP0u5A/+yFxtYLpvplGLRPgT1whlJHdChp
qdS0wHAfHSVqC592zQuCljd58V8DoDR+O7gsItryZ5oHs3qfO7zpK+xcD7cLSYGw
zXCqSxsMjQCF8PocZoDZtACTP0Hh9/4iEL9ojD8smL3/TjN9DjtVh0Nw3ZK6N0MK
cOSmFQ9yKqEWU0pNXAkNPkyFa4NgN6gVW65Zcs6huPsTKXoXsB7zfFVaZTZ2WLhs
0cOWwXa0UPpGTGOksZSuEYUc43fLYlNbXP6UlUjiGCsup5qXXGMUdZxRXZz8Pvdw
tLbR1rviQAwFxG1K0z/brrVLnTC8H/i1aM/nfv7AS4lPx32FXE70c/OJjjwJqmk1
SBM2OInJPMSOB3ahNIdWnJuAKyLtTd3DB7tWkREu3i2r4tFtUnkT7etyDrXp3k3m
mak0/2aBWXEyychaTvl2ZmC0FgzYioWbK7vH9rMQhlGCKEtUtk7T+18dkuFcN4JB
sa7xznIEgcpPks7fRNkZC6n00axVQi4CX52IdhmwIMyDtEG4uCpFvc3UzMDW7qrN
HlgZICF1xdGqXGYCp3VypDdrYD/ekTr5FrBXdYGXvfxV7QfZiJYb2NppHCwMevCi
zBs35FwMcg7T3XiEaMgTE0CO6FP2gUICeEnSyXCOTlcuWTvpXPGhcH5RA00KbDXy
vWEHs/hCF/man4tW8gJCzOV/+fpTvW9dXzzAjfO/JOj3Vy5zulNw2cmGJl6V1voe
740L9UV9YT0CnBKHgARD0AGy+J5OVN3OhHcK+x4KXDSa2OHJy9yV7Twol3CXkR44
onWIqgCsC3oKZVyPLS9D/Wz84/8iGn7yl0J0kyVGiQz20jwO7KAWlZ2+rotLjLIw
3ZD/HlWulqQxHmvdjqsDV3CIQQ93oVNoXbIMr+BtjuNBSCA2vlXtWvT/zAm0R9cx
8z6J2yPNs2OYCRbVSab8U/W5DwNZB4DWWeFTPIWc2h2kezSMTvEJ7Fj+cxRubeER
KeoFQDYXxTfNVhCmDYuK3pJe95sRB+WEP0KJNU3ruHWk/Ndnde85Czj0z5CfhMLE
BtSIoIt6L3N7WTMLwbOiQRJiBIwSVFYhmXC0toodpKKLP/yZr6/Ue19LBr6QCo8y
1EMQk+lczXMkHOWNP02Prp9VpGqSWArJs1AajovTYG1h1RQKChgcZrJUlQKl3Rsg
u4f/crEj2NllTifp3rkgMyTVIPt/R8hoFqKQH3UfhN+40vIOqb22HHbcDNlD8MOa
nZuoXpjxCc/caGne3fzmwUL9zOeZOOpN2luzDa/TVqnyw1BPuRx1quwOxvQb/5pp
VCg+vyWaJNLVaSw8yxN3KsGeKOaxOtzifG0Zhd7RKt4mNOQ6F1VP71cEX7UvLvCz
yxIyIANsm5nOFgcbPJ5IubCz1ZU8KvYoHUcIcGmZu7LGNa9xAAuvUJoIk9cPMkYd
35kFmEEjiCOYG0j4s78GHjM3t8Y48/F04nGSuPVR4w3dCtg0RAce1r8mA1NKZmg+
RoXOO8rXiQ4IX2z3m45cWDo9L3sEwgE6IXhBVPJxXSsNEYnF1RVLXQ3hfWjEqezi
8swpMcSOfArhYBXwiW9y2bUtTcFOx92axuJNv9Yy8cn37FicGeBq8s+DjZGte73V
2hcvcp6IFTPXLT7JOArRPV121RG2ZlNUJqe/2quxswBqzsc1exRTvSBCpi+/abc5
oMKkiHitsqJKzhRRnF643SLlNVv0l98zvGvFbS0oYDwjabL4rcFXL8MkdUG+nqPo
dKNvZmPiFJ+ti7YCGIFPSCQg8ELnP2a9qKnBmehOifQBY+ApxJlRxdQCmVCea+8X
yzW8tIdpyNoqcPLCwxWrwOZ8krYVOdZHgpoKs52e+1B9f1Qyfb3b5FZp1mddc3LK
GgD8dssweERujxiB+07OqUF232DpBONd3Y/oh0vXjLmDbS8IiXZVU7HX2KkbzOCv
aVQ8n0W6UQ2dy/1KMEvuSkiOIqYChSoZllQ+SpKV0axEOZ6SB6xb+T/WrIXvYTn0
mhjSPcSm27YoeEwL/5fAb1B5B45DWiijMjMbmT4vFHktMOVhfwyHbab6XeAkRtZI
LK5lO4DS6LreUQRmGopU8lR2VqfMUBcLmiyrGSPSLKEl8urclChTssPmHsBMQ6mC
OpSJPROoF3DCmg8fW3a/nRJSEI/os67jYEWS6TG1MUwH/fieSOyEfoHugmv8Om1N
xaLGWa1ZePAFRAt2UWZr0An2reoncnO0OdWm81i+KAb/UgPsS2bPytQpLhTku6/1
XMl1qbzrTiLfiskdheeie2dSXmGSSwDFEnTsP1WySeqQ2bSug+qeyGm1xUkICaj0
Rzg1H4bdotEyGAiOCr7eM6tUFXZ3leB0uUqq8Oqt1VtrPP5vOKD6ZErEeYCEKa3r
RW3hBi4BSz4xq1FIrKg1mXG1oFQQWLW/3WepIay0aYsUhl+mz1ahPsZ2DUAxkRqH
4MzWVUQ5EZErpG9T0m5V183ObZlWBA1+Za/xj9/gLauwsk3MHf7x6Mob3t+PcbNi
IBv3kxXH5K3nz2Xss0J+LMfwPGCyQ2ZCnmkUa4V+ZS3X8NBtitOGxog6TaKuIyY9
dQp0faagssOWkjfc2LcSru3+tAyYSgZOa5GXnUF7eg+4FZS+ER3d+xa7tJxvXPZc
8zVJwHloLnsWs1Mw2mk7lM39G+ebCvNvyPS6YFM2NrEyOcWvq4h/wpeJkAHhhUx3
i3ZD3j9VciAgjof73KmqiS//42S0/DDu4cjXajyTJpmZYuxwmr8ikSFdurtrBeUI
NoZ7w8J+trVVGB0RqMn+6Jtjdnlq1l6+w5WFaXIFwjbSO8wsHLassZ+NDMG6aJtR
Q5682EM7W2Vxb4GXEAdT4W+9CIROn0ienpeot9b2ySt62Qb0icekERcL1XOwpH34
K+RQeJ781sdU74k2bXjEswKLi2sMp6sPIhy0Lg2Y6swrioczi1/gNn+Y3LwMAt2i
jfbabmGQpJ6BSSoE7+oDmtc7szbpSXPSWmqkZQ2StO0yUijjAk9i/v9xT6nenk5b
EcJcw9P8TTVXRGOvcmTYasgJfFaXHpIP9tVb+sMoHulKFqMncDf9KDBV2noxIhkm
VyPh+j9mNSwV8IPJQDIeOUSnSDEF8BUp6UghWNU7zSr2HQPQ/m094FCBbt616k/d
5msKibVXhtB+HqmXTPRBBwr7VaudfgKDWrZfqn8P92ROg5JRxVrMHs0Y/yPTFWAY
KPcSTOiRr2HIa7Gpy/9yNQPSXNlZTT8A/FvtIkwsLgyGKMQywQLELYp57vBwEZ1A
z4xiXTUKjdfj+ufh15wPvswt4UfqUOq4hpUw7biuNzL2IlMpkpNV6+DQbbfMnonO
w/ml/atP4JGnXYebK03FZzcTyIWWS5Nk+OfNrCr/VLZXN05JrirZ1hZvjo/58coZ
ot7UTMLOQDkx1hLJoaRC/1gUCcDtGj9VaxvINbBgdERw4PEfnx8m6danpk27tWOO
2QcelqNTdUUmUmyiOPM6Xy7XlyWlQYcILE+zWqpBtIv2IACEEGkwiEf4jXIucEcR
jGKBXz72l8pNC/iq5sEJCwJGEsVMFl+pMDzSWPouB6+JbzH2GedoIwq+tClddOWC
55kEmubmAqrUNZ3QNgCkTkSDaZAySYAld+gpgwfhFRirhurm2F8iE5qADtcz7Bo8
eAyHds23Aap49X9a6lmgqJkuAtmtQHPIQwwrGg3mP/fmQMXAP13ETGfIfzzZyIfq
9sRbNEzijmEcKoO3txdMFX9pZ/619KTEZdmDtxpoA3mXsAo9x9unwq+DBnGSkLjp
a9K5sVKoUzpoUbjt/jRLCKuqzeKjPHzs1zqhyBygt/nK28/LrBMipFFp9US/yK7x
/84qtHr5ohDSL0heblsHuNqGV5R7mrn0aV+gRtQOrHF+BgtGEMsidZybNVlbhHfU
s/jSl6t68uphuHncBJvJy8f5sFQ9pqdFOwmhk3h5qRdp9jm1nEPGcJHFbx7yl+34
Dp3+CMadoTlWH0RRaiY0y/pQjMQLj4184jQM9i2kHrj5RxeS0L4Mi1bDPyDWJ9SG
sqnYCaQwZmh4CopPrjnOjlfYuGndkZHUp9N8ycYB1oojszuHbS44i0+Up54qVxK7
4KOdlBgbgEEcYA4P88wCqaI8zdkC1KqgVHnRj7cdZOLZao9XWStTFG7fwpjFz7WZ
DOMBcrUjwhzLhrWnxrIdT9g72vrnjg9WTSt7GlHPldqQdxelx8BnYbCdwPgEHtgc
GC2bdLeLbI3jNt37FlJJRTboXsvAO168bl9aXcHPhNPl1dOHeJK83RxVdyWIp9vf
KeyNRH+ew3BNVlOjvJh1xzJFQFJ/Zo1amOE9vs/yl43KfzgbwltZME/dekuh5f/t
vuhaCDm3+vIZOPbYGAfgdF3AKG0d2JKWBUTftNa9H7Q0sC1FornxI75MP5N7IAUt
e2VZr5FKqTAOkwpkgkVdGHldd6lpCRlr+GrAIZOp7ET6YKsoYG6FipIvc7mBMpxg
RSxFbwXXY1ta+1bPthXFnh/a7COjZ3cskkfyw2aIXClrRgvtncyET6QVGOPNsETD
2Sd92LTlkedIE6CE5z9LubV4hlfyM0swOW2+Vx6+Dc4Qv2VrR2C2nOOvD39hB53J
y/XOZ8/vjRsYRiRma+Nal25uWCUaDtmW0E5VNMDF0s7fKmkrzfyRaTA+GMQHB7tn
AhYtmXiLaJRRM53ZrSnoip7vsle4pi+/yltvZwm3gPYSSBuqWcFFn75hP4Ty7ISA
nXcJKDj8LF59kt3uF9dhMXaKmdS7vD2He7cs1ROeiXH6KJ9aP+7VMMhLOQhDp2wB
wU3Eiopq1eioBGX6L/Gi8euKdWNwjc6FxybaBISKlN/MH1WVFoZVi1vIAFTnBsYq
c6rjoAgbbkygKez+YjUteCjnD9KeW2XGukRvv7ZuYqMNN0fS9zbPkCdMHjbIhS0d
FNdjj982K4dBIyjbb3cYk0gt0EumXLzhI3So4ROOR6lcKqeUeVi/2BAg84iNbnlw
OkOxaHACTuRtv/lcwlv9S2hPoIwCwYYQW1/WQ5vH87ioL/acd6h42Iy7eOaW3lY/
gYfYhTSYFrJ4zIMP0WB2/pa1bvQs8UN9LXirx3z+LTavOktdOopBhOeiiC+Fmgok
2LyHWESNwzZMr2aPWslgtheej7dVTNCXCEUlD0/skaMuVjIUcFsIIvm7UU1nIpvi
7wjt2R0/zrEt/w4viTCPP9HKEtsnQoHRLksNOyQjLH9c7+QVSeK/Paiq8+41f0wb
n0wbTto0+4o4g9rUidr3HWK9WZZcZeJf36HdlPmOlHQigKU8zzkhtSPbnsFo1J7k
9iQ1tAEn9ywlThldXuitw40fy+oYtK9xVPe/tshgIu3hA5Gya4j9fUa99OV8Nfc9
d7WsoqKucWQaEH7fyxd88VCWGhTNLFISw0Nc/Gttpy5UsyWiyflJL61JQpcknczp
vRX7PkCHaWhlyEgilOdfzhI2yj2JjPczw+0qgKdNRJmvK50dZvL6YnJhwE1YcsPq
HjbOCmicWVSl+y3rIUHsR9v86582iEV8Mp7rDk7i1vx1KvNYYXfAPkvTeRic3TBr
KPg8/bOWRgIeF9OYCUctABLETCclHf8lNBjG2Rvh5A7aex1KTZ0vJBBkIGNMAkJg
jG/ELxVH/VDa0sgbyETVWjD79gP0gjFjeyxB3Co3QULadrtyolKbaRKsxqEvmuEr
ucSrgMBJzj18qqYgxurj7yrXyrWQyJ5dcPeMobssHv0kin/xy3FrsPFOAQEcOKdG
HmwItH2BpLkvK1BasOYe4zZ7pFeHhbWxLS/A8DDz6IsWzTxIBzWnoY+BBoy7A+k5
UKfSkw0AfLEE7XbBI8Eh1e1gDk3KnY4aJ3kLcMhuRh7UYxX2mS8se1H2XMIkAlbx
8nlQaKiZrCcIpnY0jgTdHc9Z4RoGj9opvm+R0iqrArtW6rd4ySfjglhLSKf/w3KJ
YU50AHZaUDHbE64lQ3i3qGsu2eWFJ9p8dMF8EbMjIZO9EBy24QNuZ5mQ4ylMb9FZ
KyaCOmxNkDT7GiHyLMTpgtOPpBc3dt4wOLtJybpKmp6B80HTK6Zlt/hxjMEmzuib
OzctRMpZ7diJ4EjRAUDdzTf+hIkwrPeljtq0Jt9nuoZUcvCbW4JziuUOf64Tuh/l
yxUCxLGCAxxF9/Dhfg4KZQvxzPp8naf+EpxUuv70v6Sm1ecCpNn55h+2sHnkECCP
67mt1ODI+i3NMQrDTShBK+jOHnqy4m5Y2/r0liNBzFbT8RGAizv2ZA2xipiLlfKv
cadq5CR074dVfbD8SM1s+hAh8iNHbDMww82qFhRBthh5CsBWmkNycpCBzYxCTQMg
ahvPqJuUXYHZzS8+4KryTHDDvEhouZx4IamrAZjslmwyoGNyKTcG62jgPJwpBpwx
h8AfYs0eWJ6pZs1sy4Gh0lAvE8SOPusl81joyWZ359SYj9AlfI9pmyIExYmLn6tc
Y04nsX10Fi+K/uaTIaaBnZSf5Sj3wKd8VTu8d6EKH5FLXrLOftKoXyZ6c7xqh4n7
oGXVf55OUiFA0fGkvmftKXZpzi94GsDJeqt9IjnXwGzPPngzlUmnvVWCpTnx43TY
r+ZnNFYTsw5anI7IXBrZB8tFU4/ghpBMopxWrk9xl5Amu4D9Q8L6gO9PaA1w+v0W
ISPXik5+fLY/LuF62T4xR7/aahejqVSOO+DnQI0bb5+tJNo3QwCxyhw4gbSkBbc4
Dg0N6GFsQdqbCLVifgUr/XUgUbjZ9WCCXmen+wUkWr+V44tH6TSB9kxGO8WFsHau
54ylSL0BnOFMfzPNdHWxDgMwbeR2/BtR3jXN6OYZ9jgTv5Q0MrGDBtv3nh+2Nsay
WDx8x3uFwlB9An8x0ZPhC7vk2TM/E4n2a6iD9CmTIcT2KNkOeNzmF+iVLTTDdLrX
zwvzONmD1+PdGCgBx2TBpVO/XZ6Kg/XrixiFqPdvb+MX0KgrB8SNnOQ9r5GED7r9
WlFByF1i2XpIGq1ych6xqWzkOOaBDksTZg0sY+MNzVz5ulb3wT3IREXt79Nck0sF
30XiSctEhZO1LAL+W5ZtnKlA5vQdWrLt+VZQdGiJLi4s6juSVAmNL/oiossc0HGV
ITUMkK7Bk9yw32Ms5t0HzpWHdInkNcEvQkibOcB0dfI76X4gNQkO0cGCW3UnBqGx
ibKVpXdyhrs4hz5TYg5ME8ooyP/TCqdtJksr/Xguh40NdzWh5JeEL65qgLtmAqkS
1ipaMwFzdcayY5NJ9SbMXHufwXTogaXM5sVRLRRwF2Q8d/tK0oRF3hOD/V7ndJ0T
IWPbvywDZOeA0r3+IXCQtYTxgnAMdQMCnPvP0enGKAkgXU07oYtEJymo2gLGBLTI
RsSIEKOIli2Ym7/koo2YZyaWqsl0QgerkuQ0MNGefvl+VPKjii69rJvtP41PfUPq
aDc+GH1LcDhIXU1w3AwK3j9rDE76yTBp6zLC25kbnXoDuk3h805HkW4BW9LGWi2J
G9EoSfrcQXA2a8bLTZ/kDr4yW3LR9VDva2s0AOpsdEUjAoERGW509NCX4qMtRPB8
ghQRTa0yly1PnS8ZQ230IVr81rvwRP/q3MBeEBXVHewB1urSXHynIjJ2/NgCHnL9
seW1k9c8lCuVx4LEKA7tWTKh07nwreOxedFvp2eUP6VPQdrn4vkv3NQLsWel9B9E
SfrKsuqmugUhA5h7X1MYiL0p6DiCZlsjEMmBEU6O3ctbtIsIAiuvQGv31L5CDABm
DhZCKawdKKaeHGKQOnmrLUYoP7NOORshOX1MveG7I+Y3YlKd8NuvuxajX/GOS8VH
iSCbxDyKQFlMiKc4Ww7A6KNoEWqRaELw3mw0TNhu4edUR1z/DPHXcuj2KUFESyA0
2fbWjMVQwxEDPOU7oakNYkIeZw2WEP2dJa8ccz/1RWF00KPcwl+CFDXYNHrFdrAH
m5YxtCp+6wgQoTKLhaKMNBHxUNdzTT9LrX29q1Ue1Zr2VtYWkQjeKn/aGhq2S77i
qhUJX6Gf87OVb/8kEAHcJw8LoaFFI3srEGgYEHNVtlH5e7Dn3zmiljU3GJwCFGEZ
Hemu5owiUZYCEorUF6BHPBpYqBViAvR5K344btqvtcm+2GQ6Noyrn9ioCTQoT6eV
Vfbrbfh0bOoPh57OPwUmjt7ZEfpCigJcayaMTJoXY7KO7B5N3ZAAjkQIeAoLdMeQ
GOWU2mN05M6Kwnl08pqnn3azqrvu1p5wBcBTpE4Crc5aUSMSDhUneV7PFjg8FMtn
UJVS4gEKQ+l4mBA+GJp0N5pwybwWGtkscWyQJ7nnp2tC0yHd0v+hYoPg0Mhqv9be
6aABYUBRIgVFRlC3dQzMsnJ4DIDk3ShEIOU5h+mdfwmC/qdtBvKQVxo2SAi4xuzy
4KksGQRpzIC0vO+eG0pxKEwqSdvgSdgEA08el4qcbIiSbe0VdqkckQ8E3mZXgkJe
UnM27N6ISx2Zuakl0T6nbb806Op2VNEMoZW+Wo1H2Sua/noP1RIkkKGGuSNQuatP
gHQfVg4j9SxNhPD6PFxDo1dYtkztonLSU1ws8VNmxFIQ7YYuZK1xwO4GzkQrXRG7
YmleuyKXyvfoufSc6fZsQas3fL0Zcx5F93PkuT5a3zn8okVyMlEocAs3tLQVWQL3
dRckZKUqzJzu2O0SOIbFMPBhzY7uSFtkyH3XhYTr46ZOVge7ktMtE+88SE3aVDhG
6dSvldYwtXM5QFxqIDOovqN/oetBMzB7beBxG4ULE03+z86TUH4+Zbd7/N4CQ41r
YbZUOr44e7DyNhIFP0Z1BVuHBkqp+iTsQ+lao6eFxgyu/YQYg6rq5Bsge5JJ/isO
7jKPmcX6PhR5MegeMUyUOVHNeWlt87o80BuF5ueKBmPIOtpY5jeWG70GPgs/rqi8
XXrEPq2/bi6hEnSC96MWGnT8f3A2XROQjWaixYNxSOs/vR7VEPR1a6XEbhoPq828
JTsbrRKuR3eKB4eAWBbkLg0gtCn4ClAeyHkTLbZjCr8Xomz2wgC3luk1yYFtwncZ
tZZ1D9YYqL/7xba/wq6CBxaKcLZFY6WZSdgSgmjyWYfhnerH8tWwzomZA8YnqjWa
k+lR0EU7CQEXbD6/46kzQl8Z9QFYml42nmzmElgQjq6sUYo/FPmACZ2T6oBKCDm8
XpINB8P8u1zp7hCF6Eo59QjTqqljLTjBR2CKrjsAZmt4+deHArx8bNLO+ipTevgI
xQIMNhKgpfQdsbmFDJbiGwo4SGwkeFRZNfuXgTyPSflIgUjtt480G9ZQCyk69gqt
xQgwkY6blKdZBHBusM8RP2AGoar87ZfmRoeem1D1vgZ9LV34c1zkUF3dsE7+wv7N
1iXGCd4diRLPE+3yrWchzcH+7yvGN0vKN3H1R/ynXSJTfwWSpKqu8ChoXCNY1Ssl
EbJUICHHLVbtcw1T3OoCBVmWr/rLVESc6g1jPU1x/P1EVeKn7OE2YFU7LtkmZmFR
DpraxbXxighhJsjvvxxv6vVXuyb0WMAZsBhDNJpKgbHK8vTtgKRcHr7czHfVM+NV
462a2DN5LHtaJvJ/q7fiUjMhQM1ujguhqmLmN6++PaI1+oMESqgE3veRzVax/62J
ZMFwAUfo958vfEvcZ6uK8VYLqVscoHG8sT1oLuhOw0fxxkqLiwWc14Sk/bJ95AEj
pAsn32B6zAOJTT71wmyc1BV6CqbyfjThBF4Ots1ukqAtYGSimFOOQDcpz7H3uUNi
XmW8cR54E/NXA+ZNga4Un+SpS6j10iEgesJ1IcytMGMWgttm0+M7jez+4QzAdU1Z
mMxD3ep5tWpACU1C+kNlXEtarAD7FqOfCQ9w39EyWVJjqBo97RSRh969OyCqH/uU
tczMzNeBnN5KPakZQSII4Zk1qVFGrUr6qpX9y+oQfdmCkZklQynXwIvzjTRrdAvA
laaU6IVXKD9mHI62hyPR24eT81ALZdE1aTvBb/dV2/JGv/seOHFcpwostb6uTpN6
eCKIZ7cFMgU2X9hP+ZwsB965skoNl82qUICTdHJgYsw1r40fsSysHAThl8lRHvd7
8/N31iaR7IubZR8XtJlihcsvgEMXELuOW4jIEX1bie3tjGkacOJ0X1na7aFK9X0s
LZrmf3HmNc/UarnmKerPY/dT8oBWwyT6dXMk1dH0sf9nixgtA2L+zP/S3Ebl/rAh
Cc9YF73qimhxP6K8BxTcNVChHE8MF65RKE3GkSWux8wIfzi3hJOQl4LKUW29Kj0b
4V9pDBob5x+ZRw1mLEgrg+DaSFo8avDtWdizEKLpwcBRT/JSEUaQyfXn7a2UbsLy
TFlnVWFN9J35PRtsWNUcR1KjJi98yb5yLqLRPrRi+XrzBoNfcmkTTZSUMJVCy/sx
ugJD82X3dxpLHadxcxVUeVHjSjDdIA9x5OG8odEftlXd8TG4y4cr1z0YrcDR0W2d
dlUbef2vOoDnhy0MnB7hjy8F1hKkyP5++2HctTzseQPcG/Z5pehTjlbBGFqwXsGx
mGYBLMN2zKDQ8UmsB4706vhZFZJS58KzZy62hxEW407sk3F7w6Nu29tHjEXcuQwg
FLIwLfV08sD1bnz7sywHY7Iq2ppWIVzdHitX/Gsw7Q8Pyg5XpehYpKkCkNG2F67Y
GJDtm9Wb3fedcmYTNMCinVdR58Jf+h4a6WgbzsfF2ps7du8xlUvL28RyQ8f9tj7A
a1sWF29kFOyylv1uQnk8zNJOyU3gs7ejl7Y956OhpSUVaLDVh3nWPQpSFSmqG8eK
+fPJBoYSuT28DPb6lZemhwow82sTFCAT9Pf5OEueR0kEp3hMKSmMNdyzBpCJbN0V
4bRlmV9Kj8/R/hc4+3r8lHT7rzhbOPlGJ1/7Ste63xvaMIBT5+TR4Kap0fkH1ZA8
LehWPOR7cgtwmDMRgb1Vv9zNyBnMzkyYJ8W68t/eeUgcce5QTC2TH2Hf1jppcLI0
Xzw6omYWsww6y63ic13Urb6LdFERn7xE2yn/QYGH8Mit/9mqqhh3wojXRZGFRwEO
NxM3JHi1gcaARs8mO9wtnnTtZNKX4am3iGXdyFZuvV6jFHEMCaUCxtkoiLB2K6hX
ewOQf4OAT3TsJEsR7HNX2Ax6O8nYW0ucdBf+zB0Z4CJchOauuyeOAqghdUSLHsAN
ZuWJyks5Y1FvSAK7bVHMXa51ng75bY+EgDnYfO12LAWumJez16lZoZrw0mP2CzNC
Y9r6wA5HQCu1tGhEG+prOZxz+WM6zP9ehj8VfxY6OBASFD/CyFMAIzEiXTT2IGYz
dzizk3m0OleJq4AIaov1hz2cdeJ0mqtYTn8VHi1hId3eXELCULN0aoGRcjQdt9AW
RulUdL3pn+YFtvzV9ASNEe4Dk7I3q28e0RBjB8L1leBU0jnvbmnDRVxd1MU9beZ3
zQb9jeiHWQQh+6uK5cVMMmVwuyyZL1hQHljdOBNSKCpBqWH4D3oHU6I0DCTtpIbI
6DgTpj4OPqEMOy75jfoX0s0YGZxWczuLljRna8N5grTw26XCkIweCOu0qd/BFc48
yswL7EyrzkwJR8PI5Omwi+CYhbQ0rJEZPJEquSkTxlO0dc2NeD1882gaTJgp10Pf
gOH96UbO0+PPCdfBmlGwmxOnVwXFoY98loh1etdhSKCfwU1vn+MyWB+jr3gkyETe
g+cQ4/H3ELhNwGWnaLyZDC9kdUf55giDcIPDj8Rm7uBJ8i1TKwxboAewXuWQ9lM/
a7H4l9U59oRtNTkkBkgUwk8gOOSNNpViRPI6fKzh6lTuO/vzPYf2SYQPi3l8k5Es
qH8N2KBtDdbfwr8/C1JZVWWqTZulMere+9NGkpdn+F2Aavhmv1HeNjXjqCbgWBUb
rO04Rotm21GhLim78fGGT93D14o7STCrAQ5hlPt42DhnEoU55Wpbsv1b0r3j1p5R
yBjNi+GCFRhJ/Hcm3eKTLsmi3Y9TlKE3WHbsgOE09nNCjWvqlafv8yQdrMV4Ylie
22/m+45kmlz3oELgYzey80qNd1BIAFSjkoddlHUvVW6RvyomGkSRsiZ4RW1enlOA
06lDy6s3kodqh3ef5702lv2kONdm+7arlK9PVGN8KSCWQeCirGTLHdkErn25V9PA
0U8aaNtUmvaqKDi4Z94wLIBXMKk4hpbwIXHT1CYpakUstZxMZ/GDWQgNw5Y9DVh+
LxvZHpLULOT2oP8guJ8NyAGAruRdtir+d8Wr/biRJ0VMIzMjjeHf9vytlxN8AUkh
MWLp9kWusNf/OHYTR0CoZz4TShj2hBfEB+mMYHV5WSS7NVnL2naq3hmIGsSOD40i
Hyf1rWZn86eyObvMiTCZadgkTcNSMdI0guwilk3h7xDCMTQbVdpO4+Q9bLLCBtW3
PehdjqiUn6g0MqKbN05ThbCVls11Ex3dQ4xMRrVW1l1/zy2oQwuT77ezgUYBC7wr
GMxl6I23mqlox4ysgRFjd+rMtJV1vBSOmK8wHDkNdIk469H6E3RLHa1AmMcRJ+lr
HB+VcytOZvmlgf89ImwYmiU2IDbXDzRyMyI7YZ08unD5XB5WhYQHePStPvx0fwdB
vyzanGzlM76mgcKAeUGFM0C5HKMGsza8gobRGo40IkdL1XiUE0aHWAD4oiFKgXwN
bd/vMsLh/Gsexa9VIK+kcLonaWmcyoruIqZjMFtmetdO/zTZOnGfanaYpamW2KvA
+mQ6UMVZE4eueQZ+AIqj3NE945zflPNpn10tNl3DHm79n2XvH4I8XR4dEUN8/qt4
DxuXR/5A77gDSJ+mA+62OqX/JQBrZh7CR2rzt3JOJu8+zDYxOqznMaM8RBwb9NPr
p0fFivMr1GVzVHkKWYN2K32a9AWd1HsfiL2HoqIrm4m0+5VrN4F6XgnwQEIBvgw1
s5TBhVAC0VU2hETG4kcp9Q8/ldbl3m46iVnZE24uPuhuUJfKIH1zuXUrOb28oPp7
v+Uoq1ltXnlk5/fG7Hn7nViwQkTQl40ewdSonOt9M6oErDiyvUx+xoAI1rwmJ3P3
5z1LSVBXp2TLKiVjT8PLx6vka6M02LNWT4us/yAeNeJ0IGaKAm1XpmY//KfEEBE+
Of9VEx7C62NLianWpbKpm0Iq23GWoCIkPY8PQehLKfbj/woq79uXdpJsuVOFxlWL
UYOZy+5tUFBeg7tg5t1ES4MBRQJfQ0bFGzS1SWywTIMg9L7NEDXzl3oPhygZzxs8
O/rykl5uuxNzQWa5yQpRM/kmqXrSZaHVN6nlscUohnz6vL3qw+4fsQwkO4qcX6+J
fYNAk46HEVBzW8X82UPyh1CqPirFiNzGGtfTg3/8+UR0ZiVrNQiOMHZWkbpB/FZ2
ECzUQfQkuaWiV+mXmZh9+Xrb2Rm4nOcK6ng9PiYZlcPdNKfAmfOhC04lUmjDAQCo
3zzx9zSdZ0S5Ic7u7Xo1LOQJn4tDY5Wik1bJy9iKRLh94GN3fm/mpOizbMegxhn0
ZLrVOtbaTeLHYoeH4VoH1JmvvIYFK/KbVPWQkYeAYVktSVmEY1t01nPVkGJsk/wG
Bw4PPFCqz3++wY+filC8woKwJKCofq8sGXe7wgH/V9iypNU0/2VnPmgqCgQRidZ0
zBgazbNRmCPalB6LcIsIDvDrAbrkxewwhqcIRFN81K0jjGeUdGyM//dYvplVns4b
0zMFRjvRD7i3BUXFFXL340HCrBtwIDjZx5rQ1Cumxo/ZF+TTD30xrZJX7G8M9TlD
Nau/ZyB6jQkgHWXoko0b3F1xfd4HPxMn1LiqxGGjS2Hq8LZLiE0ipr/FMyefzcrt
FskSEFa2a6jrq1oXrBgOBHITdaC5eCSrrcH/j3Qb88JOjrBR+n/a6tzvNSKHMzNH
oKEh1dyybohKJD0xnd4//iq+n6O8LLlQb2uEDpcsSArerJT9Oj1kYqJgeoI6OodX
mPWQRglOPFtZPUwzjM7mByb2TETGBI+MmRZtlkroSQVULf0d+tqmG3M5VID/Uh0w
zkuLama9y/b08TYpfcJU4vUlPG493DFpD1vb86vWmBvH74kUvYd7+H+Ir5U/klJj
VO1cKtcmAKjVcVHrdqhuAxhrxr4Dzco5ml0TFa/U5Eh4iDEraHFZxisTx+2C6EUk
45+/D6O7Ev1Z3DGtykznYllKXF19kbtlLsD/fG5syxvWCw2ZTI2sS0OSJnC0c4ci
uZ/AzS2Tl6wnZt6ofzR0Lvr9l5klmDRd1qLND6KjoYyOt/D9jE4WYjr5QlrfdCIE
KM0v7jYj6C7ymoivAtJXbD/rpV2janRjQNq8LPuz1o48bAMnL5Ma2TYKxfqFJy6l
bjmXnGOz7+p/v5Sgz/oBD2nPhCyqzQh79drHitLOfN6Nrnxj9zffKQCAcxaeeSzr
p65ybbMjFLiaD6bFiaT+J+Hhb6yNJ3vAfUkG0gnyca+6oyoLIc61d2PCQ8DPeJfA
rOlVnejPtB5qm2HNXMlbZggxGuZLOhcCCxH9c0JnUg1NXYhBVcZXrRQAybvnB3wR
tl7GiwOsC1lu0zxWMvUogzpNyXmjPTIqwxHoYF60MonoX/PgeaFiZFx83XGrXv0f
tBwx7ge6jMOlweCWP4lIaseK52QK/Sw3qxmA3wy3f63BPWzZMJFrNlcSrldLl/w8
TXOeQrZ/gQIptMCstPqCbp9hseLOS0CY7bxNeLUY9xRBGoVWWAfZ4EazLhzFiL+V
QGGGNyt1u3cmkfbV8m+N8OrIl8ssKRlyQrQndN87poirio0ptQtVaD7YefJKBDOl
6112iHB2Wz/8RpLpCVAoFXDmpi1VcllZzObDQBsjxDMBZv7y0OxJfdz/4R1GeWMG
W4ixqlKeFhUexgLuA8+nNdGOO4CtIx8RHz8Endhh3yeAsKpSbdvLpmfveoKo15BH
hrvQTR4YIfbIgAAmhxE1E5wpHsKir4JJeqRboaPUZBc5G1uIqqPTZ8BmrNSlu8FC
+7bm4WaNCKzL0iyQwyqD3Pj4refJ3JLjE8dw42mJLkctGzoZKBO1bNrQE/RJEDFI
Pm1mvDhEkcrPQ5UighYv1F5nnfCHYCzu+ZC8VnEP8fxPL5VL9Uh7c5riYuLnVwM5
Dou0NmGN02VOd8dC09g9RuXVl+Qy9Y80eW8sA5+eLPzsPol2KLz+4L8pMVMS4t6A
zNaDooOUMvu7ykHprmxPSBN2oLkVQ71DPsi+TNvOiAfBNzReJHFKOh8QOog1HYpD
EqZkyMaj9+qgzB1PnfeWsO9YudnVoIXCi0NECARNJ0w8WtzNmB5RNV2B3IvQt58T
3krn1UVdYxIYIEulUK7zapnBxO5v3f6wvBfyGEjpzIO5JtBXOnnbme3K6bjXyXpJ
ASehJfNTeTEa+huL5hT1+Y3aVLPRjoNqljTbbJB94EsuxAKmy8SNmrgUmX+lLW20
Etc6Qxn1RG9xxGdgMihWr2SsibeQIxQGx9o4kCbeAZa+kY6VuCQzxJO2i/nAK7oB
XWk2LCRZJ5ryj6/dYo/n9qPjJtioJ/FjLnr6H1oaxP5ME2ZH94VxoLy6eChKWSfo
9fte9EAH0YDL1iJo2E1tGsPfmOnzi85oMdFbIKUegf8Ae0YZjb/yiuDkWYzlMrAL
ijfDM28Jl1LIKfhrQsmNvFFH1PItTHEtcNLiiHV60H0KnxcC5TYsmVQ1Fpts9qRP
cgF0kzgLp/1T0pUepzyFByxcx24BHT87vCg8fx4L3A1eUpHtayScsvuf+l8Vgrwr
6KAbtWWKffuR3X3Cf5noD3Yp5g1NlCup7xyVHIXhwIAAa6XprYIsTnZzTt912k73
/l+FrIRPh9L1rPQwABqShshCqLy4L99Bk0eGuzgBQZ7NHcjKXQNd/cKUtmfIyo4f
Y/iKt5NcEfEC8BlSNOCVrGIDclnTnRplnSmNSQLTouRwzv+vXc2sC5KMhic3g9Q2
lfQF4G+6VRbFCyHOW2v6/BehYxOu1UZ1XmSgdHteNWjVoXBUbeYHKeTFtxJIDN9C
YaQ38yPQt14g8i21aaH/UmzsJRYsM0guX3x8xP1jMpjUq4HpVx5Fkrpip/xsYofy
LebnAjX34c7cSFEI+/I89zhBw1F1RtBARtUMv9zifoQrBtl5zvdB2tvpKWeyd0fp
hPzthqCe/lA1ZhN1OY71J+ejNhJoivktBoZBPVY6rVOXFq1HExhlmJeBBLEEGu2u
OJfWha60o0EqXagNO/jNyeLsuFLeVwRSRUTU06XLhb9kNgbNcvcFaq+GRaWfeScQ
JEMEAgpYqZMMHb0OZyKqlrPFPs1h4kJRflJurEp7pX+5mMdeJYazjchDTmKVuQY+
Pp8gSCYJE0bo/ogrgWlYuesL4b0QCVwkilY/7sEY98cxP7Vr3iLjxdnK3P3Y60xb
5F47lMV12thpM32pqBk7yvNQ+ZJ6+mvnogEwPWp/7z7/eHsxa8ALIL/LLrqNAjmW
OQh4NifvK46CqmcPHxkOWa4+iZtJTo106A9/esfWonAbBlMa2BXmsovoLFnwAbCb
nWcYxwF4LUIt9k0WMJVSMYqkz1AIpxP6v6w+yNWwQGj5WUHVIiCkZqIup8Js3x6j
ZHiYB8KoZ8VR+ELGABDGyjq58FqwCiKABHO7OMkmMedSIFoEpZW3TqFU0mAJ4+Bd
nd3VqHTWd59EJibq2l//z9l577WvdldKEGQ06If72migNSYzmby/tYCPjxyHsmye
owcZmOLWwhEtKS2bOST0dr5L2ZtvU2x/c2C+MEblIXo7rXiLXzDV+f+mC2lSdSk+
t/S4GTFa4uoSTI+5NG0th51Yj69x0a1cTaGoojZHc5dLqXRFQWMyf6uI8Ly0ioej
+DLYR7kOpdGtl3JSo3QvlD/viy0QipQOBzkhvbyqtaA30pH9wbVuM05hV48luT4U
SC9vrCKJIcwhxy1Y4+GeknzbdlT1nT54oellmzI3WZAuK+qY5NTcIi71uWNFDtAn
K7BKXUI79DNlyn7soqCXr3eMVlDKfkX9z6L4PFbGotp1V4z172T43YvNCZOp5Hqu
mwCDuRM6voTMAMU0UDxg7QVYNmWkGQDVxxA8doI0CaJ6OuHK5Y7+dINf0UOrnRQf
ZXRoMKYfUxyZzRY/lW2+iRnAA2TOCvjdtg0qwJ57lCrqM5pTKN0kzw5cgw0Pmb/a
zqCGRRVwXgwregrdP9I4x6uFWerKz4U6JahqjiBHWdbF7FAHtm3jFybylZIfmqeF
TR5MDQQCJMSvbMRka5cc8/Aro3CxGftZnWxSwp1WG1mX31RYJ8zUKxgLHoz20pHM
Jn+JChY7HCdpP3o2CmW7X0fVDAQ0ckaO0TJoRo9Ti8+BM2qj36/HsLid7LkRVslP
u3gAcnB4kQUWSahoo71Gc5DqkAv0pYRN/megj5CTeIPjgXQ/tQNm1YOAoE22YRuR
7Qa25t6aNI+jifwNo8BJHXddfUX5/X238Hian13q8gGbnDxZ69km2b3p9/ifNEDa
6e3aMz75RuFQh/WOW9Xx4Bjs7BrxiIIUDVlAim819I6VU7gQzI3QP+2JE80QxJkP
90ubXs0kMcZ5VnZjzByuVnJ/CmE1fA47IPeocPKMOOAVVE2840jXYIsX1n5kHPkv
O6FA3rh4rvFZea+zPKkqQedzf8ATof7KLyxqJNbicClzUCLz5iSPAuJYo/LKrAt7
E0b8ww+NpauTpsv2NjBxJVqD3x9jPmLq2k6nv3CpBgI3v3hiLTqEEcDQDTW9iesE
Soeb3OzoYkWR3p2lgQt5gOPSbqwzkVOkZhIyjNXz7MJTRvnUV8bGWdKb8GYRoLPd
QlRHksOHTt+YgY5Rw3EIpr3zYlG6dIwFtGK/Bzr19us7VQS7pAb7LlXwTLlZLqmY
AL9dCNg8KXvFhgyboSZtLVHuBm46qYTOQ9ILbur1ZCw3hvviM0UakFHmgL8tSKaq
A2MrQlrEkw8r0YKAKfkrFE7xuWtcoJEZxpm06Hi9C65VPh1EcFTmEr4sueEbtyjc
CeoHkFb884whDWBZ1akdnjezjYzu8qQ5aVVPFH8kj4zvFhDn74DiD0HLiee4sWN9
lqiw8yVlaofw1jIKH4NMI/xQsTOsaU6sl4gkKxUlhimCekKkrO2nPslg+Argg4Cx
XJMF6mOQt+bm8VFHulCoPsNPJYpl7D7abvTGsew76Ra3gidrw2fZc3s8hzcLZfJA
gU2kVlDFL5jIiAF8ef4pcxEyIlvithXszCtEGaQk/xONCEAIS+txjge3k2tlCK0p
7AyDONxeL1GF8ZBOcP1OOXZWDp/NjPmcuOquPzTLUJ2NTTcZ+GFOpOgZ+US85hp7
t0ykHSdZw+R0p32X5pp3/fl1/M+XR+UlnhpOnqNn0Z7zNZGmUCeuW7eDr9LZlOAc
faTIMPAm0mmN7ZjBNIW9QD0Q5ISY/VBqw8HtqvTERWYN77GQKYB2nziWM4rUWT9T
kZ2JOywIHpUVdfvNy3oQPnXPbT34FJr5Guch/p74qr47ld4QCI9qf6KjqI2CKBWM
N20vtA3FtU64ZschxJrj+vndy3e9S9w1uYoMLQKSP2+/2E3/Zo+Xi/8MOgpzkfLC
PBp2naEgC7LriIzVimFpL9Ret8Asmh6LGaMN1kHx1noQRfEpO4QvDbRhdzPHhcM+
K3s/7oQDLAwX9duczipRrxlmsbgaFWKkcmkh4Ukd1pgZwSsZ4zKH/ELbrRDMD9Dk
TCwECQSr5Uj+Ccrguw3z5waY/JzgGWpq7CKH7RsN6Ya6X07Q/B/fUdjKpDa+J9Gg
4Xv4KDl3k87701yuRd1uKY5j7raJVn1vZ7bGDgZ47xIG7EyfMD3Uxf7qRQRZ8Drs
/XeZEawL0ROF6S5BxsiXVcwa3GlsLbWCerEuWEHPVl78zGfYr57RoJHzu8uRAy7g
49wmOYgTHLgV0U58+hoF0Ot9CBi5ga/yOLpLv28st4bgPEs/JvET+ND3kWp3VDEZ
PGSfsrRAw7bI/+h0kRjOLmN/vHLvjSr0xM4601y55/tmNDwOotuOBGytVKYskskB
OUC1PehmmNrD+DZDLunMERCk2DDcdTIlFjuTar1QkNmRZf9LoqjVfq+X8h9anct6
fGplk92BWRfy0UgTh6fk1PC79lezktI7hl+1TJoo1zBASSi5bRMptNMmvY2jATzj
KuVtCIEio3ZHhLNwj+3ofz+FEuiRwZhHBPeFoJyqfZZup1nY+X9hputLX+o9Mpv0
I7aHCyH73OiAibatHBb8As43/bgvNNBpBHXYMfJP/EGSPXOZarPDVS0X3tpDx0fQ
52+TdzoYFV0PtAV6nfX/f87pa5/Jv8rz8jjO5kQvfpo5FnesoQ+Qc+HqNXO7nFfi
dJ62N3/k6nvhHHx9z9JGYL7cwl7b6nR0K3+VRXLBfKM=
`protect END_PROTECTED
