`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qTGQC0+FnJDsssNkBlz1WrjfWxEfWSJVf8Mqh2+iCjpbn5pnHgWbwpi+/Ow8fgYR
5IXwC+zvGvhfjW9accGjRg5wLDnnD8UPiH5/JPayq8Cjpp6FejO3S6PMXrHtHJBS
lAslo30YChhuYSj7YTWXAIl4ebHTgR2pfsKNU99LN4sIpt992pCxmwaw2LIn7jHH
FAib4fypoDGpeM+f/AjcKE5t8H5aZxJRUqtMVhOLE3rT6XyVwLp5xKPne3xPYIn6
txZwFN064VuoTsnU52h88E8V2b5o1BTwPV5nCBuv5QFnJlEQlBhixuOQZ0M5DaQu
9Wcaf53jy0UmbIP3X3HBxK0Tv04906Mm61WDhQkbs5xiPI4UEd6+IKNah0SREmtl
1a9QrKKqsFV0L4UhTMnydPM2B8UZ6xIeW9NqGrJUPXAFZeCUdvIklbouTCMgJbTO
RNHgkaeB2rNNGmjo1s1zK2f2VG7SV9MjqxpL94weBAcOxFHgVVGCLYwYkKeUUHIn
WOf0UUhi4oZoo8N+UYlM3D9iZHuFetrzl8i1jROQsACmp/5C2lHjVcDvMLSI0gIj
BQNy4UVs4EOT9HTySWIb6Q==
`protect END_PROTECTED
