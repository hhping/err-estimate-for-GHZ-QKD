`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q+6iZvm9lnVT404DmVdmqQ/hkV2nQQ5vSPosT54ka5afPw7+E0voBBX2Wt1eYBLD
VIrQxv5/9dmsMEKe4pAVS/6LX2CvuhN0uTbFDIFEYQ+h7CA2YqhSSgTUUcUO8VXC
0mD9wPk7dVt1a7HneliePr7D5sB6vWzjYUZvChq7hUwxzpmIxRsFJgLlKIPcjkyR
7s5LQVNhfCKKs3u5xr4AP14RPcxZTu+GUg4m9v/gTtOUTZRWvqZsEapNFDYBTygI
gFctr8BW0R0ZDN3Eds0cB8dutr+HccZpSzNYopHVZsJ25KM/XZ3xwzKeGMSa3Ti6
qKfLqEXOf6nUJH7aGDRDLuiYjQobeJiIfZK0fq/a19o4dYH0fbzEVEIhw9FXptvD
lRXHJr7ynSFWdXr7wQ4OQluL37imcF6SY5AszQ1Nk+M2eFNjsMu7/C5+QFprO2Kb
uKiCEeutDesprzTxsraVTBY/vOgJDG6M01F1GRDytdqIcyMqjFoxeckqbs4GGcG7
91+gGKAhodjGNJ+k86nD5Lp73HIRupwa1eaZz4vLjUK0aIcNYRSvxYphw+mE8qb0
VBALwL1hRFqyqa122b/JZU/n4VHvT0QXAv5cqhTAybUPiSQYC+36i3KjW12E99OY
ojgy+Mrc69ph+AiG2oGatWN4nyy+jwdtpUF/hcSCL/0xGD6BYOSzDeDnSpSS1S32
zm+qaTQ9L1AQ+HNhPW49Wf32+Jt0uFjD8BKT2GJxO7rryA1KM7FqqZcB63FDYL1K
c4IbEb+jfb49cCWHB7qXgTJnChyXiyHbch0MgdfuiejdjCiz3HC1PLlOz8KltojU
fzq+F0wUud9/TX4ji/5ZniyP38KvEHCmpJmW4cwlKJ48m88E9IkQVlwK91bao9um
9wWwGLjJ9Z7jT8DhyB2WvXTkn50OU9nLfT10jyPipojt8BX0gk18xm3ZebJVuPEf
LD66Y1g+u5oySpCNpJxQNbGZzi+A39RZiU6P0yJyqEa3XvqNnue9awfdZojkMe6E
3PuKskKMSnLeXOx2MaDyWVvSK9E7zB4DauVAdnhV9zL0/GBtKoT5YvmIo2uEAE0i
7gsK05zorL8/YKjzG3BlmJJaEI9Qob0cx7p9ZpjPebwmw4ACjMaMRZY4onGD6nyS
NwP8e14l+n1lq6Ukm2oxQYMlHE7cCu8wEMgc4qx2/E0M6E14R4oOei43ZD3SPwaR
d3AVr4uHak7EzQ5mFtqfWi0MFVZAr7luLgvZrrpHq1Xh+QbZ9S0uyGZWXnDlQJt5
eQfOQTikvNLhAgOthjq6E3jov4FcRWhUj8h4SkArCrd2apCfGeW1PduBZtJZnw27
XYME5jRxFSuBUVXD9rXe3k5gr0j/MWH/iHf9ByDevR/XpL6Lwh7Kp3JC7wwEwGJy
fjBgWJYx5J73W5536LC8lGKZTwdUP46WODp1uxI9lEDwIECRigI70JOyRK6sfZ91
2NwcTh7GMV8ydcbvmdvDpEh/Ye4Jp/NDK9WedfVSf5Gn1GOl9+q42ddVxRB4Kvrf
VkbKLSmPjQjn9br0ZewM76HY4deLIQA7CUz6AEl0zvcVLMhBVJk7fjaHbqZYL0oB
0/0Szi6VYrMBkS39RWCRPLbdy+0fNG9Kf3fkbIgK3da/2G4CEV8eEGcJ+PWP7U7o
dg73VrVj+yac9cul2WIHVmAiFJAAC5iCLzy3mVOQ3xj9K3W97lPMbr9F+lDWisy0
06RDNHyvnF56WLPhbtASNiF5mY//W6PQ84j7GIY3K0BpOFEMqgNSMQwyJ9RlrS+8
s+61Nc7Zd/3bCTHEjoCNUMDnvO9/wo5jTtD9Yij17YN5DsUcC8Op3lYP1TkBW9bE
pqNckz0SWKzRblQwyrxbnTwko5uGvRy7eMdTmaftmmVC0uqqg4UM+jMpkEv1BbR0
MYqPzbAEGDCHEvCdIsx3Wo6pbbkjtqmaYXMYlgTD9aoSl2KP4fgSDmYl+60MWWM+
xUvvd5XaE7hG7y2HOvcy/sLPIF+MiOcbNV1F+AaNEVBnLsoX9PKkWxqkDoOXwhhm
S/MMBbA3QHa2CJZMUlcBz3Uf8mfXxBOPCfVHdw7Z9eIBXReu8/e+7xFYjVi8beOH
unNpU3HYutGSO0VTJdFZGAimaqmuELT11WrrT1yCIhlclt3Egja0hZIzJvo9us4H
SmoKNsL8CJgBcKG5x09JKm0opD/bcUhTr03DMpkfpbQuvZrB3eHE/zqJ1eKjsV//
SXd3x8Rmf25KUZ5oIDrxtP/qzPxQJIe+PFVCb3etr0TOh3J+xdFFDahpMvTpXygZ
fn7eO+/o/8MAUqlYppAUXzB7lM1JNZulCmLezWnoDXESdcL8+72YvqznoLDJdIRq
KTuYLhH25jcjm/QTtIxbR740ZXIOyBd1I0EJ1eOLaXdiualR1pNkgMWDmvbM5du4
vE5s+3n0AkrFuof1WBYqJmUU/qGp2NYap8iwjKd7PHqUkhyyYJLbNEVarLNAoduT
bR3lgMWM8vWNijYHw1GVXO78HfzaguO1nDxysWs6zUJGtbDjyCUmOkHFr2xaltbF
l4JnndllZRDkXRGJ8Q+SvyIDEfQe3mMcimYpYJSi+2R7gdobOZuY/Uv2R3JzyTSC
DovzpywcbA6pitQy8EFZR1tGGvqugpuM4sy5MRqUL3uK3acxRQsdYPc9gcCUqtK6
ZpfiICjJyeC+6lH6q4dM+5uY4BBtICJu86RCC4SUpiSQtJQfzdKuWLqev7u861Fz
TnEhoWnoevxINHvWGacDCdB6v8V0Rt9xK1RyC0KNn3wB8wK61LK6tg9OwvwhIyJt
osMr+tal1qC+iu4CSBD3Dz+rJQd9eu3q/yP7J/5t6SWsylQ3PVS1yt8TwJSLFo3+
NvEfu4slh+3MsR0qpf2l1s7b3HDacT5t42jNUambIEtZMkhjYs4UdFg4qgJ6+YKe
ozb9lDfMHkIeIhwqvZxM7gYmHdKZQ6DYWeTWu9bRBQ0UdimBq0YcaQj3+Bug4+0v
SwZDReg1GGwAKQnkj0QFY6lSyTsBBfj+3KImB57y7oFMnhdbEnu5oI9whtSb7iqS
rJFP8jjP+NTJRdqUdH8/MvGNhGUqCe3EwXKwOwQ2AoEpG0bagjXzYeIvblXekU4B
m3WIt/B0fsL3hp6NwfwGVBjHt5GzjEVvN6jJFo1wOOSAB7+u4eLRHfim2Cxus5vl
U70z6RxNSxX2koHu/uXQVwTXax6mWGXS7ISAPQsOOLAUDUgGpLuGfthZ5mb1PdQm
QO0uMQorHkoyu8AGPTMyE+bL/W6xR8vTodh0DD5RKrCvVuH+TOWg1DVG6W+cU1Ie
5LZVa97nMLNf5KfsZxZMa6DfCXhkQyUjJE3tKWzM93mDLhPsmw/0diuxcrV9R0oR
8XXDZNQnri0+wicZyFkzCzmDQsr7GkNhxTuIPuAhUtAMIQPfuJugaHwD2BOkf9+8
cDm1OFsfz0RVt9E/dZua6COfhgSu+AJ5Ecwy34bNv0rIbc0VF/pLKXu4JsEKkeis
+OH72tcBzdsgjRZvgQCTyOqduWDpMFzHthS4q3psbAceJ1E0eyaaPUPc+nSZsvvR
Q7OdpRK1aEEvWsmZkVoPQ33tP+eazqQ7QWZ3Is8tQv2bCEa8umxwcYF/lxtpDUrx
BzxDjOyPneRWgSI3C71rO03iS0hq7/hc4mKcEvcrqYzMNYn0QQzrE7v3oR+eVhbZ
wUozl0tOaaQfbYMnfv98E3wdByEDyLqxzMXJYnBRlpaaZ/0mkrdrIYwYCJdXw19X
Qsf/KIvHEyVBlf8ASldL1hY4uZFhVd3VDSRmc5eG3PrlwHwkVk4Puh+roVjvo1u6
2ayqKdHYguITEJ2YOZ9OPuurdJH06JTT/vqesf5hjyJU3AnNhDMGjio7tDr26zOR
2kKSr/5q8JyqTR5hVbNqYVoQBgtqtywcxxjmMI5gpQA+CG+b6RvpVL3O/xzf2hDa
XCCVw5pxQqzbUOjMIOO5O67IQhrr/908kzIPG97y1hfWe2h2GUz9m8mXG1h9GeHn
pu+vwuah80BZ+sM+VC0XyraIb0ah9sCl3OvV5gMuLqogynExQIBdFPGrvNNMvWXf
0VEgM1bPQo4S2cQZHE+5AKWscJEEBQrfkjtoQMkJk7Y/3Kcx7gqG8M2J3I8uhWd2
4ptH0rtjsao/cRh8V2k2AEdNTkzCvU4uuvrTvdAYMa+lgEP0R7/47yIZOY+uAbDR
icirIWMhhMSnSGTtW5cXKxV8qZGk0UZL/KlOEa30ma3ZMACyAlu9kFuLfhp/nLhe
KL1RLDtNLLlguT1z+YyyMY+ELYq8Huz9U6an8m1lqY+RzGj5J0d/5EEtvFlo2QbP
kcq7Ox2AdBq2/cqN492HibjxpwTDccceGDZQlNOwBVv6Ym6HDEP4P+MaNW9WW0MF
RXk+p1e7EaQJKqqe6UsNbPcE2Pxmv3gOBOXN7caU3Ebvrzt6FFwTUS+1siNpXghT
ECowx7DcQ17S+iU2U3/i4gOEw7q9bN1b3wn2p5eORlnhiisoMWVabDwpMnQja43B
ZL6abzP1AP4+rj23SKz1U1YFLyNv3qmMBVcl9gCL+7MfGenVo9e2dN9BaZCX5Dsv
AghAYox3XKAx/wzWeRpqPXBW+wI470RqCsW4eYyHXY2Z65T7qS+6bbvbqpZAL2OR
RfT7yEoANh3SMO9Ulvjvh6LdsZ37sUfb2c7n6wL8qZcEEOcccYTTTbckJvHAjl5e
cFk3tHxgjhTSc20bfAcy1MuqZQ6V2fz0bBZRHnhRDqTU3CVFCv00iFgGsum6Spa8
BaRvYHZRNBYwywSERPFhz2ag1vKvcxM3szK465rtDYjkUQOwYX1+uv2m8bQDmzkN
iSMZy0bfzk3IUd84HT2cjh/UbqyxCjqwweeZ7UU06kscGQFU086U3gMuocxuCp8y
Fvl2LpktAI9L01pz9+qBbPjYKYsh+qkz7E0J+eFVG24urLTRLLHtm5S7Tv3tvjHx
6gcxzQE8fvGLFEeI9sDQ0DF4LU5+Xx1DPw7VYREyYRGxZONruNb8qnDhT3oE1jET
CQD5rmtJEvkrPE7yMdHL1kni551bB0oMfcwAH6g0zHTEdpaeLl/XIBVvHM/yV+nc
I9nqTPZcGA0tL+zgLvj9cDP8OBDqBEk31ackeZAwvu7vtquFbojxgSf7ghcRVbQW
2n1lnVH6uJfl0xIDWrrnDvcS49CPS65zE4Uh2of9FT1A2vjCIGVMdqbzSygQ5fNb
ZQzL/5cGj8RYGcOwyTDIPLN8ED9t6BTr83sD6b3LMPeKloN1/YgWvfpwMrEBfvhC
xQaDZe3v+56xtKR2iyp57/3LJJKKjNlpDNJ4CnAscM+mI0U9/1ezfMPACAotKmiq
mtUYw03Vir9stBTk6Aoch0nM+QrkvpPZaQNbBISljzMt4Npoc2Lm+92HPr6AaEpi
nrT9Oq/WjkgPlGehaYe4hZwRmfkd+vVXWR2h3Ld3uffaYh4aBJLSDqK3i+aroOO+
T7hZpmeFyCnklS2ECAKZSoO1v2oxFcQNGNojoNGCejC++FA9HfnrDJBwE0Ie/kX6
sSNnanC3sHbp7AmsPQHqzYJxqQMQPX3Fa6mxDefVPV3nwpvtTaqyJ6/0GZP0wrzu
KAp6FXwwhrlizV/0v7TTEGPrFGHDIfqzorvKV1cBSLOFEJwmIB7x56gmyaRqNlYo
0LtFApELE1j5FSz9JWCnxBxyIdGejkmCMmDKgY8Wx9GJKjexlRUmVvFUMgEtCk0H
rzVXz3wu7iXk4NjGlcQxjl+ovIS8fIrGanuzu/9BfIWsIHuzyxIs6AQWTl4xXp1a
8WK+LwycSvthHm5IXK9fA2HR1bXc4eSClCvYDqmz7dPk+1/zXIBDxZy9Zjz7UmjJ
0FAlzFedAILmRsmpcwdQBRDP7FP4ckSf8+o1i0NzTKUJaJuTdqq3kEfhGI+8WaPk
k92UgnWA9Vc+Rb2PYIuK5h1kv+qfUfGXZFRusnX8ic+Y4Zxljp7DPvEOedbxNAys
8nvxL+H78YMsIemcO98JrNpQ552PV2jzt1u1TfpMMvqdMCNKNOk3lSNwgWvZlI4P
zCWiQwdaWPOTyYXwZjqUwNz1Rv+PYw47+GREkmD8N18hGYinF/3FaHmbXheFbCfO
0WIC7SnnmgiaocxGAnFKN/sLPHA+N6QKuBB5EZJ9mMAiwmCiWS62MSySS/lry5BV
8eKddYSrJ+1VPSV66/e4D0NUvgU09cuKRyedldtR7hkJP+5n6sFuOwVBQA+7wmMj
YNtaTChUdGFl7d6tV+94FhxjT8khaAHU2mOldCXiN06m2SYYB0uAQkf0d/6OFq45
9EQMCo95yiCZ+Z69NllfXIOsl2EoFsliTtYrBdqEzbC4MPOdZ/j2AzHDwDe29UZi
q84U/vS9saJQ5ZLIr0SIkJJtggsdUYEMI/Ll1pzKUVXd38XwoUJWoFMB5uVC9Uj5
vbzvdOkrhYqj8cpTHsNFA/xJXDX0oSKLCEJ9qucK61uTdrhlllVo0mMpyZxksUUF
UwJGxqAzygo3RTLNKzSbKTbXui3x9w/FhmdVxIJs7iQl6/96i0cOz4RmUtea268Q
4rK5gdcwDlkgm1bx8QyToK+ZOML52NSlincQC9Ea8aM27/s/+Hu7tyG3pCy62Icq
EX5c94WbRwK20Kr/tte0biM7RzZqHrfWyWOvWSd9aoCX8K8oyjvn01oqAQJDQDYh
zKSyqDxCk4S+1suDWtazhSMzPuNuu4txmc2SVCseHHPT3u/hHgLtDluD6bm3f3yP
N4CJNvV9jYgNP3oeLOBtv+r9KcBfaX21i/51/kazzFnjdzJhs12Rzy1zoeppxuVL
EKtEyviNFebB2V7tV0UiAFGd3TthpNa2hHTm56gsS5A4JH3RjysPW5vwbcQvTUUz
ZSKa5pi3vr/coedPGWcS/PVky0ODB67YM6vwOu7uzP+3Wooh8axvudFzZLBg8LkV
waf+WurlQZMZj3LfLW7jbqeylnsAthxFXAU7uVKchLXDGNhhAYCAQREVxehkx2X2
EUxwy2vKYPuVVMK1uiklyfQnptRVaql7yWA+m5YCq887sOICaX3kMq6c+mJrKUPa
IwksTmrlDbM4xqgkbjsBWjLvXfxMws+I4sdNzMLdF699EYoS4DG2fPFIe3KNbemj
VA2kGPMSFb+3wG1eQARmy+tQzS/KcFoZMY3pQNdrr42KkM/uLSa8tFkRYNpCyWaH
rCfbD835SN6XanqI0OljgRJ9byw+Fx+rfmmfucVdVDW+J3HKReEYgYhXXHq36RSO
PIr9C+Hfu1i76Wu9AxBnpEu+EYHTVxeuCUMj1auSFY+tyKU9XtEPA83yeffWbyDS
CWYd4MBLY+CvQBZGMrFeJq6uVCR1SKqDdClW5shUBV+ir9PM+AIF+xJaFGyu40TI
Jqp5nsjbz9YrYJLOTiVqlLsP2IFHYctvRx9X7H7GCwl49xeZs9UrybeS6lL2zLH7
iUiPm9ZrkhH1ruMBW53nFj8X74zMvpoDX7ovHuaTsUlMS9DbX4xV6RP5W4f2DUTP
lq9qZks+u/NKcxaAsw+AdvB92ARBFE3h1n4nYjiUsQE1OAQJUdcKN3G9YZ0noo7p
nWgf2KXl7/8cyOTIF+QsNeyh/i0/MW36XrsomYViohbYDHKf6MKO+cdze4d+3F3m
QKRpgsAzXE3/lYH+V3pfPoWnvqKQ2WLcjyZn602FVJumbgNZrwLCMxOPPLAfb9kj
RDyXlcn4QYsLjt0S/BHpmVm5CQQgblx9cIol7MCh9UDwXRwcjnURXG47AYJJMynI
yWMxYBWw5YZgSytzI5FDBM/t89ymV5v5FhpXf+1KmpPuIMVyqCHTDscyMQID8hiq
BMJASo55qpE64DTRvwhfUDnGtRkutrdAoBjtOeEOW1Jn+4pfBybVTkwJdqVAhY8Y
GZEArgAbku3BkmLIah0l54vWXhFAA3LoI5YlMUk7R3ez1jROtI5fLd5O0ctqU3PL
ko1kpzMzwUa1JG9wXYoe4goCNe80SR5sVv1XZulVIA108veURlJwWUf6tYZF6H6N
Rvl5RldbC4M7vAr2B8sgVNngFzY04QhbPzzhD4LhelMyzZy+vVR+u9aSquVY9NEz
7jL+i1DX+xopvcI6ZPmxzSN1uQDw6G+njsjT/Vv/ENtB4Bw7PAZrDIL3gX6+Pxj8
4EERDyHYP8OpFo/+RLS9K1+Ldnase2POrbPPn8jitlShQRba+OU/x09FZ/ojVX8E
3eKkefRM67HyzkBKHj4SMTJyEZEtjsq5Q4M1ZDzs6AVEIBASDi52VfEE29jzW5oa
5ynMNP0rpGM/D1Qeze/nL9a7XfLz69ijQsHHtlSYmlfsXuq3L5XXb49loGguVCtD
bC2O2Vo0j6I+TJ+s9j2UGgGYwjjmwG2Tti+B1C7e6JG8NA9qiZOOlE6sNj3LZN/H
SE8170m42t/akgHmBUw+abdCjXYtcxdV6YT4u5OicEAUpnfHCfjyvPq/ahOXLKjq
ViESjJwAZ75IZA8FqdZJbln3wLoI78ARkuRynUA7WX7D2m9cw2GPQiBGj3CBgaVx
NMh1K9K77U896hMSrK1cKS0pXo6eGnfWQnTUP8E42Qw2DBY+fF0nGh8KOZs5eom4
SLQMZZkMnE3jTLKocN+XXZUyKWzXzzxX/l0rfNoIZXl0gh9VmK30hQ1KJAwq8WJz
0FWVDOZKB1cXSsYKxYA9M/7uc1AQkxDzUkg4opf7nqMc2Cer30IYAIwyfhGI/EAL
TuYXOPCw2CPsjOG0zQGRc8krdXvDQohnjUCH+D6zytLTtjCgNeKVdGU7B1/ipCNN
JGzSm1DVx140k3ySUBDFKZp28yTgbChuW+NCOce64MhnzpfOWQHDVVkWROhe2ON5
4TRWzYmmh8aUcRC2xtJ9tqpPiPASq72iTQjuZcotcLn6XEUi8qu8PtA9pZNz50kT
y2WX2ZlX4YTKkFMQbp8gc35dlRYsFYFH+d9/pnZIWvUf6gYyDo5kzKx8iwQVI9us
0q2aC0Sp419UjveO/X7whaQGQsS8/2lELB/XObZQGgGiO0GowPkhSFhzxC5Zaj00
9hZsmBDMegsIvnUTWTYeuLgmmuxaIfPGknifRmllKYqycA35AmtZrAuiJ5BJcQIa
uyDmv2f+TfWIQDQhAaSDimcKncYeau7cqVkKwua9mht3EnZszNk+jKpoTqW5buTn
RVS3gBe7rneirZOYah5777vMVFWYZKfXZHq2Jv0/fOJceChAVYfRjf56SsHqhl6u
jNb/cXmbsVLnRoibvt4a6+Q6d7BcWH5mAATMoZ2wRcwKhKXGUqs6D70PvpTk/Xx2
iEOmfPUB8EtYpTfSTu4mT7A7/+e6UroaOaXEqVxxnUHWlrc7kvGsvatDS49DiOUZ
qgh2U3NV1hjk+KQS334A5mwOCubzkfIaPAvfDyIa/WaRbqtFadOlZ/o1sz1Bt0hy
rpWyjsPE01EgmxrDSDkBW5pl60QkBhUtZ158Tur1tgqya7rvyu01A5RJ9cOWGmHK
SXnZ+1cEx5wkt2ApIKe+aP83qcTAlxr+I3N3DPVajK6m5Y7s/wdu/CxVLGJmdiYZ
IbpoP0z7ouzxLjlKnadktwqSPRnh6sgnz35L3g2oWVu7QYzDHOMq75Eel/SfVa4E
iXOUn0ysdhQZXgnUbvWsClMSeOnixkf5mGnQGS59huGGRcODarYLucP7OdbjAoHE
64tcC8dPpNIQ0fKN56Y1bgHFrKPa8wRLIBRR0MFLGBqDGvz8gKv+RpB7EzotGqrl
MkK83UqgbWt8mNSUhkYmYfYpZ57P0byJo7LAWYhDRR3BDco5SFHwwfLsHvyKSRXc
vPUo0abAjZvJe+g6m0XWakmzsSQV0lPkZPidV5oZXifuJS/TAV34Q2FmOVdtEHdx
IowjvfLzh5B82SbZgz9vPtDRz37ewyQt7FvBBqeAxKL1zvmwbL+Jeu1V1h+lY3wz
ypm5FW7iMNa+uYs4d7P7TBP6pdXMHsRN8pW1q7J6DLiyOeEfAI9z0mKAOrCyG1c5
fsF23J7Pn4CawLRSWsKjtldMt/9jBvGAHtEQFZyM99yFvUwCgtL0bl5SuAuAmUBe
tBaFXkQNZpxuWPMrLjYExon1JpIb+ikM6HL0xB+WAJE/3vWTiZ9Eg8zRDkQLEpw+
MnWu76/xjoB4QcARBcrwokkvQXdUptHt+SyWuApew823lZgM4AaCPrz7Eo14vBLu
j7bdR+5r+ibzSboIPIHeJrgxxaU+eVKOjKaa/1k3d9tRjkFrcGn8EPEnRbrvnjm9
8NU8D9PbmoEARPmkoPRh6WmZ24blML4BtzCWqlkkJxvlrU0AAJ7vqsO5gHrQzTdm
JpFyAXh9R4MF9ZEu0okzSFCNm1rU1UgmsqpvbJi/eD60eZbHHiGEeXOVnqHcI6Yo
hi9sauGo9js+OexVaWv2jKl0pJ1NpcN/Z/KtvP06Dl4=
`protect END_PROTECTED
