`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ofnj4mITlyy9sLtL8qmUACXA3DdYAxSibT7GS6DqMtTzFTTagooD+2D5/MHqYDEM
5fp/qJMJJStPu4lSrgpHRj9iK0Fg3EHJtSnRDec/i9HRoxoVkKBjibAs9Qxo0yy9
wKyXsnj6Shr7J8AHTmPcd2xyFHpmZ4LmkIcG9hm1Jss7cvb2g1GgmkZ96yMKP6B8
T9voS/DVjR5PIvBbyOFC1n1/uB12M0PzbAc31Y+WyWPEkvJV1mkn9kXof6UcxDSc
bpXrX+pX922fidsM3xX1Eh4ARtyObjkBYH1nWts4i6kATI90MHu+DAbx4Qr5WP7e
norW+NQukf01ZC1b/Uoc3vztzpt8nkd38RpO80wB/R2O82e1godkjolGe3+5avd/
J5g4lneeEH+PIp6OiK1elLeXJyDLT21EN4qRNKjxpm21gx7z4jhaC+Cwq+4EjUuB
1O2Vi9uete2kDjCYbgMzUCHIpsGjnBiozphg6tAxsnMCK4CDilVxMgEnreYyWKFr
wa1XJp/Wtywgo0D0WfD8REKEuDzV9Inb930gaYJvOLkAJHf+uPlP6o7ybQB66iZ5
/4DAS6Ay2FJkHNa2i/NPfH8vjipeaC78zMvsbbg5d26Wj+Y/oqOFHohfkitBQAPQ
cxwvkxRRSXB2IFViv2dqzIUoNSHGK7EIA6kYOluJoJQhhOPA9IL4A3R2u7wu0Oyr
q9li7dPewd0mttosutLSv62YuZth6x2j4raTYv7P/GJOCWoorLngnrRNjoO1S83W
KEiUNbFmEEgvhDFaNqmyFDpb03+0ilQvMvoP6LGa9HeAGZJcUpQwR9D9fMwFqvvE
UE9toNeYOxg+PFr6wHyIRgsPkCPTibEG4VL1CpYwdV9hIKKdYdWard61opZ3+G9T
tkchKv2mmzj5fe+8UUEx1oh1QC/vkhk9h2FDN+Nz2jw1+pc+0Ja9rbkk9hOj57VN
Y/uR2gziMyikx6Y+sv+2hOrGEnUXOBi939kRbK9YZHhEf0pCX+dAs6rdqCBmXAag
PF1QivwBlCwS+//aDaMeZNWu0X07ZVCOig1MupPZl1CBZFseJ2bhacmqb/jDIS+I
ummsPxg2bBpl91efeyRnePRZ/14hdW/TbbkrPqT3u6L57CbGdy8mZMLvOWWBTYet
xtwB3w2umw32snhDIq44ZytyhMslr8BbaannXkoS21ZHYF7vBw5G6/csEt4eZ0AV
A/1ri8+J1yAUH3BOtaq2ZglgBKz8xb5WY6JfMbUsxuU8+9KlASjgwXCbdgG2FzZk
Q+8jEEOEf5JOxJ8teRmJydSy+MXqI7+iDejk9fxcuMMriaQwNWsbg2uOD8nQ9Ocv
vOjuytNEwi4ZGZ884Sq4QW04ULFkDGfu87w1KSkU0u/AJOJ2Ei6McPQAs/eTOe4Q
+4krYSq1LVr4QmLPl1rHZUXay7tf1fIt/Siub7ia6x9ZSIbFF4Ce3S1L45sgQSVj
ALuwhFoqTiPRy9AqZZQUmL7SrVoKa1RVuOVHy0Y61sY2N2Y14p0GxOx1tiXUtF4q
Dtjla7hthf6jKP4V/mBpKhb72Bfql/caE7x8uxZKdlIC3gMqkYrdMINT85qkr9pt
WejpMfB8kB+bXeyuKhST5rrgvaZ6zm9C9ajINecKnNi4Cuyk9P0D0JQAUD5SBYUB
JiGQJ8Lp/VswEl8EI70q7ijTXUzmNgO7kEQDmxlvEoVPjDjBl6yr+ucytFVnoIWc
3fAH/7JF19aBCPt7MkwlhZXNSxCsv8CshGrLkrXFQZZfwv+5eK9JBdfu656yVPdQ
3yu9ji6uO2K7JXnInjCP0WaTsT/+gmPJFZc2+ZI3VYM=
`protect END_PROTECTED
