`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pAPnEDsEGv8WIcpRxcvloE706P0SsrlLaQIIJGEdo7b25v+/+QZdCeW/U7AKVTzl
HmUjYoTAserfyTS26HP5J/DmbXCTCMjk9G/7Ge0lZxR3WpuVKBJRPgh1D7YyHw93
UuwkZkZH6i6mTwqvvIEuyUjnARBMahVr7zcUTLNYQqhBjzA4SbSC0x3i4J31I+NI
tA5f65hWkUtcf0JZYnqMdqiOtVoPN0V8mFN5j5SlRCcGpb+Z0iVELhnRbqhJ0i84
FmW5us1qoPjsKNQSvut/JZuBC46Xvn6a/AHyryZEI77S4bCYKxaN2dtbOzi2C0mT
cwNa5h39WzAF8jUd1yf7RrNEbgvQW50J18LreQ8P/72kCl0WeRcj/pNT1V2SEg8C
ZYWRex/WV4O5GeQDOXeh/0pnlcTT2BhMn71AF++uSgMn60TRxloH7B4gaaW6O9p1
zOv2kj8OqSyIRWEmxZGtdr34cnAXc4Cdh2r4opbOYvNpe8b8KAunDmHagCe4St6S
oZvtyiZgNrkxqBFAREZUEPDozd0DQI1RGmigmWJGZfRq7zWwQKsQ+9mtNDLNB9VO
U2bTnephu4kB9ka5jN/Mo4EHUOUlX8syU8zUGXaGSxjkhLB/mtJem2vY2wIlBLpI
9i2dLeVkWd22jsi54hTm7ydnwwdxRypNc4EoaamjGAV+k1j8gWmIBugPl0xzgHJP
hEfC8J4hMw6YPnBLd1KaXsHSdYiLQYnDwo/L1MsLFyUe3BO2OuGzWru4QZesAIps
TCqrjtELWQrNVrMhGmZCecwSKKOMAQTOoUa9Ld8/TOs1s0fTa8/8NYgmKn//voDS
OWIgFOGxtd8BkbvsXHr+WNuzTJAQJLpl9+NbiRKfx4GjrEUFpgNaHNcDnf6gvNaA
PO6+2V3cHRV80CRxEPHCJtuoKavUXr392IgU9MuMsPXPC9LSFHx+1wjLDyvBONiR
BnlrJmlf0RxKE4lu2XKbsX2iF0sQsifJgVwAxEvaVsX5BADeOY9fHnlpUZY765ml
J7HDA89xEclTafh9kb/qUKf20tHBJruwjCWe4Z8RZdpU9lmYby3bcTKXug8YaDN0
w/H7nOujdwhJ1lGcvcI60n2jxu0P5U/0nAfgT9vWzDvl4JwkpdW/UI8LURWgPwDY
OBeZsIQN1I2KZ1qG4f+KD1fhjprX3ka0lCtsped3L2mAKYHDK4Lun5Ju8YQJlHho
zAfEOcZpPFfQuZLNB/cdZBaAksqPtfGDxlOt1ZlZmz8YCr7BhIz3KCKmziRK4+1o
`protect END_PROTECTED
