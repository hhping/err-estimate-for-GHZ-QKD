`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZYaHRzim6m0y4kQadDbVbu6OmpZtOqQBJBmzs5hbmFRq9Hx3a1HYARJuaRGNATFZ
75Ku9YlhqtmFCVcwyzItpsKf0KsGwtv+xNLQi9V0WlaBlM3FBXrqozCOuw6Kt5en
70r1GebCv1FHdAcSYlAnKpmonxAV3Fm+fiNPsKl9A1sfNeKuv93kzbpxbtPyEDuI
3OW2wifS7Lk9BKRk+WeZzQKE1vR7HP5rFRHks8O+0rG47d8NawNSWd+VFPi9hNEX
6hISaT/+4WzkoZE/RluBFuulj4AzyGAGBXDcJrfTLCeLmxjg4OVbf8xcEEu8dDna
a6iDgWXkZsjQWHz/gHXcswGhMaMeAln7qdWfH3izIUhf/ppgrTL1pOdu2fRYv9fg
ThqB+/EZnFEQHbF2ZPKm6KPtsZwoc0OmTL9xooL6+BO/MO7H/NVA4w0kEUy7bhWK
G4VDXilqfm1IMgiEr+tkab4TWuNCYmbfkRAJ0TtnGySimLl0trCBArR8rJoMgQyK
34N1K9Rf9VpnE+mK9qYRCn/nPS33286wz6zZ+KP+MqFEiM3mlDal82rLmkBk5X+t
G4/dX/RH6ESw2Ek4JIGOA5MGTgX2gyvt02I86GtzpYtU4eqDdnInYC5T1K7KvVBO
x1UQon8HrgCLQdOVTH8XpycMOpc50TfVnjmeQYbPeBNgS8X4tYh03v+dgng2fq1N
DS8nd0veOJfmjQbwv6Vjn/50IE65tVfc/1rXwq69WXV5jjmTfsgmgBl19r2/pf9Q
LyJONA2iqnGW0DCi8eR4j3klcEsBs2zSgf1l0DsOajO3a+2u8vZatB4w8vUYsF2+
rxhvpvcj+n2730wv6om8mGdsPtx5/O++GjwKNRGDgrq9bWnbL9QvaFpcLGwzsv/g
QhR2dhBjN2UosfMVCJVMA57LplBPiA3ONhzya9rREM1s3lm9Nb/5fqVmbHTJoolV
LDxZS/NTT78NYdno71S3fF0AV0gsKatQXPxSblyI9eGGn3hhwMQ/qVwcuolTP+VC
6xwnGqq29oXUHf5efM4VzCCBqCI73Mt+qQ7Coz+9zYEHJfGpA1JZ2nxtVA9V8h2v
VZ6W3svXSl05tF1tYzmXviLRwp/eaSFROxT2UoDEjCHwntgUf2+Cwuqw1HgGyCyc
3X1B8TyxoOPVPdMxLF9JROhgSN1B0pWUDMn1QdRlJkvlHNRA9FhBftKZrlZxS+GA
Qm66RrB2cxWipa3F9gE5HHn0zmKIQ4Jg3iOEyYVHCJaDFmht8VpdKFvUZDcu6qwd
3n6ySaJ9MPdZPDxBhRKpgSc6STbAmkklOIl1tD6ZAI9O6yMDBA6E34CUqqCuaaVw
5Ts+rlfrxspKSZfZ2C5UygQqDn8AcGEwPALRlUTZ9z0K5CmBs6PJ25iCErx4eoXq
78dydWC9gzsS3ujdtWnZmSXIIrF3d5NhGmArZ8pTY/HHH2BBA7TkwlL7qaXeSZVv
RDE9e+R+P+GeRRBKIHLB4PoT99pR75DMadCeHeDyVs30dVDUNcd5IbZ+Rwy8w0U8
O5YpCyaMvW70Z+WyuFhp3n3QAE6f58QEEYg8AmpxmGaHCE5CJIGDGJH5BV8GIrcJ
q/B0WhijCT2Pi1r4rr99V98uxYQBc+DiEV5Da4W0wc0GHSctaO6U5RPcFtJMyRej
V6uaSol20GAfiS8Cgk/Z/RPYmRZZPweFHtCUXp9xK0kJP/yau3zOvM+Hrs9r/JXP
WPpK9AVI/I9JFEeFo2gd/NVxuxbuTDR/AEppS+hg/rC7t0aUV6OzjVE7jYvLdX4G
25eKDC4nyof1RXwfa0VHBvPn25zPW7db2g9s0pzOKseC1n349E4AfprgD6FebjQP
zOLdGu9TjlumiCQXgkCrQZWbNHwbTJUC08opG1mcPP5npPiUQejzXZH1nm3MHpXz
V9rKN0C4xSEo8XM/d4xbr1XMw7s7gvz7LW4kxA2Jwso=
`protect END_PROTECTED
