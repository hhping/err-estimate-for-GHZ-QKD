`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dS61RPDtKUJ0kXVxO9jG0it/5eLNHxz5/hiYo9PXPikKV11jGBdMnhUsgA98gCL6
SNXojzCoLze1voQcH3rJfHsJAHB4FfLt8F57oGquNs6zON5g7NKWu5CVnLu/KQuP
RtKqIUiUgoEEB+iSyzciaHDPBhRu7j6FdQmu3ovzFeUSEjbY6W0FV1vJFJi+fonx
IA7RqXgIy4U0gejT85/akTj6SLSdp9MCVPLFtjuu8OK/ykTkqGTIVPevnxivyTYz
+YnM5dds5q40WhqB6Ki19nfC0+A9OJ5rkfPZAs/GEtYXzhsLy5XlxPCIKxDEHMwK
vf31PmX4z3y5c8AwIMcqDqaqKwLxXpLwLL+Xl39x+XlKanT5FqC/roXiJWVFSVjU
WHomDoigkY0wyNXvtYhVf/jpFXtx80O1IN4JwPpY4yU79gTGZ8sfK6QQV4mEXea4
+Etxvpi4YTalbkSwBR16B7oweKp60Rf2okIcsW5YoWqj38MlPYaW0jHRSNL5TeEK
L4zs3Ly5s9ZvaCOuatszcyOG+spLpp+YGqV8xSkSYBY5QhpbuIyzZ+mLAxx1eQLB
8goq1zUtxYI1gdv7eJRkC8s5Wzn00ThWEJ13Zr9ya8rIvWHrI1mkkPLrbfwOTeCR
FEOU0g9zXYjSZz33sh8GfiJk49QkA8kUJlIWikUARkUY3RLhjTqVVlWBEMHVMGT/
XNBi4NuoAMWvoKt9GkRBtfMuCUw5ez5xCB3DnYGFevaP4ZlDad3dBljsuirEqBgc
IXyUN5x/xwX4ui9d0dT/WTkibfcGlWKVEFH5sIbZrbrV2FuNeVx1wXjEABv0Z5kO
ZVQhZjSjkk/o3LZzLX7RABwHj2qfdPb5qNKWJfidjYzBkq/tftVOUNI+w9sFOYz6
RVRON2y43TnoXAGrk/OJv5kAwvUyzDr3324uFJshG03fJbT9cMj1LmIdRGqLudOW
bbsPfU3eWTX3+XO052K2Tm94qPXzDqn7Cccs4QSYGL6hZLpVG9lPfhgAklb5xusY
zWWqJWKc4uXm3twVugfKw4YHCzNFv/6xYZo+85ma1uMEgh2Hbdu+NchB80ErtufN
wZIaNTLJlLWBkQe7+pgwGXBEOmSxXUJRlBGVrJkd0eRDJ4weTaY0MJ9y07TKoEHU
v6I+GgJeiIEenxQDzeGHvOWGowEXqXYplZzxFOP+xExoZNOJM5criZBvCSvBxae3
8E8/aQFIYrkbZPuC1gOU3/BDqHRwLJ6BZytUwZk5Lj5ia4paxegU5E9wJGb4x3+o
kAGFwslGHdByGEu7TQLH7FH30YKgFKxOdmZeT9wGMICi+C3LG50W9JcBeYisY9dv
GjcmaaZ2IxJwld+64Hv0UjiKiR+eAJtSYalvJ/DpwEfWDrGRIVSzZrSJXoMo8CuQ
Y2qga0SV3e9dgTEsJJ/mxhjLhdu/7zmSbG0KWfrwiNNgnQni0wl8XC7TdnVkHJwU
1O0quBhRqhfYY+p0tRv9Gg==
`protect END_PROTECTED
