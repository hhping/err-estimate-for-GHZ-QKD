`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JqlUSTK0H5OYsvU5aP3GQdh9Z0m1rDlv9FQrbdise0RVXx9mAB43+2qgMFSQluIo
uS/fLuZwgkY05cgT0mX5oDGOp6k3o1X4BdUjh5P3ML7Nx/eqfik6mLWvfG53J/OV
dlinKxfvBrA+7RtWGIogQOuDsY0YsRWK+cGL3sSn/RraDntu/r0J4uOkBZhA2GOx
uwxkyXXhVlROFS6xdybJZOfbNXdzqvx6UbrB+Ou/htplGheyuEgOmUUUsG7zV23J
lzls8Gf0Set5ZYNGdazojPVVkxjRKRDa7+mG9Fn4AqNdUiuuid2kvC+aLjrLCF/b
8y4F9SX387zaTykaOamOUJiSnx32MoD7/sgdUVkPftV+mmsJB6Kpi2J+CcjcAFd4
FngoVDsqF37cgP/FBatYxM2IcwCrHa3jO1Kd4u5nEr+gEk9BWc857jHhIPiJ5A6L
7JqNzBYbrgcG5URewi3b14ntzOjYCYFgmbEn5yxev+zZjeDyEyXbons75qSjdNSN
KpKX5bdzmRqDcdAepbTQdiqfFs7dAuY92xkscSWNBcYxXq8kkDc8VEDOnP5WQ2/U
WFqo0zqo+8Plg0UA28eo1muTLHTLvqk+P0QeTfq/O6VW2WCqPsjPPuP76y9EV1FV
R/IWiW2PlJEgEnoTgAJEcVUXux3X7I8qO2KSONtab8bdRoOJtoecu3t+AUZFGisl
77ILxAsXDYfUXuQTQAOExEfegxtn+Dgs6WeJJhKnrvIgqvo1yuSTX48RYxobU52g
8hy8uIwXEfrZB3Xle9k87eR+TpPbyofabi2TLr06PbMIayNcvp9KYyvCY+z9ZWIm
`protect END_PROTECTED
