`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xT37c2ixBGWMMqD1TZT23FDk9O+TThfe1K3vO/1agjOd2VeEv7cNc9g19EDljJe4
pMsKgogdeydTjLGKUPIESdCyG9OHXuQfQhhVg0af5yuRZ0/2bVAlkvl8/xySJc58
8uQ1Xai8WL3JleXLwlbEgm9oBxsAtzi8C0W7V6jFLQfSMzCN+HrccAujMU9eOTJl
fKwrcDXG0Ch92am2pZMQvchUJ3YY4xXTTh0FXXLKeR33jC0fWM0Wlk/cw3S4gWb9
1ahLUyuHH69Bip2nqNoAffSH4A9zznhBK09d9mkEvE/Pt9vT25WIwXcpKLmROPqQ
WWItaNY0PKAJZopS2x2Q2BIQVHfcqWWaymtEwTp6Gpm71MkuN3pe7Uyf+HqAmvPB
S8pPBMFNEtPd26fjNFJ8HErgnS2ktmRXZDtPA7nRUmZ/9DAKfAJdf4kybjUm26XF
DbRnk5Q9fUUbvARY4BNYIMwdD7SkjAwNgNcu9bvOKjRsvVoy2881EwGnk4ODMTM3
mJPlc5QKN3gzTvMPaIPH2OjTAkg4axS6fjNrP2mf29s2lVdQKVPQKOTEzR5knU8G
NsBe4EcH/l3OQdIiRYbWCewju521H21vBX7CGxSJ66Qon9R97kqV9xpSskTq96vx
P9U4zBCSeBXppTINLVrzqcG6TtXYTR3c705kNAlKe6D1CqpTHfpv+83j5TRtEooG
VrhExriCUKwdWIS58Y1g1Mj+Y4gFi6dX9AY/GsxIwo4m8w46neW0kB+FDgecNeOV
v8J0zP0L028rgmucBgU5bhKgnkMLBPUhav36QJOwztxn0X61qLejxsA4VV269oIf
dzxmd2r8rKFgkRYCF5OttLCGs/0vsJ+O5JQMNY20/e76cUzSSAAEO92oixULB5+c
ErFjNj5MGTchhh1WUFVa4Aq6mNgiE1rIN3wgrjs5Xtkd1O/BKZzsynNN/qHqnmDA
k9+PtUZauiH2SFyx+J3yzQ==
`protect END_PROTECTED
