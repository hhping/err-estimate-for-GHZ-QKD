`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KxLO1w/pRNlj9Jn8DCArawXhrp66hZgqRBUrXnRg0QwOb86Z9Oy9bcfeWxMSONSa
93tKQu3lEPaCf49L54lQxIGIYF/qLqseEi69Ddo3SXOBnaUTF2Hmzl3gieEVD17K
z1winx6vqBaTDzasvGyYDqLt7xgvrWbt4go1J2C3Jqk5KtTpQfw1AvEQH5ag1eOG
CBVcJRTTEJ+kH6u6Arpu5GYy9V8argl5/PKMxYdDGGFtWA4c65u7zsB5Wauhlxtt
1HCPiHEHSDbymbtcgQ5hvZl3r/M/rGwuZbGClrdbh1rMzVM+swz6m3GC9D63PG4b
Q629/Tk8nWxJ/EiD1XGqRsE0Yxg9Aayw03xfsN1ePqB9sJCYvFXodiV/xMak+Rpi
OVH/T72oHcSA51zhJc1LPCuchIU3EW9by4urjPHE20nGscskD5GtM8Kkak70/teB
IWzDl47mNdjfKx8z7UoNLO97DNIxV2es45PXfePgZpjJIYzR7D5w8nMSMcTIn8WD
HaXN7OAV6BCYbOR9yuBn68PSvUOjVO/isXkesx62ZM6xOTJqpKLGFx+rKPY+xCPf
QOScSmTefD5enWU04sbqi5JUQAvOVK8rExIYpobU64tWf/JwANxD/xWmbkz92P81
FIbYdU/g+NhTmyvCiAf1fSJzt3YbHGoV5g1nd/J0kzgCUTqK4egKwJlbGhd0z7tn
zIOo11BXJLXHdIEnkegLG865VUhGiHljBAoBKaX4rxJeuw8FH0UYVlwRMfjvFRcr
fsQaEGesixiWruvqKzv6d2ccaHLQ/Vgbiy10BMnFUbuojlYYrskYSA3iZlmCL5WE
0k++Fyfdm8CemeS+kIHDz+a33yVvQTF3fRtefFnmgYmxFQlWdJXrbaEYFOFfjvTh
Xmy9m3Nm604bXwCKoyFTeaijKKu7A5XKfyXjrsZGu1JAYJXONtzUqh7nZwuwiAoz
zvB35rUzLbrvK9Bk779gp3lp3IC+WjmkQlMLwtq5gGhgFiB/XrMneTgGTQPIbp9i
IcrNQd3ZFeXlCD9J3YeSTzn9DirtBRbYCmfH9wmlw0j0RgBdhMU0Wh/jta9seU1a
dNgllbbXRbBlghg0uDTKMeFAB8RBOMtvhEiNSerXWbggjNCMU7o7cHK2HwVRxJ7V
CtCNx46aYcqnhbr98/041NNuA11uRHRNPxO9g5KfIAgivMIPPQx13tdMac/UILYl
S5+Xo7EtneaRE0WxNeToGC04wl5tozKiH/pvZ+5UVjRYVImtLGenNf58NhTNiaJJ
nUCGN7kUT+9k8CzASMFBfsgKYU1ou1+Br/RTBL1EIx205ZHGKFO4DJccOvCsXW7I
okm0BIVdK+HpDmbf4wVRQlfEe1mLnkgLVrodXNEcyBjlmmCIBxchB4hMyEhzKzwi
fxfPpUL/vcpOnH/sP3sPDaNskjNOj5F0A2yzUjzpwmEbqbYnRphvlytq/ZDLyEuG
UU0K15tx6u5sVSQfMrzVb2S6a8FYfk0PWxAUGP8ZgtQ8RQoxsGyzwdYhPMUWqizv
2cx/v6Qr06SFAzAFZfyMfBYwB8rYlejUEZvIxzMGzQrcZRvPxWJmBMhMA2FeiPwY
rLpFxD6sJRz1e4nWM9x8qbZzarfsu9j9OY/nADEc7HUd37pYQFVHnFDyVYWUA7dx
LYsfQd9T6XDESgTXUTklQHMhonQB3FVCN7LiogZx33XR1j7ZZQppGOBacWTz5JuM
4uQ/RLDEhOoSOTBtb5WrZMUeLbuz2xXDpMGuIeXXaAUwc9btLGWlo+RP+FAKgW/h
ABdr37SxeFDUBoKMTvZgNLSSYs2GSK7FuTTcC3iJ9mga8NhAyK/cgT8SeU/Jijvz
mk1OjCdH/X3lqIa7FZ5uw2Q8VlNbWaKSnxzmQPYxp24nwnkVWoiOi1nSGjlFo+ZB
qVU9mqZEswcdKmVbrwV2p8go2/Xd9azvTnLsEX8yYHEHL4hJK+9HEmp40pJsXdQ4
g+WBu8MWBLQvftM83g/HD1CImtgvIgC0JEmER5ZIpIxkCNJaBYiCMZjCol7NHP6w
Y+cOWhCdCIrAUPeEEFhbiD/9/niWCdV8AkiGYZew4vr3czsL9Y/7a+g3XpCKKVOn
NhM8MIHKEik+uzT2701SZTdN5sMMwlP57Kf7SKu5UF3HT/cWnYBbUiUeqGLnXx5d
VjSjXXJXbG4G3JDCBQaYFjOVqOEiLo3u9BiO8JNryAsKMVGlQguwU27SpJWnXe4U
W5QPLuUJzFyN52SNWZecP3ilmatvfD+asgw/86xxulZYNGRuK8hBXYBGdmFaKqDz
lB8NFTrS95ZnnJseBd4iL9+5J85heXOGkt3ki99I6AS9LsEP6f+NSC1rekQAJjxe
JjQEb+LXVlcKXZ4IOj/iSjZZnH4tjSKOlL0gPEifloJqiHJg7aAyne1PIadRwbgX
bUqW2dCvJTIpccf5ATUD3xc4cuQK4aAxS4SqKtqZGy4kuHwe/y7MxLv4cofid2YS
TFWYXdGB5SCKo5tDBTfalkDCmrIcbZGvlf1qjfbAcOINAEiLy6Wn34lcJ+1J94HN
0zIk20MUrW3H6liGYLxBW3AKOShKI1CcJ6TyTVvYGeivtua7Ic/agDabtK0YOKr8
DilebrdscVX0PrL7laTe5nL/GG2Dakc95KhAtXZZ8EZpWAjZs4r0ip2v+eiRcCeK
J6HGrGMSoD1JNd1zRPrmk4x6hOK2iEEilufQH9Q1KPUFrvzuXf6kS/6CTn+hOa/Q
wJ/syMlT1JeqiWm8EUABIrGKQzCY1j4hSKiaBZdsd4dY8KO87CaRxuMLgjHEbzZd
aRJIFv9H39HG9KLUiJANtLhiuIYXCWAQS9p3tHH9CiwaUkxLEDaoHXLeG9MigvI5
8ZyknbIy5lMoQ4PtOi34nnSBIbPtnoNV+LdQ8DaUq0nVjQ8xaFqwvO/wvANNMW62
8A7/ydgAr3U3pd6tONXA6AAGqFrUS3B/ekuzGpdzcYs/RtGBunDM+EROWUWeWV3B
AXbvICMfS99thTce+rQ4xdPZyHa+fqvJYfsbidKaewdrNViGW48n7RCW06qPcP6e
FmXXghg2OgpQ26zR0YvigcKja4E2FXv5cjFvjRMob1L/fP/G+K7DCk3F2INvfp6Y
lSW3LVw/y85PZhysmkMIrT0wqZy845d6R9XXnHAWX0kaNUG6/fMohTJFZsT+5Jgj
ON2E6cTI5lpH6PGMAfrNDUeu8Ysnz2RUiwmagbyc3ABa3/T3Fp7D9IlMiNd/34MU
YE8NRVxXBmYSyLK5Zx5IXHQNn/dXYan0AlBG3czTcnpDU7BRMFy7/QkXpdkCMVO+
OY6DgOYksKtMNmiemWZagV0NNhKk9+y2kKM57w9TIqkAbPX6mHuYDoWOj/Cuv4fr
jkY1GUvwt30rNHiOBuiHaLy4w7/iNmSTaMdStvTHu1X+HaLG4t6TwA2E3V6o+fQ3
Vl/IaS/D2jCGgGY5MKNGVQy9WGF08dG8XLMylzBm10In/6IcXUYwHGeWPh815csf
MaCEATGdfgcl0yy438bt/4bPQ90GFNN/BT+tTGnJ17cg9nzU16TJBSAWbliOitOv
07mNoDvz8DFWeJxejZFIPK/2Xn4gUHxhVIRehkp8sYvOmvexiqfrKCUuEMH8SyKr
FFAqk8NTlJYekhX05q39u+gI2hh9ndCm58kWSGM0ka2iIaELcca9eSqWVj1c3alN
hzYuBjH6DX4lUXvBhv7ZsH7mKd32AzDEZ56dunAxiDrk3k1ew5TboUdiwj9mxzcV
UrMKqrYlQdjKznGVm4zmhKOokljUHQztAFfO6XQsUBmqrEsUOExuinkuLst4RnrA
wyLHTieCJPEGX9i2kf5tlcnWz4nDl3RMVUFo6pg7qCCPs0X1iS/gGRzSkgnZ94QM
6ntLAbjcvPxG6kWwJpinuoeTJxsZVsiIwP7POfPDtBo2TDcSGElGcEELVOagxpCa
wuFQIInS4jFQCOBBVjEbF3LQPyhtxXA/mgK1NIAu4orGKz75pjfsQPtitZboRPjA
bzfJU/Wiz1CEOSciMzssY/CJlICUvFjjePKf4jlwmBCO8GsdGYYWC3ACA2BOfRnv
oGdda3tAUJFPXNTa74twhEUT8kGcQJWUl/k3Oe5pFuMBfmtr2zBikD6qQLO4tfce
76SWzDdCTTGTR2GWgV7UaBPbeoAp78V+oPX57WijLkv63vHuI4XDokrD62EVvWpD
bTsrcgXZoEHj9PsdknmhEHBBD/8UdvSUDA3TPIIxnFjHIf5G/CijpVJS4aq2w2jT
+32LwFc+pj6MogJePVO5pZTIeB++hA08dvd8CSm5zVTxfC+guJGhiNASe2yzUNFm
zemVR0WqIqlpVCKYEd372h73JyggyjY+Tdhagfj0nKAOBWewFzX3GV08ogGPAaX9
FFea1uYpx5J3g9hKwhu/AZBEfsRkEbDHFx7M3bMizHySQLeWBInLXrRGLA43vG/V
m4GHe2a/8+36bsoih9oKWrI6avrFcsCiIEpC9swix6vrfkS4HcglQV/xs7MMG9fi
Zkn6rl+DzBgqbqSLA853E52PnSBF2nTAKg/LnKBfFLyGQAWY57CX+Qd4s9DxskeE
goaiaOd4la+G5IncdXhbQY/kLU2b8QZRw0wBkhZb4lvdhwL78VKxs/Y/PlRMGfv6
CRHEmSNyTgy5tCBg46Ele/u7kL/3shyulDFbplNosS6zZqSFz2qdArhp6rTPv+FG
EM+9vRrCtnCg+wRBPvHrk0yyxhkT7D+B74VCsI1Sxe1G4/lbZixKU7oD9m2QXxOf
SmXIHYyTDx2k/JAB/aVN3nJACKPelMRPsga+YO8k5HZIZBSLpuGCLzq5mYDxSjL2
61QOKbbZ4/lOIR/WbUIYKLf5L6OngYIcx6Y27iByxprx4fK6YxOrBzf6o2gEGuG5
YnORyCUYh5Ss9pIhHD2Ix+z+wVZ2cMR6AFjUL1bXtYOCYs7b//iiPMl7rYRW4ngH
UfiCoQKYVN2vk+zfnJkDdF+8ESrgR/G0ayEG6UqNocGETRuaHFpU2PNQHS/uJffT
xkB0KsnH1aauuS5f1Dh0QM6KS3NVLr5c9G7PQkr+16W21G4Cxeh8yjnDNKxYtuUo
86K59R+OrzawkZSzPpXoS9iINSwLQhVWJG/3E0FVIwIADhoa1KvdqWdeQES5ErVS
acsXmqUmnbx2CwME7e9GQUf3ecBfbnUJaBqB/SAs8W7uW2a20cgKh7EpOVr+2HBs
yQQ3gNXVrUfe+eX8t1Go2RA9aXLT56fOJ3B5y7/W5puqUDnPW1X/sqb+mcquh6Vg
UX3gwF3jaRKyZwiLaNGCXv3Va4KBsmfxWHS+OaOges+OuzlD8j4+2VSU2/n1noGL
YsfFGPWpDw1po7EynhVIzF69fUDqBk/O9FScQLrorqDUEzQB6hLrLrB+i7lEVtZ4
XKekYV0Tgxk1IMeWvBwkn6l7X7KoySbdoB2aSYpzvF8z8QNlETlUoxLXtsmaorsN
ybpU405l/qRmDVOpanZ3PpLK9XD4EXkQ8+b5Oi4RJGDxbFZbIJRT+7m6NPn4NIyQ
ykRdAPbr5bXlppbeLwhJg3BEPsmxrFYvzZbqdBkiEjx5AvYt0hXVJaJjUNxECxvh
vLawls4nDsMa8u6dakH7oUe8SecSeUoFeffYfzbkd2LSM7jcJT4qdaq11Hdd6+36
I33EYS2nIGpUtbFce7Xf+yhMjQhYbsts8AkaePXTlOHXAE7Hf3JR/LE2lqcF9H2R
L21NmOn51+qIRFNNLjooD1Ed6hT2lVrgKyhBUdAHyi+0xXDval/JVGLi6I1YXcPN
p1VBO6QB9EnBpWaKyLyOnAWEGWznpZ1IOYGXXWXGxjlA7DTuKokBSJaCQ6UT25T+
XO3QN40hw0sAjh5RFsx1mLOWedpgozeA8IkoUv7RNaBfBy46LwbOpPIUMf0/g2A5
9ROdcm6vH2WvyvHamR7dDtvT6NbjyHldWBj3YJBYN7xWUET4I1m5bepLMGDxCofq
gf+m5yQ8l3D0aACh6hubugTOyS3FZB25K4kObYOn6XeYu9NPLp558/hq0t9xZWOE
E6THyf9FpXs7nDnUpSLoK0Zn+uQU6KRk8w01L7B59psKfsohfasSc2tE6s01TSxp
UKznWB7cBKQB7bT+ZyNUKUyRFS0Osv28ufWkoubDq3/czZ8bRn/9oJUzqrFrv4gh
5RfnP3ovnWdpXzAzHQbr7GcS4TmhObl19aDhnfDUownuRzM8dkezENn9pleBbF5l
t74tz3I3FO5ydGqFOrW5QhMC6EFuwvR5JB1QsIZlVThCuD+LKALNjFgvV49TlPr1
VrFjbc+yAyUy/fhFxHNJfnP+qHdAP3gMnZbSkjGkO1V7/NIyApa1Ymaj3e68kO4L
yRIMKEhp2Z0qDK65qYfABbFpiGWL+2qdBhrR4HWZe2tQ/fJms2HIU/7x+6E0h1OO
PrebvyU7uv5Cp+tqyOanL8x1I2PxIPEOSQVZMQzeuic6ipEBg72D049IPewi63hd
bDfeAgLUCZF1Ca0My3gPn9dlMw9WBgoPnBn4r9SoGmjgVYrKvxDLnAFpwY8ylpba
DsGUdnnCPhOL6dsMt4bHYCJX/LrcCFSBgazjiQuPmxexiMZGDJQmAouLHGmc3/Xz
ghi2E1RaDsHJRrZWMfxyy7zyu07n4Drm6gTQZSH39rJs888Ft/dfisRzJi9QD7cq
kVfcPjusS/GHItAZdvFtCQe+m1sHNc09eBIGSnjA9TwQ7tPBfiN1FvsRKUNCNOec
WToB/aEXkVu5pI5lfa6Ghmn7N9dQ3830lr9np5NRnlM3qI6Wzmt7raSHcp0eFw/I
jwdUJEwdjE5JV+M9273PDJBxzPs/jCBSc+a0xeJZYz49GEMvypumfjMH9b0BFK3q
x7bP+ooqrs015b98dRGwZWgEyi06xTwpcOZfiD1fakcn8DvLN7PucdmPOWuNdnOJ
u4NWZoD602X36h/HNFSmh3Rx5hTNmTxgaSRKbZojA5rVm/UzG9A1cE14790vYVHC
FHMWC7SS3Z4ZAemUiWDaXCFCM0WLhoDKt5cGaaDNz7eb5vrSOMr9Iy/W5DoWxJZH
yKYbMQw/xfrXiM1vNRPDiun14Sm0VKWeVUQ3dGmprpb6lcXpunHLAXtb4YqhhUbT
hb3AZlk0SqwdN9aTCKIvdlza3XaqcfKcGNXqQPLK5CwTf0KwRxC8L8zTyzm+MuYh
nR5hCImUp3fQrTA2yvEgVg==
`protect END_PROTECTED
