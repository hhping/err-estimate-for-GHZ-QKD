`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gs+Vu8AgSzrgvYiD7VvyDqJV4XAqn3SNMR1LMUmBLPbQg9q1zqYCLOW7HxJF9ndN
gc8x47LUv+H5okrwbmumB3zYJdEkhXWBDVAf2kGmooPamI2ayGJvXTCr/PN9WKAL
8QuMCH3DO8YZWf2HxeTHE7wh1WCyDXtx7MSyaP3YC7U/f/ewxXnI10zY/VO/6aP5
hxO1rSrViQaN4H+DEJimB9TedSRFihbPNWBnEJB1oRfJ+qiFpY7EKlAm0He13E3b
FMYiq5GyD9TTTtXGLdcQMxNPLQRJrhxgVTNO15v+AkA6QvfJaJTKt3wWqCj1nCqt
sqGRussui4I7ZXHlzrtSN+lXNM82pwG76sMY18JnZ/+ep3kpqj4uGpihIWyRwiNJ
KfFrbXKvY8oGlWMEb9Pd/ZH1pebQ84zC2arIZQVROXhsM2UKN1vnCzXmCpaRl7q1
eYkUHAYMIIwDDCk3yhV2kfo+X/O1WD9eyXJA8kTsr7O2/ZiJJzxlCbbNejPTQ1rM
dzb1FsRNGRtOgDZQ2ShEkxjVTX/zsoqtHCU/uHUG5i0kTxnZjQ0KvmkjtDCUTChq
FvILH2xHQj/ipj2ZLH3+gFOAh4lsORj9juAaqju/k5ODzNljKnkG2eg9T12KwkCK
o/JRcFrTtg2/sK/7H0bMI4PCLrUlSdM5rYvMm8zxsNlFqsk5fXVW5IcFz7z0TpSS
7xqGzoLVAsijp9neeEp//JnO0iJEQL0ZNJU6pwNjr9nrCx2eyV1o27iwhOKTDnl2
c+1JKuMMq5gp5BgCM1YO6QoILqO0tsgehHJQDwtqMTgFj4l9+hp4L5MQof2n+cwN
kFiF7CRikuHAwPhARo2Bmg==
`protect END_PROTECTED
