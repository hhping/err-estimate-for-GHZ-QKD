`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
epUguFIXQgqaqmDaEUYUYuSH0BBve/phH6yvIK3fAgWrcQ12MPXlaahAuX2KsH34
ptUdmicpXw4oMNVyzrjlwO76tPX6+LzdcjxoFzhNWSYvHlPhtdy580pWzOVFlWlu
IloFCJn3fRHPyKswojCMcMHU8L7yKdH5f/YrWZrQIFYsRnJVfY6f1ooHyF+LKSP0
xGn1cjpYxpfK5P43MbcxmVoKphijdm3RjqRrB6O6//c55OUaZXctEbwTS0W32Cy8
eD5qiwgQnhUnW55zw5G2A2Cp6LbmrhAdhNw3dMp0ESkTt1f3pYv3LBPuEB81/FqX
6TaqjdY3X2+NBl7nqzO5zEOa3sbqUYApy+AE3IOkYwBRcqdXzsT7TdMj2bsM9or2
`protect END_PROTECTED
