`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b4zOe6m33Qu9K3zjUnXLNOBz2F6DRSY74HgZZrfjxjqKuvXPPYYt1HwNjLGSstdd
LbvfzR+b4HYD2fKfoEhAjE3+VMek2tz37FwfiI6DBEQS1QzyNloD11+hOYZKV7HC
RvVda3xHQeISRP/pxdu2x6ncWmrbIJarlWbGQy1vr4kLZpA3ZNVs5YwDiUs7yFwM
4FC69UdVEW0jE+0ctqbpubEfy2C2DzEb9edB68sBsII+xzFtKsO/VET5rfotnoMw
qwcVZrzBc3bn0lb9m48haAB5EN0CdNRL9rEe42nlxyncM/8cZUQvEjGcbOMOwcTv
TyIc4NqRK00bn0AkqZhzdV0hGPSWciXrJKeaqMsDljgle+1avaYHkxbOia3T7YKf
5FWmyPfpDh1lkmkf1ynKt7XPXsqGz3BNi705wmEH19h0EJGG+2OWVidQJKgrFSQf
uvDZALA6n1sUXpfJwbPymm8eQVoe60TklG324g/OQA5m1kKoUjBH2Io4de6DFfuO
yLumzpAdg+Gn1frn8LjkDg05rW5ET/lQoviDBKjEG4leJiM5Orsidgq6So8H9Qe9
f7Ev/JOvbWtlrgZrzVtBRObqWzp4FxZ36UmDhmiTLj/mFtLHWu2hb7o2GB+5srt2
bB9pc+B8r4s0UrNpnrLrBRlRZ72ilmyZSltDeAnBTZmPQJtUzceO2f6NaKbaEtDk
PcnkADAiXv5vnQ0UhuYoHS+jFkwSB7yL+f424cId3f0w19kBNM95z/Ql1wSuZO2/
Fsr18ysYQgQoNVaf/uSshf+7gjHK18O4yg6bemRBXI2scXUf834OUvpsoKMepT2C
/Xwwpfu5hejYJNLpGLC+G+Ht1EYQEcKSQTRFntXXhHN63XSwiKQz/5aYskn71XTJ
8LVA1sGkqR9Kym2aVNulmUGY38Sj5IBDeFtLSpbjQD9CjY4PqS0pN+ARTNePIswE
9HjcnKLxuwtEg8bBETgzuH9HCb/dKvcsI3l8exv2Rncy+gsptOIDP/r4eKmt8SLw
S1lJ/XL3XGdJJpBopTZFXhXdCwv92qnT4ZO3/68ZwcsYYh3Ga6+o8zWRktnr8cY5
iqgyZoRVInKzKofOSAEIHWJcumtXRoKj9FGZd/mOVu6+ybWaHe5YYLHgbgx3cSNX
7BY8aw+uQozzbkTZ2nQ/91X1Voo4lMBFOq/Nco2FfCVQ/TgU5K89AAv5hfLwmEfT
BJsYBPN9/9LvkHc7gPe6tA==
`protect END_PROTECTED
