`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2r8sG8G4y9VopKggnCPkhbGjID5Uf17uDhFSzzIGOe9CiqqX3ehJO5fA76kPlz/F
07kh1aIyKyiuru2A2BXbrRyHM51KDzPbe3FMZw/ypOWIMbJPoj+le/BRzjFtTAaB
jOcTGRccxAtArqAdtkx1Ro0Y2edWhGqNWZEMeoRYB/QhKxAEhs1v7jquGjsNtW9h
JpsqS5uhHZzEhJIntWAnQbxgWRnFZbsjNGRapDSN2rsmUY8AdjUHjzP+uJCQPTta
9AOOFMUOWccW992iRsFAFABg2oP4wwBgWca5iyLITXuAqbaXOuoM8qk47r449K3y
ByiYWIHgHB0PU3Dm/2G5HB64zSlXC5J7/M1YHXNT+AWdSUmCRtGu7DYKe9QmG9oY
gqLtRLuqOHZSY+Hq/UG+x+ttTdqJ8OG+6qgCzNHxD/ZCR4Q3ZhsSBvuFzaOvoYbs
pqy0Ji1H7s39SClzayTAJTxec8Bqw1PuSpA2dpT8bUBrFD3nl5yv+5KZ/bmQz2Ks
+PY6fxWErPDDG9p0s8Wb5eVv8yzIhWsNYxd4hy7NucmW3/xyy2m62+F9ZafdBJUM
WyI51dihXOlLQC1OS3b1wSeCt9bIf6LQkXRcNaAmdH+bPC1k6A0HaQ7RiX4vlzYD
SMN1I1a0p8Wxh+pQYxxNnKBYkshtRZU0YJmspgMzvK0IJMRlV6n65wVBbvKXqMKa
phTS1JeaZ1TfJ1xc6ypnSG0wBPB8YP7aAIvNpcxDKingIaW6fu8QkP5QUf+OiVci
srkAiqdT/gn6v1QrYxizz6xijL3Vlu4nT5BAbwUyoK7HQ4HvN7nlDkP0t9IlNPgo
3BG5L2v8MaG6tBCn8vZX+ecDQQR342j+BXl6vNeB9n/YLxgxSVdzHx+kSVUKd7zt
nV1t6cCIYCVy4AddRdEhxOAvmIRyeuzWVv8iH6gzlsonZ873oa3e1/55roMUACxt
+arw+O/C9mK0op8MLlYWjtqFR/ZAUmCE+6j/pNo8MqljJhciJwLAzMvluNxW7OZ8
46lqv+LHERmLxTUeau2Ec1wj9td7HlvxyIjSkC2y0HMTLRgAByLmYaxPeEGfovGf
ClPLQC2h5xN0kDUyyzGejuzo7ygyMwwb8eEP0KiJ3LFXdAibvPRboGCRdg2D1puH
nvtHD0nGn3SGqhPw6ELo77oel3HsWLI5VQKWCMPnnpOJyJ+57U5IIpzbBu1wrxU1
7EmGZL4bxXN0IIPR8xZH+IzWUPcbeXcCUA4jA2k937WIAlSdK/ScoLDr2ti8WspV
a+Oq5eGT77IgPanQgEy7MgeOTQVnCf4bGNTFNFkHRKflLPYCOx/wrpmlbGvZ+1N7
dH9ooe2h9J5m8vz2e7H4/+61n/qYcw3VGHvC3ElstdttmsP3uT8Z+2/7eR8dVqMw
3PXVssPECAHYJtvJrwB8Mn0awZNhj+vmqzFi91PKpwoRKxfub0XZyJG6NYqy7rN9
3V8IAOA7rlVoAP0A2KcA7iyCdekIuxdKCUvKbpOt211hokTKUctfGced1mCg0VWW
Erz+FOTz0Fa9TEM3fjXSOe65oKvORoi/TQApAZdxVPsZmg0rM+6OKeAM2sbah01p
yV38bYJpSgo9zQaTSIhMyttDzaIFF7hj3Cm/vsKr1X4m0HQL6l+Rk6/f9RDrZiLq
Jx8HkWFXuXT1qQ22FuFtBg==
`protect END_PROTECTED
