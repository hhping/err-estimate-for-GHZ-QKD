`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JDyoi76MnDodYFP+VW+VvlrOLcOf2O3RP/yXNBlJdEemTPvfslWFYnuLxRsG/c6d
wY/toZSE4qTSWMOU6yZA2CMACmdJPmD4rbk2BMdFDvCoSrfVLY6lfDe4dRBxF4Jk
MfScjUocwCNzvx0EG1YGj/HvfhUzz7CphQC5xiiXCLNi2rAzgoUOW+UXF/DRNw1Y
oZFRx+xwGnlxwlE1TvUsjf+q/x5GNRBF9JM+wVTXd1JUt7K8lH0vtxQlOk4lL//w
s4oICP0dKKAWvAJL7HHKjbAeabldp+I8FOEoIl9vs8cRJU2kiZeBcw7Bjk4nMV4+
ryoOZENcTReU+TeZYK05lBbABs5YWknz/6T7aARHAbmHQuv5WBRq+ld5sNF+rRlc
JbM8O/jx+RCEAvOmvWBFj6z7csBjSFf4j/8Iiw/un0jWHe3iLCAfJhrJlKqRJyM0
3Pmab38z1I7i39eQ8XJTYXDmxsObKnDqlSX13NLNUB6hzZNowlVY+bW3kMfB0blW
Gafv/sk6ktxN9NbtV/bgiLe+1k0Oxf4i7LG9RIzV8CHpWPh/3Pz7sWlE2JjICG0e
0yAP/l6Cnx0SE/mm0JgUflleEq+a5H31vWeTgk8T7bFNlqRdeKdzAla3n6ZzHrt0
wI24+Ip7do3HJXWfEJ7lEacTietiR/vT54C9L4mLY/xwc36sAfr4C90cuSQjk+6o
eJqijIEO9ENagvOcbGagccU00j0pjxCAPn08lQJUJ42v3GDJTHcy5budAwMOswpj
pwpZM+tEDXDhigyZBc9C8GSxjjH79d5Bu+pOfLW25yZ5j2KhtgSDEdOXqNU428kQ
/JsbpisL0B/FtzP2D5/rJlen/Ld0f1phktt1K8wZA2RHJ0+1SMfrJelDNkAQd/4X
A9f735MDXRVNwD0xwGqE7wHJ4s/8HQBB19F4XZMRWOOmLVRWdZfZxGj3ZsFS2dpT
Va4df1Tmlw2hg2R4zOZUrCMhXIzlU3TX8uJlpV2oYwpHhAVaaiIijDliXjg/RxkQ
ihWrPfwbZPOzFyhL/ocSvfZExYNt+thyEQmKnn4nliwk585tLeDz72WBx5/ZBOkT
GKtr5fPHFwZB2hpYyaecRfFMPZZSeXg7opyS2JyHPHjgP61vrgBunl2GrsEL1tG9
5PYWhYJwLio8HpM1n2+0/mRCfNGro0yS+38yKZQPMW+W0G+OAYvrsFMFppxulezl
LFlA+RcgItq76eqnMZ2jWvZeB93v1SdBmGpZKVA9PsDc+osPsMLZfmvOc3zJtfng
wKF+3K4IOhrIDNzl0iWXvon+5zbr256QGrec/mwZZkDcnQTlrG9UbPR81PIgHKHa
2eLtaApzqwSaEAny0YCgkA==
`protect END_PROTECTED
