`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OLis0xRsbQsqSRVz7Q3wTtaisg3YEfxBDodZBy+hmp7iEifXRRSB0fSgZWS5QjQn
bMnSif/qXnmyIewLkJUhxd+UoaaKyYv3bPwKQjAA0eS3DfT9qiMzOhFVNvG6HUNl
4eigCwq8jUPY+e99raF7vL4sMKk80rYlOfPd2Uf7WIlKUtrq7p78n146MBOkvn5Y
S8TAZTU/5J5cgk1+r9cng+WFrkSr2wezWHpPUZDQD0i+0OmB1yHaHTd1CS6cfJ9j
dYVT+IFqTm1XaF75Uk1pgYjy66zIQi0UCSbNNJs/bXeo0CUwfu+4GNw+X+SzUTC+
6n2TXfHFTzzTodn2Rh5Cyc/yB9SbXNeeZnHP73mNNUV4Kfiy/9z7Cpr3vdKH8bY1
OU5sYi8j128tuLJgJWWnEqEeiKaE4FoQwdEVz3B9RHl8c+54J6E+I5e+LMeHKFfF
gOPvITrOL5dH2KYck/zKKMfDoE4zUhvu0YdsrB2ldxRQUfvpvZ9qLvZmCRL5+UGM
VXjbHeQR7OS1LI8remSkvNh6hwycHSVbIs7hzmn+T5quw/IDd/IrYREhXVEOkzBv
jjmsvmSv4HMZfXrzWwy9FmlB7Zhl5ovjzVO7pdePh+n4EqNrFtzsdp7U5CQG/3i2
`protect END_PROTECTED
