`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A6e9hngudgmiuqx3xBOmW4dNmGnBhQHJKJhsSPlLBqMmRhSyNJr1IZ2YTiLEITep
tYDkzR0+jwPgjgbMXNr4W7jZdVF7sip/4dHfDec+WSaNgXApg7x4kz1ReXy0UADR
5urzPb44GD5yaIJZ5xlN3ooVU0mgbjEnwzQ7BHWfZyc=
`protect END_PROTECTED
