`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nFY+VmBw59luqIP+Tphmo/kIviID7p6g1Ak89oa/hG/ZF+0P9Mo+RUmFxc9wSZFy
0v92Bx5c/brAPMSg7H1fDLwfot6YoyiYw0f/90MMfl3QyD+pYj+ENicUPZLX76yM
FslbSjOe5hIwCLA4UDpdlIxkI8oUnLHuxCq3yNsRI9nfGOdyprosJ7YDwRJYaGAt
BRf3Tm5S88cJsWO/m17fObnNOvmQLu32XS+Yy4u6/jLW7aRjtCNUtT1b+jnrxslL
VRKfFB8AAqf91s2rRTKE4vWtt4Ulks9aZjsU3U/VOLNOYcw6Ku9IaX3OBPMQpuvf
/sSbslGChPlNFKLisxWhsZ+Lu2+aA5tMThbWlewvoDnYUYC6VWioroPtJeqecN5K
t0ptmhH3xVpxrZSJMiyeqHwtNk3cmhm8cjsRJj9BSKlrV5qjwd8S2IEhENnKrGtI
me7UIjK3k6yhFaMSM2AbooHN1ArzEa4qPCZsa5wHPyYkJR4gc1tzcrUiccAwikpP
mFqV5f+9qp2uTkmw1M1KJHGQhqc3CZLMlu2hF9HjiGGS26Yb8YvVgN3Q5OKXo+j3
HlPNx7u35x8lkfKaBtSRynZ0UeSTUj74d4aTJfJ0TMmSkp8XFjzSUxbUY3r6XCb3
dTtBWZFQrv3N1nOd1m9mWMwzxP3YPHt9ueXRy1q7sIHYj+ur/1fyrkElxzJync4Y
UbCLkCCIyhk7B0L7hyDQ4/DCy8SRp+pkdmrjC0ULQXQTGp+Uma3zARHEreFh/PoN
C7nBZsfTyq8Kk7Uejpm2//7vXSeXLQLe0G80Oy71v8AeMxV+wLKNkIGnl4ZUMH3Y
ogEvUvi6pGtWr1uw0NEpnWsuWyLbQcUKFjEfms+GlghBRWbeIIr6LBNSK0pCz+9z
VDVrMz7dWo6ghUaqpGPo/ii4qwawpJ3olcT3vY80o93BJE5EaWlLES41ShwNvUcg
4ctZAHAKV/bOFuUSSBSFMT4/rGxJJGd4a8gD1z8HkpqkbmLoflX2TW9KF/Ed/A32
r048hQ4rOgomIAYCUrcIm4n2iOyfEPx1RNBf8GD5dGsoCZOKT5lv3K3zwFhQ+9Qi
/o8Naa4QLv5pZdxNAv+lm2h93uYR/jTvpkNbf4QEeCRN9mu5z3AcnxuGb44aK5gE
M6nmPIZXp+BTTefS509hjvDIreOKB8VJhccZxJFZbTOQgwJrjOuQ8Zul16beOdY4
HKC4k4jEnXqPMQOAeMXH3XX636/BhlTFlBMnfU3Yx6c=
`protect END_PROTECTED
