`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
boSeNAHsehumhHIMZdJvCKrDOqpWDcuZiWm5IA/amddso4quRWwrMwOINmeBtFcG
L9ZM6iFD5PttZB8YISWYrOyjwkiqQYs2Pif9kufK9upEOKQW2HakYpuCxq3rYviq
rMYSTMArLDVZtYhM509A6+Ax8VT/4+87FfK7LJKSd1ArTXPm25EiQPx6qN00z0as
2YikRM8T4wqUr8fu8yZS1vNoYXKAbMGkXzbKGo3dGgLcVKV1rTAa+2CVHQWcZJ3J
iQZ3L5ASC2MZ3qqfPFZtHuVIDlO6sh42fyi0tms7mHzIF4SL5T+O7RYp0b4HuOTR
xCvo+p85nRGmwzk4I0C+MIKmwAbe7FYd+/T4e6kybJ9j5jQLzE206jhVewfvZsls
jABWmZChzBGpqnSzQw6Ym69g+p6tnkIHSjlkypkOO37Vpizj76TxfUJnL/SjZl2Y
shQTAG5OEkhANA7LOG6AAUzhlNaRcxKRCBPxoA0MnUKuMyY4YZzx9UvLymoQZVFl
BzyJpFQfOZnl8zdz0n4XUF59rLNj6NeRJh/0l0XjTyq7xV6Agfa9aAsosF4b6P50
clED6zbRnuM8cIUcHY0oTV/F8BS1LnEoaGTNLj7pJRdm0VqWtUqBWgS1fm03P42d
0QbOBOdWKdLNljWRZG7dNqSalgeWeWuwmH2KX5dPJc5gMlLt64MtMAL0AKyvBtFL
f6o7ZLEBCg0XlnSFLcEyBnCkpu0EZghXeEHaOgJTQZyvaTsLVrfr/YBYIMqS0SN4
REPZkz3BXOt/AIVVmybH8bfynUkv1fS0veDtERsduXUjmSnw/yMQ/JtJKtj8GX+F
Q6uQqUFFZT7KjCaaKNenmZLMGarKNpuD+WBPEX5RS0NBDlMsegkL36fehZ+Ruix4
2ep7cAXtlhCRYKhqtTO/8u1RMaakQpVVE/l4Rhsx2j/2My+6lX2k8EijWodI9qjj
eCmyJDfJj4lSuzItpz+lFm5uxyDf+m8Y4nLtyQnjIb8eE0rUuzxPjJFrOQaWbS/r
ry6vxqelFlNQbVmahayMRwu/P8BjinDAeQhtYJuJkmq14n2TkBE6Am9uQLoonhdL
iNPkEGth1irBw7KOJ4fq1oI1soINbwLjyvx0oR77wt81n21ZHjFmFTVPWjbI3rQ+
C7OpMbNSZT+Lb548yOeR0/6R5DAPZH836Kmy6upMQJAndhwLOI0CLPCLqUUO/39O
/aQK25irb6ZrTpiNsXw5mNdD2kIHhb4ihHnavGKryjQ5Omha+ZUMvckSjj3ZsRJp
XkCiyaZgnZ5TrW7KCCGJUjBQzVso4eE1CpaW0Ja97G59AGZO2skBJGCHHp6UvHaJ
`protect END_PROTECTED
