`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LDHk3ZbMBdUgBh7yxZsu2MsuD6JKFP5ihA6uaJa83lwsk0yP7vvReyrVq6SMx2wK
C6twy8U+G6aozEiK3bzSQYbEzGD3sK833d8NivzXouwtvQ9XSoa71/Vz8waA0h2K
hC5uC3yFErM5uRjI+vyW7oMkagUe0STIc7bzcpzddqX0FmhHNA1WQ0RUVPeAUcCo
HLxK8DJ8aTwSUCwFplbmGw6mg9+r40z8KL/W3dqDILDYnBYegKeHhA0MXpMaK1h3
Eog8mXPxr/BQikotnoWinduDZ8KQaef4KaRTnSckpFFn6imJggQ1nP2sMB7v8rWU
xrBoe/WB6ugX6L4fpPJx7adXnNQ2kNhxr2S0ofRQxhuRJ9wpWqCH7mtTAXkVCQJs
CsfyKxpsePOENU19NYVzJgHnBVPG2k99H9g3FO4MhPjWlys805GToJoD+j1YZva2
MSz10guntcHnxx7+7ygP0XlrSHAWGGRc9xbGpPZfERsUcMVasUPYHG7Sv7fOxlUA
D26k8+BAw9iUEEKe48C1a3z83dUUYC0FKDLSlUvAoaYX4UHnkdz+Glq6zfkcfPLi
VEv2nQAHW4FKeqhBIIla9eVANPiyshyL8GbBddx6450BuKY7l5HZIKyJRsk5HVPO
l2cTxCEUfoM8KQH1By/sRFNsApqKIyqckWfrhLMvpu4FjUHhnBMInX4UdmXejauE
+3vGKhRhgdTdFFOR4JuQIqQg1uxuzIYC8nTuDkaeV2H8EFCsXsLad9CVdv3V6/RV
p+LMvCpU3XFx6kQudVT3CVoB8InuHIL6AphMtKC+3vxuVg0jtqcQsWSRT0NmcB2n
AbAdWoKKPLvnvh/lCxV0SSFlyR+Rd23ayqLa2JMwRJNI1y0Fai8XFwoiYlxElIJz
XXWE1Ca5fqfAX3l5wtIYk2DrS10+b2Q5qoriCaXYf6LhNi60VMNJhCrxVywN8zh4
YEmH+6ZTX4WP2F23EvVUN9XRhmh4D2XC7KzQJsM9yXCSMwP3MHwY10ozqj7XzNuC
EKGy06vIaj+QKbcpgSXFtvPeQtTs3jQ6gOwYUgCDog5MaIrasV8zZIbC1gGZCHDx
MyksCXizgg7q1U5KDyAdsLUJ2VCeUZK/3d3KxhbGlhprX67dGh7Yg6Xtgd3CyWD+
6AQB9w03YQrAm5o+eKD3JihsojdzqPdGs3J1k2XYd3Ij8oORBs5896de081rVNak
VPbeIdyG42QjdS1lVBquECatRUlcHRvL2vuXfPDaOp/J43CqDEQADGtsawaBYNjz
4GTZF5wIJVOu6v+LskCizQdiAv0cHO+AVvWEFQqaKNskjm9A85COA/KIb4cXhHYU
`protect END_PROTECTED
