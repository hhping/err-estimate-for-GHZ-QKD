`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kKpXFfFlrTWdCqGCZyW+hJXJ1FlaA74ne7WGeGR04BRDPLzG8cxwwWFeKTJij0wY
jRXSmarfTxO7mIUxXfE53PY4pEqLYZXzcA6htwqq9ON4vT7CaTS4bGOaD6u5XdSY
WDVhVC+gtNfa/OklhNmkQzwLSNfYpUebqBqncZC7QrAVTktjg5xZEXyLg7TkYAnO
tIwoeLskgU3/PVzGbUgL/5WGwk2EjuVyaQlTmyDsqREasDkRDYWioHfPPdq5obF6
RvaMCZzSFDVUYTPHqM75pngRqOm09ySSJstOQAo5odIiM/4CwpLAQw8pZjRuAw3f
iRtat/eAXuQlhyPZzmrFBppICyL9EYx3r1w/9n68hpOIHde6BF74LIWOaV7OzSNg
BAjbJjQhAeWEJrWd/4mE77gk8xZebrLCC0uEYriEcgeL9DpQ1mzG2dAdRVQxz9WN
nuMB2AV1eOJ1wk0VkeiiBo/dBQdqILRbKpw/LxbPWo4KRNf19B6LuxzTapla0nOd
l3mxGPL6pHQ6YmOYcwJHcqCUtB1w7u9IEHd2X8qycyE/TMR73Pj0bwk2x7fmfsSB
ufrj0i7IlXmWJt4Dk3a1qwC1uueTMfQ9w8cm3s9yS1i2SVRaUqS9I1j0DphS9q+Z
PXfIdD0SG7l62eIddXsaHXrPO7CG2SANVKhFEch2kvYFtdIsbhPTloL7mJpP58/h
DxJ04jDWkPDwzyn8BOAJhrjHEXv8wiuGSpEoctGA+Nu8ZiBeq/Hw82APKU1IzFI+
S4hwe4t+Yrfw6NHjIMHH6CvXNVKtLffaovPeuPld1jJ7gMY42C9OUE6YmJDJzFPe
hQaiboRgmzEBVa55Tyd+Pe8o59LcZDQpAbEIR6CmpGWgEt5RqG9O3m+QSBOUoX2g
cSEXR7rKoGh3ioLe+xy5EVK2k9fK2+c0cM7Ba60v2KapGjZAXQaKeuaMSbvcOLMi
XW/iNR6+hH7mXRnvsaJ6bvHTjk6Gmv2/NCw7zbPkPAlSSy7vzQjLWvekaxtTRwNu
n3l9K/jD8IHPSen0PBVh+cYHZo37/tookvBqlHQbicNEaaPEmRjheRQs38WKcrel
UXwNDAIM58D+jWPYojGwiaOIf8J0BchaoRHdi+ckjQmyw0mdB3Bfz93dMQTRDLJR
dabNbeyAvctaw0mh/UHE14nzcPpYcyWCK5IAN3TfBoJEM2pF+bRWkVtoOMOqlU3S
`protect END_PROTECTED
