`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RlHv30kEmDH0ti6OCn6RKint1yFGOP+fnjqR6n6CHOZMaTUavxGfy1HGQzDgqem/
A4XldaXeW3AUPn0/N/cYtXWBRUDPale4x2Fb2rb4+l2I5swWq8v51EeeNx/WuUIv
wNj8CgsXKIeXNkGeC+W/K5iE8mcXg3DrDGhncOHhsia75gx7fG9i/mUGV8n5j9qK
GgR2Legwm4jvCjUtlrAIV8tANvtFwH5yhSxRB2yYucYJzpkhi67H1z+1K97gxY3V
Y5EO5fEAmO/osiZLBCAGn+G0e0Lf9afiOEb6+PLI3Qs9Lp6fG7SEaGn4nkRR7T3i
2iC7HKfIvD6JSRiY+TZAziXaiHqVRbB8UQOq7FdZdlZNIBAU7c02QXg1nmLIsr1W
VdTCDN1TRRkcTV4ziriCIo30VYl0/eR9nkdI1GUtsVmFZ3aqplZZ2jq3lyFbdFn7
sVxlCe0QTnhmh5nUBOd7Qt71Q2wWYaeot/WRZX/iyMHwt5RbkYiS1uu3tTB+RBzT
acpSNfvkz3oXyuH+1k+urSy41Y8R8oTYRlZcs0TS4/h4VQdDT7E6v86Q2VnPkYQ1
nOamGrM0mqEuwihF3Vs700WddipVuTILMmFruttLPhtWzHXzwzv00eQza/QJce73
maMaKyvj0+Kxbxyg6b6IYjbrw1QO/VLy6jv5v8ZvBYsZUbNETJIiugtM0FsufAf3
LerOXdV95wQn+DUEgFFPjo/GXPpn1YeAmJ8d4gjFk9AtJ6aYKi14ESggp+RmnS8S
rY/KRf75hsZnbuUu19Vwtce5eMsjpKVYwt4ip5YID9htfFMU1+NKUZ8+/WxCIhbo
MR8MerSmf4V62pCNsJ/lmPcl6mdDckA1/Y5H/XYVBRWA1dx4oc0TFoExkv+YIwZW
pIBc9fa5zPTc3yrET8XHDoNFXwHaBgt9lOxrPOj7P4E4LrFBcf77k0LnSMhDBykH
3IusqZDDFSJ/zfORg/8/TbNmII7GUVjbEZur6OSGo6jVqXje7bOTbtMoVuobihgD
OfzU/NcH4gg7SUjiSUeqwILiymtPu8L49IyFKqnjQTXceG9FBAJ7UJe0t8Ke1DOV
9CpaK3aLxQJ0UDboUNhI4A0PiT2T1n7EbwHUxGwJ+f+DyRLR8p7eK90ounJDf+Tr
YtBcVpe/ptSQ5TWMe+RP78IfZoiZ/fdTEfzEg+rIPDVEq4si/kQqiTg3wguGI8jo
4MAjc4BfXWMvSyFuZVvSZmKHoGkLP70/hTkvhPyZtqICRN0BKq0emutqlEEWh5qj
mXVE/2nInoEy2pX/FtiW9LdLZssmymzmuwKtmaQYowY7DnAyVV3Ka7T9eSk1eMvd
`protect END_PROTECTED
