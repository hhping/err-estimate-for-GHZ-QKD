`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RYNBjUEKdyIjANGeQwD10rXk/2xXpR9WdaXHyHUTvTMJRyCjiXTHjqw1IYfWU/La
eg4QnSq2ePYIvHtl2h4D4j2kufEw1al0BIePQhm0Vq3ML+DheQxMVTnOhNVvPPav
2Cmt99C9Jd1+K8H8AtgKnGYPcWCIZYvfgw+ZMC2uwkmpV0rq+BWofu6P6CqSJqgY
xGGp3F3iVIWGoWz43au5/dRrLAoxW/CruZSy/e+gS7Brr9YVSWZ50Md6krxCtgly
6FPfVIvj6vW91OOGhSuzUPTM/Jyj3VveVao/kPMulJZ4i8WYNrQjA6tfcJ4acdOD
aLzllZZz2bGtJtMGgsVweB/dnKBkQjajwhUgVN+MuyEnNEwjCzsQ5LHqxNtGiXIb
nbmBNFdBetXWcig0KynEBoz8Cz3SFSu6vx3T5qOAzzXtXT101d4j3Yxd6JNkfJY5
DVLqFPOF4D8IPO2uiAvVizMxnhJ3tZ/xaJUefHS5jE/1Aqd/hPHRaC3CNbEA+Wj5
h+TLMduASh6e9jT4nL9gWurq+wNEEt/AuzVY+Rhh/YViJmH9yWsyieeKLUfU/DUl
7/McIYE6kLHS0EuG+Zfxy8ZmlIfLaISxFHXramr9WZuipjaWeRXIF+nx7K9yFqyC
7mpjMhCRLI8IfRZra1K6AIHIrS0Z7Pm29hX3hL0FCtF23LeqwAnmqyLb+CXsF7jD
Tk1hJJLazrMXd3DhCQuBQwlH1C/KNUfcm0U9yN0SUxEnftIt3e6vXFO9iCgUQmfL
Z62nCnQgvfi3GsmlQgQXQIDtuX8yMAK0Kox3x/3/0yHhZXf85Xt9arJ0vxa/ZgHl
Cz1Bz6FVO8VxSyA4gWis6et46/oVIJG0qMIb4T+hl2nbYiprqnByQNa9i+DYaYnR
74qA4XgDOraWQIwyvxTQjZlm15wLBFOfoPU/ukxvv2LS5vqouzqusHRa3AqlYIaR
pSu0Yuzrw7eX8DCarCuFA65qBdATIjvHSxFIvaShnLvj3RE0YIlWKiF6AXDJxjix
2dMTmjpqNF0zUej4Luv82Sc8Ak8SXi8CiQFS7R054eSNKJ4uiLB2gCvP/bHcbLd3
gXifSXMKWuQR+5R/rMpgXPmS9GjXBe4eJhuKUWFmXvvoTReoq/fQWGSqf+rjqjw1
f3cv3e1XuNMnj3SLKITxWXhjMG0vNkH+/hK7xN+cJpvGGf9CP0bXCrHrdhJB4dEJ
xdb7EdkE7itJCcm4tltzGbWAp6r05VKdDASH9i/htYVvQ4EmsTwm0N1WYLUaCw/l
D6k5h8M0EcBI4nT5LjTjUqvXWCvX1GO9aCNevhM/zbj17KOjZRYpKebjGZOOfXwU
qUYVtupA487e9jNLEe74KtqZe68E08j6GdHZMoFDAiP1LIKVn7ElZw8XQ8/Xb4d8
aF8pPQEDmVU0EpUStel8BlOAJj53SWwyHlubYyVP8IlPDSZHAbJYMzZZcj8KbnVk
Z4mh375MVA0uCVf59z9XDWQdFSZ75m2gKeor+/pfpwWxyuI6GxQcjua1YzigPYce
Imj+7buaumVr5ueumFOWFWC0RInMN+1Sj6XX6hQxNXpAW1sfJzrerFexJIbfYyyU
fHAmUwS4/f2p3etgWXk9Vqayt3Q9bVS0nyOdjmGiGZbo7IB+zhwCcqMYnRJWonWl
PC0fwMpIq5uh+tDqHvZ8D3iRfVTqSEAph4ITIk+kuTyHCuxAgL0xGoHiswWUeMIH
74yhTGzVTc20kUqvqHptXANZiWf570f1Xlcg8YxGGluffQ32J39Tcg0mPnSW10at
k4RrZO9sL9FExmIhQAqDLKqhHwq5yy0IyPktu5xrz7yFRtq5lPhg8y+AY50l66Ou
wV2NAuAwi/ilqL+QqTOGAxrr271AMKPFMrwyFuZxqaZ0Taxibg/Rl9esnA5fdeMw
dv1aKNAz55EwLkhg6VaU/QMvv4+dpCNdVETgneztiPWTZpw09/7I01gtbLVPZEqz
ChqIVGXO6hRG+do+pWhKss/ktHqLKmDpQlX7HqVyhKux3QrprCNiBjo1wAERDTtq
adV9iZou7cMADbZVdZZsedXwFqJNpoLRrPnCRNu4iEqsTJv4NCc+dyUq2UtA1J6i
tHm2KISh+hDsMh7YLbMQMAOVx8qAee3SPjoN2c02lQGd7XKsCCyO/Mh06yOBGE/G
UbH3VFoJAnQ7IaYDmhwZgkl62DCgp6SJ8EQlhJYdWnZA1sH6oUG11h7Q97EDsdUt
dmAlvSb18oyptPUVI9/WVGEXeQ2bXc2w8FlpupJxScNCf7IFsOnGmG/mk3SWeill
Bc8G+U4l/x1sshpYeNnzEADz8Iqs+mU9Vj/U1Co+frfpnlwF7cCKMBYuH+lnv+Lb
NJwXJToHCS8zjRVXoII/zL6zfqDhvG2sJdzSqAedf/AZz9bXAv55YM5beJ1WL8xs
Hs5qoEg0tNtWW2DWeBU1dMsEqjgRnn67xPU/i6ngf6dgX4Zl+bfqWK9jN+bSynh5
C7CLcd//3PHGwjsAlbCl70nUHqc7LhbFAVr07EP3ulzx9BeuhZHhsD6kCdSqw4t+
YO9dr2QV3xK5I6IqfTdQmGnui/ktZ4pakEQCDNMUxpOhzNBRqr1LHyVVsF/hEwFj
88dvrEpPaaKrCckB2y17p2DWLQ3dyT+tdLUYiIR3HgmYZH1BukQjAhcdDUTNH0aQ
miJoJDYTAgzLiXbsnkAFaQk1aJxQPXtG1Eev6cCFXQUziak8rSL6OWNMw2fHE5s2
v78i4JZvrDn8PVNrcN/tBc8x8G+ipN1VmjVe70D8+s0pT3eAWi0P2qj7X9I6vmKq
3CLZ+6TV66udMC9zbxHXxzMUxj7egFZ3yY1qEYdKEpXswvMqotmsWmozDFwx/JLp
yJ9RRKdMDnsrEJc4ffFya4JXsMXp9BZMoesoNz695Cn5qSq8FOQOaO82E3phZPYV
6vm2rh9XmmC/+iAcrrSPdvHeUmfwW3f1B82tWwRgw63f8Jl+qylQi6zRrX/KHmPG
UdTgaxv4CITDlsO7Qh0dtP+n/AmaEZkvt61VSS/BzZmzO31XQoru6/jn6jzWz7uN
6cyLzvynCcv/n+uciYkfJPe9ZgxmvP0SKhVNZSr8fLoSBnVsM+w0ZlrqHN8QVHsi
iijcfBGZ/cFmHIYFdoNe+pfx9A7NGyl3lcjJQlmwqtyjbZunF8KgIC5pQ/LOM32h
UoltKeLakJhyJjPic9KMaO/7KCnEv3PhfNNCRuUBE188Z/7mdKxb1bxx/WzsKwiO
flFLNvCkJHpFbLWuNc4hM6hoWN0ztKQOGymB5PBbGgE9iG7n8X7iSp/m2JCUfJ8f
SUFSmwf8PfJ093J//AiHQlngbcppj/Vgllqk8nj2AVLz5Sii9mWy3uz1G4DvX9EL
IxfidxhxG1ahxvndzT5Q1TIVtAnsBDiWZiONv5QBVPRbOKoCRV0p5fPnFeR+Zf04
4wA9nSWbCzpVAhWyx54eX6LjmjtdRyz8VbSo4tr2tNgsLeBRIldk6Tnn4Q0ZtAXQ
5vog1x827Zg6HausnU7HgVA1X5gQxzeNVNhjWlZYvmVFN5RvvmJgUKUP97kd79Y+
Gl8akgDGEaaqm0EuASQFgXlIu4KOdEl34yWueKQjaJm8hqW2M0eW7+u0fAwp7CXK
ieft8GAD7I2bGjeAda4AZk14gWG2QZFd6ZTm/IDgdcOicyFJFdxnCLhm01/Xu3RC
BRN58s8WGwDY/M41vCjeECUgl7Wdte4vyWwD+hBwYIg54LFH4D2rjQ08b5+kLl19
IVtBR3WJ4SygmYjiJHlIS+4gmsABcm08WE7UU9WttuOjZRGVfrTsiQlvcycmJKgJ
NuL2kk76PsJax+VwshNn/OlID/Y4KK4DA6eR5eErX3wExwQBjtAPYdJOVjdIcFIG
v5OaW4YtG6xjjfhRL/WMfd0/Holh7lX0gV3jDCCJ54gYTqBitaOFlgGLbKiaQ6mf
3dIOalSOJIVWIZvCqpEN44SE3R6ijkspgSKIMPiGj1NGrLe93vKmT+QnrCV1l1aM
4wIOYRJyDc1qc8sN55J5iYepxhVPYHLbAaxf0/24qIBMwwIj58bHZGYXIYmLTKaA
TSoFipqQSKjPycZXGYePS3CgxTyopW+ivM4Zitac3KdhPaqX7bUSJegz9QzLQoIa
G5j7qAd8oif1fQ51inCGJv+wm4jXkzYY0p9T6z11wksmEQjVStEOn0jNkaIrr4hm
DJbzu+PBOOzBoEYeHBhsWZ5tpGpx1xa18uCJ+jDUwet9rlhxwmkG5FGTRqx4yy6j
Nq2r5HWvL3rTEgKmMnlUWEbGTtLfrxDpHBfP22jYd7xwKzUsOChPnDpEPTL2Jl1R
WHZs1ItI7DLCFopnVOnawdy5L27S8PWf2Ek99o4/U7kKNTyvjf09VjrPC2Xk+0hb
f19XlKcQxn+GBY48TQzw8XQbxonABscZKosIAygcIYedooawNhrXCciBEri3eh0O
MIEyTop+34UteKTP11mzNj3lfCcYYkflBssrCr7/sBZi0JS3zqfro/90KGt+DeoI
5vFDMcFtuttlVqQoi05nDmcZin+tM12dOHXw+bo5utSURvH3NLDujVu4/33IJJF5
ZTwdNiHzhImBBkxZg+DuI2DTHhPDFq8gjCWyhkrjKxufqlrhC+zfrtiJwYN4FoVX
6DAe7qmUesMBsJ4qfls8NxM+YVVIqWKuTm2BdLJflrB9WOU+gbLMHgO2BM7w/Dj9
hmTuJ+PuX5LZ7aKutjm1tSGU7jp7nl4XRyr4sArYmh91D+7MsOczbASCXELWkn6E
U3yavKH18iDBNRLK5GteidkyVYy3SLBq0v1uIenY2uBF9siFXwgN3aHiFcZ22U2F
oAEt5/4FRsFQwPkDzKqnzWxy0b377aRN1dyxzenjIN2SG/wFubRIXhWBf6uNCl1U
BQuTIqpwt35YUNgB9INo9wtGzTQO7le3OYwKxNmW9+aW+c9YAIugH9sJ+/5aEZiB
9M7TQh9+1U2zMKAdQjxKUhkcN3GNDbTJx5e87KzOrVZlc6zmOjUN/8Unttd2Bw1A
FlaZbzixkryOByaLcol6K13RVcgON5JLBcZH/XP0TjqOraCqnPQTbI6Ng/6tvBBO
QXx+fwrTHxjfSCrT0NrI7tY9/aEf5qQLAi0WdAzoXw5e2Nqp5s4E8VYdsflyDvnY
LmL6CGOKKAG71Nc0JjD1ijbkygbyxkmdNzwXXIdmL+z2a3As9tNFZMTqD6yfPFck
xr3rAcfN0r0XfIIvroNaaroIGEGVze26l160Oab4tTEO1ExNYYknMTM1wNwxAIl7
ef7rM9+FZ9y6aVgT06477MmeY10wi587Bn6GneXbWpcobRGst2qvi0nlKGIGq+Pn
sE/Qe2XuD/5ImzhF1loMxhU+kf1Uy2hWNCogjWOqzMuAGCjaTAqsWXITaOYv78Q/
AXjCcSJAubkRzug2bYtbA3+wz438qOfK2l7fI2RaPBIUFTOQpPzCMRu9FJ8CjL5b
xALvL+2XmyGIc08SDlNeVTVnrXoOfQkDr9THQdna3RUzqFLIG4iBMbqOoe8l2OBg
PBtnwbXygM9/yK+p6RXikea74HTjCwkkwfkzxq4eVtbUMFJLVmzdG3ZegpGHrerF
PHzp/NU6R7NdmvELaZC9Ya3HRMTfWmq7YyFeorx3CZrIA0AysXldAfa2eSRsYkDl
Ea2ykiG5N5i2j1D/6bL3Tcq1tIcuQCUKPM+AAjHR/+0+goB8xfevoxIjeoF/MTM3
zvU1wC+Q/jtkqevdFxC2HsTlAB/B1R/ImYtyWfG7tfrPflysIvFFWUlcEqlTeP2r
38j9t/qmqfee12ayoZjKDsuCTVoxpwovZhbZpaxU+4NlCxN2jdNpjr01DuizXte6
JLUrPzKBXHScAy/RrgFz16pOVXK/+DE0iTQsX9t86XXWYHfq+RoN3prY5ql/hVMb
axlH8TM8Idygvlba4qEaoXeFgGo8gX1uqbRnaxznZOdzZdm5Kd9QcwqX34DlvctV
ejBqtPC949yBwYVB4Qv2BHtRQmpXCnBZKcIR7uI1IDfsXFKlmsshZdRg7t+VRGOn
N9c3xkhY9QfOm362il98Mt+nGuxiP/p97DyWkz8EMdLLqTupnVMaMf5Y2A2fx9cJ
OcL+eYcEWop0u1nFiCharT4Zw2Y9AFDwrwN1dztk4H6+4EvwnkYW+UULoAbFvtun
fiw7kcbrYh5k0AigZNUns5mfX5Wt6WpyiMaojc8zzT7Njj4xH4pf8M6Hd4FDH1RZ
JR+lnrd0rBHvrp5a8DilWCMgy8AhTHHmA3yeFJMEbV7/MKo/FUX8QLmxnwfBaLzv
UHoWLcg0W8NQyiUqOedCH1v3tuETvpmI0NJGOIhWX5pB1PvqWZ6WkwOa3OdELC/w
pgYW3wRzvmFgzxLuEUJuJ1IpzwNmi18JY+PQpzHmmvSvLg4z78J/KAtWZ+ATRns4
5i4GsR8TAUnCw1itisoehaEkhFuDDNSG4yc4EW1CiDfqEWepGLw7dZTAPFAJkPjV
wlBcc559ixoqI7nbWVelhsCNvm0dh86DOdUtd7r5U0kOtfh0FdfOLGTf00ljJEfX
SBbngkTl8R4c6TP+5vG26LX1MoIo1bw7WisxwlaFeWplEd6E5BzyQlUKXkQc772V
PyvpCP3IUhWWHoju/g/ZNl2peLo8TXI2pfvKE+yxOUUkWpLXkhmsezJbzoxdsE6k
93oXbU3hYA5C/r8DFRXtFXEMSWr1RjolSs+zqJB+25r9lvFK7QX+KKjwZNDwrwIy
sAvQCutEBEkAXnc6ClxkjOZCyOid1gQBylejpetMil5uWSpx5aimY1NmqcAKTmke
PSaUmz1ovCKIwF8gUQzh1vFOPgqVxA1MmDyKKqwCa0QgV9n90etIbnCHgLUIvNAy
rBhe3DWmaeRK9EQHnsjK7VzpUXEjnmB7mXigvObNVzsabe4HJoGyK7sfz/PiJgv9
xSXDnO8KFxjYQ2WBLslSZhO8cJ+9/n64v2IKDRUNq2n9DABDPHHpSPHTUviVfbNL
1B4jyOv3M7NZcQJhOp1Vuunv94Gw4oEmk8QMPb2g+q7koj4bENbwU5FhPFvOYqRY
LZMX8mruWnm18QWQW1cucrZ6CHSk3rhoSjqhVs+krS3WPf5i9PzfzRTE8WHntQF4
h3p92uGz0Wzm6lQ3KxqST8UQdUYRFLgQ2Kloqjab6yij/s7nitJ3ssNr8kYTlwf1
lmzJFakFYuAylk6qoFSmbX78zxx2Js0lgesSpmJSoJzXO54/MiKG4dOTMhDkbJwt
k3i0p5S6OkJz4dSDw9KccD6QSflTjxAdBhqOf3nPm8VEIcZQ6tcAtHXoVlIevgpZ
PmfVYEL+SgrhF8fNniRgrKmXQU8fBZSM4a2APTeXMjeelUd3HHQB7VvW5AZrB80M
IBLyRZ8ALO0zHdkvlig0M/z0XGg8cySFhq+ECuH6rZOog4er0pIvJxor44KaItB9
bP3cjCSDv9UaYzJ3qpuW2AvcNfU51zmXmvsyjPnYEIj6KaxnPGnvpsv2Gb3AZWZo
d7BjkVzNU7en4jxm3gpFv39KCQz/wl3visbLzb2myezSCtArVsCyuMJ6ILOUORD2
qWQkqosu4CYHoha+GBne7ZFDcdoiPc2y13OZzleqMqeobWHGK6RMJLe4rprNK+AS
xnEmqKTVviYOoi//skAN7dHUFT+xGnQIP2wJC/to6UKvmJYY476XWkygev9N4q2x
aWjvpmZKUgwMp9piwDUT9s0CigKtaS+J55QNpMrO3vhk3CLxhla+7TOhvK1Iosrk
3wSlE4I/x9gOwaaCXKhPjRF+LOFBV+HjNBpbOxb+T5lRbu30ilR2QSmxf7Jw+cVa
m/yG3MdNjbSG9y1+MOGwe8C5Ad90ivFz2PQuiaV4ZWorTIQtvgwCxkRrIIOqxKqf
W9DHD00QTa8xywRVs9Dh+ovCeGx8B2vfdkmoXxmk3Gp1zgOmv6ksT7E1CXzgkx4V
`protect END_PROTECTED
