`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jqge58RwJs0AtIzXHwDFMDyNFVu+WhD2oM2CpYjWN0XQ4HPB7f+IPR3lk0NdOdBv
/kODQom7Xgt/HSXie/VTdXKg+ZrwbifaneAnNOY7CuSSVJx0x2sJ4Szy7io8dEGU
JDufG2ZPcjMZNO6NNpqVa2odoexa6hV2MYSGjhjCcMJXCRORB+uiJnmHGS7wCfKM
nVHS7qtKnQHQYjH09KMZ/AFXLS/NqBnag46IeqTAIEAdvusMPjobDRzuszgUYKKk
sBaKFWM9zUpqeFekdS+YDMBRdin42cnYJlfK3/f0nOULp/I29liKZDucq4l4+o2T
54hxMk+Qzo+jW7QKL+u1a+vI8wqCIR7uYqycZDlHU4chDzCg7b7ynFt4fnp9hqb2
mavqCbmSYJJXZO0PDYx5RE5ZQI2ioYnABcZAlkmSwgj8K1I11l6T+yiE1q4PZv7j
LH0QJue0WsZaLCfPCY9Hw1AcUOGCjs92dVrHhrTrh9E80RFgRt506VraL0SiYAte
4gHdlAnAOU45CTAv0n41ruzdmQJfUPSHRLKMyxEaMSkODbdsbAFFOQcrPLG1+uQc
2+G6e9zJ58v7HZ0IN5UAElCgFt/LUAmJ6c4b9ixqNAjMS5hEySFqjP7FmBaQ680b
5bstVJrddzNpU/odRQ0wZL5jfddMMKqHPuQgZG+c0qmAlW5dYM1oWbyZZox9ErfY
gryOwbt2zdYv1e+ig9BgWQItdzLYEyzEXOqaftzlkepejcHmXCnmEVvITvUG4urr
qcMTLxBMsMwwsCtTa2q8Xer0P5sE5IaOC7HIjMKpO+GDO/HW86F0zw16NyaTtBdj
758ylfroaCpIIr3mqwl2zoifgWzMq89BHfCmQX/KwgvfaCDzlO/A/yH8QfvbpJWz
OnsJn23fAzVF3trV+5qzagqxtP9adQKhVb5cGVtzzjY=
`protect END_PROTECTED
