`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N1MGZmdl17ynbwP1FGWj7LgJwbXjIaw454vukFT6RpfMQgZU5SUDWCRMMlRBGuxV
65BPZIfk5m67Tvuaf8g6UtF7lhdyndZRECfY/I4rkasSZiEGkj5tEKCl9mnbhIkV
nGa44CA/eBNcEbNlEEfbusMnFZqvX9H75BLQ/+49T6cMhxVIZBNWTkEQPiw4KVsg
y5sb9OTIQoukNHRcOBoHBgfL4zlI+QCQLULPM+NbQFJV7D9/Vzjp4xtz3kdVHfat
mXoDJepVsa4Vp4gmayAabzZ078AT2T+JSeRA0sDepsy9uqxXDWLPDbtQXsorKAk1
IDEJAcu5O4po/u7P9sgGHNgJREM+CiZBSxVa9dWJnwqxXdmkhvLkFo3+BpkpEHyu
r3EQxb/7ljk06x5bPPCC2MAOhwYCa8TbF6eILWw9hYq0FDGG4hiwopMsMxZddQBx
vPdeouA2b5En59YHCdVPtjXboHBv80OhGOXnZwxh2p0ZnR0PeyRomJiWb9QOWdh6
1yKm+W7qnpPjZ6ueh7tNM4Z/8AmbGkeaOI9FsfKPgYJuSwTz7D3T46VsnfhkJ+1y
pcHgLzlh7lcNlgYmF8ezqVgNRrz+W0Sh+ia/Ho30OnL70HD6Nr4y7hemkSgfiVrG
2o204vsgNkRPVjMPuppJl9HAhxesfj/ESecgpH27n0XXCn/GxwgOSO/EJ+TesO4G
DmERg1oOPVnyDEADaI7YamSrIZ6QZuACzufBpNmKBBrQQ44+Hm3+ZZABgzlo/Aei
N27SnUScTgCx0q83qsRSpfrmnJDWfPfuTrsNKnIIKzuzeOZqifwbdYflLkhknSMY
wycD86SHEHNjujxDRK0U8pBnUYBydbT3Shfiynlhg4lUdT5zIz0Mf9zvq8w6KQp/
11f4QxnQ+W5lLMGOGgveqO3lzMzD3sq7ASV/sIVwGw2UQ+ez0Lzi6j0Ht927ST1W
zf5xHr1+IyMOoDe7PwwrnohbZSsobJ+K37P7V1Md5eiLqiDWCH4U6iFks5Py3ye6
MQscnPTRW/tpbx9xAd4d2ny3fYI/og0uIJT2P2CCYBxtvvOCtBs32KOuZvKhcVEJ
QaecDTszhN2iyE6KBoVQ3jbLkqASF1waEEFLkivl+oDGPY7WtkCHvUKFz31CbpWK
T9XZS1c4MLU6L1o5Nw2nWmfxoQxCKAHn+IF6QXaQqHvQ08widedyLzOw148e/4K5
BLn52NX3uCAZsBFGuAsvqCAPmqzae/AoWyIbW+eMYQ0EP/v3yViYrXM6nueiJ2XZ
bUCWL7is1LVKOhMDh/7GkutRJEcVCxdmVzV+rei2R60wYU7LOpQLadoTVMXtXSYc
3OQfQZDPA2UDqgjsedJCNvEoVc4IplZe0o98vMtItq5GBQW3GgujJUarAW25+KPT
WILFqZEDmRGU29CxBCsRet0PcWHM/Zn4riTQQGbbQRHRdqKiSMTmNhkUKdF2Z8mO
KeuvBv6vshHK0a5VSenFA3NyAlcSkNG4kPJcipXqZwHW9GSN9wctW+5if8YmRlhq
R7micd5vPuidaD0Gd+ytM13QBEH70D54klto8jr1GmLBjS8bOCrhrc2vYhnVv755
EZQm7FruiXrz57W7w1C71qitJOwjwDI8ujSLZBahhsqYCeBGh0ZdpQTJpF1SBttO
egfb/o/zzvyGXAogNvzHZOT6XnkZWZE7tyPUkzpMhLi+McQxexdqEnTcHM1JSaJp
S4sYsZlrOsU6z6Yh1FoxuAK4XkXA1THmWTr9mR4ZOWEMm6vHwmriFoJZE+aMnscB
wchsRIeJrYalDJ6JPkdr0p2YlCdLTlE2B5py8WX3MG4WP9Wa9qfIBd5+bybI/zdn
rRTbV/0MqF0FzPx/r/j+t2alJgHn4Q8w/LvKMAUZqT0a7S4sda8um36cdVBxciix
z4szl16E2RWSG1We0PAfQ1ihyI0MvRggIcFZGnGx+yTFiEpJDkgot0FAJ0FXjq1i
o0/vUmZ15DKbkuzOVXyLyk8F99Wa5WTTPalFjjQOhCif9RiUTS4kp14lCe4WNjIM
BBSXjyMmHuhkr/3qajuRmH3oKI+rF/Ewvb3eJuY3j/t+UiVeBR482TEhdTXKoXOH
WTfHDG75QXMx9XYnUfU0qcP0dwamIzLExme4C6GDNScNmRMkx6rrXbI1RupiHQFc
E+h/puxK9GXXp5sTKXu7DPkmGa/mVUCjsHPxLQ5HnA9xcboG3eZpUzljcmamnF6O
xMIQPPo2+7amMJylXoJLx1F+F/sKPeX802YvD7TasAbPlyYBQXUFFXCbVkXC01O2
5FkhsQR4FwHtY3KCGhagWzi92yZDqc+iRwNYAEdu3C4G8IHW7wipy2Y+wfpsKXio
7eCafDs98CQmRip3d70C232MdQ+A0Qc8y/aAj8nn6IUBXXOYi8LZxbtxp/fV6NeD
YPgfhJO0JDFr4yYHO9o10YIVhLjQu9WHb+yP5bdIQw0ku7x7Q2TnSt9lh0zweUOD
ihxm4oODOVZfCzZHEkYu6UCI7hqmqZ/cLiqQg7vqZDwYRZ3CvfqpFktTowy9b9/0
9bcQHGnOetXUFXHgwpvWZ7LXHt3fNErogwQ3AakNZ1ug/f55GJ9r28mR8L/yBraK
+1XAEzth95dHfvIQUui029srSETS6uRDOsX4+OHjXKcOp0m6ehdZfa8Sn12PHFF1
Q4oyaJNkysfEUJl5cCLgkm6LaK5Em4tpU96mrGWZskLnYk19XTUs6rxXYaVhfKnc
PFnvX33/cXpXZu6DkzNdkYTsOIEIbb/BpO6+e27x6oc2+jv/OGMEoD2q9M5n2ihY
T4P0+9+Dn2M/B94o92mPS/cHUoddmtH84etofkyfgDg=
`protect END_PROTECTED
