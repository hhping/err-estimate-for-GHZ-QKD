`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9PDfYAVn3zx46xSlR2S/rSza9zESlBtqtTVS9ctgKqVny39jRACseMK/iZSiXKnt
l9E8+xIzshiLDiwVppfsABka6lMOKrWHZC7mfElMSiihh5Ttn1CNbl8xDUaOzdmk
+clWaR1gy4ufvI9q3a3NVRlk41xBqyXlD6CniqOFylzCyYJ0Zltx4+O3f7L0n32f
`protect END_PROTECTED
