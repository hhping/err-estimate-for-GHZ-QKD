`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r+6x2gYx1uF/Ln8W8qyY0srhhObWBEwMB8zc/HV5A9v2tcuzSCW/BhXR/q9KrC2L
YVarWWrXYeUk7VaUZry64/3q6DvqhIxiQMPHaE5Clvf5+uqSV0InzLJ+ZOx7phLW
mqXA5ddkIG9N275blkdKmbQXzQS4z5dsLjJFfN1jEO/rtdHLlxQmBgUAndSYUeCw
Q981hwsqnf0P0Qw7qBn3M3SUipikWgulxqNXMSWBwNuCBlLGT8zfLdmhj7TPKt0f
D9EgerjxSP5oubnFcRu83jU19tyRo2HEl97WTlBSB/fvXYKpI0XoWwEXt2Z2JIqP
fPo/BGEK/rOtpuPmct2ACP1Qxm1G9AacMjRW9ylbA9PF0HpzzH6hL0a+vVZ9WS7M
zNDFppFB6J3aGxz0d5GSDopN0+zYXB9QvEkdfTukMfu6NCEmIW4IaUummYCDxkV9
oVl7UXFrNUfYFiy6XHN5hD8enkzIqDrRD4tBj3mtFHnE0IDIG3Gtd0tcQY4bmkbT
BJ1axgnPCNXAv8cOXRjOK2Z1pHeMSUihBoogRtWG3vHCmyn61sse63YiZcSWDAMP
EIdgHHlpkSsVnOFCXGn9B6RhfuLucKEZBjHpVAjgEscM7Cwj2qIZW7MdM/8yIfZ2
qV17EfzOlr/304mShCtb5PAFD6mNGuKJuaLtjsZMbsD/eroYtErBv32TrfCw1eOy
fuVx/FCudP1ZHBqwP5csKFT2w/aqMaWIM1hXtilyLPcvQemVtUvYYgdjMsuz5qUF
+lgih+BuQGyw7rBjUBSUIKxlpH2tou78vyTbzrllHzUnxyv58VMhm/PPdobFLJuK
KU2zXZdUzDDLAw4XlCrdpuXCRGCC9LR+UksbmV1arNiaJkEhc4oUf5kTZwHDffOk
i4W8BZVwa6Nt8XXDViR5rVulBis/B+GIs+14dQr2mhyWWSLQWlhfU9kPtqN98DbU
6+AuE2+pY46IMWiDhFAAGNReXbXcdtcFSboQ1fhji/1ane/wAjwxVNIk5eVZge0h
Obh95ZeSEr1LwWPMo5E322fzCkmRH+P95b4W4JmnoGajAq0RlE2f2baKi59bNt4a
6ApkGr1Xn+lFL002GpKpcc1GvY0mXcoY6/SpUCjAZKmATxiCbb0JJSvQnnb9YWHI
uown4ejz/p3eqaNuld3PFWGgTBe/w9aq5nus73G8qlc=
`protect END_PROTECTED
