`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R+5nQU3GJ6JBNczGqNH54Lv6u+5q4tITbkytQYeUq2eRzuLL0b8lK/c3opk4/MTp
INLsWfDfSVLvjWjOdMgxYmlW7UuGhI9/OM4g/qr2eu2GNNiUr9Fm9/IMYqVtxtQf
KXlZotFXKKSUGtF3F+rAk0dTCFLuPNvcLu+lVbjjnsI/C/QAYVrq6+WBuLZKtXxB
SPZyfDjvPAQje3dAwiUAVJNPaA3jeri3lA4pBA1TH14AXzS6gz5Pg5nDkHCoAIdX
7JROod9Vx4CdUVx7rOLoOXgjN/EnQ8TAtFUezabjEwZcBJ+VV5Hp06koK3Es7zlQ
mEdCU7DUmn8iWIJqyZVap1Jg9Qyy708OlzgbucgJ7bKTzsPbCNcxzQCn9StFtT6x
AdLLrIdhqFJU0ohj5y3moDdSkrZQoL+EI3Ez+Wsnn5x2oaW/8lem+KKFhOVH7ROS
`protect END_PROTECTED
