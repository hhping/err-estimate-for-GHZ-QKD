`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yxykR/TVTjnIc4chMR8bXv1ml8RwZOiBu9DLcDV4TfWDayjvFsPUQKvsD9US1CFp
t1BiNkDKp0QTry9Dce4tmFuQqG4psSjs1KX1wmFEK54wxu9o/4NqQHBS9buQIuQm
njFaXQwpjgTWKuxUIhPZJS8lFYk/x4wO2yAg6zxrsviFaGb9ieQukjODMKX2VLpt
yC0uiyp+FvdCN09SbAZKCyiNaSi29DYUz48hu9fk0wBWiFGkCVfj9Ft0hLhFGrXV
gX6g6J1KszVy3eIhv7JA7l7ewHwQReJ2vBTROQWnacFuiMqd6kMoxE6MhIcl+sAO
X5kx1HqVDbRXmS1zpS05vwZ5dKTaYHs5kMlb1zn9VtYncYF5GG7zJcwt1iEhjxe1
/+FqP7Zh2fohWOy94hDT6AcZPssfdTUE3CRJOoujQ9H+GmegAOLUsZNxHb+MSK7f
CQ5geMtWJ+SCKfPx5U/TQvtF3K4dgJsbF4Dxun8o0ctQ+5TLlvvteKLQY5fu+vAA
04Yxk1oR4bc2TY9AIkPOrwXJZfDln0TZdCgp4i83MwK36gTc7EpowxzsOeTiyj+g
+ymeAZsqE+i1cPK8Ax+u4KS6DT7Try4uBOSTvTKKaDe525BrV2x4DK1p02g00XYA
7C9WOQg2CHrI2PMcXpVj4BxkWYmqRbpzm3BnLwPppV4AKHlXJG2wL/H9ZzcmL8Pp
OFeu4uI3gmbnhLBhDUjOrBLf9j72VuGb94YOsuky45flG6/w9K/vMB7C5L+03jy6
NlhkYkmfRxHqC+pp+J+4dlQxgbMX/B8IITaGQGMR6aQ4jdV9JjtQ8kg+Kl6AHvEe
M3ma3iQviIbH+lF2o7s3MouXlW/bVnVsRF9xhMcliR+R3GuXD20tUE05hyDWJl4W
UKiWdHXkAOwpTYwm/1m0ga4LPvDnl1nVmh+mfvwA0Hl4sJjTsO7RhUhhYwtkamPD
mGCQncSOLSNZA1g5MlY5FVRj067ctI9kwIIAfqdxWa1FY29HIXHqAJPWjCDbtlHa
9m8bVR7jp6DzG3KZj1PGLAX+705wSg8yvI4pijxkZSuwO/fOWUc2zRNmH8vTYJ2u
DmaRB4JgRIDKpfvjDT+GLdRK/omShvNjh6UZEscY24/n+zu56MEc8srTWFHKOUF8
q10oM8t5fFwxjmGMixtOfUIEcpd/Jhqlmzxwz+Cl0TdAdW9eTZsdtjXLkqz3FSoA
W1TJH/dibBj1/Zie9gUKlpJ1XhUWb5rq2Vm73Xikq+rIUWkfvgW3rfNJp2NUH0UZ
SaSAyE7el58TRdoy52VlEHBd25IgDWes/2xYcxofqoLMJofCkOyi9OqE6Gmsrgwx
zmuCE3LqNs9TeY2hNWaX2KEDDEzT+q8160NgD9Vql9w=
`protect END_PROTECTED
