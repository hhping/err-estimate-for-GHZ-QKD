`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5ZMd5t2YibWu33t9jmU0BmZEExLeGA80rdQzfpcMhthnDJnCzv6kgzzzQ1LrZIBE
uTgOgZOa+gBhLTkASD8yAHxwtCANtyJEW2yZX739Exk+488U+wpLTzKYrOM9QzUq
T/hPpPe5Ds3nru4FZJUD4l+6uApq0gew1LK1XDL+BUEE5835mGJFVdaG4k1vPWT4
ipKsfA2KTtOv7dfEnuy4odJmV3RzHbmygDNkYbL9zQ/fe7ZWGHK1DfmMAXlx66Bu
8FJsxkxT2If1jXatta6o8L16wR+w3T9eeJGYmxIIeqb5VXzdQoleJJf+cGpog/Xk
ZaoGK8rvTPOSePMEayeDDADOg5amGQuiz+8DtVKtU7/mLKZ9Qg4+Lz3KPa1vHnjy
BkkNCSby/v8hAdG+MDhfwI50nvmlPLLgQf9ter+Tud3NQ5FpqWvQphajGpq42R1C
4488L8PS6dz7GkSgxltNjbr2/ULOHt2cPppM1B76jTWuNJkItxSi0FWq5gdZJtDe
DzztnprmWcAo2eacZVXPVQ+kPTcgkVb9nLkwjSDcVihbIh1exbvDm+CWPuM5gkBp
/jDvHxd2jAT9qRRRC8djFl3hWhLM2tY7uBRCBa4jRrDAvLtKxL2vTucxPErSf43E
gYkLgUbBo5sJjN71tGHUHVRmlhXc5BM1nnlFTyp0lR+ZyTmN+qae3GbaNjwB36rj
khyc+s2wL7wc3I9NSMQrPFkteunjuyTNdSrojD64L+YDsDXGSq5tQy0crC6+ZdOa
zrXFlTapJAue/BaZDyGZByDsGg/p1HejbszD9m4HhARjbwYbPsguwB07RJrScgMo
ahCQgPP9pUcfJydnVQG6Bq1BRqdOvCm9dQvHZF4+FN4jNprrwTLtDpLocbz1FO/C
Fy62E1lhMtUEDVfVCAdptTNTBPR9UKcEjBbDqQEmxJyodj6Gb+F3nlIzP/HUBzp1
+Dj3aXH2+6GwQumMcviQzuZwqXuEld28/mr391BeAj8P9M66TXF1aGcFVfwUmut2
g+5TJA1pfIThdh07bMRMpd0Cp+mvgzlOfSdpcegUFyKPRO2KW8Uk8PzFYBcz6K5V
w52zkP6LwBC1B2S4CEmeidPjZ+ZgutPwZ3vFPtJMSusNwS4VQx8yl/EK+XocozeV
BQili1YYH1AGsOQM5fynnGZaNmw7ZuEdxdSWsGH36AAxrPw/6ztCQNX+gH/dO+2Z
Y91REH5zGdGoQEPwKBv0TPrGRi90+MRytTGb1iV8MEeYo9y0qqeSYIbcR8qt0ZAr
PDacB079jZPiBT4XdZefbU1mFekhuans3mWleu8RqrgVHO3g2d5gFvvtYI/wY69x
sjtSRmgRkDo/hx70rYKIr9NIBv0nm9sd4mNjrndA9BfkYFHGklHcK4R0dlnXeet0
GYMJ6HbOoo3q3KbShAUz0Rze5lK1CmxNX3CDNu05XrsUBcQi8q7Zkxe0x6S4VAgN
dgguEE3OmTXfV+SjxkcbHfty0Ua0YzRf+QYjH3JB2Bbj4oOTtuvH7YJL4uQSkG/7
v6hVmJwS0truFvD41mdtDQ6B9UtRDe+zCZXn8koEaaBCu1BgSmSMxBrhAeBtskNX
M5PYhRmtB2hZ/YvEhX/OS0SHwfCSGLimpq28+aMDcJfzMVXE406Ju1kh4J5eW2gU
34owM8zXiAccZts6vM70SEO6ovKncjjyqO3PhiNAVQqgj6OhWwFJOGx3EyxtpzUD
47zZAmjv/iE/rCQRNyYZLJC//x74CGBki33Wk9ZuKeyclSrIgiOoNJuCEengEnB4
ggcWELf5erOwGcvfDwyDIzCZtlJ3pdboV4WjRcawQi1G+6TZOJc39URjA+AAQxUN
CQ3tknMukRdFld+fLyulLS71KSAXVVNgX1/U6dbOwN8YrPAenx1jGhUcwIE94xes
/hfxH06gY3HvUB1aOxE5WDnvz/oBl9GqIvG1YFSDzTuNC0ByW5Zjz43aT5RWDbDQ
OIJMM2p4ysMg+zNOdn2RHcrgfZ7sny77fU4OPBKJiJzIRTY9qG9PwxcS9vgxXd2g
igM+FUxIYIOFl3uvjo0P3oxZD+Nw5pbpjb6J0rq14Wzh50SYXp1AVJK+EMn6DIlQ
J7gr+Ia5g8tH/Q7y6bW2t9+O+E6fmZj+6OLGG7IWqVIqMUMYNkh4us4di0BiHNm+
JUva7ckb6EwcE3DuZjLK335x+ytgt3xVY/wVMPnpiQEZGDpohBpa8NVNC4OsFZmy
SOAd9Y9+bYuOx/n2jvFQp1qVZF7/GxJq5sUtOPehSFsrdubwGXEozIOZmnsiceKv
X5fmAtJOHXkZZ65RCAnsttoO3Vi4fb/ntOAEPLwLcirxkgAjnjUhRSeAKm7RC/0m
TwJfBB5OvRd35J+K4AekLIgD2ZkDPOjRET44L/6uWrHj+GmlskZvvL3CEofGVDXe
eOW4znx82fY6eDLJ+n9l5YyDlQbz7t5kcQdd7zx8r7bEr/U56VHxrjzsXCpjqJnj
1Bskicq0fgQJpE+X8yLHLPAXVbBPWmEDYpmbVI9XJp03uaOPMaFddtKfUR9LHS1p
Ng1R85eIqO9fl1KfUj4s3w/oxTMQcQ8PEHyEZ+ORx7p3N90tuz3ctwWO7PER/Mtd
CmlUx1kK2GBDjLm6a/IY+fmu+4N1ufZDoFu6Lx8F5/f5bHcrstiVW6HMJbvfL3EV
SBlVst1A8Koa+Kdrh2XFBV2zXTmOi1YPB0o0x3Fz4PV2cZAUvjte3KSbxuk4XwXV
PANmMkMU/SRbsSKyrLxwtUCxshzA4ChGa41Eb/pb1fYPWujsFmzQgxsGgtShgatO
fq8NC1PoQnJU95noum47ut8mho693DdI9+oXa/HmG3apocFgDWtbyH7zOU2TSePm
UMiGsqzWB2HsfxXsfgUQgtxVbPQ+QhomL8REUjzeYIxlf0degfgyY2oeDYGq+ZyW
hCdrViMQkZoLUdc0J/sceU6jsezfJt9UgJbevqE+HzH3LNbukF0VK2nmB2bfYQrj
1yWQN6s5cz/CMbTw0hvpFH+H2YwSab8ux6qUg4qTfbcX2cBMeH4hiCs+ujme/z/m
ZFbIBTbFvYapUxwP4gqy4TBf0rQK5ufqFqdEfOMNKN4XI1mgxOu8Nxg4ofxY6zhY
yyM5z08q4k2KrgPRu0lal/zWvFgEbjeE+N/0nWaKA2L3i6mGnzuewluiN4mrh0AL
aYUvfgcfNsCT6BXK6eMCHQA5p5TmrZvHyKMg2RKM3ggYjfPtROzPo1aRtCbMemC9
o7KJ9cqikW6RL7asHyBguqBBC39qy2iN1lKlwod9UhUZTrelKtV1y6+MrQpNFNMq
YSy+I1PGsWvI5Dk7jq729jpitF25FfAJ27RT7l75CYPvNuDQ2GvMxVWqKIKlDd4a
MrR3K8uO4AMMu5UEWeWC/A42nIOdxcipmSPWUbExdsubPNq8slEXW+fKRk+7H3bA
gaM+yHFobzgEmuP2mzYs8giFM+s+D4IES6PNiCkyuo6bYujLXnqZ17V4RelHI239
gJ+aC9c7iGPMb4fOJxR7o17nBHFWnOXiu9CzXdJrecZnNDqErZgcrfU+2p2UIhbb
SoJupjDXopNq/DuXuZc+1YuZXZsUV0XgGMaztrjUaryZkGJsLJ1HZ6sBKwGSo7cN
0YOTBFXsmv3WLp7J4TL8oz4el9zyovmrdCNG4MKm93PQ2BN7psLCkwuVVxSPwfEH
E9yQcp+/nCCCB9h0ATQKO8kTP1+lr4xuQVn500oiLtcSnNgT1dJJ9/NFc5QKPpw+
YYbyRJQXWCTGa0bIgrdwUFeZ/7GhcyJWeWe0xmg47cCzAj7JNLYaHG8eofpvQ2HO
q8WDb9v8dmJOr0H6qK4ZJphAVxSaI6MwNO1QB70oCEluyonAGDpZiIxbofUN3PCg
iz51KpyKo3vr507vkg3rVMYCkYH4TfgehBvEMy06PG0aLzL4qNdJccHKyjbXLoII
utcGMV6rdlnt8Xwmohb8AUmE3IFiMmJbFe92D2/PgajYMi8lMwWzwfMvI5qUz6YL
JDmEJVR8CxMs8u8+1+IBhYFRXmT1Y81GemSs8gniVj6zn05zxHgyy5juOUhZioMa
eD+8ppnWb8fmJfbf9pCyB9TvWTXRGipuaDriHLMf9vTKdmLfC6NFhmMhaFLH/i9d
HH1XvJXi054CHy22fsgr1FXuz7kLBv90cST/O5xUE4HLtLa9jVy1No6IufhbZFVz
KA71wDSeZ/FZ3cF4edhqtMVejebXXtcIjWfuD/4ahTLw44CfxKXRLBMF89DAuwx2
OFnd/qQB5MiBUBhDvHbKHiUO+SsyolOs3Bm6J92HknuvVHKGE8DEH0KIW9nJhL35
nb4+LMrG6+VY5ilvD1YstsvvfCDSUf9PQJS2HMHIxFqHdvUsWPzjeF1gTGzkkqyx
EqCNvSrOrdKZ+y+wmxDIXbyJQzIVuUjrQuGlIzrlF0VPELbWqs+Bn232/QClYeF4
DMcHSDOfvgqClPyBZqyBdMq2ZAkbpFxnm1UZuyqs71/6mLQ/vRo0FV+1YEsPlexw
s7p8NCagysmwP/scuGQZtytLmGBFZlTA/fzGdLrrw8uHBPjl9kmh8Q0Tjain3jyI
HYXwzpSokOV1w8zuNhIlB5at9DckfH1hnujCp010FDHcz+gITpdFKLgnsnQzTEej
9GgylxOfg9HiQtLr/fUrBj8B98IivMcravWiByyhRPfS66JYMU/XLIev3hh1n6tv
MaIdWqYsGzEUiVZV3Z2IC8Jkz9AbNEtKVDPw6NVKU//yICO+UArVqX9YeVTs6jvv
Qajjgbjs9XzFQzvyXW4DCbGEpMCCeXxPTV+McWGbg4nrIg7cXENUChmFTrmscz8Q
jHBcIb2wgfTWvyW42VmckFdQPeaIwEpZcblfzutf4lPerOBQkUZvuFltsWX9dMv2
FojD/gl4WaXPhqQjnopTtnIgd/0Mpg1sk5SOtREhuZtikB82NC32fR4XpNYPviUw
/YWC/Q/cEOs2m1Gd/Ka3q2WgS8ulUXFni0CShQ++Vw6WAjmGSV9gBVsLiyv1UhlC
AVgMsDtE7sJh+uGKqzuuQsBjKQAHExupImlKxh7qIorxiL2fI6wKE0G1TSxaYhby
3HcNvjBgwLNQ9247UFMKg7gZZouI8qQ8XJEFas8ZJdtIxmBSGH8hGNQ9Eiq/zftB
AGmxXRct7R28UP3KJFlgcv5hH2Gcdv8XUSRvadTQOb2Dt4ih4MYdg/hwfmCYSEaH
l2ZpaNy50/ORUppUzIHZq3JzAGCAAARhSVFG+C2qZAQEbdVhVGmIg8VNYTWH0ZUQ
e1GtCHXh66z9u7xeXqW39pyGZJgiBozTduGab3gbCZ1L4wOFdZ84JOTMcpv5bH0f
UeWZUvGiIz9p4NTlW4pFgqAzRDs1zST+kUvvVX89Bft2YJURK9SdY85As32oJHS7
rjl4aR1qpZmIaNpKcCOOgrXXsOrqli2MMow6dTxrcJp8cssialKSOMhPwWUtD4Ed
OHwdIH7GUpKm6LB6FH+Y+Pn/Sa8Cmj4DhLdosiO/Om1syWbcRKsVQ4T/VlsLtqJQ
+PK3owJ3HcvK+Qj2iH+gwQ==
`protect END_PROTECTED
