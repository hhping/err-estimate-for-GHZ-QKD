`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KlxT2wJufZ4N+ua0pogqC/huHee9roVe8O7Qu/U16CfGvB5Doe1Z6m1GvHYS4kh8
yq/XSE0ci9PJvQ6U8lkDRKdsb7Dq0ZMairip50DlJcY2Q85sDWAmhyMYXXIQqyBJ
fgwndHGGDSOeZDQegn18GOZA6dt8nvXCDJfOnMFT+eyNaFcDhp+KWku++uS+7g1i
imbEl/BXsfWl8Ab+yBL4Rq4TIvaG8xx/S4INrpygV0TS6RJi8l6PQFW5aiIqdZYb
PxUb3BR0sS3Fdobn4angFcNSXLsMTfTsN25cgY2CqlHEg3bTwj/dDIipTqCoEBuJ
7YTUB8T55wMljPjndgXQM3K+XlTsiSfcGPmzOPzZoK+d+9BTe5JEiO64hLFzvRCo
WpGt+D0HmEFvAN0ZctWuhzRMdDCYpXM1TwEFmSHO03a2ZdeF+yU2aY5J8XM0pDen
9jvOfM2m9sHBqC9r4w4qK4RpPozjJ7mNZvkxaQwTR4321Hu3K8d+oKDv5WNfVQsN
omdvS7mUNV7tVdOkd1SFbfsuwkfxFjpWlIL3H9XRY2YNSx19Qm9POqF2WbHtGkCn
8x6NGo76Ng0G5munGL6U8ig8ZzRAxEXR+tgpJhpu1y5aBZ4Rjek0gUTiGa8HIdQR
IDu7Gzuvlc0UNyz8euqg5H/aC2YhElXjEoKV3V3exuuAkKkalH8WFNkdL8JfAyW/
8s0I/vk20yPsISbWFam7H/Fcs6bRw3d7wa8Jqw8drqg2Ycqi3k350X8Jd7dDM1HR
WbAImfc68m+sitDUM5iH4EwjobgG5OPiLhP4eO2UjQZZbekCsbFGJymRFfYuPi2m
3fmDK67vkmfmCDCyCE1HC0OrNVi/UYzjwGL+XDO9L8a6hCkE0YGHWAD0zeHNl5k3
2P03HEECqfK7jXfHT8zxGM/ykPzMEYPvMeCKO8NDd193xAbLaOgy1DR6JrnYOtQO
saTKFOqQ5zpBJZZnekZ3QE9V53NGcrUb/PjFl6mTR49LP6rESaO/CSs+AeleTtHy
/ViX9+80j1Xw0i6NSOKM/GxyfvTtQPH3JBpIpqbQm8U=
`protect END_PROTECTED
