`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KzBfmrbKuqfVTwBEtt3CWFFBK7qenDyWqHiDKkbmUw8DuBPu5xXSAazNE7anu+pq
NnP+ZZ2z9JhT+fmEPrhd14Xjr+qglqJHhu/+rjh97poG5UM0pA8afUQKLFmb+hab
MaySmJsj6FRSziuJUifdYh5RIX6zb/i0RvIQfJ03Gkr0JtcLfo05HJKCIaGOn//Y
fgIicJib4REN1g16xcY/wbm7SWr2C3pNxEtEyud1u1MD3tT61bIZEappDxPWbQCH
MJE7+EdxKwQiSxDFGSN+VhmWa86JJu9H7kVZTIPkYCV61+5cqHzi2WBrEJLm/Zqf
hpy5rvUXgXQCn4kJvx3mh9RAq2BNEGaIXlv2wnUTXe+KQmrgox34xOQb77eAdrEY
8ICXEGRsHdSdaxzvaQzjjI2n2TCcvAi2/rJIEC2jzadFUco0v5ln5T3GbkX3UJJO
URgvlnykUH6C17he3uadtQiEN26fmmq6tDhcMnqn8zyrEBPEuzC5cG3YN3Z+Ua+p
WhUhVyA3UG0YM52dfB0x+M5bF1p5eMWLgqRHwFGTYBy6/M2CmrRATa9PvfOqLRzm
aNPoB8fQdCOUiGyoBebQIwyUog9Y/ehZxo1DYi60TOVLNC+LrlF7rw6h5BVLLxzv
V5VixKxYxGsFyl4pYxaa4/M33wHWm7pXDc55wovFUiQM8LeZACKEDo9FDxC5DInE
Aebw2SwwS4hlAXe9OYo9tfZkNznFVYlmIjpRNHUWRciFi4s4AukBP6Od21xNTC4M
fRp1tz00iKEycC0xfNgAdXSIfP/9O8zdgoEzaUU23jy1dzCinLvFPHwzfOFF7PQH
Y8szzg4SVUm5hK++Jw6j6QH2xWjjfXRtUVcG9yrG/GeW1VoC7tIjWSao3t3F/GGm
4vgmAeKRmj0VMw/DxkNAzZ9I3pnkefPStKQcUfPaJj+dQjKJT2rxzQxZ/EMgm02j
Aym7bMM7KbpkLXUkaIqMAQSsMkB41I5iVjc+2ibloxuoU+QQZgpO/QvLM3B8xhcx
TIazM08MObxpMNk0TDVIXZf/glC4cTPeyhcqY1gp7qBxos6kmRssGlsGhI2oLK37
/eOOo3EET+lM9Jc7GGhSn3x9rLIgAyp2KBVbCHlXpH8ki/eUOfPwGZJRX+Q2CAO0
ainUVJRXBIO2PPku8WU4HD7Z7uNcbjEl5luSHd0UzreE2Ho9Rm2763wU7QR1CM0L
yS6Lm6tOGbWcwmJSbGbc7j4J7iHOzrFQsjf1VHu98V8zAhKo3/51xdqbVdjDKaX/
jbTmH3+2QahxmAFIjMT0Q9W0/knOoaqErZhiuBRt5XrQOxApEsV+LpDo+s9J3um4
+CN2sc19CNQarz6Opmx9BE2ZoV8eFbZrfMmM50k+xh+EHsm8RuE2WdKqAOQLgD3/
n0Sm0dJfSWFNFmOfzXD+C/m/vw+lSrbn5mUmMyRG8Ngx6brEqyj+GLQTW5U2f2IX
l/JZ16TIkfLQQfkx+aD0KSKRk2dtQV7ijQlkO7lRBxA=
`protect END_PROTECTED
