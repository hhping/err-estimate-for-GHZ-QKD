`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kHu9O1YEkmSGgJq2EqL0oS0QLdYIrUkBIfV3wJD1RjMp3Id9nyJQDZcTtc473Y80
SIhNmP93qKlZumRJ4rlE+iflAXohf0r/bAFpsJ+jUvCI32bwSr4sha0yh9BsZWbG
th9lYsCfuCnJIHKg+FpPUigLPWhqMjc3/odp2fi5bIrDBaDbMH4AwCxtqdOtN+Xn
o9qdmOoBW2S2EdLvNQTUGXktMbT6sSGxjommIn+gH2nUFkbo3tySXpwKcc/9NE35
w4WslWaUdb3sCFvbh+UAN6iuFmNmUc/uuAzDeAfS5E97UAEVC/6TJohAcvYbCtuC
cw643ZHFEG8OrX3XVAosmZVTuw4HZof44TLNU4iBBaqRmUnadjfpOqTCLNZtBnN5
01C3Sa3bPFqbxtnyV3JgfSD41aTVM2UHNpkyk7cu0A2fYjKHZxiMg7EjMwPvX4at
kMCTWVopAtMDlEKa6waKXyWEwKWbot2p4dVe5ZCCm9KKyPOaLY1tQiAZQ87hxwSz
M6lNkRc2VLRNCrIZKWBHlgYSMmsLsk9fsPMVLmDOfugK+WYx3WSW53IPX2Q4JFnc
qyZmRsL/TGXuJdWSQ4TrP4ABk86BOSV5ZZi/FzOTPgoGrGoDaDwxpuqc3YLydXfp
BfXiYGsfKbt4qSBgsKHN4rM8BKECDNO6P/jT78NME/6HwUITExiHjx1HgXnzj4L+
Nj6n+abzuqvmQwPzyVphgkV0N7HfFyq7bQj3y1f0Z1EFOgd4zS9bIcrAxP4biO3j
LqCNUKUHzHsNhPZuG0msCrpHQJLEaq36rDd6+Ak7VCwFiNKCfkebUptwY6PWh0Sy
OAT2PuXaEMCBVtslKlWtoav1MpBiIQOjUU2cDyiktwl/e05cmxg/TXpSBBCk87I4
CpWvT2XnW32k09Mhs6lRpxbV4SUieUYLk7DwwO87yOQCEvmfXL5mdOwtGNOi7t8+
87xIUaFvQiXML8QCNyowMW3+i6+IUYRF7jwAfuACwjQ=
`protect END_PROTECTED
