`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QvDSXq8oHLpk3/nto23vkI7IGYKS6SJHg2z2Uxkj/e06q0T0jfi8k1XVcZ8Ci9nK
+3LcVRZbWnJWqeQbPZg7VktrZDaA9zdCgtxh7m22qYb5EMiTXFqa2dgKHEdaPUNn
WjuC7uJh9BENB9OcgaPCuAc+q9aQ/UfcVmgk/3yB9OQf/+ZDDblyzN8XHBo2Ep3t
GZ2mPQK6y2STzBOEHoH2Am+VgiYMYu07yXaJdeYGposoWKTrMuGL1DAwCPpbO0Oq
u7zqadCZ2V7IMQAtRwduKpEPct2EYzk//wIkQOlFRUzL7XA9w/zxknj5R2vZxsDD
FaxOVJ3DTSYG82z5ZJrcBdib998LJxxqrncRQxtyQFZwa8/9zb10/FfMBh+y+Lgp
2NwD+uc2kEBNgNojDLtiAVJBoQOPiOQ+AkQKpRFII7nwaJdys6of8NzHModTFXgq
XHDWuPrP9E5OzoOIyRDDecQ5HJa+/vrpkaCx0TqWs0iKuXwGFfUhHEoSUwSGXbgu
Oam6b0I4RJ27lwq2T64xuae5StMLRQ5pS8io+Bedyh6i46ATH1hBHw+lgfdL+3eL
oLTaLJ/NYCIt7OntfM0kGZTHAJ4EjzfXL97ehoofWdbQxovKVH8kB1aGbobGBQSF
9S12UHJyQuWBFCBIIXYHRR7kiirEBWnAbLt5SFYBnT/HneaUmyUorognYUr9A3qJ
K/sbSEkf4RlxKgw5lhgRLroW0KGn2c2qtZDKBNuIKK3V5CkVc+gVv/OYgLl3Np8B
h7IMKTExR0ZnhvXDmPhyD2SSQobH7kTlGDjTjky54eInDtMFOKqGPUB3yFjqXhtV
onOYBaFN8kWHBB9LWVYhfPhxChYt/6XIgKFbXUGZfSLxY+SnU1qdKXKSMkzcRlXS
bFsxt33h0KMgQ96jK3rgRDFAvwIBSJX0L3gcjSR8HpnEKD2uouOMF4EhvyuXDqhF
FCvzGBtj3P5DJh4TmTQrZz8Yzy6qIhEHVsX6dox+YXE5ZxJ5sktjzW2eU4eaA3Am
gJzHFG6yb+0rIKcjhZQi6iiZC2aJqVFKvB7TsiN9uOsYij6IiCy30vuk27QNmCUR
mXc87AkCJA0fvz/NkToAb2+1gCp+7kv86OThyDo1yJzQqRhjEgxXd/OlG0+qhgsQ
5ywgdWtTP+8EGJoPIAuh7a+FtQaX+J89xAb0SARHxyJIvqP+kCB+wKh2qHsJYJdu
bXlZyTJAH6kP2dhMYFFrbjEThftfF5TjM+c/H6A5Ec2t59zr0pbtGnFUIrATcksU
s/Dsa++ZDrbcxKrr8818VTOFAJpmnC/YdnH7y8dYVdKHkPO7GrAmK/mfDuH/ZjEE
nchxuDmuyAy9vAM1ZCeyhq/vVnsvXtZcOkHq22P4rKYLpGnSMFDaA1EaZyOzFLuY
h2l/psT135XZg42ROS1iSNzutfYck1yzZoDfyLI5PE3WiuwbMfpj8yH8BolFgsvN
RPYZriO3xtb8LFlRhRmYZjUPf24+O0YC89cwrgM2zHq/4mdLm/tgSVCPYwjy1koY
poCdTV+uGzS4vvVLhdppyH+/IL+m7aqbFkyBDBkUFcHDWYsY60c8kN0PjEJ3AtaK
yDxVfO3wKAuPmayoOz6seZIDnnmqXPZUH0vwQtVdQfl9NhWecRaRKHNkzK48kolX
47CiudQFoH3GU+TnNPWFHiHli/qSu8+pHYQ1m8gM+I3lc2wEPL5uTpT6HBLI4U78
CaBAtv3bmyUSMJ28TEHt7RG3S5tZbIlnsOOjkQWC6H0Vy/+Py0H8LrskyPeluRIi
kVoQE4ptig6VEMLWE7/YH2UsfpCvmqf2O9WXbzNRj/rmGmj+xJGI74ergkcwgeOK
LwUS6Azz9cHGBWFNzWOxsnuBfOUso/9Nv8yGkrxUy3Da7qoRmwAtXJ3gpR9ICuD/
GofFffviKzfrCmU3Kyh1SXRahenjWRA623iCycOvFRX1G9YBgvkjH0B8CzZI11yA
B2X4CiF/J3Q5BuEc7d6u6hCckCUky/UdWmkrYOj9/DGZ/9UTMkGl1kjd0aitFf2F
QmyA42hAItwUN3SAJKlu8EL5hz5qQ1sOFt366NSXyjJ5HQb4PsP1ohebhACf+Jiz
USclBfI92z/R4H7xKguY6TcFkbo9n7vLFEGFCy1eF3LlXHP4M/7quH1O8MrMiXmn
iqPhq2ZJYAWIjdAjUfP44jRQZLuc5ekyLYqi7emfkzylXBBEQMSE/OlbL8tMmsq8
12cSiEj9VdR5mZOe/+eDQWLJv73PNetxcjmei3BCSYwnYEYs+dwEevheXYCB0+Lj
XKeTiuL6KqNL1S64RsL+VDE0M77oC9nGvSvRo1EIRtxNf5g8K/VRAfHOQAiVXWUC
rpX73/fAsH9ORbLZAtE8iZMCOaTM9TVx0dSHqt8mONFZdxc8xpqJ+oab4UNC7ynv
ZFDgTOMd5BcxaiQP8MKg0pjGWeKxOVWT28sU+Vdo0AMM4Rxyz8ZVUBSixEMD+y9V
eZUwra+0JmtHbGwpX0UlMhPDZziQ07Kz9seurdxmk1wo4QLsm3UMqhFNtmwwEVOW
XTN9gCO5RAvLK7XhAOdo3rx4Ydpjs8ic+krGbagFD1xSAb7kuT6gB7x9Mbkcpw7a
irScobr4Buu2P+bWB1wKivgZQ4axsjg+2xgwyc+qQIrY2/5wQgYHGdlN/9hh/QYf
orMHPm85W1/TXXoUjvNZBphRstLYEW0Zh4GkcAW2YTCc0OAInOwgWKDwTksg/44N
oEcE7uc1klI16qtAKXKtbUBTCdokLiCHmAzQJ6HSo4Z7RjGPF9O5kDn+Be5Z/zCC
u4WmtxAvHlrV8h120I1ZCHXDqgM59Bi8f0K2RautHrV4TLvaZaPQNK9mh8GoENRK
0mCkw4yM7S6WEGqh/YJodggt8GmnW9cxUIoJLrh/PELyPGRqlq6IunNX+w0vdiu5
AQnozFztBPIg2oeMQWEA9Nczal6cdNyvEmkgRAqEoum527PxwXgyrK6T1YNl3OMV
zlcrd/pDwN4V8eHcav+nF5jiEiDytjDzG0IN1aXcX2MHP4dccT1tI6xqTyKydnL5
93ObZ2SOz4Vz+O79QlZmZdcVaNaxUG7/VxpnTqxEtmcA/gTkrvXogeWycbYwiD75
pJ1Z+EThCUsPLKclzKPHauO3fcJwvx9G04IfWJPEhpKg/FWNRb0p7jsyIkOFZVdQ
f1GmLWJwRRtg1U8o0XyNxQ+BEMacISFmBkvaHHPTfEFXmKK31mwgglt4lojK+A5d
Bk565yZqcXNz8WJcd2Ggnu5e5swBhsB63MNc9rQJorEX+lRdJESgdG6xwCyyNuPZ
TaE3YR7uKf1uHWpDkHLLkiJEODvXIEZlZRs2bEpPzU9i+6r8KU5ScPZAx96u/olo
Z5oB+/PtVmKnl2PnYX2luWZUUDZ9qjkA1tSjxrr6/ca5MeDsnelGgcX+Oi1V8adV
dGL4J0JnUEGflR0b4Z7wpw==
`protect END_PROTECTED
