`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NeocWDJMFpVgiADpWj9Tom99gzrPNQ1q/H09ZwmrY0TwcauYKUir0L1ieO0r5tm6
1Fb4C72/0O3RvH7h8QXLxOOb8Q/sKcIdm06gQI8WxdRYig67Ya0eyW3xZz25E5K0
+e+bsMEz0U2b2RhH0eZq2E8/jxlj+YwqTa4fsAgj/Cm1x7RMrH+n8CeK9XTsJkoM
4knAnWULbL8eXMNrlS3vAqEnmbWimMltaI1ogzyQr1vbgobaRl4Yn/Mt57sNAG4G
B6U3jXRjvwqztS0qeTha+qtYc3zU4kIW1lMJla98IGPrEFNQ9nfO4kOROsf0bITM
SwOs4Tti1KmITRnOsejvudFL7dDao8hTiPci32wVKKmFQDkSuDmkAwsr7MllkYT6
yqRmj517GpYjuXssDV1Sp7piaIQ8Pikjw6Rzvo7Qkks9BzmOf8aQb0RvvXc2bVJJ
cA1kZ+j9qHP6Svs0F2VEPytk9+IFXEz5+h+dH4RBs8mxnhMOdFWbfdCb6FGVJ/5c
SSNV9J1M6lNpUVwN/sXgD9v0kqTXXM37jFpPTVGdPKc1/9f1LXjT+miTiq7zOFCC
ZfVwPYKrOjwKAmDsf3YFgS0VWYyx/9/9nbe0yubxFyzQLiqsx2JJ6+LpTiC+Rh1u
XRFybYSlpZIqMjGtIAMbQuv7CDB/xBoTmVRetU6P++Q+Jw4d+2gP+DLAg2dYskbv
O2I1NtwcnNKyWMkXJFmrjJYVswb0pukH3II/okoVspSHrdRy/AkRaKvSMATEcBz1
kaokhwFxpngd3Euhoc1+bklSPaanVHX1pbUQcX/uqBeX9XGKbNLlEM5SPXDrvNdh
nW7yHXKwNP8FmwcYk/Ui0xUQEzlLmWl6t86CsU2pVMTgLiF3DjnuaGzZ3saHQc8i
n8RuANvW+8cRpoWmKXKUtrz3Z1WU8LPTAcUEyZKz9kWHF9wLrbc3A39CPMn4x924
qzQjUrRou+EKQFe9Jbzdij1G7io977eeA3uHcllYDvtclec/RS/vlbM+OZYlWhlp
+uZ8Y2wTQFSrjJrqQvMgAdWtNYLBTGdXxKNPufV6xQkzD1cLzZP3vjsoO9nFO+kp
YVhZFYJqzhM+c0mHnS46pJR6SlbAmWNr6g44GbgBTyt1ju2rkQJJKv4lZJHldCsT
vu87ZYUzGFq4WzsCKuZNDDIjQVJFJflFHuVW/yqhA3IsWPuzS0MTBjqSEkhlGvmO
z04lwuUQTpbI4lgc7YKX5RwUHBRV/AjxpVHHEYRbTg5ju32GnnfjcoRx9BUQF++Z
IQAB6ZN5DKK+XSoifD/4u7Qx4zNR3vWl561WWMVq/rL+OxaS8rGOLCxTJv4+Ejvo
jfpNwpQotmNcH2OQ7PcvP/9JnjzJsVlBZYbH9nI+hNgeyt4ZzHriuCCg5EYU5Kyg
V96w0SOiJLJsScnjEa+SF2LWVPeCWlXGTk9bNEKSwWraKQPHi+wK1ERmumPM9iLk
Hh5EVUO1AaX7a+7ET72QQJUtqdIm+bdWreeN66D51lnGFNxW79Yb9W1njaKD2ljb
/hjOwM8EyIOtCUrqc5Ds3GALwsLtbQEXkOzh/NSFosB1dg4lXqIS4Wc+Zpjs6vqS
XCfCrPkFfOhktcvygBQ3UpFla1/Aw3iGRbXQ68WrzSjNyE7lPdRWa5KG7loe5Z6f
l14bK9LguqQTEKdvC3W1guKjzv42Bxhj+ezXMKNO+r2nszx84EtzRouhgxfjDdMi
io4tZZLRUZic3hpxInp9Xw==
`protect END_PROTECTED
