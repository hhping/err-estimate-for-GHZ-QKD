`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MyH8wuU5nSqTWYWvWhoR2N2F2+6YNOd4dGELzMd7mONDJLuHX5DbI6CdYtnh1ZzU
8qXg/H19NTEKioX0WZDxz8NsbHcwUEbnuZozaqqVHR553BeNKtWg0R69Kvl4GfZw
Lq+rA4OScm8KMbTvAbBJ8BNyiwv0z65qRXYu/BAqSbkJdm3j4BMccpO9cpqBdTql
3RACMtCAutftSWTDPoI3HJaiy1XKGTVgFi7u4UU5Tiy0ni+DX/CBe7eRti7PofcK
swc2K/1NmFS9/g2sXAT/JgscX6uR0yKCSEBDvoFj4H86DSxyvPROuOkNsjTWpMYR
6cUz4/xRJOd/V6so+hkc2XvihfQwS2foMW3UqEM7CDzSXXk8kQYTUYXnbB8LRVGX
1ENkSr/6h6Q/cAsyj5Z3pLOvE8/ye46knd8yu9Tq6MyDEYNWuRXY7eFagpWdfl9h
FDnejQQ66j8nfqYp49jkUkR3KX8PmH2wpq71xNHmlVNrcffmxR755aAAeYj0YXC5
uX+YIe3fJqDAY+xax/mOMJOtH4Emta5QS6KC+aqBsNCtp2R6Wb8itvijUm7iW3MT
361LNiZ7GvRuQC9y420GPuZO424G8SHzbaj3edvg4O8RFQkyAruMsO/KQvC+SOB4
`protect END_PROTECTED
