`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nsrbsxMbO96asAdddmDyh9BZMlC5LjzyaNZa3kAl8K8GlO4B0KrZOq67NnBHddh6
ImQqM51oF6yOT14LwtWIBPPzr9/8Xkn7JB8y4EI2FO98fSyzPa1a66HqJJaO77fL
ibsatqT2BpnSToT9YO5/aaR5j+mjBtO/oPo05rnSjfGcAYLtlEkByu3vGvG6mtmd
T7GlS/eEA+TaE/c/ILsfo7/5nL6RiuqcTTdM5K/vKjoDVIQRV7McbvgGqb5+k1Fs
x01m2KiDAgGGAcWkBRb7HX92r9RcmuGds6bFBJ97d3yYsBQsXsJZdrP7IVEk1olA
4nSjNekHyKoIFK7gMICuo70Q0U3P29K8U3jmGYELrqZIVuWEZvOs348C5A3+cE30
vPB2LIfcjfl3Rzzfk1zq+1kBb1ixDhCr25eORc7nGzAW61uN6keDdzQLO1IFYm6m
0DhiFb6AsXorYJFpRVwaWUgWtcl1vzSfa4TowTWNGC9sPAcJaM827455xnzwyjek
RuMp4w3wcg/y/ICa51U9YwOoLKGjr/NUbl7RBzsl+y55bDYNnC5b3Rr1hULtxK4B
RhMGY5sZaiOGrQuxGhC3ZXrB6NAByTdLEmM5HOIfFN0ljbYaMm6WvYqvnsUM2tM2
nWT4WMENPQYLEwXEVPApF+M4rb4CP6I7TfjwSeRjgB/z7zUUqldPsHR+Isw1UIel
uOAO6p/PJR0b70erCp4S55+v4RT4MqxMXkvhVZtJ/Z0EpP2YuGoIkuE7c2ISFOW2
ECdqZAfNeUdbmaKGUiTMruZwD7BOKRDB0akjAEzNVMVjgyhCGqiIFaxfozI8Yzwh
11CTipnXtVss9ssYF4JC/Z+q5z2p8diOjkGkpY/Tz1dcXJyIF+Q9g6DcLWUjEhbw
TWP/8Hfncx0ZOIWfTb1iUaEHhHPTwzGgd+Gi6UFzIG8OPXRNVzzX1enrSJWATqJ1
Fuq6btZalx73buf7AbQklpe4aHyt0pi8Sod/KZYdz1Om6x3iOBKRAI78B5WzNcwg
FSlXCyMTdy0o5rEqvjfSswbmXLqGwvEDIUVuyoEDmdxd05QvsflP0AGLaiWcyaLk
Sm1kAJlJ2u3fRKCT7gztlqD33bpIaQIr2cIvgPTrnrrxmUefecST+gd9udL55Dsr
tkpuND6Y2xBOEVPvIjVH8/y+3gv33Ec1btzrIIpMepL4+GX+RZPhtK6IGgJf5V6I
g4Kyelo/2OFgc4RGYQNQJWAhzBDjgZ/WghtosLDspYYoYu7ODeQK5CpggY7nrRhk
qPiQDlQwTusefyh711SdlC7+vyaHJXqpTnU3cDE1SvJfXb8/ZZTIJr5Kn51B//6T
e1D+wRIyA27wb8a+Q3SemFmyYV4W9KdX1hyVygKuGAkj4Mf+0hkzHXZAFLuKRo7t
dMz6kniNpHuhhS/k3vF2ukbMNWa1hohr2OGQbBbYNyc426yEALo92UKYgci55wI+
Rob1hN2HVkmt5VpgG5GDG14ymCMugtrEn/NPPrrdOSHLyHKmfTLn3nHq3NIM2UrB
j+SJ8gf8ZKpH3pHVNV5sQMN4iAAktSHc1qRS+gWdc0m2wmefo8Itd4ROKIbGkZ02
nP48yHFLEZ5qTLYjMlkO9Aww67R8VKR3w1KbaUAii+Ds7P8WXJbzet5LFnY6yEhe
fNAm/TmggGcN8NeD0cgPSs/jKEZyWQCMKf3Bv97hKF1kxu/R3jMc9HEO2U/+LT0A
AYghPWTgITygK1s5+EshoZn7oTYb6VeXUTryfBjeAgYWJbl5xdWHB0W1lv3kIOVJ
6uX7+lLOYMdOESY7nb6oOUcip8KF+FVaB0j4NYx6guf3oMU7J9U1RadcGolF6pB0
ElRyuoAbt/QYiwpS6sDJnCHN2qfrB9A8KULnygg3cfnJEmLVbAOGC2H8BdBBtCR7
yW+D2L7EfJo7kWVhcp0L/rqA/pruqpv76Ft7NBBGwiJ6P87XfFkVtV0CupaJzcRB
5UxW4r+F+2NmdE2H7U+I8aMlugOV9tQa3VbEjMQsG3f3Zd3mpbMtpw1Mqz1uvy0z
ohOUlaP9Z0OH7p+jx4G0Jh+A8vCDrdhctWKbzQ1XRm6hlg6HSsa/Qv66fBpIyQ6h
EBZ5lzQI3a2LuHkoFpm7oeRZ9UsWIZ9hAnfFAlQ3DbtR+N72mx8CU7D/IgPda+Fs
ezqmJpXh4cDwf1syO6xuwsJCPeVk6J3FNpJpRnlSfIe7ng6mk1opt6ovVgEuDWsH
6YDLKS071s9QxxDlUgRfTLPwjqs5dm7dgch6+n/eVfrWiSG6bQCfdfXHXamAyjK7
ZaC81AQvQlrG71SC+dJbvDuQ6Kf1bRYqS2Ea0+t6tACFssAKk4Gf3ksNB3ALjyua
xbLfGvYpscd+eflCtqRDK7bRW3OrssIsc+4tPjpHofHOTs5GG/irl4Pfh2xUyTE+
Kgv4afpBnz2t616gXM+JZnG4NOF+9ZQumDeV+09RDV56MatX5JC1XEZjSshBOZFQ
8AVMvXmRcO+QUjox4Y5QMy55DZBMDZYw/LIyZbggM4szbNvo1MhEIJn6AyKNAT5G
p4O4SoWfwAOx8itWS+LZLCCMRkjW0GA6lzl2RqWhpI8bLR8qpOYual45MIA3+iig
ae40sJeER2nXmkC8Az6G5RkP1utBsQcPA8AxMsGeotXYw2rBPn18oTZ5CCOLiZN5
whYh8u+Fv5LFs/eFDW0CBMB2VIHLQxtC04fdaJX0rKXDwJQE/5htK7OFIk6Ij2fK
vRYHzyCCuRWznY/Q0/dUmIRov/ItekmuppQksndgveonKJBRcvej2/XGy9MOyjrv
gFVdni2/kJ+mwi0fQ4NarZrAEuZubzEGbi9nEaLtOjddvwwoVjR22nblgsyNlahH
Ipbu8Q0zg3I168a943Uuu/XvKEKXHxKCt63lKO9ECK4fNXD+jtep/Ck0qrm/v8cg
e/Tg5dOaBOuuHQqtn7OKh7YFeeo8nEnWoAgjJ4fW3MriX5pEqXLJVbj3B09tn/6W
ePTVB/Q+VITikRMo4ZUvyaPpkoRVtMiE9z/cp/jONiWcqA4jEFuF+01HO5vu7zKt
p2kedUcSFvw+G9O5wXX7tl0caLnqDeMqGPJ5tbgTuVnkJ7WwgWQcjqtcfBvvfAQl
oyCXv2X//Qd8GfPKk1ut2xrzqozHe2JgM/uBQ5ZheF2jrKJtVkvgov1QTU0PTLlF
/z17b/re6qafdXFGvFicP5/+bCMDRvc+op93KcRGISWg9J98JhS8fM4HOUayc3Dq
P2yqGwLMJqOSWN8zrnrLqXNXkInBYXYXkGxDDiLzrCwnxyqJOrQTRukOG8a8mnmx
hr7X/ITFZU5BjmupwmJcjxJX7HvqbkLV1lhLw2N0NY9gqyZre37OQPhRhag20lFW
DQEbm6+fNZBuqpTD0CwOAgtPdI5c+TuY8xokcZ4+vP7ej/Ws6313+7E1Fped10nM
zfh7/RriKyNzlUo+mJhLEqgsHsgj3xkv4QppkXAFp6MaZPHsieNU1qSYPxvkYF02
SjWmtbGCL4yBo+XLd/BaZfdrK12Qu2FbgUsCugNxOZ1LU0+fCxFNXrY0yqU9meIq
kDTPyJ36qe0dMP5mv5R6iIqjooMDD4YtsduJwFeEZpby+nQzKu5ddK4AZ+079el7
6CeW15rgBknz5JhgNcKVGpqAUC+XAsFWI8cmm/K1IzQfSFSkZ3t8jCpAU/oJHc2A
o5HlKGLQ4Wp6GJIlSbZjTxvRYxyRWJ354IskPi+lXlDuIY44qpfuWXJ6OOW26/BE
TDaO45CLwZn0zPFVaKT2soxqLBi/oDFM5VZae1eCteHsw03aiC7Qgqg55RSQuOU1
Aof6iG8lyy1fQj2bNWrRvUZxeJwgtG5jAks+Znl/l3SE8tW5fn+6XcYFxBn8bunO
4gD84WoDJzJ7aVkq5lgWk+Qm3xExWZeE8mKtkzegloFwltVs2AD9G9R70bNCtxAt
6PbmdSDwuKT43nj+UDYFHoFm0peA6ujKkC/nDw1VAM+IQwmb2ri678eQPrVt5vLG
z8OAY3vJiMx0qnDy+5CQOoGky8C94T4dUG52pf5F3wHid8w4PHQpgyuZsc1k1PP0
0DGRCHMMFkdBQcvnCTfmMtI1H06ma4udFtGKsq1MGYGZw5rxvqFtmK+g5ddDYNJJ
SDA4+TNz1l8LGjSjzxnjnJ/YDnSiQd7Dd0WxhA/iBk4YkGHiRZsemxA+OERVt2NR
jLxZeFN/g4pxW4ka6ickKppvxiprtAwW9miBeapI1jxoZHNb8OTMJ4zRlufGj6uz
Daqb6LiFGLxCl02B9G72BR185jnzozMJlr9vmwtcT7yK5fVsobC7UxX9WBaSks3N
o+ctv4TWXlT8vM2WfQfbJJK5pSW7NXHileOOBsX7rR+/7VPAmq/ZTrawcYhMs4Ec
F4nJSB9adk7B5cuaOgTliFArAte82vJ5mLKjbd+3WsITwKY3E2mQr2XuYavZ1CLZ
5FnSo9LOPuHMpLC5GlqK+FZJrnhIiu1x9rWrpWdCF7pX6pRchwUZXuF62aQs7akv
wI4kL+CYn/1XzPrOdRpa7KO96gbiMOFGUy9tIw9q+MaCvjucvwkfAogpW1Chv94L
XjbyNtLjEpKZj4qH/UepdR62o66jtsVTM0pSaVXy9nGkPA3DUsF5lNa+cOfIu4gf
rj2QYrqWodDYzRMvGQRTZC39OCgZoqAeFIqS+cZafngFTjoAHxayVxCFpQDYRo2l
LlmUEU/YQIPKJI5pUYf09o7K9fpbp/8JaifC05HUNYSnSVXIDAwlhVHG7GnnqEq0
3R2Iz7pLBGNpVmZhpCwQlQ3uFjpxX/7DZNCxMyMeAaBMR33u5Xel2Np6+ZTZTr05
ZEls74HnrT6BKd6Nao3WDL9oi4yBmpZG0BxGxpuD8IIMSvNdktBMnHHD6it54/Gi
7JQqxAhhKmDiv+1MSUswakUWYugKi2cOpvGMbuPJeYdNO2YzTf6uA3M5N5lRPE6Q
s8TEAqcmdcm9hGnJPdtkSeStBkUuuASA6oc+cXD69TfJx21utqNej9HkmY9R6wyZ
pIZa9Z1lKwEeofL157fsG4h02pvRLGVrsorgfTWqdbz/BnpsZmER6Nc9wskOB8ox
9CCGzBZyBpV2H+rQanmPMsHx5RRLSQ7iRnMQoJ7YBv00W0OMN/QRUhJRD1JAHCUH
tqCkLqDAdCMRr0XUis+o3dt2aWFIsvexkDqC19LQSDrRa8SRyA3qD7wi5s6eDH2D
pL4XtQhWETkDI5no3fat3CbqFKjffTmVRHdPCkVZ+z+Wg5qoCs+jrTqApm+noRcg
h6Eqa5tf9osbxLXG50GUVQUZ5lDY2Jex0jae3zP8mqfUJdW3EufqjjLRBgHG5tqV
eeJ26bGHX+Y1uZIdsIeL7EgeH9Bk7YCNtr6/gAlTqAppmZc40zqewW9u6g8lqFN3
FG++E7PUAE7/HmGStZAHesfHU8jVSbkj6c1OIvMNzT+UcypypAsHIPCfsrNVOT1Z
3HQ1wNiDj5kcpf+dgNjks0BBnsGxBwGxOqoocZAITHtIuqOZJLJ+7y+aGeNLviZo
G3N9YsMKrYjFCf/uWus6flyqtRXEh1J38iCvK4Azyhv2wmQj+sDsMYbj2e+T3Gnd
j+CTQB+LVkVjAP6d8nwHrE0CEA9IrHjD6Ega2y7rpR67VBwHybaHEUbjF2VDZVS6
u++hwmm2uYKUSsfrwomE6nS8neyh57WeczQsqa8OUA+g49QOhUplJPTUxExT4z37
7eeZGNxzCsdJ/08qq0Nkt6lRQc/WPaUiEWhEl7/qOPmBugWFVGm4h6WWmJoFSBd+
5Xajw9YWIDiGL6+3KPmkXvL/TldIfvPnxSEtX9fkwsJxlwCUF0D8a8iDqV30KQTj
mq3luHsA0FSVss/XB4Dr/XmUoxKxbzMCnFM5LXq05x9MsaDKlimCQEiVyWBI2Sfo
sm/kXqq6kc/IOtLsxxSwAICvXbhoaFdeYkTaPL26ywPDGxVrLmcQYwBO+SDMBFpk
MmtvHXb3/3amaPgTirfCv7dSAvXONaiughgfUn4veJ7ggZpt9gH7rxMG+wgEYo1W
XQTvGuouaW1pX0ea0OrmR6WrD5KozAYvQTGWHr6HFVLzMDjz0ZCtUOyA4Bq5XYRf
L9Nw8MMtEuVTlV0bf1+MBCX0XGv6yaM/QHliW8FSU2KmWyuBB4+XZtFPaOsociqb
cogv+SE8MB9N57xFAt5KlMMmiJSNcfuY0/sdazNXlo5hhXir1nJoTlZCFvR+tzkI
lj5vbYAPzlcVm4PqhOpW05X45/BAPB6v0IdAQwIp930GuWrOaxmhDDjUOZ/jjUaj
mrfoz5gP+kl7dEy/Z8qeJNrA6ftZD/C4GjV7f/3zV2Btr5vwkTaFlIFQIkX4PMsr
tKvwiz2uSaBTUJQHzs4u0clHpKt7xp00zukQJjCJAv43oZ1/5ZQNM/xegJaKFgk7
f2scrSuA3TnWzxs3JUIzxQBUsHqN+nnuCec0VzNoGEjgTvPU+nEk/ZUPe8GhlZDD
8zl47E/t/sYEpyk97etqtj6HwiQp9xRz3nhiP3SYBItzNeHk8hMhpdMx44V/8x12
S0bzymoDR4k10sUO0zdbfHAj4gOCsFVSaQY71BovHaHKCzwN11S9RuvpfJ5CjbHq
wZydJDMpdqS2g2amecZeNs2i2vJcYblQtQ3Z6jRT5kiJtU2EFaY+420xGgMaKz5j
Tw7iydWWV+UW11GTRX8NbLVEh+mITWAdio1mZRqWO6IRJStEa5OLahWRtpA4BJ8t
5kQG93rbrdbH0t6Gjb0QjrJTxrl5P67kox47l691Cc7e8gTKoejRfK8TdMyFYoV0
cqL7QQGohuNi2R9VnYI0bPMFRJsb7EYnW1glE9KtjJrpOtq2fiFcLgOeu6xU68rS
vEdYo/zqjAmoSJkg6XOz9sst66ywaGp8KISxHuP1gD6D6dze7OvjcG+dUdpHGjCn
mOVx03EkGNX1VwBLSs53gV3PGGsTG0hwkMATndjlyqZtKwZ8CUmbf8tF1zziHJx4
6rmtnuSk+WvDRQraLcOXdx2jeKg+fBJi6LkiT+eP+nk/QHePjs8HKz0o62uz5PA1
r4TWbdq8qERmCYw8dsbKL3DM5mTzV3Zn42JwYrkdKj8wcp1ODYQQU6h83dYXnA4z
7zTQ1C8ZO99mksTEkfnMNue6jySlAIri+fQYFwFonYD7o1CBcc9awdY3zDNThWMF
sDNnd5cF7pdcwH59A/bVH53PONk33meXn65w0r6rnr6A/NDEqOcg1D6W0m06Ljku
gQnzREXUB6jEXpYUzRjCjUpmGwKQO5PvmY8OHN0InRqViH0vWCpSAE7hfwV2SYwo
Axw7vOcg858Blhz9eTMgcpkvHiSY7PzL38XWPA8ooMRUHHA13fDu5S/WmxHXHmNz
rpVo5t0wG4ekJaEdouFk4frB2N7tjoLFUNykVOnrwyKixM/8j7vx3OQWH3rDnfjo
DsFTZ1Mpvq05rP7QJcX5ehXtQ4P+KZAJamTHigF92BB6/hF/gdOAQ9rO0UpOcqbu
XFZSzWaBFEjZICkmPwutfBnqJa4aLE/73er5hfstCXaTdHKrtirloCKwMCJRNA5b
BBEMoSxoHNgfpQjxEcOtvLZ3+vF8VF+onFr7gQJux0rtMO0tZZ83DGZ5PqViVo2s
7/aT5JcOEPj4hqJO6icDrgV5FBvozFAumR2k4S88kHrm8qzt3CTMICAfbftyfrcA
HPbTTtvUJe1QVcd4BfWaLo1wbAuol2org12IU8QTyS87R0t97tS66dWF7QNSFX4q
TcabyVGEueriUIkRvkdjbdhqCAnMCu6kz8YKA+9aOv6URSXfqnEtvyBtOD1Cw6O5
KCGAOuoN9pf0yEjwv1irF87oA163u7l86xY109N/2k1LCjgPvuSooozFrd0vM42q
2qDUbXoXjrTGiEWOGL6928p+Auywcw4UEb8pZIuRopKK1T80eR5gH1Wc+02hzq3o
4gvONxC+SxjS9LrhBc4sbFwpoemsx0xIF3mrkYqCD6MtHxGSpM7zA+XhYQy06ge+
Rc9fA3LSH8+kXiEWocqV54CqOdmUiJAGsbqSEdIvqirpFXkUtkifyyknNNM1p1s9
sog6VMdB+9aQeT0GeFxYrfTxGfK1JlK3HgxyH4Sx+ojGzWiZVR99asGDxV9g/eKN
yeEdTQI8VSsnrPalhfTN86pZBVpMszIUVLeEMV2iNlsRzevNSrvtsOKUY+6SjI1d
19TFfYo+OVFp/sXWC0VWRt29n8Ie7IANzdbCjJFzaChHZMXa+l6RbTgdW3wOkpsC
iO5xjfnth3dcFMvTZnIzEab9JgPiVHlVHHJANkgrn7XK6tjG11E8QEqT4HqcjTuC
yMP2cM6aYSVBf9SjLteTRdhOlOeCfyceX12s0SlaFjpf+1BnlJ4c5F22pubgwB8e
SLL/3K5QkE1Ff8Ywzf0K2Z+NApps0n5Q+wygvjOvr4jxERec8Sz2qo7BkAROnmUW
pnJG2Zv4prbdMkFMBLWgnuVZFumF5R08FTOGkkYJTRxmWG8i1/wsVagxJAhyAsOL
+g6k/OfsrO5u7b9LL6UoUwH2cDXpTOFlQRfi/1HorkG6y+0kVMF+JuZEotFCb7WD
V+xjw46bBb/SdjhYLmq2EjemmdjShOl+QlWPEbmdjKB0/T9oMj5XoT0G/06r9FI5
uNOVoqKMmX+bBL4Ea3lSaykMeYslIp1X/xmmZzZvtEl0uCv/IWdmZUgAEZY+9Tug
winc2JiPMYvrAvzuKDWMBLwvDVXRsW2JFig+yR84ilnZsd2pLaVliNaWFxtlXmxp
A2rEhY103+7Uaf+hM4+88mZ5p5/RUvJBajnowJj4KmRxTVKcGAZu0NImJ2xoyrbv
kvsIADZMEchhe6r1eRtseXLXm5QRMEGhtALxBEypuSTf2d9LJUdpbTJrZM9vXGJS
istLADK5VfPDf3NX1Kq23FwZeBLwI6+dOmF2haD4+3MOtwcntp79PciYl06D6IxB
PmslDSEDfu9sihg2Y/xiCAEoA/+W/goiyDvIejQI2nmr2tX7qV+Zli+ffxJCLmOy
l0WMYorA/XYlrEX7FA4kmUSrdd+2FzbNlc2gIF4A7poRDUn7my57WuzPJmHe96g7
XrWYMmifdigb3HzPJBcUWexrY7S/Bwj4dwgv4/T69BPhFV095Quw+4Zd4GXw5oq8
0k7BHrbIZahTbrH49im4KepCzYuzUbbDGO6Qxjd5Ket9Iq1jovW6r+tpmzKMLeVx
N61zLC/97wos+A6immqXZNRp136X8vll2CTvAsX/nkmPjz/DUXrXlAJYtq44/0si
vRXaHk3oZ+BFHGDl1u1v9d4M3V10dteQgM7dMl8eiBrFoAfat2CZrZ5mVfEYbqNn
Lb/lnf7ZCZuinWPRP1lnbaJpavkXT641wknhiS95PB2qEB5dw0EYbQxQUUmiaW/U
/+f08gcsL25UM4aggP2/FYfVIc6wisM22L3tDOMz67Nyo70vsu7EQYN0VQpfRaxW
ue3TqnfED7ney+YsQFhMJJUJt8i2hCKZYy3bIpoinrRWHGJO/XrEJmLgPf8hEMOR
1BsNnJEk1jmukgttGabkaiuoYI+ZtjfAPGUpuS76s7pNWxN8quIasQ3nvr8qluSY
gJkDxv1PN6OxGr4adx0luva4YyD5kJ9eINDEYRzGIzd3TgV+/Olt5f3pAJ65ljZy
xVfSyJmIAwIOMz6ZFujw19mArSUFMS2YiQ9U52GAPSeIp6guQBS+v102VCs9vcqi
tEpuuDsWTvCR0ADx92HMftneb1wCNGq2TffsjNl1/+QdQodBCmlAyyuwXvjnDizl
HKF4EwW8WZZA5xmvsARG7uoBOg/cwvniHOKl/ahNqhBczL5tqvQjJn8sVpqmZRxE
JmYBDYk0AWa1kS6OdVCuJVfJjwlUF+BhmBDksg9DqDm3e3aw0SUy8o2Pl/xhUsp0
i3mzxH4W7hpvhb6vUD8C2ZBepQSPd5w43JCEYlLNa641BqOoruTACywSJ8xmzxt4
hfl8UwUtyEg30/87sd8AnFlC0lUREG1FwJiRFvdxDlxRLrDc+r+JLS/C/su4i9QQ
CcBBSuCvEue4YRopWhd4Ok/Pd95v/Gx/dPyn5D66df7/R7t4pGYlRcnZLv4wd21S
GRYHJxZLwk2YNft2B5ajfE7q70CbQ8RbbR15UpT4F1mw93I+BGJ/M1MSpa5ytMyL
73pmDvGaORCAchjxRzc2HxAIIY44nCq+gV3gIP/JCH1AM6JlweTtMLoo1UTyRiHE
f9wdPAQOIam70bFk/07UoKkz5mpUYS96x7L4baeGOav+5ZTWc3mi6mSspljEjipr
3xvuKA1zhIzOWgEI6GBQfpSMIEyPtlx/n8KG3tJ4PHxLsoT6PVCKpUHwVHKUdD4O
CbmMzd1DeK1zdURaHnkIJAXrChQrr+IVBBaprGQzTxI+RxBlv2waSfLgU9x4X3gY
07dk1jLvbZRnTSn94vbnyPss9xx4nwIGEXgMstC5+B//n5buTg6J8VIR9NK0NQV+
T7CYJ0YC272MUGxgHfBpVwa5atZaNisLZ1TKz5nC0/VxUSTCF8lb8BQoGKMsksSg
Xyge7sFLW4AhuBbJLFJa+hvKJ5piSq7Vz4SLtoW9Kw8rDMQu4uO5b/glSHuuf3qj
tEL8vyClByj4MfDPHa8E+0+9rOuQQ4lIgY+HuY+pZu7oxy6ccOulIsXmVWqfRW4V
PTMUaYcDBKRoDsOM/Cku20e45Z+aaOkpt1VMB0epKnIrgGdEHCdzZQ+ltL+k2y7E
u+gxdxXKKZszzhgMvxbwpC8KbFlNFU8ZMpn/2TYw31KlBJxYGeoA1rqUGdqrWVru
ZhdLUWrOL5l9SPSqHYM/YEk4J5x9N+0m48Bx/VqX4Ffe/Sbt6TIt3enCGSe8ZvcL
THOMo+7KgXkTVVD1vulMAnNt5jrD06984CGkv1x7gKgTogTbQ1YrTSDQTq5MxQKP
bfDQDPmj+ZZ1Pj2ZH792IimN4V6L96WvmQpLlyAmDqBRn7mQveBaS2Nvl1nIGi/j
lhcnrtmokXbD2kE1Y2RJzGKnQX1A/mK0tNgCItHCRH9CxMSGbNT/+FZwFlkyXCJ/
GauPXqGnWQd5f9VXm9KNnoHT3/D7pN9/It+IGkhQNKDzMHCCt/LIou4IADqXDuRJ
B7QqQsefl07BpgsTE7hgntaKocqeLrbNdAjN90y36JEWYwa16Oi9qHg4P8D4l0mj
xEY+85y3Cp1Ky29VkqazZvEzCuDZquaqQR9E9qfIB1A/aVBR+5qTMh8FAVBRXjau
oyey5Nxs+fbWNnSu+voKCu4Arc48ARHP+1CBIUnXXTj/+eWI3VrZZNYVfBR+0ArR
wyFcGBf8C7xHCeTiBPXhoz8+Kvk8Ng21qNEF+zYi5ZLE5VA3UlctKv/CtYm7XD9R
uS5fhfc8mfmnVKvCb6mc+qdMIep0xFtE1LF8Vm806sdQrNmL9wfdK9oZnznXTJdL
RiMuw0KTql4JJq4aDKwranLeEgItGXvIANhe7A8KcWyTSzf1kwaG3OwXegH1D/Ds
6XI3g126kEGHx5uIYzC4i4lKxtl/uCjAEO8TYRvALzohtbFokSczm4+Qll1jXEW/
j2AJLVgjEJPckFtVgOdk/3DvTNGAZoewJO97lOXl84O1jTXK9+LH/1Tsx8T1thkq
XO5dZWlquZxTQv5oVbYmmrhNPGb6jyhWugLJcXK3Yupgy0zYSAvqtSSTxC8LuXAN
EXUohX0ofKIQVkdM9PV1+DyCZw8eEgG8Eh4dtqS7qMc7ZvT9fr0KlYqfGY1KlamT
9aYv2Ackq0LjOK/TF2RhZ/mQJMn77o03EZz5af24ycA3WEt7+/ZtaWJ5tP7sbw7j
J/m6k3ZsYDib1vF76Hew/wSBXHJuyNYVc3efpzs6/R8sRSbyOtj2kakP3y5ZD9zx
3CaxGCtmUNmgeKPPONv9s/NhhUEo918eRqNiKpPoZr7MOSdWg3ls6NvaGRdCx+dc
VYzasxja05OgJxGq+z+oIgUVidywbTQDhgSqH2/KE3jPRTLNE6SYhJsG/PhwIE3C
PsLOYim6O55+byYWJM0phdMD4h4O/H6TSlRMlfuyDyhyTRQl2+lrHdd0jr1E+jrv
CoZt860nLBlwEPOzCTwGP9AwJtuxCS97fsmfiCld0hubSGk3QU9lpIk3D1ujHVXq
S0dXYUhovuSpNH7FUZ4wxUkwCXTOtoeO3ezyC4JrEllh5zsUYPN9+cjg3wtTWY3f
CZTNRhkvglkDdYhr8fe3ysS5grCg4BFhZJXkVBXbJJef7isRjVyy4P1NvE3VjBu1
mdKxOwV7u/nUIqVP8e1tTm7kAwwADv3+s8bfQHoUIUicGFNkTP2FC1ATCcinTPAc
nP4WjiP0HML5LbAvnJ9UGlzFPytjOqqT9sSrCdgfTDjaPHln3tnVLrkf4xaeRSM0
wcKwuNluZ/xG/Wi+6d9mdmb16ELvD8qmcGazmyEGs/m9TNJmbONuhaHDujfhPEPc
fdwrjr/woB6Hd9j214JXxilMpPZA2wN8sC8G3fFpHumKqurYvlBv7qclA02FBvwf
+l6jgRF46HYobt1Y+6nOr8uUoIZJ03WjmGtdPkhdJCXRVOCLkrxOswnJLcsvyiUP
EbltdEnmZs6nwdKMchxM41Q13uTjvE1zpM6TtkmbIBGWUAbHJ3eXBNDT5uzZ1Jr+
qAB0N0vp9cZGemnu5H2tcDnvHusk7hC0oxBJqnhDO65VXZnftUtVcib6BhlwlYny
cZ+xH8/GsWAtHFGjmmuEyyJzjg9I2mUXyYY2wbqao9xaQk1b7ui0Ex36vx6pum9q
gb1y9R33zTCW7bliJpkVMebicG0UjoO+//+EGHLbCGMnBQHUYGrXz0VrCwdEwncj
dhUrYrCb7hb4MQ6Uv9ejMbUizC5byo5l+4E42Y5i+fcPrvocuHi6KNPlzzXYV9vt
kBJBYJToHSdoEKCtXoq1XTWw+eG98JRK30StBbftv8UksQPj0LoSXOi2TJLAIWKA
UTEr9ZUluM7ZpDlTqCbd4Zt+HAkE37veOLcxwzCuCJSDNxRZz4KvAmJyZmYWBtTZ
oRnMWc+77Sa8J2zBHnwH3UzbnjmCpbY0NifsaYQ27AlxnEQ/+ayU+rbrM0+X6Sux
w5l7F2P2gazXAEPzJ9wasJ4V+SSzw+jPaC5WaES+zhS4jsSemU2nanp+d1Em4zR7
f+O4ZQHGYykLuneK/P9pvzbvu79IgwqomZVf0Py/763j67kMQVsdwL4Ya7u8K+YY
E/v8RtLFZumuMJa/8FqfQ38s7l3BoquTOoSPKL6Gs2yjwH5FgvlmeGm75Uru3A0f
KJq5bMb9XyPIAbl7eulqrCZHb48JKQ2O6eMUcCpnRPDsqk0sM0k/750w7Jzv3Qra
2Ly+Vuqp8d+uYv8VlmHRbpB0hnnUKTG37bjcCTA0KngGv76pAvQ5TZl7SAIbOA2e
mln1luXYlFdpHqO/pT/ki2Oq8t+peCftaAMGWYxVqX/DnjzUXIZDQs6JjWGzSFwC
mfYX3S8aVT5/y/yVYyzgE1Qf5bayZTDud9CDtIX0mMmXdzaCqVRHGVFQn/51POQ2
tWDC/jW7s3EH4+acebg00m2zzfj0XkTPbTb0kuJpj4QnveR4vmeCSD9TOGn8VFPQ
cKJVlqu+khJgK3o3v2ATb3E2U35nUISl1+DzDDYmiSpQhqGB1YqoMvs2hSLoeOQo
Nga4HvRjRL928ytSh5dEtuPDIr5cUfqGxIVJfXA6S1VeS+LfVQmOiV0TAs/AdoPI
VE1+BLN2nLh5HxzfCZnaiB6piMMnHYC49Zplk7YXjHslT16P2fu/yZxRKZE1efmf
GbUeiTeHlbTm6WP2ylgTnfTJMnRoojlbD8vedPsOQWHIaWzgQnY9uc2Cb3IyACK+
mNAppT3MsJnFyqzG+va+py9BHNARmacKuNL3CW1H/OanrCjnjj8W5RsYsfT6j6px
TqhQWiSlixXZzq2HGEo7N+JFPB7G47bfc88dy624evxIN9lpHwWmBw308uWEM1qL
HBY+pK7RZOdsJqJizqMRTMjcjsOLCLaInCKCTDwXdYrFUtZhWatOWJ3W+ZWRrMS0
13kcnjpH1PzzmfTL9tHmF83vIrKwggVEpMot2F/EDYChEdKCP7Wg0TaM26BAn+ZI
ZGFR+1MoMnOx/iUiHo2La/OdrO6sb+TyTv9InNSZQB3TkLkH9FQqrpFgJ6nfC1Je
w43I5brkUqVy4In8e62ME+evRCqjojXuPf6S0emt27WR26Wc2GnSGsgcADeyp9Eh
OCeZ8336gM9kvr8cf1VMvzOvBn0wqHzcXKxo9YGUbf3zy+2hWAsn5Mo0bKy9c2+8
Uln4gMaFbAFWaCbRra5+7GukaSalesk7UGJvNR9CFzWv7RWef1iu+YUTWlWDtnA9
+5a22zETB4Fzl5PYxjESPBBf8rvkV6w6QQ5ACA77P0iIr76t3YXCQ6P6g+L5ihuS
k51FAORoS7OPMwCNZ4j4eBoMiqV8u0kusGHZaEz5T7L1BeWqk/FgbfJ81AL6dtwk
ncUob8cWGiXE6T5hEkc1c13cxv3ZdcXhoySEkWu6NG77l6oetfuP+3zciQVoP5GH
odc2zusDrQRVk+kHE69XfW0um1gJgOU5u3+UH93C7DZ/LLmi2pgQW0rlKerfldXS
u/aIasMomwvIBwVslf60k87eDcMFK51RQbxQMWHC0MhnADUGXiru8g6WtNkPpXbi
DJhFTinwsNXyPyoTL4g4wSZ51JC6TpP9m+lDKKgP6XkWe/Khi6Ase54Mzqj6t5PP
pROTQng+fC2nD3AZkqx46jzEqTAZFCVjeHXJUjDpxrPexHiBZ2o2T3D/plRZb+ZU
i4R223I20CRIm0Ar2cpM4kLOiI2hae3p91o0gOjHQ6FhnNhv4sK5TLEghK8jAcC9
9sGIRyIF807NynKrC4XCbKO8UOVJvnCS0v6D+930GCP7/0O7Q1w1hMnHNyvnhOAw
JrFQrNxFA+9ZPzOdPeAh/f8DAXTUKqgYktg2QK2v4pRcBeL6IrTgY3ZnmgDrS/zl
ssudEo8J1QtZ4D67mNwDnFIZesObix8tfd9Dce6JudAsorFhh+pCYXzI8IQLpE5i
p+miU6hbZSzLygtlH9dOoAmtpk0ezbd444skf2HWsl8hZc4AYBv+oEUmlSsQWVwq
px96cjcy9EwVegdcKiwXuczORogZM8z/7//7nHsOdEqOVZRf5BWwVMkLKC2Vr6cz
Qz0NCf3kPleCNUCl6ZT9OErN8IHXmYwmNZo81uLYMQK5kNEW4D5WMrMsWzGsZ6af
JWouy3Nur1D+byA/uYM7NYuoXhndmoJ6voH+BSxLm0F0Ma6ZBhhxw2Pqk/n5u0e/
fvEwOVgJu4Ski2nGvklui2KIXqTeXCUSl9Et1X3vrOidoBplUhanuhdgfbaxwaV5
+YZOzLD1wO/L/4vK7jcftmjVfCqnO9Jr86jrVURmfntuhwu3f5DZ/VClg6kqRGci
XpgsbcLqQL6WWPTePuxdeF5GZHMfKeQOm7+zBDuw7YSuAJYHY6T8wFLdiOvhuE35
jL/W1neuhcsxH7iLxKRbZFPQD/FnTdwOMeAPgcPmpEZBgBPG2Hl5AaBwH0m8WhhA
vjWkNxGY+D85Zs4yMdWSW4NKS66i4Orsjgao65EIPw5tyE7MAqacbHt+XQyBYC59
IZG+LQhyEmEigvGySdvKZpX59mU9+PUN9uUZTsn+9dKLhoilqBzg818DOiNynr4i
HGw1hn6N3StBYYveFF6pVLabL9YoJOjMWbFccvzZ22cBntW+m/SF+bNHLUhLteSq
ZMw4cTjzQyIgoQ8hltNF9+gbbBCcP2EgonU+WVf+Z7yPWazpnH/zXRdG6ay3ijOq
VMTq1YFqL4oRmZ6BZ0zUeXnBxJHz/u+KeyDdE5V8BNwnEqa3OHUadsoS5yacRtgK
JQN59Hd5xhENLU9tKvviOnZRQ2f3ImKCWzhaSvJXMK1/q1X7UxMRDPQzZp3NzPo0
PMP/rVZEq4zTyh6ie/YukvHMNoE8/nARSqsl93Femobzp4hVK8c5dCPcoHvvOrFq
9/FKTiuvh1OD4fSRSs1UzQO3MrCdmRnAtW7dVijDpDFbpBIB824H3aRQWlu9ucwF
V6WZaxLo1PclZ4TngSnf8CmEQtXiK7INl0DOw9YPsohAXTtxt0guPl08LL6ymP1T
eOiBwxrnQsfHjbNvMcfrsYnUNP2wrCCevcd72SRP8CRN4c4f5XdQHn8sKOTkFwNv
JQ1xE0h/zMe8EcBngwR2rehiUCD8mF5oTg7+taKu5fSkOnk6YsAd84X2ICeJFpGZ
al7gDcTJVkpS6YN51hxPYce4Z3Kh5nHSP+6ZBtq872gS/kfxG/oRnMlIkZ7EfvPd
ZZ4X7NRpgr/to+0VbQlPiWhT3RSlr26Qw+zOGYjxkfu8hdTEdU+Wdxm/nDw82dWT
lcci9GazueoFGnC4EWSuGYy5P3Yu95Ne0VKdqSpGwRLLK5CpO+xbPY31C493Zski
UAXw3nSByWMYa1LGHsiVofLR6lk/We01C/kppfxvXdH6bRSlyQxZJuTfnNEXSPiU
UJdHF7oTpuPlwWGysGLasqOg3VdTLs4pfaK5nOXUIbUVaue5UI1OYO1ltOSOIVFg
UlK7cbVv+5qvta4QMGXcl9LBx8xHYJhTxCGF9CxNxHg2WFluEFGS7BXTmsFfRZj1
eKjVtpDRwenUBgFewAGimBjWz8x/R/K8ycp0lZDh55Qj4GAjOsmJpi5pgSZC+sE+
ZsIDJQ4Hk57Y8pk03al4Ah+qgNHmqghc0pBrQQ3jUP7jYxq9l05J8LXRqRvt6Slx
BBjJIfEaNxrj/zKwruiWAwsarVci3Q9g/Q0bG5M20bs9ciIm/G9YV27dsjLjUuzt
sWBD63NU4+PEQNXtI8c343kZNTOTPy8nYBd+7eL/0v/cNM1ls/bHviNpiTWv9brA
q0aLPtqpCZCdIYy4PTSTq18p24PAg9XD0kJ/iIRTMRJY8rAD420wjvpH6txCLJ7H
t8tIz5s51a29puTFuYSe3oW/89uP7fvtqZGL5kHNQiw2PIyU7H2BiieIVNqKXD4e
ZeURVuu8hzxwTk9RJUSBprS8gh8D0JRiVFuyZbcTRFE2W06UEYjuQF2GFIWL4m5k
vN8X9RMEKk/DQQPpObHC6fxWgWfNdv5/Ft0mTlCyHKTK2SSa0m+dO+vbPTIy+tCd
g6zUc2CQ/c4IoOy3QFfOrgCC0jxRm5JR2z0qewB6asRsCsP6qbOs+Zbv2xMBcqBU
2DQM6PdYWWcCCZ6ZI/T/QgUc/QcToxuPH0GvWUBlF6Tn4PPdYymIjGdvY2Zie7Tp
S+BgCMEC8zR5D8CAQf+Rwfsv2iEJLs6Fpht9Utly07+mQTSXhcTJayRnPv44Kv/R
OEwe3CiHKGSq51h/oCkt8qjDmwRPfcReBR2kx6n9DFzsrMpVviiJynNKRS+9AvBx
dRrtfhfZ4XGjoC4A/MCyCrtiCd1RsNUWRAmaCErnUu5Sm9bwcIRxfhf9e336Nuam
SyVmWudzQYzmkslJ1fW2urNSlJjne+6lopxhPV/A8/HGQpAhiVBy30huZhqe290I
XIgZxTlyGhp/GQ6DuYgWmhz5Lcp8xriQK8l118CLsqnYOCniw+JHP0sXXZpT19jd
gA4STcj3XUDqtin9kjPyGrROBkUmfCs3ROzZjx5Q6qp0R9Yu5m7nmf/ANKCwPSkk
NuRNQsTONv/vPdG/m0+w46rXJzJFRAJqm8Ev/I2rUJK/1waEp7Q6WnyJRuaDM0Wz
y4OE0Hk9EypRB/+fHKb4vcyNJ1AqbAdT+X3pAlEm/CO6Lx/LaYg40+n5ArnH3x/Z
NY4mqrOUki+1KjfG8aAa1OVCZy+3f6OUNUBbJ6I/orxvOBDp0N0ytF/jjFL//gIR
NK/+ws0Xu3pJiJPFRwLWwXF3MZhPQ9X01K3BHwV0oHX2AbJawOVtQFVY16fgGdzZ
QMWWY29b5Yndl5ZtfwSmvkV6uhssYOQ6AbcTjfbkMA3r6AttdvyNPuOUkyTyqZMK
n83dstL3pD4cBWhK0zcKrJQ24bFNM1B8XmUJlCUtSJA46AZxFSqtmopLvv8JATEN
jaQPN7MgVewAmJ6tZ7+mAf1CzCwnt4ePvRqYtHc0MIUAwmLPsH42so2fhKPUE5C9
Z3Ghskds9GVJnX0c611xjOxIUpsTl3l5umUUvhZ3VIJhRF3S/jcyrnBUwYcOUr9H
4fCBoiDPMh4br1wDlMUUz3FMxHo+2czDVORCbY9sPkHVyYICyIAD8O3xEW4+U90O
ZnQi1NZ8zSlTF2t4oWpRseG84AVcEboNhwdKaWNhPN/VDjcTctaOJpbPQn46jCyE
uSs/isltTCRIv1B7uEgkCFKHTEH8q3YqFdYHPPGFVDkZZs+e/SkbG1y5sgyn9o5m
TCy5C0Kd18thVAZMpxkBsYGpR9GIGG6+xoiULmBIjyFjfqH8iE7rknQ3glWtbUCA
uUgi1P2Q8qVgDg6n+bTrPRFEsjncuFu/trBtBOjlY/XYzxORkvAkZIq4533YUXk0
qOakYECHD5livjuF51o/8b2wvlY4ZBSxbkxalKO+E+sDZ41iokarA6VwUF3zmYLt
USzxMkO2FK2uqQTpn1NsRSmbmYtkyWt4SlNYzXG3RlyKEsFoRCjTJIKyw20dw8do
2NcL7zSxjQNrIHdVBzk4iNqEq4JpjvnL463sQ0PxuF6z0ZbW0/OcVhm4CyYSaG8S
k5K3Z1ch7uP5r79ZYn71s8mRw4XKVfmrHrQEFbdut4frJcwYR/VE5qu/lo5X6vAm
voOhiJHqC7pF/1IAMVfu+uUFMx2Xl47kwPttYhYBZ6QVGNZyuzdaqM14lTTLDXHV
IlUt7VZY44w8awh6epCnW4nhI3HAeo2/bfIk4+MbO8ojO7qvealPMstfxrMiatBJ
x3DENQWZzUXgNw4zVgPc/sFJKqJgbBDXwcEiQfTALw4zB2XtzqjJNupJoSSEcuG/
WlGCp7tLFxUC7NDLbVrwucsoYZfvyzF5CTavaTm4tdx9chzx3UGGHcaBFS/j6HeO
sAN0kk16G2wrbfSMu4a2Al+3D1IbdfKkZD2Go2LkRguxFqUm+VSXKc40l6PuiFRY
nAFLAJ7d2aJrOxRvzfnOcZ4Khkko2ltIS8+XS4ZbG9hbukB+JFM9qbCoRiOUWz4v
k4QAIdSpUwdfxVLe52ntoeLneM7LOX2O9D3z3orXRuT+wbJQckEGu4ATmm3HXsLr
HNvYX38rO72c6irkYIV/1gHmS8JQmybJmAO4f2E1XuUX2Ua29h7tkDwQC3FHRnDB
0tUjy6EwShkZ1gRHUSVtaxyEMFZvwjooUR+Lrghl9Ofn5V0XZfdd5CpSWDcGJkDG
bhU5BgxkcI9MEaG7L4le6nrm7FNVkNEhrky0EB2DMn0eDXEiUfxe1B/IzaWOGlKZ
+BEMbk45YtNQLUV7Vll8DjE/MOnSPyy0cv++3iGvCu/TnyOn80O76EdoGiW+fsGi
KfWWJR27tFRxUAnIyo+/R981z8OWrVHy9AhX/sTK/TJPTOPniPOkZ337STTO7kaJ
e4NGrmIDZZcC4hDSTKjZrZIvZW7QfwG20Anmu/fVST/y1M4zKl0DF9mtk42Fsu5K
FREJjMeCxE3dusofGFTIJHZJVjhGDtiSYu0i7Yc0qtNi3fH4a/ypJ3Bdrt5F5jFG
MPrZ9cnde/wq2dppsGCQn0zrdMe8jRtOFZfCs0zltRiyjhJS79z1Ul90bhPckKB8
303qTXn/s3/RrKJD0OqecMAWsTObsGA0hIBm3C2E4kp+b4nmWpMhGCwRKds6eorv
/nu44RE/2Xi2dM62LZt2bNkGp8V7w3EA+t74twqGrog4S1PD7/hfz65fqCCM6hB6
4V+3KhBa64pZpYaFLGGU2CpGTGaduMdwv9PwUAZRAVQOx6higV/EBF/yoxJJwsEa
OF8UjWGB3mu+Hn/Z/i+rvWuGsSfJFRsb0zYxE5EwzsyFq4p2em0rkMuPgChlNE5h
/BQsV+sim+tC7yx40/NrmuvUuhdFWCjG9rEZ8MCFoCKE1F3RBg4h32oT6cafN3+g
msvP4hp5zH1aZr0OoUlMI6ydPHshCY+c3opvTcD5YsKYovFHVO74V8yGUDM44xPx
d1UIbgk72BSY+oe+Hsu8DnExnId/xbhXNUJTEibgIyDA1s63OVA4LjrmPnWHcHaQ
+K5G8Dl3OpJVcOEls63Cu4NvaiwL4DN4hJHVBMv6Wb3MbF995AnnmhRTZG4Bj9o/
TgHu4zJHJfeFC5jc+NSnQdbQGaUv8E7zN8jBLudo/GNO9pICMn2bA6JpKbtQog1k
CkliO+LLbfL/EgJpyX9bNkNv1/Glq4NhjIaqBJKz7NxaQCFs9HSLIfKqrgc8HRNG
z94S7Uyjs3SyHpyfHwzMd7hulSTSgmSDmqr4bLbLFCsABsbJNBlGMtafMZ4Vw5yO
dlJkiP+kh8ZArAOx8CFxySsU616wpN+AfmCRttD5oUVSBX4up1B0XAhP71aaWbKr
3fhVNu8O/Tw4SVlURmP5F56BFGxsEnf3mY9TohfJzePEevraY3F0n7mNoMgSAALd
pWgYnlfkp7ER0Bx/67tCIsUHsXf6hWlKkrKW8GE8/3fLYFzWg6FEv/Ajn3tZ4I3H
KmzpunVFFdaoEKJSF+FWLU75k+0B0me/AWZKT/84MXTROyo6X206Y6xNhuviZRwm
3HWl3chtulQRxu+q7ndnHGN7KCc98bKO4Hi+6MYcRciDmcLY4UbJ0S5XucLUU5bb
iQVFrh1GQrlJojgTImd7Mb4Z6mgedbQ6eglTGznz2bfS+j878DN1FXUXSwZq2N1x
gKaVaw41zkiRSYZSOTWW+R6hFMPKcsjyvhSODOdWcNi6IfA8QavK+XxFyVUNg63o
27V6Vfbwx90+ICpqwb2WTDpyM3+ZqVLRHImB0OtjaYnRj8Y4EMeenPhPyIwtvSYv
hVrO/c86tKAkyfvx58MTvRWLuKqQTzGUVoiGLWKXFBg+RTBHVX82t8y4x7/roXCM
eP+Z5tQ33YFEkba2rz7JgvaWubTJNc5zW6Kwl3TR6fNv8HFEoYHpSXjLmWTHkCD9
Ms2UnlkfwPc1FNrSiKvnGleTUzucx3V04NnIWnCoBfDZRZLIVtH9NhJS+KPCmVOz
Uo0xRLXq5mXt4xdXW1KC5i7qKIFM3JOJyEYlRVMp8YofFmet2PmQc6nDqTa03tOY
RYFVMwx0iqtoAOdt8xv+vdUDDd1UhhQSDbdIkht7Gjo0MMS7aemtMh7QvPgDxm4U
QHAxIU29pUQZU51RYEn+3j5KKH0iU0/Wb4b7Eaz25VQRTwvUSjvEKKcxSb4zyuwj
JarGK6m4/NSnpTCr1s5vd9P0mmVjfF2C/YFiMrOow1bMCcS5UQOODODrue0eZpHK
KPVT4H0oYThPObMHubEztoQK9S4uLP1ngWQJLtnswqJXcPjHIrT0AWEQBGkP5nrf
HP4jLJOYNQuj20Fb5XNYr1JY3yzOs7q5fzL1Cxn2cqsgOdUKxUn8TWbSpzySZ+Uh
s3xl8trDx2xgIZZyEEkzfoT9FXGrR2q1Xbv2yweUODMajCqXNQE+4v/3JekjbPhJ
PA2Tv6/Xd5nO0gqnEa/rKw4evxMB30lY6AuKv0gFKw81SuPNRdcMXEdF4UAOqCcc
hQ+Y/KMbNxU8qIyhtuQ0nA2D8jx0JcpUHGGHb8dQi+hoYJxNIWvBNULuRS3dzsrV
0Xo3OyRbvkCye7yPtuGcnjg4xNu8k+2fsM/+oANZzCJ0HnKFWPr+qBXhatmoLX7w
hbcDRQKUGpt/VQGXn/RHf+6ELPRBNFdMY7BQFnyi9PqlH8RE03yIIgUmlz/1jxSb
Mothc3QZjDFR3VwSciFfYd4255U3fdsjOdI537OOEYFbEwFWa2DOhdQTYaIuX4dH
DoQGzxsnH34sUq2KL0imghmfGYNzF+mjtYu71AWv0Lh/WQDbmLfWU4Qrh4+plUVf
iQ/Q1dugEh/i+GWNtoK5c9I+r/Ce/mAMoTMTuGROdD+Gs7I1RNkUgC9GEOCYs7yb
6aW0iD2mXRbwkEyWIjc/EVrIuE0RHNjufV3jwDU9YLGuHIVAnTgB84AIllUPtYSu
cbARVl+QGMSuTD0COdLeoTaUdmXMllLC73a6a18aSssy7opT4ViqCnpvdUWpoSI4
nlnlPZib5bKYNjjFiPgZFBCumLnxOqNc0/sBb4lQObboOTCn4Hlkbnc0YCNeT5YT
I4yWghKFVH1sdFMRzb4J2svWPeeoQS9MJdhGOzySPNsrPWlW289ZVB6eP4nySerj
C5/Oz39RyRchUqGUL4j2z9GyXIdzEhcVjDGllvcChllVeIQBYj7UqcRWWj4MvNSj
txA1eBEWaXZeiD7wC5ir7MBUQi9L+fpfZS1qy02DXrTYU/mulmkaAjnRb7arkIhM
vhrVxDH5TFwiK2NZDHmy9MBUWrArYApVyJByaPbPirZfQ4ZA6kWPQsW4l0IKU3Ra
NdRxuLSlpQr9CZj7oPYXm1ZS+R3BtwgmPvjkbJryRazJk/fPwv9KRL73gBy2vOl8
syvPr2bciTMveGnrb2cROqIdFsOCPTPLwFDaaETjq5pPOxE+pVFYfiVqQb8BRf+W
7/Qv++Uyi43jZSHCWXC1rgTx6eJzCa9Y8Ryo1kIYvp9nQyX/3cB+JnwIU8sL5FvJ
lKjxCuGt5NSN6MKaz/maF59rRLqViUqa5609XtGRQsLxiPur9S//o+A9aURXpYnw
N3FA5syjJowc4/jkQgqDvO2B8O9pwL3oMnRuGMI+d4JYIprFbNEeGI4WmBBhnY5m
CHe6utNqieyMC9wHIAJjrKGH9E5Gk6NZGHaRpeQfMNqSZj1O2para1eOMZE91PlH
zJIQuEgX+hvmt7CmltAw8wob9IA1Af+kBX4O04x3lpCfylP1LjmsltdHOwCTpONW
lLKYOwBWN7/Xl/t0hhz0aWZW9h/l3WkApEPnAfG8mO/pFfQww/+ShR99QPJH+geW
0rJqshjI6gC3z3Zm/2CxQKBV4/O9SS7YT/c5UXCGiZTwKjBBVUjQanyOFpbSgnKr
EtfvjGSStiK9cF2OXc5pxIZsjVG4JGsyZ3z9TTsjht8AKYI9VRywn6/8EovJbHbF
wX/IvRnkSYoB0zVtI/GJcyWWrEyE2zalhrO+6wvvkoUPVIaaobC/JbKRxa3zafYU
LkmGUAtu3VVPoBMbn2h8zR8DhgSG8NWBqa9/Y1pQFZ1mimDuCyoWdaJ/TC+FQFJh
fQXJwg84xV48Kp09FmT1wcUDcXcFAM1GqLHdcT2XuVdFoejRmFqNTKgXLz4MN6YJ
zVZ7kWI9xjNAawTP2nosYQiOLvhROn5ifebbcgNXeQflZPmd8OMrrsFz9KZsYdrZ
QAlb5z6rq772C+W+NkhDTiaeaAVbcJN4IKRWmrmILSgg6E0tjKexPyoX9xL9lhqd
fYfrIs5SGIeRfZY+lS7udGVyqLpKEhRyZiYEUq5EsE3XDDpHF67RjHlU8WyNFfYZ
ZWTpwLwOMxSKdv/sISTkaDmxxG38AkaIMsl582h7bPr/FnF5DBPBbmTb9Qhy8Xbc
LH348a8sBoz5ouLx5WIIcd/pWwBsuHtpWJDvc0mAJgzGBydO9m4h9WGNFRt1XUVE
BZjekr+76yB9Pk14UiWEprGlnbWbrluMw/OA3uDocsIKwLyzI3Nn6LZdzxyka/LH
K5NgnqJi5dK+mrLUeNZvYef3ubS5U4e/wzMdlMilqk1E5OJpbZ9X9dpUIco3DRVT
oC8CqMboTDYScOMy1pzD7+ijfBirTwvJ9fQS7nN8dncUVd/hytEzwZ66ntX7CjL2
rGSnNu1JYFQBuEifh9O87GMfPsVLlOyINyxVPK4OKF7IKWKsSUvOJXyHuiW9rC91
M0ANLhFog4TrBAtoP1ZpeA5IopBEpi3itWUearUYRuWECZGfFBBToo6iQsgh/9Vc
gijhnu5zkQZuViAp0F5CQEM/Aa70YPy05pvk8pKi6GJTUswedvIPgTizt0cwV3Bi
z9X68y6mV6SwizjhXnm8K0yHz4U8/oyiTGuBpFKSnfEGRpbTGAyTK/zKbXxapCwF
ik2zI18AqMrEBOreowqjqpjW3zOKzhIB3SXeLOkp1pW33bOKfHBnTD5Gqhyo4G9s
SiJV3TUK6XPFFA7+VZV8bzVsJlajCibb1hJbBnRUZi2g9q+fyDGdiv+IG7AoGfrX
q5QTI4JugS3/CSjgO15EjB0QWblpobEj+rCSoTb8oxOtMz9H4KejcAiQy6tZmSny
QxtmgHerJGKFhe8e3/4qIbC4rqoWTVuEIs85mbTjANrnUhTj1MB8YWlcpSf/QuTL
24H/PoWaQGbDuUu91qjh0JKGvfjy7i9EcYJQ/spnmPMISYtR3JF4CyprSnUQzBYU
2PMpK9Azmzoctp+ZgRgSWjz83okVJBOgyasCOTIOSrcdg/jE7c3SogVP9m8r5JQD
+KawEeDswUHXZXMfDW6PQ+flAsMMlr7135moICqPgQ1xXBtexR06hLEn8nd0ICTG
P6etVEVq2Qfkh9MTZdudhULuvtwb+O3hjOiSRHhJtkGeAt6ugZ85XvhkAzbTXjFn
jgUmM7VOGMjE53d6KjlXp7pUMvgoaiAbG2Vxemc/vP6IOfJDF8chZUXptA+XktVV
6wdYC2vRuPj6nEixidKyQNqR7+P+hEP/NVXHf86aVBnDGhgbW5fKzceOAwfLW9Nm
wIN6/qhZQIK7Yoa5Mnhk9dJ5SytLe0IWNncBBS3MFuQeNfTGpI3pIRTtKkIcoQuh
i9bkRK2w1JynDQGsIS53kBQ37oG0TvUbui3goXP2uj5ziPkPyUzDxM1iUvuzyTz5
Jmyc8tdjbl5ttpimD+6Q5ubfnwbyskFYDx7HO7wlI8o3I1yjuE1/4H8dVdqJbubs
FFMEDjsYz8LYYhRoBgsQFKA1u2B+/BeqT24OQMuN2mLw/bQm6FC3q+4A/h/qYHSl
X23wvzBh9yqcMc4tqN8CadzIugMMyR2MnPJ310imj3LsE3rqBHBw8/o8nNXQLKdh
mtYrkqRtGbZnol6ERO9eTTkZNTSV1D+q7cA7amYmxs6xWRxj/pdhY4K0pIl88Csi
zdyy/vWS/nTRB6SAeVLtVPVLhrcEv+zytK0vGwSuCgpfYHDQPCIB3bblE9HVKf1J
QU3wlMPj1QvIdoQWlXGff57KWt9vKyNr59VTrTOK7jGlktuHVrOL12hk0sOOIzgY
JkrafSCZWOJGXve3v8wHUFftt8WrUVwN63+44oEAN1laat8HbkQZwnLO/ZVyrHLp
yEeftDCoV/RqneGgbylkWK1C3aUHOyXTNkCiga69Ox3pQsF/wwJYjXd+OSwNyRY9
ARqjnIKETwbW3oRE7QRNmY0JDrSaI2PRV81xXyr6yDwxl2nhFdIYFkLFERPLTL95
llbIHOFP/YTbvgL3I2w9sZZ58p13H2RfDpYCU5kVhLidEIUus+qC4OGnrpk1pV+d
sOJw/eMnTV8ldRh6JcvPq10J6teaWcH9F4VyBoMqHWrWkizYhHIqlibsjjd+o3OT
I2Izvmr7U8P7DvwvUstM0D+sM6Wz/nKp9VvCv1mr3JML6qcb2NY6MOWMFPW9Saom
jJ/e5D6NJiH4cVO0g8x2JqYFd9Qm9OOTIp3DnXEArRJfpZnUVYI3fimF2rj7Tecs
IoK43gtmIyEgdT4PEXJThp9JMLoEAYLjEv4xbVgvN6wU2p1gxJecMZStMJC4k4yj
SQofVi5dJyutjjCzss8ifgMNKD2UDADEmDraPopMbP5MO+ojK7jiX01T2Uis+w6w
HVH3oliT6lEiN68ucthGRuTm+dgLqLVsEaclrYlhzbDMrx9X24Ajzm0Q8mjoeUWn
icglsbErZobPG3YYBC096cyKseo9TFCN2cfp48zl61BuzFsUdCiNccXYlwFslcub
64aMvX/qAK+NDs6N5799SLBcnWDAwAtCRfboqPWg24tjoa/WqmC0Z629icm+SoSZ
Y5fDO353vRq4l7AgTxqBb2BcqotCIWiN0AQdA8nxJKIzR9Pc9+D8SBOWBf9aE8Xz
5zwbKiKvevEK2hROxtdVduj1FUJ0x2WBWETKfRY4WlLf/BF9yLU4u0V/r1tuIgHd
XJGTsBtdqXDHNYvGcWrPgeAqDxo8PeuEsbWtEZKHXaISFs5Rn6LMv4My1asKrRMg
RQvLEBGtwSqx9uFGtEwYXUKEhjEZy/8SX/+T+qPvg2A3kYtZGgOk707a1G91+b3k
XIWBII4SaUSTx95J1WUvyZURWNDvn+Vx2eSR+qSgBTiskt0MYEd0OKa+V0wcbbC8
OS27YNiEmivnId/iG0wmWSmIrO0lsVnbhJct8cZ3w4N2Nv3RqkZcXyzrQhGFLTLH
v2e26UXexUAOZt5zoAHxEYVuVA7I1CpKsIUIl/Xijsq+a/Kqbky0/641/MYXtTRQ
eQpwFPY6kvzwKHqXGZlRsZ5YzxLKcVk/Rr9cuJ5L1pbC4xu7XqZP78uPL65syL1d
64u6hbNZKumiv7WSdNM+kZafHRp0/RHgPgqnbFISqM/tzDuerF4XX+rpPfOtVSVM
ph6fA2OIW091aBfFhN8zIdljgsX3V6Us72ElfT8CLD62n7os/eYzcWZHWsDouf7z
J+qsyxJgh9UwUE4CjzGFXt6ly7y7dfDLiy35j7wOB14b4OBQswkokvtccobVViWR
JUiB+xyy0lNk6UXfkErTxd3BG5w6a3W+chaPZPB7+sSibQQForYluShyfFWUyvct
A3IwWmPWZcDucet+p2sVpTGG4AgZZ9bDRPAh9gkNfb71zNvBQC2mG2bABuqCrSKY
n/UEexhb8cJEY6x7+3/mWlknWKGXXnQ2CD5bJhWvF1v5ir+KA76PBX+VEui9a8Pz
OECKudlwz+3qIKNvsLg6ZfA/hkO2X5iwsNSXRSXbT3EB8VJ6Y77Qj99jelhWSQkC
mW4U2W9DYf3r1sTYUoVkrVbpXbPqeKi83MxMIFPG0wLa2PC2PF5LHTdzM8HPduVB
5lDC/MzxpiATBp0A7sh+BSPI7Qn9zxueuwEPuaO8g1UlLhltBrLBI1rDI56jr5YS
/huX1I1LjMVIKZLX4E2Gk0E40LfgUt1OIqipOd17Ep57pqXyOifiEuMXZF9dHMuj
mlA8GXFClo3IiDVs/tJ0eKbVsoG3cM0l6n5s4GnZAupn4xqrD13zHNqbRwOUWcWb
tj9EYnSmuNF1HkJlsAZ3AkTlyxl/Yd0M8xUdS+FWOSwq/oUHkYERugQkroFE24fe
ZQgPSiNTxs7fjSiM+aGTvqtvwWSluF+pZklGLkio5VUfh6CtYlJXUFce6aSygvM5
GUubcu+N7FZOF36rc3KSen3dq1ECxAH0vFa6YJxeZQWrwiWVSCy9Gfnm9bmN7JN9
xp32lKfmxUwtxlRHwBimEOLzBsgp8FWFB/zd/Ky0XAj01NGwe1wW05Fs8qGJHDLx
DzgkLdFUhhgIBM8RFsrnq08dT5DwCOG3ziuyE69jV++8rjI069IynhaRU+oEbb1t
Cp65xfRdrJAT7dNezUNQ+18//1n5O6yVIoVBLGhcgMYWD7/Eq/rCFEZZOUjC5tH6
jYYJLfoYvW2Q4Bi5C/tex1wnyyBj04aB6+FAxqttu2pmLVWVrojoC/XiGH0jrmpz
nvj66e8+TFUl3d8uUPGx2ASWBbwhshKg/WvdEF5ljaANlBJejJXSeuTatcBd9KDR
T307QKukJ5VGiOClHOBhfSPt5I6fJJX72k6X36XueehN8k+X9JeaxPE9ZFgHRRN0
DzE8deNyRSUNFwClk8D1HYysP/LbNlPhOMfWIj3LMoTbsWIGzNK0ep72Acz8vvQh
6fb7+rUkgE5JJ/JSarvU/TPS/I0oQrwNZnAcOA6vEw5xeAz+WnJaGufrP7amh8V/
XlLHYmtMyo8Neh5RuxWHAdXaK96E9A84TppChNgLQLwZfUhU8GonSwRS6y6tEG5D
lc4KR02MbiPIJMieoPbtT2Fr0R+G0/Zms6aJus5xaa0bC2wk81jI2YNS7AgNjrPH
Xcu3/gZ0zX4QZs224yMbnLd5r/oszgQKiM9kfZAiy9twg7iSjN+kjsMOi+hqjCh1
y6a3OxInMroJe1YZ7clUbtz9W4+obRGeB8WTAwP06zI2aR6vNZx1CfusM/eXpt5p
rw+o3gGa5wQNHOf/zIsSELFjrF+t6IlBl/KvJGQ6G2p6eyS/ITCREyhswqsKVuPA
GkFGY92rMAGPvTTOTbT6sNhyUUwzncplTXVPt26PoHZfBWp4YT+eLcCJvPK2H1hf
ozZFnTT+ZbGPQl6q2+l11cZ9WGVo7jtH/ZQQOYZO9oJ8NFun3CjCYihJd7zO/yuC
Q6SYRE53Tc9dFyQ4ftfn9ufS84Pvc8psD2aLMBw43DiEUcLFNspOYkmPzrUKgvVs
X1iBHNW+C4jnTBh3NfJZldcYfFXuWbXdTbxWn1efMJZb9BQ+P7bgCMp8m7ajFh9t
3sfaeIwVuajn1O4w3Jru17IewN3dH4LxKcYVhZewdqqKc4tsyhyXBzv0IEwzoBnG
aFLTQRBliUI1KmKoL9UIPNa+7+8dW1362EHLQK/+Eu7hI+YL91kDlyAeztxO4Dm1
NGdAdUsaP2bh3OKQoeD/ChFtfrItsLZzN1JuWypRzAcPn02ydS5EuRrS9qC2I/dL
JIqMl4y8qrfhqUXPHXYnPSHGwNE5lmAlPzvgABhYc+25c86MCFLXQXHs1v8V1T9t
LRMtjPpndORCom6TnRWv55OGROSTJ1xIFHqsvaurX3o8WwreU8JsZjs93DMcjUyb
jcenwmEGjScNNLRya2WdzSehSXbtzSsbFE4YDSpkHSc9GVMt/kYlbFWV3joiXz5K
n2r9HshaS9nDPLxt84XUp2h7N4ooRSrkmdmKREm1JlP9XrMMS1T+6Q3XaLnewny5
wprNyTtjnZveAc0XUFVTmu6YRSXp+Y6tuutQ0CC+2Zo7WdtoztwIWVf66hq7Jk1x
ANkAv7pLLUd2xnoWWGffJ+cCCQx0bMCUGB3K+2MyTxCmFcHxUq5DmCdWxvwMsXDg
yAp5emKBI6QRgLC/ybt8/eQFqCAA3CojRCdiQBweGrFXrXnyBmjcpih59V22vnFd
I1n1YBsbnGY4zuuF2xaWXtSELTEib1M/gtZsEDnhkSY2L2WrWEHnIyHx1asaGhwh
P9fFraywaJcGsV/rX29TgC0qURz7MwahlcwrwLVyfhuOLR/BCrbHRJKTdIpYSUGP
1nvUGX6+nfG3Rm1EHyqjIACd8+MZf/B8+jLYrLeg7+fNyTeY1uPxRYRmJt2pqWap
6HReCAWSAzKSniHYY2SpICbGWBbO+YME7cDYu55YWJWqaAGUssvLPQMrkcK9pSda
sZICqYir3HBZBXQl1UV7U9aHBkdHxlIQ0cAOiLf5XJWp4i50/ZZv4XJtBDtc4j0W
7/7JLHfTcY96WCqZ4cowmXnvco7M3OrS17ThOWLOLZ55/lakssiuIfDbUEtr01Wt
7aXsDyBm4Ezz7w/TA7+8fG9xMf1f2YKLg4XdDKcfxm2U3GDzkE5jhuEVfrf/2T9A
qEbIKHW0NoxRjZQsjjD+t3k/6hnOv7pw0Co1BsAC8yb3m34ojIrJtuU87WY9wWun
XlUogSUvnInxcZ65QDhlYZT2phDQsW1wRui8MG28Oz9PYSDKe8dTyHQDG7Ow7TkN
LdpmqJYOkyU8o6rcVWCGz1CIiT/Pnpfs/3mDoeY04xk+5r4OTn9MuYwvHQcvDvat
CJY0fub2DKLQEu6nQ3Agjk7kzSliRMWk8FHJ91BlAybJdbTOuv/lAJoG2XQ9tLpZ
TDk9C2k/8p1Ot1/zJi08bhSHr/KUb7bB2ThWxFBT1Me8IV6j8D1zJ0iRxF0gvhst
xqOXtnsj2GNDEMVeybS6keVqACD7J11xH/Ew7Ex5WNEnbM+m/6t5h7JHfj+wgqUN
HUBnlRttHT6m0XIkiWyktX0nPLjB7KB9Kt3ypuKZLItQyRsbLoTHkaIA89vO0xFu
XRt99dk0xcb/akFyOycLnE9Tbgz43EyM86TajM99+vnaHoaDljhYauyHTSkbpFIv
uGjIZPMFmen206uaLQaeQyiHuGcY+hxgUzepBZ79TOzOuroLOEm/lEQZgqNQ6AU3
nU1nG1y1Szei7aBzcyyMm3BBmtLNxqos2diq/P8Q3ajKFwm8EVcU7tdrgMaRnGMl
Cim/kW63HiUlEgN4t2WnRINBcH0B2+VDWy233VUK2KZMNL61PhvChPT+4iGjU0TS
ByKTtEgobNqV4oj306yfzt2PuUjJKFIequrLcXtJYJJL8l57bsii5zp/03+ADXUq
w43Y11lakra2R01QiDD93bcPvvUKK4U9ZN4ZTivFbNVJi/PSsXoSBmj1EyOUbrQX
jOdcV0qSHLxofAkfPFVAa7UYP6E6EBIsYw1r6B5468tNupZqQeYTR5Q4AG9vkg5u
QlyP3okwqnvKHpRLjATJA6ylvuBhG63ZMVG6ZyJkMcqdTGeCDfIcV3DSCNaT2Cau
C/KSidlvPh+QOWNlMIl5M/WleZVISzNzi7D6PgpxxfR00PxEnnf3Jg03GWy4W5O0
0QpjRcudVDh9keb5+Vg78jNlozt9gIDRO9kbRG/kOui72tsbUrArKRd2yziaMmuw
7zIpZBlzrCyFuqLhZU0WxL7U86cXb7ZIRIw/hH+qDGdrxVWzyvgNSKMFVWzYbTJ4
scWecWwwxtwtP6TH4UKyOIqhQBz9UA54KRo3+Z589HEZ3iPpC9jO1CKjuy455xS7
T0cIa8W1127BHM344SZjhY+d6VPXPO4VMx9hxzlooNLOVxaivzMWnCId9l+4mPRw
VmDW+iddxDhIZrgvsDRQZHo5AX1I5iSgwACjtaQkRG3d1BqQ6OKWaefRIkyvZPtO
Rzes4uNxZ00uLj+FQXzYra8V2gDIUYfgAOgIVbkFLbx2z1im5PYR2wHqaAcNsDvc
LiOJnZEOQie0ZnmSI0D7ggCBK0dsoI37IHEp5FwyZjvQNN/i6feaY24hdRVPKUcg
J5/uJDggYN1ZLfvk3w2zRUztfXbx4NQZwoePp0fX4ofOF5A/5M968TkKsBQ+uqh3
1PTH/yXhwnE7ZK+hSiZDMeKhOiNEYubTB/9PvahqDWpCG3HWLn5MWn2zupmpOiSg
vZQzeRRWdm6dER7OM/E1MRr1Wh/xIpf4Jdj9JxoV1PSmCmOEeE1tlDeZ5pmvqLhE
I3657YLxArobZMJbxzlfP9PPd0u8N5V8w5Vu0pn8tjo7a5TgC+Rl6ifid2y+D2Vb
xY/vtooL2QiIRAKeIS8e9yuUkVH0R2pvBiwfKANFwEmKA5itcckOkxaveJqvNM2f
4lo/1sX5akV/abTRLcZVS1k9lLM/Uzfj16a8WjTM54lErbJE/76ktvokSUSFoFrn
jELYiOl7wsD3S5Y9lzGN7ShjdSvBluxQF0XMfu07ro3a4kfB/AcypSi5pY9zsSu3
iVR3h/Y3R12mfeuhdliPYwWbHUAYJ8zyaPnUqp1/UojP6dFj8TnSGRvMjrGhNE1j
IeVlZcd8fCGvm0giKaSgmQNFb/ooMjB4YSRVRIDhGv6zHhzUY+VN04b5WCYAAs/Y
LwYxBQxW5QBYbEQZCK/PAR23Tsvui6gYBG/CViKHjfKqELtJHqbaaILJhcvYa2lI
JV5y2FK5CD48L4YoZGP/Tb68Zp4QzmkuDlrh8ad+xvun/0e6kBpz3dwWVvEAbFn3
SuIamUKUuTwdpyeOOle8akUyjya01oH/9dAYylIZV91yvPg8T7ry65UBQFBzhzAm
b36qaVXptaJfBn8p+KhcJl+VNFbFVc4viRwPpJRNAkpocAKNr5PgZ0iNjN2WEQX/
VBT1bkPVpwp6w+rd737CuMEBiW2Zy48KD267qbQV3RCQ1QXemzA2tcBLQKi8gZ/f
fLuP+R//vCLXAwR7AjGBlDzrAwb2dKYz62Ed/tpKkccdIumZWcFPI2uXDJ4ZNdtw
yMGQ9tJChJnVn2Tt+FgnkMwj0hs1xAfZG/tTZGiI/sMJkNh8bkM2HGzNTwu508Bj
9Q/7xicegj8RUFxTrRWkj63s3L/Q7PPe8kfNufu/nzjsFe5wcTfzfrLcH9hft9aH
DtICxO8dtCVM9O8h8w40G0Uo3EpsNdHKq7XvFotv2tJipMYzsXojfR5yA/NR3W3G
C40EdalOGuw2ZkBSSDB4KcMxXbTDr1aX5qubX2+IZEq01/LQGhPkn2ycd1ZBQeGp
/cquUxFc/7SNsdnq53V62GLfqmYU3WgRF+JKhfDDMxFOE+oAcWZRPnFxv6IslaRP
WWjNzdNs059WrkXP6e9iSqk9UIVCGN0BsZdiUlhPx5oy3fVr3lF1PP+96GTpYSSm
mCh0LM07BWyvW7ZlWkZIDNTOSwC8VW9oJCXRHHZgBuh5b1gMp5L2FV2lM69FWKdU
0l10tAhlG5O/4bqky2fOrJgTplyL357NHTyQHZssNe56q6LiQ/+Ns9rMfnPMdAnm
cjwUV44jVADjbbjmLsclrszAqX2XB10y1khLeCxKN9Wt17OD8BQIxyaXeKBR6Xa2
OFDh4j+NGBeWMKXHNjgxImLmdxvQZusVo9VHyx4zC4B1NfTGWaXSdkgwjhryDZ6G
XRHu4fdWbmaZzkwMMJBnbiEwoQPSq0JoN8t6emi51ABUAOKMCZS8f9AsP+AbIs+B
FZwyU9SLFU50o6Ec5atzBozKsHQIzxEzmfSBRVtFVviviSKbJl85MjgGz4WOWwMN
YLTPP6+NCp73BfgafWmoqcBMSGtH5bk+XpUDYTn1L+uS0onPyKRWFYgWpUSgq79S
LLcECOlqT/L4Ks9FD914le8fq0Uob92OXqZOJP8IfYliw739OaFIay+UEfdVZDWn
lXO6CbMYFXQbPaNRURhI4c8tf7JO5yVPCf9G6Wjf5HKEFebIXKeVvPmiDwblSiog
mlRHUCAfvRQXYlnTAR7InRv8VN+pLBW8XwFLnf7uBkTWxUoBr7QlC1cdhUIN07a3
sUkNiDNOLnP8Y5pLYpcjbNjsTVPIq7XYoKYpbXSA30Wb3ciL8bblAx2RwavSSO2m
uK8Z89qrweVdST/Iw/Z6U93v7yPl9/zFpVaA4TSw3DZ3JyxhHiaNQch+GbiSnrWY
Ra6I8A4bYlNnFyl5gO0RdmckFYVqL24yIRyMJ+I92t9mnDBPGcQGDCP8wPMN2gc/
ozxnSqA2mwXFEpuPep7K+8G1VI+n+xDuItRwIuFUVw87S42EQRVYw7h+32RWlv32
1JBMtLdqQvATlGT+sGeGKDmxh8cGVB8dZ34DENLnKB8VH7l+fBgx8yk9KlnlVwYB
ZQ4iHnGTU7qide4I0ocNEBGkr9+aENQLSqu4goMq4Qb48JVHwdsxn6zyzzcgpgL+
jcWXF/qmC8NXB32XSTX/zWd9jK47XM31W14hBkqst1yjm3e8JLeKS6CM7Jkk+T4+
GMhNV6TIsh2BCh51EdaUS3LIAbRN3KMBEOLUP4tVLwfT41dppc1iMWyq1OnLE52O
P9AmZd59EC+/YUX9Do8NjFvZwDlaEn2axEqHEM60iNe+y4KVT08gyloaYfyt+U7A
b3l7INAm+7hGzj9vMXL5CCUv2xJNVpG7FTGxEHNhAmqYzidQjHYGewEFnPAV1yd6
gzSgdUkcsxps/zdNom6SgLvQBtloEBHtenGgKPlxxZGaN6d9R+gKVNj3k1PyP2G1
r1yaQue2qplZPg7+EX6FAZMmHh8noZ9k4q5PVhzGbvL0NAYUYmE9gIq4mfhfQ3Qs
1kwQ0rw2WzJPkdO+xAW8um+s4l8dnHxT1k+VkDskDucFlvwVJ9zjS/a5iQ5z/nMZ
wWNWokt+MhBDc9KL+brTyNHyff7uthJjxWD6A+mEsuwrgjpqfnmBl4IHCMIUfd85
yJK2qcbKchBw9zOkXmKPck+U7DA7Wcr9Rj3F3JUYi+8QGyn04UJ0vU/x8EVZYtFd
HPgDnZVviUWpcaNWeP1SozOUr/SyJx9eqbDpEyrdMFzxKTT0RqKBSi7fOw1+/FAI
/Jdz0KhN8A4EvM1LKYCXwmDtm/SMhRmf3k08rdMdwKqOrOD5FoLUD5XwCL4T9HwK
7COCU4rgoFhPpR8mwN2mBpBaYyMYtBFyk3nbPEJj4fMKny4BuK0wkTKF70eBOe1b
3/iwx1C5bYRIxaG1z1o8ID9Zkk6zeE6gFYbBUiVP85uXVi3gAvy1unLcbCpRIWY9
Qhk0pZe9zcNZtNoPNDg9QQBu+d5Zg/43RSqVr5ibac1yugJyTPEgqXMGeQiVLfil
1oF8WmCU+crziz5jTDc7LzED9BWRQL8WirfRpksfRU5ZjtEBtINIsoQS7D55dyDK
LfbWspVEEx7ZGiLWdW+cJ+6T6eu/b7ME7E2W9DH59a40n8XXY+bZCwThKnJk0tnL
QME5/o+yjfaNZLUqAZiQHPCXwgpeXfJE4MLVAcu5Sg975KynBFpzKv3Z8wc7qnex
dkAFg2DubgYElwhVL8S6pZwf4OVKD90CGxGs4TwUT2xhb4eqx00hQg/Nr3EB/NGc
riKb0jJzZsHeWqHsNVH7Fz4rJ2saGdr0ECFN+/GS/9Y8yjhSj/1fjRC++EQxyhNn
6K+rH+HIXfxc/POefxRB0IXSkhdbWJD8j0FgnvcpFB+bk1tbe+AXjAj07rXnLX61
bMyZT/q2zjm2fodA/JNX9mH3HpavAwPlhWSFwcyyOdCxtnerb6/RqhRQbNCSHJJb
+g26yraurWwUFZcCEskzlgT2gnfcDjxFBALDPBmO/dfhynXAVmK942kVqvpCqa+w
Dx/ebw5tixJ0nsmUO+JdBmG4oOizhy9uVmtBrWyF9RNRN06saXu62eTAFaCcSb40
wR+uvi+p3GUqaqCvgF2HUnmZvOY4PLhCskkVz9SYo03jOg56GENKEHi2t+LeIjG/
UZk0ZPSifECnUR3Sw144XtZCyGC7N7Bepnt+3rEhsas/3PW36yT17cWfd+4gyhhT
VGOAUwSbgpxAUadBZHarwSXhVdZMcQZYMbMH3ncn9x1/8mkMuJmcgKlqs2H+ACgC
7pz2iRQQwJL3AuV9o0XYludlcjU1W9Uw61NkROfLHi5q1yJre0FqcUA8Ddj9WRU8
vJKUkyZbqjLqNDKft8bW9jiEyiiPfQbS+wATCYG7I2QlI3RoHrTGR8oYFGgGP1vY
cr7du8L3hOdM6g00fsRG5uvMFJjg4YLjqVqkL0r1x9Z/Gr37ymwhfl8rAj7Uy9Bt
JZHCUxJ8lzhyxbfi4gZWTco1ifNCl+IFEE6peQYe1CAjNzH18sVQT0IrOkCXe3xs
OQLymL2F0/fM5hscTQdZmerlNdB8cbYIk44dQhiBY2CDHQ5bPnJYaRtpxLzuNGN/
W+6sGcyonjUp+bMe3pWMZ4/pVqVi109uPZuYQOzJpgmfB0xx+U+E40/geE3FKhpy
apaEAbEfI36JeHM8WQIe3+1oxzmySThfjY6iPpGt+8WK3cBpd6AFCz0J8YpQmflG
B+SRsztJMFrAbiPwmDlqhc8QUqkXUgQqZS8LJDXCABLjAm2akSklFk1vINpB9Kxd
3Tvk+QGFAKhJDLVA8cdXVFzQIipHAsAE8f58KkQq/8IkaZ5BJhdEan2TLdb48pjk
eZ4Hm7FcWtmVeZanRE30Wl+a2xFeZu9K092bu6OBw/gKd9uJvGyjQ9DS0bwfoJv7
VA95o6BtSXNRxKpKKgwDFjxrZia1jJZY7QApvC3y8pTLO3fOdI/2OS8d9VUYfUA4
1ECohaN78z2xN4yLoGx/rjFtyiLVhquRtxaXoWnPnwDPRgr63GPeXufdpVOAW5LS
HMXtnJl1O+Q/WSN8L1V62RytoJUbaiSKLf2AY5bx2jFB64nCKZ6dxp3Y9swE1/za
SIGap+yq1f2bO9rddlZ9UOSW3vd/Ufv/Dn52c8Gz4ZZzwRzBMBb6F9kpsmKj4BaC
BucFNkGaZr3tzRiiGp+wYjNqB8MTIKf5PC1EnhtVL47oK26hnCtZUbD5DKgrrrj5
iU0Sf5LC9qKMn0phJfNue2zC5xRSiIaGxf4DZdmNLd7NNrgWXPYjPWr9wGdwXzTn
vd2N6TkPzvhPTF9yQhrNLjswSF2WavMdp8InWjswSn0TQZaElbDD5I9tcwlpiQmo
qOIQIthydBAEb0YnZ41+riqMgfqpJS9Qt01Xu57/Koaja44yTeCWGCtnpW0BaLIB
L86sxHWRBLzS8spUQUQaEL2/+HLHwdZzp7dlLsDo7GjxMPH+R8Jy3z5GYEUwHXzP
qp11tCsrXIMm6PCI7zo3noJ67bGL8xrRMPVt77ObRP6ThqneygTWyUs7zD5kvabH
O9YUbPvc3MBh8iBiFC4vkR0dLeMHAT9gce6k5PY5Rpfmb/1fFUceOKhYIy7hn0iu
pvuXWSh0FaAuoznpzLkx6a++/DOf2HCziCnBNsPYUs1Gy9ioFJ/UBvx4oCY50JTX
DOY1Fi7HGsqXJuMoAoa5yMxrDv4UA4OgPl6Mx+1rhZ1Ltil8LL6xPpAE+5esSTba
t6bNiFc2ccxI4yDdqYreqL/V6XrmEyuLnlqAw9dgCG8SQx8ldpLEyeolLFOE6pjy
6DckpfFL2uNu87ZHKgjJjQBPvqH8/KcFwT09rHbTcv/EjLXGFCyMaiJFOySP2Ng5
yB9s4VpZjvC2iCUcS8eNPdKSympei6Qd4xLCrjmj3Wq5mX8dHzN0GNPOiPIIoukr
n7Odyis2EaUQAJ16rnYpU0fsZ/qtR7kLxtyfwAJL/+WUPUiNFX3Q93VVBFofsZRW
g5Sk+Th1ab6CuJwyzDxcnylFOtnhkKXIN8vFB1V4N5zyPmLeA6WiOqkJUloH8zR2
5Bzzv1zMK5JZRPxwI4/pReWfW8+XEEzkCZEMZ7EQGCrvXim7azBTNu0aUTqCharw
ZXm5hFOMcc3x5/Tr+bdRpPvbtBaZn5HV7S8vNl2UPe1jEqWtR3Uzz545aaO0J/U9
sOLQFbXxcHMMeanM2FI5eQKttVGCr2yyGqYwWm0+actsmzas6FNqxpaKxdKBH+Xm
XU2aOGkbTnMwl90T/7/+5VYV3uxD/B8LyQLqwZYcTSOr5qifSLciLQscrlDDBqog
q0+x9N0/VGHThRt8OnUge+qxn2BDcTPsjSbcyI9tY5d8P2ha0JA/ldsIkN7wMsAZ
6jYxCbGlFcAbsyc658xkNR3JN24WExE6j6ppZpC3tEtLIHY+C9z+vJovS2uGD+Pd
Uzcjwrn4nGhbrQB9syiBm75mGOkH8yWjtcCJBLM8peHEzSqp9sGNycaBDW+XRYPj
peIfAwtPLH2QJCTEus7xd2W1oBnt5CyWLf7pOTOg92gRnlO96kRWGKjJDIlIg8T7
8y6NkAjl7uWmG6pFM8wTDvcyw5Fne8eaS3IL7/9q/C2HdbXwQvxLaSBr376DaE06
IDMFpD3wah1kCXB/f17USdgIqK73tNAFMKEE6BBfTE9oH+7oGK1AS84UcgJBQ8jN
gwg+Yj1l0tHImH6C+kTIUB+uvHD1m8QMKCDHXhI53CrY8TJIT/Qk1+Uo5TGYnkQ6
DUa+CZoMw0N/3G5mWxgRrE+zLj6D0kAteQRyDO1e3OL2dQlMi6OW30+YpqJh0xSp
6Ug9LxI1oX8hrp0N5xcxvWfX/fwaS0ATvJ3z/GKpf/zUlx0qtQyUbUVCh6uOQB79
elCmiYtSns/pefXEqKbKFwtkyX1oFXyUzernwxvt9913ffFWs8lhCdLZ8bgSlp/M
FInjzXdPXKUWP068CsTfbyVGkzZceX5HhOKar4l5Z8cxBD98TkfNiBhOpgjVBDLO
rpTS7Jghox8Y4zTmRuEOgEomGKbyFRUPTGm6BHFL7E8jUIcjBhbusbXI9b4ZphBx
aItWUf5vMOftQvDHqX/8576gxyQ3DOEfnLYup0AYaxmDTExpkDALUUunViia0pqM
lUwh+vWRx1wMh14+8zE/Oc1/F/cC3c3PRht+60F0ev1c0royXMdXZMz6LLGmtzMb
UETB32J7J29QkqcDBBA7DvwwM5Y/RVHt0Tfl6D/FR81cJsRmad9oSV2msY8EWZAL
0eAU4WzqVQOYt6sQeNnAatzTnq9HWqMQfT8YM5Z3oJU73yNPc/Zp6nwrWYt1SjDH
5EehEc0zBd4OZB3hUQFi1O8ZtkMkewIyjYtiNHZua9HLA8qhJ83f/JQ/1C3VskQ2
cw/1my1ch3R06yavhQ0diBdMMcMws3KPLiroigei//70TLQes7S6gFPVthhRyuRv
F15l8dwTT1OLcNbllCFSHOfiPtDESaBJDimprMGWwjWttSzeTk9DrhDfMtamLr4I
ScVGj3C+kSQOHkIt6MC4ciRHMsv1/yggBOoJT3xdBXnCEU3DKnvD0ApM0yI6K1wu
6ehapkFtqD5zbsgz4GhH919PwSNbxJZT3xvjm+tX5aNxGHG1EqcfQbLsuwsKhrNg
pALWtjV0pl3Z0LGmKEU1SQ/0QFkLIBbi28+hlmB2sq5siLNJZ6DIdptvon5EvRIV
HRRbfq9eRG7qYQhGCAnaYa7ZVV+x5/Q3BbRiRNFC21QFCYZLOtzD9nk8zQxsYd/7
1Mg4RwdxApEISUC4CFKww514jivQbjUcCjzWQzytEXc8EnpNXgUQEtoeXh8X/0hO
+1YAZsrgwu4wIE6v9yDmiTZUOqQXDFeU0lSe4h19vNYmOzzoDw7jlLtQ6RSJAH/X
vICQiiGp1rp6GROs2OeedZ9YNhuSQ6072CsQI6VCAv2RQmlir+EagFZjMu6HYqPp
y0x3xiDtVAiHsuJvd7vbf/kM3sUaDCmXbvOPfguyG3kuKTEl8GIwG9ojUaZ4MErx
xnupz3FQfzYfKoeYZJVk90r/zqh7gshibPlXXrysaw4IuGTRUcEJXk9yx7QgeSB0
qcJiArHF0SW8rT71+15AikVA24mEdrLnsCOCZ2Lph7a8JW20PDWnlTnK3jA9RvOV
sWXKkLGp4YDEES8jMjcj5JgFXQQUqoM2dG3shHcWiQHrpqKjXyvKIQwqTG7nK7mD
NDjzAhUk9RVLgWiZiOmNP1T+DFE55CKbAjhev0oVUHwwlzzY1AFZ7c2TzTYxA3Ar
m01rIMbnvW0vW6a79tn2R+RGPkDAVykBw2oe4UnlMpYia8PllvT9GtfrJqrtN5T9
+sogTCZAgzvlgtwWQRf3lia6oTC/nFX/TaOUkI9lNjqcNcgWxow94MwOew8QEBjJ
ayYnznxVc2OBP3m38d1ybWqAQqVH+tjc0UCR0Q5wVFRmVznvx7/NGIhqtH/MxZrp
4Cpr/AYXLNiNDgVTeUV84OdQFlEqN2W40It+4tC3d1QBjX9QQvswV8PPnPs8zhJ8
nKHuyM4Cxb82sHHj6KEVMazS+6LFF7n7LKow+YoulvcaK+T3lLBFx1d1WlglEW8e
Y3HgEemf/FgwkcY/OZTLZqehL7vHDZXImImkrWdU1O3YOqqezfbahaykrvLgiOc9
52vJKZudvGlkI0RnlCmJ4BjO5gzDahPRzDxp3kxPKfs/Laxrb41u8SSi7W6XgeyA
50X6z40N8QlURSnJS/OInGogID666p2PeV6VHEDoteqKksGZTqCeB8+yoz/LPpRW
3NzHSrWfNg2mWIpl0JS/I7kwbFzIEcNZArPmH4M2gky4zNuZLjA8dwO4NCcDzb2S
vsQvnc7xeU10BtdKltx7KF/mviIcDK/bF1f991vln3JkFbW0fILBhk8rDOuG27zp
3L1K/V630+Q0rfMYfnns/ATecMvAlt54sOM7Kr60fVeZrU6aShlu9iMZcznMF9VA
XBns37+TI2cXXYMgXpnV2U9NMtBGh/TTyJv+t+zJDzeTLTbbKsYRYLpcOLcC0H4q
U/BcbIepceBQe/pGLT68GBhTxDTerJHUKEHDgos60zjQNvVIfE6W8BI4HqR30mwA
l15YULTVVjFPO8TMdRX6jnr8OvkJEGeJDBCc5MftboLNRptqrJ1dqJUtZwmIhuk5
rkuSmNPHiC4MBX4rOdvXzJaB2SPFcDGM7IkhrjFHwUhIWeOSY2YIR07k2NgjrpLR
zTBEU0Q9DbTwPShAkkpxG8kO9jUCzzIPnksrtCPHyge2XKwkcxePoJic4hYKZ2lI
O8ZliFZtdMuB+SXePwjLiEXZK3k0YBRKzJe6YKxW2JdKs2WBFRqok1ipBaEfLdwz
z81CwBt8gI4R331WTBlL2XGTAJGY4D0CYiQ3w7YFFn+7rqvn7KeUgY5ZNbdSik8k
y4clzOy2cwD0DQPX8xPhJMmQXOv5zyPceOqWt1IvVwKAEaljCD2SizM0KCXFqAfs
XDKL1KoDLJvD7n5OtZPREz0NTcTOLg5ffd2YrzQVFFBW0mPeVl0gDiDNt+m2xTDv
G4L/6ELd/slh80i/hnUSBnlxdtvK65oP/tlyeF1vEHQWlrH5WRb9I+CC1D+Uzo01
RBHkghyihVXgZyTkPGJmEoF5p6qfx618GGUfGl8dQZBT61WSNesbDkH+WvW5AmVX
A+uudpaYA7+n5kr0k2q2ajDbSFLzSZqekHXfymiT1y7OP1YXjUqEKqhSiTvsjRXL
2gAJ25WyOtNWro2uo1j1XoC/OmiDjTZHl8wfLTpJwkYYkZMQ6c6qJ3LH2BBF4Jz1
Laj0wbIL4tlXDCayB6lbHtgjlWDsK+CtUx7QxEJnwQ1X51cczMWSomie/dAiIbAS
peWZO45pccvLTWpud6JjJO5E9kFPVK6zqwf3RhE4fz2I0yRMt9C36jRzI/fDbfZa
Y2A0HZoLBi5alD7PcM9g46HtzFqXydBFH4jxUJNWWSGIAZbkYWo1jaPRegwmoi7Y
pfgXjjYE1hoc6leWWZjDaI/paZM83X9PgLEcyIzf7Tc05p3DcOtflbfxF2Ccsj8W
6mRxXWQ2otjq5e99ShODjrDrkGmuzQpVcCtixwAgkorz9gAiAt7K+WGPNmi5Q/tw
6+HHh/kyXcmQHGp6DKnQ4LgNJMUm4G1BRMBGWaHeJFWKgW1ZIOhMzpSXQKLY/25H
a8kGwUBye/QXx9qyAgOJOur2wwvW0cPhD1RTWG/z64Otd4DKsgvYkUCcuJaOox6/
rz8PvHsN6111zhWfdgKIgzPiNEIFyiWF6X7Js6CeB3zwwR9OJ70t+uklRftKxqhr
757GytgW86HTf84Hj1G/XfAaYcJoem/Q05UrA+jOOqCauEqgfdmQED1A+1hZptkc
787nlfKy96Wix31821m8rkLO0R4Ia2pKKRfi7SPwp/XlsElhMhM+o1nNOMq+n3YH
rqvPk9FXi9RWdNlsv5Axy1GfqK2EoHaZZudsTatbyx0C3oh854DP5FIdCDTfFjnE
HSLjufYQAlGIt7OHKaJM7crgU12MtJZt1w8OK3mEOGR/tqzfMtE6Z34fNvGPpr4E
R/PsBnij6t7PvxM3jp5W/iCPElJLP4H60MqSke788159nxD1LDmebasZvv/6vlH7
kZzGuGh/JafFo68n8t6UKHJbaQymAY+FUxKQi/9iG0O0RFL1puh/NN1uGaDPIGlg
PBqGwgrDNaC5nwHYrwzfPl78ct1UAPpDXlFl6Cw3LAU4JygL0E6lG/sh0pnLLj/7
COyZyzqBXsHU5IWccGrOiPpRQ5h3K71ki2pViTM/sDz9f+x5tP56kYai5YXAzd6p
GJo1MrCjuJx4UDTUCBubIwKX7K4YAP/cvFVLE01kd5sR8FGzvoEjTfn3S7Lkef2w
ywSq/76qPzJ4HJi8vXkYDDXuX47tgekWTGtXGhsXRFJ76lz4ann1+BAf+yv3Fo4Q
wvGr/5r2bIhpdw031wDHpEyxIBjZy2UbsBuIeE714ifyweyLDchPdiS7deqjNYKI
Qep7TNHAKjpPgafPtH/AT4fmCFAnqrC/z8jIJc5UN3oMs2rBvRWxOaTwH2ymXcRF
IK/VuUCBd3WF0yzrVLjWcd+qMwhqtYZfs5OfmikDVBA/IdewXPjkjM28cBwxT/2o
HejDuNwvEVR6nNHOFdlszVU0sJBHuSdiCtjW/IXxotWJPw9ir2lz9KvxXGy9JXFY
+R5LzPsT3jEcGHyUMdejBBy4/LYJDn0KD918LRdO18FHIEOldvqKfjKMwpd7zw5r
F4DVZc5+iLXXT6A9NtWuBWhOky52IkXdwpuB1z4Rhwo9FmgVUFNxOhHZZEhkSYBh
Bjvo7DbrzMaf8QoSOahnMx9k++kZreB5afrbMt3QQ6RXnSlJtGDY3kE6vP6GEJpo
kS/dn3txIcRbmbLGkzTARCL0jqRaQCH10G+Kk3OjCqdb+5Psp56J7uH9o9H6Z2my
19XYvbLMRcE903AtWY75s/yqsirGdBuUGFTptPw09GwtUbKZ2G6e979suohpDwiZ
LFqiHhlqc3VMIimaeNGYxqNqb44+QBC1L4CJE1bRxWR3ANSIIVjJrZuv5kTcVDi5
noOHy04aL3nX4K0CbqthA8OBUeUzw3mZCmIQUFnsj7Dh63/M51HWP3veseiU6aDC
P8YIwjcRX46+wDfqILRGqIqHMDnJymGafj1pJG/VflJ2dMNtGbsx0nPpD7e9U/Bi
1Iy8wta5OvBgq40WA8eN1hpU8bMudVz3NEFAJ5KMYlOX567xvS59kbKMepxNzAPQ
+Wvwz7Q7JRaH/xjInul4K5+ExwQOtSp6DRoJTqbsdC7yc4TDpO2Ha4Q6Su/6qN2W
hp+ocP1njyLy8iS19m9CRA8wy2AXaeJmwlqXe4EG2NZVLle96YYqI0NyOiQ3miXF
uRFkY4frNjLN0F4JjMBi63QsYpjbtwbXUru9de1tTL/tKhse7e9vt2nqOAMZbHXR
vXmt+Jhzq/7zOT1aNc2OuHFFKnxaLIWqTzG+/qBCj23AXWA5K4vnyJ+jz5q+s1lS
aJ72+ua78SIKgk/HyRo2ZaQT3xfwMgU0SBa0LcpBv04hO+c09fpMmBhkWc3NSU4i
k6TQAcsvZIfazR9NdaMTx0JkSHVCVbraTPEHz4SY4nxyO3K4qZU/I1jWncuhzvLf
z+j070wZ4U9YGn/veDmb5p7o7ArjG3V2iBJAgiMBFf7OWqFgLYouoKNSdBSZAaRO
aKOg1E1YwPr088+hQZUAIlgd0DuRV4zHIxVxibDLOuwtZ7UKkRyfvZO+PrqI/QxA
kuRp4IffaKDeA9gC87/OW7+TemOgW5oha/Y47QQl8vRyznaG5NK/A9ehhIVbkqs+
ih/WjiZAtaK18Td5oSUbfZ6Zygt6kfR5JxXLaiOEEJKFNcRu1u0Ej60x77/FsTmo
IGjDSRlvtiNx4mC+jmny69xpocdcVQrlJNb3imhaE79ang4+DduVfVyE0Fcq0ZoA
eqZX98y3GwlOY5qEKQsSFUeGcGMzsTN1PPzeSNOpFD0QBUcrIiZi3XMcNAlUMGI/
tO0dLRswE/X4i4aUsNenAg9DKSnUxFnzoWshN7FOyBSvvP0mnlgmFV/567NuxryZ
IVG8FZVcJAZcYtS6qky0xd6PPELudrzHpainKZ4qYjrGVkUXVRTkJgI8VG8qLCr8
iZsp2SEWqdb+VPCvDLret/om1LazcHEmh2iS7Ff0soglyBVxXr1sBsCyxhGivadC
Tz3IShPzpSzqJVgcv9rMsMIf/AE4qqODApwwr8xzHi+9sbGmb0fotJjIniW8+cX7
19evPzTgIi6/OfsrFGinagKUu4wMhBr7gv61Ixzz3kFeXublC8yNTbxzvub5Raua
wklrXiZeVE3q5iwePsPokhmAWBSu2i9byaV1/a+1hTX44cGFLwKwmnZXZQj1yFTA
HtfbyIv/d65ZamZRkHaxWLhl6zERXso/pUZzEgLX4QhirKaZrL/06foTE1r2t1nC
/mFTnkP+pbffbG4DHuSeC2gmOAWSRdt7uW9UrBmzUDyRiBM/Q/5scJsi5+aLohV6
Arajnw4fp6otIgIYb4wBwYLfdNBTXMCMP6NLr4L3TuWhOYvEiILL2NDRCUMA+Of3
8nangH5xUTZUPH4bUGYJmt9pH2jtRJXtQPP0HtV8qXg7DH3odnvzj18lGdsuBkD2
EoprQhq2uMeIniVJs164KPrigcNzTnxv5kXi/gm1pJ1azo1ldYnG0QqNZXD4ZtBs
XwMMDjuWuBiUfKcCED2YvfXvdtuwbHy//PZEtSk2KcYEN9uJI/9qJSNO7WQBtuXN
6wX6awnC7eZ+bxMrcJikFNmp7GnOmYBOIqjY1dDZpYvvWKxfEovLJQJG0GGRcCUb
WCJUwexAh3KescBeynvv1QZ8Nyk11rwsMh9cFXaIAVkNV4iAvybk1ua78cE2cLuQ
6M6DG8ySCnNPfM7I9Ud7oSgd7PxKIc+QkZW9gCqi2xYiGoRORKTo1IiUg0VopoLM
7K2UxCV7beFy77APLyw5C4aVnPtcP3XFcPwlepj7B4N1Oi/cBQHGAXKYhMF4mKzH
c028cvn5LRpBkh1n+Cnoorj1pDJb4xvjeuiOuOFqpcHlqr7B5v3LLbHwshZ5YZXy
T1UZkBWjTF9AWbIDx/oR6cO+lHtSJ7sz7J0vbmWi9RBNgg3AHWwgXWnuQorwlFzx
/SSagyoG+T9VMDZxAXhEZTV5RqG4m1754DAbI7PYF3eDuRpFGEOVb2IxxcPFrTtP
kPJ8mW2oFUrFJqonkdOwmkwW+UEab7qQvy8LXOFEr9FO/HgoGYPJxrdVNH1chZdY
+Nmd5wCDfWkSStTpKrQ/x7uhiyaE5MFSY/XtpKW4nX2u9zUI2BhMvT7nlTBTF+I8
AyMC2bWDxfU0hFBpP58qqLsBpRSwI/zDgWq1y23nj7pb7NxDiscOkZKr5cQShNHk
Vwbe/MapAdBJKYWd6Smh4xOvJbTvqauriB00Z/LPCT4mnhSbRT4okmnCJksbtYJ4
c7yAEVIo/kEvRN8pEKYxIYcsIE/7yZ5sQ7wePdrJ9O6n0m/VQjv/0pnNK784p4HQ
kWhXYWSlXlBAhar3TpbFf9T3lCVGd8q6C2sGQPE/ditP3V8AMpU7mUyI2tJVz/iH
dWDF1JJQjX7BqTEoF/oZjDLpOvtO1LJev1+Th0hThJAOd75W0CH7P092jXgI2p8e
60n+ml0ZEK9sj/SCSzqh351y2gArvWPdhzLhetSpZUHFaq48loD0yTSYzNPmRbeu
UnQGTuFdnT5NxSzlU4uEoSVVGw8F7dKTtC6N00WLWAox2h2Nqw81d6CjQTFvxwFe
dGgFTf1FoRcbtJNDCpXfDKg+D4QGsAu4rrg/ENBabTtA/BLf3CME3hI/T3ee+WtR
i5bcedJnyU0vWvMDLe9OrFobjvRSmdtZ3zWNcHqdqplp6z1qRAB5iLHQH4sqZWk+
mWDQYbtxeD7DiU9gdApu5PpIr+bth1o1UpJd/mdZMvKt/qopot8TG7wCRiKZZkRj
1dh58oGQ3kJ7AMvv2xeTiIpgqz5ygr9/zCRiEuRa+CVtpCihCIk5+nLuNbvacxL+
Cmh/aDYE8eo6bdOcySfEa55RcGzjzKginpv3DOG4X8cO5z4Y0jSXosL9D1moSj+2
StAdjfqhCPlkRVPtZMPwNBvCNoPqx4jlIZiOlq19F3QfBsFyLhOfwOIowprc3UGG
V5l7/naD9Ws6IO7qWSju1Azygj0KgNilOWmSS54DSRYEWck1Z+5tHvwV9g3cOt3L
AXqIR36/PmXs2oy7Ubt8ZRWiMAHskMF05HA0ovGgrpE+Nd3RW7b08bB3z/ffGzGn
oDoFUaKbBQDDxPpgp+VF4UHoASkVSSUZBVwQhIt92scJLFV//1FMz895PBeuyVf2
hcVkGAyTUyV8w/NHYVyHz9XlSE1Y5+xRk9xHR5bSgvISsIoH6cHLbHUni3mXMTLu
bTf8mU3mKnLfUq01yzgi+h9Oee3xgNGMDZszpmynCrepZ0Sr/0SHBBAirc1CSbmR
L5RNhheUbRq5Zc1CT8UkRZiEbOwVPQa84sEBXiE5/ftcwZTfPkaVeTL0WcADWYyB
3rzNaa+SVgnj5eplVv8jIqYC56rAeKkmIyUcUUlnCIgaoDB+utM6e8rD93K2LVs3
Ht10POzaq4OSPQlX7MiSCqFfpHZ2HXPMT3hc5yQ2ynwxSFnG3g9JpWrbtEnUlqNL
q6fNOHC2gGB0Br5kl5e6g0anE56FxpZ2RxnR7AC2Hj/KywVfV5WUoLaclkqZahj0
fDpeNIampqgKVE/c3jis3c+wxgn+Q6FMgt5UD4xIf9s3LCzAFsmXfsfEDi9Ytjua
vW2x1XWKl4L3XW5pi9Ud/wAAn5pOFHdedfR8lCdrK4JAOpV8IF/f42SDKN+7bZIn
oO81s9UR3jG2b0o5M8SYr3exVGzQ//tRu3fOtoOVfNQpWDqwUslwLecNXw6jNRGi
vlPCV1DcXBjMJeUcznZ2WO6TtElq1q+N10HfNfQ1m+sk79Usx+nNdVe3gJ0VnOGh
Xd5kSbmSht7u11IXwMeHD4fAepIt+Jx4BHlNZFsp+V4m1jOn9I4/XRQjhmBrgcf9
rbxNHUOJW668Y3wct/XsiSMK5STZlha5i3Amyb2V85Q5O5cWWt2xwiJSMirNBKVu
R7ABgll1FVmvc248v8Xd5NUQFXMoPydk1c1UcHDNzZqpQI6Xho3rhHuTTy5DyBY0
vrYXpVy4KuWfMgQB+0AMg6nyJyFoFleH8xcJuaGcIBFKzvA0ov38m+vUNibGxbyp
W0HK9K4D3jbZkzyxPR4T3zdl3rkZNlLPtvotAPca/eqAoZnKc5pKXCbLczp10cBe
5C4YBPzK7Dnwmat3WFk2DIMgU1RCHgSPAkbWYUYoFv538u9C4uGBoMf0BHnM3iQ2
vNlyoRR7unwOTGK8u8DMYTAdlGN2YsLIZr9x8UvZg7lcT0jD/lUVxb22kjQnN8Xq
yAlmaAjD2Bl2DFmSjGhR/4lf8FP3GajWdSqCkc4qv6qV4FXDm9Fr8bwJ3dDKb0xc
l58XP6zNQ3Rbb9SdK3XBPdlfteRS01NrUa2FVqn9ySodFXGSQP8FMHoIsHJsXgcN
TN/KG3eD93tiVXU5NREGgK/muuBo3EKktLX4c5u9Hy34Q6PyhFLj3wQJZ77b0BTF
+GccFqnC6VLJt/doPoCPsPUPSPcElE3Yy/ZJYkexz16wrKUdzwnlvgNU6E58kNRL
nlFtalA8SD79FwaDiy5EkMKpdyR8uZIfan41PO7HNjSFMN7rlaE68AcvOlfXhvbt
q73gYOuJKyLsHHdfhY2IihT43cW9NiAZzor2RUZJJUHLWISljpPpGHwvhyygzx3u
`protect END_PROTECTED
