`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TEXhjAeKLi18Z6BQWPtiYMfAVVUTSmNIVAS4pW6hjP/LmvDCZ6s5UNnsgMbuc28c
Knjh2zOcOneIkkn7tTyEwCcogEZV48kH/wWhD8yDrNKGJCDGHwNhcNy1OG3x1uua
WPEzzvVxc2J8ghUeyvjRGrJ3lamOD1CrKPyM/KgiE8eq1KwIf9Pnmz8YJlf2dBjx
Jzfhl5dwTxdnz69z9r3DqUBsbc3Iib4Bs1jgNKH3+kM4PTXuRkGnEoC/c8cEwsDb
rN+HwR6A8Mt9EwcZW47ucUUAFzl2lfYOsgzNeT755kCgfJPiqc3aYgyizymyUNTF
lmTTMqAwrpHp0wWQTVXlRVRP4VltSlKCQxTt7hce4RvsS2Z8hXGi0BwnMbbgMVaM
MzWUNhkjOnY1X5N1tRqCn8Zri1tWoE7B9yluur/Z/JIfbAwd0/iUrUlFeplRxhvM
gcYdWXPslWQz7MERaN5RNxR/PFRTydS9G3zZvQwm65pZRR0ojSSQnhrSgpi6OhpA
2xrFRu7Rtp6LbJOSjK1sPRBWdMEu+uzxflaXX3Xc6myQFi0fiKYkVKLl+W2B/qrb
+bgv+kiqPxspeABifKbDYDu8EUiGvmYBTHtOXhbrViQ=
`protect END_PROTECTED
