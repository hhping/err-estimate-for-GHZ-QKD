`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
07YJidFRS1yyCSp8eAD+vaixFzYsVeCYkT3ycFBb9XrrubLTOsFWw6imrIMBT8Kg
EFMDbhjIzOFymrpNAVtz+OzTTdc035CHttlXhUCzytQZm0GJCU3aHwGV9iyRAodq
p9isLFXjD/twO7ZaF8Ah+bMD3MRfcB9RKPC+Fh1Wq+yyZP+vafjkhSFAm/c2zqQx
prZjVhWy9z4HcdP7iVZqeMP3xzxgPA+XErt5hyj5F+iSG3ZuRqFDdFzLnHaU6GQk
MV2uzTW/L2mpTdugHrIcJ5AGXPnb2Nq3/ru9GP6uWQ75wO7URECl49honi9EnzY1
GLKCjR2XuvuFiNTnDts0Yim2swkPp9v3wR4t2v/QDWzagy9jjL1Le/n5rzpG/s1X
twfIfIfOzPvZEYwqa06IcPhD9moHwVat4CNUtZQykx7pblxhIIWFUzmBx451DoeL
BmhaHs88EV+N3kYMhmPnKeNaoPU8C/6O9Yel1+M3+aejpRyvAlYs70nOONUyLacH
xDgQtjBGEKWTCnuPi7umrlelZL/qufI7hXDMFP/Bx1I=
`protect END_PROTECTED
