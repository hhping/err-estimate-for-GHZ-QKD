`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sCOICipwO7oSj4hNtBdtk+bfLJwLSCjaf9xc+UKwzKjIAi3Y9BArjLJUQknqnAam
hc1lo8rfxmRUFx3B8TEJ9kt8JodeQbF+IuQpilYk4yLmOQBf/x0gd931/0fvuYBy
UQdmywisY4jLoD2dqSo5K5V5qqlKUBPExvyE6AV4VYb70dduqb2jRs/V9LYNI5oP
mcaLDuustDETuxxCJBNJPs5YK2CPWayENRNfq1X+1MW5XPjJ50avtxkGqE4DgzTK
uJtQyx+GzWGng17SLs0hZE9VZC93MjNxZJtaCub/ZWdULQ76ZBt6iV1SSI3wpgHx
zUtj/k3b9MTeTnVf3TslFkNC1vootjNpMrKW0HfG9wnW6aN4o+Ys8GzPccLxhUjB
4GJOnUANLVVf0Z2re7nmqxQeb6TzQlcUGbhCjZX1+Jj3Y3/krpmXgPI85/cpNUVZ
ep78yzcyzi5/F2loHLtfWkBX5+Fc/dLQ1IR+vhXMUyBH6eHwe2XS0ubI/qSQo2mf
sYlbwbhz7ByogtrvvzI1CqSiD6XrLS+7GIywkbtS51nmP2vEjitw75/d/iGhSXfQ
wUgYLMQb9gR3lkS7UIHrpqMdzLAzaL1Z5LbSC/P8N6J77q26mAk2ct6wlox7ZVPe
OCVS1/o8L4ikt0CgBo0tsnVQcFuEVP/1+N+OFmeOtCrppN6EW7VsFUPeGxDy/0F1
afLhxiwkel3u9I5xmvT+/ajXUXo0pXDkRkqeX7FKw0E/B2mGdJIZfso54zhH759L
sdjhHZIgD+KFuqzTHiIV7M1GXmK1BPpsCKgRL15dX40G4q81fK0Uo9XpPpmkyv7C
MYiEA59fy9VHMFCpjUS25fsWQu67HJjcVMIPnw0WWYFn8p7AJzd+lTV0jvlQLt6R
/56vA3MHM0UDg95xLHtJ2tZZOYTSlGet/tbe9wEUsNYYJrFItNmDv24O4Ke5rG6A
LceBOg5mrxl4yRG28T3bfG3X0mrrjkTsa17h45zxxDUG8qNRUwk41WkzRBTx4BTv
lVfAlLqsWSNFc9ievMxZzDikRJQuYbzHhPcuqxgfBARnjTZYqE/LGaZFF1MxbK6U
+2vGd76VkhevrHnbfKRof2jqfvjEIyc/M4bpL54BK6Msu1kKak/NkMr1eTKMY0eb
cs180zVn4C9q31WHF0BtXeMhyCKfgF5L2kuDFUCTvP0WQB9unPp5ksyRWKyPByCJ
PpyZwShuFO3SMHbDCLIubKM/+92dQLZAygzAycBgCFF/3uHJX55K0HbjzwC9ltBz
Zbx9kuJyY8uSBoOAqR78xsyZCeWfY277JDydNBKAw3mL4g+JGFM3czbE38LIwjH6
d47KeeS+PPoY4t0yP7lXCRhFtQyAxd4sOq5LrbYtRVVpAQwICl2pjge2lXn0GMmo
MlUp40oC2kKN8UGrzmcG5dYrELzs/s4cSDSDXpZpt5Zbwvl1Y9G7x/YR51HvUWzR
4tWTgFx2uhclUlRXGSI91VMooCJNtS5fkiP+vL1dHJOCTps1xaLBvRRqNXRhv3wA
axztnX6Nl48ma2nkUzJApXPY4zVJBUxVg0tow00RwLvDU7v3AAL38Sssd0vDW9NN
xNMsDEzu3pqWP/I7qWxLQfMYPPWVx5JuSU4Jrb9hbBTZB/F+4K5FTYNqcjAR59SM
QZRN8IauRgzqucQqIqUjoYAzt2A2/i0Awwe8lzhDP1SLAR89JIYkO9Uh3UiRGSWo
JmDOZEGqOTLZVL+uYfwpPmbMzHH6O8BE1mZrEmcNCCMN8r5QIEbTlPNVsdQaFFBh
6mAULpDDe617fQXPlMC1A75/Y3RcYumMMhWIXQw5+1sq9IatsuoufRXerzqc0PFF
dVVoq1lT32+U50qodYcGWA==
`protect END_PROTECTED
