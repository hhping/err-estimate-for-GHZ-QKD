`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xh67c9Qacp2e5036q/6woQXfNuLaHmiYLzujaPBfrHwQWUva27aTxztZfmMl6FYz
DY/q8bSoEXmhDc3cRNx72dTTd4UCqt2dI51gfgM8ws9Pe1AqjKo0bHFIZqwRtNa1
yIYDBzGzeFYUWegU6amnGrTAmG8/DL7lr4QwZxqZxFWyF6etvUK0wRFFOFlpc112
z+iLy+SJmXmWnF2Ninq810HTExZG4aoz4HRSlL2EzfkzwteBp5cYJlk6PNMiSRm5
eWpycSL9sBmQLS6C+fjUnycWcQOiAwUUgLTZjrh8zJ7vxqFtnyDfyCA6DkDrsLOF
T57mNt9n5c9+jLJS9D+3BFAmpbAAsyYMKiaZIEqgjnIr2E9uBo+36Ry6yZ82WgAV
Jg/3A0HutbUcsr4KvcSaalFlhquZS76CKk+toTHeWK78nZgqtw7dg8ubNqOkri4E
v6vxEIhWe6EjE/OmF6Inc4OixIH2D1PK0LaoEtuY2y7YobzH/tKk1pgD8Hzzsymo
yehviwcAuN+aL/Qv9qtKPJv0MHCOL6OBhOn5C8EIBMYRdmXvv7CywjrZKupO9mt1
3y3PdWfrJ4FogiFimRzVf8kx+VS+Dv/GxRFmRXRRsByFJ6ioI01aKnt8kB72F/Qo
/kqsvDcQrQArTYRuTOT6uWnc9jCUMa6Kg+32rbGxlCQTx83R9xc/oS+7vZqv05/g
kgIkGtuCDAqy40PBbdb8wyHBNUgO0Ma4/Z01CsmhggwIFCMPmUrI0Bieh68W+zZA
OGwk4PGPS6a5YRw2P/WDsfUH/rV/Fp3YkE89kXAUq+g5v1E8GNATKwHc5WZUrTZK
ce4YcLXHmqnRgEL50stm+MASq3JAbdH0c82plpZz/oUQ78/Kh1kf89XtlquWYX92
tpSoJFfuQQ7bNhGtEFSmk/Rm/HTBOBFKdkxmoGfQFgTarOTzZIc3L+0Ed9skh0Gi
x5ls4pwprbfbQxcJxH2wDzzKovE30E1vUh6iWdmfNu9V+ej/1PAmatN5BDFkFd7q
p4/7h9RSm9LBSh0+w2lXsbrQxc/3MOfax05PxF0/yUVcDIHBCbTL4J/cwLO31H+P
PC7owMEfSzBUU0PGp9mArjIBUVWhqU78ALDHoIrglzmsw40KrxOP1leupG3qnMTK
`protect END_PROTECTED
