`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FZDJwDSwFZdkuyfB8+WyXknVy0ci0AjvFLXmdodu4WSSngP3obKaqFaD9EgRIu3k
EmlpExjflxf6VYsP2Y5+uqwhC9mC5wmhi7lW1F+j5xMLIoE66TgItv6WBebWPT2J
8WBpxMk883HmauJLh3/+R5twZz9p2qnztSPsrSefhUfPk1SQMkD/rvXpMZhAPe+1
Fh9Tn9A0Xtw1B3X49tgBOWLf+USNWMajMj2qd6lqFY8fHL+f7jQ0021RIsp3A+Jc
haQmVdVLQ2iC+H7wkLmVu9w+XGjdz3PwE5rdFQxoxXiJ3Bzxe3xQXARPEmVzkzAk
Y1vESxGFY9tZjT9aG5nB59knQPYkqy4y69x2E7xkDG7zQJ8t8Gbp72Rp+D/d3oox
LjIPn2ljCvZ5svlc4fOgqx+AQINen9NJtqGkke/9UugxgtcH2iOoOfeem3p2qE9g
QXOEI5o83fNFcvrAdj120vNs4EOcSI1Fc/sC9f3w6rqxXde9UMUDVM8Sez5pQKQm
LohnnHge9QeqpneQ+/1iVhjHhgrtOLo44lFbUTMkRQ5m1wFOlhnPxoqrPIG+62IQ
gXFrbkcH8rnbGd1PpiXc1DgjLQM5YtK9takR6BjGTCp+pZi9quj0lsRZKP1QMMR5
A2+qevAECazPLDxg3M8cXv0LjKyE1/MV+MP9hOcLnPNMLtMY2vRjw8H9KVv8of/g
KZMz6ubsqeUgxR2wjhnHfQtYNvWkUIgwTMI5E2r3P296IlPMu8cALVFCj5jl4LzP
FjApZ3rSi1Eor9AR3r45uzfZNLq+YqDZm/45wwuTk60=
`protect END_PROTECTED
