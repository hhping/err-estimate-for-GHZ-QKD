`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TYpewlDo4KTaN49T+59AZObk5SvZzKsTiQq0FiDtR0pw8n4g14biAOlA8zGBsXo1
2soolY+lc7j5/WiKeTQ3fXDaqnqCirfeUjUvFk6Na7DrFTid0uxtpubaxl7oAhaY
7X+5QTiDQLwb2xtD9aUoWVr4XJPRo5GhibTL+RMGLLklRf/wEjsmfW2aPoz/FKup
9ARcmgtQcvCXAX7GZkauAI+KrjWJ/SePn15t8QZMRT6j4G/pJ4VxwZ1J+zapW2/M
F6QiqPA8nwd2abZ80+kohC93XvzB9hILPBYJ/zSU41X7DlLGZWnOY/M04K7K+q3E
ltRdjq4jVhOptLFIjE+A1M81+sMTzyQCM9M9hJnRXhMu8eHlZkBwQkK6sRPdqqEH
V0cy53hpQzxmI+VaR/Hasd1yTZ1Akif0swFleTfEB6u4C2b1UyUsAC/Sk2DlqkIc
zTv3d3618MORjpHCGZTTQ/ScLrXXOJ7cWcVWL+LTIZ3nKVcPNTuZgA575hpuILpg
IhQ6pJvi+YckYeAaGRjY9kRHqAjDOv4WBpOVwiJ+HWtJIV8R9GSKaCGWsKCVEWFd
G0RzBrC4siCZyHbYQiYdKPxGxeWIw4rzYDAjRwgT4WKdPIb0mU4XIOrIzDZvJtd0
ghmc7Q7s35qwzQq2PWRHOq6vmqNX1dD+Pt3O1lI8zJOnKgqhf02IygUIWXiBUNB1
OEjVur/gCHPQMyYqIRp+k1wRtKCxWykCxD9EsERB8pCyQ125UYSzpzp5XcOO3LfL
emBz7ngkegBQOQ80QljJGSj4hDeF10xFoeq8mgnq+FcIUf9smnX3Q6iIwRkJxBxY
mbquv0+ZNeHxcGb26Zgb9PEfbg5U1FSMuEqfRRyCrHiMP6hivTdydAic1lDMe8+l
ZMw5Rcm7e3874TFcnnQh2ezMUO9+gleV7WrWCOih3zfjIVeVu/I6XZikZ98yKKfp
Da0O2alU2L5iUOZBUJGKKr9TeFG5JqSpS02ABQ905wZYgR12bhtrfckLedNvy1TH
X6FQCBC3r+9J0Gvz8kv8AFqpvRO37S1jxA1JKxDfxlW7F9Aekx1RpI4prsh6IOIJ
hfbOlTcCZI6Nj619FCJBeyWomvJKK0sk+xsQfZPezu+aEzujmpy5rHqrzEX1OrVX
RTCzf8WTNrMvVHQgG1yJl0PV9Qkn7ri/Ib/UzgQQMl0DxT+09TApLMpLIgovXrF5
cfUrzQxbXTE/YQcoSr+aqEhvLGlbFSk3kO1HSz7WJFUbTZT370kSCr4fvY4a+LR7
M9jMsKQSDkKzVzofLkxD5WtLpSFZrgmka/0qRiRC3ZFHp4KbYYj8x6rXSOKsfJ5D
oaXzauL9WnJBBkmLUAndqfyS4fx5AR6PbzUl9aUQJlqZJqmg0im05JvJHByoK/Y5
5pgw6+mg8/TdV8bnB2ERRLDUInpn19M87qfUi1yA2iPfQDn1YXTvVNieCkPoOI01
x3y/gG77ealIpNOr0lDdtzd2STbb6QqHAMYsZJj9soMUW76NVSFsHkG/rLyUINEt
Z/mxs/qLIOmlhhetNYssfe2FkzITa54YLhYeE2+SkNvepJRkQrGnEethgxPEbUjx
KfpBC8xCO6+gq6oVkA05A6nADSkl1HuHzPFhaH7LOaNAL4nN5ZGF2uuQeuWG1iT+
reVgHTEqTuoohJnpIMBKYiHRLIxGeJ4TL/O9+yn026BR7AcVMqafEVGzy64Bkh3o
ZrLb7aBRrez8Zux1ifpITYPoazSpLR6bJ1Wj1jl3hYuxfsfwMznxE4GCUY6SWnWa
gMr20TTZ3aLs5/fUEJ4LJwLEm77H8V8hLLBNFkRN1PcgTgeSE4WugTOOAeYj3zX4
1dYuNacDEwJXmpaCGLdAV0oIqbCwh8HYc9klgUbGoC5bV6l9w85mdFokXZru5sda
aa4Mm3HyRXAQY8mOttU5mbYMWTUNQrM9P2eKxggitCXYNfPVZQKjyJE1rk5hVYIu
LlLpDgoS9jMGU+jLGiKQ96ld+7jFnC6IU7OzLyTVLbL7wNNl/3bTdtyhVRQjNm6a
bec+JgxvOGt/mp8Slt0JxKolB5zVDmpGj09kM66wkrUEhZhIm0FSj9kz1fFS9EmP
hLWCC23j827vzEQNHkz3GuZioHfolkYKkvbmnlURUO5jWRX0+k3VNz8mWo+sAGEe
2cRVOwbpjsQJ65LJ4ieK1y4RI1AiHZZfoU6lMmj7xBOCF5ZGXAYHiSedYnWJlGrR
uA1kX42Pd3/kdtWK6iXNAZscbDd5xmu9jQXA4bXdFqWc2CLJnfIfdx/5Ytju+qZy
2rBZvndRV2u82U2n3h3vtE7YZK5twSNag6qGSgl+gnWilWFjPo1EwbQ0UQP3U1Nj
xhJf/DMhnGYqukqS5zE0iBwThSBpng7qo34yK8clio8qpuVWzcqalqYAFSjobVKf
x4OIT0hI0sOfD2zxXM7sP2RPjMdfQU3MIiikZa0MiL+CRwg9ZFnt7+FqDtlkQ9O4
4fuB8eW5MJ6bHqTRQNj/+kyNiHg5PQSqfdH6kGhB2c/DMLse9p6j4JFt0RK8AUqc
rgEweoOQv51n0cC2cYfQgxsGEcgjrj9eFRf/n68ZN5BeDkAimYOgYSxFqJ9KLUIL
q62PvPHpIvIiSRUZDqT5EwOjKggXfsBl9ixN4I3g3Tfg02ePpDTgTaQ+yTJazSlP
cqDD7sWQ8qUWm16qOUQPn19hVCIn/vQoVhsqOKbbYPA=
`protect END_PROTECTED
