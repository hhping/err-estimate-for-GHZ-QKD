`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xEMU49oue0GdK4xAh3ydUPoA/Pw0OOML396MsDTQkhKAOfoWXH5t0ytAZxBHPmbG
oLDwMBNtvEnlxaKlWM3VP+1S+fYtAUgGj6uXudx9YG+AxntsZoBPE+sr7rb8ignh
/cWN4bFpft4DjMfSo4bT/VNy0VkXnI/kbJujrhhj+8AKGY893HBSzqeztS4CuTKf
Q3Z7balyfMHUFLPPBnaKCyjbxSuO+j7DpTo5hyBoMkE7G3GOsEpIyiH0Rg1+4pSP
ntRyvQScAien71CQv6pJekGVj2USgJVFq5qIluC8QZnPmgMm6hHX+Kd0TBrBihNe
4HrOyI6Q6C7N36g0jR2UZe9+v3F9a6gPtyiXQQ6nAK893QB7hCzqemNy2bj3GXPz
naZ1U8Rw2X2zvg+wjVqxZmO9zKD+L3Rwxw9rkvq9VUeF99ZT1WquDyObef8WNtiw
rxh+hmqLagIr+kqYgWEGZibZHqiS9aOvfOTt7aMG4RO37+pImGtp8XlDtbM/7tzI
IziG8rDBtqWDuF0Fh9nD3dwslmPFRKXON0Qw90M1H7ieYcWy6IYJExnLQNA9qnZw
DTRjOAc0OCtFeD7uLHv0yHRSoUrz/6eXW8NyPDicduVODM5/KMn6qLExG7XlgQYB
0+mUBLWG0wzvVyG032gQJx9MbhceJ4W/dyAXkIStGus3p7GInxC0dWDmJnOPCnpe
sP698VCUaBAgQhSaRUtIu6+Ug4KyFPwc3XY2B/gkGGuAl4xkPVO/us5gB3URdEmL
P0PuklPrrP7/pvVStREA1p8uyNntUhdtnLF0ZzbxrdrplSb3FiRhm14vjz13kp4n
0gN/0BYFx5xmkS1YZGTk6aXyPUnR3GeRJq2BMNfOs1t5TgKGIIITwDoNNNe2ah9q
KivKUd9xnanz7b+w2/75qC/HKVaDRvM0PSC456M/lmVPtoYiETaeyl5IhpzO/nXC
o+KYnC+p6LccpRXAlslKhITR1L8PWxtf4GbG9NVdbSbGIBh6H7LodZwkkcKtWH5M
87jq4X1P+D3dSpolaVOjWRflpJxISsw1KF3rLtbV2MhLNNsSBSPkYVcJYs5p3mbH
7IzbyBwpKCay8mVW8rMsJQ3yxsTjNpeGWTpfiF0gJS9tgMqO+9jR9CUWfDI0rzHM
obsXrMwn5xZmLkKmX6ZiIm15q/wjDQxYbtB5+niDi2d5T+G/YDnJcwdQ5Lj+98ci
ukqbJIWLTdeFTfbxNZV+VSFrDKg1NSS4vEHsHbTxA3JThh7YaOgFTRe0Y08zFeG+
6zQe7SZFrpEfn18XlRYoCi+zLxN3YVPqdYODRqCbjXTDboIPd6zhI+sFumvmmD3p
gh5o9tlue33l2z4vuxzqn5+YVOoXG/8K7BSROp/Tx0MQe4AB8NH6aNFTE/6Vd3oh
0Pi3cShUNrpCdeozx6WCkxvf5K/4wDImbkyV6O7CRWbkXS+wLRAC9Ka1AjyKC3AH
AcdKYxXCI6J39TH/xRsUibxiTKBpPALa9l1gppkXwXGTjvBd+TPIlz75QW/BPkrE
M9xzcYQIZTGPBBxnz8xz8GxjMl9ZM7ojWqGivMP81B6jcmKFcNULmb9AFod1WQlt
UO4UXvDIQ45Jv3ZiXNxu23j04cVrMEYMNsgGg3vvgdCPkCS3B0lRowOX4gjzEb+G
u8ozu+Z1z1Q9FG5Dw//v/c++37uRI1JP0dXVfmn+F7zuFW2tJoHY7U3vI3S8mgjY
1uKfxVKoBer+00qwTuMr8lY6hM63tRLHHPCYNjWMYaBTZtS8C0AJDTklQNLTvknW
NLu8dy4ics6+d+oeTObagSDOOLp3t2kHeL29Efe7n/NyOwQtdizFx4el5nYluKvZ
gK5H8QYewF7wgH5cySw2oMESAFHL12CY9gRr9KkRI0GdrICBI/2WOqZVQsRxxteW
GvHLBt8AZLXJ7ET5kZuJAGum8EDqo88+e3aimXjMxfScRlvgFpI7LzdtGCxtfIPE
YdFzAHrnLRDah86Ce6CpmsrxR840lvh4Y1NkoRNdjZB8NPGzXDmlPhD9ncxKOzze
K/aVFVjH5MRzD1WRl3gUQF+kLnDwGQpCPaHLsXYn5s/5pAMlr8XwTd3856z5szCX
nzSPY1dlUUBSBAC+DwYYASikrhDKK5oyBjxkDADMi12fLI51m565mHAMDO7JJRWi
zu8PHqzTsXfB76FfOP4tprUbbOrEBOfAxHtUsJh5l8QR7kY/yBnhRAjTf4Qxw4HJ
Oojpvrnptr8SEvO5opc4X4yrpOvYtFNnmQTRnaAlrUFtAj2e2AV3m0uH/cdwGLF9
dwgATiB4KveKyAaBAdAAxhV/tBpamGD2/yK8OzpDCzAj6wVwnlClaDlCpbyto4Kt
1HWewIHZBx4JXXBKfhVr5KU0YxOqZSi/1U/377p0h9wsMA6PiYP1X7XZF2DKypO4
XIiAGT2FB38RmAqaVOSpqT/295GrPmjphPmPRL3r8zpZJDyGL4YL21vMa956B8ic
wPzSd3q5OC8+Y6nex5fjev0Fck7zUODroHhjv70J16DGqcWOd1OlIQdBPbxrCiCR
eTpr0NCMh4h9T0R2dQlLpfN/KpGQeE84pTDpimXyX81qYy8Ee5XA6TKS0uZvk0DN
B++sOgPL7LnD4fRJiBmM6e2dpDMRLlYpSRHiEBYrLxhrG1T2CHUgVtmNU2FCHutT
NLe8BB2Ppm+L9iKIjC+YDAqv2NgrNFJBw84aMXwtFDCkF8zn/x/O47zUcBV45BIJ
iCh5Nb/BAaHa1B1ZCFBKWoajmfWj8U9qSqFJNFluGXNEtMs9wnM9/lNA33azJNlt
jEXOquJjJ6r8gu+su9HJgOER+dDQUXRZl0pbeN+R+r3EpXtY8l+0jFy3ulRPlYQm
gz42pS4a2Nl3oovuT1twMzIHqgPmyCbbIMlSPxJ05r2nZmOhEbcHLI4pt/YSQbje
FP3p2KFCZDE8emx/uGvT/GfEmsmgZtBcOVUQiM/wCg886ynhdpKtvDZCjiASGPXu
Hs28cR3nd0qmHSeNBKasQDLcUWTBz4LPCX1Inbhom1HcstChv7X/oqNv1xU57PTI
+CeffsaIcUYtkwsm5FQDLLJ5FM9USa8x1zKt9U/2+qXeHBLWaVPfDrRyjl3DGeU9
SzeML4kCoxiJf4Wquxf65yaUBzEMiut9zbjcREDb0dkSMC5ya+KjrIvtDCL9rOn+
1VHmr+C+t69e+Jssy2ugFalXDlE/LaFWuYHkKm4xkaHyYspfD0uCjlc9/QL1TuE+
yKLzXsKh+HD0cfBZQWgKnw/k1akxjMJ3aq3dkIt9MxaaMxwyU8CHOLs0AYWaT/Cq
X5+e8aNARdZmr7LTce8fmPUKkNqzttFw5YfZ+20qcht1aOsj66vSE8Kz7NTPHCQG
b5h+nBFO4FFRxsnvCQwrp+eppYU/GFJeaWJ8ai8tRsyhN67woNlH74baxp6v+F15
uiGJP0A4tbv55CqSLHXd4qCgsFX/00oIJDZ9zK1tN8dB/lhjhu3lcWcKtb7gtPby
C/VgKv5qGxGWGc6f2cPWQQ+6/1GqX6eK0nid1Vn6RVsANO/Hc1n3u86DjoNNeXsu
66YUOT6JJ/W6Zrra7LtW3hLqQrHLsSUVoZOSHNBTkJMdw3RyDPoOA+HOHDTiK+l/
saFee4DGeZWupjLop3tosgBzd5jMudBBusz+obQ+vAqvPTpTrvBGxKVnw5L7T0gW
sBOAoqvbbGuQSvjlkxHxCHC3WbPRCGhC5ye6E0UdpOAgKGZ8LqXlzgLLGRlKFRtq
amJS/QKxBTy+vQtMmc+upelL8XUj1kJ7HHZ9JHuwFTfD8nsv3PnbdqTDf/MuViDP
AgF7obqVUMePHREhNUEmmzKwSn72u5utUON7+W0sGGGRyNLP1rGJ4fH6AjRAWkXj
SDPH5qMv8phQnBUfflsNWkdBp++y+SachP1KdtBcvaCS2DkdT7+dZZl/31tu4gP+
fGsCQDS00LuNX+cOw1bvy943lW5IGN+oypAtmbcr2LQjGalSiMQL4WvCeiqvphxk
7hrf0M4QEj/52bZtDVhL9TlAwI7u4/rwzwtl7zadkGzxaIMEIZrOESUZaisUkGO/
Ro1o65HFyhSfk6qXG7b6JbiKvCKIRekO5XSNuoszINAcj2fMjl7caYKwGN+IHvMA
HohJIq0+zeQXSwixlbia75lAf/2fD8D3C5kBd0HN3gvucP0YWGFTNJ7Mlc1YZHsR
+NvqYKWWeiiblwXNmxrr62Pq5pBbWMGNVyYeX8d4fTnYrzIICCdaf9kP7LwnfntE
KuZ2MdhRMZx45MYetlc7N+AuEUHio7mct8FuBUIommrChGCpf1xor4/WROIfvdvX
AVnjZaG/0BzrlWmuzYMJaV0p31x0fTVx2HoG9Zu4LZpDpSOdUVj2H+rMkiFHfx26
2yuWvuGc+sZyXSGoTnApG6V2cZU7Xt+FXztjaacA2QdtnD4/mFa+clNpL4PFyrHY
zNrpdvV3INMAK04/xSEZSh8B/3N96rzWc6WOYdoNaalqfYS5RHA6p+4ejk6teIU/
tjMxo0oVyYEkQxCyjUZZob8JIC+78B5O0QEjoMGwekOyPtwhojscITtyLzlC+Nm1
vh7WSFYHzBqKDCmnJfFesEl/FGvB7lwUExTJsL3t6kfJu9tndRB6zPbLf5EsSGkd
YAw84dInIw7ITPJL+j85woVZ2vzLn3dKwlp0ztNdeO3VNqGDXTOazS894aHvOHB1
2EdG8RSmkekxVDy7lCCo+7bcDe9S6SYngRKg6T7kk5r3E+IYcfZQtNdvViH2sjwf
LstGL8ctjLFdQxSrY6Qui6RMnJ2Lp8DXvd41BFICkb7gsMuDw/uqT+e2BMALDI8N
rlV/PraRLEa4y1FprBEqBjveVXBCJ7QQAmFCHrw+3RNDcmKsXpebYNApvOZm8HRk
0ANue1x5LyTQEgxU1Flo6ce93B+fy31B1vcyywKsHnAL6ddOoXhYyUlP49Wgpvbn
WHzFdDM2qoWIx1w+y7f7DYrLMQmYq3pTwNKRsJjacc1Sr8q2qbGO3nd7hRUU904u
/wrXbvo7nfZYxSjW+a3ab7HegaUOY/jZz7rEv2orVUzaKc7jizSxfqTePtC0vlic
XdX+YV0m2M7F5d+LziWaMZ/n1fVgIJCYalXR89Kq4NQKOXMhmWCX4SZ27u59/VB2
YyM0PQACPTZhcX7aeUIvMGFsGkg/msxcR5d4GkgYAtb7KJWlatByrUmNSQerFkOo
fMkW1senz7g1L+6Uw5s1r30mNAX1Do9zRhC0soebxRg+QHMVFq7eoS5AHdmG5PTB
CFyvFEDfBBrQ3lpxwpsZmfXCmcE3mCamFfXlLLuEuJkGNyyaWfw2wWk6jVWvYEfD
+fQt/S9eZkI01/IrNWGH6uzLS8AWGClmLwbMfuP62DPOGpNd8JVdzU7h3/f+QanZ
+nZvEizw3oLSitjsWdoy3KabUH61TOk+9lj2AfzLtzY2330osjp5m3yBMLiUh5m+
4lBNz9/bl0GAS/phrMiT20ooJ2p2Nn03zdpKuagYczvwQDwZQF+Y/MGP25b0ILgn
i5rkXLUvULe0bvxxTuy2VwnjRvdpPKhdbUhShupogk/xnAYh6zTI58/PogJRtqHd
5lJVPLt4VCO/e78InvfOb8XTidCV6Dws9xbcKNhlgVcCiCOwpmKI0bvIm4egxjZl
gCTP0FIo/tdCoTKRO5Iyhm7F2Bn+EYRAvpp6i2tfAcl0gqg+ihGjBqRyF1UF/KHw
hJakP4HaAlaHoMmbBuIWc5PdXgr5KqKalpnIu4MZco9zK0JL11197ZzNmyJ9Ptg9
SWLmkFTyQvl0dli74XOkY3NNqHEvqZUvJz7Se94TulLFyFU5AAwubup69MJQO9N1
t4pDMhIPfcgibqEbtfR7TPBJikRCJIAipM/TcbXytCXmqAhWADlQRNWl3w50DP9Z
l+0XXPcGC6CmZaFYiRYeAvZyx8fJJ+SXVF8P73C31bsu8sj4RrT2jkHQaHVRPYOr
5/F8VJv0TGziPvnHWSkV051QUj8QOASZBmUh0lh4Ajd4pVOdwzOFkDMgH1WxwBWl
gD7dgGzyMEKJA+K9z/ZAeRCaZcVcRBlODVrqQ6Nco9wYr5vHkIhR1RNr+ZSdfO7/
ZrdulBz+xx/ysO68LqYMh7CIW6uM0vsIF+8iEtfAK3tCOSFUGhFs209eBTT9TA1b
r4iTBS2xDv9xk1LNBdfNDEA8q1ae2U1QYFtUst27dNzEcFTA3C0/bKabW87JhBwk
Qn5f6CQks9E2BSwGpR6l0iRKcXF/p2e/NLAQuN7iEYZEdDEcyPrHTRWCFOjllqQq
OcctdYY5fB3R4BwGruJ4DFBn7MxTUIbmcDiBEtn9B0rJhpKhp1b4SDZRAnhYd4pm
Mr88Z5ZtQLJv/nWinHg7O3QezcSUv/6tcUGBbsRW3iekxjOr/sRFFzO9fFjyA+uE
hl6DFjz6GPAP1OJBCBH5rQ==
`protect END_PROTECTED
