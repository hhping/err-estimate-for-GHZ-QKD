`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u8BJDtOK6TC2xovVCiL0CMyrp8VmKgK3OQTDtGm/CQnb2NhN57Huky001lzKAeAK
lnkV5u+RhjL1EsrP44wp4ThKB6vxAfJXh0s4XLF8Xhveis/uiUlBSdPk9vlv58FF
Ya77e44wWRCHR267hRfZbrJXmR15K/dCn8O3isKDs1K+5I7Cy9rRHID01NpzxAes
x/CDqb9wWa6KbhzGOwy63Ybzft8LebrdDeiVfZB702aJHr3tjgYnCqzgsdc2n8DQ
KDxbT6pyRcj2gBElcZiXsfjg1v47GsKyDXGNZZA7JBphmDIWN0tnvgwdV8YFqbvG
zKZAwdLnXVejCEtP33fnubuV3p9HdXPhHE0BZlE4oIrQVqjy1hCidUJ6sbdQawRg
wCtqnz44Stb/k35X3qZ3dJgv82vppUPrRsDcM+mr/7Lns+dI9kaMBoVS4DoLOaIg
vLAfCfz5mXRY2YjJl+xKm1sP9iSi4cLg8KOMQ4WRu26XROxpz83e38MEJiuf3jlx
NCMm0THbLiv+/+/UiMZAOPT6biuUxOWlS/ehK6QWUW5vx4IEB/SvNVPvpKaptWF2
3w2pximSn4eKoeaQR9xuGLNfTKTtX47qRSv+xZp8qvwQd+ttB+pm8y51p1tJr6DN
MKOcksbRCkLWmn+QfNmcu7Q/K1uajRzGzFuc+OzhFWnDFzZJRavmuy1qA8SH0EDu
JfJLwLx/taSpllOj7oFz+wFGyojGJx6uqNPJxVSj3ijflg++MKo2FxzthKr6BvcG
5koEVaundbTdvXjWOAqRNAp49rpO3ff1jQeOmjt7JMCyI9HVO6pCsh4wBmPnBGUI
b8SNkVE2C8i2qNivxchES2xwvX9nX1+Mp21nKwUTOpQ=
`protect END_PROTECTED
