`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JcqS+lLYyqy6b85gZuiPhkz9ptJNitLknAClKC4WYgDIzHv5PRz28dsiu6JEGKLN
/YvzM1O8EH1YmCXAhg/iYovxgYIaB7MOK2EMeuC5JzHizst0KCxigPsz2vDdl9fe
s8ukidsn4i0UM1uLCTugB7QRekEy8ePLTcZgDm3h27M0YlcrKMTj5PQXORMzxb1U
s9hzRvaZWwaFqEa1Z6bLiTOag8/2/GsX9vT1DPLTl8Z0W3yqg2BARSMsTElsTZgH
cicqukmULii6eXGHx+6fjMQMby/jHI3dsR2C7MN5BXlggrfr8I6dakcaXu/C21Mn
KLiZGgTrWuO3fYXwg7xs+ogtoEEQ51w87CPpnAwTbZQ=
`protect END_PROTECTED
