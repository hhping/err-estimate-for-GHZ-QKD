`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cpo6UMKtMujgGTDu0e86tjTYK8bsdDKIGr+aUQjTr3rCe6XBueCsiBx741dNtHPw
HbMoMFYfT2PFDKLSINojRdnT1SSaBuNk3SEMmVHFf1YhRSodJ6sU4qm4XK2Tn02Z
36lZ9J+1lKw2CrL9nZhb2fkvR7gy66L/6R0ZA6X4VuPGBFA2SxOiOBFF9ChgV1N4
aV7JKRQYMDZGuYnZFkxhjfRsWQkdYKVcROWCMVqyRECuQA4JA9jDVtbnQseXMCR/
EQ0WUiqMXmbYPayiud8L8fPzA5Ivewqzt/FNTQfemzGmoBMcCA3ksrrPUzNRJQ6a
QmWRUHybp1GUQczA2CCtUIg09uuLA5aMhBukLbzA/HbovtNYfnT8mT+/R7oT/E7t
1Q9plzH+kjSTcn0V01HMJyYeVRWZyoEIGlcryZcLqCB2D2h6nzWyVX4nSBt0EeT8
/lDw8ZsHiw9PFSR9B9KKBjeHLNBQjLCCtTCj90GPIOBGqzap851BVlWw2Tu6mCm+
fml7anodWN/GOWb2faF31ZdiXaAMY11nb/idQDVY8OkdhNNy4MEWqScMcHSbf5tI
IyrWxnwCRXdDrksQSblxUBdGipaRf/aoy7k0z1Wbn8DLM39b5JxhfVCUKX2rLfHu
u4bCNNvX4fSZ7msI2CzTqxpzRXsnbUm9ojmFfDzCxB2m9havVCIIO2NZ1I7nytOH
Snn+aLSunn+9CWWFq8/cVjRq6Oq7H9tbZ5hiCeisNKoQCDMX3P7EATpfzLJbrnkd
/lwNQ0SsZ+DhNWGb0Eg2VnaUztR751DlDRPF05V5DA1J9aeQEOedtBYoxhkYfdSI
kLnmKNK9jA2TysoVF1LOffu814lJmsA84QoK7gZrMKbq8dCTrimIEyqgikZ2nZtX
1GKEX5O4dfRZff3/G1Gnv6h8hlKttSMm74ZPZwraYDTvk6JFZ36ql5fga+br+BcK
loGbGSf1Q0EE3Ejn+FtgacJ1bMKvMb3hitqXj0Y4KYnFPYsKCOrA2sh4AR7nAJdu
L0nXp9fDpiZNGyu3sOQy7XhS8spT813P2/FGKrmHk3UGB01LC8ljab1vy2SPvA3t
PQ7FXdYDYX0besd1LEwPlo4SrKvNzSBdO/W9bO6g9nKRvMyvDHgfm02cJ2cYd6sd
4zVBs2U6rxsfeQAYHiuR6Sfg1aGK0Yhp3aLuWprTtk4tSQSHHTmrRSbP8Z6EPQ0U
LIOYtPvs17cVb2I5DiDHw+bwzT8K/7XYmTQxIuXJhlmQ6Bhi0rLVlRX6wLzKoDhd
PYVgPCjI9MI1zxmBRIhUiPM5/6GwoxuREYmv0wAzWxAJsxWChpyQe7/hWBqMGc9D
b0ZsN4WIbKgRxGGiFkejT24/79djpGPHdO2H6Nc0xXWrbNnTqvzsTQkfeEt6xRSC
wdgSNejSveLSTWcpHgz6udaIkGrOGLOwdVEDhM5Z+Q45IH9CyiA4kf4Kjo/1XLp/
IzWND9a9XqidcFgV+MR+UXI1tXXCBSB7Pzu1BZfUwY73pzVqt5DMEk+SJ+eOexkF
iabUScrn7vRLkI3h2+CXqzeI0bFFHDOCXuPf3Bfr+ha3WXrA5NHoRG34FLKwQX+k
kr4APiYygUNoxVFrhTBP6rzZhNj96G9Up0jlrBRgOLWj9aKbIuWHw5gs9vECzH0P
G23B67FNRTmAP/7FmC0GArInrULeGdoZOR0979snFIJWFmORb2B7hHzjdAU/Z00r
0eSNKeHQyDxylUVgxQ6d0dXqweOzGw8f/7N9DXzEEtQ=
`protect END_PROTECTED
