`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zGh16v+p0OpXSrJ85rz/6vZMRVwMpWcqo4BoKofz+vRu2qB61ReKBfmmPe/lvmmz
uJs+gIZJIRA+/of2MEJoAmBLBiflTBv6qKkt+0xXJmTBf6fPdMLlTHN3DBr+24ZE
NhF2CMLELQc6lMO3odt+XwH4nfQb1XQbggfaphJEx/OqBU17YfzS+1l9QLa+PYeM
Cz7vewovCbwMNWgcfdXBFYUs1I2OKzAIE4WRayyhcMDzFM7ls1N2YX6oAfQUpbTo
GolTK6+H4hBIZPesEIOvcEj+ZNiqG8c3lVXmUYpf7MuSZpNkoe59WFYG2pZRGvse
5b1GJiKv4hGLXOzR32JsMmBthgAhbQRnTyKSdmQ8fVcuxHuQ4Xv4y7tFEj/bWZin
THrKT2urcZXclBzNMgAIbYS3SJYUYMqkfBl4YG/OMGRyKX33WUkp5sP3phLjnR84
xq8jYyhuLPnk4kEAv1CFOTQlZLHei4Mqy5HgtwcKlfUXPMR4z3tNRDsc73j5s6lq
a39rjXtBU6jwXFvPa7gy9dysnvm6iJzMUc5cokp9lhFfn7fj3nYMYvDopeN4XNQ2
arfG5SZ8MEJbK9ZIxKrSLorHLn7Eoc88JR/tfRdUJV1Ev6VMEViZEk6ciAb2vXvQ
QCYhiQJW5e4raW7BrzEk48EtyOf34FNC4L0fWre4fv43S2A25M0e/Uv+jjWqMZle
TNCmTeHezyasD1fWRBfy8ydIb2Hd2mPcjPRhMEb44V042icJxjxAU3xGnWrJ1PHS
DbgZLeH4OHyTS0J2yHiylc9Lrkwi0ZoBqzLgVaph94S5ypkh3FS6oPnRA4IKLFMr
ES0B1yW58/nc+/ymDNMDxZjxqgLA7jZ/FKtsGa4ruXXjWXGGGkqVQ/U1VxOLhWBg
ECVEigFagERKFiQwojbGsPX3sbi4SLwM2QDNKDErdtJJO9q3+RtMbCl7+LRPI7g6
MkYujOBARf+uKI/N2ioyn7YLgixgDAfwz6JZD/NquH8=
`protect END_PROTECTED
