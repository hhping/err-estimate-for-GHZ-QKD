`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qlX1dtgbT0sWEm35nCdFlqM8oitTGARW0lJBE2lLOouEJ8YxWboLT3pyjSXBfySW
6Jf0IkouAhmsSCUlDTuR23YZibPRrRQlJ7YGuDIdXPEGBXrWxxuqjJs+pVfkw2Zz
uArdH24yYefvTLBU06uaFKaB07e6ntza/F3fWMWSoqrc9ysk+keJeI4UBVIXn20B
vwjP7OqOhcSZimAdQg97vsZRGYe5RwqE+2BEqviqvexroFngnVO8Bwyhnij/vNrg
0Bk95MWkXvJiK+Qpo+DZvfvyA8ogovnj4/gfKTVCu37qpfVhmNILdfQ4JgLyooyh
kIjX8u14ewTreRqq7/Vdf9/66E5TRKjd9S9Wsr/Q8rqIpSL4ts9YdweWAaGppw7K
XxewAEzwLpCD7xGMbuXMeEpbhYYJvrPqUHLGMbgpw4CZTUMqmVwB668nJzaxBmQU
RvcLVIXFBl+02BkOe93y2/04iAaujxUrAEuU5aG+cCxZ1VpAx2u/FWO4Owqsi2ia
x8O7qPXDxWTVI/hD8dmm+2eW/9jwrbUBn+htRpZvxuVzxMu3qP8XIANS4XeP4xS2
RH8lO/QSRQv37sCIKS+AZekIUi8r57LchdsiT1BK+8wsWgakW8EOklbnQhMGqE8P
49X0NtxEXFfDSmX/f59D1slVtChfPxE4Ds36n7Omz9ePQmHafDkhnJdtt4sdmrfX
X0Gh+zoZG/P41CKdnS5zxMUVJBha8+4wDy55xK9EGNfRJDR8a78E6FYQkXCC/U41
os+KGDqL0pv5P6ln9NFyLUBpgE/d5bTMK2pWg2RyHw/TVe5ju/WTfd+vhFRYc1QC
b8Sa9LgukfvjUAWP9kklchBCXuLvGvevzHH3dry2rhf0yca+cbHhQ+CZNqERlOb7
SCJ8n+Z8tboZzTANwdR8grvp69tAerGEbFmb4fnszvTt8KZDDf/Ql6zb6AcJ8NaU
k1Duueheo6/oV6o+wJJvlwVlfQ1DPQHBkA+cbmOBtEiPEFAPfOSZsfkSX5L0mXyu
YPX7l5Y06O5JBCcaJQZuoLOjIcyeYwwVuT8IB4APyI+dw1T4M0gqfoOxODTAML6z
daVurfHl2wWnV/ptfH3Ov8aRdnzOnHANyOUBJVjDsfio/fJCDLS5JqJ9R26GvLhw
+i1klha9P/FJkVu+wL/63grZU26BJ1o0AYT73Xk2TwIUnRJJzFA5QF9Hf1+UFq6J
JHEGaAd48toCcVGA9OqFEdiWrITcbkmVNOBgz3JrGO7kxzcWWHZMHMMhW31R+Gim
v7PuKRyOkriHn3UhCxPGa81C16J7/JpBJ1QMWw51k4htG8yhoftOAomUIt0/6qm+
uLAqxJj97enAFUtLsaYlzNGIDJx/tYQXzBL9199GGfK6Y5ozITlVovw0OKePNbYu
oppUNtnFZfKOfeUjHfin72NAilEv8NHzzegWb9JgJCxP1QqYLv2oSiUU7QH9mviR
gqw6oTJexWaNGXzGHDQd6BtczDEKbQSqzxtbCZipNSO3BxzaMEhm71zMFQrKikIa
7p5a9Bl5lok/x28XgFUndxayZ2CJZI+pOUKkhsYOOlXVrdaPcRF8x9l+h7821H+n
pEdz8mNTeP/56tmgNkTSYiYhcz9kqd0/D03jox5ibIoW+snZeoAzZ1nRJM/aHXvP
XMbsoqrYBewYaYRTio0MNaNTr/4prsjX5gPE/s5tSyXg1eFrXMnPyTxIxrgddJRn
azJ6vtR52KM9QIYoZQuEjjv3NaGLkn3rdd31V4TR83s/w6y9axWVkIFbQ6pRBKGQ
iyJf6ehNozIlWh0oc7ECbHub4+f3m9puKyBp0Wjw22PI2JLNduGF2o4Fcf31tR3R
pmIDyrReZPpn8KFlMA4dlpvVjbRnC2GW4Ax/LTpNESm+Cht5R7JQqvaeBlSn6Cfq
x5yqWrjOAEwPvcY1/ElUY7mZOuxQtSn4AttJFiGLVXBVMYabMgnLayZfVefHPNgk
5MRF02dTX8z5kjmPjLGDkXreCtLJN9WLCGkIbcgfFVfvdHkQvPrFFGVFz2FjSlrx
YNMHWY1B8C+VsRkElRjsCxFWt+iOr47fY9DLbXmB+F9vAOSH0rYVyWyzVRrWi7U5
uYrMw18giWUVSnX78jCKFaB2jH27Fc47L4qOe0ShGZ2quv3RW9kjD/HFP6goueL1
pD6ecoXPYLTBbTvvPsGEqmTxvU4TOff52ZdpVf0CUaYmUwnzvb8TnLJ+yuQ4ZZek
s/5r4ZlezB540FvnGBHeG9NZH1KUMsoWV5Qfy1tujsLz0iOt/6+vhVAVsCMKZg7L
wAaT6Ze/AiKVqfEkEiglBHG9RIDrtPgnPw1u33CY6Jd6BBqtgA4q6zSNAPr2lr8o
7YjFcnUq242GlLXUEtolhag0M7DMKc1soJUxcj7o+8G3xRH9AImpBdiFO+DDZ/cQ
zFNxbuZSJnxStDtYvjeRfhOvf2Qn88mBOCpBMLRk3HaZy0FW/XprmoP4en+KmMFV
WAIo2lopr/VpTIX94Ua7Uapslb8N4bTIHW580e8VTM5wy54gQDQkNr0Ob1jvdPA7
8eW/N82kvTWnom4bhnlwrg==
`protect END_PROTECTED
