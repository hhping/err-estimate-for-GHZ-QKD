`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3Fo3S7V2Tqpx9VL+lvM5QeqSRsvL0nDLlWGH8pPGLCjVhF71J2n6yC96FrpMYaEN
/imLJ8g19ONnRDlWR96ZCQsdeepgSal/vPdZR+F9+otRvytXuKPrdGg78tT3u+hX
ygkhEBzdQ26SdQXKRQTEauO5RyyKZcPyk7yrdUdNxf/Haup8ft78XxtOiDlihcCg
SnzUHlpZrkZ8b+Bg9IwRMjO9zgqlLRIjlSMF7AMNNY8bo1PfwN55p3QJkMMop8YF
MRkasiDWVrE8akNrG0mDZzFKyu93jaPmpeyNd7BPERH/Bj/ZG9GeNl/stlBpLYLZ
REGYzr91wt9gXmT7IEtgHGvR8qOrWdm/I7uVpHlsGBiq//paBKsFD0ByUQlfdDCa
n4JE7tsAkX7YaeeREUpzBcgpHqBE+SjMU/SFRwFx0FElhPW1VIhbBL4b4RwHqzvs
jNg4RybeRz+kLMLhhkld/KMXaU3v7naxR3inRj9xiBCImZh/IDRBQ14jxklDjocv
tarA6S1ezILaKjMECnfOf6PkRnOuuDLg14v8Ze3A6SdgFadWJNEzNKnjKizVzjaV
p7TegUZgLW+NnyCL+Xo0AlgMSs0TjvW5Jo+3mYrk70JPgcTrZzIZ0jzKlNnaag42
WR9oBUECX3mzLtb0vlsKPIGXCzq8kf6MkZMWdVsuf9ynwnD6peKSaY3nzzZfrs0h
6Aynh2b+lOvkP/WunWww3PLNK5LOko3+9vWJbrOOJqCBHr8VnwJoGkTUO4QEUEHY
`protect END_PROTECTED
