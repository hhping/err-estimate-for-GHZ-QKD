`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zaUBWz64aFExwLH5EvTT6Am3bAJo0AxWiIkZbvIe7qf007/639O55qLNnBEwGW3A
VKlVa2N0XHm6/qf/d9+pPzGLl45ZFkU1zTxdIpinxzAFMGadgO6T4CLGSK/L1fMF
R70M8ShoUF7fxaYkRRK4yqwdaOxQ6473tWgWLxF5AcvjxV7Q6RHUJ1qxXORZkfeT
naWn8GwPQ86jLPnGQYZ5sGQ3UMjzdSWSKiLL/atI5WwlytJh/Vy+Z72/pZViQ8eX
ddr22952DY+BcRE3e0LklaApK7DBmIIhqtqG9UQNtr1CaZDFylcyV6KuHyuT/bGh
3VQx9mPk4WluZEehREp6emBivHrlhQDxiy58Z6GB0/F4vi2CvVM7KLcd65HPaJds
qQ/SWSyOIauf7Sab5tFBL0RBDJx9sG8JSkPA3dpLd5Qa4fczWmzD5KzFUVuAI2qD
gvdA5g5ciO4Z3Q9wIOwbHpVuSJplpH9GxHqBN9xpUoJl7I8SHrwA+2qXT7rm+6c9
16Ynon1yyiolw0h5DWIXv2+xLWT1nxt5DulFa8687bY=
`protect END_PROTECTED
