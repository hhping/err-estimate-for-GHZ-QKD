`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z8tBHKPcBYXpsA+kdgf27KXO2sYiRuqPJF+1EFf8CqD4HQ4CAHvjCB4e6DLYyRK9
Tm1JN6LeGWEXchDbfyx3U1XSmj+ig1DCWMaOZSafMwST/KeCeqGtAk50vTk4xBZh
9LsRIY0wKRflS8YAFGqkoIWDkidMcZhI3EbHivPzVLSNEMnHcPM6d5RR8DBHEMQ7
3LygxZdvKC0GRDv/Jh1q3PTpXptfs6gf3Pe2Spqlf8b/ifLWw46Ep6Qanvmcb5p4
NlePx9CgMBlyYH/d/grGzLJtCABMxLIRUmjy/mVyHjVLvRac2i8ARo+gjaRSrZzC
zwKXwPVSYjuuQ1dZkH73NsJP0jAclFKKDu4vssEptXcekQd2ByTjDQf6hxOY27OJ
Fgd4ZQf2bFJiLgaINQUL5rEFLXKA8Ss/RDRc4xYFGE3hUN5tXCoc6qD66ycG+Mwk
MmWzWYG2UJvzDFmTPmOWADs5yukNGV7y5UtyBil1dWGUdZag29DmtYNvmjgKkSnX
34Xs/iDlOynRVNb4TbDHO1qTWIAabdc03Le2jQL0ehM=
`protect END_PROTECTED
