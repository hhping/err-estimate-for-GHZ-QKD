`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AxG80f4DUylGZ6rDhqr6et/8Qx5P8SUmypNpKstJusly8DIYXv7HraU37GE+g7mE
LffCNh1v7C4J260fVB7H49HAbcESHWtqW4W8F2p8fagC0wrfHIbahflHGZDtWNRm
QL70LXHY5KeO10lHAEnrqWEg5xAge+RmfBFMqpSJN7Po/0NLWXubzFi0kTkMiZz3
wpZpXQ5TqMQDEb/wzgN0jlb9nEaWp9vi9xdUDg5g+UZSeAYwac/IbjdOXuf1Gqg3
8QuikRZmc43E93ahLvqoIw/h2dOI86NY4eHkZ++cgkyWhGfRkrmEIY41pIJmdHWB
reCOLcU5m2OtwkiHLXINfQk+xSfwbPgBGsUE/tGlhxkCoZmxLRcbCST6yMpf7igM
fvTeFHHk2Dc8YGp4lJYegJTFSJksZqeklfU5KC2gQIU5Kttz+tta192OIauShs9D
yb1ZENVW+m1kDuGl56i6kKQn4uZ/UFuYztdaY3CFnCg=
`protect END_PROTECTED
