`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VC9hwbmtxpkAAAy/t2p9Vnyz8+tg3cnLQC+J2AnWO8xXDDofvhCnA+KnbYfCgosi
tRE4Y23kSHG9k2MUbQ4YFSfcwcPLXhVTBXwN7XPRSQR+3B+EzUHktYiN4xujNqed
tM4sBIPsVGm13qX6qWAwpJtZ9uC42KTmFUxhWzPbAL8bnOP2NDbc6NZA1wAH7wXf
lgPybPf5YCdqYPP7NfdjoI3+FHCjq2IqpKHqhDmngYY3NMwEEOF9n0UmSHvx1bKx
Sl/Ily+S7ZkREnNgj9Y+p54htftYWRAwTd8PQQlHqXNAHF1wQ8qD8+BFKZUtT0JP
SZTBV4t8VK+biO+h7iIEAoTnGVbg2wzGNS7Me2W8+p+pIShP3hKUe/LPul3+3HzI
huXqrPhCD2mUJkpU5nH4xZhoB72yXsdZ8+CzR2Y2fbPHBeu/mNc6Ys8IBePw8Lsl
spA8OTfml3q+pY4/AghCSRsOypNocdid7xq9Cyu8Y/atF1M/iIDiul8+NvamXfAM
erdV6Sikzl110dULzwJqnmsv9D3rUbUHOpVxN0Jra97wc2nF+U81vme3a3EsM4qe
En2paQkXzHdymooTsI0EwxtFwwnqeYx4KM8iq4RjTXMTAaHLleT9YJGb5kK9BCtM
hbXpU75L3c4h4UhTkFGXJAT1fT8nDfEBWveCGaQeEFJyq9nWAU1k//HAX6a9gZcV
K9bMe0ByEsjnElr+kwcrECIjlMHVGZ9d+Mpb7LkuXakS6swUWN6T3DnYJp79MMID
`protect END_PROTECTED
