`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xkgZi5v+UFJqfezqoB/OixjvlBlf5VyUevAL9Ys2h2x2cojzZ4BgUiUsRwlM1Q8q
QVFzpdAYe0AmyiIyjueoG/ZLR1fV+RSNV4B92Li+IE+O0NXOpPbG8Gls1IdiwiMj
IManpHl3pb6+w8GNQitzWX1Yb9fziuTqpcr8gWtpwGJ07LyUcjyP8TeAgk5vv2fG
UQEF/frIuoXy3DGA53ITjV1nogr9uUGF8Q++7CgD9Qi3o09pkHTTZ1iBWaWDJSNq
YOdAAGFIcZy3aRp1rOGz1iQAcEoIy3xZBHp7pN+VFtYvBZpEr3SUs2mhN+9F0xTy
dRjTYJ8f4LyxpQgQVwKlu7rQEaUIT/S/GYmJoV+nUhOtgKxyQNLWYv7w2NRjIFyK
xCIS1kzrT10SB+/AJUEncQMFF0F7icUdpODTkX37z1ZuG+HpEU4G95vJZayJpcQ6
7JBglI0bq/ev5NoZTY5OZICIWHKiaWCFVAFc+bciFC6/aqcYmf+HpZ192k8V/pAy
H1wjaVsUkV2+06xL9JIFM5SkDfV3CJtrowZy5jnP5CorAT9zCs3+h23BS7uQgQO7
I1ZZJW83YxZoKPQnJ+92MZCU1ASobzUtcvQcdVBNqM3rxEqJpwRd5aOVA993esYB
fm0gNA32Dclk1A0YXGl/EM0hHBfsES+pjq/UFICpA6E+7c10tGOGGvZFnQlJZq6v
wZsEAdd48KUC+0+Ui/yYwzg6cH+ZKLt6V3CEABbpVo3zM/9uTSWNiI1jthCmFpYu
`protect END_PROTECTED
