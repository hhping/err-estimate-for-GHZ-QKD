`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vfjH+q3QXj0khEBFtRGDImXFH1WSls97tk6DBgHkbAOeukkqiIxxeOmmQYjEW+Pd
Kp5VOcXmsvCK7TGBrsrP2BcUEJ4C/GuHiBSl9yAD4JSUR9JPEvSk17OFwzGnoLdP
Yq+IqP2jJELEq97rhbAN02H36GQUlnat+pQnmzF6DvaKhZcHkrfceTl9hXMIwnPM
iQQyf22FEPZ/ml+lTffLKDb3oDJs4x4W2DAZ7eKDkDMKA5E0GsgmcS3MI+BZ0a55
xjG53YjEqdm7UYMUuiSxSEN/rYFCouLziVomQwWpaL5szrgJsGJOV/Ub58eO3dOb
xaGaTvxn7cXtsdcDOYzpUizkGOIU0I2QIs9xVKQFjRSt1Dp8OGu5V21D7r/v3b5V
cZe0x9InTw2mR/Cw6kLMC6hliJriQUomsFAT3bRVa+UbZLb5cVdicnl46OIvPOyp
sl/56s7/bpeywUq+jhODfo3PzqD/iS0dR6/2aVPVxO9iHR24dOQxw7BtzsCNOhKc
1wDII6Cz+XcBhcGq6wPlLhPmZ/j4Z/Dy5EErj3UaEs8zpX1gqVtQozKSX8/DKgay
nbesE/70CSbJHqbMpYFhwB86YHnu+OX5e1LslADJifjkkXZkKMDX9J9cEayY+CEP
M9Pyb9KsjNa4upIk4v2NJRctZOJw+4NPetsvyx5TLEFwiL41f/zrU2TQeWItoqXS
WdAX7uZcd/AahMInJW0kUKIjGOTLr6flSvyDE5RXktr0IrYojb75dmFS1jx1qTJl
l+F2gZNrLjAXyFwLAUEAXo9cv2RR/XfMiq1ccrV3o1Xxee803N0VGub24nDqP9RP
zLghvDPQsxW+IEVnBcIzPY6HJDpfwGXq2Wy2pgyI0asMdN0M4YvhJprFWFSbiB4s
9Kt/vKVNDDE+g+acGp/S2bnmmzsQtFfoRIDFR+ReVXuAWCMztQO7WyHNJpnL3mCJ
kw8L/zT0Q3pPcvo1zRaEmztqGUY5Afudl79xygaehMvLUnTArCx/yUmJz+DGyaKp
eusKKduf+TZn5UJdFtttiukfp9toEq0MVdKLPdoSNq8+KtItgnO4Qkp7GCXmZHaB
V6KD1t2U2vUrw1W85GW1lvzrms3y/PrqrIVLrNFI/Xm/Vc4w7UGseg7ehSySjISd
rbtzoRJNsKgUCKZRasRfpyBP3lsgTJgQ05R6GZ0mMsG3Qx6leFTC5Mbjc88OkSKO
1oIiaoq2ejA0nfp18KxsA/F5TAwYOXa96ln6l5Cx+zo9I3ShqZ3Eh5y1JUc/7DM5
aQ7Mmdl6CBtdCLux4hiZSTTA+oW0Sto9FJmhiMAddhx6yBDWyCvoWzNHfsWjOa8x
7Nrluy6c4q/nq44+lJrVeDS9rOgW9xnm6o1LtfFlxzKu39cYNhiH6cc98w6wWosv
Vb9Id5Mqjv1FLM38ASryg9k2LNTFR6/U5nITU9pkUWURJCDBvYG1jo7Vm0+9OMxo
dRLKwjQJWG8kvYSc6YfJsIPixM9fD23ZVItb0rJs08chYePaY18QuLB+hJsGcnFM
wFxG0fHnEt73bpomnmNpKKatLH8SYDsRembfGDievu5Ie8MYCfPK48vLJT60pWXp
TpOTDAKCS/Tj1momOcsnfeIXaddguXEQGbDCWxKd9LBKwnEI5xtdZUq59Ey6VBK1
VWp02ZQ7wbVtDcY4MArfyTvws8e2+WNJzzlgKvfnQSlCrkSAKhSBay3KYTqEZvzH
S9eKzzNxMlCLPHjO0xzwFWI2baEhoDUNFcj0OxnpkIOuYT/CznjQl/R+MpcBIPvn
SMwyXt/SDcXblQQ/2CP0faAxOJgNGHJU43Loerhcqjkj6TODCPN8cNHHjBGSJU/A
Wt9CcOjECxfjynMWgske1Z4Mk8XOzJcib2is0hamW4JpuLsMotJxT3UG98pEKlw6
LtltZYAdP9A4MxJnRsCd/5nknaMnAFAPFU7jZVc0T8UHfruF+KKq7lF2myg8ooYx
PQVEOefV+hCIgUQmkTlCRu4XDieldso0h6sUbDffT6FXg3n2RRzsR8WNaWMElpHE
EO3ToCNIFdaOUaRX4g65Vq6RQEXAUMcZjJaDmFj4i9kD6SvEQhW3pGTzS1Yrcs4O
hIpW3JEUnUGo1bmiJwZO8G3kZ+QzAdU1DxNQNb64GOFEO2C5y2xXBHNKcA2HqCat
O7FFMNKsJzrOxM2QOvOIehju7zD8HXfSOqu43OM3bwnwrvpHSVWc1tif/Yo9cysK
V1HIbb7+DvvywuZp+lc9+oBw2sBbvRtnjhZJFNghyJ8P26ZY0K3Y2ZsF7XKQe2i9
Mabr8WYBhFErnmq1or15mlsqAwXNBhbmV5WDcKuuTJ1M5APNd0S9WWLhPrdtkjDD
bZOOvD40QerdhFe8hD2lWqSiqSIjkKuLzupeYzw3sSAWj81rvM/0Kvvk8hhinPuq
Lgx4CuFi9sXhNlobC7Q56zD3rJOaN9ZKgLCoEYJrgR5JBM/gfOlCueXj0EYXvWfI
vYQwVB3WKk5siywouVSqLp2l7wrut9x4Ab3bTs3ihc1Vn/0oXwPlyESfrK55SRTh
rx/q4J6rla9Dz9T5YfomEIusGHz+oQ3iULGgmKoRWHFm6G4EmB22avp91+sN7ohq
jJf2b74fB8lMn9+ec8rzgqCjgIqWkxfxF2vUbSCaU6UVhiGcmi8RhiNxTpaHTD+j
BN7rjMhBq+HChSfEAIsE4AaUfUQI4whjK+FrZdeAuwxhfRj2NgZXxp4ZqMLSjnrS
Rwzj/UWHagALWyHQnXVOnhg/5+UXMjk5yAMyclEv/Bhbd+yuQLssNhoY5MN3czhm
f4t2JEnI+B+2G7u7sxJLNYxEeLD6+RoIN1F77hOwec7VUTzk+y8OyS1ahBrEC3Jg
cKlnbzA0rSu0DrgDle7xWtK/BJm5xNEJHuReRP1ZPEZ40Z7nb2Ty+bQ1KkpcMKKZ
`protect END_PROTECTED
