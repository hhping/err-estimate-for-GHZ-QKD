`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XCcCwZEretSqGKqojSVlz88wmWXyUxXNnczvL/0tm964QzpS/sEQF/ZEhFRqcv/C
2gJxNdR9rc/VRzyBcIoB4E0fyfxM21sSwSOPM27YSVKGSM00vquYRvuELz87WdwN
pDpXbFMB2cHM9isS1+sLYXzrh0Ik4u1fry6p8giRVXXzLgpifERPvTak9aCZoK2f
ACiYhm8ILxAZJWmaNH1AhO4d0D/eHftz7x7aWYRyshFfiXQZxazakWA5AcfhQS/H
ViK4RHYbkt8/XiRsuT9jqfWdiee+oEQi96k9sVoPaXkL+SYO9IwflKSss5PBtJcR
N9y2GSiwrBlGB86AOlppu3J5gqdrwa+ZrRJk/XPEEk4l6QEXfq/jIp9w6emlPKjK
0Jp/DcNvTFcNt0fo8wrO8EfYOCY+25JcP3imuAEdJ7CUsor3OoQTJqzoHvkkSo7U
TZzvgIfQj0IJyppFwVhUy9usQH+RlUCrp+eZn96WDe1DAGBfbc9ucBLfV8a7C7tM
JkGgQQ/xjUulJhjxf6GmZC42B9sRYnZHurTjRvBvxRsiHtLvkaGWWXLven/U8iK3
2WQSxYUhdENGnCsmU4BmY2I6y0nKeIYfR/Vm0ocSn1Nby7spRu+zaFTBNLzR4aEi
dLK6tFsomu1cpBbfwziXElwunbLymP5wF+O4zQ95NnU=
`protect END_PROTECTED
