`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MVYmz5Zi/cwHKnMJuaGKexCI+A4TCYiwKRDYqdX4xRvZ94Yy4J0B9mJgkz7YJ32y
pDTRqDR3pWgK6qsPKaDT96PApYhxC3FROMaivEdgAsGlO4hzAZIw+Vg8HDATozTY
JU/L1SenfeGvdSq/VL2vdvtfl7BCysMtahrrQi7MIyCuk94EZ1lwzFdLqh+w8hDn
iBPcNcqNsRt4yZKqhIPkZCs3ds2zyRJV6pyt3MFXWEtKZsHvc2W3B6wrSSlbgnis
1tfnWg5i7U2nHwUpKFuhEWFXg3L+TMtUfyWRkVj7iBMeGFyl0FBCrrxVD0M6nFmG
Gji30gf0f0fc0tzkx4H9A1H7ZsNRbayGJaQAgMyW42xAaZKU4U7GPnUVmFijL/Fd
a8QWz0pwtf62pq9Z0GIzInr6d/rQ9hs0lORlA7wnt/XuDAeuM5VR3EOcFOAumrdW
XRdxqcAeHbC0DZ8Q15YfVgOSAOscQyInRpc+7KaHD9sVcrD4dyGDsmHhpoKFJEh2
4NspPe9FNNR3LrQMaPb0+OCW6Ekw2jsW52l5SwOh2CsD1Ky1HoSD8cRBHEHWioJZ
vmgo3cEyImqJDUUQxHzBB36FXAWARWO1hXc+wZjhPDG3Cr+695hHzEWHeKi80Dpm
VXqac8Q1o3Bt4qy9ivbAezkjUMnjqaIm/8oo/scd+WA2AAAVUbvlE4fmC3bweKQc
EFRLMcOP4NPwjAfXGSv4kEidXmlq16sQIbY1kQ4XUDKgJ1MqMYM7PGM/BBXgr1sM
qUbi04DPO1m1zFKWgSH7tYqptIbow0b0wM3siwTQ+GDL+othtu/tPuIv88szYCGx
NXutyGxdll7i2LPx5Y/Tiyr4JZEoKSu6twN1N/I8tkAogCzHu5dDa5QY4/D+043d
9U+7agLvwjXhqcV3z8BJ0RFWYLRvpqd0eotvgzsrIz8ak/yXlqBzjyMiND608oQ5
R7GQRa3UH82uzW7S/BI1LhuiIrTMojYKqs91KH4Hw4NZoo5NlIGFnJ287ntn05Y2
wnfw9hHLUtr/ubJoMqxyUmWEBlRkm8NiDGV6P8Ddv6kVqM9YygANR0X9/aN0e4RW
4dSiT/iHHHjxI0putWPm7tJhgHssteGSnaFND0q6H4Y=
`protect END_PROTECTED
