`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fFTGVL75K8C0kwq+r2OVmeMXhBdETrRpstFe4CerTSmlY7ojWshs3/VnhYJaxQRV
l3mOS2sUr6TLZims4+MxzSYw5iUD8B84j9OLqedJ/P0gClwX4FFaR2XIMQyNlvno
o9fDQp+yHAzxd0pY5iR0J7OHBpEu5n/p8yid0tHtc3azBCat7Bprl4Z/RrB1HF1a
PcH/BJbq4kTGgBkbSduir1CzpEk4qkZtiWTqvq7J5oj4t0K9KJU7zALKpKwjTGF3
WBeTqgXPvgLamSR+ok+AMWsFHB4P82S34VKH8M6bmFJausgjUEU0pJm7PzXxX5h+
79AJ/soDu8eeHruU0Vz3Mufo9yZdJiYEnzW7qNg1+XXnwoQ7bXLwv/9jgl2vzcgj
ryL5kNG9YODsjiqxmoQdLTdH3SByiQhW9YPTe31wYLBRdVkmcnzdynXkP30VY5uZ
mRw4tVN+kzjIXy1IX34L3im4UDFpYlk+p07vZHXMryusB8VnHlpdQDec6Y686GKQ
NNXlxOwCjdcV8+/y94CKFvG8uppPzJ+WOxjn8kqpYh/VZNdp51rRbT+xBM9DenbB
nrwR8WkEA/PxiFUwgKwdiSxRQ88nhvRysJIp7uOrF8/pSFO/ZLGF6SjB2qSpYFav
FP3fpLS6wbmw0NdNyTPz/sVwslLLQMztVeLfgk35oVbPAtlPF8v+DGzCVawrHEJg
voyIEFaahXNiuUpkrIMOUEuYMwdMpWI+642ZnEGRb91koSxFarew4MIIXgx90F2Z
bTROLeNtXl/FcO6AcAMIBw==
`protect END_PROTECTED
