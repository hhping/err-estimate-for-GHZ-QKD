`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uj7toiyASFnqYUPvnURlM7embH1Bm+B3H5uURWkMI6pPnPMY1PtxoC5VjGQ3rFV/
PSrUnDGZhRTOxT8wQDk90BcdPvOcJF3/B4HxlrDxdOtoD4iuPeN5ujepCl5+FHO1
HhC8XXVP7e0eUN8/ikKRgHMsZkiEGZHwvCK3YUmreWmOLI7MIi9aIIyY9bVxB3tu
UcUQa43XyCKOkgFz6FOvMA0FgvV/hQJ4vsKiPmwe9OphgyeG326Jw1C9HV7wQLfW
6mAIXp8Nanwz2kvvl8wFVZE7FvUW+nhBotuKfcRSWYMC4ljsa5MTUg2RoKy9b1IG
bwOdj75p2El6JRW5P05RARAvNKikiHSl2r7riFF5/hd+qHspShj7J7MxekPjo1kT
ynG7noYZm98xTymnxxPmwax4xxbe3jdSkTpq3nQWf6VfUmpxepqaBP7HTl0VZxzw
3SwqFz6hT/N69HcOXSlJsVeVxUjhsUM9CX7V4bgRAzts8HDXfW4wk8huDksLAV1/
jRcpBS2oGVFISe2tKS0VuEhr4hrampLcLqEqfFmlgRBWg2Zhy7X+iJLqS4+gEjxa
iQI3p6IYaDBMxRa0pVNAgHmLzIP1S5AzCMGBCwiV4OD2K0tbse20kLcl7jBFVgw8
yDW2IvlDeoNCRBCmXgPn2p3ekJPW9QadAotIscyARaLTvyPVVmCgfxF5JxQujB7u
Ja4e9HlPmmR/PQnszSyMkSRft9+Rml5d2juNjCBDcV4UbHFalvSwYrxrBT0UKP94
rcdq4ZEzIguAhXYMji8I2PXYOSs+KiA8humFlemx0/yOlN758+Stlfl1+tnIe8bD
PTfBp8q/vUA42GBfEStgvj5M2Wt0Q8N9TRz3cF6Q5anihcBAwvv+SvJTnjcOgCQ1
CtuvV8fXW3YRkC/KTCnWE4KPgFNbpzLH/QptzpC6uONRjHGpedAqrcDrr4gXFTBt
+mMcBf5ko5HSUz+F66aJjQ==
`protect END_PROTECTED
