`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dzrebKI4PfwmfffVVdc1it2e4PvZPPVW/k5UTqlrRslKxYNoFlqLkvywnPNifNcU
au9wt27LLgU3Cezi7WZv86bpDCbwGxRfWdbDm6y1Pd8fUgYuJARnvmKS/1w2azy3
hmFIlvxFH8XPIgiL/fxBBrKBqPwUmGSDRMUrBOmkYVFxTQ7OsOsD4h/UdeFVTGF2
LM4K7zFTgKc2J8JPcqZOJRSnKYpTXsbvJK8bNR9Iot3rrufKoiccc/+gXq45nWq6
jG9ftGhcJKkmY7EfF2EA0lqsDjeE4ESflfLwZ/sisA5Js6xtOdd3JTY9NjuEEpMY
BmIK/WkCKLE2eiyLLKa2huJ+deSkgRiVzQc6ybIVMJr11oOwkuh7zIIzn7N/38IO
xZIYcIuKUBQ+0Xq+5Mgp7A9swXeI6xQ3tEi4cSD9oI5tqyvJyKphl4lZO6M7DlMk
Hr8822WxATbM/FGF2usLAWRy1b0SDkObUZDJbaggLf0wOz6Olc9rbr7e+WV/G2RH
f2ROc3ViMUlA6WFwYXNGRv1qi3KgsTmX3MUyP0ML2oKrYC3HPxo466Zzf51ivexn
XFydfQdqMe7QXPeR4bHZVqvgB2+Sf8XXXsmfRZjdRZHtKrbW9JZ3s12ABIufpVyV
d6/MOvclxtKgqzZDN2ZRTmycU3orId/nfM38zT9Xgn/DoLdI1olhj73x3BqmR6XD
6p8bzdWni7lKjOvy/WYrwMfYdekLIIQYKB1erqNEWGukmWB6JNqRX1P07HA2GLZA
K8Zj6jh1hcuyDi/xTKpx2RaQNwh2EoskiXAfWLg/nkFVSaLjgXijWaqCu7dSGyLU
/jr26jhWn7JTfcFrpyq20iZnkTbghalUECHLvus+ZMG5VgwUCVHW1sPzcNTJIHWW
wDBz6GMOL7MOsNa/9+lMkD21qNGdOweQm17qtajdzz18dn+2+PR+L7Eyd6Ewb9Hv
xUczjvTZHuVASupm0OL91v7eMlIyzLS9v03keqyhk3jsgiEVWtyWsFoWaGj+a8X3
Aqh1IriDUV2wDuoXCRW8rI5RCad2Q8YzAX/7Xqo75Vcygfpd9fklFaEQP5iT3+K4
90+9DPujhKbmr4QibCRYAM93GLJsQJ2mFL5k1Y9+qgnYiYlmJXCYf8rdGCB+ZsNF
gIF4pc0jK/Hk7eHG/grEoQ2MPJDlIXjXjnmhELrIjq3HB2GVhpyRDBvwQH4mR89+
sfDBnEw9SMIFS1KBaZ3HqaMeUQxgbb6HoByrNYr/tWJuNtr0DCPWExMuz3L1oxTE
K2Mmd/xewLjska9mJ0/ty0G8gMGD9F30syEz4pyk71o1/rbAPStH/+uTNGsE8s0T
RkYvF8CW4MMahYgJXEVXaJojW9te6JQKtcHBUv7pTfLTwGfFcsZBMsBW3e1xrsWy
VT4gL8PFnKqK4nUn4B4FYzCkUvoHs/434gYawVzQr1ZXuyq8Rj2eeJiALOmaSiBE
2ZImBPyFEzRnTudggK3TvBlBVm8k2+aVbsvJHuaueOKLGYKWITJPnN4vH4P6QulH
lUlYusa6js/nX2UOx/I+mCw2y34kytX3E+U4MTGt1CC5aw7eicud1NHr1WLh3Ws6
06jkdEe937S0ExJqmLOcRZhvquVLFIk2IcoV3PSjhdZYkSAbmQAAmjl02CcyN0mR
8A1tBMK2Ose+YfJCBiWyg3cCAl1sfwdktmEuGo/2XQYNoY0pg3H0oNRTFQ415Fg/
Vu9DMsIuw/Z7V1YhogOGU2A6wWxiBd03cL/rmi3t2LZHASOB6SUsBXL4r0+qR2qX
fLB1aknmTuMv+N1X5r3CUJUALySN98q6Vv5P0H95bh93bRoP+8Rtl9i4YPc1GrJc
PFuuCUclNXlfoG/CPUUrw2WeF1duaG65/o/I+0FQgH3s89aw7fFSf/u506wvO9J5
eIDJcHq7vACmwcMqPIixletyCLX8M48eSn6aA24+MNPWi94R1OPajJ3aAQIvVHh4
6wJeFrbBrYIRU+bgeM1i1ZDZwZ00ydy3TNmJgCYvsBhBSlIwMF6ZBDjfp//UKte3
CpklFjd+dfGgI0zTqBS2yNWGKmXLgJcgekZx8tseQztTjY5yu8Npnc3HXG/50oBs
BXwGjpK2LCc8wPfmv86PBaHk3Rl6S4GiCl8GMINcENqDAXJIHeRMXKuF0MiW+ZdR
/14bSeMn/seOmthDt7PJl1Vo/DrlToFUAzLBohO15Vskuipq+wpw/U6K7Xbtz281
4K6QVWVgL+xuz37Zdm5d1YQI8w1JJtzMam9bRVVzpHR7hsioF0hXmBL+pCw/lCgZ
DWpTF2JgJ7a3RUYzbr8RC8WA/VtLvn+5AAqDgG/Em2WyQL3KcVHuPTK+afq/6VKD
St4X+QnaNiqIOPRIVupMrbVhV/xukyfB6pB5iYuupbSbno3BYaMbQfGZxzkkRLii
9NfryGM8/jt2lAq7AWgTW0OrkAJPW2Rnxdn2hbMulDdBNSgJ34qUkgq1zZkWJtpf
Nax8PuUSXWytAB+ULI+HubYhpHGhD2sSUsvVo9wjF4dUUns6sRgz4TMcHrFAEVtE
946f4RdZVsFqiYjZdl7NzTb8TQzgIfKWm2NX5OMIZCws9i/T95OBWaREiy8EJ5QT
zhJ8v9cRjEhe6bNm1GddyxX+/UElVq6fFOzdq9QNM7AtJLjZ8xzK+n5SNvrwULzM
hdtlDbANsbooE6BV0xmIgUzAXpnhxR36uG0vzwu42ZyD6kVlxOmCbKKFJYc2GYMw
Hw+oRmyJ/D8XIVGCNSfiADHOZiKpKYVJ6280kHNZwbmodDRN6cfgXtu5hqKtPSbt
UxPA7DaIz1ofYjUIjClJqXiIfdKS6dr/lIBafv0URE03qcTZY9ROmwYL8gdWG3IM
FG0WJt1GCR48a3+kXngq/FzsF9qQqYUcbuRH/76dizKzhgD19rvnJ19buGi/rYdt
8UkIJb0Iri/AwXbGdSagaVbB3w/Yag4lYRtf9IHGaeruvGvJ0GHmaeiUNhICxz13
MeBpfXLfYsKsHIinAAYsDJl3hubM273C8Nb50Sm8pD2+dCKT8PJuLN1+4j+vL8t+
ptwkNjF5H4n0xLyNTX8D2MeMZ9K19cs8m6trT6IrqfhxFY4BmT1LVenBJICKFKg4
8wKfppW4iazq0GvTi5Bxhq2YB9Df8ybh9D0yUqug2Zqinn4qn2oPhu77Je2o62sz
mE58cgrlAF8k6mn6ReU8KlljqzP8vLVsKQzkXUoRxx0bAxN1yYg7DHeW/Lh3dDc+
jNC2lqgqNAjB+4sswdAbrVM7U7oYl2c+iqwbIIxT8uK4JukyX6ypm8MfqJ/pTajG
DkgWmgt+ZzrfPj4NO1qAswFTL2KPaSwSlZc31Ov4krtPFU67BBb9JM8L6Hv7E2Vi
potJLrZy4R6RkZAz5trv58pATLoclBNZli9DGK/mMTdQnR6ykKed1vVTn7dpYCNC
r7TSEmchnUcmurQB2vWED+5KARji4JoGV/f+/QltmIyeR8KqRJGHeWY5tAeFQu01
BwlbNV9ht35kuD2vOLw4pyv/+sJGTZ6tRZwfMzxLPd24pGIalF1LfyU0u97YOCzB
Nhg4BkrNe/2gEypTU56nZXnP7ynrr78Y35j+DQO7eJYmfaMgZdWU0eRrvJlXPtaq
mr/2zQ/nmfMAuUdZUqxE1IVKaFIAWHgAl0kSz+5m1U2/9Gdt1ZWFg4aK+RyThaDV
GCRoMHEl5OW1Uoy9B+xmXJuzvrBvwXJiyuywTdsKvI4ZSpqy4SSHLYld5DcuuJF6
mPi7UEr4jug2G21e6rg/luCGrrFuIK67ACChOHjNc5JGApCdgmeR+ux1qsrofqIN
a2D9FpUHe6O57y1vCX2kGvOBAw6QTRnEvLh9LhNRQe5u9I4ESiZKsiVRMY6Q8oGA
jhXlJLYWXCppc3ScixcmS0Zb1RYKPS9YmBRFjodfaBZOCBX7GxNZax95+cyuhlRj
RjwhPQCj4U8rjYD1Ih/w4xRvDyqF7Recmtx9q2nco2OfpBMSyNMZgs3jjhjsrzAV
hcwAC0VDriA5DD+m98JfSzU6JJoFVvt8AvRed/Qi0hwgZrCP6ktjuqNTidHQpST5
83MwTkv5uMhvD7bs7vQpjGyE7VsBnAF5pJN/OCT/35B08xfmm25U4zWsFcAWTzbm
9Ov63MBU/r0LUSxRRiz9wFPxPHbgyZbPMVTTT2hvJ3iiQ6RnFFA92I2TEyG4xSD9
1y4c6OOgq0vtNequctPEnRTtPlA2yUIKfmf+Y78OwtMmEzgJ0oUfxCoLBQy7S9w9
1jO/qKrwSf971WvMkrkfz16krDebbxKg5njhCriC5NkK72ZaDB7DoGyc89TgTA1r
zSUF5Z4xaeHGgdHSJY+fwQ3tO3/7jLWQQxMxlq1GuvaPlVFz4KE/C1NOMKJQcR9n
`protect END_PROTECTED
