`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6lhn1/eKljv4PtEg0DLA8JTtr3Pcii4LngRFPcPOhmWTgcqsBTO/IJ2DXukf6Jds
OYn915rqR8IaxMomaNolPHckir4CC8TWdFPbjdWlgnvJTVZHNQJJCOWZrCVVfB/5
4T1PikviRB4Clil8WSF+ejMBWk5naTi5JVbjWcVybs615d/yh0l5Oq+Ku8TZ9GFX
WqHdfw0KWAR+lOeRtYR4QRM6a0c555RttxKNBbCl8+b+HYDi9cUxGH5RNoKhbG1u
zOWA+RYKLKoSfx4swGhzmIkjOX92ixMoIu1ft+QXEHyUMT+ygrbPPlFtwIWgPhNG
eFOOeL6pTtyEzfdUPvbS04s28cjFJ9xET/lW/RSnrlVegCTtWixWcQFwBhqUiTqg
j8ur0Wnjhvl/6j5roEBaVrQsjfAbTjMU3amVSMs7e2Wwdv138GrpagW2H7rXoZhY
Paw5B+hmL0gJ69iLFbbyejA2CvCUZqlPGO9f60eas410n4Pt5b/19MBkK7VybNTq
XS4eMiI9h5/E1yHCgHlgb+zW25nsBpfbHb1D/mao/Foy3i3cR0/WKFT9Uipw5ZUL
bQJt8sByJVUNFARRraikbdhxOIbfpS7TDxK1g52cgFh+BmhgWwqTFDVAan5wGChb
R5eKuG6RyO1Df2lp/Azu/Cn/xrtTHH762YIPBDZRECptYJz6KNv+H4tusJGMHQKA
feOcknj3AAcPwPSOwmg4aW5WR/EvM168lpOQwkVr5RysJx3NY98dj1ElxhKefwDQ
MiigR3cGiLuqCMrQLYcicdBksi1GPZhmpscmd2qtGwV5TkxfHyB88/HES4W/Oach
BDlJ5peAE+P59GVy0FLuzv0zPfu5Xz62XwVWCHN/WCqPV4qARV9yjG4ehkb9RX7n
WOMByXaxEWKjjBIIOAFoZwYWqubK+9aHzzYiMIAKJGJwfYT5rpi2W5o6+/HUtXPU
r+L96A+cgxeZU1ijzxSvtJP+2fHaY4ztNxHBEYeIOm4fbFDRaLRtE2xTbP3xPtIu
U94G6Mq1q/pbl60JVwTYj2JJvduHCXbO3mKKOhPaxercBDUxtVlwYg5CwRLNjHXk
K3BRv9Y/Jeb1mIUCFNE2zSQg+jbqIILg0cVsUo3/7YARuo3E8HXbwb4HvypwIiLK
2jWBo7Jm/a8MAs6LcbQLVbMKMeiehSG7F0bk/6AmDmT+L8H+nA5MRrzaXaPfFPbB
iFG/oriuk2Dly8WuoCnrVj/gCNsbM3IvAeGNC/fHvm4jY9fF2EG7TyguWbYXC17+
h8E0P7TYqR9yqh7EDbc0e0TWu+DRVUDaIOwGra/cu91bt7jHBH7yRxH992wl7wy5
bADBc0YafY+67UzODPciEcVYYD8uVxNchZGQvBUIW5+IfzorMS/rL1V+aMW+2djV
rWfOXKowi8j7yEqFsaFfAwqqdT9UjrTSyZgSruMuhA3zmLc/AuiWBEDQIAzXQ00h
PR+R3W5zTTPteyZ0FXZHAceuZrml0gW04zmElY0Yndf+m654Rgo9aoCNrbmGGWrz
OsInY+d7vLOL72U/vGE987UYoYUfa6k3uHSw66XpWHHX+04a83s5OJAtSapFk4qt
TcaXBO739FB9r/jpKO4oLqSXPaySdhlw1drF+jxpQ22ssADZfLmrWj3f6ufGLBS/
AzMHwzww5DsRb5H5fLCUMFQcnAo8oU1gPl91MMsdiqMcb7PFlkfm0r2ydV9ZWl9H
0ky5qvJQVxhd4lGDuTT2apC6ev1NPO+AHypVDzUQ+B+gA8tAN+Z3hZD8JmwFxTJ0
IiIJXG8PounK/Qimjri4svhtrtiRzeUEm/qICv+XPrPRPV0NYAlZLn2pkTAC3ROw
FHsPR/yiTLvhrfSWNk+L1bBYIrtasVN4SqUSHGZLHNxHq8wiq/+zgh/NQldZnXYg
`protect END_PROTECTED
