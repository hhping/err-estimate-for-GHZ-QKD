`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DCkO4hOsevreZc7PiWq+hx0yUEO09RuZkXhtyb0C3Krn9F1DDpsp6gWCeGhi6krJ
zRp9AJBEbdH83k/JfPjBJ2Bq0fVA/RVGpbuXqr0bgjSX9+tFM9P4b6PgIg1HvxW9
VIRXUOlLrx0vj/vHCsSmuVyc+n4ZXAmNnlx+3Mz8WVW1fcGgrAYyYpOFkIfKMVpY
+o4R1LXuztTKjEO3AekkHbPZN7+zK90mCWbQuaoQ1TKtUMfbjei0JcvRAnKy6hjw
bkK6pNov8/scAinNGLQgFqKBii6qOdHIb4k99FQEG1zXs+Q+6kM9uHIWPrp6+sXu
iBlBURtaXiNvxDQm0qDSKAyWhBtcc9rJGqZM7XnH7gUq0XmMAAkzIz52vUE5jR2r
lSwwa8nRJN59uyQR2vkS78LKQFxXv05mf8b5bB0MJUekGDxabpUlB2Zgtcts5CCO
0ZNLphlzWVxE93R7xt0aSnxEjgIK3ERR12SbDY7VI69UlmTYu92zZt85uHnxZNTJ
F4KZfHK/PhlUC5YiMJgPh08SsYYD6FEj8fcF4vBiL/MdI36DI/wbKbv8D7xRHzWf
9aVrZEFSvL0E576QzY5K3Vceu3IUtHf/mxDAgHhYv4dlpkxNE+b7Lob7pDDTSvhM
GBV7PTBBTiknMQN9IGfNnQDAp5Ni2Py6pHCDLPIzntnXDy83SjSRaXVCQaovhmdO
nvsWAkXSVzLAQ307FABgmULa2YnuopPbOVlC75vH+kuRmuvoX8+RZpTTWN8g01oI
nLQ86NVae9ag85U/+DuBhme+slzGxSArKjypj8GOZGEw0uodSBhGI2aK/0JHEudd
VW8S3y5wtmB2RkoJAoEmbXaiSsRzF4Mw0W7m/F5g04h/5ALRh8CjI9FL3nutl6tF
W7iV+pQ2A9iRvQPes7BB7jDzVbEJs8D8NuyYWkpiEBL0zObiFvEG+Sqjub211LQZ
7zLl1DxZ1AyF8iMqEt26ZylxBA83F5YRoWVX+WtsSGeg+dNFQM1BNr1rZGUtcDIf
hVYsSfvShaGg+9AERTho6C+PSEaAQaTGFvtbrVHIVv6zs4K1jfpvVLmyJi2ToyWK
yZDrZZHWFdtRqRPDnujJm2+ksbvFTs6cH3ugpAM1XUkqPUcSs9JZ6zadt0xhl6nX
FOqGQNNwz2n18SyGbdTTconW9OR9UKOpj45O+zqfgKhVZ3iFwL/EIT8F0e5wx7Lz
3CDdBaLpCdA3+VK9GiiWrV4UEEwOfwSknGwngEEGQSv8NKmHAJ4FejAQDCjRgV5v
TtymANc+eNTZl9qpOiRCA/JL3+LCxGl5TywnUdM+cadiD/rnLxK+GpL6c5gMiTLd
z4pAmMT5YTGM6pRUQ5JQxygwCPLEfxrAi2Ey591jB2rd7IQ0DqVGAq8rWLbTvOe/
xqU9TZrdqteyQ/wJW2EHbSe1kmz8Joy6Sp+YkEreGTZZpz26T9LmtS2xp4fbWRMv
9A4oKdJV6J/Eks+isa08ytXWCx9tMZP7KtRNRGHELOu1VWzwoqlSsbKCuzuyevKX
2Nu5xJ1tTS4VU9YIbLzHHgrA8De+06rpF9cV8y27AIqr0UX4sN+xiDvDM2hViXSJ
Ae830uSVDdGQ7XcLbNMBhNf6//nAk22FPVwWdGnz452//xiPPBIjFu1M0MkxzIgQ
BWhZSaSMO8jKg8U7c14yNsaSfS+gXXs7ISUzZdJZ+JL4QYOt1V+bIZ7as5pRPUqp
oPV1vxgqrqLKI/Wa+zCusG29PyZNyypbfMGdvVgWVgumWAPqE+wr39weYQHaBvV5
giZOGe7mSIzYrq9PROsZc+YDNoC46RodQHoQrLDb2+Wd8A/3nJGAmiyCii2/k3+s
3rXnNxFg8qdIe7MS59UzuU7F8pmkp2rGujpCNBB9n3i527Vet+Be3+kh1ifsCWXD
ExsOWzg525yi7mdRH0XJ+tCo0duVTnjdH+pKAvbBObvynldbTMYjoCKB/UmgXe1G
MIHovPNcqlgXT7Cqjk0gYWqAC5ZT59Rf2OR6fPra3jEO7HuYb/80gvo9aXdH0w9m
9Aalq1PcrWMkihPDx/iFWn8bEm+jMZgYE4zqgAXUL2fnAoQG9izfM0q/TYZLH+c6
CF28oSsF5fGrt7XfPOKMrxf2khAT+u0C33k/UEQlrrWQVhjQ63MaAAsmsw29PcgT
dHQUqT+lxZYpuE9XBkQgW4BIpgjSGljCINZ/gxiXrlNqhCuzZtwZSopTzUMXm+Dh
8XHDdl+DSshCNugULOV3BAvu/dO1jd363ybqlPZzeJJ099CoQ6Oq2Bv/hqMeJXxj
E0TJOjInH2tzQ3LAy0BtwIF03vaMx5MjWdFbBW4mVMcAeXplTvoh/waq+lbDKSDO
ht2Th1XvtOc/jxTX+Ro1KFkgJQMSXY+G6NVBoV2dUyBLaN+HjXSlGa6Mv4rsUYMW
0K0zmb4XoSj+qBWkNPseiATO1PHiGVfhvXueUFwv3BXgMwW+tX8h9zBdDBGbeEqx
6bhPY4IZYFI0vjCX3Ljwm/mtPOe7nre6jvwy/WWrN9vcT+yOXapcuPtos3VFX+Dm
MyKevuE0jT+gdpxgt5i1RxX1J+DspsVs/aBc7adkJ1FOCW4n51SaKsB4WAWxZoVw
BhIXVm1QTDuNbZ691k99G6D3szevLE5EPmJ3oGtJWrDdSSacnpn3275T6ciDBv6r
kB9bZAvSzrchCWfuZfcdPzLLS6Hc5n7o57L64k3OSCBNHZ15TIV8fGIyB+STtmtd
dKvnAWNlHFevKrUJTdjbRwgmSke33kA4wvK0IZCMWiaecCPWf5aDDS9c85KeQCBP
k4tOJlPTfOWTO4o4ZLngzlzeETpJT8Tl/FxpqO/61+ye7CR2It0GC+jB5ezXyLPL
FMPspAR1Pu3xwzxDNE8HgysTZdSE64S7wu/kAYUWG8PtB6g9pNtxcqJVmo6fDx5v
Gx290D3gaOENY24kWEZU1K9TsvyoOYbREPz/jRzGPtgavE+eR60FSEdLCNDwJeul
e/QSnP38upNijn6j7NVO3desVl/4DLEIo+6wa5p/aGprhk6fjoiPS0XS2JIVJ87S
mgLL0MLNK4L2cJqFYfR66MaltRxZZYxieLGVfAUc9yfL/ztBiWcZt5/bphwhlNnu
S9lOnh9Q9f7u0Pxsp64WbPfycI2saytyJ2wc8ETjCfJ13LvM/eNwaUSipfiDsGAb
VKZpuUABKquHw7kMWN9bMF3upg98v/fdu4LVMOkVfzAKI9IDPwn1pRmrBuK4hYEw
BoeKcIj3imMo9U1Z4mv+fkcN/VQPaxKV5/v1QX75rcsC/riWSI9XBnnd0kF85izN
S+TghhDHL8dXWTrNoeDcs11TByzahzIsfUqntvkfEiZsIHo2EbCXW5nOFhUSS03t
OwCuDZwirNFp3aUA5i5RoT1uHzgI5qBrosJ825KQCl4ZGryZ04nuoTsUvZepi27c
d0120SHIhrEu8VYOVYMJDQ9xIha6zE6EoXT6IZyuwA1rPc7OhyJ4CVyQPAjkAGXr
oL/zVhtrq0UfJZa4avu0QPqWUcBLbjOrFteHL7TywfLVOAqupy4w3Rb9aRXVuWfR
Ad4NLAn2YhObYxAPOU187C/SXZkiiYLwU5+VwsnAB5uWF8oXmBUulRVm7Fnvyfr3
B1W6eNkmCMXu9+5ghuc2skGXRIkcnmCPuEQxDH+7+c39EYJYqWISCFXrmk+LeWEZ
TBbwWn+/vCH5YbZvrrPP7TO6HbBSyNzwvWNzecmhpqqrwXHRWAl4P9WG4BPSRBs0
yB9eoUitRxPuxkDh0YSDHVfEJwqTfxtQMWbSLT7uJ5qx3qsSa3KPFUjdwtNLveHa
9835JoGuKhvWbh3hK+r8Bx9b3KFYv0K14Wx5uMMqNZ3PmCtDXZSkG6jvFNVyuDu/
KrwtseuOnXcfMlC7JN422ZpmcEIPj6MGlRneo3JYThHxGYLxPPLMXwpCpJ+oZTQn
F1ApuJB3aDLp6a9uO1YrDojXw/7CgFrPF5K9EzpKNSOoBJBR2iEjW2IdmVgzuMsU
V+ldcIb/VW2MoZZu85IDBUmBpkmbCp7NDD1gw0wUW7VeJnW8fxOU5KgpzotQfRn9
Qi1b16IFeamnTaTrXLwd3PywIqgovG2hHFxuDGfu/rDHmHp1i/eFSoFasqDo7DWc
kTzlTucRLNX/xkgy8GkAFtAac3K5378IVOpTCMr4P5bpbwmnUk5UpBN5EUdI7ReJ
Q/NraZQBHb8tK8rkTU5WI9N9f77m6WriMQSv/jMRtRmOkL20XxuxqYT+bWw/fwPy
Zx3m0T//eQzuEBRunEJKUH0Ane3dVJNDADa1RurhmONye28Sbqlw9jQwnir0W3gw
45c0nRr2kdoTBOZdY1raz6Jhvqy6t/wazsrvo/oDW8KtFV076Jhs+b0DI4vNLxQi
0ng6kT5qYyXkYJv6UXwghSb7UBUsHqAxkxDI2rffCyF9kxSTiLrx2FnW9WqIfedO
8e4WzTuLyLziMGXqVMUNAydUNaVKma28EnTvqWOJSqZrT3rKLiR8sCJWnt4pVBZm
MdFT7GTLh4w82oDMGNzvS/vzBtXaDWFFtXqPJBR2Kr3wGmG2zOVXLZYOt6JeZyYL
IhyM/Ks2ekjKSCGJSKkq0hu3ZA13zYetkyz9Hj68ZdMq8l5M/jVo+MLI2/WP+Zzr
rc8Es6ZF6+F91G2egTE3idOcqV41E7GcmhiAZLuMBUtk4IWC/dLIcWv6CzOEc7yq
h71SIHgd0RIXyTzG+oGyzQR5chfNBRuvtDHUY4bRTEnEsvaz7Q2oyopDo+erBUz1
QfW8oqNAn0kuHNVeoYhnJlVlsJhyE125RCrtB51cToixD2dHZsLGD7c0JIOUTN+n
73n1gmvJrSBohDkY0OaVhkSwlIRDzSE5ReuDGE7wYSrntNHKKBuir++WQMa2qRni
R/qp7Uhok355uRtdKvHTWBZD/nqfbPqSFyyetRXWJ/C0pYGqPc0QtlvJL2J4tkOJ
7aNoQfns4jpITASxKEiCoMuF1FhKOCnnptXGNqCvjurQDqgsjTxtJjL5Z/11aNot
j8kmvzbGHBCXq0Gki1c2mcGVDb/jzg87tDVWrX7wgxfyOtHuHptwuSE7DytV3VU5
mIixzwX0Vrl7Gc5QZyjPbsDVeWbnEgaIZ9XYN+/QVD6hnkT2ipzOD+w7atkV01hj
azjIwkQgi7zCEhHjGtLOAksA0SJiE5hBZMYF1oriThknmuPXD1vYHmqVIeF3GY4a
9PP42CokXPkkGnPMW3ijHY2zMm8OBe2T4mN3aO1DteLpZko8EeEa4SSAfRExNvDO
5ItShEHRVXTIxWHt7B2TiO8z5Xgd5+0b9np6GSw7j54C76fMjPB881RsTHkHzoXH
TSl+3FTQ4zNRMzNC/VpKaDOBaTfw2a0HpNGEkmwcAmkB7eAy9RytWgY0EFO/hTJ6
q0GKiYgVFmYWQcJE9xK8277GFzurkIvxVIwrz3Si2rI=
`protect END_PROTECTED
