`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H9yU6ssZGxCoqKxsJLtecHPhw0vr/Z72sBafRxpqHi5NUD8HzgcQXfgKEjgRmH3+
Qxg4PDFRuQ0JdwSPg9CJ/iEw/5x3OP7DPQiyw/MDG84z2aIffKj+C2UTCpExTo3N
N6q2CC8MF2DT5CxvZQAkLexm0azqf1sx29jUazkgsoc0rXSWGiSFiuhqoVLOGyPN
+KxfPdABYOmC4agUTdmdEh8yP/jxfbG6lo1c8jPvG882apVyZawlXJULlB1if+tq
3xjWWVrcrDozr1+t4ynHGXGPLhw1l9RAFZVWa+z8u+zS9t07ULKrOPHiPZUtCXqM
mOY8QQe5L1SZi3MlmpjPedqoI7z8KHRRYUWANHH3Vrq1EZPHiyfKN66QtrQ4UGdr
dvnd1RJj/U5i0+wWZf4GLHEinIzS2txGjJuUzfk4GXJqBeugoMUEF7/vMtXlYc9J
KpxSfzwclyEHK5d1NKHVh292IBqYfEH6Y5cHFFBuvn9HGQHaYvPsohnGifbAs5o3
y3p8P/JfK0Kvlcq0vvwGdviE3PK8gzAK4ePRVKp0iQxpUa8EHBI8erU7bj/Gq4Mw
`protect END_PROTECTED
