`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R1zJ01r2oaA1e21r2rachUm9ByCRCjvufTiwge10E3BMjVjwZ/3OiiGLZelEIoqW
eGmmXY1k9s06edqvtf5f4FxqfkYw2pK78mSCdynSmayUm1zyylzNBN11ADcIC8CG
xscEG0L/ftCnboYlNv6c7Oy2RIONvpR/++wxo70UOO5SX4PRM6keXMZ1ReJkVeC1
COadQuoAxDIt2hVlHn+ngbqbb4yFxrb/jhNmpbxDyxHSRd9Lf8KQiNcdUFeYQgjs
/1Dvj4UOwE5UNMIzGLPZrA1AS/GgnszlSAkqsSphtjI2mChyljhd8Ch59j4yxWRN
ubdtcHtAszTcaxDa0W+BZ+EYwAW2izcy6zPjKQjTpjICUEdR87ZliTb8BkDFvlDf
NmDQcLMhN67J8atLhIb6RyV6MN7cctX/aHH8KTdjcPB7CboheZsRr/qZR/gVHxnE
P+r7dvkNJk6eRwgT9/XrGboBWJ93OXDohP4JJxPkmDwuslWVtmG3F/Kans1Go+dD
iqXuXBEx96LgtItD8w3/O8OxNOGIr2iDGrGCDdZmY8ZnTYSdlTZ4TxxzRyI2UKo6
kcd34jEEcLOpeLlTPUl1+uYHL6nJmRv67QZXkn1k2cj8OuEZsvrgt/AGhkgE85mO
b++fkwefTR5fJ1XIK8KOfkIrlCJNXl/CWtHb/e3Bps2zfuYnXP7NNDxnEytjTBGb
kCFcLhfLThOECr0IwifCe1fEk2uU9T1eMfmBUcNxy906Kq0B6YGeMsMETbJ38970
Shnie7ZgDBbIh3pRw9v2KQid7nr1CW69aqPm+Bj4leKppE8pWMk7vH5SYxqUA8Co
NgGWIiscsyzUpHixSPR96ME/X45X0TgN+Fvc8+O4e/krQnLFl0Tthjs3y4mGJ3PO
YT0Y865jOWigthsUD2y7xa6FI76PPaN9dhUKVDUR3rxehYiibZY6jpzxyGOH+u/z
/YIJXvV5PJHMX4emR6+NgL4OqGr+O1Eou0G14Xdvb7Uh6Zhb4jxGrIRmW6fMVXNe
pkbA7WvlpsJadFexM9gkd3zCeTaZZ2ZoeW/iX0he11R7ku/J97eX8DDPiVJLXkcv
OgShsDKqW9vLIThHek2070gy2U8xiOo82PU1dysrPMAcVASsW6S636KAVrIsbcIQ
`protect END_PROTECTED
