`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cOGHMWTz9TYUHq+WU74AGjcmEiPAsB6kOAGhNb+0BLyd0w7WamIIMknAflTWESy/
MZg/9ZjW+cODzSuaAikHuUpmAPJ+SbvzFnFftEvYsPzbur0qopR+AvObYOxIGS/5
PM+jAFX7RMsb7QzYZgbvkHY+ZNAM5lY6wrhdD6X67YzMrlwMqGqDJ99LPG5KY2zn
THZjSSlDqZNqSBrBSzWtFLXwazo8/MDTrfosqRDj8xX5leVCGBsOyVM8TOVc5Iwq
tVfVf3eGS7SenBJ4sYkef1rkE7ZIocOSkYHPSl8OYWgSwpFdG29E8I0UH5A/bXyi
PB8S4E74DYHBtgmU2tP9i6hCybW+co7izsNBYHS5IM/wRTHlIH26BLZ4pult9r13
F9iiTg8kOYWoqRawdIJQkte4hqWCZn/evt6KecldYCrspks3x4c/TFRPtUzhVDBR
HleFl2p/YCBZ4YAdy+LVCgNMhi/zunpn/XNJlTOhGaO3qopfXT2JertmP9FsaDpF
Ta8Dgd/0lCtlym31OYJpso00fFO+cKcIoy0aGzGEjBvXQts6/mH6ej0XNsLPW2IW
KFinVuR5bhE3/OSW+w8NAEIvURBS0ctmNt/YRPXd8AAe3WNupJ7M8CfUjTQTFRmy
YzBD26LyNQdOnUElI1IAoLsSr1FWG0SXPOKCdzDTARws/tHR8KMQr7SjTb9aTvsX
dCK3gqYJz3njxvCRFg248ZJfACIUZFYYFr0EkH8s/RitsrAK7Q60Yi6hvcyAIp+J
XPO417+O5ubFFuQulkxnsG6Qlvpy4wos65pH3/p2h2Db+VvUfkTZdeLPATyss1V4
AHGrvA77//G9vBN8wPvcBsGyyYtQ2xuEP7EtMtihaJFPAYGTkwAsA4dJGUC3sTl5
+adrnV8FlQ6g1bVTb0RRNzOljmSScxZnLgjiIAzsZfp6mu6IZxPvXwFdRYET9Wma
Lj287R2G6sSjO494QZtW7rc+cAHURMeYSChoO9f43c8YCAMwSbxv6puIVOKfPa/G
xxccktT1YYB3Ird0DxCwVv/N/rxrz7x4d5Q/AzcRXzt9RueGLojV972IfmYyNamg
LMLEAoqdC1Nj8jur10QGTtwju6YYcNFaelofwA3zwgzCeBEQYkPBZxN3BAUWFCcg
A0/KfQQu7e1+qUglyJN8tJe06psloAtXV0oLdOV8+w11vqLjcQW5dib9ipnUP2Cz
5qGIQxRBxN9GLdLtRpco13pa/ftWGyouxQgfcRxBQZqcY0YObZejwfTnfdoVxmZg
lyqdsb/nNJaRS4FuGUeanTmDSCKLNpXB+eqQB+uSaBVVJujDkJnYaEIeGl8VvV6E
oEz+np2IPGdVIFdjpHqrLJB2oJs5V/AguKjdVXXu8h7J5gA9/Klv6VuaRnwAXg6m
71fi5BMVmL7tnF+/QfoWAMb/6pATB/mL0BoHnQpn1380llRT7ujdiGTZwFc+v3vv
T8NxBxLUM7V/sFYU9qVzFaZHiSU1L/hsemrxSxllL//jwjWteLvei0c7UGSmLzb/
yy0OszPcnYUfYHq98js8rFm+8Vbik9hb7dAcWo2M9WXXBCAlg1SRKNyGLxpJazCK
2k6l7Zh89Duaoq6OoFi5Ijie5uUnt/ERH19lN9IeZ9eM26xkTdsonnzXuKKxTzsY
H+mKAev+3RIE0pPTOLXmagmeuOT/avGL8eUpzFW5wA7DEqnmTM/UpTlTRZe0zOIG
0Uc9OjZR6hXL8jv4dgHA5k3XQKVGmKjtVgl/TRq9/ypzoJgf2/iiyX9j1vgshVe2
gPnDD/cz+eFRlTGNxYF6fqkLRRmin142XVqKJQc+TrRsEXlYQAoK1Mzx1XcM7xJb
NDcxHTFL6Ix2Rjq4qY3ngD7/pGSXSHgT3WfFCgYl+e9iVJYr2w8HvJo5RtQ3bKZ2
ZmzaKPAmm7rTVwA8BQ5PC6RNbP23gk/2oQyGRoSKaRRt+SdE2FrQq4LLAK4C78Iz
JNdbr1hKGdTaINa8FLWX4V5aIQXGmiYUqPwg43StSEI4E2x6QAnUurD1b42+EYQp
xihi+AF4U9FViS0sC395Jjwf6A6gj6Q8nUkz0l2MUgSTsYJmXjqtSQZDStU4T9O7
6z6wPQmv7sAbhtKPV0fQTHDoQZMJXInNHeUC044KRF8gpbZchz4+6u16gEbXzor4
KV0dA6iAwPO2hAWV623gq6z1rbcWfLv2SBBBnfiPviLLWfhFYjK5o+grfGhAtUQv
itvk5LborIFkajBcGaXp/ZFpcR7zvJjClSwFVNabwkXfaotmH3J46RPnpwRkspHf
4dYojCKEGgyZ6E3zmzJXHmTzTh9TcoJ9AIWIW49uLwQZpnlliys/B9IG+Zgqe/Wk
E3VEQ08rzgjN+GXmyy3/RlKPFG4Imvp6+7X3ZO0L6mBB9LSBqo6oGfIOUQjvO/cU
G0wYaxi4kd8q41663ehFRP/AcBLACQ9wwCpu8EBUIhpoJdjk9sK8IZHMREVtJsUj
GqOkAMzegS7i5FfFBW1CjWItvmeUsm1O1nyQA/4x6nr1x1fE+wjNU9PSXu2blHOe
bIJyg4QZly2fqdQSEULLWZI/D1N3LKogvvnW6M2UdfVhCDhoDags+rCbqaO8e7A2
1t2IBZgKaQjvI/3oDUqw0r4p5F/7XyYcR888vLs92odYjhfPjJZ2uMvqyZMYy2+G
Rl3I0JZoPVwwDapVZTCfgQ0u7xueUV8uCd2MIvb3N0/3VmLoACOHOqrIBMC6Wqvd
qWocDcNoh2JWBbPlsu1U7sggosqIyZNdZJGTX1n60s1iNoejayrzEjSnnqUlW/A7
WAqPn4OJWoxePRwFn+1SQWKUnAKbSWShyjErV6R29FXqZS4hHSlX9+8il400vFB6
BUlD2ZCYeo4U58+v38YzSeAWtI2z1oyCoTUSSiLotxH/c3LRuLIXnyGNznY0diF6
5Nlw10RoJJIPArrKYD6AqGklxRcNmn6dMleaRPiT93A2m8P5HA1esrxKOPtQMgUR
MxPnz/MaT3GEWQpS80EaGQ==
`protect END_PROTECTED
