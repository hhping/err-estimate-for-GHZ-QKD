`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+3/raPpsO5pnhPopJDeRvFOc82O10x2gYU94VrdPzzFuBScvGZ+7YaKe3QuAKqh4
f4QoXs6UnK4erUabEIjJrAXEiEiVy3B8vF2emTXP2uMZWFv5bqhzsr3e/p36z1Xa
dKmOaeyHHFLWyaXMD6uYV14TKbBz/Qn4EVnP7VNha5mRZmkmvJAqyyH5Vi3vd4ZV
BCOePyJcjIKJywXKDp7qtnXTYYuiF3hR5jayvHUYi4z1yzbjCEfTxuw2jwB7qoT8
cWI2ET2F+HNJlK1DDdsTJzzqOYbDpfs35Zo2s7rVqkurfbB4PqG447/pPS9tJPCp
oerrRi1OH6qMDZp4Ae7bDcAmVvslHbLErwc/5OUJzkqrZvkZjxN9OUf1qqEHw5zQ
izvNhPRuqHGLvWPR9WV1ffs8Ld/gX3lbVwpKF7SGAFKnEYEhvAKS2Oqhr8rFs1wX
IVCF1A1nZE936uyRBtZdeAf1SnTDTtitxcw7nwM2Eh8kL2zSSW7vbMhOVlttnnUw
8FeVv7l/2pZuF98cYKV1UMqgZMADtzSu3R3eEDxIimqxt3K35vKlWfdlxK11aPOP
OH6gtA5itRgX0w4l2n/GiIC36mo6n0OU1KlTnO0MvcQdrExkZ223n0BUXBzITz2h
SxBkqosbIvTlsKJyphoOZUfsZdGc4AtBx/4gEM5AmidCBKmb/dXfAnnNTlLbMC1B
ipixAl9EaSsRgGGbpZngfBjKUwZdKUDjGSR+WyAm9wvkXr2hbgQJeINh7jcBeeca
wWrhXvP8hI1Qht96tP7D9Q==
`protect END_PROTECTED
