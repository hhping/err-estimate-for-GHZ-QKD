`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TXksvyaMDJ7Iq8BvFSCyBvU3DQhv0VYIAjO6AEVgejwLVvm4ruUvpi7kEW8hTeyi
LGBl5baerLnV8X3jGJth9GqVMUrCC9L1CAWvv/RqjoC+FQ4xJjc/jwZfUFDg6+qH
9TwH/qxGm/ydURNmvPVyHDiZ2HqEncDPMnh6BsrM5HI9uJnVcMYp0w9RMnleYZyC
h5nByit5hJfF6kw5apdIcNsa7ZvjIWlOxvaOOMLPAotx3zsfX1DTUdRJBi414uHg
MfznDHasTtDJkm/e+B7iadA81MPmgG2q5seQPshY5VHAPt/2EBz80CDYTm18y8iY
co1rX+DbzNxqwfRL2rDiWsCIcKbXJapbYHXCc7i9BXSe0u2VMi1t6f8EGWbwzMIO
FNHyCQ8KBq1rbs7EM0X1bMq4X4hgfR0fVj7dWqJexjprC1RLgSiJmsbW9bQfWOBu
ZpgCNYaAZQ9T93YdHpXMavXCOHbIiKPePSCBEkFba27dzAeTb2Uwsjti9+/WPz1p
x1XdFy5/fikoUArh6bYf7+a9ubw5H7S9aR3RZoLvWXIsy8P88Uy3nFMMOy5PAjwa
aOlfTn300APGk4svIzNLEYtUpxVdYqqr4t05YOYNXQEGX/y33I+4NPTToAEh5faz
einra9flUxUuXLD6hCj0ycEr7jWjCBXXUQZWt226yFRXjcGM3Esb7dLVW0PTROFU
jMuh8yi/Qu38TVvCluDvnAPmj0hfIJoWzV6qlKH3ziVEDiT0lVM00yE9q9tT6Aeg
+u62r8Hfc5/+OkZWSS3LmvB4uf1w8JsXjjmthfqMlyurX+hGO9FgzSnSuYM+2SBc
hP2C99X1KNya9CGGsiQKcE2ZKZ5SgaVb0s9ZywJpu0ctWwOFOj/X+bIEWsk9eFfB
u5/h87jof9jf63JUQpm41OYNVajCef3n2NrU8ftEPvVI8N6bkxhHB6GXBPyM4aYP
H5ngsE+udbwEZY44kRM77V09Ke3ObQDjVCpLRrHhcS4jfB1sWwkrtu92A2S0Y8v3
P3q2QaMdSYqMZ7F+mSvCcbXEom9ITE6v6hQmHN1tKvd5yd6u4M4BXuI6vYqQhswy
N9CdzeiXvKUA1WaqSw/DbMmJ0Fx3aTkTFADytpK9jtT/li8BN3jWLlWOC8vbpsRj
qj7JexEYSnm1kFF3SkPjsiz7tp6FEkZUM1h2zVIAN9151g5CjPuglyx0v/cF9lDj
BwFPra/yPy2S2Ar/7dCr/3RxW2nMXXMaN4UL8TkEeolLJbys+cH0/fSLHxZPi0Mo
rzTXbuyo9wa1znSos580IZrKBZwf0JoupYQQwteJVwTEcG9KGwTdZcJxSzEB83hk
5dDUWualAKHirrX41CEh1oXuGGazXfq9D2EFy3zYLHzTm4wakwwoj9uvbqkufRJq
K1bWGBm7qMXmQm+GuHH3ZeX/LUV5c3ZA3IZPp76a6Y5wm1qNPaWCBKQpA1NCI2qP
mLJctOXEMd8TIketyfIer4A2CCKyv2ykvOUNH+o1aByBQHMurSWL+2AvDj5o6L9V
/DJi4t+q5Rm4JNAts0fHYwdAMr3hn0rFQ/ycWT1RVFJCLUUieWhefIGeeDQnMEMX
0/j11kjo2RN/hYv4mo1D27EjuJkw/GSLYzRqvuCi6O1+DdC0pRQGfCS5h+M929KA
Ks09aptDMRx+jkJSnASRzyTmb96Yle45AhFeujHc2gDRqOWj/GADZgEOeEFb7djW
4uxHlXMFcNyalw+XOpMZuQk3+VPCwIoMTE+bNPqcR3MzC/l4Kg+ZkQmXAFCKgEvw
51JGcS+hBh3jA+bYzeHzdpTSh1qbFvqn1xE8Qt8NCvbtpRAtLdffi99Ne3vrCRAv
OZmcb2ItGMcWrmll5fhxSjzSe3xEWfuz376lsdKY+j+lwzeHkHGW4hneJw+cUIwa
wzhwS6dd5ppCq1K9fuCFYaz3tvOxv3q/hhFHbTG8u3KUbgwmBhkjGjhcLyJ8pDS1
lVQA9PHgO9lfORdThj+6pWzUCXqT9DPQm5T+tRA25JY+7XPoMbh7iUDLw7qzPEbT
Xgx5829r2PjwAVxH3e9favSH2NM/lZpK/8xB+nKp+n4z5+AXMOyhDUBXOP7tshr6
Q7ZxNoYHUIbvj0H/33M/0kJOtPAwKxZTgaxJ6bKrjZyPM/r9sRGX1hfoCFeaBFAu
gc1GzmF/N1FCxiROeiTyJjxvYvQ6q7RXccy5DlmSFgCMFTjcRvFto8MWClAaggnZ
dzQNqfkrR9+dyxKazckSTKl5Ozz15ZWOKMQEFhEZgp7HyHHju3FYluqIIBncOy8d
uOsWA9PLhNlOrBrMAmkPBSy0KQIsgyAGbWqoqHykk5k3Emd5kJEQKcyVJykJcSqy
oTkuH8CxeJbymUVU2kxzjgxEkscPQDJlPPxtAg2ARZhIoNkR2FzfumaufgL4ciFK
Y6UjBRvMUTXMCAOTNumWa0uVRCyNa5RDosiWoZnG9H6I9a8pCAI4+xrJGHW4RKWw
xUty6YIVIswiIqkxllHnD5lC5F2YJgojC1WvoY/G1g7wVOlsvJh3jbYTEUYuuul6
i4fJMPquGUIsujtU/VdomA==
`protect END_PROTECTED
