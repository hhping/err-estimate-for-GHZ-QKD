`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6SZe9DjfNBINf4USCl8LlW5wngWpx9+EDiyAAUfeBKQ37U3MgswDkpFa7qdohW+M
wxkAONevVf16UrerxQP0LvPxGiAoEImQnkmf+AawyEOWpVax9KY26O4f+fZHp/eb
a5m8xhV2OuVt6NseL01JGEuXYneQBn7xzJ8FkXta3DruEcGQ0UtfXB3oX5pYuhqU
1blbZPD2CBHkE/vwqHuYW8y50oonFMwEYniS1YDbRPMiJpELe6jYf+FFjDWbNY9W
blKmTVHBIoma+mLtd2GCR9O6JuUCHx4jwaXlRPdAEq2OTr+Kwy+CLWa8Q4QcrRH8
R4/5UwhvuEknOk0Wf2PB5PHwcu8b2ER7M7/SvpE5OIAbs+rDH+F5hrHrxfbZf/TD
6IAm3aajnhOb/hEYivqtd4hgEOxJ5CNgnCIh1vpv9eijF80szFR7WWaRkV3Q9KzN
/qJ1VVDpbJMmryKffSk+1b64UIyltr2EHlqgNliv+NogMoP+RAreLzjVFIQ8pyfR
Y0z3F7/ywAV/LcHqd0MLMnL9JwmzMmJnVa1IwrhpKhtfYdaJ4AQplNNKMBG+3WVG
G8G8iNbUREg4otquKa6WMFvlO9Q7QT+lptKmJdUFs8q+UgX724RUt5OOXq79WVBx
1GvMnPKQvM9yR6BPw2J6fyeYBRa+c+NLulA1Lm0ELXvXIVV+A/ZscdBtVEYmeNl/
DP5iyHvSiIVoDj7TsBitZIdjgYUGaCQmWdexVonGNmMBbyhUx25CZV7vp0KKKzQr
I+HSoIY9FMXuLhCLleW9fe8ayueUkCLbpLrcjC77SIN8e0hD3IwYkg9Am2I/kkzL
ftoxozonq7SPLwCQ/f7WRAyCQtBtg88x10/7h8D+CjE2gaesfDWz6I0BczUKUY/I
XO7kEaDc2ClH/3bIf+L8xnmdBqm5jtLUyiJuU+kuv+U=
`protect END_PROTECTED
