`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r+EzZmJiAP0Y1+xV1hrdxfr/pD7XsVDSumjYQGMDl/eXoEQwtNOfrrvgasUI47l5
aY11TBFrHobgEZGpCDVDKnhcKBOogAb8rdhptuSkn14e4mPJfvwTvSR2ibsp79xP
Y0UVgcFWIVNWDZkGN2gsKGm+LAOz+GXXhq90FwY94TKYSLBPiO2m/DyfzVfFlGXJ
h/2bOdcm0HBVnFuKDSnyQdBHA2vrHVlU7thAexDT/JAObw8wkffqRz3Pz4ng0CvT
uKW1eespGQOYJ3Kg1Eem2joxfzwr3uA/T8ZjjmWn44b0NCU6FgudfiUqed5wk4wd
XRzmfkUZoeNNEBCoFQkHVoPMigaJkDGFG52wklqp+26UIxC0ZBR8CziBlz414pgn
auXNlk/FLGfHdpy5/TY4r4wnBhLuBbqNl8yJorkbPSdpOalwDwo29mMo5FowugtB
hRTql2G90mzcYeBUN8WsdVlFkD6MrWuuTQwmqfoNUAXjJh8pDJtxekR+qCndFrVa
Q5kHeJ1r4uqRvSpyF+kMjfZhBJuQdt4D3gyV01Vb+XUvPiDvbgJ/Z4I1zsm0sirQ
LSGlZNUP9RogJIrk+EO9GBk2Ws7XjTrT6fYBibvUZMKP1IgEPDHTETPNYLzJtyjf
pQ/UmFnxm7abUqIA4xp+sj8TDBFYyXl0ITJ2AjGXxH22dbZ9X80NxNA9zBXpebTE
BRGKDBIXt8B6HlkPF511b80AUOCtWB/RgoYEh7KkFSn/+WsSfo9p79vNJkyNT1hc
zLVZ074C8U1nyvGuBgT3FEQx8pNgxojP2Ak/JVuY2MiFrUWFBbDMQGr66471XJT/
g7knxDy2StmqauoRlpE/I2ssGd2nz4RsFyXWSZLff5O4J+ea9FrJr3Y3/KkIdb2J
wC481Xi+LuSW3pD8yeQL2E2epHuThy5Sucf1og+23S7bppraxns3zfEaf8foiqcZ
S9VtesgOjhCn7nXz1ocUGz2wr8DEZir5vzg4riKNnvTi2oPx7RusZeKZMVe1RkbZ
enHT8olqkBaCasZEvG5wuORE93QU0WTedUGeD9NE6ajxug/aU81aJLZUW4ahtR/F
iP7iOt14b3FKQkL9dfb4VoQG8LEmgR6eatkSb1DLsvCSv2Vn6ckBtodR77je8Sy8
jzK0gZmiXUQpyvECj4cPOP38DUhV2SYpSEGQyjKrJXI7bzJztqvCfZ74BNxqWo0O
5ZLp+ksupUzC2vSBWPwDmXze3aerVMC/1ibnUFGgUyI8dJ07hDzWtnJIU2v8en66
0VZA4JwtgyHEU/h8syd1+FJSZ93PqI1OBxTOn7Gdek9efYEhwHApumwSKvKJhL08
3/sa58xcm0URfWsA9AyLNkPpN83OJO2domcFEMEKc3zEQUu39TtkWRBINx1MVoyQ
id4JUVdokW2LqouiGXBwq0Hl2aKIX0ePPyELqq2A4JQgJljH75sDyFmrnTTYBBr9
VeeTfR2+OKffcd9eZY845g1qNDMF9iztZPzcO0tNEXhk3tZpiCjd0gh5f0orAUsD
HJV8y2wedZiRwfIAS5MWrokTjOyfmWrb9SYxl2Q+l1tZV3LJZxG9+PL/r/gh1a4g
`protect END_PROTECTED
