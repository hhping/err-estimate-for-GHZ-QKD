`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dXARXqig1q590VjawouGecaDW4WA2WHDigNsAiQc4oWJZinZsBACbNNBdwDSDNxp
9hdhVYCAjrPBVrckTAs/br46N04D1mRg4hUj1Bx30A5ML8owUQYuOAml0ooTFhNG
CUSW9sgyYE5ZYDcTunZAAsBvDekGMN2/srCcOCu8jOVgnQ1ah+j16c+ZWkT63xCJ
m+fdk7MZTIqP5GvsotrUoI6KFgNhnUN2vhJkt4yy1nvJOf7m5b0Z1KDmbNHypVlc
XyTogD0QIwp4H2oNxATsrQaI9VC4qFjEmdt6Pea4xchbwmPLojwDfSuv5qP5bzAm
SimJCQuAhSqDKXiSlGfQWq90TFOfo0AO8NhV7byo9Y151Z3d9HURtZSAGBLi7coq
XWA6sZr6rL1K6+/jmfRHzuEdfJEF7MC4GJDKtlObxhZGiBRLoxE5exOPskdBHrH9
sqjbs+PQfw9B5EoNa4JSv+BZZY/2+sWZneo6MxmjmjGidYvDRy9hB971QelNKLoX
5FeAnyT0m4ppBlEqDU8BOnFnLo+3RwTlO5iQravYnWWqQsnGGIDU1ub4PFluIoHu
ALdeojmzDhxgc68Vs4NXn8EWiK8SZwZ1GwX6ajTq8XNg5IfK1N5vd3r9RzTJJI38
CukD8LH1exb8NbPu1rz0JdU7QIktJAx5h167tlcOjGuG1H2VqQHjc5sYETMROz6h
mMpj4rrLRdL2Xyg+pOVPTYtMpd+xRwsIwRuPPEC2dEaSw8zNzgnsHKhZBsCT2wS3
5pqma3Rb9MwvyO61eMFY6YGo+p4ba4CMm4pk55m+mA2DsHFuFCFXdO+SavG6wF3N
s84BE8lUQ1hIOYEUN1FqYdhyrFKjt6XltA9AyQ1zqrw5j7HWzCmuh+dAwRGf7GWh
F2/pluJ1i10dqScF3tT0pmDNpe9wDAMwkq43TKzCKuXrT2mUrSHrRq/hSHPXgfR4
oKqQQodz5MPVkGBxXsrEllVVANWdew4tklRwZQeYvj9+xhPylie3k7FHfmaxyB+C
O7QzFb8cCOaNmAm1lLJUHGR01p8QvUX5Wx9qvLDDL6I36Ogie8lud5+66ZBOQATZ
a3NaSdXnIYgqs4zfcda4OhVx2VPDbesIt2XkVdMepnRe8y/r5LjuNQ/pEvIeNv62
YLW9CdC+ZadvEpDjFy7z6ts6CBfb08sh3Wi5mVmJ+AEOTKppuIf0A9/Vj6j5j2vi
nE6Dhk36Ayl9wk+hZtji1Oum4n9HSA9ictGz/Na3pai36YExv+JjkSSqu8yULFZX
66WlIvQAamD8RvfQ3NduhZ1uROdBYrOUbFrMIFilMpqLGUTZm3IBm/TC99/z8CKx
GIFNrEoT/LNxW6AzPtlRL/+N7e42Grsk2OyBvyS2jaNZzu3QmGxPCJLcItDK+O+o
u/pwqYaKjhozNEJBCf+FYFkrYM3cAIek2H2O2AbhZRQKyhRKnqrBpvjnfLzec4XU
Mlkux6LtC9reKyXGi3n2FYkB7wFR9Bci3XSzkadJFoOdOuFoSuR0P5pabEzykxKH
gu7yD9uUH1DvLD3QPon1hKNVI1JkSa9/hiIymO3+M6Se7g2LMY1YoV/ktChNv8lK
Kkt99dy3mcnKYpf/UeeRkNWl+E0GvfoxQwSh1Dy2/yRlPJEbKiLnJk6jhja/OitC
R76aWz7/prdtcZ8zxUVsD/oprfJnp1YFAOznFnM7TkCCI4g2ADW3hM9pjiL0vj4C
v4GPYbUF53FPYaHpFL+vvZ7cHFjiD/Hs4siS7WC1p/Re6A8juXr71opbh3nL7fxK
XPZPwhjqCm9luuNm+k6HzAefJPMJx6jsotWB+H5d7C5mPvg38pSIDywepsfSRJU1
lyD+/B9c4pkUF7J1t12RyLOojDCJ2oQxtVrwmY8yyLF2zQ1Ru15whZXC3C46P9z3
gnfdABwrX91haCkBMlBorjnoFoMeqNA2kyI90cYMqQ9nASIpy/oQZiu5D46pyDU5
ZTnhK8YgsGZpGCFJXHVqjwHjXBzGcrN0SzpXVXSRZg8soiziqptYt1u+T0qeIiGa
r2/5PLsB1McwYi/uYmq2hdxpzQ7iQzJtx9w4QUMzabNz3O+/kwxtwgb/TCnuecd8
E72U1IvWqMWs+cZSGH5TXnYAVdpZAOaVFhFGCJJuwtEQ4wiWZY1Ipyxm4ZM1DWkm
s1MUtn/+p0RU84HbqX18jQkZte7wJ0+mA5EXvQqpubH0gVE1J2NKU3mWXRGvFXFt
VWk6OUS4x9oL0whdcb3peebhqxRgE3pNjYeGm/4hH2z4miBK/eUKGsKCcKUvKhMv
Z16bnH48xAOXyThYXBC13DTAJ6eaF5rl0GVHMkbcE+ds4oZIGSgRLKM/KSuhfblL
tgfhNX8ESirCQcWfhZ3eFO88ow9+gdHpidmULlF/lHtTZVpkSSA0zEMZL7VOa1K0
C0rDbvcj7NLU7ZN2oiyn2u0MT0wkz73xYlAEmVarlSTvOu+0pzoBxcergiJxJylU
iscdetTyj69o/23dhc2T7eNnsNhsKeygBEyDVeD4FWR+jhHTi9DxFEDJUgQGgawR
ThM9qoSyN82f8lAhfIMwC18CwOGZ9sylNfelpRX6ccTWqrZc1bxRv0b+x8cev7xM
Dg19pidtl8MBtXPjSMQE98IUggfALbaTQEmWcbEUGbIfrM3P0RF9z/azpTMqjebE
zjb5DiQ3Fy4GqUzGr5RHpE4KzHYF2tVBIBpMBCbjjaDTdsVicJcjNkpSiCnNHYyO
BsqH+qf8h2V5FbToEqhC6Y7jnbuTK6TrXBSZRGN82pUwFpq1ur0WnKAVLDa89UlS
DOfV7VVX+Yr/Hbp8EUiKneYNKfw9PuZaVYfc6nU9hEs2TJZMLi/V0AURso1B8o55
eMuGMMWyubRidInC2uwOkDIQE31uq9TS58uBzU8yTnzlgF3m4p9yJJYMf/J8eW9W
TOScQYGBsjNxULxXcUItFddrFM9iyadXuxxjUsZZAVrpby8Un8jwPWr0l1ueJMSn
HufPW6u3xa26ppQpTbnaskLBu+JhzFr4rB+djKAcl9jzdrooR2pLQeJpyv1c0Zbx
v9j8d0D+7AmKCOLj4FzcmXyZ/9gRc4p1b3YFt2Ne2EtsQZ/NjwX4N+T/mfbzUhbU
iy/OcVm7BMovrUPWtfKNdsdSW7zh5GvJnPAWpL+GNTwR18Oy4lB0cxyvKxBhJmp3
bqavSHknGgTToCpVg7IjYEaVsCwWn2CFjN7rwta+/WMcNs/T22SCQlBSz/+fFevb
/hQWyEO9bUr9iKuE/Vwuz4/MeKQpJpM14aQC5F+ibN3E9+3nVH7fUFCT3NAWylSR
6u3MQ3zgGHf973BbVeoi1QBHH8MBWYTAHqusXKHiR5IqO2Ukge9EA4U4aPr/foIP
avFWLyFWRWX9gZrzb1DqLkH9F8SeiQqp7hxXTHHkPNlHEwCRndC3XsYZGKGrcVj/
grsuo6TZUPZ2eaRHMG9RRY2YY7YrGfvJJOT+l5iD4piP9jyZQj2UfVObwf33mT3+
IbuZFRzaAgDDxCkdBTJQAdAL3mLy7nnZuyvcTFQ2JSR40Q4bp2nUy3hCghqOVaW9
VQZGrY/zeYwa82xfXtwaCQ==
`protect END_PROTECTED
