`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0bOZ7Wz6mHmjeeIiko/g2LDyy4VKA650ielvDwJwheJ2aplatGm0/ogTVVgiJ3gh
7Im+HxL8jBjnM2kX3BJwmT0qrwXA/TMeyfwh7N7J1C5J+A0W2YxyeTEDuU1RxZl+
asV7GVfJoSa9qFUtUBn63kPjjSYAJlZFcJolHRfbZJQnclRcZTvQFSp7zey1ZqVc
lnpG/WIEK/9Ze1N7RmsGZFBvUyF1Z/1+oaEbxPUsgSNFmJ4eWveSiFul3oX/iuAr
VhfjCY65VheBSDQIraXLdkuk/kVUP1bTmmEPbGGHdrgouKE1UHGHsd23yi0z+ktf
xUMGc/zGXsqmHayzr14PORhjMdAFLSSUdJXk9IObpI0XxPYv+eqN73S7v132bNVZ
3FC17T7P0qMKfzSBGT9Yfrn5AxFL9aUkemLr9zLigsg=
`protect END_PROTECTED
