`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IhAxFS7VXJj8KGK+jyyQ5PWdHPfjAj+o0y1F7G7N9ZJwYDSJdM3SDxH40XycjsUz
DECxMtm/4h9PlcWVORvC3A3BHvIgRpsjY/7/mwcHJ0rQ3Rs5ux+TkbOhECJ7H4hf
TlLzCMVQxW9hoquY7WyswoA4PqfELPyU1dZRdmrWfYCvCQNO2Gv0PIHwjzfUdQgg
j5ZCSCp8xKjWv8rU7l9nxJagIUvHARX2hUpAPXtPa5g76mg8Mz09JCTe5syNveSH
OjDdDNKBheecJwDTY5m40UG32kMce+5MvmJxuBNlV1sAKTHBkoLBIV3TE5KgF6kS
ACUJKU+bK6MNurOgh4j+gcatNTiPMNv0BASy9OIMuOnT+271xp+srOjwdttS9Sm8
X2MR+tEHiUOx7R4FUAAxhCTlc0MmaYbae4iwlK8iTqwqm2KwBbY1ROCGbAaenHHe
DEEPYS5uPiaNoNDuDaZKsCBCRxTUVhxfPgMpE+XGjGPTEmTuELSa8WMhjND/kIzW
Tu3BEv1uMIytYIv9Gq4aqEtMMZLqpJSh5LseGMNNTU//+Y5/gtU0zTrpVisWtiC5
Odmadeeih2njEpzimOuuvi7MxPFMR/QrSvYOQPEz6qqB8VxS9vIgMzkzLbr7NhP+
f4HPpC+yqjPPGTY9raK0NyySrx/75QgIUfIZ4MlV870=
`protect END_PROTECTED
