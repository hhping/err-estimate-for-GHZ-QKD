`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hh1xw8Tlym6+U9kE3m7np/maxu57vc5rQPxup2qJ2ZJ5zYTzOmDNgqaR/aJfYK/L
aml6kuRNc7pEcSxOBweSD/AlUaOeArXU+mSA9wwb2Ja1/iTsdKGiem4ohruwZs9S
K8urHr+zCj/EHxqtvpapEDnEmiZHjLk3iyTfCvvYk/8c3RQRVim8hzrVc/v2vkh8
FlvS5L1Lai084OUu0wsWPoubfKpFzthaQf1cHLvRNzw743GuBtmalElDylBsw3hO
RwoJopNWSZF0APncS0CghUUwTySKqKgXM4cSJWD3cRCdcQzgvX0nblQvJcqlhPKT
39wwZUTbwWfYiCY1uV+7koyURvyKLbcpuP+PJO0aZ7zFjW6DlV1EzUtzj9xs+scy
En+HMVaTnBWifwwyAi8ecpCl76toPhZpPLKiYvXjtUYpner3nd+9btbAKWgLuEKu
2X3nNfdcgga531x9mP5/n4b9widyhkA218ou3Xp8HW2lZAPZr0A+jCENIgSXsQ1g
R5T9dGa1OQOrZSkd/msdDS3HnYkZj+A2gApcYaXB+jvf2iPFrHMRpNKHYrm/wFE5
qOu4qh6BW5Y7gFzUAk3D6M3cCeJxBilEmhzoiX5M1xfLhNmWsrJ0s/+kAmZUI8cd
J8RQg6RbNIDuyeVg7WBFFRA7dulOzFw5MKOSkzl/UcjLeAHcuv42WojV5seMye+7
aEFZqcNBMmFIXFr6HwQ4VFhcUIEUIOCgr1Ts/foidsp/Cney+7wuXbCCdR4O7Lyt
6rJVJAGWhHQa8nomomlp88jTHixQ+QIVw6gTwALlirAIN5UVKwgMu2zGIFbETMPe
woDxfGtUJyaRW6rOj+iOObaZ5E02tLc2vQ1TvuXQ7O5kciegON9sGYODu1Ui60uv
vTzxhSxd4LX2CI/aHmChrA==
`protect END_PROTECTED
