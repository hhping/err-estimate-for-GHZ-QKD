`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Y0ZIE0ze3FgsAh4soXYCRVwG9VRaBrSsGykvvdys0ShdP9120LE8zVblK1N7RmG
oWJ1IxqClNqXWU/GYZpGcFZ2gFTAX93ufu4nMcOnIEqv8NYBnq0dxlkhpfv1JGLg
1Q7UjtYdu4JjTWw0XwMSmgxkdjmoKur6hLCxHih12SW3pAZ4eCQ6ZLtGzsdwgLFM
BTEMAMH+M0kUg/AGxCPPr9ENx8LELBmLclMX0inIUWZX+Dx591/NnswSXw2TGLf1
oy0Gdi8ZN+NPGixBoaDGKd3SUbczzppBdycvJkoVSL9N8ng7YyFbT+WWgk5Zfc38
qShN/HoQLsLsNKv5dQxQcke0Qomqntc6scv7HIleNkkrihx5rw9jVH0V4QnhFkrs
pPRVMxCA53EThAZGcoz5Hs4Jp4eYAx4tKozUZN1FQF0=
`protect END_PROTECTED
