`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5dDaz03Sj90Oj5ZHb8TAFzrFodHr0Byc+5oyuoz0+3PM7Casfb9rsgU1UALbVUFK
0iDN0Ad5XyGlcALYQ98uCOynA2f66EJbIPQ8gQOX9tOFj2itnTUsABpTJsobWrd7
oDp9HbymrAAH/VLZUUIMzV4v1OMd+sKKjxxXF+ono9OxZEzw04E9X56MkS3GdzsE
07SnKnUcD4MOZ90fgojpJ04YN+0g5DErfkDWKQi3+iCJOLcsDfAnBjmwlUdwNt1e
1g7oVOajyXUaMXs0x4KEA1A+qzU19gPWKKcbs51ilrdvdbSfAiEwQMfBHCwT/DuE
FD0loiqu5C0lHjVD1JFulni3uB37X7dJVxt8guaQCMFOTNIpleSXNuY7v2rvutsC
4j/25k6Xl1rAVV3JNflXtHwGAfe9MCUattaRkNrtoEhYATZhjJGo6ZvMWEHcmXRq
DM5Yoyie5xkOxT/vpAhl4Q/7T5fdpErfbqa+Gw8VnzEYXhz7gJbz3kNIlZn2NjcT
pR7MobuakB6pm+7sGRYEJ7FMvZ0nXZyg40Vh81CW8GJxty+0H0n3MzzDseRFMNDK
fKhjx0hcoY2hXDdhlC7X7FeDFIJ0Za7kY3r/C9JovpJi1/EWEWG5KkRPZ74IB1Rz
zGFh7UJass5egOiCG0wOyQ==
`protect END_PROTECTED
