`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cWOr+iZiI5j4ptvK0KkArIfHFEH57/ipGRGM/VNRt8sMS6AlKO7fj5r0LXsrE2dF
Cvnd6L/cgGjgmkQ4RpwaP00m7Xxx54xFYzH/vyyUnqIb8IULTRH99wRpBh0/Mgf7
1dPsAO+S2VlDh2fDuIsXLE1UHTz36/A84qhwYOG9oDvNL7+UhaYnB5biNxZcwaly
iBEPMiinTGFomsnVakfTRhDKPj2AM4G87jIQQKp8BwKtW4+aK9gBqfnTJUw7A7PK
Rnau7CvyIa+EQqzXNqwQho7mPvigfa0A3cZpn4/1mNWPGj44wGDJKA/uSCgMW+/4
f/uMkroDuGOV8kMau8WLDBnnA3LE8itoWdqeFfdYBxnzr679ISgVYWQEbcIozAsN
Z1jSlqZe11dhJl2ArjLr7crCqJtCTtYo6xp45y9XIdRa8RmimxuBJcvCDLqUrrID
OnjEbfRvxJr47nrvmaHfjuz49aX6sekZAtWVPwLs++1y4qF0dThTWdV7ElFKLCyu
pWAfWkkNYjvhEctInfUBJ1VqEq7XuHNAbLBuxL5+YwEKVG+Ah6zwcGYM/Re9Wuzb
mhQiD4nL4Qck4yHBP5upDe9r3KeoKv29TEo2jeBtNvOJo+QkiV1QT0hbBxBbUbX5
A54oKSFqIvYeyoKkXhHmYefQLf3GeeyW8lLQ5Rtuvoiinyelvez+S21f6I/2CDkJ
SIqA7uXmiN3XjHJFACrr/WauEGyLpQIAISrhTF9pAeEm8hJBtYwWQ7cRbHRGcFw6
xu/+Tf+ueKqoKDLOW8Yf2pIXTP39xl72iZyilpg6L4fzNvElC9U0cXVfMWJXlFGh
RWom82CTadxLY6Wgd1sr7X6qKIcp2LRTK4M6o241PwqOLTvlvWiZc8szL1E44F2Q
i967xcVO+LDpZ0AMFHhrViX7kI3t+TrHWmIlsLiUHpGbhszf4rECGmeq0jLym7wF
2YbekGfTVVENQuuHBd1U/8X77hELrGwqPHheDuwaaufU9lG0c9muVHAQWCArSUbe
gzL7uIu/KQVRree9Xm4RdByr3rW0A4TEvBKqbxCC9zqB8eJ8Kbc2MPHsJgDwmXJU
ctyT4X76V2EIaibyPOK/WWvj7/DR5JnZFPymIaOK8l/ORL1kNmSonE4p4odp/A2R
Yn8GJ4InbWJyifBd2oLwtc4ZxsNgq+cG4yi/p+cnajhYYAZ7Xw8NClsYfWPx0F6v
YQt2nIF2QF8dD+ivfbRzE88m/Myro474E1KjvbhZ+4Ximn3xR/cc87/azw6ghpVX
lxmPq8sgBaTzSnmzf6anBwhhcg5MvdCXhPnQr7185q4kkCQDTqt0L4b6Q6lBtDW9
Vk/ePxlRswJvHwcGOrzSits8ilAQnKesZEAIUoBX3Sl5DJWBbspfvDJn7KnBMsfp
zVcxsmdsx74aMNsAxoP8Sh2SyK+i4A+UXvVAkHfau8bC+yb17dZj5s6jM7QYhmr8
hnB903guIZmfL+NghZPmErfbMf+UGgLUYu5X0COFEW3ek1H1t8eziz0rRSEUI6t/
j6QKy/gkp02O9i4AHvreC9bjHRl3wUUWxi1bni7YhblpQP1hDWLb6p21iaQh7b5U
Df2g/JokwnDl2LwE5GFail9LlIyP1MFWFdJHlZq30uiTjjTH8o7mtvQBaff+glXI
6JM/OKQg+U8XdeOrbJakQbnIZ7QmFmkt6VWuUZgwWmI6Akf45gUMuHfjA8B7anR1
Qa4UkX7ehzSdCIZ43TkCZP+JgwyILNbx5Gnk8LEfyxBYOuF91LbJI0lhrB0D+McI
2Uvwy9XbeK6yK3fTeQUcVvXhAGhmeVgGEf7hWMnvczcXfDyJPphYHobvQx1056AF
5VE/ZxGsNYWqjF6b1zd6nBZ4H5i5gObPu3k4nbX4pD+isnK86FtRDxqIqlC6d1/x
cTIGoNuKO5qU3RSuA9R0edijjKXw/FH+2O1Pjt3Qyf+CcIyWUqKLJjeBhc6MnG05
XNVS6chEmuAY9c8WNyagbINwROTcW0qq4a3i3es7J8vFZhjK6dBI1la4isqsifmV
t4gIRP2gRm2F9kxY4avCONs90GZ1Hvg7Zmx4w49qKRHarPMOgJiiGshMD/AVEhSL
Zd6H4NqbByisF8bl9za5gVioEfQ52v/OIynJUqb5759m20z+QYNfD9vBwgNWO49F
ZZnMBPcwgzkDYJwulbI5OOZTfPAVDocsu0xb8I1xk6gpZk0IfI2LjOZuICKpeLC8
8Z2eM/mV+nX1WjmnXqogf0SFpKVZuKhGsDIpmUqwWXDEflk1ujeWfhnkaCVx80CL
K8v16q7Lt3s/pZx+KpLKFo0RqK2D48JH99K3qOYFn1aoIVOYI958XQ/uyX7/+2An
SFFR4u+MMBlXANswRP5lGgstDM0vs4WhfwP9kbb74boIOHmIyoQgRkWaId9zCUy3
Osmldd1oTwu09ooRCBbHqE0dgTZ6LqUKx8l78cUqpAcnOvZLeFDMQPd7JTB0yT2/
IYBq7NWcc/cxzVzfAyid/UpZSeqFfS5bRxuXawR/iWZoA8vV898QejnyqfL2E6ED
vih/mhdX/8w6ZDzvxxlG6ahNj+Qx+Psd42ICj3UCCjisSI6zWEfkIRqVL6XT0yZN
pd687wzmHMS2OI95ipRqdwQ14mWa9AfyMG5AaXorpxH5bm89XZoWCSj7E3eP96GQ
S3A0jYSj4TGpEa01UyKrKWUvQyDZIcr+CN/AkeVuqaz8eRX0CsJFqTnKVB5sAOZt
82MXWO9QR/6OG4vsqdV8F6EYoDUDbwNFCzTLjSzFyVzSxFivSa/s54qe39xviBoU
Il+jwBVS460eXKvBXudJAgWi8PBDxldiH5WTZqqx2MLoITtBT18e1eXostOwOuuB
EuZEfORfYo9MVMgRiCuZUMhNo2oh8wwe4qqBtGh2GleT+HWJB9T/DzhFJQo18QVm
7OooNfD89X8Zwx649Nsq5vhQjB6MDQNrJ/jfRvOYgT4ZZ/28ItQT1pbJNMEbfN6q
+uRtuvVPU59a2SdZDzPRGiOsUAvTRGWCOppidZT4DyfSRAtzO3isA4oyINYTpTKH
DsoUk3k1yOYeGRUyuUXxu6+1rlL1hCM74uA37DjggO29SLmjiEVpTmqMYvJGJIFz
Tdc1ywj791kB9rowVyagCNHbF/nxu0ed5bJk/by7aLErxsqx3ppxiq8vVjPyQhQw
yX6L4Oe3cO3cFoE5qEayQekXEp0/vbXFSFfokgszZGhTl9MGRrL26g6KdXGTSNCu
ZT5+bUjkZx2RduPOPTidnlpUgbVpi39drXk23FLWKASrLx7QIbhO7ngm/XTq/a0d
lOF+lpMl4zR1/5ScWkv+SsyaTL4OlkKrckrWRybbX2xNJCzSuzI+Om/fGKftmqYZ
bR/o4d/w9f6EQdEF1c8MtNI98yF5kwrOweBZJ1bKVS16/4Lg3aOeL/Yi2Np1dLJ6
PbyexaSShoE3ZtG99vSU8g==
`protect END_PROTECTED
