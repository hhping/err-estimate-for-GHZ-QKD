`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h68spAkGpxvTnGqoIUTj+pcwOZZyo74GgZuj1Z86Zsf4eJvC6vRU/m0n4lPEBJQ4
b8E9yXd+kteUL5oKP5i877eOug6fyRqScdslRTXSS/xB8LI8wDYLV/MrkRhav6R1
siRHSSkztG1F91DUfEwr+/VmJscl1A1TlCYMzS8P5I67RUdJsBo/9XfmCl5lzJgV
853uXYP+Aq239cPooUsjbm40cdg5GnhtOaED6XW8ncMTJr4b/i29dLEDHSbhSVUg
XnSDT1bN5iWkunuHbOAPBOwipYJR4tdT+edBh7x7r41p+KclepDM5LI2f26iDOmf
XOajyVeD2aMpf+/BAHWWM0iCDOcFfYY7HA9Jkkbvvh6c4Cr5KuMnMMG14B598o4C
5u9eQYZ7QxVpA0+vbJl+ZwuATrPlx1BuaJlHv/Stzo45KF4b/VmjS851LvtLhL//
UZVzWoS0e4i5N56BglQaR5IHDYjqDdPZMyLUhj4TQJ9YNM1t6ESFNxECGaeGIGyR
Ka6iHBe6zqHYN+QuZlwwTmHpPWLXMsvWdHW+5mS75QNvLH+3GNo/yimVBOdTCgSX
ORaiPILsZV/ireN9TW9D+o7ngE34jBsYkC0+hf8vF/AsSkbjuNL33pushmA3pxD9
12rFvqbAGl90A06x8CQrmBnbXh5tQ1zvTDpm3eVF7DyvnKJBEckuK+kBIj6jZHda
PI/8nL7cbvxMZSjgO4zePImvsVcqPtJSYLB1mgur/3KUbpGG+WCUawNtvJ4/s64o
vKgJjkFbMS1Q3b1rROfuzftt9dZHHyQ4E03EbTiB6QIBAAQJNgU2rA0Z7yDA9DVm
vzJQd28KuGsdu4JoK4gmZ6jL59kfNWn1KaC/xcc31kK+kvsjIe3s2Pyq4BewmpsG
ri8b6pDc0yGFIA6yf3T74wNWp/PbdzMwukIjlMu94vugMwa3gcKUSQPWgjFlHSUJ
7gDUt8OBdQmes5PcHOhzO14tZCPWY6fQHRrXeFLB+ZrouZOAeO5QMyrZbbA9tKGM
HVF23N0V/IvUOOHDACtcQvOFRGHPIaLqcSFPhorbsCXlZ1hfLD3c58yYsXbuo2qO
MQGD+hF+F9r+nWI97qa9YHRq4304nNASlOXfv95PHCYVClsqhxkMQZB5l5WGHsam
babQFGiHFyHSAnd5Ndq3bYCMY8VXn9xLcJHm8+UrIcGFDXyQyGUdRn5MzR1/jH6c
y+d1TSWFZ5qqlrXJOAPekA9YSOibZoQmoZSx71vSWND5srmqKZl6PaLTH6ALGBos
i+PrUT7KbtOMgf4mqnPcFXCZC4qfltKlhQ/DoiOi3es=
`protect END_PROTECTED
