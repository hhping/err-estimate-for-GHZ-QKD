`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FklxL3o85nEMYHT4ZFmhyL7CkAH6RIBwowQaJgiUMGXb2cdfU597KAROJFFlEJhX
81EV8CubAmmoMWcIBuUxj8lOGTDbSE2fHA76nCo2mIIrEKNT2u+2KTsvk3mWKN/X
hoyiF0CxL+hFtuGbNB6jFT0ZHZbjQilaC7m/9cVkA4zoQe+l4MtMNKH0+ZN2WO3k
WHrDSrixTREa/fd2UayRmdcMDUOq7eOM6fuYo87j3p4dmXj2VnwBI/K05/ZSo4vr
Y5DWC9ee5cYJt9UiQCyFcYDgF3wF0HQaNNY+okWwLKVJrsVJylRGIM6QjHPmVoeh
gOjTxClioTKvOql37+gsVADoskEpsUO1HntXZeh0u46PNoeMnoGAXyZP4LSip5G0
G28QDLq6hpMb4tk/3ZScqxk4mgT+c+2smz2fPyH79gWnOx3Wzj1ChUwRhkHfPuiK
X/KnOrdeoldkkmfeBWaKqCVACdJkLEWCs0/Tz2cLkX+GH2+wgTmJIToj177Azd8q
eqAckvFOwaiKzUUJnPeE5DJ8w6jdANvNAUpeHvxai808I4/iutGMcC1E9pup73a9
qASA1Yloxksz/Mduk98uW9q+s4duIGLfN1V+y/z8UaDmN3gmrjHXV+U0fsgUVgQ5
S5LSg5e1YdUitUNK9LSpt2ZibixD085fcz2Jit5cEP5W6+nXaX5kLNJTegIWjhQP
2kEICnK/G8OPkCX8WiQSOmIn56MpHxinY6Fu5vhNtLqDmfUWfeEnfvLsR+tTFD74
SV/sXYJ6Mz4WpIsT2BAudFRH92Wg/dF1/1cukscpU+wQkxFHKG46cNTJVh7ZMB52
o0A6OTdP/SBIvXwtaL9P3L79r1r7AfhEa8zrIDnxCZgFJgxDrHl4pIz8PG/amOk0
vSZlMCF2aqyNPWXEZLiyOSEHVTfxNPdEkThhl2c7z0oHpURXZGMoNWj7ghI5EwS/
0QI+uQct9DFBvxCk99XIaEbpg7q9sr7+73tbY7gtMuxa3oPVSmENGhG3t39+jcgv
HJjCzUIQC1y5QNZA5aWiKZZCLKmiWmRowxjvg1IKr/yX/vQzqEVlBmJv3jp5rfSv
VwjtmA5WVc8pHaxLQ2g+jHUe8ScVPqpILVKq6xF/ucQ7/soR+FZE0KXf2evkwJ/i
XPnj+wY5RmpuM2cZmxB+u6RnZIGSG8eCBxkg9pxPKybCbszEIpnFHjsgK68ZKkkl
pHAMi4QFYgershFenG06RPC4w7H/KI+CTXQ2NnXJ0fMpyxaPi7hK4Gu2+aTKb5vD
Jj8MZpCZnT0nmdqP18y5Mg==
`protect END_PROTECTED
