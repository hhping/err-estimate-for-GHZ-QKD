`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aWSWJvIejEYdpehdsuJ+k+//FzxY4Y6KvPJ2Chg3oLdZ631ULSpVxKw4ptW129Vh
INv7h/AfffgZiMehkFzXNrLcEVi4CYP+jnxCiNZOTCtkIcAvZuZUr8+6apbCaNwV
e8dG9LAyQFfb9T9b86pSpgE8vzH5ZC5XNkQXUV19pZpqoC7Iy7S++AlUTBFuJv5A
ei7LcBlnhloucojGa2M13Y280WXtsQQPywmjpy+JP+THA+VN2Vln5QlJBzkoKigV
LBqUeEHb4u64wATwTsCDn1Fh640jv/IQQihVyCdWod14W9sFkopkntg8ICsalD8P
AwZKJrtkFjOK9eCS4RcRaJN8GDC4rQoXz9xOvF4gjt0luA1h+dIV5xLo32D4s2su
XiMGa09COMU3UIpfhxOAVbb9qDp6UmQPIkT7Ino+PpkkU6g5aR/gloZ0YAtyRZtn
po3Z0uy+dT50E9hFU13zEJuk5onRIGwJbZh38lAMZhVBmTUepLMmX4rCXtE3dbqA
T48DUh13jTFkWMovpWyWxwr6SMCvL4ngH6svGbN/wv4ih5DA/0Ovf/1wZbDyQV6d
IhdnY/NhG/npDZextZu2Rr+NNUpiqduXiEyStoARr9CnN5VQGocWCz7c+8bsFTBr
Fx9fVsQDprz5N06i76k1oHAjKuBBCp3CJZHFS7yv1gw1JfUV5YNlSHT8WrL754tP
VtqIsEeQyR0CaZ/mq+ZA07fn7aA+WkHxL2JwyB6p81VazKc4CoQzCfTTena/wU21
6aXgQ7xcRPVtoQLh+hzgqf4OIRz+pfimS3wdaDWHAMXsoToHHTYiMoPwzXrqPa+Z
`protect END_PROTECTED
