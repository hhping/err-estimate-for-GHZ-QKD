`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q5Jfjr77ji8/VzITU+mW2R77jSAc0hdUZV5rfppBRkKnMZJrR5HYHHf101+ufkZB
67eQ64UbzTZpVOn8BNqXyqQ/tQse67GkscL0tLeEdid3vwuc7R1XJjXCX/BF0Gyx
1iVYG45HDJYfbpj840e+/sQQsIJz2RVSIP1GdIadIhe0lmZVXY7SLPdZDY0k4ol6
jRw3vS8lT4x9oKINqr0h8hvUMIuqNQ7c9LU2JZ6O9PtqvmmJXql8wXZCRfQn8da5
3HErKsw+kayjw4p0+7+ER16KgLrqiVkLhZbwNeNJskQqRFfRAsOHmF3GIyPtGFJy
DguSm0QNxSXr8C5gzC7OIS6Jbk49obVsjooA81HC1kEgHxot10nxIAASJAMpI7lt
yn/bU3fDh6mfAwbUmTAQb6lGzpDZmcTdw2bhT1EL/j9LSoOA+71KL7pNzb35/rIX
8S0DSp3h4RCmHFjtHpLxf6vmBW4qr7w2Rkc0nAqB9yHDQFLt2SB+JuHCPdFIEER5
5NUqd2dbnAquYkMDoveD5AWQ3l5+ui78/0/VTZrZ4PsYtLIrGX4w8qSDcLs4hRgD
nLMFGImIRc9B7EOISXqzMDV4AZGk9PlJqMvvHJr867TJY9yp7Mg3z2dfJFwiDH9e
GDDpO55F2CfFt23vj/N7SbtAzhxS44k00ftU+ejaHyMx5uI3GkMAGIBPOsnk0p/f
aqDj8urVqbH/ci6j6wmlHu7dGAzmwOAp1yz2YNzjyEwMMhQf6eREEX+OIID7vnzE
XQLc9zx6jyMjvvMfcuGfccwFcSSlkiHkJ2CdAjZ1pj1grT/3sEESCt6+xaOpK+JU
kSR2PtVLi0neCKeAERGAYUI2DsWprafWMElToqzBz3VWvLvaY5RcKNzVcDTiVnV7
BqaRVEkEU1TL0wP/HtmB3cAnwAfP1nfftopev16QEDqL4+CsMkodtda71WATR7cn
VsW2eJTj1zzxXQ4u2FPcxNYC4o+xIi0GIBtgmAbrVLkwPOpuoEl/N/C2nlRE7+bU
uYaacodmYm6vBkOYN6WYQOz+nRF7z+vH5VaO+OoNhVDf672UzBHjE9+C/fcj2NLM
nuFEvodbKaBOyq88+TOkGzDuEpgb5b3JEhKla5AXwIuTUP/X1dVsAHW0euQ1pLvs
N/mNPCW6n0fVAK3KcwpR9XWmRx7kXJ3JAS7gdyrhu4BHbQqyEMWoxzTkIalx8lO0
IgpoqZzH4bic6R+vaGlZmJKRAzprzv2aVNcS4wD+IYoC4FueUB+md7chet7bqFbQ
vbBDH90+Y1RnGhLFFApXzMf/cBDQlns4gnrW22ncd/qnuqhQcpqDOiAIPYnr4r4I
8utZljBGUFg/b62MVq4Q37JyNPrzFiOgwsTh7YxeDwW8j3BOzPyRDtDHR3hcQkfH
wSRmS0hR4w6uI227plnFWKNE/rH/XZkCrn299vZoIBQpIOmqtmRKNCFI3rj8jA2n
zDwxfBo54ckpxaqKDTjTHQ==
`protect END_PROTECTED
