`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+lL1QUH+G1D9gmXU3+0SeL97kATlTvTPaG7/6TkSjnOCUmWJ9aycEFC4uduXEpI3
bkxvz71sQvlgg4MHIRYhzIrpHgiF4JTdQRRNsAPdotizXSQTBjpE9nouv8Ulk+hz
OgI9GrOEm+VzVvIEExBz56AwcmgdFyF1b2B4xMpcU2kOngkwQ+3j+bMy8UD0/RZ0
wObfuBGHraCia/nDo2J0fVzu4xpqIqAgsymlryY1DILS7b4pApLpOwWX+GnMok6a
2WnhRqeCmKIEogDN5b+O+vUIn1CbqYxsFtMsChG3dFMQnH02Pt+CD8teiVmRBuxG
7WO0Bl4jHoMcyF5y2+YDJwpk7BN/NGtdR4oDoDZGz+WDHn6Bt5MVnFo+Tk4VSsMe
//yabSpFpSxkicb6rFaXMeQzT8EPGFFuXotu/ExiLSA62NyfMH+ILE28YfH3P3bV
QBStJr2QAyn6C10XreMUx6tbctygTKwP/b5B2TsGodENryqjmuy88qeP+WQflU6l
PIKkvn6gHlDjat35mO2nn2O6fyJj60MRIoBXxy1bsiCo5LcsjSUEwKi/7g4bH5Ie
WrgAdWxhm4BEl4SgwJCU+3wGHoj940LNKcyYV2d3Ys2d+JBmYSPL8z/mzEYVvGSi
YIIKdNj+ZLMyOZ7qFlGdeXhasHHOydqEAvpu8DYx61wTOJcPIlsA9LfQ7+4DmtWk
n7tCsnKx6EdvGnAo2+ZGuSkp3uN3J2dXdm3Zlfxmtrx7bKEXIwNbvu3E8RU2ElSn
gDlWMctzi4JTC320OvfDklx5stguuEvc9Eg0iTTFYcs=
`protect END_PROTECTED
