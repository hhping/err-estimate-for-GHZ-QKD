`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kvf5S4DUwQcU3+Kzo0kb7zAKls0tWExHgmaXmt1vALoqZfQU7QYuP+FKz7W1zUyK
kDMFnuOF8GH6DgemAXq91st4jwhELSmSoSY41H3aQcQI29fN2j6utwfhDUBVCJqH
EznmLiUwuK4qFXJqu//WhZUKqcqgQ66nVGFv9u5aCNERvni+P251U8vpKkxtr/8I
O6MLvOi13P1e7PKuT0340DxGBrInva50k97k4+ZXI9NUJ3S6KFMTgI5acTRXAEpZ
i1cQbuQJvXRkjYICC7WLva9gn/RFPvkVlVNT9/9tXSqQ6OVm4Lk9s/O2gBcFww16
MXiXkGoFt3n4q9jpr5zzWaUuE5aFxSvKvKi06oU7r90kytsP/xdgP3FQMPSCEmuz
BAmHj4fQtufEQcU0MZZFuOXqfYWnvxy3BBJcyqrwt+q9Jr+OUrKhmvxKunbK8HK2
lV+pctG0m4/bZ4QO77bRApItgJ1eLZ3vqrGJAlkEjuh1csanGDDmas0PTe/Bhlyo
g1Yl7apr0PAyS0WAH2bptfrrr/gGfBYmc/C9A9cwjsQVG/KZc21Sljcclc5bWgUB
sDRHki2pUzh/N9iLJ0R6V0PaM9APC9p+NFE4mgnBw1rx3UseXlw8YkLYHdV3bzeD
WVYueu7akfUMv794sZ+LqQg03L95SfbuOQdjum6I5Lhij1UU/JJ0P0wcTJ287nUx
fWuK1onoZDkV5Qbq/u7zCSahMWE658l2pWw2cy/LRk7AajEM1lubyunyEImdui71
KH2R8VRRBxhs28lGrkIArjB1Rst+55LruEKHh5d5+/NcJMBoIVgHp5qV+HwkjMSM
v5FP1kDasH/c242yiT+a9Ob/frkr8ybxU0ZZLIxgKNRSnxRqcxVv64faiHIKyUyM
lA4hwyVMIvN4X81EuChsYi5pUH+CaW8qjJ6BbXu8J0T4/UhZGgGsOeE8IYlkorGk
IROibBb9olde7vZiOhwRwb51rURl/TNyfV9YFsXYBcJ6jMEJJUnBeVIMAGZVGHa7
RQQYwg2cIC5LxowHYUISq3aYoZvMzAtPVCNNoMmsGRxOkH8retEFkf65gzlrXnLs
I5s9o9Vheyhtz0TFxi7yQ+Ly6xNkX8DWxTsJriWmTilJnQboVpZ23ZAXuFfAfJaT
n8bdhhjVjGCslvBbT7ocLzlusw/SziUmFfLQjUNgJ69V2X1QpZw31OXhXOHUHFqm
Y7PHHIA9cLPinv6aVuzJB4+GdjQbEiavZC5Uz3sQSqMxGhOe6t+FswYKO3UHsOKn
4ttn2SSqTj6Uzux2alDZNgM+YhDTdDM01upz8cEmh+M6eP9wMWnNKen9RMYh3IrU
yn/OQN0OHBYsXiRQnZ3Qd9cBUgJ+IRZznjsC0sblfUUXmtVAxRbrQA6ts9eawY97
PFTLWb5mfB0SvcpQPfL7hE1QBZtxYozh47cAc1/sDVBXuK42AbxquGF+BzrKesHS
T7Z6L3cE0t5yRfy3XuvAJ9uF4mQ+C4EGj6VsYIc/ZGJ8RMt6ROxaRLy+Cj8zPKOg
XECAr3BZWcoPbGywM644zl782SFT3akn1W/MB94OqEda4LkmCpPsm9/62YUbbkJ6
QTd4Iisbr57qFF6Fec11gcQjVeuPlQDNf1a5TJrHJVcgPASuSNr+TjbR4QFp5Uzt
YIp9L4Qtxr9lWPf8HuDKyB9dM7jzxyBnm99qF1wLMJnKl7VRbgYwwMhgx/zLunCL
v6s2F9ewLJXBzO+fM0TwUU4Boen6ASmlNfVRx+6Ngo0SP0F9navo4FofX0xgsQ/H
9zDNj3uAjoM4klO9RrvfcTE5Tytika+8D8s6q7VLVaMAW3oI8tRmnWuQDFd674oV
qMptR8jwFj/MVEhs2xu0Vx52bUbExaVEIu6c4hhplTCsphQ2wt0kvB3p9degMsz9
hGfUp4xtay1+t3uzY9VAdefUnwDEQK24HfVUVzj19ybb5FQXcnhwl36IunA3hKsI
cgomFku3+ZL21lCndfwi6uKBDwzAS8aXsIYcNmVKx/gy9EigOaw4mKSyN3l2g0ER
wuLXoWzKgQFgDNv/c8E6YVyg7HFsh1sJIdsvTRw7w75yJHcMcFLoVW8KnANzIPrw
B00+bVZzoekyAEBMj4P4RlFnH1xTGtGnNiqDa+Ctr/aKNuS4RmnmZ4XqY5WyWwsf
WJ/1RSS7zkgTXHvjXO9Z3Gj+GZ2aB8RyAUu+3QYRaVONaTKhBRYODHoemz1y1cmV
qW38fWZH7Y79JUGu++AotWXmEjYRncNKmQILQZ1jVwYOS0lvTkmXC3kJN0qhi7J/
u4lZACaFR8yKCQvB0O1dDUtYdhvUblkvINctzL2rKiXgZEmvz80UjRoKPgsXa7be
sOdi0ms+GuRw/MnVnwLKXFNZrY5r94awQUuAjWz4wfsfCSTf1KGJbT1Fr4dxYdAI
PP0UC98SpFyhngxkUsyQ4CoI3/V+/8WzS38py+6dTwHpMAZpGDE4JhoCj5yaLnnV
WC8TdKoFSxVf84cupn3XOaLr++7PX1FaUFbbjYs/Wz+yJTIR2+PA7/8MYp5GyYSf
21rGk+t0Oao4d443B471hCd+TgwTgaNKQ+MzmW83nmNATRDuzG/plTHCiu15KPv8
xuj2LXUC2UWN3FjvqpWf3DMu2uWg2OjC3z/51sQFdjMa/ondEJfcGx7vlP0DkziB
W5hbx30R26nF1SsgY1lulEx8sosXyHGld6X8wvgZbRdCf6riS6y+F49qVnG8QCU8
zOj4EyGaqburH3gWCqvbKG1XspmLcfyCr9h3hhJk74pNJVGArNtz647TwCZZDp57
hW8VbF7VKO5c0sHxUH5ttzol4KSxxO8kxyddnnNK4jtNmLK1WEKu0t/1k6RASWgS
8+ZQGlxHrt87veAcWkh67O07wpFYrzzTh3ZaxgsdWxfYUZAoZ+DR/RsXc8kHn9vj
rLRNuAWVTsn9QGbG7icgNn2FtItj8lbyBkRuwstMwU9JRr1OxWNarr3E3vMqJh4t
jksXvMod/VsdcWkFD3pnDtThaj9G//PnPCHtOu8eDwuiWxsIpk0KjFafV7IBebLN
3p54MtGyeOAAtUe3ATYERlMKK0uZFEpRQJl//1prS0o+zFk/3p2waIF32nnuWeWx
TEvmdJfswjNuTd9Nv2tptY0iGjr27/HchNBHnvSyYUmyI5SM4+O/H40tUKZ6cHwT
mXl4YS5diQtqzsjWgT5osgpGeadx8IgGk45QR583nJQlqJ8BBlX4trifoBjIa2Yf
xogP4c02BNt5bvXPbtVMfGN/AvFZ6u6bxay684tgMDcGkeiVoOOniyJkbJVyJvKh
wtCMYI3gRyfNOvxT1Z7CcKm8BG44nO+wLOYeo+EfRvvo00z7LGiVHlPmZDlKR/5d
IHVoqy+vvCoDmT4yM2ajuwWj9UxTz5hbsT5ncNrbi9v+cPlinmL3vw25DMRC7uMr
nJWgAxDxywOxgVjQMlOzAJwEgwS+fRrEwLiN0D3Y+X1iNKfIZn8jABiaMeVb/4lF
U+Elot03ID62LCUcnwp2GMHf4gCHWulVKRrtZaBPYmPmwLzWyxotAgJtCgDDaW3Y
UxDOLQKJGpeMR4Zp38pKE5XOEpA0KXw1yJl3OOEGx+L5Sqa7KTnxj0N9dcmAmWcL
Fd2Q/cOqZ1dd8+ipFr5L1miSrjrIY78HS/4Ifx+BiLv7wSgB3NSExIjJ3uxSnoD+
KmLWH38bt6AZ1xO+hJvEKciyMgWyHH1irDwmZ+xEPLbqYnQN5gJFyeQ6mV+vD3N4
q70YP5w6sdrzqkc+OZ7XgFBfwL3PauseV+ek01T83lcUJhfyE+W1YEREc5/6iZnV
N01qjAnXStwAB088rgYhxc0PtgwPr6qqyAzz7gZtMZX3dDQU8A5AQv7mDbaGW7tX
4VNZSg5QKOUdDGHvJ5mRTrnfEriKEbOxwO/TkjaAPuUQhDnJt/41IV732B86QOhx
uMZETuUZeUqGNWUCb0q5pRrKSqp9IkFF5gdii4pv70MargwW8kgOVhGe6MBouupn
r29gYB+XuvWgEoIr0DcrJ6cT8gUhCb5i54T8YPvuYaaZG7og++Z2xxbL72PPAShG
afQ4VTLvdBIDL4qy07vO9aKF0urbllV2oYE0v3UDr7pagyfeCc8fQgRTKmc06lKf
+Kk0gaBYaSb0z6gzMj/N1bJZzPEPcMrb/0tZBkz5Db+Wh8/8msa/A67G3b9QJd2L
fMqNC2hXh/nYNgxttqhmbGOOGPozL9cGy1rMSnTXaPGo/DaWSq9Q9N3+uzhqfq3/
4jdt0F0OyOoH9FbDC5ZmGCfMpvf1h4oJkZ5nLmbaz7bp7y1igznp0HwWcBOSUTpe
z6d6DDLJzW5hgElIWTjsN8RGomfXlTK8vG4AtUzYuIxYOm2+DRo+qzAWGpwzHgOY
4n0qk0GMB6+piFh9tzlCc0mQvzRnYROp4SpBdr5BW/wlG6A3IwxJ11CXRVY1Q2oM
kj0qBVSxH3d9yr/Mv/lBdmCfcgCqtAAE2rTsTnKNkFsfRTv5UO0Xw9UHAgaw1Ayx
nF3OECTy67ZkfR4o9zBy4k7cnIV1bUT+3LfS5FM1D6qOV46z89CZavXFH9u1y+Wd
VCpe3R/U0scW5BVjvKaAaJh0lozOI/y0fPgqXf9MnWeNQvUNYg0RPBwL0ra7liuS
pgI9ik8LIw90S6kMa8gUPZRxySYpG5TwiqavgC1npgnZVkYQPE1q3D40HqsWARCy
3eUdNPirq6UIlSJ2do/Mqq7ED9S0kFN43Rimf1PuqdPSozf5HlzKPJZ6Vt70aNd/
TQxqx2XzXjhcp3uoTcRSaAyTEZ6BD+MDoP66I1oSTlTKVVlCDw91QkdHp6PsRo5d
d8tojjOA4U7SHhEiXcCNNxOqGyfhqDOQa1zCe30Os0TD07U6q31BkNO+aS5jb5yR
NC5bUt6KRA9bHFzIzzUzsUcqyIHGcn0SJwK+uoQ7xA+dy9UCLTaF/N2sPN1YWl1u
lDsohp8EMuahjblqVZr6BS/V61XiY2MmRzqUvR5yZxANy7TePI2YoNFALyjsoAI6
Z6ubeamJhHoQ50OcHbX8vxT4yKK6kRx4HgAoDvFFD6jeRgI9Q5gBdnKcNvzlJ8g5
EaEL9FO6NCKmk369TATjRtg0G78F9BRvDjkX4LyFw66uVKJET1cW4jStYFyowJMh
T/Z45mVzjAR+6VOBbEYd0BMvnor3P2iix3of9oAxDfW4K0IWnYbnTne487h3I/Mz
8pIUcWBY+Y5zgTUbB11jScPEJ6DuoXvyyHtEY9mxCWauVyKp5NwjLEUPS2RlR8a6
BCdjtxmQKXkl6A2LJT+sbDiJOhlHP6wI3gqFoL5ezhtzvqS8BGFmRf0IXUC0dCuI
rE14FKLKUy3f+Yyp5kK/466eYcuZpIXCYh9CkfIWaWkYdeQFv18FTLjJ95f0kYgC
ElWOm3Mbw+TPqQ0G/uZUoZOHhuTB1eESnkYv8fE5Py1ehaEon0sxdq/0JirA2n07
lYipWCXF6mmRdUKYAvRuvXbDdRR/5l3b9QqM4r7kMww6GKzl10Md4Okxs+ir+ehC
TMSuC15TsGHAtluZjusEm29PtL2Bv/vyuEQV9AbKJuQ4/tCjlqiLaA54lNF+jWLK
ptOi49Ozq+3wEm9aoSyn6AujqGTLVsAXK+9Ukdz4h7KtrvRUMELLD8i7wmOFBXBh
a8ma5kH4EaUuzFzinE23simHLJxxIgE/dDAXWXvZaKvMSsnYtbB/3CnYjlFtet+i
OD3ujMTwLKEvN1+Scpbe5mKfRwsqA9yju/y46Vu+QCLhCLpT6EbQP+UwI4x6hDMn
VLmGubQ9OwaqCcnxg8FDSBHoSEHJhvtRC4No00SJA77sVRJMYD7WdrvNXyUi8BFB
`protect END_PROTECTED
