`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BdNsh/jHhkoPJqcfWSJhUIk0fh4kuBCwQe2TceAwgi2ojiLYS072adKJV+1rMfdc
igIv7zC5+IAGjPIKOqGEs3qMaBCtTLSTN8XtmdXQQD/ctpMsPqEOXxd3uaMOdQUF
i0NLs6ByX6UkK9L81dl5pkY88Vv6bxXF0MO3ABk+V4VGmgnRZ24jO1+BMmiN9RUj
fPjZDNMIWOzm6/2Qlhg4xiOiFKGCr55cY8lMiQFQETRtNejEZe3ffU+VntCzOS5W
NmX2hk61lV0NykHgpx1U2bRuZIdEHpBDM0JTfduqXuawtjR33D1+aMGkU2BazIiv
cZ0TGbyhgDlzqNNfN4szrW/onbTNks4QmbUpOajV/SMUwjSrAC+48QzWP/0bVkWg
eTBWlLyb/y/cpEj/vAx1lqj0GP8fOUWBXxjpgVJWjJE3W1BUjddAXkpXESYui0IO
Tdcn01bhm8F+RzlJSzg5gokH+CWto8bPEw8PkYAYceSDWbARwSmmZ+LFOYrVOeYC
1czLnDM8G6iYJQHseR4wTwYDbzCzkYlA5YRyRC0Orso5jrWpcDJj5ibgZX6oKjO6
vxjJDlJheXKlBUUx9FFaG6Q/FVecAr9T8NnPqkNk6zUk0kNON0rcRirITOtDQBTW
YRUVnoa0HAl/IccRKl7QDX7dwboPBXFadbLXY164szjf9+ykQxAPB5MT+dabnPFZ
R6Ss/UrpyCMGB232NyjPEp9acOENL22DBR4PUsAcQs3pnPV1qx5CNN/mPSNJ3gOh
yAZ3WIBXne7iPDrT3B22h4I3i5qKmEXRtAPO0gjkZXArpdfCtjSTdDgLujF+2+ez
8QBkQK8SfT+edy/xAag9AXd5JGCsPMeEEkVnQ3C2uFMtjSlU8vtUMMUdPj2xj9e/
L5EJgSr2mnVzV/mR6rn5qB2j3oOSCe8DNF3O3/aqHuMdnrVZZtJGSze2k8EN2C6g
mXl3eFxfI8pDBJymMZ1nayHxgTKlrRo1RjpNE4Iml1V5PRYFPL8p5HWbjfXkW5Sq
/8eqVwcijoq8pKyk6KeJ5CalVTKjBp92ZNpEGyXKgrMV3XkdwpvxCDxYtEesW9A5
2l0mHfU6WM8xWjnAw586gt2U+G1g7B6rrJDG6QZmON4rCYhuZ2i8PfLT/nQcC/WV
m9xRjkorcevy6uXZmNTvuJY+VKvP2Kvf8XUH6ErNoOcGfF4/HiIEZxl1u2SoiT6R
ZxkiciBSjtyEnXZH5S3sj4d2SQgdBkIhXwweeJu6WjQW4P5EQeu36FApEqvY5EHx
3QuuY/cLvWIzTOX3j92OvgmipFKAz/ET8Yh+n/FsxpRK7SkjI539KGF4Twga/ECN
Nvle5fSvQGTcTddkE3CWkTE9clwNVWkh61rT+02qhA8pTLRCAdlCIMm1kV97lfb4
1+wlyvL7qdb8W0ND5mrNbHOz7ImsrgYAQ5E5pKEqt4vDwcaBd0VxiHjDS+SRcF3C
W1+sxdRbiyxD8FJ2Uv9ZO4cEFt5/4yFDtU4S+F694tSYuTM0z6kltLLwXLWpsfU9
L4BjJobqJTnmFPgky2G1pbkdqFlzombKvYxJBNuWrhOkmoDR3ci3cbrc9mQQz+5t
oTZRymeC1ZCLJWILTxDcKO0NJBKYmyN8w21OCEf2VzJLHemk1dJ5N3mZj3DECFAv
85HCUVtBkvInlhpnSK1ZqB3/PGhvsYkz0H4LtfmKBN0i3u/xRdSGzpku+1XcuanL
1Uhyhg2I1FKM4A5In1k4OzHPQWo1fFjdQJSwIRbNJ3r6EanShp1TDoapjBuqVPAn
IyKvwpR9BaJD2O9eqG8F53pXdWquhbPKjimn3qlmbivCsYj0BLYXF/k+iufKOi8D
bmyRlaioofJ57fVEHtSPn32/VUUvk4g+W3Ar6J42v4ERjRZ/aBwInWRvdWBpYCeV
Cg7OUtcNXXigAWy5xY90oRz28LhZQ+csi6AE3SqVBCSMrLRdow+sqxmspKrXe1wg
BCWDi64rPH75HjKs3xXIpcSYPgJjKodE3BfGc7rjN4RgF5OT8xi7i8gmYEv0VuF8
N4+tC3Me2UpdNRREbBmHZw==
`protect END_PROTECTED
