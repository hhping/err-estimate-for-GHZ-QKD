`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UC2gZV/jMtNUDvR1i8VjVm1oUFXRGxXx6TnTinArv1ljOlDV33eBtO2vNZYGpbR+
Z/6fq/iXryEv/GM/paMV2k6KiEZYqQNAfzn2hHYqQWO1NP5B4HWKr9iEtwhEQ8lH
bQCLnfQwJFJtWXv6N50jXwDwGuOxpWnKkx+lCTVQGo6PFPaugCxG5TZi7Bf/QIqw
TkJjuo1k2IoyOO3qwC8zQBOYjtcpLawDLHynRwSyrnXN9JD1XRdj43PbIjuJANao
r6MWERUidu3WtZ6cibxw12fwFhA3KbgLD6oTAyvleW7LTb8LTRtlSYWStD/WfZ/L
0peJhcMqXNvG3BOffhNEc3rDa+lVjGxtMnmb1Ipw3bJ4OapmDCbJ4ChvtbgNUVeK
jYn6pbXFnWe8B45TttMvo2GESE+K09EHP243OFV4iADxacKF7h9V+1SFskYiI9ih
R0ddFKKVhYy1RpvulODcTBowMtlNoGTsWUwCxgvVSMDV/AiGmQLuSt2LF/OtGGGB
aKTZmvS91Zt1UHp7PeJeqhFAq4tIdzEICHOTUKd6NEC4C49dypUdsDUUBO18Cplg
Y9tRH7oR18qozDGADOLQDajd5dfJJ2fQdQw74jlYvOkyfVAciwFWIwPALuvwdQy4
+H7bosNtZWN3R2KrBVBiKIDtx6+bEp9pdlSn6zG8HHnVaEOKkuaLiee6pHdsObhr
9hiBN1lTmRf05OGjhIgt+hBHJOYDOHc0ZAOSM+uoBy2bhFy7v3f2NuWUQQLONWxc
VkBs4SG6Q0PljhZ0tP33N2tBYobbwqoYXs70+w1XtEZdd1zpzdbsEocccRdTr5+N
MqpA1dC+Rob9+lXaE+ce9cg99xiydxOflW2LJDtE+Ccx2U7ZMF4vJk8lfwxYz51f
PQpaaGSTdba6qvcySzyqrg2CalJXW6t97ZfaPfhfxDBPUx38/N51b3kFx1akmewv
496hfA78K2ryI6BaBe35Tl6mtFXbOWZ8XaLiYVEaQCUhlbdrPdMu/BMI3D8Qa6K3
1X7TSJw/mZpbwYHuyO6SiqADQHfaPBLQB1Jv1m2MDrwOhMBkLwuuNlPK14tfw7s+
8HEEIQZBq6x9iojFZKvVDkK6QG+XyZ49kooF0mA23vYSI1oQmsQG+f8WpCfTLoFG
dJumtBK1jCaX/VXnFC57T2VOyFy3OQpCLqTq/IeJiYAxLH399nyktGFtdnZ16OEl
DjCqgCCvP8tmCZKjShAVENhnm3Tn4lNgTPvNd0VQBSeEyvK1FPFXgRVQVxYRiQlm
0SBjj/1k4bYcGWDbNhzXvuErs4MEftDwDHaZ2k3HNCyhvaVD6+CpXaToSE7qZBV+
3fRcaVsvtlBiz0p807KzNKbNJrlmBplitrmKbNP+/juV8iBlU7KcUHJvyzDgGNwY
zPXpsMlrZG6UwZo6kwQMwYpOkJjnOe/gkJAx39UyRa8IoWI7Q3/VCXbnIV6RVcV1
rOhEAX78/vb3EEGyGHKY03n9SE2BpxHzVS7sMy8JekdisBEIKwSX4NsKtd5sJy8q
mxCBNn1teO+AVWHOwwvrRwnY80Zax8HfScD4HNIx2uLVSdZS6HqSgWK32LDdb/Jm
8Jv9CLAg5e3l7AS4m5rMks+QVSSD1CL5awzucqD4KZQ=
`protect END_PROTECTED
