`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RDmDoywMJ48R0LUEkOL/7h6+lDqtCbruVOaJQBzICjMMrQhvEBw/BmHt2dk2rYiM
juPq4FaaeKyaQsoeSAbw9ubwJL9zgEA2M+xfJ5RdVyw2vRnwusQ78hAANjwas1cH
OUFzz/MTwMfLRy+MNcoagfW95Xf6Q0AVMVQzsUdryJ3cuODPulEPYP4nwh6t+5aD
ici5KhjPrbInwUTZUNHLhgWpsFrea9DVkxXwM2MDENLfs6AjgSDdvrotSPS/OtzL
Zz+FedsH688dFNatk7uf/kPaSYYMb8NEkwkAeSuu6DF4z9VOZ5zaRKuUe8xtQC5d
Se5uSWfYn+wS39ONlbVIJ0UB/7BssQuGUhcsmbYY9XDIEF8ThRgkQZ5FYxeNEHjZ
/RCwhvL/O3ulcdTc4RjpHnW7KOWlnpIKlGvcQnPs2K9SqXsL6hxJSflUt1mhJ+0g
NIk2zyp/NGCg7r5bJP0Sr1If2LNG2E469Toc2bvjmMev1eocmrfBgbkSOesJ8jci
8ieDKGN4mqTHrsw32utg4C8Ac2LpEKL7Ee9l4J5VTUaz90FafhvCmTNP64ZA0j7a
59UOjGMd1Xeb5aSKx7p5cR44AjmO4JXsdk4kvwo86/ofKe9DDq+znAQ/FZaupDrS
BA93YLlNwAAFSeY8aZ/altrcgBmOg1Wuw0VXCXEF4fD4hiQDOxcvL2C/b7+nm3Of
lPWRP9fUCuV4Fcv1q9RaX0mKb0TDdbsPr/5lPJ6k4h8QWcVNcM+CNb1WZqA3nu7P
8EAGSGuctbvzIBn8gtVafJgX6ODxZ8uoGVyi6b42V5KvZCFHLWtF+hIuODDH/Ban
8ln5wsozLNIUQ8SLUxft8KdEwZupbIZ9KEd78/d8BW+G7ogIYhy/Qw4QoNpCw7dl
VRjaarfkqhDcstVe6wl9lSOrOoniR/mYsU5VqCSrGDMwDsOUUxv+GnkW/W5WBFMe
dGGcnnheiha7rLtjti6ZplqXKQPxSidD0V2dV4GPqz2IgkH14fhnMEbnPulXPN5a
B/JF+KZ4muZM2cxWGQK+kFEM3NXUj2s1IBq7EFQeykOroKbi2EtmtX7HEHAPPSr3
VsscV03ZFpEwmrlqNHjFhZqYIgjKXSbUGi5fFzBe/V76eazkGrx3VEWQVdr4XsQ+
aUHgE1pPw6LU+P+97htBU0mfloq3kSza1fK4qB+DXy2o+xDwH0PMCXil8xmg2HLU
wnE44a6mEylQGS4u8ZzVQLPZWk9Flg9YfrpLjXqPUyIBTXUrw6Znty5OmoXRW0+M
EaUk619Hix8TI/96LYaXGrgA8UOPkz6wo/W/Igyxx9l0vPOgqgUTxb5gUGrKZ+Kl
k7wIF3fvuJNQN/8OCodJgOY7u3tlfsxMqX0yPRazwnoap/NhYZD65nds3OyMR76b
oO5ifWEBYjjNzvzglYPx25w2I/tV/il4ug46GU53uFkWR7QwPKf79kWbCKZe9yGx
gSumrm4oKIxBVAx6f7N2+TO35fxw8KSdDRbezugK2izvWFGgi4KS/1tkCP8JVB+k
jzfOZg+v7rjIPzsG4Utx0ms5n7SemTDJL5M7dJfNjocP4qRJYAEA5hp6KWN6IBJK
qAT3zxsZpIW6kctgSFnmwsKAIiNEgSGigaoiwIi+sx7FnyCjnGOXOT4GqNXyyUCk
oN+uXh3R9ppJX5MwTAK1CuCO6x4ATqRf6mqGLByO83rbS+IGEZGOgvfpCHgavlNl
u+RA72YU319c2x4KZf8a+EjJBG+P9JK56di3PwmZOSLvAXwgeBDSqBykb606MQV6
ZCduaBKL0LIKkVfBRFuG3fb2T7psspmnBbzg57kWCanwchfMAysCQfNH2Evftz69
Hgh0HGmXZawJU7cTE6nn5zBAk5blPmT95c3PMKBN9l6DC0TOPnthSyRLiCF9bKQ+
APrPQbDzN41uEEi3kFEIyBYFxiHmhvMbteCXHX2KRZs1nQ0je20+N6WS16PP7zdf
vQupPERumOrsfHLL7YtPzNoeW94249JCgEChBkgdHy7OwPwQAIU5FC0j8vfhuTZS
BvjrHlhq+4ca0FrklekgQQcgBpniBrJX2uhyL7ef2zGUNCsVMqh8zugZCWenywqR
fqrsaMSXSDnQhG6Q2ST7D8JDUV+78P2xILpNZwteLAlxhpgrs83G3jKe8rCCvtpg
p4A5orAwTz9DORHLOJJaZdZdM4/fQLnaJh72r2eKtZ88U1N82vXBpq7pvEwCLe2a
jeKE1mP8nJZOD1tTCeueQQ/8EUFQL/mUENFNBtrutfOCcWJUn0CledVxstHnaRAt
96/HjRsM4XYZILrwcJDRFP5sk15cpw22b1Dp0kbfvpQV23NazHl7Ee/OqUn63osr
CqXWQ7STrhrGFGUVyqehnZ5BMDs3JHQxjvRdmc/hFMeTpqabB27Q7qH3wfU9WHZA
KMJq4l0ZWJ4XmHWLBNHTI/VUL2f14P7IAkaocvOdtuFdRFejv7k0UQ+51LYCE0+8
WZ6RMDdWj4gXrJf7uQKlMO8/wuK/7bM40rtswSqx8VzIL2wVQ61TYAHjgCG9IgRJ
fK86+O8pz8+cEBNcDH+onAWL9n0/rzZoIbX9iosz25i5AECCnyjkMu0gSb3fKSsx
Nkhgcq4ssUPiVzxYD5na4yXxjIaQv9PveNpqoZwyrK2KlPhD2KoRIBYJnBH/FGoI
lW/WxAmN0bB6pTLaho8KKS4x0hCf9EbxUSwEo7ZD5E6LXO1iXiooI5rgS3xrF+dz
ZAbTK5DDR7ZchFtqGVCTQ7k+zg6j1ASiciu6t7xSX7NX5Bwc1rscERg84B5x1q4y
1OARKqxZTA5sLM674Z8bizNuSPAIgFg0dlT6zMYgCxlqgY+4WHTzBf/6QpKIkjFE
zqllIOUordL+6Wcte6b484i96Pw3E96WIvOznTXuJaurQEyokEfRt2DL0m5UImx+
Plg5l8VaKdzIFSr8y+1i87YQ3z3xW5BSVRHV/iJBsPybTKQli4wJctC5Nd1tF0qV
WmYmSXS8HDvS3FSPVei+8A013ikF2zIHU6d/9tupbBsxCMB+WbjNMxLWz+j3zNNT
R+cQwab16GMbQyycqoNT1Q==
`protect END_PROTECTED
