`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cvsGq01H1/oHhVvBILkF9lFESsmOHLDVA3+ZSqvYdh//9PIVP5wc50EbLcBejecu
SDHVsReWntV70sKC2v6HhcZ4mrEzLwXxf0vZX/VcpDXYeWsyByGeKJAVEdnglRkq
nGiW8H4ITpdncee4bmw9o1eckTqVq2noeFjtokvTJ/er8NuAyN/M36smEx1bswtJ
UVqnI2SeVT70wdZOgdHOseL3jsJP42+8irZ18BdAlJ5GSRD+myHEclbRuLZny9sT
VNvqRkBLcA67WmaGJstoSDei0ncyRvUoKfgEKjvkNJMbPcsBydx4iMRQoKz78Qoq
yK0T3/KZ3m51b7jaIiyZsylPXVnytQh6j+l0ynWBVgs5FdWgtgsN30bLuA9AkhoI
+iK+Gh/TNr3WgclFG2Nb5PXFNf3e0ypIlFJTsEE0FkL0ptyRCJUVbYM0ahinZSjJ
Q5B/xiw85Rn88Pe40t+rbzq+oZ9KoZovoU8WwwqkDObYm6OQZ7LPjBzu3/1TtORD
YLGzAbP+e0Gwa8bByimwxUHXrUbr+qrOU3P4WypvQJkP75oANaRHzVpOdu8flo2C
TCajiEn6vKcclQ9Uno+13YMS54LQnG9KuUUC2f9xnA8XPSOiTalBeEtOFWdKYf9u
OOEpWEcNY3e3vvpSdKH3/EsuTvm3rPyzEFrdSMWUfsINFIync92DLreey3VV/y0u
DTBywSNm8B96BhX04+mK7dM1pLAwVEbhseLV7aSZrJlCs7WLXW55Jq6o5GyZot0j
0pOFy7M6XAVNY55ddQAB3Qr/VESpb0qry+C4p9mYnPZ54tp5J7QQsh0EEXzoRolQ
WBIVXNmj5Rx37cWshywQL6k/JappJvJQM31NaP0gcyHeFTyHBGT4H2L4S2x3TdP9
E78QoNl7BYBwjDL+WNDUDoU7B+p4SRYNOC7hwuClbrCi6EvZdCdt6RoNRbarp2c6
1nEFKbjdxybLc06CUDkN/adW7MTg4NnPR6YSAXe7ya5xwuN4YcyLHRhMlEeUHAQT
EDNDawcGbE7x5CUynPzdMygx9T3pTiFQqJtdV3iVNpuKj170rfkKZhitg2pX1J4s
cfSSWQgNnj9DqyLLTKrJiwBf5VvDEup8RMaVN4lP22oHBANK04ALHuH9cY3vLtO1
ybYFzcseGktUEV8gZqPzmqnynvnQ0t6V3n5bSMOmdMP2K1RXTZ6n6/+0vsSEmn4W
Z4Az3uALIuxK+/YVsSyMA8/85hWc7teKJG8LpeGZTyyMARDACSrbzhw/A3lWv0Y+
ZFibdwqQOEY4QheT+2W+7i2q4T6P/O/3CgS1zKbMDp38GUQBe/jOrvOQRfL/Ztqg
oBxQZ+KoLKOx4TjYuPXmvlqfFZ4NFjzSo3stKVIN4eE+JYIgLsaMS7UNsNzvQVSE
8LEpDZPoSbd7e06r3f7exhbHlw9PTGB34R20vohgKoEd/1zN315QRjafQoTYJFR1
I7RvzPbY9y0pHeW9gAIjgwKjmgkMYQNuQ2QfMWmZ1Y7L8E25ZeeqlkhS4PmPe573
sgjPpc7fqNKWgzDcK+hYw8Ulpp3xqLOOGcxV+Oa271S0xFvDP4nnQxbqh28EeqaR
o0MVQzDUkvjk4ypMjmcpGbUhSsStwz9n6wh8p10poBGIqFwVQIbvCgJJOY2X8YA0
1aMBaqQYjwZPc1oOyvacgRtCFfBkpCrm2cugcA60PWEiGht4BvXdlVmLnikPHVph
ebN2IjfE0JHAqHv9Xk66GYkadQ7+VEa45SNdxHKnQe4sPRaspQ0qrNOGTLzhCUma
dCYmvnZ/iNVka52EnkfgK/4pqWiboQlcdGOPPCw2a5t6Hjvv7d+Em0nfoX5es/Hm
6aw1+oeYfKllGFGXEFLpzV9KhtN7pkmHtyS7+RT0snD5lXU5b+JpKq7Mfy5rFYkf
MPnXabR7sZao+we1XYduHc9fyGxLZZezNOqIPr9q7zkYxTLod6JCIV1M5n9QyY1c
5kzjdVn/jii2VLa2gJSv3CrT+FYKuq9hb+GSMPmiPrM7FYiiDbt54Y4+Vylev44n
MPUlLcJTkECXfZaOIfw5zaUnLE83pxULe3LWpIekpW+VioXmuzsrvAzPLgB8jvsj
AYySfIfGP1toa0FDfP3eJ+KVw3/6wj+NH9nXqg359GulBUFd7gkDft15pgBcs/Cb
Qx7kfr2yUpuXPdRcByXvvNvjn0L6K+LcwLoG2gqs59A4lsOPc1KDHasMu3lx1wAP
NzFKmUBb+o6e3/43tUqCslUIc/NO1Cof75o9305oNTxAHwNEj3RdzPpajQc4lkJ9
m1dfS1eSsIYx8xkK6R7TBXQl4f4MzHedIiHujrJ2UWqtG/pUzolWVIGhlpc5znJf
Gv/z+7NhFo7n6bFMmko+QVG8847tCxnfCU578WcPH741bBH996c5W0num5Sbl5Fx
3BjHAQ5fppidQl7kO8wiWa512kHUugPlXhPmJnq22QEG85cdlS5fB2q8Hfdq+2ZP
dLiAzlay8RQoZRzPPyUp7doydkCw0GumAR5TqbeZCHyXbv44IfZ1E0FYPMhov2qS
iMAEB5T4jmoWIGChfugp+8k8WPpjqbhrPRyiCK3fxInFR/kaB+tQUvR+c7XVZUDC
ewE1skmxFYTsvC/h1YXzMvDdBlmNZfpXmy0AcfR7YBOxQsOyUf43vo3EbhYnOdUH
F0YX880RXCoh1arh4T2LNx5ph/XwST7INyCvgk5YTM76yUIJ6wuhhrY7+8VhEPzM
3CCdRm+02cwXJfBCypYVNpqfo7UiQN/fAXw9ogKOsLC6NblahXYjc2+BIG1rK5VJ
fZDewfYF5Yg6OC6VG6Ra45PvcTRxoZBD7mWehC7Y2mW7L+qZPOnr00ZuMuS+X05V
2xfjW7nkc106zFCcNcVw5w21zkXvkFQBr7KN/CR+1hTHGyLYQTrhNIDZBfB8IW6U
1lUnglTQrK3iDeTpoVOfQjjKw/9SaFEiBN8VuwChERMlLOQ+75TvjUO3u9EhsvI5
g4P89JtRyfGXcHMCqhcmCTzGxVN5aBmmNNfp0nmLgc1XPsIOI+0BjabatMvuheIb
RacyMJf+07q/NJaHn4XwSZrjlEDlbS+5JGhF2uHKbyNEF6t6WDr80DN6GflA7FJ/
/HbaS1i3F9gZ10xnVtjNA54i9jy4grqbkLy9V+JSbE4Rd8NSmKEbHUjIzHiqihII
RvsmNqtAyo/LCOaI1aUHi4sktLzqLeUfxBRsIjlWtlcD6b4fWW29gORuODhstRs/
yArtYdB/pXWhX9fnvW7Yesi56LqfTBS2dJJ9DkTl93evNuZgObykXHDMxh2KV9pV
DoT1q4XPjS7lNhOY0uurDLhCLdmeZWDIhoVchNIOw5BMONl453ukpribHVdu5TxP
Qq1jemoEm+bS10rZ/4P7emIfM42ePVclK+S5iZsr23DiO2dS0CNcVGN0SjxFDxHz
Rep1CiQWH3ryBVUoPs1fFUH/n8QKWwqfNUjwRnLM4WJh3q1K5AC7GuGRLGEAzFBm
ExIawtkfOyFxLzkZ5wbSbH7DpXlv+ckESZfVtBRjiqtbFxxn9dHgTlkzHAdYOpAy
VZigfWe71ADf50VLTbKR4vNAixkbvGBc9RRU9zAyGq0ZwuFVqHjXGTSei1VQS/Nr
Lrr46q3qI6WwAM4yg+f/w+rSCw5tzX+IUPvFTbOrBU0lpTVPR5+aVgd2FLXXTmPQ
3WZKw4/SzMl00MvhyCt/iXkhm12sxdhQdzS6n9rrMiK1DomL+XCjfbyuB6uXCi6F
wMe7C4bzD2cV8L09KS6qa+ui8NBPsQtMD+jfH9A4EGnEhFmRnB8CFp9E+6G4P7fN
AjQwelT6IM1+pc/VnwTWhs13go4fEFR3LdOwTj14UjJq7nXNnzVCr+w4wFrT7z6S
z0Y1kOgbU2rUB8cRpDsaWe5RVmRI4NT7lyeSHJg46pQt9GWRG/fOwUBzvUpZdi62
6a9W+aet1pk9dXJN3ECSfaBmr9igT8T0JeI+6qf78ePDfqQdIfkXD65ntVHavyHe
FlykUP4LfML4ttIQ1Pq3TS7Ks1Dkm//7RoRQ79jLJBm3vNHnhUCUZAbQ95a7TQAh
OwnX7GXPwgZsED5ALBjEHJCWn4S1z/8P0QODGklCQ5LL6mv2VTpDBY6c4sL6XrIF
uNYj6uC1zpreKkKRWD8S2GB+BBJiEMNnuevj6klFiN0OD1MjVu5gJ192O4lT2PiJ
HfKvmR9ByLBte2LQ/zVWlMCQaF82I5ZHY9mSXQ9YOxO9R+XUD7TeeYcIPRKpLwJL
coHzioyqdonw/zlDOINUSLMfzVLzwfSb22KpLft8sSxp+9uWoeIWDaXmrz3ggtke
a4YlfB8efjELcgfv61zImFV2iTbIguf5GAyz+ZxAdUadcwgB0uag4RfSV0at4qqb
mkgP0O6IPNbPKwcOpl7YFvl02sESaegJ1PME9y8SO+wLvl7ZHk1Jw14GImcdq8+9
faTa2L1zIEj6PvQzyWjmSYl2yXIzFiGAPA0lLlzAJpJ+s/aIill47gkZ3tVfBe1n
pFX5bgi89WYPAmm1iBoTwdSkaD2VVtsMbF4uqpkoi5UX+ldnM3/LMQB2EtOuQ+Fw
E94gglL/TL2ALtZTi1CGVUaEjho5orheyPNdjUIMS2xtmWHcWS/8ESNYO+S6pclO
oy7a6FN6LazMDzWzi7VH+2bwJ9DmjylSgbs/S1JdB99RvQRpME4/Q0YPu7PNr7n3
5viOdb4NCBUMzAHwAAq7Hg7b/qG3ntHARGuCeoLakZSzwvJi2UcgfyJmUeciQGjn
ekHyml+yL9/nlVqRZhuPm9aPsRJ+kEWDSPeatLYgqFy2omIH/x1YesfUez0yFiqN
j4lhnBWtXfBoZMplmWqtcNxcZ2Lv00XZIaggs5r0JdjJ7tyD1LlsceDG3gbc35uy
ZLRjyqCqUDmgvgqxVfmAYr2NAcoD3rFl/+4X6lNHUMpHONATVK8Of0LIJHrzxFfd
3JH6SRoVC78bqHpuxRCKtFAAaH3D/c9dVLbutXlvp+9sUG3n2XlxUG7fO/LtF+r/
OPn2VtswFNYOgcvO3e3LPpQLtGzOic9h8QOeZ/iExSf1Gchq5FsrOpw9ZWw7xBEd
RupAr3qvAob4u2ex0Oh8nFHiRW0qeNU0+0sxdJl4hxMYXo9gGKNOdrPb45BbJogA
2MPxqrFHAkqK2h8TOadbxeo2uE4dNBvB41YoQ1NVR62lnkF7U25CdJMcfltn9oIK
t4WzCAfKkC1FQ8wYRGa4GaFNjcCFP2ccUpMb6hdT8eJwtfvl9QciRogPj/1dKFa2
H83oumCdws5t773F+ZTe+jjxlXJQCZzuNTExgGzThGAGD35hOZFPIlVKQDxAc6ci
rANddJniaWnzya+W7W8TFWpQQ1B/yDhABHWy2ealScswG5556Xs8dakX4SU19RNG
wEtKoHIyK+oJ9BUMsxwYLZme1Tt3awtphVe6jsGXYlF4q1zfa/HD4Dg6GpDy9hhO
g1Hv7QfhrdFNp11/jebepU9Ls/YI21QJiaUQeqUYNw4iglirUsgs4coeL8zqBnQg
00jJiJnJRmBRegkFVjeKP7WxU4jJBRxQiGcyzubOm/uN/0MuugvolLmtGfL1xYTX
TLme4tJcT0S09HKErv05K2/9pWHF/p2R4G8i72MerALRglm6P+o7Pf9cKh9Xpyoj
jZ5SqC8DcsmrqGVMdfX1Z1FBO84Y2eswKPsVZkT4/S7XbCp3o87sAWCb06pO9it5
F9wKygLq+o3uLfo+1eUDQ0PXtikLJJ5DiGXY577rEOMCpjXSUJ7JGHoQjoLtbWJn
KbYMTPybQ4yhshH5LBgXvroT+0lk+CKLBv33SSTLO08KiIaJkBEIlk9wVZip9BgJ
bldryMcvq0EseBlZkAQb547U+NnTCZC28K4CT3c5+7lS7IGKzm//HKD2McHWttHc
XkNFcwLi5B62iCAaNKX0qc/KcXXVUL7XJzXVe7NGlp1Vdlk1qOzrR2I4UAeqQIiG
HoXv1h10zf89yl3FWb+VScwq3dAVTESQBnRtN+q9LWJc68j9MzEkbUHzTRAl6aiz
jvzGJG5nefIWOHhhtuBCQtEZFdVULV8JTyEHJEuQTY7KB+2TtAr9+QnWITzCFthm
Rrtjk3LTGgUzqEi0iphnPf53c9UJaZWPOoGZVGwM7DCh69dExxz8TNyd74hCdl6y
eE7IMzG+Wvha7fvIMETC4EExJlt7FFnaC+TpJuZEqfrnCfURC0wPm/Q6pFcD8bsP
1YGYrtdmWcq3rqOyfedfhDrJAarQfUSY8q1YFAaYUxcLt/V2UV9jeImvNm4AOIR4
fHysC+wD0Ucv25beF6RoeBWev0ftp1uqFaVgzYCewSYVtASsW+kS4/iAya40651z
B2NRbxJYTxkDEpHsGE85Ltw3Ah5mXEyuPetSD0mDWcq4qtfW2+vBuO/X4mNE95JE
fIfbeuvp5wz5Jz+MhZm380r36QFq3INdY0wpvwPzBCqZioQU5omBDyQTWCinmnpD
DkcqikfHX20+LV7EDWMgT4P5DIz9px7TrP/yYAlNxxEMlEjGoROMnUOhOiMAZJ0i
Q4OZEZLbi8Rxn9owGUlKeRErpNYe4ttnEA+BUyyC1N+zJOyugRXoTUrYyjOZYjPL
eR0xLGNKc0uJ/DGQJrJ7KNWPxaYVDnpKiieayIeRG9pMewcq9Icc/Xx5q7m9LcvF
QPd1VW4v9ZqM+htw0hSPoXktTDT2VDt/b2rjs6nq7vh7r23/jAIJqiGKEl1h0MpO
q9tX3ZCjikih8lYC7w3LKFWLFqqcQ5tV/frnjzBncwGwA8JEqE3a5HeBrXZ3l5pp
Wzx9up6y6TL0JElMAKDGMCiBG9R8hX2Cqr6nX8SIMImZcWzr/4gB5fBdVL/5ZKzr
o0rnRWkG3dapruhhGBE17u9Avbx3rhQSUNrxo6sOP90nibz/7E3Ov90G1095j3ji
ElNr8pDL/4phirFLk0ETX2FlEJQ9Hdl5yxxEL0AudlVsEuxvV7dZQeNqu/+3N9SZ
KJ6jwhD+OOAQ+einvZl9kiOo8Nqg46ZmdAEEXDUjNkejVhGc8lNdtALgEawbhC59
+h0hYMughyfKAmlAexHGJazIJ8btRcC9Y6gXG857oFZqCRa1r8y8DAhkp2WrDfF8
nR6wXoVd+R+6axlBKCDhoQXHjbeihIhqtuTsKNKjFSejAjHpoqahMR85vA73jHmW
JCsKG/tK3fD0cOaJ0S6BMFGT9uqek3y+fSScKjsL/OJgLHl5ZJfO4uL0hQN1fojv
Lw018GVXnGdRceziBQtVU5Z93u2XtHek1JykNW/8v+hzOWxvSBeJ8Eozj6UT75jy
TleDntIzN98eZFJb7WrEXBLfVvLDldawSMkI/FgmyrX+mUrKynPTBhiOdvyB0PHX
FaXvrr5pMGy2KebsoMbdL5kDwQ0tn8yJa1Mbgqu/K3XLgOq4yDhiVwiAzA4255RC
tN1vPTW8oNosPtbKgTLUunMJcNuzrq+ua2iwL8x4TzdqeP6UIowxDvSySSGA1Ta9
p5WE+Gsb9p8eGoAJwZrJqNk3uYCdUFd5FA62xlK4dn2b+80q0rtlbRaBTGHokmtb
WlFh5dfn4imdM0Ql6ouFlRyRDI8z+9h+tyePK8iTbvEQ7LAMjzMnB9EuF8/c8Fsy
xdrpVMhhLZWgrq2EccWxmftJVG6hVgwHD3V2mxcykFkmxX7jQ76E/8looiuSqeyh
y+80o0RE5MTBrfYQc5nHYTQh7UFYocMMWqxKEcsd4w6PLHClYFXnrLeD+/kJrv98
uzYmHKUEXJOwdSPgGsVnvjvCXtWM9z0txWVPT3g5QtFWMMku8zUhwqYnwfXl5AuB
Ks8ohpV2/6U+J4//wnWWRnVraxx1RzUZHafFdaS5C1VFlFkIz/qiRBR+9Hk/8Ogi
dhECGZx39wKD1ts+cfh7JOR5Y43SZ3nxjIIdjptrj2iBE+u6NsyGGXhOZhkvRISp
RAaazLglXa4SnTN5Jk5AX/3gUgYscoj/eAayKElqXhXLVj1GXOh0GAOymuIbfep2
Xt9BrktBGRjr9lzfIiqa2EqG1AEPL38teEmZnbsVuhAHUyifAtWAnhErDuQOWhLn
RBKoTRtrMaVusj0MFdMDCxRxjxIKeUPlbZncO19raap6SDCVv437K1KQYgFIUl4n
jdIFhGzw28MMq+h7HoHKZUUdtTZo/miMx9RtrkjEEAToyc6lpnUtv+EN1aqtKu42
9MUiHIqO/cuTNbpfdM22g8//71yZHhh1t4OWAiO3dOj2seS6lgkXIdLhNcs2COQu
TTG26P8kwBDqO825OMER2PVgw0gzIWVnjMouNNRrCfKEwkz1Q0MPQ784H6N/e12D
I5gjBsSWYuYqAEtqSnc2nMzdU1KwemfeJZoPsqrnRI+9SyeG/Vm+fFBfr7QCSpK5
PAIb4ujTCBvMs1lQqZbqVoF/LmuAq7PIblEPUdh9Hop/Jc6jtRWL4AOf4XvHLQKL
9bdLvSsgFMMTmEkXtJAZErfKtW1Z/g2xwDPz7pgp5721QVUcDQ1Rrw3vWsmCZQLA
kfqoAG1JROScdt+ODPtZNVzavivdX0TJHxRY9IL1PQoY43OajNSIvMjx3BZ7sC4V
zrcf8cOJDN8woIxcIqvWdYemfWbIoiDJMThFWPj/i/kplD7B8dU8SNBE3cAqddqO
dhsosfB2u3NeSgD2RG2Lxg//oJUs4/OISnEfTChYKops4Vnf05QZFt2axmP4wFDA
jY6uBhKvB7wwWDPXuq63our8aeg5uGESAMyYLln9LgXhxQDDevNC3dRSjSJtCqMX
6LFgDW8uxqrnjuHaqZxsEctdkvXVDfZh4zgPtoEgjVZ3hM+UbU5taknZtBEemUeP
8hwL3nONgBBeldRVePxc+3fg6a7buPX/hwoDWKomhAvKF+lTz22wKZc6JAiGt+Gv
TQcHL9x9eznlsivVEp+rRxxMPplBmoxoS63KC4LJM0vAtVdMRRydFDdNJehPyixP
2T/cR9vs5AOrIs3PojZqEclCNfg1BH9UByrkMSJViVvfqsNi4KvcItiTvyQTw9jL
Sq8Fc9O+7yXZWKE3L5ojO4gsf3fRn1+gq24qfSNz18c+orH2Xk1bVCQ0d+3tYhoR
BkALw7nCFMxtQZIv13xdY3uXlwbUUWGBmlJv4zw+yYXkSg9p8wypvXas253Sl309
40ujNS1I7aP5VG2c2p08wWHH5lhdZkLW32Om+PrrtqXKBScsZk/vvWvpOxU/375t
QPvSZtMcZQoJgnGQk+MSTV3VhaAfcW/HvS6Lr80d6zMxLwTFibnJlhNLH46d488F
KJEGzDi725GqIoouWQeh1c70fc3M+VsayTBD5IBtgsojbXigmmuD6ZRLMC/f6W3X
s5neKVM/zDOFXRUZNpbWnktloxvaLJnT0TYLV31rRYx8kcWFG/3lWwu6CTzpYTAC
ikxQtvlXb65Isem04CE+8p2/2qZVLRW/+LXXqREjeD7t3m9KsVWzbBuLpDA/ROYH
ncQxd+fhVA8qAr3dgHll3sc45P24GK4l1aqNuaBN8rqQasr7n4mATchjagUkqAZB
h1rwBNX2GB49fmnenlzWF/EjYlI+gtuTsyoX+WDnlg2hogp3VFVsBWz8PnsH/JFZ
/+9GTfF8KE9HMT6A8kfK7y9J+0NWOEzX1BmBYCm5YCoo+dS5lUkFDnUXPbYw7by/
MuiGfg65mca0FFDJeT9Ap7NFWTBFlXtpqeK/qjQxD8F55AOjT0A8IfERPuQnf+B2
H9a8VTtUr6ju9Ph2XK6fAEOw5C+gf+Z87RmbIpLCTKH4Mo6aZrzaFSnR/iZE21Uq
Ip8YSMHl7xwn4QSiAdze93wpfU819VEmVrLghLfjl4KyS1r2vLzNU9RU15M9Ojrx
kmORFOFxhmMH1VoRHUgBuznBws7M9/ZIuWeNaNUZ98Rvtb/gcFqURudkYxzqULPU
Y/+x+FQm4V0rYqrCGBRQafGFEmpxRDZBIxBGtc6X2gvrTZ9fcYT33WJge57ywRec
B9VBR/IRTUmRQxSaEzJ+CM01NbumP3NJoGr9hZ6t8WtjUawgjbY7mYV2MfGDDO4z
k/g2dEfs8F6lZjCl8JS+/eLV9BdsrW6f2rvETXPjOv3S07o0d0gxfa9kw3BxldAP
eTu0GfNAAxHzpQOcYsmPvunCZ1pjD3mxneIfXkNT3AT/iyGA4ujeQQ4epqmNEn9n
v7q2rxTVo6mfbKFyX4N2qrvJDsjbxjwpzo4ubzrUFhfJ+sXXGxLYmroUUBRpRL0r
lUW8HFOvUEt8lkw9BL75voc25BmH0374aVtJd2T1Spcr/YxvQEjUlwvrJ4alNEU/
OJJs8qGVqi3T6Bmz3HmejAEiLjyU8LUBv9KCLjIQN69J4XcRPGi7iBzuP5RYr/Ab
kxVdWjJQ4beC17/ErNVfSPhitesWoiXW3YYhGXZKALR8BxWAgMlDl1t4o9o4h6Im
cim/n6/VCELoSzBb024tXn93zp3CpiyBs/GpxSr+iUKcbUM+ELcaeBRA+OuMQmR0
nRYZp6Q4VDwX3WClmnwCvYyfyzzrfmuLbhWbcL89IvJ0fAYEXUn0CKIRmCBSo88B
a/GqSQfY1uR1w/EpFSbPt5KmBKYKR3Lnl9YZGhFyVN8jj7gaN6nrMiBT5UucB7m+
SWKLjrkWxjPynTzU6WehzneE3rMx8VdZfr6XX/7L4eDGu6eQu/AURlEbU+12lpY3
QPyRQGATilmuivP6TlR5wphrRS8BhNMXjp8jK8rSGaWpoq/3M9MmHTOCucjZITq7
I7hm/7yLVSlh8lzdGieVFXEKxI11FhAfe+NI/bp8MKSpvsSPzS2tmqX61ahcUHoM
Z3PqDwsjWfeBLdbxmOszJA==
`protect END_PROTECTED
