`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gV8tp+poKapHGdBqRsHic8LzGcaf7culhzTqRAU0/TGJkr+FigvC0N1H5M/ST+vX
9cYD0nLfgPaRkF4i5D6gpXX84u3r4ErKfeNFSC5EI0+vdC/zCy42My4u/bDL3Xn+
Ah7rZP1bCqB1hTTO66YZRBMfhutojvODnjH3TQMpgK5P3DF/BUxEu5iS9rUFlT58
Km3Xdag9+/Uq8PHFCaA1kW2StcY+iNBhCvFJpXlsqbVTmSiK96fd4Zv0ypZ3kDGy
xM9sE1NSkhjhbW60tQraxDiz/KOcGzvpTkiUnVkYWCBqLg87Q4zhiap9N0GB/Pr8
t1PFKpTGuE9U3eW9uv/noeR6MviolkcQGcMm5lY3nKqw0YPAXyQtym3BxvOsk8oG
+AWOBWgq7xGlsgIjFnjf9r9v2J6phO2JSteOmWSE/Pfoc3nAscmfQPBkrFgS6EkL
d0fj5OGSxev7iqbN038jIenR/M1Qj8a4wgFzk5J19H43ETfIPrF05yiIxDK+Fm3E
Jdt39REsd1tdYOQ7RDiyJely7Mqb8SoHyZcSsb/8TEe1aHLvcvetn5dw2SHsjZWd
TYElUaXKls6vaArak0Yop/s4oOj0LbOKOKpfZOo8esxpX0MWaS50X4H0GmGWioN9
cbQSFXMaRCyZSAuSPx+E+AiwdpUW5jT/3l3CwXR1BhKuuSLBS/qs/a0owfM3FvjE
wqfxzztWwim9RgrSBezgBg4e7yazZewDXSnyfEnHwB1St2UwK35fbiOWTQ0dbkTw
dtqGLiwU5w6S3+HOVKlnYBpoumMJr4JVmBg3L75DZeHxg6KkFKxjRRS6gjjjolH6
S8JaPggJz6eewhoEOtRq4YOhQVSFeFVvXON2xyu03D1zObkGQFe30VLheM2H/1iO
Mal6M6gmXp846jwCks4sylvvRVvrM4d2yJNHr0EXZVQJJCv/MG+oF8k78rmQHWoH
SngcaYzS14GmTmTR8pXqnkTBo7VoBzyIxQmFY2aglY6K/X7NldwBDE4m5comqQ5U
F+etds1vfMlZx3nSKmfmgqu5lCWxuNlxK10q9tlX5XwbfYuJFNdTde2+OA6F+AFD
UHM97I3Qck+odN169odZDWbEbgzWG/n7W0fWS49Njxi9zg7z2UsZT4mAolWjlEpR
q+JiekDilV8FK+H/WJXDtX18KkrNCJmSoSxnOiqEClPRuN/hd1IH5fwhuZjH+RYV
gyFbmFS55uMUuhsA6fylILn48C7KrN54jK+SJsfbs6cHO1xG7hQNPotonfeflaaM
2Pg0BubBvL3zq3kuCsLwiAUfT9p9Lazqqn1+4/sNOzP+hK6AqSC1Ax63C9eMqxBF
Nv5BiXvMW2q4iIc5IgwlqZMRfhc6dtbgJMzMR4qq+EELtgonUAaJefVtIxUugHFj
LEMbbxNj4uEQ0Gh7/z0vpGyXKzlgWJcZhWkIMkhuN5sw3iFUxRvaAFLA1AzrNAR7
1wPLtayi5NrhD4sMkEVKXNoQot9nSQl4kxfnFd9e1O5uvDh75jKv4VUn4U+phV0G
QoWbL0z1g0/ohg1+F/iMF+71CJRQrmbpd0KkDM6oRwI/fIIpNqQapWRH0v8h1ykH
sD/VuuZilF5cz+J4+sApnQYK/HgNbo6QAA7BpEu8et7Kq3SeIZQMYRJHtDc++elc
z/+TQPkKGSe9IbVBHV1rL7ALKATYr/EGp+wrS+QqXCAzgUYYIuaAyolvA2cncZUw
wlWr+qLg5y+BM/cbGFTIEK97jtsFR6NGqHIhJ+U22S5KuCL2n7gj+fY2c4+PUVTm
xMo0XxNhEU1OkEB1cbPgY3X6i4d7Ze8iZ0TH2byZJMlEaEkcxaNggS4i6XSd5o5T
Ak9mRZCebRpa6flHt0Z049sNN71iS51WsWv1OWPIslozbdjD9N/aHr0OHGcYrZVm
iqC3kHE1HZHycq2MepC/o7NuR1DKtFdDNCkFLDaqELw=
`protect END_PROTECTED
