`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QucMTmzgYNAUJXZ7A32meBf8j3qpzs4hpuvbm5H4K19J1cygBk8VG68IUN7Mswyk
FNurZOoTmBD9R81JYKognnrIg16nt1nmMvJhfD7yrtu/PRThfjmV1sSWwKpoKpcZ
Wr1FU28GBorxwGskXffP8CFcSESFyChTQixUYBw22XzaX7ig3ScbutUQ/N4aBqiv
WZlZTQsLJr6pBG9RZhScqaHB8kd4B8URVoQJE72R70uEfuNsZ2rSVv7QRpLvK5vX
Ht/kPVA6vk5a3XFMOGHpUnE0ZuAzrpryzTAXsB1qwCbD/UhNE/xt+sleJ47lq2oj
0zFV/3waa0U5qmiHZF9YMpSUMrGUGGVWv0kUa4fNuP9+Cw8kSDeImKKOWmb6Pkl6
Ja6QnUNiTcLrNk6FilL1DR+blrsXEveXtLeagwhuXaZLqpnsqUFYx7DsA5YD8Hdq
k6X2VgczdCiomhL8r+2sj5QjHMrKZdWPgY6S8Fd3kkapbU+AWcHdEsW28vbwYOrG
fYRMOI2fpnk2ed3R6/Bf8mmmFduw6F0GSdGRSUGF70qvnaibJ8NYsvqzzE6iVWfB
39lwbBdEPuJFTVO0rDH72KlJnb7SvQYNXRx+SHr2n0qyqybH9+mCj0VjDWli5JN3
fN0fbqg0cD9Cf6d7c7khqCEPSq/0xgu+wRJXhpY2/ag=
`protect END_PROTECTED
