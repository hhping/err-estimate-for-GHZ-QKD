`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tIR3LFk/ThZ+WYP3G0kX4m1JObuUrM0sSl/SVyxPKF5ngOz2LPjh5/aXEA1ai/bG
HUteyKVe6gD+iH7b2rQWcMzJUzu1p20e9pKFxeRiFMDnUox4a5Uaj7gE7IBXnzBm
FAQoi2UHu7Rspr2W0hmvw7ygxA89pmHJZtv+R+FArRKl1wTMcOI2eunj892r286U
PZnfS+RkJUMNIcIBFVlzacGm0qoWxviTQipVkiJFDmyaRjwTfKr2v4ljjlVAoYut
kIyCYn9y8B24w71aY78RXckDGAe6aBPPv7waZsUedoEoyALEWRLMVeRYzejzFqgx
8llCI8m+9FvwL5Wpcx6sFHzxS+xpjlnMYMiswdOPTQ74ZWbfS5i8mz1vVHbmZ8/t
L8YHMcgmzG45CmswJ8K0LAwD41iDp7z7+REVklVPlHO8zRE8fHRbc8QKu15Zt90o
XH68zAOY2HTBi5Bd2z5/hLJFgAeEhAj9SkvL7Mi75EGhshddPn8vKx48OKB22mMz
iTUFUIYcjv2FegWW922PNRnqtJfTOk3X4ejoSckRQz50YzhY/liR9XEcI+rHZsb1
42e63iyyBt92QKSeQiqTUNuGev2M7LLGjVT5cfSNgXndQlpaDND/KhjsQO0E4m7f
YyM9iWUyZFdsLmVvXB4rkEfKs0subADVan65HlibqTlZbcgNoJ0XzFpUnwRj45ke
EGiRJAceiN2vTwy7jXZNw5FJ/Pfk9OyD2WCTqaVy35IrZbbe8NWEMpi7WAxVu5Tc
`protect END_PROTECTED
