`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eO5TPd9LPgBxQVAkBkckb6zKhfbEWWe0K/+x2kAriuJAoiebFm82ZejNvXWYpYjy
CqNTRSyMUqQTS8BDgTKRKoVV7bedfhauFQZ9oO9ku+qpw93LhxBig5d2ibdu+LeB
nPpE/k5Y8sF953xaf631IsF3255R9gsg+h26nR7kDkQu6D6IVigT/SYp68wPb3+Y
Yxes1BognB85/Qyc3xaX3HUeYR8F/Vp4f4EBzk4jz8HsD2xdeGV3eht5ZSJ/gevq
RICotzO9UvgjXMvbhsnab/hK+1SnwqMxKU5rPhAmXqDswHyX6ByXL3YDszbk5ZeZ
cp4coqv/jiCaEtDr75oYHL1hFRAeKJKlAkXpnkDZvhRavsK65JXsAj7LEVJ7PWnf
zZDvYPgNgGttZ+nUrl+Bzhgwo01xRPnWClQEcTeHRCeFO2xudz0KJlmZvy487kvw
mOrIYy1kNnyxiziAtV7tK1aHqvDMfVaHE7c4sqvgEF0=
`protect END_PROTECTED
