`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e05Ko+a7KTkpDIXNKFPHfhYeC64CyGsccbsMoOVsdWmxivEFsf29ZXZ8ylv9EISi
4EBhkvxrDs5+GOicZS/zlezYRewqxT+DHn3Vl9tqYueaKgSSiytmjxqKOdOnoA8X
U5yQdXaBGNFbc2R/fs1H0bdzZTEXhylcmgZsa/G0jDs2HcLHBF/I3ciTBmP6Lybh
GWbuoiwtXdr+mTxAePSFkdttqa6pGWNm/5t6RxrPlsCGMFRFUxX7JlK9PVNMoaiy
u2Ize6aDxpVUxopQ52NA/roa2aBsOWKas7OBOKSaXFI5/gmx/hVCNcIy3T56zxHj
nQftmHxEbEoXBT6Vnqw+nl4n53f7U+40E+zFIM3Rx1og/2JivtBVLnrLlqF5bAhv
m61J0lPDhShe8QJkp9ODxXBcrNiXNyLF/wgcFoAAHsW+n+KC6+NjOB9caLOC1IlM
IGKWCA1H13IkcETUmIyhLemcp8WePuR9NPghZmTmMRyvzHRC8Rwx842SA8dcJ3cE
Qd+KzI0jY3GSHV9tsHitBPUEtqW47bk4EuzVgFt7pOat2IXiIf0pprjwUjQ0uf8l
B2gzcw4wvVoTa2vbC/cAobahd2qTGdXva6uRxnYw2gHro4UTrYAfjnAd9fhrzEuh
8HSTym23KJ+f2ZiusWdQgMniBUZ7hszK71Ovs2xxFzUJnD39yB7Mkeyec7z7C/zu
P6BeHdpq1dMvub1+TUvr466qmYzSSQrwoo9a9AfB4CNlmwuq65VEVwbY08SWPK1Z
SBJ5RJAxt359HCnhE5nakRMoZxXZRWHgTnycLGpPqvprgD93MoEFOqU9wo7Dl2vK
s5upoLeO5dARMnsiDZdhqg==
`protect END_PROTECTED
