`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zl2jcXGE0lbHju8NM+6ZcapoIdoF4+NeFtIDo9SSzN4RNh4YvMoTzWHS0f5WlRgs
YYZ1GgWggW0dDVscfgZUyrbFFAbJADMCkydPSzBikyd6SQdT0GdEnZ9NfdI2JOtk
cHxiwz2MVVMYczy35Pu1rVNWsaWIOrk/ftATP81lQRUxORXzjpaHgPns262ZsCrB
+yAB9EJA2MKae/994D+PDtfRLZoUeQUsBA0TkzwsoCkqa8xL7B9LRN9Rx3OryUd5
wAbXPeYEbJelZ6XTuxfi95sIKnRwBszX3NEHajLiCTAPmnSscFmrtqhU+o4lA0XA
qBJSWEpp9qR2pGKOWSksi63su8994IoClJFuwPI2wbU27+wR4AXb9Z+e8po9lCmR
Lcm0wPUwBoIejto8/QO/GgZpNKQZ4i6L7/PpKiFmQe7VlboA4xfPAkpz+YP18dJ3
M1unfUVAx1lwk3QO76cMSpjHADJg6WXIuIvjiSGJTUoVjkgIYP70oA0yASOx52vi
HMl0eneGCKWdyevqsICuq1xNA1/TUnZgmy0hgF/zLpHoJkmLLV/j2F87JFOz7NP9
Fe6R45VNZkAInAwEVOYM7Q==
`protect END_PROTECTED
