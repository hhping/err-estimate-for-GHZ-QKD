`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
99zLTZ1X995cY7izqe+QbRqbfqu1Lt8v7vYh3mCqPfCS/+V8N+713BAChzurIChT
D53/2XjM6mSU7RtNId6VNB3UL9ASJ0OfMWVAefuHpOfsSa6l6OjpbAhJBi+OdOU+
fLE7GTn1W8x27QiLG0EdpSROwY90dD+i43U8GZ6Dr+31SbtMnfE9hCgvK4uY9YVL
Qn6tT52LYcEhY3Hgs2y5V5pFLILIEkSkLsMtlEZqJCN0CkEbXJZUpnPyE4n8kGNz
v5T0vROYLOWLU3SOjRf0jTrcTXd/yvdBGNv0Q6zpgr6PfAW5ezewCRa/YyKOeNF5
lVP/yMu0UWfev4ifceFyj13EJRchKGkgGwB/uqcqdS9+gZ9wQW12emINxSA8sGtc
gAzE/q031itzYUnD5uRmTcuqviotoIkIBW2nmFP6UiZIq0L0y7FD88u5ScU0aMfD
grkfFFi5nl8TsmXJFwaz2UJK4xJ3bzyvLUtdbxbbFcaVXWgzBgt7WJ5lhjMNz+ZW
vsZLLLFrcMtYLyLR6G5yjk4KOIAs0SQix/WgS6/yZ9v145ROyoFwZEh9/4TDuguG
saTEKd6adh+25qz4GbEkM6TMlPlZp+/zxbKQi+tLkY0qvgQrIaRO1g6aMyPWJBBa
+YTjKgmbaSY9pDuohuklcieY3oJS8ZC+UrZCYpM/IOP39aZAsOldoskQqV+GN3LW
mTys0QcXYqUqf5brLR/FKuaHTYM/UFAOipkLPcXt6vKX/Zf7L3HrIcAnQRrEEMgG
y3wxi9pAwsETxhmZv8rmd/WsZO7vhjafIYNo1LOqwbd4Uw0sTTwofHoYN7ajqr41
PVWfontIIE0GyKZ7uK3WMWyAephxd8xXuql++b59KoB2fWNIW1muhDWI2y4irbHI
X8xsyNPtVXeDGJ7iUf24NcIJVCVq8piM0ZIjoPWXYKxTgOxYnuQAwjrtukE3gWvF
C7/QruV6ioMNu5F056M7QUJg5FrDfcWuWXFj6CUAqWixpQlAyGoOYvK94uJ6Lfig
rwh3CgDEbAWJDJHprqdD6BJjW0rH2fl6X0qIFizvlz1gh7KLntjLOySscNH57vQS
/Tli3esNn+Vy3/k3QWyBjYYR/ENpvZmvxaq8jzU2kjDh+ohsy/39eodLLWf9fg+Y
kN5tTHWcDVwqWwgs3ZTvp/21d2UlnDQ9wBXzbwssU1zQVGW+0hSOsg/EgK8ztAaI
4HKpF2B/KD673a1GssOr9SicudpH/HbBZ041BPPyCzF5zo5UoU+ye9/D/9h8Qazb
81Lyz7dBC/GYoc09MgT0xPqQA5r5F4UQUbHhtbc1In4xB/tP4qvOsDJl5oj8Vesy
xntHwxotZPUuRE2aEThmlc3/kcabNq5FhwHz1Ozb/Kyqf1v47qscBrH+cc0wLrRe
VHT2k0JarY21hi4hF80y+2786HZ+zZ7SPBrkmPBZRXsJ0kZQF6bbHYWuKs6MfOHo
4Px+17ROiEWk1lEbca1wiWTrF210h1agsco7HTy76Va+imiQ8oijuQ91QD6OcVPa
yL9d/4gn0odBH7sXcpai+xmqDjggVYlveJQyK9ckLCOeByIzRloR81BTxa2WnMS8
JcMdvkiIg91u4P+O33Lc4IJpPqrVzozznkzz96vyVsN/jDdWyO1yGZ2zAWxMyrF1
1dInBn/3nlA4lfIX3vitGULV39SBAqch4IozSYo2siB72FMEPsZPOl/5Xplyggtb
zK9ND/1b3MYbVmE5dCrbr0B1gVEMKXsdQ+Hnfpl1inohJmY84+JXn46una0nVcNE
B7HWuxT6LrgIldS8SksFKCFu96MmuBDA6fmREDvcnpiXA4On+57toTsZ3XwYW149
cCkC4HDn8lut9l89x7VO/bG5z5ECLAY5KL3T6+163G5+Tf0xIQLIUkLpIntv0AXv
jjErVWW9ug6ErpLekMzJpxzRZS1UXEq/VePVyqgdvkZGGrij/CEFQcApPeX04zSp
kw6dHp031ipm9NNST8bsUeghV4Rt0oPBpQI76/UdklWD3u83/ecfU5tqekCFRKtL
yn74eVfnn/1v/Tc4cExDA6uOq42rRU2KkkUL6ab/wV2LPeGUqLWArCSslMtKC1Be
NQnRpahoLenawKnF3snNzvxmiVlFT5hxIIzVg0olrn4xTOikJy85dWxEsDdMPbBu
vmLtXtthDP8C8RIKh57vWspkdJS2kWRxiScX+iN7DVtR0wBGAyp22uheKZgt8WG+
qS1QrUXwFtdJQ42EAXVr7xJcpxsQCy9/p3OOrXBnVsXSA9/5HXywyCeiJpzLr2/w
ZtBCSJSP69WiMIDh712U0AIxq/U4arYJIAOKzV3+/fQPATINss85GRve1cJuLmkJ
iapPGlD4zvYe2KEUGfy48cQ40swwp0h5cysKMckegA++f1qyDpoBrsk2zyUBmuqg
5h7fmpVUJ9sM2J+9oHiB17uWImaPX2eFyatAmatuPFY/lruc0rNB/SeK7MHxmuvs
z1bXPG1VQ9V1zVFCsPa30MQc14yuSJEgf7ye0RqNIx0Lh3/PqiKceLHwb3HBso68
tAcJmJyc9XkryFv8dJEl98TX6SQpAi2NxkUO6HHFEc/ym2GMKMq5Pt8ybFEXVSxS
f4JI6Wnpkmq6VNKo76miGsWolfLaHUqbZhFZSbMXPA76Cktd0xgNjdKgJgWJP22q
NcvWDcUBixdWmz6oPNv4SR4QwC0wTZZvCuviR8ZY+6UZjZxfAHetfoD8ZPioNP31
JxhhXvcG6ncqJJFgudAjrcLwqQ6Hd5Z34dVtFQ88mVIZnQkjMr97QEAwzqoQC5+v
FipekQnohzOk9/G4QC0h9ZE3dBsl7eFEuOY13NYplC1UQaIx/GATcx8fcFs0rY4t
5aN6810h+wiG0bnqX7qTNz+gOl1+pBMYRTm9T5PnMoiEGhW2Iya3EUNZt6KibyCI
KE/06fpt3R5HfJwO/P629tlY7sny7rl5FKGYpxPk88GyU5B/iL1Uy3bqpBpgNYHk
YT29NNGsKrF+HB5XjCQBt1wjakhESQEqYB2Uqov4cBMcYD+PH7M+nnABysEn8OCu
i0F/0vgWgJ6fkLado6XI5f8lCAo+kVTGP4j0IGn1UdZMVvOgGs5kH2Qa+ZHdYsAE
w+S1/E8g/ibvfgia4j10DuFb/VobZZV+qAhRi3FQiwReEBJb+HSjY7Oq078rp9V7
nRgJ/AeHzFtvaQDvzSfp4WhuYxLHGSBue18KjC635qmMPT2UczYA/AqIwJh7igha
AvwufKOco2uyqNzGqfByLlbqHIQIob5CG+sOLoo/uiyiRej0utOhFnS3+nbaPFjq
w9uCuQ8Rq2RsQTkjMVtDW9/92gfBTzhv5+GVa1boAFFgINNXp3AIQ/5uXlrpG029
RXj36R9zYnSbEhdqFFex0IB1QvccrLvmc6S030M5ZGFYmCpYvh4L27V7Y8m0cjAd
CzkG/R1dXxW3aCn2rnJvaTEQSnKNwhUefvgl6pnrLrU9928ww/MYe+oy9RovReNb
plnYlkhjhI2UMg9GFYUjM5nMHduF9umboyYGqUOQp5JDqWfMRlOw8UJ3oUTthYNC
VdPKzDwRLwqNVc07h2FTMKDqQnumfenIFPqLZDQ7EI6GHHJI7et4DjK7h8Ieo4Ik
bZqZ0WYL0L5Q72QHPMUV4UArOsvUeNKW+B4kiC5Se/rJ9p2wwS3LajnnTz0xxadY
8wUR5W+SI/foz33rMoSKXn/JdU72fkYuLzJzZ8nQC2k=
`protect END_PROTECTED
