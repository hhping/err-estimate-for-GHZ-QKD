`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jHwviR/vHEqZbMwt9DtrOzpACEdRyXH4ygxrDCT5C6g0lTzjhTdRGGY5Dk0keXzq
WlXSe/FA/yAyEC9TWt0PC39nYufoTxtv1TSbm5xU+VYbkLu4Zc3t3f61pKJ0PnY9
GBdEj5DGaT+kvMB/x6r/eMwcsanXg32liZ6Fa4FwBA9GI6FlM4xi13w+mdFwDo6x
9tz3EOr0LofIWGQgZQha6e9oQ0/m7kfCsK18+eHz0ySD5UcsjirHaWGoINsNcfmL
aouGztfQGCBn47KgsbRt65wp7n5YgPDHkrKASk0F561ALgvG4Ir490PbzttNgaQW
QZrPuKl6J80y9vWdZCRJqk+iit+YfnBN3URS8EdhNS/gve0POoMUrOBXbE2YUA3L
cS7XlpqDQAVuhh133HWEmCCippzH8AqjraF0ND5EJl3kDoVbLNYvGwL2A+WcqgSo
VM++ahdZxI7FclRn+o2gFbN10guDy5AFpOYk7vI8YKnwu3roRUIA4aziQOVn5MHT
Y1Pqxc1L0VNFn1CxQ1xf2bZ2432o6dgxX/ah2lHmZs1vowJ1z2Q0ApC4bwBWUNkA
Q0rr3DWJMjr+mD1pjxFn4GbmqSKU0wQ1NdRrUFLCdvB0tDNNAVOUCXS2+cdANTEx
+/GKvOIANGvnIKrKGR4/3LT4P1X9m17xkJPPZ7PfSgf/XHJa3lvHqa32gVHJKF5F
9++2/4pzzoITlDKVptWIv5RoOsgrr5mcGkcEa9IxPgucr0Howh/WTgGl2C91zDK9
gOqOsjX0A830/MLVhQh8kHy6vqyGIMK0CociCeboy/4H46VYy2RTyaGahaOaDaAQ
8WYmQyf9OgL42EbJWCExyZEfKDC3tL1xoQdmD2f9+W71kLgoqbFBhDe4ziATfp8X
EwBbIJZKgXNrhQSpfOnge17YmRNoC4SkiA+Ur013xWqpvieaOHs5DG5yhVIhfhAx
gXX1tGt7muV3XZTVogAh+MLk9amwE0kMy7sU8qrRFc4NzdpL/LdCanUzCXfI8DBt
vZD02OS9C8qIJXRuVANTsp3NC2O5FvA4DNYtvB8f+V+9C09EwbGuYcCAGATaCySA
ikXqYJNCtBBYqphXyfZMw/dlstMG3r2au8CJuFB4n16fSqiZzGIH+326jGt5XEWA
Q2VszpB3hTscfwQUm8SBE/4Kjt95QA4gLggLIugpnMr6AVK3D79jSFXhcealw+Up
jld137G4FbX+FYre+jRknzECSw2vahPhAjY3uVqR8cH1VCDIFKRBtkt4E+i3rUhA
r3GDCv9F27pV494TZg7RpmasWVCXBXPWWwzBDS+lIbewD2gO18i1geMMf/GBHvYC
Pgelj1sYxSswrjnhoqx7SGs18BQ0NQFQe5Mav+o/XfBlULUDKpObESkjOgdh+wM/
13nEHopeSrbIfweQkn9HGgiLMdJaY540VxAPU0/aU6K6AZAnIVskIR4BI4Xf4FFx
yUQyZluYsisOCqWx3JwqxtlaHo+FHlP2siDPUbIPn1tQ7BoZ3m8bcC0J47LTNt4w
JmhCUbrb/KhxhNMncAS0tR0RpWngl49aZp5ScnxpkKrtdL7sGAJ+2EuSOFgHiMtP
Fbv/7upnybvqWNO55HyjEh2avRPQcjJ3AfAaDV9kH00eGwpNl2rxbb1fodsicMgc
sTQj7g/cPmSiEuVy66mWaIJGQdFaut/mHWSDJr2bjQFAX1/7qbPiSMfwil3ZFVGM
oZUNhNYhShtqJPeVN+0cGyZSnPFF6nJJNtoOULdmUeIFCOH6gcEhjcMKit86ZT/V
ucjAcPoP2IT5HOa6DTFdztbOITMHzgq7OAvoRx6UjZ5ykyVMFyG7W1Eng5j2IfXW
6MBPQLxDJSpKmo9aWLqL6hZ7fPlJWSS2IdNSCFSQfZCy5hg3NAKw6eiYxyzsB8TC
MA9qlisIfVNV09jmx4owi20y0ElNBfQ9kSzt1MZTfmx6lI7RF1LTPmVbji2Td+qu
xN5FuuHcsW56lyxIb2yUIeh3PM5yjjiKGOFxkSTifqEYe2roHewC1C0yWBXj/Z71
RyuD7uCxnBEEj2ZT83v6etjf/1NMdERWl68KIBABbgO7mPfOU2tkCQrjuEeoeaYe
`protect END_PROTECTED
