`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zELnKSBJkvcREMnJkpr8//cSeLiYslznUycsn3YwTxC2SueWgJkvDEENJGhiRsQL
ImHFI1M6MiGw3pC2UTpcuJWyQFiDjZCAgQSAdEMhbQ5DwGWrupr+u+u7jhL42cI6
whO66CZw9lbw+4260Hnw8f+60O5wQt/m3fh+iI88jt9V2YsKskG8ypzw19tnTAEB
WsPv8o+UYZS5IEU+niQKGcMWiYNKNJ6JFCi1AOxy/aWq5g6I9K5syPlb0+svN4Fo
Kuu9Pytm6AkC6zDc1Xa/U3esUy9Nd3RTg+zuaff9vVjZYj9hLA4i3hXDSH/hbppc
3Rfce8xgdTdiOLukiUITxyDHdRkOS2zxxIW+1hOuVkMSuc1YBuWs2sxeg9DZAZ9A
mvDXY9fDsA4tuHsQfLHTHXoJcTdWjOCjf/tHhbcdpbAYJZrUDdFy1kdaQ7z8seI1
7rh82t2l44loQsb19lx0sQkp0SHV2AcV34DNIqo3nlKph9OEA3OQBcH5PKDrG/pB
GEsO1qdQ135Xfpanatr3ooiL7jTcBv70qGE7g0c7jFbehddP/9R3E98gpu1Pmw00
ZoEtYqkj3mT3n1VVWdZt4yBbUze8lYXVXkrRJwjdATDdeMsZT0/Uztz6Th2fNRPU
3jNFGdIRvu80Lrqj6H+m1A0GW0iLoiNpzv++CxHHZEbbVqqMJa0kQCVB1ow4s2ni
ZdXkOD0Xn/BJMEWVnf3JtMR2G+ulJc1TSCxtRO9sTvI3unec6kGwTlrelNu7zB1G
XCvmhY7sR8/NPcA9bmnNpiP7/WNyvAbJJeA2n3cYUXWfLzIXEaH4VbRgIUoDhArD
Sh52fo1d9aM1ajxDYdvp8ad5LBNEIb/tyxD2s1NaHjWkZIYdYjO/XvneTye+2rDI
`protect END_PROTECTED
