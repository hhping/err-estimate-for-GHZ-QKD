`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JQeg6E9On3rVQsdkjHDUJoIAPCzC4fMlmRbxBAA0j3BDP2uafm0zt8VNfZSGqxGN
tTD5bjHNxOfF5mv3lpVsikJFSnzAj3090QubyYV1qAZUu4gA3okWFAD7tcdZnBeP
370mJsnmTAbVZSOS1uZ/cWUyRZ0PRo+w/DXKCy5BlGPtA/X9zstupG3XHlrQOgA+
iGC8WuL4lxA7wgnk1asuUNsJRzVPQB7beuDiPheYdkbaPZys4B3cg+wHX/ejTNH/
aWRjhauT+AQ6Qb3iRNsGKL8AK04vw+0K2sv6L598RUP8oVCZ3CU5V8IQiZYhnO69
fng4xq2+jQfDlzf6/C7jqJ9efnmhB5bDhOUAQIR2CEEnAR8GcOW2w1VGmBq3Zyp1
4vaJMFNWPPRMIZO9blD/cA==
`protect END_PROTECTED
