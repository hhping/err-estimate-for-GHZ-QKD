`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F5i08IAEe/+tfIF1Ze1U3wvjnwK07uVqebqNPvXPVFS/SmdwUgEm0Nzp24zsLvWR
sASsjNhjeS/Tx3ulELBKWhjMFzofmQ7UmxLHW/DlLmMtOuAHP2EbBRDr9u4U3fWK
/df27dLtWCRlwdT8CtUTQ06mxIKAS+Rby2fAbuUxiBfegDG7fiVLkKtfBFLe8vNf
Bzumrauu2Tyam1Fty50OmCEc1B5d9/VlVxrTztY7P74CQcWXClA3ag6QXRiaIbQJ
6igoM/OBMeKb4YfgsQhMhTqMzYVV9QjPdEem8loyqUqFdEwN0O/jO2Jthrmr6grc
OeolnJCnoN+uFRgMn/LK2GbYj4/ETO8unZulvJ/x5R5NE02pgMjmBXWmPsh/EBRt
dpKzkKKr2lDacKoK8ww244MKBUXpkqJhjEr4yR83nSpsCLgAGFboFtMKt8xKD8ww
FHHjZiwehGAL5cCqR4RovCWUE8rn6n293tc30LNd6Ns9x5pJvfhzpZNtOuAQ4eZk
+9nuJw8MKy/tKTaMB9dUXh1Cy0tDr5n7ko7jpcGRrdODdDwVsNttTLN5Fl5zr5MJ
p2l53rTFYO4Bx4fI/+PbGvDiyC7/ztJVKXFu6HGQZ2B49sZ7hYaIMhmY+C7Cqv/9
wbIk2jkFNn5tKZkKn1uDKLroPIQKzk6LRb39EMZiIuHw/Iw6kkPOifJSehXGQR5E
/a024lZhLVpiaSA9uNebJ2looq/VovV40teJLU6OMJaNYN2wWSKQaLGVYl4Mec0V
OL9XNuxUN4tph5OOjk5f6aCfp6KR2OuNZLjw3U3kAbBSNDxTq7uHt1sZWfbjjK/x
X93Qt/hdgoMHtC4894F0iw==
`protect END_PROTECTED
