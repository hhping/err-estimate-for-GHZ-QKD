`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NhfZEUYnRInPQJALT609dFPiDNX1BGThCqaIhB/eDoOKo41Wk5TEYNcWqJLZu3dP
GoBK+XxdLZpa50OmSv5m3402xsKQREg/g2/MjnJ/6ZO2an9R+p92P/RD2OxsTufe
ggPtKIcRXHBMx8veXsckN0TcJHOiAvk0QmKZeH4DXi3uypdEREOFvfncO3UGKeGQ
B7r5E6ks/Pc23t7lw6uh2Er7XLpa20FgQFqsHCDWC1oEo3O6Qdhb15bxc37VPF/W
biUJh/Q+jG/mAOT5L8F7o9PAlZjwOzTCpHbz540bOTUC8XpI6Ih3jw8QKiqqBEWQ
bvWUjvmRBQ8AZNCtW0jjbsdG6Ca86nPyA2wyKR+Pz2WKO4Z4HmT20QCDj2NjRzsG
SAYGMzLfanD3k03qGH3FLg==
`protect END_PROTECTED
