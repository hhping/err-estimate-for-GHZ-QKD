`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9PfnSFL4rt8adGz/q9BhbjxQb9IwIeB9LvCNzy6htJGH4qBDsorTwoXk7eFDWFVV
WzjOO/pbUKX50O1zufZMVSYHsUJOmA/WGS0iOYtyq37e/gWE2oO2tGnoOUsHungO
uRyDndvDa/DR3XXtpzGwv3gwNluQmaZdIfzCFau0BaY/W18ml7Ri8QfeUAdU3efx
oqSeyz7RLICE9Ipy6VEyEA66lGZnjI2a/NOpZyd0oujYWM6P065NFlfEiGqVMP8O
wBd6Qmy5FsYjM/P296pucfQ5tWY/n9z87iYnXobLRXpObnAWOXxYZ9TNeaYtJosZ
EzfWjVLCVcAxOV4AMNuOxJebV7Lo26V/0bwzTq7TUImoaorQYguHmDdqfMKCrTm7
pN9ZytX377jVkjg4Gc3YRRmmxuv97wVXla1g0ELdVvEXXST+mdRxhi4ZEGkUw/dE
xsSebMNJdW3bufV3BXyfwT2eH8XsogD5w2IKPlxS+u9EXnR7sGg+PMx8sw9M2hkn
xibwuAvSJ7XzfZkLr7pPmjzFCCVjUlX4ZaKd75VhQdGN58Y59JkdpiqX1endPExV
7gm/ub6+rmplYA3Y9iWEASO2aczNxlsrqLVGF/yg1ukhcPfgCnkRmwBWWQTwvVnm
3R6P4RMK12mx2v536ANI9KTQo6nz71UbuahTIixP8zaPwP9aPmfw9Jfy+T8OtEIh
A1UzB8mj7PISdh1JyTtWgXQSkq12TAL8n6rmQg13zRu4DygInQ/BvUHLW9oVODwd
Nn6HEVe8ttT/UWmBzm42j8d0t3JWInvjLsDJrMztmdQ=
`protect END_PROTECTED
