`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n8HsyKQ3ZnFGPgJHTfX8TQr51A/9OmD22EXka/mSrTv0ILFA103XMlG9OiQ7JxnO
UjNnXII+RpJ8QtlQM3/JbzGPI4KgZwCHhXkiyzWm1hTDyg+y/LU9vjCYv5T9n/kd
fhQm+uuGcZZGVNt2OESswMnL1Iw6UuEJMxT6MYHESNt3ltpofnYXY4Z1G09zH71u
SjndgZmiKiIZ3sk/PdI5JMATv+sgk5zx+f6Qhzj6aYGrJd7IdiUQfTJRoyzGvJBC
gVqFVhx36XLGph52bEvteEbNx4ceEbMM/Jy1seNQBrLg/QQkltnQJQxtXx7DVyzc
3LVQbXvVHMqVV4a9lCuIEihir4Uec/sj4bt+9BkIpPTDUNMEtqgqNztVtvVZ7OUL
fgwul5tpddslCf19SHI3YKRtbQ+MDH1zxtXD9Zpq2XCiTRFXoNBdGn1EInRQMhwO
7LxUKwJgTYclzxOp74/WZh0NSLsrNC1pwI+fy5THsjwpp3m9hTYo9hE/1rD4uXid
AAQ524U8xMV3sEhHz6BR6k1EqDIaB2Sx4K9JibgHFrxx6TEKivuZCnRQqr1VYDsW
`protect END_PROTECTED
