`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BzpnUBMeu41R4eyEi4Qt6OVUMQYNPC1GwLesuZQij7CdlUYfxLEi8/3gMmt4f/Gh
jUZCU1fZEXwUJyuqU20xAVAuRl0UAc70fNJXfbFn/WRvIx7C4qQY4VjKcW5qFT4R
J5IWj/9m24XeDcxOrHBUm60+X7vTNwzA1Wbo0YJmwV5+YPcDJjbuY0JpQwR9IFyc
fLK1QG9XVi2DQCp2hPej1VzfssMckt4HdVaCTvTeD7rOhcLkjXMVuh6gY/0Veh06
45bhVKwuv54l5hTo87+12T/Yjr/DlX/B5RC1U+UjrotfBVUaPZymQDf0yetuOdVf
v/ScfjvIrbQKYUnHG1EbTRli428eZxEDLNJ+C+73mziakc8UyLTnYPsL0s3TUiXG
mV9G5W70vkeYIKjiQLeJNysoS85d5JmglmfVc7UPpXMEp7trQquHk3eNnHs1RZha
JAWSWdqiLcKVS6U+Szb+0A==
`protect END_PROTECTED
