`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KfuHqLrVuM5qdfsvKqYBs8eq2gD4npRuysHIze1DVtve5143GPE9yG7S2UVxf1t0
fJInyY638jhLSknOeqXEA85cTPDlNnY6OlKUFUM0AWp3qiZ/D6pOFuLumwb+B217
afvjQA9ZVmSkFxaW2lPhEfKCQpanHtVDeR3u+2ZS5Fc+tQsQDT3hbynNy57V8WRC
t+/oj8agV8AljLu4dyC9rfY/WFLe4td3Jv2Zn2wKdEBmLmwNNkl3AoZhZiCq0nVC
spfCO0cIQdTmVF3rrvSTc+xBLv1N+2yyhtrjLqZYPyqpcc0Tn7BBs0dAsNGvak7J
JvimErvld0MKUSRBSBUA5Wuz/OTn8faLp7L1MM2QwottNQm72zjifot6msJDoIl+
5u7ANm/twDTwjnRQTpa7dqexqeX2ARmI2kr+Q87Sws9zx4XC3otXGCx4M2ttTl7i
lSQj2b8G9GeYnRCjNwBU6AxeaBAb5B+NvISnQMNhz/Tg0pEzeEeP1Ku0kwW8bNgN
CxcUEG2xJA3oslkYxfKUE91EyJBF3bOACwQ6Rn67KtgnBSqgMOMJNdE5I56PXAFr
MbDfF14KEVDRaU1VmnTeqdh6GC+5BbfsDBYlU1FnO/DHa7CqB3U+tsQLLZ2oecLG
bGoTtebvyZy4Ms3T736UtJ3EJZB2jQ8RUGLdGJxxdPC6TpgzcY2FDols3O1hBDTA
NQJFaGLYQhyUTHdeBZLu7Wf4Kc42/ZyohK7ElF9dAOrdEX4iKmBMYJIEl9mTKD5P
fkoMpDNJHEUk+ZMXqHqaQv/7on73lGlPyGnc25ZoY5gTVGUQ9LL/jG66s9tw3iWQ
FasbeLu/Bq91RvTDtnPjkzxZk5aLsZc+o5D9q2gjJmp06+bNuEPEYvLowBZpVDAx
bi65AE5hmutgg8vZlQ9M1dnaAeS3tqtaasTHvM3i9F0mpMMWtql5434UMQS7Gc1X
`protect END_PROTECTED
