`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QUU1jSuE3vfloG6vfmwRKEuNvXwyZ0uLZWwEUKYtxk7SRJtnGm6KAT7T8cSz/wNl
BF6ptxt06Uf+59DC0eOV9DCKB4Iv75e9EHINQm93A3aS/w4262RZ9CGgcfgxpvH5
adX0GZu1/YQi+VsEAN/oGn9VuMxGDbvFtfCyEWU0TTMtmZ8Ir/XZ2X+HEEqcBhXV
8jauurTawWGSaqBt0t/mSJOTddB4eg9wJCIG6ecGMjSAcKsVxx8DliyH3J+RTXlZ
k2Y/we1lyJn2ydBQASL1En9WQ8x3qSq3mBF2Pd3sdmXwggqmuJ7kWnXI/HuVUR2N
BdN0Ok+fFhT+Dtv/Ly43cgLKJJKz9TlnWFQqtHrERqzqArylkvuLpdoiLdRd6VaT
LJ7nZbRmutpIfzulcNbyp5XUWC3MB3OBwDTlcSem+0JrARyS42SbnfQpttRt8sgR
PybqBfnNIk16fgujoqy7HIC8dEYsLUogSsKG6LcCEd8AYSE17vuG9hVA4N6czZMs
/6KeBTb0FW9twCx+xUNSwkY6KLT61sYcvDtfFYZrHpq0J4Z10LynZqsDWxsYWCE7
crFGNkg7VZwyUu/nRTgqujIujftXu+KmppS/Psxpzff/2FgGzLPqDsjxmiYHM8Ko
EnnuHhnuZ2T/EoRPUTWM13m/XVct9CIYCATEEodfkPhYXLjYOCGdnJ8LcbaUCVeM
hNGobmZwhGMOczoN9akIvi+W9QXbjkMQF2Js22n9Ux4Nz9refpn0ZsHBCZIxgeFD
fUBMB0AMHRpJKjF1SxGyLNjB4ZSe5tQqkVKQ0dVrAIF3+PgPJ9b2Vo/ZimPJ+LQC
YI7wDK64pAR558sZpaEVjWVpg+qVi7NBTA8d/LaAU9MyAvX0QRItGs9HdJnWFLg6
J1zAyDY5wMosnDOMnY0t8iFo67GCFjTBcT1hAwTyKkWVqytrTvOhZ3s3O3HyFEQd
DC6viBhtxk3Y9FiXLPslTg==
`protect END_PROTECTED
