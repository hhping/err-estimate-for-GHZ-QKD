`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4dq+pr9/6vZ5dP6Q2G2ujWWJiUuSUUai8TWy/6TE0/MRJFA9cBcFbycz6xAQEMg1
UbeztpcjAIbdO4HiT71xSmu3EuRCmjUUjzgt9/tvfk5ULhYa+L3YJE6HrD9cC/3T
6WO6nO4u7U1Qj4aj/zaf7K5880MVi6UGgeXAENaeIfiQAOKhM16xCCGcjsuFMW4r
mUxMTJqNBLX1+/34gyks2NErxOcKKz1MDj2uxwKP5kQ2e4SjdH69FC4vnGMNWAdN
WsSVOEeyW3AadGZLh9BKwOSGHLj+yJv+4LllrpasF9BPiwM8j1NUzKOpAPp43xoy
YlfijMwBSlvD1Iv/c5/KLUGgrkHcEXdkUZV07scxrnOAt97tvZFGdSgBxM4EoPui
yvwX8q1WyWYuzypdV0go4MhpiPLeS6+UMGSkz6egHXbgCn5xf1d+azyBdpLqSOIi
xyw3UFcKW+vevWvq18JgcP2hw+UvCkvV+seiXowFEe+r+7p4u8NL0PQGn6ixTo4a
CBU3FaCq3Ujub+fxUbV9zPavfhvYbtPdFm5ZKgoxIrGHMVzw1R3tAX+qtRG8EOR/
CzRAJPebCRCTNEIAlqVaN6S3/9+tv4X2+dQ3mDOfKku8goYhxMqCJ4g6mKTvwLxf
fiNr+GveGxXQmaUzYym8+fFWenIDpkvk2HqDmAHswPfSZ8/ZkZDfCLwbm8m88E5t
I+XoOquxBrpXhJ92759hU5h/kV5IsMo7kVlCWJaYZMW0ku6/zttWMTXotXkOx+SW
8l1HleM0e30kEsY8VaAcAqZhKMxw3MDOAROXxq0c/nQmu/GX5zG/r1jbXS7BRHpr
vhzcTGjuOTNdCasKVuRm0ZWh3OOid1g6OQeHQzckmHx1oHLReCc5SFL8680nYAKH
fE347y8K/DDEjXTQlrGJ//fR/uBBMrpfxij/1eeSn/OCa9J9g/MosAHcwBaayAZJ
lPHx+OPe50yMQ5ih8ncIR58m0/nE3FqQ5kTVDcnAQD6TjgXGlSTJp2+Vo/qddAf7
V+6TC5V9sT/T1EXEZsdjU4Y0NPvTYuy0gEtTXRDYOh5dXnGXJ6ANuwN1jJ8V8wfr
ibsw5IQC0FLqOdefgJvv7GaD/NKwV61kY17yjtxQfJVVvF+e09L/Rxb+fmXXJ+eG
e+98Dnq8CpkVx6GYQynUcs4ZwpV6UX3hh+2FBxMl8PEinfQz/5a3EmIqWlUi/CNl
cd8/J9FvHa+tmTooiAGifdQ9Ks1C7J6+VElvin6vJdAWJqMHIHFnvEgPIvGyC0cK
WyBsFjbhw33HraaVblS1ArLYCIZfNYTyRnhNWj2BrTXHFfgl022Aa9aQVw4MlA4d
3QSObesWcJCDfFamJT+Y6cdVH0PqsINuHagZsCt6wxQqpozfUmtOAKEpPRMyj1dN
KCBnYefkDtymK4i1ei/9M3izXyE48nX0o/0Vv3jCLnNqzmeu/NlgyIqlBodBZw4H
i2GnU/fIWkL0KpL2MNqT5ovDDUWI/6pCVg2VKPtmnY8ktXVI3l9emK+ZkDVpqoiy
tf0kemqevz+XkQlm9FQFRmQXOXsS4dS8RjscVlTF7PGurMeCAOqYc1N2HXXWqm4S
2iV9+eUHZHiOXzcyXPRXeTKpe7Ao225iLIKIG/XwRbwFaYC/xzXDG5JOq5ov5dQ1
twok+8XRt1eWcYGoH61/u/wDEViLqhXhSVVY/0YLc31Stn/EVr3Kq7Vz71I2Mel1
iNbP5tTGZs4qwUWn1kE5sCpO9iIoDsIJAg1mRiQxhjOeWpwrD+lM/mGgnriRU2k2
aYjLuz2Wr2AluKSXSGmlccndC1eHCxGxR2KBlm8004ci1uaXbGXRwAYoSFrkA6H4
r+kuQug4shFnBjOPYzMnvt+hc5reGeFIVdEcIUglEMP8QOLgGdb7PP+ytLx/jVKl
pT2TZxzCcrQAUaTfCbmbJ1ji5R1Xq0w1RM2/QGb/lPRdgRl8qS0Fi3sYFVEeSahC
zcR0NcAdWRjTu95V07MddgmSaAIad7sISl93frwnAUDKRJkcxC2ZR0qRn2P1sCAb
pE7XIR33al9jwf+KGwmuzRfIVK6xkXrb2ZJ1PXY4i8ffrfaf+hSOlta+0LYYc0e9
EBr1d3dIx4cG5ccZPXbM4dUTxU6p629uDW4QBTncgU53LXuysvrHm2dh2Zc4WS+w
E3c79bhcHgLpN0tpkh80ieuIxkweMyo1I4sLDWV9joD+cECHZGZhKSO1V18mPyB+
O8bscsag9zx0uogftUiN6nKZqQ2vPVfWFSVSDe1VF/uYk/m1lPfKxZGxOyAYOQ4C
xozDN14V2xwSCUyK7BLehedaIKkRf41vsjly27k1VAmNSKFd9w3BJwpDirtSH1WS
IAs/Yd6MSzyoSQvro77FoFGHfAqgOWv7qp2ZXdftnRNz57s0M6D8b9VanJpBpR8A
G2BxDjGmoF2nR5H91AC8IFu+wUrkBvs5OL0s4rKJE57fZDYqHRRFsjSxEAIOFlOs
Q+2MoZwvAA7PEytyZLnrxuS+JUv97K5FUa2Kw+CwdgfWTZICmGqkIsHr+oozl09b
k/rcgmEYZwfcdSRofJo1DLNRMWxD5BbWXExUr27TGRZdPbsiq3f4VVJ9wZ1bUbcm
pbFq8s2z9ERXj7EZWRDqX8cos2qh5MFX4TMX84YldIuoxHVUEgqYTrHeNNttWCOs
GamgKo8a0/idxUeuxh+72y7mfNpj2erHFmt6l27IfqP5XwUooioRgjnzP4o+DV+S
vcAy4bV4FDivH/aHP/AFxaaLjTrrvKowE+gWk+u2cm9nWQug7n/9bg/bsDzbCj4O
gI1m2TGYVvGXxBQjs9kFyBkgavei+BxjbG21SPNEKOA13z7iHMP+CT2pQfiA99Dm
nU81dVKhqH/f++WIHcXDtIRU5BXjQOXYkUFppSuqKfNgNRJASBTCeDN7W9XN1gcZ
b0+WxpBwmHYoQm4S+slwqIutdVNfB0HWRiYTg81bXMjmfJrsvchDN4DmzViQz1YA
rJbENQsLz5aeEXyyKaI5UAYf88bGKq6CahyTa8GGbxPAktQf+olM3l5lxXhrJWX6
UhEk4O0n6YslU97RnZ4szyhTG7SH6Mvk2E4eAD3jtA27G9I+TljgmW+XhmrrEocB
Orie6EZTBH5cNmXjqjCBFT/k6yDWF+v3Ok5pAsqhqq1zz4Mr3/R+FGMy5RiezJYZ
UxdH/jEZN6IhseV6AiBBhZ5sdLJehGJr9kC5BRb+oPy9ZwxzmbKq6YFnrD5zK8Z8
6SdyoEpKe0HfMM1XK4ZGFzlJP1NUQEV8CGeUgw0uiyKtV1t04pXioi2IGSjfBlRX
rvijiSc1oDa8c/FLF5jnYnmOb27mMywb9+JpzVK51KwVO0qOkmYZyqfKFot01nlx
DzCBvVcP5uBo6HQkOquVFEemb4DW2RMZN6EAideJffwq7ZiYA0I3FFHH0l0YIkWN
EIUAy9yWWz24uoqnKkGh4Bt/GlcqsHNFfOvIXv6br+zZhgqpNZmFqCsZ/hCbBGY3
idz1coY1+t1uOfbaHiH7LjK7C1T1/WBxPm36NpgQOABNWePuMKa5TvwSd0x5YQfX
qW061cCR7tFYl+UkJAbAECCrvLVMYeuEZfeUNZiolAwU6WHEniFoWH3UUIIp0Xe5
UZ7Z+kRIa94Eob1nbsQhuGRuJDMGcE8t/Cs8Qp6KC1+Ixk0eBuNj+nP14ISGAtGu
I6tZ2eFtkmcuiXO9r90l3iPXEDYa7kybhG9b8r8s6yhRRGfEGupMUn6ktctT5nBc
+zmg9AwFidaqHVtZBLh6yFAGqyY/4Y7r0OazShOo/iuk8Qhjz3jaMAH01Jal25g3
IgoHb5fLK9vBKt4KyGV7UfFQeXmVw1hxzfywahCPvztPKI99+MCt8rxY2/xQ43QQ
AHO3Iy4GDmBlgieD66B+gp5IMlI4I4xA9lN8gvmHSRS2zshFWpjXpKVHX4mkCpXc
uYFPwy8ie8qPiKARFAwdtGz3G5gTzhxNWw96SQwF87RMeS+nEGEjkVFi4HeIx5qQ
E3I+Gc4iUhwtR2xRL1G1NocAJBAEaPolLAamHrUmAwutiL9QAv9yczj3/tWJJxKp
QGwtID0fVz6XVy9g8Wfi1zdN3YwUVRGCNfC+kL5XpNmveUT8JduLQVDmj/bQ5ADj
T+Nq9P+1lzNpdzAEqhLVmNLlrZtv7d0ANJHID2Nk8UYTWjwKc4gLYBgxLAgBxvod
ZIdoCdT0WWTd0TKCySMXlNpAIUwm3GCAXDysdfxvX/V2tu0k/1xEIFBUQTHgbOyu
Q4mxJiaCQeEglESDKqfYBVf37d8hQpwASi8Y3Mjp6vafBitqXoOI6/uj3xpRE0ay
tRE4/yp0CAMxyjxbx+v2QdwFu26e9AQujy4W/sc2TGfQYztB334FJd9OBlCcEYyR
Hh/T35guUqUxZD0JSHIUQYlRudisFQo00oBD4fusulxNRfL2rQz2kq9d5faf6JXC
`protect END_PROTECTED
