`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pVnK6aVv2ycRhne7FNCmFdbb+DRbXiSHF+b5oojXbBm1lNBk+NlQeJMYIQ617PfH
nnGtoQ3CYjcFeTxOH1Q35Co5hxU4pxx1mBvY3MsDO6r3imU9uYfWxY7DVghjqCKW
EN2PF36TnRU0LlMvOOaLawSPoN4fYjrBiYURwwvw361k1Zl+Z1PuKyIVZVKispqz
5GV58jTE2crIOaro/q6bc2tD8tUWRlXvN/NZxh9OGD80iQ593GKZn4ugPTuftPUR
j2xFQZCy7Aw5KpHRNmpktPvjZCvoGMQzjha+6Lh+QkuzEN7vwdcdtaNanP8g5f1e
Fl9bvSbPPKfbRxcpg5mRRqbTJvtcDYmEkYIUCk+sQ5NygksGu5O+1fO2VaD1ZcR/
FyW6xNV62uG6nCXAbEVmnOWPSFA5M+fO+ByvLYT2PFpt58KVRANL2rdLIJ+G/vFb
+5zn56AEkkChhHizl7OnadAuhUoj67VQ8t8ffF/I4kbhP0swT9+AjS9JiukND3/3
kDLvsUaIl9NZpLxvbVNs5qE1E/cnFuL2K9nkEqMyz0XiyXebiwtgT3zPo9q0bI41
X6CttnSYDD41qxrSFAFgJjVxVzRo5Vs+67Caax0I3a0tNIWGGCrmmONMUScQzrFa
D4usW7Nej/v737hk08BChbmPfV63w0KOzZZbbCBb5o8bf1xiKZ9S7oHwWrbRbXk2
N38GHDSOXo4AhpQ2BZhASuFs7HlKLpRJn67kVBnCZCtU94f8ANeRaJrwmuqnVwCw
bbJF3eQGOiG7aPh/L/dRNyzI4CcQlXwANNSR96+L9zgBD4vlS9dJ7NBayFjM/BxU
HeId8FD0p5QKwn29H6wuIpIWcsyoWcV4iXPuPGqGnOU=
`protect END_PROTECTED
