`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vjs71++Q4Env5RmGOWJ4U8iRAfylF63cSTDwUk9spgqlL+XxgVgjM8d6dxuzxfFz
45yJeX4yCl6Jys6Oo/6XO9+Mel4x273SxXuzawY8vsYq06v9aekFiK9sBdn7ZCLP
UXHeOCSjW9j8x3fP4Lz4cZyyuJLF1FjSUfKTMedxTdvmlWerUo/Eo/PepyCjmamE
DVo6Zsrkx8JM4n+peOy2RngiWcZSg2xlK8qglWOK8CQffQWv2IFEGJbtYVLtYhsy
P7ErU+wsaKol/KTG4iOIyaN597VfWgTLjoWOVBof9JKG7wLoYgxdlCwost0cVuSJ
uNv/IXp02TeM5mqf9FipZCfbQoPlHxr9azB9IWjfpGPeP/3YFxRRDj43Y+QOa8P9
QORAWF6P4DRpA01Bdi9tEXhhoNP5bmRJFNFocjAZfYdkUlpIbKKuxcqYp90QXfMH
gq4YsKBMabmvKa6Plx0b+zvpQy/TLg1wSrT3a/eO0q3nKM4vZuVCg2tXDQJ+lOww
MnAEQgWDdhqxmkM3IqAPW2BznBi3GIaUrgw53wawUvK4B5mpZ/YmNrlpr3Ou7u/h
Emg7+hpG81evaw4C83lf+h0T8IRNL/Wp/gq/Ohyfl8fCZbYJ/+FVZ9OWxI2JoaRw
C4W38zswwIAJx+Q9/qlG/DCQIQloXlcsLMYb2QgFPOeJMXoj3lZhUkhysN/qt9bn
HzL56jqsys4IYEXc8CLWNOQP8keRh/Aqu9e/lpmW/hNKIsmKbknpxD8y2zOmMvWY
bWGT9V7Jt4Bu6YfD/E/NLPYAFU12NMIJpsfyJriajRAivM+wQT04K2s6xwiKDkVo
E+nKSM4QN+nQydABCvJXW7xuaq6Fl3EbM8+ufDd4NvcDNV7L9i4f8rwz2Z86EdJt
8FSm/UCidPOprU6E+y8cOHe8SZqOVjtGES/PX1C10qhKhkj9PMG6SLbJazi/fhg7
`protect END_PROTECTED
