`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LdP7iDzdFfS3Op4zKOiRDSIN5mBRBt9I9Iy87MdqZ/nrhTWrDtd4sIV28DB5AFUW
OQtvmo7cSqWGzZI+WiJCYr0yibXWGTi/rDggyWP2hIoAGusX3nlQ0laW3asrXIgl
6fl8zCWWlDtkJdLEbiFc6DUISpBFDvSrKilnzyudVexyrv2F6CD3DH+7L67nA8q6
tAzttzMyb455UOFhOPvn+SUr51+nLCimMHOmK5pqOak+/uzP8EAN0lFjmKmpY3NQ
HhIs6VB/qaumqzhQKKzhZt/J/IJ4xH6h+U01tMeD0k+pPXbDu14wt8NRBfv6+U7N
eIULmqU9iJzfr51IM3qrC8NNUXyrgpDcmZdjZTTiAnhS7HMUpwdQnph6/SCm/Dvg
EX447FGsqBqTxKJkXB0lGPOj0DG4bAJT/YrrET6ke1TMUyl8ZWmfaBx4oQdF60ob
16XEhkHwcvEqbP5qE164vqGeSbPMjhCfFOP62q+BTTy2DaGDVtwddAvTAEmJmHj2
zFx3PKU7CkNOu8FReEN5NOnPlEC7PpgE/7nGH8kzfhi6zGPki25P4oOsKW9BOJUP
n8PD9a68SE2e1cJaTMsIfvaR9PZ1uJoQa8u21ChN7K3g7NdRL+TExkpt0h0P8SZb
2DYP5MCkcGO2fsC0E+5G4JPVEOJE3srgQFTdc2319m0nOiMC0rTIM1m7YZjXhCVG
bjUcsaCQVLT/cceWJUAuI/z53I/mMcP5/XfbR57culcLUhGbomVI0cwLxFmz9KhR
iXqh+jxlhiCYHUHDaF7ZQRGpi/MQTZvMQYI0ZFtNruSKxuIUVZCtvWX5EYg2wsHN
NUOJYw0AUSsW4sAJjcARObGm/h+9Ydm29bbcc+JAYRtVJcFsV/dnY5Cr/IClkOhP
mWn4i1OdqkwA4146bLT+Gw==
`protect END_PROTECTED
