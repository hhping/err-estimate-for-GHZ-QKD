`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/HqOSm17+7mIHnh6pY4y6Ps3pSWAd0+3Wm91nTx72r4OMtU812C7ZhIGzlNoWdGR
VQZeLSzpwSYikyCuPMzgV3QvPLiOH7mfJVDgvCPg4Mj2jyyswhGqbzIn/9co0udU
n8fAg/qvlpj/MK8s7iJneNCv7HXcTl0R9XoYO+0u5gEZ5uR3DbzBgn0cxl06IJu+
PLHFIRW86Aj0SySaj3Y80Yn5owvpqmX3J6XtLTgzRd8UC0O/zQMxy0ewg6bTTpIa
404/BcC9M3PT7chhYwEyLhjMIrbx4O8RnQWcu9Fchah+5356wd4XG9RcntdPtIZC
sEJgFO4KKFSJBmPoQg14a+4ZFHvwUOlexeS3yZrZRpnmLhwcSG6OIZHR/sQOMknF
nkJUE84Qiikp2EoQPvuUIUEmR6Q8J6apBinYfe/Sv/ZFuOfusRoJ26HKNQaYPi7k
KTpExJ4WY6rjs9kJtA2M2gnJVuqL7aax51uvnoTh9Dc5mBAz2q83AInlnS3em1l6
bnaxvXWnP2akhcNGCEG7atMF4PoK/8qw9SNSarUjN4R0unfIZArBy8ME3Zpp5htf
zsJ2p1TvIRfn8U++RsWLcwViwmDbAAvQMp6kWcT7LCixlIc2rjPh7RSsBwZXTmNd
PrzK2pm97tV2n2KOHNkjxkvBA2IVmgD903jxp3PY6aAUg2A2mC6Si3RfhHAVJ7Zb
hMeT8ccJXHN8UncrD0DH0oO0P0zmAnctFsmtwOIQmBRn+kh+Mayc/fmcG1x8eI9c
OLRLoItsEjh1g1idsapq2QpDPgm0IycCjfM5R3QZbo6p7eUvOnEyfcDH/honVRHz
2vD21bt3oAyqsaC2c+oThPYfNyQmSHFjAFOhqzEpHtRAqPKm2Xf8UkqA+4dZkLVl
2BC18bzt9xSsezlbsEBbzzhneCX4D/Zd/r4f0chUdQFiGUO+ZJNh00y0heukJjey
ZEJpQFefh+YckY03lhI8bIG32uepji9dAKKBUI3LzzoreQmu9FyA4E/bmuPDLImz
F1lNFmWJBVXPw8fMOYKjT7xf1xurtO6GwACS+2jygqX08rxwh3RVK+QDCZHBtgbI
nnmBsmk/Dav2d+EalPSgZmfjn8Ldz9DsZmaieLdxkKwXmHZ0wMj4tVfgggJy0TP9
ZwKqQdooKr+8ocrLwk8vLi/4T5v3TKM7srbJkRYdNWdMwcsqa/F7yfifR6O7mrot
D1TApsLa/+cWxItFCC321k3PWY9fWnSgnKdHZgCDiTf6Gl2OxYz+Nw4xCIPava1v
LD3gv600aVfeNNxzTjZBk0eJXyHBihVAzlJ7oh8574ywFT9rr0VZ82h2insGxlDg
5TvZRYfM1ydloM7e3RHc0plFnF6RMN02S4pKOtTVmWsvdzr6XW+FzaL8WqEOXx7B
RrHKoUlisiVu6tANNZwtBAn/fHaHzLkucqHYqC9bZYGOYrbXqoAdhao5hXzJCSOJ
00h/6/nxtZdq5EmywthSeu5TIpA1o0cceB9NjlySYFL/ODNtVLBd8VR9JA7WxvDd
TmYycgzUljvX3zQZ20JKMb2ec7MCoENGQfOc9+By/gEfEFZfHDvFXsD67Ngz56/F
uyHhfYhj8Y4hkFCJQEkVn601hAOc0TGt9xxtvemgWz0EUfddhjI/U+A4XMyTkvsB
h2xzyw0dkoev2ESEQ18bxwBERXoGPVtvO08r6rBcfGeKmsghpH3RB/2RHrB/ztpD
vjNZgaLVab2nb8yAATez/VZi6c39zeLw4CxzQe4TF814T0MNhYRTLTY+lRMLq6ys
Irw0YoNwe8IU3KDz4Xe2y19SDs/OQwzxM4X993OXJW5u7QCXK1jLviY+a/q1/FQy
jREE06OiTPxktN20DmiDpg==
`protect END_PROTECTED
