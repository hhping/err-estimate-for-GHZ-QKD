`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kswxpyxv6MVh+X9AeG6XMp5ZG1upBGG7A+7BUEOxUPyhysUSBPG0bVAYBhcB4WWY
s86hM4AWFMIXYR/l2jRm4r1L+VZ2J16C9Soxv9yOobqXL4I6mPb7QU5FT35KJ0bB
zudhtwGGt9dL5ukNre96vuaVqSkaPFZVUW+zwf0utgLxZT45V/ZezxLDenF8NPEi
`protect END_PROTECTED
