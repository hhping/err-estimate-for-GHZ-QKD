`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WnNlBDcykOqtRlMk1VeVKt8cJtDs6v8Jh1DyPBxWA2NnKs6eX5L+gDAQMyrwel8V
gwco2kvPQNjdzS3IvONXKezunVn9sRIGmAXb59y8YCjCPRGYfdJ5FSecGGfyhuqH
IL7atVRjSylYTkmAUhj5LBbySltfTB/pNWxu9VWuhP8yt2db15hVRI68H6Wc7YIR
dziCvlHzoXfEhTlVKu/+t2t5y62K60+oxV24PC54/LhnIN2sl+oh2cVQ8rDwS5yg
9Ryv+GvbJHU3hluvHNAUwM11poUMYBJEy1EikQuF/OsGsrbWnjggjYgXOBVf9nVH
dXPbD5hinUauPy7ol57jFGX7FF5jczqG8CafrldFdGJg7H0vsqQ4iDHF5XVNNCOG
DyyBrz1z9XmO021xY8hgYbj8JGQN8OQjyVEF3l+ot9Zr1az2Hk/GBs+keVEilMsU
AInGfbaibnWXcdwVx2BvzK5mR2YU4En+TryMCawKehyjKdCaKj477my/68WpzVlm
SB6qlL2qss2mAK022gRP1/jKSG2SayNLD+aGRWypP1MxvpxTohyz5nzmY0xWA8l5
H0jpTwJ8bDk1YGeN4DQs1l7rWIdxLWY/B/ta4teNAXmPYWpIcRMGGo47l8hNGUY4
pxpbvgeS/pg/1eW9JmTLl3XNCMS3hIY1CdpWzyr0Wt2W7IC3XvwHEAab+a+HhgmU
M5sS2mcS/hc+JoNSeaZGCm+DO1KXtfaTk2+6nzuDacQCzsuURO+znQ2KuDUdcJNX
G4v5G5tNgrUKMRREyS/dRNk+SvYPC4w4u/ybpfcjWUpBppdFi0Ck4Ny33eL5/AdE
//tTWm3oTHsgGzneVFpUUdURKOovCoRdCx0OsiYuytffgGIdKya6jwQVboAdO8kT
/Tt8RzL482E9GzctkgXKtE0nJ0cku6vUytZXvmnB70v2csMab/hi0IYgC/37BKRd
vYylcuUxrMMJPuSIXONjIWWqFvHgtaH8JDYtlnSb5s+siCSMU21Wq1YrKUtUzCEb
Xe6hZ6H776zRZzAs1TO+1jZx1aLg4NJe6iXfk5QQkbJERelwCpdhdA6w0xKnCPHg
owrc77OE6j06eAq9YqenUAFnFekrhs4g4efv3JWeF+FqwIRa1f4VO8pCxERzk2yv
h8lnDdsyyCYE5eI2RWF3zJQgMS8N276UCnKL+saCwc+kFomJCuNluwUmpra49q0l
cvGXlYZOZMxwA9q2mcMce47wFdxfIg8x5EnzRwv/l4pjwhCGyGe8RMsF/MYhHlSw
0mghtjr1fNc3WIGRr+YbKauwqaREboEb8AsEkk4icXQ=
`protect END_PROTECTED
