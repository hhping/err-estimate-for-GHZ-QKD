`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y6XFRoimXMKtK2V77gZ5noffqMrdYXVEW5XVap+q6z9JvovAXo8GS0Wd8qXHpaPd
ETFCE0myr98wsFvGsIjJa6aD+XYuWOWcLMD5GwYxTA6R+fs0N4brCk3IRjNnx/LP
OqNgTfWo080DL6e+rQOM+oHa1XRfFb3C2zPsg5MJ3AEpehMEuD6rAnthtI8R7RPe
oz43WAeK+IjePsoBwQWekkBlzgfNGFI2K9+EQzD1RNRmcVAEwPkA8HgSQVP311vz
Zw75jIPuUHq0vzRyqeHQXjQiWhpr30GeYT2TwuESwoPK/IbqWVQOBuPqgQzLQuna
iIOwhj3pQ9p+MGVEZQGRldCafm89tK534ilDDMBxzHFMkquOPi3NbmS4A0ceK55s
eo3FIQzSQUuZFqPo0dBFqCLsuD1EQepDFuIt04O+9r62f5+oVp1hpDqYnXZjSg9/
umWQyqvXR+9q9W35gwWdQfsDle4pJiE7unO01E1XyS/oOi3fW/grKFIXRTTvAh3E
I1b524szJ0dXe2qDTH1gamYeVli32XJg8guPIDb+XsJClfeTNXhnGEsseDSGUFUj
6cgeV63UzOOHiilKKMbSFsYSZtJCpH5KuyuHRRTYIqZnARpcPKcNNwAbn+XG1IYm
iZHjPDX5iGyXLdSdz3SWSLiw0jjbJ/5AADgMvYSgAchgMDAdBrUE/VYqGHAJzDZ+
ZaWVjW91t2DEhIPqRHkbMBQxTzMFyNZUJI+LG+z4m7lTe7Zzg9JF3uDduK0GKtBV
CgjBV4HggzhsP5PcjS2I+EA3/rEnwm3im+zKjqprBrnT5MLPLuRZUw25f+kvdrMO
9kynbPZ/ZuOmrVT9HP9599dolZx8oT+Xg1JTeW4pONxDsBbrfLFZs9SRLproibTI
aSDnDb5qm8qcvs277qlu27DadsLh+igTdSerzWXHwlU1oIUn1pRCRXpNghdYNHse
VAbSs31DcTuy9S36O4pttJN+PzY4vziaas2bpj/cp5GCaE3bALyQadgR20CFqIjh
X95GAnl8w127htid5rzWXlXNLyrtdGRAqh82skTFwgIleZ4tyJrB5Q3r3WfmdbQL
KH0Q6Q6soO6LQSpTzAE5TtVhGTMxYqdA66swda3AdCzZxaNy1uONqDKRLF8fbrCd
9fyyfDNpvbCAVBoZ/S5x1L64q4w3gOL9R2TojOVr8SX69i8Hav2dU7QkxRvzjF81
e2tzT+M5onmqM29op3rbBa3x5AAd5WjzWIeW8aL6hOb3i5cuzmobiUzIsZl/dkQ6
av8Ss87Y1gBMKCfWR4wlNnAMmyhEY1LIREhjN6alTKUugXogJ4mBJ7p56lJVP7Y2
54sAZQ8d48mVkWbc8/+SeuQwOCBaVGLb9rgeQ3yqSY1G9glgbSS/1rxf4t1LnzwW
I6NJKMZlMnm5dfm5MpKQxsgqlubo6JcsgSpNqBrwEplZqnzVGKeronwkVmz6mrpJ
YbQOR/qozhN4wacEiH/fJIbyQvFngoaEmYa1o3uFKv+5TETjZgYYULvNPNRfjacW
q1KlTO+h1mohI+gcSksO1tP2w7GaePMqnmWKQj0vGMoTyZtglNk1T+jARqHsqgBO
yet5aqd+753wQK9GbVLC1tgDVws9jk6bz4cAy8WzHrwS5f8AYV8pgLHl5w+TKWzQ
SVCJZhG33axc2Cl7tMJ4rNVKRHgcKcafZXjaSe/JpNEKq+avTOOh1S3keJr6kb7g
vYvi1OKqZL18nJz1HSo/Nbzv7kKsMXjHpbu9oPwyqK63Eg4Rroy/G5SDDAwoHg1h
WFVZl1DFcbygsbOHeMNNmvZWgXdOO8e6cDKb2c174lyPaWmsiLiu8QWh3bl/ZLfI
Zd8z+JS8B+V/rJZi5ovMHMHzLc7QKHS+jUJqdDAExO8G/WeK9PuW1gLHUYLXTk1k
tVlfCgtNS6jGD24pvlnzIcZpxXMv8HReezQ46swC5MJJEi14OEXl4VH7GSxXRCAO
F12mihoLFLVF0j7F9QyT1r1KzRcqo4ZXT+URq6eW6t8Rk+fkmJUgKEAuNtR9os/o
CDW7Vy6El7zWFvlj+TiPOcmPnw/sPqIysWlnZIen0o81cuuvaFkqQ+As+MI/Q8aH
oWiuS5yVDA9BB50CJgrJ+Y3iDBkRGS4KbdvQqWurXKwfVgrh98TscKI9rdlzrV+X
+Zd8NtHjqCotkpqoK9mgKH0aTlOueRbMfo8r1xhGt3knHiyJusPk/LVPyY3eZvuv
Yd9KixuDwBBF6mIyvjw9pH3wXxiviVWKz39wPBU+xQy43xG3b/rWnYqNLDYnqYRt
FSOKYh6PGIyoi4xkiwHWQdA08xNEKd76rvVqvdDTI3OjrweSDQt65t+52Yx97Rwz
GnelOF2Fp78Evtl321mH8sMWsB0zGBGkkecvAfrcMLRshtG7Ld+fhBCEPCo08spf
pGUwqhZPsA6RD3jUwghwxw==
`protect END_PROTECTED
