`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GDOloKxW1XP9oyAH2Mg1jPcFG+BX3z+Mvfj+i2y/0u3rG5hBPhwxGm6ZP2Oln7za
GNBTT6lvHLmMxFXZu8ZxdoILtlIn40Ex50Nzqeo3lMZ9Bl/tYsNPYqQI3SEgiNK9
F5BAIvidEZZkuegcRrePvrkRly4c04xX1b0EYcA0vDPFuueY5KUzI3yqJIh5ghOv
RG+W4PcX6sktDjAvJ/M2AQZ8YyQTkwLFcOcfQ46cXEr4MRRhpgAoFFbdgusci5Vn
0YqOIzwyMBvw1EwORp3IuyZkgQve8HVL/j8yvXdnJFhPCNlFAS/nrO2XsLpSA5Kd
sUDGtzYZRnnhHrMZFzSzgSVRLh4eC7sZOZ2hUlWhZAXVES5DK9tepChXyu0E9bYs
eYvgdPl1saeoqpnuRAkOVQEP/Yrouzn+uZ4Y4W1ibhjB6vY+9yAHcFzyQyz1VbVL
Xdw1/bqI4yMrv7a4YA+FDPl+rhSIzk3AFn/J/8jeTSz+buchBQnddg9Y/b/Kgxh2
FVRYc2dZFhgcO5QET+5LZBUmXyMWPBYoQW92Ig3wCdFQrw7t7Lzjm3mwtrw4iCBO
EzLAegHQ/6Dp1bheedhsp+l6wgRsUO3lLzWnVFsQZZj4DuCZ+A0gbKUSKsN46Gcn
OhlHvYZmtJR6U5Q2zfG+L3zMfzs5PXrFa5G0dVWWp5lCiywltftyL4FNMfWuS06s
ig5lG0Dq/VIDbNFqLtd1YuvI7qxmxAtKPm9wBsj7UbOjEbagkXElLUwccMPDXChX
zrkbv4uOinetpg2XUe/IYD8eyhONuOOewwT1JeBXP2Vg7uk40Bk/JtUd63ZFhrdl
OfdbSJGXT5VOH91cgPewEgHGYxragC5+7M8EVO3ghAkJDi+1aRp2W27QzejiHB/X
7OZytekmwH0SrT10mUDSQxJbJjhA4/8pz4HrIACz5HpgadSaTNZWcKBP5JS8O2+1
YpLAqC9tRj5qbjP9tEjn8s4pZFEZiSnojTg+/zkBppAi7yNOvnaAG55cFI+UP7lQ
fF5c9eaOHi17p+4zBSQrkf8sul6TXtKYOvAjm2xMOE7lJavWKqA4jT4eiOlOenH4
lrmJQ+hcLRgVNip6LXhA8QUjSXOtzYhL7kGUyfS4NNuJeZLklXKbaSOh7Pjp/3+u
`protect END_PROTECTED
