`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4ZTQh5dW9RBWkHry78kDEuOUvD1OZK3bNh9Oee+G65GFbtn0dNjnhIHeRroUDX3P
md9Z+0gdNm/XrdEyPfwn8A7hku64mMXJ+urDcPIYHUmddhUK6xTjsZuiX+wYMpFM
8tHyybdMFFGEgJlp7n+9Y4vNmZXO3b38bKmxQaNNAJDibZLgfxwCiGBVpkhWQpBi
VNteq9ACf/cAZnUJ0pEiGuHqvHmnI3OCRx0ybU6XoebHb5DmUiM7oMVnjWZclw2F
EGWZ2C4CulYeOvcD+xVsuT69vzZqUR1jDawGPs1t90PfSLoNwWZe9z64tHooqrby
40QtV+P+oE2uj3fzcns0DS0qKb0AYM1yEs+NPDzvxZ10T8r038T2znz6y5wXyIIS
/DlGJJLMYuHMjVNyOGvhfGpFqrtw8S4abmSiQzs8da1NEx1sePESBC0SsXLVAgo0
vaUHFojyQGrEdCLYKZny6XhrpGZiMMMlzfpHWmLCTH7T2Ifi9ueMODLCK/Au6pho
gknj27Z6v7NCllDpRc5I+JzyCRG5h0/0AdZghNDCssI5vYzpSYQVCozljPlKx5xE
8IpSVO1k+1iAzjwVYeKHW3RmE5tsX8Pn22i+Pxiq17s1JNbCy1hUpOPb4CWstFzB
XZGALxenwq023b3xf8kzSOjh/lOgGbiZcHzFIkWnCnoXg5eWTLnxtV8ixFH6f8wH
kbV8edUnXjhfg2r1j5fxzbfqWBgRpoRzQF3HirrGtyt8rA6iHFLoUhmHZc4huEkD
UVD7+Y6u1CGFnr7lKP01Y8nBliPWPgBQrZ8Ec3ZHMIAlJrdKUgiTGOHoRiBy23R3
3TIihiePyKoDlW/NNwUUgBadebicAR0SEq64INCy38axJqYBGeuHq9YDLfObZNdW
wJspQMvybRwKqkBFDTb5a3CQy1yT6gh7TY0t7VcklACaT4UYoJkyjxEDF14DW+6W
hP2kV6xmweafQijxmaA//+EUvx0E+4KK+8TYAs/1R47+bNkYVlJ2mxrQ+U5UL1N0
KWO1DGxtrvpW7LcW3R0oqTBO4tU6mVyATTzHlNt2afLuzjJcSq1R+liuFrTQm+5T
ZPaJJHWXym9hMQ3ISkf8lAsyUE3FHF/4vghy2EGNieDZOF42ziyYInO14Ko//cnn
g1zbiSbKMRHoyyBStTqB+GI3Veu560xpW98LR7CnvRD1Pni/2SUupXLNLykmBzrU
ouuSpbyYZofRj8o69eCIDU3id2QkeuhVsU4sGxWUwJqm1DoIckLQVnQsjCL4tpQq
8dgh7lShXtWHhM6emlAVz7R6pePIjrRm/7dCnwi4G564hAKUgzWOOagtpPs7aD2J
QaXMwwDY2LA9TcIHq35DfO2BkwZ2Yv0Hh6P0tawM/rvd7gW1Q0xMXaUS3oHUS+dw
`protect END_PROTECTED
