`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DRvOb6lcFux7yPML7PoZ5xgogglYsXPWlo3e6mABPdTVs5X/uurMukraZ5KgrxRP
sqCyhCydGjN2KLuI6kGTlUQ3AsiM3xI9UXFibmdK7MdsEvS93YwMip2YublQVLJu
gTh8A/CP6WeAVCyPkA4AnRzxlXMnVEqnZheQpiAdDWjZ9OvRFv4WK5a9FISjykjE
cFlJJF6LTNiH+83BTdFVS5ikt7afg/WFh38mFOnhXPxTiUYz6NoVxU0R28swIbGl
oUkJIcHVSDcJpZLgseuwLHZn9g84ZkuQh1kEqwa1N/UxnoJRECX13lMfYnFeZR5f
FWTtdFfk9ezKbmaglgpWUpxAmjcoEwIu4pdZwOtP1nRVnIfjXXrMsSyiKeW75HYi
V9Exwwzjbjk8i0bwt2jFKBSQKY2ei+KEZ892qoiLpSn41wgbtk55F6FQWhjbrs+I
ctOmp7eayqoyo6FD9GVPxWjmwIyJcBn3t1zycTJuZhSaG+yTNGChYOQwrPxAmsPf
v2Ea4mbw6ZHZ5h2SZ0EiB/NBm2RRE/SzAC4bEVeLTSlVDm0tYyYsA/A+q/xgYgUD
9ku512Jvq4FayvwSOahGNIEDVz1AOW4Rj5WPZpKpLX6auM6tFfWML6cUZNN95y3r
FKcNJufTOBDSU9ltDNi9QLjBaJGu0yZ41WHR6YOifUNZ+d6nc7c+IxSCzXeS64rZ
KkW43TrvbQW+c5gPNyajO/vBMMtW1c+d6OX3pgBJ8LNZFWUpGdEwkosyVrmya4iB
qnFMdeDKpP3AESfE2INkU8jy6YlfkesZd6iTy78ZKmO+JATUevFs/XkP3QSrbO1f
7sBh2UiOAChq2uRLCKpLe9hLHpl/thpykSsuB0uxgybXBTjsIOmzj7T/9lzW8j0r
tTvCFCrP4RrlQu+FmLPW1r/bF+3p6RVF0tWr+q43x/L0a6tEKdPPPU2nr7VlsGGG
C6PyvVGlLIXI3RhOvbUmBmlDm2mZADl7kF0uUa071AgJe3QDcj26khuAQrDUaqHW
zc1YZcyymVJ+Bv3wENqVyjy87h1oP/cPHZ+V9T541pvAG9gl6kb8xHcCgSGpyplk
jVd9sEht36lqwuFq2NZSSQEhdRU58NRJHSVKVw/ZX4TwMwyKeWTJvk+xEZYInXPC
RLZmSfGSkQJTKZL8SyP5p8JDR+q8XsGzALxnNcNJ4oAxFCAJQ+52Ohhn0QHmdGu9
UPM4RwaljcpvOA3k9EG34WNKzJ7vAUzSxhma88TN5I6I8gDbGEnCM9CQlgQc2+dY
E4g/nXI8r1sB3jHuZ5nGczr6uVzGHSbQpZfPiTfx1sa1gJYGOKNw0UAtsr2l6kSi
lBb52pQn2WtzdyJ0cx38+OV8018wJcqBVGmbOV1b/MhmORBZkRu5PygTaHXVI3zS
j/ujXoq6GP5dxTuRixErbOlFeDK0k0MP1hRVu01E6vWkq3lovMv7SPDs0P1rC5nr
j3x3pKmU6rqsMWLbxX+ko9fnUMNhB19oXjNEEiIhhcKGS2MXSK61XJn5xcjqKGPE
xhqQo4xNP6pl0mPGQWRsvqXki9ZUx/2na00J4Ft1sAhZf02DzODTT4b8H1Adl/Xc
FmFtwyuT/OR98m9hIRd6xDJnHMTNXjEGAjKYWhnWDT6MC0U1HP4mTd87mSAXmS/+
vzqstTF9IsO8RZrwMR/kkOIQTdxpT8DKh/0n+j3UQ/OilPXO3b8ZZu9EQShNEgWU
OsQypf+wxJc1gI/F4XmCQqf1IC8Ox7B91T1wCK+qeMVT5kgpIeuXXoC4eaWpBFVz
Wn5FxgJroRJRvUepRo97KNDFSvKuKXnVrkh8FN9xWVqLzb4xbTfmhKg8TmQtVwgB
xKddmJL2NRIzX/4QeK1xgyDNi/rbj1ZBfnkXw3NKdQTzGcVvaZa1Tx0RjwAdhjJ2
vkdtUM0fJXT+3zOyXetIQHcuRbme3bjydGNeJ7fPUtl62MECkYDG2mKpNCnEoQ3N
cdfQ5jEF9ixyzYOOIC837FlFdJus766PS7DOxr52TIpHp5WkKL3pRYcJeBE16n9f
Z2W87gJtV2DXLA/KE+uJzSrb1Hn3hJpUheC33zE6l3IN4i8h/Q2YHRxRMpmxjjOX
uFjlwrj967Ounut/+haH0AHAiJ9qNZGr0BikTnP5UDYULYmJCoUh3pZtbemNw6ae
iVBo2e7NUKe7YKkjnDx5srQtDMir9RXyp8Kjkhg1TvQN4RSKyYw+C7uINdhK/mEt
njibs9iptUATpS3sqL70cNBtDlBEgunVrbew+baxQEf1Cu+GYwcKpcuNyQM80z7F
EZIfunl9tNvm3EeLVgt/iVY8taXJhQMHyoCCB0tx5il+T9AbjRDdY2zEHgU9zbLi
+x6oozBxCj5lBXfk7+tPZ04xlypjLPnXsAmUUZOJ7oO4oOxCmAGtERrRwI119wrl
0LBH0kBPL1vu7uU1WxQVg13x9RIMWStFDFAnT63n7di7lDfIm4cMsh8ee3OxrJ1I
jmVvMZMkYXwoxWROrr57e+E0/h/uZ8tNv9k0tuiKCcMuMMc6PV+PeUrx5bj1Fi4V
V7mM7YWCEk45vMdkgovZfgJ4VH/U1TUhoTBHAx1V0ZX1GuX/L41IOJ5S5Oqk1fVK
FC765VVbWv3wEJEG/gDXGWRetCjEJtCmQKKaTCXqSHKgAdVE8Cga9t5eFfsrjfce
IoCT0V1TOgl9O0iGYeHgMEIpWUO9Hfxl/ZslbCnIGl5tIX4qsZF88qBIvpHNIzDE
GtyDNVrBRXZv5N2sSrIqSeoVOTrf20K0wtp+jiOLj1z9pz+Mddtb5sLbPdk/2eos
avtolgzI8oy4cd3q2i7njyaKqIPtsXSRMrDKsIABhxjiRrxzdlsrBcZGsmjZE4ec
QvjbEnCiH06hXiXjZSiOvRiOC/0RCBoT7eAAi4Wv5zpnItVyj6d08CuHZdnhXtlf
B/7kMwDKnlklt0zE3VQekxyQ0xpwGG0OvhqmoYkM6gnuqCxdtYWQma3PYgfo3a+m
wU1YtxWr2UqZbSCNPFkr+OC24dnnDQXEo2nrmU0Q0JcVhMdcuOgPrYy8QYQCHTX2
gF4VbRja7A5Rq+nPMYotcwOs3/T1FNZsU6bbNgFntBYbdN/WKBwRr9TOlHCAvyce
5mHhrbyzOMXtpH+RGXTs/wWztQ06376wX9FQNrg1OUfmyHC43dcL4Fk1NJ8wIpmZ
xOO27QMM0nKLsRemlD1fVLpkNLp0xO2HEvClTPQNRHOFr+xxOUkAFJb96VGzpOYc
WK4zC6tNmlp0plsOSCgzjulFg9aIbdgyNuxIraNLEct/Q9aPsF6Tv3OzDruCaoVI
IkO9ZyEjcu3B9QkPxnETlMcps005uhJmZ6dTcruTxz/7EfF0SLqdLWBOXM6P3NKl
vOCY0ui8Ar3e5KPJ7MctJSM/g/R1uld8Pp7JuaXf56poeS/W/O2Mdy+WfSXMOmUn
`protect END_PROTECTED
