`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rSkodZCbTX9NoOne955kkpXEmzB77Ul5w0C9sKMux3xDtaAdY4jbUNvHJwzFActj
L/uVFlNFGyzLz6MDIBPnpUCbTMkPWijomL7ZA852wZjdqZdX9xCg2CmVW0cu4yru
TtgeAuK9H15jXBIgxxNMiUzKbT24d0btMguJ0aESUIywmZC8SF9P1uMb74/OHV4/
SC8azaXPdA0KsIIRWoZfEHt9wdCGm4DCJa2lY5Nf7zjhpNgrMlR4zueYKWj+efTm
ROnEBTt4y4+R41qrUVqofMj7FQL+PL4gyoF4vz5tt+j1tV1xJeorAXUucnKtY0Rm
jrGEHy5X0r3XupnydTFbJEp4DXa2OqmIn1YxRWQZ+pT8n6gbeUSNU4sHdT9+rzN8
yzQL6YEWQfGbl6YOSsDgNE3yi+0Uce6hViKTVZ0R31ix8QycjZ3MZr8QRtr6b0tz
AHW4x8pAwaEZKLtl3PQtNUNrOx1AGrhEaBha5dy8DgmDJ3l0i/iDywOVkvG6caHG
ni7jA/KbQ4U+M5XvOcxyaOY0HjPL1SbdF7pBTygIuVBov/DSOHm7wDRqfctEzJg+
qe8+J/TZwaMdLDoojskpjCOees1C9ArAO3Egm8zuODGtdprnjuhRSCskEZ9dvT6X
3LQkViOL7FSfz9rrTBYEak8dycflTLLMdBFHVYI5uGy2cfaFOePKImRjBia1Mc78
Sl0SRReSaTETcZ+EcKtzGzkXcGSd/1v3sKgab75BdMy8mjs1XwWUrQ9FkO1naJ+u
rTl9Qasiij1RAefT/b6J3OWABjDz6c8qr7lzp3pnTAkx4/JNTEwqwCQCSZNr3+g9
XK2MuH6pzZt3oRUEIvLsH00kxjz2jkmQcaFuU3jLjgigSiw2VT498tkGBrljY3KK
rn2QL45eO84EfT5ZAXnlzMuPFygV7gIdjj/mIA47/ag8IGsOH/op9III3gRACmv5
dTx6sJBpJkE+nSV42u/y1wT8AQ/TRzr2oFvdZqp81WrTsLZxiPMH2uNxvSLdR9A7
5dyVKFs0ubQHmqfVtD8S9Me+1qR0DDULMf4zZRds9mJa+b3vIVVTESJ3KUaF72Rx
C6dO84Ja6SAmsW81SnmUX5ZrbPVJx4hCZsC6TB78tCxmpOKtkwzlLjTbM8mbf1ph
TQ4YDfTJj308iFiCX9tJMu1x5cumgh3VnQdFhyTSmCf1GWkw1B/LWqRHl/yBubYC
MwA+YQb6X0k/kErTIJuoJmwSIoU9AWXjsy3bZ+lc73XXPrLc3S8A8IU1vuejmwBY
6dBiGG9I8u93h75IHf0wssCAGAg3TVSOiYU+RkG66kLZ6AiTvR6sSDBdElqwTE+q
gHnL0/8ralViFnMnCbXpbyvL9RMcWOm+lKWBhEORJG1cUuPB/kWAUNUhofm3Vc2l
LSZzUvWb50pwvloEe8nTGXL7RKGoO8EhRGWFqxuBOpPHrq2KJjlqIdzVNDA9o0Be
91WX8OW6FDmogAnfcc9dyRYvzfAlkq6XK641dluHnWURp2db+MTAcaOFpRZrvaMJ
+hKTAqegP94bcjIdfQxcXm7Qz/CMxjeewkc5tZGmG49//EGLkhTQB5hMTgmLLq9P
qFytgPzyp3bT5nlnW7s2e08JPljOunEqUHarli5jq5NpCkEGWm0B3IdRBQjUWaP4
rRqA6ckC30i07BM5/QFNN+4tmWd0Xyu82kMsHwvWgnQCT2Fv0TJMZ3yxRwlgv5JY
BiCG7RCHpTsRSYLTa9P5ahfIgl4YlPtaB5g7dOq38zG9r7wAbIEhdqJ5Q2PBe8Qy
2BO0cRgeRcPbLSli+Vyg39dXofXDI+/5kZy6lwzkF52gfpdMcTpeWOsRSjXS6nDt
MZLvdvCVGBJfd0uxlK4je1Cs/PA1tFncy1Z4suYm1GtfDpgsfqPMQUCsbTervkVB
56XIVigQTJnKGhLfMwH8dSdg7/Pm2m6P36d74RcK1ts=
`protect END_PROTECTED
