`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m7ibzEo4O0qKFOURbY8KJ8kO1g3iUKMM+vVczIXuq8iM9goQQ4cMhN72GlzJ3Es4
ntgvIPAx0PnT4C6FtmKkIjdE6pou60nAIijKHIw7MYkklaVKd8shuj9OWD4yWacd
s5JOFiBGOdDSrsk+JaNpRUbmEO4kECPLvVxnkBSh8s6vvDGTVZweHTBEAaXQ3k8L
TUEQgKlec7Vl8vFQk4oJuM0Vy8dXRb76L+DPXQqr5x7MAtq0+HLVvPjOCVq8iEYP
7vt4PZ5XSfPefX6z+kYW2kHKXBtkYuZXEyNMj7jTxTEegXz6V7Roti7x3tLhPIHU
dz3baLA1JCY7erzmOWhX/uEn2HbpzXDXaBFl7GUPcqtYglSuVQ0mePmngqvwZng0
IK4YnKq1+n/tJTpJ/s/xZqStALCYfX48BFFsrmYfe11nA4BEhWhsTDmBlXTD68V7
Vx5bFnIzMSsd3f5n6LgnN3HIh0OOebndnMCzyZ3mT83MwkOat+1MHmTeT8XVpcvP
JG4WRwgAmoxuGZ/qPgsOcxHXXp6oBcvw66H5vPKJD0zuzcygi/iAglgKgx/zapYu
94BOVOatgzEl5d+EN2fkMLjHwn9pA4IAfLSombTdgJGBSbl6F/liPUmH7Bpeq6eM
H1fT18Fl8HPopERmfpLn9zL0I0CPTb1XlQsORCePiPABSkrqL7I4bJEHEHo6x+4d
XBDlS6ffcrpauzlOW/KG6WBmGTOkuuDnQfqrXqgeWUY/Kc0aHmgVwnkUihtcwHRD
Fv4md2a1B2BWQVPBI+MVi8+y56GXKrlPKXmv198yaigoUEjUfR+nx9EKWmp0jilP
0nDIMCsP9GMJFq8143bhLYC0DBOGe3V+2nsNEa+q9kvZZTq6R4HGgMHgNH+1S3lM
Rk4o60OA1I3qPKFdv6jNGsJVUwHQEzxKGcYm4CNCECEcDiidiRRCMT9eGMoDFIjg
Ig4V5NULfsbPNCYWj+gG8oyGgteJzSrK111DwdusIYyIOEZckt9ko8/ckZh9D1lF
p1q0rJfkFoHjONbXRhpMkaHxWBhRhNgKAryR6YeJKSyft4/oQK6nOvkvtYQJyQfO
3A2j0CTphw/PGoaR33YdSSYWLMBP8GnuZyFHCmsnmQ0bdfPtu5Ok27t048tAyLXu
AjXpDBNZ/QSaeH+VorIDYbPLFSPpjY/QD6zwCzhr2WBthd8cnTbmz5gQDAJomaEC
SW/sRGxaXyPqNqkgvLuj52zYIBNO79+TwzEzhp6FjgK0VfZl2kDCtuWBD+Myvzac
dpubLn0KXWYG4fkJnrMPzbQtFzBj5q0TmgC4hZBN21VIe2BqJ0fwxR1m0nG+n2PF
OvrBB5IeN1MW9HjAsIWS9GMeqScOrE4r58DibFZv/cIUT1nxvRBtAEItLmwzQluM
yOWxLDVbt5/BDLG7jtpWcXH/jwvMSgp305Wkjf6DBLufXrO5DBpM25oTZlgc+lwa
hnskhl3Q0f3pJ47wpiQXBP/w9EIi41h/54+D6TqO7tN3QjTej1LQTKdQGH/rih40
kenzfejhcLuOy8kOuoJnCloXjj2sDhxtOURJykd6ezn8pzxnosaWROoqT50tmhXL
vD1/XedUG3GHG5Ij+wyM+B1r3yIORCTQywFUkSrhyl96PZ/3YOCFfY6q7XHvfHml
E8REZeI8/vCwBLjVtTFOnvA6mWGCuWzNId75pz6Y5FLEU6Q+VVN9rRG2qCsXJfEe
3OhPDSYVoQnGL7tduSfL9IjCpWNo6Umss7pY+gUPR34j0F5559jcxYPdbGxw3e8A
Y+CGUgXI5lqc5PXg4v+n4zPjGt5y2mrzcbGOhUPRUHP9BUnwfnIgyqPBSI6pBjv1
YsyytANJX3eQZQEwe80oP5wCYucZvLrdTdUu1yTUewxcF5+sJmNGZLRHxkjaK99D
Bs8yUrcyq2ZzZ7m/WW2AkMMRT+KKfCKVy4FixRVPEd82iWeEnTEWvo0AwACneDR5
ur123aJJVq+HDNerXP6IkwUVkPlr1CV6n5OGwNu6QvGJhO6nP2aWrl5pLTneXhp2
t9aLi2WRJckizq9r4P3hRzEn4KVlZFf8/sxe1n4LT3ghis7B1fxgiuxnuiFtVAqn
jyoqRq/HXmaovoKEeq2h50wFMANpy16HldqoxUXftcA7cS8sUBa3Xh14tqhZDP4M
mgYt7TaNZLU20DnUlqGj8n5M+9HRC/M3Gr6AXKzZ2RFZTa5lSx/tqXSJqTFHnFQd
s+eidiImuN5d0ShI6gLCWek4yj6paWrp926/oON16Er6wAyHbskb2nrAMx8FeXou
zmM1N7/PFC/jQWUHJRgLFtY2YwZafOmC79pWoQLdE1qclqZbLddml/XO+ogCllwd
Mb3eujtUwSBZE359FJCVWGyjLi0Qqcn/NkQILSnCfjxDg93M/T8K7EDpuxHBdAJm
bXckBTlZ7bJ8l+g9ztR0FlM70R+9SBL0hg1LGxXugK1hPvq2Rm8W5YAiXi2430Sl
DMub+PBhjq4Rkhl1U1/v9vFtpFotWHC4S9nlgRhOO1GZym1huiF2fWVJnG0j7CPr
6bWoCvZb2I7qHC0XGIdP1xK1c+TIvAl2YG7mAGycea68EH2zFcEGg80mrrodaciC
5CMjGECySJwwZCvQAMKaReztd0oy3EzIuJn4ozmim0oWXigfpUuUPy58KLfOoV/A
x/mSqE6XO9tozwJbABz8xTE4Pbbv1r1Qcn5gESEd4mjcu5oR9Gw5LIPHye4kUG9o
/ziW3wfxsY4kWKBiRpClNiiUwgzjn1xoHDmD06Nzgx/QzWLHznWATs3StDxifFZT
oZxQeTxkGsEol6kIh8aVZlJvwGg0v/Le7bnsiyAkC4gZZrIv3nAg3rgyOqCy/N4Y
OTYsHCW5O3GNjSbBFM+GmSOzCgFo7mf0IzZtlmAxZ3rhZha5xp1Aditz/TJOSwMu
y56nwT4j5Y8daMdyKvz0FufidCmcKoppV3DQXXiPIwcASCuoA6mBG20/YwBlzx4L
reRRm6DobluH958yE4HDkjdbQAoias430f7/buJ9ANv5jkSMS9DdSJTfikJRNv+N
RMUvMlKDIAqMg3vY3WBAWDXqdG+UY74BYzFuoN0is+VLAr5IzkHM8CChE6e4R6pe
42nGYdJFFToMmBcp9knhnsqkXWhJNdnmPEe7UJZaTEsRnGG5AQk0yXjVRv7Em8xt
zo/BlzNZYWXs7N+I6GdNP3LC/WKKn7vlJsTBu3XgAbORzXOR+EuU/E5Gulf5Z6w+
eFUSPruzNkKfhA8pp4dzP/ERc8RsUsOfcZNF/mE10kwJ4vLaP2sejP1jke42BE2B
bLHyRMPeKn3pmEoFpP3TCyy4yqARDG01MWMRSrgNnm3fpN+Pqvbo9hMyu37V0lm+
3Ozs/GK0b7frtUfBzX7Rh9FCo3jHSNRtxLEdihvsV953S+LOXA5D4J9wCaTeMoGo
XrWcI3Nxdc5nJeTpk/TVkcws/l9FJh9o8C5MGkAbSN9jzGbR2m9eQsHBeDut5zMP
FOmts+eHlpCd1dn1YPdkJ3/lfcuY/XvWefKTe1Vm5h1EvljjrXINKW9NWKBrDz5j
9ZIaaZMLpWQgFlU8bJlc8n/9A6AlLklTtfaoKoc8MBrPTPol8Xg3/2G4q8OTUBcQ
pJ0D4Zswsv62I72Tc3kALPvZNF4+7me0moKAOLPmrKBCw3U4Ae9T/QCMCfvnEbw7
czzBaJrwWzwknGCxhGnee9AZxSRSA9Qa1C9luQ+zBqhOtGAZiH36GvgpTB8iz4ky
QG8S8vbMrcetpetb3Qgb7vcszJAcQlHaD2ZQ6itGu9C6tQLsRf5A0zL4Q892BT4O
kzmrLTeMCJvj7TEwKLJ3aYogzn8oKFIs7pnQ/MSpnlR0y9YsfJq1+F/BsHgnlUc9
4G3nQ4AinWNIGnks36jaq76WX9EIgvL9v3fCIz8c52j6f35t59T9VlVaL0fQL66s
Hm/44wdxa1cWGadBT/walUqWYkxzAWHVhHEYgbCqTcr698TzFa1ne59Oe31yx3Qk
eiEDRyqURj8kJKCCW8SejXMR92MRTNdc9MojSa3g3aQPSsPW2PPEHDo7yeQwtwWr
iWqd+ZskW+GNbin7hP1EQbk4bi/HtaAnTtV5wPH4kmZbVypu7Tk9o7xrJTZuf3zG
Faj0H1PAT0gIO5RqAhpj8G7hpMXR4GsdWYYzy5jOO7cWFJrC6GdwAlYYePkH4swF
hZPjI8VKirQIOobndElark4NrBjyEFaFvyVIKysPitC3o9To2kJttYhJHF1pHjMR
4jxL+72ftcKOP2fYxGVR/Gl07AclatkGW1+ywHTgkOk+MDeUPS/ZhqAdpBY8znG8
EsxdHoroLi0QesM/vB+6e+s3SjZVKFaSHdYHLk9LC5OLrEt2wtYxGptHal9tl+td
XmG75dcG6U/YGXQ8W293UP13eM+Am2KerOBlmlgGFxQGuQRIPvEIgs75nuc1ILGy
X2F1+x+Ogm8yLhxv8T10GFo7EUTEw5i1PDVl4MSy8/4onHlKXipMBTZ46WVkn1mj
+G6sjZZYlHM4NrEW9ACpPcqooKxiorXyHSe9rHRblaWWko+7ktykXQACCSgVfkma
ttuHAiB5Mk3kig4HUXhid/hhJaGf+5moD2YR1BQcf6Vz4MLMxPJWfcsJN/66rtTW
OcyNfbhXdi8z9Hfba30azaCByE3G1CB7o5ObtogTDec+ZwzAl6TeXN6YCfA8w02v
1AceAAgGT1qhmA65lRoKskYCRlkyDuhqyQkXismBZnpRn/wjSkYrDIh6hMaQsYFM
rHTnd+o9kZtbNLPPHNHs9pOHaMw0VOgNQ+AqvE+SkREr8bj0RHHKXS3xDqoMc/ik
jx3/Nj+iRyDFKeduKSAnweUQQM7dTXsMd7SKh/9P9woS02JDubhouLHK7zsEXavv
Ah4TnW14VVGBUs0UOZehLlDD2x1vrhfilCyH1qPftw3KmgtO8CVYeMyEMp9+0Hyt
tv/X4b/6KGvFGqX59gn2l+QDlPafnfYGhEhAru5C30sYqKr8QcSTcZrzbs3B+yyD
HAqFigKrJT3T5GeiwTNT+B/Tlgyhe0fn/3ZCneBnnsgw6OzcqLCeTHwlvyjf19YZ
eY744OpFAFwpUUdau9DLZaqNskFIgGsIoUxnO0OIYNmfQOxdJocP0NXMTn5WGKfC
pplc0DM0Q01xN/Md/9HTZOH/qpyy3EjlTkhYBcGynWpG12gHmeu/Fmj9VTkglHhU
3ww2dLPzl3NtjWQ6H81WG2wNojCVDZBEx/Ukq2eSuUtJ/DrYeIsMkru/h22pqGra
ZZnclDP2BUX5YJTwD7Pgbxw9VCNOsTJDc7tu4MJderP9SOBPclQe/Q6uYLYsC3iN
xk65++8ZFEPooLAu/JyZmV/XlPz1I6YAOJll6wiEfBYupXWVB81Rpg+fBMcMlHoO
0QomiUbicyehAlSXyM/huJBLmlRhswYJ5tdo2FUJIeljxt+WS+/3kl2FPH9v7PMa
qWdisVQEXfdPKk7NtOrTiaih0fawNIE8BcFcjg9EIb87Ba8UOPBdR/spthUKtSmw
vK0s6SRxzmtKXIc3rikSqAr8KyVhOJQdfkLSrHHTDkw=
`protect END_PROTECTED
