`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FdYU+T+Z9Ugrevi11RgysIDkCcXsgyafD2jkfMtJ8jHZYZgp9qifodTX+NGLedEf
ZVUZzax145NSittb0pqeY7IDEvAm0+DW7GbwA2SGi9sed21UyLCVM1NVkEGN35Cw
qC7f3L15TJwlv7zfLHifFu6WOgXJ5IsnpSNb82RTuG+0cg6++8vbjrOr/gfu5NQS
JUBzXXx286WUlUkTXqnE1s9GAd3g+d6WiLnhyjJCRX+e8x3HmKMvK6IWgQiL79O9
j5MXwUKVdhUCy9FRgGhCbtEd/CXEslZDlHd8jmKSOcwHoovMIouey6e66SoKFELj
8hoNnFLOPK/XnHnydlMcUyVYcLAHu5H5C6NWbS9X38Tj/U9bp0o7BkRcOVyhqfdP
nFKPmsxMxuZ1FxFQjLgbwuwzQUGKbyUseR8vvBTprnUStuef3LFCPPPGRU6wqVag
SmbXFls0CRcUXBNpiptjQtHg/87Dvl8AQDFy/ZrvJyXAMZ/lKosA88CtHB8XHg/5
YG7n55xmBhXjcG2mbQMQhvQMdbnfDSLvH0QL9cD1jqe1/voL2CQE5XrzR2o3a8iT
VSdQ734FHdHnEP1z13LIMuzUgzRAv6AqrwcdblnubYUDIj/Fb3wku2reKANnYzeo
+mFOAYTYk9ejbJTA9Koj4H5xibBAFEUVQhvXUAEUyG9b/nDWEgoDKfi4J21A2woj
vPIDnEgN7/BEF82wxAyPO6Fx/wUh8KdQpiQmF1nl43ceCN2xlvVjzV2mPSsmtgiF
qOHKMtbagJPyhKjfM2JhjxJWuR9tXD6Ai3awYjFQ/1CXoP84UV8eeoQk1B2j2kZC
fiBYuHRWphXFUSdpnsFW3yQHqHPLq48vJQ+1Dmi4y0INzOAlJ547ZNrmNKwwlshg
xOoRZVJd00txlHF8o39vLxOVpOehl2LyhRgj6mmssuDD0TwZ08svP3ARzhlXB2Bv
qS02lR0GGZU6RgO6WLcxBf4JLw8qwhCNBCrdC+1zTU6MAuF4WzFzlVpm0S3SFSAg
yNaoxc3lGsloot0RhIoO5W/TL/q0O4Fo3GLMWic8E4Fx73mYWEy+RApOWCgvTPZo
B95/h3tAdkSA6PJeYundbwIDShOwrd1NYaX63LS+fZGma1pf4sZjHXGVcC56A0Qq
mfFVoJox+qiGysUvnzk24aNMeMNJaLISPFnK8Gncx6ht2QpV3vodcX7mfT1vK/uP
xIL0pAhnAJW7kFGE1wKWxXNzoa263ulhU1JMcF7inqxnfeK84/AYlyj3Ncu3TA+m
oqsSJ9sKZXMUSDdxzuG3P/4mEPbEEo+7uV+41iZ2T1B772QXxKu3bgv2GtaXy+UJ
gerhfqgHSyFNKRN0U6jq8I2BCloqFjcDBphcy6nIBSDGFEOpau7vuFiTLpxTbmq0
PkCx8vW/QcwtlXXK0+wCkGoldBJCF71Zmrf2RJp5Hfxea8DmZ96pKBpSpNKWc0T0
vjgZLeTXXOy/Ob5aTg4k2IU3vCzdSJJpGro0Qq19J/yLuMYtamyYG9uygVeXF7aO
PpNNuC0HVFSb4d4VvhCq/LWNNLT9rm0LwG0Pl6td9cbKAclXyYvC8YX8/fsMnKwO
nLeYLTstGbUW2JcfFOQH1ViskKz1qJe6/30ml370s6Ms3xQY2K5xO84xO6iCiJtY
s7smI8VU0dxEdGM7xJqKbJJYCy0rhg9+KrS9w0JcbRYYmJeXR4WSPAJY4Ui5ml9N
vnCkv33Smo3bhAfheqhE4UbcTO6RTeuSbncGwO6XpTxMZeJGPVYMTPVUdTZP3d2v
KVYjGNNcL/UsYb+JDMW27n2gSEJiHHUHYOx4A6xOTvjBrHGpmgFOx5aS04aRxsVZ
lZhCXsdOC4hjRBp75lP47IW6Xvp2DvecupmQ9ydyAOI2VQe6gmey16gk+/saPdFE
xfgUddqBWfl3zO793Xh0A9abc5KPtmgi6K1LkyNwv08Ndw0d5ttJ89CXs9JzODtL
TdqtPEarqA62kvkSB5IgA2ylJr3XgBrzxq1oTisz4MgLNkkF1aYm9g/YjcR6o+UQ
kW2FMVynXjUnyzzxT5AH/3gO6IldtIyibjtSFaeIQthfUiUaE8D9q7SjSsGrnRNi
kfmn1Ldflco5HiTP6wJoWj3tcVOoiiThczH02Tgd+aTbDEK+MmdKnSB/EJb67rQW
p1IR+aIEb0J5LaSZN9edhkwhaYUL0kcYQVRHYj1yJItl3v10Wvk9j6BJjhAIjC6B
ux6wI4naCsi5cQ3T22AfXaV+V6VQNe9/Nzmi6fHCRq+Y0jLuSI0vExXcYFyO+sSb
7/EnvbP89PGy9H823qV8QcmPxfHDZm8X7uyFY6lFMsblgvY5vzRmeC70nNsFUtoP
2J33x8i15NC5mTwbRCWfKi7o4he8267vGv4JLzccoaS7ykrcbv7amxLXqwLDBfsV
FN+AHpr4/igPih7PXETosaVXPN+Q4X6+4ErmUYekYAAqKpR8o5NpQLFsAIlR0Atw
q3Zm0waz4zEa5CJPhkAhl73HAg/4nT2bVhPLjG5cSAlWziPLugQSdNtGhx+UmvUf
LIlh5XOGmReq+yMDZckVfUJRpv7Dvtve7C3KzrhaDofJ9b9jO2JUfhe8vpWiYn37
XPGBVrN1oApZd0EjeBNmcD2+XCLE3BoUEyTEaFODo0pvG9ys52iAi5dRR9186HZR
4OYy0wJjcKgKhLuSv+IxWyTBPLhKJjhBEqIUs5zO1r55g0XJsizYait+gv98i2ZK
HagqIS4iilSFmcY8x3aCe7rAvTWBDHk2b9Q1L7ne/31h1crNg129RdKSXZAuqfSy
T6DEqZW0iHbHzeuVcZl24zEhcwcOKOVAtEEtHWS8U1yM9IndCM3VQH5DWo4KCa3h
cq9lBII93Ms2DyP9X5R4wHHu5U4pzdEsypC8R+VJKsU4LdWci90ZGhYlncx+UiCC
zEZftTj8gYStDixfL6/Y2lxgfkzfGGgFNWx5+HRiO6+ZjLEi+G7bmbUXka4J4++r
2ezKj+ac01q/8Lrs1ilLsjkfBxl3gDJLQabrCNaJdhFsshAA0uZrlOvZYvr5sdGZ
ADe9yL18JcGf2kjaFvMCi5JOkYfoHmhb6UVK5DUdIdSv0drxW7DKl2waoGbZV+DZ
kP2fma4djKozA2HAYQqBuJgv4x8puyr/YObSMfNmQT+dDi+B0ugTgiHrKyrpurWe
3P6Ewz6gA1fu++l8CLPO80SLe7cO5chU0WZiCOm+BPmd/+68iiwwrFg6IjgB143D
Ks9Ja0yomTmyqvL4LxnTQBJT8v5Dp6/dLcCYr1ZwuCEIQYxqcMVkbCZ1TJD2whJn
PsGOAwm6W/BqjbamxKeQBitqsovIKFALSfJOs6JtoZVdD59Dp4EsoPVSfnct1PGN
wvRpjzN6k6NL+UPxWFqq98ER8jQStBf3s/FXrwSk1wQ=
`protect END_PROTECTED
