`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
76eg4hNcR0T+W16JvByUnbpVeZ+erK0+wtvMeoMBy01bQnRfTQUKm9QikR3WAG/T
vzSp5Xmemf2hAssHKbyZ0227bDHuFgNEV3aR4NW5mj6VZTzpR6MmzQxn+Vt1DNXH
ldu4Y8jedw4MHT1q5RJ8xK5CoDt8ZZzftWUSXgGU3ExMrXgJNvDyFcgXtkvI3j9Y
AiBbYi4dUBqvFUGVLiLno/K4DF4JfKPIlLafNqLUpkbV4CjrgBSg5FNpMsm8DABS
ilTOXiz4aUynnvFbTW7OdS2OWHN2750osqpJ2HtvFer7JO0kZRpCRu9Vzf0mH19m
8oFBiMXDZsxLIbTM8qmoO6HrSrJvApHUcaNaM9rTYTZI+diarq8RWXb2QazcNj0v
ro4j75b5QvE6wGH7isCoNhPMPRT9EztpBPB+Qn0DQDLjBaYVyNNAi3NOTvFDJLCp
EL5z0WdcqYBYG7go48H0GBQfswCLCxn9+DZobXijBuNHJDYz1LNgGGq90/2Bq7FD
sojdFIGXAP7d5jULi5c1MyaTDY1TAJ/+wgqA1n3pBzytmxVzSYt2qZfA/dIjJ1dc
mBIqXlXteMtdVrGBLNr1EegIunGFSZsB9ONaRZ61Rk+LFR0Dpp78waMRUnczpo/O
DIfWSLnynyWXIUCE5r/9E/aimohZYkZrmLeZMFofRxkRvsK5e9fnqLChS3qpjcAk
ZE/PRK9v1zkqxzWdPJF4TITT+VhJ+3JUn4Or6GEWm9zSxXlojxrWZDU94yriCPnF
TZn84f99U3vs3itjgF/NNQMt9NbsxWnnfnXGPjkMxDrR+H4iESj/idyNNR12LKCL
ymhEfxBWnJcc7JWEGopenz+9hLFpswFWF+nPvKTpZ2fhIBSWxUo7c5YhSbJjm/JZ
Qjassn/qbPaCCDbx9QMKJDkT7mh9TWvLX+iF5MGBsmW+7twMSMS7Hdff2nV489DD
/LgjpppcGWgg+EFkOctTooJkZD/AVFjRj/qan8/2SSrlCOnu0Eg8kOG0f57DVAij
FlmFriKpc0ARYb4qmBQFst02FuAVfzz2KU6EuOQCA3akZ9psikPL9cqrCGFM1sXV
Wyjm2GpENccOnUxxrebK7g==
`protect END_PROTECTED
