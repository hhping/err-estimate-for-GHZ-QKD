`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
btURa0gni2ZuDQ9n+CrlFqGa8OIlCCXv6a0zO4PuqlV1RK5d9nU/qB7uK9b8cUhy
VqxCIKVL+9vzszmiA1quNd4mlKL/8+o1qMy/g8hFc3d2QegYfz0AzrOZ6nfp2vRx
u9KDTfPqduUDZvmAy2lt3F5poGA8TS8Qh4tsWVeKWgKdsuKzOjoZiF9+LXNPzULC
h7rPXQSXOOzxPEPfMuvSQCEcrIVgvZtez8aq+tMaydqJyiD4zCEGjyAl8o+WnCLF
LfkT90pHVXjKoON91XR9FvXb/IMCFI9cZ3tCppy4o8B7gNbRTMfv6F/0yf6odMw3
Xn8oe9xXzTw+0cAFpaE0Z0CChTNOtFCRNbVTX9g65OhIhratYUYiJ8vsqapNXvwk
lTwN7PGdmmf0VtIZAJQqEsmfj577kkAebY48T6XXn3GA7WqO5MgF7PSPMWeKQ/u6
AZEXEuxlMZTJFppR2y3O9+w+Uea6gRhVzagukjAvIuJqPpZk6A2uGGOGQSyX3nMv
wME+5QRY2FKegRi2NHBxwkB/s9dYAoUZUPc++gtcxn0Bui4P01PKaCCp8fw/Llsf
SuRLZTapYbM8HA64Zz7uufmUkGgKx7PvalqjTH722rSARCqEiARAGS27bkFeeGgz
MMFzfOG1rGBW5h6EihcCbkyJWwQaWsh76WSIMfmo4966T+lraIwUqLF21o4qyKc3
g1jcaFGZIG2QfG1EXbmpwsJCOV6xrdbO7OaAq/zyx90b0eJn2JK02b+cOrbLtRZj
eyhOmEFOMy+y246ZXWOUBhCETCL0ZAkr1YVb+NWNv/PtKKiq/FY+ixSYMaNUURLd
+6Ze4CQO5/Lz6BspD0rBk3eRNRTm1fvkAgnrWNvsB7fVN1rfPZV57RUZdmRTlSNJ
tL1Gm70v7gIvePcnjZXyWvNTMOkSm9M3pdNRyIeqQHabtfXL6p6/HCzsNSoN8TTS
VXRw35JDBT2tfsTa0/na+J55428V6BHCcdbEtn9R/y6aX91xuYDtm+NVBZQjFwgn
zjUWhEJ0jgubC7a+qr/iW1GjHYuGDxEZD8sYaMhSmG0OTKcHXZFi1aQ0oyYK8jn/
7290mXJvH1btVdQ4QzhUvur3ZOH8HO8gv0II+6hkddBC2uri261wSoel/rzqQL0+
2Fu3Qn8Fr+c4BVXc9s10lCBbVKrZPe+w8KE2Zf49Rel9vjvWT8Uv9e44vqGlWCrW
TSqaCGljCZZVdtO69VBUogBCzNWMGCoc2DUhAER3w8BGrn8nY59dJX6PodlzCqNg
dmgQFHhT9Mfg3Qgh/TzL5+a0lLPFajDsBr3YxN+M8REP8+l4I5JYMkS6U7Pl/52w
Zm2F5orzL4lpjkAYgUscYTbrVfO2YtsCBgjGdXTDX7brUHaSgRZj7g12SSxgv01x
K+89uDikn7kIatv/XZinmqqHOYOo8KxH3r2p3CchIFbZoeCJfhOyWRhjcwTKLYte
E9PsTkVuu+x9tHL3+MPfvr5CvgDsP/ZMhwxP1q0jUVGpK6UVd786TLUsPCOGP8lL
s02LSe5Vyf/jJF9L9e0iH0JJJgLY5bNi3gH+Rq2vKsYE7ROW153RDwcAAm802QJx
st8xT26ds4Pmql+MyCWxxVNvjXYvMwbpsY4tQUq4/rJmPDDCYXCjxYUnYqrO4z4O
jvULs0EtX9O3NL4SvVymc5uplO7lIE83BfStkIeuGJUGSP9g2g7QjTyEcFgJYrAE
t3wXbmiEQgNltpHs+1xCocViQMESpj4S1wq0zmRhJpsHdlKe2+EtNgw08phOkH/r
IUT1Yw5y1xQG+H6ZLVKvxzDvSdpwdY3seRboPDAn9vZ2uubnYCz/Jnetd/8NeC9u
bFKjmz9l0+kyZS5kbQqfZWXKq3dDL//XFdtmw27UMGkSrnmkkylkkIsEN0UG/9Kf
DIUkbxl/H1JfwywIqf/5i7Eei1ij5b2iC11r8xITwHDIxBhGjBdwyXfl8RXgNG4A
LKn8e973mjAGVg011+FFr3WKhZ0jZbEqpaTXqWD5uRWItuBPM+1rMZeYH51YjzOf
tM4a34p8+98CGgEp7OyAGo3aTE1ovh/Q03qPxlN9P6vdJXNFPPQqcf4p3AQyJQb7
i/50UHui2D2KZf4Bd2zg79VTX2qttocyrAlNnd/Avd4UkN6tXOkmkURVKDvDBein
lFJazijkB/kKu+bQuY4sw/JOUCVTkj35l4dYHeJUMObNHrzqlW5Oax2mgTpy7xbi
o440W5zteyJzlxpPi1BGxPEoeWrvgGdJGLFczmNk1v5depvqSQmJPHu3ZNnJFH1l
C11aIfSo0D8RZZKOgLFUCOUJOY2/OuvfN6xcrBUinUHMrzGWMEFeaK0bvzwDgWai
UQIvmS7meznocoMuenTzAd3tpDN6Fq9EzV7XS03vve9LrFrx1jkb7pz758TRlcBg
ZU4ls5+gx8ly0V44Ya12DqC6yLN5MZ2WXQ3rTNfSgRSUbna9pIjow3SLgU+TXPMv
dNaBh5y1xok74CU00/X96Y9jSzkuzaw232HV6iwfGTa/9h7Ck9qp4JXbGLnPOESm
iVGmaCSqN/HhVHHXUaX7Ji7lzKwMv/EV7sie/0jRF0Wt1HBVlqcLfBuUDmIAd86E
UlXQnUiuivCgRdJoulO/AgyNF2SRVwuasBiGa5mtidJHBq1IxDEo4cTwO7O9GrJ0
j0BTtzZdZJRG5NzbDGqFPMamkRTb6zMNNC578jduFUDJW7eFEmU5EbSFsxOs5Guq
yebRMPLhw2Fl8ecnA3r7UcTHAoreCYOvn3JBRqc84fgSrhrSgYhqUmUk5gYcZyii
sQvB61V5MTnBhCEMXQiQhcvaMUv9f4r9/Drg2k9ZGRrqUT5Ouyb7xb+Z1WTgLSLS
PTmQLfpvEMRpWOaLn6jTZXZAc1QXb9vhYtw68XzPPK64rVCJu96naju6bNcnB4bA
V0PrRvtdNrzVBb7fktbfX901fB1DYBWs4oMppf2bV4h3KWTEZDX4r5bC44H/DhOE
w8fVmNJ57Ketf8A3E2YmEjqpVCqOBVLH4+k2DKrhihpwdkNojtB/8ZVSuJQY8ql+
38RE8XxIXw5h2zcj/2/P9NEEd37EEwWNNf6P4WurwdJMWcixdoh52vMElk9zjD4V
p2Sz6l20hy9VKDeNdgVZ+H4UCRfR3RCOzHAfwznkq+LHhQNGCX6xQyVrFdVkjrnv
ojXqQ3TRorY247g35lZL3cUtSi+j+8WyzRjNcWNjkTQq6S0aJwkPZajW1T/EAX2k
DdVcQhqSvZaIYhhxtQ5Lwo2tiBAUFZ3k7OV97/smpN1jwT4KbC7sjsdfnLiG384x
POIPXxXgJscyiinxT8OM4y5FDHwGEBySRQdtG2sfMsXjcvib4tbb7mSwmbDxCk54
amJmdptsFTJVd0jWqOdvf/OzVSYgkN8zUMHCgmJC+9/LsuH3amNFnQnFFyNDJWRa
yOAKVu0GlHZ51kV4GsIRoqCLTyvpg3K7kpZ/+ZjqnPysMk6onoKB62ZXFa76ugA6
MuVgidjQm1JJzHeB2/zurmQMokov95Gp+Anm7Vi54NslQPtC3HRFHMGjvC1CsVEt
/Q8gsIlM2+mW9ZOcCGZqA+GT2q9N/3IoXfAfeRAc0F9UfjhfO8NnFl9RJXSD9o7J
JMXubcgQ6YwBbt5tSB40o56V/IANAWql4ORS/jzUKvQ80k1CwgxqOhhceJQlnPZ3
Egwmf/y+RqwxrimnQ1UJWDqgC4NRYz1fs5eeSTLEsQUfmrwiKe18q1THgn8Gyn7l
5mdOhe1jPZvazbKx4msv6v4hp3vRROYKOWGjR/vuyucNH1SHoPYlfzo0xXfgcNFl
uTp+kVeoT0PjR7WHIhn8KmnOTGaIfWkjoNVCAPLaftaih7D2ceR241ghnFOWWnTO
4te/v+Z/o6k8a7vmF6WZuyHjcbKYrKeur3StcWkCNuqjowwPekVXse5G3pAIOW4w
weMZuD7l/Xu5MZC4Z/WoEZAFVRDhxZAq6z1hjS3NYlcWvJ69K5FPZeR9DHJWv54F
iq/VSUSVviNh/WeJmP+wi7KgbucYJOmAx9VQc4nYyIwmExa4kQ/nbifInXnmuG9H
nzQdvBXcCtrgAUBpl/iicY9rJ7YYmOlNGXXPGazhtlNIB2I+WunnBzFfIgEShK9R
zvrpe+WkQNzADnPaiAsst9oC32tzykM/dhrFTs0+PvtRO9+X+VVajtjnhNXbZQ+s
o4UQdD3P7Q9Mc9eT1o71YtPx3nQH7D6sN1nd/6Uj4AyshnkMslB9ojNtz3Z2aKYm
QLqzGnoYPxqSkXCPQcTgwTTYTTtqCji1bvg8L/ofdBPpTp6w4SY3gDjJJgtYlZH6
UNXqVApHx1xn2I9pOFI4qJii2x+VGWvLZew5d3xybmsE3xA08YViK4MZ7s/vVZA7
wHL531p/xiG6t/jn92DeRIh+4CAIfvfMj1UyWVPJSu83DbymedDs8hFAmcjO+osc
xKqwdFYa6Pz6w4ztjNh57WMxCy1i7g2t7g1thyx69hRl/snsuCsU2+rGZf3q1m3K
W+S2EKtG5UN3iE6SjG7vBfrTvsyvmSY7PTy7ElCOb0a5qOkHRGZoMb8G6EbmuNnc
Woc3tb0HxquSO4Pu9pGbNNPY32cAFM3plkdo0MnO2NR6r7iaYa4nJo3VLOTSLTQu
hq1d8gPS2pjJSX0RI0ofBN/fB16I+KuSfZZB4uKSzFEslHc5STxPEqUWCnvDUW0w
WLx2YH3XoPk0p63RD9p+6JgCV8edJWAUn1Sm0mikR5cy1BvS6paMHh9UvogpbjKe
L51ZYqR4KUSjZZjRA/ZA3wPYIi+RN9XxInlXZ9OlCWz9wYWyVdqCdxuqRWF3mTG+
qiIEZmY/65aXvfEy67FREAOR9icijmJL8V6e3pHUK3ayqQpBzDD+rt4ST0BKkbYM
KMgATGtDHSdl64lfPigBC/FgMvuU4vqMAeYDAPd65Y3gdqzhqfGQ9TSkcLzD7OoW
b3O2NbDtIE93PqXBd58OaT3o028lrAIpSjBPHkGAypYr+5FlsWJggVcuJ1uOG3MU
+fC0Gyj2ffUZ3WUxsoZ9FKscYQwIRTiK1mpHP2HNpv0X81Bk0KRw1vuMMaMzebzz
Chd4PUnFDsT3pvN7ROuL8xvXnbjXO9zge/ZXADy+H9xY1QJXllhXQcf+McTlCNX1
bXeNqMVLNo6NY20mxn47g+zb2ZFOyZeadGG4M6enkAP8Q1bG7i2oWXk2id2GlAh/
pPrWoVSdHuHir6g4YmcdD0yZ3y/2QKjyQLY1fuycGH3z7iOiNG4IcwFlLMh/v97w
SrnoYEAHpSxlTo7FvOVdO2Xes1Wor//36zePCWlRTqou2QLtjeCgSwbi6luCj/8F
ex72EJw1cA7DOWTnhe5wRCFl6u1Sn8Sa3NTVNjbEiivdxBNtNdm6gRKPEj29rfJw
i7aRlpWaDQbkTgmth1OtTdegSCX+JGZ4iqTQaMwgr139zZBo6RUYg6MH45gAWQtk
z8ygC5/Q8zwNnPkjcDm4bucwCf2+k1XhNu96sIXz54lSUrxau7AksYIPcVZIyRFm
ORwBeXat6QAwMN1sO8FpFLzru3sTQ+L+g5ubFYpf3H7+DOll73qLAk+7g9ed6OBe
Zf8QAxHa2LmhMzJsHbYqAD2pUndqn+UO06Xx0AHfyggZa7uxBC8itXsjrCSPYX10
Qwmfhss4Y24Bikuukf2/GPlCZ2XDl2ntWI9ZeUUuWMQI05VzalQ68PMW4JsaLVCe
KDwEGx/+lpM+E7NNyAOOFxbwnwFiHjPxBuXd0dzwqDLfWXIrfuSxKt1qK6Mi/hmT
0OluyPNJdnd8hMfLyQFNb08Yr5rTOKXwsFohpgSdxmC8PctpyFrvJR7xcdtjC38A
c6fyXo1SH+usdHpRuE1rxopFzLoK6btg4MWvHG5Dqo/QFjYkBybbOVF/M3teUMuP
C0h2zzKQuo4fpeDltZkxug8KXi+QDuJKoHN8N5h2IyTgthUmkgdiuAgFEsT2vwK2
ENspCcrX+xg+WUZgMBwUPl1WhKX7xeIBLhgX5Bl/Mnx/Li5b/tqYa9GMeNsqSPgj
15fnKNeP5HQznzgVkJypMmCQOZS54NJ815XcAHNGmnfEAnMUpTSmy98F/dOq7/AB
RkWh1q6I/UqGhRrr2BuY4D1Q6nTAGTwH+l0ihNPnhrxrE+uxd6JB57hUx/WpSFei
bmHlmBaGHhqJ4UB1Lzy5GKIaVzH3EFnPvSbeje2Ov7rc6s9oJ+81/eqKE9dDF54m
+HvLlMd0xxTM0Nyci9h9IkNMqctGiNgXo4acanbWx6riqu5tCq+kuF8GNOUcRjvT
QrsrBqYEbfaGhMGHmUXfjISZam0NpArQ0cB8VDLgboNI6OCAGtTtNKHkL2dqr7At
jahOZtTFLJX6+3QHkSFPKq6qgGIv7BAzFG+4ofU/Y8okmep13F+51J7odiiAZIqc
l08hrj/zdAcviTy960oSVKaO5W5dP29rWrRCD4vDiLdpYCz2bCRDrWPMGsNYM2jc
LO2+xbkdGThXN5tH00bpdxynuFWTeFy8QWxgGZ5QzlDVQwhpA2zI0fsPNzgObUmi
n8ZcDmcTvYi35eyYlDwudzelQBFXtuljQuCyAbdIPILFHjrNs0mt30kd+ZfzjmXp
eM2qvoJ4fC6B0kI4No+FQDdkAx05vdCUENZJgMu5mQWTljLJVA2c1zk4ARNaRUfm
DLGp1M6AE96qXdTaLfDkEHGrkjJOCPM0LyxFUebvMg/6harmVVBvecrT1NZNnAwU
UGey+1OYWwQfLlFAVwkQV8vrX/SAeCY6OuZb7xT8Icss4Pjyp796u+thDc4PDOAE
+/1xHS2uU6U4NJ40c2OWBzxU9gdWes1cE30GjDXpeo5gWgcewmM74Ai95UT0YTzh
O6sCZ2yu0LiiUuzKr/ge1cMpWuhQ9mQyd++CnsBDjSvuDnPraxyTERe2JYGKVq9l
YSZlVGd9GiX6mS8nkh4u3QPRqf7kM93AOGUtr3nLgh8jq9vSh/QZHhDFeBoCEWZh
z186vq/tRarXcys4Fouy0U1kVB/FElN9Tmm1jXKdcTWGou0hX1keYLNJRraYn2YK
OEBe8adwyy6i2rbJ3sE2XmRlkUojfnNc0S0JIanqhJnw/iXv3J2EEY30cZayyBlt
24gnJIvN0CgM7zr1K9nZ4WyXdLwJ3q9TWBFTp8n4e4gUTE1hA/9mKwpP1aAG9/zg
nsbQghIEYPtTF4HbqsX33oaEh0M+T9qH4XY0gIK5RrMvBG89u/z5y0W1PrlEGy1H
fuNBCCZhUCoJ2ypvZfq4vF+06yGrOqX+7EcdUEhuvSvwKw2n0SR12JJPZkQtJYKJ
vTrpmmdMIC4UKq4wF2BbquGjEhtWNFz+bV7aAbii9nQjcfL1W4a8daflPS62asW3
arFNKWf7ssXaA+egn5JyLJSXIsqA4pRslHSvo92ruKx7VuDVfFEMcSwzCLDHWavV
6DdiYamH2hCF7r5KGsklUBcoV63x+yYkkfQp2k9X4NSNZdRP5oQMZo8eZJBnypuA
kVXzEAXm07cYSAHv2JPkq69WB11MyFeoInIuiJLA9ale+/8qopBfEJn/pzowxef7
UgmTXNX+w/R0hNS2tWUrCKNCoWe44igWqjKKKx+jg046dHC7cuFWqsTULqwUZjnw
4hnLSynIhObGyCLyBtuopvUlRCPR76Wy1CdpJwA4D8I8/yMYmsyQ/cLrIiiokpTS
xTc1jrxRDzjsYeDdsV3upORyas6/ARRKcj0Or3eiRQNHlXpgAX8x+Hib3GxPo9mB
wMeimr82c7K4Gv6grPTncMPcZ0tEFGQf8lOceNhWtrTyLcnVqBwJjuj+UMrUnUwY
G65zu6YgOthLgtcSCGytTrsWPcVHoViCyYt6CokkmgI6EMqjuEx7e2+aFDcDguEk
dPQg5I/lPnZYC5qFIAykg249oZZ11WJwlhqsHuQ9MpFgj5jwosskYCKBQVmMzpWA
Q2hjUv7HkDIsbc4ysR/SeKn/ZUOMYSjW760UzGwGdoVXvznKjzCOwmW28mnceWJj
cg4tu+y2StM7LaSIPP+8ywvaSkknnQf3x0qkqXoj0axeZ5IojKGk9Ewg9GB6VUJR
UHufQmyyUT5aPP1WhG6GXlyz5hhT6Jaur6fwgH3DSGiBhyjAHjqs/R7QX5OvmH14
bHq6l6XYXKM3JSOxszLOiIKIN2ZZfCWfWdJA2ga0vaeFkuCNkCuUN7ioS1zjjEl2
svrieKwF+rnH5n/tdYzivhiEZxWV1FBDgluapn1vLoTXEQRL0VCERhaNuQAUBFYg
3p11121nEzaeQHmEZsv++ksJwXouRKoeapYC/kmi7BWPBPxD2NMvhpBOUI0Ohujn
juV5+9hX7VP7ZFAAKKLWhsGQ//PELSVrBxtGzEY7TjlGYh8CVekvR8GpzaCN9nGm
D4Y6l7Dj//q0jjW1NqvV195QBih2D2c25NCIA6+fbtRt61A4brNKTFNEYHZ89VDe
LZsvpIqnuWiqpfPEtNNqxDZzq/8VVbbv2S5s+QB3cfEiz/2ewFsZfGx2nHvMLgll
aNfswXy6s3NSLWUi9/FbZeWY5Tzzxr4RM0wtocVLRszSc9KmKat71wc9CTS0ncwy
KEyF79r9AMexhp6IMi8e+6AiLZ4TDEUgBmYy+O75iUggn4lFUKBv0g0YO4pf9MeX
xzSMEv6H11WY3kfPhnwuvVsGJnBFAd8htON9d69nMciZW0H00YqrIHbelvUt04pU
0bKNVDCzfzfR61FueG6hKevgZJ5lClXZedfR/MDRUWUJhMrYCBxgJ7oI/szfw47F
thjppIn9TIyo97L3k3smaWE/bbU9Bjm97vMerzdz7g6cJC7Cf/8ZXH9zqTq9JUou
e+8xzBvOTCK4QLY7g+a/5RMzVulH2h0skPU1fbDv5aOAxIHpv0/uO0vWrPtNe8z2
oJGNiV8Oo/FREdFVeGv1axmoxzds+ExSmX9Nxu8zSyXU9F35LoRKmmiVygBQLxMN
cBbokqlfNqrjQvYGnqqv9/oExVi6aTMQVglP6ZFzId8yVEaiedCGPr8aW9P1mzYI
mW7qBWIxAYGp61WFvidG0ko9L3vdAPGpvxHEc3gJhn23kXWhtaPE5ZhpraOqNtwN
r6fQ7fehTgctoWr5QjoN+aTvgAADD+CkJVVaChepl2+MB9FqIZu064UC5ASqixO+
sQeKckQOPRbil81q0e8oNVU9M19roGnzGQg0PgPvDVXfSsGp7V2913AwSsZ7uzO9
RqRgacN28vgqcxalXd4vhsCUPaxXwuWnP8m/FmAHjebV/zJ/MbI8b+HVxJ7PLoPO
+MUISNhYaNIJPkabENZ//Qk/14P0wgKTAdhHucsUhdlKor82S3B/kzymyrMcsLYR
VfVBp6wn8SBDgCifv+5rSNz61FXqvSgsCWb5h8kp0nCz57pbghIFfb5NFcLtoJ84
vEp6kWjuKdNa7QkNS7ZbpvBJsburoQJPdmOb/gEo/TwzqhkWXhNKeXyk5sybbNMb
Pf0pThAWP4aHKjywJhAk4zj1Luq0Dj0kWc7LuB1qAyiHC55ywATxTaRW9ZX8ZHe8
UZ/tm+YkFHYzCOhlAVAYAGl78mX9R+hkwmdoRtROQzulds65hl2CtL8erPEnlWCV
K8vvjsUUZL22ubYkOqrReW8KZ6Dt7MARVndZYr+PyLMhatvI4lJJbzLBIx3VIiG2
zGb8EczwqDNmf07/Cu7kG2LFOdtq6VtrIPJe7Aha3WRYf1dyosVsVg5Ps2t00LMQ
9gnks/O2LoSazdTDpngdd464yNL0T6zPpacM9AeLAGTO6XpFXLXATEKD4o5N7Qr0
66HMXs4lNVfE6jP99R+T1p5BhhhYf/oO8scEcaKzCQONj2a8mFMHSghvpLlNPiZY
J6EuU1oSwRjOb+YuL/eKurlOf5RTOUaBFI/fKOYT/9PQT8tLhyH17bZZRqfuBK2r
DKSa3pasLx3Sqq0Z7XmSWDFJhIyVoUw2/Kba7sgrClDpf952nEBviP7Nx8WfRzMk
PMI1zchvmcjwm1aQeTUNTgIN2JR7piZS7B3602pNsUKYuAYg1HlOzHZzg9s0l4P0
7eB3zC7piazJ3JUtfyhJD0flxJzkpBy30wGuDob6fkNflR35uimyfjZi+73v3N3p
DOolfFhtN9g6bzCu2Y9Hr2eDyERvt03Bvs8VkfKs11wEt3CyqBZFlrdMZcWjpKJ5
AdynHB2zSeMiiBmYf0gGxJrqPHxGZPvntNs5Ik3HZB6it1KTFkY3OMvKWVWPp5Hq
uvmavy9obKxIpolXDZ+7S03S3kkQsBKyeQ93fjCXiSxBF7RTaKG6ktDxostJaG0z
BYAjfb/GN2P/xI+0yqCCxPsJ3f2Jucr1jqt5vkHuqPMkgezyZ/cAZ4rdN/WypJP+
d86/44cOCS1xOMpaHqelHlrF7EGmrrT1G2Wjrvvfb4VyxjxjXzPitsP8ExXlktYT
NrPsomzLy6qjWwmqslzI2pN3OXDqNCMajb1V6VW5TJ7lMdeLjum/+BLWpgDdM1Wr
U+uvUjjB885oLGBFumzs2fn3TCeUjqSXFWL5oJjUUIcplnSiUcE6jBRHXPfcVmO9
j15vEeZoARUabtqczG9KSHYnk/GzaTFE4x395n4ZxjNJ8U51fGxhZcwkQwnpP1Iy
J5n2/Gt9nWxQHQcE5BTYyG7KMzAVZ8VZHTj6+vortdqWr1Wpuad2WMoNLpxm0G4i
KZu8S742n+s1Pz4KWIqRaWm/NRH4NTYfJLh0o8ypPMZi+xHRuZQytMH/Shiy/ppD
VqewEy/KWBxqUDyHM849+0E349VToRYP+tsHKUweXSCQ7EJqlC5Ebf07Hcc5V+jk
2T3D8VHpAls+bEBMjio+Xfe7XLt+Pg5m07O79ajqtAc+q8SS26AmketANA4sbW2I
MDKrtv2sFvi8hwYE4At+VvQPUL57Fr3uxeZLoQ9dP0towCmmz9en19aOWVHHWVXk
CSsEzHqdvxFkqfQ1thp/er3NyAPyqJvCSnv9E89P3WSpjBD14h5JO0m2/KfF6xve
GdoLXIiScEtBgioj3STRPAVwIPQSDNenDYf7M/BmSOzb0r35Y2Wzu0gA0d81hwla
xiNRlYvL+YFzs/spCvDloW38zcmQlG2wDrIsEolVrT/KQP3ivpNC1Feq2bI24o/R
fy44BXBOSFMkx57df5Qy2qeSYcoWHUusNTxG1mbos8vHe8w01qMY1rMIi3xGYk42
b3YH0jNhC3u/dgdMQt4tP8fTr5xVv9wvSlvh+IoQ6MIMJ46eVo4cwNUSi4zw4wHP
VNOTAtP6APZ2nMxangW8VlwYFDYu8/OFHS8pzx4jUfWMxJZi2xWd8KxGurTWr/L6
uD1pTap4wmq6emUKAdH84VRwJjGd9/ip55Asq5WE+DID88DmW8LpaNdEf8mU9Vry
RjM2v88n/QNNItEPOZ2IkGd1jmVm8nEoS3QTSOPO5sUhTBxxOhzBkCYBKjUrb+4p
J6R96D5ms1X7KM1juKFfmeRRw0WUrP2OhZ6QMyda0zOB07iZFbXr5MmrumG9th3o
81HOk1ZhbdodGVYC/TJbeCcwGA/ieyxt6hLvpPNK2Q+5z6LdRJbWOAOpZLzO/aaa
l0pXyf8KOLDYP1MD2Ox1JqtIydNqnRcmwTphFEZ2derhWA64btSIJJ4NC51KGUFB
dmcGzZJVToobhmVUVS/xjNBhW4911vCNBkov5nUc6jjPazPAd2nRRxl2B4kIZuvf
AyYwlxZxnm7T6k+jleg8YZ4W1s6+WGkg1ojGxl/ymB1sHSDqc/ACOJlPvPQg2AUz
56BuwjkI+p05wdbT8w3kLqB2oRapaNPJEKCWheUxwOJg4lxpzZVPFWMz9phQe7JG
0wohDzbPWXLw82cE28xRf0fg4XxrbKMY0WWYjA9SNG/UYUgofNtsRApbXTRQQI5+
io8N7Qy2TkXjNRbbXxveZGpcd7j5GU1dnNZ6CBtDIfJ5mTdiKG0jTjnvYGX3/IhH
D0RupcINER0AuFv3RCk7FDzkhJnTE9aJXVT7zhGFlrsZIOJhxFZn+iFAf59+2gU3
CTTZu0cOBGmB5G784G8OBo6YM9Pjt4C+9NnT8LsV8xkb8Ci7FKsKnlWCqFOo0CX3
Wr5cWdTvRbD4JRPLuEgsUhjqDCKSbNHiKjeUEZrjbWLrLiKwt8goc/77bgaeCmm+
jAVVbgoElWQ0cmgr+pOirmKXtVbnsH/ylQeWNe2G6TMNH3DCzt/jknSWwILO/nxW
pJ2zGaqt783d22GDzKAHU9LyCTfgk/UgS8mxQ5CeZdkcr48eED0VKkSZfRIYo5YL
zs7aXPlqyxW+I6VR27CpJEnAIg7xXvVzKzQFcLrGzLl4eAIbdULlFvqrPcdZFUH8
3pFurRyP5lKK3UShrY0WvZ3RKBGkEznPr78axJne7a0gnF5U9zNbU+s5uJnVSQIG
vVI7DPXG5eQhqd4wnl4sXsikOhjztVsCryQxfRMYdPiVVUjJxB5ws9oj/oo+xd3b
b/HktZ2rNJ7mVFf2qS2gSSZn6OnLAEj9hv0mW2f+gUrE0qVCAbZD9qsip3cRGOG8
NPfVY20H0obBmivZRHujf/xI7Hj//6qrpWU8wzPdwCMugs8EndvgluN28dKxcNXs
kvXvIGF6u+UWJ5XA/hQ15VRQjO68LEwIXYHsKI/OAEaj/aKls3wMCsBV1Y4SncmZ
ArK6J7tFrg934T5eXoIS0/AMm88ipeDCqRemxNR4AFAv1AacKZ7RqKdIforK4vWS
ruVsWY/ekNGpYhWByIsAz3IZuebB2AlyVTh6N6Z/Lx/XC6LUlV6D5NmGj+/YsZgo
Q8lVfOiTVw1cunU19Nq708E3gf3vIMzmvrkMReI+nlRpiJDXPzbRtTirGl6YPVx3
Kc2MzrefExIB1qHXdMd3ipf4qtpolLCwk+amExgxk8pK2uYZg+Wz6QYOph1Ui+5c
S5f7nQ7FWeakbhnSa75qE5Wn0zWrSNVh9z3RJM37U5F9ncRVFr7cOIIxEcUcqih7
Fcs/iyoBpkiWlaYTDEGgBL1r10ahUIAP0+2+VVco82tHnx1P23gcP4Bl1HfvDD4P
UawEsz+/TguQdKEJu7MfkquMJx/vm+OLAZ3dkc4gaCy8DoZ92lc7nscDEAWS+gp/
UcuI7OcwfSK3zlMdTTpx5dhtVzdk/SZ3fir9/Xa11sI9RmVCThy/LhUH8Uzfad5V
FRNcUBi2lPVypBhjgWy0feGVkRGGI/zM65lRx0hczzK8aksic2LnBpfmWnbGQAd2
CvVEUyFRN0zms50htbiAghX0XF+J6DQeTvV/R5AxqyilatxMWL+wwNnNLUEWtpMt
3DeuJjADRuCFAi+UYbBXvjdlErJNa1KYu2L7BsZvmkb9Uh9j66idD9dZF7Kil+10
1/Sp4g/j3GIYj7rylNw4fiv0DXTzVRo5IEzTX8BnG0OoCf2BZjaAwkjUo8Dxzu4m
7R5NR32SeuIPC1yXvuVl0heiYbaWjF90pa90SvX6GgnDFe1JsN29LgEKUL6CnNk7
IDeRVpgFb2I7rDLCjPBVNmnYiw2RRtNs+tS0PDaVZZukRYyCNkts2U0YA4WJA1fp
axIJwKT2re9d4XgVQX4bdKhjBifejNHac7wFEvaKSW3cI5Jr1741rYFG/9RlU6Ta
EGPDMqQj7OfWlMJhJaCxWWBerfBBStuLg1jO/hWD7rD/tdxsJMAKVMyULklu7wxo
S5NyBsijTJ8cyyZDrZS7iMS7J07UtzVgCwQmI37Ib+J+Vr2Yonp7ApOtIMjPkzPe
w9ScmfRcYBGtB7DtyxK25aAtSNDGMWRBNfnm/jagG0STzXHNJQD30Xu44NUMeVtz
CowcbF0V1o1bR2zLTSEDFBVrfN1K/hJkM+ffwlgoZiqBBTcGzcFvkJSZhQkoYQ0K
fL2780nZ6U8t9P9InY7dOmJCMdveh/wIG8ZJkRFxT6Y+Hu6dzbeYzZH9nKQHdv7Q
0FgUp7vNRm/kr0j2AcXi+O01N0NkSR8VzYnsESt0CyTaPscPn2Ih4HoxKFo0zy/v
flVkG1bA7hT6/8vTpPTXHmAahkB4pE9DyvnElS9XF0sQtz1rZTlL+lNCOPOMZWxI
Ber4SdqSnHcIrh2sgOzRDr5l9JLkXnVs5Juj7EOYHk823dJtd40+PSqUAiDTnO7C
5a6Mi15LZMJGHYhadJpf9weeOzTTNqEa9Z8/riZuEN4F29Bl6Kt+UluGmvcqwgPJ
PSMSpDtRROPg5aYr6/ISXCFXTdukgJAdNJCUiPf+SWOKuss5LDgQL8RNeacpypOw
bvYN1ufGGcuyX38xEcZtfI+LDqmf25UQHbyQj2Q605cl+Uih8fYEC44/68ii1OVw
w2VN+ts2rejf82EFjPS9aVLPIVK1acXgdwxTFF5G4RHFi4fAG+uc5ATWUyj3XLzV
fLDZPOUCPPNHhCCzUjuot8Q19kTZ88tXGPB8JnXSBzfivFtuxnsUr9Ire4Lmury8
XzgHjYU3uVdT3hg2zsFFs0fhst9n+gCTdE0MVg/+0HbEe8uTkFvi/2NYTcX8RGoT
fpZwaFYO0igr1DRdnS2XQbBcnZSwCIfHsUZH/vtqRUqBpvryVpzysXKx6GEW5fzE
6bVYirsZ5zmTIf3F5h7PFwrb4csuGngptlcCxlDGS+IAgDr8oZp0LTxBFYMWb5Hv
54XB8ssHnZ/q2CDzhw7UuFQkvrpUI+vh2X48jh0vcXskSc/Z51Re0srbTmkQrby/
nQBaQeKGBmLW7S17XtS1xpnROegzfHlG3UTkTqxRjhIKzr4Y3js1lXdSva86G600
L/Y2sVm6WS3NrOwXEJPekWIMMNilGTLtOEnWMpM2upIyVeQS4n7MFwIdXf1eN6GU
ZJGYfxq/YC5/xv0DqvE2I919EIRrTcTQYN8ckQTIvXNaUmH7EqTZYSqZcHLaHA3y
zMdwVAxv5ZVXGbp3rVg4hdMKDUtaALMrQOpPXN+Q/oRZ4mBtxMDniJi1LDNk21h/
h51vaKzq4V563w6c/LuUq4MbL0s3w2jmRKMFKq7Ww2Rr58qYL5zxvgMyLMxFXCfz
6zRCSW0DvWpV9r58+li70tAla8GbnxCx4Bu1G+wyYBU2Y0Prq3W3nhgCW4zJEm4V
FkUEE13vHifsC87EnQzKFbohWjQ0hzDoaDPgNUGSGH6xoM5oyOP29AowY1hGZHk6
aYMsi08x6WR0k7Ri472aVyn/Fmw/h2sOctoX6x38AzIKkSgv8aNWbTgjx4r37F27
SnoMK/jeq+6Dimdv3wHp8lm45P19m/KL3XaZ+TBABbk4DUKFfdvjQWcld3nV5jHY
2yzWFOmP0Ayhk5oq6+xVrwIYKMVgYcXI9q3zKKexLpafFSFzRhJRxI0wRRU5rs9U
6YU3CCCVNsHS+rDeG689FTBr4RcUvo5oO7De80Tnlez9XB4Xg3+xOzaiCnJiFZKz
qL2X+vn1ls7sM/s136b1yWnZxOLgxRFjHE/nSiEaq2crtFjR3+tPW3J6VDNqB2F4
xMSOwzsZWM93b9l+331XiXYEqFenUEOONTOnyHA3+CnT7NjhQNVV19Fu/tRDQlK1
PB42eRxmIgyvbqQySaj5SeW/wd9RCqf2E7eG71dvQRMOAJRJoHAa6lgsQkOsLMTy
muPuNIVboz+u4KFL3GyfwiIrNkHUGFe/w7lTitIbqcVVlmFE1b7TI7yXC6NbD9Tx
aPPpbxEdn2cc8ZwvWZns7uCt6j8gTFF57p4bLVxgiY50MJnWPutlYNsufnSxpN2U
+a8Aj8yUkwrDVDRxIAhvavrj7fxEKF5943z34pIO7iV7N2b/fYaJzMvLEYEHxx1k
wg75hhFWHz/HZpiFo4aIM7yEDCO1cl3GvBnh1MUAxR7yvZi7icfPuApw61OAhXtS
6upwqYJHTd19Buh/sb3bHj7kY4uc9PxXJ+X5OU2jkRGyRQ0X7X9lsnlCuZAvO4tE
j5GGhJT3DRjCq0Xb0bPtsNj+q0CmvVA2keMDLDVzN4jL0RHCxkPwu7FL9KGczstU
qj02fjaaNpuEHN7+VhwhXhlhmXksFpe3naBomgDb5Jm3R50QSC5f5lfqOgnU35vd
8ynlMM26CNVn/30B1v2j6dttX/M9dE/q2Akrk+cJP/pK6IEHVvXlREvQ3OyN56qz
z03IgXy/y6nI+FhVEL49kqHx+dEILZFIUN2dq9tA1O5hNTxSr20jVYM7goXtSFqx
6BssafRM16wOzoU6x7K6o8RnRdjZ61pDOrpoSbmBx4HK72c0kwByVlSMDtSppqCq
Av5tTEhbbAFcqd5Wb3ltjiDsg1+wde71YxThblVOhJNiREPe5RFKQuT5wuR8Nw+7
7xWYhMvk9AkDWc5Me+l2imy26UklLlbv5UzIGUn6E4LP5jMvt4gA6wM6gtSo6+7B
OCPMjkr/AbIwU2hUqgCQG9DLoHM0m98HEFWguQq6OWxQ2Oa97TOiv+yG90Mtf9xd
LrdAoY39O+8pYnA9u/sconlyB/qL8H6ppDc0HGr627/rJiOcMC7kWJ1rsfa4FgyF
ab5ClrrG8bC4YwETQTArMZAkdM8nGmu18Mei3ZnEBHEDcx0KeLZQAPONp2kHjyW7
MT4wf+ntochf2olrC0iFdjLiGa0FX5DqsOilJQG+8vseVDWlcjuwlxcjcbc5kpgO
P7Bum5Ok6ciqYMMDPsuJjuxM3byXSkqT2UFX34vLZEQDgHNSyvIZtwyWWCa6str9
r1zyOpbUK3lHNCrxGPtyWQscsXlXu4Sqry81qwZo+Bixj9Wl+2mzwYxFX57pIAKE
kQdQlWPgr3QMJycB0daWuphJkTlPCcBeeZm/c6Zezj+DcJlbwpQ0QVrn4yKwEDQF
F0qNKctuunTWAtC7CE9N3VwddZLOTlaXFrXAt2B0ezS47rIVCQfNA1dHt3Ff6BZ5
U3/rpvYIRui0siPv+cCnigrGMDr1xA3gTGVdT1Q45QGPIYS4WPKxqsvw/csg/ffK
gWa1d9unyWiTV7MapXedTosuPbIfL4zcG7ViUmPXgm+espBrxwStedGyV0sw4zkT
R2bfYHdOlmQINkBkzlVFE5QUU93QlFlawsVr4D72Lp5cpHIRt+oaIi2QCs9v/y0x
hu8q09ZFvIcLqkID5NjnNgdxOg5x2XiGIdOzvA8HX+pOKlbo9tVHBHkkJ0FJOJvX
kNTs9SIQLitnn2rjwHrk5iTrZB872foV+9RnMJPln5tHnI4zqHVWbf1pssETJm0X
kCnH2hoYFQQrGcBJXuha3I6n0YVxOMaiRuphHm/cK8W0rygz9139dEcSRXB2+E42
acd87ES19JKsXWH0Q7PyGuKv/AroSkxf0KHyEDxZby+SabnsCm6JZGwRPyXPI21c
mymLDGClvkP2qMMq87TOsAydOGRVY4PeJ7YVP8bAu2yXzy7Hvy1QmBd24UbBznrQ
pZ8HFUIZV2T7Ygg/O7nZgI6VuzeQ8K73hSq2KASb27bi4tWhGN3ViUjM4e8mZAYR
0b1SgVjN985aUDVtsoeWxd4JqPvJqY01+P6nHW8Ic5U8MmaOWBJSLug6AMJFVitg
8LRdVhOjgHkZ1/tHLKtcfqrexGRk4uReKzzXVx+PCqKrNutU2f4fadzK4bNe9x6Y
m5S3zkZJKcyfDEye6hsn/+ZXVHtatuirP3v+wIrgUK9aUQRjJ+0hj9RUDlpjiHnJ
e6m2WXmtS9iQ0NeqQNWZV1qXAZHnmRdsIzl2IbL18fe/F2g6aMmo8wCaScDfCns0
FXF7ihLPVB0ZfslNWEW576qnTsN4fnq6brhLIP4VGowHOR8uGP1+75YFf5+Hw2BF
uAqbsnpWuEiqfG0fCcK1a9DdkMGykvhcz9QOVRjkRtl+9dwy0MYgKPmKGJ0HUdd/
hfjXGpF5a2c4DA9JZYOLblcc5UuvzHHSkalHvICC63NHU73QujcyFgNwHl/h6zSf
FTcMCwCd0FMgrNBmVOq1ceVoM/9318hLwYmjlwTvR8HeUkzhLNmI2BgpFylqqwpJ
bWapJDK1UT3cnG5dWEWrcNdM0m4utuTqoizW8SwoltBIH/jxgo0UdBAaS2kg43Tu
SqKCRloPzMuZZpeXWyeCq0M0fJ8npeLiLp2iaahFa3aHkrIHMi3HA3wPf1s59fmQ
Fq4JPvjHHieFYOdujTA/NOQnDrPBH7PFZ7tyZyeufmcQ4IiTYcc2+pZzE97Q4+2P
W8an3KkkoiTUeS6Yl6UOu9u54+Y78jhFHt0aKtHlC5LY42c4ha2OfGQZoJJ4YXXy
pbNWMDS1raQt2SfC2T9rTlsU9COOZJ3ucDLBRGtwUaNSYrt3uydKSZah/aPyV+4x
LRdujZhNr/6M2eoS5ROfEzAgU/NGWS8tkpWKR2sG/4ofxp4Kb5My1sF7mAoYma95
/zRx8r5zG2KvyfKfrZZWw4RHMoLu3GjzfiE/p+ta1+ZyjDQA8peV4vH2Dcv3gWq/
dJ943tzt+ZS8eGPXckoa5mgbQyEh+Sstxqrk3VQ3Udvod2+XG24wefeOXhD0gNJY
xGksoNuuOyRODumvB8wkIY8s3WzkmPc4Ex/ctDNHoZpLpd4DJgx9xntXAzNXON3b
+6ddl1caM+ZfmsHLghP7p5NX1f7Urj0KWPLVnpwupMI3odPbtUieEhSXi38zkQt6
ROc31E1Z96tuofPhB7BdAeDSIix9cnB1OaWn+aVt/Q9UrAHPX1w+1xivYsuZbnSQ
V0CLwe9tXJv9ecL/Zn7VAldxeRHXZurdoj5MQLhv8cslYniHfa2cmSMv8U8F5/4R
ecuAa1I/SDeUu4jSQp3nBinnYLfQwFIjV9gvlu51vnDs/4h5NGnW0v6BoKcRA9Ls
3ttqPmOoKMbFhvGGIT90QRwG0oERgDzNZm+gObyRvFOTSFp5o6dcNUa32ukLrOAF
btrZ837xjSx2+vYfgSfbSPBoff3ktOZQZZ1XlF1Z4OWY5RQ0jNnZWu9+zkc1LWFR
fbQbARE6eGWQYX4ePU09JuUamzYMgMcmQBBRYaFGfroofJ4r+g5ZnffmnMEKbBMM
ZfvWpRwyEE4J+aHDtv15a2Fp51C/9Dh9JLPvl3mny/HzMnVp1L5O2LxQoD1cVj9u
NdUEyFyl93LfyR/OSnt2EAuN9FmMM7WzBU4mdYzq0DJHAafOJh2Stc2L2IpQhuUi
EMprReVxmvBKufIqml3asogE4AUlDU6T2CQvZaM+NAkD60t7JInW8OYziFcGy+yV
LGWA31EbAZnOL7QXb0dae8MHZD2mV4fP/+Lfb/pfcFxOCMsS2MWJSthGtel78r+s
cNog/7IJsK1ndz2jXcFY62PeQfubDod0UatJuu22nZUakCPTbiGSltSL8eHyT50G
b94mteKtvyEHvSiQXPvqjf6HQyzOk6f8SDVn1vmtCSYUZ0ByiV3GQgju20d87YgV
7WxaI7spNIAia5y9IdZ6ehP88raJKI1lALkiSTT7z5L0bECdvv2A4F5l0+e1eLdY
lrJCRRgd+GTgL7t+sBFd7f+G01Jmms+71cwD9K9bQPIjUeLpVgKyUountZ/13Y2B
Luy1e7qVZ2AqSSLeD8dw5whefRiCAGWyxIlo3ZZjscgpy/gfnrFLBPkvgKqsyI3c
I2FQkwCMX3l1ZkGGzCcRzV/iyTaxnC9vjku0VRlWobcI09UoTRO3ksP1yhf1QtLN
loQ+M8gvND7MnjTwTeGjNEYB8PHFlZNTcGUqmbhokUaKwYfKJeRYsgAZGzWU3YpW
5eFtvk9xy8mv7oigxhPUZoDqXVLmkac6JhGfJcOIOyFDDO9gj6zhl8bOP8NhoqGb
FrhIcIuXGIRiw+yky3EU/jND49DkGBkTFOvSVxaa+8u14pbKgh3wKt+MP6JHTOAs
KF426P0XEiz9Ozq+jfREF2sZ2ArkxXwASf2qwhpP+CqRPwFMUhkgm6B0J5I2wpYn
ZCx1bhsZvcv/B2ABHfLmayyUQ9q7Gn4Sqf7A+vCoef5cjoFvt0Y8ujrWKezTGVWH
MNp/W81YF2PRg/ong3WLNwFU4ReOkFexWHLl+byDK8MG9jKiz0e34qajto/Bh7xk
otixjb8kjbAIPcZPTXToLniPSQzoRz9iGsndr/BGSGoNGMboQDiHqG2YZArS4OqH
2cVtYsZ7D8y8/IN1OC5gqNM4qwrgQ9L2djPHmKfcwly29EhfwSIXQ6Ql692HbOaQ
fpRNpX35GSbwzTrar/dHwyS9xndWhqi6dV2bUk6ZEagVWf2XgIL2aLYn5L1qZOdh
wvwTJlT4QkGXQex6rud7r87KgHXohmzxxrFMi8K/pIkdo2o82Z0NAASmjHoijK5F
TDyBCTVriBol4uoThmPA1aKEBFemtfAfYgzAvZhLcy+nMyGRHHt8sTWEA5VwJys/
aC4KRJw7qQFTCv1AnypNDGnCvhuxGx4sbLiwHCJmstpCwxXdNPpZX0awPCaI1HIS
pDisjpSBzVtB2QuqiKaeTkY6x4IxhMDGX4/aTW4WXlaW6+fQ2uLGjv1/hKbs4pGj
9tKBDXLFm02bEZU2proh8HLBZdg30FFeb+k+L8ZQoUyWLQ/vUAwsngcTQjnNEQLS
Qk5dl141tzfoaSkFasHcU28hh1FzDZBFzVtHPZ1z3O+rp1MYeFlPKtb0tzd+SfZI
wXsOBCx6Qpt5dULTgO3GtAwtNSXsd1QH8RBLzAcI8F/AIaHVtWomHJhUgzhy+fmm
0RxAgHOPkQl8cHLdeTmsSJkm2TNWBAdT+aFv+6Nxp8NGta2C1vnmFnim1ytOc6fD
5Bm8UcgNEg3BNdV9x0yMjMsNpG7zX49U6GW3eo6PSTZS3QClvIJ5p2KcvVPerK3E
yAw0Cyqo4McG1XLOv8G38GRCutrqLrwoGLAVzC9j+RlGxB4DuNz9m/KJMf45EE8G
smz2G/kjQ785ozRQ8RtxJ/c9XT61oU0NpUotx6Oauxrvq5ah57NVs1TqYyIkdjg/
cevVlyctNqHYY/St5wsx6YunqqIkPnyS3BoayVYHNfZVZT1Lz5KyTWRF9PBl7LZY
pLqCyfMMf1W+g3zch2TVLi1oh8Qkoo0R1yssTTjQLRbQnFyzX/wpYyOx62Sidct2
pW8nA/ll+v1Xuxoy389qrWTpQnZ04qFlFwD2ir/fjlhnytKnngRfOdpvFrjWqt3h
nwxnVbm+t6mAz9cUtV8tQEHrbDvJOpPCXbET7c5Kkw77wjK9fva8SitGVmGhhcHA
ANazDWJFJNLalaAvZ0YIgZ2zd9vcQEJqOqyHyjDKw2eE46o53V0nfBEjkcgVWMdL
kRMeLhB8S6yM9oaqHfrVLbMlySciZukDLICD4jQXZaeBPu1fwLbgC+dD0v1Mx2f/
N8PqIEk3SEwrnEzhcp6+m3v7HZCcQV7oScIyuHXs7CfXnWDiFj6AU9ay+6FGw3Ur
vcsTG5Onei0zN9UuPvM+8+x820xRjTWYQ1GdM6hMoSMeWRMQTrS5TT6MRy4Rj1XI
SC9bBdbZkVb4rqMnBNZRNC/5FjDza8qshra/eXmXe+NnR0rHHW2pFedjm1w4rQZE
xjqdambkQxTTXsiM47tyywoKqj3qR2Hn2F6v5jwEWHXtaBNFnb3aoaUjMYLs913x
vZipEAFRSqz8V7psyCsem5VG2X1maLsKHOaSEmx+rhagBpk/fK7KJJtMCAcDZ96E
ddoRp2TEoy7s+Oyc/bFTu71x37AHrsDaCrhssRxD8dnG9bVOG+pef6NagQk6Fyca
+vTdlZ7pNX3zaLd88bOMytwouTrxVE4B17MBJcfIocNUF0QXcQbCYrX4Tt5Umv5f
Bi69QHX76TcfEqAI1MvR8a3itFdl9NMAGEQgP2owlG3/n2krZUMHkGR5zbhztjhV
WDXr895GvivyBmz19Ll1cvemWpcGULOOf+b+iVvJuQF0ZMxXrcZ7BLs1siV9k3yR
BLQdlg30ufWcHpbw+v3CjFh03tFAPdTqCh8rKFT3eN/rEa3HCP0lE4fU5UsRyrdy
tfD0Ywc/6BLwDutygACvRLMuILh2Q3Z0WHt1ZnDCirfj46CG5reY2PFaC/mf/tNf
6fzPd9TuN40F9a8odf52/QTIyjxHmKEDselrg5BDyjPEbZ92LOIflbkeE1Y2CoLy
YD7KURU4Bnvg1jAYjF90vRscT3gqywZHZ+EOlqJEpeYqhBiisGJdh9waiUqXcKTi
mlX70mVjcPXz1G5jIZqG4owUGB/5U7teP/bTMIxwa0q//dvznSMuBt9AvBqp9Ei/
u5Fgpa46qgbyoz22QgiL295+0BFmLrb5njVkJzLMAcAldxbIOW7uicwKOtz9sDL5
VkD9X78ArhEB1tFCcmmzPebA/0PPz94JTjfjs9Cm6BHPEfyyOzGWQFk2rRmWiuAV
cfTa5h+Gp+KfWtQONJiWfQcyIJH18//+OgUdN+j7NjEKIyUL5I73Utr1p7ZUDb7W
Hd2rFJ2rfEnA7oKUFhwVNDxUewVC43E0o51atJiBO+xMt+bBEwUpXOjdQd9VXzt8
EwNU2MUasZaErezWHAWKq0zQcba270J40gYdn6wBzctwn/gzpklcNlXdSGg+6UB2
p4jdkY4O//XlEdGY1oRLXkULMVJqS/Ve6UW8iug5sLsQZ4S7DCtgBVSYhV8ebvIx
PQibcnR0u2WYoKVkXwP8VGi9xuTEQMzeYsAwjdgAQNX+hfa2Qx7/do0nvqU2ZFx1
mHHSXrwFoNaxofmD33l7XiNpOtmlP/wiURVUGWLVoBtP/W1Pmg9WZS4WDsG0mFaW
pFFGIqiWhezVu0WvWPTx4H2JbJwkSpxmWk07nSaZ2Rc17dFEMWqmF1RbvFCMGi3P
15HUuhbunNtuFJuW13397DwWJDziD+NHDFFTJiSIKk5B3IduQ/LlkZyJaLYHjytN
QxSnfhiyLpiEKrVc90xYAmUZg4WFp99+34e61lmIhC1hwSKy+lulKRZMDO8fGlDc
igBtQHbIcy3ikaQZqGoCTRrFZqJD9++6VMyZc5hMODtKkB3iSgPO+PyHQCpB6Q8b
mZWEmYMLhGZj6PLSDsZyKWwhYOpT4KTXmizUtzZqpzWw5ewYwjtIF0WbXDRJI3f0
GOV09YISBo7NWXIivUSdMFfc/CFY0mJjHKQS2u+yBGU=
`protect END_PROTECTED
