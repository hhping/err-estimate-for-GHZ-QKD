`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/G1jHj/GBANwiDWiVsC/k7iz67zyzD1eJRAYtiR16zXBlAmycT6XAvtHmTZaQj2h
XsuflrNXdLoSZvri6JSlmhs6lxv6Ei6Om+zK1pIDQ6vMH6VkfOcPi0HSO53BpQQy
jB036Gg+LLaIuaQ10d5baJ4WG8Y2mR9u+Cc3rXRFa3p1aj/RSkZS/SHS3RgcealI
1F2fCDBOxJSmhfciUD/X+BmZtx/YT18i94AQfcuPq/02ttB+obsEYPFN9NrukbHy
e3h+IbmbtzrjHI5568vetNeA62RUn4mjIflo8rX1vIEBLWLgQ14fSj4a7opB4Vo9
VwHu2W1V3FRZrfXB5k4K7m7sUtPNgRe5msDjBUj3OWCkLYMUZo8iJtuLSWXg8ogC
0UKsiaE10Yp/jFrnmB520EfTazK4ewCxIpLdD5lu51XFyF7sxJYJ3iA7+0+xaKyr
FI90QazvdBE4Ri+AvQztBtLRgeMS4ui6LawPdy2du3x6fqes56M123IZRFoKmjhY
547ARBGmjMF8yUA5iB6jdmphxqSmqodhid7nPGgGJgDVqDj5ZVAOL2MUV85rubhk
9A8uEUFLFRPCGQ/JL8H19XpX2DwPNqWLHCkVryQkocNiv70cMmscsKGeyJpqhswc
B5kwo68hwkRYUWjtEdzYKR3OdvPi/MwbL9Nd3dNuypbw0KB3L/aWp9Dhz/Xd7N9f
g6ulf/jVWnjiO3phw9CFtZwod4sDt/FaXosVyQ3ZH53yv24AiklzqcwLcYtT+hYl
H5aKFT4fXUWe3k5d0g4fxCsjMlyckwZ/qPPBP3UzEoXN3IGCbZCwRPoE03vUfHN+
rlWdrfjq1oVdiPR8SxpaIvWahV8mgZKaJesxpjjJ5jh/sYiQJ4d6lLo68w/kLtdO
ZH4hfwmjOE/9C6FWaJIxKNHO+qOgei70NCiSQcYhPKxmRXwgSZd5hkXeIt5IgNvL
QGr4neADC43tNk9YFnhF/vlGIzJbpdOx91eDuU7G28XWj4nSK5zYKkkTaiE4KmuD
DFxXXYldzfnoEIihB3cKTZbZowU0T11EtjSyNfX9REEU+YbaV5Rpy2IAkWVKqm8b
TDVhVrg3f43F8did7ogERmlc3mOswIFf109hzpv0OXKAZakzB+Lj+h7VMUb0XuNb
s4m29VqpHyF51n/hyVd9rhTtmFP6lNOT0eJ12ylG0OOlb9a9FUiGN5EkbccyYlTC
i/aYVAB7AbmZQlFw58kSSB13NHhjDnfhCaD93mBGVcNcd+ZrnMmaw/PA0jrPQDGf
TtgBlzSXKoX8fRhYZyGNHM0kWSDRLBTT2WPk/jSCSeq/Xr8ph8NuAFN7l/mbbpRS
eCAPc3nISwdqKzFB2qaYBB5EPhNncKwcRv3Lg3yDMX7LmcjBTxPeWNJfAecEs7vB
sd5a+hONCp673zJgrZ63Cv/ILITS2YqhR4WtquWzP/g976P4zFBHQzEr746OmAHb
dBxOEeFP0qxZeXB0rge2UQ0UMo2RRJpdb6Q7XV6bAL/Ad65rg8jtF6OF2O2P9+HG
VT9RolUZjJRvwX1WX4AtBWVMtGK5s//BmqG1D4UDehH7PJLaW+beM20HeVWQwF8Z
cH5j6AB3iZfDPeXY483GjpMZSMeynbUVeAXv4Nk0rqQMBqWfVQWA6qgb0lZdz+In
PGTf0HKyEaxa8FHF/pGHdFa/2CO5ggyw1TQI2+CUV3RZIv1jP+C5ViMJUInQdtuE
bAFH32Ur3i7NU4R98hRv9tJHU31VpkjCdJn/5ebv8d4JgQqqxgB06grQIErIGrxk
jruFmt6XoRSENiI4J99rlD/Dz3IfX65tIEkt1fMKBRxLdUZ9UcJ/40QVYnh1IVBG
dJe0MRAszYuZ2/bEHnLvL9QJSbOR4uRl6ik64UlA/YvJrrojZMFi02Nn7Cr9Ega3
VYPzb83Lt1og3TzMP1zxIJ/cdJUsWu68q/LiKYiDp5ZsTzbtkwSAB0vzlWdfQHov
jRh9QKuccPci+flVtucfilDWwH2F/3I37kODB8XVnX2Fhaptv5OiAIJQKR3wlwv+
r0wDieRAjYhr7HHHsQPeGq3UXvq9JgrH0Ij9XnccMprsEYj+WzSzJKvvn6bvGKP9
yycdClM06d/5hCKbN0c49UY0nXhBH3WmU4Co4u9v8Wrm2NJ3tcR0/Yys9KLMfifP
/ewSoihkG6vHzk8ylvNYrbR4UxYSp38vm1nriCow6QCV6DvFjtHQzsKeFPNysh51
y2vSYA74Zwa+KoEzlWaPzIin892birEy+SbF2kuTU+YsPLGqNg9n1reNs7rH5HLu
082pe+rR3fXjSZ4MgnWaxP5RccCKGqea1TPEr3Drvu4XMwonM/3RpNOYM28zkwcQ
CmDBzpx80Ire0lKiH6/dvx5SWoIEg5LFyoQb/b4cPFbHIwy7m5kEhmhBXjVKwewl
dZvKOQdPOM//A+qtuw4ekmUEUaU8Cw8BnqNWeHnc3CGt9QTs9K1x/1K1Os7kfCV4
5cc5Zct1o8bUA5CrEjH+GDulJe1ysOeuKsnbiDa0DWbsPQ+HH4PmTpcGCvKRRXeu
NbmV8CMsQE+quVFcl90A6pOgPymwAfF1MQrTbKVcb2gJzZxto5m6spMqOYEu2k0m
t/WN6Ff5fDP6a0xavKgEvglIpPlz9v3KHOf6OURL2hY2dTcZbIc9m6rptEOAEEOD
LBuL6jp6+hnaFBDim+CCHKFVUEuKHkvK0aH1tvJCqa4gY3hG2FR/RKXwPuK3tJgQ
Akee8UfCd9yMwDfNJfFXxb8Yj1Og+3VuILPiyVXPuqlq3/UoMcZ9mzHVCz94tFMC
ICKST6gWFa09956KwEyzTwaKngaV2qHv9VdL/3gQopLfDlUQDFyY39+PfiJoz9n2
AXLQxk53tFr+nyQyJTQDj4Ynv8GrYvki3dgisp4S88C/KEebDlOOA9pBUllW3jQa
1Ows9aCsiysDYW2JBVFndY5JqYg9LXW/nJ33f+KvaTmXrkmduUdl38/cBhMbqA15
GiHv7eWU45rJ1Eb9p7/XQdV/8pKte3ZEJIY53guMuCR1Ii2v/vx/11izTXtyIHY+
/Yy95lUxgfivfhDSHsT5T/K32E5o/s0OWVZRk5IMcOdizfp1VL+UiFyKsqawW97j
02fbK7Z2Cz3ro/ZrRLSeF71lLkuNQaMH9OioYeMePhRdy/FFwzR18ymEYgKOCdaN
vayrJj/6kuV2ku4qgCz59l3ZfoeelI0DIwNn3DX8FPHDoa9q1TaQA0Y06twJYj+D
59yaZLGcy0vKelBkbTgD5FDAUdBLCsJvm+yZEiYtVKRrdRBgvuaCNxNf4xh/2JSK
FOWl0QFSm/C6VjgtRgHBdoge7RLOBO2igHlRz9+vzjHopRpkFrY+ckHgBDMqbo3i
pnD5nOunTKA5FeiQIEkxVGlj3ovpy5v1RwEz4NSudGj1KoZlzDJeARiEY8M9ybol
jECqwa3A3/p95trm1nrWhpjmJhxBF8PZS3OWkTzxXL45xEk1GqwwxB+2YZH1u/B/
/Ssuj2G4gsKfDz7Py0qS0ZoumcfsrX1jEE3o+tVrUC9480l+x3iZRwlLTFO+bX8a
m5C0NLQqrtGxedEhWCfQoOheB03X0k8Ikm7aXJOY0Yut0mhutOqR43H55OOm0q2M
KdSe7ziD6QTVfci7BHvkiMKFkscy0h9+orWJUn4lI/CNOoZLqTXrgXzybso4xUHd
uB0rLohkSBEILzWB2VLmvlIMzb581PTbxf7DGXP2Gcx/0PxqHItRM+xDLjnYTGk0
PE6lwwYtcN/mJb4kqU6romv2nR9fzKgrxJPZOhqgjivzMm65KGTI2g6Q+P2Qy7/V
eX0oiRyWHr2h0vEvBFhP1z8MVA1SLA6ykv1ZdW66d9tBQC6zXDrP4g4uz6f7Lyz1
0vZRpOGMg40tMt/Iyo+XYMTJCtRk8H/wurKSBlPwc20daHc3tO+XQAPwgtDl4otn
Cn1JYLjcaCEBqiJpRGCQWcuY53Ipaw8AqqNzLnpPNPd6/vm3eypUtJTXdX50/Tso
JdhbevVvh5aEEk1gBRTKmzZyHys9xG1AAv5aCsMlmATeHirnIHlgJX5Oul92CVAh
+lIPSb7lOCFRSVFxrrTvawSpGiAS9UN7I5yNX1NyiOLAHNlNTLsKj/QYafCB7CjJ
el0mjq2E0cf5Oyzj/zqPemDgvlyzZXVwLZZ2zIjgkyiBeagIY4WsNda+yhUGg9nm
GlQ2na8rA6XxMnz/Uo1iHJATN/2XmPYpW8tdhksa5Cpkw9tqtl4EWUM+ei7Btw/O
zA+zcUcwr83rZcXBCClTASZD/GQepDPLI+pWI67zEHcs+lA/HPnkzBflmvTrCheD
S7liJgSBTqy3SjVj9F5oh3fG/nSc22vWfOA2eWyIHMs3dIfx4SS4xRhh85CibGx1
mrkP+rAPk7hkyivdS8bm8mkLdDsbmdKnZoa5qh4Z4goAnrI24+InjH8SfOeT1Lhn
huSMT0CCqXx9+3n9MJSqNqOinPhBiCY3PhVFzdGoD1OgQ13+n8ycuQZcPph34aYH
oVMNiNgYJ9bRapbCrHbeXh25EZCNlzPrx7AN0Aj4Zj9rRQLzecf0PgwHcGNaZTlV
OKZ8Nz8YjrkhQyJ1m9pLlSr6Ux28VfaodSwQnleu4PluwISb0EbZxe4tXbRSddA5
LwR51wO5hkliLAIoAJ8t1vxQAlf2AVAT4fZKomGjGb32w/R7dj6/Ti4n6+8HdE6b
Iuld+wNYid2Apn4U0zUFWerMbQpqo6xQO5s5Hs+CiQqX526iu0irqIbLIoOeUoL1
jjGeX9aLYugirmhFjGWTxdtj6a9/hW7u8VSIRGWWf9yIlQF8Oo1K3HIQYGPwsq4U
tHJ+gabKxnRZ9HZgeSxmXF3Y9DLuE++VYyzSSBs7z07kkNnOwiRk5lNarC4tsT/t
nKhcm+Ap1x5MPA7OHL/kOiEF9iDlyT07PHr/kuOZhDRwgh1l3Qm3zjO6UBc4Jzcg
sKHDPwFCMaE3cgaEjox4M0khMtaV5WsCcXFq26sEqHHRLHzmPg+BTZvkMGLS5OOY
OcObr9fLiJ/Rik+qkd7AnPxsNJS8ZhBcgzRaqVmrrItTj6pwXfkfHhh+YhtRpDWE
Tm4c/gjUpjmbVfU/j49XM9VH7KTK66V7bN3bF4SzY+ZliBdTdfLp0FMrCzSGBc+K
umh2heLM+cX8L+y1/SJraNROWFcRzTH2DNDygeFdml82gxLFQmU0e+NIjT/XkDJX
7TPK9vU+n7egd0RpabVA2pPRDKS9niLDXohr/nOkGeXSFoAjTsm8oDXxAhzssVdB
M01pdwvCK45LsduApSh4GlAussPcnaIO9iymtmN7qSto/IYehFhtICzWs+9Fk+iJ
ueGn+RMBdS+UDvzjjMOfbPN0tICkIBip2UuPdTJ43I0GvMbE/9xs0CS5cIx31dTw
3wwoTn05v+UFEh/DoQVU6BiWvy0gO/MNilpICSXRXyFGTu4/N5YBvePoMGenCjHf
Gpeq4giyX2nOLXAwaHM3KAGFrIR55G0zSbEziCLSTEP7JZCwNyPciZpQSGQ8y7zw
LldZWs+vVFa4reGr3OQj052WT/TSqjoOLvo3KLfXNNSV8iqeFWUuO3GavPb8IVrF
/AMo2dE4YQSe1sk8XcuYMe1I1H/YNSpQOQz/PiIisPADYaDk087Kzsq9ssAPtRRV
2JY5yWcBxWh11jB+lWE7RQbONUK8F6+bsXiIv84Rw8sGRWrpZSe3nZdS/fdBcV0G
RCs9Gg+/ScNpihx107VsIM3rhzF8tbyc3bM4CtXfvWinapLKFjpwRiIrFBPr4Fz0
nhfB9q4oXPLOsvqnFUjlrZaN2D1v/tryL1c2Vj5x6V3S/iiUW7W0el5IRgs5rhyt
KzctFVhyPrMNfGB25odqbEts5gH/hGciFwsyQLpqtS53ot3XmrcnlyUOFRKHjF5d
Rfw3wnI7LH+GYwsNZuMJ4xooSHhK4s5xVWgLYU4TQ5b9m4WH93Y301agjxH+ILnx
DnpFzD07PXqv0U8ltjm9uodRAvy1Mpibqn73sEPKBimLXNx9mTwkWwTziu8KqCi1
XzcAlJ22A7aj8uhDIXOLMdaZKk8JpaKv3cYWXs3PljZO7aaQN7XpgOGW2Rkiyeio
igSNDyOQxmqjabClfpZ+HnkeStSUyzZnB1YYizToWBMJszE7qPvAtpmtr8mp+aYa
5lIHrhs6g6aihWozjUBwbvetSCKwUn9JIAmYn0fQWHOXMz/oDZsn21MhTyJt1mxY
HgjwBeuHK62AprIeD8esXlb6OEjlQyMV+lwbA4zPgu7rQJicpQOiZyVarVX52Nnq
viuY0E0gFSKY38ilUSmRQOY2jTgS1v5E4rc08DNUYE3zDAa2w9xxJ6SPZ3MhIPtA
WWJmdp4J0OSPawwkF9d55sHlb/FDUMPj7ZjSxF1tKj1uKAtclQYjXJNFOvKKKPno
AuXN13Cc2GRr42hKkLIL66hEbUHch/3WpXWGC7xfLeOD/bCQPoBAS90H3oSuWl7L
2WtlOUGjPvdspt1yGvMsQzLFeysyWfxVZ/NriBI7fIxPfENMQu0yO2qyM9cMcBqd
vdnbEn8zen+ritk+9wD4QYJgpsB96GeWQMjtm4isOqfbSun+iDB8AO9Yn+WVUTAH
kxn/RFtl0RsvDzmPDfHqENLh7y+NBXh64aYgepdCwJlM/uQtsuG/6M3GRyAwQhaP
scLrd8Q3iDet9dpw4TeMfQQ6421kptiWnHuRE1E0nZTvSa/gkYrYhV96dYaL8HfT
0NiAquy51D5VDCCo/t+7esfDJ7f02JLPOUhoR8LK1do6U91Tqh+hwvW5qb9tnoEH
tcc2Nlt7Ca4liMtLOeHIRydQHF9j1EMfRDywtwiv4VGncalYCEZks3rethgL13Wm
1wJmeD+tHMNtDvs2mPR30PyuuLiNYrpLbj1DUOprX9fQbZkbhXpN1QlnUofYpCDn
2pwnRMovznvwYNtb3Fk3US3tryp97Q1Z2ba6WBo31pjMdOrOEsO2dn5fNXYmvh21
RuLwGxcNMcHDGnznCtH4Oxp6hlH9FleA7M1tjwtxseFxTcZHJDJAwSkPoZgLsdV8
XBE++J/6IqWe6FYkHufakx8nPIb4CJ/JOE+diGpAcN1Xx3YPRzmToZMu9dACDQw6
zhY8xAW6L5W0HsL+HWeU3C/AsQ6a0pDAzx/JyphItc1oW8DWtoiKRLq+gWVxAws2
pEx6OHYAPMYHmERglQ0rXAdq0KShPPH90itmYAqUhZ0HWdKsy3wlIMaTq45qtSbi
A9QKgFMCh4KKUMgiNl7H0P1PHQHtzD0Ed7dRQqO8AcLSf0VWCVZ9D0GqYyioFESx
KJtTpRJTZGJ5o/XcQo1Z4xyYlZJ5Zhd6nolUpla0PM37WkDJ+NtQ1gL9V+Jdws89
ZnNMjan98k1r/4D29J0qixpraw8PXoibBp2GtBzIQ7tX4xV0cGIDBpgt8ay2fY3I
xUuBnC2ixDzhrokF4I+ct5AAo3+LYRqiwUBnKZIilxp+r+p2A6feF55WaIcZkShl
EFBxqPgrmMM9xdVEHIzQMbMyR3EtDg+yVYNxT4lMdkXWFMhe+5FJq60SAtKlj5kz
LpWrR9AIEAuBJkqcznFNXqdlQY5wBYaC/JeoVZnYOJTKT6PeDEmf/UMk7Q5OgA7Y
WM2iFgY4Q5J3mbJA1AK55c8WLwlLh/yy/YDTEEnu0hc5ObtyCW18UgScSgPWc3b4
QetYnYIJDh2yh56/OGjOa2LIteyFDfDLagrr+BbByiKgYIqGyvZpiEhOe4/rwu+q
3X8L8k37ueuHGjBPwkHEowxNdlV7CSngI5DCF/vY1RSvvXekfoeUpTw6YQqIOhCc
lLogBKWq4d5czGdFlD/VvnT3w5WDvbuOjxhN7zCOOn7njPuVg37tzTl+LRRwMpSv
BA3gVMlh4RP3tuG+AR6uRFLja7QQxoV9zV23QVYeMUR6S5AyAnxEWzbFK7uNUwie
QF+15/ayj3efBxzMnK1YbxAqkFf0n81S0shsmZb2EDQhMEchJTFeBW+h28QY39Tr
WxhNix9/OQ6HOYZ3c0k875ZC4X5KUuIax6lgMkr99cBG446cV4FAT+ml6T4SJyPv
pvgvGwyYNHayeXCYDk2Vl49weNrk0eJHkRWYRbA79CoRTVQUNo+xcn3nxYdkTfEz
dMWmceOThXK2POkqLnzu4fOFEejNnZqY0menPsztuSkYpmbGAsXDhXm9/M5fgbts
dMko/3TUg+A1uKkswhKaAfwhHogEaZ15/anjaQzES8trHVWWg2ar+1UT+YcNXCDW
fOvMMbmLJX66vDUtj27RndrB3WnMwwM1hErVpPSMZwluEFORRsbGadSbAn5yHb7R
QDKQgRRR7nga3uAHLsk7l3aq8UwgJ8+2Rdc9W48LqvjECqPWZjZEr3KOQUAJVcOT
ks+fKBBNZH6LWvseKN3ODv2wZWY7xm8O5QO//kGWQwGqFnvet6gjXpRsOIUpD5Ys
El7l7Diuy3cykp7H3fzY0BwdBu1opYbd/ejKlalFNc3k+8sE7SXv7H8VTzzuJxBm
dPRhsA+xQy55FaXaWexXS6CjWPk5MFnEWnTZ6ogANAE8tq/e8SplhmUKUEXdjM+d
jGraNtWrxT0LKdibevY/gXheEaoRLVshn5ZN1pAiT1j8lN8kEZxLDaU0+OSd8N5a
Vx+UUQKSBGnPjZcMu1FJHEedTNfG0vkHTWr0bWNXELAjKpyJQN1EXQEWjqT/Qfnb
1qTaU+2ACHRKw+maDvBURmuREFgVOaVFkQBCCOk046zhBLemH0fANDHrhNzCbxbV
fqR50HD/K+j8vVes0i6H8SRyQhck9e5z85XoW2ciPf44voGhl2vDjwsXnv3jIw/P
MBSnnQG1S0YiTyz/OrVfmNIdvZsQUbOKl7Y5CK381nPmKYV1T9BZABLHF1DNn/TS
gIx/kBjir4tDGXwQW1Ovkx8DkiMlGZvL5IXOkTN5HLgu7TD/qk+n0QqNXUsfKH1e
w6jQFs3w7xwihXzT/4ekv4//yEnnt7xul7Mst5qK/GyroU8Js02yzG8PfTB1EYaf
kumvnZouaxHwzcAkMVlsd6aZD++x3uXU+lL7rHs7mxGP3wBSmIjSpDc+YjvRpa9Z
dJ1FGNWFOL5uuXqurpQx7IClqq7UPUL3qlYjKbSijnfpcCnc1g803Ehsg8GJKMNs
6HqWOgSDt/G3guXTxEgjtLe6jkLJVNMrPAlKayKFlxaCCAcNA30UV5Jjp8qwu2hs
na80GTFBamoTFeQ2CsUwrcA98pQgFMOAsyuTQLZKUxvGAUQjxqJk8YpxXF23UpfO
JWh74O+DCpM+JiJBe+pPvyVb0pLNfR4cG6IIQHFOUvehQDdv6+Q25XhA7gdvqtMu
jaV9x6Vh/AsAOIHEPyuZ5TlELSLUN+MsOLVX7iEuEGUl3Vk+YvtYdkZLvVuh6YSC
MGv0o8tTppjd65tVKCOkBMiuts4kEx7qPeHdZ6zj2u3BCoY+GRTZ/PhlgrUtH0SX
yEE3ypWL3n5lj6FqWUPKydapPd8h2J/tfE0dzYxrGjLPA+zMuD/4hh7wGTHX72IM
3xWFn/wOf+1r7eyqqEx7l95DicccZ5b+pH+HRm1+E44J7gf0mDZnyY7Y/OpkteoA
WOEut5spRY7EtCF8fMK3lfCz98TuvZzlo5S5kZ3zktT/FLA5E6Y/OrAmbtn2XNS2
MroPzg5TbXoRyqJLU0oMnDQsKu8PXF4T8jICt4uFsnUoSiUctZicob+0n7Lb5sF1
O7sxiQ1mDe2O6jVFTnkCE9BJbMZ3epMuUTrRIxnuCSZBITNGv7SefZS7H57mudnw
g0FIHrzs10wHflBp8L6FDOXyHcOMq6KilUYhzTNTcqj55lcQowv4+Z+nfP7nX01o
XKxmrM/efVBtPi0+w/3ybHLDg6/cllshCqTbsebA0YIhaZV86bcGmLT9dVcjUFXf
T0cBXoHNC2nLl0u5kmXOiXRYGqoSNKtVGt69LvDiuFSNaUqeznBZUfybop2kWjia
Yb8Hy0eduzJSeCMP01RilWxgAKpY2uVZSsqPllebWa1gT1IfYn8VveVgyLTMDlqQ
/SRYl/uInUJTpQlbun3F+eh34/1Hm9bzFvCobS+f/Y6mq2NxHYMvJZ0Y0UvA/xij
92PzEll6/hElzRBXnFMQT2iCg61WwFJ1J6Ft2+euWY2Tz5QZKy45/lS+ILdw7dDi
V5l76bnQHhGBuWUDaYJnZbdX5s1QOllbpsyYgaXNmg0hmQ2VvKdPh9itg3iGUh2Z
2dOKjQpRP/HKEvVxW9XlCz6I70/N7auuXS6knBnO6K6KEMCuxz/YmJq9UlhVN28n
tSJRYdQHS1VQXjfCMnKUcQr2fzrW+hgTuH17QthZEYaDXBryJHzoA0qj6Gz+2vnM
bawtcgy6VbUA4cOuYOBMRhhTOqAMWWE840RAWVtr/8e3QDlYIlBEp3miaSUX6ptK
zp05hZp3bfgsAyIwsAeZNcsqaacixmi42wQhAr8dK5n54+JCIPZNIXoHBX1++rB4
g98uKDDzOm7oO1TRGFEvmScUBonJrhENkz2pqN22fIsYlZZ5yXrZGY5jgQQ6592Q
aIE4NIjrY5TvSmkEZUU38jnO7iIPnhPuIzoGbNIp1mKP0wf1JcIOxN0hdhZqKeUk
ENPA3BPfzGir04JwA74H7atT7PbChGd/Gxk7EDirnRwIlRI93JyHU3Gb6vopiIWP
FZbbzE2grUjwMt6Pqr/9+NeJbzmyOZntoGDE+sh3tbyyzD3yNOxv7+LpTNtH7xfO
vG2lVyaGR0qSofikqQRfqha94/CBvSkGYOyrdg6iAAbjlj4vtltaqnuR+cjwlR9X
CW2H8eYX6Zr6ITQoRhMBWpy2jMWQvSGMNDMSNt987WYS7tDeqwBTmneKqp9dzeP3
wyi6K88zHubg0KqF6pUCAC9B7PIE7/SpOenVp7Df1vICwCkg6IVV7dtAxacupIRd
YVULJcHQWpsWumXkrfPnaqa2mHe7Bw7763tJS2I0BtAw2WjX2tN83uibU443IfQe
cPeYe0IumECYAHO6JgrROKPHk5iNaTr5801UE3hFE/XQniunfiCRrqFZKcqPe4EC
xbnS3LrcmN5TaB93dERD0Sq1oIgA7ni4ZuBiZOVRC/lyvABeESgHvQmGGwZtU/sN
qSr/s+H4FC9AszCcnDnaZjSKt0UO5geM9DgYWh9cQ21h9DpT3xoRZ6gmru610fVA
aKgfVQgh1/lWUO2SImMZmuTXUIDrIob1abOFQAjLPOq1YRlCi7m0qw553Z1th6TM
OJca8p0nLi61udiG3AuTQjAJaLgJIKcj0a/25RSFS4htgWhiSLUx4lDf8A7d9ysa
GudXdSwcgcwToJtigDmfpEWNLjUt+fvD8yBOZCpG4wnmzMrRCFlOGR26HCN9SrS3
246gVbAPPih56XdzV/y6kZF+RpZHm0QSSsu6AuctkPbBNynx6pu1MPGikVBnX49W
uvb1Fexs/9xlr1fLBIIgbmjwps+ruah6VUTvvCpWcUUU3XfQuEoKBm87mQjr3BbT
QKWM4+cU9+nJ2axV7vdhdHaChqO/fFY5xIbKFnfS4Kp25ufHUI8Idbl/7p4vnBib
AseoaJlZ9lPQGmIV0x5tnjDfmEiy1li/l+SmBl0IUvjmpQgeTk8t3UYEpx14afWJ
unGFKVu+khkBxayQ+dFuc8H94OvUbzKA4JS4I5UX6rEkQJlEhgrDA5+PQM6U8mnv
gvceaWhd8PBkAxdkBrDsqZ/WMR8UD2cTzS02AQcrg0j4KuIz7Ddm57bnNDd8sK0J
MRsIk7x3qdLIbsr7VPXDc4j6Pz0UOgRVDsoBEOe5a5l+7Ggv0UPgNDvO+1gtqlDR
t6crUD/eSyzyWVPbYfjdkedrETTsi6C8z1/lytAiJA0ztzOYeHD965UlOV+xIXpT
EMC0jTTvvtRtK4nuEa+eiWbeDBMW5LDBxD6MOPmk6JSd2/IAArhsourlJb12HV/P
v6x8Fu/WZyixTp0lL/gdcM26lf0ab58FARBtRrPPOyQ46Mf4DK+f2osS3fjeoWcX
HQqvo04oAYyOR4qMMKH9jjDZXe4hUwW9Qywy93ws/A3wbBUg6ez9ozwI/bzWpZpx
SQ3zjzPOGgqKPxsvD3IVePOW7p4n00I7WJI9XbOeqxGu/dIipTec59KERoN5pi+8
pt50+Qo9qpiXgTjkElMVZTKP940kyRoPZFrD1+ablF13MFI1HXgCnueu+oiTZ9OI
84Ej9PzidViGX9cKd1IpUcZCJ7rC0QdIKF7pKUe/Sz+zUzp8CrMHdv6DFyf2Hv70
qBTAXTS4E/hwd1pkWfW0xq4AKGxeP1r8Qpp2s5P707PMK3o8zIRYWsGwIOjUyobM
OlLx1P1WFZzCUkvTNgEEArPBIU2s02lCsqS5SM5WNawpO6IRW723uN9RKDmUSpim
TGIBsjUSWQWkxMRIa5PEW4U+GvPDQz0opI4GNYTzo0GCgQ+F6dnujgI8Z4hZ8Jvz
5dHUGCYesRUjtX5A0GO1eKpbOElg1YaIUTIham48B00DqVdBDk2HQ6WPpyaPcWG2
N6XSGHvLxAz0pGpXD85ATVjpBRgL2zl3sqo4WjrJIw7r90ZiwUYXLyMCPHJ54D4Y
asmpLBk8AVA60N+zu9ciL7FiVFOVYAySbR5Bdi1pWIQiUPsOxt1J4+rQRThvFIqx
OS3sc6A9jnIpJkDvB8ezA0UjLE1b/KEtgb1HBI6H4DjbpdVNZxJn1qOrtp5wlL0l
l0w/3YMh4omWsGr4cIiDanTS47K8rO5/Ocpa6UmRKIVJOPwyCkG3kBHou5ERHoYE
AJZz0CHE/X4sIGUj6PV4e/dSTewgySI7/eaz/Ts99eDIXB2xQYJfkH+GtPMbOqIt
dP20Txj8Wo+cQRN+59mVaFwIEmWqTrJ9M2ChQ9Bojw89Xf2Lj3vPpMuaEGZlDESa
e34SFeTLzYRdKLiOlmxXmgMZ+xwDTMFDd6VdT50MmMDJa31mvQbXD2h5K7ecYzyZ
AY6ALNTZpP+YNrIuspUMdeTnGFXniaDfJQdfGEoXnA+t1nlh4rx4aA7bE2Vw58oB
80kiwjO0Yb/wnQ6nvpiMOIHFZ2LnUrddpx3CbjKq3FJE+ti+UsgNMhjVK2KMfKbk
HWNw2PKDGVaClCr6Eq/tgok7PqrJRkklcFsIhT5cW0ysa2k/e257zlFKqlDhfZDK
XYCxNNJgNj2+PfivOSsfW0OEUpVEE+L4XHhpn5FszkC76wuVx/g6L9PuRs6TIbO6
o+PAcbZ/aOAvt41u2Oy9MXOb0sV3isxXt1Oc0RiovI+GZee0cHaNZ0NYgk5E+QT3
UdFCb21QY9yX5oUy1U+51BJ/ycXAOL1zW3CKlfjQUNDlVxkDyg+Mc/JF9z0HAcKp
NDaXU4KSs6G4PiWuR2QM3lpi4zfUZxx8vrh1tRDZg1q4S1Oik+ZvSy8xNeKjLFMf
3qEKZhEzlnh0ji5zoJGoEk01qM0VqIqL+3mJzIVGFb4oycoYFjk1kn0eYMIdkwvX
xiX0Dd83mx58Z5CBJvt4asYHirp13MNp6k8b55MYBojWO9lNhT7KnECjKIKT/k2w
0Jmbtj+LYU35Divb4xE0WF4nwfB8yIdPukDqj1bl8LiyC7lpqfVy7QaDGn+xEt2u
l5VoZ3VBqkaIP5eAMMXOH4erpwlsCsqaErepeIPfQlxn+QYIGoZ5Z2eWKZRSPd3q
taZ5Q3ZN8A50nS5mRLaMC2IFlJqoNdqXIxujIRAEz23fuOD/CQLojFPUoceX4NKf
g1fC2ATfRBHcpd3YegW3IaWozpd21nalrqpoocZSXawpIks5WtzvOLXCKw/PL5E1
UE6N2inTS+AOD411lJTdIjzO+X4UEpvEg/ap8q5KApticLWdhVcN3GumVl3K163i
sfw0uIZiR7wrxI3b7KW3s0BBCgKFliPRZ6D4xA/chYkMotFmZnU/vwqoOzGrEy3/
K+YN99pgEGj5UF/FwVhGtey53Ny5fxg1cu8W/UEOD3lj0W2AeYDT3AkFp5u/qjEL
nNIopNAWzhlcEb85n+WSPitvgp/SfBdgnJ5I9jiz3agQk2Z5aXDUodcGnyvtSxh9
u+OMgJEFB5ceWlqmx76wiyhWe8+TSMzWbGM3FM7lAtKg409hOkqVZmrwqxN0EjEC
jDNQOeF63KU1nXJ24GBrIYytBaHONJioinrI9t2VRd0WlY4e6hzfTB1bbyb2+8DH
ps6U95n823Oi/F5Mar9JeSbJuNd+fyjKx7HsAuAtCkpP7JYsdrDF2KWTp6Qs9qeg
LqpjbYu1F21RD2pZcA41M/CzZErymdPB5OcKH8hOvgR9PRfCg9vStZpRf6slKzw9
Ut6hRqtfy+4iyk+UggNxtcrkC6RMqJJdVwDcXSgqFb7d5DgtxBj7utolmp1k8Eza
pq10ACcnCijzSuijasERLRnTnuNnFngxd+YuOENdyYTKdkLLiVNE5q4jUfC86+hc
FVETwHl743YXODxmiHVZ4i7bphVeJn2L3Mszn8DNxsEF6iFbx/CULBnoWkuPWks5
NYGtnqrvBeVw5VmDweXN+SpnlrLg0v1yG7vLpGuDg+nzkHlR4aMddh+BFiG5Oz6w
KdhDyOlJ7X9It6pHm5sxfkSqK6tmfbEbZqLRly/Yot4EopmcYfy8qJdLXAeWVHBJ
znFf2noqEB8bSu7DAA9SRxH8S8gg1lLgjDrbADs/PEi2g8AipFKl/db/cR+KPImA
H4zfYOsLR9dSyceFdBOFBtFk41QpqdcsCFyhvZ9BqydqkY/FmCLqWsi/FVFh0H8w
VusEjZAdoLvzrFUL6XO+PDDlk3y7ArI+Ibh3Y27R+zpRQ1ekTJO9rhxaF/HYSGMH
07uc7TWpcB2URq/0Z2G2jxhgIzAOInwzbMVjYPpg3nMRz26EGpmJDSBcQubwim8/
4m29ZnzQGX7s49HJTANTX++UYO1JTjk0O3cboL+dlq6Cek9cievbTi9RfR7SgMht
TSp0MhzSPX4ri343NHKunU1hjPC+swBcZbQ0U8z0OTnQUSxZCeh3EbQ06ixkdMgi
DjDcVZ15QLN2iQ9jQLjujSuQXRO8Rjf9mSv0BcfDSCN4vSQLhSD8lBeASMZYE8k0
1pqaZjxy6u5dpXo4AXPYV6hNhpAz8Zvbfe2aT/0zpp/uZPBFXWizfcary3QZf43p
D53l3+bg3gCRy7s0/Eo8JhkyGBD/dSMNBLgbDw9yTTYJIZboZyyuLkeWyWMNPMrL
fHQF2C3TPk3R1i+2ym35RTIHGmybUGGOqAS5J0sPo0h6Gq+iwv/X4FGPqeMadzuh
7heJmvcGHp1o8mWENt/mEKiOA8RIS4XK6FA+tJyEdEfODGkYV83xGJnBnslWqrjl
4c3eYgQuvw68ohz2tAf2Mmj/vYP8blq/t5p1Sa4Lat+AuxAG90ROwZ8E5FaU4Xff
9kc5485VC7icp55EWOz7cDIkeN+ydiAnla4o3n7YzfvBcQnU3B6DkRS4NI1ZfoHw
GHS6DkVjPxEGynTKYt8u9XYiLdjxTuXebFVJYiEFWBokXGuvUYwUHBEn9SpPm4NG
tVUZBCYijhk8L1IItxx2OAn8zQQZacKqql9/tnkJSvrqJ/HaA/HNnOWd7SZ9l9WC
1f7+TbGIT++UsdtbhjfvgiXZRdUl929sxuGMCcPpavOUhZA5mOg5xiYLw41q2x9w
oG37PYpb1kDppU1uRd+NzoHvYSulNCoe32cidE5dcNrMyfaCRs/LpXFlOKnweFpG
fS4yXklKlqYfA/NMGFSD4XEGvUGVvDiJSoIPiPYjOHghgiMoqzYyJNJYyUZ3fPiw
U4WFgaB88GhBvB40DS4AZ735mH/KMCh78r4pAm80kY5UZMT3ZUkzTetbg8qNs4dL
+h/1uTbjRxTfr6So1pzcu1IfHTmYXEjHCTs2OJNlw+YMWhiVIVixRsbdu5uEsEWn
GSzBnLEcGDoLHp6XolPbOQlV84rWOfZ/n2CmOFKZTU3hikD8ZN2PzWImUIxwOl2+
dxPy7bz1V24UZPSkGwjcODb9mDEhUXJRZgKw5V4Lr5nh6XT9hFdcKgB57IYOdSob
FiY2LNcrqR9OPHfhrBQUhQy9KfjvLmFYtUBIg/45ayyPmJjAYRNp4s+iTrXpjPTw
R5vfJjoI5xfC4tdZnZUGRtwuAwkDTVmY/dml4inrZjjI53lMPyXGnjHSvJaZn9Cm
T3s5sWIZWtLgue0OeU1j3cb32YstggTT93jQvinNdKN2ojWsTksYKIzbmPo6FlUh
ZYsUxXIi1IUB4LQKWUtUG1J1CkjbwOWc8umdUCGWOre/vJlI4NE5wWT+shzQOh7b
AjFRSwGftCxvDJ5uDS69CpU8ATK9o8oULQZaFUf41iXd59lty0Xdh5YVVh9phPZe
ldFCTtoKpWp3gxq7Kz7RihM3xz3nrc7W39RzmL2IUGuzike5qCsyyVAeEv7XRO+T
8TKj04y7nUP4Qa6XqCHLUI5ke10NtT8CDfdXXopHFO+cJIdqHWJ2CrPNbFtTMrG9
XtTWJHIMVOGkunFETXhwYRoGyNGc6tVvIHcKko6M+GLKpUysQPw/VcLzWll+ZVrV
wWM/6J3mVGljuxjXVq9n/b0u58mnFQL7RhAgHCI4sgShXlBSVXgudM+fiiHiQLDB
Mp6Yj0unMVQg1bsfzXRbj0eT90+rmTF7dBJQAuJNy62L5djqWjGSh0OBBuxRZIDt
gp7FL8/xrlglVDXhC5wipsQRhv84+gnZar2le2IqmNaggpbbzPZNbXfiby7xZaSU
KSsmx84+1UvbF1jLqrGZY2A/IwdhKhUdyXgptFTxJ9e/qJDuryz7/O9whE1ivq5r
Ee/REgcKbQ3G3fG0MyjiN9FmMyaQqFRcvER74bEo65S4BylN9RkunFt6w95flI7s
rQg35yNSO1MnzP/a0qfkNxb7WjnwXv4ovny3VNCStgIRUBB1vilaeOXOQr6gZ9KF
3y1w1YGeLwb1cinYRVFgt6+fiOWJJmwzdeIehqApX143KbvUVu3NLUqGkH1iwO1u
r4IxxbpgLlIHr2CgU3VA8ZCCH/uJ6yXZtZkaPrbp4tIScL7j6r49nznYmlmMytTF
C3XXX2ZoLyklX1zldEu91N6gi32NqpdnXSw8x9WCpnwouSf1cs0U15DQmzhnoWBW
kskddEFqGCizCz0LhGLZt5DTEXXeJLIfjVkzXI6bMgdg/aUNlQdmn8juVA5sAOdt
l869m8ImXRCO/8jQEDOxNa0AsB6KPGcyOBh7HiBHWBs1NVMvEjW8upXcIGya3mBZ
fXcfh6nNkezMlcj5kZhk0qr3hHFn++xj4rZkwXc+8Rac6bicPffDn9XuhHJX7aIO
yEk7u5A5kvHaxO2kKnpkQBxvAD7ybvlzA927H08K+MDuSB54xF6XrSwW3wrolNQK
iDtuErzDxHSIk7lhnn+MtBiraVKWwi5vKvJThcakVEB/Vr5ny7/xc6er298+J78R
4cyjrc0jLXKHP0C4GiRMTgTCDa+4oKxtNog2L1at1tpRrUGwksu5+N9QdqZq+I3X
lo7P8NU0dYU1xevthb4w9dTaq/FbEzY0H7X/qKARLk76VlIuEXGDtEKejHsobFqt
x4/1H5qs4FBs8xwcq2D96Q+xv2EX/oRRyxwrUQ679/jr3rz/GQ2D0q9Y7IBgJ2Zv
CV2P/RLm+CFt5uP0BgPIth1zkSiQW5BxktsRDNZbUmRIllCW5FnmuNFe9H43oEXl
yNZffMkachqpiljbdtkLQFXQ8Hg2wlCeaLp51DuasQoOEVKavX72UavpumzYPzkY
jmJDQcZ3VlriyIHgn+q0TNQp+kH0w5eBiYXsYTSp3WALU9cEllTKpUZaZZmhejC8
3LjWdKzKSIFWF95LBw/JkYUOW9eh9b4k2mNr1NYIhb0Q42bYK+o/GBvSN1CW7Ycv
vEa+ge0pV9/yJk/KGe5CIQKnD2ads744xBbBY2WrXB07rVeudd+xAja0YqND9uY/
pcTjdxxRVQVkccsqg0uqkbpAiEWSLa+6jg4GGRaOjIajIHk+Eh09T0rFwMvkyuHa
FJXaZlLmzzAHIT5Hh25jdjC5ivVRwzfcjCcWvZ0CM9dR+vW0b7ekMk3TQJiGWRhI
1Vy8yzDzMrX/uAA0hSQEAHE3+LePT5RrtW4ctAbMqARRF7vKAR47BZECtA8sLSp3
SKH26ITwZUKanZjzOVxzGmt2wMj9lYGy08uWhxDBl9nW1mdjJ++SEv3xcBcxhteX
DOucLso/ARleUHYynCuSJ/SqHHp2pBkVar4FzYdA/Mj8kb/V4gXb5lWilcsSDuEJ
F1SjWO8K/qPjEPL0ooySFOlebGanAs8agxkV4RNxmUcyT27B/+7QA5TRNyiHSEFX
Bd61a0NKYx1TaM981MRyiWeoQUTRVXK+olTyWT6CGSUgFd4o0DvyfwnwsMFZ2xDN
UaAvXqKDRtVnQ4ZWZienLDDSRsm086VXtp/ivaHgkxFaDbsj6sD4X/hfdmRv/e4I
Nk9oJLHf++kjyxB7YFdHyR7DTHEM00DkGIv+GLa2utGr/8u3QMx5VuTXZzHQpx67
ytaWNpzCCNd3EshrulB0gtlWEM/1Zk+8RH+M6o0O+wFO9X65DChv8oaz1xaeHyhQ
ttLE/AVwPN1QB3WNP6/Q09juUfLDg102y+P2Z91AH0SejDQN0MunPRxZQ2wAd5qW
c/jY+DG1c4I/OmkseKYZiZmEmwiwjmL0/3yMnz8IDht5ezXl+nXISIf7/w4QpvrF
GO3h/YRs4Q++Cnpc6Nn3IQd1ZFLFV+S4AAYCT5kMlpoMj+9cEra0x5kLvMcksfjs
veeGiR+5aX/2JO2rwsH3brC0NuU6QH0X6cQGj+i81ixpzc+WmCl1EU8lCvJI2ypu
fPkCMsURRM+vnECdrpL9qlgW+NU+nm4JLdgjq36B4i2Dv+yG3vrpfucTnMJa9M+t
2OcG1NlY9jegqcQgdpbW5E/FahUQT2Aa7WIc4KWVWLuYy+e4I/qb0QBGgIuXiMC6
0BO7bvy5aYwjSXfycls2qqyMNoiURAUsjRVHxKYGoM/oODo51sidPRvM7VzyEY9f
FQjWdotfQYIlTlq2VjABC4DY94U/R5U5SD1dqAot3CGy/EQZMX03c7UT8tfL9O40
kIEx9BCVpA3CNffYlG+55bTzirunkRkE0d9GwLsdh+fUUFxZyc4mRxK8rYnAEB7p
zEyfF8GooGkkaBM+PUn8RtN3uYWeRG5o+t9mGJZOmD/ru9bBMWk+n8MwSxHlTRRc
UwMTFlNeyLt6smeiZEHIxaNkPIe7lTOX5NKn9Ui51hpJyR6kl+1qRyTuFssTJsLd
8SzNNHuIgOrGe+SD9UcIJz7AK+WBn8LKUs7E7Vxs4NadUNl5F+sl34sZdpH9N/Du
Ipzcq2qK03Qgdj1AVsQk1cPUdxWIdurocsHoRSOWVLLGjq2i/Gd+UterAJA1QWX8
KpWYfYPidgz2Ea96tDglvPt7My0lGSu+5N2XfCOAQ6LLvwxN41UpGyvM03sTLqZm
FHmqIPMsTTxBSIINluitsELaHtSl1r21u20VuROSeP5tYFzrsPFp4cDvsbJoQxMj
MVSXWEIxDpcxUd/ET7KKxbNkh4XYvUWsgH3GBZaf5cYKoRrlkpv7psyDSDUU3WIm
GxMWt/CKoz0fIjEonM8fId7j612AvM/H6SEgDNvRTF7WpHQrNTJqITfjJ9+rv/DR
aF8/5HgIXNCoOrtdhKbhJ4oqzdmd9lzL6gKklphxTkrfwGPX1+Vhor1rHNjch+Tf
2IMLXS+xsSPE5yEl/TO54G8No7bC1Tm7wOhsdrNgl/k=
`protect END_PROTECTED
