`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q/6AxavaI6p/EHp1aeyTo8SNsL3elq5OpsRVi8BSmcSz0SWKywjp3+6Le7UH8jy5
QCTn3DfCq74h2EzEbiSfrsKMOPLVrLLuPwGFYqdA96JmS1WmoCASzJs21aHZC3xZ
WMyOtt+D5Zt0HDphK5xQXSitYyCQt0eTrMO2LFBxIw3eSN6AxqXMDgFqyonyj7Px
lW0+6FPLni6bwSMNkqltsKDuzoQ7Noww5uyXT4147mpCVRgysrD+3HeOKkHYhYfj
HDzg41g1lqsX0rOQGM4w50OnRGGLrUxXDxxLpecYuPf9qLxlO/rdmhq3TWuO5yAh
T4FSYVvRrnmbJeW3F0tK0D93D19EpuH9MkuBWRjFQ/MGHKcMpz0mYLvAlBX0MUhN
GleRRHOBQpC/W/Dbt2AWKjicWcZIKKoIvVT+F3q9IeF97AR2LAo4Iak2htZJzKy8
pmlW743ZFQl83je6QnG+/Rb44TFdTQiT1oVd3d95Jvx4+TLX+p7mgxWKWW6PWzBG
kJVgDzH769Jg4EnLkpUbbPxkw+G8w5U+zj+shtue+dJd6Qql2oFlCDJq+E0gThBj
Jdlt1WjlNbAIcq1Yjp7Q9pS/Th3L+x0Yy0y0/F/jPp+NPBvDwIiaKtUOCCtt6Nqs
uT/Loa3/KXuoI4bcF4+uHtHwHkpzhO7/MXldzN7AWIb3s1SObm3rJV7IRAU/0QKj
4xjGFCX3uj5bYDro0x5uQrbeVEXbsjInI5xUi2Bk/ZnDJ0wLOtyjVNfP80xAeJPW
wwmd2/LOHXcw0Ri7ppiV3uj26Go7IyMcDyWMi3rrDH9z5hz+3w3TSxNoCQVRybxf
TlwZAWWUOJEAq9VO61r/S2LPkgmVyadzEL5EsQBBdORv2i7kmoBOfFYc4gHvgEDl
M6CYC8GQUAwmrbVUsX4mBYyVUdfP8WygwnYk3XgX/cslf0i6veXxO95Y4Wir8FJl
A0U+Ttx5hoTv9/is1D6OQ0H+XT12G+SMJCLNnmmeYqRsb5c8Pt5ONQJua+GJKYZx
otl1L86BQe/a93svUAAIAUCx7J/6qYNs/FiLfYpnP3GShbQvqx86PEwGSIOBj60m
+xqWz+sfKTaRemqHzAHbGhtNDd4PZ6b4jInFbJ2ciW3SkRsR8NiW74zH7qFAVV6a
ffTyqEaViJBjmfYD8UOkokogKWWfCG71DM5AK25bSzTFXUmAS7LpMQEF2pvJy46M
iHLh4L/nImhsU0sPoIJPQfQv6jnTBEX9IP0K/SqYBTZF5HtWZtk5geON8FHsw/Im
5BM/urfvNmUUP8vD26i4hBrnUhDb/y5uUpYlRIW/3T4bPTaLyrbLgXMaUw/ouEIb
RBfqzfReMS6LqTMW9yZTNnmxXjS9oSqesZ3h3LgnxF/h2IVy62hu7vkCic/hxwFv
FBfm6lO9mrbzqASb7fYJNPchI3liMqggg4+SWD5j8F8GYgN0pjCkN8Hnwuval3Pf
r/HhI7Dw6MY7G4a1HqrhJnFS3c13ApJskVRaN0ndF8hoNCd7igsEN4Th4Dd8kWgp
WVnz+a0mVLjrc8IZIAnI3dNhWXl4GQOdvEEN+xqK+k9PAGg0p/+gn0Ob9Y1UMNAr
zx89YCTCLiWd2LybDLDe4txSPHjQZoNdgnjQheA9I0BzNnZWL6UOFWs/5uXq5x7B
Ts0hN+lpH3SgSG+t0MHJcFh/PFObwY5l3ut1z2C5dBZIrTIvCJm+dvaKPlmHTZbo
IF6oDJsE/8lY6WBdgB0ctu0hsyf2QAMcyITvvu3yMTddO8zHtzhtMT0vF/w4tnwR
DQk3hMaEAf2nrHdzWBgjWO6lbc5D3jotSzJPFQQyzuiDlWLycCyU7e7BeC84dAd6
sS30BTvqM5Po5h6NCchwjTgke/rzsxqdGrxkg2jN7XcrHx8DfTbz3NHTTVBu3Rij
l2ZfQVhmQY7BVWrB3LG870UUKIGXdFxkDM9xuIK0Dvn7vFCPcvq1Y9FJge8DAl21
iqUbvRvFwfkL/KPIkjQ4HsN35iB/idvukE+x2drMA0sv1ZPJMdt1fny3xJhv3HGk
Btv7w+StTa3UR1mkb2zZ815nLT4WpEs1afGMTXTr8lQsRJ4iEuatN86GxHWp5cb3
AJU0tapdGtAvz7T7Yxa9ibk4b3MRIq80QYMk+jcdEog49QRTWNcnJrWSi2GsL+nK
1lNsa92k0NnqYMJiJPyjT1Drbdy9RkojPFYBaiyWa66YJAz8Z+irxP3Y7OV2G2RK
i5wXX6ZWgC2vYTp9yZpKGkDkdh4CP+itu6e4ksPqBwV+8tIIYj3wWuyM3mki6F0s
KDDGdaSr7RebW+HSMHDE6hRXB1rrTTcl6Rrw1+1MHCHPeDkWZjc86brnZ732/U9o
HQ5aY8Hg0CoBGnrf4zkfCOFteUD9+Bgnypn3BtxXd0doCn5yUbehvOR25hmrDjUx
MoamVmigL3I0ZAHzvl8cswR0NZoEPMjZINFi5eYCwDwMOG41uK4vVxF0HnxXvZQL
RgM0YBuG3POaUF2GiCVQqRzBCz//+MQFJXaB99cCkSdVPFijNP2yapqd9qBpMsVB
QFmiL3odYL2REJ4KXToL1D0oSOblUYssyiHyrxUgwEGMKEcBpq2dWlZzMSg7MoeP
jyaFOZINzPx2ZZxnzKwtTr6LCyaHWdvEndFqK8cmMbhfWhLzv3aeAhRdk74qA/5e
Myy8O9gCPktlDUx2t/iCgbgFUNO66TDaJIRYE+4SLzfPZcY9Ib0v4lU+/jIqKDQP
XLu6g0hxd61YIynsg9BVbWB1LCvScMmlIFwNcppDFE5L2j8EaHaqVKBTCAQiMgMs
1hDmQ6PVz0vwQi0pPsPthX5sd8r1kSk6Hw4hBJchr/R2Q4nV0n8UINKs9Te+4hlE
wP5QWajvaz8dQEBlGfQeHZO12mwgGfWmOH1iiNYEEPVi3E7PkNQSU8zYTnUewSuX
OzKb1MIU5jRxBZoz8X1KJRdGKq2uooUo/LzjbYA7CSiG2jcqPFPNqq1hMmF1uBL3
6eJxefgXU+2kR1lSMO731spNHyROEnGoCO/0n7EX7NUvBHLKnGKanAFDlExX2JWU
0L6Kg8epa0tLlhqgjVn2dbwswDG6UiHWUeYgmrQomt2I2rUIU4KdeALghgX1kRRr
bhoJymahjyeJLLxMd9ZhyNBlYz5km5NtHwzOzgztAK58FRsnDDLS5jwiIrEGc+Qy
ZHQoacZBgJfLR92bcWqV9p1uH78vK+v9V1TGuIGLww+QEWe8pnYLU8Wm3Zi1patJ
0eUzQpE39HdeYQrwxHIRQPavHp949nJA0w26agIz5VM=
`protect END_PROTECTED
