`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eLZoQdA1UQzyEfec2y8FFU3/Sy8SDkPVytwuTyorE+tKSIpIFKtdNYL+QgZsJBLs
BcqdCZigRcbEpv96kEt5F2KNen17L4fQxP7WqQEPwmy8LmogGrIXjfuOMsmWOmSG
e9mPCvmLC1OhZpGw8Lw9edcrnhNkTs4Ud2JL7RrdAqaHY6oTQsWyb+fOy/J20Nli
uB0Z6l/InLDD9Sd+aiHcGHfi3nIdiHhL9W7pf/88ZbfOYixcm9WUNJBtraVIdnQ0
DCdhLMV/0EhL7yX4oCWp+jwqyIm8yI6oDyEC9st0/Xk48XYgwoB5joAoIGiOi1Og
zWD5IHPJLTQyRQJsrg91Q8eH3czeDEGBEEFwR9l+j+6xam8E/sO9FVfp6Iw+hNDR
99OMOZamUVfGVWSJt1OGjAJwI85r9LpoUROyo0B0UWwCwcU7bw0+B32EKOYomunI
OTvR6/YI8Kttcl4OMAKy7Ttc8BN1VBxCc3paZgzTWPGKDC7n2wlEExUUxmzMyb7J
pcF3OaKdPGILphDEk4koNEomN7SoFdPewbT4k+GtnELtXVVHafz84gQTMt2+mt5v
k+EyqZjo4zelL5TjtYXFMmJA1z6PaCKj5PfnHwtk6cB6dmk4x92g1US7A60jkNHD
v3EC3WTpo3MHYxogXmivEMLO6t0WwcUvvL46NWCmpdyyHmpKbo+GKnswR7+LSfvx
jHon0rqffWo6YLbhVImLYT2V7CsOuRl+sWJB2LNCc1WAITcAnlYYnyZMVxLG+lTQ
t3oTydlid0rvNyyVpFohHH4bQXat08wCTe8QO4/AKXZuxmnaSwLwi5dfhdAwF7qC
uwzBZCdSheq2ir1w3kDgv/ExPyHqR8r22pVnmukHCD4YMRfeMFLYuxOuqBbH5QHb
KGjUxcBRs/an7Ydwx4OAL++NLc7EXerQGavcr7eiCzysW/6hDYSYJK++6sKPp7l9
lZJxTOecZi5TSsjcG/2RUgyd/8chgheSp3g1mmEH3SXfVzUFrIxIkcp1CrKITcPR
BUvkN3Yi/Y/UuoI754H+Pm41BWAR3zwUmB6VSecLZ9phiWojyifr+B5uLj457qHt
G8V+NMypqNrmsEskdjdV9730JBVTEZhCIvislyB+BnyuwILui34Vp8ouLYT0xiyy
dORFMm5pba2vZ2GPkR/Rd3oVyzucnd2pTonkJtNt+tWanEPIriy4JtougAogqdIB
wArGE1kZZ+UNR8ZCig0Ajjooz2nG0kIWEqbLPIdotdAr0MqQNBRqY07mAgjsX2Ah
aDOtLUXXCqXRUt0DgfLyQECPdBYSEPZlT3oXqX0bESrl0wBBZmrAm214EqswdVGy
KvwYS6QI0wVKTwHMfuf34Or5sMHOKyXfs82D7QvlcaqxYiOhdfVKQVQtkQ9cUZBy
EEdemyxLOAAEsvX8PrKN6zOncGnlPPsB9XofzYOdrf3bFHrZ4Mp0FcegLFQ1C8KQ
nmeP/CPP0cGYfvfUOfmGamlBzr8Tv33vGmZNV4J0P+ad/3fs/ZkHXlnB14/FIaYy
zGinlx/nyUbHYNZlRGQuzsx2JbcbLfqdmoA51Z1v3FoWV/Vsotd35FdPSix5f+7K
OJ5Gm7Mc5U0BcDC/tkWd4MRb9aU8W48AqKWmQlJxuMfoiIKSewXPxwpgq/myta7X
m3F9vHk+G4XdS0W7gK2gjZr6dD+3ixyDascc4gOIBDxgP/xEK8XeavSGsWP/j7qy
h6wQ2z6YN1g4XC0DmS88qX+0/hixmcOoVdKpgrkt7fdf9/usauCGyldC8M/TDBZ3
oh7via5PRcrjvYKlIIjEz7gcNYMhd9Tp6YghQjFUVvsafju7M+u26vJQuOn2LAQg
QLFektUQdkZYSYZyPE5LfC0wC6S70dBwaEaSeeIx6scCvkt9G0sJBaEvhrl1Seg/
zob7vaCrAjJa5QTnUH5RDn9u6Y+HXEFS7LJdllEBPTdxtYupEN1SMLtSTPIrnigD
xQcekBIDR7YE73nuMoDEu1hf64WYNj51yk8eLrhPIijxg8CRkOIIGNgQVr+JKo8v
Ew7uvumzAcFoJBpnQOYNgVOxpmmXEgi5amYqeNz2C3i8jPN35hjwy8EW9WKNjwp+
NjE+p67gT6f6F9Fv4/3wi96wI3UVh4P2buyDBcNq1hCX6y8bZOgGyeukvjA111tS
FiRbZWRU/0lO0CFj3Sd3s4armu9LnOxNyA5YnUuU1yoXUed8eBB2Ax64sJWcM7e7
kuMxueRYa4tmfSkRVrazZuIqgpRW/O5ltWBMKsYkxfdrU4W9P+8U2Ee6RCOdZWZa
P4Koaw4ImMs3v2hSFy0gzuagusAHHyZrqYctF46dGaGZaF8MP9yyqULjZX+NaxQw
l2z4lCYhGHsGS6o1KuT0i9caKoCWeJ/PaK6lbYW8CP6VsekmQhZwfIKxA87cDIqz
vwzGrAJ8ToMxViFWfL+kzFuDs43O3PXXyHQi85pROhubTdzeIxvUNBBzGWezJuyB
eTgcpe09IrLn7KhXoxZjnn+tP/FANxCQZYgzkks2Jfyfrv7V6sXafDQrploZhUmW
xcL24/tsWiOkL4ammb99gPmErjhg+S6ydh/SlD0ia7SAPEJPN5cNmeJB+upO9e8p
oq3WUslr1E5bArDlDuPA812nb3YFALv4BqIaS2i6ojX6oLfWRllaZ9Sa6BZd6c7Y
hbl5VVvYz1uvPysqxdzpoO93ihFT7oD1/bHXGTzdV8vYbEEhDhsdEnZ+1U9RngPw
F9ETIc+PpdvTjCM/G8P+SEC7kfFmpkQ1dPHa4z4Ovbc2W6znnUuBaGftMaqLs3X5
66TeDznQgzsfpS8pICaBgQkhwHlXI1tMcBUk/tFAdeTBgUnEW9AoBJUWbBpqCpWa
n8b+NLkGUU8puQEFxrtsPAWcCusCcNLp+4kJKEuUOtOGvDuZ1iKMT0rGIFHg+1mC
ZcuGyrDG6Feh2Ul1uhf4eKeU92QfRNwpQip6nZ+6io0jOvCDAUc1IW/4NFab9d8P
cjiqnX0m1O4eRkfzJq/t+yHsBzByy2w+2IN5TG95lhpiW+lG5nBqducqnuXrQik1
lJjOoYWycrwc0eDurk5MheWsJvTiaAtT9mJz1Bpwulc8bt6/ng4lKIG11lv+uKD7
Gqr8Avce2a11acDwstHCByH9nSP2gM5Eq2oNSXXMw66DzSl5/D6NThUsLQQumaBq
LqhDxT3d6N1yjLDPRyGSokdO8+O7iDaT3NJJ2w2Gvsv7Fwf7x5UCn0IupMO1N2q0
gXNKtj8uwh9r+O65seE147CBtdkXKtU80fzbOh+JpNNELzRgsK4HOfGdDUn++y4t
/hgIdTgDzG6+QrW04OmX5vIXoNovc30TWh4A68WY4uTtbBWrupDhlWrBKy8ddue0
FfyyDzMkgFaVM54AAoN7nVGhuhsNNENeBSSSZPwU/W2ThU2qWetOBhD6cc5cmARI
82sBDDgs7urDU0wQAxCjWlLCUu7oVRAF6/PA2tvrmPUCWH7raRjA2M09VD6J4N6D
Zel8TM9P8lHg/aZ5c26B3b6lPcxs00cfHRWIUyUKFLm8Mjb57bELzmgFflb7PM5U
x1nCFbv9ylX1MQFlsQzJyzJ6LYvywRx09qt4njwIp7twXugERHXfai9uPhXeW0W5
FO6T2V2/aKcyPMpWKb+RIiu0MmcLMG4G3Z1sZoSXFj88G6mlrSf6EOcLD9Ek6xMJ
xWBkKaR2xwJ5mMfXafAZPsXSF0AZaWO3n9+gQU3iPp7tMeMRTZ7c/LESNmuiCrbW
Th+nEpV8LLz91dL6smuG5rZapr1vTtyi8E4ZuemKpDl9VLxlbkcDT1zhjw6RMLRv
Ag/WqcpZnhob6iFkm83N9ywGjZbtnHfkMzUHe3Il5m/4cjU0G1ujqFePXaB07BDO
Ii0GQUQN0oD/aI1RL6o/cFSjoMPso+4K99b1r+hUAuWMhU8ES1s+MuXle/+hPgf6
98w59kLqczp+ZTfV0ukOq69T93uNlgVwy/bn34EFETnCF+Z8EhAkKK1wfvyjEuU7
yFdBMtgmLUaHBtflxGqgArDdk51CKXtSUgw8ezIol/ZW1EN3qt/Dzt/tu0UaWTbz
F90APHFqJ3C3Zi/dPuisogVSmFRD7xiRZmLL161ws15Gky6nrlldD/72XYcwgmWK
ykUMTKU02RExGLRDsV8wvhQf4RnysVLpYStpGFih9nq6IdlB1lghk4R9RxpOHP9n
P30OJlQDSDb33K6qrxyzjsnsBf2WOBJ6DVR7MlHuCVSCW3zZdr7ZSl6Uv1OSSZsN
jx6tWFsEuAC7scQd+gpyZ2yJQOKhx2nNw7y0MJL2x2B0jYj4KvTwYcDeQ6Ose7ko
7SlyG+/CifmK6T4K5J3Qq+9yumkAdqXsqjkhMXoTZ/z/yygcBAa2mH21iQBoBkPQ
dsI86HM0fpLCpNQONBqV7+qMSUNI5fpYDWysnotLvRuH/FZIKTtyfpydDAEitP0X
8B6uRYmznLXu6Eq4jaCkxzFaXsJ/jZaHS+0oD7jwBfm6rVWU/hDzn/VLrdSu1PJW
uUR4ZNiZDJKM8oyAOYfr0o4DQe40UXuXDWli1ynLjnty4t1GGAE5IgepQ5/pymj6
NSEqY+J3Ft6lFkVIuWNxuWOeoi2Fl0enACOYvJwB7qBJ6ryI+BYYbw6uJ6ez3J7p
bpN4q5odF0WIUrM5vC3mLdTRdQPC5UEw1mue5mSKgUMPSLtTYVgnKyPEypmK3/vH
gAk6f48FuuXfcnMGQYQSq7CYjLkOEkXt3106jWznZczVCU2Z5UJ0ZyGS9bc3fxlO
QAHuQx57GZo2olZchfgY9/WQpFl3QigMrWDIEW9hXU1xoOQC+8brKZKmDoCDviBr
YzO5xt00yFUuMe1CcyOkHLNew5wXIwLLx/gaRFhg52TR5qAiDqzaMg6fP8rPt9AO
Y6qy0Mq/7SjwdLOX+k6Tg2FAEmkv8TDcMhgaFy0CVIS6WqmuGq0Fc1q3iLWP/Y/M
VqzczFMhG8bNGJBsz55CLQVQq87cZL8o75caarDrHx4+PIGzpK8Fib6eUo92Y5mp
irbpv3oMWDWOcMe5r6sIBPlkXBQdnIbnCVPNYSsP2DtG80PJ6hzZG2dnDE7B2bAL
INbdbnp6nClbhTKE9fCWxMzby5Km8Me+802af6XvJHL7mVGzuAmKJ2+ZMOjwRK+G
4/mZ6qKibhRwQb40vnQt3bP5zee8uDAvBZQxfQi57XBNG6yMZoh/NAtnDPmfldzp
a9u5arAyNZebEoIh3Qrzn/QqSqye3TMdy3BiWyRNDHNKkdz5Mvh1Cb2YdfdctbQe
gHJKonP5Um31shwC5LJCaOEZwLvlxVrs235uJ2/4WONnRB/vJH4cwxo7nsPiUwnI
s3L6VZ1iu3T16uFRbc0LPSD64vJn469U46wHwZoABsPwM81EhAqKpjJ7uk3wQaGV
GhAXVc/pJpgEeZBaBwnPrFc4/T1bvFmzECH9uUdj+Jb/Cd0AnMbr6aZNUKVXVygk
5X6E9uLMPy+X4KpxGhEOrfAbn/L+dTQwwHOoNhE/tdMvgy+TLA9OTRwmi5q0AP4r
+lBsjNcT3dGh4Hl8iTBeh+rOGg9aE12mTFftTDxzn4QoceTDqgMT+iQnwqbdIOZZ
9fvwfGF5rkGzK5jtBMLOIJpUENDKexcLw7TmlzHKHHxCKcCLzYQMKT/7UkhjDOS2
AsdiI0G5TlicDAt8JakavvK6vrYn5MjfA4ck5bsb4jFXkW2cIvNn6Ll6FZHAjkGu
NwWI2Eh1apmBeS7ZVP9lzuDBPxfxFiQPorkf167Lg2I/UsUBgdV0USijn7VGU13f
SF2dd5GlBau/4J7ztMNSA3yykmJBphCP/W+e769JFWgZg6ys8C+mY4ynUZ4oLyD3
1XlxdJX+gL+VvW6kVoyr4FuUlybSzn9LcOYtSEOyVJttORS1gZQSUqlkgue3hKNv
H6CtPpezAY9p9SAPE3oicMD7HRol+AWd8HmSMmYACeYHVH495/8Pf51f+/onqaWC
+MCrOcZmhOYq6ngzjXkoTY7E5VP8jh+UCjByy5z2BS0UX+xhpbAeP2enBAJs8fLD
bTGaKrSPrJ6wWUhhdtxluu9nMvzN2rO0VS71FDdapRw/7ksNake827/gtyhu3cer
nFFiSQkusgAiH56sufhV7dKD8jlzBQihJtYHI6KWRBHFnK84SDkpzeElDenLpGtG
uksTfze0CsLvhUw2kwAH6CYFREDVtKcaS2QmnywG9bE2iSidxVJW6ahqPA0kuBS2
/JPz1Ot7IjNHZXdtc87tBBrJfMvgxDVcc2i5IJcmouYD2I9C/e5jx4wvZ9MW9H5T
nvVWsEAROLqZfx8r8zMHWb195QTRdbkXpemmE06Mg4sWGwfr8SVc+XLvgZoH0CRZ
K/MDDCAnKYJTPvU6vje30Nl8pw78CUhDPO/dO5o0UBs=
`protect END_PROTECTED
