`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qFiIKIB6lCzpupXO749eOi4v0+mA3TApl3Dhxas4X12/iERgA/V0i+OlZk1pozi/
yDPpE9+PL0bh0+yejMltvWSXBp2H7XVfEPpR/7NATjSVs/+XqqBAMGCuNOFN1BhF
rRLmWvOUD8osjzRp6p426rzcVM/8Pu5qnQAJrJn7wGEAChM7x0co4EFVjYDKWX6p
M29DbHUC/Vz4a/zoMUNCbqQL78v/u3hCd126tJVTeTsUtYhtrHTDafwSo5aTEYbi
OUnPc1/owKqWA6hppdQq5pFL2ZqezJ1VzKjTgBGS9Ej9YURrvDhojnsChiiq9SyY
PdCvLdM1ucwEIVfS5LOQ2cRBd0AaA+OM7ixgQA2yM8ABTjmXKWFmTsScLN/0L+B3
YjPoBLewxbe9QGs6eAotxgREU5ittgf+O+bwIcrauxi2cEQJz+rYD/8F4cHHbnm2
7qvr6EpDfvLbnW1RIkTtq+X+EgNiDdAZSfDGJiQykfWg9kjcR0vN5BTNK6Afnvwu
Qq3+g9kHHhsRga92OmOc7jBBc4so/qrqaN+3EAn7cm5LrCroYkYzr7NMlsKOABbx
qAT6PusThkfi2Q5YF1jr3slGoqQCJF/sh8TP6wthd6EeRuw2z7r/hpHN6v94GYMU
Ejrc+DBDKIo8NRJJvzpVtvo3mZuhGluuHwCOjc2JMMcZbuxO9X8wW8DezsFmdmfS
ibNCvivm43WARAJzwRyXIG69UA8Z80uVl+mhH6XioBk=
`protect END_PROTECTED
