`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D5NsfOj9Dbi/94r04518dp8hv7v6AuZYy6MxLHwKng1M7mBXmhDmJ6Dy3syZgF0R
tvE7IaC+7pytEe8o+2bJC7mVB8+7/PIzbVo0ry8cnHTTRM0Ww6RW4rjpAQ1ROtZ1
ZzbpDlQ4mGs6JuoFgSlh/LeaUZGwsNX3dG+drUFuyYf9y+4pwU+HrXu3pLDV99rQ
a9hdAgFSk84ALIMewvGp2l6sph91x6qVzg7IZYDtN+Kp0tb9yXrELa3vb9Fc+hbi
v9Ab6vat0l+wCAWWF4VlTHUNd7gN6O3pN8Id6wUgRlYGe+0FPiecm9UHeH1Ap6ie
SXcMi4+Qc0bGp//UDmXBp1fY6FRvBzWbynhQhWnzjTawJDrOS4yJiJ314a40c2M/
x2+zAajRdRiSfc50U2nTV+kkDZh+gbrK6cKqKKdbKHW0xqshL3aRsrXMydUPOGmx
lmglxzJycKhbpnET/k9anjTdHAa8DpKLVXnh+W8ajsWw9efZ2kwz08lY86a8KcJv
EhRsergc+JmNOUdctzWygCrx6ifYrM1GG4TE8VEnFA4sqjiYrsRo0gMzFKF0NQcu
6qnnmjTqOtbA+AD6KA0Tg2Rb7dHikUacAF1lSH3Yq44OdqzK8Ik7CdG7Je7N2L2V
15GE2u0pDW3M6z2GaV1xgDRwBmI3F9cYwjyN/UA8u9MvvC+Lyzgg3JGJLK8HSbQ+
GuVq78YB8IWVzbCEH+Boqa0gk8V6w36QViO5G9prTQqIa9/AgzJlzP4XKYEfKsGg
uTgv+yI87Nfcco5/9PhcueGGl1H5nVcyj7/Z2+llO0/pvMoJ1rNsv5boDgaxZ98S
DE83DXn+qDPj7NgknL/4gjNjo6mO+5NgY4YZmEkEPizT3gDEg7xQdv1BDNtTCqHW
LCMofBk5ASatAQ6oiYcSFMn0cj2cZqILTUhaWsUl90v4y20unHs45zfkvFIJwyei
EWEc7DZjCAD58zcLcHYK/kckkDJC3YSCT8+20Y0qTsc5NaAE9jF+4UTSxYfKAjGd
RcdBGlJo2nb/0P2m7eZZE4IZZv3JEZ1fUotC5bjFyf2PX1ewQf9oYZfF+ZP414tZ
sHR4d8K94qExWgKsY6ONL6bNSWqkAuw4xRe6fxXfeATtZUz0fhsqkzxdfUJqqbnT
8lA3YgL0umh4BVR2bXj+0duFwFIoHMG54uND7QbjPM+FjhGwb5ND0SiNMw7b/WGJ
fQ8gIMXrJriFu0SZ9VllDdwxStv0NWzfgsC8+Rv01GgDIIJDyHG84zGRbNjKdYxU
ePQ/WH5WUCCJzNMSLfjNDzmfVLbaB6E4sCpFYSKNKwERgmy3keW62zkecAY7JVUV
Y/lZ+K323rPlwJc1DBIjRA/afDivHJCIu4iUQch71RkWbDLRUqjMJx1dHGNxofsG
AY2F6CWyDwjkuTIS+PKZpznsRhBcgVyMJyeutDOlabPPQca9aFLxKktyJVSDAVA3
dc2k6aT8zpLZxoekzrG775k+9TCmvOGeVtgk8a4uxV5pyEWMVLxLMNzH45lLFhxD
xXXix4N/eolX8M4lsIB32WhPzBHImEMW4IUdzyljK7s9QUBmcAbldIiQDr/Y2FRH
6htUmZPiOb7713dt06SCT1t33YIXTrzwjX9rWyIy60a45tBBhHlghgC/M5QFEIUo
rqRgKBM/DuFW+eVZOvM/r1Al/+PHrA0GQwYBm0IKJhUnDclMcNDbV3X5dU01il96
3gNvNidkqUQyAX4ppVVIO0hCQ46HzsvUgV0iCLn1tgEprkJKiM+N4lF10oSk4Ho2
dx0n2y1y2oRNFtaGTzMedl4qLlnO5XmnPLBlDKAhg/FrXbEilp8a8NGIfCkmCaQy
fsFiO+0+Jn8ZlMLGaOuKRD90V1BwQapQngwlZCvRfYKu2bkyhEH1+dy69KMnAOcS
et81gI9EejjKcv7eQtJzBVI0+tVusMaqzGs5q67KcCfQVj8lt+/ZQnC65E+vdG4n
4CsOAVRNsE7frGz+6cjh4R3InUojDXCnsUPyLMoe627K90I6C52gxDN4DEAdh/lu
OF0g2Ir77hdDU5qVWaITpn2UPbG1N01mLCM7edmbwVZQAd+aPafKYDkEr+r4UBbP
z8rLmkA+V0uf12UBXGMKiAe1x8XiWGFEgWHistR6ijeGaiWi8mqFq7Zy66D/57eC
RyNMmlMYTXJoVZ5dPvvfbTSO2l1MLFnmgFLb1c8F0t4aMafIXi4wnDpiWqE19Y5g
En6r3j8Yz/OipW1abfkOxn/6Zl1m0rQmALHE78gOCUlVIJsxgsoFfIEET4V3vy5C
7kclZYdFsbBDHKVjf0sKxw36U+6QUk2hmrhqpNPZJlEkNnFN2FpMamPUb2sgMyYh
GzCNoUANoWjE4JtrlGrKHYx3Dm5y4XvMs93Y2wbb10QYZhrdd4gX54W9whe2eVvR
oiJOZBG7WNvymZKMbirVmhwVFuF8D1OfISnUG64Gi5C/FW6ZKeNtd5cKL7PtNPXl
PhfIIKB5OxOgSJrTTLDxf3KQhnkxDkQHsxZ6fz5Cg18CyUxxRZ6wdSsVS1gfrUls
H0aIiiIQN50XT8Z/b/B8Qy+H8somEREz969sdVjBck+ECOaLxVO3ijJFWmKTmGgN
wCO7q2//qIs/xF748j5QUOzOLsofB9YPSJJtSQZQQxWLYGltxB4QTfUM6yrJdDey
8p5KpO5CP9tD44FvusGHRnuwdV8iRqpZJXYXxfqdnrXZucnwFmtZNoKhpyjmbUTU
n800pkM4lekQykJxxjDmnDhCSgX9+EPqaPd/63dOxkbEVISe/P6dNFSRc1sxmmFN
I9jVQAbp4awGQP6DSXL7nMBJz6ZFmRIKQtMhYoXkP90Qnr2hn92Ft57fu8wqDg6N
lVWTsd8t0JjFL4H4TptF/y85SjyLM00vCSthqe7U/I+45uGGVOKZi3oczOD+5+S6
HJWa8qqEDw1SB6aSWiE4t6S/HDa6MuzK2ffiDvp+V8fiKztJooTgxrZ3aWMpuBvP
j85DH9Gatlsb2Je/t1Qzwo4/xGxI2KdFZhzTU+F1opP8KjEPiAF4hkT5zz/ZVLw7
5Dvqwd1sS0GZ4w6oI6D1JDVD1IskyxSmaDq7Tf3x44wZCl6oxQwiesHmuFCJXgsH
fekvfqlCb2qmiTqaM79WWA==
`protect END_PROTECTED
