`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
52yO0fA3AxwDo7WrTbi9+tTebf0OxSzR6jiKetFfwNuABz0kId4+o8EyVI+wuk/2
mSntVeOv/mtq67StSadz3R03jAxUV4Yafm8kC4D3SfINeKB4AMMaBdZk7TibDB7N
U1gRjXuDEGSIfL17eTkT2WyLh86kKB/P+JFGLC+TwXWd4vo5VaSvU9XOIrRgNdfC
XBKW0rn33013FO3GD7CxM9oLz/VFC4/LJ+aUAm61R7jZypJdKbu5yRw+M7MDhugz
HNmG7kbAT/DWuRxPo4XtOZ8dMRQEm/REyiyJIVO/cPUYZcYx6ZEG+EX8QuTD/OOK
BBV+Xviiq6tlVbD1e7c2BJu4RerXfHkSDbMzxbkeeKgCetMqnaPKVTK+bp4iBhgE
p3erMf7JWveqS0qkF3Vg0rhW9gGVbqfNZ9+wwFS3meULguMp9zrZlr+HFJGN9hTL
x1OE4mlLfTbp4SJEN087+3vlwkVfgDwj8uziLfiWuSn3dhlDhoCVKbqgbDwfhC1x
u9WethxHQ/1YA87LrxNdXUjQUIgoZbSBvptR7msadEY3Jq9Q2C8gSzww/sgJfJen
Ois7WGnwc32t3paK/nZo1dx8yn58BTPusc/qW+GCfh5aD96OFuQ+qGV9n2dtcO+L
NbRa0rR2v8cwu/mw0TXXv/70+YoI9Jo8sClCry2P/NktSM0gKtjSOLzlnp+RFBrm
Bv7rDA3jWl1MlAwGZMK1Yr9A4lpK5g8ozWsfNjZEQCwcI3h+yf4+2mLKWycyYqpn
9R4GXl7aJuzJAzzJQ3cgaWtMPA7mp0o9nkuE2B87SDw3RK0HbhZ+kvR/OAIVeZfR
HwIT9Uwy/0LBjzC9Ua/c1IPeImQi3CLxRfVGJ31F5DOAHkAPo1eNhtmRlV2KfOUM
rkFexpYXssLBYA8a45ai16eaA6VjlhQhWfP/KSW3JEKgWgXgHmtqfk8obunLMeFt
pKUAcs/r3NgNeHSpD6sWm1kG1ojbyQBVcRxbDkyirONrbJ7xQAMDQ+Tym56zCQ40
do9gTTvKXZN+2KedWy9Gjgoto1RZmIL6kAau2EuPPjVAOZ/2xCXu43PmPErpXGQ8
V2m43HLjbyutZw2L19pPU/sqaz2qMEg1Qn1z6fSKWtN4P0axh231Hd82sw79ivP7
L2VXtLdF2jWejek26YTjIdXwhsvR/XZp//ndZVdFB+LgONpKGDPSHmmh7QROTaXP
ouWo3+SkWgIeN76FTOwErFEqxQNiHtmVww9qMhG7Vq99GomLJaNiJjPt7mo3sy0D
3OguRkZiUpNJJC4xwUYMrMI0FpIBorUyRtF5cuQsp2frvEz070IeYqfNT+0HPaFH
a8efCXO/zPnU/98f34/Enmv8cVqBLBNofpLTdd79jGvfyvWyD+iWr155nnSzcFSn
g3wxRb0jxlFDsCnd/z3tXGstpCK/sgl1hxOqhG9qC9uA2nAT+XIDJ9a/fzaagv2q
t41WLcjRBq26jxLzv4vY27ywFWZY6wubFgHjBfm+I4eV8wQSaOm69O5BJ0XfAji4
uU6iqyhsQ91UR1DLw+/h4m2YlZMw2pRBAwBvR2zNNC5UNIoby3E9rn4bINqZhPAg
74G66OMUUXXrFYkOZFwLzs8zjLlGRMxiBlhfVoouiE4Pb+DOBZlrQ5mKeKWfUzVn
9NKEPmMpE6yR/FRUHKnFlkEPcve92iTulTlWfgC/crDCi9YiWeiBOI268X6ZY6Wk
FOxVUhAU17it5vLVnyyjhoKwubTISJ2QZSIKuUHwlbr1pDaqK0T6hYOsjf6ORUbW
/OlHotqVuQXzH5L8QbBbp1DzoYaN6GWklTbd868dNkP0lcSVNZ9swzPoNTSEnzp7
vkSR/vOdb0t0u8AszopOXujsxcyuaxhGBMKS/ZMcvGgU3CCvoH1SOW++T/JvyPBV
zDb0uM/nl4/87FS58aZT1Qnw9S9IqrrftjZG57o3gO5ZnrOh4ipdArm1IudjaQc8
Sa5X28LOvlhNGelScV9D1BrIb7Vd8Ty4CFowE0Izyn36IDzhf9t70eCuz+IHNiyp
Y14zgX7J7fa6dhSqgdFWTiauXUyQBzI4dm7JSEbp+zzd7/Nw/XgeTy5W1X+KEhWE
p3CtcNXTB0nHl7dIJ7T4L9satVRr8bhSj0IVojVsCuFmn5Kr3mntEno7Yp8a9sx7
gqj0P1ob1RuTHp8RiQdKZTM1pGETAk9JCROF2/gknOyiB4i8ug+G/cMQHxyQL5Q1
s0uAl9IBD/UO3VdyJ/iTZcvt2UVK/2tSWPj0mBdu5AlWq1Ati3qVIEYkncttS2Sw
2K0fi4mI01cS+3LSqNAFsa82tmVJ1y8KXWZw6ZBY3K7GblFrqKIN9iSYKHzU/hCM
qYLb8ttaOpCxnZKkUcX2BQbGZCPXyn0O/4NTX0gCm8Ct4EpzTAhK9aDjf5g9U3Ql
6mFKiGw7BYts0Exxsw5toSG8RwOFZP0crsv4b+QL0kfgVW/JsvG5iJ8N1TVSNJGb
x2Etrt2G8/q5I3Wkg3cGx9OhkTt0PDFVrG00ltk7Y54GNWabrBAHd5iAmNtrz98Z
bRAojw6JyDKhqmhQQe1gBZgDdHWD5i99aslS8Xu2PIm3neYypwqexyLdjfZAHAym
jivVfTMR+s+kAfc5pbF9kONO1yQTzxttTeZtmLfvNU91cwphdFRdFZCxQV2OKKbF
vPRb5pS1FqjKOX64JYDRIOelqJ+v5wRkkWKi38LJQlvwXvg6QSeqZX4mpGnTUEcV
Uo2A/DK5JRlds/RTFLmEKbb9BW447qh/6RulzoAE6Xc+rHcGOGyo9p2mKMZIMXmf
jiIPilted8lQ1Nnwj9Bnp4NJxMOi1WycVZ+wra197ZlzFhUoI3vY0NJfFo3Fsejc
FfOzbPA2g8BvSaU7XzyARrhf8GlxZrqavdRllD+7zz4t1CuubodXIyBGvZl6ubiv
2TnQaZPvtoU+5aiDlVcR7auzqnCz2QkiOYuaMQHe6jBwRQu2y92oS5/o1Rov1asq
+NBEpC1Nmxk+qwibSpBcqbN9ykfNjkZVkdc4ZnHKKGGa1C9rof/30FVep/m/Kiy9
emp1LvDVHNH9cTB4ygcF6mPDaXtJ0pD2JigAzVLDmB5HmI3JSMuxWE0a1x7aKQlv
TavqHychZtgM+7HlaDpsrUgb7knuljm4lVF0sG02A3CjMFi2aONa1Is3kF+toVtW
pS7/fjEf07PtkYIzs4sE7KIfUqjF1mlL7J84tmbXvGrl8p2gRvnejTItopCfcS9O
Lci2PcJ3JqDii8jwnzZIf3+h4ghVmqnlVCDjJDQRR1lSBqK+47rAXT9aBYMlT+CS
WwdbMIbP2M2OkbBGE7s7r0y0wycdEMRwDzVUvRvSQldezAlgKfKq1GmrCPkmh/vg
G+xed0EoDg6FeA7n23d2UN8DR8te3uuFXENGIZ5qStsJREFeEtVm6T8h92wA7x5M
iWAEagwZsDG3BoA1qrT/FTiW5iztmSe5O55qGgIseGsIvVRo2IV4prn1pqv39YzG
bAzvJy+Bil0MiKoG6YOEfOVsEpo1sjSrl2UWRcqEMId83ya++r2WH8asU9iELVfw
R+Q/UX9RyGc83iG8SjMenoSM8+9ObaDn0QJu5aNcUlLo8e+zWuibuAPHGQN3MygY
VSQdCKsIhPwcMUp+BAgnVfeZYFiM55fc5xwjyN2u7sfmwKPrJ7yMeieqQz2W+w7M
jnGxxDheLPCp5QFigbBlGtNhWz5lW/+frrGtjQafPDqo6x2h9dWSfXbdnxmf6xXX
sja4xtroztRFdwuAJdsdzRcv8VGUc1vl4VwIeYHX5GSYf3eHf1ybM93srji4v2Qs
vUTuu8cEK+FT54ktlzbny5NYIlKLUs0Iix61eixFebJetXWNfUfoL4J3dGcuKd35
jpMxS4zyoKXEV8RUho1o5PMYjb3ARY2OqX3F5oCxOOC2PFC2OOWbWZ1fWaOBzKGr
VXKDWEXbTp22pvWwKzCB+58uZeKahs9qVUTh2GE+qabKdZHnaBrsSjTAvk9GSf5V
qvhhPuHrXkVW3W5dqyHnVdyRfC47D2Mp7KIpFtNZIFuGi1AllhQpVg72eoR8b4qI
AeGIbGtqbhsW7/fXwUW/YsSOVEgFfJUdbWAyP/lfhV4QAjexRziKdBgPcbUWDECc
J+ufAZaoQrg9pqKeBaLbnlASTFZFu6DF+TZbEmRjDkLUmN6rqodzAAGlz/FPietV
TrnCLbdYMh5NnR43jUFo98YiU10PD921mHjVbo8AQ7eVf1YV7dLQSkECvwe456pf
DcGzZKd1tnmpwL74LD4BJyIcDDUPeE2U9J+BOUQOFyLVH79KMDvcWEaElwI8R4wl
cLGQz2/JkXUQTeugVnzwCaDCA+SD9//7WfRSJIPbRoaLv6sT1gqQiBQyFE4x8waL
FTzub/GOU7AbiWLYAOIiClkdiB2Daj+2LpS96HzVOEXOtQ4dbIS87iFscQd7BOCx
9MbKUTiyrbq1NlRyQGmSZKL9QJWHMghiGamEOGDSlAONrmsTniqVV2SUJMF7VMlN
A8CV8kNwn9jTEg4v7DtMNcDfrg3OWtQJ5LL5nZ0orwNNPs3TlaQ1TNVVGa3SVjB3
K9M3BMmhRlUTypHRS0am/wY/ngAjd85n02e8HFazz8yDKCRGPE4r1dG7LKsewFNz
cyq0KtyhmPtPIzbA6BxM/AJ63uKjDj0Qp09EQCJ3OsjI4I/+tT31cTL5dFuNrKKL
CBzVSFiq/Q2ow67Kv+3pL2FxUNnpKo7zmBwQvpOj2hTNhlaYpOD2UhCiY3tu2Hpk
jig+DyRw9a7z9zuN7vB747/lhCLSEw5U/RIqIiRBY262vgEKxhozqqoznjhpN3ep
wj83m7NoiCzCFW7+Ff8ElB9dP8EemyH3xieYFndupk6T46NtqSSbq65eV8YBEmtV
rKwgtKxH9ieta77FXeoJcR7Cas+I4gqQrIcKqh0iCvEXojj5wLOjrp+gxtwTadv9
SYVW3gTSpwuTsEC3xLutsGf8qTMUhHFM2CXM3NefXpBAZ7TFwOU11xgv4nvw6cm2
ACkf6rBtyfomvEu82J1n6JKOuhVwrNJoH0eqlA0fkF3K7uVHBo9gdhyNUJzYBag9
kpQnJ0g2EqVv/qBLTXECsR+Ifret+I5cdxU618D8OkLE4u0Tr2t1Sq2sAIWsvGHk
+tT6vTjOzOM0TwiBi8qrR/uXBqDvChe1Dw29nPVAKxPWBAgjuRzBDXal9LE+i/SB
iPCe2+MBiWM+jBxzPJYnSazVpjPHWWn6yYDLwU7HnKE6gz0v4TzjT/xJNmaI40gE
HpiwMoenRj1cpLF49muXqfsqxBrSDr1/OlLYXlfU2dBvlnOizRjEUch+67QErvb5
j8Lv9gbneXUW1FYT52olg37AoN422ANmUoTBdP0kg5Rv0sKJrZv1yHSpcKsl17W8
w4zLhQ35G1vw48Mf4U/rvR3oERW9NrtHS8mSEIIYxsLuAWd+A1ncPi5aEr7kD7+O
eEKM6G9/5YDhB5JPiFmObUJjZgcRa57zQp7MQyWihwhFA3UL/weCt5T5YYWwL5f/
fEXYS3s1pndeLnIVgj6rk17xVozwn4vsJtpBXVbsJZOdxEMxMNcBwtwThkGyEojg
r7KfMcOzzSPNzrkNFCcvgJjY07/gs7T+6ytU+zm1UNJhV7mpNEqiAXnexHHI2rlx
ebGWW+Zl73IhoMxycOK+3kU6vArxjKpH8V3TNL7YUWcDHgGAFZYvRftuGrEfoE1q
WWyzykKnGtax+7XeeeW+dB9hXHL6OCQWkYQf9FoRWLlKWYJCB1L9yqOzPJE5836t
gim/sNzojACW/6ROexG2roYgz+SOdxG4SVswhs/zcml34vJCrTGLaqBRy0CZdBP5
0eWq5EEGVtxfaqtncMW5RhY5Iu3E9qWN3y18eY+Nh3Fc3J3QrZpLTMtFOe6gOe7s
nc+VRoqmMC6DvT1igrproTZRNS6vSo1rBe5DHB0q3T223nlPhhncEHFdf0/9z/nB
kD0KZMYavXWfD/r1Uk4qNAnW54RzJquMIpfVmT5T/xQFZMpKDCakWCbCfxkeHMpQ
Bfh2sYYRc+eh1v2ZnY2oXplAsrmhUzNNERFARehGpaI/DFuTg0mrrtzrSNTRdZiW
Cwi4Hdp1m0lGsfxZTXVQX2MAH9LsUlKpK4e/Qrdb7jM5dU3k5jdijlb/No9QrZwu
+KK6tphzVcFgIQl5SZe5hW8uSwX7ESmlDY855ZJvpjYHCnNWSFCjiyr2p8zbjwbn
Eq/1DhrsXiIxYCHu1ZZR6KfVOa9vRZ5ngM14JV0xtbvCpLiX6lIVmQr2wgjTMDQh
XDmW19trLLr7TLkjP+Ze8hrxxviRNIINRDIZkMwTuaRXdoFik2V7WpRb9qELl66t
d/mBQhys3/Gz0IzrOXaNb20jAeQ9klq3oBWPXc5NYZKDJfTGUYPnfyILrxMfxffR
WadR0a3iVmpq3QmdVeWlKzDpUp5sHXtSnFj9KgWUGr0ot6FnQOUdx+OfJjoTYO0H
2x7CyQ1YJg5R02zBzkoMVvYn0uLQPe3KQGWomGLOuoRPJyucGrbOuy+NSRy4A21f
mMYuy77EP1OC2L+X+yeVnYVe0A7/sfLO98bjZmjTCB6+dBhSPVK0vJvFBQqLa16J
VdRd/Hl/S5K/k6xtrMsAdCEV52KOf6TbIYy7YScsKQQn2mQth8aEyHo1TU18kOR1
twDd34CJ0xzI4297gltmTXm+M/nSCShNiKjCE27COgIo9GXiVt3zahJ0muSYgWeW
IBv7X9QRPD8G2s33Qx2GE+LSITV71OlTwiTNpMYvM1sovxUzDcxxl7ktAl2qCmuU
g6UqTcFlD2593+g3EDE6QN1dRatFoJdMCvwxaPst8uvMamkZIM1dD3aG/1xEV2/2
Vy8igUhCf49esDFz7H5YQLl2sClUYZJUNZcW1cRqdl1MC0Yg7dWHuH4ADuBbFAth
mVsT13GNkW2rlp6qbcKSvYIh4PHJMQfsETAf3Hg0DAq4AYYvboqZVNXcl+Xu2hWc
FxaD8wQBaUITM3QmDUpt07qJgti/NmLjUHmFaqBoYXQXSraQZof0CuSUwvxsP4a5
vqNS/vipsalNToWbK/c+EluDUt92qxOolSzCoJE1DT4fh8QOBXaOBwgbshW/umdI
0wqwtqYRjom3+pQx5JsCZCMtaZHZzSU4lbuF9Oj2JMFtbR6BuH67msuXAH0XxR3h
9j5irECyRBetjLTfYxXjOO08i1KXo3OkkfP5yO82YoIQcu7qAstwS2TK32aiJ4+E
twlDUu5wiowdGEwQHvsZf6lmAPfZ/6KTVxaPr1fLAO9R6TYcgE5Gspx3Q0+xTr1h
KFJSxRVsaEGH3cHUfaiXwYmDxq78cZtdlMKcwvvWX/NVOoyobB5/Jj+jOqggP4cN
ojygnWZ5hnv5oDYPIg0TzEbGiqnz9Rk7PKnaapEE/AdHHNCM2m8mbc6MXfsYKtzI
BkbC1TA8RpY3tkX2nZnigHHsSUSOH6YzQVBrO24URl0PU9x9N1aV9teX2rWovQSj
hH06NB71+KrimeWMT5cAZmBb0jBiyx7MbA2Ai/Dh9mayjKP7xZs6qQD8/WS/W6z3
EFSUFQW+Gib7iqP8c/55wMr7MIqWQJhz1K5akVAZs1EBo+b0ZPUyo6IKdkf/TPRI
YtB4PdZ6fBe+Z4GRM4TSqUlqc3eMHrx5p9s5FC71nCLlzAo1pvXXxMiVaPTyBjG1
QyVa72yMdtAbpyol+MkJ3HbhEimkpK96eaL/y0aBIjFg9biyfFNRE6h44AMbnnUy
HxeyWjbJO4TXOhfS+wSG27JAObBVnkEBnFTnC3M3FuHFpy7bJAF0ACXRjwW02B7n
vAbdwknlMujll1VrDpWil7ZwQhxHIsO5S25IR1dXuzPra+2m6BdY4zV0nk0HlVFc
u59PBTmQvpmWDWbHWzOrRvqJiRmhY4WqFK26L7aS3wU9a3SOYl8J4lOivOr2k0zn
TEc05jd1LPuiXmHy/je6HxqhmZb9FhXFE9LlQOoWkiUdZudQxtnS3fvAFqL15wd3
mshEdoWpMWGVOlkOL+x0a2MLbziBWDHdwVQbq33XlkWBltKS2TegRYPJFlRG/KxN
QS+/4xT8lgtXVJExZ9CR1PN/s+XubarE10kVFJq3eeVQ03WDtzpge3t3XqN9Kyhr
/pf5M6TGcKlLmNsZGhIXmGdErpmQrxbEAJccjP8g14JwpP5cFgoiA12H14yjz/gJ
SBGRH35cOWUnRWElEY7PAv4cmj66Xqv4pQoMUTVk1NqNU5hO16TD0VCoTyBlLt5g
S8TDpQ67+4AFRmTGXUO/QFzEqey7vkBFEdHeHKMNFBysDx6wwAHEnSOcLNyxDMz7
ghXSl2ueJZW3fMFnDLDqO53uCB9J+YYJiHu1wTxRFdLkeazeAKQarTfXGVTkB3EO
ibIOIT+8BSfuN4glF93pmGW+SHAR3PxPUNvqorVRpL5VnS9LM1PAUJxIHcuhP1TJ
1xbWCFpppx6vZLj/uIJb9qShkVcBJARFN5SDz2Lk/m+glDxC2tTrc4vQuYf7sONl
2VG6YoU1pupH1Nczns2TGztpEA6kII8ysHlFb3CIHA33XTL9uLkv+/jD0Qt89SwM
TQ3I9AYwaQf6OCnJG2KQ6MJUcL7jcaS/yBYuL1/asmcppOTU+QbURWtHNct/jENP
vzenfCP8LrLgl6P6stYF4llCJ+ykl8bCfUqcW8DJMtQYXwULG0W7zVMtFRh0sQMN
ESdNcarWNDHnAAJofpP5zrOCVk/dsz8dM1R0widXnNxFGDc81J7u/kpoVNj4ZJB9
sstK0oaiTq7OPIywKu2PCEgZ2UWJv7YSjBx8DtPC6Vp8Xha6ga5Y4R5Psi/F+vu3
YY2FrEKDRSn4CXec2txTqgrgT3nUk3CkV1Sn73iRetRR6mPpVR/AxrMJntWA0VZk
NJ6TQg8drmqJEnN8Jcj0yctBvTHNNyfhz557gUh3KBYWAG1E86iWBKGAjeSLqWe8
41r2XyD7o12J/VaxHHk39dPlv/txmnqUQeg6C2UkeWaz9N6xTXvVtgAvg9huknUV
mK4LMxhvoEwMS9wKocmDFCprKYo9xsDPu7un1Ok126c4VPLtvJrfhJR9Jn7LRRBB
pfKc5V3fIyCgMMdmFc9u3WKfz2dw3NOT5q5eV3w73YHQTXcannxmOIgy9QXpSVFv
CAm0DLMp3Cf9CcXoEoRqZSkjwborCx2Yzob0LDBfCD085zh5lV1e5F/ZveuOBnBl
A0H2JtlVelv1+6bp1cAbEmGPRiuRvlUXDE7ITc76YJwLAcOZDriEKw4z66kEKIPM
kSGAp+X6lqSojR3WjhW3cHvsuScjvUxN/NUsDb8kep2Xk1yxYliNWc9nwpDQfEJZ
BIsmrHjzqNTjSa/RQFRelPwiifJTdpHzpro3h8m256kgvppl/Pb+zdNhRKTMAVTJ
c/v3yyXjMdomjsTVqaTaNERV9zKjkIndr1NEzUu23tkg+foKOnaKS7Ysekf8T6k+
VKr3aXr+wTtzB0+HOSu9DWKSm2mkRTNwBj7qJZv39wCymowAj6nND1dcoCA0rNj4
Ber2H8k958yfQpSl3R+DCGSICel9K8dfXMVdr5W7fmqyLnEmKkn5OdrooHf6YEtc
169uVgp1SRt3p8+0gEU0MLfQfi6XychF8Wb31nYtRU7TUbe2RCyteGmzPw3VwvYo
HyPf8Xmd/nFVAoPqgLpTTx+tsbOW/coP5FlMZnOLVahyderQMemTecYx3v5/QXVn
JHLMt5Dh15ErBd3nC1qB8DP6JXWr90OtlDDdUxDb3/2ionLx4UKBZFm79EdVz+wE
AnAdDbPGv7VuP1FUaClAiKRCNIZMlktOPeHeTIwlDocf2ZEexFa0il5S88RNJDXb
Qmm+joruWiZCiVPXmA6C4yOihJUtsjlikfeNTrBsLhYcmDdQwQi+b53jRNen1dDU
NxXsOIObSbUqGzTeyp4Y0sCv9oP6o6YlMptO8s3312ORUwzla05YkIxF6uqRCxXc
EynvJU54lHgzhkAt58BI1PXb+S7m38sHjAvyiTwZonV+fZMIAQwlEITDyG/EkAmY
RLOCmGxjQuh7xQK5WUAXkMhZ6YOv3jDtbeczhiL3mOz4q6baYEJlfcUkkgT+SX8x
ZwM6LyfMU17y+m5nsQvWcE2NzYBb0N/DgiG7IwJrkzp7DR6uK1az4RSG2svX2vNY
YLbl5Dt9RecNIljU+JfPraEDkbh5IdpJmgc9mdK3kq2ITIqpHZd+Dp1fROWbKE5a
U7iL9KDKElGYthwt7ELC8kRKG9Rd2ZxZpm45NSTuzx7QGirE67nJI/kMvSYIcL2S
Ny2peQbuKWuaWNm+i6vukJ4lY4DqK90H84ut8iCSZe8BqQV19twc6sgcj60Vny00
bTnrnbwSkAK5ItcLkCfKGPJKXN9pHUDJV70/4wPmoKnuD9O/k+YyD73q28fApVkd
hmD29btWcxUi7P5ysrqvwhUE3nv5UZfXywbE6AMCwt2YRFaMGIJq5rptT4sCL1KZ
nb25Cn5X7fAbYlXR3sE9DbEG8Me8YyIzyeChAo98VcwxCt9wjsf3FF660D2eu9+h
weCtLUgEtKTsUIVbUfSwaHFkdRPSd1YiawgJOo7z3pPyR7VXuyMT8tLajwhsIN/f
opBNN/k18Orvk8XyTsuV9RSzVZQNEevN9c2LoDBcrTWHQVwF97csEYt+ZDfJghOI
xuhwHqt863s9cR61DHfUQMDaTF5ozcygaKGUbwefve6r9ODa1siuUBQNtOdkJxzE
VTmFWh3y7e80zR0TsWizZyJXjiS5SQvG4gmBIM78dreFVAZyEJu9E+Hs7l1KSvtE
rcjRlKdqOkJOGhSXKlRlX9VIyCrw00Z1rc+5tGe4TUw7iYCin3vaKryjvpqMgzNH
Q3FH0rtzzPE4/VUagXnf8PaPTYyIok5zJg919zb1i+e/SYxOiyqYRG9mRDfFujLT
2FlSpZXJ6oCYvnecw+0YLkUjkce2w7FAO1jdzaFmt84rIUmz6TMPaHEKrX1Q8NKl
95eJz8Wvd3tiVlqd+KW6wlax7MnHhonMm3cFCS/AlN6MfzwYgevBDUZLCf70HDjY
SF+24FLZeoXCZQGrOnC6pbWv5eySSSkS4mw0XNnxsASMwgUQZhtTs/VaN8/eaBqi
05ORnz+HjovFSS366sO/xD3VFsXn54JWrKnWl/q5h7FXitBdZ8CBhQCyWgoZsUR3
qBT7xBFt22audhp721ZHtllnlKGYTQRYVhJQrPpoj5Dc35e5tZPGY14tPABsxn3W
cGcLDXFCcVSPoBkAPzA5qVKTV7zk2/2/5KXPvXJKT/q14JEbP9fxDtZfV2ca0/n0
7R7mdoLxJI/zKQz1OCZtP0wYZJE2e2lZT7/qChLZojDgq21gigi5Q+3jole+AB3Q
T2RtaOUlj7ucUU4vWSzU7Wyx1NNGc/7HxQOfJSvElEmhQwQ3MceaJcmj22WTjnL3
kqSPB9bg3FTZnD9U6KIn/RlU5HaywsWpZwTtLvatE9bMAd5v8/y9G8MKMjYl85TA
fuYg54zh2xNvw3TamI96FMviDguXerp7tDasxE5iwC/OMuZCbNEEcw4r+8EDDv6w
DuFU7SuMxDGN2umOUaVIKvyhWsTifSnQHImREMcyLZFtHbl/+rOEnWcfmwahmqMR
Txb5wCVjAIObzzX7cZ6d53V9QryC07bY2Mps3KGqVSHsPmG0jsQJIPbbPtQvMNnH
4raYAP1xmOtXsDkP1JDSCrzVD/4o+5GrMsZtwvYT8C68TucrAtQvdi0lIMb8ME2e
CybvEdd12+GXsHLQZ9OkI0jkK2fSdg1mYvFH9/6OZ00Zx/xKPrXJnmWNq/XQj1mz
MR2uxMjoQyiIgOVtU0lxjTgkumUB7J0cRKu2Y5tDrfADeePhSYsrga9hdgaa/Mhd
BDe4YOADXXPTHNGqyB1jX477zv9gQ+BZt6Tz+8rACCDUJXhSifIOxPUaM9Affk9M
wyRdamhGG8jOkeUJ/D6F6wixcSwYG7EL9Q9I3+aPsVWuFKSWlD4KN40YpjdEY0og
ndbwNhAqtK+Ie56jg9W3Khr2fWTGs13cznyJzqciudGrebSep0q3a6N/2LXKeRsx
DflrW/jQC0cxIgmvDsdxERGt75InL/7LLwuf/0nGtJW0MSBhgXKiPA5zgmUlzRWZ
bV9h2h7uAvMM+3vNiFXRK0pIL3s2cEdNGj9jQB/u9KqIpF1h4xaA+BLrIQDpc5Nk
m3wxrgw0vOdMo6sk5Cu01huHUWyuV2VvRFQ3fmHJv0pzPjI3KtnaGxgOxQBeI2+E
c3aJZXQbCbxie90l237Zmnp+Dozw5Y7FJV9okGJxN6lnaBpI9JsdU7KjBTxwL40W
cyYVjkNWhdFYMxtr55QK3LDfz8tgtX9qPiEk7+5t3/22rVx5/sMaD6ac1/RkaDvA
2db3h0Asn8RxeOoCe56+G45ZGEtEeK/UDQkPuWUi5V0=
`protect END_PROTECTED
