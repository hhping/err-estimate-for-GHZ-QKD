`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4KVOTl/jC5vsJce086+L7+or6YDSZ9qTv+EnJUO6KxsA2+7fGY/R2Cjj0rcFEK8m
+zh2SncDIMTOyYlVe4CZ7YNTyMvVaX10FR/SOqWlNMVmT4OtUsf+rnm1xH7eZixX
L7RejUlwQ14moSn27n0HOAoYFCmS52Zs4H8W9DQ8/rpKh+ash5uSG7jfM/voz1+q
J01hGB4yjJkBXx5DCMKtfeFAtYrxdxx/d+SOrNm/XfFxgUwpPoNabuNtUEA61SeC
eTxZuEUoKN2lzKbU07uP7+iP07oBLBj4kJIBkutBtq77UoPxTTSuXEMEIGvY9jlS
n6xLf6eSijM41WnVQJMplFeyCrA8G0CH6vbpHuT25YQAeKTKQNDLRN690pPig1O+
VlE8gt/RsmvSDWCuwQ5+wka9CxM4UtCgUW1KbEIAbpcBNDznlBUEfdLRy2Jphpsy
HOZuRCVIJoIOdAef995HgMvFU4uqWIAPKUxBk2uOzz3gUHUv5Aj2S2L8m5u6tKEY
xXmjqqa1JyLr3QcmBrVcCD20iQ5YPN/otR/Fj6/AmgEdoQfSOrNQzu7gF/g4uzB0
CJDgL6MDZmLnRHEdpB9DeVdrz1YgoGPk6O+pnyt8Oa78ODM677TZPe5HfQSEL4m7
tYqJ7rCwKNXUS1LW0imjMDpYS4QPKTIrOObKJpuh4Y8jUUxzNzPXU0rEtJ5Lxsu8
lVt/2lKB85HOkXeXlN+n9L0uyGhBVahX643W8UvAZEeFjIfmdCKsFDomyWJigOi8
+mTpg7kUoN8fg2uADQQM/Ns3OdX6/XFFIaWPYyoaHmOqCW9DbN4MkSgR7cLrSEg0
1OzthSXWzbzFO3SGLiWw1VGdbow/U5YB8hYgM/wSJjzW0f5djMQpsqs4XQC6N07w
f4Boxu79/jkgzLZoBl/8NkgTUvGsY5uFUJnqWyg77vj+lBhIbX83d8IAc4weNW0S
VMym9h67LWNmamMwMTF9lMKRAWb+tjfR2MvPf1XSwlXDiTCxPjBZz6ScLyR3+jBU
iPngTMWvvQbLUE3jFVW+Ai0q+rVs0134IEdgqJcZ05eCKxYyJp2rqF8fj1AlDqB8
zqDvZOpdo2nYVwIPexx151at8d4DYXPWnVIMmXBryAtJunhHxJwJrKFY+bJXkjUm
/BlvcMtI10zOrH8tRcPE9ZjO4QoOWVpvVjXPJzhj3fw39fuGDnKE5d+ztHnt8HDA
/K3aSc7Nmis9ZNjJRY4G3qfgP77s46LKK7u35yAGLdrNIrktgiBejkbOHt5WKAQF
Br2JbWlvdL/NQ+qnQae2fiC2yjFcZ2Ikkply8NlTZLfD3NjQVGjtEzoqM1Rgf+Ef
mwirujevc/Um6QtbbyaDpxJkjwBUj7ORZkGc1QZPM6yLFv+TA5/f24OKS1RtEqj0
IQrrPOO7ZXXnNnS2nWdNSOtHd7KffsWuEzR1d7NMoAyQrZUZni9Gk3TKyjAfUbHZ
wrrbt6YxrodTvhqVLLyJVpLaURPaGsMOfbskXyJSgQTdrI8ICjXot0rvadpnlRLN
uATSjlQGigV1ql4AGEozKZzvHp6C3maB8c0pW6T5Af6cEBvkhhndoKINpXp9yxVh
8X4+9GD96fgPSW2iUMN7W/91olMnliaLaCtl1d3/48jFnJYm4h2llx01YjMTSOv3
YViiEqCWNCYlelRdOvUcld2pg41iA0o774lXQEodq6ybR6JRtLPHzSQdNhAJwk/B
Z8V7ejrruGRMO9QgGkATqcshTmyWbFX1b+l6mK7/cbHJeGYEkDrN8sCPdiUaPmYB
rBMvG8bTlYVMtNlvJdf1B2G6K4MkQgQz4lhexb6nsMZJz8A7e4F0k6BfXaMHjqyY
RJwAw0NJQKWx1YT99Tz4ks2CN/lHhYBU1RmjHfd6u19uMDOPBu7Zk4wXKpxKkl1G
`protect END_PROTECTED
