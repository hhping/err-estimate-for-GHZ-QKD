`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
arO4vpQw95Hc9SYXlTLBOgqeqZrw7hiVGeVjyDdrIGdfMGmxJ+WVYiQHo3ZTYXTx
ACESuc8mn99OyRbxDrC7Mo4NR1U79CPTIxoTUGgcRlxAtn76S7c+UC20WYRRnmxi
Roo452F+qDsuSEawlUCZ0r6fUWuCh2TOZBHZ4PySL9oa3sgzQw/pl8W3Im+JeQwt
W/DKq45NBJ8zj3caaI1mS5Dzyfz7qPJx7X4D/rnXv8lLhIfJyClRVfFFue9IZuI9
wprkBrjIjOY7cInYtJGmWFRJpneL5qfgYl3a74qbrJpmMSEPuxI4AWrzrZu49m32
JgKIl6GsdKug4Rs1NKBKiYxEAvtKheO7mWrTTEhLVpgFIB4RHiOYWPuY7k+HKxAe
YdA443PLlgKL2OKbG5N1aQ3yWdS/8t1ZK8zQPe33Lgofkvjnl/va04VciAcnFzZV
Lulq2trsRFu3XO7td5jipYmtUAK2cbpz67JminAGPnpVsP7S39/pOmSs5cnb9Wc3
H50hPwoYH2CqRJKugwpdjyioS1RkT2JRBhXAoSen9vDXcKT38iusRoqOFVrNAPkE
umSMztMh3tRs6o2pS7UbgxzsXw7hCsw9sXde3/p1K8DqBNze+eQ30ZUsac5GG0sW
tXimlP8AEYkGEjsEtHI7bdzsqTD9BxFZHl0nkUtZC26xOyHjwFecaXT1QR0s5XBg
honQ9xv7/dIegduqfIeBRptAGKaIIaNYMke1IOHEun41VsfaR+SGcZWJz9rEXVl0
1nFnPj0SCBGG6Ifu7C/JbQaMiPtxdiReeYJhdvHwjySZ1KZDB/KlD6G2Xde0o/+Q
/wIO01jiaEgBGng0DQLElsDDvvyGrwgYtCKo7o+HTjezbQHZpc7y6zk3i0FScJ2h
uFutYL/V/qzq4eSdu8sFjLEv0eZH+fJn879SQb7/LHI0dy3GwYZiTepjXsg+prKR
+8cBgX30WnSW6JQD/nALXEsG6O6EnmBHH6sGhcxz6Bh4Pk1DWCA7sGSWPTNh72hm
k2XRsfdbHMM9NZUAY2JjcfowH3EX0kE73nNh6ZSU118wwp/Yul+UOKjSAjk4Euwi
8ppCM4hL6LXrg9ISs4LUfIvk5iwQDbKAS+Y7WkxlhCspAFg1jHkKLAhxWWJ0NV5P
1+/rQYE1QtGo1aAOJ4bLBTb6+l976NgQAnCRSnBy37R8XE+Kg6shZfnMQc0m9srS
3r++Ni4IvrwuuoxlNuHtTPL043tJKBFgy9MZabQXtYU1UY9SM/KaIrXGd6+hu/J6
3KoTnPnIvYI6DCasS23A9DcAeYV6ZfPC+iCJARg+cgvRSbwixYY6Zl1v1xRSgDL2
3jLnPbCTu4RVun9azBJHFdsOZaEnirPFdekZ/SpeBTAfccDz0ZsN3fP8lWBljarI
tkcYZAuYndQotNWb1THplbxYD4rHj/zxzk2jzDujBi/e6crDiWhrdvmmRNds3LiU
HT9Ywyyd3O2UnaW+NKYHRLB34BBL61CHvRQma7Zq1zJhsBH6FoXyw6rgbpKUjSaP
JM6Ex/ZZg+sYBZ/0OWE2GHkrF48fJaOjLCjttg1bGaTMJA6uQvOpFvhvLNR6DEfx
0gCsKVCT4gn0Nk2cRuSxwAANJP3UK4GcOLb6IVeE4DTO4mq9WKRwLBx9ymLADC2G
+3Bu+4DQTTJX9nrbhQGE5C72fuPM7/ha+4NPUiMrHbggNUdx9KhiyOFC1mEXxLqZ
js/ywZ/cgeTwYEe0mXFxxQ==
`protect END_PROTECTED
