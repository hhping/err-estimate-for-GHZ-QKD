`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1zmurc+TRvD7TKQtRWX4KM+6QMqMD4ID/8hUL2sOMPfiIQWJf+1sv4tZC4l8wCKs
7z0GjB/0gxPB6JbZ/YrnFnZV9xI+nhpjemoiK6vhW/fiUgVCmvfv4tF25XlBkWXn
pqBVaQEH2H9jcxDgQLwY7h9Jp2Kx9l0vLH8oKE95f9CTDvxP3ZwALSbf42h73of9
dyUWEhqHhAYhYHaE1qBk4uYnNALQ3M4dzghr9SAPFtY61uJg/brUaGzs3XpZZM+P
pDiuImqGteHYEalZc+pmvWyzSexjF10xpMyujOljx1/FvnQFYUpGB9jVvdySLmUu
dDyYCJVUBg5/eMQP8HnmJrW4bKcdjcIp6WIoXBfmPW7GjiUfieQ94ga1goVWJXWF
8UNhx2dT4XssBOp7xLArtTa8KA/z0vFnabdMUbtvi1uCImHxAdxvETUNUjH44y81
c22KroEuxpZq2JxQqIkM61ivqDWessNsEN/f61rnD4kTGxZTL52EsLlDTEOZdKYI
M4GHyd7JBl7T5Df0JUXa0V21L7qI/C+6pd6d031cb3Ri9zzDIJptKNy8Hm5T6XAC
44hH8rlTg1+RQq4kJJKxqEapAsOfh4289P3q2lhMT0DFgzBbbMt5whw6v1F9aenO
gmTzevngRnfmhi+zpfAnX171COR5pAgH5xjQDNmWvjXWkVLfgCwIc4+Da83/3h3f
1XEE60Uvb28WtMHCX200rX4BNfbFwG8EAwR2gm0flWBPLhX2J9tJQ92I/rKGFx61
ksTPt5V5qged+Anpao0mKN5ByJLI3I3mWLocEomXtmQIdc9+k8GQa+N3ewqPKUXv
HW+uG9TxXn7flM9jmsh+TkHkwBezdn7CAaAZTkMOCUxKjCwWHCpoQTLudQi6lNV1
/4HfKTXZGsCzXWhGjsfJFGShBxtYXC8fY2ThfKqEAVpZTLSwU2R1YizUwpWkUDkN
Hc5nCXW5q5gK9tgYcC+ShIuS0xdOAlPS0Lqt2EvHJPIsfUjwIanCNW1UK69tDnLQ
QaWKd+KkdWkjvUdsC00XHpUoUoRcIudBEOno0y4nMjDrftIii13hLLx2bwFkDmUw
WayRMHoTAB1jbvCrMWNgZ3WPBrCHbQp1iNIBNJg839g/yqFQxia+gimZc0Dw+4/q
wEoiFSRd5oEYkEVCOyb1YQqmr5p99KIpcCOiC5FKif51TmtkCZrl2lGU0MrLSXAj
mjm1xZiBFbvB1vmoQGVnZMAcivK2nED2O+9QDmThMLmxmI9/CDA8X64yPwnPzkwn
iVjIKvgWEwHLqpiOUxad84hH2jsHAFTRk7MuT9vswitr1T45tFbq52mpu9tjHV5g
zlg8cWwDZSy4pfUvzkN3vW+rsL1RRzjzSCriFNiERXQ2EyIVPpJV+Ijuehu2sTdL
NUrvemtrMEQMh3qg/+lLCati5qrciPRJklzo4vj3LGD95PshzBWkHmpr64GAK91G
gGL7pAbAQb8QwCLICzI9jj8F763Orc8RNj0hViHkjgCAbge3og3bXF2lszjtc/Eu
z4KLAx3XZKP/xOA2DHm/1QpUnApbJ5VJUJqKWjh27bOzGSPMEzQTWRfBhJgkLnwL
TSxQZhlbcluV35Anl8sIRyLAsMX14aKiqepxa7VpVZv8I3zAHNz22VSrK4GWtr0K
sKnywjh6yRXd1ac88DXN7NXzTxGoo7Tt5TJN/ZL3CtkFs+OzwxpLYhbZRXpNyoXY
9tZh9gJaNkMEoxbIVwuGOb/Z/AjFQhvo7NvGvt+Oaok7ip0OTqfke9G9QZ3l1fL6
fYqXFz/KeMD410hz2UPJvx4+f6827KSKzmAKyeF0xAriE+TGufuStu1elsn8iiKE
/T9Srxb5KPjWA9eAoL4qCaLj0Ls0+M7tsomkdcfIU7+/Oj8oTAq42vIAC7EHZhMY
x+0wOZVd1hWXiQBsYXSUsA==
`protect END_PROTECTED
