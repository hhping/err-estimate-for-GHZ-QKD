`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yb3DjDCRgm6gF1b7015PokeysawSbASrDx9BTZ17T440zYBEgTRa0Wl5R0W35DHV
NEe5K0p/lyExsf6XaXyC1LCb6u0X7BarsZNV1L5FqUp8lnG9XwdOWEThBCQ6ab2Z
rxRFzc7ZP6HYpdDNkxeyCwRJlQJF2uKmPPLoYSx5RKqy5FoRk/XeaMjTVM1eQkCK
qbrsp4pyXWu8NMyGHzSqEI04Q/VjbNVKy8a7yqLKkvQllyDkWapo8dW5qdCR7Hx9
7a3atcRiwMymgFVJQGhGnxhWcFDCj5E+kC+FaQdXiXgiQ7zJORY0yOoTB+ToiCLf
T1cOOuXDQDw/P8e0d5krE0A+w/Gst5kRBNycCter4kCXkS6D3XB/z7tFSSPylZfh
gJZbTpMgJxofjO2BUjKJKaM/8OkD1GgAAkYYdqXahb5pVJi0WGi1Jesv0ndvl3N/
ldDHeSj4FTJdu1oWObr6d8HJptc8Hr2v11cAmmgEobAl1SWrkje0zXRQyYdfTjLN
jIh0ngWdh4LY8e+eZ9nTHWpQg08i3r3UaQ01eaJWMUY9zdhLmb0A+yZBe5tlgc6L
CNn2IMtAFuHqlP3+0lM3osbDVVi79oUjCFthWd2N4IwrDobWM9hVKnOYCMAE/Dhl
c4++sfDwfmuUQK4pJKSYKyaBStK4yi3LxtG1OShlwBla8kdxjoNaSKvxp1OyugD9
F7kId6klL/SqVlyPUnev0fHiLuYte6hTQrpUiCFmQOigVheTv1SS1oLxuSNe+8db
2ikL8XKBt+bm9yxgCfiNEOoiBIVhisnjR0DHGRy4v7CofOuO5rX75BtjCJ5tcIxZ
T/rUs4r0r15o6kMKvGu0TF9Aj5990iz8Cm2lFqwyNAZqIs6ul+n5wCtXh58GGo06
XD5hyUrr3SfjInt944G5lj3lb/A57sVLB88PywjyJouILnHFCUNhaXD7dTKqLU6R
plXMnfzAJT82ebeTcvl6HunCA8dHZogpiG4BLZPwWf7wr0ayjVSw4Q1JmbczUuVx
XBVZ13QHtjbsEF/JAjgB1oN5XvkwkCuLNJNsSjcNe5Cr3oxqtneEkAcYWPC3KRfc
H7qLthVsy7DJCNSC+Z6OgRJIjN/nDDIVeZCJysNzitBtRmRw47XWJDF5ZBu/DaHn
RcUozzPJ/LDFxmBpfFMNd8dtHPX59hNKPNLfj0WmHANFQwMn/bDrRy8IovAkGLcc
tMc4PR1v+oLGm552QLJlk6OHtB3HH8dv+WNl7uOQf4nYh+7AI66l55JilhQdFflT
nYbvYyPR8kzyfixdG2DAOmj4j5pv60HEvHfe9okEKydnLAvLRiSeH1Vvl1pilRnf
6o1fsqW5c/K1C3JUcOSwlJDZvvsxhTLvhMTKwK0vF0f1tBRTESKF6gYY2t5CJEM4
CpeFHKFnIqn00ZQrHHteg7rzr2kQFniwBjvESLd0bTVgLIzJwBjAFu2Ugsvz1aNo
h0xaW3+LD+YEJpg9LOUA/4RAUQ0bKQpT+lwijzwednbpSWCBm5uKtSrBkMx23ADi
jx8b3XhpbYQ0wzEuTKbmYmVOe1E2UmXVHgV3F9cl74+ifaVxbo/1jZQ4M+PSRcrF
9EmcEwKW/WftD9Z+0s7THp/IP2iSNZZEiHp0Tm2yQMKoTTEnYQFjcI4UQvOlIdNT
GFCMW37KwKs4cHVdDsPnn01XJyv3RJRpPl0E/XfrJzz7pwow/WQFO4F0hwf/JxQX
Ff31Yuk1m+hCOnwmiGLG5pOssojg7B0AfG7JJ59ZKsjZOVw3XMeiHPWyZDbedJ1H
omeMm+Gkf7Pg57ulJ74HtYQFTmmLy0ZuHI6RwFWwHMCb8MWytlFaScxd5pQmBOVs
mNJyvICcpj5X/U1+KO27kJ/46Vl28c8Ky9MsjTcOzj7qA3Ru/6kGGguuOgIeLJN/
KK9MVYasyzHYOHdMD3EByAHZFoyQbtE/YlH0d4lusHAedX+bEZnKTaNIealDccNE
i+Wl7Lvm9013CpgPl15t6g==
`protect END_PROTECTED
