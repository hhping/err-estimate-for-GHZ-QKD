`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oha02FGwox9IPEJ09SKBVieMxOQNvNebbrvqleORdj1Qit1GYLMzcBaVZVpcslaa
yDEyV3nR9CphTGEzNEeylyBgDYjHO+7lC8xKAwMBHrtdbeer6e0ntMyYywDuJPO+
EovShr2lP5PhAxTgtG/TrGGACAX4h7iCgDvNRvA6oa2APQ6/Yp1UqMTcfS1bi49u
/WbIOlTDajtdI5l7Neb4DXbAKzyNya2Ao3KiY5m4qbEw6gLYhAHUZ6v+dTMfEQB5
SJr1CeuTR5nSHh+jQAtTTlLj3vHwzBDQBfFW0Fs0nZE5gmMpsHdT3/ODlx4ef0st
hBPCmdjIwSNhNjo7QkNESeSejULfr5Zpl3Fp0j+b+B/5d5RQLinhQjDpJPKJZOW5
cbLfOewFrsPi5/33bA9j1MAlbL27BCtIHP1Qpt5S0ByuBfdjSJmJofAzNXgLfzed
xKa/NaKLFv2+LoIee0YVP5UuxQ4gOtzNf+EqKWpytZGRAEchdLtK0Ld5Y+Xnt0WD
jjFuTpRon3k6YCcbw/ZJXrhdkL7X6x/uM5xL2D0n+4G4i1G3B52FprVv4GXHOWi6
6aQTaA0nkJs5B5DR/UVoaqQdBBo79WTIhKT9tGFpiqY6EqQK+69PPMNkdJBIx+qT
791DvCJv1dcVVaJz8e1ylAuE7M/AHDuIbSHlzbHhIwN6NdkDyQUWC2cZN2PqvO/7
IYZqCUBWugzVmMAyY8JnTUPFl5P3BoccFAirUiddl9u1Em4XK2dI+8kpBRnBilvm
WbC2/79un38/U4Pv8sPItxGmj9Dw0bBF1AWS6xIauQWocRKERFSOL1byHyHwK6YY
KVWSaSaUofpdiXXuV4WBz3bJApaodZeUOMvBhiEECTON5lbdh67jyIRtj4RvdD3t
Lti21S0G7uDEaWY7aLjHZIn9mB1qwBaV9fNz6Kus86Hk5IRcQOsvGhHtZ9d4r7W9
0gCvFVJNK1KFqUB8nocHL/mR1vmnUN2Tb0+nf9zi6eKaIXWZSWTZHiUtqJOZLA0z
FbdATxylgRGw0rtTeEdcOAsM7VwDcaSD6wZb98NbC1Z/AXi2BIJ7gjfWw99thzrP
z1oiFfQKPK/LQImQQVKas+JZLJtL6m8QlVIRb1cwq6rAsZsdWyPQTUukNMQc5yWs
M3x+iIgQbx8k42/AmakwxrttshhlSB0m5ACrd0RokwihJamO2sPyYTdwsZ/eD/WN
RjOKzeLlwmUk4/QHjSMJBEjOCeskMBs51XLdV13VFKIJAUWju/jL8Rh2HDY2bGk4
yznezPp6BfORk+hkmLEPWIfhjHypW2NA6zqkzxYG1KbXXfihhi8GrqSZi9oMhgwD
PoURrN/KroJzox7NIY9y5M5n5mk0xHP1Ds6wlRh8Ml70QqzL4vd9pCtd+kV7U6H+
q3tgcolOSurUiKVR5thaFQ0xoINELVAy1PGwTEpxhTU+RxFQvXHzHIy5Yvu7tovE
8EMeBPAH66Sq4FJ8xQV/WELG3ZsjorcU5PXh+9VJ+wc3M3ggoPA1DL0Y1aKL6SQH
lIUwH6Mf66UegCRVJbhQYBV0Uhab02yg8UkyDV/J2gD3yjPaag6jDQErLZXUpA7f
X9NppAH7yuTtbazmhHfh33C6A0N2qFTzl4wrOW7yYjACxmwcyHguYHFQeUfRU+Ur
UccFVe/Is//wt79/J/7Tino+j9s3VL42xax6iuqHTWUHZgc15Xqtzwxslcioc2Gk
IUKc1jo2K5yg62XoMhyrPO6LPzYTApWyxJ4leiuxbxhYSrYV2ssyGAVF3fIvDLjn
BVJ4Gj2ZmZ9qHLAq9i69pkRj+k6mNyiwIMhDtmNHtKXeDBaP5L94cNx/4+v79F8E
lFWWLUSTGXLKyJZ7HGCq11oS9afCpNQoBlktiBYsmNR8ip860B2yx1dEI18a5y/j
CCTAX6zWof6wU+AdrL8P+N7u1JS5u7j0PeFh1w2qyYyZ/sJ1gaOyQ8k39efjrbYf
9gN2fOg0eD0KP4KbgGl24g8Umq+C/bLssFj0OXgCkJzoPkC34pgFCQtUKGX5R4WR
15C6UwD5IhAEs9BM+8uUxjdw8RsBc3e57c+5IlaGukY0TiQ45Nt5C4Q1psye4JAe
KSQO5naCMZ5zvP5eEO06sOrTcHqKk5pzYZ68tskS/BQT13RCxaQCHWedFoATYQBc
2V5GIY827kO9RUYCr9sN81Vqze5PdwJeZl2Sh7muTO7JRLaxneXi8Hm8pbE8JZN9
5p9IMjLOvkOGFzg8kjPKNI1dV1zjPeFK8EX7EoAlw0QpLFueuWEZdAs1zJyBG5Mz
fOF8+g36soLDJ+7m1NHtvQEUm9XddjuWd0wpBBMfed2U80HyZ2S3yAh70ZeX53Z9
Hxa22sOAc2f93gZr4SG51bZnZvTi5v0SC4ZMabFx5X7eYE887N+MtxUe4HPfKbGN
ZAWcB1evXvNVsA0oAd1qx9YIXK+3E9I5jrAvOxrcTmejXbisnGOxRF8DJPiJn1nn
FaR+DGXifGd09mJhOIYTWm/SXOqG7glm0YdsJIeTvwGNdZn1GNj7UkxPTYhL0YiG
FuOkGYAgxUnIK1j29UGNaCy2EapjDWYl3JbQEgNj0p3zM7lKKmCWSu/HAEYsj309
xl2k6SSU/NIbpm1RSN+zrTb4JAzO1vdSEvzqUPC1sZBVhMNGzPTfnKjFlTtpmi/8
pRE6iLQgmV1CA7CS9A1O8MDSJ+7KWgGTugxQfPSLkQJelr+2fn37gt+NdDyrUo1B
jwE98HFE79CF5nBS0KwHfbcVA2FtoD5MNlfxCo/OR39Z88j8h2ZtzhINGEZXeQ8M
Vp67lZgSx4qcJfrOvbANxEQ2JVVH8unm+d+ANkXxSJl451yorRyKFFUv3VoYpR6C
gsjDACsL4d/yotZ5N7Gkxgzd1XUhYYQymRgbcWIWHLaodm1z+gqQUM7kHOAdjKts
dDVt1E5Tr3WxdCE/J7c8umWyMQLCMr04xOHceCn1+cIRloZOua6luW95pIfLfMXf
pRuC81Fdh/3iH+hknK2FilkAc7yiiK2LUs5o4Bvc7YuiIVv5DvyrfEAG0gNgbv5P
EfsxaG/oOSJT2oORPAIMNDmSciDVrgv+bAJ4ki3hdCzfhQnbDKA3KSUUSes5DkkZ
XvHIhAhoA1khFNWKlBL8SHLDhdSBQnwpijIiuYtXYcHcPGuIWHjrCFvJyN1RORpk
+s3U6chGGqKpO9G6aLnVrIfvP8QsW4JoPdMkgg8q36R9ZN2nLYm1GvNiCEhWKAKu
/ya9cmnB3k7ULSUofdSfh6qz9y/y9CMBHR5q5iCxbBKmorW0AoENDmCtN02lzNoW
ANZtlT82Tgv4qQN5+FKhmZle32G37XUi0JaPYyA6KMWI7J6af2U2FzWZAqrzpb70
KLvQML9TdCpq3dRmLvoFz/I4CKKoCaQEF69zE36hnVUZbImzzhLY7PCJGdAmb4Y7
dZdIa2PW7FJ6eGtK3hQgR8KOguYVzcEEKG3p/7cc5KcwyLVvxg7juIaqSOF6rBDg
18TNI1YmLcx2T4db3caGWTZcxcYGvQ7Ga0WiPteeCsDYZCCWoe6fspzJP7iutrVN
e4S3elp5Cj3eM+mCvdZMY8Zo0/Pd3qhkEg4o9cfBm5Wgu6vXcqtCVQWOvucHU2lV
JOLAp9kpbqYt/oZ1yzNnnInhdtpis28kNXGLY0kpQsHqHQUFD6muAqz2v39u193p
wAK4LdAMqUkUgdZITheMwK9ZX1eR9Aswnh43RwwJnDkVUXSl29+VEmtKKtq9a/w/
maHlsSjG/H5eBJ1ix7Z1CaH5S9x923+/tnBWuo9Ez4Wl3M97t4eWn+k35YoPb6xz
1q+KxQDjmPKLYkHrKWJt+qwOR5NfUtfr7OrQfEXgB/PAnci75Sg/hsaKoHYO1EUU
YMW7Jm6jboaJVaktH/D9Dh5vRcqHDTEjexGHjz2bLnDjyCRpP9zenrLp+BUBp/io
XHS3CAvTjT32JgvhZiUnWVQmIFYzvNqIZnOclE5paQs4rCwYgytEygofj4pal/Yo
ZJ77VAyB83mAcRdnAPh+hvtKqdfGMWIIbjGtIEK/6QDKlxyB265le/8PnBm04TId
NYBkDvBAv415zIzReLpm0A3DQoCrd4u/lg3kc/ZNv+Il8WPqlvhluvt1CuOPDnNg
gk8hAJMI8l1l8Fxp9vEUiI8zOfm3cxtSmNPf5iWbbYhDklOepelPfOienqt0Ks7p
ul5yAUhY3ofKTZsxVjNpmRiwLX/zaMZZaacjkTYLiIFk1KBOwCVAWbGi4n6RvvcI
zjocbpmFhazAA+IHPKhvynoSrsJ53E5CAVHV63tHPL4rrV1VNDGrHVPvCwmUp4IM
N8zzqmZftN5dQ2xUQPT9LbFarFKOFZb17S8i35+zdxL3ynm3o/3j7tZv0do8mUrP
QqNF+PnRjcebHq2AlU5lq4EcE/CVKYgW7zLUN2uMUJ1vUBDKghyVlEstFR/JX+mc
fb7LDeMr3QjxZAfU/EBoFhwrTgFt5g11cZDJH5Dfufl+OvSicNbv9DFvo2tan+nT
S8QFnnEo0Qx+fWBz3tTLuzsN3NIUZ0xAi1aJLHLgXJEMWjNaEZAjibj+WutX27NW
TqbzbU9Y1nprzfskD4MBqYU/cBxoEJ6VKmv1m6NvCr3TgzoQ8/GiRNbK2t4yeNmL
7R5+aJ/kIg7M8gzWLpUJOvpoPatS407B/RX1ae6ml9iEhU6hYjSRgiNciELpjrrA
F1z1mKzcY4ozvw8/tSSGqfrFMgkvkO+9r0LHMnIA7MFjshsouuDdoYa33htF+z9G
6gB0vcOJ+6eW1ll6dbvMIhULQVN2y5Yn74DtaLzgrbbXaJPqhThPo9lZKSFqRxPj
9lA5RAb53/AW6lmAEba8OqIECL5xkjeHuzC5OUeMeo3G3WrKY1iSSX7WQ90I9GzJ
bpWzDlBYXu/MdcxJhjPrMD3v1Z6uB8NHFq2pOcJMfO4KtCLoFURHcc6Y/7L08WeM
thLCX9S1Ef9pwqQqGEPci+Tw2aPKq7a5r3Cjf8dDCRjhG/FzXJ7A1AdELjhN+0HS
kg+t5gopHRe03Fl4Ez4+9bVKYPqEAuohBxm1Ye7h/1tL7i2BkhMEnUvIb1WIx4hg
HUQ1pU+DIBi9QIiE5vffB73je/mk20/qT0Cy7gImiFbtr/JJiY0oAe4Z50Dc+tRl
Ns+UgqARddIf689lbKunTPmER6N9cZoUQ6wLJwcLUAwKRot5r4topehR0P3jubt9
6uQZJ1R6875UQD42tZTL0zuWHTsHnEmrtYTadFby7f/DRp7AbbnqZBzEqU9mr5sL
0FmR3rY6YI0CSvGEp/FFrw+G7iQt2cKphVRN3/kxBT+d4cz1EyXakZTDwrbAk9kU
rwJcdbDcBqGikCacMqkvPZu8a3DY8UX1NqiSAEyN0NPOkAwl6dV5581xnzWGVf/h
8+ksjIDcZR3E44qfuyMT/8VVu9o7GN0Xjlvg20RRjW4AvaMwc3o442oZOPUfkDsW
O+DfG2/mhoWM5WsCi3Zes1cyuKBrbzZ5Wf+leWMMIYDrJUw9V2AMQvsGO+ReKOb+
R56Z7QebxztSOJw55EvwQwbTQsFVQgaU7j6YQNrM/GJr8chpskYEZ0suCPAW294Q
M+C3zMWW6gozbqz3AsdYNXylDjwJ35RiqEk2F1iJ7g4l0dKcYR+0moatZl7PURMh
5fuQnXoHrOCE/D/ThfIAflRKBeKh4zEaGe1gqDNmEPg+hp+SAlC/Ab+qCutzVsx4
BFF7gTlz8QdUkW3Ho7pDkWgF5YVNsvyJlY2LI5gHhD9fmsOILmZPCyBMg+vKakos
+rmTiz+ac/z5IQYZ/4kaNHZdHfyr3plZD5UjEEuuGh5cY37j7a1XHIitt9ijoOLl
zxXRa4P1NjywQi0dTqOqRz8GkOb2jJJ1cdTGU0Z6WI0=
`protect END_PROTECTED
