`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U/wvJYtz7yqcM32ta5hlXiQXSoXdJg76gBpn20YCIhJUEFgQzVxoMqwHUHpynL8/
tuaTlyY7AF644vvxPHBND1/n0/N6UDY7YVDQQ7ILzP9pvhVgNmLrWjD9psyO3vjH
TdjvQREFwfGB29/DyvuAjvS3+0rLpY+DjAw7KmgRkp1NmUydWSyHY17P94YD/Eh4
xOxAFOKxh4uqaSwcLUaPRm8N1Bqm/+dJTyqY29r/SozjOwcH9ImLVYpDNGGfpEA5
bo5hDeNWXlPHe/CC3888tNuXMrXDS96mYb28Y1OsACtmqpdWtMDzDXTmyeEV4b32
w/eibW82TveL6vryU8iwV5sBapR+8s3bUskfSc/m/PdqdHJBZZNjykTlfMpFxJAI
KAW/KySyBUmuwNpn4LS/Foy+80S+OnBgMevQ4hWk/C+0ZWXYvxo7i9W+owaMtJkz
fIT6uxu7AgeyDDR2HVz54Sn/IVO0FHkeHuKmKWY4PfQLkQV9HbHyl4o+yHN6xbH1
XBuUIE3NpGLjqDpJK8xWnTRqVfh/ckTa4k3Ydds+Q6i9nkKLBjz3RaqBMNz4EHEI
6d/C2dsatej1dHpQfgVztEbokG6u+L++k922Fxx+jtZQ728AXc9kqfGJzzX9YIfJ
RGLzVLNwjETwYaGsQ/k382RwdAbp9mro7iOivvka3xTjsbxqKgny2WOBz7ZwZvhH
vsLh9GszVlbbA1i56dxFteNYSeGD2sgM95FDMkq1CiFvsvJhjtMoAoxZxav0k529
dlaDC3dFhDSBWtPbMz/GF/4qs48jru0W765dPS9w+C6Xoptnh3X6N4hZtLnIBK31
Tp3eKK2Nbh1xSOhh4VTFBZ5PC7LgwKahUCQ67BFAUapnYjmprEPZ2zlYmSfsGwCZ
13Ug0XOfU1rN9Aj0wNIhc1SZW3iT3qCCMgu40LJT1NuQJMvxoJ0O6/mAopsFKivE
HUEpIZlK5XHwN0DWz0YvehBPLKsRLZnYRLp9FBUaJUzxOutzLdUNOlarrdQGdX0V
sRmR430ZumSt5TQJemnc5exqWG4zHYYI4jMXPyKg/NYEaloQ0ESasWLVfvxEDc8O
`protect END_PROTECTED
