`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KcPOY90pZVR5KxZAMWBxw/PZKRy6Kg0ADLvVj8+7Xix79pzqYGXTrpmjjdx+wfdE
MP84knJo2zVtzuCPiWrh36GCWZ5+U2ckrX/HWxhVR6pGXgRsqF+ymSKHZS/NvGwJ
RfbS5bkZL+6idoW5KLr+X97q0S14JtbHCu6Nf40eyMAnLSkGiGRoHVKgkGx7xlMu
1fETnQ+CneQDn6qW3JzGWaIe/SEGh1Wg78t5U9fLg7AAgDws6drbTzBE3Eth3/7W
PK7oLaPoc7nbWDfVFwrPwIiUEPx4FInd+gyGSFvoaZIzARa9fext2sqA/Vmqt1j1
ZW70/yoXOVUcdFob09zWboU9JEjo+gwP53dlWqX4KHOMI6sVXxNxTevU99ZoRdQN
usHIgtW8Diitt72H4CK4gLVJfqYr/Leic5RaqDObC3sQH02EOGltQcsCLUSQ/ydp
kjeWGF3RGqLSOG5of0M49ym+VMF0BVPON0nb2qI/C7C5eDfFop/2R781YYiGy7a7
wGCrZa2QBwCyutYDCxKUbngMBrXMqByJzteet7jdVL0LtJWXLm4XKyds1+t+mRhe
pD8z0lbkFRGBkHqgqrtEodAWjB+tJvHfpSBwXFUuaQZLcX0BOYpQ5KhC9mcPa3da
ymgAVHt63BuFaUPG8wiWIZlLRU6+Rc/ISAV6jCOy6n+3BDbuORdn2jozEehXNN2N
+YuH4Et2tUFWdm16p0NgVB8i/BBxC1KRowy4qwPJy+vIgjG9kjOg/amMhsXl9lRf
JKeo1mbKq3VvQGMvqrMYXVt2xWfnvVzSw9Ggr9GIKare9pLHi6p7U1HS7XIOY/hz
sLtKBVLcC71xgd3yqcyfs8rb0mREoEm5x8aO64SxkcAk/vS8Lk9/TdrpTSAEclNk
FhCtDId3t+OSEF9Rj7PSt/RR0SFrgO804UEhLebx18RqVgLUVkge5n0GMLUmJgt6
i5eayqmx6aMli5dzZ0sebgT7i6oQCPBqyGrIthJJNiMWv3PsJyefNxE4V0zBGhEj
5oUR/OgEBKe+wLYoWdHw1XmbEkbOWhFTjxI66pajPoTSyAtIlFwLhvd5z4D0uorG
X8pYkxeZBYmRv5pVEbpEl86eDCRz29Oj/hswlCXLjoytvAeQotBnsXAoOlhBRD6h
QF5Y5jIegqz2/UZAzhOmTKbKy1n/um1BJKI17pNJ99+J+XA+n4EUGBnLxAmeu0Rg
DEOdchDfGMHExW/ThLCGmJBy8xgJbhHKi5PWSgZv3Wk4sABzlzCgyT3nwvFqSXYh
ZqycGuQkZSjHgtKCIgt4I36VUtUu2nosgx4R+/lLa/xwK0Kv/FAf4dh0/knVx2iv
o08xjnjZ8Znj6Oqa2jpNl9H3w6oivIymQ9Izrh1THSGZEvQ4qxh2WUbx7p99IOtV
mRe5Tgmtoa8x1x8Evg0cXcZwGWZhV2sZNzMM0slN/DYX0q99dKoBEYuQlNIlxexc
VYA3SZ8WI3dvBSlEYW+3RrIcXaJf4957E3M6ix4BAxzNjw8RhGUunVvKZqtFPo57
pnGD2cqrcMl0kw0+T6bHdb3XJJntM8E388lEtH8FU7sMx0PX580H5+3wXn+W4O/s
4CADv6dQSt3b29X/+zXp3vcgsKYB3Zo1O4qQh3e5ESPgqw2IENZOSxG0EkAerPHe
nL21fU+6r34gQZXQGkfqs3iqiHB8QSJoezHmQ64R7rhG2vwtVaJvYsImBLLoY+D5
kLphtyaD+miq8+8/ETOwqCrw64AePQuTgqmWmHAsGa8aS4HEjk+fhX1yR4xD0/3u
`protect END_PROTECTED
