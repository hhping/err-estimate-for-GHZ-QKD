`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HmZ6kIGQZI6VeXszQomZLD0jHUq1lFdVeqPcyNJgQB5CuBMf4kMn6AiraLeBrcfC
ogI2S6DkwbnPbMvvpRmU17YCYySp97vkQT1DsrRkGs8fv+/GpxjCr5uXuYTB3yFu
G1m7bW6V0OykuCMltEil3/gVXBdYo6cqlJuhfEUC8GZRSINd+i1mFx6hJXsqJGKJ
XqnguwCJlXiebhtAEbXIGOGWiC79+XOSUDS4mS56S4sBbGlvqR+nLVoPzGR2VPiV
rNkM06mNvF5IAfHuRB7XQSyPu7qg3Bw5LmbNOcyEbkN4jHXgOhuV+gMgQwcZP/T+
khbRETXPH0WUg4cfvqR8/TCaSy4BXmZ69wlZT2mShPv1H9RotRS/Q128Vjj/B6bH
0f6uLaPcLh70qoIL4YRDXhxF4hGKAy9P4DwljgHsU2LabU8zXZ15nNX7D4MxiGUK
QK7hjO7yHnVIIWcbu32Uw53vtpwIRVhfpK5Hfo91KaQwwgzbmrq4bq9Vz4DSn9HK
6AQ1LXavqnl4r7nZb/reEg4YcFbTbCpM1DysAvlyUf8VjE/2FhKd+S9aekuoXkdV
xCqkNNjRkEbHSPquOGVxQA2eatgv1KQYIdAMBzyeTo5LV81Kraz/dFJg7sWK4O/Z
yqOWUom0edmOJpOdbB9+PzzYPBWUtHSNC0clfmSwlfmhziZC7bz+2sgW5DpXlT/f
WX9u6sTGr5BjyZNjFhkA550sGiCMwMuWWs7eO1FGB8AE5GDJgyLVgnzvv7MLK9bE
iHld9lyycTf9F2NMwI27pTG7qzGH6Awsv23ieyNDsdEtAAc6iBSBr5ctJOWY/GAi
KF+9yOXRAKnnGBMzKodevQUnIDIiJFd5gGVB+bu07JFRhPvLLEbkzohES3fcxodP
vi+v6iLJvX7jKjxg38woo08/0fd0yumlg9sXji2xWWiRMzRWqg89HvHQXdyODKmS
iFXS3irtxDHWGLQpMy3cu5HdYmXLEf+oc9S/GCckLWS+yjBFhit8EiVyFIq4QXO1
w4mX1ZdX3hdZbtehpYt3uE2FjgVNjdVOGhmergsrWk03r5jwIMNzd/0a7Yv5yI53
80z1Iz8chlH/uBvObBQWOmCHON0HI5kMEvo2A/HpZgceND4S0svVhIuhQjV/zn+I
oCgu0ymYPvJ/M6Qfd2knx+dzu9XRa35sxEgXHodf2oyUazO/iR66bfE0x777mOS6
VYiWb+ffSINghqyorhgbn+odBoPq1oN5oQuIccqtbTeyrmc3mA7SmZ77foZ0kyqd
uMQvOEkxeazXvQ4n2lrIdMQSuhXuE9q0t0hrtMgrFm8H83MRaLug+MtW+2NpCwrb
szfNmsvUp+u84QmiA3+zGiEbB6lpQP3EAlxUU1cg4P9KdnN5r3D0vO6kTHCSr7oK
yF5uHZXQMKEMW1/MHzN0gwKyVj5QYf1hZU+lgDWi3NBcqIamAVJYoM5GjH5UxzvV
mh7bZQzv4aERwPj9agE/v3JHeaD1fNj5GxrupmQmCQQHWLA3QWChlnRkCOFGMpn2
uunzJaXNPbtR+LXcq/7isJwLTEep75MjxoXI/J+UA2S+wHC808je5WmyZdSUCo3m
7+M+aSEf/YKvUHU6ate5xuCdZiBE1R1wihbTHlgbBbhO8pl2Nc+6FbmF+wcbuibP
M5q6eMJeBOPWRXlkpC8f4tCKBzAlsXPOSFdmPXCzeJRK+qiQQ8tNLnLG9eoSJTPe
tL8mrJRVw4RtWbCdKSaO/IlqXwFTBYem/JE6O4465ylpTO1Lh3ExZrM3VexQTaMV
3VCP9BLGnQsWPe45nuQcR1OxjgQ1Tnka3GEJ0Orxl1sLhPvCJ6ZYai2gr5l/+Sy5
FpwP3s3ZIjd8XyGEFkmwrVj0DkPkDy8bngfSNuZrkPc6uIPDt3mvDAUZCBoQaZn3
Ty53Mr2r3m6VcmpGZl2Vx+YT+Ejjyx2PhK0SR9i66sTx0T4SNyZiLJEk12eWYy+e
pym+F/5oUT55l6D3wbVIdj6CYGugTG8iwK3Ph5hmKV5+97sg7s4nXflAMZMBYHhi
h8R5DfwxBsbMj80XfP65JDd8CsUsGb1cU8C4kbI4LJosoK8ux0kM6kt1Jp7tTlhy
yhJmVqqwckSi+oZpi0K4sc2RyZh8nchLwrRAxmIxpkpnIXpPsgQ6u6/pZfkgZu4s
Cmz+ZOMUal4ohLg9zApBqQJ0nCCd0/biKKJaD1e1cJ7w5a39cG49+kE0CsIQ+afY
OhxnLmP4I3+n4zFsQbqtg09yI27OVfTrcVqoYjYi+R1INwNmfJf2n/LZ8OvsUif+
NCRtBa/bzIglUqEMOlcxYaypEzrC+ZTaJkoQ6rfv7pFzC/iSQeAuREQ4rwP0O3ux
TdmbrZ1gnGD+6dEkOCH38oe2xlT2idCBBbSQhAUFFLyCWlhcyhqI+Ve8o0e4mgSt
3WypluuqVSw6sx8AdxwYQ0wuFj6zQc0vMJ575lse1KlaFh20xuJIbo0m4k6jmyh9
/KqWZyJ351nPtNFuv0wlDDM65Uxaui1YbNsFzx8tWWHXXkQjUz+WjHMA+CUbis9K
W2txwFIvarub3TeI6V3PoW/vS7hcb7KmYw7v87tvgLY3uj+RxX66WWTtIqEg5MX0
mM+r5tsSk5tv75A2BSomqgJB8THHgAzuss19JkbzSgtaUPqZPp2u4/BAMmXo7ADJ
P97eYn6cNV/dQ2WEvAfPKb7fP/6mQpnqBJa09IclznFCFPS5l64LAFTE9hHAwMns
syMR3r2nDFNgcq1J9nnOheD2uUKBpTHgm4b5TIJ7JwFyGISfbqzRx6JpDPzFr7I4
IbdJPLHNgPD0EENhCTviNnMkns2Ttl+yIUpoC6urb2BpCx9cxjS1WQTOAZVrDMpB
R3s7LsRHs9DEPqvDn6ml/PGAuZKoZ0DQxId93ACDESf/36s0QTHTGurcuqv5VZzq
t84DO1kNZXAHDHYucA8mrrK2gZKj7+waB1Eo0yKzjzX3KEpdcIhckxB/2gB3aiay
wXHTl12kyFZZWaQlMQH5cBjUrizs3jjg+t72vb6BGIZeWvokpMI3w8Oh53SsfelP
VscmtrnRtvUMLfXYyzUfAAaKOiQYUGmOQDmYCsBNrgT0/S1S35WgDKQNQShzK7EC
EzhvdHxTEexF5bnPLf6s+N54WGaQPQm61LOyQ/o/nRB1ictDY5bnm3AqeQy3Hrus
HYVj+DoAe9RpcyAvpxuWoqeV+ZOS6BvTHk149pXLNuArU2MvOB6iyDs1nq3raFrZ
dn7TAA5oLcxb6UC8ItrHEFas8yVpxq7ye108tKIP6+sJCzl6eUMwaRfzU42hB9i4
Ts0KKIrFp87g+GfGiO9lUvUAuT8UvfvVIL9rnGNY51NhVm2Wept708fR/y7JdUOr
rWVuBASITmUGVzrZZWl/8zxrr/Ur+YLKEgFO9eKyvgKMGa8h/CmMiDkkhXgeEAiK
8OTidSzouDQs8eoe+nVcEznyqgEdwp2XyiarXH09BcadUYBEeuOvo+5ovbd5s5Ym
DNcujeacIqdrmeZhMeFCLKFT0C5Pj354+qkX9+00pVFbG5BiqHS7hfWy5VL1gF5f
bvfs/yCkNbauUzhNE6yqVEiKWhJP48x3zUGY1bR8y1k2oE9PqtfZNGxXz5yqyEMW
m2R4sarMgzmIWKRQs3MPzsD6VCofXvGrPWnEdEhC59z476t30i097In7TrndSZQM
G79EmJ5P4e9S503v4PFKiq4Ug1nPkZ2hbMJ4HMZ5j3b8fNEtXQj6kyUNz+RzmKdk
qa3KUqaoZwB3/EQLuyKVsKP+lPo7cbi7ITH+LYikPTplHBfLI6LuA+W5wsQoNyGt
zxG8VLKbsp2z455d1P2nxcQ6An5gppEku0kC0o7GgZiu/Br6VOd9dLt2U8GnvKU3
IZs6Jq5a+H186m4t2/9NJYhIyl5Iq1VHtgR9Ryv58SiA+7KIoTYODwXTzwhbkmF6
27OEpCT/iYYGT9VCwxnZYqm5LLQyW+758RI3fwfiiTIdjSsAPOMA5zeCAMQZBWT0
ELGa7Gm3VSwh8VuWVHZaLm4byt9vX7aMAP9b7AFu4RlXN9CarZACFUI3aHQ2cWAT
40dMGihUvCNEdmIfz8D3Ubd281RWKlC5D8JHXVvakxlG6qHhOZ4B6wiDk9ipXQX+
YTzBEo4GrAL/AVsG1rexbxuKBXlvt1zKr4qXab6IiTzHvq6EQL2Pdq8YNGp0+u1R
RjW6DMF6WmUzZXH6rJ2JS9Qn8Z5Fjx6xjSGrGDf7NjVaZ1RCyEnHVF2Y1Nox8aSP
v/KIQwl5dLa87AKF0RA0/D+dC3UoWDiPB7xtqSNBgPAy2LsS1vv2DkxESAOubEx9
JMECHxqlWSP3wIRCtu+kWxMtNe1guUzkXGVOPZ0OYCYkHYvAaVUxdBUopCeg9+xr
1y6ui5DWQ6ZDBEX3acc1ji56CKmxUUu24WJM+JO4Tj0IKfdfzDOaBe/nJDPI9RrO
Clcgl8ub166dizDFDlzk1dUBpKm86oeZafsrc1V/Rq91oEQFYEnQnBaVEPsc5Sua
PXwV5uZYINoZqpWW01kAQtTyNF60bWaePmu96ueUyDRM+Yjm3ghoin3rS0eePqoD
FlNSzYwhUOP5S+rHeAl7UceS5/iAgh+Y5JyE3RY8h3Igtw48yIPMxC5QCqZGMHJB
Q73YYuN6Rokq5lvqHxxz/cQmwYZvCyQlzZDZS8ZQ+LWuEb79qPenvdtlKsF1N1jY
oThr7G82yUzyX1floTzbbIwtiYfB+IzPPeUulGpbSAYyTZtQdZ1u84denvZ73bfL
vaadTsQwqqTd3hHXr976fsohYVLC/2ElFG6OQY+8qEi2krV9tNsiQk1p66XNyHYW
apKuvYm43iqki2+aX2LRm3Y+aTnvPcPZc9x0GvFhfXsZ4XCg2O0axThJiKU2rSlX
eXBATZAfjeF12rS+K7giAIWHNg+CWUbQm9BEceAlglSkOI9ZFdPck/aBl80UHHfk
0mwqYdr2jonWAkBhDlP3Ttf30EZEB55lPrbGXnmXZalBbJBJrnpmnpx5avIYSg+d
pphHejN1BGkaX+qpZc+FJ55X3LkWryF0+XSFPVUqhqLLtslorXPIMLQMg43EgWdE
5z2wHsUc+CT8rDKB4DQH0+qJnvrdDbEYSNHlgwmEPo/6bgAF/Ne2X/gM+WE1j5QE
3ybP1mpDj2pVdMLiAk/v6IIBPVTZpaiku6SK1EK+EzZ6r3PbL1ltXTftQ3uJGb31
jLDIBVrSgM1H+b1qs6aOPU97SPCiIEwgTVBVZXdoNiLYbuBgEkzA2kw/imjTVZw5
I09+OSdDV5xYx2LLN+uaVT9blZOg83jXQ5iKVc264z06djJCXS15iz780SXDNQco
NLS2kT6PDyYNiP0xR6ADHhnAJrD5Qlu5D8nVBiWUaffA8vy5BSTHWVKQPns82qpn
+vVwUqMdbbQJB6QZJkLh7wSaZaMmhBbKUQ7ZViixXwoaLGTKwQr5VfkUQ5fQIw3R
OGVoJBqCFmlaupOzih5ZXjqUD0fdoXstNifwd5K0D7VSD8Bx6QrMzmFEwfg1FCXR
fDbMvrr1DbGPpYhn4DPmWa/H1PSCB5BZfWp9+Rgy6pswyMDf0liPbtnH4KKiYrib
R5o+19l0pAEJnPW6gkbS1wNhAX3H3he2ajbV8z1U9OhjelH6tV2rQM7OB4yr08R3
iTLD+UhazLVEdL2qhrDGXgUzTkAnTTPEwhm6rC7PfFHSld13iThrjwA7IHWmHmP0
bxlDo1zBnf6u0hf7YBye47gKJHm6b2Ql34+ZXnDWe3CkO9lZzViartWnyUc+iN0p
Z6GVq8QcDylWHi138syUmy34/6W19gYO7wmXte9IvZEvOI1YjfgVB+BnRNJ2Etex
R0r3qDrJrev3t1H+2i8+4pMTU5QOS/6T1ODmIbAaPlFat1xn5Xy0PFbnGZWliZzj
rTPeqjO9HdLVZROgWLF2BX/UVlsN8c6fs2V1wYgiHVQ+Yar/UKBBzxr3hUforj8P
XzuLXL3zjJLCwT1PncQaW8z1xWubg8e3YYbhNdmz/NPIskALXby6IP3rIJJU6hHc
wuRm7CSEpkceG59yoltKDPmEblnEP43VGnAOqFZido1ZLXI18FOEoosaarnIeIFU
eslMb5j100J4F0Cm7vdvLAS7tZ8gCA2ywn8SqQAvrX+C8JeD/E7T2Hfkuf/O6ePG
Er0fVhvEARytM0JRHupSjJL1S985RkPdEJh8a3wGUvU7xguzQ0ikOH32YHIjncNd
/w2kWrhTA2BIEikPNBW1kMbXnAZ+rWQAP0yWDGqQOCdpDLycXY7Jus6gbwp1ulWH
XPKlzaSDvbvlvXsHoMeSI2UIwPStLXUR32hlRkUbKFo/NuJHFcKfULlSrp4SNfZ6
/JOKf9OD4EvJDVdpw6seSP741JsOWW1ZeQdMyUJTuokcRX2VL787kCMBwTZO4sdo
jfZbVVjjrws3BGKcyZCIJLo8X/49py/67Qfw6I4Vad0RU0GAweVKJtLsXC/HhNH9
beYK1eaXs/kBwrqjdydyPpR2Xcogpgt5vnPPzRDn5f1/SlI5xSo9XBLmxX+UrE4h
GM26ti8pA7Z434rH3YvEA+ZpxbQNtPIHF59ZBUBr5Y8l/PXJ5Gnw9yxkTtKQHJn/
4wSE6/vSrPBYVmlqRxPpDXV/bjXkOd4o4KJivrDEh6CrTJNgv+by7xdSmelJ63cZ
7A2RvSqfwgb57CmmsgUBBxE4EA2QhWkl1k03lLgAPsKWIRm+zfqTU37R54BtbbKR
qWcR0fuv1uL3VxMYIELXo95kVUv3OsKvrNqOoeYsLeU2ng5LQ9pISLKWG9VG3EhS
Wd5kNev1qZGSEQaJ3eU1jxTHuJlVLOtIJHLmXO3NbUpfYZvqP3YHmQl+3jfcvnka
IS1VWLJ+pcDR9yY+DqTr7+0p64n9I9DstTTxbEW3d3C7DRut1VwmoQmgrfYqKgFM
iH9SnhwuVdfN6Dj59V4FKjzp2y1F+Or5Oq5xlJXDTnMScVfpViFMJisc6gnYMdUi
ajDjL1rdOY8IY8VR2hQxO8YulEcvjeNWVF2Vib+eYEeyjU8S5emActxG7Zp0+a5Z
P+vn5/LT/v72BRLeP2XvuAoekG15aNqwnisHHkO11fQLsKUvRq0CvG7k3elvq76w
lALHeZ+yWSs7OGLTOVW2IxsKuLN+fHzrPNk6yefa8qKoHdQGhGqK8SzsBvE9ugJ+
mY5wISo/VgXu+cPN6o+tUqBKHDmsGexz5a25/WdUOWAPF+WeHyVghlb79zdCja//
/6ooDhv2z61Y6D9tbWM+6ELRkLyh36/vmG3I31iampLexj7I6ADj9R/znLREnVxX
Ct+WRvHHLRb9QLHQtooqYqEmq0lWVdBYmlrwCZ973qjIqtnFtig6YuJwL3gH7rqb
mXLZp4ya/lobW+Iiud6gvg1gnv9QvoYfkWMFKjRFgqNziR318WCFOn/mQqxjfICi
yQ/UcYNxvQi5rWGri2s4bjqyB3yGh4Udq7DWTEKV9XKo/KLv6JqU8BEZAj6BeUTQ
Y8BclKzE1aPTYGwUj3Xn3UXsBUkbrn0ZjCpAPDU7s6/GnXT9nR//2s7AYYvtxsjW
72s5VQxcyMdN7MQ/JN181qDw/ACCSy9SA4UbytMb4cLKnPiQKi/jkzuTrB88yAct
H+Is0FSxPMHZ3IIcx9+uhuasedp30BkHtclb/XgKFJi8immE1f1/euNnZdg2ycUc
v5KZOEjATcZyZVfcgNlKkOV5Z+Is7oVFkh7erMm+ytWfzH8q9klxANZDbIKSRuCf
mDiQ1rxdhncVIx6nUG6dk/c9H9W3Sctfo670Y5Pxd99/QoNtqNmkzLW9FMorrSo9
nMt0K5PH10TewPtbvwIpqyZqbkz/zFNjJaiFdhtwMorRIQKOVhzHUSOsk2ZgnXv0
TmmW7xlO9ur/iiji2ZsUoZG2yb8fevc8X4FXxg95Q87eOtHbUcCkHZezhtzX+lRY
ET1+p/dpxdMxq/x0ar6R6B/IEp27jlR3mPOONDABvSN1fXuMPdp+cg9mkvMNAlYl
scp9I55GuEFMM52plY5Zx51xuawJSjGeJ+LKzwfzll63bQZ+yo195YH3pKUShWdb
QpOt9IeuPUBSCtiOETfxkQvYdUjlA5Wtp+V5lDapryu1rP2svLOV9UBompqrRwvE
hoTn+cp5aorjLYIjm3p0Q7omT7YeRhD3e+QXTq7DyoPGKCfAeJrxuvMrZs+x5ejW
TSoz2fFz/sRRLc0xYYRd1m7fWxQKc7YrX/ylGCvbAJHNEmMvbgORgjBNGs4n4bJ+
qAw3NbFoCKuYFM5l0YIHACPkYXTwm+ZBiiMmJek8lBOM5y5OgBeIMEMyZq6kxm2o
QeNQaPsBeNKBRoAp2mFgPnoAWYJQIb6unfV+CO+Suizc4DXN351GS9V4lGqgvobH
MpFkiM107rZ4pbvNu/JpUG3b8PF1Pl8TkEaGGKRcpna7mVV65x1VZkKfAt9Q0G7f
xNEH2abYdBgnyJuQrrRi/2CLjkOoC9cBtN0jibTRA8jcZhujTrIEYJtlsAfRMKHP
gWKl+st2c0nuNZCOvzxvRKxGgI2OjLgMDY7hIMUB4iCUVdJz+fJ2u3UXO2OpJYc0
WUDXmuMDu1FLXEC2jGiNIEMMaY7fZSi/IGoCFkaNsqhJCZ2VlaSKhKPUGz4r2e60
6gliivmOU8YtZUw7o8rw9sSmX/QmX6ZLioDgCpnbeNl4JDGHEBcKrPYUMohgdV2x
3R4DsqVJsB6U0XINwowSNwMHLFMULq2ReqJ8M9pBGA4l+zV4Jlmo0n92nvQqS2gZ
qpZq0GIjTRcYBIvfPH4WdukYlGrlaKNgO6JhNDDUIWHoRvr80DcJg00jj8FyXa77
wtBKGVT5EsIf92/tgT7ws2y71NLEV+5v1Q0J38Ro49AGmEmrjRkNzTC9s9h9lsjT
GtXEBqfoWOuAhxKpzAM3cEUEORPl5j8EA213NStCXYJScWDRcoSM+2PckMwUMIfw
RebgkqWCq+u5IkXnlrLBFZ+0XXnY53p3wfBuSgHMiNgIc3erAANGbTLsALGfU6t7
pMTPizXeuUC1ugpcjr2WkCJxN51vgQFgEBImhHbEZX9GUJ/F882gnytCX8C5jlom
l5D/hvQBs6CGMGUNNNUEjqd9aLpU6rZSrabJYNBkkhqaOLYjUsUm31hw8TmqVdpb
IGo4T3zwol6RCV730GWaNz9ZB/HZHS/PLrwXlBjMoESYA1ZCPkt1hpLPyNfy9fN/
jUeYDv/KwqKMT5e8c+f6wY6QPrhjAmwh7dA9qyoocJoJq862oCoRHcEYVmDt2d1b
vDOFveyH45Rqs9JoDNcMq8Qqrl54OsodkelIDK+CV+ftmkghDg9RCOQnDTSOzZAm
PqaiGagXLbXV9b/L3sQasF3wfmp4/FkiTOQy7SPxTCN49MIzVFzX6finTmHx7xvz
ANrDc+k/SNx+4aXyJ8DYzKTAxevhXNktJ/DuoJTL4a5wXgGfCWSUeQbYN1UDLFLT
6/wyOgAjAHsDiE5yaJt2qaUHo6E1/anhCRqqm1iKmHyFUs3wg+SHFVl2JEsn+eNR
0qpFFNjruae1B2+suMHbQ0pNAMAlqgiwZXIOCqJzwiuTtAKhlW75WtfbcfSmbAxK
bpOUgKLWsjPznqFvHnt86UVwpu8YKtxbwKBsWfe6YIWyRYxLeQM5gkESmwe8ot18
jgvPtQHqFEYgQW5gEaIQvLk4T1QLQv/zwK4pYWA5zBM+j/hSEfaJHtF7b8hfKU0P
ZoxjrM+R3kjlh1PDq/8BD1FlJHClC5fwZrMEGew8HCmpwlZXRPTw2HMH09k/AjOv
n/DHIfbrvQtokz4Gt/Hp/P1C2XIwSvddXpnZh3bOWRazwRcB8Mw6fPuPkk2lvXYq
3Pwq/qYJ/c1clC3nSZnNMbbTOY97n5gRYYiWXx53g9p7Bb720umPZwDuRSJLmsQi
+q44SOnxb57tmVTO2wHUEA5DIE1ZgTxiTzublCk81ZcvVKAS3ty4Q75nzGfosKdQ
e+QkOpNqGLAl3aMhF9NZalXc53Y2OdhzzaYfOwUxFBi8RXz66aGJJkaePONvCftQ
Bm7P8lw0FCSpS59FiYQfwmP2g9PtrgkVsMSPo1HDgOGwv93KzGjQX29D5vB3wLVZ
kdaH+JjUiRJ7GPBeuXs7SwTVC98WBqlyeaXL4WIpEz5pQvNqpqPGdWuQJ66YEXs5
kj5a7d8jf8JoXHPPoCSTljAoqTcY9AFCjVmp+J5zcprV8wbrXuolbyJa2XjPk6pY
V16AoZ5zF1v+mp1c/QjJVSIbUyzxsypKt7SaUgeFPig/2fUTuG2fvqns1x0LnxId
/NGq6trY/Uf22fgP+wzHV1Ji7V7zq3vNzoRcfR3++4ygnqvDHkmbSDxWR4ZsVu9/
Pd0xEPgb3ltv7FXhErpLF47f1iEieVMTi38gUlGXM8oieZARFLD0MbnvnBg84BWI
fXzAoOXsqjV/GpM5YnhUNwTkVgv4w1huPE4xy8O7WOgbQYuegXfUD2RLEUHDPutP
Lq37kU+FFabDp6QP4nNw0T7mHbZRyfk1o0fYBdoUlhU5yop47gkVH7L6etCAMjDS
6TqHOf8NF8Qyf542JzhdySyFaHaNNex+KXDaOEATKaK4sW8UgLSpjPAD1XgIJoL2
uaiJx5RDH0Nq5WChMfJBqtKwx3NaKeaS/6ULe+4l0bZHYP5wfuHjJjgKPHtZP+Vk
pjSnj7tDXGfHN65mIZieAYDTe9aDp8qpZ7r9Su76PpREBZcIBnzDFFHjCuqbubSD
bsGyk5SYdNUhAn10jqs8ae/W1jWICPe7Uzcjyr9OZJ+GcjCMnjgMkBL/qax+1TTO
FPQdPX2ck/5xALEXymLLm63cdFoF0TmOjTeXWGJ9XMP3tttvKlEAh4S3Dg5vOsy2
AhUT4eL3k7+aZ7VrrfbFjvmS3uQk/3EHrcNMca5L9v9E7sVtU3yAvgllrvUuot2M
EYPIxWiE7/kx7XSt/zQPtjRS3GVXZEpQqVpMvXMqt4nuTEJAajEAkeVHDcjm+KzO
pW1bC2PJRMJ6lWlFHQh/5IhvPmGe6bBIY9+c7n63x6trs076RbnwMV8y3gDI0EX7
UCBCiT9/SbLigQqy70BwVCD3TxxiXuPAwZUA36ILWUny3x+xp9cY1nCyXNl+Wgdu
84zEdFZFBaqGE9m9JphafLClei0Y3GCTMOrAK00NVk3RFqm3ILVQT6+7oHIcLzau
btPcjKutZu6azxvSRmyFWPf1sm7LKeW0WL29EYdzezUURu3u+xHprsuK1IV3QEfH
7Ib2y4Co+Dzwjog3k/UsjHJ35b2N3FG9y4ccna2H0I+7pKzJqs6nY9BmxTbXicAa
l2sUakTTaO1OBa1pU1InsgBKnx7dtzoEK0q56NZ7CWCe6pa69612SYsoceJYagNN
uquVL9uPBQ5bsd9tZ+BR59IGpiZn3pZ/V+BNwkPefUKXZkoRzaxqCRkYXVBohpo9
P0ffJdn6hp5EUR+uQbXzXig6r6xIL8YazBzFwSrPbpZRy6Era1jFdu6J8YhYXR2j
XT4LSHEyQuU/6IdE41qi+y/4Gbx1HC6oscIEU8NmQesTd9XhizAUDtXm6mpNAzZR
5LsAm0Z8VLDOLAv41BV59F7IUAYbKs5ODGp1rco2FZhwzSDszspq+EaXAJmO3vns
UD+Rv6WamDEJwrVwuCUd3G5tIVPJZJ7huLOV0sgQk01odmLsYEugqNQrp4Fp+XDN
g1mQFUTnnYQCk2IFJj/h5Zz6Zewjes6I3tyiyDGzb/wEaK2wNUH9rmfUF1kew9eY
Zmz5l7e/P5npduIobMznOr79cHxSct/Z4sSgLU0p2sYZAwXF51OKr7OX2azzLGg6
/4G8VO+kju+Zl/4mDPO+PLRqwTCjXS6NqAa7k4Vx9vf7SdKPYK9kWDNbSeVUlaN6
lR6Zq8C9BNLopuNGefxhh88UfvkoQH+0VdUwXIHAvQmDK+fm19f/UjY/VSAGAzNl
xSeG16wlv7fVY1k00IsD6hsIhzMNa1amdJg+OOYnzkV1vDB+EwgSNWSKGI6uOH2o
XhxTRbWM86DZ/00zpveqXs9pChfdGGFoaYN0wp4eIXpabH4TyLcliMqvqd+h7S6Q
cVdD3XIjmlTHcpsBaNS+F6Og+lYqKNlzla1zWYUh+6QzI56Br9Sc6uD5YrMatkiO
Vu5TqDZ1P6xxwO64IgJC5NVmcMXXzamuRuhHGFZUF0/S5lIy0J6kJftGDkw334NX
tl93AVBTeVttqMl0cYdj8wWLdx6zRHb3tj4I0PzDbwLeg8jDkL2DdiZivLMy9GZV
yV70G6Qfpwb2gtphXbfPXNd8nfk9Za2XACkheI2o4+Z6kvNuhu0J+aHAQ+0XJgx9
9TqEcmG2JUcJCB0k9D9ZIX6F/Wh0TwyiN+T04czWKP6m98dwzY47BxyMVoKsL2mH
brBK/JivCC9zXSAz1B2YwiDDaSRucPjt+EJAUH/skEfrQ6SBwXUQDHto02pIWgQb
fRaiPqxrftus9WFmnraaTeHtK6dyHmkChqJuc3wJ9uGQkZJn445Uaf4XX1Mvz/i1
T4wpxQlKCTa5GnGCCrPMY5ljfFuAZRKfam31mEjjU4W1kQfr0zC6qKujzZq9zOlc
gUNLn6mgYaZFKoJQx9NWa/jQlwoUOy/lRZaEur6V5tc+4sLHbWbuE5gdie/nY4WK
EgIK1ezON6Fwc91iNAGpz4TFvfrawO1xPH00KJCjeh5tyRFDnNShKbAw66n+qnyB
6g4/4qcrSfMyjFH0vXES8VgG8kMZ+QC1h1y1YSnYSq+ho1H3TLY5KVJuujPOUjN5
SmwW5TDx6qukKoao8cSUWn4+dhyzkctlOrCbwQu+plmWCKZAcOBqweQmeFeqJdIe
AubHjkZnXCGEB+mV5Zcq2Hb6+ftFAh+ah84bzld09NrLQf41zAw9vcGJhbH+xxpa
Iw5+5sG+dvx0U58sFGoVFO4M105lGAeQJ0uZpRFMGYEMMtTj1Dg2HP0941SVsHoG
Mvldgzha7jRgq+5Pe56se5z50irIbbUH0jH4h93QvzMWQLL2Xxq9Qi+8v1Ussvvy
9uvQzvnW1WnOmKA+UacVtgE5xT1xnPqdfvECXjxCThlnX2FzTzJDYeztdieqh9Pb
EvzRxcBnVs2foEtXWEKhOe8+a2raUaz9sykX3j2sxsHNMtZ9Vn/Ram7fsN4JcSfe
orwYvYPXbW5yqrUz7D8vnYB6myL1vMxAQZ8tjKsDMEq3Dk5n6DPgEKmeX3xwYDV7
mmOBOBZSP2vAXytYhUmIGCuNG9wlwC862la8u3mbgWokX/FHW8tZgnl5VZhSTXL1
xVlJHaY1R8KiShlbmlupMRn1jwlW07ghqyUwdZoFsYUYigXpxrrwYyUINdEWymx7
N2fWNG+sC4POE9tnV6FP2/wu+hvT60BPQA3k3gTWwWl3ZartWObgWdw3W8hYNM/R
DitY/AizkTWCE2pIRH9ONb88HdTJcB5ghx1wGZy745maumpBgxaPPqDWo1G8cLNc
uGP3lNM5e3AHFXOOHjcElCJgee2tF4J7ARcp3QIHkp6lpxF4BE/htERag7Fq0Dwo
QmA6MgxLU8pTTqpRHkZkCoc4dBbKnko9QD0dKOKJnLin7dElt29Kflp1keQivfP5
7gqTOWaLMF8qlEXU+jhckZTisyTqeM94rDOq5VqQIQYnZuuraLH72MdrtywrJs5L
BYIIiE52o36oZxuv01FMLs112srMPRuR4o3+oXWz/BVU/sC+40emFuoRrbUjxZjE
ULtRetveJqry19XzkjBd6+6qBYLv07Melzb4qtefgWRnlWRnCInaHp/1JG5yjc+8
8LNFlEoYNmAMocjHKJGaCLEB4me7o6tchH5N+aF8aeW/AbUOhwjzl3MRcN+GvLxm
gZ5CLiWG7y3R///OJIXTRI3PiQT2c5YCo+4++aAzxqmVwU2QUP4S6xnItKb9lbKQ
DxM/lIqCP0teiVzukHd2sLCDHUx+YI6UPy8xl+RgK5HJ56xZ/6Sa8wcK1X5HXFFa
AQWRhNyurb8iughvYC2zw1l4V6TkHGbA8qVIJSC3M3Y1A251HD2Lu2X2ZFVJFeLt
Zoy+0cChzxrKtV4As5fnirR0ixqjM5jxzIPJNB3FN1bxp1Xw2RimnD/cbdH2F5X3
kSuJE1F/bAyV5JMMHQ2hcJNwE64v7PW8iPjR6gj6V6NMNdxTvskCihL2a1LhGqrA
MvkEV/nteSELtidsMWJyZIenWUcWQtyR5MJxz+451E1GXfmTqHUs8c4grsKCGstr
rL8VQyQgizfvfYMUxv1ildEGfDFq2kdTvg6hLDrRJA3GLRJ5Jqd/4hJXGFzcxJSD
jjDhhiOt07VACxw+4m2ijeY47ESnKoc3FCa3Sb0jZa0qoO4a0dGzYjaLVebnBF5v
DeD2GhfTgiRMqj8Pf3mbJqyg2/LAmnybsT01ChaicHg1NghMwA4uh8LojWElJ+4t
q4ZXWcIST4OGY8WM2YT58JJcl9k4MGU6t76JrEvrYUdAkSBMig4d7C1LxAoLkHcA
U8c2zQZuyFEA7qOJUKkRPTSTD6Xr0v+hCWgIXKRQsjKG9XybWK6dPfOdPDhy8KsF
TvSctcWmTa6culfDssGAaSppcgVX2/PB5vajrfS6L5NryliqPCldqAPMVwGrAj6L
2janlniRMhNysItambadYwlOKc+6iDFfnQSplLtDSnFale3WsyQAAnXm+y7m+yhH
5kbgRwJl1O+8KIhWTOOF66TTXnERQOK323KNvO6YS1lfpLVtPx7bXMaabQygy1Xi
7IFFOgox8Qdh7GS2x8Ogmdq6olmklOqykr2/zr6km5yrkp2tto92O3EZLe4wUv6x
TmAFQrLAt5GVZb876Uas+ZTU9aVVl5ykK9evBwivUZnCxajHVuAretL6tpJ0FATk
V5UwebrUG6AIJOnoI2MpA1D8XSkfmcXkgUmNKFHCOQAZPzcTfrYzUbWV7ZFcvPxC
55rJBULMM4NNm8v4ZkXlZ1wWDpHmIFMfX+OxscVpnG4mVfmugMmWZBEPMTNX5VJ1
psewBoRPerd3hRXH2R8qFrrOzCYCzO+PUF/RuHDG29OXH+b9emVlW6ccac5LhDow
B9FUmv7ik8D0gPWidDLIsRzlxj2zt8Inxs34Y+iMUbOHPcaaH3inrrR5bY7NfTRc
Bwa6ctmIi7aNhv7hkVhpYr6wenE53SElYAbwp8zaqp6u2eIg8+j1ycdUqogeryGY
hw5WQsj/pZIa6oxIkSkYigMHwEgAqJagFSRp7NdjQV3WjBN1KwfHOBIgotOfoSWr
xCuwWfI9HKg1qScAZc0L9ptMdLfzmkgWSeEUeHMq0FuGlqZbRUnW5G/dJqXnOULE
ZdinVZvXL2jZV47w0Ppi8RklvA6NJyItW2CoPApiXcUWxqULjrLluCVxUMfjdOWQ
0HZoBvtqqOiA/nG6CX891xMDGOGkKVX3act18LmxH3UgoW1s+HaAlFjAd9M+vJhb
BPU3RWnCLZgMJxS/5pc7KQC5EqaGrzSlOoRDFY7ykgKnfXP7diQ4F/rQ1brHkGOn
EAw0ZnCpkXYTRbZl9AUWyZVdNeCFvMpzM6OsHUJnhLcMyKycL6w4lNJewr0lRQ8z
5Ehe0lmU0ADwdKcN3EQZ7UoJz1MNLY4Zeghba34u80q++XSIAnDDhyISSfFikf22
U37H2U7HERxHtD3zljI0EGHmPxh3xHGCPrbUmRTlPVUOm3TShUf8mhGa4wsJJIuh
yLc9ofXaHJJa4j4k5WxRY6fHM7B/Bv+8YjVZY3cs/zFT5NDj6EN/BgyW6SWdSbGV
QFlk+ltGYHvHfqf9VKmdv4lnaklzsRSCzGlXc9+g639XwJzvd5FXOrkhq6B/4qWs
W7M7YPaGorE7ICf2GKAxTyYhN9BTtETmwL4STZIWdwPTgKVxymLHexyWQvPygSRv
tbaup67fJ5ZOqNeSqicJdBNKZHyxvi4bGQJSUG7eeLVPQYh9TM2lZZHa5l3uIYcJ
TeAOr8M2UllerZKYDea3dkveJKJupmA//fA7XcnMdNs0331X4eDLVdgaNzLC9Wf2
S9KvJEaDDvf+VttfSm+xQy9MoPc7DIHjmtUi/AjPdMThs9qQB/qg7TyQBZWogHW5
Rl4qfayXK0GPPz7xGheYsByadfD+ObyH9AcS13upbcsFmw9LAwHz0ihNR0KxRMZq
9e4T33uJWroqFYsxFiEpudIG2I5ApYW2TfbD+cdb69xy71Q5cAzomzGBqLzoYGo7
Pl8iwRaVJIbJQYKXpbD7BKkUEww4WtZjYdjLlRA7HRMXV9ReOHcNrvpIOzyxXk7L
Y6L/NTvvKR9bpwEakYg/BOu8hIvYX6jJ7YP3T7EMZYxWahiRmBHMUXxArmFdDlQB
JdwZnORlqO5r5BN3rjiPVZhAH5SaAWWNjdgarORcRRR62ffTyDh2FF0bHdWf+Au5
jR9tTHM3/qS8VrHLCAcoTKhaCBCfgwtPlPKWqJke8cKk1gYXldpL8F39q6WE8RLB
SNcy8FtvnBjZ/2+0oMztC/XSjtbWMnYYvY6Fl3iFGjkE1nQ3aWzF2jZkdTN4LB58
eIfgEsn1DsS4Pql31/IZ/aSGNQOyZrIyR70pOYf63RUK+olK/1TSWhycrQDpkjtg
w5oU7YOBBWJqI9Cn/OmXAtiitnPyxxJRg4gUoy4qSDmifMb5AfbnLJuwToxmBeT2
UIU+aItn/luVp3a6lMjo7TklmB8EDXSR2H9BxLgqMRWBgye12rAy8Ckh59CyyIGq
l7V1p7Vlv00xr7bkduGX41gcIaFUDQmlQrqRoUyxsMqTXZ7gatcbGV31QPIsAICI
gDSB/6/0xYe1lD2y/XWGrOoKv4OeAi2ejq+Q9uNiJc5a60QirNgL2+vVyUxvD8Bh
WR7aG/b3ODqfEgVAxrOcuR20SkvQ5fhhg+UFacuUk6c2WqB03aBc16RSpnNrBOT9
MLg4xxjaM5rJ0Pt9mNRoibnUadUZTF4n7c85dAQPr1foqd7PCeEEa2K8qAIY25tL
RLTI772qxpucm4Z2Vxqwq8avhufLRIobqgcBqw86mRfvv5bRtH5qkSI3GPSZeyVh
PSEI+XWMibtpmDAQ6haRBY6j4PC+vyrxyePbkyguleKkO4I4OcaelQNiih3LqPdF
s7TDfKUReIY+djgBI0OlZNf7nzHck5eigcnTx/k8XXHB1oCCucwTpKksD2g6DVrD
rez8bB8QWwduT6zStJNr7TNWHu5Khv6DEaRnBqGQQoKjilqDpLd9ddDnfnlFymeC
pVfdxJ+2FMepmviqO4NGoT5vLI+3hVjtFHYxkgPgkBxeYHAKUQTHFtheIqYXVUQ3
0FihS9SD+1RyKK3ngMtNVq257f7r/Ngw14L4luDqvGrEw/71x+kE4I/EsETwTnX+
AKBQb0ddORyb+70Q6cYdI+S/UJU/IH0PFPmLvmC+D220t57neZH/0qKsQNEks5dK
vwjqoWeT0KdS+E0xtGKs3JbTkCkA9qVzEjadXD+AcjzHWmCFmJkdFXQotll2jJEY
vXnf1DpdAivqhJ1MsfHKC4gZx6jtteGwNkJyxG/0F3Wx7Ze/x71lObINYe8iovKZ
VJLuGP2iUTrPO9SEh42OTgZXFpXjuy0JtPJ+8qwia81/Cwo3Za7r6uA6j9keBgbp
MaWzW94EyQeUtZw/nitKtAt8T/Wlxsr4JamyDaZIhDic7dTc+wtdxx4Vso53yryT
pE+YaVBotfbGC2ZsPPm4Q6AF6tBM+3VBSXFNK17BOGE2zTQ5E1b8D8JJJJIxTPj6
JTVJVLHqliknjSdGR5uW1HjVtnM0/ROQcV/9FCZJQeazAcW5VwcDRR+/5aD7eurL
jZuqzG/6S7Z1c7RI5Klj75UCJH6FK6sT9g2qr7RFJvI22hAB0RrdQAc0A26S4PuR
UdHNGYo4cIrfW+iijYvLq9d/vvDVFDtSTxx63MLTNOWVEWzHp0eZGnMZSYos83vw
QrAOLMKOfhJzKFCye1W1ZaeGnLArl8vGFzG6/ksYXDYB5JaPrQnq0UOu908IHRrZ
RWHuM5ehc3XcaYw9KJ7XECtgInw9K+J/q/B7SktuBnRLKxrhGrD0uXjVz9MnETuO
DFprPA1QkBdjdRN3xjXXdjneylIvEj/Z2hUxTsK7+637nes8nR4eQ086siQ81zkG
dxGgzzvC72vAQiYqZiwrn3EY6mxWqL8m/3MFky4meDvx7K26QkT/TXzR3VkYBZ/3
znymy9mLCDd78JAyIXcrB7NAjHhPcuvAm8wKnbvmO0PYKcjGjzs+fsNmqNmy51h9
/cGNHmJfoj/lyXsZvdDJX/I5UyT1yy7uBolnZRvlVQ2eramCxGCkukCO+15EMV5s
IDHqie+rpi1zy8cYJ3UIYiA3QP+qVxcAn0oU5xNEpNvuJLdo6se2cpINwtrSx4Dh
ovErluoe7qvhDTQ9M8XF8xfwQ4xYaiPh+sbUQ5NmaR6r56S2l/1Dm9Eoce0iHqgQ
o2IjVceHSmaIISG2NPG8PzmHqwDYL6Cu3qjg10ydp5mk73FAYzAsXMrZDnXbmR8y
DX7Xdp5Y3l0wSXW29pQvmiR6HzMIuh1bHmWVhOVu48hVf++SOBZCNxNXH3bZeqpZ
KnqHeDn71OKP7J0AaRvtQqi6bipM4welHFYvMwRxvdbtVnLA8tqB0ZHydPACz9ks
PXJdYxWhZ8MEl6cXBnApsoVY8quDSmt53T9Pt1wrnZFJ8TqKsltqCPLN/jKJGKSe
mDz6nfDhbw3mn8zbnW7PpQ2/2WnbfyNE1MPhYYAEerV1Kp4FPY3DYy/2ZzYHD/rm
OJTgXzWNl3NHWhEGQ9hk6YPWqpuX6h4K97ud3TTFgmfazSF0CgcgXVAc8/dE7f4k
SvL3oWEUmDPM7z0fPMIi+l8yqBLlM1ZECuL1pi8AtCrcC4TRz0Jm+iL8uQHJq1Kf
Yd6nhxm1lyBptrC6yv99AbvD1ZTYq9Zwj4PVAB3BKvZpAjp24Ej4/D3gmkm8tJk7
KMv/FeyIrt+8S5Z8in3ENXorFP/HE21LhwozPvm08TRBjtRssNqHxhgxAFLGcS5C
m0YtTHJcxPLQ0MO21qzsh9pSPP7eKhJt0gz5/qyNNj57c8AV5iUr+287LQC9huIn
d7m1IX4QYXEMX3slzzXUG79PDfRc5/bXDESYOdmsMfhwjXbDUEAUmuZ2FxYfL3iA
1A2NJiNX91CFCzg2yUK4SaEEkhPvPSplY0ratXyKMnW+kAQ5s5zPsRXxgcGCpkc6
e+NEgV5xDBCDCQrwul9W+9VgaG3X2gzJQyF+SR08x16fAGKVelAdzXnS/Avd3sNH
cfHkZrj3zE28Mekhd9OU5I9NasKB+Cfd73eFxLxZ0WSrVXRaxvPXSs8bBiySnErX
LaESH12CJ7ZUCdeZ/fEInZJfLktxRKMQ/lLTgPFvrEIHM+mmf3AOKto9/t2Ycv2V
IJnBy6kegZL6aVVxwhQliQjmBlLR0AJCvdTVXLb74BhttQkX356NS9f98kcrSBu7
7/xYTstNGU49wm8eqYiQc7kpphi0dUS0QJt+XgPUwMjJbwpH8ompihYOVFk5/XI5
oahhM5cPFEUMpYqpDgX4FQTuu9yHIT61C/G+ACaM/Un7kgJE7cDsDpg3Pbl7PP9q
0FWz5L5HG2o8arBITkgyi04aTzhe1UjkLX9AniOFbCDb0Ux5G23fOvCoyZR8vLm/
SnI6nBKedm2tknQFrnbxwUI0zwspYNr9aCG2yiaK2+quYu3jD9Cc5yYaeS7+51nC
Bw9b4fg2iZOdiYgXvn1iccSuomQ8kEB6sE83uc24aHD5IZh7X+K9hirh1euGmvSo
LLndOM0p1IDTNBFN80mYQ1otbrlVcXpmk5Gii+PMFESqcv4lbDs2nHSVIUool/4A
ynIXSkw+nO8B4lUZo1yWSNwdnLURwyeA4O822w8d0Nb9MXbwUwglhs9U/XM4d+8z
Upg3L/obqNLDYYMPVI/agQCFYsEFKT0g+SZZ8aOg6gLaPxFgkd+L/TgZye+CtaHN
ECqFx0KiJXLb3xYQd8G5lu92yvjGXg29zlhxQ5c7ZZkCK/XouQK/zCfOj2Z7jSHv
btUP0KeoTm2hSTI1b3CGRuO5Vy1fWzmcO8HtTIlvE+bgJrwDpcKWmurLl5zgcoF3
I9VsywGR+vxVEi+oXt1lbnY0eJH405WrJaKrBrovroDoeY39ShHSnB3Il+QZ+Sgs
51DgSMg1cPNZzhp4QqW41ZLMYpRRaZ8hu/s1EhY6cBjco5dYoZ8p7v+JEar0qAHM
V9PZVO8iDX86OFjQ6Bt2Ap9RlDgrTDHRGHyBGrln8eog3EiJMypiglojiYyDAbQG
hvyM9NJsY2FPG1pWd7U1ppBIUsvRCBXwbdmttcHMOgexOQyUCDMd5drV5H04QiSG
dxvwMhpbw19jis/cpG+4t5ViUtpuyQlsnFI2byGvaonGrtcFn65NcFYh65e8jIph
ESKLrqM2cAcCm5DzNt+EVT9RHHEW//dGjeb1dZsezdAkeqT7EI13nW+mwrEieno5
WW6Untu4aaqK+F58/Ugc7Zbl7MaX7W9QKCsp6pMhPSAiRb7TdX4CTA0eYErH4FuN
zvbMKfkPO84Fkrv8QC6LY49Q0pxvf+hjvdGE3PFAkfMvI9jISWOZYVpm43D21phf
g41VII37pFVw7e60TuCPdtFuxX4i50NnMnoPm8hgjBfLFjC4aiezJwKFrPzxTB6u
PdX6/ZCsPlpGxJXujndsqIU39Rl7YlV8zfINvsj0Sggjo6xxNfIYpM9/Qkp+oy8l
HkLyt8EZQQaxVV6TlPjVZPvft6+teR9srcPFZigu120uHXB2zo9dIjkvkD5+SWO6
hcKTHf1WRynDy5z1HJ2tpZTp6POEGQXLMIEMrLSArUwDcR0aaRhyqxrrNJ5pgi6A
6aVIJ2eCEKLkNYezkH5Br2qf5MdnRA04jAwzmEE/MzOg0sHY3o1EnPGWwYJ+C5Nv
5apWEiNBQRfiPv4jpblLXJUBXxGO+NXCe0fq5jBRntxeqCaziglUgK5zWC9LMojq
bHeRmRofoTBBkVgJBWNkmKHKkmd1yv2OgbjuTUTjDt29welFQf4KkNPK+5HOFKpg
fvKxyTT+1kxRYK08K88Eol9QoXZhlPQtF790r87gozm/Fld1p9hs0foAm3gpQLg1
N+pksMGJC7RaFULU3fh0ejVBQaIoDADPYIfVLP4x8JZyQZ/gnrB4Oiaq/b9zuMX7
x0FLE04DctZDu3i3SxXeYiewJbiCNRFcBojKnVoyntfTazBtDfgOAaE3HDBJIPpY
3EsuE2mTKXJqYMPJSvU5+gnVejY3lmZnZ4jxbzBSJeyDu84gKqWB2yJqT/KiJL25
Rxgo84gk1+0G63qCUmrDRBmEH9WxqaZttaduPgOS7Bac1FaBf5KYjLgzkI2muNZZ
qEJrBMO5eSqTf2m2cEghx5zjA4bU+SpdKEZJSImmHvMRKxWE1tTAiekBaXJjg0Aq
LdhR5x8BfrAgW8Wc3i14t7Lt3nUzbxTtNSTmcGLA3uYbDwKQdm0IjUQEOfE112G9
hf6APssZCQYqj59n8S7xhD37flBi5sJpyM9OJkOVNVWAAg6ugreRR5zheuZTd5/f
90W6V4SdTwYoHCquN6EsBfl4/XznK80B9O/dNzDOQjgDKm+kpgxZy51IjX7MzRnf
rFOMH0y9713W/btS1PoMBIVHmbzgz8Xo/as7qmGz0I+3g0nE1lG+h8k5bc33l8h4
rg/egNktAzv8E8XKo2XWI92sPuph9BopWf/nfaqi0v+2tSf7Q45ocJAgpzXpYfhC
mZcwTomNFzuxrld6MbzTrB1VIQzJjMEcRyOKj8Rs6i/clk9yVrw5jHM3GJM8XKtI
F+4/grTOFQ5UuP03rApxFGS8fvbuMQexTmXtMyTJXziyvV59q741nlzj91WF9g+b
diikpYiwxJ5bhXHID2s5wouviFj7fEqGVL6TrVuqPMhxouxeqYGjA515S2WHrFci
JJX+woNAKJqElkryusjb+vDiWKpuffOrqT8HW/RcGqtSjf33DcqGN+fRPyjHd/if
U4DkEE8PuaC7Nxj3sRZ3iVdRb/LLPBYqJ4n9nyb7Vp2y+p/ajQMXe35nBvbUXod8
Q8XR3ICJ+Mxew+LLfhUd32VwWU0v6G2dfvoAh319ctdI6MLxX0I1otNgGdVzQjqv
VoIpoeR+fY/rJFc7JlJxGGDrKF83W15Te7AHwVz3EJTrRxbASkAuXpJ0/WxfaxBp
5jbkcD8v0mWnaAEX9B317Frj+W9ywZu6izjfV0QOOXpIEE0Wl/iRzgEt/P/4jcy5
/IcmylcIvi+dOHBJVkclxlbW48d1F01Q/K3ummhNHxh5rvef2QvUzuHlghbZ+Z4S
ixmKiErsoiRkeCYSwm8jsXzHHoxA+sAWOESto3NSd6PPHVsTU6/9wXgU2nLfvakt
jFAOlBR1Dd00vMTDDCxthZwHhkXMwppSmn4+MbkTNFllS2pF5sasLPDsd/koLH1O
r/Tm0wm0UG9iLgzHqtfc7kmIaBFgKzrEasmX7oie/1aUlvI5/DIheVN1lmEdLJE0
rl8eQ3+dG/NI6zNQ1O74vZpcZkrOskA5bus1lDOkZtfbSysKMJZblnitF4aDUr+9
`protect END_PROTECTED
