`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
da1J8HHVQX5bngXeXmJ6gQIOwqE9rEWrdllPIp8KXbDwfHq94uImPSnVjLXUVKAT
xfh5gYKPto79H14ZnXIkTMiz8LmL3/ty9fMOj9hIpJOjjk9AaVXsfhdiKocA/g+1
QlghFZOFM1EtgMJM6M9ScqDHihE6044+mDL/uFXH9Wk0zYgi+CMCM0yMk6wlTHuI
dCgxP0b11G7N4NPfa4IsppP+6iLnR1wG+rwe84Jn2tOh/xTsO39ynfHgfg9plHkQ
P0flJR8a5piHsk0hfyZaTbmGEct48OzpD7I/NMVaXwfgNL7GbJsD5TPe79tVuIof
DjknfdUaBq+jXvu+217AqQcD8iz5YBjzsO+RR5OuroCMpAfe5LUfwXUJnQqY3ifq
9KS9wVu7J43JSKvgw70VuyFz3DF2dS9migRf3qrhBAhAqQLjBITw1fUtnUHgr2RJ
kpz2mco8oP657Ahs1u6qGiQLOFoVXLzbFhxWag64XadH2yt9EUyLdMee7beH5U1B
2gB4OyT/AUg2Iu5Oph7wbrBLmuVwVqT+NA08r+J2uOlbxFW13VPNeZTuD2b2CsGM
lhmEitRNKGxHWkf9gLc0CSHoSzwdo+LtQSwfLMue6L/bS2XLVgeFwagcDnwqzPNv
t1LMhTvLCtR0bUO6Iszl/QTS2ZFT81OCteGEeh90eb3Kc63STDJox1Zcl17jxs0H
q81fxPXpM7zARKq9Z3dbQ22m8rq6D24VLbewYbZwBUQ=
`protect END_PROTECTED
