`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RIT68ePSpvOv7pERzsqBmOzMhWVcZuobcCly4pasgZBGBi+qegxTsEgOgP6U71aN
wdK6rdLPGut9kOiAH3bESdZWN59uyZp+U1bOvrxOg/fOzOD8g+xrDu161WdjQ14C
wPjBvfRXHsZscQk45e5BLTmUfT1e4DaR78C8wGMNdtXqJFux20rXUDiyoGNtTQK0
g79eZ+I0ZvH57FFgludhVZ+bzGIVH1Swt8q9T0t0LKlSS4ZwtlBOjFb9nLQMQfjO
JA1a3GVWnldQpiWZsVtdzIhQCioz01zs8xu3elrBX1+GwrvuMca622GVQNcdm/JI
0B8RK0K6aKAoQsRtA35s9TGU9Czkk/oPTsuA2p1RayyNoxBnZ+APImHysE2xvM14
7MictJ+09pCpJ/rbQazPwuPniItWtGzGRyKkpqt5P+avQqzF+fi6Oo8bYd80iawQ
4AzEQAs8/M/4G/n4gQ8pt46QtiGNceUwBAUIcRABTGGgrOSd0AsvzJzvIvVWGSCj
6zE5SdTjLkogy/rD4NTvYXRnWpChWPlyYTK21jpOGtHSTLhe9J4C1BeqLqOHBjLZ
YzSdjUNnqKcmaulZUeMnsZaszeaYSmCqLumcyUD+dRHs51vak7g37YpO4PAz+VmN
XLda0/NG0pOvbyMXKa228xV1d/YZrKQzp568bxkYR+MGxDTwHOUwZi6BA6NPFMWr
aMjerfCIdXW40W+s0UeQ376GFYf3Vf9qQrIDZ5IJ5UgQmsS80KMQiBV/wfDvxXZ1
sBHFpfEdHsgZNWaDvW3roSY26B5MH9em68dBVIpqX73+Ek/964y9EfGCTK+i+tPY
F5+2osvKbrWy233S7XB5oblqn0bRGxQESRjXlv1VnFK97L1adLY7k8UnA3ZvHKFn
pYaghWI4uuKOw0PoJAax9yoJWb0afTgDmvpFM+emDdUbaJUxMLiVomgSrSY6KExP
2LiZKZsAOPY5+c96KZcBKa6530wM6nGJS2rxr23yhiRDvvtZJDiFo3Io6itAhJP2
utyAxE3DAbLDgsmAUk8SmObx0XHB/9sMgd5207rAoAnWhu9FrsgR5dKA8TLpvb8l
nQlgEvIlnsFXIlxhWkLmXz/zBnZtcp2p8/ia2KBPtuyfnEICc8+zNZfBY9N3W753
gjBdqEN5pTol7n3BQAWct80eMPG5ZyojTMyGrbplEd5NAV5Y3RMuE8f/Ryx4G3+C
M39VC+1JO/tKVZM1mBD3OXumUnXzFG+bClTMDZRMJV41xjhRJABG82eZ8QfVFFsk
TpdaXbFSGhcnFOWdjVGdpzKpjH7qFkdPSxw2D/p9t7z02YwD4/3Q0ejBodCeuNaQ
ogKSVNBa6nfnCpMkVh8Zi+8nIiY1FYmnSqsfrMPGVLh5E6DJfVfHe+LLikvh8T9z
8MWpGc/FCrD+VCWNHW/XYhJ4WpqIX9tQeTH4W+d4gdPMPu2hMgje1Ka9QVZH5GiL
WWBLPtKMfk1BM7/EgK4M0XfdgQEttIhMW90CtSvOwBscHt7FjP2eWzvRTtXebb6d
lkP2rqohnCFfoIKCYDeGkTsRgPkcauQH7N8AApQ7/+ZxGDXBUV2RulhHcAJ00xou
YaI2ioU8UkTkgJ2WRFZ5VmSC7L6jM2u6NwTSRr3Q1FNqRReXgokloo8Z9+oN0LWD
J4G79GL9fwdAO2Z4fqzWIxfSWcF3wUbEol4KW2F6/JB5Ywt6gFlQd8dVymvP9yCt
Re6oM+mBAJbrtLKXdWih2iXWQtQR3LXr35kHAiWFkBhLF2SZR/elOrdPrNdGDP87
tA0UI3VZYb/m/wFxtKuSXPTBUJcdfYOfmMywWxm5Jv7VCcBh3zb3UmK0uxXpKG5l
YGnjuKPwiLY2erkUx/Z4zM1wKp7TSJhdgYA/ErS58+AI9x1aL5zQtvbxx5eBNePQ
gKbyVMjzwnDzDLX0xH1Jn2webqW06A488eC7E3VVJ4wfGgyOwgpeABvaxo5ngYHw
ofnduqmXnBU0kMGmyLy5mYrA/TffI1sQie54q5pqJweo2GlxqVqe7v16qFBKYHor
1dHo8r5cfcRgTxCc6LRppu5r9B0rzOS/Q9OHxpQlT1+Db+uszXPFkQVSBSewXIUO
SyEqz63t9sqfUfODuazxo0UWg1WSYjIfFvFv9zLquJIwAD3+1c7Go+fO3lN7VPLE
9olHziTAaReAgK47aFoleQX2Vh7ihWVIuGyxj4KdyfHJhyZxMJ8PrhXd0yz8jISn
31nyGLYjYAH5fgQHJfc0OcStZVyxcQJ8RNsZNgsKehIqAcn2FeC4gMavhD+0WpNN
2klpWkFv35O3Qhw2fkSMiiVddWFQkJBzOKJBjyDAS9sCalkV4kC0c3NDJs2YGgyd
El64XtWelO2ZDMzO75JBEng+6U0Q54ulgF3rZNBpmZHVQMjyP6h4xlVpE6AuET/4
h/zMrIUNbNZhTRTQxV7tfCvHrhrEJE+4LFJ/mAFIdrxBKkRNqPmmli9NaGfUnbvZ
iFUr87e5ZMVPYswK+uUxlt2mhGbUX6+KG1OXuNcioVYeOG4a3gNkIX80jbebBjR7
RzlAgbh3sEVoozZksOPYCgsa0ESnUCV4U3LF+Zi81VQF7XUxhiGtiM90W6JUPqm3
jbjhJleZDD4vLEKrJndPwvIVD4BpAGTU9YmagmEEVp8z1+qYXePMyQlThNebPDmr
ajBNVPEu+nQ2+/UIPDpBZluCvSoDQ6RMTkMdYbcMs7X7IdSFkeMDmnWiSXOFGZoj
/sry/nrarvhbTR6vc7Q4AagGpVU6t50+zJSZrLOQQa/sJmx0tgYxavQ+Yea7LJeJ
Z3SQC5hxdzv2CUvyXeeQYjoUXXOZa4YW5Ddwr6aeqSRVvQlUF3EiOpWLLPCst9Pf
sdHKlcMSnI8FfbTfJizYbZWM3QlKUZWs8Lwwqb6AmCfITwBC1bQc6at2TMFID/p8
CHrJi3v4+6IGzu3oQVN79enZuQStp7yk80SEMd3NFe7GDoT2h/l5UaHOwrhfBo/+
YEx8Q1WnUVpnKzs89nbwYIoOWd7okl6w+Kl+0nY0gN6Bz7Y/HD1c6Yio83a0M7uA
+1D7frHBwJgPurhENC37cQxlaBA1F8inwOs8EbhIWHEU4pBFBAeEQE8KmKHPUV17
GkHbLvBSZiuKmEdyu39ofmAq9ISQFNqfjaCCJ5nDwnvkqGh4Uq4AvOdjWQ5g93sN
2n8O6Mdc3JyeKGlA3sg+5CLA6EbbX43ZqvVVWv8+gJYrHF1CMAySG1n068nu4jMv
jxU6IYYzUR33C5JTv1It1zFsXRLD8WNeKqTo6N5YT+S65kQn8FD2GMC63sguHTI4
wwqKVd8DEc+SZX94Fqa4MTbMWX11/O5NuH9owAwzZTsYvtJ2uFrzyN6c4khckDx9
3WoQMdsBB97tU/2wudQ1mtNjko4DJ0QNRDvKjBx4c/GUGDHywN5WLLh2jOk8Rtax
BkAfCOfSyf/ephks7LiTaOF3bB7a3DPu6abVUePc/8IyruWN52d/QGUN5448i/qu
GyfPX/jKzl5RcHbobrZHyYptw3AU6om/bKQNvrdk7UgyCyftxxe4QZjFWMP0Ity0
F7vFJl49Dn4ZKGTObAHU6VbLt/zpc8DhMlrXu/eUA61qgfWKCTNpMlMclHRbdj/U
6ddVO64dKjQoPNxNmW+tw5v/7BejFaTrzHMymGhHL5gb/IxoveA53n/pKVzBH3zx
kJXY9+CBCoISSg9a5fF0BlGN9CtLNhkal9e9sdW2FtQsUgscBi5Xvna6uyZbnXxu
Utb0gcUhZAdxGD3PP3zXmb498yNbndiHLCM3ZnmBrMcnX2yBKKcBvzh6B+BhHQYr
EfPt/ODdoINhaUhkYK6zDOpn4AsOrP0oepBl3QlgOu1H6Ou/VCR5ZetllSvzspWF
LlAnLrLWyBGKUeku9gB0Bx3zxrQ+b8jcV0et47xHrlz/M0zVJMK9RpKb/KyRimxJ
p+hDYcVCqItK6y88YqqGvH8W0C8E/5Acw6ptgLgtUeDdC14omI77GOPBsdzhg9pB
Ms5euNNWFTl7tSJ//91PPISc/UpnYhUgPbv2SLkxEMoIgnXBBTFp26s9+fgIZqV1
FdDDJA/VNZQ5xlnW98UKCseCv9vZJ+evggIXP+AIh+KxDzPwBBaOvsGsPuKKMySc
NC+dqC6kiHVm9Oh1kZKf4gNl7X2VwrEjjTpqlN4W1Y12Az3DmvMjiJLDl7qnedR1
YFpdvQUlpm/S4yvQYGTOAXsJb2UMiOYc6ZoD0MVSYXuEYQWC5kl0t6PYFV6ELw2w
IqdwCdEX2MQYwyMeUhSXdW7a5pW0PGlVA19c+CtKagsQEiEcY1SH0AfD4SjBdl1w
ky9kJwQmpEGAejzeDu//i9M3dCvFXn69+whw+KMXn2vQDSvpMbxjUZBGHtxFM+MI
Wy7Mv5gGRPWmY5ycFIW6C2bo3GJvQbHioCWDYYOW3xB4DjR4rVN1hckFxTUXgKpv
NMJo6H+hCqZMZZgLmcaHi67mDpzWO4iubxjjU3Y3aOm5l0vuikbE1lRqHRCugzV5
2wOIDagnNNOmaIZ+crSEOWRW2uA2UuCOyzIpQij97PsXV2/pYSa2xqYLbaxPx4kZ
25U0KOdmh3TciZfWKjSBMn6jKWOXRjJrlWUiSANrdBTKc7lhXlRq+MLO/Tw1RusQ
NZnx46wJDzuwS2LV5/VLjvO3/4TQeBawJuXhQnBWdZktiiBkW1TktOuW54itapAH
iIS+hiF5kzDa1EeAIO7MSKrpS3z/gjxYv2WCT07Qo4YyJUzD5TToo7bhY9nHXE7H
x+ltar18WQe4WMpX6v0b0xT38arIS/eakIw8NgH/dFuBJCI+BnSyeHF6b1dp1bYG
J/wgaTsVUVR7zg7Xikg11UEcSXX+CeNE/a02CXOba6SIExHixOafTnqslaC9eNXC
iImAy2x/2sEPWDToqqwc7u3o4lkNBKi0smh2gQGcaFQc5ryH2sUgph4gyTx4uvDc
Xx53PUMNPFmkZG/8+QixNzQh2P/HGwjm/qWlUq0Ps1ArKuJG4rdyYyn4Ef5MAKwy
jazz2Z+jMg0jTk+S4jvQOVPPj47GvOUhCeDCupJzU6PasfSx4tlOErgExkThBHK5
5ERyOASfRPLwG5lFRwjq9Z4wXDmXdOwXdKslwV2y6anONfGRDK97o8GZYuW2w6ZP
OMVwm6I5hNfqMgM6T/ecer4vXYqYLllr3h2Wd7XduYkhKulZlnNLETDUg1AMSQEq
lA266DhIp4eHujv+k/Hpfo18uWolzKOzuWp0m+GYHcpgJv4WRj67nN17ebNjhcRt
frQn2VpzjekfTgak9hyuMEHw6mdgEnWv49jJgwyBmAG2jdvimY/psJLYj0nmvcrH
uRCQuKe8y+ZGtYmgymY/cEj/7cxgOew3BE9MqmL63/R65jzJYFzRzck3COkfz9Dk
gJoBRK14haIXbECfdVXzgbKTLLNZ0OYWuIOrbXUQkaiHTgf5a45DyLBij3H9k6YI
SoUANemQmtfA7kexmzoxQkYNy4eFfKzoqqrrvP6FbSgdDm/ScZX4la0H8JNnOXzN
7MNgOOS3PJF+MGrRkZPJGqC5Y0BqXXNLCray/oFhp4Fe9XnhFlhheV4lm6ukW0Kc
JbOXyqyIQOlBB0/tx+pc13XrV1U9yY+DD0IuSPR0vg0HCKQL6aI72iHa4Qh9oMt7
JRkPjykH2LUPVe9VJzW3NlxULGVAJx3MlQVurbyT0sM2UugJXxw0fBLllgi74I4M
n2PzKB0q8Tzhi1d+GQITyOldJrj464xUV7JKQwvvcisWvfkgzWVmSaV0EA6fRipe
FfzXL3Ut9C6OV2wLlVe3WcZedyD4ryecr+zV7Mypla+ECjzTDJvJszN6QAJdIfqN
Xvqdqr1drBrnUQHJe0OxNgNEZy3dBiII1o4lhf8AGQRA6NHLbby6k78CTwM5NFM8
aNsCRTIY1ZY3ScofXwzcN9YDJVoNwvvRCzGjh1Gi3X7tejKXD6Q0VxFXBMqeAVdK
rHAQWuULWA9JO3tf0T1NbSj4/d7XeagAZnaYeUdqaQ7B73BuIKiWEuHThnz+B8Yk
qXRshym+QU8FSD1JuJIyKoO37wwWRW/uRP1C7LFwFdgiL0ksAXe5jionxWAewJv6
iJLXzwjYZgMxO+omxh15s39pwow9WAQCzZ8Izg6uXNtinPnzJmM3Q74RNJxkl5pM
HzuQBDE8XrgzTnz1HLaVVORj49SZ4nRKD/yatSGTe8eXXuWqBH9yVijym+aAzLJv
DQa/TuLQ1SPS5fliZCHbZ93KYhOxoZ5JYhb20Co0qnw46o8+PQkWJArVq8p456WL
6ncy+n5nhYCGvlxalc4TUfw6Z1j2QQDX8FAPXVuPVvm8EKdpWUB5UtlcYtNXRvEa
zP5Uj3AmhiXwebyeKulGIhr6wrP87VkjFoSkAYbXBUMpxHaCASVoE/vYq44OZEmP
N0JuLd8jKFySJFVu2znZv39dfEbXVd5dlTh28fGEJz3jFZJFN9c2AaYtr/gxuq+r
ZTgct1AOWGRzUGSqKzrr7gTkpFEeDpfQbnf1wZhLevtk8dHaaLMnAbk8v3VGdq6k
45Ewn2SH9+jUNdnsxXfX2EMkq6YYBzFfvmhPAopnNaYhjL7D7+EVDe9RWQpOMwPB
6V9gMQJJqXbEQnODwQdD8RCQPsqAl7AdYnvQVQpjAl4NDwvSQpbbFIJjtKocRdlQ
QOKXBskJ4UfHQghbN1xUGQiOrVNQraQUz47t2SaoMPAN4miRcb0VPsXhGyJ6ALck
C1b+ogm2HtjP8iV20T10BM323OHvws0FlG5xy0dK3y1ci3din4Ro2SW/QofIxCyq
TFeFnJ3aDLfoBiE5uKjS43yvrONjf3xpPNTYpsmchnoq/p0KbDL/6Y+6TIBkCO2t
oxblX1u7okEpbNp2w56Z4CxjirCSkLyiixWRV82P3WziSlvwv5ivePzoV3l+rPBk
6+DFMA51MD3DPPKtDjtNRmV/Ik1Br5iAlUQVmkAvFfQxZSBmS44Jvpe67gf8ARS5
H9SlnGElxUBjWKQ/KQpcR9RgEq1OTF8jqt9mnCrcBWwnm0KvwcZcgja5+JQnAuFn
PiIl6EnBVQxmqNtd/1tjXJtrJBMukBfFlSQJpPDEdYXKWw+O4HS2Od0e0RXgB85O
SpRrLHZxi0tZfkpoldoJ3dI06DUS1SrjYVWE+4XUi6DswUPm/EVGdzzCt+yz+3AG
MEnD8ggDiOyxnqs/oPJKwoRwtOPuft0S8OgV5dR687L7x13RGjfrHqYkJDsqmllR
TkmW4dORFN+0ZjS7DM9YrrvrhSDVoPZadauccd6E0fYnvsHFtXLXID3yx7jOGu0y
kKSlCqDoNaCb/56OUyPg1RguMlPitEmPTK9VpyDPTp5gE9m2mVyRXGJ+V8U7mRFd
qcJ1UDrwOsZKKkEMG5ipX/yIhNDB6/IV22As1E7WN3VrIpYQ2S7JZoV0Y/v8nIwQ
b9xPoJwCBiaK5ugiT07IoKa8++KYlu/q3qfV3yW3gkD+fuxj9dwC9+GWioSZh2kl
JzT+BN3BF+ZcpVNBkspebRcTj0RzGAgt7mDTxcSDu3+dzetkYwDu4C86xd8wlCXs
Ls8kqB+OeLpTmZLnIxygz/hgZb+XoFpP+1YgIvv9EhjvyFyhUP35nGnRNOKD9Qjr
W4vJ0HJFczTbKbzcPJ6s75C9oXWP+2CHDGG3Jcqdp/gkX2RNbMtcI9G/icB6Owv6
a0s2agmWTMbAY81BI9auTYdbUWBpbr8xOTRLiRZ+hQP6DNv2dappLOx+y+zWMGOO
/LtvotbTdsjJ/c+ebD7ztAI9j5CWa1HdNRc58cvfPj2YLVax+6PLQnuLkwg2S+hf
JfShuAyi063RtP/dHNJ12RSoa6nEAESzrzePIvk5mt4g2sGCVOcfnOQgfdZFAMak
5DJP73SYOw8ZKeZpiI195UuRB1HOp0MrFGtJC3xs2fkaJewluAjKEKUTNlr3Muqt
VVqxkodCRrGt1uKm/yVvjTk6kMbu7Wgb45oWGOF2zt1Chc59AtOH7TaQ6vhM7v3Q
cIS3yTOQfmqyjVVs4c4BCEihawfPpQ1WPvPQQTgKSBArf+dOR273QY1hWHK+pTrN
bo+S28KKlRiVlnIK3+T9QF0p+MIAEWVUTurQlImN8FyeoNkEUuCdTiPu7dVHVnO4
djecCCFcrQrDDd3SjIElzgSPKc8oiVD+VL+wmOfPATSc9RVJp2sk2gGkXuG/8hFX
673nT/ynMqo6e2H86o6+nHEi2g31hiWeF+0n8HWud9fVzZFeO0m0uCclIogO+o3e
3uj9fU5KN2sLEATbUf4A6xVt5aVvTvnd3yg9vBaoHznIu3BxvKXvLZyIKjhupV4C
xur1KTcN4ULRyyoLOWJa3/xlkFqbL31VXTNPOqhfZVjlzDT4N+eVUd9hPj9Ivu4o
LUghrxALcKiDU6ka4hFpi5sz6RzsZ1g2f9ZbRR7iXXKCAW7J6DVv2/LpDkK0zCeP
zNX24agCReKeYCWrpJfds5hqoMZHduE5MmFJzCKQXCzNO0LOOPbp7FEQD3fg/7bV
r2pTUoRWUvvbx+8gq3HDahbKnfjgAx9Ysd15Pddp+oMPJQEY2ybi/f7UvoRkccPK
ztjlWtt31OKgOxRTICJqM3STozZgPTSVS4nhd8B9MBrIObvmb3hJrPdcv/M6QoR3
u7xsDedXhvRrcFcDKacnmuMdYMhPni994aNngCwtbH0Rhp0EjhUj8DeMtiZ7Xhn5
TveEx76ltAY2CWmts0UW3tDNXkBQHthJM+6ca+nF5KgLjujThp7PQ5hyVa2jqBLI
EAhu25SVzhGO/gbdqCMxz+3Z6UxVSeiapU/ANqyp+pXLny7mvOsTRzn8HH6LIs6l
ug1n1OT606ublKamq8cJQMUedhnLsciOGl4mfZFrLlLPUP2ocFlkXcDZ5ZtSGhqe
pm7oikcd25idlAvbt2UQ3nIoMXvhvOEa3JrkRUeAG7dG7qni8DSuVYTR3e/yd/hh
VAg9JXELPE9qdD1QNiEUlKy2Le4WhfFaW3nRhX8JT2TqYERYei/wd19zw8VqPMMw
lliScIIDsNgWRayVhyOmff7Xn32WutT1pwAxKSb1qfjACZ3Yc6npwAnKDagYVenJ
gEo3qWmpNB7MTC4LC2mDOgF9RazNCPiRpCILk5Rchy7CGhxY0wM1wVUXl825SI75
lyAubiykilRAyQzj2APNP+f4y6P8dDqn1cQ56Qf8fObGfaqg0njhYLPb3Dwlfouh
XPVFxeZgtPYQdcCGjpZqnmLQyMRGMoWaxmbJwYl0SPx9BEB5SpEmS5rQi6nq4SE1
L+WlOiNz1LzrBRirnGBp3f5QHY76gjogOk8J1TLn0yG3rUBLAh2Qp43XAvhkQ0Bu
vEBlgXXmm5AdhXyvs291BU02RJ2pnGGsa001euhpIYaXbU9mbvOAhlslT0+xADTj
ntHuspNZx++vk6eJRCwQ6cuU01l0Oh505MjFlWOARblHyZT3Dqg1ekJHlVSNF62y
DPrHhCwa5bfkTVWkF3kdmXZ7aLXCMhOo1Ctvf4ZiOMvsqGCXX6wGwmm9dXdC/zuT
l0dze3Ky+Ci9co0kAffsx0g91ezoHmiBoHCL6OyXdFsC5TMC9Y723RqErTFKWd+0
+3yiVel+XUmLT6E+ceOM3IaT5y26Uk+DsdaLcsZ33Uezi6fvJUXukHVbFdLVd738
6dhPq8WMfO57r38Cp1si20dayYnvDuPQgYDTE7lOF62xymz+hvg6skwSp+jXFkaW
W3dz6e5PJlpOx1RwfLGakN5EZfG5FV9UYRKNjhlUMe5UJKVgZtKECkDm1NTAL2P4
VkygdGKTJp2UtT3XB3c3lGZlnqdUK/QPBS2wSbFHyJIosAYNHpjgk402GUwnLBXr
nk0stnvUygxixENTuLLQnUk4WFq723wyp7VKkkkWPRSI1qwNyW8lF4HXe2L5A1Tb
k5BF5zgEXXgpT14YbEhvR2vMRrjubiX5gdO2qc1wyn+PX3Bwg0Etk/4xlHy0spbF
IYeUDQ2xp+iicp5Uu4pzE2GHu4+8Q3YfLKiQgEhdbdZHwYIgBQN2RxY2bPv515bI
7Hv0CBR5uTibGPs4rfbXnxF4j8pD9pIYcsbsXi3fY5zvuc2saxmdM8OFx+hwGtlH
d3WoupsjuCy3XEQfJAGAHPwvqqDhBHep/6wzQ64SG7QxZxb9RqGa1poZb17EHcX3
uNeu3NwYh950KJLqIey7QhjHBwzL8U5Qxrm0cB3B17EAa/+EZ4nxXRXrauNcVdFs
BBv7Lw0m0XXgLdj1d2r2YxZDrD6zMc9H+djGFNz14Np5aW+BZlc4VjyOzmjrAcGJ
S/Q6xZscSeMGqjwfHeI7AtGq2TYAAkrUlke2v0QiP9mFL0DNtm0T2YB7+HGnfaEc
B28CYpP4Iwp4+qN4XXn5Dmom4yHfH3zmLGfG3uhhpXnxQeQtXkDa6U6zNdsNjEst
mPZ0W32SXm5+TlCstsCd+S/9iumYHT4SoUFxO9iUfnrDBi6Jq3jjOWtZxR8zDDKe
hVdfSgNzNDSR8bb4JSPxJOlalJwH3o6rk8RGsgoYdfNqAX2obWKJ5XTbj6JDv20T
PSZH06Vbt0u9ZqBmFys/JHHuUVqG8A0XgTdDlvtGGGUFyuMu6trVD0lOGfiPBijK
Ds3l3FiUeb+f3wO7/R5Bc8HjHwhlUwu5+pf/w2r0JfAzH1iuBvcJnZtpKjmE47eQ
9cPOkNFIyk+Dp07sqm7FNoz5DNF8NNOQcZlqJF2clgOB/AnogktF1/1/HKQ90UOB
Eaj/T1b83T/LUWBUCQmYw5Ln0m/qKC6CH/sXrhl/sNeOFG3M3ezGW4/7XTqSuKCZ
c4v6Rnk6+cq0Lc18i3Wc0unPqcjW74sddETUWgkqVfggjmThApKOex/fzmxH46uw
OH2rDkNLnNMVapWu1YfV1UIGDBnPubCfPTw0qNMsI1FYwPojiUxp1/HulMCMI9To
GDRDP5O2L0FSy080SKh5mkes9IWRgafHBIRj+Ne3vDZKbht0y30jvGtpUpQYg0MF
HvsnJO70sfGKqlqIMs8L8m0NZ8H8rtPuJU8eFI2ABSAGqqSnTQfMHgrxUPbfXZ64
4yTvKD/VdU+fmXeBxHW4LOTNGM4LciZWwUHAyVhmo7p+KKdJfHFjT+PVCQ8xMfv9
9aCEWBaT5VC0v6quNq6Q4Jpw1kVMyZrh97SDj7rTEJgIxONyJvK/ngk7WEvkjEk3
2tmVF1FgxttidTN6dydrp5PO1pRvHwknxcOaEcWNSJyXEPkjyHRsMhoxRCexoyCa
qX5K8Z6JfXf8lJ+sLOnHnqqxAudsrqZcTjAAcxxv9J2y4lA49rzcFsMWqKnPxSlE
kKqAaCG5EyZEjRU9B70Z9fyx4+1ASk7tgOZxo4GO5SibyWgQnKVSruuZgIL8RJsT
wLEaMPKYtxP2/YgBvX7tKwpEHtbhM9xK83sEcr9py75S3zc/EBNLXo42QKTs07i+
/CeBggRlDPcv/vTvtjsWNT01kyT25dtkyxZJDAooHJ6ZUON2D9WVpr89LXqlSKiH
88CSuPJIlubYMPHxuijaS0lqMcizt4ruPOWk8idGN57uQ0mxvUKXoZalHg0yIwMB
taKdF1cvOH/9beJSv7LR9XxB08zFnc+6bN9/fEw5SzYYIhCPLYbLc71nj9RwkA8y
0gE4ResqBfA290SM1Y9Jc1KZclx+BlLDBCyVH2J+z1xMkkz545pffNRLgGGswFYl
BejAfxd9lsDipzCTTGuHkfDp1Wk/gJZogiYMHU/xywOC1liUzN3yVnY5UF03t+Zm
pr/AohN0x3FCyfCFNOraZM87Q9PbwuVOuzjhD7xcxIsaurc1CQULCZDX/9/Z1gwd
njE66fWY6gKgl6R3IRO1iXKm8qwIKAikneAGLpNatxy3hur72JRl6KN65wlD5Ait
3fuWIosaAACzNg2CVGjWvO98jiyzG6HAJJjlOQA2vo3plKYYOEkKKulLURv1RNa1
ThKgz7Q52P7QjfhZAiTrBM3WI1L7Ffve7QvtYkVnQ2QcV43hZyyO/WaOP15bOMMu
wOBZbZo6/NYcNtVxHBX/QvXYRhSTOmu+WdojOxXzJrYv0CaS2axtzWMvs1Nk4lh3
LIXr/vdGH692HXUzgOK7Klm/BWt1J40GSi1Y/miexhC1k1uFm9MnX5qmaJQOeDnL
eNuUJLqAyKw26YPbnMfOfH4a5UkC3yeCePr9vh+aJW/0gd5FvI09JxX8OmHr0kfQ
ovUDpWdqbE9ir6ghaK+v58yRwUdyCulWyTKPAUIORB71ENs6AAq1u4w2O9nqn1QD
PoCOHY0BTkJ3rJH48L3ECuUjaJcTEyE4XdkIWUECDaoJoQW/PycETc25hZKCIYnf
gb33FRe0vnfsql3Z4PBkrSN2LrgcKvhdcPeVgbfIZz4aZ9U7TW30pQlLJZ0aqGjp
r19MjREQ7pkmGeqjOs2SDIAyDAir7hsIe3TczWJJkSdilKkuL4BlAAI94cgfjG5l
FyzsyVIzcVo7s0OFmglY4npytdrq3Ueo9CMup3jzsC9cdRMoBIQSpYMpGJ/vaU40
75NL9Z6x76BkQkwQnZTDd3pyLIAo9arMPlltWIRyeEgPS5E0RS1OzYyu3BqxhP45
TfLNdjEk8IFnfnOJ1PRdvwwAaUF7EnXOj2LIN7kCeCBjMi1z7B0PSHBCLdzV0GB0
bu4J7Q8KoW6yqibUn0bzeXd+kifgaO6+5pVEw9WUuMmCw7Tialel/gAU2VfzH6jV
EUnhMPBOk+S++UUvNYXn32HXKpX2kceUDv3u4vV+2YTXCCTqxlphBBYdBugL6EEd
faeYDJSl74v5W0561hxzUAYABD0WD5nfpub54o/q5XJnrF7/hQW73NKNaE+gsRhT
pfYoCu+W9szskhrZhwvkPexmu5I4SaWNhPv096NuwC80Yq91HxERhNavdNnlaQlZ
jITvhdtiDE9syBuLQWtqRvC/yGKl6bMhEcJc7uxdLF+7KIyjctlzdCwORsRkGWSn
vyzIRYOJo3yb8C3ztov+2hcsVjDtq1f3PluplVqlQnmfzZwcDUGVjPCNhL/pALy6
VfGqjVWmcWKlZzKmENMMycPIyZqPv/RK68J7p993D89qqUzf6vM4/qbumeLohA+O
qxr8dm/9VQhYwMUWZGA/ZS4VipiuHFCrVgcaUhkkXhsl+K5LxPFi528IJp28Q0eV
HEJt+Y4hCAZlNg4c2WrGgwRq2csb6h4tTRKOflrYSDhVs4ohndLm63qDe3sKoIAR
ztI0w36NJ7QtpL7TPBP7HQvRAd1HiHTLL8T1RIOTZtEx7Dsqcb2BMkzmwtYnqDIs
1nehbjgyQhoN6quXYNL8NoOMUW0yXdn1Hw4a/pbfOFTolr4s5HjcKnhgk4lQsi//
wqM53eJVjrhKxAjqe67+Cknz9/UcWQmLjl5SET8WJdkC/q3EP3avWalLNnmyg0lm
Tn++DVqs6ePAvSEAhtDhAvwhibFckvhY4GmN0iWHW8yvKn6eX9YHkElksr/7XcBL
7/LK6WkvVTW3lMRB7S2y1S+feRtQFed8BbBLbh/j/9ezjUcbUpgPLC37oFhUWVSP
Pdf2NiSt3aYNTBO8PbFian7bIZeg5Kj3OCiqj3p99N3MJcK0AYxbCHRGnixgS9Qq
YTxANKRZNpZWJvfg6pli5AUhrORdcBwe+DEdvS5WCLMzKN7sLuKHJlIiRAVpms3y
BnsCSTH9Z+N6lzjyCYsr2IAd3g+7fkKcd3r2WNa0BV1cEIy7XyIvJ+vUsi8/Q48P
VAaxc8LeOiwvLPWDuewDPByWyo+3ZizMup28106feOHuKYRjuAxVLnWubhafw/Bt
NDhSzw4BGA8ezeS+yPKTddDunJlg+KjMCsGQ86yn+gvZGREHzPEJi0GCgsm7quI1
FHTwk9tDAChC8jj0uogdu8flZPFVUyc9bzhnh6EPeAA+HBu79yc+Miqq/TGyehmk
8lDev6dPwalNa/YGzgvPB1f2AEy0gSGcakwVX3RVgQlU3x2auYVN79j6szrMYx/d
AN+xIc9SoB/5xYej4bzzjPdQinB4E0Mmh3mubWWXl1ejNVDZrc136mHumRO2RaRw
8TaXXnaHuRN1F7G0r8Z5KuLJga4e9hrjY5ndsJyA2P4ahwobginkLOfHbikUDCz0
hyHx6ZTb3VQsv76WO9DUM/JW6S7DcYaqOGywP7gq+HpJG0ke0tz+AW6XLPWPSLL3
Ig7z9vEf+SCv26M/jdbOl9UfdR7PnGZgkEz5jnhPLgDP+4sNAoxnqNbjfSZV5eHG
jsAs0SLei4uzVYpf9CrcKo87VzMPJAmzDyc5Qlp1hYK9oqcmwYamqFADwe+0GIuQ
GWaFN7AhXL69OnvdUgzwDQpVDJieyCLpddnqieEeq+8zQxoWm9UKY5NfsFItPJTC
+YWFHjZGHGAUVVXi9VAI3gDk2lRLH3DeZTtfyo8IrJQR1lcRINqSrKLocJfkTWkK
OAyIWn03imgtzzO5ghinYLZ4FAaiT866MO6+c4NKedAjQhGFFockCww/emwkSPoz
Hr9f790RsJ4m7TpOQBvP0EsSqZXnqgaI8O2i07nBp/E1E20xeWzgf5DTLql7gmn0
mXZXipQiMXv7yiYuCzhBHMvW3KnT13YE7uz5RSu/ddZPQhg3YPGTkWHOt+oKMpoI
hq/Gqz+VicGjCCErJbYn4gxZsoN3uNN5AFomsHqHVXMCYLBUqLCdX1n1ECnljrtK
Qi5pCCkUDtdqwh6O9lxzEvibtyzpbMvi6W1eBgP/WdCD16vAcT2qWYM0JvybjAgd
ZQPPA9r6UPwKlX4hpt9qJjMsPkaxPT4X7hyYjmVlfBfa1YlwANn3v0zgaj62yeMn
AGfJQnLtUL2UQyJNB3Ug0Lm+WVgpKqYpriXNUPmW+0fq5vS4DMkhKJkoSWnehA01
bRLKKe9f4DngZa2CiiOPyFHlTKkek+D7RSP40PLYxGRCAaItLaXSSe2Ps5SwkDtA
AmaFE1Uq9mhnZ822gs/9sSnbLR3FHjWt7n48fF0D/kruH+8vafDb0KJIon0XtdE5
LXI6TOClhBNaqMwCMpP/xsQ/JFenn3m/hAtvXZKyLwgN9+9Mozkq1wj17Nx/Nol4
CBj8kvsSJCcywFkKuc5T2gjPVm8jORUkOooxa0UnCDdejCtsXljdw4WHuNr8bHnC
g5gwez/5FGXxaUAC8NwtEcf9ipavwoXyaosMB7O4PwFDO4q2cjcxgBa3lTLxzJnJ
oWAtTmGaPqNfIDtQHv5P7EoxUrMSDHptGf1XiWmvsl9SwSaQRVcWMOch4S9Dku1O
bGsyXvP2uTmnyLfyGHyiysvCzF8a1XifSCoPHyjwmO8DAE+1vCsArWJ8afPsK6Vy
T2dzE4w7iQRroD7PxZnQ9XRd0/wX406x3fkyENPTloqUOe/yY9z7AscDhJVakkOF
Bg+9XOxvWy6cIMu19G/I0V7U7D+/GYdrxR8XmEhdlTGICQkDZ/QJaOvzOQQSHNm4
/MiJduqy83wguvGlZnM4Az8p8lbQIe4EhQ/U8p28gxjsNC9GefTjnO21wFGZXbqe
AHUfVOuTqSfnFj6/hcCHc3B+2wlARQoF0jHCHJGizjlIAVHv684NPywJG/JXNWW5
7zEcJ+3ehKcNVxDdfeWbuRUM1WIy3LXWjKJU9Ubak2/cMvBOnierp1UvGZlu4I9w
4+2YPeuav6yLIMREcepioMGkJuQThRezi7+ldwLojUYNDKiXOfUEgxwcQoHv234s
G/yptBOiPBWrr6AfzP+5h+jQQZx6jah1BL3iSWv7Ap5egdCmLU4+Ya/bVaFnSl49
BPkH0AQuOU5FJiPPNttAQONEVJCY3geJRqTwnWL68c0X+L1G72sCH9x3dVhB3Mz1
Oa1wmZim6wEnBZzEJMIGmR+Vdh6eDv1GUPsFQjego+bbUgzkDK6edhN7cz9pC4w8
O5LNc07g/p2M0DqxKj8xcJXp8IojSdcXdvAztVF7P4hA900JBLXCbEmAHYrB2aUD
VDJlnC6ZugBoOkF5wPZmlZLbb662U+Xb8URwWCCGB5eRLW4zf+5TIc6DYG8HrKNv
+ulyMXd5iyzVagZmGXRWAC+VQGGf7mZCznR/P+eYGODitM6989Ga251Jyogl5Px1
ZEEmFVMHPSoW/WY64wIMDCAnZbCi0Zn4E0TnlUlIwRa0FUhgz8FCST7FPGdqs53c
ymnjMw9xV6v2I2Cfuck/ZUBUolMK8JidZjDk15HAfR2Capsnn8ntKmnhdHp66kRb
S7EBVZ4LvBDcBwgIg5MNsTYH0GTB1bClQRwszhCD+iuil4QhojfAJO0o0iAUxboL
w3r/9SUyXICLaNm6CQCWbbssDnMAGFQqQWXfF8YHN6JMNqA49WQc201PTR+76dJs
eCvXLhaZjm0YoAX44Ms4kgJdiX4FXqzotLR6+lxfLzeNS9E9uTdo4RAEYXp9ILUF
fztipiIY0TH0jDI2DuPOl8atq5u5olvRNPcgm/Q9re3fpIVPRhZx8M1LNndeKi7t
NWZ1ri92F8dyW76CgU9vFYCToG5LSzyUcC5YyT1PHTrvRbQFEIp0/twBuqPEK4Sc
zBqJ89dzZIFXRyUf6FHAcBjsw/IXwKcLN291lxGW5hh2CQ7yyy2/pnkU/Tad3SEB
kjAy78NjQxcHj1de/zgUnpi2aYjdN0kqdwQlNPqwE79zpQGsazod+c3SRkS16RTM
HFSYvqKIj1SEUpgH1dlWDgye8CQneRDhwk4daVfGN/VlvdqBr7BDPJaBvLjJxwBs
UhhixGpbFrmAXLPQWjcDcWs1mIJu/NBtySVAytJqXUGxNkyKUtQL/OUB8ABMopVu
olXqs3r2thMo/sHQtdj+Jd31vU+Gz5s6mkvTAJjPHuuO7QupEbSzrgIkKB6DIAlL
BXXmgV+Fcphe2av3SURAroz6PoXtJMR0VUz4NA2A9XAiNACrYXzuxRBLSKRj2tDV
cvjWFoVrTWCRIX9HZLIcPirKqAfEnIV1WZpR3OMkvxRKCh5yJJUiLzziiUNLr1o4
zx6mrP4BuiJg5Xw96we868sOeshINkYVBT8VVpemX8qv2f8VW+mnB89TMskzo9UZ
/ZQ61c2nzuQcr0bOWO4BCDisNAmVeXbS+/opkQoakLrJB9yhnRdjl+ZJlmuDgJ+f
Fi6AYS60TJaQhG+zkdCsGUcTD+zI2WFkxbYB7DyIPkuHAf3WrHJZai4tkMK4ihRb
DWW/jNJZ3G6Iueuzzs0s+1xZokJTzLwtexLYTQBhAd0eyK1jraKQpIU/9qZOgbs1
cS2oiZFqXnDBBN4RkKfxK0sxLGFjsJUQSQr8+gNf+DoKAXtYIvA8sjXEDfyCfrHR
AWk+a7xZNuCy069W1xHEKHFE6ECgHafN5v5MnR44RdteZPVlD/wW6cfzfd4yE5wM
N4rmktoBys3lRrDTL2YMSzM3NrCedwpEZLZWmUMsBn6cwknFKzrbSOIzuGgDbI/H
Fu8XFwg5NpcJkBovI1+XK/y6lp5tVI+QqUzBhzATwXM5ELlR2hRFZcUwZLk2qxcd
IMMKzGU/F7CfDw5cwXIDFU+YWk6VwIC5xDP3B/Z0K7eOHOEv2Hf4gsRkO+ra6kww
mjomVZZXiKEKUOSKUPIxH+EAzUtyE6Rx9UXpmUDgiBGoi1Q0PMjflze0VtbRAwPE
UFcNp2bBRJo2mplTIW9nkITXHqUICIW4aTJsHahdoXTI/yKE/3XuuTfxAdIgt7EW
iAipYEUBRe7eui/iEBEIHs/RdKnaVsJjUktQsmba96pZHIJjyH6Y1qay4lZnul2q
rR9JWJ8xq5JScuS/p4M1p0G3PadLWxiKbSPzJ67kxtHJi292EQ9hCGo/Y2+TCgpK
LXtxIhf1nushibFu4/3/B8shwZl3SA1a+3tzyyhH2FgNkDLcITji9RT3vpV9lNZR
R60RDSeVvKvfET4PHG5QYphVEMoDVw0O7nvdVvCiO2KZnGcntRsirxfKIuS/YKLZ
vOgap6SQRZ4gN+u+KDrwEnPNO3RlcZWXnUWmUiMI/x+fD4LSuRxQ9sEmi1dJtIcC
+58X+139GvP8owX3clZqpGwh+Q46l0v5lyMPOBnq9KW0XkZ7aqAEYIvaH4JGMt1l
PFYNf4QaKRAm+pnyeEjNemmbW26FS3MyaQ0BVvd4ZS55XruYaSjRZQ4lD64rm2mo
8G+M5sjMOKc9R19QNbkdHQuUhUTgZnp24flwNdE5ag1tFgwatz0fxFg8Qv5qae1y
A3Cgo7ZEh3wELAEIEcGMFUOo2/bBT8CMDWr/4LhvrTB+N7M9tViCjy0ac7deBKYo
CzBGefBbUAcE9JpRdb85P7v7OG8rUCc47KIoo1XttjJ+N6/qlrpdXMCfQZG/rDuh
2ZeDLET73b4YnSyh+nXVYDFx9iCRvcThLCpF3cJBa0yMZR7EXlELiyqAauvdzOEN
GAuuAofPUZn/J81Vaz3x7HXBA9BshgYhufJ7YGkt4zof3qvzLpfrxFcUunebcq1l
WhUxgjLnzg+esSziYwVZrMbaOzDJMUz4/nxTtYGYuuFpmSab4oNH8QjQLCfaUJne
wdoH7UUPh3wIu0y42cxU3d1xHzWIp7P+g92hDi81DOt6AYeSZ75O27t18MNxUQVx
LlI99M5SNsgN/ubVapXBo0VXyhwm4B2C7OR+aO+k+TbaxrHq73T6xEooBTG0zCja
Uo4qESrSmXBZXs6bEg8aIPOI+5hEniQxWxg35TNKQ70+iHV95zhSir2Tzca0lPla
nXcqldIQgLDVwtSdD0Hs5IPW0tppcz+UT7tccUkTp9R7PpjZNzKAWLGPktsuweg+
ujRfjGXgEM4bk+kAjCu4YMp4dNFg1xFk66DVR/VGSc065pWR2fnYI4oE8HDORKMQ
huMrlpIjk/2V5wa9jO+CB7B6lPVS3qh/j+Z9AZfjky/7CBdhxFK6edukHHpAPdRs
MnYioezia9P3UsASMl8MzAOGoCCK9zq+bZBVu98JvDJj8hoiNher+qLg09TwB8gd
Ec45BvQaLwX5L6AN9e/iTIjW+KEaVaEN4aPqvI3XP3QtFYO/sAtyXE3dm8Z6nCkn
T2ATKN8LO4QbcY+cUVYGfzclGmRenIf5fbLebipY1EweLp+ounMdgdIv7AzFEvs2
7gft0W9qbRvIUO39xjYpqUBuqmzmUXfIiAJx1UW6mW3p+BO7TSFhCEXylzN5HO1u
wqLcBdT7vebKUaw8hkZCU5kLZgmIg1ryAWr4RZnZtm1evMNDnl4JNMXu9f6V4Txy
sFfoO1Mj3AGPgZW7L/LxTZIxgVj1+0G+6LF8n7OhQEx812Uu6I/amNsO5OzNpQti
Z46KZXRigcnelEUKQqhR/EC9qUVkVDKwuBH0uPt1duq/kxcAx4NQ9um+XJuicXuc
VlX9QeRUg5fZVzqUMlrYKwg0FvNSrZAAg+KN7U1n9qsfW23XqVlTuJNIjco1rdeA
WawAkvxsdkBxXMyeoNAkJQkUWpodpLit9/MtRuEmyEMWjuZEHdmHQqg3Oc8EAk8X
Rfe04R6ipo/LzjKdawlGr3KIAv5wrqI2oBgLfBHHFEO1qOWWHnr0WXvVPCD3HGoa
H+RtGn0T9i1mV3maHYXYQkFTd5jJsZFrFgTwkpl0IuGhghffwWIZuEtY+LsIPUrU
V0W4iOrOHoQeloK4SbNn8zd4La0kpob9xlG9pby1BDWlhy9C/FqNZCv8F07eMgUd
OtzvurzuFDVFF3uN86NPnW5nd9aIZzS+FbzlkFKQEeRgwZIsh9iW6texAaemEzQ5
wUwQEXYkua932vdsP/xwfSZC7BoHe16MLuRvAZq4lUvvWDCYufcXgxq5+fj/pHtI
k94prwqlukzxriO8fbc4dacohIbUSIaMAh5IJSGMNmZVI++0PDfSaB4rtq3em33o
AyeFSjsf00/VvOnjrqFecTm0ZKg7uC0hIgsQBFVujjZDu5vjuayCrj46iMN1E8GS
XWcJkABn1wa7MKmB9NwlB/BAC7sgGtooZd0LxsO9+nejVx/g1JgAbkrA9jIv9Dv+
G5aQqIAiJ3sbZueSRD3QjU6zTLZR8UT42+HcKM+HLBWnmcFqi1UF/F61YHdlko7V
mR3/c6otVLJvRBJjix8Se/8X8KoR6G9Qm4Sla2KuDgI4gKzsoq1fXDyssKcek4et
xeZTyYnCtGU4wiqrDOWVaMFfMdijIxHkP6NNlIy/dKQVURxc8EYOonVrbdaIhRVz
NeIuae1q8OY8n2BZm/TVTIgFrpN5t6NQSePIbBnmYMpYWDb4GkxJRaZpckUdSO9F
f+MbR25JTtyBGC+I62pmSXe+3XlkNCyii/6X8VnutJECNK64ROyApFBuVxFdndVG
IgNVE8ctfNUo635cGUOZwJLxQeHlUHrYbOadYk8LoTaU1r0BVTqYoBlZO3QmqXV5
nhdSWKCZHlCgDtJ50BWd7DdusqgVG7iGb+fBOpzBp8q17+Tps9kS8IJ+T6CF9gzU
Mko9Zf778JF1IuzSPSvOFp4rK0KIoaQG7+TnVy8eiyvTkEmeUSFp/04Xc44VPRXv
Ax7jYlTLNTQNOLlKzRtNQ31KqZVdITUQ247UbRtQajWFUoig2dRkMLQPmmdkDizi
1BrvXl08053gKW9r2WmuAWLd3FuD9E1IccWjEr+U8wmv6jS9wuYtRay9Qvgz82+P
dCn6ypLf8dXDJyDU0mymCr829NUeB3lBAcm8kfeRxGVykVG7knOqn7gnROmWO8KH
qi/beHSV/H6J5VzmwVNdVyUos7Na9nH0F3NZGzXW4W4XQwzoOAFfY3ZFtLXZ3RlV
LUsT1eknkrZiYQFcdlb3GFbbfQ/o6igvhtJ26pOXh58+VZ7wuLrfja311vsjlMdE
hCmpFo2pPKbppCudOeYn+Vb8fMQI8lDo45LaySkJT8CFmNA4H94C7r8TR3N5NP2L
539thFuaHpU8EY7qFK9oLsWYqvcubVHQEUhqecesme38Q7Hm56yKzIr+Y0RN98mH
6op24t0NEDaEvHx0kDKuNFeU9HGxNP+HbmeYGHbnBCg6HFYyim/DnYJgiwyDfBN4
k/vhGDtpJAHZjvY8TFWpif5SCPpY3LnR1HuirPfZyUJJh7N5PUt7noMWl5QRdza6
hkvQ2Bhxk0Oy90kRUpHb9SIiEpnuKltj7Mv+BB/PSxU86eKw3Sw/GoMW9S2ox66W
+AlNMfmHuBy6ro7+NPzhg1iiJ2afT4wxvR6n7rs2r3S701y/L3OHanTVWPSNjJo3
LHIDW2D4wTz9fYnUudM3rO7KWop2jzVkpAV0mQildkYWWtsbo8VEx3aB4Ygn01Tu
GXnsgID+K2ENUwR5kNb5ZLLWYWgUTeIDSf3Fk3JUAPCN9F3kjuAq/SdLnqbm///z
amqmQ98ZCIEMPFQxOEsoO/BKxW0P/VemGT4yJIHK3bcBzO/+zsv98x0czlqyNglz
xYdTS0Xhjh2b47DpkjeWHfCAuy1PoplphGu27HzsiTZ9ehhneX7bSq7yOj0sIBDy
AG5nXTTswBVxZxBUbCufszLpUotCJIowWi2KAtHZ8aSWKsw8MdzN9ekKrCVanoh+
51vDDvgcHQi55fmTWjG/TFrpaoQ+UXZ4suObGmR4wdXynOW4xthLJMTKTDZuXfn8
zar7oyg1qLOfRmf1dx2174ZWOIkXKk63/TnC0JoF1NYa3//KkKzbcz0CsaACIqXc
+SMy2vV7WuPcY09klsooYOVuXq4V8uYCrlk4qyyF12C56TgZN6W1YhKk7WjFmnEU
sf91BWp63hOAuC64IRgvk8is8BiUqN0e/+I7s2eUQwg2OZWwdDxP2O+JZTqL0Waz
aDfZx2jmJIUqr+4jbWfTNRmwuACuQDCtbFQIS0T7mYfOaU5srsmyyRFbp7n0btx1
Y8dzwt9R1DRc1p2zd1qIjX0WGgrmJ0HAdydpH7soIK/OtYG/rKMC27wGRaOw1p7y
SEgof63d+J+7f9+v/zzjZzK5Uhr70O/d/tG32ceyqdLgn0XV1hCRu0tSw1jH7Mx0
R2pIQWxqCy0MiLRF9qYVIkPeiQL+EakGkgnGeLYUcU+Lv1IBlxY/vXDBsHo7kMUx
xstCarPz1Pd2FHSXfJQBduNByIlUtn81COaDQltY1Ya/SVSP96GwB8yIQ43oNDT7
qlF95hWuVV2PhcUCXh02CDOFhsiUISPmnMJ2LbzxHbQ6trKBKMpsVYp/Jpoxydbs
ZHnkXkvHb8VfdzKeA6DZwqmipGU6Nb3qGtZZRr83aabXRHP4wuOiuODUyZmK/nYi
cNQofsD3nIAOgrW5E74CaSs/6tcNktWHMHD6N2q50tmljCKbfvmaq9KWULtELrc0
kU22ZHHZT6pXoEFfUEpsI2gZjmfCOufBAY/87SxkiruyFtW9ZIdWl0GDR2p21qQn
ywg5IFAUzlIlbU2/12Qc+c1PPVMKg1qScv9/DZJiFVoEnVWvZj4yEGJzWtzqyqJl
oEWrYbB6+rFPnKPOMGagDOoapFLoUs1Ho7dseT9PpPOYJwouwFINtGDaP67+JKm2
Zrp3P3q41zesq9YH0nNx2DaI0J/6KZHSAiJ8VEUCmGa9McUyKvJiUV5SA2HcE/YF
yRRfgjKoKVRZC55kMPO0YMIF0IyT3biPxYsIhStKc/vRjtmkTX8sDqzwvUjXtHa6
/eo/qQGmVq5yFPK8Artky1DAHuxiyFyTFIsz91yCOz+KhGFlZUR/hScXhXIW3Z9N
PVQxO9aL0zksqYiVsbsHylmJtuSHb51r9oEmOU6SEM1jNxLx923N+p2JfS9xJkxu
fwKa5CYnrafp6jIit/e37Wf9y+pIfMUCk9G6zN3B8+w1mnlnf4H5A/1kokdHSm5j
wUc5M7StIklCcjQonLoeR8jmYOs8m+5gIjMGGqdsvog/Dhg3LbixHISjkYortGjv
g+RVyD+uSmzGGo89HhivUbUpQF6M28D9LVDG+VSqcPBw264mn6jhFGv6A2ovnOuX
n0y8Vwu9qDhQBPbDaVLv+5AaMG4mfLG7gW6AW/14zlDoB9k6V3ZKjt18qYXLrgj9
7dGhjOdiyIriKfi0pQvNWewQhviKkfWaedCPmj4iTOiia7vyM++ngI7/toFn3WjQ
ODGg3x2cHie5GIIRRki9v5nYVs3Q68xp98u0CTKJB/fl1Xy7njfCgZ1iLLKV1zHW
RPVJ6vVUp3JBy6wlFzpukPb3zbo99iEPyUd4eFjiaRog06DLiE5YA37zpZaAXHSZ
Nxtq076V226O0SxnCrI8A500zg3bxkHQ3+g4CrYCyaK4ivq8WwVefbbkwrbl8MG8
s4qsA5BQBXBuAyB2oGbAz8RrI2yUhQ2iYfjnZiohtybkWqHlphgiznG5zSqhwaSK
DlAmqxDrxgVxoMWpFMQwYScqdpi5VeI5fXhatfeS8tahro8C0UYpwYcsnvbPa4Po
hNlPugcqzSPynzm3P/uuPZajrwzXPU6e7ppHtLcG46j7uWSd3a74+WRytj932jU3
mvj4QL2tX4s1VzB57d0IBO/NFxNhG+at/pM8tUP9mcLUdpN+motxSnYHYLeQ3mgo
cbUKjYyiMjqbqj59ku4/YhLhxZSHacIMTtsVhutGEftj4JmTkap6PhO4AMJQaT41
AqcxMH0y319vNDkZmthxeMlJ/I4lY02AyTwgLZXtufCIa09MaKtQJTLISHL2fLWc
GsMpOyEsgfhVt9pN+viYKbR3PSDSOYu2G5GU1dSypP1VLuEztXRhPpeqYybAsQRi
xPQ1Krow7N5ZCsz4sJOyh0f7kSjC7vcsqTXpz2Xi+R0FD5lfzf/ZYSdcrOUMQJ4Q
n312wVcqJc3Q+80wSjzrdQhH9e4j68S+GAY7LDh+y3LEo8guGWSvjoNEe2zWwdRt
DlCU5Ni7kQmiL46dSWKodNzZRUuyHd6uG+G/jk0CzDsv+7fmzoMuyTG3tNGsXJbE
4+wDVgkvLREFe2KiDpwzaI2F49o1PoW1K6u9awh+pnbqz+B8AcWzgyaydek5qhwW
wS5dQHNcQHrBm0GQ5dcJESfsBJsaRKVGvsVzJ6eUzNiYNzlP1JRHw1Z5NfxX+Czr
Ub9Ar9g6CUkGIr0CCNjFeCN3hVrjcz9ja9gspQDCyJcla8LoQ1GcZgPQ1PzFKObh
efm4WUG92l9yZtjqUD5pZlr/0n/KDPKRHsvLa9SPhqAVtAvwH355a9lyZ35Q1trZ
YVqGxkypHHixZwSfmTRdrMOKFU0c+HHPQcbnT7maMYIpUniEEaPRR6fukgoXno+x
OuHHPy/lfiStcXeksX8AMTb7D74R+yLK8Cjx3W9JL8HhBgBcAP60vsW2zNiE2J2O
8b8T8WzWzFBR2sswtooDbsh3yQuLUjUZc5HK7MOydYHO6zAGEw2lBmfWTsv9Brvi
LGsFD5H4Y2m3k2NWbpXzHpsTs28kr5AvQfqYcmluzak3i6Rn8IRFIg3lurNFE57X
CPINOe4b/d0aOrqHsGXExfpbcluTXJ5YnlTP+k4N431hto0yuDDpURgAodSGInQA
/RhAri5U6qlUzXWFLVFQO2bXN0J/NttZgoWSnTUFm6pShbbN0wK3wItXqRi5QOxI
jV49wJUc7Qu/o0GJPJmpMF7YSR/08cpGRFVQjnhcM7CIlrXUvV+VMrZJjs2rgDW1
K0eZfPjnH3g1GqHl5U36TMOPIyRWlPgmRojtKY+ojIjd7+OWqmJUmp7qqVNQgQOK
Q0sxGFcA6RY+P9VpVS6ZBc/9TqYHy5aO1P4/VnmQFRYnlQ76CYw1Q2Lc/5D4NcY6
me6ohjVI/o2s3Y5n3X9L++GUN7i5Jsx+zm6Ag87AfKgYdQnQ+SlbicLFphZGBy08
6g85Hqp5zQrlrjOXlcU22M/T0PrY2DOYkNomHb297ReXMNM1HwEk9+YhSm9YecNA
43gJ+Yl385Wv6ssxVcYlUFEDLlAMpLOAWKfjmXlnc5FhLGfTAZwURW+YlJ6jDIIb
YwxNU0ZqFnr8bysV9kB501IjQbDibatTI/BzYnph4xP1zuyPnoZfSY0Wp3kHXrcw
cNdwimQlMgRCB7bL7ichSnA2vRSj5C8SlQ3ewKsVysibdjMI7w2WF4gxIEvKs2Ui
VeTFpszhOy6pxGbwqka1XliCEWPyo/db59RhP6wP7/qjN98RNVC8ZjY+fS46/Pl1
0Wa+wm2JDD+XG1qagHwsdPIqzXUJNLy+DE/IQW/vvuYKyAiACwMhJYvOpj/g6ocC
8JoXEnL1q27KoniCAw7nW0jir8budz5z2Cmp4ukV25TDlLaSthCIF2wSRJazHNtH
D7aVsaRc63U2lrRlO+NXc4gHrvSCxMazJ6s9NSqFk706711NgwOEtmjE00nKhgya
lJAh0Ynk/M7ecyE10wiCMSpEfdtQb1TeTeKm2xiL1GtHonmmN9BCDytgJxGoOxao
xFDSkisYO8jK/azVao7moeh/ZF07x6EOk+TK6gd2LohWOmI9BH6dWuDGodD1tG03
GGH+zd7biZX19TRY/na/kRtBNNo91KlfKgZtsfnHZcqQKmhY6yoheQsu5petdWWd
3YGdGHo7SYjdOQxmcKLxuNPzDQ50vmYluOuQ0+Gn3j4f5gs4UKm9RaiDkLTqQSZu
PBTL1er/otcFHDLAHk9Hs1S6hem301rkp81Vx7D06zDi7U1OaqzekTf+FU0s16xS
3L/4M806DhZn/dGFNkSMQlhfeQBpEvkNBnvCh8e5SAdXo4k1Qgh6WvA3OAcQ29MZ
ra/AHJMFyE4QK4qx7HjvalSJE2v3vBZJgfFh+auDQwuQ5nR+3ynvQDU2vY1Q/4wr
eLroWsnOEHUT7XI6su+Ilt7G3weyNq+OXTYJKuiN8kNy14Ogrfg2G7/HryZ3pg6K
f1m84w48b9dDCggFORrZfM4nZtXubi/zahIsIp2c7tRp3bMxxHCum54acA6SbRmQ
J6dO8+DG8tLFbUqLzfBHe04T3g9hSJw5z8D0GVDDTY9kzL2+zFtj40FHCz2w8aki
RSlX+4PzzOpIvhPEQECLPkjGrvsQK8wkznBry4GwunGI52hRMPgbVBDZK9KqcV4o
6PGw4kKHQSJNuTmsHC0KumL3tX5eq+pDKqq9mCeIOWJujOsn/+3EHntOZWbqky0s
gDeVwRWOAYalr0tB0mh0Agu5p14f3HIVutk//eMDTcZVR3M2D/DFjlqGKshUOruV
nasBChhu8gMKfC1OPOAHNL9eFGK2Pk4lsnHBokt+jcbKY6PT0l7fFsEx1pUm6xps
lUCb1q6FwDnrsmJBfSHGvx3mM98dTmNXp0oRofvKhDR4aw+GOUogQ2WqblJ+41rP
eTBm17YoRRL7C6O9t6/vgHkQ1OlrRKnFpOUTJCuolkJtPWKgZfsxTxjourMRExWG
ZrQAddviqolUaYBaTs5hGoan0gB7gVXPZyBUi2YEywhYrHB3Xr+BRdpXMaEfK2Ou
fI005C1i/TUFmiZ61retS3bKuoFrvLRGUBL5KVKvh5NGjFg+gSFJ16ugYivSS/Cr
GdvGWDLqlezBfx8Yoac+HfmKDnmmjLu2ieap+GziTCJNQJ+J1viPe+Q6uCuujCUd
DlY4k2S4tNuv8VYYHv324kZ2H3fbME/ccGPMFOxsJ7uhHVL7SuP1JkuoDh6zNgNU
LIo5UUF9GsDCyfqPhVEP6qhA09N0lBFPEgkJAUiJSGo2RP3Gq4O1hsLCkKRfvpIv
Ex0oqn8HPZf6NwzTT7xbcIWDdCt0HfljdegkM8GBFBbzoIEV7jb8QB+TNCUcdxaj
juq64T3cmMRPIRjjGksdAgOLZ0+5Ta0td1mCBf6CMGITWFnmNKEC08+K2eSVEVY6
Vk8vqiOpzhpByGWKAPO6MTFJD3nJ3HgEbgx1/JprdGXwPhcwY8+QH7ELCueev+3I
3vCEvfzev3Ic1BXxPwA1Q8IxzTdokgkmRTm6c3MqH6sySO305RPX+nh05Y32uOjD
UzjRrLLARbg3JQC37QjHRAxIbcinztEdACrRcV2EXawGPajvHY+miqceOG/r6QH4
l+tR0obMXGS0Cr6XlSP3IS4WdhnUzHK/DrP5OBf5ES6VYDne9IbbWmsY78Q1zoFt
TG+bacZVZ9jta48AC8VR5DsezcTJJfzOlamhTm/QC3B5VL28Vky9BbKd+EeJJUAl
u1eq8Bb5KsrZbkFzYeL1LCqW1kvS5XWq+Ntf17KzDg6HyzV2zhsWXVg3/VXnjTzI
8Er5BewVD59LZHep46yE8xgzNVZDpnAqbLBcqxoCKl9OPZ8X8B1gLNPQcc/v8TIl
XrCXqoWr9Y85Qp9xOyND9GafRIUfmEO/i8O8IFuKVOv2aJ+ML/QnZUmnoDJRTMve
4/WDh/NxpUOKrzzvrAFQqSyk/piwVUJewUpmApaM/jOZwUVHvTMb8vrndsxe77bZ
gcbqvQvGxacWxYmI4thevdM3IGHip0m57w6dD/QZMO2lCuDogTsrxF7KKkUe2+X7
kF9HNWDEuz9aXiGlHnbDyiC1xPMhJvaxZZTOSk2M6sV7asLld/ghya8R72vNIYDP
nV/EHOdryRrGAr1EOnU9J8TcsE9ph704Y7hFgvd60nlHqkJy1wqvsPBDPokRB6cg
1psbBu+GLjtPDB3hHzuPaZWlW+a+yak/f81TVvqJKWPk1B3Z6WvGnj0RoLNScqgn
Z57D4OyndI3k+2u0KAjuCpvp9E8XHUSmoxQ9KhjjBTBBkGqWZSv+42A+t3F3oQ6Z
jdX2zhAQ8BwqfOlVNq1kccyCrLKy828Ls0BF64+mltmRDwAiFRXrvhcsVIcfNh2M
jGcYZ2QapnDQXMFwoBATckMrzRfdQXyZQ9akb+I9SeV64wuh2MbpS1y3kF0eb2Mf
GJj7HriK6WJ9d2izTnfu8Xy05FrYsSYtMvKAtlY+NLYbTtPTBd7lxZzRA7J6C2Bh
2Pq+c1zv8U6vbDJtwmVPRtLk5D1J1EV5AFtjbxVYJSCEJoJ/BYK755ZGUoIoYEyK
piVWFxF8SymyENDrJ2YR4iOfXc/q7O1V3Wue+RmWcJszPJFYIOQSzbaAhq1YJmmg
O4ElG9LG2EPIQSwaVXw/I0ocz1l8x6f0HTscuI3AaCtfOtBJYzE3i+zCPMulbiuo
cS1xPeICJP3+ZNwYlwI5gsSbjjkvD9sNM7xh+lJPPH/Vb4LbSbCyfEbt7ePVC+4J
abskFK47pqyavJC7VBkHRd+7DcoNBtln42Bj5T/Y02IdFpcVk3A8S/QpFEBJvY4A
G8FDRs3HFeVHHBBpU7drXdAvPrMSPHJPxbYAdOG39cpeyC+Fl20nK/dQbAn3zaal
3RoOgDgx6n9t1Vcuv39Iw+MbCWZm7O7J6qSpceDc/rIxEdpW8juCc3Srf0bSAUtT
6xCfARwR4Tq9g6DfVKCO43tWz6YDVChVQ6GMnANfCoC9SAUiQJOfszuMDuNb+6AB
0SHFRqkFXVKVfDiRTvD9p7N95IGWJBJfYU38m/MmDrVrpYXtFa7o0PmSxSY9OkOt
St6IJKG3/GULdb+rewtIjEV02ePRpY0kXmEeQJjZycsKaL/Nz3cDCqm+5fNicZBQ
DrS6+vP9CqC18o39Y4aCtf6BtPSMPd1kdlh91jexYmobjAsruZcIN5X3h8+FP6Yu
Wyp6wiBThl+mcVq8pwQ9FPrTWDwGvgE46k/FC158CAmJhIZ0ZXsHxwHOCIFjuV0b
1U8OdbzoEMrWbKXgq1KqqZPUx5/8bG9mRsRFAEqgFs0ta+admiBooZDmLUnGvJXP
E4CDR98H7VbkOnL9rdLuOE0k0nSLaH8OHX/Gavhhls/xQcTtmdq8yK0t+dHmRETN
/+YSEVwDURMfX1XudMS2aOG0l/3Q4gPde6BhBsp609YP9M5/BieGQLKyU3psMz+2
cSoQhbUE7k/fFTZSuGx40afqye5z6PRKWuQaDGFW//+6/+j45973OU+Josi1YBvG
jwzF6TuHhDfhApEGFSoRqv+0RiLIlqCE7/J4wcDxTsI54rIrbWTUIsmnKjtI003h
D9g7oQDv4KvnMSK+AhlxK6gfUssP3+tMnqSUhMdxzfvTfzY6sW2qzGpmQTR8V09E
D9bdDQAbROiBSCSapjyVsjwLPhAPZuMWoHDxMpQl6WmjBCdppaO1hbQLt8Y/pF47
uNBne2E2esn7+2lsKoyHws8JWaB3rNvpisIFr4HCOTnhMSus1o13ZS45oF/q1XST
WIUZEi9isPWj9qU3inOANs3OShbggTSSz2PEhT9V0w68uGuq0KBDF5fhlPanXl2j
YdsBMA8LFsSqEnGhKr+mh7eS11Ud/fSHY8OiPBaSn0l6pKjBLZA1qIvX91B04v1/
/5nDVmQ1VHowq7lQIygvKG+4M7wlq47OEGWunhg4uGLcmGqJ6B0zGtx/fnfUYopS
PBLvVVV/u1YAhkdaRY88qfe2CZu30MXjBWyfLjExrOXHjulAz0NMoe4nB57u/7jV
4LjCUdr5x6jrhZIovouZbl1DG/IKG2uYxJRUg+II6+pFvysyYYuKwTl+85IH4TLF
lXAKkp0AkMYVhJN9vQl8aZ+rBH1Orf0AAztgM8i036ab1f+6ws8I2S1nacJfd8qF
z+CLm88TJuk7b51g956gmW/uAAR9rmaSO5s44A2tolevRN6A3CVOaRnTpXrmAtT7
qFDOpQIw/L1ECwX/0ji0KDKR2diDygtV5YNrFBPvJHkEmzhp5knfjBLksbjC+cOO
jW95X1j8i4Hlb/A2qpoM0hvvv0T7uybbysYDpMu5hfpgrmh7UbrIrFBwHfaGl7D3
gJAZAW6NlKQaS9rwirDMdFr+axMapatIzUj+cGVfLHacVifDPfOXL/L03K50X1EU
1mEofB+nFRIK+d1YTlVmzcnSafnR7QJIYu92d1ixkajk+9HFlxOc3woWvSL84hTH
ciBKPSMWYUM92nlWL1Q+wc6jhvr85npS9/XCtMx4/Jpg8ydN7Tbq4Ogv5hrS+Bdd
09rsgNSWYasVwAv/qClIX75/TQ/RWObyJR+oGQciI5VSkMk871dDzvCe7V6Sufig
p32OTkWmRU3GPduppPMLcUkfH+XNmzUGiJzBOEWSZ9KpH2NUUQVhqR/SO0m5I49Y
c+gF8D8HRm4oqniSiETrN91fTBqKVu1kvfF+3JcdsNm9HSgiyyYJotL2S0WAo4kA
axBTROaysOlsyWBIauxXz8NmdN9itXvVd21BjxK+PRh6UK2r3Qdycj4a/sf1My/+
EZQ3zDEvZBcw1cwSo416tXWu9R0vVyguCvvsnlDBnQndv6bEiOSvHnthgzcPi5Ey
qgByxH9BRUctHbEtIL5/+jnr1lC4Lx2eZraB7MBdZdYrKzkzVB6bRTj0iWR/l9rF
I5KD5qI/OE5yktdGMCgl6OQT/i7uPsCFJkkwXCFB6kd7RHO/B5kd7vIwHtBI4ct5
Xm9zkwcgnb9+DPjhdH4kr6DtuXgSnEcIayOhMdHnRGeCS5j0VX5N6+2PNYQou3IL
WduGgWHUQy76JbbMA+CtrEFwZF3MaYPyS6peWa3RUI+DTugA+pjsVAUKbfU0/gAz
l1ZYiGHxYR/hIBBZp+cyLzrykxgvUKOC7pkykvDfvvqEn/Lu6/eEgURcSPLXLh6g
jj7tbZwlU56jf8yLH/yh/Xx7L1LW2aXs7AhXCv4mqyufqb1JCkTz6d1e5HYKqi0j
3oYqxFs3M60asHRps+9dQei3ujs4+9URTINUh8hGOwapkPHVwSgTF+mJicsepQgJ
UWozTQg72qTjxEbDcD4KHkQgvzSGEd4F7GR7ciw/jhHlXiBayhi+kObnqNgP9Y7o
tPJrlzHbtvfSCIkWpkL0RkWaj4x3ZU0TwQmTKwdtyOdNXvsHOe0kg/ntcIO6nqgX
b3w12jQJ4i5qVLh9bJtvdZ0447P16jbWiw5jbZP0FmIDRUV7MUgxTSxtZl4dDVXF
UVsT2ny6EYSUu48jU1/ddJE0XxayAb9qt5XUtXklJ9EWjTdTtehepCD4O/l2BtbY
Tss7rzW1BHWHtEORlvvrA3voWXtYW3CWCtLcP8RnwchnZNkl2GccW9zg1ygvDNcF
+hLPkKQYy/73UwWlVjM2rA15s3Wp5qtxiLq04QLhAthCX9aRlnW+FMDPSqO4Q1Vv
yKjEoIfPUSTGgXODacoNVzS7/VHw4o525uzRz69yWBU6cSKfadkv/lzumsCReiEk
tlnk5fN2/7ieygdPRSqtiO5tYS/x9NMxHkn7KgILpbFKPy5okbzQX3MIEaWgSYZZ
dDLPoafuou67Lfb9zSOkhlN6CQ+gIIxIt945s69ymiEHA1jjtK7VnqWMWYyEPE8l
z7nNs9oq8CJ6thEk5lvnRWMrWZTRp5rp80aMd+C0dyX0yPtJYqhztL9l9Qkit+f0
CRYBdsIJqgmSNXOJBj7hFrwydsuA5Q4NawEm7hLQMJnHtRSXnEcLnnpxkEWmUIKm
KHhAZN0GTk+GX4IUR+LnL/BBfEVaIZLbdvWP+nNE5SI8k28HsRP5lyuPml60mzqK
7qhYwcrwCnljJyvXIdlLjmjX6E2hg/8zU6TKcB054lDa23XdKihtjo9e63ncppYL
69DGXAMrIbFeVYqBhqcRMEdPYaBK0CTOTdxh0838iX1+XmHKJntROTx11xuARtce
XoxZ1s6vZXcOceJyA5v7jWpBLIaYL/MZShFOdzv1wP8ZcSMS9JPxcj/U3dEMxvIH
6SkOHv+7Wk7WBqp1Rp6w2WqdTymhjGwF0+LmedLeG9PkeFV/dLsg9VTykBhE/PMW
55zhRDl6ZqzckE3aQrwMAMRFu5CYEyIcFwyU3rh5dEfBXhGnuvhO6xmXLzBdg+Yt
KEuyNFJb2N5DSXhw2Zm4XFeWQePtw1kimAXaQXArBNfncfGDtjQUS2DI3ZsHHtZy
HmOmd3d1RNbvudRKHmJo3GSRjuTvItNQGKS8AnKl6sM9yRWOhlqRU96sBeDRw/q7
JuIamMmVYFQbTXoSEbFSOSWIeFiD+3GRFJSwcNN6xGxQx2TNpeTEOscPhqbvyuS9
nog0Y9CRLOzTEyYAV/J6v3M+oewXmR06SxV/aET1Tpn2WP6JfbrtIbpBggbPta2U
H44AM6x4DiF23QfVVGDeaUgy2jM4Pq/WgvTBZ3QqxDG8URBuxZ/1Np3jHmYsaIJh
zrFcMGcMmy9DqlkUlvnKeumAwTRgeHDtlSQDBpEaccIkuQ/KahS6x0b7A6MPG8t6
cqbXbaKX1YCaJhaY1wmeLYIo6KlUOw1Kg7wAFRafy17LmGf25Vov85xvd6Lxoflv
qxn5YvK6uo3dOSHy2Ir6V66ZpZCeAVC7GMmGhzKkSfVE2iJ/a8c7zhhq+BhkmdCH
b/DW61DDzm6/VS0q/JL+1+i57RAcL4W6AS3M0+sM24702QcV6Dr6ViplfGc5+M7L
baT8ZK53ZNmzMSsDB2rmMYQOrerO7y3Tz9UZaljGI0Sm7rkk2g6EI/aC+DRYbwRn
Y+jUzwII3UxCZF1XHS2FYUqj/T4Z7Xk1Plj8fZLs9+ymdzHb/WflymPCzgJoXyFx
AVZ7ux+AiFseMmuWAosG/IwV0mkcTq4OX+0hvYOzIStq4AsDtxGqpJ+kA/VwVcNV
AsQbPHJ7VZ2Un/wTqadcLFKjw93x3usu41Jng4hy2MIdxH1lsUs0ffIKPAGH5Bns
2CpMlJWIhwG39U18ww/WMdnL5JeOs8tPcRXyGQKfxKv27Bn7HIggqW+TZ2/4wKpy
JK2GgVEeLBNA5ptBAiLzhVY5F1KqRKrhr2nlfKeyzqkwT4f/Wwg56GIEJtqlQ3FF
o49955of3yL8oUc4Hn+djW/cICkBvQUmY9smuPjCtWLWEHI/0BSjAhMOTHEtIBSs
pi1P4IGqZXFboIDXZ+m19LfmYk4a4kLOisLTeBDG245QVDfNPCXsAEmteotHvT7a
Ns4lJxeU1LWSHKUvBgJxc6GNgzRjXcwLQhlkyYO54NZzqie43te1IbzNdc3ito5r
hvJZxAy84fYWV9rnSg5kekS6ELWkQUfGGWHGzFv7IicqOdSzXr3XzYrvZFw07JVv
3rTOHztZ9gQ6SSQjBbR6VggFK/QeXg42XTtRM2YAnpZ1DHeO6Gp9tM3R5I2tUoyb
gpNCLHEClkoo7zYiDM/3a/GFXgUyt9P8nScG5kWd2+Y3JA9R5AbP+uSL0QGIY8xX
dJ2G70QywPrz8rkJDAHGDd83oI/IxpqB2ViChraTlruuGiMTvdcpzt/1qiE1c7mK
8KnK01nfb1ZtGb5HNVCRywOrxDX5G0X5EiIP7qj0HGZFf+qqME9Y1YA0va8g7Baz
jprD+X3ofY+H9ZJpP8lL0GsnMi31jK1Kdiy4RnM20zCc8sRzz2cQZpnyXXL8+ZEu
o7Kkv/jjhZpEKfHdlmmItmqivUO7naDsmxAFFpa/k5tV5K6b4aFNY+E0BuhAy0vn
LKciOKT3qLSTmdhkJJBEfeRI0136ufmA9xelVlyIJAYOarqJaQNhTZLDC5I6xorL
sta9deRK9OGxfccOxdjobS+vpG5v30u0sCIh3kqcNLXXUHaQbdfFaKZVUpO30rtE
VCZo9qHlzeM96itEq/YuTuVATC5f6jBQWdRj4mVNxaKm8jCZ4tyfjtokU5gyfvAW
YeeLxXMeasrHnNoIc2JFQ3U0P6jn0GXmWClKfn9P1sCZDd4WxR1NHVjia3Q75nV4
uzQ+6u6V7ofR4bWSclWB/OxNXUQh1QRHwFoGi6071Jv4QxTq15sTzSItHSo3bT3u
kiWPtRrnkRqe2R9YB9Aq3HsqZQYrw188eiX+XRKK63I+m7d5OIJvmXAXjKb+rYlr
fqae0py+BKrboQYgmRxyEwImJZbs5dJXUXF4WnHF2ZaTyLGcpGx/Kj5V7jPW58CA
cHSLwmFlpublnT/1dVlzzbmUr8zusWwQQfLN1XRZTMyv1aaO9LsQa563r/lbqKK6
YoozcSjCxMgh/5UUhPDULrhDaUCnr5nVr15C8sH6ySH7HPGuP7KaRIh2sgbnNTqf
3FoLhEls3rWdWdIpkxBqkrtDvkpTnkCU57Zh8MVct3PWXxH3+InrcFnllCpxxUre
8rjG2oQpGtHBg4hDyoeYBjn7Ls8a7lllv21oFoq4b2Sl5lI+xbz9RnIn9IlZhXJ1
4NpEu8xlbA/TGYR584f7d5uuGhlMLkUp25O/R9av8uzr0mIBNDHoyBbfs39VcNsg
PbNTjyiBqLKNHUsmBUub0hPpZ6Zsj+BykW/VyK4LT2cVehRqYqveHSxCuQDEvWGu
sQyR6mKnVkQ8hLO3tNuVWRj7IpUpW+LjLav8q6HOVynmWHy28GfkQ7lPxCh3gXn7
vdLtW+OCoUI5w+9jPTU1o0DinepzY9PXzZXtzSeQf+qIy8XCmIB+0UXEljozvE++
aP/VTBO2IqBob/QJx2yexi9MotQ1KruPbzSLo8nPWeKzXiDejVKDmOWvq6Hidj6C
FmYqTdA8GeDE6rCONir0DidmHzsG+FEYOm/9WL84mykQxNnX6bdwOPQyrvxJITWW
SRewp66OXNLTVs0B4PMxoTIhobGZpxyjkZMZRVnVvbyLKzVftWrxcDpUKRTCyLx3
p1Nlzx1fHE4a6AoceftN2mQLEGN1hcmgjsyznL9xB3YozzLIQ9S3rA07r5erZ6T/
K2UcjlsdjoMTbxU9b78DsYRyobmX98UWuMt79b8zURhZbWf9rUy2jm6iolQKWnEF
AavmhdxtP/1OClT3nUcYfgNnp6UvIb79EmFULF5cqUDQXCE7hmArCJl4ZeF4Zb89
sRo9QTDGurAePS/WwW1jfeEQ95r0JlnCpvre96ZMzaQtg2GRjLfB6pEGzc+ynGbi
6CckU5vEowMOKouUxT+zBVwdVXzdbq8SDTcen7I9dAcxYg9NXXwQnYtiDqXLoCCp
FY5wqj7csALVU96njrvY2PucaPb0kZE8T7T+KbsqQrM0syqu7+/N6Ix6qY39G37Y
KtSmZ7e+lkxomwuM0hHrfD1anMHW7V0qALtTYGuhHsXzV6eYGI5JHGvf0Znct8DY
tPyLfdmbgZhOMUrLUKlANdNBpRhkoNMv5Y4oR21xJYeWff6rCgOP0U6j0rDLfg+A
UEA7Ows/0Ej5gZC1dPWVUJbcOGtArmEfs/ChhegKtP6YaKdSB7nflEn76ESEE3GM
hprS84AAne/hdichpSsmFPRkaX76Qu7XOA9uBC3aqq7N++suHQInjO/FJkQWm0iD
OgevHgJmJr2UtZOjQyPavrNxWurrgWXhaWPT+x0mcpeyJx2e1tU1a9VOpf1OufzR
6uF2YJLgPA5WNG7anb4Uvu585NbFkeMe1UAY6OOiTIVfYPzdQEb/7oQkY4XzCa3d
EXX9mh44vIuaMeW329mL5X3hWvHcgsd6+fR9GMBFjNPsvmWB5VP/CRxJui9k0n6Y
K0eM/aHRq8J7/b1uzmxBJjr/Zcno5RXBMb7+2Wfs783l1uorLVQ6X9L0SEZ+7Edk
0c0nk/7URXs7qm3PUJBxPleXboDTQSG8LGaZYyFkVKECtJftKv2Lit6WbDB+xbYq
oBj/CnE8K4vJzRMZ0Ccbz+o5p6vLinDrP4Z5GJtbiSY5etZZy76+HAO6bfnd2pl1
08CDc9fERC/2Yq8OI6jj2j+ivDsZDS29GxSH41A2Wq1bC+FNwfRDl5KdqHxAJ6bp
4a+DK/H//wI6xqijz76T0IvCy+jicrwWpO7BPu4WRVVb6F3ACdrSy6q7+4QDuFEs
z+QWgYBMcW75/AOo6aQHejh70rI4yXKPCJQAG0OiLmy7do1yYRFEuBj8/qUJXllv
8d9tOl0VxjetShXvp7EozITv6PyIHn9ouZ59TIl1MlztreMX7GW6HKqQBqEPriW7
z0ohPynmvmK996+E/VgMtIK6KzAVSW9ImUCmOSctPbU667A15rZj19MWt3mPdGtc
ATlZD+JrkSU6qUOWycG4r6vx8pcoWl+AYZBi3d6owGZ2zBRMD56KXs42z6Dfr9tm
htwsD0fye1iMMt38UL4/m+HUWZIc2WMAz3yjfSmWk9xL9be9xsOgJi+Ieyengmxf
awcQrwcakQodQyvykNWBW79Lt4S8H4K2COgyjWWZNQvT+mgT32o9/Q8zxJKdzIBY
qAQ9yT54YbUFueGLR1CDnX+wKoCg8U+phJXwdnGDmFMC1BRoBffokLX1CnC/VRZL
nl1Re6ZVg7bw49IHHZUzCBtwD5E2ITFEJFexjBwzyf0zx/8AHljzOYS0I8cMBmxi
SX4DD6u5pwthQyPUvqEr1ADp659T9qJMQIe1FhaYE7Bg1id1j7uP+qCn3H1IpVHn
Wr6LQ3NAF4aMexUbozYKELsR8VBgZic2mU0YHH7RwCHq/KDVlqqZwmuJsntIptHF
XOgXY1XudJh1F2V8aRohQb9CDGiLzOqJUjN+ho9sa40NIOjaqAKCWPZ/tQECuwN4
nG1xCty/5xYEpJxs0CWCZJ3h6qjjFG02lSz2bGN7WHAg71zeRgXe5KYnpPvp8AhI
VXKItZVfc73+KvbO4LsxUT1B2P2AsAwJIGzT07tR6/MN/OpR7Ng8EMeDIA4Yx4tf
8M0NtxBZUiSUjShMy10OR1ytOn/Bwp/lC8Tw1XKyT2cOpH6b+QiJZY4eQSHTPaaC
hbgNmkddVXlhNR8rnXGtQOeVH55JJM5PQ86biGd3Kd4jRsH8xyEcoz/ihz/1VvFg
763iTHeoE9KhMeouYAFu2skwEHMGqxutxzBEBZQuOrIjTlbsO+xF+c60nQ9ycHU8
kvUTBC4BSC8i2OwsK/7M52XVy7y3nMsRaUedWkv6MohcTE1S2fOGH1pUSmJW5rM1
/ktv3N9KzXsP4JbdKVaICM1esfnF/AYYu32Ew9ELb6Qlble3qX2EQUyLr9GoDxJ0
rjneYWtMQhzAbmyaVrK372YrOcgd2dl2mdHbCM2Yfx31c0/4qxHMTjgFeNmExrBd
5Lh4p+6cCSUk9ZJsEAcBIv+UDAFWDCoJk6RMsR+9Kk21AxHm/MatPiL5uCHBdtgr
FbMA88cCXUl/PDFcmZaZoRkdodR5fY7gHUEbxzRiCTHA/ItwxT5SXlUMm0K+ZwZm
OvMMvH+47Z9K26mmgmEoFnyvPgoILcqzW4v4KK2FOxrDfOjjuhrYtm1y15HbIeTK
aVuc5hQuQnhIPuMisKEfT26JkG8yg+hcZci/fXnTj77d95UKaciXyOFHWRjQno8z
iwls6MZnloBzdEA05/hD1x9pv6UrT+Cjx3qfxrqqVCo93pHveKvVdckuxp8f5pzt
MkzzdxNFQb90ekuw8NE4x4JSm1nfnbDeDvSY2T6IeXPhC2YW7+IWXSJL1M6AGR4S
QxOqKnYh0yyhyKoAQlfp+CPd4ohqDBM/3gJbadTDP7EtlkMGAeAyUFVoCXdNw9Cb
q07NlUIHFSdghQZt6tpP9NTD+WR9z0uRvpp9Q27FKR078JwFDkEMq5Y839l/8FZz
TrMCp2GlCmeVnbqePWMma0pkmc9mupx5KXGb4UlpsYKGoyZ+ETbYuYuhMwfyUNbS
NtqUxbo3pzKErjR89qJBChjixltzPOEJ3tRKiJ0/MJX5cgnjzAS4WucOyaY9qvY2
Q9sYL60q6h1QYafabhQG7oCUsSczCxiLF0dURtshOB3FALEqEf3Rz14hGob21Iss
TxjfYIKim3xfwUkN+e6lGFxIsNyKojRd8+oE5dUvu925UPZxRSIqCv8PiDa6LiSB
xKBPckx5CgEqi0q1D+ygDENRkTg3yLKBT5S3Sna5ScGbp2jIzy+LSGqYamIdOlkU
MJ0j0493CRtSGosyFbMniO6iL7Jm9ZJuytm93KpjxUbCW2EJS05IFMfpA5HdmU2N
kZZUXQ9NUUqkrCyoM4H5FYMhR0xA78kyANseL6ZBS1hNg6Hk4gFzcd07gIgHEGUx
uLdPnZO4ZGu/mn/UsUm2vMtDEPG2KfOcUoFGsuQ2FrVIuJe4kKPrevm4oyXNWJle
xOiLAqSC6lmKd0cp+OVNyFnm8XKIso6+xIhgEpLkrzWwkkGI9c12Z3qvb3iqjvsh
o1wVKKMytwqP/N8tFFajZF1p6JlnvVx10QqsdtgSikZdN2p2wZHqTJMLe15JQp3t
gcvlUTJRK1yzo7yZ7YUC2aC8JtKPhDw2bWRnreqybqerhcBbV82Be4rw1phyfhj7
lLYX/Pnqd94KSXHuDz/G97bKWoXMDU25fGfRRw832YQmhape8dnezYd26rOhu/DO
Usdh4y8blTu4+Znvb43WrMj3d4Ast5xWb9H04jveX/XslTG05WidvLwnO7jncaU5
xlMS1dy2X6MrxQ7RNnCXMujxm/Uxhf59yQTHSxbJWIuVaj77NW1ltH9H7s/MvZlV
8jZ53pEJ+5AKRR9Tcqdb+DaVSALYJL/kpdWL90hkamYAkbwcpPNNhNvJATcuh4oI
6J0hrFRNn4z4Sj1Qb0fCWjj1MYwAjN9eE/9v5g91J/bgwk1bb3+Q69RxqwL26b90
IPQHZorIHfB8oS66BSg7Xc1mnZ8FsiAq+/CJmxy/7TEq78uBKjWAU2Ij3QV55cQj
uVavurVVIXpLeo4svQFOJtUj/p2gAVB9+M2JPlwf/CXmmmiG+UUNKLCfD8Bz2e+s
tJSeouyrygn9PtFP9ynSbl0UFUKtntn3PrTTD2es1UnDRkFr7UAhMTFUpjIig4Ae
dcGpvTBXl02JtAkTcdL1k76QHZH3coa3H0HhwySCrZc6laWs67rY6+BK7TuExDoL
aq+G0x3Dp+OZWtSnIJMTbTkaqqvFcHv7gVywuEqEjOEhYwxfLJJfIuKUlebQWkpI
Z1I+BIS0/fGezzBJoD1WsxlD4BOA2oWNv9/aEVOygwjVw1sV9HCakERF+Vq13wwa
ccqn0bbzcHNGtMiSc3UjIdBKBtZdZIIviJm6cVyU/0lMhavpB2NEB0F2FMFbWiV3
i0JXp0N1QXwQcKzgEsvwLPhYMXFllBFe0uMvtDa7RRwohtKjOAnhM0P66yo+1F1a
6//0Th5BwuGqzHgFP1Bbdi7QyNeaD7h8H9JoXT68kvu/Q4gveSx6aHRsHqr9A/di
s+BWPTXq3nC23wnQsOcp2SpZzpRDZxkVY0ZCeGeRTuO9H528vG2EevWtKxENYZ1T
XJ7EYRL0qRRE+UskUMkBvteBWcyoJtGw8u1AP9yrY3Bvc03H/IvTtLXK/ehXUhdr
hhxLn4Y97cRYXynL/wRUjIN2Kxv/aSYvToUWyFhMvo1SR1O6hE6eOKgkOqPzBqpb
H5by+q8uEVzpsGkv26gylarja1HfMcN3Xlx7n5kPMk8uOdFMQoBgXtBCI3TpAQSG
r3twxTOg13aZLLlIabEkeBJ/XGRGV0dZAx6fXVFW7QrSv6vSNhyKtX3ZbZKg3Cct
cP7T/sOqRAKM+GP4Od6KPvZudDqlPdnIrF2ZtMiJK5krG+1WsoSBkTxzVVFZnDkA
RBTNbpXRMQYfFNu/m500CcOzefjUQGqSVXRXMpJaxms1Mz55m8ehxWTZRimH7ccP
FJ5AsjMi497qhryGYCRfoZiKZpxih6jq08xprJ7ayEybYVaaMKKjGpOYinJpzr7r
MaSF+XWS4fzVpWEdkg2qaAsMSSAFnoyWgyJ0vAHdGXI1D38ghGH0WCyB/v/lGrvT
p9XxAvlkjDiNl58hjkYQFLkYektCAp569fZYv0ZYsfXMb/6lNhRrENzP0xViiqeb
zhHNnsYKzF/IN/Tzki77ATjLJj4IEw5kWIsYRe/ukXkkjTGk1FP1S9nKIlX8OJSJ
eocigUjBemJp0l2zTjeyXDCP3mzEUh3nwVgBS1oUNTR50T1qZep8vlLsymBEcXrY
R9MlsnPkPer/g0Tjx5ViSXJSSjsU2BLcvkkZDEIH98u6DYpnLXPvpv/BSuc/mCpI
BKVuJSbb8aYi+bz7yQKSOQDDdivqq5UVLapb3PCkpys+3+HB/j3MGxhMKEecMCDI
8ZLmVkgO6Y4y/IjZai8bQrTdkKEk8QcePuL2BJE/xv5po/pZ5elsaZ4jTHOe7CPh
KL/UCPkE6FffSmSb9duHt13OJKEXqMoPa4N+1GT0MyGB1KWXwlW9MhaxJShcpnma
4Ioio/DOMcmlnA/3GbBRlpnAR29FlzpGRbRa8+LrJW8F0UFXZxNFCAVD7iXf98VA
l/vUV/aUkhIO76UhJ4DPW4Qiyuu18CyhVFiVNTywEFUfAzEj4SkssiYGECjzCOZQ
zp29DtaQkkr79BXQ2oVY2fXR7baQo47fwao2GxvJ7CDQrKVSEzmYepv0Er5xBToD
6hechCGCARkWd4+CLOLbpJyV+kjDTboK45f8BKMStAwYzA5b+GLRxnLx8mlw9mT8
m+mIwkm+pJfxr5qrggb2JoP/hvr89gnkUj+sRd+Noplw7Pa2y5ahS49n+t410HcI
loIbPwY9rU3kOir7belBrK4oFNUVcRcyOvXC7dfEv9HTao82DOv246h2y6NCTFuV
Mg8mnvs0g/UvBSCaqbWdmL2PjSeYYsKbalTRiT51UrA3SNRO400LNcKJk4pNo6z5
68J+o3g8aqOu4Y6mbpdDEyX7cN+lhARzM4NZosuo/2XtIlIaqzg32lG6akK2ksiN
t1KA/Sr44s68mEoTV6gb5jKvcPU5QqABCQJL/t2ETO6q6o42BP56fJ3MlsLpruWF
b8wXhusZbrnBeWzt4ZvO4WMfdxejGoQ8t2YuxJF8r0Rd4qlpWBtYQO9BCrvZDdL4
WnmO3o6tiWp7yEOWnTxGY4DVzKkAqsbmMhDT/Yc0xAYt2MUBC1qhQDHyARz5/+y/
AjPPvbMcPQi+VyjIQ0+/CJ3KuZhg/ZXSddV9j+y/KaMLF0W0ZN/+fRwqfcUcXH1k
aQOZKR8ODdluI8Y9fSV9wlp8jjcTmbkGT9QEKHcZak/GumBNKMYTTusZIpdraUl/
91XN4xVn4geypbJTmssWCfFLdrv5y41C6NH/aHxggj60NjaEi24fGPB4MdcLcJb0
7inLxWmAEKS2Blea54gkZhsVpCvab5mjICL7Z29RTx2wpxeW1W6MYP9YTAx9Wbir
AWR2Eb+Qj1AtyfO+9E5pOxu+oD4DVp4okco3/0b+orgEwL1t94e/KxP7x8Qjg4+R
vl/kidH7KyLpRKQCcAN7pGs87muoauBP82+JEGfxgkZtsYF8yffnqdU99+Cw9H85
r+HhTshWbaF66XhnD8QAimOLtEonrNhGAuC5gx3JKwjLX377zrDYjlL3i1DFRp4S
iem0XgSwXVl1BiTVouJClQo0wubGLJkEvkF+Jx2rEqLEzKi5moX27GHbPiVjHcOH
6PkyTVueMQva56xA8CyrYflbd7srSFNF3Y1iB6SF9Y+Rvu+TDAU7dj2ZIBm5SSli
5rDVDWYREq5IsANfzpTZGaj8AfECtXBm0WFFQKfVnKRawg6KAx+9fpJiFn2s9ehF
C4LzC0Pgrz+Si68xF/dO3JxxKEIBIs5YytJrWi9qGrNge5nSmCZMcLsCSlFNJDJq
Xaj/gGL0Zvrv9Uq/rQ+eZiqR3SypsYwkMJwiDmTtB2KsdOBzzp/JJ38v+A+yrPvb
6XmL5zV3QQwIQghuuB9JhXZhkNAmI/ZuP0+Rs/CGXvAFdjXkujSerCPh1DVZJOEM
Hd4a++HofhQrQnWpnIUmjGaLxMKPMXkO5aHO/GO7TvQgq3dyqufPJyKqbz1VBiQt
Gon4s6DMMm1fXtfUaqbST4ih7OtqLZzAMXYH4yNIvmhhrG+bfflGL1SorLbdFVNX
KazoCvprxRFVhgs/RUC/fF5D1V9oi892J19h2FZjx/IP/h4LPVJUFYRUhhxI48Yl
nxvvgNjINogsayjgLclnf+iWAPeXCR7PPslbotDk+8ZlwdIJ2qGhi48tgbuX1HyX
zBCxOVJmtvzXzgzK/fqzPkS2VEhYiCdYrhQxDFSxwk7hn2LBzAfq2wirXClx32YE
wiojrVRgsV4+WhVhgBpQWHkxCYs9SudpSoYrlwzCOZI+NYWpkkvFRTu/jbxhYeYb
DYStt4ZZpAqUHi3XXghEc97fujikp5ZzsSdJCvpaA7N6/WJ6cnl5I3teBP08fDf7
JhuhvQ3wNZDsbHhsZ1sYV4tGCw6dP+i7fXG7sqb+SIDSBqdHErlsXRpHiYHxuIGt
DJnsVOeIuHPsGxfeW1lsds5PBqiEprdg1Yek+boA5RNeODmg7xG5yiu6MZ2faZze
hccOA4lnlOXGc2ZjVL5Z0PCU0GaL/mKURekajg8zf9eNfpDWiSCXjT64cIMTbbjg
7fogoNjfQMkhRugG4M11/Jic06rY6uKUuQlUwip/owhBqjiOTA/nB1At6x3kh9oE
8r8Hq/3E/BCEVCPDflAdAfrKkHP4NvnS2Cr2JbJcDDyzeh2zhGbq5oaCs5FuH7kQ
5YWqLlSo0JovJPcRIigsZyv2/8wWfQY6Jvb6ux85h+UZ0lZZDLg+Rf6U34V6myD5
BFma4gYmVoiv15MXlBujmzBkgVbnqIzHtMX372SGbx9OH3UnnHWzqcElHynkyobV
/KfFwISqCxW1Oz63iJ+KuzwK+fbZV7eomnHGt54hdLtz43pfHRwjdjNkfgQrxq0T
eNXleac5FNU0oxeN0ylUaNcJNBjLBnzeOxpAqIbfqh+ZH1ZiW1eL4BbJW8+gysFu
Nrgy5OhISNQZqrgj+Lnf+Z6Q+B7/Y/eorhYaQkl3qqZYQgY+f/3vmVDsiwAUi9Q1
7zCOOF/hVUASswehz2zWKaxiiWz9HVf0l6pF97xw3bFMx4iJLEGtWYp5BOERBVG8
UrD06YlNDhddAxVMLT+CYc69r2AGHbkwlvwOM6HYIWqRHiL90IMEGIF4y2zhA+zd
vwJmxRr34itXiEd3IqU9mG+s5VBuPUP50fmVnU0p6c8ZK3v3O9Hefba+3m8ZFPae
Y/6kKRT0PVKfWDvzlWUuoFOBglzodEPMDGRYdSUcm+YdiHbVLa18MhaRtjlYZgfw
e2vb+cwMY9gdm33kHPk4i+WFnoiLJeYeWL1RGrGYXybIgAv3qsOWGGu9CAAigZ2A
GvrSlLGHKcuBmCX8Y73IAN4Mvq4u3YnmClMydEftA8bSh+Dnkx+1XFqONcCWUWrK
ON5vl9bU+bkph6xoPV+gZtez3bJfUZPQZiZaxo9Iqn+IC1O+EHU56qCjxQS+tqNz
eCu/fGbtfztir1Hj2UVmbHMB/g4NmOBbY+NQ0Y53xkODW2af8hNek2ycFFgSsq4P
T37PyntbsReifSmiyikbCzwPNLKhfSWwm7zFZgylAmFU/6cOz9W8RijpgSOSDqNz
lVBuuFTL0Davb3YDjT+lWoslzYhk+2k+XQ+PtZiljAO2ERJnopGwImXzOU7v/+2Q
JrgAx75huxyjSm/77quKm1a8le/hXi4AxDDT/1u7TqA5pWT8ot0BLmUzzxGl//8E
x9qnjbIWR6q7nCPgCr7sY6AVa9GNEDq4dnMRKV2y1FzqnzzyH+EaTTRfBWMWabCp
o8vua8AXACfhKCWTNBRqL3hQPSs0xjbMpDOuuZgk0ISgZE37vD4pbPpW0xKVhjsx
qFEaAL1MDiq6WSIhsDRWM23Z4gjtS6z3rg7IikcuHhbSQ0NWPoXcILoCR0wGqsoV
Ojnh0Wev8qNkaM3zFGO8KDKHVsASUWiksnUa43P7MxgBHYvZL2vTaV4WoisfFZNY
d7m+QxHLD3jY2NlaydCpmFlBGyWVVK6nxQa/zA2Br2BV0zEcCx/Tl9M+qGxRtxFb
6JeJq1yUObxtLEx5rqErwJNLhHlEA6kcBCCmD2IoVg/av8pwDk/0exBjcQlVwXzh
Wi1fSvtkL4JWFDUlknxnzd94LyHLHjwEciYCS067mHTqBSGh76yI6KUtFO/AjGW5
uOhLZR5MLsVCfrBEWB604CZJC4q8LFy8UnTiasnxJypl2iM84+22odeb8fLMgz48
r8hqDHsxjst2eoKv4aiJgaUi2rtgzoA7/E1iSWDCKrg5xHOfFqv5h3gxRx3W7Gym
hh28CfNOVe49fdvwC8eICIX7/q+XEVXAwnimeZuke07ALzJDwpShsia90NHwuFWD
IkHlYacbxoMWpxZi1m4QzUSmyWIiGjiPQM3dZX/zZ/g5NniPaGpnsPPKGteKPzwl
asboF2IzUoTa55qDzeyB98kYYgdLoGk/9v40YN+2DAJlOAPCx7xjnZ1eJRRWJZS/
zywM35ORQOl/s2dSSiaNlLHgPqvXyLh6B9RNX6krBh5m01PBj9DamN0vxNwKQE8h
Du4PsOOnJ7diyuclwBtn/fr3EKQ3Nfi4bhTzQsZM4nuPyjVpCneEPX+hG//QEOWn
3GKGudVmUe6Bg+E6Rp016Yt5Ck5xmoOvpaJDPOk0bzi30aEycOOBPoZj4lr6347F
Knsuy2wW1BKlbU1qT5+a2wyJtV5jZ4QRrTlpuknYIFRang0NPGpK7yiq4axr+XnQ
oxYE31ATNziMRTNApea1bV48tB5ohh0n+zY00IfdAyjm1SUrk8/Ith79d9RJUjCA
Vc8aFjJ0PC8ptKIkRgBfKt9BaRkO8S3qfmirSZcuYE22/qcr/8VXMJ3O5eVD9IQy
Rr3eyW/x7JQdYH4yZIRWyfoAROeQojPcxcOnad4lxSLDWysNC3pm7mIEtRSLOe7E
MDeranr4PouOUo5yiYw5mPh0wah8q+3KAIgdSxU+IRJzngv2BYsLKPDst098iU/O
qy5Ag9Q5i17rj67dQh8Z5/gf9fLHfCz+ck9GuAK0qIGZDuS/5hSq5FgpwTLYaull
GvYPdI+Y1oPUIjnkCyoWd4kE2pL4Z/QX1Zuns/gTeLp6omSbGVtf2NaAXYXr0mip
N5nzraABUz2Sp4aC8lo0nvEO8TlzTg+QstqjgrZsrs3RuZ+2zCHRXEc0ctTe+Pxf
yNSqDFGKD4i2aa8ekJwSnCvJdXoaBwEDwoAmoPqd5ky67o6J0X+jxK0Ha/vdpNqA
1QXy5ohmVusHs916udN2BFnH3w0qdnF9kjZAuUubjUHuGMPvB6O7i8zuqHkg195l
c3f4NqxaW4nXQ15gT0w3LMWITF1gFy/gPe2ZTDRpgF1gvZQpv9w6TdUusnu8QAEc
RCE45KjswJyj1sNRBfEuwjIOqxBJECzuyjLOTjBZ/tYYf4AMtSeC1y6R+R6lW5jP
eZ1qt6Ebr5yfGJWhmsENZbKV+THgedIlZZaVdxrY9kKOyq0wpp9HNLAoB2LK1kOp
BGyOS36dLnxDTcCr9lsdujCO8B7nVrC3ddX6TpzxbLEj26nmIvtAlntA8pdzWXxJ
8at9qbvoxOTc85lv+kaMpUB3t8lGTpFVreq/uvaPP5Sl7f4CtIfXvda4y58+57eU
UVc0erhdAflZzA3sgyf71/EBq21gqK2U4e3YBOfVZskTR7TVnXHINTqlprVpZsss
d7tJGd22BcFylIk1373OeePEmJKvO05CfdaT8LAd6s7qK/qIQ1gADCbaDxvyP255
6L5w+Ig1ElacgxWjx2v5f2bYoXQ0NbZ7horkcw/ArZEzkJS8TNxhYpOUJqxcjpxw
04kS3FE7VN6vQgUDgQUts5qq1YCMC7tgoGvpZVJmrOvmqncdQ144k0VfYlNrRZAj
9Bj7AqsD0ngSffDBouaGCkEYkFS5M3NU8JrKwsAueQ+wnkC0gqZ8oJ/V+Q+/7DvV
Ta8Jvx3FW/XnPJ8FF46hdSkd3gc/GhXp2G32DhoYutYb/VMcuN7NCq/nw0XTao5k
Dczd1I9wkU+SU6GvYJZ5cbgV87fHf6WjYVHg1UpnP7d6vqZAfGpCANCCnhDRXg3K
88YeiGDhkDMO3Kh4Nq7T7NwBhe3X4h7Epje8/XkGjTFMBuzzTAIsk0SzoZm2+RSl
iNPFhdma2qte4kn5w+FkNPsaird++5+foY5ma+G8JSkrXpHqtFq7Dgnw1zEUaD18
+/GcWayAMlQoggxkmtMAx32z9YcDJ12FGlbJ5QZe5hPR6XTg1pWWriRZijs0YNlH
owL47gliH+tl5xPbDwvkL9rn9NWhUrYcsK0trBOHCb8/bj3J5VSjXcx7z+lFY/W9
uwE2qDZbL4deGKnyHP0TXP5hmu0hbeu59VL5U3/p9+KvJgGHEWG/FfTPtBqqR1rY
S7mZjPEWsLTLfMPdWwhaD0FlduDx0/e4k5uLXVQ6SVyDzVz8r1HvPllQy1RDik4K
PUoYzt959jb+3uYmfsYDXSxRiuBKqTIyQ52M/yf8SLcdHbCfL7c5csQwo234xW1i
I9l1wU50lqsjEY5BJvaobRAiH85KnSAzvrF26Q8Xob3I237hScS2f6X0Ygs6prMM
zpSGCORMKHsAuTiZ9N2SZ3kKbuL4FNEI1fN14eo6SGiOdQcrAYHOkvVFvS5TPV73
F3UQRbf7vnLKrZk2bxFXdK+QiBo0w6e0RJj4PNJv8CTcU4Dv8ZvQRTMFHyJDkIT1
LpATA2b4EJPeiSiOwX9S6TnVNQdVmIchhUe14Yc9TAhUmwa+pPWDMMw/Y67hphdY
BFK+jc9mHSoeHVoaaASoyUvd4iJf3z8nQtvfTHRx0PRO/Kug4S0lQ5lxqjWSLEZb
r7eTMOV5ntgq/DAj2CVt1TcvuC2CfQjULIMTPzTufl3tsusAwz2SOX9Mj3Nulys+
5G0m2Ag8vh6g8YLNRqZVnmEHmyPeweT8yQ+zk34hSf0Lb4SU+cipBBZsHMgb+DG4
erz+AqfSezp8M/S8w347WwnuQUnl5KlX12U4w9C/wIPoz8viFMiIvctlAWRMbeju
69at7lXIo2fhuapSzFvpDT7oHQDz0+9YTSIO39boGrA5qww+DU6Wdwp5yb0mxZbQ
SpCnD+wbaQfPwHzyb8pr8zyJLhqGUhG6TrCZwx5qqjQEA2FygdOsCrEnmlI7EtUz
eDbR9QIYmXiEH35bvQlVR55jZQImTLqtnF7GaBc1WdEn+Ue6QoqjoVHPhgGR1RJF
QsvZX/yRnBNC1AksMJFDY2CRLMjVde+0jJaysiLjAZjbJgq3KQHERxPp4ysd+WIc
jUdWNnRnQslQX62zULFO8cXjLmAJpyzOeo7PyytvOuPnjtdrdeA8oPr0MSUqe7G8
sLwmK9B5oQr2VEN8SKP9/hsznnOaaL78zesOYpM3+yDlhDa6lwEWYfbLkXSCKqfU
mjo/Vp+IuSBMebJtuLRg1jPBdQaeR33388eiHkstAX5hcdgSX864UHbTR2IqczNZ
tkWoBHVlVK9A5+pp3N6kjRU5QHirhUX2SUFdSAkMXw8ggVVVr63G3ORfkcr4L4s/
mCV1HJM/kc5ocRAPRa3BPvzTP7Fs/TrwuavAR6GtVC97plihTFlBmBq9e4bTl0iH
YcS20Ie2DTOaTnYIj8e1z0W5HHA9w+0RxGEWUEvFauJBRJtS1IN8BzV0OKAfST0u
RN7ChHoXnjTo60V5ktRYnepl3kTcq7Mpjtc1baDDs8tEkAq+L4rE2mRpcVcJ99LM
SSqTF5HGfwZnzmdDWngV4xaX3ECMdsuOFmdY+6ibc4zU0ZNwH7pRHh1JbLh/OyLa
pMglczR+gSTjuP8HPcPOW0g6dUz1UNrswsdc9YcE25r3B38rOHqvF3pDuZ1zoGag
td7ManNg551jaIe3Q7mfukBljlzb6Gkn0VAak19bvtNAv5rpG6NmoMzp13XIsOuV
TkHjYuKYXj6j+DO3FFoWZbi/1a+TKZzjps6qkeh9/47iKTmcDnZh2OHOV6A1HdSx
jCIFwr/fB6KO4vDV0NmluyuPbQMgkxDhIrq0nIW3a3y/yzATChU9piKcHiByAlku
TKFXry5aPJXYPpRyHGAN7l2FXtbnpw4yEGh2SlzyLawCQE9bepyPRWV+tnYSU2cy
jFny92Q6aBF340B+fU1MN4SsN9xkvvT4p5laVFoWsQBDsTv1gxTxJ+ooSpgJ/47N
whkMLENnUNnL7Z6uyShGOtfEMZVZYRSJPWJijjDXRPxeasJByhP7ApY0UJ+g8v5A
zZ6Hf20TsEhp4Iq4LM+RwojN36fZt6v1C/SMBzGreeIlnGv+8xI9KyZFgnIvSUz+
YlpZU/pAEw8M8h2lhm3XYMSqIhJIAtMEwabiCYfbhbYqU5llGGtywkT5jRHzni8a
7vMJ0VKD7FT5J/kXMF7zRocl4DV1SHK47N9sfLtmdLQydxQrKOB4I7GaXYELJlG6
oFC4XmlMB1FBE0onEdkM4XtcFUwl3kfOv5U/7kZwB+weCWxKXgZpKzqv2TLeMubM
FN2uEu7Yr2jgLo8TJTB6AlV9Wonti82Py06tn2T6IISMEviIgzb4r11pU9/EYmDm
L6Tf8DzLPPZPjYBZoCwFc1RS3AjVSAPN2Hl8EL265ByT7Rq+TTJNX9aW1pXDOzjc
MluYMbqgO6lhUHMfHljvUaCxLy00c8xMKB2Iqi7asUw90LDGCnGzM9ZWqtatT4jx
z7yXU/W5k8zmcOHuNmv86Ssm+EdGLENnm7YWyNnzPrr3pNCL6cBxio4Y5LrIYB4S
JmJIJ12hl4AWkaxrcnScZFEE88t63Y7lIwb2cvoEBruImG8Jf44q/Vrcr4P/tsfT
DNRnos1ThABkSLqsAIwgY6FCFsbO2cLSndY5Ew7Ncu8UBPmvjmgcGD7NaB3AJrqv
r1MPnhofhkVY7od1QhS7NMlNBINW4wetJuMHrqUxf16KJBcXETWxDOdYaWOrVEoe
LegW8P1lzAN6yYqkfxjINKg98eeBYimnSANz6B1vVQZkzxpCzDgjrNL3K89NkfzW
M/JWSgnoESJckurdbv8h+BjV1SKliHNKYW6/3jnfwe7Js31rgpS6MP75+Eqs6W+c
nxy/9Ko+F51aDSNVEYgROit4HY55Rov50A3YHUX5wNN9Hl/8+IUheODMPozFozjD
7Jx4lEntAit2ejK2h5xdxvPbgzode6gpMgbdvZVNnEddlzkQoEpBXhG/VMyXhiNa
grrEW8BDmUz4TvHCVeY8Gqt0XQ+BwV4kAdTuf0a9h4dBs+4rGDtte0nA7OHagL6+
DuxCjtg9FNkCLY0Ef1fFrjnhsxWywANDbFHES2ZePK0CrUNj05nVR/pgOijWC3WJ
vl2/Mf49FaHafKheJhme9CVbRCsmQqMlDyZ9+wsmjucVlxZsX5He8v12lRnyIi/z
ii5a3z34BLFjIjqQoULk5Y+RjBiNHfRljDrHIdtS9rIRutv1VbsmTcjX/kzS74LC
qJ0MLfcJ6wzz1sBTVBDy0YVZyJoWA2sHUyfHa7Q09IUCgHUbGSuLpiNrMHudzVRq
xRRau/PZtHYMPBc199lQeexsMqTO4W0cM/W6cgjFfXseSJcC8Px7rESI6yfIzu6z
Nmsx/TZvtvGClVDvN1kNfqzUn8ZiprBvcyZFmvy7Df3jy48AVmYD/ZA1ppL4GYjt
si/3n2uLxTvjgsnVxxSQWVxOe2IVui0YMpQ5D7ECB/ZBOyAGTHzAJXdkz9daMv66
MwJIAl3UtENhb0oiv9xVK6sou/r/vxBARuc3zHMvng6LK5yIyte8O5j7tNa4V6gu
bkP/E2oQuMy0cpPp9rWlWdq4A+vn8DiVZT8J2kMdYkM7T3T1pXYN8R/bLtcaJ/Jh
uSSjDz8n2G2ViozufD4QqqXNj3YXzlRdG0y3kT021Ktq7lRsu52ImzIiwN6QUHQB
yG/r2ar9UF57bEhoWHpD2wuNoMfb583XRFeaHQ4z7qTSW7xc2nFpQLuOX99gov/l
hy1V/Bgl1BuqrhedKfL6KapzwjN/PBd8Vox1amI31S4KLeAqax9hzgb1xT3YrhES
LhLZ95PaoTxBL1cLMQdQtqIVwMeKKvpRWI0U1HRB3sASXJiZB6Js9F1v+r5xkt0G
zXjLDMcBzwFaYVceb+jTLyM0UaBumhYRxJ4hFfH7peGSfomuWeMYSWSQO5SQWDma
hhGskHkbhzxo0WyJZ3ac3Eq6kvXJzovesphTlGk7wrh/TMICzIckz/pywFlUdigb
yK6VTxr0fZqCNdnbtLTR8ARwuNVOdyfbFoR20eSBdvQqbh/zl7uopzL2DmQ1cbsh
AfU1cs5MWzWoNtq4MUDNJvc7iD5dSEvta2e6QAB244LUjOPdKafQSCh/BDSoUwWJ
AAby9H7dDisxIXAe2kkou3z0inygkKsvp/mrXvlFnvSb7sVrMF14QRZYgMx11pU5
GxdY5WAof+2LYaCmI2Yqgf19rMcE+Gjl3HJgADVMilndAUWYr1cDQx6pN8nLDH9G
bjKzKIGEHfBkO6IdpwW1oK4TVIPngW7TL+RbVKCAJS707ycGe3tny218L7cEQj+t
ALjaEG6siBGfITh9hCBJCr3QgrkP3xDivIW0JBpltHGWS/uQ/r8+WxtHeRu1+5km
oeOqR/VeBYYlaP9RncE0NMxyVoZMSFaazYvYM1Sv/TwLpnxpbKfjto4jgfG9vDjb
kwAVUMENQLV8ZpIUmM6hFGSW34LcD9ts1zt0mRgaqBsppNNYHEwCX7UbijPafcBt
Y5DM+6p2l4pc573UqAEOybzAwGOA4/8c7fR6mAEuNheFfyQrnwcsN0v5YeTQ+YuB
/Lz57kU+VwOwyjUFyWGLMsg+WI1y/vVqU5olbGRfGltWY4Zl5gerld02op4dR/Ut
HOM1kqce+3covS4sYFpcxmGbCYjKLC7q28z+kOJW0Nd4zaaC3Vnse+/HHy+P3xqn
Hfz0yAJdNKPZDXGJl9ROKr8YpTc7ZvBQ1SZtgrFFRTj7/fxUF7ahWxLaYETwGxWi
nzWeDKpbZX0plskpPNfMSVA+AB2siORrwC3iYFQKZ0VcZmE/YuYBY61fSus4s+C1
t5m4sPAGx4bigv9hm79iCsjzn8JJsKzWeauTKwY/mrYG4QvOAGTm5yU8oBt+zBQk
Gxcl4CCWB/LSKUNlee66ioaS3GYhmEWJt3voOriiPXM7ZrYw81fYzBuOkj9m6PcL
jJ/Gl0390kCPW+wF5atPtZhdffLWDOia7vyicSHpaJ5SK2RvtPSfDT2lDqMM6iKH
Ya3ez4InhUu1cJzb8JsDCFmfg4L5nDNvwaHupSIc30MLWbuyLcjg3Xonq2wySg0X
M6LtAXV7lzdVz7xiK/ycKU227RS87jpF3kg31RsyCmAABouGjmQqGGeeG4ExbJ9h
X6k6+0gxIUefBukDPNhjLZ8lu/Ka3zwaXj+HWBqonvQbAJsQ8tF2Lmy1JMuVx+HR
FteSs98s6ueiHG1M+9GVBBDmH91NsB7a5v7GvmGYldr4XvMheo9p65FMf4oseUW5
DnB0FhfR+OAYXoomoTawtHMYbk5WM3sm/+Ej9wUlmzPk9sOKxTuaDWR1g0fqlnhI
HGClctj2NVNbfZ47c9zG6ap7vkirkLiocwhiGh+DE/jJMNd+jtRV1nBgvTpp5e4w
PaNlNmgWykvJEF8FkrOPgezEeo06sUWJHhwdzkii7d5yrQBYuDvgIS/hlFfHn0tZ
rXqYcRgaau2ENNV+Q9T3GHO7HQBAsgzG+wcWLYlAJc8S3mpCnQzNOWVZCEzMZBo2
mO17tMYXJ0o6M6sugkJdIWLIiGK4jEk+LSRwPgWXuP8d/h860W5zsvYXlr73z96P
zMppUVNGR1/rfiCNbKzSbR8Tlsy1D5NurGzOwzEEzb0gmrGUMBaPXiaZzgiM/aof
6BvRISqKw5y/ye06VgnyfMLxxBuCq7p3vhaPIMU4WPct+TQja56aT8wI0ceZMO/z
ORtyebpgkmGZ8v4iE1CxMleZSUnZZbRpQz25+iObp59qe9z5NCRRk8rHRBn8FjF0
G2gp5y+6UptB8jnlARPiy23C3TWWP6S/u8LGVmjU4XZltGtMIkzKKoh6KFMHwVYR
yGDeVc9omNgSQv40JvFirfNkcRLgORwmFju5VsSk7dMIcXRttsxcSlxZIuG5SG1A
sU4RVUL8cnTWzlpS6+UlFtj4k9XI+8+qWgdOiREC/g/i4yjh5CRNmzY7BYCYPjv+
kqTjJyt7R8sqbTq+qUfHO43EbO0NAmQKBQm+/m7A8mRE18OfdOHC8S4K+d/LJfJT
9jTwlH5NlylQdA7BXEWlKFZ6bCA2sQqy2Dhr2+miOvOdsv6WUYrxOvRvEQmkMqpT
v4G8jTkAJitgKXkdVF7lMRXz+nuK558xT6InjddcCijxWMYYBhkIT3zYb/5H6xbX
ATa46BZAbYxHZ64bp6Zrw/ZOKBXpMMSqiHIT872eDLQfc4f/JfZ3LyD0Vw82FcWW
jmcCBRhU+NeDpa9TjOOhlnk0ZyCxLevDxTq5aB/pqQi/TAZuXajrlJAR4iA8V10U
Ypqd8oyNtYbK9Ta3Jb4Z2eKBXecOiLT0PsSQdYRU1+G8f4/L/oeC7ZkThbgZWSLX
GZVw4Q7drstA6Q68U+BmwP94n9XTjeJ0TVCLyILG4tJfXu1Bz3SvWVqpudwC0+vh
wpvo2CqlKhnNvYwJRyLCzt3gLAgzZHvudSpz8QYpc4/Qr0eePgGPkbSN1JHWqG4z
FokWzAQzAmdiy5XlMfObfcD7NIdEBGzh+uyKbmTaQri6C5je9DpCELBPIwxuSWyn
iNq0H38A7lx8OmN+cPHFgtM09XBpB1G6BsJa4IYdB90T815FwOqtFe3pPGewJ20k
N9fyHBwir3f0B0+tXzOXsdgaVDZvvBAqFSiuFb2nokKSFGCKD/WTTQb1//VSipEh
tIeQwkHF5lWdCoA5CB3qRz1kytYCK89udtcO5sF8JRFpELaG1H3eTw+AZvTESELv
2lab4UY6cGDTSNUgkJwPZ3PYUhcTbLi4k4I8CJCoxLHeeWvVtPkW9wcbjn+oWiX2
YNMkzjSIYx0uLjHaoMTb2C4sgePAXr4SNa75I1HL+2PVxHj50GEC92J9Pf5OPpRR
uNoGzmt7Yc+kDM7zKLF3NXcwZ3Kg+ZyOUAnRP/V3JTy5BVlezYDEGDnC7WxgkpSi
xwCPjNX9DO+VpTSu+/igLdgtIRLBhsEGjYm8dkWsW5mknpf9PcGbPvwC181Eas4Y
SuiD0oWF/J2oga3RI/wgQe5TiG3iBsig7wEKfDa6U7u5I8otXUGxoWXdYYkTZ9sm
6gjSKelJ0/zGlhkpLtuuqIg7Oe58a4xRmQJ5MIiFiLaF2EsWelaCbUtydX8aT4d+
NtIhYd6LEf+uxrflFHG7VyflKsKdDlPX4UNok0u30r1+r59RNJzF7zqCxBrwbSqi
g1ouc9HRaPJZbPerfrjTVU9DamqGmS164RFl++PgTl4vVCN+aShlsiqBzs86S+Re
TqG5dorZXTQ8lsMPavCS9yN23lpeL5GTPwqRNBt4YvcTZrgNkEswAM+lTFe7p3kq
6eTTNvdZf5ED9Y+PNu346Rvj72A89/2pHhNRD2OuaLMyU4uMDcvkX4W9bo3wV7AG
Ge5MATEGb4FsR0J5G/5TeFCW3EsUbVLU7gdkxN3xafwk6TamA7kHtz/UuneJipct
npHIop8AyhcdZ1Ru2cLc3LOmXqzXGKkV7X0qbQ+I0q/lX9Kw+zmdf2GlOBlOsM2k
DEdWrNCeJGY/wd+OcflkH50FHyRcSUIzOsEBwKmlUG+Wqizqa2aYLl66q4dE/WpX
vwdM7GibiGDtZ1HIUfDDVTWJ4QK8WHSCeBtxPJLhAD1iwiA5luOmyQSf9wj/xpgl
FVP1W6qFI7EMZXNM82mBMvhY+/X4cUOEz19XNoi4I9xvEH7mnchntEM49yOtRI43
7w9CbFDuGZF+ijcfu2utCsjPoQy9/+7Y92aKSQllDp9UJs/kZLLeY0PPOjTolESK
lp5tIxq59IKATpROMSWpsGtWMv7VXvjdoj5F6rvYBq6wVbgJQQJ5nVgaFp+7x0Rq
SRIw/INt+X/V7GHt9oIa2AAh8xlZ5ggwVFWJ2VkKQese/qzQ71BF6c/zhi3H5IoE
8H9ADYF64zpech8TrdsCLvXb0m23TMrMZzIdZBjfSFfNULndjyS87qJVh4HOcpz4
gbvv4nNklfKUhXyh3enAiji9pbDz3WFPpMLmhd49wXvP8YeeDMz7B7Vs/QEYy1SH
b2aiXiS5xVasPZpvLY5GR2N1nm2ckhwrl25gXo+BjABh8H6a8Kzigz4ZfMQ7HrBl
QoRZmFEtHTjM8xN5E2vP4QnTqSnd4AgcTRl33LPjtC+5gVZsyHSbMKp5fvfIggc5
H2CRg2NJkrHJwMWnVjTBR2pYPvAWUUvrP6no+2dDYZt5I4ia6Kbl8S4HBjMUiyvw
njrSjU84HQZjZy8Xl59Gqw9vo9PcUCkO6dNq6vnrvJoXvA+0G6MbZ/fIV8QgeLum
7WgU8sfIlFaOw/vRfIjnv68lSFVxs1DLAFDApYs23ompHsHi2MEXz8JfRAfG8fTe
hUZJcK79TFkPbL7/yR+RLIMJeXqpT9KO36mqIV2cek9PbJqebFJy9FmEgpXs6y+t
b8lLLvg1W2mRrtTEAVkcaeQ73V+0yHGNUy/+U2DLYzQZZ2Mj9gLgnJBeMeLv5PWL
yZ0LsqRdZmLMW9gGLcOU00rM2eBnVVJokVbAP+u0baw4tU7UFUs+0d/6ceabld9S
tgknYeKJVdSJUeTLHf9JZYAbSgAzFnIqg8LHP+cIoGWeUiQJH/8cxgeSKW7/pMIZ
TIO47BP1MM4OteJZB61dg1QiO/DxkBq1JabIFXb6YeCvvUY+McW779NEAxap18RN
cRFJMplmXUm2v8BU9ApCuGzAZ5HhQLqcfjiLJWPDGJZyhHoqf/V2oIEHoCWidV6g
sHlbOCsWgqfcDKMbj47Vxyemldqt62BQoPYP67NgJYpRbK08DFQosEU1RuIc2wC0
SHKvM7qug6gxfA1uiJNCTpFug/nchHgDcSvATz4hSw4kczt7PnYyBTXzJ0KilCmG
crKpnYl4ehFqafd6QdkZKZXJP2oSHjYFl+pJitrb/zQnRm/omyfy2szGOqci90vK
zPeRUG7KwGoRjTZtA6hZLp/QSsSbVNIh01bkSA9YaqAPvXmTiUQMljl5qbWwSN9Q
/tGD0NufWju1Cllz4vnY6aXbRDmkWxpelWgdj9zS00LGOFUyAhd6tKF098q9/Glp
dqrdYAFW1QB4PMWXBiIS4M4qXbEKzS/tnF/Y7Hqnxz1e8skmiv1/3khc0ZcT4IQa
bbdsVaJUKjnc2W7VuUdK12A4lveOoW1vjdf6n4hZMQKCDaYm/a6u+y8w445s2lVe
DWbo/xkQTiKR0QUPbu+rADo6WQDlgKbMCBF1k70sTDlRJVdt6d8ByJcml0BXSlHH
hBTdRc9ZHNrhfUfccLmuEL4IxdbcXrOii8QN7nyN749WQCV4F2O+k5Fihe8FLEdm
qD7gG5SXtf1LfgyGkwVdc4gRSGxmNT4snxIbQ1gseyPtaZE0AVQONvKTqpZEPKfd
7akSzoLNF2HixGM5sQOX+BgrMLVyKl9h3iTzg/gPtcUYwp0fRJEu5/6JKQTuyIYl
igQ5rIJoP7VTybPyvavsVgNBQ1L3SnrT/cRJKHYaS5hs6QaBsE8osD49jIWGy6Ho
tyUs+WgHU1KSr5yTcBkqFI6Y8izVAVMraA72pkuvCpLGON/YT062Zb0BnFP6NPvH
aEmRB/VpHmXrqThLgvxtrHee5Herv1IrYO/zDdP2VxOPfSx6FPjF1sc4YL5jx01R
srBNP03VaXUBYNceuoaFMrEgTVAbpFaGmUUJRNhIeU0sXOPxi+ndCkmrpNfZKSXs
aSPTECud4WrVGfprrvSm0W1eHO/Ge4a0ZCNilfI47UA4/r5SyXnnF9O0qUxXGCqD
bE0YKw/VyNU31dc8Md/oeGobBkkmEH9KGzUONnX3d+7rwbLPqjzjcouSd5z4UbQp
1yKKrAc+ZDaDU5YW/urPz2CUqb0HxGLGc8V4F0nKOpBaJQ/F/USrozNSJPIsoCs5
/vz3XU5r/8rA/Oszc6NS22nSdnnpkuGpTLKg9SDXsUbYnMHD+y4bWK4BHWXnJzc2
EtIKwV0toVrrZivZONb/QvEKwOf03s2fy9l8CJNfd3dgoVDNG1lNuSXjG07E7Ccs
pmnzIrXLv0/a5OwaQEWmaFaPmVAr5kuzRCO+Y85eG6hefMSR5GPYRW/t6zI1LOh8
kcolZI0xhP+J32lYR39SgUWfsnNX1qaIpntVtleN+29DacrfIn8pwJk35uIdsciL
cE2Y7r1qPD60qQ1j0DnEzEmbGWQepcnjNeWTgkFwKUpqBwZrZFqTU6ukTTKC0bb/
5NEgrFab3jFk2l+4hvAlzW0VJ4U2JDfdy6pRud4P/hZGUFSIFV1OgwRFUOpGU0ax
6bjpLihzDuFwyFCm+LQ6h58c8xkTjRMsLnke86qK/8JoYorcn5hodzhQUC0seI5Z
cWHcw+kP5aunn+lFMsMerxSXDzsXWw+KTJG6FmeSqbey0tbOvNOQWpiIu5HmAliY
OMHShF2ramzTKI0SwLKKH0WuFHYuEGO7GqmjhOPwg9iTIySWEcDQQtFxxA1XFkuC
3wLT1D7pXWNOauljiWfLrxhmQSQjfHoTBjw+KSLGiRbL9loUDzREZnKRuPhs8O39
uNe1WoVUYDv5NqjxtJVikHby65OGMLlqtux+0hJsLdmhJrQqnMK8xJmk8S/hkrxF
SxmXoibbj268ZxflXhdNjmyDUSnmAQ0w+7kuuw0GmyK5Gdkjo/1qG8lXv8GXVvIY
kBq1TxitXf1Gdx7jFVd2CGozf0pJI6/8rUNunVfRS4Ak7xL8Y0gIzPCeSoJACzb/
PG0Zn0f77MCdzx/Z+Q4gc3IIyXHMlyG7TC6rCks0SctxqESryEdqkef3+RBjZqPr
MBwMklcolxlxg33tWDCdh8QZLJ56dj0REpzfss53hgDqoDonhJpA9wLFrGO8m07s
532uxdFXT0/Z0OTAgTymvDQe0v+8iI1LXP34QcGJPp3+q7K2JAbUGI4ZN0QBneWC
8Lb/MnuECNAzSq0D6++tcoFJJ54PFVvv2UHTdscU6eEKgBADACjLkEtHPabBdFMY
AHqGn73lS32G8C8/gTItryIoo9RPz3tVsJvVsAfdx6237F979k4+EmOzf4Q2i0Dz
pkjJ243OJJ95FBkublyo7m7Pk3k/DaJ/7CmhFUBYdFBRmY12Q17d0V+QUiXcyfTn
DbuNL05MDEPf4uJaCSMkRwczEwGvy8Vgxegblt0ORQHXrmHLISd5WGgOzQHNYpeK
h9Io9nVyPblBXin9el1ecxzJceFhY8rEg+jJMdhsUTGttV82sqm24psjHht5Tctv
FMKW96SEQNrjSFA7SKCae9Ri1mVmo8u4CHlMyLO+290/M4EPlCifJqtWuCFXqw+1
2/b3F4L+eVWHIclQkpKx53wRZDP5aJkg1gSxOkabb43x3GAG5oQsPcj2sD/NRvC/
iRGPyZNk52cbPbipv0/fgOCxjYtCpXk21QN/WO8t00lJwjcImMldB7d3xro4ejL/
+Ouvqd6bgjYvuH/EUVscjjr01aeXk12jMgahWnSXCg0jUBB35RasLVS2dixfjiqw
6vsBf7CmCuAK/oG9oGm050e1utjna2MAhbg31AevypJdGzrRdGVvFv8lxT5F9iOu
Qx0DDPjulRrczBVUhEzKNGoIxeIoGYYP12RsELJmc/l43kuRPhqDaiVOAeM+O6tq
0HVRFbafGSIqVgajGgy3bxXnuvlytEjo+U20wlS/upuI/+g2Ir+6z9sGl3VmQLM7
XwUqdiR25IDE4PjW2iqw4ZYPWJr30apd/xplIRzhJce62WwkFr1H1ZmyvgSX5tA0
ae1sFCkF124avaFzDGzG/UG1mixrdgIZFGGOlL8DpspKT/Yqjz1uQjWl0whtzAao
b4YSV6+UWG0qHh6iBIF1GWgLqqdYzzxhKSKWRFzZrj40jpMPXrTqV2KZCSrGuRFj
1yisVkyGpr2mo3Ynn0blD/WczVi+IkhiUUBprrkvPsTbMicabCk0dWWfFybwKIKk
0yypPbLMgGyqWmqyixl2RMz9B7azuQ/1RqFTLHK3nxztWJshSZ8IS4/QsOjigFbd
Yv+kwwVzFZDZzIF+e920Jn89gGu3dpKu8DfdmlPzDDfuer/eGuIGfGaQhTlkjekJ
fqbT5hF8IxskRu8ekRnd1glU+nF9zW9yIwdLnN7X1gnisS0M+Ctf6bL/4BtQxmF3
J477iTG7g6+iF9Mwmg773k1q6uBB41cpw6QqgR47ZDT5ZMISmiGbgwczecN/iHi7
OneIVW3QWVDDdOVVkPZ6JrHL7rKcB2C/k1fzAnQAHQ6VGYLb2Z9AAbQtB+7jPHyF
HqymAWPkjo0DQV6L31Zb8h9my9teoKEjp15wM+jnK7i7gqoW0k+tGQ98JDfgttyv
qBbVkLQ21RlevxuDdqpFpRApdIJy8AP/TaNQuCuTySPVSefPG0sN0hjapgwUxpgA
YKtf58ADb3SqEIQkNAp/w8lOHJXNS1p8t1aBaW/In7U2fFpSLII+HRkFPudk29G3
MlTv/Z1G9Nob8GSY8HNoGNuCThBcmWmm2QyebKjQn2Xx4CtmOYT30MAHeREw6uhR
1DOZn78zHLqrTW/8o4BKJMzIHtN/EQ1tli5Z2/gTWhcooxsCjf4RXQT10r4Yp/wm
uJk1qBHGxxcwOtA8hOjWWoAnPatgzbrJqKsTWntIfvsFrw6CV1KM5vphtmaJl1bx
eFF8y/jOglJlG6Faqy6/FSPGHlW8bFVEOOiGZW5jpo4hd3UxF5+RWymrEufNWakG
4KdQuG9nzD2iAehCBqhGpUOMQu74AhzAg8n3zvoiqQi2ASHqCB4nb1lcA2UB9lOp
ofnZuS+EGoLAveM4EhqF3I4UD7fG6OHcn9RPDOQL8SgsVWBvd16b6xQ3VTw6uOj3
HKhUPtUQk3SuT00ZObmBLUlcTO8RuKtuaiFwkHqG8RhOGIpU2qlq2dOfN9+8/iqt
JY4cXZ1tcqssu9rFIQfx2gyrMGGVn9LDRU2vKA0w+IxjjgtJ8dBBnAK8842dunF0
254oe6A0kg04Tj/9BGvkP/Y1GgWg0knI2uy0pG9t6FimvzR4Y9gfHWHgRs+R8SPL
FDHALGJbkpg1dDCiqrs4dSr1AcpUcWHqBGCIFaLuKc6F8o/fFVFxwqIQskFd4pjD
CBKBkPNAU34kdTX39JuYlmCCdOcRUz0wEwBuACGLVv1wd2mG3W0oJWe0/hdtchHl
yGQb3LdCcd5nLRBAKbTKo1LfKJxIUSDOxTKByQjT953UdtYTvRMHCpEi6sxdAzM7
S2DKtbcFHSS70LzthHDSSdKV8KOwreWEkMyO7c/1Cxt6RGY8IJV1z3HftVyZ58w6
k2UyhkPa/tKcVItfoK8ntCfmjg/+JfA/MLUSS/GQCws6TfT/tkF+62TdgL8a+5oA
V/0cXuD9q9S+sZFqnNU2XazEwDw0Lt6V6VJdV6GiRHXaaMmPrIXDlEjWXgK9T6fH
JZcG1C9N45qpoeI1Yq3JAkD6bgn2gKnOv28kTPGXF78X3/xkotfAnGzg0vNslqHY
x/E9euS0eOaECtDUBfI8kr7on8DQ0GvQ3M8sC8/LwYTf0CqEm0ziwLdtkqWWlGwz
ICTEaQvjj9T3BrFMqRslywOHOtZzFemflXhbq2tEmU2xWuy0vPrGT54JXGF7s7nh
98ArJvVngrdZ/NWqbqQyTepkAWPbVBDjcNKAesf/yKnZ6CL3NzxR4weFWaETmv2G
2U+WFPzHufquTsNu3mVmu7VnVgIutWCkHqmBYtHz2RIHAVLUDSB2KSJ5VHNg8LKN
Uyw1j+/46gekKZ12O9IMY7I8dwCLMfXG4rOu1MzPGc70i1Htuz+YGeDWWZEm2m4U
uHFBOq/xzeLKIZim9K99TGXl2S5lCRVNgknb6qGfjEIzqd+5Bj8eSa3wCobjDfph
EOOnbHGFiJyAqDjydw4dRdOwC7eNqdHr8SiUvELAt67WvqT81keotsHpkQVyrBdw
3yQfxMqR3h7H/48x43JhzEysV4pZT6ECHTw2JTpNS1g4G68hHXiyc7DeLG8HKRJQ
++3MuxbLVizJUPt6xidwUrVw0wI3UogQ0j3QGKCwtvSnKew/Eo6vF8uW9v5Huony
Q4xZ+AmG7YM+dvMAhv0fFhWwqyKEMFGZxl4jGZuPyb63mrB+Wrf5YOg/360ePmtg
Bh4IUvdUMZDBSbScuxmVDMFcSHU7E9VIAj+a/qOqvQmA7N8980opt4+qUjdCx4gm
KRZgIJ17h7z6r90bwnAn4g6voeQMUf1YczBaIGX+8bwwVJHkUGX+eO5w+Uc80D0Z
E+fqceDpLiYJoeJNAN9c06n45r5ves1Xz3i3asiHYwcK4uSaAVUpZiReVr0kk2Tf
CAyOFQMmXV6gcDupMIfCc0rQZBsy5F7imPEFj79OBueVHwTcACcYcmhXmHgEZ3kP
HwmVvLTqODirO5jsmvs5/AYnLfbdIwa0QUxP/9kvxwC83RblKOxjQR9baJM7Eshm
ZANbnVmhKP5oADsJhdZiFjTjmO2+5NcpW1QQQCK8ez9eDzcgvtiA0kwAPDTjVtY4
k164rstcRm9+w4g+OuG9m2bllmHqeuZuH4ie6M8A/aRLYnSDN6yTnsSA6Iwf89yg
AxIo0cFQhdqs7tp008Oas0OS+bdKrABBb1tiq2cX7Y3e8FY3cm8hKaodRkDZHAMa
FLmnFJGPcWBvVqY8d3eaC5KIR6ke1a/UboALsHM9OVKdJ6Gu4RGwjrDxHPzm8d4C
P41e7/C9DNNVQgVl6/4rgzQMtPy2TWGje4YeLplfvm7RVSmSsywXlyfhUilWf377
Xyv+LGnusGk5gv3OhzHgUONH4uTGCVOw0KMszRPH7ode/mPC1AaIGUiy4VwnD+WD
YV6AOQ4c85ckj8AljWUGekPrnCKHWxSz0in80+2rAmAfYNquUmE6c83Ey2xdsOZH
pd35M0cLptR19jld7OK0P6UkbpkAp9XUGf4b6pBKgQS+vZkK5eG8sq0xQK06M2JZ
XJ1Wn3L5tkwEFaxU6GfOd4k6XAU8c0CQBTY20C/I2MaZ7XA3fdh4cV+ClcvTxa52
dj4idlTVJOfDbdzqSAmiVyPYKW9JroIsQRfvQ2KHJXY0xsXyyWaVdV4ms2BpC7Ko
bF2zm4jJe6yP7Fwf5oCzbbKabeyCHQbn6+2BE5teSRnNHiwKpAiM0SN/ksQNoi8p
TUXPID4/uwlCbHGXpfioo51tPflsG/M6bQkZcu5+rlanzIHDGV85Gh3OP/sXEvtU
bRlcsLpFY0FZ4ttDm8PTVskPnzIhdWw+Q3yYvSb8gjeYtAplgpmWAXptoTnn6LN7
8ZWUZmCYJhPWFWdRaCMgSy3yZhZL/t8HfsLHx+OxhsWLlIwIBkti3OWh1kCe+Eh0
q/N0c02NlFvGAVOgyLIAC9d2c6DswhzJf5QFQRuh10+skiB3BFLvzSdFYsz2us3Q
Rf8Vuzk98do8cHKu8nxCfahqcUU5cooIl929SdF62Y7/q6dcxjwWogzS3Qqod7MH
Lh/pXryzU8cPm8AIgBYw4bsAimOsZvvb/0XnhWawqR6iE11+hSh7BYydNFJAl8nW
tRNXRS7hBZRzb4YCCUGIwyKPL3l7aswHAdBLSvm4tTee8BTSV8Yk52QQP2aFaYI4
DP5sdlc7YAriiz0roAGaCflDxViFQZZLslkiH6/wrlmyNS2VqOAEieTNYHQRO3fy
WCE/aHuu0N9xoIQRX835hCVVtqaTJZErEXxpOoO+uTZt4dETqxrsK5m+ymmr9IQh
TpOyayq8gpe+xbh54il4ECA3w7rtFjzoXo6eez/H2GWKMWW56VjMn8nhcdpyBS0P
2THCQIdttwH7fpehGvqYPh7R4nfNvSRycbsmXzFi/aikP7FZq/uEnnLoLuNEBhne
Q4OhwZZVsuS1587vlvR10LMgymI0/1AU3KSTs3zC/barvM0uU78sqqtjeWqXL9/K
80pukKx8JdCdDuQwmHMhKOJQW/dZIKat05+O4LimC9dyC+DGoc21TZkkda40eD05
A7UWJn6JHW+uckBR//DbS3KdKI399275kjDt8M0qg0ARiDMpaK18Ayr6nb3A5+wV
/asRDNENgIS5mORcEQsYy+wChg51CfKHvHXwI9nC9P1ph4UElfgQ8IDthKPHqmgQ
bZYdMuw3fjqSOnh2Yl3kXilJLJkERC0nww9PI4ITge4tNRaeUoVlA/RFKC719vE/
DHzXaGhTarTReFxUFeUistNh2MdD/VaLf4xZ96c2a30UT7EfTYLTn1Tta4Y0a1bI
y3hiYD2eWTb1sQ1eS/O3cEgOd0zlQK2v1LxIfxXxLWeKBwvHEgCW2uRqYo7ZCS6Y
yn8/V3mGjobGuxxUdx03czGg0bkgPYwpTVb+pkAbnU/CaJlzfnFl+Zmay99iOo6f
RU/GBQkuLy63sjhsQVW1YYHNljESv/Bgg444fqkT7/Jd8jZnL1I0P4bGcG+lli8o
Wl+74KZhlz/UqXt9aydOgXCzwBx0jVQOWX/SykuOlCXgitBfUyT4EYR1E22VaYsV
DLdUap4HVEWm1IIt7JocGOukGZgmeFlPxGB0MIoSbKO1LYDIG16eqNV+TU2UG2X1
0MrRHs5Fc7lOE9ZPcN4tysP6lx2irhra48MMv+8Y0wXwJRjWLhO02DaC4iZJTDj+
DhKiigpxYfgvq0MzLE0oSkAeLW6pZb9rrlu1yIMhnNLLtVbIi0Y+5hE5b4ACeESO
RsMJG3ESJ6W4txI1/en1rxCarxecl6B8IaUP9yAK6c4aDbp09P3Uthxh7GzzkQZh
FovaJaAys+XlAzACkT3Mr5xIFKWNrlHedG3Xv9AQ8hV7hEJXMKm8e8J/lmCi5lyd
NHlWZuo3h5TlaRw1j33+QjiBUAQ7p/h3Nt5BcrOrjUA6LyMViMKL/c8EciS7Xv6R
lWuSBQdJydSww9k3OjuQb4J5v9eLaBpQPzzagHnOaX/HLeN6Bc2JZY0pvcvkLXbQ
Hqia+cKv2FLcDyuSX11NPsnRhQURQrW5OOazaMLTKHj2NCdSOtWr/5SgrJ2HKpgZ
ztrEmwBenitVX1cwlMdCsfjj6kuVcpYYCr3urnA2eokDA7OycxcG3e1RQUagZDo8
gDUtYtcIk0JqgrHJqdxWWXCznX4XKG6BJ8dEQGnQWhLgtFhNDlekuKp1jSzfFJNd
yYn0AboEcsHs/ULlPWVH0T/MICFqMGN9km9gxXBcubzo4lOtjBcITy/adGRMn/sg
K0n3QDjGrsI2zmjB9l0btjdOKF/VKPBq4W0HQNRtfeRMSnJnKwGuL+C2XHU/lAR3
wUhBWN6G2mFRwmwp7EtxPCpriFrBAYhBDA84+z2UEo13vrXi5W3o3Nkhe9JSJ5HX
KhC5nBYef/wQl6Iny9EJ5uQ0UMmAvZamNMoHQEViOm5LtsGfZFg9sjQaDuKMCSTJ
ZCrVoQsN6GcltEe3FbXwnYEczlvp0aejsqQfTzNfH+HdpL27EINuLA9XrxMqWyS2
it1Ik2NHp4jp2nerFrtHNyf5cd47tb5NcbxkCH8/yl90Pfoo0efaS6US5hW42VwT
xSnVFnbA3AD0mW8q5tzjdetxKJWRxfTkaVQ80ppO7IH6scithGA6J/zMTJTieQSe
s1Arw7RN8xr0SwVIoBc2gatfhMt5AqkOTqIrXNBRfrEmXMmE92rbx1wKa01yLs1u
8P5GVx6FUTdcVbE+GfqpC57ThVrDrpgzwZcfTE5OAXUz3zAaDskRve7wQyYhUd/9
sqfbQ/HCbyd6H1FTiAklkFLXJuay7rTCk7Ing/NR86sqK8S6jUnpJkKYogiIi+xr
BL8qdAy9Yey9jg8XqlyRbTULaAK8IOmrBcf1B9sv6BVALNPo6yiCIUSqJzlHuH8h
KIfIB45xOojxgYpg+jcZWQTVOMJa3fz5wQGFBEa0pmWryMhV0mmGRmwHjeGU+ON1
SqMOaz64erG/54zPufvAhklUYppSuy2xhP8Tp1kbrt4PhD1M2k5BACItdV0vIM+H
I05IDx6DkxmMDu3AUpewi9tKsHJ1tRp15X2OnCYa8/LQrU4bcnWWQMA/pq7VkylZ
wZ2e46qjMIV6bjDo6GJ2JnSWJHI2uIhQe152oUUVXq8/qWupxdZ8eZaOqphPVgEg
SUzUIrG1boiBEqBAnS/akKdAovQN292soqHhHPNUWeGdqrgC+s+3yYF0L2pCVvB/
YTibmIuhdnrg3WOeoVlAxyQ90hDyN7V8gs1Ns9c459yXNbk78G5f9kTxVDIVCgfQ
46YFi0sWnpbhbquwxO1gEHUgdyeLaa3Rjo8xu2AZBclSZtWjk6tlAaDsLXrbXHTg
+aiGUfW7O0ToCDvx/fexV/bSa26FMZ6d01wtAVrKnvTEbI5/GgOD1WQYpPl5lUQh
3C0onthgMv2dhC5uLGEnhkr0b6nLz9iBI21MYjC18cB0E94kj813w8siqO+/DfS6
5ElWrp+wJBMhl+7MGexwFknso5g6OTdgrk2b7hsyWXJZyZKbYfMjwfSs0RGu+XPh
3mvqK6qfH+RQ/SWjv8zxmppQKu+W/Bb86ONBP/4iPJW8Tsq25Z9Lr3DgziqVAcSD
n8ePYjc7C4/859m7/YLe7PWrMzqE51xiM4TW/9ZtBP1VqKt5d8w7NRhBTQfhOwSp
N+h+oQf30nD3geKFbVhcX0pHJ2HK0C4nk1j9HJKgIFM/qleCUhKoVrVaieZzwjtx
Srd9FJYsK4IO98TT1jCXEV/zncPjJBMXyi/LcvqdARN3ZnDQtb4GFm5X+/ECo1X/
Y+1gQScXF+GmmZVGRhSHo30zm006jTXUj1Kz9lopo4ZcrM9FjoGV7RvD4EvAPj6j
i3dSPhDhNdt1QgaJBBGSSpZCexwyEoCQCwoMVaN2lRZhmYCSrlA2Yw0aRDRJOY/5
4YJ+uAksuXevaB9GfTH0zUgZlJkAoSXZJqqObfg8qKOjastu13Dcrd5ASMaT5rul
/4u5pUk3oqzvgEZcgesoKZYMHJuAWxtiwliKcMCtbZEVUECHlZS4HD83svq7qtg2
6s57Cdh+1p2pwC5nXgLBJq7aJbHXXKCEMf/Qtw+7StSOq//xS9a9SDAxON0gwVPs
0WPctHtNe5BzVlyH5YsJm62j2VPRK+A0pg7WJ3r3/ZiFfXjf1KTGbw7vitpnKHby
J25yuDoxyzcZnML8Ln6rzkJvHCw7Z5BRljvCCJcVLyM67iWTAVG1TJxyeA5oRrAm
qdd8FZ6RCose9WfU+NuYGTH6A7YCElpgJC/XTXD3VG0SfqvBM433iVGVaDWioY57
J2FMNaRgvbZPbUZv5NHtIjClRdv9jiCj8C0HFsBKOUd5Kv/Kx5i9ITV8z/jZO12N
SPQU0g956FLv1nwnBMOMDQrzjqrYijnF9aBA3+2UB8/aeTKFY7udFP+nKrx5LdJY
dru0W6vMk4wFQ4JXmQ753XX76dRiQzFo3K+OU5+GjUtENMqzKxvE4A1qbYd2kSe7
IbwRFrenl+d58CuMhmb/YfR22L0hdtGMRyD6LIIC9D/PBUiHm+QQ8yT/yaMlYGXV
GmvSZBxeChc6p6CzmBft0iu11nxvmBH+hUM5qdLO0VdOXXBYv4ZgTsAQEaiQ5K+/
g6AZN8WgArkDCj4W9CWlBsROVYcd0/kPoiHpFSVTVodU684EfXO2Es4pkZSH729F
XvGuYAmWi1usk8IPFddr6ZDCRpeeaXfVO3X3b+Dwdth4k+QI4BVwH47B80xPXSSG
OYj/kkZY16/uy8aj7/8RN8/VqZRFODnc7ACmTSkzJzjhHgJYu25ci1QVYjJ6kzQJ
zzk3sgpLJjbXjimH4fv0RbVlCuOP+MYcq33m0eWqFXUH+RF67kMABWNy39led698
7+tL0w/VajLMse8zORmi5522C7GdNanHCX4gVaZu3uNhVjGLY38E1YnB3VZ7uADe
8QxgFnb9cDWphj6TWhCeJpgEV/TY8Jofl8m1CrFjl/QSpgt8z4BMV5MXzSqSetJv
RjRUUYUuEdwqEt7316FS9w4HNVHRY+MQ/JfJsS112W6AtUPmcvS88eLUA1r5wud9
QWqxU56g7H70cj0YAtWg15lAuV/zjsvWXku2Ik72J1luPiRDaaWhTDPVcznyqqTr
+eyDab8MZSkfr40bPX8nPXyZg1fUF1Reh8NNLHsYstPkqHKwpW816xT6eprO8V9S
HI37w0SgaRIjWbd3RjBpIPYMY0bghDJNP5EtRNEehbzRB7l/xOTc1hJ68ujxuxNN
BlAuCFa/W7l4tcLF1ooYgxx13i07T2wIwKlRa06y+D/X5TrLwluZRK2v+G7tf1ni
WOOPgPvF+7LZqaSHT2YcPFfUSbCa8rsoBft8V1OxH0RoYuvkmDNkQy15SKe9xFmh
69TgM/eF3JnTUNZUwRx7ZuSl4azYkEtSUyO3dL+BL4/7DH69KfTkIVdW/KcTPPkF
fAo6boG5I3/0nkRgOUzuBLFF45dgXemD6Fd6Q+EmUJMJe3AXvLk547U9TtUKqw6B
Bz1q1B7fA55siiUmvASkv/mMrMWfc9D6aWRY24nKYRoE4F8SLU1ZpO4WAZtQIKq1
C72aiQFrEQp+blNN7xMRaQxO2d/uOzQf1PZtBrSU1ZCHiKKx4p0dfQerQyYu3PZl
7w3GoNoL5ZAdZzxknlv+mU+a+KdTeht9FrApFA90Rz8K4NZOubxPHFvQh34NVFzd
IPdIoaJU5bWEWj2tKUY4WCRXaK8CGH5GnEahw/rrC39gfMbD1oXyKyyoHaecc3sq
eL+jsAofdOGgIj5bOwyx7a3Jf6dklpxgECcK1P9u33qqRDXLaAcXi+HouUfO+Od0
E89FhlmDxen6zNvtn6yOsdp/8YEyKZngrzro2xWzIwrnKTAViaXOxuVSv/gZ+pgr
REFS25AnwhsSyX+ZZijYXpm9QOm5b4ga4VhVet4LWQbYo47ffnnjiTOTRBygx3pP
eSfwbpueg9CNwC7Wxu/rLqz1pCYJSvoYRj9Fx8s17HGKNzeKGUiv95K1fZTa7U0i
gzZtdfM2y94HJGLne7k7tDAMX24siG7SFMxhR5ZPnTQOUFcfEpZGkL4yXzonc60C
MNEcBCl154d9B1PxoYXgaiSnN6f8qYPHlPsv/GppkL7XQirmz2cZZOOx3rvpvVQv
7o5LIY3ZwnzQe/xMeFIsrkehWctpNfNMd9iWYtryjJFokrcLG6BBIj0O6XV/Skud
erZ6NC45EolATGhYTCmSul2Cd2F5Q/9PizsaB7t/RuXATevhvNEEO/mkiRCNSjW3
8p3eUTi2feiaoO0VGKrf93ii1mmIo4eGie5QopnkdyGzI5fN3RYR65/yVGNaOMyN
Fw8n2gbmKBRZPTZSimTCu1nA/J5mW4JqdkVgqUlnge0rqcR1Yaqr7accTuonQ5jF
dHkyzMcRPTDJnca9svuJ8wv3NIFYBLxyZMYNgf4brleLY3G1+BuVb5iaDjoGQ0/y
0HY+R8m197OJgjBPot1kZsGlOQl6zOWEIwASp2FL8NtVJfH/0bu84tRt/5hdYYB9
mqlja1gZV9PrNVQZGSVK1dc2k7FpIHQHDT+le4hMyp6ml9qrnfe9UIJHh2Sb1TTg
qJGirqShABeX34s3hKFGlvrZtLKtoGyTuUhMxkDjGr+Gq1Fxtv1YQJ9HIu9geNsb
t7oz+chy/VoI6gl5nC0z8Ws9pYWs4YmW/xfpBj9/n0oZFZNOCquYtdopkCQEgZkR
MtanlyEG+T/rLpdKam5728n93GRlYizt6/iEVTiFgDYWWvfjVCvm1HanO5NGDOlF
785Ysv3M233Xlf6vbPcINFcMlARgcohYTAgfae9JB3dBnqihI9h91qj5psPxK5og
+qJxnI5ETo16PVdVvAPCFU/5bSABmuzzHzg/JuVteGIe7mzbhQetv/DvK+U1A6T+
ShdwSSZg3fvJkriniHW1rEffh4dodzsqULzKQli6QqmrAEzE6yTjTzq+keuMN8OC
K055D7J+Osha/n6lADksC9/LxKlJgKj+Pet0H2EzsUlDYwCznV/g/2hAClEWShZk
LO4DjzXmqbYw8hEbjyAmYFt0x/C/pGVaTdVxH5pwzjGYkIcwei/4LbQrJYzUdwnK
pdbDmyQH1K9oEqlEDh97nguSbRgYWeKxas3uC/X46mwV2qnflUliiOZ9r0zX2pwk
m0ufB/KpZlmZsirHnxMqSDc+k2ugg1kxl/H1s2kcq9OBJoJwsr6/hSqi7utGsJw9
IPU0RGHTrWSev3CYuPMMdmPclvrC8GZm2K3Be6tru/cdvb1i3mZoUAjY8HL9XxRT
w7sAhxA3iYl8ePs5Ctydy/6EsWTouWQOG0L32GrODh3blqNgqWCueBqBRZi2S6FF
`protect END_PROTECTED
