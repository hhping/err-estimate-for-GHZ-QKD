`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OEgr7C1DZ46uOojYExLL8wGyfgUFE2U48Qd++dGleYN1JHr5CXly8wPcuuuSHZVt
4vPef72OMjUcO/WsVcY9z1+G56yTP+2niWgkABAG/6aOZj6GYPEEOaXVVgKtEGk/
iEchLDp+bDSHt25kDMNuimxmX45tbnjHmBx90WyWXtEc02FVJXbIuJqWyl0cfnJP
2LBpqX051dfdZX4KMgnazIMMac33Q4WU5Xey5ejDclEJTpo5g8DK3yT5Y+pZg0MB
2oVdKWL06p7Tn8mS6tiw7hekHfVJmBjaY8f1YKWjdVWjzqNnzYnOg+c3cktUoAcC
P3+/okNnIB8gEhOgiaRDjX9NQu54ERwo37+6DcTlzggF7BL/TLUTP4hXT2E9AZkS
y+Whr3fZ4Ue3aWEHPUZUlkIabLftUWsGqQh1Ij/rWfAA7BRFZan8xkmLkRjNJQWK
a1PjCAToDXqHpWgVSRsCHURs7+6TrlFCDz7avm1Z9SYExvVvbL5MUvF6L0NIQjyD
ZTXbumBErAWHzblS9H26o1qFGyJQ7jfRz8DiBRu4/B8cJRLIScWBiijcIoUPRFhK
UUazjj9Ay0nF+hAprVBLG2GugEEpaH6FQy29sajGdSsb17Y6/T+qZu6H/OA0tU8y
6Lf6UHE8rjQW/IlNDMui0tSoYZI6QOujMJRd2x/COX1+PasYhAP8W/pI321f6G7p
BU1UOFfSc+MSJMEV/cUF4yNbYFLd5I0iLGgC8ESXD/1lxdc/iDIda1xQ/EDnBoQ/
CXFl+WZX+4+EOoQ09tl4jwCJIOFwZ170K6LV2+jzFw2PN/plXgEwenXOa04ynoNQ
TbBo7C1JzhPVxjOIahMftqgLGuK6kG4HezOs/+6EBEh7TiN24qnZ8ziXgzC+1EVy
QTHtu8NzXWAvIMCV9ISBS5g81ncLa010ON19nSWgS8yhMFIrSILZ/IrguDbFo7BK
tTdZbAQVOKseH5ddr1B6eXROHFwM0XvNOTubZncB7rz/xykK304ViqX8YeSk+nBJ
s99PqRTCm245W5rk6mFVHqfKF7ivjoTpIh3SNkFqpK5lrOuy/x36vWNYt22Ja505
7AJxmSENssXx+5rhT/7oTXO8Xc65+AUX0lNTY9LwRoZ7HEfCd3ddkGLUiGRSWcLV
P6bgYZmw7F19XExKMF9mJ6/E+J2CP7Iuj9shGo28f1upgFvUN1VBGPu9D4JtArf/
3JNaUs59B4lqi4YxL+FCIGvfaVzQStO8UHXr+5X90EsS7VmyFQVWpc3XQcaIe54V
AtNWCn9voq1j9WuXBhRX7jYGmRjVBKVenZ9clRNdBaL6FAHPOvvPTSQOS7+XG29u
GEu+qISyIUaWJKNP2lykaIKdMI0Oh6IWzLgiDXVFvNOWKuVZE2Id92mxMqEW3/H/
Ip+F4k0lb+jeyrJYy6mYzRPf0GTOLhX6XRGBHWgJRT7VC42lfZWB7x5Al0K4Vbif
sQJzZlEmLTiXtkgWwAw0ZyAitnHaxGny6dpqi+tkz1934jZJaVST4w37fzafIzqY
PH6E54Y+FBrbTbFAOga5Q8pDCmgSwUtp1T3QL3a1OstsbpNZmHBKiGozs/pGnatA
pZUuGmwsU9H6D9JU70P6IM4hIpgAP5I4sLneqG2cPYCEEppb39WTmh9sKR9KgstY
M4aNQETi7FbQnTNO73X2Rl+Yr7tbdzZX/dNo3q7cAeoWk5/DwqPIoPGKEb6drTuj
RFX1TgfygY4IlH7YmdV+eQHqYMGhSQIkoIYuYQmx9Uwbt6NVv3VQTMBw+OmqOWgR
q1O+HobWlOn1LQ56SI5kSCU0e1KfQKzGfrRz01kLNxxT6M0iWCXcQdXVi54SiDoh
KGQkxm5WzxGCJ2p9AFFbyawEaa848AflAVGQgiPu+Mz9dHAqWSocG2mtstpY8du5
vm6Bgp0qUxplmp9E8yKxUVbFwJsjqYFNq5xgY8UEK0hW7AtKzUQD6LJyWeaZheCK
YOHHdNpfZTJ11gSHkLoSAa/3/NtvfPUNQV4gky4EIbF+rhSXbri7iacjm9Uj9sV6
os8nIRQDjkiL8pvz1XhSN6IBUf0a5H3hIZG/feIvBx8ik97EftAup+S1ae6kUAiF
Q9OpszrSVPgXjLrl5naz8To5Zu2kqZ5C0FmAB73hTzmkIWg9VS6ktKnVDOuF0xjW
vZun4EYbcoHQzxim63vVVJKNbT8qPEGey/WQ3cI0NMMmUmXtW4Z+qBBqJ/N2+mS/
NADlyBe+ehf09v8oD15HdHzjfTM9xrc4FEFctzhIJf+cVgU6xzzq/DXCSukzyccP
g/TVsTfY3prpj6FWDHFK1BONVYgqG+v/u7PAKrNcWpfC9nP9EKHSiMZ08UJCucDM
nokCIzTAW3bbPNuyfUUvSUSp5nmVFbG6gq2lcck3z58EseGt0G9ow2KJy9xwaIZV
XKmPt5d/6+jtlFXOJ6njv7TTpJUGc/vg5rARK15xCR89kVniecNZmyjasVBxXReY
MNpA9ipvtT1AxYzol2rn20YCFpP39+s6uRBfcO3+wSTbxkPPxfrSTashV8htxuKK
NEJQLHRejboA1JgmT3Esly1PWi4QTzoT84+DPv2iOQWQ/t1ZqphWeB+5XpKwjT/J
ajUN75fYUuJ075eFaRNVDYYt64QQmWHJZVmnjNd0gxE=
`protect END_PROTECTED
