`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XNg33vTqd57lMrZ2psYAQPvexcQh548DGsveaNZa1Ht62vx/CMVRW+tUdldbREEs
cHqngvHXFwEJoyKifeu4QxeW6PPAmULXfOAID8T1KnbncKdL7ci8he1l7w6v8ler
V7TZHUvah3zyuY+V5C4MGWqCMdDnNQve6au0Jlx3H4/RiqU2bz9gQQrEydZA+VWT
MOypzYkhJ8u29KKZI386IBU/hy2XRMj15HgRUCzNOqjhAdIt1C5ZWhEthBCUswtw
jV88zwMQX89TAXW5hZfP5Dx1DEfUrAJwL9Ifep4g1OxODkoL3BwTVRAJGa4J+oDP
RDc3qkFN/B+gmgJzNimpQMZAjJio8cMBWqcb87ILD3RVedcYJpfGUzey9uayKxgJ
6F6xv+6ZKWyO4iupn0ZNaWff7b/vwSN80LTcfuiQxLn5RMu8WiPG/mfZouvhO1qw
B77g5uK7gQ1/Eoo3Hyxa9Wq5tdaWP9zbnwLOl7T12nGYfPZZkB3jVut1WKKh+QTN
QJK8eUw8/Mn15SG4zuIjMOKz+i3Ul9XBTHmmrGXoadvMvdoK5WP1FaZrSeC/u5SS
e4KhuGtIB+nKNoALIkLYLI32MMKqny2ocOWbvXa4hzvCM7S5OZaNRq6DTmuGTR2i
xOwQQWu1gY7+QEPNqeGpnDUTuI2SU3Q5AFUzaGHZeaoJmxvjg3w6XJfWEguFoRfq
B2YK+cRxbl9vCTCMfWrHlFrJC4Dmr5q9Xs/Q5w/N1Qqu1bc8V3JAQRvpYpNXAQnb
1Yhl4XXei7/uB3KO4brYsxy6z1HiT9DGvcQ7o73rr0QZE0Eqed/yt6WVyO2Meeb+
TtdgrI+Bn6VO7RXMF3zdgPqo+PaXjKOGfkRzUu7Ba7U7MlrMCm8+6iCwI2CPBdYq
qI9Wxo7H4Fj9+GkoDl+xUHOdg+A+HtBIc5EP5eUqSMkS4h1IG/JfSULaFb2qYO33
jLbgvKOx7pNVsikWviwioVsTp5a3ii7NkGEPgdUOOCOfWmXakNrLCEMweH6jmzzB
QtV70eUV8BoKgQUyfkGCZHOuPNfyIwfsWMVf0mgubCTHywi7iGyWMJaHahaAJmf6
llChHmJqayXez43Un1y15MRHH+/muGfHvFw0hup0UffRV16Y8uy3NTv6ASC9dW1E
9PXjIaZX/8LS6o52yWjumLGSM40TJtPvt4GYrN3laCGtyTVCQSeGr0HXhjh12/Kw
ZPeX3MugAOTi8VvYovnQPePLVX2BiBq5A/QATrvsA3A6jz/bT7vPSii5DD3V78fJ
hLX8fMZDMMofBk2aOovNJqXJ3f7dJ2wDT0LsA3KU7x41AFhyeuXhxRfCON62sSkC
f3Le5EiUgIn8kgMPA1ml75mL5birPo7TURRBQpMvDj/0Fn2koJ902ozbGWk0CVhb
CICW8uIi8x5aiEQcxC/NvO+unL4rf0RRMHO8/s4dYLBpq7jfLNm41B0X3bHtMZar
+YSF6/U2eW1W4UhEjnbTGhsfrCoaUYcLJ4QJNGaqP7ai+6rPqToObkfUs2+KtQQE
Jo9k2GrqB2bPZJhw3zFKMHA9Y3Y+GuSubW+RTIFT+p+bRIAyw6ZlbrJnW+jFzthy
7dO7Fes2HUwRrAeDv8MzAEmWRapxd5uteiAscv3bmLG5uvxN9mCMtsT2deBszc0X
M8v5v84jxl4OW0Pvk46MFx94Tct1kKw2FN4/2sRBf9KSRaTELJMUbj7MFuXjeKhe
lWLlXJMkgAUJ1wdzcypHnYKu8wKHlHMhEZJdt0/BPgZOC0w53s4Cw70zhSozuaEb
QPzfNYflPF9e7Ak0rkpQwCFTtVeBvajjcE6WSuM+3O1Bkjl8Wa0RbQuthbH2QxOd
SGsgdamPLCRpn7z+ipOBlNxKTV4Ds1BnzvQRPD1ORn0=
`protect END_PROTECTED
