`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WVedCPpqdL/8GJXas8ByDzaa/9XanPKRD+L0Pp+4+ZqhyFoYc4yiMdOuoPugEtGx
4Skk3ngDhyKtJ43THqUuivGC4xDlgC4k3ua7ZWa+3qKtI8rtx36W49hJlTAJcDKh
fetjemTxCXUssBz+9WN3Iw522UddxZcfi9T+pV2GX+8bnGavurcMM495Z/IkYT3z
B6256nOBQrvYyJ5Nb1Jnjmy1cx8DncQL/yXjDwQ9xAjUyqot4VXbJqaVex+hEiF1
J3ZkqIBUfKrIloCkUVnI4cHZa4t2djwJf2UpD/w6ixlh6xr7og2q3YfUuZQRgslU
5C5B1K2ucffkXLQUmVJBZE/nzPQYJKuLjsBQnFtlnjD7JaD2ZL73UEKWezn3cu8u
oql7poxTYOFxp6JHVvvDN2Goo7zQNdPvhaJ6HwOynElr18Gc9/6ACPkMmZ/1577f
I33yQ6t8PvmpPcSNGmbi0Pu4nb1g9fOyJqeoxmW/gL0B4oKkjn08GtortfilgJ/U
svb+qZ5YxfsUg4uopgA4xE23H7NQFFq1bvt48pz2J06mb5+LLTgpOdMDs4EHdY4C
d4P5FGodRzJZhLargFeKAxdXqEv5sn2rWL1KP9ZpLfVBo43ad5I0n5qneDVPgXMP
ePjTXU5PeV1uECoGjm20BggQHOxC7HPBT4z67cjeC7bRGh1MsrF9guRCjUNyFYcW
PbeLfa3qtLxx8c71AKSzd1NRFWnFS+k2cDt0/5GeW+iSYjpyZgwXUgpP+8uwO6RW
4twg3QmIMD2Q4tCJ7mDlptzxrMbxo6z1H/EPdDbalS7B9RidCG2ca8O8dGSqetQH
iT+hW4mFEYaBux0O5UToCaQKh2AvyS+tL8CDVOAvik7V+GtvyoEiCjd9ZGCOxYad
qzOLhwMit9NwfZOSj+ekaPuw3H3C5Br5reHP8BzWgBLdZTMeYWRJGISi2ABgjbek
8SYJ7oIO7eP37uOxBuNGy46UH5n50oMthnn3aeeyyjAsbzxsQw8cpmR5E3J6sH7y
cGWefg6gjK8K/X0bmByGHg==
`protect END_PROTECTED
