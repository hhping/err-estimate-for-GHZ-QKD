`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ktyUztHPCLSAlBuuVbKpvjSjl9H9yrkHO1GEH0Zz22kn0jQUthZ18zrSn07ikmt4
WgdhhXRbrI8fFXGbOSMXdgoJIOfVMgUmmZTYB+FQKLT/rRPkgOE1mdGo3azGTYwa
uuJw45vH2PEWqnFyabrlndmeec//GP49oSG3hQ1U40Pi+l7cdq3UFkjrZ/xQvHcS
6IDOg6cnx39W6RtHFGD7Ja33uNMuDYR8dlJVFg15k0G6VfPc8Jkxsulddf66fazl
t3qvCCadiGJg0BvkG5tpcvgt1ehXvmZf3MdMBApBKWDh5XXiF+5vD4050rYjuhFz
TRc2XNv95CpLNSHQ6fWxgfgOfj+IR0kz+IhL9DmBRMed7UIdppOulmGmJsOF2KA2
FtmeVKjR+csBdLiuGLIr37ObtzyMm61Xa+8WZU8YMBWRDq5JOA7G7Y0eOamUiBq9
3DqCeCYTcxNqOAL+qFA84KJUDAGGrqTCWEChkIhxSa9SP/vpgB8R/cSwiUbumvEO
35fgRJ5h6zblW4G8HfY7v+mMRU6Zy36DELfEldEDDOnyVQLXBM8Zd34RrmSGwPh3
6VZPHRV8HUSTN0AnFDCVhDs6xpoMbsFipk9l4nj7STK74YP40b2CI+RfAqt1HpR9
r36cKVydo+MNZt7mNqtEuqZTkK48f2Vjx7RLp4MCpl8Rfj+j4SLbzHpT05WbaMGj
WUainBUfbZPi2FKDTDBMsLOUk1r0IRZY74WVbS1iG5Rob9X5dn9nUHXweGAir89Q
9zsjyNXybWEhl2iV0w65o2r+R4UtaiMKhwjNUmglZVwQNgRZJCozf6LqAJ4qNzdF
gc0ZyaX1ba4XulAUGALYZgRsIxt+gLhfYkyMlMFGeEp3UpI71VGZczXvM5INqEUY
`protect END_PROTECTED
