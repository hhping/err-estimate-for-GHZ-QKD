`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x91nkQU8UNmwzKh1CQ5dq4RRn0wyhPDj0IUCZUoftLk0epnFMF5nHzDm55wdnRG1
a1CZaRSMcUYg2IhHcDhJASqCm+9+wVOjjW32t1rKsFo8lk0Lp8skC9UiV5PpKnRD
pTpP494m/Hjnw6m+bK554clWK+g3Odga0V12X96c+Vh/REV1BIQh/YiXUX5LndjP
nkjQoRNy9hdTpnl2SPolZhzZE/K4SV4R5jka3DpQ5kUKBKIO67Ax1FgzSx7YgZoN
vjN83DXAD1Mf94CrVB1ekcHdLvCkHjYXtJQdoM1ZcQLWSKK7J+chO42fe1Jdgr0n
YOhu/GmtR+wfyLeRX1UEF5y08X9IBcxlxTjyQH9BAV1kyK+pmwzcYfZfkvaTlhzu
gRjwKOzOYARllLO8R8KgWpd4Bligy4mFGmVRfQyIHPyFx3myFTQgOs+iMmuQBdrA
ofI8kitN4JhdySA7vq7wVmdYL5ZFsZ94WFgJvFJr8PRerYvok8ZfOYhfKBs/31vX
dtBf8P025FaCk5wDAEe06gnw2GM6CnbuQBe23CFkL/eKK9Jw+emkP2zgGT30lkYN
mxWFX2vAsvOCrQYg0L8ROClnxEuwYxuFEDxrgXE5wlsjK4EjQ+DyGqV996mp4j8W
/ZkJ+m7tZFtdny3Q7MsDR+xpSWOMmVHrelYquqJRdG8=
`protect END_PROTECTED
