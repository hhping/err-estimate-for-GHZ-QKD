`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j2V8jFSBOEPhv18x17NYYrrGOyXGAVAvErUN06dmjlmJ1UX5Nt13Q3GUehY4HvNP
pAlBqQjsvVFIOK6HdHPbolnMHma11/MqQt7zKx4fzK/2V/dV2rg63tjM66ZxVLwD
uSKXxx4VaS2xMacNr5PB2om0iqFqpRJtxSLj6nI9velG/0EMzU7Ad7oJuxSkzgq7
7kCka8imzutY/wV7T23UL9LgsFk2ouXIic3OMqGKvFFH1zQyTdnzUzt+uMSUrZML
EXNkr2aIAraVBZyJHKGrJgQsZh7b7orH/3GQ6/DdqdgKAlaR9b7aHA1aqYN9OJ5O
0nyZtPKc4rB/fzHFIGDhAZGkDIuos0xjyo+wZqI/qpTCZFEM4lOmq0tZGYmAAocn
55AuMWL6i0vxP+m0cgv8+2Z7ugNbfeV9r5iYvhhjrCm9mOOGeDcRRzlNDUKAAwp1
YYneKv6z2I7IXYMO9PU4mNV5pgMQtxOU0yIu24mJjD7HQk3SPVKhe8nn3xbiz1D0
+vZOqzwUAtft0FTZSB7HbWFOF0miJ7j9IN7kOXsGtPkkhWRzA+R3VjcfX9leoIbr
OSbp1dG9uyEwXzQ6lStBNm9EAso1GNypxwipMZ/p8AYxj6DKjSfmFKU7ifBUQtEf
6nunCNOjKvfzUgHursB392Yxz4L/4/Vr7tMW3oAnRcITlvo5Hy5Ta3/jh6x7HIuS
PerqB1LmVkaJMJ/euZv1eZCZ9a1Zu+PKoKAUwLgTvpabLHpMB48mYHSiWk84Cyb+
af6lhhIDS8vcMiEhbj7AU5pyZcTPH4BFAiOpw6/BLC1HndNIYCdDM6vtNNClUN1u
n0XBX4/x9JDliS1050oqgfNED21GDSbRi+tadsac6aQUBYgPPKvQygMB2roY8ej/
OezZ7VcKjneti+Be5vczxTl5yxDPuH0H44ta0/bOhnRDej8flK7g1cq79sNsCv8p
Lc4kUyHcYKptO2rhrB5djTUfYPzBhEcQrKlUzHcl7CV3uK4Yp1cKHEZP2/Wt4Co8
BHaU0haSPHEVq64Rt9QM4vxTddkNOLDEBq48jNPaFpnUPNdyhduYHXTd3WzS88kh
P5gPdr0p/jn2yq1ET+A01uugKXbwpYQ0Aj42hIYzp1s+kWQmSKN/9zJLgODyIiRl
c24T7dTJrd/AmlfFh1qYx90ZicIl3H/1eITxtg5XQ4WgdkzqlzUQNlvpehVYdFPT
xbjJ0pQAAS4JPRNmFBX6k6Sd+ePGQ9mF4a5VQX5BkdUcCAEGyKjE5ZdD+pqq8LrZ
vOMHDcYMxMfc8Rpbw4hJ2hSFYiT9MdqVdvWQClKuaD/Y0OVKUREzSvY1/pjtVM6m
E4KCtqQ8MX0R8tjoXxD91Msm+phTRiND0fAZJjrbRMN5jxkemh9QmcXDBqCc05Z9
tNuLE9mXui+8Pt+n6NkaQajS1VlvxjdCn3N2l6UPT1M/YEzAyP5gihYK2zfZqTbk
NGXcK59/ou+avPplKo28vp55Y6wxXOldTNwJ+/JZL+H6WsajUbyNlpPoY8HmnEof
DLj2bj10SXvbDZCK3nvKGIiI3Zxwsz1TlG4pAnsKYwwhHn9UbUtwOc4TOrLfkUSE
bEgbx7M89RwNXg8A7KSjxYotelDlhByLmWnz0QLuO8GFA16YiQXiMqPtegc3EHhe
Pyeot+m8GM1bGuSD8KScKw9g4fexfN4VGav1Lm/E7QhxsM00rCFBC0Of0fW5yKce
7bQQuDe5xNsV4zIlXc0wFpiIbwzBP2p8Ker3vd1CsRbheR33IjT+0j7ay1OypiLn
I93G18pjytSiKLf5P/siBmbH4vBucKtsKPJMj97EGvExDpbUWalke+jSTYamOM0i
ChfPhhwS0lqVlMNjsUEd21UWFve1jGrSIJo/7l/dPNWcffWkkGUFVpqYJfwLGBd1
HejCMaBZC/P+nDZnhoQw7lhIBGZ316Ln//b6jf/Q+xGXJXqCDk6e/QRy3TUa4LMY
WyVoaO4MFswaPAwE9c/LEQxbGOJPC08D9jexM41IiknxWftqrWkZ8svHC0yFN/hh
iFcL59j/WP0QrJb3MfvSPJR3sWIq+cJQhNUtQ3hRS91u6VDz8zHawtHusD+HwdFN
Nvylth4ZgAWBvULNPpsduWcrOI7U2CUot0SkWa8jukM=
`protect END_PROTECTED
