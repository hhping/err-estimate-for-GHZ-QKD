`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xaqg/bqxgNWLIp31d6f3gezNBJ6skUDvhwky0IS8Qy+QKJ+i9zeV5QSLHE8svWZc
MTOuZ+ZUhZLyPmqRQV4/95CsAGiSiu/XGLZEpLfw7wDeSsSVpVbEPBlIDwXLOWSn
bYLnQKfx3R822906bgu/d6xSZ887+k/cXPYg2wZhME6h/19l1fzuhvQa+GrG3tNZ
b2+Vp3yxPaASnfpkbMIRtSuZRGwMWk2pW/cPM28AU669+8U0lcaOnsFN9fCUeot+
Wsk0mf0eHBPSUXi74/x4YkMUYoRuFEjSLCM13prLYCbmZY4VPpqsI2YJQdDN9AM7
hqB2w4MZHkHwWLxIixCW7HGO6gkRN/2cqHygz9xJrSgwq9LJOh1ydvDPSQmWqtCX
8XN4pWP6rv47mOLLmYIf3LWtfcwlMgT+mFDtFKL9511B513gP2e4jYqMJOOQJYrM
L+FumbvqWSjQS5gHTkO8l/k/VvwErW9wo1KHSnBYLIRoYG3gzXXEh7ButDY8QbRL
InqiXeMkNPklRE1nAKdllnRFO4V8sxVMCzcoDkVNy8i1NwTVnQEyhkyWmUefISPn
ApPylDtZ/6qKGwVL31y83Uu4upS5LX51+p0PS59s9oQiA2D/AcZPIx7HYf8Xh30D
emTo6z1f5DruCCmy6zK7Qg/+SnD09NZjVlF/5hQyFgugdkEPxDRQ4/1+GygXE8NY
5LB4NXOZvRRuIifv/wnx/q3Ku1+LvBzQNUxsgz1RHhCJ2KgOHyyIiwgMT6yEKvBo
Gk0FeCGiNWXT5WNFhkBn1gpHf7uJaO02kIam2wFNBZeLMN07UvpXPhOEdD9d1D0X
eL98Lh0bf3VPhuUqrdRWrXlgRjGb5HnblLBn2yA5Uf0M6Ps+1Dy+FMwHBmvmoHWv
mOj2Y9d0hflgJ7jNXqhVIC25j9VSEWYaNnAUwXK+qQAICEDYjhHpZKhsoQC7tHm6
xAJXg9apo/VEUgjIJrcD6OOQ9baCXpEhHUGI7D70qVHxWGISNL4rytz94RmTsYku
PpkE/2C+33RIyH/vmeC7NDhhU/H9Wi+g/r8DQLl+tNu9v+0sPpgFJy490twwyOvj
w6IgeWTFCd0iYFxIi1iXYWZtoCInlhs2kse88DsFzQLvOemPYoQvF5xW2V1SZZUO
FiwQjgCOQfPfP7e09Z1KckrJiaNZoadmWu+RwhsaDAacduCYnsDM8t5J0kpYo17V
6qcEF1zSIFs7DREAS7hAFn7ElnrNQK7i0hXcpRLdLfTdHjTgQZsOQTFoxa9uF/zK
tPY7/xG6T1n7sRCO1e1+huAnEjcIwhNRVytXIktxLeXAiYTTHoOQRbMB9VaYEaix
TXqBjYUugTNvKaSOEqQLEsYBY83TEUzozOQ/yhmeXr8y8pkA6AZ9xKJsV+kYhnCR
3e/ng+dHMJm1+g3tRWLehA0hbWknJEaB6wa63VzhaizG9vbplma3E+xCEOy159I7
+lrHzArUHFAtUBTkSxQuXmlrdCvAszEWNQknqvBvPUFb06corjwTK+gFsJuhbjbD
5JY4WKxDB7wFhKSUp+wD1KMxw3saq4vzLhpr7HKgI+npCEL4KHUd76RTQ5/pJPc+
zTUICgIQkOpGrT7ybvZCQOUZq2yL6bc6lol/EDC4sMNpMsqOS0MOQJIzXC2m9sGX
SPmtQIUxmXp+xUA56Tujeqfo/cWdZQEMl2/WtdGEKZlsUJSFVJPRi8cr/3Ic3TiY
16CPLwpDvpO498bW0kmAsuoJt3mC2iVaF9uKOOxhi5/6aWPVUHAp6k8WRJIexJ52
wKzJbZDjGTdefenmavQobw==
`protect END_PROTECTED
