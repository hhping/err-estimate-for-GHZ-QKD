`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cr/UV6FEEDj1EkYFxgHpFZmNW9B+ig/qgUcF9NvxenniHNjzr4BymYdB7Dh+nlS9
0T7QE2v0ofdRY3MGyqFd1vqNXB5cxtiLOz2lLDOQ6Qo8lt5qk3lmRDyXYKbS/FEY
NydO7pDRs/hVHSNmguGFpcimI/x4GdWEixhkLjbMoKgzJLWXDdNQTbiLBIWgwzyC
yrYXzL1ZB4C1720kkrK6he0BOKBwyh3FIPKiXxy3dKNNdsmuSQL+9QP8Yj4M349w
UaED7hjcUDS4tCBGLOKJ/nkDEmiXNVKyv+ZWceFskZkXqogOEGSKGi732GVOco8z
b59CeK0kzTtbIED2MkkvjyvZdMjcpcCWcXzhmWghzoOr3yYWkAfiwxwWJqnn+JMu
Y/BLrEssxZpz9z+fwC8ZJuIQnD3aBbEkr+hy+IONidZM40DM2icsY0bksk1+Q/L3
Bj/ad2dr947V/LpD5naxb3TlHZf0D1PudqbOKMDHdSQ+hOXxsuVkqc2g6PwgUWsQ
OoGzJORiPsg5oMPbjIZ3s2GitYGKjhi6pF/1WRFVWVfr8A1S9+iolUnhO7z8G2D+
8RQqY0YOLKbT1XV9m41puVAnR+C/5LZ8gp3LTsoQyTiQd3XWbQDsLXLIi8m21Rxv
uovRK0hT1l5NTy1QmLYkk5uupdGAhbIU5f6KMS2dM8ytiaQtuE+UhIPyOAn9t2wE
RnVzZfOTvmmFQ4n0DbTgk7z6eZJRhfhxP2wQB5xHSB0ZxG7AmZoTTlm3I4f1opaY
KNZbvTnvv/U75sl3a2j+RJW6xgez+5reD0ExpSCl4fKM6dZ9/cvW9RHAt9hBLdBM
N5/ls00EkObnYY9Fl72K7MOPNoH308O+03xBq85uDXTuwU0iKVekp+bMfsCPssbK
qYR+Q53GNk3AlLJEEH3OobpsiZe532Hc0uLNNFfpKzXBrDS2SvCvlaaVOvgzNGoR
dOMpISU3niV5qH17skipR91lFjiiugXnuDrEBlXpI5A9qE1d2KTCRN4jIMaYZuyY
SZseGrYN8Tu4FmteW7NrlouNvBZ4543xdFCvDtyFHJD8t7+rPj5SzAuRBVCLOaxN
bkZOMJHYkLP8BWDHeNVSEI5EbKu/mSeXigj5k7cajdVOPXuD34KIwrh8WC7rZAlQ
DvQTRLsAofLPrAUSclZUlGVy5rzz7xz9XuxT1nYrKHMohzBJ7KfkE5m+hpnZ+tTl
1uy44XyWW7vy1sTBZRE5kgq5luATX4xUzQDn+wyftbfG6LzOst6YRFTzjAkz5MXN
DiJ2pR0Cvib/8XqJIoWd1x3FC6M1CnkGZMxrrInNuj+Zcp5+5Wfjwcqz2aY54+H2
qSqDM/b0zefDbQMoDzT3pSQKWTGkmdkEeG/OvAG7KjtB6VCfKnRhdu0+LF4muvve
HsLltC1vymYlxmoDB6oP3sBaww+GjzWQBryCVp7a4EaNsQhgUB2S4TPg6kn/hiva
DjWbrL807jZI/jiYPbFVZjvVQ/JFstW3rq2IRh59uNS3o/nQE5gjRXqvrK7CJVJq
J8Pz5+wVlyrPndk5x3NyPFWwFiA6vW82Wjb8j2+F5X7KBwbpqea+Z5+51cXP+ung
DjlRYsQ8JGNgz2UhqgzSUf9YjOrSyUp7Bghdu+VPAzbqIGmf8kdt2eNVFxZNg0Mx
fpfC458tcX75JcPLDqev/WZKyIDg8e3pj7cCC7nD+cwzKg95G08PIeXkt/qi2qFo
6qz041sYpZFUi0UrBs1MAkMV11gIhvPDDayijVi+dJ/WcNaeABVoX9EJpaP/hdF4
uQY42HdaVkg7tBK5Mvs+Ew8RdhlPIn3boSg48CUcKeKtePzH+IwDox4nrEFvm3cD
rOvKirrac0bxcWNvWyKPkQIIOzksW9QLE/O5ghKE70EFx15zpR9P2zzQqINzujX4
DH6bAHiBKFjwf3rmB5v86py8HFic6wnxgmgixpreOeix2Nd7I917fHiJIEvUzob4
GIv/vYza8Mm93joSZPnqs1wzn0hKj2XlYLT2TCzDT/+lBEp35ZNa0F2y1dFlloye
t3pGP7Lwnrje6LK9NNmAabKh2qpi4UGjO9/+/Qf7bEHVh+nIREUK486vRheFgWQl
R2WrW6M0OjWCzk5Fiy1vwMOAMAh0ZcUoinGfiEg/kEBBnF8nMGshW5nNCDswbPYx
qnaoSRavlEsIR9MFvdnLweXO/8KeDI1NSGXjscpR5UPTATkmBAZB8AGxH+aWus2C
FuPUt6zqu3XXPk/MbMXilGneLvSJJ+N2t/xc2em1AJttOKlWmwbvmds+94un4gXN
e6sp3eq76M1KKpw6J7iG5ZnwFPOJMZkRzunITnSjPoFTQxWJ0g0eOLgR0QOULQMu
fWwX4q2j3FF8A59SECHZm2FWIVR4i2vIrHvHdMbrrZanw//bS8jcP3XjrwgaTw3T
TYChS3wDNNm5c3W7OoEZtEwcY8GgTamMxkt2YT0GwwhqlEh6I9DMo72rMkfnF5Oy
t7Ikjvk1cSqss6VNSjLuQ/Ww7ZXjVr0y1ZnGveN+El4/5VFEHE96QVw2mM4eW7Mn
dHVpD7CZk/adSLOq5/7DRLqTk8/fJhQXTbprD4rLY/HJAkKtxghZXxKTTcjfOIuJ
rVT6DmNEwvhgPmR81Esgz2vd+7bb/eRjpgabalWux4monCfGYeOoUFJjnTVoe+zR
nUyTMhFEsDfB4aViNIfxaTV2uf0j2qjiJg1cp5DZZzRVR8+ltMM8QKIs6lCPQxRd
DqWXGwIWVCsFStyh3iglI46eW593n132o33ehKZyxxjaOmechjSHj/ligo/h8RJs
IRJSrAXhYfr1Ij/bgG+u+8XrSPve7eQPdC595DQozkHPkik/yb7kJu0z0YKDmUc4
eShQ4nziJ1i8IFJmF2EZ5HrTfzK92UTxy6R3PkWjNMmRXCdRlUE5b765ZTBkzsWt
ytSfozF/6u3hH+1tfUzfz+Et4IzxNxUhmyYZ4+eu/GLKRwU/JyfOGNdh699FZfk9
GOq9o7ETXWZIjM8RGcOcqwGctRir9M3Fsz8CisAhtAipuyDxIpWFa3eaWXT2Vrt1
xnpt8W9qjaJ8kVJJ8yVGbLfpbpRtQPAA7TjeDWtT9uKESk7eLBg1zaf/Au2FGgJJ
O/PByBDBqP5OL6kUuZCa6QdgA/jAbaGAykDunnDTROZBeT2jDc8x7L73+RjQYJpo
fUYfOfsz4yXShMvzr5+MlTwHsXgZCjOoJEQFT9M9GwbIG610OHx5PUAp1u16ClQz
zjhFRzaLe1CFyCwA5wLJvFGCgT6YpVMVsvRbYeTEB8Wivykiy6XaOevbYonfX/lg
/2RndBB5TWD0Q+r9kaC7amKvYaKcglcFPuvl/QOa1E5FcbIWAK2xEhoJUMIU/8ht
7N0k5FG5wGBFnjmp7ZBDAfZBtJT7ZiaTMGOH1YvHVSGLXfesZPosOfDyjQoOCYnu
1ykDsPd3BdnKwysGAwmZF66b9Qftj79tv8WlkjJcEWR3E3kznu3SHkw+qpTWN9i3
XXs+lzGF5HsqXWxvjWm7+gb2E3TUs2wL3L8OyR8QjylA/GKOSRJvAaOhaHQmuk0m
Z2+qNW8xNF3g7IhCG2uZk8sMiStILlufEvIbPCssSJHZQqZyM4AdhQRl1dg2ShAP
/3pOsh0W2DaRj4V/gQxRferKGpI/FCFjQvUheGEQvinGbrsjbUO40O9Xz0Z9s1I/
SuJCHTPsUzcYxDVSkLMCqqqqFBL8CQ44Br7i6AL8bw/Fq1CAhlFW1xBaNrAQ5qqU
hmJzTo1yS+M2syheP/fJm9GrAceG55utWOCwBIOCyT1K6X+khy97VWJpPwkVPeuN
nFPTnIPI4IBGjPgoxQ5fAR9h3Q6QMZuhJmA56aTLss4B5DbTjyARBOLR0bpozo7C
yhKvrsoRIrJSopApsL6Owv78tioS14YPvopUFU3f0ztbg3mQ7kxc3CNcTvmOVUXy
rCPzjkUMKcfEiSS7fIej6y8mMcPaWStensvy9fEvsHul8X77NTGckEKo8F3Bf3Fq
9jVJSJwMG8auLdkTq0Ra/a+fjcIhNrKxrgssCR5El4nzgWb+4y5bM4EIJ22Yk9NR
WtUFZMPxSTFS7y+B+B1zIrn7VuqcnwewnfYknBsY5sFjlktAe9WX3rPVIrMa1SB9
0lhq2UJRjMO/MIau7gdFTDEWFyUqGjWbqSkfD1qPfDqy5mlbW1PNZpuVxpoUJg5c
zUF+fLUYrSb6SWAhJvoHB7aaLCQLzGwLvAFf3FqaBNBft6dnoYUfHPStDAncWF7G
Xx6fpP8DgCD5uIFsVu54Os8vSMQ1IAMa9+30y1QjzMLBGSaCmS9iWoobzwEe/tTi
f/VXdeDs58FaHf+C5poOucKM3UJxB192cshnWHrkz5T3oM1j7/PWykF1ZxQv0l5j
gNfJCMMmOyDjzZTh9/YvAHQBgkNj0VmdCf8pL5afwLYj2ITslqqCCx2jnNjkK2CJ
65x/clNsK2IGd5TzhS9zC1AmpoCK3loovxufiOX+fHcSsrFlHAJrZtehT+8kSafN
lZw9cpqmVHcagqfoKH/iXDPOTkUwBrbaEw5jNYUzYNQbOzQF/UWXfYXyQTeT+3MG
JXPaUF05cauw3zC5dRd+zk8pC0z+uIIv+Sed6Kf7ZgWm77vRrIsCfVg7H9fNEJhD
oJl7CexTTGWCzL/i6Tr0WunqooqZkWlEdvhPUZOe7LaK/ne3mvhrSKiaaUp1w5VE
/CqUsAWz31opskRMItu1PZOhk/9o0WhTaVXaaFlQ2ulXOeHEqlWFat+7/dP2jg0X
ju4mIwBlfBVepeVk6Ol+L0N6AYSAPll3yYd7E4pbOVWW+e9ngvhKZ2hpSeGaRMzQ
4WEjvGzQuFtWxJ5jOfy59nPdfTsGmrw0DEJbilDO2SjvFoqtckMIahCxPCSd1CI1
/pSpleXvwiJ7EzU7SNmzv02DTQvU8Y0/CtQyjxSMq75M6nSeSZdFsumsmotWPbij
iTeuPTYpGpQl3CvZ3P1R/kxycvNYccESn/KE08F9thPQbPxDaQl3A3OUmPwS8xvY
w/V7dARJv4OEZ7fHwyCZNfn/hqHoOGo03jnQAkSjV/bxC04+4GurNaSCBy/cZ9ag
TxQkZHOeUTyetDUh/z+yIwJb2w/tWJ13KdKObI+UEZWVBTbcEcctOVGaI/xj5i6H
vWKBGk50LX6rWc4fSbjSr2/zROfosSf98fiWkuluyjffv2+m5WX4s7fmTfeTFGG+
JaPASn63sQjNdFAdxRyuDBb4J9RAkw1abKMS8hM0MHIT5EVcrdmo8wx+5OC+RWMb
yvvQ4h2HMojkBs71TxfHWbZK2CKj+SM3Aet4QDwMY7dA/hbP1gBU0PoVKM0Qth8d
jWznki0Zgkd0PwvZrSVNshe416YrEQX/hMJ7Tmkcje2sbfTZz6t9Qh7vfR87v4gH
YQcvk3nqvOBWVW0aha/H4dIhf6aIIUGEJNKHPRP4/i2kbMPMs0lelM+hhbcqX8IU
w6md0qdZrAqoH7o19YgEccGX8q3/NTO9TZzP/rhtxz1Nqvjx3cjhqZtu+hLJdtCJ
j4jDjnp7kxgVuRK6M+9ECKvTjpiuZ5LLTxMSavqBoZa9S5B9gWnhS8SDBwcJdN7Y
C5JxmAf0uwVRSXi5JTv8EMu7qIWXmieodRr1ppcIrk0MZs2xDH6JkfaxHxejVXGj
/95VI7NKPUceZdum+7YvcrFrRTcp+C6kO0K+Z0Dyzx0kGoY+rmob4w1WLZVsr6ez
/eohZCNXn0yL6nsYwvgjwkzAfBMH2muXfMSSMKMPVPfuMNCiVVDfRv4EyMmdiEGy
kvP/GloYxLcOd+BFdIWd1zthZAqZUIUUKpMhepIWsAgUhVd0vPyZKjushD+z4grR
V4uqis1kxS3G0M/dK042BxwRGBix1bkCVSKPPGesOLcGuWLMPZOlSxG6oQ99XOUS
S+vEqNnPlAl8WGsivcnrsLZh5B5nGvEymIz1N7GFK/O1FVGE44fzbPdj8GIJ/rPd
C18eFkEDvMh6T7efYB4qfCc/cjrTRH/Q+7Gfl2CaQWYgs9ymopXsw9lMgSg965K0
wy+qJOhbkgR8D67MRjMdeIi3GDsrqt8Sye135bWqXmBnCBwm9xoV8cxN7UFeHtPX
O0hh8yOmZif9JSKFLVCm6aYZmmUarCO3ilKPqisSX1LrgswrDVGgGB5Gfwn0uPHE
adlLwFAudoQdDNPNXTqoaK4VIgbwOweJK2ZBI4TUB8eEIFFFW5CJUnxpS8AW+TJo
luxblpkR0P3C9CAhgcWiaNfYoR2kj1G3fZhYHnBlDiJWbG4telHxkk9CiyBAG5NI
9dXloxC5Ut6LudQBwN4sDnQ3Cb5ZjeaqfHZmzk8hyumd04DGVfhGF/oBVVNn0zkk
MrW7rAz5o14teKTOQWkssPsDmS5LVH7P5ExY4ANYVPaj+VGhWTXoIcxin/Fjt4jM
jy9cPk96lAXt7QB0f5lI6TylPDcnwkVSAFN1AlNfpc4yL50shwmOTfCR20Bw4o+S
4OE2bypKL2Xc7PtuF5JJNo2LkItusMCv7urEwcZbX8LcS9sVZSUG9zT1IZdi476h
+C11gaWvpZn6t0/SKbHn4Iw7wCpFF3S45il5QHXGAnx+1Mt54EY/tNjzInP+Eavc
tcj03L43qQCkv6iPhOW/7VG+6anxPuMxgzsBnkhhVMhu5IyBQAOiFyputrEy7RZ5
tr7uBig0Y9IqEz4CmvbWEJhGTYkJJyv4h7yg8Tyqf+7oqbdimRFvhAPhSDgMF97J
ca1sbqT6Xhx8xqriYzf6Op9YwMolO7EVNoQJW9g5tTZu+dbz8Zt4i3/CNN7ksJdu
feWjPoFypWRjGGULnLMoJuLe9Z65FlggEHauSlh91KCHW44fd/0T16k+6xDVsB5x
xaV94M0sabwbYFeJZH7dh8V5WIWSvmkVt3zXdyt4xJ0w1/zho6mUOCiaaI3OHHKo
S3MpBkGkudjMTo40PakWyIl4jV3zTqaC49sL2La3jv4m061UVUCRFeTfFxJJUxJz
ZD5UJ+wqfC+Cg0zvAwlInayIuqWJyXebCwwA8ye8WAotEMnsTS/KjSUKqCN5Wzrb
QPogsOlJo5u23IKYAu2lEFRDcdIzgRq12ibo/gjvxGUTNINu54Sn89RT/Rr4Rk5E
buTr+9Svcxyb0fA7mqMEN/S+sTdDx4ZjuFWdAfJBb7fi+Vj0WARrFK2GRxqV/oNW
1TzOYXffmI0IkgHt+Jzhfah/hPtdbdT+pcRSSSGZB6xHRgehGeAmUk+20K7+6UZi
ZKpb8Z+msnvc36gad+0SHmByGN02OUcn+XAjMTH2j9W3HaRRAD3+aHY4Yn2VQJgC
7wakldmq+PmmS9VxRKbVzhUBRBT3anySruDGKIQTe/kLK4D+fIxqLVBHyMVfPEPD
jP29gPNW50a+Awq/IWXvZvEzb1eIaHw18ELRtn5S0IzDtttIuWAY/wBvGs71VrjQ
v6PAIHxjc+jg0riWQtFgCzw725B5aDFf7aJ7ZLS4I7ew6jJmH6O/JWf/6uODduBE
nYciIT36OapOBIW3kk9LCcMGlC50LOYkEmbXA+K3eZzEkk2F3HNDFYWrUxwhBww3
e9x+8zelFotr7ZUbeUVu56lifPWQJOUXBm1pMCm9obR9HBGMqTXHK24j+wPd/Kbw
X/YYVP26XvR0wwX/ZEWtL/2aoXkZLSXleOjMbedoj7nniywaTr8hI0nKoLiNQQZD
IlobsXp3teVtqdYPRr+HTbE+p/hMLP646KEDY1QgCNupF5ig0YNbsAEfe50HmW4J
t+yl12ihnOJIN8vIqAZOHDIpQU6p3GjAIyUDbzx0p6YubBDKIFNovD55aIw/Jofn
9QOQ6dPmHt29x5OXt88MM438ci4dEr+f3qyst7phK76McdbdRTqHEQo/WH8fJoWo
ELUqolti0fDNH6irmMrXlvr63FpRuXriUzsGB9rrY39P5btxajLqpH4YoM9JHUW+
+TibQbX8A76jr62rPFcQTj0iCX0Z3m3DC6oOM8CVuRH0LNUSwKYLsDTPPHBFHuTS
igMxrju/nxFVpov+ATzml4xjS0un/NyYm72DKh+Q0lyDovM3QMxv5FhLjLw6bDaY
/UEjxekk4IiUSuX27lxhf54CLMJHvCc7yM0S+6LrIKM+M/ZQnCJGphsKKZ3GRQ6o
nB2RC7ZNmLpsIruMoG5J2AUJj0LA8Jm7vBWYHug1uQGtZBF7z6l7RTQlYEaYVCrs
0TMhdpdF+VJO3e6Ala0SV9x4ZSp0ObkHaWXRa/w0x1jP7Q+PN7uWoh8Y8baBAvvc
ZulO8GT2wc0XWMinPdoYzvIFnaC9yWKpoRr/GELCYzDhyBZSLLpDvjK5MHC2Ixmd
em01oZiNwWgfa6jfyNtvB1H0hamagpB7dkB6xPB5BmlrgzcwyhEULnEMUO7nnNuu
KNXrCrZHcW5QFq4jTt0pv5vi02Rj4BadZ7jumKh7/i1f/cv3CgJcogDG0zdf7FnF
+NI4CmuukccPumWTtVKwD+opNLwgFbzf25rc/LQQ550CuUbfZmA7+IKTPZtgVedY
6UVVa/fDRWdAINRBCqGSD/h22mz98y1mPAhy4b4YWGMWIzc8t+M010NfWuIXLgjS
q9B4I1R1ktf3lkgKAdIDYS3LDfoHEkA1XTMicwVcX7ql3nYEFOR32Vb8R3sKbefd
jN25atUaBrisV7nBkY0oXRLNOcl3H/LlWTKaHcBg/0hjYv/Vh3Bxb4ijsOS4NY9l
fyVWJk5UMf77iGaZpjNiK8pYHHWFPAP+/uAbOgOwA7lq4brs1nlW0Xc1gK6k9wYR
WTgB/HKHkP7LYmvc8l+b/mKC6PM99BiZRZMpGUj6rhSIoBFny6scbgo14zHZtmKI
HCxcXsRk+eE3JTqdk4qBf7GILZmoDtqtuTGpw/CMhxwRCKILglfIhWGX4wDs16Qu
LeyJ2AM1/1Q968nlhlu/zltLBe5c4rc4gLdWx4x6zFWHzHrzPSpvaBFnnS6Tpm4x
6ghyoYnz9m8tPPaj64rQ4zEOQf6fTojesn/s909EFy7S5cahI0zitR71pCW+08Er
iUS8LoDGd8W1li6zrbTwVaDi1Bl25AQMVMnluFcI/8+Kk9hX5AFE6AJTbrCaM3jR
B+9wRQomvj619W391WnDFnpcmZXahXPXVgXOzF8GsLzW5SCCFpIh0Yty97b8duSZ
y35syyT2rYPFVBFzwYcfgPKOdgQ2KGYEoZuwGrxBZOKdD05OLBBYWtYTmMgviLXD
0jvzEkSv+JsNJyO0DQ+riTQVPlTHWtQj+rVhMDJDaJ1it2sXzp2zbQy3GSfdlpaJ
jLkB++ShmiejJo+fhGTX0sCZiBNhAw4IiObraF1Lnt1gocD608HLbtq+z3TPFXeN
fznzvBNadikvEZyP7igvBsq1LDY8JzhHWUjxtleT4sDU13UIwMd3JZERRHjg1rWF
NLh9nMbOTwULGYpFcrzBGeHaXvpJXwoVGZdG4KEfUYioDpcdTTCmxXqSzaR4F0Be
57O+0tZKnu9dbofsDy8qxfuQcBizfWjceCtOs3+LzL8xZ8QGXmF4yTc27KSe1Yl3
GGnXM/c2PzM7L+L6pbCMVhzalYEM90LeLhAtSNVOlLQ31V0jjoyWyyG1aGWB9zvZ
FSfoK/9sbQNECk+h2qTbb5f/nqJyu7UhMDClMfMJ8n6TOsGiXJyr+mh6Kl1uy3Jm
vf+aWdiz+fQP7hB7Piu4X90NgCCNMNP7294ABAAmb9LBZ+m6ZDSoKIZVq7pPQgKB
fsHFlgnUOd6bYCLxEx8R+wg1liS/2HbnNE0srrCe8TxHrTDJpJCHqQ//i9iS3DNK
/60F3Wklg2NhwNSUNiCF5EtJ1XDJvCLoPTsu2SMal3QvtAAvq9NFtGGLclwHu2dH
HCMG9+coOs+qR38mHUrHJSTBQjK/WNfgwTt3eruDwC+tm1HeBb4u1r2qjTSxhFKx
QvMNWb+PfW2IhL6YXs39iDyIFdmHKOBicsEOKSyF98UOxvpM5dMdyUKhjuxxjshj
UxMQbUdBzhDET5EwUKFkT+wQ5AAq7iCQ37dJkcKmWW3vZ/zrUadCm59rwSZL/Wck
MIuTmi5daLXukic8WLYBKLOlwmQa2TtpXK5ZqEE82+9REE1EsYKQI+593zT2kqmH
5EMaP9OEjSbUyEe1Yu0/L3J7H/tVSp9STj1E9WsBwJjJYES3nJYb/oVi/kfb9x8m
binl3zTsLoEk4GMLlPxgwPjtcJ317/0peKspnr/U1s8iPQJCnZLQOljLEuncG2on
vVLZaPF+e2gOiu9hNYgB/43TJS2LUZMVvk9CjKVTkZWbqgZXSjoKwVmR5QbOtP0s
v3QBGF9DN4SE7P8Nu3DGVrTDDMcXegctCp7LDAvtQJNRgNqsqOCvI67Vt8eL7hs7
Y5z/IjpOEbw9JgPVz46/jSWQ75GqqTPQCBOX/0cC4rFhgqUEgV1nS70lJbKbZGwN
RLoQPuStOY7prM+BfmeBzYrEiz45Wu1M5FD5dEUoVAh/mnMN3C+HojYJdFXPWXKe
m16PaRigEBdkJbyHtHJ8EEx/YG57R/ewc9KNF1nCVqlOfvdsseZOrZFF8yv/11I9
yAKzef2WxrgEgXjmTzowNy/RhG947CFk5iMEQSs2FMa2CoJ+HQP42N413SXw8Eh/
0ZGO3mHoeSUnMvJZwJY8oCZPLSroxVmhmtSc9vSp/dPwYxctyjpOp7zh+AYJUP9c
8v0xL6v9pZTzn9V7BieWy4x6THRn/9UdtJM7/A5RgL0MUoetjW5VW/yEXeDZLozO
gVScDgDXYtCpjdIGYeswcpVYcaQY958Sfoqnmgp+E8uMRtv5yPdLajM+W8vtgrbM
BGg/VX+plEP36YEnJbIFdKuCyN1ofn1kAOSozk4gHgRtNclv+ZS/alQaeuAMJJgc
PBtxVRaZ+QIBjDCUO5k5zjGkJK1WD/WzeJYY0WXDM7jx5ayQka4y5ngfHIpewfdz
VdkFCfJhZJYbwZKenCeFGcHrsGnfb9xZpMYHGruYPrU6as6bUDcyfg5P0KxG3SeU
z9uf5JbNL6ygXHXBOk/02eQEPlqwqHvXkGmRTJP3U4iPy/ry+N9lq167u5+4e0Iy
B4HipvQKC6LH3ovCwjSxbAmtjusklRG/PUV5eKaKrqarb+2usotLbuSHD+3741mR
Kh7xP3hyuqX7MLm2yYh2maeq6yOlYzGUAR2F1C81pIMNaw3cJIUtf7tLraZsz+mx
I4iwvwFhoqZPrZ6LYHWBXevonODDwHeo7o0f87sPAtpFdJSLwphhqSh1SFVSr1G5
bMeOzBgjtAcm66XrEjnCPBb10P5TCwULDtd/D9NZuvh6QCv2ioNtwi+XXeZSNPq8
DI+BUZb5ih/HW8Vhfs4twe7GOWlgEOLui01iP8jHL4/ws82v76NTEU3oocPW04Ln
TbNf7VrTzIm5fEsxV/PzIpICunLDU5nu3r01ixGSC7d5kp6qM8FtbFuSb2+xWyiU
W2z93KrvLkT3bKDEGdyTiYg67ZE1dmM/jJzrmG/6pwWOnEB/D6iax0rdJMpgtEzw
SAN5m86pgXMdDaGIKiLNbaCl/4dwP4Pbln/77IgIDy1Slzur40rM8eH3pIwMDzTZ
KdRgITK60s8tAv4PeVO9uwD7siWuGfjqAC5PYz8RHFBUThgSAP8UEZjfC5ycxz26
JZjCes5Ceqjobv+3oYuEg2xpBOATKMirxl8BWV+fLNb8gP3Oss55UfKQOZ1bq2Tz
fiMtll7tXpoL1f2+RfPtTOflK//NRUvWNWUYhtKTVJpUCCvy+G1wkjuk09Gdc2GI
xFPbCWZd9rRscs+ndKOS9+0wUZWHh5rnXdpLpmIR0NSnnZmFZHPX6KDr8v+Qvi1z
ixaeweWt5ZQIP3BLHQQdqAo7NHr0x9bTcTqmnLOiwMJ82F9cJsI6c78Zy/szRVKU
KqV7eJB0bN9Ts4MQG2EoEcCHpKapqNapCE9h7NGxpvoHvyW4+Pnmm038mVzo5c1S
27l6+bZBypdL+F/hBypLTjtiyRgZb4kzIe/lGRNATWHAT4iZYg45o9ex5sZJ2kOF
vGOJkIdD8xtycrGJqn5vLq8vCarlAGvBfRWW22wISF5sVAT3RzaYAfpQX+0nqI86
ptZBbSKyeQ/xtHYsur7WzKhidQn/tqDuwjgIDDk20Qf2gYF2msdZ2Hogi9tc2jXr
yZ4G40ChjWtrrVmBZRFZ46u2tkn/Vn1Xkcywiss9+iUmKVKuJvAwJl/gMP/h7avs
zUf8X4unrKmn5nqeUsO8rzLKvb8APHfAt4fetFEZ7y2qQrosXorjSId3XDIVJYZ1
Ms0Zc8K0NFOAvgd8DocyyAfB/stCa/WJpAn3PPz5oia3DiNXyTPlV9E1ses3wOhq
3EFzZqiKIH3d9PPgEW9ZI18FA9E96r7nq6EX/skEiIDIPqNQXRzSwL2DvAgZjHgQ
S9ZR6NKDmjaSGgLc/IyS0kuLpEBj3OXUyknxrSXEMiov27qrlsVri3RSpFbnU60b
AgdAHhFmWK6kdtzzhBsmIE2jNZaXl3avr1+pyGR2O9BFvV7IugNZ9LtXgP0kSTDM
Wz8vBbbFCcCcihfUbCE504mX7CeH+aZMZvibKoA97e5AuK5eMUzVZ1eNM/Yvboyx
pwPytcPPZHxYmtPmN+rPMMCJ1AzfujuXbqXrX2qprQZ9LTVoodFChRt3NlvVsxsd
UIkcZYDwtgjL8MmS56hJyXjuZ6CZvs/4WNNpUDjbfq3FGAkVks3t8272DFpYrEhX
FyBZQmOY7QcyfeCP1bkANz88VkjGelCNTXUsHNRAk4jFys++Hg+cATKaApGg4isx
mnq7A8ECPVUw7jxp4keKaB+5/z8KrBSM1VHDXpWiGpDAypA2zx78qhaCzOML4rWA
zcM5dgd9xGf4Bwc43G9AiFs7mUyJImYRv27RapeLSnTvjPLr7RpFU05gxuB2pSvY
ATq1TOzIggtdMVjXTZlAlB9IRsoJ3jnbh5NDZhLFp/TeuYLOBhA85aHvvIRPo2m3
uLbosH0vFTTd6HwsBWgLpeIMx93Ut6SHXXJk1pHC+7lQTgszUqQ2ePTPU/ksfWEa
IlpWjEXxfGNkbhS1ieUuUyo3aP/hrrrlNko54q9r3OwK6nf55ar9i3TTNWBpzWeu
Kqk3h4MrILLH03VH+nQEFmWycqfA/i/SGm+43O6yVeajiDEDwjKkM55ehSL7HsOB
IxJIbOj9sbrjP3vN3X/sKX2sbOB/zWdsrv96MdNUnAeMawkU3k5RMsFZyBzy1+Uu
VBwfFGQDfbbpvhnzdDMFOUwPLjXcAAV+DgYpQLnqyApplnXY0ElioIXVRI+ic7xf
ndq8y9Kwdv5Zw5uBhTTApSyihK+kRky7OW0cWNcsczVA2MYtvvxGt3hJvF/lPsKr
u2lFBzuAzwOG85b21OaPjn8gbrWc6BdVLbsqckY8plPHk2XWVHGW9I/U5mNySfaC
CZoOdFEgWN5HwPN9eMAoKtoEjPDsxXy6GvjjhLu1Rzreq5XG3Yhln67ogF5Cjlrj
M5mqqgNOpINpKyIlfLTALYQYIRjTK/v18sytx2/4+yR1CZI+mzJ5EpJPWvFJaePO
k2VTAi4xVIabyGPl1pcA0yQ8LX9MxhqvO/TWMhy+WstRmS6l2mcXaSeydjGWYDZb
A8l6lA5UtVzAipboOAtmPxMPLvRtBPSuG0/+DWT8NKsJXGlg9SQjiYDKrn+OyrbV
NoE6Z2tvdgP5PSMOMg30Wl5fDSfxRggupqYmI030iBwLW2Om45+YUkVnafjkQxVS
Cfx+ArI/W+A/bpPeJYWOjb3TOMQIxRFrmVbK6Rdk17pPg+AsRpXAp9+X0flBrQ0Q
0V4aLSvdLcoXDA6IpvNjUughDdkdLFpUmozBm6ukCEfeB8rd/2Z/mg7PyDZ9hoPY
04nvtK+uJglt/maV1DqwBP7nfCXFjd3dMYrE5s68cXkVAsO414IsIahQZ9erCcx1
6JwXIi8pRSE8k9aDQSxx+ljnmf1hwY2LDJpdxJ00xvllBfhWsY4/6CQw4c/BP7ke
kai/uyKJyCzg4GQtpN9DgBJIG2MuK4RXBLfptc30ChniiZ7loo3U2RW3WNElLrpx
5io+xh8TA7PWDv1+KsT+UZ6We2BvUkn+o31xMz7ZV+q7cqjYiibkOACmChbsPpmz
FnxSOUJQrQUldTJ+dHDkvXoQEAcaribvaRLIMMXbj7bBRSfUivYT3ToGGx8tL8wv
qzjuRK7jUwltO7a2qyF40ytqgHLj93VUnu2b8QK4G+gMN7GbtnNDPKkQT0Q05ECZ
wmkavPbCKz0uxMZFqGfp3Lbc6uhCv/q0NRCHYgCIL6DWZZw7XCII+V5QBDkgIIab
mFmSFDWr2MEkeFYHdXEMH++16WQLZl31tlGbyuqq8V/2EQ5YnuhvLPYS68WeGy+T
LVAMBLWJr71wH1WzrM4mIIcHnxddfBSso6qXFJt6PoErzC1403esQvZdqwRByzuV
kdLdsRNGQhFv4K5eiBGpQfg1EuzJYSNyia6jqjV2dm9e9yurJgNOwHStDr40xAfn
S7zAWyx0y6avpwHv0lGAAwLydJODUOwiJFs7Hcb7MAmzHQdQU2g4d5Q8KNFmcVDg
bpVaEy0R2vezezib0Ap30UUQUxmorCXFQfjVQkNPU4pI9ysPB9PBrOoNFdEcypPm
qTVpVcbzM1f2mFRD4M3AlvbvOAIiKDu8VAnxcuuuubnMENCpscfJ8ywV800MfWVQ
pkXwfCajqWQSaUaqjzyVQ7yTZ87PyFRXZzU6wQOduh3KG6F1zZpPGL5MCDq2NKyw
/o1f6+GE8CSM/ky23QI435ti5/VWCVNU+7MVfYz2DlZFauTTK/xK/WiFQYJKepWU
QjLNJoX2gl3KMgr1sm1eNY+D/4jPOVwSq0Dj+5d/+xtKVduJQwbgOTzH5bpTKJRt
a+D03P4N+3altDP40/R6UaVWR8SHuToMFlZDv96Qi7eNZCW/SZuw24OBZ84xNu2Y
BEPw5fT3jqO3TapQgPA3/5oR3NfCoJfFAUKCobUIM247PlYUC4wjxgbK5YEUsqwN
9LD/VvV5J1uSILNJHygrFLdbSyYI0krsiKbAiB3gnnq3awhYSjj2jxMcXWddabWr
tCxG9RV01Ak2m9qgfFOZJJxvCPalsZav7K07kuVdBM1TjlP5UsCRnsvsltEh25Uw
wiyhxWFw7oCB3j7vma9aYiV8VFpfpeu7cu7YGZ4j5gWUOyUkc8ocjufHcsSayFRs
6BRelCqowAVpGnb1YsQ9uvtoUyzQ2VXwfM8v3qmOU2UXygjyU4nm4GRrfv/4Rp34
5IjX6rCC50qgpH0zzLQ2t1ipQ0fEQHSsvleSu8kKEgXcxnC7PngoHVD5qiDW2+8X
ozIOiZYVlyaXi6kjcEArryjRhm9J+C4wqzuzkLgwFpKl5eE0zpNAZzxn/jKqU110
P/QM2D2wytz81Jfnx+FbpdNchqQKCuTKhvgTFJ2mkyrwUQwl3vjUVQzbYbwDvSq+
7GI7sMlyB2jxz3n6+ZhwtljmDqf272mmuCGJno09fdugXBlmF710sjbMWHoN+mUB
lj7MIfS3aBhhXaSRrJAMrsn8FlKa6m5Hf4N+YpviN9wuNWhEAxyokhYy+IEqX/dZ
2YBI/GRyMu3sBM6zr6Y/yDZRrjhnOZ2UoktvINJxQhLNM8lQAhpvERMG4dm42YTR
3yrcpDnl2mAIJf45Lm9MWDR/e1IqjSROipbfGGOZxLd0O4rlJkXIGci1mId8vOuN
mdh8HgQ6bYwMUJ/Lulnj1wxCbIVBojNQbDuHuIhik69Wf3eUKXHjg5dDlfs5cMkq
8vGEFEiJbO5wBPpC8BXdJDGhdMajFVP74W/O99B79FO3kIHsXmyAlrv5+8Irvt7h
4MYxkBOs+pguVS1ftH0//1TgdDjlb5G4jkYHRbV5FIGIaSt7jAAl9dXEZvnUlEeQ
kPzIHcbZ5BzSs9PrFU8/OrWoqaDpHQfzbRsLtCVWB+j1sz1HeUeHcFSmYNQw5Lf/
8EOGLlGzFshX4fc4cRWz7P/fqVtVeBJ/YhbzZHxa5HxA27IMJUI5gQnLEjYa+IYv
iZ177KFT9uu6BguFi9gIpzpjkgXQy4p5VjJWmAvCcy9pbaI9ID10sXB/RNxWAYV2
KLI0ECSEnxmWIkEPepcA8cFzVSgsPIbZ5X7hrjkitv0G52kLuUDjkRpY76GYAUo2
8+lrt8sNMe21mL163whAaXgKCoSMOZmiOJgNlK/yBHgezK5T3nEZjF3ORPNr+dnH
KUY0ddyVJr3CbzCCCbxs0+NWb0M7W/YmSw8V6rmVUIxiun4g9X+sBxRnvs6X3lNl
QLwD1lWbywR6xiHCQrmO5CA17lRPfIRYptvI8Nzq18h21V379UFqjWLOWtIFQ5Qc
94p6rHZ/dsiCGFtG3jEkVjnbVT2gSLVW9Qai6Wh1BxqY2Yw0xpRPLc9aoOvBnYl6
AwTzx959YtpB7ULFuLT4Ql4KnCJOkBIlJaJg0oaGPV+u6P2SIR1bmqbGIpEO+4eO
BiK/gs7f+qfyIVBZqm8VEZ6d0Ydx/4p5PLUZ48fjXqxGmuGy1PiSR+KVXMhYkRpG
qb88RJRqOd0+HiYmlMLZCZb1b6PxuhsbOypSusnnNNe1yXgsX5lEWDyly9Ixz7IZ
VvfFPhoAGNuellDdixgNNm29UidCplbYI9YnFfwwYA3+kA/gg0L5LUhawpsdGcul
LLmLySt/QeMB48tszRtcCPSkCSU5KkKP6KbL24ESAc+Az1pjA0DG4yhulBX+PWkm
vXlVkZ48JKIjsjtcc6V9bMYOW5N/eb6lot8agxd/p1DJhsDyfbHSKHne0ktrww3O
vfCUo3bBiKw0e1bDMKxyLSv3LP3zgHUwwEzPYr1Pf2qjE9RCi9Uwx8KlsUnOf9hB
m6lMpO1bUFA45YuLaA4eRMFwqS4OucEG8+xrh9J7nYUZjvhi0TvgQbu0xv/mJS6g
XIaF/HxSuQ/SREpa1SPIVyPZ2xRY1EIhZuwuhhA2Q+B6uOa4rNk3OYUSrKDCnRh1
EuC7OL45JIgBOdOVjAtgsE0D5ETG13NkTgrLqwfMyYfBR0TNTopz6iYZ0CLvVjV4
rHEYVXlRwHh5Uq4yddSob0H+9o9PLfFvaUBc8+8iiKT88pxBGjk3DuQPyOVwiiO8
IIHVF1oLS+1Ut85PT/xmpQZfXMVRMwrSy5KAkZLc8XASbEmhfWih7dFL0AzykLhX
abBuULEdnraetyY6nJlAHgrqDwCw7Wb7FPXzR8wqzydf7854XT21lxnFaQ2olGrY
zz6yx0hVQ0IoEs+1MWRGC8LoaHFkW7+iKL3eQlPxBzN8BvptLjwy2K8Q2973KtQx
X6bc/PouElPz5INYsF4lXnJF6ZHO+Okcw6xFwI46NpT8gumKb0H1SHmJ1BtyQiCZ
a07qkD+z00Is3+v9XTtcCaebj9oVxrdwsK+A4f6JqhHmLBoGoQFeJEYjk3VE7aEh
y0uHLzWwso4raTz5Xt8bE1ZFQXx0yqiE1QEnMImiWm6UiYgLs/8cmgzyUixYjvgG
ncJsv03BrclQ3VZUewq6KCF/1b9uu/mtzf9ulUx0PUmUX0owhRluI3icP8Pk+cJF
jZw8mK2015tQIt86sXH7cx6aIakDANYJgAKtoPjynkLzssT6kPEmOk9SfxIw7wbV
tLVJ2xHYXun0Yqa6OAUZtDdxDzrzgkyo79jdeMZcE4dy284SPc46T05KJDygPwUH
Ck7c0zj+ecC+ioYvT9IeEqPobbpC8Ya7YFpaX7OpD2F45VfyHOPefn3m6NRea39z
6aKIUa1Vd3jn9Aqg12K+RfaLcTFovmo6NcmaqVzbtJyhSBOpaNS1btttpH9B5KS7
Rp+sCAynjYeH9es70VJ0S8n+zlBrfDUJ4XvJefy2QtWy/4P5gISYdgb7r5O99vdA
7Y/n3jHnjcBx+Hn594pSNfahxPcT6yo7SHgFwQD3LKuatdvFPFnfhMSs0DAltvLz
W077pYlPHcGYpXO2i3k3iSdut2imJXwxvXTbxaXWLmTVt8eQ1ySc8o1Jv7O/dQH9
2E+ELoLCmZKsYCk6Pb7T74aXSjV5Suml3WWZbgINeDGThrtjMxDWsg3zyBqOP8u8
zMzLlbmcEFW1zPeswYFy0ctcvUL7DEyOYk6qSRyysc+vDcFJgPkHT9BlEtr5obLf
hZ7kWXORnB1/Re5rEJCEXg2jLq2rcoOOzOeP/oERrwTo6q+SzQMKYTpOim6LjVEt
QWxc/VAYo8DAUK/x29Q4N7gRcUo3OSiPaNHCNSVwME2VwWbb4r8x2OTbE4iYteUP
XWs7hLy5RXdniYaTRkbELb3TTPJgRb7+tzksxi4s0sfMVtwzM9a32qha+s/Ofdqd
KEx7EHNwylGdf5P0vOdMGJZuWaJtJE259Q6H+kwaoukwB8O9pO6A+nHI12BbVHoQ
LIM6RTRR/QRpMWtEGXIMNhkrD2V0tAs16KMTaLJinhdAtFGn5ogeocdpjTxBeD1/
2Fo/FuJorIgTdKHSslKuSgFqdrx+OQis1BGe8R1WrNuHVwsttaxG7dXAYCcqBlmU
hyVbYUii8q24jU22xKLX28tU13dkUeBVw47P8jGZ8k9naZ16l9CMREKw3qfZLMte
C97cO6Two/P8wED02PiB03LcJ4/MvB/ZJCED0XkN/98YmgZDQWc01XnTdZy2D04F
U81KNiBisHm06D5ylsQbooeaHkpmnG5/TWCV8jpcfVaTJFpSMmi87RmweHtdt+zr
gGV+QaTlpzL+l42cIGFSPeZcUfIlCZYQWBqSfKH4oL6FZFV3A9SX33JjH1MNCz5S
CT3rZnffmgCi/r58mD9rsX0GW+iA1eLfTLv18O6XSmh1WOrrLermbrceUlrTWkF7
GlHgeDAi1/KwJpGPz6Jmcz3KO3s0QMVwwXPgHE10ojoTS5YTVPxhtrFKsOsi5Nak
2WGMKpEYJQZGV340qtCCnjBlUpWWsXifvOZDeqybno8blf2Oj9DqBQyRV4HTyBfZ
PCG9xOuomCbF/6JG+KON+jrVTj/7eNJ0tAvTsTptGeZu0N2sKAA0kiGw+rQk3Yf1
CJIw+M4OuMsKU4GDIcKX6LzMWJgcEKDP+RHM5wJ9JkNxTZtS6Nlf0v6SaWZeHo16
nDZcYGU1JwIMbq10kAH7vXdfDU5prJinZQy7n1AQ5FHcofaBHH+rEqpe/qVc17lj
UZHFG+Jq0lPi30NcrnriFZWT1fEn+TRIJcHQCPyf8ER9jDofaVV68oQPYdDRaIm5
rqCo5VQJkPE9Z1tSQy9ipQpFUkaKX7lRv9qhn6ddMVmr9GRIFv0mS8RJVzQ0MY8W
TIz+rmdlclWkrazgc5axcN00lxhaDbsRAZCEd1SHA/vqqOsYm4HlAqPcr4qNQURk
E6hlX57FByRpSnG+6ggLt/ncN8vG3Bgf+/HKCChpLQFBmOkVEO386HLk2Tqj95c6
PrKquG5GjBibZbAvynprFAD4jLAMrqcCq9AIgKZBP5kMXgi5PLhkl0ken77iaa9r
iLWh/Wg0EEV+iadkjDxej1wc9vxM1Lcr3U4dHMjxOvqhW1pW5ME6BfW1JZ3RBtiv
dJtp+ODfUUz2QEmBxrkuFJRheu8QDLqC2KKPpp6QUYofYmZyvIM5m6KVkJw6Qw4D
GXAY6rSiYN+AJ+U+xy5kyCRZ/be/NN3Z2veMWxwYD+vrx+eK9aXPcPm+JGvz0uLI
Kaias7NoXnSRUk1X3RA061Xq8dYIITggbIO6gbVMTmmOWNhBAdfy1lOY4nt/CzEc
OccPdK94XKvbtbJKRm/cC8nLCaLqtW7hqwmi6JyMQO7xX2utyqJToqdj831GI7NW
iFXB8zgOR8opdj31oNkdkgI4vVrecZTcjWyaSIlTOPyKNvTQSkVULqKi+6r2LmOk
50XCFLN4PJb2n2omo2XWMqXdQ5eqUsY4BzUxdvGBbRBVIbR8kC3O6650dhroDsVO
GpdZ+DJTFPHdfnCQSD1mqwfT8GeZHAOeFynPdnclVnBnPXSrsWfgCeGzwoRdv5bQ
O+p/655wO9aXOLS2AeHEDyiD2qhOfwIkBBvhGnyqwetA4Ruj/wI1Sax2OR0r3aNr
FXiclF3ekTefgVBX4Pi6AWZebrVxS4JlezUYJ1hVcEbzToTrjpzhhsr16xTYp6wQ
tWKEFnFhrvAlb5hV2atx89DFkZopErKHERC49Mtw68Enj/F2eqkilHoWPMVjjADl
LlMxy6PkElaFxJLb99rOABgBzp5+3ydOyOAo76ZzBE9YZQn5aiume4Fy0xZnaI9Y
c+BpRpz2EkSzkOOHyJfR14crLT6CnvbCf5HWuyR+qkrO1dVXBH51viXBXHXi20qL
4OdmUJGJZsRes+T3L7LBTtUm7GPGmgP/dEE3yXOdOwMmXKF1lixxyGRSsfYZyFIg
ljsNE8EOUF2BKQ0haKwqGktoXpgAuh58qDbBKm5z23nDMJPr/P86nykuNEdqvH2l
ni2xkvUCc3tn+0X0MNQCxp+kUUaWtMEkmNFnOviJIIMjoYNccG/ofMunhwEFjqoB
/60e4+u4Ms52oeApjjYs7aeUI5v2hKP9ODH6Z/X1T9sQXFbeNV/78ksoGpOurkKM
dz8+/k6qkpQ6mSrwENVxKoOM5tKr/4pYsGs01qMmEx/BDJDKaqcfDxOE5eJuXsWq
nEa2cwVu2xRtJ3cH2VxGQGJ8L7NjvuWmsnkondj3WC+J8xLQ+pOdyb3UTC24Y8y1
BUL50hvoe5VHqCUvy/Nbl0UKnU/qA7Al8RDJgH78etC6mNmkt251wSny86yQw7nv
w5hLZk59qeRGpM8izjpBTufnIkY20yKWhs02H6WyEV4GmJXyW9oI/miLK1PAaWvD
TeynV5vrAkjZvnJbpPYeZ2DT5XwPC/EYpwrgUzUKg1pKhxAMmhK1mlpwtVnfhx8L
B/07CcHZ79N+vfZeinazGlV2/heL+QgG0iBkRn0tR/IhpEaB2UPK7La2Bl9MnZ4N
eymRIKH9rmbpGqqR5v9JI74o8w0R4WlRlQQDMNIaW+URqCj7E9hXVV/fqMELjLFf
G2p5dJBf8ad8bOzmYayP5dXE7+isIX7PVPzzHWvc9m6MqH1iH2yrDF08YmL3g3SL
pp2sqhydWI54tWiYbXuIIA6cXUTEIwAtIoeAI6CSKeHEnYTMdeeGjcN4ApclRS8q
Ih3wY6Kllvj+y1KPLjup6mfMO6K7FgToIKeSxmeE0xApwzURi/8IvaTpqTUhabS2
XD8IzbD3YwA5NXoxQ6bJDj95nEouH/x/++LStZxVQOSYKtkc7HiTPJ6IKbgH4YiU
IhympUFYUUfX/4exIV/NSf1T5dYNn+xG8mUsT/PLzPYpEF1fAk+PCDJXsmyWgNhe
B+nrh/LSFwze87B1BJdBNSBi8T/gB3PKoxbq8wSlBLLPecEJ/02Q1lY5cBudi6fU
gWCGfCO/oHn7hFj0JjsYUzKNw3McD+Ez5uCgZsAfB7NZpumb08UhPQMt+yZYWFBS
QFs1hVApXRyacCmyK5BORmVkJx3WNwT0mFeam2rz5vU2qfDdbxaHhrvJCWsobZ4j
/TrzDICeGotGqNd25EaVsdCFMyFRNi3X6x7Anc6DLOIjBADVzfiQPW/pIh8TGSPZ
Quyr8rO/RvyCcAwLqt65cDJgDec7gQS4TXf3nSahfZ3DKfyBsYhkdJhLFsCS7+DT
XSLekn00I18WnUU1ElRuerzZtynwl1G26QHIWZMzTcqLAd+H/ehcHa9LaQOhWs0m
0mi20mt2bCEOE89drzuLVwhelROPobBbRCyptjgxWTSK6PF+M9FU8e/IVqcYj3uR
g88VIGHfktQonDmL0zK70sbljx+LSpVqfbMPKthQEAETSYR2MeEW90NKThUa6YhX
THXOriF6k0uo+HVbjU/QkICWrRDGLtWGmhT8pD7f93wJpRQbmdZm92RKgpJ2mdXc
ZbNN0QUypctAK5bSKCuZj0djrEzVRj/Q2W+QUqR4jVuKIhA216SDJF0Nh5LemHjB
vXRbT6PJeetYocgMBv/uV1/fPzA5Ol8HOt+LtuD1/hkoIy8ZaF+12V0YWX+Igu7n
T49Z73bTJlHDKZd1VYGuGICqy+UOODZCzOP+Y0+BONA8HYQRr52TXyiVTq+cblh3
YXmh8DQlDpWdnFCm1VtvD2hN6qy28F48KVLt/Yalm3xhWUpbBJV9z4Tul0JkHeLC
OXmuZMDZiy76DMLkXjf6yFXgpCBagB76KdYCOqek+m+z99zNqo+c4M8Rh2UFD0Eb
/c9bPBja2fEV4yOeF94ixdIRqox0KFw/wElO+L2CNGqeF/17pIUxqmPmXb4QPLHW
Hb4c2rRYz6sTerzQZyg1rGixAg85OjoqgDZwgcgEMxevz6IS3xbxCpUZmRK9y48q
OSST/4B/ut+/yzgbhoqiQFlT6U1xrqYtGafAwztxYzjexr3hLOfPovG/W5NottEg
h37pnpw5OzFqn1+pBEWXcKcJWRCjSjTWmWmQrEsXyXKys36zb88l18HIR9VatKAr
djadeupmo3faXD9bsOkbCkCQL0cg0p6cYWtePu+uESTvOn2GQzxdTRHdsm8krFOq
UEBunBZQ1vtfMiHUplMDjbx2qZgKGrrvhqCLhLWIxS18ZDHbvKNlh0wprsSVyVZD
jqFcvhBQxLFeiqNx6nj0iB1slSq1rVpRuITMevpP3sSujNYiVbJlbVhPV2hi2Pw8
emhMByyEiO9TN8EMaavslDV9WXoIN1rjMzIei0NMK2NzYZeXJwbw4Jaf5pe1M4kV
kCVBgHU+83DO5vHqcRQU4rwIm02omMjvqsfnHRvJmkZSx0J3GNh+w+Q7D/kGgMt1
vK0AHCXGnogIG2dj8GrhF+nRXdo/16y46sM0j4eUAnFuTeBnS0Kv2w0fTgSKkCq3
cVQcyeHdeBRGMlAZ+ZHzNKkCSZqOlUvA64wIEbrDvJOc5Vfn9NBhYfCXqQk53r3a
dv3ZBX76UODjdKMfE3iYFtWgnED+q2h1TvXTKELLCFDQElC/qGnZmpMp9amwbH0b
zlqGUJnl84sfnEu1xyxp8nKaI1CKcNtYVAnXRIas6ZSsDMZFY/8BpNWBBgr0yx7z
tE08wATvYp21eu+gZLQjnfx3+tnfIbZodr7WD4m+V6aOoBsAbhzq8sGM+Ao8Wb5q
7T9axFsGKSm1c+d76ZxWxH9ctrESJ8MCms2pyP+H6GHmJ3Khggbjqr8aoPplvZLD
8L+/VEnRChW6TE/yUF2BQxrI31BMjaK4Ms5ZdorumOgj0tYQsUURU2J19DOyTTBz
PKZjyA25pWrHOIuu6iLnexUCyW6At/lMo4Y4vKYtgZYQbJfQjPD9CEa0kW5zchTn
WoaTxHBZSXt7s1XyTzQ+IT3gHMlkdmNALlffIsWOYjXo48Ovd6rfO9Z1nTr0X1Gx
sEBuj+9qtGkGQKBjj3QvkNH3Q3/OXRnckWhl1y2WGlgGuf7vsWCltR1XaaWXpSR6
si+Nxpmae7kBq2IaoUCWE2CQZcB9KgCv188UqNhgizpIVOg0UpRo27RfVucx1+sm
uK0gOZQxxSHJoAkUrUEbpI4uEMw/xPrImv2dMnheAV6D0CGQzSd+bsbHwB2zVmBu
E7zVNGcBb1kf+PYvFYJvPk0EvLKC8kzRrmIVdEL0HCbYCiknGK5/BZb+2I7nJ9E/
qWDwVCp2euUzLmy1QkdrJwnmWHgdlpra9WuwRsFLQa/YabKSaWM7ZdkaMtTu/q35
LHVsgj86Z/vfn849rCzzlPRk0wCHLFXSAvSjJ1pWiHyfDohCywywmvRo6dqYc5qR
zdslIijdNGbWa91uZaYvTFCq49SGeNCDCT1JleQND8AbCQKGdv3TELog5c7m4bKG
coCAFRx0f6dbn4q0wpAmnnkmjUSX+FbIqfwNggrnB/eEKUGkrVggwFOwxPRGPhnL
Fz3tkhU91rzB22tY21sRs4cy/gB3ircEaxUKU+6im9NaYqHLyTLTHu6MiglXR9rj
vhdgmWghALwKCIX89vpqrX9sG5uDcv96luKW7N/4K27at/HPWsWRA56hYnq3ZDKW
sXe1/6QdZuPQBM8KIgF6qiR9Ng2nANao5pH7t46c0Y6G3a/2W/CDKQn8JrJQLPbk
tXC3E4wUmJps60yOwYNYESUacnAAQv9JSCeUvUMgDfhxQuuVar0ulzh9kxrdw1y1
mtVmSD3YB30D12IlTXyx7L/CK4+btr+nI0nNt6KpHlQ/QAanmf8pu0DwYssWYinH
BFUVPbQcDNwKoK0qcWw2lNAMDb2QExhE2A7WOYO0h7EbzcxyznsY8krZ6GUtZzIs
Bir/gbQ7KftpC275FF1DjpaQxn48i1aArbkyMsB8fL5+HH7+vmEzRHeSIwuRNusR
SQV/I8bFifWbvBnkTul7Tkf717JDTRl4ouJOMShBmlB35uGreQWBbWxo4miNPOWT
7N64NsO0nOIZgjJ6RVMp7q5A2SmDMbf+r/b4jbZVAcYw5y4cO/uurLi4OTrBI/+G
/YyYcREalJhOnQOxPP9iHzN8bYDMrGQOGC1jFVe254QOngx9zH9cV4qJGGm0rgF1
pIGBz1kpd/FNNw9zHZNAnZ0DV9Q/eohD7EOTO1R0MbARsnxLhMMcxaIm/Z4jXB1Z
nIkqVPAFwwjPmBThg7Tdzptog7lHpSMTRSeXRIY7x15YbvpeV72tPHO+F/7JR/Fe
zHNzGWY33QrYE/cpK4mjE6z7KoCwc03exHtCBcqRuTYRpZ/8mz3Qr+sf0mPVnsJt
M9bYeQBi397tMqYwrywq6Af3uq3fHQ5E9JBFC+0uc0/+OYkKOMkuuq7NTj7sdug+
cjEI7KnTSpsxF8xABusfdCi2vIyt6Ip4qRCTjetIo3ukib2oGboiKtREUIvXDYQK
8ToVIyk9qNkDHTeTpYJQVpkWyYfjIZ3WNHEhNC22aF2cRzExoR1hA6HuFXxJbPEf
WMV20JgmMG+HEcY2/ExF6Qqv0Ha/+xEIEEU/Tz65tfw5vxbEhtiEYHfQPdL9zJT+
13Qgp642eiU4snxZ7LdzpgtUhgoTCzEwlWvmpwXFKV2G+wZhpLoye8Emied7Ac1+
A3RvnIj7Rakpq5awXjdGB7SniaYXpcCRfRno4bjiXV+aJlA2Gi2h//NH+eKu5fDq
6X+GszwFIR83mbF1VAaPvCyZ24F0cOST4SGmz4+K1GXXcER74u0P2fWZ8g5q7apC
T3XRUv1qSWAiUsYr6uHxsiYZgUMRM+lGeFxmiuuNELHurh0VBXwIxWdnqGcxftSG
OdGs/RDIv/RBswIhhbE6Q2IF6FbkKjSw8A6Iqk9ZAeoaW9QH5o2Z2IVolkA9JaRn
BOL2wryISolov9n0o6Lre/b3Q20GAjFn1QD2Vf2L4Gc6rkuXaIJhSeA5SBvNVov7
lbXcbtvo7JDQdlVKEum4xNAOq0qlFj9EFXaT/Vc9LSK0LuA38VEe6I1lvu65xQ9F
KCpL6YIWP5+/LFEWnWWOgeWYSXRPgQQXgznNBrWGD9foqYFy/z64/xf9WoULKQX8
NTGYJxH7U6Sehnhbn2UiKsi6BvdML0mvMU9yCtBSLmJdYGRXlr3bP9r/p1UVab/d
0mk+0ZO8I0UsprMBa50Yf/5Yn3f0Pc4k5pUjiMXieTnNsxMta7RgrTu/nDPvvdY7
rggt8YEjICP9i/7t0Yz6SVW32ffSWFHdwsSvnk4MFGgsXYz1v58eJSyDleW8Iz74
ra+SO1A9iCN6sD+TnIqgqT3KNF/++CKAe3alznKPsCmebfcNrtT0kHg5KddmNQj7
9ZF36Q62eUmFFl5dzp53CB/J9dm109cMOfVhPQDelTXVdvYGzBv9jYac2lkrAmdJ
Z1gfmNH5pYnA1bWD69YXRkXOVpdAasAu1FRapO6KgiBefEV6RZGXSvok5KbXJCgX
WUn8t1GU8C8LjcQk7NSAaPnZPY9IpU8vLtfXONcSA5I1Zi/TopdT6QqyqGGqSbLV
WhGTmKGiDwaDaMc1WG8mkQcxFPPDI0kDYaT6t8tt4NspTvAzrmo4iEaGkZ1RUAv4
nPrv54V1INV7tD+DhgU0vN6f2e8vo6FJd7zen85D1PdRLIDu2i/+/7C/KmdQdHNj
f2mMrFJx1NIhP9vvxIguqJzdKaepJpL5ya3ewr7lZr/ZqyX0HNNMmpk4dNV/N1/d
xHDjrDkLMp/eYX/FNWnXteUJ56iIeTPOtq83NmM8q69B58ovEgKD401AXh/CURUe
Bcm02VS+LlPtbiTw80HrhHgSG6RHFWQ3M5ia6HR+IKHpxFgTEC1FDTAKZSApkY9y
DUPpgA1v2KoXk+KpkKLDn2PYRGKvv0X82pNUiHgmJFdfgFtDuXMWSINMq/6hLgmZ
4OC1QaY8aNa92rQtPQGpMClPgCXG4MZLVHAg88Y45QLBijYl/ILOcteZI0w7miez
sU55+Ek+rqnrmWHbMeHjeT7MZZBlAYvDbHze8MIaDIF2MLHTgbFFs/ivrG8fNISR
ny/s9SxoDB3wCFLIJO1rFz7lG4xCtFuAfSRPyeIFT/1RozcGtBvOYwn0QFVEvSAQ
xaxFcIawvdpKuoNDzpP0JDqeIrpxOsx025xs+9H7gmIw+z1YiAqO022vGzp8fJyl
1kW9DaJMMWVTqQq/gWXhaYS8ON0LChkInbyYcg1X9IzGmjHxczqK3nL+AodsJK7j
AU/PVCiJiB3mQVshHB9J/G52C6BGnT6rJwVze1C9mrQKfxopLxX5ZY3raOzQdHk+
DoJCDG0JRgW2KfyyogqMk/EWycA5MA8c3e3Q+QmPr3/4Habg5EAQDTqUs1XLyOHa
XrFpfSD4UAKlR/HObM+vPjeaTMJZ+nK5JXnLSs3sdfDc9F9j52DTjrN1xCPNZrqF
oGZuUjOreO9EfZL5ske2MQ2eCwkdTnCc0dfeyQpE2Gx5nAv0TAyj48HqeImGu076
iVYwFdPPSOK2S8rQ6j9jJQJCzWHswuVoNRYJcw0gaCKMDsGsg8VGzfXBzOuQDro1
6GCbn6f/zhPGlXENRJCjfhF3MzLAv6Rr3Rt+Te336D+UwM9beUx9qXtSb6lli0VT
t0Zr/Dr6B3XoEbuDCIRCCy+beOQ6yH+k7D+FapXiecwtyxG8PwVyol+trOwv9Rxo
UeKVIb4hBWZ04NbXMPS8YLdsF2VjxvVplPvI77MfWgk7B5NBAl6M0PfeBlIU0Ijb
KFuJkucWhprzEEGeG/5qrdLM5CvQElF5cxoqe2QM12d6zgaBJ7IO6i9kGiPIK9bj
kgTLQELTqmWlD/AHD593SZKfjyTQwmuGH0uw3VMHOYE0/kI9In+2q+FHZ7Mh1SIM
skQy4p1kH89qOUVD7aYE9+60vDtwvso5uBz0v+3TMhBYHgbfhPK97mnupTv2GtiF
98e6Sg0IsIGTUecLyoM+aBh9IXPLy3bq9igGA5sqr/N4/CRXjOaM154KNOkVAcDT
G/LiDczhkJKrUvKEB3GLO3dL7XREodjgVlyhn6uJPeXw7cbMqQy9dkbqknkoPgQM
ezN86KfrWAp1pdUjcksdqL3yw0Rm48G3yb5W21bz+hxRD6czfsjXyaPu4ogadOlY
3WBkav+jGah/UWfD5rx2frGqmwVLDb+Gfv451lKJ+W7eRSymZsNs7fdO1I8apTcp
GGw7iB4g9DjUHfbQ8gtpWIlqrK7dyZ2SdFRddNAWujMbiDf8Dp9hFts9g2ByqE9g
zDeJWB1OX8yarXltLrQ4TXAsdsRfQKxKPkrCzoemt6XKhCLpDIvLSBf+N5sdLRuC
HZAPOvucIQHsN2REpaaTQ2/mTRSH06jmjWX+kCZ81YsrZUO6J9V7TCMKMOxwH80K
8EYgmYQ9iEPG8WiaqyHCamzmGTsAiptJmPXhRX0hNrZJ4+AJbK48v2HNyI/YPjk8
8ffaWS3MxyO48AQ7d1d5Ixz+pS1FRQ3dK50sDmpcsnmPZQ/oKxmx5cvJzhsfOg24
KZyk0sIfkN5NopwD70AugyKn1vDKyiSkYI+A1SP0IjxjmvtxdzOb5v4zXDWhire8
0/H9T4qfo3AscwyQjDmPxvIclQ3+hLyCAaT7h9bEujsCO1Hk+MbR3lXvbCJIaWia
/EzOlWO0byBl9ftpIk+BlRBt3tIQCHEDobXilLZNO1lSnaA9VhATWq4LOktEOeUS
x3P/YH3OVR3c0adARBVo/cSmP/PBM/adhimK0VvGlEOC7YAkoLL/I1MmcORZJfPz
l+Jy9Qv/hBL9MgoeCNPcVy+lUWUQv6WpW+qBFvGXRQP1gyhl8hWu1eG3iY91e6xv
Rl2Rp0eYaC7P2K/l4f0PC78OEnPrteYyBoLh+TUjln5qlQ7VMAgeeKTIgp2BclbQ
K0vRPCB/1aYGQe+TIX6/vX9XucQo5g3MCuhfR96h72HgAg/26HU7zmrHfDR686AA
ijnP9M+lyuk4T0ltr6ke0IPofLKy3T5D4tNsYqptb0RYe5iJXoJmNKcw7vLU22iO
BSDmt2kjDvQ+g6i9HdQ5uRbiPcgvUM69pgyoGL9J820Jiau3yJP/NmJH50ylWnII
ggt7TNMk/UwPHWAmT1GLXOQY9+pklFfWMN6gasiX7+0c8TmO74MiIwZoj8FmQ2Fv
eJD9hXTrOStQYVH/NvQqTzb5ORA31sEn+Cw4O6RxZ5HdwglGZPr9ZpbZbD3HopuU
6tMF9kQ/9yKe2lp2iuWc15cm5D08VG3KtUxatTECG0nf8iIscWgfcgrzU/BdQf7N
j8PBeplO9Kn7qivv/MOE3eZeDEpYd9PlGIAfQ4tLJu3neSaRSYZJ6xf642Cb5ciV
dbGVpwuXhwY9ajvgAdSk4uWz4nv+mK2fAV+vqVb9OQiKVIGPKsso5cWtgqkdWlLL
2b2sT2gwS4c38eV7JVVNMGN5P0tdgKpaGu8tl5Ik5uWzk8WFWEtRrHGDD51UBygE
9YcrQETw82ydOi+3axBJhB8ZiQ++VNhDuAiHWiMFHQKmyNHhXMl9TqnuzRUVKHk4
bmZ+P2QsqcAjBwsCeOXVklpXKjB2MAJl1mI5r+ENU0M8aUWsRa++Q6KzCqwkjpXF
z9lFsC6Frnk3sFBx3/YHDbBg7bsImrnX6wgr3nqnCXAaXJjGV9T6RTpbGTsMru2F
yFoX39m+GWU3JCfl+uAkpXuyBUEdte8qr979pF4lhG+vEnepodcnmNJNtA5V/RTz
W+HtzGNWfcpTmSEeBxiN0T2M68Xr2xqiBeg7tadDmsMtIbI0CNAEXyP5j9oZK14p
4mIPuk+2Ah7+a3Fujvhlfi6GF8bNnuZNGO73+o1HvLL9dVSAzGEWYIzRB2gfSD3X
KboNaAXFvANiVs4ig+QISnWcsvvRgH2y+XaHrBlbGzXZ7uG6JjYdTzwEUSe0/BkF
o2SS29t/7KOr1CfvOO05myYz3bZFdcyKNA55K2q1r0arqSL1WN0F8cnkdhr6bMte
3Hz2tuDpKG0VP6FnDYlU8pcTtIKQpW92U8LxhXQcQw8S4LsHsVPm1wVfuMH+6EH0
wNmvR0vjpuFa8pVEmQYTpTzfcnrg4v4xDKc8XGFJofBXyPdCSJVhZpF+ggnvumZ/
8ZWoJInXaBdNU4SkuEgGvp0lY0qkDGMp9+r35hQosXuxsiRHnpAB1jocbwegvlAa
IsgyX00Rolljyl/doBJtVWCV/qiQhFSU4iROpnGcaA3xnmb9BjHKm6KxbzRMZ3VU
tqa8W7j7F2u6R4dqzOOHx4Eb84vKw0+gkFHyRCJAxo7R9hWcpB54ldoQhisbG+uh
RSDt0eYU7NwTgkUBPu1ZcLN85YHZcahc9WuYciu7tQmDoPjHU2PKvi1mvOuFgotD
VJ6053EVzchrsbqHeaMjqV0d9nLMgzB/ImMaKOohCdYKZduxVGaOcOlU75Qvwimn
1+1U4X35geEEAYmmJK/GjYo9po+OJB7ANaBwdLCY2b3sPaOC6heVnq/7x68TX6S2
Qbmzc+l2CWLMbcjbc+cPRmO7INUsoGOiPVXRpRxp+CVHB9uYGj2lVOaEa5cT7AgO
YKCbcgFVAdlPzhO88MXD6ZsE8cydz7Q+zGrroFYj6zKKp0hUfxbwCqKboZJydY83
JT1r+2460liwKEeKdAnTAJtHmPB/7N1WEUlVDD2DRQ3JXtO2Yn01GlYYsNnh/HRf
D9cq+nuM4gnpFxHN9hj7yJ9KX7sOfsu22zMWbpL7tzdyLPB5sS2nEqHZw+P57GS9
eeKq8HHDDWO0K8ZQFgm0emc8zcePk6RiGTSL2S1hQALT1q+Ihp91m2l2SN50GRZv
QFSHQJK/pEOOswThSKH8k4vG6Vmkt80Rw3t4dO7s6pLgBJvkeTGNBChDMrqUzr6w
HDlkA0kwmPQfooOcfOtBUV6Vl/YH9ud6WFxGNg4q+fo5PfNSy61lol6RNxu+O1yg
JUSkwRiGYPThIOrecXwYRFKSxymvlzKgBxP3SbTNC6/CV23itEkQVJKB5gtv9O7Q
VlUrvs6Sq5YpO1D1Vh3IX6IO005dDRswXvDZz5wvSZ2EXasoJtI7mfhFMQ9Gij3Y
XBW6FT6+qLhLWhnzwSnPJXVC3D8h2C3jFRutKXtBd3yd2QHgTEL0SV2be3m26ETf
cDQIweAXfTgiXE1UBHjt/4IJ/GHFehxdlzfgMe8q8/vjoKeDPjm/RHVL96ZNne4O
Obiu22Hu5lSpqf47kAfCXJSxmlPfZGOd7usciaM0NkXoFhkNCn0Nmxi30o8uWKdT
rhWBg3tiqC8vPjEN/lO/2vymYu5Y3DWwm93JTfSvZMtRH+JSoFZRrOFer/J75OGf
u9xQsfR+aJgfi1wQZb2dbg2DCblCDW2XZYA9bby4uPMmU68rTRzPB9gOePQmie4u
fbiqd25nt4HgsikRqyF8l0UEn7YtIlaeW1e07j++AspJZ0GwPB8gDCEQI2ec+igX
GAx2AquhdRAKM+oKX8TmVXbIpOTZKBNUt3LgdPaqv8kTxfpQwFUlNl1JWoQ4AEzk
xu6twyrocGEeGoj6qTZvMm1utP4IGfXpTJOIOm5Iupy0tGvwH9p2jZyiyaz7NKoi
giiXd6bTeDZNDIjpyGG44TU2L5JlpnSRSBtcNsyKTIdAG+CGemaJWIY9Ma8fHozc
86i9NG2uxRBhv36U4ggtDW7pbaAxP0STJw4wDoNi7Es4HD8ZxNrv9w6h6e8W45Cd
W3C//J0LtFrSf5S5Yg28i/i9tLMPVed+0xusHVgzVG6NmHiCp+HWrxnzWvXQX+de
9gshPt9y6icVDzzZRir2EBRUKO/xVyxU0PaumDazU+yKwXFVTE44kbcr55vRqMYU
fKL3gp3/FgSXoWlY81rHpPNyB3OW7dCDOmtnZ4MX+uPrh0S0WWXndYPkf7Xbc85r
nC989XtafwODzY53kpXLnVzZkPXLcWLnWsV8/UcWolD6/tbw4NI6Emm12B6gQlOr
6FzY3D2pDqyHYdfy03iCh4MqlsS0f0hNPf+ZICJrIdQF98wY5+w5FeUoiHI+la9g
ys/Aq1eOgwCDj3vsNoLhYKc7XBtB2Th52fbttXp0LSWKB0pN9jqPzqtSmBaqDPDt
xvEjJtjPWbKD2iQV5XNAoYSO0RY9nvz8Ol0PBc5GErE/0bHQYQBJPLxs4TD+vXwE
EgvSSGNVhVN+yg/JT+y5YxuRnrh7F2rDkzTMzpQGJ7Iz29G9c0xJc6E+j30vcdTV
igcWU8sS4sdz+RBPsY8Czn8nYwcb5rLqHS/5cjySraPZmEwvCAIL9vR3o2pn4O4s
AeI77mB7vqDtQzIBbY525lld+5kYsstu7KwrIHmaL15XQEvU50JkgG7cM5yDHYg/
cp9mH1BjQ2Qhz5l+3OyZu2Jd/85LjVGU8zoTTu2SkMk2EdhCT9p9959NcO08teKV
y2qJ023kiWRRK5fl0IwnzkLhfJ7fng67BZSaVR884sft+K+IkjEyrD1xdmQ2HTHW
Tox0fj5ppZKaw9LepsXLiphl7YLPaIuunxnqIFQIawu08SCVrzq5Kx+A2y0nqbTO
5Czdb98ichfsx6udDrO8tP1BzpVaI1pik9kM+wCUQVBHfijHf0rexLfQYaxSe6t3
kXDL02ucyDpgg55h3Qqbq/srYJQmLYfIc/8K6pgXeTWeyUMFr0qVOmDLAKHnTsRG
2cJ5OKgT1XJ+dn7VkkDygYjk1STO7yGXJ6AAFTk1C9GcRYvnIazWkEUi0UsEcp3h
+xA5JW7YHQgNhAVSlzYyGDKpUry7eMHPn3o0vKU76QmKsbm8xUx0d2yb3wcIYtag
AwO/TB/yxUV9oWE3d2rr3XihiiJA4aIgYNvGKOH36e9+z/CmAJreWDTQtxzunc1a
ePzBxji4EhpPBOs9nxvK/SLQLoJS3faI3/igMgohFE+p8sMOnd928M308uOewMKu
cnkjL7832kvNDUH1AdOVRwKpjbf0kJnENLmm4z3n+2D25G7MnZY9+LQMhyA4mmEH
x03baGV7DBqsCHuUMfHfVhIYC3EHEXuTO45PY7+F8vHPr5/XWU6lLPK/N1L2z26m
CIdaycXf4cBtZJ0xfxo1Ci91Ap1ZOZfvFOraF2G5DAPFZQgBZBejv01bt2O/p6H7
bdB4l9N0DLiuLatCc7KovQrnSqn7ofLoa5EM7MzG+lEs1bz9yPhWRM73EoQiEu0e
ZPA6pSwsyCbufCu7xl/TqNsWyyE16/Y4viqxwGuhbWXXfxajdXE2UBg/Fb2gNBIF
Ugurn/iJgkDbS+ILaZRudPCk9LABImeAiTx4Y9JBaMKwIaeqFhVwCoBVhAwT8hYP
cQ3yEU5II3J4MJZC6/BPIxc17J8/S8H+VCypOJ/VMJu9rfUG8Ynbo5OTSQ32zLzF
+vZ+tjBuboXUZKi4URF9x93gouwnovdlysRTfGw8DmdiFBwlb4qOBKni1QeMw9UV
Q/pKH7Wuk74z5q41GBmBd72WmoWEpcg9e7avYfLoirJFzaRG6RviC/5EVco4n04w
dIiwFkRteeJzdiY6mOT4Fzx6UuWiAmDSt1MkJPI4SVzKrPhJdwImCcbtRG1U2c3c
dvM4d/laA4jrHwlc3lmV3VXWT0cMkAw5JHx/R3oS9wfPr4lIvHQsnxB0ZVC03LfU
HyWvwRccoBmnw7BB0GNN6Cv9k2yfvmZ1IGFS+BT9j9CPrjor9IhfNcRD+ANTGT7s
dGLr5jYNqoedN2qks32RGWXrCZu1YzidUVC4+mgiCEKQLeZoi/slGaqEUljt2voi
SRwwgabQub2IENKlEQUEU/L7ZaWnTPKWPdo6MHXONSbVwhGNTPoxdWsVNp2pnlvD
9slJalqRyJi5HObOREYjQ0yCSHTW1n9oW3kwunL7djT9qb2adbr6/acTuVrUAv8g
ROVpSm1K2hx7liqu/7CA7ryD8CasbJzxqY+ObHwFsSJSjcLrk/DVVpzARjXR7qW5
07a4jCUoXET4yzhAftY+hZgtl6qJJ5eVMA49k93F9S7rc5dDG398OFYs80nXlL55
AnxZVa9YJk18iSgsPCtG+JugsA1FwFydO8XBTRTvRk4yrz3Tj5PQ2TkY6sU25Ked
wgL6ovDyzj73/fjIo0NmzIIanwNvQLSYVIHjPzcMVxZtPeYD2e5wfOEYHYXWyEb5
wDtAdUxX75xa7/XtswiofK+4eYmHTdYTEq18lnwHEOTQu9FjHtbcnWFVEW3+73Iz
ecXajbkMmNyq3/hdKWx9oeNbAPulql43mP5EaTlpnqmh7SU6iReutJ2eux2Q8Rr/
WyOFtqUvy49RfIJOfdhZL52ZuYauydzpDmnJruyV7HfIcdtpt3z+Z+gHSI2Rue3i
wr8Mko5q/MbRb85586vx3wuRrPex9jb1uYEbOoqYKg/qpOKbrmWs6HHGG5EHgmG1
MK4LUGuv5IxqwUKsXcX30Tgw29otQsTXoi5kjpOy+I+CwlcLpXHRsjhqgd5sO1ZX
Dvc/SUZ9kbhRVmnijoDxrsffCPF2NdUq9pNi5oTyianpcxlNzSiM8fQT5JYEV4ER
CXtsQS8nlYIchNpxdVWyEvuzcekPOwdEoX5SwdTVl8YDejreYuFPIJ8+d6Tz8TSa
cE8jCCDCR6D+lSYwDDs4UOANZFakSaARAOvZxM2XhDJvdge1osWpeEmKOfJ0zixP
hME/2D26Fvw2oBwQL16EBbasc4ZZfVxlc9DEkYlG01MGUfaPC1/Une+9XFpNNsfX
bI6Cbf+7TeiaU2a5TiXTvOiNreihSe5SnMgDalJee0m+Ji4JRJ6CSXZJjUe7UOAb
Z6PvGrav3FLzlFkDR6Qb2uDAghXl0Z8R64QhQGmydgg87igokGPJT+HsSPewY8An
9qA+o6ykJAmf+lY6VECZrXV2O/YPlrsBoM2JqDNXJHVfJ+qMsR9jBCYu0ubZ+CDX
SeG42QW9mmJgqF/Os3az+TPvCq9PzoD4eZbYHbNaT+C/0MaGCXML/cMAVmHsD/cj
GFqRkEG5W4WK1e4bDKj49sMD1dQjsLLfwSaWZOf6qUAQFl9fOENoQciahnC9dKSF
J7BevChufYrbCcHSErWyk2uSasRm1+rmg/pYj1yALf3DAeTPknpAY7hMPF7EUd71
Cgv0n5c8V9ygpor3man+BEKbkyKRqFDeuhyoL3/3yysZpv/JcOA12mkuAMCAR5b5
MZRsXTrkg0jUr4f8CJlaSIFfxm5LmQnI6COYaQ5ry/9VJDyUkHEGGyGKzzI+rdDP
hwKQWckKeKyq6hbaB338gDkJIQT4cSFNOyJIwKMdUum8qVHRHAgB54NvMl1D+9Wy
WMl3IvurbUi8orlqt7tWTE8pvtGEEqgiVHgqX9h0ObLYXcgbPgOyhiBG/yVRzKk2
VsJZmql++72mmIz2L3mq0EYaEjE//mwZ5Ap+kyXVSKjaIpPaM6HehBb3lUeSxGHn
NP8ZLvJI8PgzpAHpSS8v5yIXhzRBzKJIEG84OW7CqUfpxNoDmLMe5ikAL9Ytggir
KDumwqiWuPd0GxliXzvQ+EZ8y8ivrapcezqewepKdsYJddxqev4N+0R4YyG+yCDL
Og+g6vjUsgkF/TmVSHXyLNcxc36iZ1JdUNrWgMEbHac7pWoscW5esZqmnlYHFsRV
g8nM013z3Y+BIbh0gRWk0PBHftK6hVzmQsoC0RYgL8N30IDD3uf83XTzNYIhF20h
401ACV+NLoVkoFKVDj8B9HFUAgMwh0IqeAlWH2neDC3dsETSwsssSClf83M4+5aP
bTHnwYThEtiVGjkfX83rzTlbk7NvUbejIfPVAQy6FKZUqe9d6L4nOrmxnMpMoKYe
zL8FAZjrbwcU/d5OFNZ1YNxoywDF2oxFfL53+45WYLsmC4Td+lrPmqUHbamZRrCj
/Ce+yPNKyU/wK09cRP0NJ9mZmYChP2xR8yKPCgfdknT6KO/sBP6JDcqHglePJmac
gaGJzIUzDhoH2weRFo7lBRFTufV2e39Hf2MGb4HrFU5XURHPJtiIrqw77V7IlVQf
tZxk9GsL72+GCQKWaW5ptxQmPcgVXc4BB+5BgQLz2xqbi3YmumdzexNMzh1CkEYC
TDO7suRBp2TRHBke4QNuKRu7p9HCb5CPjouLiPIaLSjrvPmJB3haZ1pGiQ81kJ5o
jpo2XeP+V4fcv0Jfs2tym6+5bNdwpFeK/cFutXCNpRABxbJq6VlOgfDHIvgSX12g
t+1jATvGl+ntdT0p0+O2bhkxB4rMg7ymnjgoT+ajugr8iUu62cYM6HZpZyxrh2hm
juBWW/ZCD9c1/vih0eBhhXlSAi6SZD5xHZBHRyMfZ4CiwP60jbOZNDdXcbXDd4Bt
hoBILCIR+Uc4JsTI8cRneKObaX1q3sqYjfxCIJFlshN1Y5P4C5LtVzQRFPRZucMK
oB0k/U3ugDyWReOwSfTRAlSSTjqiELIhPVzdykhJS9IIBNr4LyzI/fGgJG+SqVh5
5ZiBDeEXxY8XtbddvWgNyMjiIxLjH6sUEz5SAQMEd8KGxaYsmXwwpEWeCdZLC698
HdB97GBzZ3iPonlNJuYCuw4oOhQWgJXV4OoJWS+Q3RFzMOwZ+NjeBy8kwBTEqVVZ
kZfMkZvmOw+HT1atM/Y04rYZ4MPw5SZN6JRp62zDZfR3N4i9h9NsMUzdffdR8mvf
KZrJ7pGEvm/JIkenFgRfOUPxZwQknTz0bq7il7to6gk+q7SF9C9w44RFtpqifTq5
jpYYCMOaXC7+wmsRJd0jm+H5GB4dOJf2k/EVv7MtCnW/KJwqtXVGPMPk6Pez3gyv
fw0Sn7H4+gRhInXswsuYxeQTF6U5mLMjWaTCeEmrB9NCIiqDMWseQEIclO1oMRoV
PHKnFGvtnxe5HmsX3gVszjVENRs6irVHFJWIEsryjFL0byn0+z1cPmKga3Q4W0nd
LYuDJMNIfFeIu6tAyixZar45zF7cUAfaozb89PTAmwH0JhAhWOvARpqB7b9DVSCd
BsgpW3hCQbHyCqb+n80NzRidsZdAT14BBl2lk6/Ww5+GT02MVtwrBnNWLvTJB86M
0lz7vUhQvkoAsKx4M0Qt+YK6v945TZa2rHFvPAzNT4VkpJyOdZT7sLKrVN8fO8uR
k7wDrka1Ek/KTjfjHRzCL/MJ2O+do3oiH/w93sR9Z0jhkeehiC7lp3sgoposwQHS
V0XSoBHo0Ox2drzKlS589AAnqAn1RaeRrH+Q1lDeNeNi3m5gzgdDdW1f4JUPK9ZO
3tuTyjdFRRM5n4DMkvKdwq/1oNd+DwklemFFTQhRBeIJkStCrjNbkXatgihl3AjX
HMUVyp7F2sJY4BIYH0ddHZgNqjrR2t3wi1sdV+yDRzdc6qESKbppqGDSpzVAhMKr
1ocH5G+MMYkRBJEAhhlLdhisR9HJGeyCbctzoX0062xAAHqpcszeJ5ANJn74d4y2
gry3/JpwVwcWeLMOvY9MvB/THChocY6yXmn3HJvjzr69ope/0NRV+sEhudASKS+8
gcuiLLe1unQFRIjBe28gmPSwz6+j4ipmv67iJFIQm5s7E3JeY317sv+2Jh9tf4d3
WTPaY020XLFgY2ebzAL+/EC5p2lOgGo2EzIRiHn8cFUgOUjFqVKMqSIipxES/t5p
TjE+Q1uYBhSK2ZTXd4P/YH4B1PsjUDFc02Zylsto+Wkv+PeDRKs6EqwbX9RXu/Fx
S9fpJ1SEHTCtI7NOoay2XYzr2bladNWK0Bye2J4sFbFRZjkrIV/98qXu4V851WTx
yU1HY2m+W1j6DLNaumU2wAqRJ5pdAdxS2Cdxu1nz9zQSl+nKNH5bwZxRxsdkw0BB
DX7dVEeswTzJ1LQ5jNOHUYtBpPTZH7LfOhijAJ5ojnPPil6e9ARDpgOJta1Or5/k
JGScXueuDPcCqdE0m0jCC92jmTiHRcLMBhsSylmIh06DPd511B1TIcMjnSO844nU
H8nmA3c9xOuEpfP3deXr1t/3R6U4IlWLwRBOvVNqlg0Y7Lcrw1Xy5mTbVu0EfVmQ
bQezd6CHBhgY8+z+79GS2lh6tOcGoRNVgv2nBbnQ9Tmxx+37dlx/YMuwh72U/hh7
A899lLidS2Gf51ohdOEryHDJ17tP6JTG+Hi3IgwV1cMb21GSoV13gQ4lK+5jPKqV
98v2jx80iEVLab0M6GCCpiMNafwUGs1Lf/hrV6OZXc9ekRKpdRvIvhWoc27FMiE/
nSdn2Eq+rOg/Ckz/WwiqlDTqJw6Qjv2yvJ7ytdcnaE3vCyPk+CRmnRy6IcdK9y11
30HH/Dd/jU5/nbBt3lmTULJgHMOyw06P68Fv0KlkO0JmhVk1g7UXwjCIBnd1IFOa
c1NL89radIOheSbKQk0Q2ZS/EKEed2eLJGTt8hKmxQZURQtn85Wl40zYMN6jmLaF
IGQhLtgsEDtC5gtdfHhP5dqLEgxD2wOjZ+PmP1eBqx0noAQ17/P4oYeuGAt7dIKK
dlNtkWWbyMdQt0Qpo/CCSedOjWaIwTgv8gVulugKcEijxxi48v1Wm2V+DWichIgI
hR/u/QHp7xk+D04jrrup6Tqz07nB4qnWBc4J52oiNKHPJ0Jjti/AOcIZ5Q0wwHZL
W7rU8QlSA7i0nwpBdADpNPV0n9jRHt0BMxrfXAoDsmCJVs6bFnO8Ez1asUUekg/p
JAlClSgYN4HrF9oTSrrPiDm0dhkfdu9/QiCGRl3ZkV+l04vrATRdrOF39DPr+pPM
p+q3hl9BaArbrySKIgFidldW/Uve+lNyySQBP6L6oGoxasz9gDiePEZ0VWuTeE1t
jZX+d+YSbXED6TY3HrRPpsvuaU+rXS9mb8d78Ex8BfgyltRXtprPYXbE2hISi0my
dme6XSumVko4NDGgxHGbqck9sbZJ87bAOjU+1JnxcdafL8xNs+k/p28OmN38yM5o
ixP8oVMZKYAIPBMFLi5MxCIqC9yNXuMufC4OR6c/G8kF+Q1QfqpmZ8Qa/ZshWRxk
ZT2nzW/tnuUISNDEco9PheV0qnWei1LB1jWVi8bF8B4Rr1/F7WaHHd0v2xhFaW7G
89QoxXfurXScefwsi8f2WWCzeCvzK/fj5wj+VnvXO63/er5MAWS3q7CLOp+sHSe+
TUMUdSN7k4oC7Tz4nSlYcZ+/2sQjbHheOLXKsypQf6BemQBudbXv5B8DIaouH5pg
e2RzqbpoDYI42joZMOckkpDs/4d1J3UBgCB8PPQnizUTtjESA9p6q3/x1tm7swfJ
yfAtKBNI7bF7AIlBLLxPSEAJqGAi2o/hjOQzrAIXirhJzzK3PlVA18SAfLngEL+9
y7GT/MyA3znsMR4izGwy7IGIttPZW6CqbpYojPIqlqFDpQvO6poFggtO4oEjuTGM
D/MXXpvyX2P7G++6hMUksFEApMdP+tCHlneWibaw9wZPzzCSvjqlpTte9bUmiGlo
VkdoSZ143dMLcLjlZ2MmuAxOPVcUHe/tK90zPqhYPaURkyS4ifARgcBfWlCZRVhu
migp6A/CtO2/Ef/cnGk9Sa+YL1DMSOL49pNsweWEhxOjUjfSy2yBiJGeFqjE4Y4+
uOGhd+/QDg7P7p4v7mFvMKj5MAnBnVufHL4cHPWQPtrqrnt8/HWi/pcpU/9zmp/+
Da5R4p/eiisb5OYuQWHU7BH29hqWW5LJI7ea+XGOekA3A/yucnra10vg2FBD8MMx
/7835Sqm+tUEGovMFu/820c6u2T562PCvoVGXSAX4lsg7pbOOYTlS9o6z4fdgYob
XoksiWmTrs+PNpJ3RKN8KNwnbM8MWjAkDmSNvDvDIwmTXDOS1/vQ0FFuBdKlHdEq
zoBo7vyUceX6t+jo3u4Lu+HzjxZbpXKxsIIHe7917+xUzlB6CAiZDVkwPpiuY8Cu
HwfnwGKOe+tsB7KHTgqLq7OjvBnH5GQVX8BgmUt1eWJyxv59zQhDisjbLnb1N9nc
dkuQfc/hZd5MjIHkDPfCJ+ocv/plW4hS8z+w57k3IZtMMiVUw5EXeUwpklN00TTG
pS4EMkS2lKwhGR3JKhF6MFL6+Y+y8SNTfVmT9wZTF8NuTUKwGbhvIThlcZpu+GfK
KFkvj2Xl83nN7NPNxZAPJX2BCAucWjpSt7VYTz4xGYKvzJzegSVcwvuzSbocM+dI
QmU4MPqSkBtRE5mKu2ELJF11pI1XTkua07hKDeeaLw/sWDuycHw0ZoYwUKymOa1D
GFJ8s/BlPUSbaWEUIhFNmrfg8FtUNDSMeLGaczInYSA5MBpMdHFy2BE4RbikQiOa
+P7W6VTdo7GtvOr3NogD+melvjUiEDLw6MEbSe66lEpKOQefcRm9Xlgn98Pvcjx1
Yhg9Xhy4UKqoGvMYeR1ElC8VrM4/Pzf9Xs8763/sMu7Gw2vtx6FRm1j64CZcLkje
8V7GOPO20zsxJP60iq19sUrRC0gn7VecKh+zFTYHqPc3HW8LxcGI00F2Exu0cdL2
MO4GqB4f5/8TroisjlgC9tzlWnYsj8beXgFoXXBBX0920D2RdP27z6u3B0GQd6H2
2SwuoI6TFTSE6Z84YrbHK/HfQVkwJmycRYbkOCEUTzxooSU+MTF3ExZwkVERFA1M
fepDlnqhVPhlyBm7eH9xBNGZXI1A/OZMHbYO9isPeVgQLBLAxkQYuqTv29UM9nY8
7L1xTDkuufUVSPVv3S0ZYTXYldvH3cCqkmzY11IrA9aKzyx8ogxlm18FXf4Q+BqC
fxhtzrHuSSfo3YoGS84fAEqxA5hPt3mnLt+nMFdIcuQMcJjEv8HnPDnura2mQYCY
R5zIwgAHGW8JYAIY9eHDzCns5scH8uq1WyE1I3HQIFn61ahEg2LZoNV7NM6fx2MV
u7wyZEHnvHAKn+ASMuCm9EwhczgbrunKW43tj00y6EhBGR2E4QzKCs15STyEbU1f
MFnSbxd5fHALrVSLy3qW/wLTXvRb8d6gqINOYWX08Cyv9YGJxOZYLwS1sHKDgDm8
0eSqd7qY7KQ7AmtbPT4l2oIyq9O5vFaiwOSqeAKFoQtK8BTNHR4W+f0i6pnSdxs7
XKYK7exNlFI9JUbGUoi6Qq59CyWqr2pMOqZWyWxwWg2vJU07dexfGpBQhenstjIs
lbfcyGpkVaFLGwThthMGW6Rkg7kWMHEsCr8sBrvWG5owUwfUiKNC9AqXqQPZge1l
NKm+ax3DKAkzJ56xTZVSuL3nV/pfHNKh8jCkhc0lFFzxnboHj1mfTDuyDOGnb91T
Wh04XsEbIRp7A3By0tnOUmXvpCHpD+2TM0hI1Ig2MbqIYwxQxkAO7aVYKooZrubt
UI8btsh9yBJeI9UyN29sQdoEdTRpyjxU4fgBjKYE/NC5tsFDAvdxv1TyhwM4VvN3
dIbkgZ3xJFOs8xZnKGKRzX4gdBpAOv4S3Akr/kuqxSmkkLYZv9dp/2qpS6QOhb2z
Gdu8Znjrn8uK7FcDzD8w5e0q9yiPb3L8z5/9teeEhnLf6o3KujvUum9gtT90Nk0p
e5rqfGghWKgneN9Re63oMCAtmE7xwOp8p40yKo/1HpoRBgU2QyOtonTvyoEjbUBa
buyA2z6/c3r3fBlgJQ8vTRPFkqJPt3X8n96nkODjkfawuZXdiN4iSzfc30Q4BUpR
KgoeXb/hlZphT0PzNhKAytObHWyA3H1Za1TvquCr2AS+JxVsLAxEJ/OGutwFqfwy
fYA7ieUMvhQc7W5BGFr7+zOqarhDKV/yOujXcHRWSWjMA1EkvgKMNQtMy36zCYgH
rGB52UdTSNLVtogVGwk+BEGfTXJhrLQFBU8vqNBjOxwlL1TLc+oH12iAqzVLwGZM
D8FUnhOSAF2d5t7OMNuJV/P6ZgIeVPP9ttlei3BaxdxAEGTcpsFXYRB3mgR4UGvS
ooqkKrmNhS4LvbcJw+VzfgDh7kZgspSnQ0+xymFdjSHL0idIs75h2nJ8E5O1dUhX
u4ciAzJ9NbFO9dqyDNWkv3C4vkdpyDQxMidhMNVg8LIUdZQPoOuQz40udX2QgmDA
I6if1yvpWo5BcyFBWnIKpCmIfauA01QCrnhyQwXzJOk44Nh2yGWws3qWxaUSSCZs
NrVSWpqsr8iQZD4J15Zf/0/dbSgueSxb9VTVC0YsoPQ2/eDWcGY1l60dNu5i5QPW
3oAhIcp8OkEBoo9AdneCis41FFo0YTUKH4TDTnHIB/mbJLPg/kE8yVA2XBfRm+5X
C0Md8Xpdu41lHqDVPboUjG78ZJtxy16zxfdalJWnvm1QaHiCaLT/SQseEP9Vb4Nc
hwnzc3UtKG30o4EGqx0ndYN8ACdBMRcoJq11np6rU7eT79kXiOJBn4RPFPTmv2ke
jbeYSUfHCyJ99PPdsPK3ombzeqPoEDb4P3v+jZy+85zqG9p1xUY3Ni2UwbVEefiM
SBLaBOEzDdRW2IKkQ3no0zaPc9jwVL1uH5jDo5BRKBrzW+O8jY/BIVxNq1L9jg5a
mU5pXzyvv4x2eZH6oFx9LBO8jgmkhVNvYCDUylI47ZB1W3NBuU1W7fO/oo0iNbCF
0kiVZmkGSxcLOhLE/L8ebN59tt+IyzCTAZAn4BR9rbmVOh+eIRwIjdtJ2om1iMFX
qDvWdKsLrQNLFt9Q5Z3vUMyluowb8a3d7pHshusClMW7R0XtcvOMWSjxTnuyK9Gw
hOL9npdUhXAGVaiHxIeJrXS2ExT7Gw3ZKK6ySEjdzdj5Amx4CCL89tyk80M8Loqy
ZK6W4m9dbV2LcgjGTxkCu+41i4iav2fZAHxZDlW4sJycgg1u63nbJu0fsEM2lbWA
CVJdWKEELsPiYhc6VmrQMemBtHs2tYzR2PhJQXRPNHjh9a5qEoP0ht1cEdYmS5+r
3On4b8Cj1TFLnfFMvpOnR8U0+Z9VfRLCivsG3F60R48YF9wAJlglqZ3e70xtF610
Xalwx3EjHNbEzh6pASRttvpPXJ7cWb3t2kq6l6Bs4DyCaz5AaF9/hgsdJQ//FgkR
CIkHLA4UaNMoBbtAYBs8xT7moR7B1fkNKvkjG2UWbMWQChob2HDBu5U8JILKda/D
h+/gmK3KJPmxz22ihxeUOhhph4dUAPc92lXU5Ln6CbQGf6sP7WDvPo4vjN7OFvMR
+xsRv0ONawburxjj12f1UWhbj5olCHF0A930OfTqPka3Pr2RXButxLdkbRlofRKk
ud3clqFuzFslMtJb+SugTdLjC+bDgsdtyg3x9NPAAu4DKth5LPQ1ASUZHn7fYeqm
5nYEdV1mB8dG5y2Sj0eabfIb31EPrHdr+9XCHjZoBC/mBgMrukIkNeRh0rSCYBkk
zRBJgVcwI1Oe4TQZFvDJio3/G/JKfWNRrLOy/GNHHDuvWOjoAONeNn3VNmhRTDFG
vlzS6LUW8gNz1tshhIU5/0269WyfCqcs7OiAR8glW2oQQbGBNkUSe2cTyclanImx
Br2mckTWYCkozYqcZy0Au6TMzBxifkFeacrhvnzJjix29XV2NeXyvLuXOzO24CRS
PTdNYVtfpgFI3QeZ8YWyk6OFIxenxmldo0p/UY7xmsXh/6ZX6XEQTMqBPDhLMb4s
Ow8TuqnmVHR9r584ed5OQ8fcgxUG25GnllGOVzC1/Z/LN2mckrx0W8Iaqx8VUa/w
jS13Bj/5hfl1uBz0Hy+CtSz6UHU+xA8wFh3mCCA808kUaGFTL8iXMec0Ik6YWH5/
LRwjuwmeznC55BxQu1GfMr933toF6x8pneCZcVYoAIP41m3GJ6MhHc7+5YytozKz
EWX4z9ajyGA2hqTz/DkDoqeQEazLrjKsEh96f9zVsAM6JKEO1qreWA2MwqqFt4x1
DbFvNhlsa7FCN9MeHuv6nVp7arRaL62QptTfGRhgL8I7xUWxAnZGBFdqiLpYA8os
b234c+mPLRMpBbUZbKMf3gPMMELUUJcCwpi8Oa22fFOzfIcWW3jbdeEKMZnHdwJI
mjxRzLqcMpUpWXHO+SKBTEgy8iFkrFs9XdCylR+xY1HTSBzI03Pf/1iEr418gGx7
Yiq3+t03LpK/zFrC/D4l34miefecTrKJkjMOwZerg2e7c5lacY+C6CKIzUnueuXs
MrDslI0t9JjPZTGE0W8sV3MFbjMORredmpk2HORYxjfMzVWPOemryqKt9P/0Dnby
3tsEQdfExYIZUGy4l8vBICB0lXCtQfg9meV8DOknH4M+p2gkhwEuk05MDZ+bP2b4
RY1jVbT7IZPhyWR4dhlHzjAaWgoZDSu7YxvRPiVgzc/p8Tv7r22YmLGvmvNcw7+z
qbrI1oSP7BENC5VjVnPfPlPfX8xMzXwxMeMc9wb8ilEx6WkCK6zX7pdXki4im03f
csbm90W5YCpApD+hBZ3KlsnZOGiO3jcjGVx5oaB709toAz94ntMaQ7TpUBBEHfj3
klN1WhKSoUrN0vBhlvQVChPKl/jeVfOruT6NysDsZQNTF2C5yRZjFc3nG5KmAXY1
wDClDBqviy7rpsAAT7pKWtUQzradzSNrn1VvJfVr3W0CTBsbMwk+B9b13m8RxGwO
1xyeJ39xeXFdTLNLOojWzlb6H8TROWfPiT4dVTndQ6WmUHEEVd+7b+j70Ra8g7Y0
aL+ToPNgo6Hd2i8OnFDmjQyb9tSfpFZ+8t7FVO9nRT+rLcF67MGQG4wLf7gDvviE
Kb/ULBH9dGPaQMZlslYVPWinC14hY+wBZpd7thbW2say31bwm+eGF0h0lpZxyK+Z
Btzr7n29yj2fdDQ2JrQKLCDygtPH1W8U5YwdCGD2rYopHuagvfY7Z/PObwrRghth
H2PzPcB5BpQAMoKE6U5BxChDYthT9oUow57wc+IKVpEwi82dsyLDnzDQKtXrjLOj
ZYd2BowDjyxtbJ9FKyg3spKRbDXAz37CPyZYPM28FfgVVgSKpriEFa2zfQnkf1qc
qW4/z3aaHqTU1eyYb3QAnb0f0YuUx5pflrYb4guX8floo+ZxEftMXd+L8y5fcJEx
5qqe1Hoy/HmqPNN10idj8eBl7Ii9DlPB/WcyGjiDwCwNcIyJh9tV88/uwWMd2K+2
f+Kb62mr8bbzpqy/VUc3WhamtvoLzJZPA0TJrhZYE8QkgeePTmCZNiDRMVmItVAc
jRyTjgUxk7uv+zP2R0dNqASwkxj8tVSE5kjwl5+9PNty/XKflZmcpZu0sHtBzIth
TeToNnR5D1pyhBXTNnvKFbzlNIoJbZ+OsEjBBSPgsJAv5w5yaLT7epYlnpQ2VcrW
DayBMWRJPC8vVHhBtOd4G4qioInAJcYztNTR0cyAgRNVW8hE6T+gJ5xRzAAiwfqI
hbx38KkD9GnvSl/HSl3DiZbOTi7TXvx62mkf/yUD69gmLZ/yJnK7XSXfSxIZDGn/
a0WERUsYWIhkmJwWMdh+RciUkEhmH+871dtbKaod6fau+VKxIVjWk7Tj4ARYjHp7
BVDf8aNhXwoDAG0GinU6WYl9EKJcJCvmxw9C8+JJPZ2/w91XAtDIMVoI3DtjQ0pJ
xuWRIBmdlNoJZ/LumJYofeqZRkjBqNCbRZPOWn80nP+UV3hG+xFXr0Ggd4DfPadU
t1UeEDfOHnYu/crMwtjks7lEbwhAZNInq79bh5bxQn8bbq6+Y0rgg7YQjwweqG9Y
VJWtk/hkSwcT3PvAF3HS9LkXmcsM1hoKipYQBsbLs46UaTV/aAJsgU3G3fguCDkE
VT/X6QmpN3G2UJWX0BjOWIPN/jzBU0nKJqHz+YUTZdbj2fNRai0Eg7hbU8tKlc0h
mYJ+1i2+hpot/F7vkK8pqqEg3/udIHSVx3o2dyjXb5HH9xCNpKIDiG9MTrCI4Qnj
/7/EJo25P94qmBynuHFkekEkt8NVI0IDaxVOKjOJNAtyZFDxBKBhpGppd+OWxGRb
zuCyiiBkXSNaRTCU10+mhSrB6c0kATDcQsKAmrUYmwtSgd4Qt8gO0nc6GLIetbuD
L2/RymdF05VkbuLBksHqjf/ihoTwygKEYx8Bh1Ry1f5pQtGPHgsqy52H1OcyvycG
T3neOG85smmyDIi4Sexwa9eHzFQbcrzWHjGu67PyGfIPMimQroYCm/har+2qn/ok
ID4vpuGZAwg8ttAkvX80r9GZ9/JX3slSJHwWg6Ix0hlofv1umaYrXltptFs87Jmf
McKDH5VH9mv9KrP7Cu0qkQ27AYTKq4OV0Q1uWEY5tT4vz20YFWODcBT46EOT34FK
jNZWlZ/OsZH+sPxu8GbD9sBtP2a/PSOmDCN6VbloULIuY+k4rU8zX9lasu0YAMbu
nsQaFyx1CHiMtqJ0oOkuXUEJQYGCNs+udxNWTN/NwJxIfrCz0eWoVjgqLAKZ3xg5
ENjrG3vPC5Papk3B3a6fIsP6IcYCbFduzU1h+DEwhRTpk65Eba/hFihi3QmDpo09
jOladIaPfmLIAKO42qQcXWSMZVOSu8SprSxmeKiiK/AHBUt9D5/eVBKJ2j/qBgW5
503YN4qyEDBuC8RbXG605PlbMAwFwPgRPAE0QF4tEnIgxkkmGqfaUTC5yNeAUEot
iYAfd6gOay+hfGXfTEj7XfSviMpQRXAY4VYtrJ5hYbfS9ZXtytMOa1u3ecOu9rMh
7l2BiaqTig8TXZrvGsywrp4ScFDay+720gtFAKkZTP39g5w7fLGrJh9ALRc/iWKN
8m91jWPKjx+/RjGeGI0j2Oc2j7QfKaO2+UZ6d971R85CrPJnBKUf2dArDOvoESUX
Avh+nHHYX31gsfxoPT5Jiq7OP90BCgTxSEWPPPxnxsnmkWX1cJtaV1AFFmtqNQWp
kWZv068PIngYlY1P7Kw4Y0dw+ek/7IriwTIF2VPSJUbOtUnLGeF6vqEuWuhok5FR
pInYPkyE/6XCrPDkbYcVFf2gh/1h6UNPx+9mfGKY4EoLkkSsIFIuJRklZp5Pmz1e
yAuO1MSmjp0qXztNVl92+pDDuO1mcQWnylwbclaVxWJRu263bp0szLhr1Q6zF1Uw
KF0G+BVG8wfHErBsCDbSjqYIxnszIAUQ+4zQYCOMBP55ZEJeCesKeDu8NQLpRrB/
Rd3mIlwWReO0juocNGv/9sY4AC5dcj/yeit5TX5xjXhgNFps8OD//Ugs1+FvW68j
4tlj6mAkZr4AKe1XULFa0EfChDb2pXk3TEXw5Ybs9nued8k8ivUYSmLmE0PSDJc/
DzgmL5ktsguhvjM9s02VS+Fzxy4NCHlg/jM42ihJ4J8PW29BCCwnufVbRH06aVRZ
0gMhykJLRhY7GukofpgvMIRZY6dTW3RB9iWPQ2vPU6DFtPF6f1gLaiGK2w6qL5sz
EiomruixlckD6z2oAvn7V9JnnRZR7exQnaNig+O4+7WHiSYzQd7hlU11sOjE7ufc
DPqCgxAD9+M7kdH/E+3V6B5oJOQn1Gk62856ZXNIA61GI1ZeX6iMNv86arLxqvRx
TN8noiRE4zcJ32/JmhHAn0I/mSY0TSXs0si2citglnTvTu9qBYgc1odGYOzDBxpk
DRW9cqcd/Acn+CQfKZRPV1eqwN5JgLX0S28FLWmqqVAj6Yw+/ihNofefODxAkZpd
NJQ1oxujBAiW9GoFEUnl4IFyH30VmzHbGnnvvj0gi22H6XEDUCMHBKCNKGDo0VEm
fc4NhPbBPE/YUirqQdddD49Tdjiz0dSS6RzmrMFTnHjnDZKKzrSyXXQitP/HH6Kl
5OIGC8a+a8qwTgaQaMTZvS5G19xAV3jRPvqJSyItWbyVc1QZuXPg1eSPVhZrRDMV
a0OvjjtxXPKlrtEwb9dmDWSKAOLs1xmec9tYdVvmcn7P3W5hqFz6SRg+OITZeVvI
e6kBYHenpxPjQ+S5HWqrPYkJMGsxSUfcYgV9PRC6EP7IwyVFpsrnYVdePk4CvpYI
wo4aAI27xhJl3Nj0qatJ66WGrKaNGwj/mqqs6q5PCGMKDuD2tTPpJfkP5Gr6PY/m
K+nWoLtUGTFRcZJy2ovtR05a7vxvyqVAvhQdrLX5C+V9EOmusyH2z65quJQ7IefV
9mx7ryI5u2j6NZGNLIFBzHXPHVzHONxKdBVRmY0oE7OrTNiIS//6EyXf9b1X+7m8
wk7dOgXi0L1n0+haVPEDnPnaB9vOX0cl+zP1rnzsYdj8yYHDU4p0y06OrS//JXPI
unYmhcWX9525p95dM9LDJlQVSrmH/wBOX2jI6Qz3mJE97UGPTkqNUMJK/SdyVaca
UYPhWm1p3mKJVIxBwqbdFZVx4vmLU/h5rnIiGdLGeUHpizXLjxvyHcqZ7p44J1XF
EKEY6/NdH0FdO4C0JIzGNvrvepd2XlO1Cmys02iraA8SgATWo1H9i+xcz9iosQCS
yPutj3HL78n9GBosGHjCYEO/yn9aJRWajf/dFMG9dHzrlfxz/qBm0XKmjBWSbAc7
HjE3tg+3FsBqa6WRR0RtJV3vlomwADiT58zWSjIMSeSORyORkjqIz0ge2XQErgG7
6hiMqifOuzkXDSzxwmq6XutwMxCMzJn0geIUwOgCalUL2Mo8hM4vd/ZvUyz1MfmJ
NuYWH/uD2yHmOrhiXBZXt9f4FbABjZ2U03LrtSj8gVBVqmafnTxKJ0QyFJJVMVi4
XhqkwNXFXW0LhzLicheT+unfFUeSuCbCO+OwIrz540l3Y7D6UiGX8dF9ZpUIEBTx
18vwVwzBMr2JWv7CvKJVCZvqny01rbME7IYUn0wviyZwZUCyubOwyoHXxOfk1ljR
Gjte1IIEV73yHpM13aW1rFg5cMfH0p/zxzptUpyptH6b3zq6holddR0Q+j4oowrU
qM+pxuqe+xtwu8Wf1y+b4eg+2n3VPUuBg2Tli86KbnttShURPsWNatInLsiCPtCq
1VXAcJr89CoNHF3+c1XVPnczM7J9pLzwyrhr33XLFO2PDlnb5Mb6QwbbqZJF3+gY
qRwmahZfJ7XHEAO1AVOGtphm8GJ7JD6TvK8liP3fJ6Y2N+mrQB55fv2nKp+5s9F/
Wi3o2a8FJVp+qRW3K9WWCHgzaBcxAnaXGZzH07ooTeI7AMYae6/sdC4v61OUY7FI
0PLnBH9GeN6yUu3VN03XkFs9DWYPuT+JOOIkZDB3LIIKh93YR93WKIb8CqzeFrPO
+yGWjD1V2ml8KeF3aO1B030vV56XyBchneENAv1m6NZv/jR2urC5vU1iIwjmwch+
ehNPWClPuOgPr5Wi4hAV4ek+RujvtLp5UwBlNFoZc6ZN0AHg3zumzq9CmW+SRpx8
EYuMcX/YeM1iXwQshPeudQAZ7/XLMkOgSAKe41CmL+Y43/ZZ/rMhshGZb1zMwY0u
ZuGggmoFUgpgRxFsJZkzreK8AYzbCb6OKrwnnLk99h6DWnhCpnGaqzUqufD+/tRi
9xLaR+dl6q3cj7T77qq0TazruJWv9XIQbquFQiDi7g2bngbKBc/KKWubjT1EucEw
wY3tny5ZR2mRkpAoRoDB8wZ9lB5AqZn7OBzYMB7KdQ/a6dxQK5S7XRMMC1oLFAYB
2k5NyuWyDJ+/AP6LPocWB11aa8Xe+J5CB899Wtw+cKwi2jWMgWruMOIRMOoSjrE5
TfGQZMGJqaXTJDencWekoouy3WH6lo27gbzuIGb0kzilJDbU1Ms9UVuYffvBazL6
fxPj9hDeSOsIHMmUH+iKL3yZuQj88OOJ2iXGxIUASPmG6xPJ3e8WcO0n+v6+eoav
jWXt3YIawUIP1Sxn0ADI0FdiUKa4SgnIHf+Os04pKSSD2/RZgS+mQI9vp9xH1Ujd
JBwNUlTPokCD+ZlKCqNmoxcWroikF53l2jsqN+u51V+InbgnZZ8x9UkQkiIAU5Qb
Xq0c86qoYrBRxAo1TLTO7DkdMJIooB6bajcQTlp8bGJs3rIFBNC3RjYId2ncasyC
mAdbfr8NCqJQ3k2yXh8uROc5EKY7HpPylLEy7VDlYX3RKVW9z4NBrjK3rQYqnA2T
m0Ktf4X64TUU77liukrX8Gh7xP/MZzhxOkKSHK0ZlqGf4m/mjUOnYIUWZozUayxo
t7O8cbiWVrkRTyFPEfIjHJAM94ASNuSyK9iemsv8GE3Hne5/DBAjFLn/+PXZxWhP
4aLb/T25dydoEwU1KZ1HiyAmEZANIxrU3Jbu3uH61eLab36AGsJg+iIRYh+JY5A5
NOhvZG7E1SKfdO5qjiKRrQ4F+psuZIDJZ5l99s88PjJ2TZthiS/UEkLP+nxlF0Dr
WLHmy6WQbHAn++kURpcoAfzgbaiq2OpkFfo+3TaHrGI46QOCTf9G+hdZlk6Y8jw7
Dnn143wK7FT00fZgriOcg50GB40PEZbi3ujYyUviLTEirrWFydVcDpmxb1tjwUdZ
IyDhvEfYH70PucmZbwlYld98XnKg7mtwDROGFvsDgRSebzQgKLjuZ3N0kyJUeYGq
PQCs+xP9PfFczEv4ONB5XEPTz9CAu2tFyjwfBhlkN1KW050I2eyA5kXLhCqPRVA+
iX5SCt8sBBhLU4CBGqfiSBvnM+0RxA+eGpOhwGjKY8xUzbqtY/uBjoJe+iFchi+C
mMb5wXPdAaCqGMkKSWYCuN7mtPTerVhyBCu8Q/yB8qjVaegbAIbPdt4zPfdrR1ra
auBxbVofStbx28wUHg8UHEPx3l4MT08wkg1F2J4LNqU0pOsMNUYYgL12Vj0OVkJW
8CSu57GLrOnG5a8JT9LfRFwxdWClAPO+Y0gvXaYxnoc/wwBEVgBIOfNGQrKj+Dxw
SieCJO/7yPv9VUptGwP3w3lGPVb17OKFaLSFNC6qYLydamgox4hCMOpAGzqzIigG
73ajTy0uQieuCQbnQQGrQf44EPA33P63Hq4KCbQqVmGWNKK1hclR8+lUWief74ty
//r0gFxmlRn2T8+WhUOaUeS+INW/GaeL5vV6otgXroDzr6yjc1m8clcitMAEOrD/
K/hBgsFdzWGB66RVkh8uv56jgvomLWnuV+w3+WS0nr/WSxvjbyRqclztnMTneR/j
Xyo5rqWQSV3b1LYirScszBzNrjakItmf4heQbxVx614WFQfwdilnA+gpZDWSqlMe
EZWDSaakIXnMqDMordfxDwlJA152KShd9fPYQsyTscteV1oq8lZES4LbbkqQCstz
j89Qe+1nA2008p/tplmG5Imya59YbVIf5xBksUUSX6dUav7Jtx7mUz2mTCYRrfyt
ku7SGWYx8bjI5ZcNSLq7KRYg1Rq9dl/bNtL3s1gTt/lFE8pjzAtomVyLHn+qRhEt
j1LwFDXq9Pmgel2BKIjQr0WPSetp2aAgFYvutMAEqRb3CGREYDT7kn9DGfLLEowo
C8lJGq4HSkDU7Fii2NcCHxbNJYO6SMYek5bCy6TL9L4hq11tq/W51fDHqk/FpEDV
z067FTDTXQxkjiJAXwwiaePvrGs9hDhr28rMw6M7ISuZVm8PqbUBYL51xuc44Yjr
qQ2YDvIQdWoJAWt+pxYn3I8baww37CTHCh4+KonGw20F59ZriDiADMYHmx2Hr8z7
TYU5/r1OS0lkpr0YyROYJRS7U8AxEZFc9C++raQrX/Wq3ukZjJ1W6pSnQ6MYb0YW
SLHLA//dbk4NOZQS2QwjfLnmuWgOncGubYTayzNwyl+lOvfvEl/YOTYZtIIgC3hy
Yxi6BrMe6PKDtddGxLW9Cvbou+JPm6qb6Mv5aC40SE4c6a/bQgkZ0pA1lA4sRH9O
RGFEpEm614vXWyvQd/unJLkb8B9PUc8f/JAJPqya0dn3KDnefYmE7R+E59+MDvY4
tynfYDA6NmzZLQYcTBIGYUgQa074gs4FbZ5njLcmY9Bkmrq3BLzfn5Fg4RfgCnDi
QxUjDkPYBDC9hjR/7ULx2Vc0iefafQCAlz0wRHedT8AaxvowCCSXLrZKrA3olD/n
BzAjqcawCqLpZzflrEpT33W/tHSH7KX+MGYkRTovc4kdLVzdWg2rqQRYNxpSRc/8
OFQHq7ndmWYLdzsOOLrqQrw5ZKEQ1ZtHHN9karhkujlSScJ6M1sHxWP2cw4E8O2a
ygiXogWGeBFF1IamQR9xTX0tvgK+XFwoAMPRgYiQUaEs0pIEbAzlmUiKCOgqTrSx
Yw5L7yvawUG8K9GWp01AETbgJt+U4alx02NpqVR/R/1PvXDrHf9ofa+1UPtoQQau
dr9ijVydf9tQft1vjVcuRO7Pwhtrufahe5YITCC5f2847pH/xYVxeIplqMYO0lmC
Q2JMJjn6hW/NyXgtA/2LEDzNXlpRBPRVhj/qHVySgyhCFaXBhaSWxQyykkuJAFH7
YZTbuZP0Hqf3gFqbQbS1J11tmrMkYfXwR1BMSlxBHJvVQkZO7xsi5lkqE+LJZkt4
mWnDSYDSrcshXwZAGWE1+7ivY17khZ5WeQiuROHtZpRzg5o6Fwusr8MjwcGVx9Fg
y7Nwi+s9LZBJvAeoefbQsCV82ZRVTiHGwT9dY+AaWQeB9d0zH5tM8SjdnbsBRdn+
kxfmT7J9b35VGVWbw5wRyXJk8bdXgIjIjD5RpwVtuunMOHIB/Foj5f9hU0wDh8P7
xH22RmuqFVcQtgOyjiN45yABcKOAP9d6cZCK87pLUlakr/H01i90mgC8Xj1DQleI
6/2B3TCZ2eWC6horaRG47TZGHSdTU+6kH5lnnGfYj0q0GmFsHhwM9iAU9QqEjppF
ewuReKCWl5EJA8egihiOE96kBnGrEeLTQX5Ts9c3xrYu+huQPVvtpCcKpSyJwCXY
Rl3PVvIjaip8f0pY4S5ZDZRx3U66QmyWA77q/v+A29hEH59lowfni5Oazfj5yP66
WR2toKDXgQ8s2TcgYOQ2VRYEvpZU2/9vVk9RXb6tilXIS7tbXUROuttyo7muDPUH
MA4VlZ8r/lEgFnA9K/dOZwpeOOYisxmfpJ41bpYaZmx6ny0gEneklU3ReVWmjO4r
f9KsOq1jQADjynR10AUoGUDhwJ9a2SotBjs0GNHrpm24FuVgo0ZC2tGFz83+YxTX
DCSylFdoY+jvqdVRHKhw5z9NaiP+1DpRUwMJ7w8j6rLeHAWwxYTD/Ll4AZSMN2LB
5Ly+WazCz2X8iW9gpnqDzYWOoB6hVum73BTViCWBb6IESKzogHg0JISwd1vmg0/f
c9K4sNYfkoCC577wjR8tQ7Qf0OtiURmT54uZPpbmA7llnhxMq7AZ8f6gpTWEEHIY
r1tkKrXKesJOw7PCbPTh0m8A3p6I/AxC2sOSYDSCRLuBqYYcRqn8rQHaZtv84ZvA
S6iZBrG0SkQty1FAiE4i+zBq7hpuT94oylxAyRff2f/jZgZC4GOY4L4s93xcG2JH
n6fIrMB+Hfjzv0Wo4uYUuVdhyBlnZO0oDPAeq24TpGKpRnSTk3stO5LLNJ8HkKeG
NbB3RZN9m6te1wXLk215sMMMEm/eXp4VBLmpOSOaZGoIdvXKO1x9EXfsOCn313ie
OFxMxAhRCnFGoLk6lTY0dvhxCvJeAng0FRql5eaLmMMULt6H6UulUD6PcUG1Rf+3
/jHEW7BTTCNobMGlJ8ChCy/SN8Gi19Xzk/CknhVS2jmPMsuklwRR1Vg/iImS4n8k
R2P0C6pR9Ff9ZHb6n2BO3kZpzk4MGW+RLK1cuMUAYLjxcCwnEXL9MhCgNxDEYYFJ
b0+jMHuZ532lCClS1gdG0k1Ge2BvSicC2Qb3eP2XNPCTdEYSBDA3IVfcUD0v9WQv
DCZIk3JSoQGTelB+1HXSlTk5fpQ5IMjq7L37eG2xOtnpLlN1d2VjV77vZpBSM5qo
k2KP/fYq2/qqLyCMT/Mx740KZj+EFljMIgde0JNz8gBQ3e+CXHBZ/ceb9LpC9CaO
c9h8BQegGY3ESNdSSfxfghyfTso7wWzSTX8EYZqBR377gNZfpnrBs2zVPxZ5AWAX
Q5WCjaAUjcV76FZg+wAH5Lpt/K6NlgN1CWJ8d5u6qkRjfGB8rXn1cYNi6L/m36w/
anokNCjUH0JAwrmlOuMD+8Jp5kAKuHHNIsA2Adi4HdQLGlhdBehkP/H3Wkj0SIhV
lA4xBefYp6i79Qmf9fN8IwMrN6hGK3M98Rt78OkD5ouQ6roX74zsfO30yPvmmn8O
bh9IgFB3j6gxwzMLOUkARGbo/JWvqtEHaEsF1M3RxocOk85lI5Xr9CCb/9dAAGE+
6Zs092NQ63o4aiJFrJ6QuLqri1vvMYrGC1PBvGBj5PQbz6HI/j2OiuppZ0i2N5WW
I7sOsx4tQ/A62aknVRlUeB2H71VKBVmc0XPijZjkkYkKy5Wuqbq1oZARp9zDTeyK
O07+2cqfPgh/M1p/axVNtUsvEdMhGLyRZUSo+4wsu8WHYCFms6trrBTa1Px6+GDP
0xCMVFBA+vqkwUqHEAB+5u4QNB/1u0PLV18kf9ou/1oVJQt8zzZJzl3TG7WuY5AS
IFVZSTe5UAA2zGQCrH+9v+9gcyLyVUdghLJcSl2yPUQEgIJSH5WPzQheXPYcCi2c
pX4MB6qhfZArofVG4jYxZ/3kr1Rb3Rj18wPiESCR7j+bPgWEUCdzmvLn89na4U2e
NDyX0yhE065F17qwq94daZ6JUYhgPCMOvHrjwmbpiqIZO5INXxcJ5UsPX0M3MPAD
jDh9yuihMqOpE40lWFay5fVg6yLETP/VbSzxE4Ugl+kOq+JSl8e46Qc6ukc3oG/X
qyqqtUv1E8EGGEiDZt7WTYUh6YGRE1F4a3t/m54gFC6HjjPQBItlNoSp/eiGNcO2
jTyy73E7SIqnE9NYMjkJPWz5CtDJS8A2FgwOPQ6gT6CJ8pbL14xuAQ4N5zybjHT3
Z5Zf7pctD2VaIwNnvH/SJElAKeBdjhhwVZXCKdwSBT7tYdRw52oqOmfD6DMEPdwp
YGEu+S1jsdyxit+6Tt4G3YcPpZahKkw+keM8ZIh1PIEntTQXt66P7LmVIOoYF78Y
k5QZ0UvbE+0pxdbC07R1xBBfRxfTYXPGdgFmzyit7wQpbgFzPGU0JLz3NAp9b5YJ
ZSeWQOMznk8p1tYjsC/J+FHTWrs5pGC//2Fz9E2V2XZa5TT6gijysv+FNbnoujHa
Vr7aSArtEdB2xgF1Y8L5uf2PvN6I1yWO4JZLonBJr679/mWe9JNvfaNrZ2EkMlfY
PbQMS75sPW7vjTVvJfbhw/fkAsAt0et2NewVCRrX6zji8ZATIc4yXJyCMkfj/W0M
2Srph9oX0ic9MGMOMJuzgGOrJ+2gYtzMvp+PcCwoOY7ut5+bT6swBayReh0xY2kv
LRAq8gCQmjEV7052aKzRpsyuJVsX9rrTJVuROT93fNzt0mZuyyX7rmWETCXaJ8Lo
/JX2xp/JgGbLbshpG5oY0h/OK99VMEwxYcgNo4xPXJ7PIyzBk7TOzkBNRSOCzmT/
dN62cA21AU8vCUYRz9hZoFWuzf6dNDzyKP1KP2ebi/aPbb84R5VuVWbEaouJeDP1
VSY89V+5gpzTXvmZ55YOVSQPBA3IchUcs7FVQbpvIL9ylnzje86KuOPRA8mynUGA
71BE0tOs0WDY6gZH+wXyMiCtJ/aGzZ38zPswhYz0qJNauNY/qZqkkY/BS4YOYDfz
OncuYwVIMYCE0+AobW1rN1xWvb82JP8KigwjSf/zR9H7r2yJJCuK+bmhm0FRnf9f
BRawHBfvEXKm2d1zmoroadcSZ92ThdalGebVP1Khycqnf/MMci+yKoLss6YEiev5
VhOSNrqvTMQYYQIw9yQiwTjbyrb1fSYzd6+dy0wYVJyV2bImJW70E8JPU4n+jyNX
KUlHOGbwDxX36neFb64S+uNr0kQLmagH7BbUQ9Gg8W+oWVZOaqbU2cJaa2Dx3krH
G3Dk5jejCq/8Q4BPuKDoTE/xZUlwbyBBTX5Be04hqoz+f8ExlphyyY+Vu37jOXZi
88xgjrlLOvQHCuGuTDhsOVBvNqyyBQyvXbbSYfXAyI73ZmLG/7CsNSwjHscX/jex
ZL9M6kRdvKroG+/W2hTm3OYAk0UXzbDwKzu1U19D2Sa5+hExLtEuWwG5Kn+Nvv11
vwy5KtgTlYi4zx3wWJ6yObLLYFTEYLDk47LAYESsFdqdgKJcMjSNhMI8nka7BakM
ZzMZ4sCRNgJOJULyx8iGypln6+YElI8aFlwch+1xS8oOKRqi73/wzIbnnsGGNQ2o
a4zVinUtQzrBO+6QKOCMT6JMf7pRo35ldfPNRATxsnJ1snFc0NiqkvT9XGHcris/
VKiNhHQVlSYykKmkzMUUcs2j2SzYNKIcGN5bRp73sqn+yj9xD6oqGraueSpevy0g
ZSpu6vV2cLqLk7rtz9nizYyhfhAUW9rOkVaYDU7L/U+w2e9+zk8hAECxYTR+b/AV
vbVA7eUmITT/jDcrgjhadRe/qtCd+BmQqJoiBQ5XMcgnlEX/B6jXCA1ktZayCl13
MZHIDnj5j4rP/LqJkqTqtXH0q75Vs3BjM/qI/qK383qrvF4D7YEwGnWMdMNbNNpm
xkWzvEYJUTc0y1v8tzdJ0ZIkKbWt4oVFcLqQElG+zGead/GFtZgvOyyojs9V4En+
alBvFn3aRayhldiEXPz9fSvZQSJYwPp1QmE3BbgnFSs6Eep2lcPd5eIH4zeREhxY
zDju+SzUN1WHzOFgjxYwt/HQF6TNPCsGwbaaO13UzL5sq5PHtpcl47bazh+ut+pI
tM1c8MlauV6+BPRIncIg52Lbju8/lncLtRK2+Pxkc9tYuXrzaY4AfHSfkB4gdtlc
6f6ya+m2PMg9WGVlFOAoIVoh78nZOjY95mEVNqOEn5f2NDU1nT9UW4C4AyfpT3nc
C7iI4CJOpnATe+7lhQowOfvXoaPeY6MfbEDrcQSmJYYtS6TZ1kfrR/nuHLX6SLog
hTlarShk7r+8HKAv1pzMyM6U/v7kXYaYDwY5xiyPzCGnJBoCMl6HalfZCdhkkbd8
i74j9IE7LjRNIYUZ/Lw346TBZ5g/y8IaFb4YIrysC9kXp4SNavTrg/9KhlWOTMSX
01VBO+fzrSTIWfYSeYcc/gwASqKzrDLWW7mDV2mOJB7vQgIcxtSy7OW7YTDA041z
MZCRzxs+EuMVE3d7Qqs5U+cAOl673dSy3tLz4BWMNXne+WawHgyWrnf9oUo93UH5
8Pfj62s73hzEXapGBukBu04Xl5Z4DSc0pnBBrJd8/3rkCAb2usuPy/NfbV6tHwH8
QuEBEqU7i8SSXoJdsLCb+fas6GcBVS8mfRlJe6zuIBbyZmXKnGK1Af+bBAujpkfr
y8mBOLNb2hQ9eiH5bYHObOWh4h96IjygBT09701QC6TqTUUp6p5cjKNYiPDnz5Bw
uVFzhN+eVCwFMdivc/Dnep7HlOU+3khXpj3i/MbcRIPuYDNmGVcpWbbanH9wrY3D
6Ry51W1IeTbmmSFJPBGVcJn8B7gWXMxi02wGPRMk2ZhQQAMBfiNLmsrfgPc5rT2m
CDolk8VFE+D2Di7rvEG3PNQlT9Ylu/PspZb04uvFCmlKrEipZGnDopUIctZMObVV
VH5s9Gvcw4NetpAzjZyqVlJCQSk8ITk4nnkbqWkI9MPAswKyBJkpihePyVwD4ftP
K2mAU/RwuWrjyGRB+0oGHexgfNDYn2KxaLQHnCJF+OvsJgCLh5B2C9kpzm5OnjnF
c59CsQ2UQuso/qVVcn/kA724RcbC2TAODkXpqEsWAzXcFMcW7wM0O+rKTnUWoUpv
YX/WwjoswaP1BteFrcWsKbmKmPw7qxf/T+mmkoiTDPk8d+xpl5R9QB53dk8Mt81i
/Wf9e89MLkqAiu/fl1RrHmFR+1jNPSyMEhU3u7/84xe8+6iHihK35XsnTz66RKLC
S5x3vrqvk67jQ87mhuNnU2rSGlxLTe4pKjEJmPzUul4ummja91F9o/wZB7S2jG9x
rQ22iK5h31aJpyqJS6Du4ZGAq4faRRMkGt4fPiPbuh0R1pu4ti/q3OwhCLHiv7jS
HbIjW5Og13z9F4gzFti2fp2VSwE570TnaD4tTNbayrR7kkWKzX6AQwGh5JWsosIi
9lJ1rqKf2IwbdjyDeGTgDBXDjZ+1xhFsd7us7U5Ip34YAPP0GW0FVZT/OnQZsVbz
q6M3DHIsueniiiQ+FETdLGN9jSx1ZTe1uscR0e8GgoJCJAt90VmNQXx8Y2mt4RDw
d/letdYkVRH8srTLIdlhQwG7oBnQYsNc0AFS8Y/bnHySmzkP3/yCkhmrZhcbL7sn
zzi7a1qZH2FGqbUwRRqAJ2/xt7ieNDPUGf9PnomX3+yb6/1ibXYEr3xJkLt+COtC
t4ZJXShbbUAzwFhK9x1dmHRX5XqVNMrW4j6IMAx7ez8UW8hoElh/S9/1utY3lJ7n
CJBgkcxgWckLV9qti9SmusBhWoTDRrbaU24QtL4YwOStRzIiajPzQklEnS9RR4CB
PFpKEULbi3TpvD6QoYnVMrKA7ENPxlvjfx20D++14rLNG6EzmqtKkQNRW9jzLjDk
fkzSDY2kql6GFMeOuE0uj+zYr+QDGsuBlClhjh1XcfpqvtYQfaUh1viq+5NakOFq
tnxZwFT0in6pvWLmORu7LK7jggFIHwmD/X/Wa7I6Jjvl2em+2lRN5jl9BrmtBO5z
F/QoVDtRXryzCa9sL1j+fIl6Nl849G2+EV6AbVHLJrWR/3NHJwPe/IoFV9YAPSwB
A4qHgcl+Tb8GhM9zzH4Z3f8FpBnZ2+6eb8Z9C60/Q0vKEAo/fiNYWZArblZ/NEQR
8cOPZcZpFe5Q17DaCgrXgP2P98Qgu/9J2p3qHBdXNBydEmRMvmRaTNXGq7wzorKI
TXrp4R7QLuU4Gwl+qJR8o3Dn7Qo14vaaLJ4IFt0ylHLCHQp49zSZoA9WqC3oloUY
vvQCnOUvnHvX+QLinrOIIUOegZJhDaZjHxM6KEBQuIQUKUynonNBm428n3tReZQM
Dy62lcOL0Z3ynnEMqXdB8jc6vygQlx82TAU9Nm8aa72ssRTijPHMuNGpV2Ql5I+r
a+L7ctqqkPHm/krhIDg/w51HkF4TZzEsErKuZBBLBZ/e+HHl3CwNjPsH6bIDk6Ae
t6i2t5QHTXD5FYP9KWtsy3cd7oNOE9wk3vh8A5gukHPSxHIS7XlDJBc//x7oyKPJ
TZh23NXBgu9trKVktuTVJaywRvz1wa/A7MZ7PSUKDI1be7gekDNm+j0T6FLQMDSO
v9/HCY8/0a19XFGFHAiXg3WC68cw7CZII0jpqlu2eXi+e7YGOp+FzII028FAwn8Q
7L4uvNp1nX1f4HqO3P2uxgStQAgZrW5VyK5gqit/d4P3f1VRQ/ZlVh7z4+Ws/MBc
Ba/iBYarxiM1mQB6mJafmRUz1Jw8ZGVJu91+GubFuSBsmtMBgfHv/BmDYzk1Km/F
1PrNNN0eZJPsQ5wJdVgvCd0ds0VKV6s8jC2yKDCTZpa4MZNOm0lmwXsCZ3vE/wYf
+XEGZjcl4Pj46dsBAelo6njYCgzxjXpE+jlQocohIjsJ8etzQhV5orMCN4PrW7XJ
0pgyIK/tcvnKLYIwUAL9mClc27ievfEEQ4U2u9Bt2IgLpgLTa46bltZQqJtLxZDb
v945JwQv9QOagHOsi7TngBJhdK1wPkahz6f3rLJZ02hE/uwCwwkWfgewc3VkLkuG
NSnT2So/LNMfjsLCdCdPQP8+bR0tpJILj2QlBTec9sdj2XGw+8AMax+jLMDRazSS
Znb67JlCvD0uepY+mKFsM25RwF+hRYKXQszCrGaReRuYtkiVaYfNXw2Z3Jl/FsXI
soKi33QtmHI+/YWbnBRKPVxVpvs6XQ08vKeejcqIN+BJrscaxT6PAceeV/PGsJBS
ro30vm7RzW9Lfhoug0W7kqNX+SoUyPtqQ75JOTohateeFJ7Hr61i9+tQhINatoM4
bheMp/ILw/gfaGEqOxhs8mMfFDM94nG1q2u9cYe4I0dzKjhmFZ1BPK3vKa1s0eGk
IOU7PiMEltNlZmkkIXY7TQtav1+dorirqNA8TlBSv1cyiAGo+n5DZFCh3e+yvEW7
LYAjoHD7abgqcW1iDMIosb513jtBNpAvEpql2zKX059Y3f9D0jeTeUe1wPUgncUx
FVg0o+iMv8m2miEnozYyyTPQKOiz4B/7sgC5NSMMEYk+xAvP0VfEQq8UZav3DlqK
6wiHZs/hMSTwJwBboHPownOaNVWnGbubMdM0i9P97LXNhk9p38J+tBCTP69E3gjy
y8BYsfqxDZPci8ozgi5ijI+81RlK2yw1FDbEjt1YtLK9lwap+VEcNcgUhJousr6x
BuseR/eOc5M5RLZBIRr2wk+Ck8Fh2ALKmlVsKTvYovkiB3UPE25fUqkRKPOxxs4m
CvGNWwmTZ/SADMMnhSQMnBEOIBYz65IGsVDFBWAJ+IERFxri/+R+BL1ImEMRUaj7
ldSo6Is3ponmZBu1LkyuVQbUSbGr5bcP69k3jSHnUvc/EjoWx40XOEhcr+pwzqp6
qZjHz1W5gxPKZDLxrhL2RmYtDUWvlPX3jPLLiS3Po6a8+RP9t8Ge3JfO+vnN5Q6Q
lYxNyq08vXHZRgzTtFrV0yC7yjEWB6EFGmBoZ1gT71E/Q+AF4dQrwJSm2+IlpdnH
+nZTMLbp1GMmPBzo8kx+Jm3S9koA+bP0Pcfey8eXSUGLXlffge8oo3rkIkFFqKl7
fCdfP4hVr5fWEfGkDEaxWpOWZ7vc4nMzHgT3QoOIoSZzGOklnM36K1ZfdWeJw7YQ
tFWCCk7P8mzXj+NCvB3vl/6NjGPTEbujXhSNGvBlyzzXgux35ETmP8h0+HrSK85k
uX95bVKTu/tPD7ke5Wvw6OP9sftYBhw0Xr8IwwRGFEfUCSKcO8T15bfLxUDnATph
JKk+E8A5MWeH2YxmpiJ+bD8baJMOFiSdwIwM9WyTs3wUvrxtiyfvVuxiLIME9bGI
ff6Xwu2fn90mmZquWtalGiBbl7li402mO/OsrMcifF41++kGwPRmcJeWTvovHj+5
ellwVmuLegqYD5L/XvO0Z57PI73slUsVgyi7DtmDboJ+S0dA33kdV28/NR+qPcYM
u+RDP9I3nbi5AZpNS1HUQlc0U5qJ5aBgxzyouYLslfuOCjwNNouvT0d78Qvp0D9A
z8Xd2obXqJyEMTmQhTqKV1fBgD7dxiIXES+Ve3YS4nt9L4NX3tjFn2lY/1h7ivoe
/kktHvfi/M1pDaaWFYWb1tl+IFwQGfyr+J2bLYd2GMGDuB4LTY6JEYIH5FWLr2yI
TqA2T0m+8Dm8+UIp8tYyL/YSyOiwdUcvYtYL+oDM/1fk4nkBBKUTP4uw8okmA4d/
8NXoetP0KsiHbo/NNnhd+j13sHGTjntQP37UPoApnwlZeugM8UgOM87UsTnXpOyG
/nsEmIypWJAyyWjSmTSSsFyEZajegm3cbsz3vgphB1SpuzhDuE53/TTMsLmgjDb/
uKWmsTkiWam1EgC2NiaQgS4Z18C/QqobZVi/xnYhxMSH8KrSnbYvo4ml0QMyzrvJ
GKCPKI4pnl2tZPZCkijkUitShbQGlKd3dWq3SW7ziNemxhBcVGCLtd3+nr1W1Fwp
iOedMIkPCUBBDDAgQS/gFaZkUhWwDGDF0U5oH/InaLPadmiusoRtp0bj9q5g7Fag
VX/nHO64XKvhj+jRlUbuRB2fs5esMj5gJs5Qg9o73tV6t3GFfILBOCoWutaxZB04
DbjeW/GUFhdr9mMD8h5ccwrSkaXt5DFx0X6+Yha/AZhHnqjI+LYGeWri9hyMSf78
09Wks1fyHWH4GT8vq/FJxkuuf628FJ1OB4/3BPBd7fGdoCowD7Uxu5zQ9JkM3s7v
JA4kIhD8O/aGSaNyRUBwcLt0avLthjfgPKwc/zLv2o+Sl/Cxqc18ybFWKEcnpg6H
gB6pETfG4Ji0vrtFt3xb7qrPv/pWME9C8TxDi7phiCVCSvChmeHi5NefxPd0MtmS
WlFJtyT+aBJR9yiQjaZp3s6t5PueYNXUVKeRdXmmvbmfF5A5fg5u+TI9ZChCKLnR
vLpwbf083mbQg4M7/0+lBQu/G2v+BKyI4ZAmV0rSnOPm2G5gA9mDtz/jAKBx/myl
8RkBaXDtvfxh1AJcWgUdbQC3M0j9ZJWozP9zCIEJiyapXyy6IVPT9YO6eCWwz59V
94XPKF+vK+cTuqr5Wmw0uu7VfEzd93a69zsnQPwWay4K34MUuaV3SZQCaSFihnVz
LhtNr0lC4pqLB6aUP/Hpj7oSccx2TYUIE79+3PUgFa67E4gQMY4HCv7Qc6r5Sku4
z8pytMcVzNY7BbJs+/6h416lhoKEz1l8epLbSIB7X75/70yytsD2l9Uhr3tll2sg
xOzfS8aZTAkzpRNe+dd+U9XADg9HP8rqtqiMxz/6b1/innDl95dhDySQwSmArxuR
HWkXv56xWdsmr9ohvH05quEOpckQEwo3DDD0alzGrtvfTs+pse7oe2QSWsBoQCe6
/fdR+l1vBpOzHVHOVqm6LRR/YtyopTpAr6CBeX7/fzf/eD23QWaRpndWOOlPFU46
B0d7SrA/Q2Ylu9wpbi3I71pDpPOGbeu+Lu/uHplX+MUp7Jy4RblghZ1z134HW8zp
70vVmq3FntMkIcsPYWQfx1UZqunRsnotb97uJik6hJVZ1G+OqDFNbpN7E9cEnzQs
jHFtrT7yle9aYUiJZt8HwjJEzoefVCjlG2umFXRlQeunYQoXmy5PeOZM+B8bUDtU
faCiPcJp0ylDJQc0KrdecQrmz4ytfNp1RdF/BU5nGCI857GkUuvywAIT2ZQrinGb
WAnv4rXnPyGJjTj2rQU4zJvWHhplku9eAkXTvCnALcYUIW1HlV5V4+qZch5B/1ZJ
dI6RvSlX2t6WGA8YT/CJFgAg+M50GLe3TwN0fv4j7RtlQBzZ66zKtbveusJjlxJs
rhAfe0+BIkYAAuutlGFuZVc5CDwax7NwyofjPEq+7oQcrIxJ2/gHwGOpXDipr1aj
M2ru9BxCDQw6JNVYUnd9PscFjwC9gHSs0DeOtaIL0E9Y+lH1AX8TQFsdMlQu7FW0
+hGDnGOXmJT6R4OndINxSrhlJnel9z25Jq9zOoQDz2I4Tng6h0UGPFDrqq2Utfcp
j4FUD68gDGblDvtT75CvnRV35OGZdSKVnopJjrrTdvsrMQEESiWwnx14RpIaBsg5
UR7GUE52sNj6iMcHKOoRALGCeUEgx15wxsYUWm0vfFGwWDX5mo3HpAt2K3oSBjSC
xb5a424YZkK5lYnNZsvrh6pySx1s9WLtiCXmVVE1UxBtoI+tSn/aIswvmTsitvne
lsIGrjred5cznaGbb5H72Xm08/jlflfmjf/KUA99FZq1Mnla3GVLkFE6sJ+LudG8
u6Ejn/d1MFzBm6jlAJvg2Ctcsn//2mJ3g/GIcvqJzYYMHVPevFUQWawEQJgOwM0X
H3HAY7y9f166Dr+0RJfJF+1NrxwtbSBNj0UtpJIaW4qHSSCjx2DSWRbcYNkkuh74
84slbTxbDCAsMyX0Oey6HuxMPH3dMp2O2/mMUhwtFbTLwqZQ8rtZUSOzADEf/mBp
xmjLosUf0AJXT+UmdjJ0z9luT7zilypiFZQ+lG7JDHGqrL9koNXI9iSUBIo4Bm35
kybdc5bgJ6gpviTql1NaLj9jpaXkwBpFljQbiufB+TIONKAf3N1WKhQ4IWll4gNs
jyKqwqZPRdmw76eafow6UFWfWh/TmZsNRlRwhBugUQtjvkd9s2HLmJSDVQRbF5e9
kw5ovBst+W6BFdoXEx5wytOf2iv5XmHxqY0KAyEKSaw/wrO+s4i4PJ/adNbhCTNT
/kq/KQa6clIWL6fhU6GPt3onVaWnOIhXQWqh4P9dj4gX6nVvDSey16UH1TN3b/RN
IaoBbXUUEbdJSKIVrwg3qttzi7zXwTGKJXv34iMydQA59CzQB9WJya9oTpTk22iS
EraWW83iywLrAAW91MgjDZJzCoGU55voyR1CDahXXd7MrVDyQY1q600ipenzDMwP
XqN2gE1KbHgl/ltn2y1Fu1AmvrPmmTtoPymGowdscyICn7b0UnuzlmK298NRGSr3
fnLbFMQhgSfBCAW4wS8JXWkBGHxVM4EqSIRzGHiVht96ucwQXgfBl5TqGEt6CjPy
ZrPe1lF+U04x5/ifvPuTIHgVf31axUIflVARVhh6JaXqstKRC9LhrpRSd6ifc1Ig
Ka/s3DkMwsXnpAOthD+qJyUr9gHFerQ062YF7+TdaiCKyhGVOH/5zygdGSTxPu/G
jJe/ZiJn5u/9/dXAlc2YxPQ8QjL4BHaCRyeVJZ3szXk1JtWQr9DW34lnXTDtxKU4
AGPc0zMfnsPtki7LSZySv3sH1S+G5XF9csFdxarhxMbBl5/yBXerB5OTuKijWlej
QjvBnt8C5LywCUu3kyq1gI9JvbWuOUtfRLOjJYx2Lr2vT+yi3O6wcE2mmD+XbxNP
1kylcDL0m3Xz1dpEPx8xFfNnxQX+yBIBvvV3x2YUOP0lzPBOkb04/K8yVkdRITRA
ONu0lrg+1cccK62R3RKnIMcg9D/Hz9CzRAUckGM/+XtBUv+Wk3KVlDvhh1tiM0H5
Q5qqDiyY+v/SSXfL4FTT1WY9zJCoBCf81PQA5nXtZW8LaeuZDA9hLR59Y3CebW9Z
pK6WICT4QBx6+dkBbPGvNXH1GSbTj0lxKu5Ema+7sPQP8M3Ke8w7v5btHeANl92F
/Ikb1oc1PNNFqKIRb0MV+yRB6yr8g7yiAs0HpX59BpNV+ZhIVRS6u3MW6eX2RGWp
+TA1vuGPp9HUfVj7yWkaNFVbqGG4ZA1yEinXHJB4AnUMnacqOD3i4yWAY0pN1ihm
cdjJwG3lZnRGwUlB3v0Cex2YRw99q+QrXwIELY+iY18fTwLe3j8fuz8svRx7F6LL
aPiJBqPKwZbcYz/nvwy/xSO2JxWLsumWThV9+y2HV7OdFzG3sszXHJJ9GhI7nG7A
+Dh0JK0nFx2ATVcrS8kYmcWmkKGwUT6UBXse5FM+S6RahRNxvgovfaybDefDYRRf
ZneG5uiD/R8UqVHVOk+vS+9Jg9U/VMwb38uV2LF8/VEgix7Jc6LRjzG1IXSiyBZY
s+BZklJA5l67DMELRdPN/AtaMFH7LInKYjvv+r1b3lLXI9YUCjKIJKz3G09MZpxu
206AScN2ZbW4q6poucZk43xU6B8dmwnEryOp7/gI0NeG4hEdSUGnV4UTU7H26gdB
hB87ySXk0tEqnBHGziYUqSdONK497FkfAzj9NPgPg3zNebV8wx6opvfcxbG2iKz5
mFJuNpUKcQ37oRzBF8lRX9KsSsd9ie3Q99IwTKkjPrgXVOH0dOKqzDrLzK/2VfZb
yZsThyIVuMK8SEmoiDRnftBsuKyLTXLryu4hB2Xg8V7553BUHmDie4xlFeQn7hZV
BUW7HdMWn0frQ+kgzJY5jETsM2XHNSQoiBJgVIjQuc2Beol4xZAYBvleRNSUpVCT
Ojx2rOewd9JmSyQPSXCPn0SCCo/sSaNbSdYG/bJTq3WR0tM5ZsSiS/26euDEQPx0
orx6y3Q6xg7U+VwGlbn9hJ3A4KtPs8C/jynkiBhu4YzpfJyqMlfsVsxjPEUk7lJy
YfslMyRK/ae2T0B+cjfGPjcIMI7pAlezNxxdrWfqS9hS/x4mYsGS2NpYJX9f1tXs
++DJnclZClMM73kn5m5TlyaX50Dw0Yg/uZZ8rqbgbgvpe/+K53ZXgrw9dyaPt83Z
gmTEzfD8zo7tDR9Grhf/mpQOsBH1kttIzTHzl0X+f9NVXPlF08MQ9Obadh10QvL9
wBp8GRDKnluaQfwqHSBQHnIQ788MAgC6AhjhoqHaQvvUAZY/noKhGv08xTDLmvoe
mfC60J4v8D5+nd21rD3X++0avl2rlih2JLYyhZZokckycqFS0L/NIKjaX+ja2EmV
8H5ZjIMLrfhxKVKYYmPmyUJ+ki3l+LPMBwoffoKkZppiFEmWlRlo0eFBVuIB8qQS
yY08jG9d9AOi/WvRfz+ZYvg3tKNburBnnDXFbDzeNVG8pX515YRk7Z0ihTWQG/bw
97Gp7akhTncCryr2qOYJaMvmmho0Ik13IexhMyJNOEb72bus/jU3NV0rKnS8Th1s
abVArw8Y82ZkxggwGTHxv7zJH17OKPd0rxOpzz0iW7sAAO4B/+WbG3pg4CfldC4f
+rvrCH2m4W7ETk9oV26BgHG0m8ySNtAGMr7WurXzM2kl7bykorkQ7Ye+YlBhpoOS
bzclpLAoF4T1JjB8ZdNVEnLm1y/xl8E/UlyQh40lAW+keD+HCjreznD2sdyuKuFp
rlgOCtAugK7jeofiB5YJ0E0t4xaeQFDeEAJWMbx+XWCOnuAPMxKgdl19x+vE4Xi9
7jOhUi180Rbo85LpCRwTOBsCxHFAmaUSQcdElerSN8HyTtF8AHe7MBe/wZnIbFxC
C3rZzsmDjH4bVQDBus5ltTOoFm0DunSl/hGTV0j9SPWaYPwxEfTBOp03Aphlm1ZX
1iAmGOlbOvWKn/CjX+nYfiG3G55EE/gIUEDKhZ31V84NJGQHflZitIFbOD1uksNq
emxXoQ7tplyRw28eLnerMnHg2ykjTBB4u4rQRwFY4vZG/33uMoDeSIO+6+xXBxsi
fcNukkqkAQ9h0a8hOtlfRPIcvTpUX9FOqWFqjxhrYkiyxbWqzQQXneoCRtZFpxE3
pJFabtgu3Uz99AGjjMIG9vTsVl/AxV8rY7tvxoSW0TR5dzfgpWF3SmfRBF4O6nsw
7mGKQoOkYA9Kqwpx72w5TLtI8I0THERW854b+swMHOr9dTv2Q3wHFmTWFShxWfeB
tztgPU7OfRFMvSSeK845laTdd3hoK47ZFLmcYK0P/caBn5ziD7KIiYFoy05iX6eS
QDM2yLZJOXOZyNf5dfqNwdgGg2G/QjgOZ5rGqKGou/4qz8ymD2TJwbBGZmG8qM4q
Wgy/McOHYKdM73iOHtryv4z/AbAVWmSaobj7DvLSF3JPiafqSl1eyA8kjM0awLbh
MpvZLymq2GevpzH3LfT+dG6KL7hUngWGZ3kUarlzM9vria+278DbbrkH4PxMh/H9
Z1vHeUbeV2kI4QVscFuQ2w2ImvD2VFG0ojGZbiR1CHu5qEn06KYGwaGSqDOP2UbT
J2/v6U16HVr1WqlEY0yyXRlyizzjE3eu2s9VISU4fvn8IWjQHhHJMaqG2qNGaxVW
1N+BcdoJrkRIfMpzdCRBCEFs52eksOp+x2cgOlvkem0sUJ6UWCDA8GicexE8m+IK
EcQWfgaEns0jWSbOGe94YqHvK9DGEBas7y/l3mwicNfnwQtf6TxSy4PGNuII3kjX
9G4hjgDBJbDwUW7c+PnHepG5WINsIoph2V7VfNETLUbjj4m1iaTX1T2Ly7jFDrbD
gB10+7WrBPx42Aj9wOF6/CsJyUXwrKBosOwjFf8ufulmpIZJVSYrJc+4YERPWj6N
VvHua9YHfbIHQucuxhRs684NKUdH2sMmljpffXt9cem34kV5IS8kFi7RuWNC7WP4
KIoLSzHYMhAlsR4jDhYHa0R71uh/FLwlUF4Gwdn/gJqeuj1z9Yw2vFmvafzxZeki
bkqqO9vy/G0Fweos+fNILJveFvL62r2zDqh8V/eIUH+IYUQACNq8U9sNxKQ6r0hR
yCjvxkwwi6kyqB9l/yN++cmHDt4F9h5kTMu7U9Rng5IA8wLjgPPMqTaBBRFldW91
aikhYuy4xd/rybNPMV531SlisFRj//Ao+AWSIbR2vziZkm06fDiOwENjSv7eJQPE
/y9jrUSXtj2WzSMSy6ZPWJK4ivsW5GA/vTh4pzOc/3ynAwZs7SBpVs7NA8BzvvHE
1fiKQ78EvD5bx1iIONYdLbHV9vID7MmgfjqeeY7ILEFnvbkK4RryQtuSUUuPjU8R
ojTT1p6SurA63Y4CowfrkDcIAbc0KobKrNemXraxyQRvuZp/ixJoP5ylEVRxrGgu
h0XnTmYEm4uhyvHG14jNlHJ6UZyGx2nvQU1uEibW7QchDzS1SZhhLWc7fjKANl3M
cwTA1NWuuPpYDCOYGxAr+yjr7z0lBROO04zVt44o31WdQSSKh1DRdjEaQRicr9yB
XaP/ZRo4XrsohhxFO5f78IMXUVg2Gejpg0UL5LrwwqGUGZCHaDaitu5LGZdR4TGg
3b4raZJyC9HBQYIIJYWcaipJqs7ld/4OXNenMhBsNEIQlAPpESFZxb10iuuoo3zz
h9nCjFJG6Hw+yTTgH0VB/njVtSOdYFOr8/67hLz9203K86vjSWfhTCzS00F42X/S
9sr5Ks712MewM9rQopZn/0fkKbAxVYztYI9yY3dO0VT7UHFK6syXUIbbGWdE5Eb+
OmSOjKSsDoCIZWIBCGGDGTxJupy/po7n0xxSFBoK43BiKN6x6PVLZGpJmMMv6Fv/
xdccrRCawk6gTDS1N76eLcj379SJe+u1HZJXaqrH0xnd2EwIwtf4dRoQsoB2AUqH
AXBJ5AF+sNBtMNS9lEu5zB8yz6q6P3vEkOTGY9NExOLO91fnKzr+Si5/LS7wpH5N
xxM2I27Y1TwtP9LZUeerCOBJBIDa4Hd0UAol8tSLPTmM6ZGdjNGn3Y6Bmat9tvvJ
BDPVE1UIqBcTu2yqM91CQoFccOHGSgrJ6LXjduSMaQeH95Ujktxqtn5Ax6UzbF8d
rztM0N5ckRjjcX6tZI05k6gZTaArmzPi0weUe2fleAGBP6WzYtFejInBcIjbUWgN
8ZQI/fEUCU6P+cKgsSXjuQlxFBoc/6jFlsNQ2FRpWKpkAC0vyPV9K9VZPpUSMfvn
ncpMHpWeTvfWNF878UORy6VR6uzlVBQiZXcq8wa/wprNQub2jFUV1E25t1CwSqiK
+OEE8HUS5XGOdP/nD0PMnHco+q/7uG12AMtw7SsAAalpjelZeJVx0Y53kUZOpXfN
AWHHHPOqBMqLHc1FFvEEI74p/PHrT8kBwf/zBVdJhWMEXUG2TBaENjwoaFsgasey
ZNNiORw7vf6BhAMsZbAEdujdzFcCjjMo137IUGCS8NcRe4PDyU6pP6TkL1cwtxaO
EmnVkQkqRMzfDq83dOZk57DJICVDPeJ5Iq17l984PJFELA2qfF8VexkgKBNTLiXu
JNZvu3rsynC8Z2XSv441H+6FWb6LHNPeWyy7S9N0wX6VDw69ApRJ9t84hg+7XC3N
JpLC4gMq2X6sPoZNGgYGvVfcPrnmIt7Wvy3GPS6yZZEchaNMI3HMHj1Zei8Zre5K
3Z8Y8fPVuot/Jpkfjw0BECiSOSIme9guj0yUyJVJkpOHQRUUnj3nai5BuhUivz8I
b6TNQnajNLNE48ss98rhGZJi9ukAtOGkgF88LJXmEBgcg1yl63zcZwwyRPKuYAkU
DHgi9E8/eoUGXYa+JmGE6yNHcXrhbjDumqsH+7m0MTN2fbRj/xtv79Jf8r3DRlgy
42EJcPZqEegnc0Jrs+AK6Oeg+WlWB+uu7c2AR3EftVj6GfhgWwr5szj7KNRaXcVH
qZU5U/qQcIbEbEu1ScuyH8iM9bKPRtnscfOEIDHVwY+GbulRzpBiFn2dvFKPcmDT
7u2JkzKjOxcKmnlNHkyHDI1XUJ58KFVJsYTs4uzPcoy7ccISsxsnMun4aqvfPZvB
OQvXxti59UqcCEMvo3+J89kJkoyc3dbSJC0SiMJ8EE1+GiI3Oj1xCjxgVI/lsxcc
5/2o13bgHR9YJ+Us51XhXi2lf4Q5vQJA5yOoV5nFKAoHNMuNSKnBlxLFIi/TeNMK
1uE+dJC0vuHz+3nGHh0nRblMijG4tSN1AE12AooDHS4emM3mNe3XiiGGkJdJcTl2
2emkCAIWF8qAZFCuB3bO0tYCISdohggCPdQ643D6+Ro/gDmdFoC/1VqZ63nmyyFC
yWOLr8n4PIoNkX1H+PlGMysbsioPnw2SpnAl42WS9/slONdZCKDj8mP7mh3QgJUN
E248SghsL4PId5JfmBtddUwRIHjUErUfvBqQmTjb5iSiRY8Uoj2SSvpWPANuEpFx
bAI9gwhWCEJHgaPbWALL6ScsL4mg9anh+Fm63E7q2g/3DP4SaAzpgNt612/k7DQH
o3sJ5RFYUWnk5lVhnmrZ5ZVoLZQOidqX/81Bmgf3bQNMJgN75AxNI9lOlV4SHfXr
TfLFGYnN6udBIrt26Pe6AE58FFnpdwurjF6THlnGZQPrQOZr4a3MZU84H7hs1COH
O/4LXi/wWiKPAnoUELOnXc5ipXe283MTHw+THmGcoHKco3n7EtJNKCXQrwhJAfRc
E7iYtLMjujsexzLJNTKg0I5c4T33YzzK5tukLkmFciZ06jfg/5Dbd3G3NlptniV/
CA1jihEZxEssrZSGGVUwIvCQ9smKsLWKTdDSBvDYvKumhjHVzrm7GK1hxGcwt2QO
klNtKHHVLZUYNkgFifOsJM5yRIz5lQBYvzaGKCt8dwHP7I+hy8tbGRznSHt1elt2
vje51D7jmWVzWvNVkOADm+ehglvFis1xLzgVVHvnQRA29FU3+mjFqwl3oVa87o+Q
4RlgPC2HCZu0Kn1ERIc54pHtL5vCniJ/VZsZPr8aP5YPLR3qsMfghdJYnoSN9MTI
KDaHRfQhHXkcU0zGCEklSaZz4ciFQLw9oCmzIjSVcsRxLQwjjRq5dkF9hFtWbaYh
yEfQt3Zm2E3cSfj+/Rm6KzsoJX/Nh889hQTXmFIz83bO518SGzWZLNEvrLmtObK7
PgruuGfTcNjX0uTMDF64YwjXMFER24ACcyVDN0ZYJwU4YGpIP19oVLbHXMjm1vza
h3g7tnBU0xfVYTPldVU+Y1QGHMeNaYQZqjhw0vZ++0NJxhtJEDenpPX8w6kvqh68
f+yMmqVb35jXGOAniXcwEicglOD7OHQjfAapr3VQrJQ2EB01EjsKbJhXzwatlgVS
Vsa1BWmsuSJnZW8v2kJF8GzhYFnx58VWkKtdK3KfYqQrx4l1f3dmpuIGcGi6L7Cy
N+WOB6z//lnxCulE+WK5Pnm6CG5O8IWqNB2D+y/zNTMtPJxL/xe26WhvJTsTnz56
ndhHHJlDkujuLHO3lBkAwUzCPaQwimS7gcDCBYHkg2/gemixbmY1EemRILuvcZZn
9rzLKOpFQ1EcSGVZ496OfWiTCxScBIak8suSq49zYa6oCEHN4pmO1W/i0AHZARVa
0NG4jIFjPdo3R/VAHZeOsjj0ADSXDEuc1DovJuaL//LCqGKHD/uU1tr2h5Dd7ORH
hNj1t/C5RM/Zbwaf0uPiFVY7pXHhjPu4BVaUaIftOKXhxKv85i5/j5rvnicGuWZr
w6Js1QZ1vJ85EcLtQF3JFKC76RkiEIIKYLJ/eGvS1T4XnQpAQlfdl9fcFgvLI83Q
nrG9Kk8XCGY9Y/+t1KS0QCCDmF9WMT5En0W5YMl4/kVmZDtOTRoFjkNoYQVJOl1Z
RqQivseio3l8Vq3RoYd5QTAP9h3X65kUAjciYkjc7A3KBs5O2jYhzuq8T37HtkBf
XMNJkF5mJOVbw+Yr2CCxhI7WSovbRgl8w4jLuvQ/jNroS1Vy/XL9gXvI8i7nxUd8
vXdeBpsiBadri5+m9rUlspB6xcJonlhHXfNZ7czZaQ14bsLHXHNWSpNsVy5MOTjN
gN+i6nkmQBfmFioOhYTlg/ImF6IqGpioCxKrDiquyC1RI7j7WQ/IutqpMHMXhNWm
9jeo187hfVzGGRjjSEdEEnAX8llmv8+9q6LKF9bPne4UIKnlJRTP+PANU7C5lt8t
z0zfyr8TRLdOijeniL8/1FNxSpGPYeuUimQBsu1qr2C2y1A/YHGSvWalV1YX5w46
XolkUVB9QMEclPP/pojAvKp3dEgMnIT5gElYAQh4n2W0s9gZgAV6kh/zBOn+QIwi
7MecV+Y0T80/2hASTffUAHMkOFF/yiyb+l+hseNe7gi+BlQ/PugsOC6nPiGcS6LL
F6GAK3E5XeBX3Bb/wC4eH+GEXfbYYqTVvI+yISGG5uQ9zqxguutZY3+DDmY0ICuc
+Nv9RFI0RoIO1NEUw7khu4olYQ/TL1lBpWChzZBUQ4C/Q90IYOG72sbdBKoFZtFh
IIFWlfU/a1uylnyUPV7+MaRcTStzWy2ihVyTiTQCowZ1CTWyJ24nKHHq3W1qkInB
cTeUH27AB8i2XnoO+r6o4KDVoYHSlyzsmahEstB6PUC+Ua5H/R4rhMAQRzt4Miti
8FlAmAoXpY/69f7j1dBNJDerrKz+4BZhBYj1rD9fGnGSTK3FO8tYTDnsSP9dpzna
BqFtKr4vAEBPsgeCibZyal0Ggl3kySlzb3mOaONaYuEBmTltePHO7/ByPooiSDY1
xHQ5y4ThxwKC/TSslQ5jssyWnt+S5wKQ2NKvtC+KUYtQ8QEBuoRuMV/K8m9hFmCG
MQ5swkp2WqDsYjKiuT3UOarCRSy84DJWx0gUzOvMHezgnjYAYO9G3t8nOWZQm9Ep
qIatWsIdDXI7miYDk3+89DfEy1EqcxkzvkBrnrwk+Co4ZnveJRYxXhL52oQP9fE2
J66yZq32/bt6fq/nkidkeGX2nRIZ/d800NCRETE3Es8GuJcAKVPZZ5RO9StzJpwL
VxigxhUFcUGxVYB+oDr5rlQ9CWsE/u3h6+oVUsYKrAW5H3f0b+v87Y8lZIez2nWq
0RHqZj95axYNMGNsa/aADcV7l55czkDff3Wkl66wPNjR+iCsp8DdkOQUFOdzMPbY
+7uehEb8gZ7ClkkRDbq3WT+SuCkVIwJkJnLCD6uptiGlRwzX3DtNbvb/2I0z/qmY
CeX91DJU9vUwSZGfK14CStMg999dHqQweIklDjGe77tLG0gnPaeD5azIojsHLHCb
ka4HBcoFYIwJSwfr8pwFUZeBEaDIsIDrHHrlv+1mI1yanAG4D1jBSg5Ck+PVaIeB
GwTK8eyD6HmrjTE+RgDs8he2mDX4lmuBIdNpIZdfYAGEpPD5jwjrJ5urzB3N9iLW
bxkarTU9Wb0bzf052EgKIrD60dA2ziVmOVecPtKt04CnH/0m8o2zdfbknBg0Uhbx
sPFmp79c28eTWTSyQyXg576H+ZIbVaB7lo4poVIRPL4dC+oFnppwbxardBSYdZD0
120jafrm8glHq5S6tEgiG2SFwn8mo2Ie4W8RVwRDk72MuGSbCTf1XZajLd1R2tW9
1uiijiEeSQmkGRt2GBIswt8mIC7IJQh+PwhQrid2i60OjLzvNxOxWXCsyt7pN4Zu
jmBGRnD2wjX73jdSKW2EV7MqOE2mQPwnk7JdBW1cWuPqTohbKmVSgJn5zmrCjJ0J
MXlIb6iU+9sJGT3sbWGJTrA4i/eoBveDrYLzXnX83tdULV+9eadqzI6ugTvS+eIM
IvXRN5HHNgiwcPHVHCApg82wn8zOohSUrzbMx/43K+DhdcP7EIBdCes17S5wBmYj
FzBMJlO3T2Rlbgc82yj0Lgu2yWm5iItnPLpigU7pp06IrcN5aXcgEuUTsvdB/EfG
dMwnFf01vtRzojI/RYqR6ZaGlp9ouJFUgxuVBrcpzLWbqmUhwb7Er3j4eJKQ42br
L5ANVPKQs2F10AWglb8bYPOxvG98vuA0bh1QSqliFnk7FhNbm3zVt+GAe0j+Ejjo
0SWtmAonLUpL4tDf3XLyHZOei86LrdtqJ0ba9sEE0d7FO7rIVGazHqZPmrsIR9/G
GoWFJH7yz+bCrM5SymiRO5fcBZdCUA1fvAxwfId0hmU17SyMFVTEHhY8B10IK4My
bHNrqiN6Pm15ZhbWEYqXvUD4UGAARWWB9bf0uGmt4siec9IOCXtxhAP+jcOD1CGg
d5Gfi6/p1DbPwrKHRljbpLPJm4Ya7nSPtOlrawWHhf+8A7bJmW4pJoXLSF4/jRtj
8GLFY0RoRJ+o4QgwgUDMp02km0v7xmx5eEuKGk77iw0IpuD7Gf8URY6oFiScaONZ
jx98iy18ZoxnMIJP6yk0Mvbeel5L25+uIYOtP7VonrjRbKUW/4p9TTvmYLhT/TNZ
Sq/ELkFtbIVaInESkrOSeP/SpLPn75AOvEvOSJmkHcvqNG566b6VJO+I0QnH3Jqe
4K5nlmSMi0tlkbjSrvPupPcGtqJez8OtETkGC5Ta2ghrXElqt0OHtNjaxzZKPbQ+
1spzqIbGv3RVOmORFB6mV2U4hysuoJMwS/rTV/OKBnKiI8cFK1JQR2f5ahrieATS
MF8isD+8uo5SavhdKK3k7INL5OA02+qN7EQCXioZgph8X4IKuJhv4HZfa4UU+xYO
MvyFPp6Gi/8YupVnhKuUkJXPzwUnSFYkMHlzgjZg7KyaVUnem9onOMRqMg0OYQBb
JCTInZ0IC28c1DIm8oldVsV+Bd1k2hjdPCPhB4isQfxRozC6HZQIq+hDLyz6rztK
uQHczatdznqnMI8XqP59Jipzv2bWOU1V7BF6V/cBtkXc2whK0MnXRAVu5aJuB5DC
Hcyw20LbW9Jknw2k1iOaNIAkzSb/ux9Du7WHlsO9XiA0fMQYtyOl4lyDBBwLxCvI
V0IXBnwSxjXwCw/1UUvOnsirsQRO/WZPwJKS0NMPQS18X7BtelascU1O7r17/uXh
NMggbEBVDHeKeeYQP8kLZryoPi2UT/xgi37c08zInQgh5ayvsJwZws55gFA548s2
d7z93JGR6Tl3kdfymwm0UFhDeVVRovcmq4U7bbuxruKVN8J29pnOhd+FnDpeK2/4
ceMX6Onex2Jw6RZ5NxxyS+H89PvoA/gULn5VM9yKyjNlGtzIZJvba0i1PIzDEGjB
XNBgLYWXoT9fzfsBb2k6ZaLOjj3HWMX/f2t/6+MsJrQpWZC2lb6IL6TFoXhI2j06
mV5nNQHMn/1J8k+kLHGzybCz1fHFkRpU9TCL6gw1jrTheMCqIVwCb0RMOpUjLXNH
3F07RdZp6aQ249J3mQZq2g8w0ppKXmdzFx8I+WfLeMAKFrN3jJNcTlb8IFvI8aqb
PuSdSi71ojqiarTTdvdesGZ9DooMt9pmIxkVZuo830INbSYOkZxVVqkpz7Nj8CDS
o3fYQTJ+v4P08gDIUxCoQYnF8xdnYMaSyWAusgebM42dM8Ojl46SClz6x2v1xmPz
cS7VqKPaCgaQ2+FK9/gN8tY5Z+BtABsh0dLd82vFLwX2yn9jm1WcHydTAYmq4Bps
YhsLQHJtq3hTTORhHRO2GLvAAb9fscrUQ33eE/p0XHV4XdAiPkXDUWOCdhZ4rMEV
ePZxyh+vMukcSekYxWlsIE7vMxzXmVxvqTl8a226F1OA2Bx1x7oPFEfN5Pgzjnyi
e62ZDGdWqi0hOtAFzB/rwh7lGQjR1wTYD+iA0dnVGWoecQj4GV7wmMZf47pglyz0
0l2BywLGWQxoV126NQUlsiDz+fEtjdDbNhZx6IUlEjmfJD5F7RnIolSsQivSY2AM
pO3jk9XqOHJZ8+77ohOh4Fq3AxJz7yYFSJs4DmhoOG1DTIEGFgQD5HUYw51Csrgo
vWQH2a7KCEGEhXS6DZTdn4559a+5UIoKpvZr/S5t9/p0xe47/2mlUGlAXr18SYwa
G/k13JkUeiURtqVPLP+8G+X/v7X287+zWUbeQ7+xdd06bDuHKg4tCTJyNRsaucCt
RaIjmtaBhsxSUaVBYN+5HzAPLG5LzMOB7o/kG0oDjqiSXHioRAMoIcqPvi/zkhlK
ILz2xo+Hy2aKAe8Cx4DlKA3gPZoQFi86mTSmGqXdbG+IWeGmLdCsNRcE24LWZBo/
Sv2PDUClFV0+wqxspvm7SdsNS48PiIZ3NVU+/gKWugf/2617KNMd6jeMrZYFTxmW
txFpkEP1CnXtzEG9bk6vuAdZIKXxX9x8mV/WS1v4wOogthP7n6YvOPF82hKMX9gb
w9i61iERsnDpet4vNwPtxJQ17xkuSldcp2jyG/SycluKmLvgOg3T6rJLQfTSbIOO
Q5Cz2it9UToRXFWIaJ0cp7qHszPhO5ltvNdsNUsv1upmfaP4YCoax1FRsnpJA6hv
dV0LLgUcehno/5vK5VQBo66ZyxXYRYX+QOQBbw9zhiZfSWNv3KlhqfZDR/LUYpEj
TR+0ZREIEZiQ/+tT6q7WZIyvBF7kyiZJW/IAOj8szvutrfmBU0u6JmsN0TbOf44+
jKuc1Hk2T8bVDUdO1TR0G5XqwFueFGm6O3EZJZDLiyI8tHXrMCwLCvIA8/tDRtJ7
BLFo79v431vHWqARb2rUIxAIqaFb4FC7R6qTUHRf6hiUWUpRx3usUQpK8m8yWqrm
SUcI7g5LoVC3Sdqf12TIfecBbh/diddk9IvKa1w41g4KL2ojVF15iNujHnM9WjDv
OepMUmc3TqVomH+D8ywCluzqNGMwXHasLmJeA5wuTw28Qor5KqmMwcA++RXFdWYB
CJWXm+spN9en0S6GgLEyUT14D+V6s3geOqvfHOKa07YI14dHmsFweA49Pgs52/O9
Ma6NiU+1PvdVmTdHvAIvcNlXv5XQPnhgLan+GPi/qkwt/UjqBqB99QIj2aMZnkAY
Uls3NZsV98T2YKJSdkcCCGyu7Vv/LJZ8x7ovVm2tD597JRFsyJxfVmBVgjUD5Gwv
ipAss76/UF1dBMnU50v4Uaqz1oTrKJTIk1iuRUrvu1dJfaDlsPkQA9UdVJZTPq13
NHILWE6+hRu9D+YykWhPfAfqQXGdYF1Jp3urH9GCNXF3tkYJoviwNmxPXa0i4dD1
6uxoQc1IBIP57Vj2mQ607dDNE6Zw0YTgKDDoAlRyTeMwW6//eqYp1TYC1KvZxSQ5
T64njzCwXp9BzvXTdtsk1yHQqQ6Yt2Et+5o3ExQ1zyxq6CAciM7BsuYPobo6aIhD
NthaQEbbH5ZvRMKXcJb8ksJzpnHYp5Vwgt+PDW/4RIkL9QnLFEmGCG8lq1Vnedk6
erIf2Kssl1t7ta0gLgymE40EKN5A/UDZIWt4U/wRs6W4sB85vKpCg6WoXaiPLjtq
qDYhhmL2JAN7LAYtoB19spgMdDybAxD970Jth5T0i5F9uQanguWot9iLNk8BBV5j
USLfuuNMQC1mmk3nikt5x+fNGrfZIBpwv2ME2mEIMYKAPZIUnwPS557LbSCeEuLO
2jcq5Wmlff6ltEu9cNQJo9GDVYEly5SJotD0Mp129Q4Fo3KReKrvmgNHQFSzcL3J
B9EMeMsfTmi0q3mMB2/8OWihiqQ3/SsZs2T6WXiBLOQXPqmNWYDytMxvbeXM6AAZ
jmi0bDofbXTMTAFwD9xIy1GkPKzmRIo+NeB40xkNIBTELaFiKsNunj0vP/peeyBC
rC1Y0G9rzvbmMFpIcvKR86yzOGMzKM+qBuvi2NWNW63h+Xlo5NtJQHD+V7keXk6g
x5rGZZYSY0LRjGkkoyb5QDzlmLMqhNjlgwIOpCf8ajyNHVS18EClWaV0SM4LYdh0
UMJmhrFFa3zu3So37CufrU5eArhfIZVbF5dpGinD3UNj/P0xTlkkmOPjk0iDSXaf
KYy1NL9Dw0Cfz6uKS0WOok5PcTID45r0bdrEfQB0r3YunOIz6J3kRipxUfhHpIbi
v/+ODhbc0e8b04ZTeL/7yAP62l/EuetfbIMFhvvBWgBZKBbiG7FsMa6dX/mRJKEI
x3B/ZR+KKgGrj/3R/6OZrQJ4637ffY6nnEA6fZZ+Ufxk8TrIthdCsDueS1RbdI38
QFMZqyj9MdLpfJ7BFqzRjmfD7MyAwSV0fC3603iyq4339TVwJhyFOJLK0sxXcMhI
w61r10q08pCP3uZF+7D2SB0nxHJimnzDF8RLDgMkGTwxyASVdczzFYnnv7mKZ8rw
ewPgdjdMhP033JlS45pjnoHl5uX7+ciHCc4SC1II0xgzMAqtWX1UcWhle24s9LvK
IuV7G8/ze5VttQZM63UygfGQLz7IeypuI/jFznPiVMKrPQAmkaZUyts4UwuFfrpk
/OS4emHWsX0UYy8SLNSAoyTvcFo4417zI2U+ijhXVEo+jfCQzotjOo+4hPOz2NjF
/Ih1gE0UP9xZ/8/FPAp4Bacs63993oJkBuVHTeNOsoCPc7Ucoj+j2yeybvweRiPm
DtpPco/sOAdn71muGxKJu4CU/e9hzA13jD823t1wMZ+rhkUdz1LvsKMN/zzD5jGf
W+t973ffwplwfnfArpYCWkpWZ2Vb4ht3N754e+TNycVD4HLtybwEPJiAAQvMdGa8
nvzdjsx5YcU7D12S9ram0yF2EmpbnYk9ZyncwGLfc/lyNpkOIi7uu0BcNc/B5ZkG
2VIDc4O/p0A/MjdOyT3NjM0cl5zTnTyXRXK1jcVM6b9YQw02y5MpbnmQKZ38JxC5
a+cKA8bW22EMdeyH+cVRv2o2byS6ZXioNuUWqfnUQy0Kl3O54jrL21pAcdp//4eZ
IQ2ilemP3LCLnV1ZgUwKQ8T1s2Qr+XtCgMT6VyS98uUdK8GeTYuAJ0fcaJE7Dlr1
whktadjh4z9GioCzk59b7mB6qRTazasjASk+BJMP+91z6ucUjYJM7lGD86o4HO0w
V7D+OOqUTYc7w1TPt34PAzChM/WRkJswtlPeSoOuqNBbHFFLKwp5kQE+t7XtDAZS
udLLyxt2jtdg1vdLKZZyKpBHgjaZRHlrb33Inx2O0EoMSuCQy5aZyLhK8Kb1vXFS
s9SLlxmBZ8mYhMdkXIJgvEdjtxgsqR6QgK4knlfaQyhC7cke8UaRwLwoHoELXPtH
sw3p8lCm3aNrf4wueNY9I4yjEpCx0IsQVJohYHSNMyz50b5A4AFQYBklOBLwXMab
jqfpRW9YTKvFNCso5I5kibG2XHRfVE4JG2casj+HAqNM9f6emRmcARFw7bpqLv63
BfS5m0k69dIEpz5gh8+vsOYHA7Vyp45BYDxJLWxakEvwdnOEDadobpZVs12yDLNu
1XZ5FCvuC8tQaWszH/ltwpoT2bojbOtIx4PV+egWLV9Z0eTCs4i/ZVWHh1xQphV8
FrIAqL+gT9ePuzKFWLQ32eH8aQFc3k+OF4KR9i+5GI7+OEM/s93ibtl4HC+CoCmG
1iIukCy2mDNkmwdDJ/q62MMqqkWKo7lMsWy1naYA0w93i43byEu0WfHAl1+4Sjwf
mfUqD+yZ9iM3UCEPYI3TWO9mICbEmNEXIIfjkxbXz31KrbwjK1ACbQ4y0Ns9UG0g
H9jRQluKbbTB+MNqPc/2TQ5tjkvjzrjWqQebqm9mcQuHaCIiPdD1x7Rkb88zb9ut
vSgbjQL5XFOg370v7OOm+k+0/Ts237UpiCJUC2VnQDsRnx7c4nYGGV/sR5WDHbjp
WxaqCTM6kRDLFvYZRZXvvhF1etQc3a9FHzENq6a3kuF1U0nev7zcmCRgdrbY/c6v
SjtO+YGeraHOs2mVnBi3Mw8Zpp2NR0EdmMIwGbFbfMN+I4INLF6SYI+vqXBYpveU
Bw0D9m/k22GAlh7hbN0xuawMvDJOaE2CYG2HA7uYaot0XUsjNOXPoGdJUn+1o8VK
oLDEXVldpUm7ApcuWb5htyZ2XP9c8u/bONxEQtN23hvNagWh0viE4Pz3ffkCa2fK
h1Eel16F6Nhd3o0tVLv//16eD1AVPRKUS6r07JeMRIh2k5V1lQZ539SxSl7uAWKj
np2ENVuTDHHc1LWCWfF9sufjpVh83CQ2PZ32Y9O1PBiCGBMOSUVcmZNc1aVylt69
u8JSl+jUNjVAw+0VbpvbiMNzy0l2NBg44Pz7Q+bFiTX/ww4bhQws0AjXMfWTbSs1
6ZNbvWSqb0O8N21Bt9vOLVqN1QEfwQgxT65i8i0dZ9S2bLhoLxub+YTvZswVxVdG
gBEGby7Z4E3BFt1XY6MGsYe6/A6+PbUbYhEohrzqe9GbQQroK074JZi0hTXP91bT
n7Jphs6cGMvVAKBVc2+D4C4ZmQXpWd6mqTOI+EpFQnqs+052ErJ4hTEUi+k3EG4l
bIsG8rySPiU0GoCRjsf3ecU2EdUfvwrKJj6nYLuP/XCOLogfdzXkeT2FG1G8TNSx
JLGJBWGX4PXc3Tq0Fpwe9Vau9bURubF+SF4bw0Z4R9FJasE0dxRep58e+kWoOfIp
HhVPd5+5sdbvGRu6GHp3IllrpWaO4jjO9LLvcNhHos3nCOcXBo/lUb9jHXzgGahY
ibmBz423W9dM4piWQvG9FnCWxErc/+BmgcCh4jPhRng5ObnaKng44u7s3HZG1AuP
aPvxiYmulh0ok4eoDBaxBxaDJa2VPTvN+uDk9hgawj4zEl7Cqne42OnQsBXkrvbm
xT2DZaI2JNvrK01bwDg/0pDz5/wAlfNbh8wNhN7kGGuQ8YxeY9Od5rXQpCRm/ZtE
bSEK0x12f4f9C03hxsLC5UBX9k9zZnVcKAWz8v6rm0Iw0jEAYpJ78TeY0tYytmGX
hHiqy8C3h7F2gSbE03bid5jGR7usGkJ/dk0es3g+01EWhDEEWwr6XIt/EUSRee5C
UXP8Ny+fu3b1/aHlLFXLePw1bjKCLEVEDItSrVLAZEgrf/bMw2JZ3LEfe56LUPhZ
qb+//VrxI7YFY2jE9x0uhI8he89MGVUL5bZYMyeyYpmH+V+AJIWNDacXkTbT9xFx
fIddI4mv9d0kf1EiWSno+b6kaVy+zwOlqvfldEiATRNdEGw7wJMKrT0OkWicCRQT
WVJKsVXqSZ/TJhpfeRUDB/O86d9+jfHtbIsA/6gI4ZQpEQf7hOnSSdHrsS9tZ5NX
tVDVH5CiuLHVInZ7tY87TSRtHnwahEO02Db7Grem/lnrwUQkiFEAyOgNTFmDeLXe
5u1VvOrZ2VEPSxlqDAl4wT+/O1OxfaVFk4wCtgXZTns7UjYOkhHIsp+WOiYs/Mrt
WhVV2oC0ppGd8DSRoBtdSksy2wfsZgJfqEtIIzSOfBtVR0m8/oOfWmYgXHXc2of/
UAM1ORh7t77q2r9yTlsH3dJAkbekpY5JrvAsQvTopsAHoVSmyPEMGsY2pH5+DDij
LPSBE9agQSQP0WExVQrpomqkTVfnJGbFmzJ+tXrtKjTTFQHHMybCwYhXD5jP2NuI
UCSpeXtyfEXmP2DI0Eo2CN1owhvKgUh+CGNP4/ajrBx8prPN7cYh2bpQSvSgU0vR
FJRTkmHu1sD9lLcEo7Kfwb1ZXSvR/dM5kPMcY7o/kvQB023FYqa8x3l9x9rOmu1I
4n3KKWpX0a5gLcrSglEysI7wA93oiOOiZMOBpPDC5Q5nudyEHp/lDqWk6fzLihKv
WE6PASmmmlSHSFmsx/TZaIZepkqAiFRlpH1Mv47Ti6GHq7imWIlHdMWLuM0WoDz+
ZtB+oMFGFDwCaMCbEDrzHs9M8n0CksPvLUiM+qs6pl7x21SgOelIYneuLNEUwYQn
0rYoaQ4KSd+LnEI/DTRNN7pmyYre7rCSzamt2yPX8zXxPj4lxpF17WC/ZEpGgeL4
0wuFzvDqq1TNMpbdYTGNXrNgAZr+oLXyXZebllqUh4BG2b9pgZpT3iSxnJQx6Pba
grzxHg8SltViBe/jgNFFwSf4tTfCjbd5jrROwHtp98x269CBiqQUS8wiE5wdBt8z
c9YfqHDlSCLrx+sreS4AOYdD6IedNXyradjkH3ahQfPqUlkDHQFrlaGjM1U9DtKX
20AcphTN1ao37k4IIHArkWqCAXgWqBitUDyE5grTcigyfArSw4pAUtEfbAZrajxp
LXbK6V+prIz9oqVL01WIpGNiVVNJrs6dx/ECoCsZFDHmu0CPup97jZnSa1PkIxC2
maEd8+D+26etVscK+NfpAedqR3IlpDgvSiArB0fOC35tfPR0Qckd5s024eSIQsFD
RidEoP+/iuDVGtOaa4gzLRUx2y/6G/a71bvxUZE9I2hCPTCZWzQuUy+YCPl7UNFX
5HAtvO7kuRa70PUTKWrd5Ug1KiS6ahNmtNmma71Cop8VI1ITzmBf2xxzJOGmdnPM
EOx+Kz0Sk3080fxfBMU0m2c9nq2cmmUYDMmbBSXEluCd9IJV1DElebvopWIR/DRq
M1yQYSBxsqPJxrYH7wQ5NcN18ciQVvFJBETufil4vWwtcQFt+Sx7HqZotiQ2Fyzd
2/SgsnkU5WgdMBy9S4iVhaDYXat4J3+o2G+Zq7NpQlzJgGeLEqvwPSbDDvAlMAhN
Pfhv3tYY/AX3utCgqiPw7qyJ55q/S7qW/SS64/ukoGj2uKufG8L9ttTeZlcjWooK
Jz2WJ/tu5VyO3xa+JI0VjOEWCiz6kUGrm18h7tUTHoNGFVmXWcpJOuUzEJSmtjLD
AFZ/zP4IsipjthCbTFyxFb4dfZgucA866lOiQFLCaYE0+CwOAPVLmEISnig+ZISb
33VukdtjiGyEMtSqFgN99yygfucOKEZkt9oRt+pl4laDf3MHjOF0AWQErF+cYx0V
i5mpvztGJr8+XsvmfgXzYJNZ7adMNCOy2lUnYxXhfEVxtYj9BcRJRaB5lzURL1xb
iGDt5WFGIpblrLWpnpX26+qKhDdJLazEFXph0hHo2AH1mbWRVCbnbzDBhyMENskO
LOlOvWY3hcgDuFbIE17lyUYD0mZlWe+dt+iRit3Zhp/CCnAnVFkWYuaqUUWzf5ff
79XFVVUPeRH6tHAvy4I4T1m1lY34+vsUQs8Zdja/wfxHL/LWyatZ9/tSiX+3qMJp
3oud1emEIzdMSa8gbSqmBqEvj4RZqJNIT88y1O/OwfIVpQci4M6szTaQAgvSh1yX
LvCrKZBrCm8RSOyGS8PrxgLK77M/NwA2OTkJhhmG9uScFJsnvU/Djlw7TPtUU/vT
CS2O5L/oSg2DP5NbduFZCxawzovQJbFqh0thAZiHwCl9Op55wYaZsywx8nUzsn5c
NcGQzRxu56r0ZvuOLLGoYPzdeOsWnyy8iT+3MRA68Dlje5wDG9W5gmDn3JyYpONO
9ddR0W6UG1mcUHDQiQdOTbaY1zcMZJBsCZvGMk5agEjkzNE6UcjxnV/qlUOdhYmJ
e7xgNiOiogdogAjrzPkEuPI3E8vgNWsRPRRWX0wOhr7BG/EvZP3Le5VPvZUY2KVg
xwi2fhhw0XDp7N4W1injD67OmX3jR0zLgVdwFhVQvK8gWGw/LYjvr+Q3RN0lzX7O
o1mnV7/5Ualug2UqupHgMq52qDD/6xzsWnT77e0gtaoTyRFtJjGq3ilSMBQIJMZq
Q1i01Mq2ON4UOI7+1lrd4UcSciUDwrfVSg+ag5hDuXUGnrdOnnzV1qnR7l2KBP0V
kxI0e/t69BLXMEwAJPItRrAuAKLxAbF273Jr86Hb0SIJ151u7t6rqkyULINjYMxc
2lXJOnDdeEzXFTPdO7xB7TCDx2QoWYrCC+tzEQcluaQT80mDVhvddWS1CZGqtYgM
sQDEWvay7DhZ2TMS7QPmqVephfIdGqn8VWF+HiFfeITCZ/5lt5Y2Xv6YJfDJIqTS
3BNT/TYoH+JiMgEElbsQ7hjHd+QQMmRDXx3HcR9+kVvfYWaMMlKpb39udnKFu2YB
KXRCvBx7eV9xqniRT/ye+glzQBEBCjJ6VKOyvo7+l8SAR53aabNAVO5befQ+Xw7j
HRKq0zP+SvM+5W332YrqcI2sQkZjGR12sdAcEUONtwvARAh0Kx+cIXY+pIdGvUEj
CQzIoP7dk72wS1d/GL3jDz8CjJtxXtzZt5aQYVzb7Tc4nf3Zu9BBhakLaLCUH8Td
a7DgteMty5R/T4N9qGUi7Y+grN3roWUSZYwZMcNXQIgUuKPQy1ss/TUM19ZNpp6Y
25icxkxOpHExrr1e+AhycFlWsz+XtG38ci7foWnhYo5kitKbl50rTG+0cdEt3ImH
Rp59vjnFNXJKKkfaBjHwn4g3dk0ce+nhXIMBVRJBJNkSi4W+YLBv2THjAe5wdBvy
9H+Q5Di20qoYMc9W8cwfoDyooohJl9UvpBeguCD4HB4mOIWVPIjdEIDvuJ9nJ9TO
Co/WybEA52N2o08gT2Gu5WXWyDco5aIeOhWH0V6YET8sdH7/NtoyIJOl444oNmpR
3Cyr0tLomsRMzmgSeCRShJd2WSP07ms0FuEX895F5ADs5VnwdYPJUA4Ra1DlFW+b
EPlAvR1t6VegYkImT1ufOX9UH9ISkJpQPyKanBpz5ceippLVdZwWLmw8sDsM+Pil
wNz1AaipFmwkyyaSjjr4cSMBr4fgqZVITcncwp70IQXODg0IcwfNdtnWcXVFd6ws
hH+h/gZ4Z+inwhjPj5/Z7jLfN9OCRO7zFQCzAkrr1vdSZWgWH9jU2n0jXtLQTT6n
OsmXnQJqCWHM7heeWHYWf4junBnTGHRb3pZSgwJsrkGCxsvyCpCrhWz9mK1j3Mf9
yaHmyVGXo9EU2xpfVzjIe21J3OL6xCcO+xshmgKfZGf5hXvTVusL1CcI0ufRLIAe
ygCdRkbvtA+/d6p2XLqmotatIaL6UeS24Ikmg14DvuyQI4mYEMMCDmSwd9pcfUeY
86F2fuZeBdkLQzD/agdx0JoEz1wSZ9oRcA89vow0Mi1uadR+E4fiJMgDtpJlNF/q
pY4ufmAGWSP0M2q4CfbBL47Jj+Z8Zwl7VlzH7KK0RWSPZpGxC30XyYMOjrRc/ddI
LTiHH5Lpuey7Ve/PZHi3YYDZ5G7UTlo7iBn2X5ZO6SNG8DDqN9LImauswhLBic2b
r0C3dlhE3GIsV4CW0DSHjwIyjYVrvJcJLyZjtMhGlVmL80YjmmpDz50qrAp6ht2t
FjF9paGFccCmSVi8zP8EiEgu77wrJU7pMpX74jh6maS6CftjRS2K0XcEiWZpRt8e
AioEwmU5Thka6kw5u2nQ5JWJ1uWSVAMlOaPZ862bkFaHsduJU3wCm9xfamsUEdoC
rXQ5T2hvfXMk3aewBQ7DKpORALjStoaZFWXpp1VdFgCS99feBq18oL12GkmI5GBp
3wAqlOl86At/rOZZC++4D4ieInk2e4o9JcgYJj4Quvi8lV0MO8BOdvCa5HHXuQpz
3M4kVf0nPrllUdRESh+aIZ1XDpHOG6sp0RkA2C8EJEaLqnjR5iKw94wAjUDvrEt8
+uSiHB+icJJDg5vhaqNzpCpiNVVB0M4zUqbak7Jsi9e/iGYR5Bdq423pfOF112uv
qAYLK1PlRyuCLfwRJ+eSpmnS4lt/A+oSQWaZChKte+Wg4stI1vVTcA/DSmXWzVFz
oa3d9SUgcei1icULW/w7AFjH86vnopiGmTISACmRSqFA7ztXZ9Ft35IReDINTL+i
i/F406DgFrpHA7cs4V0uAFC+FbpMMBGpbGYAFY6pja+iJ9dwhlMfCsiFQsRMt4b/
QLw47luMk7/OpwODekQ8QsTwY/JgEd6DAD+E37FIZB83uJ0c1iGEAMtDCmJB/906
LuCM9J2ElBi2Tdx2MHlsHq3GFZP1cnwDbBjy2z86r8RIEnNxHbRuwHhnFrzJJ3ab
WW3DkyvsuCNU7EYsvtqM10Cg7p0NujAov15WfkVlDTXavHqVcZF8AVFoNxcPgMzc
EoSDXFeTD3RiktfPmPx7BpTR/L6rtKybFi48LwMQmksqlSpIyz0eh//qjo2XWkCv
DVrBHzW+beaZM3etYbOCQiFW9Zb3P4mS56D95saXdOHOE2cutuQcbr6I+grhOuwf
ypVH3QRKJdbM9ml6lz1u6sj0pcl8Kq7mZJRwAry3aimB0utzs2lK+kWc7Ucn8yfE
NKkCFIFIe708zH/+5e1dDdVwYxMmXWfyKzR8WYYP6eRGP9Y5i3SfTbd3iGRKSiY5
D7kQdEMBPKF2zrw+62DGPCX6ihzqqGYo3+qBfauOaBsLMk767M/MnMp94ZnhIJVX
XMGN9y5MdbqtBDgPRL2s29qkafTpj4pDhp2yLa/vWzcYcqnxTF/ba4NsYMG3F9dl
OAF4KyQZSgodFF5FyV/ShLuvtk7HBmGLtdvz87Fjptxm4KIMi08q95VQBhqN5GaE
22KjZ8MzsmXB/5KoR9xZfUzfLJdmBgXMM7wlNBImcQn6PWV1zye1wm2F6z+QTBio
87+xZyG64lvj7cBuzjL0FZzubbEcmH95iFkPv1JM/fyJS95HnKezI6BRWKV4Fh6p
rUFTkVA5m4xm79GgA5O35pQGGYHnNJLV0r5lNhNLZz1ZfvMS0W8W71E5Vbo81adj
43A/0sjPRx1K9tt532Kms7WuH08byvrU3Gui44hRy9Dd5IBlE54GHmISJrHiN3Y8
LigEM8WZjJCMY3fsx8aQhlo3khqqvPmEPKlGz7vRGnf98dKuuJbRILD1ohx5XvHD
oCwT38hh0rPjdnPHaoFy+R0jv1lhBWfkN1atVg+on87VPu3c3cKwYhET664crfL3
kNMXLaDumiLDJEmQ0LoVJq7fL3pxMzWU3Np5U8rhX0hDJSVu3DX0E3Fw1CEJm0ik
RVfVz9UP5m2xtVT0Pu+OpinFtpMTRiQU21lHwPzH0M2Qd5XSDSnd1k1zhHWe/PRT
AxuPhB30NolRyyry7qhxN/PmJsmHvzNae6QvWPpGIlzTzZ1mOsKYp1Gm2OEm0Dt3
12rFeWJNQkfigbnXral8igFcfs5kB8Mf84JxnTCxBtY3cKEZ6kKFE6zWZMAsw626
nhzqqp3G1lCyjnn4Uqbnb/GCBJD6Cl/t8C/n3+BdVnIZEn4toDlMTGABRO/YVeHF
jeb+6HC1MkCChrTXzamnkgkJOIzQqCTAgeplTnifvCx0oE+1kASSgdxLPNyj3BOn
a9zgH5g3iyzwSc095AoL5bEpP2tGyCeVPych0udmXerO6oEid1wrbfjSgtSCsZ2y
1wUuvn168dB45IDWOa5wXTJyvpq8jdsL+uB9jdCPz4JtWY5kPwx2aoZImV2C7FM4
bSysrFqVTSahIAeaFfTmpMLX8yednvbRnl/6DRsqWr5liMfqVQMTB3xw51B1sskr
86gIbs+Wh1cW7D/I6dagXuI5KOXMUDrjsvLTvgudn3Op0lxtKPoisYynTvCWkxCl
Nz5m5yvaRObfNtfzNPUUm59N6G77Ezo7lDdcXenlAg2a0Z6HvGsd0IPmZd7uzhTb
i72X76uRICrfdnjbGqULXtzPM7nGhLWIxBeaml52kjb4FYMgWwicakjpZ7d2hg6F
YuwUvEtlxxO2LDB5b7Qc73hRa2EcfYSvoRFvhlNT1MCX39ldcoHItNY4eC3rTUpI
v4Uc7xwQo4TiFfrvTJXTExXaB9BNuUdKkpLrWqWWLP/W5BRFrG/L8MytVR+oJAc0
FIwo8+usgw2dFzPAxq3+C1lbWUaSRpkaAGpjFRe9YkEc1jDUP6lPDZ8Cd+6fZhMJ
yyHq+rsLaOYZduAkQyRrhz6JqdFqOhRP/DcRrhkitCKM4+3MO4we5tVim0UbGsx7
tbx/EzsAaxoJ1Wg6iFKO4iIYE65lD1IjqsKxJHQdK3aVv1iQ/l3Pegn5xNvpQs8a
YWlmFN1a8H9jPtWNmFpfIRA1JuYHgMzFIxc8mIq5oqqYurBgxyvgi/YubGt1j95f
o+QdSj39ub9UDkJtckLjh8XOiJ9rveaHxb5j5TeaV1ne5iKL62dRxPjGBAkSoUQC
naPKiiR441quXv4v5KDI9CJCG2bLh4bIiXOkKcBSXPChIN7juJJGrk+45Uio2qXM
RUE1xun+1P54CobNJO1ImXzsPRFkHeCfNxfb5e78Ytz+Tgy3mBFSnC8Fd2CvzART
cf/PRIJ3C+rPG/MFkd0+XAvwNktK9Plj6pHnIsDt3Rr7yuhXoBCZeuJ8YMZ6izNr
B/7BZmTppdb+dU9/pQQYhLlwmBO75ghoBu25ZDUVjhidCyymc/XWj6T1RtGLW2pi
ESRk8JcAfqvVmJ6widlYbYPfbCUEe15h0gS/InBPUFff+orzX1e+w3kbdh7XEwin
NTjktjjTHGtCen9WeujUdTsfItSN7To7j8uNJ5SBHeqDtkPV+JSbLWe2TbKvPvlR
fkYwT3SxA2GFlFUwvcQHAvwuaRnbhCwycbUH5Suu6YoINJHhspn0WvbSXEUf4sFp
hrcip3E5rj0zWkRr/Bhs/SLvqkUm4TY3AtWvSQLDh8bjqNt3d6uZtBJl0HfWxtxT
hwxmZJk0G0PIxlj1+LNvRQKBhnDDiAKxV7F28srH4h74WiYhOz2mSfdS//TGcEtP
cPhTx+8i80fQeE9y93qpXvgpJYXdhzXX4owEPgC+7FxSdjFPn7KLH88y51q1Kk0q
T33pNjDjSiMWD+2aw230ZQHK4wW6UBIjZvjH1KccQKAOV2Nu7XiHPtp126V7r4TD
EGMKgRqZdz5gQcJncBvI3NsWAkxNY12W53O+3gZpT3bwsvca9v6t5c8nXNY51qzr
z2DpuARSIAzyWtHRNLjznVf42raRm7d6fzW1sQ8EBg17/5erlI+kE/tXd0LwSxpL
BqsPi3FBNdNFLpmpCtq10zDj7ilE7sYJ5uvTBaJ0NBFQoYNW0IVhWzoBlx0S6nWy
zBfHiGxKV9QbuCkc1us5nWfSpmhfzVb3A7ccoP0qVYsWkERWAAIpqB28UeJgUBKP
TSB3JvLyi24RSZPNetuZvBuOgJp/tUpVrAluHHKt5Lgcx/jd7yGQGJdEzO7ToxmK
tZw6gZ/e5/7G8RtMLCG7kQMVuKyVTcpjmqFzMN/5ogvd2VDtRlnj+kaHGCeCXa3E
0KYdab20QJh6/VneKwthIOhxczU+zjABhm+kMXP+X263RrENcG9ME1w9C0gKn/c1
FHf7iXOAqCio/rPN60JJTqwM7wunmtYAIb/hxji5DSzx6Sm/dN/iAlYgdkgHR+d8
8PzuecZ9EbzgqdIGOfz6F8n4+wpDXyhMSJ/DUyYgxI77hZZJtjUBGMu67Ts3TOEp
bUkvQVGPjYCN9IRpW7KCRnHeH8pz9aZIEWWSpQ8POYvRZyfclZLc8fZMQW4ujGK0
pgSQdgbEMpPwVt9GdSKswq+cDWbrw0FzZvYAAGVbw1Ylf9eUu7rxHT6Y9FG7xzLq
4rVk8kmgJ1+XqRk84V2R0puiPGnLtIOg8hcK0378rKNvfHZvdaEAv0Uh4f4sodOL
EGn/mIjlpecaaMA/ZEJubohHDKd/oqHjYMfKyk8BwD/IHyplD1aQzAVxUg8DKEO0
iWw0UYfajlU0Dp/OYvReyTkWFjePja4tFKDXhkBbHsF97LygKpM4Ii19YalZPwOk
ilIeYu3nRsQ2/PBD62clpP7lmYHzdDthfjCq0vaa4Ukn3nWg/sJap3zzRxk+2HkL
l/p4ew2ipQKmSozhA9Ut/q/Z71ymPHVah8TVgLRoI13MXaJufuoEJ0SwoHkz/sbb
gXEunPJc1YG8hvD4tc3MzuLB6URaZWf2oIfXkMjy2aaE7rkMekqoWR9BqZtLdq4/
QTWvpoLd/y7e1FYq6bVDGV7tXErTy/2F50qOeuba9GgEeI+Z2+Qo91iFV7nyEm4J
lbsxgn7eVN1V6t2Gv3Ew1k7NfUTgrQfyPOkxOALXp3Im/OhZapgJd5hTErHY+FKV
ZOreTFvDvxqJZzGc7ji38a0SzTNB5TldFCiD9afhGJCuhhtWMoawSAHaBhVEfy0S
WX8XbnWYGHSmIh1tcx8sgKEFgH94Gvcikwj2eGyxGg/YIbtvdX5Kl/WPaF4Ozmbt
Zw3bIqs4UTlQT/gvSfOvkLx1pn36MN2jq1hepoCOfoxTlTXFlxhxILRZ969Aapvi
NhYsQ8rb8eKwUu7UB6rj+EYdcB7AR+A+ktePMmv9yIbFRnoCvTzR0yAfdgSg2hJ9
ZtJ1EZxWeQJl+gtBMokaTkfsPAXf3v5QjlR5/V2rMkxePbf329db72WkLqxnLVJD
DRgZCiwiPYuEEuhdEKp0ZzcNzkMVR7kjEIvj0KqAqbdNdy/pzi3ko8FzwrqeHErk
cU1hJOx15yAtHX6SJmhuSlvFVJqKZW7pOSlRNLSxJ/oSHyH29DGpjEuo1wtpoR2r
eCtlJMnBRU5R1gmPJuq9uIauYG+sP/aYi5FfPoAD/Pd8bfpszFsFQrg/PgLaU1cs
YvTCNYI41SmG5be8BfvDh3Bl/NaamYToMSI+7iuPASd/BD7BLwaSvocjerC+/nbU
0sbcJ1vYAXxvBSf6UV7QpkP0DDCeqGlWN4IsGkRoEzMUb80y0T/L2VdX2DQJ/Ciw
ClBeJX+/eIvDkyXDnnQ1l917MrhYqczM+3GQM2fBX157FQ5vDB/PTAdYPMkU9jhc
pVM3qKApJHeOkWt5C1ZRxPFGADToBwWHQcmsuBzwqTpyKyZ/3UTeYyBM1gngidJP
/LDaKIcga8dDJATDeovudmtWK1Tuz56Yh4oeqag2GBER/xCYcXjWFbcNVJ9DuYp8
CJE7TooRxwLGsGdiV584/uV+wfh2Hejte+LUa1EigYh1CiPALzMwtLCj8MI+/9Tg
IGbNKLdQ8kXTm8qYKPuEikYwe+NC1KL8Hx6RWGM3G1pfZfevJ01hkKXTEs7vdti/
Sixel88qZysDaKuKV7zz27Co8rWoAJZMiFBmmKWdz5uG4s1Kb6vPr6lYR84YAKII
+ZgrRU1NPquFW4IoDN/ZJtrK/aAiW+WRA/2rq9XMVrrd91czQ58m5RkkH7fw2oef
TsA4mvczzQZX2U8pnzh0Yye1WTnx5GAj19L+eTlKfqkvQBpEWs0GLTKCWU0p0yg1
x4t3BbbRrrpMR8o3vcN+FzV4AeH3exfHwYe0+0iToKzhGhTQGa1xK6RSz8iYL17A
x6hDcVG0+pMBvd2KGGdwDWpehNf/jq23Ps2j6vWFKnonZeyvpuF/p0sdCL0T8vBy
a5uKdnnqOENKJdlnjYE3nRydxngsu70ZOvmj4zUHHyxfxeGfc43ghoev+eNByuzu
c92ZJUuT9Eq+KLcOjcfbb+1vRajQmnCUP+wilHcePqNLaCCJCwunn0qCJE26NlCh
Kw2t3tuLnIz5SvgnpOgUWQcCP/6pJLIbLlyiwoUk6gbgfgsiA+ZkztLq0YPttEBa
OU/uql4TV3BWyYuhoh64/8rKoFXoug3pk6RBPFLAF4NxbMNX0VtzmH6C6GdvTzWT
5RTySDd2z0dRZneZ7ndQPb1GPeFAtdOJRNYu6PnO7RwVtBV+9GdYgSIcErlfkCgw
sd6PwxXDn/RD6Gq+uqgT8HqK/PEgsZfAQj9GRv4ZuCyt4UxSxMIhYklmZ+ryFGkx
aEA2v2wZrOBkXgXDzOG0j3K8oWKD2wP9c3UOwKmCsxpwdFs1c+rZajOTg3qhlwUo
w9HisBgWUlDIjIeSTP7U+yKXNr81/o/VjQODyggBktEAygJASGuLVKzCSlVviad1
p7+NsnG+I1j+aZAXvUItxHuKGhQeW+1/jaPAyzO0OvUaKD/K3TbQRnW78CHskFIb
qOsKrPxIstrsMPPmfKodaHzYpEb7ZL4Fmvmq34rL9+mGXT4PW2hwoYaINC/+SOM1
uyJx5OJyNfTwdmnA3dTAbmvRH6ypnebaPohLQvl8CxW8IyghimzAxhlLnXUal2ZK
XkyARDpiKro6EqRYmPcibHW5Jx98/Wl8BdzA/KRQbJXO/NInWNUQ+NvhxReFM6Q3
ZiFlNX4VPjx1vFo76B/EJBm+j6MirFzBjZMR2DtXP4xTgBYviMC3znDqR1SyqkR8
49eQWtUE5T4wo4xqLGtpHetND5ZTblWsiSkoxWvnSHakbOqeJ7vp3VA7uoc7XCd3
rqoF0i4Tg1V6ava0u8jhshm+4fr3MWRoQP75an+IN7pCT6E8BFumQF8BCnnAXk70
iKuf4zuOsNb3EM6aQGGv+ATImTmOoBXWoDFhkZA+jKMRGgtAEfzdUoEQMNpdrFvL
ikiA65PITCd5lKcj2mNN7//tX231J4Ntsl6zs5lwNg0gG02eVRyd/LgG3ggfysbi
h/YVeUYcqwm5mLRvN5t+eoG7EFg6E2Nhai+RcDxd77DOWkRVCSrw0rv/Kf+2yTvf
Org4GJoPDcB3pRO7kyAiToiK82OvVOppT6Xc5mmCGwfaTAiFCieFcCXXtczY7k+0
kEDwFQcO6OM8wZ7qUCMF+ygSSczSglXTYVl8re4makpO3TQUXIM3WrfQmTsJN+c8
MY1msoKWTXRjZICauzg60sy+qCgDSW0XiMNMz6Kyct97Kr3exRVCcVQ7avJKX8uU
cUMId2jGpDoOxIGD4VP/h0fun8pOg8hG39y0aCi/nbos6OG/Ra6Xg2fsaIeSz8RK
CcVOWNZPvGqx6bhyfDAY0n8kKS2IWRIG34ZWB0hO5UPPgxeSJWF3AaxvgHZ6oHI9
b6XeVfnw+oJpK79GBNlyQuDWZPV6kNAq4hTXf6VNZcfKsT5JkSDzqsKA8ljz8gDB
31MaLvOaBItowPfzTShAgWRB77FNL336yZLgIwnZEhh4mZY0HgPMMPmXQa5apkLF
U4GmaSOeh2KqlVp8nCGyj6zVY3psLL6bCqO5Yngr5AgzcMvExnLdY9wjVgYVdKlf
jIa4T/2v4qUWwgo61QyiT6z/KIhhwH95ouL6V+J7cE23xR8Cj/1JPczCsjjOinIW
Jf4adx+gvdrPQh32F38hOF6l/4DQ5haNazKMKfXW0AgXPJvOFiaLkMAWrothZJ/N
q/i9y53OH1atH5wIKVXmdw88CAQRQ5X10HrMbPlUB/yU+aUfSIPv1sGAid5eLg2i
MFdLqVC5/piAXx5nc0NeeMViyq1nlOa2uU5ng6B9Tvs9wmUxFCpZAgH8/1xgBj4W
s7OXYG5/cmA9zpNBqFD+VOn7b18lg3gOlr66RfjFc5p0Z0dHEHHBIX2Tapj7ug7R
cv9CM+QXovoN5YYWukRzwAuHv+xJWDNCnen5jV4EadL5Nr99e4lMrH6oL9l9GHfz
U5M1gnPdpvfFxnOuiyidiKL1xBW4AIQDq/ZWOY4VpwpMG+cqGob/mKQzrItzySex
/yUKQuvzKtQ7WCfouObTE0dIJexrj1WRwc4I+tsZXdWRVyMur5T5TkyO2VDbfDGh
0A876veb0Nbe66OC6Fidr8QlIm11dajirb0Lnyl6CYy42Avmr9fm+T2HthGVksFH
gXcux9KNlMPIV+jPgQbnKYeJXZNQQOtC5t80ultzlRjhuBXA1rXfKJp7TOY5uByb
eodVOc0ccCoLalYwoqSbrj8gcONSN2ihBq5aTFzRBFLmmno4ng11f9eZ5LquXZVG
GMw0fG8EVc4NQA+JEQSYynvkWTFXBGuyU3T7WJx8j6/G9fP3sEhtp7xelyRbpBhP
STQtGRP09lS6lNDiV//nXKlGQg0ddglm85figyxNxyfKe+BbUyH2BpPt706h4eu1
vNVXcrIBaDUTOlb0DAx2U8LYG9qpMSEBFX5cPtB1sgfLJ/syOxxDYDT9tviZJvpm
s0yYhKHqcu5mFA3uiy25bywF2F+eQQYNhUVWQwdHAaVAxIuANrmR22Gulc1yQUhm
g864WMOfnXdjqIApjiXxgZIvdvH2lRk4ilo2uluqOyqZDnzYBE732M9oGdL24+Nf
AGx0XXcU3lWTeZPgGaJ0qJUvSalryozGXFc31wfAobiDE+6SOMJxmyVwgtQgydnm
3LlT22r41FBmxtaPssJ0L6QTgnSBA+2ZzcQt0Ws3m2X96ovIQC+0P60xjnKDcrtF
pkRpSnQ09wOASke5GrChDjupkWlgt+Xh9Eft9ssH26eZUDBS9Pg2InKS6fAVj68I
h8t48NAwgHTis1WBlX2xeYMCtqTHbvur5QkhbwZjuYKRBGvqdpa2bj7HnRbdxpu0
XFGVGGZw8qJ9Sr8YOUOF6houQ7JJir2w02XBYfoLfQaqC7ZcJejGiM43lnY/KX04
NEoDTtehBko1Yrj13pW1w8/IZUP5X99ch4hJ9N4umb/Ve1EIoZ7By0twMqYLpI7T
lChRGyXX91U8zAy/GlALn4HMEovhcUtY+GLuW9cxw3uh/5oMXYxrhti4NP1QXVH9
zyl3zOoejQvkG7yNbDjuidrs9CRsSsMv121InY3QQGHIp3OqObnQhs6Do7rrKxfJ
UcYaXWmAYfYuTM5g3GIi59QgbpzCtk6GYdbgnrJolOFvW3Vc9p4aJPtG6Ur3MyaJ
XxIhZ23Ye/VpVlbKtw4pnmHS83l2C1voqL7Oe3h+eJh+q3V/ShsVZRqTAKYdZbVh
Nr6NjFxssoFcDbzxcOPgxyUOVrF3vFQAj0Gf3OQdjMEnXyK7BKxJ+37EQK2ZxXX2
/l0+YsWlMbQ/3d0TO12o0gdCw/thyq5qq0RE0ZQvK6WbGIBryWfViwrZqXU1dHMh
LMtPauluX0bD+imoyGoDmOrKYGPXqUiGcNhsz8M08L3xKxWqis/ay+8nEXhW2j29
W7VHuQEIO0w0ndGJiWvJaXklkIeJs8LrSI1aIWsgeUIkup2C3XYCBkf0aLldyIVy
mN+cNv7yLxauQkH0iGrgZ8mcO+i62P60nujVRdOJkC9i+tJmlcN8K3tG6bOyqWWU
RIZgIs4Pgtezu2vQBHTGNgf31BN7Ytt50c6PULuYlkr3B48rsvBnQJqzhj1qCaen
4rv9Fy96WPHGG+hwIzaL5ftQrRPAFWahUx6xSarbJVICusJI6cuScgIei2Nxa+FN
UVQQZaQaY6/VT9Epc8LCyXSk/UII7A40G3mEdoUHb/8oF+zaR4+wf96TdPzqJnxO
U5v00xL1p1UTAyHyXtisIGqSZit0lmZAqNoqg23ji1dZnSp9jE6jmh5AUH40KT0W
CoGldL0kUQwh8u6nURs4ZUBBF4kc2ngGfqgqeFJfgKtqsrtH+BySiiCPzb+FH9HQ
pMFgmxnPC9J55GYyeFAyTeK4iCUcrYCaN+lW7LpE4txF94lSxaDQ72OISDAmimmi
35jGQjh2pATtVIv9BvFi0sQvTnhoofT56bFQlzAnGJSJUaC7rG5SA6LOO91bf5DU
i4Fiu3FPrvs+2mfQ4a5TVZVoGincMShF1KhMAnoc2WugupjiV5g0QeioV1hRxBz/
BdHiYtbhIWflIjhgSGlsmpoOXf8J3JhJRccq1TbB/pNIg77v8nXLt/Op8AJVkjdz
Y8272XQA6ZSS5nGwb9UTpXIV39qs39pYV1+4vd5yILO2E1Y9Yjfw9AX3883DfVYO
Ba9xqbWaeRe4ny8AssdUHKAqMTO881hzZB4INwW99YsOI1N3sIRfpSASHpUoVg/l
ZRAObv318B2ROzlwa7CZb2XX6Xu820jhn6ulY9BJBAaHvOB3Z1B3NtzO547GScSc
fWdV0tikbbGuRGRsMzjxs3a9KtY6QZ164vayesxv08b/tXglnlSQnqWA7IIdbeEz
J974tba6YUJgT+fzVfJ1RB+EpGCRs0UzficTDpg0oy7qODhMwCSUCW/A4onwm04b
yme2wGqZ1RyjMJX6iFXJEDyL874NA4hn3pVtTHAlhiNMMuwWZ5A3IIpbU8hCFl9/
YS+VTHlKWJ1H0+ibuifwhE3xKyxD6ddTLleGYAAuqIELJ6kchj491KUIF19mc3Z1
zvXmx9nMa1COcmL3uaw4GE5wxbIkDWeL8qrSEl2NBzfHnEVHGLPDoNxQI2RhzsON
g9ZZBap08UZ9RmtzgjrTkMJPSlDmNthALs3EgBC2816XyDaT1owdROa9UzKbtC4K
Umo0kTmjVJV1SoGdttTRSMYHScTfKd9lrB7A61mId6JKHeh2l2PUwgAI9wbz9+/w
oJgpOLmcYVfIgF16VU3QNEQTXMPEVzyYfAskx4uu6Idf7PN93sbC3Q+fPf3n4BWA
st2+tPeLHjI4HORg9HPVqghzSkuxQSKUwfpkosSfDEpNQPS83EbTc60BsBKt4o9S
wcahcRSjpWOHxEm9i6KASOITfciYk/fKpV1XhtMtc5UxeCf581Sdos5bvrurPDCq
yBK2sQ2LfaqN38ssnXuVKheXEYSU90xopdQf7/T0k/Ftd1Ab/TfA00vK1jD6qO15
UEONjB09OzC52UdOkYlO4u4AIoaL4LNITi/av/4/fF0WHx9ANnZgP0wAwMLbltGE
dMx5UdF/Kppnww5/FxE+tLHsG3u6yh2E7mwFZcw+SPeLmZa+HCeLi267uDjhr+E+
BNyxgu78/s4kQuUfly5Fmix1FVcr271E8cTjyMlxY66+Q0lhT3s42bjlUtRzpR+w
Jdzb1LzLwLh4fZjvL1jmpZmw9jPHYY4il53aNKcXKEA5qwANiaBiYhuTEiqXrXkV
TEVYBV8M4hkdE9aZkzbIi7Bff2N/hA/PxOHmOuqpDUC1ziNwbI0O9RwYfVbDjLZ/
Kq/DPn3kkYV3UZj2d5a4eC5rkj2OzWVRnU31cX0I4IDzV9grzoooPL2PsaFDxjN9
Thwq9zLlZbe+V3Fgc+fflV6VFOcTjk4pAn0unv9fvm2e/L3119Uho93MjwYI1uIz
k3UHeWC8yPFo4iWSL0kn1jume4QgZ4ETpOpFnoKJHLvPvrZNfohfQmeQeikTsXX7
IojdiWJTzMAE5pmGw5AD5+2noYSSpMdCk9FdoNo7cQQ1V/saVTLj6y5Wq3MT579I
L2yR7gYJN/mcCm/7YtqG3I6pBEPIbMRKjgZWx3Wu6ielGBURlGa632ncuj37zLou
Swvwsy8nMI4WLJ7q6al9zVw3tkkvMz4qnnWJdIw8pDcc92JdjdBHxo2oUXaYNCQH
RjSzmltQD3qZuQmNFMu2qMMGlKzq6/SkiRGp7+RQgwq49t+QpV0sRqW2jkA2GHtF
ogwaDnvgU+CIBfgiJokoCSBZ2JZUxmj42cFU9H4kbzHQDyVXBMu11rlnAH8TMrBU
h9+c93HTOgnx6/fNstOnDJcyPsiZRbDIDlOLmRTHod6YsHgi/V6c3Z/EtWED+TDI
6rUZl4XsuYFSZuybnioGnYVTX44A4mzIXnCpcICp/RrMpsoZJ7/pgqSR2pecZtVY
LHQ0CUuAYYaanDs0rFKPHxVrk0AA6D4ogUZO80UTV2pcJsEazTwu7L22U+rLJycE
5X0aofyNg+8u+RMODRKtnp9zFlOGGXzYkF5EgytD09wW0xoexlND2Vcdahmn9pQd
+Joi8x1JR6efDMiulmCzuKpzxc6GvzKDus/qcyJrGjvJ71rtdFcm5WTweQht7Tmy
wysGbkDWYY7oEN1XL5qMHK1B2AvhPl5NIN1MO10bjZZf79n8CO+ULSzk0i8vC8we
2hEY3k4cdtn9k+m+ye3tul2v0a2RhA9Vist30B8GrGjhD33hA8pw4kgwA8jU0FRo
XdIdM3gky8CpGuhbsyLAeQMORZ20yyGblchinaewIqt2Jp7fa45mK2pw1G91FusP
Cve2iNUyQVMMabHXh0xXC5N3HHQntEuKizq9Ci1boCwWmfqxrdMXaYlZKtlWXK4k
Xoq2zF727eWLplV2SUKVZh28z5ezQ40RaVc87cRzQVtUjpNjDUTqyeBwneoBim+v
M6gTv5GIFlZyUjFCiPnrKpXHebmQIs55XkHMY2QPEMmZ30Ge0Wq1Ma4AvdXpS6Tc
2qrvSC2fM878hao5O3IrkQzW9p7WSwB7Bpwb43R+ELBHRL/LmViBnxMl/TL9w0Np
Cqu2ye9JVc3bDOV03ukTrgp43z9UCigZuNngtF9L1T6C8jGH2jqJWYICcgj1yTmJ
or7yZUWT+trIpy2loS9jZY88TitjIp/Zpe50KEm6bkZh+zfgA2sEUmR2SazLvWPO
9+Oh9doiDSl3eY8KIwJTqLckFlVrt62IwNEfnaVt0kZRnTgyQpJbZPMyYUw4AhNs
+dOMDVpnkvU89cbZwnLQw7bRSZFPrRqQn+DiUl/ScM8qR3tYitG8W2Ugdzvec3hr
uyvGZwNrA7CueaktyhVeFl+c1TSTWXzuyJNAqpB5Elk1+RQrpOMDqnG7Dl4wFmRY
A/WHk1o0GRWglagIWB8v6VL6gmiQHc26RisKbEowuSrKGpe3WYrNdKYrNLti/hiN
A615po0oW5hHGh1UFnlqvwmk2VRNq025H1XuoZL90mwHiidT+PXpjSF3dbWp3nMp
XkP0YHOao0zVNwUJJAKFZDPDxddwCDVQ0flbc7Fw4t84dfvLjxm0NR5y+0QmlFqE
fyOUzn/BDrUR6W0oDYCoCnL9/BMR/vDXPdXLzCF5Z6+Bc0KaGSF1khKiwotx4osn
caCKtEZhA4pljrAAEikLe3oFs/1sXbNyhwB9dB2WK0D3WSQE1IMQrOFDkeM5T+OL
gZJbE/6WC5V08aWZMW7lvSEqAFE9u7+q0zm+7WCHU6CggqR6SPA1clHj8D42K4W5
BGBzNagWdLkdVICyBK3nHzltfy5Pum+C2X1QwuwZ0i8MaBBDYPWbqAsnUpUIEF1G
YGv30t5ciXt+kwlOtS5BEEIW4Yo/UTmAebjUsOxNFwkMFRhpvmuYYsNhenxI8ET4
KLawpM5G438hUdiZrt97JuYN+lzLwknQi4wcvdgPBU6RM57Q7aBnFklxMOvT/vIQ
durc+tiiyuZfq1u6NOun9UmdGJOaW5WPlrwuoce81w1l68/rD+Q9nfIJYo4nfdqe
Ywx990l6nhDvF9hNapiBsu6dWdKidjLChzRNzUwpCHr0wjixIctZMdJE1GH/LJT+
f3XP0fI4NBQ7spmsMLaz/ui6C0PgiHLneMRwHH0g+i9Gv+RUHpuP7pk70CCdebFo
6JezNbEygpD52oRRo3EfIiBX3fV6ncyGTNH5fxFJs4NQG+08hxFYblD2FKhYyT/x
GmgtSs9ypT112Kw+GAFFNhjHjkQwuNdqiWmkFBtSt7khxx4mVD82Y0EnjXOQMhb6
4AZ1jwajStu6kna7knKTRsSxEB47ej050HZgesxPGg1JFBl1J+GXwMrAfVVkifBT
BMDwQU2sF64joKaYkn0Auc1A8YbPs8OJtfZEL+vZB3xQCD9pBG8kh12yqTWgCDX7
MaJVm55+M2KGBvEZ/pfgsFFM7QFT+yLij7+uDHb1+kcM+4Cld5VnTeGNkVwMuUDf
B5eJGg/XjG6UmIgUxOiFGDfVADU5WyxAjCiFHXAvp4gDfPK9NpJIN3XXvHaFSGRI
Xab/GMAIbTg92y0iDnxr9nQrna4zN5pwxj6lgNbHvw4pOeLJi/le+fwN6p2pMZ3O
OzA3tPYTsn1jyETSNEpHwRzWYOwQRTF1RRLz2VeCnql1GCa/8YJm5pDGcJTG+max
VxO5EWycJRgxH/fU7H+qMgGgRU7LlkunW2en7S1a7JJ7782iD+2EQebA7JIUNoLl
+fu+vYymEr2VE7BFxBpzYP1feq1YH0w1oDEchH6cWLXSpMsU2ZeHdi1SCXkOYw9F
f1ts1SFIH53f6Ymo4/bgX+9mK77wIjSvIqvsYl/HRPVVLe/yq+/56d7aCsFi1i+P
+px/OnFm7Pva3URY212oydZMTMD6GBMKS4ljVZ87mgxBJpKRDtI9UMnB5O1ab7Ca
0CIAldgYG/Ueq0n35vRuBTa9PpDWOz7zYXtRLyY9c9I8+diXSFZaQzUjgQsNPavH
/hPHoasglPBGCbRBUqfOItmFO/6KxSuHJI8/3KU9nFET+9O/IwkA7qPGOoAlTBmS
Gg+0fZpa7E6K+EhD1jahDYY1pib29KTEXOcRYMvpsJysirkFeIsIK7C7H5xCd0Ru
S/74P+e9vPb3z9wvKabvNI0Xc0hzQsifvM23M+c/f/rdp9Pic+ceDf6mkTlg6G3R
H2UA9tr2juJhViu29c5knAHR2aLp3IpmJylLAspAl/RgNks/S5MIjHcpPbXlY2w2
tejf/6LYmPsFmciTaeu4jGB55FSiZykvQThuc2Jpn30Gc7YoK6+ArHsAbDixSxff
rspVt7QKvpPD21Fp6uO2DbbPwI8BzsP3JgCQ4UOlrOchDqdxFunTDBqz8aQg4l88
Ax6GHuYbdqUb4KLDTIanujZ+iI6GseD7Scc+/KILo1rqcP1ximKTOghp1gz98+GY
2BrupdsgE9HKT+6Ef+qyD93j4IRiIJBrsrclN79RUlu4/eS1/m/NCVAsdioam/UG
gVqOM3mpbTKybdl++Fe/Ot/HecRwb76AcXTpHkMK6sJqBCEoV2R+ORP43sFlxIW9
tCoj5pF5IQDQ9o5a8yEPqUtxRxOkL8YMqEvFnKbMIZXOQaGnKjkihXV4QslUdfMx
If9TrRP9u0O+4MM5t163N5uTI49oz2KzqArhq8CycJufEaZUL3FjOewLFukLJrOW
RkFq43SbtNRRIweYki6CeI1nJeSrvc2oaEKsVnS/nb3HorlAXKU79hhD0jWnEH+0
1NMLgDKX6JIWBnfs6jzmp7nOn8Zyy2kq5spCSyzsNKgnCFjo8WFtUlOnSvakwWyh
2nY8RVnDwpBFv8GOA+jcFqnagrE/KzgVW89An/ZTjG9T7wdtTXUPQwee+TffwB1x
RXSmAyZQDwwIy9F/fKSWU1Sl/d1PlFyOjufyMgTheIyIQYxja6AoNmHPwztkK/nD
RFs3AB5AC6wYbfStntCwiWFyfgUpS4QKoXyLUNtJpjdrajMzki7J3GYzTZwUWsMz
TsMvzPFMdc8PGnFSaZo78Op1uGAVrSCl5Z6xDrHDW/u3l8kfHSzKkSDsTgNqgQjh
90/qQRGugfw4hJJ1bClEeCcyKWYHGX6TMjeeThqJZveACfAZskmtu7GRwsFbqqzK
m21BmXw9eMaOv0MdpEQWDB2/xG2O0gluxmkNQWkGuPDvgZQgn/dsliR0pJWSaM6U
2kFoAyatYu9hkt2Gc3zxUYFMuJZXwIX1rbj9bMqw/S7aST4OnbhrejEEeInoG8/z
tOTbzrXi+Yzi/j+rSPHzm1UrougL6s/sEi6r8yUI9frZVvhdea74XfFReXdyYRpI
3VT+Tdv/T1DNBaxl2amaFvhsbmubfBLrDRRK/DxccBBzR0q92jrfXlMw0Iz0WC8K
Y+cf1xm/lxVm+od3RfCKbX8Ekm19hNFFJ1rPNUBhrI6WGI6t364PMzLXoScQ4kWF
NQu+hTxbUe03AsHl6OFZq3uEAJcYqRHwCqNQtceOrareQf9xP4NaFjBIhOkTnDgX
kv3qosB+pQyxi/lIfCwe3f79uKzvGO9q2gvTun56sWm8Zhye5i5awO8zLya3agNN
wItQ0Yav9dIndcpwwyh5ReEpcAKoeDh+/ZDS//jdTsH7UCdfzQ5YXfrEkyEI2kjR
PVVQTW+vo1OH3QQVxN7WcCg5DKSf8C2blAXtwDObMrqUKsxzNlQINTDdGjV7Mu7s
Q27JFIm5oy6s3qeMAhIKqyVf8hnUFRWjZtX5vu4wBgarKFVduoqfRjlvZ089Qskt
JOFMeS/vC53tKy3Y2l11y90t0d5jvCJtU7KOsbMZFfDL4RhxBpoGFJDqPdALWpSa
zUakhohrjbQ0MjSYlqdjxqiOrNrb5nkYA2EiJDz5GYQbUhkV7hPf+hXenRoYp9Ju
tBO0zrIZIhptucKdtjon6OdpR/g5nvY21aKMOdtIwhnvDvNWoXNrkrcUcqJglFY8
d7+iIGOdtfW090E3h5nn9DRGzNdqTevlIl1+AUX6A3EtnfWTGK5LxDJTydC2NJAz
+l+QLtkXPgXz2GlR3ZYIfTVTRUpuNUta9h2Di97rbM/Or0ZfbZVveoI4RW1hyn+2
H901bul14O9vcr06soZy2gnq3SmHrcYUWwHq0PoXiGmAwdXBG06UJdBNIIcTapIK
Ic0kPBy4YsotpIDywLVH1RlCZxRW1KJM6mnLGLzS7m7szK1b0EafzFuEOUJEkkaF
qJqLewnh8OtI+I1WPtK+amX5YfUPwyTLR++qGqVA4497laVFzzsmJH1NhKk4PyW2
qMbKXaGbNWjjiEHvbRNMoDZ9OAeD7ceAhdDPDRZRHKWKVqPku6N0nYXtknT/Lw+l
k4eEyfEmdo/hp83srFKbObZqgIyrr8Tgtx+m1xfDNHOVkq7pgzXTy9J6492TP+jX
hDIZklj2mmzMSxzPa0RZli82nUHSvRo+LZyg5CWiWq7s8zgcVt0vGJhRNZNwezmB
0/TUjmNNbbLHOsdhJp3JvAE9jhSz2ran9aj3IxAPX0nfeEbcxWnZHn3lJ57WMVul
4HwrVGpT2pyUsXEO83aWsDrudzaTDn/h9Bje84HlJfKElxfz40F/zorMewIJx5qZ
rxrvGTtI8FhyMzeCMRitNmgiODOoYHXxf9Eh7eiUthENV/vDPOsmL7JyYyZZrVA8
6A5C2cx4ZyD9ZWnWw3CwmL03jHWVUOdA4eBMW6GkQswj6x2ldGwr93xGH6E9LRIB
3Xe89MpsoDBgFxZQJH0DXFBywMmLBvaW247H+QawDeShAXx8G/dKq2jjPjrhKdB/
Wc6Fm73FlesIpU3DF9MSVwqwBHKTZqx15JvHUinQi0MTH0BLf4g0/2BlulYxvoM/
Gn+fHGCz7pSpCC8HxY+KUlsM7Q/vvjFS7aXO3GqhWS3oV7nxxQb5H1RwEQeV1aqr
Pc9yz7sawgx7RSCwpFgSsROgChe5ZisHDwh4GtqhStPBnB9FtC2XcGxjtpO9YMCn
/3zwYibFRFXWKJ9aJUBylZGx5ag6iqXbmKdFn4grO7Dg8QOW3cw15v6gXqqLIepo
a6AV4zzaSZ9fDN3JtUwS668Ivl4WjLbS2ToBZWwseh69EgSUVrAv2llFXtQSWxxO
cr/drHEOTV7gh9/X9llWt8Jeie5M8+zPXT7W1oAiEfI+5l3/qdiMPRBTvOOLRlbd
LOrzpEKsJ950lxkuRixh+t/vvfIP9PP4Kr21hpwYGFHBJHOBI/HXWy1KkP5JuehF
1g8wEqYcCgbOKI+0fPrxvk+kAj1pXT75BEKH5LPG8kHW2OuIwtzoYXL86xCbUm+f
KZICMbO1cIm/44Opz6Pk8AbVYvr8bIBcWt+FsDeLFnuXPfWk8wF0ZxA2tk8HdoZB
D1Ucj2myIUKa7Y6OEwAWwWjyTuTgfZfowdR54lyw+BHvODAqGnxL1Wbyqua/I68S
9ZBRbo8nzfDTkoP5+k2v28ML2gA9zALIx7JSIv5ZYv+wf2IXISikQbtzxZlYeCuf
niBFCkXh0PermfXqIQ6pDEWFQ8pLf5nPElXD4X/gaML98g1O6Drxl4xoVTqmhZxG
JzLc4xGvze12eZuC4c5igEQOE41nGXs13IPQSBefk7+WqkxxdtK4YKi489/npedi
1gu8YL7PGAah/clLfcdgdbWenDzy/nYGUtz7PDpwg5G4ymAnXTTkZ6bhUGSImKj/
ksJGupT5bGb9aUmQqzkljHERaqiK6WhoYDeYwx15vOuKt6Nqs4zUSthF19ctrE54
z5g+sqo6wPPF+cHZ3yBKszfJisDWHFzG3wn0OLhyGtltd0UAyVJOAVSCYcbmmO8Y
yISszLfBwrCEa00MqtqbVpFmGzWwsuhgQIh2Eb3njOtMBQeytTLFn/C1/UnvsFSf
JDvnR9kdY+ZWlIbtw4NS0sEJagEDghmNt4x6ZCLiZfNXIbEizJtkcdVNcQHrblXM
qXthoKPIgS5KiyHzquVFtj5jpbCAypi0KFYNXrghoAk3G04RRtdSUgRSEiuf/z4H
p4vkhj+NVen8wM1n64Mb1AiTKHUP4CGzXSzeoAY2qfkKWcjOEqYUC806FeF7L6+x
A+1HGtlsSIufh8C7mISch1UGcHjjgZ329qXszCOJf7LSJi8VQ48Kt7tqpezV0YVP
aIbn8xuAJrzvN01ExJDVV4gEkxjOUplIUQuGVuFoIn0kJbidI5LFZ1Gx3yVB8ogv
5MAUbqEchWzhFF5CsAi4Hp9cBnSWNOCAK7xNY8drnbpBWu2UrIgocmWGkzrekSe1
Zikm2oEKxOIjcef6Q2XkP4mV41q2rwrT75+RwZz1tRtbQtSjv4Pz1tIzDu//Wb3S
D3RFi70bvl5C0v5TfFgqVFEMa0I7jyOfbHH5rHr/XX60Ix3CN6GIV8GLEFE85/2c
mV6cfE1kNCNPhfG+VwaEQmm27ugAumF0pFJmSLOpDxv1e6IYz1FfDXo/6m3+wu5n
2hSD48cnbrGM78nNJPC2ytIgKzKMGxgXvQVQy6+cHPvYJJ8YW/0fEVp3IDI2Hsg5
OyaDaAnxgT6Q6nK7ehSB50KOac6T8K7GyWvxQ6BYzY1ldlFxb32jfH9Ehr9iWwY6
VHkY3/G0/pYnLJ/Yo4lBCQTS9cMiIPyrrEQ73WptIHbvUZ6A8ayOlRMGgs8cCghv
S/iky22bhMSrlZ6s+cX5hgaHjQvYSMxGrmao/y1zsX3PB90nvetbzcPZ8NHDp0ST
P1+YSBbPFj8k9UogUXT4pYmVG7QKBTAMK8K5XBmxdl49346+gs0LZWAo10Cnk5qo
W5BWwvWcFrV5d6Hh2rVz4R1qfmMsT+nmRf2ijIJr3KvCcstEN+7/l9QHn04G2LZV
WbRNlNpSFIASGKAf8s5I5TCv4XJkYNHpTNiNyYrAXN3OThVUzW1uoC9rnBOyjl1W
AMsnYMrZw+bR31HzLUHuW00EdYOOYmbZFCxfAlxnVA7Kz5UYd5M/NG7Vhe9aZ21S
ncg784Hxd5l+GObhFQ3GrwR/PXGbQ1GREres0WAI2xY5TklhLRzOdqhYgGwuyStn
GNobMt2/NpLqYqCteBrlO2ZAdVGwTMej5evCDmewDMogFGoCOH75Kc8Uuj514HxO
cdO3dtaXdaabjBSNkKHdtlsH/HRg/6kEf9yyWCqz2mNR1gdy+utzW0AR/iM3FPCB
CPiTkDNjdEBi2+EqgNLn7U6EgZ9+48mDhkoptlfzTcp11vQQIzwpH98N9EbNJK5u
tl/ftos7+Ro6O4SiKRUwcjSM1ISdP40bOn9PZHRNbBjH3glNDHjpzK3EZQDpYODK
utACucbos5H4P12oygNV076aZS4KXjV9w4anQRUE6qHveJIFQvjRAMkTAqrMT6dN
3pBjzFuLevJUMvos8PukI6f3Bdnp97YtKkpRYHUB8fV+E/PlTSJWlrTOvcLzSfdC
REhFHsMX18jOSAwW3sTt9uZsDY5bhzZe00ijlUHUVOVaynm1xtJ6KwRtRoWaqNNz
TRYDnc83auWsjBrQYCftasja+ThZmIVbYZ7zVDJ3xI34Y7JwI4YSFaCBqdOWrUNn
8LU5H+MKMmnbsbdYH4gLwgJ+68ic7lyCWdU0RsC/QhLDlhiLpqFFjXFImD6YjgMr
EBjnuXV232R7X1Ykv/key95fY75GqsuoFXAn3o8DXy6/YF8wXLbmIwJK4OOClydK
r0yeFPattCmqDBZ1s9kg8Y7LisOH6CkTPnnS8ezu8UjJ6j3HcOwl442cS1xTpPDT
HZtBtAGo6DnJvgnMxUK76Mv/DNfb1ZJ931A3VlZZHSRpNYP2NnvHfEfZfD8FzbkO
hFXvuK48LdGn7QHCX10nMrh4q7GebuIV3VmapGQxrZ+xVr1YakDKhEw8YW8/nT/f
GDKgmCjDSkFq0RXf4syr6hhM0yaJwn68sxj/vyeSzR5VrZQsaGCblfrBrq8toUxX
rjIVMrDm05T1tb/O+bnOHC0z1Mi1fd8lMFvosmIpkz8D8rg0Yt6/UmzxofRPHbTb
rFzpl0QXCXVw2U5qxngbgc8q09YL/LPKr/vv5XM2xjHp/s5Iu5dAhX0uBRsX5IoY
llYdpPMQgEujvc+V278ZDEj5jJ5K8VT6P8bm0XQYTiX29MVYt1rEJN314KRpXCOR
5FoYDz6NExpcqtSUXW5YPGvRYvfcS6A8Vcm4zaJOl9UiB/ka4sjv/qP779mv1DPy
lgXrfgH+YClu48dv1cQ18ChyrIzA6Fl5JTV188xB5yp8ua93T9/jelenzgWAknme
rFMHTWH4O+N8O8RbeXrnwE6TUp2rWObtU7d7Xor1rbwqqRxLE56McD5RfIZHKvWP
sPPWNmUiG4dlmAZGkUUoi5BqV2SCAvg8vNJ3EIP3bsyCAk7WBpFXbUI8yX7cKWGy
xeox5LbZPFQDmqxiOT3TeIjeG1qSyvbzbpiyXeGm7EAk4Hb5ZA53v2MFQ3prwc1x
UV1e/52x1H3bZGHH8HZmU4+gGmKx5adGNPNf9APfBcagMC0ayRQ8uYB2zIMXJ9Zv
0fmvWpWx2OmAYMKxi/BNVidOR7FLaLD3EpJ5qQK6QRhIJ7bnKd/TnMyIIfSPgeKJ
mjqGxqsrqLQryWU04NJaBelyb1CMPNNJoASAblj5nNU1oj2+V3XR7rl8/V3a/HAn
QSdxSrHinj/aqQ9D8JuZXvFEb6KnLvRuaJqCW9Bu4DjXtaPyAh1IvgL/RaVq9mSS
bzQxbIg9R06oUT8DOsr6av37w7TaQTYnygjFEtljasgFH6vBeBaGWPkzrfKL+pOU
UJcPqSHbXdb53VdYWfyPD/bUKdB63taKCHKew3EoHrcBchQX9bNYlU/y4hPplhVd
r/1TkK+5lg/HtHyV4LG/iTNDUn0xNNpCoe4KC0muHpfWsfp/5rKfL6ds7UxPGkHx
L1B+nWIVr10FjZy59sAZ/KN1XlwiA904eIph3EICLM9mjejuDY2M/lav5sepLXh4
lav6eZ8Ti9c4V3SwXd8PtTNalHznvdaxR5Fsz3L4dfkoiabPtcGQTaAVmUZ05Lbt
cOOauLgaf7zUL/L+AII10i5VYXjo0lLqz0bSRIh9pzQ/LWPtDWeIIcYNyNvio8MW
0XbuB4l7+AZsf4Du4FEHP2M5mqiq4OPISoWLgdNzcsqJAc0YQTPxm0QfHgsek6Df
p/2e5COBeTuiOpblX1r3CgZ+5bPrcQhtaQ4Mw692lgayN4d8PUenhVQv2OGejtj8
YE8YJwFfBR6qZrcOthnykNa72ZB06YbxYqp7ORkOVVxNcWlMKtHpAshN9NfUdyr8
rTuKe2fzHxWmknF6Kwl7k7p/YNXyt+b3woNuDexEfO8D5RNd857TMqY+DlkO8AKh
N+PRJFxgEG4eCA/PVgGcZOGZSzFYdFV2msvhScyLz5aTOn+af9/BWrEyCv35PJN+
kGxxb76KvSEiRqe9cHiYeKtqeDexJ4Le0Fpze9/uqALXVc/RzN0ZEQnf3hPKBy6D
dd9GiIjqK1xI3C0CScNGiJGPkf6GdQ19lbutcNUT15/HqFfFCTvYdyCb2R5H7kKS
l5B5jBuJRYS6Vrvzrs+t4aWBMf97x8fsHQl1RUv1cRSBU8qg3scnsWtDXRPdWPCc
2mKN2hWlCZ+81pHhYUll4fvT3LSke3v60RwxwUvdRGcccyeDOX6z5N8wKlAO+ElK
MVUDSnl+EOkVaoWdIJxW9k2NNh5A1lmIY+tmWfOyBRnjwy2aRQrsoj2Ztk2/u5/C
oUCa19SzhSys9oSZSOUplqmHE7Ibl7H1D6h1NcOrSi4L010503UHiRc/xN1xS2s0
/GFVsTBEPvuwA2z/6aOsxzMjhCyCbQ37NFSZzkocIrTqdJm1E1RWEK3wchZesZrY
RUyRv+OZdZmy8KLuiS7kqSnHz7cSGWzpBTAcLKXXADw9JUoR/1HEhkl8bxVjQ4H3
4+mvnJVJ5MtCR8RNQfNqBbgr9VffyCdz6gWWqCbIZQi4wT6/IU19aB5+MXSyJcva
48fU23OItIuueq8nzxaccbUfHsOOuzyWYlZaI057Q5jHgvoBHbUCOtPEdpjLDaeJ
X/8wq9IwlcFaJRPPbgOpl/b7jrJd5lStCWeu5xWJrEcvBQxHWiazyZmqo1jziRCg
r1Hl0qDjmyecI5MQvHTgoG8WTyxrge4+3iiEWnMQqnuvSLg1QWB5B19GZz82k/pG
7yW4ig5GzRquwFZf36PISc53AuckkbrsuDliQdDfmaX90iPjv1AAocYC6ADmI8/Y
1XwZ6MzM91S5VweHN/GWZ2J/nOchiHxry5cENJpU6EIXetZutb5T98XUzk1AB4he
ULFPodxuRQHWuZTi9oUwmVm+LUwIikXFWdXgebC7WCmCWAG6co4K7/x8pFQomNpF
7dQOf1AkyL2SWbOs7jhKOTj9RNJMpmlLWpJ5Xbxws3Kaht7tzSGW2N35wIKqTQ0X
iuUk7mjRAjivh4vUbTcuKa65o+N49XwJPjr3ZNdP4WdMta/Pl/8tXXEK7poyDMwR
UHj0meRbWfGPULBFaXHhuykLTxIwFmzEeRWEiYm1BM+GiNe9HfVSP9669ZoOeTgq
BpVxooduFdxfmKBQhoS0Bf7+PtQca4B/L+x0QjxNtoEkQqygDdUVZ+jyFc4x7uUD
kLjS5BfSBNhy7GJjtjQIWxgJQLPqwg/E0uMrUb34uNRonLtqtDQRt0xIxSBEGQXV
VzSOLDXEd82OknKVbu6EOJx/hT1JY1qyE1tPAz1kgqyetXknZTvmH2PWb5Ubb5h2
+YwY0zJYMu8DgY3sqwtE6oHWGFl01ofZ+X2eEEFiv87MZAWLF/55WSAi80d2NF/A
yEwMHesCeYlqOlklpJR/JALlf8LgyKwvDSxck132h27t5WyCDbZikgPizgDCTL13
isHGZjfeqo2MHCaAxMZgBVjZP6KjrpF+hebZWf9OIjWVAPDnNo55tCtKGqZ+wrpp
rlN1l22GIBHTd+v/yabXASQtB0bQ6g4s3J8LqhxZrMJo2/QRf1oTJRT/zMuqONEb
3RhNO4L4U3Ey1lB1eWnS89XY8mxFJJKWivBteiAnX+WvbLE0Vh95Vxr+CcAa5wkr
7JQo6tM8tMZLYbocb+YonRL+xgdKX8TaUuU37O21fOq2mbyIukUpPBujKT8nL/NR
4Pj7YkCJgGDeQ/LnV3AGIBeIFqxpU5R5JP9NRciaz0YeoAG6Roh99XQbCs/sWAks
vrEnEl3ro+cLOxtKLqedqxCT369KnkhUWjTH8XZ5JSRd6wzc1QYEzdPq3K3g7ZvL
WdQlm36v/TPWnD70z+GKwwjigbK9dQvRkfgbA6vmpMeRmQYLksO2tZq2uimhdROq
ra2kufrvalWPAizMfL8RiwiDGqGnjXjluvLcvje7uy90IPo34bV9/raoI0OJ7fWt
SKCK14YK7YfjdXT3iCyn8Fv8qeHFiS2PZgx3w32+axI2TH1SJr/jDrGIyLINEfuu
HhIrjY6mHJBzG64zluzPWhYS1w5tWrNeYlFUeuM9gbvVr8b4ihYO22n8JP6IxoLR
cxfrKuncFJkPmA3woJ9emD5hT6r58UKfxwL4nL/TLYEJIOJcFbHrOjAFPP+89oWq
6AZri1tkrQ8WVkC9ikCg41s89b+2CCMDZLFwuIlw5CHEPBhvsyGQcWjReM+BoFEw
/GtvGHVg6j2WeYiZyIOYWZgZo9oqI4otQjtG9qrLH5g14S3APPYJRLG5qz2pi0fC
ZH1fthCA/yDNfiKyma8rPhAziQY8wBnJBZDahFuxpTzB5h1npgPB0R1nf+e5goSX
RWz0T0/k155k3VAVWcEXi6BnnmQZJMRnENh86KIotPmkzEH9SQ7488MqHH1RWP2Y
3weroRxRXTqSJZqDYG8w2MpiZ++L3qU/09jcndUqKuURXnuG1+PpMdcJmttBmIP1
TbvOTTwf6B/Y+Epg3Oq8JIqPu1Gsqn47Tiq5vznKCVYfoth8bOp7lcn3vSeu8KF4
qtLvwy+VNw7XYMkm+jf+4vSPHPPkJzXRAI0gq1ZA0ylrknE0o9dbb7ND1Iqm8zck
0/wGGoI6JMSB/uCMirJ0j7rOpwaZ+knGNk/nu3XizwfczBgVS5Z++k439y2Yuems
ooNGgOfwSbttALrKLFRmRR84WGgbG0Taj2c5DIoS6AqZYY/NqZe7UdG4/ueN91HV
jKPb+mgo0J5RX8RpSkelLEv6Z02I2v07e33i1XL7nWkpmUOYNSt6F7j1kH7f6DV4
nf+cJ8e4gMr2TgBptudtrTu2ktpPvFxoM4k1Awve8mv82DaLxs0FTVyRfAVGWG5V
Cebj8l3aY2Ih4RBNaDX9AlLONk1Z2c+Mlyi30GA0Bh6BigMHvPIge+LQm2VBaKfP
IW8wxpq2NRMgAYNOlkKQyytYAwtnDKAPBPHHV2WwAgIQk9WQgMqJCjMVZoHIONRm
GvqyoxHkjpT0NZmv72Kj8/mAIvCwpr/DZt2c4QN2fO7Ua0Dl9HVxa3FiZLeXxf3B
TXZ/AS1SWgTlqhSrdxv5kaUhRIuKUNhJ15lbbfz+zlIiYE93v2ERrHZer4cp+vP2
fvKYnKhaq59FsLVWG/K0dUmQ88G7BFVg3BOvTEyO3BnZUar5+IqBtYtMhi+J+0/Q
viG/X9WRI8wrLhIXrSWnBFV738HUVvf3p85XJ7E2nXqRaOYh66z9/gOdf84wwmg1
K+/uEvbOGfnjoWz+wi7AHbFUUuW+PiIPjWEA9ahoB1vW/1is/m28Q9/NUFZ7ENMo
a+wilir2otN7BOEmNLiJcY76nccvJbpsE9vazPodF05a79rjFb0AfzfNObnp75tR
AZRsuyE2SB7qapDAta8MJLsp167mqVAAA+hdE1teyRXn5pHRijjaceLuqmyaMNAq
NUNKmK4jOE0Q3GGfcyhZ1uDFy/0Fk/8+oO2TjRb8rzxaiHCSXBuF6o2UdzZgM/kD
GP7TfsBWkahYLKEYuBrNyqilVnu3LO2FaZVMvGVWb2tnazYbWkHgoCeKIefeZXcE
UhRsqlNtsz6C6J/wpAtgDQJQbZkz/2SAesMaiAG4+F/7QqEdKaJxP4LSTTwhexld
292m/Wg0Oh+t3luOS7DFa5/CEKStxl3+pIZgdFgnnIIN9UltZoAqmIL1/eUvyXTV
WgktFDvhSwIQJr+XkeQeoljVH/Ew5pe5/mnN0FATzegCazunKWxtn14qW/SG/1CZ
PE7mTVbZGaqUQr0pB6SsdJyjRCaZ7bWHuh7yxEBZmYbg0+OdyjyN1PO+VTfyojV7
R0LZJB64jDR/KC+ODBbrWIG/r3idSpzNe1BT4OqJMJMxz1E8qb3/WHhOLhCGeRzz
j+acjq9UhuluhmtAkHV5BCeHRXPmazLr8wMuSBCGmx6SVnVUaFw2812c0LB8yxEY
CbqEkoMynZLa+uuOVxcFZCNLGOx+fd00Xzwr2NQe10S3TJo0GDVmSBIPylICpCme
+ZlimsckRvizutBDGgSH3fnEyMjqlmeENtscYbcNG6j+Xg7LJZ0iL4amSxKTHfYD
N2sUoCLNxD+/OMd7ZjKjn3IdFvZajQWzK4yWn/6QYwfy8+wj5EzVinEblb/YGNge
8uU6t1WDYqcXB9yVYVAfpfadPkTzUsg8acPY4UeQHgO9sI9ERAeZftZvBvKc8MCR
iDvW5rwzRG8b3M0Ke3YXVXTB81zWRRAGL728sy0iGp8fk7toxo5tBes/AoO9HRYA
g206fDIn9W1fw9FxB0h92sI+9ylF/SwXTfOuWqYHFfjGOD56ShldNxr4n+53IChM
6TwnnkTrrrh9kFMCdpuL6tcM3HKMY/CAHPdE8jSWtfgVWBqBLYABVcrIIqfpvEUc
HIMUDxikPn1qYBhAJNhucJX3Ja/hl2RBkKhXmFt4+2vCRpQCcfwZRWdCOqkT2jTu
UVm3xa1jblEQyWwUkFalRtqs/W5XjRpoonLjQYshlCYefFTxJQSf43/kGAHM3yBN
Lg2QT7i48kFNjLRTyoIe0j1VwTi8a0UBP4DqnZ0DeV8GVuwxLD0y2wHCC0yJnLpH
mFmKZhCim35/z5TG10Usg28msWOXgx3j7gKP99+f34gCyvSc6yyo4Upce96cr9KY
yN22cUZtC5cCknZbF7XGWBADXFC8IudVFTKdhOd5bubL6IqdAaTbm5JZqlcBJRTG
ZWSMjJqX1RRAWimMrWmgLMen83Qc4sMVOnPMGEaAdl4lF0OTzalan5wAiAF+nOLc
9ByxUuDCzdwxMBHm0JnIKuOd3mjMtPj8gceDD7hTB04sIfVfhWVy4NLVoQKXPKFO
iUofRsVBUiBtUA1uWIhM3JjV0F4cdKnqRiY4DLJ0/+9G7TpDj84x4ty+t2mopzr4
q7F6rMt/r3MBpTn6rv155B53wWdYhyCgQcNVDYiu+RU06YpgO3yaFn77lY3X1V9s
ZfA17u/fDi2gwFArEaatEQm7SL5Z1zZnKWiJR3Mbs/N5W+ag2Uokcp9sbyFgeHX8
lamiBh5RSLIgH5Oe15/jQu2GniFu9PLCNwsaVkwT3rH1ivFFgWeAo72sc9yX0YhM
20kE1DtbLKDwyuJJO66tg09gRuhQIbK3TuuvfV0TDBFN64z45fuD0JsW8oVAYeLJ
6RJZBpOvbde4/STsuJPL6/vT4AndxBgypP4np4MzOCyFp0Au9j/RZT2QaIu1cDkA
2wITO27fmPAF3k/Fl0dMlKtnmyOklXBiMvqBozHK04ab2eLDPtMeOyhcvIDIXuhw
F8yGer/OxwY+HX/HSq5UHzvN+5HGId4HSH3OjTH7woIYYfDil0CW2HFT7B19rIxr
lXGoXwJGTbGRLaXONDdz/VUVWynQ+UViwB/dRsmMGOuqmURSGt6K8w63CRezHQj8
b0svmLueVtNSsJGK03QkzK5SO+T2wQdMUXEwqa2EqhgJzz1T/HsjWzplPw4xiSmF
NAmOjoFD+DhgKpNVggcqdjCol6Yy4x4Sk32xTgEFfxCk2lle0Dy42bU2/0ChMsdq
DHXtL5VaNNeNltbXFtYksWZQVm41sG/VrEmi5qdqUJFG3362XKDtsZ9rvcK9V/aN
nNRAp9cCQlmhsniPg/2jts28uHj0D1Iq6J2OQx5v5afsc9DfO3VpAp6eXQb2HqQR
mUmtzb6lxC4rzxl6Q/zJIkBsF5d231kaxJlnL+mFtZYyPphttD+3Czbpt97zh1QB
Ymd2TrH8R5TbMzEtVeYPJJTT2dN9cTgn/G1mQaonAVyTOAMzqCY6ahw8ekxxxuWr
WUQttB68PXrXqnwoxP+naD5hI1GsYWGO1NUzbfbqY08s79mcqn1fyGE5N93ecPur
UcIjBQhoEQaWDXFW2PUY7ddkG5J8aZlzpIOv+krVJtWockzV7Rk5yN5e2vYvESgH
NzvgIdLmMlYzqzw4ln45ZIiy1lK/z5fEbflT5g2S7MP2WGFAJ4bU7ir/cuJvk2KN
gV7rUnrxJ+ep/G+2P39y8SvZaC2gziQctltcIxbp/k46OJA6d1/aPlEFyVQ75dKO
jhQltfDJ26tbN3ZX6HtTEDKWTvW/cT1Kh+ZBtWR/1+PCvXtwCFoIvcUeogWuavST
k35BNDZrxRlLeehtRfgxa6L044qXLv53i5YZ3Q5tMCMK8Fbrwybu/7xjmZe+3nER
wEhJ88kwH+RvPlIglwRS97gYE5DuPlic3HO+nEbbSNy2NLUjQH/wVQjQ460pXCo8
KBz4aEzPh3iIB8sbHOw9Z2FM8Wh98GiuZ03+VRZoFz/dQt6hgckorS+llLDX1PlE
NW08MzLbmQS7vZAAG6vBkCpXpG3eWpnwN2KJuiJk3NP/PZ4l+sO0NSgifnNcH1cK
QIn75AxZJOkT9oCSoHpMTyrUMlWl6aJCMiEFVNmb6An2mjVQP/lc+UNoRqGt29Wo
IrP9npWQzSSSvxOFokVQSbnVKYGlzteQKXU5fo356OTtwkHyr/nZnDfIn8/P+Nyl
ujU6+qePEGvefIkBiVOL+Hz6232t+WGFHN1FFOA7PsfEx8Rt1EASTrx+I1vlNZLz
6gC06PZPHeZs0i0lPVaRpyzRWOE247/T9yHXAcM+NTJ3hn2Y281ksUIw7ufrtZbq
boNC9MlS7esOeIs2/be9HVG1IjapjvRtEELWzDQz+bBS/LAKXJyC+ejiUDXhDzz0
5YrSbDaOLpExYlPvkvw2VAHiAwGA6qVcISRUamoO84ykZy+CCBhNqpHQAmQddFjj
hh2QvsKu+GB+oMlunkwX42KHfYBpqdwQ0ZzbGAO+wvqqas/t+V04NZX74ZiinScu
6w+h6pEOQAZYcg26OK66f8JLD49UWR3pdUv/iNXMH5Rkrn9o1pOLXaCs4As4CBt4
L2DjYn9BrKaK6VcnrA04YrQWoXu3Hzfac/7BG0F+e46da0FKbxxjQp/LqAP+HmrQ
731wuRTGSUfp1KxSrwfcPrHX1tHKcJnOZYoNvzr9AnoZDncn5LDwxHRiomMacpzB
7KQMsVsTwvLjPQUZUSfJrZzFMd+ZPbyUwp5b4sstsLtPuz9GhA3uwTmA8SYfCzWt
hHRejUzXYjLF1GWYFvsL0100XXZPvGPpHbzXJ+jW3a19f+O4EQnf/JlpAgkrQ6uQ
9puPJNAbR2/kYr3CS1yLZNfH2SOtTfZCK5SQtXrNOBUU+E/dZ+kYk6IttlSny4O+
V8gkEjg1j8xKyxch8wUmHcx9H5m7NhitKyXZv3NK2tPoKbUxkW3ak1WsB1VgTC/7
tguoNKltwSsmE7+YI2gdd2dIrI6y/l+nsADw3TBMlnplRzipON3nZl1Hi8os64G+
QWqA7ZNvAWnXL/wkFPE9PlAUT8skGdN776nJI6q7QGTXHGFD0CrSP5kmPM0mvUTp
XyR9bKyxffBhTErdcjNn1ut45yKIVHlpoOMgEq1NLqmBnwEZAs+s2d7iX1xFr4BC
e03Rc7iwMysGuMT8YTvmbr5nkp7qqoyaks+5WuGTaruliWyiIniSrLlObULb/xcr
sKrqG/z+9AVTJViQjx+Q/LFkkoXHvQdGnL1hNiUFFOrVarnyhdTINvO1JJOdSo2v
5Bduw/nazm4f26FfwwuG4u9k8cKs2P+eAefrV0/St2P+PkGY47WX60LHIhHHXrae
EW/WdT/aS/gyTTeL+QDIPHwaELEbp5t1wVmIBOvBbtaePIO4t47W5kJlNnD+VqMV
kvESEzpqh5lLvvlQ3rVVIu8nMiyOT3PvooZLw/2vp0CgKGfswmN1HJPF4BXHzdtS
/M4vM7TemURrQ2gBtvrFcsqZ42nEsYMp+jfLdABL6CRfe1TeI2zpk48SlrCEzfQc
78Cgma/d6Lt6dZ1zWpSgsgOT5yqEY+h6q2F8YJYsPWfXCbz5km5QVu3JqGid4AjC
m/a+MMQd3kPHZ6rk92VxmrRcni0YGqhl70mSlUJ/X2snECmxKWkqvdW8PRiWcW67
NY50EpOOks9cyq6DqE9t9qM6Pz5Edcf2c43DUQ+tah1yal1ci1FO966TqdeVzzzq
OVsbWow3b0GMZw/Illjkk+G4yAB37lFcFdI1ztbcM+WEUKoc4OhsoQhxPp8YJqgQ
BKuEqkc/SWncN+RQWopqbnSpQCv3Uspw0Q1BCpJ+GNH24Psm56aWrHeQs7GcDAdK
qhBeOjSW24xWLZVesIuR/KnChlQYlkVNpCuaun8mBTmP3jJFxjAuHNaONSzHGjwC
jXgJRO/ezT3Ys9CC57MZD1ubdzoEZ/n9PTgOsTGLcPv6/UsuZPUSoKd9Mjss5oph
IwV12TRYo1SemEiOCtrGAIyzrjRY8wL7xSEwfGs8BVR0vZjwK/J6Ba8hpkMsG7ul
iRyfMNcGzvE2AKWobge9pRn+/MsJlelmXIWoQp8HI1cQ/38qDWjQrw2w9wkHC0MN
vBYGfJqxJYJsQrZadvLkcRwaZOv6ALFEagYWc98AxFfxmiFg1wNYaZEdcFwneljp
a9BlGMkd+KsZndXeKTxh0xCECyo3A5a4g1hInJdyxphjsJvqxQoFOlEvY2KuViyg
gDJ2aIO2ZqSTQlyf1KR/O8/95iNM/4pLaOWIiZOZfOXSzZsfRaPcgfp+tmB/lrVj
m/Vu/Vjadj8OvleLtgw9QIySwu3mUuUKpnkOlG583sRAeuCfBOtqvR/zmHjQ6xQf
Qiw1dxUiCrERLy4qIH96/3NA2nSR8rn+z55laEoHaZ+KPOVoVRI6Ep7IknVzbU6e
eYYuARZF4AfrfkzkW1AFnRho8yAIAKQ2+PO1/ZoWL12IKYhkmen1v+23oRHO8nSm
LjnPywRDk/wwGwiRnj0GZt4BUoS5xqFxLH4iTU46Ib53zi2RGCIQl+m3iv5qsVDs
erzvWBZmwVcVNeutzj4bYisZO+0p+iFW+KIoYSualsjsLACWnmh/PJhHEDTUXyY+
WXR8I/pTGDzIJ7nOd0Rn5zkWnfnFvARPcPDUe+DsFNHmpsim8RgOLd+j74FrwWDr
8RFtZ80FypgaNODMsfa76BwxF09h13sOcmZuNpzrrfsEsVUtlwWT3vfO/jJiwcGO
8bOQEabUelrijNjXIEW3WJg1GxCMJmNmea22ZPEPic3YhQ1jQ8aas7SpKyldF+ai
MxsvfOHSaDmrSaudyITPxiboaAA4KG1ZMHhRhyZilzuEHpRUIokx+GSTbHAxXunv
2mhJtwa65tL77lCCkwZONQKpNqrr8AoGvKtuYpaS+4YD+AiLTTqNHGmjPwbl96/s
0T8/odq4jo53hb3uomE+Wj7jv+h6pFnJLuYkrB3vDhenKulEkkdLwI8t7VKw2ZGD
p8RXTZHeeBCK7JyjhJG7XR6O6XK12QaeVMbphhuXHAh8s6kZCuCD2cBf98th0o/Z
7YI73Tnh6lh/HwQDQ5Li+IomXqr1SuOr7vcXCTZN78RBJRLRnI/FA0Y9pt8vNAA4
acREB1iPPF0ar71kFdk1b1MuZFPtThcihi3lEqWYjNUnEYoje89NGnK+n9jLTTk6
fgQHKVCEKG7uDKKKb0ePnYbisf5XtYATDRH67kVot/vcFewaDZW6/3YGAMIwDZic
ZOKRRUNw70uSGeaOiqNHasoqGcxYYxm30fYtP1IR6iZX7X1pTUF6KQ7cWiVcirn7
FxsLg2YFOHxfXK58LkzulohRw5+nbTl7DGR0Pg+uR31JSKWyagebXuiyqtVLFnjL
yQWw11dG2kqTybBbw5rWBdbqf+9exoLWv/wm9zW27kcOTILB+CDA5S58bAu5BvMb
8p14UgzjvEPyekq50BY1zAiug7ZuZXgPR4n8QLjPu9OHfajsW5oyYvS8FEugS9H+
IU8oeH9KaOaN3g24OD47QFzoJOCTDD3zPhBUk7TgEsEFnjNiaZ0Cp0QmB2y0AdgQ
nRw72p2Gx0n7+eV43sPYqISpBKcAOmWTCAyYBf8fnH2ByaMtz1uQkhThF+83knE/
1w1B8oifxK9ip5+tbhFQUgHo0o3yLmK3rq4nFHY39rgzD3XxfpXjbVw5vVX433L8
AxvaDNNkCftOrm741AINAhtsJYd18fKk4l5nhK7xzhVF/LyLspbTcHT6BmkAvTT6
AI8gb4JZidruH1kPsdXdtcN9uEvhSG4BLwQvufsHN9E2xO7lRxkJKrysh33lZKbF
ouL7tSwM0jZVZMcPX8ZNjVrwCE7gZn8Azl7Bq/WNP7D7b+gcFFCq7H8hzHtdPdi+
YjDspRbgHJ3VcRemjSqGIY6Lpay5JjuaFeGjhhm8Bwupf0FfqXNrHrBzRcR8J7Mq
W46kGJ/eiQgKqn8qv8WsIPbIVjdnl/VPu+Zu6G8EguqRthwGg2kBK1kupT9M/e1m
YYv3khDYiJNYYTE9cno3zBoPYY8Rot2Dms9GTya0T8EThviywFFP29teIEeWhJIW
N3h1swTKB5EBr5mWsP1xwLGl/XbnIlIu19dvdiSUBu1BABQ5LSkYZQp9HpRmH+E4
uTkZy8LpEjj4tYUklKkYkIzHz8Vda5dkLEZcJGz0YU189m7q50n+/Ac35KZ35aDN
xMgatkGMunljDekGYI0XmJVzxNVUZLpqjdeMWYOLZWH7yY47it5BkGG/+ZFQIhIc
H+8VCk7gML2mGQLwyAWhFKCETQCpXx7I23n0u/GpEycS92UvJAw9eK7a+fKbARXr
b5URMTuhAKW1GrH/EdFAPhN8zxmJvYIaA31p6MITMvDiHooGopNHYAlTfO5XR8hz
WgZ4DBHKr0phjf5HjXIn1EqagV+lAs1pWnHPjR1TNzKA6IAeJ1K/6SnzbsPV8VPJ
2iahDbD19+0GbZVjJJZt1zgd4ZnZZ1mDwUsGZnKETg1PfuRJtJxFA47MgYe/caVl
kR+rYw1fKZmQ6rdq5h7ZjlGV7DAE3WhXde0ANxTT8dzGSU7OMTIUscBj7+z2kbLb
NOt0imy6GDYl9k8Fx8rZ9xCAWmzjbE8xLHBQ3fkdtXzMhhdMk7QNEgZmsk2Juiyy
MYk72U/KuE1QhPa6+960RS+lFUgdhZrbhX/EMPukWTHtEvkFFD+rysHred0TAHNd
Qs/UrHWXn0ZkWglea8Aqp7hI90P0MOQIHD0E26GX06oRJ7voRDNYTRmiSC94iu1c
Qg8KJkcHodJYcbxJJLzdlHf3mp8PyOkgwr3OlkanlBxNx+nJ0eaYsKB0LbjggLQ+
L+EXKM+rXBBPx3T7lZU7/XGPcUxNJPW+KFdiCVpnG+UmCEN+IXROCDCfy6tHhc/n
Sgkdolk1Qq638bEpZLL8mEtNuSTjbFl/uchC/4a2oOXFHGhgaxyr+ypgXNKblDV6
zStNgw2fmvXQm8W+Mafu+BqxBFsws28SDYPyE7srp4kLB0gsj5/IZTbSnR7ZQ2Vf
CJJTtidzy5XBiJ1dhHy6mml5RKF93fDJRfAadZciUzGayohdORF1qnBZq5IabfSj
rm3CI8Q80J92koVXC8oOpieNZB+qv2jMwweb8FQ5ATSLCG9s38GM5FDCMrUcFbC7
gFDyFbFD3dtIXo/O4ByfbsNkz+o8Twu6o2y5mJCMSZEob+10rfkwmA9NY+gPjI1x
VLsHuNOWhuJ4hCK0rVqlU2N1vS6D+1ZImOSwF0tCRmKSMiZMWLQACEfGCZ6GNx+F
l5OXqtRng10IEDtnpWKqXGswf5dXoYsAvZvRGd5qJ+CqdHUJ0P0bBdBAuXnPGpsk
fKtW98/E9Bmgtgo8etMK1ZYMU1LV9u3kq2xOgULBRAi6ixN92JM51LNGy3Lf8B7/
sbx4wtPqdCFJFjHGNZFkdWYxMrtO7VCpIk44Ni5DGJo+SoT/UY/NgRpc22rw8Rxk
squ0C+lhP9h/5i4gx1RPzMlbufYJsfvuh4hIf3VeGHK3byd65HpPWJSu2fANZ/m/
vgnQP/+QTJT1jrPkQ+2ct6NjIkYdRA7lKfUWTIiHY57QRWrJqImBihcmeViarrDq
UTp9VUCivCitaQ/mgzSZkA5WA5O93tWsLzPkCYF1cUAOHnauSLAlRT9UT69hla1+
prkK/5kob6l/nY7Xk6V7207JjOs2FrDMA01Ff3Evyszz+ZpVPkYICSbcbCqBzMXU
eY0RYVvsEz6r5zzY64sgOtqrG4soo1tsmtldXuV2cYD3K4HSYlW+9WskUh7AL5Fs
KVtNpwretHcWNnpSGWSa3MftKV7cE/qxperNgian0L1U5G1Ur0peD/dO8A1uSxj6
CTO5qu01TYwYLP/QDHpP1BdUAaepCm/1T6bh7q1n6NEr14LhQ1XE+U48MybmjMm/
Tf7WAhcesCUr1Rw6zz6oboDdgr2tUwBqtzuu4uiso7trJS2E+IxUwOFtLWc9cBlN
XbrY5OZDSlBejDBTuP1T/r5qeYGXMVu25jeo9FyG9oWvxS+9pR9mqKQrE7l+cQRQ
QzO22mc9Sp8TTzngCmyT7+pluj2f22bJVST5sXsrQi1f5qHWieZRgnLKVuXkv0of
WiFcHKUKl+hRP3EFV2GXSghlR6w0VIzdHsuyLSST6r63GGZuUor2ipEb2teBXtpv
5PbOTap3Ayh/5AeHh+VxtXI5c9qdWemZhx2Mv1dNELuDKwDuZGlzHwQ1tMe+GIJK
ic7vqlaIvRf05TYYwmSmXDpGu/JXXQYYiuhYpncY8ln/Sf5bKt3l8U6oVD2foj2j
WHyABF13d1gqQzKo+9t/4e/H1n1337LdcIRCPYm7pfXqJNPtuGScS8q6OPcUMpcJ
BJ8pdFTYdQ2qQAG+oKJd34Jny5S+4H/O7tUNKd0jFdoMZxER+YGzyPXh9kov9H/a
1h2zOI0iyWTv8dIl0cy9XcGGgWIxXhARo99i0qaxcvA0opfl6hEIzTWRcjZYH+GS
uicFxM+1BBlcKfcdytsjy7R8csOEhqlf/WOr6VKRYnhI6BaDWzDlzCLsfank2BND
EeniforEPI3h0cyN/y2xH2fqxbj5u1dPU9JCtZgr6yHiyj+ksf8k7aKqU4Yacz4I
ATYj7/dMUDPvIGYep/drMk/BGZ8THVXum6n1C1tcsVzC0eQ0tTRcXx3//ne71F2d
jL47nA/qBXrHyL0I1we9liog2n9LpPP8WxqQfSivOkM8+n2P+m3MXHrsH+XWizw7
iWxLGqLy9AqLT6yUqAnPZhSa5aletavlYgQES3J7ubbBQEV/pbibXhyMxcaZUbt2
XUZzuZwPvqft+hDkjrsWsvxmYrXkk7JX007t6AqqJigSLbr/oSqS8zFGeDTKt7QD
i3T+mYVD+Kso84KFiN1VXettID0zd6tSAtRnoWd4UDBmGcfErzQbVTiffvbpv841
N9/ytbIRQzd2EFZc+JqElbqxG0ZMnqu/1SpedbmB9bV21OsLO7JiB26KuwqyD3gP
OIbLPai501BuObQPxR9pUcj67hCNWEO2aFxzxp/XbCGE5iWO3jt12tI+/LEGRiUC
veDyBNqg2rbOuk6Nnv92APVT0pM1tqGV0zUEZYjPWcSH5ZqCXoixT1R7mcSYwcSe
5mFYy2L6tyKxxn1xfjJ5sHLn/iJjCM6qp8rXitiMoiQQ8BtqvOvjRNo40Z+db/at
q6zJxRHYvBzE8mzQBHjxJdIpbCtD6B+r77GZSPi/W667hMf5YYP4d55L2DYMP8Lf
07dBXvI7fX4VuLNJIeMuaU6XKiGkabv91/9IWv/VjEo6V/xrOpoYjSny+GnvKSZY
fWSYs6EGhsaDX8tAygj3QgJKwDkEi8DjZLglWDLI/sZ3wjiyKYVdjo3FFwupHr8C
V6m7EsgxhDofasAZa6P9tXmNHa5jdG8LGHPMDxs1oJynfvACc93OISsor46kpK+7
OYcUeI2PY10VQyKuIFnIYCHJcr3IlLoU6yxn13v5YynjgqStWwuHCvaxZnIFm+U4
6Yao2jAYGEUn/+bT/jSiEp1oZKY97oA0nSSYj/4QjKrpsfDdMwCBtO/wQGmxc51u
BMuMAwwfOAKSkBkYmjZ6upoLorz1mFltvFumQmQewTsKsMW2BRgKZGtxYBIU6aCJ
e1thfjYEkIEuNHl3WsvnHmiF8zXA0ek61xKoawukd05Icm72sk+QPgViH/JOLLez
7bEIZDObAE1j2V1xKp7ClD57ZvOGfbEgRt0rkFaHvCE/s3QlYPSnzZ6CYNhHVjpu
ZiUzhIsTuRuhlpgKF73EQPWBTHTj1saw4EJem4AukZ9y1U0qdJ+i8uI3q+GBx59w
H7SAruK4Wid0uPdUjsHiw9NIDGcTzAVUtv1fqA3M946eQEc4NAyNTFGuDoKgEZqD
KKDHga+C746ufWrt3uVCgg/3qQb7TUNxgMFoKwcPRME6vzYmZK0FkDrI1p+TcBY4
3xKFM8h971pjQu8Uj579C/GttvF2gjLyg2VeURSQIo06BWuRUR4FR3CPr5FPPfcS
12ehgdV0ilc83+EOJNN4XgmIyslscjN+C5vAbPvz0F6n1UGyqZH1yHumPNScqUuz
/FW6WDwT4bR2+E0/Swglx6Vpqr4bVskP9QKFm2+IVetA51M3uAX/jZ2rteVlTRIG
MbugEB7NPcwP4IcGujmjnGjSuJdcXlufo8En88ZIgbN27RZw3KeJpjCyNCAwYLTS
gWVNWxKqSmrPqVK5JbkGt8GcUOiwfa+eref3Q+g/1V6cXJbpX1LGUhhEeuBSVN8/
Mb5sF7l1yc3cM1pgJPhf1EJ2SvEFJexKh0ySRlo5lY8gdSaZ1K+Snscv2f4FzJmb
oJBIc0GdI+cm+JgmloKa54Vs7oJOlWVDwAMiIleWoD9UVUkq3tYhd+YJq8Vb3cVU
zZctdDT6qFJuEINUF4fWFATXoH6/17SrwZM9nyJxqMEgFbsSFM04ogO7YuZ4I0Xg
WVVHRfoRNarcDd2U2Kz0BGy8UOEJd8/YjepgvTgVMnhhRoByiODPSwS8pL70Drsy
kaSOBS35JgoQ8BOQs3cfSmxrr98d9QmEF0L0GCvw68LQNvaANdASQ8uxjzKtBDjU
DaLyfu5BBRLxNoouQiOEWBAKspZ7i4boHQbR+feJGdOiW9yvPV2iWNLhELV0T8o1
CX7IaMEsEFjDBeGAwS5XYm82dX8/1IXBldQG2rNq4cOFWlleG52WH91wguBssn/F
uXedtjbBXb1k1y+TqL/Y6O/4boZ2YY36X1HYx8PNNlajVTrvq5jSgdePIK0cuQ6k
OuuezLxn916ZME9VM9v+QD1geEWhlzz6Tdaw5TuEthfA9nDskjptPAqpSkhx/H7B
eVv8N9ukiNKkH9+A0ySGEtUW4tlXT6fWutNmPKV0nBu5aymwZYInoGJkqzLg9sO6
3717HLuWv4q/2UhttqKO7qp8iAVdXVdXVoCuakSwBzLu/Q51WB41uEio3uVSIsmF
4c9f0Mj8q2fgRLcsuYBPvNKWErkkMzaeR+YukEn5Aa0vQvZWuK2tCREmrH8lb6Jq
sqrS0IL2FNITWraHSC8imjGPa3HokwvBNoFSCabrr1zpndIrEeF8Rfvrp01FYdD4
nf0yYuRwXNGcvV3U2BHNPahoTuSZhgSH6n7l8z3dmwPOY1bmjMgd8XEp8bR7kfl5
k79rcd0+KhknakqmHthsFKeuUJqyFhiFj8EtJsFbtv0cCYkIrIodi+oTZMVZ2pR7
MferI1Wr8tMZSUaAHlpX0v0M8KPw5eV7AFXf0YUq8M1I8YA1HmPOE+9oedaTN9mT
HSS9Ebg7YIa9kMqtV3baHKYut1rxqeY+LuAq+cXlu+7Evn8FsJxqCyUpXPz+hlX2
C64Nerdlt9t2qhtO4GU+HrYf3IksL8Ccn6chAwH+/E7MnRG2dtQ1cxbIajux66Wp
tUmlwUA8XLNhi2XQhygx3qIFd17RNjdqiHOd6sxQxx/CdIUpQSTbeuATzXsbEnMC
bFw+gGaTkCyn1BblurrtH/30YNf1sjAApuofg3zwO2OPQCWGwZZ6ocosLsuC0QKG
YGda3AkB0iVAcEYkQt4c6P7kHwuhSdNySal4J/zKngIutpk62nQGZWzmhlYRWuVt
KPS5uK1jlMbA8ngVRJ4seAvSTGqb7W0kOZOxGgPE9TM0bldmajxjen5ZxN2Hs5ox
1IaysZxipSDpkh0gMX31KHjVGYM7qeseAhcDzn67tPijFsev5SyARtfv7qU1+1B8
wp/vq8XYBCIl5RvNNvhR9sCXR4TzPMTD/3fJI45PJ1F8yXDAkyNuiqVFZyzV+TbI
+Z3VYJmojUp9Y+jrLrpKIdSVDpnrYFVmtUJ/u5XFmSq5zlo+CanfEPMdxR5OkiUg
cZC7Oc4L1hPEIaNF8FzuXks7TOAqsdM6XH028MAUqZgFVHG4cXv5NgN5v7gVt4bJ
AjGuW72kXcnMuDHvLreCNTDgv2EUnZ/qGk0RagrBpLRt5cxtjCQkyt541s+sjFnE
FfuL62c7n6ScZAvRQnKJ3kiUAzZRxOUjikCdDZm6XsLTcmIjXk4FyVIyPS52m0y6
nInoS83b5DRvYXxTjH69xSMj4JAOMaIlk7Sx7JmV9+uYZgX+i6y4pPqJGboDakPV
KDa2V7xeUzlrhudNXUzudZ1HIFlh5uHkawBVOgvIi39JZDZ2JIa/rMzdspaJdn8J
PygZZkHLXBsJiity/SLxpf05+iPgDoCMEAdrMzKa7vn95j+Dl0qqdTaK6AfIMS59
2ZicVmh6OwUxPKF2Bujgbjb1FANdEHRR4+Puax6TNrpUEB78zN8CwFqsoBD2sxV5
/HK65Q7iySKXFWfWUeKft8kfVha8fvMhFOSxhn2+Nr1WlgKUJXo7bJlEAgzlmzHn
1M6oM7ko5D1WAFVG1RmQgDSMYvWWY/lFwTbJe94W8latb73lXLBDOyzBPN40eFxU
bugVDlm3bTAQ5uEO17SQP+Oo6Co96B+t9amJrqSkohnfRKITT3RTq8287/+qOBSM
guvRBiRf4RVSpF3vQpmTI3sme7iw9jbApp/Ds5nLtqlT7pALXmefBqmZilhdHNO8
qd0LKzB4jU/pJkJzEebhputVhEB6+CVQgURRQHITLH7nLOqaVNzd/BXR9EUfskQG
4D2bO2CUvd0PE8y/pvy5v/64yRa7deq54D0OxMxYtK839eFp7UbrCvsKkWROzcBM
U9LGkv+XxgWM/9LAPeSTst0kgsao8tpAXlj0kHOInV1mOi7OHe/TRhT5IqT309xH
1N4a+CKmeS4z3j4Uow2N9w9w8iHJYOhvKFRRJv3eQ8s7E8nFezk9+X8/ftqqAZ7Y
3lMCo4KPdmGD5NsIY67mrigGD4Nlreyx7psardSMUc4Op2T1yqDPepgiLJBESlT9
GRn/SnP2vhXnk+1Q9bg1bkwaG+X5hqzEL74d9i5ene5hyEPMHn8B7++lIqQIrjJN
MNCb3dAqjR0ml8AUNO2gYiN1xGiMlR3xd/tQkKxSKmqdJnyql9edqe8xLjZLDjRA
QycNW+mcOFhYhyD1DxTgM+JHiMtWU0FXtCW5xajGggFzGpYlhFzkfSIq5brAUbLZ
1V3V/vNIo5a1QBQAz6aITThOEYbNcmncerqzSlqrDm6lBHs+Qf1Ux0Is2+afMcta
Llp0I4eucaZbQuF8UuBwZCONzE28KUZA/pBKubvDOQEISxhv68GjjS0Za/Lzfv18
ou7f7lkM2plyTuHiklOybj5rheSKGzNagoOS2FejiUj+H08/l2lV3wDwrCiDTJIj
EaQcjXwF+Giyb+XRuw/C/50KkwXeKv0cn1X3Q+6RmPzpoXsPXeO8gbC8EJ1dfnH1
fo6dEH6AtMO/wfcpc2UskyrI01rZUftrIM4RnTKNPXCDqNYZQBHyNUVRMUN9OV95
gZdkQ6zdtKei7Kg22Rw5x1RRjPCIOi9y2fHu2ZrYJgJuOMTAoHtm1w5LSsexu1im
lM9qYMMlwUHm0BiLpPSLWkaQuUvhBgtT+1lKMYTnog59ZFD8tBbX6CAVbNUth7GH
I1RO+/VeFrirfxxBwwrTNwTzLzvlKHRnjrX4pAH1Co8dTZf28895lqpXglJKMQDX
chwEOB+FoxOzX/X6Fahj3Z/vb4VqJopxu0rvolwOGy5Tdpjj2RF97nmAoq2K/2dU
lTqOEMZRuDW4gAaWJCW4A3CNPwU5iQBvNwU8eSR3PqkI6hNHD8VJM9Q+xoXxTlOf
8ZZ383aAAJknh+zXFTWDPFKTTWp4qovbR+Lp3btXuk9P9+5axLpxIaWKRc7PLcSu
G7l5+WpPNetAYvfByuajvsY01IR1IVLfzMskJbzfJL5pSlTOSwOBOVkXiSR91467
WWSmjh/2MimT0Fcl22tU+D8ORjUYKAP5HDQxiBUSWtwj+xmp9kXwPe/asIa9bKoO
SnrOtHRwdg8jAdRHfuvvvYL8gJt1Run8WblnT8+tSVknrtbPIitUrPTTI/6nHarf
BYa85UwJiKNcPKloOn8LLKD5v7abPbqCNC3S5YBvY9CB1Pcl982y1qCg1SwsCIkU
dC7ZwCvXAdBgWE8YWUO0Vqjgls6WsEb106bCqDLCtUFE/vCLuF071wXbAfjdkokh
I4KHdhVZUehPkjVC1EGiQQf+zHmE0SMuXNJUJaEAjB3LstVqsINbHxU4LziXANRD
ZDebx4D/G4TKSXMzll5BGuLDzW3JIrGz6rihAgxJqc5kQMHwVFf6OIKGjkNOvEIK
Iicls2LtJmoUVYgJ5/qqLb78HbG0dYWz54KGm7Eh/Q6fI4zqM1qWYnndZ4swD49H
xKFhI2J8AAPFVuP6LFwXFQg63DOD82mvxW3r8L7GiyfWbzgkujr3fU9wnvUunzSQ
ofFCmqUfBp9gCL3yzz5mUvzXxh6o6TJJJEFPc7l7Jr5M20MCzYCNw15rZLlfryDO
wTvmsXd+fAPdIT0C+46y+oST4q4mH0Ti6U2st9JuTZ15PwWnvhnUbvX33wZzV+FQ
V2Lg3CNsQ4w0OtMM5qSLcHZl61zZrmCjAJE2WF3trDaYAHVB9Xieb+C+gdRkrNdx
C6fQ4eImf/whMPKwZM/SMN1QBkCdbBc0pn5iOt5+25Wks0wUKLsdCCHptsFQykLz
P4Xb/9oe05W79KEtus1rrawyLOi4nPAgY/PocoRcYO2yz0C3EFgWw83sahsuakRn
XtJeVXGlwTjnNwuYPpEy+JaPp740aajTq8HF3xy/Ueu0L3MDjrdXso/cY2FQ4Knx
OPH1yG3lJhykWF97nlnWXHF28RhGe1shiUAQFU6ZSiMbs0c8JuS0kOdbUk6Jfpkh
kVdD4Anple8AKQZY9w85R6I/wuJrfucBnx5HTR9oxQ+4a2tfKyGjfVJ+5SuNyd/o
qFfMDlmAlL0UiU06RkeK8zm6q21CyLIao4dPf4PE8TmlARTfI6sZ0YN+TqVqjFB3
IeSi9pW/HreYZHLkeU1DGjLXy8ojF20x5qH0xnpSwuPLJbsAeWLGEIH+uzlxrRmO
El4bE6TqIDn0sc681a0QWeKIPmVfNWdk9n6dG6mrSeukjsf1E3wjaxY8oEpQ1KMy
YAhGCzgZIc2oZxB7bqR06nBDssesXeqFs6q7pHp+BEaQdwt8Okeo1YA1OYWTLVGX
m0ut7Rt/ucOexT5MUmsTWSeurLclecfxzkQcqys2KrYNSlYBQVcwIZUsD5HO1fYa
fd9XQpBk+duJfjff0pQdJrd4gPf7bIy/abd70uc7oL9ZWJoko1hb2s1ob66AI/5N
s5hL+2sAnYh+E/PmOoU/JStwDOFeKqeWQ2xUnsge1Cg+TV4bPnz6rDMabEvFMGmp
nfdQX4VcZ27FgqXmNfYoPFQyu3LvrH/PYF3Jari+1g7GKGu4aVpmT2P+eaLGkXL0
1+lWZJ24UCaS3KOjwvGH8iDowtg9/+8ngW1IZKUDQvZCbZoQrqRbiUbvCM1Ixvvd
QCKMSMrMwQTCmQYIgOD4qK1FnwE+0IpEcZwJv96fmdm/et+wZPCJMnQgwFPVaSMW
GdD+Pfz5p8liudejEcsO2eLv+WgAG9ALqe3HnPog96XTFwA2Z6A5ejsQQb2Iz/8J
ewTe5sz/PAoi1YrS4h8ISQ5JhXwxT2I9jsKV6vRGDS0I1x6i+U8BJ7dQS1ydFZ7e
VyszFqII5WXOnyNDQ656XlE8lDvV/Yhg6n0Zej8/Ux6uBqLeD5E+1mfrs2DdZed9
wptBC4kS0GQL+O8OAK/pylSXvdTVE1PhrzpcIkCpJ5NQnoTL1muJ6HitI020oJZo
LurwjaTArTMdmQw3QR2bDdWMPJ0nPDGqYvNLnlH1D0XOugVC/hHtxg0WtAZ89lf+
1vgaVMOq7ZGeFePdIH4mtsmhsn8jQk1bAogAUrfsD8ixceHvydl10RjKkk28ErGB
M7VN7CoMRgPfhf9hXfnUZxPpVt/r+kTWnevr1+D1Rpk5imjTEH3tVoOxUjJVRWF9
KyDAVbfjXQNUK/zSAqaFWBLv9v+6Dbhy30Q6J0TSGIXltafkoAyFf1LHDQQyJf7O
kSZkAY/mFmWxkK7Q072/Xi+K/F+QE0Uq9BQtaE5VxBLkHRqnkHZBSikz3cbFiXJf
4Pku3gw/us93JSusXUvc2J11c+CusJqmmEoejrQAIqp0HX+fHcBBDdB0VrbJcRNl
Vgdb3soo9R9HOPfFet/Jh2jhc1GhbOyfzN4MF0ZwcKqI3V0Lt/p71hNcvaiwkYoC
pkfs/WBieaNERJW6UPFUKdUdKtZgMHV3NIZFe63zukVasfSY8ubGStTqml5exoH4
OTeefHLlKRl0AY/Dc/TEUgZU40ZhJKBufZwSQwWzEMbH6jWSLEWmB4WapDkDeQqQ
y4uYAUOYQ0AOCu7mFQvJHf42g6ll8dtnGRp5SH8/dmDAjQ2X2dyJx5lNZFRS5OSC
djNMBGwijX6yUz/lmac/djb/QPJmsc0jgxSqusnR4HsKgOuJ3QXu3KT6bI5EIsoS
0bg1TI6KpNDYnypjm6HzTOxmwNuWSmHaGRIbmrIslQuEwVVTJyNDZp3MZMYDJNZc
kxryNYnL2yClygkDL15PsLQoEOiGjj6YlBbVQxz0awX0+RGDf2nrHJUOqb5CJd96
Y/nNtJVLF9+qn+ZW4CbD+GIkkJpeanjdMaDsx4bjFh9KGG6pgfYwJX8/55lS3zAs
hYYYoVuwZqSh50iVmYR2kKSeiBfHuontEZB/aEA4uXkYC/4rcGfHPFv+MnHmPmga
7pnrPZaLukx7BMGBr2ZGV7nNsw6Mcw9QLqHH+VLXe0JsIIK0KvhRHLzsGg7f7LQ/
81BiHHy8uOAp7mbo9+zeIY15Ut6GiINzbMFvaAZITf5fCX6uQxWV9H19gw1GY7UV
/2nsup8vAKdMx0+KJM5jdnvclrVoDw6fooDywkBP/2Xw7cyzRtx8taY1AtGKdfdn
4pkJif7xnEAcSF7XZg5vsgaBjiEqB9+mlAx4VARvqONTnWRR3ynCoqgA5nlmsn0v
Yvn+xfajfoe3TJLcrLTSthuq5Kf7GR9F5eRo5YH+B+5EGtQ7tWGQR9qVaHBK6IfM
ZKjVZZFeRocQCXfxnB4cHjx5J6U442OOjdd+lmEyPxQ4zbWLSKpLoewpIPCpVIF5
GjCB4KFvSksKfJS3vOiQGhnyb+xp1GJl886H78xZJKY7UMefNTrdS7yGcI1SZe/T
741rYSQV1KhvBbqxaD0Uagb4FY1xbwUxkcBiG6Q8/m13hwOAMwKJBUsA9BDmFXRi
xp1GplzPXQRrdNJ/HJ9mokDh5HL2PeDmOJnLzgyTEXEkEz6FSIYZMDS5bFWLg65a
4roQvz2Bh4fGrWab76Am+WCVBZKk+ind8d+auCME4+8rjv4Jhuz9AI04ZGdUdw90
AWFVOI76oFoBBPX+61B13wh5AXa3NEujVFRN2s/hkgm05iOA14btk9263pD5IgT/
hHTlFP09i5vTyPqzDufslEA9mHOgXVruV7XBByptRE+uB6SDjFoXM8P3mskN4JVC
rMbC15TkoKO3mvEMf8mgRFlZzy5grOLn/E+sqzRMPvMac7/9kozutQRg6T2MSz47
8USYXlZ4PQSRbPWcE8fLiWXGyZ+3prS8htRSQcYwQ1T21Dun1DjgmKDroNo6IP5l
ne/cp9MmWSx4R0lXHjg6H3YXLW5fyMAu1B1AnVif3ROMBfE+6PzqPZhpZY1e9m/V
yKje8nLYPjRwlMsNXGgV9a203X6Wy3b54bZYNys84jUPBTMPJOkybZEf70nR5Req
SnpKXaLMhcgoDMUugqtmzGSUXKGaIK9ClEGf8H6f0x9idvLfwSHe53V5lz0/NlBx
0WeZbXeALsA3jqxkz1hbxQxvPeDV/MnVBqyPqhjos+3DnMDSZyFoEGdJuUzTS/tZ
Vq+Hd36NGf+qDtlc1j9MfQNjd2OcF3DawwCFSvd3/6NFmYkTWKJl31bnq8BSdPLA
/5J1+8wnZBn553FQdQweQ3Y7dzawJaRZ0oejpdaeJ6BiAAEmkWWSlISdWjcmgtWJ
zEqM8RCpXDVaIgQW2ZZvDctfMIxtzeiZsNenz1dMTGywbkBbOfjFWMjfjOFi/o5v
ERRs8fZiDQoMNxQOouInbVXmnkt3zEV4HiprwVUTgspmvO7LZFcJtLzcba4IgEFW
fS0+BK2J9miXM34DB02HZrZdR6C2se4Cuf+HmYhnqkVDi+3LVAuM9MB64mu53AMb
Eb8jT+VN5LCLsg1s712EJnT+BrNudU2YsCt4n9ll/FHDSMIQVavwBitpM6ji3RCA
6U7uwMwADRUrpqNH+vK0eGraD2/fh4hSaqN7uWpoik3CLTuJVjoPJfWBG3sUP2s/
tfj1NzHE59qNGtag3CnJz6AMZYJVMY/z1ECf/DucTuGtTKLV/z3Q1db40YloqrU+
fR+MBL4OEukF1B14BX3BAP2QiTK1BHYHHK0z1LMMGAx7cMcgQ88sA5hxS2f6RKDI
NNEzeHDOr50n0S+9FsJA/CZovvcjp974b5BKJp8NE+5EWLtUAF9DZNJsqpaMhvhe
5j90/P6KojRpCOuCRRlpD+Ty+Gs+l4r1pVD0Ybu7SO7Mqr5jfuZZ9or0y+RyEmwR
P7yoi9eVTj1YVBn2fkMd0rU4fVGntg7vUIG3QjFr34q8/ImGKisMZZy5if49ELj1
5O1qXeB6haTD2NNFYk6cGzScDQP6EEOZN4f2sHGJQ/pjibkbIU7cPhtHEcBqGO9l
YB6vYI3oHOcEMqcTRE0spNC4vXbjoLQRwIyDOHkgAqCFlP/aKYkMFC90QqHwj7tc
vxhTvvfCfUOhai34idjGL2auivUz/c6aSP8laqQ9kPN1FBzRP8iqaN+o/M3R/xl2
TVepnPoQobJ2PfbxV5c1GOtGIxvUXQqEIhT5Rfr5+lS42nTVRYAKYfA4stuf0FH3
jul9jndvz4A2nsoExWQ5aJzRUnzWn/Hh7jeQ5v5tIShZfmHR/a2TYtxJ6Lx9oYQy
+R/dhIuR7Mu2ZEUo9ThE9qakwdDVnPh3AXKd/a6ym8LBIAbrN7B+KnVlnyIiqhv6
iMhyfyE4qqwbEDBRi0PxDEZjgA8GR2WFbH9bgTcRAl1gr3aMnH4YMOkeu1HaDI8O
Kae8noMGusf7d/22DlNh/AefBII9rodc96nf0KUchl6wNSWr0swHsdI7djlp7MJ0
fZxR+6g0EfgzwDjfKM4c6xnXfZJX7Q6WQhxAnxxdQw2aIr5qsKBdmx8ceG2wTmEC
1iYNoHQHYCzhvPeLuTCIG4AqCip4JToT9VlSmMEwt57DdKsBfALXxveb2SEe2EoZ
4NXowrSOLUe1hL9/tOU8L2Z25Nu7RYm8OpenxaXV1vmVD50urgZ//JUtxWkZe6SW
mKXlZeLJVPgl3pmBJVpu6S4dL9eElTUk+BiYLApNUAyF61vBQKa532K4++sIE96k
jrG/BH+F+uPC/LbN1AtCpMuwcMIl2dhXGHmOIyWMuNVHS6gJFOc5XNtRm94Q4SB/
azuexehMuQoRTiyYhg1Kh/Lz8p9088COXrSw9Dby7stSSMSWX+QL99YIMDTCMCo8
Hm3O1P3B/C3wit4ilcW+zMcs/A8Ee9oH1fBsbD5pU6S3gGdfyf85Tvs+LcKGiKcd
Zce2iOT7Sj4082NApLFYAEtekMXux7aSMGz3bNhKzd0JxTVqz3258ZQrM7V+Qw4o
CfE5Jzq823Ct+s8ZIBvuPJP4wKPyz887SUGe8QEBHXMKMvwfGdgZj8wbRlnwqnnp
2l1jFuvSYbNBPjRTv83oFrh/YzOchY3nlqPr+Yo0DMLVkKfJjoXYqZHOQssxBs/x
TMPY4nLnJHkMZrTHYbJlqmtH0MWFTGHoDSK2HMD4cyJNbE8l2ca2omllrLyILC0X
xIs3qLXP9cjdxKOGjrKTPD4/UWvnmeziB/oymijFc1tqNN7hzD05kn+//Gbq2Jxi
8jcGVeV36d09BrZfpUEddlX2nhTqYMAIUuGlivcYUB7nwwvdLU4sqyleHaRqLl0d
YayJIwXAH9gYDvSyU/20BUx2tpKCkL5ckADU6+pwV30Sq+iR60YDaMZWSc9pSjeL
x8fzFcciIFgnvmxT+ZeFOeuCFrYye/hjcNBUEZLxQytE8uoimmemBUbu0xSfD6mQ
lwut8x1T3Jzqmuq/rKpi7iDmQRT2/Vyn6zzivwWEvXlc1V1k+mDYWhl7rz7U2yM2
zGof/ASiNLBXRIDBLXtXgGuNaeKwi0xnRvzRscvGSzZ4/mHQYr1dybcyKrkAuV8F
ZzayY93+zIKmJEVm1ol+e0u8S2ipaAsDhlFmffEai2xlXBJBP6VuExVZzkLCZRwZ
BI5YnASsg/GCs3djCyGqe42BnHvcPsrWa+BPPRy/RYzoMZNZBFdMfMo7Psfm1Jfj
tR0Z5hbceH4irJyhs7KWe4/5GOwEBqApCfGptoUZKaIbgZtSpZ866Q9Gbb+vYPiE
lNdAU6GnHOTcqjOzlCWcXpAxp3fH4EFB8d6NUGYQ53HD7iFBuaOXzxKnEZSzeaWF
/jSkhihJeGwbTNdR+ujEFBgSkCA1DVnGrXkQusyrf8l2lHQu2Co0rgDb3QXs37nH
cIN06aKzTFW6rrUua3URQ1VRfxDn8FkC8ju06PoQI280V9OEKKk8U+r/StuQkt/5
h+ziuRYKrAEmVg8wvHocWb7OopScOjSviQ8OIDayfeydo+Ozpw7XeQl5hX4hpwbT
hYFLHVurVsbpn6QZ/oUeaP4fs/0XJMx+BqaYPEs8t0suNbEwZ4yMtoXQseDJFJyy
3krxeE9wpfhaTgW4+V8ag0dwoqY5kVncCIRxoiDwWSUhmaBAR2aIAuXCKRcvFzyJ
GVEUxSSGsMUsCY+WIdRlZ3GI/Ki5QpbcHAmKdTMuVAVtpSBIdNzfj5qYCxHrKtSl
PeufHUvWC33q8Cf1+mo/RGV1P8TjvRcpPao2oxRac/Uzm6cBbyfNA/eKzZJQou4L
9EhrG/oocluR/LyDI5KXCDEZWBL18ND45lp8qnU9fd1olxkmWvWHWUx16E0Pw1vP
L6fvlfNFKNtkMY8t721poSmO5nzApO4Tp0Nq9Ts62Z65el+41Z3q2ndQozA6kK7Y
B0wOrgy6w0mD2pe+hUFVG17J27qKXSgLP0KElDvdRxUrSigcrGqAMeGgJk5sxlS/
tXJnKcSBSYD8kDRtpzIN77bLnwLocvoQuj3JC4zk9LoqwXXatHbONFsaTYr45QM0
jlty8JK3huo0enlMUX6CUIH30Wug6Llv1POkFkBJIi6ehPkatPv1FgpQB54GLBIj
RsZzXeaVTVxuEX5J52x6AvVzmACzrDigLbbM6VjHrLvQ0qXvmoeA2fS5uIy4WmXp
cjQRVI6b6/IZP3r4PptejUR4Ao5bPQICO7m74pSTyUW8fLhri8gjF3X1G83gIPwr
Bi/8PntkY1U6lBTJi42a4u3VDRBqh1VyzAjcPyfobVYgg7lWXUZEV9q7m0JdQhjO
+XnNqkKnDvWJxQMeYpAXO7D0YHarBlSJiJeIf0ttYYp9BU9GTB0o3FwQn/jrVd03
HGu4Y5qWsYuYVUUpfLmazQTP2negIlKj7p85ZW1+q3CBiKvWe2L8AFTWTtU9MdSB
/dCk+Jkdkoua9K82wO1TJeEECF9jAIbEJxZPfjg/fnn/BBGy7eMxbw4OODE0XNhv
11J9/1z2oeOIeF/SLf+ANI5qRDwnEUjt+R6IH3uwGwYSxSgTU42aH0JqAiwvnbPB
cMpdmcH1MWXzKWc5MM7RH3W0Q4TQ2PwZ7931VdSC0cZVAqICL+xeVNo/ezl4mzmv
HD9Nsp7CPK1OxwuacS5u7CI816EMXnJooQImDQgjSG+DYh/1/XeRnvBHm0B4WrNk
9ev/Xthz5yLKOh9wh5CjjXoljmIa4ie+tz4QFPKzS+GF7p40gPtTHStn97ColK67
8WlZH2u8NOtkp80E955OnGz1mySAPPSn/FPPNJWNOS0SR7qENsLwh6pJxsFqu98s
l9P9ZmTJLlGMBK6ks1EBryIZFnxWQWqR4S52VJIbVKZueEPzY/9QYzrrrJo9fI3p
gr04xc3gxyuEU7Ow3zfCuQZ+bmNIdSLQiMLpyq3EX/0L2lSr4dFx/gqHoxUT1+Pe
iFyD+lTC/bfcTor7FKu+UcShWjS0ukUxdIDKmEtikdNWffzl9HGWZgxw8ubNR1TN
tg1CqnLwvuWsvoHhJthuL8nbkJS7pPnkUJdbaZMQzuktHf8hItZRQYM5IsMWpmOO
z4z0VuPKi6+sy01Dd4d/ot22xXSwQxR9bx/TJP/0Kwy42kPqBAbFANtnWLTX/pTi
+M5SySI/cTjk4LVLedWabIw7xJpzEvTJlmhhvaZrO/tT0q92sH9OKOnHB5oYCqDh
UuqIvZyMcZ4zMrbPEXO4XUy0q8UHNyxvs/ZqvuHmXD4Xk6OyTdxInAYHoz+8q8dL
EEDw0VwrmMyEEPy0Y5sU/MoeUr73GN6BWaADACugJ5ZfgktOjKx1YEZrM9hp6SfQ
ql9lhdnq9iCQDM862qI/0IeC5ByEgz8emG/JV2IJ9to57w0QF3X3+363jdV1LRds
rrezsrIHNz07GNvdM7qAC8PngVTOZ+leHfK6HOQJSQKRjhmT5xoK8CNazcttNxEC
9phmLy0fZ+uL17dJhx8/8FEDJPprF5fQnKKQVieTLuHV9gg767qBhOVnoofk07q/
u54kgEScOf5pmWsb4594/KxHXbGUANBU/AsGO1o9iZedwRgz7NQ86xctchQJAe0F
gynQJ109blJr1tlCOrbaIIwokzQiXGGg4E00iFmveYuSuCRd+Lk1PmOd3dTCGZsd
Jzo1NIgOV6DoOHmSz17hlf2BRuECLb7tPy2FaoFgIH5YgIWDk5/1bi3fSlMtdQqq
QfDx5QLlN1d4Gxu4HD7+DK8Yc9EpylNho5EIBiok9A/pznn87OxBNHmcMCQNlLQ6
CS5eq/I66/4GthB3cZKj+i0OHTfZ9rNBu5EiYnDu72BxfZsgOeuy47cbTupETKn9
Xx6syYrKayeDK9tBNGzSFMVMV7RoA5aoKOcu3W2S3YZo+xMOqrxjyhyras/q/RUn
RqmcnfB9V4jI4krP3jIJQizG79gBgLcwRbXZIP3FzDxOGTtTgyBzaLc8FB9VpfTw
7oMJLoL96kKvwMyA8/gOHrzKJ8Aaax3R1nQ+8TOeu1g6VFPjgeQxTypR8eZWglNc
Lra2MxHHkAHCwsrjAn33BwIcwRUpaGxsD9H9AslrZ8HbaOd8kL33GWY3lGEqhCck
G5/L9erCSlbHlAvgrsgGpfU82g0ykWFBkBcWzCHk1Zc02mq5mrqf2R1qQ4O4ntVY
jCFqct5HtTL5tLley/VwcTXjSpBGz485pII3/hgFHBGWkCcvNOrrOOzpk5ITvrDi
4oYodkTL7giprjPy5Sh2q+plJCUjwZbK7XnMyWJkrWcBz15N1lwGeNlhDG22BGJR
mnOC1HFvv7cDjX03dFSlOdx05NjFsppEbMba45Np4VK2DL9cs9Vy/FlCQO6kq6ZO
2gkbIr0EWfAjtwLyuWJeJJ82YZ00urgKobfnqAosEKW/PUW4zfE9FR391p+0wkWr
B+T+CcEH13s+ZNfgFlJ7ggAb2035eabPNU8iX8YNjHEl8fO5pI72kHGvkB6XJ8xl
49YPRyB4K6yo8+XHg9SkRvMphIkpOVLfSWgohEhxSXzRgfuH89kpuTDeGHeBbLUm
4AayAVUNQVoE8QNCDPSn4+ghJWEdPD097hADzxeFH9E3wRCrK+Bnj5rK75PXtS8A
wkPP891JYl6XJbzKkiRBCp3TB5hC9dujhzA7ql/jTUhHMpnIuAs9ImMooqNgoz2x
sMGmDEcIM5gwpYJ5Y05sSUdYM/JXi4ongKZjUxTrxJHLCy3NvulmHyhRLRldZjMa
28wucVQ2EWjmPbNrqjeno6xlHFRmh/NtI6saJNmPqYsHHEnOLjh0WdcBBNWmoKpj
gXecfElyKElxzSABnl2RmZHE4yZdd++ar6d3+CvTadc9M+MzQyO42FWUTarEBIHV
qq1laoKn7oZ/cNHYYj/Fyu/aPQ6i7dGgU24+amwZmj+FoP6vtNYiCsKjuu+XkyVW
kFvnDILmn3+RgrzrgyfLNa/DZQVSSnmdmjMv4KpSN/M++6U8s73bInp3mHJFvfzq
pFRoOarQNGKkIS94SkXIJYdMwmSkTM8YM5ODtT+Sa48VG8E4wq0pyESq6rtR92jh
BfkdMMIaSZX9LaDUr4HKsitW48CICZqbatpW8iFmhrKPy6LmHcoxIsHJ52Z/xcvR
RWIZPkiV4VcU1oxnVgDBkg66vLKLJ29qEpL2fgZBjPgzw5tA22KXYxht1he00BhN
5dH3cut6Ve/f2/s1HTr84JbEulcV2HCAJIVesFcpImzEneXPIReuXmTUSJTqJr6S
L0lRkeUTbq/U3oXJ5T/JEEa33bjp46P/iE6sh0Mb7UHGekhhhd7DCkGry8wTzgOj
h63GRU+SdmMWEb5L8TKI6M6imD+kxxFWpEdeQCaO/K+cT+TYLo4m5PPE1dl1ufmm
ZxmWUOQmDUYNr8sSd1h3zdmyqtP8Ls+IwLe29BeHsbx3qk8fbsKdLAJH/Fe3Um27
AvT5qx+TAqaI+2tDCR090RQWtbe3BfaQS2ZI3CdWmmqyGx9MG3Vw1Rr7r0CBSPnv
txAN73NVKPSsUWIkv6gOAGfKm0LLaTsobpDxSFq241sXTTST/C+AzFNQIwPuWZ3g
rn1BBYM66sL5Y7CaEGrVrQeFyyDrTga/EnA7VPqyroZBP7XNM4xJLwFBv/ZGvmi6
kFs984l/sHbx3ywf41fawKQ2X3RWsGQfNBXfk9GeUMBcVYFHmXWIWD3Lyy8D8HtP
ERcyPYBBGn5+TFq/hlGXRBfZftj1GvhC2DEFOCEICtghRvofy5Uc+Cw/Ys/3eR35
4togW1146fGuRzPGAE307Iyr3/HZHSODmyy6nU4sq5/QnbhkeqdlQfpoU8o6DnRF
ohBtl+ph2z62d2cPTSq41z7pAjWX7bhEV0bgAgOzBhJ8TAKigJn3UYz4+yz8VzSl
C9a4/8JlGWtMfr40ElgdEi5aU4pc05ldP1SWOwzaKSv7/J5HoHsEJdXNs7+PtjdL
QwZ/pc6gJaWI/1e/0CiFp2RH2qOl0qF5k9uZjiKFQhDyiEHF6JjwL9IJOsLJLKby
NyuFBfDGxtyi3BP0Pv3fkgY+RURWHnT0bfIDu4J4Q5+7cSUwUged6ytjheYwZ3Gt
F/JkxeTZ3VHv1pYpJcBLxwNKEeL5H6HW5RIVsJZ6wT+KZ46j/En2tLZwzq7dHmUk
ox7IEWuo9NPUqnRds2T6k5XLJJMjbe/MDlY+K/5CYOz+YSmNyFBhSD37BLjIHzPp
Y/weD/lqNxe5wITHNIoqaP9Kp9wOb+OXblWJJj77oVJedurIIT5hOOC4MJXjnQPh
hbBD7jMapgbA+SLA769xLz+7pD9069WC1glb48oEyhyAomRwxNsCxmhzFwi91k53
LKrUt4fJLiqMXALRQ4bCFBX6qq230qBMQQjixr9bCmlrcbkG3wdbEMBCVr1e9dfD
pJIg0cRO7vVkqYCyYa5gLipWaXAK52ugUAEuEgS9RLJXg+GXjMzGWPRsxmien5Ka
SebmAo+V1VP/0wTuZkVF9v5xDb5pLQDDE9ezKbPWOFlvaANGcsI6+YcUBqA4V7mH
iPaNKDWKBA9pHBQymKZIRKo2jM3PHJg+1dMNYai3cpSjuPE1muEtXA4HBp+fAwsI
uhZo+cEIuWbASlc4f4DpBZs7Dx4eccXihPPLXQYc07coi7VNyEkMONWACHsTZjie
QDsnVDIXp6mmq7IZYLqRbLcmkkPn0Yks+7tLSf+t4acb3wxR4xeNU+lBC5mDWFrP
W/WGnL3zNI5OpVVDsM+gSNxqBLXONqV3slJwhJ/l7Dy71L9pemgDlIOYs6ngaNw0
+EEFH2166Lv0G6+AzJioMLwdhn2FuXypBl/LKbsC8jEhKwwQbIsGzncpdNsR39E0
wM+GzApKsZsASt4ATYpMOHiyKjhkDnjF7pzb2fAEb1zlWVUihsnq0sLjza2Hhtu9
MuQgXKEVIdyWPNmBM3FbZ3OyJwrvrzdlc1Qnx5+/G5NZtL0c23Kw3DB1sUp/ugj5
OAHDs093joCx62JGCI+Cbu4Jikeg8M3SJC9+cbcAOPM1Ioz8AGPT2NXJofqwnzb8
eVx3l8d2njLyoOnVFJfnpOuK87wFzckBGgK48BOlxq/og99EY03zrl/+PZPkD4mT
W4R4+lvSxDsMzK9/0z8lvgVEY6oPYcia8c1g36o7/G73jNMPC0J87AJy8ClwC74n
DHRbynzfMoC3BGq/EcdIPKUF5OG0mWpa8tB3J7fI9s5pATuNiwktMGqEV2ECLkHk
6pEgtFDrDNAZkHAD/ihlGc2m+isteKd9SLfHxGY/1oXzRGPZoL/5sI4fR9PUoqqz
iuNbfcLMO+/dCt1cJK5Bu2RkqB9gWbW3gXECRK7XEKZ8eSqzprHWmnVUVMpdurdo
nW8dQUS+E/8r765zdgVGxZSLgjTFJYU5Lbq7BF8hjF48HsAWJIAJ7AaqhevSoiFL
aH8u86+AcxTnJalNiyuNXGX880ReHD8LZzwlogxNlPeAHU3+zb0FX4cWoM0VT7sC
YjdenczHbDEDQWu/DXlCW3Y4nL8RmaBapLWdAu4gATX970BYcrabbZx6vRa4jeTV
/R9gT9pdoRLwPDNfe7XKJikWrp9Qd446+bNwF8i9eD+UwcbtH3NsA81zC6Pyctmk
QrDD8HtdHrydoLGx6p4Gwc0jMYGHDiaSAc2dEQ/swfa/9Ut3Js8vGpVJr/weQZGu
dBmV6CzBGHGBsBi+eTwuCb/bQgl1/S9MGp60gM62UCUUIFtL29olxdZbzBo/6o97
Wc8X0sReo9HDUrLgwZ66IqX4t5rlF3uQ5kZT9elTosQGy1TWGWxad0IOnhRVppwk
JXF61DCy+f1yEXKG8RRA9IWSO5uzuEg6nabSdsZ0Qe0ekkoICo0HEfeQUucsA3mc
13njMTnH6Z96MmRKJ1a711FJsS7m+i6aj+2kwde2ZHg2ZqDF2lQoXplf1/VzVmmJ
SlykL/k9RGdQWCIpVHj0Q0z4ry156FX/9puKrLFOhlmIXQlWXnyzlbUXzQyb9Enq
rJrHb4v8XHGU14UlNgWBYmMWu5NHtqQ9K6oFsSPMs1bHaxu4OUwj5PZt+SH5shfF
RU/oHVAsX6X9st5eCgxCRA1n9hSxtlG8Ol3pnmZgJir29RWpoaB+dbg0rWEUWWc+
Jx1y6q+3dkOJXh0/8ZYOeovL3bn90IfaQFUurb+gj9ecjehZyfMdyQT6UxXbnkwK
4iCFF4jMylbd/JIv3r/uVtvWBS7fVkKSjiVMSx69/E9gSk7ltRw2De0nT7NpPEEu
7u57RfDQMbD35sSCzeLkKTgFtaU0UiBZua0EG/Ycu4wxJj9AbfFt4urQxstav18e
iInyr0y2t5SCdk+sl6STH5NXft0vU3iIX2UL837MTw13i3TMRDBTphbUJNTtRVcp
bGI+FNflFxKWMLN9TCc1lZekeiWa5tWK2RYNailBcTBJO/Xl4mCfuqag8nNQkrap
UhjpdlEw4gtjEzpiZxjITzepRK67Q4JchwPw7JMQgMgvlkh3WLU2QGZ2jNI6pKNZ
2KR4ual3k1iMik9vOieq2IGRfdYVKiRjOd0FJ2GeEn7NH0kfYY8blPQ4q/G7xbpy
jsIufkbwoXA23/zMVCZAOJqmOPK9Y2QW/90La3HSRBi3+IeekK69FPCaMhsgoNkg
HkZLhF4M0B1PvaUdbo1CnFpaFp1j9G3EsqEw5uVuH703z7iAxAn1lKKcQ7u9i+q8
8ly9fC2Qe9Ru/zORoS+JustnVSXKiUDNKR9FUz3cZLbFYzE/4dENncj1qd1T7PiP
vH/0hBLRceppaNQmCeV579CJuCYPzpSqx0NBOSQ6dnyGmD7ZEfwiYTt97zWMQERe
nbQNDwGh3oTI8W+/xf+avQRbVwAxBbFrqoTKUXlAuJz0q84TyTv3stAFx1V51rLV
CXIRIFbnrYHFQGK1PI5wMKrrY8VE4CpCTL2aHmxQzu7lVw1SjH5nuKnyfUEALmpT
ZLzV0LSk1Cp2v1UH6CwvKumzG01PE9wC70kR5UMrTF+Fp4W/TCxcPOlEceD16UZE
zgmopWQV7sKIkc/3Ix0dXIVvYQ0boAQeHjGanNyd8dMOqoLR7MMNEBmC0owRNRDQ
aCTqPl2+Ugh+n5CYD493rkdmWtckz10k3SFs3hzxK4RCLE3I4CMF28b92eXuXq9k
KeqhWKvRMPVM4nbKZKytgNmrNRjcoxVb54Ygk3HZy8k40qNKmFBcCwmghfiWH/Tf
/YYIEFgBU4EKsA0hpcxcCw1svIFzJb5ZiOHAXRD0hMxkJOZwgigYWf+Zrzxwqb5z
BQ2YwyjE0mKCsMLnR1OwaTGEZLzlBsiLjbroXOJ93MQB4+yeh5hMdZVwqSaslTGu
kCt7tXkz1u1Q/oQ2meimNiRolK7L706+CPpUemcG7D2s7N+Zyf5Z3+AWbBkhbknM
sNxvq8KNIgs80/tj/481YnJ6yGTs09VxX/zY/ra+JbaPfB1PqJRmhHmWTCoapC7R
dbypPzLkinMcpNF/hYjrHloUOcaGNACZw9ljKymk7i+g9L27cVjPEQyM1MEeioix
zbVmd245IEQ/PueB6ysuLlzLlbXuvkPm9LQvshik43P3vuAJgdJrRcPIsfoOGU7f
P8B/7+H10Ih3hLhGuBW2MJCIF3+oEFyoSrLUuAsurzQEA9JXpir6mIEuqJ7+zxDJ
GG6N0xCHlOR4QwwYS1qYvqdjpxfGgdYiE4smg36SLzNv7hmdj+ScN4cHwUIe4BCs
DvgghA5g7fzzI07exafH8KWgHDvOnpV/55trlivcwXfISbpnsFZ4+5qWPndLAWI2
z2fl77GM32DFdxDD1V4RAWXnX08EtkAAwnGs0UhIA/TEsvr5xNaxCKIYQYGt5Vp6
A3X533AYKtDQ2arf4qiDdShMouAExyX/LKlz5d/n6rLRr6Z3ynsyWgcFBpBqx1jH
VRwOC+pVFDOO6ui/sfBiBHL1+waczAqfWVPPJjjlDUgWuuXqlHMi0SN4vyx7V7pP
W0Hb5JnWaSPF1uV9VHfCrZZSZLxQ/tItgMftMyhF6Z7pReAR1CFWgrjNBpGbks58
6DLFBh5M1jrvAfX3v2eWnFR8ihiz2/I1gTcHf5/9roFunfweY6tJri69Lrc1YgFm
yJp943KHMg7J12pH3qHo0Ju07gOafQmju2FrKgM4hac+kF5DJmVAxPlGAWaP4EDz
H3CeAgbR/o00qfKAhF84nfMtJwlgscVhoPiE3YDEKkDNeydyj33NdTkzLVzgH5+j
ivXUoEsTRET6YMu0Mo9TulKN5q4xPnGEbifH8AgA834pB0uwdH1xuNQ86hHrqXNo
2NrT7brxq+u8Ns0SyjZdSstS/d6wpxoUSKk8R/1ZJEbWmwGTFI/6rxviLTT6o19m
hV1wKLQUtVLXVAWW+Qj2tsZOoV6KTfr7kttlLPfpLLQudfqFzTZsir5vBaXXyugn
4jczz2WFDdZ0oqCvpY7MPWy9b6TXkjnqXBDMwEw6ml5egz8a1Sga/LrtGSxSyQhz
nkmOkwC1wzi6NZLPUwSmaBx4RaOMKaXJtSPCmN0UiBDDy7d/o4wxvu/nPwlypVbw
U8onHxpN4v1hPC0Lr+7EJ+wZjCUV5d705o/6svkk8IaiJCOUXBlqU62VdVx/jq7Y
ucGjcLamqOpDHZWzZiTyfRirBK5rfsK6PJEUGCVwtEF2EtOcXSd+yRTuqXVwDZ5p
/logsIvvYm98N8bDyX6dzaC9tDPrHEtpFMXC/s/I/AKfGRfntwJKkZ2jm7n4Lrx9
EkC0rDGhpypFGMju3wxNCr8eWU7cPKAf1t61qAB74e3OyCxfMnniIi5AxUR7SMbH
f9tMGE83Yf2e6TLO30oihFh9rZpUiSZa9OtxXdkyTnJW5QiZUPS+58/IMjOWNKDP
fCjWosNLOPraBSV2tm42Kpb+81U9vivcwzgvOEyBQ1sOBuotsOKFYlcQUNgIVUWv
xc5YEwA6YLp2MnWfWfaH/PhiZQsjta9UWySPKJvZlrEK6kYL5M339MdaXqqx8Npk
5FIMSxMx8YdlAsCVKjGSMqhIHeAfFG7UDkZF5LCgX6aCHOhcVCX6gRb5CGv2JQ0j
lpzqTtTsHu6nnUzEX/GIY4HoI0BvwD9jzyNjjl2Ek3PUX1RxScyZVqdQb+i1mJsy
/Ju4hUwUVfk/8VB8Y3CNJO6HFGHsMYiTIMSnXo4AcNNLKjctHoSq01pkDA1100zp
mjwy/cwf97zsaXe9/d0GBE/ZeVtXiSgC0SPbATh8lkuZloHwXw/j6uyaM1fn98Fn
b8hZB+0XU1b+Tz79XqZxF+UTo569zzyJBSh/XJGJhe1wAqbOwlzxbp7/38xpMarQ
PFSGLjkbu+DIxzdIegos0ujZd4VSQRBIho5xmdh0zk6ab+Ufqrn8P/tlBxreD0hA
ZsHkM2Nmj1UI/od3QDndsStFi0+eJh2EaYINHVlT6pmcnptV0e4O2txGuxtrmGzw
OSscPd0sq9xBaQco2fa/N2QEdrd+bwQbCRwT0DF5R84DUJMhfOO3dCZ9oeTZ6fEl
IhvnFYRUNZuz3YFij9b+kaY2jm/z05lglIY7arj3fvBQzPi0+EiYB9IiZ9p6b+MS
f2db+VDS9bxZsO2RIgBQWXJdrWbNCvMKYKk0rDvmegJQvJhCHSMYwFwETjRReqoA
/9InmUoizzDbgSbubUJrdeoTXxxCKovyF2WTgdLZvP9wx+bDq8lPgvWeE7Yu0CEo
W+9tT4eisfuYk3YMDATeerGUnY48S16yiARqZjDHr2PZjjVy4rfRu9xA8p1JW6a9
lgY4HOuf9HCC+fzSN7ORc4sQ78sR3pFffSS2b6xG2j/k2TnkVAXTED+BVE7u+aZs
mTNb2kqZj0i0eOzjF7fE9sC+sofy4gveEg+vd7/MFr4ejGg8Yh90kPu/3+xkPKfA
cXzan1Cgx8hg1t/mgfR7JA281KoWq+uWjkVISUhvR8//z5fP6unVwdBLwq92rf+i
wc6zvnP/KB6pk/YzTCHyVgLtOnBvG6W5Cqnd9cslQCRlVLXXllYWHZwCpXDGIscu
G0wMOtkfmFwHK90r8UQ3BCDilZRtz1NYlIHzG0Nby4AklM0ErQxk0Uy9bwOaLJIZ
Zgv8UH2/ALI1AMa0OJIteUzoF0zsBVODs/NVGzRDyLcE4b+Grm/XdaZTuKsnCsDw
/+q6TDEPrfl1NtWZcdyuIZX4hmvTAvvkvqkhlx6mi4Gvpp2K1lf20NmhXSfaFWu1
EeUF2SNrVo8QIN7N+q/68hC7ihZhmaXoInosLs0+SfhpSsCs1zlPndu9voKrxYbU
07bwKFhBcTVDCjZBsvOiD86ANXdI6bZAaSYt3MmbN+a6SlZJQME4/lGdHe3ztwTd
b+Rfo/fzbCcYeobhah2LpV3Rp0yZdBCd8KzUS9iJPyWLYFR+n+hVe8u61XIsU28h
o1GsJDGTOXTaKiTR/VaXgJ56dVatEA10PSPAH3m73puo6/L+zXbC0ob0681R9+DX
hPCLzGSdRQQn2j3a/76tSLZfWKucYW4mp+PAY/0Ao29/e+7dtYm/Ter8wTFFJd4p
ODJvJAXNsAzKhBkzKV4p1JkCICk5MHBXXLzMB+JVU2zZouaq1dlT5J6xv3N3V+Ly
j6i3RH5uBe6z4M3DLlLwCDlgHlkI6Dxa4EOrBvAGnZSD/JkVVHEQydIs9D44D38L
BL0XRIP2FMOQe+CBsHORXjzPmETetKGWRN1Aabh/KMBE43iQCrbhRyPLhTDY/JpJ
cimPFLt8AWP7nqdm+VsCnFnXc8+DW2YHYmRYkYrzJPB4jMSMWx+V5FVNhR6JkNFe
6csTG6ecaWPMXaKKwJt1Mc06N7zP4GsD84bW2ryXWeNsshPsCDTTexKL7Jw4hiqb
KtJZXa3DuVbbpehh8tVNIu6MYjOa8HWG7OcOwl+xCOMFkQvRaxdvjIOWdi0KBdw3
FTMiJ891Octom29v0L8oVQFy+qYHoe4J0c6/wGyFY9rjx09wD0FVcgh5LCXtOPyx
I1T/wbEbwdJRxYPs664ScLI7NdFbUxX4orPGowgB+iIVYfkDAFI6JmNAYVgo2NIf
+0arITe/pP3zGOopQIr2o5KujuafCS+w+8S/A3HmFnuJAcuUhPW0xSlFzyh+p+LW
OswVks3DC7gIixmZHk+Xp/OVgqYZN+Lai0zZb2iBnwy7aNvI1hvFMoI9HyTeArh7
tmYDKtgWcGX2zY9mpVPv43u6KuK8gnfm81SmrAfH7u9MjcQWIsu6kXGy2NRK84Z/
MsaXGnXUpdrRg+WPCcehcxw4yF9ar9O8kMZCgfRLZL9M0NrlgpWTHK+ZCIXLe460
rOiLlIARE70t44pWe4yaKxG9rv/KZzSHCOMr6F8c8b03ElVIXrumJWQWQArqwGsW
BQY1Wp37E9GMGTC1Ex39uXAi/oZSZMVa8KW4aIDTxtxB6i/JNmRHNLXtf9h0kLFt
bPYGvHzE/U9ukCCHs0733dkNTOwjdey0YG5zvzvhjbA6sIFAevuuGHk4nDVCLWaX
hAcrl1NjFIqcoS9VfSnzxI7+xLXV1bQyw5K5WQXzmOFh8SRFhBOsSwIwG7Znc4fx
byqM7U0ykSXMe0L3lOA3XH/8zYNCEc4T6b/YWIIYpCaOuvriUdEkafIE9/zwJ/j8
ncroXCC9CgNso+Xd5NRw5fcQby+gDUfeHUw99OGBunC+sTMWHIi0GGZ7fEZTqiDj
kkjnc4xqcHaZ34HCjuvx1tYklTttkASBgSgscIhUwhKiNbzUF+LiCZXSdQ9KPwDl
id1C1XcZOTNVRXhM0IVyEltb4o2aWJZ0kda+ipmN9j2Jx3+HwET99Oa1XbETVRCR
gJQVHiQBXDpoLeBG1IYau5uAWU63seK8yhkdXQ/QzHA++eprm22WQpIo7bi0PJBr
N9QAMEf0A464dMmmh6Q5jDT/OtNQEa0VtM0ERw/2N1atUlLSlA7VCeqv6ya6Ump7
9BjKSxJNBrLAEpMEpE82Kr6vKIfNqDOxueTSIAmjol5BUXxqKhBhPsXB48Vx9e4c
AXunyPGFYJk6I94BAoHl1R/TgcjspuwRnN0rcmOYYra5l8dkznKqtJCVHIuIEAy/
sRJge204WrfP3+DN1PrVLHp/S+sbT9dpw6fq+NdCrinh/ppBYxd2ibcqcUQEGTrH
5AsH30H5FF4c+zK7X3yxgaO7h0MA/OeRyBXS/5gg9w41yCFyrM+2aW6Twa2R2ZWN
OtQD+Uf+Ot1HwWL8501154RnKddgTkELnWUMOuJNNHJ6yfZLLupVPJVORk6nVrEX
irvXGK0eRo7uV/PjPYAawte4opnBFRHUbsR4PAxLcaVT7zpWeDIH5VmvyVQCkLhF
qolCCh7AcASuHrBck1KVsKqJ84rQglRVeTbXHYu/0+GixUtTCqiiuf5BEfYPOMQh
HEXzvWkjupN/VG5LpCmzVMHwN4FWoaRALGWqwhGkJ6bb6/2W0M0S9FWa/wuKb8yI
+mPs6wdsuQmf0CmnSsfzNusWKiO+bJv8aJJ45oVm77lE+L8H/vsuLQ9hMwKSLQgP
9s3l124YyE2U8d0VdMgwHurc71TPzdzRwTdvptUi5vtaXpqPDDM2Kp6hm6eNkZe0
cGRxFGmlDdQaSUBqCqdXo2RRihDx+dHSyqpzdbJFR4qou8NJp/p4G7IL5p7dI/WS
EyTlomiqdu5BbAzwb6GtuA57w23v6s/55w0Mk8Fg7SpsD5DHsE9nKWKDXC/XPhcr
JLqgw5L5/gIRgebkseHA/15eVLxgm6voaA1BstNLSNOUc5CapQteUUcndZlyef6N
3BMDjynM0HFENAcBBfvmXGJ4arEFK2b28n4Rh7xo5vFy+flBSMtZoqCf/INFmEie
vdFhT5r6Qar/VDet79bf/E8n57WMJ2G+YB5M1Rov7CeB7ajhtoPYX4rFgZv6wtP4
nnFs+04v81tNH8PoxCEwZUg21tk2N0sA8CDxiM9fPHvLL8acP3HYW4+z3r/2JgoI
0YHWQMidOCLNEalGgZcjgsRenF2IXcLaph1laALkdpLonX3eqE/Faqrxny3x1DcF
aLISCVq/4ypaf8vVHz2VkhCAP0K+28lqNOy+6NdOT5QLxUlqVyAnX7kVl44/XlIb
7NynAvNGDHozeXw1758okG6aL28dnpcR6fUc/zyDn59WUbW9uSwylsposA3kRtZ9
nquijVVmg2pLfuX1bmQSi9BrElcOsg7V8eYUyfruY11OazoWylTPggGx5xXWH+8K
edfHC8cZRH/PaYufOeix/15sSOPMYyhhFk9lEzQGvEokgapp4SDwJDVvD4LD06gO
fYylbaXSWF5C3rgM+aGehKbUwEyS3d+ph9m22M4mVdpPfjFaMnFNadZmIooDuNsR
FEWk60gIOfgur1xSFdUSX+zvXrrX4gQwHu5ipJEid4Qp8EmUG73tCGFn8pLSpSM1
9x5ELd0DkV0+hIyQ8KpKJkZOD65VPy8UBVh8YOX/c5GoSdyXLNWeWjFspCwjiLYO
81C9Uc6qK5xxeQE95W9gunWz8ZNhNmr8PnEL+4T+eKWoZTMhn/pA7FytrqQqHmRV
T58H9gX5ov+LTUphQz6omQdv059N+5R3JCxikDIGY9QUgiz2MD2wS5yPICaHJbq2
S7NvqGLzhyFHCArLU1mIT8GUHQiftDRUsnnRVg46HwjkcoH6e/SKRbwQIAzZTf6u
KrhksHmxTeXC8uJpaJg7rMoj/GFriITDJHWrQwapcH5TK4j7ECQ05YRak4DGp6Hm
sdBnVRtrc7WXeWRLcA+M1yNRZH+iNHXzSNgTMdubNBJuA9Q6txjNeg7SDfCsZ5QW
OWzInHNeUsaitjAl6yxvKrVpryn8aQ9r8Kuv3NdKlNUwetQ3tts9j/P0ydrgwEhE
KBTEpbu6U2oYZhM7l8ewi0wUFI3LkDJMR60mfC2mgrEv+Hd25E5GVBMLFRPO904f
PYfBsXwuyrKUeQoF+TjrLU2ufIgOeraJfFz35hQoBLTpSXz9oPjaszVzI/svSHnN
Tz5vFqZB5cTj7U3iZ17ohBVhAmimwjsA9N6QW4Yrp2SFoWoIOYhDJzNh4wUW58NH
Uk6zK8r1TqtvS8s4lXriiwMOYxqQ6lvJDtJL0Jg7+ghfg8mgqgbpQq08pfmTeWrH
lnPzCQnB/gP+UA4qO/W4+7n00E9ZixwF+eU26Le+gHPLQ7d9Ln5BvkLM68P8jfxL
9sU5au/Ed0yf2D91hkfKlKVeEwyp86pBUu0nwZsswv4uaF191ZRuR5KD/l+kVha4
jrcECGwOQmTht7rxSmPE+GMOO2If6ml0n2dYjhQCnMxaD9LteB4ii4OC5z6jjpOV
7cay4fO+jAm0xJL2Wcq807I47hf1/8TyN+COC6KZft+jJqcdG99ap4Hg2Jw3uy6f
mNp4iPzGtqMsLWuH3CarnDIigEaM5MaQwwZ8ZkHnfttFh23FsqG4RJFVx0Dq2tbx
aYEF5As8Vm2eguopuQcFVnhhannN5SS4e19EG6dXOsKvjufkhNXOfzQKZGRbqDiU
jYBTtuUYCvDihs3HT+898/qK6xIIiunKtFsznwJ0X49WkcmyTA1Njwym12nQ5dY6
XrYjJ/rJ+1QiH+OXoLu5F77CAiAyPoJhQ0im63enjHuQXDrWoi7zJFoRnk5G8asT
ApXXtJvNtF2Vl8ArbfN7VfaIvG+3kSs8Yr+oPFM0JbaopbJg0BZRn7eRyZ5a7Wt3
p2uvdsfhaQPOWXrLf3udmvQAom8cbP2wvBLYfG2ZzBLxR//0qtVSbt5m6jG7V1tp
dDIdrSrcWMFvXOR+JhqMLU0QMayrQySptB+8CykA2n3bpMgoBdyhojKA1VtcVBdk
2VZkoqPio1O+wjyEBBesNCRn0KI3JtazYkaz7DybakvigBI8OKmhRN3lT4cMrgno
ENa862w+dnv/uoF4r5KvhYizGOSjwvr6XCYScTYpcF+TKp0thXszOah3YE4j8CKd
GZabLUXSZxh0ZFX8gGnXvRUIhDCKkk7pFmyYWFMT4ajGKJUkhT+TDjLp43Z6/W4c
0BKvLlDPOXMmS8PXDDL/Xgu+TUhFhrMKt1RBmxiA9ECUD4jQtLBwxZ9BCeHAaEC/
FMX7oQt+mnKePTdK0x5/ueJcooZ2YmlhsLrXjo4mBnyCh0KjuKMdzVS8H7PFzuYI
LLQhWp0H7mBx/kQv3YowM23zxRECgyPfzHhCXfk7WGSABQZDSK4mnUT4WedZu0NK
/qTWl4TUhh+5o3b8Bl73OFCbTLSoDB0UCGTv3UwhTYE8K5X7p0rrg4B7it+UvBN+
pppZ0AM4BRs5kijRWgFFz51sxptH40TVehOcLP8iSUraVVyI3b5ker9VtzbHqC/k
rFULnQanOtOH0fclKQdVg51pRFVwgLb6niDKCiWS+HJgTa4lJfjw6Db0zDlATcjn
A0lLbMVe+XmyNVlSKlVqZxwni7rUeC0zm3XylPhmB4UXkclzO9JUTZ3aGIYhRvmt
VNVmVFtASp5VcMXVv2wjXf53SLUMZPQTmJD5MR3UyuPb0EKpNd2nJLh60WsdOrUF
8aepzax83eeF0wQpgcC+qAm6T0oRlUKfpgnRiRmSpntofa/Km0GsRto3ByRuWG76
wvX8MWgYLgcoStt4506Inq2bDhcnnwWxCc9ise8skIxZMJKTa/aolwWK8Cextc3C
DrNnE7DhhDxN6DwOBpJMMDAjUYFLCjhoLnsCoGVPHPoOfdfkzb6clqh7wlB+N5Zu
wZt1dK0cdJJ5m96xbG3xt4iBgGROyEljpRZcdasP8/hDrWrs/DaDDo+NrCLUaDuR
m/XkFG4dVMCCCmQmBClesr0qDJLNRMqI9/EqtppVNTnlf6+d9V0nFcghhPNRP0Yh
WRGC5m4kHmT8fOFCnygym0gokUyUR2sCTseUIvt1RH43cxUcEPAXKggccdorSjEL
vQ9OUMUpUOruAAMYsaAHecym+zaK8+tmLVGNyxOVdyAY/xOC/tBJjtpDrvenigdr
ExArkDtwY8MrDdx64+GESpV9r2SVTxvo8W+yXzrBqLCVPAcuDqrnGQ7Kw4CYNJet
LByHUicd/TqERhvj+9HcQRKy4zlcgRQyflyvq2gzCvLvM6Ts3KFvOFP0SWoEz7P6
1bLoH7dVebtLzKxgT9g43O2wypFfWFG88mdGmpF5TeWfgK9IkQ5kih1tAqOitmNx
+47UJ0bVcaby+gf4fk1dJGmjiJIR3KrTTrewNg5f0Lityx5Zj4Uu9TWWr1wcTUc1
NhWM3kDgTbrETfBPrNh3N4Ry7BJaMrm8s84jYKaDP8X4T+GQM9uzmbos+QUBBu8s
rGR9wUKQesidbhzP3KkKOKFEG4+YiXGYWJIK0xughIFWRcIdZ3Cy31uOMYTQPi8C
GK3K8vitVC938SoziLOF/mu4LWDfvZzu0X94973C877CB0OqGhnq/XcOWAqnLQZ7
tp/aEBH0F+Eb05mQJxdYJbvGngkLAF8QMCSY7uR3bzpLUutqoMNc/2OdmOgqQLR7
Sq3EM1bQWUFqGgUsDxCbEFC13f4d9AlNkj9cvUDaW/3JAafx8Piat0rzEyQ+tmnl
b9yS/vJKX2AHXjCCHlzLZkU6ynn5h/yi3MDu2eP6bzZrOzDtx3CxfuPZ6oNGhRYd
xm8tftwK9ykMzL1cPXbOLWX0Gr9nhDHQUnugZj1+Hfn3E/3ahfZaQEw3BIaMk3PL
eTd4wymqpVHhM0yEFdOTst26JPbZTrMO7l195Lk3L28YCcQbvcw/Wk5mLCHv3Fld
U+sxoqOdqGJxfagaNCSbATYAX/IzMXGqT5OaRGR70vcGYd/TsNlaGsg2slk2xYr2
YZXVCa7+j7SNEw4oxHYJrRMHq6KWvJX+kqzJRv8u9GysMH6P4nGyJQSSw4Nianak
aTC/FO/WuG5YpOKoBintp0h9SqZayram+SmS6+UwT53mzmGzApePpby88LW8W3op
QVmSlv7He/pXfc/q/KUN4d7EazBrWN1VPnoI20aobSgsyteZWKmJ722ArG5Onb0D
YLDasufDt87grvYhdVBByOaaXV5QXh6zAwEsuviDH93Nhp/e0JvmCXwAt7R4NbRK
lnFx+pyn51dtNjFtIeOny1vJSxbURpiJ9ojZUpOeakOVdLn72zfLpXenid7rYVaS
NjLTUhIW5KKPY+1v/3UjmzFyUbJ5vZehrBKcDn0I2dOQpFiapMM0DJG+LzE8YhAr
lqz6/+DvbGflFRuAymgD5vfJdVZrQGVW975ivb8jdWY7f4Vja3iTZe16epq6ovHo
gFfjgHGETWqvVdwa/+GxGIk2I1rKYNBHjG//bKdiEhU8Qu14AFmDjfE2wLGD/PdC
cbYt2inNOlEESjSuCF2jq5zYjNHNRNWy96IsZzDW0IjhmauAOjs4ZSVUZG3+s7MX
waoM9EIC0JyhmnijBHJIuEKMQ6nCZqUrauvFL5dGkcONOt7p+Y2WqOocdDD4NsCz
8owrkJYlCagHrcR15EbPy6iuBZLjrNZqlRsYRSR0AY1QIwVnMCvY1SHXGqaZOgEi
nPo+0H6s+9na4Dob2E8ehwBaHxTudpzZOs3uY63Wd4V94HnEqEtemycpWuekCYOy
8WLf8h71iQ880zXN4Pt/j4OgSxB4/aBgasu9mNrnOdoF5LEAAiQ7HAQvaqzPlZTG
fbxQczp7F1HXYAOJHxj7X+x2Xg3OZu3VCMZYghXJKGM4V2tD8xwbhLaxlz9CLTzA
OX9G8Yq5twTgEzT9SIaIqXyODLA1HGvbsdnq68bSvKs8ymx4tRBT0bvTK46HkOwJ
rWwAyAx/r7f8aL21jbex0H7QUrd+qdBOm6or6aRrf2JE7QGwMeTSzNmykge1r0HB
rMxrk3b9D9dSymI6D7ueBg+shdsquLYZufJmJtD2a6rymhYewym3Chm5AmZcPk0l
UmF6uIJKgqj1+GwDoSeo2XjPahmuUaaXiP2PVe1wCY+sg3CEAf41wDWldihNhbYl
kQAA7sp/UpRpwGXuF03yQDjoAgZk5JXVakwGBfMf9gzPcIeVhOmDDBgU40CbyjmR
eylUt3lXq+5YoquvrWpTerako9jwFU2RYNAMPfLohSj0X3aLN/++LFCrZitNy849
nimgqBCePI296P59NL4vHpxc1vkhApR7iO+plK2yApegh6hg8n0VUTiJiJwImZsp
GjX1jH/nBWb/QriRFBVf/jC37BO6jL7Flfq3gFF+hxZJ/ACOn0sv11F238KCGjLI
t11vxUkusIoz0Z85a8/BGNIYxQs/Rz3+x45h5CLL8YoAhF4LjZnUDww9dDH3o+ql
knc8B8iUXRrqCsaLdw1NoVjq18qMFfvzUph+7FH56dZA41y5oW4TkNvGjLU4U3eQ
QB0jOywUfIgtTAZnNF/dI5RN2DYvhbjLWLgKpdkw2P4TO89my3BAP9XWJeHEJDFt
n4IAGyL3aewz8YzQJSOCBI8qZszitSPN5R9d+aKpT6IPcir+MoWsYRxj6T2bIHtu
J8cFzhSqeZEGQ2qy9XzM7IyddlROakl+vXs0yJ0ABcd5xv5fj8ofetRsu6RDSm0A
lO6bFeaPg713Serm99dkmAC5h0pVeFFPTTWjGcN062baS1r2BcBqKaCKEv37Lom3
DxaAZKxkn895gPTJSuHP7OY5W5DSANtw/LJh95jh8kfIMreBmg33eva2w7iNZfKs
oFgEJRyskYvat8Ae1PHOt6Q0LYKtmPq38BxdtomBARh8a5K8wW9fMY4UB6NnUy82
vWadWfVCPmnnbKSVrylX6UpEEEqlRzwzXKHJ0r/nfshEa4SGU8OQfzBffQKP+wbq
V2RfaS0fNg0FfWfptzVZTWKLlPSlU1LPfCfQCcxyeOFk9Y/c3H8pkwDVQAY95D/O
ZxDgwj7jePZs7BdlSmxA2QhVohf+oMa/xp3EKaR/CQx2F6RkBkz/T1UIuB6gXL1J
Qi85DsteEOF518zGG4K1gctijVfY190zN6idepj5KrNX4PEd0z7dKUm3EfaBzQtd
26PglPSFFMAXkNVD0EfbcWECRvbzhBs5623VxqJYkj4PlIrMVNR4G1RfUYKn4byY
PbD6LDGG6XP2WePqm2Wlaw5tuyYv5mmAuLX/CbjiCRupcBzyBXq7u3ms84bnFUBK
UXE+z2IHi+xLYwnwYM8vxDoL3hylptKhb6WzsztBusM9it7jfcZ/PeOdXopJ0vWq
1p0NZogfIRQRISRsi88iAcal7rV2Lx4t7QowNdISgxzRorny0Y0afZn9+6oD8SvB
hxPbS4DrFBWROE8zocmqCCkG01Sf5nLE6zGkEU6tOpZUchbwrvJn49gk88n0hrXe
werX0V4R/dpdWFSAsNp6BzuT0Ms1S5R4kCGSUJMvFptT+hMuuSpsG5ie3QW4Puwn
exGISn2iawCTodgr8jOJR3kRHUtdUJIRy5H98+ZqxpjWfi8hdAZfAym5HwMP0YrY
FRUKhFc7KYrCUGXp7a6ZX9IObUkEKpeZyj9UO+K4OlDm/hsHbqAdNQTKtN9Gi87r
ihbvAr3FqcO8AsDEE3xG8p5zpVxgke8X8DkgYz9zWe2BkEvzfe+BUc3UjGcwfwlM
Dn5azC437ziZV+Le3oucsyEbF0FQzIoBSibdcR6EJ+ojdcc17EefZZtcoYW/DSQh
fe/uxwYWtKjJYu4rnsl7j4IWol3eWgZbNAlwjRI4JIl5snNlJ7j1s5+sLxcKrnoQ
QAHBH2y3uQ8Zqua45XQ5FA/ZuLbQ+3rxAWe0E8YYSDKebWWa0f+ESEdVJ89cIAVC
+Rji1RdNYUcFj1/AnYAv0brUWOrf0i1Kz3kXsDv4tvv8ksHtMn6osoEW+gAlD0W4
Q7wiaWRRJmHEBfyO8zjjrCeelIXcmE16CKI8RUNojA/QtdRB3jBizM/tHyTZqPc0
XM707fFxwuEvFympVofmjzeMGEiYQgSuJf+h5Wu+Ka/NHWdwBR002wt+QOPwM9Im
qoGXuKx7womim7iG6Y3D7qkQHltDAXWiqAqXwB/vqbzz3NEXu3nzj52keiuL3JI3
wCvK/bxD4te54tDUkZmYM9wqeNJJeI/Cas0Htq3K9JwiJgpbbRCtAFw/1T6vWDaj
+D7T/zqYZ5nB5org1QmKdHLQq7jVfeks2ssXqoEyB5uRmg+NABKazmaFelvIeTn3
HFcaEHSarUg70UiMoJzcK3I4seYreODfmGHJE6OuAZVbLRU1H4XRsmoKffheXmvO
vBM59Ae3kz3J0Kpb1vH9y5Y25yBjozNO2JE8ss7JpnND8XrbWGY2AuWyPCtVRm4k
1ACcCiURkPk9VAPMNk3Wub2T1ST45g5j2yCHUOLYIeAaYQZtANx9wgPkr85vGkXG
ydmTmFWOHmfvwAz1BIjSqqocZgUrUtWL6R65tjrqpoyvOcJbHRK7xy25lIzifgDp
9pesneDr1Qg2hjI9He2YSTQmuwZ4iOmSoMLquZgMBQrLx+9SxcYKz6Mm+Z0tMlPu
Nj32LthEZctpdKpIqAKkbHGDixxRDC27aNjZK3+Z/q0WK3lrImz9yJ0xwLus3/qF
XoRQVVTpEH9+JPXy3oFEwShpm95q5jaELpjmUEl98XPGMZul20ct0lQOD8p638pH
oCG1vrVKCCW8VUODTf7JBGx7C5bheEnkGWCbAibKgYTefJ3MYW5JDqEle+Po8Wfn
b8CAWd0lg3mIaO9dw8PK27XpU/FQoMWNPDqln2gNHNva/vd8nDruPz/mcRO15S6e
1jHrCL42eKPmcYzauX8nzPNo0vAAaEugmA1UUBJ8kbg7EZ9cq6F3zIjLNEJwpB4P
u4CukUaqdzVUQgjSALYGKNNh3GmMJV6o1tfnkcR2yF2znVpHJX4zczXlERnmgGZd
EOFzthKX13aKUN6sGvTiWRfQ47p+S4D4VJydllK7tG89YGy463Nf001OdaxgpA4o
YGkVdaA5ERNP+j7kXUo9Q7z5Ev3sbnCDHabcb3jc3v36523Lkw9NL8wWkFpFS4Ak
kkoA5r7Nk5c2R5o3gsYZ44CDDF7j27drs9n1yJwkDXRhZsfc+2JmlhB96U2faoCw
GvCJAM0XP8P2dc+tqkfdoJNiAPhyRQeYPpLxP2u10QQEcO7LqYDYbeGQ5ykSTaIj
PWGP8oYD9QPU9jqXQ6Uwy3zZAyF8A09DryxdAteC2VyEaoluoJlm5ujPMOmdzxy7
t2WOSpXCN2ytsBsYn0BvU4Ontt3eQAVi09lunV75pJSznxdimUyDjtV0+4VZ43Jm
BsVY9ylzgNfoeBVb8T45J8/EEIJcZsAOPyAZ/q05QyniAxCS0n6Yaz/wWWN1+Gn3
/PtaEGxZ+431FZcDdLJmeRsI7XOzt7NVVLZriCZ/8u7jkSlOXo/e6Z4kPU7Hydyz
hQGAYhzlxuF15J6sD5Wf/z2/wr8L6Vhr4kHs9TnYf2LiJw02Ti+evjv2it36mbXT
zuwVE7woBAARw88LViC9H+eHe0RtLR0L9ZJK0OHzWg/H+Rt4VB81scETpVFItdQg
dOAyWv7y9BbuQX1NgcTlbHddqUQXm6PjI57he9W173HoOk3fh3yS5Ju+BCqBzdoa
jmHqcP1sBF96p9BHaIB6iNuI4+JKYqYv/TxrZohizH05RUosKlb9q2fL14hIxY4Y
KsxB2bg11vuqX6FHBfFJSq32JqkYWzwV2m3Jci3BL2lGUoZrv0pY4mW+jgnytxcP
gWHNpZVmGEj4GmrSv342Sq2/XcFhUR+l2jtOXNNBNxxJc+9zdKynKIm9/k9oIIjh
6HhiOjVSQVny6i3kckCdrLbSZl0BrFcXeTGJZawy9NjBDOgA8Icc2f3LpR7HReyu
v7+RN80ajdGEPS5A29apz+p1Eyqus+XjFYsCik9apu8k+tL512jL3fdFfv7ARAqU
E2AuKHqIbID5l1pUnTiM4QLpmehJmmYKVbBzXFUF05QOfGhT4NKW3B4+kg7CvOIr
sp/NmYEbQWbynq3Z4Rnwy/E2kgd67SBNcFa5Y7nCod3kctKNYTQCoMqxtY4+yWvF
NHwwOJE9oduAcEcWFThbDv47Vmjc3z+s7Qt5D3gBGnX3fKKFMVLP+GJ6WMlyjySV
ryVKzDSewnxdkWs6+OstVtnKSoM86ZlFb8M5c+os1/cjGDGmoTC0NhwphQDAUlBt
qvixi+OPhSoYwW/UN0uu09LBubuWcQYTChLrbrGIIo8SgA6/qoTnQqEZmLDyWTLe
i1LOOIRsiC3AsWao3JJQsoeG23m35UdQtvmEAWDQNiOj25JP0MrWAVW0kfHfdDV2
PKUdBooPXjoumWmDMqcN3BRZ2UwhQoasoH1B+jssxmR90rPcpBqXKTdfCUC4+25e
mfLCKMdVjShKnGwWDfAtoo2aZ3isTNUjEwyAry5ly1ii+ipgMbmYrDCvntMVe7KY
/NFd+U17jz9Uih5Y1IelyEdwL+CM8XQIV3/SYMGAKQaLQi56BRFOWhHY9WIoLhxy
vLMexfoWa7uklhSPM4AiI7rzAHYBEVZ3kmS5FyHB3RUrAsZzTI0O1Imx9WxM35qn
CVgUWvrOUb7/n4zdq6GguMTDJRgWFVIZjbt0qc/WmjQVlXDIpBOG6ek4au4hDxwh
HMWUnt9HHLab/iQaNJhw823B1eryNr0nzca+TuxAYVzd5LGAlullUQQuhWbMNkhE
dhiX4rH/RpsogWjutMWb5LHDVYPLVmtfz45s7Ja4NMff3OxlQGTydkxBoIJ/n63A
bEoyxWzbSg+/Wn6ROFmWmlP6XjngNGPe5bvro+rxdsIVUxONc/0TgsXKcCQyVel3
mntMvalbAeagIbwlcN7eHdwYDyFaNxo7i0C1NkUUCjwLvwe4U+DY3Lh1fx1KkYR+
ynyKurTScmsBbDWf119HJIP5gnRLDQstWg1uPQp3ThQ2QJvlDoAMvJU8smbeNfS/
msoFR9VTPakMEuV8I9X/FVZzS9+wtChiDCbcvMgB7EAjb2ZcSf8SQDb510Olcqlv
0PoPWmm1D3PFUNikzJAD254mJwVwlJx3BeeuEZ5RgMb+0cwKOrGOEPjJr5q7g3s9
vEGfJhWpN7fvnXnDLwus7bf9ivq6k0I5Mcmb8d/q9NBsKmdq/hATXe0A5GD7XcAV
N7z/rlr2Sd577w+Q2Qd+Bq6S9Ad7/GAv0vajHyEw7Dg6JXHibh5gQoBsR2FcZynK
XUf/JJJaUo41VB7/DNf4+Z4PIoZTDLwi4li2ArH/6l7DxW78dl5FIFX1I6hmeTbV
O+BfTBnwnfw0BMs4mxmw2sspVBCB89mU1LmnPN++06oMI2gv30KiGKNR3TOTV0hb
M60Jqcvufi7CPBkQKyoysIcDDxJWPP0TlOv1t7nRTW8tZYcT/EmAH1smYQrtXybt
30U5FJVnTCOy9bY/acEONhHkg9dDjqGvb3SYbiKPPRnweXCy7KZrpwMzYRJ6QQKb
8JVnCSPhGVb2rRuoMqT7w+qSu8Iy9fSponiYblfy+SHpT3M6DXxVGrBk6mGJtX/6
NpYS62haWmDLQDhMw1cuV8+0/1TDhhVofditzSijAlSOT85DhkqEoJcuETHs4s8X
jtwIP++o/fj+7UszjavOMr5LtXMHtjkK18df6WTYhU2tCjZssPR5vYyegVAbi7ez
6CpqF3U3oEAKjrtBgNlb8cjCgnE50uboKRUPGZXS+a0/QyTor5jdN9rRVPmp6zPJ
P1jrT+BtuxcvmBSSREBzpYNv2h5Wxa5U7dEb83lQ2yI9fxDMUQcuFVlDJB5mXSv4
BBB/VAtGDdfIRYqnAebkdm0k41pPNMLLFPwFs45YVbkk6Zd2TWjBBh9kTD7yPWCO
dmOHt3sKFHH2DvhWNJy40j2YG6SpzpB3CmKWwXhuFmi68M6zvMkIKB8hkcaEs8Gx
qZdS3s8BBsBKr7qWLNm+maXN1PtT/538kYLBM1DdnJU0vynj2C6KwuaFdBIzYFAe
3RP+J3i5iVaXPcpFZYcTOeDazG+hwNQ3sOeOs5YLYGMj4pUnk6OD+bOSdhRtLBm3
YWf1RGQ/FRifmozhiIxPEBtDSNkfmPtAMveGyK/1A998YL1LiGgO7y+yrZBEcLLn
gryCIdbreIhMtB3t8aPt5LbZ09xIS5tH40Ak2EeBekLRj9PNAwPv0mPBfA1HEsSC
K3jNsp1umq0o8JVcEBIeSiTjv91N3kthJtbSbkiez9ROOpZ1AeP9gSYIN6WT9YkD
N4B+slOvbLClW2rZh0rmomPUlfVbvT1pWnq3i+qmGITSiKy/ihhjvIqSTsgmA0ff
xx3oOgu0MB0bWifgouIwRMR2hU+pOPmOwsJL1ahbFy6I28WqaRnO6oepU/ZNh+/B
prkUrrY47miEjzeKczqa13WYFXozHO90tY6V6oLT2oeYwrU+WJgSpaRVMVG+q21L
2R1Pn6/yKb62n0HeOd3Y4+DVTPhw6OjY72ZHC5Zwdv5E6rkh8nDXrfFYChQsRlTk
QKCrq7V6+xj5L/rhPRr7CWLIM4g+2uyh22fXdpJO51tmB7+55xLcfNRpg+zMugcZ
Zh7n1gjsd7qt4xvBa81oGIAkOxjx3eace9ygl1RjSycwptNuD4U/8Y6lFRX3wBTy
L3ExtpYcTMzw3zXT3PNqH4tA9ZHo43Y0j22pkvH+QZaHQlLbpIxQL+n1MX8dAkkL
+htxF3XJvA3c1XRKI6jbGgMP/X5oWcADbgtBBB/gjFn5AWH0ZsI8jXoZkZnGPOVV
JLs/NfJLGEt/ZYMBW7qaGmnoaKLMG+abMvOmR0Jn4d/RVCTZbKRFgj83jjOfekhk
rBHW7BZ2NYvtJ4nLY2wAf7UpiRPy0EygdqceD064trZHENI28YPbW7l6QJR1FDzH
hK3DwWCi8bGFfi/0AQ9XFIQRbCMQb0s+sR7CCVAZK96GriGHArHY1L2zpgM5gaOl
PdO1SiLadTx56fhUHTwi+H+qXDqdr/kcwLDUqBAG2KVL9TCFjoZSElb30FGluVIo
mZLGHfB1d3hL2To6h9rTb/S1l2iFuirUeDrsGK+QJg0XDtpsWNuK8Ent5o/3WLka
t2mtfRa38+oYolL7QSre7nfNPSZIgijw3w1qA4yZuwGIrN+rjue9RHe5+R8tXnfH
8JNX+p5JmtGAL5e2EiX93tLl6j/JAOBKBY04TrytMfd/05B/KZepk40wnaHsnCPF
5x4JGhJLocnJDBkYjN2nf17w06IhPm0QEq/wm4gjRhzCtl9ish8RS0pWpNgSBhWW
Io+bIPh9Ysi0cmYxVXhuCplTPew4JLCw52hOo2HA4kre2Bc7+7y4gawxq9N4aU3U
UjqA/SE/8dj3OEQACukERRAsRB3KK/WK6JHGbpbzysTymaocjdS9D0jyI1+V7ubV
WVwaJ4tEuiSoPX/sY3EXokHadH0TptwzM7heiz9dXBayhc66zkl0NlFjKP4yteM4
+BsW5R19UEVSZXuipf9bzKbNb8+j6zJCI8Xo30YP4yVp/A/Obd8kFqanH434ejHN
2dE3dC1nvp4pA9A0hSMgc7iOmbTWmDYXh2QPcVOqUc9Is/l78aHmq9VRUIHT4Fds
fFVz+se3yr/spzH+kobHRIFIFZkeiKaxFU1GV/PmBfXEIfmOdmjO5WuKLXIEpZrZ
RCU+h5j5nvtPw7c9itaGrg2l3o0uGlOL5i+FxBKvlaiC26qBEobLBTbEy3d/DR6Z
qanEk1Q4xTf/gyuyimn1RDy608Ml73RVLe/7Ea2TZVsmf1NzEJU7OrvFCKdkGkKz
PrB5MMwo/y5Rn5FUDmALg9SeYBZtkCcaM80GmqPFmhxJpOGsGZyWyvbIHyhtod57
E2IZ/yhYEi4r5stx0YUpF6KZlhTfyf1gagO5t1Jt0aE+/+E0DkMqud0pHyIb6Jfv
+V8wgvIbbVzjCSwNZ5AHp8c5Tp2NTf7mHqOvAQ8z1KRWnwIzmliM4lxqKiBWapQI
SMesNVVjWBjt3xDcnXXABFDJx6PecPCDIco/KapH+Kzwu8W9WQOrFzLPj8Nb4wJ0
vQUbLis+aKJrVZ97gXU6GcYKYO8qkDIDbNa5+J1XD1dVwAATlWYbUfUOffycnuG3
WHkpEIifpOIgVxee9CrP4Lo4tX6VcUw16+iPSj8IQeF3kzGY4QwQIRBP87G+jE8y
JrK5ol1oPzcWezJAFDVL+fIQRLm2njzY1EL1s3JGySpkCSxbZ0GVt6IGlw+O04RY
eoFtBJEhx3r7p5qVr8O7NlrtkbdfTnHHQEi4PvV2HRCbMibwxxovWoBDUOyb571S
QtwbHVyqSlpsbpiq+atY7JVuvKYca2fEmoGvCmoiS2W+lg3uz+N3VV+6S/8BCbRD
ZQ3DBfnfr/YBVTTmd9FXJ+cwj5xpxnEplcLl5eMRVLZmmqDDAONMitetgNzl8YfL
a3A4YiFiazeCgOFo4lYvYATw/KarWC7JYES5gb6G6kLPxT1EPFbp+GWyOCxz+Dzb
22LbCZAKmUGR+oAuY6RbE+PffRw20jAFCZx9FofOm2fD14yg1X6IkY3gzLKZSvMH
m8WDz4PeGArcIe0BY0CEXvnAYoEI1RBGEEmB5eBd2EaqdE/gn3MseCsVCy3sW0sK
0Lq+HTpaaPm2/ozGWU5t4HsKy8Wnqkory/4GbAklfxOI4htaNfoPql9ZH6XFf/hf
EFFU3mlpZjHYisX01puNp3WqzoJiaGyY2LOGlBH5DV5QmQO0umMmIhOI3PUyqWxL
/VLKow0cuYmemojUVrEvCLAR/Enq1rsnGnIKGQ63JemvbSEppxJ19vCigdCKaeVx
UCWTyoXrgmINXww+SFhwY6PbO81eKIXClY4Y0LqJKQJ+dU4GLk0v2uVy1dl52lCX
/Ub4pBwugIv9myeKVZkyPPrtssH8y4W7p1cZ0dSFwq3VNvrisOv1EZJefy9niiuQ
/IV/cpPAUqKBD7LB71qK8R37rAolGkjH7qSBYedVRTswzu6Zwm79mfvgfGk1ecD+
pDIwTC8n2TLxiRaVxQAbtD/Iyu/P2k7X5glr2SFOvpRi5gC9OiGjosO0BSm0G3qh
45uHfNdTIQIErA25Fv87JAiHJFc8rymNUEVUKBojQQsEWtZ++HBPUlX1bACUkiW+
frlfhnwCwENGn49Xe1EEQfFoRiVsXaJ6qsgKBSHV/twIly6EuXLPJCnwxVry6A60
SJatum5Vjap7UccNj22MYDGTUh05PhLwkq3brcPsgpK7LCVXB7ZONZaL+9TnUj1F
uBHC8kNEXVmdIk9IfcC1iDafLCTjpT/q3tLnlDDKDK0W1qYkRN6rR1GUpbLc0vaD
iaxc6bdWhumZIGmxj0ru25mpHgfWGrwI5IZ/NM7nD0E55mke+BpHpIw+TMskNbBL
mizWLNkvIat88fzUSW/7xeQ9+gmx8pb1koQA0GS9UjfSM5f01Kht4vrlq7GiDEaW
wNvbMKHZs9SyJkqA6U2ZV7jMq5iqkf/+xkrnjyWbJ/H+izel0QBK3rmQbSBB2sML
DPM6qdeo83m/i48yRM0xHbasY34qZgPXU6vigNWCHQMDim9AIYsvZyJKb8lGUn64
YsaNG42FWrIkUakJWhf+RNWFmQ28f4M05mDpkFMukw+j9Df6RkoDeIQAxrndQE0a
Gjb2pvLRBjjuTZH6Pn9gA3F9s2zB//YVNJRoTvRtjCo4Z2WshiUcZ3KS3vBqAzTD
f71ssAfS/Roox8htQ4M9Fjtn0AiXpbTZCu0zV5CeLc434tSU+ZIusQ/7eiKGDJF2
KYTPh9emkZIpmLNN6mx63iqs2g0sBdxVw96hm/uu2SdcidvEAN4iVe/Pzutp8maP
ssx+4Aihhgtue9yTf9JLnQpfOQoer+NYR5LAhAgGwOeaJVa5Jw1hlSr0mUd3mynZ
WC4X6AefUhwtqR/jlnn2nrbXvDsVde0Fu+c8dv3lu+JtfRPDidQ+J1sSDOSNzEXq
FXYi01x59p4LdS/K6ZwRynfAmBFOiNKI2FEF7xir1ZsJlg2GYF8pkAWwJry8M9zu
SMuLFePKJrCCIUnIGcwoA9E/QfvDW4mpKTAILVYT4LqEvvT2Mocen4VQEWZDpJIR
Afl3/9Cawk3yvSsi19ur+ObelgmHfuK+EkhS+57yRz9FcMrIr8aORFmwPZpu6hfI
R51xETcdL92y05Z7UHu7AMF8HDZhqfPnjwn+UUGdZ9O9xmxAHY5DPqMZMnUGrw1J
NtSX2wn/OCe7CFeLX2BMCF9hwOWCg7cHL1N75eEDXWumvekd41/Dfg6BbceVFHwV
PDOfELYeeWdssLLpr/S/i8cPc0kolB1JBtCdgZSIi6fq0F1lETJ0nWkYNbfsT6DF
H51tmJvUYpN/Onae75Qv0iyN83yk8oR2ZJMCkWPKfdKP1oi2+gOsqale03j982wr
tRD4n1dGG2d4nCSb5ReCyKbDPm4KT1iufK2z2/APWPuYVXGCa13B4BgRCTtL+Joc
MmL0XDEz47MNCza0VunCGH4RQEUbZMgDAS0s0FsKXnjmsE8EYkF0dupp3GbgfFl2
ynOI8OgcgUAckH5QWA3GbQpW56dXC/ftocBti9UN58Kfjn2Nq/0Qtx159Lv5NSgS
/AR+1mTIl1YQhE2FCK7HcBRl6EUrldW4kB+jdi4mpt56+d8NIuQaha2sglwILhVh
2PdDSV7SzDE/TxGO1UOjwdJombmbhPNXejUSVFMt6yoMy3UiPKF44feeZHM+pyAw
KyGNol8JOv0MCwl522ZgK9Lnh9pkb4nAdzS4dDeiw7pU7uPjsBo9yAfnx5lDtmCG
mZdzqJugQ2PUzyo9hzp+xOnJFIrnDbHR+x/QVh9rl2tMF6DmIbiY0gGtY7hW11Ab
dnr6hfzn2cT4WUJCzYRPbIHAXAm21cXq/EK9Y7/Mz36YEA1dIMOZI+XECdg+wVo4
NYuuI5hcuBIhAu9SQ/NusGMyxXFEXL4997Gf7IVydknBKSYV8G+7Q9Rq4wuivCvH
c6cOhmVLoMMSRw16SM0xmM/01JcYf9VdUj+ZQXfo2WEkdSrUYbVip5EWOpeFuU7L
+h4eu8bDnKnr9TwqW9qk5rmWlQ4r1WR9sTLCt1WGbaTedbKB+Bno5bL1KHKGM1uU
/KarS4CzeL9TztvkpjuVn6aCrM28sWCM1mOOLiKAwNbLJ7BIZRxUOcGiMIJMO7MA
ily/gii/DzAgiLEo3i38E2NqHPhT1kP6XE1dZEX/xURdbhzySy5dS/sJBzHlP3nc
2P122KBMUTMPJB1HCFTCG/RZY96v51/g1rGbifLVBVyI8I/vGirf6nmL6Wzsiqih
gc/9fjS7+cWiZFUsPlXttYPsHtgLkPimrGCOTizDPe5++ZMtKPmnuykTMVI7ilO9
x6qx5vBwFOEIuKi7dRPLqocUVaOr+fYc6/TdSfk6sr83gmRBS7mL0cWX1k5rXSyo
NngrE5dqRENFfFxYGfoAlJGGjEuj1evDcJ7XDFmtgAYNhAUXNI3bZq8A52+Ctvyo
IiPRzxReSuj+xAQzofFFY/XEZ/NLicwHJ+GwMvX4iojHgiOGMM1Q+kopWIO7ht4A
vRNBedUknQ04Fe4Yg6jYGKJFRKxkmty+6MXxjCSZVvI9ZI23SyGKvm5jH6bZQhc8
/TpUC7BVcODpFjRaPjuSZTLhQryDGFBjEswlD7xLrjoh4JsKZTTotdEzniDYdIrs
ervbcyMdW9wmVgfiMO00ainCq99hW55GMJcsL1OjlmDUsqae8ahxNC5z+9qXrAK5
EACk6UE2UC3ElKBstR9w1upH8Yc4H2Smv0ixYftbQoXKufSspqhEeAGQLmlpr76U
cejBOQFldS3zkhTHGU1pgoULzLBZdP3w3gX14zmi9CnP9XuSNyQkSGnpnKA+BBDv
nq0vDQBw6zW3g/f6K3Tx2+4huathmhAEMrVMwcqt00PB9I2o7tc8XiIC517I33wz
Umj1CrIbeMM3Dq7zRTNWA2WtcPTFTXTO0/Rlxv3vOHZCZRy4HTw/A87Asmf9jpe3
Jl5ftXsh+fR7vNErXrnUj1T4xDBkb1ciu4PXpZhOb2WNcP+GgYCepiWSu7I8vLb4
ci+s1QoufllSuTNDBN23D0AlFj8riM4BYRlit20ymYBS9xBd9n1cvmuvaE9C9zqR
3D/PBd5DK6aKa8D5aYPZOUljV1M8Xt5fh+jyjcOy7Ml/YMYKw6ayz0IlgNKtuqPj
A4Om7s5J+OGoRUUTBm5BgBiDYkEEw0uhISvn+OkKWBqYDG1NZssSyUx6nacZtIut
uZNUXBldgzc8xkvBH9/07MH1djWns/cpuhkJIllIgDKVfSgrQqOns20XxKQxsFcH
t6vIJU88nO9Q8sHK71EZe1jRNHm+tFFqpiPeZB2Z+NX/g38zT9nThfDdr1V9L/Ae
8D5Fg/tCWnF7a2suhcy4WplA27gBY/aFBo+NkcV+tLoJ0ZKJ2FXJWEAfBQ6utI8B
tKvKtR7TLnMHpKX87mgwSfY1c5HG5kcL+mKVb8O3XxyLP5yqNjY7mNcY0R6tmNgs
b0ST6ybfKXsxlBg0nNtw5YYloppPkZddEI9zTds1z2/7ffV46sWyNeCehjjWl7O8
UrCKybntKFlVl71q303G7/G5MghNzVMNWwzC+2uvuBKC9hruSshnDW5EcXv+h3nu
qLuam+6OwNJt2yP6P7Tscu2X0kHtBPq/Vjv1GrXr2s+kcMVKshHeoEFo5l8cKWEE
S4UjRYpCwiUrDYBMhLOZT2VfDorpNeJS4G07P/7GrryapoY3ss5a60e+RMjwMPyV
pTQikT7gDRbkqPmrD4n3qfI32LuyOFOY02iJzK8K8VDIwCzojLlLjLPn32d+a3lR
r1Z4QbqYwUKqfW84PLiwtfUtHtfVzcG/qQWHZarYma3TXG6G08dtAKdGI+nMZ9ud
Y+Aaj+G+enXOm5Ifx9b/eojV6tWQiJ6lYLSKqNmijCHggl72t84o+HtPFna8i0lk
u9V8PEAOsAaOFKavIx6KrbmPujUFE9w5JGaF8aEd6QZD78uDaLjSV7w/cyiXPpjS
KFYrnno8BTWJiU9iPorTjEgRkO7GHSTN99gj8Y+R0uoqOF4IAnUiKcOnXzuzYR+d
VgqnsySIc9A7iouUM9w8oil1smkPsUcfZzh5elbCHLPvFLy0x85XpyeNvrjIEGCo
OIuF//3OdDj6WWBxC28YSA2WjcZMfdorfYTEbPmeoPq3fbly7OYeN71kmN4JgffF
GRo9pbz3HXw50YKiyy0+JLCWei2+cUlWQAHn9qb7/5TIBTu/R245aMwvBmhwElS5
2Fl8xLidLHzu+KYombej7uJO9giIMX9mdNJ34jQF8kSZ9ixCrJ1S8nK9SEflOYSL
YjE/pMZADm9vnvf0pU83fHP3kwlIHUKffr35kA9/ZFyOVLxX3Pg8mSfHJmmJ8LqA
vAOWwDAtg0EhbsLRIUFFDeJz9wXHtaX/oBysIitvg6VjsIdX1837usiYLtz8Kxaw
HKE5w4DAXEZczuZneP8YSMa0eax6JRhnhiypF4W3BRncp6W4UKKgttiexkzKcDGw
F0tKoTYTYWo0I+kG7GKX9Fq9i6/KnO0Wwtcaqbq2NWaGuc1+caU/9aG9VI+xGoUN
K8sA2WhHgTO0u1MRLqHffbCN+/tzL/vAEaJYQ5igWyKlwb9IFhTh4iaSqRNOjQNq
sztfNQmreaUPthHQNTzb8VLyzBicMpIU8EHnxtkZNLppfg9yMdo0uFTrXGxtzc8w
LUxwSPtnD1sQpgCJ/9Lz1FOX8Rl2leB/LClLdZSI4foeSClLpNa44hWjDIA+AvaH
uZ4dFv0QLC0LCzPDTrqEhMvjYkMTAys5veE9I03yhTenFiTjwfz7tshtZo6yt6Ct
pq8zOmvQTZYyTq1weY6Vj2URy4KP3XqugXQ1tRfsCcZoWCbniwxqRGwDCtGIi2lg
lQq38VMzL1N2Lotl7x+fJDAUAcf+5Tox1ZHqsMgDENJaye/Rbfp78ICQUS6Uic3N
WbhfAAsw1z4siQ4ZmbdwOk+c4PZm36j6cecxCTihZl2Zay/fVhxaCSWxe7xhP/hf
X2me1UHHmfCoQ6Y51GzYpeM0yJytVWbNMjU11CEuTzzi9LQisyAZorBbEM7Y2dnU
I6ot07Ro0VqajezsRdu455/zyB9tHmbahRqiOLSDVs4QqI3xA5EjJOZeECNmzPFr
RBf8uc/IhomZr+UrqhY5vyFl+USrrxGSZJZuc7bUHIbxdAREsLqRRRi0FYMUPzHu
6CkAu23GyFb6ycakidJQmpkd+lEQrMgU0ht/EBgLv71SiZirLq0UUjjIj1AX9Psg
a///85HqizbqtUSwY4quTm2jO5p/0lnIr+m1yA9OGEPUmXeJkc0AqnZ23T6/G6IA
VUctw0h3Z3y1RH5CAh6L8iDPVKcQ8cKAOEqlbmJjbLayoFvCVLlWEFsn/7Fz14YZ
UZLRqFBimwViIng7uS0BRXysgY64p1kuxK6+7vLGSbgvbZITwy/cBmJbdQLQVKP1
XPnxuVZ7sw8Yma8xC5F1dHu0+CGbk4j0fzzf0OOdoe7YSwDTVC1vo+uKs/a6eubg
XbqM47Bw+3HBtZ7/dhg946wANzBopHMeYe6nXSXbWp+WBsmmvLyuqYxpoaMSO570
EsPedCeNftJSxRKctNZMbLivKkAOW5nVl39nuWZnHFU9D4H4ei3MZ6/H4DRdzOU4
i7s4VcqVBBFhKWU/KpoDrvWDkd6hKr1tDZyKf8Y6CwLQfC315yE0MWcw3hInavlC
WX+vdP3cfLr1pR3ODhSXNk3FkQowJRgLNJSLY2bqRbdAMEFbuVsqZMa7eI0yAH/l
VYRITfdW/Asx6U8l6CHTtR4iarac//GherO21RIAxbqZIo7JXU5LqjxBMXLat2ib
FRTnYZtSurrLOS4+d0dLnmyeKYFCXWnJmxvss50Gu+dRdo019FHydXS0g5Xvt+vC
d8DDnIWqWdagyt5MgXI0eZGb0N6GkhpA80Sf0VkYI0mrnQpe/373NPzgaAj/aYqS
ONiGazqD8YqPCCY1IikCFtsZWBcr7MtIebA3LhxLyGMzI2/c94DmZ/4HDX4plKvL
37xmmkOCIz9wEa+oYjclsazDVuKGoPx/COrIOCNbea7FeuTnq9Ai/KsELe/Sti1m
dqWgh/XP5KIjvabISL/v7HnYPRzTJyHMbxKqg1cH2RpxzRrSuahbTj9lr84hs74A
fAS3ElPRMyJRAvGXEUuv19UmO4NNit41itcSuNRmG0I9wFolhQacveZb3ATwfkyD
HKQaqMSlT3jwuWTpZHUlrFLgassXzXq9rRrQy5ql9r9QG4q9cpXbh/d3CgNyUz0I
Q33u/UFnlTgKynJjzNtdlQMTHMCiOAl1HktMa3bbtU9PObd+FszCgu2dQRVQpyaj
dfZzSC/3TiZfS52POiVkMtD6ise2BuCApHTFOdnoVA3G4UkJdDxV7p1QdyvrkIuR
ezpu3qplrJnSJBZyyJG48qaBeAmhjbhcUcYKci/EOS8J4wqx0hu6kqiMrczUfJJz
K3d5pXjjME3S6uGD1s3DemKNkAIOAG3ZI3Zg1FnUHMYbqqBXMj0nxNNkgsP/Ra5k
MNNcY/qXbiOUmyxGremfxsbmEVzIG5iEQPFNYh1cBqMme2ML5kSnKPPPD/RZi9Op
HWk72OQrQP7s3T3s/IYOdcZJMyOmU5M0oGNlgNPDwgCKu66Z3eel+yclOfIv3CrC
fwXU4JYl/FzVCH7puQPl2M+0izIXRHhMQvXxG5UwXIHZJH7t8dkQcVpMrftnoruX
lIJTSPQ4hHVl8C53pBXkgVfByF00v3CD8Kjaevuk3qNelEewu1M8jMBt/zqGjHrq
YOfYzt9Z8l4a4w75HH4G1e1FpiqWi8De93VmaUMtbM0ISsg5eE3aIgLU/Lh5URFV
5/1LVr7IZ4KsCf+4tsa8MDnkG9zrKA4V6wrc6M/tC3P6TpHlxrcSnXqDAHbcW6+o
cZg1fkLqNnefGeu8ncPT9FlUETWuhoorbJKSNgpqAj3hNpI8NB5dlOrx1joKOaHg
1lI7obPBvrIfIZZHzf5RvMr7OMIXWc7rBUoK9OV3BwrASPyb00/ntFDNVpxtjZsu
l6M4q5zp6GKmxMOwGb7Owvm5nl4mLZX89mp9EZuvEL9B8mv0YKlliQmQfC6uIPqX
kV1pkAyLNYVQQZUktZ/gQfvTFG6OPlwwkuDupGPWargPgQKVlqmLijmskiwxieSg
ovo3YKC8f5uiMZ7x3QEjzN2j0pNBLKFTwX2Zym5kDXgwqgZIvVQl9KxyGVjb1+qC
xPq6iAMjzDHBA8TgRTTEVmsc+ENu4XNfZS8azsT7AteRGwy/RMYVYW4uvYf5kybw
z8W1bqh8CexoBWoTaeRBX4kF9KnXWYctnAZNRIK9C5znF/V4x7XLvnWLI4gBDmM6
S81dOX1waz9elzsUHuq1BEq33yH1ot4/fldRJqPjsyJ5XKR6Y8IdXHwrDkOk9af+
xiE+jRunWkAXyfc4EzsI5pqaA+teJRgwlge2wLZK/zxa0jRXaEwyGyAxPVX628XJ
Uxy4DAaFnRWnlg63E/l+pa3ue+Ji45JT3mimh/p3zyLFeg7t4doohYz0Whc7nxYA
D9833AR3CAgKqh2LhUvIjyeSDXLZ8+QmcID1ZcScIJBKRHgMtDT+AHDO/pFL/QUj
I0rcLlaTEEZg3N6R5d/NoQYMb7n9M1pwXv72xdq5tofKYXWp/RcBcAJHmDputO0a
RFN2pyRkU6lY/Foz8MOcj774X/wlB/3JNSbOI91Bh2jyfmJ6hGbMdPXdhV7k7MB8
5k6IekKEpilIKwhKhN23MZHsDS64J1MFGgqCrjyyczDO0/wAvd95irMcUYTfGStz
7PFhWQ8j7Q1uOyxHpCSps7Pf2I0v89cRaAZu6g0fM3vC6PBulQkwew4/CfsQl6zH
cnczepNWyWCSW8LZ9oZqqoGHZm44gpZcebT5gQlHZQACevx0IqjJ2UM9I61+Ok13
8lZKx1ROGoJXnIzkX6hZ6M3ltXsW3y1SGFocJdYjEUL0MlVCDX2JmdgRmTBrBU/C
ZGdFs7bXanOI/4AmJeeh5J4n/MjZ36Nskauk0qp3bd1PbqxuedfB1QpwdKlU4zMV
oWQHek+HSXIooyG1I5NrUj6wZwDNIbVkP4qtZj6SprGjYWi3iXjrfiUFYSUNfGdS
T5IL4YUoRJunBEULO5PfFRNuJpCG2hgd69WcsZ+6uDGmgNiSPc4N1wY7kep2KCGx
G5guPtWaBGBF0FKEGx9xCxsoLJ3Jl3LkgR4hs5PGnBQMuPuCVLcTLyyjoMi9BXCv
aQEIq8oCcYWrRQOyjcDZOapgRlrlYL7JUs5omgo4/y+JTTQ6lPO8Z1HDxWBAkWI7
xyLli+5nek9PUzjGGg9TNZlrf6J43LVgWszKAjrWQEL2Gdt9vNIcZ3v/Q/mVxphx
nftt/afQkTuowo5RtHoipp+6jSKZJrapqokfV657IStiA3Y/y4bWmBAEi6PmLwjq
D+DHWGyFK67atg7DgrYDWTQpoPGom1TOHQQcDKKg9oKftoaPaUgPiJSo2YWfqCb2
EfLwTV3OkHBPB6X/dRU4YdrwH9ueXJ/wBhtFnxl7pICm2BaoXZ1yJ18f7avKNLK2
Zl4nKxXJPFJ3SAlPufV2ouQ25MRe0mlVCORAJqpIRpdVOdns63nUT0LAHNJvP10A
sbYyom/KC9jEtWVS2GM+M+kk+ka2p9W9lpY6/snLHi5N/o/8plP3H7ieY1gToyED
GBxtoR1/5ncj2N/FvGgI1yNoQ5/SMoKna/+ZnQhHX/Wf1W13kkz7fVJVM4SHGeRq
xl7Dc4Hay0SkcuQQJWSAZE2woBUAQ3lpIi2BakfHS1Ysh4vpDcMNnN2LwiL7Fo+h
A8Q41AuJs3JUdYEaTnBtwyF4yumxJglXI00l8XmJit1l7WNGi7ViKIF5awraUglj
EQIW7zW8C82GDdIS6LHfHbIDb/fMjM+QdQvIb4ezbGPlilTGV1IkSaXwL0qTJSuU
LkvYBzBtZL8AEYtueDhnnyfArZ1RbRXefn9ihyxoN5ha0E9yJFfECruFZlguzwGc
3iLPnNIEiBCjcOBRedWs0nemzQieedli/Y6HS38396D1JQ1yXv+4ONI9sHcDSF31
j/HNhDNujGVI+SRB746gBxz9ZnflA2/gB8sHwB9zxn+0rpJZtZoljrGZcisvJbc7
KnslrpkyY33ruhq4Gb1eya/YUbhVuQZ+MHG9XZ1GaUhywCcPMQp0wYhkPoT9Ifbq
Z9lBEp0mqFASvYZKLO5L89gTb1OsUwBelGbBGZ6BXgrbit6UE8PBqZYlyABfuNsL
uWCiKElT/mydAFrfyzVUoooOAG0audB+ntp4Z1g+IszwaFBpKVL59Ni2F4QFwnn/
x695ZtYDaN/ucsxuJFkhZQDuYK7lp4tFvmkMI0Vz+pqT+AB89UZSITimJbkN3Bl6
KZMe29cr3cU7argcPHU18739AAfhaS8P1u2vBUKBWDmEpeTgOoOdASjw7ZGyeetO
Y21OobIcLSiW71wkznY3ozT29YlgmMbwA//MSSMStB5n0zeT/Txt58dTnI34VRa9
x0jDOakO4wyc6Cf9JTiSsezaP4cjz16zuvr7j/fVZRsJzaLiarrY2osV0EOPWBmr
5cnJEKQIUA6fYbF69e73mftwDk+wA2X5IWfFWQj56wfKAXvtIWohZkwOp2Wisi0m
e0/FX0ubTBZ+E6aysSaul168Nq/WPg8owjnIVzKoGeEtPV0WWaqZPH+uvMYt9+c/
p3ra5iJmxaiqKO27UKOfn2zbnUv6llr8nAaI8cdJsRQcBdWtBw1TFpp+1e0ooEzn
QAUp4Lzv29f6MMv+U2WWZ6QMV4hzJcP4ZocVsFQ7P/lLoVKV7FO/KEvkxA6UQVss
TLL1PHbj/zuU3pbOTJR+eWjtc5JxWhE/4/xg52AYEoHO7hiUylkD1K6ptZc0Z00c
KX+PkSjKXqnWXWaP6sZpDWvQ0/PonGzIQ8q9Kxlwnwb671IXGhA/FqLJpCbDhsa7
69S7MhvUBj4fZOZc4WY/FLatI0YJUb/5Np4hsW9TwKhDmJtN6LRW6Peww/PjRFwO
AhMquo1F3zHYoKqiCW3VgUlbDl2OwZbkpqBQoAkdGWo2ecvMfRKFgW/xyAnE4Q2o
FaaYnmMfkvmGk08dnt9mcEFyyEWMblRryM/tLsLlK1iPR+Bh5bJnGekfOKNcptN8
MibFsQZU/BRjwS0IiTPl/vC2JW5kP3JNog+Lg2BCZiWVyncYRh3Le+lcgo+IcVMI
Nd+lZtWTIFzglFayOAVk8ydozGH8mRT696H/Y4NrgHrRi9PEA0z7oX8WCpshuDCw
ibHHKeaUPs5fSigDaR3KSf3mBq955J2qzfaw579gOxJCVW9Un0Yn47vQvfF6XwkJ
7+UUxJBNw1R0CDoxvFGBv2iwXlYoPbHmn2aYYAEUmQehLMIrdbdPS2nq3SqJDwG0
fem+n7u2QJv79gtzap28CN1IAwbFXKMwddM4j8WQ5g6Z62nqgFGnEtCDhnqHW75l
vYd+dNSPWew+W1OALAjgckvfDSjg9yx+M1E/d1zDfUnjL9Qiv+ECvn+lSR0vZDjz
u/BM/r/Th4PySnaBLtQlA39HzSvAnzDnKhUFsebAGsLaRCg5/ynHxev4+wVVpWfo
wyFGIjVCn0JkEMjBE/xZFW9rLNEOKPESyfyf/YhkNqth49LoWtzeZNZ1TvYQZ9rB
fNF6+fbRTv+znZ0gr+fdysLZ22JEOfW6UIdNM8Tk9V8DjA3/dpSocSIiDVHIopSV
+CbgtJS2oSjwELS8EyL4/LEOhYyp8Ih+SQEMA4+SWYUf5auw2ONa4OaZW63Nwdy/
dtrdJzZ2nZlJiyKXUxilWW2AH1gatoDPNxX2n9VBvW4xgHzR5UiT/czSTTu20T1c
EYYkBA3DNfq23tpsee/tDb+Y3dYvBmNtIaWyv2P+orPehcC6O6nRuIx+cdnJiC4I
iEpZWMz9AFV0wz8xxxch/52s8ppwUOqqyGBFH60JpxKePh22+gKJQcKJTU/C/IMy
qUdln6TRVVI/SzDpV0oNX0ngSScY+3fsbIkhCbJeGiQD9Wz1KPKGyqLGelhlguRw
Jk3sTMoTb+cvKJTGC1xoD8sMnyyVfyziVCUnn8dXPkiQxzCeaII8GgpXmzHjcIZL
ZIPpchY9uximdZllxWqvYl0Qljx9ZiSCO9KNtc77d6visb/lCn/+uoiwe+QR8HOi
FF5jNIffS+1xXmFncXFImHSBA4YQedxETfLPFX7xwCMEqTrKcnhh7Y5yvnpgEXVL
xz3vlOjF3nMQ6xqI4LUeKl6j4UIjzfFKInOean1O9IFrdMcZwDVTpEtgL3onpmH1
BCzGuiL/UgqwgxWV5nMi+mAPJYNBhCg1Fs2U4Psy3Msu6jmvoA664iuhf089enP1
uVFbAS2s380tY/jKu7pESRzmvImbk+clIdFpo1T344mDgcZnaPLCcDA1TuNjp9Mt
HpzkMkBrkqoAXFeKxVnmSD9EL57yGzZ0M892tk3dRGaaFhqlxbAqCS59mqmtOjJG
t8pHm6kz+JSA2d3VBNKUVeDBV6HxuGOB3Sp/qK214kvBpEQPumxRlXsdJWNxLZrq
Yo/JHfCKc3k9xWnkYx+U+DhluUWri/knZL9VL0aZWWRy3q0Wyv534zTDRFtNDDB+
cI/bNPnNROGuVz/HvzDxsZZ9HjEHlIJR4EQzxVgrOuoquNJ61xr7+U1wT1kXFhLw
IEBncgwDj9dGsuvtuA7MQiAziw2Z+WkkKoBuv6tS3JghYzoW0S+fTytHCNEjDPPU
c2DVk4xJCOYFa092Ex34RxKRcMN1UcQFMoF6j8oG3QSZUUqaoRfudCrDi3nazkws
0qsoZxtlTJvpREjP+sTTu6dbm7BER4ppXGuJKmP8vx0n3WF8QZtBfyADTEPI2qIt
zGXwXX/zDJ51/qVAKeGbt3tV0uFGhQdetm3m5HaxaFUSqej1LpHjjLkvlL2lYbNa
Qm2tv4AdQ9ovWLg1COmFjiUdMIo3jrHI1t2cqBpezNXv5slUDhZ/Z5d4TyPEJ2bl
X5tb5WP2/j1QeTQbALpEMucJZ9FJ0ow45E/BMwmMrH6kHZotmkAnAv9EUtLVG27w
FuG/3e0haWSDroXvG8Jjh1pR/9DZypUzBSDSHLjgUwMRmgOhld6+tgRdTx+jb7Wm
LFKuSTAhCHtkTpYjygALGhVGJi7MwXsL54HEsW5NoV2VPl+Ex1ZVOpIqW3OwwIEu
Dex/BsNSTIJD+OLw9ksJ6x8r6dRcfxqnXsew3BqVPk4Ua+N3k2fQAx8A4jcu2CYD
2H6GVJIVqyhnI+N19Ic5fkZcSNXnxFJuFuVqTWoO4YnLdh2BQxaN224ZbcCV85iI
uQ29Z6tH/IYHcWEfhqQvN6VMGMd0R4r4nKbUZ7YUxMBcStSLNMw1MW5VMo+9ZZBo
T9fECNc+Azi3c+VMJTJKBmmBfTucV46d+sHvYmRDqsLc2et61sD9oZ5Ya5xv5rfo
nW6dAUHZwvtgI9X7HaRumA/OoAhx2QqaaqRtLUpZZ41h2DT4pudTrn2ZEov8qxlI
uB6UjxbyjWENewmN52DhmD/aU52lbYMu3yCs0unOv5i8tnZcH6SYRCtuaQZl43Zj
rZOIuKnpWuyCDqFiuebBvwQTvquxNtWnEa5IWHlA7srHOdzY1G2XWJhz6Gg2aI1Q
wPQj2a5GCq5F0vNIEYMzzrzXXsSE2feLuFtdko7Yc99/EBNdefEfcCKNDmgi6WlO
osHnDtnZttIMEPAc1Su3KYEvLnfk1Llu+Ys0+4tW2iR29u3IhoqKcfZBv16JUNV2
M4UlsHSR+SDJq4gLljbgJZMJFWzJJ+PP8yx+SmI3AdHEbQCb6hfo21VmrT09eYp0
MIBqcXTKn+YacCtK/2nBC+EeKar4sR+D+b7dRT3/jri4/sFUyrHhC/Q/cF9Iau2/
vG4maUPmU94UNA2P9kJp3DCXS7bPSeETLYdebcnbyTFbNaJ8rl5k8SZSbAF53zIR
2OM4chNluvC+CVui4ApykuL1r3BepeBQ8aVEztPfmrf+fJIAPdmDYU+7Q42GacLB
PMAbz6P78F3OwhyK7S/fnKej04p5NSgKyAqQ17m4FbEZL4C8iNJTY1BA+Bi2JxW3
e+MlNk6KJL5Z/gclHnzmVtx5iRatqFY4jM7Yh3Jb6gpYWhIdxIXAd83atUG/fTTI
CPObG1u5gqBwzLj48c+Cca6PQGc/QxhRSRtDeM4P8X0+lEIaUHWqjv8IJq7geC/j
EzML2bAabr2/oYXa45pdbmUOYMibH47vFfUL9pEhyIMWr/OD/z1YWFyPfyh2KSVl
KV6JbdU2emWcAPtoLxc3Jq6CH0L9qg+WQdy0/RevW0kEpqlvoMT4lavS14KVWp9m
HeEbVNiryOLlp+A7jRvLKNoFZdeSVADJUykEDWNYHJ0bEg8UAdKLfmKaoDDL9GnS
aBrS5F4UiJznrC4BI14YdRzG2sEbnnj56KXGP5Enk48exQSNWtq5vS6QqGUbdQeL
NuYWMnuOX1Fiv0LDvg/f/so4HQHGR9aNBSGWfGwwx33iAzTXDIwj5PisyYt03/cX
pd599kJFmxFXll0/4NgCF3T/rw3Ca7yFbcvR+/S4fWzRyWVQAKHnwrrO4Di+EAfo
TVre98vKnf1yoQ3S5mq3Rb315gXXPdIgWzbiDW+BNy0nL6LPzKQTcarm/MHL39SH
RimBzfKdrNBGKxmf1/b65BD83BcexYUc1qvTFJm21ul5bGuSAyAk9AU9tbkoFtOn
aAoToFI1AIMeBCkA+W97lSC3ya3t4gyANnRVK9s1INrBhr5KiYoNPQpYc/s2ktWs
8bg8Ct4FzoII6Tkmcv1G+/HOLNRuRBUQBTje2DR8lfWM6cBptvS2mu72w+eqvdEH
ytX5qH3fHsKrf1sxabhkqYGtUW288xBFohYXtrgQ5+b/GiPBE/9pF0MdqWBDX7dC
VhOYqrhxLP1WkcCic7w6uYZAIESg8MNnai9SlwfVt4agD9yRGhvh9rSAutp1cmNK
+tXGdiGr9BwbMbAfpwU2DQpQ78TqfI6ssmwVAabdaVUvQ27ebeNpcKyoY0fgCSqk
HEWMiAGpIjlo7dhr9V9v57EuxQo5sohrHdpPctnaaPrr9G52P3DRW+zYDHxv/vQj
zHmC8XQ5gjV+JfbSyQZFHtGAFwMdZYlhwo0dkyRGoAUemtqwDCcnF+TFrL66iKLj
e2j+DXv2UDQyF67+fAfuH+HHKiT/gsdhph7CPh+P6g5fq6eGIqpPdyIl7CudtIEF
osdYb1TQOz1l/Qcjh9vwYIG9S8b4zksVqzvnSJg6R0ZO3V/7BytXi+eFY98KXMon
xyj5CxoRVheqfBxHky0M9cOuBrLhjEVLrhaC7OaAXv7HeBR7nRhQbQlwOo3P5ZR8
CRryDyZ/CM+ToT1zLzqf2KgTKOGyg8GhRhA9cMPnfpECh12GLz4oedsed+5W50UM
5eAmeVeoKlHJEtjycqHb/qsce+Y4o1VRxhAhz2hyO9oYrznig/MQQimW186ADWHf
As1Fj490FUqZ70gEPhQqYQ0Tj/JcTlFLI26Wx2QpDxH+sFb1dack2IAkzGOQP/1D
TKApWh4CV9/I9DfbkjD2sDK5S+wTkL+5YcSSkT8r2VOZsZVq/3OTcEsJF/rlC3Iv
oYkud+4kmdjnJ06ZHnP02gA7A2yUhaA4JIu7Xwmzq4RDYA3afjoiMpIGAz0DL+b1
2zRRs2OdoWj71rOVKvQB3ae+dCHfTsDO+0pS2iPANcTeLsCDOZOY5cnGcntply39
4J5FHtNdHlJPZCFPSkuZeVq8/XTXVNzCMuHHFS4+TL+pTx3tCMSpGiLyG4FtVrCv
cJwUCUq/FxO6giP7pvdMNa549+rV3eO8guJoMsRgUAje2+SE/r2KcPx+QvRityfu
0EghDReSRL7HPaPXB8wQ6O+hTLf/YpoSydHscNfVVKymHtEEdjX6GpckTzvVp6OX
mTxHiuRD4jzObxBuxc5VvYidVCddk8sR2EqgsQNj8QWjMGC7SRZhVH3dWjYy+2ru
ve2YE83Kb+Hn7uXx6OjyRkbkRsjiBGc9w/MeN5XVnM/SFt69ifwgstKoaGZLOArn
f411z9P/0Rr1d3AwzQKn/6vcEcyHT0GoiEmouQN3EoImxzypXhIyiijq/UmkzI1P
oKDTMyrIuoLVcEegvV471o2Ay11DjkKDiwD7aeJamcdCIbXt1stRxKygn290dNpy
ZcpAuOKH5SFMCzzrjJNE2VNSoF7YSiA7vFOx8KFW8yjm+Yj+rHCMxOeud/RDUQkG
CPSSnJ+j2aowkMEGHY8UGcbA//5yoO6SvfBS3PVIMq4OaBdfyjXb16inX3Yb/iVQ
HYHqP11BkUNBCb1JkCJUbaaYJ2njz75Rflpr5yKlWRpU9Ipqa8t7eGaQ7KhiDmes
X9EwCx3VJThh2Jdn4NUSi5f/8Zki1PK4DTKLiDJ+qPaHTEkOObkpuBmpvFCmkhF6
vsVWudWwWFvM0Qfxn0y+v2FzgT74rOANoL8hZXtxesarDUyoWfoM38yI40bEXxiY
Z+aw0FwGp/yoBlwuWaFRkn9RLhDmPwe1VqzKP7V6GGaHOKpjsn4W8y9sDYBj5YxU
9TajS091dEgEZSkcicGOwfRa3CBLKsME/clQP2Be7fJonqAn9SCrmVLUcoEHjo9s
mg7I6HyZUjqIld6PPgOD8rMy7+7wT05IAB2w4B38fR4NkTHtIGUVdNZOG3fun+zJ
xGNSGEqBYnTSwF9vXLzZoH8GA6LOF6C51tSDFlvEy9AadefSP1smceonshg0T2oD
k6q24efFB0R2lDL6Yh2jK/7EgsXmR5s+cpoWwxSBt/1rUi1ZmwvBv2Fgsc+0wv21
7Fy4o3/lsC/OobKCVpZIfY19RqUBUw/vUGsYKfKA85mf4fyrqAvdIkz9nR++zu3o
J/rxWXin9DVC2mzNMXSI9HGFGkyOzk6gJNtd4BsTuTPOMxCB0Gk9GHAvCc6DaG5r
9wlqhJ4SLyFdTwjWmUEd3tLqtLj/mqxRkp0yf2IBxXMjZ6kG33Ynyxvc+0pKlq1O
tJ3pLLph5aGOEt3pnUaZ8m1SHs7RRUFIHpgo40dmVwWcBmaaM8M1JM6w5c+p6x31
cwcA/LNbfJ5wM6jxlsXwnQq6lCnaVZc3hz7WUzHW7T1UR7jOUTwq6csxgxo5IkmK
f0HCAyvdYv0o9rHJpw+Vu/kb1SlpscxlZP1ltq7ma0UITV3ZN2amjD2DcyIZMIgM
UR6IS/K1vZlv6eTBzQKS2M3J4/txCvLzQazO+mGxXGyRHvT/A2pOpvUnwxXT+Eqo
iJzAuDrEG5bNytSxTZN9VuvircxODHKDJ4bKC7GyqGayjhKu0QbKNcNI0qAErTpq
xzEy/YNK3BjH7TzLSaRLXsKbX7g9hi9dJLG/t0wGdfitMQGQCmce2wyQobNRaqlR
Y9Vzq0OrnVLEuX+bjE6XhAirPf8srPu3S32oEsPo91JY0Xgn44vsryXQeteeVHlL
ckYxQcJ5iUYzDVBYpaoAhhZE0MGZSTW5AJ1FLJ0K2/XSxUNvZ2BGVSiyEcLTvsu5
hwONfT8TcgZFsOZpd9hvAUSKDSzlgMOHxAaBGYlUDjGcFgRKuhMD5ny7aKnOeVdh
yUobGg0gJU7SKdOtqFGhSqV+gNQAIFgUuVlukyir//9wvgu0n2iqIvrV9xQvbPYA
dTi7li6jgsnbg00HLpWrZequFHSHRitzbNEJGaO5AmA/W2VfE5S1C2Nnwbgi4MvU
5HDxwLmfiwpxeI7+M4pdZ1E5wxYacCX5kJsAQSfXFBop1loa78UFmqCFup0cpw91
JuD/kGGZh6b4iEHPbarWMAT/pscfZN4PtNQd6nNnAeOOpHlGhDt1puIykjEPXa0E
2z6F5XGxEN3DuURP8DSqkAycwtAigxL0mCsLsQWU5Vq/8Q17HD/KBjs50LJXDHI6
uHGefxtQQZGlsyssVwQoiWbbi97HilToxBEEM7qT8LT50x4AlF4bVN2i85ybD/kK
PslP5MUY3MCYPyeSw+5rIaYf8WPxCzux9ItBavgx+4wcfz+f/w748OP9Ls/GfpBD
qServvxOSNjnqc3RRGZ17TxowsBPcpAed+P6doJHg5abxh6VZR2A1LKy/5RCe4nZ
XYP43JlIvTOXod4BqjE7SnP27aMhw5zsgVNwZOA8kjDYicdUfN9vhRiPRLuyvtNZ
AvO5FB0+rYsdhcsdapyKAiGL2XPeq0qN9dZdhv4swtblFqAoo1tRJK++7faiMhnN
3mUBOFq9qnzToo+FXQp6zCxB76G1wi4QqNBQWBEgThDjw/WRhc2M2kZX0E3aPKYW
E02k8srFtEL6SScTmhlxkAiM023AEjYgTZFOvBOTGf3LMygB10YFj2bvqLN31tGQ
kT2ZYSF9wlZSpBXV+MZND0I/6uHCzQeU3Y3P/340gM8rfNVt39ZNXriUqgWMmgu5
/9R9eDAPL/qJN3ZoNJBijjsyRpQY3mha+3jC1oqw5/5xb4iI4pqiVdPlvlnMKW8T
th+2P09802VmgCKVriEaM1b2dwpwIjeQKDj+i6EkyOZ4m7mQHpDB753Sjo+JC+tW
NER0qvY3ullkKAPkdAmFIcRMXFXTSQcI99d8t08QJtFhf07dFSOgCPuxFeOgcfin
3Lm7qpRx6kA6xSFYQ5/b0tbJUU6nsxuIXJYHGnjP3swKfzBT1bjIBgoniJoIc2IY
DwJurh1mDBqcr4U+pVreGcZfEcQhtOVpNORAOyn4PuEUpi/Z+HU+tMl3kwkILkP3
GL3OshhE9ontV9AeaN/O9w9g+6A1dUaLCD/aXyxn2t6ZOtyHUiWB/fypuIAz5uKV
N+uCjFtWkxD6Vshv3b+m+cpUIn5fqyfT05i2x9igneBtbAGGXYv/8HnSZ1fFLB4y
OHBg1mhLLKeBcpEY1wcFX5oLKeG0jdri9SGF7BxrZca/otS+0AY11knZizVkT8kK
2eR2Dfqfviy0DjKFV1Kraikq/AFhyXuiqLvkSEwzfXmihaGQCwsX5OWOCPF3fJW4
DOIpajRAqXp6je5X9gsskHN2CWN8O9SD/RSDvIq+JLTL5xeSe0YKzyu4NnGFijIH
X8kL8DbI0G5MnOhc41mTKrWRhrHE2yMSv1Cn/3myxBWXQGbDZeviefVo2rjoaPFP
8sFt1dv7s8N5DpJ6ACgRg2Ikm5sZYI35wQti1Wlbc708Cq/Tgf1JObkGTgy0SNBy
2LTEvDlINd+FUniJb1kYmHlAkwKB8yBYcWp4zVMcO6jT5MS8hh0nULIEHge3Lu1+
jayVCodVr+vSkf+6g9jdUCH0zUvwvJDHQh7TsPjMUEYb8aI1b8mOp7/6334B53QO
Hs04YRiVKD5Gm/RXx26/2Cc0XpBMCl9imerw/zJcL4xEq3M/fKQNpMdVGNQGZuBq
BzmU5kJU0CxosgaLN6ZkWe18JokT3ss51hgDtFRYtMbM3dVVM/G4hDRQwcEWw1rI
HtAzpYXK1qiPqq+c0CUhl0YwvnOJC/WwUSjl1c7xvtbdkTYCG8+mc+Muh5bzTgts
GPz3Dk+5bi+FFgdLpaBIrjfzvA6ywz1lD5HGlg5fC21kYFLg+tewUGYU/8z6p4WK
Bsi0wTCqBoab4RY4yc3E1Hsdi7Hx4umkQDHGQjDYceEXu+qhoPsiRKTBgEZ8nH+w
G3ksLJygiOrTt4cqUnrQMpgMIXhMhNLVznP9899HbYk/Ksf54Cc0aC5EPv6RlVLR
FjKksvpyaEkn6WiWY1rviH+7AMWRiTla/Qj/gRNkmrwsa5KVWKsKfpqUPFVPMkR/
SeAUEnltmfJ+JjxkmPCcFxLE6NZQZ5CfOQyCtMddhwsht86Iq7KydLv4R0R0aU+J
D2ReYqWFYRtXTQ5WUEZX/OxiHtoTax/bbLCf2wMFOWmN4RXK+FlDh9mNhckOwCtJ
6pP10BSlbas6B/R84AI4zD5LCW89wBrf5YANRlquRMURQVHUZs8jDWmmxDGMIzDt
fPSSC05ErtYsYHkO7/AjZIPkQRC8gG8jrMJTdDXfqnGHDd+wfFrPkc/6Y1LVzh5E
RPz/W/PPtLVJU29sVUSjDoPwAZw4m2pge/Gk5wamjZ2OCojIY+Ymhy/DWH+gseBX
qtsMrjgV0gtjzhiplY+62IUHOk5hxn0nIzYaXOt0tNosx16cjNJ7bllOurZOYnCM
vPTkjjBMF+ofmgh0LWCY1Ag2r9EwHXoClc0ZzXjmPqQjOCHvykKspfyZYygpF2uy
lcL54H1vm8vqRi95MYnaltwaVr+FceIwHK3ytei9amQqakwOARW//loWYHWqxbaH
q5Q+HixpoZxbYaDzQrLg9/ya5Hl5atWpKY9jA7PB4Xaf5OaDKbUKkkem6xHDthqz
qFaz5ZKwaY4PjtrfYGO2JN2wDCMzui/uwM0+41bcI39i4kTnRzCd2FyFm/RKxdJK
cB4/7lR4Q6Ufx0V30VA9LZl7p+KIEAemeAnDyLRitW9eXEgvI90DVw6YHG+g8Z1a
V6gniUT3rH+ProOwWVARX9sZPmf552bmqm8y7EM6sU57fC+dKIY7vFeM4KzIBq79
1UnAHtN1lsugRNDoAJ+NV+oPa2XyQjrpNkV1XLxUhMhD7o3Q5CHeoI0zI7cIOzA6
W+niCWyqnJX30qeSUiG1dYMgRP88aXQHVk5zwKEJCNLbRl2XwYbiWLEhCxovtqIX
VSh+GyEbvFM/t74NpaKi2UUT3vPFciYGFGCdN2Qv9MAqoWN23N5pAV1abxq97TK4
jpOE3yFJT8mgMAIfKXzsTCcKxnhk5zMiAXXErnvigC4BoX+eN9iYIKPPvZps2avE
dv0O2shtkE8deoA6WM4Lk5vIYvWybwDPe/2RapuXn3D3N6p6R9dlx7K6Tx5e9hvw
IEpx5cyj7bzZJ6VqZxED0jD/H2FaubicfcmV0xM9INC1I1RevUZDu2ag/bIEQvOS
ZtwjIS9FNU/7Sr1bYCV203lbk1TzpX7gXhCBHpZ5QPbRi82Q9/stvH4kFckBmeTT
wtkrj1MBTLYvprnXGRpmRxOagZ4+TKxSw6vku1hL/SSVeYUfUnfupJ5kzwqgd1Qs
oTcu7h9oeqr5kINzS1AjKu1gCBCPJDIQfxtK6YnBUywXuNbFVcfuKVDxdn5cybAb
6HJRZd1ep4IZLyeOQSIXLgSCXHavlduIRQLo+dcTmlKwA3GIva1mbNMMTp/M3k3/
/5h24O8ZbRIXB1yj7TxlvUDSU5i4L/Mt/ZOwWP8NCRT3SBVgJ9RGhd2t60WMv7BN
EvIRtKI8qGOm2fkb/pwEvqdywmP5tKdiHkrb+21UFo5nySd2YaJnPXjM0209ya0P
E80cs726DT5+rGRPlifH3b9QPhU3J9dLvQbG6EDCmtE8tvKF0rTe9HiJehPIY1ue
Sjog6F3c8pPsUdYPd6a74JhHSs389PjPaazauqmePDEYhUbouRBtHI8os95aR8zM
HkVwm6n8CrAoUcRccltfsENcwpvO0L+8dN36THS8F5fcPrzj10gLSKAziVcpPuTj
x7ssUZYIcRfxZk/MZxRhHK+43OPxQGoG6ykK7mwA/xkZij2sPUXTjC7692wlzsaW
rY0RU8Gb4wRblk8XWx+o51gZba/34fBiqufKx97KC3e57kYknrK1n5Gf2uhRKgy4
rgqGb36BGSyay5Finq0t+O/nB3W8yHdzp1wenGGZ9cKElrYQA9vvbsHCby+AKvtk
RZFCWhyvgMLy7PqkjhK1apoTfVX+iJWnKnuR0OP8oNd5sAt+QU50Qu691jrnh2jK
XMmmyQfD9Mnh1YqQTW23bteUjnHSKJg3zU1QlBeqrlIv6LkYgwR1GqLRB6u6JAqW
gKhqDQ+2rccXPcmmJ7ZLsUJBJE1hX8GvW1uqdKrbq3Hcgp/KpTXm3BJ3Rv7iIoVp
oB8PJY5Iq+i8JEsymhlvS+o1Jl7nZIXJsZqxnek6DQY2eLq4azyPENdTcXiSKwUK
Q7StYjwiNFS3KcWjyWLPJyNPXSj+4G2MHd87ZrvdJPT4n+Yy0IzR/BnqWwRfs4+v
5EOTioEZ8kxY6Gi1/T68283DVhhiR0fb1XSn0iW8ljClh68y7JBbkgyAom+HUMVa
VJTnaDsUMF1xWRDfXKWeOtsB7SJjlp9dY5Z29Y25WadNiIq1uaqXT4PVKWE2NHHN
1dLhD6eN7B/YVDchFYdIoRt1AZEXd0pIvqmQDDJ129LFfivmOiZ3s53Jwu/qOvCV
VZaOnejUSTifYKrC9O0RRKwIpgK+I2y1lEzPC0gWXM1FzJLrt2MuEFT7gMGpHo8R
DfUNp5Bvf6FrJInpfhybh+BMvRE4e4NyQaotYyN0/sk/CWTYwrB20K6xql48GjmY
PELOhJczeU+vYRBQ9ZscrOBg1mooo32P/xy1xQRiHo64EiVYDuEoFaoGeU3B8k4X
RFsvl9Rssf8cSZHvKrbPMPAJ6eiGZm/ZTtwcKSE2b+Ph0g9POVAuCQJi7Mfemawb
P7ub6grySw2nCf/BgQkvCKEKtT5qY6SKmN7Bc1zZ/laqWBpL1/DTYtazaVFRmj3V
P/2rJIfL2IduM3opNBBG2VQQYwkAth+EWGkvCrNuj34Z82ShIXQffd85qDTocQKz
sP8sUvIKH0bJs6M34rI6N6iK2z5oPdVL/ZcDx5yxHhnxW1qarH0Ngax/jyfMAjYH
mgAWhHZVIowBu59wrr70MwS+LFRdukVBjOPW1fr0gTGr958VyUOISrae6WYatLN9
UiUUOyj9MUrlyb8pfEixGYEYtuhBc6xjwLFa2QPrn0sxfYGYLJqYoeHyKxvB8NA+
fM13b/HsAOZn0zxvcOWGVgp0vnh9tVrP9As51fVnvqU5wRzN2VzDdOQDNDj1mbQH
QLWB49mS7MfMIFFaH9PD3M+7i+rm8Nivf8XQoFtN8Ev32/xw1G30HaaLmBf+8n/a
KMc0K7t8PH1MGTMu+aCWnN/J53MZ9cbfJBEuCdmMb4PVGMI83DBkWXj/MIhhdpcF
2nJsv5GLTqGEd1STSvRsuWK3LrXg4ViOrY+KVbx84mCwv9wezKeXHxMODsUFQ6hF
42BMG3RQ/3cJxh0n/HK5cWkfO5OaO8NAnM/Inkedjg9Fqf4BQFsubX/5W5vryhAx
CSHzDh5fY8fz5dlgljqIU76bBWhibZ6yOsR3rTpCh/bTZeFbN0Ck1yNx340CuRfh
ehlO8BNmAoGrUvFI4G5x0yBT+KWwHi3Kw377yBNgHknBppRQik1iiWOSIpzoZtAp
PeHm7jATDO60LMlEHAmLWQCPHwkIjj1sxOnmg9Y5v1ogfQSDPxz3dbqN4fzonlOz
QY3bF20X9ELJaWPr3Q0q5MaB5ZdRHmE37fmqwtDdyJGbvMV7/tS0Pt5FEifsjU2U
JuYmIWCpG1zywCu6mExIXD0CG9SEdM+gg9BSX4zG7Y1c0A7sOegyEPuzks+UjYip
+8sWZQfqN0LxSvSH/wotd4UdqKF5pDOj8Q1fro6BOwLdsbaMyUT54XI3mLlhdwM/
4FjKqoukizviExE5IB5UPuC4FYcwpeHdwZfoH8JBSwN+t2wG4LoK7O2uykYE3M1d
W3/LvmJy/aQTLABjCo4LUaQuPTl3uTeQW/5CJ1EUZgriRD+i+ihuAALR4FCglzrG
s6y8iWBxxpgI1Cs2AY+sUgi+xr6H5yYKEH13RryckICpdDJheWLFclSuypG0fMOF
YUaeQoTrpw//qISPJSldc6jzof8lM/2K8xGzNKNp4PJgj82zQuO48obHNhabvfv7
lbzQaIYLx9nZq9vCNHVjw/MZdxFX2iSA9wKGypwgTmiaHom2YQQehDmHPCQXJ7tK
j09jw8y2a8J1qiEKG11jdYe9k6kuqHsvOYCH+d5MPU/C4wRk5foaBdFCWvjtS+hh
vT3CqvLJhUoIyTA412hsASdjK54sW06K3ey9wc3Sy8mGen58rd1xFHoG97luJ0Rq
mLS2McSRLqx+kwrAztbMr72qnccMYcAdpn6M3dQP2jAYFvRRswe8b2qUrEI7d6rR
gJ6Ozb7q1JwkmU7ev1ja+b8pMhna0Vm2UtWsf0Oq4b6roeHaN6Dywjqvu4eAdCXy
elkaScr9jqPIdLWm+oQcXdusynqw70c7NtjtgmDsnYJJBbZLh5BD7cyzENl/0h4l
hjpGXr5N2+z8NoQTM4rOrXxZnKBD3R6+m7zE2eh6vmto1IRCcmCO5gvJSdG+Snb8
hLYocjQkKRCXlO3sLh/gZPU1diDOELiuDNQextu9umj5aHgIx+0e1B42mgk+Rn0c
svECpHUvKxV7UXpYZGAaiC9vMa3GvgVdslhNLHr7Lvih2evKzC3OBpOdGbmO3weJ
BBqdMW7h7Z+/Qqmnkjfibk8If0d6Tcy6Bejqf+Dy1OQxWOGrzvztWBnN4ctE/V1u
nv/cnE0WVCdlnfileAs10UA0JOxsvxnsrPQj7WFM8fGx0VO08WKw82GeEZAiCp8J
lpsmYZgGWrvd+BwxP0dP4rxLEdH3wrMgIDtugA/44Kf2FSM0NiXRaGg+p5sgldyx
WvemwTEPZlWSm7xPZcj3+LTi0hu08ojIBdWM0yq6CEbdWWE5kgLts0Zuc3dILnd2
HmggBGJCco9jZIJ8lH/Jt3Jkw+hO+Lq3GgZcpNjSkCP2ksyGI7/2knkCAMt3FjHq
5WmuFbI4bMx0LhN7gXIDQJaWEzRRgC8qHuQLTlXRt7gBdmpxxi/UxhHlVB1gxmGk
eGCpn5P6E7BRV45Sl5dGaaloclu5CFD9Bh1Y5JZ8hBSYUcsX2TBj7EPjt+OBLple
OloLOx7uv4J+RYydPi5UdjxDNRzls1mnTZySW9now00szb2LCxo2UWz37qVzFixR
kOFCrh6yBZ/C2z1kKU+rcZfhJ6yoOp2IN+1tyB9jEWf2qhvQMFwl9fLHgG0gRI8E
qev9uqAXi45ntSjdc+Bq5gZJKCQWpW11mlpBD8zxk4Ugxdp5Kyte9EwE9a8X10bq
8FlT3f6Pcu57SNY1KXsktWy0wcrOn5fRzWHgxvZlqapYvBkkaPBQt3LX86BUSdyX
0I0Zmf9ZEryyIYHyxo3WbbkvSc5eJQBdc2QfZxGlxiV49fS2U6TodX+ZaCQuGu9I
6kV/S7M4o5RTbyu7mhiHYtZFtiO1qeYdjJgXCusvigLd9CxKhp/4EWO6b31t4B9z
l9bpGGYY0CGn5CFnJyd63eIGKUHNwSWOQ+h42EZUBpgO9FYL6vW4wXX+xPhamW0t
ZrvvY8ZinRJVtGKiNjBhLpkvJmRlehPJfNTxLVomlmOR5yddaT3t+9WGTciVZ/CH
Vzb9c+2iC/knoJMpitufDURiwCTPgKRIfKUU0jhWBg+l79VH/2xPv8+l7uE/US7T
c6WoLJrQbWr1xPCELWMudpXsIDOPHr3vBoTHOuvURed9ejGTyQp066PbsoLI2RHS
psNshvSXJoHLPRIwqsGczBYX8TW2gXbuK4L6IqPTMbKfVFe6BDbckGEjkZr4eJNZ
Uj+FKZEsyUIsWquopHxMaTl1HaIXP+47BmCQv92qZn8iBFZoA3/h0BqJ5gpViAY7
bhLfsyoLPJ8dU8elNujHduqlpvfLBxNUM1eLIn9QRmT0B+VWebr9aousPe3/VVCG
EKvpoaSv4MmhkTr4/JH6s/LBaqQpN8avB+SLW4MQg0ohfTezeyFY7rLOFLdhD6WG
ZpvbrAePfjhkvcJByUvrMsXkCQz0HhXbshlGVQphf7k5QGSaA0tZqEWHogxQeBHT
6fH0mEF35TUEnr67HZ9v1ZWhzWs1RLRBz25HgcdU9pVP/H/JyOvs24/uoBbYdzKE
elNnQ0FtsbHc8v74ysuIwZBTgKvxY+b+F/WYdq8YzdKWisgXnNSYe3k+d26Av1B3
77LSPED0z0mU/nUT0Xn0x4+tWDCtCk+jKCAXtUfqMo8bO4G7kfKPLfKEBNBBC6a5
Za6HqqVbgAqA3HUT+slhD7d0S4ivRoSGvHvWUg1x+0yeph/2nKI6GMQGo6yS5fEA
vtzNZa0F77p4+PGngeZ9WbkFrAlVR7PhQVe266CvjCanZD5/coFT1llGBcwL3MtH
YtK0KQrQ6vBonhgXVr10iiOMCoR4dMzQIUt5F6zBqa5jGgDSPvVmeHrPFxE5/scb
P74DE+Rq3IKtXzU3Ub5ofMgrUOyvMKMElAR9ildUOsyV3i3BXm+M5IV6m5OAlZtb
ug1GrwVcU0Rym7YvoatnzX8tUffqq0sV1Es/XqkWLigdqPXDNWA4f4su92HatW+S
0IOZ+gQMNYm3+Hq6+8VCUsFUzbxOpHP89S7ORavOsnFpb4Rgvgudh0gt5LlKbB6J
4MjR5U10WkUl6yoZ1k7kapXBN4+aLEhCurVjoJrbntyWJLhmsdskIqWgmtPYSmkY
Qm5IfUTmPRdsN+jnbJp04yWYguDtnwrhOCGqxj89qucj9Yhe5SbMOnoi4DvGBvPn
45tmC8W8S7D7apLMHDDg1d78X5pT0lTowkEZF9uR3AkKpg4kSCLwpZZeYE7mlmqg
tKSlv/JzpaNO4UbTpr20U2M3g1RX0XZdbK5hFOPksZC+vxJikmYeVx9MPgiVVOfe
jDgECOR/Y3Ux4On/pK/n15UhDvkekNdnug1eHOFDRI0T1tA+OqVsWa+sTHYDfDZg
DKYQN1dFSGRmbTXtDzESYBoJM+XpM5TrC+Oj8dBsP5hOZ6EVX0/IBfh+nynPB94b
i6XoePuaZUSQwrNKxT3LQ+ADOzFSlyjE+audQ4F00RMGPn3hZW5pLuLDrma9T9gD
BngwdiMLLK7SHHEsUfx6397S9rBRxma4aJKY2y21d13G5f05IcrjIB+sugAKGWvk
sONU+0kZBUViqS3B7Ojt3dCCkG7zKiiHAi5j51EH+xNGclsKBxjV81K40pC4k7pf
9cgBtK58RgVHI31ndFSlghyrwqBSRTvQIyjSA3xEXyY5K0xJ9ocl0wCmyhwtua7P
sbIURo01cEttF3UoWYa+UXpZMeg8aygH8+/H7sP4SXM4un2HJYAm8XuOYwbU4pf7
ceKLPTuPxqh2/qSiAoS43t/n2hCW/bGPStjmO8PYXAEybeaf2Xy066XnweVqmzkM
QZC7fqT9Nvfqf5GswGISo/SAEq717qSx9Ohe3HreADClrzwL7lzIvTdU7n+mORXF
nNQxBTK/KClt7z+mzGmjfNutQmLvc3lV2DsuXQ1XaE/y5/G/wd0luFrmM2teQif2
RTdroRCb7qVGQ3VRHrBENfUby6lTNmWbQpTHvgG+s8o2d+O2SFpPVZuyJupSIcDF
UdWpwRncouyjPF86Et5NMy2itYqqyX+UTxqtwRkrlWH5VQCtIfC+Ff6b82fqEdpa
gQ7z0bAMQidjMCRB7JGEpWFD23iO2K9itcHRaWRK2odbdz+8010jQfEqvKTGGoo6
0swjT3tQd6FcojG0kv0lQwRULMN3J0jM0x6xerNCY2yZdJ1J21v3R3qZE/ztU3op
7Ln2DN+5Dlhrz2LtWGjysqE3cJEzhWmQiKxxdq8MQNkiKcGufYNjRCI1P6Xhhoak
hKHKAJlgAROtIP0Rg7QcGqDTfmB7fZmHgKvrEWlmTYhjb8dW7drdptOMcY0N0HHA
xOIV6yvxrFiixYPNP7eLIoGMvG1w5TegMrujXWZbb94gvQFT7lwo/bfuq89oVD9N
hp7hzSGMRhFU8KNgxLSUVhnxOzJA+jyGKxtumBeKcS/3yR5nrb32qlwWyui9Q4i0
wy5yo22NGTW7HHpKcS4cWNxbhE2ef8BP3RnNSe2g2QV767tjhNcCXC4bIthrivSc
JehpDrpSfd75iUgYbST6bu1iOVRqmtUylbT5UL01K4tnS3cmmlhrm+tpCD7wkvCd
JfVUAQh8JqZIpm0D6zKMIAA3af2/kbwGtulho6s7Ws5AVuYxHhufZO64xJA9Zksl
gOzCn34lM2e/A3W8MtMR0fggelAYJTOc1hfqdri0QC54NF69F6DV+/Lv0Tl2u3ww
8dnCJGNFR76hvb9kNoX8mCIPInMHG0iJ9oPONr5vg29CDg8FQ9292GNq5AKOSRe6
PiDoxRqoceaSE49W0E4Ev1/p+qTazBfTwOrGH5t7jKALqKUc3lWi+zc1JnG9W6tQ
DqfKwrpaIiKE1mzzXnClnoS1yeBumlCE/BLTErLbmd5WV46vZsOAmTE6wNqMjBiD
VoT20exn8fPyNMBOOQu3Y8kPjA8Kh/PSmvy2bIQ7E5znOUwQ55qW7Mqijud/o5Lm
IiqtJRehojiv7X3OTjsOzBYSE9ktubiWeLiFuAsI2bXFckZISoWe5XvLSXDvUUkQ
TOdpyvZKlK2NegUlo4OpW/Ns57qgnrJnZ3ulE0GDqguS5WlSTr3udgspx6ZuTg6o
8XBoVRqXaOtgTUl4cXFu5vgIAgs0ifByUkNr4ehKJ/PEJ17b0Tjb21pNwLTh/Sic
ctNMzDA5PVQX7tZ/ZKhapo20ioAjxBdMfYgI/eAJU/YdIDLb32i6lkSTmMjXYhQI
rHk0IZrNa/ZGCAZXkwkja/Mf4H8pNvwSSbnmksE+aA9SB5vEEjQAe9U/2TxttBTE
lf6TkoRqN4O/C1ycDSw1ThVZglrNdsqWYjt+5XpXsPhZJYZevw1VpPp5d71uYFyk
vUpTZ8YQYcS8r1bjbd7WvCJsetepghmtcVSsDZf3IIagr4hcIgcqy2WhKYe/nbke
MOadu1cl4MhwfKqj4nDXirjGcK0yn9swq0qTBmEWPxF1/ihFaRgCz1WNY3ujItIv
ttTjzLP32ryVPNzWCswjlynqQ5CxMDM8BTiY2EDUASmA4h+Cf9LwE2I4TT8KnIqh
reNg5v42Tg+V5Cf0+n5ri1vNGBletC1vJsUe1YIVjyuDeappOjyWwc2A4zQ3Ovc3
FHVS7qAphAcjyOe+Azlf+TXWcmOLT2wfzpZjlFr77IcleL2D9gCN8VuDnTq5E6Nw
kAY+3+lAjnRVg9Xz2HKeBPjCQq+tw8UvEBbPEZf0ATyfwdgi4xtjVFao7R3ZqQ0r
XhWVIqSheNKg1lfecOGB1KrEQZ4CRLc2nacM7zsk9hmUCFEvGSQvRhm1W/XhwPX/
VKMrteUD6PyUNPO9UY8tATw15+/UD/EPFwhy8yRrSEzCrJV18LCPiRTssWVBYwtc
IhHklKBxuirFjcYBJVb2E+qiMuPKmIjI3y4TAQauWyfYAvUvG6Ct1RTYX2YdBMUl
1TfopzfDOe1EOeU1n62Atgx/DOjpHFYW26jOcXDItKxOVNvESvsz4g5l2EuN9mZD
56FF7bHwEkEgp2oOLz+lQ51a3YcHd49ZxTh/IbvoogtWOZps0ilL81sAUz+YOlzs
xNQw7sYLO2qUTkOdvyFwx8m8t+aFOt1cENmsRGLTKp7B5W0hPj5rUG76YnZ/HqYy
3xRlw9y21F9AG0JUoxYGV+9BlADDBedEqzXwVZDB0Vh5Sx+ReZIAP9cxyshm7zgP
+cGgzkXsWZ8cNOJ6uDB3SPPtqLMI8U4CH7/hU3yPUVmZa+b7T937nbvB/Lx6wKbf
WWZnp0HAsmBfyFMH++Uq7JL6ZG3kHUBTR2JyTmbSTqdiYKM9G8745PRQUc20/AHB
qzx9pke7GhjhSBEUAWYvqvF0Kv3RHKRGoXqR1ZabERKlTnDxh7vP7e/WHKH7cQWI
sqUsjg3UJhChh6paXTers8DiLZu+Q08y/e73b3HxonTdD8RxmglPVmg5thmvTvYT
kl0pDvZi9emO8SauJvkrXct4+n0iUB1Ym85TEtdUI1toxRn+BlnaoMnn1xR1IvB+
Zxk5cLGFGgjg0M7ikNaBwGX7FaLRITtxRrDBHV7Gnjt9I79TrunMUQDhB9k+tK34
pYsIdY8UvD2uB9W5/zEa/OXZVUPvrwAnEpfphF3CoJjJWczjcd51RdU1tzzq10qD
Jgh8/isfkH8MsnQcRGpJeOUKPxncm3J1WslQX15qF8hYDd9CkCBF+2BiJWdVximj
wPoNwVgnfkje+fRliXV6Hb6aJTE9/ZLf3GMZ2a79vGiC7gO4B6LKtBj81fLHOdJa
hirHcGeeEYr+m6SmfQiuWwCcigYREpsogmgJBesqp6vCHRHbkQ3Yfv7t/H0+hVhd
EdqXzuJjaAi1Gaemh0DarZYlNbIvs9Y1uY4gVRC+KsJlLp/ns0sgyPGWh9mU114l
6SEyhCEfgoAI2fo7kXcTsqHikbSG7GBiAlsYZnsj8hHhaxCrzYqEEnU9j2eV8ekr
Flyj7W7g5DFQvg8Z4Ki7A5wcBpBi5tqAlqefK+KQu5l92iW2ZVVmufpd5hW5GtNS
RGYeW5N7xbt/hPhke6qUAMu+gDapYAWCHYlgvBueGfun7HNdMNH8almepu7QxDTN
/LiWP22IDl7xU0F90sC6WUNH1iXIg2PqYMSgXPUZc2y6Qd+5l7JO28mys8aVr5Bs
NcnybUZxdP8yAlKK/5UrCPpOwMy7s9tvhRveJjTYn6s/PIfhj0z7zCHpWrT5/ue0
xl4CtiFNCbu1UZa5IIF2/hncRh9stzkQhjNpsya9s1wTu0gAwmUuQqToWuhqyz05
sGBvr1uAUrRtpQe7MGX887yp/eC8sU2OKsmG9G6J2klyjR0V3WPYaPjqL1jgfqh/
QCrGgwPSIJ9KcLTjUBm0I2MxQL+/8Es3BRj/GRi7o/6OY3TEpgZiRp+v4Trwbbaa
Rlxbp2J34y2gYk9oHPgVdy+XpkjVDJmu6t1Hms2eueM9K8UICe52ty4arqvbPCtt
JQkl6W4s9zPuNNTZdIgUYP75b0xwuhNqbZlsaYnzan7qURl241MGxEaI3KvnGg+p
qTAHWseF+U9dn+Vig42FLLCihHv/j46szqtrqwb0dTNZRS9PhEmc1IGDz7p/og7w
bqYP5jB6GlpG0j2Qt7dZoJl4GLXZLzyADxjVT1afT6XgHZLyziuL49ubA6mXyqNL
weHVa+xXFe0TNmYA6eOezLVXX1fMmMBP0RbdsK2AYGn/3mBCRuFwfZuLuVOCLE6G
RstbW0jKNgviEggwVGsBUoopWR6GgNyk3qjxsENj+snzMhGUQOB7ohH7rRD+p+iR
KtkYUuA1hCO2Bg8elRrszE2vaEV3hqVYWFaLaeEJBQWOr0JxXahHcX6NmNw4GY/P
eojGvYeGKN6nZkkQkIAdrEllvLFqOOfesEX6NiCdoynrz8oXAi+o4WE+YWCGazcj
P6kg0UWKU6OGjKoAMHKTt3Ri93WqNNWO0lTg7KZaTlYi6MpOYkfnvqJDxZl0DYMp
Mg/kfh7B8cw+cl+EAXenMT7owlUPlv2nxidsaEauwGTqqGeK0szWqEQVVewRkKZQ
zJxsNAaxJZB7loBVkLRYTFDUH7ADlqSxneBctkwaHYjJ74OBBDeE1Mh+Wd9FX6/Y
USm3fgw5Sa1C6Xf1tfQ6qEodYKnEL9t998qT8d9bOPoGO7I8rLPBlxCf031Hi3Kk
JGhg6XI0TwTgWcRLfDEE1Wd5i89FLVLJmbJEIrpTyvJ+H81ErEaHRaLG56vlFa12
tbirABhw75HRZrDyUhkJ3yGGMQW2KbhccC6OfMBa6RMHr96TMAdIwFmaDAvP9jJr
jrXtGCpYSVbu5kRL3pQ8yWIeNVY3EKowceQryKyP7f+KmUFlm5adI3Uh1Nhnv45s
49iwTjNQTvHDvvVLGJVY1BfleCc7a7QGvVuLREWHRJXOgvHknbvy4SfYH8yeiFrX
zpVvjvdvwuMhvQ0kMEepVRibQCU3r3nRoS4hmOc6xZUIvYEe6neAld1e6riTuVbw
uqYNRE73oTYdeo8Dh029Mo/F5ONeXop1gdFh0yX0pX7NakhwIbC6eUQFWlAF/J/s
5w3x8XSV0bEAqfOTQbvXjaoExy2y+BwvlLdXOyo6SvgBqbvCBHYmvoyq/F13jz9Q
d0+H5B0P5avzvZoYh2t4925X/FLtkRrtQ+pfNrjXmAAgM1ZVtn9KFl3aQRN3h1tZ
zHu35zaJ1qvvBbGrFQnQ9ZMmmTuQ5dATFidhXHZbSCBh+gYj0WjslrEZB9+jJl3t
Q0+tfEKJP5EtvgCYxIhtXueclr436/xLfazwX/yq/Y6/oBOAt9jD5effO0BFqztg
zXl8QEcVw0+DkalEAyL3dH95cslH30XqTHwxWKNEkKx1dB9q5z5L8+Hb7+f6RoTB
FAj8TdXaJnmFht1feidhz0XNSgj7Jbks/gjwjDKh7MVL3NdxoHshEA+cvh+JAJfy
FKsmvEo+9yvDR2LQm27DSbf5TRPAEEEXGlBMzSy/dkyV/Dsh4+YlzwS7pkwZrE5+
HB8VbKSxtAJt7GPVKE/endb+F/tQA3rAsv1+waLrrkS5x9aNECFRC6wDQL215tf7
zwh7tc74R+vFYYKG345Jbhw5R9Ds5mqY7vUAciGfXOaStw3Y4LPRLgXNftz0MRMd
qdfXioFCWYp3vwJ98M7WLSL0Kiqx2aNBvqH7Lp3fctw1pUVUsUI4iMvgfsKIR5uK
/HSzfQzAoeXlD5Tzb38eeCEWcGHJz8wD6gCCkBAoqT06E3PIMkKT8YYMvojzSExQ
P3hAE5TqzC+77rrCVMNIOffD4Y4v62L6RcwAee1QhNz70KpZoSqYXGlWmrAZ0nDx
0B3Dx8S1FJ2KG7RPuYxDNwg+TNaEdhAj13hYx65hu+aIWsCoaTSjWVYqGL2dxrtj
37+P9UZ99TZAnPbvadqSsmWhvGVcixMhSGwnoE3LHR35NN7271qxynV7YkytHI6+
pxGl55iGlrzHbihcsw/mSGHWMZ3Ew+LMP5nPqoBN0yaD8R2u7stwb1TmwCONkrHe
LgGcUJYHyZWLjwtjRwZ7/CbU/G2ikfT3ykyawiGSDdvr5DJjF21aU4b4oihulHw5
bYu5Z0Z23ELAg4+2QvuAud6sXZMSM/XBr8/m7n2cTpzZKaXA+YtAJH4NCCs2kcKh
PRU8kE7ifsz2vZVjLOAPmPgn6kWNeoAcyVwjI41nfH9RN81EHTKy5UzmSeUwKpRb
0N3fPq2J48Fkn/m0OVhr48qLyx+DhWuAoE5FDKdnQLSoR6Qg8ss/5YQ6AoGGiYp4
OkDs7YnLdsyTEd97x8n9nFN2GOlhqX49BNBsbBLnEF2X1E34vC+rCDdEgB7lGh5c
ga6ejK9ozKpTE5E4N73JoFwGsdO1Gn9h43fY0HlxNBYkbg7ZCZdk3+y54RRH0nfy
Bf21dHAyX/+hHm6U0EsO8ptJ+PaKYLkIEas5pQFycvGKAcnjzMHEhWQ3kWyxyjZV
ywkLD1J7m2o4yTjxmHY2yvs9scTONbOzpELoUdCiXmfACTImRMO2JdnlmDLN2Mrt
tyac9WZKE7Ybu08/EMmfed6WnV+OLFOhEbNVWRFNw2ycv+4yTbu3sYony1fxnhN8
ZEFfKvQOE0WUEudX2Mq40RgzbR/n6wYD0TVz21xPtaFxw7w8YyZCBIRN7YdbBu3E
M0qjb5M6IwNWPz9xj6K/wv7Ols0j8sgaZ3Rxtbdz3+XrMqiEhlWD5xZ5mSXL1RxC
X4RHCNuuO55IGETOlaQ/jvYRD9UOBd2ZXu5szFjjB/P68cnG6//UicBy8OCGip7Y
CLc+9MIzKxz2s8e6h+HBa+Ebbr3WVCxAft7hnDHT8l/HXo+DOd/2rD8XOy+glHRo
1ZWf1fu/D3G9/1z2h2tx++oybRpi3EpQIPKmTwN0gH+o+Q4QYg3bbgExPLwJlheI
hu1HDsGntlVkIzgvoDDhFrjITBy7/wQ0TUI4Zyv1XAFcirYPCUWO3t7+mTGsfm85
t6E65ZJ7CE6423Ds+f0addWB7Q4epnKcVYCBC7vEa1DG6F77/mZnEeGXpxDgCex8
Y7DWUGF/bXkolOaf1KKVIk5a6QwSeYSooiO+8JS2KFwDhSr0Ur/2UL0JCXhIuf8o
sfdaPMFzgJ299La8BXZPMI4NSlrnwCS+G2dmxiSzr0EsPgmooGojNACR8IlDkhBj
npjJzdohpgcX9YqEUP23c5R9wb0YzIEZtuaV+O5FrANInjzm6zeDyoenCVLfytwd
TzYeCXrwDdM77lTBItBxndx2SLGpQ48TWKneGjuzYxcfChFoouE1Q6d3bmukg0o7
GKLmawpBlOYTTU+4gKIDhI7Cwv7uX6WGGu5pDBlrEZql949g0annM0g9nKRSgj1p
+XzvEXbYdDGeHVfAMArVEH/im1lrHpmQ+q5ifbWfA3wbJ0t5XsMoU1UyJVtRt/hk
8kLMs+NxjBPkdvhSMbXGzpTII3URdPumyFeArswcpDiJyTXNLlXkxFOR6f+CwdEH
XzkpenidzqsrJsDhyt78cSWiLhQ7GAwRz/vNhjR3WvDXXkYPjF1kAmWXp3LqaoVV
R/n5lC+SkQ2JY4LniU6tSfN4bIOHotDejlavWOc7VjEM7GV/XJ2K7NGoYt562XCI
kIAa8JAhkhzhqAFB4BWKMKJMMKEZYrg5BHHoiVpFl3NseJ02KjUQCq9SrQwASrNU
ROaMfM4+CkYcy1/vLsUk5FNJxrLGxzTpEJkAAXMT4dko7J9vpXdK5fEuhPqTg9sn
lXv++hdvirSQ5xjdcTlTjSLgzNBgBRSqWCSrb//N/zCy9czt0i0lQRJY+wHbBAlS
d0IjyE1YYOh7RpZXxTCPbHknECM9Tolm5a4GGcdL9wM1aLA2tOzNBIkwA/Lan47c
yHfuO+34i6456iNznijyny+M1PEG02a1B4YA9yRiqb5WyAzuMddzO9eUKYDvXOsN
yRjs46DZWFsYc/CfMJX3ZHGOsdOLmV0ULV6rJ+6NqTbybpXjgHVWhYFGgEfeYyWQ
O2BJUSz0zT2VQDfOPD9K3sz9PZaeRTBeek+Q8XTL9Jm3xI+9JixqsdpFx+23eZOm
OGIp/TITiLciRSYeMJulkPFN9onqFFy0DrMXCU1a/jlos7nS5+EwT/hFf5La5FCm
AqbHu4xns89n87baALE6vc9hMYub3SSNEzVTFs3i+K5XrJgwJWZ9B8LhBbM+R6G/
+z6d1guuEpbEVA2IM6wQQwdsrjfDYk5W1BO4H73xo73Thmt82mWIUJJwDcPYOnkU
YC1VL0E4363IUrbpD6KFm3PB9oMxIWbC+REJ1cw0fT+gUzhBazPXvyI3hMj9XZCK
4XtAa2OMA62L2gHPqN35OIZlQ192WywamViYfAVDYM/S4dssCygidduC7WXKRVO5
u4Y8lcm+gyPMWUFDiNGq6NkNhLUB6SmdPfk/jZZnlGSS6/wjdNgC0FWYp4YKG6Fy
Fvoym6bpedf4e5w7tr8vv2LkhllpUZQJwYs/lmGoOjwHh5CDwtE2GY/FNUa/nSm1
IUrvbmQRJ4UwO9X+oPjqTDn69bB8Z2/m0rHkwhH0VXPwXvyjFhd3CusJR/P1Dn8z
WHmGEO9jQgOtp9G/3EgqZRBaFHPA4CI+SOkrXk38Mz8u6uDa/P5RLOQDuQ13Fs5E
+5+nJ4yFwswMN2Fhfla14oNnk6BhzCEFDEYM9SdmN7VA9bMC1Hn5qiF/O//EYxf/
XZkMdcmGNRuOuGuq8ThY61o/kCUvxZVoDeyrYVdUDKOu5ZqI7NtWwFBn+Km/Q7WN
DsyJ6P0atK8LFF09BPGiiXTYEZYq1GOi6YM4n+H67KsJvbrviO5st053ZBC3Ydro
ZJQktdGUxy+ln/D8/FsZm9tSjxpB7Km0cX1/3XehJooAFyumySPE2HF3doBRHais
sxB+eH/Pk2c8QnRWfi0Eebrq7m+l7TfhEFs88wOOi8SMLkbVenALwtF5ql9fWr7c
IPTX2dMH3F2D5eOc0DJ0qLC1gsDB2ZJhx/7gyk9k+OxXVUb7U2duajcVIyfkwuYE
Tt5WFs2isVjzxzLWHpCk1zzsttyU285uheMWL9wUglk9SZ27rFGBaJQoVVOhdQtu
FOgN5H4u4Y2WOOCMkjDTfnbUT0p2oImR15wDUXHl8aIjzFy9yuvUifnrxugcSWP7
tKFZa3BLuxZmef/4/cFq1ZYTMpmhKx8wCUtOTDMnsynIeARbB5cQZydYliOGdcTf
9xQ+qbcJt3BbwxZy3hBiYAM4nFv/IG9KB8svDKXoNgk/9NStRZNWG7oFPqP29oSx
KKfmr3VNzoBo+6vmXVfzHJVdbXypgVTjPYg7t+QVJOGl5ZlkNorA23XZSLlmFWIA
zYJEvisp4YUHlNLYwv27AVv/2W51FnDYVe9AbYLvruZg6w/CkwPqkFjZt6feVMuO
d92V4W2bLqRRbGqrYKD62/j0zDMb50WWpTXOqYlUCFaEKKWWQJMd6HxiCU6UNiyR
Lo75rW/OgD8qusWRg/SIyLVaek4vcszD47m0vE+PVtPN3XGuyDSK2i4q9MJJQXTi
vU+KzOP74yeaCOLR+NzGJPFUnqwVKzzJNvQmLPstJGwJZsCcq/oxhs3Js6STSETn
QwHi8ffjL2zL3V6SmdC3dfTpugsQJAYimeN2gvXy5Ed+T9/udJ5KyiWpWPc4Wynw
Kv4BTsOTn3eq4/aX021JVTev18oTa+ZHlnUlqQCg0or6OmMSdIaYNESzqoUU3737
qzSiKa1Db1wCTNGdil8wWa3VO7s6OfbMS0/QvXXFYYeEquM5ozRU/wclLONtQNFD
QOYixTkO0G5XlTNJy51WzYS8lAzHrw13EOH9qdK3amz23gf+iga1a6cXSQqmenlq
Wfo0GZGFzhkUaGByu7RV4LfoeLvReceyWxCVv71nDeerMxceGX6uSCXVR4QQr1Ir
CIsNZZnFnwYYMW80safEn6j+5oYecfvwfH/EZZnVszd6/LA6TPNz1+DR+zWP3KAm
/hcZXpRjY3X/0SNntdxVyLStGIwVpZMsaguRvmBRvNZymcpJ75W+GLDsxIrfYKWI
cLRFCYnxA6+Rpqrtp3c3K5/DXHhfAgcYBluWtJCYsX9N09aNuwpmvwvE7pNtkrbI
EFE118J3YId9xCwfeMfVigjXhrE7LMOQPJVFYjvxm/LZjq5iOsUu5IOeYMy7cuc0
i4XlMLVoiDblSCx/RWjakR+p0aaUddOUkitO9bGHi0feYPPtZMVuUHF8y0csB/ez
/vCqYbjlejs6+pLXH2wxC4B6LosgnXbTddI0K2a+AaBz2+gO3gm5yiZClGv9/pnT
NAI1ICm3Acac1nvm3KT1jccojOC8/pzd1diY8QT5Krcp9pwUVawwtgNCUCHhQOxl
ouF5llgy+5Xcvv8beGB5psAKUxo/eGY/G2+VktH2zI50FA7V5vqDXhPRradDExQP
y+8hM/5zNJka6wDo6EO440hAtYZS2S6VmF3iCjmX23CpMOLel4fKSuDJjMACnlv7
CNZv0ZqIJ5/QCS/gKqCa2j5Saa7Ci8s+HgWlPBpD7zZ4uQXhxGEXmASQYeD7w8uX
EKuFzBEvN8tGQBkz+vEZiCzKPqhNg4FsqZJvROwXeJpdcb1OidTD/lp14hnarx8F
EiyG8YkHwLAHLyKO8km+ixeblfAkJPldenfjFrcIAvcrE2+WgUu/EZBMV1J9zqag
QIdI1pJIpd3J4kSbsRT/yUAaMh0sUUQ7/AoJ6XUhiI0MRqC1mzzYyolG6UGBn3EF
wFzNe1YrHsCCsplS5las9HMfIVGIu8/nf0HATARGhURhbFR4Wsn6wFVWonw/tFuK
cO6vsSgwD2SZ1u97SZvUEELyFH1Q4v0KcrWCBwfsEtxiV84BDLUpIA1KqY9d3H4T
k7UHdoUZ0AcJBeFyseRPBP9cM4NiVJITkK/4WzrPrFEW+yyZD9Bd8Uab5RXnN/iM
wLhCw6Z/bhwtu2MLHj5wkOzUbvlQbQiKUWrEwMF3BOqqhJyeLLoc71FLoyrukgLz
IHsVUYClIL0Dqh/9LItbpSv10tVs2QAPSQaJsySwELa39UlTeIVMqtvR6IECk9vD
0B+qww5/7Y2Wz3Vg03MaEyiSxN28xzFUcJLxcphhYTbtmJpmLW9JxT40PgF9HfCP
Sc/H7ZPXrx2F+4uzPj9OCJvXwip8BRyjAFC7c5A9mm7SnRALDglZyYTDcSp1ra2z
zbczJvQKp35gRf9JRzb+4twEatE6fDTMr+YnTVVuJyHQs6kVd0WQcmgj7BY2Bhfo
WXHXfVbwZ31L5HsJojPwo1zw9DIcgRqQjqRbbd5QgU6rZvx7NUq4EHx8eo/ehyI6
eSQ1T0lnXeqPERXJrc4gktHYMo1tV5sBajyCxJQx6I38vXm+FhVO08JcJ4S0rLOI
0A6nww99iojPBzR9fpZXCicG+jxSBnJ2pVan9vbTxJ1Gaq+grixwH0n1SVokuSef
MqmghtehoyC0Z2Ms80j7mxwjOHEWDcZJN+PYZFG2jYctWoB93+Iirq+Ibyk17mLV
QXBWMfPyyTUoiuSXHvAyBlzsdguO9+olZrmqRXo8CKq30b8L38yyiGHVRAEW4YXt
8ySfqYOCUo/kOc8iqz5ENQq20MpnOGD8b6dAQxTH0Aju6q8lSjOvFR8+g8sKEN9c
nrNgpsjxI2LkQ+IU8gy3d4PANDxxoTknRfOnJeoPCBFSPGzRRWrHqT+6sV7vyo5Y
5AacBffTpIE6ILWos6ilhlzNi5ew/JOTYdl5pCgEV7KiZY+jYVd4gd3/1tROSuTz
NnTz1o5oGb8s19gjdBVjgpREblwO63OiMZKjUU8plO8iO9Q77+rRdHNWdgTES9bz
vbBOV31wiQY2usiQHzgf19BuJw0wJkqXwULg4XVYLwhuFJqsuT5PMsiFlTjY7NZm
n1Z2cYfLFiRpa+qPUSvLa9hqKf6iiVuuKxqrbzTm69H/36avK2FpY+yeY7Pm6P4z
JGD/4fQrDi3URoC5rswEqUuqCfeM2tFL+kbALleho3rvH9UIY5Xgyd9eb6ZyJ1W4
O/H2ZTC1I1IPH49YQbVpDbRpAhcdxeTNxab2AFC3uVOwXIHZ+Jcrwp8P7sr6nYRd
oeMDkoJjiijTK0lVUqf/M3KRCV6fM5v0BGHv1aYQ8cbHwVspp6zYeokloxHFxpWD
hEzaWSjxG+IhSKZv+vw+bgFHh3pLLMKyNV8fX309+ipUVIc0f1xvE0HcyJh/UO9a
Nd/pyZXy4LQ6qvHQX2A20VmPtAtnc95IeQb3uR5qt5FyJAv5yCAjumKSb/KhRuMB
7xQ/QbkGxbE+seaXC02Jw+9LppnsuzAHn0dfNM+MZK4GMEJVOnmZsnvpQErAl6ML
E1tLau4b1pi/mSIk2WgGKqCoDdy+AO7qSH3Hjrwr1DVikX9UbbkG2r1vBR+T2m5i
qyxXzRmAtjz2OWP+CYI0es4bYMPCHYc+iMZNgsLgRXUN61U0LT88+DHfoDpMU41p
oRP4q4BUmWkKHJYF+O5KBT0WQcHE0MnHWdjrjSmsqy3TW9UiQFkRx94wvZ547zyz
WdH5yV7PgRlLoUfepQE6rpoaANiryJSAxQ77mf6fHnPU4sq4dPv1nxC+/p8w3b5D
0QtakR/G1i0R3CjI4JelfNzLf1ihPRmRySXbg8HRASqmg8fVFZ5EJU76pEXiaR5z
hU8PTw4H0adzU2cD4KbMjHYGhcBda2n8NC/fyh7DpmpuA14EBISpdkh6fzXoRvWF
2e3YpK40dZOZjp/i2cODvUULHZ2Ldp9SzkWlet/wxD+37KR9kBnAGcZZMpxFAc5R
R7+qyJFtAcLCsYvDyVVi1KqBegNeO3rdETR497uM+U+8YRXneu53A5KMcwOGRDPy
4Y7hv1XqWYMZtDYnJaK4nq9GZDdaQQctbxhAht1OPTSlcjeuEcLE9lZXH/rhI9rW
P2MMONV7ROKw3GSWgCZi3B3fgPE9tFarK56nQB5PA3TEx0HRbJuCGuvtrMQMFqsx
v7JJWDTX/BQmp15VBsXxxrHepdCxKyVJOlpzwQ50niMfCHF5uQO16yb+zcU4q0/W
8wrfiwrcXWIr52oWdlMnPSE7cD3Xz6m72fbFTFOyJIrhV+UAzo+qCxSJi/JNgtSF
K8dQXKAHZrSnG3nYdeH037gPeLJesq3xBO+Tp5YSyxb6aQPMOO5BqNByOnho0cKg
yXI5kWyQV9flKjnc8PwJzL2hqNB7MIYmBGe6REv1BXL7fIRp6N2Ap6a+SQ+zRjoL
Py1LFbAizO7AYUX2WMkByHLjcaqg6HFDpyTl4wuVdYGXgDz/EcSy07Ifrg3L/JoT
9ShAsoDTzA1sp0+q7gh/fyHpHMRNku9vrEFtTg7D0m7mOiju4EOSkLHc8XAnNthw
XLekLRelU6tv6ltxFmJJJG47ftx05/LrJHablT4lNLm+mGX8Dkch3V4Jnl6st2Oe
L5EjoD34FiMAKO0IKM2gIXQwwxHq/QE9iYjUhNjcXc6XO9dfW6YqZvapgpjvnC2h
x9LPqJ0oqsgLE5eqDdcL3/XEihDVDXLyitONR6pF6ESUes+3LDcIh8BWXg98pA2J
DXncBX0bH4WLK6Q1Hb8TjdnOIjE1B2gCLDXsnPCisJpCrOSYyk4BxtRA/kP8x76c
F76CZ4u4PHPZJgRpVJo7+s40DJ9UWwOhY21LEkB3yXZe4nYBnVbJFAM+pgXZNIVw
QWr7Oh5c4tShWcjnMcRmhBM9B0Yh4FNrkYt+GvYD4Uwr1NynrNh40lgzfkAO3gyK
q9IBnLtQmuf3T8M29y4THI3xcqPfpvrhVl3i9NWHXkLSAQbos1bQtO30IHK3IGEF
zwBLV8L3YdYdL6GMyrsr2terGPDO+GlpAve6mLKRjD/4dnjle9wte6vBnGBvfGFd
q49OW9QxbXlVXHyIYkLu2WUCTm856yzKzsREjks8rEE9W3UrfMZr9qCXuIT6nBZK
DXfUzZZR8BZtm2jCgXaciztHtqMBWLpIIgMUKysrqOU+/YPdu2ndF+b2YCH8ZMV5
XA1EWodSBuMSuToKH0X5e7Ez2B5e0NuDBfPRnoE6pnpjIVrvA/k8klJH8ehLSc5Y
ijhM24NTmfXIX0+9Dy/FmxZiLqEogzg5NgCfFA50Rosr41BO76HVfsKWlQwcXUKs
PX8pTUwp/LTaJ1TBWj/03yOwrB1kSVOt7ifYM4OuqGVOg5y8PyfR86X9Tv8zwzAa
EzD59Zvs3/FQ4y40bmH9aZW4SeOZFERKDeYZAbEBdlwSEIo0vCh2/5JtiKMxXQ+v
UTldal3rIMn9mBk0sGDYwdqidgnJsrlyoqx0DxMxK31mREME2H8bi1Z/HozYJ+uU
9n4I0YhD9kpXZeFA5F+C0l0HMYvnwCVAAiVR/xaMty8ZAvZCimrTR9BrE0om+dKn
miyYEc4p5llRy2W5FwP5y+DZiijuGrL+iJ/DBjSp5/Cx+AtB80pqwCBIVsud7QRU
1U/T3mDiw6btGgmTNlvbs9S+j/HbqpHZ/TTsOGfhwTZ7diboBJnxcoCrGfOkBQ4q
z2eMbvZrte+b8zpJeYylex7dSKJMLUFsMitNnP1FsivcRbZrWApRH4S9A9IfmuA4
Xp8sGzmxg+FgM1x9Y/qZP0LN7SxjmXlcV6ZNkuTNI+D0zD50e5gMjDKEG4GGbSUv
71cwrJb7DYAXoGE3Ho5VfAoea+iB9ar1QUYK3ngTvyF/k4STn7GnFHuU3JQKAV4l
kDWdW15d8VtRhHuZ94i+41ElyADr76Gc+yDaN75JP8ZUrE0BDyvfX18MW61l6bm5
V7Pak75DkoIlmbRwQiVt2DokAwDhH1iJPT+kOTAMybLXSEujGegmdBBzRS7nCE3D
FPqRzX7n48I2zUzMwMJqwmq8gWm5fmVil/UI5GvHe0bn9xRncXQzgqH6ZNsCj3xX
znkNvlddVBUgT9SqzdRqFUATSGrz/hL0nG+mcA+nGLIztZDqKvDTvH+s5rHAYySm
DYHRvM+lyq8GvuMebuV6XvMnFIvuqIXWpGAueuRvts9mSjt1yH9HPNJWfRLoBPk7
I+JlUNkjwdyUJ6MjoFt2CoY0ujW+2OQ/8WRJAGkRyguq5MfBIHh+SlWV8/Q7VGlr
kZc0kgXa+HCXSgMF9C/5krMUzVsj+ygxmH4IfXnE4XuFv3JBmRc1bcZFa7XcKo9r
nEPnkgAzTM5cC2IVCjWfVNmMg0xW/Tn6o6LC1sIVRrjYgjE+rBwqfvZteV9l98zy
XmF/8kMJJP0X9G6xLM7U1HQDiIy9DOqTKTYzM0JXdNJFC3CW6NupUvC81OdIu5op
zdAzdoR6say43fVfC4N/K1Jrb3S5p4sgeD3N5PsoVF6SIl2wpAY7OEyyutJQmmmB
VOFguhjz4xXbZC9KsRztaVppRDrmYV2evPwAAOSz9Y3YbU4Hkpd8kLP1kLxPceDv
wmkRHuHtoDFzL1NuQbD3aRkVklLjDWPxgJJDZxpx2NA9mNGvWTBoMzF3+TWvYIjC
1F/+pL/3q3CAAE3L0wIjfllEXQDo+mPnqKGIZK/xKnilHurK4nOb2hPfi4BDUTPg
IyKOqgz8i3ZgYAF3Cug0uIYRzM59n4gIGJChqbc7PNHKrrkCQafjOM0bbaTZGint
0BPiT33c53gIt4LLB/Dh5Lj1/ZzGJ8dFxl1XCnTbOmgIPqCUnbfLSyftia+NDGSk
vkFaxHHhxFHfkwjDvBT5MM2hJPii4zGY0IUzg/4EApM6SqBghp5R0x/32zJ2rYWw
6i1/N3OtVI4hw7j+/rgvMt/4gVWHvUwaZyh9SmJF8j1h5Kgq5x9Nh2o9vy0fKmKe
5uq2fFXMNhoZaSh4G0FGjAwe4bRhdHf8P1HviE8eUokc0XA4Qt84COuUlTGXgAiC
k6sBtudcNT4ScZzimLa88vXpuCY5lrDOnXWsqI3Ry9bVL7u8pZgKSzxepqnffnWx
F4iKdyIk544hvvUBxOzikh7G8QgKxTOok59aPdLBvzSeqbfJYt8/E+VG5PahZDT9
vjpBvr3pV0dXeSuezvBiJNcaVz8wsT6D/vqUykWmEuTmCjTzAD9IhCc/GNFiEHlP
UqZZbH5t3V1kbo98lrRAVVJbmx4bxalLBuYfhQCsgJMxScLrsygKr3SxoeeMbuIL
hWlnQRLpYcxUXUSKUIqCMT5J2bRxIeMQW0mfD6vio0YrfdO2rBiBimkJmTsU6h6X
nOFEMMZD3lAYoJcu0nuEYQsAdP/kn6GkvPG0exiXLwOs//2A9nmRXpQ66Rhy9FOq
qZTzK958++g3kVyCU35vCqbinPkZBHUlXE6Q/PrHxeikmFl8Iwm6NlaObj63Cx3N
hvA8xXIeIQoazZq9OWs6djdamBqtmSjj0kS/PWdU8vAUu/lZJDTdcgzFx4sBloMf
WGIVFi0KMewsfr8IUTtZ8Y7EnoTL+I85CLRTvPTbxfRlNHuWk5iZLby4v4b0xTXF
06YpamCTKqy+xOKdw5C8wstd9Y06P7MrPIBSl4aUzmPC6B9g9xMjWUY00piBwd/6
IzPGJQv5jqV78qqdyKmC012n02ma6q7bXTReOrjGl81UnG8vsdhUWFYfXAruxHLL
2m+16njUXMBcY0jlIqd65FITPW6LX+HrR0Q8JojCGmEOtwBmWPGIA27SSDEfdVRh
9i5bBXdWsVbOrcnEuCHSvJSRWl0NL/mlcuckEglII2Us5SiIS6YlIqhhnKteLvzC
IqrATraG1yUxMjrwK65lUw9o5jzG2fPMHSLJf5puM0jXs0FPTXvll38+dofysaQm
oIorsqpoxajKu8p/FFDi15OvYMn7AK0Yjtcsm5vogQNay+Rwi+n2FXDYgrYHP38Y
F6ZQOs/vqDt2CQbTQ2ADCAI5N9EqUshAwLJJlSJ40WeZ2Hk9BiqilY0xPYPBGrHI
S1wWxgDssEt+9MLUYjjYoTEP5zi5t9xuZreuRo9FhvqvttdjPN6ZG376Az3tqkzO
Owgt34Cpwdw0xjYNbYVyoCpSvXAvprnvwa9w4zsp6YudxXG/B77B4SH240I1GQLL
a0PdqCf7CEWTEKaV0xYfKDWeB7FhFeWHqxBYKLFwlvDsRr/30vYG9QWix/56isKu
FN1es7HaFNOrvpuAEJ0Stfm7RHH1/Yo7NR+CVAvsO1C5nyOCzpg31ofpOzvReAzZ
gAjarQtA7Zf31yWJTZ2v8ZDNqElS/sStXcy0nrIKsj2CRBt0EKRaJ6LTjtmfsLJC
4TecafnYWtaOCyKgeln4QmxPoQwPhX+0lWHrA4mslPVkP0km2L+zNrVlWEUfUKt/
MG34YR4IvqN5hHW1zy3sP1Im/rz5A8C7X1Rqgh+LxC3OyZ6GJXeRrrjtI473hcNW
agm38+lX8rVPtkE8pc8DDvqesBtTnt+HfeSr+Fji6V0oyugmp4akrKbTVjO19rd3
DI3XROIXQsrhv6PKXgj5ZFHIsBD4bPMOvlUsP80hzWMQIvqDSyzxfS1ofXJwfgxC
MsJD2yw+gomyekRTCK0/lkkHVPDABPHX4wDAnRpaCol2OHaTX+HSmFQsSE9ZfG7e
byFJv7TptrzJeR4NiOq3QQd5SWl1BvU5MP1+OHlaMKJ8nrLNmh4ef2RiN7dw7+Pe
HcYzbEibo40zEDaenWj69QN16bP2i0jFP18VxY9IuQZSsxy6zikGN8cxk5Q4NnSS
DYNjmsTd5QMFcUrdufBljWoEnNrCZAuQ6RqT68Md8p4AGoA1e+EjhHnDK5muws+3
sjytqyLpYFChFIeVXGPdiQuESIttQtdtOCYCkLw9gzgYlDGP03MmdVTVPLvZ3M1u
Lfg56j2N02JJkTqz3D4/nWJc8pZuIuEOToV6Akzm3zO+buzDlRAhn4a3dUsu8zlN
KUSW18Bu+K/HRQSKeiZ1hxta5EuPza/n90xnqGlXUX+mLA36+VM9rYOUOzrRNR2w
hsCkzgvcbRpw2mONBEvuDfA4yEyqRIcuqqDBgK1oBsoWHIyUTrtkkhVznCiTwu2c
Zm2072O8kUDvlEMotoeYnUS1llFgWTGsptS10bVnouOW5FImcDIqNLScVUN9sKYj
ko/5ILXOy2r9mdkMPC7/44KXyuaUiGoEjQ8FooJpzlQ3a37wR3PwD+pZUVztJ9L3
x6VFhHaf+DA0QnDYoFunqZUsmmSFVeqgSbd74qaRrJaUVTXKLStFP3hGJ7Ea6Ut/
hOqgRvw7kDQCEhR1HYw4LdBbo8w5NAHNtq6sKPMh/emN+ra8fkwXbiL+M24IX9ri
kz8/U64TdrZPwsc4iQF7mg6y1Nik6BbuhfSPuEZdJYvg/1uHGDJrOli4yWKDkTvK
1K0PauJylioy+Wx1Xs9bXX+NbksOpFz9PuyPZAChTZw6/pfYkosr+qbUBNUAGV7h
NtBTApbMWHIOJVhupzk77Ughr5wKqgKD8LEiHk6vJEb43ME27EIpGjLKrJJZpIU7
vzCRHSMt3DkUUgRS0vuHZc+6jhOjui43Fh2NgrNkCFkAw1LhU7xE43nBZRcFpjF8
x+1SsTTK6+MG3DgA2XpiSGWFwnVF3uGRdZy/C09F+iuOlzFfMGxuGCiZ7pQFeewU
oFdEN+eLvBnWtm85gYb2TxaGQi+xa/BcYtgut8TPdCU93H3WaYMWPQRcIGNdfeg1
dC9doFnvJajmUgHDox4u4+ylOQPsiVdt9NA+qT14Ec93R/uP6av28fnKwRqB9IMv
xb8Q7mjyCHZT3E4vsa3WnA/AMk36k3yKuHDeH6k4Gv/IycT0iHT/8+FswEpAmqLZ
yOeWW0EhIXfB5csSzL/N3ocCRDiIJeek7ugQkZsbr7JlQh7qDc4YVyJ4PuH0Lsy1
67am43ZRYD+E7xPlcZWa626AkGYNVTzZ0vmD9UJcQL2I3dRt0v/rBnnSUZ/bUHqi
gld0kOxuNZHtjMQOYMTMfALfOjuFMbfhAaAFMXp4G+EPxAIpkx+pGIoX5ocVtqab
WBYCjk1Kn7HdTS8Mr/89mxMxJM1l0xf/EtF9uDnIKgxIXCIe4dM2Ipcf1R8pnSuG
oc5icz6cStWAVfCA1NDiH86ITn6aPq1yfcuZi4IA4RB3/SGPB3n3PYkWvGl1dlmt
fx4mdR0tgxwYbx8TuNEY8StSfuFnpkR4hpb4rY+lwf14PiBLKkp14Bu7raFrzFTY
UdBdrDuLAb9fnYNgIfm+E/QcJ412CmU8fcZ+iGgkQLm/wymzg8ZvgQg+oKuhBE5/
ieOcY9AM+mMZ4V4M+TxHVQRVJCHCkcozk1JKAb6W+uXZBhnoGLgIVuteSgXjwGpT
2hAG17T2SGcaSfHbL7Faot1FQA365ao28PZvOmckq8MUK5s4nrj2c4eOk0RUq3O7
jB+mZ7AGJ9bmparBl/hpQ/6iR4Jd6hXNxLJLiFbAg94qt2uKTpf6E225RF4c8nW+
8sHoJhMWkpvty1hS/v7yUs1Mtyplf4hJbHokXEKH584n30n6Wk9Z2t8OfMnnEwyi
VlDSYf5QkGsAhxqm3Nbop6pTCdfVxcBjJUR01XuN9PH4vzmSF72sMSONSEUKmK4q
Tdn0Nk22/cRoddL1+l+p1l/d9B1T31PbnJ0MkI2nE779+yrZNItimgQBkoihd82f
VTtikB+jM8AyHSFDrBoAtboDG8dk9gp0PLHyUhSBSsD2hP05eeu3xWGAxqp4P/p0
GHoPFOoST1RogY5+SnCfQja23mQvnvT6LBIqI6zAVpn35QPm0y7nsHcTe+PpkG12
jKp6I4IW6mbjhQYWJ4qHLLljMA9/GOY93njH/hkg0iOi+dZ4v6PMvvJJJ/lpWyS1
fvRetALNxSqMJwS5amM5JuBiv0FmVsAsPJ7RYmKOsLXNuK5jFjYRLC+Tko+TN8F+
CSjyfNqaKNE9B0Dz2QM861S1ZqX/6UDW6XDMx3qEXMkahThf+T0CqJpGC49aXyiz
k9PMGnqDnCaEs4UmFuc7jGgl4CZEA1X1UAU/0+iWMPk6k5xFxLinOHdu44myitqW
EnUoYVeXg7cLWLALUgpSe9Klcvz0Qs9hEpiF1fX9uDBWyYpMK/yrS4MdFISDa0FV
jua8eZLrcOlLAtdGQ6KSeauhJY2kfb4hTPQYcq5gsVXX7ZilQVc+4TQ2+AQGHjmQ
pn1guMzutYWL8uvVnz8LrhFR9tRo3wvx+GE6UQW0ibXLY/ORYmMfdKHf1sKKaZYQ
VM6Deh9BgxP84wPbsNOG5c7k3esOtj7ofZxEPsAAc/sf27uiMri00fQAqb/nUGtV
QVPR1jSJoiI2Im1NAOQt1R1HGONs+yxtDD/xnaCYD2yw/hcAnfUkHBVa9mS5NcF6
R4Eol5MpW4VTqzRlV+TYzrfKZorpJRUjZ4r5+M9r01AOu8OqnwwbNx6fsJtP8Jp/
bU1kY4LZKxo4gxQ+BiHXrGRxrw4YpuNDD/727pxWek/qhuYsazo9LpHf9hu7oPP6
rqEMtZy1wgDnCM5Q/KAkGwLLtGNObmYB58/TBTcbpPTUU9Znaf6IchMcuTFlYdrr
ilvuAesVH5zscPKNq2LF88bG4Ot/QAOUXiB6+AUcmYJMJdvXlLhBQ6xnmxGuJHuW
sQ4fHhmDCN7OO8L6MtkMu8K9/LGUI2MGsAubajuEffnihu0Ve6JbA9ChJXh4iWgD
JwuSbJIURgmLjmeAmFo/MW7aXV2kYlQXPh8PYZi3Ud+b6Zk/EftbHroLNDa316MO
/qAVXunn3eRTG7KJQiCTRv5I10a/ZzqEaNwNHb2dWEEsfucijlrjpcvasd93tI3q
u0Adl3u2wND/Fps14Cpjx1u1OvM+2yC6CWC0pA+7IpNPGFFcPZlBULfgcoOsEmK/
aw25KOVAeMQUdMSmN+wNIp8ZyoPyIE6ExJXM0YPzEw2t8hfRebq8EYutXW6PJ3VU
i53gziTdTACbk7MUwnAmb4d5b5+cdHcgp+5tWi6ISWFQK0l+Ctw5cS7W+dWQO+67
Gwwuig7LzMZCUHOH3B8BWoXtVKvLnvoS7LJqDudNNK9lwCcrfptnthAueEDeHZgZ
pruu84/BcmHnbmJhM0QwP/ac9xojd0zICIVsxQMwYu02yx/vrAeDRv0GMOs2K3k0
03w88OgHndx7h3doF71Ng6vnvuoNTwb0cV7CzA/iPzThJuFebfH2XmIyhjrR4R2p
N5wIbwC2gR9yJJzHWKWPQTp5V8ByEdr4RHk8JDBW+PbGOIpuzwvWG3QiKk0FG7if
kbE89umqhVozleFs0JSmM+ztFki9KTK2415SHdEHoxI6vnTmaBK4XzbYhlwx7MgH
g8mv9JWuCPgYvh0lvklgpXCYMl5HfX+INFXeG+w2IIlBXyt5gRjgB4FjcFlbZkeS
w0zv535KZBP5LUaMypjcvXFYB7Gk0ZXxx/FeZie4/GDa85btT2ADokmMCNgjyLnl
Wx3Weu12m+OWFBpXJBdq5SfXUHsnYxZITj/7WItXmlzsNN/Ref87x5nm9Yl65HCF
sPbz68tfoxxtQAiSujzxPrkbEeEPIA0L4RejIXsGqzyBI1hTnhF8jzJcGdq9w8mf
ck8txHZqTOCzNsQnS1uNOWAfRiBHNacGPKbIGg4KAURbz8wa0Ls4GU4Z2ouQp0ud
58LOmUBCLk1fP7ApgrxKbl1gMRrSgUUAfdMp0JQgGIjvs3qYBK/smTV4wU0Ce2HL
FlF5ZbsD9TSrwVMbuAyEzV3Rz5wJ/fvl9RAofJDaonOa23/yHK1vzEYMH7s5xMSs
1L8Cx/IdZLYgSrbxYo5nbeNIrkHTeAZafQ3xw4ZjNFcJsJmcor5keqBUR2U5dDrs
5CMf0C2NnsvDeSl14UxpaoLq0VkqpfOJnRczaXNwNZJkZkkRt8tHGlb5mpwSWhjj
EbD7DStgyR/+d7Cj/yDSH7EyN4jz6myjKwkyZ4pwhGzuQ1+i1pcznaSmErew7iuL
ts3y1aimDw3/SuqlwcOZMFfIRl6DT9dhK1ynF4O6aTN0cg5jjJs0t7ET3IhcxzNh
OcjSkA5o0KbzvL2RmU0VUhTwEDHeGLShhrTf9P4VUpCYdqv2t1pjHvIYIKVdJHKq
3FLSuq5GCdjB4qBXPmVGA+T5YfoVRBri6F9OoWlurY+wTZyy//3FGb5XsEWrdc0H
Kd/TODgy1q0Fu7cZKOBiI9nrrsOc3Arw7ZScweBV4IbwWOpgoAAgNJ4kx8vmm+vt
koDR1V9LbjKPD2KLftc33KkwY6NUcFvUw+E6eoEGXKREdRIg4QizXAkfuk7EnYrM
/qCTFnQQQsOV66VUQz+gTA/M022ZzoBXbbSM+KfldILld4ysRR0x7JV8sR2DquHU
T67+6Hijgo1aetq4sHcHKYVrfFgmtwn7CJsE2I376ps+9ADGv4DA8cemjoMGrqxy
bjNsXE/H4qfKofCKIUQEXx77cm51hIvsEo8UDdt+8dlVoTfKq+M9gMEYTAkDrOkr
K0wsG1y27THyhh+7Q71UWbHy0DbD/UMl7i/j7syDZ8sCwtiYsMiukLNmleBhGoDW
KM4tBXPyhx4lkgP1E+3kLHuUEHvKEzaERWF2GlFEX1k/+mXfgf2nz449tO94IVRP
NSQ+oDZnhWHH9O5xo6TvHaspmp1AbBvrdYq3Hs2fpldWfXdkQFTX8RM3q8WRqyKi
E5Du29X5AQQlSqUl4ocVZGyxsoWplO31LWU3EWSLxFivAnz+MPsfFeuTdDkKRplj
hGXWb6+EMI0M5/ULHcQup4aZPaHi+uMvxgiaIWJtQRq7oyCnb5X4UBW87LJve7kT
jypA9fRd6s2MI0z3QxtFcFcRRDY+pvHnrevYOshO20STJqBlZcipFWq4bqheRbN1
QzSP9YCRe+R8McXWUNb3PhWey/raPgcnM6cNDfqvNMBeVTSpzoKP7ikOIjTKRx8p
7vp7LnE2/KJM3Kmfvdsse2VpkNRhGNe2DduLWDrMEtDYRt5gHN0I28O02jjsFPHg
0dmPV5NKpgRXDdDUFtMjMlDfXCtFMsFKZwKRiUf3EqsUedLFBLOLlWUBfOc4xpik
xSocVaNDYEg5DaGthsUIg3GtXFy8XydmyFMRZYk32RqVbud1vCr4RFiQUrvpPF27
MA9GhfNgZS5+hymq5MkUBcWu9aD+cTj6LLTKjDI7YK/heqiPOPp0XI+zSd3ERjs8
mpAGXWQtTp+BTdGnyiEUh6VgdZUCHgnx2bVT5wxvNNDsfAmlyZ4aqAUF54Yj1ITe
+Z1dYgBE/Eb3Nlj/FKl8hVntmR7fdYHfRw9QDvdhohc/zSWfxt0XA+V0dBWDI4a+
2bxqYtYcDWTwdo8F8CgfiD021zh8s4OIyhVrjFC7iIOEsceKNvG9FFnTOzD7kXgy
Wi+yQWi6d+pX750w4s1yK8RChufdK7vEyui2xsks4fXoyuVWFXEK7YIg1eKdqdgU
9VPwEmOOM3m0qdRvoG6oViC1JHSIM/ACCBYciYD8ykS5dfJnbHx8sbVXBjItzfTS
q2FBGoiy2mF1py2Sd6fPZ4OJjfdVv1ZtFKokdTNyZjpGsWPoYMpjbLmHOk8XHouv
SsqpOn11kzcDL9V5rC9relcKT77zfC91wqEObYbAegEu2JorOe1CArwFDM56C6rr
iQBpvrS5JzrVKoHXN3PfTD3ZgEr8bDokW6kLoyhko/vLEKD70qNQMgL8JjVTOsz8
l+F6U+3p/wc3VAqJglVwe6BRYMtlLmGpHVwcmt/vK9JQtT3R5mZ9OzY5iMkNT5f5
VM5/qZPaGzCD6z5fpJAsaYMM/pM4TLlq9eiVXxZ3+WJHKj/m21RP8GcNz/SEpa8Y
SDbxeHTRa0KkSkJQQNZ2Pe6g9qlLymrt7gmS9N+ZWmFqnKpg+qHrYXT6aaa/oXPM
f68gFZ3TwAHprlI6TZbZ+YOh9RPSX33OyNHKOmF3vc3JR/xXKT1A+ECrAN7NfIt4
73y/V/f2UNqeLVUj8pTXX4VFhwg1x7vix6aLYeQaTIPJABlIVy1IvyvucZoWgbFI
NKe5vvqp5ebh/ti7E9BU7zMXDacsm6N4fFtslu4W8o2QTzXEFqWb9ZbRnkd8qMx1
fAqBc2DdtTMu+MnsvjCFwXcoRNm9aRzYSfQN8BwVU71gxU+seOSZHpr5WcemHkB/
oZs4OaumTKGfi4+Nrtgtx+IqSxvSdy1BtTibdSAun40E8KuFkHfLyHNY1+0j2DsZ
+iP4MOQKZVZTkNASP6jbJGdwSLoO7qIIds4cfuurKQNYtUh79N+bPn9VzT6QEBkl
cVxszUspDbRFHftRCY4Qnt9agzeAD43AZDIFN/fqEhwT1IXoZcVbzzODMNSJmk4t
0/pLH6szwTEAuzdPdtvWCPq35Q4ygrGgIeR8VGlGtvfiJid+jiQQKkubcUtjkZZI
4VSk1stfUh6U1UiMJGTVvDXjZoF4l58ITUS3OYQNc6n3xU1VGAvUWJnotOiB+yyf
/MOoQaMUu+IVaOVHMNV0B5agzyLJ2GNSqSeoON3A8frX8xAGvYFa4nSaxyBJBxDs
5c3IjVBjl6d+uAuwXgV2lMG48545YSQ0RXr5z5nbbVKX7Huib0BglMjs88xbhFtc
d2UZs8WrWjVGh5JIyC9PXfDlDd8cqaivJcp2gNOcF7u1uIljQ5m/Cw/tKnRX79zI
2+8nzU50/G2P1dywXws9c7ctMdjsif8pJVw41Gx8Zyv9iZQOckDpry8DYYD6O+Vy
H0fyxTO/tyyg/rlTo+jjKHk1mW39KI8W2kS7Yhy3J73xUInm2gLq/2BwtSWOX6YP
ciwaro7AhaXd5SYWGSs0qXs2/WmUDCvBXwOf8xPfDFAo31tLaI3Q69d9Loet1Uti
4p2MPwFFyusioxLQZbqQhrSCl4hphrkOACsl7WBcM9AUF6hCvl36+0kYqgK90zQm
oUh4nLo2qInALMCGELi+iRrle395OfTe7mFxRMVmj5oQlT+snZq+WJJZ7V6CoJJW
WdQJHl2v6AzVZY4I0WeAT23ULj4sz4Bqdir4Q2m3PrROQYwN4+K9G6wUGEg5au0X
ynJhmi6WVLyWZyrcEgGgWJcO9E5yJmd8cD9PamUsbfIosHuR+m68SUocNEYxaRyU
NlOCQ1ZdN+zJto3TtearelNipWUYTDT2mIPnXxiMAxWsl9Xp8D5dYBI32ACrhZE8
aFOuZUsZ1nQcSTyUq7tAX8ccEnZRMHUlhlrWBWekt3IeY3KaRvUE7LydBhoX2u2O
y2PNPOAWyRAS6xYGDgXxo/2MdyuZHxZWNUMwzygtNZjhXXNMgSOWdgnd2nsCuliN
9Jzt8to5YURyjgmB03xQw83EhtSzpjIjR/bVbDiwxpkDRY/DAq0UA9KXHLDn9XG4
vUXnf8CjKZFHOoZW+08Sfh4o2odocksKF633hSXSRAA2XsoHYs3sRQnzO3X07Mkv
0eV16SJGFtZXkrwEPMDqiBly1S7u3juf/Ln2+GRpcKROeu6iX144UAnnXRaXgsp9
XOXdGoFHBWFaMpqALEW1VTtbRsqarWjyLaEtoUlopp9yTA5gyrq1SWXqWcK7QMnJ
Wn7Kyg4r9s5HVYCa+ulCS8usdagWIAwk2JEOCWErgeHcA9tnIWcA3E1Q8xS2eg1I
ndp4ZWo67Geo1YAzAvj0aJw5hDK+erOZHwlrLlW1Ye/zxMSnIj7pQoVI5IslmpAy
uJ3/Hu0J8Ec/o/1XlkeiYvrOjd76CaLXigiwnHJnxKAwxiTlRYN9VgbmoNivPB5U
TiYpIiL5w55/zlKoXGiIN8SM7U+7XYWqWW39a8ze5UbNCf0mOtBH/zURD4Wxl2gP
VtggLaZTHHvasubWQF9SJq8O3cuR3thSawEOsSz0AnYElI37unwAgQiH7UQW7hey
vNV4cUgQoQytNYzKE1KczoB9GgmbySBkKBjloVBfItSeYez3iNW5kqQ9G9PgIGhT
P2mq9hr4ZjJH5JWJQYqsaSrOE/Sw6n+PbpHOkEbqfnEoBjLqtFN1Gfkx11b612Xx
Zq1xBrN/JDNcLJ1Njmt8Lifs2YbWwiSooWh9S+C5/J5MwnYGFACH7N05T5SXmahm
HQsbayX4urMebgaAcRKo3RwZ60LTp0n61+gf/ZZbZO6mI+J/8GMvR0IEtzcp0lQT
sHtt/05L3/lIQq4EU2lF+Bed00rsPc+R84GvcZs7Wy96RPcmBRox/JwxE9G33HnC
DZzfc6ljbt4G83HkMiiwhmAQHUV0iDBwapTyTQVWmJo7cgw2HsrR2KAOFlNSfRMp
IQkl37LuTV0EV7UzEQnRKdpugMwdoAO3Vdc8fFS0zslAFpqY7o8nCuACo5kSIZ5q
5TDmgDtk6SpF55DlPm8XGWykwFQkG+6+vl3any+BAkDDn4eAmqoyhAZ97hYWnGXg
ZV/Fq2p23Vi/GRGpIhYkMYc8mduGtMFul/BKh/tVuYVds09xInge4hngjG/nGJGW
KTlJP/chj/0FANBJ9XDXE96wXlN6N8xoC/1IerM5fw2s8GGzfSSF9ETKxO16qmMk
x3MOL3x8aezDHT5Nh8v2qym1t3UnTdD3l6I3WQDndGiObfQ/jGFTsiuuVOnVD80Z
9hkEEz7X1tw+qm8yg0vW9uWh6VZFLJTAcIhTPskKWairFSoB6w/0g5Z/AWIfNlU+
lJ8xEpUHYk3f0YeHPupBhIshi2GVa/v8eKqSU55XykAn1FX/mdFtK45PjWREwSh2
xg0VIkmTZhZix+SxXBt/1Fe072vnUY0eo67j8JUtd8lfBvpEg5gojcuhZZf+5qPJ
rSqYdtEwi0yoYHdCUxA66GOqpgNaMg6HqQ8bcdffRZ4fbstIYAlGp7wBxJ4u+QHZ
AFUNylFNN5TenayzyZIPsrmVFniaUHgjURaNxUNTB9fvv4hKTy4708ufwR0DYjQu
hxBNN5b5dxbaW7XzM6YNc19yzmZjViq4IPENUMg4azZuCBv6w2Yn/k1GgGFtDOZK
HkpllIMapsoQLTAmvZET6XhMnh97J412c7nQG0SF5AyZz5rX7jQD5beEN+1YdJPZ
A6K4p9AdKM71McQq2ioef4+v+SbQA2QOtgkKiePgzeRgQH6iQrZiB5IvtXfLtIj1
QN66UMJvJigTyaVVdD6koagveX8AeySmUs+XPk9xrAslftqbDJQO+zKyXC6wmbmX
CzxETLk40131kp42uQcbkLR/TBsdM2iAKTxB57TrzE3fvBAwAVe1llNwHxs5bwKT
6jxqGI1vXb2DNZKCobWM0lkYro8z8LIanx7na3PahNwDFFmtX2yPEDHCJ0VZQiMr
gex6ITd9mIvF+IC6N5QjRwA58zqzxRFmUQ5v0PnZuWky8W6EMueM6lpHOVQuinZt
rjOfsCSJpzDrlugWlQyLt4DSTNU9TDzD1OvAsyc4oQAORxV6AChIDG/7dDg5xj4N
Su97YQhWrkfziGj4UFYE2przOZiGQtAwEyXcFTBfOhcUXBwXuuaq4ZlLNuscSPOL
6Zrmy3SXvVjdyQ8snD0MB6ryi6wLaUhiBNNb1TNPltFqdIzxZCg9AYifxfeC62/z
Ixum1hkOHSmxcCqEs9H3BiR5XhfFULwHvVmXRyE6CqA+kvm7N+GhcXIqLXD1WJVM
WNoQnozn1ljmpHQ9N5Kw9dL9yr4hlrYKaqLupRc7Lt2SL1X3P85ChND7eu74B/No
+Iu+0FVkVUdac1AMPFdldgb17Euy5vjueM6ZozXcR6XklDKGGMnqXCB7XWOvf2+I
U9h0n7iV7UOdzKoK7OKCLET/qtKRziAreTeGM6qmWIG+6XH4rwTWmXptzAPfLp7l
yABGmVNKt8Ss9RY0HMo65naE9je9Rg8udjZgGa969QPyTdZJB6Z5SV3Llw1YPuDt
nFdycxO5h01B3Fsi5+G/TGvoj9MnB/bYQqVeayGLmyBF5oRhhqqF4dmcXspLhT7n
yWpqMytDBOGzDEQxjja7zyKBiNbmshLDvUcZBbtxsKBjdBqkUKU0skjCuELdeQ+9
MS6DRWHkMd8nUkxYDvEHe3FT0EeEfPuaEfwfbF7xhg7fW673hLCWICLvm9fG0dFI
nb5HtJY0urcGo35TJzc+/cZyR5gHo4t94xVPkXlivApy6BDUGA8SDPSGSAfC1DGn
/hMkizeNS14aPN6nU/RDxkbCc3pZ05OXgJPtnk8H7FFuTMiDv9fzEnF4YBPk7q/c
iyoAAT6h+FFJ2zp2HHIF1sFUf+s9KiYg+yS4SO+6JGNvxkedw7wItvtkSWIpwpnm
3SOvnAEyXnsC9QOysh2kakfPvR3btDOE26ONqwAi2HwP0KzO6GYdNcYgUvz4YISC
6cI6gNJ2OJSE2Q0vGY1Ejx3ftNkknDK1dqznedy9ui4qy0RY48CDVp9FrjdA5HUz
7lalQdTjFC+nIXyU3e9Lkh5+jW0AFhCDIbT84g30HVgUlF7tO/55uzWRUcpq/NQ+
bAxuAWHF6RuPYWqAmtzTOKGD6dLup0nunD5XrcMizpp7LHReXo0S54yicIueTiJz
uzPg2vn62vpllG9RI/qkiZdmqjYboQlh1XG/MsfIyWBzPEWF//s67/Lf8Ahv/Azv
sBTjw23WsaBSMHAjvWJsyo32T1vVuyYb5gsstCuhbusA4nShWT+ZpD9fshbBhNSh
pVFOgbTkcg9YDEYeSZLEn1VdvamgLLii0EfvYsaT/QLE9WrCJ7owbA9xhDGEUtlI
rMCr7hv8MAzg5iBIhIAHUrFzpvaSxU+mno1Nuiyd/ZmRMoLH2pSSAUfeEdBuQbE3
E/SwzPJk/QCkcNM+5R38fCXJODCciaknwrWkl4FV5btR9kcI9xJk7I3jwZxX8jcO
7hx13NBr++SHRQd253FWbYGgqZwOAkAJQ2s0n3lAxdhfeXPGurCeKunnsUlkrPpK
jXF62H0UbXzWgOIKqWg7+bm7dkYYcqc77irkN0qOHxQ+/uv3OtfE88Eb7oIsXqGa
A6c92oYGKp/RNWhL36MC3nJdJZLGsTI5QhEDqVE1AYF1ydNDZfS+QN5tnN4B4oyy
EWiXl0Xb4ABduj2w3UBgFImmciwBcYipaSqmXv9+89UXl83w37XvINHIvSiW0dN+
e2mTUoQnu3aRPiNfXdUxoNg5G86HF4rvR9PxBZgNVr96gFU1s0PVhTS45NEyanPo
Hzqfzrkytca4oJmrrRcOabKWbXehJLRvxN8xQ5GARh/yjKIkUBZewwv8j0NcMyzk
gn9h9yN2yO+Xe/fgXjsX/m5CDrShhnzHUCnl274KEwDD454pJtg7KTIDobnr+7k3
aPYAES2SDN0M/ilaA5X5foyavkA2rQPtb/8/AZTSTn8wCDjw2CtXEUX1qjY06+hI
rDh4vDiYmQD34Nech3A56IX3+nzZvQtS2rpaQ9NpHA8QNPPFiahyL50UH7mV7Ts/
9Fr5vhgAlwIeBGYO0iIzwODWXyWQS0HNwI1ZNLoCgFWyhtdEzyBIU7z2mieHIxXu
rmvUN4kD8QTuqmClpHG4Z+tnN0G7nfS6yV7AVGC++y3xe9+Vu/2ax4so3+sishCk
4/otAiIxSYqg11h1ziV/xV5ZL4Mb/0IJ0QWzRJc6qERoMra/pgZzLwL22OXJQho/
BHsSHEvlqjFXTHBkMGZAkcZZlUoq37NdNR+SNSFUIv8iKrMf0jbr6dY+dMhg9/Z+
ClkQi2mvC8Bgxuh3e2Jy7j5lmGKYL7u6wwo1mRIX/fDzHvdFORcgwIU4myvztfCX
6HMbGUpdjBNxbj1UERxoyzeZG+eplw0jQn3tlGYw2h5fx9YBiwO/tJrCZe0TIvbk
BYWbR8wD+2cPq3C6a9yOHeqyh0cH6Z/0AFevvTsPzbEB8H7BsCzhVBsPmFmkMc22
eiqrzRvV3sJ7qg9yJwakM/9vEDtjuEKWy/n2jsZ9Dok5fYEhxuA/YPBzTLv1dcmr
mnXBgk6nEcaG5XF1YggYZdbVe2zYqN2qvnnL5G2A6ygqgX3o1JaAE5RRzvqbiyRO
y2gdHE2Xm9e2SREjFKWWy729sPzAxvdSoMa65ayUktmWmcU4vVppSAJv/MBQcVOh
TtzqTx1+iWzc715bNB7LDjuR+P4UM64pMFih3FsYSwXPUlwoobhheWUaXnaRdl0b
7wXkyXe62/PUp0vCjsMATlKNEfD2wPgP6jV5RxMHenh0+t6G8+TTFAGBHvbmDQm0
jV05TVOgpNDdkiGWDQEyTFtqPEPRVWI1242yLLSLTqo4oOajSsSgXIRr3yx21bMP
1kdQQMiA25PU1U10+JgDPd0Ftpy0Vz3hJi0oNY81/lyEGNcFAtnTdCvj4556vJbE
QJsRuxZ96obHDGkkN+AH/CETOxDq2Ic85u83tFtImswfdsy86ynIG4cy2NregKQf
5jAoOjoAmdsGa3Y7oi2ypmSPjxPVLodxwvJaxXJj2mwL5wUvy4VZDv/xp/M6oPMs
7MK5rvbvpERZ/PWSvJymlh3sT8U8nTMbRWWHp6XSDcoal2J8e500PcVoPBZOqx80
6CvHrmxrOVlnE5NtpQomK2YDBcisrVPio8BW7CEmNVOIPH2+B+TPi+tdk83QhgX0
AWOwm6VaWQqpINWgsdCG6H0kzdCgehAa5kpav6T78f0jH57ImZAwcWbv+i9oui0t
87FOZ5RtxxJQfMrVGQAPUAJnaPh7LCGWU9eZ7VjOTqYS1dwuj5eQSRTossBsLQJW
IOlWDjMKkoRLpT2mswtFO7hEFOUG7gKbw9BAHj3wTakKJDrrISnkFYzq9maENPH3
QFvMoJiJ7wvZdbdC9K+jsalDD85mJr13WO7GCL4CKNnOmrADgKl2LdqPSnNrg/7u
7QzoBQb0ss4v2ULWbNOEfHV6CxqCqz7Af4/TAQBznkNERBcADG3+8LzSGdWTYwM1
S28oxTxD8sETrHZY+x0b6PRi23BjTgjiP8jFkJWO1rNqz/W6JrzpeF4HT9BZEV5K
zEKs31lm+h9V3R2jnFEIQOy/flTkpi6rl2Ke7ku0KRSkGHlX8Bh+j/NXHZSEhSQX
gy1GBlUXmJPsLB5IVJGn7UIvlL9C0ZpFou9SL3uB6y1i/TeFEbUu7BEeyxzRhlM7
5YL/yJe1TAtaG+sV9yaeK36IgWQ9Pd5xqGoQVbBeae8AR3GXheaPijH2/U0ypnWk
LRHo3nO91dyXgosaMdPV3A0DDhvJ2F8nrUqoCx7hcN4o0pO3jb3OCjCpvVz2DkNE
CdWGYrnrGFNdDS2UM2WrbkdBfhGRLZz7FYniYTLvt43w8aXy3UJu5TA2drMvAyVe
VzJxDKZwpcIkOYzA99jgH+FVQhhxdVY0nasKxybw5sRdSCQGyNdi63D1wH/71gq0
mqMDuOFaNTRYBT+X0xt61fIxvjjoDqbhoVDAC400VhVV0biid0bTVf1vBTCueTsC
Cmd9peZSA1Pyv5yaaMp6izxGnwGmwYd5Z0Hkv2Fak2mXXXEhHDiE1kIVGhu93R74
ont5QAp7T64D5Xk2vg7dXOD/U53FGtSrxpuxggKwNzJ9TgpkiNCGes+QvfRnxSyU
1FPyuJ6kbHArGfXYwO8Kk2Mhk0bl+j8ePAnX5xguvgP1iN/Fh8UQkElpNBFg/HJ0
zq03q3zp/fuEWdVsfKPcBvZaUy0zFPNLXtrNqgJXa8cBBf2yQ+g/xAIuYOiBYXSr
+FvOA9LmpBpAtFcKn+qSoT1Fh/5efjqKhEgyKmxeNTRy+pFOvGTR64dwIRemAPpI
GmToKvVoatZAarg9zKE13dCsXJ8AUazHVnL2uOHoSpaea4D95FwAIMmtAj3k1BBt
UMSxju44YJl4JlcF8+7uLVO08W9pLmTMXH5+jA5j8Tolt3hwDhzEbIxdpaTlcw21
Xf16bG0LgbIChBjT4yxbiZ1kto2anA6f9oYzqAfX8IRDLbvFht7hFKBzJiokNX7W
ErVe2sMF+AVbDZk1A8iTQ4V0NFhyrHwBfVUw9eb52RbzRgm8t1ep3+snV8GB0nl3
dUXM7mBKETsZQmDsVh1H+iIBUbPVbdtjF0l2e+0q+q13JnIHYfYhOBNxVV92ERWt
Rxm9oCvRwpTfaiI89z/Q9Ec5injGaMRlwlv9/AkR/3dULVVDTesZB+rjsolfa2aZ
MYOEOG8zRk1F/GQQW1SEAVxZTqrTqDXT7hL1NjYU1Z1DF35H60JIYmFKqAforLAt
uTXT4fnuXiyHudpiaUY8UOwkf/ZfsKbrrNAD/wlkwXZMev8G5RxIJObc9HgIZHAh
0ecun+XAXCx8WJaAVav35bjkbV4DTdN31E8I8/dH9plY0AfLF99Ba5VNPeY+sAsS
2wqWVILaUVu203rBu4EXgWLQ1Re96jiYw7ciLNJvenuat4r04qvZaTCzOYttxwUj
mYS/TOnWbb4KQmSbGdlddSdoI9bomlgKxX9N+Bp/rhdaywXECMPFxt4MCoBeXuEg
eX6UbQJiV6QH/wGTZxmhIBEFHuYTKNsL/QCBMnOl9bERsDuzrjmjB8d7k3+S9VVk
uvcHVcAvSi/oNTQHgOx5x6ODt2/7VwuZ4ptf2u1Abcopa1hvF1F2zcLUGKei5g/c
l2Xom+3LfVOoEPMC+pVDbdJz3dUnjZJhwnx9/drznemI5Oml1nQdMhxt3aqarpNN
83O03mDwg2aW0y40DmMbCzdUfk41iJ0lWoC6iuZwyQoAh1K7Rr33sbsao0HIyY/c
1PPnVq8amOzjZYKFXNKPZgSW1ZQEVlDjikWkmwxuFXwJaGgFkgP+h2VmcLmatp1T
GlglNw8iseo4SEoScG0sK3XqHhAbSFa+WJkUZk/tjJE6NNsH8STA0n5B3QsenwYG
nnMlEuiy7i1bbLmSmc+e6j3UnLOXUMoj67YsVav/D0TRO6DISXXLJMRaOTdR1ZbQ
Aufi4FCgai4CWqe1ETaDfYARHakyNq/ciEcKsBYOGtnRysVzDwLPrGkh0qj2NNtJ
ZPJHnjlZcZV8Ca5sPszzumwr7l4H3NUd4WpvS9coMbEqPsgG2y7pCy8134TPdM/C
0DA9U4yS1/IscGIF51TCYbfoBeWZG0PveitRMIbb/OBd+iT5rCaPXGA3ToMEWA4x
14UWAYEBoL/q5b9mwS2oykHmenz+O3RpZxT3FWuGmDiYbjqTuLQXIpg9kngXzLpO
m/5O0+xW+WFk30nwSUCzF94s5iz35qeNnN030Mz75AdJ/kCD/x5q2yft5naV1DXW
sMrzb4FVxOVUzel1DDYG/ujwNnv0FQ/hep1ylQU5PHi1pbK1jDcE1r1yw6yyZp1s
MsFmIADTdSzA3PJQWy3MKbWElGFNKgG/dEQ5O598wpl+00OC6QJux6EUuv5GP6RQ
3QD3YeZdaL+aHi6Rch4mGlP0+5lh72YcQ/utG7uUd3GrjYuyzLv5swxh3xhy/Piu
7D8nXec5yR9Y4g9tPLGrCA7I+EAK0LZOW+qcaWpTWSNYoWsMpRykUXTa7CXfY6DP
uj3i89xE1VOxSwd15eCZFGS6+VQhL9HUBqnR2Z/zwB5Ggh1myzNgXdw2DMFmAx8n
/8/kUNt1BqcrjQzYbMnHZ0Ce8N+29SENEg/6AStuuB1kOq3gEIF1ADuKaJY/Lzjq
p4xBwX7aXU8VayK8PzaYy2j0a7hRMIQcVvPyTZ1xyGaPT4dJFqCj39Ts8bKhqfZK
bwX3j+GYBNNio2J8Z6kSmfswiL3QIuEOJOBrDPmINFUCFZt6hudZFgqLHqV+J04Y
vrDUM7WCgutUqku35kn/QiMjCQpnNmkeK1FJmIjfRIXRiv0ET/i6QK3F/u4kMqEt
sjJ/2obbqUbZ6wT16TrQfMTX9Fr+u+0wm2sLO4MtPBGd4Y1NlwuxoNowLDmiDrbp
OheomJZ9dSdJpET2dIqcB19gNbouuYYX2RElhy28XzZwgRx01Yu1PP97BoZSCwBm
9EDKyWnbC/aGIwLbHOiZ+vahtyBDvDn4C++LQ937S83pYM8EgefGEq04tn+yrM96
ECJ5zpk/go5b+PnO/bHE01qbq3tUocqy0wBxym+BD6xJbn/5p//iTdo+USiJSuxU
8Ciu3do3KLweYv18tU8K1HMX/VT4MyUmaldGZaHQ4i1uXfvZAgZdEvTbtxz8MzMT
4LSNMA11PYR2LCcO5c45MrM2e4y5Ssn5IMEAZaToafsoSBnn2TQtfQzlJJuNEmSv
ZOEykYg4prdHjtvSH6tISa1QmaLqC8Fx5TXAOklgK5Xot8XLMkeOkAzFmFvcQDlr
KzitfnaD7NIN4u3XQMXRhk+LIcPGdHshYez/dPzJOMg64nF20uaQAidsn+c9VPoO
OwbU4w9VpnSy0KeKcvEwI5wEWfYsAOD3tK/DRt7tQZDHCVF0g5siNSDl6rQotPOF
DYoa0tswa/0bzq2NRBclS0ituqkMR2fyMLCXu7H0dfXoWEdSmf6fkcbY4sJ4sUEZ
sFYG3aaVbakFEsL362CWmVZE/76awUGuKVi7PgGkM/1903uaSRYIlhUfad+u2m7k
+6gvWjEKPof5sCtPA3/kpOFhW05FYzCiqx4OyZJZwERiBv9WfX/eNfEh/j7KXhN3
E+iBki82XgJQHSqz5crCFE7JKhjfNz26rIgO06fBk+9xKEHF6HSDiMLrGZ3OP7Lm
81IkUhexbuKpH4gBHCUMN3e2Z76UTeXcAeaSS9r0IVQg4etPv15E6HDGNfhVv/Lq
KB6nVaA+bo7TtmjCh/ux40Yw3uo0n6ArTt1T2lOR6sf4TkMD9sNXgK3fY9ptPkEs
h0KNU21afxkc4uw9Ce8uQ4qebl12PYvFQFA/0bHlri2LVRAdMjA2UVpyxXQUaTfb
2ErgK2ccL9YyokV04XCUyoeb+0yZfmkG6w62iwuhX1bP5MyAhJ5KCL8DJceJFJIp
+P2P4wELI0mXiK4CVtD/5EZJjWYfgaPnrTPBYOUGDDy52B5DTipPWzcEilguDIF2
rdNdpW/pspgtDkkfo/yEh91UwJA2B98LmzeSkW8lrE84R+G7pC7w2Y3JSI76qTNJ
9+Y24d0rMB2blvVEhJBWQF4B8UlZ+VwBA2/pwxUajopMjRk+i6aXXdgxw2rny3Ly
766vDdqc7LFz/q7lys2ZGWR6AEOLPft2pdkVpaoWLcSKpqG/PB5f4GhRt4HQ7H+d
eVCLf5KTbbW1WZ3qMbKq1VHmIkbZHddCyXSsr0tDzW5l+RI9sfz1KmKv2cX0lXtL
TRxf+1rTS7+Su9TOQcoYV+R1T3Pa6CqL9YND88NPJ+BbzmRAYoBh/HX2au/Z/0CX
MtMuwsLpDHc8sD0WsP3KSxgfhD4k2L2vjYy4X5zq7FM2+9swwE2B1j/5SqzTxg2d
IYuaHV2k1z8UMClUkvmxF5aeK8z66YS+q90QMKX8GQZMwFxv5EYbSUrkp5jUwAmC
mjs0s89ipl8k2VoW8VN1vOyTL9PFGikVGaJk+y/MMFZSCta3547FnSALjWt0eH1I
E67ej9j7QybQnW2yYpUOm4CxBg4BbNgMmeONl1G+7TSetiSLxPlOBYUvXH3bpnjU
Lg6CAodPRjLlnEM79A1xlHAjU6X7h2v/ik+jbUPv9YsE92PbzeDLUd0YQRJIn7xw
jM8twma+o+VoiPbIjydZzaHFP02rKT9o8DhO+s6DlxaLwxHAB+XhYmHlJM1cw9YC
vUAq8lIRTKrA18HiBC5pVp3gzBnWbz0fhAAYYEccRX0zWXregA/qq9ZekISl/SfR
AT56Y3tHLZh3dmunF7PDkpN44ADHmPBG+ExduRQbJAFhztBkKhXX+Yf68uQNaS3x
gREhD/T1CTA8Bmz1PA9MYjb/ROocUdc5uEAO7HN9HRqZk1rYPtxHBeeLb00i4+ra
UanAGbSoRpcyC2odiNO/R3Dl+SNu6ZSFZkdvv9bieDPev+q4+5I9/vl5powJIzwk
xT6BQf3YohLO4bqGDJ9sW8/U+cAEEsZBOBazmoake9uwnPoi4OXbgpn/qzznvbw/
fGicV7ZxzGfQDtm45bJevlcYj/a223pTEdwxl5YduaYLdaM62//gtNarvIlQWqSl
/nAKmtT8gV1vSJILtn0SBsiUAZdMp7/IzAZOpo263dUFuLL8tDZw2ey5VXY9HdMr
cr0Pi9dH2CWVOQwDyJ+GAGEdhg/nloQCyEzjt7GwJ9PNn49MMhLd1HdeMiRHqVg4
5S1xv/6TL0u3NgY0O5mGmlrN+yjG/OgmuLuVay3+2C1AYYqhSnHxLWngdpU89QvR
Lhx9VO5pKteemVYDmC8Pl+1AsalZxKaxAWAcW4kzNVUuEsbfu7YsrXmpQQdJV/Bc
FidmxKgMWymoFukdb/BD9VcST1wkO+gjcmSpDyKkPcOS6XzSyN6HjiMvwZLRgelN
kEO/DkkziW/ycJ9y3IaClHeOx23z0BXEeNoIBYZ6wVAVMeIzwUCMmo2+g0VfViRT
DGcmvH63yGzViSixM4uolwMfBFUI/e5+RBRDWEEH3c5PW0KOK1OO8LdSXMchteQ4
wxjN6w/MoHb6bJdsWPj+ntPpBKGao49pHxUwKaD4VpgzMHXjCvoB7cg0Fp98oOOy
xn6gmEu+1YJjpJ4xAU+/WQRsVyWpEbxUvVRyFOI+6pdk/kdZJt6t013E9r/yJiWc
FjoGdvHnRm+htm98Gt2ptiEDLhW6YQA1rKDGaMO1Kk/MOmCg3xhjHF5Vz7a1jCjP
IMs5eMBJFtmNP1B/7Eh9zWjWXdwFu27HpQ9SHIuEiCHnwOVdcVn6eimo6tWKgCku
0QGqRbwy0MgXSprydv6lGiI0wgtS53l6BG4aZiHK+uv1evk/7u4GoqkNYjpGuS1i
D0H42eq6bQ/PaIiHtDda3aeDm2UhFNQIzBHah7GK48FKhg1UOwLSGCc/g8EFQu0P
xF3TmHlsEAiFQJWxhwsVaoMPOu6sU+AmA2qd7crGSKUObz807RJBgQ3ljnk2+OZr
GiBy+cVXCjaMZ9z04DXAd6p/B4XtoGe2YEk3R1on8q0PZEyPBl6g4YKyJN0SPmD2
DtDygZl0zmVLp5ZsfFfnaAn067zHUVXXhh6JtSBIyNh0CdrPSJtDtXWpM5diA6vC
ck/ejvdL/uAk+E/0+KEnoCPtJFk9Ihf0GHxBWwrgNkXcl8D/iPyvgr3Kal/kk78w
S/KLgJDg1/+Zn3I2P7QUwGT/QnTs3fXZ6E0e+/zlhymkKEo0fj6aykW1kZvj0+Yn
ciAYUBqoLV9GHfaMZRh7jzl0+V5EaH9FWIOayOK/3v3UJNmAOFn9Lw/Wv1HZvalT
vNZBSxLojPuJj8KIAI+q+NcUXwqx9/VTerRUudk9bTaunGhF9IOW9uHnHIF2a9Oo
sSf3rJnH5yf7XGW2YYBmcBxOocpSOv3ivISkHvqQ+Yet3ZbmLrylxiC9wztIvLfv
H7WGcVYil4j75LU015M06/NT62uIBYc4NkN8KdKWMKJr0vPszzUQcY+q8mRYfq5Z
LVGw6PJIqrwBfdVpqW3tBA5mX5SxufiUiGxJc7RI3Hs089pukhtn53a2Plcn9GmJ
1jkPDfTP3YE/nNgRQZSulYehjibDfV5OKVBVYeK/+AeH/Peoe8EU3n7OXseSHXFB
5NsEU5KNHxAAceHTMmCAz5UD1sGmxzrd8JEF3UyPMZZMGI0foQ71LBcCYWTnLHVe
BLp7zc2B1KSobkOghhxCGuYZN7MEKJvVBP5JqA2ijc8s7W0aNDK9c/dNET+riFH3
wqQbiS+wVsgbPP4FivKX8BYLpkb7P1PSqUtUrklZ9DdQgoxljQJuoMtTwLPWfRIz
Dw/h6pPwDF/8S1SlT2AHPZZmaDeHiE1GbnnxUDxmDCbb3TuWknZL2SIxA0LDXAzv
fj6AGFJYGUzpQoLbJbg25NIEP12YT60lC5k8x+e+482oC0wkI3NDl50wcYB3h2mz
rWCFAb2MYSCDCvQmWO/NuVSJ8rCBXNCcG1XkDAbrxSE56o25Ud0dj4dPyQPWHK9m
5aV7AlwSW3/R2hjPtmlaXIkdP99blf9MXjmDgcyHhcyh3rGt88JyalEd1WGw3naz
/Q25IDZmTwI/oEc3FNM+C7UqbjSBU4JlH/Eo0q/5TNAscv8PmTZX1NqGbIP1Wis/
oxo7Pg1PqYpVX+nBOHRYw15bXlQIti+711UYH/Go92VAcCB5ILmQ8ky9dM4/eDHT
NJMOcQqKIfuqPmYNHbbPoitayD8NaK6dEi5MAl3F4xHTLphqZpSD0J+m8nZb8tDX
II/gDd0MUTCEKso3rIEquSvNjjUK1Qz0TcNhxse1AZemT5+cFeLiYh3fqUhkv3Ne
DsRDDI8prcLeBjEdsNMQpD6lp96PkaRISTfM1XO2L4WIKU+1Yzgb+cNoHUBBRYp1
aHN3eb7wNqiYphwqWPqvYUHytClIgLc+r4f6ALe/D33QmNb/OvHaMeD0lgtwCsE5
VZB4x7MY3v8/5t0OoMWsGGokGJanNaDLGdoUB4PdhLvr8NQoEaO32QZabL7vhABK
BUhHB9cfuAA2SwZ16JqrjMQIhPg12fl4GwCVzIHzbSo5e038PWMK04VnOZYkdslZ
ZtBZ4ipamRayQCH0kbVfRZsYR7QKfO77cnXer5AIEWzMk6tI0v2sDEs11Fi3LpfY
Nsh4XMu6u033uJCOZ+ThoZcNAvBdYjlvMu1s2iwxqnCI/a7x9d91gFKM64I/RskH
qwHKNiNmd1O8gbrV6He98lfmRGddtywcivyoZLU0SONVcYmTxpxPGQjbZQFkZMgf
0lxskY9rDN5hA4X3fLAtaFxZi76zwQTmgXN+tIyAI2Cm3NDEP1tbSIoEnLh0mXLE
RyOu6B2PcwiaSa62impQ6YT846FP+lg1WKfJU4gF+pl1SkyjhEMNJETzm/m6sZkK
MLGQTI7i8xLgtifhYXVWvu7u93FDe0ggHQpYZd9q25NOZ3CiJtGQl8opHafZJYe9
Nm/UyfRD7t4sIex/ZtsTn/tuTJK7bicxoI3RMrMb3QFmbJ8OVcRKthLIasgXH9KR
2lpTtLQTb7664eh2DwaV+eOD3N+f8l/NiIjBNUaUHX5jCML2YrNHUGPB1oMvvSHp
JjdfbiWrsZaYoAvG8u+uvmm2+OdpcIKM/8RiPCT4aYd/wnnzE0XjteGExnwUkgco
ecHZwf9g+HLNdllKqLP78P6N7F/ilI43jqW9jKwGGmI2PjCGALFQhccOvJ3OUSlt
ww2FiOKEWUj4Lw633S6AHaev6YeW2COmrCRVK+aXEgv8xBKmP3MrZAM9GdGEtfQ3
XE2e7ri0Gczl9HnQ2t3+NT1fiZfz+5UN//4UvmNgNMD3rQXJBXmZgh2vrC5GG+ln
CdiEyaxJoXx2L3FrPHe2kI6NMFXTQzvuBgEQv3/JliA3qIOMETQFpodp428FauO/
v8XAbIYnMUUbQeh1iR/VjHuD1tiuD7a9yEnZjT7YslUPzG4akmlMw28sIBPjeBLX
1diHKP2LNnFsFnCgBooJgp/90QkwFXLiDbMqbLsD3kGZIROrUALiA308zyc1BndA
gFis5xP0gKhNGsqV3vf7/ybE6ikt5vNUGhQCLGF7Ub8EnfM6mCBtlAhIh+7DhE6R
Wm9E/87uUkYs19aYL8B7NeMhroRJSdJ6cDZdqnqQGdZnOgy1DvJTfN41W2GpYIwa
Hy6mPNeQ8MBOd/HEY8vsEiEAc86tuJPN/2wSTUpA5+1TzkX+TOopT+Ln3YlvMUGM
ovuWB3UgrTka0ULZxRDf19Yx1ftDyBiUkWWNn0mj+YEwxc8O9YjcYHQcL07FQJHQ
1nvBJABxCwZxfvyOi/FbFBjj288L5lBGtotWSSnelC1GzwceiOIZlEmR98KFHrv/
JFxKc9vqnpDEEE+OlBkqWNkSgqOqj1b6R4FKq0oqzgUeKHfx6hiPd/NaWo4sKaWt
0rSpk/8bprQx33849d5wcqVwh5fcPPIqylZJrQ6mujT8cwGM4IF5vC0nKDhzcBi5
g5yshEVAI6z5jWkKojH28lZkY5qUQ4Qjhs9qtCdx6pDI56PRx+ck5mM4pTrDy7AP
OAnvkLqqsN03MNQuuAl89WCTY4T2/hUf2lXMlT5kABWC+AqQeUkcMV7DCJLNpSxG
3gsWxdtexUjE8Jn4Zrwln8YXNyeDjmaHjdcPvrRJgvDdGi3htaQs2R0iC6bCV36U
9ZfkrRRwbDkHpekdY9vAjndBhJrBeAeFw0CABaHQe3SHrCcWY1/B3VwaOwyVKuW2
YL1lvnA6uzVZLoX1Wmk0C67XceWN3x+yYj9wLtToOzDaYmMtyQPWQ6+M7dXvOeow
i0Qt2ovgWyh1eADd9pJ0j4GE3+cyBZXJiaHGfOjSK6/T8bMBo3paRKngVkIFcKU4
ENM+FHJ55rH+/Xo/VbFvR+CTrdFAztdxp5BLFowuOrdRL20QTNZseODdwBJcr5u5
sQj59YVXG7oCa/djDaZaYEQ1ew6Ztl8+X21s8XF50zn3JR0hhKfvMorKfuyNJy0u
Z5/CL43IFv1/3auwhwKcMMSTyNrbcO1n63mn+eGo8jLg164PXEta44yGSV+x5N0B
hJWTQ6Q52amWY14ZGn0WB2aVRWBxXcIklkrgqIFIyqXe7sSCzeabLU+Zi7IA9oSL
Czsafkc+O1sQgO2GliY3PB9t63RLLEjt6C/fuPrdwxY/4vIngif3nr4DqA83GmZ7
j40r4CTTEJLdrxJFgfVhDIo25KbHdCVF5NyBnuZof9b7/uHbVM4/Hy0Nm7YZ2bpY
TlDriQQYS86lLGQZKe3xFOBh7nTJ3UU0GglegMbG2tV6lIb7S8MBloUav8uuqu9q
kvyJVkRc1ZxdWFLcWid9sSnuH0jGLn+iR95DDtwWYR1L8/bOECXr93ZG4gXvwiMF
SLvOLTCfoausiQJ5d/HoV+Vgh7xAFQ7voKoOZ1Z/wBkLKxcO3kaett9O5nmTR+6s
ObU2x+lYIu5KnoTOXW4q9+FKHtwcVV3/dpeiBghJpaTd5jxBzM7EhHmaTQgGMlKD
hs1RJ6Z/A5l5rPJT4OewXrNwJ5wI6RJ81n3r/OvsiTy7GbEm7thqj+LQJrC+MD2b
YevoCxWNf+vzZ2j0n+Ztu3ChMocTbKC4TpsUfgCxDnN+wUHIo+RD18/L0Blc09OY
ONM2aSPIQBn7AjvUnLtJ+gwAQeb8ROGToQdXulQamBnUJPv+hzuHtKEa1Ei9tMoO
yKsA5f2a+aaABkDFLbgDEDeXIdCRGKCktQQL+i4ynnU9KmFNWjkmXh0hv7G+F6Md
qgMczAfV8yRJRda7bfIq54tZs49v/FMhgUrWwZemaB32Q7NzdS/ytLD+aLPczQVJ
N0/RQzMuBP7lmW+0vX9eJ0pIChns5G1SwE/QVTvNPCVkF1qJSCdlaECqXPjf/TOs
Q0qe1K7Io7+Knn3/dM539/8wtLc9HcIiIjI6x9h/SbW937lhnuRavG2TW1iU6DmO
8pspLtWUouuWMiqPioq+46Z+qpvf/X/T71OKB4ou+pJ3/0PVHZq0WdmSH7NSo2E+
p8Wg10jQ6eLrykDw72y08bsXOLoZthC0e7KfQsx+QK/m26uwvxp/dBLflYAK1zOh
OHiAgB8lIyxfSzImmGSsHzGRWnhloev2lrjC5SWQor5Nt4mI2dxfnylNiSWEUs4I
oAIpCP7iLCDkZ7wbeeki+U/R7AMQhvqQYnpGyDraywnrUZYjZpK+LdVBRq+94tD9
B/1+OmrsWisS8PWb+5yM+q8/Kn6cIag3ucA8bQLTPdVQznucoWKJhIpv3KlAP6KP
PhJvYPCWDHIQTcGFCjH86CoolTE/HXuiK/FeQTjJOHSF1Hx8YhWdrxI4upsIWCxk
1Wx6XGGUJeJxPLDVnJlVjOHjXWwkhmhGDN1OZq+a9pAI7h89VyUef7HubQ+rIxOE
ITWzMzkCVakdlhGsljNe1AZ5IHf4IcKUFQ9aIhdI4hVXvN680QJhAdXN8SgJXkT3
5T2q2PIH5/KY/o4dABRIPjA1EIv6x9Y+aRQ/CR8f5lwvKYRH0FJRIB8BeIXnboRb
N9if0fvvV8khMSLXdYfLCK1FEw5xet1sqYH3Zd8kH8ekxsaRi5vxH5V2iAEB/1hn
WupKuulVYXsQiHdXJvkhKNGUd6Sf1niJgUsshozLMjwtiJi5AGSkMlbbNh73EiFL
lLm/6q6om1rNFPLi8p6X4+/5EmHgp9dgCa1JA3VcauU9pNdjeInk3lJwzpYqCx6Z
662s+KzxUTa9xoL3SArKjtp5wknp0zmoUbF2wW3BZj30njQH/cLomZ1tbznAIOzg
SCzzRL66RJEo5lf01gYY5rNAqPPnSwjqA/l9kR2ZCoWh4XIdhp2Z5QRrp3aSguH8
67beQLZJg0szYTB9KY3NiaZqlY5M6d6hY4jtNHXqxTacPfliLgoZvrhqBx+RSHCo
UgifKBXQjh0LEbmAQWDhE5p7Tmggzx248QZKUdRXsaCjRHFpRHZOb6GZiLelFgOi
uwU1tdbZ/sC55EQ94gUj6sdWl+BtGYVeUZOgayYfrZ+oH7vy2rGae1eAFS/k6WUW
lxEmCvS1lvKMwFTsp5fY6bcBz79vIDAnebetlstzdexA3vZgF3SoK9OXYAmYcPTx
z7XxLSXhwjiATvxWObulnlZQoL4KqxUp54jea1Xiq9uMiiqu5D04CNsxMPor/o/J
ShGnYD8IjT2fJ1xn26YOr6yxC8Ln6J2Xeh+eEawq91j10rXKLb9auE/Hiit1tlFC
1J4bxk0ncIyQx4wFaNzlzhU55VkDObR5QMVBTEf7mEX1BB+ywxquJ5Sja4zdAMdR
KfK8Px48C5v8BisAF4vbCJjjpuBFAUPosWe5Wb80Pmw18KRPlsbD6hLyf6+Wwsxt
lh9+lHNl98e76KX1GDA70O7XXgXLQAc4Ga0n5dityyRLo1J3HSEoF/Y20wOy+iuD
gvu32PLPyqjP27M7lJB+FIXQYXYIbBx74+q7t8h2jM+2+37AM+b4MW2vV33Cv6kH
ayiw3dbbq//h8sxSCI9kN6ESNCCoZKzX+29q1spJ+YD/mII6OK+ZFyDuLjm//UV4
Bp6Rl0/L0wnjCaX8NoD+JsqX3/dlz7d5zg+T8aaKI1JBzbsvdbQeGSlfCkaHz84A
p2VMczE23jpOznjUZBvZ/Kfo54nvki8zxxvkSqJCoe81O8ymuijFfasxTccjWdcR
BcEBNeOYmVVZRaf44kyQdZcLtiYooHkvOviBDxnXsJJF9PrYrNlM2+hvsauMKVcI
AF6qndfu+VC7tHZWG7LiuIp+3Ofmk33UFN5fo2Fbpwk1Lr8R3ZbqR92vcZyzQgJy
7IrLJfkwPfeKcULiRLr3iyDV7qiiibl6ptLEH2gXwORRL/w4kkjO4mYsiA+Z6JG2
Z/dkMlazJglfKgVGDPcvT7FEv9Xb49b10INv3czbz6Ot/VuhNAxAgr+S/hw/rdQW
9ZgzFFBkFDLjdzJuQ918JX8mTpr1twcDZhtwxv3gEJl/C1hwdLcCXbvyO4TcSZ9u
Nmr/n10xHznRVx/cYkovCh1TtehwvGKjMs6ppMBzEhP2SEEaUJH8KEdsi5O0O2Dl
9rWJY2+TpbSMjAtC5EEmev3zbO5OboWl3cATX56LWmahfzAf9oPlzit1OZkSNH0c
Fg3tA2NvD67V7RvHL68pDhGpF5bi3XbjmPMKNGambBNDUHivxIXkEqKa5BvGDG62
79WNkBm0xDB8lK8x67oTAF3sMfwfzg14oxLHd0agLJDM2ImN42k3M0HBAzScjDiD
PQJ/O3tzWqExZ3CBZtygXsUYPbxykDD0Ot8//ZZ1QNUBUUOiYnQFRt57ObKduGCi
JlBerqB7xb/EMvqEBFFdk7GBhH4KZPEUZ9n2EPJQC9IOXrKwb5Hx5UjvIJhNBZqg
te69qwZvwLK0oCpk99zWjHBxsdCLq0qXnryQqZrzi5/lWy4qPVoFEwgUtWpvdkjL
ufR6l7xh6GMCmJmb5DjBvb1v9jpnCg1W4ImB2giKV6k3N1g2PX8B0cDn7DNPsg97
2mq+ndIhXiUUmF8X6Hc8eWFiZYHti59dnleUb8xoH7PJQNi+fATjoQHm0vtgS2lW
GKSThk3RbuY99uaeZzrvWXz7bcF7ngNp3V855gck49baYfeLola84YKLJ2cNSvRE
LJIW3b1lGxRV5DSncurLuljpcOLWMfqsOhi3iAm0x1hpXcHvselRVLwYacnOjB3H
psqL0OoeZRHlQLiVGCclQZUHH++uHEctlt+kwE4PrBkXU27/pDJgS8pUfYvvO7hc
NNbABH8NcYw2EpwJRReSfIpiL3gvOy968BsVPiCVaAFo5vcq8fVNDIFLGRKWrINE
Wwp8QGsFsuFMHrJmhWnxX3Sr2uT1pUfhyLj2m4FXBPSriWFqO8I5ZvF6IEpoLa8l
esK2jldaHnnKNHmrE4zzZV+HQ98G9kwKlPWpPEH77Bbwqw5fG4Y/zhoDdkP98Wkp
8TZob1R+d8Ft7JT7+nzogKDWJ5ZzTyozyPWU3f7htjHywt0Skp49R/B0A3dykVqa
rWgswLogXr/1VHY+T0YNt/KeQTx8wh+AXOFTr/HwHXdY9muAE7ynyc5pgx1l+IOO
n0qye2PQi48rayiLGQV6cnzG4IBPvQHcFfXjsN3RQ0qkcSU+XT+H2VbwJDSKyGze
+vsNznx/tt04oYAvtjRaVvTdQgSUrOgZNwJSR2VJANsu54ymi9zb2YbDGagFBlth
TYcVXQ3iSXht7l1FO9e51f8Ax+VMj+7PuIHID1V/b6ukXa7PkO7LUhEPUF5I2r35
zPEsttS038NlXXxE0Xa+yJFQ3M+X0JF6xkGICZWAkimhgD89sA9LfV1GgSmAzvhB
FIll5jZO7TdQOXQ0vdKDlGReEAYqdyjxkOWhLSbIW0wV+/b7I1ydk6lmBZG6RLXr
KPyf5cy9kgzWDRyo1Rr8CMjjUVM5nqL1Sdln/5+PvkJxCo9fsWtLqu85naDZZNTt
/6D4+oHDoBsvQJb25tOcDIcxVG4HONbPH7miZpmZUE5ten3EJ+qKJMSLTT5B+dM6
UST5XM48QX+oZCirmX42Eq5LkPajDYbyGdvtqstFUGpKJV6xpobyZoFXcynNtR1A
Bj9YLuClAVlcQtETWLvPGsJdeZ5K4VT2t0mR222B4UQya6i9Dow42VU/Z0KnWyBW
gCzMaW85hUggQLa5RaQwFf7WVOnMbApbDaaHpPRchWojD1VdxCDribT2ulqZu05H
Onmts4lVehn/1nMFMdgD/ikoddNx+dWTDkPV3x2Sua1sQrkUGxFrhkMTIT61kHkr
KkCmcljX+7AQpQN8wpvZOdTYFKKigOCU5y2FU9sCppWoVzjZlLdVF2jSi8ZTAOX5
IXh7aBMGxo6ehxPELSTJSzWCSNyCFvJ0lCQYdWThnKSGI6PjZHfwUm3sYDfKuLxP
tEt5ovzCTWUF6Dvkjbo6M7RGt/innOwOb6XGplEyi91go33QA5VTWPZS9+6oQNp2
RsL+u5dWoqjQX72PCQ5b3J32I+mom7dtgot6n5uCkrb08tL6XMXw1T1RrD30xQck
5B22aHSNNH6+E1VN1vQMP0HkaLbzQGha37oYhDFesMY4iWKa/KeqaeIJyJetlGyT
BFFY5tiOIydIL5UQPSt4YEXPa1VYkL2w4zCajcogGZGi/OcJ0jIv6KWyGvfszRqd
O9oHkOIVIG1nFl6f60kQ2JdsO5PH9FZVIKUBKI8csO7byk7dQKFrLP/nk6/8k8bT
TODCZ91/Wn/MRJ8+zXDtGZkA0HIHNYraNsDk0xX02KC6m3vAMBLOF9XJqsHU55yo
n6sraGmGay1wAzY/9dgLXf/mcnH+lLuJf3Ys+3O4kJeOBxlD8yuMryLIThYoA8FZ
LIPYJvhSrhCxamZz2URJC1hKmpKeNSmJkOqKiWuUIduUV9spmsj5cPawmGqTTQ7+
OIbcfEwLvnppmd7aLjO4Tm362ah1G6nGs8mND16E0rWbpxVqI7bPFiDSsE4W69Ig
8x763NWYZ6h8vkv3ngY6c8bKQ+C1e9Fl6C0nTz0HrE7M7SXXyTWgyFXWJiI9ApUh
03ccOZkUiKP22jyzXQInZBhPApMSEK+2CKD6LASgT9A+X8uCe7/xOcI6dr+1QW0n
maw6feEn/cox8dXCR1Jr52EYoo2p097EzKaHAOY2sei8JPs24kkHCxwd+KJsX0Fd
pjYSnW/eWWUyfoASt843tw/asLKQf4n8KVGjdKwcSxI/qbm+gpZSqi7pH06KE8WD
IVfq6Eh1OrtbDYKBRiC3dxlRZKsbpdOH6vfld+JCOySefqaOxcETWfAtf6AwcmJD
KEGL31cRDmnA7LlZ6s8PdNH44VTV/sY+6rorKP7UxtSdGM2hm9dnPGZ/66ha209F
89jp2oGX9wqSI2EO8FbS4bNNPirxLMp4F/9s8pMj2dUQYVljx7rU3EsMG+d3wV27
lqJwUv73MO145kem1/JLUE8GBkhccvu6bdJ/z8rWlgV9IUrKOBhjPsUyhNiPtZX4
ycnpBuMmJx6lKsFeSzl85YS22/ezCKcvo+yCmWnso3uIOmrSCxw7KOrhpZAz+nR2
X9P6BjSjGpIztEdpAuzLaSKVaP5+sYNIGLgRzTYRbDBWooLQlXNcHHMpoQ/VqvSa
YsAjkAfqfVgHSSfuLWVOkrKl7/J3hnFWa9SQhMWns8U3NwXYXYkye8iku9Flh87p
YIqyOWbvG7eeQ058k7oEwGGBerl9v6KS03Zi/L3kXL/f5xM8yRNQ6Gi8SAz+fknK
Y/9tQCXW11sxZBjSqmk7w8ZtQsPpLZpcWXXGhlqjUQYKDgKiWyarBGiZxUpTOOYI
5EeVd8geqTxPKq7IWC9gQyLR3r82svmumCtL2E1vBjpaMQv+VvkBVHzqQ1u7wWAM
7e48CwHr0GuptsbVEZzCdWfnErwSuiJ+4tuBRvfweIBW+ZmM2OX1r89SqDh/j5Ee
Iqo1JsTy8mrbptKUvCMxOye7Wefto4vjpwh2/DCNBAo3O6L2KcRq4WCspRE9aNRy
CVhswUcGA1KlYbHcz8iq86qOlS5JyroFYpUhAv1aTSwr0EdAx1v52NXDCV6pEAFF
MZeg2i26dp5gnWPvXkbUv4W7koyPzNYayJatFPlUy1IqN5jhnl0Yhosyg1of12XM
+FJcnBP5dsJiX8o290xliYX9QWJWxpmb1/IUWjMKpplaJCvxeALWDQyRBPSWch1M
2JqRj3/7Vj62hyVgwJ6njZ0LJPkZTVvCzA4ufNtz3hEoGs725Wgf0b3BkhdrfBvG
ft3QIGhT341mKpblIazou1nMBB7/jveubedNvsi62Ke9pXLEq9Id/JZFcLk+vgyQ
QJAaqVSdYSw3FLM8Z3tIfzLEPuv693iftisDqyjp8yRhet2ZxfL+xxYdigFztbbu
ATGai2ojnLxCSztB35Xa0piP4Q5RiFpA+UuXvbbx61KbOpo8eJcMh/dF/jI5j7t+
d0CJUW9iE+mjPchcPwV9AokC3IHlLGShCNCliEJRtPSUIu+YVIuE+yCvfR3ntCHY
N4Ww66WRtimyhDGGJVug/O5/aPYuHRHXrKu5DYHC5j8L7kd2gs5IUKdAphYTchHY
9VI5zKxS7kIfqiPt7H4UdJyLd79A9K/xH75ug9GB2xHS6vcy3BZS3zvXg6j3seO0
RqHp4/F4jigzQTquV1w82Igmf1areYykeFANHkHTPf6WtD2AZH3bHnv7U9+pjTUH
+sxHm+tsZa9kBvf/jAZ4IW2PezmpEg2KUBnTPWWwaXjeJEXN3W7dSYrWP8zL2ONT
u58j05XJQF2h3nXV8BOKIgCTV+y1Ii5Q+RnA+eQ9JS8wZgIp7TshTkAMYLGmvVc7
LI7g2+YK86PBlBIMiicosJwori9Vf0uqD5A/S2jwBJRDpWWyWoWxuBxGjVglPn8v
YWJCdtCRSyV7cFoblogaXpp5sif3e4O0VOJifABupu/aTmCT5u5fkXp6uJrD+pXl
8JDUNkDUxjb54ATXMgLWThDyFlkgq2zwHQqROoDnYayb6kwJL1CktfhNeCE48xSW
qROpaJ4J9XjLVzZja/21LjLNmO8qE6UaodGGWZ+fsD2qzCbCycZuDvsrhCWlV271
0T5/tAR3RLzThNJWSw1Aa4C5KRMuhjQc6qFL72FC0/gd2qeMsaN+axM9xiwHIXGh
VpNvspyWRRAq6kArR9dc8Z4oE+wfTRv268R70MaVP53h8i2ahxXc6KyDmsG17yLs
eW1NTdSCA3wDkbKhg/0BdFabzO9dy6ZDFhtivriWnTRnAe/L3mhocv9Ysw+eaZbb
TkAeVzYAV5VftrhsiIb3DeqcEIPUJUm9A1dObHHETgaTZuTCxLMLwPTIpi7jcDds
Kks2N+0C9dk/GsAgwGVAgTjh/S4arOzOXSVBkt6JIzGs1UxKNqeKIQ5nHjZEZ9cV
BweC1IYkPgFeZW+BSaZi7xL1fbq77KWTq2fAXxNHghM/dNmw95PNeObtrfNw6Iof
BlNAUxK7Yu73MXwCQpZSKK2NkjiA2/cuXllC98rlltp+mASiMjbtWhLegNvgYdYN
J8nVM1Fl8PhOpTynK6FRS+d5GfJgNL8uxut3aERh4IhwLJt0y8yYaZPyQ7drctPV
nPnjHq7AoGKg94LEdCG1RMmZmyBREqvuxxRVXvaouRHQ2zoHN1LixDm5gug3BpqL
uqeor4PKfCAgh92HA/lzIm4Fzyirk0RnLVv2Wni/T01LxVqDL8G7HVo8pv7GrC5n
NwMLbSNkbdBsmZuyBNWPZqYbrNNn2GKb/8exQ3kcpnCVPYe9aB3IIQiOfORnOc/D
0ndmAmIe+h88AsZJPrJoitUlDQbohK7wehOPgp74pcnt+a59SmM/VrazWG5QnTKe
40dzc7elLBP3W1cqfuz+UHTvb3iwl5KKDXW5TVXHvfeXyo6O95T78Rlx14DazYXr
KarSIBVzyoYJoKYQdr7Vr2fNsTlgsEN9MYBkGJMcMnxMOWtgOOFMd1Pl5vF4EXir
xvoxD98iPgHCl9KTgJmwTbW1wUEj854/VYygDVlDv0J5/vMnq12e5eoxNLdNa3A6
vQk7cACGsVLK2/f/KJ19nG3djrHFMjxhvpIOgnYMMFjkQO2OnjDbRFTs6aWIO9Dy
ooqUzGTWiOUy0MZLC99GjXa0AAp5CL3p6wkkn+swxmTnSzsd4NX5pFlRk/TBNQJL
qWjLfG5LA9e/sRoc+JmOYLM891KjBt0ElkGX0S0yu0vZYRNsafR3hTP1QS/jCXox
nWXUq5sLdzFP9GzYCYp3nj4ZePa2JXI8jxwD/fPf80XdOPGM0Cp3GbYwJM/SNhyZ
BF2HhAM0Fc7Bc229ISeuvttPFsw/IR1wF++zIZ/f0lXSH/a0B41hlLyVZZtZ3B6W
HB4u2kYxDVilMAqdP6men6TpoSoAFDoG0w94RR4+NGXig9y6DiTP+f9E8h8NYVjL
a1clhMaG0OvNtoFEDb9vO0CEw2YJymCicmC6/Lx9TIvOkj8i5I0sgIpyl078BHkZ
Ntsonz+QgT8Rka7MCBpdz11l8P+lkT6FxXJ1uZuXDto3enyz00IjgwQ3bIbk4TOL
0Nzg0m+EKnkuR69k0ZvkoNFguovTU5Ag59/XCVmmGcwNtqRTY/WVUxH1YRMU4kV2
Z+RS4tmy3rX9HhPms3P0xLrar8TMf+3KRN4WDOhNrVKibssDbiFYmpqyqq8ClbcE
VHz7gxiV8fYInaHTteNHS1hdfFUFD+0+iNwA36IkhQwu4EUXwgE4Sm3eDcvbpBHp
SfNvIJNfowdb5YQYOJAyARLkfkN5j3gupgOKvfBrdoXvTMa2dWf2Lw+T8+KPjFsO
w/o1ePi5S+/3WbxNmjvDOp6T3yRO8VnTAYAvpgmy9RMHiRjxsx+7pXNJS6En/GPH
OpQjbe6kak9Lln7UIuc5ch0WJ1e/JCeUjfrZcx6j63pB4qRVx46PbshAnzl03rnG
Uq9elFBDwi17VHadwaikfG/rQpPCvEmCt3YoN8h4YV1Tv3PvL4eDTwWrlG5DQBfb
GwglflCq4e301Do9YqbdaQxNxMAgpR94mcHfJDJFd4tLaWlFKFQR7s6/d+yKCLvT
SWoNA7NypzqKgAZ9JXZrRqFkTgXoHL7X7D9uBwdPP3imKCA4DLRpyjmWGjxkdBDX
op5vUYLdPP4jf6avJrUhL1jplmm6z+GdbOmAgp+43TxT2q8gtO+MzGq9vPamhXrQ
1SZ4SxpOI6ayGE0S2qJGhVULnW+JgJwhvkak3y8l4VvWG6Z5upR3wzoYvdFViJiM
raIyYcnWN7nyvjIXZThlakenG8v6VtACOCpeL4IfMGnnRgw6gkbkhC2286p3RWhg
jyDagccWWH6X7v+nYGyjgPDNOkq+rcvYWnB0O/foT6oNlP3drH+MwWM1rWIobUHn
6OUBDl+lbuwL3/Hdc6cuPGPxArgwkldFW8BKZvRUuE4pXKYA03Ogr9L6ghPqZSm9
3ZLfc3SorXfd6dGMVPg3VyzYK1F8tAKM5JPIhKmzvmvPgC7wMaTyPqzITOI0Px2t
kqe81T/5MXaXpHZLHqUgyqnM61yHhc+hqclmJLSk3QEJh++ySsGS4/8GXnD1Jtif
jOGLf5mN9CSNuQfXn91uaKb1bxLN/AR0gSDchJ8TA7bh4BobegP5K6cC9sPwD/d+
64TQiuyv28/GfMlTiAkbYDeqXD081kvfwVjeDrU8u9dvf8zI+UM6Jp4r8Wy8d7Db
cpN/IcVRDHYI6cBMY5QTnEvQaxOu18S8kjZLId7WtQkRK4jUgVa/1uUwCyDpixjM
2FMO8weq3uCkXtI4wUYzK0VOzAhBzlGp94PYdM0PlefuCnWkPUgNxXPEkFGgnldJ
DI/Fpu59pFza9/XJybHbz+0/upBm8si4YQtKF8DN6ujbQxyvNoO8ZB9C0h4Bk3GE
9bCagyStS3lQnRs/95DpbdNbovyGnaKvEKHRjZGrxboQSHIxv9pujySVRriR4hRG
ImSVPGJdguOoYFCoCIrTeWKvKtp3GodQ8/tNt5HS0mcM7es82LVDn6TB9l0TJ2fm
uy2XMap0OW4dmkkWxtv6s1yXNBwhzorhaRI6CEVDnBekr8FCDKK5owgPj8eZl/1o
r9qxR26EExE4FHsyI76zvBJWp1k9rzHyVE2aSb9+eaFTZrK3hRNwS5x7HUOWZ9n6
6ex4ucUqdS6AyBdCIbQiiWmHMufp2MiZQ8+hxld/hQvibaoXbjWyJPqfzC51GxDx
9+uJ6l7jba7aoaHMrwY30lE+K8yZUNYv5bTlt57kYQoN2Ch2DKvsHevEUBIIK9l5
ZQ32/Rygwx84x+uvA3EawpxV73HGI8nwuxZwL7gajvEytO56giG6T0DcX67Khffj
CF08V/+v3jNh7ZU4MQlSrt8x4Tki24wZbiWdGW+kuDtYz65x0YibCioK/Ux8Amxk
m2OOgoLY7RQxwGz3UWaj3ESt3VuQbOZBLyBWprkEL8bmiOAWxN/Uka4/NqEa0e6F
i0OmT+QYx1TrrPAJxJDzknmiZ9wSbk3QeF8GzQQsQUcAxmdYg5YziS7GmZbErLe0
Bj7g9WwVm4iznJxk7Dmb1UdKIKENBXguxHzLvJyRe1krlAvYJBPagSjDoDkqTU9J
T4v6GViU9u6hWXy3f2KEAw+eDiAzYRCdzfq4zv3hDaFfJzXwGuttXIKUjgCzwzux
MPqZnPqQ9fKhVWlSZJDzdTCtgEnYDNStRimVdznJ2hZUSF1JSG088DzN5ORcaYM1
Em5JtdKykIITHesH3/5ihkYmMJHB/MWwcxBkssNCod0evMQd0hxgOGtx//cQlew+
XXFqMI7kvqpiI1zZamh+2n1BKUpnKh4mtP44TJIft3rvq2EJtBY/Rj917j/Wlbe1
BiD738wQPBAo97v0IU+J4a+eZ00IxmuKIfdXWoPDR9dc95BDqThoriK6vOcLiZ9U
uUAkKTX5ntRKq2oe0HetsKiME9ma/uVgMhlolXiccY33Gv8xMszWZNi+fes9xa+J
vuKtgpHmZWqiJ1QruYo4oMfO9wh1EYDE1bj+LQbOqYmBw9KarVajTaf8ASmCpMPk
A8HsYLp4agu6E/ObJwzVXr+lG2ObFfoPQRcaMz+MqBLCLUcZfP0N4Gs7lPIT1TPQ
aYmhShvxjrzv8n/aYTY9upWJttQmhVVsLKgOXyYeO81rFaYkHyCe7uDj+EvZPssU
2391V9+wNBd65D32h0nGbPAQmPzMYFecp/7ctJAiHXQWQyIXnhFa4yq8QS83Iu1n
yDUdEVFn3Eur4gxuNZhGENWvCvwrDBM/HeiyK/ICb2wJRZ6bsWja/eQrDTvCKpkR
DmObZSDcxnj0gHcs8ddy5nfN+PjEBkOUbgaIaWKgfgMMqguA5X378O8O3OeUAuM7
Bhvb7vYojI1QzdCJKwXNjVFpn6cL6iZdaUIiUiC5j0r08KpEsLpOMVTLEfRvbp2z
cCC8BZMseWGmaoDEr/ltNf7Ajk7OIxMNIbkekw6Ho1PyFIjDjRYESL0h10f5LYd4
LNyRALYbsYF8lt4mC7g9FSQBVPWnXy76qwn4LLDqKv8hd/IbL3sLqMbPtCPUvNrd
A0/nZjmTGWR/DgMqHSuU89fO5E4rIAU3yw1Z0LpB56LrXsUUrqdvKASWj3Tq8CcW
yteehQhP0fLbwXJvOAX3OIB1eHK56hpHtfKJaCI3wJuDP4XWSIV2/gpJKRA/z4C3
9Yzs/bhZias8x1QfuzRrL7e7xWkVG8ZjUO8tn2R4NyJOPOyH055AQGyRWGVckRwI
9JxyIFLlZ7OhwpYA841HfcqmlNYVykn9te1KC5lk9SqWpYhlW5lYISjGJnMTvP3n
A2P9soga/dKCd0z/gzAdlnganTMjTMDU8TJ0pGCVXC/10wX7CU+MYZ540E67XrwX
CDUwZ1GyHbSup3F6fsTL9w1iW93ardfx49YR7wZCD9tHp13qWzEvrC40I9Fn6CHF
drLo+CoHiWNisAsAWQNz+c5Fr3s+UseckwxrlhUqdjsduMiCQ0uHeJXmyOqQqell
TI9jcQjh6OC30vw9k63zgCf+DLr5iDAXZOCAkQGrQxGf2+frCOktE+18huAN4d7a
ofyoadVpww15VoRm3bGCaST/F64eTmb3b17+BT0mMMolh/ieKJdgIFzrqHpehgkm
uyZRuFWaVwvHzWueip5Ve6NOBK2k6Q1pS112nyrtEHGu69RDazWB60rmYk4fFQ7A
J7n4mw+/xHSo2wJjcRv9gqfT9VCMwgKl9yw+8lNPsFIw8J6aOPZlUDP81+SYbCKp
J2xGkI8W6LVQTTtiLqt3/4BYu9ihaWsjTxkURQV6njfIfCsoJuFz5gLfM13rqlyq
NvKo+GAIFtb7tFa7TZGuf9dLdoeJBQcf09hJipb94e1ytjUXuW8rtywgIzANXwrl
GPs6odlXEzTqrgnWxskLLeRhW8EFElx+iw6YdO0p+1DNfPIoMsgcSooiSusDFXFb
ykMK0KhDehpL1FcoTXO9dYGNYHYmAU8Zme8sstKKbWIHwspJoTlc1E96l0D/ZmWv
/6qGXLKDMiGdTOayuRyAKNonn8xTH7Jq30v9NPLahEaKPmgWB9mEcMKOldaBFDES
Zwpa0QinHO6I8inwCA6sSPkSMLZoVL/HcY1xKyQvP1giIAf84kXKb1ZOmNU+OLPw
q4jD2pt7j/8wxiOw8otndwmRPv28h9PFQ+mFgwIzDO3/xHokR69TXzK3hhvpZ4If
rgXiR+d+fpVxVFBZvNBrVbwhtTykAhurlQyEBzlnlTzj4EwXr2ekI5/iyERNplSA
JgZ7k+juYIhKGRatOrP0zmWp+a4Y1qLehcab/tuF95SNDauR6fbwhIazLr5yr2uk
qJjGj6bIp9maLV+ndYbnWGfn8SNY1MFbIHYg+vIpU3LN9mHrXNNcgQoMt3EXhiju
2igXACzq1+mhqK9STRukdj0gXtX6AghZ8UTYX9WMWvP3Y2RcY46osXR5GKUjHUwb
ZJGSl1Vq1hUjPGvZpe+64il3TT+uiLB4Og+7miwV8gqwOykAFy6T/6MDIAbvzG/Y
5sUuWEdGLMB7M7DBlb426Z3RT+nNXdNF1STrgwOkjGJ5XW730hGAi6BHejjyog06
iu4R6sUoWdsjnvINeGKSr+FYbnDpDPVETP4tSa1h/Ur6zs+77EYdzE0MBcJPZ0Ms
l/gR0CdF4u5uYb03eiUz0bI1xwfmEU43y2Ja4fhZe8Wa3qv/+EQwvdok+7QXXcPR
vtIo52eldAg67JaGoOWftufS2T4ZzEHfpuzCPFjcqJ3adhv6g+guYXeynzafUk9T
HIro++FNYZ6kW+SFSzYCC2KJx3lFKVbnx+DAaYCJorM2kHOSUnat0fGZpCwrQ+y/
ME2qWCIXE5fty3d6LWBBN2Sc93Bd96sxTGIOyY63Ixk203gnMVEfUAf2wBjT2j8A
lNNtaZzhKdxrEkgQJCiV2WR+GBWgh4LOBMrAkWgT5Vv+5nY3HNQurA57xccnJj3H
VS/9otzjnKydUifWoDG75y/WDRoRDTb5rLMs4c3/39haY+vTmzO7JURdoh7s8XW5
lxM1pJvUd6VGsZnz2VwpbtwPYwQtv5rlmvdJsW1OeQ/8YTPgv2H0snRR6WdCItgR
FmMMvLfNXltsq5hGZvihbcFL/zCHFwA2A4Tp8jvR0ENht90ty8VnPGNRPElWuegv
b2azOisGpZWaPTRr8jdBo3NAaM5SwQYAT59vwBw6zcPcVa6AnUoX2zOEvGeFx5Rk
/ciFfYXmW4coHv8UrhRA1N42CGrQKPXL64NwJI7Y1DAZbA9ZG02+0WrD7QmiiR+U
HRreQGNz1AUp0cF+R6PYHa/yjvNxiYLflPe8sVmGpczO3kfCnL9qp0FV5iCU36Gi
zI8AwEKPxBUDVoNMid6djr2mUWdydo3AZ0f/heNPtwfUzFhxwkLA+HE3+qFlOz1k
4xWeI3qw+GJNmfpOT+24iEllUr/kokuW9NHkrZo4RrPyxqSntjE2nBnDXjszM997
vVbsO86Hc5IjrWm7WvVtZSWPsOv03ak6lOOesjTILYAP4CelleogniaOqzEyD41I
JE2IeRKXobfLQALHjJXvEpUGXFs75kSdMbP6wWGyQwF/xXaIrHdD773YBsWTc0Tt
GA9/Vs3FCDuX2xNmDZBdBWQyrQFrCSXAfiICsWMmSqdDNAlYSnB1I2ftx5mNcdNF
sqp25x981u2fkmPqzyiW6qbBTY+tSjyzLCvmV4OrXA1n123QQ2HR7utDCJHM/qjS
QVggd36015bQnmhh1+AG0QfIoJ6/apG69LABlHGGwBKoAZUzcL84aCzQURwqRCbp
da8aBMu6iwDTH4xe6/8qKwCcszQBj4G4GgXpYzUmTQWrP/brkhC1GmZ4Os7WQtca
ljlD8q3vor0+MvTIj7tiG40I+2GYDFnQMsrkEu9fB6Riod7456f/jvWE3bI/YvMY
eRQF/bM66TuxrwOL8+DROp5f/17/D6M9uQm5j3zvJv9PLbKyBztPBn6ql8vDH0GM
GLn0zDyhTAfDyg8rsJVie5Dq7GwpnbaDelx1fo2hFWB9RdwWlXpQwJMA6CzPB8uT
t52WKR0JKeChiGs5GJyKjuYZV4c6XjvtmQL8DtglqQYnbsQEFOeYEvr8O1oMH9I2
7uP3IQRkThOFaCOVpMbqctCuL4+ZDw7+sVqMJLEUyUJ7MyJyGaKOeJBAPYYoaQ3y
InQokprxvYeCSi22cOfANrMleJCv5qlQyLbgnMocrzOWuPPJU8NsRJkn7kcGHKYv
QBmrBZvg0UoKBsGVpKJ31zHv+aXj77PZZgdSdeLPiu3cPALJVjN6RHZw0JZSSssu
ZD3YP3Hb/5no4CykJIHytRH4mJ752G6EvIVxFE2v8iXZJ+fSeZFm9RpnNv/kxGW6
KpL7Vg5iSaStqof9vnsZwZ58GSnR+xKcHkrn/5GPBwSzfqTFqgG6QarDhtOGrA5W
+jKvC+hUpCoyviWLFPdMknxdY8RrlLPy11PZk065DgGpWRGWZOsFuZiISyVjsFTC
1dyIREzaJ8W1BB2CHDIFnKWNqzx6HX78qKUxHYrn8SAQmo9CetJLCwmlK6/ZqHHU
AcPtsRsMX5VwAHuM5ENmcAl9sdVCKe6RmGVq5MSsP3ZllB3NF102m6FTfk80Q9pV
HWGoeX74AhLwN+2j7+KmII3jLktCq1mt9b7aLxFSIzTaSd5p4WGjUIlXmvRdyeWl
ACB3zLrAfJ1Y9ITgeYrMFyd6fTChOczLjpTLPAUNH51+KStLx1EXrMELdFxs0Qjy
uiMJwmJgidRhmUbfGm7J4iklXxYI3FQo2nujHyKLhh1lzPZww1OXBqxmHsNTWnK7
L2LZCXyRJymkxF9C8Gj2yrXvn7I4IZNtn5LDmyFC9UY4U09F35DTsdY4svN1r/F4
xPz//1NxXNOhNxpORdxhWG4Xy+hMK2uKfiA4ARkHVWYdbzjFtes5YwNMIlp2yHlZ
7lgHgtaeBiGXdrPCU8yzlab/NhPpngz6T0piYIBAS+4ZYoYmH5mVon8zEyHpjpMB
hW8pFxoPyfDUFQb+MV42zWJNnUy4/8of4pTFemgMo9oeRjOXhhQxnrfm83jcbpmJ
GcTOyiIIIKxcWfWFn5cJ5QSRE/3ujSFEQ652+wDtjWOEo5bZ3zrVdXF/t6Rk9xeo
d2BicezStZJntVLqx6upu4zTNQ69kIgPbgSRZxBfDwm9ph4LOVJ6qE54n9Aftrgm
d3gvk+qLfGIgz5xgaFJQJq1kwzFI78JPU7/kMpALHOk8O/nLL9TrBZAW3QHE7c/f
+e+SG8qx3NOKlPVY5ZBZJ1Yv43keLeuGYmC+rGCgqrF8FQqoC/ZKl+DrV07jT/2g
5QcZ/kyITRC5KHTEe2EK4X7gQtS4/iH5qcFeldKAeTErn6qqM4dEfyN+qRKWkD7c
MYJw6hUYN+nQVKxToBCaD7dAI4oWnzNhLfjgCzwaII8HFFygRGY+Mqz6eiMV8PGo
Kv0O38Bwy8iEI9mV/2kbNyXmvBq8kx3WxiOVBKws9vNozdLfqlbz64pecF8oIWos
5TOhwncAAzNBL09kjGM/dT49frJwPpIqGp4K4IcROpz53XWUwlb4e8RydUxfXI7m
scUmxtWu+FOjfEwwnJYNyN+Jl+nVtoEdCQnrSQ9WZbTC3Yuge9Ga9tm3goPli8mc
UeKQdI/FRKafFI6GkUiVvBXXwS7wmiag39EGbt8PRfZpdBztnu1MTZOTE/4UKOed
ko2pvbjxTKNXmKbpEqid5A7Un9e/nllpmgewzdSaen9aWC03wtmgDDGJNZ2OPSHd
qs3ry/poDyFWcmJTrloed8W14/pO+p83HNLCdm799hENO/9gNpUq/8HRilJTnzKl
WWBYEYcHo+EcHLaSrF496fz2EGYubGdoe2+fegx5iv1gMg3OyJHaLfnHqcl4XiO+
47gu4m0IEUux+QNiSEAoRH9EUzQ1k/u56ug3GQBlFPBmaZ48b/nB2nd2yyUGeguf
m2MYLV1dbQ7+lo/+GOZXVs7/om7BQOHBKGiQM+6FmFXRgj+yvBjnTsMNiPmvwzkr
hTIMIp89zdGy3el3NmWooMbqD7TPwTU3gzb0Y1uZfyrqa7UR9KQQaJ8xh/qolAzR
CgROgWRk1MpDXuydSi3cuLWcbHDLSbLnFqUzjKhfu/2QdDZ9IONdxdTuwKl5Rq8W
7ZLAOpWIVBo2ToQea9/9hFcwNnZ2LSmtG55fTTgHB2MxQzOpPDSOlTNEiyopHPDn
JrirhNjSnhhn35J6gEcGzggihbIqjCQF53dFAfaLGiMl9eGFNCjo9noHT9Ayxsff
P64ltAKGF2tBI5wdIXtsKvqJjQcyhkHwMa3ulb2JP+7lGuljEA6e/R580UoXxG55
ZEEqR9ojvUzb9ToXq5rr7U0AVkzooVyESYfhNWOdCpy9/6goRex1a9w/F+T2fQQl
+JYeiPZDCGyNQkE22Uf7XkDo8Pz0bA05S22q246DWBmuJhaCh3Fg9XI9lCTOZ3JP
RfmNX+jo+m80Efi2Tj1fvFnfuLsfg9cGWyugWTaCW/WXWWYCbYtkaEBfSnjtd97R
4LWSmIyj3UPfpkEgejSwUAZJcHdD3IOVpwkVDJUc7sT63G7Q4PDZNXTpqt7OTm0Y
T0vT0fUia67iVvCJVr6AVTRyyDtS0sulvucWMCYk9kY/1w/orbHxs5VcVTknSRSB
xBpvHBLK5CYHBNRU8r60ar4kLFBK628MfOEUSR61rX+9c6s37OmMyDHrIBZM+sWe
8RPYWdZxSgmCwIAuGpATt5K91ayUFkFiGBRHk99tt+AxCnNABhSgSlK45VHBtRYz
xvKrHQVFZfER/G6uhsvTOusIfw28mnjqv+Wf/bdcCVMCvvkqpdQsbf1Oh7mXXi92
phgDF0Qeig+dFnb5mi2RoA084YlruP1NTlU2PM01LBS9BNMUri9ionqCYGaEaJo0
qoruKXn7hfTQlKGumwcojhNyCrhas0C/94T+J3imW0oIsSPayg0boeDGpJsl+wEX
zsnzlGYrBSZNBrWumLEkwOuzF3zGRKFNoFtaBHZpgknD7q6ZndQlIT8hyfItv4av
yqZOoNYvORndAlxZfA0b3OQGgtEhH1q9qrQQBJOvRn04oXnNMo297E+vmJLlLgp4
RZeLHFlVUCp/fHa62oOdLexFTYHyCgN+SgSt59/nNA1MmFqECyx2c2zFN1lXhq0U
IyzpEBg5X8uBVF17mxBUh34fULMh6c0EEj1kkcMyoheGV++2MofkDygY8I7Mwy97
mjow4HnZTIbaCEuol3Jkj2rPIDFkdhSPf3YM/CKaG96zTqVqFcHLhHdZkMJ4chzf
qeD6aF2jygOXKW94pts2NgB8sP15/QXFy8D5olidpfUdzfexI8Frudk2/wJ4d3Ok
5d7HkH6iJWNJE3LgyI5DA9xEQhJ2n2XeMPB5UG9e3kkpFcJ3jf7w9tU0pKzn4OeY
2L/Im9VqEXVGOH3kd9sQuytoHT+suwx3cqXZtCcLtc9kLQBpHlKM/1RukJhcehHW
x49+rqaYBQo8ypJEJylALsVwoFvoDK9URVHXRw/hp2JMEAaGPOT1TPeU1nsv8nSg
cl+7Hfr/EL21eAu9QyBi7nZsxNnFFzQO0XtpK3FgDjfX72nN6+UWjHaLCHTjkMdy
+9sjL2oGW4e1dsWNYGoJFCoesIwgHNzW0qYHuvDuLGGIS+jmQE+1X6f+5AWfTpVO
6E+pvLq8/Ohra2Q4hGIygXrfs8F0owjJ+/1ywnMFndSA83Il16vor/shfyvz7eO1
FkaNYaQmMKNDdRJVAUe0Jvc85SBu76ERVnQOOH8vdYEovlp7TuqXVVRKJGcie459
/CW82GGYG12JBLwrBfmr4mKtVmR/MtHoqsCkz2dip0zi3F2blSA3g42QbRah6Zuy
KWhykvy+vSQSuXoFaosaHUh8LXcHeLVv4OCWOKdg/Rvd/6E0dmNU5q5qlr83dvbI
DCagI+qJ+Y4dP9C5L54MYfOFgXqd6l/Zra2G9+0byn5Geo1Za8MRc4DCdxvBVJkW
yNZXeKHNUJeFSo8fE/qiNjTFYsnOwvvmiQbxawFDaB/UqwiffexqfZyinIDgG3Ft
zvg9KUfzBM5vnwNcEaj90XqqwO67SA+cPtGrZvbLqRkzvHeLVFHZ9afrnP3yLlzz
eQjg8PqSKj8pCpU89R0xhA421Uvm1NpxXjDoQ/MgrCDKpw7kCznLdGyr2a5VlhzM
hC6RXMH9LaXny4HNNxGiM428+hjFXA8krHxX0ORGRwCGqXjdSNHQxpacWBuH2UfI
Y07gTNs5UraNJksJLndqlNdQkZ4Z2ioO07yhP2v0aE+yfaML3v1wfo49ULaZHFoK
BzfOBoU+nCIP7y31J+uqFbs7cAQPNsMTQT9pMC7y4rzLxpqccbu35JhiE67Sivio
oHkzMYF14OwhIbWq7LEHNuL3ck0PhbLmk3qc2pXs/DDYwdGedWCHZ/vebo62U7cA
jjtmWP+0RDAXbSGio5ZI2eSqkWVpDLuKA9xsZXi7u0+qFPEJJL0k6Vn/Lx2sZibo
ZDYuUPfbwV+1p3We+byh6utgqPE3ufST7rlSgvRT/WURhpgYzh4tUn4IHkwNIglB
JoWjbV4YQUzDq9WdB2aFEM2YfprU9+bhCZzN0jzZX1fUF+Yh8iHAS4Dnp+PqCEjy
09dCbyFayxrm8taYFpl1sDB+1iybCni3Mzj8xishByDuNsAbh2Djv+emzO5lf7MK
DSM+CdHgcuvHifXUN+AhiwB8yTWIjwLykOnBQa9FLGpkRNmqnJ62SKjVwHbZrwI0
CswnsygZXQvxzq6X7Acq5Wdjt99nuEFBgX2SBY4Z6+rfKwzg8ZALjCqUkhnp3WjU
TfZ9mFuToxTXgOIynO1bAwNX5YkSMXSm+ic1wlGtctplVR/ks8pKUA/SiKCRSGIi
R655goswvssGtMvCrKbhrw8/WwiTJAwIQZZEWQMqAVALTKtXoFdnwdt3BY/BAaNo
kenj3hFOCsA11RqVkk8p94DidHb/5UbHXR4/utfq+XOl5hcNVonHWE/ujUMFMPN0
jiL5SsUfJiIbGKzq6/Yq6cdNI8/+7e/AdJIxgK9Zkr/pVL3+4+2oSbuEklEmcEsQ
wi0iOzOyc8o/yoGSSqsOefMqG3x9Nx0+C7wUtjZ1ZhuvYIU0hzKrImfarAwn8pAi
EBSPCi7eqwNfnMtIw9OX8eYPAFDhfYHV3gKE/EL9uyfCErHxoD+ja6lIDt89Q1ZO
SNLKjgwWvBA4OYmEZ7qMGbtLW5M9eyQMj9Nl9IMAgcPO/CJMwhFjRALX+Wf0Suvv
0zOnqWRkDVDusEdzAUBxYe26OvIuib8ufaANaksqPiNVSjSn1g/VuVdAoN6URwHg
nw0zvHzcoL49aVLUHbhdnzg8EclWvRVL7KVug+Ggg8gCHOWQxVvqeXV3f8Sl2Nlb
B6JVwiemzdqYRXzPstqB1xHv3I90oxUP0zFRaJSz8bv3g19y4Wg4YTFNJLypCxi7
nG1MQ6w6KnAaXxm63FQCQHV4eVqEdDgoEk8LLvxYT3mfXmdnJ681nmPZwLuw8H7d
aJu9O5lXAwIYuiGz25EXM9MwuFa3YwGufbgKPCRPrazdsKqSvB4145S3yDyYxO9s
TI8WPIauCvULOlA9UKX/XSbyeTc5zkKtJ5wFWJhLOcpWsQihRV+V/CipgSrBE0Zv
a1cD/6RVj4jfZRtTFR5ZL6lDz0aSQZqms0OYaR1/nc+9zK6/OacufCG8HE5mwRw9
4d2YQf3Gb+cye1IxB+ilPJd5d/rx2AgAae2XZnROf3GXkM48UIQJK6IyBz+8lr3h
qTktLed8XD2MM9fba1Wi4OlWXwMU+i4bmNPU312/0RNPvGDyothsi3D46Xr9bsCg
EV4xW+gR7ieRtd/MXO5EoXyH59/du296fRuWO//5y3h3Lr6785ypISPVjQ6QMkZe
XMMjlUj3OPtez5tvQfc8PzjKlN9p5vlX9wvpLKSOgv8TtFVnttG7WhOPD3n+Otcv
NIyZTRp3rpA/LtsET/lILbboAexaojaTEc29Yc2Mrd95/UyRkfSVjSljq7O78G/q
RuYqCwGZSBajSr9EdJvnFC/ZXzTNj2aEaBbt9IsfKbk7nRacKxhOqVjh1tgh6xlp
eYxrHZ4NhAHl/RvlzJ2cyCokkC8RcdYR06xnGrgM6K+vXTiBszZOkP8Vp85cFDqk
lqQ1WJZKq5lzKQw8/fJLsZBR+1yYAKT+3BVUrWp+gSFgi7Rjor4E8KnHjkrOtBeH
hD3APSKaKRej3oayPakv5x2up8sX8qEQySdaDbCWMtUO5Nsw/Mg639i3CT4OgL9/
cM4mhtKDhect5t3PTpG9rA/J5kk5V2byQOhuzOjXnxPEtEEtGPzl/2KT6ZBkEVg+
+wGBpEeTLyF8OYLufBf5XiXRvd1fHe5Krwkz2AH/AP9iTIMN5/cj6mK5HGdxaRDf
RkKi1zZnpBoeboYwljZK4tUAS4kxECmVZC+S/jBum2D2SPLH5bRxc2DLoI2yxzoG
8h5rKh7YsPIPEu32bTsR1X3xs+sq3h06L3WDwoZiyRtLtsEwxMiUxukCzifDK1aY
Oux6SdNinucLBZV137/u6kiSNIyqu+YmDAKPZJxIyMa1o0lkBq5OvNaKh0mQBoux
e+IG9WW+JZ1glrNqZBSXUkz5VvIKmWPJLbHbbJUFjtBGhXsM3pxvwcWQZAb0UL+B
J7QcZfOIwjp0EWo/FML5sr0AKHHuwdCalhCA1U453TmHDeh497xl3CG4laOL4bni
QutTtAMd6pDVAF1Y9J9zbRYPe36On0OPvLp17LHkEdxQcQzAHLa3yc+ygFfD+mi8
7kkWKF5UbaAnwBNE4p8u1IdGPKUdzW/vfWgo/HT9pU9uBuCXZgC0PM6McJwfpCiv
XvXpcRQM3FT5Ma4qDts05PcMbbYT8EHNv57Fedcn52EWgRf6b7FSdA4aagiuYD9e
MwXE1FppBSZZACBvVwLgX43A5euxL+gKGuyoTuyLkIWTmJeE6icRub+AEIGMXXgD
AgiSaS0aXtcV23VGtLyniKfI24iumi7RAzp8rtIpPQHNGvK1fJ5ai/9yf4d8xncg
msF+XLC8i8n+e00HJI1gw4TPscdAvou8K0upYKv1NQiE8culhzPj2VMr2MPnLvWS
aTXAuEkSqtXym4wdxR1jmk2fPqaeD11AYAYAiKrzYG50+7Cjx06gAozIxL7mtEIv
WmFPzz2sHI0zBXWZjORYHMARFMsaroznN+D7FYjacgBze9swQHRRPZobEwo61GZY
r/B96POddmXPMQE/23IUg86Gn6+dPpbt36ne9UiNMqLQtAoE19r8QkdT/rB5UbEW
d3xEPhVmha92EywKWpVo1imiopsDImexepZWr/WbB8nHO9xxBkbhwNv1OhLhDjMW
/TWp5bOkffVTFkxKvszsQVRbLobfU2OnKLlnfuZo31Ou5PCssQ88tF5Np86RW+qz
c0byD3HKJFwaF1xNmU/2+uKUKaIRtl/kSLzL8+vH68Af7DTU9Xrx6oTszVd++Mbi
2etOT4LSIfu5fyWuo7sN9Sv15vheU5FHTxbj9+/ukiZCwrlAsK9UVtIOGtp63Ioz
nrtp0w6SIUUSh3LHoIA0xqplrO9LUMqgikA3/L3s6wmhdWChtF4BBEakfBXpFMF+
VBsB0GDdwmhvaqHyLYtwYrjjb4dbqdZ66ntCBGuAdPzXhnkUu0kgqOpZfdPWSz+a
Hyf5vsRev+3AkQ5uSdEka+M0+3mNhdIgcmioO368Z17DS0oaPZNuSIHMlBFxXhNi
VlD8Z7GFxHSP4x+RDma1wWEY143eaJd7tFhosDy/MrD2Xfz04qcVk3LZLbTxQOLc
sBGfhsSqouS21rn/HhNieJLUDlVfK9ZKh6GlirbcWe2f/qPQXglaZVPNvIXTeDHf
Sh6Q1+i1FiSEazXqoUSL0DWmyXn3koJKUKzmXEUMS8BQYyNB8lIOt/KWaIjsKYR9
Efm/FXY5dFQKRs61ej93ZQVd6ykPVn9IzQRnGa85zTj9tJNOx8+4+MXFkDAcSxQW
LldawniisCLtaBAUovobKvfa/g1WhoOH0w+AZ1ESsjIZIHC1sWk5HsFbjPNBs/t7
0RgYZ0/dEbWobvkYKQkwF/gUUXIM0zsjH43g/nKvnzOT94feMeoRnNS5YZCmWZlf
FIFWVtD8GvUOT5+NAUVXA79IB1beqXDlrwmoCGefER0ByO79tfJI/Dy7rgn/h0Wz
yMxOfAHZZnB/mfeDWTJgBYCiNaGm7bc8tTHwVvlfPKY3xPhDv9sUTWAbowbrOJCx
MGKDJ4VrgVjCdccUF/B8Sa/X4TwuD9iqqn8dpdQLIEQ7yI9D3CXsBJTr8wcP8fYK
7mqi6iJSs4krPEckqfcQ1cy96W9Jx7l11TBAaGeIaC5U5mwPCVzIVc6qrq1R8lib
jwBGFpS0ocnvXgxIti6+y72E6whjVH2VvKkpnU7MtYz8WC8PjZDG6MHFey24Lcla
95deSfTXPOgqpmZH9pu0CncDby1iTJ27oJwvhQ96W/3Gz9w6k/RJhdSEygKHRd1P
JW1RJL6EWpuCRNCecjBP5IG46md8Ghw3y/DTzf6eMLYlC8/o0mGgXOuh7SB7/Ycg
5rysnEMxRRakw2Nkd0SNJJMbjeQfQq8V3v1Q27fXSjH+GF2Ne4gFIBzkGFdijdh0
2eKEryLauxaEyZSHVWat26qub/CLHml8CtsWNgJ3X15tBI5AmFwCEbbdaxhbr2vE
aUSBsnGRm0wgHfAuiXzhmk+Trj8jFdRmDx8O+Q1gUROrrJukTm4LcZIw8FxShBPB
G5ei15hNJb9nenqWBDnmmYaD0kkZ2LdKjsPBAmQcsmrK6lC7AcyH13cYUaMdW/hV
rybIvhiyxRlm79WF4iaLmZSetcGpRSRrohoiIDvwsEFLKtlLN3/UW2/SRI0Jv6Me
n1u4XZLgU8/ar0kAA06L/2BUAvufTrpIDhWzPvS4xYLRrbHXpBWYXyWO8bfKp6Tl
ChPKjXbZo7BWKya/wibYVuNryQPoKQucA3ZhqyfhUVkSBKC9VbFR+mEtmQ308W+Z
+vGGqlmcVpb5h55cOpcv1SH+7KWylb5qEH/NJ0J/2cBlfrbb4MB5E3uJpkNwTFUq
rxCaCSI/4+8Xl/2Wsc1wFRu+4P0hlXwor030fnt5fw16jn/asQB4XkAZguGL6dog
f5XOQH9K23WXh8HSHoXt/MhEzW+VYb/mzNC027rlu9eCnMZ6MqHi1gorkrsIWbi1
JWWvPXXtqNclMtTfh9keNaSnDZPySINpRnExPQnBMA8TCgCCyjbTpb5UpHCUsPRJ
f+8uYLwOZY2zVDff8EGMIxXsSUdBzDC1M4QZyaK3a1Hcgu1INZKymBUpCXn/fb5Z
+XUEtUyfBrYVwmsxr9wgRToilcXDZGMA0IaqTejg5LJk55NWeDwEzE1PH8G/9qgU
jwjcHX+oiw0pDSQ69Nw6tubHPHxb0LYaglYhTKw6i/60KybHV3ioZLlmT7MAwHzX
72pjzbu1c1CSV4Nz04bT14cvuZD92nZiyVYcpo2NURmLjWDtSrEpIkTiVW7seAlX
RsC9I929WFWrPxdyxcH5ILl4y6WWpuqG4uPwPbbZP1ozSKbbkUGIqh+KieonS5DS
LINn4bzjXpZb20L+Ib3Lh91kMbgFBHKOTtkcPPd0NazP+yJI0T9uuR3n5CSebUfg
82kE18yu2CFd+ujUUnVj7qzOlBCI3xzI4VrQzrizyvrCX1MRYPS/mxQStNrCmaBX
iMgMjbVGBk8muolieIwQg/6CEVxXpFUurl8oFfOhVFMfVOGtEGfAmfZL8Ro+FC13
5njLCF8a1HdFzpV1aRzT8PbyWKLf2pnJ/4h6bcQOIOj53swmh9fNGEjKVM9Je6ox
exelAdR9n1+SQMCCxTf3yStma0if4XevMm4V2+v45FT8kCR8zRZ4Dz/XvlCZwPEj
WVMynX20jAWQ4EIosGEfB5i8d5XWDCY5HLHT3lrf+GlVb0YoGva0zILZZm3KOIhp
thJZr1wvB2BsLLHP/M8svd3CJ59IqnwqTPuRbjK1tH0XR9RC6X3pya8SFZU5oWkX
1h4wfBUAh6fdAu8DBLPWZRtIDJ4Y0MDMI48NNzBdUKS1S2o4XBPJ7b1e9nVVkAX2
65MBxgGus+fd078zbvkM8ojHb3tfElVHQAgEwFGEHuiNuExsH05hzEikT96do4sE
ZItEFRXZsrYoYGhCpfB0KtL+37vX5gSCNxbhfPuQg/FocFDQjhWvXa1mtHNaDo7C
4p+rw7V1yJSUdk+8Yesws6vcoTC12pnNOaJi+Jtb76MeDzXktmfp7EsbaKMtlrLf
fUm6YRk8hFMGrnbUd7tAHpr0fbzMeF7NgY+CmW4Y1T9A1jB/Ymz/XIWZQIjYUqss
GVXP1GjJOUxZ0zefPntiSQaHr5Kq7iGVfNAP1wqyK47LZR+xqq+YcVYBIXBc64tK
LaFG8PvCBLkht2eRwoRuW4WD4dnn2oRlZX4CGQkFxPhs466bwzpl7LN7do4d/Wkp
wmiLP4ryz7WG7NkoNHzJoNEFAMCUy26LK3ZSnIQj6zw5Q5vG6++8IcGenSLE8y4t
9hSVDa+r9cXC0Y7DkQZUIxYBi0/LJqIdIcA6w0oGBttLXjwMXaoWZBltVVOMY0Yy
9jykFDH+aDiHpZXYuboZJhrOqL7Jo4YSfpcBh/FEqiJ/2UJ0+WU/nAyGQccPa0wB
723XzqRVp9or8h9wb5yAYahu8CiJnYAVj6a/NAP/oYUrrb/u936J5+/pb8NYLZp6
hdRGIvILYOuTpyXAcOuVhgR35Ah+mYyH8rTcAyXbZXj28punUAgpxZd5azHDH0ih
38EHms2T2tBH9TW3x1bEa57zkl2VImFfTbUY93GMz69P1ch/YM29f/4dVZrnS2Hh
rF6eTN+38f8NXINGVvhVotGtao63i0qx6dnHpYHEEuINOKMurjZrHABhvgKLNbvQ
BGT3rozA4Tvb1yGyeLPTEQJO5f7KkKx18CmtDi+Q3SqETUbJXuyl5DZIUuDnJ7Z0
NhJCxfvByYfbOyq9k8Hq6ekXuNx2By2uNa1io5Vwgp5MBvclav7xAzeGnsGIlFU+
FqdoYqeYNhW+NGSWlTz5TRMLdbj7ka7XHcBPQvs/bMsbtlkVshOSUMOK/oJ0YDFf
smjhrwFqOhLQhQ0HirNfgdkg95ZRwXrAeCHKvOgukjbO5/e8wEfTbFH11/xEEUGV
pteF7OSTe4V93GOOU8VPRXWG6Aq0K6AYWPqfLWkim8ZxfopZgdB4R0S3NIwfPFAD
2fy85LmGKvk/7i8xiCT6QNc+3u5RvsN45a1Qz3z/1lSg5BaXjk5vIstrRX53t4nj
SYewWvL0+fKNMnyjR94T0f+T6XkWP9j1lf1CWhHsYdOAeWD9+3Z8Rv3AUd/bFlI+
Dsf5R8FG9QLJaJ1M4SmB1M1qT2UHcqlL2tUGMoQ0HllL8Y19GtG7hKENzLkB2r+q
8XKTAEPcwGp0FXKFrBrLq2NnrylkTdGwLcHs32l+9SO1C2+9X70nwefntcZdx1Bo
I0fgKD/B6MVznb0i0viTMPMq5/hUKMWu/KWah5YmZQglpE2V80SpBRPPncCalw8I
X09L/mP5s++3rh2+rfUH2AC9gmmL47zOt4ozgvM081R9rEUkiMF/HGFkVxyS9DUw
YGpYjpjMvKPUGTgOdy3ziivVNxH6eoilLikNGb2EtHgrNKlIWaQ1QNmYjLda/mUJ
XEgMtQjv1o954x97yOFEDNDImxtXBVt4/Apux+qBonDdrEYjfC9ty+c7tQdWzeQK
fYIs1b5xCSsED+TR5eteYP2ysCT+dQhSAffCWsQJVep+O1VELZqZW3TI7ZPkeFo6
9VQ3kTwAUUHfhHI9SoqMGTbgBsZn67Qv6TUVGeHswBkg+7yfFhdHnZvylZFqetUM
AkQIx63vCQtkCmHqVdgfae8FkSFAenmxcYWioMskg/K1jEnpRIVE6mW7jkRAFAGp
P5UrbHbyqhMKe/2dVdLvTd7BFuQaEAOUar3rz1Jfm9SyhT94h5eYiR3ahfy4FcCh
Ofwr2l6DUoDInSwrmr6ryxB74h+o2KGiQjd/I+YvBePQ+esDZDCN7VfPn3XPGLJI
dt+EWM56qWzcI3lU6ndSKI74KMgYB8hssdBTNprJVA5GAYJps0NihdU1s7yMATYF
bNjOSFeZY7iG8R2Ri/r+ZhQdVTuoMosqYooSFsdC2vQqX6Qwm9/tNJC2EzmZ4QUn
C8Q1XiTVuy6EYwNP86CRm+KEWhvoBxJwqx3htDaTff4l3Kbeuv7UMi9635BE6czi
g2maXjhqj89hnstDzh5RupccDVes46VvROSE5cHllpVEAJCuk2VwI3mHVIKwbl6o
kssuKSZb/jKoNrO1Pvhu9uaRXLUhRXQV+eGj64Rqe58VMosByR/S3pwAbZ1NVCJM
/AoBGjxSLIPYatW5x4SreLWXpbEECwecg+1xubimoWPO6kTJnQ6mqG6BmAdaW1Jq
U9nru477wkRGrFeEM+G+owfgo2oa5J2HPZf5sqmYqSo8BIjKEQgRK/B44RgxIgUi
omjGo9HUS0ULx5gJKHyY88Ee/3pGFIdABcWrkGhs/5HtRsmS8R85J60fDvMrPZDT
RQ2tJCpNVtqUzsCrRWG2vhSAfW3GhkFUFv6yYGMIupqyAV1owoj3FOtC8QfcfVuG
eIRvfhOhFi+PXTMbVoIfnMsJONYFI+XEhxNlckaBfuO0Pt14bPf0Dck10Fu9buMw
L+VobjUcWGsESYEMrliMpS/kScosAOTQZ6iqWJf0eFW/Xq/Xy06y7mDwRLX05EUq
HWLL5/pve5z+FjCcbswq6ciVFJKx/9pJvS+04my7FwPoTBi65h09PYTj6Uv074Zc
Q6SW9Gc0oCGyE4yu5jdnbub5Juskwrwk4CKeV4CUprlSf4hIsjSTWv7S/sGXKMRX
WqqepA6bsrX0plhx3Kl/1R8kmpQ0T8az+0wZKd6uLb2rc9g8Hqs7b3dweBJh6Tgx
BxLzd/DpVZtRFpjuaRLzQnwi4563UmB6WcIUp5Tmk8bN/3hKzkI9amb87MD/+suJ
UBHE6IfovaGxxAj+7byzvfNGplX+7Iv1PxQVKIcd6BDVegcvqAqZ0XWf1SI46pvt
ciRSLwGXTpQa6itx0CnYLeLRBwIG+Us13jEq0Ql65QaxxJ/zzeLuB/G407+zQOww
a4X/VN1dbE5okfr6lwsaxw6OFzmmIckpDza0WI8T7G9TgAxCqZNZHklrJlF88jtr
t2tJLkg6NRTgRW1wzXTv0nitHNdDz3O6BPj3KO6Bo2KyrHolerYjaAxoS15bF7Fi
UyHmLU34C2t0pnXewTB4M8eTEbiivbJtXUBJGHej/ekKhkAuaNuNR4x8Ihr+YMqj
hY1rr+4Mpdr8V4pJJ+eUV/xSN9Lpt2Vcy3vApJMwoswpt+4muebIuukD7QE+ycpC
L+IdeNeByFNJrnANdVksSh1y3+ilPr6sjdFnP2pN3KG/wLtZlfA9CNjcWk+4A2WZ
bX6335YosxEq1FI1UbHjaSWfc2J6mgHCS99XiRJVIkOik9e73JynQqCP0fukqm9m
VkGwO+SfICR6rnG9CedeAk4MpZDdplix/8QYKz09NA/0Z6CHb7BjT67bAu2e/P2P
eEgwiIzYjfUqRLk3Fk/SxVASVQ6dQhmfDxTtVJnIO/+pE1CagpkytV1QbkP7sfsv
szerM74XmaLyoq0k6DfP5cwAmnScAYSEKGHlxGxRcaupEX+ijfkPgkqFVUeSC0H1
SEKnzJr1tgyEbgTqRwhtEtypFv8CMmt869fqSTtZXum22dr7X1wawAU26d2mMl8z
gkUilWMubqVFhp7OKa3zyU68gzwA7ObiJJBZXgUNBl33EK0bLccvSkEy20CJ69nd
wdxi0GOetX8hcIjeZ3MEZu4uIYLt6tLYc/isUwkPXijieiRnw9mAUydm883DIfeK
zyL6iKOXxofXLvpYz21b4Ru/lTC//CUVUNKO3oKaytKPE8kHjnKUJhDRHG8jFD2F
1dTEoLs4f+QrhqYV+Z63CwnzdTeHk+s+N9DvQKMlUY4WxoVBvegYxb1tCsLPb3w+
IB6N0JOj3ytMTv90CRCLtSPT7yFudwS+9yUm/qDyJRxZlyaaWgNy4PqWeCwmYt8O
UrlRRraSEjE7bPtNJD0G1mFwqMrJvxNcGPhSRxJNnQ8+dXU77gNFDf3PdkwMPsj1
nHU4IgHcVX4CKpGl0TRAUAT3ioa3m16ZYJP+b+f0zxyFAIwih6tlMIVDKpsehJjp
agN8QSRMGR2ApmrYPgkLvJTFqLpdtiBtSJ0cKWD70QbpPb3BhJAVg1ZHvvkpicPS
DiuUX98gf+BhDuNPf9MCkcpYFmTujGWEAB0VVKCAKQELoGpgHLlKg3LC5uSMTP81
f4edR63favQKSH9aNlCk3MlzUhIrPOWF4uR/WkPh7mGN3I5gZI0XYXyCTqOotI3r
zD1l9W9b8NLky3OrsuTRcxp53Am4WIKPkZFJLZ3lOVX5o2Ijomzicw4SSg1bGcfD
jWuQKCvysAGB8uKkdFYi8/HbvfHtQhiNR8LWJVRT0d3G7aLmjqxN8oCN0PzxtVgD
0fYm8CGxjf72lfnfiJpSrz9F2a2q+HNrLWaG0WEfP6ZSsQijE/07n1oi+zg2VyF5
FPEz8OOSOBIzdwPG1Z/bZyvJz2LYTiUezSWAUKSclrJ0Auv60qGYvW0J7kbItcXB
G00E8+ZuBQNyH4btVRG4omfDf6ZEH9P5nA/WRnzbpYATseAfbpYfQt6S/xcj53iM
iF7lsT1JIlIBIshpwepCUjfX4Ys08WY0jJc6SMo0Ho23tzxIcfYbhxg/HYLbO10X
7lne1pakO57+BpnPIssPZH2YojTezxSYE93lG7LN8QgPK55d/S6trzHHds/6u8Gq
DTX5WnKAcBlp9Ylkgx7SWYdCf2IyL0Yxl1rzBofAXdJr0gABFydX25bJ4PdgOw/B
sCJpMwzF7TeuOdROsCK8qyJ0UCWUEgmpUN5txSW93itcjGg3XvA6qQ2Vv59qdUCI
N4I/SLUhFL1cs2zNmUOnwm5B4VKNuget9s9COuVko5JT5YNvCQyO3/P8ssq7orSY
vDjP4kYTsetQRdCOuC30PfEy7ZMhCNJJZEAiXYbT2xMVtvF4tAqjaiiss9tLTBDx
9om8qEIMW9RVUKyshneYaP94dcSbjjY69L/+FNlzevN+8VOtjkNkI/MX7IVwVYQd
+JiSqnFcxia3G/t2Nrbrr1g8f/BKxW+QrWWX3s4X3WbdP16QC+cmDh3HHvtYpUui
oK0pVqna4zr6EE4lMBm8CXoHUVFDPD+rnbpVxrDtVvaWqu68uoJgfJuA+e+1bUz4
wTSP6kQ9prvJzeOG2LgfxFU0KBoMdpWIrn7SpXHHKKeJo7fcUY3yptTQe4Mu4tD6
Y04XkaK0MKGCfIXys/9hVWE3qOqzVQwgyWIsNh8camGQ2yUHUWM+cJrlmtmydoy6
EliLb4o/e0u6xB+RhM38nGuKFiqFY1gckFyfOmQNMAMhn2q2KMBxMYqwwymwUF/m
WC29kGdl8rvS+R9R9/gwJFh8B5RXZ5EqReDOlPh7V7hdq+zO2d24hHU1Z2fXiI53
k5npxXqwo9GIwFvwM/us1j3oSvrBMkEqg/Z1mXodjbVMHrUzrOf53mT9fT7zQeic
DLgAHdfP9N8ZfImZ4VdPax0KaQZaeaflIMzFnUcD6jE/wInanH8QQFC2Zfp/A5NP
nzS1GzGqD2DTJxpTfQpswqyA94dI2s7Du6p9hb77F+C9Ypm194aiwGB3TFW551Rc
C45YS6fAbnAPuogmMAUYJwpN1QJwy0akUQUB/xuEm/KlGGHsvLMDS7T+a0E6NsfD
U1cDSMdI2cySF5FRM3S0tEuodL9700IySzDc08ULLEGJ9pMJNUZ5tYeQAA4ph1rD
SWXdwFx7jXJ4QEWD6H32ujABnaG7YXwTWp6KwQQCXCS9H5WLI+KQ6lOME2NrPj/I
f3wcXG3kvAvkduIEdnR7tsa7QbthGAOpubSVkHRf1HLJYdm9aCEgt4mq71YMPl1h
UI4oOlv4BVkS7S2X8zraAukFkxKgn6sSLUQU+8+FPtNttDBkrIUdFflZQWNr5zla
cBBo0TDBLnXqsj1KCMd+gYngD0H5nybxEW7xKBq13zpGvJ+/vwNs+QIvUxyZRkjf
ZjmBorXDJFDiRFlFGTDHmZhMWgYkxZvT4I1oQlwAkvdP1n85fpel7ebciLXpLEYr
ikkYKMTYHT6Gk9BLOKJ3fICix7IETxHrvqa9CRi2Ti04wTW1LQ9TdBTxvrH16nAG
oW+nNprnnhDBrctBzcUawMH+8naOV6e3ChLROZPCKtZDy3tsgAeKOQOSZo5JUNWn
HGiqmWZqIMN9rt46hMxk71CCRhd5GvTGCRz69o9RHL72O8uj7qBon7d1cx4duxyV
WksU+GLgQyvZHhbc4sb3qKy5H/V3juRM8G3dP/hRSzhVdKjzYk2wBJtd/+M7KHAk
Bz6Utu0i/y1XKciwteiFvXnM1euZn6hD/fDiUIkRB5jBBFaa9TVklFIj6Abvb8sP
Y6oYbjGrMWps1qUigbfo5s5nK7uLZvLVhSv0TkdVw20P5ZWxDThlwyfiy24dsBrR
DO90DXAT5Y+6JDtkhWwM3wOvmlKgMGbiKLxE+2OXd+NzOJMsr8o5PX/O//9Gzg2a
6QO/hJMmdvHW/jrBrcFTZ0ukBiGowpkOxjduUMx2ICGAb+NCN6jsDAEBIimOYcV1
4swLQTDMn51+YUH3dKuDHyJJQuKH4IgJDxDY1uRVdMirNBK7bM+1tieK+AqATE27
FXJm+JpZ/j3ON4oggKM7SVyFeJZhXK2SS3g3D4kV7+sByOSpjSeFl+pzaiWqY+X7
E8EBToBisIvoy0NlwcCgHnUyG0djP6jzrsmCCQqopQaOk7sRjtA/iu67LOSofp00
gGIlFnSHmUU12GuhDRHWmBsl4zZ9sIqsJG6lpbeKOq+h1wBaM2ZAofAqDYSUNCsx
5AEplFQFw/Ep8nf+hpxgzT1NPDKhZ1rrinW4cRLxF/jb11OXhf1UbL6UeJ9Cbcui
s5YafSSNvkVsD7UBO+WZqD/CgPzejlvZi+eARVVmmwW7GTmbT3AcQDADUfkcAqKY
l2HChh3r6/GNtDseL7wWLNvzfQfl9peNkF2ViWS8cGuCicmh+FhXHHZdcnpIgcD4
MMe58MNvU3Nf/8l8I0OuAT7n9XhxlVXVhOsVkxtNW7iXIo9HX6I9KTEr/HEjGy5S
V/H/25PZypJo7AAaRG1i+RVgYuGHgvjeapiH7KNfASNjfA/HtetYxmNSQ6UagzME
V05D0daYqbpSdkyOjNy55Hqc9JjUXAmfO1o6EwEm0+5OHfQBJoxlIi1PoGP0uFAm
BYGXPtkgDjuCAxrwf/ypwVdyS3Ut4a9Onln/kb+5MT/5fLW8ThSYZk842Wo8jLz8
v0FYGTP+dff04e3Etyh/MhV+ykmUmWy9jrU9xo2prOdnkxSzjgyFW3qS4lurkXOo
F6jInsSSQD7b+PRnt3EK4q1XCoa5V+5x7NBX3Cf+v9Sdxlljd80U0FKRtGbt3Pkp
zYLb015BJfkkpFAFNJ7YHdIoJJs1B8EeLBORTuRXMer1k2lsmXh7cTj4IVkFjveK
3ZJX7KcjgzhpbSOccAwGXVnZwwQ3ZtLldJl6ofbzgRtSQc/U83D+84qmRsWAbJI0
bO2pLFYkaHt5MrYPtNFD2AHNCfIob3v3HagPIylylSVBh/IhK7aNAQkMqMTkfGQE
bxlYCbbJam1JTGE+TNoEEdEvDsK5HF9nG+W+VjRCn8c59sF/sP/nBuzu4p/zXz2C
GUagwTv1q4P0sSaiKx83b0sVAemSSk2mxp+MKUf19Tux2NbFriZGfVGC3YPobReb
rRcB9ocMuZruN/rQ1knevwfi/+EF+nK6ViUHZ1fD/i0GL+Z3gASit8QQ4ZQIAIQG
Lo+EDbZj4sEg+qh3uekejvvomaK2817Ro5e2cmTIZa8upwdTWe34g89YN3Hs+4bT
50Ou5TDRREYEBhgP3b0hR9YnGjlEUtLlefZ09S+u5+FwDXwkC9sU0tiHsX/4ROah
idxEjR/7Co+i2aLQXckZyq9bexrdngA6+rGU4tsWIb4h9tzR0105R2Cpd0JgDyyY
bLSPEw24Wh2dZ/uo/YKS2Rg2gIrC/rw8DCv4v5sua9TYWdxChYbNYhldB1JOzVv+
e/iDMfMi65DlZ6/SMiDL5NDAXMkzV2RVwCMMTaKX/9MSFiurCWxMdogK8/OO+WbF
WoivOKTUHhGdI11kzPxghWEF0ftk4L0rS8/M0VcHUWMKi0iIpBjrciRD5gCeJ0xo
7BEv/fHNymhYvtfDF97qrqUKfNHP9jo5qwmmpbvuliK/rTJDzuUzhBGnwZlTkpcW
FyNKbneyKr4rCKsaoPg/daPe0dUTewtEhDlcUuQVo60CHMKyAn8WrERcECMStMRX
DgNBO0pMxTT0Cw+8/xX/66vMIKuEO8Q5q5aCNFs2JasIlJ7JeEyhq2d/vU3xyjRP
AqIQ2qP0cwjZ2xdFtPQNMqGXnKkbgkC7Gi5R8+LAf9GwUPtWFFR/tJwOimUv4837
89SC2gSk3mYF8WPfSej2tcaL/zsotmz1gffPWjrgFiCiNBbjw7k82yUrqFL2M8gh
UO+rFctOY6IWCnVfaFvQGBNyan8jcystOQJ4OEQwUscJUk/w7lGaI2uYI6wzaAPt
gb7AYpATlgZhHbtjBEty99f8pBPzeL3i1QQb6DW/MvLyZMYuOW6qSXbCfOi6OTEs
HkxT6YAzFYc3lmTM0WhIcvdYqL3NuMJKobLsRZS0gvOsxVgWj4V3UuqJ8YHP4QSI
ELx0hKZdJ4+o+gMAgfE8oeA+vvOeeHxiD8Xz7Tx/vOk8K/4i31TpKFc28ZD/033G
AW1LJKfMxUVFCZqjh4UbuNxtgW880wnyN6O4YhD+JrPIVqc+nUNXwD/vdpZiazxA
qj5+24CC6tzFQ2j7QofPzuuSPdB9TgWtPNbUKGR40c9hLIdEbuL9krXl4GtvR+H7
BY8+tlDRU6Nymzc1o1AnzHQTUNpPuq41TeBj/NoS04w6E9+yl+790rH6Xbm3aCmS
i7PPulLtEts8YItwx0Ce0UChbAaum7vBZwGJN9w677h2+Kct6pebJVU2e3Qf5Okq
JjLI/23lUYqAfuSuS1Hf8PBlehCqpbUVwPfOFwW4RX9L4QPf9NIehw7ZIkacq9OX
j+HC2ZtvrvvE+6CSyNKkAt6ucbjbGscbIxiPX7UWY4Pdb81Rg+IpQfytsYw6ChGX
NQkBU8W6SoE80TVvesNRUCNMj08/ERbTJcM/45CQF+fo3JjGqJJPSK5iy67n7K+B
QdPayb5XvQierJbtgEeRFzNO1aeRoA7xvfnQYpAB9kAd+Uf7oSaVip5XdxAxejKY
w8+ApPIWO9x/rEuSYUd8/PXSOfN+Hmlo8yfS3/bWR/VxudUTreH9MWByrWCLApw9
+CYM6NzuPEZw9V/XouHtrBOFZzxd20ks/CZ/nctJGJHSB2XoqoSpPcwkUh78+tiR
C2uUS2kOdvuNhJIdX7T3tHZqe/sv+8ahyEzlXxe9clacbhKcgCZVbWlSD3I5nhws
xo/93E+tCKAx5qntg4IquD1TSxw5TFYg6fHELcg0x7Rzehy7ux+UEWprG6++jj+W
aNxO+Z9z7T3lBAFFNbPs6IAdhtyRhxtcohQZbFvad3XW1ZgYYNX+87s39l2EC5KJ
i7v3Z3zj96/lmkvVeTsllh+uRTmSYlWA9m72MlXiuMh0tsecujUw0FebFPBj+aEP
ThKS/kGMy8lRfP21uTDanSeNerNDTkzcCaDyiVFV6IldJEmOvAiqiXjz+AY452GG
kKO2VEJzlN2OKsSia5ga9neSIb/h38WqGiRY0LPfQxrkIlozPPI017Amu6T4FYGS
gsW5H2h8rfA/8auX8N2guUtUKo+e9wvAz2ivBwl4jGat9zM83V34ecbqCtYq6J41
5xzMgFcj6VYdJRCPIq/LRKsK5r1RlXOxrKEXnLH7uMc89o/AhpQmn9nT3DYbZDM9
n5xdfabSsjBoZEWl+9XvvQks6FFNs9Tvk+d5ObVJMnBOP4eFgPByleAqeUg3QgTR
WK/iW9zDx+HxKiQ36EepYxaZVJeksoW1z0gHb+ZplKbUnaBBkhgUhuZEB9wB3EgD
jkqfoF6qaHcZb6J0d0qtkKeg7XZqhg2MFUdlp5bvJlJYSe5Yj/TtKXEkyn8ScG2K
xouyVRHtOBMjAjDx85TTiMim0EoFCM3mMKJjyvFODbcIc3XcEAtaAHqKVV0C1wOI
cdtXAWd4Sjadav5yRXH8dGNfEI46xDdQvf0lzPDUXxxTNx409N4yUAc1ryHih/12
g9PzEkhBu8I2R+1zbl6ZFjRX6COlQQkuaiZGbqRSUdqXvtLq8GmkjxwlHOob/PAU
i2D1x6UaTcQrBPYBnX+GuW5En0Z9PrBWbkjulU1tYqGzY8tHWQEQAIfEKvP+Oc8g
XaTU0p0+1g8QdXOAUsWodgaj4Ez+dxdhsVcQSnJlpP6g7zt2ZC6ItR0xHYVQ3k4D
VPwqM9ErSrhRrdQdVEVHSK8TqXnS3Pzs1Mr8am41xocs6STCxjdhJ4cR0Dq89Iis
QbXGdqODHnSD9/w8j9dFtwVzlLHX2emqLEUDoELeyggYsEZZkSknS9irJ6GewILh
a7hQLn/c92LyCaZqjBhYembauoQXnCk+65qgZcv7HzVTznheJ6lylgryO5Q9KIX+
0FnETPNn0pLoA+j+3Ybp9gpIqhLraU3Zxh0SBEKdnyKFXCsHygyuhSO1UyptdBtT
xwAPf2Bl2B80RP+ebJzKkOwoZSaPWVuGrdeht45xmYZWsOLfAwvnFgoaTsZKTmIc
QOAsNYV8FwRXQ04T399HXCv3Uz8FioViYpgvmGpQj6KykPXu8xot7seeaG/E80yV
Je4eri5TTFxQ0DmTeEMFMM/T8JNDG9wcJM0wkw5DcDbQzs6G9Qk8hwCQuyeNhiKP
Ejo25IkGWa9ozXKvaHga5+6nt+vVuzUgnMG4MUha2GVvfk4fs1tiO8AQjgHRESc2
Hz+O66+NrLB8ZOOoIFRiK8IgR0t8kXOh1uKxRPlz0FcncD1n9VYg69kobSv4G/jd
kdG+1soN3in3X9UuH974p5hQeCU//AnLNZKknAUApLVMp2fcesDqJedfBZitkJ/W
eAnCi6ogsNB8cedqKEwYRNXqDCu3tgQE5FEXgv9PtsvgqCkoJnS1tiMSPwA8exWy
iumcxIiheoid4GZ+Vy5WENGZXc6guHFbXdVyRBvnqH+AiMLCp7mK5mhtktJA+DPe
t7tzxUw8KwQfyTN5+UgeF4W7esiZ8DDxsCSCTkqYuqtw8TAv+rwdv0Vj4c9Ab7RD
9FLZ9Ch9g0ICBnEuklknbT7ByVQeCnI422voSarpLy/cGglIptw62u6VVBAsZvMW
9kTzJ6B60gn2JpZVSIEf0SQPvDlNBf3fD7uyd1we596nC/M1SVh5A7WzuiG9f7bn
2Z0RoX2Aa57aLAFqdmYmptnarFph7VtNKDzo0yWG4v7hqytfrdA9+5wPDz/q/Xyp
4TF3Sov+TmPWDQ7tRkya9f8//kCaKLALDwqOoYi3JY5UOzNyw5XAm4K0NAV4/gZT
YUjgXd3+HfRYtXOz2sDovbFPJ+/fNC/LCk/amO6kYg0PSQwNDr5P0mo9fhi/v17W
cYVsfpBmm7qnA6G+ebmbrNYAgDYvR/+8I/HWvRS6AKaAuB2hJlnMFUHX5vVXycG9
/iR6FO1fTPt+SbSZMqTvpNv2Jg4Rcd4cmPDvDFxEhO/ITAa7tmPO7sNmiRmCC/te
xnzz/1dy+MViYKCI5kYZA7/JqB2BZroy8MQGTnRmTuStnI0i+EqxS5aia9czp+gs
mH0hV1fnzy1G50HiLONhqAsWzkIN3alOclI5bQuaQ5uXfQanjK2l4pdZBxK1Qudq
tmR83bzAVJONB8920H1zjOmcRFHIOwz9zgaxa3oj6KHm3+h2Yoy0+d0pOnHulFCc
tAIPUvyTihZgT4zIBcLR0+v5OBePkokyAYmobaRQO5jydbgYTGTn8QbgsrR9QzSW
A7FQM+5T4SvYmpULomNcMI/a0oYT7WfcpdgnGtcIeArFNFQ/fzXUTy/qOyyjxciA
XCGJuO4Qg7axywsfCayDGGu5LFeL5snPGfjKA74ct54wLYlTvvJ/sfZkeG2kg4/N
v7jB3CF0LC6hVW26N116NQoJLKT6dZ3S4+N/Uy/SpkSOI9zpS6JjInD1J2PEISLH
r+uoKPeZvamI3S5h8AilZ++pn+9Kqf+rFj8+Y8+pGPjA5jgToh3IOBTbMZ8XIReh
tvM9df+lhzwfbp5K5LjX4u2bEx32TWvase14izsT2hiPhvg7F1Q1DmIBzjviuTha
3auAdRfaRKZaguGR2Mn0cNhDJEo44wfEJb11Nj7u7b/qb2PbPQ+JLX13+M0S8KhB
QsXV9eyhU3k6KxHPtnondNv9KGHQBye//R1y1u1r8SjvpWjkLEvNQiQ/eNPZ3ggC
JCB/VGadoIXuY+RIoTMJ7IOpqULUWuomt+5s6don3VoVZWssYRL4Ida5jwrldYqA
6jt1l+Y7iJ8ryUHDPIji1Wo4hRVlEfWQjKwB7uZrlQ+xcTB9c6BQpNTb5HAHcyG9
fVCpcxS5xwA+z38XrMh8EWYp0dC4GzkYNmL4IBXv5kfV+yfmsiUxBjYsSZOLPA4K
uwKxsJW7LmnNYQr8ucBH9Hcga4VAkOCvphdsdA4F0NwaVM/IRtn1NqMmUPGM5bWC
K4+hT24gD+QFxYAbG+vn0t27gsqPS6xSXUIQl6W6nLbe7c+JHMJV5Is+a+IMcy9J
aBCTIMz+gCpksnFf/k5PicBJSQBIpXgzZGJ5nIiYl/+oigCaS8PGtcXCAaC3YC2z
sCEe3u/EH9hmWmwzbCZEpkLImh3u8eLbulvEBq7Nr9rlNNFaVcwuDHviR9f6JV7v
atIquMUXn1sj0cZf5Gxsn6HxGP3PlA2u45L2wr8ng+XNCxUjBZu2sFUsCJ4U26/s
6/MwxFA1pLfbiAwXa4lFtxw++b36/+zw2bw/AQPnNAvm0QAeHL65uWwvP5vw0X40
TU1gYwQGoRIJw7uOab3VK4wDQG/mc0BXR7miN+5hpBOmTepxVTQjpMIv8kGlCxZL
Xt/wStH7RL08+5XxxRC3uSwk2o7zaj5C1gV/6Rh80cOdvqGTLDyj1hOk3tKBmt83
OwePVYbIobfK+qbQpowB937s86A+s1+MDdI+2cSOQs4h58ZwFcRT8Xzt5HJtSMLF
O/nSqEFEobEofskvHpWZ4CHvuWsWCpIKwIL2+snvTU+GPn6xP8nSjai5kEY9nqom
kivUtzOoSJXX3VRvjFR6OWih9UJyQi7IuRTtGBOxvsytjgAgyfz0fXimlqalR9OR
A+TPuOfNcg2l2v1ZxxckRn9TCqZuL4ZRYRGKFLQENw0n3vwJcXLHlDTNTANbCGQt
Mm67ieKu0sVQLr5oozpOmQzF7jzh46xtAL8zp8eMgXrtG5UOLyOMxJmI6gNG98mD
jQ1A6dQC7JWqZY5CsZZ83cjxRip8PJC0iMp1rrLpShHQpa90Vqm+vnmdPEH91uq1
j3bqVqnzX5iMSySBZasD7O4GwzkdA3PPf3TV7qZE6X0D3IM/d5pC0RMuyFZcL1rr
eKCGBmDjeoP5Lz+/QW7S+b5FZ8ojQA8OB4l5L5FnWXzDcltav/4RPlx+WcfGEMzp
v0sToSIDOKWTKOhvEEenggMh8xhzNABijzkmBWRt5Z9k1zb76W5LNw229uvCwUia
rwiroCEIAh6hwCgN8Ba6yhRAwKVjfz+utcpuqOQHMbrVPMCIzzy2LG4B1MQ7cTd/
Y4b74rmhEQicPXbKUM3mX61VNjb0REafHATH/v/mt31LRuHlMd1D2jegpo9TGdQ5
/aSdPLEkE0OgOFX+Of+VGPXIB/y6hqN4qJveSasJkzk+Sggxa5ktl5esspwr2DGF
CysIG/RCk9r8ImgbBMeQA3gTnLGI/QOmH8STe4P3kHgxBJ3jQXHIj0LwWyTTzAh/
vTYX6e0blJHzY8bVMrrAHVgPc/KmRlkaNSOCIxYlpEsQ9TbOjCN+lCV1DcZibk6h
Ygd8peJqw1hz+2bvIfgjiasGbNY8jhWfURzkibh/UC1wDmxlGU9k6Jn18/G2Aelb
dYiTeUTSKQjcF41JJI8OoxBa2MdQg8dWjBnFqsmhSb4Ep12tfiwsyU0SLv3cB16a
J7Ea61cL+nDtsICFKsaZ0/x0dGTp18olYb8cAKpDIb0uzFofs+28zfo9THGYVVop
wu181JTRJonk5U9U00hXaDw4KQa2pOB7pzm4OI+lVuFcFU7WF+Y1xVv1nhP9ulUS
0OwJQX+zyig0zLgoaBrpHrg0WxlAcQutPGPBDwyA/txQ6Fywr6Ito1JrJk3HnRyE
RnSvBO1sBXY67RY6rxw7zwVhiiNU0Vxoj5NRc8r7AmPWEXvmvmUBePUfBfoC6G8h
mke5uUuJnn1XDUwOJO5QG6c8JpIGKvO3/PWzx7hb+8JZ2dzTHlnZcZ6i4c1OlbM/
gRr+Hfnwlwy0/dXb0ND0Xfi0PEQOdLtyOWLBBgozqxD2+oW8cnSJhatv2qohGwjA
w7/bfLEsoPDNusX7IR8mvCNaIcEAB/v1QYbey0mw7fgv9KEn9LiRWBW+WLhy20kF
iv1louqeRxTFPYNOigYUayB7ad/VfvQtMBejTR3U4vC/tOcPRtAcQljAKduUoaBE
0za5yOgPAPK626vlqunsf0UPLlH39FL4PlIqKeoUYD8U+ZlcKR1kpH9N8OQb+IXp
ltaZUPG1WkE5FMqTk+nH2J2DXPc4ZpGpSvnd43rtsIBd9+DQ+Jluv5xsp/GLLY9V
rIJTvodWUhikXZYtnn+1YZeOkOImbqJvPvgEzeXBSGDHlw0PfUVkCPd0zzhSCbjT
YuQU84K85M8M1hI6T8WpGgRQT1Msr9SIzndIqlQRDGAUnxNQz0QR5pHPjyNsMTrk
7HzLYbi6OWPjJIRA6H3TwcqVRuEVcgJn1uEbUgK71oLCue0Z/6RiTpVYyxT+xV/z
KVIsjIJigX/zMNITeM5/IVxJzWYN4/gT+MZ2FNzNA6xUOql6yuiIhtpcb9c4V/JM
1cOri+4mJeItY6pMfQvOajz4f9ExBXSAsVdHTT9eRMI8swYFa7o7kT+p1AT1daY0
0LW4AiENn35zhJDgH/XxNGIJePi/HKrujOA7jkeeZ8mbbouwi/WNksaGfx4Tyb80
bw1brcx9b/gEQxHs1E65uz15Le2HIQhqdOIM+t0WjcHDtPfMUr+SV1bB2PoLVQ/A
aTtvCWpCb7Lx6x2Z72ErGia2g0RoOvvvhsReK6JVdaRI00GVrUEDVAVzQ3UT9t0E
P8A9XENk6iQhfFH1pbRXk/o17cL2kc0iJCfXo7TcSTPCLCVkuugHPJm8umEfaONv
JIUzSIACyYzik/4dQabiKTqMbHcbztxweNqqVZIzvcFjJ1wFlDboCTIsVHfcrYRi
SsDDELj4/1YF1aSmOwFFwI+ajXNyPvgjVjxGoDF4eSrDR+BFg9es8NiQ1+gvD7Mo
edArrLh7uepmwqqq8sdsWl8vM3LntNIyXy3DdPidw1rbdDqvCEB7zxEhR0omWR0d
P/EAg7L5Rh2tPnTXpu+jURours77OZvWKkkBXrhthyvomHMTd9UXG8CTtoB3uu3v
FYaHKc/NtOvBtJ1eK8ZbJFtofjoowNKOpng8Vx2IFtiJaLBqjOiaZutkXzK8CgeN
+EqYlJk3QYcWjfFJlEhmjlGNra3mEOOCgxljwdSk9VtEuGQRoCYeurhpNS9y5g+/
Dcph8ke/PefVpyn0Tc++xb1AE/0S1iF6HA9gk4r0DERmamE8jfkF6rVeQeBngM/c
WjJZOo7/LwuWMFr7VeSvWPrXENB3kmX66GcsAKyDICif008NfRYEFmsyoVK7hXZR
t8NiZTL7xhEPCJ0NLhT73m+6hMx0jzTv3q80ddlQ/ngZuj120Vu+3vhQNkpAWJci
NpTuJU9vhshqK/CpnMkUlpWJNA+AGXCcM3+ETmAuX5mJoNrHQHix/eGEUKzje6J3
71JXxf/lRkjoXskDSYdHcLBj4AURLQ6sHSnTQu+yKJ3IV5PS/GhXPoNorSGgve6N
MW1j6miKbq6heO4N8Bj++/lOtxMIuyAe7vZw8VRmWrFBXcNZyLUdG6VBOXCsit/e
VTClAMX039PTTWzZKpEboTkNCj4JQ7l3PE4nXTHjZ8dHA83M0ssroFYa74EtpWzw
oSrgQBEzOZ5K93vYLnm7YGwh0hKEcAERyyU7iQw0J/DY96X+kEd7xh1r9fFsd5VQ
YvmDkQX8AGIT/dkHy0JcBB+t8E0Zl1L1WMF78g5nWtoCkiE5Sy5tqKr9GPZ5JwVf
tlIoqYWTtQ/ErJPzOZLEBTrURapuUkoqOtQ00eJk3hRMw8qf7JsMhNjzEa4sPLzk
+QgNc+FYPR9J7D1KMUo10N3d+z1ZFhoZA3EUfPY8CDqb8gGSfZO3Cd9niUS5lBph
26dus0fgggw0yPycsK+1VkuiQR2/5VY2oWHQfjVrtI2tW2hE96xjHlOrRVKadxba
gm0zRrVtCgdGaM/uLz8gEiiPXASzLNyRZBes9DU27VAs4+fVBAFbSyAlAasvCFH+
s3jsVaPwh/nxLRPqI7Ps6illtY1vu1yMKDvVsGiKcpL3KSqhxVC1R6qsRtG3M3vC
uDW8XFJWCrnsY/urptde3M3s7MU536JX04pVWmIRzXe8wBK1Z799FDwviNwQ9SL7
xPpL76MivJs3/994AAH4fQ+q48bacHAidJagbMYLzu6UrQTgv+RowAAOsCBiHhIm
m/kct0D7Y+t/DjQZj6tZ9+9KZuXoMWTHBjw7SjEe+NMaRU9s0CDiQ71d6/y4OmjR
8mEAZKEBw8RhPC9I52RWgSHPRVb79RylPpR67WuXsEV1uj4KuuZozAAW+DUQOo8f
mccyDtcwqKj21xJDU7Ig5NtrMcH2OiYyyvI7jWJaRBuAsuFrKijc55n1NQiPbaSP
ov8zuV9XlSiyxFZwBCRT6cfkPMTmpG5HdIygEXpNiG8gX+/kgOO42FWslfMfmhec
K1oDSs+a0erjGIuejcW0VhgeI8fTvYkVHsIDOgUTdQ/HD7RH0pYGn2gLU4bZ+dVL
igrGbxVWT+pZvyozlMPhzbRN8b0j4bnx0MxzTmhhUMJT4bhVmN/NhKZ407+M+m6o
A0B1s+rwOKRGFZK+iDIgq8XPuByDyEuwHYWFJ+5pcbFw34mPRum+0nujLsG0sNoU
WQ5Yg8Ha3mLnKN8NfJwkF3DQOy3K/PvAzWXkavQqjzhw7a1/GzSzbDq0OP1/Op8s
rqwu0iFdYUsiVABzW7MeWTC/a9C4d90uoZCtiLIjxenqIl4IBffDo1bN4lSvNlXO
Y3TNnP7szEQ3XCDD4buA3pVjrgUAmDrCCckm2uzHBxKSEubsquc0b8EPzE3NSlDX
6G8Z8EtciM3BxiRGTXw/wv7qof3dmVQ6EfIpDUUNeiYZMt7/N4q4M0LYSOjfPif+
9oGkkj3ZC21S/6EOc95VUlNpFGpjFXGZDfrk8w9Q6C/x9xOr/cFqmKEQKkDhXJUv
vlw4lfROH4ZRo4PlrlHom3uLn5nH72NrReLBTQXnWIhxWovlHJl6YhNTcxyLQgW2
7Lv5GctFJPDGHNkMz/vaobcZjTykrhDGrfwieQvenvm815tA0dE5Oc6sGOjK20yj
eUacExq0GPkXiq83IuvellGFNJqcRG80vxICGwjhUBCTzOOi4JeO4ozk9GMmCDv5
Z8GWaodfr4Z73HbZCdXjRckymx7ZePVhBc3qcE3ih5MBj+f10Wf9kBwlMGAV5InW
kPl296jMgzO/vWhoGzWv2oJAfBSe/tMJ14XCu/tIDpiZZULP7LlWVzY2pzdBHi73
KYjG512d00QlIYKrnMd4jEtL/TY6OxjQYI2WArmBpUPZ49Q+ILutL2e7eHCgZQlw
RefZthiPe2TSoNrYESEJG4/ccw+qI4x7T7nGnHRvppo3XUQ0EO8YZE4Ck8h5cCZ7
ka8bBuhivdBg3MP7KUlFU1HdX/nrk9qKgk6wmFHp+jr1tJ3OI+Uewp7LQDKM9QLA
1lI3LtVUev4+/XennNt6Nhyi2yBIXzVIEN31IvM1SC0SElguiOzosfpE/j/3eHId
NXV/GxvYVEgPWln5iT+T48tZVdz/dMztlbWfgwEe4YcvTkqax2m7gH4l4HljeMP5
/5SjobKAgvr4La13+LwxJBh6HSu0rZz0InRYqRNhaB8t7VcFrbQ5i4TlAFYO8H3q
NyAA10Qp7p+x/d2fqDX16okVjjS7fnjCAm7UONdHsz3Hiohm3yeimVDpKfoD5rX6
rX+Au0OZHGJiwXeuj3aCMVaYabSYW0Kv/xcpt4I0sFrnLrjS23Bvcl34U7vcZ8Bg
cMukQ14m2yV3swDZzX5PVF6xrCjJ70YuEy1ze+gXwHakGPEayLELY7zB04S5hkiM
D5A3ARdFOGaBu73dLxDgcOFHWh7N2wDFrprtx2m9k30UE6qY3PoTWd+ruV8XVFP/
5olRzYlS9cqXvVLUjFoyyVkDBZwt0S3AIZOnQ+MDF8MczlhS9cIG1ipFjPeM+e4R
WQGlk9KcczGXR4d+MMMdoK1VBEi3JReO6s+xDe8dXKvzYGVmd6mlOwCHcW2SnHb5
yTTTNSg4w+6kIwTrB6Muvu+oFyynUGVM7AKY525U/fq45lRkw7ZJWmlavSE3S/op
dt6mKUSHzjN8FQjqeX+vWD/PDLLpd9C8mGwe5aV1kqZ/UyvRkDII7D9EfFSZuFDl
L34eSt6zGGea5/a6qvBN5JcXe1PfBo4d1jwZDmIJ5QysW5RiQeg9u1KYSELmcUJp
rltmVpDn3UdpQPRVyp35HiAopaC3YMsfxb9hypf0mtWqF0qXkexl346pWvd7rVPy
Tua9ennSUDlIur1wUEdYWcW9DRJcWrSGAESoV825z7ZjCXvgrmg7BUtiY2FtrD/O
QxDnd//ApsMmxS9EaENr3ahBNYqX9MhyTx4ignqt9N6cQGkp28XrhIIWQba4dmJL
5xSl4pqeHyifWA8pFbfew87PJVISTBdtS7eUlavmUej3NEk6ezp+AP2isNH1BPic
tnhvI5PS0kr9FXbJ4QpHsnERsk4yqvEQ0Y3SE4aOM4FsyV84fcT8em+6SLfdHHsv
i9100rAVequJsmQM2RGAsfaGR50KDQot+PfkUd2z1jehB59I5VAsUHvx7h1z7nvE
yD7F+nfO2+EaQ0D1n5raj7QtFKd41aFC8B/tFO2dXYqc8ZtjtIPY983D3Pro0ovQ
aN0kpfjB8QPCd7CSYC95LdBIrHDpdpjxUQi2+/2yiBtBwFAGdP/1R69MNpxjmrOB
MvFGVkeoakPjuvrjZGw1F7t0Yw+vL8Q8Bm5MCs1y/8B9mgjJNR8NnT21Y65I1vHH
8QjnY5PThyh9ok2LbeBWUbqEYEeHdRcejTNZFvBHM6ikd4kJQEm07YHf34uBn6Ih
izrWSaIIW5EUgcNrn2RyH7Dozy4EiDGttEljfmuNzPNsUYsXIWoAJ7g7bPDWlBDw
/WhAgPXUjt/TKAmgQAgMnfKLcPRpm6XPzTvmAlFayAuG/XddhyyinOz1dWiVapgr
cH0EigfT+s8SvJoL6WcU7NAjByXGN89Boz181MJlF3rS47d/WCe74FgC9FX/AlQi
SNUkvOvmh06uzScvBbPTzl0h1FW/G04j1zoYGqU6kzfnQwd5cjrr1LY5pLC8RRjT
6+H/29tAjuWkZJI6fx5pDAzHYfg0HFWyDEIIZctNgnX1faGiNWW1FkI1sg+cx40b
z9vIUwdMtwI/ARHA6jyffU/Wdwz7zlkRJRUpMGdHPp6VmQ5oiFa2YFTgJso3HQHb
fm8dgsCPjohFFmSViHxXmFNaNxIs5pSVMCzFTS0Rb6hRhopfIoXFSWYLFjxuWWSl
wcEf74Ewf0aQj9T37Q9965SyNhbH2Ydxl3h1jQG32gMbQJ48/rdndqijgk/5BUcd
4R7KpPeQ2I2XHFBPLfpnEg3SUAdj8qoRFzylU0tDqE6qvNqC63QjLxxV+FcR3LRa
3ibLOHC1UUiGJQ8BoJmc3MHz8iHD8mH601vXCrPPyBKR9PuS5rI7SDpIVIC2tGoa
Bfg5d2hrSC0evjAdmqKS6Mvnq2DTN72ohKh1AvWwuMPi7ZXJvDOKtc3Wa5q5Hc6K
m32m7Qmo97gSbuurjo6ywjiJwXXchkgLP77sU/2GzB8wNSq2ZR3cf6CJatcLFHph
QgCtzjNNZAQKBGwezEgDPBO0A+IFJyEvqGuuMcLdqOPKFrzi8pQFV28UwjqPJ04X
rhRQ7EMN/WgJwG1gjjeT/aeu1OeaGYT5H+iuJkYCCU/MTa4OoHnXJvy8ERhFgmEV
L9IxzDa6ABUEyOLzGZ0fvAPG0sF8J0aFdDGxvz2fKL3WoNLovxSCPGkaFjUFN4uH
TUV/DC40w33jM/JzvCb2EDuJONkUmwxl1cmIDL54W//+caEjJqsc/UvS7RDZfwhm
s8nT8u6niW1of0ASVonDqbQlqorpgGKWtIbhAbI8jeygZaE4OqiExczpN0RRQDt1
s+gqifEO3BgTHYQaFEkB885IZHXKWqnEfdYRhN3KhiWUQKiJPFxJubgSQl/M8U5r
mim6orX5Wu1r1V5B6i69DXwtb95LfxB4xrSkq8z0hoBV4GteAlgy6rpZc0RPbFMQ
91iQ4c9DIHxIeBne49dEoPbZ8Hk/cxuelobJhNhjvaqLfwb1JKE9yPeTW4inOluU
0U0a98IvU3nX9DIrMChKuy8F/2AFb5Xye6+vuYY+/ujvSUdN5yM01UPiKDeBGi8Y
aXMEB+aZgf/hkfd404JLUK2Kb2sEuzoFuRc0RXYgNBL42CG4Z8FBkkmWQd6pWQbh
wPj8aqCB2ucBv9+A725mpi1O+/Nxd5xUTfsDInI+xoPUrqz950kZcgekCehjyoOW
SQezJt/EVHEu6NHjAO99BbZr+96b+KmD0AfoWsthzP/tj6olMnwH6W1qjfLe/jA8
MxgggXA7ZSlJOCBB53Y8TJTcjiCJgtrKNSpmQ8jfpSpKaliC/YECxHsMb5JKVsZy
rxSqmsYFbcemshgJl70oXoFVGXT7+tDy5SLab1M2EZxGJdnKif6jzYUOfoQ4YQHP
EZr/ReEFLifMf3u855wyXkAiHme/7wZq7mYNoRMLQnVWA3HMLz3I3hb+rLbRDWai
iCR7eFgQpvXgck+7LVUjdchVM4guU7n8OplL2yVEsu1ZK+ojC6+W6IXrKmKfhnMs
T2ogclc/90xLHOJaLGADFv+R9zgSK2EY1yCD2peUCa/V10KqorItNmWm4ne55FyE
ZlcdM3/sW20EB2zKiKID+99SaDBmyJE9yW2u7rjDqYWHvV08IpdcNUVUXp1nFQiu
ORhaoCgiZL+baH3bdYM0aqzHygsu3zkFaKW6pycdLyVMHgQI7pk/HphVw2uQdODs
JiRgRcSHSszeULIv/mv76/TbeQGA/WvacuSeECB/YPsvad/sAudz2rnLZK40/wfs
7l/bsUFBAWL/DL3CSMM+i6+ioa5VMAcXtDQHVG5JM+TwKYAIqzfo1E08AddtK4oR
t7ogZd4mdP8NIUdM3tduKVr8Z826tlrZv2V1AbUJjwkjxxm17xsPbdytFXvB+QKI
k6lBEpWS/4jz55RUs+xSvxLV46C0ZlgPwXYFUlLf/73sF4qaMFDmGrDi4RWIV4ot
UsyM7TKWYpS5mcEXVK0v1c279baWkGy7xl65MoGujZ6eLO3XtRCF5uifNQTu/loO
CaLrXpHZu66sKmtHNx7PEXSbF7UFsjmCIkw/C98i0nP1YAJCKaZiis8nHJ628gKc
FQuZfg6gslWkoMCSZawiyIgn7QCn998qPoJM8ZeVrXWkGe3/ARrxkY3jQ2vnXcuo
w9Ku1HUL1RDBf/sRik3tjcSEs0H2AJ16DA08txfm8MOyY5zMXkXKP+JX5T7EVlYV
yZiFDFsd0B4CJbhQVZtDWEgWEx8coOeC8IF6X6ADa8lBD0KBSr2aSCaCopDTrDB2
ttURnXnfE/GjET9etCvYwPAYdLgSdTC3rronh0Hkg/+qx0QYme29XB107tvcM6lQ
lRZYwNHneL/XVXlKmQSgxnWms3XOs1nWFa03uJ+P444p5Ewx/SV1gNdo8wyiS3ck
qCSjXbxwO5MsOJEt6vkTb3Qhg96Jyl7GsqSke48jGpeViBplE6VUAJ36m01NiF1d
3RR+qeFgfXB8RIqBOTKLdBuIKY6gbCFEpLnOI+cfD+U3UQOgpXHsAFYCBUJVZDR9
5GDhQyPKD9lynyHwmTOWCIv0jZGLmf/x0JW53RhU6advwOyHpKF70rwENxFAdeLl
GLpSkNOgH9fMoZ9FSAS1Sp9+6zKnL6kWMJ/dbDQt+IzAKwoW3HD8qn2b4kp0EMTH
5aJ3VG+ldpcyomSX5MhQmsdYWATlP7Agj2e1+Vd43+2mOwu+lxX2TPUcglVPto1i
dC5fK1TXgWbscn3kADDdWoCVg+/WgdJiiHi2bAo3NRcOXRZfQObFzsrN1yNa35+/
T4BPSZDATCV2tsfydb/0Pt5PYKY22QISCXz0qMRIvU6+YjqkwesBSekXg2KNdiXK
gArv/BuHcVOhqwgpKXtnG0OeMi91cT+Yu2f+dug/iAD+iElPnsuDVwfnoMzlp5sc
a4d+niMLzNaydtbviE/UG314TMqjcskjlLb1W/KGJPZz5NxRteYGtrzrqVEQwCMA
1bK+JQRqZCH0jfiWMFPI9w1ia+9WZYWgcP1883tj20uwRnbC6OJigwrGQi8oTwww
pGCl0+FVKv0Z/TuoAiHwBV/gP6obwOWWxPHf0xb354EWDmci0XpSmOZMbLWD6zZX
QVyeTVAOM13hfiKFoJsnKBBhejIQAXD8+2CbRJM+E7BV/fGMmg6MMN/zBfWmzx7B
DRuiexovZr3AAsB0n9ZCNk31FFGyMsnqGECrUwSbC8FLkwbDze1TEHgKkdlsZx/x
10H0kbbFQQ5GY/qbzlbOMPJudWBzNPSWkJa+GVKgonEFzk8LHtGhUVDeGvRsBQDM
qu8ttEpX+2h1akOaJ1b35imsw3Et8XLzJhXU67TqXgA/fS9zW9rglGbGlgI/+mU8
GAY9DJWsRbwsnl/ZMSsb5WqvC1OaryASHPSWkbqcrK9+0779Fsheps8ruFlKzDfJ
vhVmiBpk3EVd3IJV/evWi4MGXGRrUCljWf7Z64YD6mBjW3hQmiHzn9RLRgShZLTO
Y9nAz8hOwi97BlU8yzMnqBf144H9Ut57TKcChReF0Px0zaJzomqJZdMOqZ70ket1
HLcn526ewUiJEgYT1p4+x0jwB/fN70zJCml56kwRa5npu3+bXHE7WOyyZPdcvSm8
bsPwJlSgx3YFYQ+gJIyHhsZ1p37MSdl3SbfZs4VKoLXzFwjo3vq2MEgNaWfbXomf
HC/n/pAP/btISYBm/X/qEevHZa0LYv5g96swvSaN58trcodJ//0sLxIr1QNTXsmV
kyJQ+WRiMzYwcNAkvz7JCM/cGy5aaSBAMA9/tO+seeTtbR/lbbkRrI3dgIGbUbTC
rU6yd5/Z8XNFL6wm2uu0xM7i85OjmQW99nakUjO3HIE1W8cj+m1k+a0y3Pgng/wa
xS7guGc7J8KkX4xg6s1NfAv0KGYsZy1Q1XAj2+9ufyxor7L3TEISD3f/XY75Qdbk
xkgr6taXSGDbgaK+iajmKe/bT1IYQXOn0jzsDK61b7hGHwQxOHbBy7v9E4LEkN9W
3iralEvbfH8Pie9xD624v9JnL0e+3DFDLIoi2/bCHN83MpeTITA4Fi7w6BjZjlpj
sTYtMX+TYEZzMs/13wTffmvmQQ3ftK3+AhC2VdmJprjh9dUKYD3C6q1G38wMgGdL
qJKMz03W6gHeIB0nHD0KsK+CB095jP2I0fGKKMZPPJLrz7Xgjiyz1+cZyo7IF6O9
nDDs5NKQHPL2xOPRazKw+e1VjTqwgX4mVnre662BNxXz2f0P1y6hpjDDoR7jwLuK
G3Y2H2VbSPQHZXy83AwYXdqcZTpfvfZVvlM4s5dsRPJgTMMl3KDNlC+9/cuNuL45
bPFN3+jiXFyNDjSMySGoJJTbBfB71fC4Vhx6ykAcDJK1WkaYwlxwNwSZQAJ8oZmF
UWeE+GnaOKrUOsSDR5natNtSzxzga2eMtty/8I11pIBO2RVlXddWLmwgmezCsmHH
fyllThQ7lF5Nc9kouNUOLXlYycH19SZy2o8mF2Ha27EuXbk5xbFe4TiCI8jCs62T
OjeKTSrAGdcEJgbPeTS0EPlarwyjUpjDdresSsAZQ99eG/Qotrbqyj/bplrdYifw
Q/1TMMOAqorCKn4nhcg9nM70RfeGW23x51pmTbwC9qqUsajKC7HdgpvfuYuAOTS2
TnhqFzFoAmVDATTcj0OTbMdYbupzysS5R8i5TQVXiO+f4GVqUcL6FXqaxsv5mVCK
vDCeCc+DQexciC1sOnSUcidjvTV5FxjBVDO8g5Tk8/8w0OpSOORYY5Aa2L3TAyb3
iIGIJXV8g3hu6tCLyuHrE4uHCAoR/8x5tTOJesLFq2KXmUXO/JZwq1lUIbkKfDts
N25CrgQTu3+T+YUOVVli5FFg9gqZdvLbrZubnpbuPKkPgyX0eTMnt9bStk7HNmkb
Ry3GNNCjJvV871mdGLwNq7ZxtiFU//dLmrM5T0ug3wK3yXLr/9r6LGMRQZK95Yx0
wtlavq7gXauTgnCqMNatJMSQvY6hWMjLcPPZQbx/kI6D4eEIWMhtSlhTpDov9SEl
zt/WgW7rskgDfOsqN81tN4MNlIDhy9z5zEyT/uqpzZ1R44IUxo4pq9G8nU1Ynrvr
CEB6U0hY0+EiiIuWnXpwWk0KQwIOuuzwgafdUQDeyAz/FvYAKIUk5mGg65OF/dXn
yQeV16hNqbHSvJcEmYVlKgVavsXV8nu9fWVjno3EjjLEX68wZp6u+a2f/eSf6dDf
7gSMyFKtHo8Cc0qeuag6iUI4bTQ0+3Yvcc2CcxDPPI54Oz/oKRlq5dSkQyaz6vjL
rXWLP9RAWPSajZXDLGD47Kq1AZmaWRVIRxwEQnOgr4SjsdTjMBqFBU9xSAzhP791
qCS7wSqNz7+rfrRMq2LINvtkecz3rgvc7YY6qjJxeNGPyAI2/8nL1El+YD+TapiD
oOtCUpPPA1/IfZqk4AUivM2cVy256jE+0heQ6syfAZw/geQuDefwLsoo4eoopJUe
LgAhs54+wso783IHdW8UFJxxDG3furvmQRQHZkjsZtpC5qSFEg2o6RDiIFj+puk/
lNjKlFFrkLc/+sqdbeSDYu75vDfN3EHxYEFd5l61j/nFA2hk2zLF1fPqfJ0kWWHz
ZkJfaKEc1lMTRxgFJxwdmsCmGUdjHHaD2joGh2J0UusIKGrmxmD0SnjgygkmBz1E
OHVtfdvLX6tDf7cwvdQGjXjh1AhhkeRgyHpADhsdioga73XjIZEgVUKBCwQO1tlx
BHSfv13J2gOmbXZV6j4K6ijJBDgGXcmKRfd06uEsVzdc4GsOm7Y0jOQ2f+OjvZxo
EZAHNWeWhydTENuEbHUTw+sk7hT6dM/8/iiXdZ8juQKrlrmLIeV+Un6qU3Y/KA86
7bh8hpYfoowInayBd6wUVIFoeTtkhUZddJmQzsWy70aXFxvq0uTpjfGyyCZm6jPY
vGwaom/9Z+3ObVWhkXIQeKMaLNoIDCPM0qiKiI8VSdMBMgg3amIJ3EXlCyJ6bWTQ
XsRL4AiikFrfRd+wmp2rXQSqUtZzPE5iiEsrIFsjevihwpftbo9Mk4Xx1xGRx272
G/2kR4NxE/u1P+X2Lqvj5a/BciyUo5pOnt2hzQfqc5o0BhT2Nj/wQ4Fzo488ZlhE
pkJqhwEi69DXO/Ag+QmZjaFQSckS2TDpFcgyjpZvx88zBM9SPt7qYx/a2lg3Te44
T04R2YcHX/BZWKxdu/Xlq8RJM5uUMUWsM7hzm55h1O8j+lBAMGoc8cn0XNbXCpG2
6glL5YMrsItp7tZ6LSJsd83XF2b1aHzv/HabC/Dz9kECFGWDicC6c5lk8mCpyzys
m6mowA5q2daYeS9IU18onuc6XWrETeVEgH2BZHC1dg5vXRDyGGVJ3JcXbtX3O7/m
5yrc0KaBmT/ixBVGDvIQKfP0AYP/yGixGJvZn2bonYehdYBjaWxIZ/6EiBBfQH0f
NQrBC42NHA2ObP1ETuumXNgAcvocdLB1ttlGjM06VODw/4JDtwZOdq2iSBpmwgGS
txY4O288FFh5Zm36BcXRX/Iir6ENHk68KN2zFDeygn1CF6yzR5J8tJb7GNP57ZYp
AD0XC3Ra7nLDG76/OHky0A49DiVOJHzBtGJSDjMSkc5rXJLBNaGLmUom1Wf1qLxm
9DsQLXaCAx07lE+pmO+IaPYrbcZ4c1Bhy6GLPDwgbML7t0mMWr+EwXu9nNykNKOM
6qzdNb3ADyTSBIzhnCMC83HlwDnMMDoN8CVkXIaXdyFvdDtJ3y3QVEI+D4OUYe2E
aTb7CuAFr/A0cbJi8XVIELdT9zcPBMUyfzz1jJECJoq4beefcDWS+NQbi7+ScSwK
LWi0AoYa4K2BHS7BpJi2k6KyG7s0UwflrjcmO32Pq1raYihtVHjMSxUgT1tFEz6N
MwrrBChZS2urbnQUZ8yQpyp17ivEC2xnTL5b6DvlbgSPIW7WmLsSLz1FFSwxfgcH
ZCecAZ3F4R5RwCSLh+h1hMuucKywAJy6hyEAGMdhKyXOA1WrzAEU4nL1L+E4A5eJ
/AY//bYQwWml9j9rdBGgMH0BmwPfx4mryoY+6TEzzNoEInZEG/Y2LNGQ94trgYI3
7CScTuaNBPb337zK/TPYxMpX8uWiHtlswCqTIFwOmelNqWdUB81doTxvJskFFnoT
xf8M6DWCMeTwb3YpWlwK9SNNe3fdOkZ15f9hYB+h1CEoUMYjuxH4rUZiV/CnQ+LV
AQtC00iRBTqRHnj1+i1ye26WxCBpRpByMXe+w5srB2DRV9HJ09gdtJJoHkqnZO78
4Kf5agJ6yyyGE/FpjuQqpbS5VlUdZb7x8K2dMexSw1LrthDDvv+LPVYjV0+OqL/F
0Lb78fjcuY6+dv/z2dP89QaRZ+mqfSK7pjixPE+NYTusCTz72WIGSLRKzwYtPcX2
t0N8m2Zp5O0OoZ52f8ncLb4KF4N74K06HBNNo/3basSbQiraLd9a3RW3agy/e6YC
bKJNt1U0093AJyZClJ+gLwfMd/KuPCRllBtTMuM0A6rdghnnlqMh5IEED7zFw6f/
ZZ7cDYXIs2w8q404e3SqRivsTspRm5zxGfTy00T92MXLgB1IiggkCVThSkuNhZmi
j+Za6fGgL5A5+dGWqFEKexPX9RKPNL1k4bOazL9d8/soNqjSbMDKXWWd4kC36sX2
U86V4liIvc/pkgcHk3b7Ir4u9YpCFIZY+jO87l5AJ7taokh1kK0nP1DWmBDYtUVS
cWu+1y7vQj9UwnmpansE+lMqszHoYEyHFKAGAnfqgspHJwMlRqBa0V+RwpNrFrS3
zdR2NZvr+y78HZ0eK91RLgsYiq8I91DR17r8xFTs/f8TX3b/hqMrtpyDJIM0BFTG
OvIdpeyqatQZZ8Aunz/Uw5lwAAqhIkyM9EuVQqpb/QyA/Cc5brzNvr/mzXmlLO/f
JvGHFEWwTCj2xBsJDv7Sbw0Jg7uMfkpxleWv8smOivuDjAyuPeMW4hPhYQwSrMO7
JMulN7cukJnO8lg9rb2FAqfLUYRCnbYfgrIhW8iniP9bd6S0ipoNyyV3I/V1KeaX
WU1uGVS9U0kU/Ott8pEwI/OJJyvjHE9dE6bvaTdwGRkUHuyekeJ/MBx6eEWiYB6Q
hSUwamJSi0JzPoud6yprK6zHIPgpvu+Cwvy7/Hup4MEEdXNxLvHY5CYrHo8F8lOz
dA+sW385HbnHVGMMrO0h1J57Z4qAc+p6z15zwaCAS/KPJBdD1k81LQ3EYQeCUVAx
aVuoPHh/Tywq0bU91SW0ci+RjWXtdO55cgZ0GfAcPCBiv1Q7Ha+OaLap/CCuilzH
uoY6ustS5P5pPiXAn7bM4YssPhwxJQ98DKUyykCrIoMtrByKcPmSLArwMMl75Mo3
iMEdxiKEadnlCE+htfBc3y80/GhXlf6xuCkY45FFIY1KNitT4CINykBQcc8puTW+
QrpEYp2LETXEz7769/J7gJJyexJ6gdnVfXISWPHyq3LqIh56Vs8ZTU+wbnmvMtls
71zgyHXEdTjGa347H/b/wG1QQRRYKXNwiQPvmv902ADIkuP/z+0c7A23XK+rU2Bq
e6CERkSSAmpqfoBfcMPjx1PDiDmIGwzJpuTVmGxqnkwgTDIZ9UrAQCthkdFVzSo4
hP+ixF2WzNvjsxFLSyAxxH73yYwExbGk6MDRmYGQHIBFcvcVDSIp8KpT8cTPcohb
+oxT7WJW9KDngeDC2iztgV8RL6qe+V/sNf6+6o2QBVHRycQ/WpzkLsLSGJ5ORyjv
kVqniuC/M0iJ+7cKp2FMyKmPudFXOpMqaCgzXZb5NxqOfgLsRjFWuuoeNhWg4+eo
vOHyRQ247FUtxQEr2OdZIEAiEW5vUiINAGigaya220Ky5yXeH72QUs1Z06FWPYnS
cu35jCcgDtOEFWbCxh8TSfeaCViqvjk/zCta+xS0ntxK+r8rUmKx/D+sjTVTaG2E
9Z6Px1UxrimXXTgQr3UdNKTN+YQqgfAar4W197+P8bAjFAVIQKKHmmKLxWofoMz/
rJc4UzeldwzOcd/1OfmB1h/MSa1/n8b4RMFw2ls9LUVXNIaASJ4Ut1IBewGlw0Ox
bG5LO04ZG7+qu9fX4jJi1OOfq/Ahy9A5Ne8kTRxcnhnz46cgyk9UN8hFQEVfF2uv
1Yat3pgpPO1yJDntxFyJtwMW3Lv7Mo5W0+JWOJQmXbrnDVak6i3Vx2B6RDysFZxN
JDd1MyMj5Dt/hy+6n/xkHC8N189nh50mMeThpPuS6n4DtWTtotIQxX/wQN9yIidh
aAr2yyASLXTTbQWVdcdUNLz61kQwIf1R3QbES/VYkNEp0EZ9N3zmCsIOR57xI6ZU
RCUgNI5+3c6YukaqJ/QKiiSYzerluS899hJ1RaPHLsMtRit0PMYUw7VZqrzbWXpV
sepTJi+c0R4aiKkD6lpcg6/Wn464eGXB9YJuqppnxNpR3RyXUEQWXfXPh+uihArC
ofJfoARYKIgP2xPgI+b24Mb7k7scBg9J9zUrkWkN15AyGSsx1xjzt4F8e9fyx8gW
pu+E0q8Tw1TJ/DOqX1tRdrECH/CBHjONJ6gVqegsjFB1vNkEBlQIRKnFwyDvbKot
RmMEOEUTF9LrzLz7r8CgFrenmekGCwmfKxuKCGvxa8zivG0Ruu/5cLK9vo578D3j
2UleCvZcxEJ1bJJKdA6W2ipadOLH2DiVZxWzvzRn2YmjOSXbUnXOsD5CBbIrcHNP
nWcog6aG8zNsWmZhIQWDMzT0YbX0U9CTnwY2zMkHNuTbv7Jpw9ZLO2DlOGgt7iBr
WXpMkL4h/POisfqv9OEQCeavzGp2g8ArDj+N0/i43BYz50sAyqG3FG14Ii6ZzhBO
0p2uKea5ZLMpassjc4daXF+bcjc0P4BP0r0MMLVsrFU88vwAJ0fS5IvOTBcgtEY0
lLY7+NcETb6KmbF/Iv/42WacHMMUuB2y8qIlbloOqQ6uabt7HTbfEAsqH4+qqtN2
ynXBBOE+dKQM+86/Tm0fyV33Rh/V9ndbCc1zs+Ap9HqR5X/FMEVjiFz1HbtdedOX
ZCHlmPkFYwAlgYwpn1bIHMQtkmrje5zIp4RInM66lVfLw8HqmMWSFmed4Dc0BGUK
ZmLhN81dNaHmB4gknKnim1HBxCYnttI4DaNug+URuQ0vkvP8qroK9vb/1Z+xYM3i
Win1zMaSytCiL5k/Yb1yGJTGuvTdvyL1r+VuBljesHrYGQ9KPFUQVHCAtClLMPp2
LN2rEfaCGqjhpJz7aIGpKIQP5biyVlSLa3sLo8NoLWY/YstANAMoDzi3/K1TbHUR
mISvVwQOUvNdt/q3mY8wwz75ORlsuBU2fEnwBLcBPOAePKq/m3DKCqpexGALTc6R
CxaY6/9ix+k6Ui3/AWD1+OZqeogiDIUanXYdjaN2VB/6sDuHySHQ59xRoagy8BxN
+oGf6l3iH6iBjDTzK63Wy7Qze6jEHVXKY/EZozNg5Yi1oW8/W4Gw9NCIAXEeE2R/
1RMh/rruQMXLVij5fyp1+uoukob90J0UcAm6wvtRg59Aj4IhseEwNND2FGNPyDyZ
EngqgNeszHx3B3jMF1INJoyo/M7lyTSlgiUfPtgBwYSG3bu2qk+mqqZpL1WHlQlA
BdoxznC0HZcIOwsOJOvh64x8sS0WFEEAQiCsbycZp+GILgPvT4WZRvHOYfrXmKNl
xXHJDuEEXkRefPqmQdb8gvgKFVZx+Ap5jqTbCIZ0y8zRPyqEh5c/5+Q5vkwJQaeR
Ni010TaQ1hNYhIAoBVIzPlOY2vQynogw+9MKO8WJGhAkW4WIKUTKBPP5rP4Fyu88
UV+3pgEhxArBGiPoEPO5F6dGazaK9gddvCrEWPUttANwEHzrwGUGr09TiYewgciu
tQZjOpZlI55cVIekMrgFKIXQvZH9VQH5fv3IkB7Ry0KcKxzMB6GTYLxJrBIZhvLs
L+VhhI1/3P8cXWg3c2K/ItTpXrVMXhB0jyL3YEUbPXU/OSy4J4KMAABUvOXhnvdH
ZG3DjiJVpppk861rPDFMlv702JQUPH/G4944eBiA4/CjpZviW7wjkiPpIjh7vgdm
XfMGQYl/UKrEE/NHWl9IBsRTcfR3PD1iUposq+KIW8EQfukDfPHjAdmbHrxSnOPd
gddemfg1JywGzP4sip21juz1X5Afyxr0m+R+1d0Bmte9YPas7z9Mo0zEfEqHeQ/C
4G3egwGWObkT+HgFuQlXsfU45Q+WVLNaJ0baNktatIkrXpKhz6DfnQjadnW/HlRi
cSAzjG6C/U0WXBc1YuL0aHKrDUzJ94sgq1tJqygAEV+C+r2S9o1441flmRzJtrsr
77MDlTUgvgMD03va8ePuND/svy7ZLNa21E49nSgYuKl6P33OIZzjMGiuukbM4dOI
SlZYMEXLClEtimVVvRb7QbFvcGi9DrOnZK3tgpUJprmLRCEms5kKQXhXn5oGALNs
4hsbpB01T0zCbSJCy8oTeC+HtwHXILM+L2ZQspK/g0EgAjD8AzOoEfooJmJGITn2
VLmMneDR2CjGH1kU5QrYcZ8U/2E6S7qFeLDn9dlPso7tb3GEnl6EvDzO2BjZkiTy
MGhLqTgiY4ATeNihlyX67IZKLMvmMtsYBbdr0m4t+cHqY4VbTw6qiwkaOXWSdJTK
/0KSPoDpbUk2vlIqgbXOuT+DKw5QdcTCo41ocsSEDU8eF82CwhgFCbFncCU1sXNI
rbyvRN6gEpsMxe6XeETfB3r7ckcupvLesBrbR2/JKxeFg7Adf3/WunU6LpQxGt4K
pk3foTESOuz5bChFzAGytNyfXdsAyXAuR35MXV+kt/fnbeQBX5/18Oh1D0aAAeVu
s9yyPyXeLcGTiicN6CLO+7sBiliuUSFskZK7QuDb+h8pZ82/dTd0greBxTvmGNZP
l/hfsEJ2uquaAfBuztgaIkDVaJABI44DTgvoiGG7ZAanR75OmwnR/9JMfafI3EHg
i2hXO2TfaDf50IaL5LbVxjWRdlst3e1uenKPFJCkwS6USh7b/5lRDmb8lWOAtrbY
ShGm9+MPltlFbYYMYEf7lDcnfWep7ChiJfUFtz/QUezk8VNvP4O2RAzA9lSEbszk
yOcy4G2WPlYudr3AbYEuSGzwF5xI5NkbgBrIS0ZmlF0px7z1BTnleuBmA79OLQUw
1BWTlN4j9XQ8cdEokt5O9x54se/zf9+11Mf1XCBzrBcYwkh2CpL/rrdcsu5kTgRt
esmw+vpFLjE3CTSnYqHpaICkO4WOzivfxzbFS2j2+5Ppd1qtlip7/dGSOP5l2Bpp
bOnKqtbfxoklcuZNbx+ko9/Wa7VMBNmi0Bn0OzDS+tzj6u4+xfZxtz3Exc+TUVxo
iSxMCqoZjqppawXD90dC3GY2NzOK+CkYA+xFhcmFlGgjB0o1PuO6Ik4jU8s7xcJT
RyOrslMrhd/IWhiWsfLEquMWxT1m/AuYxuJzbZcVLNzi086XhY8D29ocvS8hfIkN
gbgiqUw0doIpWyzeh5mZZwmv0L+TAs0Y1cKrXO1TR/bNhnf9UFJ7HuaAwRVUPV3O
ZYgwGTGJwl8Mx+R8x6v+Fb/PySn4YCZ+DinyZscEZVmgokTJrIJ4mk2yqOPZdq1r
t5kYKtSlJWf71nv1uLKiq6U+YBmVkhb/GqvlFMpRJAA6nZWaxW3lD3QYL9hHhi+8
U4nxbhwgjuJKmPGeA7Z9Y70dl2jJi1W4TLJiYyI0RHSrEd4Aua39hTaalbRWgWsK
4l39ep/4EY6EqV7ZOYPPAZDL7Y9WMW/K3J9IbdeUWkFzYT32vHDjexwBlpXqjk9+
5RAl/fyoWrhF8Ovq9MWdE+IhoTSAUHfdbXoTyrTxIc8PlpXt5NS1Ua5CFFLNU6x+
R5aZuGaDElsT2dCDvGPXNjT85sj3zLBp0328mKeWO+a8ENJ1td5CtshBxjMNsj0p
PxuJbhjY4DXK7BAoRjxIUmNvJG8BAnt2CCUcfNA4JJny4JbElFNDJOHN0H0Mz6dA
qYIepLdCZFV/4IJLx1/cNbgn4kLQkYdlB7BM2VDiHFPZzPT476WwQUEMxmMsQ/Xf
aWC4fDM4juVDBn5XmgjnM6QEHCJ5RBpemNuclQcKyNYJ65KRZ/irBpntMoGxua/z
3rPtX04tHuo1JA1e8Ew5diF3qK6u40j4HXUSGfFhkKfi0mS4X/tSGw/SItf6GQJt
mUVTumF4sTBoMEwJtWYJ4VxbO+TCnObdvJKE9tnKl3+R+mcnd2izJcaG0havrw9S
pMzmGz1PCFctQKgBxSI3Z5TFaVe8os+G7ZbJE1ri4lIw9J0Lxbx7nYqKUAC9HopR
jWO4+vWHzDn/y5vH+Ya7zhGM1tUA18D/R8EhMH0SEqp2NZTBATe0Xw9CiAqf6Zsz
zyjuyxfejorzklcvNRy3WaK3pXesf83yYoSukQcQXjQG4sZs0KNyKN9sEEzLx6qE
+vploPZc8rfyFhgAvAaBSvyl4FVyOawLZDApwNKZPpn40nIuJNqhmnOlQeU+Bihm
eD45FPHzOl+9fXmsgQqMSKgmosjwQICwbC6AimlzdxP6ZTjgmkq/mcvepH8hskMb
6SrB3i8MeykPhf4nA9TgnUomyRYALHSRyxobEi/6SOKeVB57xXCy/aEqXWyG5znZ
mbrdHBzVyDMSaX0sv9dRJ9X5BRE8s3yBPBm3Jt1ns4jJ2VYSpaW8moVaHt646lJL
iPN1AKbYVxUhk1ZBWg+dn0edhHYQ9x+bvMzVrkdT1YBzXHyFLfPR1PJFNp0SPQAS
+ggvqCM0ODYBgUnX9ngICx6EeUYeJ5Q4IflVlDtse3XMORudsHi82AJBavNTpGdP
0191RaYi13JVYfpcr2rjZ7ANJ9GWSXhSAMKhUffJcR39rxdSiJkGD0UoD1LzINwt
QLKetW94ZidhbUmAI2EcrdqUFP62Rwm9dF9dCAx8bQh9dEF6cV/9LiPhu+p/6lh7
81gjgW8pQEGTmYvUWmFgs69DemsOV0XuRbZx6wxRj4O8JKCxfFLVss8BWBbYcwk6
HLSi4UiQPXNLtmsTDvgeo270lqi1jH/rKE427BxXa0aKNIbgXENTZ8SA+HfYSEvC
3lXYVMVpu2siYJX+TqR/2qyO1cgRIUyTAZrcIhpG6jVyFtQT1+cwWGhkl4ndSznQ
3ps6p8JvPH33jnfQKaczfwUdL6WHjQEFxS9KpNYBZ3OqmbUOwBsyR/k059ZTzuyy
TI94AxX0TcquxuVlPtHmM/0fuy5BRNTKqLvuzHXNFuz3qyVdmpv/Hd09rsBo5mmF
SnzcFKJz1X3Cr6Mwy2PCPb0qqoeIUOZLrI1slkr5UGBW/RUYVJ/YediGHvx7m6ih
l/RNKjFrae/id8zDEWTqwTN+BPuyEPIdY6U3qteHPjCyNL7OL4Vx4D5RJ4HPVXn7
cvGQpMwCBaBRejCt7Pmv+6F3RTnpvj7/r6QSmNdko5fFv/StnaYiQlRI9oiKkXa5
XdxjnlVw635x2aRA6nKyjBdOWGbJPpruORBJNHwIslNi0MhhNoaih7Aa5yFQPfGs
I9/dIp7IlC75FA0DkXYD7WYQTiS5s2UI1y1U+ixCb0WDRFRrH04epD9KWVx0fefC
1KyqMsiMbjWvI8s9aGjToMYnWlFq4o63oeGvzfe2WF8x45jdcn/aBBunROgYd/Ff
R/UIorKe5783ZLNXC9rvCbBNk9V0IoXl+DltkKxHHk5X74OFqZJi6/GgtyJ/hfUL
r7Ml3bUihLMjyZfYo2+q8OBAuTj3W6FwJzZNDEt0DumvNJAtAlhDCD1et78t7bOH
2yvz2kOkxNKP1Sa9X+qwqQ9o8pEIDeZyMml6s9amjuraR/SFCqGht5jCQZ8rzF6F
GHc4NaPt/40RHqI+T247P4gwqWPNumcq3ahNJrJGTBMPB1JIaaAkKFnCb+4tsoJW
p4kl/VZ1Ix/n/CBEJ85Rd9DvgKQPpqrpQFhgote8UPWhckc1hGekw/QBa/UI0U5K
ISLy2RfluWjM6VF7wkZYyA+CLzzd9OgKDc7OIk78E/cIla2cBAPFOBq3Ym7GNXaE
DAKFg4Ecl0avmTgfwx+7APMwChZu2xUynTSceJpJ0jq8gimRuC2md8gH+o3A0w9Y
r+5qoCqACMvy/JzskEsW9BHvI2+wplSyqcX43HsvmoJ4sTK0P7R4uPP4E9ccqDOB
Uu1LQqZXr8qKOUaY/Y9IB2YNabbSS55wSHj/tsI+33pAXkRDbS2hIPSFFM707Cbi
ZNztNO9TycTCem/ldUvMU2+/B+avcqqovL37yuBgEPYAU5/1tp8n3GSZ0dbjUYmI
xmCAO1NwweKFKY/v3dt2CENKbAsXrebmtqu3htDqYgh1SHGrLML4wcf2f8KtQZUw
YdDnOtrSGsbm5QxWN3hbSpbUSCYaTQfJWQbNPOkLiLhIoD9a6Z+R2AGQvO9GNB4r
+jYc1KJQCYEpzbVS1oGOydwhgcflV0fQ62YjH7wuAaf7Ee44+oIx+vBSJv0WrBxz
NX0lYYMyzKtm3Ila56tLYk58W1sDrmCOCM3lJ8KMJPKw36/y15hnDUv1ApIHnjYc
YhSjaKoHtEXvWWOOs6KyhC1km2GJNLNQgNvSjTzj3ylEEdudf2I6/DVenziAaJF6
P2sPRZGh7jtyOQkfa+w2yT7DDRNwIwgz66C9TQJomEq08ikh5SwUS0FqlftQQ32q
GxvsjpozcZBMwC71pme0TAWFL24VHHWRA610iIX5GZhYamB5/SJRu9FlZcyi4tFz
dJFq2wsxQDry0rTGhw2o/Qsznuz7Eppbg6lerFQ0DakkXOGgLC9cVmPA8fUdvgCV
9pc+GF3eR8vkX0PRBDJtouTwukCZXcRSawmHp7+BLxG85/ke8l93uP92dD3zYTYU
bN+/UysAZ3GDu51MQc6vtyJhKfxtY35NcIp3ElAZoSftuivtVXdi2vfx8ARv06R6
PkkYPTP1IC4xqc7OTBGqEq07cD818wojR+ugo1Em5HuDN5xKeGxAdUKkvjK1xQvv
W/UUf5GhhApw1gf5KRDxbnWrhaqAX9smetmh8BWeR7aVEyHW2rPz3atVu6BVemTc
XQiNBqMNnuJKBG4tJ6wUra3lkBe73TP+Vyg2IzNo3KoRmoAi08aXEKGSg78TX0Yi
JNfPkdRWmPKi0O1iaQ71b/R12WmaxkItRQpfP98gcAEzivNKURs5UaL+X3noGBYU
ZwFO6ci+YRCJpfdNeNjBOHaglputPHel6tMVVldXs7fKbuXnJPakkSR4kviRqL1L
lJsbT9ikNx9Xdd+9LUatxPVUSIfrTOklJmu+cw3fEnWe4OEzo9EqzC+GHIPnXPkt
Wz0q1NP5lKFDrnsA5AWPna5HXCJlwObkw4v/HFxTLk0LNiODcOwUHiRyDAqJiw5s
ATN4oq1SXOUcHbcI33VIjdTARKdz/XIRXJokCspWDaKdQWq0tW1z/388eI7OLX7h
lSTgtmfHMaPXxfOqRxLo3Vkl8Yrr/XBRAnsQv8xDRtVxtfpdnnKmTtGKzEomslc+
GHjrUTNXHPYPNAGRQk9DbUDQmAu38N++2Yna+gpHNiv1kgBMZolx0uKGE+4o0MMR
97HfIiFS7JwRMcj28mnZ2wHIScYMq7w9tum1/hVLdcgikGVtiHXm/y8wp091YtR8
H4dJMZ8/4QEk044UYp0ubWeRPQ6p5mEQ5IJPxEuHdy4T3NypG7BiU3QZMpOqCxub
P5/gOF2diyc0+27DVFqcSeYMcjSCrJR5XjawJMh97HwlABWLhpRbTXyuoHXyRZ+2
z4FTbjcyoKkprNUiUtuvzToJwc7ymQv+6LiE3mhS6Y86QxhAwMalqsl0c5zu4Y1/
CHL6IVCpuRpVBjM2aFGDMKYmGyp8crikvjkDK5aaSB2Yu2Y/BMVI+yZYksun5ShP
l0b60oH6TLrFWOZkXbzqkz+o3krR4zZkizZ6w40/1AYzn9gpSPz5gnMteqBH3CHw
xjr8wU7BAtmiRni0pkQ5giFOGvgWqsiulYQwjAOZHpPOzBKxNNy3J0oCIUCTlZUE
MZYOlwcPBSdwsiY+TP1XTEyyAiq+eE3fRGwf+qSF4H/Vc9S4O25HGq/REW4OpwiS
UR+XAv+uwXfs97WT1VuwjKO2IEerNYsu1leg6Rjk8aLnZGVsafglpvPIPBub9d4Q
Sm0g9N2KRRSsQ0IRb4fsM4SRu83jaXAZosrXpPK53Hvx/xwEleIuyxccUD2yR0tA
iFqo4qatgb20qgY9zguaamZxdJ1orPhzgO6DdoLPyQ1FIqONIUssUwrwK+lYDE2L
+xh+wv3NPz/9qB7nKO4YF2xsjyknPlXXUz3T9Z0IG2CHrmuImJHn4B29sTXv6x1F
9qbHuwGvM+zp1w46LUfGID7EOu1mx3nsEjfZwi9H7pWl3dG7WDXLCW5wiZEqbfXz
yJ6Tb1u0nESF/A+mz2nDVD+1wYRjGjrRPU5Pbr8aGXbKaFNvpmcqAqadYiGjCfmy
SUUb10elkzy9hIKs9eJB1wH86zLyOfH6fI26fom0pKmrLJXML3jPAfSWlFwAMMtM
s9QNKSUfqV/ED0TBxJmupTwCjFVPDHcd1Kqzo4x4NgDybyloY6AM9o8oVoGpzOnK
c+MOMcFn0ZfLcUn+Zcjd9WPpALUei7Jcq+BlZdcYZwSoUX2lja3Vh6HDFnn+Rdxh
bivVdaQV5LC+UZFMP3LNONd4ghnPXy7594+u4aj5JfKRnVx4VH1s9Xm7Fjb653ie
Qn90k5qvibZwV6dBVIg2jMg3epoZBnTFB407MJ4ywKYLU/xX6pJAA4ePijo3Ja+B
cNBBdrgp1n5jpK0HfygK0ntxQ/s8GeZM2RbnVG/M6E0AqiVkAQVX4RYgzJgJ0Lrz
lXrKKLnxY9rCCzvxgMEoRxcr4aPaVLM81NV4230sZF62QLoYleP9pU7WdhmcgjaN
QFsaFjoS9FC6WaedBcuQ1TAezUeiv4pR2NeEN5p6/pI0YK5sDwW4gS50VjX6vB3C
1TLlV/J28Eo3mzNjshmkxovSF9vHDMaeDmehogZjJM1AkpRXS8rVd1ctolK+M7CQ
LuluPoXlrswf/p8KmNROupLjCPBm1guRAl5XneNoDjL+rMlUbXOjZ57Yc8spMpkw
IV6qHrqxp3tZNK3s1BoKVF9wDYOUGE+MKFg/XDkaZ1M62RcTzRjzozH07oMayEKB
ECD2KAy8qH2rk6ZmIoCDfu8jJdix/lW1vSGJmnnJ2C+kNl21ZoBEzaeY9brQViXr
9NM4Lh7uH9UekMrt/LTWIXXliWQn0haSau6hxvUa+oS2zW7wTEbkTZkbe5zJgvaS
qot0pm12OZ93LhI7svmwdrF7hRujkaaXgHJaaegDrc/F3Hu/nwvTJhOnBaONrtcT
0u2V1ubCmOlxOZPxRaaPlEmIIn1hDCGSmK28QCo72rmMZHXiFjXjpiKzrykX3FF7
xaLMEZuspXmTl+q2UogKvO1xXXbw7rXXoVjz15srgUGhTCqKY4F3M3jC+9tEPfJg
IEWzBE+d5NyF+Bgz3wK8Hpt+mNkaYn0EPfD6NlRZ/X3kYWpnCMkCAWAQs3VzHUiY
nYLzbbv/Zz4fHoJj32maeBNv3zIX9kr9NivLuYInlUItWuROwgmMaKmysuenqWVR
Od6X9jlURvl1yZE44VDoRKQfj9eAOon/d6easikrbdT0ZRBvq0zdfraVqR76CyX4
1uhQP+tpMlpqRvj2wXl+f3i+IWavqQi0c+QEZj8KWPyqC5Nlwj0uJJf7RR/JAZQ6
cv6MnwCfj+2cqBA5N5SBe7YCgZzu0R1ZmVaX7T08lJ0kamz0BKc1V+CRM0iEvJDF
dy6PnTU/b9fWjht8YUR6VbhJ7gZhdnm8fVZcHS0fLQ81ZAXAEqOtmlLy+hzGRHtf
RbLOv6anNAAkrkk6zxXJBO+be0TQ+loKRciH47vN6GTdygNbUm1UUi1bdjZh4FCH
pAWn47jnDgW8PCyO9/FqZNcrLKFigsFLAJa0QfnceEjOzHEcG5/Btn9VVBjpHH3p
kNJ26Lv+awdsuT4kdM6bG15Gcb1EKQsJOy9IPHxavlsal2dDu8VeFiMVdabZMYGT
sA86eJvY+C05Ny8eY2NdpGJRQuLyjX0iC9cbC2olxqbi4M1hE5cDdm80AmR+HhxK
aaie5Ovf3HGtBnDhaCMXGjv9wDvb7gYJvF/9PRH4TBni1X4IWYOKGOxCe/DBx+SY
wZrEiEKusYLDMpCbzbDxlsL6M2oTqB4PlIlsGlvdg2mPvxBz6ZDvjz85xsziCEYn
p+WVma1YfxYeZEYI64urvvivGiM0Yohl3wUJEVvI1+U25iS4gpkibE6REvwMLx31
V//o5N25Z1N8WQ4JPLNhiXj2gPZjPOeaWMKiQGz5Y6Bic0ufnya0jKdBsKyTpxKT
eu57TlRlySMbk2ODp0bCGC2jM4nqkeR71aPCrFJYa9OVf/zN81/qvdkGyoZfRqz5
zO1t0dJu7iRUqYmgDbJv7JugxY/fauyTy4EvyUvBudr5I6h4btp6b6SKxVx6lw3y
x9LLmpk2S6WMKPZzuu9J2e/HmQEsg7+pkQxo+BkpCHcg0RM5qBrxytNsG3vyejdN
vFpTaBx687mFY1Od1f+t7f1wQZo4id/A/azwPoaNhBXDlKYFTvuKjmmtP/Yce3eO
7fcp0vh95yRWbchBTkG3XQ5/3Z/leYDR52Nmrz2iCLf4wrr2xe+I5PO7x23SlX2j
H4H54/JWOgmrE2OGYcetgP8YWGlnyVmyXTojKay3phutSAmDVTHrrvjBsJE5+/RD
SRqqJtLHhHBiEhyqrWv+5Z06IT3O79X1tbkHawhBa4Q5Sp9KWtZh/jfGXmnu2sJn
6vTLXnwSUeRH5EJtcD0IMxZV5rc2QZosYKi3XmHx4/H7lYxlZNi2c50st1HhFO8p
p+ZLGwouHYC4mElXlaCbZ8R3oqD/BNb6eovl5ZRZznNjRC7En98CVhnSUbM7aZJu
RkJi2XR1Y+iOVzwHxRabI10JtDwEEbvSSp+kvDRsvpgYgtHOYMbuXENNZBsjwun9
Im0NczZcOfRvYdn3UTxxcFCPjDeIu3o+I/ooQCl75QRCzbpnx7N+CYltNXWyBh+Z
/Wg0y26tV9vQLT/3zl8llXiObWovzN0yKyirx0dGiqFyc81ebSTxVgw8arYsnLdB
IW6984BYrq+U9GIWRFF0ds7rmTrkqcRhqLqW5JDDIZIjsOZ0U4GiP8HgbnPeRBav
Pz+3KH+odP79WSe10crCxuFK3u/YmyFkr8kijTuEMXUgAqrB55FWjcZdx+vUAio+
ulclF8aCQWkbzK8OyjpdjEcMznLcUjt7gwO8+maXKt2gznrNvHpDNgguR3zFhfjv
vnmUpaVIcaAKKC8ZsK4n12hJkdKaVXnwc7n7eE5o0BF3Nbwe0SPFA/pfM3ZG9R2U
6xiGo4C4wjn4dlHyz3jcMdGOJ9zyFRrpbLR0uoNYixe/a9ajVyYf8b83SWohtkOc
DaLAdEvsI0xKIVqKScz1F5R6izhtmSSxTSuZJqMK+DnFw2Kk8l/i1jZgaTOXDp7y
BXoHfIFpokXVGS4uYX09tl+xCZbTUGDk2d886tCEysYMLMi8b8Quey+Ka84kipbB
srRxZ40t3hYNMNvgKXwVIMvigtCrWjWEtDOzRsMKc/STj75EGwnivyNkNh1u/RpS
2Qz6elKb3c2Vg1zbSqtHCYqmRnpFI9VtoV7XUQ6HpxKXSBJilfquebKiD7N2/+Na
/SMmAw/g6T9iCUtlKC1TMM/NtSLUhjefUjJaDPWRqKCsOCmuLp1kxD/aC0e+m54Y
EEu4RceqiS30ZIrGl1VDPjpdtmQT6mS3LEHMzngmP2Z0mwp5rVQkK3gqWDbUqAYH
oq90Gt/RsMQ/UBRBxtmYVu8kEkG+HaVRGOJTew4SC9Wtjeg+pBxbezeQKAFjs5IF
OYDFo8z0W3gdcHSrkTQ44T58LWWzlH7vJPhv30t4A4+SY5bbnY8uBTaTgSwT7/Jx
hjN8I4EtR8ZO71Ue812vE2g99Yu2q5G/HTSgJBds/tWRMp07LOWuYLIsP0O3PkUF
lQLXYd3OuXcUs4MEvSAhvPhwz8VyjjhxSbi1dMm2SPyOilTBcxz/qw+dJeT9A3Zp
o/y5hU3XiyoCN7upj0kt9X/x0t8wC65O5V7ZdIkapDKXeYTtkmwWzVcYiZhZtpUD
GYmNCcPgn0ViUBtzPVWPeX56WVVIi/My2gwG1uIBq5CLg5cUARt+dZ1IbhDSBZ+Y
hMEs10LfM+ws4d1h2CgYQI+kuGWtA61NbTPhvF1qbySsLLf/5G4tayoztIgSK9lM
H89HOms67v5rPAlEQPGTwAiVGLqkkSwB44AGnwFlNtB/PthgjK6txr2W/KTOU7vN
HD/rnKx1nfQxfyi9nx8pUquYRy8PLipJTXCWTpRi/Dh9OANyx2sf7FZ6b5Yt925Q
97YAytZ4Hq6SF/KE9THpvEkoe8h/jsX4mWB0SqIlb8Q4EFgOzzCjYwiER33dKNaw
DDeEbKRmWXnSIcU47kQLLN42i+TYC//EXhajF0xKG493zQZOg5lQfgdSvn0rTWVV
nZHxP0LlqkjjMQL+lsTDK+HHCNLaVU+PvzI2Ji5Y7SMgbI41I2L2prOm16qwzhbf
m6pa7MGKYtpniWAEo63vNb0iyLaxEy8Rmb8mkbCpW5td1Fk09BRO1h1BgthTCs5M
XZlh5s4qCGIYz/W0AJYKNjbZcjCiInuMHst3/FQ6uC/jlEchND74QhuGK5+/kQ7n
qG9w/jH9RWe0quqsWcaaBKfLasegY55/47Re0d6dwOHIKkQv+a2ELvpCiwuJJm6Y
OznywwihpiFlwDRrnNoqxBFQ6nebgTw8GnhmNfafoA5k3pL0CKuA6EE6IYyJ+gZA
GOtjc6D6Tg13h4wWTDtNBsj356rYEFSgdolzJGQmvGnalnwF+bepGYrjM0ZoIUQE
nkqQR4dNBKgiYUWDILavzhJUKyHQFigoqqwR7W0zuuA2j6wwCI0DH5SO0zcLqusg
VE8rVRrtajw3LCoHS+YZPZm15YdmVGM7Oh8kOCG+zgeK3KH68+7rXd1rZmEZnTsM
OfZ19L7K9C+eV/IIBDxXhszGmHBYpvtB24lPv0Ub7pclRs5TXhU+UROyda6jf9bA
yx+yVbIb8FKFLB7iwQfG06gsBHSOpJu1oZFO3u7fMgnjEjZ7opNSrc39He2rn37Z
DSHhYRPDt4WI7ylQ9NJ2Sfjoy11BnMomSkQYNqPsS7dFMvONQBK4LtGmY3Y7BHbP
ihu7q0esk1T0BfjwGjd2YCN1bmeDooZ+KM9B5yoxevlvtSMyN5NqpPaebKTSYbr+
San6EpV0cKNiiu9NXo7tB0takOwr1/L/8h5kfIjjdY6JCjdc7yNjw+BY8Zw/IHm6
AI5NfZKgkMaHShrKhsTnx0VI8D/3ft8TDhofnuRP8YaFXsmF3Q9y8s/dh6OZOdc1
K8dkRX3+QT4d9aJq7WTq+b81a3AZMGyalFYCUV0LZfyoozd7TekqdvR1U0CjWRmD
tUSb9tbX/GTt+s84T7QPRJwXWMlSuqcv0D88OkrfWGE2Gmoq/41KvfRMQ2rdGJqP
66GLpMp5jQOYKjatNZR3aZdy3UUNNxeD/X4yrCST/SknHOpDbquXbPaRyb4EE2Jt
eW7Eszv5L23I32rSZ763vimrFytQ9kHzJs8HNkB53WmWBcqN2qO9lXhfIgIkBYrV
GEyG+F2AOrpsGRvsBMmlNqY6iRBv4x4Zq/8mkBXs9aycpVmUPi7HwQGUBKPw4rwk
9apEdzvMh6Q31Esjf+GnfjX1ct8gEX2igX66lDrresYoy8Y5eNQW2MPhBc4nWabh
PYsU/n/1E3faKUHYCXS5Qo3iXKh01yepAPWEkLsCm7bS6u/TESD/F2TswYQCPlgl
0feIw9Z74C2Aw+RjITr3Cd416uyg0CN8xk0leaQpTutb+VNL0gFxjZFGAH4S1agk
4+tK+kfiVEhvgF+FHM2VvMLCj+zruf7BkLZDjt4xVRBt/G4X1QKyqgDKDOltTDar
noaFveVuwheWy+Cpi4O/fMbTQbYBlI6Fk8T20rsZwi1z7WbmTokkhv2wipj8ipie
NpnNtdKoKUW/WpnH8mVCkT299kusQLCs0aQRTpgGAonbBlRB8Fiu5qYB2zE9gyrQ
kR9lrRXxvfj/TqstKQfxMf3yK2J/NHwA9u0Y72n+eA2XDf3x41lJv8Mi1iNlElPD
79uJdxvJt3l3ylIqzLr0fLZEeEdP17+GLslnhEYDgRBKStLeEhys5v5nl80+ePNe
oCkrWzjSHiCcONXIY4g6XGrBygeQOz6wsG7Hhb6uRVZFKpsUaQA1KnpIBUhjQmjf
SKVjFFY0xnTU2Cq2LBaBubSPvPomv+mVw0jLKo85sjAz7IKSR8lHZR1uVHUcHR1C
gUTT4fMyxFb3cgVR02jIeAu3oHyKDwcRTh0JHKUN6BY3fNibwMmSfn/i3q7E+vfT
F0ilA+TXC/pzpb2jTFEp7aMb+x1Q6a9kvjTnorpcHSCkEVBZBjjHafJHOqhfeKhI
ldDnHqcyplF++MFBZBqeqUT5XZ83caKcUfePSjmO9v91+AZ2ENjJrtViViBz6TvG
81pb7QepuAkzjuc2HJ5lMyJb7jX5zrJSBZEW8etaINEZklXteKAZSLPizSGcCZ2i
WOETxbLPYTXvNMXswuZseLxmtgsknQmokJD/D0Il8K5CHMNXEnswpfBNXADiK7i3
JaYbop4/gZcFWNG6idpTw20NwUwiLKlPkucJCSxOg/9v0XDYDFtnlQ69I2BKe1uk
CeIuU2FA0T3/WE+UTUMFjAtGNeE9Lqwo/ENRs5Szcr0GAE4UL+B3DHxwjuEIL3th
Xp+pi8uhbOOVe9M2kxeBaUZNvIjmjHXO3BljrAGUBXLdc9AZ8wjJ0rwktuuUyVGI
1BF3ldDBkYBadM/E2HyGYqkjMD35HEbCvS4QEa1v32MMxj5fXPEYtV3rIe0kEVtE
4GcK9lv40Y9ZhDj7oXkpcsp7qEVfQ04FnZXf2AhlZ/qKy+m+4lHW2ITdD3LHORUg
9rD/3fxK9qcn1syBYGM28gA435qZYAGpkgEdJh5JnRYi0iXCxJG5xd3q3/BHHDhd
Pdr1yCuZhEdT0ArnrG7kcShLRfQqHS/52PYTuOI9nYpnjHAMSxEgipoex/jGfglj
b3HdnLJsajLAnrwFQVUM3WWnH4esbcreCVBbf3IdhwgDajy54RoYlrYBL3Q0llZ2
Tu+xyp1PBcd0BKsISXpdGBu87ZuFpLuzI4t33zEgPCYMCEOHiEvpDrkjKIz4NHId
vd8PoUxRlqkAzVtlT/Jg8+uCcd/JEwbRWUPksJXVYGaNrv2/hALz7L4WcPs09xLn
uambiZ91sYd4PuLPuEk9ZKHyuYDkMYSAuPG4IhBRsejX/1ls83Im+xCWuGkscfKQ
6/3lOQwQdIrVhy3La4Bliusj1xB8kDaIXS1IWeNsGnSYFvXmSyyP1UUmpv93bYvv
tXSOcM0NealqQUMdJ8GWIkLQ6LwC2oP5rfS2fjycj0SVJ5tkO9WbmnbfJkzjFgok
7XhDY2I+l4pV2peAfXRBwDR0nR7MiWxpqHs+9yVX+BPzJCGIzlQSQYetmUBu5Xiv
bs7ICet02Dgjes3a8/Mm2cNqWDBTQLMWJeKJRWCig7jwxxY3laFF8kXNN0COzPFz
fJ9zCowoyj8i3bX8kmNJ/8gR1p4JTmWHvg0uWuvmCdvqVO/d9p/OmtEbajQgIRCQ
HOLYGwxCrd3LoXmDXyIvL2Uxynj2fTRoePz3qQquTcsnb7R53zoJld5r/6C58KbO
mPTb/xskdEuUnAeYioGTdvzD4vWxXoJOcBvhgf63uiZaN62/PsJDaTa8Dtsokeb+
ptYkENkYDu0jLF9kBRQZVsbH9V0OebV9ET4Ggd98bJP+v7xF670SS+LKHNSMRnDu
zDhmD63mklJxAE1ICkfgWI/X+4ynDcpUG148QYB6CaoqIBTqA5CsOcSUq2vfWFp4
xjIJNhrri8aRPlxRNmixmLoOpF0qXQ6dxReObxNiDFKI48lCHkGdmKQOTpddG1Ne
XMft3cvLxfeDeiVpNPFoL7a1XGhT5DaZVVciMwkXyHzCHAcjmkJMOmx4m3PGzQmT
U8Afb8KorBec3TYKl7cgZOzg5ysL9BrwLwhJwSZZYx9umDrXFtC9OsZP6VIES5qv
lyvDOsJrsT3TO5TAYzwMDSeYDz7XmKJ8d9dGGpOQ4KRCGBkEQTtkfs78kC3+HcIO
Ny8U9UwpjpSJqyoVR2W9jDhHLCYQvc3bi4sud29pHFnFT3K4jEJIWNLDeUt9ZOng
muxBIh3ueo9rKmkFgxA/ssmKRbVCUhuCGLHf2uZHqs2TRDH+xMDzqApWWsdoFw4g
pn2oFT0yQgmjqKL1IwyCe/zNJzg6WczIinzVVRXDyC/Xyh9mjeH47yw01RajAvnp
94sUkG14MvFb3xQqeODle2vf1kkg0P4TBFHIixumJFk9b9Aw68MHqp+cHy3RrpQw
t7YB3pRmYU7PBT/OxI9lYcDJmPT2ch48C6rwQjO0suOLxY1j8Z2lzxkGhc/e6qiF
ay9d+9KSiFfJpch4LsyPxyqOT9SRYbcn+Dpyopr4usCRGOdG9gdF1wKRgU/pUaG5
TMKQvKn3bQUSrLytvVWN7cHCuvbgrdDdgDDeZICYcBDaQFx/5WTNqfc0oCAX3ukM
oHjnyuyjaCEu44pYJjGGXqmlSCeKA5HOeI63Ys+mSQCzrggkPCZujuwkse0TAKE8
XVvcUk68lJP58EUURwShx4oWY5cGF6vSV8NBN9qWa1lbXuDs8vPORbm01v0hXvHp
2Os2i8sKXzUC2Vg7RRuYDfCHcqXfBu5zHsNdby0U8nAbO5w+wBNBHm1k3GySOjwz
59i7IV4tbPgaehtqmgehM14ftllRJ0yWsvaS42HPlM2edXUoEErG81ps+rPI45CZ
52X8nymBttPxM/BkKHNenL8cP5BbD3Q69T3m4WSDWWXcWbSmLe2w6eq7zqwld54d
gZ3+MwiAeXQFvqTzYpikJitsSr3rakGPZoD2LcsiNu1xgsnh0h082wxIcvAbzFTQ
sH0hcFkYTdzBxKw61HFjXt1VUcPb4bgQkH2J821S/c9bwnNL7TAeAUgkQywxocIi
qP9zf8IxIrOWKNazAajxI26MsWKNXbkOco9TYkCVHfsDVuMsmsbHpHatQTbxoquP
Tbq6xUUrREqWfBIH6A3ubfz4jLqliHKFRsjUQxAppX0R4VnGSLgDvz0p9XFYYJNz
isM+qTxk8ygorViVL+Qpw2fGJIGQtU20PdbAyOp5MRsmT1VmTlQGh4Sd0Tj/5xh9
oCMaKWEP0P8cAFSyk75u6dBwcDvTW9YY7TTvql6obiadRejd/Sg9B+TpDa2DCWjw
bRbdS8IGyGsPLBq0zH8XDX+EY2G9cIkcOIFieZMsqr2LqX/hnOwQDyKqyVf8ZXof
0p6dkf9ofq4bAsXvnT0myfFuhxNP4fwuRfGtaZrWzgmBwPL27osXtn/IZozUersS
QEywgt+W1sIR0mrsXBoOTmchZiq9xImTn22A85RL1yyIXTUy+aFdwEymV7X20cPa
+dmGvm2zBRF5U54XF+L+AqqSHV7QXUJkSv2Q8Ryr68KA9aT25BSM9n38obK4qzZ8
RwPa4DjBUw67hFbq1tXRGkVEQ7z82P6oZ5sm1zmXl8Epbj8a2wQkj5V8bUzkFlal
CPGoRNISrj6tYr1QNwH4Z0uIngLrvcIB5i773r/KS5xSsRYryOc0w56hTweSjknw
umPBwlvgbkHPpU45lsCy/BBoEzoDQus9hXcW5G4zQKVNjr2VmSkeoWLJHuqQux/5
zuD8T61CWh8BhNCR1BwVTtzjc6ogMvASI8hW5LRvM67t7YIOIQi8JJB7V2leHbWp
t8N/Nrh5fIKRoF9kz1dNtKngJ5GQK3j8u1ho6i/8t/vok6LpE8649/2a97FOle/n
plSJ9UfCAXKSY/YQvsqEjo4H5Iw38xqut+Z8NRSVr1/qlsBxyRNY06E5B8ykNhyr
vocPB+gqRdbui10p/J16pnIqyXyDqeA/NLeWhrj+1KqqvBgO19FV2hVGY0BuBR6Z
2w/hhx9QdLQ8v7m7dzUQgmDDvQFwvFBriEQVhr6DJAnc5Sat+Gpf2cu7X5yNcV5c
ByaSQ/fSpPIKWdZxV2Qf/adWXtT3gV7nmHzBLQjfDRhI7OZ22jjJFqRH5iD0XvOE
STbA52eyzRgpI2bSxD78mYhBATznp4z6e8OoXZ1qM0T9Ng5wvuuPdMo8peYfIgHp
XGYTf6Vg96mz0GtAQC82v2/fSj48fvyzaAVhV2eBgwGwU/oYlZfQXzTSKMNCvkLP
BJWpcWtqfwEP9J81e6RldwkZop7K449YRtWSv2UJkuJOZZrtZeo7flUzr1bEehH+
5iZSQgbJdwBSpeeueeBHGciec+Hd3G6AyAFbCxynKgoUnYbD/6TqF6jcmT2X9Dzm
nQOcj0pE0akcjLJOOH789A9TEMhA13tDDoDcpAfQkmCxA/psTgofGl2DUWsxJjz1
lLO0mW2yT1O2K2suB/QgwuK7RSoAwW2mp2nbfIMmuEDspNrOJY50dgwSwbWT7a0L
xYbeX+ZWICuxBRwAF/G9+HzJoWmXgJK4dWXqIB+vAl9ow5pi/QGuCa06e3yPTHtv
YjNnSAsRSmvth1tiJxuI4F3oaY/R+/qIN+lcbyFzf6WZqAs0cIwFNlPKFfGqrwJ+
0rfGhi4aMeX6mgUXsqe9OGbLkW961Y5cs4azgf21kXHAXjkvVNsuW4p/8Xg8yP8D
s9uBKBwnjCjuMi1SA57wP0sz4qUnsiQB52g0e/5z526bLPOw6ArodnQ+U2e8UGG0
4WWyXemaciticY04bc2ULGQo4vsFdZLEssRYa2vaGk4ZPyma1gGYFzfndsTsK3kp
BpYxA3qWUpwenQLBsHbgmDCuuIBBV4ZziJOt224alPIVP37ZLnt/N4b0Br9/CM/e
KxQgUPk1daoCA5wij6gUsTeG9ZOsF9BJev23V3p5sp2WyCmmS9kXpmuUD8CCbM2o
ft5W+hNoDEztfxLbqKjO8um87Ls1kH4Sg/6dharb6ZUal9TbcnyludAMQ3v16m1m
vulh8xhvzyk27B2Kifb0KpPLdYoqjzxZeXwYiA99p1zrSvS2xxB5LnDX8TjS5JDZ
BUGrCv++sdnTiBfo8lZTv6PN8Vn21dTy7cbmFXLfcHidSV68673Oz29s58G+yTfV
k8Iihyuwnzvh6Lp7/BxFQMU39VA3RYfQ0vb5JsT4vF5M+/ZHuTi0lRE29aV/Z9nD
QbDbnDgcCBy/Q+gZeMTH3kzMzvFboKb/238nB0gwqHnDJ8lruRmWyIfl/7zFfk7Z
JcUl2+DWJAUyzF1gLT1CHAs/VxyOSWWKK5mYmq8UrhodRcSpDp2gIE8CoZ3C3L1H
w+fo7paE8krJ3tZaueW4ITdsTw5v1jxmZD8s/FYMSKqBF39wdeHkIVLr4WBKCjij
nzSRFVv60qBvrC1q0JhY7AyI7NsxvU1f5MDbnkgGy0bfZ7/Xf9dz15zhWGEgwtXy
ybCzR6XEHIYefiT9DTw3d16WImBrgGl+ChNVbZq8qi5gP9Lh97VeAtExxJpfRtMb
Hg4nloRGbDIyqTVz4BWwnyAF047b6OH5i74lmvLhI9QOv9jy52FkoQWnTY8mdplG
y4u4Hz+IcsC5NTgNQOS2JRQ8VxufbGmo32wdnPmeeDBghB46n6G3uHSmvz9WbVd4
WKUEH3waxN/u74y91lZagNoA1WXBqNoxuEDu91+Ie7YjkZjbMNpk4U487yPSwNi8
VaXFWzmD3watczzOMYHA6jHHSs/AVzLHMmUFbFwXQI/fOlTXAlwCj4oupr+RaKmP
ssiCDBYzcoGbTpVPNKOeF0zKCWr4PZL7UHzEwQ/3zHhoNYNAVADH89ZZemvhB2Ik
/5l2C3zbj9hy/Vgj6aDFbaz1rki8AirJCywkWtqaHlyDOddPBuSrbeIrOPMvRQgo
yjzDyRLQj4GMkL35svONUGJl7dKXBAHCa1jiPZFKhN5ASiBVe3lwGaRQgDnJ+Rr/
SjvqrZU1LdopJILTa5gvHPBxTR818F0oD4b6y6qQGz+MeYsQ1HVFKSQzRILQnuJk
aWfkTvLZIJ9wramngDy0U7kUo+bVsNFT4U7A+1FjsdqwdqvmgwJO/z6W0srEeOIs
ZOS/vUam05IRX7SQ5yLfXLRRgZ10hksz3z5VRtBAJNEn7saJoZruDTSca1Tq0Gww
DjcGEhFOruwfJhlp9CGfA//uT989h2wDUS9PmIk5OadyfulVzvk+XNpifWvpUTSq
D9ZChSX28cZeb0v6WKF6KhO2PTqSVXEwbVNKNTgmoyEnr0YBjT/5NMhEzI25H4Jt
xGtRluySKf2dk/Y8VEUoc6OUnB2+oW4odJJCdhADcbtg8is9e+GLjoVOvAk4Y2S3
VJOVqYBZXncW77IyVoXY5E9GG2lTg52WPMcdEt2Aqls6U9Z8XfH5K7OXH8w77ySa
9tpPU2MDuiFr8/jYtvlwzi1KFyraQrsbF7hYwsSmhZRnyH79sihGM3cekwroUfdX
4u2lepBVz3BxhRPZSFH4EAUnw8ejgbm4EOL28WeawyLIJQs2eNiT6DodzxM+VdPC
/QgFhRDNm89owanBD7+X7kaZAriutuwPcTU4fztA6xxF8uwT5vIWQq0h0RaiIB0A
sPuepLd4GG6IZrcwhfgu/H+fT32CW8VxyqpD6u1vmzZBDnYHezwesfxZf5w8GO7K
lUyNO9MUS+Mo5nK23BJwKcfKz8WsPWIQKxqsMwAmaM/Fxv8Q/my6fWAsUasVc+gq
h6ahvNynkgG6OAw0IjfzJKVmqnMIESBDt0Gu9a7zuQWQQht8c0TbzHFjSnYewpJT
h5MLyBQ45lW9qVEz1KQBeWSvaAuQlIW2UGzh1D8IExzl2Z/Zmv/eE+tj/OyP0mTq
8ZMF9KekGr9ivOOtweunRNfyxAqLVT+d2ncl0Vcylq34QxREgB2//Zk2625MU2nI
VrNXHvmehWwZiEEeN92Qt8JqkuelCnEmF/2Mhy/hUvMkoexoZi0/V9lSxVmzjy3U
cgGCDFW5BP+WxI/8XNTKcoS07Tr/Gyok6julzl4vfbwkIl5UFZio6dJzwSAAZY+f
DrGuPJvlvmCyol+hpw3yG1EZh9uZe1zIt+oD3OP51GOhqqDbSUouoaodS6GrBNdd
B4RaDOudcYnlWuh75stXg1LAiCu44tNlXbT8l6uI+SX4Qx5Ckn3vwAQmZGBRVlKc
s4K1+vxNKkIUevcep/fPZ1TNpLqqyfDfdH9hcytzv0jJEcILGWwqmlGByhc+KBJ2
dvPARY8PTKFXm8XqsbUnPc6nZ6kqOgdb82nlrLNh8iauwFMtgUvJ9Pv36yzNNUo1
y66HTSFpCZcjCmZtOXxJ2h4c5g6z+BhJTC9q8J31wKVCyBuUBLifje1xaqUeRCis
8/HNW5mnCpMXSrbYtazgYc+2OftLCBe+W9uMTV+cJ+542w3hpFO+3ABQ9jxpi6Ey
Q+/KaEXMhEF803xfWBM52loV+F5crM1wEjR/LXssm2tm3GUiR50+aaRAt6NTDE70
974kmg+tkygWXlD53DvDo1JmdfXSFFXTE9tEkGpt91cj08X4Su2DGRmgpYN+lBVa
GRjmfjR4+NGLUa/CInRjbAWgqLx8XW3B6jOHwp1GDeAsXCr1gesnVYiTh/4WZEKu
PC1SQr+0aPJ0yaWDGJkvWYRwC1VXbLpA5L8v79bz/mffmvY25SaiHsk31hpLmxMj
CnOvSQqDWyn2bvuH1c79Ye9oXguxjA09OfsmmMQZZF9GxDyyxL9luGwszeZcfY4G
Yd/xKOyMPeVm2V/FpfZLRtH1bVa+Q+onRCSnqDwnu17jf9K8Q/0e3jtSkIhIvFqZ
AIOme9M9wcfRTqmJx7OXPBSTkT7hk9+xNXR01qghkUFFuA2jLAgx8Gc8q4a307Pb
q6+FYMTKhVLPdfBydLYULIrcNdo9ciaDdylFjm7xkRsz1GrlkTYjeqLL8T/iEgMK
PejM4zJvVXqRYffcPOSGL3rBPT1R7qazKwsCLv2fU+3Hbt7ADLLyvW3lL7R8ZZk4
RZOznvnDa5NeExe9mHX37E2gXXpsUqmGIId6PrEIPh9L5EjiLJi79x9PA8kkCwG4
LzgJvfhc0xtdBqUujGUxaXHnHJZrl6OV6uHAtN1yvKXbfx/P4DIMzKdrHRKMJEBb
jch7AnMjlFi14awKO9MuqeGTsSqOAa96DM8Nuup8iJraocawn2PDmAIVOUKje9wl
ZKOWJKXQhynLkfnB3k8EjklX8ddny7IHQ0aBtgIVQkjMSKXSuF2aStrokRlIjMqy
ifJj+CMZ/dhWJdAQbfAr1WahdTO788ZgYcQ2LtMbnbWs2O1zT2uZB+F3hRjp9L1d
0tpTG641sMBt9kLrSrok1XNi7vVr1Kp52mhXg0a0jmglhG9QIiPUDj4TSwRpwpq4
j7ywYJboAXQK5cvR+szH7ioWDOLz7ohnJ2ENEp9uGUaSa3XVvADdar4AcIAW0Pnc
iwdgyozbYCSLxupZ4/d7ejjxZUvWWNyiwqsNb0r2HtKzwO1cUPEVfVDKA0nLgG2N
nioZlh0+h2piYJZLPbPqZDd8yYGD/Wop1bS4ARzuQlgDipe2t/FNjQEL6acnxLGF
n/uE/AtnwHiccfKqubBfj3o6nuEoqKB8Ik9ozUcSdOMe+We/rwSbidJ+/FWCqgX8
DsEABMvI33/0KutRB9re686PpamEa6fnxE9tf/wHf+uJQd475XfHRlfYwBFK6sHt
TIEfS+hpVmBV4RV7Wf9xFzg6DA7HwB7WYkH9Hc/zAaPbgQfhS5S3g3OosQdLYt8l
EXKKHYszKMLJ/B+LvqKe8+1UOROaq38pl1ynP7q8V2duiV5sQmFMcNr6fNPYH57d
xlVGpqjmmbxXvOCuxJqfHz8EuBwR0v2ukn8PrTLm/t458GXjscVegm6hdjG1i5M0
Ug3wM7H3BwPZeB8RlL3E72ZfaAZYpSL2iAN4w16KGFVXF0LAOPRSsAHvarHE/Exx
WcpDZh8EzZkve0hh1xmq/W4khvKyXoMPl6NHGxutGZDAAUl+FE20HeRTH8b7cqKG
XjQ0aLQWqY1skbAzv2EVF7IFu0DQCRS4kaVAqZcG6LmJkL83rRaqnc+0tCpmTneX
ovp7lefFMFtgqJKdWdnTAA07Zh9G5IdFvC+xi9WbNa4z5DNBsmcppaAgyHF3nSR6
wBGny2ZkXb2xOGuzptC/wBwfZFuG55H2D61iKyrT5LyovYng7yPFlMxlrylmQMn7
keM10XzhJSNeYS6nZLER1nrn96id4GM1qnuQWLmpGKt8DSFqhL1DdMKHerVBWmsP
gvmOx0R4SCiqaofRvSgF6/KYx2aTtB+Za2ljHjC0ok+unF6ulRkjLNwRSNug+3Xn
rkbt4V/Va/wH0VCL4OaAevt7JKJHUMJyj2NgquCiEJgM7PFHchMvH41nDSql8W/9
pSnZjLRUMFLDs3QpxhyKLIlrVzf+V+4NA0KgjnSzbjwSczlWun3rWN5dJIw0vF7W
dIPKyaI0wCh16wpMguv2i61iQQhp/JXfCF2E+sZdPjxRxmK6/CMGg8J0ihO2lekD
czz7ySp64OGjKChJe8nFVpcxxbwG+dg+N1mCjsHhyY3z9Sv64JjTGHB/XdahbQ2i
Ai+hCEpRhCiiEegdSrDhHAjr1Ev2gJPoDyMG3ZbYtIRKTq9aWng5AWD2hxCQh2U6
+YcecoD80DpVZB1A4YAGsoEKFrcD2fDKbl15/ltS1oYiZYFDfy1j6Wk0UKLZ0O1T
VEUPzED6QbV9NOb0iXByr1s6m3GpWnpNstpVsbF/8Lb89r5Tm0Kaf4uCWg898dGc
r89do1VHHfIXv7gz4lpZdkqzgvrfS2FlzFRHVU8lx5AhIKUE6oJJbHlZ5ta8uCS2
OqQgIoBbb0fxzV495ZlhFucBILsaAp+bbxryQcC++XM9u/xVw7xkIWKNtQ60TgBb
59wxvFI80hMCYxrnUTsIt7/gfAtHBNrvbSdpUtBmPlIBeRRKmAi9pkZo9ic/eQQU
5rd86s07Wlrxtl0NnZhjJD9iziSzJScsy426p2vBjHY/xbbR5h1KevPCvOA5BtVf
X0bNsfssQxDvuZ+AzEKBtt5BRfDoLF6/TYZXaOuDN1iyJmwaPdzeIAPxeWZLrdZ8
9pm76/TGhGotHCIZ/6YC95R302apnvEakqUppRA8zQpIyqgMsGKEk+wrLp0SnzOq
+p4O4xhbsGLWCM4UvwKToTZ6D5BV+8uHoWGmsYh4GEaSIc6GZU7EwTVK9WoLV01s
hFJzm3f3XxKjBibTRGfjEdqZDTxGn3Fxvq5war4R6lDhahGA8n6GBgtOH3hIsLHX
yr3JZg9gmNLLQwXh6j3l5J2WUgq2YKr4uD9knjNhiW4vcTy2STiZfG5Tsopaidxw
WdEAKOvppGqknvDUJpQV/+7ShuYuI2eZc6LcIklIDg8AaiHwvWedgcqDO190mI6o
jNfDxFlKsKOYUMqmMJaOWRfmHF6/YWA2oMzK+oiYWEOj9SVDW6skNcECzsn2wscX
p5+54mS92mHTgB08GzPa/3+iI0r4nTTP3IyU12OqPLbFWn44qCGxeRzL+PeTdRIw
ZQ2O4aHARc0PoiLjs4b8OQoRlOwwB1ZCaw+Og7FyB9Y0imdQeVqDQtnVcxWOeo2C
5wZ1TzgZCUcQJEk/qh+0cie+9EqdBxXA7swRjKUf7ehBCy80Njb5IuK55THStr0y
3uZsHfZ/hVfjkuw2mpeg2jHDE7RSELftREN+POyshyE09EiBmDEnbojNkjTO65Re
AI7yGWagoVu+AikT5QTqVY7T1S6/Q8Q5QbXSLuv/qEKEu8ML4nSlj7nhf72dcsDJ
l6wX5oQLrL8EOPxqAz7c1WM+tGXdnoc6yr/hHdXGJJRs3KkJhsUpv8T9kvE8KRw0
/en3gw+kUBn0xiIKcn3iqMmlyuTMdyAsH51sM4vKRDbQYudP0hFpTCL2zvcllVSa
JzmbXnDsQ8ly7xxxn7Hc+Rq6GFf6KtC35z0LbxCrmnvUI8P+QJO7auYy3RXBjZoc
VeuYBuIS6smTwt9A+YMrFCkxVdrCUI23HOGuyleiO7QCb+5FwTBwxG92ZtjA6flb
KmxZaIDXPGemxj0IqrOvfW0KFOcpWJHi38HRYtAL+tC2YaweLjt4uOhLFPwhbb5x
DoUvILP/91lVRjzxtyStL8ldnnlR41zbjQnIAsXoG20OwSCN8PcnGOq/nR/PeKvV
WDfeVwwd1Mi8QaddT1zCCRHGJtk/WHiF1YvWzt3QgimdijaohRmWQMSobLG1R30M
vmkUwcuooklyNFSEdeQcbRAPGNCd8uatZgdJ6MvaiDq1sftU+OVgL2ai/HvHq4fu
Qck7gmC0eS/LPjcksZyynkcDVfaRznrY2PAOzDX0G7cSwYz9j7mmiz8NXterCeDr
0aNuejfZcPcGrHoe3MlbLJlwprCRTzmHb/Jp3cIv3ib1C/nWWjZd+VurqzK2d1/f
N3Q7tTlR3C5Q8sdB4yn3eT9uDlifLyDZtcJ5aNBp7NWAfEkBtk+aAwQjBU+E+ozu
6+/VZvaRmOHzpGGMrMbiJy8IqiP9CZoGS5CVtPKbDF5/QxLNv+ShXG3N9ITpBtlQ
pzz779CopOrHqHNSNTJQkIodOlEcmQlGDH/5Svl9qhOE8PCLtCu//vn/e8oI1yYU
LwEe4bHSOFQn8N0D/t9gSumr+Qkp4CGR579tyzuSHv33qOCwNiql19+TxESN1Ply
anHpJNO7UW4SVdA/FJlCgLPsQZ57oc89r6mBqc7d4I7WEIelpomRspD1h2/ugjKM
6qjsiBTth1vtMAkGFmUD4cdxezIKvcCfQFAggy5N+sni0Zq2EKVPG858dq3nKsEj
BBmRyIAY1L86NCe7YAS4em1i7CcISBw0VeAg1Z4VPfRX504a8ow0Q3hE04m8H3cr
WGOqDB7+gbUsrph4n/ASRaSMRppl+bnjCOv9RDu22FX1nQ8u1+J91AbSu2/inFDU
7Dl8CWOiFxzBLVHLxF9erUY26qTNo9IIAX6zPM5BRd5jVP2ekOsotb+8zMBYSMoY
g6Z6GYS/xe0CFSjg1/RDwbeIVUlvhvudMdVe/XT8mYaFzdxqoCU+3RPeuriPJ8Zx
n2Y9UyPNv2BcJJA9i07dP0CSxw2gUB2lsG/dQ3lpLlaFF2yKqXTpPitbPrefB5KE
A2jc4acy2j4Sa1+0EdBrgw9xKqVvG1j4X6NW3QyiIijqn/V07PhLhv6temySo+bh
ZFNwCWj63z//rq3vzCJy/zm3h84JxrKrtJA0WlUaBebQ650UYUtG9PVXlTC7Dyeq
+mps13OZ9RcQC2+ITOmm334/52+RdNYk0TNvpXF6QlHYjSliI4et1qrcg+EjikLo
E18nFnIkWV+xPQwLH612LumhdtS76uMe7Xx/l+SDtIxDCLapsBijcWHK0nsUjUIj
UkuCCcI9NnCUhKCniVNpPGWXp2JWCDSiyHsWmlOqUsu0+QpzLxj9MU1YyQMdd8qv
y9DfMQnNVxeWLu+dWufkt3TjEWxA8osIlXz/jeMeALlbdRuRVdqAs6Omr4SCiupH
hQsZjm6RZC27fGxhoWD5hBYJdfUlSu7OSPW3/Vp/OcMYLstxeOJr2sjw9eWijj5Y
jfUztshYljWSydSPPdTSjtDgPIUWnFZ3bnAsVNHjCWMBhDVCNt4P05ZYgKH4mJMR
orHifXi6IhQwCfaO5iWmmAHwubrhPBuGQgwBCjxaopBoK2sXZQDyYEokexWmZpNZ
Eok0NBQPzOEQMukhZYr5km95V3OajIfT936ddsm4mhG7mBcjKyp5jqQP5EtgCw5K
ue5lmrFxHzWqsibCqngwHwUAKHCxn4LBiXc5tQG22SVDoE1tUWcX1IdKOojWUTC2
Y8bLj7khXaYn4dDaCwWOjsm46pAfZ/pmFSNtnCnIYCyYSpyDlDRnd7DP8yQ4EMqL
kU9hp/XufnkMjOtJ8EbX0GIXzg7PbK/7MH5Ldewg5Wg+C9bXeouSZ2qOHfuha0lV
NctaDqp7Tq2YWzKQox6IbkDDUAwPyUORv5oGnNGLuf0Wniizd3126a9+TEdKI4oi
dUtrMFDQccynaOyKPrnh4RgLeOngMToJoXXuEhCb6FQgxhLef45VW5OgSTYE4w04
bXuuC2k0IYjZFp+FSOr+zVO3RwP0zVmwbEgasySc7cpKXmJjUHGmSLA+69FrGfJE
7rkUa0mb5uHgetnBDoNuiKZRGsz0ZRemNAM8epQSsVLylOrdFCGDZloBQl95gkAb
wNe4q47Bk+qR62KclkFJOUd7kPAEiDV3FbPPWlP7bIs2WOGIBRAhnjlGbRx8fZzR
+jqSFlvCiNaMh7qsH5TawH0Nt1QCsmjzGZuCMiW9I8Drr0JymLFG1qFi/fdgRlBx
JVT5JrWQwXKOiCQHrbSx5s8wl5Cq4WciVoxNU7+veVnH1xdcu0TSfVpdTLDiSKYs
Ib35O3qJ+RHRTDNWpMTGmvWdqhqAO5aXyEke9t1Sy08gjHPOynpgrARGucAXUGR/
UmhzvlLzlhyroVbQ/XZa3C4JqL9M0HlX7c0oqc+DMyzaV+Eb+ai56ag46YOVBQlf
iQUc0SowdErEmlOC/TE0WeGyqbsnBs/L/Bunt3Fbt9dQb3KMDsggFdNYOY/nygEx
gXQin93LpvvAoJqrNlv0CihxEysMS97tle+fO26evcT3mjVi3Eclx5MF+BfDcXZG
ZBh1EJXl2aVacMNWKWoYq3WUgnsZQ6HuvNT6Ipg0DYROvtWSm8cYjdRaxF/KuC56
qTyqTS7TJnD2oBQ6KxmkEETUJVF0vOmGqXTcnrQzDCCyLH1WzvCV3pmYADwf/GhK
+uYgmM9OqY3FUGskxCZiDIbDXkJeAi61lOgQLO+jODjGE9OF7Uc8D5kqk4fKyb/D
ODEFGM+z5YpTX74hNN3gLpKFxZ4wif0L0/fBgKUTpOiTYLeEQNmOhWXYYgGhm2rx
5/eYLIl6CgyHlidBAwQuxUqoidH8E2T6MwCKdgSgXdCytBUtVb05OFdSyLJxp4Av
HLprybgvXjvk2dappQiwWsnT6yAcq50CXe6OJSTa2Mr1WctF+4Z6cuOIGLyDOKlf
uHtq9G511GaN+pyc/svwEHA8OBbBYspknXtkvWtjzfBU/kWie6SarqHw970KB9Q0
Zc9miXT8KbppIY883HzJYX8J/XUfdoYjOpaUnokagn07QKJsyEjRUJgC4XSYPLnS
eIJB9ZAL/voDtnzX9X+IbY5DdHzonq1w95ryOKzgDyC3CIBsQ3tddNmut6LbeO02
+9kfqz8fP5ef6B0IwhsBRH5uHjTSk9nbZc71sOIBl4bNqDA5TtMH2xYBR9dOwakP
RrHFYwM1+WJE4x7M31BxyqVkOYlNd2deYTMXdfm0eOKppWP2wLAdC9fF2K8c49h4
Su+1cx8Kzw/cCbAJPGP2Bk54lgmBZDW1qHf7BEBq6PZSfbIUOSN6mWWqExpwZRaU
ZD/iUCSn0PfjWMrI1BxnhnIqcn/b2fnVAYsm13S45xy+8c7VMf8aLQ6je2c2G2N3
I4MWzJPNuXXlQy/+QXfyp9HHBbpCVklFhC3S/zNuVXptewUF0iB3hqZoX6MPlmd7
IS8mK08EXrNRKKgP+i2MNtGw5b+M6NfgdD8FAJJ6UUvzU76v+kUDBMJX4jBtCrfH
XqiRfm4In4/djJHNY+IgbIrCKqL7Bxv0f7LgrOTtX01BxjXW/BD2RPnDNw2x+BH5
B9ykq4H1RmDeFYpmAJzCSVwZYmrCYsGR2dReS2JF9yBnP0DUH0o76KztJp71cu9E
ol2CEhzh+BykZTiCN0ITDMNLPTJbFRnGVLNRBlD0Vk9EyDMLa1hgaQJ9HMvHyiVm
MdYDG6YjSzk3uzVBpdGl9DOEJnCZ0uEuLxJJxQ3I+SZP7N40AFUa7i0GpTlQRjZo
ezKU86wA7OXpIzU2EFNA+iHX0vEL1ZcaHM5/f/ihbjPZvnJGgAriKxTEoF6UNXZn
Guhom2+QvDE4luVmH/vbtZUP3q44UfiWCN3Z9b+Eg2mKm9HaQPkjZS8WIyCKxEoi
hIP2Tfp30dYLuJ11cyXhxXyfN6vmzHSDfINkKonJA020yjwUGuHVmlHuiHyMcAgg
7rW/5hOnTywwW7L4U81aWIQcZMwR+GMtajteyvgZ4+dxthH/fNZiHrfj8e+5bMeu
tFbs4lLkS8+AU1dP/QIUfiFScP8HwfjmVb6h9xWnyU5L0UXV9wTOsa8OmEpSp7i7
Xr5QLIdzETI26DZ69lOzVlAXLLGtjsklrPVCl3uwTxer9FFdD11oIQGFVLPaIWZ1
hsJ2UAnGfjvWlCnvNfM5Bi3R9IKHNZ1sb5XRYa3KM82+D7CJfhnPeY6oxgv/1mmy
lhVYJtrMf8F+iKmvGfBXuWE6xJTWMZpso/nv9rMamH9aqNhbGvrqbn1htwm4Cbt/
fi9HD6m9dvHEXaj9G4C7ltQnunWY1henBaFQyOLmT2e9vSDYWF0qI33pmQ12GO9d
hDV5dhUTXnNM8yi54EiApitpF2ek071uFtwmThMIq7jOk9TkCP8lO0tJ+Nai+dZn
4wBB9EuTvnmdLDBv670DXUv2XRl3zlK2HYKPzVkKnj2c8dnxIHxdkAFtVBfk+DJw
+4bU6vcoid+C/HQdPwDzoP3c7PVsh8/d0Dr8MFz8/3H79H0eXFrtE5J9+zbE/7mX
3LRZlMYkiLRqzTfVvmgBpg3X2Hh6BuwKQBxewKzebjj9RkFFF1DDqc7bWjeuoNxW
Qw4ELy6XTIas4Jw2kBYaWltZl6+GlygfrfasMh2o1BA12VGc2KT/iNdkTK2jS4KI
87PkNuDh48qeifil9XSN9JG0lsb33ZotSls3FgA5DZbFmS3h1uv7+wL+MkjHDnUy
R+9CguL4w04XXmTxNH76G6A7ORtROi3K5apVjTkuBSQRcjM5NPh1nCNlU/rp2PEw
KgZutgzLe/d7pVHPmCVwKR7DlHqb1vrMXbJX8VWwwBHE5kWUT5Nl3/68JO8vAg/i
Ag8f1HPq9LggaUxmx2Ath4rrFg3hIfbKbPKns0y1PlhX9iFEHPKc624ijQnWKNjf
j/j9S1zS9utLRDMyLKXbgtk9BMQsZ1NjJ7p1Vcf0XL2IpV2QVQbH2MRy184y0bdo
1bFg7+tVbjAE5D6YYsbAoDt5RNHgA6COAikTgAhtVf87jF+zAK4oCnYDXyyHcasT
p70aggUWY0RLulZolRh2Cu9iwpliXBHNxgr2lOiPTpmwoAAqqQCSMRnlTAzCSkgu
b9f8qi29UhhF6srYzeoOWpDR84qB0HEIsnDp+1Z/ns5Pda/1gePBm/Kd+3bZUEW2
Jd3z6bdBwYAKUKPI2nRXJQXaM/bHUGhCKU60epNoH9XdjiU6wFH57ZGPI9joYq1o
/wqXjb831DeNpNh7p0jhwu8fnRxxqZYLkKkqxrv77e9ELd+3h0FBunf0XaBb0UEs
A1MEecxOjJEEwfy47fctrZRBDuzkFJ0CDGlHSnOarMy2d3LlBPDNjtheBAq7NJBH
JLFi8wJwro9/qscficAsdaKYTbOaOD5p+9nnsg63tO2rPY/Y/PuX5JIEMt1MVLwV
RXzV20bkf1auloxoMx2sECmswkz7hZoG+ZHca25wDAt37G1VFzzN5hXLFNLGuNt/
hpp2tjFAEzFXpxetLgd908DWS4XC+2sn0+ygQoV8MVJ+uKq18YdP7RHI36De7kPo
kLZbUO6oiH//bh6zLFTQJw25HtGb7wcPBprTcxIsEIphImX7g9FjKrZtRBBcKDUJ
PfvguB7+YcVbvy/6jj0uXKP+VdK3MbkiKt91wmUaFmlAqjvgIbcIjbae2kZr8O4P
Hw0EVSHo8T6at/WK/L/mGUuVH+W3hW0Iw7CgxSkpMbf6sUxu8wJGcdPxF5x4PIiK
WLqcu0vJ64NeGOXwNKf0+M9nm6AxSQdLKM/V7g6Ayq8nh95h7s+kTAiqZCIl3Egl
sh4EvAJu5D8ui/xmZe9+IpTIX9cpWOQTPqHtfYx64AARrtI04KRdRjjoak4pHWWM
174TPx0RafFD8q8djwQ6GOXqAnqI5YrEzHyf2OH71SRRE9Kf49JQ+KkuhgKHNMNI
o9TTioD3QlAKn71GRjhed5Sf1ule4fC7yaFu9Tr1vQ+DZpOTHJUAEoI6mIpFDpVE
hgFr02ZiuEeir73gFbiR5gK/0sjeaTsuC0lrTjIq7JeMxrcSzqHo7VBLcgsDn9Ap
xhVe71hkybrh+nZ7PNCf/RU87NV9ugjW020BrtzPkuThBrn+EAdgkV8min33Utx1
7jzYflm6M7GB09tuYjOoqID2V+KUpU1Mj8UBd6J42OiQvncc7nzRAnn0zNtiAjH3
5EXpxRgUEK71OLsA37+rZl38fwl+cKlfTc1PWg75mo7r5afZg685csC+IR7leZGM
U1XnpV/4xU4eBWU8yPGyixOsPtHzIcNVZTUNrvED17ROkQIU4LdNMlI4smIlwk2h
2KNKeZTGru2aPJnA/13TsCDyTyb7zQ7pgMUl1cvEWugnpn7Tvca0Edhks/QOEX7c
iHgMl32icL4AEraqOLXRpzDpfxwxhKx8PXA8L5VW7H2YqhOYTOhyEyd/Ris9CZu5
0Yi4RMdpUDGWgZt/THx0VToKKEl1wxkzsrbcZN1SXAndlnuQPOW2XXk4BBqlpxx+
lwOAjUqD/bSEA55fcTmyEV5M5sl8RWAkWLiU4QyxSy+S4ApzdF28DmojrFx/4AV8
qlcFi+QzFS4hNG9AX8WADeCoj7cyUhWofyi44dac/SXrSJmv2rps5sADTqu+42Ss
9hFN43diNDfNo/Ipc+urqC+YaAJ5DGfp/q19IMjCQHz/ScjstEP5mnDgYFJQy1ex
+BUWNu2Lb5Wsn1gp/hEPN0he5Qkqhk64anaoXGMoP/yItSxkf95DZWYMAUXbgZ95
TtkprRafmL8aQ3pgi70JcomFtZWzoYGY8IJ01XoQO40D3w/nDU6Pw4Jq614uNf4I
VJrinmL0wptoPAPvWTLwKa7AepUeSbD0JDB1oEyvIOXNWDXJbOu97grzH1Vkq09t
bgyc5661dMCtz5zdvHqI6gedKkaWP+rocsP0iTkt7Ee91hVdm03v2/wF9r6VOWj6
VdmEQCgI62La8oeNc3sEmwLhroQ/gCr5Y04eHsmGRHPaYHIeiRmFB067Dbqk7n7n
869FYF38Ef/6MfmfQCKdQyzAT9pkHn687d1RiXezPJkoK3TvWVozdYDcjBlF/7wp
jTUo+D1YDMLYZn2rz0TOF0oY9s+gSu+pfhzBnOKRBPUezmT0zpMDT2OZT02HBRdL
DoZ5cuPU1x9sdt10KmCg8PjTk/AMAMnvTP+LAf82y6CX9/AIermYiKsx51ud222V
1Br5AZtqfxn527SNlzPBlm3QZAiZsEkeRlZ5fbqzgvgNoCQg9q4KJx/WZA7ykgcy
1C6YmYv10tJJ+VYOM2c8ir5nvL7B98Xjp7Fk07xaV7/75ot6rQsvNDHAT+mi+IH5
iI1zKmPAQwIYZJrU2alenRcKaud4KtFJ97CIouUamiMqCt3qQExYMiGmD1fl0UnW
+3NIKkKcKEvSdQtPszIZXcaaQIqXSWxSNwB/PNhe7joxiALssRDWaCOldR6KhaHS
ar3202Zy3Uf9i3q1zfx4WhC5dMe0XCnOgDJkVHC7u2KrFC0fEtMExNTxuS3+WS1z
JfKf2hW1oGcYtYS6og1X9j87jn8v6PzkZ23IJteYw+WqqkwMs0Q4lj4V79XeNmQI
a89xPaBF5X9/xAXSbiNdEP1wQLf8Tf42OeB+hsLR/aLSNAAM4tMM7RqqNimxzI1h
RNlabw722CNoWbTOEzmi4GG8BqWVetomKJsyMwjKPFmnim3WS8exiHQCof1x6ad4
p5cjQUNVVnkYJv92eEbfsD0TkiXcq6Zh32NnSY6i5lTOaH9gpxKWUKe7u5DqNQXt
Z2qU6e5zOtDPk+Hnmt/ARD06mJWML+caqp7m16Ri+OAH4IgkwbjT6uu83rwPVIeE
8cg8k9Bjt8QHnKtlmKzS3lSLfQ8FEPMpH4awJw0TdIW5F5F7GZ5k0Oul6PhkNgA2
Pv7ybV8okMKXwiL+WuYeMiBNZdq8SdcgUsRMPMNVzmLCJChTTnEqpYP/TopGNoOF
Kz6JDJRTX1us6usz/qsIh3UxvBHFDe/XquoK0C+3dxA0qCJtGEZRLQVSEdVAK7az
Yln1kMYRIQ+fIvAwT9VG1B9knvNocmhAz+uA+NLjD79IUIwvqaUJqN4lTnBiNCAf
9ZrebqjfeBoBYLp5yqBmVcSBxIwwyCM/s3GSuA921wo6VnXoE9VJ6yUri19xgBql
44afO5qyuK0nLD7Per2NXTSRgMMkGAdaQ8200ii9TT/ywFiDIGfA5Usr+qA1wz8Z
DhkQPcY7TBZrT+Av2qEi3ImLkEdNxAgjJaGcW48wUERb8w2rdOOaMsjvwnJWLrWl
8MeGGTk+Fb4u/++Fjmdc1rvH+ixmyvwBkvd4ONjXbuFxj1Pb8s1K+zwFjtbphPOu
eC55+AJFl8VWK1YZa2denhyw5ZfpVzFkUUtRK5RQiByAQbs3ZsplUEQOBkkvIldc
rP5k6JyfUfVXXJ/GZi2Jt9Yg0M9XNvy34OFHbDFbchurRcywdyzRyqz7l2vdZm/H
7DmZphZXUd74IXt0SfW75LcJnyBNqkPVhXg214owX+hosnUrgcxdFrvBtL51aQp+
a4I3Cqv8XqHxksBq3HKlV1kQ6Li3Yh/tBIzMYu5Nmyyu6iVG9QxKm3rZmnJx+rpy
iU0KTbUnyj/TxLlzY4BLclFHcvYeCpb8mouFhgIq/cf9H+/NW22Ua+RkWB9pLS1E
B3MZiq//ww72lwCnrPkT8342TTCQqu2ElLwQ50zCUX90vcBQmqY/voZ++9dSjSgx
qN2m4iXrjedR6zSam9+IMzO8nxVhvEsahmB5aKxAa2TlIiPnLymIOltbhDufb9j+
77LCMpPqe7BwGQ6FgP3ko8ucAxqTOupEMqZ/TX+6y0Vs/2Ark0a9UV+FqqM1bkhK
xl1cJxQ6O1mq5iV+uRbStNGb89kfXDTrHUQ3FEwTiQjGhRcZiop3YGRJ268lnkOs
KrBvctYkavZUaljxh6mtDfg3aIl7db+9HBEEiVsiPiObjNaSO89/0U9UiieeaA+6
nlxzGr8Qb5uNeUU2mmddvFGDSFBHvB7oYnpxDbBjywG49MoCzdkWjJPbjHY+fjHj
p2oVBiBtZwcJtnFL8m4eJO0NAiLOAZLdHPRymGIwAD/s0DDCbM0EY9ETB6s9qKtI
DmJxSp9gGyVVRy4AxicGTAe3BytSoKKUri7t9wmZSMOyZzPGq+PZSgAk8cTdYH34
w2I7vajXY1MmvjXHlep+3AUe787sxqyLGWP1j3mbWNLTWNU2STzoVuGvKNtkG8wV
O4S7Q+1dZgkAqWZ/c9ua8JzJnXG4a+1dHJsXGPW1PlloOUhw3PqGndV0yjjFdpFV
YM9FwmCL99yRkYZwinchtGMujfjuj/0xzi47VKSlAgO2gSvIVjnQNH+maI9Ne+MD
kESntOndNgWjlOj3Wx2xTYO9uAV1gaVwomGXX1RP0S1Z6EJC9JtzaJfoDWwYgTdD
bsKoHH8s51e7psvsAFwScncakPk56ibyB7B+PWbVfxSjWP45HKkLiDGONcehusYk
VOv4zlMVkUJhvUZSKsagJKvyhaDiA9C20br1+laVpeqCYkxushCsOy6jSNHcc9E+
O1Ynl0OYgsleQCuLS4S1s/fNMnUk1R+8qYZnlHbz8J7iFvWZ3iA6R7K8SNBxnyjw
M3S6nU31MP3MDbPy4Zrob4ky+Uv5aUbXl8vg3ebHPaLl8mrdZkEpNcuLR55aDN2B
L1KKhVlqwaRTnW7rMymYGPGORNzMa46moDy1I45xK3VdU7P48SYwvXcUegbJPhVV
xB0IMhvY/ga26sFKZESNgwlM5sRDoHQQkVC8aWzr8gM76WatudunLzdlWXD2YYBW
YBrKguIG5MRvGALzotcSIiijlFpVtInwB7puHoe7aswrLKJWgGcJNMyISiilR621
yWZ6FdNV7wQg0OvVXwHiUgzTNeJHW6aB57DdCct7NJ5c8OMNMrztmXR66yUKHJUW
5iELf0pThNTWE73xnSdKAuYXLnSdOYlHthbks3jEjJq/yOo2r0aW+U5DnmUK2R08
HWCsED9gGU1QIXp1ZqnrcoJpwL2HeIM1xTuKD3+PR1BRSBg57dCgFyI489eViolt
AqxM587xX4T3sketKpeHTPv+rVBqkh8Cr7ddb/6QI1hvyQQTcspwZzPuWjxoalBE
PvegOwajkZ0Umjbu2G0iAJsIbZaj0GBFyGD7+kbweJI+gHU09NhNJC7usD4hIwHP
a0HKGhx3qJyfF7Hbq35fH0KJ8Jk+fK2S4NFkCRwxvYf5MfwUwpARI7pJK7Epjkd3
6djxe4Lrp5FjDQXbbLy1xGV7S2somU1KWOgTQnr98GmhMVy/SBkIpWexGvwpDof1
cU/us2eEpiniFRn3cRAs+LmteYRc2CvFo016pMkycTMqOcjI6Yl5BRnjoxnWK5jR
KilHsd+8oNqzePpWAmrPXhHu+E3IkuSPiIjfUlAT6WUXB4cN0cXA6Adi0LibDlqu
a1EXUFitzgDLsN8VCp3UPO14IapQMSjFm4R3Ym3MhleE/OhC5yH2plF7SLpfFRfB
w1SV+9GWE0n3x3Jfmw6VlSAmpsKO6HFOJjOZs5Q17MzUYUDtC4ZDruzCCDShsOv8
lNjl5VdV0MiUiIMOqGpYWEeCy6A0nYVXI1KTpe7KKyYuXnLOMvlH/YPrrJVpQoMZ
wUM0Sshei6CiPi+dBCTtzPEV7uT4uF07dDe9Bhb8mcopjNxE58Gt0bLPdCA6NzsI
cLCQKbSNlsHUvptrlx3MAsTDiFsbTDGrl8KxAR20zZxw/5/I1hoJscNNCWuTZxew
8a8DA7zOQoV7U97LlnG5e6yl6XJWF3+j/WwgVan+g34vM4+zf/tzcaKm/NjVB6vj
HTWNiKD3ro690PyvGTp9wj3oitjJ2TaS33Q2JO1tpkQ7AOqFlBhtRrAVQKu+a1jj
AnFJRc1hpa7uXRKOphrG5RyjwSNbKEWQIUGdBWiU/4GsRoqgGpY412X3p51PyPiy
MFEiArLx7sC2c/Ct5sUcOC2pTqznm4XC/HRgryuXm2509BFEZS13bXK+ZPtri4fH
xcRDCsf5RTKlt0BpVWOHXC+JbXH4xPnJOmoXLNGLlI0TcHU6GtdJwiJkoYqNQx10
jK+XwqAqEKzXjaEDdxhneP1iqlzJsX49ohFLqs+q5p6etW5YQaxSaeaplBbChNSM
slWcy/QYoJDzin6LC550QDAbrPy24pEUjhMUUKvRQ2DhmXC1DIj9hxrJ4ZqWYyL/
0CyVQFD/HXNcHh4FYZEobh5lijFJuiSU36u6URy3wGm1BeXoBIUCGLTk9LTvjBq9
NYJwNDsvU4fcldTaFVgZOX3WEoeiQilvqIr4OukCjmch6Wopq0h3C9SutaXHu9yM
DVt5w2T/WwaP/S8ZW9RG+POlp6bpzEFKYeOqwKkgOilN6X4lJqux0E9NFefV//Pj
7efxBs+MApfHN2RqCcr5DhG9mLrxG1FAHimCI2hli1dzF+fFIyiCjS9drpJx11Gt
T6mbZSEiCAiA09WqYLOX+TSmysSLkydPeA5lty+0XoYL5UdHulipHPS4wLpjJCob
GmxSm9goNveIn6XCvHsLJYbkaUOLiNq3NFoGpN9ICmCRpcHnZ7PjBONbQjQ+dANO
d2zOwNHIgmIHpo3VramcNuse9HQ3pNaFWrDX24C+IO1zvfU8TkPBjHshMlBHTNEy
A1Mb8G1fIMJIdEB5WsgaoJvJlVlYTm7ie9++/Mfnt26u4Tsw1PudHB8mhjohWWCR
4V4LM3fDt8KRwgdil0qlTFdmJfxDHuBDEcYrGg54QmSXq6gVeSYtqeKwXaL2cSQ+
3Kr3KDRrORtp6qy78MB4utrTYA6ZTOOsHMlRm2Gt14YFN6OyHAl5EvMxsrxfLGnz
pzvKXTKJwCGxzcW245ClSfzjLtcfpjzVp6gGI7n98CbtKRg2kAYGWixqik5gRiAn
FD8hiTmqOevygNqke3zRKGSKSw2lDv4av2qUkZN4uShZfQl+ZM63CBnQhy5VgP7P
P+cnspxDc2JzMqDaVETe3be82S9qetKNVWLBQiFcgSZadGTZxUuybrAdOUabvtSg
3OFg+sUI1a7llgRjTvAOJKqll7Z1C9XvAJIMPckH47Zk5gCU+St4Om79Ysj+yJWn
nSOCeh3Ue2+/ervAKLuJX/5tmZPAef7LNE+rNMqVqQ/x6N2yw4/usZB35STZnv0o
+XLQ8GC91iNGUOs/MEYYErJfLCNHOq+vB9Aakw43v88I2ZXhmmrgrpRwIwM2+5AM
GfscZb8d6+l7CDlz51kiQyr0R+D8SzzdlTMPOOFoZ9tKotSCnGdFd498bJd2OWcr
5bv9ZyOCdkgcC66tzmXOzXLQxZXbEQTQOr5ZOHimuaVDbUEBnd0uJOET9mEqrMhd
ImprA3W8pFiZ1YaF7sUkGuoo9SlkFHmk8KneXUAD8CB7fFkNAbyUJlSLnM+mMm9m
uDxH6KlVxu2g9b+/jW+qJhNT3+nGfBVoloOdUmPNGilVtmLYFKOWJQL6zYEQ5hxJ
GCPJ4Oy2obduBcd/ClwAhSSh1/ox8YLZ7/bNyV7+/Z3+qVJuEetY4C3QwrA8yS9P
WfqYal+GEOBQQim5WRx6ASbJ4ZC+qziXfC/mSS1TJWGKmIKc14hjJk3724eZSb8D
6ct1ptxSslyL3NhYD0kXEuv7GHZUBe0DEhtNA908Im0l4nZTnfxqxrY7rY9X/4v0
EZyZkn6VAM7Z+GGMTo8hjR/VvV7XemsG1R1IwTfX2f2v72viun7OVM9qQSQSUmWR
gZUGW+lCx0iQx5LtZ0f4VbDdpkND0lhhPUPX7VmRczGxvylo4tHnuGDoDncLrw7l
M4eMk4rMz7CEZ+854siFPnzADP+SUhklZX8CtDOboBSxAkBxTtOUjfsZjZCiMDVb
eiEmtX9J/UYQnrAyN92dlV+FxvwbarFjArV9T14NG2Y6w4pDHABiHbNuhbBUa1nV
WAoUCNbfm6+4mqK7iyqerR6RLmrQ1HoW7ZGG4YMOLjY05lkpOppsAMN37s722aKj
V4Z4S771p9WQ5zfFLwkuKRO4oxiCfSrGVdfYuI9Qu8+G9SCgdVc6PGG/Yr/2XhHw
Usjro8iJWZw8umvQ7jRr/0K4QdhvgKzKvyYCNh58pQhlWY7b0dYRCEvVJNSQb5WP
haXgRsvfMqvJYN24IlNERuBWfAdYIYFAllhmIs1TiMSa8zEjXK5ma57eM0uT5U/K
NRy2fC2mAkv/gupDa6A34S8nWJBkJDFrf9fBgfWgAD1aDbER/qVlk2igk3qg2w6M
8x7WbOSsfG/aEweIltbLrwfoG/5RdefBq9PhtHftpfBEYNgvko3UJvrrEREI0wBs
hUmW3XLkbFOieVt88JojhF12md3E36s8bCFMh6o5N3I88IC8SP6vGmDLQfJ2XC3g
8/WmKWt2NSTWrB7T/UCcaRt4hsICasoSpsd9HpRZaQSD8IeX8JXrazsY3aWSsQTI
okf+xdh1puVqCtTS8ZJuB29HH+vgGmd/YlEFD3GVPN4xzxxuks46xQtmAvItEyhP
9kGp7HSsmhQ/vSTRNL/Mx8iqfzn+QdlRwoT/2rKaxt54GaAj6YYQbrDswjbiQRqA
xFqvobBT/LE+Op7mbDRGHfH8y2oqCjzK8gqO6EmZcPc15yEX93+7RQcZzuzbvdXX
PVHBwIQ10weqQU8kIBtWQ/4pg6Mkmxn76d8MZf9gHmRkUqtqVMvwsIOE0OkA+yao
HAFJKhXr6ZBEwIQ9HpS4A8gvOMUYlwU9616HcdaO+bbBAIFAptDqeGHnopIid5Kv
yalYSRMFR9gqXo6UrVxbm5EZbbjVtxaXqq1ok3kM7wNRdU48oPFCMDOjn+0ic/3p
Y7Njsrb4dzvU/Zaz/vR6G+VQMKa+lON/HUdPq3adWL8SkrpliEXIxpmWa/JMZW62
uspJwyW7Y7bieXbYct7P9pYQKGIX+T5N6KV/irz+La8zz+s9P8ZwVmsqfEdxh4p5
P/QBhAaLmF22jcNkrMOOPTCZwrECjiVg78wG4zZCTsdU2k4bY3cWwycrnivH5fRK
DwNNkMkTUi4VMbP4SWk0rMzIQeOsoI2KpyUGbzKzKQL570K9KRcQWt85bV9kerta
VUDvYvE/GQqjrimrf67sS7r5i0wUe/fUBJAzLUBOlceDo0saH+3TrWXKmY80UfMK
39wafICSgUJZKg1k2jX7Ipn6Ob98ocbc7P93wI3tCZO8kt8+HwbUMUAFmUZ48Bo/
tefEaQiwu2WjhGtSPDgxa7TbYLjUXosMgnZbXuLrn8INPMZkMl7oeyVwvp39QPM9
qL0gNkQbGqAyDj22byrHZLBPj0dUI030rf2Emd4ssyO+B/SAHD9n1JSSz5Atl/Ay
ZbYO1i5YLYzIXbcZPOw5x2xhC91rFKHXPWvrdtZlAoydAVKORxBSiirZ/LkCpk2E
z/Ip9mH0ed+VpU/lAJmvjwi3yCSGKVcWdVuoHxcS+S/sIOQEiyHa9QyCneBSz8hZ
mTpf85xlQHS4rwbfsUAfIvxrInuRv93cWrvy2SUHhWd5M/80Tle/viKZaTwoa7jj
YemASb4+0du++Uk0AbXIMs85PERt6Dqfv5qmBhCkgv6HRTUV8g2NK01prQTSpM1c
G1zYRysFBWpc6AYnBZiy6OH9+NpaChoizxGlGLyJoYBiqVoAySqE+UIZl0/K4DYh
zWOCblsvWkVyxxoUwCNSeq87CHV4sHKgQd8qzE+DGYbLaIpWPVYaj+d63kMSRlYZ
N+xxFiGZ543jqIKDfYebjdCpWsMMXvSPstJYuPebKdEHqCjCbtVzYWu7JpzIjzi6
EIZ6QYrlJ5y3EQKHefkzoGQb1g+DWPN7+N8xRbDZu7YYWAhyjUw43nLQy6FX4OvK
8999ka4NVCCkl5n2cu9MJr749C4Q6h31pd25Oq5ykIizQwqVsZchi7hoMP+WwitD
r0aSPZLmOij5oIE+5VTWTNr3nsBkOCG4E212i+r0Vd/Yv7JylJOAMA66JloighKW
FoIj/05GU73Q7P+G4nKTZ1wDrItF+LzXG+0VcXT+xfC2e/vUi9Qd06/5mt6SOCEh
+GvW6hJQFK21Si8gIyA2Uj4TO2uB9TnvSggSE+bq4QNSCjtO4DQJoHE/MDoyTuL6
kouu2qkkHKDhJvq3l1CNGhC7X1pO273Riqf8JmJfPxHORuUV3yy7CXKcknSEAYmZ
zEaBdMdXt5RhK4R2FgSe5qHuAe2ZZ8qeVT3VHGtFbBCyrJ4pvT3Ks2JA9d3fycXA
yg0RJHwq4lMvTinAmsq0s2nMmDJQ5FTIxMNalrSqG3KWRNtqSiwcigUIgMtzAXog
83R5+0XAhHQsvJTMTW/lllgWbvn9mor7Ih7ox5/GzMgl0WS1BqXpwzPhtXtEIUoY
Fcfp/PaFAaLGGgKQZSCAtH4iPsP7c2o9Y2Oyln1VdNmTDB8M80xrxcXMB76QPHQl
JD2wzt4FHXqNqroPgCrxVEpJvh6MoLFk88bwt09xRMZgOt/+GaArVlTEVO5ku7y9
ErwzyuMqZVnxqJfqlZ0aP16KsfniDImPa4G9Kr39GgDRWl4wsZmJ7rR38//KvfQP
ltIVjj8nG6AC9sEIxK4rA5WP+4llQYutHb+zjdjHXKZpt6jDyYWUL+Tczobn0oVz
RVHQAC2/gsAqDJS1r7eClk9SxAe26Qgb7HmQe8nPcrwbwicFLVDNBJhCbpxywP1+
C2Brv1G+TEtlNynLvHpJpz7uSNSG7Vi+DuskiLnxj6rEFmiRzL2FX3gaehZIy7/z
uAJyXVmbiY3N8bLpMa4dAQz5MIHywMzWrPjc4v+jwYzG1iwQhG06AWgccXC7pHzG
VMklfmB2puilkPJMPBEqaXP6ADuhKtv846O2YG7krSE9GRgCCnEC9IN2JMKTxeWX
AO5vry5MQ8j3LGkU2OStwPIrL6O9e4K6KZ4rJf4nRFDFddJmwW07JziK4sQVBmKK
IYe8jVQCTohOEvcTnWM5A66MHlhwPLvM8lqfgZ0hhyF4+YH3ftquy7IIP7msagTb
CuGS4VxTCvGZL8SYKtKvbzO6FUrYr3HUyMecYhXErCgONPxAmnKTcT+eDjuRTf/i
Dp63YHVIkCyutkROekBK9hgt6quGPJHyr9p+Bc50Y7En0SN3otlkCG2CObazRYDA
ibQj/YPe9dSzoIPitL+EWPPAlQm809NzVyuSx8RPgpp89QgURIrs/+H7vshypqT1
uHeZ9NDRcCZjb89DSCiXrAth+KDe6rqKrduUGqR7CY7338vGoaUY28SvJCde/E1J
fQVvpmTMSOFdyIGh9UMjS1IBjd9/5qCHWJbglLvE8YaZrHhUi+9PWIBk4RCSze4k
RymwP1ylSAK6f44wHbuInnVLdltSZqWEy13wizewXlPkMjyoaVgqCJAXqRPThx1o
zL8ThbKJysGBJmM7s0APUfi1O8ribup12hCTw2OfyFPxWLM1YGD3QopiJqUYlxRg
tFLMqPIHkL3tXgTMskmWGNVCuqc0GxRojpeHspUUJDMoSgCEJkAIb3nxhnwEaElA
JqvAi7H+eccVmnAAVL1qJoiUdPVVn3XE37AuIlFCGNGU/jE1hZxNXNIDw/WPcLMD
v2g+X0aHNw/k8TEOr6PdlW4dYHEldusamW3/eFXu7nhcroGMaU9a4OWjILCWHnpX
ahaRW48iyqYhNIw2q8dR9kgGyvleDvRn7PoctN6zTCHPf1ZOQuvcAhD40Ocy2o6N
agiANFMf9P+DrRJq8X/8YZWx43Qey6/a4z4GfxmPsNt3b6kp7Dk2RRgzdtTan3yh
F8+N7LLZP/6Jfl+SYoPflbXzNUOxCk0N5IT7tk02G0AxQ8lGSJiasknUlv7rSA1L
Z3dS0Agg1QrX4eh6OUICMoBo/u5UMJkLllj2s+et/DLmo/MNhezL0+WIU+YNvf8X
gpCxHFP4/eUl8BguDIno7IK39mGVgLY2wgkn+Xijn+cwLqjBiuI2pNw/lf3sZiBY
+jkgDJ+dvNfKs8rsvufdL+F7Io9ZHxNfkcSIQ2GsSyjL/YDNfGUo2BtNhG469Fdx
jRh5v5r8aR4avJEwZGTjqmO2JsiSGvpqF5wFnTvNw3x1BnymnBrZrYo2bpj7lKfd
q/oXgyRGUx8xSONrvnDs82QgcLjpGeB86Qn9eurXyUyxPhf5qWMUXasEE8MI1GQg
+OYoYMTxTbHM++xvUhpUB8PPF0d0bt7arv7XQSh4KrhxVHJQYncn8NjCiLtU6hzW
17nLQZ8VX2lM56dmN1cXbj762JpxeHAgYBXY/l4X5xTeg9T6zlify4N34W3lgq/t
O0fq/Ydk3N/Q/N5k5r74vfZ2cOgQ1kDkjAmJgz1siGawNz//phsxbttuoZyTmVq+
mvDBJ8GyoqUfG+Ul+M8N45kajA8BXtyy5Enp0RY+GaLq76g3YZ4YGiRaNYGsehvw
fx97xQKbV6zcuDBoeRBJdxilrw1fco0DkCJ6RR26CnUrejFBmr2+ft7Ixoi7zwfr
C+O9cte48ac5OLv6DlvIMdkyLcmHiwG+cWIh+SshHj7DGTiTmBEm/9fdU8LEsjvo
au0nd7IHvci0Wq5xB1iX2Ek0SNHe7031F72gktBjRpl133YaPSsn7pwV49r3M1OP
I5oI6P8eI0qAzfL9/FoEr8YjJcz9U+bpcCN5dKL4GeWT8HaBQ7LQdfyiCR4t4A0t
dGHdS1J0uobBxf5UgAw30r71Ye6ndEso1GAN+2+1l643eKh73Y5hK30vxh9Df5rY
ITfg8FwA3uz4bhbhMs8Zte7erALCkLvHzekqp69I1NxyfP/4ko5r9Pv6u0sBU0dS
3yu7zOw6z/eRbmY/v+xrAO0+HkqSDkkOaDW+ft07WLFPl0fHXQMPouQaoG85MHq0
LBMbmYH7XWfvxwSZDurS5Ad5LxBlihZicFceRlKit0jJGtUixbBl1Kh+OQoQA4G4
k292rvOyyEfWek+vauVkPifh5ZIiKI3TaXGPNaS3CsEKSp2wG1/ZfKMsXcMIy2US
kc7U7pmpOJmywjREgw8xFBESWZZREqicTKBMi8Q2gSkShIwY31JFDuaNtIYwlkoj
2uCbx9eycu+9IxB1m7fvPRiGdRGKyC1VFGtopwb9qaZAz81cPaiBBwPgxD8eek/p
9uxdhKHs8z7EisbJ39MVvGmz0pM16vXNlOJAQfDh4UiPxPxQMxVicGWS1n29Ypte
tFZ2/BfhLEpp7TzfDXC1nzGHBCc5ytTge/VecoZkJKThlebz+pZJII52t3Zg+rQv
q0/4Tfb/r4qrl0csbTrdElKo3JGkkhUV5lcop9igijCu/D8dezf8fb9d7TQw7r00
qepSnw3uPx4FmnaljeijJ8Bu39oOtAjQGjPkXV2oMY9GeszfoD/O+HJAu6MQ7Up8
wFXoNAm9ndiFHLzVjgF3SllV1oYIJ1y/a3I7OugfFmBBiGcX9Mk5/i3r+r9fquFU
/YgVgf1uZI6S52IaQVEMJM5/MoEeQ/L6fq8872r2fI+R4zMLcpNgnzNDcrLm4G4n
yW9/IJ2QzsAVQUeoHvP3deMtPQCf8QcSjtL4xyWw6Ip4S23DYSdjO8L0dikpwNki
9QRbs2e9yfksqg2FaTpMo/hVEd1Md6lwO62DqShCb4qXx8znSlD+y910Uv+eScFA
qm9r1GAG+3xC7WRwHDYCYsaKf2DWLgDAe2V8m1OxN17CxzBhsAUCu9LKbwBeRjwr
ajBB2CdWdXNGoOSlgIIAoLaaijQrjc+yk9BoBtwyj4R/r7QA1Qd8ND6uaeXCxM26
HMPxrBAj7crSHo4fiOJYlLBWUr0KoQCiox+qqcUuIAfOlINrbrSxWwloP0ADUb7Q
pI8kRWThFYK23/MUvtTiJpXXkniO9ChG2O6//ZVx9130jnWeObv/Df7eJgCV8xaP
lh41Nr0xP2wIkQPV8mZREP9RfOyCBMyhgmhVaPaRBHgiv0oKmZSIVKB+pDPnw3YD
f1kpmzrJnw0t88FkiOF5osivoSfzcTb6OLdgw/7hLxsjycECcHpWt/3WXb1eBFoD
vJ3VZLB5AUxDP9aMQa+uca8J4W3eGWXPNju0cj2OwPnbGM+CpLtjZ4i+6OdTZg/B
995IVeRHisQCFuOMXadmFV9j8TJ8M/s4/xtHkHvVupNNhZq3OP6xykhjToLoKK5M
QluXQIaSjJo37rrPYzWx88HH20loBdyC4aPq3yA3VBmzYgkp7XbTihnojPS2ef03
W06yF9CelAQwAkIPZhB6n1pWLYUjkjbDWHI+xfG4sike56Qt3VDOh0LAyuVp2dt3
kJIPGMdkR3Rb76M/BO6ar/XItcKkckHuC6BbUylJcV5JjvdNwcAWjCQNMC0RvAOc
9WlqBgazRuyavjG1BBnAUhVVmFIpVGWELMLw3Ad3ZAN+sdTFyPo6J1trxwKH9t/N
kA6+cljkfYafkZTOE4VSVGQ4VYEI8PKrhE6xjOaA86/L6VQKXPvBxG4q8AinyoSB
KrGeICnARnHZK/UiXDgfBBeMqgm1XaPwN/i4jOj6atc4jMGkefe1exvxlt/Lzp+/
udK7cm5oRYaM5Sg7/ejVc98yLd1KwBGnZRKj99RbCQXMmLZqNO0xYWThjIUGpMJ2
sr98l9iQd8jXvp5T57UgqQlUNSlLUeN9GxNdta/N8UshEKWpOljAgfL/ljymVkfu
TwvCWHZjmZG+A8Fl5RNm+QEGqNidpjIGvHz5p7QjCcEC3Zd5DUv8AUnunYLqGQSF
jzD91keiv9q8hZ2/lOHvO0zkZ1gUYNPHJ0xCwzSSxwuvNdgMFkmkXa0wa2BK/TXS
Z9yJZztYJRpkPYvLNuotTC+JrBpLQDVMGe+nw53K5yxISIEOc60Uc5C5+nxn+919
O8Rev4RBYV2OOjkreUFNctFTwKj0pnlabMh+HsB91jJ1chozbE5MJx35HkWqoQVO
c4tiPzqzvJpmJlPkIaFb1mnd48FZcZfdWQuB9UNpHsjLkAx4B5Tg+1KlyjAzdvoz
8FR/epsGTnoKaEyvUiCXstx9bSB91Dr5pTifhNFFiXviSdrrXG94uAIsmylbQ+wc
Ws1qJEuAPPGXJhx5dIeicWbvh+IVr4z46rogkm3Jitx6YQiockOCRWyl4zAIT1Vh
ol9/8phedna1g2V2O34ESx2qR/XbRzVi1avgmFYfypSY9BCh89qz+wdHyVeWoRu4
DfIRDQqxGFhNY6qqSI1uLxVEG1Xb2agRDUTDjQE55+m1ibzZrud4UDQ+Fay0VnPD
dOlWPzlb+JCUw4vF1QS0kvfo4nheRGLttSp/RyxwlACt/Jkumhu6ygGsIIkAenJ2
RrJjWXM8UiPWecfTPZzr2XPK4W8+GHopGG2VqT2JjvrhAY75ymH6bO9kSLimX+BF
jFspoKZnMdBb0t3GoQJ6q0TTdW+xouTzr4eyXsi6PHMP8nJIDYUoe6aBK2EA67hJ
dGf19wD5Uawrxgnv6M8fVyhzwCk/vSkj6hxoDxkZwO2OnBPDdT/GGyCbzdF6Oroe
e4o6iaARbOxMv143yUmLkhdUhBhTzZI7rJxMvfo2iZVdnZFbSXPKZQ8v5OmQdaU3
0ZIfNu0KbFnKvFD6HjdPo/EfpQ0WK377bMnWz/n8eQpmnDhUqyhBVOzy2YqYFnGK
7MjQS+7aQYKT1vjKlphLEpTpP2sxjGoXqK7kvJNASx7ipEFBiZ4XtwEuA5+e+mnL
9mwEmCGuOvnHEVO4/UlpYuJvtkVhKJz3FmrHN/3NtM2GbICCGeaO+QvLzpitAd8M
f9Uz8npDqWvVGj5uxzt6VXDjHY0aLsMlfNDUTZm4VsnAGuBZoyHRAKDhRUYRHqk7
Go73I43BCapxXkhmBan+uPOB7XoxbQ3+bjYui5sWL+0cldXwKveoI5Ob75SjAcHU
rchHdZ4Zxk8x1Wa+yjTO+BkIFKr8eUOiBBn+mSYFrqwYZG511uZ4WEHFdGQnAXAz
R+sZJV0sOVf+TVfWXUp/pY3u2PUATAXg3Jg2CU0WBmXctQZHpa0OoCkFuS7YAnot
VRLaBhSNWbPNygERFlf+jgam2Bvsz64+ACR6hr9kdqsFrZClsic6BcQZBBD5cvUN
r9EgMBzkwtFRFSfTKRUyB5J+2vZ4scMZvL7R9qCb6qcQiyc8jFbPyMNX+70rYYNk
H+C2o3+jr+Z8WJPvtknD774CQu3VmGjG7UU0zvEeqpJ8Nc3W6IJY5HccKYnTOQrm
O1Zv0j4+s0wRNzKjGBqVF80/u7qgso4f66rDsF0hMDMcmXrXXuuvPpHSVOZoJJTY
5J/j/Ah6BPaM/lDMNWISYQ5SlFScR5YeGhe2PsATyaiRxGBac1kxTuyKIZZqROsq
g7EsxS+9/gufsGVUYcENRfnb9NR9WHEPJyP0HwXyewy8kIXTpWy1aFS34I//F7G+
qMLjfbGCxIl0ip2ZqQH4UMP3suN4jOZ+9TSxqwiGh5gpMFEXBUb+DThwYHUt3hfK
YE7KYsG2TD5PM0Z5by6oUToU9zvOzRlg3hBDDdDWFwh4E8/E6JZTgq7VvUDvqxY4
wstlXdEzb1L5Hv9wLspw48V/eSgMI5DeAn2aXcv5yn21xyl89WCgfMiDuQhK9YAX
7iH/99VJgF0T2BMFV9by0sAkSK8FvH160WsT6akDuWGLkgis8TkcaXxe8pL2loJR
ihTClSxKKISDDqsxJKrzGQFylgzYIpe/sSZdPrp1oW9lDgiSN1jNTgi5XfwyMXf7
aod6+P1xYt3RmPV9vBI/l4gJNtNjB4+8IB94hZjqeXkjmNp5nYLuZkpdJL6nhwyR
Xye9vhdXSXvmcpXLFEvvWKq14wlML/hqF1e8l2BiXEPEKJnLJQ+iNoDuOrL+vlgL
KmnpeKOIzqXyGC8CoXKJqC2IOKtt/KhgChDbsHYc8gz/p2Li2cB1aVxXMDdEAk4g
xwm6ldZ2o5yRacSv9unu5eWpTAXqYF/NxZKtmyGrzRensfSu1mXik9eAernFx6eb
thjV8jNTUAMSG66Wh1bMBghwpi7iVIlFl2LgIw5/409vHJmDyJmxif/tgoIniczM
8JyfebBcrEjBAsydCwpY1wt+36TvweBDI8hWB7Hee9iVf1R5I3sA8gqcYn3m6kFW
E7aC7Lo/VDF/QJqP0/rH5nSJ9ReXf6pLciW/WaXwLz6mDzNFKQuz7RUaNh1DSvdt
0UfAlnfJ9rSfeOvWCG+rEr4bKeNstQiOutEGvx26SAGsy9nFcwf4FRrlwRzFizQX
5XUpvcNz4/1GO1OQzp96lWbdJciPyYlxz8CKrYDJBAZEktPKENRpK5fMXg4WjZeo
Aeicq4rw3Y6or44dqTo8QKLo/Qs4vKq5Z/V/mcxDTqhCAcZ7nWYsf6ORJYzEY+bW
gk8Aveu6V9bT4J8byzZmRW4qSjMYg6E/e8vBpmFoSpTVJZO458dgoBgFe3nzFCNA
EnDhIRjsUNNFqA3n1lWlURu/a2rU6x0WVqYlRKcmR9UYUHBqht9tMX6Iuaapv/9e
0v2AHh4Lj1Say0hTlhVYD3tbb03g42hzAx8oahG5ZMx3ebuUTruyG5XDlaxDlm+J
TPS3pthMs8DQFExoPikO4FpD9ApQy1zrYFnnHZTwWbsZmsqxQtUs9DE4wymYvDZy
LyQN05VISF1MOB/QTW4UzNwJTmG+vBTG4/WSQCeVojW9YLLbg32LmGlFsepMlW28
UWO63gUPfbqDOKYgGh98yuHGRt6qTF3EocsJdiSup3e6k8hHQ59JfuDYK85ChheD
wVf/qW0kMCQf3UiVotmojRhbJEfze60/vMgDkuQEbyVbkIc9yR5VTevQMARpSM5s
ISjmC5gB3uCJTj5U0l6aUVoBQgwWE/USvgXbIadLvbgXNwpVsyU+FQfqN2X/vHfn
a6lmJ8qmAFXT6YH8OG/+tMXyLxUTzoaj8UTmVWOG7BWNS90plwhhq08kNhVy8kjX
PklIxlrrkOVVsYhw0Nk5y03Q8UIbm1ICvRS2XBlzLy4KW8+GUyWmM+E4EGgAtmxp
PDcdRUjLS34tpzAbrdjnrYnL0Futxkq73uIuJPwHe3fyjN5il5cS55LWJjnp2yeV
L/a6ahyljNCYq2npDJCPTw/UDWzhbZu8mc0FkWxXDIWctRLalRLRGz0dNH9bTTZi
KmSseTpTRhGCQfgq1v19jfRp5hPHkV5Oq7B8JkNaWTST2/Q5sZNEkIg3VxPBFJvl
FLR0WQ776sLoQlneUT9ravHK7ecd9N92W6WcRbC7xT2n09WOWALlSxW44/i0tvlY
yHZP3SHMe5Dnpa2Blm62x+jwDKVQ9YDV7IM0Y0fBakCDRxQpHyqQcly2i5vDW9P+
3SOxjdmWO8+s1zCZRuukKYRSNz0/yLUGjR1Hqm9ZodEtb/xOJYV7kcjVEXRwbMmS
K5eN4IpuSXZ3/Ny4XgwREWHuhQHFKxHFbaXjYar+yBKmiz7K13cz63g1L1PdMO6w
GwRx7JUUziGZRAF8cIv9vrK54bx8avhSgOhc/ESqS+o08KYt6i0jVMhSaLtfoQd2
Nr20pPgz+pZEzgtHoX+q9zTaQzzPFsbwDBAQY53w+WLvAsfxmov4P1uEVAVHbhvX
JzTlEodQOxsFJ4CtLYKQriMjkZpaH7Mtg/E/a6icABv05eakIbMwDkTmxbfWwptk
D6NORdvaxfc6QLQcdxjs1OOCmpj0T84w3rIbNGiupV9vVOBCbKBNb7C+o/py3Drb
3gtjLcjgFJMTUBf7ju6JKjiwSXPVLXAnKHauutRe5u/Q7Yvbx0d10yjWHHZwLGV/
yEZ7EvWXc+Sunf1mpILEcJ143ZsORU5HdT1jCf4VXfuVheWRnMUT6p4RF3WooUPy
otKVlHctWHEezXaysIoK+EFA3Uxt4yJ5PmPuQEMctSvqDlVS83RXK49aaOqRG6Qo
oq60EQQ23XiDz1a3IrnSjt0rUDZaHNnS5pnqE82jVlr2ZQwhLN5lmlwHOz6XIE28
XQ2+w7gjJ9gwiJHOmpQcC1DMzYYMGpfapGLLfDMNZQZ3Wg1ziZ3Qaur+D6kE/F78
f+yxa7mtqrcFlDe14dKlzUy/HWzfIE0GVKLNdYq3ObcAHlznioOM2w4t3PG9sEF3
KJiakJuFT99RtpG511vRZhdPx2JaDdb9neQ678vo89AUpu4SDU5hlnJdM5EHcrUp
9WVOfuv+q0JLLk2dmKSFFrJH4kkfV+DHuU0XCQF42GhZZUbR8Bc/gN7WTjk2VHKY
+NAFHOZKUkXK6y2XdN+dk++AgGYVi3PCSGaLxKnnebXw4M2EX3xegoAawpLsyY0g
+ORPQ3lcw6KvcLhA6qZvrQht3xDQk2044aquBGuwCGblfvHAOTHyAyxH8L52D8+Z
fVFv7B977v909XNi7K0ijEbFtl9DA4lpw6gL5HXWodur1F9T3Qay9eR8JgT2c6xk
7qiCcoerUM8hlJfJGBPiMZE839R8oRrvrWAT98+M5VLL+b0/Roc0ojLNvTpqSzFr
aGTp5tduLuUGF6xCLkHLqTU/+zjZcfXVAQnpeqyD+EbWEZhLEUfWBCQMPFpuPq6b
Oy97bn7jjSjP1MYg+SE0Zeh86QrlHUPby4qvtOJxLR+l6b+vO3yC7o0D7T2JJf6Z
LlSY5aizuCKuzHUGIs4yORIt6T4kSf2BuC8V975jl7AbavKkWIVmYY0AELqN7Vxw
iEBNMXjeVkSHI75ZZYpL4qEPVSzzNIxpiyG2Fe3MiNYYZOE9l0SAO0Eyhh0Lxwmz
P1f4Q/38dizCJt2Nt779F/+su0ZJXQff+6Xg8YNSK2HKMGWqgYaVqoC1awYzNQBk
3yg9Z4W4jrp8UN/9dEh6ITCpHIsDqeXUZzH+Igi6vpwCAZP9ecDduxNvTJ4m0958
gNc6ZIT2bxAmqcLD0OnqvqNoSqKumwC6RyXFpAMK8YjjTYtSB7EuwSSoTV07Ln7e
0wcOgR0S9oFATSGU5Lj+YS1VrZPacQnN+AYgRQpi+UodhGBjzocEDcQ//Mof1STg
uWLlB6xp+fdvJTHj6RtXC3rdHSHdTzFceh62v/gapei/w0sMZsyIYOFRjZHnCdAz
dtDzyPnQzLWCq/r5EjP58VwWA0E1ijtR0yoalYznC/6H8j6AXk0xNVqpYbO0CEON
czpo7uHCdO73l9pDqStAa6TNIaBw4BT3Z9x/03ARIwVDDOu9V8FUTJbCH22LEz/J
6+W6vMT3A+/1GZSL9rs4IorJCZMrJop93UABLAtdFHbeoUWwezlPe/XDFEGZkZE7
TyJDY91TyalqhI38eaRCXcC4YUGGw4L8U0nxcJcRQvL3d6H/Ln/Ayf12fAdkxm9N
da+hRdfUeYPgn5jGlgA3AvmjGAzAgZsM+ce3F9Mc4tPXW+8euHp+0eQ/t15FmUnj
dORfl8jQu1SDqyGJ28D0+pwzeQy8OibIdNF4kT4Trzt9f0wctRMzusGlD0eWE17V
Vu3BbsBKaMdRVAKVUTnzLJztA1IV7yH9mUw/hVIrkjlINL9OFcdwPCWotChmeiHz
yHdc3DMEyFUEkiBy6jxW4vJCPgXHGUPg3ui10+5bfAm7d5Xbxta7craYJxewAKE/
ie5nMxaRC6jxMD1TP7bBOobnft9Zdkk2NWTUTVaYJ9Hr9/Il9hPU6yVdnSWWnpwW
u9R3AmkHGmvsaSjlDnBeeYasgPibZrqbZ98Fk8BaxOK5Y7hD6g7mx6FFIdnRPBz0
BtUuWHAKoz34tcHFaCQfTO25ipNwex8U1XJhv+oL+Ui+0uwLJf8E713g4E9DBdlk
AfyD5rvhOxAKXJcqB1L3MvoO2jxO5m9wbmzRmBiHl5XPS29TERK+T1JRiOtOM8Zv
TZOBo3LbB1eBwKBoylkb7PVClJFaolbyVuRJbx0Dk8AJbIhwwVTO92/9hQbKyiTB
IcdGFOj0u5nZblg2zwcF5PgjKq4N6hgFTKiJiO9iGLC98az1gNGunJt4HQRsg0C6
BufrztIohNtRjKJXKhclsKeYGZZHRDKRBBu5SLaEDSC9kRT+aj4A2ADRjcGeoLYV
Y3OZSF9woYqHjncpIndYvAF39RKQ50J0lnS3vqstdltCV0I26252Rl+5n24yjcIi
ljIVTdF7zyXpRJhwHJipV+sxZ5EBODAd1zO+sbJw0P2u093DjMmKD1tJ25WHR/hx
RkFNaKGkbIsVoarIL570Rs2t9y1IEeHIriaz/LmMC2E33LFgC1URNBWXIKA7zKmJ
LKw2dGUeaHBpLbZ5K3qGmjRqS3Yq7pCE6wwv+YNdR+Uf3sn3xY461wgTyRF8WLQX
EgrWXeaA/EfbeYYtXNb4JOHOyPhjyG8bXcC2K+Q3fxo3QdOpzX4zYDGXVv2NyJLT
mi0iWGluQRxTgaC3JxLHYyCVrABrRhdzPBtYHO8S1KkAlkjGoZeJgR8kCmBXfpmo
RCXUu++h7iaiK88jvpIFh+yNqUvj/NIK/XXrlBlrkbXnM8EJpeLXikjSfid7tjXU
gfxMKDfmHNSVZuK/bWgmrCZnfgEYFOayAAKxe9eJ4W/qF0aewWYdTn1SSwpXWMlE
IuQaoRefd3qPneJbPRLAFhKrLeROJ7OWDrhTYwEy/O2NfQ61MYcyV0EmtkKuSWW7
lD43FBHlh5rSFD0xrF2ntAHIOFsiziu6I86qxd4xfExEhfirbPnq8dFwQaFVvE1Y
DiKjXh82P9CTmJIStShb3TUcJ9Sqc1dapZfln7HzCdjsaOO1FFSidDEiLkts1U5u
iFG5FR4hjh13/0LLYv0HjQy0AZKNc8qu5LyU5mkgaUFBDQji7hDwLAxxTYPvb5Ze
9Jpatjgf+4SAOprsCn9M5qJqG5oo9EugRxlIEiK32xbNHKu/m8LG5DVDoDpi8Vo4
ciAh0Vm8vEPi14gGOH742hC+1vuRP0nK4IgbgD/6d0ztfwhGYUDO/zT7UIOhufgZ
L0kfUZbsngjcCAPRp0kyV+Rt+mC1qW8VHP82ipuHH8UIQAae9+3Zard6VCUQa+bU
egxhLvsUm04oGJMFbOHpKtRFp8F3O/Rq1q2vZee3WPcooHsegPCo8ny0nn1S5FJ1
lWNiIDxb6S0T+BVF2iHfwvy4gkcryaBo2yaJCBYeSyISscFhhhgB3GG65VyyOOaf
0YD99cfv1WIkP5W623NDUD7GaCBiDaG3zlLfkfPz60gI7Ghi9LL9plbaGT1cyCw/
nd81UEV3PVWpBphz9rZm/qi+hMzThnZXWu4AUsnmoLlF0uz2OnY1wFC5QTQZl+3h
sO7pX/x/wheyP8Zb2nook0fYJH2pE+Cda6jn0XPw5ReJ7azKpzFweav/LKFGR/Zp
lqcNo6/WY5xbyRqTBn61MTmcnPzPEIcMMXSMpUhRCW9EoAWm+v61lhvgy9c1rP3L
JzDXAkmCiBO6I9+J4TeKE16W7f/2IeqW/D2K0UK15GHgxpr1Manc1jDoBLKhx88N
NUnnE716H03DeGzlKaQqhk7AaaN0DJLWkHlSAXLmM661pp4avsR1IZ43xk2NOk6E
Z1rWhcc6wCFG4KoXN+1BHgWUJia64RTGq2uNHFmFOKEc/vRWpYcZimiz5wC6mHkf
MVztdI8GTZw7O5j04JLRIs7bC8XHDPZiF5WOxJ67mhDOxH7w8eBBMnfWWdCwD2B5
p7LZkeS4CHTMzECzlHBj+JaLydRaMZOQPin7vGTszc/QaXGch/SMEeLTpWNQYsVx
lgWFPhAWdY1hhqP9KLg/5Ah7OeDx0zeXewoUlvK1M091spbLw4+AYt8U/V8wNZsu
Svc/i4CSfv8n2jb2ScY82oEKo9NJSd2xc8PPtPfSsfOc+ihcmltykRF/5XfzBwwG
fcJzn63HtGuPES+EzF27oU8JGaPvT0EEM78rjcq4BdCEJ1YaiEK9b2k0RL8FIWT2
oAJVHAYgWUI0dL92n5vaYb3BaZC90b4QijS9eJM8nIFjllX+OkBSznB2OG5NmcjP
YEfzXTgY58WZsrc5rSvpNyzNASWUN6+/k8BpPB761Fpj7FKpCnGqejQVBHVHGz1I
8ljZ8hf7HYjMcBMoh4jxENdXMSQPXgIOAHXgAqJEUGl41px7VtaDoLq6dli9n43h
+oGimrzKKhWUmwLYcDMxbHSBmmNUgkENcjR0eVh7tm50QrMqRERhi5kwnG8L8tg+
1rLboiGYqXnZ8FgMEcpLuhPteSXtYa+WW1qQUF4Zj3fwctnEuqLRThoFcVsHjC7b
YbPOse0PFMeTcSpOXNAsDluU7dXTIyljuF0CjqsHKzOdwl+Jr5OCo8YPy0WMw4I5
ADOc2B7lmwoCMLNlPzub//RJAYwAoj5QxK61NjAqUtHWAhoQ+wzOH3BKJC0EfQe7
4Y9nNg5HtU28/aERw4Mc3FsXmY5I+2M1brDBOOtx1v/tAaWPz9HEofYr8K5zfayc
XawRKn4Og36OW5W/4ci4pGys4BkvkyQ+GA5OVEQ409H/LRHCApMXhO6vLFDqhPbE
keTOc6/gCdDsckE8PQY6mwYoZJbswAjAZzMccPaNtrC3d2rqppdP4qoZ3Jkj0ahB
jQwd+mqtfqv9Tgl0PvtiiLhlfhbiTTHg2m06holyEnIR+ZWgJ35OJUPq1xs5cUKJ
u9gv1pFxrmiUtEl1YY95feVLr0x/KB7j/xPfGIqtfPALcMoQpH1pI6CF790lFinJ
EeeMIaPwwOJnDSnmDsTngz42LyAMWjM+InZ7N4cyYNuLtWOAL8pyCtbXys4Uye6T
eDlr12JXQC2Vs1qW5pE4s1fSYUfV/nRdyDD7FnDhHfU1x8UG/p40HFpgCVvBprU5
9vQbpqb37MkqL+AwgeVmMDvvf2AhOjIdRFv+dA8Aibwgt3wkMYtzAc7vG/3kqgk1
E5b1g3+e1C2xdrXMg00EZyygKx1/fThwABGOG4Qn1e/eRnIjOWez2MqpHLTjSOB1
xLhojTtSh3IlQQoNH2h0LvQoikcnsxPuhUgOaZCejtCWk/K6sZ3mIkYuGLS5ROCk
6H3kDK7fhIsmO9RyPxfjxmOfxAyVXK4l+GaYZjQhH2nVGMwq1hfrKUkLdiAMc9i5
qILq0DSXvmTfAf5lq7rcke2pj4lX/falPJ7yHhuA7yKLfZYBMbnti1Nzd9xZk/XQ
pmW/p2i6jf+XvGcp9slNzgME8ARCwjSZzOElaxEjOEIlZFxSS96kaiJNYIt3sLZe
9Pa7RXd39SVds4ANOjHPuFG/sTgDBQ8cnxogDsmr6IFhGenf34titx1m0Wt1/W38
iR5X5jFPvqlEkajB9IBn08/zFX3FGmipKrP+uYL3KGUgAvYlUyPNOEWiPHhvULMP
+LNl2N7i5ci+4GHDVR3uWkhr6Cbz1APzvedFSmyet3PES5r1YrpOAYdyfAVoHfWK
IINhpLp8J+75UxBDrBdhgT8xBAZH52J7CqiGYdQdbarXoRpKMaj4qyc9aVyehRD+
CHu66/TVZlcIzQWVjmGWmKJF8EvABruZJ7oF3PW7i6R6qMz3J9OqG+8BgoyZ3tEi
SvLFFnAbz3NRgXsanRymUHm2TTHIFa1OnOUkaZdMw/fkqK7nUrKnkgNsaxYg92zc
+kYMm77LWd6XHJLI81/YdbRzawcfvOK4l/fhwY0Lel7+qIkzOmp9l3gdg4kJdTPl
KQLM1JLlcXWafitWXLKnoaGPUunkkhoSKPmeijoJYPA8upJr1B0nmuE0VsQjFvC5
sNWBhjGFU1jPqrygPIdCk1HQCUVEF2kS/+WnydPpsET7O565Mcy4Xsa48Wq31BZ4
jskvyTD5/Csgb55Ht45PI5sc9qT8TEW3Zq92SKKRMDTFcSYlxxlOkdNPlxnR7FyD
mnI5fyE0IlYxvc0pk0VVkxuJk37CY/tuPvtWBqbHDwnOfzNA7DmxACZq4UnvgUMk
5OUwJQaWh6SW837aBKu/vF12+JtSojP/m/Qp3Epdy5OTNOQ8NvKVnf7jvOTM3oc/
5ApjLFeKPr+dJY4yhPehfF0xxWUqG8eQhbUriFVMEkUcJizIUQEmh792bvi3rwZW
J5qfrONdXgnPRMl3Q59HuPoW3QRCFm6vz7HkVw1ZlklgjTqcybFbLuBqfhKhke70
H9+JYU2tbjyQ9AODYZqq9nqZQTYnHepp/wfYi/dBTOSrSqEPD85yjargutd8z8fR
wY1DHvD53sQXHtPHmTZ+Vaa9msw2ytE0cuDbtnvEFf0fYY4cF0AaXGsEISckSDn1
qBqRsJvszMxLxhIEGcBkuC4KjUPf/odlgh1Fxaz2yapX6Qq3w9jmS8OG/P1TBS7I
8V6ENJALfhsh5R1KyCEq7a//a/b3dp7IXnjfwyX2LUBe+9+qDp1lgICbgrSttiL5
957qMjqzQ/8z/WL3O9nUL8hhLguVCE3lU4CYgBtP0WOkuMuDmbQxnPGJqhQr8Z/W
+vTqsuBt/fWQjf9KaJQldWi5bcLvWQUevZJ6wqfbvPMvjemJmFjVhkWMpEWHZijj
DoPPb+Gfr03p72LTOgmg7gIV91t4VnVXgDMOvaJb9thQX35+37W6T3JClao1OCH/
8PHy8x8OfwegO8CeRa+R0+TlSYYvY01ifH3zRDltm2KfIPpfXn5JUNiiigaqgvgN
nE6p5ilDdZrgCGn8g2FX3IZK7/VhzFhZptYh8+XhlPWl3/rrrFPvPbYoeRaxqZRb
ciXUfhMD/PNIOLFhlu/9geTnStd2dtYiKrBbxq7VCwBShfDCfL2XdjqfXnidhqSX
68fMhe0Osscu+cy7+TdrHD6w2/WLjaX8yUc5mL6z2ItW7nunePZOqXEKwJ9bXdCv
S03HFAN0P/zvFt5i4TatOgJGRg3W9plukpIksI564aq5U9mZbVRDXuhMpWioQ8nR
YUmHhGStdOkPMVZjQKkyUQCP2bLN3TFsNYkGLLX6U29FbJ0hVgb6/9J9ZDTpjxDE
RAWIPYxT+6fFxoOIh6Lzohh3vfAdLBLsESn3OivxC2JK6cpkkI2pVqEyhmYVGT43
V/FlPpBWiHpOatMz8Aq3ua3tUGREmE1k4vKSfgsY2c2jGPZizhktYUbvnn3BSpq7
39t3zb+bjRiN6JRFVVcpu6PNk2Q2j344/Z+VgkYnUjSCMmpCps/953mklLv/zPvV
t63CfPXV/croSgXXWV9pppPLk4sxAInzvdn69VvPa23E4kVfExzMObZxWgDOL524
lI0JZlJbzAyFJPRW1B4H9YiF1mCEJ3MqqEAry7mspHZ8CFvKBL4AyiUDPfKL6mGl
Oli9D+Zw2ah/eK1cpVQYrFGurX7/8KxyTyAqA/gH0bb5TrSBmv4DGCw3RnSU96dO
P7X6xK/ChrGpcbhgX4Bzqk4QetIPXI/ui/wEBKBM1LMxoCIZSsyReZsoTKXZshZh
tkzG0iG9IK5dJlHRgWSax/Mt5FGc0AH+ou/KTPN6op8ka7T8b+Ac9cy2eEEe678d
mnUUmHg/Z6KsNAWKrtXyeuJZgA4FcvdhMF+xl2IBdSxXe44P1juL4SLpBO1VwEiB
fn23bd+HdRS9i3APdoBM+1HyQglcrfzAVxhyopH3cxzrw2jbQXJMj4T+oyy67sNg
4X/feQdib8kBfKOBI2txe25UHWj35N2s58Bj92BsYxbtX/28dD2KFHdWnQTeUMUG
UqezNqmGFCc7wBNDykzx/Ihh9fSwiD5OA776MDp8qHiYKgrGcTk6tbXtlPIkjyNH
k/qLP3qJUFreU3+zkdflMTPW35wn3cPdcaNpKPOcQVRkE1OvLko66zejDbMAuxn7
Fd2Bc7WK53WJA80OmozQh4J5Wu7a2/8ssL6Q6uCiyDGWqlgIscmgsGlWhMYJy+6u
s0OnELVj7McTBqoUsca/OOZpDIu/9PegTKQVqGri8cs4SXgR7yDyIvnyG8wzJvX7
JQpqURTNTM3FeqbMShJF8YPgsPDarAEO8XHwaF/eeHSXoK5EMYQRWWhffDPCBM/T
azk/AQ1HbM0X8LGHxsfx0F23xsCtMtRvDPEmLjEmtX5IC9HSqugJ76y9vhfbSAtA
w/P32B5FjoglpxRhHRCs50iWO3EBDH+oXHiFtvmj/7GtxoZfthzKYTpEqaNPmzgk
VEFjk3woUouUZsxq70T4ZpQV/VZ/vhAjeyfciVoCzXL6W+Xs1OMnxL6viSvNbkZB
6JVDat9WaaDu+NfaZXj+Xkwgsqkvni9/KCpr4kgM0n1XhNoyDH6y87IV6qxAISYK
rT2Tognv1UlNqJm8TU3IBYEEwpHuqT5BcrvkmNzdKr8FXxcSpOvbw2F8Zn7fQp7/
25R3v6w57sG3g6mHfBsi579PcrNuJUWoZosL3bU7BbzU5jHMHBvxs1AmPljFYMnH
gSzyBEykqVmFQDVBGH2oHrKMzLEYx7f+M6PbUQHDtkckOqUvlFVSlmAT1dUejtSK
DIF7vBFeEUEOY27mGookj+xqkINEharPrUpWUDUjG72b8lK2Fle/Qw/cy9eWUnwT
r9q8fAx4QxBnwl+3df7HKtAhVGdL2EwVwK51oHVr8EjY+Q+fU+weAMjuaVb3xLnO
Ue7J67wQ3T3JXk3IY6uB3tz2WuCfSUzEZXMIDrCm+nxZMV86Yu+fdQ+svvSzRELv
tYusKSOnD8go6XrKkO4P35o6e3ylAdgHKYjutcOuqnC89bqaiqQQHeUGSftWjYh0
IwN5yDEdQBnxvY+cizwB9XI6EDUfoqIgeBrC6VbHKIV5gfkBG1RgvamUw3gKBBnw
HXyOSdVMkgRLKnCTqb78jwNSpheJzvE5zG9Dh7WRyGyRMMEjQZZJ6cu2x8YAX21r
iEhGZKgIT1q57eF1gCX1siVQkGVlQdzomAVTGG3jDWL7FYfw78u7Yf+FXPE8789D
+ZpHg9ANl0lqf1b3RicV9rY7I2TE82DGeu6I1z+gxKScUk/Zka2AKE6pTJGOvljz
C+AFHZBRK8V+WRQ8wvm/OHlW2GJP1UO2PnwpNP0h75ZXBHqNKBC3gC0w4qtUaCUh
flJkMTZ5DZuveH4ocLSLY6zPJLSFKUlc8WC7NHtFWjWaIT4uyr0aukTU2TAbez/d
FfhZhcmINEY9YQWaHHCHbGrLU5S7QZX1WkvggfJR45Thmi6nhBnB9mg36ev/+4Cc
2GeQfgwv0eyfOridTCl0yNXjGFk6dZnkbeuXeSqcqqLzDodsQCmAn6zx0TrQfhfW
9DOM138wDydxg2TEpVpfMfMDMhwq9GqQIdEbXWmTfLXmIP0a9RD+OYqlIP0YQEMn
pvH0+cM5k3pXJp2w8GkNAa/LLBb0YnF42vOSFA0PJVHPJlbDqBEMy/zeTsrhuCk6
HYRBuKVeHppI0bKx+edU+K5bYL+gcf4OA7p2jzEnVhHPQzpDZBOXNrONzWOofuUn
f6ODJq0hoUjWBO8IH5J705GFEwpnmTKZ9AenCrvTNAf0dpqU8wgaMx/13/EHUtG9
wTLxQdjT7o9HPxWEJvIIDrTST17H6wbK53qMx7OYcbBJlf5w+T/oWGRQTZ0mbkgM
1uKEm5mJckCK55wmzKtsFsds6MEfhqksgikkYW9uaDlmQn3vvPk2p1EFbDaad6jY
4vaDPBySzpC5soJv8cqTxD6cocyKVPvhwJd8oDBsuligM/Xr0wmeUbqV6OB6oZqJ
NVu8NLm0WsKnWSVQxXXaM+rnQZ449czbi/zeOtcHbWZeLBDcrAuOtFZUxPbYvdIr
K2QqabzyjbkimPphF5bEK3HUZwUmtPouVpf2W3kd6sckQIuQcztrjl/9xpFb4Vx8
7Z48EqmfYZQnXaSxpSqPY20gpiz/QX/TLSV4GchzlRMVfxJD63IO/w6OGDlTKTPi
KOh/6Cu14XwJZcl3pTjVoMBp1uzV/0ZFTrREvFkqZhhHpdMq3fJNo6pvNDRwjw2q
kgKhQIJYuvuVLsjsnKRTGgsiqPeRL0TUpd2KQzRh23dZQf8GZeDJxSvAdpnm2ZIn
9sSnZV0cEXfc9Nq6leVI+DXTjlzKEHCGdT7EX+W8o/PHi4uKm/KfOiQbR/45FJ91
Vu0qzuo88Q9Pl0jZjoFpZ5SmJMpGxmsLXBmv/dxGGKvfX92pNSjaI9+XtM9abiSD
SGdM8HDvMxcWDr/jPIieyxew6TkfCZ0mxx1pxicnzmO7w/ArYpOqYElfuS/Ka4K3
Wsd0wQlf9ynXo2GlyZoqoFswPG2y4xJ73k6CkC16g5FT1XDX9kGfalIAo6vKvGWY
jBy1pEggrEdLg433B3duT/oUXNziD+lFcqeTyTF91zbtXgrLBlYVLxiAbkeYAYAx
fuDLsfRCEGFJoThpsZwbhXJ4shVwGEshMlGpW/yUhRbf8pFEtt2WRA1YM9/Gz++B
Lnd3OH7pKni1sRTDkJQMWHxBPbNQUlocdHVdvqfNL0RiJgPHoErAiBcZP1/j3s5M
mC+VEnqGQZ+ihevGCkHnxtLlDe2/2Lr/yRDEpDgd7ybaws5Tcyh4GywC3ZeZRmyJ
mmipXBvrbIrY0sv7M4oKlBmUiFu3vobGibRaBCwO73jPwTvdMxF3OPdz2myq+HyS
NIXEmpvEdj868QVpW+GHaCkmBLA5YLKc1vAO3ZnZlBh/W9N/6hJktPBjBEM/0TZj
03zRhPsIqzvHX7VJUSO0EEoZkBd6/aujLMVvke3K+W/pvTpdSlBkEW/K3SydnBzB
vUHOCtUhFfzAKwQ0EhlTKnLrTvO861C79hXzEnqLfKXAYEtPHw/f5Bf5lT1FtJ21
sNdtIwO8avL8Siz5f4IfKkXPH+ACJyBnVwwMP3+82WOiSYcby8oSeL0yuYldHSAI
sHKSlUNO25bxXbaBjmZVW75ay1MGf5nVhMC+g0PQI3UemNA6uC0cGfV8Xf5xf+cl
KdqBFZ5i3I0krIsdOKsoJ8s6w5/0StHZsYyXVJIpHmvRJLa/QPGhT0b88yPVgWpi
1j1ti+oJvmxs/uz1njxssyyF5CiyPnTUhPkFSHoACtUuIIYoDGvJzqT/q39lW/vl
xL62W4dINbNCCFvifauLQUADpMWEDCOw+bvdaPXaidxPbWWTQplw1CvU9ZGtzylY
n/wmttfhiFeKozQ3KI1nJx6l67+CnsrAG9T9mOBOq9xyJOSQ27ROZWIwGcOmTmtn
eV5mafff+eOWFzAH+0rDFWWbCfioOOOskS/ZKHoS7QPcsHlalXsywjpDDF4LjJ5p
xbRgy/iuqU3qkavuUS0bw2CyRun4nfVjmB5NyRY8GseaKVsNP4yAg4Ll8GlHL/jj
WCJZSkdMS4/kpVszJoQ1KZpn0fJrQQ581j5MyXt1vcPwQQA0IMemEBowM1GTocs1
2MyNHTZ7N79wyzlqRssCw6LsxnlWbzVdQRhaOBxMkThW1Us+V0xZ5cM+8+90NSHq
2+zBBoM/s7V8gTm/iSqKifpjm5YDBvAF9ThM0dHuIe5PdFk0+NSDtIbtx6tdpIlW
zCjUKO3ybrcVVHooRpWvhiUBJTEA1XFXw+iSHmyfTRgtxP+GVyjbwatRibR0In2x
StL86hllJZ0la7iCKYrwIb54bZfIaYnfc3qQUqjZk+Vf73RHGGr3QWUd3WsR9Kbz
6zWBR3rL5iIUxVYHF+RImwHugEyhHWwGmjM8bbTVQWJPeawCwQZl7o3YG/Dhe2AL
q4IPy6v09lm0oz4rntAPdbnuL18xebGUD7mKmdd3ojAaSBs5Tf79mgOkSBIoO2eP
jwyv6+eRqw4yo8/A6+RP6lsvlEZlg+jpnSbg8pykrhvoAUDD60u3SyAbYPue+a2l
28vnGg5wVKhysrj6t+WkCmgSnIAbpQfzBqJf20s8Go4wqFpHPyD6WuGi8ACt9B2X
eiFX2ukjOSm/un+pesAR5cqI2gBGDgY5p2wUHa8HGFPqCJi7qAyrKd9a6CRqqPe9
VRx9cyINRJ3UlpN1IXERr3NOwFpGO/42WzewvXGOcp3S2vYYZuO+JkY3ItFZ9SD0
FTCHIOKyTXrzjjSYCKQ8MQYSLWyD1oh9vTMGF3lAUCuTbBT5uRCIR+OK8wGOdROZ
l8Nb4bhE7FdZdegu15/v1QMO5ekftSHPbUU2/r1Q7zxxKwRtWY4xX0AowRtnlx9k
sm55hUATIPsk9kfAQ2ZUBaTkjBRaCx8GW3j8fboyif5OrOqd2/5Wgad59sg5tal+
UNLxbn7c3PkrLH+CIMsHYKVLJqCVfeYK6wa7zpTO+s+Su5Dt+UoCsuEDR7fnlO+4
PVq2Z4GvavDdR7gLR3NS948M0J13S9ZaBrEmdA28sl/BnaewdtPKmVXAIcVFs6FP
FpbmBuj63/ORUF0KqBTNb8VYVgB3jlaoHsOuMTG5wNPKBOf5Ay3jdMTMdWebtHtd
+1fkF8ZSoxQthb6ibAOmyJHSYSXntn4zgEfE7AoZv14w2QOHbFsFpu6CfixC02n9
peSkJTMujSfgphWBUKsPUqWOCdTJUh0P8wb2zmPeGWKgQb2ZG4/jvhNwxVaSDWBp
yUnZT+q/8C6GKb6wPmoAZ3ychCVeBSnuE470rjsOMxbCspkdX1WB48ECw7xODOxw
oW80GR5EW7p9l3rJJwKY/2MkY00wGB0svlgv0MaKqN6eEIIYSfo7XngVv/Poqby+
ft+Mfd2Kpn6L17RNuLmH/IuUQ/6FIoc1u/Axd+qZfFuACFu+QPWgrXZZAWkcW5na
//j1uagrqqOExHcmCp4CdsLsWttil+FDW98wbTq198Bilygx4uQtpYr2li088rV+
9+cl12wz+utLNCsDyyAUmiKddUVrvKAS/dRNgxF+j+5E/GsKQpuizovFWNfKX7rI
VKosT1weq4zK8T8ibt2StkHlEV6SD/XrSZ+EB3V/r2oLOzX+FiJr0g9DfmOHMxQO
D5pCZextGR4xwJ+FSbs5AZ48RyTtoHfK6x3fJRcXC2oU6apeLSYx6idrv8ae7foQ
DUaTDmyZXnYf+s82Efy5rGf3Qmkyg/CkjGDHLuDUtN0LD9ffCgdM+vZtGGIhdM28
6fpHrCHxqMRTQduZAf/R2r6q+FfSpaf41Xa3bW0bzLeD/IUpmJ1kKdh4qulpgFYD
GKK2Pkj2meWLSPmFPW3HC4FlIhCz0sa/6VJsyWRif6UJZaF2hz6RnEuKAVxK9jK0
U/OND6xATZWuwq+74bhBqq6Z5am3hITIm5hHZ9lPpxZOtbtCypfsJmtdxMzoQinO
nxCQ3/cSkXPzRTcVfKAMwF2njzKD82KeG0qwQDZOfcwsFeHEeh8+V+E2lm7Hco9E
Xcs+wtRGV+UgIHMFKGal2sZfce/NXsBkfwXqa2zBZi5iEA6iVUw8hcrvwMx6Pe8V
Gdkkps/gi8vBwEd0zk6mYlYSHaA7cJlZGa8Gom5rDsOLeQfqydpbrYrEsP0k3dHY
rQn/sMiJOH1YQ2eCmS2LjeReMDDZgtKdYtIdkhCPAqCNEsuY8AgYlyGpk2Xkw1Q0
jlp3hzyUa4KQLIbjqHy79KZzzctKHszxls8SDou5Ib5s1SMotnMvLfUenTvmh5Zr
VA1ssVnr6DLKBoowA2RAE6J5HAmwkgCOMiUR4JtgDXLze/3hymt4j1uG/puJWNV9
3L3rdjJUP13MPg77w205aKWchRvu8vDFOGnXWTmquUZPBPlFJRYpSfujQbHtLBR3
NwP8czWeEj7kLQW8rJ+QukVZxVklMgc+Rqty9ulJ91/cAoZMh/Mu8YnO/cAmdJ0Y
FDccvqAQ8IeCM7tHRE2sCc+yPXf7SmyiC5GRyOktitC7ovREgwwoJGBHdQkPDBHr
kj+6n3PFTa9TfVxczqkIonlp20UTRSWPlOonTa2xRXKuMesGxqifeWqWQKbPgoW7
IMRT6orLSeRRj7SbrKgtsal3JN8IuO7R/M1BEiDKboZALuCxeTYV0si11F2jf5q7
jgjWOHEZRdycOBIo07TujAZqHtHtfZ3rKX0FHGlR8ZfJnKPL+x5rB22M/0bqn0UP
QawoG5ZUq9wdpeog8Tkxkwtao7DdR2RDNFCZ/tZv7j9/qSyw0mzRfCM7nY/pUyq2
dTHyFO3tYkqgqgyVPj+mKEcAdc2WbvVmuQdrE82W50AUzR4oA5fXQIoWkLj9YDe9
LumVHX4rALmpzADShzIijhcMAqa+JWlg4i8INgTvDpsZ61In54+VzYyQ6pACnXvY
32y5JkXm9dTCHq6WWU7Og39kMbu56q5iP8qR9ly+DBqETry2cW8NPXhpCW3oqy2R
nhVsMEgQy/Q4anK1jjDfwZtZ0NMYI2X4Pa1Vfr/lMlJMn3dBlM8PCZdZdENL6jUj
TatBwbafizP3I3SCUbvuGGcJokvz1Q2URXrBG8uEA6uZjgE2hAF3vbq08HH3rtut
QmbCKJCJU71kw/qzFsOeRg7MR3znOsiq1H2GBzxVIMvUlL4+hpJl9njNFDeTzzdH
J6R+Ms8nDZaHx8HxHXSY/VAlc/DYurdg5nUFErav/QEP9qsHs+THEeJs8oCrPz0m
E20u423yFmzFPUajO+zCRa+z/hpMaC4uD2KIL8gD4HQ005lxOapLAZLWt9uAiMNk
rFdgiGJs27l/0gS8spwmwlQD5e+BV0SEChVrppufK/TZ2jX2O85lBD6f2/d+X+yY
rdbhhiyF3kDBLpis9Jry1JxjOCmTxGNvmRWy5bXLZG7OXGuoxpotsplkrWTYPdJH
ynP6WY3EFvyMUAmD8qXfooTAdpxvR99MZouOQGjU60IfkOxUaRqIhaTb19aX9Fzf
tm+OQB0mfaWNlGCjNvOhvRb/BHyHkuxgzPkmNAN+7IMz35DofQwdBPoF/P8JkggG
N2O7QTFJcnXt1nXO+9NNb5AIJtK3xzp9hWCME+JIC7UPVu/3P6fi97aMlTQ7pxdx
3d5K7Lp1eJ+J+ve6altIJazAnxOma+vLj7eJxd7MBHZDz2t8HXnBp1mCqJYsrsPy
XhnfASfhDOyl4H5zkd5Fnzah4BOxLejADz6LBx6yt/wvbm1olJUcROQ5oFAmf7Af
vw+tyONqwHe0i3Vo88RIkAz2op6GJlvwVXOqssFCciqxh+AivFP6ZwnlEYacl9Qf
o6P8ityD5MZsQ0UDLWQY6UigJqRQZQTyqfMqr2pdRniRe0RcOXJNSFU83xe0uuCc
5P3edNnHtXOKo9S4KyljGq9wYwY1Xxf1VzUfzYFatmko1Z/7GVgosX94Dv2Kp1db
RN0ci4LAPHlM0a4fCCzZqkbo1AVvx3KEMpgcN1LN5gRc8ca4EIWUKZNNsO3LWSuG
8Rns+87y/2F5JGHv78KZuJHaB+QYQzOWJuv6pZlctNUMTXzOlCyxhxAKFEYCY3lp
22DviB4/KToGAPI2Yq1H/L28ZOrzZ+rep6tNh3tsXeKQpFXz+F3V1xjRfIjsTWIk
rq++KCxKQa79yhOQo94rAiMzujWTi3j3Z61Pczq6CaPxws/rCokFQWksoipkUFF6
dEyQo5hSKSZmIKBtkC3e7cSCh3B0tWhhphrIcydLrE08i01kH24EeGjGhKDrP4sZ
0HneqmzAqNnM/T8u9Ir5DOQBQxobsxyUrxoPsvoSo76NPfQ66zJ1/0kdUtfhby/e
tNsY4RTTdfSeWZQx+F5FcaKTTtvueh1qRs14ljUX/njGdc4COGvUpDfAZs2/cuwv
q1TP9tvyDz/OhVnN4+XGf566JZafKuYQwAO2bK7z2j1h9eceRwiuBJ1C/tUQrHVv
+6rnaBUzuiK+qnRkgaLePG+0s6IhFdQk2LacFKH5xFqzSf7W1rUWiQt+4v4B5Ayj
kDchwaU4vB0xjqdln6919/JYz5tSo4qjnKhZwLNQx0pFhQrx6/SudfgUStojZhc6
G+pT0cUapWTmuXUpPFBJ/9Nfj5Tq+rxd5r20xyYrFPJK1+e3cX0Czclfoxgux7/g
OQPN9SgMgw9cyUs65JmE6SZ8IEa5hfYgyqCTWtgmy4ucPJ/QlyprVDLTzjAp80tn
ZWb/vLU9jaKhLVfqs+DlrfWW+QSB4gzJ1wcjKShZOtUw4/4tLkF1rnBqsDvOP0BR
0CIJdc71TQdrt7LI77JszmDupWOqNYJe92puZQWu5LdY0RBdncEg8lrFW0OqPxKY
9o91vOFYn+BGlZS9UwloGHbN88NW5azZQbYJJGnv1is25Q19zyMtYouXP1Ocii4D
a8i6YbrPjaEjpAc7C/DVi2z2ORqcsvs324ZfdCzrPZsTzvoO3wc3npYvX8T1O3pt
p/fVGP0/jstSCmlURbc7ZSzEU02Cw4NjRp2iaiALgn8+0RmhT6HOSWrKUz0oInWn
qLw1grSpNzXvB73HmTURlvqfgw2vNl23I/9O4buG3B0qs2hF3GWCeuF8ce+PdbsP
pWcTKwp1HV6Lw2Pcep/ZySDNBAw8Y1Z8qn2B2aLCsNN6h65ht40viXbNzkNxh5IN
R/Jm7ApHxoOy2BV9ZAuiHFlJY3qdbHMaloxhnYqAOy+NzRjYzjwXvUnwHxam+SWU
tPZr56n4cvwiqFNof8vp7q4+xgcQw9Am2iCkEglTeoWmOg1Az0f11jwifruUPsla
Neg8POXye56ybxnpJ2mAy7V+sGw1Zq/+ECU+KJQMPv50De/xGnuaxyY1zNaUbjTw
m6gHWjyASW96NnV/8dNPLLUtQMKkTWHsCzBjfY1LYeuwh3iZFvnsEr2Z6eQKvR3j
uv2GyxyhdXtywtneVdHrDCtaWDtMd5VBfRgaX8R+z/ikyfib1L5zvmAVqR0sb1gF
HvBsO1NE7NOyzYPhbLk6kXeayZFbeA3MTuswyn1lNSkgaq/0tPZUwyblNGavwnUI
vhuRdP2pRgrRlnu3lwd5mvQ+xiprwG73ZKmdxTnJPwdprMP2F71PvgjYrUBVYScl
PMhMIj8MG140jc+mX5cUz+HQK1kTtw5iIHZ+u7FM8ugpm7SFyDHR+sBqGaQlzlS0
PRNKbkuGLvwiMQpXi30mDTgmVNdJOCYz9IVTZrD+TMTHRypNhqp/+G/qArIu6+fA
3X/7faD8hic7ptPqNifECHGoU7ELioDCG1bRy1QFBkXm1lkdy+SM4wgE2RGCloxf
rer2/LHcXqS4KMww5Ib+UGhIOJpStzScJ6OsrGJGSmc1YCsuzJG4M56tHlqzTLxu
9CiO8ztCfYFOzTpIeAHH+F/hOGy7YLz+aKQJ4DqVAqdcgJrwIfQMsDtyEr1I+rtu
1afjzfddjd7TfEEQRveF1OlIL6RY0xUwhLhds9tuo27KcfYsWc+NzD9ez3UMrQOB
D75UF/8dAL+eXkqURpi17YtHHJPT834MxXbDra973k8IrsXAcjY9+lC5xf3dnSyA
pz5HGwAjJ84JKt7wICZu7p0iWQfIbe2IwVlOAPlM7bTIQ3n2mmS1hB1ev9vJUQ8W
yG+G+ndvegEFo/wAjrHQ94/SxkS0BCChY2YFfdQADJxu/87Il0chla+ii5hSMR0y
52KIotNoXAZymQr01rCmMsfYMCkGTUs5MZmud6V3JnjpXuwqAFeZxobHi6EOxZ5G
56m/W78h4FFtE/S8O19dEFhtborCoW7qKTUN9Qx2Ou0QV8WHJAia97HjO5P4d3j7
R9tEH64OsKi5v8eDHIJJWJGFo73l5b3ipstcLYHkxjIZ+crvlAja9xhpqSCT2Z/D
ABLPwdsizYabuv6ZJtqs/shcQPQrFrP9ztLjSRAJvuR21bG52rXlxup1QibFr+jy
UDG8NteHM+Urj/hAtqfViBcVRKgKhc6bajR/Emc0MPL/uJKSYzLJxKX3RcTtP3Z6
3STz5tCDTPCuF0IjDOopa6KUC0KXHdEV6uxnUb9HhC5X1eF9TyfauODZoDGRvRkP
ING8zg2DUr5dCYu+WgU1pQ/RzriWHoe+NP0IrU/xaNhv9bcGwUKFMt+YQAA4bvEV
XJBi35Tg5UA5Onaz1zYzmfTgGGmholygbR4eriNqeJ786n2qOhsKmzXM7L1hkCD+
47/+P1sSb332JxULC+8z8LAivpCk1S370djfOXYZrYE7vVmfsf2zH+38CsC4UaSV
NHHkK7tRos7ldL50DpBPsJJWNuYJyEdZ5QfvWfRG6d9b+0hEtoU+amTz6X9ZcrqE
VfUGBljEnF4JplkgA8rdb1pNjgHAJ3Nm1Wy0XWthVZcrXJHKOcmOHoA7kXV65iSx
bGbQU0C96TGMcP03bpiDnJ7LLvvqaR7Jmo1nY0mKcDC9QTGDkyTqfKMGO11x9ZFk
r3z5/uE55I3wmbkpg8WxiZJkLCbbB2pP4M1AJTIQ5XOoOFw5Ds/wH2Qqws/jPu/o
VbzLTMRxXdGGl8QtYy838pgpoVFB7+5XR50fkuJ0fU0wFGbNpacvaGpUfxxvToom
t9WmC775Oq2HBShf8RgSJhnhWju+h98Hv6MH/zb17oq1GwRil7jui3+YCithTXsq
RVMbYmG0hqWIC5nE0YlY3bQlLIcPpIkZYp3RGsqHhpjrW39c4kZTybJ8G5LLbeMf
kgZqiPiMPYwB3++b814wY+sDH8ef8WRmEuX21ECVPMmaEDXxDTXY2spe+VkXAKM3
CHftNgNuDiHr2tQ80/nENtiK7n8qQ9GZhAG3IqMmo+OHKgwdT7g0V8BeqshbG/em
iGnTWJoh9OWtRgaJS9cQeFmg+BC9q7xbB5xA0QnvHbelWCNvgS10o2w4M+QF0Kkp
IC/cTUMDprWJqvpuvXcn0QCSzXfLZSq9kZ/gm7zcI3X6g/Jl//RI/bwlrqv66fY2
KbTI3ghJwdXyoQVqRZZCZ1LHpbYbu+2AwEDwJd7dnSuBaam8NgZre5pIJZsAJIil
eCIhnLWZvdxGkO7GCr8+t4OG3eTIZN38mANBdi3WL9rHZLgRH7QEMr3dtFmmP46F
D5WDpXFnIHFsOuJ/K9+sdixSwW5Q8om9bvE0oUqThElCqC5zc5/HeO4AsC0/4hsD
dykjmEKc4nj3hzdl2M6nHo2dtI2HapsVprdgVfVSDCw13eBv0ZHC6Aa8YT8tVZ0s
GceXm5/0+61hvuEVbtZpGD3Sls0ldHH0JupvCa7YhNyYcRmkdb/kvbdp/GWuMgd9
YDIO1r0kC28OicinYTRy6y8oaZJ5Sz4bMNZgLQy04XEmPY6dzxKHGjNnVXZEYKtw
V8zwcZcRKpygYmfYlwsB9bRBkBfBj3oPQ2T14EezrTYm83/7Cze3P8qTF9dfD7Bu
f4SQUeQ4jSKOh22vtI3l90Heg1frfnY2eXjPw0PuQVFtKfPvC0pkim2sT9xAZpWN
Q8b6JfH6tgceDgqsUGpTwZ7uwWLX93ITyTEo0zEkWhV0ozeVX3hYFffHzsrLdpkm
hvN506y7KpseYl6ZarRl7GUUhyieOZPCsLsv4Jw+kXIBDnnjVjUPFyQtj7ISh7C0
9u0hGUaqPDZkWIM+eRnoEKZS3pnyeqq5mpz2azs+anozbnB8pIDaJfWZ885L4tng
7HTPcbrxNB7y+9nDMUwSnktiZ4Knd5cr091F+5MZVn6GcNQA15xOLXgZE0apexDn
kghoOcCvkbONe8AQANczEZofOWXHr9f+j2FhpKx1tybkrI8Qtz+OhWJDijzZVzS+
Sl+5dtr4Olt8BLzoECo0enmA9v7rMo8JgKH9jay23J4zveWZyvzoCzAFdNR7WrgU
6bVYsu0lOpbTbTwLWOe9FBwx2mzH1ICmvN1Qqa+glyZTI4Dg/A0rDZqf/9fd6JJx
pwpu+Jx51rdy6YOg/Bq8Ch6U2BeKGhjlYw1X1BMy+yORL5x2AT4LXY0X99NRF49c
fHS47TZDzwJtzxHew93KgKh8ah1TY0OVeWLFV2+Fkj7C1boaoGPO/NDr8DAPk1eY
+rXHw1Kf14F5G2n8gToR8kClFXk6fwC+nwPGeZfvT8OxKcGerS6ybm/O/YLnORTB
lJUD1INpBYtG72+GPAPdP77+MyfXCC85inxH3LmuxSxxhNWygPUL56ocVTOP9uHZ
+JyPK5fbybhHeKmfg5vtJZmZTUQaE0zYO/jifToBiZHpBpXIuPfubvZgLIYPx5Z6
/lQQ2G13HM4EG/kyp+gLePGV8rvkYMR61QkoKBJhvCRaejQty3URtsYKoZZW+6ms
WzMQqiXIsi00v9zhn3+i2HnV8+IZ76yT/MgYsG9W+2eJlm9OCf+p+7iwPKmZQE19
K6q5YiVeR8yBkASYx3rMZAoHPadA2UhReZjpv0oibTPaXxueuEu8yvOuczJ+isYj
y97nIGNKaAFkWy9NpwX0Rkyo2x8um/pTzieLDUaQWu7vBJxA8TIpOfexPR5/bShI
oGrBlgIZPy5/c14xJ1V6u/dL9JuEWKJlmvSKqJGqozSClLCl5gM9K1d4YhA79+Fp
1sph5lBQ1j+EIDRYLUVBkc6civzQVtrTC+T+EMgxcgJ08uN1e0Z67DOJ2UyaMIe0
35ZiB4dYfyvz3V6fT4EsHE7vdkg8PyIg2hxUchKaOQmJ6EsHqGIumB3+xNN12rVb
BM+Dx1admZNYGdamFVwoQ2kYPlkEUQujAXMlUiOOJQ5wysOD7ueUSUzrsYdxGzT4
kDsWVu2dyNzbYbfBCccASplnKvHxR+SXNVyYHmkRhGKgBtvgVCVSsk77YtcCeWxd
xHh9c+EZw6TTKn0b1LTXxTTxvFcpHh+9hSjcrVYqAi6TuYpBF5ajOHQ2is8bIfGE
+hvG/mZK0n+dIStl/VXtmi2pB3Y43OK2GKCnYYYItXs0gWOyU+ukd9E/POtzlvpV
sGiVNh5sFX6j9K/AabbqcIGmZioujTJNgya8u+glDkXnHpeahy3Wn/1PeWlCTTNA
gKhrNb19MygdTcM5b3uWwQ+ePqSbnWwGFtE0KD7C6JaXteSciUt6hPWWGGhxt3f5
RtHmRHQLT3Aeq9gIg3nNC2IwNnIkLrXpMDy2gKavw6rFtSOeRWouy3aCclm3ycBZ
skJw/peheoZmPwkf8kAKal1uuFP+uULslgCsBhchsM/a7SYzWu6Wf4Bn4tX3N8mp
a/omzviLej7YYcYvhWKySuH1rk1uCE6SWO0pbiJiJChuLnCBjdDTav88xKX0e7hE
0lFKdK4paXRcr77ecaOAGWFfbFQY9T64Dh0smhyp3YaF0NTolBQzseohbDLLNceh
NfFUHzPcHzv4KERjRid5ooZmZSzLGEeTRRwsbKNacqPgF3qwbFA9HPB2NYM1GFuH
xVu9AfQTuhKvYWBrGKvBxuiAIBsGMVshsCij4FzUnmqw0aFFx+mNNz+IG8D9DdQq
EAb+jWmoBQzQ/R/Vz7Y+A9l46te0AwzsUYAfTuSrGksxqbzQQXwIlPD/u00KBxSS
QbfJXYoXXYwsD+K0JRpl3Vj3ZP5fO0evZr3wqduBG6HESJkjSvc4tKuiRhgAV+SE
g2Miqj4ECIZGLnVKSjquKyrcNIm260TGdM505k/rZt5jqX1+TNgNoIhhCuPpKYmc
bVEkxnaTq5yBo6coJgEG+LgGybQHkcoLLnh1yFGx5/r+unHlubScTMdpQ0717YCA
Y2W1A3IJOTcMvkqlKjq+/01ke4Zsh2bZwu2OBifud9wJD2UTTc1mKvEZK7A9INRJ
Vk8L11r0QbjJQDWYwFPedplPnpVUehqoc+Njtge5ul4dP4yZpeu3M35xUmWW4Wmm
6jJ2htlVvtWe2ECYwDaw6pBavfgVwdVMQcA8Z88uQcQPG7JklaoZ0veR2rbYW9u1
cVi5l/ER9DTexFKCdeoMbHHTUxbwGkoGbZOqFbme9BrcwQOIEzh6iRmgpxyDIkLE
S+CVaASnFQYHmf1wjrgfMEEQEfEOYDkBiC0J7NtvYiRhddtKIpY9mEQ+h4MMuTGC
3t1iYQSa51HO5FvrsJzx55Z6sdaaMtxtdWODj/77H0t6zSjyPS96/jzPdIVphqPm
BSYbHJ28bhJaSTB1kJrHQrnBfmHfGNG1BJr6hNZGAXxB8XX+Sj80lLUjvZjSiSP+
iX4U3xImYNmyHT9Xkuco1U9qEbpy3XUZ0OjVNNOlIsP+b2/F7ESoeQesUEOAcoHC
f/5tI+LCpTehU31Jjc9YMcvXTLFZ+i3Q3rtwM5VDLKvtShzreEw2lwdQymtszHxH
Zm0enq25oqPt/zGwqhkcGPC7qSWuyEOp849cRaAm+e09ZSmEiy9cy6PrlMr0bsDc
/w/s7erUGVO7TYOAoN6CwggVgWCLF8X/3ibyOSfX25eKQmjuX64yM1exasdkQaC0
qZaVvCJs13ybJtzrdP4cW+3iifWAIufb3m0138CKYyrdbhKDjsjDLNppNqiK9DZx
yit6SPF6458QKqPYcUGjW9Nr5nLQC1wST88BpyUx3Ind01VRLf3wWPQIePRSxi1O
COj4LGf8mdpUrEgpSUNHQ9hnR1kMrZIxKh2i1W5gzLAM6fzqtWXnxHa5k8jLJJWP
T0l4FFQZ5zfRsDbkBhhMK2fJZkRZZScodFh5s8DQLETw/j0ubUqTx1Ui/7CREj8x
ksxKa+tESvMInCjkzI1DRJ4XJnRZzsMMNWkWGccVDvmpkN0OHuAACCCmmrbzsF32
aF44PeBcQJ0OMQcO4gVLWbfRQZNEJ3ZPErAWHtyGtBiImIy7SfHWpeqwrc1FxMr1
Tn0eGV4NwyeufW7Ca6azCtfdypaVRpHZqHVYEIMgMu55SyHg7IsyDi+P3JDOqtAu
WGosegtncCrD2eVvP9j0nGb4E07V+t8TCQIzpWZWyTlgNtInnEsv0B8IWATJ8d7h
8Ltm3BWlO0rzJ1EhtsNbMpPRMB3c2FCbdDEj5ddZicC9NWuwvL9nU2SBG3uihy/O
tzzrJ/VsP934K8xDgsxcEKLmOFEuDTUe8o9d6h/bt+jseoYHL+FUoT3E98b7U8ok
4ugRCA4liGTHPvu6/06Q/LoM9WljTbvauUcxklCq8/neWR0Aq/uLzkXs7pPDduPn
hcaoIsN5QbtAUFBeWWU9lNE8Futf1pASl2H2NUF6n0qAuwsawstxPrWaVEKAKSDg
6W/TH9xT8a0/Sk5szDKLTktRP8GX/D4HFqxc3NTc9mQ3PMaPpqb8xggVLbfn111g
DQMRLAiI+JboI6NbsGNa4EE2RgN6PCUjjHobVXz8ylS5SpJS6M1ivj+xPdShacOB
2aCdQzAmBGanMugRp7lydmoiqkT58O2d6v1m52W1W5+VXE/DFhOtxigE6iumHDGw
AfspIrlUoD1V6/2ZZ3mIur0bSGudSJdzqlf//w5bT53F1nH7gagIaPkcJHtW3zRS
kt7Rh9Bmms9WQbWIHu/zbI+9ukDWYgZNh1SgjTbjjWmzvOAHCekvn4BeP/OPaE84
I4hwFxbYQgvvQ9K0ZYUa+g23w1hmh/mAN3hmvJ8ao20tk3mfnNn26kAoWdKejAKH
+5p7C9d4xLCRAKNRXBvHQs9AM0QzKyOiY37wr9EKzFlkybytNE6xGyD3kgb0rdu2
sEUJbPCA+8SZ1Kq+uOriB6dUOc72VJIBpI8/t73Yu8Un6fcoq6NtNVPgjW+iSUSc
mQcCJRp277kRf6LZmf1txySIM3tso8i9wpTEwJ25GovYde3rc1MGCXd4z4ox1r03
PjrpYcb0791ROTmVOpKwVu5CkR6yaAHeMZ8otgzMDx+jOs+VlcJZXM9GPdeaHBJB
WnCRY34txN0svF62M27kkIR1YwnNhPyXW28eOoH2L9zhKm+6w87Dt9NeAxKyK6Ep
TXql3Wc677vuXTZ5oIxIh9aulk9V27ix6V5Civ3HM7tz2Io0A1F+6rphSnQoHEIP
uuiawjUGz4kxoz6T22eN0n0nBSI78GtVUmokvAaREcn5347Nz1QZBuWUsX2UfCLN
WN5JeuSxQBlLc+E+OWUjgkT3zQ0oQw78V6/f8VI15zFXA8LYeeAiJBxnb0wzvco7
VTaTSE08Udx0E5DYb/9YKj9Z/NlTq+BUBkEM5QGiBDLXbfFcKicVuZw3yX13V94K
bKhQD1LBInVJrFVB58vcM5BNH3uFfAeypwZPGRNQOCYvx4FNvo5/5gsBKr5h4Ize
dwjqstMneETyNT+hqGkmAyJ8Y5lnVBnrgq5bjgAncevQAMVN3gUrrOKT6+PAgFme
bynae/ZecY603CYws8RPOzmDP46ZrkTiFaewzeqFhTDGNZ7m+HXZsC/eay7nRlhE
u+fUGKv+o82LcBYuz53VUtVoWOON/NeKVnTFKL3mMtu5HJ0j2NPR6erq6r8V8y8K
jQRWNLwUVJB1jCB74Sy+iRaQ5u8DycFaLSBUHas6Z61tGG18h2oxCw2FUyzsJkpL
WRt3IHky289eBxpVB9zxKg7pYyDAa2CDSY2K+ljRyoadknir59H6Ht62ckO4LEzX
dNyHqUJqsy1Wteq9Jrck08EhH/YPVLXSO6D01N/xW9vtrAf7hox/Ackl2U27WfRw
nlpL6+WRkzKk7dAKuoeEkY9Jky+lbAfJQQpOsVlar8S5te1M7WAUfbGdxl+BgjKG
MLUUwE6sGCRaVs0kDXZueres8U6Y+d1wD9rjcKZkXDAArb+Fm7GgFjyxWo1u7aXq
s/fLlps8LEyB2iv18Q00xwUBXDmgq9enkIx7ozodmsU2Ah3AfFzNRNbPppf3AakK
l31xyq1ZJ06WwpvFLCqjJMvUDJ4CSl1oUqEJqIyIZ9CQ1IW294jAbbChp+dmli7I
Jc1Xu0QCQ42XfF7qP9dYvVRER+hJ1M3VZTe//8Ma+Hvc8+gcmGiJuv1PVhbM8+hW
auPfrlzejI42EphWiacAMhOWfiiKDumiTZH4Q2/TtwuG+D9x0qP7Vv2O4ewOOkqv
SVMb52/4edxH1Bd6RerPbwFX5f2dxeOsvHKILfs/xQcl37g88QtfLPnzQtuJYflt
kHA9NDHQ5FKu9d8jJ248ijbkLSxPKAdkOFpe4hoMiYrI8FmT77M5TliJyJKbrHG3
GPGmx7ERNijz9teA5pBp9cZowt8Ww8cCZEoLPAmH15A1jRFAdr0RLqEucYnHIhw/
ol18n1+N3jl4aIQOqtWU4v9XKD4ccNlWni8J6TBiHvIBt4Z6458IJwnA0wu2OGSr
tvAZoziVTLVo6s9OtJBSPubybU/GcEPop9RSPTTFn5dB/2NvozG2BRBzvhJOajMP
KMPNYIJ5ATpSFKu1ZfJyJYqQM7rKwVfcvfN+fuu04/9E5Gb6NpEmhBd5xf4F9z6T
4Rldh8/oXqZcySlNG2UVx9CLyRQDkaMvwJqvV/9fMd/DzR3NeRiWndyzwxNPE50+
3gQxg3fu/4IQ6oPlboVzSLGuF1D0sws1EkeT+yj1i7mOBVWAn/TKG8ssuB3uig7B
eH0qq4ufMWN/P+b/47a2MpRBlJMFPZIUvZ/v6CY3Gli1qE5pRt37TCnCBm3fcDsZ
f0reKRUuOq3X/tI/7GNHRePB6/In+clo2Y2PsHSusB+Y2AQeQc7eI6hsGXQSIjva
aat3aJUqpp0ymBM+dE37UK1H8MG0AJPlsG3lHDavRR2oYBGd+UzCvRFLbmuQaBdc
xokP745ENhHyBwt0Z7+SarrytkFYWP5BsJqEPRICNIR52LNaSlp06+m6+PgOafov
hx+Ve3/udfvE4O5OqCpxLjoEKIyABfEOGIrJeVMSNrz/muVoGiMFQw2p9fgvsOlt
5gIoY000RMpC3uwEv392I+8GRFQIPwm5wxrAScaz4Wb3hx5N9Mms2hnZig3WrFo1
h1MCswRzW1u2S8KIpMCKdd9Iou2dOlKwI8iDYXmmHskKkFnMKHGjZs6H8W4ey9ir
dyJWZbkZ5eN6vhGZHONK5TuGCCkDBuWHkAUFdPHEpxWYSlSfInvdCEmZh+nyer9E
7blcQlPuwpGMTLjkIwz3lkcjdZEKbeEGiLSl4/WLv/MV1CxygM6f1eLoHh/wW34N
hcj8naOd0a0n6X4QA8TZxAWKl+8k8FKgxjZxVzuMwAy9VUDQH/RPPFD0w7i9VpwQ
h8vatlImGeuZUGWEqrXHThYqupqUKP5lCAQPKXsttbu4DoSqbGHzNeo0NFZmorAI
D/j4JeHVwHp8HcOGqk+X+5SHIBcSg8PNcCn+Ouguw9hcMC8miR4Y3vhWSqNio08P
DE3UcQ549pHq6cZ0WHsKngvOKl62R/eGrMiMeHnm0eWkpt7PdqpGeqTwVoLr0EA/
i/0mqS9XyuKNT9JHMc8ajKJMP8Cre7PpRHOxrNNQgjGt2n5dinTrAVA6G4RllvQd
XpmbpXZGVbHb438LQJMp+0D/9pGLNozg/HdxXglDhfMUioYqNXRplWMBBZTfV009
TQR14G5eXPO5TBfEyFwGaU5Pr+W1iC1PHUOCY7qrdR9BLm+nAD4aOxZ08VN7eSrT
5dOI5nixecqcowKkscV9Sb/PWTSeMiUZexRz8dsVxd/L8oTds6pxQraJh5PApjH+
FsMHuIZ1tiCqne9jqv7S+EVAxaNZ+89idqIyNLKLx071YhNogo+uz5XXHWb9ZeJz
tXURkKsXR5UjB0VwxoAzPww0HliPNENWVcl1yF47yZJwt34jbtaR7n6xy9iO4ww/
uqM0PHzCVQwYYCwaIR9VWoDk27mEbYzGhnMd59MDSOTPuoNpxyXNVjAUydlYB35N
4A1gsR+3rXYbt62oQ91yE46l7JgnozhgjIwgnrNWQRulLdGe06SjxjO6TSoU7whc
Ml4et5/pboQbYzgdrVAV40sFyFWICtJksmyVLIj473TJvT/2CvE48XUeaS6l55WF
AN/NA8K2IoNjT4t3DTliHyvwEo6O7FA50zEXDM5ySljfS/WVNLkH/f1YMSAqSVW8
LZ22g3unqAmLjZj0yx6dQqsPOIKwGL6HoG0PeqkdgaoiDURTYoeOV2kYfxwXaHE6
E8Oc/pZddO8RhYncY5s478KGVgvP95XBIBzwj929Jczh6/oair/7p+LzQsjfpOS3
V2ZFkVHda7g66Pch5ZuYNOifok1Alt+3Wc3TorYR2n6io9ecNRajCWxz6FZ9UEU7
UeBa+r0W+6nwOiBRECvdShidfE/jaSfv4llQjIYm/EGstn/yKGird3q9ch6aAnQ7
3dBYmemKVplcHdWSNKgeaZ5iuRxe+qgb5f45rQ/HqmTeCz7z2rf4OKJQaaxETmqp
RopSOeyofW61wSaqOqnMLm1BWpnJTiMvOcuiKHwPyAOEjNXoHgwC8ik4b7O8qDxX
iJ25g05L3BtI9QUMJKUJ5XouYpxJvC6rVtmtRtwtJ6n5y8kElqeFcGUTkxPQtoXV
0zYUHQDcjbP3ccaWVomy4QrVOce+rEim/SyN+wdM2ySbFD5RWIbnnXNLPrnHgZvc
c5EtHmtEexpxxVs4zEyxHamKKp4yBymKKGf9T7p5GIB94alxakDY+ggdHEpFypJm
i3ozhr2Hhu00AjZpIG2QP4f/flfkAz1MZWm7HDWIk920PiDrBIdWN0kbASke43KX
QU7pM5KBVAd5xzHLMFBMbvsj9Npos69wHlYZfKKBARclc+t5XM+7okJtdY25QsvI
lXZPgcpLZ2z9ilkhQk5Tf72cbjbuCBO6GkYtdxKuTmpkk0roOzML0UvreeEi0oc4
5mkjipLCNnc7HHZ/eamWrs+FBFGmHCGGF3mWuj7wxp98nuZowL/OUENRzgxMjCPk
gw2Q8CoySpn3KYW+I19n1Yc4phqMQvwByyfWL1g0rtYHJ+DPdX4kT9H4nc42aYef
pjkiFcFjyvgr4WZnml7xjpDgW69sMKhJLOK4cXMeTu+5/OWKg5FA5lr7w3PhXp9q
o4DCvwiwq3DP+Ehs/a0cCZd/o1gy2zsi7VYZ/7olTmU/lVW9bXQwmWuEMbcXkFiM
r2zJCyJCsY124A2ZgnBQxG7eqsphNPXLhBHqmnb8OO6f15xQI33BrgPqyYxSRL1M
qbzqQNpptrxqvVPLn53i2YTzN/b+v+NurhkX5Z5nukDR6OZ8A/NNCzYou7VLqDL4
iSbk0EroamNUOFFuAv4jhp1os6aVFOwFfragfZCw3Vsh3x0IfA8voG+fmWWqaoJb
4gBmjicnBZMuLnG7aKaaTnI1v7/fPH5mi4ESyTkziyDXmMrclYGU/aZTn0Qujves
Hfn1DjjK7LSKoIpHBqZ70+jAP/KSD1ULGuh5vVeOpEl/kWABujIDyEDzXEIb7Fua
7K753v1nHiLQ+Wwoe1D6A8DNELwu/HQve1oA3tJb2XsQcPbQe3qjZy8EoLEeUXUp
EX/X134aH/1NkgqrLF/zAqK+I6NxCYaPCxNJePXuBQlp4rxo65I5OA0KcS2Zev2H
q18TgQ4iPCgtJcrGs0p6w2z9Gi8a8X3XbM/7gMPj6B1XX9I9Xi5BfaiNvg5xoEO0
ua7or3xSS/90B0WvISYfjsX9yLExAQDTbRa+sepHaf/pd7x1ZJzhzVRXWPUSUZ3b
fI8EB4Qj8Q2VxJ2ixFFAYDrtbVAyQmW2xOeoAq0Gdr0zsdon7h4o3D8I1XLC3BKK
OvEUSCqmaTRbQfTKSlnO6eRWqHra2fonHVagkostcuR3MlcNowDYkP+GkHDm91/J
TNZxIElsc7YzsQ9rgd4CnZHU40Ei/qntquUfFdknAsfxs5AIahGqNrvjT8BkK7hH
porZf7b58f1if6JNZmG2j5cfNJ5G8nP2BOBW/g+KQrKTpQfd8KwgExmishAW6rIb
bQW7TtG6UCROMgZtzpEqVN1p+MuH1cKtjYNg1xYclMt+rTTX/k02VeWhr9l1zz9l
6MoKtro4PMYIFR/cnQayVxSUnkzxlis/HbdMEUYo8VGFVXpk41/zRfLMRcS5tAln
fTHAxnXrXXzfl4G6EQF1d9KNaxhQF+cyzNYdp2/g0fXOe4RVp0XGZyPSYYAbxyxN
ApVTileLDunV4BlH6Msv16gdG0tCU5FUgPKYqkxa+frpY1X50m5oD1rwhbXasYNn
DxpWS19V39fNxhacqIabI+3GWjKPXxb9Honj8kiEwxjU6WgMZT/5qeb0d/8dPa+X
494MtBrCc5k0ON0t7pdUi3RV6OoqMl20DXOYOcAgnEwniqjUF6TFRBd4eHbXbj3u
lquTl+of0Vqe6RA5csq6wOMSJF9jqvGtP/CJpJD3aJGOEyvD1kF6R6FVCENW8rkU
a4fAJmX7xB320t3/GQnny+Q939A6iIaMA++Ydd4gUBjMMmYhCKdsmm5IymbNJ1fI
fMwbqKrQsFW03zOra3ygJvNbruXGxiSclhqkOH45biECpADIofwvZB7J01Ej1ihH
XwFqzbyjDo2hbPwM3nLGvVFOlqx3GoAcsKbgFrPZiPbuWzhUq36bxmcpAXtWxdwp
XIYbbmdspHbIDUNxdxPvnm2p+8H+taU2kkIgNO68LRtaYkpkhiT0hTOjXovh3grz
ZPpPc3/8fvlvvxoX2mlYHREfz9AKOtrbPkiRvSqA0dq2Sc9tNJmdWFxr7eF8mWgs
cI2CcpiJZFqwQTYtUcCm7BprHYpEXfG2AudDBseG45KMmHBCuc0j2nMm4Au4CSr2
WGrEhEzgTcYzzPmWcR/rFhDBaoJCRsRq6RZNZgXxDM2GG8rzhCg043HCHs8JECmR
/8a+clFsgxZTJy8KE3buY+OEuY3iWK/3J5KAbV7kXDDsHev900KIm5yAVmjrwVnb
/9PDdb/DoNUNpMUlqQuQrcstrNesqQ7lXp3IssQJQIfks7AE+B0zfv67BK5jVbNQ
HXGZZo2rFjRp0/30Tqlr/bE2zV1fxLcHCWX3udXv7QRvm4ieLHN/CJBEs5FR1WRM
UnovrIY4zC67qZ18wvL2qj0l4nFpLoepP4mng9V+Xehe4iH1gw0XYygGMDkF++na
9YAi5RFajy8GHbGjo4eP5Cvqu3XgasfYp2j05keKKVb73+i3tWSu1V7tb4CiwQZ2
YYsgs0txasAtOW1zm73949162k6TURXJ/XF90gxeIFkY8q1rGrQxC9Ot5U3bC1yG
jVt8laeLHNm35n1Hfbw5pHH2nLhhPRwILMkAvccwY1kI5SfgEkeNrok+TB+tGPpW
P7g18ThUIXw4Gl/oVQKQrbnufOs6IwWWUal8TBQ05uGVxiljtCa6wp3xtyFmfpjk
Yk8RNukJ/7/o4dE2DaGOw9LAc+3dN95y1dPLPBRWz0CpjGe7thptI5vVHmHpLmym
J/xLj+SaDp14T3Qcq1vqtGVrQOk/GFhJDnTXs8T0DixIzF6LCJ3UZ21Kgntz/Kcj
7nW6fWKpReSvAGCaGyeJEu2JvPjLJ834VysMkNtcHQ1HZjdwz1Pt+sTFS/Kgtuo7
0xI1ak0NoNoZD1co9Rk9f+cS6T9FzWNQhj812vqU3jr8J1dmxxEWy/a6vAl1v59B
EPeuXoDK9fk2RNJLE5PQGMu98udpJMm/DV5Z9YU9Mg3qQZqLwK76PJA38T6vCtYv
5AtaA0QvLjnUVsEQPn5ZS9MOiz/t0Lng89i2tbBcEA4bv7fqqW4aZ+R6n90nVKE0
2bnkDA47jeW2aJeth4QNqDSikMwAp1LOLMVyzqWkMpOJ5sZVBsiY7Cw0Jyn02MAt
EbSecGeAmGWT+VATAN8QUs+NfsRQsJ36EE77jlX7/B7FGmifdEt1JUM0TLpx+474
2SC+0PgzA3zHS6/L590xkmHLN7zgw/7QtELeHhn0gx5pBrUATAtanRVA6yeJ/CNB
yhTQbsYKQC2vQ10weWs3FrfWMwqhxa7GrJGF2kcVBdFgEJ/gAOxz6V5Yx3Zu1mDW
nnjq/DeeVrd8tWOHmF1IaQIZIPj4SXLEipusa2YJmzP490FnZn0d6EKhsNPPbab5
Z0fJ88ZPFCmksqO8JgTMj6J7XuWoeQNYkx/AtzBy44aXFsOx+jxH3lwskikvsdbC
6qn2TBDQoxGn7XhC5g+wyApPcL3RDI7VAjZ43Q/6HlSgkJe7OKU4DY3QUwDe7IuR
4SjmAD5o++mUuftoCVKnXQVrnw4rp8A6/48ELEdTdIItvWr8wbMnKrlcWh//yeS+
o/M7JpBd2ULKiyXeZPjUF+pR2TmI3kRSCcedc/c2J3hY8Sgh6YBAjd8Nk+o1PZNy
c+opScTQTvXWvuNMiANQX8VqlfelxqybtFIpmpXVTz5OSbWMaW2dfb8vFE3waWhY
Zi9gn9KTKUJXe8TCRNo53mToU3TyGNkqQtpSe49yQHHIHlFyEVgUQzhBIrVS6lbR
CMKUPKnWRGVjJzBgat9btWpbTagKT1xVzbrTf9lYguzDOnILtodLF7iBV3fsfMGu
AYaNutq4a7OOmpRK7NPCgrawxg39jgmJbgfL8oaYoHjD8WolruC6zq7t15pyVkGk
hdMyLcZM+jOajkKRBB58WNM7ame9e/moYaCSJ64lXiuUhV1UA1kQa3Sk45DRM6pj
mnlQGw7tFWsOWIZe1bNu9Xok5C69FeROcCzp8/KoQVbsyPi0K93CnXoUO54KmNeY
k1ort8CWQ88Fx6+Ie5N6gPaM8klVeNipUR31N5a3bR2LHm47cf/EDlHDn/22Fq94
P7ay60r020EYQZvD4UvxB7KWehVFOnlHI6bxrMBxUWAtWuXAN199VBEl9bWnJH0p
L+jNK2n8PPsUVBLs1EqhrRmhfjEMVaE/fmFn7alTKRHBmLIitl6PwLM7RNrBsZmC
4EoVik+WyIAlWUmgwiggUGvNW+0egWNjL8gB57Soj6L6KxiBKKwf1pXi+YA+f8W7
OWp82G1foMi/kk9Ug80iUmB4UJzvMva8PnaP7zvDF1hGbpRCM+FXtJ5KpKXX86nF
8ee+eLhQRHkKvVVH8gnl28lpbXtOEbR0LCMaqx1fgBcNDQKVTGUEHy4Pk8UQaudS
Wq6nhh5FYXta1520s/IP3XIOiGE165p+qtUNFai0lApXqr7U1nDEaC5W4gSbOxvu
ir2bmiC/0PU5RsKmqcRm1AnYLGCdnHX882Ip2O2f9s/ewaqiFfUw0bOQShf7FgZY
5P3O6gxH/5V1GPSvW56sw4NRnSJyXfTGzvk5ks8FVPYTJkZ3eSlt+z0sOTUHeCWx
nm6SrRHTGQ8GIhnOqAG52alf4D/9m/2sdOj9TskutH1V6kE0/0uQXTcsLbAjH/oK
U0ssdTyTy+TFu8ffeuvTUuQHwTHBk3HUHeeaSsq23qrT2qH+LhzeVJk2CdFzIyhC
ms4+MnKjmnV+3eXBSFF2GmQggqUyGi73MG8EAXULKGI5dOP96iTiRnHSbaQ5gION
UIYPItOxnulsavXAo5FajRxR29l7Dev/oTe+FfKMyaeoEV/x4j8/NEIVVJz1pA83
KvNwMpR+r8TOio9ZWhNUX66nJlUO+VavFQavf3h6zJ2/qxlfLoopiem5tGahvU1M
l/5TAQdCrm9jFdsZ8mKS12Qvd2/y5ewduySNHgY9TGBBumZBxDEzIJYc0O/14Kbn
X2OfDVCQompHEPYPcC1PisXG9iL6fGnwuJB9f9fVX7ONygjaCV9jQ128HhvqX8T9
hFbpb62lp2dUJFOVCXUqPKZbD2iXrGAO9+cg6Z61lHtj1EoWnkM1rGbTgfHr+mCJ
hqmz4YxUSerKdNaej8Z3xGqldl7WJLMVJKglDVSK8vmSwd4qHG5TJriK07CB8zB0
TdQbleYkJkmC2Bz2eH2oORIWGaSHMJGRIzRS+UbcSl9QfNeuQBU1+DJ7/UoQy1Zk
qusBLUGh/v+YAHfYiKv8KlijyiR0WGVn4BRba8syxEZcoo3JUybu7uboxF3kkdv/
jsRmu54xOIwkaj/xpCZ1KFcV9eTcf+ubbsSuSm/iZS7yvA3xsKIi7MLY7tAO+nqu
mo+4cxmLCuXY8W77hE9QyIspty/Cvxent7wwqv39GA1uMVuwc+pID80evdScesG4
RaHJMwama+O9m6zRuv9WFQR9sfUUmeSAGHw5cDMaMoc2xHSEjWUTAbzmlt47Po2B
wxy3t5gFvp3chFG7ZAjYWKxjYL4cmjs+23jEfSLTjbGRf0fmxNt8U7BZbgIcm5nz
OwUdxmvyhkuwY1ZSZ20Nk5BnJb8T2qnRKDwJQUUoQPz/E/r+MnETDxZpKAb9hqJS
4aR3D39I1TzTln9Gz3Mt0QKaYqMRSG3gn6rpzbHpISvVuNeBRHzV8tqq6djG0a96
6F6HNXVj2bL+vz5qohLsRDReS6n99NRJgSJxS2yFF2cLEF4wUIvEgyBkuSwOU3Td
emX8ssaAHwP1S4PSLGVC9MUTdeM2jYD0yCYv/BXuO+BwqWw3wr4WMiT6zKcDkdhX
dLVPO/15bdlgpWp4cxU3ZSgzNvWpllRSGlZFNlOER+KitFxfPNisSXz1FEYNL6Ib
exLl8MbT9MxXekNsAJ29JKClVP/KboIbXQuRFdp+NNpCewYrNPqRI/1BejgyU52C
4gBiRYb5OdMpIs3woBgdkL9wXrpi1GPnB83gsZWd0bN5BMvcRWktcuKSz7ykHb2I
AYIaXAmQlmvxmj3RdEMlvzVBZ6PWdiAut45IrXToEZF9w4qrxi/XkftD9GIkGzNz
70fKt5QvJTJL3K0mCLxzTduaZ6TzNAWdc7ChLyGI4CdQzQMBD9W23WfcKwdv72Bv
9D3iaWznWjUFuihGLvdt3iYyu4ef7k3kcuEdOGpRgTYJWPbDIYp80vu7mQp4K1G6
Q3WUnlnEvXBacSEztyUHuGgKiI5hiPYDqoCi00BASnNOEUy/MrtJaXOXxh3VS/iK
yrrLKyCXUYPxq/FjXD9042qBI9yJaY/jKp03i46SBCs27hf/6/LW270q5uz0t0+c
EvQ/sAzF/TaiLQT3Hb9/ZAkic9kmt2fTQfBlXbBSrg7VAStCbpHW1LzmJy8otXcU
n78V13FLlWJ+Mxsdt/UWZFx1vGlOzY6q6TODhOafi1bQVdxunrYmR2OFKysyfFfh
5rmzNBBmFBi9aQfA3aQ4k8gTkpmPp9X9hyaomi6dQAG5kt25h47IGvi5f9q63PoK
OmKMu6RCrAfio24vD6b8LJCFcCRwYcNgFljod/eu65u7TFeVVKMOrjIJOKWTKB6f
Rs35gHCUaCBxRuWuMGDAXbVQjy6/IOSz8j5CxIjwlRYt3maxRMEQT6RX2T1kmXKH
EEGl64EzBlMNrX+TtLRoxiB936570rCtN8L0zMvG8jWObtqJmkzQQ1HATTgLTTYo
7n5pQScbB7KQpCRWUegLF413pVpI6/ck2+HwVBfhmqjENDA2pgI95NTp+x1jiotB
Js0eRMVCF+ojxgBAoSEnCbupZnplWUEfJq+RxYyy83J8HJc0+ACZ6xoERHWk7Emn
bRbBeleQnTXolAA0bZllLLZZpnB1UZ+uz7sGW9lJohgmpMJr5ToCamycdrJoZHss
bo+wjstqNlqFdg5W4g4mVoyZGPJvIbMdMiHECmjW4FiroqbrkOQQwEzPo8ePkqaT
nO3ie3gaMXifGJ/SmZ5gEfqtAHQ0x1a0orlGgs/cG08HQdt8OlTA3GQRBTD/ojj0
1zT+YHJuRpUBxIXUpfgoSEHMJrxOxXQSV55DBYQ2GCXydrXJMUlASf93ZUxGHjmj
z7M34TW646YCQmru5QHWyOxOmV3aTcQ0DrbD7DC64p3vdckOjLIJodf/4uVnIONP
JCiciVXQsyQOAm0sC/a166RoR6WvKYyw75p8/+6xziK7JWmRGukUUVzEf55Rt6s8
EUtG8cte+8qMSldA7Je2eMnrvTlMLEPvs3yU6e7B23vyf86V3Y28o30L46C5I3O4
2C/LoHHJBtDxjDeriMN8xgZ5XiO/c35fxt86OrHapYGRC1vrJoZFtcsnkM84EZ5y
IBfSc7ULRmPrc7Yxz8H2/pI52v3UffK33fkrl2R3rYAYnB4tVSmOwZ29p3U0UtTk
ZS1lozFalewK40NR2rYX/pl6847N7lx9P3izh3C1W6twhXNXYY09P1MNHU//hxi1
TeodKPuF1oLH/qt7oxp/+sAyaB/gcRw+gDbd8tH5NImyCjTm4DrM9trtkhcPZJu1
xIrwIsjcIxYmeJHPu6IVaA84xsbj6akj9rAKwRU7yyn/02pGPcwMeeHGUCOjUkxq
RsEVo1+LV7pWod7fvufAwSyxXCcrW3m3xBmX08Pqug+TTms4v1ghqwCl6QCOvuER
kh2/bFp4VKcKaTito2N37UQxKo48eFmWkUnBgnumbSc1GbsFalbvwNTgYar7Cbs1
MEwEoMnA1UvfZQvsDyQstVmqxMEN4764STtjZIFYVowhZT4D/eDJlbx0QZPED577
bAFse9HtSwbFUVoSKp0yPUDxrhLUDc1kgWNvOwUVoSQduPTFDdPaJjmYfFVZlgDM
DAyZz+WaZDvgErCEH1FGmhROnWw2BwyNeNHU25D1W734osiZsXVDAQoUf9W7HTMB
lab7nJn36xMEbXSNcienrci54FDF7eRdu/mk7A9FKn3+QCClrmx9V/EExBkUA988
k1USy/0LxAxKQotSU0qWDuuYHbHzLmcHa10nxeHcqST0KYyrDEmCUgNfAaDGbjl5
tq+J/5QcuJpU62dwZxeHow1c2AHm8C1z3P0QmA9iCVh96tgUivyZce6T7pwXG3+s
oHcdvLMWi1OXIBG/Dn+UrgTzeooGZFohgMcM6vG6KbP2foxqjdW2pHydVSyNSWKN
cgM9ksJpA4QK+pU7Qiai64IvFvgsO137LVi7vE/JVwk32N1Gn93pWuO+l1zHcFKk
1YnP5mF3H+XhJDqAVnhJYEQdH71M+iA0CiXfFiSEaLOuPabM7Rr53kKvZO362xym
F0NItXHKc2YQOflz2hp2yFpTPBLmvHP8AC9lp5RKqseRmJVBz16hSHqAgsya4sJQ
jQVw9lDUhTyxl6jgDx1JeQFjyVmhWMjQTr+ETLuhgDyUxZGEBJUvmbcgnY2kyas6
BGuJt3E5x3aY5JjwgUsnA7X5HyMYRcd5whlgh2cZHeTKwMewX7Hhp0vmI3teUcgP
ZoXqKTIWuHB9kIwkRPSU9HytfABwcF+hwnr1E73fpenogmMeSQrAb7CSLgDXxtKQ
IigAzVVQrp7Q9ImlAN9GvQUa2ybrXHf0u2e40Co5/7bv0PYz2ap+MpyarlgEpczS
XIeFy9zztAow9vq1Sc7idJiAC7NjigNfMfexDnEr6AB4pNajN7xto/p7vGtus+YR
jNEIjJkbngmxRk4sjSvhLMNFH8aRpYPR9TE5bqZpPax8to51c+gE4WWLj/SI8xFz
Ghv5wpvIAvUAIaD07M5DQORMj6U/pwREyOoupXUTTb4q1+D79pcOcF44NuLY2gux
bfzooAXkr8k8KinVumxPxZxuQxumlNR/unV05cKbsHB4INzsZxwPDro1fyd0bHl9
D00pIqo7mjB2JSgNS9rnyvojgDPrHH+YKVxwtlFPuiQtZaK3YJ5+ML71GzrV3mij
SiOXn4n+FZ+xCZrSz2Td66z3v+Pyrawxf0YayPOcMGtc3p0VzVcWR90qNOKdPWoG
FiNFAyq1+f36bRN/llO9cQLS6ms3Qfc1+JVkVCbl+R0lfAUzF0X7oINeK4nrmQhe
Q4TNTuCambVvQnj+VwYAvmNvHKPbsTxxPf0RYBo5VpvSOsIjXgy2W1b+wrToml1z
G/7LzlREesPVo8d6K4SKeUk8GNC8aNOR8EYaZ26Q/+jQkt85bpm2eK84Fi/r4CT1
DWS53ahgbYXUfy6a/bHSbnZiOhnINYlkRHYLZB4bjYVGGBAA8VMrOdEo9OTOo9SI
/qGV+jY4159yMeLpwkk1gHyThR9ZvEqQsAkSbkwg7I6VWyBdzHP34J6IF3ajiloL
RPQkcGkvbj8VSL8dCzgYeWUBtr84oWtnOR3fg9tkjb39xkPDThCAxZOxbnd01giw
ZT+nQdCI/FPHVzQ+FZ3ThVcmABtmFhVSk2uxbguNX+yfrmxO2yPOxhTkN+othLaw
Lil3NaaedTx7qgGVY95Oc5hXynmnk8VtRVOKTEZ6N2SM1p4rOapLqoUDPb1Fr+KM
5pQ4qhTDir+2M5pU83ANkeniUrRo5mhMZ9QcjpvA6eFHUgfx9US6W1a1byoL5yCZ
MJX9+ow/3CtsjzbVt0cnvnG59VhGCQ+c0rgcsP3PopnZd7Psdq4UxlNdSTWDX25K
+SAd7iGGUr24T3L5YoJ2HDg7/PuotMZHw1LUyjZ1F6lY7XSXd0ParUtllGr4tkGS
eLY9WugE2wSkaYtpnqiCl5S0IQxx1tTsTXH1C7eRUu8xhqDKv+LsYlwgh75jRBSa
et/KeqpMu/WghD27wzal8c6DT+LWBmjtaJFSAV9KE4PepZojcpkiI1L+Y4VOEwiQ
WT6VnCQ8Ov1z07GXlLWj6hSYjbsUz0PIDWea2PuE/FhAoS2c1vUXoBAlrfZxFywQ
9rcFq5q5ggad4vueoWrKKh36/uq7WA5+IYrME3dcrv6l0BI7Cr72fwI5Q9B2+8mU
F7fDeh4fPKz/bCX1pDXsCU8DuXGeInWSLnHC/7cuAVOhmHD5wd9J3oXJAG06KMD2
5uB0wgEy40K34U4IVkV505uMWTU1ZnAVWC3Y+rXs7A5pIwzB00ZSQu2zLzJDSLA9
aTqFxBlUt8rUwwUFvWuLbtroGGY6uGWl+hWOHngRIeGrcxgG4QQntZ6TbI8Vv71N
yn8W0/0D8hQBxhQR/f3pGc43gZBVrzBdr3ZYX3avLBs/KBeBDUBbGFRdWEWMDn1t
rgbizb/Dm4zoQRo1Le1gFk/oG9l/rQ1wxqPVGoFGk1tyvg/+2H5hjitbExODMP4F
/n1SDn3O2ITF74U06gkbkO36QaZeTHdX4kTvyTY4uZjpRg4wcM4mGzXGAs9W3/C5
v6tc53uLcOjnisMrLS4UQL1Q6nRfwNB1V2GT/laoWoXCSI6VbmtDzZ9NClVGTWcE
w/EzjxC+Wed/xrpuA9kwg3AiZ0tP0hZYCBtMAlP2s8Cg7G0rEXaw0ypmBPwygSXo
wtutgznlxtCUBOF3x6T5v9KcOfF8smOhN1vxaEtjfSDKahnyBxdXuCcDJw3wCl0+
WbDdzi7RGuRYhRrrY+onRhg4Yvfzsg8wgPGcG1IA8K/xi/TWxIAukLdyM0fQs9Gd
rhes0qvRKCZ0yW/IFmaUqn0A0Hll6BvdQ+dTxrlG3Nt4+Wmf63hAOPQRE32MJm5k
fTpn8g0rpESbZEksHxT2nYnkA8G4kV9JGOqKJJ6B0ps2uT7bPSK6gDiBN9oJYdtj
u4UoOmUaWxfSMnFNcJm0W27ZxZOuVFPAgbOm9e0kWevH3jpdWijE9Cd2yy9jQ61H
26W0wIBvp4ZvaMl6F7gq07Vu3yDTMTRrjEmgwigS4aO9hfRL2hTqueXrE+ikJ1gb
YQIxbhYfrY7ZS6RZM04hLB5+qXw3YoenriCt4h9CJ5ixPLMX8oLqO5MyRFkvfEs/
HZ5JQGdTmwvFVm6TZUeR6bAuM4/el9hoGql5sGB3V8sj/4CHk3K/iOXPDBY6bSQy
v2SNLAKE77LVj1bI/wPdcy602kCXtKr5e155GJkrB48fxzsxrC9hQSAPr5VlvyiD
FGGmxNL80B7FmnEb9XPGEmsT8e/hgTIibKVLuZVBr1JL+OibueqmUdp7zZdbEZQJ
I5vmwZ1/kvH1/jMGpRCP+JoMP3xqrYtMUWmjBhpPf+HB/iF47Ferh+opeTLfI+bU
L0zWohXVUB37ho+h7W7pP1EvuKO426t19j2OlQfN40sl557ZcvIpJV9rQyhIPRIk
VmOsY+fb2gnUEvx6qLwm1d0QJ80VQ/5mLlMZcjcolURbHQ/ce8UfmkvDXtKm3EwV
MQNAAaqEcqSOs2ye6ZA8G5/xT0AeuMINCzZqXNiv4xjuIhqkZq9AZXCkjjwtVIPL
b68NJY/v6lWAZQxSoq5hC/B77Ffx5vtMO0oTdBNq879woTgq7emanZvwaYBZmPq9
Zc26pNZHBlaJtTcJzR0yGRRc7PJEjaOJQfg8cZDM51tzau7n/z4A49GucQb4r1rq
DFbyZJEQQ5YyeVAjbFknmMLnXvGVQbsLxrbCJWRLdZZFxwiKYyQjSycts3fIGZH/
orZyRattcj22US2fLco33hgGYgDNqAWyQwK6wmYcA1f+w+9FDLIMaUQlVxTMwEJG
nc30Same5Z+on6j6jvDaBb0ImCIQqgcnU7QSEMq/DoCpfEbBb3sjtOgqyHUPqEgO
te2Eif0lmGXvgIraA0M0zbnk/eLNyKs04LqcEKw/4GuoT4jFeHrKxLTjLCoP5dWF
zDz0y/2TlUgqPvlUObVgsQ++eI6UB7JeJBPmNX5e5yZykn0Znho9zbUQeoEJHc6Z
Hk7PWWqdkxWZOKiKnhX/AooPE6At8oLCt604Es4Sau43lwS1wMKu2yA2lQRguOyf
PxgRM1xYxqm46rStSVYrWM202rM5x/j+4wfl4nXSiW3ngGLRTPMxxp33rYSmPj25
FZ3nNC9x//2D70n1HIqM0sraYlqKkKYDw6r2syQVzpBGIwOyhOi2lsVFxJjqJpTo
U/JvUKAhT99ItLasDG7GBCwQ4DP+7GsSNK5f5zX3VPhqjnR9RomaF/T7Ayoq8huA
zJ1Prvn/1Dv/SC8uTFNBW3MGBFGIrdNg48d6PWVOl7LRZPI8+SGsaBuzqbE0qku1
EBhu0meOuq0JXkIdeDjiwlvxshysAbWSAgFEh7fUpjxDI+3moIDwQSlrNVWAUlRf
OtygUUHgaeuR59yIQPa9vjNI4/tD76pSctnS445CCp02PLAVyV8eX40FpUExGPIN
jJy+GFFUQ4u4Za2p62zWYq8OGEoaO8h6Dmvp3UQt4lnRjQRoRp7BTrl9NpJ4zpct
/1FzAcHlm5ubGxrbLIfRhd8kYmzvm5yP8fW378K95X/JkbPnDAwX6vtXsNhG4tvz
9Imdnit34oUOs8mKgF0qGxbarFyY4cBAp76oWv9bAszLSWmasxuABEOLTB3h8mUW
7xp6RIUnaJJ2m7QmPsf5gwSy7Geps7II4eEK9APJB3+1gs458qpyujM9MPbwTM/r
VRfpqld6aZu9Q7megCdDw5SX5I8cZ4JcKcrC3n1L9s1amVs9a3IeS6OCpfPjf387
22eoBDP9OjOHtEG3Nkr1a3MRDxU5YXDAowM46B+urEvJ+fPnVth4oh6+W0aG7Lyz
wmrKeOcsmIAJ8RHdsp4G/rpKIeIrgVvkriM7C2zbykdmZjE5TyWVLYiiQ93MDc+8
yQy4Vzw7aJw2POWgc9MBdH12ndzRO3YR5jPv2z64dYzee3vfyMOLMTUPngY8qT3k
o02rncnGl99QD9TjbtMbzgfufXF0lXaTk0lfVzgNT7LQJIHeZSTir95LC0enZYMJ
pIEYILMtOOipzM+tnf3LIaQRY8L67rUHuJN1v5WFOY9MSiL2KPH5VgEBBkVkTnx0
v8yflaeVA1UEiYDpQtsqih54JZKKq4FsboPgg4v2PMYBGXBwEdmV5luvVEtqQ2uh
jffWdVKF1YQBtdf/68T89d34KsWnoe/yn75bfKRHeZbszb6azVFmHsXMSYyJi1FM
rZygsiGOePOqEomYsJGfmAj+TM5khmHXza68gswmD/sQe1yhOrt1uGCiLBstUwBj
ceT5qUiBOgP6NGeDHPwYhrwPfN3mCZfFh0fll8rkQQPJap22AXAsnRgj4WLt07A+
FmMOxdVFy1vTfdEUC0hIM/pviibzXo3Q2oRJyV3wg1fSo8o1AQgAhfs1lyxoBoFC
rV2tg1GcNcU4SHldOYhDnAp9K62qqmUlJ22B2nkJ52ODETkof7oK3hgsiUh2NfTL
09cdn47eGFBmw/ZZr7nRkgfmTgh/Y7ruCRm2Fyk/kd5pvPLCuyFPfSVhpLuzk8Z8
slxsppC/mtyYY4FQXE2H1xq31ums5Y/sYixvbk6D5q0O4Hseaap1z89YVWT+0EHk
h5X5Q9au5liYEyAkuy2jAwJIC1gw3FbXxrkCMVhKMlCz2mm7EbusT78yz/BlssoW
oxiSl1jT7iKq6rmEjogeeU1rvXgPl+mMg1/pf0tkOBJPSwT/ASBZneCTbKofd6Yt
bG598XUE+zNk41qAKtjrcAqbphuQmcktk9GqDASbw/KgOf56CLWWN6vu6cdkd7Ql
8oEraGvVFoDfvI6QsgdmlCVQUPH7kbBBPn1ZtFw77ZeOh26WRTjiUSToC2hKN4Af
ZpkX6yeIugMnnsF2212D2hggMdxPYYzYJa+bnesQiUwALWgMOd6lTVkOJA9XHNSk
1s+f0FZbCOTY7nmKH5rZT0z4Plhsxrk+ajKp0qm8La34RgPsXDx6uaZfAVgDlArR
HfoyDOe1DMQgQ2x+sXZrVvsbBjVUMs4tOjGQowvhg1W3vbtn3GZ6o+Ku+pFjUmtf
9GT5QT5sniKnBtw56vcK/jBlihMjdzqW3uL0WEfoV2hecWwok0ejEHXGSTUqP8+1
Mowl4ssH25JSyv1UtL3K16TtM0z2EWZqUlC1ksWAF3vANuH6JjjS95tRkEIRWsx0
f4+O/tAvOFNhR36oa/8U/KdIEsiDRhc/QauiOTVix7zYJJMNr6qAGpSyQPDgNSRb
eoaBKdAxidcXBTecEbjr4BbgPo6iEMEOhugiHUUcRV5V/9k1Frl+VIIr+nQqo7MM
EFG1QGEZ6KWHX0dBmP2ACdMJh5MCTmRVmdRo9ZzPHtHeINJdlnLuPju7Tutcf+b7
eRadsgVySIm68DbFUQVdRMDFXq/XzdSO5fqhYEOlK8KcaylrMGz0kG6fEPJh64O7
BNpQGkWaD98+KqOro/BttSGyOm6gik92Cq/qDfQXITXuUj3kbt3NNNYPoquWzRQU
ux1Zen3wPVbUOREJZHS6hOYqQqQ/y4MbQIU5ILMhZjdottjhBunH04GGevlK1RG9
+zB0kW4IIn84B4sPvGcG++DLerzI3UC6niAcHKfFO6n8qQULoynP5mc9T93BhKB0
p+M5NVLJJzeLmmnpFKdrUkhoIJUFFPe0Bsamkw2OyNAc6xWXCibd3ZbRldQSlflB
SKx4ak4WA5h0GwZElgaYjz+PQSaRIc5D0T3Dq4wVgYT6w12dSbqvEE1FmhpdghgJ
jHqYvSW/rltTnHtZmohY6REWeGAfl06KRuMumjzNnA3DMoD+8ENFNdMqvh/7D247
3PaWoO+MEPza1bHOaHVotCcwMhJTId7VYQ04BFca+xWsOH6Ja8/aNVSLn+Vf3Xsg
M34KsYHcEjPBoCKcmGzw42ZXdOLWLiqapvf/EN1t9zJ4yihr2OUkKUX4vr78IZcr
bMzFlJtXNoKKNKa9gCaFM73ywaRGwaLJePnMH6Qf0a480U1WgZJsIgK6nEFjJ9YN
KIBBJZjS04LzwbHfkONnvzZjiDunXr7sWE9knJLen/Z+QnRHVgtzgpx9waP/UqFZ
4og6BgS6iOi9clgaBfNfkxHkC557yotYkE0XS3KhysAnzRC9MXRnrXVOsmLdQm3s
WShogulnRNZE20Jk8kZ6UWNROru/dJzkY7oevoouQdTxm6+6pHJ04MtpOmLnc4tx
oMvKv2ZluLtrATajgtZTUVoo2uDI/OT4sN99jrpc0fhKeSUMsg+2r87bBga/hesD
8QeM/K9XMEV3CmRBykzz+0OigEL1iX3phBTK1GoyMetNOG77DknQUj6OUDiWTo/s
+gdivI0q4idPNRORW826//9NdcWmMnyiqwoYEpM585FT1l0v6DZE//krAAKjXpGV
T3eoCrkf4hOEF7jfZLxKc2vLw+0qqFxXaqHu6CiLz0NLKFANk11SF3F/h+rwP2PU
T48pw1FzW/vN7egethM6IWFg/wDXQbXCsYP2q/EfPZlnYAp9SOp63K1u+MHppTGm
km+TLZN0WHyv4ItDcS9bkC2IJ1ckjDcoACLXLTbCIsZZN6ZKELMpRvZoVD3JjcJ9
owfeYhcxosMVoUClRwA62tWx7XCIG8fqv5E46Caq0gM5dIn2R/M4JZptOQfXcyxs
paBLEFKoaS2ELxGI4E+dWfqMTHu+AQ2a8NCzCKPM0J6fCNbh6Vp9d7JYm1d/JRU+
OEfigSC6c7vzIo7ZG3BC5VKF6ZeV91Tf7pMi3cPb6l47PvqZI2xNha0+LSva/hRQ
YHc+TBlMH8sUQ93k2yvi/8JPlEsaODxoBuAOSk9aJLefGHClOjqNLcHzR/6dQ3jC
9+d5RhHjZN67k2/kRroxT8i87LJBCpJKwCOBRvzIAiz+Ii8Dzk7souQ2v+//ZulI
huJiLFhpQ/FEPsPvNSwSPWe/e5P7voJkxAHq3r5IPGV6svQ9wi33dyqo8CtDR0Xf
x1qZgkT6oBG9tG0VopQBlzIb9+odnsBCqqGiqhHqLL7YoOLynNFrfpa0qnguUGTF
E2GYb7YqLD+5AUaOlYb+ouZ8k/Dert4Rk9Xsng8DQYhMs3g2H6ierJd/fce+TS19
9EY5upPDX2/ZkvsZSFn0bfdB0uO2TQ/yTDwEfOdx3VoDND30u6UWWj0O+wk3R+1n
WGyd07um9wZHaCgSguXtorNtpBm62cmILz3vTD76tDKJRSkKvjrS5KOoLy4HdAq3
eI6T0jPpcqFIUUG1G/Hc+zEdBWZdxeoUe/DasNnUOxb5Qn+TGOC5uErKrHfLl5UI
3zp7P60L//BZPOniR+e9KjhYH7T930gIXTY1w6HvqaBqNs1lNKMPxFYkTjPrXYlk
u4Hp+1mS6Ort1W1J62TKOoxnig/QThOU3H3X54AtctGCjAB1o8O2TZ+73NH38ulg
0PuZkgyyXF6RJ6vqz7uaSz3p2GdGbF+oasyfOgnaDl9OJ2CKKgHcY760mfccABqE
41WQwucjLw5NkLr8xWXxDScvhj5cy9aGoiF0b2pPjNjqTbgIO+sp/+E7frGes/Bj
+4mpMU7GulCe7DrbOo8yjoVNMnv6PwKLcZgWhyi0gTnPhnh3a8PsIc6HLK4c8UIL
E92V4ujnMUp87WUxshX3Z13EuQof2yVUKz2SjKyygRDIwati5CyaDVIK/tTf0/mX
2vaQjQ6VGMbPTbauSn4RGzqU/jqHOZbvlc/zh1efSPGq8tF9FzhOwfz2xdeVX8Q7
IUhwsNUdqHBlw3L4dweJQulHLEJsxVeGu8JEvTzYeeUmJfMUKZbqRrtU9OS2izLd
JHBc2duRAIXvUc5S8f5z5UktkMxcQ3j8ladYR0/GhIE7Jg/hnZ6986qaEFP/4MPL
QoIaeoIyJHmgQk5jsbYiuzU21C+5Xj5hGdW6TNcv87lOsbuM99foB/cpIIgKSn3P
pQvft43XG5Ixcg53O16xX7KvpaxGz4j4P6/ty7wA0bvxwxq57IH+7QNsiAOjBtZE
zc6vftSE3m2EKdIyoGFroIGNSBAIlStpLfYGh2D9b8SgcpFgUX3Q8D1Ecj7At6FG
2n43Df9hx69CwMJkRLzdHzlXQqCrhhO1ja/1+z+M60VHb02Z7hx85ac9BGpj9mGc
2JTSpBr5Kvi4TbYwrqb7jmVdHEcEpnDdrPbt7pMGzyi9ahzMAnWVMsChhUxjX+OJ
WL+LIxK6z8TbdXXWyG96I9CSM4iAYwFVdQ5rEFkG0DvRx/+bGJ1PytGM/yr8tDE3
CF8ROcgqrt2EYZMGNnr8MsXDqgvjGPkNmAN3MkWAYtR1jULUxDjMiaJ6byC4+SMA
I7lEkJ2C0VtV6Yrrv8F1HXlfJL4rIwn6DZp4J/7z50U0wiMtdVEiryUpWV1CePyx
h8+J+LH0mLhePCBAvwzN+U3imMZAIxAQQyUBNjTARjjzl3nfpHaOkwKXIjxR4WAQ
JyxuldGGAxcp6Rrs1VKG5dZZzDfyN1WwO+HRxHs2vLdXkBH98BXVjHUJ3cPiQBTO
qBybMRdTSQw94pfwzmsi3ANmrUItjykq/IRocVepU/B1TbMObfKF3R03Q9zkvBIA
2QP9GVw41Eg1wOWA6fWFamLDfQ6LOiLf4Hmty5jy8Cb2BTUkh+S6vXXCihaVSV2q
AsVzWbWtd6SH++XO58u50M8YFFHX/pDBlCWSa7oDsU2IeDdD3Q9d99BRNlEDz88Q
KoWC9waO0LbdQUyHDSbGCL+3Ul+qU5xM9luGb0pScBPAt4eqv/MuDrkB5i2Fq2IL
zdt47mE9BM27ck+6gyECDn6oMAYrMmxHGudhZDvrzPt/CaPwYukQDONRKuq2f/bq
QysnDa+cqy5M/8f4mNxDO2yP2mB0KYWBgRYDrUoWSYEnpV8KleMP9SX09vMndzHk
RORTE090mVB582vgruV2N8p+2EcGpT8Vw0rvqqreMHFWcphgtlFVDfSdKmDuATpt
6WUPiOyV4kDoQywRNxP4ur9XfypCYMZ7xMr9dLM6cNnhu1TvfNI696CoVaIgSR7u
v/2Fd0+oXyUsbNwgBaa6HWswc7+dLznktnGlNyI+zeMx2N0eFSqkxpPUBkGj5886
oKDPDaXojYQCczvTSFMM9E2Hm8OeOzFkQVD9Uw4A3VNAPDL5AQHWXkJ+w/cqxuRV
0Q9C4U7GR6LOsa8CKBC9OvDbgGDHpdLsDHZOLDzUDk2ExdcFyDPCbmsawRHFnzAx
zsJZ3HNZBLd+yc5LhSga6H19gQ/XTJj0dJxjtFfbRtQavQYiS4LPYoK2cnFVHXmd
nPYjcp5iQcxSyeO/cF8n2ZzrrQEPEY86CKf3IqgOZhn3yKyelvEJsOM6qtzo9qhN
VgWCTT5pdvWHSimIYECqKNAmDGnja/AvECUhACyEi4euBNQXt5ZVIc1NUH3VHOF+
gJvaAyZ0Lc9XCvEKFGALNvktJdJ9KjQGvQKka2ImREU55aYQ/VNADnsNSeLAyMP3
TCR3iBQ6DYucFMUHPeXvFM8VJrM+R6uxBaqQG01ZowSn0aFSAUFXDSHMKJFLlXER
4cgsR2a5/UMICbTOTbLv/yrIHIBcQV9yZ2KYmLXsObwmKHAsx8wzKEMif9mtu9+i
W4TA/RVEnScio6KJVPG3ISTAdDd1mKNKMqVMT3vvwp8KIaH+f6jxfndV5sShBD39
Nf2dDNn2v0uNrlg7Ek2m79cQT1VW3S4aQ/6mWGFqY1Y9xMqZA/nBe6QZeyAUmU5J
JHNgqkMLHpWg4ExK0MwH0ZCXR/yo2oyjbr3mpkOtvzroI7oz4t6qz4JDNS8fttyB
hlcHXQm8411w/eXfkCIMsQCqcqAck3fybiXA+PbkrGTj6InWsQYTwH6r3G132IFE
VKhazM9u6xylPn9jAVgrmCg2SLujTEPPqcuMii4DqzWNS5Tv2wwJjeylfjYtOMKd
M8PcrJ/gQ7Ru/VtPibpoNkx1pYHRXmkOfomvAMRIuwUTACYb5JEBFIeT+YaovDD5
sR6zBkfpbc5Iw7giHH6RJu1SYJO82VSuWXntkdlfXoHA/tcRElpX+3Fp+FXHo7NP
WkmeZ2xLjggEsQS4+qmSuepv70myu0UrtbIc+MyIcOyxSlZNnNYwkZx+Slq52qBx
ZF3/moUEkBmpvd2zG3olnyA0+7ET2xg0vr7zC7tCVK5dhP+827jbCC9YEeX0nkRB
zKIXTX4y2yu4M+05AACDNZe+wwmvHK47SxR3SRQjIcfnS46h8IiVTOh3qGu2XPi4
u2HKavgw1CKh8uY3tve9bGQIgvuM8Y/FDJXEAIECMm0DyZ8Sf5ZZ3+8U1ympCzgF
lamxX8g15b5+duwNgAGmzSBitTaobEccJWWEtJI+NkW+3iGyXNH8uUh0M7ERVLq6
uQDd/qPixL515ZxGNpgZAS7ovTtYcSLme/K/HTYbEamWVi76XqYfgDK8YU9gLrw4
kLUZB7vXyZtWDuOFFpYXJ14n+y2A7TVJGsl/Zbh9mQ6KR9KRcAAXu0gFHPCoiDtt
eWLodr4+G+Xlc40sFKAyAG70GVBk9nJ/SHHHR92uw4dnWf4DXlWPFgpmoSKRbKWI
SK48zZ2IPex1Tdr/sfA3MlaWOSpGp77br8EPrdq4B8vZJy+9YlHdclkBymlQfc1j
P2KjeI2KCE0ETS9Y6ks4dw7aB/hjwxLqvYZy0IxkdJJlsieOGRpUqWFa4CBmNjme
H1f5X+gZbBbZ42GejCl+ryOWXloij1tdO8DcIJK7yfQNRM8oWRancrYBRIyixl17
ERIr56EjROqzptHC//6rtDdRzcuS9kEFE+jNKisbGXsKr1GtNWszqbpXciYQTeic
6OdOnsLc6Wyr5lBItFCNrRmJXQRJuPZQhurt1Jw8A+2Yu4X0/1XYdjzXPR446vCp
FgfkQeleGKUop6aNXOv0hZfFjIB7igKfsrtkh1ye/B729WEh/3vUkOASlOu+o/a/
foFuqQpg1qfSOAh6XSv3PgFz2lOGFxuKOkTNkNji0bfS/7xR8WHTf0JY017pPuox
ZR8aoQKP6kBq7b7HN3G3qdq04t9FHjo189rxfklCotjMJYtB8RN1RClRzc5S6zTa
TewwowaDKijBx6zSb1SCmTas5JhZLQcGIGxeVvOq5bLcitUZejhznaCNaW4kRCpV
L6xJ631eTyB8GbFzdt3BwPFsnIpD6SKYwYEd4z/mixNZRXlmnUcDsvt3GBo0R05U
I1MCpqGnFhnhDMoEFBlZiKVJIydZVAbhisx/9T7QhTk7tSKaFgynr7ho5FtGV0mI
7tuKk7Rwh3AMaiUoiZBlhfzFE9j4ggNGyq/oXdOHjORcIi+6mxYWjcj7YXaznOOm
HpI5UrepMpCeIxmRPEyLeWryACXsQVlk2tF4pPMgcEe41J+koGdhV8mBB5dd59qO
sE9mC35Ra0Jzl3swkrF1KN5zAXhI9lJ/w4Pt4py1Xd3TINnDiGT3yzOOpwTcuc59
4pXB0kiI4T+h1R7aguwzpECiTrfkcwzgNaPRYNaIkVfBWeHVDsI2vLRlRSeJrTZe
TRrNVyssaqxw2lwizsOzlHqyj7/sbFdRYvw4dAuhI899q24w0xMpBUxxabcuHas9
ZTaWSPoKD6Dru9UWsD8vRyn2PpXo1Q41eIIi2JQWHFiB7ILqdtorvAfV7CWIOfBC
6BkXGzvMTY2hW0EK6Omzka704J66gbjUyJ/DKB//O0bn/8jI15516YOhCGyAGSwn
sfbx0Hvnw3l9PCsJnWKUpamVCV8t9a98XPxMN2+5oFbih5d7n1j10qdnfAUYBB+g
HzWiRV79VzuEeVIJxxUSaNCdO/pG2fEq3iBd5SlMxNarZM0JwdxfwyDRMGEtrhJq
mti4O7JKd0/nWAP62YrO5L2BRIwViJGz6L1R9HzVwPdFK3oPyQvdwUs8X/CHo1tB
TgsRIH5K1qQNxM0wksrJhNVkalUrEKUV0wQVh6tCOhlDw3HChq8r1b0Cxr02tGfn
Mc40l9lm6oOPLRaqqBskFemCykx7OhVRdAiGYg4ER+c+vU0yh3UWnui977ShpgIN
mlkoEnm/RuE8kCG7YIn+iaZd5WW5+BMeWidMZk4sKSbLxDK35vx8dM0oI7jqWi49
8MlwmPh6feTftK+3RNYM2WjefzjjGeGPIMdIivs4YKq5z5jjlLkfQ+c4TUJgIFAf
B8Uw4psfbwGaNJLrgxi4qY06yw7/7gzvLEywI9L08LCkl2yTdO/9eZ8kv56xBtGl
HvZ0zfQjfR9vA80atLuVQ4P5V7DRMYr58cF16eXye1Nn0mGkwmVME4DqQ5jjRVrI
dAWhqeBpsEZaR0LREJvaraH8FRFn9T1DJRdxYR3HXChTpTq8ki8RMSWEN+spO22m
d54rlO5MUX302nGu3fLJaYD0/7VFvR8gQQB1MNFi64bBZvADsReOCjWqdXZVWUUv
NRSgDFGGAaGX0J9GF3ogXZcjWjzNyzDJGAwjALB8bCBIOETZu2sGLYMAfkAl01c5
MhWNiNBI76uKa/X40+OmCjtuZmcJBA7timXCwiB9rsLgJfqE086tKnpLl5WVr31P
6xEMW+WKvgrZ07bJ7Xc2jHgSUTCvUofGh76aJ4WD6Idj5P4GfXc9cVRDTfHhxDQX
jHGTb2wBR7dBI0LV/XfSPq0ixGnst+ABgY6b9XwoQ2+e9aE64dR6LWxi8p2UhklA
sdRTEYIgoPcMC/zXIrEMZ1W034mCcF89lLIt8II400RLarT2CWlva8djoQZR8UPp
Cn3UvE90SKfzboq0kFY93sS9wsME1Ie3WLUrFz7C086ULXRiggWTGYlP4PGh84+9
XHPCtm4zfjWxAXaG95HLvTc1o41oOTUCGJJVJPEWNnNtZ6KqtPeXD6/e3y5Ja8IZ
PvMn0Prqke+sL16HfK9y05Q9GD5Nk4TcRGK79IjVbUDaxrNvM8vOSlt+aKnAbmbV
oNT6Pyjxy5ukyLkCxYHcqNamvUFkU8b/n0yQehoxKf2DAN/clO2Itr7gGOyAZdQn
tBC/MAlqmdy30t4MlbZHvTxiGRU8RZT7WizbbJ8ZpZeIIvZf3AGD6tXdjqka7jh5
ulNlPsoYaLoupgMxJXxs5iGqpEFMngHlCLKDJkzH8nMVY/1DxwaaYKFS0YZyFUS9
50zhMbmW0TgdbpTZ1Ads4zY01iqjQUiskVXZAyQMZDD3MdRrRl428tNgH9iasRCR
ldDoNb4A6riM5gdqg0xsQiSH5tq392Rv20WnwSop5iqUWD5NmNDrmFMthz6xllQB
A9igfjvTCk/902oRGQ2mkiaVe65IM4zOU4F1Gu1bc9+pq/++laUAYMilBFXUPmhJ
VewZi33V+/SgIEXw6easRmSGrdOOJBO3bpHYa4nTAVP+hTQ9C0kn7DdWM8L0heiP
/+rccjUV9Y1Hs+s4fRJgswHQF1vkRIfdH9aRt9pBNYd9qrU9lN0Ux4x8Een+pgQ5
uH9MG5RkAZ5pkramKNKj4w7ucdfPX/YrhQ4CaqK44Pnutypy4G4EDRSJ5Jd3Od4Q
JWKN97CoIjDCQCoJ2mGHGILFaFV0WfxSd4Waf8dwN60wKtVEkcHV4ImPP7FfjpmZ
viJSi/yXYLlOsgGirorzZt86p48qzEVRlyvgwQBUORRDgLcGA9kkhPcUSw2LNi/a
EooQRG88GF5CFq7hD/7jRmYNLuOHRvCPuH2VmKvxNTHVLS6eA9FwXeaa9o5xrB04
KRCcKF3dUjIYEas7D71u5oFf6ERFVFdLvzNY3EVt2XwNrm353RDNTfpXfDDYu16E
IM2DlaUkBhIpvrb5cTvl/lN+wNTc2TWpvIGtgOJbO34KQagrTVG/BAGJoUjZorkX
/2oNv8kwxrh8XdE96E5Jx3J8r6yHgL9At5hohmO+pu/rwKYHQdW4wbdBFRcs6EP+
sfvXnYhM0HliLwVyHATZYKX2+pe9bnkZZ/uB4BEEE+HWa8VI3pGQf0V7rLna0y6u
DO+aQSf9VX6MbFLdyft7C9XS+uUIJcdnSTHfiy8HnoPTVVDl9YOPqkhQ0VpjNmoR
hzljf1y9RDZwhP+7HehBRWaaO0BxL9YsszJbqaoE3FEXHkFHa9kPEjjR5+m4dY3s
5/EtM82Resb8GJKhaUYciN3a+zRUwPnDlqxbZCnQG5Uc37U5jAiis2XAxrnyqPLx
lkn28klYUNJx86gn06ktguvwN0iSER+HM09ocGg3BkAWARZM+UunJnTU9T/nry+r
GmIoIyQmpikYG49oGKeDkhc4A9mP6ZdLghD8EUGc2e45fRZ01sBabURDxRvnQDF6
3QaNnfy/6guSQ2QJms8QOWNDC7e8klyk1PcUUPqv5XNf24of+PUdb1/7d0+2MGtz
nqS/uHXkdWQM6A7yMAUb9lAPvDPf4ph/+pGfet89J4jxtvdwiDjmHvL4n5ckQTlp
VlOt4/MOnMeXdOLe0xjLA8EZXAxN6yq5/oExtkH1HSF4kx0Zg8EBxvFTehM0IdyY
lDw4Qy9YmEVLfpOINLlmDi1EhG1vDM3lEZL/lF/oo5+bAtW/oTjOFlbmlNlZ6w3a
tuVIX7ebLAmOhzhHi69gclZBCpHaaYhOBoTTWfEBWB/E9Zr9GYKtK32gln2sQXcI
BgTAuC7dS93xHyA1ZbSFmPNIEAwfbO4MK/cxAihZN7yVg0I93sNtF1vWAStsa5B2
nQmpoyBTeRvY/ZBT/yPvVTFs+h++zsSNtNvghLCdiA2U91zwjSNBqmQED5N1Vqqb
fGULJbHmof1SvBYUTUfdffX6FkKE0wo0vEta13ImQOVVsMznhoodUxdSfF34bnLU
9gmYZBCGCVZSdsh0sx+5MyDb7VsayZF9dG0+d51zZW21If8se8D1FZkI1G34Qh/Z
5EAxVr+LUpDWve/QhivhbZKxeBxVLfGiCPy/NBbO9c12tcfE7EMpMsuhErGkPwTs
agNJa1MA+jzwkGv7y99EEYcUu1EdWOmAiutpXatYJilgmWHFoj/TuI+KoLwh3zJ1
YNT5sBnfVl3PR3/GiWZ071POliFNsTf7HvdWPsrz/E+5tSygb8SctQWh7QiWEvAP
yp5BymyN6dtEXHtUjDCD0mvG/zvXw2ZYt+4ejHw+S4oC2gF5ymdzHGPOC3FvRyZ7
9eSjE5BtZO/SJxB/th0xQnNsW1e1WG2jgfZhkEfJ35cV6REAfPTANVsvO+ePH1Tw
A8KNzdVnHgLylTE+9zPO8RnmQR4HyVkNkT/8DvCnsElaJgOUUoaOiTnsT+Lbkpqq
BKE70g+8Z9+R99cF48txPIFdJPRiSpnLzhc+Njfs0utp7snWJ6qlxo9Zrk+16hI6
qnXjN4wf+f5l2sY54Rx4ah+Xvbm8ktLNl+okzix01y2lGABXZzcysxQDEHVkA063
gLFNR6D/nb23KaoYP/MWJSezW/F51oRkqg7fWcupxyDipwQdEUec99G5o5h0zTor
oukhTKHt24ZARpUZAHoDm82V2oWOt3L/5uyM4SHdeorCqB2NCZHNAzPKm7yuTzYS
S3VUOXVz/87OWhW04LeVh5Y2LTiqQUzVQoDxMwPCV5txvb1ibIvdzlMlq8or2AK+
I4RcHKow3gH6RcksQAQ0xUhYAy7zRKUHtfaGWekM2JHtXJ2WTrp5rMqijguWxoEF
iPNAMeN2kUa5ELNubHSXJ6pCYlk+/BohyDA21cDdVgdQEmjnr90W1lAEqpXkyc9V
y92t8QCzdCoI6M2CZCRHWBA9236e1oEndA+lOLK/aSbY8g6KO+FvPE4RCAJEvbz4
Dv017ciImlcouM9aoj8hgVzfwLPfChmjiFdwPUhgjQtvJaBYeEES9iZMC8H8Qza/
Tss0oeuR0CuQV205guW3pfyzFn5UyrhfeCKZzMWQ3Au+WE7SmCXEJZZUbpa4fpuo
4SJMgBzTWBVzj2d2gNXtbW0fHYuqKGDskU1jyQdJzr2yVxQbZhSBhhE0x/GcegWT
fwNvGizgs/Tb9bq7KvusDWtuSxEVd7lFIIJbIPj8XCuI7PALt3nGlZ207GEHrG46
gcv1yvTQ5TwFqUq0jRt4H4lNkqjCJpwHGJs3mPKMAcqdIdueLJ8h1OKJtkYRL7yO
IUb6Rexb5p/NMuSC1unT9oDkm80YL+iBsiurIbc3sT7sX/L+ESRTWkzLeyvVs44m
7M1V3YI3pEunWyl569ak4wuEBlVOjuSC1iwoKpLIgeXQ0mmQS7HIOMwVmMEhsVS+
OhjxE/PQeGA1tFAED6kxztO7hSkZsFDgPJn8rKWhe4QIgAyTYovDavy1T3s9Mphr
5zC+bUjishDuw1fJ49uXiAX88dnbOGYT8bhke/Q9Rnvy4oqNpw6oJ4BQ/c7eeSWX
WEXoGcvAFVgAFde6/uwFojtXJc9rTMEj3vgYJRKxpfYezujTf/8ekQszH5BLTbEs
bePZkSULh5rWBpfsjdWFGCcJ83mhLXFMWA15ZXey37/frkKxBr9SwOgBverYQ3sP
otoMzWuMZCl16JD2+G7I7kLqUXnbYhj92wuRDs2uYEphZnjmhMOpVkRL/Sq17yqF
6Ad5UX8iH7ug3rZkQq8aMc77tDbCi9yetk++EEkNxbdvB4Q3FNRk0mudui/8Zmx9
AHYBd018NhS9Ju7F1lm3liw7sW8RNOydvJjoGjFH7r8UNvQ0K41kNqm4iB0Ls2CA
MLmK6gOlVHMe6ubeVjrSN1RqTOxF4MEMDuUjaX5tY9jQc2K7EiPxibppg1KK0hPq
dexfAN8nx1pcOsvbImV4ritQu+n20ZbawdVnQShm759seF7sbY2QmyquDepl5i5q
+XjjnayWB2c1eHdmm4NyUknYNg9Rc7yoyVOndtzOCZ8SxAQ5WeYyyhByUj6MVRba
3R3or212OvtqKxHDTihlT2lYihFk9+BrN0C8uWltj+2+uyootQEguSLw6X3rJJHG
s6PK/8P/3VeGX2dupKccwN1SWWRT7KeQpG3Go+HOjM2YCc/NzerLu+agjykfGLPE
VmDenKqW+uy5rnusfMlKoyIpZlyD12iZkDUa3KtPcmi8jqtW5U+4fuox5WCWbG7W
d60Pl5UsDC7crVEJ6KrfTsgwYAYvsXZVmbeQIDaQfQzvQt388/H0D83PHWt9y1Fb
Q9O/0VtpfodzkwzGAaf1ESngOkoHMa9RXMuQl2KiySiRM6XuPlQHMQyS/0l4ltKz
UxCQ+MOtsuh8Zszc7qpQ9f65rAjlXE8wU5JbifVwjvGiSsAsfLDyNtkk3f0rVsqe
8O+2o3gbfU4aI4LsPEDUgcM9/usgYpgeg+tvBVe5M0jj2KFa56BmDW6lEo+eSTqZ
qvHhB/4xxPpxYUHXw9V83vifAap87orJvSgGEpStl0QH+D9ZI9KqfNWQKRhpUIY1
CySw0X7AD+38fUd3c+Ju9D3YECbjp48+evDspw1a+bxbSgAJVhzFII7ekUbppF+6
EJNARYxFwx202UlSXRK8bhkHpT9LDRholAR2R3We2q5XCnTDii+CQ373VqzftkCo
863IX1a6IuuuUzf0wid91tMimAyCYFwIQpDcnCy/kNT+00GKHbWXvTqsEWWTZB/P
v8xQJadjdIb7WkS4hoe2CgtFZEQhAgW3sIb+t+qsfiij+u9v4iCEuJpBrLMOEYWF
Bw5Kqf62K1OQl9byZmf+pDmmvmmVr377cGZpSz04uUyP+ioAABEysbZ8EYbDFmw0
CTtPPvcZMRf12ZTsWkcKdqaKU40SW4n8JZD+CkINV0TutgBP5v2jy24ZXGJzN5Id
nWRJg8bMIAHPfZdjiNndpVEWM34myRlWq1CSsvU+eMBVGvYzBvPXLlVvpPVTV+dh
Jnlkr+NquOBRodjvgL/zYDsA9OZSzO0S3ItdU+yi0/t5GDXZ4/V8hl9Ck+GuyLvP
lR3vaqjSxkJehn+3fKLJMdxAmImASpFZgTz8FNXBS2ndri9C5ZJLPoGIOUP0GpHy
zwacFtsWuUms6ShLizcnlJT4jr2vrpzRSUrAC/DipHOGjLx7zv4VO6wZp7LWI8Lh
KIGKppJkS8+bIt+m0sOfuSd0qfUmJ8SRAaM9rfNj2yNnsCBbTMWdQntWAUGpSOG0
0ZiNqsP9OFIytjs4obwkZds4RLLeFzKwEiMJvzsuIyE4zDLeyZM1NfDD4lw88VL+
xJBdxCJUvb3ElsQffN8DNpBt4q1WHneNKsUfC1g0/GN4X7Dk9RGPN7uR+0DYB9IS
j/b0QKRGUJI6oPTTWqlrhNdVaNUz+p4O3MDZaLbx/kjPLynVNnFEqPhKbI4ZRkn2
GsSStS8XsmrqvmJTWu2y3tAJGtMgruXOSi0i1WO4iwPLpU4F1lFcMDjG8sw2uWN4
pyA6QrdneC0KovPqe7oQUQBt/k3JrMljaQP/nqB7fr03HUZQXaX4B90Hw38RmGoE
oAFmgHlhUbY//EuB5WFGIgRTADseFnorbcEHMgtqIa3MoaxOhTgZVbXy/32LHD3E
TpOwLZVObgmLS7FD58Q7la65xdSNzAAh6qovS8UliOkNbIXjlGqj/INZ5CePuGXK
Wldip5wbLzU4meOSQx3dy1+Lok07BgG7SdN2QXppwLwo3L5rAJjbpaCsyRtu9PIq
T1WDibkC1bfwetb02ZnE1ZEeWMIP1C4XZ9Vo1g9DHnGKKOLD9V4I5K5k6F81SZa5
mRK5aAAZG1yPSNsFiNRY92ysYzKcM+D6lzkGfU8m6GCwRjsP60h5+QqQC64tclfD
tqG8PVXaxacRMo6Z08DToO0qwmkhywN6/7EZ9+Krh7HbLyJdbHwMfyughHGp/5kO
3qTYvh7G4hjPqaOIDmpPWhlp+0PcEkBY9nMcb9uQRn7Z382uiaQmczaBikDuYqFZ
afVBzvasZ8/GdeGHfeKRSxIMcgBHOPT5u4u0LwT9tORhV2HizrlqPhxh+9m1plyN
qhIYeRK0wXnnwNbhWXxsqxY1ej7yIFOsnRUdCEcaDbCvLMggsQpFqBjpSChNkUD5
WD+4HP3NSAsGqkYi8E02Tl9tTqtzAevR7zaiBByaChVSqO3UUnB7hNBWmlwkRVg5
vE4rBXQ8xwQwXaQE2hBfuUnbCONEL5/S9GC+uMDU0R5c7edN3F7CEr061G6hne/9
3tROOg37h9vNBZUzUVQ7rAmZwK9egnYxL0oHxCJAtK9HESSOdvuPhT9bPW+F8hrv
KL8TEaGYS3+Bkty4tLqUTH3HggMCRSpgcFv/n9ONNf5nMWGucxYUkOi4eCjwDwWS
1xTJiEEoZPUGZn87MB1U2dN5KcCMz6wV4gwzz117llaZWrUd2F8kvmCuLUyziYBF
QIJCFcU0YO73vmR4xzuV7b0Y6+yv10L94/sBOA6LZ9H05EXjFxYaISai6RWgtazb
peym3Fdpla88AZO+iGGJiLJLIjiqKmC1f2MG7KkkqNCpeqlJPPveQYN2p+hg95CN
z4piPw4y1OyymZWWmHxxEb9muCwIE41HsWWJCZSNJEyG5PmBHjS8Ty2jxMXBInQm
sijDei8c/OcLMB2ogBmwQC2fChu966LpW8TporWTuuoX8XQc++lo4DZuk+70jD1y
Ms0dsvQ0L+MYWIoLq7jzDhrJsvRjpfYozVgS2XeHvfDs8XbyyKxG3EAur60XUjh5
NDyc+JVF+Sd+DTfoSXj70FZ9318/AF495X7ZKqZiyA7gzx9fbZGSno+Dt9yp2B/Y
BPAfjrzo7xC1dtOvd9AYuKv7O8+QScLtSgmvzK6N3Nyowq25OMv9ZtsGNKsBprEm
AM0DZmPpzZp1tvwBQbs2b7B/fsIQjHYXJyAJX9NVaa0WvNZ2JQrAvd29Yr9nJLSB
Xjrsj+V8XvBY1Hj+uHhVR5roq6F9aRHlGSevS0O2rffyx3CB7f7lbKGxde4cQXu7
V1DL78XW2g5XyQ5xrCkjqmycBX9Ubk6Johzdb7ScIwMEjxyN2qewhUXASuuK9hJG
UPUcEMzAQfh6H1GqZO+dAR2Qzic82hiakiO/lHvo40qMFQLVzMnfrIQBx2JWjC1e
a9iKMCf1F1C/3BD03ypfLWMTGHLo3EcZ167pV2FiUoAAwpx+UoLzE4loSBStkIvc
aDr7N4RPIsh0lRGXHFL5bJoGyJKVg0mW+xpJnM15z2qOt19F4h5407bqoqsINmH9
vc1ocC3/bj+o8e1E8VPIwu55k42Ke+3BtpIrrX1GrkhdkjhXUPbZBuTJiarO0i1w
ojAIdOQ0ahV5n00/F2fYz+icIB+kEY5BGYeHl5OdK81GAdYjTEN0rtdETkJX0n5l
n6Sbs2SMQHAxwsni+NMZtbdUY6RqPknwLWjE7SQpAQK10KTNbFDXeNTqsamfygBK
sVr8VS/dbKYK+pbULCou0NSUp0m942t38Itf7M12IQ+lNyZy9k0XFIgIzIZMgA1V
TOeG6zDRzAj/Eu2N43jZUf32iw+jr5xSLhlYM+/FfWZoVI/+yDmuJKXLExIBjwjP
+FByuozNbbWTA+WppuLLmTQvkWOR6MkeTc6VbbnQANke7xHXPNUdP3VNv7cU4JRK
IUgEeOrlPEOvf5tmvod7CPlZoPBcCjE1IkEI/hDvGh43yOpij1Q35X0gYyerpvYH
tbRsr30R6+QfImJ0mSykt4hsBjd9WXtCkbumk9E4U26WjrFg5umisVbOijixmxda
baRV6rGjHJR7w6UB3bk91qmwvc1oizL1fT9xYv8hAeJSFRpV5xkGkkEvvTmiUoBj
8ay7xjiw7L7aYdwphrifYEbupg2bOc312j3puodVul8VY4kRXzUaEvxGh6/yLfkY
3tr9GCrnVO1pAOFBqa09JwGLma5YmHKtREIp1QP3rB+wpxudWPx5Rjq4LYQR81gi
et4BAjGT8w3zO4s+NA9IwpDWaXEj2EEfcb1vVqb7qpcY/sJBPIMWY52bML7J0bJV
E9sK3qLAzntTtTX/xbdXbvOm2PP2kUQ+YAaXS4LdHMb+nFMBQIyNWOv7nSVg5ywg
6FRyYqXfuUO/KYdI/zynBXFBCPyDgIBKkhvJ3qozhSAygWn1ubueWRZUfV5EiSAW
ftOcgqS0C8Yxz14NQ8KSfZPQmvYG8EEiRJ/u8jm/ydVDxc9orR8Vm+vOorveavoC
Vxf8xtvG+tfODPNajHUG6htkrPmGIq+wCUH3cy7pGTBZkalCewrtW5MhQw5p14VJ
b9qa1pkh6lC1VOippDFLe/hB0464DLIQIKSHRSnkewX8oKlpUhcWjFawc+1Ke+Mw
To2ztxcCmS08sCx/AdA75U7WTLXYdaoTjEXlqXW/vQTWbMlzEJNkWS+4TsxsD5QM
VfJPLVY5kzd72rFXnxRKppH41GIYkNJlOWEDJlRFbx4mcU5h1jZFOD5A2fvIi32f
D0TbM7Ipk7MOuXVDMk/BJc3kBbBXY2JGh+2elg4XHaIzkBhc0LU1bTpDE+1U2WbG
FNvhUjH2DJb/p5UE/RZoXhZAEtL8ZX+uZP34zChnwEZVLAgRUHCqD0NNhnIfhulj
atmLnu6tDngZ8X0VIP1BohtpRFJbemEFYUF+Um41JrCK848TkCTo1VJBNzwltexA
5a1q8oaxm0b7areBSwAGLdmuGzmioBx26ky35jtZmKMVAuop4degvnrDSacjhCbV
pN0andWTWLLM2ognOQ17W8u9BuEZPY1VchHMJxUcMMvLys+gK1tL33Ko+YLG8G6D
T1kGUruDyv+L1S09kU/0SUjkGpDvpdxWVke8CMIBsvk96+6LaUOWi1JsxlgBBrV/
1/nHBT2Y9Pq+OBkVsOrEBSTyv1f+TWRO6vfqxzrbeOYa/LKxfIzP6GKQYTCG9Rii
qof1Smuz49G8sOK8PYnGllA5aYTAto7Lf4Sojf0LEEEe8aCw+TM9A4njK2Odz4Jf
1PSimnIPhW0SJhF7vrb+lcOXKxPJFAdCW2cF9mdKaCYXK6gRbokaJ/1Q2aHQYQv7
tuqW8vigOrCRj7EJ1eWWgQgBOEBUlF+v8G4+D75gPQw0a8k4A8ov1rIy7vfdIsJf
4wMjpUZlJAWagD4RyMNoobp/9hE/4oB6/+K/z+MDjfa+xgQVtD16bnTcoYKunJVl
eWzCBziOzfFQ6jNJAbbcMnQ55nTxF/udOtkdba1aTVSHuwrHYbyM3I3WL/oATqeS
UMywCfdkdmHuo/6d++eC8bjAAfajP7oQaD5kt2JGvBP9tSOtmefdQdc0yI08H+f+
0h0gGmmdyauyOpQZlfDKwExvwaCDqyV3FqlbiBCVxOntzBNBActf2WOqgMQHEp8s
zC4zcEQBZTOLUK/ZELsV7WPOwjywH0fgbVN2HE9B6N8wsrgSKaqshh4xurppEEzn
+O4LHI9F+PG8WQsnL7RQVpugB3aRxPxsbEyTykjyejaS9NwcZOoU40rI4B5EONJd
YnpeHvFAsNjVA4Qu1fBOiS7LK3qeLyrqHLlx1v7cpchndlUlQ6ijSeQ8zZ5p8jok
/jVekCYeUu8GFlpMxjvFYOEji1DxG0ioq7Z9zB2CnVsi/za36gfZidnmQXENUTXe
LDSdsyiKW0NPPZq3BJHpr21D7IpZldWSuyB5LZp3bsXzNF7OedYkHybskuoijfLQ
SDku51QNWnkY31svGqp1xASuUd0+yuQWDxIY5t1uGeqxoAhmUeIc75l0sraldm3F
uhagtep5ADk4Ys8VmmMt977DwjBXjnG5XfnetAbFcjt4U6rlpao+ovuQjO92tYGp
W2CdRA9sygcNhTLX2yTJxKMcR4v9f44iFUX/6KLU4vs80/+nnnFQ1ujL2Wn4hdX+
2eYIOw1qDMZpI5IFw1zDs02qEeCpjnONTNInwyorK5av36w783c69IvD+BgMCzdL
B/8Ulr0jn9Yk4IT/1tfMqFTocAB15ncQ8/5RcW+xggBd53GPg2X6xVeyDijegviy
NO7KhEao41pW7Sdf/4HPpmmSj0FPI24WMgPPhpjAY/PLyBsW3QwL38F0M1yjTltl
73Tvp36dDO03Z1wAs74xlmKY5zSHRFo20bAnzkfA9wHgR6Urqt2WOnMErsJgBrXh
OMLQhKq4NRem6uoGoocse/6XvHRiJhUazuy+Wz/BlCNiMTpMBRqMhSUsxNRmNTki
tAVN1iBZyF9+E3EzW7up5hs1m0W/ELnBCWnBxFPutgYBD/czDYHflPPBHBYPiFMp
L/AwnjLURXqT8I1TEAS8s0ECEJ8I1Jnj0ygMM0bnmBz8+0KAk3nZkn4jNu3X7l00
df/4mcAR3AHyd7htqNtXH+Snp5cDUhYN/rddPOlLojC9eMxoOZb7cyezXA/iBmw6
43PMHfiDpV1EzUYQZ5dBTQ5TmYcr6d3IwMjxve5OVja/oE1VCogBSUIhD03kl2qb
IgxnyeNEya+MDd9qZSAuv9InkuvcGdtXGV2WQV7MChG0yHbHfXttHE7S9LPHIn7K
YON0AwW8sFYaoyzpSSYlugCTK1alUWhUmPsir2khSamnyfEOcI/KOaxy35sQ8j0t
IJdwbbG4JX4VFGdQpFFZD3zNaNJ49FDCbwm+vbKdzo9B2NKBrn1J/QkAJlW9GLM0
iLDB9nkJOFY0IYhuBtAcQoT/s7dyHdSyvOD2yUQXT3D1tsLOlEh/IABmhq0fYVAe
jTlbq4Xg8Ns71BgR6aaI2oIDlZa6vsKpY/TceM0j+iz24oUse6POTRGBY1rXRMQY
spy1KyfgC0a3Iytelbfx/FbRAb258Vb5c45+bB7SEKwkfTz5cx4NOnlxApQXGoEy
iJyHLeS332yYDy8KbxNmvcN/hWJlGcCJf0lz8lOQuXCqw3kQ+3nsV1bQM67NggeR
gMxmAH3vFtRysSNLXInaK/+kx3JiaqDoj6zUQ2lc5yjH3Ut6sxOGbW1LMdJP31O6
NST+mh+xbhY+ZqVdWGEYQnibCg4ZmSJXOPQIgnCvZmHMKPkm/QuhWc4CjSFWzKuB
ahxv8dSi9pu68mKCO8eLn9/wU631MuO43D3xjESwhirCmsgaY7Swt6Dx7jJQphuw
FOeeGIO4I09GLNdA7Po7HP80rx3ZgSwEy61witzxcejyrIGto1t7gta5PYoXbSZ4
mZcqitOJ4b6qoPK0xHriTKdzUueY0SyxA+WV233oXN54MOjBV0wHDb6drgdT6NMt
HUvSUHv4cYZj/ZWrwCS4dfWLHRFAU8oEE4mi0a8+K4RsTWdQ+DflkEBBY7atpfJd
ATRaR4lGpK+DpugshkqJPDfy/crajEjfiJnsRjECXdBhp26pWFkvYG2SuzdBTMb6
P0gooGUpaGfG12BaTIbmGmLp6WV7aG685VmH5868g9uVlppT0dGWvT5fuvgkjX7H
0qVip6ux7m5NJ1jNi/CKcNyz1FJ0CUs4Ajdj1Jm0D04IVYtVzg2mhfoYks+amcZo
3I6tdNJpPxr/STHlWD9+DyBJNHt5c1phkFdGJ/kCgxBnlM6q6Ifew+3vfw/+nmC+
CJAClMNLaDfPUjHOlkUhHepvXhPRRmeA4ghrV712evVIHeuOuFXA1BDnv58cIT53
9lvVqtTF1njCNxqIi8QSZk8x7/QOKoxq/TZzg/jhth2gvhLjGtuZdGG79MBPck4l
qYjUEQMZNwljUBY5ZX+ovxKlAPUnCdn1E+GGiaHly8aoHLj3R8Yo0CU88avWQI66
Y0Pibt2fZKoclOPiVO7D2WXASgOtfAyzroQv5OpuJJzqA/JImj6GcghesrpuT44g
HR5AQPMwl43IOWueFmS74oTBOgql0iUp6VsDDrjOf7FhQ3V1WVnNMhVs03nTeMh4
q1z2RX6u3K+nCMfZCHBy860/WlnJLTBNjvcTJm/rMl8yOBr3oKDV5dTko4yq6+Wz
oztO578U+1RPw9DVWsr0Yo4h1pVg9P1XCtEnvnnKLLWoI3s9WIPQ1z5UXHTPaiv1
Zoue5/NIQruVm8Ssw2400bwx3buBekfZZE/yqbUlXnHZ59aKz1vICmXQjApmwicD
xjxgN5H4P/c0kELDhkfCbwJa3FkYoMY6NL18zFGIJ0EVpFPvdrhnDpJKHLVoEu12
MZLEegkxG+UW6Vf3/c1thILTDTt5ZWCG1/O4IM2/KgCkFVTCzcmaGdjwsAXA65Or
frLQNnlBC4y/yKa6tF+nTqFrwBe5HVGpUhkT5Uiic/q1vYjWu9RCBnE/RmGus/Fk
N9EELPYjzawCik0LkaeeKtr/IWu/lzd6AZ7xRIGATSScXXYUIDCeOZU8fMvDtT77
I8tB/h7GvuaWcPH6snmKx1DjNvVQCuGUOq3V3ITSLdmwXmxoO+3nH5o3j+Cac7RG
quTkUa4QFKEJqxy8Jw0B3tJDedKwyQJzRfhpLn5twggTZWqKQQ/0F7nBHnILo6ui
tqLCxhfnR1PHd/OQPyHaxQOjPoQXszHggRLHTc9TgM3nGQ5Qt/rauVVRsm3muymY
UxI1oJcWv90QrR7g4/tCyvEyBjq9dBjTWsrFhtfXw3WDKxwxsHUGbFgszO2RNhzd
VPkp/0E48Q4wVCZ1s0NbtvjFvj26mZ+49FOdoaKPXB/yUJCUA6UmDgipT13No6wW
RLFdlLWIe8Vm7WhnZmQ7OBW0zt2X97WrTnhBFJDozV6sxzyNicF1XjVyiW9a3n1c
otFPp5fvqXSCn0l3lW79+ADPAnjuYzlWPLLVtQfks3SrQxP6RTIeFmVmrw8ToyPf
sOjGrdWgctYnKlkONWuoHtoD1iHwEPeADlv0vTIIHC4Qr8Or+PDRplWu37bNZMye
MX0pdGo5gF3xvpovtJhezLMiSJIdw93eSQmVtkmeW0G0wMBtdvz+IOTMHFUYaY9M
MLvWa16ghqj+gjwKKf1ztJeWB60HLTJvUMXJVFRRLg4Xeh/AQTzy2knUwisWfCHV
QxoHLGYbKL+TUQF4QiqheK6lg3GbQCkthNcg5tgIzazLn9s6fsHVuC3uvGbrW0Qg
6ilPBYO/vb7FFW/kl2cWTZ06klEmDIRam+0JR4KMheYbwZ9+Us3YQkxppho0EeoN
C97DRe1ucR2/RcnKSpq+hCwXE+mMgxyV2YkqRtE0Z65yQ4L5y2W6jOXJiqgZjk7D
27V/An5YRupMlZMfcUMXMlq2HDqyGuId9THEOGSn4eRc1h5Amfs7FLSpI8Wa3aW6
Gi/EviJ7WHCU6iJMf6x7SQPGQpu4guhhMDu/v18j7AqO5LkCd9X+gyt9N2SftzCS
/X+BxhsH4FnxPGJPuB8hZOnM3QRMHzCw9RphuskRnx1u+s//CPVHUgGRvToI/GRg
LLYwdsUQk4xYyZlY+/1z2vN5d9JGNKuGaNACTtwojwRJxsDXbBdTKihG/ez3EcCP
JF494oo1uckaMCD6NyAZREwkf/eDrY2uT7RTLumlErbjYKUx2gSM9G9F0l6QT2Ke
qzxvrAWOyCKIjfZbIU9vN1GN5rxqmPBztSFndZR2FZ3dC5fQ+3d57FK2CDZA8G3H
bLZ+/OQ3I58+fBj0GnztXQtxvHNjkxEh+QJej6dyKwdjxNAd5IqLiTolJfsc2LCv
LCoOysIw0a/DyyjaQOdKbkODdJknMUAxfHfKKNSogHOYV+kkRFH0HVmLp0bBL9aW
+QKgu8BjKi9+/dqJZ4MWbXoNKxxc/36J5bG0HpX3Alx08F+LGn7CsGe22EYyykGz
TRJkUOmpkF4cpjC6Q6bnx0kNvYjRXO4t/JObZ49bCT0zbrKIYzoyXF3fqO4d6ULq
VMrUl1vo4TUcqeQ2EF0xUU3rT4/BTaiuQShzyne0iCqh3F6IKwhWUJL2+LCk5w/a
kMiVs7M4cyYJLYiZAJ68gXlLJ5iDcpTwzyhLlYOJ8MnGGoB0rkIqH0QMcHlb3YP0
b7/xpNNHmEIbZhHRUWEXqfwGWITTNGfFY1GgDBdg4q/yWejC1/snyQtyWKYSvGhi
878pCunphhIwgGUTZirI8LQmtufDt7xlJ2RaujL6in5saQ6UOG8LAdmRgHY5IVBe
2+8lJMhgtgVlyHU0QL4Rwz2w03qzNzz/Kshph3qynjiKvuO+mKdMCEk0biX4Gezd
WEr7zf9s1P/4VrpOs23KDvQI1oUze31BG+me6IyJvG52PGywFheOVdLvVclKa5h4
Dkgaxt5WAdkBs8VvDKd/ZkoYaidEA20741+4ag1uLrDmBx4mxDSO3S8Hf4sQDJdq
TlKrQRdA+y/iUaUrlElxeXV9lRE0BRk3JpVKICGeQ4V8g3Qbpy7R0G8PJdI3QIDd
PRSNB7Xlhu2Ltx5UopKBI3n9m0+6iaF9JOBaEgfi1QSXjUHELE990kSY6Gro76xb
2Pctg7IoqPIVGtRlRtJn4PAf9xVox8VfNalFz/6QC72IqVhHJIs3EoRnCqZZgAPY
Zobwx2v5Z6cQXVPRsROCDU1NTh5f3GXdjjRWl0wTWi82kURIR1Gg8M+4tSDQCS7b
Ku8cfQRgRYKUtJSFs2fza3Rwd4NltRLyP4st86aDmGIXLgPu8ZdNkH7fXA6GapZs
TD15KM/sBy+JssYR0AUZe3z21tEcVh0gY0tSf9Ffyt/4bcbxvh/yL/3GV7s3EZWi
ysagJzwWUl5WgsArZodEkLPyougdTlSQmzEG7an/0kjNGW9U1xPuRsHUz0rzfdbL
EacDAs9PZGOOrdFzQDkHuq6zDPx4qtg6NFr1HhGCemxDkJD/zdly9FmkcMExsyZs
UROo2n1pIxUV8t8QArhpg1RX2vk0+WQqOo4DRxI3fgG91kQwAT5Nsey9EAPnHJkA
fS4gQjkgpWe5PaVANmrUrv/ZWDGppHLueyJ8+pUBVEvObPyZEyEVIB/ms3Gs+UsQ
/mMUU41w3502L70Ry4533Jlio6WBL38WkbdhlaP2u9ok4y1BIubHXg1ELhuWAQxx
K7D2kolN3np9CRIsrEIEkxpnSzqQ4Gwom+ks+A0Fx3g4hs6VCiWd1HE+D6pPInXq
89htn7M3mCEQuobu2H346aHdZNcfOmNuURHtrhy2eRNcw7Q5ToIasrOMNyX0a5Kc
mZHbW0C+eAUunrXjaOnoZRvJy7e78/jBkKmRoj6G6aHFAEGVrRq0T2LQh9X0q1mq
Ub49SS12xutRRSp3ImSSL6f3ilblq7WsYQwnQvOJNC0k7QCjhjRYfAuIdvEZdpYk
yyFtRWR7OBXjpPrN/uwoBsNUqNhKlZzZZXDEqM/22E7EUd3y1LPOSJTPvUtOjO2j
z9lX8PKtYmJh6w0VBv3YGYQONaLyuFy5mr31sy3RqCypUyv82A0JZ03SGEKsqaca
e8W3tFtIr75koQVrEuS8qnwQ10aKV59tyiG1Vkto9nDK66wWUU/OvUicdry7RmSF
g3VxvPx9mpMrak8QU2ohgYM22n95kTAzajPCHcZXVMe2n0ZOwUJG+G9sXgK+EwUW
+vUYbi9yMySlYQdP79CAS5gt8oJQseGhyQQuAbzcKLtec2ZEOKP5x8OjrC+8p8BL
wH6TnW8kl73X/6ww43phQnZQdTVkfpMmDiV45Z3lXcm6ogCgJAEtTVE/3KV53joB
yR6Ube+KXTpuLBRDvAt6eqNnHLltA0xw9q1KQLAI/3plFCRKlROCA4tOnxQ1cOY3
fV7CQoc6JSVPTr3dKJiuss101WsVX8vMowXE9k46Yrv/0HK6AQId9ygnEvu/Npze
GaCVqzKna+CID/p5HsmsDAqvOu/AmlgY2Oi8wbCyPHrBZTLG2h2blBpceh8cUVis
yoXTSxm1xWnR3gfTZO6814PLtMesGe9ZOXeGX8a6HdUS6GIt8eHPvgV4j5SfzmyR
gTX8chcbA+s1zYwZqNAe99iKmH+xjdh1uzi1Vve/bxh2d/+ft7JIsT+xBEFDcza5
N9YgG3919+bEmIMNfDQzrnRgFeqpLmNBEoZYhcPC3AD8WwDSNG1QHbEIr1+2VLMQ
ZYH3RmnFya/SFu77iQJETIrgbzP0PEfNEk1o5JPbZEslKpeWO4PR5uFHZ39TcLRb
EOeMzBY6TfrlXkF/FfzVE5VROUIh7SFv8SKxHS2KXfMVfCLwUbYPdTrh4qKW0P/P
ftB/sVCH0PUNKLngIDVD3wAjx5QH/tfCJrkKDvBOkaUOu6cbjgbg30L++LjIVm5U
0cUzV6AWoTMrf1lNUyvmEeC9JqJOtNsWap6x5NFthrD5iwj0xqj8Ij/PTLIS8jJH
bVDUQtOXiAZwxlCd58Oa6NRbBkSZB7+zAy7wbweSZwZVXEJEza76LQ9skm1jp9TD
8wExx9V/OquYYDKcfnN2+e5LLfld7JPbcNSoWbc/14FO6vEVVZlVe+1Lo2V2UQn6
ynA6KZQ0n1WxlgFSFH42ELGXidqUcOK2xPiIMsL3t/ITXIsEKRxOS2u6TIjSVbun
RhGKxYwgIr43tmL5C091yK8DvdX2MXiyI5WOntrMdQMPyEioFEqM8+ZuLP/67+Q0
olskzIqh2zJ2prCyY+yc5YuXf0Cei9DnCM5mauS0QkMnS5McWu5uzfY9El29wACI
P2Wcd1xfO7SFYfWgx6f7AC8iR3aIqyxmH6H4ILkc+G3EXrYhi/OeCTwUW4TLOPbv
KSHwEi5QQfROm2FE5mPPljJsWBMhrbW+t3AmLuo4CLXf8u7v/ARHGRGrAGrg/x+E
7qLVAR4jbyrKgTLq4Yh64jlsYpRDoXGEf/TjO+OUG9ar18YLohUPLpgib0NJPxMf
VFSh/bn38bei9lEOg/Jcd3+5j9hke6ZPHb99rc1P2kbbhQQXrQF6HpHnAsQpj0K6
Z5D/G4SsB3Od60QbOMNq7tGHynEMNlSG0gGCwkt+MJSo8X42EH1cTQLUyIgRw8nt
GJ9XIRa6dvailtHaBcW0dZN3fAXJXsxQW1ht+stZv7sc7xb5vdlmCZyjLHFbhZ55
mhFTgr2x0ZLos0d0X9jDYg6uaaN7x4/svnXeI/WrhJy0lb7+BOWqI+O+caQ/Ocw0
EGNTxZGGdJ1DCgpmJyT2yMABgfzwxrP/b6DQhNshWkMTwOyVd4RIq4nkRkXVzeJO
1n5+Il5GA5WAGRrCR87p22TWOpTge9MW0R7rgRkxDmXADw5FF08KDATVRVb1CmdT
YC7hLmGUBAXP5o5H5mK6qCmTdsdnhVsuBofdQUMRWIiGVvaVYcSgaZK+GdlnJAOq
h6EOPl8C+IRLuJIHbVHm1Y7mNDmmrALGO1QZOajOvI/ao+KaphG5AvBUobh3cpy4
TjUjooWJYubDLKcTdafQit4XM5f/kvkOc5eZtJHgEe353WUyCTuaHdewFqnX8mbt
6EQfyKBhX2jvcDdOpNta83M6Myyky2j5s1tNGZGif3I5R+dS7xhwnksD61Olsafp
21PqvASyCRaTchHt/eoEr2hqhsJDbvI6neCefRveRJHZYwL8L+aIfYUfhyEbF1Od
hfh7O4JaImgriOuko5M7zolPvTx6lq+fix40fPPwxtK3U1PZLvuazjUT+QcgPxTA
1q7nXLQqme7ov2hP9UMLUM3YbLx6wwgdTt4Yb9mvIQCjNWadNNjGep/WjeHUIuui
U11ERSYrkPFzz/Ju6+w8Tvqs/0iSBrTbbqboQbKtwKr9lG2XUQl1r6urPWREApfP
fyxFGG0/ut15VzoicWtU1wQ7JBGDPBfz4j0hXz2gG6uIeEH+ZEqDN9wyInHdxx9B
RC/bZwvLyDzP8uI6mbae79MxpGWKY+TsdgNilkVnxZ9dDwSMmaB4+1JfVd/o3Jjb
a++l7DV27AhnvdfBK4GAc6Defwd5wvPvZnIPXYkTioFbY/ZP0d64/P4EGaFJk5mW
kBx04vpPWWWn73RgCIcjjY5QXfDlEklW/FNQhKLIuIndDUwyxXc8p4aF0j5N3bRp
XfEJpefaEybaa7zXcjdUZCeSM0W9nI7JLlax5oNAt5zNnAlsS8gzuvi0NZgreXjI
F9meYy5AnEPcOlbSLZ3424kktMhCfOpWTk2oVMaWFx17860ttJjSGGJMj6sI6eDV
dEyUtg/Bj7NiGRYBcL40u/uB5jK7a5Q3ysZp3IWdcNiqUrYcUbwi5x1O/hY4aj6o
EK364nvn9XDHjvvHahUupSreAaUN44/lEreJ3ewBoz5uFiGKCjnmqI1S84FyDiGF
3PK51WJT46y4psv8Frcflv4cXECfEbmI4A4uA2wWMX3MmnJaISnq+D1knE8sqtSu
94k5N8onv8UE05XUZcxQnvq37/aiCXIw0BAdCmWtZfrI8fqCUaOVfMXXcCb10CpR
XYKf/T9SbATzaiisqoqHBu4Z1prWl+2MI0v0RqzACb45ZwWyC6951yoJ0H+oV5xF
EwmePVbJ7JSjTF9Ca7XZu1RcayI/FxVY8RhLaXFWTnNlkuJ+5xP3BVSExo6IRr5I
gGxEKJjAk6fDdDNciY5cU1gqnfULnIE+iZBRP7t4xSg2JtOzA1bcKoSYPc1vGSKZ
7e8O7HF5j8IoF6732jsyvH3MlEgghZvY5F8l84fIu0S1LDwXyXGuGu5fIXFtxB3h
d/fZBl+0blS9MQrvTxfqxgKzDAcQ0b3Y8D9fBag/8dCkFHDeP517KoCr9uSjJz5K
ZwNY/J+ngm0OucZCJD3pjehL7csVY5izf1QfTMexlvAXAml+5BPXc9X1jh1wm0Aq
jMobl1RgOolUHP7BXDiKXWTiJA6YQuqPQ9BM5IYi+Km4tcQLFLGYNF1N8s547R7k
m5GDuvbxwZLnj4Pqsnvlb7k8H6RE1xnozPAC1CcUZAt1RoQr9Pys7C01PYrcnaM2
lz9pKngaRjkq88PBbaYcvWwwsvvPPMfC8QqYQVe9ewRqLR/p3GI5+cyrO/aFyxlF
Hv+rIjjueUFLIrpyoB8O5d15fetvAS4Ioc811AaYlFyM6et09XDUoQTVcnewbvVb
J0b8UzvaCnL+FHX+mwJwqQ9NlEJcbaP3N+bBcM/fzUV+A/4bG5IzSvgPwQ/Mse8r
ZUhwdInCDJM1UDFMSXWGxs6U6kJEKjUVGy8XZFOMZgOw9TKfK1kyAwoCj0hFffYV
Oe4dMmoaI22y3Lib7EvaoggOnv4t7cacDgCjbDH0wG4ZhV+PiQxIjeNvMVPLTMBn
IpxnVypG2SvMBLrmFQMmoYXY/lx3I/u5Se00zTOMrLr/4jMIDPwotOVsxifrNYzN
lmVVsRYEiAIaEBVVlYnBLb1tnUMk1csHXuSYA/uUxtosvzqay23vs6LZ0G4ktlsj
DtGAJjjVcw+MQT42Za76FXGWILsanYc+80lqzKhRetxGfEN1qGKvPWchSwKxrxVP
QnrwFk068Xv/AUIM1EkWABoBSBkYqIeK1fy1xb7ecQM4Lg7nOELK/f12OEJTLsXh
L+GolftGWpojRLv6CepIi0xEUs2fk/unFs3jCRMaFyB52zEqhUN0m0HT3Uc8LihU
rcXxSUSQ6lPddV/Wyqe/5R1k8DjyU8VDu6dX1IQyZjeQi3HAQHaki5chlZLWAHEV
vXjISNMOW406PjQKhe0HZgM/wM9ozaHGZULV2wE9AupNjzhqWbz8UI0IDrQEXewo
eMrQRIq6ZoqMhCbYO+WC3ZA4ApP24zKTrnOzu/cUXyNPk02E+k6kpKH3vSgpSc1i
poPBhicBioMKh/RqG2SMHpyaycM0kT8S0qSueksvQhdLq4hKjKyMghATEyJ4zpP3
SEyHinDdTjuHS7thgtYC5Fry+JitiiJ/uWLcPl4v4o2zN2DqFxPZLuYuHQ9p3n3q
47CB51f8AzKOaXBj0dWqROhY3kzjaoF5iunX8z3jPtEM35Q8wSE3uP54W+do4SA+
ZLP3kUPBpZVMYT4r7LUErequyWHl82HPKEJ98AWqDnFXYQGL2g8cGKWAYAzj/Wve
GKWoVF7ogDG6J+66sVdRVKQbu7mMgSPzU2vmhWtyk3UsmtHRYD7DY/zPsCBXgaes
sys501DE4yx52jKcT9k8m9LkgupeSRlCY26Enmz0+aszfxfarEN9Mqt9NnRVvCFO
HxiKH1gkkD7vfzY8mLmu8KuCTpuyq7ZCXKp+6QseIQtXjCm2LpvcxYTUc5AiaduG
C3hsxCDDPcovMC/q5qfiDVMrxHYNaZFaBT7BsMjSvOLdRy0GcRP3oEHQAmSW0Byz
kCovZ6w9uDjK59s/q2AK7MBjFuYvgvuCYSbzkRr1lX/D34BKnmoHqG8GGpuY+zsL
c+GXrrj7DrlXm+f+R/Gv8Z7AFl1SABZBEjUrYIr1qW3IDuUSReQN//fE449amHS0
d1kLAlGHR3ys3X3u89hbXScuT+PM//jKzp7dIAsuccUz2IJPYJ8c4wesqV8snHwi
uEMQAuzC41gFKkpeCtfM/D62OBSIj4C17ecyEwF4J4uhcVTytGFEn4q34PsE2QnJ
gT1bVC5nXl9aml5ANMDFFBvvFKuDxXnayipbt4ILDbubJvvTsKt3RjwUjrt286/R
sgJ0gg5gbZGgfvVChlLrNITKsu+1LC2Pb4nToYa3HWxtew7nqj2GvpxFqOzIUmGP
lnb7m+xnbpD46fOimNW7RAqj07pSvvQ+tUxbGe9kyZfYYxyRyDGXiHAvk328hnGU
RDW9g3MXnn9djCUxyloYqSdKm2yDn7L8fgJxlup5JER8vEcdlbIX5C2lgBxKJg83
rx7Szuar6Bn8xaiXsg4U+1nl+TEz0k41cpdTNZZG4MPHLPYjU9WFFzN+dG6AnkhM
bqC7MRrbQ4N5l+J16Q29026/CND81H7reVcBszBU5V7LSB7+UvxQy5h+5cimdPyj
bHCRjDcVQnuam4K77MvmRs7gjnC+g8U+97kkIfwjWZyFpPSCR1N8Dqrs0874hM0r
DluKdPiJOTL9v711Tm9UTAVk4XexrWJ1F7ho3lcAuApFRD5Zc1ZXiuX2MTq2D4Df
4CoIYv3TP/dVaJCmOFuCi6doWZPjKwMj9BjKeIpcwAjQeLtZf5Lp/lBn/SHKcEcE
1P3hLh6x8uAHnZ+Y9GtVnQurQZJwzEKCj35/gjsZvW8YLDM116rV9s53P9upj5cj
iEODPNHUw8l3Fy1sRGxcFwQvmKl7zGiQxS9D41HzGSnPe99GxyhtiECFXms+3Er6
JLa8Q7PyCJpx0nQWadDFtyyBtAKauOOyMEHbYD4S6NWxLdmRqtmFvK3oag3YQSx/
CwOzCVFkQ60Lrl825b0pPdCjwpuB3HZl61lIQ7CNs0a3qu3ZgSSzBG8q1k64G8da
EipjGDjSYX5mbmvPw9drObtZNO9f4InoTxjoEiasKM0onFC1xiQRHQCIzin1+YcA
+g9CdG5wkYj4Id+NeOu1qFbcwsS07VU768VEpxIPuC2M4EHVOM+Ny6bGIGHAEXLd
+o5vy2HyVT5q4eKzXQZZ52HoxIoUJs/uSGcNR7e47QRU8CZxTcFHzS7BjOkZ5m+d
1FYpeQ2t+tz8e9cBh4Pj3CDsQAHtgMLnZBcZetk8dCQgNwM9XNOe1adlxK7CqvEx
b2QSc0WuS5Azo0tRZqRmPXxtzPmok6apZR+euI1jxQptuAA3KHKQYfqL1QwLvOFm
LmeColobJ5dHwqsfGe/uf9SBIFcIumtIQ0/nFhcdF9VrhGnatd7iPeFaMDc5PV+l
p7iuZqelJeArXPFXw5E/nVYKbvsIPa8sP90lgNNr3OujmUJ1X3NNMlfuKfeycOIT
WXs8vkTdQsqSduxMrD4JPNuBP+7Kv9OAQglck/T3g1NIXzI7yglNYSOrAsRKd3WB
6wTz4JJsqPRGyzLkd3iH2yvLYw3YaV8+eRYChm8Re5+mZYyxylHzv+mW/1DskO3k
xjCMGJT3TzaSJSN8EOtebNHNg0yLFjycNGryborgF4wU5sOLtLL9xDvd1h6E6oj6
BQITZHFyoM81TMZcJixGR6JAVHAdhcutx9xeNVo+698f/YMc6aMQmnba+QAeWpr2
kedP8xOZu5odwX6ucd6acBt/TF1Qlua+jHp1IrZQJPBodzPSB9d6oU/STfbVWDpH
CBiu1ONguCmiOkPngZCPkXmtmWlybwxfl06HbQq9pOH+6z1CKEfl/j4s0y/JnuKw
xSjm3bcG1dW1Z2uDzSaHK8qnoz7v8uoEDOsDn7NMqSMrPfvw5AxevYSO3uIzYLNt
0kRD5YeqxWzJLXVKf9iliCW4vkS8YOOlIc3zNbG6S+oJMdenHN/q8ZOSgTLn1CZl
qwALhm1L6ib/pCfxx/FVQS+q+ZWiunPtahkRuSZ4mDb+o14aeu3i557uHIvPqueA
t6j80U8wW3uYVoaHuhP9QbSomFEl20LJU5tTvlLS08W/khuLQkst0PiXHXZu3bfG
mXRDQIhu16HWvy5+H4MnTg171wCkle+6MYB8pEJk8d2tezlSU2ONZu9VDsdrCGJk
Ds62NF5PKZYnm706Cx1okjsl3WD/r2e1wUisqtmP+W6W8FWAjG6CgRqfYZT1QlhO
LAoFuu1bL3j+ldTbCZQ8SUyhRtGJtrLhcbGIdmBBvplV39sROqTRuQ0cs9jQIvhJ
OA70jSvQPTxyrKmJ8J9tdsx/Z5m0D5g4uSuOpJDx9P4PcOJujbqAue26l80rGclN
YRbwHhvyR6IBXF5NFxHhb0f34EuA+w0TLyha740jaDK1N7BWUmj5Lzeh2HanTcfv
pLbalcRPVFXaPVyJCkhykiTl2AtNG38+Z6jUY5Za4ELzWqylMBAlwu6fuTPWx3La
D43sNPrXOAlSQxMHRVLLaLA49wT/rt25TatCvR3zwKflB4uqhKgpZZTZ8rVzCcYY
mDWKCBWyXSc/bI7exo4tXa1ZpV77Kq6wJ79PGN5ocjz773D07cfGqng83EhsGNCF
cn1VQ96plnt3fA4gAlYPapm6rnptJ7DPIbHxTGmXZzfoaJPUgd3txgiOVI1TeeaX
665y2Phf0hzpgQj1iGUBKH5ryQrVSCuTwFOpSENxtPa9S1vq5WJIhO8R16i3bUqd
TiPPrZbSNjvQJ9+Jci+wGXuDoq4h1dn6GPujcguLw3xNuSOp5i6tuKveWz2GpHtW
TrswygwGY1kEp4DzhpDLiPzf8ei7rwkt6gttYLwWf+z6HY2FmCX8FMxsG6z4daQ1
SddeMiHmGvOLJL9h9ZHCMH8xU2hQ8NDrIcr4eqsV2+nI7nh8UE+2bQ4w/tV8tNBu
3l48o3x3A7YbmNAfKFhVhZOHQCBzsj9JWjKEalYtAY+nV8X/NQxcn/zCig+Arkdm
3Y+AuKBS0Fz+bHrqMxcrdmddg+tKcQEjrLmryMq1j4NqCoOXY0BARGtaYL4ZS95I
u9wtBaLWN9IF7Awvpd7ukAGmowYAPDUEfRlgI2SbTCiPOFN9mZPCL+glazvuawDB
R2LFo2CPHu0l0eviswiWOP9oYk9M1AAG2XCZtRsw1inX+8sAxgd9REj8EqCJE7E7
FXN9SfV4Y8fOxIARRbNM636JD4GlJLOtX31f+HjWrYSxBYCwzn9DxjQAyB3zyqe5
0lnaRkDqQSJXkJK7ImftfQirWqF8/txIkTHY3jDtkinAGWfKO3zZIaWRce8UyOsM
1N9TST/6UKY8Syb1u0QpA7EHPHU439dMec9NHtxhGLnsVMzgJdZK1aTCGPU6VmiV
ILC8ENnkvqJ2gK3uDYccC1rGiIidfzgTH8/CyizDNIAGX9Vmrnwa4zUzRa1tfitB
8DHy3fpLIlI7jUpLtEZbx+xznmvBz3hXBaNmEXaQoIgf8Rgnhlrvx5DvO66h6EG9
kjx3gl6wXk0Y85uJaPBF1grjcG3G9vvphlAxSLECt3vJt1UTj7CUIFxFNVU1jBjA
sbjufKeOcfs2JGXqYXJ9kdxBzIwr3OEc7uWs0ZtUPwa4yXQ+8v6eOHayZocGHg6X
AixRST7dE/USNj/4MLyEjDWgUx37vK1xh3hewaNhu3F4GhKGHD+hvUQ9WiZj1fJX
smkFE8VwhQr5GDj0Eph6WolYZYr/7cRv/D1PmRDUxlgnHzCGkGQJCLPddmNFsHsY
1y9KRExaiJO4L6LxeqnaZlEEbySXE1urDCx/nawEKIJlTLobRpH7o+RK1YLBzZ3K
ytUAA2bWeduMJuV7UPCcIYaEa4SJkUYzMrG3jAQutiWu2qHn4S/CB2GO8Tp/HYCi
LdeJD6jnCKiWDuClIDp9a6hUSagZgyt8VNaWSnpsHScGBzdRbeKtVMadW2Yh1ptP
IZjtLg9DOGL2gOwRVsLT4+4dnC1twM7m/dVfZ9KjfGSPwdohyrhvGTmcqy3ye127
p4Viuwp+w6UXir/qRQIKo1Ao6M7H9hwApMCGFIi9/zP+Ytmj/AuFvCK4cH/uGcdZ
QojoVfyEj/dw+Kb0Tkq0RvuJHrWYCKT89qRPFYk/Eka4Oq7/GSlFUd3R/Q9SG/Qn
mSp3Qy549CF71fA6Ppei6cmx18a73i0BujkVYCJWvjgioVjL50YVApiJ52yz78cE
4CHP6RY8IU/LvMNCTGO1jti7LVgPaN1t9AsMA5PI7yT61gsJJ3BVTNIIvDSDSwix
qyMc4HkLw9MpHNbAvWxmauA02DlxD+rTs/i1vDTKMdWH90FcboqfJRTKw1HzPqVT
UY9mJmicX48Lr6RKuOC4gRsmAiu0USbb4jpzf3/bKuOEF0GScBNg6zQu0xBbDiW9
0nexVW5ASrv/KFxtSCUXz72lnPmgYNXaY0U85W4F8mbJ10SUne6PaXHwGtT+4g3H
dHSGOuSp7pR9aIkQBOe7rNbaVDfy6fbAtv+5BQWiRlLR7tr/F6bYkf3c3RCUeacu
K0/Dh1Zo7DZdVyvkm7Z2IKqBkn95gdAit55oOK8rPyMLA0VtfXbFMjYAkbBYz0YA
ierhI1bzVApJhx2vNgMdwTiVJJCQ9Em3ZID5yYaAZKL289HVhWHpdvxP8HJKk+Vb
X4nqyoxfMSb1R3sDi2rQvC2XryatIW86chWeoJJhEdTBZEPnNPlEDwAI8LrCbPGB
ESmvhpJ9dSmZtVqSDBjfopKMpXVunluBOzLK6BcnjvDNT/7SB1gpCtK8RHdw/MOr
p+NkHWVZIOMx70h+5gneTV1L+b+x1UlB2YzN4Ai5+LFExdvFx5WsEB7v1gjMrq38
JRM5CFRDQrKU/XdbOIN9cs0NXlqRaqeAnIIbL5PnBbFPip1LJwDE02s6wOZvu/ki
tOcSRzJYgeR/Oz0ZCDEXLfPIsjpsWFrj5htP4WboIyilxq/3FZs3+IU+/6p9roYx
ClJL8gu6eyeXZPQpFS1rz0rfT9Nlr60K6TkKX5EBC5+cEWALX7/T6Tvft89mCSC3
a2S6VVAabfNApLdzL8HSOYGLlMoj5ePlVU4lWPjcbIhVhCbaaG8iYKNfkSBYJqkd
HsEYGdeGmAzyzBVOfaK2PqLY/kE4LmBSkdO6q85sAz/Z9C+C0S4LldxS2r6dbOke
t1joETgez45wR8HZZT+Cp6h1jDoQ2Ys98buk8652JfzU/EeHHkuuUWt9kxnkMYYI
TlCVwT7/zbxnmkAKIb16gvZBDyD/BgEpleISYvMoBlvwPcE8LdHocUQGofGHAqmk
nZRjzLyJm/Q2zvErA6grZTKEiEIdvoMeJc4OyPEuv8DkZdXjbojinMrEeJrqYlYi
xJp4jCSf6xg0NiT/Q9uyBVmxy9TJAnaVE2eLukcdWP5BMZRSaUd6hc+PxSVMEYFm
w5sscl+C1ppH7g67/ALmts+bCQ/9NACWjF9UTW3H/BqKwRQ9IlITmsyHjqLVyjp2
GOF+7wq4lZhCsjpbTt2Hf/W2M+Crg3WDVUr/2722OYxBHdVYdpyaK16GFdpTJllI
GxkBKOcd3geZ3e27IPyMk6721XzYVtAn5Dz03KyRJ8GWukZ2lRmRPOcjoU4DpvPm
glcSnxyC0CUvkzAcfvKb2R2bPiil63stms+meBu890/viskn1eXLW5WW6ED3gkCP
A+FseKppPPBgmcY4PfW3kkJscffUmgvURmLBcrgCCKUewRYqUH1b8oQoHe6rKJzs
v1FZQkQ7qpH4sGrcxJ2eSg9vsDTK95zX/Eu5vcJUguJwzIDgY564d/TvCN1cjug4
4iAu31VpIAbdcm82lTbWxJvieH3GiZOtqCTPwskkokN1Xf+Lp5eZH51NqXSVk4IQ
ouB2pnZcrsMjoQ5ggcogkwyPu1g3V7khEK5kooBgafC6V268U2ekv0vawCx0xYew
tSgqMyGZjdou8vHBgKzhwcF2UE+UAoEQFWrrceTzKjLFrfSottSX6x5z433lUCd5
sCwuLn0TcaHbSI6Espqx8yBT0k4OVe7Ji41HQhqcQFvZgml5TAf9dEz+htgmMNJf
4Vk5d6SMnblRWkM0MB+SNmoB7YvSm8EOOONMBbRRqjp4/jpnYinzeKspKT12GW6a
3xOkFfEuIfcA4u29YrHMufRwWqq9fdnXRzBe7AGPykpvxxUnvVHV4WOIocIYbELq
yytkTfGq+dP0JouYhxj8dOqSUyn72GEAnCTZqlB77k10OERbKtroyb6oeWdvn04k
vpuSIlVqNpA2y/eplv0CERicSoIrfJglainHWARMK4uRQZ4LbWO2ZWNOAuGmlIV9
oBQb5aqI1PGDQA5veCw1bVXDt7XanyYpmn/CjDFEm2ylc7m3Lf82xP2Uvm2NXXN3
HXzjvB4iFVFvqxJv5nzzTVZItDQHs6O8YWis/1ffLb+e+dpS/hbHsqbOHgx+gdkb
16VqJ/5JpzOQvu2w+7EbRmxbs9lElY62/nWnzN5nYG6M/tinZAmZDHHcjQCFkaPH
eY+vculym6ysUXlN9dXgfdy1d9B43LfQZhC7WdohHdgjY0RPKcO97BopPq9GGCfU
g2VH3FwbYFgtj4tRykqDLieKvODNOh/LY1skSN7rqHJ0aoicQcgFZGVB6R8aWvnz
JgDase1/UsFZIirHia34HzJxW5tiSBfBegmVauol3+Syh76TLaYd7UHgLloSeWRw
pKPAjFenMArOFWHrkAtk0lUm59NFpx5phmmzIan75FvmN5Sds1Cy0clJH/shkvfa
a0qWMfuXzLcsWQw/e6SCvHr4ExFc2CufI/kcOXDq6dg9INDaQITPYfsvzG8qtxoX
uPTKCuAQF4u7qTmI4XLdhNcmxjnM1Y8CWIvU7sw4aeNle3NpIPuIl0YH8wvgB3SJ
XwI4QxW7mD0j/VVCjdxmrfihzyxYEyow/iaFfeEg2CX4wr6FU16zWEjo0LcNfaEc
IN+mcrQYT4d0wPWpggBHsTNW3Maa7DaIp1b2meL2kfIs0zG2TnIqL0jFFks6jf6d
2HnYor3Mc7+BCYTg4ciykJ1xDnD1HSmAn+F3cxVIdMD7uP0PCKIxMfwQCf2thmyI
5EDe63dj/TjTofjaw/3oTTqRRYQCjQRfizmREchbbniMtgNsmCmxSt59rEdbQDWR
X3owRieUDhhIYGY8XlXhUHNOrf410i/Y+AtYRZ2Nxr/10UMTigtRRPhopyT8sEK2
up7E1ggqiUgX//6rGSdaLPYWAaXNEmPdgl0xnZVfuNXIKxs/qOYHHRMmS9H1+JrD
hd44gNlJuPFQc4dBe137wHvHTy98SzeoH6D06fkjnIJ3cbT5fr35Jdv8N4GP00To
TAiGMviXrGYdAeg9JOxbrNY2Wx+Bv4ZDe7VK9GiTv3pnvHyWK9ddhWL+ChVWZiYi
jqoJ+XC55GySVMzppVa3G+tHn4CoYiBSvyHuXlpNnwygHXWfuXkRlVNtTSDlxYYe
JMTisHPdQXlgv4+ctFThk5IABZH/nucNOEp9R3gw6O73bfk9IT+1PKGPAPMeq2Ak
YtLQ4b9b1WAZk/PBDIpnV093qFI5iNr9HQc8R2P7NocXoR9MDoM2K2ig7tQVbyu6
MbSVWwDSe20PPVV4HhZ7K70ab5RkcRN8956kCx7fA0NsmPOovDyXwpUWl2PKd8Hf
36ayJSzYsroyUai2kvoVhjApYGSwFD2YJuRcQwicgoCwkfb+E/q43NDurogTm6j9
k0H8SoxiyQ3/yfN/QAPnYNkKPVDE9lglfUJwQAqJrJtjaEzzh0k8g4FoikQzAuOP
2ZMuwHGbLlYP+03jiE2DFxytE89lQruEVvHVm8O5kQt+qBW+kA26utkTMwTSqSW8
a8PmBORCkKyDhsK+Gy1CnTG8ns1q59x6fiuvRSkJpEF/TFsx4El9BEY52Tlise0A
syknW2ylJqCYiLc79T2bWeZ3pRGKfOIcPjOGouCOCTTMtbYC1olnWxnjoYRzvvMw
+zsN0us2iekbvrj/sAAy+HcFmg/F/svT+FBpn5nNTBQ2W2LViiHghEE7I8ciymlb
nkOoPE4QUQiQhwktiS0t1MYSG9/v+2zglnYlnZjpkj6EoDcDffxE10FwQa4cr8sb
BXwLh04WU1Px/g16Fc7gD2LHnt7JRjdJJSIWTc02zGSu8jKw5HVR0hUgweNq8T0B
BTOBa/ohUACkJQXa/xAeqbAwus2t/QavVNCd6S/fxMqc6awmc97BRSxFsQAiNaf5
v+enDLdunM36/LxmiGdWmauR/dMNhZeRDhTMJowVf16SOfMbwZvpoRbvUSfQ8zzi
MGXlWkdGzQLNM9AfhL22IUasAsy23o6G1gLAR9rWiagPkjGiFRu2IY3+/StTmLZX
Q9VyaecOgGB9+cE9F0z91pf84QcYAO5ytBH9DSCz//EXgTcTEnVaRl2jun7COfym
0xjHJpiokq3arUInUra38Bd+FHFj6+LCukceAxToszL+mRHB7BsFR6cgDVmW3Kbs
QWNd6ezZXRRnk9i1QwyvRnY2ituVE0ypv+S44or4/SY/oISH3lcAjpU79Mb8nJkO
yjKEy+Tv6rBOXdRyoTI0AMQOn1JZxePKfn72TAgURAprsMVs4eITpgeVM7F3KB1I
gU8QFFcQX3A7qbmf7HMMLYZb+sI1olQpHlNVYPz9pZ/t5bf5paC22eoppt24DWUv
yFdWGz0uyRrobbt5QaVl0jlOEj/VVc8bO32aqWmLnUuk7yVNHagTb46VEHRsVo9Y
QASETslOl30KV9SeSHNBN1oVwqg7+9RYiiKfoY0TGAGUsRt2znmP/ky91erCZkhB
lasfpmTUZBZQFhmWykeeyJztLliL1mZlcOXoA+AHBrxpOCg9jypjaEL+XUBBafIl
vHnTLTd9qyZyDkokIroQC3+vux98rJygeLLbW1jcCs23ANsdlX1adYhdbrF6czrr
956+/j8Ed2Bq4pQYKUTf92FmcVRhiVW37QGr2cEsK1v2GRaQbB3Ykfnfi65xAGGw
anlEoVEnR7HZfJGPDfe+Nzvf4fjeIoFGkSIGlKm01+nY+iDzGjOPk+yuqbEwYf3w
hT1N38W2svJp3rqTgZ5lmbIVab9epqJ8MTwMs6/qoEV9+eXMSQBxke3O3Xbe68Vl
MRENgcYMKI9z1pcxBH+G/IAdxovPVwFcOvthJh/frGE0LkXAeL64W03wF8ZCGpFG
u9QFKmFAuhQoMtR/T0520ujg7SYA2mPPswmcH1U3ekzYYYnAFKfwyFuxrvCMM6Eq
Vxvft0S1tg70nPGUndtZDY87M2x15XRIUGlEGDHp8pCFJWJ5fH07p4WM5n3+eaYt
YdTNo3QsgcHFv36GQTnTeEvVafrfuvJEkhP9zE0/yqZnpIp1H2guWJ6qKbV17dot
V9IS2+rK5tI46WsHafI7vU3fwxwftH7u/Q0JCOQZ4XQgQj2YvlH14DZSMXBbZ/W8
v7KhwF5wIEkcZ4P7VHsHjc4bma6JcEjCk2rimlz1JsaxNY0xNnKqwJgyDLDkslLn
wGoZl9wpB5xjs9DFEoR+qzC9D41DLjh9VtUg2+7OpexWhA/FyvMO6UFUzFGnn6Ok
+yZN1+ma/KTBX9y8a97ia/mcsKN16wsd5OVBz67rEpdfLYculEr86ZL3GbgKulCN
NX5basqRO7LUEEJA+r7Pi+zyI3o/ZUp97bpkDCXWp39Y5wreolpcGLDBaKaRznh9
gOmWjIqfx0bjLTSD/V2Au08kTMst8oBxrMEdWJlQIX2Q8yqwnXT2JuNjxIvyGc/k
CTYlU28Dl5gtwdwmGsZedyZCxsWYLN1CfT95o+gza0qqtmIlTUjtlu3/8qPui9Td
KZ5vbKD7+XFCobvgr+scitiHa6y90863cKmvlld/918bEW/QvvyTTSkAvHJ9jBNF
U10rV5P+2p/fhBINd+bHZQhSw8Dllsv7J81CClcjpz4ztXogC7Gt0W424QbhGZ4r
MTY0v8sNbJ2hgmeFAUzAmkXKd9+INSLS++6dG2b8b3Lzn/WTOHIgWACGXvdeJczY
VyJ+tbNRE8/iGswnEzGw2HO/XEt1XUJYovS3jSud4iHe3+vpUbsfrI6egMGHijX1
ExVudfIpmWoNmLwZt8o88Ar3ihzn3Caj3pU3WgQf68dgS7yI97fYZFIYyQA6tOXS
L0JJbrcKlEN+SB71CDJw22j/9Qb4NQTlxGSicGDiwPnkdnB0RlUaCrxBYIEBh1YK
JLg8Skbg00/gtGCl4pGFo7tWeFC9XbI64XKZJs90Kfdd62E4SPdlN5j2eOZ0F6M2
5gExH4CX8NNv2kKqD6f7Vs3cUPgHfMXy6wAz9hQ7ZMed4X3GS1N31x0HlsfjaXTR
7gHFIiCk38dPzPx8xBoQRQuwFW3fa1ZF4nVyeF1K79V2aaBbzpJ6VN/m2gism6F1
4gfjy7FyOb33KvB1i2BI4MCLigbNqASq2iiATkcbsZUTtkRI3a2nIqGLlZqr8pLf
m1hx4VZyq07fX1zjRmj90EyS0uqmcwy4ATR7MdjJVE1CtjgOs7wBbpY7nZDQAV90
N/MLtjniqUCgRGhAlGzmhP1nP9iWzrIfKap0UaRr2obCRq42r6pq6lo/vjuSRMkH
2MbeuAV2o7yTRVt0zrtPnem4gHA1EsUFsK9PkWDPVa2/niRqqIKn00e/HTyI2lCF
hFsZznoOI5xQdtbpecshUgVtB8Q0ReGO3uk9opG/o7m/ge1N5VntvSYV8xHZ9ezB
1qAbSp2bWuczICCHGZUZ/iNh9vdmbABFFsdOUGjdQoNk7U6dUcXBFUdx3aBY+YhR
Q7waiiKzhn211FWV2K173jyqKhZO3qjvtdcgcTZBjvXFehK9vfvkQOPxFWMPyNpb
pdse+EUQXzTZrXOZOig2feoWakUSA2AgQiGvvcpzbUgym1ekLkEg8A3dUk9NGHcE
FOD/ZNzAqSR/oOCzAefL1zLKClBEAVwYrdIMMe71+lT4ekFoW1I6HBYAEpjcYPlg
SD1f/QS9pSsSPDUOI+jYD/ZiIGonkGB7vIG6O4AQWNjyUPVTPVhBzgb1GF5H4TrS
1bVNDNOKEuGwzcqtsW44zKuGH2NKUwYiNs0Mb0U2t7kkqGm+Wl9nuDbu+ORT1woa
n1r+38XlN7qTuJdzWxsQzlHP3HmTzKkE4b+vSCnoplYphYxbqYx39j7lLVk1Qvho
zfiRYHMBTP/NSyZjX4t/DQfn478eYs7ll0x4KgfA7hrWq5D7HjSPl9Z3fVZu1rwe
u2K+4RrrsOvvkbH9E9uooQpITotjq6ot1IRtSs7YqLEgf1lQ3iGQUQUhN/P11Aw3
ZKWQgIOt7iaLg05Ue0Rn8NE6aFs5h0mVUSLTn5VKU8BKJuSCd5Vp7t8O+sZkO8YA
Oc2zFISUwLiSNHz8PhcVtfIPuT/I12ZDItoknGv+xtO0bIavvoKsvZOmWYFFGFQ0
EVmGrGMafNdxl0k2/UpXIx5ZKvBz2xntYdtnF72AXQ3ZrJJ0gGE3IzVxQ9hBjbf9
vfm7uyouTi31O/w5whAo4Vhur2+9FOzGMjwKuyRuqs+uXUdq1smkJQCR1HAp9DIX
mV7mxjEXyS8w/k0vePaSQzTD9aY2M7NYy/GMpwu4TiWHJC0+yv87aKAb8qs2dZ9R
dZlM4uABdgYPSxZVqcNC/3+QM0AOUYrOKOepZAg3RpyTgzWPr/M6YcuUe4rf4BIv
il2FNvWiGcBfW3mSpBASNh6YYE1teJ3Ux8Yq5DuIDOvK+5NMQoStZAUekDMuljyj
aKfuxZEgZj60nV7WOFltGuOg4VGLi6+Mb1wpm4g+0MIeBrkJmmp7XflFadIbNlAY
ImPk1CMqGKOVCoe2YFXFCQRhIWcE2fR5hYZGcGK1AgSCm/wGQ1GVAWemEnBiRrKu
ILuAMgD+N6/UJsz2BFpWdRETNjiOI6XfsPt8sgf0XgfEHgGeeWXoBYNv+TKx9zBv
4pNM+pXknuiigepOaDXw97Vu37VRcRcL9PVTBaabwg78dJiNqrkSpWI+8XzmgARA
7IIb7lp2HqIRHw1JiUmc+Jy2gree0yK/KsIGIoKav8IPYqVW59G9xIruDcfUZb6l
LZ77eqTSmH5iP0aV2vicQXg6G5v0XeAUxZAK3k8SHwmmsDU/4OUT4XMwYKvwGIQ7
uYTDfk9GDHH6HHJNP51z1vtvUdcIoxxNMD04RDYWImakaeeIehqN7fQUb6XIjbSf
vHezgrE3556j3sXiN1IhseqAIgpGH36iEmr6vHmi8xlPKJnnGlfMJN54rcui+ejz
uSeYerz03MGe3ZQCE1ldUuOagiVeBFPOweapDaMntq+URxOsYag5rfVkGnIOrIE8
voy1/0YXvZ/OK4Lv/FqeJXK5Ay7IxUwukcNlZPqbJFdtCGfn5z7ne6NLS/ykNJ2Q
b5U/ppnjWvBSCUdguGRtqW+GhoLl3LNMP3LMLm6JjSVTSwYYy8E991LuMj6+o4pU
e00IXKQjhb5agtscSackzpPCN/9sDlzMMZWiRCgoO+mvw1H+/CSIsGpuJ1h8RuoO
tg6oi68h9RrSS+SveQQtVEmLiC7IJTu4UveCFe7MWR1FVvuUaipAZ9Uqb/AUoSS6
wqZXvmMn2LM6rNrt6QykQUmfrxtJ61RxD/MsXW09xZBlkhLhVsSPZsDnbodv5EA4
xIfLkjDUW3x30iyhyIFCqzF09HUGmXxXggayfiZLsC3oGAcT8qIn6qWgErOTPQTA
nTx2flTUmhsYam3jvGTdr1rhpzKSE+kArw5wN702A/JrQuEhtAWF3IExf3lIUwko
BHZ8oFj1+Fn62KHnaJCuJpy68knK4Rh5mAaoPRaEr5LoSFWwnva3lik9wBm6O/9r
dLnusd9IaU1Jqal+FmogimXcdkrG1yhK6oRhPNFydJn1Fotba7OMmND+WXKI6f+9
jS6LSw18Y3kY7U5zQy28d6nG1hpSlTM0luiXKd9Y2KUXmh/qdfilm0DafkFx3Dej
TvCksj+5SHzcLwKlqnp3QuLhelv/ymeWvXQVSHOJ3RX+Grqzdbo4pJEoiD5OEyMH
4T6qhvCu/hbasbbOkQ0xe1RSQPqks6R4F2C4OmNYTBSeQr8PDtBsicMBUYdx6I6u
JIUq925wrpPhWS3eJvORuktzNbdpZSTzVPeqXSgnVpJKZF0+9CvgyzTcf/grNj2s
0AlH+Sgm36IxowD2iu1k6ixfUAU49DKSbZGnvo2pFaU5GhE0ivwKN18vshRhRGcI
PIeaoJLHyIMDOZAsPaPRWKGNUi23BkQqnEAhviMzM3nclBYd2yRYwhqNYZS0DXal
BudO2g5SlI/025hXzlXFE+/mObb2dSONHpWKXneas0Jyuy56qlGdIdKG8Veu8Aix
g9NLGSO/GnTV7vcBTmZnaSX+ASbzvxkeMXV9pPKOLE/V1nRSyv/3Fq/mkQkj7c51
x7SxuL01i/houtAWvvpn4fmzlakE/3F2lDsgoJeJP1MeUdj+Nd40gr+KmaeIoK1o
VqtWvlCI3JHGAR/vKHR3IRSuIfPxTvondaoFvM3qS/XtVhriQNCx3j2pI9G78whd
0RwEyopzcnIwizsZ8/EWVbzF28Tmcecuwa+l17vIrlvASMG2ErABFoz4LiQzNtVm
nX3zUEuwvR6w0tSnnad7VBveonURc9HsMXvprUC2BBBG/ORHxfOE9RvBllt9rwBc
e69meT2b8XvwJzZJ0WnUCFHCIik8e4RBhs+4zySdM4pzmxIQFqgwbSt2BIMJhd/5
GxYwuSQY4qkgt7wCgTqml1eSVlQCBsorgXgTGmhmietivumPVQYd2SJjaAT81kGf
3rprl4L3Ga4m170HdFQpDdjjtrpSfKzHnbbW0vPbfB0/vBtyJwocwsH54Pna7ZDV
rfwB+H+3V/CNyf64UyknW3y3CZWTfuMqEF3HohxN+dTtRcx1n7sxzEXDIj8lzGI4
lcV4Jw252iZlzJOsg7s0MTskR/qAZY2fU6j9jjX09+Nd2mBcTfGqgaayXcRXqpZK
lF7V33KxDi/BmGp1lFTNqKPmx0uPXfk3TQrCWSc9l0jKtl+1ErMcsaRnrvJRyZPC
SkEpt5bgOq39Tp/76wajX+uUZPecJoF+QFFbljc3rAsgrNFF+C6S2aMzxOyXgTLa
gMgkUbm0AWLzcpQFs1gj+OyADEhXw+cAiI6zP7qtpUhjNQaMmEl2/oAdKn2IkO7E
8XKeYucjbe4484v+OxrjXudQ25oCHXVQkYH7jSZAETGl2HFAh62dazdy194gvEPI
fEEhemSDm3Nfd04LpCyvSP4neYGpWZ2LA+utfsrF1JiF70gRwnkjy1KW+8rxvGgm
8gYJrxLBM7VwOudq2kjO0Wma6enxadusGSdJAs+ARnkb8OMBuI6ZPHPy6CJhAlCB
3dsG2+yDKxdegLcvXQW8uKWubm8OgFy7DogQZkUpGmJVw0ZRWOXnImT4F64/olKN
karMM4/bNzV078kb85PZ2p5AA3TeyLwtNk5eycGqSLadxOscz8IprMXbcihUqbjo
1v2EGRw+RRNDWZpsrSFGCGDvp/fIUAgmWhLfSQ+i1SwF/IFpl2I4skCLS+0MDqS8
mWZB2z7EzR0P89/UOtJ2h1ib+lluBxKwXx0qw5hDqudgoVg24UqarDwpY5cLcoKm
WErLd6oRLGoBDwtef0egrxYacVEJcXh/Yz0qPT18QHdcBjZa5+kR3bAHD+NhNXBH
8WSkryCrPuGtFdfScsy4hpMsQ6o/AJ8TYYNrRJuPwODBMB8WN22fpqbvuHbZmfpv
SnwB9OPqwL+94ZiYAcBEwA5kmyWh1g/cz1TXGLL9iWpSASritL/VBLPCHkyoP9T5
bH3wrzc53Qn8cC5H7Vo7qt4hdL1Ni3wEpjtCzD78A9Ou/o62U9ZQawpd+JVek7sG
qiGmrM/JjuW8mX90PPt0Tb8ifI/kyzU8eEUw0FSAZHmtu3TFB2i2AIVO2Pj3Cboh
BGl67VmmzpgXxuj+UR4aXfwLD+At0ZNPPECPEnJUiuMWa4gL0IoQIMcY27Aogo5z
xRsNdGAZoqwIPewEV0Bf0uvTeRFfBXZFlS9ptQcZLF71zFV9+dXfHaP15PzxeglK
mEsEnVmZ70A/s6khDwNuSRwvyXPT43/hnJPDeF0vzRx4GdivuanqDiIK/bUn2vZW
/LOtJgRXH5CnW+JchelpKeiSMjiCLpZaMaVYgtCSbshiN28mt1y7oY3oEXaNy46e
JAgqlfxTPil2lhplDd30je86j8L42IA/jlVLp4gAliqQR9OU6WnbkhRlLr6wUh+/
zZ88fy1pMLHRmiedQZEStjDLtj82JQANwTN+4du822LNNgMVKnX/RGYZ4MbyyuMv
wjLaeZJLMI2Mia3IWhqmXrhuJWlYfbwf+18Nnbjb9tHzo6HDmqkNcWlHkc2pKL4B
rlbCNlOacEThRNYUyerYinSxchFVYj+NfIEKKnq/EgXdcZAUW+mnZWfaWdMIqLCf
QYwNC0bho/vcrUkXKrxgz4yWBkVhLG50aoA/mo5qKB85L/pQEFHKCmTQ92emNiQk
GnQ6vuGFf1GIzw8PXEsUZyYLzsXeXjJDsb81MV2mUb3imMpx7n6gh3a3N7tI0pAW
O6U7HkxA4isR4muNlT+8fEWwSedWIL7bukJ/ig1UAcfJKoXWcahopWn/j9xwjbWk
OFDv7H/UY8ljszEnt0wSsN+HAjbfj1OHsw+N3okwWNH5kXvskB55HuHrEGJA5aar
Xb9bjT/wJhA/vFrnh+zCY1gwFP5czGwnZU/wPU0TSeOCWQLxYY8eTSO4fAyiKYFc
8dh4g+di1eI+1ja5msJyV1tAxEa26au95TMDoWHlahKssy1FUmlOXtr0C2zDLPVO
+US+fU6V4w9mKrRekgbxmHsRWE2Dap1E28+G8u9/HD7MVQW0gHhCI1ibk7mBicp9
GDY1D/5Ez3ZGFxLfGparuQx+rtScjHD2+JiVrtZL9sKMOf7nJGAdwieaAjoNKniS
7IOnurNzf3EIl/T4Pdnm7hAVqn4EdZX0gOKlcWeVGPxYnYh+3ClV/Z6EWHjRjJb/
5y8R68Fom6zjf6buv+BvGHtrKeFTM6cv+zsBL/e57jB0WB9fvNLnvmzKcL7vdNAe
r8Erxc4bGUcfxgEXoLmKVm5H1JG9StElDvTiv5CXWiuo7bi18rjlYtw3QMcu/ROX
+JWEglIGmZWZSf4SGBj9lXhUQ+B2NS0xMDwgaiGf7GMpuXuVOeQfKKNJsz8ySXDs
CF8Aj9CyyfuoCY38u1kUq+WTocTIpUbDztZRJxauYwhLiXH9IojB7M65HzZlO8N1
Ihu5MT3u1M+thEaj96MzMjbwrFvIbLrZ91cLoXR2m40zY/yfE3ry7Hgq7eSNCyh+
Q5v9ucSAYnOnfGlH3w4WiL2aNKz0+X/odQZPfDcvLnSRATaUX+6V70lwfEkw+nzY
b4CO6Xz2520LYMNvLLlq7s0nSzWzFT4CKxV5rKFjj8ngjarPmjc/V/Yf2RT10rxA
c7bCu3xoUWGeeMgxbR1Eeb/chvtgSrFNZ+0yhwNipyXzaQDLoNBT4EOt3DITzI4m
26q+8NSkPY4pXZhShfPp2Pj55Za6wv62xqwHXBn2O0T4TeqR9UlDHQfuASKOZmmm
NaWJLniPEvc0AAxQLzEGys1Ljj+ylQArGhOrX7HctGg0ano2qOwDmd9e6/sVvbJp
lVlCCGiyh1vaMJDbTWY8/HdJ5fhMz1EbdDlqwT1dcT4D3BwWtAvjXi4mFiJIQRS1
T7xumXoSc2qWIrwkNpGVh8G3gbKnAW7X04eR9TqCjSn8rVdpAGb3/Lh7YUdYZgv+
xNUlZ8s6rPj22jBB8idwjSieLAq87K5/8NQ28EXHX9YK7J1AQnwULBSCV52t3n5B
ocUMXx7vMQM7geFNOwua5kR0eDoKWRQ5BGiKLffPuQS5QsjzhqwiJiHB85FuoVaq
s++uonWm/wQA6JW+O0uvPtlAh/yJv45keghmMLaprc2AEl12jw0bDTFBlZya068W
9WTbnBuO6r6qrbScew0Hsm23Lc3EKa890FHTjyHDeE1i89BvuxsJ/mLlXpcx31Nz
gCecvjLgN4DJUNgQq3nLYQua5oRp2qcAOybSp/Gc1/hFrIfsmIkjLaaM383FA/NO
WO5Vljlm8gJj5ZeXPtwQj6AQRMU6gcDjX5OAN9dU8tTCHZ3+49EReNbskHy6ro7Z
2ToryeQA4hRr+kt1jCGyBlCUY0YVP6SVk5xWJlchHMgSHl5jDc+aQzdNxbENQdTA
uxr+kj/Woi8nrq9gu7f7DvrBnf9DF540apBn9oJ2UFjGupArdbUdSkBmf658nObd
JPkVCBert7werpKAgP3LYdWcM1GvqdEsy8uAhRgpzVERg7QgvqMmPl+Lzp9IIU8B
fPTRD2cXYSx4NedOrWhYhdTI4lRNUEQxU3jORcL9PWbpYsfjrb+qZi1YKTRDujUa
AawJm6yMe24Veb9+jsVA6Uj9g2HmG4Ce5kOaQ0jBS7JygcfbhKEuVBqwqvngRBos
yUDtUCBRvo8QXjWclvj05NFIwox04t65ixKr1mMPL6DTCxlbik0H/K4+GfYid30W
d87JeRxZzstm1UyIAeaiTwS8FyQwQHkk6Pn8QhqQB7Lv3ZkLz08IDd5qM00Q0Bs+
RsllIAhRXQjHXH/Tqf5aqWthEkJoiie9/mhbcBTYpqRekJipSZgzbc39ri6wtd/s
gymSlAr0VyN1GxlZ8+QBaJnHiyIQfsV5qnbg5FoLyYpGnaCi78vGKLvmx/S4IHg1
yUqfEB+Ad/ogY7HnylNi9JUqZgk55tlbJH8O+pLx1PD+c3BeuQeRodQr9fLF8CrZ
e/T0deteuX64l/wDnZV60kmyN7UKPvoc7kPkLy2O+kPk80uTIPa8PHlzbKhj33/W
FsAQEXAhQuaBXknV5lXrC5VbhGWxx/5Z3JcPzBK1npmYe3EK0Zn/MhzuobVgLFGM
NrXwCwHv9J4EJWdXCUaiFPhIJxNBGtCktjUk0vBmkUcdtVslkF6X4nfaj+ESd8uG
efOnucIEKEgzN6BlYOsZh5+uYP5r5V0Gs0B5uPi20wAeVcIbOQr+NEc3AJWGdsoF
f5jJ8NIsawBYW325N+TQAHEUWtysnb89KBL4AR67u1dqUITkAMGET/QYA3uk2nyu
ZP8C+CRN2RYWXMpcqa6tKo93SztVTTuzTIfyNLTZJ6Jadod1LrPQAtdgIG8+3PIS
hX7HVoGJg/C6SsjofbGOtlqpNAmYRt53Suo38nRQu+PMy1jPX+WIZu7hHuh8tNnu
xOLSuwKwoOnM3owJ7zYfzbMhQVBmaTkISbCrRnq3D6sxSMDizv32dSOLqsnV3583
FQDWyhuxilj34cFKpBEAvEwI+Fxbd5fSIHlfCffMSCtL/u3QmgQb/vzclBSkhJBz
09gH38rb7tGnFnxiiW1o+gtmc6iJWfRDDUq76vUuvwCgacsgMgjUJ8oI2sMi6sbd
QsH0zAYYe890zpO+kdSulbVdWGvZ85kZdWowvRzZgsIzZJAZzrkNaegs4T06GGma
JK66HnmHNS4dfHiLWtYKcQRZf7YQOlp4L5eWIcIJzwNDNGPzEwiaq2j15iLG9wNc
QP0GbfAqTiLuFJMYh8VY195zmP+VhpIUNbR0mQejxpgeV4vNuxnAnP1bMxrgyiEB
49wZWLofnyIScfUyhiqMVUgXg2AuoqCUD7UDsWNryAmPa0tItaRxIMMjG3f53zf5
yyB5s9WqlX2z6bnhrrK/MTjzXmuIAMSSvZYEOJd5m0oM2pym6eyxDFhHgxH94n9r
JNB+/hW00jaYWZK64eKQSGe9y4S65fqIWk69bx2abIKzlIpx4Ut1bIatD3N/RK2a
MaQghQHxaNbcqv+bOCzi/IZGG/sPos5guDekkROobCDLgg+ujhuiVEsNZfti2GKq
ytNfLIEeCZTz4968qoBWmwjLK0YpTBwONGrsw8m5R0LCdM+vidp8EQPu6sVgBkDE
nqWCS6K6GT8Sw6W2XawvtxRxkHuUyx/F+a6vqmrM2P6cBo5f7dE/tVT3vdN2t3cy
kNNHVW2hHQdle5Wt246eC00nKGwnh0oi3vfZfXqSE2hx84tnmyIPyjVBhvFVZmwI
9uzhz6d+3DvYoVHwV+GrZM5jdf2O2sS+46y4IXjvyfBF8+G/3NYFc1uGL/ZiKjDn
Nhqz2wWsSCA1O9q28RpoZQekCZMnOjJgCIZcIAIws73iwQ1gfepKLNlYEImBIF1+
oIYu9n1eFMh6JjGrE+UmCiRR++MqdMf9Nnc6oo7QoNyExUKR/jNX1T0mu2NOcbrj
h2XKw+eqn4E/2lpovt0613KGszP6UoNPEHmgWFw+2EV1IS4Ocfvk+uJ8eOvqZvpl
BBRYe7B3GyvmTOVsa9JKGVNkIxdnfKcNQ0eitDcse+PrIsq7+H3/+oNUt4xe3XSU
d8MU4BaQ+NHPRfGHyJNWxsGza9ra25FSuaoSQuEyOQi/NfFDgWfCdwOv+hift+bs
t+UC8xNUyW/fkux/on4WN8ECQhKT6UacYa4vzJET2fOr4d7jm8nWiVY0+8ZEfYD7
uB9dKngXA04G3ZhNs48R35zYXXvOy0BDbQw+XsQrO29UEzLmP+SWvCtx2JwbQ7rl
hAZKLt5wiXuD+HvwkBaoeMCW2FKuJ4OMRjBAb1LIep3c3iGjjlB116ExgJun+C8t
hLjUHt2LLDGUTVBBRdHlBhartlW7Ga0HBOQ8ZcdXArUE3hAU3v19pLK5UN3sk+Ik
tBBii1WJU010fFWL0xnjwAIAmPDctwTxp3UJWW3zEGHQesF6UV4DfRRHrJcawGv7
KNyIPSXVrK4qypemPe9Bxwc+ks01HYvUB2mBPlnr0gsSFGr/3n0s2UkaiKM9vGMC
QsMwxEfwAhB7TY1NOa7R8BhE/z0rNABfHXh5stYdBvcQoKdUXrGHi47OcChPwIsq
/UMoOtI+3jf0c5NVmcM9i5ENrDV33Ew8mnLRFViswwR2ztj5sEhZ3/8XjWFkpFks
SZDop6TLLX9jHuG0IIdm8VaIk5Ac+VId8KCB2Tp9PnjfBXwxRAT+70J0gZ0h3rmB
KOckqkE/U8r/VoyHmamOGhCqZ/YbZTSsHflM0Kjbhxt8N9YwCj4za/xpJWdCE/Dq
Go65f1HUNH8HH/LGvbco1ggUn5SPerJzZYNVJUXDJrc3n9sNz5j6xYEdMGfonXIw
TWMbfx7H1Dhia/HtLiCYws9rF14bdL744COToTqYkLMDMi5i3xh2Z4/I2NOqDR6M
FvNAOIbNyOAdU333v8nuL7TRmdHLXZT5Xm7+D61NIeUiL2Mp/URFDr7c1tWDKJW6
SdsUaYlZHMnv7asS3kbJvOTaUFwKlhyofCRP+hNzcqlS8Qlvgw07JXWfu3Ma4J4U
447okPA4xumvsrJSoVnl0ntGMO63qwBHr3Ym5xvKzviPFymQSW7/7/ZP2Ynu43mV
+nO7AMTm9hJ2nOfoFtg6FQYchpIYnImjuzuFOcFEmgvKnARFDmRLM9r882Oi5rWG
bcCikAI2jiauXwvB3YI9BLxVs1ndYQo/9Gv+n7UPIAR2+sW2JknZFxx7FWub816j
QuDyhg5llIt2GkRoZZszNAu9IanZ3wL/6OBahse7tqpxE6GvKGU5oFlLbJon5u/M
3HC6qAFNeLm3OJx/67bzJcokAdH8rqIDzp+m0eGHB4YirRBSh+rWfc7NYmkkCw9H
npjBfVvrbfnRHC7zKgZ+bhiHK5F2KSyhlUhIUg+FIVA+g+s1Ro1t8ZpMd8WDlsG8
URbPvt6XmeNS9DCowdtMv81y9a0vYzQu9uNEdyu7BQpWPnXgFSl9NY0Id0hKJ2+7
aRIU+tQA9s21MyqlCjtGVmT3SG1fHA4JB/rS6tmaUMgi0zfsA7dcclayRPk9awDP
jgFW8ud0cRg04ppbQ0UtZRtBfOs3h/2OPglABbhccAoQNdEHS2Ki8NGQM8aWcrKZ
6v/J22ZI9XkGxvvF10hLT7oe85FUVonS0GBS/E+2H39s3odqZkRMCZbhR/V5E/ZD
SgPs6l0HADG79+xgCDA/T7Wl9Cn2UekCvBXe96tK3C9fE+Ube1Qz7o4uXfa8D+bL
JyxjCM4jH+rtCIe5fAn+4MOZWPPqk5lOy07bjJRA/MMB/o2u0fr0MnHlVTwKTEqz
yHrx33LkhY7q0EAPD2EIs+hT0DrtP3Sq73wQQh6HuXjLf+YqDfky9oT87cma3g/b
r5kOIUYR5jj+wfqzpcKdlWVDzTcz2MgAECVKlCFxTJPLY4Cb5XwykRO8SJwzP9vE
UAdp9KT2j5xz84Y/e/2F6aXMaQ5YTCu/uYdU0DEKQhg2cwT6stsh4guO1K8v5aQ2
TNpQZbhMEIyA5KEtU22BU8Z/IfqRk61S9lLhz/fcUSLam6fzCC/xqjCO8Wb4ZHyN
E8UWIJ36yFbPBviQFS3FTxuMxuMndhTcOLlXHXO909GYzNuzyY0ub5Y+4rUJHtJq
Z6Ui41et8nJ8vd+oznYC2sL/+WlUIyoxYHDPqoiNywfgGufGhGjtymjiEejNTNiv
vXa7lygdEb5dQxoAxi4TLD8jsQwkNuyFaYHT8IuiPk4KZucrHA5cWi+Z+jfq5aRC
1is348CNxFujRKaMy8LWh+Bq9EqYsRKK1rPdgh/YrICidd1h/PF20nhEc8xHuScq
OYJxTchz6OwNIwCCq5gmwg4lw++nSsvwZCjaEHu8J47z7JBR47CYQKuG7VLlYDiJ
XQF0qLTXdPfQpXI1+8sW7SxX8avYTq7lKU+TS+9BIGViiNX/YHI2WQFt6eYM8u46
428WkT7kc3gnHprYZcypFf3C3uaV0yLNL7f2g2rE6opWFckps8/gY/8j1V3e0k3+
l3m5FPR5jHmi4PIJHdbkICGF+RlhNBInYtCIFUSFSnc51doqrk+GExT2OAA+IKum
lPsNywhXfSvs8WEqPTO1rRKflTCIbZnX3rGdakaf3+Lz8od1VkHSnbIcmcDK6PZA
L/cwBNJId9F/9lTgJtgHWZA85twqfYDscmAQlvM6P+kew8mTG5EaVonQaoT3fIAD
H9xyGjNC4r8XhKfFW9Ns3n1mvPiE8TqhFbe5u140uBNjxHDwIHcD4Gwl1t/37J2+
g0AG4lv4+GiPX6K+xIkfooKth6dD8AzFCDkLuSSnyp+nkrZv/idD/kOwnKkPpytB
uZAzN2dy5sHaUPaKQ883GBrzBxuwDuVa0iPTg2tMeKY3XqUYbsRe6Gkh30Yq0Lr4
zyKLgL4IDwz2g9i0FCh/7+KV4TGf3WSK3sYwIIcxF3hRyAtTltGJtVdevAePWpmy
N6QlaDMvAAr4JHxTwW0tQ/ne01BlPbfZwsY+8jxrBKm9FXMa/fG/QaCDw4O+OyQG
OpVOUGTKqU1OrhGjS67/mRg7bkZLryaRMBzirFJJJmlgo8hegPRE1dh30+gz/NdS
LdUsJja6OB2leEa0X75vEhMOVnFnrldjgT1+32B2ZHpm2HHtqQSzfzC7wUdDU2mj
AUCqa0iU/i/p+Imo9iOz0DV5vtMlGCwm8NpK88PmG9MAOQoawJbyKCkRr235kx+n
nzg53mMQnus5mW+UG4HPA0WoIL8nPoRu5sKlSj9X6yFOKCahbH+u4gbSgp4xP4oc
dsyMDXnp8gdWQORZf6leCU8BFUlyVHaeGX3TajG4QFUHJQz7D32qu5n0/Heo1P/W
2w/l8Pvluhq2/gpAUoCNlkg/vaZCyNp74E5M09qGLU/KyspQUP2AqoTKV4ZCnK8l
+Ht9qXjFvovka3vyLZodO63/EZCMvsp7PndqgYEbjfDGUXLoHlSm1J38XaIf6duB
wQuIHTfxqQlplK+Om70Twzuo04428K4pROaSGi14EGeFKlY5CEur/DQYM+5RuwIW
zJ3PmM+DHsNFco+eCtXHvK3n3qDMwWjhhfGp+bgv5L/mDaqUVCa0zreSrIqtdW4w
RGyO1QxUbLpb1nwBGhjEGDMYNnV1NFJ9ArRcxaf+/grl51lz7nJk97cboS6u4lkL
/evRWA2C/hJ8SrAwqiS5xjpbrAZI4Gm3IPQfVHUG/ihw0ePpbRI5ms4aewZckeSN
kFiZWB7xI8XWCUgp3wm74HmjSBM94k08vuv/D8rieghfejRZfPmIBTREM9FtnCot
peirfhryX9sF4Ilm7vJov+csU2KFAIRqbWZC3aaoddFaHyUdMsARDog6uxI/kyUq
RQ9+eC50ItmGUxfVWNei3oXpwI6gb0zFrrCU/isXMQFdWDE2b7NA9FjeXaVYyVwN
KFLt3IDv2uAfIthLPXgl2euTykp34n8LS5cffBBnh5OkBOmRlWs6AMrvokH0eFmR
8aY9tDNGvdxy8Zz0yCXHYDepemWhG2ViNJcHK5qB9MJvxy+vvqAo3gecxX21C4Gf
nhF82KHh9IwHKSyLilPCjn5fbGDe1qUUzfCGDpJeRcTMbr1G7Y4flw+UYPm5NkHm
gJHIu8qnh7nzuUZ00nzloZWBypInSiHQdB48hMPEDSFNvnfZEtCvMCGROFLtZSq4
u0OlBrqAtmBQoqrISTDhmbYyuHOSJMrpdyao3+LaH+cNNeRlZ8UoDwptYPXr0Wia
Snj98tLN/mVuFCJxuD/UsJ83rl32lcK08r/c198i85JOEgMHSWyjbgjsSvnU1tNs
VdqMwpP7dyXLCv5EOt7u//g4rWLVmYCohq1oSJW60fhzSivJaS1XQ2xUI2J11NCV
A2WSvawX/h15We/TLy3cgEwNF9AYOPLhdLWJX3gJnPu+qnO3x1wZFbYUxM69deh0
H0/2j1TK2Dc7ISdTkKsUE7Tjswfm9gCOHfhidG6zipRyn9LsLWsU4cxH+eQosB+U
ZU5R6KQ6yJyVFQXNMcbPfkD2NjZ9/Q4OvkBoscKlPv5i1f2OnFAfbB9R0d3grjVG
wzw59BguQ6RpXXUrwG8/rEyxOjp/XCmlO1BPfLatTRQpAWU6E3/tVrd4nVyJg/vj
Jl5viIhsYKA7itJhO4+KCLRkhrNrSqwGGUTYM00MenJfdFz0HaTiEIjfDWA6Bfwu
Z/7AkuxPJU6h58dUZLjB9HZVNppvWGJxsjKq8myGCLMyoyESGuNnlwy90GD5MsLf
xaOPYzA3FWFetfd6kl1mMpMhG3oNIchnedmXuPTo6dimdGn/bN5K1bMCuhyS35I5
slO9TjLSO3eSKjRHCiXAauy7/t3+UwRrVvd0ifNOs+486eGGzC/VZ9cHEiseU1p/
ASCS1fv6VCd3inZkD1Rp6DNIbc59CPTblRw9rRcEpXeXHSrj4Nm3dBqA9QywdQ5f
+YXT4a/2K9YJDdfNUVPMNEp5EYcyxpnOWoqZMFSqsOGXhYGixkY8KnIr1YK5x1nm
Wwa43+E2EJ04ZY9BJsGbmyQztNrWi+ky/MbxjB0XrjHjZNEg3GsB2GAcbeSQ5RgN
5oO1f3AHtw+yN0lDMtxMuqlUTGqCogI2RWZl/3vKX4XtCJ2kt/bArsR3iflWU9Jm
uCNFyufVM0Rnv9lnqB1z98e6JtgWyXnFnXmJnTdGokf4XguQsNph46wS14qTXZZB
xe5MHQjF4bS/wEqO/XxtpTZuGpM7j6DhudnFeNBOu0eTSkjBDRlDLIf/yqus7s2Q
JbmLYhModhnEf8nc1lMNZV0NTn7YVsNZV4UwoWoGnIWyoQitTNa/5hpzdjFKeCFN
YwWe7unqt0utLhDs3EwNmPqdvuVRMozg+NJO+YhypcyRH5pk6958mtV6A6IK1+cD
94R9U4MOfFV0B87ROq1bG50l5PwcCz8Okel5ik6HBBCate5R/eLe0XC8sMMDRvvW
d/AL5eiXSy9crwzXiYvvgefbgei8XR3hG3ZgXMSOtnoEX8c/xpRnzYzTFMi/Z42S
VaOk2u4Q6zaSw+6uiuwRZHlhLqUra8xVwgqGGPPlqFcFhmoBS7h5AOOSnetv2wSj
muABB5rx4tR/VLCP/NyJ3Ylouf7B2a5OUtZTDzaVIRSKfihAMj/i/6yfy/De582s
dcGsQDDph1819YWVjhYyadZfZ4V3Ek48+Y8Wyy57pJWZFmcaLyTg44OxljVHY68u
1KvwHcT00maAw7l5BSaCm4w/48EmeNorYUh8c831wVg3wP/KRsLB6oWCW963c4vY
xML6t6D27guSleJdnfB22hIbtcBf6lVBMNptaTJCINCy2piusEQUoAnXW/fn4AzD
pEaIxQZ9QxczrMw6+LROQzXVrHsfVehgqG+sq/WQM9G3l4nENVKXd6EhhcQz1FVF
ehZxqTcqGqsqbq5+DH3CWbnBo2RFDIsDMUebVqMF/BVlopXs75W63V4D42p3jbTZ
FeYDPftPTMfyDo1pRPkeLDGQ1T07fmhs627Rs8Wp0sL7bf6k3JMnHYXi/vNSXxGV
GK1yse/bSXwL4q1m1LAIU6mrsGrDBlaYUutsHSnwrAFHhCRsz40w8N9P/lyhbkXe
t8d3bJN8rhEoBx/scvF8Sog9lBnnxO616nEfdBJgJ+7aLTYVZdTFyaldEGbftbKB
szxqb1KMLFlrDVLXe6WgvqqPNfx230X69eDLUt3gSXhA0RGgWoPt4T66ux7/XOlQ
+zCtzcf097yXRkYWod/piRsM0ZZ3Tz/pBS9YnTllT616Q12TKHW8OUHgOoHxpPll
htUnZeT8RIsILC0u+bImk9qDfya7yPIioFHJCi6fy00teSE+zOzjwzB3+RJx1iEX
1tbqaDnSe/P322GjXu5tpJXbjDwCwj39Ku8pFd2QCgTrTjPCKNvXm+WGxSukYpB1
M4jNYS8TYNJwojtY4Qw4tFI4DkaKA1I1lUFfAwKqEelXpd+AARStNGbj6RU19yGP
6DYdaSVIzBqKWz6MaYg+C2fOMAp/Az2GVvVGI8qTkEjpv7SWfvfSkRSjZ+DoACHW
i2oN3qLLXELVjg41ZXdC/i34kBf74VW7H15WIA/V7/KWYHmORgzvsjfug/bl2hQD
4Z/ZZjjJqwcMeTTymmoteJQb20lH8zdKIsbuhwEwGCm/7JTBiW8gLKddngpuqa7p
vmNWXJaDfEB/7XU3zcO/l8qDmC7NK+DU7wNeHVC0iwoy5k5zVvExSGnFggCqRBU6
a9PWMaBFhSnI3W16ZpK9pBpY8KlD13s/gqLkZ83dHkpjTZIWSubpBxvLTnd2HmhI
KK4vVS0sh0kSGfGTuzfSjwZZAMBFvkAIqgli8XXjBRcZsE0p8ZcP4vIGWatDmEBp
MO+2MyHUXVuIpfeCPflvSUHGzMy+pJoXzB+s6PidWVGJQNVn/WtPZVDc2oVvH1U0
iRCH56S+AjJgAJAbEkFvGF1p3wN+hWqoqHcPRqFMq+81P6vNlravgI8SVh8GpRuY
+d3WjjaVQXxpypxjdSgTaac/yFe8WHlnghztwjrbciqJykWnTxbLASk2BVSFQGEr
b2HPDfx5CLkxIlts01ssV2sG8SpnWaaAYUTNNUHzr7+3AUXeWSoxTs9fInf1O+KE
dNXJ81EuP1zyzMn7z6ec+IQ+Bsv6ENTAEYDeoEhDb6uUDn60FW2TpJj6rbDVck7h
4tShzPr3mPwrDT31fOt8AwJNk0kkMQghRvyBzgZkOxTdTGNMFM7OgW7Sy3XwKgoy
MJKfb0r7m1b0QRjNygTvU/l2mGL8bD4c4xZ04gffcDI2yIKWiOkMkdFY3iFpJuK2
fCwmxIFB6h5LIqKPyUyg6n0wfukeU+eIePbkho1cJPCeLPqikNgRipV5r7TkDGAr
U2BbBiYaV1coh22mOMGGP2SP50UvhFBxA23dH9dz/zw2RZ5Mb66X0GmWhqErh/UD
LRJRmkzb9JgljUJG6gcul/iyiofxeMvvUFan0BQtKQKo8kEy4L8D57Zqa8//0Dk3
Ngqj9Ncee4ghYDaScpW9r5T2mrpg01YR/IBl3giSQZeqYpJKne0jDkScYM1JNzbT
n6graqJuzTXwxvhmInDefzi7wwFs3nxK47FKLqDIZuzUUwa+K1KAfVZ+HfXpPmUG
/Se/wZxTiyMOAlxmNcTK+rZpZw6MFVzPXinUrmDLfqbaTKzYsU9XbHJVJ+IzHOXO
Ya6TwDCJLuy8vU/8Tp6xc8pIy3EkV5y8Lnvjs+j+E/sdl3qxEan/jNYS7W9rkir3
pGTyv9D9gWoBaZlpbraeSgtVxzFFQlwatnD4OhOs9XhSiDrFSGKG68dphqMCmNen
Eh8lF//X8ySdGULhs+RPqdkHV9Xuz/4p7LtUI6kMDYYr1TLAR4TZD/4WTzTK2mTR
eiVZy3Ul6xsevhwJdM4DEP3wWA6t//ulqgVC1dWNhXMyNfWym5QcQP2Ay96fWQuD
iLXdovYWlnl02drFAhYftzIbhYgKFn3UYTSP2P5YIxrkNcsTPQQ3hqCP0DCE0HvU
v1pbKdQqBFi/QsNi6TU6wN6uJRRKGXswCUD1CTknt/xwKz9kqO5OjdhExqtBpMFn
YXoRECb5P0zTz/iuqu7ZU1FI7ClH8esbNqN/Z9R2mpr6imHUnxkHikFUzE4FnDmy
cXxUFxIpM4ivMaeNgkclgUQyypnKhagRgxzs/gXJ6A48GcAG10QIT6pj1kAK4fVc
GHrEnFvtaQnO1oeM4p35v8qswDDdXtotH7BhPlIpvU7dP/cRZ/4f/Zg2bVaKJ2Gx
uuBThHOEZfkRgeJgf1gHYZbafnQfp2K/JrC6NTDpTVNs+YTLSxaz5jYXL7YeQXAw
GIVwjxQo5Btv9ObCU0E15UJyhs/JvoWSc3nyxDnVE2QS/h1BhoeuF3zJ4UVwD7l1
/iOzbgjXteFsA5Y2Y7BqvaZ0Nyc6g4vRCDvK0aHxu5kvUIQlyF5Wkz+0xcYZDyIu
YrYC/o4dDe/kIn5Tefy0gjGhi45QcwklRHgc6xnl/F6NUjF/WLi9KMNv6S1xRDeR
EhOpY6nl4SNXK+sMmB4tDftF8Zwd4Cs6a+ChjCN+t8KaSWVjH2kpqcmesaGDGH/S
Uq7sc0FcQ419lycpE+YfztemB8B3IQ3seRE3Z1KwICKAadjx7Xnrzbb2rwM8VPrQ
PmHxzK3skWpMyCY7KLhhh5vr3dvYVuPnwZzTl3Zv00Qq/54fyF3C/rs3Mbhf68J8
rAL6VknQqCOD0Ph9XTRzEMSq13AIF1jVNbMlJ7PWVj4+G3MRlYVl8MNyQ8gYSWil
MENcv4vfyszbSdJOdwhz0cD1jnOUM2ndFnpYnQFmNBE4N97XJkf9/+XsN/qe/DmE
FI4uPPDTw5PJiEHVMTCLvKjKMdpPfYSjK8vq2B3wm2ZXd/Y++snXz5xfgondGx5e
pPaAGvmn/rw8124nSN4Ag63cvs6/rL/rSI934QqA1UA7R3qfVLKCUTHD/fkAPw1Z
pbd/rJ0oUYvSzeSQroRJbuzlrre8H1W+5uF4SXEYnUaYmMN4r5MaUq2V8TXARlFa
12GYPoektFMKqaEg4+ooa615vQg2MvDbepItzA/GqG/2E42Y2rmqD2Wa/X7/i745
mBYgT67InZX86FTKH61YsHe91ara4Oh2KtRoepNaTa3yclwvB8q1l9PkHXG2JlUV
ArFrXyGc3AhaZmIU0N67W5lovctXGM6K2fAuI2yRiDGQWOP9den6brEx6zDGwcPY
yxvseP00PrPQ7wNNDASJ9tjis+MlQN1a8wOD1k5nNNjowXGUg7wl9eR5e2KL5cGN
KShQqCr7raSsLXV6sIFp91+YIuP7C2xX7qk5mBMexZf/jvq3dS3KvKWeflTRPKzT
dPUtCfET0A8XqzlyqTV0mit7M2b9pJcOkzfB3VQ0Q+KNen58yC+qUV4hNyF1GyHo
xGZniZz5hSOdOJfXBl21tNn89TMTYhTaxSAPmAXhk+WTjjqGsLp9/oHZfycVFiwM
ccO9u/BW/0y1nvIIJa2w0OlxGhvUe9znNYCJuBpM7zzZDF9FmfpyoGj4myf8NTPt
6XOWQWNKwibE/+dMeGS3BCyZHrKAcVlyA61NldA2reHm6QU942x0dsNLzMghii83
u+3mQ0r+MXMn4wXis/xUZSoAMQQKS3z4A7EMR/uDIpDceqPtKusNB+S+wFWly6lJ
LMIGDpGc+uB7zXCKOlsFvDL8OZ5SOHo/NQVsTFfX7qYlN8fAyXa1FOR+l7UrJhJ5
QiAfqAr5Tfj7PxTdPXzAvGrvv4ClHEG2qHbA6SsHTnie1o80Rub8IUX6z+gZyPje
Aare+ObEzWHA/M2K3gmbzy179NQtVoSbnjUElE+7oKB0X+bTYXyv0EJFXWpaw2k8
OBDzjW5pGh2umDxAPeeN7Fbiq0BkZ25UluxYXNvEMFntlokyGNjQDeGPSvslEswq
qkP1wwmy+/1MYFoewQ/+9r8qwR7SJnv9MlrYKQLW4oTrc9jgun/+fzeKjp/H2EPt
UlzVb5ZW+OObCVD5d763KGQQm8lytohdkg958GWhvbtCSABFEIhaAFMzeIKrzbf7
CY+4EQWnWbydG8UAy4cXMtsJwBpR914QSCVPWcEN3lrKc369/kT/D1bsDQqAgyIr
UIeIOHitTbOej9KGBSr7lRcNrrfWMNn/sOvtrKVzXKQwlJaChAfOcoi0lwFIh/NJ
7zjfx/2CMI14ScbGyiM+/BvVojUafDriIU9VP728XehNqfrr33lBhxHtsIUyY4j8
LxzJKawmjcccCSaBgtg/H/LHB7uSH8pMHLoDxN/JXBkggqPC/nUpHc88BoMNTcfc
Dttr7hCnuMSHdNAKBMEHUp7d7e9bzCNGb82RwZ7Ewr+G+124rGmS8cnWjF/2CUgK
UEps4HiAlVp/tPb7yE4AOnT04WWHj2Pvb0EB4Pod9Eovfsgf1CVAbsBo8K2RcQd3
HIKjINZxXa3/wOGllPTM2rZm5kW6gTMxROe4Do013vJuucZvq9tvKPtUI6YRJ218
bzgwMNjwt+vZhsi5tASurSjBjqWXBKKd2P5eCk2kImN26LGhcJvAzOSRgIeWgtkI
DdjlTp9yXxZJPZc1/1uASt0q7116rNEOo/nIHrLVkzFlt6do1Yy3PPBj+OWaaTtq
3WupzHRsxEjZzq43O5Sat9WCkBiVJ+mMuHqZurPT4GRPM8UMVmTg4k8klOlUgg21
hukhdLGKM9eVOCvV1qWNPrDuZYj4qxIUUZNb1RjdbNmju8UU7YMzEf4Lh/2F+0BZ
fg5xWcVJSQVyYd3ou1kGlSJ/iPtTuTuUR5Li/RbB34kLvNgsS10iUYn/idkNsOVf
QSqMWxxCeg7y+oG8L+fmvRyQc3TrSLZUXAax8SlX4KfD6ddd0zLdNnHcihlsROns
k4k51Bnv14eVDY8sm6ep/ikMAQEpz+35da8fw8GszQrkCoY1bVCrH5X6QT4vwqJM
n8dXCyVvXuYq5Likd+I4vfZ76v9bHzNJihKr5XCHDpYu01/XWiHwdVIKkWyznzkx
U5POcJ27hOn3SoqxkXksHKIEpxW5MXDeGN5GuN0jWsXrSefnEi5rGJzDObki8rMZ
d/1AM6RJOoehh7ohiPfnZOS5UC7LkMCB9u1heJ2ZcTdVsBrbYobMEJydF8MLsUYO
Yx0Hy1O+Gf/zrOrlyjuc0n92m0z+hmozCIjUPVDAzGxX1DJ49h/OHbodZLQ3htmK
iZp76+KmBDh/WY/YtHTtgV0cSoh2wDNi4yQYHPzMIi243LUsz1qknqWlh/uvANCl
rlnvI8WerAGHxObSNU64i120XpdLZa/3KFAZRYGwnxnIM7EGr9Zaby7Kq5X+oxym
L/g0frYsUMj1pq1HZ0LLFwPJCEBVg3YP4W4VEmoP+SlVWYUg98rrszKlyAvXi0/t
bbPtEtt34eFCoUb3gvl/V1H1BsA2Zl/BzuNNbYJcxW2BoFXA5EFILDFhIN4VYN+r
4Z+oaF0+AHqyWwI0Cj0wDHRY6ESN/M2iXl7yQFsAqkuxkuJi5grSDUKRaUIFYj+G
q8+jX3/yx9i6V3g7koHYeJh+TJaZ8Q2VJi6yruF2MUWB2a/xvnbFuwlMnV9wR7oT
fUqVvTOSvK4fxK3aW+l0ZTyZYsYz9eDn4+6af+dbv062CF2l5flLmVfuF66ghUcd
OuD9pPf/Syp+ZQSdr4b8RBTVpimwieFmjdxuVyed9U3a5Nk0sukq+rESSMVJrlgq
VjfBPSQn4CTcJe9kGxTcUoBvfJaLv1xUTTiG1F7t+ZmgmjEB3KyOfhXKosu9aIDA
AOMq1x6tjd3NlVKi9YpMnKWLMjqloPuPwDaLYPfM0lLEVn3R1m2E3jhZ3zFDzj77
2oXix9LkFufks2GU2BE1jLdam0TXlMm6LOHcw2+aP1NVNhjLwAdz04p+qdo1h6k/
y/FqyRdvXqvBeCZUtaLqOeReVdw/1m8IIxNf5sHfmt0dOslIsaNhW3CrH2INsWqc
HKJqVPziyDDENI5AC9IyhJ7puc1ut6qs23fQ9eWrYEoTS/21bgTwZIIna21pC2Hq
+WA//KQ4GZBLPpr6etM1IcYhPNxikgqN4wr1rxnspcHO4zlcX1MFFqmhuSMovyoc
Ru0mm/tET9TMiiNRH5VJIe55twr0+2hxIuGxbH9w+URJ91PwB64oWETQjccFhjLZ
U0QH2iCItLssnapBHPVeD4N0hWeiU2d8Hd9YzUm8eDDVgaxjNJ9iWJSomoTNfVpw
1tjnYag0Jymxqo63q2MVMfx0m+07UVolFJeC0ImTf6qax6kTxPRd5ZsJOEuyj7Nx
zoPzw4L9DRXEvbm7WpXlLg4UgjlpogRdwwZzRaLpu4WifkqVn+HK4JTos34XpijX
QiHIZ+8hyprOeuYG64r9mQlRRHaKuKLGSHV5ZoFM+VgSkmd7cljZnldNRrzNku2/
fCnGXDUUmx0cq9AqV/z5l1Y2mqa24rRyo89W6h5FXJ9/8kdeZV0NIcTvig9dXOlN
oyuKZCJYV6x/KzECZBTuuNaypValjm5dIwcB8dVoS72hpHf6hMzRw55muK3WhT9I
WFYN9CV8oXCtGBNpzYG92N330BmJXVzHqrLo8ZgWpAg+A4uxubcXvhrNDiNORSQB
qODZkFVRBDLQHNuXI4R2A362DvRTBI7GY12mo4f+P3VmWqYAlkvAJSqP3I4DQli5
H1DLm6iz4ooiTigD3vbABLCT5hKBqorJTvoy9QHkGJF3FbqRDFRrnGvUddHoedva
SdP26Jox08R7oe5UBJCKoGuS3W7rqYBwwiI5wMa9G9dG6XlV3yPNFD6oxDimVGpX
ElICb4tI2oVjG8HRpo1jejJWpY6F1Abl+7DMlQty18mUoBe+14t1mG0R4AgBLy2g
k4Nkn+zEUZMw2wKzGp7RD/Gvwb0c/CwS+ZR0lh7GhuH/Kyd9ZWFBfcg+0ijeEenR
SV/63MSSzJertrXeV4uDVLTB7uFi9PjwPBPJIQfw3bXFrPGHO2eczYkkaBFfAph1
T9C9Th1/HKbkN3p63a5LjmAU66TRzgm7z8jJVEjodvnfgyRWSIAbJREEBufCVgZO
6ijenBspV+YhuQRIhI7kmJeG+sUWS79De4nzI5SlqEFPy/w6GDhL19bdcQZ6fsGI
WJyv/VwJU3YVUUymIatCJJhaIbJLm0MmQQNCqfpHkbRSwGTL2vFKeL8XuRoXXad4
b2TfgwpmEnh+FCk5l0/fI9fPaRwRQBI2rwgIYjq8xhXsJBrkssRh2Q5DbuRaueEP
MUk4j0NwS2OIEv7D2738O9n2fypUYhu6/qVNbSxOOKPK0DZODaB/He7G3xYnKWN7
4NEttTWF8YZqGBic4z25wKrO6j4tB76hs4F7km2zV1xQPva/2+qJNbUQjv8F6KyV
LyC75KCAaRaZB+qEAc3efNe1NLJXKEiXa4Vv0aFXRI1Eep23HGhzRyCyaZ8E3t36
P5Ae0rbSD2OvdPA197y7S4my6MnJzDXUTLXE8zDjq0y71rDlznx9PygXZ+Z+H1GB
ecGgLryXoVrnw6fIcfSlUFtc0qqcAbEYIIbtoKtauaUgZREH4pYq2b7N37m3sJFb
mLLyWWlZoZNHvm3blRz+w0fbujDLCtJltvpkMGun3pRsYrYRY2+0tnn2MtZhOcjv
2H+MpzboVruZrILUWBXo0w95eof9YpnsxXAZU1dvUE2oBQDqwZR7rGdL52y+7qnj
IZQBxqqdRClC5vHCh44uV4NlH085GWpwJY3dbRIL7hsHxFRwCDSj7XN+mBXi5Vb4
IvBxAt5iYiQlmlkU0BIheV2IqB8ogwg2x/I+RIQ18uI4FiDE/liIl1UvWh3onJ9I
HlvfkjHMOCFfK6S9QYggb+Va2twTRpzkV2bWMWbn54xJtVpfLN7RTRNid8jJnLcw
KH09G9PnBfxpWOWBsbVZwGstPw1MI1b+DRkaVsh8Eyd1+QvE02P6fYEB+zMf93TM
Br8xrdTFr+dtgX/xbPMHRUjtB5Cmc6WDoUMJPbdIv1dSmN1KayuFlkSXaaPJDtGn
KFHCBEgvg6p14ALeewxXnghT299NzMTj+JwZVP6i13yxGO1/p8oePqHBmUiPpCg5
aHiN8C3F4ZVAxLLSpZZckJnCmlNbCpr0uGUlP0+b2v/rvWMn/gMXqI9a0yUDsmHk
huliajAQadksZlEzORqoTabZyIbamwdEWAjA96psYD4pZnMqkjmUvnyS4qCT90BN
59IMzLLbICHg8Bs+BDHNxcLfU5Axo9XrmbMg+POur40KHlZzTHb/f2gLOd5WJN2N
34IjAI1nKDT7KvhnTIw1MB2hhbxA05BuGnxn7eVin/e94aPiNp1aXiC62jl1gpgK
iG/Mw2xWBxtKojjHUyH2DUVc+CWB/jhKZC+1TgGr06iVsxl8Zk1ci7Wjl9Wn1fyr
AOLchwhMy0pdHdNKbXHNc/L86IosjQVRNDhGo7yfDcd4g3ma6NyUaOdG6l7hHmdU
3DijOIqIOEL04BtCEYxmNX973oeHqrIutCJlCp3isURa2BzlQ0DIUipFi7kv5tRK
Fu34TUzqJXdfW/t43wm1J8IiF1p9XDDPkc37/i5e/Toqb91FvYVoi7xrLR9vw7x8
DurCxuHjlibHof9YCQqcxcGgY4FjpNky9v7/mWzTu1rFNaigx8aWK1wdPz73zRAL
gW0A/V/gvQtvYNnZvUdIV9c/UWDgqe5nutVcQBB1uLroSzfQqDSQiaQeObrGy9By
Wsa1l+lhIRYWOTZyja8ZLul3FNX+L69KddO1feny2I8Q9mHHvFwwM6iX6iRPt+9h
JZgt6uxhcaI38EO6SJfo5MzamGzGEq5EHT3t6vlyO2Jw7P1+WWug9yWZpHleqa1E
wBEqGrureAGlCfQJKN7KAjy8Dcd2a7/gXeEe3LtJH13fdP1x6HlPGnx5oc5sz2xD
gkefHuwzLELF1xXy4sJgUg6IypI/RR5h47/Kd8N9AeIB3eeHOnLrET+5BBaemN8f
aBGww1iNjxt3xpmC+K4BVX4AucWHk/sGaaKyfPxmoFwD+ovtcg/vFrbLknfHcS2h
ZmJitRbi+HyCsGOgyT/QUQ6BQjPs43VDuRisIfUW29lQMku67bZdqrcJ+zaSnUmU
mQQryx6gQSuh76w5CjG93Dpeo6WdUYFgMSyLTlxIr9F/cvvTp8T8mdXXB21Mk6HZ
+0MkimFL3Xr4qjDG5cY8O6iXoZWRUy0tB5rAJDnkL8Ig52vAjOnaDTuGv1ExyVCz
dkSRd2483hsJWkVs+bq/1Fy+GA+oSuS6gZ5Cv7ONw92gxT5U5snlJpWM851Aoh7x
Qada32wKH1OQyXmYI+TLtTD4KLym6Ca1ZDiIFkl2FeL5ObGqI0PHfSxnk4JurCoZ
kY06EofoEJsHWEIPxpyoXZWao48jSW00H12rkfMbgjaW/i3C/ZowEL7kNkANENJ3
//n067AqV7kzqEh8IshS+eaJGCqXWw9MyTM5dFXXai2MQjIJ6HA6WqBcDB1JOD9s
0xYk9WNgDdJgDImFUtee5/fN1m78wvuv3tJzjlZoCRPV0PJfPqj+3MHNYs1xTpCG
p0C8E0PEzKVnPRduWfR9Ter2xtragldknACX0eKYWMcV6s5z3laiNhL3YlBbqU71
6l3VxntOVhm+HGs46U3IYEG1lMLRHNrjZu1teMjsAejvzE+owLx0hhRk0s9U3o5B
hN1Wwy5644SgeCZHrSBo4okE1SqtbCsmogRU3KPtzLoB6T5x5I+QkZTHxOhqHiEx
5Uq6kSVwY10kefb3hNvQ+PAXXoMx+6PJvcpD7ot5kFbuwNKHAj+S0SdpMb7zOIbR
dbrw9FabVBFdrJw4O5WNEje9Hiyrw2IGyyQ4S8TVzlAalr7pfkRPDcjclHof4m94
+ERbz/sOIRRareFYVcYxMHnDStvQbdlh38viKlGfHHUP95mrb7f7drtpjCf3vuGr
hpfNTHe8trMMmnTTvoyedX4vVGP7qtlTi+gE5y4N4zh57m3VVmfbrNrK1tpkQD01
88nmyWSXFM0LNDfc4M++7UHnA6c/2G/Eh/pPPZ5HnsYF+jx5vpn9EmTLYajgwkeG
wkulyuVLTXkq1d2T64rENQJuImJCfYWrYUmSGi5E2pq2qwWtUOlFCKQXGPhfLT8z
GbbNNiC2on8OTeCWE25nMYcUaZPsDyUAGiVjSChP4o2xlh6oL72qLeG9XomuktE+
tiWMwh+aPr1+IgpM8Lujb+IQWfVF/Aj1HWsfdRQ3cH60N7lF/6dwsvsLt3UjBrpO
FICagSq6uaiS9RH3Dwks6xw3qJQ6CbKTlMMaZtVErgy+DgKBDC+JzSxq7+QXDsB3
XCTnGxfV6Z6zaDGRFYSEirk2uKLOHdsjmqncLFBdDIxL7bfwrmf1QQt9btYc6iM2
YsDVSdjd2l6Bz5T04ZEmxiD7ErBFKOBvD1iA43yVBvXFDt+a5rhnzIEOgm/e9CnR
vXQp///Rywh5nXjYGppKUwvba4q2ngUnOuzIdCQ9FhfF1VcV0ZlWcMjnMKVgbA57
8+eiBp/kWr+bjFOhzfpCCECKMjIkNZgSYBjkjVIjPRduJtb4P7lXAUhLMtQeRPqg
RMJysY/sDFAvw8CIR0GxVXT8a9dG11h4zKIgbxCpvpYVHaoUf7Ivr+lSVou6v1e9
PxdarIKyH5pJWtdyPjsAqvdbm6gJsphRNFVf5nh/BWdx95WgBEgJARTTjEZu3CeL
5B3rbM35yy5MXXPmvEA6oIBlcZZX5Cow2KRQEd79eiPnEY8wAiYQJGNXFDZH5oTW
ZzQq41F10sSXwTW5JaSZv2Oj98h1xE2eGvRmDcGRgupgZxRxA11gzTogGlfbgleE
HSCOg0Q1U+BJh6sJH0vyCj+5ydGLdXnr2QsE88zlCNu4xoIMpneNdOL/mS+mDMr4
CuSucGWgAjX3GNGSdUe2cz7DVWJE+cd894eZAffro2kVE9luNy6V0E4VkDlDdZNT
D//8Dun4LA3drq68vvGPw8nuRSHwan1NwL5Ly0AytCUW5E5Vghwi3Dhvt1OXeGkO
sQo65YxhrmSfGyV7qcR+5HFijGSoCBWqWw2FLvMayy6LnQNV1mFN8jRyzwGdFL2w
sHdLVwc1bK8UYYpsJBaLm7J1C0mrMPnAmQUvqiYS7wPDcB9MbCi4vPdMR41om1Pd
KfJl4DIQXMp72j4NvfRtdWOMLYPOVNbfwGRmBnxvpJ3F+vDUBZF+J0PR/y7iM6H9
P1Or5i+fXqPznjYoOTNWn4Vi2PDq2f2H0LHRWJKRg09vHbLvWmCPmxxrZAkIMTxD
XoJftPO9C/RwyA+ltrxadxGJSQLZZ18H7sLLrTERhii7hxwmN6A5jbgyVoru3FMC
Gg/xg28Ek+o5o/TOwIwlKSezIVq9anaRfUB083STWNSlqjLMapmM3ZU1QBm4qhk2
RmkqRJyOhHZM6hY+j160W4JIeTX3+8xf+FT1TuKo01PL1AnhBPst7BbzM85qBZ+z
W0KBHKLUUA7IlfCXnJzdVnbv0jUp8+CUKSadmKxJ3PGz9cmlMJ0idB90sWp5tPjT
nX27BD7GnQbTbqEHddbGUvQZXk6Ip1H1IqYIIkF5Xfeb7EnqxSOGbshAcFPbiMOh
81dVckwJ0qVLDbORWIpe1y8wGni/E/vtoyPgC0WS5GX0dJxsC4o5Pz1IWFZcnsyk
pxibr8++1Z1FJYZw/nOrnBejNyCcFpizlbukazfWk4oXoDH/qHyTI8I0+6DgD5kP
XIrgM2Kx+qUAb9ZIBRHlrlT7NGItHkpvmO0EGBI1afIaOWuvrADlR+q3JXCLucGh
v1+WAw0Jn5REvJGZC5LSCYEtL48Z/e2Tk/c72QfQZQATZpnH/1uQwjX5wsF+DAlE
I2QhHeivoe5VR2a2SB2HMzW1R17/vN3rzdXzcR9YOHFY5lFeT06MyWf1a363zz44
EN16VEEPRPhivsB6a0h4bSilWacQL/xLLCae6NoCFliNUh3zjQ1iVzLLSio0ZPP/
Wpk/Fiw9n7Yy7bnnxCWQf/a4gLN++tgQYxBmzVwZwND4cWA2zfU6wM5YOUagHznO
wc/jfdhfuy+h3zHEiOc3yI/Mj3IQ7gFspWRh/rqaDZQaPpuAKT1SwhMN4ULYEXgu
IcY8Hp05jbAErE6M3Ch7qVcAraBkYAto3AGzmlHbVKYkLjtM0s33jKU7goby7MOx
oBM18r2R1WObr4jgD3+N5sAMl9xAitGEVq4mCRetdokHwS1ZdJCHI5Zo86UIZ1ZM
gE9MXkgylzgK4EzvzXnAhZP2cpSbNX1ZQGuiFskxL1g6AfkIbIxPHHjvH6Y5zs0C
AIbIShVNR7J32OFSj2/czi2pTbUhzMZJm4cRIc97eKsHrf4eGEkotmxS7R7IqdXd
I8RqPDmkb4j3hL2p2OArFEplh+UBKWbxLuVjmB0LZ9wquoc/oQcXwJsqL6+mHiQ1
bTFSp/ML6AZdLkLZ2bPETRveRvC/Fm131uffBkFEbSmMi8ABnJWL3zM+PEic7V0f
jdtwIGqRn9SufNo1tIvmyKIjoRshSevg9TD5Pqv5tjybOIR2NS/HdxNvNfOwBplA
hKviPPl5NStuwxkL9WDroFWvqUybFT9pX3KvQ0d9paeA+ZwwVY4eB65SwXXpr89H
O3cfJJIBd4fzzIyYxSJr4Q/Is9RpYlbS6qYtK1pprFlcybILGWlmqcyhecxQL45d
IjFhkk8CPhdt9aDp6e4Vyqs85wWU2AjZphuGNHW60cW7TPrliAUI00fggrZsgRZY
/hubw3xMG0ynPPzsYIKLJOcUYhcLyWk/XrpnotjY6XhxhBzocXuxJ+Rs4Xc9blHI
mM5ymO+7eEkG96mZEyfpX8PnY8qkH1WEd1V+4zUPNncdu6+brw6RW3aJ1uXS6aEW
LFwcrbWHGXFpH3vRiyrP10Jo9Sh5Zw4jQ5Qqqk1SsR5RtZs/h570Y7gdvHrvYFIJ
bSaR8AGvP9WfTeMHvOOM+4LRtpu0e11xW6TwqWXxmh/rx0orbq+4U3uXwvWTqjVk
tVDoxpZGHS1uFecWtbn7owj0ZyH+F9LEpivhylNCuscj/qk2sDx2N4ZPtLGX0VGl
8vcc93cB3fjwTRQ/CQCeFrv25utyTdANOQIfOcegcsZwzK+9FZElzrJgQJLZDHWl
0fsAhhNXd8E4QeFRc/T4NH+t6uT5Ek81tpSXlOLzhwELZLVsFBgof+P66A7o6/c+
ZQZDJUuFSBnnVyCpc/myD0IgyGg4CUWQnXnAzTcYSvm3CE1FUEsBu9kan9BkSxJD
U7oShaJ/cU8fkjt4yxeXumN6reFd+2AhMr2OOffjCIBvAPmMam88qX0y0aGI910F
6GZMD78ld8yNYDQQEEismsZFmO1wTXdetK+w6pAnmVQFIW4gp5ds21CQgzheu6/n
13dTnCbw2Pq/g4I6IMkTEbR6sX8iX8wzEvAuMXAJPKO5w/W/Lsw7mN2Xjg1A1VkJ
VOOJkxDrRyHpEjOE3vqhikVgdMxPWoxXmrD9GFLGLBEsrleifBLg9/+5nXeupfRY
kf+BTGe66J95HEhjdPf6JB+PY5IwkYH7AMA9ALeas8CjQHu8j/zYw1vLAikjHiCW
1czy862EGp37sJh4edBNIaaIkR1kZ9ZUd8PTjbbnrT+cUJXrPRopfMd/VaKuHoa8
vXd/mim6SNUCoclyba6CMpNmtUim0/EDgWwfUPDGUE7vZVG8ADWXhHulXCjUuF7h
/tvwPDuv5FnTgSbwixDbBa4LyO659e5oHtoQOiPe93l7ukzKjDZPOcIpuquqAm7y
Nj7qElM/n7RseYXAlY36F9GxS+IuQfyq96TpZPoIkfedExgOmAMxZkZDBN9u6xLj
Reqkq3p3saeLHw2MzuzTgSiLlo0SHjftqAtfWa4FKmvCSfJ6KPDd/ON82DLTwZX8
KB6PfcZBj75eFDGUj8xaLf4y2h8Iqr2D01i1xOBAv7PelsldTlIZd9ADSLgoH2nj
RzePsmo5b7kops9t6UCdQTkM7537Aktn0b+cnBeKlxmGPhnWktBTCJOUHuwSUqcR
ar6F0R1M+r88C8WZ8/6OzLBz8PrSQl7/MsmSRFSAA6JKA8KQ3SdJJ/XvBsqxNIeP
vzNvaL9WvdtzswLER1mlncoO5gqhjipmvzFL/UVQyQ3ZbLvvI1eNcZILABs2qSTt
4puhkFJDkHYH3g5ZziAT+z8E0YBTa8RAMhq7q3/UABYcg1+Wmbq4W7Y++gbOyGan
2b/F6Zm813rqnEQtb4c4y84ciJQM/vHl3qRDrZm3Td0Aj0ETHZ/qLgOO/9+T5yOT
ZXk2EMBBj+azruTpT3QS7J9imUlurnmond3rcyQuxC9tSKUfxZS7kyT5Z68Msykk
l45PQwbiGsHJxI4GWvy3rogcOqZoo/cfqmM//BTGHR4pDgMwNRxsvGyX2F5R6jfl
VY52WqLsXPpDwdj/dnZZewELolaIp5tQ10bAVPOmCwJbA6r0lUmTvWGfVU3v86ag
39bf0vOEQ/XvxGZwZKHXzKbx/2J9aewK4/sdS/fuHc0J5vWjjWOSLZojToWKAlwl
QOEZTbSw6S/mLXxmIb3tVvmP6MYPdis4ztqBNbK3/y2HhhnyqJqBcndGItTAnoaj
SDR2ELyWKEXw1qRqOpfX4tNauuxHEX+rOuQCnJjfWJM+LvEv9wl/EU1bwG+lbiYl
cPMSro5dFPcUuRWH7DvCAED/vGPhMi0800PiRnI0NjoHtb4JwXI5rKWLDAHM2tuJ
QzvzHdW3aJKsRJrKgF+LprGTi3R30nhbJoTsR02slbBxTQ6Vn+HB1Zk4cac7tSiL
OOMSi8+pAQmIGjSOYlbolt2t4FP4Z/cmN3pDs6sHS2yO4lgf9OGz7NA4/j6xgYxC
F+MKTOs1hgzV/O+VItRfbljCAD+Vott3R47Q9Zdxb171lH/ymN9/cpD0U3eSI0O/
IKvg3rXLiYIBXrhC9WnyKOVkscIASc5n0cEtEAI3PLDSBE4hqhZRIB2IrhKSDnoy
NIeyk6oY4PA+ianNhleHYIN0rHoY0Hh5/0jwHpoRl6XCb5I4G/yP+4fZyo0IBzPn
vTztOZ8RNuCIoxH2+C07rmIbiP/2984ic0TZfuJvdV6haA+tp5sEmwGmu99KMQqX
Hhy+DppeB+x1rxk+9+k/FFhz/BkbGXWCoSUnv0PTnOtdDQWKYIa0AzFf898UgILB
Hj5aij1Zd+EdaeszRnJhOCX8MiHHIocpyd8h/ySYdllUokiG5XzNa/BBai/NAEc9
kbE4KQ4+HEBnZuURa585l3t+6gZwgJBKfPS9a6JahpWaOlpHCJsr4gSJahVDpsPx
ivqj1isEPBmqLZkcHwcNs/CJyzwYKI8EpdQcCJrndUUnGkrvMPprp0DkNZ4GjhUr
JjZCTcNcLM3zN+CUgw+RcCR/ZFrJUg4YcLpKHBvBS+qttnWsc975DbzWYGi5XnzB
pZJoE6OWXe6zZVdlEdjZBS79MSg3tRJYY+STPZW/kCryXyv2sumuz2zA/ogFQ3kZ
IB/vYillgjbkyhOw7Jd/l+I8KXnG5EHp0HenNJ7I7NEn5LB7FCiMI7QwM+tH/ocv
6x+B2/M93jm5H+Han+ZvEGS8MfeOrvH1t+eQywSVraopbzVLO39PZ316Eq/nQIBr
gSGTR18hh93XA59vG1R60fzLbiryjcOH3bAm6zv/qTUvvT9XTCG2zYQMAIz0Zl0b
IbLt3JlAHOH7UqtvxuuoHXyw0riWIOwTh84vEuudLgZ3eYXM/8W4DGSTRo4DsDCZ
s57GXmeEL71moh9hIa1chXej8lU+4xky96i1jcml7joC5PWp8WF/XiOzRjRlLWx8
DpNxi+H5p23staPE9Sc/3WFsjJ/tURwd1bRVABKTYWCm2+Kks4XCNstT0LpL69wa
RDh6JwEBFaolqo4zjn7BTOjLfgmlPhjioI1H9k55VDiPMpXNE+munjpAIyTXY18U
v0kZ+SiqiIZVSE0yz+W3Wm2c2V7QF4+Aq7FLXj4KCG6sgU7G0BHvzESRPqO8MVuc
fVtDN9hHAa+s6QD1iGGRtI68eVHgwx37xGnlVM0VsixFOGY5ghlhxPjpanL3ayD4
KA3h5EImQk0ocJ4cxpvv/AA5L+BJhQzA7OtrURdkWDSjt6VZ1ildffkW6QX+8ce4
tYjC0722c1N0LvkETVRXqaVBT6QgjYfCi+95V9K6/SaCqG7aMEumJZDnzQC08pfS
ZIaONsgjIBP7unrme2gt/T1OevQmTdin2sHA5qRfp7h9EAaoZ6uKlJpcsGdYaNcx
ESoDfhjw5JmOc2SsC84OBT5uUrNOUjHTk/6tz3ueYCDyganUmo477VH7psHV4jbB
JaVn5x5bDXq+iyhAVTz8Sy3r1VvQbZW4zl2EQsY2c5FQ7ukInqI+ePC7PPVmd3/o
NOJaxifjIogQjS/FGrIVm1i4nspucIScMQ3ka+rJ10O7OpsZItRr9KRC3TDOCiiP
nG7AlQX5PmzyBDaAsATBS/QWvGfTFIkzrRIP3nSI7F/sEeYfoGmNNwZtPnx0N39u
8phYcV2GDU+mRj9sw+km+RSse+9fe2uYYqr7PnPdAfQDngu2qy84dF5bHJazv7C9
1hAKXenfu7VpTu2dqYefgXLcoKrvIdWUT7lZrsR51W3F9JccTp8jtqCwkJyavaay
hYNwDTejsXq+tPor1XhEfHhBMWdP0m8o1PJKwwa48pN9X1WlsSsFKy/H3DQk8qQc
2n/HJ/Ddrr8+LJW1/ahXdPlPReadyhwojxIoWWsdhtc3QoILneWzzAt1/0s2Jasf
UucGjjReBGu+SdBIeEmrpOXyaEOggGtbZpl+lGeaNLxdKDOvasahx3tJg6p/cqBr
5zzi8cg8L0xVdgXS2LDbUdlNU460VCpIAoVJwRbVR8tOhr2aWfrcmzQM6VctAyQO
e+wzfz7XIt2pmAVQXry7A1p+Fp+94rLfmQtSXgpvLaE0Xxatq4gMkq71TWvthPRk
Nkf7MpY8fupfSWYdx3IqOzTD7FmVkS+xxBq3KpIPi1zBwXIep4lAB6r+RhFqr5jo
UbGdAhFdLh65ovGALnCXuSrdzYZRSIGYlg6XDUcD0csHA+m20peum29VqRKWmeh5
4EMcu2dR/DoDqyq+DOPUjiW8vqs409QGOirIOYpiDyPJR3G4+Uruy8thcqkdpf2A
nshorXj7fRr0+vxjaJqkCxd0/6p+lgMJi/NICEwPUFvY5eIJfvd5JmPMgQG36V2V
oRJRF9SS0j4EozSg39dqhFyQHj2byW/E9DiejmEGCNdtSUh5H2+D2wiMzN57nWOV
6+TJvNPDMzPIhrs+zwEzUPsaLP7J58/HguAk5kUr46gAIZhr5BMEZpfniZSsROuQ
/03Jao3bVXi6LohCwFpFp0YG09pO6komu/h/kKQZPfNUJbd7rMaA0AKKadkGjW3v
RezQ0X7TpBGB2clsYRT6ZLNNBLlx5AUp470+bCLhUwvTQSpM+0EvyBUWQ5JgCCED
utfLWCFgMq2N5zefX7EHd9OYsRjEjm4G8N2PF+YhOAYE3quXVFBzXMHhwMwz/zI4
fdHrGwGDNjizkImEigdUnX/4NO48p9cQx9oDEWs6iEUFxcSv7AeSGGU2xWzX18eE
38mkd5LvtI5OinAbqIlglh9N9JZUfH1a1whWeMpJWJG6dO81zneCUVTizgDNVZrN
V/QSYK6WaqcRWX7Fl+X74MmRkiJCP08CU87KAnA8VcQknE558wlqxBF2ybvdvDUY
AP0Gnqr1oSC1kZvsQSfUVNctJE+ZevgZdbdL04IGNquqyKah2bof7MXbnLq0+wUf
OZRD28guCZVTODqBUcRafzZlThrsnME16xTvKMo5Ps/8R1MSCHBtiup2yYra5tpL
RKopyHajR3dMLuKyZ4Lp6JMqcAs4GJn8MMvlIpNQsQznZuQBdFjZXrDYGU0vRbub
LIe05qCdbY1xQW6j7hqYBTx5owFmNQxocQXmecamwI3bw2CB7LNPti22Xp6+wXHA
OnyKqcFxvzeO46I5A3zWeY1yr5W1ocybBM0GqbwZkHbB0NVZjNzk5NV6NzIm90iE
I7vwGChmMZN5Z8IebyFiQu4dLfVEru5Un1CJA8nrymZXsAZsgzFLv1FAJx48N6xy
aegF0uL+I7v2SwisiYyQjO3cnViOz8XpF1/rXDynaq1wnYNduKM+iJmlddMa58d4
l2Ctj/PpedDsjd6WxUsrk0UyR5Llfvjsb3Bk+uPXR5qsx6OsIXjObJjWKlBhwLRI
qQCHy+qaQsb48Cmyokh5SYW0GcNRVYg+hfDnPmdZOPknT1en+k33vpMp0r52MKoW
b30j6hj3EWlSqawGsHYJ2151ga+acLtzVG7BXuUBd/ghU0tbFHL0KPaHx7EPOfY5
OHgWJdSwErdXynY6yUhaUQJG57CAdnQs8LN/zMHugF/Ee2pIbwAzC7dTdChWom/F
Ss7Os2WLDPQOTXi/q3yg6TR6nwtjBj4jbkrI6aYWQihqiP3t0ntx6ezth3HDgh7/
0oYTd+FFG4PTyHv6FmWP0M2VdPUBIhp/PzDaMi7c2+/q6+/x695bn2i3lBG8sdAW
TiqpYEkoC79IfB1MRZ1Lw4ysxUBXmZLrx/kvXa+jxOgy+Md1Kykc15A2VBDZL7xI
ATNdHJRHICE7GRIdR1eZcvkm/vJXDrj+qOYlGFaNZcd0P/yXApeI4fUoKmooHL6s
043ZqM4fSasVJxCg/0Yn1klamp5Q5nbUnnkgTPOzmAxzHpNnJxZTxJaplxSQQwuM
3bQesUUYpzhA/WrxgPYMSp+eipUy9wYcF0MZGrR/89zab0Dv/7eq9BISBy0Lp2zi
pWVng0arIfxk4pmwz97/hMHD8YTvefIaIPGdUIRpP2MKyyx615e+SJIi5O/JC70q
PlOo1dl3SaalYhbZfJM8ht8Iwz1W7rnQkvQuINlOdzmzjZ4zRx21FHSJxli3He75
MYH9tSKM1vmtWENlBZNsRI2h1mod+dy6+2Hkb0fB2RHL8Jc/vjR2O6d0ljQto5AE
h5wDO2BRBF/xApk8Hk3woZaOlZlIJ97CZzYz0QtoaW2Jj1KmyxDLvUqp3M2/fOxW
8T7c3HhFzqyAmpq555Cw8EcaEkbCYh9r/I9GsGU9W7xa3hP/HzDjdSsITKpoIpo5
+LGzvwMQmTwgzeo0YUW964pQhzZsxl78BprdfD7siKDQ/Ba7NZevE2AYPZL2oz+j
kRTq2Fe5wePrRW4h/a5u2cwQ/nCrlCRQ4c7iWM42lFf1otDbkvT2/rmXfm4vXB+/
8vUpU8OUgm14J5iZuGk760fv9eEjQsJssxGfy4D9p/pTfsQbzdXB/He+FbebkH9Q
SzY3xVow8Aijsy3vAOBMpyVZveypX0m0j/keiMm+5qwRRuiQt3Thi44LPklZZnyC
mgurNInATSDJOQ5tlEAhWkLskBEZbaSUPEthICEFtZdJ+r3DDPU/CN9/MksK56aM
0uvDs+qDQw6Dw86zOr1Pt0PF4XOKrXz+tpyycLXdAD65xoK9KVunZJNOjBN8q/HQ
00VazXO9RXNFSeaYtr71n2IAXT7JlaFRRG2GI3niPSOg84V2yDX0Kv7p8fG0nwqP
r+eZhXXRf7N4mgZP8gL7D+3egE5fxVIGLprF9RrltoUuyUoqBOUwk3tzKsJsZiuu
RtsAGbiI3vwUODcqm7HUOBUaFVir279PszTCEdoPjRCN3gCrZ7sYraptPBnjYUdN
ELGEU8It4aIMZqTJd6Wc/1z6ekJ9wESUxu9yoXstuWwg/2GMXWSwBet7jJYAFm40
Rdq9G9Z7+2BxQpcHiXVoiaqJPLkZkk0cvI9J+lvH+ZOhqy9UZ4RpoAz7xMAa8A5D
CZgBAJiyXiHkRulwr/9knudTjkGcRhmlMxp60rDVx4QN2GoEe/nMyE/HSaIcNWia
0S930k+w2BBO36PWh4vJczFupMW1wHLORUGLNDYhassvQ8yq36aUbwKywRmQLXML
iz3s6K40Tu5WmrvcR8hM/xs2t+8NJ0mXQuzM363faP/iiTPaiuG3w91NaqFjOoqk
XzXT1Se+eXaVFvgKEQgWHFuC+k1SXI3Lgj3hT2sLp+pGTNp+4XxCD6aBY0v3jHH8
iA+kgqZN9aFTJVS0gbyVzNnb40xMSwssSOu9yKENXQZD8O7TQqa4gXQoyrKVWmRJ
h9/eWNttMqcUNHu5umIlX/i2XWdlpMVeLXo1HW4GN8L46lOpUi+m4/PaxVy8fMH4
+M+nJ2O2ZSUQZ7ziZ4bsRKrzv14zsz/i56z6RX4OseKDitzX9t6MEz4IxgbTdwXE
V1OR5mGyy67aDhKS/2PCgYTnCGQHAOa+9CxfLG7HjlJsLj48CL/d3OAsq2m0leTH
jsmVrg6Ewah5lOjgX3pWYuYSBkIGboGGpkm+hQWXNLHYE2dmX5Ylj94HJ+Y31WDa
irXjFHO89T++05Rlf0L9dYVE57eAtDEq58t/kuV2nvZw/XeWXYi+H/pcg7S7lr4t
7XlNWwZE2uYETcv6/pUwbgi8IO7ntubR/ClNKPtSpPBMYGVurvONINqZRK+/iKpI
wyqRuu/lU27WnHV9mKC02Ea5zMVklIVgOrNQ+mDVr5T7QY8HHDeP2efhOBWjxsOU
ob0FqLfgA18YrlYdGr5Skd+JlBjoBu+0WXZjBlf7qEnYaHnHkfvK6mpkwKZz+iYY
TjM7ZWsmlVnFI/LH4TK24M0DA6XP5VkOKkBMGYchJcuzB09Gqf/IHBugTemZUg80
uk2hCR3Pw++Sv2mv30F/EYLi1BYawpkAN7px3q85TjKj2wGkrgcuXOF7q9oPjG1K
A4j/TVak3b0cL6vDVdT4WQ1r5zVtA1m4jpBza0c9p/NRUTvaryioKEbrtgG2Ayv4
3Xz6giSkDd6H7C5s4A8/c1AukR9pvSu9d2DV3tWZ1lwuFbcjYH2OJHyrUSAnD0zG
UyMPwJUXetTfggp00g3UmDfRCk+ri4FBHV/oamOLUyks013I/h/6YO39eE/ZoX7o
TTLOAn3ceOfW4BJ0Smm9bLTJv8uLREwI3kOvegAi18BLk8ZTuxtxbXkbBOUJp8g9
BHnkyAP2A8WIDMer7+lDO7cT4xlsHS+F8OWG7NMC0RYHeIxuQJ2bhFJBpuPCfSJM
c7Pdp4RFxu81HBH1L+XM2E/EqBsU2CwAH2+oJavfLfUAqA6ET516mk2eXfoZNIBW
Qc06BqqNDiy/dvR8iTb0zs0BNpbJ3uWEP4IkZWNHhDrGW6/k71R3wZGM6Q+cgAys
TLxIg8cVGH6B2OibXRf9VlTEXYQYL3QfIM9dEKv/ZRLpHMHSvTI4w+XX/nyJlK8O
4apeV47UEDUQd04ojC4eLaxGrCPX77z+5G6j6uvtQewPHyzgBYBAJHkPUcx9P06E
xzNYH1CSy6azNaBTspZ77VhZ4bEKeidUHYJIOTuaXzjkeMjZN/H7vT37Bz5srfqB
dVakD67zJEjvkjVJJoNmNFgDMGhQlDf/zpt6tiQj4h9ZI3a1Z0W+mJ3UWPgP3GNl
vg5S8aqMccs0c9tmhk8ycD+3a+/fS/FirnoSKQedgNI/VpQhhqHU/1imqRlgQhDw
x4g28en+s0hpilSioNi9jmu21z4Fnqg2kXaCjM5alR3ZMGMweachaRNQ7IupcF2K
taKwSh+QW2m45TpmFKw9ou2Q9m8LmRGx1AqufpUGmaaGKY7VzCB1IbNDb3SGpXcG
gw1iu3iiRz0ruVgX4OOCJFiQU1f+YKi3kN69YBDsZ2P4jMv7sizjM42pf05oCd9p
E5IKj46sCFTnBZP9/yjudyqqB8pVajptaGBZghChpuyrrw+AQ6EAzaJAmV4+cYa9
P4eFDgyz6TVjhA976NO5Y89FUSUuFdy6+hr5OiRPRl/nBgqhg5pIOXEYYCcAJC1u
w2X6vgumUQUyRwjkTtJwynGPdIHMDA08al3bJumw2qojYoVf3eD32Cn81Hz70VHY
kD0pxc+DXKYQkrWV5lslWK6vwt89duaq9zfTMOzilzhkXl8E2mqkOvpKdjrqaw+8
8I9PlWAtpHeupOx4KbHXJx7S6PCzli/fzPLTbzfJCbzSD2umlD5m2epVzwp6Sk8V
svGsdKOOxkWKWZascrXXaKijTUZmobeDOKgVX3DNrSX9KyXbO2cV9RWkLVoJ1DEG
nWNvlkwyALSho3HfxdmGMwhb36mBfEKACaFk/MKGDZ8xGY0u4wqLniFhqpFb7k+y
mrPrhbUB8iX3J0w3YIRMfzd793PIam/iDIgVQUt92IVveJxg/VqN+WRnLV+kZb+R
//33sYa3VpVgwW5KfVK/rVABlbDbka2zqfLaJaE42y2ET6f+x90snPCa8kE9rhLQ
v49myx1JLkG4vvMQZ5RGHscmSFebtMoCOa3biQHayL/WNe/4K+GLdH4heMnrSK3T
RqpHswvsuY4XBjEUpwizJDxJ9OAehee0aWwzO2n9g3fYtr7uj6pgfp2B1XTkBo0K
hSCP6zsOCeq9dQh8MC2wXjfz10Mfo3PwJojM/QoICBY4UdfC85r6mvnDiozpG+qC
S6jZ0Fc5UrEhexcpdN5zjnIjkat5Fog8xVZR7aPm00O5DxrxO7MCqmNdtbdJ25+R
CuFdYitGWYcoS5tHfToiiBKpGcEWPFXbUm4bHigf9j9W6ZUB31HtZfB7wObLH4YO
MeWGC9JE/Mz9hco5NbHZzPLNdpBLh12rxnANf2rcxr3KEFIWW18/+mSKycutNA5a
VV/SL1sAlqmwoHgzCLC3OdmzV5Eu2hnrCLq3vIVe1UfW3sSCuJ0keiDoI609evZE
aiD7HMi+dh2QKSEZnF3qwxQzIIeXWwi981YGpRg6qjie8Hzdvg7VO8QLdVxRAHpg
SHs91uhUcYlaWXIXexKAFJ2ORNPY8nJ4zGpzeImC5nJF6MwSwlqf1uEOXGQ+4Gjp
TSKV1IE19OpVqF3t8ZtwFR0YHzCSDLqORx8EGk96+2y4Jj2mp3FVV2lulz7jSbCG
uu24i+QyToqLZ9Kenp4Nix8957IE9V1n1ujgh4Kip2aMXhL9/wQRf8WrJf92OwdO
NGpiLp9P2LYqprjmZhq4U4xYGVfr/PSatjoPWePCgdWJuBlSLX3S4bHaQvn4yv9/
ziMjP14Z3II0CWfxCVu1kHWxZ5YnuFGLBonmucp4sX/uBjjUsB7BVxtMeqfx9PrP
5HOfoWPDyBgX9mtym9d8iygLpIgweutD0n9+6SwNGQgPC3xEzBQU9M7+2hTIWaYY
mihdtG0H56MNej844XFuCXgxYG07ACvjDLMCZssFnmfGhG44KG8znGr3xx/NrRMD
FKQSeeGRSugcEgQCK8aJsQrS2S1aZ4dgP2ujZ3MYpAQJg+2kRSzRp7ky0vYd2smA
XVA0vYGKeBK/O9Nrg2mzkUep24NIMrPo2UaIBQ01bNQaw/8rEuDmTVRNncYqBH3H
eYMwNmRmIGB4VJU0WqqpCZfSxPCVLwSvTpBQF5VWkm5IUSUTZS08tH5GG2oSAerU
C9dQfFzZaNBd4pDN6yXz7slzjR6SW2xZsPyhgtN4SV1HSE5Uer+PuKb9Xz6vceBf
PXJlj0QAQVgn3D+T1EeEkdjqJJXqdYQKOS/W5GTl40Uxx2io7dH1iWFeaU6Egfq/
qY08/902ZgDvyQwTVbOcTb/OObrKJE710uPPjIRHm3I6BhOtecAb0eMOyVU3e9Z6
IDPfm1XMLggbkyMR3ufQ4to+qf31QYePZdWWF1pQIuCMe5IeBUlmvoBSd74A1fOW
pwob0nYixnopJ6Nt+fEjDQKshghmPT+Ml0hIvxtzidS2dBbThSticZTUBWhNpP3b
uVmEQACekjHXT5/RO2lj8Jy+8SmfXdxJpp6S3e0ADBg5zj9Al5VfFAbTnZQ1pV4Q
beqEeUTh2Yx/3IJaSulgldYNHbJaymUJHpQdgwuBYOtgcq7X30Git/XMDS/0BD9d
gdeAteHsUV1kxKQdHtFXaSGODO/Igg1EOs8DNrHBCw3uVrpavuBkDl2p48f4BcGz
Q65FL/+XESMYbW86EIYCR00PPC2U903OqQ8BByZM2MOWz10VLB2sEYJ9MjqC4lie
3pO/fpSrHs8Cn/Y6CQpT80HuoR+0gKM91FOrfJI+JZP4oEflE1m3Y0jg2MGdKkNw
MB1BPFEHEqzA+EP0FJ8KPmIS93op79th1rDGZ4SUo1crewakqnDrQjZ2SgZvhBVA
EZz9SNfNE1iIpiUrowjX0jJDy0pdfNUoVJ0491fTO0M0K1Sffa08xdpiIXNB8kyN
oAx+6rwJaGoB128tHgOgjzJQL3/yT3YjeFmqZdFSRhlCfQJAaZTt6hrvhweZDuZF
66+lWvqAF+tRxQgmJ+0zyLIoi5mHEGSe0+gv4huJ2b+eM2M/o4pZHTA+DRK3Sn8s
WWsIv/m+w2PCcI3ErsvhCgQIaQto+E20W0oZNtXdVIPA8m0vIMoagZ7azD0ahUQj
EogV48ZpHM+cxJX3j547GmJHY4BBw2iUnO343PzC/StECEKB7Cn7Tgor9IT89SD+
DC9MF/D4sYnOqfu6dUOac+tnnQPZmvI+Txsz5quhjglU5cPPLNAuUr2RbefrW7JN
e6csqVYZU7s5egY49k8YVqSCQN8/2T7XBbXweBT7Dm0tCFqDBzgSetXTAtsHj8Wk
skBBkkiSjnhDFBc9HdtvA0TjltAMaHhyUPT1qCgZ0I57LO8Nm0BWVdvdm49Vug60
b7hpTU8uSXGoRZMwWPXUQnjrDJPwZE8nx4CH92SzordEio59/YIc4EPlU3cH1ADX
vsYxdOFhNThwc/SPgzHqiUq+MJ/H62lqR29WqZzgxdam2POtnJ/lQblMgCJX/vTl
zZXwVYBtQLMsj13sMmLW1JPu0IfD7ngImpV6vg1P8wvoN25sjcyCyIOJq5ItZUcD
ExbcMknnOuBxN2bOLk5UbC7iHDQFcOVLilGQv5CTKRiIfV6Tin5SE05LnM3s6/CC
HQLNDYkDNPpZi54pCMpRXXfQwkc98RUfAXm6ZypQ7OYdlMGgD91gT5ItaYI0iC+L
Yy8sH1UMUt3RHWuzpm4PWMvNgvfIA/+ls4Bo5cCXghHRxL/3gl/JP3f3ZkVZQRxw
9fxIyDFZ8zvWNaLBpyjfW1DDNfjNHRPrN7cCwqNjFU0G2SqnFoyZjfTrng9ch64F
DIDTk4IPblR6YltmKIE+yJk0zBERDq9Z5b3tQCiVO7Q0ZVTi1J+S8FenX2V5HLik
nQTvw0J3Zb4G7hpp+JokDyxVVgtc0SpZEiUUouE7qDyAiW0Knh4590d0MlhxFkQj
KLDwY5tEfdDnPnjekUceO5or9IfWpyVDqot+OtRd1PgloVp6brJQobDiDTXF434E
2zCcdx4W40nMSHpL81DpaKcGfF4B4RW+ZOLEZeOksQWspkuvqm2VxU87K85oJGWZ
1Bt8/IXQkddnZkAvWBWBT5PvLMtKMcERSJieqeQGT4Qlfd5ovCi/Rwgc06e3+VuI
b69q3DP3KrtDkfJmRMKunx6oB9Swui69OxOFYvfXlYfc7bTY/TtbqgyypxWEy1ID
OLS9Ub8rAwdQkoPLiUm6xFcQp5BZPBg04WMXixkhge7a1BMRPF3Ic8dLNpXOQd98
U6BBqxwcAMOMGLI0BfRIHLuzGbdIVaq0NgOZ0j5hQ5qoWUS0kBH/PwcA4I4tP74c
1MZdrWjaB+sIM8j0v1jqkeTszXM//hdTDC6B5PRfu5qZtYMjj+gy8Z2JjRWLF/Mz
ksktogmHqL3cij7LhyMrsFBgoVLawFHaeO4Gs/e6w2HkH8Efl1USMfl30y7ITNx2
mKlIVOuVKfwhNPW0XnQReBQqiibmuBMiGrLChD4mByH6nQPxPupZZtLhl1XF+aSp
SoxYkGR/Ta8/vO2i4VlyXFRTCBnm1C+oz497xy0rAbMA8Ikbt9FTuT/JtCmuU/WZ
9aDME2r6u3LaSpZkeBpVNoxV29kEh8JNjcXXNq/W/V06azhm/Tgm+v6OoqmSQQNY
wnLfZfWOBQE1wzoMtH+AslA6sfsX9AjWpkRiwJuUH3mUX/0YvqM1Xh6P7LUznXII
NZNM5RXT35o8wsjApDSfwI9H7PO6OrNxV4B19vuzLQBLMEab9JPAeVcJXoYapoRL
+YxuU1jT4AIbX/BKntJRAPe5q2NyWZdCX+rRzm3ffpjScGUZEX9SBaYIvwR7b51s
4Xw8t/qUNejuWmrKnyGbo7ax1AlA3mwD1K8EejC5jXUoh6Cz9I7+ttrZvOL7VqT0
SSKe1Y29MPvAiED/QaYhTQR/58H8SR54ByM8Azm/7G0vP15LiUGbHoBa+fQzOE/5
IrK8IGhwn1q9yOW2pGW+a5sVkDEIOFv/2g8yJoTxdeeGb8daSycJoEDLYD7MqUoC
BB9NoZ9kb8El+Th1RJyVLyhUjV+b9hbgWmVbA7i7vMxUBxxkmUWIkWLoQ0A43mWR
XinhS3zexbO4dzMRZTKkSTaQCBcPZCT5IbOxDV8raeyDtpQo5tCQ0C8jUQ6nBwCI
WJnQzsvDAvFfTfNkMW2fu1lKRJBuXSs0vV2xfRAuSP0Mv72Xjjvjt1SZjaK6UmPE
9XNdAZw2KT4vPmHPw3IdrcMPGvvHs6Vv7vMPieelTZw26JVQTfdw0pnlLg23vxY5
KqeSwgus+P++4rnmo8ZrYw/30AP8x25k0zYRifCxZe68um9+h8FMpPFovclBxiSr
v0nQiFkopTdEYc8D2nWqGGITIRRcA8qAU0YbGyXVR4J3AXwSS8nr99pvqn5DfX3u
+k/LYDde5mrB6H5+AzMDP3JLun5dTxpx3eqfCvrFiFOByP8FhfcjbhBiHZ79Hr06
caq8tIa6UiqbS5o0gNfYo1V7H9LjRdwGD8zwpISKY7ZJcl5U4ro3TXyEcmcB4+E3
gJvnRbD84HwnXCRt0cZfTHm++GUb2MdgtpwHdcbhYR/IVGcelfCSf0rdVP0Z1DgT
hqfJcqqfH6fOorgWVV5zEjUaANPKTHi2+HJH0bECubEtsi+UFCPnb8m61ENwW+sC
bbrHwgYqVHHXOmYy+pXa+aT7YDE6ye/b3SWRWw7igSfWtZT+KcgJbc+xkXpJn8QU
zlFWEWwC23hTy5/g8btT/BfSZ+/BjCLCOPmF/8dxnP2KbrFQwFdlMWhwKqJ33xKS
wL5ynj9HRqbLlR7VKqFia6Oozsc6Yz2bMcfjsN4/oAq6oeIIFD3PwHr5kH3pJ/N0
5DyIZfU3lYwn+v38ff6K+JS447YEyVg2cXEMzZKIAJkDmrUhV0HNPxnz71gAKWsM
Wx+iJ2lI48u78dHwbibHvAXfzaDZBtN7m1JVt0obYlzDB2gCLE3bXBLzJhj0c/uY
K3TGk3COwshBD8lIkEowz10YzKqeqCX9nuSmbZciR1rO4pFuWoEa6TlQqs7Mk4LS
tN6CDgfRFz+JnE4tryh/87Zlj+wgq7JG/9NtAu5sUS+IYL2+kGoPlEnCDm1jj1A9
WT8gQzAT6C+NoVfcsYYKEh8G+Y/dmZgNSY/rF+ET/Zzd79rGkVmJkVTtHbadWcKv
uBYA3tRKDfq39/e1vyBA70EjSAldEqAjwSyrJtyP2pTC9vvCiPCHVt163wJaBjN+
+LhtgPUXVJl95wbAOG7/dtbEUlJFR7fo5XbpNp79USYJ6XeKZoLpnEKpOWhHXF5v
2M6eJadYU9+ep78/v9Z+m1oZcF4emkL1rm8H3Tfun7kJ/6eUkKaHwZp1gL3VGIqJ
FW6uunniT6/LEPhSlxDGP0cSZCx4KC8l42qfM/AInFwpCh7uBRVuJqfrdr6FLuGy
83ALBPsrfs4s4i8ZWf+OalCBXDlFfjz6+uysFmz23pPcrcMEp1KJOZXpXJZWDHhs
SUskG15E7icmtJx3EVPaYKg0SlAiQ0V5CQ5ZF9bKJuvoIxr85PzNrvtQTnz65+71
SjEb6qxDuWb+Q/Z43jRfpPHacDLAO88bmMqqCA1thHPVczQYS1xcL2SbLqlIa2ip
b74t/KeaDV0ebjJRKPm+rDAHrxaqMWmYjCLgA7nVffF5ZBmzN3/MqetBiXeRJzZc
dWzBFH1ktqXfuBOc5iLNAlsq5E7xlKfKXWrp573DWDDPWvIHLkLgZUoVXBFBheAI
Jq6ulwTU6raKq8yy2q7AfaP4vKC0v0DgOomxLwz/DzBN6kYYRKMoICeiYraAVxXY
UHImEdl9lVFBCEdUwuoOTUmL7I4+f0c8LKEpGf/dYpdIN9GAVpWOqNtRP5ACXz4H
MXXwJ0oI95e+oXa/iBxhd80bEMYWEBWZhK5Bam8BPgHytEJUCmBaFlm8VhT76yoo
UaDVtSeO9SM4AapCqSADBI0bsZ1rRV4L3CTr6mgPQ/oAS4Cz0C6RjCsIpoSku7v4
4m/2wC0ADfLrXrvaxnK9WnImCSX0r72I++3MbVV50i1w+xSseAFXHOB2LRIqRoQ5
q/JNh7j0taN2wI77qGVJjU6ecEyT8Nao0dKF2QDsT+kKjGjyr4IkjSXY2O+9jWeC
pawQPCzgyGbCuKb6+X7Jc95eZNBWvygGe5W4/csJanwcbL3dEGuPx1dUyPg7X9aC
DxQNTJXkVOF/CrL9i6tCOepKuOWU7a/qhGLl6XrOQTE3G+u4MuJBC/lm6RQtIUGW
fMFtP2CW87YPVJljMqbNj/sm9qjCrsi/oB0Sk0VNt9Agy+QHXtYB3C1Unc3v0JT9
wl6SjECCtvqwpQLMCQgiHHH1imMI5sYDqz93/pW1Mn4MkldSNswt6KdzQ4HoC7Jl
nuhSKTika71AnlRWfk97bW/lJblASmtZdbcmTeO6sTz2+ZrV+urH7DJboqLM7gKk
rC3RJmDTEDJjwzwARgD0ND8M0kjlMc7Ek2NKy7F07y6mqh24SCXZk4WFxqOqaPdj
1bHGbet3IYCC0Z3/B+hnDkMCMT8ljUwU3kME0syrtECGnfzPS0Rrmii9DZ7Mi5au
1i+i4hK6U5grnWTgt2Wi4jeOCr1KmZgpPtcbbAjrV/0v8UuGD9GrlI9q2O9tW+E/
VZmLZdqBIulsrw7T8FSyfGWSNjxQy50jVtI+9dEeBdLuOYpMWxhOtH0k2//cMIBH
PCAZIU0gNv5CR8cOrhOKoQgaX68w1LCZFcy8hwaCce0ibKzgs3na5FgXMGXoQnLT
ska5jPXxkDj/+vtcgCu83m2lC9kyluzw8Pqo37RFWWagdKBRH3KrdFRnObZsgcvy
w3BVcGb7sJ7rNkGMQiScNy3qLG3mH5GcSK4fSzb0pOBvezekuJj5C/0xqnxvNBHF
IbQ/K7kINFZifxF4n3WLl1Lg6+ecJNZd10ddjqbyx64dccJ2KRUPsRdw1tFUMOpn
hfiZZKKQa+OSRMbEFE8kTTtssIVOBHTmyWgvFusCcieIYKZN1waVWqIQ7rH3Z2MM
CadauBqGapgGGggJY7jQSZ6QQOP6PLoBo6zp5ZUR+l5hGglAXf6sbtKb9gka7lXG
PxNQ71oRnVej7iPvXZ1kbbshpGi0uPdhGfnO8z7vg7oyoLK6Uu4W3jw1X0sSUjf1
BLVDhmZZt1x7OnzFuEzVqq+wd+OXDQAvH+EoRb79i4jlEaFo0GnLIl4aYJZQGSXq
gmm9XMxoKZwBRHP06Mc5OWhBT9B5F10kijZE5vlYj+nMsq5gQjbBiYbJ1fedmJSi
TrO/99hNDkctLnCqUPVn65hkKeSFcuQQ2oLhUm+Y0H4TlTiBm6jqAYVTE3Nv/8/D
FDalBHHF/m6ZX2q2pjAN7GKzmygQQ7KzZY8EMtRVhpXfRQrnt+eQaMrPtfJoZYNa
6vkchHj14FuWNK0rAbB8s6WbcubWQ2wqAev5/uIbBy80WoKxSqiu0x5sv7PPhusV
Rkv/E73M1hpNUjnabUr3Qx8MzCaCfdiu6zwxQ6vXkWTJDAzhScUWCKkMZTSv/lPP
ATBGHsXBhD9idae48nVNjxYTtlKWyeXO2TdD3USldLElKmtpVerQVPhU7Z46gEvj
g0Qam3S9ct9gu/6AxpIg4twChh0S7XK4bBhmy+qOeltylLDTzbs38zISrlMBhMth
17Zrk1jZ8h3a8T54PYD69nIO74MhFc+PI7G2gPZe9oyH+j/Ztiu2iG2SkPJ3/DZt
2cE6Dq6V1e4bZ+JUZN50YphdRnmey3nGBhUMuUyonEgtYO5Fj7lFCIb3ohw8Z9zp
aDxygIgN/6OGYJGoZafKNoDvDRllLvcywox8/FKDEyvpwzv0EvDpYVt35M+qE2FB
nP0iJQw+sVaXMQezPRO0Wice5tFa7ZAgo/1c9HFGkmulKuxCWorqH3RRjot3l57V
g4m3J0o9z917+tev2Sbbxt8jzxQM2ZLJs8JjRlMQ6ciDRT/ZypRqiJ72pb/vetCH
vCZmHzu4C+GOLdPmp5N1IKeutUW0aRu9FgrjuRmfBUWYTRrbG6k5wibNZYfAf8T3
OBVVN+dHbjlMDa/0eTMOLsTTCUFxkzAMSDfHVSjDBreS/SIEQSy8kg6ulRU8Od3m
9TUCapyKOJ8hfFNXXAXXh8WoELgZj+hSMcbGolyg3W+lBi8mUyKsqRNUvkixtX36
e97Fuisll0owAFLl2ZBbiK5oaJTk47g+L0vg9+fgotPjq8itnlxKJTsZdDuZ+Qnb
CbMA7eVfdAJv7pATGttRldAGmCejMm2tCMncIzi939J6GWChpgvL03ZhZLyoDvfp
tW0wzZveumKOL4kJHHE5JGjGaqTmw17hY1cMZNANcVI0IPcJjlzqGnicNg3yjatZ
72uf0VEuxoRR00Lopur8j3f8YTz2uZdFvA8WoBsfTQfqQW5QFbK5hnAxmCwgnd9i
lwt+pxVHXpPHCo+mMAgwEQmfs6VcC79KEBxMzekZtpjR2NcrFyWlv0xnhhWaOe0l
bsKN2rld7/sJ/wn1aUF7xck34C4aXhjH7rk1q7Oj8cxfiCpJsWnQGTjJf51kvNsG
0ZC+QpM7x22u9SMpaEQna4CfvX4P9upfgmFauFiPqH46i/AXt9F0EVfMX+diJm1E
ymJGwWHIYWjV++/tQgh5QCE2hhe8n1jXzvKipqOO5buqDcaCXpal2nKJ8MWjNKtK
toAaDd1zaToK6PW380+zaO4savgLEgZdeI3ol78YOEhMpfnLgaf95qG06ahkprNc
90J2JrCQ6cEKRnSuVt6sE4MfHnXanJqQwtEz0vl25E1w9PK1TKSYwgENpji7liVF
z/c+y04imyb3OZPe1TX95orM825tMc9OShExgbS3OwZy3es9L8ZRE6FaPmdxJfC4
C1U1MVbOUQ+7SHIbTsCYC2nEFe2VW6MvxX+RzbP2APwJYQVi77zEKz/mj6HT+A+R
vOSJotpBAyn9K3FWMmgMXG7EWFRX6VLzxIZvN2ahFRIxyPVTaQKNBVE5Z9UlsdxL
tDCQVYScdIVjKOxK5Er/Gfb9RVPDybcyuXvYDI3AxAnzzqU7X6bwpLbpMP93F15w
wRob7tudQKGXJfl+5pxb42P8qYFS8ZWI1VY9p6eUmO+ihma3D+Nw6QCi9ylGI7CE
P6uQC4znEyPP+DVVGOlp0grmyhq+LWEym8KWve0nXnQjzG0M8umvdtK2xFCZANVl
4OeN73GGq+6Y4Xr9ep+/tBPKZInpi3x2C0nojTUMoxnLI8c54dXBpoe9J41acNAu
eDZixJBUBiZzMPwI4N9qwfKu/wY1box1qCCB958lubKLhXxkNTSTDh9lr9MBFM2L
WnsiEX2iMSMRdz5MZDBnZme93a6PT7JZWWlh/vT0foOiTwC9x0yTfvMhxDIUw4BT
nQ5aKIhaOeJ40NLq7+o/nhtrJIw8gPGZjwPaCZbCFYhoJL0QbWfOWt4LPn08F69L
+SSIPniki4pL4layHz5gOGjWxi9rXGu03LN81aIFRg2RMa+w0Rtl9oCb3I9WUp3t
cm9bS7DBZFAGe8ws8ZeIYMREZpkjUEiRvUtt4Ld4Yq0heMRWBZvg5VRrAFGard+M
0Dy5A0SKFzTFZHXgJp1QlTEMeQ0Z5pePVy0StW7ltzCS1iNX5uDLJsC7rH5Z9B44
BL9UmC0l/apYBw0CI0sFSU4mYbEP7gy8v15WTGzMPNKjizf+cd/gkQggm/2zkxNP
OlOCW7ytWbLZJpVAI5UhYnCKBF97Uc3Hj8DsWF7XH8I8A5KHA9DpYMKST30mWZch
jE4CI743XeAMLjV9ugauo+v/QmUhZZJkG3GV7hGkiSf94/JBPqDQ3fELGQTnulnX
xQl896bs5mRULeJqPn791bw1K4ieYsn9PwalkveHrbfAtGyXEEXiUEj4GWeNXn31
AgetxZ+Gv3quiHrfwi4ehth4AA3lCXL4Hmn6rIW43LGQIBdYVq66ZhpnsBxFMzR/
jLOpUDVmvArU3OHCUBAy0sSZZKBIjhIje/AxRM7OgxfNbl30hpY5TkVsvBV9U5gy
KghttUsixfSNy9o13ybhvSgvGXPhyy8cJBmLEr0M+yiCqL8zNJpnsglpRdGSWgLe
1ahN9RXgblWvzG2hvE9PwiJvqkxOHByUxv6wr/10svBRExu3js+6bJOqHyirzVaH
KoomCVch/StsvVGBQ8jhtNAgP5ihcD6z860tatUyilzawDlbytNVST1fI5lcvufO
JxPRoegYs8VNlL1mTlr+0rdNL4BbzTfKvWLerZBf0YnnRJrXqug+aCRaAexujaHH
7YTn8KEIMqLRH1nYNWtDy/OF7qYRqKZQ4k/GruaERvE7vdRQO2K+fz8cKBob4lYO
SHQd31taDLIVd0HIzPRlgy23hLB48TOI8u6HyBqW5BjsdK9l4wazOliAzMrrfRH/
R8/sbsCrtBxx8V31yGEPye8u7G4vfyE/TQSqlfO7N/dvqaKqwUTP4xq0D7ls0iPL
LGdE5t4X/tnhiYQK0i4DZxD7H5zljH4OBbR68ZgFwdlrO6V9PlXgid2XvPxIjiI8
fedm8P7D6vraO4XkOfatKCApg4dPngug68YWGG7xycFVJjCs+dTYDjhzhLVdGSfG
k4+jjqBNkSXRdkGyDaQhT/IwXDK0DbDrjv7cZaoeai//qY8WVzwnHfLeuCL9bw5i
UvNtmGc3sBpOpulUVUHunj9KeW75m1WubDfsGI9orxabLSxCCmJLcHaul1LupaRf
0xnOsYYpP1iCwamxK+dSzAAFYk3JPLXtTXUu7mFyVResUknrDKoFxXeXfBn4Orqm
phC4l+2h3IZhe7NWPlVvNelMx04U+izZenQG2lMc10e8BPWaYiuvDyqgDX+x/mu8
AWd7QLHRh7JBVdhak3fdjDpCPvbhx6LokQS5QCwWSbYi79GEzbVKMkVraxbQbs13
dfDy+EpGCmsBVdnAMGFVZtr253oT/Bux5mwD2aJFBlamBQYLWk8rgJ+GR0NtOjRB
miTNWRFLru/uhVMdEqJiR+O4G1jKWdv7Apru6jbvFnpz3GP6NqJvorSfyWQtKHuZ
+Jouptsia+zAKhlOprt/IBRmlYcEk/wK6bOyfbMFSS1GfLdFOL9JPtcU/JdbqPL8
rLQla+OUnapELVqN/NkHkTVDGrXwA1SGgQxDiygvU8j1PY9dLWiyHkSOdhGhsQgS
y3MT2QPJ6pp498K3hpKviStY7dO71X4Xs8tNxFxtn1sX/9WqAxFg10hiJlwNh3Bc
XKlPOQ8NYeThjymM8eW5oGWonKhqXR5OYPCKfZSnegDkgGBNID7W7QkXra25agB1
umrj1777eDIBcH6FP86Fk4MOygnYqghdSv4FwHhHTj0JMbELHYNLA1Uk5pr4z+cs
IOoIuNXLNesAspphNkf8WdIODYMtAcUVf2ASkVUEVzUkRhsc3hhhnBsPH72Qs35c
MPR9kwcEl35vDNGAuDjZRNdMGDq+vk22nbB9rUbImXDoAVb8caIhZP7mWtZxsS62
UOSv4UbvTXYTF1ONUEpGSjKwLCLg/wvqcl1DDAF/ePXLjMrREbmK8/JyWLfOxKhL
u9nQMrVWxNUHTl89g/iFfck7GTRqy4Tt3N5o5AAUFfd7O58iVoNF3jk2dbwswH8d
/DKM7Vcwg21wTWxXUcnROZO6aBFRP5WKGurxEHrcnQemjEXW6PhJH3vcJMzsAEeN
eN5+fBMPwm+008hlvTtNRR6WC/dC3VRkQ3TI2OTr7JPGP/c31vNK1lUESyZMTU1K
CmTUs8Le5iYuSeGqIuXJobtkmR8VBEEICsJmJMlEXs57/mC6xE+sxGPCtDpl2PDm
gJwT1cxRzs20xdNqjECyFG/jvHMQwHRerC3H+V9g2zI4ygCDyiB6ycUET4/ypIYJ
0dhn8T2sBnYpzTAtGEHayoNbSNnSdLJ6eHsTQU/SeGuakicquHuED3J7/zK92+Fw
ssKN/SkMhF8fvivmktmol9ZcshbOJYRCchbyIg6bYK2Etk48GZlf0W/Wk8QuI4Rj
/OCcxt1kjkfBOxzNFLqBW6tnBz6x+yGgyVstc96q2Rh+L+CVlMDWzCkSdBGWU3ty
z3cmpru8LyZ9CVzosu90gvdFkburgaI+sCaRxsyLTAlzAtIKxE8oKv9gDDrpH9yi
XJzIWSmaoSMBrpdkKnzvg/u+goIQeyCq9F6bPCY+dgPLEi/BTb6Gwqb3pTfcYsTt
3qS85ieCw2nZTNkAKQfCcCxyBd3d/PVKQhsE6BvxhmBFKvtjHtMYT7xr3cLgoFRk
bOqRBF+0tH7d0u8WoYmTD/wEjLLNeCuen1PvowUAa7Ud8uzZGIRaaqjILJtnSbkI
2seGemGbSL3AAHfbZKspbT4MvuLpJnwQ3f7iJKiBmJQqYE3nJoSORwwaJXs0487S
RWMiQjjUUNTagMxq1FpuEwkdNbJoz18kyYcRmELpeWITZcbx69aj4tkJcre7k4de
s9JDOoya+1llSr1w6XpIx95rX9HfK0EkJ3m7pSRkfYHCeUHBrOaakQjrTBqzOucN
0oquA0DgavaFrogAKYDu9aaDUaSJLQKTHWQLe7MBIKuRpunC+HZRb+TxJbNTCxSO
pcmI5N0soDELbC9vVWUIb5gLAApy/Wd8QvWntnyryU6Kv6qz/A8X2JyJxV9nVj1g
fYCDfgsm3cYJQ6uoyWHaIDaJYpX5d1NB37W5ZwHnCuhjVsT65F+k1veZa43JJJJ9
R88g0Bh6o/oIQTvvQepDhDhe26xLIekZ0/aROeklYh6zxPW0a/RHYUU34xK+AK7R
Ji2645M388FuIcU9wCfVvTx8I8X22Czo5nG0sNMboho1FwWodaFQj1SyBVG7rRXB
+1dSeCi7GBJ6djABcKe1JBMbYtazNmA4NKa/KKBETnWbBiC6fEiUo6UZ0FlcrBDv
aFMDhKHzPe1AuEYI60xGmfB7J3Y16DqNad+fGlfbRao8nn/3rqO6gaJaX9axJjSa
JaAMEgGgXZoX9bDlgo8kFiqY9uNAslJrgD1M4O8dG0UHdB0XTUBCSBx6TcmpVVNu
Vm8NzXnOY+s0gFO+6YOXoTB3OqATa5JLEA/11xUrdC7XX8pRrFp0itjXi1NXrY3u
fAD/bnlVl4XTpusoBVnbPjs9U+Tatf0C2b3z9mE4QR5XgNVzq5OH0MAv57R3TyIQ
k0Z3RAqoUfse/mD2NHlZ+wvrTSnFYtoZU4eF/+6kChR8/SAkHjWGaxjtnI5vKewr
n7Zp/iq0oSVF/iEcAu8G5piEuwjoPPT/+hguZ1DwBk9cp3wHIRsxZuAAlKArWAJ+
ep2h/ZLVbcT0WPFToJlFX35HKSBwvhcAtgzn17G1Y4QpASxYSuTzcwjC9vsV58ZO
FYFG2VlY0TkDr+6TlMkK1WsZbqTOdxu1yxRhTOUdq/KYmgyw7LQDjzk61BYD140I
k1IKTJx+vXDfum02QhhGcb1/5V/7dDjKzuZ5j09gYXVQ+Pqx4c8UgQC/0SFLEfMr
e9Pxgh76cqCyte8j5B6vNiRqxRu2yJytgpZ/CdVV0wAf1z9caqWQWliumHtDXw5j
djbpZ9ZUDdtSQgx4t+Bo81jkw2cncotngT+PyZjQ6bVMfXQi/CeK1z48A9NwWy6r
9GuYt3wh8SB26Dk0mV4uoJFDeGYj9zcXrmFlnlLhiEFVjdJDTBVS67hVwozgyLoe
ua4X3exClTxBFNNKlofwCR5kXnZ98PG23x5DE/00QvP7n+7UtZaHvXEk5im7hgus
mrTQibTE8iaOT8LS6RjzYA3W9sssMMbp9/71UY3P+jEf0Te0KUNt8uhHBDxm4h3k
tBbXYwzLtPEzoIWwPIWgvL8cL4ZcdNABrxhIj3Gxub4hU41Gkyt9lEgDWnSxweUL
VBHo6LAo3HiVRzyYVfLCUhRE8w4iOujTlgKV/h9I2rlxvxSmybx3IoZiSl42Heef
iXE7fWe0/yASx5EzURROwcGpxaHBnAHOeNN6VJxtWeFvJaccKDc7ZvjbTq/yHUCm
2Bu0QCmhjjnSCDzHWVyLlhE5jhaHit6E8j2T1jwDr/t9seho1Ouxjv7Wdk7Nkob4
2a7C27xbWETfw9GlyGn7FxxbRijPXbAvtjXlTkQiETjYmlWRHEzGQga3Ve2Oi3Mm
eU0oh0Yz+2qGy9pAwZ3V71y/WSa8jtmfhgXyThtm2RSoBh5hYYcFx0CzrKdTkYFp
fdu5kaEFfWi4jqQY4wo5evixtAyHt+gXFAxWox/vUCxXv89zgiNc+vQpfDnUocuV
iWqbRB3SJ1rjZsI67YPo8IGI8/htfMtrJ/nJbrrY+G4bJrpwNF+QIqEHNvOI4zR4
+OmDuf0JpvVuVEccDj7Uq51AIGXly+2t/9l304WwsiqJ8Bia2cjZXeaMb1E9RC0b
ALQQbsy/XrZeduR851tctOrZr19vlQ5byBdCDbdqoRwZNIeCLulaSJpNP+noDYKg
smgDPdozI2Hx9CXgc8PppuC8Nqwoz8nX8SanatIYjdcDMmG4Ide8m2XqYLTyUKFy
XI21AtX6Y7V0/r4cPQMtVXz+P20v0kxmlF2PuGQEP0Cd2e98PPn4lR88KU9Y0Tda
SpGh6C3SArqcstho2l6dfp/WpVRk8JfIsMeF6YdP7DXJk8QGdTWJcoYoGj7VtO4d
XcKCWPmx0jOETigZjkKZoNBWacs/9rFvRUjc7XIq5eWu768GxlRNOVHOSQaIK3FD
hEt3aZFjF6+7aB3EbcEty511wEJ2l5DYX528BGPLF+D4KtSKplXfu5Ine0CvI1M3
pFWIMaBMqGKE3IpcwsOehM+pXJ9xK/86NZQg24ZsVOGZJDWr90dYocJZbEZlVo65
OX5RB9hH4uwWNhZ3NGcXW1ZXR68SYlb7eTgontR4qeQ/PMtQVO8oZ/KvQ6RpY6h0
8twJMsLf7uHP47XkwNZWDQy2k/YKoglsGHD0u/xwIERvGLXt8ssXOia68nth2oHG
PiXeiFXJ8PXRTcXFLSeJTnBNlGQ/oG9mEpIy40maGJTkh145R2FWKOSdoTUnSz4e
/8X5HYiPF/Nx+94AMef3A3MoVBbVLBpoAQkE0cncxQy8Xj4ysYC1Lb4gBmO96T/x
CAwaEgL5Zh9AieLDWoCV0XuWM5YJSqvl6JiutGXxoRU2yu7D6qoARKrJ3A9zW7Eq
+0ndCr/wv/giPkXQIEMtu5b0E83WwezvgrHo+oYtycA8WWJg7q8u9KRFOuOCGwjO
BdZT0KKaOeCVmWvv52gu+YdNI9Zl5BzK2A2qioI3KZs8gE1UwgzUDcsDyMQAj/Iq
0b3aaCIEcrXb/Es2JJuBcdgZI0xeIhPTElOtfl1lQ4RU4QBeu0k9n/ll8loE9b7q
ueqzonUCgdltHim6rLGtQe86hm/pT0lO9Me80TjVSrVkbUpQwj32NEpJrHfR7hed
7thMNsgP7iOFgK/UDOQe1DJwe4hY2qs5tJuJOe8+9+8EHfc91UlgTk5VCk3oqoMw
A4pLW1ZYTrg+v588By+v/xtPv5Nl5WO830a/lu0jas/QXzXLC7rb6cXZEiN1OvSk
zdDAlNq0VCnCYu608NY1v+tvW+CdV8qGVIpCqAfUuU0/pPO3D+BTGID/zu5dDTkg
RbkwHsQhtiw63IwjOEnMBFWwcri0rJQ0gPK2LU0PMV4X0N47+SihefGxVU1oadaJ
yhOxsy9M8qZuQ25XqXwVsF7xGJTo9VSdIDgUmM/wrJ3nmq4LatMgglm1sBuKyIdr
0CqGHGUKKKzb/cqF+vAPPc5v0eDI90esicYd8b+RqHFNmJV+3Y8ejQOzx884ut7j
XftP89uH2A3E8/X9WesrdrqgY/rqn2dvJp91coLSbdE9cLAf4PU1GXxFJ6GcPOH4
NiFfk1kkr64hhDGIpIWpKwf8nryekpcpqn87fgj1wv2TkgmiapSIS/6KRicBc/fF
is1PPyanOJBgEXgpv4ciVwZVW3aQ4Dy5jAqjYeGpB5P947fY3NBsb1gCGayMLq/n
HhkF5uYu5bVYHre6jnqHZ/RUwE6TR6ckualqOmbUtajmizHvoMY2oICZcRHTOM1A
wTB6rVk89TuMNwVWuQhpTxS3jaFHUylmnA40RYRYqcBIMOum/AUWJCyZxGnWqkm0
37HNojRgvpmVpP6Q0w1+AdGnqcckY6nfko693Nsf2TM8o/zHusovWHUUC2MlMyXi
55VDO6HsBemCeqyJSJS5WfrYAMgDuIi+2omAiqAfsorQOrjUyOPzZ2QybCdqmWX7
QCqsm19s+iB4VMeVr51e1LGKnijv5yPGAa+LoYLqJYzDHFEQ6Upke9rt/UgUcGnj
twdGKN4zSqVsUnsDc6Y21ZylQh7ijBBB+s/cEM9I98DwnalJQyLrc7QWCw71tbmr
LQBAh5P9u4qQRMFkpWCkxDSqxIboEGbFoMb0lNmi29g/+hXIHPcReBtjXpXVOCIJ
51wUl20eaTtRl40Zf3K+E2Ze1plOF9eHELAcaD989AMgZDrmR/wgt4iFdWviuCZy
B4hmdk8v+X8U9D4D+iVArxHnqVyNbu9eM5OrFKDy1mzgpYHeSSzHyhgu3NrcOScm
mVeNAAlmCn6BwxYA6prVeOYGGhtnuXMMQTH/QZPAjaIUpXO8HcXQtcFxA9v1VycH
aoKha0XSvkk3LoEMsAvG+8MNnn7jA1swX1ECHapfw1lnOmwkmGXB2qUU41LQ08Ea
0Pklaf/l3nlUyoTLE4iHg9mzdrUmpOdB5nVn1wWqdJ9fCFYxF0gRI4c93NInWm1W
/E48e1+BXOHtjaywejgaBSwN/O9v9+QdJlP2tECQShtteP8AmpATOlt3iDNWTWDg
tH2BXBXNmgxcHGxZKvRbCfYXAe4hOJ0RrDcqAThd7O3sqndvzBo+RTOM/Be3MyMe
MbtOKuhYwodxeKkjDfoexuHu1bzN55WiLLzXkLxgyx7latVscp2qdY8ZH+Q6jCcT
9h83K3bnJB7ZYphGQX2Kuqt0sOfJzzqNZhiF1k2K9PECm+Ms783HyAXhJBpCQd/G
/ZqTfJLSZShFHsSQ1AhcX7J4BI8VbITewxhCVJTYn48oXpKnTL6mM1QWHAAP5VGK
Iz4DKlEtYg+fKnWO6PdzDfAiKGgzZb+494v81Hfh9Ctph/ShrG/ukUNDbYOZ3d4A
AofV3XAGc5iScMIruIS++OtEgN3E5lwYdfyoiRxdeZGcJtSEjkZLcZbS+iV8DJSC
rWAc+m4X+fEd8RWzufGl1tvxdPnv2f0fFiR33cQihw/l55Af8i7S74dRtMZmW1LA
hREC1bYT5zqU0FcXDANlpCdB5oteGJ5XUvEcDYXkzJaM1YNPEzgA81vBCSSggZcx
XQodMO//qM+loriBB8zls2fb9Zam4hwxVHEB7FWgKN1MK+1SizGC+ggKPFyxis82
NIjYGCeR9utWqHRIQPeVq3OhWBf5Rp51hfwx+tSulQZcI/2y/sxRf3WcZdR7OCvn
x2mqgMsYT4T70+RLWbK7nMEM6rLSq6vcC4mUAVNQq/z8qnA4PPOJSUGhEhdwOPZ0
kaJOEIvFAeG+1PwBMa7kQVK/WDPIKIsjEgrS9GT37S6bla8R921Rc8SjxlMaGRKe
ANUUHIDt3q4ILo+I+QPhu6LH5YiDa5h8q932Ut0rjTTbjrXsgPKD3HePBZluCwJU
5w0f9k5A3gGkuV8Eyvia7urejseT62zsYPZgoGFqH6qTillfv+C2Xpzyn+8BeHPS
T+HzS8Qu7ANb49v7MexKVaaDFJ2VBG1VhDqaXXzVCO3uifpWsqXXCb6AcmxTCWV5
Vj8FV1b6xKYLpwoGAoKl5ZlNJC0JXAYEuFE8Uu1RPCqCJUz1UDoNrVCs3wmANnM9
Lq8yTDES8C667E+WZZMM7PfLVDGIhxSfv3GgMSAwO/D+61fOgKqInih+D1LCcIP5
H0PNs2pgitqMAln1q9xWaieTmEcoUC1n6wRszLe/TVbI60eFB/Mf/bAlBgJHBZvJ
ccCeHRGjFktCJUyhg9c8LaTBWK24FG+tBiDmXl2MtQG62gldguPPnIOUK5+7m02m
vxdlB1Vqtbrj6SQCKcTo6jSuksg0/HYW5t5I2KxVMyfbSq6RScG5mKyaQqz8GIeM
AuZWont6a/JTryjnP7/YwVuVrvmMV554AZzT5J3IVVZNMbu8vhehVzYRbWrDETU/
Jy2RBdKoOxbdTaMZ2iXbIpVD2QtkOxMKT/6pAiP27+sH3zkPkqddFDGsLCzNdsEU
kihUVjRWcupUz2sTWR9sIIMo1FwF3BN5yagovrDwupnNELkvkaFZLAanb8A0uc5J
kKvN7Le235eKFpCYNSllpgg+hna+TcBrPeqOagMWS+5ooFJk5YOw/EIc6cGC0XVF
VxppvWvvI8xX6icSbhDeAo7cvDksobYy3lfWWZ1TvuKoWRKXFjt0tSIBZ8qx8ab+
iQzAuqPH5AzE9bMOwbxG/7P3iiEob4UcA0xNknpzOR/7NzJRlA/oazUfrXS8plWz
GEhCAVrm6lbUVU9Wt9/bE1equCrS2JxrJLNth0nNcUoUo9lYUL4uZWNbDtnkNrH2
gtK9gjhrZCER811Ht1OEouo8+0XG8PeORhf35Hh/Iu8S9F9wFEM32LMrA40CIukC
wVtpywqLOO3aZbyMO2pJyicgS0f4aB+ovRW4CRvDUuGO/0TtyykiWMiGB4n0Ef0G
WT7g4DLLj1CfYdIWKpBeaf5y0gZ0bh+UeaQJ91+ngQ28eEWKe3QBSfJilIhVDHFQ
xyhgighxfZAclgUDiIPByvdw0uaA7okBCHXIQ3kRslneH7Fj9/VBTxhcdzDvF2tc
l6QIkiB2bVgjPZhhUxQHYUFfLazAvef4MGPc0fVo5dGioBLMs7zvEEnb1/G/vKk7
xFJ5b3KsPs5taTTnwT2Rkt1cc6wG3PUmJ5OlNAFwuSQWtJFxOGo+f7uL7a62DeY3
BqsxYTGuptqRdA3cR6pltoBl2P7ICfkpCGsNlym7feY3suuk4xZOnzy7EiZZ74yo
47yMz4KE03roh+v/M7PybU8IJawbeSe/jymheOr2XsQ/M9ci/z5ZRytwPCbScxJR
Ek4RXq0eceeqHpbLinBVQm0NzyyH9HGXTPAcklC9Wzd1p2As1af2W4Lp0Rdy5zfy
0OkgYEfD00IG/ik6Kel+yXMfsmv2Yh9/7v0xnhj0p/gbnubah9TB2eoZVz1VGr6m
0pTCJcYvN0caZ0PsUt8bff/A48j8KG9gPejCWEZZwS0+K1YtoaETUgdNrJ9Sfqle
RvumBthaFbrgwDrMHoRtiqb5jUaskrz0Za5NF21WQ0epMTZoCfzWy4Q5Fr6hHiox
3/916Phh6Hkq0IdmcWnHB6IHnBX9TonDO1gQcR25GgCwinO9gX1BGQZrBSJc2x+k
1z6qkJ9bdKU1Hwbo+49wSEQJY86xwxcUfNWhVfR94H42t9XRCzC6igMbCdADjB9r
d2b948pg/XRZoJpjtg2oQITqGu64hJORy9rQSIfyiC6VrtTH2qh9uZpfBAthGouC
uP1l77tEZ3oF3NsbFYc4QGNz+0Sea5n43hsVRudKfrQy5ZHmEMLWN+cgMpfzOd65
05sN980bKMG67TsVXGdwHiwQSSQMtUKYWfydaIUbP8Sv4e1xLV4NYX3MBeFJDhI2
OjNql4rKswr0pRG42oOuXZsuVlj+DQaWSUo+6fkqtMAsnu+joQ14QrGGuv1hD/kJ
DoafJz3MxYop4qonat/qvONtoohiSqCqqK8rrMft1ioPCD3LDG9AJKZTekDgvsHv
d2Wn3hBH0ra+QbVK0nw/nB9LFolJoGi0FnetuC3y7bKBFGUn3cg5+jKiaJsoAnEx
2RF3PqXl5lgC1H0KeCaTZfo6Ih+uNJEwpJJxdJGZmJCGShQmej+rMo5x34ceezIR
Av8sG/8zJ9K3yWpz3sLr6kiRoFhSjcryliaA4Un+QydTDZRQ6VTXTuVM0CDYuL4u
d4fpM0di0itFUqRi1arMD8sLCVfS5oorJRQc/QmytRb8Yg6vf3EO4CYz72co0dAm
0lPh9VWKJEjoizQT4TGGsC9FjqYGaELEtNoOsEfiFmVyvo3XjJhgLHZfsvUmGKeL
7Y4Z+KY5afIn69xr04SWpsOLGWBIp5szR/oLp5y0QBYk/nib+tQGdEVhXJ33M0pD
LhYZJktYFqZipmbOLu0H1nBI6hpthbLro+RpzHPe6sdNh5vCWi/wNA8TTkGoBPc7
BqTY8enOb7ZPfo3vt1Z6NYPBkWmcxF+4WBHiCBMUAxsF9ovAQcsu0H4jNSH1VNpE
5qgdFI2a40LD2rUNgsNydxQzdED8h4Yv5zgDgaEY2O/miDToTBXHpLhCYuekTSEJ
ZlhEmeMIWUOk+OwUpOXiWeB8cWlzpZXPtiuXGqmJ8EaXP6BbYHL1+rzjnNcX95Px
daMFdMkfNRV7vnzFvLX00jYnuIYLKP5meAQoU5K5yc7CBAu97HUOThg7I7I2AGtl
0rAFDjvqfG/P4JT/aKkfrK0wmxZihzx38bstmxBybOq2jt2rPJPO4mw6dMEAQfZD
vBpxfNJrAuhgmGaREJNHlmaoTLfnlV9YSmXb8UPc0Jr1oylqjkqzK22AVdMHhVy7
mK3Zofb9pihju2YckWd73cDja8q7dGLS5wc6KX0lr1xMIKU0WWErMvVsjRHO/yNr
3ZX7Bma7xelVtQMqNeVzL96HQmX1q9AJTFvMeu1jqwS+wtqmvaxRSg6i44bPKJsC
ZGZIO6WZUvOeVfoa1Cq3wg2CuKggwxFpLqfb7lcFPPdnn//m736TT5N2Ut5Z8Znc
RupS1pNlLBJxY2A2UlQvPAJGmDg5AjKJtrozzPExArIQJ5fvq7VL9tfqkSZS4gFI
LLYIo3nBpbaUxYlFC9k2H/Ks69rkHFvnRRVJbnQ2/8nlClmdGxZ5u1IEeJglgxMa
k7Qb2UdPqtiSlhgPBQE6etZlGp4cu7QileiNeGVgY3+nFN04JxtcpaMa7DCsAIMc
zJl2SyzQW4G2pyDYFmoVJuI9BmWgGMiuoGoIA/ob8JhR9/y0CVfajMQQtISArBE/
F52l+rxmsADllWdxlRa/fJ3aHIYyIgEZlGMWZVrZY53U414xMMStq8dkxSuXphRH
dHv63PyN0KwTVVLG8qRfQu2tSuvDZ2TJ5tpX4U42hNlN5A3C8IgXNVYPWuA3Mzcr
p9+dt4GkQMSKWQ9BkKB8Q9NDEDO1VE/YbHdxdsU3KM13mgzI2u4/LRCn2qlPe0AY
gDKL1O6w+/LXSgKEAJtnSLJ93wDdhVGehk5SblE88S+Q8PzV7yG6FKP0+IAO7pyY
68KrABct915Y0Hg/0Nf8/te0AsURS7+uDY+Bt2T/G/2a2QS178Q9mskAtsr6JbmU
nuPL+Xc/YOVgH5ojg2M9QPQ2SEb+/OLRwYK6yY0kvOGCS+wemUFqqpQfpeMgwaRo
N8J6G5WYS9UIWc2IxQK/3ksJJtLpaeuDcxqjDhQ02XVRv/8I5IPO2k4j4R4GlK22
T0xTN4rXa09TSmfNTW194WhTyKwnL3EIOzI/a+7DOG78UwIj07vaVfZuP+cGb5a6
44J/skwoLVS6g5qtqt5oReLiLwjNRA/Q/HbgQ9I4DQjkhKJR8Eo3jxKuMwU+Wnds
0X1sJ+GqiKmeehgWVT2k3XsoXs6m3jHeZXzTYEcxkp9hPU5A1h7SfWn37sV9+r6A
HUgzJhm7qmKSA65OmyS98FlHZ7DBZVXHBdCbfJv4TB4i5B1lZe109BdPe+szROgB
WvcUrZjRd43Mp125h5xL7YH/9AbJOAObijcDZJFr8IXQmIzRJRm7/nknWFxzRi6F
+oXKYp3tNcbtWFay+0mfCDUjugYEl5s1XJaUqOqgT95H4lS/c8I1f3iIfPTWfT4q
D+/nI6poKITLuhV7eAUvlYM43ViDaH+JpwC2XH9SDmgLBbO6ypZF5EUUVMn7DPq9
A++26dxyDDrKou2fUyva1fgaG9wa7VYFMnu0dFLA81utTKR8bZNXfvB7nYhHuaV1
ioUte69LzG0Z5F5vPDIIgk4SLytXiSSHBJ9wJf29fFkDCE26pbrD3/HoaPaiJSt3
dZPbgLpmBvXXgA04auvMe+yxmQ1ATYc3nbj0dvTVrtF9GchztvO7X8Zrs48eH7EK
rTEjagCSpz0kH/oI7gDJEjMFwYCQ+5K4SECciOVH0gajf79KVuHMo67YznQLmGT4
mu9fzkQF4ETzjZ30byFHIhZ9z7BvKYr0TfXHbkb7JQsyW4Wu2nN9V2M4IG5ZT0qa
mvhKQhsuWQ4FaICHmUGx69+u/9vVn5QymGTI9Op6zCTINiNUPPjZOz0iUx0DWWNA
M0Yfpk5X5HhDRlhBfdpLY0e6rfAwvzWomgEOsodmvuebSaKsCENLSpbaPytKhVrh
OnJFw/Ue3+GxA09b+vOPEKIYzmEynN5ihgXNmdeRgZPlp4y+xI6aR4ZkL5DLVvr7
d5mipY9fy3/z9lfmDGcB5G+uvJnhvpGWg5AOv7ALUKxV2nhwlpyUqcfX0OVywSCL
7v0mAo3PoCmcfEbbxAagr73v9jffTbqCHl07cMHoMDHC8MNffQhoCTXICkMVwCBp
dat2dWsTHNMDj8mrSdfl87ru9gXi3TFtH2u4BOlKYuUzgw9Uga3zw9EB3lE51pC4
TDmXzp3L08hbsgd3Oc7oS/Dimp8q+RPtbyHH6GSTlGFmvWGdV/FPyAeH7vBoWYKH
6mxrZUAGfZjqq4klQR6RfvNKPEVkQbWeUFFqfR0/a164yfmPKwYOZLgtvfumiiek
gq2CO/qXgMBaJIGZ8FqK7rENx3F287clpr9/E1Dw/pm6MAv3J1+A77ggxlAUBNFh
tgpdzIttzIeBbL3q46vpJVqHkAWPNrRE7Dogjq8mZ59a2hsYqtHdZYuuVJMLrHo/
tDFjvQ5Drrp2X4KN8889Z2gaYGQRGdotyU7K1HWOolewB5W0D7PiU74c6eB8TAOM
UnYqpKcY19SAeGarsaJUu7S0pY9Aajw2G2hj43JAwCDibK76RZF5zXp2Tq0gV8nn
uMaKxyHOoed7VQw1e5IbwuinpHdf1ZGgkynRHRYB6ElQSdL6M61GxuHvnQv65bVo
27ItpOz8zlENwVnzG2D8rozufpAXV2nTh4e/Hx3zduc+EN7X3zNOHT9yMwsBC2fe
dA6OgknDiLX7JsEojruiEiWt7BaovucAzalQUFwjAHOeG4NLXB8Yvp1Avd3NzfJp
Q1w4VxLQXtD0adh2RI5ei137UfYLOSa2biyowjWmAJ0hF0WrHJ9LkCdsIl57vPpN
dL+IjNsnNcRe8DW0GATX0VF2V8tsNQYbqZiG4gwOq9ADuhGCdDHdlk/fAvIZ4Vlz
+VW+ne4BqKSFUNvPv3Gqrvjdn6dE8nV675qIIy535EAzvNguvbLVpptLnEAxcpQU
1owW/yieC/7/6L2u4tZSlbr5EGQHeoNPNmiVCa38xOJtcQbchGJ65635E0UMk0NZ
2Pdnl6VUAjugXhQ8uHiJvX2lXZ+l9fhENSq5Qid1LM6sQ5Hxwqug2et2lrVYUjf9
AM2mFQ+n3gu88rP/xyavvCEkGXNEKdSQ1/x1+oTxRgpioGnbGu8jAQFqZuG/G7QV
SV5uFAjLMqRLpx+HdDjPglTGqW3WliiuY0Jn2o8jQ2K33ox2Ty1W82Ocjle1QVdP
Ao5C8VN0mDQbv61ksKW6YAlezjzlJQjGzkmM8DwGp8ersCerHHWkQDM8ZMLjs0bI
XaeBY2BEXAGFqSshfJFcA7b4Sp4M+eyzDJoPH1XhiZUiPiVlQ0x4pzzfsTFf1Q6V
bEXEB98zSrsF1d39cSJgDe3/8fqp4wAeEExeiw9JIbWM9+bvOwPAS29J5GAzF8pb
+HxrE7jnv99T9PquI7FiLHAYbz5PtTbfMz6B7rCTE/UjzIrf/XeYKSe2XAASgA/x
Nu48O4SbMpYOJSbFvzAO6rG2kXMJp7xTA/Y0s4ZQf2+dFt2Zmn7Kk/xbYi/7U/DP
Fv9sJfZPfQ5NCmHlK+TeT+8Gtky/NP28qZeEx8fFkS0aPS5qs6RMrebz9+YK7A0J
GeWGDzxP9n9sMFVYh8kZpUrZT8GC8oRHbcLjnTpCELyQxyHnkcC36q9Vhm0BETfZ
hvbuU0NiExZUUEDEKNejJqCoZ4wXMvBe+oZHv2x1i3UbrZ8caGAwlrhHFMsF95XR
4OfCtV6cXRtB24tPWANYAq8imdXxeNEB55+a0UTLYNNrg6AwKOt2k0QTdHJu0PoT
Sr8n+L/IV7IQV8kjgqijWf4BPKsysybkq7wiQ+oi6K0izyfMW1TchaT+mx1cIhz3
R+MkJpL7HXlyED0iH3XoUade+wZFmVa80XKptvmNNF1EpG6M5lxJk6DqGStPIxrg
RcUPLQr+zt9waSZ5Ma1pN1BD+8gsvN5TOTOMmCwjmQ2XT0OhC5pCh4Goaq52deAs
G0OkMZMG2avnKj0Xc/jj9bIiVEizaAeBUeNdcdtvAYNFsQHqyIJI9bhlw32uMlJB
VPphJaVTIJUI0ZkqmxFmthWuJcZdvJmhH4mCQsvneWKhjYF7Fc4qo51NxGJ1vDWn
7hTa9htUac6OZ8V1bhJj/39TOATockhVZYyI3IL4SCMBNR2IKJI1SoSqZ3CbKZfi
iHouprPMqiAd+2vg4s5Uz9vl6RXPJ0II5b9OxZLXwt3bsEBAWDgbtZxix0XHvjP8
j2wfUuT3Gc4UdlDdP3TqFXwsck6UXfOIeQxXu60OQL54ASIRCjI+D8qe/oMiMWXY
McgLe176d7vvn3mDJlVJzHlN5oNxAWFFwMV3Gzp7JlYjoQaRxHSFRkWK4cDPL2bT
I+/D/wjM6Et6t8DeeNDeNRrjmpEX4HObl4NgpTmNddhP57ys0tPTLnA+Hu3P88rf
b8tarxqmjuyAMH0dJPdBf7yoD43qqg1jVe9wRcdw67FKaJ0T6202xk4YeRaZr8Sq
zHMH6MhNkuGJbOjaOAPBH69t3BGm2BcFN+Ce/5+qLiAx1Mq6/adou+cy+VOxbGM2
SqTJlIw2n4ytboU21P0WfsvAugzSRG5euEPyaK/u7JjcjgQkv7sp3FXkiYmNiDOx
zDvhS8yab/ledka5c9EeGTeVN9/+yQs3Mu2IUKC3q+sNh36eMLqOMw6JE63DVC5/
OllQvsVwaNJc8wTCNHq1Uu73xg5e37ZECMwj2SOhw4M9Ah/ZCeStLAPkpyKk5VA5
ABj9gwxhs+crqANYpVw0QnBZ63xEa7DhNYk2hAwnCsRsvtivkDIMm6Sm9kk4858R
G/fHZXEC5W+EAjntkhFtZZVWHSXnw/PvP5z+tZogkTiedpH2bwVWMmCNNQXH9qW7
CSSrRHaP+/Pxj7dhvZH+NC9ZPyUdLaEHcqaXoVjJ0CS1BVfIA51u8VJxfNVErNnF
N9rVZgLLo2XKWxM03dAQjGvbfLS0mVNnEoFNn7gNxsrFKbiFLqSqHwLqK2QcvA3q
v+O3niCFxAs633s/tC/KjPhZ38+GNc5awXhx7cBn5DKdk0cs5C9wyAq50B8gAxXH
LILqnk78w5x/OE2qZ1mNC17Y35aiAzVXjc22H4FtSyPgJX+cfLEWpoSgiddFavkA
SwWJSYDhIJCzK5L7PbF0UPG86OQyduSml6XSL9u5iGMhLqrZ/l35SZN9f+83P6ef
QqQ0aIB0rKGHISZApNPlOkdNkipbQaF3BDLJP98K3ikCStJLSUKHc218Oi6Dyil+
WAh19cvWqIsosWBsr780+c7hmNCuOYU97neTE6gemHgm6SrFOJ1RWCny/kUW/tvV
5Uflo5xC1qEY2qN+HKri+SP/jwe4CHLNzcQxw7GpIQlPYqBsicAAO7DXX224Jt+J
3DELak9Qq/vhODUBCpjM1791qcmiYDkdgSzgOV7NvEjhY1KXZ1BT3AN5rVfE9Bnw
G+53RAnJadJMNNVs8Dci9TOGHcGVaa5nak3dWc9DXsRH9HAMxxVEdg1qN9OGpQJ8
kLLBkd/HNC3ODtzN9fKg15fpNZrM+v+K4K/e3Xu+sUEhBOP9sghrwnAPl+UiHEZh
LbInRWiRY2Pr48HaFdw3oUubyNxLAIEwNNE7NDvcQQrM4wrNVrOyrW/Z0aKLX43j
uoLYvhmMg2PGevEUdk/oXPHHhY8620pP5FrzZSSdY9dhciXUZGWXaUOwxHxxMvJE
HzFuM6cBJDlFH7H2qziFdP2oZ1AIHffZA35+469/euqU/fvQyallRahL5sgv/eBY
oDiFCkCErpus9NangjyyhbYTCPPFHm69CEQCQis75+GKFMMx7M1blIaFUMnSvM+U
gXQ0feqbkUNLQA+s7dmPV4Qc+9/FzmTUy3N/iatGiahWz3cqDDAM/XFNQuCgxxOW
7hBVwoNOtYisaV4JjDmD4XJt3TsBWMl11XJDJ+YnGMD+H448P8xJCHyeULcf5/rZ
CLyCj8qvnO33Xdw9hQdE3etrzlJv9TvuBT7P/S1yUHgK+3Apq8H3/dcM/W7FRUOx
MXRP5w+ROYBu/0auoRr6p8Z+oxr/4Z2Ld205/jo9ADL9qOV9fvIsbfmp2nW3tUUy
X557tD6ur8Z9xs2AQZKnOk4lKaVUvYXmL1hYajhzWb//4f7M2mJsxsH7zwZRnwXK
iarmMevHAlq2CuHi1ijKZHnmzk5Kz3+4m3HE9Fyq25caIuPAgsgO07pdY/vWl6D1
0GQ/xC5ugPZX9wVy0HNzq2c821b6dVcCqbT7TeVUeXxeW0SnNOgTdRQUzTG5mY4v
8srlRMIC1H7zEuM/PeIBJdqlCwjX5VmCwj2cg04UEDt9Kn2A+pPHZeaviDxF9FVZ
m8vKRRbX8qA6AkX86r7BPiXE+Hba+S/O8DIus7VrjmFNc4QLkx+3YZceihA4xnx3
T+RULsnwW12TnDu+s783ckeTk6NTPOJcv9JiHa+loQctuiut3d+1oQZJiKjmk3mB
3c29KcJBeIlmvkW0Mu2QIniJVqeGuQH0X2R/cqOoDfu5cWkueJcIsXjrLPJmIA1y
DCAyemr0uKC6+eh++/5d94we1axVwrtgrIsSJS71H+Sord9Xg6H48zavhZgTRrGN
tumS92WBtRYPavTmf/YBGXH/CkQjSsm5Kj2Vas4Z84TOjh2tuTHcm3lPoeQkzTJO
+KRNvLwvtjZ8PD9vKxWntFP92FngbyzDXYXjy9O94Snp25X3D1SZCCmJyHSJ1gYf
94UDPkeS5AddetNoLhkmP68V1pYLqUWgR0Bd0NMkMvjFCmss/JHVIefKwP7zEwD/
wBYaA1llQ1uBtIzsv38woqD/+rH4H6XeFu5wO2Hmv5WKTrW249/LUTBwIMbP/Zg9
EHjdcsZvAsIixhlmShOK0QlU1QrVpiTMYPTFttECvw0WTkG+bMt8IUo87LHl3aB1
423EJTnv14QOpyWSBcavi7XbJfo91PGBD4euuzTbYli+wCgnHQQ8J6vmmGf29mqS
77YWyplADuxzjIvmLA+uAjs/ygyfEfVhNHN0pvH4vzk/LgaP/dM2RCtgMOarRMPU
0S6nzTDgxlvzIGPhCz4uGgAEEY86k9Ofnh5+hHUF9nJ+BBgb19HB+NvujkT9OGgc
SC6B0bHTJnxxvMtgFJuxoy1aW2+D6LvmoDNV5DgVadnGycR38SUPUY4eH108yPnk
XroOsZljn8vE5SiagdLiNPbABWTM8a3LludTTT29UIraifYb6UY9O76HVnzf8aiz
hDcqn54sASFIwf2NETYY9gogkhX/Mh0KH6gHg6X4OjJr/Re/U46/h9fKY12gRbCT
Le4cKVQqKHBo0F+8Dz/2crMGBA445Awz1YXocGQRfWLY4EBfSWI3Kfd2zzcBOe81
vIvEywh+v6LdWWolQGh0Y8PwPWs4Axkgo4NzjI9/z4bhQyV8cipg8hDmlNxPOk9t
SQQjj/mfhxAwcrQmhIDy3pG/gOYvBVjvmaNq5ou3v2o1EyOBJPMGGZ3eVRTwrhyJ
y1iGzIplF1gmKxjk1XadXAJDxSsaeiZ23gbLBCOrdZ8wvqzOC9foD2K3tQlWwPTe
YM8hNZscXMylF7KOrPyJGovYbzZvuK8JswY1bYrnWNw1dzhDbVuc3bdDcjIY2Ywb
JK4MmVJfLg1pmjgEwsoH6BUaKFXoUFLKYMrDOHQgzUVvLnOcjYcRr+Hadg0wn7ak
xSZoMVQbcWuMHyWqbCEcS+c5R6pWpJuglYIIoPHV9mzgLA3TnUSWwOzrXAhkTuNl
LPSJeRWJJ7vOVlsv4FCZK4TgdZHQt2LINu1cPpACKMR1qaQ56gTe1ByzPU+f/xeH
lu1ztFKQzWlnmYDshCR2hcbaQ2yiekEKKZNN/gOjEMeaPMoxtDiK6QfWi+Uj3U0o
wdgoQz58ULeuVN4RccNcIO/gCXxzcOWUYUFwp75BDg8xZOdIk0OTCaPZ+1HN3MdW
n0Z4oPRpIvPMV0hYRT7mcdvKHbV76EHdwT5MF1utXZy3Lj+o8skrDOsr4xaBovYb
Pw5z3FbUY5ALvr5c6pgaGybySFQAuDG5aq3XVrjk7wkIzF5L2oYVUO+TpYWiZuMb
Iify3ZtOcK/Yq8aJyjvH0s5Ie8rKNv54zIX6M6nSvLytrKA0bua25tyoDotyLD0K
IcTqF90ntgTbeNDlxx2Fd+6gsVHP12mXr/4lJUMP/SyOY7D7Gg6wc+IY/PdfKbA9
u8LhAJ2ACdTN4TwHXni+f3/IKF9LpA3x9kr29xwo5FIVxIyXf+ALBUKvdllAM55c
Z7sHyNyqIZR7KKerAfdSzqYnFvQEtac6hsFnpl9cgXlujTNAvVQclK1brG1TdwM7
I4BMMgUuBTlq870aVdkYKuSNhFQuqQfrFKWqgiQl7qBCTRFhCF6FY+r4CcQSXeGt
h/XnXr5J317u0SogbfSNxwfI8nkrgv4+3WioJhmyVEqFTZebzr2TlWavBxfI3veB
iYHkDqDZgV4sOR6khafB0CZt6ShHyxgWbSRiFsTnIQuzREChwxAAD5wa66ypCXMP
ZGWHyONu7KPMNB4K+XuIt9aphrVijuyDUHEqpCxB44NfQbRyDsXF3gPstuYw2a6W
OuMBd01Hb+av/+s7oupVvuVm/ij4gg5PSDIYibgmA4+3pj7DfH8mrCtMhKMsnFRs
n3x/zM4fm3LFJDk2Mn5D81AP1vTmJ2S8ZzLWmJd/yiZHz78qZDyvypl8GmpgU6Ck
1phSY1bH7a9c8NRNMV6m34M9p7D+GJRnrZJcZY90TEpoEvmiy/4fZARoXDdm2v/M
BMWToTznUuGyu6DBZ/C5JgYOvovqr+5R4pHpH+ZRHBmg67W5Kc7OQKjS4l24uIbz
5qWv1fkh70TxaAWPz6aBSFyPRKVUuEjSUM2iFIFpMxBz8E/pqclFm/fFG41eI3aT
Mjihx9tidPLGz1jmsaBdArhKG5EGKu89M1F2YT8all+oyNTw0UAzwhhXNjB7UyT7
JF+HEfqjcc2rmSdS6J40noQwA27GMAzdg8AedQQP/GjbFRglMUgqMnJiPc5iRR1A
brZKxEZVW6oJmrqvUT7LF48TDU4ZcgaPgR3VQgZT0GrLE416r8KEscZz4Ap4JM38
Dp7KkKgsKToKpAbutuMef1Z2CCAGG8DKvx0iUhsFP9k+X22uUXRygsnmfCwMXTj1
8mlEjlYuIRSRIHGmIzkFK+aukN9pvTWo9tzB9EeRSVJrD+tFe1YjhSPNngJ70F3a
VYWfSgziC6GzwQjCTDz6CUejebNQBqhEsl46Ml1Sspde3T5aFfPujmfcYD+LS2jO
oIT6bpWEFL4CFP3nliJHsaUQjezMz8I2ox83g9YeDcpFV1oLSX86XhVaePm2oxAC
mR1+lVIPd8Zd8ffLnklF0EoQwxcEDx1dtDUL+x43sJiVFP0EqmBHs3XlSaS3gBlV
av3t0PSZwY++a35dr1odaOWEzD4Hx4lBNfCVIN+8OHDL52Uz+HlhyWdzSo5Vl7Fh
BER6L3zebNIY4wqj8SJ4h+/4Fj4Wz71jnKNBN54W+5mqwJU5X/mOe+nHnTOi1NcS
HYrkwIm8av4Myq+hry/TQVgSu0Ork5ZyqMF1EOaQP+ulvfGLsnhfD+WuxD1j6vJ/
LjarBdQNlTUv7sybMxAKDmE9skfSLelFTci+b8MIuQ4YdV0xSvFo8IFbhNJyu8aB
vE/qGE20AV3/qEr4FcT5t+AZww4Gm1kPIkGxMHE/HBe1N5LPfbp8Z0nTYYkVc/u3
YdWpKU79TK50e9L5cQxDdvoGDgf6Pdh7TQ+P5Eo9xGJ/MO73qptB6JRWpR9lGcX0
KyMxr6Z+io8IXS5fzgHJVMzY4s8U9++3ciffAFthaICSQOEjgDm5wlLi/b9oMyj/
jAtBfly2RsR7ovRnXSf60Emoh2BlyANyyClxmGn/kMHjHXE+CBvlMJ8T7YaFTNum
ym0FDnI3ck+Q9tN+Nhe0zFDC9UcmOU1hLvGhRAe/z4xk5pont40xB4txljYPIFem
W5Kg6yrp444cU2EcPU610ozGInuNmV6MwXZwVEkQKPoF0egZ+W/o3lUgvugZSF1/
DXlRb3TtvbxCRARMr1XGyUH8be6BctUfmU032baqOiFtfsBC4wJsUbG5ibkoTbh+
3dUuajlXkrmY9ffDU27yoOe1kXpdZhjr+s5MaaTBzhxKr6I1Rp4qVulKQJBUO+H6
aedsuf4wYl9fZKXZNtZ5gU+g7Iz/b/LFcFm9GbLMEIW1xGhVxeSVqf8NL+Fwuj7s
1jnNyGPC726HCmmx+mGowd6xEQzMar8vmDcNgbrIqM/bWRmn2qQoEVFNPNc6JvwR
cI2cD9Tn0M8j18kV67CQMm6C7plG/oIBrml+teTPhrPhVMi9UsgsyiFyyc2sbOdO
H5sH/xaX+sBCFPyLEmv+s1IuzWQv6mDElSiBNU+SKpNVtFj4V7xk432vTb2IyiiX
tLkjnoo3CI4+5VLlqXBRPkv/ILbK5kTkrmnbykV4MHyKJ4nSyJ75uZxYh/f8mBCf
duVq0p5us5hRAlJkbV4sfjk2sKvdzVCzr4IwxtxalH2gjG5uR+w+V/nZePGXWcez
AHEh/oRMytxOknZ51H1VlhZ09EZ3yWy2jZ2E3daJTLYPB7zX7Mc/ZZOkRlI45z9q
KlOVvxRrK3OxtmpgZ5sMQGN8q1k2Mvx6oGV67ieVoxJead83wqACm4GFOgrhisPA
+G50ZT8zFkh+oiwnSkmbjSkOaFwQdG8pJbdtE/uTlMjsOehOMs11mpuqoFZhKfto
LkWubr1guiX0EN6d42i1aP0PhTDtXU3NAIUOFA3V1Y5OmaJ7S12mgEl61PQyuS+Y
5uUSAuqtYDYiLC4Kazy2Cj+iHYqAClCJhmBi9QR6INSm9JlxhwaFTwGPEnDW09h3
z/rqEa6SCAc979M5QwlOuiqAFsSnahlu6WGWnyhmSmXX8OdejnoejNSipZYjn5Sw
AxKU5DVKODjECoVRTYkxI6BvzVvC0JMLj+7Z9nKY0sSreK0/53S/3Tn7UGTsKMYP
+RR4nimzCEMkM/DOiNoKDUPydFqDtJ/yGWIoIB2UhyHGSStO8b5M0vSf9Kvil4hr
NgEd4cAeY2DeNW/JYRwPQHVwDRSTGcefplyREIn++y2M+2OawQkXP8HwR1x2aaGx
NAl/ikXig0+7dV14WLY3ilejPD/7Sxb/lWNpq0KhrJqiixymK3oz8lkV+6EB/mjh
plIOn7EDF6bGWkkwMynNOPCPTxoLh+/Gaw5D/LhfJmplHa7VQHW8RIl1kkmoYWwx
JTNoCe2nPtH+xgE7QE3UH/BPxL0Mab6cZTXbdjrSB9vPRBtUgiYclyu4J6ESlXwJ
22kLM0z4JB+tqaKDTRCixQesWM7RoEZJRPzUYvftJf4q8VpqwC2+Pdy5UeEJXI6L
3dSsMwW2Tzne4ttx+RvqQX1jUOPodGFnysrTrLv2FKwUBjHdOq1qWE4KrE61OG7s
T262ofv4j/DohUuOewUwBr8qHnt28hnzJbsxv1HLfRftZMLezJloYdBCBMyjUKfG
fFF7fGMPD46ru8rBnAL/egr8odc5EV0ElJi2NrpcRXhYO/Zvv6KXFMhFqbFgkN02
sdANq3D7pc6FzNU0XENhyDai3zU9Z/XVuvBOBdf4xIzAjcXyRnHMTS0+0hx+SuNW
3EqM7oHhCKnqQKVAPc1GLkb24J9inttJ6k2D2dtd5vDSkfwPQPTI06uMaTf9R0uL
Ohc6alf80WIcRG74DvzwuU0rdH48Ilk9ytKRlzP4t2+qLtWBO3kJsHqMN0tfJNlb
55ItBB8BT/8ydvy6opRIXnCtKcUYkwqM/RveDesn65PI+c3dS/e3VJjF3ILTFtMj
ppvTcCoWvmXy8hKcARcfFloOtFBa1kAzN93wHH9jAw/Rr6h3BctDnd4fxxYyxfCM
pO2xAK/mFL7DSDASU+00XlkwYtaxJdUlvZot4Wrks8a86jhIbYj1q93eJjtEMHq9
yRVjlY8eBcNge7a5nuNS+tQyVpoOozHyH7MifYcxzLLwiRefcHr7vco/83OlOQZM
OCe7IeA0iPjr1FDZA6AtC2qeaQHBEUIJsYScW5CtJchEO+zckar5Y+ClwNHxBIGb
dMmiXgIXywiRWTwEVGtaKlEdSZCgsnx+NOhfJYwcOOQiBSR8gyrA5XeElrl/XnA3
5K7uW8GXGHzRNi6Embvxc5brj+VN/dIm0eFA9AtVPXIitK9B5tDphZWNEt7i1u7C
OmHec4GEcFJ7ZcYdcrBTN3nZZi3CknX+u6fmGOOTC2ld1GwD7fXScjk8n3L3vPF9
upTQRg7GZU527UiJZIPz2XPDMN3dk95cF0ydKq8bkU49aZqF7iXLibwutaZOHYtv
lwqK8J/k2+cyJgrFLUCbRPsx9p0Kt+DIlkSHW4kYbOO+G7TKWTVZW/j2lqRmUwAE
L1Gyy5ks4yvPbX1bgDdHQHykgjDSnW94VogiB3nlTougIoEfisYJ5bh6PVa8HQNS
g+/CnSGYyh1/5zb534hCz3cVzpRL+WKRd+vzB503vouOqMOw3IsENgj7lrYqQIRp
CFY79IxNfriqi4tSzzR/9HIvLuYiaDabw/6JJppD7nM4wKUK0lWDe4OFMhNpVFYV
W0gOk+uFvRwBGdUXbiiSb2qevhF6vOvytUBYNpvekRWFtSR5zcPsJgWBMUvxT2Rm
1lbEPG5cnKaBDZdyK9fniTXbWRTYYI5O4+f9I5ZeGerVF1uZKzTDPv3lBfvY4rPY
WfHMfCHxAffFKWrZtZ+hsD8WnEyYECK9b0bxuiCIW1c+uPz3rwX2jZk1YXwegK2l
5hZ0UtK9swLKHPUR9XbDWJzP38mTLxvSGp0vDEY3koApjGVGp0bk6yCeW1kfDH+j
z7z+VD/5xW8zRiEa0zPH39AJU/CtG6IreCut/Ap7rvk6H5U9NWn6j4pB187uqfGv
heKV4WMAZ+AfS3XLw+1LiuES0lIhAoF1eFn16EkEScS3OA8Evz3UL39AkjzCTK4U
hikvRraMvtIR3DYLxo86GRI2hplDtEnZBa70frj3Fd8CGKCJLhT4Zo6cNAqNu4vR
NIsJ6z3Hz3wV+f/ZpbstOZVGKYhXFScN+M9MxJm4TuyFnwQps5N5sxhH4iX4wP2b
uoc0EkXqkLAdC6tzU58hporAwO23oh4U3U1BlSq6gCUx0qbZvtN5LfSHL4g5UZBM
ni5hP74AXmzEGslO4S1msiqrwRgGOC8olPhOESam2s8fm9Z5qIZ/SG+AyDHxIdtT
/9kqpUxfVAaPyt59xjqTE9adEmst7RFcwHBK8sCK3aw/eO+vHhi4kPEIQNgbQnpR
kSgVu4Kur4OscIfIT5qXihc0uIAs09QaNNjPLMXV4uSzP812hI9dXePmp1UzWVGD
9Dg8wbpyZ9q7MbM8xrJOV5auhQiKK1XhmagWJhfiF71Ty5T76lpo+8NHWvwzW7Tx
dTUxCD1kgWGWSbuwPJ5ibQluh5z9BVnGyZGYuznGYyD+ncYNQ96miskPIyvRBdgr
aZT1lQqUbGQKdKRqgmgQL03+IFRuIV8Hezp6QOpFObQ/q7smE0slnn/vyntV6yWK
LeGOoS6Q31XRn5tjdGQhPLZuFN9ttqnLjrvkmkcW63D4XU8S8Ig6emB9FIzGuZMQ
0FZZsYa8Zbtvo/64gUjxx+LMbyY7qDHofld7Y3+6VIPT2JDQSutlfuw0MIQ4SFJ8
pwCaaLQWRT+faBXkGPv/zJfbJ9dpJrGuz+65EzP0WdfDn588KKp34Errlu74IBaH
voYZAFw+pRS3u3CZh1TsjXRe+g45Wit+oRsyQyitUquFYd9ChIMjovFTeYWfGQYh
AODXjAl+NqCqJEdT+CU4LI/MBhj4kwkquPuWFO3rywlMlqyMBtRLWcIBm8xfusFz
3FGg5g+o8LeG7dtkUnoBypIu7OjjBFuw8exkaDMAMp5szcop1B5sZTgD7Lheebhr
ZUmw9HwsK52sI3RCc8JiTQPw0tTWEyGn+xwGpyz4q0ghQwO/Nxy3xUhI+GNaLahg
b3tiAYKlM4DsVR+vuf7w71UweM3DeE51kBC2tmKH62lr8LkICG7G5qvAw01U0Y6J
0MCEjSlcpisI8QCtjsv4H2j6i07l2v01sjWeosQs+CGuyzFQ3zLuhk2/n6o3RG5Y
VgGHAfWxDgm2PbBBEk6VgLgA40rKCt3ESGcOGGXZ5zGqSn40ALRJA2DoSghGr5aM
L41hhszU98lJIBke9dH6MgFqplR974QieaRj3fXBbrrTjX6aXTAdVTk71PNcDb1x
Dp+E+qJFsS8RsCvnKcZoMOvsZj/S82laGZ61nRN0ajAUBUwW6drOlY2W3NSt+ONw
mdbfTU03D6SnO+w9LnIOd/aMhuljjxD3e7cTfaVwrMfEbrIfBop9cOyYI3CQ+W/J
SyLdli6kX2Coc3YbXCxtfs0fEG3pf5pNtSKO4mi5r6Bp//U9y8Pw6PZWB7XY02tP
isQRvOE0C/qR9yFSymSY42O8S+2+wjfsg8yhniXcD0sm3c4d9VPA7FfgtLfsSil9
ObVfD5++8cbQu9Z1eHXKQ65DikR0puSUCFktBC8VCE4BBo1Tp5UEirGfXQFBcItA
ffHjMLtyyn6/gEng0mhvs/PXGNXKYQt210DruFtPuY+ShclXKPpIb+JyB5eimLbh
aAucoy4EaGzKIJ054r+Vj4c6DnPRZqJAd7f6zJSBnqmKtCeKofEcayADrfyd8O40
hIu5eYlR7vmkLHwEIsUnGoQ50iPL2vLvlYhDZItjebe2FQ/XimBQ1i7PYDpLlocJ
sqw5/aDW+IpONzN5IIRp0s4XUQQeVwk1/oIdwckd/gO+rqYKCnAMnDQhFWwZdZ9m
LO/ClT6YJtRA8pa7hs1l3N5GqA3wLaJG9Mm3EI0nxDZxbhPyEKhnqjcsSKXZu+7I
d1nP0adsKFEwxHM5q8CppZEjQ/ufoeCrv0iaoqa3HsIfukmD4yZW/HObBZZCuM4j
DtQNmXCTD8xgxR/QOkeE6RWDVunhoQuGVKVhwSvAYANCDIMThiP7ML8kCwoF5lcI
ML8370/G9OBDfQr2L9zlaKvr/5IeFKZb5YxgwYkOGoX43McdqbZlWcCDFgv/1fHV
HhM9XuvLCfoiy0QZgZOd+lA2a1oc3NPewqYRFpWYAVjCpYzvZlw7aRTuy6S6zaT2
rS9lgcBrWJWAqLhmayx174P1AeE/BFq4Q4uXgmVh3doIk4BrpJWGHyd1PXOQKcH+
VUisiSFp8xrI2gDCiSduxQoGftlYEMiXLvn7YWZIVPlfaZ3OU6HVzykqsXAsKCR+
I6CvZSHVrm7KL9ZomY+AbRB1g4MbPdqDpy4DCJ4w85XnF6ACL2CD5BYkhEQrKnVN
R6wZOSagbyiDFWg/a8Jr6BWxxw0GeDPJhF/ZlZyQu0gxGVio/uYRKCvwdt2qJbgz
VFL9qiqbNdol6/OBUW52Vh5315d9xmEF+zDQJx/m52cZbmCAw/WnTiswFjS6mQ88
TEKW+KDOfK73fCTwMrw6xKEbE5hHSnpjU1K8dFDqGIe4LXF4MRTeHSA71X+slhGR
NRr6wKAgyEQe2lbzUJiL3tkhleDWkEHDYKD+5pbFHlN5OWLp0c2SbkSoV+3RVY5E
qMUX6VBVeA7dbP1lJWBENcMKOUl5qDp1I6rrGEI1bobNIrt5GhyOekxuhIHK5k9c
BaotuEzIFNVn4/BtMB87C23MOp/Qw1Y0hZ3tiKiuTTUhrRZqGHo+WLGKya/XgOS7
qjN26vs8pcAQ80TJyK6UchVxrgv0NbxuzTyLtf1hKeW6QTen3xmYvacPWr15IAqj
PasKZYxDsWRpjLPJzhK70kzUxEQQEIRSZ9rd65IBLyp8Kjv2NvmX7Mn0elNIgYEH
e9tyiVhftH0Nep29yrJeJuUIzqVdq+cUzeRwpiBc1+3TcxKELUY+kCrDO4dLbasC
X61Bb43MGD14aNnMYwZNz5z6CFbA8cLesUpbO4A750h1aEcaSmocz9o+Yu0skMPc
XwIorm7LW/Gzk90q+eyb7SPGQHxNBCtCUK7KeaP3j+x2VFmW4MocUrMx+g1qQAdx
KDkfFbHtdPosIUU8uS1RaLWj0CjcuqMEQ0ZOynEqAr6spgGqiSdASobt/l5sYGL6
L1e7NsYk0yHRQ2w9NEoTU38GL5wmKhEf8P0+6V3qDVNUoby2UNSTDwsDCDR40inS
IhAGbogLPjAlzOVE9KK0tDRxR54LGTwrDjmnu4RU2nfWgd41abxEv5fomjFa665s
/4us6+xWekx/OY8bVCEa3Nx0PgkQnApzsRUykOywXnldXJhhntRam7DEo+RV+PE9
B/FhnSZzkW3L2/rNnBxuzE2VN26l7vvXW9jZrxF7TRP8jG4dxgi4v+4NRtEixShV
1yYRkYhujXRSF0z/yz7Xbrcr1l/xUkmVcqGK1RtEOhWt7iopmpbP/ZUDdZxlUwsy
phz5pFF/v1jROtM6nDVdTtOqaEoRL2DMikui4Nmd7CtQGo9m3JtSlL46nzmYj8mM
uo2PPU1MnMvBflDG8YBqcDqKRn/g+B+LUBg5F23r6J6w1oOxr3dRtYrPgaWAio0K
/6WDLZuDkGpZMfELlNvHTLXba6hrz9FR9jpA3KBc2nOoWGM7S1lisyw5D7wEZ1yK
GQWHMxRYC4eS0RnwyY3F8ZzexgRIg3ziOYgdd0LypD72RKQSGXQPEHjPkYLBErz8
gvs6jjSVTT6mujwSTp3o0pfucZeP9YNZhugZhwG07iRmfkuNnzHh1SdFwCLronrn
n+nSi68bJLKY7qjNeEiP/h/ub2uhJy4uaOXTno5yfTsxNqjOxxRLOfQ56K4lHivd
mrOqdR/0Hhtc3hr/L6rt1e5aweIi3tfpi3agFUKtGI7P7HYoZRJGEMneB1v/aVDH
5Yr2wElQKa2RQo1+P/Gv6pFX8eEPhUQexZxK0kSuSEoUZ8Dy+lXaC0JM4/jYOrnn
Rl1G+5xrm2WkdB5r0Cs7WYzQ9cHT/Rjew8Rffq0nVCi3ZdJH08jVCXu7C28FV2PF
DWcCVCc7fk8sZeM1XqCD6V5tA56RZOesXZ1fpXlPOH90zja72BTpAQrdvxY/nn1f
S0YpdWR2GnB2Pc8RL565FSSsK/rhXcbxMbF4HjQ50sz/PyuIylLQ9D3CcJO/M0X0
3RHKfp05ulBN0ug22N+WAXVyRxIIjd7Xx6sUSIQU0Ioz0chFz4xyQnJEPR4scrTS
9YqF4lRQJ1ne4mXcrmEKyylm6YVPRN+1DbhElRaYZKHA87nTIssKyjR8bi6D6KIB
FLnyXIIoDWR5qSUHMVC5ti4GgCb01v3MpGfeBqV8fTmoq3929Rf0tHtWuu/whUCV
Q/08le2ICYkh0g7ezuo6N0xdPH6NLo3vDiPpD0PxVQwsOGR82Dc0TI4aFQjChKoa
rZwumGvZ434pGBrX6cTEb/EBuCSvgkz6hJ3BaWIqDpuMjdjle7EF9Ycl8QawUB8X
p1JHd86TrNa9xKiz+0iluQe+QVGeLpSvtW776C++bloa/rpVbnY78yBXtJsGcBqC
ZEHh56E+L3xUCYeoQWgIpHvl3PNGv3zrT3NJEB7P2Ko3B6L44aqj2CFoY1hdDsXY
P1tDmlZMwWXoyqTXO7/dHUD6Fynxby0Qj5ZJwTjJpspCmmKl+WJX0D1cNFue2ERd
W/nvJdoCXY+FXoywZ3PsKkH/JgJRPUNeK0sAgJK/klo+DqJP302MIJfKORhpppEf
oZGUv25v/EvX2LilD9Tbq34cArk5NkUrkSn95W4J9q30E5B84YsSmLDctBKQMdZG
J+N3B6xEY7CbCO9gNjwVQLMgzSi+UG9+omUEgN2plb+HEAaOAJ/w1ugJYo0mIjZd
JEoh3yhIeAq//h2NA/hsVZpcZprYCQhqArJYg0SXi5LFf0HYQZ2lwciiaR1zW6kq
ZfBgV4P6Jxuumlc3rr4tZHrZDQE0JNvioKBoiyVhqi+P8BiQHIg+4jxFyiPXT3I9
c19LIamxapxYpGMkSqxMotQo2eM6AKIs3ha8/gNwEqz9XernhBSVbcjyA31sU5Yd
hePXjqQQbP7pV1RihNazm7WyR/XJrgAOhZDppozgaE5Yju6TnPFYbaeZav5vRTpC
GR10EuoDub75JUhbW9Mgyh3jt33ffGYsg+yBixiexsE=
`protect END_PROTECTED
