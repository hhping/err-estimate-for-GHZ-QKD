`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sEt5b50ijZTPX5uP8L2+KlbSj3y5D8jwUIjQtWPb5LCioXV/AImVQ+qQ0j8Fc/KM
hg0RtegYhReZjA5yCT3clm2kDPlj+51fAenkcXnht54pMPao9cT5TQT+rVQWOdjk
W/3A7pF4OkY+XsGTebHwsiHnDHGPzPAGqiBv2vujEU3M7bnWWr50wOC8IdaHwH1t
v0R54iB4HKEOvA6vKBnK2sU50R25mHZvqOlbNGoISebA6SnZjRQZZlTV2BgFVrnz
4YzbQNrl5qQ5zkUcnhVonLPcw7ZO8Sobqd2PkPIbL2EgFHA+q/12wvBkBFaRQLb+
9YE0cn7G7XV4b+/E9NwkIEP6nuiDEwuVY2VXPVX6nRYYs/gzkInXwlxzT2zNvNpv
UwoK5qi2N3p8OwW4NG0oaZcTz/XIsuDWcpJO6fchmQ5MQqS4P052OpGbzITuZOq1
/YJLww1d0u0eijcTSm0kM/lMMXLbXlpdV8qmqPOgcX1cqinVFsEiZ8RzJK3CKGCk
QBU5leM/AUF0d79CXQ+yws03bS0A8inK45xPYWRtRY3R+4KvjCvf7csMuarsA5Kh
J5KGgO3OZ5JKT+sQl4HEol9OD+7SB2fscKnVEAYyOC5zuZmiJ1M1VAa8rGzrWk2x
Dyly4fR2qMI06ind2ofdr9GOcuN6tAZLNLar6kyfQDLHALFXIyLeSsWYAMA9OydH
uIUcT9HHryZJgd5/j9J0Enp+kGjZmm0pimB8VfvmFU8VrJ+REJxPrwX89jYuRqYd
XyBxc7s3lnElaL4Y9RrTe1+1XNtsoS0TYYy2DlgOUEFLvhKBnOHQk+jxr7DMmBn4
IMcxgh21AXOBUSOH8ko5fKC6KsAhgVsXyW3xT2fvaqz7TDJIAhklMZ8mqrPGgM5A
UM80Kxo5w8jM1ZBjM5OR/TMR6BsAwMAG61Vxom6w10YlDUeDeV3kGy04h+HBV2Sr
YZYgj/WIulZV94iNPyGVN9SnQN2OOYaWUf1K9a1+BP/97YwctStsiC2zX9S+ObVz
Ggr3VuaabLo3mGG1K1/QKBmZ9y8qHEV8iVHa8JdAJV2eO8StzX2oqfFCZ0KBqFLh
`protect END_PROTECTED
