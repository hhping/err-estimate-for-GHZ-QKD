`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nta7MVN1Dx/6jCI0yEHbMb75GgDDTaP1Z6veFPQiEJ7+yw3HmdeCGrMdXDUkNTk0
QgTQvjNR10O/qeGSzMjGKMWGcN1n7M6ESaTD5NGdt6Gas5dwqek1VQ+x9yGCfis7
dsPuz7w1UPO3mxA4t9AVVaeaNsQbMhYAS8ZTHawbWLLG2x1N/A1Z6Zi7G7zQiIBF
I+P7aP6zZrtdN51YikEiq0aTBr1XD9nA0OavteVUM7NK+M9v9sN7Eq8bqXRUmUKs
Xt5AGfMDzYQLfI91Nnqb+eNvgs7cNllfhlo85ojU07Phwp+Wonz3Qnr4iB7u1DtD
zicbzieyCRl1MfuPUYDb1C1hMp8/p68e6jrZBCMBE6GJNo8mhYI7FOAoyDkpucsy
tKFBC1sKJHHwL+RYOi3hzp6xbAAYEfSOR14JZgiEsRa6R1KZgZXK1wmT5s3RTfqd
psGyVJdBeKU3n3NimuT16sn/+jgeQR8ZVxVqJrKIJvEP+Z3/66L5aD2wAR6efJnS
jqNkSHQy6rg7wHPgr0FHo4LLXBRmFoMAhtZ2AWAH0ApTfaNIvSCv9xto3XMYJVMF
wszHc5GIwVh9NgQOX/8UyM8bINklEtwXC45hWC7cPj1u1UYaoQmpBBPqFvIRe1H2
/ZpjCmOhRdG9O3ocozDpUhBYbHXW/dcQBWY3r2Jy8jkFZjLTcMi2VH+tlZTXEenz
awVYpTbeo8bgWxUfQ0/8Fz9jCKAKp6GGQctltLgg+6vvaLHQrupo4xqmGJDKeAm8
b+n8J1fHWi0LgJuKaxyDaJvKGrt9bYO8ELWf1mSkEy98b4IByOspWvgkOKhT86ER
TYRyRQ2d7Q5sBu8xkQsNy11tIo1IyNDDt3VcOh1rrOLZPUcL4IiAMW9RV+CwqMx0
kv/PCbTNdhAKw37SC3NmB5iSfIKpIWw1VKb5/bhKrdWYpa4+ZKAO5wNrLkhBJSNR
66AyZsUN/kjCL9JrHLd4EjBNu8yNQTuOCo1M/8hdZ0YbO/XpSvTnXitzhyVaeP35
5cCTBoGIOBlYFMb9/rwYpl9ToUAc73cLAZBGVqGxxUEHhkJqgf1zojt7PUA4RWvl
pVEs/JfHwE54s2vVVUbHbS/fEu71FNFN46RqDuFZhKJIk9m/aspUQ9UC7+3lEQAd
o7xS4il+ZMVUQqYR7ZOYEkY1zqsuBQrxwufmxbNafAfriFu5FUZQGhUcwbnIo168
dx53HtgX7QYsXbtc+hELwk2szkQjxXQ4dRhP7CUvpuVibpKpF6Tb5TEUjsQlqAGq
m86fHZ7mb45KuzgvyxN+EJ7hojWx+Hj/7E8qw+sNxutS67pITUIDc5mCKKUjcAVr
z+w9yMm9ilRpFrzvfztwhgGideoR8ZrFE+i5sBaVLjIk2paVtd8199t9yHnoAiNS
HvgmoJC6U2lEOaXIXUE3q5++0NXnQY+NhiWy5FUzgw5tfp/etOcD1kUAZ91muQoT
5MHUK8dzC1/7pYPBAZ+lYcLBvaPccaUAWv0nTNvxJakr+rrdm5zYKx/t5i7t1Ts9
LNIlzY/xfs2ehBP+CB+9NLv3trC/s74sHFgVX6CrWDNzneaJdJxyDGKsDRoItFPs
/hl7orplYL/KBP4nalKwaFoZrX3+91q2sliLc16/e8LAMU0lwyLQ7KMyq52JPsIj
Z38wZ1coNn5JyfoWlcVuvDCEWPXKo+i3lg2E4GP/qRAI0qe+EZlSXYKlipmqanoo
9IpIQRm9VYp97wtPsjO+6j/2WYvXnH0ZSC+ZL6zxWTwkFyQP4fGVf9hGZKVnR6lS
BKtF+JAXPIMYmf483CU4e8wazs55aC67JUi/Y4kzbGOKqHY1516nucOfM1/etjxY
FGWdHDBMlwkysJ5WH2uVrwhl7WrWb4IHMDgVc35foFvoT6UNXK95sozT6Y8jXHiL
BPcb2/hqkJQAjuc1NggqKxBTm18Qa4TQMOW8qK9oxn1n4lfGX8HIKMAwcjpMFu5W
Jh8NlGOZOwG6oUv3hbjftsv0CNKnpL5D1IDp7TdOoRTL0CwdQIKf3rTB7BSfn+M1
7rZKkMW1Vb0MqeBpM2Y1d8KC0fhyGAkhDL90E4RIE1nGTRVXo+g0vxzos8R7Lar8
KMYGgINdLbs679toDICibcu2TTayFl2jL8JAfdiI3hsOv7jOc9To9IgthTVyxfPG
l4AdpRXUTcjbMd8F7Ol6WobPHgl/wP7hhGnLAcL535TSDrr27kqEcBXXe0LqalcD
Rz1XKc2CKeXQ0WKlCewL8WNRNttolgGe62ayMGRtuRw3Xc0Ylx1/GGpqnLXN86n/
5L353b/EEzd50+VOW8Q7PhP1rT8y6rzjJQDTBCya7zveUOAZOXKVVMwAkMOyyCzZ
NSisTDnq7qdsNYUp9rasZqTY4PR/YmQer6Yzsd0HS1e+PutZBT/I9eJZhjS8Z0xZ
NpNQHRK4RZASIQJ60TJiuvsdAOBWLjA6t9DvtC2boR7pOK0eq6u2i7hx85H68/Nb
/UwLRd9HxEFqFv2c0xqCWlxN/dZG689QDp0qRFCoB5SfjJ654tw46/jcVpi41ykW
OiddLf7vRqP0nR29dGs4r+wJOSniL7FwXrtkbSpq27+UJMEtsdIwz7eWsG1cN+qw
`protect END_PROTECTED
