`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NZDo2VnjwImqLn3+5Yi6m1neEEomcxNxkuRQfbeV4Afn2bWjYK2vJwRfJSVOTGoj
3So1QIopuOR2G9gle8WjHwmq7DiCbyzEpDp6MUOfsyJ34Db89M11YRhC5htgvvbH
3CJgIOtIvwYRIkmXRk/0T90DR1QUcuH8QuBdq+P24becv3bR5ePIzFVZLmBnoiPz
wCPdONzidJQla9+gd/6g8CB/FfivD3SlvdXqGYWnybA6nVfPK5xvc+VeuenD+w1q
lcjki80vEXvHhBpjrE0V7ZCe+XJWGm+8CBT9EHTNEIet7JstnMrWga+NDywbK3I3
wG/ugs2s3inJwgAiFT85Bre/h1ADMvtnZZPv/mA4DVGELx4JefEeAXkyLv+LgO4n
hAPvPc4IU+w1UpaFUX//Wrp52/Lo5nmAv+EK6GBx7LesrKr028/pah5Vfkt/f/nl
XMZBDtuCk8vFNQ+A3QiS7xsEiSMEr2YO32etN+VNWIvalCnjAWnsafeNUF89ys4Q
N6MLFjBHMK3/A/uAB1C8Q2O4YlzAEVb247QNy34JE/vKDXekATf1vnTVUIbgyGKh
Nw/rMpUe5bN+CgygToCizr+lSGQCoPtr91ApNdsIIE818S/r4QQz88OoHpIQA8Bq
B7JG2LtGEAI+V6kdq5Pq6mrrNoGLlFbS3IffVSkIHnUAJOUkgHElSCaFeTPJ/hVm
jDGIqD/uuHxVO4MjKHuD9FqkMxFnAYi9AZb9J/RFPbIPs1TKkbnl1uifYHhFEe/n
SySwxhhIslq80e+OfCK9LdiopdQaDKO7Sq+8TgUojIjEgVNa+T2TkhVBDATqJ2ln
XlBhWs7QwpQGLslXPj+teaSxIyn8nX3c0AdnCNCkvL/XD6OKhNfQH2+VNJMSLvJ+
HOpIzO/xFfbZefvXXMOv80bE0aO6cz7wzzvuzDZF2ndSJ0WnCxtT9JpRjYRtLxh2
omoQh6zEtbSdh3+WIXCsYkHSIAxiN9tzOM+nOuLp0NUHlDRm1fQUaY3dgbV2RFqi
DMOQDbI+TTCMtvJmUleJz6VhQniWSTm4Y6Uy1HBulz6jq88KOvUJr+9sMmIxcgm2
J7p6QJZgZ0a5+3I96EyBi7wZV313Bgh9vNUmhx96srG+FJ0+CnmulzkpC/xB6/t3
K5rF/XRZdR5f9ht46pZ9dNy+xzBYgWctj5EGV/2AAH7729pH2uNNpOuSWduw9HCD
IIKFzqm21QFlIu1MYWvQAAALGjTBpwUViv7aL3f5YZU2NyNENWVmpYITBqY8mhsS
clurO1az5Ft7rx8bIxtAiIDDn4JlYSKX2RbUol0eGp5jSA59IZj6XohaUtIQai5i
pedSsFl7mmTgGLaShqPl2Dz/Qy8fzzXaKZyNJWSD5N7hV8FjzSuYdbADdjr9DyBP
oirZ4hetUkRjsA8pcXMNBqeATUkYb0m7Y4pNEYLi8sI=
`protect END_PROTECTED
