`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3iyZ1Og38qZBJP2Sbtl0L/tYLVSl6xIrnqrSRXJCD56TZwm/v1DfdJvsc+hSY3/c
CnvDpaU/8DPBWWNWM9gFKgCgJDaXhpbpYxwItrsA9ZirgsPIMc2kynOLCP5ec4/t
5TLTjfs4cWuHx9CoPP984rVKi43xKQ5sB1fG6GzRGOj2GZJeMBfGwnnGRXBtORDy
BNg6njbfyRCYERaCWq/3x2E7TeTGBx0a4aHgkmuhz/4WiUCPQNymOKnSkpJEfaHt
FmZpbIUZsx0Lv23RoZBsB8POHLglhlXVl1tG/IuComVlBcwLqoJpiWUcBsPBIFoV
UJ0KvgLh8obmuWbspOx86iIW6Q8SkAXQ/d49uZsii2oB+FDp0RTL8xFSv8VMEfpY
M6EBT4uajSp/8D36AOymMNldnZU7ZEBvmDwo8bCMkSFF9HOoCAbGPjQOj1m18PO5
PACfu9T73GL79nNGgTiwT3MHQxGBLkX74gOSYFNrYeIeRU4ujl3WSwNF0wgGwdHD
v8uCxBj9SuS8vK+h1y2t67vLa9NIaVTUJLLns5dkgSqkyZIEOEyBSbiGh4kguG3c
sN61eNiMA26kwuImaarcsTx0o4sYMdGppsyAcJnBxmToIwy8cKArxs7NikJfYBB6
2uacEh8UVI4lArR6w7NrR8ZZma3sMEk6CHLPgmLVsR/34QId8FjfAcJ8WgaSd4rd
GMIEgyvxh/ryY7pUNVdJy758KvNksqJnuZjFhqGe1A78Y73UuUBKBzjvwhzq894y
B315Emr75Hny1ZNAeMRl1c6ht/KM/eiGZaIEEpQ+2HVvXYdbOS3cSBSwRZQKxJ/c
oIVs+sqyObLvJwiSLaObcz61X/7L+YLB0fJfPBODtCZPXUKnfYfbFC22JBkbQVFu
o7Nwey1iQwLDR6Z71CvvG1zMQBLRO33w923wPiYfCY6xiy/6Ma58F3qykbFRnI6I
rJyhnfdY5FzF1O7IrvpqJ62BSKqsI9vTQkYK8nM7WSIZN84qY9xXbFhx4awFYYHX
ImDj1VmQRZa2lUOuY1sDHqVkys5sq0wdTU03pjhLZjlT4TByvJlyb7QM3O9hyQFp
Pks2d+SXAauH7Zpfjl2YFKtczz8tJ8oxroCbLEp2wopniAlyBxyeVAsNPkpgkAxI
YTrh6PMEci1icF76saMZ/fPvdxhhRZxzvrRBiZ+hXbqPq1rRjHW2TiUwDls6h+hq
J0YWVPuyY5Y+KsTEB6AFBfhhxLUvaSt2AmTawESuYT9OuF/KTF2QJer4qUtV3Fk+
AX7kmdNYu5a2Qb7oj3oUy7/nEw79XzoSlQ3kWMM1cLkMfX/WiH+ACK2CJ7xY2V6Y
dyfEe3/hOBknCXUAclCdnNWLHfLleREPueW8h97MODJaxxt+uZ98qdDf7sY3DaHa
M5+vs6D/6KyLcnH33FwzGVjjv9FL7W3ETXVSZIswhqoG45AgjzanXTZRFWRWAeQj
YXh8VPZIn7UFFYd5vTgrobls/jvs7+TYvUoBrDfRUt9E+AoZx4W+CWaQxkY/N8/N
5E7w0tpDtosZPhPmI5wKdBwCDdUUYT05pNzNg6X/BWt3Et49WdLWFs6ESzQiQfxU
HJRNbLBVgfpuPk7C3G2oTNdoXj8AJnAnqNQRwUgzK1I=
`protect END_PROTECTED
