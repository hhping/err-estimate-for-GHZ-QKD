`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wiwve2O277LfbfUyKoxOwgjpo8kboLUm9T5Rq7yBFHIHDdqyQ2/QT836EbuhHIxg
03dLpBencZF8pe4sFdB4vcuSvdu/5GVaCTlcEV/0MMe+jaAbmF5qWD7qx6T7tqTc
B7i6xcnrSSoGsIhGCUZuJZPg/fHCiV/HKOzRIKdQwu1a/ANWHc+C7zuWnVrs8l3z
6mxdXXB6giwHmsUVRt/Vw0xc0mv7U23UJ0XL/U7EihlaKc9reFNu8Qy6nBuwwuFZ
sRsgjcLa6o3388+s1vqHlumvCfakXY6vGcCId2zR1w+1WinsyiBtR0kUQkcHPYsB
obnqAWjRVX0T1fif5ASnyQMFg6ivc9j4ToE6zzjUolbysMvv6wZPYSHDiifJ6z8a
gqKjUYDaRzKm/5pklCL5Kpsf+B1RBUcPlhaTfRpzcnTiaqWz3sBVw71NML84F2I8
5XG5CB4a5qjD8XQ1AhkPKzwl/iyTv2CmvevcrmKWRnQo0ad7B8o9MZah/6mX3Af9
HfKt8x9PbdpkhhLFakySX3B1DwowMQyEOqwkbGb1YTRdP3czbld85ZYFwNQ2jmEr
hr8gae+Apq1DUKBHKzJlaTiKTL338hkrVvy0oLoewtfB/KbKudLDJ1eRDa5uaGIL
W0rJpMA4GI2sk58UkGzCG/653AZb79C5eBpoe1lM9SVEZKRHDyVyU+dpRvGsnaIj
w2P/EUighkuGJsHbCp1iMPyw2JhxclyhdVbpm/huiP437yQIcjkRVgB04d2lx+6C
D5iQF2PfI13KPyQmBy0SStcMnkFIXBl6HyxKkKfaiTyQ+wR4McLKRibAD5C8p6qa
pTWKpyjpa6YaV7LlnVLp05d6hLaDk8yWFhmxuApaP5TKYJ6r1UI2CbV+wkInItiu
pjPsecBDZydjJ2IQvXu++SiG6gLCBKE9eW+l2eNG89ziAyGVTQTQq/hHiT04ZuXF
QRP9bc2AYmY34w+fwnOyPHQB7xA6eFseoiqYV2JAU4D7wDGG9GfaThH9SWym2mEJ
GDMXiA2rHkMqheeltT2EEL+BrxWT/tRf9Hvb8gx09G9Ow4RRSVeAgGtAuH1LXriS
CUpLVZeFYt95zZJKgJ1W2BYRj+7X+jOt40NSGVuwahldv2+4M99eJ+EQLCiX9ESN
jhJ+gsFb494y1XK8ZUI+deRHK7oGsHtHY8MqMUJXA10dLlL/JiOHsEPPSx9GjgfX
tNQNm06LNVnBDTPzSqInmt/tnplsVWm0HGIXFh8Ax7QqnD68r/eSHB7hNFUYSi2s
SrRcpfSq8+3Brk5EKW4d+CKZhNwyK+e2cqACFAFGajLyHJqm24uOymFntWFbLHHB
/lUG7yI8GWWMwNlBet+9zFR2Ag/+4jZiDgdjt3AExS2QNFAputMD9HfWhXTdFx8/
gA23Jku+X/IMj36LuAmTD9b4ZVS1FA4NgRsRZ2fyf7PRn2P9qy0c4v/kFmT7rND0
wABECevNLFVCxaAz2fMGikqfechoipqQrEl3iZDgsx3tj7bojOEmqwX73j8Hu/Q/
WgwRGOLnZsO+9ChclQrTymCPnosVkNiKJsaTVljr78pBZjeG/6SRrwDj7eZ3ho9Z
/Jfud8iw2/DoE67xNBqMYsQF0mEghnZFoeJcMaNNbXhkOWV0UIBvg0oUNF0XmSOp
0I1iSyafBIVRCVIm4UlI/khhRsdR3B11LF667WhGhUlxzUMdW7c99REcS9uwwNUG
8zEhgwlHUT6drJ/aOi1fsVVSCsdJCtw0z4Wet2vH/3J8yma+x3xi261BmR5E1oJK
c8kAeQ7MsDn9rG+vmqzNArnlSNmnLwP2shfsBNQFdxyrGcpLOfYM09Q671HxNgSd
ruBD4ki7QAux2Ppo41kP2aklIq4mT2d/Qm2t/h8hN1wip/oLp4iQYGZ8puN0Gn4x
NXAJNIAZNPhpnO6Z5oYrLm9TRrJXOetL45jh9UqIrVMMxJXAq1GwF5PpE3GQTaK3
nvuPYOBpeNSuKdlwYaOjEDzXIMmrSAKITn/YFlSarvfF/4PBf0goF2uuVTsa9LU/
24t542vRBzJk2HCRJoCiJiaixwaObTLmWUExGGSt/lejf1voAbFlOZVfjy4eqMXg
gqMe8ibj+tto2odyhTyPKLTbeEDwFP8oWTaxFQ7ltReyT6rvuKflp7IqVY0hnMT+
Liz9SEzo6uPns7N7UU7fT/9RwnqHSrKxi5mEGaCJg39j9AKrcXRWypmEvwNGOO9D
Najhm52RjPqfH6OnMUIdVyi/2zsYR7pBPoAcLcKwm37e26vHT9qh4UjMUenLeozs
1namM4C/zr+u/KPfcAdb5boic4AN4oQSijE27191v15SnAhH+AhaYPK94LuwFrIT
yUpyz92XJawSzr5USns6rQLb/5RD6Bs2HHLefa5vWgN//hDk7TXBsaKDYu5g06gk
oMWeOKf+XFvFQ5yMVZesvtf88a0mqZOPC8NxKXeT53DUsYeB5s6IY5SYXqo/cL/Z
FLuwhT760fPwmtcOK2snMMJoBPDN0b5WjyQ+BvwbVwtNRBPlRp0vDtc+WR1mNKsN
5RK11KEukrstexpeBInyJhNlusbG9BnAKvVvdJ0eQy6Dt/5yZBDGbqKAJNFSYrKg
zhK+gf/MZe2jo6rJHpuWExYTwpqilAP/4xn6aCNqDnyx5m9GWgIuli/PNd8xiM81
RuKRbqlGWuCdWPzoRbmo/rVPR45xH2GiMXw13Y1trZSWkjhePkylsbSF+2YFK3XB
n33/Qjfyp4r2G9cRE/E43neYgm+k0b9ALhi4CtQ/NOihn04MxC1WAK45kXDoqFLb
px8mw+Uh1LOe4sGnLhTL8n0F88PutN0zwdRE+KysNiVwgzCuHJcacuqjcNedTCoO
VFDjGyfXqHpzq3ff2ezJUwpbQHoG6vtoaT658FFgnXK3xSnj2waYnvUJYSQ6RlKk
mMtxNXrzrYFCT/uSuAFN7tutXM9QX0Plxe7g7npw7THOC0TfyfhiBuIFRJPa+eJI
Af/TE24+rWxkyHvaINHsnO0UilZEYuTd7hcsSwaEYncjzEk1kdmRP4vf/g7w1+mr
r97AK/9mr42J7rnm675CUo3PI/ki3wKEevO1VTbccONSlxHOYAn8kjcT9F9L5DSq
I6G12rlyRNdGy7kCbTMR072DjFqTjcXN8CPIwtGuqc9IIVyvulw6uJ846wybr6i/
vyEflK6bQFenU9i8j+IpHoclNRdZiDfs3DAkkZ81Ew2uAa08WHNeesCH6VflD1G8
tPg161eACkXKzmKNwtUYCeU+YDKEKTgWBgBtx7DeNGTPXbYDa2uUfptl8RFBs3SJ
Q3gLde/G9kt9L8jrPt36W+/QFVG4AmSatL2Uda2IUEyNQku0aaLn9Lvif3FXuDeL
8PHvSDSDhmUZQPQ+lJOZcl8a6W81u+3JaZbdA7X1Et6lJKg5YSZ3kAxBqseBHMMJ
r8gVWOb4J7oOW0TzLke8yLdbhUaGgLSCEdI23fK5aLwsTaQXKUogExoZ0H7PzcLm
gjui0uJNYpYNW2OUStxnQsrzb2qp0PspCJwhVHm1UKxD0i1bQ1UeioYaPwCiKa9u
mTWOalB7ZIxmhm0WneqXMbtd0Z2EVDiR9YaZKGiDNIKXo0ILcjmZNP8nzqCHKaiu
h9161amoh2g0fWDgI/SQKjvZ6bzC/P1NjxxRxBUmnBnVtFh4AP22OUzJD41hsI9R
cEua/+MI1LkEOO7dNWFLfGu29xBb2Z8EJ/ak+iHUJwW+kA5XnpaLHEZrWFS0ioht
WMJNQGIVeB01lbJnAL6+5Wx6fZsVJw91suFGd7j2AHxJLuuE+26CaCBPUrcKutKp
Wym+Tfcevjj4BnRdQAT9reT37JBsEkaC/inlLQEPBcKqiBNFpUz1q3w3jqO31WtE
p750VvSVW/reIrKTk5ioP/1Im2jxRAaLKkyeiArJmJarQyAr5kPxPbKYmex4ys0o
AJIQnaV6M7uT84n9EZD5QfaBk8zg9dPEjkB6MnNnbjlmGuAYBqPAlJgX/UGAFVeJ
noOHMXXJQA8i4EYLcDIqexGuj1ps1y1eOYaq4oTrstfZgNu+ES4E+ovDr+5ZFxcN
iGxV9tpv3SJ9K1IWzAo7J82S3WgutCjxAKzEx7PoZvVcOltujOJkH43mbD3gr/id
I7RBz1zbrxIi1SOeVeXUVTduoNWACShuLRn1FIBbs3UCDPmJeMkFgeqKAAgB4z6L
EaI8DqSpGkqgjw6uHepS7s2jW4OPt5teOozQJEu2Dm1Xp/8Oy7MNzH5L237ZaqyK
jx6mKDS2hq+NQ0c4zF01V1HYWecKMZs2whzknFUa/q+rdRS17sltW7he20MSuOLr
fknLXps+r+kDhzXvtp4odk21BP5FG66JkVt2dNlwWPoKc9cRSBTZe17tVRlOZP7T
5S+OLkOa9mQT6dNMs/LOmmry4ERimEqvSGW39Xr6iEzYjDxHYnupgTq9onEGQXZI
DwpJ9fzETzzySJTKhAsOSWhcA6nfFiQ/DHsMVUkwTBT3AjYM/iu2BmgZRny+Fauf
FCxWTs0fvUosqQra2/uPDRRWwmFjl/ErBnRfMbm1OHq/+BrvS1coc9UvBZldg6Uo
I/aFb97vz1xvI7xI3PfsFyowIEdy4IzSxZ3PAIEskc2m3iraYKo6Fj3kCezOSImf
FD464IpgaOl56o2LoB7GPlz2aCcPCD1utSfPf3EmeKix0ynhYi+24RtWrSZyhCFW
Td2QkEIsLNDno+8CTxjU5wFN+nkFWEsxGvhE80F5fWnxOCxoYzoYERnrxrXqQPmp
gUPaKstJwTlB6Xa6Iazqz+IR2bV+xVJapbCHfVwGQCLZqJEd/5PSqXFe9dRxZGOw
bVG16/ntC5MOg9IEgHqcpigOqaoyHBEfvY+l7PAINCqOBTMsoSgrmmmSbXl33RnB
zVjDXUMNxK6VenVmaSRe1ummgoAOU4301Bc7dhzFkHRQ5HIH9qYc1tZHyy/4vYpt
c4AmC0N10siM5WELbNzW/kcw9MUFndGwFc8xymdecvyknFGt+TuvDnak0zxjqA40
wA+aBAAEYpwOwnmDFkrenXovBmZSlMCPqsjrqNzaspn4fwX6Ogf2GaNqeTpDuIrE
2ssT1mNnZiCH/KD5yz6ajJH/JnCif8//GtszYrRhEtC8c2tP49oE54gscD5qwo7H
GSjh0dgXvly6I1hHOOTH5rdA0bADjdMyFCsLREnglZGOA3xCTnk9xF3pwp4QJuE7
XfW1+EaRw0ZhM/GIqUlFLoNE8vvpIlla3FUSQhRB12OWTkHqhporOj35X+Tkw2Aa
OQ0AFAWUeTkLuGTL0Dj2NSwtm9crQCh5CiC4/Pi78lgcOL0eVc8XOeNwE8MMIxkv
s2CflOHGxzxAun1a3AxMGLbn/TNKq/Jq0hkDv9fGwcM7Wj0DodWZqDW5ciuhkGSu
hhYJTdo6cE5FHkGSfb+uu+clJtpGnNMpWHKg1qEsbTzZ+psOJSibkJvwU5CBDAus
/Ia/7/DSyRoZG26tR83BIVuI7wcP2SAilTWhIU4IlqKh4Pf71ck/sFux6wg1Pfh4
kUqbypnO8aZH9Xo4vDS4sXZq8Qc6/X0IqWwgOZ5uVU40/ZTXMp/Xh3jmRNUoDYmw
cEGfk38YUAWiDmkby3tcrF94uelEwsgg/Mko1dVcFxt92wx86ARKYNb5LGe8Rl7d
OYZ3UTI+40Rf5addw7inuO1dP0yk0zKC94VPNiH4Fj5KGBAibDdEYHgXM44uxvHc
HrK/9nIxfhZa6KOWK/3uJCv2V3PkHuXVobGSMWPLppRkvWYxDW648WFRCuNniJdp
MKJBq/ZSzH0tES6sBxi/mtAidFC+b45ww1WbTVyM8BH93Qsku++h4PUNtp6OHWVR
OM10FHISYzKM5GG8UveSxNBGsR7k6OSVKD/FP8uXvkKS/qbJm/XD/SL7Jr7LkzFg
CxQpkR1RxMab4yy4wgwZFevw/jiuYOTfWzzSXwiDVt5kh6nlFcq6n/5OuLghhNoy
Q/hKzevacAaYF4xzAD+/mnWkt2bMeTZidPLIMLUt6XekOvPSMhGN0I5ccRrnGKQ6
NmdKTjIFr0DuKbVA11b4pURZx7b+ITtrSgZv6orun/5mE4CV8ex58vHpC7ve69bb
eLXGTFFV/uWHCGiXREoyMMaJFFVW2qRby/7JtAw7c+lHv9f1OEnkKl98edlTXgHN
1K7h9YMFztR8UhM+cUsaDiA7vGuqCEwbo7n94YbOiCoFbigH3TtznzC/SdnFRDpM
FpFa2IWFsB4RmPudBQQp22ST86Mvf7ihZp7oaAdE8gzdvwOvT12CBfuShJmDFJMU
+TiONdhA+tXk96u4Oo7aqI7ltg72rHX9uHbtcNUN/zHVHXPDnKlUBcKBcc9ktU5E
qXkYV9DvS4LkIO8FiESRSzDuX92guFqkRpURST9V6sBF7lxzcEdZMp6bPg+r4D/u
geTWChgatE+DgPN5pEiXtU0wRK5bHUIq0bAwFA5/BEAT8yNAKlgQbwanVQ884rmn
OX8hpD66vj3QjLv43vuJotjYG8ZBlpoRIN/b/cxTLcEBrhwCldPTt4VuYMKkRs1z
ipXt/Hra+uY1mdrWsh7dhwwFxmgRISwF8f56QhTfWTo4XCECqg8qOtB42YajXxcu
OtFTfIANoRpd+2i+ZWSpFCNXRcym1yGZNdf79n5j09KNw2w296ulkrl+bQSuhfgJ
mpdH7u0UZQYXNuLnANn/derMR0wZJOjw86AAf5zxTaucnVXW/PiXYo7ZxtqTU/Ra
2pu7FRDBYNn+xtk7KRsk+g0q6ImSSV3UTqJmtL7LyK5oUg1Dwttjpixl8Rtq21DH
mkL2S2Qn71fFDeJQ0DACAsCIe67rNfGcKfwJIZhvyCCYKoiN94e236qFMKp+PPUb
GMNfurn94TtHT2CCv4f7J722E2obJ6m0yYDWCTuoUFGIkN5g7jgqaLFG1gXv2J9Q
DcpzEGTdorvjf8BdaF2TbWCsyadL+gnEKP065Y/E8A9/Xc6KtyuEKpSaBFUgYKx1
bxVr0uYJ9hrQIwb4U6pN39cbvBZl27vY/gF1yategi7BHFvByDxcES5fk9qZJmfw
wKfWSJZ9hahg7rWyRQX2GDGzWAxEiHurBzorqMf7dfx4Jl4rNvhV8MFxNB5B30mY
571bzUAYd+gptCr8u+3zZI8lbMwfRW7Tf+LjRlB9oxUj+wyaQxKajVbVGhMR0s6k
AfHyb+zUOTTJOpWiy5+XAmkrte4F3nI0pB6greGcGN/DgjAVpoe1aFBjstUCARyT
fpMuIgRb7Xg32saJ89hJeS53orx3JcYiCeQltMsBeBjGm76EM+BzXowkYO8ZpIBa
tqbeoSTr+T8S3m6UntXww7OnVzvc1EADc3BJHjagy7AEEe1HfEMqEKWbvzQCPIEv
E4Den5SYB9OQ1BQy1fED/NipSL5nD0UTvsUaOgNLKXBP0iPyxpLiSoXRlUlsgMyv
OphbM68Q0+6sRWhgdhV0knb0y6HPojczXGTEfaXHMkkxY3QXpATbJ56ZlYvN/IT9
dqP9SXcVU2Pth6pY7JCEjZNb6n5sgZ83NvbKkHO2fQ4/WGIaH83m5m+vSkrdftvV
wIrQ2zvbWcl8VvB175LsoY5lY7ai9cmtswNmtBOAuEeSWi/0O5N4UFHUmcd66b0x
wdkslZTQRuc4+usFm9vT3cx/cQQmqtXvDzJ1CfNxwomFpoOtnrTGJixG3KtHBsns
pGh/I59ApuESgjMMStQXKFBr4aTWmX5DaPLRfi0YjMmf1M1piEPbtbFhENuNOAoe
+rRvqY/6uvOSt20YBXCPH2WdvEmmlkqdVi2jqqdkKUrpGhF+g/nhDMIKB4x0vxLz
AGX3pdYe8kH5MlxBEqwTfUIVBrHQPwHI4sGYs5ZP0GRDJ3CDyMBj45bjbvmBqKd0
H7mbFuYaAaS5a2/aSc82saZG9ay+8GqJQIFD9EMDBXNX+yVMQdI9Z7PWFj+wwlAE
2bwsyKFaUb3cQKTazYdwvt25uG8XLr/XLA/ZKdr5IurA8h4LAXCEbgtxE2Ak6rAp
mKyBYK0TNeSFj3pghf/pKo2Vp7ddvdMkwXNjyU2duh3eMflj6kZcL0Bt2P/oc8r7
Og3K7466iiLOtz6fcwhEPdHB/DbuIXuLj05hYp4ZkwU1yj+YeOQp5+x3pe9Q1Ul5
6srKT1wBmmW0RO8+GCjneFYN8dkNnV4ZC10whJmI+2A0+lbfeg7LK+k3tlIPw3kG
fQpMFF0S7Cs8vCBIg0XDKls06i8GtGW6djpbCf+uoaJvA5EcLWbUSHhsAtU81loj
bn0dvHQGheydhDJlYd7V8A2mcyxIKYp3D4nH7EojUDeoHVy7TL0lDItSTwmbTWF1
HXV+gCSa8nxN+JFwm4jlxFNDn4gkoxGnXFxOtRhqp1oU3Wiqre45MNhcGNLH6hYi
3AMp+QkRHwz3jM1G8Xb8Bl/77OFaW3o6n24YoFWGqVE9wuLoZwRYIcY+qkqKpt8W
//oNJAnryfgA5LZ00phvq928y/OK7GPU5/1A/m8qIBvbnhrSaUMZB8VAI0NfsG7V
4EP5flyhbLHa0PJPOjIjR+w2LZOw9jGy2OK2rJn1HMqf+IGin0aVUxs5DQz6TiV+
VJBflOfq9EnX5cugqufp8VlAR+T0vvdcIWh9o5Yvgy44UUkv7NZlVb63tFphv2nu
aQuV9vzjtSp1Gvf59JVPOWVXWtVPA+ZMtBtmlhzwFq2GdJ1k1LT7qXmskZMsqyfV
VBz9Rbl7MoHfmMn98vuuqwcViqFMmbs2bLgClMjIDkL/tprqMKVGj7PJIPSqB2lp
kdd4YBLRyk+0LmA/7bY2uxGiQt4bZ9ZvtZ4xW5vAJ23KaoSqIiEgwsiiMHXBD6y8
WxtKsW8w9+IxMAbTtlgZn/5ZvnBvTBuZ6QXO55hhaVhv15XZ39ILsUwKMXxOdMcd
uqC1jaPgS1p3i9yeBaxwdk4fcMWOapW5QmR+3tw74SMyNaKSuMKB5HzBEdf0SO0K
Rn4kcVx5ADaRlZhBEdw0PIkqAHYhltF6JmTxpWX4MF0J41MBZrMIKb/MrFMqNd2r
XpNohtfzpSsCxgglSghd9byyXF3iZ58IShppdyga1l2KBgn7/YrAPi9VxXPOu8yc
q+0ZUn6NKchOc+vkeAwbiI5wORH7e8fQ8xLd/44wjpehcVdYXJVuBruMUWf4ohPL
fGg0OouO4iMMwTM0uuCZIOrJe3a18AjJWRhCVd5pn8b6QlxI+6tdIdAURNy7DzNv
ZZ8uZP1G10q7tCLqA9RowGTHch2+BR5KpNgAQaTBvKnPbIwXXqFzXifwcaJB3hNk
0MhnT0FO3l5FNBdYYOP8Wq7tCeA5NkWNFfICjlYzOHoPQa+od5EQ5ItheZcCWxn5
SS/wMvAEsfttmm/dKAEvyjN6RPP5FDmV5Hr0gYZkGQBM5z4RFdT6jErZFbRmQqcz
g2knbAg71GyejgwIyI2p+sTuqSN1xdxD+LEGy1vrTP35DUKdPm/ZJybQHxSWdnrd
aHZ1lkyrM0ha6n1yswBb+9Nfrr4K5IYofPMc3h7NzF06x0f6EaEGZuDzb1q2n9q7
J45b2qvm5oHZDsBS2QcY/dX6WvQ41HEX0B17KEcpsYxBtgkacpe70Bk3GkWR+7Fz
BIVCoof7m4Z4uX7SmRurylFcm+w6dIWOPYMtvaKZ86ujTWU+z8zA67BacdrOvKqS
WV6JtoRMU0NSBhYB9XH77ufDzRd2YFFdTOUsjSVg1yhVQ6t0OF7dGI7qqBJYKpAG
lhIHYmbTLCEk0tLu0vXXnYZiLQDNsDoJGj+MdapBWc30I9l+ddqV2lhoacFeUn4Y
TOY+ZktjxNsXdBwnkNmaoss1wwzbIQu45OHjCZVQtmYGrtlG6Ym4W9lYP/sF694g
qQCg92nQLJDbxPRRfUTMeejWaUPPLgUB/U13bbAXbo4P0pTahUlbmnwThFvvpP33
corfHuVKYi+FJq/AMEOS5AdEpMkLY5VMDsaoj664L9DZSno43gAwGncWxuQo2vVs
smcuArUZXEM3n6uFCHuHppL1cwtNVoHsgma9ulvNSgxKEghVcI8pEioz2N9LGtF3
v8vmc3UnBXY816+RU3/S/Ig1MERYai9JHPB45hXeZbPNPTuxDF5Beve36H3Hv5Jw
HZ+D3eDxEcuAxLGSVwFxl7ocrUWvznZyZhQ6f0q17KQ3XtV3UscKsGX6etsr+KgD
1R20MheYVCABSbz86vOLMIKquX3ga9s5mViz1FriXRxsm3PAQnSZpR0JWmf9/XDQ
Dqot+TDgYzHcz23FlOelEcbghOMZOgZWeKOG+YNLMHWn9SI6Py8WVF37izHKWitR
EQlLGn7WSwvq0GB3wAdWS7dRhqltTROe3zMH1eX/YXgDDvKUKuuAC17KJnigpIBl
C+VJddwSce5YXwIxmRpmlVH6OGWYZ8iS0zjYqZ5g3z05sFcWyHULawuzOaLBQbfc
fbJjVf4NtZKCJnlcEDpz/RhqFLvNhPPO6kQUnmSk/fdyHLggAC4BM74b8I3CdY/v
EbLh3JYK6SzyJiXSsXemxWcUxMFtmPwsaGGXYDwIpvxRBWosaVINf+N+p5yNKssP
zaKAwmCS/0sLGoKwNcy6t/bhnq/FB+Iy1l6d5hxzoICdraS2tzvvrCQcDGKjfJa+
nEMmdOofpSl6SsmKmxA+F0poQqb2mYqEllpLWE6Tn3QY/vveLEbwxrX30E3i1Fj9
GfglMDhLlbCCE4IGI1pLpt4e1vspjoldCLS+RsRubeThgvdEOBz8fg49/TSIyR8f
0L1NYH18Yur1bL5eqrA9NdqYY75LlWVIkx7TMCmvcnqKZqIKrxUHo/tLIPIWfNFQ
UNyu2c1v/oCoKKi2zXZM5uSLBueifhXpEc5KERZrQXs0wYxxFKP7vSkHn9Q3vc4P
QjJfQd95ZAhy6trq/uHAWr/O0cFxnfZYBnuTPHEdOiA3hPYoGeGtmD0nKMGfhAyc
/RaieEU9zIs0S5ikNuAuPYkKrVk7Mu4W//vdMjhHv8dQa6VCtCSHqwwomg6qiib0
M7ALxLAj9+RkE+HXy9IgmQ77x9HpZJRP7ijwhB1W2aMCvX1WDN97mMaLgyXob1aI
H4C3uWNr2HJuqJt5m+4LngF5U1zub7euoJu5iALxzAamBBAP9t0u0KnVWf2npUzO
1Q2+VTDRWXDvl8uuo7H1PGSbVRvDiOump+5+AlWaU32CsGgv8bP7LO6T8DLt7apn
fD5I0GlPpk294iEl38OPyu0MWPIO3dLE1pLg7Jbs6+gzGgg1E5OH93Yc6vrdbHuw
jOTSdNYuQmvwJTj/Ed+2JYO3w4vxFz5xj26DTRCQRJzEFrQy63O3j6BqbSbcxM6C
yfXs9pKWZiY/6jtY2rKUA1sjVYjlYaYIq2qPbDSV4dP2rfHz4mwqzMxgWkmk7x9d
cbkf+jzE729W1PCLXtxp2lVWHVP2J/oEXC6OhxWlqfuhSl8N6KaqjBsgLc4WZ7Ec
8oqiB6mDAWOCjgVq3foZPln8sjfsu1rQJhiMHP+x0jrb02ohGxPWGF35NxEo3M+Z
aNORMs1wPR/PV4RYcafQyzyhJw3jScf5070qSu4DxJ66rXYqItV7+hGI9/y6vAYe
GMZAHuLGV/ziDGewZ8h+q9XUPJUkprIRzG7awXyoaMpfZ1XvFwAncVTIcPJbQ70y
42+Zz1lDNdqh5PlAbEEEQLAbdOpAVatygu6ufvjxbj8atmU5yx8Ig+P6D2OhrkqH
Xkv1vn1bjG9Sz1iC5zgmiLySqt3M8h/WHjjgjzDhS8OTGTUbtmMGNTxUGN+x1UQU
tOIa4X64/7PRLv5kjIgsCjuGfREAQyLxDSPBkHK/6Zmx9EINWFhAdcTyI6PcnlEf
x+h9m4kBw0qz8dRuU2TCOuDZRaKFG93mdOb2DqSvxhjWI6E185JxGw345CmcOvgX
+uk7DIre8Val4YrqqMCs9aLyrLU17nuB5R96rnkPYVLyDtaHTjRUG37tXEy7i6J2
FRBXJPB7JOAa0Qm9zPwfq1QdAEXyYq3NhmIAjrih+28WyswU5gkBpJ9CaorYIr0G
r0eKVowLzP4cKZnobwxggJu3UBCQIxvoLg9JJkwiRpKaqBiaPee6c26IfdKE48Q1
7BcXyHrt8WLamRWUs21zQrKzkeKMSFc6S6MRg8X1zfTk0XoZ1115sN2nOt4NsG9n
mXtRDNY67VhE7lI7z2WqD5ImH0Tzt0jfvmpTuin1KKrj+1JXD8SqRN+L8eltCa19
Q8wZB3V8sJgVxIpYoE3oKvY/lse++oTiYg+KyOJSGEiUyhEpZLJyfzqf9FY6b0Cc
AktXgcph7191yhCJBEp5fKrTt0UDJyVwrSIoRgrTPkPTKbzUkZdM8NcVElkebFP/
mtR87sYekYPJUyLtikyAdjGm0j1A2e1Pq14NawoP8g4C0BMfAUZ6rXXlWbyDSQiY
Fih0LpegCzz1roIRc4e/cjr1G8yd4qAV3RzVHSewMmIoWUILDLmJPivTJTHWNmvy
tudtbZdj1kJ5E82JDecg8BRYxUoxKZhaGLCI1ibV7HFUdgJDV4D+bv7c+4c26UGY
0aPr5yzeQvPRHjTPElMIO8yBiUGnNb7IcU4KEFuZ8UAElrAGENtMErP0UzWIGBbk
MfpGIhxqTCEfWyW9hlxEK3zTDHolx8q5AYX6qVcthEGIyN6KY1kYcOWEOOSW3Mjk
r7nR404jjYiBCNl0v/8oHhskVDtbpO67hZ/IcPGY+EOtW21VZ0obd7cOib5EKjfL
5ldaeg0l/+FP6ZYGHKr6QJ3rmNx3ZULrE0RXicZPfVx0n8KQmoMHjbSyFze7/eSA
intICE6UkO7rOFWG0cuORq3cGrorItdEkyuJu1Zo66nhK3Ujp0pNrN9ZaD5K/fCW
tDYF+zQEtByMmN3XJal4tJGd3gtEyZO+SrCpKpU6DUboAIUNou6f/wSe3WRK5zsS
dZ7oln4n1JCUWdRS0I8LqfPfY6rY59Qge2wXNC1X7F4ykgGI2uUdjnroyrG++W1h
iQc9YMR+EmLNxfczIonACZfR8eFNTnFL7dpqTkGkKx9UPUEbKqFchJWPbZunPIll
4enu9l0Mz437UbAjKwyv3AR0W7YTHt11HFLMo4Nt3tunTShvWjChkcZjfHJrbfRF
OFMQ6MmrPPc+F4kxfWdjHKZIy59/oG6JvJ8PObySoDV619bjaig8VT/EfNC3G4OO
/fMfXMead7nVUu4ipjB7lEmoT4QjzkbpD04LSPMkWqZ0ywL8a3MBaOkD2GMUSNIF
X3aVsP7cLuHx6U5fhGDGcCe8uXl06StE1sWmIqkISxTtPulf0I+YHsj2YUXHHAVz
QBZRcy+l4wlT8UQsjVE0xGTaDJtLMYRTO2u/wMzqXEUIRWMFDiXTsp6M9u4A49+U
ckL76PUlFgPnyi5jq7Huv0a5cEItmWKlQQuzBiI2n5QxRVQGDPnKUoIaJyr2uXyb
6+HfUo8wFL0chsNSsrdw4la5nc30bfOx5krFPhUTOb89nb2L68SGjbFTQvI8jJO+
4tszHqFzf5/9d2fLQ6n57iYHvJxMZPL70RDivf9Yr2TD+we3/KpF73pKFtvnhQNQ
4R3KUCUDk1nKyYPWtksXLis5+JJAR+wwL5Ffp15icwy34ZVhqGahtrKHrq6T/nvM
J9bNUVIRGh65vMmFBdwF1320Sb9GPwK6M/SbofZgiizmPoBHcc3Uq4angPHASwT3
tSJDu5f4VzJNXt3gBgR1wS3/vcCaowc1r3dCFpONx7Dd8MNg2Ctf0DEc2/Xh3e2T
H2gwRkgao2pMXjiz7ndTxxVKXyLljRY7lJ86c3VGrFI9xUksCcha/KwVyIhGn14Q
3u7RnOqII/0Tj3I6GeAOXr0C3uT6dG64aOG0XH2PRqNUNOeyr4m3XNsgW36v6Hq2
1iMFY6g211wUlT7jtCZ8zCU+4a4GvV3LWb/AbZ1CAQSfPjpi4JTEBDBTRVmU08vp
gwQMlkllfVpucChAkCOPVrClLENGMOQHOHvRmVdlrCTvpNa82ErTQEKXiemeQUAZ
JftbKzFaQHuswT5UDYfAAFc3uM5MdIoWlqYlTLGsRTZ9C3ndbQJA54238zPrZxKP
wPMLpqF4kV0zKTLOvp69DAbiRi6n2WVuuXMqd7vSRhuqtVwBtiPEs6gjoEkO+Nkb
gKl0xFnqJ8BQaXNtgwG5zMEwCR3or7hYceOc7dTHSZrtoLHkvJ7SjZAjJo2m9gNP
KYWX7cgFQPesTQGjn2sWN8mlI5ywES/GGeHYoFCcYGhkZq+IgrPKBi4ubqOlklhf
ppF/J2D+9zzZjLnKRev4edHjeaBVljO4Pjwwr1dB+avsXvCExFiSNDg6PT/a270d
o1IRhi1Mlfze+twtv0YIDNiyr1wKSnY6n55r9d6pRO9NQH1GPvYI6KbkOqMsiFfy
YlTmxpRa0aT9N4RLGYfPNILeRMvx8iVzmmoHPPZtHKGT99I6ounBlrXTVJ1U2lbW
3wdXV47sCxxj1K/PXUADtkkSA09jYg/5dv0HGA4tw3rh5xFOIRTl927U0IxMJPir
jL+VaA6feIogGfg31gwC2Z3F1gta9tRRXKbKLdM0AnPIscN1kdWfN1tFsSIblGIS
VlaJ+nmTrHoXdqyTmbGgw27Ze1gNHhLCwh6wUu5UJ1ruo1owwAWLC/8iUW7iON0b
pUq+Cg7P3Dbi7vk3dU4eNYJgg5wROthe7mLwNAN3HAZ7lx+VqeiF0OsB4tCcT4tO
9UNGDD69RaTYIZr+ewHlr/sF8DHmYyoEPtzJp6e+x9KDO9RebS1hWrLNqXYHoh2Q
ysZ1vqm7wAVCESNsTgQS4jJUJbu8rQK3b8QBY5mTafOgLWz+EmApDkw72JYk5fC7
q+Z4LIfJ/gDgYBUyd8IOgeoT/rgCnZ/heHia9sQdl1fhMtRycZVwaO3STuw+b2de
FpN6C7Qez62sN143KddQk+cED+4RxkYgHPA4EIJiHRZR29R7UaAbQ2u/vfIMWSFf
EVSTEpW+Hzwl3mhPrBXwNk4UwkT/mtLUA083b7q+nH8lWhbnzFrtUBdpGKxKeaI+
Ahe1qFDa4tdtneNwMqYcJcDujcJIisE3Yp4Wxn2095WivteUvgZg9qAr1p7Y1SDm
cICAheCz9T5sBdE5U0bo6qT4sVXdR7Z8EANRtIzcRnSt6zdSVw0xAc4JzTN7vCMf
+escYhSGRXt2wGq92knd7P8Gytiuhdl8/sCySvLZj1XAF50GIpGX8fGfn/7gcqFl
8I7v5YknVDf8FxFypvkeKJSoZBXv3tXlIf+eRRz5dc38ma1pINXbxvG/BgMkOsCi
Uknomj940Fm9TwH4pF5FVX0jYGd5pkrABbsAR7ZHgTU9VIfK7BgUlnr7CT/nQl8+
EEQskvqr6Bg/KX9MR62DLOj0/q204lvmCX/60ABwQyamFTYFDxbB5ZdgSj4pL4MQ
aFjBT49+KLI76qa4rCXq7lvOLgLYSnOlvOgJFNNUKTr6lds+xzGNPEp1Tsmb00Sq
r2x5u9q2YjOd0gDDep8Pd17ds6y2Hhr7Wcpif5yyBJq3+Aub90ZFi9w/3M+77Ypr
aBhJPohqq+fXhL+ZXPY5G8pmC2gDhmFCPdlxeufOfRU5cfqK5ScsSQ2eXZguJzZS
8py1kcI+ir5qrKUMRUbUZs32WB0ptis5+ep6c5J1KJFN5UikVYBzsDnSh5GK64wH
GCIrl1K28Vv//4pzE1PiX1t/gbQZ2uSJgGVRpbp7sL5bvKKWFaXIMvu5jTeSGyFs
85mCzPbkZARg2wT9Z3e13yZ6PECleogoE7zgo7sKu/4EDAymOrG8N++Nwt53MpUk
B9bKA2FJ7IMfPXDqnqV29C2xyPRrarW3loVbw+0F8CdjT/eHPPQq4KncjjJlgQBE
Fc37d+ZjZkxCKLH0edpUkHs0BAKvTvUTwf/7z3NBr0ONyhNT8z1BPd5jRwKG9KL8
uBy8TTsA0y5AUc37Tb13W5kRH2OOR75IIdFbqeUoXOmOQvqu474BFZevYxoD2+NE
hvirzJIyQncF686Fteji1Qu0IJ0Gek0gpUsfZbnREt2P7IxZEsJRL+0OMM0nWRjy
KIqq/ejtME6A7xVj9nVc5sI5nBi0g3s+hHFhdpYxA/LYfv1Ef6Q7d+flVWnGFnsI
kgHlPwn+3fUtHWDDrqVhTZxC4ZjMFV/8msE0aiURv2OVjJDzyDlTmH2HkI/DvgtZ
/hFxWwuIoHEU0OtozUa9nEhtHIc1NmB5EAK0iziJk2KfPHxxzAiNFee5piTpyL+3
FFbzBvM8ZdWr+SpTpjCDQdZ+XaZvKQVxsNAHQKNU1KAST4W382Sdoumze5Nr1E37
v3Mvx/RoI7jjSg36KU+Olpl3eQwyQ+WGqVwpRJUv8Ghkh43DXkhOApWKv9nN99tb
/kSX69vPmoCOpIi9b8Te02NyIUlQImRATcBLYWZx28CwgxxLt+Pd1GzslfcZl59A
NBEfkqU22mIP0Vd291T2n8t9aKwqf09nt/RjLN1nCz0iF4RmhlutwslZVMwYSWVr
UrfqaolvF98w/W/wZVWbRTlSNpCVgj+q0sPsqDlbLlDsqpLiPx3X+zgX+GrSbHHb
rSTFr81Ep2bGtr3L10o9DK7xKjoXkJhVIfwT05wyg/QH3ipHBJi8TLU7fUDXTBhG
9aaKQQM/1J4QU2jx1qmPGcsGJf5QdijJc1P0Vc4Do4BrjEOPBvad6rOgS44H4kr2
4ti5Okbwf36mtMFLBsyUsXQAERuRKNTPA+n4GRoCMqDfWtn8Z4oSwk40hyX1HRmM
5TLo6I6jypW82tIRQOOUvpb6FFSvPiPkfZA3zKboKtfsIb/ClHfOYC0iEWN/qZkI
P9I7MT5aGRHJX9MVMr7IlWSnsZIowFLtb/aYdqymDlggWPO6xfejCiRGgv5wscg7
PQKAU76oL/ff1TSLoPv4vXnubxeY2QyAlA3errpuNnIt85ELR2TNhKnm/1K9eRkI
XY+7VpnB27Vi1ahothf7e4cdxXlknNIIWjnwcvImnXmg6LTvHTVztC+IJmhvKUj+
C7CUJY8YqbJdsX0cMRA1NV9/4QSud2uIZqsK6r0cQ2CUXfBFhuUztpeSagmkH5Lr
3DC/q6LRVJq0Q999c2lXRSx8ad9HjjlyCu2TMa+Mc94HdVolapf7URt123XszAF9
6NjZ7x0hKGZ/swJABgyP92/KYtaAJ6ehf7AtAsKwSxuXwSbLvSUc1wzH5b5TAC7Q
NbR/PpleDTUIYbMSZJxTFPKctx8GKH6xzd5P59AsEYYpcqgoHmSSumjpj26EMYWp
vnnYVqA3rPh1HO5erdn1efHCbNTRdyX8CXhpWAtbY17KJmfm0WXx1YiBjNgIC1Rb
Q9LZMmTXyqsmh2IDZcPEx/r/RzJB5LvOfYcvqXtwtNpdTQ3YGXC4JGz1FOq+VYwi
KDrk8Vva5GSzvbphC64N/2RsGuiimjh6wVRlPuNVE8DHUdXebxdMVEzT7UUalO2p
72aYfxjqYouPT6PC5zF/N2/Y/JQT7CsbK/uIfqsz/CKWVkgrSfnpdaHF04W1sDio
9FT42etvtlwkQkXP7cREIhBax9U2p+m6FjdcyOktJMqPJgLVoIoRWi0n4HhDm9ir
PNwEmqADN+E8KDT3aSZw64aTaon8JrBRmPNxnOmiSdKckbGe82g4cE1pV6wDgWMe
EVz2jPW1tvwnfGhpvpDvbthkugRhjwmwwHfEfGdxgig2+ArHqL+e01DUggypobhT
KQYu3HUARE+VuIkvnNyKnPVhLrzkz9uq0zaaT+lOuclyA0eMK5wVXLBDVoIAwfBB
8AtUfNT8a4s3sbiji+SJOrPkLSfl/OEeLmC2NJhxWp5EQF0GADVdFAGfkyXxhtH8
T6uzv24ywc6+ZqbNSVHNqqxWaI3X70TYUK0HJ2nIm+oy57akxAUuU9VGwDpfJIeG
q8lXL8AyRkpC5aCWnldyDpgMNn3XCF3VhvaQv4DAh4/NYti4+2tMcWmQfUs8E1ga
M+9bWRi8FO3zgnWbngKZhL+7WFTJ7qz1FsrGKwrZ+qErqwoC2pSLA0uxCWt+2G21
Z+EUU4CBh21dVE0KmIrK1C5rDJAvvKIoKvFLBhgUEc2QbZBYFs+J+z8oYF0I5zqp
TzI5N2yuQBdl6GR9QNTA61yfqoe0mHcy3DF0m7J59jjxTzTmpHZr+ZREryQdLyvu
jhGKuq9WcEAEl7Slbns3rLxuXl/X2fvT7bLT6U5sVCeqPCkouQRbuvRUZXCVgfDb
4LRT75vOvYplM4zQOLiQLz05X4oFQvqm3Nb8UZKr1riMAFItrZhndmI8OX4V0Nfz
qf6QTGNhVYBxLPjre6R0Tlr3VrTcugKS7RJloFn1WFH4BC9DaNKj2wwb0Uwop2Kl
aQKP1G/0AkXkdqaH+SXrXxv8qT9ysM6SVAy+WgDWbw2jacXR2ARLHSM/fKJBWjtO
9h0bISu1cfHhjOYNXjxX/JMhcAdJ4J2ipg9q8hVS+VEUudCdDNnQKxkTZ85ZOUsD
EwY5E4R5w/tWHuSClACLr7mu62Lmw5EDDc9/YNAqf+Baj0CtC8LE8cDHz1gsFhTb
AO4D6vyCRq4jWhFln8QCzVvBjszysgIU25KX0bDzZrPtLv6su49ca9Mp/+UDhPSa
uJt1v9TrtKbrxlI/loHtgxG0c6qJqlhA9DovSLgHDhDUWOkvRvGy1eWWyQY6g0gx
td9dX52qIodHiJGx+PZRSLyVBwQAGpJdUtf91UkX/LVdlqQZUlhMa+1mCQcdtFsL
8A1bTJVazOQHgikFoHZn6Dj2Nf2IDsnLBKw+Q4Sa9+9Omz6c9+7ncWmqTHgMT0Ci
/hPufPSFtlENl2qGi7e7i0q9g8w9aJ/cK9xFTsK/cLpKVzAKOombvVg9pwOmteAg
yChC6bXwe+OKPHqb8yAcxjsH5QjYPa2qOn5Gu1jcPmNJw38fMtuk14t7gU7Okwtv
dnmrc0pcdWcnX8lD5kC7f/kKapaIFntWccP1nEuOC1QCfzZxV9UHUfHAlh7XuPGF
NhCuKtVcAtHwvn8voZ9WM83DPciMpPoNOQtnepN0ACriLFuZlMcWc4LaimsSPyKi
mj+TVyzT6K1hC4QdW7k0X3FMKzZIbccvj6TkqvKYHXOcDXM5XUr/8riLgXB42Rtf
2k3z7IZu+2dnFJQhBmBNJnT0qrtSEFzXmTNIEXECdIvH5iDJL8yHio5btmljjVKr
D9Li+UjR4bNbddKOLqDgSsWea9akBrjQr3t88jMnvJ6Ggjt0/kIzADVplrCf3WSl
7bqT7BEMbdpfYZJ5T2JppYVdiMhXVSy6QZqxCy8t1tsl0o2aBw9gdECNP+xj2koJ
A1m+JrsZfBbjV/m2Gn6kZ0dCDzNDjVLh6M/+NoMNs0bER1qjLELLfgxfFXkyJjvO
rFy/rMKkD/08Sn44DlGlCITWb276YbA9aSBIhIS0UZ3gEiUyDoyxgSA/gKN/HPfT
+2SZ3Zeixbc5oxFj1f5Lyfsi5si3qoFPqdhzZf/IpdD6me+48CQ1eWGH7scHfHh3
MX/FZPf9ql2dlol8j0ISBVGEsVVa1gjJnBTLkVTPrTK27oc8P1mBK33RZrCOb2wL
fHheZMwogFyqdaxZy1WP2iymFxVEUjiI6wIZTEWw4G3rzk46feRq1Lqr2N8aBGaF
My3tfUlBohM0PVcQOSMBjOJ3KR7zVCOE1cOmguDKPv9itd2f3llSqlASqtUTlk49
leYMgUb4Sef8ggAgE8skxLbQc4y27YWD9BD78qDWS1dg+ePWKpZO5Lu5Ss+St0LI
e4s6d3VlVYN14f8uo46iR4REVAucAK+Ntd4QcRqGkT8IrVHkeBC804qbk1QsDRwy
F+cq/T7cZJ4omtTLAnOON49WPnJv1MvC3k6aHU0mD0R38L7I3SoQA89SI+TD4wPh
83ppScqOaIdfDflemwGbwQZQFKxXaVZo3EE4AUI+cy+MuyY42DQkVet4EfEVq3g0
NKuMkn4lZ6ezQJPjUtXPSKFrd/PyAeDxrSGvPsXC7gXsJ2wrFgCXp34WAq9b+ru3
mf9oE1RMOIFrOfSLb/2utNXngYRy9v48Nu+DST2AXCL0N8ddS/qUOjlhzkp6Tzyy
9a7+SETyLO4A7JZwCRcbY1Quq+LztpjY1ryhD6Zb0VplrmXO1Ko2nWfvo+TPW9uH
1cSyq+QSITmuG2tyW0QXaBb7ApWdE+DaLlK2oMcDLYvGk/nxhtl0lySTYi4XA/aU
m/s28XyBVboBT2gGBDgApqlGQMEidhqg95g/Pj7ON3+FXnnU12MVvqDICB0xovqJ
LOZGxsX6fnhj6UyI7U2ckAbxaeTN1KiHiPqweiKWiiN4FLjwc4CuCMtRM6igc9k2
46cHyQyKRdxZP4e3wZatGjZgtyQV2KcngQGZDrShWmxKtjgFopLr8gbY0xxCfykw
tLCbhYI0yHNQqqvODJjiMCuLLURTaT7yXOLekDccfUAHM2JdXZq/P20SiN68Jid/
9ryWnaUIW/aT1Kjk3ybgYsPrZNwQHgGcBwJh0rMBj3NDZZm90tXqDIiHZ/EfmyIU
fV8x6mVUZsJ89UNA48Gi1uv0vezOPBcPnKzuWdYRAFMoGW1MVFkX+heJ2zxc0Ogq
xMv/Y/rrDSR4L8Xv3vzdYTtZWgtLS2sTzyHJTTcBPkQZC/BamQAY1BOsco6KEneK
+jbmvKr/2p6gY2Iq+4+f8solw1Sm6gHpfzQJqt8o5PGbGzMjyReYnFr/0aVOTd32
KtBCJ49GX4XRLxPvya2RQ0NHuSaO6oSXz642Un54ccgHBdvdiWNcyrZi+Fs+xjuQ
iCJ3y2KuvLclPRfFtf97ehdK6SZrUJLFdheBVRjC+KhnIj5D8OJVywpNpt+IMmxI
5e69Tdkh1yFB0rUXQSDFnzI5bBZHyzgJeR1FKVmJ53B8jj4cd2A0OAWhUxsvysqW
i8zVTR/wtcxehYteOYkk6fylLXZv1CGmEwR5u4CPSKL3LvK+z2tVJOAhc9Gwjbgy
WIiYCs3aKirbJwDcdYyBXZDOg3QkE9z75utllFC7bKRBa+VHRe5G3kXxHVqE3yYm
8BQzIZMfgtnVA3SAR1G5G2s6NZlM8FkvAIk01BGuwI2DAb9CzJ3V8j2aVIoyN5RX
Md3BYGCwJyJGPjGhTvQAQbKOkEk2Zzz+dURzwswtjscdGhuiG4w060fZqnNNWvOE
/P9vyB3clUGG6/LGYKyyUpgZkziuRC6YJBzT4Pn01e87kasU6Vj8CAX0ylXGDN6k
EwFGOFDSOFNC8DGuQTmI6G9vrCT0rAlNuvfIjUXEOtD7w3MJGulxYIrlavHvSKgd
ctqx40pjWP+LUv2W+VdCwdUOf/+KtuXOuPRxOAsqQ1dH94VPLvXMGxmZC74ifFYH
RjSZuMeEYUfuSedOnfFqeA7741HFuJvAMcJSmIyl5wLOUwsjwva5gUkhR8N2LSKO
WgjlxdxzKHS4N3E2PTlZLZm6T6NnaKRSOZNafaCwkzlh97B3ceLSoUwi2CdBn/DI
6SAL5A9J+K9yWLrZho9vhiDS3+tVh0ISODUU+dleJab1/kdGe6XXBQ1aui8bdHDK
PdHhHFgBVLmWrBCLxPd3+6jJDXZLlwFMWUuYy2sMi46BFF+bDhrqbaML5mSWY2Q7
cBBm9cM2mKrRfqKX4W5zGV9opZKI3awn/BYFszcXfxmF8IYO2p+pGv2SlFsXr6uZ
HIxURESPs9TniFz6AviC8JMyceMLPA7z/4q49ANXmHCnTdlKpgG3ocZVpfKarKDK
blNQ4o+FvecMhdRH8B+yDIVB7kDdBeWUZATBa6BKCKCj+/kvtE2OVLf45w8PIDuj
ZmAQi90sHCuCjfpM8lX7JqdRD4EQauKN8sq0dK529CnHeX7sCuEk7KZL0soIYpoX
lYFy/Mdh5RKNA5tHVWj7h6FuT/vKamVb3jGZ3kOXRB8oBOGCj5GxpbS88wVruH60
ylZEHDYgCyyli2bfqb2ZrChZ5/k67qxR6O6kgCL4V1jgx4MatRFHBXqfRMhm0Qi0
PK5rwBZxPFkTzVMtyyx81JXFQi/CNWvP3VQwCtGyfXOTxu96f1RJI5oxGufvUAhG
TjzZiCMAB4EU586DkmR6FZ2/D05Q+OPS+5fG5sLzXDYvb6LIMYcaHu5IpzmVojd0
hRm3TSzdJag2j6r0nI4WnG0uveOaMZkMMJ4cqYhWW5B1PdHRlAq4If2QyMYJ9mmn
q6JCkZi/7SktuXByYNOGHKBJ8ZnCjSPMuJ1SsoceBFYHA2WnS5eP0aCrnvxnEVLK
5scRgjzSscyIbiyEsGFHQL3kfCIzaDhOmXq12JsvaolljlXB26loaR/0krgJMRiQ
gJOiZzmPylIYYcDrJXr0qP6V14+11e6qcJwQjEm5tv31z+ZBZQmCG7MCODKt072k
YebofYzkpKH35qdwj024M/5bWmwmsO+zIjMuP3fIJHf1OjCoLkCAPtsh0l8MbYaQ
73Y4BmBt27xvWn9NkxQRFCIAmGNIHkZZhd0p7EA6rS4ObbT+7C5A2YKSatUDQtcO
N9j/JT8F8o18Wp1Y+NFqxwMB/PSRqOL5+y1njJYXD3IemWIosAVBarapSoji1KSx
C5kGzLbNNyfMYaCwKc75zWOeUFLNr+9lMCN1DFkNX0nyVQnx4KvOrWoHx5eSM1IE
Qxjk1TA4qPndmnGuIxQnOKHc3DHXWhAXaNmgn9xbrkw1V6SiYYbip/oFEVvSw6q5
xeU/Ok0yXsKDnwczmdPpIFZgFto1Jjm+6MqUdXtY3zPeYuM9z6GaprKMjsJB2UpO
Pyx7PfqAWNa97SMh/wvUN2a1X2UgqMLU/79dPtCTK/BvB6gwFUu2LUOVOabQC+ww
JaMdjjKStRQQrWSsbApkvqUbt/NojUph9xxmoCQGE7X+EfJfg2fiIIkRCAcfuz8B
klS6KToKxTx0B0FsjG6lYEn5JpDv4S8tiA1eiqjB4Fy3ECxKv8aBduDiRDMZx9HQ
WJkusp5PFU+FWx+oSCOM2zwqj4VxjlPizesJ3IpMuZgIBA9EZNkUtn6P6G8y4cds
/czfqLnjPvwnwm+dcRUhdUduCUhkbiNcpa3b9ts4xCc1lJzpsRSVgcIyJXXnxFpy
VI9icCyqO29Xs9mF3rG37OhMUMyb3T3e1u9g6IpfP9Fbd7u/09uqQBlN/h4EwS7m
kpRmUt3B3EbvXhCr2tPU7vvjwOowN2by7iBzxapDLUQ/vibFXqG84GK0Q6bZ4pLx
3HNS64/qMmEWCOLkqiJgUjN1RdvQlrKhO3oTsldiF0DbKzfEOk4WEmX+EaDCTWPT
EksHpO4kT1PZJWZX1zmgY513rST8zQACpAwByAlxLzfinHmy7FOu8XznAbVIPM7R
liZdzty+T2Bm1mA3FGDHWVbfQq6Yfm85imgzwlCJApM1rKv0LAmHvtf7XJ7vtNGk
BqipnR4sogtVQInr09KsGHmVnvkTcOO0p3lK6YepskZRoj82WozLP/K0P1gRnFOf
fmGev9GT62EbuZeQC8UiVazKrnlBEb+za7TK5n0faA8nA7wRrFgztLBoNV99RM7+
9HX31aaNonTa4K8MdRhPpBqGDmz2caUl+yKta6gjAa7xs8PMIVnetwN+Pau7CfdR
rK4PQGz2BRQQQOH3AxvBYjeVux83d5qfiXu7CUGX8pEqw+mPu0ZOjyuqwuK4Cy7f
dKl/e7o6svDz+fL43CAJocr8A9jTK2honxrWCcAfJM3sKWTugCQwqagOvaajpwxy
A0eWx5SxU915ODmnoxf5c8KHQoLvziTYCqtKFjvAe/mFudeDfe7By8V7N0Wfpsn7
lIQbxDTlhbsGJepVwYbObPxYcJYU559hWTatXqWPLpwWw1wipRTZPSq8g0kamXJH
X0DttFDnCQxLRsNqL4uZ23QcQkGq63yuy6LSMtv7Xz0vuLFKjn0pSYuLedVhBJ/+
3OHOXOq5E45w1H2zphyACdrxw7WqYxTt27QYyRTWHoJ8C/StBxEJs5Lodv/MQW5i
Xu1Ou90p357oyf3aG9fSuUcrIC81aFVgPYfvmNAeuJ5uRIpb/J5PmBIGI0npVqkv
Md8bXtEy7iwCf/lsqC2lEMnaXKjo0QT06XW33GzSx8PldXRRUCNzwkU8ChTxCf6Z
E/LMar3gGvgnl+7B8QAfha9antcExh6nqsxVnZpUDSQaVb2bZv+CMg2fc5f11sGx
Wq++z+oc/RjI+CBYdIkE63DasIUgCe1e4ikOWLbvCSDHQJeQBN6PTXvBaVEumqm/
IGmcUIowf+3dfkaQYZoBzuCVM6rKUvl4/4yNbM193GKcIcGRLQampap087FCu7VW
gd4171ZQVicgtYHB549MpGzi0IhY6M34sVACHIhNDB0EAFgbbwWSY+2oSKswOLzg
sOwI4MHqUcYL6MMckuiEon7OnOtms4H3/UbpI9KU6k5mpdE60rsKGvwyv0VTb/ua
a6QL5e930RPeRYchg9e6RMzVWuULdVMLgmQ5DRvUbFnbHU9078+vBs3fHpyiXyNn
UyidqudAGqAHjNsLlYnp0+oXhR7YWcDNTzush8jplduiGkgXW0g94WATY1RNOElB
wZkKdasvQwxyRvUKbQicAJvrPAq08STScWRkFV8Aq0hAmWAuq+wDeM3PWHA5Rf4P
c7BrdbOSGzGGGeSB3rXaKD44sbQhhKc9lGz/1elICKUDQSuqJzY1a/+58LOZ2IrN
RomlHABOgr83kMKaoQFX9qXdL5biD64Z1XuuI/joHImdHokZS5TEB1rzgAz+ZMvV
aw/9lkF6U5KWcMbj6fprwsakaZ1HaE6/wDwpmbADKSV3D+l+nXiw765ww5AX1W4V
6SLOMCeOksrbQ/dWPlnB0Xlec9WYssED0Hx/yw6Nt7JKSIj/jAl1KYPwo2jZnMMa
yDPsBIwhavlUztTO0o84/mNcezfr/wP3MWSj36YypPoenxmRPHzcXET9cJFhyB3Z
ZjZmVxtrgzFXt4YKnhsaOBMMcg4wHn4SF4vs8Yz8cHwxzZOlf4RuIFMjY364Q0MD
A9mmPFFqNW5w8GHjFh+lOAiktqgWdTLhCEx7AvkwB0LqawMf85DrKlUrNopn0OPv
3jLQ4C3zvRz72Gajt4nxHmjGoSqZZul4MWND9AO67GqrYsmmjJVLKImU35a8Qsc5
AnCe5Q3Z2xWKUNhiNRq3TASdiTodZgQbkIjugwHE+8RVZaZ0UXTC/LI9v1kEmNby
PXVY+lwRpj40Mf2+1yClJShGTAAf86Zi5N443LIRC36HstNE8vRsWWTt/FPMEekg
2x0OrjvWKQ2iQQ3Zeh/FS4MkNpX6qGD4u3RhCq9Ohj8Cq2PZX1zGq1nZwGujpG6N
Yh6qkj7KodTJR+gdGt90NlTGriJM0iRWUEn4+04Ko0eUJsyWZuRlxdKpjye8BPxd
FPNeFRaDD1Jd6K98uEPSMlsDE+qEIo18WJjGjzuY6HWFfFrie/Hp3cgOBLlY6ba7
NfsIxxzNtamq3N8l1oqnAxvh60/vzTZ608CYMK7dAVPGuhcIig1+TjstTLR3dFAq
vI1Ifj8xm28dWx1IdGWMrZpDEl50KjgjiitudtIwe5CyOuJBSMnkSr8YOpPndK3R
Db+06rGd3Hg9SogN1J0miCOhyBpB8LBKuwGSA7ykGmYWofjheCnt0hcPIDsbXthV
KVBAYhh7SCIGwJzp/F1IKVItiJTMNDBnanm3x73AgaKlyfXtwkcWNRimXDnPKIYw
vWTr3TmpgISk1RAlhUaZoR9676bUhgPNmRGt4NJVNglvZchnGirDedRntinPN7br
2LHuUsBtOtpD39foBTTxsZFMQ4WJ3r4XuUJJAPhuqFZDxFh4PiAXyD1P8GEef9gr
0POid2sm2r6rm15Aoy8XCemCpkXZTbDmxDBUqa5DaoaxAB0uZ7xLblA3EpowqtF/
e6mSJW+CKPHZtRm4P85d59X8PN+krcxdtKIh9kw9CIayceOdhXtwn2FqCHAQ9fsL
CnrP9LKaMs6VJM0/l1iSW2tdwpEsjI0Bnpcq98DyiN64Me7S1bqFzBTN+u8PWBBJ
AwQPVuqkjDxbcujlJ8/wp9001ZrOcbu/bn5XAyhvvdNhLj6CwUkAOxipZ7Ip3nz1
yVlGEqWr2Re2vxz85n/xDLdjfu/lOGO0nv8jBhO4VJHtVQDmbACXIJrzNLlotjYJ
dae5N9xMv8pbvr8j2pUxTrinyoo/mkTChv62jGT3ldbL4oKfrU8mQnUPnsvLmsgD
tZZL+/HXpC8Yk7rVoP1qdWIetYgke5bCd9LqHEHp3SxJ+9QN7qEDkbw1sy9F6HPJ
0Ri1VdcyMCpgd2xdS7e222Yst0fTSVIrNJ2jNUQeHRd2GhJY6uhjCw6wWndEFpyu
jZvgK+FK/7g4Mp4k+XgvHUbFGyO80Onf0L/KvhQgff3OZNS6vX0Xu9zJyplwA2Wy
3CSmoIT6I/nde3PrpvFkX8HgzNxaAH33PQ6M15djD0iefX1sER71UdWXKTA/WFYW
gDTi7xkDhjPl6obLWBqucfAm5zVBDN3eELSHvdTWfcIhKBBIt1oNXJDwHACBVJ9a
t/u1RK0Hul8Y1fQBXAieJsQ89wlFcVuhZ6VMc34+lgC4PdrO8OGpcy+/fFEA3SLR
VLB8FArcKFy7hgrPNUL3UAlFGAhIfbuh4lXOVEIKeblE90R4NcvpYvAKS2Tv3dLd
mgrmfaVjDOsyz6GC/RUuSE5IYbrUOdj6bRtY7Ls/yhES/ViUFZK9M4hHYniBaC5+
H4icqHgG5qzkxrPWShQrJs+///nHmorI2peGHCVRPrzVDpxv5C8Um+Crmkk/6Fg4
xPkl5ZSn+thz7tKslmOZs2ZPxsEbqJsuwV9Y/cY9M/zgabIKTpz0YYNBcr9sgFil
KWwkz7Sf+bUhvO83YcpWivyNMrEiXB5ct5Y8DQFB8ZFQzP7xU2i2puCm8Ot1mFef
ar02IDLC4zE4PSo4OIo7PqCg8YmH/cXARxwykZbKwZYjCnjX80KKvpQXmR3g7YXi
2Ta3zVaNIDkUco1Qp6VXURNQz+TqVRxmI4KRj+JQtPGXHKtxhHN6gg49DFkpVmsT
U1V9NWKGLnvpxQvMkyaLMuH0nbiO7RsMnXXdQEdbr/F58XocSTcWEn5Hdibp4ou+
bJz3qmYupCDABw7Ny/Mf78/4MRbdgAPRLGXJmSRy+3yKewLT8bq0K/9pZqqWDY4q
Q/Esoi8R9QsOyOuooqFWw7giHcUHHNXIMika5fxJwVV7k6bxoOOQKLOph9pGFs2J
B27VtpYBc7CoIqdc7/8DzrJBwgSmKJ9qKeXcWYozYS5FZ7nGJdN/yyAlyMMosM+L
5vIDfaFFexjjo1FrhVkQEcjNzDn1IGB2Ig5OqQ465FW1BGfbvOdKwyQ4mh3YIPaR
jpzKUMzGGpvCoISc8WHJnkKbIMNe8u6X282NxVYPz2WCbUbJX3/3QXfaUbPScY5u
/DA6A8vVbS11Zn+WzCUi+XsX233W9IpFtLp3888hmmGDJRMMYGFt3hP82v14+LcW
ersjtYiU6hf/IsqoDZDsg68trvR5Zn+PbY6TLAUwpo4gBMCfLaNLnF5VBg8bpExh
10c/8HTn2MdMVyU0Oh916in9MqRpJ+m49zyXieV9Hcpy7lymFCQoMztGiv8wGAxt
d5t5IKcwGxF+YhbD9eVKrCulHXakqSBVGbwu3MucGcI/TW1GNHSF+3zwzfUr8YpT
MW/jAxGQrcV9w9WDkWeRhmVCied8X8no1XOvjLl57JIc1EuSfQl+i3y2tjfAjoE8
k+ILlnQEKYoAXv89H/eJIAh4nTzp/aNl4D+c4xObycm+qkxVYvyMwgHu+F2B4AHz
TyEcktYcKovoJeIsoxAAnURxKWZOJqfxODhjH8uXcOMC3oGm0TWc2Fd6rPYLvQiC
XM6S/wtYIUn3DLTQmIImdC3a+QwOd+m6HzoaZsw/8w4CB8h/s9aXg5z8Bg55knBO
OlhfouoLZDtdAJkqLgM8Zo7vFB/bUSGXv4S+PukndupC4oXQfVYFAwqB0FRqKmcC
ptIYp6owque/Q5RFwn4Oyoe3fsRk2y8t0ogEe487THS2obxsPJJABk7EcHv2W+vN
H8vvv+v2DCBUuoI/3RFff3hvjETQ8TPY51TeMu1yQUUjA1MeWVIBuvq7Bk7hFtQT
dh2bC2V0WWppbOOisYo+xZ1yVIKcICxfX8w7c/fxvA6fcGX3KGakPUKs0bL5vXTs
XB5vwIXaefIRNkedn7L3IbOwFDtFSTwMIvd9BXcpLc2ZjasAw/4y7/YWgZlHiZbQ
ZOvghlUjClBnNOWhralz8cmhZtd/UAl5Rbtv8yfv/3bJT4dHSmYjhwhcOxIJIEXi
OHgzPhq76+NL6y3DeZNNzr9CPnGh7Xio4jRLodjF7i7E9XMJVIaBeAfv1SFavJkX
V9E98511gwaeSFC6SevW0mYGA7v/2XsVepM+yeVeImtrO2568hOD5rcgGrjXaw7i
gIrC14kZFslxcoQv7obDfIf2hYy4KgkZGCiqSBoi0rnjkl6WHkpBBFg3BZM35LIb
3LJ68aOqnML6BxH+2SS0tauhSL/dyidkUi07mO9vbhc2qNenN7rk3QF06lVY0deF
gBOhcNizq9KKh6M9b2QqVdAoSE7trsqG9DcOquP1g1qxYf/h9zYHmUH2O7yEuGmC
+yu0Nwf0Ai5pd3+uP+Rk/wuIaVVdnDOoVJNFMa5AieveaCiUT3X6Dm/dmHvBsWj0
bM2zxjY/8PUwbVaNpeOQKX5k+uL7VN62o50fL1pYWPco2XIpH9fgGrURiEcwrfWs
dAvDfRqJEDLihPHYgLZiwD6ZQLkbigdO/79UTkBJX3tqauYq6hSeTGEOI1Iqbl9q
fH3q/gtkQjuU29K6/bnjIadL96cU2Ig97EZB6i2JcD/fI3NpUWRB8Bkq5Y2Q8YFZ
o36T41zPwwPObeR2RqHvVbVHQY8YrxZTYO2hXrzaNQKl0srAZs39+iFodSNzK636
o27zD+fzCMxXbiQiYroYJGZkwHAx23gGQr6u9VhDDP9nidfPZ7M7XVv7Bxi9aYx/
T2fc1JSRMkGb8a2N63JAexneKMRebuvJqpk6c/Xr60+DSkCWJEqh7ysTTO/i9vuG
7KrAO6Wu3hK24rB/8MViAI/fj/RXasXLTqfjmfNE9kxxAC3/jbC3zRk4SYKan0pH
UFF/PTbP70KhV5hwHvxGMFn+iFtbnpJ/vSiD833J35mjMR8R+eXNSbCRxQs4LCsb
zbJHP/9jHPP3dd8qVNjV+hjqyJboUQ3ofzMkYiHlqCcFqDAOjUk/YfKrDDnDHsVZ
wI5PIPkCaWWIAOZ4UzdqPJFwm7BZAteYECylG4yzasLzbkmS9TTwKaTU/R0ELCVl
7hg2c3zcNzWFuB1iww0g4RnxWeiffjDXerq9BbWCNeuRKYpII2e5hAb0ZwYp7slW
mgk/qnw4OFK/6eVKpVoFFXYcPXu8zMb+qwGZjc1rhluuzzWG+L75pUsDnTW0oUkQ
8/zEGRqLiLUB2HnVpdlfPasRVj/MhoUnZl5AuoUI6KlPxSO5tjdbB3sp+D2sTnLi
YB2PIoHhfonoGXeBsT7VUw+IjSKaZ2vE6XW0We+tk3gN5SgDGQ8szt4CKOIJFq0i
ghzlb8x/osgCfFXkKCnsS7sQdd9nXhhGlY6l8uIIbo0yLLv65l/coo0eHbZGkrvL
32PUjhc9nZWWKTwEFWt7uzgMKiOa3dAobCsqMEIFmu5CTJB0Y8cGuNzPAmbfAYM1
rE7exnGLIq0kehRaKEKNx5O10o1r0RHs3YrPCci80ZIasAGySNsmsMd09J7u464M
wB7u79qn3gxv3yhSnU14noVs3M8L1fWu/OmdamFiJko7utNa7BxQEz7c9qqEG0Mw
MK0KqTD4/TmZUBQGCFpZ5bPIwbR9WpRu2m6IQ99WQEB683FmqzDCywzASvcx2RuZ
avXGyerHQRKSNexi2KvEc7OMfkKXe+L/fdbhMdVOgRAIWMbmgZEE4W4LLLI/l+Zt
LatuM1zzNqM9HPzIWRiOxYtv963ujZjWdtlPXSf4KaXmm3F/+IuFogbtqa55ehNJ
O8nkBYOMTuvaP0t8LpwnXBCyX4NAdrIyP369jGtFsUOdHTcjb2b93iAumbAeh9Ez
rSzpggxqLfR2BUsSrWYd1NefL+5ZdZnoBeo+K7Or8m7qpUeXzf8uW9a2bd5i6WVD
QJv4plWirL6jbd4DV4dASqmOUKUmeIssPiEJ+o8Q7uks16eeyDpxeRKOA07xal4u
PrLU8tFsj+yt8doRyJd/soZqxYq276qGPz+XxkL+VKRODiFzG3Fury6rcW4Wq07S
uGfQum2E++8dzk1unXj0jh7dhmcOoO6p4gvLNGuXrbCKnopDGv+Wi8cFEabhFGdu
Kp8hyhPQCUFMEOHek+9T6NvM4DZMW5MYDLVfbgONcVDocMYrm/iy7ti+6ZyNA4sn
SUJ5wJumPusfPEYCOiU1kSf18hWv4tWrAIxEdJ+GZH9K3tq0WWYJfRb9uvBFU8zQ
0YtxLpIco7kf76gr95mWK89+74slGZM7T2BjZPEoYoWWjVwPzH5L3aG3vvZU0C5z
P+EQcwXyLSeO7fDlJg+i/F5K1IDTtPv/p2GBk92nEYNZmmxN4qn36/t+tLe5re6t
BUx1pVBF3e/AHDzlmeCxOqzNzTnEDjMTvqb/iO6wWMbItRK/o3RErCj6X5aSL5bl
XRQ2Zp2sSez9JzfzrXL+1btkfEtjGYOuuUsZEtzwlwrY1HO/RRbjHHs7bt1npFBr
iunmCdvZQ0a1Qk8XSCXWqX4flcU9Qxh3koGPauwPDnS0rnDYNlb45Rwr3H2O7Js4
vR+duVEXe2OIoeQUyijVc98nD5RhATZ0tCbHNUMbcdgY2pP0/2xqbl8fPyUP2eva
Q9vUQ6JKHFXQ2r9oQr3f+5Zw1CqMSnuyxh66ZoP+CSB8OKCbU10cVN4iNdumwZt7
o4sW6slOmJP2DB5DGaeBHpTtm9Q/czB+Scc5d4woTMMvb3t1QWqoOblYn9AEkUs+
4wwSgfN4laag2WkNs0tL0CBkMWFIsuBQP6hoV9qxxE50wsR0CfWxiIJVE+KLzwVo
EzCD6B+QpoYc6nsZVci2lKUKU751yLd4f57vNGspyeUghJrzbWvDdv1vuHHs++9+
NlAucBhk+gq5UguhXFfjuDpPZlHf/XzUi9cdQXZuT8Z3hQs+bUU+aL+XPwDKOYK8
RVFDUM2RgzDQN8gJKHqfCqYYLfvsZh7pWXW6A25bqOjI8mXrlynxnFZ19PtKL3GC
bif9qP0jGp8MY+cd4Vfgp0S8e1qyikPeBtXVdvN2sjI9GFkFvvevscIIWB46zvNE
XGsA1VDJWUXER4p/I8gTJGCm0146VjRTyS8Cfe4HTm48q9LOcPju9X/vVk6Bf12c
mT+n84xe+o/koDq8ZhQ1KesAmvkxpCGYkN+Iplx8iOkuTJa1gyBUadzTn2gK4cZz
iO0mi3zOJgDpI66WFzI7ib4FdLyqZpLGZDP3o6vMUfDROqPs1f5FsA6TSI4+apih
x3G/ML3jVbVcKiA4pwlN/1x+dTTYd57hYKe4uoMzsjA59fP7542f+3FGc8I5t+Ek
P1z2m977FNl8YBAhCaVXgVjMGS9XtGUrq6CJIukyuE1uN6pJOFmBnmzcU/bJCWFa
5cSyU0zh9y/8S55wsmFolRIZIoHOwXwbh4ruwIIpPowutQdAG1CTtHoDcOj8k4Ww
MvQDK8gd1u8NjOm0z4400Rg/jBTasZuNnSg7wvmvkpR1N+CVlr63FrlwIwb6fWok
IVFx8FXd4EzJfOr8PnULNdVKDkGbORToZ+83UzH2TcqeW9QzsGnrJ9n5AB2uFVby
nDBPQcLXPyHTkwX0hYKKmebYtyJWzRG9EdEyl0WnqNTAITq2E2IMCQ1NLVp4dWS3
nXFk/Lf/JbQSERuQ4/YSD4tTM8qWB0vvXC7izJNkAmWD0wcDbM7lU+Y2w0XUx/e2
J/gshKSB/k6sePgCWHMZ6cUbyIJhMmGxwYj/8QCZ3yk1HFj2+svKE7N8uCgQXfjf
0GGozR6N+QW5vZNRQkgh35EJT5s2/C+/A7+LtSc1oWSIIgB0/DFHZNdQSh421s4m
1LAwHRvHniSVOcrarDPubOR9uE7Lk7cIZ3pSm4yHeMt513zi5dCJs0vKPnoNJmlE
T5pSIQB2fpO8uRGS2cHby4cHTnS4eXS6sFpQftO3XhthHqJ2DPRfWP+3HwDdfgPi
wjpndZcyxRHo72/iqHBxQBeSH9LMGKAbukXapm/VEwJ0Urhd9qv4GklsTfA9dupu
LbrNQRN/+PH/lhM8xWDzbszDVFIzwJJxsMAMR95WA9XotL61z6TjAnT/iAqp28aY
YJoAdNeRQdoOUMqgo5HgSrniG91h1XKp1FcHwr8zL0xcO/lT50vT7UcTyirJP+a/
kQXGWkDrmWmEXEGVxjyhZ2K7iWyCdhoqrDSHgDYeHTG9V2oNKERYfP6f7mJtJEE3
Ck5caXrD6FtLxcbUxyg/Ji9k4t4bMISm+OpzmIF6xcMGi6zEE9NlYq2yKiN0EBN4
Vk0kgYdXiq1w7mq7iJe9FZnaiHuGX2feIFloKwl0jj3XoxW33HelNjqYGohMTljF
IcREyaWZKp4gpAeqZOiSYrQOd2An8cW9SYrXb6YzRbcffGVhQB6cyf2gy2nNbVCS
R3+6Akp6m1Rs1Z8CEKQ7lOqP+Dl6fkz7g2//YP4xG8Jk0U2Sv1r0RMbjA292iOu2
IiH91pw5Xnv+ian0KQ/MW64v/lRhsUgnPoTYv0wpeZ9BoNmo5grK5EZhiUJzYLXZ
DIwjrLLLnsJa57ocvMHT2DlWmS/gz3c4uSUOi5yM2gKtymXiLTszsBY+zGCaJHHo
Z3pVtSP8mOwpEcchuirfuY2IvxzM6FGu+t8kuJnm3tw+F1GKScZv6L92D4V2y+YB
vqg/o4hX4A+OzJWecGRjueuDU+pwqvvmQ+ZEC+tacza5XbCqKEv6ryE9KP0v/xub
xXhP2kS2N7LHx3DUqFltfcPugh6E4ZdJKegx8D8a0lRaQ2QB2ZfHJJVDgUYFafLP
2CQ03w67n3GxT2wZkNW0cW6k5kEVC7GPiu+cQle945ZprhJ1FOBagjVt0qJF0tOF
qZ5gInR8qnSIhsivMWKN/51EZiS8/Qmb1joPcb0ooO5rDMHwQ8Tmy2RaFn04Qhpr
V2U3Hul1RF/hPwG4lhcxkYr3tUV6LWOON3QZAMlbiw+yRDgOFNgyDmVr1dPj6K5F
zhjIYCsqFfl7Q3zGatw/vJhj/fUd/fVpw6P5vTf9BK7mN2Gvr7NNSKxQBJVLSnZE
IcdUuKoGLnnotcXspcOL6blTGYIMy28JV+p1smreL0kl4W+YWTvYvogd/R8au/g4
K/mGVQ5g5D/NE4Lfif9rn8s7ZJwZE6OUK5VRb6gU6SmmM6xsaVecZAwyklhyEiWk
DYKYgU//XW/gqvpBNNv+jYbibOWJc2OJRfzrX3xlUn7bjjbqlzTQFekiJZU/UwhZ
+t6KlvM5fXBhBBpFR5i/+Koc4Q12/SPSrhGYquRj9UERILmxGPXREawaI47aefMT
koLxok0kfMO+Q/yUS/bxLMAqSMNBwOrDkG3PTdC1yvKWRf4dAuhcZvHJRF3UtzkX
/7bNonhJoa2dfq0AE7SQv27LC24A38U+px5FlR+qBAVqi/ExiammmaaUgomQwG+R
fc9UsawU3PmimAFSaJFL0IZiEfXObJe1QoCY8qiVBdE1FLrBbWZz93sb8mLjWHi8
exX9U95A5Xs3HZ17iZXdeCu/10dqxABaXoE3gqVr2Z4V3V50P6u6xmOtqVhm6W7G
/ykNxdAKZ2+FR6dA9XkrVgR3XKYtLmdbac/rldemqiUrsCXESfZ9UM/8MOYicsYh
BECE0I10FGw9Pv6eD+ZG944zgjnxuhyXSSGq/KFTfpDd43F7jKcKyvMG6V1J8qW0
j97mGgLbWPPa+0gxIh23crhsc936zdcdyrFphvzeKLvynsjCqkrlOsHlwcIeQjPb
mTMMWZor0P8YxEmRbfWFw9K/rhwny55KuWjIgsXpJJbeLPdp12+AH/HZNq/51eh3
+Heu8ecOlCm6qAHUCAvTgUfn+IvDSNuaFJJ+f01yQhgoy+Lb8tWgbHs/Ya98/0dC
cKY287LM+GSUWuLCdUZAdAByPNbOLzK3H2YSbPq+NP9PsndUO2RGh5oH3JY6wRAl
zGzMkiP7Khy8Xqg4ziVrbueWQ0J2lw+SQyNPsuJ3fGjWGyLrvM5U1S39d5dAUoSi
CA2LxGAdp0B3/15YfsmzSGSjwubNYqYfv62O97wqoHAh1LYpj1Qumj1x8vr/Vc+F
8iLAhIIDr9XfsMMNMUqfkeqPyRY7wkv+8H14ZRbnrJTbGVPzxHEeLlZ6XXvy2Twv
THRS75OJgq3uw40X2TwCwa7MBHnWIXoax3xV+3XSwTFYR45gkb5XeSwkuqvDKFL9
KwwjXuvhU/cPerIdB+PZfb+Q1n0kDIPlZEKexp72js3Sg+8WQ1I8J8R05qUGHHPp
EzIXhBmbtkKHihbFmxvahY1fGsaOqeVII2JwpTTO1J5XRyKCqlKH7ZBPwOqpIBNL
BLw0f0J+oQty/DW0sqFFMJpaRpTHPwBGX0jrvk07UiCkJKqeKnCbqOqFleTfVD2l
v49YVOtJIU5jTrdPBiYc/9T7JgCphN9zWPPOkVhk5o8S6DiM/xExcmouyxpqlCdE
kackZ2SbHhBCUzP83DtiDnHV++X/Cyolopzu8hlfBhcKvHjk3Gfw6BMI9wKOZbTv
YnPjzGwgLYj400hAYOH+L7OZhAx+sXgWoUxRT9fwjKBpRNv8wMRlmyVHUUh+Y//I
Di9swe/dHnANVbwXfpiiV+2EjrdNCnjDjQdVM42IJmLIT/w6SNFVUtoNpsjOBHjW
g3jOp54nP1zq/yj8jaEd4DlwlZOgIPJQrNjiWdSxVYgoYh595xGNPTlYhecT+wQS
tDaF3UmNs5H0lWW5celnsiaWk210lymJE3aoYY81ubBHiCNBYqaN/aC89ye9hqTx
S0phFyIL4gXcdH9QGny5/qKOZjml+IQZpYPBmb78/udqTgbTakIFilugVkh1E8rf
vKe8n5eW8cHMKLTgWol+xuBH5FLglS+u2hnSf6fJ+F2RKXpxuF5B0/3cCTFraS9T
bU5aoczPRe4wrU0eUSDvyHtX12akAVgkbuyawFfL8LvRQUla5xuVGvPs0vQjRxBD
unOi4hPh+eq3TUW+/SMpC+EOv8JRhCRSpdhG/Mpry+b8pBGd4zMb4Nl6cbqbHpNh
9yMLVIwGBBcLjiloKiAEcrXpOQ0Y3OZpRAmJSxV8MpSZ89FuoAjdQ/MRVzuAxsew
W7QQXeFGNUy1pe5y8Cx8UniV23qXfa0eY/4C1/OWizUMI+Iw5cJIwchXd/H9BzFI
YcynOejDZ+zV/n3tVVbs6De3JrH0HqHzZaDihs9Yxj02q2WBl+VbdFFzME9TebVR
j0sXCJgzLoJrXFbJ5x6znmR2KefDbnAqh6rZ3YQq9eWYzQMfQE24RMA5Xhfa3j74
zeILN3lkYp32v00lCEATEgPvvSrPDOOLRrfjQdiPOrvqqFedfHSkYPOd/o23r6ey
dl2e276rOiwzxTBnKqDZwuZtI9pC47fWmb40DUZe0ou87dazP59E0I1RM6/GQXmk
mh1tuXYPyh21/RixEXhb2ZUNP975e2WrevTs3AWbmdrmb4wBfKZbsi/AJ+/OHJ7P
B0H0ao/0phpTnfVotD3C11srdkD0YE9yfKJ2PZtI3gP8IM5P2wCGHPdiQlSqHmyi
YLmf1Zs9laQ9Cgf8RXHbUM5BAkBj3Dw/WbcjImjL3xRvbXIfXXaroQCQZ3Nh1bWt
40/n6BcHVp2rsnB8742mXRslWP3QI3U2TRFupMc+ITli7JLv+NYP9uW0o37hGVAh
HltWDiGDPkg66EeHNI+DT5Vg6Bpa92jV8q53NQEQgckAPMT9pyPpekAaA2qpd4yw
UqK0wXJRdUSHPcAyczOB5tuWg1R4s/HIhBeKfHkOVfZv9dL+NI0nXCUQA+OfaFYM
pL2AhyQ9DDN92l3kY4gr7l6pzdOvnx0dGoyTen+5Xr3aMrzhro1xGoOrm9dPhyV5
Zuu4MZDNbl5SmnmXeNXV6kxOeaREslKuydAKKAa1gR1C6Pj/Lt9dU2+j68tFCjM/
8Zp5fjmJQckEHN+0VJUKbewIyyXUFjLmbOFOgL0jw7zg6ZZwWx1T8q9N6Rqb82Rz
HExOoMulKSt/qfZOZdLfq8kygJq8xl7JI8g6HlV4vlSHKuggRsfKqfUox1lIKEMy
PCpsfdGdZDiWRp/BmZswp4eOrizzx5PH5uI/V35/D5/vSrOc9YhAnGkUbg0HrCFm
nAfOMVHOxlfvHKsnHGDGZR2xT0KHPSRm/f5to/2lLWxG8D5V59WWOFQLW5c5j0IG
tA28cp0FHf+OMzQKtfY9j0IkLTSfyPZ2VB1PHYgjNy3HCbtIf8Od5AUsv5/TPy9J
rA2VU6PqcduI4xk7olBSpGoDEztHTddmRVtsU+UHQrfUX4vtECnDjPB2znQh09mh
/rm201gC76arKbE/WWiuEJBuC3IZNpc26D2frXA28m6Anx/pa8gGtjNM23h3/Bd/
gtDpG5j3RxuHq5sz5KsU43L9EIJnpGYn0Wh3l3OgOAIgqSMNe9C116gdPrCo3aTx
ximivnOiT9eQuYD4zKDtd4iwzJKtsiFrP1Q3pDM5/4BcPrHkpb7W6RwUC08J8L3p
u4xCo98Ix2UcyXVnGhFb5wKm95/sVCImdbsRRFrNP703Bjxpmgp+omvUK/GD5NDN
a8eZxTzokExv7oFobLauhVWXF1+/el1dwE4qE5kamh9hGuZsHz9wD1jWtRLadODW
q6ZDh/2/+FNELsla9b7s95+geZzfr34steZpt/MXnPNsFonI7CgMigMgcDNNwrW4
QaXDbtKWvDOBnqWTBqOAfpgFjJJW2gF+C7lHukGHrwFpXUOoFsCFYf2RaoHG4OiD
FmH9Ksy846R2hM08oWxdQlG0uNiZGnLoosDvYmPctvQgtGt/LDTsXGiMRFXUCiUT
GJ6Gv0u6aMOKBeMQ2nNYT7W6l+d/UftP1+IiAPJ4Qy50nHbwqidWb1XLR4NHquQE
wTClzJOkBTG/wrz3gidxS6RtPbcExHJVW9QkVyrcRiX7jT6ZGImkHewtizWOGcjT
E3F0zGenTikaS8H5rz7VU7Q8t3NgWq1FFMknlUFkgIs4MBupjk5zOzGdShnFIv6L
cgW5trMBlsJSIiJP8nRrmbNgjLffT2qCAVjMNMWm1JVxOrOIDeI3mLgI+HHWVogu
ILJo12n2GFLT/tJxwb8lQx9zNLCDRsQ1Dpfz/XIpCll+XTW0Rw3GyjF8vFC0k/Tl
eE12tGo7gS3G+72EB6+WE6Oi1aWgUYgZTjPu/6a7J2yZDRzbca30CWMrkBnnq45R
XLAjpA8t8lTp2ZTMs9gpgldnExTFB3z0i6UpLPUZ2PFPSBEQoCxuI/LvgDwy62tJ
pXTLgZqZMBt9rVULH3cUFRbpingHd10ArnP1DMtVDV4q5FBFpzp7U7e13lcZy8dP
ka478Tz+XxZUepHAMLOYpT8hfvPeyBn6322GZ4yusDzI5zu/UklDdR5WuYWCk25R
3Pba3U7U1OSlGfgarLAIoVfNiCkLJIP7HDpJYm4Fs5knEXC5DdjHude/6bHzbh8k
E/nmdb63jjcWBd2YIuB7I8btJImOzAJ2GTgFSHQgI2yZH6XyLcfKGl+AwCHjZSYr
UH6xgsZDH8lllcKri7Ev/yACVf7+GaX3r5I4sduE2Nt9RqqI6jKl7y6byYR8nenj
UwJsqgVtkpiGNWG78gkFzewUsSZ3MHm6Gd7s1AHF60xEGr/smN+grPLP4U126DLP
I2sDx99E0xjWCs4v32J2uSras2sGwdWFSJdNii7vZjtKisSqe0FvDY7K7sfi8s9c
KAS7YoCbhhHBB0BtwdIyIYr3UZBIhorYUK9OwV1LQzfjoTKsD75Lh5V3MA2Lxdto
9ia74D2EjQSiOHS1EJTXwJD03uIdK/Rzex0Ujl5ARKDvXK2GRllF0A3w1A/b4jNf
WggtLUItW2w/g8z0/DUuIsUx/2lUiyIFaE5hFI1fiCjfo5OW28bVr6HBNDX7Lchs
LALklOgANh4PCv7APBhDci/CILF4by0AgBy/mPPVCOMRMwCk5AzQTsKplniM4Txf
3K8L/Wp2bSuL6A1Ax4++hKSaAfc0+lKx5wkFil4F1/xCL/xSzSR5Twud8f6IczMi
/QdxGpwjDexGvtvm+kcAKtPREaZK+6h29EzCDTleMqBxAcJjz5imS05HBobpFNEn
SLE5BaVSEpGOdt/I2WB7bY7+PKHVbZ0hZ0U+yiFxHvEli7FdvK+e+cLzECvpCf0z
0SLHeOB7O12sEI6z4iFIlY0zLNeKPX7qHJG8+p/yyiLLJ9qq27NqQuObu4HgqX4y
J/mcOVonVhYz2/V6L5zZTCytFxnwsLcbTuB9JTBsJMt9uyTpH1WI/dtCSc40zng/
/jnVooCWfqPHOiUhltwRIuEkTPy2nn+r8rdDYNsx2cvrUaU52fLUBBVlt7BOsEpi
NoFcKMB3cXZDSCaVLDgcni2AYh3FI/vzykVpyg/eCkNcSIjUg7HIzngEORSmZQ7L
CU+Ul8OMvWl2bwCYFtSlM+ZTmpiEz4JvavkmRxetQUAi4kJ4fAnlauPdgkot7T1p
/4rJYfzLjRfcHi1jiVGJ21COry35Lzo/yqrAuNXOdgD0V57QYcD5BJWQFpEo8gR8
14+ypKKMgFl8y7Hdd1U3rnZR2/0z7ORnYwxEKJ24Q/Gdws7THe6YPX7fgWyq4BM9
iO1gMzgcHQ0c/Vjy5xJu2SwGXgZaMs9J53M482kPLHPK2bqK4C7+d1QvdddnsBya
Snj06C4lxKf9QK2ySInwHpNIWg0D5Km3/42SlhRzoz/3AYAVIELnUym+H4iZmCpj
n3DrHBJ6YRAmFSyALlTb8jNgLqPdR+2pFZ2kkyTyELfGSGR5kP9AvD67q91uvp2q
6ttvO4i0AH8hZ1QjXio6kUAvm3oYtrhUBHoLs9QL9O+2tU+PoHibxxYPJbcBFCXN
WiL9btfGk3Pgv2V8XtUdWqR4xCoox6153qQj9jSyiyxUpMZwuwWaYRt7gFEPV9Oa
+hcXzxXwem6EP5HOxvnBxWNABP+k3KxS5V4y4s7xwPnAB+giI/2iTVCvefXAsNRQ
Wv7PsXIbFSY+xJtsmtQl9AS+xRlmGbWWnFS2lJYVPKkvqYhvHB2UPcyqtU9a25yy
weMbyZl6NmUn+7cM6cyWls19lHJ75plrhbJGkGlQwSBXMepVfkB3hgIDmN9t1TGG
SIY8br9M0SvfcG/zCL4e9RX365IdYSeFQ1iGIATWe82iWQe2JbRIIEYwi4hzB2mv
oFhhheQ87Ym0MZJzJ/krlGhxXUtuqVesuznd2dcMshRRYVu9xXp1pfCnVQggdPM4
dpd3foagP0dAUzZrYYQA+sd4+VCChTGRh4nnwrTmMGDbGgpzWs62aL7fuARZ4Tcf
zjYcM1CVT0FJzTl88DvQxCHq0vlAIBAuKyRHbw1/DmKTeJQbSyZnRHLCZANgbzVd
skxJKS/4BCz/rqsV2xjiWAaNo21RQ1MFjfV02RQiXl6Iq+1Xm3yQNMVeqfYYzSzG
msznxeWiGlOw1CdJSZpA92N4FQXrQJEUKwL0kMo24sUsLUZoGYYXqH9pR3Z7iZMh
e+eccDH4nf31gFQU7FAXoczULfXX5eocQXihL/XJ0XQQxny56hBz+01i5hrBbJXh
lz/8CHc2qtWchT0TcG0JSQawHwejnftN7iz1TEKsPxVvrutTVW+gZdq9zeww/NIw
JGchGyNjpBC3OnYqEGqxxWVltT7WRbwYWBs8mQrXQJHQUx6m8tuPl+GlZtW8dvzb
W1ez58A3CtcBV7MuEe8nDMzxKdKxK4FcOr02Ars4RoqIT4BVh/XYPf+QKneaOsIj
kiv+7wIIWUqmFsWU1PHdfXl9JwxhmayKnC/dHa+eaV7SBwbpx+2R1GW5AOU1OVL1
GPa9HDIwSOX0CwCCOHMoP18yEM5gIJbl9UJWi18zyWHoya4OKWrMsjCBUH2ewtbW
tpkZ7efkkWAoVt1+3KnrN5QRcPsE7Wzs1P4YLq6KYmh56lOdtRTuj6QaeTVD8wtL
wewGdY6qMcuf+nygz0QZoaz5ZdutpBUhaewCNcNFBOzXPHA6wsvetYudtoN6GUVn
OP3tZK1iTjiSK4JmKYr/R3aof0LQOZHZEjhUnYDTzFokQdBrMqDWQr3X8T4NP7T2
UmtMy/sBXafg+YILxaLUOH4HWFPoq6f1rHeRHL7+hOuCdpqxsPxkO/9SL0BSlFe2
0N0gdeWQ0LaHDxzgA+odRmo4Jy4ZOf3HBClV5Z9uyux2eZj3s8TDkN0h+Hf7al/d
zcgB9A/SRr+XRU3BfAlF1pXgqjoaOet06WmBrXZ4Yn1D6HvfADrED2qTtLC08MnR
oSAxJmw+qPIUxH/okhwgu6Sajp8e5Da1JOzNZO24gusGZ7s9lEMM9b7Hd/hVVH53
U9W7Hguy+6uwnN6/5QkUcgNdEj5paXXExnepW+8SF0h2u/llPC0ySdKV0wmkfQ5Y
N1lg9wJa6evDcWEzdZ2zX8puAnVFVTojs95hZOeP9/x+yGPeavnCJTb4FutNyRUC
Udu1Dh+exeMxz5oo3MnRuCTDmViWx0JrIgmXvmqE7vZzMuaRivJmPY1EnwF39fin
PfOqrGl6C7dYHJTyLpBuUGt/eiKZOqT1QDV9+o3xs5rB81q2IDtwTLN5tTIrkgOA
yCIc1UE7ysx6S5yuETBRPR0ZzmqqXPb+RM52C/2xcFva1LqNfxs02eetr5QSBnxs
/KwzlLfEYw83RnvbOpRAKqZD4YaHVEef+PioKgvdAswCO5WpiY5bUK/ROCxVUO6B
sc/4zK26x4kxlyYP45Kd9NsVC6z2IP8Cutb4wbGu+qYsyl5cjQpuvj7fWbixcEsQ
lry8vkX0Xp7NNJUR/WLrrg4XM1XTjj41i0YsI85tQSAtzpVW9zzU661aN4t077g7
qIqV1ToDV0dp8vfKNCGDcdLbxVHZjm5uadi6Ygetrr/NSBXGwY1sFjjLq6rFGfVo
lSkSENiR/1D4B0Ej3VMkg/DXT2yYrFK9JRZ2HXma4ZsLiGnXDeyZX0fYncyEXKQv
E6wroQHKJYbdYkF/IM3t6EOKZzrZsusdsXS/rucyYlnXpt4zrCFve69hv5Ox194n
GgzQqeTBRDQwUIKW1vSfLl3YDnt92mSADujh737WTs01RpMnni+Fq2e+G2bGuzNE
50yMZ0mxrXT+AGtUQCsZ7V76ytzIy7HZzM9vwewom0okUssul5+i/ONtRzY57CHM
ypm1cGTnVnhVomHhCjeMj1CMsP7WWXnt29zfvvG6DSen/SaXXaJRsm47Rq+ycMIu
hLIImQPZCs6F+UZ5Fob7GMoRpFrHqMYL7MdxmM3yJ5J0UTvC9CkGjYRG6mh3onEZ
sdMPUJoRGPEIpsQFRencOOy8c1t1Oab7BuAORrvTtklPeAjA5LtpgIjZLs7IAwrv
QrFxRKqFftmMN4gpdHDBYHdn2uGVb8ufdnY/quHrq28JyfI9LWb+VKzWDaIx81te
9+IgkUy1jTnD55CH9W+jvFEjMb7pTtLi0pb5CIjx1wAdp6jTVD+XEG1+4ohPCy81
jM7Me0K9df4yTg2hzPh4xleBU/Txdyan3UHS/XqIgLNRVqlGEbwyfqHli1bKZ/iE
nd9Xt2mS4vnKaxcel/vNO2aTvDQESmXegAevFEwXRlYCma5s52NgRaaPN6sxB93U
EBTguMM9OlbDnImEKJP+CGkC/kuYGedMDDZNrTHJnc+5k3KbCe7t4Nqt+hDrisG2
C+4lsUHVaBMwIiuKsKYf6Qt1DLD/8nLG1PnBI77D70zxkoZoUx5pLcDj7uUdGbOn
y5XSm5yFTyvn0EsrhJMcOS87w3oto6LdfISrvNkHd6xoel7ZhO1UWnVEqI4eoykn
sGvDslJZVaQzxz7pN1zrDc1AAEOvs4YNB3m7p6wQiyxBdau3xpZIZoiaV0ZqTEaB
ym8uO2D+NqiDFUKor0WxXq16ZSR5FJe/jiIw9Qc8y/EKMywDMDQ0lF69vsT6nmpa
jx1Cz32IxbZT6RdceO3918+oPQuzK87dxuo9V2CYUy85O3/NPu6vGVKyMlekBxFB
g74Bc7G+05kgWlbxWPNQHHTztPvUpFmYRpOxX9s446zWT48lWMVtGG93TLCXe1fU
ZkIPM3c7ssoRMfMFvfKcMhOzRqd/yE4yPFsqfrzZI8BaV5aKb/JH7b9r8L4oIfEm
DXnjSyI2tO5kIwFHjsYo8gMO50bSztZ+bGMpFy4f6Fk8vncNj8Ux5mkED3wp513N
dbfXRfm85/wQmfhn6CX2u0TrH1McsvGPQE8tNZn2UorloOF6n1LxoB3ClINFY1Vt
XUD3ZHtlJmVxhALPbUTI/1H6LGAByALXj+RC2sDA2ZtkVzQ63hH2n4LZFwn6F5ZE
C/t4gHBXV4Ug+kbiH9QGrc8Q5foYyfxrKqb9CVZq29dOC2waOcVqn1MeXYgjRRYF
JqZKfCNGqQ6btoJEtt4ZNocn/OgZZEoLh4URC8RRoJ6mUxTCy2UJvmdAVQ2ZYYCF
9EWmmFnl+NxhHv2Hsi+O0PaVbJCi5qYS+Uc/xLUs6autblr+WpQ0RM/2pD3jXjnQ
xgPkAvzQTfndvt6kdLPr4wv13PR2TNj64WpHQ+bXg9jZyWEFA5adhMlRVIrhbNMv
LDQYJ1J35PHVd0PW6d9Zkd4RnseLQoks+nA/LH4SmH7mpCaUTNWq+N0vmvjQLO3i
C1CjHfP15pQdC5YDfQU210iL9UaIPG1A4BKXBUz0RMyEiwFMqiCpAWlVaXb+U0zX
l2jc2IQbYrkYybT28xOq1wGsIq1vabhrigdz6rBj9OnIFBUip7SU8hg3+gxANfWl
LztSd3xrhrI22Tigdpz9111ajzXUQ6s3cmxTjWit/MZBnqS/PRW1eL2X6/eyRfsu
sOQT/sUJ27Eo0vtuWkNQP8xDs+gMvcy3ZVJ4LeToyFTRJ7ropyvDSCsfCeA6T+9q
SQWUAdqqxVuHni6HXYotA4yJ5ANCPxEWBqzLjsvKlOgo8VqzWqbpKj4VjE2qp4Lf
uyEY7w6OsyT2xA0SZcaHYCn1Gngg4PyTJZxRa/FYwUdF4zb3Q2KIyICaHayXql0e
8LSucC3FZA8JDtwDMg1UumQs9lAEQboeQQrp3clvm0Ib1y2Ex0HR7kPmYWdnAac4
QXcfyhyAHjHeOTDs0J1blb6cdfXGAzDgjokBL//xTHjRG3L24I8/AvD54CxKutSq
oMVeaqDa03G4VdjunCam14P7lcEMI/v+w9E8mQqjMjLS0BNYTqnRhNrHDXlURuCT
Sob8aUTAuFQ2EulYVOlj1Ck71ACesJ5/LCc2e9L5SOHDIrAw8yb4m9X6VcW6Ivgq
V9JLYDTTi2IOBT55PZX8R/J0k4nEm8g9pCz5unT3eNu3//SGBxWlawpeiy8eLBJh
XvrsDq8lMUQTvwnlQkwOfSHdWVLblh4oaHwLABVnf8r3eGWHY403iyPOI6/gzIKp
jTaEGZ5MX8hh+OHUnyzeKLWAlGuvKpZo6+JTKqrOcX/QE9J8lO0WQulCZtbv7tCd
sbEAcrzGA44jX8mPvD/X6qOOYR1lT/W7PfurKYXr0CLiM/TLYNzvNYaGBcP6YFLd
7H7oD2bnKRY3QZigGylROnr1FyQD/3jItjgjt3/5GETH9X6kRSK/Ypk7yW5kq84R
R7sajIHBlBtKAIZq/Pm3+trq9joBpjAFH8QMNWQeNrt17+sbX+re+fjWqESnwqOB
DeHFl0HlWWV+Ku1ACotigZcw2EJh5ipxPaoY6hjzSKDyP8yR5WNvOVUMgs3gpZNE
jB7OwRkNIy+V9jT5fdwvLFpJYh/+/Zr+kxrLEuW4ik2EAG7BoQdITKoEaxnlLPBt
TtCJ02Y8nRONrZkOI8yUDLVZbIG152swsR0gXIn/RDm91pMNeRLgGQtIulcl4s6u
S+TllXALcUOYHPWPYOC6kDIXjTl6H6Z/4hO0+ZNsIj2wiFEwae9X6SjgJYU+0vpr
5dsVTGqgm+QnmUCDMZrIzCo/38w+4vax0PLrMpuo1lHFExgQ7QwOTm2bGEcuDKlG
ivTHx55eYBoImqpiAPzFBRfxNnSVY4euZwOmYun+89dXH7jxdUwMa7yypgqaDn1c
rGr3Y5y15PNiZCLcYdWFNU+Km03YYC2p3BxsBF15qpbJK1lKYjJWzHUXU8yA1bKw
4XsV+VbhdJTrjhkMt4w5d0UScjXGLbtAVWhtKCkT1Qtb9w8aCf9hMGs9fH1g/0WS
i+vyYnKOqVHXyvkgGBgxGRirSetSWnBwzdJoxqRgFYZ0U7gyIuiqB/M/HcrillBE
9D62rcWL64PNqCb57tKxcyXn32nma0wngKOYj20xJh+S1KF1/jGg3DVzy+Z04EBA
a34ycYkirFXNXpqwKjFWjFEoMeNWxjsELLYu7iCoH80Ofz9I08LY2rec0wB/hg5r
zKQKIJaJWbUT48gBhMVA8+bqjVeM9WX2Lpis9a3rHOEolelK7odZxqHJHMpTEZr0
ia/oJEa8oi7HAbJbfjNEtbG/guYpQTsbe6on6+sH5AI1HzaU8TSL+FUjoWWgLGOU
Eal38mIho98tUKheZ7BBl+S/WW3psEKFGyB8T5+OJTYxAlXmcfEP6y/nlmOmCjjU
z/OsRtdJ1mNd7iOz3QZQgyh6oIk8UuqNDAmkghnPmzjV1yEl7v3bQHXNxbqofIS/
X/2NZVWWqba2QzNQnAXHAu9wdsCZOmddrjs7fPh7zB0Y4PrT61QIUHkxt5mVmRN3
71GATjPCPOqs0VE+tovfbM+40ernbMy6SDPdEeFAjV8k5JvF6rC417aGBJVQPAQ2
1h1FuUqCFN9AP7VRNlihr9ZAj4bW7LPsoLCk5Jpz483uQkL+2k5tUK2y5TbK/wX4
UQNQq95YwyeB92NgtaY1/Ut4ejZgeJQNuFHHLDOibY4jfiqOhhDiHMR11/pHGtgD
yF0I+dFBTaCJImHQR8QfD9169eYlBBiymjT4Ea5sSzsjOvsrN11XX6Rx7O5zc2PM
6w+ED9ZTkZVxlI+e6uQy61Saf4g515UOg/VCP53i/GVdN1cFVzw1Zhay2LbvWZjG
m+SiHE+pqx9ncua9lPG3JlfJkH6NE2LsxIQvGjTtrbsZ5+38oJvz7+yGmPX60kmR
r861NKsddhASfQwuvmYoOOpXnBs07BFb9h1YeNmA3KIqeybt2kM73CI4icR4MokV
8Q5hp2B2+5lk88aUQc78hqft2iBN87G6WjnF1rlmL7sfADlv+Z6PQr/Z97JORT2H
lExH1yb6HerDozY7MelE1uXw4HCAT7BF218C0nJL43Hp0kMJgFwclWlpYkeKpN6C
N+/pt3XNIIC+1cRMJL95nZ0pqVgB4JCv8h5Ai1lXUweOKPTrVw67JcG75QFjH+ne
gX+3+mYa+Hz/t4duQRKeRsTah1bM0ZU3JUcmUWqgkpSSYQ3M4rSjW3EA03FqB/B+
sY0kfrjV6BK/WUPsrkD+r7nq1qp6iDunJPIdEWwV6mhxk6x/xo784XmZpw3nOzoz
uRDYnpUELY7nlCvtM6FoLEMwVgbI81x0HQTAmVB/I/RB7c1fRST3Y4U+iUwuDQv5
PVVCfRaN6MwlmXu9zA5LWVNz2BlxiVndPDT3C4HMs6aYgiDcHdDlW9cmCaUS8HY+
RZgX9x/7JVC4GuwmLacwCgr8o8OlApapvGGlKE2FPqFSHpRVbTgSkWKc8FUygcq0
V3FWpwQaAaUGzbz9ZCY8zNM2seyV96vYy50lZjW95En5u9Qez4qeBHqH3URXkaTE
9fi+BwEoCu+ys0QNm/DMruPg+E87K6h9Ba9ffTy4fcZ61lMz80JOYyxvVrAMv+kT
qgmyvGnAGwizXCYNxFee/P5kdBva8bGDb9ffhcervhzU38SS+6i4X4arWMR7i9hh
uG8xy0etIViXIbAZwplKMnq4DHVRs5FBBRkV+BEbM67RrXknavR+PLYpwxifjEuq
LvDCpAK+K+JCFXduK/UlH9xgBPxl8xNoPin/U3cf1G4zR+lg5z5ivSqMRdLhG1Jy
KozYjDHZkkY6qj33dH1Qx9uNh+3oNvJL2mxPAFWJ/+bObLG77963/oAFT9v6nWqq
XmwhWWAHq9v+RHbc/UXXQNplY2SM0I+8Gsw5KxPv9/LgswRoMif557/F5PgmrXGp
qYzLyODuLJ3cCbXkt7Jemb89sTwZ4oX/7eMN1bba4bDor+vGhsudl+3l5QjDcTZC
bPKPzOhWLPv0dZdqtQtAbk5E/4yD+pnrom7c3NUwW1tSu3K163Z8wqEcDBoitF23
7r6ltk1KrJIMrIsTSfjunbD6P589Oe/X2vuY9xabrMrbiV7TRowqMD3lq508mB3e
c05369wd7JfX2uz+5dijbC9ZMhIOFWnAWCT4iZQUSJHjNKQdTz9iNsgM4wOMnwlj
c8aP9Zf8O7dR7cM1DTEzG+nFdxdDTJiPIG9VUyacA2OkcMA6vDjRJILdkdjsPJZ1
m0Xw46xVWDIY1VGn3vBVkAogEncMHnv604CMoIMGyZBmWF7zd95VPy0O2fCoMr5s
RL1U5iVE2KV0TnKwjIvPFwWpplG0s/4dl4FCgdcBc7bJrRQD9KCUJF+o5ivLxA7q
aYDAe9R9pE+6LdifodAXcF6A/rzfAfeMC82g5dwxmFNyk1EkZu8Vnyx4kJAfg3M3
9k3aslqaKwYnR5z30fJEB2FMfRBpjjndK6AMSoWDfcXbhP/xhJlJjNpi6n5xXqH+
PYkQersuaBFVtMZnSCVrHqsyONQwMuSoQNRtvLZUCzfGTMAxmibajtF/3WuehMhQ
VGybd9mfN8nRjGSqMcoMncoJHHlk7jjDLp2vhcEExLq/etymfvcOIaDWf+TIrdWb
fX6x9OMlY0QyCT9UFjjHqSJMMkBvguiPPGWGdxyXEtfseNK+N/W0zroB2B7ByH8D
lEBOZAdy65dignWFuHzrAwrlNJvnVvRVtcxXSQfuKHNGjuo6sB+v3vuhY8jIqFa7
Jw+2Kapb8A0/xaXtATL+Q6+B1fwltSrx83Vq2fKd1meH5bCVqmjie9xwgmARHO8W
ti1u8fodtLM/jnwup5omgNIrDkz3uZ8nIJ37gJAF740jOoB6tD2Xu7dpSrdlvDlu
JxEubPwFEVp4tVwvHQ2VWKg301lQdRP2Nyfb14rKnEoDczEOpkCIA/wxzbKdosdn
ujBJ/M6HUOWsc/ZdZJuxGPYkBI99+tAwel1R4ZHNTmG8Kqh1C87pzWn3kjD9SPKx
jRwPFVNiAu7RXrBg4E8q3fHQVFQPVzCTZBN9QnFYxyn7AUlrM7HohKSQVpQjruOx
ZYKdrvOrQ2GdEl2JpVGFwFcR2DV0kuPdzFgfl2ERZCsF2fD+y+izUV+pxgys04UM
9bnzc1lyQ0f/7upWIgNnJcvY/lD4OFFPqNwysE5BfqBvRsnovuntgbN1rUzfub2f
TRfkVylwNUO4p3DxV5QQcPJM3pZ5nFQe1c9Q8f1jb8x9e9xUVx2cPWL1yFna6ioS
4L+bJKMKXoNx1cDoAITJ06Kw933p8SlJSz1vPcwH20uWUzqn0UWrcdZkHmYDrEFe
bhlornNRlroeg1WEkd42f0FUqOdOPhuWAoX48psQ6fKVS8nnWX0zErG26ENbu1Km
oHlaD3gp3LjQrM2ZOSWkw6dCl8f4XrE4EC/6GmJQfT1OutEaoMSbepbu6Q/7mEP7
cjQGGbXjnABb0EsybTK3tCT87l0/WmaXD1cWEX7QfJsK2olOqGxIjeJMzE1k5vpj
P35mcCa1HNqcFkb3hPu0vciPCevWAXiOCF/IO/zzCpNjooPTcgTqAHb0IoUoECdP
SmXKGZv2ZCArupJsoUprz3y7iI/1NCW8CU2vNoBNF2i3DSm8NxZ1lnddr8hcxFez
E6ggITAASB0Dkg/i9uDPCLRFiaiwVFkAse93IVz4HOHRoBaJKa+SH3l2udj8ysY2
rLkKR7ukoI/fQTHRBTNLBgeDyWKUoikww6TRnkHGj2zvOZkN6l6+lqaaivIywPGA
9KW1UrzlxsuVNOTqPp+pzTPADxcL4ZlF+V0zkt4rOLk8ImZq3CI3BtuEox7XN940
ClgMktLUpjXdBbM1CrH7F43jSc9RLT9bzDod9BxLA9VtDsR/rub1Dm8D6dhDJVT0
398A16Fg4v+CMZi7rFinIoUEju3NWPy7bFTwVC//70bwvM4YAsCQqUHTSz3Y2qw5
p1aqsjJ2adM0iEFl2hu+qjOhIAUBXNeNAqPitzjrohZV9Jlg/5gw6MEtm38vp342
bM/lPgaXN1A1mB/YKmXCq9u77BXYimu8/uFC2b/0CNUm3M0YpaUJRsV+rgMGOz/S
TkH2Ao/3N2hU29ZJ3IRRGBv8hUcTWYx6GIUeqO6PaG7Ka9av/MYVIfZdten2Sh3j
nu0fgrd9ROzw1xujV+YOp93XV3woHgcROlYYLJqbWbCwWARLP/znOqvGoK08Af1K
KwfhflOfhOEz2UIsRvDBZm7TH1M2fup5/yUXUSQrHZ9hRVz+1f/hixKEqfzvYY5d
ixu0LOOmIKHzD7/Ns04EVZhXd7cYAX2rL0AqetPJ7LNls95mtRb/tjYwDJgOQpib
EAurs1NcGtLGSLhFD/pQTRZONZU7jk6H9X39/15t8f1wFPZbGzEneWPwt+hL+lDD
0p3TBd9tGQtlNTxvYlV9Pig9EqqK1TdsWdYePIs5O0vAee2SO3u/TctXDGOWf9jY
j1So8dJApkaqViOOygDm/HdDPZiUEmebQnRYW7XLHl3OB4PqvCl18y/Lhu5e/4DV
51wTYM9mBXX2yIqzCpmMpGCFusgKpFIgt+0oNX3GhiTtDPHpKLmCAp8wbot7Xf6A
HmXJJuCrJXpBCGsQOk2j5weePlb8G2S2xc26tnnd0MWvxlFiFlCVjcChLeyCegsU
I1GesjlveKcjakQsDsqajBLDvKy/RCJM89lvbcniWVGt5OlnxrW5INxy7Au42f8I
khhzeKlSifOgUQcO8nUGFEBYYvVYNyVAW7gZs8KbrWf8zVwwAqqALsyv5KZROgFC
xsJwYa7Gbr5fQjViGnw/pu39+Y9QNv1JLUgOPSHWxSLdWlsTQN5wJzabGCCGdQ54
oBq4ZedlsgP/Q/8M5SxHp/ArFUppBpckrz3PHLksnNP9hFDgDrnDxzLH/qC/TDKT
O+R1kaI21hx+kkQbESqYMeQSDrQgZof5h8iw6UJ/DFEP6wlfsGByFB+t0q1e9Egv
2aCDW7W0bDTPDn0lLHx8C6E4jIlOL0n1ZvaATFdP+NE0VxncZ86NlTA9xlo6BXdW
rbyDsNK64+F1Y5NbPRb3mCm3d3fYbhiCQqgPgTAKNA2llikpoGvFA2xQHI4YymvL
kEEV4ST6hiUlPiyrySbIhORD4rsZ0lL+Xb4jcj36ltYmIkEdpAGKaDiGTdSit6a4
tDiRx27+0mXZcDJyAhvDI1VzOAIQp/kXKtsx6JHLaiQ8hFXUY8UkaYTstvvsqiNY
BRddbWXCfwLwZDL/py42satunYUjnUYvKYiNTWJZ5jEos1qCtFxznOagne9V6DcZ
yRvIimRB78uqexiUUqSHXVKZo2LDJVC12k6/W1C/oU+Lxp8v6JE6MKQRXB/2Lx2t
7KtGfVc7XwdqjzSeRjt4CUpK1w2nKxbf2caDXHGS3brQ49LvY7L1T9L30qeFJyqK
0LG3lDPUF/i06ZBiEdrSHdgrCkNNVZa5xLcvZ/GhJHoyIG8Jsf4n/fbi4zP+p+wz
UFIdgrVYbEY/jJV2VStjM7kYdfdkulwd2zYcwIZnIVWV9XarwopvvJyE/1P4yb80
UzIU12KEeN/Q7UQgrtniDwC9g4vGp5E2OS5Ikg8nO122vo/h4aHFZvIGTcfn33lA
EjUQv0SDzcJdU4VJ6AZWI2dZDWN/lT32mV8HAl3l3K21+XSpgi/cWslxxW01zkG6
ZEy03ZFVk8WNhLLc6CMw8ntlt73p3W59OXRPw3IbKUVN9xTBKaKAePXT3Mp56lcc
d3M97JExUVsmWsiTNmpEtr7L82NrCCAoB1maIRRh/Ybd6DMa5pLTDNk+P6sUspAd
aJGV5OIS24RGhnnARNJdl1wkltIz5RZ0RTx+CS4V/k8BZhWA7pp6sU/PMlUxHOVi
OSElwwVEtMi6bZH+zk3SeubHrGzCyaCNxjT19LZNcxlBvaT6G1l29Z9aW76zjrBr
551yGTSN8U5XR7hr1e+2ExL6AVtiClVZB0vX/QHDdu1NIueZYDYQNZb9+ULeFQYK
rVA57yA8nIwmZSVEjV15Xn59l45mqPGu5DZMiEh/uFcw+25qDnnn4nACFpXAKkJx
8TWt/l9epU20MC5Det+LKVT8vx/cXpLQUg/radg+TSR5zvDJGr6SCIoVLXfG71w9
D+Y6YbjVRdboSuVaruKK+BYMaFX16hxLTxzP4VZK6Ni7Q0d8AOCmz9XYBpohZM14
5WZ2IrIOq1jK/wZt3JAGKRAC+DqD1xFMLeLnVqBaJY4qK711fH9XkCPqpQL6MmO5
WiSeEsxAkEZphPm0r/NaYh9eGp9Px8Hgf8Uft4UBTDWtqiBne4tSs2XlH8tBcIru
/poZop06xmHHiA+IACRD+ECQ4XEaMJcpyUpFelziokgSlBlGXJdTOz0PDlorDPXd
+WVQWFpyTLbw1WJKiXVT4JSZLy4MAyt3Ty+hoiLloWWaA5O1oeLCGpw+ct39YhZH
gjuKzFgqb0iNnQOqrwUhLb2UyHkNF3t1MaUS1nJy31Ye0JPYRWVkQbhgTycFYi5R
lQy24txuIOcYvUhOwilM0BpiGZUr7KlnGFHb2HUKgjh0PffSiMo27Euuki5N8/5R
iBS+tIVh2SVSKsAeYA70+QZnUCy8E3udSzzDfq+xA8wZkr+dhJ7a7htXiihy12o8
XVemGZ77PSNjpdpoXzHpH5x4JV6Jjj413ZD9eynNXbj+cUgbZJiyn/tHBG/t75ej
+rRRyPakhKlKa14cFjM5a3JxcSil3uLmndmm/I8oSzeyJIPmxUKBvtn2yhGGYjye
X6UxCKAMOaQFCuA/h0pn9nprIFRAz32Si8DlsfzSADraugGE0qnay5C6YX28S+fr
kc6KMfe/KRIZYYtXDNsQBvZEyUprYKnjavSKRe50oUa++NuEVbua6M3aEfVJXgrG
RJKxFtQNwtGMTAZVZKczuDjZOv/LWXWEiQZgkeTh6//ItteK0AzOEwJVm5hXTmGp
vC8oWMOanvBe+NN4gtspqmTkJ05WiP2PYBUYAH81mxAJHro2wfLO9bkuc6kWUfAv
mAc/35wSeVeSwH4oN1uVEzoMYTybEllfUZeqxfxYC3K8wRAcPfNKdBqXx6zXHLnd
xSMoJ2L59e26zN/jAtzBQjedisax7EtAlNXWmw5TUVtYloQr1Nw6sexxT/3/bO6o
BDaM4GOI3RFR8iv0HcRWV/IoAvg6iSB0wQsM1BZq9nXm0ArwWSwLV2Itqm5LA4hN
NWS+GEhTRZWAm/ieOsPslBy1H3yW+TDen/m4RB6MGC3D++m06UeKpSkt6n/98tkY
MAP217Joj/j+aW+PObuEbLLkteEoHY+btbX2eEAWCmz4jgoGzUbmHbm9yvgBiQ+C
6rAZw/XiZMYIy4DlDh6cfefAxtCuFB+503BeXjpmG8BHOqFH/L+s63FDQgGDX5zX
d/zU5BaKCpldfBAdrB7TH7XVnp17ImFKVETF4QFTc8VnamJC99AuGC3yGa0W1fAE
jZBL1p0yQjyJOC5e4/oYaOeU0L9GaR+AnpT5fUdlBfTY6DK2lKGyw9WfVJUyAMFT
Zzx7Y4YWD8ODDvbT2Obl2ZPF6xlGvENPr09evFiLsGVWAVFGPmWUq46oIus4dG1B
tMYhseII2pdQ2bgWSiXKNbPceN2ocKCm7hhAjxi6RYWqPSlCdghCzKt60oosvs+M
Xv0Ko/8gpvIRxQArOvpFY4/SXG+ol8qknW95RNU+BVXhMNj5gu+1eudCFjoQKWD4
g/haLtW72L26orhqSg6o5rY2DfJD+fEutEPymd1nCaIaAYcI7w4M2BN7zDeQOTV5
A9dpS6a8O3FCd93/o3JzQhsyALPVBkN1l5/M2uPP0WZQXYGJIO9ND1BVq1lUwJIp
cr7cQzmQHggYLpvX40JUW6tsebVX//IDTNs16gDKiG9qIexN/+IECAwYhS5JINy6
r+TfIgehSq7bhxYX3i8N+uuT5ujM50tsv72Y4Tk3sH3xYc1NLeXKaYt1pfzfFnGq
hzf/Lyx4obgSrgNA78XElAAAiD7dFTTxk+SUmZFXBJZFxW50q/LIIN7DuATZJG7H
vtgljXAnOzSnWQhsXyXovYllhImqT1O7WnU7eH058jxJRYGLOPO+U5zehY9NfARS
w7DimK15M3DNka+6qBFmlwDegw6Ytk4VSu836v4NpjuzyVGtQP+kvn7xizoP5KV3
xr3OIDbbMVHH+FRb70B1gKtppq2CBC5DFgOVhnWj7g0UJqQIoBQZThQ3AcKxHOCd
H2jf7K9h4BefzseLp0WKhf6gJ3XBpet+ETmFlxppGHKA2wR1RhuIlQ/IRgCAssVA
Jgxk0NGKxX1kQinVxnou1MNDclC8q/vl+A/0Efynp2NW/wf8WdzD+S/5e8xqqTDu
s7aMyqelwGq8HoeonQskJ28aZ2j1Vf+lxGlPz4WtsjvyoScrgiboIqGc8yitt3kL
Fim35Nx7mXvn3t9K9RF6ifzZU2F7AbnoQ8MJY4wJISKNrBw3UcdlkskhBJc9d097
9ZVDcqgXFE0vj/z9bRZpQ9tCerTYcsIS9g6JvKUf5brPmZg8hTLSlV9O4RpjUK72
4kvYciblFCIpO3CHVNRcEma5ORCZj+EVSFhAPPoGWTUdoUigyESdx6uEDPqmzPon
1MpvKsfZ0RrJ+/e0wLpTOBHYPBgg4NbMC59+78vGLYb88oXkf27iGyRy8G9pHR1B
bC2MhHJNM0GBDPutaKJVXgPNGIZTPTgiIqFyLQT8fQcMmkJDj83P6VnyzBMh9pOO
sI1SKaEsCfDW2UibzlfEIdAzl461YPS1T2SlDHqNiCwlHIUIscwUtnjm2qfWmjA8
cxu2QFn4SYvAbJyco9KTNz1G7TDDtcwYoM1vJDvQ4Nb9Vy5iRM6gd7X0VCZbzUCK
8uyJldO+CxX597/sK2tq2wnOgceqv5fyi078z1cSFoDwCVWYCg68sR/PmfH12t41
fCMZoK1JOk2cvFGppRBZhcFPtrXWLiYGmNJlr1t2U01iVJ8tVLZM/65OXhWK/6VE
ceR08QABI02C4s0a8Q+3AV4iLLIT4oQQRv7hiRr5ZSm4f/LsTwH5/cjLKrH0lQOH
/wSX+RcnACjEo6kNSpGAAjUNYMkho/CmWUatWgHq7Imh0bI2Fnl8QpNkbE4XgEu0
srRTlAITcGleeJqfXhBBdWCLcEH+LZx96l0z3LeWvmtG9uUxo8ZUhrwM0OPxSNmq
/bbm1XCwEvNEXyBgNgZBvhv9W1/Dv5QO4D/VfKI1x0EZ6gUWM6l0r1lqbThU/C+x
5AZ0vToHSqch6xM6OV9vghu0L281as/i7+pad7rDU86rDH3pocXAbHOqco71fh/p
YzCqzSSlEx7sisHUPGqrBbrZRq4NaZyZW6YNC3IIqXwCtXLgjm7JT1Louf6RqFbw
SyS1q57knxkum6FZDjSyunezs0XzKDlZMQzRCG6ut4pi2YObzMLLQcqgffPRgxAh
fKg81Pqun0fpNk3n8sjqlldpOiox5FVmEQMXpGcS2D/6rRiUyb4XU6bJ7HE11Huy
hrWGhJl9iWkeZnN4pEWPfgbGpv1h4exxFh9P5kmwFF9OfFq/afyrInyV+CStY7eL
yC4lLAi1hIkLr708mMfn4WFFmMgejuAj4lJJw6jyhHjTuqZHnBpw9Qn28VBbgTIk
jKKdeQ/2lDCbhSxRh6sSJ4LHVm3+kCXVgIa3n5kq53+VagnoT3gCaaRysJgBp6m6
Sutiz+bHx0s2OEuvH78jv6m+bftJgFAYqL50ziM5fAR6qqjaXm4WJcqjYgSgHWj8
QV1PQyja7K8aMNKGop0HpM6cL1DQKSstWK1zcnYqEKwlet0kyof7wY3SYldQBn1d
rKIsftvP0mJp7nciS41Iw4b0odqafzgbQgdplcmC8n6BnWdQrpaI+ohYNbtH7cZc
rkPMMTYV/+iQPjWHhMvIBJ9tTKLUBfcByin7qhMS7ufIGZ41JSe7zXGvb9nl8J2u
r6ffg5Uu2lVtMde/WXaSoLDxVGewvwEutZbcNqxBOBXXNxGBjOBcyE5LqRHICyyQ
RdcENdDg6BOeUk5oqg9T2SD5n6HYb88A4YZyTtOhY7BHTKV2dTBTE+5XkmHhjuvA
DEPqqEPHatdmGzdp0rtFNErHbKVdycAOJjUHp55ZW/ryQrs+R4sPZkgvwdZH5tAu
d47Q985KD0pSGV4gok9VVYs+piUudgthujQR1UmHnbYb0+Gj9eQZ9Nmb0e5Ppbgn
HxzF4E7Ca2/uJJU6sUCDq8kmQX+B5s1nVyP8P4NoiO3j3D5xI37mkWM6Odf/5MSp
v2SBB1WhACFM/Vh6+ceKB257UwL0qPdrFqchQGcfF3gmEjhf54lR2O1DM0iPp8Yj
u3uB/nKEafT0GVgw6QCZSzowphcoPQoa6UWxI4wd5/kKhi//1pSUbriWlBxKKWUb
NGeSotOKpyvNabwM0mXmY/1EjJkftPNC/jWlgfAhIwhwc+MuyFoEJyetqf8gDEl1
nEhAQMI3x4umHRBicfK0exyM1G8yE4mKWkLj3nWl0cjFV9gTfv9hZEikLHAMoJjZ
I4OH2HTO/f8JyNy+xvA20GJG0vL80G+sPJOLJTYW3v7jDg0CX96wPKebX0U7mbx8
1Vnb3c4VPpbJI1FJ7BjbBifSWG6zba+WxmHD3/jIi1vyL/VyQMDJWQHjfySGUT8t
9NWFavVLXAyUG2RMSNXiKAVQ0LU66i1J4MqayRa1kKXNxa35Ey7i6keCkjDa1g+S
81OjwK9mPi3zqBsPinSotcQMbBduBfFF5+I8/QBcB6SHoNYUHiE9eI2wT8PMljAs
7vVAbOsvSmwxiyzsTm25WuCJavvtxEN1GM9OzlX3egzPPjf8YqcLcNTDegSjX5Xp
56tcuf8wG+rAU95jh7MCOoQk0RNv0CXikSW/RrXGJyWakQ4VPQf4XRDYPsdfzHeN
jmbLEe8SI7YNV61JAdlIicxp3jMS0KVwO4IOTP6XH3fI79bp/6JZMMwCj0gl5FKW
aRHXbTdbugRJup9U42mlGB0QmAWBgsqT2A5bB1XkeU9utn0I7tGptyK18Vqro9ke
OTN5jPVR2c7Dqnzn51p6UVi4qMSeN95zg/dVUu9N+wZYoZFn+4P6uDK/zLb8L73S
wujhrAxqKFhKHML00xWKeO7LY7csxv+sM4G00PsRop5xyjsLY34pnxhAOR5Az9Ao
p7wFhFK7GuI4wIAPlwBW3SzixVxDuRYG7FUD8Lx1Aa94LlYDSEpzaOXRPRb49MtB
uMvPfLnn2GX2gPuZpZc5ArRSbQI5kDUQ5ZFgi4cXXAFl0+65YmmCG2R+9O9t3dCn
cn7VrFUoJSV+DeEu+es6XlQMWpXSyfp+bSgdDx7Tp2wweR6IvvzGZX3Lbe/Te6OK
nwE66o4/vfvkoBt/HmsW4+osXVKw2GQbuzjy/Ce38LOIN5EBZzHLnFSQOfGfhWFg
eJVitui9ayFN1kTN/RHBS/86Pp3N3PMfwRFjIDl55gCS2EZVIBgx40hDu0U4ZtLj
f5W06Q/hffIK+c8HSE99cGhm/vfg9h1YK+6wHsT4kEcLgbG3huSmtnXAUBjmX5Wd
pBmEDc007e0lNBngCCIswi0kTSykPeH66D63rOiGL7jmt0XZq2UmAtH+WisVAFfc
DYqLqiIyCahDvRpGVDJAQNSbxmf8pVfvJR/PRezhJEqgT0XWQDt0BULNYCBwbAKb
jZiMsekh70FrjBfZGRNoRlLbioQoI3JrVSGlC1B5yBTjwDyjE35G2Ndlv4TyFCdN
aquFdNJ/4hBe9Xkua//KskDLdSgOaehwHFxHfsE+oO4VGuDtkmS+cr9vgzUBNyaG
0L7tQS8XmAX4C/IgKfICcqPfA+qzNaDHe+1I00G0p996bjb7aFRw4v74fopVrmgs
uAy77Y+PY75xq4weD/9FDrl1+MWpmft7Qh8HBDfueSzjLwuGjtgKXKf6LC9HHyEb
cQAzalbV5GFHiw1MBVazuBW4otgHjvUf0j45TWj17F8HNjX/ZyhWwnbrM1h5eyha
8s21K097g5y/UPyg3O2brrnvEXs5GG+Nw1M5qehUsA/LzMbOws3G9X+oWAhkYJ8h
qi2qNAubfc4ZPkocF2sqfdntNL55k1EmtsdGcX2lIGaG2I5OpRFLk9qm0S3zszin
LwOh80szlbj0fhfuTZVejKVdu90eKDKiAGKpRVXM2tMY+kdRJv3SFRH1xPNbmr8q
VmiOj48sTksbyXoos9M6/HGz/UDPDdm+BTqEcwGlQEqDMTTT/xIUW59tHozCv3iA
JBcq69EEo1V/SIvWixVnHV3wPJIfcM9MWQIKWiw1Eh+i4pqqsfP9SG0XAKyMaUZe
iXnfvHE5WObhrXNBuFDKrzMcTLiloQrWP/ac+DO1OlZWqJuocNXNgeKKL767IsRj
Nh6Xqfvg56fVAPOWl5DMf18//xoda1zyRUxnbhZEALjSdCR8LhxIjAJN0tRw1ruO
PQ/93v1YctzFva8c+vUGC+KyrAnOoAkDP+QWMHoTdOUK17cKWtmEXPtG4Dr/Yd2B
17GI8+kpKFlcZOBdnG+QAQpUgmTzo4SGlDSG+a6iVu2ofdwD4tPsyM33fy5UL19+
vfRnrzznfBhiEh3BunFdYA6olpnYAWN3JBIvUwucN7ah1L5LAHq5LuLw+Ncz54hA
MZE9WmHLfkDXFjcIGvFvZdhdfMgixLvmBz+Wm26cFlWeqZYpHkxW9zK9VPO5oFtU
i+trUUIoy1XznjP9ZFc5x9Ee9u/WL/09fT0DjSOcWBN1vwSD5TbTPHHyCFiRwXMD
c1XCZI+Zo8w8CmbljoQmU8oGeJ4cPagFygETsTDXBizJG7q8R5bzwp8GSV1UIIfn
pUcXcFHtME+cTStA55f2xd9WFBHEY/mIY8x3kU5fneSKNMtWbXwbqtYJLYIXvMlF
tqlZMJ9LTlkK5XrJRZBifPFcrKYMbH/RgJmJ9UghgKrh3Z6At2wZKYbN+P1ENKmi
dBct61/R//2TB7ihUqL7C7BWm+etJrp1LF48pTH3owBW9j+YcFykExrOIYiGXHlP
Tr91YqcqjBq/Rm+qY2L+ELbb9JBfvqkyQgkW7CE5CsuU/ftZDP/NUtfT94IcwUJA
tGFW9eeAL5UWZvT1KqvnDDqucjI5dFaEH9td2dmsgcVJq0hCeHcVTnRXR4mvLY8r
rFs5wtPI0ZSPOw60kn8WEDyiyToklBKB7ZDdcXBqQ1mZUerZvCvkXW5RBu1ktAH0
O8gwuntuC/lILxz6SY1BAVXKlkoS71wCmdE4g/4odKjMr9bQeQQjw9DJtM4XsdJN
pyW7B+9tB/nP0j4GDmJdoSgDezqp+cfZ3m7en4w4F3h4BukjZH5c/fFFJhV0x27o
9HC2/Sgb3zpghIkJzXSxlU48q998EmcPEjhFWgTgFQpgRwt0wa8hRcXusO6brSB8
ImiV9CLvq6FFcqQsarp21iG9B5cpENkGEAJ9wcmTpcec7plGabs+4ua1sL8cNB99
YOztq4eGIumRIQkbITh+ZYou5rWXz8CMjQ57Y2BjN/7QfeWLezw6+vDdGWdT7WZo
vHEFfD5Sh0GmfEcKUtlUKooQ5zDY121nKcO+4x6WPm2yKS+ybD55qpGwa48XOOIB
TKWb4xr3b0BYEpGaFa0sF5ZZsPB9aJwtWNeDGlXPZixiId0o1pJQlAvZhX/bsB7Q
HfXfZEXgvBuqlovjmVcYTDAeSvOGp/+PqD7xP58UPfmiYGrQ3leAsobjvuFFHhTq
Slievwz6FHowXOTQx7LiEPpQnb2O49oslFFiiZkRZ5vX0khBPDUSbWcNTC2wtEHA
hy/9lhXzjouXzBUtIBcPdhqnFZc0iKFBFSnyXMRADYePNGY//ugieqK9Oke0e8hk
jeBqQzGvlVP4h8c0jxqHQbwN4oGSbBYbDXW90Cv0fe1UMs+8QZmkkFd4i02WV9gJ
HnWJ2UY/+ZxEZABxwAYFwMAi0WoqkPIr2mw/Tntz8UTxjHt4qgZTqeTh6PNF0sId
4mAQf/zipC840ht2xQ0lOukY+0XkiPgk2e6gAmU2/vx9ncRt0MT70AX8xuBV5iXc
DeehHWwzWGDF6W0IVTJyBPNeVaHNkv8CldXFuEzxWlv4fhsHdwjwsyM/d8emE1lj
2R94yeMGqpDqU892BN63SlSRSQn197cU++gW1DzZVr595pR0yqJb6sEkqrA0Z8X4
2Lci/qVFUCMtUIbHn0h/lT55gNoVux2c2LmtH41PUYfjvT+EKGi7cNfkubpdrdaG
L6/+Kmcf1354qrvSpNmR8msvAYgAyFv2E8y0jMlqURYz2XLsuYXhPY8LhG5Bcu1M
rTJjbFxDAnYNwODUubIzTiq5hxPGInB/hasgfSYhE+8FtsDzmsNSPIl+aoyfVGV3
eIvsYMqXkNtLpWwcoVeHY/0CilOD5BGNZULmjHg+1O7R/e1V6zyZjix3WT9p04RT
mT/qU/fx/GD5uyHamiLTbzct7kuHxJNXs4Dfq+8+Qcg3WydszOeQ/dUI+deTPXuC
ietQRaYSs4loihNI+OKfTACpa0Suapl/4oLO11tvY0yRieBd+IhkhgbXDQn+808B
oTcHLMceSbPuEbBLSmcX83KwIhyIWIKLdZBTBjNlmw6VVyf0mbiWg02ts7jnPBFF
VdCFHtedAF8AKXlMtH+XZn0kQeUIk19fUWe7gh7BjX/gRiIoJLzdvzHyaCe4yemY
VVNpTDioqmwrdnyH3HjmbB5A8bytQHzQFIsfLzZSteFd+Wato4r0h3kSDfYR/vqs
OEFTf08kgbiQkgay4wffnLDfkHuwKsdQVRrGquZkwkrDF7PHwpNpvJ8KerH2g/NO
glG1+v2vB6sWLYvZS/HEEnAvRn5D4vtgii+UAu7hulFj3fFZ15TJSSdyjN6wK6tM
mMCzDmsK6n/be666+p85pLlsNO2Fzd0VFPFrpZOPTqLnlHfJ3ZGos9QM17ka/M7A
9qbai5HZJKJWADdm/Aztu4U68ZpYVp8ShF6KPlLruBSOk/x/gWftV6oXabBBlloo
MXg76rbrutsvFDPVv//RGIlIdcItc1G3FBi/eOJwkr3HAYMjXztP2raCqzljKCRs
TbLd1yqERfP53FRv4nV2EOvN+CyyuG1qn2qcZpzYvcKc5Dsvp8/kc5tXoyavRyQp
kgMBKUw1UT5xVKeW1BXJOI/5fCt5n/L7ElNlBFV8sq/NUz2B6u4dVf88reQ/3f6D
OLbSQSK0KC10QUuZeGFaUyDHiq3467mKtKFFh00mVYbIqr2ktKQhMB6rVloOFvwD
kzSFkrmYNCNE7/sYFfBv9ftw4PXL6h+2/h8PqFpfLgbSdIKM6vc3qJTn9IlphKIk
lp3MB6YiOnxyINQM9BDEEuEIBp2y+PS04cXMJ7hzcfotClQs/Cusj8KfSABt9x2/
2sPb07LGiEDRjGx/YQ2w9TxX0Lj9aEQB3V8EeU9/zQv3DXkhDzjoQPAjTePr3Owe
AszdMyPA1YN7SJj3c5TM5nM/mBCQDGx6L6a57OAjCJBPtuo8CA7Lc0kTZjAJ5Oq7
Ca/VF0eDSJqdp7En9loHIVbkV9IljTBLwdhDhr1dVicuPbWjSZTugkexAkQRx4+2
1cvzp2ZeKFjiexsZp71CKCsOcWlw8B1AEoI4pAtLsZF8sYq7WM0xi7shm0j09Cg7
vMzv+kf4IGM8G8yxuxWrcKYTNFq2xL3VncXwqgkmHKWMlvFGUloZMlD8F2ok6zPG
4gnL9cWvGqqhlDTtBkO+HDWAsXll92agXTncYq8km4H7NHdPnP7MIthZEOTEbqo+
w8KZIPzPPBEj3Xn9VhPbsNaR6NsWIRt6kH1LZXkLIclWkdRCrGuImw53XRngCpcP
ZnZm9vY3FDjsCz0RGt5DpQEH930UeTtReQ2qLJ5iR7dbr2qsicVQzyQkP+QFPbKH
ylY1URyuzlnkkkFZIaMq4KBRUQw/Vx6YznovKhVqiIG3rlIzval80CRibzJ4uMBp
lyyYiqI7TmsQsSyAoT1/6PFgSJqNBiEfgzyf+xx8QJAzycjK8sEdPbL0zUfPx3nn
cVGzhLZLB8n/NLsy4T/FXlZ0usCHGDWBKVFrWBBDd+qux3bCy0PoTErv22KMUNOn
ZZndWOBMPRolwnvV+lYAqOtMOIv2XMFVw6pGS/QHVAE1Qn8yAslUbUS3V0tIxL4c
VDzIfGlemOEr+lOgYpUEB8pvIKyH3ItrhUTd8EUIJAsxb0ZsEgWFhjOmc2Ht3NN1
2fcsqYm2PnPmbBjwZTguimwHWFtGJRLqYMk21WkudqR90daa1sBJPRCiQ1vOLcOE
UohIx7ywf93rZ9NAc11kpQUwXqkStKvymxHtxyMBkhe7jZgOixof7Tuz89ho0DeT
ca14loY7clhJNVJrEGx1ZI2HiPflmIlSaaczZr7ZAGvTOe8Wribi9UpGmLJ9OfOy
C0r+/AcjCoBYRSxoP7xU5RqCo+ZEZWMJG0w4tSl8BG07zvd0IhDaqEtcpCq0+Xdx
3JxhvsAea/ExS5+nJ+G0UsXhwyJdB3K5X3iDIZZxuCp+F2vutcAyTV4Rsfuw2X/3
drmKcHBVnjtmfelKOphecizP1QTl2WXMGUovDERcrN3RZjZ270H09981UK02ZOYz
ffsXM8ZZcXNwVr9NLSIPaOj9ykPCWVCJ23Q2hGt2ieFdX9zx7oDTcRCEMeOIncbS
u/1Fnl1zxwDtUU0Q8YNaMi4jiQg/htigbv2XRzE4J5D/d/CsfMnX9CfmDVU1lDnY
8lAWqpmsYK4vusWOGyQjbnw9tCS5jbM0t6GKVWh8HaXwP0LAOhrZNbEC4nkDkN1c
bM09iayYyr70+okcPj4G0LLvHESs5mLmmluJuO21nco/16I1Zgk1mqyFIUnU7r1u
SPzpgn1KI68q+gTDt0b7hqbZ68O3EAuKpjs5A8pQvBpkokvLlUXMGx7lKit7YRKU
lq21MLUXxWLkXNGFaSh77udczqIDeOBj+TTg59dnyNFtjQWIyd6k/Y9VZulbvcaV
fHWpBGYmDZgBqJhi2emChvF8Ln71Q/3kFdZ+rI4wjjV+Qb2SWZf9///naDjOtVJZ
8gJqmUGpZc2SzMfxKgk3waOu5KRwTyy4PZ7rxKHL/Dz6EG/CGofttr+2ECyIaQhv
VWusTRaDaBllPceEczSI9ZQhK2rD7GR8O3R7daThzEnHPQoT9TTmjpOaM/o438hz
9Bcwm3JPbiGriWpfvpxs9j25t1iJcXMyXKQ2AcpUkoO5O4KlBW+J2RrEYCI4gcCD
LQXvS0BfwhylK1AvZUf7UzrQrdVZh2/5WebB+Tkvu7V8ool+E9C9vfbYwdtXAe6b
kEgaSUpBiHENQ1+aB/J+VUESaqkFCq3FIGjHyz/aYf0/ugxVkhtz7Jki5TJoYMp+
CxZLv4gzJc3EGDoSL5WWubmBkU2ay+aB610O1W62JeI3hz8PZ9Wf8BCN11FUa/gQ
wsQsTuKjGcRZBu6zVNBrWuZXfRrphNutSLzQ2eoPHvAhPcsPouX538FKStxM3F4K
BHKq9HqM78wnvBqppLKqB6y7TFvynXGL9T+DzKTWPhEE3giMT3D2uezRbeZ53TdF
7iP0PqM9Sh04TQQjTDALjZHbjXd7o+MztqIu9AO6Geo3it6ODsHa5lXQOFvmz76z
k/WlAwmHkHGfT+KNMtE23MBrGymZv2DLQYOh7MfEOPO/JIUPMHpzzq+foatb4LTw
gdbx5fPdBk1YQ2MvEf0ncRoghNpXS9fqo6dix75MM/xFc7SGspPH60Cn3WgI4b8G
DLU7BckfqNe33EmNYIZK8RiC2neVwji9Zqx6OwU0svqzbNjMOGRbs4TFQR7lHivF
O+LvKjWlb7kU2baPwEKQ0A==
`protect END_PROTECTED
