`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7uM/Ntzh18nHk6nViIiIa5asU2Qt9ea5gKL8PWKz/6n7Quo5odRp+OMld5Ab2/Mw
O9chLYSg6m9wg9DdcsiAfBQxkkwKiSgP40XC09bBcMZdv41kLW3/K9R2W3rBk7Y/
vaJEjofGxqjXcOxVUulbb4sJKkU+5Q5ps3Q/HKmqq+BbwkhXV/Fh4jHiv7joF+qR
5uCWqGjTOTPS+i4RAsWujSTd2CAQjAOs4WhcTHyQEX4BhrsWmWDD9MmzTzCCiR9/
Hbp+T85OD0NQbMiRz7fZCJjoBQLKkY52YGg5b148P8NEy4Br+6fbUqk7KoHyx97t
qZIDrlOInFFjf17crrmmXYVAdj4thM/a5n7IcUSyHMlLLYAXW2ox6W6BDBt4SCR1
9Abw48C2+szqDlQXGn1ZG6mK8DdtS3/7NiJ2XliEvHW6eqpOq57wk39bP1NCLIPZ
5+N3hFYtBlyCyV0giZy9Vf0pSN23crYCdaQamnDhC+8KWlyq6c5xDhKZxaY6kjer
06QFQiKCD+nDo4tJQq9gOxi6tpnZH/U5WAHRK1f48Pz4FxWPv1SwWhafiiVa45e+
iDBgtbvDEZ08ZmT7m8VZTqfgDYGIrSksUAx21160fkXDQTHInx/x8S88i92oxH4E
EREoxkT0DQa4SlutuqbrINRDBU6gH0FOJSxWIZ3qz6TBQBkIwwpvCDQjwqGLT+oQ
ArifpPIn9+Xn4VhoXdKsr1lfmjsOziy2c7cUcduR1oE=
`protect END_PROTECTED
