`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z4ekGzL6y658gCdV4Q+fYYOKmmJvHNik12c5QxbLhX2qKOsmuwulFuNwV2kEj30U
BK9UkA6/T3tniTBKDQa4blQxgwqzksJ2ucI6e7Ifz/nEjeiLn7cGDhDXN2StsE3i
9QlkachiacI8GfSx7ZV/z3qYqfNf8y9nMKMruiESjAlaKtzjrrOsW5PVeBGvovhU
/jreMOcM6kQLbCBOgg5y0wRbsc3pYldXs6rpzNW1V64WRiWGj/EaRBxhtbD1FOUe
v75ZQq9P1GZ15WVOErmITjdY96ZZoL7dm462UGh1X59PCUhe/tl7by7TPEq9+IKc
MsPadVybIRBA4+tftlR/mfEEhJApbtRH6nLNOSrSVgWkk1OufhIHcZeMt7OcAwsd
WGscHPYjWveDoZaCQpRUZ1I8qOh4rdLSaA3RHwhk6A2oA6NbUtI5fCH1n0ZNo+Zg
iHKbeJe3aWhE1PisQmyZsAa0xxJhjtU1zs/ykr+jbdhladCMAV2Rhvn2CkLLlpZs
+9DclsVxAdTijCsJJqL5a4JRo7rY7UJrB3rJTgMRQ6LllPalIdgtJUn6umrDhJN8
E/4sFu5PxEtP4gCwDh+1Ve668rbjR+tiS6JZIs/x16MzJyOZWoJt36MVZLes5S4r
0Z8yPeSKQd1G2xNk6R+KKwoMKpSpiQZDT79ws/d1cEdVJWCk55+GnaQ0xvudWb+e
odAHZji2RoG0KqnOj0MBow3Y2tAFdxHnE7yHXQxNcsFIYXtgzL5kCp4WdfOQ+ZUo
ngxrfq3peHzIgKjIYg6047CHiujvs3anIiLFye9VicUB3Ey1iESlgPxWuh2bkVLI
jDiTb4dr2QswD6HaZdsgRIz0LZbrazHvVngjf+jZt8ceobZtSoWyCAqV0Y9Io7vx
nOmp1bs3J85lV19W8pyX6axpMzufeBqqjIOgbURy8xJkNCZanuz+gCAGXekSqHKu
FL2LMoXAFAc7972KcOHs6QlDilTe6NBfn3+xb3l1YtpZioLoHIWjeu9RiAZqcWZf
/zeIBKrCqgvsf3G1PgOCCksz0Az085Afav3KuTXx0c/RbDuTu+vBQSnrJcouNSWd
gglxP2VsvVSoI3Y8BlUOPAPjgcWzA5D7D2ZCaFCDpfoqL2FIL0bIzkTyVMJ+3bem
913eoBd0pbzKuo9Iw4bKHE/BubOJP5Cwhh4banMWwab9PakPmWnsLwSvwwo8Q4/U
5ZODDSqe+qUzNPS76datoc/TY9graJ6Xev6LVQXhAydvWgnylNCGzpwtCSm04krc
R1AHugvE4OU8fEdOcIUpyKA6FSXincYzH9cgeX4EWmyvRdSYTdbj1x7aHgQuGNjO
v/kAdwKHAuCOx9S6LyYhun10eU7XNGTG2bYta2ROZXCHSUk2uiA95JiTlaxIGfJz
VKG0Ggxk+Udq0TrxQl0cO60JoGTEZW/ir/+JDb2JoTICuXTV0J0Gu+Zjfk2yKRjC
OgrAyjqjI9xYikPhQO2+V5rdSrTvrY1VJEeDN7Frsh13uJW7dXOSjCJXd7ZAXdsK
jnIKx3T52UO3J3LzQpydRCOkU/MGkhTIYZ6JigWYHLElEyA2fPgo3FJWe6eM+Z8H
37k63dAxS6qCoXlCexJ+X9CLMnJdRHtDUIw5mMEbSxBk80AUCDrsbM6kzdHYq5fx
w/INM5AqgtpIXxqQjhEhKhH6XS4MngwMWpZo7YG4Ee30BptXxfCej84x5DO1I6Z7
9JPNW2tZ5cllvpFptSi6m4ft2iKOVUc98mXG+jNH7U9E3FMbvRpCGUIblan9qSGj
x4gqbVoW3t+EL2lzCsWcTATjfs7yAw0+8OudsgBUj6pYsKY1PKayVqputQnKvmiW
VTEUgHQgRQmY/2JZx+aAZEAQ2OlOBFgQODkv0JmUGhA8C3z7bd0O1QObaKhfFLxu
GH6olBmhgyBjUrGLaR3pMn85F+kzlH9MzA370zFywU477jCY4Bs9f/iTUkJT5RYS
dTB4MS+gUPPRNM/nHxhA/coW1KIX1mbiuripWjg9wDJJ9SqwXhLL/TBSDk/BS15u
aqZeyTJ7rHLEnTupkxSigeqUayYGY2IS7RxL2PjVm2We8rAecQU95VR2NJX7/Ury
eo3OrVbZme/bz/8tuQhALaZMUbM0KRiip84m2NHWjlye7xZYj/ymeqn/TmcwEsdd
jAIcgUMlbSf2GtjnbL0v8DLXEJRiUZQcLv+9hbN1758PXP0qug5AkYV/PX4jsMEb
9gCftrAKGfsSPEAnn6Za+fCY7Ahxg6RR1tigLTbxwfiJwSQcQwCLo4zPZPC1xAbU
9v65iHQBTH0H2Qp2A5rCYj93RCiFccUF6ydmeVuamP5kSeEdJuOkvFIbiteutYHX
q82sttaM3MmEAT/oXfbBCTPbwh3wO44eNKiPH9lP5vM9ukKLJ6Mb8hKi4CR7fOyd
nCFWORsOjYl2OooOMsnZndu6hY0nAfz3uaTvguP3x4nOolXkKQGbHbLIzG8RgSaU
8Tr6fgW1b/ThsYwywpE0yx7/Bcpb5YTEzvIrSBAoOEF7ivr4TrV3GWgDZGxl6c3q
dkAT9jAXFRxgVdBVyEvxp6dqNcBxewHNF5r5iFlzBkwCplJhoEo46oBiK5jD/DJf
1u/Za3zMQ/Ysd3dT67XhVj8xouYGTYZiZuow0Ugn44BcGILbnEOhGutq3/O1/xEp
3q9mGHJpdlA3JGkwNr+PBdWo8ezvBWGRXyETB0NpyxdtGtOE6hOwLAraIayF4I4b
6MQks/VH5Xfg11qdu1jT+Fiu94CpMWZGYohoNmc757jVG+AILTsWrS/1DnWWJ/kq
qeUEUxfE06uDkXYxwUtzNmuQPl6ddYatMhsBn8jC/rokPX3hp6848OuY3L/e1sDg
nKORuNWAgm1RBLmMyvjyB3vAu1TVN+JNFLUo2bGbF3HUmocJKRjL6h3UlvkGNqLn
x0AYitpR0/E8bkeG13XHQeXbU/R2rS9ypcN+CpwBShAeC4riTo12cqVoKVtiRvQM
DPh/Nxpw8pgTGelGrkCL7ZXLumr0SNJ+oCWcZLbPhlgkxakwG6is05Cmb4BQjrZ0
qrp7wA6jtBQIMQifPqYnE8lIIKTMQ3MfUAfgH0YfIRQgC82r/1nSce5gUO5HDZyA
2vtlSAfPGpP+xz3kayvxsRuAYCM9/awIZI83Fms8IhvpzI3RzWdxqKUTw7Mxq3qE
CeBu0Pht6XArTMaYKceU1Ts40/3gl79Rkxs02J4tbpyZ3hjB2yrEt4ycn1gvhR5T
a4yqyE3DTjkM/qwNT+cZMfwZpxSW+7CYSVrAqCIhNfFvfcxkKI7cikW3TMSd5DfY
JXw7nmxh9EfSPvknATsGU15VLE/kADefSdFoig/C1DIoIisf4ORDLm518OLf1jLr
xukG2MzT+Hk0N1oZvv3tgrFEf9dCRb0qGzU5XnV3BNY=
`protect END_PROTECTED
