`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GKKpKvquIFZksmh064SRcpHD2ixVt6ip099jltM6LetdcION6Sc2OZWzTO68BwzW
gLfDZlyN4PL/flmPYziAKy1dmnjDkrdaTnyxr/ERrdE8hyEOFt+1ptSB0/xT4n/i
Np2SVJayxKqs1emaPkRusPb9ZAaCuhr4l1Q3Kbr6DOzynu1PT0lCwXmvR49QSgJO
PJufzo4jeEszuKoEDtHbCyy5cO3bHoScYhgDb5I2JSLe36IQ9X+XpU6o99gEGigU
TPoJi9U1hSgCHX8XoOAX7hB2YQw2P+qJRsscHcTh6jUTPWHvTUJWJHvU3x+Z4Ox/
OWV0/7YDhnzcOpmB8nbz6cXukU+/FoOjX4ats2pVjF/WkidJezgwhBoy3S3Ch8e4
X2cTMP1MY/d+dfhnqVoXJglcygKwpPd0cMtJ1MNtncylbeUSEBU3aYQCnsksqtba
YOsMozvuGOGDNuW3y8ftUIGNEZhQL1les4Uw0DqwOwLbEwsUr9eQrgD9+zeZNIOG
`protect END_PROTECTED
