`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XeFLwrSPtH7/DSZrduOGpSqlGvhH3x9wrOrHcw0700VhJuADTpMlQZy7FxJt/1Vh
Di4wzr3RlXFKEEu1irxxkEQkUU7mIpnAEIZ4EEpcYJd9ZQr44syuq6oU6lVbEkLN
5JR6VrV5kU2HZsIwQeGHs0YAkLZBGeQ24GsneU9iMMLjrGs9O+MJNUPgtjNZI+bl
GFvScYHV3HsXC9EGfqX1bY51wDALGvlaEigLkR9EK3Sb4W2yoLTpnnEiWpvkoenl
U+eTvFKwlwy1mbceSzO8RlbeQpF4ytDhaqyn8oix3FE5Q0WwqiAbHyY/8mFqSqqm
YKL4x3FOhKSr6Ny4QJ7p9Sbe3axHGur3ryQv2vFyBOYcexZaTifHiCnmHglXS9Y2
LHqv/578a9wAtUY/ixDcIwb4UZ2L9nig5qym1b6913y68XavMLiYthEaFS+XoQL0
+Uw69thl4quPNE6kapuCIwJ2gUgIs+lIjh4A2BJcf4GtTGKDoQxl5EQ5FTmAl06O
tSEl0voEcrBOf/Vq36dBnMx1vUR8m/nOjksQF4lNgnrdcB8BW46TzOPzqc2X0rpk
Br+zHgSXND9Fat/BymcAxObqrq20YYPfwKOZq/UjwBitKsEwncxegg5ZE78Mx2cl
zdAuvPUZrEdL1UkS+VazNIFtFy/AdCqQ7iufo+0qo6WwuIsYzxYNUWIkgPVEW42A
taBAPbEguZaYI9iAgmFHhpLIYT1BqxAGELA+aPdo8EqruXfTJmTtMza01X042rBk
HLMdECP+UU53HnhW8eEddN421u976Rob9eTUV/DIPMr0MFHcGz3kkWLM/4hZURPv
cZX24CVW7X17Wgp20WOxxxLY8850WlvRIO6pGPuoT5wjgSir8FKMZaYraq05qYqr
xgkis2Ji4ag4qDyY39cA2lglxsYswNJbnIVTE+Hm4LR9qnimBwbJOVMPOaIILzU9
l3H5uActhMGefcdxMhDd9qYRPcB/OAI84m+FADXAl3a+7AeAP7nyLL/i4jVeAMyN
+hUnJys5W0w8SGW2F4GiEEgnaDFQv4k0E/UkwvitQ3kSN0e7H6by+V5G5qezc34o
ocrMVLSvCmM8ocoYD3YLIKfzndTleTMIE3SRExSFKBinHQ99rKqtxWRzKQRIlTQR
Ub2ARQCEc4VtTSrzbHZFYmym41obxIWhb0cCYOsWXIVCAun3b3LC5rXF69BVbX/W
ORXsRfnz2dViHIGpsUCSUXhAUN9NWXcpcu/3B1PSUXBo8RUn1OxGOJ83tv0NaAU1
KlbOKQYmUcYvCtD1wo6/IOX/O2ZZ3xxOREz32B14Eqk=
`protect END_PROTECTED
