`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fz6MBJ4gGViMWybrU3Un0BSZexZ2MyNsyTBrGu2Pb+jNbIYSYGd/azakVSsZVYdH
ngdCEjdVizph8yLcjewFtjRCM+Y00stczxX87Rzl1oOqQI5Da2yA8zcRe+tKVXUr
X2pRf3mAKZGde4jgmaVSrn0YLmWRv/dBrpQXTEJSWxXr8KpdUgoeU++bN1tO/k+S
lKUourKkg4yfC1bknlUPNcFbG48xPXrsrHHTaSvOODSEwMTNUq0gcaLPmCbfEmGi
iZyfPcS3G8vmXC8hcEiVutp3aVL8Knb0KyKb0j22f/0GnhpR4IiW0URqSuT7rr0I
dQK4JcW9T0J82kpCW9mzhS6PS6CDCHEUN/sLfihf5j2KxmKREAO7RG8ubRTTvnWY
PMiadKKyKYnFV2xpY8NYzw==
`protect END_PROTECTED
