`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cgu1N1lr41d1jlEVHTh6jcBt0Q+uhxGDCH3mejeO9PdXs2OalDHsqxlYSqdBerD7
gkxQESQXrMfW2/m2hDPuOyP2VFFa0ejHpGHexmsTM9qYsWdD/tMDjEOTH/S4bC3z
/JftXP3XSzWrA0XUhB6MsKkXfRdLcskRqqQkaRuSa5IGNCoTdOoqj5cXyZWl6saV
zGtZkSq13EGJAJR4rubxdsSSSX5qCa/uNFO+QXG3SKj/2Vyg97lSX+esUcNVAyN4
Ov/WUlrSrgNOyqil0gH82y4u9UoM9DeTWpf7HH2XlkF/VU0qjNDAYCPmHn3XUP1V
3/lCXUheRkQ4a94cyJXPixIIK+6T9BdgAlknnjjVxIK7TMfD9Z0NcD9ZEk338Uff
ahzlScKMx3+ByTje2LJsQuW4u7nJ5VT443fKReL1uFAcVcIP5bL4FiXEDV4C7j0t
le3XSwcaUpEQegK0QcmiPAM35effSeK7Xrh6TKAMX5AxOxDiypA8ITBNMF34acw6
vjQNiAOOSaeMS+8dZE0kXblb22c1mK2s00AP4c+0tC72fMcGR5LF0RUodQoqP/sJ
y3uj39dLepGE+5+W7hVOqrRt4nUTQlgFzoqsIKLWvJRw86GcIetUQ2+9CMGZZUpE
ZmWS2gOCM2HQoTkLZHAfPVKycLJhT+CoIIUsVk+Zxq0ZtyV+7WgGmmiK6LCdM9jl
QG0nBtAnCL88oK7WN4vdmPNPcFVUUWSzQ5ODrJjQtBY=
`protect END_PROTECTED
