`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kkupbgp/CzKJMKSM8D8vCR1O+TbdMOwxAwt/XazloxvpuplJnzys2GOhtKlRXHDd
mhrXYie9CpyGxHQ275SiOJEv+fU36z+d6ZYBR3CWcuF0Omd3+HlTgMSsAU7qXWcH
RgZ60B47fCHMacgAj4bB2fp8iHnY+TINNEC6zNMdLw/vIaEpDyyMlZEfMfaZ01Vz
0FBRRZlhflaQ2pVKcxD0kZ/lQrORxrDA9C3dKO9SXp2ogSmv8+1yGD89EfkcQQG1
pqUrE8sBosOLRJD7D7N0XhNYnTaWDG38YdB1Uj82uHB9WY97wml8MBmCScT8s+MT
RL8bnqoaXYh/W5d1Non2Vx2aDkzxJQ40pcdoyzLyX6MXtS/jNwRqg2tbOKYE9hYi
3LORYFCEltWIij+wvCx7vQW97ZhbPinNi2XRkjeXAnPZp1nlCbY+UOU3jK2pEQbS
veFEiRPhdIZyoTFeKVWjJ7zD98HiFJB1P3P7OS2qBr9llUAGukfXGR4GsaWak0kK
dY97Mp+WH1lzftSofSLOUOiL6LkBHDJqJEZEJufobYxbfLFTP4AZqTFb1BtDJmTC
bE8290Xt1j09Cq4713Y5H/VqYXfa9rzhefvcEqrzD7U=
`protect END_PROTECTED
