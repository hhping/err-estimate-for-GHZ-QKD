`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PXfeISgeA+nNpcxS8Bdj1VRoigy5JbwMARqJ0ZpzkJVhRbUMI7Pew1bnjJZD9slH
hupac9hJ02QhpVeCPQlVD31gt3aLXefINV2xTXjG6IMdRUZ6gMPeBCMgQq/C8EWr
wKE0cCu8wapQhAP//kgSm5dsd7tikP8bd4moMMQwWZHytrj/YY4reUdR+U5420jG
fsA36JAiFbKQNqRn4Uw0JvG33XYaS/VzdxJZv/PQ5RAWcBHChAGlBT+GEBlmnYx4
p1+bRfgYRe2SZiz3fbG8CvXVQ1B4O4VPKCnTBK/OI45ut2w1SH3wNpJPTYYcBZtc
8CYoXu/3oTwysQ0MPlurzjnASPvxafX0BNGF+/EMkQyFd/zkJjaDIlvUcS47aHn7
+xDos7GSLMHO6Nd3qazJOtiULoUpiPMUHg3axsnp15N+LQvtMOTUxz+9wqd71MXa
`protect END_PROTECTED
