`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
luYpizxzV2uk1qJzDpzJBx5WhFQXuDShOoJ/JpwkDr+10VK2t70EOgYIYUBkBVKb
YlLS0vPXQ5uU2BQXF0iGhyhubRaQq3xekNQ0681rfBXeE2gQhQ19YRs/OTHxsAQg
RwS4blmjs6H6s6QHQNJDdGaGFTfTFflskjUXDqcjmpeq2a24UTf0aTQNp92OknWW
q7KFvGZgRZBtESyhhcVpcYArhTdQiR2G5rUX2RuWfGDuVSEjliq2a2pDtD/Vj955
Lmtcf7gkUAX1YWYKfyy8fuf9MwdJhk2dxjAPL85wAnR/z59XgmlTdhjSKYj42Ktc
dfDQ7dx5fK3/8HYG+x0KrRz36WgBm+L2AsjqInKVgHs74qPlpmkp7twe1Fy0Xa0s
exgbVZsUxQ+jk78i17+ElxttqJ48UFjDgJ+vOoGZrw8GxvMhz//BmPfg2rfL6DM9
ak0NIyzSkm8JWHIBUkCQBMwF8OhpeVsqVv/Bp4krLRwlHVkoDaWHWEGbVA70XL3A
tVaMzLNCiqtZSNAKh1Q8nYEv5oWDny6RDyjB8MHj/zvv75q2tMCKZj3P3D4M4VOw
f6HWu2HagTempnG6jEt1MNicwR3+bfrAyxE5FFdXF3aQS4OJTKoO4bU3pmedPI+7
W7c+GpVn+HcYgu1WAjWNwlPtPfJqXHbCYLWP1ABLHWfBt+E/sbQNpp2tBQP+6VIw
RUn06qSBGeRBIsB/cUex4dBOvlRDC8AAocrwYQjqNIsC1UEZ8KUtXZR6P/KjY7cR
9s07dQ4ghN9Iwr99Et5CjQ==
`protect END_PROTECTED
