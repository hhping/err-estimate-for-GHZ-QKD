`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SC+nYmjji30ckSEvo0RhO7uGbuQjQgETpWgV+Rst/KTdtTklYHo6+ViVWxyDerq8
M6mZQYNYzB7+bxb/K5stOad2OGJpEbVyNKOoiLnEQs2MrmFNd2pSCuO699Z2GgAH
O0AqwlkJIZroyJYkacwPhCzU04Nw21inQHx9GETaQ1pJSehKZJj2U8rZM1zq5pLv
q/CkWAhZuoJ3wOqOJ6s81w5qeIb8fibDZMPFW59mN06nfgJAFRLlhmHlDIoXK4+p
O5egi6kgAYX7Pg+0c0+MKAv4L5G27eUoZT6MQY9rKybOniXuAZ5oWQNl6EDh/51W
OM+eMoE84etmcCQ9w4gg5YvbMhghPltDpLPweg63aayvSBLBrYbhCHXv6jDOQAsP
vIrMze0yPahsxTBCgP6G2wNmvqB3Tuw4e1LY+BR1cVtdLjoQYV7K6piKz//B1AgY
1zsasDZmubN7tvn2z5G0thZWJcsbFxm7QD4xSz0xjOtt2L8mNTqi2JaTaz13tjQp
WI+bPj2F8A19tprH3REqwCBwA9x5zFs5ghvrnR3MYOOgLgU6CpCvoIVfdYu2/5zt
iPHvssOxs2K1Ckh7akv2Vns+Cri5y0WziaA85kU5gNNAw9XUtrxtmT94dLGjRG9i
tzKOJeTHaFaEYQ45N3XAr3Hh2OYghimAC0mkcbnibxHTjsD1OxIv0c9SmE1AaXMc
hfYqG9hzx4mkus0DGld6O7Le/iSv6GH6XefXH+OZY3dbcHUyQruovZNW3XUsU5DF
AzlTFM13+a3X+Y1y2m92Q6JouXoEHFK6dKYiSMmNI4Woh++0p/bQDYFsOvgQja8Q
BbGbDoiA+SlAoymWk7Q7o82lzHoIvPBaVjb8mayLh//nsbsIRAFm9UKpXI0FoBL5
LqofJUM3Lvot+zN+Rlo4qTXtTTvKDvLsuSIvXva7ByYGrvFraEb5nXNqxNTO2WZ2
+QvoBA6Rpejro964jB9CAYqYkSQaZbKJyW6Nyag+hq6r03eXReV1vhpiqnad8HpM
sDddVFjShWhZaxeWcyf6vEL16WHaLk7HMqw+OooAhies+wT3Numyk6XdYa2lFP3v
riT5M+9cidMWRss8M1yjK//pRnhnOfZ/K8el7CExruOfSZgwVq1eNMq828sk99zN
gDrR3crykfNavnAlSbpy06N43rV8mUMupxe19/l/kLeMeQdoSo7MAsRzH0rYDNnY
bMSwouZB0bVlNfXRxOI/i3CZ1GT2WSKibrbbJb1LJnXGItwgXw6ZCE2oBwCitjE2
5rCje+KiC4rl35jk8C78Ct2dmS8X5V23nnsa1KFKy1+5DYpvd7pHCAnSkCbh63QL
jIJTGdXkpNCWebexYQ4mkCjGY/o7SXu2DgA1nYEKsajRiESqx3mPAT8iZE5Jk5Ub
B8F5ud+sDC+Rw5et9GDfKkr6GLNtFr3NC190y/BjPNv5ZTlz4XoiocAHYL3akbN8
rf2dsLI7+WY5BVC9tKdwuwCDkVp+XQCPaNa1VVwS6Lj00xXFmk4JW3gdO/+TBoO3
ZDLdr1UQrBrSoIIy3xGqz0Q0ZFQ+et6nYdVgYSA/xYLSSQAR+jzwgA0HmDuRxJJS
UjesY5YcDbmKb7YYhNNVa8l1TVTDiTmTUnjeojYiZQIMOF+Y0JGKWzOakFoaxgOq
DrTFOFw8HpH3J91zM0/v8YNzVn1J5qdv//s/ZD/3iBQv7Fn6MGN4txDGZx6yN/dh
8TQsAsC5jHVc5ncPIgViv3JDLu8C+s1M2jwfvJQVR9+1gwLd0SQmsCDczrpE60U4
2aBJ/ebFdBXezijptLz+vrRatA6hINepEjSCBgoaWut48+6BJK+mM5U1jstKkFk+
d5+YiLXIZBRouVc6rFKkPr9D5ksEpuOdK17B9wIUDqHmyYJCNF1ga+JpvJMtkNP+
FJZmMszG9iwPWgPRHjsD6WDBEq54SRWpGXWI4b8Ibkjo5Ln7nu/MoXM3+RpKkHVn
vHlly6UV8WYZwFUxenskWee7Oyl3UV96ieVhLqopHY96kp+ljWHXCDpLh5P+Sp8d
U3H0+yNWWGPBeFnx07Q9O/diqoUUiajvlieFpmIptVLEv3MRbpN85moP43w1lCBP
zngow+3/Jkwy59v1WEAIXD/PZX//PFRdI5nODODa2lfsKYwD9H8bVn86ZlMf+SEF
xGaJV15WGZwkFzDy5068uR9cDmo0THfXThQ1XA5ROnFPnbeReYtkGIKNef3r3Wbj
bZEhbr3DkpQA89a/yT0wBMicUymYK9FcdVw6ZKfLR1M0Y1/uDhK7RkE+35h/2tTt
0KPGGb33QPoHQvaQ5U36Sn20R46+/V9l883tEerUDxdJh/W6KPX1pTTtV2qRsg7J
TG6J/BlS1moKdOr8v0TRC42oRoE3mvNT4XOJnm2epkJN1qS6DklyH1zCoL7geQzK
mtaSAUgfOsbGcxOIMwjKw80SFrosxVlGDyuuQv8tiKv063s9DmOSOvOqkux1GG5r
W+hhmMv5HgzFOq/saIPyTJD4+OidzXCrK/kMXJOMPL7In+Rs3T4G6SYtuN/7HaYP
CjQ9wRvaeQN4+nrpBuug7Ddem44kF8fd1rvV58EnJEHilDrB2pjW1GlcuYUwm0ZU
qf+qQBegUGkNCbbpVfTNP2R3DN04VkdckALPTPVMp0E03JaR1zejLRizS0hQu5nu
/g8JfB/m6AMWebThOynSZBIucHxZ/ovT/e7eBs3/7F4y7hWjeZPhm6xqV03BiOTs
BbrtEBcrhHrEhg43gxU6XoORt9SJf0S02QxAf5e44xET/7d2z6iu5/1qY+5LumfM
Bz8cyudG6nDrRqkJigICd9gxovslSd0G0MOLlvM8MSKYpFH7tdCEcRWPzYfb7Z3x
N/qRBeJSIX8/7c53UGyWiLsXW4k8h7JpuW6qbIwePYk++tF0hU1NSM9wYtr3cL9I
qsfnZXRkqkCHaLaiWnNhbczm4wEKG2rlzxVk3gBuoj0lVh6DDbdMqHunb1Og6uKu
MzeW+5rF53hOsSykdcYatyPoY2eiI+/n2upWNFfPizKvPVAn3YZdCsdhubQzWwvE
zikcXV259n5upXnAcM2ZdDtzLJhYJVRk6cfqspg8d0F7w11g+ODPTDtpMrGAE916
73fFF0IeKZ5Ze6fzMLkU0BEFCdoo34QqVxFpSHc1cCAySDWtmxn+2CrlM6xx13bY
aOSvukmFsHqOXYB9jfxKxnWmI+jE+vfRl4H6QQJaOTb0QT0YisDS8qHguOp6SRex
hjdrfVv0hhuLjm0lLj/lTXJvKAcBvW/qq6GKRz5OHDz11TlhaEahdoAiUCxSfpOc
baPH/92+YIF4MDx5J+SWhm9eMlrcUojIfkqdt9STLM/ekMmdNA+LUvLw65JgbhES
0ejp42iJgSZ/paz31YSUhLfvUTl+kAzYKn89RtqZPQQeFrmnZzsXXFJTZAW7Pxd/
Oe0hOnovJQqOHvjHPK7PAOtLYNhjXQdM2Cy5bevV83Z7lgRGIAzWxxR6RT1h5CMF
Q86wVJRJuLS7kC2V/+oCbxx8dOOBd07XofbwaPEjhpKQOgmyiK3fltC4eRMq+7vu
QOmLNu9Mt3CcV6xeTweq24xqLIYC1YdPMwdbS6my0r/d9CV5C5TlFyWiYTSSco+Y
Vc1tBdvz2EQ7N75zAnEBLHolsSr6SoCR3OqGgR1Yw1rA63FUuWnwFPElB1upEGUK
murkkhhjCWfslvtu7BS4xeSY1YKH2x0HrNaGg3nM3JyW3fCCJJwb1ggXlWrzJojm
5cYKsq3/Hl500UwGVgpSrZseri/b957yR7BjNv6sHxAw7oXTItT5o2gYxBimovXf
HTaQZKmejh2ne6iPk8lu6B+QHhyH4jIi2Kw2d0gh52DmCRKB4rk8/4F/9Gykb3hT
SFbnDZyAyO/wyAX97EwYSCJr8l2hnj0v10ovz00Gz5BPXot33NQU/Ip6/asKtCi8
m/tvHFGRioGFPucg55bYI/8aLd3SIoOnZCXVDAU1IWbCFLT/WMTSgxsQGhwNDSwX
WImj8l41U/L89nH9Q6EDByPaggBhcc++2roQ56it/E3PC+DZ/Dms1sjpcYQU6K+0
1F09GJIR7Fn6FBAFvyMumfTMbqoB1SAKEo1K9Y+fC1aEiuUUlLtZJk8n4dSffZM5
03+ncBrziE+7YmAjagPecauudYqLvgvQwKgP6OkhvPw8hns+VQ1ajVBIiPJFjLqQ
5e4nvAuuD2eQhiTCNH+cEd1LvlrZEF2PSIAqxd6iGaJ5w8jisnvXELuy76HHv6Ag
ZiyKLgfdTaLgpGa5eCm6lxF6Ni9pERZmazBNjAbs2Dehe4t+8irhhKukwZx6+h4L
orzy6X7ST4Bb/Hz7vPx7VZ6iLdGh8dI81VOadShF10SQZ9zuPWAPjfN1nyj9P58T
GUy1YZtZFtm9IVa03jrf0mreJnCLKyvg3jAfydySnC5jB397A1fcDdZ+Xgqf2kju
RkzxVwP68hFPGqvp7GgWG3qrM7dIGIZfowJtxxWTUR/wtlMuDE7HxfjcEthRm2VU
+UXQR7KH4EtIR4fNMXRP37AkR+8+lvKrnSP+qVlrluLvYOYmlojR0BnvN+NekNsQ
Rq3pgRX56qjmgOn3M9AHJN13yBNs+2xEe0CGKi08f4Ijv4jUEqvRcEjjzJ0Rs2W0
SVXHEjF7fziQNWI1e+WtDQftsUO1m2EONJrclqueuZc52mf9JVoRt5Wf4XmWUlsi
Db/sLR9dx5iOm4s0G4FrzSc+YOq2av6RO9BkpEz8lbfOHCcyK128BP/UF0AoDpyH
4sd0DikqB6IGa/ZN6qmfgkeOiuQSkzdpa40hCYTNaJntqwDGy2ZpmQ0uuojGrP73
BlBSDcYc68NOr3KmTA/iJOXFKqWJ2BezfRG/yOtK3XhJ1Q003wtCW72CdYhooW7C
nOtpJ9AeCFpuTSDMCKTJQp6mHP/V9+rNxDylngTfL3ySVmvT25vCYuwnagzjtkr+
kBn3eELCYEbQpCYelglxk+Bf3BpZX2nJRunUfqoaicqb37FV1nlrtpME/rzypYSc
eja59KUUPOV8mZhsENrEk1tPCPw9uNdv5RSZ1g8P42RAwxQ08xqO6S6Xh6Dhz2Wt
taCYIks3/05hiIF/CIYvkBwoQKx4eOL73N24K/ST5aOlg49yF6WfFDo4a6O6e3fc
JAiXBzIrfalY2qqMP+96Rngfzh/tFSIV7OeuON06qBj2KH09QoxdtM5mF7kyxiOu
t0UflcPlSISnHaTdeiia6bD/HsHVdgYWeeW2PYJsJiFYHcKJGheXEyb1epYP8xfz
egfDRI8I7vaRZXWstm94Yh2rL+cdM7gOVaGRgevXTSXuOzOCanU0YYLqFQ67xS2K
QsqIJD9JBUIjYzV25trb8/zgX6dSRrn/nPex5sMUiQEi0+pr7p4iE6tH9Tk+i6LW
uWqnVJYTvnTEEoGOermL/LXPBizoMpBDAFF4kYZLQUZFe94VgRwjhbpk43ter0XJ
IHY5bB4x58xwChaEnDK2vQW1C3Rh66Tt5mfNhwYMmu9F5M0nZkKgQGb6jU6lUuyq
o82vUd4FTVhaSzF7hTtKEBwvWnQE/RvZLsl8fQa+/CH+8C8a4+WRyzpS6W9JS0FY
pr1vDR6LF3m4sUqemMJS5KuS8X1LH6fupf25UbZNlvn/j4WhCNJofabNkNnbFlvd
mbKgn6mJVa9QKad2GKvwWR7PHNZP5/fEfTLkWmsjcQs1USgq+7WaYwAuI7tJ7t83
oCrxavZF+iF97Bsb3pbdS5GUbMNgu/8P6IoxYKeWstRx++/zeCqmYklDuZ7hbUNu
SnlKCf4HAsxh0CjpdDpWHfywW6Fl4IsA10Aja2d6wMRrmlXE8l1DSlCp7qiLDrFz
h73+3jytpvuhLgj35bxdfXSxslwzkHFQPyURBZAbW16u80WaQXF2zT3UxH0Mo0cH
ZQOfFOaqZBRbFPIrCdyLa/7rxgi3DCRRR5qZDpqaMVozl9CcIT84iY/ioHXWUvCR
SWX1rmxisixkyISXG02vMUmD8x9IWksMq0W+asHXptmBXRvskPBM3g5HsO3vVG1S
jH8l9V0B+jGfElOkiVgvQifLrv8athh7e7RyQOAjGNwso+O6SUlcj7btauNUeNey
lV6yyhB88UL2nDWE/3a+r2zIBW6NTUGnCF+dnQnMAkvWdfNTYWN40taTbp9j5iYy
rRodtsbnDRg344uBRI6iyLH7n3FFlR1Nc+CbvHwxHZLhPkPhGYUpTx51izrQ+usB
CW27tHCLX+P9PeU/xGz9Nyp60dJOvAH8gr8Y0CT3E28IfDS/QCA+H4htqz1Fi69i
y2uJg1eedFHYa+YsAyvjI5NGvlXRXLwQgYhFO7jYknk3/gf5mwNlAzPlms1YzX8/
qHK0bjIN3H6HM2i1cfKrLluw0YfJ2uuoa6bP7YJBwtgH5cNAlSMGNe1G1YZfq5hX
vc3i6LK8bnNQGzCqSsC/+52yn0hXwsCP/YysT7Y/NBBggtfCuAtznJTThvkcsNQO
k/Kr/D+26Q3iseLMu2pLGGyViUeMe6OmLB66gHOW1oC0MT7rbKl0/M0VzqtfRick
XrlyPtWaN2+ZWiiYR+Ea0PXZ3/UcRLTbssujSI+a9ctmT4WJl3yGK//+152sPsZO
Vw1zjSfE1RfIjo20BGG7vpuLpFTZP19cfbiWSCxD8i8ucLEVcL0sE3SFaeWnzT7R
sqXQ4fROXRERgTIexjGBMHa0Pnw4Hl6jfojHN6AzRrzQdLGO1LgXGNCvraBjJ6VJ
+j8j7gAfZ6AJ70b/zOASjtlCaDXekxcwg/5brPEJOyMFfjcGq9mIcQ9n+Zcrs+hY
6HliGm2k4Em7oVqOZ83rV/OIyIdqZ+atHGWEfT3dVGUMb3Kq4GtKwqNau7m2Q+zk
nLOHr2XbQlf6lBXvT5NXvu25r3zsx0d+5ECA+gpTo+tac3r6XdCC03AAKSKjlIAq
GtVLocbgfGO4xOzrvjtE+hLIhxX0XTQEfImcMtrGciogmkMB2Fo0DFkKvMJJEjoL
DipVYuObCwEnDMIbY1xyq81w3AENDD73hvEBtBwhTn4=
`protect END_PROTECTED
