`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LsuNKljVHCXO6zcF0Y2TenSLL8ozhDw/Eh8v0VFbx47IukXwTKuy+nNTetLbk5H8
GUefoCbha4hlB8+Ym08835+eMEKinFiyS6Ot0zzcnk/e7C2L4HRtaL4/asOXN0on
H8UxWhMQgFWWvr6fmGorCoSbtF47fHv/oMq9kcJZibj/VKlWFYrxBSuAaaTxMoi2
pah/wqNPuCUxcDDJPKuQp6LUKf4HbshcAxY5s+kK6+ctJ4H7q9m0bFiGuklWEYEA
fmkLQ9cGXBoWrQsyp2R931cvg8eHu6IXCW0cO+sV8xp6u7gwr7oxelg+LLUPCff+
BpdAuridMmj/hMxzpRBvvGYsEUB84BOLt5zAFu+0nxOXq2BuSYQwVDjkHWf3ycQP
8625FZmnElPBFSt4XpB+wgFn0VhKl9ar7d1o8A94DHPkh76fALmuR1T+LfEaZoFb
1gR3fEpZkt2CWwPl8AkAVZU4Ax6ReDLz/u5u1+2QLb7qXV8in0bxTblzJYvEd4zw
lWsLx8dvUYn9tyBceCJ96Yh5fB1ZzZ0Huf+uH7uPMXTrkCYQZDvOmoDPndRRb/sI
x8i0LR15HfV0CVT/CpRIRvC/3G4by2LnSKn1+KvdQ00BTQvWmOxomQEgeIpNkVBl
`protect END_PROTECTED
