`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y20XvWqFiV0/JMaxtLyBGKba4NoEH9Yyj/Bh//M7G/0G7BSmvmikMoepBaGhAWQH
sjTuKBFZ6Pi5Rvl4hd2jKVVoow425lx0pmUhvGIFLgCK/bKdkhdBFLadJ14Ii5Tb
M43jCfS6P6xOfUN/3bMUgCOaVDzOCFKH88d0GSvLgJRiEMpRnIfhC5NSPp6+8zTR
64kUM8ZcEbmxMIbpCraQ11uvPjm7KzfjHVvKmwCLGoUil1bg5y6EqRGtuXKMxNUQ
CNjumuf0HvY/Lg8lG8DJ/HaFRFgL+HQe4VnvZj8WeKJT8UUIPVjYD6YTlHlC+ffX
PowOBwaSE4Pelr8zfxy05nasJ9Eo1+D2oKNkckELEp2DW0rYMvrEsKmMIh2AybtU
2uBHp6OqkbYLFNRPMmfJdRwqZSkjtf6R/aO37THNLfH7oecY4F+iRvRmfMclrPQ9
ZsVrpBtRo2TMbzT+9546UA==
`protect END_PROTECTED
