`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a9k2kDT7DOwvfX0nExRSKCa2raQSTq0LXzrScvHPWsoAXERprtAgSHIc8/ZaXj3d
9mCkzjIrikm0QSTDhkbG9HXRrNM78OCARYzABQ+6R2ohFOaPmXWAFim2h6tE+WVp
ZsCmXpLdDoMkB2yUUaXC1e6ZPiEOFvysSjQ60EUefp+F+jFi+EGOVnPH7qz9lrP/
qxrFbeNSw8ubZ7cjFf+Gqnuedfz81srw9CbwCHr2rHcqwqZbS2MlU7d5AHChSS8f
TeApNQbZAMI5crNzq8gALf5fUNSxXJpH0vqFyPT8aL/O/9BkvDGoRZAthoxpRtQS
oc4tiTK92dXLR9myeT1n6GV1sqFGR4i0b5ymY1bF3ZEBPgHdBmtH9r9/7h/yf2pa
bEy+vVWwU2qjYGe//XLkp0uS1rnTroz9sfWyrtWrxPiAjpM7ViQEMmsiHKO0yX93
vfqF5ZWIdjwBkLfNJ7pAVXWZIhhCVJEQhUBt+9LTONB3qvQa2W0QqSu5SSWNO4Mf
q3dC+sBaSStjae/1kdZkDjU7tz7CkFHT9AYrG6paUkw+/UQ3AL+yhAzO4ilXs4A/
p/TOZrbmbiaBuC3jjx8lqiO+03LiFSOmlkIeRqvVQy77yN0+SUEYmF6VHbQJmMAu
Rgurpm7ALaJxE4zyoIgHDLMhkBfmEB7YBLTznKlDDb28yMyFWmzDclGGj6fHtYfU
sVCMOe5cxhkFmRbLdyFZFPam8k4Xq6mOkkXcgSjmRblX62aQ2vWMqoGOiPnmj0O1
sHPFfdcseP+XuA18ovF0D/2+G93Ezy3BwNvrLoZny3sNnbiQ/D5KEaWqMmbsE/EH
Kt1Ygsxgrl6MIyUOie028pa/HTmMAFs4Y1FnQRKv0c6GBZMC5IxHQ4ogUhV6znbw
VZcb7pkXrH45DXT/0fEGIHd3OiYRleLvpA71mXXFKBCiu7vZzj7ZXsNyHYFAolyC
OQHH9WFFkqkj3EhamhgJixz6yzGScvvUopH/1B1kSM8n1A1zPOPZDDFcd8Fn7gCe
/b4UKCeWNpQQORgsomBvZSP3gvHtrsoUJtNK7jugpCtkO41mwhebuS8s7G2IGWFj
OebYYVbI92cYKbFZrAbIX9tPLRESToRP9aKqzWVF/lKBXInCoytvSDYy23EMkgLn
0Y1QJVqtUbhW2GX734cHKvdm7UpMAcdI4P/t/vy4zB8Bvzhc29pWSKk8Hi6M/vEo
BUWl/wjuBTT59TO9sVDrOwWs3uRFr5gLOA1cLgWoBs6aJTFHD+5cBDY3XsHzNqqE
81xRLh+qzfSGJUfAAKGO+9DZGv2sa+5rHut2JmYJzZVwH6ZSbXgfjop6aT+NQ5BQ
ZyWV7O9Ck3kqrIrnLIzjlOs3jNZZZimNWExa7XYM72+Fh0fNwYbb277g0B/6eOxl
RsoubAQZH8g8N0lC49j1uXIH2NEclEEHh8k+mwEW4+3l98Y/bf2nubz7DVLVwX7D
8x47y8n7pJVexl2tgLqgJG33r4vzXbIHE4YyV+Qvpq0O4iGPW1jQCq5dlqDQyEAQ
H5ODrkp5fnNddIUdluU8c6DOoodlVQxNTRAGekPkyeX9O7zieQaIYTkoC/juxh4v
tlRkio/yjMuh1qrPYTVsvxmBltxZf2hD5OQwrjUb1tvSch0n2hXRFkyYWBYu6mB5
eNaMSFpRUUPDXcnIw8EQMA==
`protect END_PROTECTED
