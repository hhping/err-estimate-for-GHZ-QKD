`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
buJ2yEZQ6Y47sRt+JdSKGTqwTcioxViSYGbwGry4hyzAzWOWdjobUqsYnfluwjUE
G1XqmEY433YcvR69luKbYAPN2VMWJpEL7JJK2B118GUuOIuyeS/tNd3Nd8mXAm9p
f6eebNGjmjdM/e/qIOSHxTYCi8q4xNm6kRlr0t/47ofyFpt70hJkDLdyw5VmQius
61wK52flltO/dR7RTLLcsooEUMo236ACaS2sjLVsu31N6Kdkg4QhefGoSieXWwIg
cH3K3Vygl9qL0KhdhrsCFAv/FlsTVNKH+rKUg9Dkr+i/lomeda1eW+jYh+j4uvgw
TALFGV7DVNwxjOMTHm/tALM7yGwA4bwvbK/OV6m1o0e3+cfWhcLTMCbdCkAQfhJz
BENMkO1gFWCe7noqZQgyt00Ujzod2xGk1voxDaRTQacddU5/tKLVv9ZTJxByOMZ/
M2R2gyplo01dOs8sjO01LItQaUn2NTN5sALRW5suLfZVAlLgmVnrl882wKCOWtPE
Knt1nD6Y6e+G5tZaRH8Eobpwl+4V72/NzPdUmcqktDJo38Vd7YmyZoHQB2EiLvqd
ij6YOQB471RaqQaeGyCFLn5n5VcPIoi8lqCRl3ZqDAw7tf4S7wrzedeEOSJEuokb
QkHbJFwBwqHzUzBmoCKirZbqc5PwNXy0vmr/46no4oakFtyamX97B/D7DIvdW6yt
iAZNXsKSYb9SkFEpJw9JcFcNFV01Kedt2oAJo8G1yJv8Bn9a8bgTrpho14H4VAXd
l0TyvsiXKK8HvVrOExK5SmqUAR8b4uB8IAa/wCgHrgKdYRJQZBQ6sLMVKfSrMhmj
DCWpU10yi8O8g+Lx7akhTH6CbSiq5TbqDU72Lufe36cuaNtACvRpQ6fIb07O4Bpb
YGhnOqVC6779bZnvqGdP2St7Q1lrPzMWLODK00pcrCE73sEnDkmXdw9jUIdexo7k
iuAk9XYwt9gclTiijaPW0PabDMizqC46qBLafBTRlIVjrezAMGNRVc1X124dTE86
E1WvMUjLelGiSqiTBN4QusCr9GKZBrXJEPk1tgE4B2WWk1f94DTUdY3xm2L8sy0Z
93ZQNpQyuRok1+XUizpzd8/WkAB8zvIL5kqhlYLTCH3a8y/9abgiAc2MydfA6+3p
0ipsArWHIumkVBjFhhR80mkeHEL2Cy/sv1N3/xbXCpy3R4oTLc0aSvF1OcNibTgi
Tv4xD7NEfZF13NFLYSqXmKmPMcYNA3aZwwGc3mCLJY908nttMXd5NRufUCnvPs0M
Wt391yBzNytDLFRb4WXxvu0LGh9icvOUYAzUn4ScamxWZrj/deyM/8u0ChRSqmRv
mAQApDXxBt+lSmu3IqCrKfP4SzBNtPZwY89P+/f5iy718ubZ9t0KsGEU52WgzHQU
CHvADlG56PQMJUt9LcIHTvHxp8cQS449SXHZeS3jn+QxGS0zTmOmZRlcyQJ/L1nP
VJi97A6mlsdVziVC2FI6unZiIGGuXHFEvxu1dj4ufZ6LyshDievO5sKTz6hN4PqQ
kWUCKpxd5/lWDCYJWlDHVcdatrJNYxy63xXxI36tzSYmOYttTy3ss1oJvBHAsigW
qvDT4QR5SJSrl2axtTTgk3/82CDC9VXGQEPU4JKLUSTt9brfAN2LUGH/pt3zFY0r
a1Cp1igqm3727886KoIMvpTFb2mv7rCYSrZ2dUJoVc1htwPtwZ2g2nzUFmPXDc5E
wgyZbOedgFdZ2XN7DWUhjqw0sFpsIXDGotsIC3dP8sQHlbXNlySMtYnsFLqhtxVc
kT6AMQhJRo7/i+nBpfD5jaYfLLmZUjxhgLbYrXlYN69ZNv/52+bNYbnWvTGO++63
/UjBChvq/wnvSjY4nz9X+dXx5CBvLqsAJfOkD/WGLkvQSvacwRMcmacsnQh/5zDl
atHAha8hAqrGWLM/bxNIVf97S8JNpQ/8w3wDvdNkTWgw+2DKc+wdQGDcRwAWmAfh
n7ch9kb0qlxdDH8HRdUXLGTOtvryjyCkAQkO3tDBCqyvJ31nA0yBECWY3bIK+MBi
Dlx4Mx2BKrybBVvu2beobWw1j5E7/ByHLkv9irwD8Czv/thFpcByfZrk/E83p1OG
NRZEJXRljmpvlfDP6Q+wTYCzhKeD6lVMlO1FLX4DCyU0MwidJpEqxr6pAU8EDEBO
ifD1hbJniRDczdsA5fm7kDjr6fslmJtnmNjrCCiX8CphTEtKAQXd+M3VZoerhI3x
OUIIkQaDDgS2QO+68neByh++qVd3U4kY6PeEfc0NbCqnI2CFvxO7K228i/WKiU+c
LA8hy/HFRrynyyrVmWWWD3puwlM1FRhJmO4A45TbgDUfS+IH6hN7OngrrLW/3g4E
7DEmqF9yC/feBmwsM/zuezc9NvuwztwmpGeOCY4cMwDEVBnNjY/V3whwXpWMwBGp
SNyLcIvnrSpDnHowsIK3E86UJt3Qm8gX2HqcJ8aYrxE6X3dy4n3jYXlss7P9Ue8/
lloPblKCeAdMvTrdUTYt/08Q9/MY+5win6ue5dSTZEKQh18nFybZqB1H2g/KJLUZ
qip/nSjKrfcf5tTMiCEqcVnS7RgM8UFhpATDxKS0rzBoH8GsHPcFcyZXfPDOnCoA
s2gG/cC6vrFn9Go3MYnKaj2LlhV7+wULeAQ7gzW4w4wXYHAopFX99rnijkoYJn3M
/8ERqmaxJc4S+VkIxGAZBRUy775SvYfJj0nNggSczEDQdKrNj2BworvtJqY4GX/B
t6uXxq1hyruQGHzzWRnfyZm/11N8i8Jbns/8bIAmDeVMER/02EaHWqP8B2/ex3HJ
Yh2yDLkzfX82Oa1vDo++Q/BoQ460DAsRNumaH4JZ54qbM8gCcA7IyMOALm2nLzbr
gUOd9rYShAz5um5mXO2fTVVwIlZdKzfuaVCLmruJz0nPXVMKKuikc0hdF+RUrQak
clAT2Z1EWia9RWCIjlh1YsyygR3ivFL4BsL8Pf9NBQXmiryIyH6eSR1dWRrB5XbT
xpctDNhgzyOW7bX7hatcGZDStEuan89qpn11J8zwNHvNuZuKdNdZqTxZpN9UKHFo
YNSyIGdaLi9GJzXnEXssEvaM1EWGfyXu09U5BqlgGa/dmgt+i/xt9RCpkcnkU0Gg
Wz59OxWiFHvSnhQQblyjDRJQ352Ph67YjgV490Fc1jrpIulj0NHWXv4BWxPPQjDU
nssykkGFk2II5hwJ41D5A5SEyhy1NwZiE+iWhS7i3NIEM9BCSVAcV1oKYG9Zm9Ge
8O/f95lAiW0vodNqnlOR4R9F5XeO9BEfipnJ7ArZgSLx5Ay/UddNzft14FzV5QVI
mR7EuI8NxbWQk6OxKlpizhdOv9TiDPKYZ8teCabONwi2AhMfVAzlC0Bg96otObuC
a4t0QrREy8XtS3p7cJ1YIK2a9SR4FYPfWKOOadts31CRPqur021fzF+IMPkPkVrB
BoTRfyqMFk2t6bQ0brfVHGnI967s8lQ1HQ9iUSBElmqLX8kdrEFeL/xDS2qYqDa8
y/dq2yruRL/BFhCIRTK6osBISr4L2SEjuJDdAARdvp31ixK/F2lprgkqcGkJKm2B
MlkCLvJ9ir+Jd/rQCPnrY+t+0iRLy4RvPlyL0Ip2ieE9mDqF2drdvliG7S1COMEp
Z3tSGZlGvtTHyBj5GKDIdfDiEgEbNEiiirugllIlFejCqHU9VG8RCuQpr6QXcNhx
lNSsYs3K2kCZvWCqZDmwnXTaMHQ69peiZQEOk89hULrdkrZk2D+oJ8nUQuaY0XJY
lliaP98G/YJjgbm2/5BtH8O7TF+iiuLJ//a/W1RzfrxsOTJCF4ei6mGqwZtmJNbm
hTAQn2j9FVRR10miFtF2L/V62K3y42OEPNK2XFwC4xchJ4zEZUI4+ZQFUBu9Lx+k
cVLpjY3HoutGDBOfma7+2BKEfOV+tsbS/V3dZmeR6I5IiBP7Kx9kQYf7voInN/ae
bKWjglwejnhsELuxtGN+3BbCo52eVnw5nZk4wwEPiMfjxPAwRDQwgFE9l/mF4TYw
RuVwbUp+dVmumYGY0OSy+3mMEErG+eg1rx1eN97T5UnowShS78fRo6qZaqm6wEys
r3ZOM1ZhH3lT7/RlYwFfZvXlMf/DCAitj9sLuWwXjmPkAL5RC9QKVXhpRLJG1Yfi
PWTlYrdkU4DTE8ZfLfdj4U+jHSlFlgLZuMgWSADRAgc/b9WDULgTNrR79vbj+T64
Jgj7Z7u1mKvPRrw0azZBjQBTVao93u+/zAC+ZupGavR8tSTGX9SMm2Is2icZBIzl
6GXC3oC1cnBQKiQD5U8UQQ0pb+T0qdnXTZEsKh5Zj2b4/fB80u+DPW9XylPPv+i+
dw10DYCXb0TNqBp53pHgInjxc5GfapEhRFc8siyMfgM9lli5v/wnyazfYlAj4Eai
Lyo5buCDST3e2HfYkQ+ug08Gfvde/7LuMUxVGBD02ihNWIOR0Vgm22nWkZuwOSCx
3KLzKRuw1W7dlegNgNWAXkbbq1sm7huBBWyUeKOr7YAEnV9heq0FGUWNQpqgRy+V
NzEqu80xlo3rNjX90z9tfQfp1h80n7lCctrLsBpTu27yynCJ9G12QQvxJvNaG2sl
zGpA+1RV75I0L1WuDGwVdJkwpylRwwcjddhuwHUM/7eL0VRr8RO0Bx+Nt8n8JP+1
Posrp9qhTRILT0X4yrl02mb3eyXme/94TCHSNpda20fnNOpe88hhP6Z8e9EllMFf
8UON1LLUS4fcwYDQ37QrPONqsDZsupBK8D3zPtXvRXG2WcQV8XlU4c6+2Qr7XoNL
4UALYsB3mldM56ab1NHeXHjdwJnyPrNsU8aYJd1Sb8KEJJexwYFfIQ5Zr311itMh
jpXSq6ulN5LzedwlG5hFrjIYBy6VdN4svFhZjzJG515vAbu9FaGEPLmhJWeASTAB
lNotHMKhrIkPn+0izx9Bgy2pukA1HT2oMijj0FE+rGaunSb0tY8lkKNpTsRpSVCg
A3C2zQlcc/NjlUZto0TgLGx+bqDEjhr0moGMK5qCNv3libZLNnl81lecdlryEH2q
IwGNl8JgLZ4A5QdhYJ0GzDC9J/YCFrcDlG01HTsZr9zVbyzXTH0cxlo7VWRTfaZD
YNM9uDBPUAh+wXVkkXtM/DuPHlxIIhQFfmN3QsE2YyWz0O6MWjCvFNz3HqT7mSNb
gDNn2KpUM+hODv1A2CR+bOkcws9jT0WFWR3QgDI/SLCwXzMLkSp490QjIg2sgsjg
dctPSADbS9rGpKJjsMd5FRyzNBQREl+Vi5dhsV65M9D3z5nx8f//7yVwZtwr4AXg
/RxW7OFT3jTpRaJAa2bH5vVlOneXaubfTowkRla0I4lOF+J/fGhhtSqmx6bD0fg0
FQ9YTtXuL5+bI80/X7ECe5GbECvFnLYi2FBPSWVSbm6wM8BGchpHA7B+YOPt2+Bm
XwOdV8Jb/hMwYH0jn9xlj7UeSTPOBg9GvYuvfEhheiAn/DnjvkxYl3eDyzudVmOx
AE7jTalZKukV6+mrH16iXB9FH2zziMJSnPMuIacvqtZC8xVgO4bfybxO+yi7h9tZ
NkPAkI4mioAFIDTW14xFUK9UQqug2xL6BPLSKis1IabibR67lNs5/Sr2/vm7KPNs
yFJJYl07g1W2BsJfrw4pOSIO6ONA8xJ6UqWosQvPRGCX7ski0FTSEeMTS2vAf4wl
YGepzv7y5hxYxZEkYGfWZ4/QmTq+PXLPa3fNlzGmgqZpBCBLdLaVrP92cJ3MxLCp
qHT3bLntQ2xgMZDzLPyDM0h/MV371vxC/+juHznk5at9xW+6PJYocNKDLoxgeNp5
Xm68PcjV07vbC4uQsN3VExf7WD/t+RPlgEageTwmKr9IOL4a/+zGCCCCnjM9YiHY
oWYV/uvcEYu2+xsdlDO4DoVFXZKDDC46Lf1MdNRqQGvhuu6UubwKJMQudAFVIfVK
HI5nk1C5u9k/9yuj7rWDd5m9XgZFkVkJLWKsk1pbkE+xvR02SNrLen3+gjmDmkkd
Wt4xSgc0WdACUOnvmHraiyx7xej28lrpIStr3Q5rUV1BvtyoNjKUy51w9SG4TRwg
0GYEDBVxfUmcXA9ByQUNwwqiHmCLXSX5O3OpBcerJu2LQ9OFlpLxY0J4c9xjKndv
V+e1wMrUMCDLiSKRawR5YR+g2IN2x/xBJjO8EG+zRkgdumYyeX7oCChuWla6nN2s
jippnELbkqe6B+Cfgapd6aoM6OjV3L73dNXYUmn2+nbBrzabI/81ZHgnQ8RxvM0F
Ku6QK4riCmYtvMommeEGqmjb5TJejIkKhW6MzmRCVwBsZ9B++OO2n/MAMEmIMcjb
2vAS2J1A+mmn/kjyN7bxGRP5y8LNNSMtScN+mkWnROOBr8NEvDktPSM0Bfjl2big
O4k0WVsIv5K0dD1ilQPj+2LwuHU9b55c+jdtXwZqA+Gl6SSvO0pvtfvEmtBVOf98
52Tp4x+8mNLJCYI+4tB1UmmxNFR6a0y7UIPQhvqriyK/ESLkZa8GmAK7rcUnmShX
6GW0wZ9Z6TpAb5BgmZcEOZ8/c7Vvxqr6GBUtIoN8yntIgq4YqNB8SzQ6+rkXvcvs
r+lnCFqfVQEoeviXBAfdstyAxLFyM5KBiNFf/wAi6q3QzpDgY3nvC3IrtcH58SQJ
W0RFHC1QAsFJ5WDC89ZxmMQYMRDSiYlumjPXV6HVzczVZh9nuVF5biS5ydn/apJF
9bPxCuwYuKOf8cEW/zYy9ilqBd8H74s5rg/ZtFkoJmqJvPb+81I5+vawqz2yQvMV
G0rHD3M+TzOU9Xl3sYb+RKmpz95noJIRmOLZwmkTPlY6Xu84R4MfEnQpc4MM4xHf
YDGri09pOnICel2WZ0/EwIt2/Q/XuFEegaAw3XK2kbF58ntOqtTHLrqWouM21gWg
5eBqtSFUFHgX6dTmyoRZ4z4MZivHHR5uobkLwMlrKujd+WWI+QILowPBKIUIrK2O
4Cm9o416gWYZ6XDcBNbMC82q3FdKMfKil4SJ1YNt5vQlEY41y3zpB+2cRAtMfQ2+
M1Qdjcwik5sGCtqx23PuCbOWua+PCgMTEI4HFGXYV7Z4YL312IQ4idrLUXVoDqws
RTNoCpREwJycCGu43pzwVRYMr8SBVHkjc2ii6ufb5KtjdwxfwfqXGVhbGnQ9xOS+
NeUhMYFBfkLTchSLGhqFKP5wbBXcYjXJb+Pf9jeP3HMRRb+3v19MLAztw7jPNkS2
0U9CvqT7S/rTiR6eiUXFemCaMQaZ7sWMJL6X1q9hCKazPWNHIOoxWSy95foyxl60
BHvWoLVaZCD39hhiFnhNyqr9FXnL96Wta2isbphQRvhpTaGgKxYpMrybP0CxnF/E
7h/hfiZh6d0BVqTk1QUAtAonuynJSoU2AGKuU8P3i/h1F8nrZP7+Pgsmtpz7S+S4
8FEgUslkN2COCglfikN7ns8QlPVqU6zSb0zfLnOTn5yLjgbVKdX3kykzBe8luxXL
grqlq/hUyd1whwY8YxoqCQ9zXS4IO92ZNiAKAf3i42gjzt2YX4PaBG8U9SiHU2qC
C+TT5dyvsP+Lucrqi98v+zswJIW2DGqhAaD0SoWMYyyeUqOVm2QyvPZcTdblD55q
0Yj2Yv0nH9W74+bLwpTVoygP+3CjfcDX+IUsSLSlQWiy9m8wpsxxayxEQnIWOdqi
XFZzsKuH9cKxSGmrMLoC97nRI/4hFXggQKgblDmQIbTCtWBFGCqqE5kjd3aCXgqh
/S/am5CALlDlVPl5gLirCE0/06xoKUp2MgtGI8s0GloJ6ok7wc9zvTq5P26cYlYk
+3T9OuOU97tYjlltvI2hUr///uajvqoIcxmnhkEdu+b+hg+Bu3jtN3KbW/wQl3Gj
3mLcyrxNmuqhMIA5jftgSigohIuwPmfaU/jQjTYZ/ATrPeXQCixrXcRlYgMatvKw
biTamjJo8JRh45liN2/ttYU2hgGLYTniwiYprZ8S4+zw2VfRe1jtBNHMKB48E2qy
yv+bQ+20nOPknCqStCf9cQltK+SLpVbT1K0uodpMoEGhyaXVP0Iq5AbqAyrmF/kw
qc3pvHrwTZdJF/8jddTPCelxoBbQvxeWQZHqlmhc//f+Blz4E5iKGQd3Wt83lKw7
1QF/MXeJdiGcuWTHe+LgsOcvw32r4rU8PgtHmS1zASRUygSFCEsQvGCTIL3oKc7u
0wpI2tyg5UT1PhhM7T/9ETwJSOdlHlTyRkCSwIe7TcLT+w3wpdE6ydB/knTyZYTC
mEStqUKkBw2RWIEfbuqSNQny8p+ZYurQHqeQADvF1QS469VfO10C7XyYJVkcSZHl
L4J5I8Ddhs5aFnVw6tROJTH1pfh1yK1I1i9My/J0VwcvAhy0RjeP1+9GYT7A41bf
nibkD4W/81kUPEenzR1TMxQLlXByTLnVpU2yYi0WJya4Nf2h7EFbzOUmTDjnEg2P
2kmFnkcReC3vnOCIpmFZMqmUyy/QELTh4AeR/A0+5U+fJAMDHaqg8cnQ9cInmaLR
ZgMcu1DJn6XH5WhUzAdkJ6K63d3sT9Zk2V5lX+o387zGZzH/KUh1nMXCkltmQNiP
0yXHtrT9Y+dhGNtMY8EYODHsgcc9gVxcQwupUUyEymfyx+hLfaO49wX2Ym5RDyXr
DUEQloV5mzMexR+ZDAMq3o4EBeTd8USpcd/1sN1HALEjzTWrUrYnpEzIvOxCGzMD
uWWJPDJna/DiWtTkJjwkRnF1bE60UlBgJUm76PNCXfDYlNAvIp1gKt++SSuacsE4
wWgvSznhxu6pdse89+PB9sPdQFGWhQJJLsSZjECFei3eP6SPQQfDm61t3lSZzhkd
yVTMq7+0o8knh5b9GlAb78pylXtUSYLQf7o/2h3gqoQvP+0O5/IayJy0lXoS0oRl
2wlq/k86HMU+LakaSCi1XGbT4DmMgZbeMnAmUBDaqBJoMV+6nglA4BRzi5ToSHa4
RQw66bLtVNi3spyF/HAVTL0WEo3HfWKo799v9N2YWE1gWWIpDUTwuv41lqs/olgg
rXntRlv3VZnrZBAtpHCLJBjuCymRvYcUKCt4C+rzNPp9bEPJHxF/RV6B48MznGnT
QQFPQMppfs3yRxTilKX/OCHjlQS+GKCvTYqf3DhdhN+kxu4VVIvmc5a3YFSsYdmn
B2Q6tWQloUlDhz9Pt9ovf5w+XhfLpRKp8LFOTuYk278JeCQzSb8Hhxuiei24Cjbg
zhv6xNcKCmXDKrksxfu6dBXdadVTD/Zfre07r1jm1A5EiuQQ2+0HEVRJa6Ny4mfW
audHcRkhPfmHyy0jrzsYiruagyYzWRDOOBdVP8PKlaULt5C/baXH0Ct0t0C1WglY
aPYZA/eulNvuauCdCRuv7OWqH4DmYNjqMMKbyPe3vEhSUasTAUFA26KJD6JYJ7r6
gSIuEFWJk5wVnfaLQBk+wKI8BatJ638yCYvTKlzXT41gNgp/hruQMx0s9dvCEqcI
KA3zQ7yERm1EWzFBJTX4NLIRXGrLucb6ByErkp19Z9MzxG10kqHZ6cdjEwx9RvzE
sqOdc221BKywMwT6Cm5vDewjcIx03A427wqY46oTnwwbixY4BUXda4n0t4fPG9iU
fN5DqSaPxHO+8iF3SSDicmD0RzTvBXEhGXkY6v7qVq6Izv/3MdmtZOg4bNsAgQTb
MvkaNTKl0jAjku38+fx679JFrNz1IKRTZxv+Qyqc6Mnwqvc6u9Ka+VQHZqbXNLbo
uHrOIJ4l7EmtYchJdJzLYipKOIP2L/kAywG40oKRz8mFLHAl/HBM4Z9py7sais+m
SdnwE/nICYg7UKS2nUkLuUDNQIfSnGPQZITHJ9U8xLaT4fPHDC5FXlaoYP6RSRMY
wupTnQkqmd/bMWWapsSAUjp9lqEnx8DLl/gRZxerYzRfss6s+wQJ8CD+UfHNNC3H
iWVEImcRedxFOm3n4EdE1eK9aFPZ3tRIS2Dcj2W7yL3WMyrh88h3fwIyNjoJGJQ9
LWjIDXaSiMLGieequKiLfOq9sjg1SymeiYQ1r81TlTkiyMrWCFkpA+2kOR8twUHF
OmvxV8KbmJhuy9jU+P1lcJYnqv+Cn8kOkn6QvmPUn2PxHPBZ5+EC3Izq82onCQh5
sOjkARwgBs00b6dOLa/EY5naLk6FhtnkXmDYkHvYfjJTGe1cSTq6NTmz6TgKE2xt
pHr4k96xHgpkUz5hslvh6RX0nPXJp4G+T/U1ThK/L0H2S8pP6BHClYMn1wLl1P5c
x/iQfo2vHx7QNTYCMx66w5pDnYWYh+U+NGBGmHFx1mJYRu2lg1blQ/UPFM4XyJmN
kgNHboXObsfch7oTdEVITTZvsmJWX+a35+EZAyI+pRq2PdcH19BWeOOxjXpJtoNR
/KwBB1ATJpOYjixENzSLeEyzanCKi4eHbQXUXupLYOMDZIpaMQYSMfrE1WyxpcrR
Y1LOQAVC66l0BObFfYzQkHLaNt/pSSKk5vUBEEdJgXfnIDQNDztq+qpeOWDXtKEV
MJnbzyDlbitH0FUGYPEUxzMCqsBYfvSt9B2PZ5C3QwCISqiW3KImUtNFKdJdJgAZ
jbdvpm7CnQG4Ts/qZ7O3CsRP+5xvOPeSifvG+krvl1aFpCGYjx/bUO16tPLo1ECy
8gTgDHooaehPVLlFox2MbrWAy/O07b6oMPWV+aPguNK9ziIpo36mnxzZtb67+YYX
iPfzOcHOYXW/vSOd58csHAMBj7t9zUSvPqaxQn5O7jn5gbb/623SdjxmyLriJVAQ
lynVo3T+CCaHcky7sM3ZjOOsQykjbPQYKbtFREoiLMO6W42XAEuqOAKXG2IrKlku
U1s8aHtUdTzszZTP0zSqcD3AU7V+dVWnC/3TbA6G5yFUgmBLUq05mSQW+9XDS/2p
+jFQ6D5d9eD5z6R5mwyNYXg2a5o3sXlngchXinKV2SXCVShCjgaO7UZNzMhON3Z9
lB8TRdoQwGT28ht5gAaJuyug6kMfpwre9u7xCa3ER+91MYw85mq82cuj8nI7QIyQ
In8Cko0kq4jtJdn1hoM6EtgymvziGuExgd4lwizUrNzl8+tL7DFFCzRz14xXLYTF
EygycsXL0ZHJDpcfg4spI0kHXyWA4Gpm8iNdStcUEaTrNBM/OCJwE36kxxRcWFNQ
bN+uuT5aJaUg0LTtHQxS95MmeWqJQKGJyWNnV96So9zrxwcXilxjbzCDXDeyBgMT
1ZQh+I3EYgHJy7GX+SJBVoEfx3DpF94WH8TZOovRkBJFQWq3gs0K/xP6Ix0XqHKA
vLxNlwBzvirZAurHjd+t4AH7IJg9UTsZj/2TsJCWarJaE/l478UWHQWzDawaZENn
xyMGaPvoxE8V6GzcXKb8IQf18k7cLP3V4MkPCXYU83KY+KvkoEV4v4eg7qnnvHIC
kZRTbQusQNZjafOwHiZwEtEeXTZf1Gn7G9zcOLogckjbR/kqsAEXzeRfAl2uLpqz
A1KNAEKvHLcLNqXhWKOyXXK7oOYEnqtb68K1rcy1uRRIEvuWKFHYL40W5L5rwKWU
TbOmmS9VIFHzslRRlJtpeYddzf99nJ8nrDMECGoqvTA3bLuRz9oxCvk+/8+HVNDw
3b7+5biNd9ehk/+HnYbvGpsrfrqlI2qzUc7dTStb2NPzFUMC/twYkzo+gtszflkQ
xMIYlnpseOH7mA1/F+IGYtlvchJurHg2wRpydviA7cKgBTprJ8RgLmYXDWPQBTdP
PjPOyu2tBIHFEWVUj3riFrnqYEuyEAvWq/wdPcaBepIt06tnwczvSA1OZEUQ97Vf
YRzI6j5wT612qLRj/0XmeKc5hev3PTdiC2dq85WXZxhl6OdQCCK4DQuVzhUPmmWu
PJ+Rauq4vVwWw95dI02NgY840xBRRGr7kkcz5X1LwoNK7JPUu21Ihc2JGaXqc4Tz
l23kZi5+8E5nvBysFBu1+hJ+ZfPiP86hHKM5wm/lbFG0kJ2Fsb2RvwFbbN6XTQL7
UO2vj08k3pwAiPkGp4V3cW+XV4ktk95PxnYoF/z1FGonMwtw2lYPg0TA5JEQK04y
qtcqihvfi9ZAPC7LNML8+CerZfo3/RRxIb77DbcsaOy05XeObL5sC5qi3IKkNGhy
rqd39WxXtCNH+ett7urZvF2JJEVax2HqtR8My1JYlYypfYW33ooP1bnKt5lT1h2+
J2mRN/0jun3P32P0OrjWSHWTUhqq5rC8GubyiXYcvqarprv8HzEvWKy8+Ae05tTQ
hNHYVg1O7+aXpQxmtUG5jwziu35/I+DWcKasN3IR8t1yH9omDLvFdWwLLNyRD+qK
8ssvv6r9N14WCjZNrH0BlG6XOqAjaygdph2zTtenlgG71rUNDJpf4U2RaU8HP4I6
ijCW+ti9SzzQn1uRlcLVMVT7Ex7oZKrvfi9j72Ll27qs2RrIxZYOI/CVHECN2Xjt
mNn+u/XmDs0RIca3NO5/o0V3HhqGXpKbC0IZEL81lcroNJY8s7AAXr+tX2hO0Ewi
TpeEUCLVGevBp8Tgqt9LdDmjiueszg1E+/bdRjfXMxIFQlbzN72xJKXlO/+kBMTh
fMvTlTi+R4wpeUddyFJcXrexQczjPGGQPR0ehdp0XWXpl/trK4agwdMAvzTUSXo8
vGquqWX3vGLNX8usdncYAzMJAcmx3hStNEzGTGtL51exuVllrE56sMywgZqEbYsC
DdlE4L6+tKhfOBUFZFGs+vNZWQSrNEuHWWszUc2bRZkie/u+FNdZjQ/0PBIk9slA
xpGoWN16RxpctIcomAbmJdD5TguC2HOhNv5eHdG5Yy8JMOZSLZEc+rnqk0T5GeB4
ja9yJzHoZJAFGi/nA3GXNLOO70ei3CXLJuzWUQk6/ZbUjGLdVDAuSbrtrNYLYjUi
3dssO5Hl1q4jgG1qXuuJMHTPRgsg+LBCBLbCCEOWMz+uNwcoolMtYVVyieicdVTy
2e37eUXxPRnquEDfLrB/gJ5PlwZqwiZbIdIQmbryydxjCd/FBtzWGvefXZanxJEd
4z2EBcDya792IxOT53l2bbE0mhEhJTqd4vc9BlS92DKlBJMyfbyS2MA38IRj7DbW
YETJ02EhLfM8Wk8cgzS1BmSziUrRjg8Cwt2bcNEjsIR70M1o0402HxW9fmL43Lq6
mUHlqpGC0CQoRmJBOPIfMceb4vq+K0EphfGlKEjzbMAEhe7VCvInischzRkTfJIa
K4FIz9XPerGHNX4pyzTwj6xhdZIUUl6oc88TnSBoSc0vSCtBtvxN0ftHO0wW5oh4
OUiOI/PQbwYvkh4weqIyJzq7kEdmbdxzKBzVjVLQOD4PlKOMObqo1Zw+kRVQE0ZZ
hBzYQ3tpFMlBlXLdiGvkPuA0qkFN28lskCxp5rVpShrkJQaGv47fY6TUCGknaN3f
WkpsvxMPYtB44mVEcSNl9wCjmUvYwoxyJ7+BnAx/+7Hgm/1ORao+r++IVHicJDPd
5CVLXHyIvThA9BNS1s6n/QwwWbY4cEW0snrfJr9ouC/vqeGhw2N8JYhe8Aza1WSx
awqE2hUVKJGq7zW/pXoYAK0MqvTeSCAtxD//Zx5VPVmdVks3P9/R7M3vE4tFOGgL
5AoAkPCEQNF0qkc4Abh33Oead2mLyARAO1eTSbYjDVjmkEME0x/a/v7e+cx2bOVm
Fld1cpef0NC1yzgJZ/vsdutWe/L3kNjBmkuVDKQpfEbWYXMGYcj62wE69PZ1s2aW
psbHseX8p2k4HzOdQa3MBBz1v7ro03J2n6JzniSq1+jWewnxUhHhaFMCk+KBGipV
5OWW58HJRKQOZV0hH0ySpVoI0Icpn8wisS3aZapNADYgjeVgqhklQHCL1DEKGSX0
V5ac04JiN9XZMCQKncexjkBFJ7zbwBqbSQg2Xi/W8319IZt0ddnW0E7JGOGwvTN4
i7IMiyGllXMC1oqm4mvMxY3ZEnFdG5DI4cpiYK3OyWvYr8VSKZtAPwVeQqvF6+r9
xpcsx0coR8OhyY5PRrg0DqRyGUp8j0lZdsUO+I/ZLgObUdyL+sUcuuI4EL+fz1DQ
Kp+g7EUO9ddrq32wjN+l6EEGPlkQwuWyZbOO8JObwv92Upo3Q8nTzFNTFe83PEgE
q6qqCNGTNAiP67pgDwFuOjpPNhyEJj6K1NE0J9q+wUq7NFLXVN2xvDu6oziJCZT3
ZCiY2hGymkm5jXGQ+JiIJxQ/ZWplDi90UtiGLqNs79TPJKCLZGN9P+DF2sWU4fW7
iNGl6ptatRg3Ein8yQ7NL46WZTlxer3IEmN8bdEuElZ3HVhBN7q0EbwmtoiQLlcA
EHO9NDl2YS4Tfx8sXwLYLfLbYtJbzLHYp51Cc+hfXorIW4P0QMBlOMoxrgTZ4ufT
sXzB9FiZVGvOz8/zyyVqcm1fm4fd26arS+ngU5Zj4794l97Ii4lTEQGMupoYA0xj
bsGfOlfpywVtwKNK+Z5+bHWNccfoRChb3u54LyJwh4L1zEIsD0K4YeIv1v1jpLgU
E12yENUV5Gb1NawIX7FPEanWs6R8HPz025fhdKPnqC5kRake0oYOdIa0+NQ8emam
PvFKws1xkRa3bSIXdtkQFy+vr3Dom45vjMZRAv0j5ENsoOqEcdXAkegVY2B29H9B
qru+UvBUUw3hZQ2WosPSWRfGJKRCOO9LG1ssgQXtmxPLFPtoK5n8Y70nTotYMNO9
ODdG+3C00Cjai6/uDRlOIDQ2gIm/cF1eG7l+y/lHX98DZrBNj0QtlP1nXCtpikdU
igKEchUq7fQrJ737LhFeTTN2uksbNbVgweTxWjdphk6Yf7EgwBQR0gbo2HMaGm9S
SBzpFh/C0vGsFU9Y+MF1bQL4wzEm5y/touz7GrbYRxDca2IYpaxZnX7la7Lg4mTb
MStbIXYlZEPimPgisMYmfh4Imq1rdiqky3K8VvLimX6+P/863J4HrET7JYRJty3w
7P1eZLdvSes6SpZ9TN0og5cGu6o9H99v7XQdKmYmL1vQ0lMD397AgBUjyUP5gL+c
jap56y/3cgJb3UnD5A8yTZ2GHS1y3aO5hwsy2ia1LS7JZpLfdVVnpBJV9Du9iwEw
lyWMDYmKkGDTjbikZb4L66AalKLEmLrsGJYW3hzP2WN+S2z2CCeZabzt/NAhYzqb
mjHkO//O/ImHG4nbEq9RgMaR8zUH7MOEt5fQwkDrW1Wyw+34TpGlm4k2Vr5ulqrq
ORCVtCt9WW9lRag6/vbfA6nfVRt+NB2Gm8OadPIMGJL+E6577H3cyUg2I3vAEuRr
6EyJYlWVnfrLGCPesQXOzeidNPBzqyNHVhxaIRiKZv+x8wPX0lvK/hCtGZPl/ysG
SJ0CvE6jzSSGBT8jrmxnIi7IdstN6ldmkdNd3CqaGsnNC43hvQd1XiirxSsh7Xib
I8V45ZLx5C+Cl5p7svRUy97ciNgZPWWiC50dndLJGVgLUgveRDCNkOYJZGmvhGuZ
4KPO2WwwV8aji0HlHU76LZZwclTQyFv5CG8alX5xmH1MCpilGJXqKgaUxr2lDLoM
VQnWITi48B95OlBEFlZvD4b6ZIp+pmC993vGqBfjFT5J8pcuMwgDxAo0GkIOXHIs
yYEUcJAZ5lcMCQEAh5JVjc+P5nPTnMX1UtVM11YR2FuZOyfddrFY+3STSEgwvFtC
WQcKLvldUVfipxmTFy8Kf1+nbGn7DrGUklglq8CrXhswOG0bH/RPWqAvVH2nDP6/
+ySXE+74RzgJSHwK8gLFdJDZzoa2yF6brElq4IIP0yh2BES5Gab/UGFKOFSPp1UQ
896sQxZfQ28ytM4j/T0e50SiY711iDGkYb80MEnqEiacRF6tW9xo0XnA9Tld6Wjy
ZAdWlgwX+gRjrkGfakKWKSn0I1EuYf/Ht72SU/XHYCdwBBabwAOg7AhnfUngxlSH
21OGEbXJ3v6ypNrkCiSHiFO0ea/Nb7RdT1sFl2ChbBhCXieeAnoCELxALaesScTW
YXAEHT6iI1Z54vTi4OsR5B7NM8gYBcrqWQjHdj+wJHdPXZRvAGhmv/4Fc8gUIyM4
5Bgl2g1qiIvLIsr8TuV9B/wEIwPb22rBWhR/dtSCP98Zcd6LovvdABb9uOvTOHbG
vBWapLbry2m1KNHSzgfWWFv99t77C3juk+qhn5jy7A638pXj/wwwH6INAoy7+4kr
TQx4xAXZG7fFq/jCns3HBDbNQlmMuackaOTN68jfqUF1ntK/RHZgg2oyUBp5KKg7
NJ9EUuET0/GS4H+DGlXqhnxjfgxUNBxj7whwxzDzxFekw5pP2HZXeiCEfNo40z8s
KAlssRZoULZ7Tu5NSD0EJ0buEh3SeJA1sYIDgsQXqSXVAmxylvV3CxGAGEsC7RMK
Zix5eCuQWovxxTLbScli6t2nmYODJztzRgEuao8XamO6ReTVyUJ/Iel4ilr8q7Xq
589wC6I/pGB7pTpsYLAIPSpK46zgrFaMmah6rwsqvEBzDe7HutYbmOSC/qAfQAgM
ZzdCbqjWgcxArQ0uZi/fKROtvYu/t1kGWX4HWEwqzBjERMLXRZiI4V7i26NhF3O7
Fk1r6Pa81MJXot3e3Kph7Rk3X4gtvI7Hk2suEThMPuQk0s3kp3Xs0UuGT0Bl3Hyn
z38Liuvy06A/vuxMRcPAec59GkSxLcXd75asV8RfJwhva5n5sZsixkqkVwfQia8N
G3q8B1xEFJ/+rSKmeRrOUuvOX9y0Qk8odRYPoniF3R9He9ZB/nlf2eF3qb1z4LVX
uYY+jU3fTBO+1r47X++wDkTGfYL9qzvvo6CrAYmTfo3MobIh3H662Yv7/lB0G5Cf
9pph3SQTynRbyHwB09eNYdORTVk2MphG+IggrKx1+EvE7UVs/JpvFUx0mAVWNhCG
6cxTf6VBvphwIqTUTnpmbUZPE4NDk0p74X9SkOnheTHnLHKXrjrmwjZQhuLrtI3G
pUSV2EoJLUoqbvtS3CQT9ca4kVQ1bhIE1YI9xmiUCT3Wrl2jb3jKO1WtB7dysSHJ
ZkRZkRT2NXuCphBh9HxmadI3BZ9l61rhJzAITUSRetboP2yJW2BwsqnRGK7inovu
y3JxS30mo2zuGOgJV87+gDVeavC69yufFu44QzK5xg+ygJ/Fm+BWnKmMr92yn79G
1sdb0RWA/wceuMhsipzNTO/P/3IPYiNM52qjlJas2XQGNnwF0rZzYuJLGtCTwsxE
7uDGrBa80nvGJhRUEiXLOplj7Yo0PYQj7HaYwrhOJsulbD8nEhzeNGEOqJG+SSRa
VjkDmve+L3z1PRsLirr6dUokHBN9ad3BnADDDfTc+sU9TiUD3COJJHjCj8OqKgus
a8TrBmAzZ0f4NZZ9vXczhDk6J/teTe9vBG/sRNk0yx+W9frOu0fhlSLHWkg8r5jW
V8D66UJKqxcnQIYjJRW3VZniCj9TyjKOKozqz46nEPpvj9PSjKaj6yP7T9GvihNj
Smgq7jSaYOd9qpfAwDRzIxotjIB9yW0jFBkNpFCgebbUUXThBvg4sz/lDXByc3da
svnbDLZFAEMl40BeUELAxIcDlJ7+CNHbaTKgHcOXjfwAQVELneFZS+dowdgsr6Ne
hGQ1x6LRAqzfS91GrZZMiAaD2b8JYMc3X/elavpYix7cCAt3Prf48D5kxpuNH3ML
1R2OvRy4txq3IvhAsl9jvlwouhkHlWkWdQfjSi8dDDfbyIL2yS/G0Fs1iiDLtRTa
wb4HFOULGWwRzRLgksCAs3l34quiQTasaYNqS2oSuJDUCqSAPldAIoARMTNLUNkF
WSCOJBiTkvU8r3WJB3Qp/6vpFg/5zNeNhq2SdohEIMxd1I4s/QZUlq8lgxrg/2jz
jx+Xbe3wXKyiEqz4X5E/cCnrW4akZFK7En1b/6pJ9IMjbhKviDcphfQeangVKuAp
Msty+Bp4fT1foa49DCui9UsghmQ477IQfP0vZA+D18prn5TjY9dcZKpNXgRYNPto
EnxkUw3gbhCJnhVKI2lcCCVnQCmSRyRSU9dDrMBoIzGc355kwayKOxmQFoQJ65Q5
GYsWckt5FIPmbMj1WXXVOm3Zpiq0fZDqMvMYUm6VhlrM9FJKdih5DBQikrAA5wSf
fNo5JXv7zUAFcAjH6+KHbpIVgftjzr0S74A0G0lOkPyr7uR4Rqav2u7h8zpA8MGi
UoAKjEOkFdJT/DoTnfySjmmZGSWfENWNOtSSl0N+YBCf7aIGQL3hHJub+fYMmj8w
CvsIoW1QXnpkRXnkitZsRuBE1ni5C7CR8OBgix+TofeXo7/pWWQhE2DgJ0U6DO4y
Agmkg/jKWswlzdJOGSVDIYi+Pvay00CcUShVOAgCh4gFKQa+NOWagNl2VQQhRbsr
xWaVGCRaTLPUs3tIsqyLnCGNpIsKPJIRYlg9RoVzlDSCI4LNfnjES25RBIt6zSf6
oOQi1gVqbjjQ9X97VmQmiYUGvmQf2YhoZxtnV+RmY9T6nxJFpMiVmYEbDW28YGDf
Aejl0+FA3zjlM7/jz+fYLPc3IofHzkrA6cfoc48wzEyZWY5PnY2jJpdoNShPo6jk
JYRDxjKAthcID6ZnSNne8WElbfMC3KHHEP4dsRzpVmxEaf95Xa39mH2AGs87MfTI
UoVttiIKUyHQDBHJEOs5v7sURLUoB1b1JTPs7corkPsdBHYpgPG8B7nxAgZ7/hat
mebWgBx451gtrMk9ArDLNK0HukcvXXTUUrNA7Q47PByZOes1x2ph3LjUi+S7dmTy
TI8gAlNTSVPAPM8PA6H9K71E8rc2uumTwmlEoABPiZ0rnaziLaK7jbw44keXMWc4
qoLGBkEvJOpl7jhyPsLzHoWFkMTdfvI2A7as2IXU/CbbKESBcEIz5994dgC/sL0R
orcEUmFeykbpEY7+HsqoHc1AOzUMYfeagbTu9+9NNc2+ribWHZkj7kZ5CW64IkWW
togbv8deS2YjGMwaqM3kZqR9g0BCH3hcicrsS95K5ImKokfii0hFUOIVofWrnIwR
2xhKKlzgT9WenWV9N5vFObSm8XeBIfZEzudMFKdW6A2qIN28FOBdGxZkwYfOgLzJ
Pi49SQKNIvg5nXSEGWjW9d0rgivuPKVc4wQ0YfRESsAkS8qKApLe73PUzyn6EKB8
W89kz6mQyCITCypZJzTwByAClLYCDUgmL8xguumRM4bqjbaMBDRBMZIxaeIUeYlv
vItSbWIup0whp/qvdrOEKcZ9Zy0z6yF/nYgNmC2N1wraxnVD4fCsC/pEey7wIhGQ
Vdk1RdLi/Bbp8NOO1Wipxp3Nn0IeKIyVY/C6WZxZPnXfaGF+hc/7EIDWyZprJuef
1f1u1sjsDoqCecLge2GYhWPS7lW1zFZHPgRrJbDVMgZCTwY7cJa41lsoXWrD2HxF
ClO11WWO2vLkWqqkBgA49YM6bkjoNoPqCWg7xFBRKROHkoPFHT7CmZ2Xkb26aAmr
Uc5YN9OV2xHZiIE2MAwH+Nne9P5Zga/8Q6WDWPmq9J1dYho/ANp6uJxyCw7JcBim
LChaeYe4B9Ws4/Ooe/bETg0l3cgvEBBq7C/BNhjuamwI23d97szZQmYen6QLQn86
GEMcCU3SGXuh9z/YoQzErYI9rYfhLq4brxlaLKxXdd7Qs4e9Gutk5uIK+ou4gEmH
Fkx7bA1eQzJwuriilcZ0UUYmOYOYxf+spFwIyRWY4Y3dYtdlAJf6V6/rTO1qYxwG
CktNAJbwx1eFOmhnfO1tt2wb5R15wppt0KzMvLUSxhew/6O8jkTKbzjygzdmNwVJ
sos/az+UnPIEGMrSgI4rUIIQ0lA69Tjr82c38Jck8na+EPLeM4z/NEu9J0s+l/QK
icN1r0oCnBgG9qTz3W47BmrMrJpc+Rgogptr3Cqc7h20TQ8aylNNgAjKHM8Yiu41
PfN6WsItUVGCBhQP1gwa/ygTEyXz2klweoGXIPCK/rEAT9SeJhTjWxMapUSL+4Ce
OKMSdM5K1gX+uqVxYq4GEMAFhbL2tehVwMYxtSHVgtXufP4UturgEb2ntpRu0lJe
TrOfooavl5DhQJtbLthMDEVgQSRPb5J6/rfy2dUE94fLLMQLukKnHEy7juWTTnZa
uxE5dA/kAhIJmyhZHvp7GmK7ciQO8KO+liQLSYcPN7a0Ma9iw/KVTB7KBrKIwTd7
UYCOAd35XQwT+Uc/g90X9ySzFkmFdjXbHQYSMLY8cWpy6t4HXBtEryFiy/rzyXr/
Fu/yZ6s126YmZBA2DnmVPVd640kI5BtIinnk7JVU2KjEVrO9WEA+gSYKF6KYOI1i
nIJ9zh92rQgglBvZQM/9XoJKamaqilQTjRsI78ZejasSIXxicJfjeFkdTZWoAsob
O35cro0VdDQSn+Oh/szQjrq/uAUSOTft+uCClDyS8faBBjx/MqmdNEVfWxeLO8VQ
jMXkTX0VUKDYJ0oCcTKP/uaeJNCQHJM2dvoXajzQ8QOYDZ77uLP7+PBzWrK1H1D5
g2Qgx1juREHSRMr8KwStQ/tngGqzqsCmz8hBtsTTT+1W44bLFcYsr397POf3cxPc
C0/smZ/MAzRUdiILrkaOOr+/gL8FLEgoqBQwR56r/Ph/y/6X/Jy8iq/m5jncwKvA
95pAZ4ysj/7FTNktiDRm2Wf27RljUNdvtgBwctuvlyHvD/2nj9SDEz2RaftBiruB
InjRwk/1hFVySz77CRAIUL/1ZPCNEH4jjcr8NRyoJwIpatJ7DnhCl1cqFkmQYYo4
H/BiZLLL9l8hxtZbe47CHdQYOmtOj/3XV5pU92acx8ja/lXFWWHTDt4WSd3XjnYG
1KpO7iGUfSKdo+pCfa+eNyRlQzsHIVCWgV6Qn8fn7DCdtpjMnM3DLPSSVhfBKoXE
iIYjGVYjSYeGYtdlJAStoEKj6E009HUbCYiHDtPywh7AeFKL0dkbiZdkMp1BXKxt
8qRhpqR8iT672XR9ybq3TZ7Wz6M9sMXRKvDVtteLfp9m8/KPktHTo79PoHqUIw3n
7m9+QN2lHPQ7k0XPhTg2sdTZ2MmrAWz5J/2Ghd7puee9jB83KcK5IrbzL8ZZRCwQ
KiBvAeg/cktEqWtp+mY5OfgLZwBKtGyPBKcBtbRw6vo2U4n+HQ9sPWNpNLe6jWyF
JJZhRKR+1ZRMcGzmKGBB7+hqUhCchvpTiWP3SRoNho4LHqIsMsA7kBkpl72Y+EY7
1rWfVyxKYi9o59KU5aBTbdkwvmZDvcw3YgMyrleYzwPTdEdMlu91e1QySw/KQqw3
nSBWtjSs1u+H54UulLGwffm0VK/nTeUUPDwP+1BXvKgT7BhTtpxBu8Zs4eM7pviX
AhUUkThGQs5dHZe++LwXH5Wzpq/WemjC3DxFrbq80kLUVpiqKisZR6QIUnLIpk2k
HJ80xjr6FzmvbNfBkpc32qyPIXocvOjXti1V388FHljzmw6kz1sXGH/TQ37uAcCN
rEOW7HGYR/oscGKfPchryZV8dXdZ2HxfWiCgT5h3KSjBO1v0ssknZMsBky31Ze7b
wUymk0stoqFkM+zVtTncp1A3G6mc0kyaQ5KTIcoMxA9GUUzeH3sDSWN1H22hEBaO
JrQlPGZT7+1UqlpJO7ZZrl8fVgY6SU3hXY6Dm2od0EOUWpyiICsootHI83a9dAnE
v/tJ0cAtuR7t+j1WOMiuAbWyhPNEzRoWLXXzRyhdE0pWYksTAoN15mpaM6/5QanF
/fV/o2NCkNZoT8uhGuGAxRv2p9lM7IO7qhPz1+d8udE2o6NneVC/jXhZLf6WgoR/
trgQAgajCjFBJ5+fp955sZiRnDOzsY2B0IKFV1YqKXxf9O+LK08rD40GvMwMpkUu
yoIz2pXAKegfgJPWggC2b4UrfVFOkcPkYhGzaknzWNdO0sIflZuaGloA7w/t+kSe
AGfejXqXCdKBDYRyjeWbSXQu4r5Giy0rhG8fTwIUv5J23D37y0F7CHGb17efw0wt
qPNX3aJPi8D1mPkWw/Hl0i9eqoJQqQrCVDoR+TobVxP4fT27eo5+Y0g6PqbXbhso
GsUkQ686u0FgbkAk1luLPt90j+FS2nmJdy1dM6QBNMP91cWYtWKQ+ufuT4AQX5lA
Q+BmxLKn+72toKgjRVHrvSHuEmBX9ij1BxacSqG2Gto44TT5j1i3j97JBQjDyUKp
lotiryl+7QOYnCgDVjfvUrHuo0R4SSEWiCDO0/wbdbGt1GctelVi34bz3wnRR63D
7mFvACtBQBsFhBnpJyTGVJDrCw6KOlcsGs0tceiNuIA1DwVd5nMrdd2lw6rjxw8b
kfuG3Y787Dofv0OUpMoaEmbmLJJFfYCQE5vtrUnpoG98oMtHLnfKm6lq1VoNPNZ9
3g9nWGo+6GnUR+MVVFZ0V2nLV3iwYsx/Rs8EzV/MZbeqJbIio56rBIC6qRJDf7DH
eJcj/afVkdsjyG4IcFWm0UQnXmzLER4/I1EM2p4vlXxr1BsWln272e29Tnnv3IuG
fKFfFjdU1oT4t/GF5JnGXdCPu+m5GKMK2+SqAoY6uh++JsHqh8BhlXLGdc7uWb7V
RG6qxqqcdmG77loUDZRBWFIPUgyStCb+r6OHItxq+2lDDxNByOKr5FjMtogyWf6y
vFcrp8CsXe7FUegXIOC1Q4R2MJzJ3+i7o1e6QNNMsbIboyxuThSO//xBpdBveCc6
14orILTpVOP2jzjIBDANdR67K/D0ZD5XGaZClOAfO9pmnZIImiM8yks4it1r+Vdh
aYPKku3gFk+hY9B+3E6WSo20ZzIKrvvUqTF106nQtwTzOL32N0IVY0mNp+HoUZ8F
gvuA/+BkLd1Ba5yPun/otf9nj9dYnFLUKhG2IaJD8b0ELjVLLGi2libzNBIlkF8n
3U5hNyn/Hj7YFBUSyEhWCwBc+PT07UJKb4GXz1N9ysK67ZblDg2P840HRv1gtvW7
ANMZRI6wGXofCMlgwOKB40a07N9ibKT5L6lX/OEsd220g2znl/ZOxwfUc3cl9Kcs
h9+6pEGBDm9BxWSeaTvu/118UGI8WzgmbLMMfz/k8SQPqOH1ZYgCOL21X968z3VC
q9wY0dSnAXI1/Vg3CBUYiS85TGaZRg90WvjEvJnQHNw47BDheBjXFvMx6I+f4juv
U+87Fi5TisMvUghUDoscYMs9f43fG4BGC3/n2IYvy3g/47/WekvVv0VQee9RNqeC
8ZkdtdY8vUNzwt3TRjmVjDXRUPnI7fVgitIWOVP3+idhtDsml8n0TAOS8rtpGUoS
Q9yrAGxD36dUiC0SLdKn+CfABK5TsUCW+eTmBl7kUg6ozASt0Pr1nayI3/pFnzC5
sA7151t8rH28JbYP3LdbtLX1gom8JXEu8LR52Rg7q9ZDbIeJ1e9wDeOojNc/q966
1AmR7NrN4Fyk+fkHQSv/+5dH6cocFlF1jJnMo0+ABhY6Vcl6IGPeuz36Y9w3bC7b
kX13p/EszO+xkFd7M57IstCWtlAqSKG8z3I4u8OnmpD9/MC/rf6lj3OyzXYctAUT
+Eu+NA+UleLUToJ0mw5UbP+a9N+zR2Z6KQm3KLyMuQWRkxQBC8WJej9Tb9vgu7SK
r9vt4jd2tUFipVXu7ObweBgtDB1mMqQl//lciQnn4jxoMVE5P+/DFKVc8CbXnciu
v8fWJ8BhtW0rNy9BpTBg7UL6Ejcah7tvraEYeqqF7A++zpO118ZTjOdw2c8BK1uq
Viyq96IqCUqDDAaXWSXtpqYmm4tVeYkrC12/QNsjUkktMdmFXBMcgnbI5CxHdeHj
Tz1DlWNKMr9DImJ5jn3lDnpz1xwd019bqhKJn/tuCcv3COuRwicWNOkMXPaygwU1
Pc+tVnbrso5dMyBQFE2xzkt8XAfGNX0HVL7/TN/bwPl3qxoflFKlFLNx0Jwg+O0T
0X+LIIqS70ZCMJIB6TPIfej9nQPGZjK+6OunOOIbgaxBmTEeY0CT4zSg/DbhZRes
naxtlJNobI8RGxxsjHj6+Xct/rhJYGugy0AH1GG2S5ZP7sOqilRHZyi/5lrDj+P9
sURQTKp2rkjzXjGhZoacgs7Ffqz9lkWJXMdyJUN+kksw90KBfoecPgnDqOI9ZdmX
AI35FF01RM7GY8GeNG6re3C66w9WN64KU5BjZFPUsXSHb+HOA5vGFqF5k87U5gZ4
3tnHMkzHjjqOL9ArjG1tf14NWudIqchnkmdvBudT9fDVnOLI3jsobla3LljdXs6e
/+YJBxJpNxcr1SZK4Z2gKHWSEgJp1R3fBSUO2QmDDVuaTJEg/a8RRWTbiygXU9GO
qAOmyxC6688ajWVr7TdqlvnSCqn6P6/ClFoBX76cHAEhLPzcW2mQ7YIBVNAS39fY
5x2u0HH3pba7smcBlyYJ49tFZ0extgw/fUlhWJar2C6j91ASzRaeN2e9VdMIdqgR
vhzmyBQT+ltmFN/xnC4VMcb59I7COV3qo/BUqleC/+V6iSRKnmff2+QgaFBMTR1v
r8CsE21bb8BHHN4TVCKjWyIAlIHEBg8h+sjxQug9RqdMrB33KG8cxu0k5iUzQiLg
4LNQNwvAkzuy8vcDE65aUdTBQ4gPYCZDGsXYEFSi52+j34MVMp/qCIHONcCaE4jy
jHXGetAvRbCbVkYCMQ6f1YaP1f2Upc7cWJsgfBK0IRDSHn0P4KCuSMvu6Y2WdLD9
/aGwlv49YyDd2l87AVagRWdiMnmEVwRjPuAzqWq/OqPiyK1eqZgxJmbmEWTKEVOH
OCmjYo1N2Rncu8Qcdqs+UNLHHVSOfYd3W6hW2piNXOyJkEZORTGtVMO4a15FHGIT
znsGxorKS+9YVXlwBfTTtZqCtAna3KWbFSJERNxl4Dnp82I6Tc61XCDeldJ905ry
lXjBt9fzSzu03/Zvn6RCiwcG47PsD1eek1r144nHFxQVPaWAfQ8K5dzaToa1loEA
vGTW53FsfvYir64S5azdZHtkTjX6gopolkV/Gg63ApHmPL/sLjnhwVeurtpdbacQ
ppfKfc62jXH8PfgTYeAarprIperU7JJNYruCjh54bL1mXGQngAnuA3QO/91D4wMa
uCKB7g+e5ce7FSEfM6WnDZOBk5JVoCLnWayENrDwYi8Y9dDFJRa9cynKgRKnOSos
YX7FD/yQRa5+DD5b/NYj5uidt44XKhR7hj0yu9uljoe3UTMPtThtj+YtzoS0D9+L
CR6fubZhwGdt3k5ZOaH/3O261ShEOrdM0l6ulGCMQ/vYJjOgdoIie5jHwPQLfFFz
IlyCyUh1Is3wpAZEQt4RlSmdJGf7XUmyKevyd6NbL+yhCZjwE/EZxI0tMpmN5d9f
BXTxGc5rYgVK6zDmzCdPOvkq57BcnqfKes28Jl2VT4akXe07jz79vcqwJoan68Mz
l3IhJFbBcYiHBvViuBCYyOKLwsnP7DJoofY6XO0JcIoPlwpZvr7sRQkVmKtwrAEZ
wzKDVIOCKbQkU4Kyp0f4wBDGhuP3SwXz3GWS7CbZQpBlAyEO/KDBxjRSq/++RQ7y
aTes9aWD2HA2njK/pR+wstmGEo01ML+58Dz/7kVKl6JmXr8uKPRZhcH0T3EvwI1N
ACmYDB4tch2gIIFxJgGr8GWZNaYE+Zcj8TZScHlO5qu4OgUj4DDlU2HinVmZn85n
D4iMQQ2WVVheWOKjPktXi6sB/74kZldJtuOyH5SaqKzY6hanQBVO/r8kq/46Bamf
VWKG40Gy2RHDqd+WG4noiQzlQBDn8F1p6aHTGIy/XFHjwvb3yMWslzt//aAuS6pi
uCDaLjcCP4LiDr8mhto2s32pE5+NoxFgvWvECGy+qTxemVL9tn3xBT3KnTP4nBbb
epwDsTs6tdUFnVeER4cFOCnnW8wZlDBUl2Ij/Rd5hTkYz+RKuCX4WXLk0EaTC39R
5GhUbJjHlqtps3WIBLDgtYQbjlXWxi1aX8wFOQQ68+kgN5Utvst6YoFlHvweM5Ne
RQEkVeZ1/XFvL1yMfQI8mv2Yj17/T5XAoHobLeYsRhlVFt5gZ03qgWMTu3CZpqCm
DZYTb9wXWTL62/UYxLyHoWKozkNqJ6Iw0MIUFsl5CheCLHHwbVPnMAIQiaOuu711
j4XHDyq7ArzuTCMq/hRV4gD5LyOhrBaEiaU26z2jMqbvPAomOgpC4JYITC/rzZVz
KG43Tmiawrb84HggNGieDg3rIXKJtVL7a4j/PLzEi2W7WCMZKRDHzrxwRWh3UZNj
3qyJJkIqAtLT8W+wFyiaRJk92cBljsyQGZpfj6ufYIpXHh28jGAZfiPjb04BYLe9
lhNWlNHrr7V8xHV1wg28MJ/vJ8ved0RgLFuUpHKVBsn/dpiZbpLr6VlAu6RU+ZQg
0mh6MKlPP/BmNcyO0rfhVpNNibxLFsDs7F9VTntwAYD9Hx8LnpAZG0mjIivF2IQd
bAlv/fVa6uJofRlAQRS6hILMjqLl6nDYdKXCeyVJGxh2omxvWnQDg7kzFJNseAzG
xQ6HMw9AI663mf0O8aMJgRo6jRVpbBxKd+TkS+cE037X7k8FJ/pxCWxzZRUnDBH2
xoeVLzuS0Fonb71RXVAVNOGwWGX53DSL5F5fjoZwbZuMMgL6h7np+5c8Kyev1Wc+
Gfii1mc2ntCfE17Ehs6ZO4Dia4os0yazM9X4UEYbtQRz8mI0CR50HXRv+pqnZQpk
CNn+FLSO8UoICQtHiZDLd/cYiRYWAZooI0HtABkmQyqMXMQswEAkcSuOD4LZpgKu
d/IoGluNcgsEkAQu0f/Z48N5Mdtg0RTMPo8PtfErPGXBFOH/fL0RZz4rVorGgnBJ
rkCA/poauCCOR1YB7r8AuQZj9WG1ursJbNjIPDmL1dEOpCbQ/YC+Qn918cOzTJzP
CBFsr5ryb9ZvbzTgYum3jNao/iHEqyKJetCclcBOeg9JiJU80MoLrJ0Qr0azA8Ry
9RvsLQStwbcvbUz9yW3zo7gAHHdJoYP0DTjrd08UHfRzzv6f7X5gI3GcHgHSN/9p
3994Aii+vPjqD1/LaTN+3CKtQsR498DwouPaLRQbpNohXT1eUzZgIyex8A7DKDaU
x2kcftGtY5XR3D1eiTtn7TVLYuXF4hscXWCfm2yYNubvCt3dR0Cd9vK2PW7TTD8v
JiItGYeMyxjPqXZ3gfn8BzZyWPvWWgqenJw3wNosH5cG8OQfA4z/lmlBF6UuMPmN
+zx3bg0jhV9tvciycWRNCmjjUxjZIW/uq2RW2REFWxxi8VuQLdsB7YbyDpfe/QN6
231U/tkl0Qh2+L5F10/1MlBPPL3pjzm/3KFISsN2BolRIzUTqEiS0IWZVL3ry5i+
u+wx5vk8E7/3HQXEgkrn7UXQ3620OJ2O/bK2SVPBnoLESMcr8jZbLooeIBX2PeGz
tgNp7TkNohHMOCFFbLa8H2ZMw+lax3x6E3VLjysjcmMOoHN6EIgIqr7S+lMNHYXZ
9Zm+d57r52C5y6lLj+NOKUz3CzPHPTXW+8NXT5iVsX4Hwp5atNeBFmpNkuSXnuZP
o3q48zCI4mnGBkJqyYjNtSVkSs2DM2H8pVSwsssIpgSilDJdzRqm713JrL5hTmCB
2P8O1Uy9vtldToAoSOm8CmMYwn6b6OfOj4HcQYaoVzWwhSKwq5nLcy8hUumgKbyV
G0sBGEX226xU04SoSvzMrrUrUIayl3Vv48SfuGozvyTy4FlCOL+tR148KDulMltZ
ZEaEBg0RB/EMrc8XiWp1u5PWOCN255xon1oSWBfsDehzcqJEBoXuFvd24eS4lelh
+gbRalnlNCnCU++gjDpCxUDeOCd97ehbIAkx2L1PXKDEsxcSiV70uwXmSxqvACzy
jh0cvWlHhJaAag+JPsv7sZOvifo2n5o9RUD6xJjVhiEinSxuPxm788Sq9g2i8Ktx
/ExXm6Met4CtMy/R65Bw9ra8H0ECtv/b5T2QWrFo496sCf/EYbkhDNH5H3t6rONz
Q7RVtO8DpzsQSnfze+Lmdsy8FruXPuZEXJXnDiPP3OrVJLj4AarjKCjj0LQMSzZy
hAWrWsoXa/jqjjgakinkSY4OycGptloxIdJJBIGzY/lZMDj+dQvV9h3iATO1+Fky
3ZUGOqvaFY+2mpxATl5yNmHBw9GszBFTEVznYNGOTKfdfW7o0w7Joah4wN1tMv4T
M4qk5qoDfUqbYH4C8PDfSFF/9xN5n9LPGxwshl9qKT0GYKusFQW6rIWebuq4POU1
jQNVA6IjyZ44gUzxstFR5vsWEakWN+NXjKwvDTDR8DdxPbQzDYLuraNiWHtvDNk+
34Wr8hto7uaB5uu0yV480kGxTsXtS1GpmVByceC7kRCRd/Ln//7z1hmKtubV9vcu
f2XXC1iT/bGvArQfo2p6UyUOmk9Gp4TasG45draPs3x/ATZN2JU/7dykTWsZsX2A
y+QFAyLsiHLX5yGWBoEthqgA/TRpdcJOpAxX8aSQ7egnXVNlU8mNj4u9V4WW/NTI
kU1bWbMsHq32YVbyzFJXfhDYb+prFFladfrjdLxR8GPGsA/gy2JkSbJyvUXTyD1m
+rUn/qRo2GyZxDV90IUubFY3M8kb7RcTyWz2B7NRzsNjM/c0TIwLQ6yEyblDsD5v
zxPrRIPuV+sJpHPs02BbHHhZ2D4QTrHSiNW9rPpPb5YulfxbBAoNoYNWGYoLo/j1
mbSgf2m+LKEGEIOk3LOebTzn6VolOgWeV7u89vpLZNFSwyvdvN73BneGRatIiIBO
RxezM2Dg8tizUaMPqPlPLssgEM4gaFlcUsZ1oHVErpD3m3H+BTmFk263BjFNdtDK
eah50UmSrs41//CnanoLnLKLXAa1L9gY0Q0ozW3LqxCoekMuhgq/HEfpEAWgfebh
T83EA8BcunHbGxLe2ZJ/xfbPSn8kf+2H9nC52ZGEyP68uJx67+MspQWO3mMe3rUe
Q67vHQCk5lrrQ6HHaoJFXUapBJemP8JpS0F7Z7wpAfLON3yf2p7PMzHJAxOnidYg
p2FPl2RGXYVQRIvaePSnuSTfSpKOBpiVmBmICw9Gs60wWmvNe/DVAc3B2C4hAGiI
XM5ql34UcpFdCZpQJDgpUS6J3/9H5LcNl1PFxhssrgvilnNAdqMkMkFGSJtobST7
Bkt+rnxpbRlR2wdxxHsmQX67KzANUcywLeC0wcHP5Bq0AibCVdRhwAI/NtKhT6Wp
Xtw1e1AXuxwQ3DWHuU7XTVfE5NdsEEQ7KJyXAPj1MFj/hDS+bq4aEZTvOL3gzE3p
A6+DdsQuovUfcMQH2rNittnwXP81tihsQrF8waqkvhZltaFGCmjz1635BkBklsnt
TLXN4fbBdSu9N81LRRGHeZZoQNgL8ilTkFjuMAzYd0N3t8auiWQ4Uknyz0xO8ai5
T5SZbeFpeDUD8SZlJad2rMc3KZErbgrVvpba8+jqx4QD6B/UN7qG0wvec7swWw5a
HuhT1vUkbBA5kcHnWx5FZPaLHW1/EOZBwEiMD8uVWKhSc/JJsR1s/m9z8Igb2z03
kBN/Q/3HOoAVe0S5pofpH8Ka/xqNqzayZjHYF+SZUVEFCQtLuoePfCC5AChQDD/Z
VbTiEO8Tk4BaYrzi5NR/hBgC651CHdUTa+XoyNKvevmXyXpoRfIW9c2dNovsQBeQ
WKJeVFmmpgPfyyCZUUy3UXtwBIVBx1JsrJ6Ubu7vpiGbxI8y+P8UOb0kvjI6Eg4d
zSV7dpn+WkxpAOQGqS/XGayTfjmCPx06dvR7l8gSp0UkKNaTHUmN2RjowwcO9FGj
4w4EZKIyE4QamC2MsT4A9cW2AZiNzmLFNJopFI1DLtVigbr+a2LkSOkKpGthWoAB
/V9zuRgzWOcMaFrBkS/3MY8K+xxl5OXbts4Xa/GUjQp6YY1aR8nT0QNt9n0ZfHof
L8C/yEQ8fNRUtpf7VM7gb0xnmdCe91QhANJ+gDUQTr+oOiz3DxKc1EZJLQpgxNPz
chaVouTkWGaPPWSvV1zSF4o17n3TCnohQIjkEDdfxEWVxbfgbe3ogV3c5q3NM+qn
1PxMUEvaKrxw+sQmbU7DQjp3AqHUx54l134nrCsIzZ0Jo6Th5m4+NuQsU8HDy2O7
uke9hZDZMHM0nqtnmV3Bca2I42Xo2bdji/8pLPUVeoHEwsIodZfJH408PGCmrPaP
ttA4wg/W3Y8oTvQ4J1Gln0LlTgzDeirJykjFYArIL7bYtDk1aHUJP+xtpsX77FLx
l7QL9MglNZFOTBgzh43M/ydq+g4e/FMppdGmrXIqWRWDkG1cox64M7L+5S1mLG9z
DJQwsHR7mFWwUsD8RJDPJFGhaG0SIeK05pSgr+lWWy2KlPNQVEzAOpyKtx5PNguw
u8li0d2OIKGorw2GEvE9yhsSYNE+HFmQDdnVYAsfwGlJxcztG2pGS8ajTTtFWjEG
q9I3sJWoDm/1/snbW3IYq902smsEwom9Y7deUOPfBZ1wNLh1QiDHrmHvWmu2k8bk
czcoP41IfxTCqw6ZwwC/OMjzfBPTMZrOmBCpocJTf46oOc0nyojJEXvV7pQJK2uz
Mt+1QeaVDLYjW86zcumrgUSujVfAhlJXTYSWXCtp+MgvgNfBcaqreC0Ew1paFuL7
Jer+QatL81CUIfy6zimydvqkR+V6eofhIkQa3FNaidzEgyDa3dSKb3waqHckfJDu
zhQF6yWPc4hsuXHrgrE2QA1GhsHZixwpQNOHFB9dAJ9QknU9P6PIZR6VyOSYCyiI
dXHnpbAVkcjv6kdGMablZieZh94pAtTub3OTIij1BMlnVu8yR3HgPFQk+NYedAtr
Pv0D4ph/TKi1RX1DJbO6k3UHBFNr56ATkiNREtYxv4PUPvS4w2jVNSzcUejXbWFx
LZ4XodkkYOk1YjGKjHKeEyhJcl/RL+0Qmy9vuda4Pq6qyy44vlXbIoIezjnCVK5M
KUoO6VIKtoSeKJthJiV/o2joonLO5mTOUCQKOb8RcZKqYjvAxsWg3WfYXhjeNkQN
kTabZhNq6EINddy22CVOqIsIvkI3GqGG6DqzHQrqn16CzRW7YPS6fmi5RkmeQzHe
dHcw8FBlvYZG0BlgxO24XKv2Xk/zPlpnUkW9HFhfHZVavwi0MfEaqxx6TMdD58Xf
PzwgpA5zDH9/1GDUNIVmzXSJfmQfynWv6qFX0gQdgma18FWSOHBBfAOF8Uj7vEdh
Nhat8PFqmx+hdsbY4BsUMGmk6NYzFO9yf9gogzSIjaHHY+VRWDPV7LZl+GjXsS47
F2qjG1GG0ou1uBnoyDXT9xmgNz7f0uHNtUIb1tT5DPzlvmfZskUF4tw8EP5x4oDj
UMA2Ly0Z2AuaxcJdcvu9zJobsHc3L+zY1/6Eom1HVVbxu6fWJ8V5OMhUEFiWL+Va
snoFirVdRq/oemsGao1L7ci3qhfhL0IEMpD+dKPvn0nNt8q/nIgvVg7K6y929D3p
UWlZv12PbSjQcp0sORf7FRvryL+atafoVNY6aqNj+blOJtOCIN/Aft5RarFBC1rG
FUolR85QvGwptQOOVF8TY9Fi0agaTDmj63bqi5/qceT+gQ8k5Mj6moW1KkiSbALb
oXnRJiGtYHt4lOWpjf1QcAuGx49RiG0omH2D4BP9BBnXX5EdcEIZWQP06Z2cu0M2
MY3x2G7eELkCBFBKaZoAcfsqsxCKXn0nyUVWOfg+zyTlha2lqpCaOwFhkvx5gyTE
ljZN5qrOd6VeYXhvZ3W4AcnqXCrrq11PvtAdpLJRhWdZIzy519dJezMGSk00/NPw
5Xt+5X/TPfh6QSFcWtEEqFXmcL2AdBGXMklY5cabNC45RtoHuQgnEpr7YX7ub2CP
+tdnDCZNHDUuWFVoNHXoyaoo4P/h/jBGRflJsug75Gf61dWr7PhqXmK78n6EAtr/
I3MP+53DdlHcwC8LohdU7Zp22PShoM1ajfX5c54NCvFHByAVYZd5avpY2difLTBl
KdbsNbmtBsyPh72dBKDiWDt4TRNIUQnHACc0B4UeYeuq5k3mgRpWaFHO8GK/DCb9
/nOvZOqp3vBAPjeRfqZ7YSHJkhTH04afOF0kNICx9iChdJ3jGwvhoSbPDnPReoSf
q4tyB7EoEi1lCzda9NdrAqKX9J7Ysx/GXdhRO8iTryFFY/TLN2SQf/TjW4SKl1JB
vbLKBzyuQccM7u+rzq8S0SefSszh4jQMYzzsu33ep9qhz8BIputtcHk4sXZkN9M/
SHL7iHEf0pRvhNHwfCquuTT5Bo3M6u5O4sUz5uIUrB52IhkeDTQ7Jfrx7auXTWFu
M40Znv12302aJV95U7kFbiL8g8CM/Jr2SRdSv2F017G4WpBgYZ9Zte5I9sBKHneE
oU70DJZYJ1V3Nz7Z0sYeePWuWUhvLwZ6M99xMwxHfZukDjUv1EGP8Yt4Pc4xPxWu
i5CE3NsF88wNzFf7zF/7mNGLmLOQcBLGmCb54cbTiiCvXFAZvkPaKw8IteM4mvBW
m9LCN/XkmFmujHp9JTL1Y7iEIUFgYJRAnTlUo6NELqXATi9vCgZnb6H0mE2aAzWN
inaqyuhegqIWMhQrGGqW7M1JtB9Op0TSISj63cBlnGHf1zsO1wZ7MKk8SbSR2gou
w3qeG2wrDtY7gcgK+DM3HD4ttiHpQLgDrZNqvmdFp6lBUriE3PujweWthqMEcQe0
+ZaYsBgU7nLyd0OIsMGkjyUED9c1PoSpCEST5OzOshf8tY6653h2Pz5EDayO1L7u
f/1b10MnT4JI8Q+U8D36RzdEst+EMDyo/TaP8vLwTHc4T6xIqnSn+wYcPjJZpWa0
nAJeErKpsclLFUQYESRERWBvOwXJwEK3tfse1WcV3uhRt/obOHYFJ486jPV9J0uN
ZbWlY30bDWf8s9i1sEJzU9DdkqsySAnzPF/C8S5qtdhs4PBaRWnWE5hWdj9g3TFJ
BP+62R8yjlqre3ve7Km/YEMuQe3a1xTjYzfR4y7gBiz/hGWjKyrSKbcRyzXyXzoy
PSJm/qpU8bFhjkkOwfA0XKVnOWoRe2YCJISIO7frGkJCX14FhWW2gTrxqv9Rr7xU
myyUyvYnmU9LubgbxdJK72sY8lqG3QmeKtHk3rpwUcL/D3UQSProybCQAqV5IjR+
CFwfGll4M4w6EJ2Ftac6QLrKKH+aD/zGHzZfH9HD+d2SEamUxIgbk4MezG/D2pKi
eyGEepW3QkRN2zaSCEKftQY8hr1jRPgb3X6NpaGIfynFNmJLhetbCOTUMoui/pPH
MwD45JGyeaPKzkd7sjkcGfu3C+IEQm/UzP7ReirG/SlEWesXpVOUqfiebOQ7Kh4C
PkAe29jUVdN+02Cs3VQb/rYvrd8uOPGcxD7cL49vR4Bt4njYC+hdGeSzG4iudLgl
F0+Xd5YLrUZUk0tC7CBGkfXGYG706o9bEQ0K8KvQpkFymhJwGxGHmaU20eAIO0oE
75Dirkt531z2VeIm72ecGKVX3vgdp1OdO5i432ZIT/HiSpPCTtTJ+WPRxBQzaKGi
6h4D40WNGu4bJwONBWZAfVYrLDZ0S7/sh9hIJE4cXoQJuFSaU7lf460YeFrL+8L/
HwCQSwgNU0rCxuAltjK7ClWnzpwlmwuyqx2bxr4Z+CEjLrEpq6z12n5FW193rD9t
pS8tz3b8NCPzoHFytSMiZJ8nrYqqzcM8cjCb5Cm3QKVJiKMBD1LaSvzo2yave+Og
yva3YW2C+82YG3dZQuWu9UAyuCYJjtxwdrIYLOZEMCwoMNEimwEGzIRPabnJas+m
1butnXnQDPvY1Rhw7NbvFkrIfYnvv7de4N+PCYzNgI58vgomwQXleKt0wQpNtryU
E2mXVgWrwFnEiNChbkck06nMTA+x7Y4xXJkkfDoj/XcPluaFABAQwvG3IzncokhP
HhD5iA20eQoKzuSVb5CjZbd15JV4WKbmA+R5k5PnDEZTRY8mAscls/rVAcKbU3Pm
iI3O8nXQICJic1jaHdnZqn7PL3stLo7M6FYSJppH7I9OPbGynwCjKnYGbEiewhpu
K4Kqspd6TvsCAOqkYDUMf7w2Lf7UsuEBw8/WmmiqoJFDHQaFUUS1do0nIKfzh0ow
6eHC8oDTf1/VprvsfaDZZkOOVEi93K213rmuQVMZ084OTAEFgfeuvhedlHVg96ce
suIBZQdFNXFvSzNxY315TukSzRP9c4pKze/XUHRvF2WliPTKimMogghYQHX2eAtV
246Yl5mTX77Xqb/CzA94lVyCmTbtL9cozd5V8MZMkulaauYw6e+wiARkRfsfa0wJ
DYhDsAm4YgsTEx1MTrL06kv/0CO3j39TJw9eAtQKf/iCgIG9jRHYa0ahzDbPLNE6
tfzQCkPPP4w9XGjZ7sQIywt5GBpfWhHu/IiDSeafuQijUEzVFaaRIllL6rPkIftj
qoJXLaUFlUnvyn9jTHYS39hZnfIidtbyGXd4mD9615j36tQcumuY73rj5rFxCtI0
yLuB7oZWbByTi1odVOUsXCr0I8D6Huigl6gDoyFTLcBMGLhFkrnnu1acEMRAp6z8
BK5twFOyxj/5weiIKWUuO71rsY4MlgPLcTSS2IyNtSvINifM4fEEp6H6A3+8cJci
tjL95L/7K5W957vzZxr9p1AQ5nlhWw/J+945Z54czUTu9XSaly3H36u+onOgKuN8
lfsOnW0SvS7VTccVKgLJLtnh9j2E90PlWZCr2be90Ygo0peM1SmhxRfrtpuylywF
Mjwgn9BxUBlz3EQ6PA/+lSjxE3QlM85TyH2IDRMvej7iyMJm+l7lIfcI4qBkMcmE
ZSwU01irSJpfb+2ODhH+XaXI/CvRw1+niT5KczMBzWw0GzgdK/huP2Ix6NJBPz6d
n/rpA4t9y9F75gvS7ZT8J6JTz5Z3zP8ERpoXdM20JnZsx3iBu6+nzpuYUCc16q7v
/EJZSXkh3z/GYdlrxjNLrMNSaSshF6QRwfOsWbieV2DHOcsxg6NZU7EduxcpQH1p
2MTX4+YUKUKtNoCt9XOP1xa45BooZHsO9ilBRae2H/KiK+SchOOa2+LwRPbbZDSx
LjNroZhAHZ3XFv5lti5ccJ9PYGbMFOWfWkOJCNuEMcrzGMaXCSNqrJ7DwQ7wONqv
vXfi5Gl49GVprrx5onQRmF1Gm1LnSJGnhE4Cq/3SzImkD6gTJiN8ntRC346M/PEQ
SRbr7wxO0ZFsqCaGDWy1bY2UBb2s/p/oaDvgJFojA41mDVTbLowxX/082JLMyMp0
KZt2B4CKNO5/CwDgyVN7jzzhz5HqaFKFzo8xTDzP95t0tWSG5bvBLon3x6eB4Aa0
YKYGq1DFtfTCYFmoMv2fBtTrs/oLCoFmykvvsv8MpPnc79AEubL+Ky8BQY+0Dqyn
Uyhm/sqWLQnJwGW1z8RlmoCp8hYR5RS34eYECsvP7k7wso6c0f3LmCupY4F9sN4X
10m/76NojB3K6boz/T59ymz6plP2jCUIAvt95uRtMucMfI5yu8v1EB6VdPj1RERN
BUghplrv8WLbxuvpKKN4ag1mSRMY9RRovNZb+6Dc6fe6j9u9YXydSgStx9v2TxP2
eiXft+mKFbmx9Rgkr828xwmbbc7y7A0evf2fpaxIoNSKrlQy/k78LiGqA0LcTlG7
68i3g17FD5iHixO4XX9/NX/ik77SmOfrg0QTsj6ieFyA6IlQ4mAkfIJKYJ0g2OsB
IOn/Dov7i14dlp3IaqxT7oRhmshd7N85U6HWc7Ar9EZPGRJnh8rpcoZC86mDEJpV
DC4QTL8Bvlh8mxzOJ56JNBnVbIANHgXlHFEjt4DwCx8MJ16Z63jeTI8viKE49vG3
gPsuC/WoRsUOpIIBYRSa3DeV1+JK/TKj/SnRzXQBEJGNDHeaUBJ/Ge6LaUkwNR2b
6W8jFlhwVE0LTHmTMR8RnmcPZiOR2ghvQAsWIhTNvvD7qwjigYv64nZ/fSj4OwAa
Gy/Pd/j6W9SlFUML5zQCgfwAa5ogq4OX5AKjzVAzY+IblaIXGX/IGJJaI8UvFscz
vYcKf2sIyxH1xwSbcqtUrGo8MEq+2RekdM38WBFaJhLe4NZj/QV/ZSWlrDnqZcZg
stzKrwxl3djjttmdRtlBTnICfgl6yXjnrXqI4SufmLVmoZT6tVC+qx10PocVsC24
1aNbezR22Bx+HJiOhKzUfoh5ckXriNwQW+6CwqLlpC7tVHpcWlwIbK9PBOqDWdbV
kHEvB7oLWZRmIGSapO2tHPVCofm/qoRDVkRafGCxjfa/iwkV9UgRaDNCZL7no6Ec
EXfOVtkMQxLf+oRdSXjJJykETTnELgVrDs2QroPPf4cTSg+3KZKDwZytwZ4+z7u+
IS9DkH/ervzpRWxJQe0z3oUyTxCo6u2EZ6aHwtpHAq4asLZcIHGMk9/6R8t8lqm+
U89ml6r28N9vAvNlUOqOIWB3vIWGLqBqyRFb8jbELKh6FUx7aUQNqeFFhMvev4Wq
PrcMTtBpsOOG+M5808N9RmFjvcpDBBCYkVUl5afxEOO9lWMk6slXL2I/7pkY2rAs
ouOH9sW0MNnoJgas75ApI9HizyF5bFqGDyWu9kovm+fN4AxoR1/PjTIu4zpuYjwZ
G3++WREmZwQiWTfzz6086UBOkjF23H4lWfieZH01P5hL6R4y3pkWShfTgkXLIUUm
okmo6ArTv7LopmipExIDouE8houhUA4rJyS+bkX5Vw7Hbn4fw8VjW1tPfXpFdMw7
cAE6r1B3VRJrUj90glK4AaEVh3HUIL3Jt1OU+JHCCRP/mx2YCWOLud9VvMQoHZvo
N7kmg/iGcizjptBhyi2MxzktaFkhRL2ERbgy7OnGaYYbcdJL5BiAVJklSCGs4tsE
ixFK4NVynuQK7P32vk3eb+L7C90VA3xea3EnBom9N59B/23uvrASpkKbOcW+Ds5j
rYNV3PodKcgz0QJGSjmrgEmEHHjdbdcec2clKS+P0JfDbVsa5sEt7lr8j5Er/sCA
o1bTZTFgN6ymIXdLUNht+pzzo9sf2SDJw+OhENU57zwZIBYcK1qIBDFZ3LXxyJYW
BOzKAkfft1tTWtDvl5elZjEKGLtkAH2x927h4iEuyJBZUBJ1mf0zOoAdOnZKIGw2
KuJssZB72fqt27yK3VjD0VuKqILp2FEs+dwXSnPOdG2Y41xaWpC55XKpbwpDQBuH
PfPgKXuuQYclUK9YKlxrig1MEZIm7BQETCRva86T7dsYHnL201xHYtrVsnSTtmRa
541bTPUxT+eJBsN+YtHoFkYh8HhkskYrud7L6CTzQ/k2nXzwrvCAQ3KuXKHABld3
9KSDz0m6W1x7Cs+nFrZ5uwgQLdwHLfMgUqGm2GVNNuSxo9AYvAM4X2UMoq2uUNk8
1dchhDS1oTRH0QK/1/vPTFjfQTLjrTKtg3VRDtYIwgrt4pvUZ4C1Ed85xqPfQlA0
Da31UowhBl1dEDAy4t6kdLQOcflgrckKsRAdlQ9cpeEuX3ls3WhfyytL1mi+XhoW
XYiMgnKdAhhdFk1WJ+gRl77ZUjoOstwXBrChqcxf+ki/fRFv7tgB5IRCn/Jue2Y3
p42BEdGyqbhM/UnQScXQBOqHXEURmtOgLQ1exIif9lbaMh1NVJzAVKN3ivyWK/sA
RQCFpBYzaJqNV7X58ny7I2c5QdVRRcsYIreq8Jd1Pn83/xOo72x0AJQfAIve3UG8
BC3hVF6CJkk5ojEMdLv3zoKI0bUGarL/MYaAfj39/nos3RXPbYETf1swTbmluR2f
j4WA4zZ9emriyWdvE9B7Hr8EexFQcnce4H0OO5jfrZp4vOGFjhllYQKlYewjGJzh
oH7UDOiBPUmZnl73mGvZlz9I/wlmAx172veESAUbOvMMXdx9A5l5OWRPXsG0qftY
1lDFgC3VfsmhDKk/MPk9XkhfKAmyXH8Ze1WClPN5tpuNNfJ/ql/gD8X+W/V1REld
8EWxU4qtxtNLtj2Q+4vmmEALrRcVFwj1pso6R5rSHRimL7oW8RYI2vyFNuXy/XFS
pGKypLOYgr9PQ0v/2uwtdGANoTiVKW8hfQCPh8FvXeKPxPJbAYC/7Da4Zw6ExK2d
wWgBLl7VUWeCDemvA8uLLgfjq7CKLYfejO/5By7pr6tY/hQgey0TH5B5EzacCquA
dufWdaDvldrroIAiOQTNMdS75iA+W1hgm/Bf9VS8GrjQSJPk0vXtYnu3ZbeynC25
5Yw36fZuK/DH172IyoVjM98ioxZOor2z912b53L1r9GDqq2nwORNGMPc0100ExUD
/9NKKz9viLaMOYSx0fFpkxwwFhD1XylXgF0nEYe2J9TWgGngM30O4XJcwEkTbbsU
UB5Nbqt7AZOq9M+yppb6upkf5iSuR0nhFpVgoS7L9RW3bM5bUkLHfeTb8GxdO+a1
kpHHXXyGyL7cUb2udJI7pjfXYf8fyhCwVh5mLlkTlIQC+nYjmML0cZq4u8tpAukp
MnowirqlvxlfcnigrtKnsP+n+z6AGRFltioGFDhkMG5X2NVSyB2U+dl+5Qo7kXS9
YT6kGt2+r0LCsaRqBXDHaGz1Znsp/b5d4ACBOBsxFaFzwHc7Y83AbCAEp9/QMaRu
L0LaJuROvRQgORyG75EtBie6iaChysacBqL6LdIMG03hPHuiMoAEMENwav4rOsgF
53RWnIJOg2hBEx7RGEPId+kVgUbmsIe53UahICituiveKXA96lHeVNcAFJH5p4uf
oXmKkqltmTwJ8T6kO35IN0FBEHOAzw2jTXCoTuZ1vutLrD3BsZm7gQNLKGQlmfXM
mZR6rRR4+HwdbIoqac8kgvcQozycLhRNAQ+i6k5bqKGpEsm/IJnhk5NQQ5dxBU41
K1sTNzmHKeR2tASzroMUvy5TV/1yt+5GkWoROLoatjDeD8XvzA48m94XYX6HL4jM
tGqcRRMfUqschhmEK7sKDJmIh/PlYhU9HE1bRt/H+w0NPzhRqHl5ncOA568oCikI
UObkQ/Z+4yHv7THoaDujytjvLMdCnA+KOBvI8sIdjHK/hHqdNIMcHPsYOIAzQ/bj
Ix2T2KvMDTF2nvYwt0813MgGxGRlOX49tK/70yhNJ3A6GqH7mSO0qgF8N8bB05qR
fIWZR9RxLJQBsAG7/UvVgzHkE4YJ1i//kND6mLakyp7chxkDPMYtI0vHNsPG3Ceq
U4A+hdLw/LAWvwmNb/yK23lj8bvUTEUbwUhajYGBySj5NObxbrVeUctAvZp/KCP7
g7wSFFRN/Vxz9RvumYk8C4SCWcJo8wH7LLf43sKDaFplwSkodBTVtRTkSqo+O47l
wmU2GR2UlHCsK28f4UX3KUzHk0t8X5cv5a7c6x6MnK4fbvSL5fu6RFTty4HlRyn+
hu6EcN4/hw8sR0r9M6Nh67Z0nUJg8vDLzp8KxyKp/3ZjzDW7XyXZjorTbOcs/IZT
PAD9PKg/NBjtRELHvPZdbAslINSkk9SfMW2IEy7lR3nlP4fHGOKP6nv9W2TdIpSp
WV48DresiGqLELW4ZUXOgfP0+29hTf21vfbg6Ojpx70vuh9fgwVJgM4vIGrn6c2e
PrJTzXkpj9OqCA5aO8j9WEJhNvS4stx1cewawEqfQp914Ef+uK+5yv1WGD+patX9
EuPx/1GFHsizvI3P32zQrOQCPfvnEIgmw+1yRgWHtO1ChcpDkO/IPhoqlnApWkpq
Mt2+T2GAoleDW7rirNWOCXE78Ffv6+Ir34W/cSDEuEnBAjd/Qj80oiuf+jxZ7xSa
u0q6Uo71kONFhFTBQNAcgGTJ5LGVKg6swCpXpeUOTeY1vhGiOsuGkPxDCXZGcj9Q
i4NwbyuEnscaSkX8BCjmRGTuyeD7P70H7rp0qtQKqLXmndqHnTmrFd2pzglqlAM6
4zjUL2cLjdSmkVIl9NTGNw0pqE3JsEO7yTEogVRGI4l0ZadKeU85z/3ILs7pxmrX
PIVTzhDCovSoDPu+yy3oEEDM/RfBry4g4Zrqdmpy9w/muhbVTE8IiZ1QWqlnGGHi
Ju1QxGFVJNZOKytAG9RjznueSmHhkhhzstqV99eH8aNnmCSrckkHw12lZf2JjDUl
XZ5uq4zIGlP6743yy8Ee1OjwjMNNLEpM1rszlgCGdF+Ul88+9gfkP+JlatkkzuA5
qiam4zHqwcplbWOnosGGa4MuqhF/0bdEEFW/q/TaxZD7QVJXkJETpg+ZbYw1dNEy
ANoFefCB3alC+APGuEm7Aqgftx5sufg7OmQm6EAoWGbSxicSWVd0gC3hVdzaXQkS
R4m5pk0yOcXvG1wXC3A/HuJndfjxgUIQ7ZZpGbZq51PU/2CxOhgBnvWZ6+Rzypql
gpYEDgTK3vjU0mNss6wdI2Q3sPbMBDQ9eMx3b4OVhclBeLuM+cTVJfFaW19CHszy
6pg3b6n8vezrtCr46XJ1WiVSeuwbIJA0LihpuZw/JFoo1Nxu4ned7oPKB0Ts1t3T
T2qGP1i4GVmV6gnPrnwY1RnKxgg5DlFtRSqvEAct6G3LQ8IUKrQvkKXFsInggaiC
j2AdLvuGGZrCywgl3ybUnepe2B9nMIKg/YRW8npo8B/AitUsLs/n6NlWXMsos8ei
AgH+q0MK427Axn1f2dX5jevtaB6/oQnsmY8kBNezuoWZxi2XA2UQCKHBzymzHFML
03HPcriefY25Io2Hz40UnUJtLt/tr7GOmmvnDDaQ41cwDYYhKbYXS/sjUJnSNJA6
6u+/nWhqrnvga6RSG+AeJ3cClUPpbOKST9zuSuvYW2ISpMnmM4o6KM6kL71LH0r8
egBP1htbJnerGM3ADGGj7HeuMoqpfi3yAT+NofZZga68je5cf6k2OfsEt1CArPUZ
ZwSwI4bK+QDzRKoltR2L0/kf0s2d1LCZzBmFCYVdKurjsmffJe0sYX2xHsfYUOcq
39xNWEqK4uOFEUq9hlxVYN8ramWdh9JQ8qBv0OGp07jwxgHWaLvVccfW8gTfUIly
qHLdByp5mTBqDpaJ0Zyg3aS9F+g0stDgHfTmW8flodN/kSpJqidxRvehF+WBsYXh
eTc/TBrmu7PXsT/LWvrQyqeBTa3oRYnSoneKQo0cvvSlUaiAdAuYVso9CwRIUG9A
wUXT+jMuWiAp+EFZlKe0yPRW1NbiRN5q/T9N1KEaTLTzVtZyR2QfGcCrvGFE0DGw
u+NmJFIRAFHHnhBDWmhZJmnNycD2OfY7NOZklXQ9BP2eJiWv1s9MQjfeBlrzqrGE
QU04wGY5dcbu5cgehA7I93SmlyzxyOHui3el7a1eIKFQ4ua24oSakOc96dvz6bGR
A7k6sDFAz/ppgGbwxH5tAt98oe0obrGYASCQ/oSsSoBymOYxV4EwDZcktRNExwFT
2y1pYKVGz163S3zqO/5SjzfNPmCjwD10V9GVv2xZzFZBUlnJ1KYwjqEygrBaYq/W
OYChqNQd5ILZg4rn9Oe/+WIPfSP48DBfM0s0JE7aHL39Izq0SdbdKDktBqrjQ81P
vVWxrTUzZVkUCx/Ila57FU6av4cvgm0frA2/MUSKpQU6WMZ2JpB8YAYB+YYOzaZ3
GcjNG18btVOcXNRUtwlCtu+WBHlI3KsEPY/7CssF9dOtsa4tACas0fmItc9Vxkcx
HpShMCABZ3+3e834SQ3/OO3IuLx6AiMs/0Pqw4krYgSv5j9Dm6fBprHMkjh6t0J+
IcBbenfEzIBaM8LlwK2nxOxuHfPmpe5mYKhyEhAnbTWZqpxzvX+AWtyrnqHbmV3N
rBXF9rb5PpcKis2OWOl/nhjuCCUz6E4CPyDk9MxPEk5gwRmctI8UKqWmSVDhYQvA
R4ihCsoKCB7ZpFB608SmtxadWbmQJl1wD3Lvkpo/rlGw18xzLo1mLtKIs4SOsBbL
4UCfuqrhtx661TCjfNBPisqftX+CTXjx4/Alx/WwsutZdpQksbIRPRWGJ41ynWy9
FvaoDmGOes7L0q39uPeHPpTkkfJGon+QkY46O821Xgxg/n2q+l93LTE42FGnwCKX
MSvXPlKZCRsQewwVKp9WtK9gP2muqnDlh1s0Pma7S1sTE+CUEnS0v9QFAG+a0HD+
11sDzK4U4vcbw1lfWuONyN65LHmFKIEjjIyvDdo+Jvx4Tna5QgtfQa/B896LpGuW
oVzVPtEwuLzjLUYjsvusb98aODs28B/MuPeBWyjOk/ZL+v32Y4p37JYZ2HgNZ0hU
WETYNzABeP0K3/sCGq6VgX/TI2KdMxlkkQODvOsaMFhVxmn4xinr89Rx40GyCc7Y
tT/4yQ4+VtIuIO1lO9Ykb2TJ4zfpYXvsA52wNZRS5yyopG9W9f+BxvbzI0IJuOIY
NN82/a4lGA2+y8z4u1EW64saJIhDt6ShCOqMxn3N1Wiq4pFbIFIZuao1ISxCZwJe
JhCKVLbc9JqvW0SKZht6oahtD9XXReW+L45nVYvIrYWwVkDVp1Xyh3aGLJzwr+5R
RXNglArDtuCvdw67GVQ2vixw6naKqLC84JY9eIZZATTvy8qGPaL+61JUdV+n3bOB
Osp6WMxtZkPy+UmxR1aZOS8lkwnnk9sscWCHX1n7pZNSE2Lef7s821WFvwZxg5GM
voBDMepnHP+Dv7jgCOBtbYigXjKdjlb6ntYbnjjFSGuQtnxXxyUTbAxTWyVT8gK9
0+Ml22EWBryhGKwDNjjAt0GXC2jMJDNuGy+F/cjJTEAuV0/QDvpCSMYiskfXI1+m
h+yopOpWSQ2gR5dNFIhoyp3RQk2zDTE4UHKLPY3I8korgtf35rnEa0pXG4kyVocx
j1c3lUbfZ/Zo1CrfHMVx92Rdu7mHfzw8gRx/WiMtvuS1fMHpvqQSIsno3a8rGFjX
pNNoV7pnrxJ5+CN9Rm8z1/RW8U0vTSvd1jnNA4QPY0A9MH6I2hivYlsAsMgOzp32
Yikk8hn0q+PL7Otk4kHWnhSxtfk4UG15jirbEVCMtORZoYavQqrV08G5AkEza251
aKEQkTcMRhAsejIzKGCJksWxRloamypnCo6zmrBzeYK6OZDUJ09CcD9H1jVbs6aD
7I/K4nd5XajK0LQkv/oq2oKhaAk/kyWF21jeGwGrjveCBrNVe3HbBKsyIelwR0LG
AOXka1Tr1JmHu7Rb0gPC9cwgfA/hZx1A15i4X2GBmrZOPSgeAL4DBqHqWV2jAWvA
XzuxJDaQ3TNuhRzB68B0Otpq7M3mPZ48y4FnuffgDPE6QauzdPtQr2gSYBb4/45F
7Tu4YO4iCxYBzQKdWt+82nTYdAylPlgyZRU3KCc6HgI9Jef1BwipV7ijU6+8ooZX
XQBNjajTLUNRaPnh9NJ8mhiyg3bSBzgrN/EOcVzUxClqDcSf9vZKGA8Izd9vgHEx
oDXTXWOcIOdCRpUtSGdaSZ6om/9+UTmiK6QznHh2z70tzpaNhRosgwteygmyF6Rn
u/cBLCTZ+fWJu0mqQWAG5d9rzM0jCk8RJf8J4/v7xY6Mq5MiDXHpHfuAysKFT1eV
vas59tTQTU9EBmzzotMec9Nk5XNJryE8NYXITJpoP2F1fjSAACqwwoKrk8WasXhv
fi7ZeQ2dW03Up+6Aomg/OrqV6DLw/ln+dxFNmQk5IuJSQ6yk6yGQ7pYU0G62Ppxv
BGRLvq6+12iCRzGj1yIIiXP8PXvCsr/eLTcnXE6NnpiHqErTwf7Fdwv3YJucu5Rx
jIKmZpuyUqp7kpj1efDws6Q0BkZu7P5+B+4/7RiwiEj5eheLTNToMcrLdXnxL8FC
FkE7Q6boRnU4TQ0IOST49JncSUSu4MkropgQN72dTctcariHoqvo1f9pJ04xr7jk
Je7AVrv8XN5JZe+tWpuq+A0NP+p+ktELG6g41uYg2lMut2dFeTaIVDhFIkC6P23k
GoiRYw5jQNh5c/cqS4VrKuOyzCb+t8oVLTQVoJhpaZ41761uo+K069DgePxmaCk4
Fiv3qHr6IzudkBL/A6zSn8KT2iPPWjOR2gkxar26WJz+sxUagKMjUQXclA9JsHQP
znyEkArI5/58BuuBnC+9DZOTA8t1csdl4quuP6rcdmQgOzH6jTU7IbEb36VH4tgr
pNlPbegtvX9bsiJiwgW3ZJaD4pqw5kGqJ20s4lFJkSqr+0cZlzfERREuSgtZEiQ2
ZoOdAvv6oRcpsBL+X138UU8/njfZy62f331u5gsQ+Rd9WgqLDbPKBPRtLULkwXra
CXu777RbvBXGw9yjKhLEokIPkZ/6zr7x+Kw9ueUaIjKQK6AkwjBlcVGB63rYNejW
QyKOtkCgTOo07kiDLHGIQt27sTSeplErkOEiMx1CGup8fIvxQzIGCiMG8iFlEFri
WVVu9H3gj0zoRXL5gesLycx9ZUDihSlVHiMW5YiLRk5qD3DwIXFk6Ge3Xh2UWTSA
bESTi7n05CRuxY7/dc/n6BK8VRl6euToSz3QJ5fFeauf4Co1wVC2Exn80/DHt73J
ZYXh7AWCdRqksA+yb9bn2+mIEv6mVIOpvWSf3Qf5eCQp/QeAOWCW1lCFC+yWarlN
AAFBgp6p1AYySwUby2x7UGOvV8jDXiAxJX7eU2zHrflGunBJ4W5exA+MV7oWqVMT
xRklEiQTNS+DS6RMgpbuhKdliMty3qA5xiQZg/fCfFcogOrF4cQw0pap8qyCZz/0
3CfL41/y8U3bXRdbCvXnpWnHQYmRTEgBCeDHy6tDOGYVtzY8THMAigZIY2+Bn/OT
0XcTOFqlWeaTFqYyZOb0HjhtbKZ7p6W8ekkw3S+ZkyPoPibsCR+YlcgrgLw2B+km
bhX47YIkIkQXjookg7kEbRAl4kkYexAspwchYzPI5ZAn2icE1nOQ2Q4koTMN4JP6
eX+OImH22CMBer9hamMNGp9ruVuKgBtFDgnuDeFBCLlMIlW+eUaXuVY7jvhyCw7X
VwkFvmQvsIFxjRcFQ/uQNEm610uk6T+GFmZIuOfyPIf70IKF0qLZTKzz5W9Jabw6
h1S+AT36g/mSZMJwl+KzzsO0AVJE2uGLvgCMJrPojTzqI6sPqDJpw5gR/Iu/72na
JOg3HV2a/qCy5br0PrVqxk6NKs4XYeYYzonyhoTy+U4cc6Vn9Qg4le3go49Zracn
hSLDdMR5S7zVXsjR3ZuTw9buR6jzxMYLdw0xG1UjCLo4HDGdj1k34Zzxop5A6Ov2
4N34m62ccIfAGA9L2cCaG1ug3LphFLmdDjUtlg2E8a8I0yBrP6A+0AweRxbY3es3
d7+ukPNvp88vMVLpsrx0dI7wCkifRE7dxFBTr7ElBW2M+Fs++f7qJMGKoecgkGJE
kf22M9bO4rhyAREjADEd+BdTc0ZYQBherBwFGGwRiVCgEPXafIxyEyZ/tZ3M9VSH
gLTfJsG9fx8VuDPKRQnzBBnAFpGIjpuWHle/U9TpMVwWx2QATpe86dpLeA89XpKQ
LJK12hVwuOXzEZYGfq0MwzXBcPGfKxFXqCEX6PyheyZX7eVhI0/fzCXHrsmJkrKh
V1WYkGeyZMMROz8n+UWm519OAOB9FcfPWjpiz3HSNg6ezwtAuaDHlW2eCFCfjEKI
G+qCa07eK/ylTTX3qxm5dYTwkY97LE/KfqKfNJ/2rEqthjS18dV9c1C73gSyu3aw
2sEHePRSZbaU5PJ4PWbW4jBEU0GzP5JKwPNSDD0Kr47OYynr5rzuTg7R5XsuRkmk
v1Mm3ekpGNDxJFG39pHGW3MR7ia7XGru4eQaGH3gVuzFxp9DlW8QXMGLOJKOJyij
vgzhtFrzw7twK2FW48dd/rVaHtoz0tZOFcIk4CFW3dqIZTtEeaDeyK6rUvnivujd
CU5eDV0Jfka/LhyDsAXZjSeHhrydufROkqpv2NnYEVLNuP4M5EzVCl1oDT0/k0ou
EmA5lUHmK6C1mX1SKt2b5pgM50ex46AfYpA5ZTnuYSo/hb4DBZfjd1hgLtjqtkRN
J8Qqm6etYOyblfknt3LXFeBV2jeE8Wp7tlRS9GonpKTEqZOQ0cX2t27e64giDYb7
j/jsXz2mAffPhG1qnCsLlMAd/LZDyBnZxiQF5ReQkqN5GybgL1uROE9k3gNMY75U
PMWAZeLmVP+ZDGUGT4E9nXxSFIYN8GGy4PUOHEpyhSymt/q2H3LRAbSnVuqNrhRD
QYvdQxZMsNwPiT2O5ep3MzL/boppjdOrF962XAdmncHkXlYQV+jtjGhpKdJ9UpWp
1fTKNcFqWZrNlzWCZuIagMqax9Wi6zVkTiU5L2wjbe9ybN7cSsC8NFwUfzmojFDB
EnlGT0h4XQmmmXsK+h4evjgaGrTUgkIhFHohRh5MYA9D7aMxGB1Fdh/AkeYRmI5Q
1v7plVgJ0xP5SQBinDstl+fHKADGf0JYfsCtfG8VNScsBHEgUxHH/gbic3wg4nrS
QVSkK631pV/ww7EmRO9oFWgoKgvhctcGv9oqHjL8MuzB4QGLRUofS4x7yee78wTI
DYpoVI6yKAF9O0bdvYls8wpO1BF2VhL1C5yWNO8DHb2FGpZrNgeCn7Of92hUeYxF
+ufCYgRPMtogTmZFPk0sAxaIWqGt3OTEnJHiInd+vZeFeP66WI6bPSJM+EMnHc7O
iJUmrbEZjXz6DEORbG9pqgK9+XkXFkJGHfR0ZoFZSEO6uWp8bUS1vzWn2qSL1Vf6
S1ZW4eY0BEnwQq5qfu9l8DopBhHhrp3IDILZzOQxdIVqC+pydXJd1CBU01zyhecZ
2atJu84TWA17DrZOHeXU2YBkZLS9pD2OVsuhNFyceyUogN3Tif1e2ADvBVtNqNuE
YFrPAtJI0idYPG6eZTpfh8pIEnn3lQ1+YLL3l5fLqEFu/4maGuNqx2LOl8/BAW4o
NArT5b8bmBGouLPhirJQBUhZjKb6KCsrnQyHVu5qrlFog0mFIEODDB5AVcTlrFj2
BUF47TiV8O/5hGHrKTMZEA3pH///Q4YNUzmoWtehVlQTrujzcgLWuoRRehXoN+45
klWFDVcr3ihI6fZkVWguM2661p8CF5kLenT6MyB1Et0wnzEfHxRUfZqCCxPL7O9q
r3DKBu9SlVgDA8ZcvYRcNhY9+alTeSWaL04lx1kiO1u+wDClfmx9qrihK3AZOjZb
WCJJKGREANQ5Iu+ixcT0P13pYaQv9ESx5GnCC6biFjo2kULZNrG7FVdfaMY/E7dU
RKfthIVDc8DPGTgiVDpvkDW7KGFyoxhJua8U4xiupKYVHyfeRgAr4fvavpiNNNfU
a1gIzyd9+I1MNza1O8NzvS1dZ21vCS8sjYL+Y/++OzH7EGdyhRwIO/TqcKcm6nR9
03ocg2cdxazrMoOYsTtCLsmt48l9hk1AL7jy2mtdFj2k0V+P8/x4YkyEmevC2xdY
L59xGt/3Iy/qbDpE15SCwWXsQf4+RKW8tzs/acIU5uTFps+U+yDRV9YOuXcN7jW4
yklzhadNJYow8tKHYtVH4eZVfyFUys+1d/vWXC6XI2z8ONdQxopc1+pYm/29kqA0
K9r/yn6X4cpvU67oTQpsOIPrEZrGHLEpAvuIsEIHLnCPzTKmk4jdEPUtjrLxaGch
Zns0xhG3JN7jqtpwSmLqMG/Ue6is5lZ0xuwKpBrMcaZpgg6HvtVC4jOx5smmb7Qd
PvLSY0d7DgDA5F9qqFy0Vj5I0+VpQJPrHjII/3JsH8wmnR2HSrm90SF1cFVF/HqN
EGt6DuAx4bBgkU9Dwv/rxYDirKkh3eMXYvhWF9agMf6uzi01nPHtNJshr/HnhIXt
X4kfsC5Jvl9FJC3M2lKnFaIlps3VfQdp/cmcLMK1kSl2ui0mYIqdGRwHtGN0zDzE
LhBkFEF/mAsJoufq7gJjjCi+Gngy+RiiycY4mcyhzy6XxEYvkrgAi+IIdGRWc7fw
TkKoQgtUOp63enKiAthxSLYVWo0HIgtwhlayJxEUyQfAmR4+QMbGNYsY7YTwUObE
A8RVYjOmpc4tRZVcYFRPRYcQd51tJnRijJ5VS0wKwJxcpi9Bq0s24whGzrxuXdPI
9FxfoNzko95o/U5Zuv0eLItn946P6yitnELNMNHAu/ugTxhrgdAxGgy/AghLiFQz
bzHCOFxk9SiOHQPJ7Yv8sYOA+2tiUUJS0Z3o30MHZ4bTm13N043JlfmzgDcBubCV
58TZ548uY6lfAanOe6Vz1qpkpMk0zuds5W7+1/shd6KoIFHl4lzpYz/uulMkXlUz
6mF88jpJ88IhSTU1+WUTsAGaYDaB9ayP/veK2G/5n/Y5oIAyxCZgIUmfQqGW5xdB
Z+wQg7g/YqFoqonRSQY3yi/HNTWaWW57JSVyV+yfL6CdVqbonHO6qjd/tKKxZFCm
YF+lxY71aYmKBV5w+ylofxLcGEL8ZKyKhZYSbRaWGprlD31HYzQpjg4lS10817yO
/VUqzwPo2yfevS3SixjKwHIjVqkOc2NBGtr46kY2CofO3vhW14RqLN2dKod2UNzv
PY593QKzYu+3WXiB18BoNaXqZPurANRfk/oyS6QhgQrh7zU10T/d6sVWUFvcd7un
u/H3xAsbVO7iTBrsgp7HiFuZ/of240fUFP7Rk1zx5I4GwBt+Hp5tRaBB//uXSOkb
/xtlUghZkQktFKXK0PsSFCwWjTwJ9AUOQ61xV8VOzyZFBybYZtSxmNZBBqe0EBje
RBYF3fZ6pX0HJOUVy0QlWaJcZrgYEmPHSu4ZWnKY+WG52x9XtMJceIBtH7Tq56gp
9F6V08G2j8GEjbzeDTYF5EE+XVcHmXAlR0UQukSEPiozFHMoYx0NxW42nr9DyhLi
15XUIBviT6QvHQVlMIVe5MLQ5kCHXCjux/GkFo0dqeBI3baN5t4ohfqlUv3zxt0m
HmdFy2wocg8uYB1OR7aEKbDiYs944mLX0KhfPhYACspCD58rKcbiGEgYACNrzFxU
Tz7sjKjs8Mr3c+xY14pdZyy9oungMrpkf2XjJGjrE88ooG7SGFOKQ4PFbrMVTZ+2
1rksR0q+52eNyc8nUQFB7F2ruhMHOfgyMpngbcZRHKxlbhn0BtnPPsVw0nSb1J7O
ehFSy0InaER0OMsb7yFa2FfcHzvassSfmzOT4l0tTd8gwkgtgI9JBEVFcLrtUl8z
wKl5+MJ4cjgEjM/gzYdX9+DwpzktRMENFCkISQlx8NOv0WWJpeSoNuGXmNMnDOOT
vmvvoBefq8eqCSEBtNGklsNDKtqlNgDEg/iAyQcHlLuHRu85fd4Ilgj8Td0gZEKh
60sdRFBtgyiLUM9Oiay47OYP1wIcjK6oZ4m0r+G+WFczwTAcap0LmML2x/ncJImL
aHJHQJEf/mclgr3xvCcjIvDNqb+cQTHECdqGJL/j6Hd/9qCbqNRQ4eBIRXB/ZMp+
GG0ClpQXE3tZMkYcFXyppPU3SdPijU0k10nbvYAN0chpyyvQgxcUWRGp04SqCI6s
Ewbk933dSWo238fvqh63EV5/dI0WrYl95NH6lB+ZDH3SKl87HL4xP5+5bW9/wVBL
HjtFcRjAsRqGLF44YyQJfyJTW+wXDnWNLHlEaHU4y/xVY6IOsiHObzrb0jJNiKil
Alh9KMOjcyX5ZYFYjgC0YN7ffqbLBf5Xf6k7n0lKlx6x5cKGub80Dm8X+zN4HtUr
O5UXR0XxPs4bumc6Dnfk1SU8TGjxP7Vz1o7M+wlC4+M2U7Vgsl/HD43uTZDFPZGr
M+6jKEV/JeIZI8RFK7ieZ45wWfgRue4oWczbjOUVX4amZDjPp2ICZ8Uld5fZk9D6
4hOAIv7LSqU8aNhqJYkFM0Rv1DdIV9HlHmXSE7NpwqQ4oW/ErqthZJBEfKGjq+68
P4lABCUgV7sCTwWmZ58scIOHypvm5BEu5POaLoPK5RE/8mqlSEP7tgqIhQ5Er8oo
ZdCzK8ku2nMWi1RGDUYn/dL3D6DLqGcDDbKJDFVhYbb2Jx6oQU8rC9eviFZqtxiQ
EPpKKg/16QJlSyiE3OMp6bQxTdBxQCRj1NfjPVakMUHdhneBZGYTZP7ZG3MvkPv8
4JIZFrYGo0MJiDV27cxntmvvuwu3NDSbFb0MZ3r1ZFIMltpO1Ji1f3cVeCiqFrfp
OBFVETnEfUJ2YbfMNbHXHvgJMdvLz4bVIguQcnXDVKSJpRo2E4g/Eje3R+m6k4tm
3qfoQjGrxHesBtk3stG9a5xwVK2/jxF2fEg5DRLiAXqro+/Vxo5sk7114tex+GID
QujHilQbPyM12mp2DDYCfL98p/l6seHEsR17x77HeFPF/mnVB3zxMyPFbYGvQivd
MOd73gOBe/UbDO3LashtAfz7JWzeuGKOwF2bKOc5Y7dRZx6YuZzB8KHI91mMVJW9
oZU1IbPQ4zkaMNdtxRRmVKqMYas6CCQld+LOUBqN4xnKwEL+9GK865Oszhsuamxk
i2ENmo34VZbtypyrHs3lvh3kH9h61V7sznVziN8wddhJ4kwp6/UIgc6+iXuIzvg+
1W+3DpzN7MedDyr+sKF4EUsBHQCuVBpipPEFpdRZOIRMEZUwXfk14dkcmjJU/ove
PkEvSHN7Qa17OnEbD0g+8m14U4HjYN+Vu4fyH2+P/8FmTfEHZ4aQftuE4KhzrW2u
IGUE53KLBDl9/lG5FEtPdH6c1W0mRb2xy/el7jhIicTCIiWsUXmeNUwF1Mg0ckKP
81VILK7Z7F2NzgYHb/wa8dEups7/VV4yBV09jFNZ7PPM3oaHAYyGt3ypaZnTFY0C
V6UnV541vLjOj/t95I/tvlIT91GNVfgoQ0RRKLJSxMGECXw9KGJKDBUU4wz/BAnO
kAOLDwUQGicZYkQloM79qZrD7D+lPPbtg8HL+GlsUwYjOdwmQepauLASRdvV2/CA
ciu4KsaQ2YfisZk+i04ckBHlQjPMG0kDGyuAvrmPqb+9gBu+Q+Q1vcMW5Dk36n+l
J8VZWK/FEPf70mVujRcR/FPLdy4oC581K2kNdA977xwG4cIeeUqGpDNjGLr1Jpir
rdneZKVe6ViW1BAixFUjoakWIyMTpDile0BshnuAuq6aGynRp9rDQjNpDfdERYYL
xY+vRxodBTvb8lJ+z068B6Qilpwe93pGK5NG0DUhi4/2M1CU1hF/t6HWrmtVCwMK
Hnw2PbgXbdug49u/VhKPCSnDoNXjteVSl1guPw/JOA0Y6fZR+C596vofa3UfHv62
+rZ5R/7mgWg6ik0O89meoqQTEItqu0EjuLYL1h1wD9B7Y1MphpLyzGzcCpNkJJfh
AF22V1yrgwqkKKA4kINdRPb7bCL1kOU5KT9YL3QedZzddX2rfmOmS5N6n8GO4aLc
/CChvxquE7zc2K3tBWQ15ut23CV65T5qs4ADqIN/soyrM4D7ns0Nn20j4oBZ0xtQ
NA8s0X1oAnUcTuy7A+IxLi6w6tLEtsasMju9r2p6JBX73Ps3I4GyMUWtkVSvPElK
0EaBe3pR61mvhZoJVVYQa88TDYyyhgcj5UwajfBnEhWCyLgaXt5JOngOMMT4a/1v
36wIO7lxMEn/WCAjb8COhRoxmFLks7/uE5VTvCUOGfUg8ggnT7zM+x9IcTdetMbu
Kc2hYjTn0y3VL/jVl0vMrNgM/abhuaGrHFV5E93O543NMFkMYulbz1fKroYgXMST
mf7XQkAf5JHwQuZMwaQwjcJwbJyH0akfcCcZose0juwwe/cf5ijK+FBF/e1lvj2y
iW8cVeJcTnqskjmfkG/8uoeB6xsUhstkUWOuMX18UlW7YLsSpjDoqCMJCrVQQzcO
a/u/Z/D3Bsja4E73q2vfc4sI5/9xrY5DtDG6roTSllOEPJ6dTjOw0L4Van6aBlnw
RkXyghMv5Fv7u5edBAE9oZaFTZAcA8HGQ15JUV1S8JxSCkVwb91HygBpOn82Me6J
D/jPiGJo3dsd1nJrL+jqowXoXjSbowsK/InNTeloq3ZPZQ6OSg0pYsJX7+SGPISk
rvyhDW8OHbipYzTzarzl1uf30RYYDc79mjpYDPj9TsobCf+vb3ksJWLicwaRdObd
XBqK8X1B4JZh5Sm73rIqhC9QqOrU5eC1moOtMF8Q8zRlizcZ9Mvjn9b0rw/KRgm4
JtIooJbYe2Gw0zZCSzKYqPR/D3w2M79WE8q1STZw46fM4VP3C/Fv92Us7KndhFMF
fmd3C+xo08GA6HzXrP1saJvLHa3d0qrUL7dWzreipkR48D+Ry2QXmWHw6mrsnI3Y
agdME6F3CDLdE/N8HsawJtJEU1gmtEqP2J9Uu+OFp77YmTusjKNRRlFTucjKVn6J
AIa3UqJPevms9LOfsrXtnsCueqRbpKVSv87/4wmbGSgeYEk+2ZXVNJcX3+dqkNYM
gxVjSPl0G6CNG0xtEyKm3q06jtC2r/xMb4rHiZpOOZq8PBHM5wTnt4mQ8CcJmku+
yrcupxxmFZJpR7sERqoghVKAa9mc894uxDgAo9NvGWEXM5DtrZ570IHuhHRBID2O
AqUn9qkMVYVZbO1gfPOHWyVG0yKm4JAY5ALJca0qgOVa/ASYNc6w3dsnltGv6DYE
MgW1L44Z7fVvtvwgEqCWg+xRa6LN8Mw78NIM8z9kOxQEAM+yqJP9Tltco26tLVlv
riiPm872MBVB86meiNS09x5/Qngq9GsMMRsWoie0GZpm4nHFi3gEG3tTe+5KApPH
vzgPvdTuZB05S+7b9y0urD97L6FR6qhvclZooAfgIvAgxDPy0+LQI5E+ScsgQGmK
OHUC4xkaYs+MPy0+oAXrKIq31kYPy+GMGVGIyR3CSJTu8BSQjGZQsYD3cEszbSeG
ZebIQjrWnE6BVSmdUWingDpm0VptQR0StePDxXqdajf6Do5Xc2ntthObywNnKGv/
YDyGaoMIurljG70RHZ1QFTT88b383upD+gZddzN4seIWKkrfVYETxdp8VWq0GZti
j+Jji4BOrrY4z5zdrr82D2z3mtngxrNDd/oaIuQnUY3TkyeMuJjZWpnb/i/Sdyei
jjCfk5su01bRIrF4pHxCluBUkfqNhjvexOn0v0NyQ2Zg6hjt66/YalyoaOMmI/oR
dhS103vyyGlP8vFJSK9dshxok+Q/H+cEg7YPDzrfdambV7KLqrdkZykUqTncc/4K
9N2Ed+jejYc59f6GC7yBptEfuussZYR6ld3pfxHcy5+KvXP+yJtVCfprYWkiyBgd
HMmiSJmRKJM9bn9zgzoFFIV+XDgrKDWYuUZgewu0uJZDwudd1ALhT7RXYN9W6+ZU
Polpbz5RTkSN1QUCndk8Kug947yUM2nAYzZNGJ7GAfcVM4zhyviwSXg7A4jZUIbM
ojGcG/Qp0iTw205zQW9bbJcmaEx3zfmEMkNxhappzo2/sEScnhCAP2v9/WqQ9mJU
8dTbaeXRE0LdyaNAJpnZm2leL620F3hwraSNs6htanDDITX1jwvJwulJpjC/HiW2
6wWhuyEz+hedRblfLCrXCak4TMJrz+SIY0OSdzSzAdHq0LjieEDuFPVf3iUSfxcZ
h5o5+S+VvE05TSWpuoKmLXyxWtfw0nlQCEEZR1MnVrHLGkJQUUQ0c6LTy2QROA26
RnCurdtkCFU0ChkPz9bqZMTagpRxTatHLDoLNr0YkupCs0fB9kO8dkAoSvJwc3Om
4uIrMQFc01NDK1a95etj3kIC6fg6v+7TMMWZHsJ9zZKIm5q09SESuwVnlryO1Mk4
CH5ZoZ50LLDIsLHLK2TwdzXrKWugo9Wznni5mAZWA5YYGrKEQcwkn5pRAGN5qsW6
T3xzT9qUNg18YNWOeSJpqky1zAt1b1fu0sFW6qhwis2eRC8S574OHW48hENS6q62
oLZQ9BZ4WevtfSBCS7MLpy82U0G5RmWsi9wAOG4eo+/uvgb8SRo4srqU2EVyp53o
4w8vvWljQr47bWAoDIe5MwghtfuzWGvdFSxkqFz4HhYGh3wZFPpGrxkyMvFuNk2E
wOp8E6Z3s23+JfG4Nf/JmHtqVNffVh+lcBW74JfukK1SjM7HFP/etjPFO9K4i920
9qftfK4l6XJuMNw7qb4vywl494M5NIDG9s+hx1hV/xhk0nKMo7VbOuJuFLaKCuCf
ukbwUDFYj0VzXHqXbZmFlJ7kGtLfHBRTK2/FalOla1ie5ZW84AqDgXWg4HYhAdiG
uJ3TJ5WHFyjf+xsxnQnP+RNNaEaGnSkm7+1JzudVIPwsqlASz98/quhNFLSgpKEZ
nMWTuffe1OME+6Dyj5JSmpD7vHxBd8QWrVRmAXoBdkwvzxocFc+xR4qP7uFbiw4R
tF522YLJQ4Y5TS/OSsscy9xUyt7dgW+QH8xmXqs/3j3xRFVpKtfOsctEVuN7zs9I
AeQ764ig2SCbtGLLMEKJJBXblqTWYmvvHaWugWo2Tg8z566m11OQ0Dm/LLbTTNS2
m/PteokKvSGeI7OUDhUMWWihDJAaipQqQTolXRU1SiS2whOptAQxAZs/c5NTlvVs
Qn2csCrDcRLBYeeL4EB8lzSBvollFD8F6+k8GBpt2S3oKj0/fhn1VGUzw8+ylpDE
3B7jccV24zI6PFYoZyAXhfjfakM1t1V3JxHIf0JzABwoXoJX+EIqmYnLhLgF/u71
Udfw6Jy/msDOypK0Edpe9wBtIaEHNA8+ae/Vwqk8MdO/rJkEYoW/ydTYGE3PSsfv
/aUDWhHudquFGvKyIKDH/gsljA0JBq7KYx1lEYBcyc5hQr6yST7sM7X/775QdmmP
RYBXlUCuySXkDpnZ2zHeTFLDfKhL4EQiuKq3Mx0EvU3A+5m3AcVXAxJ66OcELycx
FfxTr5nifYFSi2LxSbF0pwl7ZkVxf3MRWV36qiZPgmZrhkYGQjhEEgCz+zt6AkZy
tvJc/0c7nxBHQs83zCoTG1tZXpR9CFRNSdAY31sIQEyCRknNFrJnG/C5ZQPqc6wE
LVK++u5Xf9QAyn/ZpC/WAqCmOaXghs8ehnfjHXafhQ2XpSyN+Sz6Mrr1IpHpbg1O
95ycmv55moZbWTqfSCDVH99PxHELg3hO1wlBgYhtnJVfevLUO5Rufl4momh7qgdp
UMAMouwLFGqWwD/8ljd9efJu7qnJblnC/TXj4dbch87Aj0J7TCDDW5hFT4MjmaC8
AbzL3taAmUcrPkDuf9I8E2QP4teA7PulW+Olpho3P+l80CJ8ZGiBydf711ijQAB4
S6bbBiGzeP0QtM1Nxo7h3BUTLDSQRBG/qXRzkZFcaMqVzXD2ZKT6Ljed1geinqzM
TdJPU3ksT4JM9lmxp48Gt820vihCj93usUTekLlnzfaiZ6ssX1iMMvzxtw/jxH3N
9No8q9e1wvgeW03y8qXOK/p+EGoV5EkevytsIyeN6ut/FkuC35blhP/cKVh5Z9vr
got1jmt+fszOIwXwJJCaLl5WuZOFasGeshV4548KNejC3LkplJXEapYK3XdXhbg5
xb80Ils+BErWmOoDjoEG9UaH1+o0ll/4g6QjqHRl6yM5COAVtysVIwKD6vjGNpvA
SQFQU83ly86Wh6AOvtZxbzpf+Ae13cEQJMJJuV68r80tJLdXWqmiemv94cXE8ftM
zi07JvgFB79qdyBKwjuW2u2iaaZK0gQ7S8sHtDB/YC1SUvfSBByRizBMDYj1fSiD
7Xj8DDx53c2NiVT41xo0bdqRHWntSg92WPaW5HSVqS3bMLiMYl+RnWYTzq1a7eHQ
2bMGDNuuXVsLKNYAY/OeL9yyjJMgWxi9GQ0DQZm6mP5X31Dia0YV/Ooqq+oWSfQf
39JwY32ViSqo17BVT7ZEaYAHmAu7JgrTNl6V0rAn9cwVnN2fl1KeD2vImMAFhDBm
vAvbQ7BQKAjQVu0uSa6ktZlwe2Nw2RSEzmHs2LOqBXjiz+H3VkhRZxioKJ0Geub3
CB0X/WU+aWJ80FCJCg729Z72eUxaPbccxFHZ/ELhXtVc9CJODoZpND8M27KjXCcl
3ibs9QMkmszwv+/GTqdmJqmLjjafqVpzPZfrgsiFRYRZTJsindu8v3ExBeH1JryG
NOcYfL7nXZxtGSnqTOMj69BQZZBwXVXqAizPlbU7qBRzjA0LIIi0D8gFLDA94Rsi
XeRj0oOjJAqrssEsoCjRplqn2Wt18ixUcQiHhtTNqYKhjNwl6mqg8nGzHuD7N6o0
NlqFJyaBBwoNWQ/oHjdoV7o2mwkdRDWn9DqC3/DWlMnRUJEAdFk6XuAdPqVZzjj8
GTrGdu/bulA7i+6MHKBMnQfFtVd3HC7iKnhj1/5O6U2hRri6vlQwbwRYuKhTpHDu
ltUQt+KSo1Xs7c1xaAktpNQnnqX9zeUvUF6qBMBnYb2oeSkZljA+RWx5SVar9UYg
sU9woZ2gDefJZgZ80YZ9qsFEB8isNjCiq6BKgsoiBjTwY3K4ZtB++34xyC/XJ4Xg
hzz2R+qa/VMy4HD1pi0nCFeZJm1R7UbMaMcXw2jYwIqeZSrGU1K4uOXFVrGRfUhM
3js9ZsuN35nYr7sDstImBLagwo3YAAbnreVoVPvvS9EXqD6HtzCI794VeiTBgT59
xnqZni6NuGOFIo1rIHMIO7+LRo4hLnBrm/TkU11ByD+1BG2zcGn8am+JRW/tV7Cx
6wLKp4Qf/OQuKYwlStUT4kWl83sY66nHKHKtN+lJoanPaK1Xj3E7rV2i3U8LpxCu
KPxTe+BDBv6/8HZavv1BMy7YU17Q9Mou0Y2RjvcDzYtUdHQjC2Ry+WB6UgSro0Yg
hU8CAYBiQOqIT1/ys9QDt2/9371iPNQlWvEvxeTLWbeNuqtJ/Jgs+NUqlQc6G8lm
bezAJJTjqksh+4dn9zI68B68HbwK9xSKJbjZZRoenKl4AZ0HCxZ2TDfwbaYiagQ3
H8TKvvl11CnaN+NI/D0LgK6ktqkY8LKE1mDOGlIUvwLak9DB8JwEhmuYEG8We2YJ
sc4W7kT28/88ea5Do8UFdEzx0CGF9TEZ903iRUOiJwEnVWtK0oCgIGbyL53CQEWM
1IfyUkwIz4AnsRAgXggEI3UfZq6PmjIZ3eF7wCwsEPHkQNeTpV2CtsCJW1l3qed0
jlBH6ediieqcYNimt8gA2eWivBPzjQEwQgb6cKoUZHjUt67qI/SMQpMxL1szqVrO
j/pLfe6/H7sZiIgzFkXHLTLp5LdYsZ7BDXMLWkdWe7k7eiPVQPGuOX6ESVkK5Hpk
IW4G/rpaMEGDilSDPc1LBBflt2KqgzsVeTdH/sPdZY6oO1ZTDBJnpZrX/tJqXakI
yd92C0/3W1IaZQ+I+3ZWi7LEZys6OrMEBEjyfTfeGJYUlB56RfTRb7qKGiEFUAZM
PSgxWMmeB+4oXoBIuBhhChjtSWoHPLsMcAkEFgZhwC5Ped81lY1+D7D3U27ZVNc0
o5gn8L3ZthCDSntNJT8QVMKKBGabF+sD4IBbAYlKQV/nQxUjNd4/2K5f2SXFcwf8
UI/NyHgmenL9ZBSsYUexzVHm/u1hZSchT354/QCgsvB4GuCDa3dIyVqv6SOU0eK8
ngh9DsTN75v6PEQbPHB9mhWHA8N/xEgBm3UjRsp6e6CVhQzOmz/4KLz2ZWHvSnln
RM6Q6qCLVzq2iSriVECLlOpYUEndG8jXz+NsGY+P7OCziUElKXVMSdNJinMqJhJh
TAOIEeYp54SbzcIN4SyWA8lEm1k1eIjuwtujgZ1a8xbR+xtsjPoh1ra+Hw6k4iVM
kOvwjlkwJ+TpuvqXVl/bPiLQUO1sc3pVk1mBF0gLTzMoNV5NdBAZJGS5YTo9n2rH
JJxQKSJxsktas1EWdPCE5wgg7FRFzcLIKy43vrpvUXNgh21GD8EZDgHgT6wNjQLw
wEPWnXRg2fM1Pyaf1rV5gkrYzhRSvJOq9JRZ/sjBhVYnucnYl7ljgHaPVKPMaD6v
J01jQlNybIHb/pwE7bpV6SDN0Cc5L+l/fC/eBd20HS1yH+M80gn2bV8cdtbZHJt1
u65CMJmhlnXJ93zDp/A50jn/BX7u/Ly/nbSpCWuMjtBoAYo14pmlH5jUjXXMNLK+
2zWH/sRRMy/iFeef4mEQOtvofW8BLYAr7QC/NjK8LNweClu9GMME8AkkpHZNpbTo
7joT3uMJ8c1/0qygLwaVlZfqf6FxiF6ZFKAnAgknYHTAHqC75z7b0FH2tizHcGEd
cMmnp/vmuxyGQBxrsvtlthVMCdBIefeF7ysbt8SS5jm7Sl16XDI34zwGxOL224iJ
M9fFVuBU7ZJSASsr2q84m19XnTCrclrqPwRyzjyMrvMImN/w2bvuAg9D4Hi3Qy2U
wEadscdOrKlAmc72A4mtPWUsCy9pQvg5qpjo4GKAmYGOMMYyT7zvOa3KcHmt9j1n
lQs4O9qPyEgrU17ZAc8tqi7xthxh+KIuc0CJdBfmscSzd21FR6NhMCzrDi1vPcG5
hJyhtxjsoYjcwuLqtgnvUJJ9D/uijbmTgWYoUXdGM+Dx6jMbAtY+dONQYOCN/xdV
9Ir9LTIVlo1FAeLTrRbbjc4YzHDbbgeXF4oPsky1I31n2WXRI4zJgE4fV3AYg0wE
S1gRBPgM+sd22FLSzVL/quD0WIbDhh8hdgaihT4rvxFQt4yTeqMWgAY+NSrtIlK4
Ycs+SPwhkeJKLxuSIogHXWLmWpDCsuJIoyoVw6jJfEtlwn9DgmRPjc8km6Ok40j3
lAlD1l3obGjZmLozYJomXmiqhczGhXKl5bMA4B4pTW9I4PCEzRT1CGeDINOZlVkp
Yw0TerkRzi2OVVzyf3lzTQjAqbp9UjNelavsYTUVh3MPuGKJodNFh8q5QhCw71De
Ub3i6cGXYISu4VNYAeeP6VBAetgkZdFK+0Sjtoh0TMSKq/CR0F7dlqanNQk6JN+d
Ay3lTnbr80Lwpzf/aFeEpzE8TZOg33pf6ZGkU1o13r2ZNmIDfI6IUmc+qMksl16K
gZglL/EQ8CsxUdWi3pKk3698+1Xo2dSntv2Mf+nX2Ue7igBw4z26EGxxZee8qAyl
20/PbbxMj4vQb0hgI9++NQTWKzhCoYmSNqDa1G+2dqt+VTcchT+q7szTnZ5ElB/z
+4vJPQ5D47Gx8Fqbnce+iuZc4zJ2pb2v96NshRRrHuG30hWrmtD8wqW0XoMde3hb
tbD/rh42UTPiaCxAqENuh3W+VOrOsXH9uT+LcU88+VO6c+INm1VCSxr7vxnrlUpc
9u+bKSEudtWfffN3Hm8NkKSvhyUzC4hYsyw0sjUY3PpdSTTF5l2RJcKZR5B2bvxP
Dh41GbsT8Erd8PA3x6sP7HtEfj2IQUF9JfoZosSudOdw9c6WSxYdgaF1NTWmhFhO
ChMHD8XMZImWS9+eYfFVhJ/YNELrKlyyBxnTqOqjVVteinnnFcrAuIwvSOcNLW5E
7KeUSMUChdAaVedX8M1HsSx389zxEk73vezoEzErqIFNuAIPtHps0V9Pusc/7lv2
a6Mrl40ztMERjRdsM+p2cWtTfNiR4vWbMw+wDVKEUn0f1jbS2QBHCNCnzJ+7saa/
hGgcaDDYw1DyBLEm/kDsu5PRTRjsYPIWj5QfIAKNOoDQJKt+TgbsoZDCvEreAY3j
Vs98CTJbUTwlCtfmk2Vt4nBUIujVIzq0h7dspxr+H+KKvViKQ5RGEMGPAwcuhVvL
cGT1YgAzi+w96/PJf3HHHWDpLH827Pnx+aAa7DHVo/vm1h63lecC2fPoPlZ8ALCw
nb0GohsUa+jUSynJ03Y7BLIYTR+Qz5wpvOsPz/InWiTyN+naQDjjriSOHOvwY34p
ecBly2RozDO/Ctx2Rw7M5zzpwAw5KTq+3lAvGnIrI/QBEP9L2qansLm6zCUHKWhH
/dAn6pTv6yj1cP0jE714lDZ7Bxgfvk8SmYG6parFduGYtFdCUdVN95Hc8UrPbiEb
uSP0Rcyp23Rxk7n3d1g/JA3U8LgY+hA7l8zPm3nwmunZJk6quOr5lRU7iEEW4ApG
hu9k8fhx7YlOuA4bc6XC+J28zyb1Ely4JoGUIDNlj04jaQacxTAoEpRN1lI0caLU
ergioxalELFfvu6XxdAYOxRwU2ArV6phTwoy+J4lxjhLKuq06ArW315nomsnS/cu
ExffzWCqnC+prLGB2EB5gasoUrCNj499usSINBO1Uuxc+IDhYfk9aEz70FJou8pA
XjruRbyaoXlZcSjZkO1ymMwGYZUtYI9B50hvwIcd1xa6YfoLnvABUJtLo27NKc6h
BH423ADzDJXxTMk1+PpRFfpl2RRY5Gn5FK2OLn4tJmmXpvZ0hCEU1axA5zyA7aYJ
cY9CJ2363Us5gb9iMahg6ZuPMoMmtgW0o3kzC9nLrwkzNFOyI0cTkcu3ufbM5R7M
F4D2iyb8vpzA4LnFg0WNIbbSVdo9wclD1qwzm1OjhYTD3TkavEDx4OM8ePSJudAo
md2KZODbzLkBtqzHfi9vN48rXJiqypNJQLnBu9GNBogxO9M4b2N2y1yXUEa0w7ZW
WSKTlujeVfkqp2I5Et0TkyeDrHjH5muM625qtCruwx7H4OOLh6Zta41bfbmYKYAT
lzBrJAMPlZPfObJSqnbnM7+KV44aqdn8mfX4eLtyJ+FnxYaZnOKS2gkEQVVKpZZu
BBQrIJdCydrsnzXZalfBP9kZkjw0p96bV+zBp+MPAn3Yte322tqUejkoguVJ3jE1
GLAzk6LmbW6u6EHtP1SynLd1zlD2/NzuAI2l5WZ9WrBnvUZqxCMNzwGobRyytiL0
c3ifNXLvXR1cRkjxNy3wS7A9boVA2fQIv14o2pgxZqR6Go3WjGiVKxWItckCvKA4
g6xaGuwS15vwO7jEHHunfcO4fGRYOJBKuJTq6Z/IJbwsKzzGc9AFOHh+ye43K/CO
eaNPoPfPTWhHz8iiCu8eVtzWy52wYfdcbQXsg5uDl6jw1F+AlLyB4gkLFxKZewXN
HNkye+3D5jGX4CIja+mfIUxhxSmM1hhKNc3pAOiJcHganuQeQZ+CTJp76qcffr4o
nq2KQ+71dxG/OwskLmyB58ORGadpDDNa2hbDWnlSKlZ3RgTUH4kcxQpMgVbtHCDY
gpIUP8DAOfHiE8kia9l4qigXoEvYrjjk85SrOzASdf0wtkRr8+AwFSLwRCerSIGv
YipD5hTQE1z3bMAuG57SOjw6l8/ILSL6qbWGWlVYSjj2CDJAQoa9oygWbLty6YGi
TagZjtQDoPUFgF0w25fdB32HxZfWWd0N9Ne1cpc2UyEaDKVq92ROzhEa64+aMZd4
ZRY3MltclBYVtR+oEOK+gSUSDcrjGiHiTZIIl8U19rEP+HLY2rTxmRpQrhZ0pVO0
hcDCHxteMKkunK2XCKGbEiLVA+UcNzn7pIi3b6I+pYEr7U6KBzswXTODBKln2vnP
rXtyDdwMPh71qNGsRasD9DWAyyynUczejvFSvb1YIBmwYxIIJIk32CH1d26hGTrI
38W+qifbXRkCtZqa1AKJLSk091/CeLXAul2yJtqB0Qr5DQmoYSpSHQo9KNNT2RpX
wGR2XiIfR+x3fcCyxi/i/b/hYRqKatsZcOkC67v474k9PKlGJGicMsvM1iRnRenu
T/fyBSe0C+CnzVlkyEPkO3Pt+I8VUazY0hHzv+NfzyamXq+gcrX95VJ1A0i47KBB
e0iYAqsGaVh/JR/QcxX09WY7gmbnyWTHHPwZyuczC6lC8DlF/3y6oshSgexTePU0
1li7vxRjDTHLZrXR79/F3l+KXAATuER4tn/KGzFtUrxQOyo1JgWvNVcJ3hBOHsrx
7GDJufIITBVPzWjE0pa3w+YfArkcgYzRua1+9sVN/kYeCS7D5JkILob9R7vsvSuN
wRZAqPYYNFmPlpLfb4hto3TQupLUZclRsxs0cv+tCJ3QS0K68dP1CyTi7GaJGgpr
UoJ4E96s1Ch/Vqwc6ID+JOYe4zJDCafLic6NtzvYIaqvrgIVGDPnbPJ5iHQFTchr
Z1UbteTplBh0Q0eck/uFpUNntWa0ebbYXqSk0uE8pNqGr/EiZb6re4m7aEY9QkWD
2rlyfP3fLGUXdCCLFqet6UKdxctn573pYkjk2dN/86uKwIdHO/Bp11mrUBZKfPom
nnx2yl6jxfz607J28hSgVqfLPfQWsxnh47RUcd4lLTDEO3ovj2gwtgPFUzPEmgUE
euCIG+NgiUMN0Js0Vg6DCJdSuoDD7d+tVjG+tPx7Opr1zUiFCsffxCgX7k4sJY0X
MjOnkBztUvVYJSqMlgBz/BPn9w1Mnp/r1opzedeakRoq0nnKe7N1HEQ/Txm9tZ8/
gef3PHs3bP7LayPciDiuXR9FPw3Nqte9O+tsT8xQwf7gjG18rfYmakvQppzoTHeE
bnzKivZ4WAXL9xDVWGyX5SvGjPNANDSltMx52IvVbpnUXC1N3jw9k5ku7YQgBYV8
hwdAdvFJympSLepjroQcqiMT37AA4OE/2m9qTlKSkvq2qrV+NwoWULG3sI8WuQIu
+jb/OZa4OO5sXAq8+0i6d5ckV000XG6ImmkR/aTANWANRsqevsAQa9BN0kol3Wro
ilR0216ORqs1FQFQSbXVLOc96jDPqY7k0CcP/iGexEdNYOLsnX14dBkJAE9igWve
azVd4xU/RX0Vl2iKgju0lfhaGBCsZA5ZQv8o+NLBPieMiQ2UWQCNJ2kupyYRdfrm
c8KmOJsYJJ2NXT3EmWTsZG3ZjGQ5c+59Ihdqr5o4qtbnx42V3Pp/sVKW+u/mAUWF
jNnfLCNdNEKoJKIDYyvy9NoZVWNYrrM9U9dyok/zPgg+iSyT6kEoPZjx2Ee1WTjL
DsvhQ5brpQa2dphLL53EOVmB+uul/LrMAC/dHFNGOK6klKvs1tp2mbBYuY7SEPZw
bNtfLiAUVAbXYMfK4wNYZ+xZkNoeB9XZV4wpXYf/hRjAOOqcFFH3yiivwms00QTv
mziY16EoG1X8DPB1QpPb2bhOkF28Gw28h+xiuGZSYGfXROAVlLczJ3P4rQ79MgB5
hkBgaTPdlAFaJyjFBap74j83DNjjOa6urlkuA/8UqG3sSDLORyM5PPnBDLsbzyfk
Ele025dW8zBqwl1FDNUy+VzcunVRKFUC62/AoAN5Nfucpktnn8ETpTiZwcn0Gr5G
YnsrUBsb2LxQ8kKAXDMiFWkrAM6oMJe19ryY6FQaXwVkrcWXDaVYt+pVeCICbuG3
CJwwEmU4TrcW0zEhYr6jFybmwkPrjuie4aFrQ/yk8E9WiNKu/RzbiAlWtjfVfI4e
f2DhjGb0mtLeQkYW7OMOV6iATO65phzpt5xibMuVB7K7dDH63+NyY9s7RLfOD6lv
Sk6S778JpzoW12N7f88vgw8IVuoNqNQ3qw4pYVVwjMjS9/fssSktX3feiIa/2jJQ
5VdXxj4FdgVd8traqOr87c6qbMlZ1In0euysxYbIWoiFzalmXTm0PnBFugZFBXDr
lKmTFyq+LcgVF+8+BoVdggYlTZKRQ0p6WHlE2KaEC35yC0sIENa194zEpBGDtpIm
8xbNDtfXaslLv7DG6BqshtoqROFjwxb7EYou9RSxxbm8tAa+3KLft8C9AR2Z2kDv
FFZTkMxvv7Y5zlrfdyRi+RQ66sbjH+7PnBa/sxkFpNIA+OyjkKBveiZLWdrGs3Ku
3ipM6AjTSKtVa44MUrGldx6iLS6/wX/dPabKU5uYmVbOUzTWw2NPWKdnn+JaCWVh
H4lFtEWo/tJNl7Rj0dEtsr2INlLLqepRn8Gxo/ybDUoPCXmyVWx43OLW1l2QDij4
k2ICxeZKRxB+mueqZv0T+/fniLTcOAE+ODWQZxaP7xUpONUIK7k6Wn15Kxoihrxv
GKzMJhYWvJCZJLvq6QI3KVVlcNIcmgwW1iuKhcvihftnrW19El9b2AtbloqNctox
82C116pVeTWFO13gcGkIWMcLNsvUII6Q5zYdKKpQu+RRixBa1m+W3ttc3EdyBtNM
Zo+YPxs8H4IoU3P9/knU1O8M6gQi7uglnwbFs/Tfea5MJvgfpSA3JOYNUWSIkDNZ
KpgrcMP88+OJ4wLmNX36hO4AEfSztJiFH+qs4e2oiThJcpPaz0bt3rqwq8PKvJxy
lVsFxnMmgyk/zB3G8X/M7zWqwwKySnc89dTbzCDIVFE4s53dt+KwZFpdmuNXrBZF
TB7jZto4+d+pQV2t4BX9875IBHi5bB7I3/kn8xA5Ed4IAlbcQtd2o6DPW9eYRaak
AmoaATZsEgZx3hTjpEvdV3QYC3LkGPJnke3lRbDtN1DEXBIfVbsaUrCeMJOIUeec
Wmu14OZwThhb0sqfqL0SsWOhSbTefbA9bhPkBxR5xV3HwUoCQY2oQWj2gG1obrXs
xbcwPXe5vuCaFozPnirLMyNHAlzip/Wha5172gDwJAkgmXM6R6Gbc2gLC26H+8lu
Rtv7YefCBgcA0MwgCfBDoh15JBCTFddpL0+hrPwDdWJagj9i9ZEkGglwNtIopOT8
qqS4pitnFldk3BxIIZrEL0HaHddSZFV5Jmoj5PMWmnDmgGL8TF4Fb2bi4m8Y+8vR
BvXXkBslJ1HU2RdzkgZkxEE3iIuKRVVk6jm0w23ZyQn4l0IKadX63lxmwtavvD5s
lXzTL4pM7mk4mI3WvOjXayEEzsHIy80UXc2TSEKfPZxjIjdtCvl+n9kSs+b3DAav
NmEJizfQXF+9QG5NRcU3eO5sMoeSuNGHXLSmqoGoEZe+Z8OyoWiRr4S1T9/Im/hT
nG1csR0DXN9QxP1n0MvwJA==
`protect END_PROTECTED
