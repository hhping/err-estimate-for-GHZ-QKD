`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wJEE3u5KdJZ5QbnwY7O24LqUhqKVgcTiQsXHp9duO+xJ9ErlMbkFJCk6yHEWgmz0
ASQKUjnuiK3w258JVE4eCgfVY88N8cdC3jJpfoDFPczg5vsChXkybQRApToCNoSV
W4IOrrdBnVKsDQ75Ou5He17PBSVFTUnEgNAlz7yMQPw7GQKDzffULz931JB4NPbw
XISbfNuCTcnxeD5j+M/bMXFzNDCGYkBI/OGILkuE0f/ralqmogkOmX/UNlAn57u8
ws+ddZEj6ESvItzhtS05OMgyqY96Fapo2cDAjuuINTQCVnEA0ywPxDdte7A0Gymo
iLM9KhWmAss96XgsqKkG0jt8QxHskU/9YhYwD8mHQLPFISHnTA3YIy5BHkIxa6eY
gVt5fNwDFBO+M4skMSwbzb/Wn3c318bUvn7xII/JbZM+4bdSd5w8XkRqKNyvXedJ
f1/+/tLyemNXjU8lJAJOM/xG1fQMo8gPyxm/bowjH7YvCMpTQi3xbQ11psmavyKQ
`protect END_PROTECTED
