`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eQXMwgVSZxMmMy5lOOEEIhuwmucl982mI+mnfituI6PJSKwuBTqN7kEMmI8WTfKx
+hx9ZPkCRiD2VFXqy86LVdHMPbiaYjXa19qG0DzfDMrT3Gk8bKR3GDHjAxwWdWj3
rm0wVDUjTeR/pMDqaP5/QDfRAHS/64MJsESV18rA2mV9y89JqpVBT8W5TrRUyNtz
OcYpXKfXaxxSVBPv0YMR0KIUiYvPWgLG4slixbms6xVgl6snoTT7yA3W2Isawtnc
tGNnJ9qLYyA6NHYFXJvnQa1B9MfmXlAOL0plv9nEPU3VAFLzmfWBVwjB8wJfPEK+
oZRQsb8AGtclf07jam/EkNxw0UnBAm139wlD4Qynr3GaD/dbw1ucOGSV6ODyyhWU
Y94Xpu7A8lfv0Nh0D21h4xtCizIhBzhLeiwzTB+Gg43sBd5RIhSUOGe/jB7aNwNe
9VWdyB0HMAXxSyDzN9rh1EGsp6k+nvimJOxdUfyBQS+O6GE7TZxRn5pb0buIvcS5
b0arTJ0FWIfH3dlcmlTfHeo0IctskVqxjXi1It3PNtPeQg/K+VB5/OAFICEaLnRq
ldOFmleu6MkGN5uyf8O4eqriYjAfd4gYVGXs9hqLqExiK8cm5QqraM+xvXjUh2Io
YJc4Q60qgxYjRs2gJhX+1fEXZHxakjejKFkZzmB82J5h0s6C1u3pOfQ+8zI+Zli+
OFGEWEogLwc7hGJdlIIKT3eSFHk3zgBqZhEZYVCZ0Qy8dwXw/dzsmRRjL/6V2ULZ
BqM4adr4ruC+htlV6iGxlc/+ik2AwOrczctEMJ7j2BxC08Ueg5KCcDu+7Egfb1Zu
QCOFcKOAeBpPvPKYMuC8ek81EKesYP9eV9FiUw33cHbscV1MVRER+Qt9+JiBgRA/
Xl7wyWW2y65kaidy+MTKlVxKdruTTQy2YdBtW33d/afO6dNMik3efHOwjWUF86na
2pZROYPyUGjtU2wigm9sOBYow+0rZfpyKb8gTy5uTGEQ7SGQIJja06HuFLA75Iy/
NbCGLq47ofW0RNArFDats5d5CThKgOvBeQ1TRniyj2CxRRsFtukKEjSg5Oh25plb
IqWIhU9wIVXs10vZ/Fj59gU3qXlKAdk+DkZcVoQqukVfeESSwjb2u92h21Wn4gv2
OG49UyQzRaj1uRHKYAsbb0EM3QPQAmCXoteXFSoweAm7HkkOmtT2XaBj+ZUSPxQk
bic+9ecBt+SkEEo2Mq902zf4aXHILCqJHWAC2CgxRhSkbbqAs573g/H1fJmLqead
IiYwtpVy2LCGUhprMpXSK041lyePk9L+nULYlCDySfBxt9O12sbvO6t2Z4yWJ0yp
i2wKFNf0FHz+1NtBlYtDlrIQOxjraipJ6Cds5kmGjZxS51tFG7MxU4YTNhISIBq9
dQkviVTtj6bL75NzCTNOQbm8H4Rb7jca718KjNCyZ3NKhSVL9LZ656ghwg7g29L9
4wPDsQkI2+9T5SjH0y6TLEffEkX5n3w2iAx4lxoig2uHcXTMaf9jHBfUHjNqYr9f
F2xK0bmsEkiCWCoVQ18zZtpFMKPsESDU5pMcVFXsMO64zXOd/Pr+IRCvswJb0L6Y
dHXWzfnyZgYRl02vD/BbFzAkZ4wisngGc+qLL7BCv9aOBzNTOL07p76+xhxKZuOL
hWVBIkpFzK+0UXIQX15U1pTlEViUmKM2Pei7oTzMbtenUkVzy5+AdnaaOQHIaCvy
kLysI2eGvFJYM+V70xauBpOLEmw3byr2q9V+OiOCgfFKTg18sZ793whjWmLORm7a
HWqg/s5TwPwnN/5NdHizzpfT/964b2gF2qJmPr+345sB4aOe63GK3fas5+9S4s5J
azu154dLQWGchohSpE4xyd9IxV5F5+DgLQJfpYr1YhagWaZ8UpSb+oSMJrBbz0+H
BV7T2kEx2w09VPucAncK8fg8x9+8SG7eB0LKrFRPs4Bq95c3d8wfXTa2iw3iInTP
G/LTfDVkZLSGRYq7EH3+PctfBls6v2GHcBNVpuIA0U5ftYI+CRceEq16OSAvPXzN
L8sjCOgsDoUncmi1W5P3GQ==
`protect END_PROTECTED
