`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RVmuack8tmacLO1r3JNqgY3MRtGtrfHPNbw7sPzb6pdzNMyC/sOd/OHPnJNSd5a2
X7jKslg8u0tQhR0/kykwppardfj1SHzLMkPeiANhtPcDIX//gwiUV273bfQoX6p3
PEnuQDh+IsFDREKpy3q8ZzP21hzK1kKyekF6SsP4X2pNK316FTmCLRAEvUYeuSYx
UKu8rniJgRaQnTNbYkmAcliJodkTjwUsgOmGqGekyeCorH0tRB2v8MvthuarTN6h
L8ruQTQubyds3TbGMVu3mg1JPgdtOYIiyLxOANskl4cqHjHclplNxz0YRkMh/RQv
EIv+CJ4upufQoc7ZsNl7wXsgZXwPlSh9YSUF7ipSdZlUjw6pZuBHT2TWpt1J+2ni
GL51lcyJgAX8wJeSrKiC7b4vXvcAm5BBk4iE2dd5cXyeVcAXvsGVRW1KfcuSmXgH
ed9XNlYcvAj3iZBYS4twGOHjbUfRYX7EyKHgCI7WoCP2rPbPBBV9mfOenpR93Vk/
8vmBwC/VePiEt1GpseAsTA6S4gDw0uX5S+iaLyi9Gqx8Y4cjvWrjIvgg0LqaA793
4XTAjOIWHj7o/xSGfCCs7zRR5IB9xbtHHwTx1TFQV/UkNMKtOletoPlUiwygg5CI
lGvi8gi/yzVjHfsecqEu6qdWPrCIqPpu4KVFX6XjWVjQZeoq6lmhQprvYDoFMnCL
3QLtqEYAPEXbcu6/Z6bVKIyZn97zOIPd0QQesYztx0qAibdZhQWjWjK1W+ESgyOF
U/1KBe4kN2y8sf0Z3p7oH/UkI7/OBwxCly0e5bPJUmoi/V1VKrmVl8fi/6LkTJHF
jIZ2W4uSg0O+x25uDHbU/fQKJ/AtKgk3L5PJ3fh/QtqHE70aS3xx4Q5VtzV/niYa
9YTfizyrhfBQuPStfb3Uju16MAqGiA5KoqhKZlp8tKyxxZCGxgQAH4GOi+wgmTl8
AzdTGhvRav6dfApJfhWlio28LpjpkZ6YADyJrxLkBsVeB/tYekbdcywvFf4SP3qI
QRV8fVI17yI/eELjwWJNAG524vyDQ8sVTtPFjX3Z4hkMWQXIEG/dU4/IXsQcuzCx
`protect END_PROTECTED
