`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n3ieL7AqIe//wLceAANJleT5O5SuVS3gKYlPmhqSalWzJaSSYK0QamRKT4voZenk
OB9UwJM0brwQwdrhW6tjuySQusnOGYUwK7jR3P4cDDVsjBqw5sbUgNECoBg9TuAe
zUiN+sTKPktpOAK9qqFKgXvoaI5OiYlQC2qqyafr/TOgP+5m/Y4Il0vR8JJnjHo8
HvJ2K7yMvqEzFfrZKaZuV4dntHN5e7km8I4xY5xST5NIN6XDkDOROqJJd4CteMdc
azuveIQOpTGdollLRGPHt4xBqFpbsW5EeFzH0NTtCJb2KKsrANZT0592fvk+regW
dW0/4q4rhOqar0/AsfUOYiD4Cs5ni0RmUZDubNki+u6BzQc3os7HMDUSWjhau5ud
1EWfkttjPEJNF8kVECvD7YUJl0rWRsUYFYNK5Cl//CmrrOAxICLRpG1Q4atuA/Hq
e5N9m0ZV3EniexhsQ8SU9Kh1EYuwgU8DwxXRv4QOzmpoMLkHJIzcBC3QQ//TVhs8
q/Qcg1U8eVYBC2KmYvOzqgjwqAF7/xfMJEIQV/EZARsLyif+MqW8SeO1mDR1IN76
LjH0jwyAIWe2UaMUPw1Sh4FIFP0ZSR0JemwIHBZkrEcyCC1k9bmVXKrFbcZr25nc
8yWsCw+SqCZvj025k/BqYe/yAR+Cp1Z3ZtbcicRTmSK1aVOACv0MRBAir8fw/SbX
JYvpCOQHtLfnGqyoSIa187CvT5euFF/xEQ1vWBYx4RV1Bze5bsI+MTEVk8zGpps+
MYwWnrSiWlGttBcN8Ga0NUvWiEB0PL/q22i66E1PgfoiEvhf8qnxJ/MQr2f70WQo
fHWHKUQ6xgkAnfqxzIGrZpUwmTMak9/bpQUMpvVAah95B/4B/mm28QWmnnujyNGK
Fp/ElcIkld0vR5bK5mGRqMswA5vxlGltHQ8GWHoki66fk8hREeEkiyEpq0lrVUCS
K3Wl2CKkhTQlRdi2znZuAHAwBTXGaaQU8POaWz99y7BUF3hyeuMzRSR8wv3SCogc
mZxnOLuWHGP0TpM5iogpaWPhW+xNLjdTjXnSXBvwYULASBGyqXh3WMnIyiB33rZb
oZHCFxxzoJkmGM45iX0GMZ8C2eyGFZV82vffkbI++aVIDFT8pEpjt34CgSLZlcTk
tAwD3gA1g6QEW3kUUSyuOPUaHEsEIhoByBS9PCoGpUKXRV1HRNwA6IZInp0YjCFv
AUP6WomVV79maEIGM8Z8/mY2OnNN/KQ9liwuFpoosu3cwKdyhjtbp7IQcjWj35Sn
iPFfb+NQhoE22exxvgR7BA/nZsph/bWhfcYObWrH52EqCxle4IQuzOsUCM15whKL
I4q0gOurlXRXMgWb9LrQPSuMtRIJlmhVeQCR2YrsXf5DxDfXF4iK+f6CimFlxa79
Vw7k21CylEkuQn2Jp1XKtTuWYTPgOuWhLk0melfmtmAZhyJNF5iJLwqPtGZDDDjr
P01rVlNbc8TstK2vzDQ+VMu4gycjReGxzmhEox7iekDKWx6jn7Oz3K7XFJ7Wjz1h
B8E+VtEnTiJ7YyGApMd5hnoaJI4QddSymB2nXg4WjzphGxvHF3dTyIS0c8EE3A5P
M35IOAyDETakBaq3b9CLJmWw9qBEyTZOEQ5dKT73nrjCRpDvNT+562gKSa2YUNsa
A5TPwOPoWYb9YHAH1ss/pkdUyYBMF5rXwANQ+SE8h9YQ9ElJ/LbnfM+Rq3AkDuX4
Spw+U4oZ9AJLz6P29eKaL3KOA7yR6xR87mVLedLqbpSo1rmSReo6/8/iYCr1xIQQ
CTmeeMgxO4V5NsiksT8lhwmnGCw5gCBlJM4P7ukcNL5CRCjko8a20MWhhBf8UWmc
7YUbAvOGo+C1iT+zlDlWj4VHRbBNMJVric9R8L+lbt4xk4oYs55J2Zp5iTZLROQr
cvoB5+1YT1WvgOihbBRlMe+YXONOwSw4D1Ylw2UvtqoQufq0FZcIzbO+7HY/lCJa
FGTHHEtH4FcGVX8evYUeNl/zbktekwzgVNOFlovZz5m8x+XqI5PNc6jcdWUgeQed
JSnsuI78ccxSjRC+UBqTjFDpp/vDzis+exPb3qGjuMc+45bp7CcVZqwIOhBa3Cht
egLZKAqckVA6j3V3e/xHBiuzaZD8Im/OGeJG/MZG3YJuq/NeGf4aaHwgLfxUq8Aw
AdsidPZWbQIlXTd1teR6jbx29G6wKWJix4AV3Wm3M3kcvX2b9JrTlOq91DwrfYe4
/3NGKi7pgeDvuO3rl2dz+YHXK9FwDAci8Xv3zfW6RR0FKvd3ONkW9AZ+DQSJID7q
Ymk7zkNsT6IH3oAqt/fURTxswMlAHUv7OmrE/+AIxTSTjdIQ9ZGewzHa0+pP/7p1
0Gl+SjOQZ/HsqJKGLch0AsFcGiD+O/wozDbZU2wRFrIKNODkYjfTyT+2vVEX+RGi
72RGH/NtFHV1yLv5HcZw7PT2qIvDktg7pRT2j+Y7S7x3kbB/UhD/I/oE8SM2hzOS
fAuX+Wg6xVa4ybN2imhsM+jhXE8FTpnrPGb9C/jJxVRHhBqbWJEuenhV6CM4fZ2z
zaBrA5/NpvtfnGJFoUDNssYmbkHbgA29VJ6Wi/lXUcW2H/wjV9ieHDZzGV/Gasjj
bBWf5V/tHJO7MRXGFQRqOHGTwns58s5zHgHabJvDLwFqAq22x+ksFYYZ2vm+T+fz
kXDngD6VajwnQlEgK6Lec2C+XZ5C92ZHIC3GTy+CuT9sWE0sNL6fLer4O9Q3Mflb
i2MsQbdIGTMHFdFkw6ZE6FZr7d/KEOJdkNTU48BIH3DtnY/0M0Mejo7Ol2tg3bXj
IJE8sSTl170a2EBWa3gOIOcxcJcC4WNQD5Haroyguv2WAYqWAkmntnU7+8B+7l3i
qY1lQpaRNyWOrF8frFpvSFJeeXA9Ts5wnAHqmhUVy+om/9M/2fmYvGzdZxo5q3Aj
D0e1FNUFbmT3o/9AEVTGfmNMDwJu+svc/CMy9cL6wJ9rHMjmvZ0SBy4qXKcc6jr1
JfPDKg4vswRVZ8w2GuTDXnc24KwOpbeJPKBDVFVFpAkvx3XQqSmfc84ePZ5yWfMJ
1nwijMC86m/yxNC8xq4pFVbZM0F1xT7MI+DY97l+E/qSA4+Z5IbDgPlFLpmc4PTn
Mtj0QyBqVBq/9MxHB7kvqN372HfeM2WUoQ/zZiEMjILvyoJ2YnNjB5MlxlC3r1LZ
MwZJE0nczxK90L3ivGXUItdWe0QFfqFD4tAS0svLsa7Ru7Kdn+LEKisZ5sOJ/kuQ
d2a/WkJ8kToqnX7gi3qmewnEAODa8cBnDLK5X6CvomXYtBRAmzLlmeh6Vg1Y6smW
oEhYDu4xMSouTakMlAFeyE2scbrmypSymBMFOxCJ/qTNRGF0ylUhTdqlmI9nJJ3D
ijGd+GfTzOc9RPBS+HH3avVDC1d2TsVjV8EoWfcQOUF+9FlTn+e9ER6jsNGciwgr
lgbJFWS8tvEpyPAn4t8oIE/lYzJT71HctOKXvbgXSXafeI78af0DFQj9x6Cjd7xM
iFSb8C/ha/FwFfV2hcBqumnD9eTcw+zJDG7/NxTjZErA6DI+r96BrAWPAD00Q3iQ
896VV2n1nH4woc3VnKkD4nT1KhvRcKiyvYKpa/JlLnEOtiKyyY6FsYs6NWhW1BYX
siXaQ6TBajMAsRCbZhOmvQ/IAGGihxkBcINNIn7Ul0wwHps327xE1yYqY1c7H9DP
jPfy0wqGi5WMX8RGt3QPlQjHm8WGYytjtcP8WbdBAKYBLK98NuLMdAgkdug28h4R
ZyczQbgADKKoNCCSQjMHi4wIWM0vM6KuuzNPBmVY5G8tNnuHB9NtumRUeDTk8991
jD+G4rGPh7QDpTNi3iVYtSJf8RpAvImMJ5pcf1FKSKMd6pe7hDaru6DvCWjtb0U5
kPFf47TeUYAUsifVZZztSDdssv86PdN7j72kW6suQ7sHvIszZpzE8jwC21qlJHDO
Rpp93BlSNPrAddDYJD/0FX0TiAMkXNEa4kVUjjh6WfbNwfGy+BU4vQ5npoD5gIEb
ikMhIQvKmrlq5sNoXTwyFApLAIs6j/+bzxUituPDh3jV4XZcNkMeBUv8HMs8dcoX
jlIkZr8y6biNvTjW6+TadAa3RwGOYlKm3Epa504sSGxHLxCHL5oGliwn7vzbDVFR
Umm6l8CYxxbXb8rUArc/cHrKwtUO0/AHuZFm/rkDojlmhsMwDPET/E/2l4jIg5lz
PKBPb5CKF3mcUgzCJxV1hd7ZZsrLM7hR/Pb/Lzsz0m+0H/IunS5lgvLDpcud77/8
63V3Xa8y4KXDEmpfFA9lthyfQ1TmBFZ5g9KJUUHIQIXsk4yMaSVAzkQcj1p2uRfU
0XwTPSvvZNLzmSejpU2nyKN70NKXFSD0T31Q9jtKuo3ywf/6cMhrpE1a5eBe/Tfb
uX1m1gOHTKZWGSi1I4QyDrdHNkIu7cAKRsyLEjz3xvAI7fL4F5vg2IwD31wal1HO
qVtXDScoxtCQ49jFYJf0p0IHGRt8wpKVcnp9RFcY3HjbiyQ4hyxBK/5ljmm8Yuby
+irkxoUmjOIdbvEl7RGK9LTzCzyvMfuUWRj9VJQxrhv/kjvx3qPS0kfiTfmWuSTM
PQ+r69ZbV5SeKrySpF1phfddm2VyOO4fLXRkHuOLdNaIOmW+IBo6NL8sUAydY1jB
exDKzump05dXRfIMOhwwAC0uCQy8vBZP4CO1fzoG/gcRvu3ykMrWltxKVNz9DYly
I0ZwLTEtqCiiuCLJr2kMaUPLOKlrL6xmnVy1kT5m/CI0N8pqR6r2JvHtdP5FYsuq
uOLhE5xeSYuJySit1VVtmV/5hWUSWmrUtHu5CcXcCVL46r5OJD/pnrULAdaSUGpo
AvIkOYl9CHMIK90IyeIe+JrSMOe4DF+tLImIK+hXFOFDjpcMJT41yan7eQLyivhZ
Eb9WhP9A50y0ZQBl9etGxCdcdJJvHvrR18Kppig8z+0cL85WyCsm//4BOv+uiAg/
g/S3yOwEYAkfHIkqbLVmILZSNyBHJo54lfrl/Y2Kq87ZzYJN80ciLAqUHRkhbqop
o1dT6CX6Mx5/lmsNcfQksDbyRJOTKC2GEQr9RxNf798Lc1UGt/Dkyq43pIaoBL/m
rnikDOBlOr/FzCQ56Zu179oAR4RYeqAHJ8+JgNRUuSc2sdvXoWE7m3j7ytNYYI2X
la6f9I9DSLIVGOqVbqGufD8EMJ1YOWvn1AaXZjAWYbt5QmHva97RlUWkztaX0bF/
zOrFOs8x0f7LzxuglfP0mmn8f4gbiI345zbRXzPbpC0ctCuQlazi/8ECihAgU9XX
1+2jSIVoNzFNf1jvAbTrikfN1eDROFlrEQ03vM+3TFNoqLo4b0hKFTDzra1Oc+db
KhJrUJZ8uqcgt8AnP0l9I88/HBmoL5QLXRMmX74jirzkKHiHvFJLLxTJCZk4llM2
0ajE48a0Upm+B1Gz1m2LcxH6W/CgQf7fYJnlpF4iFnx7eUd9pvnbLELcM723wQN0
fgM8sVYXfutshAx8pzxhm93pQh24xm/NaebYEAfTsbU45WI+LdLOW3apszASnY8U
Em+KCF0p7Vbm9c5w5XHht60EsUJa81MPnhAiiBnDGKaqJadjQdA1qCjaLurrdk/z
q/5YYa83UMA3SRK/G3UhLpt15Z9Is/k7d2TaZq6xUjhprSVLZxRlsRKabcsD/WSE
4lcYEV7ErbN9z6s6GnixuhpAWYPoROI1fpEUKgKwDxqHnkLIWqFzlgJUtkEBm8If
ODh/AOKgbOFRKhtmi/p+VikgHe80/whuafVbMDCQy9YbUXl/Ju8uLLOokVfAaY18
rEDHkVi23GzpEetWwhLwzDM50KcLOGv/psyMJAPYyj7HR5p5dfbO83zpyZ6+l6ZL
fKirt1qvsO14YEkuJpD9oe83b47aVs8ma0OaLaU2YU8/sWSPIdl7BR/scyH7gc4r
zGjC0fg5SLQrjOqyD9Rs5b/tDk9GOVnsBKoyr6FaSR0GWj0Ahp/HK7wxmINiawyC
kaYbkBIMOTOthppGkC5owfjHRyR0ZsPnLLHY7kD6cqotIxyoZJX9o2n0ZMAl9U3d
rArYpxZ9At8vmrKIAzXroJgWxR8owAE4URAiGiqzKT9Hyt4LbSFQdTuuSwuxW1e4
C3OvvPLEEkw/9DDaejbA/2qIUoDRYnpVYbv6YcN85KAQlbI6t53AL7bbKnJc+Xhb
tDPSI919wn41yvDc2yE4PBozdpPiNApQwPt3eyF7rNhV0tuM4/0wQ3zNjaLj7pmB
eMs1yKxjmwbetf6qiibrQ+s+1GcFnukuLw4uXueGOLoeu7foE5kJ4AC17ZkW78s7
zVGe4JvDZQxApv+wDnWBWBBUUjDvLawj+i5JPWyIhGkU0drv2dfXaSvBBGUB3c1g
07e3Ac6x7Emuee/WDrHfFHJ27LGXZ2Sndggsws6VkVJCU8SSQom+bWzhg1raC+EW
ACf82+/WfLXXuSx3RlVzmhxNO/eUXFiyjxhi5UQI+ajJWvYog9CCBh+gjcJwojJM
JJu0q3V22++I9dA3NrfsmgHBmisz5HEjtKhIyp1H0PgKabW+KeWryDNz+pm6HOhL
/xnXfbgQhiwDJrf+ABoX+rlNC612EykNI3eo3+sv75vrqwg0woIzSHPvakGezWX7
EAQL7T64KuOPPqDmAkgBOA==
`protect END_PROTECTED
