`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kgLuqrLRPLDsSdVRYILMS9BFhONgZdW7uPD+yUqmYdqdyiWdHC4L7FHBwWmVbDiX
t4Lv3ZBeCt0TqPUe5dNaKbGtpnS+2dOpIClu78KRJavYMKfxn8scvWVp+JrwfG7G
Dv/3gTsM6Q/Z5YxxT8voX/UnezS93sxOgCl3TS/SG/nIxYYnGesRjHzTuiCXFzyC
Y7Ct1FgN9X+d4sK3U94Q9Sro0JBuvpWVW/uGmiI9itMzWw0rI50wlfErDBhLmLvJ
9OeXldHb1nyLzIGjRPaSA93e213PBtFgC5AxxSa2XafrFyZoOaT3gIsxpHP9IEsY
yhIEXrwYxgnM+CQWvkuk+8bMnX6daV2M3xG2J3pI7uC6tAcHWiy+UAz2Wq6CUb3d
HWYD3sTGFc33wJ41nk/JaAKC5A+JsPL/kdgE3UPw1sIWHN2mLIuUKMu19Lsq9V2F
SgE5WukMeY0ENhqmDnp4+aeVWz5QLPmxyZWcFL/IhWYTgELNmcfqDF8XLkjrHfc9
z1QPgeaQpRKdkTni+zmwGtKFhDC4VTHThTDl4FlqsSbKCMHt8sXEHGdL5wK4b+PJ
JU3AKcbvLNkpP+KFAhQjWfe1N83+LnCVUEAtKT60yghTzLuPxEPonT7icGSG/HC5
Ce46tMyH/79gXRnz+WWZj91FQOY8JCpS1VI7L5ZRyF/H9SrUeItKUxlkfUSbllY0
QDtQfmm31+UP8AcyQeGYeyYSexfc769j5/ozVdI9tDqSVFvPxJ1NoM0g56gSJ2w7
gStKJ8Vy84zP0ZiBH9iz39Ma6aWgXCmyKePGGSGgMU6Hs1hh1OAOGMLsVAP0labc
Hk/czzzhfe8WBLB/ViGPahIpYG8QMKTm5AHdaBG02lwur30cg7PDAgIo4WQ2qfND
XcaayVHq61c7Z1XdP1zWPMB4/pK1DRPWlROfGufJVGvT0AqF8SZ0JqDlJ7z9hB1b
TKTzzwXdMRbpagKBe9nthsPPiEC15HFMc4atU35VyUswauMB1pl+8Q7+/wto95Yj
h4xeFgV9MMxtWRu1XpYWfA==
`protect END_PROTECTED
