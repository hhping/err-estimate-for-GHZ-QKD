`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rdRska+p6ll+qI8clTTsYkeCjvHTpjQapalqAxxqbJPM+3w7EP3YSTQe3HylQSul
aYYbgu9C0fS6vp+H3SLxR1+ZtNWUm2e5DhB+4qwfM2W4gDKmSRfKqY8SWi80leq0
YoX5fi/DLRqFjHOkKUlpTuJXcOwUyKYxmmdlv0WhMrkxJn61DsOAQyCVS7Y1I5zT
ekcxMePHOW6bEoVVdmMndAg0s1cXQ2zZQSPNALDeVOGFWnzA4AkbLo5Ykkp7mwjM
eNbyAX6MBHdCzLEp67dT6mg0PHNdFrZqH+dhejSMZwGwwj/HFXtIiCNOI1+w1Gn9
s54qIYHrls/YM/limxwzxWoDLlweVOsO2qlX86LwWCqGJY3zEkL3jUrhmAQKnseX
mGPBMtCNZjLIx3XKr8+NWpTHPusEcZzR4Z0b/G9J+z7qnAfF3ch+iNSIXwrAAlF9
ER/dCx6ocjy66IriSy/UTOrfRUJdi2FgaPQupsXi5CHnO7vD1YlMCrRBqyJXDDBe
Ji/ObOGX0Rw7IGyY+ylot1SKgi7z8y/7U6pDRnEEgr8wqhG8znlWG8zo3CSG6zQo
VqAytSMCAB4AkkbHDQSElfJSW4IJXC83eYRg48bAhVZ/8TKARoK2IEyD0Ehn8z8M
UScAuUPTiqldAxhvi/NjNpyD+U6/xCHllGfjLV6/PLJMkcGcAgFWP5takKyMfhLK
KonAGrhL1piseHIRouoVTYFfjLo7YtGXVipea/kxYI/2XBesHBsI5hze9FtEa4lC
SselRU8N0NyUVQ7nNuoNMjYSae9HU15V4EpJMNA6OQ6XohZ4pMmRekiuiiqjLA1W
5e91bEzRIUzELsQbsRAFARa/4Tbu42RRcvH1RCgvjcAjLXxZqxNM/Un0RZZE+9+M
1AWTZL6ggTSw71zxKmRjrfjohjMDtF5IwlfwLCG7iaCE0PDv3Il9YAaS8b95n8vp
uLJnWe+SSVIywpjp3HGIFAjF43W8DQs1kBwAFnUVo9Gyxw2rJjwQtP5WIJnU5T93
HveAyNBanoYYQirzpeOZalj53W5kmeulfGC2jPXIasol8GpuJKGLUwCazF9M4R0G
kF7UFcZL+Tm+X10Gdv+wkVqnr/onB1QFP7hbhoFCBB+rSJc0Ueug1ZzH3aVb6IFQ
wZg8UL8qzjmQtcB68E5SVm9lLR1y+gzqLO8yqHBXT6SdtZhnlZ4QK6r4IuIthvVf
RZFC6ZdX/wPdUu6d+IzGlG1pmAixWQA0YNZQgd+1wz3DzDLrvsmrGEcv+4iiG64O
Nl8uXDyiWhNtlnNHmqIhSTlHkjisvINtZS6YaAtQ38dV0zC1GjIl0Q2TW33pNLiR
FfyAw/d0UhlxvbFJ0wPSRRUDk8EKkRG4Rx/OI8BUf9tRp4h1mKSnjkmGskwtBy2V
DLaLnXD44Rx5wWqEUReCmJQdiGcgIytU2MmrviRF7Ho=
`protect END_PROTECTED
