`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b7IsOm29mr1dWzbwVRh8rvUPAtY6ty1MJcDeOvtlov9KQhPNHuwaDNOSJ37e+eWa
m6lu9Jv+pTPbyqAUY1h6glyux04ktuihmzcGK1bpn11w5KhUTdOhthlKxjqTRraq
rsp96cl1/vCuBCILHW8/nHaE67DbK2ZoZLYtyDmInRHpbsAnKmTcsuiP28TcahJw
uT7jysr5uRcCFdTgXPHMxoo0J/8jnCswVu5YGWmHgqOeIXMZRpuYbYmYLAt+yx4+
ZMrx3f4AxN/n4+gyEAI3FhpEfKTidTpQrF+aZ24S3T69VzhT96YB1ldua2qlAwpA
UIfg6lRJh5dHP/PPlGaGe5liQ7zxLBRe82JpyBPsTvQ4imsyXrL91rRrYqlRPE0X
55hISoMorAzvjWYwUxO0cm3yBrcABYSYkNzUr8VrEELpdF+ZLERITLSOoSQCdPmo
9MeZpvJzxMEv5AEcoxAxKZLE1ry2ps4D4ilRNtm9wkTwfJnSTQUiHSNeD1ZcTvSb
fQD8r2GX5oEVEKAvbMF0T8+4jxHlSEm1ghnxLg+OwAxDeqOfc2ynvSaYrTNBblAA
K2eTDJfcOfKdjs+K/E6O8zi8c7Lv2o5qLDAmYL42D5WdT3VxXjOkbvUzccWeBVFy
LJtLdyQfacFx6nMPpwxxpHW+0FX4VmF7nH1YZ339eWw=
`protect END_PROTECTED
