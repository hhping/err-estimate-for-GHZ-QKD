`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n5/t3Or+owbuw6qBcF5Euh/xy7xYrWb4g6Mqfcm3IQxurO1JJFK5h6v2Gkqqo9up
KBkktVsVQjsJ/Jli9xR1MhgB/bIkrQL54vF/MkkaD1wcIOQP39TO2HoojKsty8uN
meHxSVG95Ru3mZx++VKdxFufESHpBgU12ZZWN35miyGMDtq5MmLeYPVEJwYvQEar
AA4MfWMpnYfVaLGTQIXrCSXLmXpUaF56pgJsqFu6bX0hnkmGs6wagmoJ0rY1+VZb
PkF88YX2x994QgIYY+dByRYSEmEipdstk3q6hM3a6e+Ittki2GzNdrUtP7w+HPI6
xE0dq/XwnO0VBxGh1g04hp35T+fq9LtmZGfJUmz1wJ+ydMFzQKyOFuqOjZQL1F9f
czCA4VtOmYF5zVxUEnMJIgWYl7eVDu25SCS5coehd+pWNjRUrhMha8MUcCBirzFC
nKldmkmjCEQgln1tuU3PKd9R8cKxSgHqDaSsbCkDR1njY1o96FMMWW41LxIbUWbA
Db23ObkaY5nlBYXUqSt3ZTIJFmJbaviCNW/80kN08N3PshDannwl3fEyDxNblEcX
wklAjmEs93t+2CRXshEQv4oOkUs3Loi26ssPZWDjrMwlemVo0BxV/SLjUrHTWOBZ
2brWqKnDforII2E+XE4ouCoVNK4me8RIPIMOmB55FpNe4JZgO+An4KjeEW1K0ftc
PNYm72KotfqwI/XQf+x/SdNVnC7kEPg7YvUfo3v1MDwCQifIve4ivJI/xcLcDNIr
5NIOPGTbS/Ns8K+nLdhFe+8WhCxOzW8qcSQMrw65RXN89zCzagaE3JNUQ9feNq1S
iJx4ZuGzjOhY9uSrNjTk4nt/wkzh5WFAxaSYBnSmOq6oytgwRxoATRCt0mSj7/I6
hlugoik0we7W62bXGXBbuz/M50dzxzlJeYP98UygPXBHJeNOMSiqDKWVXA3g099D
j9VGfpD8ArTGLlfFZ8qMnrG64B9FNNcDMA3V9ulem4hHox8QOMVga78SABll1iTy
+DwEzO9XFrWfpyyu4KTgpm1PYSzwCTcgpzwH5+6WDm24ZRsAVMGPPUY2p+6HL8+3
hi3GzDopgBmH9BUYSzo1TXJR5Bzl/hFGilWL6dxQRo+18ZgqGDfGGQKLWPaEmFvG
R4GhImfXaIOQ/N5+I7b2MwcVWKx+yE5lVcym2HSofT8=
`protect END_PROTECTED
