`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b2/NefTpUU/J/flCJcEQSphbM5p+eD7p3PqrOs5Ouz5UKKk9ITWYZjZfodQThPxR
b+gXFN/WhyaYSUyF220L8bkaJHguAjk6SAVlNhGz4uNwEP+AhQyNeVHM2nsU5tF2
YBcB7vemQdw4JhBEdNsdolzjorfZ+ve18DM9PknVIZwRVqEKWIVi7tsN9+Z8MMFA
bbgC2UTQgru5jsIgTIfFxe0gdcis2UGgsL5UWXOzukQ8poqe/cYtAFmyIrK50yzM
5KfsQB3G2dT0i1vCxKxCWYPox3zKtZljqWkUzEEhAoQt8b+6kOOOSZDb/qqkXS8e
xMHmtMT3p2Al+F9K2nz5asbUXb085McCF5ySQNBzP3vC9dvBnm52h5W8wZpslvPA
GvYIdWsbQXnuWkekAFulqZU+YOXDMRGqtkqIIwfp+gHcI9QK45WkcE7lSX7X984u
sZvy8/eE1x4nu6rokufnOVb854LbD2UxWvvOrZRZZgrvDCpndyR/NOGhT5vD5kTv
R+27GxtLPqlRsL2KEJNLFFPC28AomdIM/TvFArTZ2vSbZGTl46EnY6MoyboDsfQT
PlLI6E9AbJhYwVEsMDzA4qzyYe4tvGc3sumxxGxWdT6ZQitx7kWInOadX/SzVv9w
bnrQdfeg2xfscB3j80YNtF/oPKLKNeZnPXp1uQhSZ1b/wFgrYdnASJTuu0qaSbUM
8sH78pNDdlX/aZuvhJp42eUSbjvdtD4Fuhtplo0ViWqKEnBGU5kZtxLe/Igb1yXe
dmxbdr2LvWTQjoO/iiD8JRnwhmXgki/yFs/osdvntdTL5Ndrhb2S+ZAzxW+u3ilo
FP5a5O2Y4rWV56wiUwwMCunKR8h3SNvPae/j324ytG10suoa65KioinlFRDCjTaH
/niGDLMna2zbKKZIS5/qTMo0vrEA3gBenx7PYBKCXxsD3YZJPtdq+ouJueIbZTt4
xzH3wa1ApfMjRjYwqz1PUbJhlQv7ZeZgVPfxX3M8VvhGgslOqzcfpmUYQj0qa285
WyIxlWBdqdvhPjg6Cdf8toLCdWPtZU2DEKWHVjpmcSsXigXwV+MArzlLpL00Txmz
lKyjUn7qfPrAnGH35gfRLrCyPubyOgTRuhR/Bm5h6YV0PKd9rwOm2tJtlyRp9web
Nw6oyLNCy2k8CrAzxlk683r50SDOxan51L2Rczecz8k76ItRVvkWQiaPJlF3gPo2
LESdqCh0eqX6jyHWzZPaaEEFcblhpAb+fk5oXfna0zroguwR1fIcUtGfYerkemPP
R89ft0ot8aWt7QQFNCnXtm2/loDWxfoVrHOWNZC3Elfdx5RVjypjXF4pgzjtlucG
3B0URiHE+yZ8GrytRTFVjBOPpXyPpaU8Gptd61CQ4AcZe/SYsTYENO+FnuAF/EXU
K23AEoCs1ynv1rcxbgwEMz/3VLhFtQ3MAwRXw6duwkUO9zq3uUFTB+GSQu7ephbU
LBYtx3yD+Yclf/AU4abC8pquThlsumPuKgwyhssLvhXuxOfR28TCYB3lQvHYh9FK
6MRecWP+KmclidJie58Cp9HrrAvQ5oZ3xg7Km/3wu7hsYmc5/De1JUt2Aez8aEII
DE92R+X0MeJfkcQ1FtB4BEbGX3W7TVhenVt+lk5njKCczwCfAapoKYQQParS5tb+
+sAGH7+ijWiP8j4bQw47XegMvb4SbVFfrAY1XVQDF0jP/9JJ+Ts+hpmbwmfkJnTV
R4ZiWP9Mpa/3t+eOULwmLp9Y1W+CGuWVHJhfxMY360fEVeTtXBNQxL2r/rd09qTk
o+OnZrKP22cVei2yAm7z4o7GETbV7m5nWlFhD0mnZeza0dvSADT3q0w/vWd/fUvh
d+jaM2jfnfziJrF96WzAI7ZgYHMUiS/GRADIiGm/B1KMm7uEaxV2r2JY9HdkOPyX
iB8YEVdVBxvjxH1S3o0Aa9z7INA4/Ump4A2/UVnO/XRplWnXQqx0P7GUgktM50xj
e/gc8ff5BF00a3q8BnFTb3TmXL69cIqO3lqljHhKaMOrzv9P3t0qN/eNqvNzclnK
xOdeHFyOQeFpwVGV96T8tJ4xTlzMc3yB1OYt6nzwekilpc9rds/2lqR7dSmrOOBL
N6RShD43KnK8egibpxz+1WYr9Bq430Vp+59B++bUpqIYWcacHLnmvCIw4jUZwSzP
I/h0gOxE6WURafy2SlQc6HSo976NrQSU2oWsGHHN1w8D53UUfbkh7jlyLmD1J8FR
Ghs6VUDvOQN5m9+yjoPKcM4zJEy745E2EwB8KZnuiBMCr8GSAfMJ0uu0qyf0JqYj
q8ZR3Kxd0pZVIlUDJsmTYthA08pO2bjOOQKb7nc2fFjGFlo7IQB2LR4jkRrOhDIF
5OJXWwhTr32cyWr1+C3I+8cDrgSxqZY7M1DSvSfHiSeFAYOEB5dZaq9uHUKsKCp+
FuFAZ80HPyApFnWAghK7R32SSnNoAvTVycQcJBGSB4PqiKV/op48wWD1qh6Z+AZ9
zqv0vwQDdcOGuWUeMxx53+18RwvWYV5CvBlOrdPgOs9puvcu5N5XgHoDO9/Nb3BN
SgevJSTJqgOuFy9WGpupW9vFQTANL/6d2f8WIwXTJT4BnmD0LDNRHrmlm6LZ93p6
ox84zUnsFiahtzeXKpoUTRJQC00s/ZQzxXwpmu2g353Ch0mv2Q/70E35SpCMS3AY
fXdI/OmcKyf4T/PmLN+QcOmmFU3jwXQ6EYCXH/1whNWvzLu8E4ssKN4AlX+nq2ZA
HOGleujpKaU5SDFTyjPvENbcKqcoXItWJ1dT0kgkxbp8taZzUB6L3AU8U1TYyOoW
oz3Qn1+WUgelGHQWGoxFTJcqBsoXR/mMwtuRM06tORHF7CYIgjSRwwdv2jM2GZEf
2UZs0/V21FLJudQomTgzzmWpL0QehUGXyaHz+ff45N4PjmsEj+Q38n80i6RFnL+0
KbkgOSWX/ET13El9QPg7nEFnTl4EueD7EkmN8bheOewerbipAn7ErnHVB7TsjFZU
LwCKNXLq/PpzGTSo/XWf/k2K4lu7d8OupodScYoDDnSi2tNHsUm/lBRwYTX3LRgJ
8l0uaPZ6HUsb2vol4zKlqZF2b0MQoapewq4AhMXVFCcYr2Mc5YtT6OThPFCWSImc
vRviE1BXV1XTDHpTccurROr32upD5vVPBvxnEpp1KY6Js/I6JcqNcaAvRlB3O1bX
bFcoQTggpPSbCRSkJFj5m/yD1Gk6hKtADwx11p2XO9K3FhzYZJK090sJAkV+K+b+
cXkrAxfz7wiEZ+veVjpLSdHsDNjszm40zvMzG2UpSGqgqlUuoYgV5TVTdYtwk7wz
SBjssFoLW4hjeKc2DC7vgieY82BzsiN88B7EaVVZzJlRtcIy2YdLjksoBphJPUzF
1A+Eq4sRfDU4OZARyf8N+DiypJKI43Ejmgv6i2dg4cfxWk4x1jJtT+Mty8r0bWp6
N57O17Ox0WgdeIt6w88GcmDCmUMuL2Hu6C5hB8D3Y9kvXdo1n/w/jtWTWJeK6aEF
C+QE5xEamp25mdHk1Ti8v+Yhmct+ljsOmHfXN+is2RhA8rBKj3hcfepJuqK3SDS7
WoNhg+CQMGbQL2hlIw/FEQ==
`protect END_PROTECTED
