`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uM8k63HMIdSV3C+lbZQ9uSMIcU7Y7DvoihzCZCCAMAC2bvpoP01+HDdeyB4V6N0A
i4I2rVhwqZTy7Gwjk7s9yuElh7cZcPJrVom/LCZV3icMefzuVrEzCLC0eKE4hVnB
Zkwg7J31I6iQyxxP9iP9cxv2PN4IvJizp3FDnuRHPuEIq/6hINgqZpgHkBDEGbvu
MSI7m9amFx8gQTG4bGfutP2qpWaHlrjg44gFxns/E2ZvnE8db0RPWJPil33uuq6Q
EZ3zuGnt0+QIeImQRI9xu9dLUdn23dxgvW18tsnkSICb6Kr87pNiOTpW3HttA/x/
zItnSBXgqvl7DdKNUnNWHWMVwbsGWD4gy8XS4ohOeQ0WNRYJHBUGc3OtyfPAHV8k
4ftPD86S/A1e/QLqVwuW+KeNbm/pGDL2O8S4bv91qmcg34ojxtmqg5kqRocVJVnh
+uFTozqOlh5LfusEDx7GDaqIatajbAI69Qgb6huOWYSIRUO+ZfmdgIdotsVDAnmd
dzpkaZod//WQ8J77QgkoOvNxPbiUksfimh+fixdDT0xd3d22hQkF6QL4xA8a0S22
Z0e9+BKx/VyoNxaAs12z5JY9YcteuOWfYoHCnWdTwFq6pI5q/Xz22PndFyCDLXLs
FLopcDTaa48BUw39evJaPkgBP2GKhN/U94nFrdjdK1LPVMDpsjlwL7eLsMq1xuJs
y89GW978/gZE94dweyErrsi6QzZkHBF2hVDMJdOppK8We4bpvP9Eg8gALKb+IiEW
IwCJTNhV1ksFf2iDcU1zMy6kcv1kMeHUUS73YB0cW/Ulw1NSx1AP2DEFbYWaTfkp
fFJNgQczQBFF1BEOX+h3oQxNg4d2qfH6WlIVVO92lNkutPeAwmpFDmA+RXqiHB0t
yseEQD738l+aFmIBv3++iySVaGojh2C32OZuw+TJke4b5H16ht5fFrh8xQgOH4kV
Wj6tBA5Q4e2eckxqknsrdiVd94im+qSFUyX4WzTZcVvjWgZpofvebvVxIvtpH7av
Jzg18sotiDK8+MoCCjTJYcBKzs6/9z647j6JnTlnPUusuXLtrSfQ6Yf4Fw65wM+A
6Ogmu+Za+r8NFTCRnI2z9dPEJZuyOPdHCJP4neoY7dYzw4rKEUayzHdAM6OR8vwC
kO6qcxI5jlNBz5Yt5LwJpGYsSyKu8D3L1yXmSoEH+b6jY+32mvcQ92mK5ZXk/ztF
65VKg8tu/HODCECEVawXSNfBBcZB8vnnXCYEqFaS1k3/l4PQGNcIVHLOmKNDYo8p
E2LUo8soYeOy1d22YMT2ls/L4xqaRXzXij/vx4Pn7Gur6n/ZezUcbc6Nq/T27o40
6CbFG2MAkYx3FNx+yEbZZgP/nMVmhA4XkrsHOSVTDFs9bPutnKhPe+rVmI3m2d6x
+tNTn0K5CmChQ1fBzFs52XMhtvH7wZ/Mbsg/UOPw7/9jUFGhaI5TdM20w3RNQwsJ
pNoQRtK1sbEfjC93fiAFt9Py/C0FhHju9RoTmjAoC4DcA4wpaEAQ9PQn9zBrV30j
omPN98j02lEa4ze+dPOPUz5Ni01ORuSCOMDr83YSmqqj2tgX0RNlTozTleiRQR27
C95P7hTNekY/gnwJkJ1VolanrC43PAKyWB92S8D3Z8fJ7FJdPjKvLeuhTISAixCP
rwS3Dstx9NpmkQYQ1mTFwm3HjIK/O05UvK7CYlOBOJvF3W4GuLlK6d8qvQbUb+dI
/sEUfOetxlFYdSN5/4ZvcuSB0FiW9AF3UfuV+SsGfMGCtNx8YY1oihFcSn2NF0Kt
OMYk6OCiwTq3isy3koZHQqBtls4UTmTH0GEfsiSWPPqdqIo/cRy06HQ5xTvblypF
69aS/EQeR0sTvk5tRhADnmashCnTo5xgcoNu1tl0fapNoIu2o0RFfv0RjLk2TeTx
f2NcRbjKwDfHW/ok5xURTgTy+wWmsT2C6gtI4xGrokBF07DngKVhWCiChYtdj7a0
OoId0oB+XWWa5ikwNlBYiSFOOwd6bR9tMrCTygAN20orr9GogMIE/jj1MrqfW4Av
+1/t1uz/XwqI8TsPwzNSHu4d4jLj6wl+7Ubz8/8ANLFqm96do+FgrXMadmYQa29a
1Pv5008OR0D2XoeK5yfn6CuFSxgGbvwPnFxLvWNnub2FVOG0QoHl8nuLi2etw8FB
Qs1XqU5pmuaPPRtQzd+XUnFw8c2y/PMSEUZMed7MNOjkGXK9P75blDLrR+2EX0xi
XZtwPeJocuRiaB20u8iKBuwaRdNxj+JjYcX6rBuvcOtToLyjwZ8XxQ6Ixv923HSb
ewDSGhE9gznVukfK3Zu3mIWHr/II+aLMiMlYxjwUXatgbRuhLUASPtO6D8ofXuWW
efSNQHoorElKVxP69vON6XWEZTdLohVp8G3+P2WQpVFWoBPxtOyfhkHQmPwBLs8E
KpLf6fj58zyQv8lfTrpbor9Z3+OnL5/kzl8tQAJ3j5YdJ6zNK1gUX/3slJBATe96
lIZP6nW2lkfbjhvZNxTaqFgxTX0hHCHLNb4hhO5rxnwuzt9vZ+bJwOSb/rWIaetG
W6CQFqylkg1aeh0M5brB/+mASIU+a67fZ+6w9QJc7Jxw4XFx0j8KVfgvUZiDuHQg
5nw8zzhwGUW0px1VIyC5e+ZjSqR5hnaFBXYLYvNciSPNjayxMUCt/BS+dpu31Ov/
8GYBWYRYWHtAMiaQXAJB+2RFO0UPCbwGM6sLsoWz7tG1S/XxoanwdE7e9sEoQDaz
XMHWwTqzyq7ICTYUcAgOX6IWq1GfCsq+qWx+HbPX+0SwYjBQHRI+BghhakN0j+C0
ntB2033H2WtgqkbPYgPbeeYhOtzGVWva4IAMszIubNRjaQPTihkLSANSmn8PAChm
bWPzHOyvE0Kq8P6FFxJtyyS2jzIdKp6Fem9YaWcfWJoH7eX4QtdanM7iI5+wkuLl
U2RHg4Cy9yNd4J5ijTLJS0jglopfFRZoO07FzIkv/yxsSqgvt5HfqWeR5SPhL78/
Nyjf8q6ytRm0dBmlGWYmJ62rBY+a+ofRcW/Gxrvl9dpIcmEN9c3iC4Cl/v1er1FA
kAnp14aqcmQdfT44joCHUHDd07B9sv3c5+hHx8HqGLUWmiC7T//ZIibtMs1OVEH2
TJ3tW4ARCQ+jhKwCphHB/nwjoybhw1zeNK9daY2S8v0feWooKWpjDzcKx+cfWQCC
pFLWl+qgC3l89Tqjz3xHf7pO31VAnyZsMmKfGzSa4YoUixO6q7ihqwYwCAhDeF7J
0QTgrL9niAI5t6WMfY1utgu0Fdjys+ChlGdaOdA+QtAE1+z1SJwmOGl4sf2ZzYyS
T+TQP/UIUEg+utCUo9FPsC+zAYUM9YQLCQXI0GFQocyhUF8k1b/FpP8rL8XBZpoP
QivqPzZDjmmge+rHuEYrSIX6RnlmkmGmppo+7LJc82gijmYNzGe2oqmxPMTH3Tbs
Cu+0cKga2qLVBpmtnYnQD+ELY6scGCSJICr6mdZR+ftZUhApgd7wSm95Mwf+m+E2
jv2iL91s9Lcuk5VmE+MiDFz0XLkTmQ0YbNy7ldHEbajaxxXakE0Yzzr24P69lsQ0
4IT4f0wE3ur9GER5YmdFvTc07jxONxp1coWEH0tSSkILAPFswt7w3V7xlRtGCVfO
+DLVxMibdts9239OIw0mAaC/l5R9zUq2s6uLCIXiFyfhqDonxFaF6PFVO7MgmNM/
WPdjsihtbrV1CNScBzbDAuA2KJwg9VyV+Ntv2yThsIFWXU9BheaeWmXrKebhEhkv
jUC6o7J7ujwIfzMAWaVFyv6OZYLOW4ByHgzbM51HJlE7+aquLp2h0/C2keQJvRSo
wlJNsqiQFYw7pb0LP7opH6yEeQeuCalTKgTpOznYOZm42QropriW7t16vxja3tzA
C/T9YROgPifnNdzmm6iUsGjLdZpao4f+PUACySByLg16dknVIOet/ys8yg+vGI1K
aUtKSRCs4JEP1SAo6niLPuzWhtbs9MqAR1Gkh9QasdS016iRIhynruoKOXEO6s0F
y9i1DP0NL2zj1aqBXTUJ8O3zGCx0K+KGh3yxFGNQFNvZygnHLaLE/81BfcGXtPA2
xPP9JB0eM1btTk0w6QiU6f/ICfm9nIpK3yeQg4TYrdYDSFmJxkcCcioIqLGJkPWV
GASCy6axZqV95t4A+RKUs+4Is4GimC+AYbTc88t4TLt4U+VDm26rNxvJBXZrH9Gr
G7G+XuF2aZ/ADrwkfs2ratyur4CSoKIPy2ElYHykqHI6YRjWb0E2q2xJ5Nk8xvdH
gctc4FIIxdQ1aexcuQhvmNkcRJzKUyc/fESpkWoW7n2NHtyqU6LHqc4f4qj8JKcE
G/WbjIG8/bBQvOEBYW+lnk5yxy4jEaNmhmW9QtdSRezQwVz9x64rQrpwf9JpJkSC
t+HFGUNpajX1qI3MY3T/SGb44GXTDDNQwB1EOGdmMwNp3c/eOAHUKpPHZmjJ9Uwp
hWPa/ktGW72TUbMi2O7023xKa3wYUqVBd163FM+RTx2JSMaIEa6KerZa78qmHhKb
F+pBvvJo1sYaZ5NCt9a4F3ozk/r6sf35T/QsiFrjmXEZPMMCIYSTHaF7sQ1zJlR4
99v66dMRQplX5AY/WlJ7+d57CVFeR3OcA0wFz1F3/1sKnXIAmBavJR2pB5qGIqvi
uzxsaZBMJbzuMDJStmpQvxkgG4uZr5TzWOAlDzRkm1XwewH7DO2m+YXUYYFZNg6H
qwWqaDPz5spx2JXhMxqdOQnq84otRDD3Zb0/5Ji8/SeCdsVSVO82+llNkQg/k+fA
sAM489ja2EeMRsq50OBL6Y3KXApLI5gi7azsDP2DFsOeSyIt08MxpyzaAK9dD7MR
PqrwFdYBrR1435LijOvLApW9sXzJEgUWGYRlMdM0saufMFUhDmb67LnHp/yZN1sd
65snpE9ipT7KII3UbdkuC2qSolT1L3mbv3JouC4BnIuDHySJuBwgr+YFg7OssbzM
72aCkFmPY4TuXfZrS0gAIjqTtPJFF+CEd6ddQhZlGFJYkrkjjjJUn3ycVFvdfyrC
CuG/+eadN6P5n5w2sBjOCT424CrlGqzImMRd4QejXKZcfBDHY4cvAW7I0SbkgEOb
KWz5mt/zF1VJ25jRez/cElCKqoyMlbe5eDF4P1DW8UFwNIXN3LjSnnl6007hMx/l
wlaY8Q/HCb63Io4VTMbDfIhTMC8i728RC1RRcPxo0FzdYcNiBe3fvxaXcC96A9zO
qYlu/ZfMwtc6XoCC9x0KCJbABRX2Q98fhDmyUSw54deVCgPG+P/y+5/hVWIDn+Ha
Ij3sLonxeohqh0n2yOPfAdG1TVuiXbWc2iYIWjaOfg16diVSu04ifSHb6hbmDe1o
Bkp9VB+rVvVy4joBsqmkIl3uE0xjyqUGOBEpP5Yk3kWZDkPbOKFW3kv5chnvmPsH
LCBOHMrZRpAcpdynLgDuDqbW3s5VFPrK6gn9R5M7oEI/dqcd5TUsz7eaP9T472Wk
iaYruyGGxt1uLp3RSyXNaJEOYRqk9ltbhzncO0li+MBupOYrLHB8wLuCrejmLBhQ
jthV6XdDpUx20T/nagpz8jCEVxWPxsypcC9rwVetAt/BxbFk6qot8ltmBE3XzxMh
Xe678NGrgqO+0+9o4/+dNl50/+AQrDIpw5gmWu4vz4WeREisa3Neku5NXaWlWYXM
RkbKKw+oLbRcng83pfwFMR+OfIKneJl45S1SL8oMeXbADFnx3VvBemRj3kSxDp2c
K76wKCVhWsfU/CxznVHYrI/1vMwmkBsr56NC5CXgFtQfEIOCDz43VI5+S7OG5Fbg
YhLX0W6SGxAdg7IYlpRdN/2qPeHX8CxueiLdKszL7jp1cecavf57DB74XJGnytcS
fU3Yxw+5DBpw3DpNdtcHOtZUO8tBE8CkT4Daepfp7+CKzTEPW4Z2+F0BQYV9uc0d
pMQcxclIjjxHcwdjVfe/gQunChC8U3w+vqIWBZSx8rC6k3on9t3JjsFqQNW512le
vL88teZpzjsBrSHUhudI4licCyv33YC+qGJhHUQhce8cRUkLJyYbLqrxiFgt/JCI
t6NYDhbfYGQ2HYq/uCDoKS7jPzRvM+0QfNFphoSNyQTAafISLcD9M6Q+SawO6hTS
8MiJx5X85NWmv0vBjnHtzk3Z1y6XbWHLECrYm6LAEEplSm8LY+CrY2Ypql96OrqY
mLdO4l0oyTGg8qbpYwtX6HOKo+ONV+94oQibJZd9coAK8bReM2FqKlzAanl/HJ0C
xJ3jmTh8d82Jh8D9aHcSrT9AzraP3s16YKC4u4bmZieDRHl6ozo5WDRaJJDk1ikb
Lu5CE1jSCjPA5ZO1uki7HLhY5mMn+Cx0wFWA+8nfmtxRuSo0Gcew+9uYSi4piaI/
vBuN9SK7lVeMHjhWq4l/I+joSn4OP0FRIxYRFApvZ3b67hA9xG+fx0lo8JFL4TS9
TF72YSzfBWx7UeyJg82hv7SWlXOdrjUg/LW0y4hUyG/4VgZUpD5lU8+TF4tyBAAp
jkdowypJCK4JSb3jvBFE731j3WpdUB1qLBiaxOfMb5x7X9FMWQX46INIGIJK6Rbt
uEW7yr/iSuAu11kBVZYKCZnQBwysmKOpc89DGga70FKs9LnZVcYQ1cuzzPXWvWNt
QBb/ox9A4NhQsieu2oG1R3wJpbj7dB0qhFSARunnvfHbmkriEbBQL5TnvZRj9kVn
bijfGPjin2vNJpx2uoW7ri5VJe5QTB+tReAJmDxVfAj+DpFb5mbUcPC23eBijwBw
pMoXT4ca2DopJIpwuiDpEdCVUm6P7YjxaCbvYH9naDfREfWRmIdRzcSX6i0+u3ZB
BR/NVlWY4WR5fsclpaBelKpWLvefDEUEL5dmnd8uFm/qnC3qRmWmBLUAS6iL8pWd
ufsYrG5QXFd19nomz8Wv31vMST2amzSW6mkb1CWQxQ3PqXgm7rgGUmWIBVkYXggZ
oyQMMvaJ1rY1lnJgbo7oXtPdwFvVRBHAKD8BkYcu+A/pkB82prroZb1jij+yLIET
GpheNHXtZzEkHj8PzL4VXi27EbCrli7zlref12+VgvRjhkeWutLCQbYV+asR9fo+
8zhORU5JUO4Q5oEWe5unve2tWWAWQNxWq84weiCN1rSsTCidRrVkQH7AeCIYICpF
+RWntjnsRGfHD7AiWox1Zl9j+LaYUpgLopQa6nW8pg4+jUhNDvC8w4uAupuQF2r+
UNAoGUbUAjNE2QNSeDlEWTEN1BCvZy8dU+Z3rhBQX9x2hzVbdKTBOX7bX6LdmSIM
d8vktPbZ1otnQMebfkx5Qg04AYBq6z0eBZZzbTf5JeFvOgxf4Kn4pW/dPEzJnzI3
1l3mTDdt5bQBVT1ftxn9vMQLXxvwjuMLGqrD/IBhhJEfC2pWv8WE1bSsMUNj3xY/
/ekXTnfmbeV4b0AdvPQ8bPvVQ1b+nXfyObZCzavu7Cm0DAdcFugtPZ5S1fH4DxqU
FqB1rda4S8x+pw8P/mlhfHV6boEhkHcUrriQoG1AZZOkMpJBALl2Kxr8M3KYurot
JqGw4AjqSatHQGZ/Yt+/ZnTS1aKaoeXLz+//nTiyrNOGffTL05vqdL+lIWB/g+iI
W5Tpiz9oSHKt8D/SpX9sCFn2irhDTnVvjkVEmbGG7M2qel0K3l9PLlUJNgxc8Y3b
oLWuR+fWgRUNCrOU/kQRpNpD77e1opLpZEV3EzsTuIE9+w/UIu1jyse1G+hfh9Ct
S7okQeE95APLuxTBI1Mi4uIoHPv026CuU1CROxFZSSFldzufSwT0xcdbLnXhKTi0
pLtY87V3Yr8P4J36G+TeJ88qO7KxreSsFtWERMz6uLa0yCe2P0DAPvfhUBfj1yfv
GLXwbhfz1pNShtbq2PnEQx72H+/dTxm1aXWyyq4ZFA1aW/dcfZaAmrBZSCaMElq8
Sv99EOwIzXXW6rVpwsiFIQgLl+ICbVbZMPkpc9ndEmx60Gtwqgbo917uUJVZ7CEi
BR4clfuCb/1bQcNk+ac3PXuHyfrlXPox7iN0+KqLdFG2oWpvuHo1Q12T3U1FDxHA
JnF+d3t157WzqEw+ByhsPNDfzWbJxo/nrXi68068/Saa5XWxlvjMW4NjV8QTN75c
f2t5lFzPcp4EsDukKz+iEB65et9curlLGMgSZsSMjsWg1bJ2B6u0DN+Y3ggSUu9P
tj61uIXNY3nPOBBh9A3/mFcqLBkFH+/YlAGEhdmubkKiq30NruNGub6dDl1oWUFe
GFoiviLscKfEBxFejthCTGF/KU+t9RO368jwAlpsGnSMUUBPsdKEDClasWkwqGIu
zLNuudYrE1Q+hWXtCJL6Yi/74ryU9LRrKWCcogjsEUj9T5RYmOnC12O8TGb/iEUr
I+Rxxlc+PMDQOUv4fucmGwsIWTTYudvpiv4szQ1uFg5qIzN37EWY2eJL16b7WpRd
dzYtHIuxceMdvXbUpWz9n9tPDy94aYCB4YaFykUmo64Lx27lFlk2/rKx/8rUWzTb
rr8Y1HKooShhkhnCzVaEEzSOe/I1D8DykNdk7o4War4v69OrV09bZLOqh1wz4EJK
JwvuaT6E2y3qpxmYQl3ysKigRp9SUoGpDM6/v02TWNJSKQuAhqfk5mG68TVMFN95
6XuquX6B8aNUL742lXrtCdZBab9OjtO7kwKXH9Z/sd/cfIFzBw3t96bzShjfoXIW
syAFlQvZ241jYF3lWsovF6K+HvotOsfE9pU5ljLeQquOtWyqb7akw+8eeUpgliIP
wmkWt7qQtnTtXx2vkuMdAYTbQiD5u2oCTyhJO0NiEJsq51pZ2wE8nc2ABgOQtZSO
YG5NOF0/aOP/VOh7WduZf2Dr8qAGQHHITyEk7P//9UcL/gOyCD+yFdLjpbz2P+uE
Aw287cL6ctn9V4KXwO0ybJUtMFYLLWyxo3FodV4vthrq9G+hpqODDU01RBQ+2Hea
i4JXJe7lcLv6IgPU4tYh4DDavLe/oYaURkSIfThmRuuqNE1EmGQAGsRIW2z8foe2
lK+pzuR7vcEpSt+SqBpy9An5SZ09KocG4jPBX9MWlJUTNNWBe1+kxWwM+q9Fvkvu
6GROjau+TrE0omAuiZjlqQOThUrFfRDzZ95uB7VDjKPvuQB0VM8qymKmgWc3vPa9
g6irmFgiTDYoiXWSkqXXHbDW8C+SPKAr0E1dcQG5Eqwes98B1aE0Nxchz/HjWnd2
6UqOJCnnunBzXW3QumjTibh9iKy2pYQpJzQN8M6iHyE6Hknzv/hrKxv8cQ5jC2Iq
8QweuQ2vLpl12nl3uun/3NqJqVrqTuGK5+Dp96QFvvwuQPnOYXKRs2ITZ6RRRa+E
t9txK8RtLlDmHAPHLcYbZQJgxp+lGMe3ZE4u4z/1ksTNDIWtnJcjqmUFnnBXocBT
/Ow3LZALz0Wxcp1K4yyBQtd4Nv1DxPyfYkaWFWmw7NrZRzpFfQrT5yPHywJ6U+WZ
tCRSPsLXRrkjSX+K2urFrCidrZp6ksZjcjVcyDYvmIW3O+8fLRpEdRBnbfAHTW8+
ORyrrmQenAz29xVldL7J/qtirtEMBf3r1lUUmD7yraZo7CHRyCbnN64toc27yxf/
hvWS4/ew6ywNhPR4YmgUEuckqNd93WGHzpUKdjyaWMXBHPh8SPYYkgCVYU6fSu/G
he9XvqoQm/miGS5IojpKGRyKty05d1knp72BrfMhLNRdSBZXYV9LDMLl7t43rPjY
DDNHupbT1mZWwkudMrt99SZ7Sh63/+5leCQFq94oHAKnRe1WXXrsQ5+qycJ8UBlv
xRZxsdywO03Lw7BQGGMeCD43CLhDQHuARSZon98NB5lFBw3hXkmBkwS2it7WxN7d
c1r0Tm78QJg/Ul7fiJqQx/scdA6fgyU9pdQoAWsp7+udNDa6pIpdnTlt9y3HILhT
93UlLRQsL1wWNclMlKwf8stuc68G6U4xKFd7yAdseplsVnRT3VZoOZaOdEmHtTiP
ZfcKKg5zz2/YJJQmrBifCCMa/j3QqdZjtmR06tos8+XUcxus8PtupTZ06WGPVOia
fFnxg7nTjd0eEE3xci1AhfRJ4YjsCbsFzuyGp9BnUHzhFpbTnpAPdp6IPC/jCnta
7dgZv1Rs8fYkEP6zRXO7Ld8W86fiGlxfCqwjeNGBhOpN8mZL0yKmm+OfvOeTuPmE
6kMzUYxklB5v2hScfSwGTPObOWoLTF4npMwo7rDUb59flzeZpgTad9pJppq7jXnt
KDFpnFazjxLXn3tPGmcHma1U0tMaLuKjJJ/UHddQ27KS+cZ8RLjKy0Eluj7p6iUY
mcDPAWCKgxHfXDDFq3SCt/L+W+P4wqg/PvGEbCuyb1SiE9RISgXLAbJr4BxJ96Yv
zbFVHu7+MP6eU2QYGd7x5IWz8KX9hYzpQK+GS9B0xd1dvjh3h7F7WnbPRmGPPlhd
MBjrVzFAM7JWswIFVMFL8VxYmh1QtYxqXDq1nIZn5Sq+wKz9bg2vG5VcEKyn5GZE
OEDF3ESMxapTh8vMGrzxF5kqsL7lzgHH6u0L+yO9SGvCNFrpQjbS3mx/dIzKLvQr
fQFDYH9FAAUc1sz/KaTgRq2BXnTpi1qqA+cMj+UVsDEPzw6OE0i2Lwee4BHRIA3y
GN/oDvLR13IpHUbQBF7owBFmfMEoNRh8+XSI+BWkzoCeLTmfp7Uj3ESqOH8oKxYK
5JNKyakuqWPQp1UTdqvptXGd/boDJd3xxL6WlNizBrcj0weBvZ3g3vqK6UGk9CBF
SnQZo7fdxXCoDQle9QZVK/8PcvR2UI8csDk45tcTM6lvvn/R4JrKenuwAVmqBh6e
43N5/8aBmRPkYsAip6qq8kygNfYz1Nj7Re114vfvH6G0T4hplgDQGWBfF0grjRIK
gdS0+iP8NANEMCf50WjqoIaHKLJsKMuwlq611MH1RQ3w7dLwVPdA7FC04089IrLu
JpMZ2tQu8CrxH5QkmbHYFjnJwlbOtyEgHAm2WzjWfJX9ELibbR4/TaTU7I4SQeMq
9f00XqAlStDqMOTGroBIxwHyL+iiYlJdkiJ0l0J/WqdEO2DzvCN4RfPsbzpht/4+
Hc5JaHU1eyimXB3zF5XiCF46wo9lIczgknpJO5hGpTjeKVSZz35xdSi/n+I9KGE9
/HSgnRMC3aNYV9iTinpLBTMgbGnRFrFvgRR8knuB1c6ZWCmrNv31hVN2+IrX98hK
AHuE/eMC8I/7LJNiBy29hoGcv+7uytZ09FuHVthZUNwU+h+Wt1/n//01Gk8L53oe
0I+X2Djf7Cl/Ad1GvZYZnmCvwVowUTKgzBd5uRzpNLAfSMvhSE+uyarcdxws4Qzr
ysrt4tXZ0CAi3b0bHYds5Bg9ry9ZAnzZnp39IJNKdRMQoA/UjZP3JGtYrHZTAHFP
OZJBHElXWJboRGplHWzVrDon865X0no3bce4i004EQarAFAV3ojuYF9jVDRTUOyH
ULB5zJDG3u+IlS5mtc3lNRyCn1P9uFAmaNlG4cHnL8e4R/HA/VQHt5UjUU6j71AM
oXu5d/2+i7nvs06Ef8d0Fn7ISDuSez/oSQz1EH2/HR+J9WOyOIvPy7EZH5sMya7F
MNoPXlEcimkIw3hsugwCecqAj/at33TTKG9056hVRUPtHOpLCmlbsGGpHIH4v8Qi
sjU0a6+fWnO/KGwhZJLKG6wJTF1mr1QobutUzMOm6Wdyr9jXUeMArFSPXw62VXS/
9c4O45IkTRkpYJA96JNCzlBTEVP3SuFBNXawYfMm5uoFEDTMuYP25yMfENtt6Un2
K7c/I0NHCmJ4ImmZFuoN+bRK+DoR5K0Z1C3ZVI7ShdqrCLc4apBAWuUk1G7hcnnu
fRHq0Vm4soGpsk29pEQDiLC75qTHFmF1E5mLoX6VVuEZ829uNuehLfOtg51AGT16
6h6nSWnay3NZGH+o6IjFkKqVMyFRCyJvBE1KQGnE2k2dSxMSsYJcBO+EgnxoH5UM
Fvn3TDiE+KHb7Xv7oDeX+iwFYuH0NQj0QAqZcmJ8XNKGFXh4lIGMP0z+zaPaVc3y
yhkyB8XPxEoTEpjS5gG6jKCu+sxPvldcwKtJHlDYsMr4o9yXdLPuSAcCPNNqKSsN
kr+O5rabohIQDLY47qZ9x85+ln5Y9+cKsefqZAyuWzPjd74J3diQF/23/vnaytve
uhHZbQT8kA3HkZ5R0CCf02zrtsHKlnxXx9gq1NFJuf8EI0pvj8p1h1BvmH+gGIaw
Yul37SSRUHeYL4dchfkci6ewiB45I3tcXx2sS8W2tNOlgThtY/L0ROunzz2nYOYN
kaF1KlwHjFFOu2nv6EwfPYzZR/Pc70Mv6NA2qnDUnwScMuFHHo+sXwpjMA5sLDqW
UhdapRjQWgN1sg4jiMSEQOnyKuq3eVrSsUGQjEQHY3EX6bxd2RNezBWuzfYCCBRs
9x+psS5DaqX3BGpgMBoCczwmH7rRlYKi7Lc7UknQQ48UeSJg5GWnSlcNbzlOkx9P
JmOzT/oiz9Gq+oIMns7O2ARhRkuYc3TwsULVJ0oecQA0Xz+oDRVru/bucCJchKbz
SC5Vr1vx4BJBbZpiAJL3X5auGX/JAQIvUCm/W6g6c/RPxIrVsJONAbtKo7t4r7MW
ZGPHyTzkdKDWY85A+4k6jB/jGu7sK5jJfLjSIx7R2r1GUVl/p3B+xnN2Vbmw+LMh
NfQHmzB7VAIzuw+Z9gmuspt09rNLduhoJZIWmXLHtukCPJwCTzCNyjILFs6XOAHC
LUP8X/o4T3O5r9/09mPGhhZ3y+kcts7ea9XFejMhhVjJUbpUUg7lMn2kRTUY5nLk
gBBWlNYThE8OfzSYp/U6c8GzH7m0XJct0cd7AOjUUedkow2xzcPDnbLslTY4xzD1
F99DRen0ZFggNxwfy+f9LV42gVqPzBLGtNf8B74UzWuI8OM7TovH9n7uHrJSLfT1
gkyqvOBh+oqVIAh++TMFCU42TBrK/Rxd2nQ4TVGXjyeLMk0ZxzxkdJbDApf2amXS
vkRJX9w4LKElhgaSTFQ7qM2lMARHcbfKbLssYMYqNuZnWKqjbTo8e3XCEqZFZv4p
68PVGVzPnC6rRI+SvPraOzKEbBNAdXHCs2PyOYmrr18KqGwDnQQ/nV0x9vAuasWd
++fmpErtTrlCsuoXNvlM94vzx83zFyGkGKvMg+TZANqqSchvS7XCy+vgTfSHGRwm
OmSK1HIURu/P6+hyXvb/QtOYd25Gy16GFx8vQV2yq8tAHDKoyFMb89BUuyOgzge6
/RHilzwUrlGVCHKG5RPOGvlq54UdckC0VwwYR4lqH4iAO+chjp17P5tY4X46wiB2
DR9/lF6MwuqBu1OMVGbsF0QJWGElabNqny/of7Q6dqU0Z4TA+AmZvNGl7elT9lfz
viDV5/pC6z9/Ywuc0YmDDZAB1fxGwwEXLf0K3c7WlFiahjfTJSN2ihp0hyexvocB
JkLtX7xwKYkUqomJm4k9ivOmCjcGeefaE6kDoMtIvPSvPXd8zWiKUMdRywcV2tLF
f026TSV1hIHwxTflUf4AOeYTBrLmXGQgQGVeBt+6QleQOJ1XTZ0G87y8xFN6L/5E
QIRmKYb6qg74Ew7GwYvgNuDFRKfbd+NqXQ6WhuXJ3D4ugwhxXsEqLxCf4Kvr76Ez
9bEgBfqxP3wuEOza6plCj+wfS4qZqUhiduUQWZbTAwzofeCEMAnJreTGB3gIuvCZ
glwCeoWHs1iJrQjMKtV8tUzOAKTv/TS2buTJwsE+SVXRwnRdt8tBu4ReTNUyqKzU
JfCeRzZWMeRx+jjgLX/HRrEIcZcOR3MPjl6gaeBA9La1FW8pVzLPIf7xKQCVNpdg
cFbbPP+rn97lIIunpGpOYzl4JUWCQvFZ6XzOY1vXE59LrrNonfVab7T5gm1PagfD
O06F5bezy4OCBA0EMRGXYpMZf6xFJcgR5Je+8Eml6jj+Q1LQWzsgIU2ZQXaHvrKY
kH51zk0RWhY3/rg4raNQEgLIFgQaFh7oT6e9suyNHnmtBJiMTdDfq0wpaZ8iDJvU
UysrHuaKtRTojTZRlSIQ2e4ixtO5/npGr1DMOOBSWoOz3px1vBVuDMOPcI5m268R
iHstJXC0HiF9CwX//6tyou7xZt2Z5K7o6kijrT6cBIApV6lvASGDU8ZKm+l0ioEX
JyIjgHE4cbUYy4hHKwCXD9ZvX8Na/rbW06WF+0tXkdfHZCfUOZRi5HUlSp94y8ny
/eqwMBAZUDCBz1w0xIG8zon8F8SgT30Sb/pSanpDh8afoAAGGKVYTDmg8ID4ka1F
ZmcOarGZW6MBgIu537yK5E1XiopeRgkasSNZb2wa3qBBH9rQuWpAgp6b3jfPK/Al
dZFcHSuwluOLXGJrXrm7fO5gnAVdnGiL2aNuxBwOXpOo9t4vf8d94qIngLc7i8KN
8QZjGK/g+CB3bNkyK/QSC9McdBeIkBalKAO2zb89zf0XaW+xqVZkQ3EKDJjU2aC2
IICxVOHsFi7YuV4VklfJhC2j/uniRg18sUU4PijrZAdXKh8zY0Lh+WsATCuiySCN
6Xnc56HH4OBehoz2yWwFih4HXEorSPaJSAmb2rLqDt9BOOXHtytT82wwDFZZC2XW
rCiMJrfrg6uJ42Y2/3tc6LhtSYYOxj6SJXZ68fBFuJsIxkgbOsQZGsdyStMwpZtK
ZMlQMIodMxdbXmlkOWp6jpZr550oUlnEmr6bf3dJzaJdto021Nwdfs7er66vGjSn
UYY0LpPUAR7E0Bkdas5M1mUO3bPUvTKnCcMNIRiiSZvyqZ89KYhTDvjiOvnQ0kWH
yKSgXBa2Dh8c2U1035PuPzAxS2AyqZVZRbhuIONWWv36kzTb+AZeVLrkOrVG69z5
2jDrTFyp8+S8Z7MVG5EeYb0VHtQqEmQ7+KvEEN2TAYYjSG6QGph9MEJhqHfEWD7c
JpLx0chYcjZQrvXLeiy0pI1D5y/2GzB2qWaYYIGZOfMw0H8YK7JOp9lioS2joW6N
Xih8cGHMYigXcFHjl6UdwnXNfjsMb6BJovaFe0t5wY0WqG/6WBHLhJrr/uthXBnI
A6PaFr/QAvh5DBX80FmQDzt1fiVPqftt4uaSnxs86m3Xywo9MEOZ1vm56DwLtcWU
fjHfFa7apON8DUr2LJarcRQvGukR1HMWh0YgPBaImY8fg/4pzbqZcxkFG4ZsBgi+
AybUf76sUjxMfcxYcDkOxRrE0Ppe2mJGJHvV/ngG79Y2u9XAwbt+gap89qiSLr3n
YNpxL5bwGW8pJGTC30l1e9c9xgKNe3wnZnmLlCFbmlL0cjmvRx+KlsFXS/0y1ZFP
MEla4ZMrYMmID3ILCA1GNxSmfppcNBzBDhUyP3t/hCp3HteR62Z/MBe+jMqCZ8e6
Ms8RZqfxWbptzY8M7jMzfIpwLV1T2Q5M7HnK3Er5vHwUAu32HwV5uc5GXhbwxHg+
rlcEmycY2x9PKj3TtbFHkABZq+pOtEUasmQse/nzIq7WIOqXQANW7IXB7LwpO0/x
vcJ69PEtKAYcuO4Wa7kieNPJx4yz0oyMbmUM8D+UPZDcf11z+TcfjaNetSDdwuti
Pxt7x2GMgbhmQMj1IdB0d7ldNdeVpVOtHlWGBXGG+6MdJ4OV7zFeGeyMjQ0vqAUT
Jgft7dMN8eWCVpbFAz2M/wQ2z81MkNJWqR2VNsb+LO0vG1wEFzzG+5xo6cXKJjis
qOjE4PJVx/mpzr/KVqHxKVEt4nlSIqPxetqF9/FQkih1kzmrKsCbMnUZIREbnm0T
VD3tp9BCSF/m461OWCDxICOQpUcVRMvwsmZeZZkYEHezGU3We0MaHZQ3NI28R0bw
dJ1ZSV529fYa7R7IZEv0ESG0FiAzag9ijoiKgf5qeVE+UGA8jbjyGZM7fN+sSHfN
+iDnbL3YwpGQwikkWtRMsxtZ7KOj8oENbWTJPvEbwp9aJrtQMqa02UcUIhqb70n3
UVwsHLwYe82E8fKR51Mfu9esY2bN/ofSHBEBmvo2o48BpL6VBT5MrcfyiEPrcQtj
qbGpnSWmNxCnnNZ8yMiRN8rrEDT3fJLCpOxDl5eRjcwGiAEV7lK6t2nXlr2IWctw
yEnn1m4KhiqUwzMqfKPjHG42H9wtvVbSivMdLTrnO5SEQxExzuDoBQFAzJSzzhNv
KxH6XYG0asFguJqEbj452l7kWv1PKBAz9zo90hFRF1wT0z52B+VHprqWAlSRO8uR
4BddUIOUgkNq6ES5HVzi6fxh9/3KBfVU004EJTb1paDDUtCflqIQGLh38vqlICpH
5xoMZD8tS8acel9Zn42TzZovDPpT5UsAqHkWhXlsSUlHJBxjnAA3eRTBqoKDoeBo
AxGEjA6ERd0+ZGgIE2GUHAUrvPZ3SgvWdOIfdyxiamJ1dcwDPwjbFBohORUkc3aT
SVhNC2uqOkmrAXXmkKjmNPnP+cw7HWYAL+ePRnEzecPiF64rL4lT5/OJdb/Euy/j
sJdXnIqnohfPNR5WdEYIHm6l/TOfcCsFzEtwDfBds84VUgoo/IisRKmM9hoaaIWc
aB3mF5d9bVQaEYc62GFgDWgU2YJtFZtFRDQBPYqdhtqiNRVH+uqMxTcsVNtxeWRj
aSn+XO23HrhrG7Dq1aRc9mz4mi69zm3P8NDZSZNDBn+1dnNZ2kuh9Uxc3PDFAvyj
ma/0GaspXNJknP0q1Ch+WJK/JWtKn5WpVsQW4gpfwa2YZ1oTBtgOcgTufbU6buiI
VVTbu6l/bGBmU0sgCNLPnjsE628Wre0k+k/hksGpQK0YijKDOWjmf8yEnkiH+F+p
mn1fgqqcHs4tCb3VtY/G2BLgVqFwfmdKeTYmZxfIK6iSZiGUDVcaqGeXF16h4G81
KsHtqnNdpDJKVevztcgvFyH51SNzL+LISzhou+mduqGY/NcF3hcqBqmYEU6PR3Yr
xChkrzagYgZeCySSbxu75c3gUdfGYQorCuvT2HixVE4ogZVMTcWsG/ZOu9mokx2Z
0p3ciDLKQRdDJi9jVpKXVsDV745zK8PmFOvFmHQ/6Q5TuFcy2aCkJmiZzGt/0DNw
VdTLkPRpBOsP3rZs4+kcMYN7rrqsaGp5L0ZogEnStWOpxna7Kjzp/k3yyQ3k/hRN
V0nMoNJwZgA3HcJKvUdq8kSY6zcX86JLLHB+ZjWfahxJyPoulxLV5S7hYMoLAZSC
fmRW6XB6S6MCcHQowNu58tTOvtoJI7ZjjXhT1GTs3JPUdzEkHWIrMUthpiNkIgJP
uSCpTqQ1yCF2c+V9APeKlHsWGO685bwJYQwgUhVH1bj1TdIjDvi+mZm8LBNfKGrG
XfmB7+VUXO1JVvt5H6JgAakIkDrwNRJ9/IyO9w8kc3oFGWGDW63QZw/BuiIebzAi
zin5GCdh/rmOzIqikEcu3m47JLA/7WgqoIv8H7O+2MBKTmbQiVHYV23NtwGsFFNA
dZ3u/HxKL2xWeNEMewANKy8o9UsXdSL3GIRQjryHfteG5zq+5mW9IAtc7C5v3am1
7LInRe8zQIt5xEzu2ykNV82UFw8QRIpeqtQG1UhnjKvpyGsswhFEt1WG8BAhXeDN
hz7fWYMTZ14NyJXjafo0E8+TXJvHJeaHN0aylpPkzY5SW/UTCHg26e1eI+FhCED4
6kaDJ9Qp5UVzrcjqWjf/rcF61oqzVxsRzRv8YqR8YorSKMJZvvNoW6YMTXVGoRRR
EHC8+Wo3gJtS0MqEFwKjL3sS62UQYiRTzAT+vRJ/+IJ9Rx8i0Y7zya1rvR5rOyYa
4UoPionyF+iIeGOCFhzbGPPAwUcYys/9SwFcJF+JCQ4EtlfRE92SnI7FydmM0q+B
p3W3C29eVQVJogpuzMOTWKERCWLVeNIYXBKZeJDhYjE1xaqWwSQdGFrb3QVOpFXt
vycQ29xy71XU8S5tvd3OsTmSjPWVy34tDVUbmBbwyCUXWu1Dw8npa5MQ106rfQcE
xdjrTzzH1bj+M30k71MzfeL5EwtwQ0jXnBMuPm8Q/7+0plAxT+wHOR+2hb1CCvBZ
Pm+NWh+j22KVxGsXiWGTldfSPmn+HqZjU9xqT8w6YAa+RW5FmPrjwFlwMJsmWnSC
bqyLpdg6edbxDTAWsqfJthKDi3cKlkfyWOUB1IsB+P5fy5ipZt2h3NknHHoj/QSe
2UgNUaT7P5rrRNaCn/0uY9NiF+L45fWPPgVAckPRxCLMJW8OVMO7hwZS76HLdiQJ
VU1MG16QLdrYejZX1ttULGLLrjPwA30hOmbathdreAxkV8em2Th2QZ6PtefntBwc
v4jnb5+NIw6g17FEQhspZJspAMpE8Pq1vCzRg8H1XribqBYeo5AYj26I6MJnOW0g
HBB9E+UqQS12boj11DU4I5oCd2Z2hPzaLQyNSrCntNWtW1r2CR0SAT93a3+cl3vV
9zj8/haHBXSF32fFalV4cprJZgxkM25ZsFGYvxZGwh8ZxFsfrKO9FJsG0a4otZXy
ZcSyHS5p/pOqx0rAEj96cA5T2d0+j2EFUdMlkbyYfgKA9BgboOjgQwKJ5shDDe+D
zMZdX7MRWfcW4xeQTyVYW4B1q/ShY5Xa0LOcWhGVNACXVdS3syAqJWJ2KTKCrOUL
ZIXgWzH76ED+HiFttpc6YkHPh1wS/ZrhDkh1hpRSmt8c4h/p1wFLXT75EuqVd5wV
AsApvoFwlL8+VoSpi848UmoWSRorerTrBu73Qt2Q4XF2t75xhx2WpvSIWGqUyP6q
/BbfrL7MFWYLqmvDUDEBpQG4MdchcsAkupLcseonOl44eKoAzQcIdSxTKnLQwKPy
3Ffh6CCJZiCK7juz9SXhrDQ9ytg2IzJ9nKsgENChe76NsOWUMbVjM+0f5uopPPF8
jS+fE1y5W71nBgud7ZWnEHmh7tcC0hrf59Ypm6hApwkRtFwHcz0htLFSuW0BON/2
N0pLbAzXlzi1WItcNmSAUQLkvgtkLSzfilcW6XnKNHJ26QTZOoWlkcI9WKKD5hQj
XawSZ8yqGrNok0+Dru9D/17CDCD9R938Wuy3GqxCcsWMBdAnq3+egAYDjXBcg88Y
H2YbcEKW/JFi/0nW4Kq//qCPaMsn7bmayoo2bgEVpHhFNx/rsXGDnv/EcuFx9zSs
n381vmmLuFhkepdPJMsZoR9xJoT2AL4NsO1J3I5Z19mu10vkWNQD5yVPiazMOxDm
sI8imdKwpDDTuFatxQDQ8mVYDqHaPxKcXgqVW6aI2R2KFqIo3uB9ZJhDdyJ2WV7r
2ZxGbC+wpWW1/kIhV2y+RLaGQf9FlfhyJDd51pB9jIeoocvrEvY8R+nAASBBRBvj
ySbmW0vRfCVlUpF1pqHwNiX/18gbYyzjloYIWWQH4AWH593ab6mKm8a4/tb/wKP0
rwkD9c1nNb1INWNNrQmAryI3ktncKav2jjvFI+ISrHwbqVfkEpMGYpXCd7fzn7BJ
2ltt7D5nG9wfeW5QzyAd12FHxbtCrWyqUT3RC815BvTLdsWLhsiHUWiO4oUpStIG
jQ0A9EFLJq0fVP2QqjyjD8nDIze0h8+TydOnJQ0k9qRCArY2SlcauEdnGCnINHqY
KOwe3MIIOKLeEVXymClZ0I+xeBbjYgyTUURNL+1uK18IUA5zYYvbkjPaRI48wark
OEjYEZaWWC18lVYixmL7fL+4W2i/C9qJnl4jIKZLm35MCG2vuOcx4+CLRdMxvPbG
1uvBHDAsndVdNWPEhM5uqlN6VzLynluEnvJWaFUAh4zSfrGGGi2e2diD4pY5TgCn
KejMD72zJbiIdy+XfYVNcSSFz1GrN9M6ImBEj7aYhetrGe6WnUIOib4v5hm96XDH
Ne5HMbcwnf5D3Z+ZA5gkAsKrnCFytOHoUjhjekUcMBvgx9ou3U9X8VN2QCGEYM4I
AcYSU4Lid/TklAEQHgyfPX1GOuLPTmjyuwiNiwg1KPYXSsuCJ88IoKaFtbJ/5Emr
hcyKfNPNP4ldbratSR+/DVvLS11yAcjlyW5YIX6s9p1wi04M+wrKYkgp/8cNZc/2
ACXdh1uJ+8Y26HwhHyXaH2XbeMe/8qe/zfnhQzN7TkDrNl0L/UPojr7iZVNh7D0W
Fjblb/ZYnjOiUirAxA0hh2v9sm9tJOAQ26wYv78ldkw0WY32MexDgsfeGekyvhQ2
lERBoYt833tG+lzLFAstRUJ/Kg5LQJWyyX1kVU8vK+Py+uYMEq2UcNwb9sD/+oYd
A/mIAJsj+F9l7QfGmEMgG4OZrfuw1KrmkNR1my1Dcf6Sb9o8Q6kJFbAaUEKYYvxd
9k6NUoepnZY6inFnRSp2xLCcZQBFpT6P5bXs6hUpQxysMFKidWy+i5Ojpry/s4vZ
fngN6cIdusCh96Cyi2BCz6gGWs/A9cbyefQVgDTtrTfV6zdbBk21AxYMuUBsh8eP
0cSSxEe7Ic1xs1BHxhAqYqs2g7ss1G38MUoBTs5XiGckG3cGKd5o4Paud7h6WGPg
mYKuQc1GZEhTmoRJOJLZmgsGs2eOdfT39kYSGvQmZnfv8XE2STMI+WaXhxJhkWvA
1tMIEtChHda5XFTh827XcFymmO+4ORCMTd/F72xDoX6B8DARZOn3tKfLShgW57jT
hCljOeS1hQc69JF1yPEXiRQEIEMgrdphLf7OeKQhpws2ymXH7xvswQuTyF0i3CIy
CUg2etuOqzN/k0LraVU08Xt2JZpeVpuEy0od87noJoM1Y1/mpiktMB/mlAMf/3kc
URT87MpP05Y8RTwkQO73yzmg7hoNq+66gkhi0FXx+AmznRa6LjXSXZjBW6oWfl/A
Bagjx5fY6Ao/OiJIy+OvLHqaSdYSiK3vzeYp0NJSH51Fg9k7F6BqLxKwU1E9Q9fP
9gOcUtyI7AhZAZu0ZkO9zBcsTaKYWb4Ms3J6AsxlN523vxooW34IP8w/Ab0DDKOQ
krUjipGVgUeCd7eaL6PjX7dqhPT3Us/dy8msk+Brpzv7elWwRaLI/CcnBZeKLxDO
Y2Aw2stPXq6PRlB0izSLOX5gl1XGA0DYWL6XDVd2H5Az1pioBOJ6FhQzZ22lhc3h
DzeneNkFN4Y5EcvW6p8ERBUancf7HLFPHqy+bgpk/fl6lqh/KK4aZP1/qhLz3Z6w
kuqFUMgiZCfLJFU4iqwdF+i0afGClfY3T/PpIfrh9au9H6nas8pHA/renYJtF481
mj6xu5EYsLQublHABiel9+qJql8r2dXKrCpKKkcuB42IZMbwlo98yC+bylcBTfVk
IKuJYqVDWKXpJfJLxvohpXrXOFVywGVZuvpEChR3JtnEDYvsLsbFp9vIJx27QaxT
Ttw9LXg2HdolJHsfTlXFTMNifYUfDOzMAyb7r5T7dgKNh11hT1zyc82d/yPejbQY
orCqZJBXqHjN6lNi4i1qReeIMfK0oECBBCptDzZbF3gb2ZEE0uNE1ECwrXJdowhr
tcLRzkpvK9pXQHzZu4KF5yDSm2JPIrDgqFHmHmIKaq0yprVB7ad2qxCxWVFyJpFE
19bTqrt7k3U/94XaQ4JmeXkb/C5RApfXCTWu1Ct8Fna7Z9guWhxYFzUoDeMtZIGS
BJaK9HIhXlRH4zJNtG5SPkpcYzsca5Zl9IganB9YiAUxmxSF3XpX/w2LjojE2khT
G8OGQBTJC3ZZQHOA2MOGo9N/nI+fbt3Z+Iefd4bN9Dy7wpC1JGUQ9AchbvUyO/6e
S5IHA59k4eoD61LaVQs2KeoC7PXwnmXOLgwx2K+pWJERNYuXWkT596FAv0zzUmFm
AGf3Ce/Vh7biriDQNwa1ZL4cBeR820uPaWz7KkwGA0RvzlPM9tb+W4hdLIet81z5
Vw/oR9QzW61xO8U25A9qwUkYs60uDTtNCG30oPdWduNDrr2DcdCfWP19ACjyqY4m
r9ApPZ/k7W+J5Dn9XdD/xUKFt5o57Jd/UtzQRr94cRAzEKd2tj5KFnoeuViM776t
ySozzHKMAcEjgLby3dHCMDuxBgcc/r6bi2n8gxXnfyghPgdJnJzWYFh74IQWm/Vg
bjUO/SFudvangpgAVM2lwhn0x+0cmyhW7Xs+LVYqkT7m8J63hp/SoisssilsUb/l
WKu6qfQKalbV29RUKASP2CW62MMJ0fwVep31415FHaATffgKiSeCrFLPNm0yeh2I
4hWc5Rf5AKuWb9yNCKa36p5sXrRXUYzM9S3hIqIho4GIOdnadBX3Oq+yXZeWBsZF
zLmqWosSktC7Epu/XBIn1D3FPD60homQWiAsZ2t0+lvmX3FbGpCX6q6+qr3qVXue
lr9uryZ9rTwSx2jlJnbYq1HpBQVw+JqAvuMFJhtFPo0P69qVepm8YeaBrXST3LcM
2NA6/um3l4Sx9nT+q/QuL6zyLkHnpbsssPrGEF7GXrGE3Q9Qgv2o/kH7viBbwaYR
x70hk3fTlM30ffySIbzKk8qlPPODpZ8+7MkUr2L1WqJhdhZAfN0c87/cLMm+nSHB
dCuC5SMtrxqgipkFybIRQ4cgEuiEGG0JCHWKqlVeYLk3ZiuS1qcpC/abcJCWUqFS
Si4wufDZuQ3Ljym35vZriPKKdulws8lquhTFm4/6FovgZBCVLpDXYVKEgl9K3ii7
2uq2BhtKzpdoilFoIcTWKZhk+tZa0fTdi3qppc/9jFek3wl0D8znHUZaqHotEeer
UHtJj5yrgKqgJ5yO8nfJEDCHGXEMov2GQ0XF2VoTfB645puarlTeSN6Y8nQEChzn
YIJC3in6LYZecfYcLRcLqea6t6jns4Yk2xSWApO2e2VnM2TGRMnpTCHbwfVRq2lx
RH2B71P9LQ5QAhNVhn4uBWpn/o38GqTRArK87yDLZbC31iploh3wz7mzDhDfREpd
2HHiXvVlox0xeVRN+mJQc2ZwM7OZ57z/AsZnGieG1ODY9aR+EvDyIBd+Z+rqpugG
Ex5IAF2EZZhdbPDKTt8RWlSdrJZw2zF1se0qPDtnZyGAZY8Y0zkhX5UZ4MD+gME+
qRBQfILInqxy+8xF50XzD7n9k7e4rka1jcKfN3TW5of7xGObj/CcUb8Gz5P+F7zO
luhX669M6i0hmmKSpBChwya3C5VLoAmUQIsH9jYKkSwUy6Ptl9yc+yofGithJ22j
YAmBVVwbQ/ldOKO0/DwdrqG14sPuq2UYAZU1UAWniqEjspU5gSps7VdexXKmXSnt
hfoW9QbUcx6HWqVmPJ4EYWMZDUwR9k935jeya+Rr6wHWaUWEEMkS4J9f0g4vwFmU
z4YzshWxbnsUxW/iyQLzG0RwNtMHfjdNp9g+ebRuqGCFBA0+S76Lq6En+hisv028
67vKMfohXF1+HRJRvvfPQuJHLYFDVAxWq/zd8og1PPzm3LLynWDp46wllGa+bNPG
HExLntG8fk1d6kAFJffz9M9pbUjDHcYm8/oYNWRUpKYyYsQ0iL9At+LH4BVOLaf5
9mJOkO8LdBnjmsSsoynqUTzE6lw76LKeP/5L1dgRsbs4PqMx/4ZhBnu8i0G1Grst
drB0ky/gG+ikd0lBqKQzY3Cgz08nVUhd8/9o/pi/y0XVd4fGcqF239TUtZ3BQjp5
/KL1DBOX8aDTJ8W1UIvUirVEE44/R+bngSQhow0K66dJ8jGX+xVRWjEXs3X/Nx/D
zpyzbfQKG6dupEQiPkRUSAXJfVeGp+mlwGrlG2AGrWv2doxGcykcGNtwF02BEzre
puXbNei0elaA6pFK9hKFTKAehpt6MOCj8IS0KgJiDbu+uf3phb+PThlfEupEkFjz
u4qYZ7RLXWuxCSs6bNe3c3jPjHZIkX6sVg8zWxsH7a7sCswFh9DkPPsUgrk+5CgS
7OvLfxXO4SUqsnQw4O3viDC9jwZM1lbURmPN7PuBM69Ke/z2hYurtA5V4LuF8MUV
bLsT++QN5qjZuRbZI/eTEFy1AT1wBM50DU10If+h9fJ7mKM8dSO59eEFKJSdZFuw
adwGW3zpqKYip90PHXzp7FRMYIqenGvtFbR/XC8rMTT1WzRsAzoPuegjmdExf7rX
t3jPT/iYeFlJPFmRUQ8uurnUdInpmIBvG2Oa1R0r32k2I2LjTH59V/oXoxxQPMNQ
oX7xAcutq8FYeSGA39UxQj6nkMicbXt/yPe6T/19FLiuyI9VxWtJn0UoaPxlDbAW
kziNFMSe3hwpYhVOsxQ52ykm9BXbD/xaPwOhnh1ctedatb75xdjjFXvE9885++Ct
QZFUbdyD04t97gq2ybPQEIyqXxokBolNCVunUJeIgcN8qnY1B9PBHAfpgmft09kt
R262zBg0k1msNycmnbp0FjZXOreybyLpGIZAzu584JvIUGa9uklRDGrmIzDZjjMu
Aq2t/9stPHiAfKqA/MeEQd/79nun6kiw974XVpadWrPopnXHX302LAxAcFkFYQtr
N+mMwveN2XQzO4oiIRkR0jnndTzmSk5SkxDQh++tmwDusRQaU8Yo1bMo6YN+hv9x
iJBF+VqiO8Zyt8jhOaCrOi6Qq6Y/ICdFt2ejJq+D9yhN3TjNOB6/tMyMCVxPy5p7
oFY3y0Gsh4CI4BcqgPDe8HBFdIuOMiB2NrjpvoETj30PF7/wH2b2H5wQlpUTEUB/
5y7lv69dc16oP0bNOjrPOSX1OIs8wGlzFLOdZksMt1/XSxNO6MLposl+q7o8F1KH
Zr0HZTfK9A1Uf2nHtpXu+ySmkhUwju5pmlkSRvPLSAhNkWUBZlyjs7bSN7Wn7dSR
J+S9pu1xBDfNkEqBAIR0jMoq5B8WTGTvwbYNPOUwLsWuTyloDXDeVMmDXh9O4eKN
gPxasgIKSKHAiJK6ewOo/1KVpnImd9BT1GVZkxw7+EVWDCNJ8AIpOGpGMZ0N1d5d
T/zyl21tp6QS++IAJtk9aSx1rGHHNxOEhBSGA3H5UuhI0CvtEoBezuUF9PR5fRUd
mtm8514/PbZ89b9/y2Nw7km1Cz378jDaC6aoN2EHpD7smf/5SMXB5cFvRzjr9b5n
mSgtjRVjPGNSkWLMKXpNWYvA1WK6F7yZnU0bp1butHmIcb3DdI/d9ElxykqfLl0F
q+AIISYVhFqbMhOcYM2TbLIF/dTj4xlcGSWc1urWeIbKuY/XJArCbVQ8mWAAr/oh
VjzIngfq88WqrHypqSzxn0J9bpHf/wNyAu9UBocS/Dh/1DKC7BqZekqRTB2JwhiK
c819non/K70aMb+XazYDOuXDxScigCNZRk/EgdmvrkbuQ8C5pTjs3SeDypXdpzx9
I4XC4j34O8sjEzTIwjnTiYJOlNVZnyUvsA5oCgwzEntqaD9PcIBrNDmvOYPBG/SM
J4dzKzUEQ1xw5O80Iu1KzeEh5L3x15V/LJKyn8uMMBiSRFB+sUy6Y0RkckrDIWJK
TV1D9HEh22mkiOStnbxgLPHQeNIC2CN3gz+S5ioHQ6phvmdCivd2yADnIlXQa6Lk
e29ruSMkFWW+HEusuQd6Pta0m+hQ5hshHmIyjOa493Rrb9hZaYUfSCeXCWHm9G+l
6+AnG6x2mygjzb1NfyCvAV1sDqdUhQYrxR/9orm8fYiCpRTzNPDIMpAkJ9arTCH9
D3D8kuKBRrV3fAn3PRQ5m/ZERv/q+E++Y4TzXak235qGgduupsRmCerYfrgdO1NC
BdE06O6h2rFCsQDhqgVaM+Laa+AoOcnnRcrSR3sAqD+onU8vTYPTnLKSbgQEHW6X
CDogXz0QG8M9lnLZ5KTbNhmIBTSMqbbNhu1pwH1o4yerzjgboWnJeeRjhENt6+4O
fcAWnqxdUbGHEYoDmKTqvZ65Ocq0RQHWWx4vL2eYKmLxKJt+Y3ti5ik5sMfVeaSl
aUTOgoJnJ9gchCOqedCdLkqE7w+sabr1Ohg9DOpETbxQEDJsxoWG2nJ03Rncmz3V
Fdl+5OnWZVARtKfi40Oo3RFKAGUyMZio/sUi96Cn6uqVfCcRQIWyv86LAK/IAv04
HUQwiiRU5b7F24I4PwesYVC5q4qJLstVB0I6R/pge5SggAPhIvhvwPBobFgyZ3ee
c+gJtBmhFizwVWyG/SxXLYLLqWFlw5ZsSf4xNc84jDMqL8k1WS4W4jPC+ZCreqNP
Y2pG+QMDFLLlRVd4j3mtPmn6SolpyUESDerpMHpIMLSPMER8r5YmcPIqu8thXei0
zU9KZhS+YV8NR/YS5grrRN7E6St35ezXoBz7JMCbS+imERIoE76fyyNJFIloXS7z
nmtlAWsUMoQZlcwLVBpxoraiQ5NvaG3tJokHln7AhJtc/ZgsFwwIUCdAu/gBIYtz
cdZpaXnEJ64g3cSoT9HgziSAK8eufyoVYvlZwZ2YUwbijbRg1waRX84z3VDfls0G
oL7RXd2T3DQAwQZ4U6AwMgzDFIrdIRbuzZcE+EZqLVIBDm4N/pSJ9fd7zCE+4rC8
cDbLThFE2l6Jc/Ht6uE6H6sQQq/UuMt9P02FJzpiXj+VpSrWt2m2bDdyq3ZBllvG
VLmZZEgt5PRbmureD/GQJclS67wJ5Rzb6pLj1XSiaq6OmMXegxLfDZmT1gEwMxTb
+lKyqpPqkykYLoQQ0yKGEJBXC4HxHZUCt0lCDkZ1g2q6wyBnUz5kOzoaqBk6SeaM
3o7xQgW5o3+mMgoNCBVQcm045yECFnp8+19aATrwb/7kuKRwNe0yx0tO1n+fPpeS
qx32YLHfDZ38tStiJJ6dBa+LmqWNa4wPDfDq3qPMOa4h9tDoWNyWFlih64Kxs2Gs
F8xpXp8RUlpzlm1MqVch1HkECFqLivcoL6zKajw0Xy+e0OzJ2IyWcd6MksJWM3y7
/khCWe6c2DnJLCQf4gs+W0iP95eKOphhxcUbkdQiF8cmroztlt6r/0tNyXvhPyof
NUZpmkV6fIsXGOrEjcUEgXLQ4029+8nHxVadAyUNkJg0Q8T7j2kSCtKzv6NBvo/K
WvWME9Fft+uvYsMe8QM6bqzJsLd5kgN6a3u7XWYSaqJ8vwmSijnk/S1MiWvozxen
FvuX6oUx2udP00LZMAP03IG3QjuXfOzlTwJA4LATw2Dy25Ycf1EEMCuAlZxDcza1
VB9fB/mEbU2zmgnoXFxRSa4WdfQvjxTUTigbBk+63aXz/BkQwfE8kJ9lpf2T+lEv
hIzkefQoYI9R7gyK9yI/lc0Hm4OMgoL4ymKBPUeWm9qCPljo7Utfo3OWX9K7vqtt
ASlo5gtvKlhPzen65daM7OvqucQElbt1yu4dBDINo+T4lT7G+DxfKnjHI3gCbX3q
EX1SNfbL/wpyyQUESx0ZV8B1odU6sz8GUzva3IkH/PO+PubjkC2E9aC8Smk7Q48m
4XOlShkDuE1RcEahpVKtdUPBTcid2egSquIFfKPhxKQ9Ii5rBr1vFD2Vgrl1ncw6
cP4kzoGzFYu57Sv4/3EItvAJ4vX/Jga2M85rHAtjC2j57KeHjBCMx+q6HVBMFUka
O3IKTXuKPHZrIXP1SyrLE++esWmVeDx9qn25N6i/f67j6rPESkMmgGVA7RZqavnu
L5Ck/gjSLf4XW2Zs5k/ZgyzX5rtxViwz+CioieI++0DMBNvOsbRuyrSuh6KoV0Ia
yiUujbcY3OO9u7ZIyqBeKliExdRGN41wW9BkAPoPLlwIsc6KrwAH5sn/+t1jdDL4
tle86YG3PgcwL0vx8iYog05hzCaoLll9eGzCcbD5Jhm3JJ2e/+jhePcmRF0Wmyib
bpeag82JZCX5ss8bpZZ+xxzKwulhfU/gOHxpC3Qu4Ucm5s3cHyd+pxPk932zHU9X
Dd4gTcXt3j5M07Bp8xn/BCgLQRf7qytTc0Wtwyzv4eRRKSSkKZelPPFUp4PrOi4I
ROs25VIjj/i+SwSaqiVXlny0QxyZVBAgAZhWEJkLpHRplyq4APjnV2pB+mJ475Pz
8S/8wltANOG64q2bNnH3bWxNgLh7nO1+5o+LFth44X1ijD0Q5kwDR3jQ49oDbH63
s843VWu2n2QFxHbX7KVaiXcLtkuUjzZQ55rOGJk04m9IdKeiLABe1WpZjscpxrSm
LYVyZSM8S1MdZydnaJsAy2ewDeAsIZn5XmzzK/shWqzWUddg1AF5LYtYQcfW2kJZ
B5PKKfFW+Kqo1vAwXGe3w4WHmyDxRV6iqtoV7Rku6ny0eOfBMmODY4DY01eHjojh
udYRbrXFUkW63UAH2bJYvnp5CaAC/WNcfMvJSef0OgLSZ0KvWzURHYrNPn7+zwYV
vdO+zEcz/TOGrUKLyYabx8y8ylteyfnRcmBQ+Kg9n5V07ym8tpLY8tbE3idTT9Vx
TxG8+PbSgvCFK8dpu6cHxyTInpEF3eASMTFxH7FcSPeowaCU3HhfOApztzQUNLEJ
+n2Jwmy0Ey0DLy17OUiCMwHRFwr1aBgzB8ThQyXxUIaGsqQJIMNzFIfKHAIDxuUl
TSAZZcoNplWkjeDCqZKsDX+hFWQq+2xDDutNvLCzl6KLsxQinibhsYhicbjUxuya
brkXGId+slrl0irzenNDUmgZFmZemo6WcfVRPAhgE8KecXDLsjD2rE85T+6poNNf
vdGV/MFQ8nQujDQvSomMt2xCI3FnIVOcxUE45TzHKIuFCzm77j8ci4eUfDcdnP9K
NYvHVlzvv+VyITpDCD7ZsBTWMQY5Dha99DHoWwnuJnz75qTGj6G1otDco4nEOGlU
d3vVUqDs2OTjqR7DwwagaUHGn1J43T7ux6YDzZo6p/NxhV91GMm/Mvd1QjFJPLah
vWs5OpAtVocjOCqYqCkuAQzNHlnaKK0KzaYRsp4AcdWQDoPpmYX2UYGI+zOV/u4d
cPWLFzbl8ZIoDq68rJgFgUVvqjtXHOC+02wCFjeyu/9hOGNU6o35QaLdJbaPIKrY
TjyDPYmt9s66Fo/4HoygUwcx2GaVQU7EcWiwzv9qYzec1gmjW8EzbXACvmd9gy+0
24q9lA+3XnaT+FjGbEZpsxnNJqu3Ct8pHrSumj925AMTVZ3e1R+FVhTLYV+Y9+2j
QqtMdOLYt9IaWYM6ouOG7LYdaRKjDQS+tQxXtV4/aYl85JcfqkUyG1acZMheEtkS
/Fap7OJJkOF6JoEhhCALB6y0xgTAPW14fLgntijjnm7vDxUE9laiKksowEpGU4in
Dv/BZC7TeOFEwQJDVALXT+xuvYyVZiyMWpLbO3S3bmQYf5yaZXkVUuxAEytJ9oLT
wOUcGUhsMKBQjIDEmgsX/QPvQjH6t3FamdnEEHLanDJAT3SPM82ivietg7E2BXCP
mKUzSFSDa3n7pKAdTUQjI/xHaTgUg001kztiYdRsXL4cbaNSms/MrkUL61vY274M
SFC0hgUhpBPoU3ZfZH7Ca4fIfszWwGXhP77g/3UDXx4idvhFkLB7Mu7IISBfJ2JA
Q2HNYXZVymcjBc98C017Zsm6vIeNLJPCf7OWI+qM28SZpOQRtsgiJ7x42zLG2s7c
nTEjtuk7Hv+AdEfaykggNgG4F3C3yZh12JefDmStwPkjQ4+HbrwDtGkxhPYr68yN
9zBYcdmtCcHZ78GTcnUsCs88Rdd6vfx4AyiBWxVCUL0gydD06HcVqiGdKFLY2s7D
NHhTQzfo+GBEYkHUpBtkxPZBprVMZ8r3XFcrI+Dst1KjU5adGMSXjJqJ21vJ4PXM
lNgoYb7YJYGODLmok54LLAjvjqqgTIbvGA5duhMhqHwL+m2du7AJcOVUyD1q1R7A
qYy8DNQUWxR1ZlniaqdQXG4U4adsoPZm35chTsaIvUfIIUK62eNxX6hgOru2+vqv
tOFUzsNUWIdU0bsrEM2vUQo2IoXx6zmBZ89Orx0WxU9v8M62hKaJHex7HKdeyTrg
JOHR3lF6Rd4Bo/br0d0hHhGefVv0AM9kYkLbxnSxN7EPjjx4oAdTAIZT9OgtB1Ax
pcMmXh/B8lioQTNIZT3LxlEXmEj0DP/4MId1zsXBKiVOCZFa0CUP8jAwvBoxRJ2p
CJmYhNMqxmqe915VPzxA65ZCXqhL0phHRhXRGrkjRcH9o4Zn2tPAMjGEiZJp+TE/
1EG41KjUtaSddowcLtV0N4X8SqAQzY9Br8iRSv8mvpnB/mZRWUQWAF4YiNLWgLj9
dGE+Eg/yK/eJK34n4qKpZoxSatRkWH5Lcq+84nEn+WtUDUswadWHqn9t8pMxcxWN
Cn4IDNENt9hMCx5P7MFfbDt90QI0sduf3Vt0NTH8diBWZeV3bCwk0DANTdiVkx1R
AwaEcjuFi/rzECXncvze+hhp+ekA2wU+yrIi+VFK1mujbsiI9EapMY4uBKY/c4j2
5WQBbvIc6o505VYc3h8CedSQOEQz8fTHKFggkNQ+FWD9cubnrI8Ry1ydodcProZs
g8vkQkJ2AIZMtJRhOIx+otTqKgCIvMXl2yTGkFCowjUO5sPocd+878aNMGj1TueZ
Q9tZgYtRKMx2xt4dKbrmAkkH4Ta9nVoOsnp6jooACgF70tZz3pz3+EdZRjD+jx9a
KM9cjeyUczqW61n8XTLu+8soAHe5FgOH8kP6IzPKiycPS1VJO2/vU7ZGUHHO6LlS
RsEHl7XyAUkxdCPRBfjDAx2eisbU49EUBiAgY9KMF3wLs2+xocl5C6nap08HHPyB
2c/aXjOOfwuxvKXsQbeD8Xu+GsqtpIt1qsigdCXqSBbzTxtAra/g+ce5KuIYr8wD
hR9OwHc52bdT1E335Zg1NF1OkKkV0rc6N8FPg20CmYmrmB+4z/SQkR7U4B3UUSwm
ubwFFMu9vEC8AZhoSOqhV7ES/qeHIEh6ut4WsAuxSX3NAjlqx54ODgD448Pubgv/
Mx6+7vWndYxTY5whG+Yf50sQ4Zc2F1UPEK07EvGbqpdCFSh30WUVT+1tkwS4Lu5l
SHuh1+tRpc8Loa9lYkXYzeemNgP6vYMZ2Sfbo2SNgQ5JVAy//+P4wH6vmX0GvjdJ
IMwpwKWlGkkAuvIvnKURj49lVFpf4Bvcj3OtEB6QxOQA8AUFLj9hWzHH0yY1/p4q
Ry90Xr23xy4b4KmoWqG1etV7bBqHmtqevqLXiWHv4EC3i3M7UBEEoKN7le7FBlMt
bFeG4YGW7wbafLrgTJdbVxtK3H+uPORkwTQsv+bl5ss8ztp2QqOkCcFJNcQVAJs3
mQHZ3j2ePB/yWD1xi9ozPFtyaLt2rimJ885OqpV0rhXH/OJgcWmwR7nQHUOS7AQB
gPUpTzzhE0IAP57z+Ye84LVksEhjf9vN+Qwwk6yL+k9AfA8VDslPMvrE6jRg120Z
kNRz/Dvu2aF3fMk1GFUjYaNDIa+VmjSlO90WBh+Hkfb/qI6ahG9PZlzwfnNUMSYi
XdcFbRSBocBdpDGGDTc6aFhw9zp/5Yso4yPWH/HiOne73uHfshKmmKwUp+7vu0aM
x/mmr+lIGIOT1gEtZwMH8QpAC5WvnE9HRxVSHoaxAXklXbehNRwoUzSlAKthbaeF
qwpriCgjIQ4Cqrb369aSENOZn/FIpeKnnIO42ILG2QUQLPOalu5kjkc+aMP48aYw
HiNkdoP3LR/LkdiGYVZsOLi8hYr9Q4K4tsPz+KqtuTkGk3l8nBhUrShU1ffanzrx
nYo/NkP1s4hj7mLqlo0BDSjotBAATuad/H718c+30R9LT5Vh7EzUewbz3yPZuu3g
ADg71hLEL5YmXdClPPltzLaAogJ75HPdw5Fps8gjWhxsEVMgdLWCdH2q+gd/cGuC
kXqOmxZhTXLkem2+WbPdOvPT5X6EZAclAUz5GzbrVn4VeeDqHQU1XspKGEdNe7A4
11OWp6p+W3jIRoFk72JuZJFqkDSK3fRyswrMUHLQjMTLVcUdcnwKjWP53WX471lt
8SVcufhjgkOyM9I1J9u54esoyaaV16eQpZYyLnE6zHqetIdn+oGty9NM5+PSGwlA
ulh8e5O7H0WEusTG6KWbZ3v9j0r956703pNUW6Y3wjuElfojw2XJFTg2ifdIkonA
vSAImviNm3cLfwfovVNXv2VZm2SW2vv48fDpSjF3hpU9+cEuoWxgGFvtYjWM7liy
9t9e3NpyTOOog2WINPuRh9SFcag9/ITpXvjUMf8x4F0CTlMjylbg5hg6T/Ivef1A
p5ujV+1DL1LZBQXRwGfArIBecPbNvm5yQwpXZYLXFS/MYZXcdD449YhtvlGsUuSz
qTtgghCURB7mhInp7vDqvKFBKG0Aogu0bL8E8jnrTmAHw4hCZHzP1C3QyDZiWJyT
4Vy2Ei1BCZcciMxMoTexQeDmwesRHRXfayZwkuGKsEwa4qdAHFcApzKlLWuqgi4S
O4L3ZWkkf0T/h/BKS6RVZ23JMfVbu4LuPWDHhqQWOiRiI6iUxT6agR9UccdbXlQZ
Plf2PedBsdyQeRb851k4NNXQCD+ecspmB/NFqq2vnkZ/KZtn8/B5TYPT0G2q7dIl
akiydzxcrMN0XxRDB+009JZi00HcVZ8cZpSqZT0e2rV1TPMYYCvcjT5qXtBAWO2k
yInwdyzX5S3WGichRfHt3htAQi/5BLLzo2c2Cj1LM6zX9rDAKd+rEvURvFTEOi+P
MWb7WEhTtZSGzUCCx2gUmF1JHm8JU1BSt+dm0zQhMF0Zn8YNN7M7EjIl8u3N7qeb
fUDsy1Z1xO0IcyPU896ntpvzD0r0TlvrjDwDIiwPwINorxf4swnDzK+alr9dQORo
waARporXplzWaigO0KytWbUx08n9Vo7D2qpZ/CS6MK+A0T4tjyRjAp1FGxxjKLNu
ZU6Sxu+x+u4gEG33ogzD5Ng2FpXj0WbZQxkogUzyBT8l5Yw03osOMlwm/Bi4ZAev
qq5TYaLvXv4wAB7m6RwXnop5lSHenjzDwTbECQWofheQTwjoL9bfYTh3+EP2oKET
HkMJQar5ME6yh/E58Bgpo83huOPt6JCBHb2MbW+D/654Hp0oT6EDBwOASz++bok9
rI6q8ugOH/4fYVLIjF7hFTJEpPIvcwUruCXWhnXmMgZ4QLkva2hWR0Z5IKk1wzW9
W2STjcawTC8uf0iduykhjJ/Eb010JFiPKMwF+Wwj58lhljZVdrsncFeAYITvpeoO
uRL5IM4WZlpwF7iEd1G0hy5kt9qWYA+xvmG9+s6DhVmYhHNXP/qK+q1WHlrOMAaZ
GDYbZ5IjmxIrHxexCDOBOiTpd7Fo0HQp0IvHHzcMLiotllHy63haC9K8DfZPVhh0
kt9+Kn2GL30qa1Y1Lm82GlJdFxdUZGCXbUZf8D9rGv/bTVkGTMfws3vPXRmyWpjY
6p+TCmC0rbFZ0Oi7gLKAt1Z1UrIVHbgCNRUrOS2MJJpAPNUM/FoBVl9rzXubkBPK
9BD06FBgtnILMUNC6rFZt6Cbmh4QOmnmVegQoatzObAr+ydkKHKUMdxzRb8gezxX
XVMsdaC/QC2tPHtzS5dzqWOI+nKkY6BOt2fGq7nHA9PTfOfnlgIlchFlEWFrxqmz
n32UJCF9OWMHt3Sv2i7/TtEjmEh7W4NA6Ej6I67qBLSO2vnTz35oemaVnIfQmIp6
K6BCiwN+XVuwZVhg5dNF10CUjsHPqUWunvlJb8DjVIr3w8tSclyJ1yjGzSAfU7j8
dS6wl3uJ4ZMMuu5f1TeEhYlG/6jYAvc0DcjpDlakfwgSet8ZlL92DZAA4UPVJ0O2
zBFM01/7lbWYNktUujq1Zt2YrdWDDybxJclZYDwercTvhG+ZDBdt3/7/EKb6MtHW
eayNCfpU70uZ0QKk44jwLYucsy/MRzzVSlQj8zQS9CiaLq36Zx/6GQhCWnsRGAl7
qQfsLt0DujW/t4OwVM09nmHE6S/5UyCxzDrZH1glA0YP1V3JRE0uOVKdaYyntMqf
RcOgR0NbA37dR8QQo2h9UjEszgNw6YMhG3U/lkYxRE5ObAwnblhyCrzvlsyYQVSy
DpPxHrmX9Lt0qrbN3jP+fm6sm0wbp1Kb/QzJwlYyQs5PJA7ouoxLx+8P0pPpMpLa
h45hmoglav1uqY0vmDBmGMCv/IAeQ0CaKERMvvopQhfFEwWgakZWKQKL0tUEIR83
XsRAqvj4RbnaHHZHZPwuKUt0/aVDHzCeSXN2zJz0JAnfBLOwiCj0nyQECnZ/nm1t
Lorg7OK09jP0x4o9GN2jzomXckZlxqBH6JR2OsY3lCEmjmpReexCZWSnQ/UP/5Ef
fpvzP0dZXsN7Wv/0xlTW+GmqyF51C6KQVS7DMSD7lg++79ICNlQrHPURVymceE7m
yd54luR59NcSj/Ads6nIQtoRBsb55s0wj+FpFq/xGzGVWojfvUzpVXwHfHxf/IaQ
0RiOX//BTwT92b6esWTI2n8pVBWC5iZvwRyK/Rb5l4bIK694h09t5tkLc9nBniCN
5AMq0CLP0aef8evGW5HO0WSr7ISni3OyNBcZpsFApU+SL00D//XunXaLlG8Xn/xw
ccsKSZP0ob1nsO6FeSTG55Kh3L4Q1pcHZvrro5TKc90IwLQeYlNK5E2HqFvot0c9
MzatvAAZFgnZG8ecJLZhdPZ9I/DmlbDIyiYOqqdvFqTKV7/CYawzB8vGTirYNRLI
gonGK+1hpQAz/3MFepZHuifI3Y52woZhRTwLfVGA0mp5juN4IDXHbUXpMRMc47uO
ZUogvMPCp2Nyo2YQ8p4KbT8EEfoejqTErd0ehrxVnXFg4nbOhyhV9cGF1nAwTQUl
ngXmtwkntQXjoDScwGEZS2mCYZH7MR2dVwJgqz2LMWbQ5Nh7cP+no8IUtogGyiIx
sCsmwrfvSzE74KQPnL/xT8G6LxeqUEFFkpTT9DPmPZYYRIHAUvaAOuFn/zYEusDP
1342n2V2G+7v6csl/ci6Dw+Q4/Vm9RWPUgb88/KpOMMePEbszE73kjWinI+0jEgI
Y6TPwdwPv8ujaKrCgUQ6u+CpfcjaqNUB7uCCuVT0xIPzfcuRaq+30mdTCxuOn9mN
M72gpX8SxoaBb70CRH2cstWN7a27xBgvWpff5FHwItqf/N4t9fZZ7TOFutXRaFiY
ETCzp6BZqBcOG00v8WZZ+br/xgy89dvBMZAtcQkP1Uw4WQv41gHXNpdpIsshdGIo
F6bTEMjajU2pSZboTr8Unb2n0PteDhgoZpfBJv0tj7qJYN8bpZdVMq2ONvC0CO1s
j5Qj67/z4oZYPX47kNxDQnsOHaFNDGq91pPE25weJEjUACrSm7UjgnG9MA9QjUqk
9shrYIudJhVa2DVqU6irmFFyX1qiq6kshfAlkyxIh8SS8l2miX1HiqiW2cI9fKbs
fq03PUVJG/m0zAsib94U+uewmT3IWRCca/98qA0KICF+hPLqhAq64nXJAiidTZaM
6gb3/nt+KbvzJr9Dsi3x+N3bwgBaECpR7vF9B2hyTRbmsA9D6GX9xulUI+wWmuU9
T5tFG9l7uGDIpjl8ZsH6mK5mx4F4PyCKwZ6BUYJsayJaSxcrjo9zP8BGeHkEdfsJ
wvgbE0ipMWRXXAEwq5XDqHOoS0l1oMc9T1HP/sKyP5HuzFOqtnbYyxE/DMRUQiey
l/MckQ9iiuc93UR9bR2CnEyJEM1drzb4xv4FZzGZqWKr5darI/4XKq2Kf1BLWygK
i0bN0p6LVDIdM64Sr/nV7Q40a7/MqQvlm4+ZNDumaZUETo0P/Wo6WJobpZ61to50
6vYhY/bCWGCLO6rAl0RL4gmDubCeAdJe28PU6ehFJUeoWk4gHvUurEyJ+qUMUB64
SyC67XyJg95Hqh62CwxdvhYjhs3jp5iiYe17xQ28EywkhkhAkrBJbA7fJxCSDSoO
peuZ7AdMXyb/KuKiTmz6KJtdFyS2D+eKhEEBVjcvyvOkCYYy2nVVZSkZezfolrWn
HXA3XVRFKRUkHj/8ZES8HvbCs0JfnkfKYKJXDdA0S2W2hu8BKK6TZsdpVI++YYjP
WVoNKPx3u61L7azLQX6FHGNqCT/jGpSMdotU/i74nnm4CYb2ZriyxemV3kA2rthX
Zz3hxY94n8Wja/b8dkshDhoaT+SO4WTpet538qFeA0640RIUHlkt6Lp31W77/2q7
6sXEowQwBznPgJpspSkIPzWdgF5mMay9r+v7+Euc8IccwWwFJu+GK9KSuU0dZ6ok
WW7bCDtCt1BSasRDqPaO8ALqZiYxB7hVoRcC41zxabiuAG8QUeDgrhxQW+Xxccb2
XD2sNY2H0DEpl0pu1i+KLIIMqfvaN17U31d4p3QZfccc+n+BQtFCXHNaXkBpohhv
1LatTOhGXBVyzgJtx+FLq+uIcWeuqUGVmNNyfyoWPviOHK2e2uQZLN5fCsbJGFN5
18MqHPqr+tG8JHsOwB0lfUg1iGwzMPU/CnuVEZJaU2Lz8FdzbL8YiOVPyjL6qNxY
uum5UQeXJ2+S+E76+PXKK/mj1e/j5y7g3cFiNOs8TVUukuEcyGpiPEwxJW+aMMCK
PHOKklJzDsWEtwKA63i/2mpKk2RJ7hC6FNvi/8ZEpQDBLvkxWB2KXcaEP9Su1RfM
wD2PAmXCYnnb0Na3NfBHmzBCmx1Ck5cO1UkKUzMe3Sk/7/aayKIzK+Y3qeezTGKK
YCQITnKS82sDoeRQFPtRFMjyfDLlP1kMvfAsMnOBeGTxZuWsYtcbUYCXJGe/Sf/w
qs2TVp9fSl7beN8qBuG2koaCi1XvpxHIYSq8qhPqwy4zzuR33DnBqc6AIa8NvBw1
3jG/d/l+ALBgOJuSixYTnoUevtuaXlB4psFNqvrQR3l/9kP/TWgOLM9R8FzubXu6
zCD6iY+IGRKX35cU/lZVydF9pwX1lOu8c6YrJ66Enh0/19mmrGBrVUQ84nWdTRfh
QJ1Nz6Td38lJb1+MMTUxcOZkCt+3hu3X1jestk6ScrFpIpPKrkvFXz070Jk9emrE
6v2dhqvWtxSKOdrMMsD410BKVP1uy5yej6nAPpsjwVVrtYLuohc+fhbcKza9NAoz
WMEWQ7qIQEj0unBWdYzO9iWAObOj49RXCgJ03JAY4JBUeiAgf/eqwZM9SgYSUJxJ
gnpCWolx/NmX3buneLkicUwupW8lhZWARs5fGqNwfBcv2r5W3NGbut4yDjXOfwZL
IX2JVdufy1xUT+qXkOFexDcKjcwkClR2eZrsY1aHfaN81EJ2BcYWClXSmCTiBi5q
31/lGQFlwSoK3st+SK03XluTBjYXszZv5E+7SZaMe2F75kaJr9/XgIuqCZZgbZ5e
odd10Mtiz+xfjpWwZR1IkAopciftdk31vaWUbalR6djsQaCMJUGm19YFriR9SyLr
yMPFJUkX8frrix4PCRPkxKYLQXM9JhRmOzhk63eJIf7jB3BJhTWuRYQGtvSS9nFH
sIGDdKnV9L8S5tjQ8KyS99vViGViQ0UNqf9J54PsgQZWkOyzynSpBfAjlZZ+KR9e
TCQQdMuV7oyQ8ZyZOdgGaZp3RejmImCU+5GN2taZQ+H5BXxyl1JIJoQh4UZXjK5h
dpauSTq3YSbJ/5LtCfSfgJMkELWBqQXh2lBMkIoD+Gaes8V59asiuJBxU/ecy5n+
Bp+PPAGIgUSKkwf8HLqnfCi5tYtD2mwA59vXHtJ2vA5RwMFtOTy8VeE5EYke5H3N
b/wTJj0aakCc3+VHkohiSFzu2G9wq82K6EeLlZV66CLJ1feDu/t2m0IlTo1PrpV5
1hfVlOS6WYgPqv9eobbRaTG6dXgrMkO1maBJGHzQDKIACWfHuu6iyx2bDiB6nKoa
BhFcEqVltGJYPNLwbHSJLPENoumyo04oSw7DRxfGXbsDK4+IxEVd3aqvKiFvqsGx
FTD17X+WKZnwzrm1zZKkU9OATPqGzYNNM/wl1sR4+oXcJm/Jx3xdiSfNuxa+vfUx
eJRyP2RU9B+XEX1A6MefH5XoCoZbosVSnWeOaQne33if0ab3RpHystrn/xvCF/Os
qkZgR1YxC+Dg9iY62i2+UbaRmS69LgKmrLXbUpd+s4EloO8QF3Y550Z8rFP6DaAz
QfBA0PSA3iCxLob/uiZkjZtxyjypcIJQmOxN0E9UfoWApWlCwuYfCATzEVaWq7ep
mySNMd5tkx5VawsVUlgONF+AZDn08ifuADxVtky1v76PazyaxOpMCj9qL74lf4sj
G9rVd38wcwdI1aP6MMwU+cjDC7Wtk+UsrfFlpzO2aJ1F3+nOQWiVHAQY0hXRvCKp
0nrWPwfnq/qqOnseH8gPwzjszcaY+zFHtIsNh7210zp43C3uyixlRzJ8lSI8cb3E
DtErZQygSLKToi3wtdyKC08YrT9jVGyRkTpT/QOIXHACApkrcP2KoRSnJ5xZydXW
RC8qFHTvp8vGpj5y2XxEnhXFgPnIVliaVnhtwVoJa6TBXd8vB0P8eglKVmT8txtk
ggJ9u5m9WeX3sRSx+OUIbnbhmOSmSJdPJLB/JXkJqfWXTLQFFDb1zfmt9JVHQL2E
Z5iiSEIf0++o3TKz03mf1fzVUEKsHbsb4qY8/LFjioEvvdZMwghmW1Up06lQr/tj
DO4mBSGDNJz4K5J0WooKm7Dn0Kzwocu2GAQ/cIEItKjgPNJ99pfM4yiRxCF+VmB0
7VJv2o0sUoAFgoSfLbEY6dbAZ7kAIqAFNgN1MZmqWxBoDPqPnCSOvGYxMzzP7bEb
bJ4yxVGVEoJYHTd5Leuho1s/kN9AOe8i6LqQZNFXUYO1ANEYt5gYBmxnw8HzzLX+
4V61x0/BCv8IIkkTGDZEBYRieaGsMzzQ0mnQOdyy1+lfKPUNcUJqJJbhHftbiA34
fQkyjXDRbKRsCSYs+8WW48Ljpt4ik8QZPEFIsToQpICGU5Ur5ohrP6DiFkswXURA
DGi204bimTt/oOCtHi0Yi1AT6hpLU/YgfIJLkq41MBRTH78YcCo8ovvweNqXKPdv
sj3GNE8o+ohxvy2LQ1L7OZEWW2hppiphKZhIj+8zFwwcSRN9/1hXPIcX61FURt//
p6psCuONyolXx6EySRnidS58vFFjtfrv56zsIciHM8S0QkG5TvzXJuGtHWN+DreJ
9ZmD221oZJ/MNjE5Vbkj5IiZmnD3jiKfm6AH3McGha8hk7ejewN1GWQURSJlhkgc
Qk9WQszX6JxzLVe7Hk68tmBGfLx6pw1Xt99M7+3BhRM7dQsOB0S1h2rpLwfagIGY
WFibSyFQ7weHCoROHlWBKWHB9Y3+RKtnWxQEn8A+poM8nfeLVw0UzwU4w6rBPbKH
jUPl3oro2ekwOkHwMb03gtckjkU8X4Ri89bQmgH2f9ZJBOH3EWPMH5MBBu5VOqK9
z3vAWyqdu28pGPv9B4ugpjKTji8g63OAlxJM8galPFoRCbAQt0Gid/zBJ11Qx5Rp
F3m3pww7giZEPxksBsJxoecGEptjtR4HbozetaeqmUVEQL1WrvkaEEVocwe+hRSb
1y8iHNdvcJVNYHnhsQujJsggVP5D4qglvf8135Hfc9NAHCqQ6FHv7RUnVTiemH6Y
72L9iPlGDBsfV9FYA2VQBnL66gSazhuymXr5zaAPaC+lSvg6Jc7Cfo6tP0kGost/
4u4vQqQaki4emVAbXpM3C0uyN/Gk6MMPRj3EU7biAfi8lr7B7og6D2ki0nMhy6g0
SLAU6Sg8rn7Y4eSrHolQxTR+4KR4mDD52A21UpCKmtOoyOMAemDUTNg5XylZ4p4g
SmuI1cAHO94Zpj2g07lhBrxrko354+D1wrUovgjPcp66BfPwpyE+SU62Jnx8+f6W
u7xDhMbCq+ISmgqdBmHXgK0iGksaY+YiSaIcmPmn2PXX718JwluoxI8zQYXRGsq5
masUb8LXpdClgtcpSPA2R1Y4l7YAHLnc1MDxI/2KWEgIA8L1r1HMFUTe2i7aMnux
79o/rCeBWR/fowfs3a94zMtbLlFHRgTifC66DJj8U32yx6CCVO4smeYwqOiU+96/
jHg68aG/yzcfa2HjxwC7RImaQiSQ3xcYazRC4/3hU8NadFc71hjzEM91ucC+ERRn
f1WSIH3EVzW75IFbqRIai8z/l2mo7JaxkBcBaoIpyRhrq1melsky8PZI1fVEcMSN
FRCBpgDMsTRg3dMIA4tuPxiXQkgCXyWmFffZcdpJsF3686QIvwZNQ48H20LhUijv
rD4fOezm6lF3AWnPuNwL3FGMIK2RWFwY3drVnWe84GcJdkbGkQyQ+KdgBHRMCoPX
IDocmXHuQCklpwoTKQgKGyVESttaF5+NUdWtI64bTyOL7T89jKw1WeLcb2nkvVHZ
Bzqt6WwoE/zpv4Xr2DFMtabQMdQytcZ9MFo48p6xG8qTMQK8D4lFRmQ5ELUE3Uaf
R+8BsN4queyXXg7ApO+lsKfW+NRMij+o6c9tbXq5VIcYBvPP5tZjZ6taiNcNigdL
3yFJQNAIYTBWlri39nQnE4NlC1gubq2BWvYMHU6fJCVWeKAFZlYYy7ok5bQxf0WK
C1qswXSqPQ3m7V7s1eVREQUzf6xiz1WZ0fG990aSs9vRSznacCSYhqIyMYGa7hSx
iUnuifIEbOFLUrV7pK4p/LAEeBd/AJn+DzVe2avBfH5d7ZyYKvy/rmrQeYa4aStu
rxX3dOeyye00/asRlqo7gBUT/+tMqIKcKOqzojBQiddWWIpVaRTIcrPvkSrXiW+p
UZRMb7Vczf1YdKsDD/JTUg8so2E1IJH33ghP6gxBVx352ioJZO6+nLBxF7i/klo/
Jn2aESfNptShoBauBFso5aTTVVzM4y8Xhd+5gOY+KQ1Kxa+EuSh96aT0BQnlV9Q+
vUtH/LFiajNbDa6q3l5ILUqdulX5V/zGXaUhhAP+s68g3XdzfCKS2vJA/53QXrju
jBbrhKQBAq1/+W1nmucGFggl+cjiPZ0TotDUcb4s3aywmkfLCaRuRYjULPNYczFN
QUQb6bzcxlM0qpX5NDmW5GNhn6EJBdKjOw6WV00OXaFJPrnBsL3pQolSjQo6EnVX
ZzuEntf3Oj/lxljObgPDX6c7Ih6j3BnGujsbqSWMvKfyBTud7DlaIJv7N1yYIyRI
swew5ZyIHJRjN8J+LjvatQyArGuCqFJ9rPnmDRzJwiOZdQ31sJDCJZQxNLMz98RQ
twqweA+g+fWBOyFn99IjQwdAyIk+N0m52H1fsZoXxJ8dwClsa15mHkS+Qf9iX1/I
5gqtFOfDwI/r6zKInazm2/FguA/p6sDVhv05fAkHosK00j+5U592q+R8LmxcmmfW
xUCr1Y1kVeFGTLU+I2IdD9SezVPIYk1TI0DDsDmV+h4HoVy+E5AkE/K+o2pNwlBo
Lo8WgJMPkmfz8bm9Ojk7aQUCzG2MGXYZ5QBtoXj/iSTbVYLNWxe70XVzDzrxzLmy
aOZnOKRJj9tLCcIhp3TK2nNz5JPHj8Hg2lMlSub6H8QpS8CsRG+hd3jqaKwjyuSO
xUm85XzoTlOOMuo+RS/4FBnQIAAA1iS0HaiW60zVX2m9hXRjmWZOTkpJwHcoNhpx
4CD8BbLkqEw2GVFpd8SQE0TtQ8j1xNzz3Mmm2n/4w21LCVdD6Sa2nQXYmC3Ln+xa
DsXvjS75CP08hGZTjjxQ5xzzg4Xd12jkRtSRHGRy9bifsW0UsG1e9Dyt0L1i+weh
qAZ8/7DYyqILaAxT8ARSKuCJlmM7/KOltE3bG5VS0wtSEgF2trVoe4F62opVL2DG
iI73YGGHx1B4xFwXhmlzPqk5ZSfWtnEpDkgVVLfoa7jeWD+e5D41doQZi22f1JT9
j5xMC5aJrgM1JM0Dzcw2iXE9ohkSqKTrhKdvQ1wrSO5iDwE5aUZkRg/48O/Gb/R4
jCQCVTS6alyuQh+oWSpYUXkCDUgTHcM5gZJhOjBTTyxoY6LZbxi2XFwu6SnKppZF
1ixsoxnyidaAqIzRePmOKCFYqHG95IZsyfbqtm1T8uZ3PHiEjnEnOABJZ0EwiwDR
tIF87F79Vfzt3tngQwni4TJMubqtbz1uzkoxGNOhdV/mpOrnZo4NqgTU1CAcePlF
m6hUNVjEK9lrJlktzt8mqQ6nkYNQx6nbGcU5m2hzkbxZT7vjuONMdbKsHkldRCYZ
856i2IcEiMILgGkGvuLhYjfhuVYfruh1/N/0ltNFBQgC9+hz1fKAJpvr/9JK7hG6
qFmPeNsFdMida4KC1DjX5pecjXjnsmXPF+ucqQ25cprpHe3RUBO54xBg35qzxwWG
jlK+A2dd6R+K950CYdaUq2gaJnNdTMBPPXLodcDfQFuSuM/o9rrzyTlT9RUUFYC5
fSK/h3K8z3DoPjt5IRljMA/3yo9YdW7VB6S+cp5TMpRXvBw4dbWkYLAmlmaAo60p
Dxqy3PRNWNuV843y4GCN54tYARydYm7CwXEMA82sX5tM4tSglCrQPJmgaTcgsryP
Fo+Eu93KrEKj/ZoiyJFf3+IhC/CbddxZxK3udWLwKNR+I55zcB20K5yMNy8DmvBh
6tZr0cbkFJJfPsc8wRiC0Tlia/pL3bOVPhfhzPdJH8OmQqYOKOa2YvnUR/xHbILT
P+Db0gtnHglX2JvPdJo+GE3pmHqmUrHgThnc4fyRQS4aSMYSt75jG1U7u3FKf8Fz
ibh8riEtmZrm+RS/pz5KH+dMQ7QbdRq9at9xaYrpoyvweDwCPi7UDT35jo6IGP2x
m2Ysrnsj8lzuwrV8PxSYDHbY0mH8LFd4NnMV3mmX4uvgrFl0hG3yFHYZgp5koTcC
6gNWaRMU1VOVPGXmHlOQOJr6RxUDPrKU4kHiwqy6NpoSLhOefpqtebKwydTq0TFU
LwXijVZySqkrzb8vkeGg5zgyEvKLEDaYT8Ukx0/jZC1+WhkAt+/SvqAQVT+KcuQK
FvL9BQi5gXFyahTa9ksVEFtlJYjRDGWp21WG8kHuJC76B0OJGPYWAfv+QlkZSqLe
fL3sZqNYnURrWlOPcZx4qMCpGtyk/eJKGSIiHDG+R1+RN2oXOWtVxxViSfQsr/Jl
+QywrBVsdih4bDboQyVlM/9DNexkoDrUibkAOb2v+54mcIfPMvGL/TVuODuxIqQm
+cHpC5elUWEYTnBIESPpEIoGkR5xKMoDEbRaVjvOAkB4K0eHMJgcG2jh/4RCi64A
5iud3+mu0b/0++/CXp+eCZIMedxyjqHjJ1phpQlty8ELvXLY6g+kDsv+eEsSdFpC
gACXU0jpesZ9PUKNdufnLpC0fSoep1vnjrY8KEqBKdzWMS8pOhhwHY4OMs0eeY2W
uNygagGeev10RAJXEULBxeDkModKeZNS0lq0QN384ESL/6jBafEVGgNIr02nUYSY
PahXKQASfuxUL456NQOUXDTKZNqJ+2eHDRE7sxGCOJBeafHVvrHPfbBz+5P4ZAPW
bSSHBUOCpU2bsk2GxVSf1K+xRTYrSz+bXx1U3RtEwz3elgHFaUuNGT/uBfnF/bdj
f1wq+4nDOr5NNy1/8UlVnj2+pm0xo4qtjTW7xMM7JaJlZ3Pa0KCwIMQC4IdujrV+
xPwtp+o/JlCM8ohW3dNVqRriBGOnQmUYoZfPvVW10GpVex3eCslpwd1mMRW/08f2
Jpq68ooORYUOpEVS8nsZUjuw7c/eZxLRUwL4ykduNHmzkc2ivzbh6dZJrFUkB3Ca
Pvnxmgan66Yp2ZQFcJK29ZWJLy9e2agYoYQi/0tKK+blNcHCL1hwKyT5YqrSsHHQ
SBRgr1Y5tuo3DaxEX3sSkltjfCCSL9Bnav3WNQlmUsuGzuaoeWl3tW7B+1Nsta2h
lsg9l+0ZQWrK8ROIVG4polOOqoqziWKTpEpQyIQGYIRzw55LowLJrhfE+OGQ9dPR
r8vBZURhc5yGg2ZFApIJWaTn/WzZlLd20X+G7kEh2T3WbCtEkp4P3HY3W8SaiNYf
Zgh1VOHokZgbLIsnkiOhagtwJxDgdSpySMMR77WayeNfUznPXmSQDDrvZ1AAtZuU
SxTkbdJVHxx9WKDrhBGBKv0ayWWBuiBQhBHgtkrHdV8H0UL/+wRLCjnpOxfRoDX5
JuFZ0/ShKWJE7IiTFeeEalM/tsYC6KsdfFmIbHBUrTCYjn+y5a3u2rZ+MfzA0q88
9SORUD7DjfbyTQzyt4W9e74QooAttsyQxAqgY9oht9RwhvWZD6LjJgFH/SpR1O/U
gp2s1cMaQVNBTypDBpO632pJpA8yEyymKWlb9iKOjGMwfi9HaTmfhnfYEHZNsPeZ
G6UBfh2aOcrKRRKLf8Wll0xuHPkPFcXR/Tw0KioO5ZStcFLfXpo4GFZC7KLObU8b
FEVuGXvlPpknYfJH2XHlbS7aUJHHSZDg9KXYL5H/3AqsP5PPCmMDC6JVcMwa46TI
DxpOO0L8HCyiVbfAvdFDfxZf5EPRuGILo5OIR8m1c+hOZohEKdpqtCS5Fwuz+gvS
Z+qghR1KJjwCfAKWjOInqr5OPmB8CFMamHAGTpzJUhf/Szi/TbRG0D2DwIS4B2Xj
MS693/qZoq1JXJUHSd/dgKVIyhE4DhY8sstsBsAzshUVKba2POtvkxe5ohwTVpbK
+uY3rLM5dFvzn2OCxSbPPpGltSlDl1A1g4lm630O0rSg0nhOeeH6orIbWDviVy8Q
vxVVajVqtXubUk7CQg50pZA87nsDem4DaTi0/D98iZW3gfFBNc7sB6q+nRXQwanG
Jc8bQ3bYgPpxX8DDJUBUv76eaHQ9F451O2NTb8XJaFLkRJcBzY2YB0nVtG6bbFGF
n0Askz1SkzzlkpvcoA52Uwru08K4vLcQ2LQeMJ9BxCc7NApWOMjyHJLl2sVJWX1K
P43vwXxnfJPIPs2Er9NvPiuuPE6gdWvAto6cBCLjX+lNqM6LEfsq0FEwhYjxCbqQ
HffRHSc+6qGqJtjpyWCiyQEQI55QdH4UNLl3PCVoTEe+DfNP66XIDBCSPJNAYujF
PO0sqateIkTATgRWqIY1w2VK8peWJZyiKLwce1PIRTVxVdwjGUUQun+mptDlclhw
2zMBv1vCv2141xoWKwvkYZHW2Jc6v4bsSI5KF2krjZhaboIqVBrPKNKhy5IP865w
WgZ3ODh9jHdX26/SJZpjwt6PKh1fAZdFZn0VtlZhcb1mlxyweOMI2BIqIbQYmae6
oLFXYbkl55OecydmVwwo+BGwXZ2c580DoLSfWCWJsOw70jR4LLHE+A69RidNQv5j
LwV+Zx7Wz/cmxmszf7D2Y4pMM6RytimaN9bUNnJFxChEHkMClH/olQrJ/bndl7W5
P2jSpHKNSIWUHrQ/rX5FTMX+CS4GqBxzx1Oy3NcjQkQg5YUUgQQnhuk5OCOEqj20
XVSfg27OydcS1lKg+tZX4d2TjuAtDwIi1h1MccQ7B5WdHhH/rBlgpunM8m6HQWhf
zfSO4lVF52PwvOzkwgcdljUMyIi12zBkMmxVRN1Svm49qQ98vmSq3V7u11sL+WNv
CKtKehIOQxE5uws2XSaQ7YWawl8dl2gti64JUxUNpHNIUOTMYZpk7p2LW1qMAx3D
u7IYyViud0FeBwuFPzj+jW4CfhcVKbOy4s2apUi8nHmqB/rOEbLLIJ9hBmD/q3vX
FC5ExxzBTAt1l6Q2vGESZEzWMW79xpSeHWW31ot4duW/ZgOgVjtZUz31Y1EZhPnN
AQZ7sbr0A7HtPp0fN49KlEGduS8qzZLGlrYEa/OqpD8NivaeAc2eI2tjBkDSrqn0
Ty3+DQciMDCScGx2E6e0gELno3G5JjjimV7eqEUGCEVnLcELE+bgMaPE35tt3rBn
pHnhiRzb0vOW7pPFCDdfGQFww8OdF5edxGVOBybDc4MgBri+hVOlxkWVBQdp15KI
uEBPzHEQUXcWW6QGhn2qjf8bDoMtiPu45p6hKTHmhy2Kjf8gB23rJqNMZXBzxvi0
hAa4fCsgN0p67tiSZh3cwC+RvGy+Ss0sZsTqFUv9neEnhRikaiwqJSRp+IgUQNlL
JFse4y2LgYTeVvv6s+57R+ed3Rh58xNdvYLXSRmkyGnvWY8eVXXbWKtNB2Wn3CmJ
7704lnBDba5yap8Abjfk3dxT27lp+cDEVOdQUFo/+/3PRla6Ye9ikcTQX1xcI47A
+AE65yBkyNtFNnsClNYWJ4d71V8qmdl6np0dYyyjEuqnCmjqX7xodjbEZH0ysXoW
jYiAfutwMQPdh6QFKydDMTNdiX34yjRedrXeRd84t0ONpVtBAOZj2AANzgOViLxp
QAxBVBVtR/iEO7g3ndbh6B2HbISgr3F7ahSu1Tq4QyPCiV0Bnyxw+PRQSbCgUzwk
mUkTWxqa7gi9+X6ubm6HdKWwEdyr1X82p2f7WB6DZMg3mY+tzS1dX+2R8ZOIgs6e
ghhAwPz8mVHgCmrkxwkKCBPtNg1bhFWfvKEVYyOpoCg237Wu2a6lEhIdGN6q82pc
Xu5YJGkHW/H67RyGoecKIEiOIDJJRo//8m8MTSPf8OfjU66goMWBHqIpSotTDfJM
2eZhI5bHTf8WrMHzGxua9kiYLSo4tSob5+lEJx7L7gLwiRH9qwUWfDKnFacJpwGo
AnqMyIpiGh1xOXKQ4i7QTaF56BygXvgSSM6igcosCcJyHaboGgQTmRECxwoORZ6A
gLozlkEq1nzAbAH+Bio3K8thcbWUqEao/9PdV2ijGJqfytwkzw2oT976aTQiRw/M
sj1ArynJb8W60C9Y+eepwmEmJ0ObGe5OuS3YHSJbMkEe38TgWCgJ+E5jwN22Xk+7
M6AUS3kkLpujSW4jCyXnYvfk+TbnsLMyV68satDgsofZfUISri8QpNaz+1cwOd1m
TwSaGpl7Iz6Dg1CvXFS2xxOBkRpXqnFiTr1oNswX527hw3PTNohwHNvJX0HIJltO
0rLQnlO3725tHaFlNzZ3C5SeWuqopQRL5wFhKv7ZrZS9OwuACVlZz0FPDt9mji8g
0+y+KZRbez+jnrXHzRDZtt6P4lijlrbGfg8aJCj2WbF946GuyWvH0osAOO5zXLbF
/yiCA2BwMoBZ9/6lR0YbVYnWsfPHPiC+D/Fz6peZ6kQyOpw/zDEbwQXmtgAjlSs+
DX2OiGX+apx0OB6CQhSM76lUc8M9S3rj1KKv8U9QL7ZqHE7CQM6kZmQ9+7Rw4ofZ
thYI5j76vKM41oHMDRNe1SW2/9zLtLizKqzq/mH/VYiZENtlne5R64tufhg8GT7S
FXf3zaNlddbREqHHT1S5UJ/4Yhf1WY+k/aLJiyy0hsoDi7b7DZooMjcJvuMtLwZn
a1+RK6Yb25jRgHO60aHyyW09OhSGH8awwUnFqM34YRQFwfDi936bI7kk1tNjZgr/
sxb7jLFlhM8jC+aV7k+XiLp76uiqjpeQRCUBC7NSjBMqKnxjQv2ZWW2IK/goUgWq
2cOmNxggHOODudJoZNbH2jWYNThv6GEYsephzodrJTHlofO66AADUyej4QEiqG2u
zzIFPOYHFkc62DvzghrdY05V7kXYBOJrZPYkgYUsu8D4qmnumrRz1ypXzQ2/IXqX
kdOmQe172KMGm1UzugWGfQNTMO7fY+wfp5bavKDqf+I1VyX27z2tCdJSr6U19rCc
J/f7OmwDBTaaLGyRIjXZng78S4oRzVird0zuE5UC/mQfaNDhINi4/Q3naw5P4FUQ
vduN6cfOaGxrKbl8ELlAmDjVKg+MlsIrtg3xzdGlK6mzbrwejsPHc6dNugrHC2FK
kS/gKkyNDdudywNM6TlB7JfK0z+4NlIZsTKTLXXlsOa8WHDFoH1Rhsf2TyxsY81m
2B/gtwvf/AUq5mmP/P89cuX/KUT8wKwOvaH7GKckK5k+dKwC/LlhI1Sy+t+Wk6kg
Y855aBZUB/XFmNenB4w7tdSg7/9KwqZ/22EKjDDm7sz22wEWgRura9dbcdNDp1x4
Czmcyr89RxOVpgHfD8mJFp76+d6yB7EaARi/lqgWCe5hbeOCLtHXpxSmRtklxG/R
DwsD+WmSF0uMNWsBCif0pvNC6BvfH9PHveR6y80Jth91GK4BKsnhdOf1aEiGyAhu
FCd3zFVA4j/3ALpC1DQf1kyFlVTLq+ny1FMKUR69TbIU2CL9e9Izm1R1Kq/w2O46
qGABN8yYa2JBVQ1HaZHdf93VlE+dLcos+8YFPmEavhCsCBPtyzsYm7mkHl2Jm74S
Us47M0N9KoAcXfq6+Prhfqym5THbVP6m6tDz+n/Zy0ZfYJkzakRanR4ne0drZrJO
6xTf2SbBg2CnTOXzZk6l/sVeDyYKvot4alBWkYYJDC/SyIRXmOCfXWKCLc8t5xMJ
HpRkuNDK3ksw7zq9F+Sg7U87Rk3piIYFfGRMz9qA1nIQGhb6ja6/kilxReAJvVHo
uZNHO7JeLFYSB8rMP7SmmhZFPfNkYO1Oc0jPJWRlyxGUq8HLpWhZviBQwF7VaB2x
FAab8ymSSKLmZ+yiMOvVU5AFDHWSFkKOA68WokUQD936myhVVCeL35flQlTHsvnW
u4H1YO8xdcZcYjHcBBl1zjl4eHjEI4aZ6Sva5NhFP1LdLIKWo1SITHucf9DVaiRv
5CawYWYwcooApahx4XHBGCURj/QO02MdZ9Cb/4ZDs665naF3w+jvp7QW9zsu3v/v
AFDjIwm2PGGX58udbFt7WLcKVQB8I6v6CnbpBpWgu8+szS6+jaMocK0g4Aej0klW
HM/u5ksAL3Bjz3OhdSdwQZHHWfYaUWpJLEnrMtCcI8QZo3q9usFQOAiWTrfYyBAT
ZaAsMHRpVbJYaFM9bYW55pcfgYQ2NQtWG/SiApqjAr7iZMXCrSGQgAMOXlJg0h8K
8C2tBTs4j/AKlj8hxG7CRwYbipTddbhlAn8GdNRUBVIySvmdH+IjihkBVcySXzb3
+isnvedGt8g+YamNhwKxz6BSroc/g7DuC1GXG9EHEsWcxndbvjKSTkYp43aZukSg
72J4/i1QBuvrLAD3O5L93jIATFfnmLa4zS8actgZcc3B+3ynR8Vmrb18y9mIpIyU
rfQaHiOyW8DcMx3Ygf+vJZSJmBYE2nI/i7o6gOFaKYetMxfb0yTCoam9f1B9ZJ7H
RFewP1NKS4VHCUhDiwc/6ig4zQ8zIc45cv7GxA4z/SBK58dG4oPOTOMacGeRKNjE
epnlqA1z+wM9Crali/ngolIv0pjMoocPW/t7c4KaEPnABIpzYqd5shYZpqCBxfbP
48EL0Tk5dfagEIdLMEKuv1w9wQd5dfyfHlt89C6DTkWDyHgl5DLJE2Cg1Pjj5Bw4
1pqNVE4ws6j51WZdxb0Im2cDzqgwEb2om8/wR9XnttCbblrEtde00uCcgznH7Cuz
itB9Z3g65TXPWrqhO/8WBUOzqQaxDBgb1TGtjU9uD7/pu8QxYLiXYlwxZeRbl9cb
euOfg1ZC2OV4vp1hBtKKF6m9PT/hQJcfP4pMf2v0yJ5vee6cD3icaHy5LBr+EPuU
ZjOKJXnwxFSbAPsb62V5liB/BDyHG57h6+HGTIGY7vPkuXQa13R+G8+0Iduk1kJA
+epdrIiRkb+/BW36unTyJ62Vr/fX7OUGToG1NeHaOIHof4stwWtHPwQiHG599OLH
Cix2pfkbWsi4vJclfJNzJsgcY4zTjVOXsaKbuy34rCBhw8yAWrLZ+mGPnlfgQRgX
MABH3FYWHdQrXdaoEh21+UwAU9vkhA7D2sh9rFEK7vIu1l934yO8FqaqXIPMdmuu
BEYnEAcub1t3vrqLYaDK2OSSZpPU7WhR0TON6zFd9Qw5qJVABy6Yele81cG1AyPJ
IQqGeV8thqzcj37zY7YQt0dbgVvTMAWIG7f/xovHvA14aiA+60e+YJckvuYKwuHv
uOKaqwhkoUEOXvcbK62VMOKruNTZcaubVzmbQpvk1rQ7nHjni0KZKedy2Lr27Wgd
hBb/Ttz3EEoC6zNi0VWN2k/00q6aaZCY1Uo88FrrcmM2RZkW5ve3QtQxuDsGr6Qr
WaGAN0OISojj6wtjWR8yVFUhPEyCut03+uGocDaMuDp6yLTll3RpmL1TSxa1Dva2
e5cpUlu1JEbtq8J/k+jICCBWQ8qj6wwS0RDqVMLGlcnwyQ9t2R+CeMrCo5Js91Hj
6b1hNKmJ6llP+O3qF9AmkOGt6PYBj8V9A9QeWhnpv5+1BEKLd/OzmD6CwiTgtuqt
X7IbqOsFodELHhW9eqTn9+73C8bXclNlKgcPwWS79Tey7/Y5x6oHmt2mSPn0CLgM
uzyK+Y+T6R1HuypL8Jb9tmcGK1YJF7QcAKDoiHx5JZx16sKvkQcUF2LuTfb6HIHT
UNrFlQQD8B35252kNcK2bkrEdeUQw8IlvMARuBNKRvwO0uR3VHbt0w4qzV3Xu+Fw
8XvGmVtalQHGnYK3E33yW6KWMka0tkYrsK4TBnbkqzhy7eL9s49ey+E2DjRbYbHW
6VKn9J6I7REl81m2omuZKcEQOANQ8CEGHLKuADNwt1xHINiwAZaivtyrf5GD4Dpe
JF8+RGGXH60u+VQCf/7E3Ffe5jmrdmJHm3jyo6dAlSjK/fG71RPbPuqio1XM/wdB
vWfX79OTBQ/bquttVUutn4JhMcBWlTQO1Onwk6tzF2rp48qWqLy6qUOT1i0rWp5A
QbAQbV9mASh9F+EnPfA2kRWYYGPsVYVgg9R4hNbC9jb1emue2dXgKvOrvAO4SoQ6
s/SrC6PkOO0+VGmb6j6PwruHEQ40hfZ7wUrOKdID1nI2t8hLX8npILcQ7D2apY53
GdmH7h1o1fKmRN5Vkge6Ym9Df6qdqfZJRBCGTCa18I9edD9OgZDq/zVg87t2xe14
eeEcn74RU2WgwNT53nmfE7k/MkgwU2yvFBRlFLbDQP32QtMAtphCiS0k9AdeLB4C
i/nlwsiZKK9T3q/4Rx4H+yFvC0umzMl5VoTH5LifdDoOIlxe48aQJA2w3hgt3Z0w
JgeA0EbfBBeWIsxE2wQ72TFxWOZu0D5w4PpYnRuO3mput1aNIhk3oumUaVgVMZd7
p0efemj/R1qdZMdEXZrfs3WkQ8XXfv7TU9pVpEVymBoUPST4HkqxAiihigojWDaw
9VJ3UBFiVg8SRvKxEsU68TCwf+4LCS6rDi4eTmyvi0Kb0SJ2TiVGPhcauq88GIHQ
wrK5cP2PCnIkGFQjfebat6HotOYt3FWNI/ka7BmS3PxbK8QKgQijP++2hH+hVp4A
Xu9Yc9ahHl87j3Lzto6o3WLVwaxGjgzkqZ/1srX/m5/NOEZWukOGVYQw4Unj6u1R
qCx1xR/+Ct/d1GQc7vQ9R3WSk15t86lTrsT7izF4dSYQ6e6G2+cLZlUuga5x6dqt
FIq1m2q3dSXbcj72w9PFDWOMASke5h2q1+oJAXRG3eSEm8BZCICkizBCHVUHSphg
JrkQIOrtZjdkNn2vXHJPjm2rHIdxn/fpWL11RFXj+R1/pyVxkPWaQ0ndn3/jwx2j
ie7f6Qx48pbk8O7ixiizQg2y3xLWQz/eXGD64krqu01qUgOxoLrDEIyucaCKh+7u
MUxVumuVsuwHVXdmsqJ4FtOlLJzEKfJGcq3FnzRo+S0zEHgbu4iXRpe1HN7iA+j/
9KGdW6BbUd7XqNqvrT9BfVcET/8BRbj4resO+3o75PFHjMKMRSxHwO2IVuOpFx+j
2Wazag0uLCUwwWi1lR6c+YeuS4moDAvu28aSdszPojwSLh3dKUiF5fm38+9+PuR1
0p1/jgHozScy2zAFxn+MJ0/+UCQRvr2WkzdnZ0NHzfGoVXWJ+49F2CbDywarJSNi
4HrNP89AyXrxi1VMz5ZO4fGQhs7Jt6ZEd2E/6Pl0BLPkbCT/s7UbCJeMJ/ZUC0Ar
9/QqXgRaBJ3Bmevl6h2A6LU8nSBecc5i8IdGNyf+fxpbM156TwNSKgZQOKd19+o3
MYqXrvsRYf1CwKNYe/OYLskZuWCYtKyh1FVPHOymOSc7f6Q4Os98R5X8m81loRlR
8b5KivE1h0ICND/x3G23OpaSVFoNrPSx0U0G1qbTo+6i7K7JCwU00n1mzXizqhEw
sRdq4kJwCYilEidVZUNQ2mtfuKG8zm61NgAGtuOdG3jYdSqksTpfH6hYczJSjaB9
0wghbxoqAe9OjBB8qCE/ceIwXkp9Jp7BAgIyvAIQLSDyD4YJ25PBjAVikbKYy+UB
P8lChftCxg/7ZTE4aUnFZsSdq+WWXh32HLw0DiH9WSkodEdm9qqmdL3fYnLcSzVr
hjqOzQJVZYDdZVgO13dFcvy9P2lBA5F2QEb5EJjHdBh0x3L76W/ZpSLbGnW0G6rR
KT4YU47UvCnq7XX6LG7r+73uGhf+Ud/eYx6YuHhWSEu8Zp7ZimXVrz0QzE6f47HP
1/REVgeUMR2A7xgupGGHtqwmyuqdioNNQ8qYz3EwheBHiyID1ltMewhYP81kEQPW
2bpK36321FRi6tuqVZG+TswzozyWKCDE649vjtxEkx3gnp6qMiTjeQGtkB7AuQOn
cvpS9H636dLHO/nL9qwNGQf2ngZKDE2U0bKq9gwVUwTes992045Npgk9IstveFrK
2ODhRrRJOj8XWRhAJoLYE5cEAzPva4HdQ08dRaYu+RmAUxblw6/FQGwGxTnFnfVj
S0le4/woIf0uD03G054vLiNBpWvimVvI6sZ3+YzZZBEOL1k9QXRdlodDPPU9e9vK
y3cDntIhkayXME5pTTb44yhJcq8LnXnxqmYW+Lzv0J5vIv8W6+jsaCjtZApGTgHC
Z91jFBB2LV8myaNyHJX8MWis7iWqOrSyQq100aRFnDUrn9KrP5jNexOdVBJLSFMX
RgoHbaU86dGYVa9+STOtY/4VV3BW9Q8DaP9uX3fe+2t+wkoSAU7rdwr0kXUqm4it
BKc3OYAxW638XSh+0hwtVJXLYEYCSdxrWrfGINsQ9j+zmHB2rNa3t6WAv2MaYf+Q
7gyZJW+wiNSsib/OOhz/I58v8pJ3h8ostiHBOhtkMpbal60tkAy9SrvtNR+qkO17
+SIj+FFL/Q5V6wZMudUklNUGb69N/KcGY/gZ9ILde2NeaRZ/AN4GY5gETUXWSsxS
jNYeYbwMwGRiOj957DSiyEY1OFTskhwxrs2ddyZe+1/KiEabOe/yqdfwUdfPS0sa
h+ZQvG2J0URcTSDSAoGkkmzgmqK9DhCg3QLFW5PFitACyBeFbjXj87oqXJc50GUW
h1YM6AVwxr7o3iCZH828x2WCa3x/5Xw/ibPlZKqXCJu8cCmK8nKQFY3xxnPJxF8J
1EZB6fQfImO/24HMarc/VPD6D0/B1hB+poA3mzyKfAxRYZGi7SfO9hhvVbL50pug
SgIxBkkGKPKBEs3JlpIPiCCd/jkoyeS/JB5kVwfdPcvRNdWZb2EZjn6NtIAts8EV
zlT+MP5xPqEjQtlLjgPSMLossZ/6s48B3BPWjrTtVxE4BUHFOaEpRAF3Q0TDHxjZ
G9qF1FBfjYlIqjOIwAnnB+kQomWANLAY6sri/paO6bZAt3Pq1SyHeRfrTLG/8+wc
mKt2nFrI/FdcAXqUvengMAWMT0Sy7rgaWBfa0jW0JYq81uMbxbxRz0PGcMPsqKMu
cS9h9cqN0P4vHRLhKejdRwBXUWkTNKkgA3Yt4Poy82zrjRbWffZdaYVAw8QDk39c
UfM8+d8t7e30E4KwlGDsQeiaNBjyD/LD+VvaagWANl+pHpflHo8tJqkZdr+BqR8Z
pB1djRK3qIqa/71PfR1dczqEA2xlSVpLPV9JmSSVjosO6J9QiSaUkxbSF8ykmhaV
E9CxfXhOqVXhWkstgy21DS5bqMpyxCe8aB5p04vrq8PYfw3BcK9wfq5iRHgQEuWi
0pMiDUqEBcHIuaWlCCJsKkT8A2bagPxnfAqTG7fXlxarqvdWx6yFlV07Ox+qSD+D
BnzDB6gUa+G6KY/mmIjlZMXOd2q/CO0PEMFvrU4uc40p7WZGw6s34QDSDJNw/NUu
mFdH7fURHBp6D63DRau3s3/Kmtwou6rT5RmtL7Ei2dT7E2BSHUn3WTG4a0fdKAsS
WpNzCCc4F8ewoinjeE7Uc57dOMDs2fx28/mbEc6XoshA+oaol6c18o5ADuRokT1m
vojsfwmOlvjlPBGDUtcTkpr7SOQ8bR4mbnv2mXkeRa4keQsu4XKrst6F2dQ1OCsm
uOgHbqYFkl6FK2VurcA64eYoqhIkZ4ToMAI+zcLLk9R/1nHsPMkscOJyUEFwclGn
dGD046+lyBVApLt34m4ghtsg/X5uAeucSk5pIUBtQL7v0sg6/8VZGlv/ZhecwxMi
T+yqueMBm4Scg9nI8//aCmORStk6UXTk7Xu54GR9153stWyw9fb22/aTI3KTopFq
oz5T/NHsyrb5TCgbKaZZwGKV+vq1g0fGxB2tbPsatByw00oyGzATgVnwpUe7tbJs
QAZ0vN7o+kNb7JTwXPbIPvmdrneNRwGAr1SV7izSOVfFBLqySY2G1c/yp+tPcj9K
2JbaGPM11+uSoNrlLeDTGlSrX4n5KSTVJokbJOe9dAavtj5F3r4ELsFTiVJktA1m
xrg0vbLmVMv8q8KdJj2WOn7UhYJfLPj2BgLp1Fnrwp+09efCjLnj0Fm0BWZ+re3k
A18gP633bm9A76RjJ7ugh+excJhhVbuIS0wIem7amdV2ebEm8BjNd2XX9tIqEJT1
RdXPPN8BaHYRuOB2NQ8iTdxQgztrtNe0FlHhiyCndq0Ri8PzmQKVQSbrqNWIVrAh
yc8+5A0+vp3qkST8bgrO0ZKhZY+5r/8zp/Vg/hKYrVtz2r6XYy+HaKne1z2S2+2D
VZdKAXpdQY2YWFcDKZoQuMqEekJ7SeXGLNRsdIR1iirobOL5oKUsCOz+5Sp+Nx0t
IqTHVifVq0/dTp0fiEW5OfpiyuEIBBfuvQzOvIq3qDrnTNr4AEKexRo2iBEjQceY
U+df0pMYq54IPrijE7MuCvbuuq5hGzsu1OHJ2POfTCl0Y53IQdR86cQec8WqHDPc
qIS9D18qorrCS+OSj/7dmtt+Ptm3olrcW6qfYc6Dnty29UU1pxW08eV1AjN/RDWY
8aX3qgCdJ/0+Ys28KEniHabm9VI88P9U3tMcvjwf4ykMV50DR+vC8H8MfA7grl1H
jFoTJ1OkUUi1zESuMm+c8NxEhJj3FVwvVemGTyKPSPwsBxXqVhaUEiCfPtWv9qYS
7MmwTDlSXuSFm6kM+XVlF3TxouYcgZDO9kP1JZ03Nc4TTU0geAa0CuyUth6HqxGq
TQxiW3IvsnNSow5XoJAEkRe87pbhHS6wv+OgRxRoFd5JfMaKmYD09JSKtYzyloc2
EtAS1jNYrIl698F0SZbK/QLm0ki6vBvb4ED+AFNQqNA/08rBtkSM8tXv30CYbPX7
zXY+1j4SN5TpiTz9TTTN17Q7Yd3FXo9OQqUQS5gZfa+mlw8HXS6dPcixLmCDl7KL
GJ6Rl4wIBOuwU9jPJX29Jazt2EW8a4H7885p/jswtlUbS7F4hHNPWY/oKHkDY8AF
H6YKiI22Uvxs93vHVcTRakAgD3sOGUiohnlUu1LDHhhhdmeJMiwp83uWGD7NGY4M
bLx76WQSzhNaOQ39eYLzzQbLu3P1jfIxYiMVE8XhyARHpKIHnCL/1NL71Nq16MjR
/jwo6IqCeqPOI1SmiJFsgYwhQJV4iPOJwVFRLOdap5L2GuRgPWDQWEl/PUvkkk/N
90PpYk9w02QtMUl3INBcxKSVa78bZiD3hiLZpM8ANqW5VFxp53szCcIFaKXW1WXr
CdWjHxigiEby2PpGUoZ6ahcacshxOJ/bBKZTlOCZyUqzuIQPZtEbYv0DprRMlG2w
B/AiTtaq4H8OfkpHxJSZQc/al6V/tQioK7HYzBPr47+bkcWCVlHgjxnVDM1+BZHJ
6qu2sqn29xtLbaxPEg2ENsPW464LfSy0CnZn0wcz8CRkY8aLyff/KCWCafbN71E2
L+1ooLtuOED3brJ7pza9rjl9hw8gZ9GoiQzhM1hflAUrvJ1T2p6d0uLqLFP0VR4k
14et5ktNg+h5HEaiwq1SpE0oLNMuC9stobQEJL9O/qof115N4AcFTRqZGCgCsYWU
nmJilvvA8JONg6EZfig2o04yVy/ICVwTCfLSSejSM1WSSQU4SF59S3/LDQ/UWtKy
LBM9YkY4rRuKICYlOUOy9WjLZkOjQ9CPdXFsUqBOoM13jA2Y7OH9TEhMUc7sAY9M
44gO/c3um0biFinrQ/rbcV0u8mMXdJ1LEwIoeErv6KaTiMhHQS+G4SBI1JrgD3ro
hPKs8GNzPjEekIm37NA8lggfjKIpXkTxkc8aA4oHm7PYg8C1bcmo1E//NRIjU846
U0cP5sWaov1jth95gkZqc8oBIQ+1rR6dH5kZBD257vnxUagc1gd16+k1dmUKkkfu
Yu1kL9cddzrGWHz1m1XJM1cwO456xO8iZEJvE8ALowr4Qks+5ALc9JTLrT4qJxti
JON5AFGLNuVTwbEKzC0iQt66TjbH4I4mxVCj5kBw+kBamHPXNCwYEvCTqMbS9UaR
/RprEtJvcBosHen4jTXRGO7P+aj6BwTEUMkaRN2kPlFn8+esSeabJVWoWJfexsh6
k4MSL/98JNe/eyM6CiYGoOyUerROvyuGhXufKCzfUVeOojdUFwktlYh6tY1Rx+V5
CxoOlgNKh2yQycG1uiUY6AxEjr4hzsFDjlW7cslSofXZd9ReINZE95wEBmMxOWz3
OXWdNYigYSqudzaYkwVTFmbbYWjhB4+nKbqSkk52fy1J91k3kvh+NNid3cUPxIKH
iSVMM9aTtcerrFXJrD8iKaqrmfOJW7Ixej8xNzF6/BSf7BsOFnH3APIcTOwwK3iF
9iztCiTaNexGVkGEt5mOuHDNW79wS8Nh6mAP/34ekdv2/uzUarhQlUCOea/LooXm
1IufmbphakbEcqz2YUFN9tfL5cVh7cL/qX9oR313xMFVEEoCW047YAqMSfGMeuDz
od9JEi9K7CLNxY9IjapT3mXYh7VMWCW6vud1PwzgpEu4x4A9nYzz0/1xwdJLDpES
S+YLErtf7ScMGqn8Useov3mwFyk0DJOWGTNuSCXgifDwU4pFq/jRQwX1T5Vmz3P2
+v6Lix/28iX8cR9nrvovZPRo2f1zNvAytkRFYFc47M0FyaG509sLuqxbNYNxsKMr
VbrQZwTZn0fBISgGaesfz8mD+lcLtZVEIsiS+D0bIx2l+DCOKMo2zwUYcTmRGTVk
5jCv9y40Nko6UFYwm+uev8DX4QSDJxgycv4dLdHK4Cpv7qIs8pDr71KcU1Ir1GkO
4c9lpuTjqMO4UKvEByXVt34mjlJIF2HTJa4F1X/d8RHRPSPKEt7W7QhLlax54HpU
2ekMXVxiHFLL5ZaHv4lXzJ+Bl/9GaD0TwO5zfPqKixdh6HOU5DjkmKiCVA8PtjKr
A05+8osHDgDmQ65ZZj6lwJ/1UmSeCx8oPLpb7cLOHnnTIDCYCKaGZslMyeY8fDUU
TQpxC1USzabrDmQPpFPonupySVySuLmKntq3F78imDk/ilB2YpwP1CjyE2CKRMOR
DRFjNCm3yGxdgjirI0rRxV3ruHg2LSfDYCJiXCqVz+M+BAVRN35+Vf3OVt4f1MXA
M73ePUTQJy/EIjLH7GK779p/Wxli6SAJdLnwnH2J2b1nJEHrGsIwqP4Q67BUmqf6
b3S1qT2tdODvhEwnxgx8od6nlVv/uauDbXBSlHjX88kWu9BqNqwLWpvN7rvVme+1
MtW1kLRbatRA+xS9M7IrjqhZvtD15dX4ngDTviic6lN4v4WwqKaZgJEX9kcjloJD
xayHwOIbFKJSp8vLqQhuyInBaF4k40HRfxJwMKOeDH6yo/TXAHicJg3Du1Gh3wF2
f9yzlKnC4jKxBGQw6Wu6nyj6/Ozvcyr9XhNcOPuDVTkUrCUUy6fyiYb5ZNm8CfwB
4WqNiPXsRn3TxWlZEPEX5YLOMHQVWfvpyR2AfIWYlRGtebAM5Z9cJ+IZqWJwhy5Q
HP75F4nf4gfbkGXZboqYViu96pvX1E1vzLH8Sxr7/qFp2uPnEyoIerXaiP874Uot
nDM8mwufqFC4JvGOeW2p1HOdmhSu9WK/zkImbCZ173ExreiL97hZ3yPilKTys7NR
+p4Lcms5DSrXlg+yQLACUK91z1ls3kEB/pan4U74E0jqzXRS69aj6IOJ6GhgiBf3
i8aS/0fLTCygzkz1UqeNly5FGcHgE8lhDBQb2vc4dIzDAm9H1+2CXPp93uwCVXur
6tbWe8gd0YokGThj/vY3A5UCCix1oQ9FqjwDfn/xDL/860/3hdbcKm5p7kbhLUtU
pmB4Y2SqKZ9XP9D3Q0TfpozZdBRkzcvGa0OebG9SPDSGIgLQwSup0L9phzOwDJBn
35ygV2alsbSanemBxUlGmZC4+tyzo3yVhcLTFo98IzPkAwoI6qfN2rwfIc0muMOn
86lV+l3Np1IbGoRB3B5bQKVKGEM90plbDysMzWnS/tJ9vLA2o8SOgYjBb2FmryeB
yUCjWVbV8E7muIblAA3t+N4cS0QAQAf72x4fSNM64OwqfnOFYEFH39i7CyqOY/bY
85GLnno+hIJojuFsImUXP8o6NTnEWHsSMSypNnQtnFyatEQOIXAWE+thmQpKBGVO
cyqeLIOp9QwXARsAYx4Q6ozXT9Ph2jkEnVjtDkllcDpPUfcZ45h9kmQe7n34SvqL
rRY4dO5xswdjCwhTq81qNHJZ3VwLlEv1jsIMNzlDt15YoX5wCdw684op20ddvtxx
OeGlxCjvKnLrYEk0iTm13hqmT9w+6q9WAGQC/GkX90WDkwFKu4GWEQQavrHv6MKv
L99hXHy3o1/mqXqSvOWrCpv7CQjRrU+fNLwa5ySX0p04OsLYbzlxQKk82jZjBU+W
5r1eMYiTuBGnN6iNqLasN2nfkTZWUzGVJPCHNloI6Ny6Jyz+8SAP7qC6AXElzxY/
8AIq5lg6pbbE3JEkcNMuW95NcS8tvAJolHDlNTi94zN513FLMD//hpNno+bzVGo3
rDRQ/1IY/1jO37u/SALurWIFpl2GETlu9rL65g2EDKl+928FddRsHQ2kooM+qwMO
BHwKs5uhVRtKUiZO0vrclTDRiGccNZYsyKobvP3XIrgdehclWmkoMXfjRzoLWW7e
oL0MAvDIVrk3pVuqbyawUUKWtMi4uP4Vso50cG9MAaFJDKgEzHFrtsLlX3FKSEVT
kkpRcMGhsvkRE4cXR0ru1VA/xIwy9XrUHqVZGLmrBl9tS6phIql9MG1m9VVMVSSm
1Y3/I4CEU30ExGsH42KJ0xopSaXddlsbGxn/AtljrhJnMENcq11fb22qSB38Oq9K
WybN7CE8n5Jq5+H/umKz8iGQ8KoR7aouGQAcaIlFYeOfpyDVV5hX/JAS0Z4OojcN
d0nKhZo1yDM7sEgIaVeaLnAyjoqOiJnSXXYBr4xZ/tJtzIbgsivbsiA5HkY1y0ov
vj+2hv6n/5+F/Ub3EklFPjR1TJLlf4Sjt8aKS9DCVXDpt9N9HJ2eLuIIk5qk69cZ
zc/ThfwiC0S7sE8AEBXpt62nYZn8ym5jGOUJhx5qG1Z8Y9tFjChF7sjPPi7Xos3y
k14RCHPBWKZj2ny/Gado8d/wXomYufaJxO1xlYuUb2sRVU80mfbLtd1fuEVaxtHo
+xk0RAzsVmAs2UAhFv2nP4zA+DU+F7iqnhvDLAK+YipqcWV9NY3+xSp0i9zEhZMm
EY8XmuYVv2iNbM9jtqsj/hu8ulAJDGjF83H2YcmoPt0MoPo/6UcPouHqtLMhqxIL
O9wi/8H3H3mxTqJqQhL7rQcH0hYL/B3upLqTFBKtpTYM52zLhL73ahDrRaRkFGyG
xoSCVMTbGHlf/nLgZ5V1jtNCRyZSCQ8T9yYcUJ3gfzEl3KFyeSCCQK2/HlgosGjy
rPhex45myxar8yBYxhZ7nZ5LFeIFgVdsaIPARAb0OVspUW0vvPwMB6yNNUzGanE8
lOvcdVLyejXqXISUE+PwjSDT0xMnFFfD0xVVnrQmYTohq2BlB4ctJv53EREjImTI
AHe92WCnm94+QmsPyXMg9MzQBW040+oaZ92f7E3v/K1Ud8P9fLv5MtDb1FO1pdvt
QvIGsNV16z1JbR1/AkuCN99PpRyl9hpO6bSgSLK0Rs+72BmTpqqFD02SPMtnuL72
0DupkLQ2KlcS7ld6HHikhVpvYHjmmyxOAwEiX2w5Jbmu51lkzSes/hbIwWD17Hnv
9Jnc3NALgB/iZTpVP1Vwar+ibsxMqK91FOAY61xBm4pHDiDoGsbaq5DhjvRnpOpO
lwT8L/NZT/pmwwbr/m3fzwNfw2/90w4Tls2mlT8/48bwcMakVrsCcW4MAJ+38ONo
VxSmuxkb0bwLu48K2dXol2lt8PQ+rHTAvKR8iSuMX2ovcPjsaq6QZR6uDzgskELH
vMW1/5aBB1oe7l1LA1UL5v2V12Jm+BE3ijfoJtefvRJRLN9pefVuiSS9D0KWl0qQ
rF6huhmqqGyG9nCFLHk2pb7q2JyV/V+wyLzLnuywTiMiYCj0zfOMmaWZWu7K3jGF
FihabuXDgPAXINRdM7l91zm3J7XfHENLmSSrST7EguOy8wMuXx6mzBpjtdpo4kGe
QOjiP7uIt+ZbfFdZC+P9aVVvxp1a5pyUDSInU6Tr6hauoHwOMQMMZcMrMNzXHj5w
OR7n8TS/PZKktP0X82vAMJiciMCUd2pmCTzhY6vncokCYXRW0NRUnjfb0RAnFeKy
09+zZ67znx7m/A/EjchHi1uPt/gpwfYw62mkFuPvnDr5yYOxelaeVk/OlNDEoIgN
F/kT7CORcvODuYYILpp0BqjwkDOztRRmnth/uw4t26vYpPLw5htP502iH+4a4Rbw
3JZr8HhiaB7K7s+ZHL8Dwrw2d2O6nSbSqk9j0vxOqBT2Ox64bFylN6K1iIOR+xd6
ezKXfrphwkmFJwzJQxXgFyJJ32A6msYPCsUFr8EEYUBj+RswxLBFcblJytHuVc/h
AaCC0OgOtm3SJ++9paeT/RCvF/zcGa0aP99assx8GujOBopJwRHGQXtdQnbyv+2m
mh22rkJMOTEZm2GpXInEf84U6EzUoR07+mtvvTkIo2RI10OVEQ+jwYsBqax+YgnC
C0uaFQp/PpEbx5rr3mgDEz3RBNRV7W5GTrOYvPu+p0pcMrMt7TM9RIbyclBCMMTm
1ACX55H4T8oLoYxnuqjADmerHfXzAqlyZhJ4o9DQSQ9Uss1bSw+hWw9nTj4jic03
2SAKDtofu+6PbSirFY4/Z0R2q7ERveT3GBEh17xiVBHfVCf9ZzVQ+fJonoxPAj9y
ir9tqdW0QUcMvPvj9Hj6nb4Cc7acyIGlPzLi+UAKTMFXCgtMWUUg/l7nJQvTgHJ0
2aNowUDQLfEBeWTYMp6VyaIUq23Aje9XYSOE/ue2IITb041CDgd1KHk45NTMApq/
Z41Ix9Rs6pWrNEI0dojQmPzU66IF9+DpQmP5tmR1IFh9EAy/tylyl3DwmTLTULsm
ShpqwqJ8qW4zrOUI37bdyV1z8UCrZXIpfAbqQ5WuftDwO/yPLo8QgXLHdJXiZnUs
sIeZ0o/5MNCz6LM3lmc+eg71+b8v1upv601Ulx3T6sP/4GbBIPjPPUb5HkumaVEr
eKRzP7kPByYy6abXuwozeBCiCQviAgEuaca1ws3XbUisXXQEs5BXQxxiIxmiLxe1
irMyQuo0JTm1o9OjwdxN+wvoo21dMR8x0Z9IMRugsxhGvKW0BQT0L15agsBoZ9C2
QwxVCFPqpQYb25wshtbu8Xlsm+vx+dfi8RZbdTDBzhOMXsL91LeQpH5VQkJX3UX6
6ee8ldyFjRhyKXAFyja2rzd6yHq62iqzQLlaLK+mZBeePO8HI/oqacmURlb4px/x
QLbe2d+Hxn9VsO5NOkIyuF6haxQIrEEsvWs6t8CBhwpBbvO0IWsKyWFlOgutxrPi
x0Ym4TFXNFVHdiqpBD55H6tVxBNg8Uee1xiqiXHiIfp6VgkSMSV+SIpgjW3O1DD1
NHZyTNYY1pCvtSp45AueQwoSajBEoReoboExhZv44UFIiDnroMGFzjvXgQRyv2up
ntS17VaseGIUgKWpiQ27l6GhCuyuSIUf9DbwhPjC+JfPDedUm4PrQYBb6soZJM8v
PhCB4xAQAwB6rZXo2Vv+VBq14to3H39JiglTBeR8xDzY9Ark0cxxlzSO4LBmv5wU
aRf2y4WP/p+6hqltBPTNgdNFOSRLwXvp2Sj1HKKbbzVcKnHMdM+AqB7zGb0dJcDF
YoCW3q35od4PZo6yz7L2NGDVTPQGeEmmIH2J917UxRNqOAn0jqT+aQz49dPZOB+t
GZlMUkQxm+LXy1B5FevTXdv2+sTwk+RRXdLWsZlk9zcMfqROw8k2P1jARgI20GTo
oMreeGpaykJqHpuDGt6HPmNy0LpTcsY8KumYmiovG7TuWref5VLP5ELJ5KKSW3yh
Inh2nfop0EJD7qR0Rh1CiwS8Dbjx/oyqXCqr+jban+2lrRCH9FdSwEi2yyQseWSS
mkqGuHZxqs1AM3nqH0mp6q72v1pWL+l7OKyPdqcBEK0yPC6Br142Aiw2D3cdbAfH
sTJ4SDjJlrrzLcmFEOwsDCV/yZWWZ3ZbeZ1nhPxCy/5/6w3HroLhCQClrRu9NGSU
upcUANt1sRaZderpsdSQDeYgtlDzFSiajVch/xiGDpUc3D4iwducdFbK1C5M6XDl
aLyFlGzcJP5JHxnivrzKqej0K+lVFtSkuU2Tx9EVW+rfjFUrx9ezsAlT6Cb+L8/7
leYUDAFxocxSJzyJ70X6yNW3y8xCQWMOcQe8kCFiwIwpV8B/mZvHgVabj3B/U7ld
G2QiRCSDbkGZYrtpxclt28QfMqwK3P3mPxs7T5MEzbrZl1H1TJwJZ9512LIdlkwK
eiqR7vJaz9nHK7r85gmaYjaopJwF2pq6OsgvWzMiKuzlhdBl0SUmnUUTD/OU75uJ
G8WCxWvo/RlXr2qMODtzs9nXZZs58iCdrl25Wq4+/7wS9V8FtBOXI3JujkvdSgLa
oLpwpQLwb1XnxTTGTm4QSBRHBbOEhuXP9IpSG/Co69DXtAJvtCRO4dSDPjY5Ha2o
VaR/I48m4mulQ3lGHuzEliAhoiWbz7iucn8CMyz/Lhze1ebki9xGebrKl8j/awGZ
Pp9YTA/PSc0iHZ4phvQDBU6Z0BRFVdoU4yOcnBa/V2rXGVlcZS8IHNdQTRKnnLkv
7m0dfgGfQlqExyOOJLbBZky9tyHgWClqyoYoEDqfd1/UIbUUsY+TuRx2asm5ZvKB
8gvrhh/2zuBEZ5C0tDIVz0YxhiI3vbWsSaCz0/gHb+Mmo7w7Rw7jHzzUoMc/kJlk
qyix1cOUmNzXl8ct8zgdcp5XHM2KKtmVFlWma7nfwjFDSZxmR8NgU6ENQhAIC+NM
vHGeAbXBMZEwWjSHYUATpCQAYkpakoJWDOgy20XX+iqjf+l04pDBvHmwONxoNrXw
Voik239OtrZMWrtrg+vud3VjV3EpKv7vVpAvltowCdJTmpIP/tsEleXoQB0Ts12o
2RRclwcFXP0OAnepbwjV0IrpgyHja3ydnveIKTcI/nO91lfJcs2hdjakiBJ3udcj
TR0LlVf2iDJK9KCQYof0jS6PKMT10NwjjtRLHsDyjZowI884wDomf/rvludaL/jh
Hch1CyrFtu0owv78QGBqfMRqKonVSGNhCWJ/p6y6v22oAl2V6iINADjutUxQ4IFP
qW7sygZ81zJg7XI5ilRCfbYf9J89apWAU7VmJn0eP24b1cw47fITuO5CUQ9VUXoK
Sqjt55OS7RofWZt0uaM4P4cQBZCV0HqRAGBiYLPLSbJnUBoRjtdSCRK9e24v/GGC
IH4Le7Hjq4WKrx3xl34KYZxjWbGT+vR4/ybrp4pWrxl+6FVzJXNQZ1N5Ql3dkf42
whVHxH2b56MxEcDZiXloVfCVPahdcFxgfYLhLJBg3TRRK93J0+ZVaVEmOfAYm9Rs
+L5Ugc/vaSor8IfNRFbUqk/tgAL62yArVyj7RAC61qRHYu9Yc+Vysz3wsBi0/8YG
cOpRE1aphjV04YsdvTDzV2rCcDKliKY5zY/82Lmfx/sX//xIBerhWr4bqTI1HtzI
b7rr/e7jRlvoOWob569jqU+jX3HRtbXmQVmWksVWS8FuVvf4XFC36lPs2KkD79Iq
Oo29Yk0YOR+vSzJHl4wCkyjSnf2eqJc6G7SRh9iYQoY4f3+/3PDZo1uL62T8IpxN
WiT9/ku9rvYybwPewxFiVQMi0FrV7oZlWvYsaCYiOy4Qk9Q0Mfm6AmJmP+RzC+RI
aLW7LFxgRBkxwZr3y8i4uRKLHRwjy+9rX4dqjwUfYB9ipt31K2YAH81iva19A+5r
C/6CVX6k2zvkwfxcCWymwVavs+I3RvtAGq21hvxY09w2ISWJfHkNV+evQPP7Z67D
JfuXRk3hQmz5+hFEV4PlbixUXG7QS2Dfvqa8X69ekuZKx1PDDGMkS08D26kmzdKX
zY+LCwlbu/HdEO3/Ebyokaa/GzUGgMMdEo6+I+p9vHEzPmID6ElPDngAV2fSyl0l
03FUMzPgtHLDK+JrbC702Wfhde5wFl2dICDl1QMEACcdcjTanS+/KBEiH78Joi3R
D4HzwbQeKQ8+pqaoNbwpk7ZlzRxAftYUPq2BCaptqd2atfG4hhhVZJD8su0aNm1F
PZwxL9NFGwrQ129SXkF0OOGef/P4siSVBxsg8iSGkZsB8+FGy4Acj1uUliIue4Ws
DIwSN/WwkrxWVt5UaTwvY2WPsqvYYILUSOuL9G7CzTuyQO2MOjhMbOl6rOUX+JZC
xwPmQpDerjTdT2wyMlawq1rUa2V3T+331l/0wMhFF7aeoGEouD2P2fN6CwCQb8ol
MxO/tTFD/eqn54v3RSK50QFkxlm+MjospRzHW3gkEV1QUQF5ylAkSVRp0pin2kCi
X+Se11ZxFDvZUYQYtzhwDZ6XE6TlIXhem8wbis6BpDF2bi2uRiZIAwlzFV/XsQxC
iMiB8UUspPhnA5HCmPtZcdgW5v/RMWe2s56NRF6gGMJsJ+2YGKnZ8/WpBOhAjncO
P/QskSLFwMDNol8cuLMeBPD0Zc4DnEb7+hfAa5AdyJgs8os/ej9QatL66a37y/xA
cQ4N+B1kTxPIIvQiTNGmBH9mI6I261oTgS6udwXKGS8NQd5Mqz6tZJevXL4/GB+J
B+0h4gYiBsNqCsPcbE1BCqH5jGxzEteZk5pPBJsr6O97bgmr27JpPeFo+JtEZ5ur
r2Z4TsmjAFNSJh0ctfVB6h4n4ryKt7Iycr6HBHzV+XS+NUGmTy8tQz4sqKEAMjQV
r8AB5jgFK8Mv16OvKOKzBTqmNX9jkNNK8Q/0q6Y0hOUfNnNvscaAVHJERZw1grd5
y36A3oKhiJJrqFHuHYJirgGWQyseclkyUjSKcPlHzbb2EZpfjiuhWUsVSBI1tMhs
Ha5quntLoQW06Zn9YGKd44gcOcKSaHZXItzwn0Waysn22Y3EmpMRUf8KIG80FzIb
Xidp3xph50bh96Bpw5u1OkxYVVV6MWGXqYItpw6YiWtx0X3kbswUTcyTHqLgs9Uf
QOA8qspJhfE5ySz2EZR2krOygRj40LYWI4mpvg/oaQm4sKczOFvWRqaOe0PdRht/
pIkSXMmuyr6Drdc+q7ox9hSgK26ncjxV6KId30fHcSKR53G+gi+QIcnC//IPMoTX
Y+B4Xj7YNXLV4r57818Bo9fywcPwhwkYFCnV0Tx/fOAklhJalhUNRru2M4KP0sE/
LEkSC1p6hyiDTC7opxcv2Bub0hJIg1TA/vXktSSdUxNXSyODycOabzMlC+jL+dp9
R0cXC/TwUy3B7gHzVr/b9F1Nu3FQ1w5jO+ZvLVvEEvUdIAsj611hcXWhxivGn6gL
7aQXNYtdgQe5/Cqy5/JSReDxXXxgjm/YyufO9xo/u6+Iz47uZ/r/J3/010mumpu4
xKfaqIR3FmR77UAcZRqsXCrZMqHpASUbuHYEq551w2L0JYa6MW+mG4Fj2LXyoy+1
54cmF+we457VsAAV0Sar6fAJPpovkUVnJhH+TKa8CuW/SZRS+6WEFMj3utojmV6j
d1EaL5WQhtPFcUz9zP7HawS9NTiplngBMnA8kMRN8rNCtb8y0B4BsnE/cptY7EFs
CaWf2dEMB+04gXFKk1RzpSZkVR/3EEj82fbdm6altbWT+/4c1KEd4mEadNCy+Ioo
3wpCf4eDnFUDZ4HPJaaHefpk3aCqkoerrab+LP3PusXiEG+fXwH6AUrN1HKdoB2V
fWMWfTpm3zctVDIe75LNVfTesu08ZeWtCHkFDASc9nCaBw6r3wiKlCzy7/ekcQV+
4pSb/cIEnbtGvYzvnCTSmhlZrlmAlLXHu9wY81GdTFRIeE1JrWutr7PUGSYucCeX
pQLeubrjCZYsPxmO6XrSpDPLY7ZAoLy1l13kMPftJEV3cFlSPov9lNPTzLBLV7Ub
bqaVK+bo0mMRDa65DxI/Sme5J9+dgv9pARgrS7gHRK3VrzUtoFu4z6DI+P3LobMP
os18lHKhTCdgEJL0D+Xt9qRTHwRQp/fdXU4wL85WyOi/KidTmmku6sAnVRv2s8xy
Ik7tTbmsAimimyxPzoUzhOeGM1kJ91PuMiAmO4mYGb++BBuSCot9pfgNzasaXKWe
x7nQSN2JU1/MIM2IqE/ygrTc2oSZVF3AiaOh09QqkDl1T+a1sMUinDJOMD/47i36
zS8wFZyn4Xm8gWIuQX7Hpl1uAzPyIYVPN5iQqs/++sexE6dF4//kDCZg3HUyovVX
g+02H1ASf8UI2LtZWKsYEqbw1Uzz6qUVOQgiBQMaonh15xkI4p55VTV8tcjjmNUn
moyWObsrl9ErBMcUw19mpQPJnYbl56JfltMijBGj1i4xXhNbSLy14GTA3Yp5m8Ub
0KUv3a0gYLZnc59X/yvKG6GyCgp/HsSIc/C9dsebdtTuBrNqAbHMnADgiZTpDWZB
ZcgD1iG7hPLIseYLH5fV5YzRee5QhIN1Y1BlyY7C8OFPS8lL6mv3Oxcc8WFVlaGW
Zexr5xpXt9xQnp+j8MaXWMiD8N3F9P1sEEUyMN1hmmLUiDjJY/bPRteG43q2wdp0
j6z3/yGGPpVyq7JBk0IfbnUYNudQ6dhbodvvmM3rgD80zLC1/H/C9Qexjr4/AJ7B
8pLkk8IXpL2hB/hGqrw0O1Z97GkIDm51Now+BfJMNn1D/HWIScwVERmC18Y/x+dD
Pl/mvbitBiynXQ1CdUbT5Wz2VEh30lt7G5NMKz/ggZ/wmxIHoPizjOYvMHHV7LE1
lsKxavfTufAaFjGmMxBl5bIzrTGzt7BlorjgnaDyQm5Jd2j/pNajAmQZmCdkMCtC
Sibs82/URif6rM4YO3h07qzMb41bLQwTjNhnTbvBmy+IZLE/hWezLl+filCRHQR4
CKdZqKGFiHy8tkeb2zV4BDvxyL1KOlRtWz1ZxutA9s6OcV93MZXXs+Wdup7hB3iD
y3fgtmrPDUu2aPN9GZ6AYDdlyaFClFqHY6GBFmPcej1DFVxthAN4PI1VAYETtAkb
jOqqy6DPAag3qBfRmsbeSmghwvmirK9GI/epmOw8A6du4sKosc/YQGOhormzw+n9
FUdNkuKwSEnWo3nSC2lk+faRsJjSyIK7Xdc/FUQ9pJ022GJPZkPn10dbWQwzO9G7
jF4fxVyFGtB7GsWrZHtN2gMffE8IO/2MM7Di/ceFyEHiN0nabwc4CQLnYKfwsKBk
Y39lKWMpYucCv4FLcuzXuWLdQ6xoMIcnAo+PElKBc6Fa2ppxWGLo9w1Agjpw7HL4
eEC52Br8lG82B1Af/AV+2X6b2ocwQJs88SpcfKWt5U1g9V3+JntDwOtayg34aDXh
GPennzceoJaXY4iRIHCdsYzs/KkkrbdOrZNowbHM5kgqGOTthjnJn5CyObf1lMpB
NyTbYkea3daP8CVHOfniFA2gKjV78hq1kB73eAQQq0A=
`protect END_PROTECTED
