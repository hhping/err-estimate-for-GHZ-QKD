`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DT4aueD+ULaoG7Grj6nkVhPl1ytTI3FJYR5tXcblmh94hl2ZT8T/IU9vInq65mfL
0SSB9B8EKY7TPA5H+nV/DeryguWhAOFhSca1G7SahmF6CnoXfv+ZFfjAHtt7SHkx
bx57fGFsGig0OqyIj8xMUuf9yHp+xmMo3gZB7KO4kBN78tfq3jNeGji+XlcP9WNG
rN/t51He+sfQBlFeeY+yztH4XpelUq6QC6gY/0POrx32J0Y8MqEakRIB2wJ93Hmu
4TPI/KE5QmhwGlVPHGyjKjnngZuUVurYikkW0Gx3u9gPYbdmAjOT3QBXuTmd9vXo
MfOrWUhZMZ7RiJRlP29PHeIt2SoBiHli4Wa/yJwB2ioWSqc8+on87qpJzr4b41wz
fyY2ARjYePFLguMkuSFDU8IBUXiYUZiPE2ug0NI5gZ98/ebvqMk77CoC+fib9Viw
dxZZYiuLAA6Ujdku3jywXQLrEQKS9BEdouIKYJTsk3aMZkQCjJKa7DngsOMxrz/F
Xc1nf0K9w/3qUgOjqWWmKyIgiaFcWO5mmaIJocPMonZqXSr5B3AO2LQKUn71qcwY
v+tVLbV/Z6k8s/X19333LSGfHUnHTZeWD09emCo4obM2WiSZ5N+l5i9b5JBdKM7T
GtWXBNAXFOimfMfFBxyZPIyC2nGN8KjK1zS3q4oRH29+JFuXUM4+gg4MiI/4IguD
PRX5DYQfTPFNj6cfMORypRjes6BBtv9oYOycpwAW0eZ0dL6s75tjS+ZI8/xKxh7f
QAZk1/RdzE/J/kUWKhuUKL9AAJ/Dn9lh+S3skKJMJoPes5YfocS0w+BF7JmJyj21
n84fbT6lgS5MNNzCWAGwljfyT4m108lTnr9z3xLT5m3Y2tKr171soedG1y17iIIA
ODgaTK+9Lr/goVZEy7nGjI6cpeXYuVSzu25Mp/MLWjS0RX3EbKVGUbViUBAw0+OT
u4pCHEVTWxPGBc3++ss3hFKPwUOR+kuD5PktamfMwgh3Tjlv9NFzN/fi14ciUG/y
9//cdhgfnRgDG3R2y7Xd/78eWIMANTiG5xu0xkIfGNC1sKVu5r0MyaxzwVTb0OFc
dXJqVDqsxN3Kr6aNXWcmp5Jbx1hw6I8cYZ+9O+CG2iBbQ1Ittha9m8TLcVf1hg3v
znnAZcfi5qyjgjDoej5kAKHrfRJVn0bZKhRR2vNe4GaNWRvkeE5vD9oCyrJ774Az
/ehGNnZLOND0RGQYnrjaMPdnEZ6Afu33mDXnVEUE/j4S0gGGdlGx+V50MijmGr3G
POj895x9WI0vsPQhIBIAT6WHx+4mUf+Iov8zpcloAZVg1w2ZVx4PqPZiMsStWpbt
lHIPKR9cxP56IPorUXtOjf9NVnjANWsjbMpLuwiOzTK/8kNomhWLNwJfk/cp9akp
TjmEAKk+5k6Z8YkDk36IA66JKsINT7konEd+294azcfMYkXsRzwZkFQGb5K55uDn
KIyXuoz414W8knP/Af5lVaHYR72jPJZJr6YySkRfn60bGrpilkaEdYcfIZGWr/ZJ
guDAVwLVr39heAUPZExDH4IXQ9kqN/ThORfSPPmFXrzCc4GLNv1JnH1nZorvvDuF
L0mCbrQbDsCgVMS/iXw1T5Ek3r1tkR9v28BfLImrzI3OQgfAFXwhJaXqzAFFnh7I
uTzsU/qFYO9Vqg5eynnL2P1Lo8ToPBBEhmiDut+wLLNORphc+/zFRyAXKCYiEAwQ
xr6WRrKrOi41EUTO/mGhryPPcYyDJ0iaty6PfNUb6vsMZ5Hlk1fGx4MFuNSWVPhE
L17wbVJJ7KnG4TwpG1bV9r376IlESJTBu/JCmYD9syESC0eoNMHJtJHVoDKg8LV4
1BSws8zQnWW181Brxh42ZWjeSookre23sBrxpHycCSJse0YfOOU8W5DT2qykFWY7
Dv25gEkt3dgk/6fgFe/54VA4d52CKxln9K5/cRINAOMshS8JLSRRXPORU9LXqbTO
fefjsthjoqoq2LWYz4CYK4ZWGijiyl4tB8imiGHAUop+QtlPdhvIIkaPdDf/aZOY
st2BTENqxQjDycKTxik9+pLUFbud/fW8XQM8j946KhZzkL9cwHhQDprlwXbPKNPN
CwxjuQRL7LyQeqMTjOqC7Yui8y1TdZWKHSO3ZJiQ13n4m556AJb8/QeTHXK3xAqG
ixaLIwVpkdtRk7U/nBjBGnFOSMYwVdHQMFD+EwxuadBJWqOUQo3JkTEc8KNj4/lJ
+hcEchc0QGtlUSvmC7XrNck7DDArlqASpfOJhqZrQBm27C63i/SPPYT0PzmLixoZ
lSQ9VHJrBB1LYjgaCRzngaA/urVZbe3SaGiQbXtaMPo00lUrtqN7nW8C/vY/wa9Y
5uljz65qA2WqaJkQMTjWWqTRbXYWDAjZjb2Wzd6t6unzzoNZymJ/Sz+ZCdjphYcx
KkEgl6tj0Bci9aVaaV6AznOT+y4yznugTbEJ6YBNRxkJ1WsidSj/e7jZJp8wc1aX
zuTfauAvRsH8H12gsbA+kccPs422/hGTHOTn0P7aPyLvVeMez9wdV+QpA9AKo2y8
ivR8LWZWPDH0+T1xJ75hhhftyRbokAtRW3IAt7kBhMj6ZVm+fCInqL3hTiPRdjom
f3mKd7q7jtUWLV0cJ1iiCBluQCitpgzyF0M+XB2oGOA7UPATEjPd9VOSeSTDnehw
8hBsF9v99qXo0guJUctHaAIlsnvZ63JKO7sRDFZSLkJRwB6gcsUXlot1LrXbyQ15
VeaASJQu3gKopqmtXVf4R5Rdg5BLEAN/ob+AO1+Artlx5gPY5CLfM633Uc9QVx9s
+povG0ns8R1TAcPrxkhUaFgpFZUyuxRZmVz/jIPVNc3khDYnFsB9UnAsLkL+HQuC
KAXnyCXwCqGp2uVz1uRfNjyfCgcgrWukFbSAJeqHFQcXruSS1UXAOWhq6j1ROQp1
pZSNaeRmQIreRG1madlLIIE20EKS2QPxwnNnuJGn9y0dg0OOvAmBptUZbeXRrO4L
yVdxlZ+3t/3l6p1pAy7zXeoDzINlPRL2BCnubyOSIhxkxluDELuaPZNzxCtxDUJ8
cBU/xuqjcAj6TrFeFsv4q+INsne5vuUvzJEfhB0Sw0kAu51VcOcel9v0DXTJQ8GB
qFYx6Ia13Kyp/MmtZsMpeTqLTYaou4FoLjj2rC8Hj1G2lgDIdzPitLy4StNt3ApQ
PnvXiqFKZO8lRmMfTg/df9qr+bZp+mzHiupw1TeFVO7H44io92dMogfoxgG5rGK5
2le6pGeXAJorHDUk2yrZulp+ZUgqeCVNNYXwGpjUXf9ur3FtyYwIJQsKzG9zOcCy
WuLMkYUki1+QhggtXrOf06E8UcTbPf/ByjMMbR9v5D6L1/HTHc4UEuESjntb+iYM
mD7VyUg0/ZUP7d4T4LalC/i8Kwu4rq6EP8glFSzw6UlpSnNXC6PjZBmNNoLABart
JNVx81vgc8sBkBoDMGt7i5aMMh70V5NJU85MjG+auRHj5/Vjz8Rso4rfAN4mve7+
56UdexfuSKUCGH7aixoKQqoIBqKn5HbGsNNUvvJDZ4OGm6w0uwTYoXnBcW9XyS9o
m0VBQju4QCpcbEifu3ti6JpkeFV4lGNMEW+VwOCxNCt5vWzsWbYkeJhP7m5MgtOM
IuZFokGngvybhe7fAeX+GEq4P2Pr4S2w7XQLtROFqueIPrcbGHKFeatMlLKNplJg
C9fy9QlHvUDzIv0H6rBMFg==
`protect END_PROTECTED
