`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+16xrNkfQb75x3oBvRFwQ2Ht05RuLmT3pyJqVxKjCOJ4D9mAcU1apvFdjjLjNpxi
oak6MJY9Dn9vhmDLylvxIDxWZRHBBuAb22tYizkQPJmeCeFNquFGNkLeTrasIHe4
RtdZ2mXdi6iJJYRICnAozPq+TFE/Th5RE+bIpLVBJUzE/+1pHI1wCPhxN6Ewcyci
aFB88tzpl/pAY3IN94fdtWqVBa7v0Ev94eZ53QaF5MdGOQsmX6f1d/B0Q5r/owAe
0tPYovI8llRvE3QIqnaX89CyocimKPPxugk+CfQ7XQydbQTFRabjaRY1ZpNQzh7o
rUpjAb7gSA3miXQoiTkiYdXKL87EdUp++MwgjZIopQxQ+oKIAE0H0XN5IEUoV+ZS
fjnPj/G7jSJyWpW1BnDrExsK1M4UTBcdatRUL0e6Uxribw3O0CWF1l9v5qQiH8L2
yN0ez7v66RNtC7o+Y5T5d/utkhQezLpN6DpzHYnetd7G0wl5v7WOgfXdj81foh9k
0DxJf1p3lyBnlG4FGw2813ljA4niUwqnSqVLEwroCWW1a86a9zMgVOxAOp2vaNu8
LyIVzjwvRrwxI17xWlrqTLI5Q9PxbgWvEqaN+bIP2xbAbHpklxyFXqBDpQqdYNnq
ToPISgYMaZl5R/NMB7tE6mugaHt1g2eAUNze6Oet7sSWxwbawGCx59YBu2J9jfpr
O9YfSAjkmLseOYYjTWjciTpDN+qEk6ldbz3sN2HvAPK2EZswjkCz15zRv4grLMZY
IWkOd2m+aEIhjHcSd5jPLbTxWK7VXuRoWbu57YUX03B6w8WV52r76UyKwcDrLQnB
4Cl8fZK+0fpnonhwagEQyw8++TMaqPN6Cfh4kqNeYSI9J2L7FWV6ThS5o3HbmQdR
wmScLBL31V7ZwdaaJGoEDzvLWnM27+Qtm/wF3/TpaiMeilkejNwosu2rMeIa7PaG
RPn63gIE+/ctdprMD03rwMk/SJqh7Ae0el/Qdp2UNO9c3FdgzOCRot3yvliva8SJ
8KwyW/1EMRXSgtSFxtDrmbyBs22x6FRFS//fmk0Tl/3oKXcrWrnwWRI7+K6732Qm
`protect END_PROTECTED
