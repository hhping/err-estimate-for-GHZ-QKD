`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oit6LA2DsLsJZ8imTvq0Ww1pRf5eWHMYLFKYu1spIu1/NSH1ATzBp9H3XeMMg4zM
kO4kBZ2Gm5qdBhbQ3jXZGwn5WnKxvUlIjYoAvsY5CzN5Z3B8Ptj+9o+pAyA14+jh
Q7TiJifTNKHqkbtmAKkTWiEN7qtM0k+5EGftWtuot45GYKN4VOUWqK08emntafHB
tCkjM4hjmX7WwaevqHdDK4tRghJ/uN+DCPzfq6yo64cY9Yw/rp93WmLWbLDPYnoR
0DxKsg1kNGbWsmtA4D1107vKdIyVXk0jtqjgMAAn+ReUEtJ/eGkfcdiyiJsv4cXW
XlrleK3FC77/0lV55J36tu6XiHpo9sO9IhspQlhgZbjlsN24GuDJSjNLDebINQIK
wmP875Uj01yH1lLMAWKyGPC3kp8329jPR7Onut10ReFUcBeBkgRQYNFmC1PvQ4k+
z2LZs9vCOuzzjcyfatW3cQ12t75NaN1X4CfXXaG3mB6DBH78Z1aCTi514EXfhzjQ
aVOHBAVX7w0JuAHqtD5ZPMTbHZVLISkwvPTRvwPDfGXViWBD/8ZJsaLvJ3jER1XH
Bv0H0304CwAsxRIVbGScliViHgN8bG7N3jV6+95CWWwQjj11SMSFIxHOV3jNqEkJ
SAVuMEnNSUY1KMXC4FmALHkRWx+Utwo0PSr2niZNz0XqLBZWlnW3FFz81GTMPBNM
HUh9gcjbB8nli1nT92gZHi9WzbvnxmSFMe1s+RyICnjjDEpgFSC0oktPYXexhAuo
PcGhH5/8I6sORzVTqQRWiJbHQweXg2feCi4AcvZFHBI7GABx7xvbIW4SyQZlr7/7
fIRZ3UAxi+lR04e2D99nfDz8YYMe0T0MWGbwaVgZazfUkpLOMWm13CAS9/vxOws/
TUi/iWx4MZ/vwYX5r1Gtw/ro4wUBxnc9VlLEe23lmg7cJNUGcu/VcX6G4kHJ5xcs
iXg0aaKZiWC07C7Oh8DXhlZISXanUPiF4IUz4JLtMbL092Opo/6CCuZAvtppHGTx
4/huvebZttiYxb4PaE35aZFG/5mZIIVmQQligknYl20m49W2DSL58ebRt9MU2+t6
Q8si7QM77LVWz2OZfM3nBPpdGv4IHIZl+8vWZHD9Xs35HZ5H+52ltKheBvNDSBDr
nXnpTYkh8t/1g1vvLLNm8guapcPlDTlUhX97UKVqYcIKsLSP3rI5d4CID0iAHJ12
XGOx9mMhJwpkEe+06zo+xJve2SOQzaO9d+I9yJs4wDY4AKo0eEfscMi9Q+zip0RX
g2wdjGV5/QdPxpsOyoIVcTJOBi1B+BtAxv745ZPgm02jCbrBLA+3CoeuB3L/fsCt
zLhP7A5iMf8q0tuX7U7/jpbUwENyzwPMsyJwiq3Fftk=
`protect END_PROTECTED
