`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cF18RaWUt9lgUpeoAJ/oErtKCvGH4Va1jp8v7NSB7H8owXbvQ/ggjS6+SHdPu5yN
1ddQhxDlgg7uai/L2Vs6zjHk9dE5ksYxZOwv9Aps0rpktRprMLujSIUT0zzGO2+r
+IPGItmHNKjkXosQVqvJ9LCcdIY5XtmallYLHq4pSzhHQPy25lXLQzKBYgJRkG1k
EwWR83BcYHrBIafPX3KVKDZNRZUgKUE8sKh7746e7mFijwUvheV63IjuissJiRq7
cybv77TIgG5P2ZX0HGoDL2RdaJ1RumdlbRJGzs9EJ9va2u9tKXdcPeaWFMY36XBS
nh/f+Dv/fJ+rCsxPBkQPBOyDeGr3ysWNBLnmrBQGyRmI6hewXFZLPDG/TA3WG+dp
cTNOmZPDh2mYPW4PoPy/RYKEI3qfrNuXL2ZdOaV9pLVOfVoN9NsjV3AaV/kzlWbc
EhopByWwkYbP1htDmAF9tnHAZ7xeUuaqwS5j0EyfNloRDuQTv4Y5OgVbQukLmZFN
KiBm6mIN0AFQ43SBuzvez/f9FlaNQQ0Kolc+fWmWhN+unUtRGwNvTnvz7rRDo8Tc
x/Phrv1cusogCNQ1lpX4Rt3Qv6DNuE5kEmjM5ZRl1c2EJLAMt7ASoPLwq9WEHTpx
iSkMuuTsKQt+6wj/awPrjRIQBEoQCnko9UQj8OBmHhUG5s8jnZH0yOqWt/Ee29WU
rydgfsZhN54ixNcxCkJKWxIGz4ArDkVNnAjWJhRh7mMhU23NyhAk+L2whlESPfNz
ErCsVRuX15bUgMRHQCNqWYln6RfSEKqbvyT6KCm1Y3WTkR4gj6wSMqkwDdZ9lSTD
tiD2e54TYjQHeS3qMC4btWnrpEmNlhtQei74gDpx4SZ201CRBmzudyGRRzUUf8TF
`protect END_PROTECTED
