`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4DR6u3YO0t1SoVPoWSsPS5BcAwObbd6tfu/LpzfLrVTN5kjElmj9xgz65bPHZDSW
Wrv6UUE8CQjeLO2C+jp8PuGod0Zz7+MbJrKZci5AX9kBVSGLnTDu9JzrzkXOyN/1
pCjn7Z+6GuqVvfIqVmt1aAZ79nW2pA/XdEQi2Hsm3TNwdRhZzFKvuP/u0bGB9379
yuojjC3GAxe6EO9F0cENO/l+9MjfuhEEVcozzZfCIMXWzeFUn08VrcCq+vxs0Tvm
1nBBo7pb6VMCMs78uDht6betrYrKI0mtzLJz9rPyJzm1eHbRHdfWXRlT7aNrJWY3
nvX2kHMxF7VAKQty1YrL5JZMZh5tiS5d7+sDxqAmRJyH469OrSYGsu4o8LJe9Weg
VXyTgmIZKQuKyE5qBpixWv6tiu23w4C/99kFJqkypzuzL+53OtsPTVeETfuug5f5
foQq3N+VfLW7fVW1IdSvdKGN4c6Rgqloft6olDpCItPBwHkmsZc+m8Y14qFYYUzA
SjZmIm+CLOxdb6xakoTKHlZDs5S2n3R+ZhBfMTdz8lzPowR207j2hkL7Rz6pLA4r
nPxr8OiE8UEDZnNKlGSdYgjf9tdV7fDNJ/Vbkp1pLut2KXAFfvHGfAPT0sbjXHKC
+NtCHE1RJRh/En4Ef/qeqRWNBF+PH8w0Gjmc8Sd1SRpm3pm48kXsq0OOGCwIn4iZ
0C1HMyYnWdJgmS2xuXNehazxZWWLoXj6muDnaNQDo1WmHezTanYDx26xPkK0JFiA
NErGZFx/XeZe+Lk7imSr8smxwcuS1m8sO8pQ6H+QZ3L2MVLVl48rFaOZRdHtHjgc
68xgmaorN9HzpWGKipkxLbySSgh6IoD4Ww9jiBVbYsXYhxgOB3/KvXbeRLKollw0
r906O2emPWUKRUMmblAxY0s6iS6Uz33nqpSjDSt1M8sCRsMtBiRW5Jb++3/N/u5k
VXHm5eB4KFQ0vBCbj5WLGGxIme7DZwtmNbLVzd+R+k7d6ufJUh21GFbUuQGPv/Yp
jpJQGIUxzYAhL31MawCzT5INxzmIjlhLD2+n1I/ze5JLRh+n9gVyEh5ObddMbJD1
h/X6WCYqqUaoc33i54A+zovNOB2Un6kJUcJy5/BnM4WoeKOrjCE2+m+oUOhiLIDP
GMG1RCNcFkFk6i/JjMaIUcLd68caKN0J2FPWHQxZhd1PEhPr1Wg2OrcI78aC3Ilf
tVtf1Uu8Luxddg+5T0uXZf+TEG9OWs4wZ8dNs4WSzBfDUIIirwJekbHUgv6JiP6K
pcEPnvgRpCu7SA3e/X1YOiEpV/fY8O9+qU+tDPUw3YGG7AzF2DqzYvPpUkbMTvKQ
mdMY2kO+nvrt1NvcLg1sGfeFasvKcwtJ9cgxz01NniJBNPXx8BrZFjuJNDgXxykJ
mUYYyufLHj6B5Y+XwSKKgPgQdetIFDtdZ/TEmqIzYX3YHAd2lr1hisLC7g3hU06z
pGxLE58aMfFs0oVbn5XQ8OexdviwVi1QecaAA00h6QVeAIwazAc6AoFB9y7jxlkA
K88kCuI9JaF0ET5Lqb5qUtecAb36OqGiEUfaE0JkA8XDkU3GWNCM7gBXxBauR/Rm
aQ850kXj4LOeyaLs6TNBPG9XCrYaMiLUAkQ5Hht5mKeGqaa/AZbbwSKD14SnQbkz
jtIjLvaK8nqtpC9+0Ee6mSe/Cqa1iFydsjO3MAfIse8Fbdo3b6t1ylcSaBqB1rdS
pCruDv2ifGv/u1ILil90a3wYhqAWRl+80pVN2Km+iXUXDj1W2SjX3msErLksY/5W
1IaaOIMqW6vp5uSsBIXsNApT45G1hykDVDB3ZGozwVc8YULTmTKBEBhK95hI1eIx
0xR9WERR1rapAGEegjQ2eu295Gdmto8clyLvJJTfxhSQtygQeKKDxhb3lwVaoRAo
6emVS9de19ZovvzAnTYNi84xLBGFBg8N7whVaEY5Qa5vmi4kwU6sgS9KXWu5XMYI
MEt8B4qc7pKJoXvZjlAw+lKKXSnK/gnHn2JQt10YSpJ6/eKMAg5T+ssDEkKTmpP0
mzNN7FDME+foz/ZRrOtiM9oW/xw+6oX0Unk5qmSGrhrfdmfPnxSx5FTqTvqHUTjb
9su1gB/grZntpbBXQWxUcgW1DgVtwj3RQvph0vPIMT+P3fIZ/dgYZqsGAEiSgO/G
4pG4ipILdF26bc0f0JKrryh95Gmtaur43cnlPv9RNPE97gS6bKjSAjsdVppTJx6g
t/3+hX/zAfABEg6YWeKLnpoEJ8FuUvzzAkk32FauF3L8jH6SfcQzsR4mjj62DOYS
6w6sXb6okCC94L3gRWWxpQqVEH90lr0TOzcgLdMRL4c1toazebROlDZAPVkQqpZ4
w49g3USWvIjFMK08H0HD0Pm1ScKpg4ss+rgQJGhCZ8u1hdlaJGTuBWypTfS7xUJL
DKEtsAN8lWd4CiKfhCMO3/CvuoJtdsVDMNUKoFoICyIjy9vg8zVuZHXt9BXm1XSQ
TQtXh57PM4EzdzHNmp0FM5s1dxt/+cyVgsymwXyVN1VYx63Nvxu85MmnZzUl8MdF
Z04Gsmmz6bfXRVv9bnnYryemyhqgddb55J4fdTn1BMMpPcV37NpiqAgp9/zKW3xk
kkBo9y5TpSzy8vTXezMzlf7opmjOxD6TYO8d6FsSwVhUGn7NUmLLeNtafRtAUj0m
ivq7PP0W25u68FUgXFNBZBt4X3N3qfJW6WjuY/GGOIpVMs9iFc7dKWztv/Qf/NBe
dvP/NqoptRN06lTUgRcosojk9Zodi2RwDt9ZdQLKaDPasHen+brGnec7tOI9i3e4
NnKgjXD5RDD4pyIT8kdReB8JkhWJEsUIfC3w8mKuncAQkIyJruzJliUa4fP3L4m6
1lZcP+LpZ+ErzaeL4A6Odu8OkQqUjZ3CLQJeaVww343ygZ0dY0me6FtgwHmH3xl+
XZEB5D2C4qwU84KOPT7LEh/DJimWSnN+I3YDC+20jJzUhV2Ax05EU+Iamho9Qh+W
8x9qzXwgeDuX4iBR5lpEWxO9QKtErf4c6vAud2/f2g+Nbgrp3GF77mibeJqGRtmR
q//HwT+gGRjJHZEujC7HRdTxbv126Pu0SVQoZ9b2T5RDoo5ldWWmkNpZWkMt7f/0
dnD+ufMALmC/3+g3QOy9BYslrblxGXRXy8kDP1206T7I+U7d9OrvlWw3Zp2UCJq9
H9ZIFBlpO/UOTEXiRTOiVQ8eZHDzZOID7X0C3RIOZOjbMbqTT0PW2AROvK2UKWwU
eAbsEFPGz9Vadv+hJqeo0CHvSwoiFQwGItBWzTnqARe5Ob/lurmXDgfv65KcuZxA
bptghmYKUrqzx5/2l9ZuEXOypTWVqxg/ljQc8GbheyJVHlBkN2wD28uo2G23Tmuk
G+TMnLtwRVOKGVkh7kwCLfx0UfG+KfWm9ZuSViJjGKS7rw1abhjgYcMonegBSvP2
yZ1NFh0qMY1rsQjkJ0yQlr8J9Yh72U7v8w/qAj8hnj9JA/cqehFjUml0KK4jieWt
RhO7N8ia5SFUE0LYy1WikWqyv0Blh5s6wJEue+l0ByVwTyhOc7DCqih1cTmcprDl
T2fSofT9X/QCl4P48zklg7PSIElg2gvdeUl/7vCPvFdy4U9kfCRQbUkzqOQhGN2t
3Aa4/Xe+IffCsvw2LmNTO+8N5T7eu/spCLoYlw90MHIyEJHANEdA+gAdSXaV5STg
qKCZO88NLnlOVFuHJwETiOTR2oq2A0cawz37D/U9MdzUl8/hLqdG2/iHf0/N3mVX
vWBbZdFnPwafnPfQxpjQwkAVrybO6f3jjRteFhOym2heQ7EE+vf7ARVyW26EqRjf
LbeRjNM4APcpBBZDajWt6HDtNPL27/+pTxhMo91rtBqrXJakNKhjhvmPnJlbSIes
o8Lanl3gHDzcTPMTyQFt2m0o5NYkFNimuZPSVVR/jRWEuAZ0hfI0RCuySSIRYtjV
udSK8osFqYbRS+fUq0umVa0IJkCmEnmXsLuvTHQFkNO6x4HhuEZmYXOyR79DzfeX
iXQV/hbR7xJnszepLHP+6FxBuDQOH8qPn2dKwbFxAATmbQNBC4Wkgz04ltow6JYQ
MxWJC+/G37XCZyU5juFjHQaM7uN/FsLHgEoOMvggpOfyW5IsmPojERQrVU1LVmCw
iljjGkeho66X9KPd5X0qPNb16cECkOVXNfzvD3k8LWjI5yeb7z4nmSNuZiKHkUWm
ceu3ghJJAgXN5m/p3rqeXkrcnTGt7bUyGOkICWHxHGu2/zOkAeYgMn6Z9Xes+/ah
KaAY6r647AzVpKa88SD3fScLB9TgdEsii7k1wOFSf3HpoHUqPNSP5cwTh3yiP+qC
Mjz9W+FlGo4SAVQ7/hXD7QgUo4iPfRuxcUkpJIHWxv+VJ17KuvPwSQygB3BhpNmu
j4tzhgv6o98+si9EPs0nzoQuIP06/SMOwZ7Ei7xoEs4ZDViTIL4yo/LRUHglGz6B
`protect END_PROTECTED
