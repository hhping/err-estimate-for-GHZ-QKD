`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n5ycIVsX1MdZvUVn4Jotqdg82Tcir3MdWu81yI4GZ+YJIbDCeJy/ip6EN34BJ9xh
ipIFA4xacW0GU0rNxbRmhg4sA25eRPDVjxlg6Zf0uNZbEOvRdKEnl62X1gHkQpaY
SW/i1hWOh/0KEYggO5lNrCxXnjmbcBsXzudPPyfLYugLQAhxtHc6M1gkIrxvsO8c
o5Kj8dSeWkDepiDx4I5to1VUaKf82keUsa61Gf5mliryXzCampmyraNHJ/orXgiX
L3FSSHbnUaUtI3HrHJRN2n46vASGpK72IGKijpMIZxGOKGnUsfRkKGY48wcEmdBO
rFnKMHb2h9Z7iltmrs9cwjVE1gIDyRq4HALPv+vwmDpr/SZ02eig4bdsAym62zHe
dZG+jX2YgM0x1ST3yLw850gnD4JNSo8nQj4d1cUg+Zzo1Kgoqr0Nk3GIujxQsWaX
dFybsKmI9sDAMPPu0JcguCFM4sUlMWX9ZWzAZZvJ9nOzXePVL0yCK3sLOtabYztX
nmFjz6AC3DjKwBjBsEHWwQgLfT+JhefZJrFuwKurj8/g98ftoPijdrwYhQLhf1J1
`protect END_PROTECTED
