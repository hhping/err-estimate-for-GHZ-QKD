`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J1OopdjCpVONTBo1qq9YRC12dQWKBcrVIw4QmV6KUkSBsGVWfGp0rd3vfeYuFpjs
mNxbvucseUb0BLE6SAZuVdgx9HY53E9l4Wawizl/9xD7N3wcvfP9YFN+XBtpu2Vz
swmxM4AwAdPIgLQXLoeNRK3bc5imEU0LPmFCp2onVmrOGYPvzDmumsd8mW1YlS1M
Jip4NS5dGITOsuED7jgrw/AcsHzAc3/gQW3DQLOeZavEYiOqusZPQa/6XU1eyhhk
67B7Tslpyf8JQMSpX+AMvVM7aHEjyXDwWYaoHnQl3miqCYjhPGKvh0nEEooTS42X
9EQYfAjYtDKG+vYvzMiEYaEWx/2jYXAD9SHoYhIhxYT5tH7/55QkGKADh/f7IJcr
6Kpzhu4hOiSoibCiAJruElEtNykeEQVwr7XbDu5ZEZx8tK8juHORiboiwpflNuvX
zNK9KfCMgTYAPSdXFSaPhgn6CQN9rEoxlHm2PCqIZGcldhE/si1qBq8lcJ00xm0N
EYshGfUmDNoJfdPHVlVnmbla97BI1Q06tdBT3huBCjbaLQ6o+m5H64xwfJH2Wn2+
Ziosf1puMcrRPyQbRPD0WQaUNknFDaRsUAA/m7zd8k5yVmCEGl1grVqhdtNvSAog
M2lLEyWhNx6IvA/8+k+yPbiM74WBHfMAPP3DWUDqMztpn0/ZHD+Ezt+q6L1OonGN
65vDMToudLo/JimJRCvl2BMrXXIn4Tez8Izh9pPt1SrYMmHv3PUHbHklQV1wI3ii
VKIR2jD26JQCvFcScAXt7ChNG1CkymMYucKp4k+qlfrfXZ8q9eCln7zHTOfz/Fam
OygiWb4pIrQ3FF/cCfF6ayqAevS5u6raxRCxVMHMp6nST3IzoCXIXpwIThqPp++b
+X2LgbSxWnYNLG/vsyZ1c7CaC5SCuwbUtao8ivH4OAJiEcO+aD/jIjbhbx+eymy4
VQlZn6AYQjLo1DmhVolJcwUjsggfvrapzYPU0tUJ9bAFN8tb+/30WjUNSHLPE4eM
dOz2BATTgi+L+tB94Iw6DEgnj8ZWqrdXXmwINXwK/TKlio3aLROn0kXemrKPuuXP
bV/sDi4e93nwOQTO6O3tClBbWhHXh7KlXkQEu95bJWX7ThvPPciYiqvQJsVALZ0d
1F7j8Y/OmkiwSXRdbc6JIAUUcCZ1uFm2/46ZAjuxyN0JLzYSlOtYx/paY5i/tYvk
3/ydia88B2Y/eCcCuTvKhVMekjEfBk6BtiOZtbtMhxzUqR9Tj6Zcg6Z0gKU6yBUW
lxEUqrFE7WhYzvPf6rZ7fqaRPhfLVLBJ8X6kwiXRBqeNiM5DMbpMPIoS1gxc0u/d
Lv35y2SCeFyugas7rqxg/JPIWt+/H8boQnIxMqli/yPzc4E5EbXN//DGQ3EEXYVn
3w4qrOM0K+g8ytaRAumsfu1yZu5fJZ6oQ6vj4nfV2ntLWytDD0k+u4v8gdqBaUCn
BKV/pwTQ9gNbdqiUCwxnLMWqpmPwCl5A/J46rvzhItE36L3lEmK7LrWisshwqQzN
xQI3l63kUFlMmPAfqqV1m547CFIHD/jaGZHf54J9ZDsen6uMKygi1IfEoFsoE0k8
DBsG0DBsvjVvMme2xMLv0Wj4wUBG3IHAcNEIk7AbXAVwsPTyCN/b8bZ2/n4+SN1i
EkUYPwSSrzvqUaxkJsTTEoTyYnAdhghw8kUgC4LroOMqEyNrBrNSsClc7Y80DGjl
fB6UljdxKHgcC0e2oz2vprbli6rIMpOLJvPPtFyY+Z+/aQrRzBIJIwM/nIzVFpKk
pQhNgXBLeYD+tbU8yOnOdjDWwADvxNWD6TvenvRHypWKvdqz/zpTS06XFAiDrAQC
0JlWfQ6Y8RoqkWhNBtpgAndEvBKuE2cG6NjVxXB9nksLeyFBYpUgjqxJkTB+T1uW
mvLHH1T0oy3UkVasWumbJ6ImgzNnMnVkKMnbX2Zc4UaSPw0RBjaf2K+eAlwud6RL
peSFOw1v/lQeJkcnRjY5dtmlMxoa/gQudbzzYb2n1hXgzvm3xDdQdbCzrMNi/fvJ
rapzl/X81pOjPpEIHky+LFRyXLJLFzVv5yue6sQs/Sr15glCOS9uLfKzWjflstun
KiQvDxT2l1pc1HT7sz6Wo2I0YMryQmoisNQy17IMN28L4EkIEHh9zL8rUFlJkmGG
cUI9Wm7M1Lv2zRzuJhDiiuWSlWsTU05uIB/FWaP4MtU3c3onbm5A4GnQQYrBo1aN
xTL5W7h1hq7EN77NIWzbwaDNorvHTqruhdflupFFzMNet3Cl6XdYmyMTir6v9Bmg
BafA30RwE0sL9ofCYKp+757rRwDoAsuOkEGuT00YeDZyZiItAhY1dJlGK9SrS2YB
B+c1h4SRNwet3FaECY90mB7yJJZJ+efWzjrWH2fM/RILWIbX3eZ9678dhPY067+4
bfxrE/5OrUD3gW9qYhQ7Vume8D5px9YAo+UFmANWrkG4qtitLiHGGTEeVkZlR9Gi
0YrxQ3xf1EWbik45/zE4/MDVGzO0HULqR3+2eO3LPKXelHR6sZBPq9FZjGFgnDtS
fCcjPwKt4yaDCxiTqJx/SKcHK8MXLdsjsixbRhUqFRtnQ2SFjWn1I0l55hV6Yi/e
C002yYVXSZ0n899mdsjyBsQBbsBQLSaMjC+wmIXMPB3FLZM6rnCPaMySZWl+RRZf
TURNm9vzzDup9j6fo0jigt65viQmpGqMSYhFj2+bVv4ALC+u4uB5bQJd8nEjmzu1
BiHHFZs77zDJhSPYn7/iN52Mw3OrPqt9lza3VeLqKg5KvZBd3ZKijQfSAbYD3Ekz
MgNQz6gchi2S3JiHlNRPJHNgqAicY8UVnqskQurCB0Tp1RlqAnNhpcoRKt5sV4r9
XeGGGUYsyY+TavON5gvMvw5jCm3tEiHNF3Xh8FKnI2WFTXm7VVEUgg8uCYIJU1RC
utvSFNrfUH7oOE8qEJkiFO/tCGD//MLUpi3d+WFB1xERSkf9bDXUuxMzjfwZ3v11
KqqqfsFARahRs0S7sE65TqxZX8Nm9FWn8MhxW3nFVglJJtEnWGCDB38HZ8LTDwC8
/L0XjrijJFMKqT1/NSLjc1hPiF7G+xGUJJp5psuQajvVl7cMS77KdcZ2ZjcfUoUv
vTgjiKV45ZzJxDf+AbmBuf2xzFIGKDNGOhtQgzRkjYkOazIP/Gp/6VknSTALrHFe
JCms9nq0zN7js9UVph7gi9TiuL5XH5WPIWZ9Oo9kcEYJ8vOfqO3b3dJ9niTiuw3W
2z+Gs35HHgFOHWm316/Slbe8mVbo5Ctv3cPvuvyaUxTTFYhheSX8fBf0iFNor62Q
jze2gakoKa8ehD3vw3Eh3lxwRHX90WOJjkhU5ImFXnp82JhKgp5bADMcg2pricfv
1Ny/erfz/mPOKQf2K2jzPg1FcnDTSjjQniQ+zurAR68WLLurJFnMswOCqv2F9Sws
h5USZX9FEgWHvMOYrm20XopTpuQlsvielfngWYMnk4n0uPwcOVm/aMn5R3yujNn4
ufb2bzwj8hPnPddkHxk7Yz289wLmWGRk7ZV8jt83Q/b5YM/kDpfQ/ykNTzR+1xfi
omqXJKZirO2OTi8l9TQ/rWdm6dMVM0kQlqDEHdmh2CTxQFcAp4cg3/SCs6V96C/d
zcmoAC+tJ9ui0BWLXioA6SGByH0d28E9Nk7msD6TznaT8Ua1mE2HFSmlIaRTlpJK
LcBWs3IGFQISiz67p4h7vgg5ZP/rhJIjRIDnj6+9li5A84nW7CO1KJlB3s5v2KSq
uqOcd+sheEIRqqtHeyKilJRJ31tVKocOb1aqatB1eTkRAa1I7/1lNgdwFL4SOokm
kUV46rY+TIzI0xQTCOqONhdJ6JaZ5pjW7BocG1qB2oQJD5Z7Zkg017S3SYmMx7jP
0pIy+9uNSXde6eABvfdrNNkWRZctI/Tjc1ok6v/II5jwQ8VMGXVAJ6J67zApa5MT
siX1fGyh/Uo0SnZwn1EVstzFK3zN50cE+V50OJtal6k3DCQ9BHVITCsDWOne0se9
fUed9pYUj5bayv9Y2JU+bRfb1SP4bjpnVTaepsYadxX19Beyjo3Cfwv4p/VPPXYw
nKBb7v07pRMG0x9t/v8xBmcg5UQmP/fTd1DN6oBf7QCKaFsk4dRI8QsnASP7Gf3e
hr1DyYw2Hd12UemZUEM7BAHuN1+UXt3ZixMC6G6eS6fhZcbK5XiVQ18Ycq6tjUPo
8+8j4+zqw6u8JfXE4XOfBZoQoKLppkkOzDFM//Baav6JMr9CTcN9NWe7a9sSd1Zd
2u9QVTh9j9NjFNnNBa6rmsBs9XhkULa+fizWbPTOFvXxeTkenYg3pt0TAKjMir2h
bmEU5xLlksIR+VlBKwM9N1dyPH1UVJwZg9wbi+VCdFv2nS6Lxw6yC/XOvYJz2Mo5
ScO9z/xvh7LuvwRPHM07hdIm+tENziUt3CO/lzKIlIROBo+PZBBsfp8mvGhckcBn
K1H5K8ARwjPvvCFzDBLLbVWcri74RK/JoAHLhhFFkzI5mGEj9ZzidtSuZMgFDhpA
hhc+xwnqDuNHiuo6n/qW9Twfk3Udr7SZIaXnW0ZZ9GH3yEGo40pZr0Qom5Ra9+Ej
8OXVF12iMq2aC4g8dFpPycmVrPLm80YlVsxXq9TL2HHRy5Hton7K2rEVriLqdBn2
aBTAeTqPlbuTip9ZYoKROcaPQcrN33J2VfKmuSw2fR6dlqZeUV9oEf1ptKqVrlmQ
Ob5rqa4u8yqaymKlbLzjjUm3gakNPVYHcnVO2eGjqILGJTxs0NZecgrEa3kWHry6
D9Uu6HptOhGM7rN9LNodUzK3MW96FgB5eZysYwrunnlkVBw0s1muL1t74PqjMMHB
NmoKpO5Rz5+BPAG7I+lLQ7wjXtC+LW74sD4NehF3/qjT6PNnHJc+MA9Evkgcjw83
DxlmKwt8cQAVqVWIEs8BHXZ8f3jbfxMweyzgF48r7SOZWPHPkMWfIpWwibNYZpqk
gElktJHh+04CrO4VRafDaOhJDM/9ORKcC1NJQPxkeGeOCdS+8BFv+BK7niMwBG3G
f59g6ffB2PTYYE8gPmyqevQZEAmnwD1pk2EBNtG9Muw+TFmFy5crNzN48dyx9ChB
E78k/L1qayNj53eu10+7WeJvTT48OXNLbM6Tj0TRZoigpAFlezR+AfZeoPOpRCX7
e543QliNDpCC2XXyqF5Cv94mp/i+z2oseCEnw1f0JR3emn6dP6gTitNrU/APr6iT
kxpC0OEC/viDDHokKhOlWKArPDEk8/s7ypf+0Qfn3if+Z7NgM+ywMYCfw+OS4N+j
YqlUUbpoOWmMT9lFhHWKB/ozJNRNg5C8j4EDCuYGSy9AYtSyCl3NtOKjOWBwjihY
PLhscrzcIQ37vtOpHA8NTJmIM+SE2DtNE1wqTXKnj1JUg4IE4S6kdNcHJnTwBUDB
oaxdvYYRwvSapG6R+ZYG5qkJuMoGcZO7j2PwAoGR/1w=
`protect END_PROTECTED
