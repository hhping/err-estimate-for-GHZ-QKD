`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EulpzFGC0ythn9dX2xYA+k9yTTIRoDnPTxbcajZTavl1Hlo/0uLKnFkzHa/Ehzic
G4d+bxJLB0+enK9a8DsWB0bC/h+yKzcBTAwiMksXj/yyTwqvZX+OsXH9upjh3EVo
TSXigqe3K3F+N5/0Y8PQOSDsqRcAefv1wXzyKEBHzEcIVA2/1zFh8YPmw8Ifkvw2
usu+t7odGzrraDUcDa97/r+TiwF/oJcKUlnfzhmGCFAWHkUcoCaB0CHCUHKvD18q
ReZelDj9D6j1B9EfHKEC0mFfTrtQGKhjZPKJHVlWbe4T9T22EOu1BZ2p4qbj0mKI
8UXeVD3e0j1S5JN/oxJGXGDwxGIr45RWHb532b2ePlUW4+kMBlDk9QmQGzW01Br7
btA6nm4ge+1c5EZru9IfveVQ7MrEKGdu770/1JSyJ8zlmDESBZHDnpzO6jj7saiq
Y/JhvsbdMrwja+wam4YUVjYZg3Na/KxFQmrTBq7jTYngK/SOna9AAHLQlCC94nUw
kC7VXH/hhgJJxv0eoz4q5Vl+5/uQ2820a4yuRnn9Kfgsj8FuMOXXlS7RQltJIyJO
TvcHlLBERU/75lggq8Dbf2O/cuDW4dKO7mAby183ycTwDGFU17vkguetectEdBYY
bpRPNVt5XIrwuKyvMsCVLLf0h9pRENCzBdAlVe82YGL16QLjd6P3lZjZfVJApwiI
rh9UlaC68PF8TstJ5McNqEgh8Mx+cLHhdo5FkTrLgBUC2blK8sYFPw3S/lvGqcIH
flN2NgUmR8jkzkmrGfaioHbB3R06fNcK80R8tW1wRUubr+cXPo/ryZXHsCmTZqSc
UkIc2erIE20SSjs+6BQnHjiVoHnD3lUk2eU50i/fPClManOwq361Nnsih11yQ/ba
9oijuUuk5oZltoyvYwp4LRA+HWBakP83X4969W6UfmD8BdTomWkWXMSSzAM2QVRW
mKg8azVevxFM/YlDzWW63qpZTnzBTNesI2NK+DaahCy7pUvpBG0viIkgUEpR22KW
JeCOLVdjYCxQSpuUDTVyJ8AUXObPchQdBy/xzAXk0lPbKdTTfV+S0SJkZUIBwPQ5
/1DFUeqo6oyAgS4GjZVqrr/IWAM34JRmA+KmuElqMIrT/pxxpz18hIuea6p0wsSz
BOIrHJzIyJSAbsbB3TejFsGI4VnwsFQG8lp0Zg21v9EJ1MmwAg8m6Cs6EBTduzXa
Im8RKITsTaTmkm/pbHD1PwQuQbTOqTSz4PA1nO9P8MtFOtDNB7YqazpldU2x3QgD
RyIuZ71sR8RCnEOBtt6ozuLp/8w2al1xnSkEiKeEurE2BD2B8EgF0t36yUZWY6kR
JypYfcvwe21AI4XdI0UYarP3nBVGPpcdnnd9mbpl1XH3h3PXA7Xbb/b7G/f9TDYm
W5FZYz1hYnLbdaEqjHk23qE3fVo0mwxxrPwxlfnTpCs8p/gheTctJfuzMdPYYLn3
gj2IXUwIi7IYim/PqOCDugJekAfUvTuxgZVzhh2OuymWU6nWDM5E8GfDBgmDlQ1S
7JZ3DsHp23w+SNsaSe/nfKSGR4QsTQRUvSj/gCl0AFy1Iw9AfFNyLI3bGaxoQJia
YzyleM7fHdd+WsLfNOqbXNPXxPBm2uLe3lZkN05gNAg3T/HGy2XgWp96mupvQdzz
pipHhy48y76Ozk4JNTC/xW+tfNHo5e7EZhmRztjdW8lS4JYH4H9nCYqBJWAZ94Hm
PDl5P42io+ANl0JbII2Tq/E43QQDjRMjAe2XkO7qaOWfjQJMJOp0pCGuTUVqX4VN
FZ5GWf8NIDf/HM7P+8OtnufZtsAj5dlyvO6MqPb29WcbvSL7A4VBgN7QdQTXivhr
jB7e4wUY5rcYPi0HuO7YqBVRNb1ZolZoSk64OGJOvjV4q1sbYd8IUCZ49RJE0ElB
T55fsRPF+K8Fu8XLZRmUMTmzEeA8HG8DRvoOZFQw7c/pwCe22Yrm+3DVlnZUBoik
TQh40dB+D/oh8w1O3d2pqh1Ten9c3hz6zPGklFJOQA4B+2kg818GKrIbBNeKKEHM
1gpRsbT2D6+0Q2FNXhbQZgm8uzv2w0IwmMW91nh7upilmxNKX5PCxTUONQCEFdzi
sAbsrrQkQIOMqIa3ITAXXykpbJzXP8OVSNzjVLvx0wqPjAK6pOYdpcAQwnhGjTzd
sV5wzALlCS72m60fkpDVdwkLhMN4+msefDYYfiw58DbOLUz4N42qAr4BPTo5pwla
QGaUXuE4fOdF/YVtPtIgTSFWh0Gur8GlVBW4CDpXvfVyKaPpRZ32/d+sMt8C2Oeo
9v6e7Oh4YSkIYZEESZQ6e+CotBoxKAXC77bXaqJ8K/V+fFDuksC57XUgvQTMYUUA
wMecbzJVz5kh6wLchraAtIRT5tMWftjCSUokTbfG6p5tByx+2yI7u2SdQHXTTg2C
0COEIFVi/xnC52wegU6QyJCVS4ul42e5miWTtS1y+pjxcw6LYhgt6ypWAjgEsuxG
BG11dBjwxfwKrYhVLO98898W7JCeDHom8lRVlVXm18wlYw3lfuqwWZAzxTizU5Rr
RWeO6tHhQwvCvTxObs4hxT0ukkYakEkCK6rU3Y5oKUyoUtZI1vjA8nGjSGHKkOOC
j/JVuzNJPzQtgqp1Mwwk9otMx4fDlDMZ+xDz3sZ/WLJ3yw09MwT+L3qrvM/fK4HM
spkyTQvVu9zcmIAyEpPbOU4WauVctTq1yQBQsAgB/AKYAE3UgZ6AGK1fuIFy7lne
JQ87lpOu2A573zC+kAEJ/XZKZxmL2321pwrszmS+XlU9Fc59LaJrJJNG2pH15ybk
AhTGSMcZLqEwjQMFXvh2IE3LaruxsXmgwlqkTK38CA6a1l2Zk30HkVjj/p4A/kti
HIKB3knKqQHP/SdaktpqTsXnFudT1ZaAyyryaSd0tIl+cY1RHduO4TTBdT5AVQ9s
EuFv6/+lOYqNc7WdNrRZl/RS9o1NpPzdMH4iYsIU+pcK5DLb4+Ph7mjoxQVoWSgE
SGAcJVNZYPPq9gJr8Y8pcaMVsb9no0dY4i0sCWb76JTqyvB12ZCEIYupHeOo7dO7
SLYKzBUD895Pz2Y8RvH66A==
`protect END_PROTECTED
