`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dFA3+lDdLz5ppTcBypz9RR2VCLUBPhIHJTauHJTIU6cVv3FlX7urQY0TMkqB/9KZ
6kvokmB4qwiBAWAXhPSZ4cqfzTYGMh8iacI0wPyF2xee7tKOjCUTbdHcGaYLNbyu
nXYZjVZP9NepFn6N2U8jJmXEs+VuXatDB1jT2qnkFesFdq2pRkOiDH0WwiQzEZrK
7Yt2rvPH2hgQ2ILrBmIEgmI86ch68m4eXSIxdtbuD+uPHwjaOUEr/31kYT7hwbIB
2W3f+SmMDYuqcOn5GXkh0Ds3z1O78H7jGTf7SUuQurVxUiWfJFoYZCnzKlPTD+AK
S/ekYGMugy/0MQi3+Gtl6GkwhoEiHpO4qrgiDDqlY9BNZKHx+89waoWRJG+O63wl
Abussr6pS/Enp+2srcdu+JI4bCdDyCQEItDtUAo1kOe/EpEMNt6QBnwrX5X0EJR9
7W3puoNNb1q3DQpF3gtxOIqpxNQxdUMxHPmOgewSOWbpdTFDeTDnv2Vgusr5Vyxm
PXb3fkhifOShc8cPKhK+6vPa90QdKXRcKzFXHl0+66ENux1KyZEs3ZrFdWi1l3k7
1kMktDyD8liOvh6wXgjYM7NLInoAv69MpiUW0qtT6NZFFQB0GsS2710T5zq3bOuT
MPkfi+zvUw+mNk6aWzXxgGqNZBe6S8t0iKjzX0iOawGWwiW9gXhk+M1u3pnoJFPb
S0cBrYqZ9sy7oGFlmEfXku5PnAZHgEWERYd1Y8GZc3wP7+9mtcgpRtzaZfRmOYVa
UVEqOwV1038PVS2KaBUFiMUsx/LSGqSriCbvgNtPOJ5njj2oZcmWsSZuNSsZexCf
0kQuc9Yv1k3uIVdWvD6mjucWvF2TX6eP1UT+srmwViK25GwK0VmOsKNwBQ98VvZO
+vRZY3n/PWP/IAab3IQFTUhgAB7su8lf06FX50LEa9bDPWfzIHSXcKuWUpCOXoVg
qTNFXp0dik6QC6gvY8q4uJ9dQJkhbmnU5/vGW8tt6GSHkDILqEnQSAFIU8E+ddfP
znc9ptamZyv1Kdt6RhmEX4T+KKZXUJjyW7G1Y+jXBYupVf36OqNDRPs/c6EL55xC
aUXFwS014+BU2wD94fvPHHzMQU6tOCDN/Tq/wwDcIejJhLZ+xtTrdu8uYGWEOi89
KtLnN/fE5ztSF+T9Mlh73MRKM//6BicUpyaLvsmvju6CArJHWVBU9izzSydEzAzc
es/lARxB/DNWjQWuwu5d/G8iuJlXnwUyM5iPOTqOUcCaTKve/vG/WR2cveVOxemd
Xika2gcF1jPBf/UhK7JAtOGDLQS8ysAvn5HAGDrxa2QbPmoqXFXWMPyxZH4SiXkd
Yat42buhK4MiZaxmb0YR873emdePgxMVZDthQrqvtk7eJJTZzXqI+mT1aO/5EbQg
ea1oERvnGn2O4H0+FjANkNlyIjvrljmGvTh5RzPiFxEe5HtA4ZQInpgfBV34ASXl
FjTxBKxmVaEIXaupQdNk/HlXwIO5y84RWYPGPDq7YMC9aSQA4fyoI8PVHL3ADijC
1BaypWlZUGgZD4EEbIljPasBX2zNnwNDCXdHW7fCM6GLbn+h1FqCPeHTrV1LVNby
Sxo2Fgo6vwNgGIhtpkMYvJtzDe1ynhY8/xqEX/3Gf9pVzZsAozZFkFYA6iZBDTAA
EleZ2E74bAJXJjcbouE8eQOcyuP8hAlKIrTRjfgZmcndY1SHEGWfXn12nEC2x2YJ
LcSB1PHmy+texX9ayzzR1pPpvPKg852tEHcgTMDiUMMC4cCCtfJ+uHiKdqWiwsnP
nXPsCZuA8lqAGc70C9q9hQRrncyYIMTn+hc1o+lk9iTqfJoleg9RbE5EJ97OcV16
vNd+h1YOFrxM6NFtSeMNVQAVkEhRKkafWgs5/a8Pi2D3d/bwFq9KMLbebAwfYvYV
HPvE12k5a9nd52EJbnD/fYmmPuDuhX2YA+89tafzVEpe/D+cyqKt/nu6TM6T8HqM
soKCDeSzR9iWh3RIH+TPf5EhKH+JcOeZ5NdZ/bJIDJA=
`protect END_PROTECTED
