`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tw35aUdTdbnkwDB2IkNwzZmb//j6SWVt7A1JTVCTrdruIFEykQxIEyECpwyjmOU5
jgZP3hFUcvbtvHWNOKI9GX8KH2D92ecQ90BWMj5DaNWfV+YYOmnqm/VQXrk/UxSu
AbE9VvsWxIMu1ajKtEP/R3HCUTJxqCxM85EmuEwCTvZOz6OI4QJ3UXpAv645auWv
uaBoP2EC0gmDzrZCK20QrshOIsY/fLweiiOS2oOr0dclH2kakLLTSIUzk7T1D3mc
Sj56g9jZLYtvskdIzV5crcDE9YYljfVhygNBononQKwQ3o4wHBbRNGz7YnLHnql9
GAegRHNAN+BPR5+zgO5Yseuw66/ISJ4uVHo04taTQoiZhP7uFm8udzGYf034AA90
zuzcDIEkBEZKYj5Aj5fXNyHQcnZpUCu/YsPeQD5S/Rc=
`protect END_PROTECTED
