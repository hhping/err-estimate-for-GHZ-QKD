`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k3qcZ//8d5JALmdA5poy5/MILyUlov6voRgZWds739Dvi4gw8dLKGIsOZNeOyEsd
8DgrzrW62OB0+tYknS5bMLsBJthbB9sKsy5bxTx8wX4q4yf/20RD80n77guR7vkh
MBEFZAZYyt4+uAWBG3pWBNUJKcuiisGX4Eqfpv/K67xB/BQXOh1e/SHGT2oe/Vka
XHVOYu+IwYVjowgAeyLXZHHWjVgxxH3rZsYgOS42dpkq1eko5wSJMH6/etnT+8Al
FsF+nwXmzTOPoPWBCWPJQiFosbpvWIl7648DO/8ClAZKBkKsn1qeK4rUn68lW6cZ
s6a9xP1PcFcHxetSkvkfjEW/ts7PFH00CqbvgvGV8r+dtPR3ULWfSm7s0a+2+d8J
XKCfJjNN7iaUnOnMY0zXVYwKpBK7C7osJpT9qjvXEJxfQaEdIQNA5/qwsJGBJQ1H
AiVtFmWYZ4OO/Fgme3ULIIeFrCdK4YCzj+swdZ6dGG9jIe/BZRB8RcxWSDj1jmDB
HZQw+k7MMdbi3Ro6AF6hHXwMgkU6hmag3qepxafSd30PWS0t6w2V8/0F9WTN8LrO
m1MWP4tXgsL87YX/CYuF6g6RdlFz2UsDYCteS143w5QBS4njczRFkXNSp7tps16s
v90HfdeG44+bj1/pHjsuJtYNeiqrAZymlQt4CkbORGIp7fYLIrafb0JRAv7dFc0P
oM7+GZbTTAt51jnU+hbC7k3R3veP/u5MeqjDCGZbB3E23yRA9kyZphp5N3CCSfkW
Wr6IiIRwz2+0YtIkC2Q9biXEFaDgWC/S8MFL76yyy5GyhV31tdooW3NeJGPJrDlq
772jv9W949wWk74ylv7qLxkiO/FqJZu55aY7P6ML75djvnT7pybwYVUFaZ/f7vyA
0rIVooT2LBla0KrmfhR4FA==
`protect END_PROTECTED
