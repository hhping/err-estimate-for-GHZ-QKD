`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6jLZbJrm/E/SJ4cjuDhCDOsKix3Ix8RFuEWtrHppFpP+xG7vjMcjWHcsLqM3//fT
enCKvcad8Q2Zwr+ST7naKukLxjda4PWwrDqKLsCsYadqBAOh70e7qRiYU8alHE7l
c/jaFUDDF2lndANJrfk+HeVbyeTUVWnL1vKvDV0LWKE1gDoQYk7XePp8oElgzaXF
rFL0im7zjwoAZAbCLEKCu8ECtOPT1lQIgldAWNjLwecWfPMy3PfC7L9kK1dP+DBt
EMvQiD6ssFRAZRhKaMtI6gAbrKZMrE89Kb21E9ckhfj5Zq/XlPLyOuviWdZXRKD9
A9k6h//tZg/e6WFftNPnGOGUL4lojdd5Q56CBarJwvGbpSPNV3ZdZA11l/FBgJ1R
3XgMF9YA39g6FhX+XPcou/iYryN3A3Aok7183bCpJJho4jGSLwnA0W+AA0B8OBmJ
6MKvJG1FFITnqgpzin8YOCzEYxeB1KlqwH6oAg+2505J3bdyPL0GwMpyudSI+ZQL
LfWZjm2hirVbcDbjrGOcP+wSobviaSHMCmflufU4CZ2pqPvYVOkewgOq7q0Yjvcp
gs/UNdsLmmBMMGrIQPziP4T8uHs+eRRWw7VWtdDhadVwnxJFAPlO+Zl1yYf6OCDA
2gkC2AEc/Tp703dHF0jsP4e0FtrSUMI/NJQkpR6e7+V+YhamX1KOg019kbJ2SORV
zIX05kDNcb88Dy5xTvATJhWCF+9r56oQT7UlZ/WWv83T4jvv2GYwDFx8OvXhjXW5
FssjMWpfQcJKLEc9MNnjAFFjfVlwCFeMsOk5+/kQNkwBfLmQ/RvMnWOwNC1ZVZWL
Bf3A56dNNpXVLQVK7uTi/BSHylI6IT94qzxStvS4A58g/P8ujPvia5RVCVSRrWmk
qBOvyUCUf7hlvEtWjaR/zhdYgtdK/k77tQg/cDKFfrqFffYCOomgSc04XWBptHF/
1YWt+jQjwXXfcGNddVQtlA1JNZuynO+6W5RgvU7i8WBc8U1+ntD8CeUwsIyvfDK8
V0As6ZExonXTxS238Qc/u+m6IU/giMG6fh4C5rV8kQyS9NWkE1hj/kYeDPueqOtP
pKEmu3Snz36bGZefsFQZMp+FTHhTBOw8tQm48saWSMFscNMyewXHu4v2Wn4sDuJP
zzvl2tXPaK6u4kc9geTtME6iGPFiMCRoRyOEbbNqEZX/wG5FtoHCcQ515HxXG2Y3
lEw0hsWOgtdhB59FtyRMqxoTA3N5bnO63LzlXbpSiEnuZxMonR4a9WuRZ2A4YNd4
dsmhwdy2uC8Or1PJbnTUky/TwknltzZy09DiD97X5Lppfxniu87u4Pud25dRroQY
SBx97yPsAE/zEJg/kD7j/10fgWyqQdYTegc45Qzsvhh7ghogEGlR8kPvuRVCqGsU
q1bPJGrEmoUVGOl+YZciwnZYB1J9EJJuSwSpiel4jQkofXmMtzWEvQioKfPQmufH
TAMDx2DhIXPGrlP+h75zWTGFm4loCtBh5mK5F3grSyW3yagC8sbs+iHiQc/Nm4YT
weJ/xVtmaBLvKJ2ECyU1RVqlCgmJedFw8+o8lbehTxIehyhJAKf+BZnOS07etQGL
eSWL/tD8eXXId+S1PrPh4g==
`protect END_PROTECTED
