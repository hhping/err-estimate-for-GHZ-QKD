`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XvmbgbT6MaBf+3qxn0nq3f7ZrBJH6Go34vMgxvY8/KCfmycgYiJCsMG7hQeLs9+m
4Uxa+gXRznlk8Ytt4n8pH/653pw0QYL/GIpD23gLv15RQBPZxmplndzVWCPiUIUE
zfBwDGqXdx+2EIsILA2jHO0OClgfrVbx9Gg6qXgZH4PcSDp7jPGRNuypXfFhwgjR
9RaqTM3OdYbZv3nWRDtcbjQPOn0NVQAuQAEyMsO7O1hUtsexxYbcr5oQJkOTFkTQ
loCdG4+LYDjWcPS84zbdkJ/Ii/hGVJDmg3qRoxCOlsgqDVRPJS+9q7wDutT9QkAP
C/BpVre3tqIvvYP6kzcAdhZTEC/Qz7ANQtppZ2uZItMdM4G2OTzV+BP0aW8QXgWa
5D6ilv91CStucqPQCVxJCMBmnOTGNQdoJEaCZGu204Yqe3aT179Z9sAizn9hOAJ1
C2wkBg3wbdYcksoRcrUH9RphtFA9CSBiXVfM+F2P1sCtAiHMxz67iEQHcVEdTQLI
wOnVd18pyvIGGstYpHPZGw3dAC/oylbHLL/64GllrOZlXyE6WaMLl9glJyLHiS5h
2okdBqsCfi5NbAaIHIrF0luv3JP0cWdB7ifFy5FVLIS/DAFWUEd4X5grisiNQBri
/1DKW+2e8pSZlgFp+iysQ+o9NlEE58DDHoZ0CK1lRAIkkkadBaqza9E2MGn+Lvzu
4EfrDm5aLXFcAixiz7RRpTvQ8EYepyteg5TmYtSE8YzjC7L7J9i1gPtA6g3Z4Bpa
NOUG4L6kSIbKdUURWbiyc/BTa5hE1Qu7/MDv6NMs5k80r8J4ucaGPZ0Q6Z53UgFl
2tuXfYXXj1FhydMeIq9QUOj/5FSVIYdUF/EX0vK6LHrW5k75qygJf1rKOdfmqmd2
bBHxi4BZEFXNFNGaxlUXC4CLwD/Ewv4W/kX0rYE3gJfL+aOlLWN2Feq+qFDX1EuC
wzB2p90IE/zSkdXHRuHnHlMG5q7MIXXMrlxKcs8DZk5Gkm0+0+kEfxDqxBSvBq9K
fhEZ8H5a2Y9p25uK8EqjKroYOzEgw23dx5rRnAxTsAf0dzzlqwJJ9Ro/YTThbqiQ
LTIW5EzsBXxLTu6ShlTl6zj5YGxEznd2jv6MSUQG0pXZJMYHyBiHGfEt5w3gXVzK
HYkmIoZvtUvaFjkgQQ59j+AftfGABaqw3c0Fn4bGBYbALaqeAbHU4XgbonRcrSNg
vVPKFTb4bJZ53EwsLLoV0JuWLlZNEcSMXYrOg4Py56BWMBzrFsTHU3fxh3APwJc0
R4cwf7yxnZjajl04nenPyuKJcpFikgvnkhR4YSBM5qWqSoBsKCTp62mkpdn//Dar
JEUYyegyhUrrOVGlkCAkTRzeLBZ3TBKxm6edq06ig2RdyKYWSpOK2yzTyAQ1gBKr
g0PKYaWgK2ryHHNyk0YrIr1kgnNcvyKjqB66DohJUicmtAhf6iqEnmlduQLyBaXe
l7XjZS3dEwiNIXTDc/UFEA==
`protect END_PROTECTED
