`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VOaCUukHp11TQPS2Pp2cVj9JOZBE/00Ys1faEfal2gDLByHaUiiO5HX/S59lu0dx
y1NYlYLhyHsieRHg2wbqo3W1Bj/GlZduGxGO2CVeglYeOKlwLJkXHYiA6cV8z2hr
mJIFPQZ9LYj3FyaBjsY9O7UnHdHhW5PAlq40uZJ/POxzRtKRthb/gtlRDCG9OOHH
MgBwzQn7CqrNmzjG/T0qHZ6nduCosTO/HCDdGRXDm0jNFVV5auoxZxsGdTTx37gO
FxwdGO9NJg5QbyKjIDaPL1xKbXAe2v1i9+oVmg8aDY1gIjb4RaMm3Vy6U8BWWCVd
714RvCVnMWCcxb9oYExzt5uFuEMAucqav0+7OBVSkGRw3ZuTLfwuZ2fqsBl6ObnO
vyr6qmou7Fr6AhOaXZ5dyOCBXqKYBcTH0RmUmUdDJcKwyy0rwCTmbfzV3HroHzZC
af9Rlo1b9b86NoPwAMBDwmGL+bdT+wKUKpQYF3iGlzRvpOoSbxElasYCnScRtgiq
bPIkZPztwNQ8cGoSF5w0iSqYwX0jJEIDVR2fJDOsGjq9acUKCF2ZejnUeO7kd/Bs
kwm5c7H5TTpuLYh7mbm9TqLgi/S6/7M5l3ygoaKgTrU6Nr6Z4deHTIiMVG7qCLAh
E2qnKeuaYZ0388yZ4QvsBekRJaXzdYetcCqLEOu1tr11asCnf+zEiTIQ5tuOYazx
Zk7Fao40IhfznrauUaajRO63C7MKYH1krTgAxHkFuHZRjTYqJaX1p/4zQkmMPJYD
+lV13xGGm/usOCyd/M/hYZ78GcML+kLnfEF7wqm+0QBDWNdDTJ/HFtWrqEtrPZGS
DbQ/rNEKherjYIgpPr1Uf2gScuw/G9oUeMrVj5iCJpIXUZPl/ijN0iot4niwE4W1
iBY9lm0ODvFTZsOXeegB1qMB6lEmeYJCBCbkoLXp8ZV39J5CwRNLBw0A1GHJy3s4
oJHK5D921Eupv8ob7UVbLua3bjzsp0CRkxBr4lwbpKz1mtihqmtGUXLMRpyZI0wu
CU3GE1hOXUJhUg3H3xt/tQfth28BzvT9EyINhzvcr++3MYiGMc42CQjLfnrW5jam
tCPHNP90m6SRsAOiTqE6eeRFgxgbnnmKV+ipNo9g/dveMsYIsToHtEjJWNB5F1X3
CAgd9lhWLNR/Rq4s1/GMHnjFZq6TZF6sK1fx8oBv2Gz5aqQDgyeDNNZjNHwcsAOF
+qFszV+OZGZbq4fbGvu/ePThuE7jPSQ9wfzMgVl8vex+nNDs60tUxPe+UuYFOgFK
3QCA0WWWgTUNBxy7Rothm2OFSg7IFiQPCd82itl93afnjp/CleNVUpbysTtRwmCH
ctNY1e8v2hXUBB6W4t0xf0HmyZyjM6QT72yQ4pBCQc4BUNLUB2zTYZiIDok6+qsq
WbmwnQbVfZ/GBfh93FKA5K0svsdKk/z40MP2b3ASkjssjf4JUxrPsCQJ+O9yp7Ws
V36m3TJXa0vd5uQey4q22wGK98S54enczg7qkAMGfQ56my6tvPzXUdgFcRlCTCOn
Y2GpN7ALzNmUx1O/4exkbclihb6xknd19EwavLWTZG5S5I6o/uQ3f6C+DT9wnZXR
I6uTJsaamc9VZlHvM3HPh3d/Z9Lli8x8kMwUvLt4r9nZVxnfOmKrLQYVLTKFuDza
aV2wH05ogYBqQ8akGDR9HmOZn18KNzbhVJNIQ9gLaVojO0vYNU+kzfx+AHF6HL/8
srFOZPm3P97xQhq5ultNOOkfBdYWvrUps3avYs1HFM6Y2X2epiuus8LpP7O27CRL
Y6gAics+y6RCkekP3VW1sP7R+zFcbg9OrOCuF/KDOdMjo2T5KtKEXh8EikRLEUGR
yXw9mQN7k8f38wtDfFiZStZg3ruptfladTSuCCW7XdKIcNsEtZj7DP4T7pXJaDeq
A4isrlrfr9nxRJsRYsXOZ/v6kstVImBEI0cM2vPjtxF2Mw2H2+eN56/J83X7XJ41
EzCKr2yVfYjzgeX4efFmohyZ/uxEqzNCYgZXNyuVOEFEwNd8qIRiQZ0XDaT7stE7
g7HPchOGwkVl/CnE+quFzkwHwGRZHHsU7wv8P5jiKi95c3NdaBAyDDN1s1JY0kcA
BmrrU3Au05bD6XKU0prFHdQI+xc7AqqIdoAl3ly2EQ1Mpvqiz2kSNCASrtdVc4kt
igMNpo1mFQt2yTTgEvaHsJEf4FVlLkxZpxZGyfTko52gjibTPqX7tVkRuInu2BF3
2uHCkM/qyw+ogQfBU28RSAJGUDkJZyXroYOTW6IS8s3v1IqSkhOhtRHmZeHXC63f
TmqL4byAVU3yTkuNoAsO79vul/+VW80AoeAnKyO1q7sboHq/xO8EHaNsSsV18HqD
BSmx9xQWtDHwIjgSlRgBsegXWUE4DWpWzvlUZQGoUN/mDpsi1OCcVzSBblasRHIB
nasKbQ4kJZn5THKtxpN5gdoebr1Y9CRBkbYsTfuzNxLWnDNk7tjal5qu0gyI4ww9
X9pt80YBy9SJtupDiGUvmmry9B0avvYqNGDpbYHV0nHvB/kmwTnnVJfJBZrA/sOc
Aduj6AVQDoML87ur/9rlj8832GYyeF42zDw65tfHzxiu7J4a7s63tTatrkxRvWLA
kIae1FYtoHGh14LQ2W9bdYq1AcZ+ihjTHTL/u43+8sQEoKTGzvILsxbORhOpYUHA
IZhiGuRYajYDL4lcA+RUJSG6nVkjkhR08/MPbmvGCHpn4BpTpA3XJw26IfAipnmM
jj12vjaRJi9MDrNkK5ioQKYeHnBgh3Ys6vwMpbvag372B73AfFKU/5z4gsnYd81U
JSh4535PHTRlfq9r0vBdSRfZN92iPVXLj0FLG9jfkB4gnjhtLR8bS6j8/FbvXJZk
oGaeXKr/IV6yNEreFSJHVeB0Z4YLTMGFfOI49YolZ8ZwwLzAQZ5YOm0otlfqR2MG
ukiuX9R3C7XrMhPtOa5HduRECXl8ygvolJcIOm4HmWJ2W4jCmy5ohiVKPkbBZBe7
AdLiIBaLl6Ec7RJpfTb4CGZ8ZHGpqIwmPhkio7wCvk79wbrk8VMd2Q2u+0Z1vRVJ
SiYVOKL1DW4q++0e/jRIEhmFMkz95N66ERxei5ssc0Y7nqBtK60ltcZsL+xeEZZy
S++aRqH8UDSyJA/RC79RoNKT044IV86fQw2nFRAonUsZS8WOOhB7qiImu9u2TH8n
y5O/uzyVGH3H1Xuw8kcf3u6YxBZAaQKYm4JFXm7Qu+T1i67CwgvISq1s/zrS3vXc
vOhwyalEp6Wslz0vCK+7fR+DR+JE9WcKFXB5aV23MztJX3LrO7VG65zWMUGNLsNf
eSirVE7pk4IedmMqjtzYMWQ1G++1R5/WSnGovna1wx0rXSgjjBwLNr397GItPM+b
WayEUhUsTaD2m8LmNBKwGuoNvkZcyU4qbrnbEZWNcDRS6++fLiDM00hzenxAeoPS
+vgsuhG84WdI1UZMOmSZRAnwwFeTmcnQXlm/ChVHUlh69X5zJs9MY7VKnHt1CVGs
WaQNdcvSSyi2HMKpsxUZcjMfXaVhfW1POuyzU5HEt8Oc5tsbKe9NfpWZuwZL8jhi
IQFaQCMVOWRdvF7EncWKA5J6cCrp/SEtbq0J5fDwkJkuPJ9CFe17bEokhtd/siMC
hGymDFtOcRlhVO2aIjcW2FYKUEecHirUxu27fsJEQg2aTv1OCrKhb1Bj37y3zVvL
B8FHGbBExJBwljffT+hLWtRZvJV2+fyCUZZ86ivRHlLRELBjTIfZ1pkmY2LSi4Ja
GNhvskSvKYylg03a9ZdjFVcwfJK5wpVZ0q8L18Nj46foCR8uZMbwvZTjPxoYRb8w
PLL2eIEsTmjfmGDdqXrcjJj7arbUVVm3mlok2YF9XnyABsqGMP+Q8Hsx0HC8fX0A
dmZRRSvH/CMy3oLDl1Anu7+l9OGqz5Nz+Z4OnYzvH4SAx1ZtnmPEP7wTErl+3Bx1
R7ZOXIaStfRj+dnzwlPOWU2dpiFy5GpTxT44fLVR9S3d4imvnV4vnyoBtSTbLigH
FIQKswE/LjMvHSB+WXZozyhPbAnwgweL4asNWkWVoV10rGE+Qscoxzy+Mtass9Sq
msZUZRUD7pxGU0ZcZVSJoMeKS8qsjQ2ikFF4C1qOnd3HKeP4UzC9IWoocGEM/QLR
f02r39rxqjX1lvBOSxykDSnuVPzOGHjLVuCmLMW2ccWs7bmwJ19r2V/u79Pp8UnE
cgVtD+QaJziKmU+NdMp+4RuIeY9/q/R47IaWSCSfKJHTwGWBC2KmK8FVCvIvu1fH
A8OWAmT1a/WWHdwd1q6ofkBDejIMp0ByX23t3sa/Hslp/Qkfk3qF5FW4XVTdTir0
de2QnbmKbeKFetZckBGW5pZHQJVJ5K8xdA7+pn8TMAjOG8MiZEwqFxCyVEppaDp3
pFJcfAA2q205yAkNyE/13mctp5Glf/BINTWfYWHeo/NXGVw7Ui+UlBF540jhlppY
BGmSBZQUOEaqnSKl1YTAesXnGhNrzyYcvEmGNK7iN4mW/WsCRXeEO1FPSzZGOb54
Lvs7QvOMjBnBkj3HZWD9SOTwJvI0sMxFsYfJ4Nze0vbDADnWTjg76ZMduKGCb10j
SSHzvdOCyJqnCX51a998eXMV67HA6W/6vOMJzhzxp1o=
`protect END_PROTECTED
