`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xVbt58HVjy7Jm64KexisbtA87ytWrBC+lNAt1lrAiU3uGd8Vgh5TbgyGOXSqlN5N
lFfuNzIX0/v9ZfRnlHUDorjgM3I8h0CSlg0u4a586kfwL9wZ7tsX5sbU4CaHD9QM
dXbpeHP5Y0YvLpCaX/OXkUDB7BVwnym9/iXA7yKaGXfS9nh2tlQKMnYVM/hHomPN
8LkYS7I7xRAy4ie2chm1k0RJtuyNf0FUAu2TN5Mak54qUGf9tXSFB24TIH3HgfYa
L4jMXF1YDlNul/OSKS1BnqzktdJzhJG4WQb1y+zjICliaNOCd4zoVvywT3OyldgO
+POZOK/R0Gce47YNz4Cyf6fdl2hTurGkEUV1p7TmtghAS8lzSpDLVYGHiiyleaMQ
GuL+pemAX+/x/NqnKVYY1jWdnzXE19V/wYCqsA6T6vcpkizsyRn+AU4qyG8c2eB5
R9guQ/AQ0S7bpDaEVzdiUEF7cxk/JIuLFKH8S0HluAir26uqH4nEZSSzxPM8o60p
eDLxe4UketnNhVtnXMpeLzCLiB3bck8seN3Pr1V636P5lJtPOUj7QjuKiwlqaGaN
Si8BeY9/HYgHGoEQX+7RdyikdU0wu8yYzbKFfJ4rHSZciyr0NdcEZvCIVWO7SxyU
RHZrAcdOY9XA2YbW9JGSVO/f+zrYJ2Yz3lMwe0kJf8u2rVs3YuWLa7uP2tRdvBSL
DNaO9J/EJQbrxxl+QpiCQ+4BQvWLDw0Pb5GIMjXXasTzc6a7iidbL/J9gfu7LwCX
Gl+auZlrogbjSNQGbZNTjTpioh5BH2cGvKWK5jMRuuEh12fiyCqyIni/LovyR8Sw
EF/y5YYCAhPLG3D+q/fZCpgZFyNm0xsZDHz09IHzzMU=
`protect END_PROTECTED
