`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r/rfzDs/LmxyAPWqdVihzR/bkQ+PHwKtfmf8xbtXoIR2h2deOjmKtEuxfX+tMHSP
4hf3qOldfwla2WNcQ3lKVimkfJy00HRzHt1n72jXwSBqTjpxOR8/iAJUhrDF4HWC
NNIU8W+aUDc6V7hqNMztcd5qUdTXWgFHefDH21oMGoIiQQNtP4I/42IdwUHMad6m
2PXiWzbpOEPZeZdb9LZS6o25n49VK+XtYBMxr2Pgbm/xEiG/rIN8MakXLyVPV/mu
wAAc4p3Wk1NvpKBZTXAHo31wFcfh0kGTbrid1kzb0Hnx8W3Pur66ze+ZwevDwUFt
JOySBS0r4ARUt477jymv3lAk3bJrlMlOIHdVyv94DUfgiTWnTxoSk31EHws/PDO9
yzcl0HbPdu+WH4lBde2i86E96rkH5qBjP2r8/3NwVInujES5nQKOkfAk36HeNRSg
VU0bx8j/XEWhJwNsZA7CxhpG24oz89F1hHWavH5CQW5zbd3llFuw9++6Uewtjb2R
qlSUvOAL7nI1EUPRfVDLzd063OdhIqSHKgEgxwpZZ6+Hlx8aX7SsDvhWK5g3BsRC
O2biPL5h8ss5Cj7IwQHKb5do94bcmSTyepqHJT1of7fBBdOIq1fEpsUdfWD1xzew
Oxb0esyiFg9gBEP8qYZIVHkpnV+96UtlGBwmHsHbvuZhfxp9g8NzMyC8Z4Q5kvCY
eF2L2jpYlSjfXTl1Hf5YURzEK2ICRjEZM6g7ixIFyONGXF0eyJSB9uy17/4BpVTI
M8Dtr4V25G+aTgVUbPN6LpaifbwI+pnnAYgujPXt6kvCk3pxaUvDkqY83OQ471j+
aTOONKfkhLLEfH8gyywoLWxVnNaBBPUvjDp5qex35x+ySQQdE78ocrux4G0zXe5j
5/87fRulHYj2AS9EkUNvYuNSC/fKCllysTXjejyEqoPJv5MEGwAGkAOIFyMs9S6h
MoZpZDgOAfonDZyRaBS7/ujZU9FPtLhOssIq78Yu1p8WtNkB05K9ywOtcg6uRAiF
IhhizyRCFxbRCZTFKP3Sh9Ud4bzM/ekAiU+rCqXelnAD8OaYuhzaVhnTpTk3Y6ki
UISN4ZtrQdSv8sOpT5HpBBu0fGj+psDF1sc+U5ybsXr2lKqA9lA3fnWTX1Hq1KAV
HRFI31617EN7rkXCo1SgAu6oSxCggpMlkBub7qtK4B92X8a8BWHVeFZz7DQRExL0
YR8/McigXAfQzGf8/qRbXhMMF2SBvzn49jp8kPuW3wW1Mr0+DqJ8E3ULytf8T94/
MxeSaC8QG95eEiFa9V+q/S4gerVMsfwApHsbwhCXxRwENJB8cTTp4N2396nWCeJW
HG63jwgF9A0gg9APH63dFgDs4Y4Jn/DhGRk3FOAp1hD5DGcNeDqlD+4kxyNJUf7x
vfsSJh27j+ehbQibXcGSU1ZuHvJUbtMamFdeSUXUzwNidn9FWP/CnliT/iBrlncW
F6sKIo7GojGsLKmV8t3g3dZJEmdrC9eiuuy1zXQe12snfuknrDNzimQJj99YXrwz
5knVKRUQgUSxshW558CH2/7aCj0qzZ/ezej62y3yYzjE95AnxWDMP45I9KfHoR/j
VyCw+f/MIhC598r02g9F5ov9zn9QzLsgsisMrV/ulHW7S/Kw+IdJTtNdgCKPDH+9
ffi/vBiARLD4qEKQlpCu574QlDyEIQ3DaQOwnCSvkNRVwO8intXYJ0R2z1PmIWl+
/M/NU3LLcnZmnYXO6wmHxV10DdK6NqQI6aIYX+74hUMV3FASnUNd1a4ah+aLsCKO
JHeHPCm8RSMeHyQS7MAlydkBF+TniygDZ4Ljxv049CjkJj6UbESztwvNX/ymJAwf
B5284k/soQCeWHDAVCkLuu0ujkA5EeuDiIHCwpKKsSigh+uvIuFHYWSJy4DFI4dt
aTbJyVRQdhpIcR2NVs/IOut4pvh2jLTd7TPIib9djiSzMzEjDKahwVrFtHR8a7l/
CPldjmxt42VR32u7384ZhYMggjdPgyt2YPz3kb9zPlSZnXspS8EITaqppbxZsF4i
BW+3aXAj1IdJoL79z1CIKMT00wg1Uz6PUnjhajaH8VjBkwuwjoKOt/DRsT8djQWz
Hm5GJf5Q9dFTi1JX9vEIyGOssCTHJzn2N0Q/Umuvg7RZz/uSOLuj5BdG4RMqLC3y
T6ppKMWroBXYs5a5ZQU4El9xNjZfe9UH04/GZwnQeTeViASLtJviYW8ZV2sCJEhJ
6jvfEvi2bJN037Bvf6zx/2kejx0Ofjrjw4Ll2dKac8/WQVtcjP4JSjhN2ZA/i3W9
KVDhCSlgV2oML4ozgMvPhV4fM9uowCBG6jMnY7ml9Jr3uXIr95YdSVn9FFdeTU5p
bTwu/owb66c6kPRqb2reYVMYQrUWD+hjAmrGo74Vnctg5Da4sBOn8LTaM6PwFr68
VtWHTIl20yxfgd1VTQR0LpCD3YJPKN1XGkZrb+Wf+j6o4gSeX9Q/qAoRKyQKBvy0
0sW7n6IehXBlKN1a9yWgWaNFJfUFpgn+574fIkZme+BggPYcqN3LxlCixjNr8p49
egaLszb/D8su5dkpR3PjCtn9I69bHf1myxzmZWoVCQvU8+Gv909auHunLtWl+yBJ
gvETco0ATSsXnuy/EmR5KiS+a1k2uZxWdCmNJ0Yj9yxgrfaNqQt/Um4bznoHreCY
mkDnIXPzs1laNhhhYW9UG3GOfIpzmKruTXCNPwWnChYHauEAf58M2NBvR7rkBdVz
DHC3WppHJch+YveR0BJZhtruKvOCj2exJqnZdia8t5gca8jUtQHnxmYX/gf5/N66
Rx88epyR8xMLHnReLXNGQLd30j5H42JfMu0r6TtrHguzlutEAi5eCWPP6866OJ0R
uCkVt7m5atTi4qghHufh5xbxUOJhEp9wpuZqhN3PkOEkncwtvG+m0XIrDSNcrEPW
bDWIadUlfy7k4WJxrrSOVIrpnSyYcSHeiqbOERGqUgEJe3L+1dwZtqrkDnvgjVDa
bZGlBrYY8G2nd2HVPn7Jp8C5hL+cnL3cdyplKu1FiTAZdqoWPO053261xQQW8dVT
Ubxg7eGhFW0l9bYOVo9kOgdfaQ+f0nw/cCf25EtdcgJgol+QIDp7wabe0zES/Ks/
moXEnUSKr7oTwtQCt6Gof8wdpZAwMva7ZKQmGRx76++dfMPj9ow3tx6GPhX6EuV4
ZrIqtv7HPKKZCOiBLG6RZNT8Q2c0T0E4aXc/Vg2WmhlB1gm3Zq611drqvnUAkVYQ
FGzaeQ1w5njZ9tvDF7XfYi6Szav42PQw6qjybtg3LSO4sbr+F1tZ+9dtZTlZtFRE
kH//4QdiQ1sAKnc2N3xghUijjF3hlhBtOI1fjIrepr/lKtmRKE0/Nn673e1qgxOU
+hprJET/fjSTyrKd9dclxEnoUktWw4Ve/gHABJbp5mn0azKXclMBv9nzKBJIfC+3
5lvISTbJhWMFTY7dDm9s3/++O+6hmIQPDgOuT/Vybc5nlllOADIPgm7Oy+kmcXtv
o203yIK1VianKBL+qhoOTcunNl2F1m9OOA7nBTc5wdJcCRgPjiYCc0hrH8DKYVi0
11dABJdPAUbsmbkDxg5LM0AEFLG+TpjCaDM7vjjzdKMI1bwafRFheEpV04XqJde5
29tZ4pi6zQa/ijyC5Jyvr9vYvbiIB4UbGjkA+ozWDNyKkOuo4LvBo4jyMT0V+rDS
5ef+ooZHGxQq3YFRlIO0Nh8e9/U1KfJWVAL9gb/2ZPmShdUmm+CvEI3oq/xfa4o9
CNV/JahlAKo7mQo9q9/3FMh7M9RcUK280yE3KSAmG7exNuQM58qOjbyLElbHf4iq
s+OXRNvL6TUZGfKik7nkHZG1utbCHCbTXDVLkhDKCD+lRPQhoE+w8Dr5Oyg+T4ZK
U44QMLkpMNym/XKyK9AhMjxfDg/kvB59owOTIZHM3kSdn6nPoaO3IlyHzMO5ZPZS
iUSeUzAj9nrTWLhpflaHh/Jf0GFXa0y+rVJNu9QNP6kiBIPOrNQ9JZSyLZIRIcKM
Lhne/w4HyPZ2cuslhvGXdxmznA5O2sG6oopDsqPRNh2EwKXpRR07vbssWLB92RIb
W9gZaQtr/YIgJExF+wgyZHd0wptF7417B3yN+DDtCmIH9Hzgy8K58MZWKa6IzAXD
j8hetUnmVthqBEKBQkfhvKX1hqIysy1oJoLv0DuBwjsZmoxy0gUkFO2/PvhKbtbk
iR6pOOqVYW2zcyqjTtd2XpxKTlSzEoyYxGWK4WjMLm6cjWF2mfIvt2G2grYl+yY1
nSqYpDaJTlUZbDv/m1v/M/vY/9EiPDJMQW0Ike1m+mk6ui8jZ9rErzpY1+Nplbcg
HQDD/L8llBqyeVj452WtaKjNhTJMqnrI3J249V57MY75oyvNUdztTDdS1zlTK0yj
dZo42lpMYzzU+zRzwz2RVGDikI/SpWCaOUjJjfy5jMQRazW4KRRlrmJexFHBvzBX
mqa84OrBLMqj659LLIRTL/1lHqDA39afeNIyh6JrdiT2k2c3cHIEsa7GE0v/u+H/
M6Rx/R0OkD+jv2i30lU0DTeFXRCO62PqIvUCl4X/loFMyOPZFsu/AeRPAA0iStH7
nwkph+FiT4D9BtBrYc7LC3IboielPZnkyDStLo4Wnj4PIZzgLD8xriKehmHKRtbq
I3LsWYHGQlQGTSsD9KJGfjRtBC+I5rBYYTCXuL+QsoCcA7/+0n22M/QMTf4eGH1D
lWmoroAxdPolrG8bo/8WDMM5bGdjO63wv0kCCVSSdUiuZ5PvEtNXR9ZNKlKEjIEb
Tt5FfjedgcVuEXSBucdUbhpym90+sqgy2IimzVb9xFEyp92bFUxfi6CB6ULPGV+c
IDB14CGcKC2Z+Fnea0yJPgNAH/sGWsJtxubSEEu7BlVPX0Q6bioAhNOsjbl2OxsV
XPAu17o6Y02DbYUxptTTLA==
`protect END_PROTECTED
