`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/P4Fs4IwnBcdKV+r2gFvCSZ0nN07MPzLhupUrKnG/ae7dQn1B57HqOC5eeDo3NnX
fi99yRJLjEfkVHRC6eMJ7buUdpVQOzYoMx24QTU8WjU7CWMHTZ7Ol0fl3yD6ktt/
zn1OZWlEe5mNinn6loPj6lxbB/5OyLYtDFjm9JkZYwkpzgIri/HVWfogVY79Vmfp
XFJVX2gdGYMUFIw9TG/VxTwKifFwgxTd/7RZk63+lw169Y4BDq386qH2L/05V8+n
uWiX2iZFW+FCGXejZEvpBLcY1xiJIs0MSjVQFyIBz0DxfuaM49EzQ9zU6w2wLk3x
ZxMz75e8gv94xcbB4Q1fWNNX8S5uDGXX1vgQonn76G0HrwVlx4euMAkmjJPV66Ns
/aDkUNWTDycQ7jRMphiIS27T1OyANoVL6lI+Bw5Fs/89r79fH0DRNq55mLWOu8VX
BSbQOS/O3rllRUSQrPp8jIuQRDV275Q2fruos7hey0fsK9LROgBPbUGNdpCXjUTW
y0G6tnR+aAL9A46O5hegM9Mx2UV573kpT0xC7qfqpexVKvR4m8lQX2ZVwlqLh33Z
kFadz1orQogGzumTYmAneeoDmE9LE3eRB8hmq4zzqDkx03LcuFBLdnl4gQ6muZd+
yOOnkLlt5vF4m6v1cAxWBG1/LdapB5EEhoqqVNg0hVbtnMs7eo9CbB44Hrzrufkf
U9dwEdZAPARMyEcA7fb8bc8CUwh61+rbeEBJVnw1T/sQk2FQWjKuAZMNkMe2vPzi
WxRQkcHledIB5WsS4UVS0zFtSxGZJU1Nm6ZEUL49+v24svGgNFvRog3664uaewCG
DjKJDAYlbfwb+aOcrCI/9g==
`protect END_PROTECTED
