`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jLRSv3af+1AsVVXIAe96+jdW77P8fB5Gl/7UaU9MK1LS0u9+DzK16/VMcd5PfNWi
M7Y0HK7W8w1C3n63FaUBYFuASWMniRW6P4SPvZti1IYreJ2eJDItR6DdxuEai3OV
T6nFSVNzSkabFEnep/WoQ/0WaH3MeVTMeEl7UUE8aCuKaD1Os8qoeuSTgaKRCak4
XdVg1mQhjhrSmLqi6hJ/W/7ejmrFrUNsWjgMmu5aH2vO21buXDaog0MYGr+9hLQw
h+wFimG89lwZltdC2l3I52Sdeittv31r0akopWX/rxk++Jvtx7cd9Hz29wNWHzhu
XSoFQC8HjDKUYiODU2QWBHqGDW/RBImgykJ95iJvi+b1G+8gLqQBUapza8Lti3ul
jxtj5EcwxspsIXl5Wm5QX0L6782+g6owAQk7A44h+cAnZ+eKrDAbfnX6MmGLScdd
RSfyXyMYeVzvsIzbiYfVJ3OGKapnWSvwxLs8LOOrWnQ9ATvl5AHQC1CGD1YzPnKe
QnBwQAaE1wU5hch889oBrb0vkzsnunOnuOD5jA4iPShZQntJwwdjQJ5lFEAMgcnW
EymfOYyYBP2FEAKBGJNSUqoHO0taFZbqhKyftnwazTL/6O+gfAbQjymqAyB34aDy
KGsqAYGA90WRH5f8k+59Dg==
`protect END_PROTECTED
