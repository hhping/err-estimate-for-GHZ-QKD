`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RK840JHvJUS5Fmavq2eY7iWiqDJ8DDXRP9N5k67RCiA+DxWtPBHYNKnGrHep0eXy
V/ShLogD7YZVR0gQKSP0SNb2mUNJLIh8VvGevCR+AfwMqL1n8Vuh8qYsRTXIi8no
XT8EatuC4acC73f10lt/KqpNt8xrZEfbm56N5VE9MnDvKnadfGswYHzFLB9/XRhi
XneN6Lwwc/heNuwmiSOu1g+XTCRyZ9l0+cZ/Ph+KID3bjJQJ9g6LVhJ4xqocU2If
ZQKt9Lg2Xfj8JMNzvHhmUOZD6bSy73VCVtB6IZ1Kwq1FyMJ/ISQSDA5dbiB2JvnW
QzLy6DTAsy0k5urNUhFTIzR6c37bhYSpbSF8sdMXBqK1bg+lX9koKDt9ZkY4/Gr2
RBWW60k6n3xIxF3DcoDkl3CgHb7FxiRuZNVF5+PSiqb/ut1HwQ7hWpXzvKZ0pqHg
W/JgrTqqOifdZTgCo2qQ1RQBBDizRuEVlJbL2MzscIrbXimnTT+o4q11ORcDjYxg
E17Yv1mFnZ03AXAaGUxz6S+IABg82KHF7egGKgY17G+yGttnrujkyASiLUbzVSTw
jzQDvs2BumH2TxkD8hrKGOLgMJ4lg/FJb5XVFXWcfzEM8fSHNiUsWdY1ubwUIicG
4/A1wFKOAKEZWbQcHRATOVMhbFsxzHma1WQwFc8j3FrIUJzFmdrjsFwMq7njBrMI
`protect END_PROTECTED
