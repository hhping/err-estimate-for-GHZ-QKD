`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tFJipB+LyDoFbOtb2c3l2fUDLjvHb0Whrh8IUXwS1L89PoeHckvyjNU3bhvM/gA9
Vxl+yY3f5Oe9cF6AfoahLdTAT27PTVLlQT3oGXyM1g7VsGAaCPvP/ePVzqnC+gmJ
D5P4k7sMm7VIGHh6Jz5rIZOhSzOHWAEHVB0Tuo69P3LD+5Uwds62raD8dvo2ItuO
DqC1NtQLHTJS0p06mpF5RIry3WmsXFIMx9ZE/+6swuA0Ge68HnMZ4bpm+rMJ4k0l
H86C5BvZUFXy9I6n3TVFGAJnfDmmbVs36nFC8SZGRxsyY0yTWR2g5wk9rLrGCtbS
ZuF7jBiJn47pwgCBWss5+Hw34To7JDNJwjMNyCFWB519NQfXDdultRQL1Dz6h7a7
V6zpxmkLVkmLWzXyfezHF9M+LkMKOFpM27Ouhl6GSSBHssKkgtlLhQesqWo6plLG
hjbDjjQX2DGFzBW6IG7vRsgcryTSOEtrg3iDHw1ZdTRykgqgTqvgCj3AMvUN/g00
GZkIhadFDSQNSJSFBJnWs8CI1H4TugKOaMoe9zLNhlMjxTIENIRoxAIiiQf3sB8e
cUnTqPyN4jhfFZhqWX4uhiVVFUDoR84O0kD+mE0/KhmBT2t9nYGyEjWzpTrTeg+I
u81KuSxCl1xvtcO3O8nWXn7ylES9zhC1KoqJDNAGRsjEnZU7/GUl9xld3vURXMLD
uKAYhSvy6/1/lbuZq5fe/+fpq0X4NuP14l5SZ8/Y9+p6+S52uL5JwC1PNHNMqZY1
g5b1i8NJbZPRhWcEJLL+Q7uOm1cK5MLR/mmEhNSk58tggW5FE699WKydhHtx2Fuk
tC6z/qDRWPYlFIh4pPNMfPh5bN4VrUsaYnIvTysYOlFsClXvOpsTF0aMJDpd7kXq
6nD34sVL9zG9Zas70JepDo5vhH/jN0dKaKFCgdj/D44fPH0IJA/RiAVeOiQNZlH7
8qKnrMlQW/RrYIx5Cwa9SsY+ey9GHvReavHDq9X5sUVB88raFvQGyKrq+Zy1jYn6
g/1HxftZbIH+otxhESrDsKKAD7ugCSMPE+t5D3nSqvhjDQIbliCF/mRGmoB0LC1j
QKkddNaKc2trS2j7Ia+F1Jcd1NLCBp0CJB90WbF4UjEJ3r3G/xlhL0li0IOp9UGf
4t+Dm2rgCn4Dm/quEQbqsoiswa3vGFJyJ7UFuIiAe5e8pwhECNZda/HsQh9cQVLI
CBTxgORbMSkMoa+Y1VcSaechX4L+Xg/aPzVkDLqU4NmWbD9xm8NAKuQvM+FihotW
WFdGvgYXLO+UYsOJIegllT/RsgBKp3cW6s+0LvVhTLheZqRGHPToekcGw4etIdDN
Ic+Xsv1TDTbOZDWWjI9iMPkot/t6JKb8NpLhgw6NmmW5CVQglGpsbvalskPgAJIN
ue1qJk/jaTAgOpI/NEGgiU88QTJosbx/dBmqk+MfmkqoXUqa++7P/um2mkaHu7Rn
1deg1h86fDJpRUgaqr6jmW/HcYOjH4dExqDRPgBWLQsOSRtr45XylrgjKkcgvaIr
KJOmlXehIOSLXgqUp9f1QGRIdJALBrSATO0rV18tCldfrU6ipjqTr0izlSpHhf3J
zTjJfAv7WvA9SMp5qze02DyWIBuTxCn8eCcMUnLTgbrU+7xFJVz557L2Gu/Qhj7+
wGaGeQOP7BDjhkYfSKl11fGWJ4jo2pJnduL3YOtaL4HJPsFlzux6+RJEjYXMkaAH
FLQiqnCqLJ7vZojLt3DJs66YCgSPv5Q5C2oE6rPtrjpHX+QS//zedTdZFHkuOlfH
AYERxK+dbnyIrgsUUi+V26Mp+TXU0rNYLkh5PqrAZh48a2Zj3oWHdhPkrhZFw1b/
9SPRjaHffO1F+yVGqJIR0iwk2PLxJ7lZE9bH6/fc8wHyWetqT/nHuFT1vpuZsxpZ
ppJUg0ISBZFLOnPyKczPUOyh2Atf/JcxMTLsSpZ6h9M6jwnbl3EwVF2j0fo6U2mh
nwOk8EIx1hvjMxU5V87IdYxYMsKTGqqTGqB+VQZ8q8Nlab6BPJv5Hqp2lWkDbn8y
8srwM1821CM+HxB6NxFwmNK2N0dlS0POXWDWoJJkjbZ58auq2sKFO5refYH3PUkV
LnrL05ORMG7SpAbohP7+YID6EcUd1gKrX8mwNJegu+mu0SEq2hDWqF4nk2gC0d9J
8J7FIP4bMlWXE/k0ytTJD6WyQR3/I///cvjT5HlV/7sS+5/wV7PDLAyMdCoplq0f
kYLcrRt9yUeciLW8+tiwHNDlJYYDPMZGuOZFBdkPpYUdSEFYYbW+rKOmppTrNq1x
cFLymxXjoKhfmAY2NAk1E8fs6HjWdRRR+pjXumr3maU=
`protect END_PROTECTED
