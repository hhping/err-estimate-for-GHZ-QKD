`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
igbWWoqf0hIB6NUdXtFVy6O/aB9yN0Hu3sh3n+adMSJ2biIMPdnYN/DviPm7sjlJ
Kj2m43ejbmbrACdbLN2TH3Ma2K5NzWG1oz7uwbSVL1SpIbcPuuwsAwxcjlJYsofV
EfF7AtzJRplwbIRtFsWobSauWL8+cSUNmAfxcCcY6XI69JA+GyfJ5n56DJJSHN3F
40M0cdcFpNNVO9JsI3XULPo3xik6KCmn3mANlivJpQlDKGevh1S4e8dwtqdCobmZ
FODDEnazONFhIcjucqevEwedY/4nS3i4KIabO3a9xnAB+sRtsVjsk7+9RXhCnJJo
ynxqz2DTm3NOntNPnwwmWH7eegVvEk5ySmkAX/KEBFhe6qf3iqnKRBZxw9hAHeOr
NK9oUAEkkJZWrEAWrk6+UX7AO5ffeUA3/OUMcMMYmUAsYRiQvUohLTRDrcUktUFx
n3R6QeMozqc7174ULnGqcwAlWYSQJHIVPSjF5HEHvIVsyLKiOgJ3Kmj1H/1mfBMT
ns+67HVU1pANDUpfKKCDG22TPRsaNzFGfM8etzRlmd4/ilosKpI3GTeRs4QbsodO
L3fHip8LSkkz+BgTUzfIY/8AfFguDFDKdJnCHVzuzKaZ4noqzQNN2+bzOijIZz5t
CB2SH1nXr2PQ/e4WGj9Pkf/1LQ4Aq3tPOxFvyzo8VrDpDEcooUNqk8yBXYMdhsXM
6fb+YaRJP4hBQpAVz3Bb3PUb7DsDYntdaTMtZiMTBV9wBaLz35mr+osz/+f2UrJn
zeGDM3LMjoSF9um2wLzKc4JMZQVcX95WmoHHu6po1AP9KkudL9jHhRhlw2P0U8Wz
qkzJVntrJnF/zjd3QH6kCb/uSatHBp4dLCIf8zn07JWnQmcffmFUOlcdZQH9NvSJ
khWYIZDb/7nMhGlZjSWpNXEXyGRqksFf79YRD/9rKZmdU7arRrjDsbuvJPFuxU99
//5aMwGwRvKlxWcQhVuXhWq3jz/cGqm0a1WzrYr7oOAJqghaSDTPArZX2UKgzgnV
dmc2UezgwQn3455kWDL/RGNlBAuNPZYvkA1s11ziAqsaa+CNe2c6rLoA3iIzk5I9
lDfqyjjFnkLHlLCW28JHoe5VUkiEC4FKKAeMTPoqpBNOP8MhLY5HDQ8+4hwozJWj
0FGAEdlCn1VzZGlmUJKa6+s1c3VpORbcFufg43Wmv2IfZQ7CJKqUOjRy7byYQAnZ
FavS7VfUXdmkqsqTZhPQWxUmQaL97O8GZZRqlwtIkEsz1HHcp95e4yfTNpkNbLku
VxbQGn75sZFMdC3XSaz7EzA29XEIWBfSalC0VdpOX1ciqAyjB0QbSerYGm6hmk5n
2DXVtanCRgAWNxhQklR1+TI8Wj1n7fbNE6zESw4byT62COiKbQiEt5H9rk9usQnf
fsPrOKa+kbY4veCJ3griAW6/F78qUX55dmLyqYOVNuqxlde+8pagI3YNnXJAC6aY
7JLzQqyN8ZjmLmg/u5scxzy6sTW8XBXCQko/ighfumJqFBBsWAaBJ/HuqSNoH43+
/B89husXDjM0xGZRqUikYM8Zch7QdiZUeZ2vvCRMlXZKIjlOdfPV5IL6dDuxZRcu
/VR8MloJr6txDaLFK62mnPgDsBAaj58kwcNC+0Os/VJWecY5Zay0Yfb8qq7QIrOp
kIr9BToh+9alc5LM6f92LczPSSuG55XIp8sQxuUiWo/zvoh5IrlpCg4h1dLh3uEH
0gmRIscq7lwJYkEE8mQQAERw/yrBmNBX8UfOjYvcvq3/HaJip4wyJ0hitj0zWEot
kFeWutDdhgutQGLSk/An/KbHqNtidTND7eFPra2Dvogn5MuICUmBkYBcca/eBhCx
5wkN7iwGz6XOiY2DYmRcY3VEE7NGRVfyR2DraCxHWEV2KOjv/TsKOse2s3Dm30Sl
OBBQcWiMsxevLM2O8lD8L1D5gtR9KSLuUpuV3fGD3lJ+J3H/fgY4i9pTbjVyUl8t
dDBuui4HHzM0txzcfRaotN8y6KBED+T4b4Gbf3F+p7gjDsfoCsh3G9GbGK+qHP9/
eXAmhq3q3IKiegDX1aq7oW9XIdUdThnxvyzbm6V8QAGQXU5xd5IiGHvVCmKaqiDW
GsytfovghYHRFmhl+b1zSbxnaV0fp3LaReP6LC1P+5leORrlInEiJjo4Zzv1rEVH
c5N5zOPxNNChlovRlkD2vdjaUIixIfCg0JvKaAzF4CNp+VRpFQ0LCf+TdLLmBXFj
MER7MGSVk2LH81wHas+jH4iEIgg6Y5QDa+sOdtrwUZMdJ+4m6IQmdUdbRAfBUxE8
iiPukn4HIDtb3nAzr8e/Km6PvEgirqtxTDz6mbPg6XNIDw7bE2KYeJhSimS2msML
fk7Fv3CT3UjlQKyRrDCfFZQTqNn+YsKNZGU57qQ1tju+FKKVaTCPEeCak9RfEePC
65jS6QdoYrCWdxeF29uSrcp/MpeyixtnQj68Jmd+YMcBKWUgyhli8vckLyLCWN1/
9yt7hFoA4NVUKOnrKH1zYq0hV79tycPO8oEORPbElii/iXDmPA6SYxUERBbOgz1v
9oCYbHldUHYWw60CwasydmVyGNR8i3SAkvb0NhYvhKMiNCXdner5lkL9s4Pt5IHe
Yv+8AYKfXI2398u7uEMJbavFUgyOnAnDqrKDF0sYCrKgeJLebu1z3A6nNgV2Yj2F
/zqJsTx5rEwis03auBnw9cIdz4A2Tcvdax/+lv9nxiWiiPPpU002kSp/Annq4Xal
KhUwrTe23TusphWmm8zeQhuOdVi3ELKbnWbzk4XM/yK4braDAVUimT3RqNBKY8lS
kQtdrEsH/INwqX6QWOebX/6MG8zJvnvln6lG3Uf4d/Cvw92c2HIpPc6A+NJH1LYp
WgFGSAPbIG5Vc4KWZSfk3icOJyhBqx8YUA/2gkrvI225rTTQuyZ3CaTuzxUdJDyt
PXzt+k2UwGSbPBllNRlHv+M4ojPXYyDGqiukid1XOOrg73boErmwbytH4udExc2+
mVjxRRQhudf31AqJnw7yYNg7teGkLGWR4jLWuJWiYs+mcHSdk6Z+mP6NAMkrf4dC
6Zbj9rDq1EBe+PKUuORFve+Gd0heSkMZ0EkZM6mkGVWVp/eBj4tKStki4gKzcT33
yAXjRD0CNTDLlRGJXGOTJmOKy/Saf0UrlFyr8xDwaxkrINhUrU7FVlppAl1uSMv8
`protect END_PROTECTED
