`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b0QMl+D5oVZeIW4/8akXSpp0hD/yjnMXfRAaiaL6fJC+7/H9H2LdR0MHgQSC9sZf
CK/+xB4rbUSFL5BNEQyMjY7Ul6qnObXeYvDL1lsl3olPfy8iQbKmwzM+4YqV+F1u
kHynWF0lvE8mErYMXhNmjkeW/5rLlQIvUoZHOcPLLqIovx87yb3xyLtiQ8Ydfko6
4ldFEwnjTQhXqRWz6+laJTfBbuzgKGAktIeFKS4/OoHAa9TFeAcBlSvP6EaTGm3Z
Sh+3uBDCc/5JMtRcR5dK0/GWQ70sURjTsRAGrvkwjvJN4fSMN2Z20y1wX9SMAZuU
pcGpVDiLXSdWTODnOx98kB+wBJOpyBo0TERVNpCj3siIRddNBEgM9CEbn2MyOkvm
DUvf/mIcp5Orjf3Ca89qF0cnxf2kOCnvOPeotPqtfQHud2p7PqBNtzaqd2yQitjG
NqLAA/a+wXREj5Zj8s2XDGbFhzxXrzHCbGyUopL/qUgnBcsU7tZmUz7c9cA9isnw
LfVeV0MkKUSAriaHCVz8SV06ODoqtJyRtP6hEVrVAI/tsMxspa8AEM1DWCShGblK
16AxEftEPtofyqX7UaKwUE4Sb2alW0+8kGVgsb2cRYTT03hys0GTT/YH7EOFLa3s
uBQFqXVHgTrtJfkoOFVDbqFMedOD44fw2A9giUFL6ynylB2Ha5rZ/If8zvM1UR6O
D6jGza2bm08iJL+4elJ6gu/2+ngSegxDy1abJfSLe4sUxRFBV4rfNd3GrEJnhgIM
vuCpKZKmoRIKoGv9m6gK0WeGYOJhDiC959wH2d2gWOw4X7Cf3VU8u0IVHDbE42+6
0nS6TIW4lVstGmiZzthCRQsno8y0e63WY5uH37DpWBEV3JfS7MT3blvZuYp/+fSX
u654kTyMIyENZqulZvd0FCQBETuHIB2DFbplZmabpsZF5cbByrePGOdffLwkA2V9
4NtQ95hdLtVsETISDq9JNac6R8vrEQZ+jkdC0lwYy98mKFdG+bXWCcRKpaMvtsIK
LerPAAZ25taHyn2h8ycva5aDp+peRCy+bjDPRCuorHOmv8LQEQbmLJk3rosf6oSh
+EYTa0PCMY6avLVB7vafxwfcY2gqU5eVwmPH29twUo3lul1T38f1xqbDJ5HdlFR7
Xk/Vw5Q0IIoTC2VjjFAZMgTee3lI9rWDcoWOdc24aURzLxVCCooQjYYWG7nBMPeY
Sq4aPQfOedsopgWJXe8OlCG4lEhMsbWYN8hoWacHcgykXs1eTvfzcNy+COiwy28q
XNKDzu0MUoMq0u8w9Wp+0o3ENTGpgNuFhIFriLF/CGk=
`protect END_PROTECTED
