`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ReqNKgV7LRTU0dZYlqpgvvL967Ptf92ZXhA6BU/sErAdqbnCpibLqQ1tfj6j5Bfv
m3VehlDrlOx8A+yT3OxtaKh1tzcozL310lNawPgjn5oRIwCR+8cgHnW9gHH6bpVz
+568QZKIKislUbqaktWuwUKlPj07Ai56BkJur4qAUGgJE/D+loI+ZoLDuG9t2369
htOfE0CIlQnCXO6pV8/dyVa43Qua7wfln+G7PzBOkCrU4wFGkMzx+0ODVo3Kl4GD
XZWjuZze6qVMA6++fKXssAWFWV67//ICe+hPbraDHDqTPJkaJuzh+rRUyfwAjdbm
6EGJ8WvaBkqBYEG39PLw9ZcJF4SQPUaQ8zMW//fqzdK/pKTGI7g3ZHtws2+YllRh
orZYh9udXNns/VZ8r6kTG0PMKAYXeTOWajV1j8F3MY5MY4xXrWORh9QV7yNYSxDO
Sp3vU6mdo2LeUYfQg64gtQPssuaFP0ekGRQIMZCIscSTuo1vTljuGb6snVnC9oiT
0OcSQtICsuFaMVL4+Qh5K/ph+qccuobzRg4ulvspZqDQW3Cy6PtrviWLzFx7CNR4
WFKB9Cy/sBFJByYgY5g8Ya2Qol+AAuYqTnHm2B1lk0n+D/FVugxwXvUqhZwG0bBb
2cQF8ah0tHQhKthzragKisyCvvyHu7e4KlZreK7V6OzjL92GF9A+OH6d0//cOu5M
brQdFUONJcym9Nxgo6iUfvhCxGmoXJwpG//AWUnoyl/aMNVa3npEPxgauPCQwfdw
9tLL266SVBrzdWkjizJ1Cw8V5fsGk3KRXmacCO6R/CI=
`protect END_PROTECTED
