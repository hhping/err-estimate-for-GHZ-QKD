`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K6px1x2MCnV6Di36/jU2MiQ4GLW7+wIJm8stdeAFc/W7neWvx+qbTiz234OBKpGT
e+5SR2HSAn6T/nzm/PnnHicmiDvCMtb7qzSCWJJXFSAo9xPbzr0IulfJxideYbr+
Pg4JI/rdfeBSTzJs9nwBFSalGSkpkxuzkoMNQQMz8E2zQy0a2kvpb/sGtLI1anAN
WHUCdHBlRaM2TMmrDYXeanzWRjdWx+P7uWy0J7ZVnvfM4Hn5sYkAwMlfYtcQl9w7
yw8KfI+YKwY2oX5pyKiUG62umxa0KnHKZgESnpteGjRz/eBQduAXReeeTyt6Imnk
/ro8E/uw+RhR8csmBkP4/OjNPv4fKtBFgy85dK4CLsm6wMS0L2pdJ45cLYg9lETI
+jWjLhuDhRWbP03wxNrZ+M8O/MYkjlDsd5qb06txZbTgf5h6kx5VNtZN+Ph6gwA1
gEjSrCU+0V6gdXYBCgV3hdstQGxCnR//atFiOLRrikbxQNSHWNIenss0qtaFznN5
taHCaSBf/GTbt15WZzcFaeLL1rU0RjUF0PTLCFUKyu+jVlj6MLwOEzAErdg70QxP
zG/HDPO6meDc0RbP1xoerzeQbJb8yazP7ZtQd3aYJ6xaTeGQlJMAcw5fyzY+YFib
P4sOLN9foI/DvesNGqiwLDJ6hC6iGAzZK3z+7EOuS0iYTsrsbLqykMAM27uB5gJS
DQF1UInCAeli1VndJCWyCw==
`protect END_PROTECTED
