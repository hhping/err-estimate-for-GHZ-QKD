`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DbwVBmsf765iadngNJcu1UESV9XRtJSWXJdiK9B7lF+jzASkHcExSXrDJQUSSPpd
2Kr79fsoR+z6m9sgHkv5S9ecHclYUGptyuIfGydAcQxQEpW88HMNXNU62IMjI6td
LZeG1D+R3Y/CFX20HKAL8WByJhEfmUlsOc2FY0Ri5GNO60YkDObwFp9rGo2kJ27w
dPq0UfJ1DcZjdzNe0mkoy457HfcCF7esdHOklvYaIH/nrp0XSSMjGlq/s2UrO5XH
wrKQzSKQ6Wckzcc48atAE39JLWTycd5wx0tCLwz8XgFh5o/aCBusJhYNkCxW9eXe
J6CJtDwD+BcHbTTUGVojkbvxdW8C9oB2y4xw69cMJKPW9LVx2rOgTk9ahX91rR4T
8Puy6si8kkri8rc82MC390wWRT2a4O39p37zuuaLLNCIbRnpsapcEdUBx8k1oH8e
W0mvgRYKGpaOzFMcWgc5kyArs0+Alo9TAwDB6myvsGYFinth0gXziixSHszxom3d
rjUuN67gLpG7qz2w6kcisBi+Vsb/32eEJEmbxa3XPhfv/O98j9HDrisZBA0GOvDw
goghYdj78BTyz+vxXhcMH/NR9LhEWfYldGDRRXycIcBb8eymsg9fLXaQfK/GkLFR
CPkGE6Er6V8lsQMpVMrwO95dzsrlrRIZPi9fE+arDZ2gzqpTagnUIQ7wrwNnC2Wo
l1CCAurSOIlYx86ZiSwcsoHUJYCOwrtihsIZRyDs5eYJMZEa3ngERCx6wQO1wUy1
Ql0uVJLBustTUppHc6s2kroV+FiPfsmDxrVeI/d3VjMs2JxHt2SJy0oEdXa03szU
ZId/famQ4pxtoHuQSoJq8fNxufirlcM1an4fPp52komya0yqlNGwPVoEl6u2kYDe
3330ONAm67+ccgaXxTEVIGw9ea3O972GcmVFaI0batep93hhYLCOdhW+u1ysapXX
TD/Bye1Bu3Uk97wQu3N/S7ZlFWYsVDGdLWPaVmPZTQAxtASptSW2Apgn4T2dQlJz
s8ssRxWGCYMGXPvmRE7ybqyjuTAJqBzeWG5rV3TX/fTC0aXOFzbGqznLJvZnN5mj
OWObFpUG8Rzy4vaTQBToFFJzHvMG0M5cQ3M+SVgux1U6Lay4+954T/V+1i7gDll5
V5/Vtp3EFzyymAUAL1idkLQHk6zGjUeyyMntraDLx8HCCqJqT5/yUZHu+SiPq4vX
jsAo+Qu8VOsU1X2R69oeDHU6/84vLM3nR3tPjikb+Ymy5KUmuBruX1Pc/IY4i00T
ABDMTGzzzgiVx0vkmle1JBssxFfebidk6Wt4w3wkgPLLN2cdmGEQDv7rtB7MIPbs
utaaizKzJvxSFjDcbdHOnQC8mUQABaxPYAra9gl6Fy/MzAKlkwdJoRfBROKN8DtP
oreq2513H9eoqPeDa5ef3iCKwOWETfWWcE8R2c7KuVN5KlW3uOH9ISQFtDbmYkTw
P4hosZpd0aqh1Ly9g2bJz+Jw6HyvbScrXArlLC+8irlpaKrt3It/lIQkLF7D2vBx
co1TcnTlt0CoZBtYyBVxIfHQoBDQdsTgwsHZmbjLBr2EE3mpN1WdbEUq1y2STPCj
VM0/XWL8ls8R+jPiw4EPsg1GQ+VtVlPa2Yn7BsgxM7dDyvXJQk7Bh+d6wn0tgUNg
hK2LQqvc4T6V5jrGPvpu8+o0iInF9xaj6ZMilVzLYdg=
`protect END_PROTECTED
