`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rVZcwMEwjsl7I8TRzkMvOyiQKJan8uvsVBtGptmzKmTNvszuORuW5o3JpLpSRjmc
McI2Vsdf+fWWi2p8GHgcmA1vwhSIcw6YssR2jrKpUB2I3iW4fS8w3JZKw0QEiiR3
jSZCN7HQrgeDAGLcp/S2HJez9uLKJcn04/7e5HRYzBr36Xbd4N9BbPwqMZfIrGui
g/NEUw3GpgTFtUOsQTwj1zXhatoYm2ZsXAnAmbOjoTOWuEbmXm5zi0gkR06qy9hs
4U6KlaEeuvGOpJCApfAgq2OwvC9XKhnytumWfuu/q44Xp7shYpiH5JkT8vkRZr3M
TbaFIO64MbNqts3S9yzPz0KejRw/2olUh4cMoc/Kgrs9Xg4r8/fTh98BXxkgWNO0
fegdG6KqzV2jD7aVKdYV0xNHtuKu9rUtnnhcWEkXoKCPdpgEbLoRvjqTtLvIEBdQ
NTi5cHq73yfdqrLFvT1OWXys29mp1bHfGwRo6ZT1PQp6KMFK7foQRydjA/MMZZjp
Gsa2ByrFwronmHYmnfIxPS18zImccmMGEOZI2HFqNsMkGOJXQS7+RVyNDI5WMghf
tiIF/Ysc/nwrXjarl+CdH1gQW0Jj8uD8qqlp0gOS3/UbLeReaecwfTP6J8w3Vz1N
lmXuLjx7CC8G0p7IGu96+j2l3LOStD299jJSsNbblAaJzdxBdUiJJtcjMzlWKn+M
Lf/7STSVwU7UZc5iW922hdZuSSpT+qy/jeiSqnzQ8642Oqj4pm2Pny75OSuwbAiR
GaphgOc9CLu0rphdSjG4sWHRLzoA4t0YL5bNOjrHcfDg7GqOVUxzLwGIfWgQ4v1d
X18CT+TnpIehtA4Ewf/9mkUTEA1YSrsLUXCkERGItJX8UFUi9cEeRE/mafUm5+mN
DYNI6O2JsOI4Blvdg1HGQ+2l8/2c0FsolAeZ9cXw5EydKbeV1QeFU2m2p/CkshUg
lYtIbZ3MYiOSki4oeOH9Fa/DZrMJYWqKjg1C7pOU4GQL1Lp88U1/Do5dq1NBpNNq
33/uuGOm9jATHbtjcZBqHyUbOFR+WlQD6E22iMTlEP+mmpGyYfrVP45xFZhJa0aX
c9YmN5ZqOIZhVbRtjTaDW3ZkVMECKYKyRI4EYGyw/EwDuhpyfZi7RIWVKw9pXsB0
snN+qL3Q/p39cxPscIKLqpxqMRJh00RBteYfbGDym/c353KjMbFrBhhx9Eh1NIMd
RF92n+LftAx9gl4gfFjVcn6Ef6fv6mkrFghcGGci7IzC4DSQHb/NxYMcHeiGkYIY
1FGmn8AaxNE5wIVxS7LmfAtYNC/E/pDOiS4xiTjEHcFf+J4wubOb4Wh2N+tOcsGg
jZvh+X94LJeQHlrEhQscnCjKWpL914jspbZjSujVljA61/42tzW8+ndWlcgwWZ+0
NBxKcDjndiUcPko/m5WE5qEvzlb5rK+sACDRpWsEAeM5YDnCB7SLztLQhw5ybKAF
DdkFjShO9VkxZOJCTOelCrBc2sC58BVnkI+xFNfr+ngixLrgEj4KpJinaPHp6+VD
NPjyJaEjOswx1hinp4c31DlRj+rgQF+IxY9+ubjJuWdkpVILkOI0sS5VxLge9fX2
1k1UXndCfLIovT4ZUU0T++uQ3lq393yYjqHjbeK4XdpSdHwYIQr2p+S/8YsnEyjS
r/w/R3BESiEFfC7vrxMHUxmiNabJTfoFj9TKbWDsSmUSuEvg2zv52+oZkGHk0+Bf
gPOJeCA7+vjs1fxUX2IkJTvZjuWnQ4AbJdv05EITD+U76qdgDPceRD/TMtM1MbIR
FmZ3qlpMEIxWKrMbt0NbT5tXgULqRsdHgkJQIvTWt+jvFj+FP+v3p/GaVO3ubLYk
ljIl2iQYOpAaWHbFjdC5N0ONXA4X15yE5SICS099tvNku/Ghxch3BR+bqYrWnGac
jRGduMuL98TdMGE5EEfz4RWWBD51cqA96VLbhApRzYdglfjWedx5JiieEukyz39I
0XnV+E6qIKyT/wCHw1+zR+jVLPWU3hv8VO/TalBQZuKg5oAfKl/WEra5DKCoCDXq
811Hnmzp6sWefrY9EyjYnTrz+48rqcp500Ym8DJyHJTcfzADt252ObZ54JbfOjVD
SSeT3jULCNw0KJUSFaOSGt2j/4pxFC+2u1IDK/yW+R0=
`protect END_PROTECTED
