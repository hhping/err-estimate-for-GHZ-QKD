`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M2s9DUm3TOk4tUYnAOedxUjz6vAoeHRxbrdKvcx3YedVirMySUyn1In3VF4TYBbH
aVOKbXlmBQwtem58Ye2ZsdZl4UDmg8xh0d+/WLvObhKW4rEU4BemFbsP+HuonJGy
ZHvSY59ls8yYGXOv3KhoHeNN3muveTzyAA/FbRlJfd9hoMli4Paiuu1FTVbezUYJ
FPsX1SsO5c5aFFy2Aj3VQ5mwUIN2CPp9kDJtrvpJRpOhDVI8lKUo8BdtRJ/ClYzq
Q0HAT3k0vXcpBuDbR1vSZAdndcDAxNhH1c1dGjpkqhJL+EDcwWf88HwTPPqsHMMN
9tQbvkXm5APABLfpNBn3pgdlZyJHAUiwUMTEVq+pNdZ86GSCekAl3A4RmeJQnnuk
zYotmBgSU8AuEnCQ2Fjwp8tTJk2LxyPcBEUEy4O5U1R6DVGmGS1ha0Snluvh9d2U
L0PTz/9bJC6SBbJNELUHn1IENubw6qi+0l3kZoe77CpqDjskwyQrOgSrSQmCHK/h
TznvMUx3yXL+ne4IIrOAdgeId/l9LZ9eUFAWLqWdkaBPHmUEAKy7SfOVFkeYhaM8
U2vj/MBOJV9ZfmCfCYx3IGNXSVz2/nlJ7N49KSsKktnP7bN6TmqCHXxaJR7KFR8Y
aHBbAPAeORNABtCh/LzYIHCXmtheNMGliZT2DbGynC72/nKxIjEmkQzeb41vvbka
65aRz5y1HXA/zOMT+5VTPHj84gostU04bKHCKFWwtfdtx/VhRmk/SWCZZHSSS117
4ee2KxcRy5oveJTeDzBpiOY8vzNaAknqhoQ1LSVhtFlZMZtT0g61qRjL2Qf2tkPc
ExKTZJbeZTMwv0TKn9qFDbvUE0/lwVjH7FlM/HzAYMgs4V6T1JlEvYi8SfFt2oDY
KFU2iSGHRDRdN+Qkk6GPgQ5q+BLtJrQnxVluYNJxYSmWTf3dcOS9J1Ap4wzDwhGN
NzY9em0rliVaWyrwUDpB8AWaPtdqFD8g8ZZ5TwNPQeRarB2UmINpyaj0IuO381/o
E1NDJeCykTD7ND8jApZhIeO98WHmAGQNe/XwY9F2eBgaHt2DZfCKYr4gBqXiJZVQ
lbzWHFF+mnshDiQ2cFNlHoFhHIn9xed/A+sbjOxLW/e0avuBM+03f97a8X0HhFgh
v5PWmEjrVE90T1ZSh9IEZZsVCjGlAK5VhOdhkLuohM9LAUmACMz0YJDcleSTvDPT
6MDtuA+Cc42TO5jhHBJzbZhR3w4jtnDW4c2kFSLnJJx6vZyUNGHS+eG66wiDyQvF
OH2Hvqkk5Ca2XUHx1iZUEbYnDmdhPf6JpkMTW1GoK8HVKNeMrypunMcNOpmQ/vnD
+W4Yd37HluyPfl76imhEOk6qJiBO+BYnEtxBBVeRmPY=
`protect END_PROTECTED
