`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vwnb/h4Zv1HyLRfFMyArYkdOe93LnWEA5p1G73rzktCyl7HzYnBHrCuSEA1VLQ94
NvY6xCLx9lq66gM0xF72l+IpmeyyfeiriF1FdU21RsSDbiQqIEZRMmBMUBJs3I+Z
gFJZkyVHgxQ3T9ABdt+V7xoiMh5DsbyKlSgED6lXIZweCgaeqZA+LfJX8sA9THbs
OCYmXW89ByKu/5GH6xM7tji222KRs7haKYwJPB9zMqO9bwJCnz9kGGsXdF7/5f0d
rFUlC81pC7ZWBuI+ZhwvZd7qSJlW/z8VHby77Zjtd1SSF7zMAxiNy14bm1I1EBdm
WtklHp+1e3lQeRIzcDhmzAPuoaFHHbRZX3DirPY/OnrR1GnDx/I4eKuqJW71x0Fn
Q0Mq84mTe0p2iHAOBchrBZSxvjDP6hJ9iSWu3btns0jeA5TobODYeFCgg0WlTiYE
ZCKQO6c7VYYrkuH3u5KZsf8+2SVpwUC7N2OfNuJD3nVjri0YTxfIfKMKE5EO0R7L
16GdFZ1miX5Rye10jAgNuhzKZDEO3/AUnjZ6xc0DWsKCKI3qa07M5pRuLdLIIpl/
+lC7ebbtPZyJNXK98eAbdMOW57z9kmpKB2Kg6fFZCTdRgQYZAangCcn+wYUtuagT
SKLPNpWFGT3xR+R8EZlYeuxdSGo6jv6Rjt/zS9HX6VzYDL6c8qbfVdhUvqXJK9IN
/vbj4kAKUL82d8nqseG4HFRfgH1Mh9tuZoEYzSnrfQ1mmhBMJ12NAR+uV4LUpKIY
558F24we/53wp0f98WgLU0LGwgG0moguv6YcgPeqDuOnQMVVhJQvDkvXvtuh0z7j
OuF+uEz0nmZg/sf4ZmfRFYSilxoYAaAmL9A7DLovmbYLgKHyNfnIWMhKEM+RK8Ia
EYPLtuof1JGbJClQWuyz23WEjhgX3TKqhEUEhrJyR48WKegJhcisVPEZBLr67Ms2
nvc3s1lPyGN045qB3WOAAz+I9Jguf6BluDGgv4OOZfBHwDvXuNb/1AFkq5Jlvh6w
nZTw6Ayzzv/wsmtQWKo1Xjh0hNnb+gzqP3/wEpoOV6DnadjM6xbEgVsjFjJ+ZLFw
xOy69pEKlD3hJ+TwPggH3nY9kOt0QohtavtNhW3cexfKuHNLvXXGS/HcD9qG3bGg
3Tk429QxOLlzUOIiyL5wDS1z+OCqnm0eTEHnCrvG467VF3Cgvun9DWSyLnBARA+t
6KLrKGfGZSBhcUtZXHrwFeFj0/njjBoRb2Np94Vg5gp71TwVjXwR6i4IK277B/zu
nvv5f+mAD2tCC7lVTumaJQa6Os9fc2Twu8ByCPYtj8wNcbcqAVps9ZgdAMQmbbjm
kMtSQNyqRYNlRtwJon2kFsGnHefqt4Gkqrn75ej/XzIASlLuLq7BufL8RV/ZCOJt
tdozcOhOHCGS+rHFidMIYP9/4VY8GMoZiDxV2cxIcBpKddLRumr8AQzWkXSe7ndc
8b2hAY8zB8fqLdGuiKPMomc20s8a8Zm5kJVb6HARNEZajq9LVuu1tRjqdbM8IZtk
PJb2XJnskcQJBo2GZQHzaa4+Fxa+cPlU4zmt6HQzRGUR57U9xF0kVgyzmlvzXBdL
OvHBfbS0wcJaqxHr4l6e0t76v9Muu4/LFOA382xnPJNXtVDrEIP85BovrySfRplt
32QukuZZ+mM9cqqlw0A6gV98WWrOSHZhFXVtwANYtKAu6bpdYPxOGK14bu4vWHiG
tF9yF9gA0Ldj/WbyI3VSIdTC4dirMm9gxin7OTCyI/bBAHbzhFVf7HKhNxtom3/g
jtTF799QJXwIoZADACsxev3sxTwyBteHp1tAIh0pCBQJNKnmfPiPPfLTOr/GmOuD
oLTlmZgP2bjfvvmFIXrwcgH1fnVXFnjwHMM64PVDDiub0yghvOr5WhXPrYqYIWwK
JxrKJbdulwi1LuGIAQjMOQLA/Z1uVe2lDMyKtToRCJmGzDL2jAZEOK9dbGJ31y27
9Hm2ScDMl/FfJvNrdbjidcXWVj7njQA5tw9rUIXKU5jkEPm5RYBx0TpeYruq1YOE
GscuGykrN3Xf6bw+NORS+9A8sW7bm1ejVxpzCGx0cLsVAyfGFWCbQK4EGEUY11Tu
GBRZvCn+0LEOZ8errHmbKYk2eQ81eDJvZL2qmHdezYbh+tSVrVq40ZKNL/Lf30gW
`protect END_PROTECTED
