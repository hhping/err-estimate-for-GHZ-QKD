`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OdVzbxokRNRfpGq9MHFn9ZHhbNAZINJ0/bunQhwBLklSzY3lgz1Lu3tux2s7f8eR
yjJjlGnFkaFpkGplNurexAhg7WD8IQ4gvDMOWP8sis6+GSYmKXQCV7vGJoUmXy5u
S9pOkf5ILxjRWq1XovgaV8Y7UrupsKfPVm7qQHh1mm4ynT9QnjVDuCDYEn28UdBC
02CLfdi3iCy++CdSKXiOeg9/ncP5iUlUPXJUEOHN/3+7GvCdf0itQyGceyjnwD2H
ZD2n4/kUlIGYIAuZsEkMANIVe2HwcOpOaQjXhloQktvIWP7fbdixn9Kg8mFzY1F2
W4tzGB4/aHtXkdFdVmsZSWBoXhi9SVPeynqd1IEN6U0r51iCOi/PTTYKQVsF0CZ4
98xHWtTC6W2tFFJ2C5k/BWUG2cQCKC2EklIfoKiKezxRxORV8kFhTIYIqIO2nX/V
pRkeh7AJ8cZM6dYNBAnRnHIsu9MsjJCqfChzyqYszVHtVOSnrgiNNjLfKWrnamRS
Zol6OteSrUX+A2cNNmPBgkXXBgA5rKxHbtgC9MOFXtmKEs6Xrf1LmP29HaTjdNXg
GG8A+Or45W3EZRbVtX3QIIMlksvGzIdDqv7TPPHprJzW51BfvafOzh+ij3KHdeU9
TkuWrITojQEn0fiGtMq3zAHocnlBAurVtbCSgkiddoMItFOcw7CX23Byd5Tw0R3E
e7DS6myvEiEUPe8cI5OAVrF+OTvQI+XBEmCv28wtahU=
`protect END_PROTECTED
