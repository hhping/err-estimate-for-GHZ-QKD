`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9UTnK5qS35iroU2dv/TshW3Dw0eNxTOt8XXUpIJ3hXQYRUXjgV2sDCPHEwm2dr1q
YdcvEcnZ0DQD6NSp97bXIEF6gRT3KXYZPSq9Zc/KWFNfXQ4pSQapFt8jf0xdo0DJ
SuhUVECHJnlNllVle92EBfRZsJwu2uwHGe+e1UBJkX3dopVbonp73+ResnVm1jbX
0ZtbIOSxbbEu/cfmOW9FiXwzO7zkE7CCm6dEYp4Xw5Et1Kw6k0/WIajouIC0qlTQ
V3OeKv9gPhwxiZZPyQxS2x1pMxURWz+NEadPCpzBQ15o454yjbJIQR4xaRsiVH55
4WKB1rZjdie1R4VbCzYDMTUsfk7n+1mxIOv4e+jj8pN2YJbujzUlGUsljRVhb/g/
gI1BTbyrudmZIXSLyvO00VRJZWHsdt2dopYovwGHjBrCXkMBMxFb9p6ud/1UsU8+
OAxJ3tdhFP0txQFTwh4hPebrKemYQCUQplp6TiGtaQ9kmvhGCE6t7RB/8WGMbb/U
cKQmhXPVDqloFjxsPpwcN8uBvA9z5Hhh12EWOJxeVlGZQg1EMRi36T2pWqpFjnTl
VMaB6tqBCaMikNkAmPtgAE19E8+STaJI+fhhbhieGe4MRDHLsl69EmD9i2OzBf6P
XKlFfC/fOMQgDbA7NZUmSIv08Dm7g7FTJlBTKpolj+kz+TV6D0GTupS35MZYplvO
Z6KvPY4uzmPJ+/pGxjsq7/Fv6hcG+n8hy7PfP0ceizd6sAPX3UU5zaEvA4/llCoZ
z+zb0JeOGbazYkHGvoPcL6TAz4gvtvZynHPAhTR9RFIcGAOoTYk3TWLFb9kipTi7
Jy3g8beLeRvYK8bRPVq2+gjz4yFtFGUMgODS1Z+nCCdOyDgc+3M/MLUsoJ0AI5Bf
THiIrLUwDhqJzXfte62xrg==
`protect END_PROTECTED
