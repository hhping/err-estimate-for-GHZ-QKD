`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rzlDrg0e3NDMSELox5dE+sDZHRSMFaDvGevBYTcMP42eMcbgoRsV83WCFPGc0FmS
wN7srBresrsTOcjKtvsouDtdncfnpIfFjvTl/RVJYynoU8XRsRDVu8b4NMOgWJf8
i5ZSEc6TKWxXaLBhk1mgcuUI/N5cqvQNjR28zzdWeGZV2ZjSgl0YPECg/5+xxFgc
17duxb2HPfLeEkW2lVVA05T1lJVVFMO3wKPSBqpJ0kVv8JwN81Tvj4jzZEjZ5AOJ
3eBA1rOqVAlGPsnB7LhDvkZPFLq8t+E7iuzqvcW4rVuAoZfIVBi2gde6Y7VdaHYc
4/BZjq4okDZG97wgd5aaE02MtYZn1hdtSVxSjUEMqotYGcZvJpMDzXcK9XY136um
g3fkT0ulbDjRHzEfOntEWDj3HuYZ9FQe2RnNdVsGPxgigHwJOGVMsxHz+7Cj348Z
TT64qxrK0TpKpSYBEApPptFLBjOCYUNhmhyaTJVi1hYpHcCcFDvG054vZHswIz2a
DoTwkLgaHQiQ8OdkRtTV0dMhhaIGWRMAIz+o3c0bkY5pJT+IhyushNC+AaQ86eTP
cfuvyIqTcJSJTprjio1uiK7DAuXu/6GY7NMf69po5cbqceLREznKSSqLO3G5zpvy
gcXW0k4AgC2nymfki1UC2sToHASRkIJuuM1mqZM6CKGqdm1xwqF+xBaoTghHieCf
WR4aiB7aRAHfrmW/8t4AFBQc7Efb3ceB3s/batz307wawiMaLX9VaTky8BPBAt0x
v3RCBAxg8dYGOMyYiCHvTYz4FzV4znJRokBVODpP1ro2AXtcMPOx1t+EweL7X1Yl
V0Q0HVG914f/2fnMkxwWIkWuyTE89D0XzvxxTeyw7nerA3buuHpdlE73S1M5f41T
Tac/5xtX41V+zK2xdfxzztVPxbIZsoErsiEhznZGTcE7aw4bIEXWj9kqPgN9B6HM
9ksK2l3wQVUBpjpQo5d8sNomPzwzE2QHB6J4JA8u408uy6tO5VeZpMy6UoU7UstO
arnJGSTI7yeZsJYfEaGLLpa4XqNJVxe9XLW6zuOCWWIdFFh9FLQTmO63fbVZYniR
rGvuzkxgyydDVhbxPnI8cXJEm9rp3KgRomNoiDpxoeGoWqyyAR2jnUe/gG4O9Hdv
XxP6M6KyU47OyCAT0T+d01krqNOdbKufcQ33xqo2px3Vsy4A/qZl0jwa165e6SR+
xBAuqzXsHk0dyorTR/zebMVT9sqV0Mhk3Z9+wZJukmP1f9NZE5WXUqJXlT2GBuOV
hpjP3wZ0+xtXZ6ngKb65UdOdPLAbvHZoDWosgFdME8qEUcIlR8W7Idp2mY/XT5cu
MQ5JgaPsSKxidU5J7+WzjfZl8nWpM3vWIo9NjiSTB3hUwEXagGQZoP7cJ6yofmp8
wKxXQv9zxvi5R9++8fnHHhMGqkSEUSYL6yX1pLBxY/VGFC7NGwO7WZuht2ZENRv5
t1akcHJu4OpWXfwtarkTG2NaD0ZBRHGiXGgBIkXUwQr6sr7bA33bIEfdcuPw3/Gd
7JPyi3xuRx4LS5ZKVEJkWv6z1b08rzqu4KITAWEsZvKciPLCpBo/kzO7jHoT8ANU
4QrnnPd2EmObbTJSmHk0S43rlml+EDOAbXMY9sDrZc2723vgtOvnhWhIJn11sb7j
0tk/il+ZG75EGdvbA9Ifm09zuPRpjn6tJko9+/s4ezVH3Ca9Wp8w1Hxm77GNpry1
6Av26W2j5YF9x3puKmGxJY5CAb+xukGFJVYfE36XE4GWBQtIvi4AheB8aRupm/8i
GqiyRo1UiMwM2uhROFFbTNWhpkYUGzbDRsIzLMpr3QWXTmc+OZx/fNwGwsntDYmD
GEawzxxtjSZWHWOW4/aQZjD5+E1IbdLIfY0xRXBn+Xka/07+NQ/mUX/mlNJQaBWn
5pW36T8hTWZpKjY4lMyyFwSvKxQexaar54YkEuIgQ+dPP1ShPMVf/ESZickZlMOs
7wA6R+LyrzUVnq4VHLaWbPu7AIV3q8zV4u3nV3lEoPU/ZJyu0FmgZNHTWi9+7Ua3
cgRBsIidd9ilL5BJ7N1BTWJyD8mBAWwYw2E+VOxLmXIhkg0W2u9DUx0IskQdjeGl
P5bgn2HB1Rk9T+9mSEPMK1w6kG4M5ybxIbi2QoRtL26EPFx/32vx68ZqHcgBtvmk
`protect END_PROTECTED
