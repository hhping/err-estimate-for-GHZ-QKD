`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lhgwDVGaCuEfWQBDbkLhrUqHr+njaPVgUavASSptckC5GpI+ftbC1J286pSyjuic
dtgr4ZTRVYQPcJSKZMNr3XItjWjBgeslRjYQfgZPmOGN2ivvT9jMrj5dBYiv3hqD
g9WJG6LN37P4FBG8DxmmYqFLqz5cC6rtcuJHVdMRaMzK4KB/RgwhEQnXNOA2Wk2U
fng/Zq4FbVaWXWgwSFtY/KoNmi5tKx2nsGc4UuuUruYp+OX+tAbTOfO1X05SzQ+r
2H+BHwdz04XA7mBFh50rMrhhp9taSSc5Kul46fBfnyCz1d1+Yuq003rn7oxvgGvP
yyCi4JURb4apBIIeFeHhZoRn/SnYlWuoI2By5LxO1A0b8Nn945btZ148ahvlLX5Q
cCxBw0JhTK7DFleJS3KKCWcMbURRz/JtTtFPYLU0dnUdFbGi2H/BfgUa3/B8Y8/R
TsuLXgXMdEdJl+sgDHoiTudeidJDmMGsoSl/jKBnpkmmTFNl1NZpzTsYVlio01PE
BHuBPtU8RXFBM4cdfelUQwDYMQtfbpWKCWbPVS557cW9527jixjyj5hwnv8ecOQs
aDuHqyeMGBrXeKkmr7x77EpKUCcgzA1cqKVuYXuyyKjNIAfm+PvVJ0su+ZhClR5y
JtBjZ0cZHpsbn/rQFXL4m4MEZDae5tQBn33lTW+k9srQ1/J2eRiQahw5H0uv7yAI
vj3l+qctZ+QU63fV8kTbkYopJTeglP7tEbUQfbsFOFUnYoyRW90tpI5XR5wbjfb8
gb6AeaczcjweuGXULfePOlq/MNPqAznBkS9hCHKQtqANhGErH6EGd4EZIc7P0+24
YLsKUym7fT5+mbrXQtMdYB753Dc3r7ELG7wqS2s44/hUOLmdXIiHD0dKmkVn4ZJj
tz4PAu1/uCHRTB+Ybdngs4JEgA4450Fp3CTtomdqFZBIPwzmDh6Z5J3GFIDihN2c
oQ1jYffw4hcaepxjryKyMEeK+NW6WQqmR3DS5Uy1dHKFNeuQFLBcXJb1AKaUfYdx
WqnIi/9UHxG6VM8l9x+aRGrgbaHLdUdY7ow27xJWvqdFzbcDMh4Pxn/lurFbd2Mn
RLEeeyYfWa/tUKCJ1aMoOg/DHkMnF+we0084Ixa6csvkfd89oKUSflID0oy7DHeB
lvKlexLNt4mbO0izuCd9NqC6aI7j146pKNAFHepE6rwB3LllLyLMgf2CP35DL1zE
NrisfF7JoeoDmIFnIxGYMtvH0KrPmNwO+mMOjp+VKQoNcpgf8t6g9C6ufWouo4St
whS8DTgjHEds1CYQ8HRx+ttiX80nC10xRSktdhwECwpj5F3Bhf6ZVludxVT8/yyU
P7PNeD7AfxUnIIa/ihswjGZYo8XdEIuzTMV8UUV3uYEhNPDdH6ok6xItbDLbKYu7
`protect END_PROTECTED
