`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TPmhfGJ7inJZ7RQwayQeCbbtv+5o8BbCjz2hfpnS9KVFLRm1GL96oUClwLcWJEkm
2RNW7IRgwif2lJJHGkXRJH6nZ/OU6ZQa/+Py4N6HqL6SLZ5SSDMIe5gGk3IzegFu
pi/Qm7bvNtzu1x+sSLA+23cl8jsOuC2LBtaMsnalj7pkcNVnrPp5+AHHIi73e6PC
O8oRfzzUiX70KIS8hHmHbFK8eAEnPXDCxffkWm2yPDdJvkYypQsVG7tVy8cVbdHj
Z4j5vGYyKwW2aviWCaf+5LtcFPHugm5YYY4FZnYXt/95CeK2p2TGzXPV6Q+Px8fL
fvNgxpDPg6duNqp6uYMQTjuNKITEqfhNkiJWuL3KBKnt+QohaoN3Ol8B1ZuYmZQA
H6k8N5gggZXN4POrTdEhdiZsKdbhUK8yVwyf0li9aCYm7nBpqs68T+FN4SY4gTvn
yWuyLxSepFkapUEILg/kBafGIO0CpC3eHhBA240R5e0=
`protect END_PROTECTED
