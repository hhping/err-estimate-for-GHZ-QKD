`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FRBYbTWY9PFS5ER209MjcxyqHQhzbxwP1cF6dCFb7UZ5e27L4beGhA868PyXJuxl
q2HRy2yE6NScT8eTmgOsHHM0AA5Eb/Mw/omnq2aH9tWebyHCOKrlferaIDMcAqxc
nOZyuhzXUKg+LZwo0H1Mh9UK/xiMiWTrve97zAGGmBPRebjnAuoBd/+BGMarcxYo
aWXCGsQW2ABYjeTZBRHixUqT0iZU3gkBCPTIw4Y4m2tReeOYjGsuOYXjpD9Bkkkk
UupQoDhXlCJZmm9cemDIO9b31m5aBjIrBvePOtjuz3InxmH2NicEbFznRPwIEFHv
BX1ZWfIqcde0BR6RSOdZc2zyUJcNOzipvk/pbkgdZhPTrwjloO1CXEVchE4nUJbk
YJDD0DAdgs2SFCn3aBg0C7sO7AX0k9pWevNWhGiXqLi1kyj5WuBAF3AvHKdMnSx9
I1cc7E4Vce5c5fqnx5KzkabWPTGE/BxVx03xnndsTvSEJtlPajMeyjUndckOJDdg
eFdw/WzfOj6op2kLAlnJc5pkNlEodkQhuq6i3D5Yl+TIsdcR7nFku6Ly6ADnet79
BpveEqx97fnvAoPCM4iabIMpPFK6EQV86XjxOM+3epSLU97T9Nqec1n3cPrI6AQI
qJYVCJZDtEqBIFAYOQbFip4lvlKKrIVGyF5ZL8yvrwoYvHNzkiqghbvEhBfjL7H1
ttT3EdJ5o18GJ2QctJXsYGedpdZun7Zh9zsTliWxTJVCnRF/iXxQgKDQ/yZp9gTW
AqvD5QPqkSJ2i0rMMGwKKYG7j1pLEWQgC1YuZm0x2+hgcmq7VBCleeng30MOM78n
XAkLsdODdY9CrCDOW9qWINAuopj7j37H+Q26DarDQqMJ9ycpMQFpUCZfGv40gpvJ
S4WzmtwRRT3PCnrfzyJay3hTdDqAUDWblEreMb/ZMc0Uy8Ebq0C4rEFloqJJXuNq
AqYKbTLflpuUG9bjAqN6TA8zilfjF/Zli/S6IX56epborBdUBpNze9KHrZsQgMu/
Latb49GvqU/JVNISVriY0pl39tKBnAqyKgBczfl8EDvYkeCdanV2zhsNYNPLVPvf
y9ir/Xrt2IltGtojhPnWAimSKZWUpO7iRdo5XHVfqlOapBni2VmLYW93ZwMjwvzo
P4nmBK9uBvFyjzIDqgDhL0EMu442pjHPU4JM4s8gyRszg35guHurpUWO4BtByLZ9
U87042zGQHfvUaBlPQHmIPbrDC4CCqBZPdrRcXGVA43fE3Voi2uEXxoEYtB/hC1d
I8MiJXrlqXnVihHffVuAWuYLgAKI88Kfxsefue2Uv3zcaT9OF6lCze3fXM+8RaZ+
PYyXweO+EMJfWxL+1euC1tT7EocbiIG72+29vcuwSqkcuJ54wmovm2zLzhh2jbEq
9OF/T86leaDoUllv7SmtplZOrxar+rLChbPwuvzfPrnQbXEpUVGNIn5gJhrpvpUL
4Wp6FptK2Nj8LoIliCTTfO+drfbtE4L3W0xbzU11nUrQzPrlz0pa574I4OeWMKrA
ff/d2SzVvGi7BAcQramA/89aUbGkWz2hj6Cr0ytFhLzJg4dAyPlwPntFNs51lVdy
RJ8URupdIRowLiCfd/tEVnXDetRxs0i8h/I3hl7U5W9ZfzhW9qDI/A5+25A2h28D
A/3PXeLIk+DI116d7ksxvgILJpoigJl0yFvJxHbr6K5wB0G4ikHevs0ZEAoGXDrM
3d9ssDHO76xXjszJzRALem4y05Em/p3gQeM2cyvxTcuh1J6iTCk0XyLh8a2dAKP7
lix4invCdbdlWEyqheKcvuPp7ks23tdXN3cZCTeHJDVphIaqIhobDZAC+o3ocmj2
NB/+XpAns+wMRcYrAOcqjqU3orrbJrv+yD/mR95j5wggN3TE1ULoEBnE8coEcNdV
NM6/on5X+g1Ah8T2bkD3TyuEwHLcgzgKcjVEs8+/zY5PjEZOFbVItNIqcnjaDNPQ
e5hvYoAGL7cvDK9LyDggj5nPbHhpPbe9A+dEy57vYGs+Tkazse0Rwc0xd2TYuzgt
E0t73QP2K3LgQ3hOVGgYUH9IFiqPgty+N746qV0o+bIJOYsfefqB8cD+KuTobMva
o3vfvzABwpbGSrMU10NDA48dt5FCtf01YCKa58bZkCKnwFP4OY/58Zr2FCJg5Bdz
iZ8T15m149yWzcq9HoF6o9DT93LQcmNmdv4pkzbTCV7rjuBMF+5BvvFYTLLVwcWG
OCUJ+rV4e84pXGvuRRyM0Eef/8uKuSPzUrrVEnO15py+Eo/p108SGNu80L+bamov
KG0tdA8/c5TEjyq38D64FZp7Kr5l4ff5bWTJ7+vHrotuCJY1PWtjR85NJ7+lWz8j
Gy1MNRdB8zEGPAsjBKGNHgkHsOPwTGHbC0ksoY5GxOW7qL9vjpAS81zGr3tcLuim
lEoC/w7sW0/varjEjYXmxvV3TQnvrqvdp/mDXPwmHA5mWcZ1b68m4/Re8PBZQh7x
p+Gaf+vd9CuLE1a1uQybQe3b5pwsTKayZgCvpIFxtg8glYFcmRZG+UGOox4DaAq1
Uap5FTUVbSCLKC01cfMXK1mNpOp615X+WUWBnEknxOr1TihnRBY3sHsIH2hwZ/iO
9rRwNQDZeMpUMQQYWGq7NcDi6yr2jGziJZXFjoxGVPn9DQp1t/imiTB8jIFe8x9Y
F96BsMZToU1SnUSdBkO8+A==
`protect END_PROTECTED
