`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SY0euTZpyX0gNIYjSiC9oCXrzOb8HIVE8GCLmZX4J4VmANOAeDACRx3CzKdqaaVA
NTLAkNB38ZV6BUjNvjOxxghqGl8vidhomNLUx1I4dktuNoOw3WVh59AS15DCJBKV
zLxfJPZ1LIr+0xZsZHIlv9HwtKpZjHAbz0YfsAHvo+jk4h6VOCcmzvMG+lQ0wFUV
mIxr9hdskUqpYU/KozWNXrh1D5hH83tURY5A8CdMY+pobnkvARIxk7gi/qY044J9
L4D/Gnv1BxowQcHQkpStjrUD6SXKTTePTtLa/anQUtCwLdb3Ro75KP49ZADIMYz4
d8Hfy9GC+jOwhBE8bUwe/q5kQNNdHhT4l4CFy5btFbCdsyK7aH5kwUwvsX/r/h2x
WhJvnQ4hSM3Op/LGiioRhbGaK4tNuDU1HeDiz6ren21NeMfgqvMJ1ZrcXHehRcWM
6DGAaPKxIO6WVWOBKfLM8xKalNU5n8Y7gaj/F6rEJduEVSYz5U50KS8lOt+k35BH
UvqmmZe0lvtAXHz+dMHE7PMSk0RN6S7vd9lEq6F6LmVNdF7Yikr86UWPGQTUMGPD
R6v4gggC3B5M8FqbZnAfTwsom4DJimnYQ7s4g6HsTmP0BdtAo69xdAWMV0LJkAw6
ite2Oy5clrbMpHrRWRyFqzBLX2vj/TN3oDYyq0kq1tWPQGXbvyHkpLhe/8WZUSAQ
/n2XsS5HkQV0kiH050evuZ01+sfFXcxpCxcrNTaKzbqMNVctTuhtVLWxOwFP2bSm
YubLZeS1Y2iHcRpBg1NcU28zX+NBfe0ubwi82Qvt45xtGwD9DO2ecPQrDJfmV49M
F8Vg/YM7aMJBT2B1P7yrMRfTmY8cBfLwcvEftkPHNhT1LwiDfgSVr+13bvqJ/r7T
0eH5vUloGp8Rt1KXOBkT7l/GcMy/PPCeDcB4rVc3yGs7ay172HDSZm2GrqSkc30V
ioFIYRcjkEiKCfDPDML0Ez1/ql3Za9pS9DVAJpsKt+4fT1Qi/iy5FXQlCPSBak9C
d56ZTQOMYDBsI6VTO7NpRMRFGzXprGNxAIBQSpQeOmF4LtZsQ6trJ2Oe5zRS94kr
seDR4Hm6VByJ0sOtoX+xCxgbCMrwFGLx7Ji2aGBp5PA1t8/Q6Jdbm1V+V4u5rJzw
dUZUt+TD2ji4KT6YWqra7SmZ9fagaSsgfORBwEws1e6Hn0Kd4gNagCJlLoHnbPAF
Z+5gobRGyEDSgGhjcvRLPMASnRp2bMM5oSU4f44/cFofA2TfQZ+7HnBOQSaj5MjY
cq/OQ0uBgY2ynpSLdINyiKkQNXIG8qISoS8ZwBoOQHWoocnC+W213MNFoXy7FHVr
SUp/VyWJm1tqLJdjmh0+oKxuO1su3m6ZeLCk3WTD1l9sZEkZa0hqQgSATXQvVspL
okGoUscJXokJBVSv2Wks0RzZ1qvqNlVcJFw7mwrTgESWFmIXnG5JEdwKLJ/j4NGH
GUJ1hhROJu0oNpFQXe6iNCLPRR5XcwIZvy1umlGMZgXdKGJ3QOy87iyxhrt8CGPr
YYYSpx8QQaKOMRaVAuyQlpqR9ehvoN88XBoDxo7VyNZV8paxAAJe+PJrAB3jeqXL
/0211ogNqQ+rBu+igu//lF79p3zLOyh6nFGNGNeBZNgLi778LYbsNLnnix58SBsY
7U+40RNUw/1xeSRVuepcffL24fzlqNP5XKZUhtQyf+bCNsxKZW8aVARCwb78TK0y
V6TMf5CayMjWUNUFVziJnU1U9MWvdC7HcGq8hKxEYMqf5c+ZMeqVVh4/zmMu/nFM
4QFD0D0kcCgTk+I2Sze1ukEcXJyj3LvEUhOHVgygqV/VBZ1oF+WQsQnib+s7Dn4g
yN4+okW+WsGXeMNDssJ/xeOnUzxo5spzc2WOV2mEbnMGDw8aZ4cgVrVJ5ZJUWTEt
6RYKrZ0/mwABNQjihULBdcu4pXscMsAAk/DTAkG+yZ5mw/i+Mw/e8KMp8L1JIeSv
sBngJRMj80fYru5/lihL4FTCRFyPSYWvfn42hvojrb6nMqxYfLx2RSsT5dQYLF1Y
RqwVcmfsK1yOKW9FV+Zah9L3oOLO8Y87RMMWDxBMoKXuREj7tAKfzQngN5FY0Org
L9TS15bHmHHUCAVjIUAd5zQ3qZcr7kDCtn/xLZTU/Yk=
`protect END_PROTECTED
