`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iflAc3O36aPt1Vqz2KBnS9C7zMNO7fDiXznIw+nslH4tRK9p1abZ5X797f45cWcs
KL/hiyBgVeg4ThWRmNrsskThQbVoxHEe2Y2S9suAX1cRCr8RmUTpom4f2RcCzr3p
BDpf1drDJrqxTf5IH2mRZhxmwlAp6MNtzRnjLKCq9YfsB2ysT0yu3j9s3woCDcbR
CzBJ3HV6HXdqR0N4wpieElfSoJUUc/Vbz1oxeBOVgf+UCVWW8mWGo+XTlOdSmVEF
mPh77w10M9AUEW+LQ2RxGmFUIuRLHuEp2VW3QQ6LBSrfZ1yM3vfmpruDzt1xb74I
J7RlDcMUHLnsWlMCf5uoE1QXGKYVHkHRYv6cXs3lTsThIv1CyAxntfvddwWeY6R+
5v6J8KjkFh47IFVhWzyD6+AlSITEoXf+gBLssP9GGIHvEP3h9RbU7whZWfu1oSRN
SF44YhyWkKDwGJ11ATEarhepMhiqCYxazyEScDrEA8nwwTSExiRgN/awnK2Z55xg
6dOGvDNjtppWaYjjzSjJLPt+1gg3rAdWRiDO5T58WdWsqGB459OzBtjKMbDp9A6e
0DFMdoj2ne/7r0FWsRRASEOOTRIJrKBYvpW6sZ3uUix8th15k1DfMLdOJ998iDwu
hihxVRvW6X92Jlw8LoQle6gJDB2+MklW8GHK8Ac+tlBX0G8lWBW9GRYxg43ye+30
OboEksihuEbpaw52pi8JsxnkfOAhb6ALu/jywWnxrM47AQdq0gzC+0nFzlS/AxMX
kN5Lh9fB8tN30il6afFZ3pImSbMfOoaJUCSYmE0evKly4KcTYOlY1Q0RcTaEcqAK
MRfD1nN5lowqFvYcEK2lzV+v4sSqzOKQRq1EKri7FVpLxE2ufDLuk1Em08XoZ21F
P3p1lxNaSNofG9kkAi86P0xgF0/qpu8cxFI4/MxNJZZpiiXRzMVW5XIE0sSxw0Ph
Gq+1ifJje7DRkehjgZW8I4bJomFAFR3iSlEcEbG6lXRaEWzg3bd1698WMtZSeSuD
iSdgBSBpis4zMG2cCi3e+Lo0ajHuTtm/WtuUOLCLa/iiDgytLF2YaoKifYVt6GBG
Bz6J6Di3X6QxCk2aw6Oi/+H15vDXn6TdNxXUER6yCyNli8bU79t4Fg/ZYwZl6uE+
5U3QpEeoQA0aBGZSEqbf/wspHbEw7VoOlef72ueNPVLfjQOK4uDUCnxUpcp+HMvx
xtVSnY+9DoVzqwEYNoB12CzgvJ7j3WFLxbHm2OTzpWBiLIbwoSVUibSk8WJNaY3z
/LYIIyTHte6hVGPNnI67zRJivP+mO+cyWodduIkEXvw=
`protect END_PROTECTED
