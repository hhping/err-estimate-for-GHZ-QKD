`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cyip6A7wgdaZtz8ue5gWath+hkq0yrdL84Ja2WxAtfhgGs71+7s7GYYPhc/0A05Q
VPg8DS4r5FJF/WD9P50dsADSqaw6x4YVz11w9WLerNoT0o3LmoPMU1PVtdDnP4kK
LyfhLGWvEVrQ0CTnmo9S92SpU4MMlYPO21BvQMjKiHxrW2hRg/myUybDGd0Zqr3Y
4gRyUnDeKicDFf9nBrQFsIMvERiBSvM1qVCmSJc36CWU4KUwKtZQS89tSU8aluAf
rjdH1rZKCTv/9e9l7JGrP836nljyH9o/m+J16MvCnsWpB/aEsLPfp5teXFKLaTJZ
q1LdZlo2s2qakV90wa87i0xtdlCY8Z6FiVwmcbWajW92oG7sRLxbTkWG5yztOpt1
gN4+XOsibOnhRm2ahSgtPOPimbwcq6XUyabJ4D4ZfuYTf7yXfn3BX2dEk5yLrxG+
j5/iYAPUNyZpZl/U0hkzm/43OHTJ3T9RcZUIlPdkWkb2AgeSbbTLGBlVLdG8iyFR
`protect END_PROTECTED
