`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mmrOIFj2NH12SqyhAJTZdCJOTAgnSbYYhtpSV/DZWLmliapyDeDcfFP4W1i22VmM
3XUN/ciRHqai74sEN4ZSAWuZMLN/yVJ+LgIZQk3htA0mEDZk+omZa2ud3WD1Mrau
xhIHB0HmowbooadJChKW4CpgGZ8tp3BYFWJdJCnDurswFWBAzypiiNbv6uBcwWX6
592ogQV+h7iBfkjZGiun77KztOLdoDH2Itl/hyLd9iumdNrqK7fjb9o7/O0v1Ytt
j3P9Vlt7NxehXSqGqeaMmyJ9DQnoCuT6jXxcX5UsuYIrtV/2jEw4RmcItsIBEvIK
BmPVTegnk7cqj7BH1pmt0FjytX/pVlLbB1cmkbnW5peRUfBl4sEKBQSO8fZKuaK5
wvLHFF+rh2PnBIqEtkx001bSdSpAem6Pifu4W29FukuxNWtYWLJOiH6e1iKIjdt5
PYuus13FOmSnPneqG446/g7yLiL5ZEU8K0E9Jhm/xeXmsvVtg3VA9xdgEMQznHlH
CXfOWQh2UDKRuMkhMg3oVqfVCsztkVP3WMGVCaW31iJSWsjchUQD6fbI/cj7UJ2u
zikZesUhvvsg/RCLf1CUpRgKv07mf5h9yOnnDbw1Y43gaX4FyTd9sqdRxMZXBaZV
7fJeCg0SVFgZYhk3z96SeQx6L+Tmydz/v2e2nAYMkMfMt1V3y4k3wEfQgcy3d1uy
WOthgTLruX7RKsb3opmh12bP5pSwnWaDAhtWAMA9oIOcpchDkbvOrbNkMnbSsddI
FMFxcndJAQ5yE/FImyDc9UzT9bDZHBR35ridUWC8jB8C6B0HcYmxMUqw1riiJJyx
M1IiHg6lGcwwuJBaik16PHfrp5Yex6odTpsuylKcWFEjdJJHjSe/QkFTT3Tq3rrv
pfkBUH66b8MlSV9KCwoPXmm7zq58OvguFlaEFgb6HCiecWtXWfeh3nZOScpphKe7
cE5sjIh798sAqqJAiiYgeqM8nJSa8cyjJCl5X4RJqaver3qrQ3llv6BMwe9hGMX/
jkLM3fRnwOStjze+WHhvlKq71dIAxyEtDQ+WXX4Cy+t6ljvYbgekHyd5TUjEGS7t
tIq+m62ldui9MFKtt6KMzmAkYQj9QVat3gaR2H73j+Jb7rJWmk4R+KqOzNijyeC6
oEB1bLYHLnaKKxJrpClw0uAuCWgTwV5StKIOm4frEkD4nV5/ulWK0QhS+EG42c5x
YSzhQAO+FMszmhWm14yl0l3Yx3H7R+u0dWlV3SQPKXnaxZOm8gZfHhMjCSoh8GgJ
Y9fjgs4nuciKUydpEpx0mUbl8j6sGQuGUxSUa+yRq4dOWhyj0Mh9r+JscgucFl2t
OKA/ZwmT9wrzv7nQBqB26hdMzAqqC7zjL7E24lH7ZeIqdNcfNvdcajeiPXYfL1ly
X9E15zvokssPXt2raSirajO4jYtn/ntOYzGwKWMmO6QlmI32YnB1Opyx4tuR3hvn
KpOtx5+t3vH+JzSfvrdaERBptpDKPOUrWuDNumtFX2tY4k/0fqYoo3o8lxEVG7Mo
s3NisAYrA20W/CXOZ4th+8mE2Ng7u2nszT1b79uOy8/YRaLZPkStF7AFWtWZ4Bzb
1eOyx1W/2ayNwn50SehatIReaMo2DATDbFby54rcWdNF/PxKREB3TJJpNrWNbhZk
R9pMPVGssIF289s6X0+78YrWlWKpr4bRdvDoKnEmyFrNE2aGY+cvSoHWe/fYhDpp
LmFVIr3wuO5KUTplFilau9DAPjKZV5uHVlBi7nD2Z9EzQUkHi7zTI0f8aYeTCC0c
5QWfxYOshmRUmEqocSDHtcn+bc8YA18W7MKXY7ig+7z+vdR+qLReFrzuT3TFGEdo
WnJG0GPyAuvdUi9CJay+6AZQL7MWQF2FOeogk8f/yMpamwBBLckojhpR8sDkWujR
QFPJp39SaD0goHmULWUTeDyZANSLe8fV+SfQWBY6P1YWlMxFB6v5y8WcgAuu0yqI
xWhvWmbhsOa+5f85OlXCCEq5OYGQb+dvwQjvW3LmmfzjbrnNihElgcUxbHu5E64q
3VgLakVraFoTAB5LNc329miQPPcEElXlIkBhMH/aTV23roUPXCvldXs498GDwzGG
Vh6/T2CPUInFbQwfgLmvTzU1nR+GlcGt/g9nAR07IaWvuELJlFsslFnHs5HhPFK0
n+5MHGhkBBXfSfsMMxNOWHB2rCAa6rVBKYqhbKYCvFPUc2LlC4L6IM5pfE/zGv1y
yy3UtX4//A84Wdomj8VrONTMSedgwji2csKhlVeKW6/zSi2dDQuS0IKJxnHJyQOR
wblcd1c5u71KQ/IkaWecCauQSu99/Tq/eHNazheMBUINPXm2pjy2peo4LqIlYpfE
OgYEd2RyDU9r4NKAnsy6jeiER+z0jraastxNWZzTWhTDudt3LAU3VhFvic3MBfNo
ydUP40h9v+ZpsyeDjg0nUpuggYcmDq5A4dJ5gqMtZt2MR3oe4ZCTy6EjKTJn1iU0
wkVhLJmHUjTnr77x23jYWbHjqxm/d9dG+5QxKLhJLcU9OLt+WdHpfK6pvV7SjPWz
fJCl4HEKRhqjwRkMloj6fia6ypc2yHO1sPa8LWXWVzegju1J9IPvlZTvMrhH4CVn
E+fsCxpj3XzM1sJbyhp7vW4gCD2/UleEms0LKkSj3jq3CedrXJnSGOUAXIFux6fF
c5nqJzigwt2JiLVaR+/iGIhQgTqE4Eh2dRB3s65Tqugfvrnc+2zl08A2HMBotNfd
3pvv+rFgb6nDCu70Lo3/weoirt2OpEix79iG6OPVOaNRszhbBx06pW/OWdCfpGfq
RguFGzq80iTkZ3fW1QGwbHVaNhzM21+7AVn5ORk8K8NNhTmwYxcr9dzQdSYq6Z7p
QrhM4wwXvnyQImPE4yOBm4Lj4RRpsWllVYckKR1UZPaFIZmNSlQ2mpOYufabZ5T2
21tE30l2G0yVc1YGbj/07XqOpUmJUMT7JhhGfTEyVi3+NU2eRNsdVELl3T3PWvTK
ohksKmeh3lBTvwYbJbRgfWGTxiAidE1cdLiG3CR7n4k3wOONbkBCKZJAr395p2Pw
XneDs+Vz5OGDk76UxJZn3kHopfroA/3xKf517R1UVvbtBoliSmHwUKOtQlK2yWE/
a3SNHkvSbA6f5CupicrjWN50oVPcmMV9zu5XCVuQ4tZ1T/HUe1FtddhPf00I6XBA
Cgxi1ght6fqUJwz56piGtjNaDemMeUrh/CA9h0UM1YypH8T4PnWv2E1dd1Ug/RvG
tV15I1Gkf9e3oOiYi+/y0y7dFFsZ9SR0z/CO1BOzet1A69VSyz6+qt9iXXttcYTK
hJQ8f5JJcYu2i9FMe9QBmWaKTPjTMT0G/Sq7ZodHnJpRHe+lz5Y8xpYmlg73xObF
tR0V541wi+AcODv+hMbqlAZc4YdKP+/ZTu9owToyfTNfdjaN+nkoKQkLtCKSGkLy
J0G7DJNkIQswrPq4ONOF+78NtelsZlpekBzdVb4moFxAxmEMEwe9DODT2zcLy5Ym
T08r4psZGBc+rY6pquJ8gEQOLmtrQLV/wtMCq7sZByM1bg2ZElECUb16baXySz/S
XTh5tuM7tl2TfLc3a2xCGFjX9avmY+OA+oXw2cuRJJX1QWGWJhVebBf7L4fpK2ZD
zpYft8l/0MepYFUUk2+TcNIB6jk1oc/eY3J3xSJOp/cx5g7IbTK3v3AmrwY8XLn1
lVtWFrKHmRp5WpotBreuLu8xBxwfqASSly9R32OwLcr70vjo5sOQjux/cvjdZ4R5
q+R91RiuZFuq7EDgYHNZ3+YSb3VRKmXIFXunHbqDedLmygZ9UOlHJ1ovDP3NrmoW
ad4xDIIwodNM+v5rSBmgdSokUIf6hZIY5DaNjbbvbZZKq4ynRCleA33O4fBNdH5o
cJrFRzD6F1lhp6PU11/dgc99O7BYfIwQY/xHgOca6yqtrBuEUDWiHVJTDJ+kOBdG
Vg4wvTn/t9rkaXGb7OK37zk11EkXAeTAoO2hYopWDV8+E9ESm15/Luj6HpVXsNBR
ptw9t9RNG95bL5eWwp5N/OtfapUjEP2hxuIOsB0lUY4dLmaZC49zkgHwQO3VUL+b
HdaMIH0bOTKF579W+w8kn+kmoEnpLxQrWaIrTgccdkMZhGWYVwhVtpcHtal22y7o
n4eI84zx994CuJYrcQYtZFJx8mykCGW9mS0mm5itl2nqNBfaePFXak+BAnIgZST/
sPhNamRKNG32CqfxXuFBHFRTTOlI6J5ah/m3wZ4hNMqVvgSJDkYjNAmCveRjk18G
WqLtM0Jtd5rSCfFw/e2ggcQlyVugdudfrXNrBac+dWNfgJfZalxgeIHync4PSxnz
Aq7xGax4+BN9/091zUug5eaPB+yMJ/Z+CxjHV+WDMMTq9fkbtaDHj5s/5z03qWBi
IhydGedaSybxjAuz36ITua6IewxOT6sjj/HrwT81aCNgZsKecLybnPc/XC4K/pSj
KF9Xj4VpZiaXLL8Cu0gOvqD3XkKgwMEeUkztQYZo+qmsS5OZpu1nJ+ZYimjB6OkW
wmthq4aHpyAW3+aA/v1Svt2hDZ/nRO+KJCpdF96w35u4PMl3j+L72cz3wJDAkKi8
oq8a6v3FDSENvnKAOXtahXdbdrVLs76GPg8p7rtE4bO5LAmMvfwEJmn+IyEr41w8
ZxmtUW4Ooct1Q6dmkzxf6O9u1QxOTsjBqBIWkdKkk2O4jI1Vj5vQIUUe9PdZ28iX
NebCdDhN1U95o7TgW7nVpa0y/TbaySJa+gXDcVGUlNN47rhpi/BZVv/izdW6Z+fT
7IkdcP7uCMjfU1aAN2d0FLMt02XaE2C7NIa+YwLnBiVnUI/rvJ7KyukZRgEoD5Ks
zPMfzUh7pSvq2VejupuBqQ==
`protect END_PROTECTED
