`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
twj1QRh0gRMvmMph7jWC8dOtgA8ZBjQr7WihCz0V13wrKg0jJQLMRrysShc06/fc
q87U1vZYbxBCZDS3OUFjPm4PkcA29b0cAyFQLOjFDaSyJw5WDj53OKq86CThC1Dk
XGzryNUGPES6lu9X6Gjx67nLm2oiSuelbQz7Z+M3jUu7I+j5e7ahlY/8a+PIKbjy
psWz6rL4Q/e37LV5vXQVmQdFeq/mfEAB4ske5aT6fM628mPaKqgjsCY5rSBRhllt
UuvtYe+SMAYd7IZrNWe97nfNc8XHA83h11n3m/F0yxlAc2AkHNLeXi492oVJ/Ahw
mFaO+vFML2zfAa2q5WC0AwpwFaBYilH46m9Ew1utwMoTuRnSiEzPcywP1A//jFxp
+x7QWfGEQk4nYyWzWmt/xld7wIrSPUIpbJkaZEN0RI0NVrHWWITzd8zm5EQ7Q7pt
`protect END_PROTECTED
