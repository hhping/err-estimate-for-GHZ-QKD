`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hkSmHk7FsEfgJPGrCkVq7qvZuR2D7d5A/FJ8805F09pzB/O2h9f/zOkXi9l29Wzz
z1mr6k9jb14fTzjl+8Njn3fQROxcJ1eVhgP1gvnU39IeqqGNkQPKzDoubwDxGdtF
bTp1i/cbjJiva2uPpLjJrB3p1zoDp0Kepy8bbEZbo7o4ZnHKiLg1NwBsD2xm0lM0
kxI4H5qfDj832szu+DyXkiNkPTpiMIkdvCEnJ2uwSgjgw8/qBGRwG2R5zh/YggQt
jV68ofhMNC3Nl9j5PJNoUCvJtm9ASPBIOI2RvgkdIHCD6EGdODOvQR/G6nqsCqnp
NrMem8Xbw9L6ruSTm165NSj8J/hNK20qfmrYjzhuU22RSjYw/GJAGbGyyJXz8qXC
9bSWJ96ufJ/0NsaOPUXdld2+MphdRBUxHkqj4EimHK+j4M/gmZ4ZzPnZs+95yFr/
FbcH0GS/yu91ILB5jt2s0ZSu8NCtOWp+Hw1qFjNLLt+hA9Fk2rsrv3YZ8l3Vk4N8
/Rc+PPzrCNFpIFEwRkjEi4ysENOEfS1LpKEl8JwNQnD425gzgo2VyQqhDuP9sjAW
oo+M48BYvdmrHZIUkVDfRE35YvZHZEsEOId25ceTvIU7ez8PQRvK81Z/FntgyHSk
pXscga4XRgDH1oM0bST7+4Q2eNtcDpbUQS6QO2w6h0oJuCh5UGVdzKZRYXl6hxO/
dIZnB5bsFWDdcaQ2syXKC4olobUk1qIUtBDYzHzuaXR9Q0LgXftmtycNx1+/ryy+
DGVUj35SuPy5tUY4ZVMO9N0IxoPW8lpV4dtq3+mtMT1SNNADUPRlsHI8SJAaivN2
cIJ8x/oGi/QMc2s6fb/jvZYM2rM//FF0pCr5u6UzQ+OjjFD1QXINna3fL0E0I7hZ
qM1d5zwXVjcBzujQfSrzP6mQqqJgqKHjOmPM69qJBhuvs9itmtnhmNe9AKVPfnJo
wOP7RqifYsT2J7n3FnHegGWdBfNUkpI4Yys83ekZvTYm49VNUfYxhw4Az3GUtVcY
dT92hCM6Nanmg6BOu8mKdVDZ3MwoeR4ascn32TEoIZJuw12RRXKX/DL/K9GzDTqN
LzysqzNJIHVYG5nvT17eDR0LrDLGFt8yslsbWE6JkJc6RIgKA7hRpruWU1zvdsic
IYPo3J44QCyJpmk+oHm0Tl0sMUDUdD6mfS4c8qBhrn0gPHG8ivzzQn9rJ+XIrJoR
BlJ3aYDRLQd2r1lwWt/FwVu20Fr8P6YsG/zLdSIVY7iyDEfrRsla2I1+6owzv21O
QwdIT4n7xxhq+ZEcrxpQPXkLEAMTWNISXPzKIb3YnMiqwVgoNNAFzyBqjG2kbuxq
0biFpn5ljSFuTas8AtqQq87UOWDvetQOfdaMFijBoqg6HLsuwKTKZ4yBCvRklKYw
aQkth8S34n5bjuE6xFfTPAKRk2X/Ka555JQU/a1t8XNyf+xntU+WEmtoIQUJQD+e
8bw/uQzl0AKgFfPdTBhXyEsQ6HhzIuF4Am+9GcOPB52NTRFPyVYqnwN8FF4RhEhq
h9+HFoZ73KE/arQcRce6uzshnlDSCBxpB3zb08v9B5Ys01wMdOMhqn1bAiXKO6+E
mrOAJRRdodwHTxUkJDYlkkKI219omZ6l1TFayn3mrCfNPPGlC0sUfx7m9n7XQYAt
3PFP16+q/RUTU2etDjZ0e0HYy06q3hk3tfvpaIeipZQA728OZ8UHuxtJSySVzfB6
Q17Efhc54wUUfyv/aOir3wqZK8yC2lX181Ifz5Tgy2SVnrUCjNLTOtYT2Jby5lz/
0/nXAhWJKZ553D78YIzgnsFr2ksZ9ZaMFJGMjfNUk+SzEJtm6OjRMTUgP4ImQ8wy
5ega6H/L8hbbVDdnHYa4SBRByYP3PSTCC9dSe7nia2XmBDxWLFBxDctxB7xvt+RZ
45pORH+NTLDvWZDg5kD67EET9J6fiyP/9U3RxCgaZY+AvHD6WfVjxnJ90giEaPhM
edpqGgog633kTz+5gtdHBxASP7tIh0P1eHfN0ZmjZTO0+9GtZ2n2vV9vf+gkrJc5
t067S+jjJbgWXs4/ywuj5pwR3zHV+C7NKtHTiFVLjYKWINom0237tsUZ/YP2e8j9
evCOn6FzwH8jgZMeh+DU6KzlGlDfwlKE0dLi6sgtcyg/CHKqVALyOilifSWlg1Sd
I/1JyjsMt7Dc2aSdV17juR0ZFmHXwWI2CL+oGRvDM/jPk+C9oJlwJfGXamkSf2sy
ejtKU07jzpuYzchlMMLxon/9RxZm3fZn38TYJYPupdvlGZvlBR1ztl9+PArBfg8i
yVDjyzQc9TgGGxbmHp8prsgvcmCJvIDfkrTH8FEb0HQ6Qz/yI2QmcJNLIL77fZcC
N5p+RjD3h2M5//w4qW6qAS/U/vz+F7vU5kk9T7WYbmZvRRkf10yYFW3hY3WKm15c
GZxFK3/Y0iTW1tJgaa+7+Tk9Ka6V8IG2NGh4mhvFU55j8Ko9PtpoSuZgnL6x5I6o
Am0fqbFp/lkJiBcMmCwPYUoCL37T8IP/fCmnfCvUFWzBnI/pR6kDk5Lc/ijFCiQC
kDipo6AroNEI4RMpAKESPmG7W3Sl8n4jFIxuV1eZN+/MJpsUje4AIaEW5YI9cFfZ
hb2Udpd17XioYqn7Zry7+6w+mnnrEWYLn66TLNa0oK3n/bzhZ4duX2IK4CsP6TNS
26iNig9JM6vGx8rrg8U4R+CUM9q/Lt0hq6wSuVQMCMBAl1TERHIicSc22o54qn1+
hA7iVKExiR9FRWEk3/YISFDbIG2Gtl20laeJg4Yt4jfgcy0vOzDKiuvFkiTcO0yB
mqP7Ix0+jmmeUFW52knA+RUQ+ng6VejMTw9EI7g3WFDgDaDqMUGJB39no5nDtE71
0fd/Cjwa1acnwsFt/c0E7vIIf/ByKI1CzQ0vJck3o+p3VU6GvR6qtg8j4+lb3RfU
s3NBbzkC+v/e1V56XE1XSV/8Qxt3OnKieSsTRm50dqRgBGYsPZCISLQo4lRz75hp
O8N5jX+1atHPOn8EzQha2fuOH58KKYj8/waoSFiMDwsp0c428EIuD0FZokLmJhAA
TCSFBjpGJJ4olxJOHkPAwkjE88OeyMsopa6BNC/LjyaNKiYBC/TMr2Yr1zPXzcZR
Hz3bXUJSB56dNSCfVjm/WQ+FfZr7+3ndqJLAyyKRN+Q7RFsAE6IxpslKNsF2NxiS
CfRBwTIJQtNVss64cP6+Lw+BU6Pii7Gc32jR26Y9jdPpDf5HCZa0yTlMU7qdu6R8
ixZ9fbh9JnXIHK3W6A4qiq5Pfoy18UDEkUoYa3nZcGld4EtxhdhO1LnTNyhpdmtw
hcfV3H0O7F+N4oL48IsfRvU2AgGsDK1Cb+cMQ9yhxmvPqRhiABsV19oOUnGoxPSk
9tk8uuikCBygVq/m8axDWQD2etTDj73MM32mcIS82B9f4QeFtOpGZg7LFwx/q8hD
tQeNkfvVQF7ZPEY8EeKN44uW73qixY3jqS4BkgAnfhwybAH99pU8R0rAE9yvX2Hj
bBt10SsiD88ZfLQKEKls0fZ7y9qtVyZ82LCCVnh5MACvfmB/nCkgt7yKJPQCf0sN
gdNt13LY1PTEl6I47DJ2EzsQvGM2lqbBVwK02JaVMMyO+jCT8E6EJkVwl0YsFQ/8
NCVc3AhR8iMFO0/YROKt5b1/oO8/6GaZt9T9onpgRtii1R5v5sWqXrwB3IgEGkJL
NSuNdnpT34YDDHQVNJyMfzWw6+YzlR+YYkxRcssw/DixjPicxKFFuCbmMnIFo8MO
kn7hbTuLXseMxegy+KcKVkOkGFoB501INJjRN5e0mOkC/x0lyn62udjP6acs3bDF
hNFKM9u8wqYEOEaNVJpwjegUvz39NWEnVZziKe12ee+gQMDA309kyqzxq1mtZeao
jWbJGjHi3wcQ0kGTmPO2dLUvVbdembl3Bbk5PFN9JCpLEARxuCkt6+ORi4V6o4Ft
1pEaeq8OUrHg+xBrhp4xyRNuEhr00QTVZkWu0AzpoPjZFwFSqRGA/tD51mHe3UGg
EH6k6YSRe1hwt62FH7LFJeiqDGcpg/4QxXhKMYysLdxrPXzuEWVqlq1BO0fzMlN8
qui/C5n4mmbF6EbIvsglF1qTzSgmZnpdR3gKpf9nqfRGVYFKgRw3WBbKmXTj774y
dgR1quoxIsUddkuJwNp0uAULQiiLypLWQa2inEmY392YMs4ywWZm6WaoJ6AHD7yJ
h42UQMGwIv5c4qtsD4GUsywNl0R71BsfCfCXMwEAKWTrkBNEvhOK6poTPD3YOclK
+q7PCwPWfoxFjGgtsUwFeaN8ROl1zbvG6y2N3utRRdT1bV1rCs5F+9//z9MJKrgg
HN9UQLzQQkOzN1VqxCb2s+8WwBJzewlBjus8pAR2/qx1aH47y3YRkVnrvfVwsmra
xABjfyeUNDNGvyL1/Dk9el18gwfVxllMA1FQMDm+mS34kkDBOPT1W3ODzKkXvReS
5kD5TIqGzBTvU5/V8ZZ5TFzjzIPLb9TdN3ELlLrTVz++xaRECvJqO634QuPRfcy9
Ljr9t5XJFx1O6EdLOUNnyj1B1Q01IAIoQYjAsY3CkTkAYSpOd4Yxc1bV2+XG7pc5
cGTqSU91Rz14ACzDn33c4yBoK3T8qv0787DK6Z3LT6P5xeQxkDRvtdXksgRKg6AQ
McCpxJk3iDhQMzFemfS19rkarTjnmVxEEvypZw8hOXe5eatLS/ThSOfliwJffa6g
ZOoAjkKVZcs2dUP+ABOxdT9z6bAi3fSgjdlFhcJhdPAr0IGg8QB5gfviB9hNjC1s
gr2i5SHDga+lC6JgENNnu9wEdhyTG02iD58HejzMNVACJxqGxElXio/LOdANZBMW
hM/8PCe3m8MzaA3ghvSrePqgz5pLLRd2P3JsD8oUP5iXtlPNfCrG46YzG/kkiAhZ
KDfTssmGOWFzU1O234r0kGFZjDcDLiKqDZSI10+Le00gbmNWlDmn9ZnPsnFSALht
U6o4eAwiN5Awyhl3JMdd2UQKG2VoA4rOwZv5eCqSeDWdXKDn0H7yHhAFWGE1F4MQ
/j6UkJpjYlDYp+TSCJquVIeZVRcuS87SyTYgdi9URDSJJs4mEEq2NSf430vBzSV4
L2WmQrSKAa1/rwC0UwOP/0HB/fbUvK8dWwd42Om944XTk0Jjj/TScLgUkZal5XVa
6/vg5tOOBDYh4j/CCpPkPaQY8Yf+oUKl8DHzZ9lvVKIQTKm6D1EF4bRX6LsbeFeQ
7fjcdW7DZvZjuV1Pu8/uyXygaie2S5kuOpjVDu976fUuG1BnGjVaT+itwNj6df7C
8iy1qKn/2YM8iXvS1Lf4WTmju1tBGBPRyudxE2Htlkmz4xOi3ZVAI2iJVq1mLEz2
fi5GcVG/NGrQdbjdFhfurStcqbopNby9VhxRDxKN9X9vijMjcvgN7KSNd5tNy/nq
IdFKHJz1EnHzTxU4UauhM8320az5KQiYd+7NavvlRpykoJS58ERbE3Z+Ygx0xWr5
vOgMvRnt84vFWM4u79e/ITnaV5YYfseKL5nlQpSdb9ZpUcN7CsQGPod3D8Xy8IBA
MAInpkZu8oxSUtZzEgDkpYJcVbT+7TNHNa9dGqgQ+wlhMM2bDD189ZVxpx9sjoxV
EbWITIbuR3CJnmzUkdW7a64Q3pvi0HkWFr/m3fF6JUoam6SXjGs6EW6RbaxnnvAL
ljzxlzDC3H/MmfIyoykpbRRGjIyu4tg7HrDBih0TydOOcTmkLCCow3GlJTEi80Zt
IB6nXumAFkCXVMIUIrn0kYCHe5LEODlUoKVfyg7fr52BPH2U/AFSefgMHf5lj5BI
5CFpl1v4CqaNA/BMZC81dbEOzWIOG6/ySDf1QJI/6NCfnyrl2mDyXdg7anTz9HdC
zQCi/hkqZSBoXEHfL4mbGKm70K1ut+r0Kiv0KWNb4AuORoqQUSbj30XhRCBNZU6l
RzEl0l2vw6d5gUTcB4ktG/r6JBHs2+GpEbS3NC6t/SDtpTQB0xKOz6Jn7IVlwFZL
1HDKboSM4dLa/Ja+aou/Nq0Zc/9SoXUanLZ1wMZQVgNTYpajX7NLOIJmU0k5MVtv
UjDlkFqRjwDOhA4n2TBCKd1SilHlxtJJQ7gIHz/gflaEMnvm6YyXfGEls5RLlIxj
Bu889NyKd0FuID5sDf+DFKcl6UBgQ/waCeVljq3ATSdN1B8MJ3SqoNWk6gdvu3TJ
qYS1BfpiV7xkyWcP5t2+6AkZLMctpPvy7LwGMNgOL4C58eB+85KwN6ySVck5RFFe
6/KGEAjmgduOMaCqoavWiC226C0KWMT4PWIsz+EDmOEA4GYHHfQswaLdUQ6gjr+N
rbgHBr4iifejyfS9hfIKspUFqWuhIKVB4xTKMBE1g4U3nPux2GBb5k9N3oJLZZvl
7bcv97TNjPNWDWMZws1Y8krYCjc8YXHantxvq+cSXCHGQZSu+cZgnpvRtGzvk7MH
i+BdnpDbB05vygbTnFUGsxdxYUXFD2aYI26WaqwPxaURjFEGCfUtx9epyPeA/Aq7
2c5/RzBeyW4wT5yxQnXeidnaTKBfPsXNVGpzEKW+YlIYgHaZA3Fzt/QEH06FXghE
++BXrCyioAu7Oi8swseyYeyhGWGoBx4oRmUIr4b8IvXusRjvw0e1f3vWQQoZEiOM
Egg652n1lT1T9nBXUE83LTC5HY4aOFQPlpI+/782NV9TtmGxgZDICcF7IR3CGywD
rbZGY/2P8hX1lKDsRb+NwO8bh/vkEZEW4f92AnKGr1NLGQGoFj3sXyBMKs2rabzd
77A12VhBsGQVcQxPg34czb9tlw21qaU/y4Cif2VhttBBALAnGOVLgSsnqPWKTv9r
qnImZnX+AvLi0tvIHfaw9fh4W53NWY5kCpcaG/qOyF/MrzkOqjD2lc5FjO/YB7Cy
4/8gFjhrkWQy9Kk9HSm+3zOPvnaI5JyBmQYU7zEV+rwYf0VqRHavxygH0YSceHg3
ZrmZv+OGRIZ9HnKZXa4zdKC/KUaEUhGuRU7BdFFU/KKEePMMSdykHKD349+ovgWt
gy4H7ycKYEymgTDn21AGzNe9gU8IaIH78JFltC8IqbmV2/IXKXmRj84xE5dURkj+
lcIPRZ1eZj+HkFEoN8MBtdtV/OMXW+RhTxsjVogrCrZel48IbnS9rkxE6Hdo1dzK
qkGi14KS8W4SX59zXM7SuKt5ukCd3JocT0n6gFBQ6ngrrZ1CejZvJTtNlJ81rVkf
GxX/LzQZ7+BuYNkSmreDyIJJ8QcBdtOGoQ79m3yzoXpkmGCTHlxehpsKuxrLgdAK
F9nrgAOHWeQw5PE6iubanu2+/3N6w5rLzmAb4BL8msrLTJheEG0OTh30QdkpYAfN
Cw8sA8F9wDGg4ahpXv9JDtSfCloB4lEIQQSci0mr8PMpvmdNSKxlg8XrMlFzIywu
X4bvnv1p6Ole4Ysn4XnjfIqh1LBcizsOExs/Fwv9g4P2YDCFvH+fzxdJjqjd2epc
Dd6JXQD8J8s1kJ8E0Y0Wh3RVMOLiTfvHXK5htJK9JVp9ZIm/eC9UN77kLK71a3Ye
GL2QcPQY61yXPuCBxtMY/cBDC11OWs5xAkEteeGZ0mhZXn5r6YpQ52GUWm0Nplbs
o18cCiT1oVfvLNPYfM4Z948hs3btHX4iMNf9bUHMIGQVRBUG20/oH/ViVZmkDHRC
hxOiXZYvCS/S9fpov4igiBE1x1BDXj3cqT2QMj88Ij8xsyOtf9hXSuorX7HtpaSm
cXH4+Y+wIfWkyZRjA215GZKvOKFyY1vPPnB8JbU7CxwLN8GfZaR+Tsp0yaZxcPmn
oVVu40PN9i2zlGf9C4HmXHdhkqAUe0jfrkBeTmBzJIv/v6oqHttCdmEmMC8H0T1o
JP+AMHWtPai6ikfkHvEyT78rvFAnwN4BjE0+vCrUpqnqW8EMxifGe/wVV36vsOkE
96q8USNUR9D1TozKFz89qyBTcUch6wAcX6IPKmjDMfdgrJEY2O+sWq2R4W9v0XUv
LfUjoM8L9tR7Db5u6kU82qtvCsA2+929uJ7ez5/s96qFCRfsmq8UXot3wIzNC4bG
ERqLG59nzH+0FReQmZ/gMEXaEuFGgkrzne0wvLwJ1o6svAn9Ulcekl8VAMWjkX6z
F7arOC+gVXl0d+1gPqke0l1vRZIo8aS2XcuEftcSkK3gZeEYaqkB7jj0pdDKNPTG
sqQZFHKM3NKLFweu1eK5j9drB4qYGBIuE5or5aV0FeUPVfeK7LJhmK08lDs8/FiV
0SBfdlV9m3CPd7vyG82h4Yr8WlMhvH6o2ETdZtDe03vt4wJ2uhOIWtCMHsqutChx
evVVme4p63Vm+tA5lxVhUC+0lKA1LjehpfkMoL6RynH3pkQtE/hBh4dAg26y07OC
3CMWTYdkASyo1NPlmagD27IyArKte/i7tqwCpnvqPSzF4oTA2+/7/4P68oGs+JiF
pQVfBOiQexXFjVVJjSeROjry2t+dXa+uABu+di9fyKdBmrx7knDF/FNMJTiTGNhg
2yH1fkkkn7sORGFJumLJ9mXKM87Qfk3hmOOf97UTfoOL3mnal5mNbPtLXIjbKp69
/XIAE/Gfh8dkwlP4MLSVpE44Itz8nwniH8GcqxOgM4zSfrZTELFmZ5jmZ2aE0Gfo
JHxsm4YDE5JwwH/pyaEtIqdDeFpJj+RSJY5N06qimeTgv7+cYOa85c0meLeVglVq
OQcE4fdzCYuiJxQiHLE3WDl9VAthpevloDuQweVcYnTfsRCZqI3BkHoi6eNe6AZu
lMJFYuLynX59pWO/daNL2SNDili92BOFfaphJ5JXERM07hlYJ+0ApNAKJ8lUQiVF
oXiR1Dd5UnfbAZQUBWxLoQl6ylDfeJzPGNCKasIjiRp0FMOcilWlqunxBlnbUyZF
Z9LRDAh/3sLiq4J6MlJhdwLqy5tWol3R5Q/uUH5e+fXo0DRSddwydDFJVBJA3O6P
vU9JkQhZ+jSkrRBLqIVfDtaVJt3beUHietmsFMG0napGw6IDe2DaLWHzU9qVcPXg
bwWZxXZuwAnx+ynFFriOEzboa46iDh3Ka8xMEjIDe6oVYycYpZ20zInACIt+gXsa
c5pGkdlM4JUaToJF9T+gzk+ofOWx92UHLFnQOSfPOvQ1cV3a0dpVG3PkfHUtixZ3
bR9MPFMKblJCNC4DOTvOJMftGylwKmJjgxZxS1BvdgjlFoJTxRwGXJh4s8Q9QttI
eHrA8cFoYhvWTsh9gJsE3UbIm6eXKz+7f/W85l5hCk7yUtv4vL5ksTePsteyFyjf
SA56I8FTRIf79vV4sDfipH81scxVkqV5PG14hdD51NJa2fF9qRFiHRjJg/lXtO7V
wUQBQ8ALGt4ZrQC/l34ZY8fVe18snGFCtjcmiNtgGrgeBxPXrlQXY83hjts+jVfU
7Xx2Ob6HCEoLfo0+b7d1M/PuZenF/zdJa5lXLb9JZgUBgpTy2tYKt4upvFlsTRq4
O4QidzaKkTtzPpi/c5vPVAz0O+vYLyTtKTm71768adPVwV34JWo9nUDULJJ1Uun1
ddhFDTYE56xfvsFT9R21RHh6l1XtcVl2a198cQNze53IFP5OBBtzPzSK8+MIizMq
n7p3fUnKpOomF5P89Mnp8WmQnmdN7abNaqMEm+iw7wsDVD/LTfB+QXURrAg+UpLB
sMmcoK3QzigoE8VY7L6bv0/b3wWwEX5AEShN8mcWKO9x0PGc3tUpT0D50HIQHvJD
fO9dV0MUUvOEVlBTLmAgMnlv0C/pXv6wmp+PaxW6TfnIDKVSBt3SlUJuLYZkcpH9
lte9/2jwHOBzKhYyIjKcWhCCwdMboSwAcRSJh/38rmI/9yBb+7bvUtgN0/104cN6
qsUREhBV8a4TE5hT4bsJhKOr8CGzbEAA/9mQ5K8NpLtKJUuJLaMhJFFJhsuvPlVt
mjkWYxUbDmMXIAaI14n+G81/SMY9h5eqWHz/dvelsqgDCSqhEnAFNTResnbqkPRr
bkhE8sb0yquddT1q1uSAsJuAYMoJC9mlzlcant7PWyOe0feHHYlGYRr8M2YDPWh8
sfjaqwTM+2I2OAcNUNfzz3Eg07RwB0nBP0nYT71USqO4Ga2RNxeItDU+4Uo5FtC+
7Zvqfis63JWqljPrXSaa01ogEmmKd+BCudJ9225fI+Ttj8vfAxrHmYi+Q1VeraEs
YhmDawWDUBeCBBn1IEDQ4UNoUF543CEYUuhiPdxnTg39RMY+4o8TTrEMhLqSDmo2
9hGvuLQHza4Yb7tlAvU857ntAF3izxMMUqCXMI6Lkf4m3SlgWPzVs+lORIZvgnAt
7wqrA/DB6b784tSqx7hqyyFWNkITR3S5Rg8aqBSz6A2LDUpMiu9bzX7e2zHaBMu4
CTwxrbMYMnf3wzCjtXQkS0uSNaZ2yPekewqNIoZFh71hPrCOh3tiZAvv70qDIHri
lV7YUVsFuMLbstaQBguCY93Q117a8xg5Qaq7Z+38e+B9nNDW035U/NEsPAV1FiC/
43XhTXAuHU83K+Hi4AF+LrxhNH9Z/ndj+3GzUsSS7u1aYztbWzU8lYo/KVYl0Ks2
rWv8rGnLrq3xZlRvRS6tcX5W/PRjNMlSnI/53Db5b68updUpE9MN+JTqC3Hr/hqf
yJV38bEZKjK+cSYidGIjOuIuOuuX2KEHKVR5HvOccw6Xsrs1ekwbGFBPEjiyMM1m
l3RbQe6AYaXu2cUC7k6KOs/Asekh+p87f1jdjFcePHWPXIP9yEmZUm2YPlpuYKBZ
2TFGRsEcdoGvkGKFK6i0As+t5ZMeUrgbKWoQWtsjk6EL9aXAq5y3mMna1h14x/Lp
8T7pMN6vAoG9b9B5r85pGQkxieG38rkHY8/c5zgTm6xamwEZFjjKmHVwWxtcIR+w
J2IMjauqDMNCAu/MT2Xq3O9Br+aHDjefXW7bJFWTQyERI64LNDe17JqZOyIUJol9
jzGJYWi43SJxEBuhvYnCbQjTRtHmt9zJqTp9dsU/Hf2GCKEmPw3YUonrBjXYEMBP
xc9ZWbprCk0Ul6oBMMl0sNSc65q3B+6BMVvocfnMQgS2jdPUTyfsRn+Dypj7jTUM
HL/sh7MrlM62+5i3++M6CYllM6IQ3nSoDPR/4LTVvqqG0i3MxZMeBTNP2aeVUR/A
OPgDY8HHy9sdFV10zBxXU0TDpzhO8xtl5B6U5ve8ek/Hs6jNAYfRJSrb5ZPQ52bs
dUSDYM6EbcDv0DWaJGzINdUB1dxZT79dqaJ4Xn4zBkfmtv+5ff2mBMn1qdvqH/hp
HuY5LIZO3YQV/OfYgqbwHewi97J7hkTDf3+GqiKywFT52gPid0ldFZNN2OxH4Oss
Il+dBEq+W0k3k39NS+Vx2wOm6HsDVTpT3dJg/9qumsDqoturj1rFzJu42H6fmVF/
XVH+pr3ZeE/FgdHELyVw0RzPVxGB0r/RCrfmFUUgoUB5sBQgqYGY3HEtdoQZADjJ
31CiSz05SQmZ1NJKlpD2AxT+1xOGp0azCuxxK1SuSzW+SDnSMNHvUhi+0jgbWAnA
QThahuOTzhupwe/a3FY+tNoFppOnJu5gQnErqRWiM+QzbTIzyizP3luH8fHm0z6f
0IOafByCme0jkaT/6qYIP+377uOcKp+2kuMqYy1VuBI=
`protect END_PROTECTED
