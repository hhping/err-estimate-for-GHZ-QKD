`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5R3POIrrzjF2MVJRMqRTvN4RB6myO4O8NLG3Y0Y273IDxsnuepRKHyQRmhtDNJ49
TFEZ4x1q0rO6hszmaoKNVVdeKgxRaB26i1QsNyywpJVdg3MUDRUIAAsXTyX46fCc
EQ2lsNA1Mfv2kR+XesBK2CQNCe2XC6Gm4wIjcfsKa+ipf1fEdQtf1j35Vjpn8zTQ
Fk21eiuGu9EWKBQYjEsMYIpBj5HW44Hp2Ny1ixKz5b67Rw/VthtnSwqr7eBBxB8Z
ZAxQyyfrErz1x9bUaKS28EtbHtkz4qsFlycviOXZCtSE4CqhSyTEhNfJ7y+WtstL
iwmQv77NeOVRXN5eJSYUdd9P8HUO1blFStjWNGaFL7qkPpypA7MtSQ8eO8MKIqcg
KQ/BPEgbE/KHtx9HtpfjwpKuW35Ae2VtmKUynDqG7xiQoGoXUp8ljXxh3NrSUuJn
8DFJ6DoJuRWR2AIE5B7ti1GNdjfABwXdgE0QViPQNtovUoI/oewb1ALTfcGDndVT
BYzmBEDZpybD8wiYVV9j0kMOtVH1EDccD/Ymwsxsgd4mu2tiwjUi6wGg6S2XmO84
85Atzi9NvCyOZxhCFdapgiDsxzBlj0uuSqb5D282ThXXBhDqYZauokoMDYTBuxQQ
Bp6RBLVh0AeQboF8YY358Birqtpf3CGn5v/Wu/405FI4sN/OIgih0XXLCFwC/W1Y
N/2dME6L97AUyUfwX4rJlOOO6E6H4ToqHmONMuGBdXH+euGIt+bXLnyD/nA0TfjK
6qHu+j8yOqvWkE2omYPxc/lgeBl3RfGcP8alLge2MzXH0kFbdqGpyQxzZf1/Gjb3
+RKEixGucaQ4+hUqXDshbXjT6lUaUN1CM3dmTv+TTl6EOqCu0dvInsPa5zA525pZ
gZZSBTIkQwYo12sdAaGxHSDY0lVQdhIYEYkGBBusC+3fV0mQifAh1OJu5mQDS1m7
0gt7Ikzp1mGW60xU7Lz/84dN1S0PyKF59DXCjMmi+nzjKtby/McvEEpLl2mi61cF
ycpH9Kle0vi8SbJPWiqqiFkRVEgCTu3X0RenPtrLmWdsSH1+cLJb06vr92VKlVuM
8mS0bajzxITmAePw+WFUEDwIocP4/oBdO5hFR6QoUXkfVCyogxAZcFLytpRCAgAm
xNUzWK7uJYdKTHNpsmLgBc7YUDBl5TEYKSkcfzI+VVKgayiggXWc+rJWzTY+Te1K
ZSptz0Y9r49GT59q9qdbD8dV5FRj7xW/ricHEdlVSH+hwecN5zpry+aCyRsIlxF1
hPg0ezxCvY38MDCSba9iq88CzOBcC4mZTRXXB/jVTE6GcZupht673vpM6tJGMzTw
rT06ATCqPFIH3Ch/kCRb3LmEzsMLgh61Vqs6yhAMzxRJd7k8gclrxnwhicDtcgQp
VVdt3PU29m5klgoG/lHaQX5WGKw5Dz7lAh4aVKgrb9MXt4YGdNwPi+mIkXecnybV
7N8En2C0QUH41x30zF3wKjHDorYgsYx2T5yI+k7b0HwzZglv9qMH/U4I/ZotVUv+
vRi0EAqNqP6f0QU+V/q9rw==
`protect END_PROTECTED
