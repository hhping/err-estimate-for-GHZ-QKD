`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bAfVDp7XOdsikSuq3AmBa0RHG/7l5k+Zd6aeqLFMS0GUBFTKihChsr1Itg16d5cp
N9S7wGAZIPGXezxajSzbF+uubm2nZmnoqi79tWMUR6wbrX4XH8ewVeqhTxx4DWbT
apL7QJonuboNhMBXegeDlVypR30VPKJUnCIgmTf04yP/F4a/TrPGPPm9ZZqBU1W4
aq85M99bTQt7/JZVAYDf3glxNicLMBZHRUTLuOL3hg6+d2cpnz3cEnS+5PIIyH+M
EqWq9wIJ2pvPkHIXPZNcX1qCkHhLgd82wjeeIOMOJsiDfl5Ms83YmRK2A/pansed
/x+brY9mzpM4MD6XUl2Cjrn9vnqDFkaN4aG2UZskSf0iHanixFa5SZjANitiLBgT
VJNaSEKrqw/yQxSOw1INWCngwHavvUuw4mWWUNm9VsGHRHX3E2PNbeoeDhJP2Y9O
4cxz6nF5JXkzJm7YRONe6/8TnozU3UyIKn+5Be/XGPB1mAIZw2WmChaTvKei89RK
++KngORi6BK5kiv9V3PLehF4BQkmDfxysQe4kxZ7tnGysNsllr3aitwgv+nvtjm5
aEHRG77tmEy4c3coN0oTi1BmQtuAZzD0MyE0XZ5B77US2rwuweoveQFk2EPLODbG
/YolEDaL9xI4etE/foBOQeVeJD0HVqxS+WEtQs36BwfhcPnUORnuXrqr4nMdI2HV
7UDGyl2ADskc4zX+9kLh2BM4Rl7p7aRqOign/BUyTmJvI2SniHq5rA8hmWDMwLTJ
2gkCufZutqthM1+xu/UUgrXTcewEVKEvJWpIPPEdcs+AfgNgkX2Z1vxLlTzqyZB5
CpgiFEyx3Y8POr+6N538B3pHtB2Rrye8TctKCB3TqvmgeH03MSNi4BbFezTJkXTg
cDB9IOqzCzGY3T9cwpDvg/k5Isf81gzymiUyCCrFgz9hUrC8FLcVUXLUamaHDxe6
vKOcpxmWgW1IgIbps6vVJA==
`protect END_PROTECTED
