`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EdfnrDYqHQkBRxhMxGMGG4x9woe9r1Oov1oVLdLZ072WCJEw58CquLH/44eXjuna
cVjg1yuh2Bnsn4Ii36QEBnv8957sIJ9/ySJCf10gO1qDC988wMCn/W5/2bJcFsXS
7qyFrrgMVSjv/ICNIWa3erB8Q4EW7qZb5rfBbbhWYbJMdLQ3ljuCLJurooJKTGtt
mO4w5mxqyHVRgpqFVHQJkMgy+MWbt4YhELVgJmqCEMdx+lSVwZvwRNiwCD3CqtAR
ar6avU6PufXHmHaar55e70gr4GNQOqoYOORQsMFPfCgMfO1izlCfVOtlARAr1KBr
Nxww7bpv/mRfRbG/XZ+859E65pxQjIYpcoHFiql+zTQQD+jd5WroFOKUW4qnQ3rg
agtqNYNXs6BLKJIAAy8lEHRrzKYeWR6fjK4TUEdls16bBmMPHgylfI06pBX3bnuy
PCcCtXkdesFkMk3NZ+YCIueoHc8QbDlvfkUv+VkLKUBz1VLS7bIIFd37whRIy34l
2KooJSbb7cdCMxDd5FMNmlaqE3PqmsPNqvw+CPyQwv0+47DcSzGpjxpl+I1yxJgN
qrx/4lTFdRQxXLDkPqq2lswZSspOdeKImZkdKVC7dfVbPg5AtOR9yOX5gNXo4Orw
/abdSeJqMXIEglGo1pu9NXF5t3YZM2F51e7nrYntDmc=
`protect END_PROTECTED
