`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y9sUytofEBJXyIYGmuPxJhqBW6UGvy4J7iEEsIa0o10cFpTxleQNeGKmTCvET8wA
uEWEwKgfsFADVEYkr/F+SIA7Be9gy94BbCSMA8emGZ5U4YdObSof4uYs3i+d4bO5
Wih7f6XKveSx/+tCBvZI49bbyw/4ktMoiEJF+AoFQEhnrVKIJn98mvTFnX4lLqmF
K02SZu1ieWJ5WtXKB+7oznEBZzw2ZyyPZ96JWGqv9iH/PuwS5AEJmeyLVQlmmdEn
8IlAdmFhKuveClorCPV8O+7ikMuYKp8QtqvtsB1nEFRBe6xlGWAc35QRnsRn14Vz
mTY9cEU03Lom2ObTv6KtS5b/bKnr9ClMwnXAF4xQ3QUgR6WKad8CqKzLOQPskLOZ
AYp5k4egdQpUN8BgZWnMPN90vv/+64nj9kZMVmwKosqdfFk5Pbw4U63UDr04SVnJ
rfAimglzHyKg4KllWvq1KgHupLc9HyuRBxlH+x68IE4s7NZ3inRuvMBjKviQZslg
5Mb4ykfDsFNrQc88iBrxixoiVYoa06SoBzY8PhIG3cBx1JewfJrrEiBQptMnJFVa
WU+cOIvurkwe0oeVS8FfN0onElrhRcqBvn0i0OZOFRidLjmj8hKxtFINC5pGv96Z
Wuc9Xmkp/cJBRRwQ+x1GhS4A0vFq7vXgGpoWW5YXM29fZdQmrxtjSQqGlntG4dHo
WmiFjMWphePHiC2TqB4mNZ8x5Nnr8jOMMT1QhkKmURTBnzNLfA5mB1B+6+XJ8IiR
Scg+XifD/C/VfQHzp187L0G1un/tjhUR4SaY2AXacyLc9VW+8jCc4PuUC9Et7cuh
ko9Q3/kr5HRozEoNGPZ63ePY3k9MT+TCA6OsNX3CLEAGceStg3EfodsRPaFfslSQ
LWTxbIl96d7Ghy0RndtNecOJ9D3iaxdgzNOAWsvYo7PQtJwyqpsIkrRH+0FmjPJ6
arVszzTdor2PqCYgeg+k9uTbrrPSC/PWwpmz5PDh1mTwJoGx2C2XU2U82TGs5RQG
RFkCOAQv2DnaCdCq7YJryk4PoD9cBO24dAY4soRWiys4x3cuejfFUZCTEcAK3uuH
NJSCOGlZYICHFY96j/AzioBkm3kGiRFACuQKPadvt5f3J5+fs5PmiaCAxLMhdDfc
PKizomD0lSqv8u+dEFIFfLx1AoQD5l0VzSH/7EcBkHSoQGHVNj7VPLG4RUJ4BbGQ
bs08qIRBBL/jghwT/Ym05sqe6KYEC10/oJgeHXBh5l7V0/cxROeFW27kNqYSzhgc
kI11yVN7MNhiWMAyLPSdz1PnTgyLjhdZYNew+SPBjiuxuMRQiXu+UqQ7s8kM+ho4
5JzfQ0uHB2Ps5K/zo97Jw/M5iNWDP6Fz7lxErdz3RZnlvG4p+XxoAgNLyYuVKXuA
+8r6yVjkGOlddRSdky6iXA4weiTT7oO4VmKOgeTDLLJkJk21wCr59pQ6BRfggTGF
d8UC9qntymrKFk4Vq16/eipUIwSdMAr7yKqrcx4ldETEtbSySGXn+RcKXtUzf3OS
llML4IIHf+Ke8D+krC4Or+SpwMIm42CBehYWF/cgtp+YOG/Z5LuBmUWY9UQx25dM
FvLKhG7eAVJzJ3RNROsQ3uukhYe5u9ePO0VTXLAoF2sUUpqgT+Xst8PTZ9ztBPL4
R9mHiBE8nHKKua9mxajdiVcbxVRmtV8OZ1OGziuEGrBxYTt7nuFPQkY0eB82ctBB
OOglNSHUcloeNWkEYTjrepiOQ1mjuk9ARQUoNrUhTWNp6p8DYZuBloAx8mzLXXYQ
c5JDNIGyBeSmJHbSyCbEzMxMttdcSiGUOp2FWgH1BtmKcBdHFRCrhWiVSAZrHC22
/VXqmFCP6PeEEjoLY2CpQd4IywEylfSsWc5w354P/1sv4iRf3AcCBmeOGrvOUrHb
srqgbgRnUxMjt9QZcexjv2SOCAVpr5G1hGEm+eX3jxftMGqRrIQxRvGgQtcycrik
H1OKP9L0cRWmD26ay87Xn2yiMN9Rbu7aWKQKOsBhMh1CMpesAXTujW9noE/oqgSQ
JNw3pPoP3ZtX+GR2bRkqLcwDK4IK/rekR7fp8vNQEDy0YLB8LXXx5BMQyJdQLCGm
`protect END_PROTECTED
