`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JV00zOfbCv+dWtBQ/jPEc6DuyWBVC9jawlDf6MGbkQ1M9pu1fkfUsp8BkgQU6lvR
eGKkXCUnF7crYmLnUxmwdb0KMTdMUzIGoUZaEsYgwvyiUB49zWREn50Z0QhrZZ4z
mtMdUqMxICCV/Ardwz2HGyX/FUl1lvixG2XaiHxlgjVfy9ebID+r3TCZ6NQBdj/f
b9wLOGe/ao8XxTwbk8CGwXAqZcf7LTkwm5qaFaWxqV+MzFiDR4AGWhme5W0qRT0t
99IRFIAtiSr3mU8sVFvBxEGNZKfin1r02Wg5B7FagjcvyE3xbQjRvUNUm+ylFrpD
YZlIfyrZBg/RVwYTitKt1pz9yGoWENwKczXscEFD6GVu0WeqT777X1z6FpP3aGMX
AGlegeHf2UVjwSN1LRVSPhfQKfu8NMOT1z5r+6OHGwlFo9fr8YTS8TS2sFcXqNdi
CAhfty17h6ISGwPjh1+UiiIKVdIAgsIy/M0jZH1jnpcWwxBBhlm0TantAR5IbdaI
rFp+K7dGv8ifIjboFwIyir052TjF1T8r5a0GKWVs+SfWd79d3go+hyQsRr2wRCM5
0bc2vlmLG7y1CkMPYImIbmTGkZlyjQAtTvfPpiiDP7Q2YflvWdH+XNA1jFIh5NTo
nU/KCSxmU2ente3C1zZkwLgfIp6PJRMvl95y6TiJTCYrWZfJeOnigpGjoQ2i2No0
AzTLqdPRRYpHzHFggSncvvKCtyq9ofNOj016/Mm9nifDVmyYVszttjZMV5TV/Hnr
k/6kFULS9R2x2Dxu7oJZtR2FtzO5gCe/nUW8Fv0FfLgMMOc5IHhEevpiYxe5FGFF
Cyu7CIVw6e2708Q09+FxfkcaL2Zk2EdeETpUZKJr3Lyp5y25xI/yBu5vmGOlIZbl
VQf0cGi8nuMkYZdjDi+hAgIZzkDRic5Dl9M+gYsgSyQPWGhvflAzb9esOb4X0XEj
`protect END_PROTECTED
