`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DIWFUk5dOn5TUO3ZTa7QFvjR1SPnlJh/6xwEhkbbF1rLd1x4eIQKdmMv7TVwofb2
qQ67p5STa0Uy3wApRnSwKS9/LH2uKEqp43E+P544f5657TN2WfhFFkuOdtM6mV8p
Kncem0xrWClvuQqANAv2H3TjAby3b/bEEqOaPwKhOqLl7sqLBPxfSD0Xc3ra7T0Q
1mRNSzLMBjcR47Nj/ceRt543Uk4YTs4DWNgtMxse1am7aI6hOU5gBjJsm/xeooNY
WygkVZExi0rzWLgsVl2eDicarQBQcLN3Fot8CBdoqlFGfLn6I/vHNYIzTXkgdi+D
nhra1mebVARaGqYXyJq0e/yOJb4qIfpKlIjKFl+JwAh7gaObeECwcQ2CZkB1WSA7
s13FQ3MLjbTOTCYfrF1Wy4CFH8RDoEIymcUpXE0SvBkOpYN3GjK6qL7RZJ3zsTVp
WBOHzdx0R60cx+/MbQTXG/N/bZZHMhulu/HrI+/o1lLo3A7vPEoYVZ/zAdbn9tus
uR3h5NYRV2HAIGwxA+92zVCce5FIUdiAIPn+DJGewZlQQeap0cth4e+UTm0AfX6p
zQ5CTmMNlVRBvfmEZja3R1DSIFdWLq5Nxqt4mngv9v9BuHmGR8ij44tC98QGx7I4
fs6qck5TeoJd48+JEIsWoOznBDqphErgtXljYj0FU4w=
`protect END_PROTECTED
