`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xc8i7pKDzZicn2DFWeNHobbDnBHfKTnjMUgEoLdhZKB+GXXGD3xB2eYVVPJvArOt
MAXzBsfolbpiUtScSj66TrNoQQyUW/Mx5uNWHAjngKuf3vIY6S8FNQodinsx2nG7
izuQT0EVxvRBePgadH7R4bKeLMZq0gQZMPj3zyu9xThh/L+p/J1d4yOGogwg77a6
NRZjlR2fSdHKvuGBG85bFjL364MubWrUuK/2MkrMct+wW2MTFPARUW2cwPR2SGtF
fUeqbMH3WR2/8KcfhB2Qn69gW6lspRpIjBp4WY5ehtdi1I3BA1LWOrLKJ0OArwbt
IIk4/uZR5hcxCgBERGVzQdA4RjGS7D50E9Kao/K4Hv0NZpXyOG9AzE9RCpif5SA0
e7mOXjhXPWaSor6chfHTc+eST8a4qGdQs8PmkQ6dEhzkOP3TDQewDmUv3yHFVoQ8
wx8vU0vez8NPcf9tEImk/+NtEJEeTC5pQClEHNWwqfFAmNBy8rIBpL95rMpGuoND
OdRxSy2wvcO/fdhD2gtwML6XziDAh64J0CPby1bHK5ICs6NaaLTQHQOo1SDsheHm
5L3D/Nny5rRhXBdx2SNKKQlY5SkFMCQ1CG0MBCMPlvE=
`protect END_PROTECTED
