`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1g1AgaVOO1l47TENhXdS7/fF0ltN+UrP5JNvsTz7PlhyRRyrxf1bp4frtkGZtE/U
+dV54R9ezPLpZ7Ny1HyErFWrFPwRfFhmyK7ZXdFXikjlbHGuUKhsCaQTPRyz+PmQ
75UCAcbJm5URFG91nggnROh/NEIENJeDyUeqAAdK64HLZjYdBBaHEdBYkofI4WA+
Lcjgnlk4CT//pmTdKe8fTru7FHPEPT091Z/MzGEhzY0NVcgupFOFA9XmUaEVupC7
tfaYo/5hiZMkNOQW9g7lWAbnViB1FED1bMIF5RGA4IPBZlc1AMmOQGlTfIB0XYyZ
J/5ZFgTmdF6fNwTEZvZPH0dPVlpUI0Obnyoe53sx7m1U/pZGcnUtdpvpZPqd/Daw
1+AnWPbXJ3ayWvFo7tpV/fmpXb2ptOLJXmKorVW0obp90oDYcMrx+mio+72dwPMJ
zU/2Uz9U61z3bxrb8IT6VA==
`protect END_PROTECTED
