`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NFZExAnqphtkTUQigDeGdED3nY+R70PWgEfYjGYAa8u206TSBMYXKc+SUH04F7w6
3yZFVbn42yn6kWqb/yzqMD5DAsMfi9tSgAeDI91p2ilpSNPM3wzF4cZwtYBopkuu
+UPB3FPd+DZF91usKRxy4jnLsChuX/jaTclMPmDfczx5SVUf/s5136LI0brELFc8
iag6u1Zy+VyBkmwmUuoLC7PdvY/EXksHArr41IEkmDyM1HN2iOjWS0BmwCA5OH5Q
8JFEFzjy7KQ3oJDd9QtsBuDyb35wJk36ld6G39Wz+D72kjGtjKc8rl1DDa4qTn63
gUsP3akeUIuxtN9n7QBP2yM6sgTDlIj0ltZNTCS660BzNv8kv3Mfl3QexxFXHmRi
CEqCgtalEnReLrlAF5NQ5yqkarv22dyeWnBWKJtL8rxIr4jAs085UkEeMeK1rpMP
Gbu0rXKjILOq8B7SxN6LEw==
`protect END_PROTECTED
