`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dDKxmNh4qma61HDlUvZaNw1u0xF5vvr0ilpXJWJ8D36v/1U13LqhzygRubzxhyUf
nOM/bNP62yHg566wPYSKgVDYNzYD9oGr/27Ad4aurijJJ7zazv8mo55G/fzlhOoG
p+bT547AqzJPgp8Cq9BFrgRxMuYlN62iTjBYm3/seSebRIDpH8ZaLN617az3yaBa
ncITAMdd/5yzImHoseCxr1CB/3MJh3mu6yCXbI19GUynrdtAmgt+hBQHoMf4CMHE
HqwTcOYKhRFScBhTSVMI2Dr+s+rbwYgjBGsO4n/Vx4qX6epKkwm6SnWUlqEU4efu
dKzZ4hGCrDNh8F/avyVnHwirK5ADtFwYqM4SuZtQ0m9mUwbMD0z4mowNYri3fpT+
yA/HegUl17EtZmjZHRkQFe6MqQGcb+XqJbNktoI6TB1hBoxUMv4jp90B+lt2TlxS
7DgzlUCgrPGsRaxZ1fkKjklbLtjXzzUz9cXyBHvC8epUEj4dLNJ+szOOnk/TokB0
bzdVK7taZIJ2BbYqVGIApbxkRzd4wBnMNgzjgjY9MYOLmFSILDTBh5nH/ZkF/sxc
7oNliRul7e2lLt3RO2eEnLoHbkTaS1DlJQlNS5O5uP9TqpCMda8WTy6CT1CKFq6G
YcgOdiHjZuS+UuNKaddC1i9qW5yqeM7VDsFsFDWzFmx+AvFdywVg1yRUXTHWYuLA
1ThkrrPXomoyWst1snybKx27q5pVHjBy0A2bs5inRNkoUe0UdhR6br7TUHkg+JR1
Bbk3BIAQHxLmtFTZbXU3l4Eh4KsGsCRgKf6N70WM7LQp7eP5UFHL7HIcun0Uj8qw
uQM0IdpmoStbpKm56Jx3sSOAFDjV3Xcg0DYxmar7hqe/+KDcN9mrEuO7BKlrXqvj
axgGuMKZLSz8Dy/gXS+/1RauGm191jRQwpGoLkomuiQ2C/CBf06Y6trSJveOfV8p
up48Mq1Vu2e6jrm7oq2qVvJScFpvpGuzAg5JpIYHASWeaDad3uoAEgbvJD0zhUrh
i2GWhf58yVTlx5+TDSAG1U79m7dv47KiYks+harRZIEkWUUELMcmVieqbSJ8WdE2
waDYRf6ytc2nmX0LC2DVCNNcWelqDs2jMqbxHK8Y6PlGuEj+mVeU4Ln0QLaAJnOe
9qXZqEbBIC8DT5p4iCQ/7oB6doUnUl8hjTxDlI4uLasHETbrj3qbOeDgfKnck4zi
syfddD6xORtNzor81QM9X3R1FLEKBGZS0e+brE3lR59URgJeIXhUd/6/k4IArnNl
3cC4wXOoKpsXXWzCtL5Mil1cpjY57S/Mb5KE92/A4iETNWCrgGmtUQvbneWuHNTA
i/bDgmaRpHXSXzk/IKAV3sG71ZJSHrrBBf6JEPwIMPWtgLtI03tllyeyNsrAwEPq
LeFzjncIal7zgJ/9dcU1M8JFkD8bmko3783+oeyBgjm9ow26xjnQv06iG+/hQP6K
knhvvtrSXSYQkODS+mSOt/JI2NmDEXiBi5fE1mL1zWlK46gDMoYxd+oixaFzd0q8
Cf1o/Nx5eItO5aVLwjsKExGFg300R+gO/cwOLUuuGWPMtYjViTsOOsbx85a4VNTR
0wPwtlU8cfBr7jIzXLsvNVcY7kG5fGMcLzHxerjuH06CehpVBjWtEYhSCdLWKWtc
Brfw52LwFk/GpjZJaTdn72XWrtaEW3RbBrpLlgMqxD9gpnYQSHqezjtThg1XQles
kbULrBwIPXGqibnEKpX8ybZSy15d6Gzr9B/nBF63bq4eX8w13PLEkHP6X/loLLUo
j/99YG5QRxVBtJF9ncynFixICpO60hoyyy2416ETcvU7XBxIDM5rbWlri7kx1vCc
v3G0Ofgcz5bEvckuUxFF7CwSIJVN9JhB/zRufTwj439EFL28xpFZMZuPuiix3E4V
RsnP4nTlr06odiFqdabx982MdgQHg9AHgsvFjaAqWINiqhSYtPi+JiHh03IvdmRm
HCCG/MNzpJJBPioSpePKM8tFHDrO6/AD8O8pvK6NPf3s+TruBqi9WJf9HjcxecGA
B1PRzM3NWqd2uw25gkLZ2T0ODLd3vJ79EIj51V5kyL7e1aHQEaCvKrjaktwAs1iN
uSZVTZ4yrRJk5jAmGxVHvzkVuidO3Zk9jw/po//ChUk64vH7aWSh9fDYQiDvnFnH
cC1NuZh/0bZGNmNhclte+tHAL6dDsxq8ht8WUFCbKoqmpvNtdIf4EXcGU9cNqPEH
woLeFEZWs+SMssKwBq0disEudlDSeugjfYwOE4Gg8vDp2/F5nNaElbN7TZUgrk3f
TMSl+q/NgchUAvGgCHEDmsOgqN/sey/LdujRx7QdVCTG+vR+CVlqLLtVp+Y3aXbx
1EoFCeEfqmMfz0Oigiqf8JDT/AC7mNto/1s4vi79nmIfgkAWRbK0L/Ul1Xocqdwh
xbIhFks9+RDbqWrYogxPmKdONdWw41LQuVTZ5llzBwxu0kXIz88wkpbstyixvrUQ
Ra/Om/Y4Kkl+5xwOEGUIuwW7y5vr11sKU3zByXTEX5USKJ4fv1Arx0cN2ffvxoas
X+sO8ZKJhg0XfTu7C9aJ0F43wmcBapJJ/xlV6dH8sJZu7jW/XkXDvtiKfGsS6icU
WFrNmD6mo5XAVB1wiHhHAw+mKJjaOku+q/hyS0fi1+Fjgm1qEgWq54qyiTm1wW4J
MSrXS1SevvQqMC6R4RTmkoQ13BiUYBG93d+hdvB4xqUm9oZY8syAMe4PbUEX2kvR
ZxhuumSefPBU1KWd2JXlWJWa7xj+gj4Y33xVs6+U89cL/ER+i6QIdTXpRJpJR6X2
Ij8O4yxOOLt8xoaNvZWxvUQ18esKCGTx2jRTwYAiELflsWA5KhRroCWP5+5aWcSP
6+dSIhU7xACs2SPPMng0Ja5WTyOhmNlt+3PpdGpsIZzWo7ZuY3DYhT0XvzG0kuXz
iIaDbNlRApo3nLfEmrIV21lWB11gVPMDjxYrVm08DObyo4ah8eo6EmVBStZiaTEF
eZunqqiQGIMThAz87lMVKV04/cfaeAuUxV735p8lbu3JEhoq+DIUFZ2c7uILEi24
VJ0FVvkPbfR951Zhb3tPmiRV6UtiPFM3E3aAyUzZs2NnHojRfW4zH2rLSMbLbsne
b+rT8LO3WXeZcdjOOkuBnWVKKCuHH80BZn3fgCYa+BJiqKA88k6Tc9TOW13wbpu8
LzfB3lRE+GdwHwU23mSOCAxu3SIjcewWUpeE8ZEQ95JUwwn3cv9nmDIM6o4lP+Xt
kSnP4iJutQGtAX40XNe4aSHBLrUwX7P9YU/15AgtFp42s7D3O4Ihg/Fo3veBvrhF
lWs2okOsQw8qpLnxWKiMNOZuL3UG9DKhbpTU6mYV8iHeoYtTzbTYEt0FPaNx/kzs
OKV8t6xuhFW4iWxnQFfPGInndodcuaKxoNRRhN/iYEUCmKpJI9uuDGTiouT7TN/F
6Xrt3k3Ey1K8z9ep3ctaZKYInVJoxxV1eJ5ha4c8ygnUyKRudUj00UoqjD4WQxgF
0ScEgXkAk5ylb3Q638WJZBHbRGASCV4e3OdupIf/xkcAeBlNnkplnIimG/pgCG8+
p3k03ve0FMBPpcafiyCerRFK8ZKNp34qqy5HbovBRYpbaeVk2OqUtBkM84lXMtak
oRNtstbG8rGbPn65jvPRFb39GTjs5ZFV5hdPpGBgognUc895PaphFtnsUrj2YCfw
OJLdngeCgiPoDIr7y9ywBU8XoTAM9NQpa1qShEFdEsQK2/iLyZfNsqWLhXBG4Olf
dW9wj5AWFy0N2UEF2VxdBuThMoE3XhZYXfxRJKMoK+6fzpa4amSYIIIPujz8oDbA
Bz0fQAks9VnE6SR/PqW06qcVzzWf8VbMTZVxGOZMl4AsCEfopaBVWk1pOUz1L+vg
3xiIoKvBOyOZ1CDl9u5bFMNnXQQY7XFgu9GRt9o3CL5DfgaDENI+6UV+nRrkSxxK
t33F4k3XEIJbL0rXX+zYyuzY1xxHT0rQUoa9OH1sSIlO5AnQkEQ4Yusj2rNrK+aI
2vdq+mPF/FazOK6zm84wxpenTHusnxvc6bVl7HWwWQCcmLrSXc5HPZP7CQqPyVKb
gFPokijolwRS+r2YYC5uwKzO3KUMaGzJmacXWBAUxqsPrh71Gask4SygLzmG5wWD
w9OjXBMByQCEitJGAoDv0qrUJnsvwPHIFtIqxHauLQPmzIpoYJ+3JmrtT/AXO844
jeiea0lOC7niuNYBH4qdABQaS31zJzJ4/Onp+V07pTueyr1Ilu8yYcq88PFoC78r
BnpiFh7LBY+2qE7qenKSNZDDT+UDJcO1p3KkqV6vyvRhhx8DAGSamSw+l+88wlr+
l/59aUWohXGOHKl7qo8PFTlbbMnNYOPGbSpxZT1qt5ZlCy0J9AtANsewc+fwnD7p
kFjx0idC1f0B36k0e0cqaXgzB5hUHwVyVdIBvykUqOblIOevWmjCEJm1GtzfoDI3
v2cwgpUvnZsj08KCCfzUhnCzU7n78V0aEik/u41a6C9fHq7OLIrB0WqPJIakciit
oWqap3YNzQO6QqWf5m1Kf879i/2MMsGoR5KnBnpL4sIv9OuLU1F/MqtxeZiNTLZu
sfOhblekfEFpqE6GQyu5GcLj1lWK2HJFLvnpqafk+oeTqA+Jz3D8naPx4Y16GuML
o9PZ8MfYmmI/uNaKx3IY9NW7rkW5ig/A7yiuuyd+iGjkMbeZYXs9bmiFLH3jUbLP
4yhCUlsok4x1VzwXC1W0siuLRQWkEKz2mgLLf8qNFV9uG8mJuyO7KO5mf8/zYF3q
5+mGdwYPkYz8ZHgEV+1TRt/hQWzYFZYXDdqSBlTmZ7IDCjtUjouejpoeiJQHcFqp
8awwV06AVGlRcOmfE3mFa2Estq9I8oHAVwkof2DlNjH+EgxM7jaAT8XN6jAoWrjs
PbR4qNzFccOe6IwkNbbajN+bswV7lyG2X+60pfmKmmGSEa8ug9uwSLLsPzmW5uxM
pftEbnPrxPjPgBqe1/50+/nIdpji2jmkhLDcO4pVP3kBVcw4oyljzDQ0JqJFsMuz
DlJvon+xYuB9xrGUgsf/aqUqH7snezs7KDecEzPav8Yutr7aeJh3RAtFAKxheP0K
UNSpCKszaktFeZIVKXsId30Z+HWrIWPgAUV97kLKm5LodkLGySc54Riyxy1qlcLI
Yz3tFJI8ELUi2T4KoJ6NR0ilu2pbD9xebFxykb966APTbVAICo3uwtXvDPJYP0he
feaVUH77buUH5p1c3zkMe/GpeLjTXXxT5yMEfPdRfN07tE4CvNGk/rV0kT2gXOQD
uE6F/4yByoFLEtxvKTDKq1qpyT60LuhpfgMyA9S3lhDQk2FmvJ2ovIKFcvKnG33j
1u56t4D51BVqthmRVttGm19Ta7Pe46pJPE+1BmQWTYEuKqJB5GLw1/5ocDS/Xxv1
/8IfP/ZX6Hehq0s7wvFPGT+m3IZqG62yloiwoglDhzBQVm6mcKIeEW57qUxJsdmF
XP3nNsnRwQOPZ+W0ZUbVUwz3blTqasxGATqtDcPxiLdf+lWZOtdHDU3TlCv/Ya4b
Ru27LU09ATA9qY8Eqq+quOeMXCwmMKFu95XD7zZqdDUSTGlZ7bbhqAViJDKfcW65
1BCF3BiMlzNGOMWnnEZaIZ7V6FCOufChIwmwvHmRLLBMCUMv+Kv6aOX1iJnjFzvW
iF5UYkCBl0yCeVDRnFV2NnGqMqa02p6fMBKJjJ1nrr9Ex9daIat4f7dd/Pd+dW3a
7Lj++Zrsatihedek23ONcUYW5E3pLzHNsZrQVUxYUUl1tH+Ck3Ru4o52FORHVdKh
FBqK+MMXSfSDnczdOp20XURacSh2Q49fs/9wu6SnmyeUD+w94wE1uprVlCbBiLyO
G1XE2wzg81XNRxAHBXGF6IfNhcpQFrAN5pkby7YUeUhv1m9+bAILWsy4JnvKcc31
A+BvXAzw6z4BW/L9mpQs42miGG9NolAWZiU9rujl7g28RauLiY4NsteXnRNpbhtU
N2oNGYMa2N3ltEAbn0yaxspG+rZXPgjF2cuyJtnA47rMXwurlGHmPuJWWZ1mo7vU
Y+XwEEalwgX+QtxI9TPvwamqtXr7O5IBvnbIbBwjQB1twHjLXflKfFsBlSo0QYV0
4pPTUXLj2For5Ha3EbsudoOVv7fPO25Hkt5/mIn6ci/5kFtgAMPsp5l+AXQ4iQ88
pGtlPbE5shbdy4DxE67ua9SRI4kZPCUB0WhUs6DWq+rz9poqtmla/waRtwqJsFYb
t+5i7jojW/vFmDFn0j2dtUSBYIzLYcu2J61ts9Hv5+KqsswP7+QbbHCK9DmATuMj
9xU43pc2eIlvXDcQW1owGTKL1GFRrQJFEB4cLswyWeffaf1i1re8FABWXn1DYAsd
i5ee2M0UUEZ2T1Ci+q+9ny2JHFovZfPuhNUalBfxr7RqaeWMDwoHtouagornyPIK
YVSA6RP+7wM2jOxGDbrzl5js7uwKiMFWMQeaKt8O6gDFl5mRuBNlrvk25drcznZQ
SIsMO8BfaJQ/F8vTliwvQH0wBwn0Aqao9k1seeO0YhmZJlf4MmF9b5iHIgD74Tua
YKRhN3L1up0//i0VNWEF/7JVr+rRta5n8UnYwdWAiGc8Anj0tXglCQXYYcU3uOjj
wlYykwC17vhxpQAqE+HcbUtU7j7tCOfc15f+FWvDeleeYEx3AdKuiTXUwYkbZppx
0ocmonUSjXwxguUw1/SvfOpKParCn5n3aEeSNB97yXAOImRxm0XwYH7cc30VHSvO
1QAV8NhQmf+x5T4sbZk3l2qtGPhEYxfNwBudEqkcGzNSYGct80IECY4vy+3UgqzZ
sb581IMbNab8QEo3Il7IKfDsKnJEAKfhnExpGQTL74lfOeYqcD7+tWP0hfDCIk+5
QxiAFnMuMW2DLMkRLdaQMwrbZbSLaw5Egec4GkZ8jKOUZ0o4TSG9kPhmPiDuPdzg
yEwQXOwcxQutENfLcTt+/mrm+n5wYBlfMSAC0LHVLhDzN0iZ+87mKfFgoZPK4Ce9
WZ/uUFP7PTDNDMzk6X29vtuVSDnVrYmTibQg1WxBnQd6d8CEBYG6cmdYb9gl2rYX
LCSs1jNRg8u7g+Ih3bZYTimp/IzFcdZtdr9YzjKDWjiBreEHBLrhhHaM2TBg0zUG
tkssaXCFkD55lXJzxBCSkXyB0a+h5Ha3U0iTaJ6nam4guTDpNvw2FxOJlQaCq2Dj
k5y98nEqpC9NE7x21E65yvb1VhLyUOU6XvzDciN4nGhOEy2st08aWQR8T4D4trJq
dcqHPGQFxOSnxJzsc2b0Nbu8BSR8FwIsrR9Tm/lOoGmEzR+O9Of8lgNjlZ6ql+st
LZTfnd0fQmLS7qPk0ItdOqCO0kkVBrksY0iZR1hX0q6GQJENMmwqzlLuxDR9sYAy
dIFi1vdao9qpkQKr5p6CaT9N9G2fRuVeUaP19nHJiLyge1oMYVjBaQmCepLA99IH
wAe70b/EkQOwMnbC4IqoC1gkKf9ZRUuE2+zT1QTIf120dOVhye/8TRp59UHQakMj
VzG6NE5mfC/qWDl5oMj9Z7aMg0TXU3Zt6zIVnp5C84nXfn93b61WWMpXPdgER1+r
A0XljCp+3T1POK0uGVrM7lRbJruMfKwhQqu7wC7JFgG2BALVfBLCBO0D5YQKKlkU
mdiqnBS2KIG/pENUdVzh0sdCmPG5fJrHBxaxs6uzI2u3NmzFpwBjfyPDRNa41wnO
OrSKeDBHi/jbdq2gN4a8F0Q1TW9rG/oI1Pe87bM+Wmjz2LH4kf1pnc5ftohffwg9
8NUV1uErvkSqNqHycR0tgdMLZNFCnzjqvr2VfCNTvMcx/CWNpD727b9s/6fmOnZw
0aNLf7rVUHX2yYwC5Yqb6xnaXEwYPESHpsmAT1oFM++pGEAXk1YnuMvkzYG9wzpZ
8EyTKjW35PLcsjzF6FFvruAmfSs/rFRn67r/2AdzMyPMx+KxCXvxg8u8Ru553iTs
mqtSvaSpLRw0FxeP1PSaWa/T42jH4DnPIYPj33E11tjbJL4L4ccRo+fEXnY6QkxR
+kNXnTCH51x/l6BqlXxVTDDlfh+V6bKUxDaD6lhPn2YgVHGTt4jsjam59njWDDrU
0HW/a3QyJGuhsF9wQNqJSC78lq7t7MZASVRS2d+CGE+ascI0pd4BPOf3BZ0eTjsf
x/rtjhBVhIrQFVjJJa5visnd3gTYfcxo/tOFyHu8LZuBLjka40PPRx2IK2UxFRZA
sAOWuq6Z5r9OBUen3HmprGYWozq2e+nYroYVYvR8bpHuIfHYaQjtlKlpd0v6Y10P
Ge+1GG7lQzFRPp5P2ngCl3gLlq05S5J/O0J74o0m82HZuWcOOQ7sJaC5PzWUD/yP
blE3mM7xT1jRvipt+sv32nGR0nGpUEthDN0put36EZfi27JsjUd9PcAB9kxV8WSk
Gz05Mbhnl6YzrOf8WHOh410QBujwahGzWYTxGaTUhFCqEX8pw149pcDbTNeXhSFi
Bi9D1SLQjQLHXl9hoDZgqAvpwZl9EPL1H4ImSxFmk1myOmNImxUJnRXa0FuTjUwt
ekHxW1RF4+mGhvA/nZ1TcOFWlNl+GF+Bubl4MO1u2xm0ahP2GF/uGFk9welUhIwb
1IxdNaQXspo0FrgSkVHgRFbe4pgAw4WaYqpdBVCKpYv/DpUKdB7oZW3zDRvsGhv/
ss09tq7A1XcHsm8yrjtHuNNLsZdzsxM/eHwXUHXna2g3KizbJ0wSScCj+b6yFMHL
ZmwyTXaRAPIgAKgN/MZFO5v9yh8q3UYy4oOnBlYzI8bw5azBGkEEH/7ehpcLqSmN
teIcFiI/YgxYDpcQj5WdhfFjzJUayK4NSqPboBNU4NW9+s95WNajVvrS/zXNVh5J
4G2vTNBzgYGn9xMkh3KaHljblv/qSI2zhkuNQlYz4DFrJIXiyEajymEwljcDfhbw
A0Kesw4PJ1dANsCMIATEKuHt5JmJG+4re4y40eVbUFxKH6XQZ67nzwGsElhqMMyz
VB1IRUQPeujq2aCkKPFH2Yig6xj6MgLLGpQRzJR2JIWwfdbC35xLC/P6oPmKkmqx
kw9u5Y1PvbO72trm2loZl1dui2oMs4rGwCHD9JEYwcPPAIFsYFzl99Q06zChUezk
xd7NLqiup09KdneMXwCQmgoCD3+mNsoF8PEcoMGrbjN3oTJBeloBGAXKqUeZVpDq
vlwPWUg2Ia6JufC6APTuNhFXQCHF6A8+DcA739MKCyIrm28Erpo7LYwtSxZaap9f
Okp5jh5NwkuSrSQDdO5oH7zg/oF9ZSdWYm2eQmtAsKAsgtVHPEdCtr58+JLMAs5t
YvWbAM6y8Xa9n5HkXJs4r+HDwSr110GDgw8J0P80yW1YRL+0LeYiCP0r1LSu2KvS
0Z74ojQ1Ez6S9sdPc2WPS622YRbwelXZlApt0XwC0XxuaRS8kA9+Co8ETKY1YfFH
UctErA8/jehQ464SGvoPpF5F54gVhfzISrclcoT51AbwcUdxILXY46/R16H90J/1
Dzfa/QoacpWkeRkDnj9Pmct1pd6mqpsyv7vvxMNoWn+7xcm5UWSDE4TsWHOoN53p
YIMHYxrxQFNQvyaofy3mUb5nmKeoZS7+GZz/5ROZFQ6BVb8Nr/QM1Mq02cGelaeT
f3tqZgnMoxQ7xIQNsddwopvdeuRBKT+SMKdOXPEx/MZEhQbPfvB9kpk6PQERNnMD
ZtyQ61NLiibQmhUfjWWIsXA3sXctDQ3LaUNWV2HFrdl43riR569kUV4nMUUy3/Dk
na43mOZoidiGmseaUWC/4G0jDQHX9yArVPZAqdzLREGF1YVmeTKcioe3h0nKcyws
MnPr39jlgaMVf2tg0ObMvSurkAftd3gNymTYYCDxkOi0oDubdEXHYjSCStNPr+lu
Q/n06LEIenG5ni4DEuXvzONprQr8J6by3ftKYfgbkVY0fqOE2SkmQSWXZ0KAghz7
FU7nTG3c4MQ0jGQmjsnQONjtkwtbiCZhj94d7EBwgZ83oXvov2MW+6AhSWq7719s
Mv4FJQPF9Itz+JC2Ne407LzrLUzUGMc1HED81wjZ1R2O85fxoF6872FTqSlfovje
TBhgZe5Jq2poldmIL99lo19iUIaweNuZca8+23xYxm7Fpwf05ybly/JgScozGLw6
S7gZMCZFPszXXKOR+Nq6nceQRbHOy/IuscjLU9+3w56a6MrjCjauNbA4rjbCQsaW
YpLVvitsk8yXS1UbctrCRBYKpvCRKtzouoMgKBcSCs0njgfGbr9/R5zy2viK140S
thS26V2Lzho0GxlsbR3ZUNHiBewUo2Lm2q7q2Lz0xlbZ3XxKIaULFLkzcV9JPox2
iviQSUGeQO0TXMp3KRAG1jtLDhr/5+0yohwQ0me5xt9A3PnBC/62e4BbI5AajjgY
mnupaLfcXsf2uEn5z0ovFpXBtWL/sU6NkAtDBvuz23Law7tqt+CU8f9rnCbWJTvW
AdQ8gBKUzBvsH/open0eyfaA+xDlSC71vs9D4lFr5cC2bWsHHb1Sktp0Y7AGDJsj
9Y5ijufqVfCOlO3N8eZTBQedwKpjo1mx+VIZVYXIsUM19V7gH06BAwNsKiSZXn4B
TV4PMeD9bSDXLpiwAIeOwFSow3myVNTLiEHV1m2ZT4JdR5TEBFbv/sEuM7pPQCRx
Vt9F69I3hdVRQ7zg6fDdIlh/6kK4Q86Jb1dogtSCqaw4se7xeiKQ8aXvgOMkfX5Z
w91FcDtIij3VPrHwEO07QsSudxb7zfyQVGigQZ4ReFOyZEZvkQcnEDXvK3itPaLt
oGtXseTiiR4Y75Oi2aa4DUVd/j+CYUvMGpmGtL+aIPsO6I3CkHuBgEycdW09f3LD
vWhoSMYUeClxY6pNQ7boI37pA6QNEKeLEM6YJHg/vlwA5kCWvOEqtYtFYwmUp/Qd
t6A1WXW+OJgvTCzytdPmksijMqbQyF4vujr4TilQvlLBHCyGa9qplZ2yoylcIIvC
DlYlh2PXgQErw5xJqKjgGH7f+x5XBofAVbpeB0nZzCvktSCr73dqkWcWHLMZuQbu
MARgn96eKljqs4UX5oh32oUZ2bQeEFQrbp/klDVV4eJMPP+/QdgGuByx2tzIZ4Nj
9nhlGJ4C2/n1qSE4Jt5Xr71xjPsw3M/Nj1rtKa7wOrWnO8MGg/BdqkuLTeslcmb3
mRzcYqoK56bk8Kw/4begeMce1vHpnTuRX8fDa8y9jniUl3Rsih1as9bL8bPiTqPr
A+RK13qvtErXucemA5pNWgcd7WGnvJ4ldPTur7U1FvpBoeS100bE4b4C/xmIPxGD
U3qnIL8OmclIvwrsNBGHJlMAXDKsrIO4iv7FWvzl56MYF2ke6zX0UwAncsHu2hFF
YerhyOrToGctXh3Xc0BaQYnZ1vKOSSfV9aU3dzZMcZsfmnvFFVlzsmaUh5qvD9Lx
Cekw50QQ0BZw7ZnAohTRf81bczPhy5VeibYVTlvpzzydsVoKP/5CgDWygmGiD9Vm
6LQ1jf8/9Nc44IDMVMoFZjlJ3q7tzSSEeBSA5jl1onUPCYldk9m1sW5pCkMAB9a5
VuX8RZYSmV/JI6h3Z+c4ZPDZu8a4R83vX1nPj/VSPRr2CtKU3iEtTmomiDnw3TBq
/jfpmDB3JFjcaKGi0rC9bU9ad6Qih5gghbN6mtfBOLebddkC4yofxy+aVbZEzyj/
avlWEEE53pB1w1v3jR2VXYUoVmlI3eKO1Bj2Ftj/sirVXBiWmnHjfcwi4hvFZkNj
3MSpyrXZlOfys0qaUP4HxpNKjg04kToyHkqWZJHWcK85IfdufwzaljG7fTmUDXFR
hkXcqUkALZP9wJ8aHe/X4wYIcPd5GYkpXTuK5nAvoHDrLMcJvlSfijk/XmzSb0DY
JJ+WrxDudmLS9la3pJu/OcXU59o+pZXRICDOS9rUptqdZx1nN2FU+TrVVTSOKbxQ
Zbc0OFYwVkqglgdbNXCkFAbBqQTqv1HR1dpID8ZOFz16yFiccX2NpMxRClEbaPgD
tWpGbfdQAzrNhbgz52mdu6JOf5ZBVm36AM4/8LlbAa5fe8Eh1VAql4AqTpo6LQqB
AmI5/lYBQakCMW/bcD1P+15Rn2oVGcgU+Xpx64c39loOxpEuA4vVsRHRGaNTlD5n
tBPAHR2DGslF/PHSY4hrmNZ9HcpcUngtZ/nLyzdEnBrW9NCvA13iuG0LHeqD6UJF
TI1/U5Gotn3rX7MLGgmSiSDncBPwaQ1PWbK9ARwP4X5C2WvnGRHCJZtPPXiQqcBd
GYv/FlBmHc5tt5TanyRp4m1EKUGNFDG5gz+bk7Myh/fJPK9haRPJkFHvherslZv4
BHq2UWd+lYIfYhmbhdIgfKbaYhlxIeqtt11xRz51eiLdieVM7gSq1eC6Px2wDlJk
Vsxa0ZFm7p3IEnIzqiaQ+3lva88ICH3Foy58m2HC4BWIbrP3wOBggboKDATwBzqg
RmNS84m+MA9JpxSH3rPRjYPq+UIFPL5hLjYgDumVxIEPxUkUCpVBwHSpfWzzoPGZ
wtuQF2HHc0H+Vr/FW1EhTYRvn1GW43pf3SipgAtoXaYGJJ/CBVjb/9dXrNXMjHAA
Ib9WDdVYcoCxN0nHc33dPmlXPREmAd48z0DKUGVTnVaY5La9zgnhQtE8ooaiAxvA
2Y89PytMRGxVb5kq3YBkpiJFchaEThySzlsXAu5LBNZGi8oSo01nAFQ1YZGsQUAX
wBr9IxMXVxzTE5lWmVoUtDgr61Yp5ClnuXYA1tkYVKgEitQheFCFaoOW1xLVN/KT
vT9b1uYTwsa+pVHb3ssIhRAFFCGXk9a+O698JCQUEtOGj/d9I17kXac7kC7NC6lR
uEdUhqgDhkyL9nGHCrkCweK9z6jgisoM02ziTSslShoPbSQMYCo0NbKgKtFyLUxb
ms/MtG5fhp1z8coaZVHTtoFbEsWkbn+V5HNyp8QTZArClfNXxUPXLQ5e/I7Cuxfx
DJdmjqCoCBvRt0kt79Kfi1UD/aLL2NxHagd3geN1me/B/DZSUzVCC7c/vEtJ4Ixf
EivPtGVAktnWIUoqTkf3Sazg7AQf51fnTDufLCIOT+uWIzM/On3Oa/tSQrw4zOp+
Ebbhfpg27mdBabRi8b9wVGc5fbi3dOULR0YmC6+SWgsNhbMXqOqHNOyRvDFVqSgY
gO45qhRQrKAdy9Y29OAXn49Qzg8CvC2FrjIHE8oPW3O7SLcNzs6hSgAVCUN71+X7
4xMxTJxFk74CRc4ad0lx9ouznXiQM0SCo9uviGZlDE9E3CCp32wmjLJJbJT3iJ5n
RADl0ME58frJ+LejWQwMDFYbcvPrRtBTemLX5jn9WSfSY7PdlwJ78nBgUHQFLy/B
RIi5KkqAVjYJ9MFyKEz/WotGpRN8KzR9zCniXWk5nhR3/t3hAUu0ssu5Rfbt5E1E
fZZrl+xg/p+NVbmlyIRqBgTWa9YHFP7oyiczhhSlqnNSA6/u0Q6h2Wth0voX3OKh
LDRXGxb7xd6o2FdztSWWA7rjBML65BDCLTycy6jIwDbZEBzqJX3EFsEXGq24BA6f
E7okTHYLnTCCNPhw8eEOIpRDJy8XSij0M+919ISU4I1Zyj+ylW98gALp/Gzr29pO
OE/yZxcv1i35JssmfKotVXb4f59zgVyew7Ew1GGfXzKKTo8zO1xBzz1KrtPCvDCz
U+aLjegkliCkCfFPTzPhdULY2n0KgjKKnkLOuWckBOT/gFulYjDf8zUegd4NfW0U
yP90NbCpeZ1v1Sf4Buo3LVICfXgSEarDDxpq3emPRuMWXakMRr3A6G8ubGFf2otT
rJRfRN+55zRFJrTTBb4IC/KNBH0SwwBXT8BRDkUAfu38ORg8gYwEMOVjRBNYYHkj
bfWfa50egMrrc+KeXOXcw6n2wz42x+sl2Azbl8vavpUOZa1ZD6bIHDI6Gt+YYLbu
14gNl35xY1gePqQW85Yx32e+z6Q3as8RqEFz1LaenYOyrnljzRiwoRUDiGVb3I+R
Ct7Ne6hWB02kVK85RXm9lk44jdcBaYCiMXzDf3HUQXXJBX4PPSpe61YJUU5FIvB0
ZTh3PVLaQgQJ4AzAYfwmpB6NTb0pbu9GCb0ItbpvdRCsNyRG2saB4DywErb/CkqZ
jUqHw/lLH4NcvR6VdcmGmp0NtOTbk3xk1smlNKRvZni/kIdkXOSQ/l6PHbDHNXq+
iO4E7gzDe8l7Blu4zlvBR2t9/wUgMcD0SBbSjSISTah9m9mHfhh2hNhu//xFCVzu
/8yN0OUbjyXcj2+Jv+pqoCPL3h1QveevUoDXGYBD4+75WkmC/eJQE/+uTwHsWZBK
HGyeSUDNb1hfHJHUMiShC8lPeGey/vT305sBYrBzmjFVzqBCj1k1G66YQNL8txpI
uwGZMsbH9tSQ1UK6IkJCO875ZzvDatzhs+gbaUIL0N241vv3/wMe6Vn0l4dte+43
JMEMxNDCtSK5nxPDGOvVzL89hGq62jsCd8hio/6NXAQfejDrPWqFd3lIS0z+tG0D
kYznRN8om2CZfr1gt7d/bpVALCOH527wbAJns7FBvkyomCNlfttoJC7me6p7G/LL
4QT7u4ml+U/ByTkUI4nlml4Yp5V4ViCKb5UtfrX4F2CsZ3YD/EXLMwrin9zDsWRM
xSmjZvU/6/ByXQYB35GZ6rvGahDp3Rpjjlz3Zc7bzUzNfQXbyJ1sHdP8km2Ub8Sw
Wp+D/JQVirl6QIqgbuT+19PJ+On+TWixnsXP6hkKz+mnDWKK94tyRLNfaTpm5hu8
Gth7fuGo7Sl6ajRam2IgxSGvVaZlwXIqanl9kso5A1Ljkzj335rGdKgExxX4hCn5
Yl5xCi7CMDB6kYYMCYUhUcP6nEf9Kls/47JEdSAt3VdPjV37/nakKjwOgtC2ZReF
Ju2LSMWX55D6gCS9TmBOeX1JwC6lCsfqdjwiaY27skA/cvimJEZM7B+iBWNg/XI7
KX/cAWZKhGrjD2AcOQ4TXGVrNgbmW5uIQgocqM2eA8WWRic3Bj0rFWAriMZ4qKIS
UfZi8JiMRVYkuDYzNLfeSgLxQabo06xrNEVF3VK8c+Fr+UccXjdZTwrYw5L59BMo
SGh9tg+VURcKud5iOpHfZ5gSH5dcVT2FhwoT36MXjGw5qEmTrGslbxI4KZWk9eYb
cNK5AK6wHowSNIcgA8IRzOyILjDxAgTjPJOT7mNuqBY73Ba3RUg2JCz91Ch8Tfkd
c5Pcbw0ohu93xgw/AD+1XGoGcszISUNj/f7E/h2q8k66uGzlamVyKxQUnSjuDDY1
INscj2K7FzdCqa4vAj7/8669iYtMZB4fSjSXVPumWuZN2lOgp6+ecq4GGGC+Krfz
rDf6jlsNWGgCOhWlMgrE/d4GHcqC7qd4Q9JjmhdCIxoYmo5rg/9Jr25foz79+RdS
XnowAcXQCnsGcXGcLfKE+1CyI4NVRCXhJHfB5OCwQxLyJKB4k0OBW3z47eQDbBda
iFgn1XVyrvpRXx2GG18h5FehGDUdCgzngXzChZsaSvuoTc2Rz2GF8/rjwVO9FuZT
0d5YPSU4JAogTmbpDlVvC55f4RVkvbQdn0LqvWLfnx/K2WapGMhFeesQBCvBP+zV
`protect END_PROTECTED
