`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I/tR9qyMYkPuMX4pA70yySjaqvaAAFZPC1ENAyDVk/myxVz9EQ7cA265fSPLdRyZ
MezNOyJMVmIngCnJE5t6DGrqjIPvicvOueenuTpekaWxC3YGgvNMoROUhFZOa2xX
y7d/gfZlAVQlNVyuBWmvh4I/pC8qtqTMvAr0KtJZ76L6UGsVy8yf7h+lrv41sYLg
lum0ptsE4lcy0x12m9IUfF0CLx738lDejCWd7lhenl/6EAjI2unacQOjoVd3amlb
djTXaBpP4MHG/Oxg9UDm4H0Gd+fQlGRCavPhLW3vTCyC6/Y1lMSVC7JWyHdopSqf
m/GXXroOfZ80rojxKOsbrXiZBd8cCVCSAd24P1RJo5AqLFpQrOINtEeeBgFAfWOZ
O49ADjibqe2PoqUdV2exBbJ5VIYJYlab0fyjGvMxIbADDRLrsBtA5Q4IjiE3I8nf
tXwDAbVXshuRA/oPPK6DIUJj57uxnyQUn351E3TyeijONvGApyN96kAkCBpKlOKY
Ok1tJ1izBsFX4r25IqbIRlwfqoMbPBEGFkttnd4qF4VSDsYWTnBWxovS6LtITN4x
ZBi9vpBmMTrMgyHnTwLUztB8uJyY3+Ym0Y63tE00TCsoMlGWv8MvlJF6YMisvoN5
/hdVuk9QjXvqriqRh/ArVUjSjEWEYuHVEddm4fwxotcShODC8ElZ/CGaK1CdHXow
aoNrTe3SmC6/rDlHkJABH69lhQMWW00Fgn8qEKAWgbV3G/gFn86yZgK3+AzGSXFx
7OwHEHYrcHpcUcLRf4/FkJLwbl43VvheB3itY8l+kel/O0jD/E7UdvrhQFjf7VXc
bvbRaZ9jy7pDxhJF+LSvgboiMjdX74FaCR1MUnJKai6WXWl9HwRr2W8gBWWFm6SJ
tcY+c1GGf5PYLodu7gyqafFXMJyphQXL6E9iPdLlFGQ5f85raEX2d+7zdK1sQfNp
qlh0QStcbLRniVL+FQ85w+zti1fEjWnL+7+lLTyxNOk+KP9Wa1eJOl4o5Usxg5vE
qBGrX6wzLO867h9WXSVdiZ/gA5wtNKAxWhRYnf3u4nGE2p+0/GjJuWCJhmUdfo0A
VH4U9Jg92IhsB7w0ho7OD9JxB4qSHy5i8clrKNqJryzJX+xNhHHX6Q7EQedf8K76
7Zx8x6aISwsVnF5sgx1VEqw+T3rQYPguJ+tcPexpYZNEFfMMuh0Bc3KY33jFDtHI
epP1NKYqdH7NN4pe4Tc+PRtpQpZjm3vgvHycswvKo60+T7ulHSE2KdZCr/n/8kFY
sn4s8wKqzP3gxm3vgaAWZJePXOtmabr0kYARt1JLlMLs063MnuUjOsAVSUMhCcvS
KUKD8u0kMwxl1hxGRLoGKv7snRN6Blmb39KLbyQr8kbxmAsnWb8AWKt7zi4sDeW8
OziOdGNgEg8DRxzUJS09sHTk9EzeBPecvFoPzvjPE88Xj4VgPjLe7/KrnpMYrk8h
ZzaHeLnnvBEWWS7BGyYTI1F/IK3QT7ku4R16N314mYe1foGISUC2CAPvBVZgU+uE
3E9ZqHpcUbtfta5Pal5iq+RnDC0EkBIVj0KZTpGNbXJJ0cewz+uQ3gyf6DKLZ0Fo
Y5rcD0ksfFvjU2KAzGbkgjdan3aBmzhl3JA2RyLobELQKJONPgDR8smATmXxdAYc
OyvcKWVV7OrZc9+Mv1StZoLpMAszcuIUHjF7FUuUSk6BEeP2Zmywyw6I4Mquntnp
TTjHhKoYf+eSKO9hzFg+d625s7ENOpOUqFyp//MLUE+Gli6818ZXZRMKgFMa+Ncv
SnL1xCt+RJBYWz1rnRWm1OJf5EuFrD5FVDHWLPP0sLcvhjzyAxzAf1ZmQBXN9LR1
3ovXOVE0JmBNcgmUpGNygXIZkFZbfu2ZYjuJoaPf3cBwloy9Sa9gdWdCU57I32uz
/WG6T7/dKoaYb4AHz2QcDE54xxSTZecewmeQ286X4fF5AfENmpqXfT3yKsDd58WS
JD9upki9u3d5sMInRPWKRtifmSrWfE5/5Hev2c4hcHWe5OaRkelqMT8BJ5GcDkF1
sGSoVVBDwZ1pBbadRClGNaCYg7BNmdZ2u5F+0jeu/Bn3rEOk5kC8ij+QUCWR5zWD
S9WwDmkTaX+rqvzlm4Eo518F+BLAZWjnRRFZKJqOGM4jDpS5+g0RUEUQABG44dpZ
K9aC1hacI6TE22WmDsZnNOR/9/n4uiT/AWz87181vxYhpI004zLIhDKfMBMsS2Xr
DqCm6KwiMJce3fNtKe+gJvT8LC6ota8Ibsq0Q0MKdopai8nBgb8Z9CSxuPdgVF2K
zWj6qENk2TSzgDt6Kze4EGSrrN4dsmjJd7Ix753jnZ4WrpSd6UBEnmn2hBuxsLhy
H9B4C64hayncSPOtldW46se7LxlJRkil0r7mmhctAQBKV2zI61x/r7bweQ4fToNB
pKtTykrrkI3vLK2JWXTyyhavMCweEIezUE2WmO+/aNF0KjxNqdl3a858tlMlbnAj
SwtylErenSjb9EEybMbG9eBgKLftDOmcwb3GRs3w7Gn7TVNPt7L+sL2njK+PXzmc
SUVvOI2//Mjn3WJ0wGz5bnXVisbWJdDdWPonzyHlERIsJhl9UXaMuj2FUU+bi6WY
zGLfadzeZkDBkHj51MI8ACJk3PBMLhs++mevbpo5jcnTHJrttRYgGu7fsVwcCwDO
VLrpKsmmsE27KHnUuSXrJiZ3hrQPDl8Arki+3iYWAUnRpGCuXzSI9UI/hxvyGWL6
enYcCNhmhIGmYTTTA4H0/quHdTkIEdvh0JUY8zY4vFWdrJ745Pt6sVTmlNhxVxCy
wTqM6X4HZPBMYq1RPJwmuKUIJFGsHwOYb/f3FWGcVhghydZxWsehAHghvKsVK/LJ
kO5zHMA0VecLz9KrB9+/CBeDgt9lrITRsSM03y6ErSW7f1ivshGNdRZgXjS3Ji3v
3UqWuQ9IXtBtdl8OVPyKFZKW51WDtFXrsEDcxbzBTPSkEy1wfULRqUNd/IXbqDan
hbcMzMFd4EXwJ4Hjlf+Ta6nHAVCfQs55N4OI4fTDu6i6VgZs533JUSK7lBb8uBm9
hwqMvtkXO0rmReBQ2FCzMrHxQwwqwpnlCT/QGyodHjhfXzl2IaumdvoxI9m/BlqR
3koqouxyRFv/TouTjNrI70xu5aKfUhJs3lUMrZeZawkZXHna8VsMNC6lCmy4CDF5
4rlKGryO8Lz1FtX3at7zdNnm71/JMo1sXj/I1hy/kcKdkC8INIKPU4GRqd/PTq+D
gayRDoaECs1NtDUiE6mIhlm9aP0H6FI7caHzxMWhNtHOamLeHPY/JzJaXLdEPx2k
RzEVPEqpJK988wVj6dK3d8AhXL21o6vboFLoV+uTdYvbhEbS9KT3ijUiUWVviq3b
p0GjTihN5fp3EiWx2nl8cji6VxmDRYzxYSycEp2Fb8t0mcn1QUu+hGneKcBkVnf+
RJIUov4rUDOjrq1IRMRP/axo9m+GiEOHp2aKDt1Y7uk=
`protect END_PROTECTED
