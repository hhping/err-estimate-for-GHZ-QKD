`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TtsIoki/jf2M5s4Aw390WrRly7JCi2RHc5IzVBp7MhZmv0g1Jk55HYzWTjHn1Gxg
32gc+BV1ih2tArNK2SfyEkV+UHoTlL6shVV/sv7qBtqqcukuOFUQlJP827wD8xb/
0ET10I/e+d3yuaZIQSz1X6u+8PDgbyTSJN8VzycJZfA/nd1lvbK8B/s+R1pbS/67
kC3f05g9jT4fmyu18BSX8uBKQSlQZL+P7NVPagg5rzP7bSDZefhWrIe5zJCB+kTa
z/gIi/sp+kE4bwMJ2xVCGEaZtatxhgQl2CjN2+fhnO6l7+15bQQhHVRTmEQfE8JO
sRPqE4odHL62yqu4dU582BktN9BSTiJFLradFojX2hShqnNe3QcZUK4jqx9Dt9/g
XXxmHJC/yA44BuiP0qU6MCHPt2NuYH84m/Gh+5rDmE+4eKcrh+40iclDTSUOWfi8
tWbixMXCdO4w8JXBpsk50F/6FXjj256ZPYl2ZkjpQykB/EAK5mZ2hQMODJtnFQcY
CrtgoMesJP0uKwkRR1GkbL+IvXeXP0aobnQqUQu0iqO6d18F9GY5jW1CEhqjpu8k
qWIxP6I/Eqj+NMKoCDg9QOix9ugbzMy3GhI0CYM/KnSFP1HCVFByiqyO8CIjDdiY
oDekqYy9/nCT2vTn9rg1Qe6FnM2IS8q6Vo1TJyx8jpTDo7J/6Op8yrPEk0lfSHzL
HsaHEG63OLQcCTgAp3ZHvH3Nuj14mLj6F2S67FsBtVSDu3yXZbS/FrFLKb12N/i1
PnnJc5/SvNk/j9cw10F9eGbyur0EZixLun3ekxH+h6t8nf38rOOZECIy8pS0WDg0
KL73pf/tqCASe9BDn8ZKU4KPcq78AMBe4W2dfo0tonKEZ5p2Dxyx/6rZeGGPZUDM
C4vrYsSosyfKyInoSY+DKA==
`protect END_PROTECTED
