`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6nZZpZiDZkFBE1nYa31DFZ/y746FqzQMw5qFZvQ7s911jnb8OEMhedFu/xCiTcrd
4s1C1+hjTia94TQD7SlFY/OwoAXrakeAldwfM8vt9x7qppZwD6D8H8oYX2GvJvli
LrOq6TsgI8NDNVuMDGjAyJIRht3jRkp9ZWYJdaWi3Aj297cNfg91ixEpfp5Ir3AJ
OSdJe4TZTR9Fcph8ZDm1UiFySF7UDi1i+IO0rv/AsqMcR6d3yUz+Bauh4JrEOOfr
Thcg+hcYLLdP3HrXu1yt+ceN3VbSGk8OyLHNW/xn9Yk6lVoAdnqmkqWDOaur/s5Y
n8R5/3WtBtOS9FUPMgH5f9jLdE2bwN49Mqwf8g8kNbXg9WsFHGZOoWIMh+RwT04R
k/qqMYiLvSoCV12MAZLZIFyiS9+/mbv1xfAnOKNQGjh2vMeNuybG1X6y7E7di85i
Iyl6UVfLdmqJaYWvulpPX/CGVaanxDMTZY90+OxuISkJIi2iWmJVN8+qBAHYU6Ik
BHxhKjXtNO5600qCmavbx7GW59wGA7qIMXwrAesHeeqagzAzaUIBmWrvBXfRgv1k
dyBDpCDr/wWS9wLmZVdVfC9L2VP+pxb97OCYPjLFi70dmCj8euiEXUFYgCY0jDEU
J+e04lAAxfrO+A6HnZf76UVYdMCiXlgfd4q/ySGjLhinWI7XzrnblyhNAeWZRGbk
CwCq7nYIWhjrXH9IDjw7yD/UfpLvq8KPB7KgeSmsJn4m6Y1rmWpMRkzmlZNv8CNK
UazbTITpGElGzRcYT5zTFc9d+oJIge3dU4OEgR+q8GLDrRVn0yFc+5VXssKt1Nh4
8NZDrez8TomwsSKxNhb9HCcbZfuB25A/I//D94o1894IF9UH4Z7Lbsf7BkjAn+mO
OHRyE/hbPkEYC6ytl/IxX+zZHCCp6mDLpla2INP+WPwRcLABAZexygKrx+YzZUeW
TwGkRV70qjndjRQSczqvUrVRRiEj7tgf9V9NmSXWLFCvuflElhZR2twqrRiqHbrM
ZT6t9GiBoOMhNImslSzgaVgRuBDVgsVuuEZ8YBlX99zPo5/TZsntVcmtU5T+dfFp
CxPmYaBOKbkU5CB5gZNd0pD8xDOpwewjA0FMWFI5kKoXzHpgKOVanMkwPp/Z97WW
7ZZfVAUw+iq5gZdc3Hg4JAQeMHmk+t4jzFLoMWt76lgCGaYbNCDayMK7gDlpsgfH
J9iF1rkm8aF+okFnkd7YP8HO7I6Zq8JmhXbb5iogTH7NTuViD+9Wpoh+O/OY3MzU
p3YswT5V/weBCLXz7EsBwlMeCX+dFhEtyfjlaskakHPxjg9zs4kfd6gvdmVX6gzT
l0eqhwMQGCNJmZq2QwQ9OmkcYSEVZOU8dk9/GAKi38IASR1NEwMqMmxlpOB87M89
svt5HpEu7CmH7decW/lFFR9w6UswSe2Wt0nmn3I3uYpEP/zCXmW6Is4XR+CN0DI1
DvaBXySCAx1feb1DDT/wHVY2kzIv3/IeCyZjCOHDzFiXU6qTck2Uj6tL0gPMwgMz
Bmwfl/4094BhtuKY9j0uh3/QtdyANS+IF+cmjymlvUyGVhsIQbib+Xr5ExkNBXhv
UeO23VaWlDlWs7BVtGhsZBFqlglF/DeX8gCls6bJrOPUtcbIZRO8I9j/Jd0oQGFB
xJE8RdmWjFCLC5VjfU0NvAO5krrYcjZSVkNCgFb0aBIFhJIS2uGZY6vOn6oYbhs0
AkppupD/mUxD5KgAWWNaQqgYyIkIPWUvcGi8LUHn2bItqB4wjcQGfJa3yA7zWBMM
/uf+RLGnGoK7VHd/0lpbj7e6dXwiuqh5ga8x5E6IfgwBy2AipXxBxbHc83Nq4jOM
hHTgLhNoJYL6gd9sSF67ilOsXwTiL5akc9XSqG/l0dSCQ9bXV97Qz42ddpEO5TrD
pIMZ44WCpfKsDT6JhHbWzTjtoQX5O14C5w4l2SgPmb73wHcZuzQRM624CMVsLcvW
zKyMGLZDyMgTCx36ltj81lQkpWGpHd/uzPMUy66Xl0dzp6XxmNihfKxCd1iUxqVA
JI+peennn7MBcDIH8I3eGJe5q2j6pP1Me6jiueykG4cxBpWgTcCu6VIvEgdBa1BY
ncggJ5GPJb+/mmdbKLjOQfTI+T2I4YV979ttbtFLaiN2h9nBwNlD8CM7Sr4tQogO
4cUIP2r+4q6ayjdh2964hyALS0Au5ZB/5pkmAvBx4/b4LFDnNSHi1hJ75tAvug6Z
LjZZnmohDoqF/mooz3HVAqWgZweglb4awEEgoM7urSaooD7bi2iAfXJrdREZ/iw4
UVq7KV3Fz0kUHbwUOvQYgD8/nKrb9KmXpIBhKECco5HiqJ6lEYZJmkaZd+u2TA9O
PLhkQvSeTaRPX58Lz+RzE+SMgIj6t/x2Z6VkBuNPdNYBezeNuQCJh9u7CBTIrahS
jHa7deE6+thV135T6+a6EWcQ23IJvzOUtMdWOzMFghc6ERiYwrsmdmd3Uu6IQh9/
KSQwGKiusPWcEeb8eIgg1+TY/m3Xywv4jebtpgQtgu0pv/TNxO6q1/pHdIFzGbXy
apSnDbZ6h9yVK2BOPGqFFmhHLuPQKWeKPC7VGBq0uZXMY5RLnvwI/Lk6IbW0GNS9
G6tE8I6TQc4z/llt86M05351yQWafE7x8Qu/k/Fmz8SVwpcX9MoVkxgz6DsDzoag
N08kJ5TT1lhjz458eDy8y4utr6p1RTpZl659DIXfxrI6j7EMCxAks6RCGsebeV89
4HsY/nMFwB5WG8YHMZ2VW/5rf7qlJbd1neU/LZHxkyQgFj/5xDpfj+uweokLVgSo
mUBO1RwhE7goBFmKp0rqih8xfxia/t7Wi+NTbWt5jZlYvL8ZAbh7T33wcJOFNANi
JIwMBogt3mQd8HMZ1lBpvdA1nGKKUc7qNoYJBBmRLzAlhzyhHmlPciLZeDhYZ/Q5
yU0gmUbLOjWNk0T1bk4TOm/L0vH0AJ6UIQjEVTvf025XwEVfcMIIpQdwTBz7qDOu
Mvf3Jx2fg0fcqil7N53fJI+YpYqxMC1wPyBo1MxRrqwP0bRDy86rtBn5gXdqUV0a
xmcxmcmCe3qwo3i44jE0G7SgZbzE2/bgU6zYn62VsVkGdOeZUMHBbXgsQgGA6L+s
elpw1kMba5b1t7I3cQ7VH3OIIdlIoBi0qxaICIZlci2Syv2ZvnBRmOH+/2t5mR19
U24asjUBRuFnLP5OZ5wc7Sp7djwltfvq+e/u+OlEKyxQdspdpulxUJlibAKsd+r6
eADyqc9fWGYrAJlssoy3D7GgGrBh9om6UmEgYHtf1UOO9LxBy5LC4eb42vSAUF8I
nl4aBgdz3LKw7TRu8wmFcruo/ypZ0ihNY73DqlT0UHMwG3ypL7YbNA4Zh3iNL06C
9vS4NfrXGpRiYoggatqSyref0fbMdwhqdtcAjSioQ8YjU+8PTLyYmJzpdU3ncOdj
Q9KsgZcEaNAwge0tD3j93V7tPP5FuNEsHwjoAYxMVxqXTevFj+V3YUtw+E+X8KFt
2QtlymsaXjYlUbvYVbCKwJBHNtdE/6LYPPYDtUiQ75R97BEZN2L+HDl6GtONa1/g
D20dZ8yyi+dxc+ohU+8lb1NVhLj2rfU7lyaWVR8q4r25Z5eqNn36vhPF5I5jqPK9
kbvEtslhy31yjupNLhcm9xq8OyM0R5gqtPsmflhasu0wbA2NoB0z7+MwS47op0ZH
NrRwXW/PKzpY87Q9mpzdBTJV5ch1gGtXFJ/IBZMHP0h8VmVpMf/PXyIRfGDHeyj2
rgr78S9m42wTk3D6U0BQbAaVWGXpRVQ9C5eEKFIr/U/kuCcaJwfrS3lWN4MeNpIm
MXBvezi+0FueFt+9sFo/wDdVFIUWrE1OVzdrlf0A1J+h5LDfgtD+IsgEfJN4oivv
dnr6515xVQ3JfH1QT/aeTvpxJ6NJz/EddFCP6DkLGs7F+IbERCWKulsMhpbD1jqq
GyiC52mlGhrYqEiftGTx0Fb/4NWYGmSQQdZO+DYDFFPxYQSpAnWLeC9zLwLzYcuT
3eg6oHW7F6ebO/dHvpKLqzhmTTb4hO3iuXyCP/EnouKvLaBxIEcIaG4CB9J9K4tP
pYJ8Mue0zldj8wn3C+cZqCvVu75+h64KW0mD376CYjrtdqEq1mPiXXfb/RoM3NYg
GRTZQJENqDm5idU5AG8v2C3gcp97AYyAbxtgincZ8/qD/nxATKJm3aOcim9I8+BJ
hpS28XGRFG2cySTZDliQoyMgyDFVUBWzj4rWIZTu40V3aIUFKFTsAEB6bVPHDi2o
d4VX6A+dm4KThauxJzIcjTIzirlLQIjeDKWIi4cClObjcMN6GsBZO26Z3F6uiQ41
6gwd7d0qGS/QaTRbx//fAhQoxQ9mHsYmfQLSrLch8lgFa+gcKnZmZcZA1i899RuT
8cWPYRHY3eOpAl9uL6RW9NfX1ikGTh/ch9y/1lN2v2hqKlRc3zgSSvxPH+cDse91
beA/zqn6eccoeC3iEHYSlNMTq6j2S7Adun5VdOPh7xdITee05UFn6pEDhNSOXP68
CZqr2McQPH6pIFpOUDC3VKSScLYm7P5GYEWivsRfGM70jfthEQFOQlE/IQlbajAu
f3AlxsRlheFJFTT8KL0I8KgjzcOGCCAtjk0WfZadPr6zFx6IE7pYu5NLJHZQwr2T
6218YPhT9+DqGbbTnXmzqkaOiVyr7oea1P/nLpDc6ongm+aH0h7TkqDnQbArA8Fn
OBT+5rlrREGz+flIYDm5eAb+tNkzpEWW+cfP60XNu0iDsVKjgi7m3G/KRRXwZ0hG
r6epqkITOPotTsiDRgfg3gPE2d8W8Qh5VwSF0ZEXCOasWKwAQov9+zGmpaCC3gt0
NkmqNMAjcFFEH56E3bHfrcGu1t+JmBGfaZF391NWIxAWxZqfg3vnMjglUdzVBZK2
ggL0nYwlavGIdilH65ylF87Wh/RTuNsI6nvD/4KpgUjJP4PePpt3IdNXfMHmVADP
xyOPpq9bLmm+d+yVofWJiBvdE9rgjFGapHw6eZYtb/0htlKEVz7g2czW7Mst55ZJ
oS0BscZFc88qiu/p9x9tyf8uSufKm1/F05iM1o9qUElt6NQ9ScykR+4tW620pX1q
ApjA2ciIV4DmR7/lBX4MbldzTDM1fZ2udIWFfGmy6FxR5ymdR5lDUP6h6Y1bvvdF
M8H2J6yFAJKcVPLGXjCAXZSYWIokR/9MQyjSXteD+t9Pjrnx38hTNVLuuS7JDK2H
0Okp1QLYeT1yHOE7nNmsaem2ZV/1Pfy8/uUfwhh8TnXwjXBtZQZW7O23f0eGA5ZP
4hBW13tG/3W2RQ++BWqsiJbwv36VDo4xsfB5bvJtXhdSasaoIMisBUDFXilwu9z0
pdwCqd9vnsSxI654JwPTa8m5yykrpRLObIiAEwrDVMzAq5Indnpg9Ao6txTPX9S+
HvQyBzJRxrtcT/HiP2EgDYwaLB/3rq5KysxXQsrDz4ra2TJ0OJdcoHun3eveGDhZ
g+NtkQfky/SP460p2xWyx3DpdUZzprfEEa/52WpOEfJ6Cx53N9nxUYk5whgVmYvB
1IE45ifZXByimtgX+a+SJYaoYFFUjExDUtZYBi7n/JMXU0emBFvf3cuCbC4s/EvG
6f4ME1AW7AXCgdPV7u7tskWza8Oc+RJEbVd12zvxTV5T1J8uq/jP3ZA/wFMPEVel
YqytQ4GuPxsl8d+xSeWnqtxLqKCTwc7TGa5oqvEg1dT8EpFeYOzx4pDcBnoe5/L3
QrfEjDKbPN7hZC0DLGa/7mU9lWa4XRM5qwZJMwpX+YdoD9HdUs3O4KYbVZkTlAzT
C2w+OT2EESGsSbDt/mVRihqECFloK7EdtdK4+WpBfPCsMyYCOf72F1H7qC+TuwDl
mShfBORWbfDlysuPY+T38n5jQkSipRYRRWeNI8yUJszsG9x6JoOKca9YqTHIQrGO
2G9OLDGEY7BJQ3N8R+uyyaBhwmB6Yh86O4Ki4ucvgfWFV6V0JHeiuuFSRLABNyJi
/ibFZe1kEDs5/79gdc27NwJ17TAocs2MJkovKZYznretmTTNVU4HMA3PEA24xf67
ngrjSiusYeJn1850/at9knpPvH+cHYrFtT+oqgzLOwmw7RDNSqQ4lycNoByxR8eY
QbRNMKPPLp0GLfWaj/QLdD9S+Z1no7SfwDxSbrIwmMgat9ZXBDlQd4M7oJXUyplu
UhLnfiFvVIcanHwDfWL2SnrSJwFof0fktsBf8H1XYJ2bgasl7MiAnY5s/vussHMD
Zq71H+xSKYYSZ/Vbqm6dMTy/vLGrxizOA4NReE6pEJw/rCT+97cs4LatESvloQN1
MLXj6eyLQz3402vfXs2OBveAbRK6xdLZANm7SUuhASvzGdGY/s02pvfybZoyKx7e
Y1AczSmxiAalkmyR0GHFJXLcZTK97HVbxfZceE2olTYPqRRjaHJTr0q9yXDx3cSM
+T7VtsR62BI4H2fZwjWMCOJ/cDG0rDOA+S65DMkvWdYk2yXTHwUTWx4DHKkBML63
WJaSorIu+20WfPVs+O9IzH2lY7X3+aHYe2qM15VPE9ipwyLIRY/wG1warZ3FKjxq
VLKl7cM2Vg5joD1qASiWxSkaA9yBGph6yR8V9+2WRNvX9+Qdtn88FKPidkW3o9lL
QR/JRX346hSxMgWaVpLUcazv6RJaST1IxWwr2EGxxxjnIu+j/VGHAdDtEAuSKO0f
SlovjqWO6xjJG5VUU+8cLWXDdLb1Hv4MJgFamtW5NAklFQfcAAgMMcm7lbQO7cBh
JEXiVrNx/v9eeqgJ17oE1C5SYgpfc/xwedaLLn5h3oTBhZTj85GDemxr1HHioJZa
zoCx+mTO8Zoy+0G3+tNNotLbiqVmw42HHLf26IZLoHZV7yakMLXA1f+Xk1I9wseT
g4qM8Qa8991ct4dyw9WUupfIT4s7aEIJmkkKaVDp6B1j+nXM4gj7cw9p7J5y+bIA
WPFymcJWteX2P1LGt13BQgqLMjkej+fo0nlJAmFqfAghhoxPKZiVhu7Ke74HvpAt
J2F5A3YOn1NFCLNX2Cx1E675NjH0Sky9NPdxNJl5GLPsUZhV198cRANTaC7vFK3E
q16jH6Y/JM7ePhj4I7d/VPmwlhoEsV4b3KeelQ8kdTZNF4XLUrbq8O47fe5THAFi
IxnBrrSNNJcDHFS758GvFx2NZRqYqk4PFFeF4J0ENupNWK2t9MVvxuuEPkE0tQTS
bifEAn0rQWW289WyF9mRRWJmHHkNbSq+SHXBmXqMzf4dWvkSmNtUs7Vht2nJ1VeM
QcurczJdu2M7Cr9JO0tJe4smVqc9337hTlzmUZx6wOIDW9zL3CwkFg+YnimM1Fis
lV5QalfyDmlYJIx4xK0FqD1Vr2o2xeDP8s2TsMTnZqRCqRLQ4xEo5Nsa3TOAEkDq
p/X/o3gcFbgA2aD7AsGgQQmAXqxg7PhCwCutHMh2L001w6ECpB+s8OP7zhSe4qsQ
hpNTYr9KAleIc6+f7Jgh1giG/OQzVE9bbVF13hVk3HamnRfy3lmQMDyAvWhBR2xg
uAqSw/9MupqUisrtLhFiRL9xRJi+1c42zjMvTm+WfrI5eGHL7bFnfgjfsmB/ZP1T
advCSGjfAtP9aCRWuuJaWAIh6MhUFxTkUqYIPMgU+dIRnwTpnL0sIL4xYIU9ePJc
AJOOjTUb9afAO4rHXGSAPArpbiNVLE4vRKbPi4LKG6j+VYzbFdXehhWVIz3V6ZhD
YFQKYxTeUAKZKG6mH+M3h79DvysHfECvusE1+dyw6JhR+8/f71xWhhC92igRiESD
lfXydpQd4q8tWJPnhjgYzL0YSKflhSg93hQyuhzICllTwEFPkiqTBq+ZpmZiQ978
8q6/HVk9SkotyrefBl4G1v+THmldTHDQEssUkkahyyexkihcOqwPvt2vKs10yKYZ
O0j0pNreTfk4d4qvpD1177d0VphIqMXeRtSw0AdzyG1tViISmd+0aDQUH8FFX6gY
8Y6Hd+0cHGitakZ0vTp5CG3McA+9zShoOYOfILeclyKEyPgIqS5tEHlUIFmsR8Ad
FuPCHY3b4w/EdnPxaIN3WJHejImoM/pdKpBrBx4/eSJG1o84kk7D2QolIMeyZY7v
Vkk5pXkKy6hA6Ukym48hdQOqi28VNKowW17CD3VUKaAwOrUxUqC6DVcxQg/4+Sy1
p6DrvIhSXgTP3Z8yWVWT86BfPma2MLnhtWYIUr05lcFY6xMm54NMw1SWsFcP+RSR
AyAtSejYYfMdVO4HFN6vKjDyn5RkLnGKpkst98E4mBjFfVgvPDGoSA2jg5oFnIYs
b90y1KjLtLNqeiyvlN9AR82u/O1GpWsv+MKj2bIBVo5j2YP99Zn6BGl6rxYzIV2r
xPUQiYgJXHfjllKqs8eRR9Zla8s/Ai6j0OJ14HAqvgYZ94SUggH/kqvA2UPlTrMy
GMYe8l2tPXyhcnFPq1+UprCqLNjRDWsk7ow+XjKCpeUMTm/TZxiFyspMvomWIRXU
3hCtRtFwzQZ1wo96U526fTO1lIOujw9i9VjHtHuIILmHerZoAuPM3FnNvp3K/lHr
6egkROPnJdcRkaGngXu3e88OFX7wlDucw0STbpg68AXWcc7Eyk0PX74o3CkxT0wC
QczK8nLAE7AURzNhe1wHv5ZX1ZNj4GTN1A24Njbm/viX+01kfr6HlUsXraLxpa8f
+IDIGdDZdredTexe6/3LM6vIFWzkcjxXYf3p7W6nMXl3+GC7FmwenG46Dy40sBTz
XtZMFrNopciMJD4u9wXdBKnKUqox1Hy8WomWIy1VHSkJ7vecQq62jJTBOZB4zxdf
msy5XHnxRHSeW/xdr/meDn5LDvgh7UJQ+rzO57qU0lCk9mRAb8QeyDmkWNWdAxm4
51uHAEFnDJDQa3lzFVAJ0zkMuhAV7MguBDm61B/xEsyxQ052cH1Nv89sLycjZ7WU
Z2cIfs0WYXT1wpmATWy7s8sq1iSiKuf7S5w386cJRQiGI+OdpspX6Upf5Y0S2OOW
8s0ivwNMsCC8kLivcUp3CTiB8lORbuVAy60A2HIloKldybcu657m5vnCFbPFoaNN
2pY9sjCmpZL/YhGWI/uMty9WT94TKoGxw5bL5IH/3H7TgjDuOzmA6ivYO5QLWbAz
w/zTqLlH4gr+t2Iv3J3Rd1IXSIvSBnl6zLgZ9deoKSBDR6F2ASoP+NAwJfXLrGkp
PqU93qsQ2m6Y/vTDi/FI7rwIi3kCeZI7yajwnkAMJOC6PODlXuGBhf7sdF2kvzyn
dd+5ODz4oXKEFZCsSFQ3fkR1LixFeIkIMHHBdY6A8rCOPHX7y6gA+LL+1MElsXtG
pQNiQuS52Lel8FTZ2Ol8XuIlMmFECWyG9VZAQ8I9PILg/hOTk0/a7NvI9qY2vzpu
KV0CUXSCCo908WYZZWqNxUNCpaE5OhAJt5tReii9eS9OPJ92rJMWatYo+l3LKMNf
ntuwhBWno3OPitSg6DmI7P99YzWj0+UcGmLG8LwjDEzkE1gk6TNdVovgj4G9jYYd
TyOqyQkygaWSlAcmKwVx9PZugaFHSW+3PuL1Gxm92UlusvpYFG2zg/bHqtzE4WVc
oIjf/ovKUAb3duknxaZM+dHQwzIBimhHE7Ry3VQ6Rmq/QQKjg6FNMPtFgpXBonNS
yZfC+cWarGntho11U0JvzeZuoqKs6VqOBLn825R9o9Wx1tBqHPN+MT424L0JT8Fg
BKeW5pf+iPQBAQj8Q5ZUvxPP+/d+Fe0o3B5GKcRo4uw=
`protect END_PROTECTED
