`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bo9zaPvbWCFSsIpeuzTdRZ4Yvvpo6aPyT8V6Wb8a+8vFCGY0BnQsQjQ/gPQOekkk
JF0PcxRantmmgLxusKuni/z0dIAf0vkOHExsifmvhfOJPz4okorF29w3x9dtn0Ev
+jEWGizy4btfXL/Y/DeC0ta7Sd0GwVqgJCMBHiDozHhGRiGIwqX8FTfq63AlxPTt
K319DtS3C0f79Dp2GoAjT8ifYmccLmEPotq/oOYqX+xnIvX2OYpIjMK3/AHilgm2
dk+tbBf3++TSYMiY2BDVrIjHfMAaGHUb4NtALn8c7ETpOYXsq74ltpP9LQb5/8dG
IXs4rIWN0nKKQT5mdmPLazQVA4nj2AFRiKD4N7Ygds5gsfXvePnIWCmQrcfYdSEp
Jr3ENnNK9QnqCeZlxikFf63BItZEz15vqGyjIk6vV1ACVQWC28EaweXL0ESZd/q/
0Cryiefm/DgfftePeCE+iTVsY0xCPexu0z6LZL2fN+BoUYn+L44OoZVt4uzLOuen
4MxK4hVKXsF9IgYZtD0cqhCknBAmMuECVxFcMYpUD18Hw/Ite0YzTU3pra9LPQzv
kdEHrDvZoPnGYKRUBKJpmwryBFItdAUT1tE7YX89ozDkrNXEpTKCTfh5dAcvx3GI
grxfFO5dy5lWjHH1kGF199Q9D4Ba4PAHb7nIiaKzrjlyfEyibLRXbrgJIuw0o9RY
bqHQe7w7xOAZcaTod4xBTR5SeDsd17HwkNvEZOYpVgY8jSVzfv8sn5ASTjrTmkjd
33tR//vKMJj0C56CxvDiTSIUjnR7DP0wp3b3+K3712o7LnFshRBPcaaRCTe+XCJm
FkreueftyiQ+rNXdnc1Ws1Hh4KC6GcEDJG6oYrNJerksgJSEobIXmqap82VGfjgE
vtT/YpXDVUeLwo3qLFYbyYtb5xRezT7rnEsZVvGC4o000T9JUVsrthscmHneYVbK
xfrV34X1yJ/1DguBBDztuJlhNU6eccqudogr9rqDenvGg7PUy8FZhIamuwQuKUwK
b+667vxiTANpBYsbVuHchBWsOU2GUFGAsKGbWgw7iaUKeZ2bvMqOIbhqzlCELJXg
BPjYLioV+qQ9C5qsiom5fwkk1AQFj5eIv4XIpPlqld03VSo2CNW3wTushbSROPf+
AdNZ48Sc1FZZb8607si6px/ovz1b4l5UHDqiQGWdfL4enMNCV8CHaW8tYQZoOSNr
BDcb4qDd2Gx/imgOQ9NaoTWEkBfdsXuxyPwMMl+FE/JzOj4xly9GQIR9g2C2ICvA
+3u1IYKgN6N9c9cIR0GihdK5nc8f9Imo2aa+pOUrrulQtV+Lzhao+ZGhba52OFfU
26AQ7X/2mtoRkWIKH/Ihb+f4QO7iJWb2gB8+9T5kkKUhWU00X8q5yT9ktv3jc/wO
I6lZ5bzr1kH3gJI9l7kBVVJIu8msA7yrnPtSdtVD4fR5eU4iQgD+M0lmDFm6/pKO
bZV3ophW+wN8+UffkvwJ8Mr1qd13GdbSFBfZmVv/RSsDhFzi/OmA5wbNgmKDv4T7
B+Xd9j4UvOfghyIPzZdotvyK/xhi6OJu9fmWkUGg7k7LXgVtnrgC8bUAwk2H6CdK
SYVbdp+6q5pGnkJH1AruhBBgtXvA1LtOrcmHbdSJGsgm6P3TYC9L+q82YIK9lHOf
wpYFCBp4A4rlb2lqDQDdZtCfwKDcaMxCtVZ4V6lf3lLhdmYoDu5TDryWa4HxecE0
9FmDiUokoWfXFph+IUvuktDYzRAAgXpWE0BrN4booV/r2BFtTe4kFFADTUs5tTU0
lGRTOeM/Rfpob4XhnvWTNGqQkVBpc2kqIgPAloT5K38kRez9ShJQB1kJm6I2m+5t
4RtQZ4ZnM6oh5SM1QvnP75cRjITmE0rMU0X59eqBEqASNZ0dhtYpj+XeV17+U0DU
dpXIpAqYbL49XIgX9fnM+FowsmJrrJ/qTIiwHcmPo4v/4n+gqy1JFoc/86fNubo6
ed1qWpMlq6rNuPnlF6/nW6+YLlnEJ5rDNYIn5rcx1W89QfNMrTHSDiMCTg2FNcrs
oRrDghN3MWn53A+q8cAn5uciIrowZP5ltTHWYVo7LWE4i0JTDBCvbQv140rWizYy
IQCQ9nvECmV6zHSAK2U9o+4lPCd/1fO/W6KRV1G59/FqgtJM9orlM3zx4LO7DAOU
aZJszk6knGR8LA81/9Z/Gk3x/nmFQVsQHjBKAY/Vzdu+1qMdUWphHdPajSwlFQN6
VcFRQ4uX1R3kQ7dQ/uGrpFLpvplNrn5MZWHEx6Sj8KNlJ/Q4hH8+CtckGShaLFdV
WkY+JOJsxkIvxasjNpeGjz2iVD3U6in9HI1f0aJTVeeCXw4tqO5FwY2RlCYMeLd1
WixH/diRHM3LWKdXqMkiMy7FFnkVxTnSiqJtZBa/rOCnITFGfy88KZo2i3SuSoV2
QBqMtlE4neW897OmR3/9th13A0TuksQBc2zU4GWzGrg3QUq5amFY8MYgcvALbz0I
6AZgUZxZmvXbNdswwJhYjcLC9KBMJCzuqnFhsOWbg2txh6MgeTXNQJDBagUG/HSZ
LhkQecEB3wkR44fvWEP+5doJW/kHIsrMrZC1Pe6bsh2+s8RQ8qMaAqr9zMWwUwbN
kgF4Kaunp1Zek9pLQnIvwSIYhE9bw5tqym8elvwE9CT5QSlCW8FMVhOyDGkhEBnj
b3g1Xuo/kozaaUjZ3nG4rTIP4KQWgCCNZdQjRmNxT9lpGUfyYkcD9Buj/lqbZx/d
iTqePosr87Vn5jclSF73+6Qdt4V4gWKUqBzJtdCTjFY5XCZCbP91c4UqOCb5Wka/
hlYvNgL9ijkt125a1deY/NqeVC05/H1Nhl7LlCbO15iOIHN8GI1mg8knpae5qsBf
7pfOQFBLtJEIfr8QyIyXFazrKOuphTF0d8sliynbmoMoNpLe80f/EkE8A33V6Y+R
cc6FQ4fRKmPpHpbKJAIwEcAkbtLLOv0gEli6Cb2WEJFy3EoXqXF02piVBGTFkdVe
15FvdakWL05MGXkKb9p5Usd0Kw++j/DmP+vFTVaVrJW+6oMUqW19Syw8IxpdGaPP
4Hmc5tEICcAJg8HVGfrJiIxh8VcCQtc0JYu2Guy/P+SVKOrmS1pgcnyPUpVIdfDX
mqoKJH3wt5qDabJl6ZsJlYkjDcTNxB3lkStLJVGUpjEjLO1Z8IwKIyzlp2dZEDUa
4NoyvFS2QUdjmfbH4+cq60v93GdZXKeqfGUhn5njjadmCddFGpzJv4zzHBY+iVm/
RiV8VLLBarYENrk02scXMOF1KgB7+A7CpzRqpEaQyKS1bkW0RJV75YAwSMF5PxMn
sf7FGOfaFV4ee9+g8OnVlEgMyNCcWlhP1Qjoi0G/MJnGJBKd9omtPzOBn2I31M0t
hxBCTpMKN4TpHz6lJkh4sQ==
`protect END_PROTECTED
