`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GjREnfE2yK0kRlA4ChKtr5wI6yEvJxc5+QGmdogBzl+dhclRHZAYWZiesUe/vfpI
K0unx41VTUxm+0uEvWNng6raBAcP/W6m9r3WcIigQ1tGOSBnBk1f1nFXvH9Rd4Ss
quz+eDudDv/OqDDiudMOMWoakVKCdhEZuUGdrq0PHvFweJ6H2LhvrpRNNv7NVx2N
H5OV5CqF0IQQ5m9wIbkYIcImA6/PPNMOwpht1z0Mf9h2xzmYLuLAYIft8e9V8aNV
xmDgc38hAjp7xZp3QMaYxXqLX8Nqxwr0x9a1c8xLDSaOSEdjmQo7ek2P06/65Fds
PWi9P7V6lRocE4zY113BryknA0gbe58a1pyEXAdBNhgrv9zR1u325CWX2JdzEktr
M1dxXwiwCH7yQNBJuLRKr06GIYIDZknttrauo+qo7Z9N3aXNMjZcuI3WRvHhAM2C
AeSc74XUcgZWhplopoYND8ZLV75yrjhZVp0zURdb5zsYJZAxZcdBRiRDQ68awXjW
lYf7QELIDwzyNmtmYjMvZpiq2QGqYQr/c2EEK2rJQ/lFkXyQ8+Uw9yc4Yv1lRiPU
8OL+5ETFLOTFPxAbdzg1iufTTOFjoVgJileBPDYkqPKrMLNVy1BBmf3PLqKQXyor
H815NXRW4fQVwoj539nUJH1ZoLEQ2I2h/msX1PmBGBXXOLZ4ZjQ6Qk8n+iyuZbV1
uHmdOyOpvlCu9KjJ7jLSb4FhcJxdRFItTa9qgZY4zok+dEmxwbLiu13LHMNgFmiK
ejOycby0I26xmdNptE2sfwOjjboayWN6/TT2bfB5dR7S3CyQYTdejtlRxLwtT9u/
CCQ84C1VjL6l63WjchWqEiFiE1bJFxthDJ+/onuSaQjQu5KnPiLJUByIaLKVjR/x
Lk6JsYDGRxiDrrHmSYfIaGcy4+FdcDc1/RHUfz46Ki3W+6rKD644YTvXHqPvZVck
x7MEcZ6KSoBeTindeAfB4+4vuccgqoUi7oQklKbQvTCDlfbNZu8PavcbuQ3p1KoI
LYQzhH6ivQ9KVyBEK0QmMxHzsvJmAqljPtZzU1qPrfwJwVHD7fuc3er7Oop5txqP
M6f2cCqxBc6hC0bcBn0g6vj3BicuSw6WxgBLVcRZaT8QPutQbKV6YfU78VohmbPg
y5d6DlAqdly6P1m98hYNshE8o9Oo+qNmuU0tQJttds0P36CHtD1OYGj4F6ahvM6D
poKJX0QhWzZyMc8SaaPmdTjBZI3Csec40wkdZp7G0tRIsiPxYuVKvjfkNmitWM9N
5JYa6sJHVUK+YKLouHVYsvklWDtQj8tM6nW1N03xL56AQ8bb+/8Hn9OfhAOyqXhk
IlGdiQwWUarcP/APktm5TrIefZKOSqxZIRgZKucdMC4wz8ABhFAzLTEBCeifECvD
Yt4RHGskiLk2iuEQB5o2NwZQCc1KAadUuzTxUCKmMxrGB6XmD12FjvgmoW+H8cUr
XEVYgsLnkZ4wWhc9sTOh+MLiA/POhgC1r6Rs7TiNMII0Tb8yixfcVt1XympzLUgs
`protect END_PROTECTED
