`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0BuJtUF3maNqvWQVO4V87UcFkur3HGEnU7yu11cJi+H26j9pS20anMhnLnceqXWb
i9YWguxHoWMXskmF+F/FIBf+pOrC2B3GiztSn/TTVzkStaKWIBFlYDiYMz2r/H1l
N8Nnx/R8n1unucvylx1wUPEDggKj4vOkCaatDE3KRT5OUFuJtER4NaeNgfOi6X7a
iIAXsP3vGfDALasa1RzvoTk5EBO1UQMoFBSRmXCL5lO0iVapak97W2hXGQw9yzOK
0tURbzvdgGVSnDaCZTuC+hg+CH/mOXwcUjI/gcnhdcRZPK29bzriiBDQ0sbvSYXr
TzQuMKJsQvDqkZ+0d4baZgyLEawJGGJU7S0fn3rCvw483hzFfvtNsZYhRSdnQO1T
pG4jA9Apw9nUwXPlWZQWb4Xsi/e+j9MYaZnIz0FarNsmFEBk/7sl2P7IN4VcfsTa
dkb0pHFYXIg9nys9EUHmhap1qMF1HxtHGbF9MzrLS8+AZcyO9HZRJEc0sY/xYQUs
3muF/0qf4OVMx5x2bSbPak+gwmMLHy5zdsOfhqCOgnVgaAd3wgEZ7UxW+Z9OboAe
dpb6HHPDjDDpb8JJ4NrnkB7SUKMtAwvj7FrLVODIofsOr53bXAZNfAqlDMhWBRcg
sdQMSg2SeMPb9UsTJ/fDglBJAtWEy4YlpXnRKjNdq7ZJ9DS7E2n7LQHdtEh6OmC2
hBGtArHH00kGZYmzj8AOXQYcdGdAoc42sTLEwqL9XmhnhEW8Wk4IGfgYp4Lk3g/F
jEHyciWFx///ZbOhDwi/8DKoqr1HgooreooJUwhSPRS1XjqhFccxV0koaXKTfCed
I+s7l74BBVFVIfQ16WT5OpKHB+Rgprr8hqS8xg7SMglAAc7B+pokNvUwMg5U6e7y
ghl2+rwT24Qo981wsUT76mhVb9Wk95NEIYnYQ9glVrGaIbZclaSHsueYYoTlhM/u
kzGZzatRh07HOi1vEFb4YLBYKBUiLnuQauyLIQ7u56zMf6EISrL+UzaxUEeKwzdG
uekMhC1msjnY2tjSvHsc9owDiv6sD73yq2gNfEcHuNFrKJ60hPpLEP50tI8mBvpg
oG14HMDJ/hsMPDbvwF9Nqkve46bRN7vtPGaXd9Ns1G8mbzhd6BUjJ7nb0Vu0Z7ZH
iNvrMC+kGnM2YUDdL8v0YeBpyTLGzps0zbO+qjn4a48Ec5Dyt+KpgMMULH+5d2f6
mDaPBo6WoUBjqPphehXIdhDmI7Fc6RhptH4qSvhCQ7p1iacD09i+geO3N89cMPIL
ZxXm5iMt8Pah5ASH60n+j9eCBZDVsGBtIos1pVa8HUgIBdyPcEAQ4aWZ622UJWe8
LCrIqd4cMm3679ZzTVNpcbR+DEWV65qq9PdSteh239FPXLp7EjtJlaJmt1rhjfPu
nM3CCMxaFm2ngNIOgZ+uQhKLCT2QjKrfj+KIptdK9skIhTsbDzOZ2z9PeyDucM24
`protect END_PROTECTED
