`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lwCIqR887TgSyhiV96kOwxfALnFeOr2XMg72pbeOfg+V9u0FMDyszvjAn4/qq16i
8BGV4S0Zee0NSyxSjIP3Ti9H18hBVLRh/0V+7r0xv84tmR/Qm5U6CBk+IEg8/1y6
mhCZn3i4cHO/2uWxj6/DBFi6ZN5MV8oB2eEl9M5lk8xNxpqlkvroZkRQt+y3qeB7
ZLrjD4LfynqZFeO2Oq0m5q/+t7oZp+QckXhrTdwniJJPscApTx6IcpXMxn89GKFn
NLFBjZh4hgCaUGm7Z1pPqOcZxr9cgxocsbKJoXBlXczx+XwqT34FbSdgryIOtUJK
B1yaN1htUhI8gQEXr1SzCVWbcQK5ytr4qrC31Z30thFoLXb17UsOZCriCGpy7Qjx
KkzzzIUJ9Txqv3f3w+BYpENpos9sMjIYmOYY3bymVlw=
`protect END_PROTECTED
