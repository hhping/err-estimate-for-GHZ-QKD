`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yRh/peyPhzqnIqG7yHwT0rNRD6XWaCONlrewQ+GPQTAnbrGDxUNNYe6gE0C01mJx
vYdrn3R1LuQOwEznRonF97n/AK4NQQMng8eDlle+1YwONxI/VQTLwW00o6oRaHxU
0SaO0KkiYwWtSWWIhriqdVg80IhTMgAtF13iKDRQ+xaCr6uX+JqlYd1s1KPeQ/si
ZlERwtK/cXt6uq3707bPrIUkAi3sP+vJQnHLBlbyK/XKt0VWxCT6MVdMjWNivQ4s
C2JFHjDczdy0EOIN1X4Vm2geTjsPuFxf3AFVcviuxXeiKyiZWetq3l4PhA4MmIrK
+U4+aSTkvM03GY2TfDcyEmWBjV6YJqycd9GSTiFt2htlDuge3+993r6vh28p3aew
IUvD/p3OThX/ERaIoLuaJ7lEU8daRm3AEnjLO8i+IfuVQ94SB9yreCAw7zQnC+i/
tCdqvBNjaJAZAaBQrk3HiMFuF8pBtFvjVavCV2ilqsRuCV/brjLAthYBhkBECLf4
YkoNB6YmEzZxyU1g26E56yquXPQHNEjtuDfkGY4vZw6V1sC8jxU2osMpijUqyylY
6iz+Jq8v1rymxiUZUi/4Gt0O2Zq5TS6+Nw+5fcj2BPFOD9snyzRyHrpPOCD851Gl
qk+2kxVkqFTzFnFEtd+iXBIYXNbCGhPAtBeYIEWQ/f72KXINKeuTCQCferkiMhCj
OORUhT90lufTHFLh1zJ3qWpebF0ByKnxWruzaMEljDUs55X3VX0udTRWJXOZDI/O
gzTVJiHhj3kEqtzO7IUDts4/NL9PbfdOdP5cP+2u57JAoPOz4VcsrnjUEbrjQY4C
/YYGdmsuqqZfgGvkerI9Xl3c5zZQl1Ci8fnNb9lweaN7T02HRPRFkSScnOfw29i3
DQi/Dzc64ttpXgTLX6QJ84P4iNizbwBcVrm+UKLcYxnMlcSAtC+yoa/CSKTXamWb
KQoytk1YwfnVaUJfelgOgA8HsfsAevy/Czs6Rj2W1YNFMqBuGPbTENCm5ujwNIc2
+Sh4HOGWqUG4AzJh+3uZsZIMOW3Pfg7TibhK6cyIhhx25bTd47iF6Yyd3qhYmMRh
Q+2yzn5gxRieiqChfiOJm+GU0C/BtWqXx8l3v8BvPUyUt8e66/aSwk3pJ3eQgBlo
nG4oHIamunVoJTyqa/ucn1ZKnU2wSP0D8IRW6+HFAyAZRAdXvqpnOBovdIyzxQI8
+WZzFqlVb2XYH5jBW9EUuKlIdgt4yiAqbYpl6FtXXp7pl5u2bKEFZkqN882YHkmB
N0Zk0VlpV9cZd7QbklT2bBktrj26A/5WMTaLtPOb5XGpwqbns3uUAu1iNbREP6nu
wS4BpRnL5IvJe6I/zRcuBrBkRAhhs/5eV/0Tn/Mjs8jdNRo9JaBs/l2VinUQqIoh
FXaM0F+MY6eAnADvuiNjDItkdaz/BVDbcdXUcEtCwjLf3dvfhQaqhbPS/0nC2+IH
roLAz3EtCHL9xHzG6SEbAPAruVfZWDkFk0fOj63DIRtZsWUqQboCrPwVHzNevqZk
6zQMIVrIZJf2blkFCrKic2tWPqf2JBDmD7cTwA5lU8Abedws7M4F8q9a2wMrAfX9
8r22C1mscj6MIZPfkdMeA4KxiJTpVrLOtGpCpr3OIr8jLPUq9oMMOQfTC1usphqb
rMMNvf6lLDbMeLHjGOQVaTDvZxxE2pOzuU0O28KyF8fnUn8BJZB6nSPxer8tnDxX
Ggg5KuT1wfvGGLz97OXoJtrX1D0JcZUu/x0lt/nD3XpjOY0SyFBafscxRtYC556c
98jpsx+4G50YbtF168+9ZfK0zkcZQrUDD76Ldh1V/sGZhuyfKhL1KuDZd8kuDLx/
b48Tte5WcE/fBU5rsl7m85ArtZtxarEtz44REzSUfKq9Boo48xVOCMDAPMmHA3I1
Nhua0qcUk/znVXh0qzV+9pkLe+A/BPisDFR8n7io9XFyZLoU2tVz1ZbPwNA4DP+c
DQqMac0NE4XsN631e2bBjDUaZ4TIn75yjk13jwiWEr7CD+TZCHMGFH5OpIT19K6z
q7Pp+XF31mjmkyayTa98fcgIBgd/UV23V1r8J26RCX5kM4+ZixT5HGk3j0hjcHZa
OjxwuKb3bIx7sKqKPST/QG90JGC+JhJU8P9W2gSOcZNSiGAtwNC8LLo39eW70V7N
4OKGbnLi+Xt1NBDFeUxbP2c1ptNkGAaRWDfQiI6Jd7RUO1Yt8jjoPBlksSxBBSUh
FQI2QyeXwEYST4DvVsJOEN2kYKca3rE/ZATRUJRmdRsu7i6fM2ytBQW9b5N00L/Y
i34B+aDVzJWoDpXZ0A34bUKTLnYwcruGidnGexSQev+oXuTTgL5zrLDNJpxh27xT
Vl9UB6L5fDO2ehKfbMe3SIvnAaj41cz20rXRjRsrsSArdxzE5EN+FVVUXiYHyGDr
5qhar4AgT33LqNckvand+CLISp6aH/EeVfL93fikEs4Bn/NdSN+kTE4lUhLnz/5p
XuR2W2wbQpvNwkje0P7+HDSWtFOiqEV9kK4sTrw8JXsMXRyVdAdWE3B3SiAyD8Ny
SgBjiLEz3s5tTPX4hScjOX2E9rEGOSODf00hZmpDrt3QaI3cbv9RxJLeh/ScXohq
lDhLInpFf+0L7CWANNdKKh7pxkMvCsGoXKRIylFS/JrW5bVRiM5RMXhueT2DRbCx
emsP7Q9lvPx/cN6B+qByFRWghZ+H09Odq524lZ2CjkkRsyndffvxBfsQWe11r7z1
tyBmpEHAXl1iKEYkRrkOxItF8v21vidtxFSvMMsh3K/EJejwW+wCDG6anDo1Ihs3
KwFT8RNukyXj00ystNWbqlxnIyPqQBVqTwfZrVBRqhhjBSQwF2+qGXq79+M/pJRm
9siyXFxHgpaekHKSwCQuq8CpQ3SNJBElXjnBA+A/qQtloqo6oeJ6AM6zMGgwczUj
XnWYA8xPWRMHfnTrLB1rM7UH4bIESxEJUz2W8PeW2rZZ6cfXZc7YHAz0B94qF0iq
zBqXQalWU8mcJTwRP2nrxJR8mByloZ37PvAQi4F9M4vV7volslnPLOA4d0s3UvSD
SGMJjL/1Yu+GkfFIkEp21H5UqIdanj8ygp7uZ4YU7l5B5St7PnLSIfzuHytRHKL9
UqZK8ATtAlPh6fVuUlmeO10uoy0ExoyjYcFS3bYragABTMbr70mVhU48VT3tvGFI
QN1GR/vWcYW4I9zLy4ZWji0o/kaow9AS8U7HJDbzBuj4uZsWhzyxBNcIK7SrKDHS
uEnVLZ3fDQpwQkqh2vVieAp/kiZI9W76N5bS63D9Y08ebdRDHZSGU3Obs3uGYP7r
V7oVkv1DSesMeu/7qZ/XOGAgJoetU+dsY+srdebPlv+gY8U4ruNwFN9iWM+HPm94
o8kMnN8b+EK/T0oKa9jo6MSYoTdqoe5R793WUxXGVea0lgoS7MNrQzioaMih8Mql
vK16xYvB2cTh28DZq7kdkJDgaMcAzXLNmPt8yhAmxPzyJlBXUruCIqiL/aaWcR9Z
GskfMZnECIWiawgxDVO4V7miBms1pEgSLNCY3DS9c9LYMTpyD9eYmhpEH36cokQw
EJNu45brzatwZ0szpUsx546AnHFIRB84cPspXTXgYdlUdeBfVzwELvuwb5XBQ3Nz
LnpHvlihi2yevFDb0u0lBq2kHXUsG0mbJKaPInrs5CEzxA1e3hZlBLS0Xwcrn/Vj
ltuy9y8uXwj0RVBhtsIqYJFwG4nE7i8fenz7YkAnaCtkR2dzASqNljcH2jLPyZks
q7ZGnzrTVZ3x0jkpg/cxG4vAjm8yGPP9/Tx+lqDULm32iraTVEOKnvTq0ZBa9gNv
ZkSPFMo5vb6NfmTAW0F5Yg==
`protect END_PROTECTED
