`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L2tr9tv1RYZsilGwB/0D1q8HFVoXTtqs5cqLGEnGQZ2CuspS56t/+YGarFIwB7co
GsH4i+fmvq9SVOM7f1llSWJObqSzP5sSh22OQqPRgRhqRxLOPIOhKhanbrwK4wQ5
jiv9Wid4ovIpiE6V8bPc06hWqKGAc6Grv8xWuIMwEIrMWe8kXPw4+svQu4iZ2P2O
8MvXoGlLgYJqVf/eOHuQvnXxYQjfR+C98cvUkkYuZFhAHIYiSg09cl9ykzO/x6JF
GMDXSfHko/tFf9y2BCYXMVh7pjaMULzAIvAQFLvILat2GEHJGnQAOqOID7aKkVzW
pn3xMGFAYcHGVqSjGeKhWdG6LBqK1+x+qg/Zgp8UmmNQbt2DaNT8OZ7mw7OgWrWm
dE/JTc6BxMQSc0k/vSWtRl7T0lzfM8W+Am8EkMsCZLMgwBTGtOWnY7F3sI33m0EP
9TCOqczEo4mKyuhrRfeQAHFfmr7MiQWbM1dBc1TmmYDemqlR77CUhXdn6EuRxgcE
Ps6nb93VXHMmVX0fBpKqATrGMZJOMWaM586hY+sX3r//k+NP0RqFWjZYfkjGj3TY
2AJfiRRI/Z52+S1i+x0+AXkSv4RbWP6eTcmdA9oKeVKllKFVmbnMM3wvFx+9Fs/c
OpG9+GanH2fxR+7hKLaCRIgkYF0sDpofcQZrjuzOaYVpMwZ9iiig22b0VKLWNhfm
qoB32X5NfIRKbXuSOEZzYQso5rgLrKk02K9XRHqAaduDZHhvacffrc79lXgp6DXE
`protect END_PROTECTED
