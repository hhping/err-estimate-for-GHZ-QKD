`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HHNSxSvrtAsuID0LwWPrZqeVoxSbBnilPWq/88vVJJCx1nVIGvs1q4lwGJLANU/0
7KxTH9vNWyKX6tnCir4wXM63mug6/13BbCRb7iDsnEXvLvl60A+ztXiAImy98UXw
PHdRK6ZHAquJT3MaEhuwdncFvUl44GFnanNMOmqLKwHIhreu0YYzLAePljcSCcKB
PfmrnhAj7gF0WTsqNpjbTT0PP30C+Xl6ZayDvkO3zKV+yHSlXlIHunDWfAu7BVN4
ZjSpyOSqd9zSp51uiwKrd0qbHHwTvnjYU+6PKvt7D0oHbbBuZ0ekx4aC5Z+W1m1c
Grywjwk4Tuu+zz9NwcUG5C9WL8dlkN5tDktobYZHyPS1Ys3ReTSU/c2RwuHs2bqJ
`protect END_PROTECTED
