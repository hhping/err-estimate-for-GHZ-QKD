`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V53qi0EhD/A4MNZXum0gL8lM/GYPQ5uek7Qqns509Ojo/DYWVRhwRzMvS15wcMLL
hdssMMsohjSV6BpLw8FrRWYmQgd2Jgf/fuP57J+v0fGenFdGErx9RevQXGz5uYuz
v4BasYA4O7B5HOaGttBRMmvzFJvEr7LzqhA95mjIsvSeiaiLX/QtXzYa5WhXBOAB
SRakOL0EUR2tUuRPOhE+K9pOMoIVNWs2aUV3MEJRRq0Mi8UFTSquTbd4y+4ljBIV
0A95MHRH5ndowpJ8diLl/k9jHnwX5TcvmkvdmO+vikRWUB+soQnwCz+U4Etbq3F2
CCrQjBsrMMWyn7dlCT/qXyNdz2MqplHa//yIei1mNH/z6atvxMbQ6SW1BZv+4euZ
`protect END_PROTECTED
