`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OH8b+R5x3HD0TblHd8BBNXZFMSF07P8zk4ELKkGy18GLZ/40GhNhnCdAIxXbcHVV
VoTisFv2N5v1VtgncZbhSsRfzRAQzh5U1uN+pRXa15VlXtJn7l9912NuGDjvW98E
0hgulcAq/+1LdIxHGjgluzERX8l5DSEA36Z5pnbs+qVNXYdWfTRmhQ9RqQ4TkSHQ
PMogLRBZqbuONOXU+GBrZlw/31Vt1dCFcygK91gmFoP4dy3cXV4yvmOW64OHD7T4
Se6yv57sYPeHnDwqkNW1qsJwQkLbVnSK68WyIvFi/BvTMNS/IeXaFRs8jgXd+V68
rxC9uCdXzuwctw88ieuJZaAnEDENDpTn8H+jBaWeZsNiJvwXhJA8TyRoljt+hk+4
4rCSIQqEKmn7XlBd24xn+FSy6Z9dIqOi2tnFHAbvshYSspCIhSEYZEo8I1tXS9Gw
ygkreQ0UpR7dGH70Sq7Guoxr8cSAWAvWEEriGEimx+uCP67URX1rEH1XNSRxUE09
ZnpB1q101z5P0HuRqky4kFxkxsrs7Q5WbAWqetP1j4e07FSeb81jjz+64qi1+4fg
mRagitJVn1GgV2bXvMB6glbv+wpDZsIYfW1HmfSG0qFqliV1ime3fkgg5ucR2Ztq
EG51LSPD1o8NYbl/pMMQVFnQ5tTOsevjyK3LOW4y1pmRWX8t+sC/5ae6va3pij+x
pbdUfeRukI7Aqf57hcP3f4G/F7ypUTmZssIdC+Mm7HxkSZXSk88oVWykwlFFT95q
bmrXIpYrGR/KLyWynXeinMkvNto2wk0EeoCLTY3sF3EWw9L5R0or0X8fuWD/yVx+
6ljrOLH3Mh1ANnAKRYbtwYTK7lHaWE8ik30McdFM+sEuGPmSAiBXgstusx0xyB8H
2r+H5FGoHstmSBUB9b+pJ5scZVm+gMfIYaX1c6FaCIT2dmJXyP13rbj7lPSQzWNk
TsP1GsyU263aR4beAapLcas/TvvC1QlsZhGXrJEAbXYZFAxq23FRO5lfC9/yVXXd
ikaRXzTfxur2kJOCm4SxmoW/SpyV/tvpdTDYsJK5oH1ilZWR8ZRBzN+0Gs/uYUUv
Y2MQK7y5hMreWFTdW6XlNH3JjGIviTpLMZpu979volWfpd+FTGKg66mxmY4aDVJh
BX10Cnkx4GmBp+/MoOJ9mr0OEaOhW7t1OMg/n2X+7n28smq4doli+hdfBYEHU3/x
g77wpsQin+ibz4uIl2dbhnfb+KYRpcgtFqX9sPgXnjFaO01J1vuzVBrWep8TgYAy
inu0kk8OsaMmJRDRMP3TVa6qcVm5m4yfZMEwzKP74upi6BIKBcdeSAhJynXEcCzC
4qIjL0qkANwqkchJ1U0EQVolE+rrYb2NJ58n3qHVvX3/NpAgw7B5G4DoIUfws9Fg
EUMYrM/W9bHAIMv5rtD0OqNrcFDuGQ0t82F4Bz8lAmQN+YchsCbf5dn7I2IDe6+l
ptQaE9gn4+V3DoSqINLVWz/2l4CrodVhUrXLvgBdbgLOlYm8cYVzBlNCebUzlEhz
jNcbIq3ew/Ms9lWsu7ZXHuuup/5KS69Ezdj0ZZ7085jJQBQ0SH8g6Mianoq/XZDl
OQ9yyH5iPOxvG5Codmt0W7pdJnd9QWdGJaN2606FkbVuut9ihK9ufYMGpPtSHsHO
z6zYvACf65pbWtcxbcFT4rE4tC2nm2QP4gL/7Oa0NU0zQx0hgLBsDX124sSkfFsn
5pKdyTboszi6lfqJQeWYMMtCXB6fbHFS/DR60wwvt0MTwQD7tK/TzhYHaJyLiIA+
vKLVmWf+2mkxB8gDFhXHFWtSkrMIqUiRgNsC5/I/p4Rd/QxKxZQ1K5YFkLOrAAXq
wHbvhILSFGVPG9UJPnQgsSMyTszug+6xZ87BWu7sxEFouXlUr8CnIYqH1Kw9Te2Z
27O685S8GkDeUyQmubfaV7U6pcoGYczJSvQ6GZcKCUrRPodVRnd2DKyFDTnXclR+
xQ4tMd4ZeqRkmCOEpnM4Yi0GeufBnXRRfzgwvub1jls6jzu1loaa207jiuXcRVmS
vvAUTDhjzsqOAhoffGUntCwn+3EX2pa3bxUGAsyeCzCBp/R9dBhFORopj1wJikg4
Npbt6yRUf1FofHiwThihIAQAIE1pqt6yvpi5/lomAAe4nQXwD7Dvwm9EQEuA+eWB
NKpCFioT7djdT/upzFbMmtUDjnbA7MbjbNRLd4kiXQo05INoiL17r4lTbZY5bWoX
6wpuh55HQLVqUpNl0YkwhvUsu1y5dmUAT2cGpp5IvIMyraVoPXCMqp5nrHqOgyZm
EhC6OfIkHef4hE7d0Qi/8GpyzKD2DS4gE85cD872w0DNV+mNkA3BJzOe+o/5TyQO
r8rQDZlhB4wUamdywpmRaRcxgggpI3J0z2Ct0Q3oiE48s7L7y3AK3aWfazAkqEE0
GtYrpaS8IzI4IDyGXccnKRUwReG+tglNrjNpY6UB3rLpfkVFAWgCXo+8jujfmlXf
SFmP9iDrG/r3pY5rS5tWh+hk+wRPJ+HMfFIpv0RkE/JYAt8H+lfDRtSWJVZ+GNrk
GZMn6NSRUme9haAujD5DnLf8DEQCV84i6CYT/EMoBmpCbEB27ckzQ0TWSi3Oh6zw
SiPJDUTpxSt+4ZvJW+0REiOP5cQbxjlmfxAabkugPam2WmL3kQWkijcsVS2WYMEF
CtNcCmd0RrdcYpWaL1aME4O0AyIdhWI6W03O2d1cGX0=
`protect END_PROTECTED
