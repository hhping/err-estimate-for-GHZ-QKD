`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GRIBfCOQvgEo0jGefTjVScpzop9XYNKGxAeopU79FFyojDLE+hn1dQqYQyf0q1hi
BtkCJYdmD+Hpdsvjob0erxeAtczPAlE/NAhxcqQcpxMDwH2nE8aIjhyFEisXBPi9
3v0wpgDGLbjxP0eNYEu+6X7+W9VWWGRli5W5pFGpq275izRLRscD51abNTi3LrlH
FOtXvRxjXOpvHc+2GymmS9ASglTcJYhWKsbXShiqGfChDXGsRhwsVoUH5GWofU4t
WpNjq9QXOOLhSyxe947paXE7kndSRW3KlYMAM6DV+cBZOMRI1WNv183woXo5cUAC
j2QYfjvqJC3EKxw2xGGlOzNG4e8JLHoMi7+5kWK0zXshsPiDKJ9E76SmiSgm9PzR
WOKU1zfmf7wPMnWgZlrlLRL64GmL1u3M2Uv6tzMoZujztcsHOeOdCZsTH9QA1ye7
+/q1JLJI/hpLbftnWGn90+78HTaXpZB/gPaU3/ZYJKbN9q2ZanuAfkKQqU72iYBf
8/c1gJF9bGeplDuviA4X+pJjbjQLRf4y0MdL1nDI1aBAcP+eYhcTCbTK6lukud+R
FsgCjprSIs3WpQXo5bpZ9VR8XpbtKLGFtos9XDe7g6wRU6wAULVX9JfKUlFsT36j
q1KKqUYLgcVVAdjZlxZZ6tGPAWcXsb7YPykRUOUH1kXeyPMOUHkCAsw81BWCdhZ0
wfQbkwxEDuWdoHjd7o5+OJBPIKX0HXTOtVGWt22ZjyXOw00xU5ypKnm4rjVziFor
RqwOL3VxAmc933MUpDY4mxzyD0QTey7zaQ9iKhoLngzUQyBQ57UIhJ4D2yvSx1kc
CJHK3Cz/AnB1tbQWBz5Y3dbBnB6GiUXKyuZO3SkQbRjdpjJxijPG8gdyVYNjwkmx
5aGMHn/QN6IvVORLu2davdvXYOUf9pWxn/xuhhOTELOMu6d+aNclx3M8an6j8iei
xRp8k24hAsV++af+6p9t7Ia5XD8HpTv1arrYc6CM8leKg4EnKwiqPtDzyjsMkeKY
hDVj6BmF88AOI0qv0FV0hzjzp+4AwFO/veNY9WzNMpw1maujHJuUhO0Twu7VEXmj
2ML256xHf7q5O7Jx6ej/CFS4WVFCSFqD3ku8MiiPVLp9+EZwHN7wrKMLn08MIicd
stYhPWCuW5NBSKI0mPKhACc+YeZGH6DUDWiUsWuIv4qw3V7neNyK33x60C75Mt02
7sc6nHGRMSaOvESlZ3VqqbDDKy0Eh3gCqB8apE7dREN22U+IgwP5oMCQwSjcfHXK
DrTCjORyvZd76WcoQLj+ghQyAwSi+5AISQsKFaYdAmE88fh9+NL73tqeLWxe/T9p
wdwhbLrb2JGOzXtdBrBtx8NWEzvEsgjjPcDnOHHd85P3iG8JB2a/49VNkLcB/7rL
CDeFjvutRY1L3Xue7uLbgUs4pTveg8UC/tLzFVPl5EdMoeTCoXycR1vfUxo+WhTS
cTqyEvJqS6Oa3tJME2zb+jljGMnIqGl6ED3MJ2rIjvfZp10AZmn8wQq//46cZ9S+
3UKYm655/Q2WTiR6LNt7OoePY/KhexQb/6pRVq9y8jOhozVPeR5fc/0fAGUivIsk
yLC2tW5nObv0w9NNjNHgUYk9cpkuvkTbr/n1H26RbSD3USF6yQd7ax4R++Zudh6+
4FX1CsUfV2eX2Zq/lkc6sMmYXDy4GaJaFWNSE+wjZtRwttpyoj0clT8XzmYFJo6l
VsI+WmncaU/RDedP3xg7slLP7l4Cdcje4IcCCwGD88Kl4KyNXtxe6In1z9hOhzK2
ZYKoqZv/h+BGK0MPu14aPGFXkbOlZkU3FRCLs2mu56J1tT3N+yFQwM9n9Ne3kaDn
WSddBnDHy8zuGeSbrgDpeNpjF9BYh/YrZbIwRFj36UVtYKOx2jlnChy46rGsbkR/
LEQLkw5/IfebKe4MpfEZxrQPsHb3+cOSX/EbM66+ePUhFDku4Ztw7MVpx4irQl/q
noAoiZ1nE3Cx4VUPGxR9fgKVoNRQd5ju51u+wPkgHfIcBxluZTAJQ67+6vD+Vt1j
96GPYW3TrlD0S2GGESdO9RulIgZPN+y2oIs/fYGALFKn9RzmALecZRL2dJ6Ofx+0
LaWVO5wu15pKHhwIbcNfVyyk33QWLKsDCjwzXRttxl46OfHX4veCcYkHOZglb/M9
lX0yZ6UjB8MqYsT6xUGRhPfaNnNPNtpDvP59bsRwP0YDkF0M0QkvAqTPxCxEJVYK
B85KOpIRTwKI1oBPsjX64cTjDBC7B0aza6F+EFUjAy1fg49b05EwEC5R5xClKXAM
2E4tsgmTc+zuwy64597n3Ck4bIMa7d0OK355UhCoDiD9Xn/IPcG+1oAfFwjdwedd
xJey9bD3fmLDIqi70eN3vNKBQQvZYk1RX0R1diSYYmFjukg6EGeXlczO0qAzviAB
x5P0jpR9faQxBef5taami9oC3ZZytKUOW/gWFF0B8oaEdOkTM3atdKDRSSPXwzZN
ZE2/aqb4ro+WaijBKi3dEzAHn9xujYNMe/no13jIrkMT64TDkIRPybYv3OxRek+t
AJgagJ5eLsCDAeVuQWHbfuhLhp2M8R8HzmdXw4Hos0Mahfv1e45+gA8e0PDl0Fn+
7l4QX+nHgQwo1Wcarfhp7XgTyqTNSj5rDMBwf+4ynS+J0F3Cy3O+DRXoRP7RAEKu
CuA5o3UBO4DoMogGt3Ze+Qjul8ZoBslbqXabjF+FByIPx33fZ5+W8I9241sqB7TX
u77H1E/EOKQSmM9Tdy3GQbDZYuCBKTMA3jZiVWNn88P8knT7Gd7MFCuUM657Wc4M
nLdglk7eDVIhY2JhWQXvTjoxNax4JRFRai6m0P98WkZEim3Xpi102qugZly8PJiy
6aNm0tR1qAT73NfBWtLTHBLWCxxJ3nooHxdsiZz3zOTApOaLMrmJMymMOnDCv++7
0dU2OEUzQ0LGF52+kwJywPXA5f4EJ+5P+gPdoAxeHzrpfg56zJF90dBbh+SjJt3t
3kS5d/cMOoaerdnx3vdV7sw1w5m3VUG2KUJ6FQP6rJqpIFqbMsaXUTlUmtC4bMeb
uUhS1V9b+o3Zx6sd+YkIQFXij54QBt2msHqWAxmWodvbSdfAlnEZLRIIoTBgnMhC
184YB2cU1Vk3/+Tx5SaOJpCdTLIR03XIab1AKwP54b/74YtS/r98pMoLiXVvy+uL
lvYU+lvv2WpG4H7JUSTSu05g+AINdEvDdyM5zen7X8+nxuZZzhgQy4jkKDIkv9Tu
e4cmG4fREmJEiITMPgnfwiKziXC75X88t3K+dKJh28PEGZ8PUMEwhNVnZjQcnn2E
maVik4taCU8ey1S7a7tTXrYZ11DMxmP1JcbvEix1EZafbs5Dw766Zrk2W3Z/YWbc
+8PMCxyVRMRbrodbEpdiq+8s1zGzfCtB6p6Cwusk60rRJnmOT9nPT9Lw7eWF21ME
wHBK/aF9looJgkXg5PN0OGlVZjiMO+WgHNho9QAzN1ym52bCSs35bgUh240zeWCA
RogUXS3Lg12r6b21AZ9sJ+sNWtliICnc7XqzJY/VlQfC6iUr4wmQ3Py8W3pcvJSk
ibpOBrIFWSXY/oXq/q6QBhvAzVe2L8xM8RAgo9uzIQxPVQjlkKYTTEhBj073p5GC
E5mrVbL8L9yduxIF9xrjHmUvXVRNao72zMWjo9aU90qRBzLYqLDD2ztLWrtMYTfu
xiVAVotIGnbzkfUbhJnLEk6/reUoJzKnOtT7jQzOP8xbzfE/bUjJC4zkb7jop7ei
IHBC9lfUbye+US8Smre4R76km4zXnLkeMCfWZJha/5jl0PVQI0vQQBE5TsBGPE95
Ne8F6pMmDWQvfas1WIhrnhpWw9/TyRBlCSz1nzLV5txBcPCv/9wIE7o1ELdleQrG
sxyP/nknDg3UNxKc5KxlCO+FiWkuPpHzBoy/pSBatJmG5tHFqVr3sOsHjqLOYMsJ
oa6RM7QKshEqVDDcMitY8wu6R3B0iDIAnKRpFnmyagG0RcxKaPIDsS1CyrxH5m+p
rfD8D6CWnEsPDxbyaUIMSLBCDZo7HVvDhcdzvhTe7EVnPVu7HGe7iYeXISKqFMHd
mceaglz5Kn3fKCvkra8b4r5MYAzHYvxhLBT8kxCNoMf/m1O77wCsx4NtX4nJmbmz
hnwDtmL1xnSPGns4HO9phatzKmm0dxD+Gv1YkmTvx1jVb4xJWTVgsD9XrsuO3138
hvZYzXL6FJnqu1dxea9VZsDp7MWsfLt3CAxgROe4KbbtRNq8M36sDhdGThgOWWEG
19ypgZOa2bd58l09blaXSYF8htRoyWYPN03ZV5R3rW51aOQ5ZOccGfJ8A8QPA/6e
xqpznDHWSCamU8jT3XHk+WWsnYouHYZtzbnDKbX+Z0aP77VB8mEkPyFhFlU1EyUg
y9yUcu6pu3pT0yj0UPscsziIhcyEcnfo/JNQSNhnLtD9OtphUb0a9l0Nvx4o81b/
982qKloqCc3pK9FV35tZdpZprxGsVUyHT1CB3fI4RBbYJ2iSHigeRv39n2BBr2eZ
AOBPb7CIb1Gj+/zchzSWHq8eKWd/RxpGE6sD1od4BbD4ObbbGZZ1GlQBGlkN1jPp
EBmgiYilpxk5QgoDAx4wt0jGpvtxYtalCcTQp5q/o2TSHQyCPTH+3dBxCGsVA15D
3r9N8G32wgJpCp4miFjj7gNTfnhSglTQxb2TsjM/rs+ylPSqvpNwwjKHUcMJRC6P
N2XO2v2p58TqoFIi+Jbwx35ispwNxmzD6J4j9rnfdADDJ7bKMPMKM6B6nWNQOasI
4duUkKZcuyh0+ZExT0k1ArUc8n7urDtsKRpiCxnCfK6Q35kDR4p3P2vPsfGf1Njs
eNP4MNvLofoUgrjFxb9Wpfdlgi3OZtRSyRsL3c6loC7hifD0D4ZFBqoZfprFhdOi
ttA1v5nFwioBA25lW9qOSH9zQJ+uNfLlIEmnWxDzeMklaNTK8N4w71Tarct8fbsc
t5n8L/St2wl7tL88UnkY71L1HXSIdoiA4Mm5vgtlGOjloyU8lYWzLK2mlZZppDqE
IPdMX2A3ZYGzKLsZ85JqPQLk19K912LRAnTkOrqtFZ8EaJgD5pdTkj+MvSItTmXg
NWYWtojRb2IGAaflpmf3azCwalx3q2YTKi7YfkCmVbwEvD1VNLp8QsmRe/IjI83R
CGHcXA75FqNuyLrvcbI7icaKD13cbHqShIh4Rh6mNyYzxS3WhKiQERHrT2y4mbwz
JG4uHNLtVnsoaOvJSoA/ou9oXTv6R9kXNqdX8LPYZ9JqzLxNfr5mXzCKD0m4pz9O
crjM5stjfTENq1yIknAzj1hIoKZ7/I0QL3PCwSszNSAOkxPus/D2OKbkCMHvG3X4
2xd4aO0RG7M6n37a7yGjsvpLbF9WAWxpR1PNvh9bycqIMOmpGzajp0VRZiJxerJ+
0HQwH1y2Q9aBMk+MGQxuKU5VTQP52JOD3a6kSeofWrLnuuHrTZjCXKCWHYu739ux
T/HZd5F+A3xHzKDpm/AmjFfwIu11koGzvtVZXIO6pT/e7MV41F2ceKF21bqrX2fZ
s1c1agial6Nq7+D6IweaA+1RdArRukSo7IUJAwQSiPp0qTrv4WXOMTqn/D4poXHT
1j34PeKJ3QVSHEvgMLDCZmp1DakS40uVfwSBY2CzpmPcpNko/zBhwwgH6Zj6o27x
i8WX13T2/ShEwOUMexWZ0sDjQLZ10rlf/ZrwofS0YVoFknDXXu9F5wc/iB5t0OCz
vc9SUz5I5Rln1/lEo4Xvxmu1uKX3HSjSwUATZyRCKfCVRYf2vOMQHvPFTc5uRUTL
Sqezwlc3FBX/N1uee3c+1UznGR6bhUswGdtTEpUnUXaAQE3KuvfdgcE2NCzcmmI5
phY/u7iVEOfTKeBKxZg/uTUttNeQs2kG9Ou0EKFcqMm55KQuv/A5WaVD2iU7bluC
n/+7QQQP4h9woO1Guj0I6UQSy/zsQSLzuN1D6PJuMs7nSFLclMaPUQ6esx+Sbn3P
mDhT+mrmFOrb7EVoECdmA2C+amShe2Q4nugUHCzXSynYJx2apOeL7KqJlO2SsT7T
MxmLBQDzUBZix3gis79LXLRW/Le9g4/1BjoYY+yLuLEAjd7XmvsO6pD6NdLrIGFP
RVJ8UWbZZYNGCHeNqLcka0nacqwWWf+YfSfZ2M0RXJuMrskOI6Zh7oJoZNDl+1+T
YGsDDu2iV9Djq1Wgekw9/yHx3hbmk3EVnrhbUA/X+CUxGZNfspOUNYhW8YQceScc
3ewsEwn3880ufNm0upDrnj3LsABAY+ws71eHnK/Euy1AudzIozfdP+QRVSb72uc6
HUTyrJPrSukwMrofABfedwTd3JzCeL+sj4Bvj+tJvrI85jkCyZGIk/lOkvPbLXQK
6v01IagC+IGFOuF3N1atOnXzEiGTN8JbOI1citXIuzJmyDgmubEXzRVhQHsGe4IE
KaYXPwrjokIAU/Acw5hsKlv5R7H5e8mvxq4a67uTgb1JpQUOk/bwGCnIqIg3KCD/
Gl+iiw+Ge2u3kUK8o4DbM4FnWrg2HrZ2z2mbIgSUCRsurWVajLZYqRvZLiV0k6qo
nraIr0/k/UpmVgvvn6rC9+WWB7FUtFT0OyAyRCGGu1YKvIlNffGIaBNURoD7Nmco
XOMrOa6iQCh3VUeoffUPzc5ZPwDhVvD21rzlPtu1nTkZjA8G/Xp6HTmNjdhxw9CF
cDwjRyRrZawDGt3SRRkUmKC1BtYP/QIn67ajgoL43lTCFOZrDNVD8BaYr6CFueUE
M3mLDy7jo+WU7tFaYGqnkOHXCzHnxoMhytUCLcM1fiPVxqkMkW9C6et7KYTAdFUW
rZzK/HxiLCeEjoKhRR8KZpfSQIO7HpJXeNio8K4SAIMvI9ZUYHadbJjmSkHoL0Bm
hgxUGW8szGpdml24nQSl5QJt9Yg8v8gQfdd/YuGURtt6GBJINomlywK4ZugOmfpQ
9PnPeodaVskB+FZR8eeLEFXIxkOrWO0RRd36vsVmgJRmwH608JXQMsNt0swpxBWH
1eD6mlSv3ovpFtj1SPfsyIDvIKku4sbDoRGBTtiHxpn6ZVHi6Xt/97aNS8IzLnWV
IxC3GDa8dlWVUQywDu1hllxSNNN28aTcXBE82WMXG1Z/ooJd4OpFrsfZhnbsZtW6
bKVyIkYNvCpXiQGJyva+I1PTK0QWo8A9fTh3X3Zgdd+Ukl1oGvNKPY1nANMu/9AK
VJVho4MgEaCHNn0AUoS/5gouqAxH7y8ATwCYqmdNbA2P0S1nYEfUZ/S2BtqV484J
UFw6IJlxSMyGfs5nXo3SjCoSpBr/5dhdQ+3RIf8isdRuLOWiLWqytuOceV9Yc1So
Ln/T7o6HbClmRIn1gTv8fhOf5uLGpoltEeJBAr9sNl+qCE/44CQH29Rbch+YPoU6
tCjNrztNoH0ex4Ko3cWr3pBcJOaB+z97KXBTz4fIivo1RsIrbTNS2B8uKjEagdUc
Pg9ifVuUBomiEKwVp9V/2HnuCqTb5xMMBm4UoQ4wIkv46B8xnfsshykjNOwAE0zA
PTX0THix/J0w2BwpNm9MNBHSjZKvvXxBPVucvUb47JYtoRUJauzC1v0NLHuj5/6N
h1dIsh6Jav/+6YW5f+VxIg1oXloB5mHrr49QVgQ7TgrgaBNt7UKqT+5GVjeUZu0g
q69CbhBIUOqR+t6e6/ARmyrmckUL04wLoHK4ewcMMPZiSBaJWrVkVsvGMkvGCTfW
8a35PB4+WcaBsnUeHIB8hW+QUwm9zGFj+Z/PlLbxeFHkoE82QZ78G7FYWZjGv0cA
joNeTUfItUqcrAHMuiluK35wAEywgU7Hyb3WJaTQEIDSh/TBNwgufkfenU0nagJL
NKKINVqH4o7DmTQg1IAl5yqodT64m2NCrj9wv4m/NsbsFGYGY3SNz0THHVdNpP8u
nUd+vQdFRg7r0MzDwtdNMfBawkjaQFmdMr6p1vGmzDC5qu4SjIIwEtvJKVtkULQK
VpRtOn+RobKt3mvzBKejPXfzrCAVtJsIVC7MapSO2fD3HRHHqq1WeGDzPowSdT2p
xx8A0ak5AEI+ZeQlPzWyOZ0xeJS9yYPTFncK4YjGh8h/gT8cG5oGevyh93BHIXSK
an4m+0F/I128DtfM3BoDcPr+BbPUaTMAlumJn2iVCxNgfVyUkpQSzMozC4/YP2I9
aY5ZO3swwu9dtfptGW25XS9JAL6777/z5UfLPccAfB4ZQIx6koMDu+1s/yEgmpBx
gxNmj9ErVne4guaxxGZcWbeI8U0MPPq2pQOxW/SJybYUrv+giQHkJS4OxG2xkr5s
0auGxBE5HhlL05GaDS4iRlukAlteFPejMxw7RGPLeu4uyS5udFcQkACcHRO5i/id
H/F/bgd8hTrwGyonitXv9jGT/f103ezRbt0YL9BsCw6z3c9zn0OGH6l2SRV7eebH
CSPAExR0N31tYnCx0DLwilIh5qA6mZs6pDAnUxrwArRP829UVBmLik0whe4unRlO
E7Mtd+dHxwIFUfr0kLtJ6+G/fsIbZTZhJJv3PgbICM8MgAQcAQy1kGzHhfJF+kVJ
zPYH8WVZ/N/en1ZU6AYXn0W32GQuEBr5VxT+DmwFK48PZGX13WFpKuegc9F3dvZT
Xc/2UdIHUYuOqfEQ05EhEv14+P72QaHXX6DxW7+dEMcbFWRHhdJi0t620qtfFGSa
5XYV7Luyff8IQtkz9PQD1Vrs1xkYgJQpRFRrRfdPiGHKiQf1ACq+eIIYydqaMkjK
bIFQA9FSUx+YqOvMaNMIjOUC5Gk7ToX+73ev1VqMXzS49fQdc8xR3DBl5r5uyZ8O
OaQnH/vjoju4BfPelDDNDpvJvXx8lRmdIPp5XIc0ZcpaZObFWhuMWRtQr75PWyrc
pxz7uG50Z0ysb3dL660NN1mXSXxJ60QnuCZvQPSmHeYEuIeRCbxmO5pVzjCIkh8F
t2mRCF0husuL/YXIgW/IqleCxQ80YF4axUOKhinikyZo3mvFj7Xi2Q/KaK0158ty
3GYLlXZ4qmEX7HH/7gPVCQKrDqzWGyKMLIyFGEO7tMPEyhZlnM/M5OV2lU1hb7Mv
K+t9/LXbXRwgDnPsTiCiuZCz75oh9Q+NvRBgV91tkoVFlEqtTYFOZ5EPJBuFoVm8
CmSsg+XE3Yvi7pS6S+2NZuEnIxFxYkv/oxJsRwSi4YTVeEqSDmPrwplZ/5F6bHzv
epvek2yU21qUF66YfGcCpvLq5RZb8C/YloeXewbVmd3MpIKL9wiLcoEyGwZ3EEUA
z/BpwtXeCAz+rqxb+2Yi3Zx+Ww0x9I8h9mQhxvCNj4bon9zOEOxAgVxzmN8w39rw
tt+lasV9Tc5loHGXySefrnmyuFjkhCI9r79y+D3a1DohmRoMAfEemnBALqEqnWUB
dLb6+2bJdIA8fq3mM2ngJC/VLtFL5lw/4txCwyiqdEZqoeyhtkgBOFU11l7b8axw
phTTOC+teyAvZ+iWkmjDUM8NLH1B3NkIUMNJD5IbYfD0L2mSKh1BZjxeGMij560Y
ayr0n5iwnUIzeWSA4YiXnmL+RH2+bEWNhgsBi7Kau79iFisF1CmKL76xNJ1hwCKd
QQ2iIjdKmvgO++qxo1QtHYXsbP2IJLrcBy8jny/56+YDeCJF8tnnNCzSdqhIAMh5
40mnFtWx4rC5LM1WwrDlvXm46RaEPhPguIGVJ1RgL7BDVWguBa8cOvASAI/iwcuz
M27DUXkL4aIpJeB/55QWIvxpmFAr+7g1g6GJPV2gMEwQHJZ6VPAOBYBUAHQQnkuf
aJQeJZZiQko7+pmedGgJ3X2eFke//2RU50ZcRCzDWIQgLz96VPaeExtX80aflabJ
w4m5l91fJoh0y8gAxkwiFXlocuMm8VFbTPm2Cnag64tlFhZWh0UkU7btwnVtNXqX
Nhgh+pNpwOL1ZDiLS/q+XuYbO+Slwje81QdQCACEBjv1wMYVRvLB+k7Fj84OZxG9
foWSZex0iv4XTdAEIX7Z+tBSsaEao4dwgI84JdCLMH3RTzCR+F7C2UT1xJiCBecP
26pUDdwyZ4Ivev1CDkvFryZXUPf8t7nX6BULlgUWYrirHjZaWnM8/dtWMWfO2p5s
OpqnrnqtZA6jliIpJSUZ1+T+xwH5G5K45K0s/ZEqb+i9sQJ/DuzK+WhvbvWVYeWY
zXLK/YnFRgmZlSfNUlUpZYlNU3xZunLCPjmaEJHGkTxZtutLeaU7reMVLcZPZbq4
tX4sALrMDvp+3OyfF9iEzY/eOWWHEy8BnHx+kPRMwIQ9oLAlNuepwvDtynidEYc6
Qj47XKai+x1m6C+jsKJRDfwrfwKlFLbI6/VuBuBrOr3aARFroUojAipBI51aYuD+
IaGt8AgeyJhNCTMyncJNIifFt4lpLUXEfPC88kiLEXKdmD1Le1ZqjrLVYAay66lb
zF5h6C3GFqe9z1rSNRLIni2UZ1jh00L5nLUXTqCHT4y3IONIGY9m2V00A7vtJ9hR
DRKrglPKo42mA0NiWcM62tvjGc81bGKFfn/KWyMuoqCRGzRKvA0pfgyi41835w3R
DEepAfZ+HEk2Fi6JVzfW6Gn4yNcfwlbJQ0X9yfYucJ9cS9ZRRmsojpQHlulFO6tK
cTKVTNGwWhluoUY4mVJjyGL1Fz1uM7s1JnW7BbvawISO0qFxWFw5EQJpDp+kU17a
3PuhFOCJbKZoIVlTGJcPGPTT02/lsfyRQnKmMxssKdnFE1e22pb6lLE1fXFbDfEE
816n90wVw1oywbIXfhRIvtmzaJy3X2O/CdM+sDX587FM8rUVh8/pWLqQETTfqHTU
bOP7YlW2nd5CMINfdGeOtxVrO7LVs5X1nhZMhwZD4ae0t5c4zv6bYwzLyCAFouQC
4yiizUbgFT354fkapPEHV3EC+k8sXj9loH/IEzYsfDGdhyoMmINwVQhKk5EssXZW
P3DLcDsrNp1nnVkdOAKgKgX3pKRQv6y2N9Lng7NE6D1CYZdJeS1MgWe05z4Hkz6l
N0yVtnvEmIIYO0ANJA/0WS43HOw1z+Jl6PrHyw52Y8ow8QWmwRsGTwfySCCApUAg
+ZZQeOvt+IjRCsXfLTkYO3VaViqhLxlUDWcRpoOak4YN/Q7SB/+cWuI84w4MvV58
pfvTLi7Ky4wNsCx+KROI2YgmfMf2K+Epj+INMmXGR/2UcG28sKfNoJ/Hv/Rc65vh
1/UGefiwlW+tenQ1syKMnfNZ7tAE7rCx0vPe9aQeCZuyJ/dFFKBcr93BqoPSYin4
78DfaavQGYNr8CRfrAAq7l86W6AUh3pfzLWUpYuL0tf3RpW2T1nkj/nYLhzPYW73
gsrvUTM7oG7sZ07fDHE4VvBW0/NHG3LU/fQnNSaiOMASudTOK54VkNY6l1EpVJ4O
E747ya5el+kqwELhtCd1NYk5yPwF5251Ayv67YsscijHrB7kamhnkcL9eAhoBHrs
OsBHqYGPfZ1dZ10Z1qILY+j/5sadceZmPTojcxYolEFuUQGGBuPGBOtbQyEHooKn
Mrp5umJGlk/Jm75i//LFoYa7quh1DEDVhgWowN0bVPbnbe7gyTxk+2qGWLuLGrYK
vaoKvlE2dH6EvvFNpxlxnwlBoLmdiXga4fNx7XYxWAd9y/zx90sSmobkM7sT9dXl
74CvcY533gyDJvAbe7qGvDJ2iRtVpVCyCPE1KSWSwy0PE177vJ4sKIqgT6gugR7c
TIUVFulCbYULCw+QaskvsGez6xqSN/ASwiYNuycvt4uD/kLszPMeg/Pk4eL3V5iC
aG6bX3EBA5YtLRIIAgxeNrgJPTTWkYdco5drFP3L6PArWIcXWw/EGu3mIaocOze4
9c4YvPq1CgFpjoaVGeh0Pbbzg0tsMnHR2Uu67rD4EO1SmLbmyvkdWpcZsmuXqbtn
rpoI5BTYJvqx3snQRLn6X+V9rmp7hlREkQKMwNNAod2WH8MgL+53zP8vMP3W9vNK
6nbPAkPMf4Zp1nEsyuTat1LMzjCkwrcps/waUawR2AuT/x27xgrgthTkNS19OdK8
KI1PlGAQQJMUDWOASAOwCdLmAO2/jYGWZ8H088E3t7vCJ8m6aJtBIsFZtlFreAnm
0kVSg/544YhmV6nQOw3dNRaDn2UqCDuTbM5ADgkJ/Afm8086xsfcPfaS01qnts+0
nKAlTpeNms8x03KZ0QL4w7ek+4D44WADIKydJJcZKaQnhaPvk4tiU0eMspLyqqX6
goyAMyLAet/rW+BfaraZHxRtDT/41uKf/JZjalDwx3sMXcHRuXTYKIBZmeCMrbky
Tyo1NNiR+MidKmZv4vVVXrvptI7zBH+uOoBzD7Lez4cu4dHDi8D92GOU14epEcyB
Xd4EiuSrq3HWMShcAdUs7kWN3ZuROpfMKpBwPHutBTHN+mJabPOJHSkfOtCa+gtO
a4yL1VOd2lFQxqJuxS6PtAoDqE5Bvr/AfiP7PyRvAO/5t/68Zx7huWDbOybjTx4s
mULdWmYV7DEDYIbL93jtneYrqMrWvMvOsgfU6XASXn3aXyrC7oHs6JG/dqht/kPH
Gfc7SzOz6XDBfLWpWZKOp2viBfzzky5YxIE7OCOslYIsV58aF1ZKHyeBz7s+u+FK
OFXUJKDFfljPWiZqRSK/mAm0TMbbpUZFJBUEUfIS9ifqZoBCgg32FHQIkqTlYlr+
Rk/6U6QBbDO+3rUFyeQ6K1s7gMWF7azj1KmOtvGGIFtFBwgN9wk7XTcCBsH4DlIW
qIISL5+w7K8ouOqn8Dv113zfqRcfo+5/bJtsjgVmwugUgDDNUZiXqjlrlV5P2zvs
mj15SR80NPJU5Hl+xHEKOXITJWJb5cqNbLarKwNlX+oU1DQEecLmLE/GzHgtMV/u
2pWqW7zVB65K38iVaM8dk6DuxkEFRLiVhA9tEBVxtpTd6hvBLvCGaBkoI+eKH+PT
XCtoU7pjzWuhBOryWPDIEsQYgbkm0z5QMDPIXR17XWQZAlamMS4GCQZQjigRlEur
RtgIQtucWd8mfvCdILhT/6lleF/OFMSY+Oo5v3lvv/89wSWU+oict37v4xxfzzwS
W1GUQmVmoveIE4nOX45k7hdiTRjVEJ+shExOUMLWDoqYaA5Ltu7EX0XrdmAmSkOz
yD5ZwPtUVHv8E/5kb/EPQiblL3LpRDUgb8RU7vz2NK61dK41kVGLqzGGlsNtSneD
a3JCAPMFrO4UVFmaRpUKyGTa4/a51WUDwcdqSE2Hy92WtkxQgTbWqZFuy6i9aSSL
07XeD0AMsw5ygBT1bzgvS9SHW47oHLxFn+IH3Pg6ltK4RmswOqykiAqMMLybKaG4
bFAWMwlOvJ99ug31bVtx8UjTOHRaXtFBWDfsQp4wONfbxQBwaJjlLJniel+K/Mlp
B6HLQZT0eW41MD5PN1daJwewJ71ItNFh2v3cEG5bLGCZFTE5hJKdzlvZyIu0Wt2p
1mj+KkgR0hEfZc1qEGDqhIdVeOEaSWNWCguV+f4PyMgPvdXOTwWN+GNhGcN8KBtb
WwGWh1KYAVUVZIEfyd2OOg7c6ICvMD8m1H1yCsWii5hd2cOXbZoFUXU+sNpVkE3Q
FlKiFP70nFO+gKafXqTZmgQSruq8Tt/nFQ/dEgInd80Lv/foWbriYgFPnizAmPw2
lw54BU+5Wa7fiwM5eGa/b3LkRCTxseZTBq+f4zuK9arIaQPGTWFt4TFWM56rvzBI
qF6ZWurSaGS9zMJvqY3GD8wGaQqUJGofNmCllAIAkspdYLcM7C3uwVs6fuD/jVRm
KZ09K6h/ECUUpnD6tL1XOq8kefDzMmrK5ukIb4L3TUZANLyq/Ca91TKA+VFcqARY
jhWV//QQDAn8OUaw2IU64fxY3hTWZLqJbS+iQeFjIPC1Kkw/e3QYDZTkey0NK41b
S+xmq86pfqYGSvx0exFNJldQkdpzWGnlEgWTRAXVu//Fopzl1vw1TQI3YkoVKOAj
UbHooeMAqVNT1GCfNmH3az5FF3IOvnqq82xSltYpeG6IYmECJUenTpYfrgSh9JQO
8g5DS+JO3qkPbdmqkPguMCDrhkmP3poQlfUJ6ARmvVIUjnt1xX0qo+WwedbYSDHY
L08GHSZY56axgbHnCmFSrJDU2zEB427dixMK1w+2mD9RCoGB8kbP4K7eMceyKpgn
ivgQz4bSi3YPAhnoOdghpBrR8NADgbuAxkS+L9aHTjany7vwGEjIH54DxVjsdq/+
kCt+X4cocugUFKjFw0LP3HR2ps71dER/61lPcXAfNxyAKKg3K2QdCzXCciZAa07H
8u2ygbh5tpqxLgKvt2lSKUXw5rexf3Oslt2gbgIiJs9C6DAZf87yY7m7fXTFee5D
KibrPIQFBf9tJ1/xy6nYkEkJ0KV4+i5W+jVGauy7+ZgKuFYzbKSSQAMi+9evf/TY
RL9ds44MHtLtoM+mUygEYDEXVjEjITotrJmOL1UPtn4UvJxz0cyYQwg0KUhYWUKS
lIrr2bKbtdl4jXeECDDtAw9320sq610Dvj8AQhhfoJkDHGSgELOtO04XYuR1s+ga
37ZLpq25LeedClt6yjIXqsI+CfEhS2IUgVkGkr+6cckOub22SxVN1OtDfTPqnDZp
PPw+ZqFY7OCoUrvCqtssiaXsrq0ad2GnrQSCQnNt3JkwNKOAPU+OD9DetLhRReND
d5s53Kzzz49VVOO5hR2Y9XWTJ+kqJD/1ekWipAhT+oRO1rkpp33iUl6lUauml+1o
BBmoeAGB6/Mpmih2s7lH/+cJNLRdKmMwxw3WdMWDRl3bXSkaKlNXJlp8TH/kGL44
NtKqGfFsy4mVIDtJEowRxm14KhQ3PvC3ugKSSvql0f+/XvBTMlhtBsXEE0HwvIDO
gMTeG10V3jlYx0TKAry0iU04gXigfDw5JmCbO3HIrJWOEFsoVcQm1hrMP1IfLugw
spfDzBwhYRgCr/INM6bQWJ9LVGmbXhZP9WTc5tRkQdE1PIDcFuYsQUrPchH8WBWr
i9KLBlOyIniiYu4a/H6Z79L5QnK1SSJMvkUwKUCXZf4ONZpPhnQ+DOkzbacS37b8
81KD1tnHP5RN6Lqow2SyBvd/zVTiwd12sTfF/deTLc8A6a6T+e+gtOWFVniHgxRd
/BpwbmvjEOk2Vi1geJURViwKlhUhCc+CbFv/c8pE/srpF+YDNX5xmNDJHlnJBNvk
tQSpihwzBBrmqq+RV6qRy/fOJWLTaeZ0yG9Oo+T4nq5lrvdZ4cb9bJg142GFmYvr
VP2S3AX02ZMvDDDakFnKibefufP4aOwVcnisOpVuqpS3RU97dl0ko1gAVGFDG00k
W+IGlOO8XC5PUL9PKMEHVHvr4nAfoQ3EBSgiW0/7nrHag/HBJkx7oG1xHbIysxRg
MUGDcfP+SEzuznaf/WOCEP48JbKl5QGob+k4jP1nnZVJ1LvCTrZ4yZbvcFpc/bIR
xnqGcxKmI4KW6D4zCSSUHRaFLBNPCN3ZF53vSFlAxdMv82WcP0dNktxEu6/KnBJF
Du3iYXuKKJaEIV/S9fQTPrfhHSp1ubpXc8s+Y+3z1rH2/CtxZvxWH8Ep48qv8EvZ
pfYuSrtvUc3OpsZqohX9jiNzYAHFR9XDUh2O+7ZpwCKhbZspvMMAGTLUKIsh0f/g
9hYbdTRVxUOS+0PrfPRSfX++Y5TOC9w1zEOU6gqFTElg4UrLRIL7x3ePJSa3NSB3
LR5GHiMdgF93yEFyDZmljZBenoDF2z1war7mMpfrtKhxPh9gUtqn0q3A+TsFZNBO
+ecQhZ17Xcd8d+bhTHohlc3FVOJujAfPocq6kMSLXg+ZsJdOL7QDUYvziW1xzljd
x+0YTkQhTB/OwuL83+SdPOj/nUK6YdFQe+OyGAQGB4LB2xUUx+rtCcjXo3VQKEIU
ed+aPJcu+82scBbpvBH3nul1IELYtZuSlZy7GYFApu/QwBtqG6F6Y4RoVSn5uHgL
pr1Z8yTJilokRMfRmJoTQySLsL0TBnUb1Cnl9wJxqniSMfCDWrg7N54HVaLO2dPB
Rh6VGGxUf5nEAazw9uIFSfFlZTDcjORKMUAnz41yoP3b8BMjU2r+22AjL/vcTBBN
mRR6SAeKvXwEhDv0jrcnOO9Nec3X5ggMC8GaQ3wltCziugjdP5K7gXv3PU1nTk/Q
NZ4sEfoL5w2lix/KVR/hTIrFaghH5h2Sipy+0PNzPOmrKKaNpVIaeBD9Jrwz6+7q
PFlhyTwwcOs1xSKFPFfQBQfZ6j96MSOt5Kc1V2pUH0zjveNPOUvYPKDhRvwv4JnJ
aoMWJln9MwZyIx8e9OhHVWKhJ4HOHtFB8rD0zNA1MPNOc3m/YEWX7mQ4ue2sdCCK
DNbZfLou+1SX81RZ3kphcGZT1VJWraqjVdt2vnvBJNr4/KUE0VY47SUSteCs5crL
hCvS1iw+cR7aWX6pu1XegDcg2dsfea1qcRoEuX+bsS2xECiysQ3+5TcCH/30fZha
myI91r/rEFu4ux/fZR4ytSp+md+y5ec4VGWVTraYoZS4QIuKceaMNAp+SZVVjh+4
msse7oQ16FPPpVCgyvZjW06lTYCFGanNtESs9Q6mvef0zb7evLBGkANEiiEG0qdK
IfySaFuwBJ/W0q32BMzJsJqia4DbA0M0Zd9+xDHLO2Y99Sy+/b74ULxCf6fayF2G
RhbGKdhrgN2KhigWvsD+bx3M5Om61S/R6msfekZsAuoc9Wioasy6CHvR51Go7Ra/
i7M3sOpCaU5ChINqgryTlZ2E9Ze5KKP8DbvicZRFxhefUvwdMEhTOhDZzww19lWH
O8ek6jQbN9OvTE6g/IdAPRAEvao8XSlKEXbHybx/NqeaX09WOcrWz7Ayla3J30rU
NkMoc8hcIHXEr5SqC/Vp/33KSZZtXjUT40upPk/EgQCBYqiXKGfblCslJ2sSqc7O
SdgghfYqXMewhywA/cNd9USWIWJAFZ9WidZoP58CNFRLW0GgugjNO4L1y/Ie7fOQ
E93UAEtECnVUfmDpVTYKHhcfyvjjr+8V+MJBAkzxQk2rAeMUEt9XmGRLrexbWT0a
M0usEECXMk52/gBmivML7wQWiHHZLZAV2Il6z5JQd9xlI18dy3QBgDdgagCDqOde
kQQh3b6XMKKxvg6nWo5xQmxCQCSH+sxrdyr7PmszasEJmLd9ndCiM91+ciuUgSCM
kYfH0p/blCCLR1b7Qnx+9bXvBrU3g7wDQCL9UiTZcwRMQssBaJaONL8PBSiWChwi
YMe9th2+uKqkRlA8oXn/kn7ODyc0JYFeMCYfdnD8WEdsR5ycbkgHFYMAdcVxAuYb
Ry8OFw4Mg4bbrVr86O6JHPHg6PZItoienQITnX4Q2irs/76haadSIGBwSXrM910c
1yAHwhC/CWZdmDrxjweFmT3HyLBy4LhFRft2gUj0bt/SCaTQ3CEvwRnJm1UthYjM
Vslo2j9l1bqTV6RNEZkAbZUdYH4jolXw6PhSHn8E+YC5f9e8yMP4Dfx4rMvvU70n
qdMgjenkXnQag64VVXmawFtPOzNlMfcqPxGq7HsAMe+3h1JXeb+5OkvMN4Hicgq3
AWHP6k0jAgxqwSGnVwH6BwqMYXGQdc3bbSZUa9/aMKtaKdJ7810Tv0M3MgVnOucH
H2vEHhiilgwdPqfvZWqK4DTCNo1dKBnNy8Ue1cAXVmxQlGbTNxzPPi4mtw0iP1SC
TvJB7V4FECfWXt3jVJk9Vvw3AW4n3qOcTJ5atF+HanfBvoUACRQ6TWKK4RTLbwMN
nnWncgt/tZlvjXqyz4X306dXTwK1VE2LbFC/9W8PQWLAlB2gIfsse1MXKAbFonwl
z0rDOqKXsqxCvnilbnkAoGDLFMdSCxASWRxVpKySURh7Pr3/uDgSsasTwFHFyMJg
96Klw0vVCi6+Rwr8Ul1PGYoFvcwAX/3SFYCU6WxSMbMYfJdNVgVj2Bjy47twz+hq
IIra8/r1vwl4ItVFRXJ7rjiarIpq58snVDhqKUTqDWpERf5Gr7Vt4GHdal+iBeJY
e0s4LF58TscCLh7YN1euSuCCfeuvASD2kL6ntFxNW0C/uwTaSFHSbGIzRd45e1ts
sAyzZ0J1YzPw9xmDGxdMM8O5opjvgb905M53JlMhWuUhIaOSt2Q6pggSBWqegGRU
a0fzHffWOIdi7RcQykaKK36px4ZSqvlhCu/3reENSCHEaiQtUUbu8Ao52DA7W0c+
103mJ3KsxPGW+2ZHCGilJYAfpfO537fv7IEPkel8ZSy2R3Qnxn7ybbhl/OPimbqc
f0W49WvGA0lqSfCf3J8Fae8iklu0Q5umrQHcKZ1fTJbCCTEbKxDbL3D5KpIXvVqn
FAK/PM2BI7VU1MvkJ9VFC/qbw6BhpZ8d06DuRUBcIj6enoReK7ccZ0P/4woPTIZ/
UWmYIkYRNRV9RlixwDTML6Kw7C+4qR8KHdO5Zb4snrKW1xUo06F2aphSoN9CxBZ4
PGHkrJWVQYfGt0A7IPcx76fHTwykeFptUnc+I3dAeyaR8/L7eL1Cjp5aqm55nw7h
/3Z9hZyzaIWZZbCHVreAlES0l1utq8V7NSfA0p/qQpVK+0lnr7cCjiV84KCvraoS
B9BJ8CNGp4ljMixsx0MttJZTSLrUoHZN2h488w5Ro8QJpH3cTtYxYAyIaMyo4dFX
8oEPalFqZkM2+xyn9FR+aWeaT+nyyPrMiC3EEjIYyksxK7BTSjOp0CbsnbLKumrz
zLTcPvK9agaE9vA4JiTuSkypoGJ4o5npo3Ryr34xo6q4nk7DH71U5tervl4HFBgP
Y3FT4m3ZiZ+H/ZSqV+Ft9XMi0KeWWP5Sd7ocorJ0GtFSGaCtIQIarGdF7umUZOcm
E5mE8sk9rChnWcK4gVqyOOIuIU2+QDDdywT8fLvu3bMMQWCTA5enDvarkDa15qkN
KaTJTYNqSPmq81qcfD5iSrTe8dYDoi838DYTfkdvRvqLjUFA3R3Z6JiuvkkuJzHn
U8v6VM0XZRiGYouP9JxaVMpb4nbGrmW8sNs4RHjJR3S/WoUQzKZT2gFYGnmHUvwL
INntZAZ7WcSxv2aTITbFrWluRLYkm7oCY/9Q6ihToGFD24UWH8bzZ0NX402LbMrw
8siZxZqTNzD3y89BOkwoDtMrzbPScJMNcQ5n5V+SbSAPnzjKX55clOyIQbV9LvDA
oeNE2lCu8p0WwuRJk32LjTGhxCG7Rn1W4Yn8hJbxn/iiRC1FJF0azJ49QGPPmQxF
Zz8CUlMsT9eMaiI8zHfcsMpA0QRsR7a2B3JMTj2fJsdkXJRxBpT5fajkO7bVtScE
SD2d0y/0E7BGT2OQCG4kBdB8WNyLUeMuNt0b8q8AzcQ0POw0pwoz2UrZO3sybxNq
NEdLMLGF/9O6+BOMs9UYq5WrnUAU0Ile5QrgzNnD9EYZF9n8S9Avyzbuj8Jxf+50
aK/jM0PQPjzIAlKylUKE3P1gM73eE1B6lZ7R5hgsUisFqF3gwCBhil6c8EdBIYux
8Vdxd27rDxJ+I2LQ4tFylQ0YQWmb8DsXgyQLU63fEcANjqDTc5IuiWuzDQvNQ6MI
cfA0WgCi+we8ZnpR1wzimj8CQC6l0TK0a8muj8/SOeS4rW6YJe9HvgK+/ohlYL+k
IWHKS9jEPfyfoeThwOqr5D9QocNDwKw7Li3Y0tXZv06r8pQZPvBId8nDRM87qbeG
iLOShmCAaha5CjwteWUurHHOL0qfItuoMQqlGaKOPozNoGYDyC8FD7bYClt9p1qj
b/F/qTRup5QJMaG81VDTtvrHLhXUqWtj4OUhVRTwb6zjagGXde8JQHa/exaWQEyh
cqQRTXOsrYWH2IMpyFJDQIQ93/lKZQwSiPLD1TTF9j6O9nW4wgCgYZXET5KIYbOU
09r4cXniUUmEKcSW9jrTD1p42ICvRGNMP3kyiiJQDdR7qeezxEp8ykdhy4owpNi0
pw+6hk+dkk0jyfFmNvnZyE/rIFSFjiHS8XPTbXDQyNv+vC7/Q3R5yBBwLl+malKG
2K2u5y+bwqy1AZH3RaPyhnRAk70cZgq73p40OE0295GMb+cyVwENLBuqFFL9woXo
FnuPCYSApl+tZ1M4u5sPTO65UeKe0/m9k2gB+rDndDr2vLphsFXAIiTdoOBYWFVx
hp3lUdy85IPWWjkwbE5NmA4bNxcPrfUehpdmPoyPm/PHvvPuDG7hplf/NpyCgzsq
/5C64tDykV7p9IRLjNz2BYFthbi3PJWeko1rwYNFzOosbFiWg167aW8pZZ5pQJb1
kiZ4J7r7O4WEhrtoetfqz1JmZ9UhrJvR4tRak/T8CwwBo3cBRqKGaapnhuO9FCu1
uRwgXfbHFnQQ8/3bQ6reU3r4FMkLTeYNgUysRzpz/DLwkAy/I1l4HOUDTbhyOADk
3AhU/mxlQ5TBZEyYM3TlyVNxjDU+di0t80HHCTe4fJiZxhKbEQDuoiZsvVsoDXPJ
ORoXpdZyoCBosVYJFsfgmi+r0ez4/7d3+7YRav0MUGCYe+l/HvZOu42UMNQIBUM9
A2XJANwjh5upd4i7Px10mW9VVLp/0s1uGXOAOcIJbEjLszksdBayA2ols4lUD/YK
Jym1aWpUPMv+AjFRSqIa5FWUsQTMa7zu0r1vHNTriFrxxcpTBasxnNJRKL500kPq
W97b51XXgoisIyRAMztd7jWa+fb402Jk/MHzscd5l1lCQMrWHoLxk5oprZM6hcpQ
r6vL1sfXdiP3agp6Qc5DNy8M+mnZbKwuUHEH4LTiQxsaw8nJGI8GG1fp765ji/8N
NMbCBP9F3RQHw3IrcjlwX5vm51vycam9bnMbEDkSHqVyjOM4PJXqfa9tK4po60ip
H98kuV3bQYLjbMBLecVxb8bpo9N8N5lcVVytWJyZSuUPgOERBoMmYyRy0W6YlYfH
Mh+GcBAwImN6vkjq/pJ1tm+7k/65hE1JxYG2ZEXo+IbRgaE/llp7aQbHg7jldE7q
g8Cencw21Qxg1P79w3ufMY5N2O2iOzfRed2HkcGwPdKnTbT6S8D0fOlFTiObErz/
9SBY0aQzGNNQLY4zy+4P0HF3hMKPTdvA4dwcniXZIhxs1rNcUIJkqY7H3M0q38rk
/LcDXxCvGyOA/PggR8wt0xxxUTNxzvfejTxwpDAr3PEgP7N+X+X5Wts+MuVG1fxq
7BQS/6eFlFpO5Xbl98Kpa93FHVAxv+0w57KMz0brc7RQUjTj20hU8uuxcx60p8cG
4+oYN98EfCPFfRbDCArIAPuQMZHVMrzZ2IO/wSjbaPevFP5nmHvTQo4kQSsa9FaT
t0yP28vY+TRgc7Vq8dE/MRPeFqxN5GRYraBkqoc13cBxeP0giVEpa3jCTL18HRpK
LjQHmJ3YSw71UVQXcfLRgVt534pJeDOmLgfPkhJd/feRFxfd7U5NuW5V4Mz3KXK8
Vn+23/BftXNI6OOaEfOxa4UfsxEcticOSpnehOLxV9H9cN/YBmC0C64xxCIpabuU
liK88yYJRgE8n1mGBUANP/33svT7gEUEJGPTNxJpEtzT6vAmZjBgkWmZwPCLRIFD
8TBQU9W8iD/86yeUH+lItkq5CKNRPIp9CCuNcIDm0gZGBa8VH3T38zxulR6Kukfh
BhIFaniPW1b+SjBI1jgg8c2l5qBFbC3SkroQyG2PoOF0iNTB1GwkwO1yP47uF/nz
SOKkCxcpC/Dfw4hnhE5E1qYtxRlvy69AylFcS2dT15gD4qrWNlxj3L2BlQegq0Rv
vgYoUFdBswmar6E10G9GU+PGCaxDRmh2I14nHTeMJalnHpA0ON0+DDDezxYWGdGm
MF0gj+h34HmBv2Z3smyphaTgN6CC1hb1yu+4fiIW8phUD8HVDHCHCFjHUIvLEecS
QpfcLyEeBS6nCyPOAcfccMKcd+ogsx/kxfwrYClcOhTX2pdkSwoZKrqj/Diext07
eFUE9mDp2W2Et9EJSOZ0J2Ezlozj27Cqdg/U6ttMqT1Oe35YeohegktWbRohWmL+
xzjGARs2iHykvuT046cbDFESepSv0HkkJLMLJXetZykBk3Tz8tvOuGeYZzHuZ7qh
kcMjNXF7f0C0mxpt7Z9OWBf5Qb1xe/C+h9CJDQKLEVCcBXke5kOqiRxMCzqECAsa
hHADmggQZ6gLr0Ai1koYtYANoZATjDbfR9jNWUXtsLrFtjHRTuzyfcwTvE3oyTuU
fWyETchYQZXx0zNxLLfVHZIq3/ThvpqYnpMEuaalTPRCnkHp3/AkWmS9MDlfbE6b
2sl6te/NCTu7Vj9QvxmoL2/Q/GncfkGF2M/Z0gz0ACRYusgJz+74mjvK79SwmmI5
xQFSxM1c+gGdD9Bn+meZXdktFoKubNPwoIco5ehVlPhsgv0HsbEO3s2CHf9d1p5l
Bx0J5bt4MaC2w4EP78iLlCzEjIXx+dZebcTH+F7NVX8ePphmgpwe61PME8lnSaOa
/nJ0ZhQ3UW+BETW2j/JrHU2rsBArqMg50iAnWQF/Urh/q9l6jOeVVxfEeKDR7/j/
qSTG5vNGPnO5ZkswqGI5naA2vD8ZppE1rxm5C2d2yZwWW07ewYbiOnL9s44ACBAD
lcEAcgTZJyIrnR5RhR+84LXKUVzn3gQyPTjVSAbmg5+eOF7DrDwE7BdwiKR1Mbwd
7Ju12h1hQ+yQ0ut/yeVZRR5zcbD6dc8rP+0n1nFgdQ7n5Tjg4/e6GRFqcMVL2RX2
X2CL2viAooRKbZDIAHmqp6cMQUqPXIj68YbBM0DtylRgCoWgLb5YC1AjZa5Jvifr
7EuE7R+ErBqKYQgCLa4Ai7Gm2vS5U+AAOK4yZUP8um0yHxSPwj/fxxg5PDQSG8rc
WY5iKe0CvQDYLM3aa69CtqaVchoZLC2PvFOGBMhMJBchf+0OdrrshE9C05wt132F
rVwcsDaQQhogWgfJtRvKk4gz9lZWMg/yxO+40pwtGFEYc7vg08j1W2ExWfvJCQVE
r2kU768s/ywtEFhuP83OovACyIUg3hVQIZ1mMPKemvDZj3EGEgFVEvSTkRPwULqQ
LpS/sU02/oFGupUtYeSEJf6hRjUoUxn1ncrbJNheJ2HzDkF5mDqSgY+K3wG6tBeG
BqHFq3h6Ku0lgq5Bg4EF8OnsEAxPsbpyFWYUvh1vzlCOqSF0qiUfcu7QqPZcEvwT
8f+5CGHQ+zVlsWMohECBjmUxwxZ32DOjCBYX5br/aIjXwkcNG6xgPzBpn+Uz0/TZ
W4kFzhOupnsup6e6vN1/uC1s+ZFIJNNQ/pitCw6P6EqEClZph0/xR5uYv+IpgJLy
NeblnuGNPbgq19zk9D1ZBvADUzrUlO7GcWdBpRmppjncXoY+NQluYwKAsXqYp4tv
b+gZCe/2IuHX96b6RYTyk90Ro75WDE0iB0tsoGp4J3O21QFwkPnyqXywWp3H+JaB
qjWj5de6bKkl4Ur/ulI8M1zBxLEh0j/UQ2lNafIZ6sn7EYoctWIvKFuS0DO9DJX2
jsZW8sFJfnJDJJF9pjOOcEzkQE8RkT5/CO34z/ShXmYwJRruetmexYRrDzwYJ8gA
XW4918DVct6Qbo/HSEz6tSkHXLThyWOM2NsY+gpnGyqJf6OjwEWcMJbvPZumL8ay
HAYfw1fANHN/toJ4yEmUf+zBddxsmlQk++/KMriherqQaYSPxZQmpAOAo7FFuFOa
9Z1K4oXUEfoEXWraNOJJl0HJXsN9Sa1etuUTSjAIXLunslCJDxkEWTY8NTdHH8Rj
1C/BdJprqLiHeRavvAlyaFMNKzUrVrYrLKjFWThh4B9fnqqovjJ0nX73Cso2pzfb
06ZYl8hM2pIRi7DsRKeQPGiTeTAvMOUQxt4lTdxNkmveflY/M6tAGtuZzqwE3Rze
Im6z+5z+3aqNqDPARmtjozro33L1M6PQmEGYrdvwBgp81yMOCcFckF0zeA/wqB7F
DhSbHeViWqe01c+Ge2G8zVVutdmMksFNOEWgHdoT5aG33io9IJ6yKHXR7E05cFek
7HepFskDcxVxMYFFyYvGP6KKTKOLXWKYopT/bSToapHu/ifXvPnq1mpYcOgN1G7R
RaRTLRhXSjQgCg8ObmvDKavBn4GrdTDbgLrTqPMklcQSqqQ9WRnNW5CH8W7EuxTE
Lb4mr02XvkR9m8xl1AP/atPxQZ2ZBlRT47mi1JvZkqHhBRtb/lxXbbt85hIGKQ7s
vWsIV1sXnvJtJ5gjlB/EudacMw56ZZi918EEyz5W06kQctQgxWYi+G/D5+++iKOQ
v8JmAEoo0BWzn6a27YomwTx9k0dcfqiSs4r930ndzonbkf5SonbyoUF88DY5iUKY
do5BHpOn8JyC71Qlbsc1sUh8Oo2HWkMvLoSFkLE4DrBTz/QS7TysmH/ifFkWihiL
h7oer0rSR06Diy5xauPbs2UDsBwRxSDcd/ZKD0NoVqRLmYccSBl87pXrXjznjSYQ
bQFqHgNaI0DKhqjzX1cVKPd0RkEDCj0wUN13HnAXzWZAWRazo0NFWOibHlWcDqFv
IEECcpAl2Km3NJg4JKDFEi1NOa28AJDQaxPRAqphWfL4cFY3dGo/sRIB3Nj+YInC
ZIACpkCeQlZigdoFwt9lV/xv1873BuDSCxfa15/wxlTX0HUd2A0rWtlVlLX57gVf
Zg4+mJXTiGP6ut3LSkGYCJ/gSZRnsQZdOMArvb2EHi+p55iboE979YfCIXE4FkmF
au3A8KOwha9JdmJMCrEQXdW9t0WZiaxk6g4/1BWPrW8f2WRoAF+Z8ZFxCYJKm7N4
rpRc1iIIHcA91V/OR1S/GB/tl/P60pfXhFyIXF1DCghd+Cp3UtdLx/7sZqwKwOYQ
QzcgEriBdDlGVpIyjMEXC494s7FgK2mPlWBIJeQdGGZZrVYMf5dg0/2ljFufpweC
2hD9f7NfvKLHckAQNULC92MpjkEwISrQTb4/DfTHhlR8QSzdEHBvHLqDilcKsphk
1tMFpd+zGvxDAjvZ+0iP8RBEW9iVlC0RkaO8xTCHF48C80M08STQnCTXwgoyg37u
GzAbNoJz+dcw4mSVI6d48xDGh7uXTBk/VIL3SPlafa3bUtvm00fHqctGv8Vi+Zjt
48vm+lpXhO8gEi+UbZrGRW8o68JpKgd4WmEbIkir2voONiUz0ImlcPqAFGWy1GUR
6XqQb8cmjKm2dz8BPUfNdwNQQrSecxU+nL4hHVr+zhYc3YtBvqK/agueMtMi7rQN
Wr086IOCLX9/YOoIUe0LFSNNZddJuCBPQ21jYMPrExiXcXyDwlIDWfViTqPnQkVR
St9wBmZSlIbj6xY6fbHbLRnVj4+324ReWDIiato5ob0yRV/sTWEDsm2VLWo3i2Wd
1f8qmKzvA2JDILNcu/LrO5d8AoG6WnBKa5IhPYkQGg0aaliUw91d/nOeNrKJuUbV
8/a8I+/0I6TUKpQRV78Ky8H+zp6iBWlokxTYhHANryTdNVEU5/x1BwNOIRfx0QUn
YL9f9WfmPbbAmL5fyGBevjwgD4GCXNXot+xgFKzkgpnR9Wxjo2nzkJdSXA5cEPJL
yWlL+uBGzEAHyQj1PG1tbpjW+JdzqyeynpFpOR/S5WUtrk/sI0dB98Mtvv3QTRLl
GbRkE7R2yHQXAnms0O/Cm+RZPk4rwv+6PLUgY4FKMty+y1vDKMNviwHAFxu/DzZJ
j6eDxb8Hg9LZx+tqqa4IyJGSmR5A5UOPFZKR8vqgsOnnKpMKHhN9ijgO4bvHgEEe
4rkgRJ6CPTWIkDpI4ZY0zvIgt9Z6g0rRQEaOBMHSlLMggWOs737gXMmEc28wwcbh
uEPwk2GOgjUBt57JBCfzrF/kuw4/GQ023aNRhikm5Y5oQlGUUiFiShEBARwYMhr1
AkzWqgzA7ACan/d0mUG2OXHLyQB6HmZfDWKMKakKSOMiU5QPVY1b9E+JECANxATW
vTF0+jPJZo8+bFn0DOjK09PchWucBz7g8vsTYmAbL8Cjpr9MzS9/1OrcHhG9MNys
vM0kWQdDav2z3XNEjPem3uSA7eoU/y7JUPq5Uw6VxLlO/JQqXY/Mb8SwbDQ26SIW
ccBC6fwrAAVSckRdw0XPrwFNxNr9+7xfwBppguB6DFNCcPcw7aL+Xb59ak//3glm
FGP39bmtt9b5ikxZMo8cVwVXK7KiQBJEd0kFrPVr/ptXh9hN2rlOrCNMRwWqzIO3
Zq1BLHnzOXVnzUKFbVuDCC7nO+nICwtUMbW8tEnMPbYkUBhMMk5VenY+eKBDZy+K
pz7ixIfhIQhz3l62NAOm2KG/+8TZUBEwJ0AMwsdlxgEcnsWtD3HzKoi7Ge2KkdIY
PdrXoIw8axYX0zy7ppWBuHEl3qbsoqjWj5UG21FYhGf2w/2MiQv9Ou67q8k0yiTH
4apNa6u/AgVkWjAZF2LZ286n5b/muyhPLRxF5D7OD/wOlRnRgsomQ8mO1iy9YqDM
oNTvxF81gDuRuHO8K6iQNNyUK0a+uTE8E0WMh4sZrVaGAck8aiBqvQ704z9RgQQP
PLl5EKArPoUOr/RMVVWSBXYpClSQ8Y67Nl+ojLgJIQ4njFThJ9sd8JOlDIZ6BwV9
4iK+2/ZObOUgette65i5Chet+h26MvXHi7Lrxq/5bFAKL0R+OovMhWoVlOZofS6V
J5fnYurzDkU/viM4/Azdcd3J4mdMuaB06rvHUBEwMoMeOnuSBwo0b7FDlZwQbAFg
QI9MkwJeilimiB6Unfi7gEiLcV+k0X3wvEn2udvFH2nVby5ZIjVshM7VebRm2GUb
M8eQM7wHQRORg2jwwTs4EYnaTfxNBE/o7zfjr9a0+CGbk+5XFHyVJw4NS1AeL69K
+GJzwK12uo3yxuCXxHMWODL3m1fz4XqrvGu2TcZlCAdFcNR/HScG3o0iVMhizwdM
PQ8nwhO0VGkEuoGtGshg8EW6Dpz2VIDuiUEW+jNH+vcaLuiQXI5op7D2k0ioi7zh
nmXEFIiBzTE4aysULxdgsVlILJv0JOfisJDkopWEB2FtqoCQdGcNgTGWM57BKGMv
9Bz+Rz8QxPpq7Nw4ToYF+z4kqSOrENaVjiLmdlPTvBt1fWRNtD9O9VPhTtnNbRlD
ZeVcuVhUH9Z8Rtgt5sAl/ZCcyOxO3dho2ZZiL50J1s9zSzBEWM/3ObZD7Li9f7Vy
p4HKuFiI5mNx7HWA33sSJJ4ioUvT7NmWhjD43I8KwN7O8CaoBYdPw4QlKx1avJWQ
Sg+/jbiACc3KYqL1NRqzzxr1NXJDiIKOAgyxWAi1e/R2xFBNDvO4nDfIFxYB/wDS
QLL8a9P76/2GxUzRBSO/D8R+QVkQIBrVslD4w15Mhcx0Wv0IwuRYujgJ90baJzt2
2tyhId4lv1asGeVjKJcF8sHE+x6yle8zHQvkRuJiZqw0r6Ib4DZ/t9t1d/6K11rG
Q/HGAdMpM7KkuJyJfnJeDxaxCKMZfp5KZ7V9eezvhsFTnEpWj3haEMbhYHqaQdKd
bH6WtOD79urr3SwOdQNNfXhws4YfuTZlMfrD3Ec622XQwv0pBTQPmecKRdmde5dQ
LSOgQY5E1CRzUOf++uPla/JUdeMKscuvPQmrbIWKnn5sAwxPIy9kvS/c7dKzimAJ
6oUmXUbKFWtM8UEgkMEU5rtf856UKXO1CY3vX22pcud8IEjSD37w3j6oxsZKwEGA
mjQLPEG3Q0F+bk7Chwf4AuDhg+bf9cy37LbKejvO5A4VX07dRpgaEU70OA3uGXFy
Lg5H10y32wo3J4aDUDh29V+GUwM5Hbipf8XtQo5uhfKROS8XYJ4jvNVqIi4utVoN
b4y0cDwmsKZhhpA8OBoarVRljjA9iQWMEC/QiY9S0A7s/pOlG8eoIEcf8K6MOV69
vwaAW+k4Ryz1/O3BRzE3VFezLQIeD/AZc1waw6QSop1Tpnvf9UEAeTu+KrURF7x0
AoOQUzr7blx+ADq9lMOdSDpK/ZRKfOAPCCAV8t7FJA553/HqrrClwhUY8jFm5UZl
pybvf8YdP1sZTE1Ewy5n54rLq+dOKKOKvR0O7d7rZdDlwo4sbIoioKIhZP22dNQy
FN4SJEoMzg0nTgjSK9Qkc9LHzuNS54OYtMW90VKIN2Lz6mdoCC5kCBgU7kv3ITgR
6ds0ep8LkcEpqckUoQ5AS1kGGN69mAcRTJPkvQRn+i9mFIle8agaTggg9mtahsRp
ssbAmHNqdVnxjN3VqtWrwH/nt10i27VtCOZKenzikjVGjAxrhrhZz7oq6u9NzXNk
UgK41pBYy8yYsNzr+lI1DmabzOY0avn0b1Oa10e3jcK7eHE5603HHvLqc1Q6riLF
bFsZq8TNGPxEMqR5d7ZwYpAgR82OTybicdLfMrK4VTElGSxSvLw6j42xqImM14tl
dccF1pBlP0mHq7BSNqIxWIR/ICWXOKl42egdteqcqbpvJvTNlnnQ5Amd1CakHX0s
K1xWgf2/1wi5uBreGfIfgXrTgYApuLosQ9KjQKlZnkMUnuVVh1MbeyJ61PmmXnyV
2ztOYUZdrRVauBcNCJWI7sPXh+X74l2E7+1aGUVHwsWLiAcR7lNiBINWIsv5m2YV
DRbCghlIip/cFyzGCbme+k5F7IEaDJJmwcyHtaj1gwcd2cznMMJm0Cdi1LhGrlXo
QE72w6JcZI0oTTJ0+x0k6JjsnG6SIvCsP+yyR1/CzU26ScJNIpN53+8DTrbw5w2A
qcwWjPKMeFQE/wJmrhjR0R7K0eS1I303yuEKaNNfRxXdupEs5B/gc/r55F0B+fUF
RtG5pIX+Jzi+bJApkrqBKeXhQHxd4qXPdvFxV5Z8t06+HOUYtyxHgvgvhmbsvT1T
AzAi0Yc5pIK99hWmAROX6lByGQuAHAkTiaLI7I9QkOKDdPXtyyCtyan0haDR13ZH
2imNFQlQlSQqQBVIDeGt0EvfRljZfKlXCSeQhoUe7WTy68ujRAG8Xa3nqtAVcRVF
xKZuAwPc3RDYzAuCNYBP0GbIF8IyxVrGwPNbFTjA60Q/++b8EUrdytOFKtkPiy69
n3LTs4mcVnnfVYvp37uvEjCACnYZozqlWeGFJXwseXWndMgXJRtCYcu12o6DHRqv
oVLKQx1l6vDdsuHA07qljo3AHMY5aZWYL3TND32f1rz7FytAwL7fHWoDtNM5W6zi
KlOtV3QO3DmF9/hkAuYCES3dI0UvDjtcjam2foeEE5obUPRMwZBM3YAsLWsd7XtQ
ETIkgWVx/OqHJHdCfVPBEEd+OR074OSt56ec8PvyqqpAXRiW+mhqT+4dzpxtsBPh
p0GWqbG6CI3zixrH+mBXACnKWdUjpo/2UVBFCPwkahw2acQ6wjxXp06ekSjmaMra
Z/eKFd9QRGYj5efv1z7qinVkHLt6/rRsfhw0wY/zBU2OJG/ESJLxmUpB3pEZKRlo
IMU7SamtHf7n+lsssOFlG+1S6kab4MOeY1LUfaq1GklI1exv7oPpDhgJ2mnOMQQB
r3ShPWjEFwSWq8MhCyj7a1zB+NlnBK7lks56FFJfVssalfN71Ph1Eaf5QeJt9F8V
Li8x7jRNFRKFIJHB9Zmv1x4j1Pd9ehB/of6iKWD5k7vNsPkESY1RRldZnMyth66q
YbNmBYVeZ5h7TU7OoRDmEh5Ov9J6MLH0e82tIVRHsZx/smZ5/6OgVFr5R58QhhK4
OWWY+FT0gMHHKtxf2TRturykwqKbRnd76ftL5kwlDWjuTBz/tIdiWXUDNp5itORM
hO8egFSLU+xRsdfopgucMrnwSgMAY52nKWD3H+03Hd1F9IMru7SX0DzmaVYlhojG
deR+ctX3kW2hM+WVErPdzbj9PiXbFC7qtKhr4uUCCmNfAD5cbUE0I67YExXIOSQe
H7oth24sjYXV2cIGLNodfWc1seeAfWUd8/lij6bUAMCgBjaSUOVxKUCbT+3hSu0c
vIxm3eW2XTxmdMhZ3DCXTM+z8AMOB72KOSys+HUvraOf5y+NV/mWbHUM0ohmeK5y
/fVYWQ7vCeXUa6xoFDI7VHN/px5PBtGYsS1KWDEOQSumlpTWX3oPLlpjJWpliFX2
GD6mx7cO8SvSo7e+OxR8kTW6pLB+t6kSdDKQTqQzAQpdSbq4b+ZVb6OJuy97ldQ0
3dRfkGRkV/GNBRRFY9fqxkHrpR7B6MytvveDq12CG5bWNiO9Ou0jlEhEcLbAToTC
ipy4oyHTnI4crR/N8pybXdPrn21JpDy1vuzRsKMp4jmJsDtnKSs6vyrgItzRi8Qz
2udJ0/BA0DTXLJ7K9+lNXjkSMhjcaioHsBD/lcNZefATp3gFBBAQ3zzlD4cdcfhg
VsKGoQHVcG4QLnud8TxeFM0SA5q/6UnnFkoCJe/IPiJK+j2XiB6Nvq3JedaM/wFz
vbrfXV1tiiTXYNd7mXH2f+C2h8uTweg5nJ5DTY/KUXHO8mlkY0awFjwhA/gO+jfh
AH9VsibBwsLxCkTsFujfkOtZu6NroCmpsYziwG1Sfpto/FNYEVkjNFJmRB3m1l7c
zlUo4CVACClEK4y43rSK7/9C/59HNIxFbjKeghKGiyY7a3cCUG9axJj6k+yC497J
EzzlwNKE8Yd7ETB5oRLo77PzrKcwBPswbH6eRnfL09tFBm+U9e+J9kgV4Kd8/aP8
REo4fMS3pAoFIbmRzYgRm291hSHNn6EkISlzpgT3iwtL9xAmIa1QbshNqDfp0WBc
F6dT+zQrjwxavBALdzynmuSXL+3NecJfNCVkoK5rj4MnFQTAsxqvkkbQJ1XyB5zU
9PkhYEz4MT5WM+BV2oBERyhJjDTPprT21Bxisw5kocR//w0RvXSvGFAICrnn4qep
fnOXxF/D11njP+POL50tTbvQ9FbQTk4W1hUrX85DmpGqMIJtD6xEnlBTcZlQ06iG
wryWz82XiyCd69uzWxKzINqm7/E0hJTq1bxZgE/MjJoQz88XJrYqJz/Go5GOMZsR
YlOdvoz5r6ojAc3g003MySnbGgIyi9OdB3wOMKw3Gu52qRsL1MG9yKjwNtyR4MEu
WeG6MDBvBSwdJJq8+vwS7BdUBvRW80miZPQ9XpJYGHsgYP31+TuYUPXS4861c9GU
ruQdYcYfdRIuMNkY0Ex0bHwRKEEWReFyX24C/NrXOm8mcGUFKvMe9mjg6OGyjjyc
vxn9UhIj3ZEe5wWFiHPBj9GUvIsA5QhsY8nqb8rcYAWwZvn50QC61O0IbjG70IGv
M6hntx0M4ctMKAezqW4G/tFWpkQnoXzU6wOH4yIBslmhnkR3fUYX203Qw0W9BX1J
pDbAEap5kwI92eDjr7N1WHh1Uq7TP4fEy5RNrBYFaSNtqDtQKrpMwarRKSHdGXJM
+QpPHquns4jKPCiJlT/ekEZEUccx6if//PdC1UQzhbcLyfNnE7xzX+3jG9q1R3LL
YuouLS6iZRbNkQ/UFVnHC+gwoiTtGuM4YC//HJ68/fD3gg/2rRvtxTpPBxN1MEfc
PDtTmqp+YvRmySQfr7rNgMP6GbjigOwK4DpWWTxyLZUH8bUE9RjlTXnjLqMqEJzn
kGFfxwxbciWqebm5eGiXiGFKyEP+t0IvtvUw6bLSsPY+zIPjrXTo7fiESk4LK/Ws
RWzK2ELFC/66yvEqMQgd7GJRNEqof/Yrh+xZOZhYi1n6ziFnz6merpEdgZzaDS+H
zRAWbDSVT7BYmnKnp9smOFmz5LgKlA/w1MSIhEHw9ELqX6gdQPrNdAekWEwV+zcw
7mTaZL8U8bfbUGzB2jPcfj0SVbkC4cVMDNjHnkQWfZNInnupoOL8ZWOhH+n1PJwh
zxdTxjVT47UHJsGULoCdFtcjaeNIk1svTI8RnaLBzrs8EghsdXHAeWmNVAqZCO6r
P8YUWHTIwxCYsI5jl/C5d9AUllbQ24TmPH8TMue4ND1oZdhaBMxeuIaRejo6Zvnq
AZ8JyEoZyMiZdhbJLfm8+vWKO7SQH4JuCT5pXWyGzJG59K1/wz9O0ZhBlARJV7MT
1bhuQfEdZvacOiUbjrJY87qM3N9F7f/WLbyAQ4zOpyhqGESkQj6OJ2q40vy8Hq2Z
QByJXyfaIIqqJibx44mxiXwZFqwtu5sIVkDmH7MtbPqlc3sgAUfoCian3X6Mx9/R
lc7nl5GzsvIrrxglW+XdgYj6M/VK+0HqeLDFvqvRaZDed/pNFMQtUD2K/6fj4ycI
q73mYSIJfN2bz2opPK4slTDNsOEETuMTKa7UjGK8BXxPvywqgQw/gzbEWhFCZq6E
cCq2HrYQfTg83eykEbTnjMpTEZnG+U7U63EL7pHQGyrO+G2ucaAVKbcQioMJQq9k
ok/nV/lNXt85ayjg7naGeOVIVIY8mJQ4SbH0KZiz9GH5qTW2Efp30er2FqJGaVsE
+8sqdZRKoppRW870T/OMldkWjDnMiiRvYIAwgmaYXqh+OYes0VQkSyNv6mY8Kz57
0+CTeETJ1iU7rSy2oV+AwWgT0H65KaAeyasL0qxzdYyBNHtv8SQhbah+joWQPJt/
lgU7p1cAWAAB48tyv8ItMq+DiyfLywZsIbroUOJOde37g3xoCVEe/uqWYhTTBnmO
+o4wI1fEBAVFZ7ICXBE7q872PJbqimR/5Bw/hNq3WYEwn/fSq9aQp2XFpljpoY+c
iOwB2g6luZXn7ZZNaYMQpk3FTDM/X41AKmcS5al2I2wSo17IKqvs09GfzQ6fW/L4
1OtcZw8kUBETaUMiwLreWqotxgjDTVFvMIcDzbzXj2ex3xXrmiNDypSVKQfLOEVt
PE6/lI0jnsB1fqfRCycoE8FmCtvNJubX5gMtSza2lXM54FniP8hxs35hIQWW3ScJ
0mpoJkOEPLr6NembF6cejyRY0QLBiWS8jgelxOexOJiBrAEbUWuu+YtMbF6GYLsQ
D2AeJuET8nzIqCl1NHleZvfD4ZPcHj+TR+2tqKo+o2QpnkOWF60P4FGJyqX0Oo1o
UfnQkW6LA20mlr4qHkeadd4Xu1OlicjAeNU86nKwxXoEIxkS/D/0q3m4bqA/NozG
Zw2LO2K9MlZSDI1rf1N8YeM6m1jSpQaY5+fkqTs1zk7DwQeVJZa5Liq/Mj8wvMtw
i1RigDGGybY36zd9jHDuXXYRBdezGiGHLyAu5PwXlco/zx6nLxE4IpFsbERNg0HN
HBKlqaTj0Ovdg3qmrjls+hCdYGTc+gmom+c2Jnp6ZcCaChlz8Pbi64jVctMChsZE
nfU+vwweal9rdERi0eZbrDD7U0jblNM395JK1l0IlQNcGLL8/x6QQgsGG1qndE0o
Lj2+AK0rmWqVoWvYwZwImItB0a/+Z2i0AhSQZvxWPE+YtJT28p+QU7loZhJ8LHPB
fXpY2F8w5P9wAWvUqAvjFRmta83yg3dvQgJkjogxoogMCgp4GwWGDW35kTEYg89D
ftWX4N+tNWsqAyLOP+Z6WQyZl2MWU2gAxnoiDbYzMPmk/Fo6U7VUbk7OBPu/LoQI
h1Z0FKISJAGykhPw96FaviI2+XYmJLQyXswE8WLU1Rfrzk+tZmUCh1A8du40NM5/
J3cWgVyZWt8T0xQ0IaG5GVFjzysvindnU0f3RqRs69gBLpiBtiRMTn1o8wl4k4F7
EMiRqHPe3v/cmg8B6cjd3VlMVxN6jSYUAHNXY6+JGnrEkflddwbOU5sMSeqoas9g
/8bSj2YqQAjFcWgsywE2D+2HFc28VFjCaS9xPqa16WsyqQi2eHcT5Rpoaq2mgFHp
uDGqxLY2fbw4Dsx/bBOUXbCXz3BOrxLPUlvL2mWDdYzmRHyA+IrSukDvKeDrkPSC
NjzB1uMb9XqntO0KxZbW6MRoIg3zHJvJdeFs/uolBvYMxQJGA1pBJXxkFLNrQ1RA
t+fS7LKNWuAo3fKa2Vxw0xfr7GJe5GkZXLx76onln0NeMu3eMpg+ajZ6+8bwzy8T
gkRHPh5HieghoH5W7M8YPGsTCcNWi23F90WPy4nkR4IslEzycD0fniMp8uF562kr
U0s1KhEv+X0WJtRslyBLykx0KphKjW7vaRB+s9PUwBd0mKVfibt3FttDETnbKcPX
zwMa0GRbI3SL4Cv/RDKhbvn8A0cVR2lzcPEooklvuhxdO1lYvfaGTMD2rK9VcHBT
FwcMzqzqjcg9Q92t4FeF+h4VCmA6EuwC5R8gZdkQdNX9BUv/fFBO+CGOOeHq/EHV
EwFJxCYG0xiCzfVaTIeTjYqF5Q/0CxomAP6yCMNp3X+rnyt0gTodZDnslGNU3j+A
S6cpCUWHMq50DhaLOxJaX0Fhmge+JdfUk/x0p6GEcNBHKwG+grvf/RAj+JGVZfED
jAAkqk8XFPkyLKqFmOyT4gcDbM4a8v0RGkIgkmXrf0mqITNuLX07ELV8j5Kra7AM
in5Sdv0lfH0+iHOnjp9Ckv95tZ3LBV4d0h+w89pHGHG4HRC/luPZz/uc9iF1jhxy
CWY53fP2cR0ikKJY4qwSwXjDxQPwRylw/DcBZvUG/C420TPAvtstAmKF1hK/EcAx
oI6ecOtL39+DmzFilXavWcytCTHlrTbTClbQq+QCCuypZCIwskgufLj/91omvLfF
QMkP1GdUWXChP60uq+RDLMqyePZepvVrMSuDTvk/Jm43O1+94qA4UMJLr1s4KTbU
0y94T9C+NhZetD52d9WSvME99l+0tOIfkUhrGjxC7xqSLnrYZ987IxzxYJdO06Ot
QfQtNfqbDqNVm8RiSZ1B3+vYCY8+iwEV2EpdxjCr7/wpDb3XAvs4Ss7T65l7EA9D
+qjrghy6FAD5lFCjFSIJX1+IDeoGs5uh7mL3LJEbyR/75LaZ6kcNcd3uUJ/MG7VK
21H/IPUk2FJIoZA3uKq4SU6Xrnx6sfLheT9g4DV4JeuqVn4xIE/r1MiSq/h40daF
5JrxdbN5z7jGCF/iIjBKSX0b+tMbcWuYSrHRpLYoxfxxufjjB4+alu7RCDpXyC3G
uF7aIxTXhccDjp4fodRi86AFgVq2PNpei7P4U/jGWjCkBiWX/vsy4Brb2HmEbjUF
Xkiyk2Iqqz05UPF7FyDHUrBgarGEe0R441C5uSX3EN9cAP6VmoWwHKrWDf+ayxdC
RF7RqEQbEAX9bzuELE+tMlrJFdt72t1tnvwJ8uA7B9vMLhBaM5MJhDKn+EGERL86
2PDz1/sE51Tp9KSP2tKVdD7tLDCXZo063Mc/rSEjSnzDP1zZEvt42C5EzwuqUXM7
8yb4fOAht4n6bNIl7JsQbHGaVAmpeEfLsD+XEj8HT0kFebO9QzzIGTyCCn5i4tXl
J85SMAZKRc4AXfB4e4m5bOGFCcHhlJT/M11c62J9mDyWA2bTWdtveEo/eTlcE9Ac
bvmAl+PjuTlQWZjl8MbfLZCtPmnQzvlUkH12jNrY7kjWn29EkN8Bg9ZZJqqcbLyf
pJeV8mlYFMeEO+CrUnncwd0iLlNGZcLKBbvgAKqS6LLZ39kfwU53gHe+ArWKopA5
Y0gRwePae7KnAew4O395Y5BWslkvVVFcx1Z9XLOBhW3CgbMgj9HR6d2fmwKUWC56
3YdLorcpaTixk8O5vK9MzkbHbLgSPw/emcCg5qvhSjxd9ILqmrLZTZVOkGWWN8w9
tWlWepzgra1VcVe809EqEpVKR4KF6zo8s2R1x1FV8kB6LJnbJhm+nXjz3XvRaqQp
h3u4ivljXuiuQ1smplrEmQxAg83bn+UJObYKHVrIOt8cWub5L722a2APojn8YXpn
Q13fTE5WSGbHmFbha9HbxMdVfp6FWm2sqHiwS0slpPxRy1ceIFTu59ab+kSwX6Cs
zV6geP+FaEeocnqQUCa8yYklaEieFXcDgINvz9glmBvL6aahzH+TI7EmCZwlUa/T
S4JgQ08YMJWa5LRBhTwg/J7acU9c3laFS46ssYCuSJy1G2VhxOXKXeGj/Mwm0SSN
Dk2nUiul4koBuKGhnRrIdgfXpfQCRM4T5E/dxQXsI1kufTOOhkjE7QkqTITtPswS
6jde2HawaIk2oHPzdHMUg96X/b1Dg9MewQhpYbZ7QdbAIn6OTxs/RsRwPvsxeeAy
z2jFoRS/5IRulRGl5EDVGpKG6pPomhf8G8u3xDT5wyPvBUXbQ8DPzghlye+Iplh9
M/ScTPEfuFezz36WVdZBBoZsIFYNtSTHnXdwSheKloHTYeGN/g0kuIKwWmm6/TJk
vIadML2Q/wa7k91lgPUsOZKFia0RmDT8wRd9YyQpxgDW4Uv9GjJ1t6yMwwLh6+eI
zWrX18AJ24Yo54Mh0XWahol+tVXAnMQ67tzFam2IIot8754zdGFHsAlPZit995vB
Ua6S7wFSo13M3bbLPrg7N/EuL/XZm6r+A0NyigdboXZWVxHq/Nav46fHgnw6kv6P
dzXvvAdIe5DFs8xJ5FSGvpQbaiFSJ2iZ5WEuWi7j8BpmwkKtwvh81FRsvjAyuBY8
ToCwf+Wy/zBydWz6YwFH8v1I0yHhA7V4guyyFoir1VP/FzyxhUC4pVCg08YikVZB
lm7xFixBvjC2qb7i489YDZI8THzLnSU6rRAWMgWj1FyjDvXB7xE59IEI0KbE8i6+
L0Dv0SI0CPnOmhDJRF0CseKH/NOtL5XH2GShMmB1WMjzSV2/IzofJz74Bb1C6bhg
e3YleDt3ylPsnsA3aKL6rLz/uaPkXYpBzK8oGu/m8Nw51eAkgpKbvAHFBp9jBAO2
a1/5pqy4SoOHTUrfLRIiRPt9LUsw/aZS2pxkaCinPUqhpYf0BmUFKMEQilT6+EDB
CTSQbFm4b8ywN0rlAmqplVHDwxXi0RhMBY4Lq3kZ8IPnGaf3v+sJp7Ginv1sqIG6
ZFycb2Z0GNhI1bzeLIzvn1NHYl7Rhh15X+joetH70s0OV/NYVuOdmvBsGNbJcq2E
L4SsuLNNIQp+FQCxTqPSf/eoC8lsoi/Ljivg328Y3wgJUQrHBzae0JZVCMOj/RMX
2GFDj1Ti9MF2LlkFM9nBRcAqQSMuo0Tv/hn6DEyoR7R/OSFvg378r1rWaFsNbr6P
4NjlI/0PLV8U6cmsdTvPOujPvqLpwht0ZLukrNMZoOP23QAZwo46u1GE1DlZsOck
jAlgSVGb6Fry36bHD2eKiK7wUGoihf2n2j+7Ss5GHE7KdboQ/0w9IZnnTBRr1ARk
flNTCNb2CgyGVgTq1kOYob/zLIoAL5LSK7sYfNQnmzaAAvOQCct6euPCsNrPu3MF
+bzYuknB8PPgCL1H6L1NMIwVyEe68/sBsM8ll/KWrhjP5JkFTaBfmkyqzSAyMltw
aucvIhpRJW1JQGktPKDQRZ1rtcqlL8CAo2gP/8dmzxM+6xcTMmM1VxQEv1rAe2+2
MSNxmCjv1I7gR7gU7y8JjAKhR/vA0/g31ijezAQqaahDapmod4rqFVGSgj+clAx3
rTWChxjfNpJHQaJ6EEPnB03u516RYPWaiSuB79B086b0cgKwz/InVaX0QLEbiWFp
UGlo4wXnJMgT1kHBnMGlVPTRU1STBF03MkQsNfVsMBm+vkD/flcxKWrEfQt0/vEe
mJlekunpp7Ea7L/eJ9hJa840Y4g14tpNXRSo8l0p08r6ybs1D63q6MqCS7G/R5kk
ESMTEkXo5jOstxgCD1uMfecidc8yhXl6EIFk01To+7InXRWzLB1vVjRjIfoLnOEQ
Z5uEJxdat6/LVzHgXBKv0FJedSIiiIEmSs9VAOfmn9NsAXLUt9Ln2Q63SDmVmwcD
wz9Au8J8IDJGQROgq88jnQIfviP0/GFLKTSuvUDxPRSgwJgaEuZ6kkfBhmy598sF
Fh+2ZCVVr2q6tQTx3saKDRERViL/rrwvcl2dYQuIf58xgmzCbkA4qALrZzG1Lb9V
Ezy4FdlR1E7L+424vxekD/oQ82sohCtI4HAD0A5Vr21bKh35rc/u4oo11lXhdyE0
LTsrE8Y0tTl3COh+lYed1011vaINX1b4kYNZPy0ZImnZTs5Nb46vKa7uAmHyK5r0
TTdvtuaHzZtrzzdm8WBEUYyAqBaekI29bcdRnkQeejRyTfY42JtMobAqrAFd+tgh
xAfptB/a94dV4RMJ3KyvyvmU1Hs1PTq1wNkO0rlQMn/bhvO7X16PZa6V5Fjk45Pa
1tPM2Nqd02nT+xUoHeglweZ5JM9oFSPqjegyVIztiGecdRdje47Rax5QedXDR89V
ojSyM67fDnJN/BkXneBv4h3RsYkJeME+wWyWyqAJZxmaazsn19wUwYa/NztPswDw
uzTzomQ9MZLpbUPrR6EnGa1F4HxXGZDcZDbcHeH0GmJbFHn4RiqwMMPCB/gHVb50
L63lwUwAtU0vO0I+Owjir5gJQwtE9w7zz8Kpi2CBb8tRzn+2YHC8bNyjWTlTacUQ
UhBMxcWL8dQcDzlChc6sZCr9vQz6bQ2dpBUkONsAzLhetgGisePUzGQRO+T51nPA
mRvpZapEc+pVikZaxAgcMcbrhiNoplCJqBJPKHi1LHpqK4XiLKtYYcxoa4tK1UxZ
MGfKE8qtPKQjw35hQD3PvSI8KnP/G8DdyOSgtqdgzEkpKmBr0P6q3bal/TnuUQlE
42pvzTgJaSAz3Nly9s3FNVSM7AXcYtOXyxfcDcTa227P1WYESn0ZX7qcN2LLRlM4
CqjnM9UIIkI7bmDdJ5dAaS3IKOzOrVj+NXMePuamcCSUA6bAluUKXqJWKI9LK3Mw
XMUK6NswIJgzwWmyDeOOeP3Pe+S/NZqoLcLLzk+3056RouLcnUeVh31caa4r3hS1
dMRAuNcFl1GBSyYjKAm7Z2cgTOaick6KrX+h3sfypG/KmySDGQbFYxsG9AlpeVHo
d+rMWrdn7Iqh1U/I3jlLOyxeyWnaxtiTrlZH7kXn+lXMxDCjL+1eUOv6qjVB87aq
Gm+cMrs1JI1JzK3STwoZdGW3viuB7TFHZRQbtzFFhFwZa1orJvEhM0SRNqgm1pYB
xp3DsOvBXBk6K7CWwACOVVurA6lj5a7nHlkZgo0XOlTHPhK6XySYX1RdOSBv32ji
/j777uozX9JNgPuaFRl48a5U9/k2+7wVhFsAuXzuEtSWY9xpUQTwvBteK55nvA/2
BuufdJVTn127WQKTu2S1dApiyqiTmGBnwBpW66QujJRAMNIqj5nk3jGLlMWYkGtO
h9dMrcM0U6NScOTlgYKs4nKzVVlPpIvic8MPDU2g8q8Hjuek89I6Gr0SUmeN4+wa
XWo9YnI7HruwZDun7FZibDYs0ADT4xfsnh2g1osb4haFAcRlb6qvr7Ghdp5XGYbK
9XYa0/JwZ1RaVfGamsXS/O9gzfi1zAonnlI9agF9kDZvZk+7cynWM50gJKKziixO
RwNkuvFAiDOnOzESVmk+7TCSYSq6O7wGnd2vJkKAl0NAKLtFxwaQiOkMVIQuI2dN
kbJsVSKkvUX3U109e6tg7a5hjohLuVPeS4NaL+RQK/4ASpGJDnyReFI1iLAIQpDX
T3zoyf/BeGqFVb1DxUG7w7gvrEIpYNn8nsM/qLevGYgoUVHTxIAszSBLzVPe1mmA
a+ttg2Cu0izybwwhOtp0rcH5pkA09DF2QGLnbyFcbiAD7moyxKp9wKI4MGISm7uH
Ya2XlZ1azdeDiYp0rsdwie9KdH96wuWhajZPOvVdsdoFIB141N6VLTWhyvG0ev+u
VVq4YzcZundbr/Q1UC86VlYOjrvo072fzNDZ/RiTtx2kh9hl/iY3cV8lYDS+/ub7
aiWxTcxkQM+cJ/fpBDzN1vwL7dq+6M7yLj3U3ApPmRi66gHVHzJQF0BJE1Zd5efc
9fj/hRr+dM5sqKwyUOBW7WHx/5/q/C7tdJ3qIu7d1waAxShPgqpBVhCshoZKMuo9
9wAuK0tQfNP5JYeH3Zw/J/rdqzOKcsCy1IzNxxXaSn0d8xe5JJoYlpDBfR90BSbD
m33qmkXF8L9ZMP5v+C79poI7qtud+k+M81oMRA33i0op1g5RdvmuhgZuQwQmtDzv
akwGhPUTqiHQq3sgfw5tN2q7SJF/77W26d9Q7fiuZ6ilytHB01J0G4jsqZOZ5lXv
05mfIbe1va6q+Q5pP9Tmajq5xsY578my/WMEBrg2TyWJA1vwgJHxe91bVW5AfhVp
MhIhp59xkjQVCqsCMohjZ3fkihiNmCdXKOw2n+QaL2Vy9kdxqkx/uHeXXZFg5w5E
ND5QyeLqz9/7AFTCNSgdT94EwgrRGRDrkf45X7eiRwPyVBXxbh6x8k3OoQbLWtb7
u8Lj5+4+YNoCaxib1i3YSSSV6UNIVyi9SZavOUgxAwM4XpHLIlYNJ860E5dZfCMU
aZeA7cHN3rNB52avk6hIqP5qxcrIxDG68M3OCewjuatVQQoHnJ0pH2KurbcWYlRs
GQ2mlgGqaucBeiJoJRREwBZVhmr7xO4/iw+/FCdE6yjRTOOV1l9ArzYCSsrqumCr
zAAFc2sGkXI2EaeU204gBB2Ac5Put/1WrSa/ce8dG5uKfUE9pjrWg8Gfxab4R26X
SpfZYvs2YmKue0gt4puU5tThMtrg4zb0kCkEtPd+2W2x+EfUZFF0QJATED4Q19Bi
KGnp0Y/bL79vhyiQ0ziJgN90e51j6qnf4FL1joAdXlmw2a+bVncgHk3Fyp8sRMtQ
dGUf1LqK8X5UXAi1ohymO1VesmKl16Bx/PZlZ50gVhvtpxKTaDCnqSGm4nN08pB/
RkoYD81uU72FSkmtqKZ3yJpAMxejkndWMTNHYQjX9EnvX2F0sA99Qb3RNnbYDG6Q
FacKOUIXLPKmPEGCGdfasAuGE1q/ShUZLzROcgPwsG1wcGcLHbtJbYzH9wRoX7DZ
0s2aSX50JU9kxOHO+PgOUvoSSrFi3e0W9/LUkpR96gvGao1XO12VN0lYwyIclE2s
0veBEjTpI3Frvj/IN619u2NvztDQiEfm+NhezQNT1yhNCPEs37PcSBfskVhGxK6f
OKfTAD5egJT+a7YO9nn8Us0VohnHVDUVwWHO4R9Pi6lSfx863RV+AfNYy1eScuIL
cP8O2SjXdPHcseV2wpVaX8PFmi0+YrByCEP4SjpAa8CLxODazmiBGgP8cu+89lKJ
gcGr+L04oEsdGryf7aIZnAyKcrw81crPZUJM7DE9FYF4mbI+wHLheelXYV9GCTxx
mytS1eKjq7wQMayk33W71YnEgiUk4daZI/DUMHbeF5OUA4twuHg37/S7U2FVYjkw
PnF2EZpp5x1DSeYuspDiHK0oo4KoarDznuEcpolU7iXtAgsvfIUbSm0UqY5U4EcY
AWwFOuiau///4yxzsiUERNFRm+zr6ggmo2wizFFHWj7sxkzmgVr3rhz6StfqUkhr
aKE3/6QfvWT+HTDwwux8cDhCrBwm2hGuTrxSgTqzDCGpPQbfQll6N6pLCaDjOpZy
UoKO/aaoem6BN6qnXSIY4BsqTEW4JVMXsoUL4KcB1j0Iy8IEf6RN3lBaVD3AYK05
tfYmTRXG1G1+uS0W4eYUZeE1pvTa0DLM+eDIIY9WTDyXE33Z5U9Tu/xhmLtaGSz6
pnk+Wg9M5sFXhHi33Bzs0yA0oKMuAGKS/ZA5555bQR9gQCpBABKbFglveVafE4N0
NQTlP+YBBvZsjiv9rYFrGbMutbUW8S+DJjABLUIGGSeOChAUPqv9LHnh/9900sFz
j7hJzoS/+PDYn4LLdYXAenNLEi6iwA0FMMl7KRS132tLJasJa1yzJo03bfZcppDL
vP8v859fK9zfLViDhuZAB+WWPnC62+pAAKvbVBdsfGN6O03NZ2iq9Bm14ZMLNRTt
KoYhrgZnqXbYJGjGlUYr3HZEXd0CprX1KV/L5Ee4H6pFK0LujjTxm2kc88vIIVmr
Exw81/74kXI/E4ETo03S1jZfT0yWYR0qXmquf5LLL8v6h8rZxkSLUDjYlb0ySmJU
Bw2H1TupP3nBOquy5KhO8yVjErqHkuGIVXlGxdhUELPZ3xH8Ipd5tG9iY0dBaB/t
ullVsiEEJilzPnthm6raYTHy43B32otSVtVcbnxvDaRg+XgRFknlXoT5Gqd4oLSa
SSwps6eFMQKNrwowuXbyypT6k6xVxSaEXPTWbZ3iIRzWza7/SZu34y5MkLpbjcGW
m8osRyURpN5I/fuTVnpnKJ83Kj336IoYYyx/6Ie1U6KUxMgSlN5MQLZJbq6T8qn3
aG72kzkLj31YflyklWuKaDD8smaq20+KshnzbtPWHafhalHOKCaW7/sT2dLBfQuW
GOJbqsXccdCflknGuyXD3m7jnRItGJzQf4s5sKwEvGHVdxlfgHICbq+QMUJEa8Ea
86PWP6EG5QzlAdISlNOwbq7Hb7kQahvhyyQ8nH+xR6zrrFnUStteC2BLAnSsqMBT
tQqBPaE9/oII6wDUPhF9b4MMk/cwgOo8UFJNHUQRfO1f/rky3k6t/hqdXzmlysha
owHTxNWY/L8SA1BATi8hk4mmNCQXIBjEcycGqhmAkQQUkih6d63tJaFSTD4F9ZoM
/8CJIOojBMFUL1OKyEzFEAq1qdf1UppQNDkAaRtlWixgqEypy+GbmMsYHoRFXfT/
KnBZOPSFCvkuePz+qGPYU6mINLtYtACy87etCv6iMDZwI8bys3+I5OaKBzHdkemE
mRgckVsK4bg9m6UPfUrpcS1nn5rqxVmM8HA9MB/c0DQBjUiGQ5GkWIei/Hw7r8YD
ZdtwuE2f/n77mT2GctAPdaAaNRK0bYrvtuymu5RfDx3mZjahqbcjIPDlJvTU0Vl6
5IN6aKmD73IqrLXTncHAwYWaVArVgZu+Dgkb3UCtZRnp4BKRt4aNXmLUUjhdavso
e/q/h4Z0bW7kSgYdORuXPT/6HRYGGCX5gqxz0PQB8NMB25JqJnvAhdprmi1uf4KN
axZ4aljJ4N4SwkFFXYz3ALl/BjQfMUP+fnJERu2KX3cur5QKb6WsWcclAXuFoeqL
6EuwL7XQP6V+l1fzDU2dDEG9X7jxD3xwsyvVErQjcIJxhEBYV84/GZUYUzuKvlgX
EdU90wUgDmyvXzdJ6Fd9k+jhFaFkaa4qnby/FOgaTzewMUtISX3jzn2bkP1fpJ6W
vZXz8BDTqE4c1WZqY6FI19uqrMSF9P5+tjMbg/bgpXMx+Zmj2KKWmq2g43AZYxm5
ugSu5Cqr9febOzXXUSFpEKbbdbzAkbodf7cJ26/PHezx0ZCQDrdzDxwVXVVf+MKR
GdxkyHwfRuY6WUyBYCKH1nCCKKitNyzaNUIOajFFBkTv6Ms8RkAAdWfWSHCrzkbI
In8YtHW+nyL82SdER8qPZnw5Ob5NJYyM2OqLfsvXfNUYtgyza0MqeNnN0c06WPD/
JW1Je31SoSEJN8LoqHnKCEjE9rBE1WwSKw9pFx9+QAlRUNPAB3LOJkEViJ2HXaTA
YL8TR5I5Pf29vx9DERqs4q6nyRZXkqxRz6j3RV3dbsV0EGf11EzkrvLFpk+dqr84
5IQu3rIwDO2tvujFQQ+Rd/fpaPvsXy2o8p+ZeKDJiVsH342q1c7NFemMKUKyj6i+
uwLM9rh1gRgdasY/Kem3r++81eknVqzgupPp4NRnOKGPTV3PXXP1AtOWuuc7kHGA
Ocyh7wlwehkI103yW59vTqH4cARa/qYJ+xP9DbBcAJF1+hLmKN9okBUC+U/O2euG
mfajJn5PNBsJTGQUqzH19KFxCjZ/WxCMJ3WumtXEiXW6jIRxmhvOZcP82aCArgoA
ASQjnJ9VR41TAggK6d0U3rE6UuUm9iKKIsonZMnX8szJ5CghMQ2srytYCOFQENiI
5k6pp9wjCu3OqQPjfffdLOKy7dl1aQPQ9OKw4rq3LF7PbrwtQ9blZedBqBVV5r9s
r4Zsaw0YS5Rvqtfmxiy7z/1WfAe6H+oWWE9JQfSNWT0ebVxaJSiSaQ7+wfD1X/T3
l+u/MVlaDx6gQvDL92OfWvhetcVlSbk/GX/D0/Y5/r44aKtWk0dt1AexCdb30pVP
XFKugbHtsAiLJ6AQJw35I3z+lY2q0OXIHroJTmbmeJ1CeWVRi9Ufx0vh82YdDY9m
c4xvHiOozf+Wu3y0F6dv29HNwgPRNrL/1zRaXaOK/EELmRh05QS1uFf3LmeyYFKV
sMfBeF8ty5YoNd622YazQjp6sW5FZTd8XRmk8473fVRc2S4yWC0v0ZmpNyVEf++t
x7jEGrhzxtnRGywfpc62nySrkCj1S2LZmWsfPz5wzxSGDMgsMC4tDHc4ZP0OAz2A
mhxZuKaraN50B2E5blSxSwE2+1Ov7fUWNa4Gx+jFTTbLmoVGA4xG8qB3timnyAhR
7NsdT9/9zC8b4fXcxqJth6177TLRPpZ1RYTVLrJJ2PQBQx9ESAyyi+wehYX0Cwbd
+JB7+Sxk4MZCjrzU/sXEQRNw9NPzUj2TLWv/bhx5D6NeOLXQBy02A/G3gWo7N86R
4qIkG850HAMbRYRY83/D01zvxnXwXYRbovmxUZtJmPYKI331AOz/uWgNHFxlUIig
UDqxPEA5s/oSk+1/WIKD0cMmrxTlzv+C0BctAj6pp8SGci1gHGHGZiMiCzShmPo7
c4wpI8ITaJL5YiRAU33KHKf/geeVUzuPWPFCjm0KPoi1ujhy773SUlA+putwjLr5
EaeHCWt4yZm31x62D/EbKWMcTc1bya5Z7vmG6TYEZSEoGfl8T3ZKXVk0EyH0ff3F
2cze3fCoIow2KX+es3iRBCnJR6uAzv0g0iuPByB6UePB7wtLMkA3SZ39y8w+7WOZ
zU4Np5my4oQOYjnWnDmFDsSDecdmWU0vlezd59a/Za0swXFomZNnWvzAGZF/Tt0M
ERgFt6x/wSB1QR4o5Kq02n8Ib/C0+8RR6wxze50IBYO/RwK8b+j3uO20afTX8z9d
nzR2WDzrBdxr9d9Jic0AmwHvbUsABLfHn3zAripgu8vYtLFoHdNUMr4KazAa3txq
OvvUIClm1Jr8uY2U11jWUgDmkT1/mB/gKzbI1w5Me3uFgTqYT7SquOh+eVW7AN0o
jmsqGtIgaLpZfUgPkOW2K+HLm6S+pcYjAmGoRwx3JRww30BQCuiRfPtjaYRwPqeP
OfagsBqrDN2kFdrYVgwADNSLKzf9xsn+ZN1XEXY1qJjyncdz4EFU+ji2YATXXSfr
oYqBmXuUNq8cyHrjq/tN1HjhcASlRw/j+OZxNv3SJwqsfy6++k1z2UeW0pxgEhzP
cVgFcpd9dwB32OzIp2tXgYtpS4uRUcZrzledjy9wbL28WQYuGnQYrqMTRiFRL+TD
Lt34u2zsSyU1ZxOpLAS+J+J9fj+urFAldpCRJRrvpenCc1kZQzWHNyby0RyiSRt/
45KDc+e7xBDqddZqI90uDdMzo2ErUpVBYN0P6uZnna+CwGL6W8WISLodh0XtTB2F
468iq5w4ayqKYcY4mUr/ax6v/JJ4pQcaa6SYylz3DfeZzPwYu4B5+juro+kwT076
9mhRDaYD3AU7sSZNys7x16ndaaL8Y5OT95Jn2mqM1wA89iJQTfTASNhMWbO80OXt
NFN7zTDv5VQAM7PTrMD+xPH+i0mNRe9GBW7g1tyV4ZIUrxkgtFJ/XXzzsIWvBxjQ
NIsKTz2iOkIqoTtkqVkuTl62i6LVsjh091QKI5qgKBs3sbcX8Lkan7pGThTaXAaw
smFrJlRI2O8ea62mpXGfWoMNRZ0NSIGkjXxgM1KieyuErt1V4HsYBFfI3CNd4Pvs
+3cDu/GnwwrUGnNebKrC4o4xhyBc5lBSfHMvPtb47YWuX/d5Cz9/mweXftVWNxwc
foCXsFz5LBIAGCgrUxYfNH2ruAkomf0eIMjvbpM6ME15t+k64d9nyiAtV4UfzEd6
GZIAjw740eUOSvzqDUpOlzGjIckUChywmzA3oyAJBK8NUk6PgrL8wbXF10AuI/1Z
VpKo6/FsvmuCUtNYdQLUiknG5upMOd9O+ZhFU8EeW5scTmu2hdJiGtsIvDb028BS
9o295uEBeNv08OmRIgaM5k8i2R4aU9NYICuWCG0mdHPvcxwM0RCpd8BG8YcKuyn2
ycChsMPwVw1PCMRyv4FLmn2o+ZStp9NBRvc1LkzGqtOqCos+0s9NrMr2UPPiZiDD
3AOO6j+/ky+sNx+s8Pqf/dXTc2ykACJo9ILZpbRy4u99H7qS8rNkHT7GueJhXSV1
DutviRJhamimrETOLdpgySFK6XUV+bZfQmAX7Q6cAnhhZ1rGBTOEuOxiCZrjZsmr
xlkXPki+RUqVDJcqGEAnYovPLA5qQakJFoCvGPaV2IKkTUw1gll3EvLinWt5GPib
KyEQ4gcHZOOmJ1+PKniXgbZFSr9ooMCWIQjYuQD+wZddte+fcz/2Mlw8S4ztNl+Z
lhYqlKq+jD8u/0LXSR9MAGcxibNqCPY+O0hqAfMtzjxiPJWAuy7oc/rstt1kdFJQ
Ndrjeujd3rvnx5iZda6V7magKPXAxm1PR5RF6qN2ZpnsOUFBthzB19E82JR1T1Bv
XqMB0I1FkXpQK2CzuHYXFa2uXsHEn0ebZVeNKAfj4Rp4lzmiisMpgQirz4h9AxJR
ZDkP9pHo5tFQPO5rypQfXQtaqQC9JNIqrMQ++wm9fgL+HxvqBi3p7GEOHweEHZjY
Ysi4zIeRhUc59kYIBjBU4SaD/cGibvzF+57RaydOKsv6DsWVfV42FKbOS86gaG6K
sARixro4HOTPHb4SwoTmn2IiNSxO/dWb2EwTRwbTVNe8LvkYbs77ZN9bj4y2V9rf
9+m2AocJ82idYa02cUA7U1pzeBmnEYXBPv7GrzkF3oLbKnS7k/0LGHlOsFrmlH6e
8omkpoIqaCA8c5VtTAGztwXWBFwKaNmCUqmzIFlzQIk9j87JSkvZzCrt2ZkOVYBC
QO0GtSRfmwMPjTWc05AeDJLOIt4pqU+vDrshR1S29NWwAlE9bbva1I7U4BjnBJqN
8JD6zGYPX5KsmfrtHjCEFNTYbCdD5VvVWRpn0vPUK2vNJHbT/LbjwI/5PNxb0+Bt
v6X6RTrjqE8j1qn53Kc6z1yt/M6bcCH/7NZYgknaxa0FkV+bBj8b6JvbSGks5JeY
AfUnFPTbXBWwIdpWIsJypXsCJSeRbPIioUcSzbkO4FSMw3xlJDUMHFDog+WUkWDy
P1EQsQpA+rI6zRX870vbN+5MvvLcFZ/EYo1XE9EU9b27r0KugjJx/weccCjX6zMQ
4JLunxZGjLaLeOEgFH1MfZgNbhAG7ZOp1bIRH2BA54z/+gL0wAnXE9U61H53TCWs
yOLySu/NoCC+ynQzS/nxVQXFyGnu1brLL+0RorwR7KN3RJoUmnR6WjKSnPd16dR+
QFgUsfodDWPyRrOMXyI4Ed+J+WyUZt/fJjO+QeG5GoaaL8qFIVQ68VnH997lhdO9
+Mo+QDr+YvpEHwh1X+2loZLz9d52vwpqWmNBKECyF39yu1OhV4yT86LHp0xpVBLH
cSj+pobPL14rJKr1B0Lc+S5/6NWbl9YaTZ37xC1ej+CdWoqXwI2xVEJ5+XwPUxbt
I9wBy5+QzyL1diSovrZNoUWfNorD92CWXjCN1vmSmZgxzi7FIdhdSuY1X1vtyvoD
bssLFPtW+Os7J8lsHe2dnNYM+Uk92VbUv0bdN1y6saTnupFpM58/879xz810QZC7
3rUOEQ2x55dMCPl4OG78k6OyTq0nV6afJ7KQ2WFzU1nEieHJdrS/YayXzT5whsbX
+/kF0jDI2Mu9sbA0ZK79bXP9NC8KI0XNxPAKl31ExZmRutT+KuUKSXYYDFwi0fOz
qrm6KmXIxmvo8PTWG9Nz17PCnt5u88/IuK2n2tONOn1CfMDOAU2g8VzII6dmzur8
2sv+ElqePO1/rWLstUaiESW0JcKe7PEzgf2+gvKyg/JoPh44OwKSu1jmr6KetFXc
QOBBkq4O6spW2YYWPN93ZpqDK97oTkIyxEu4puHbQtlhaNVUpTD9g0+5etr0vzuz
z8Erk+UxzxHgOrFSI4ZwiJHoN2QEXcWT8nkMee/r0P3VI51lWMSEcktwrasP8GAv
Uz4jI/ps/UEQmbjMWFCsVNXsUROxFQZo0AHSFTUqfHwxAKItq8ECCFkq7KkrxxQZ
uGEyWrKg8Ny3dpK5AaweNUdroABOxEjDMCU+W2QWkBSmTWzII+S5xkAroMTum9e7
Rg3kOV4Yq2x21PbGCZbGmQ1rJCFeRMW3gO9OO4REibtExJqYHUBbLAaDiRDXL2cQ
dX+9DCkBEW/nPLJn+rGYbsoPFLR/bD27o6Moa98fSmkjfVrJ6SvxlZ6lN3bWroGc
0Tgq2pcLb0G28I7ilhZ8Aq7BIUzqsEXvjGvCFBQLjFDaC4IabZgOm+SlcFQvhT7h
rJ1YeM1CkpafW+bpxJDwkMofGOOnPWQg6c1p5FpnyIgmH8oKNyCo5F0PEBhPq2eZ
FOcL1cJUC9kiBqqrFtLtKN6KqadXL3kWPz4w4FbxmRQRVeMiG0yKaJDEsfaLwaSO
nO4awTCMylriYGkz4C47xjl81qAq6rT6puHJqpRbNHMiCQHf9jUHeTJMJEvTxxD4
e4M936gNPk4BQuL+10EwQZQfWO2bDEIfP+HxQnT6eLwkzTnbd6T8Yrr4JC5G8JlA
obQ78xAAF+MtopKYUmWha1pxvUZPvz735tHH7MluB6zAO+AHNiwjvhLR1wkHSgTP
8AwQ+V0tnTK3eYYjLyzCo2+Qvc0/LgYHY+LMmiHsGTuuHj2ZHDBr2e/ObiUlninq
KiS9zlHbAKFN99w6kS/9ydGvDtTSsNiqQFMU6eWPNRJirMgjzfGt/8YF94V7qeSe
cj+bPlAFlL0CHqaZ4MBs9HacW6lIyha7rEvKAhF7w8IUYhmZZ8vNbLHXnqEhsZ0P
7yDx16UU24oUQund2zE1aUuRItLj1hP6stZ8Frdq3DazHrA+z2ZWxBOWPLZ11ufx
kaFllDkJI2mgC8kcuggMc1ALiSKxh1cqEgYbRHp3F+n/by/gi20xizQ1w1ylyTDu
FW15cNzoTuPU+6kG1fO7ep+Jte0lZarEwC5a3gAb3/FYtmAyXHO0XjthwPA1XrDx
aUplJE9JlseoEua0iOq1EeIxTMNPKHZuBGJa6JSPGO+Z12MuqlDgR2MFj1ihSbAq
6ByB8UOppALBIW93w6NyPv3sNXjW9NkZrGxhSdtzMGPnN2OgUu+22Zvak13gcSXO
YkpXA7wSvFHyrrpY5tUbS/D4ml3tHYNHQ/FfQ/g6huIPXwVzgWg2OCnSgXCPgvAF
HiaCbheyJpXZYZZbX1CN9JSSToxN7Sh+g4noXdTdzI+X2q7hit2bOrxINMVwVewI
AOhtKI30QoeRaaDwmetfIx2lujfxrzRncIezNNzBWbHgSzcl6PFM3yl1d/c5vmYh
0N8SafBRv6e9aPw9Hb36VA20WO3DoCamST5O6ANqSlDBp1bcZxkxaEVwv9gHYRiy
1t0B5ff5rVnhMeC1QugBj+/x+/2JNLfVC+/4AnymniWTDqcpFtqBep1AsDnbhFUv
GJm3SKN3z77BP6ffuWVSnYqHNmNykf/87rgtyEJyLdgXJC95chc/XMCY6rU268IU
AGHmOhlz2y6AtrKJVNhm+0Jvx5pNBugReLC0YoKhWa460+HoTSvSbEC6M6ZfURJo
+0CzkKjrriNqd2qXkFajWqHdbkJT275nmf8H2CPghn+Th2I0JieAi8+DBHh9cQ1q
z2ldcId2dTCUUMtd4kZpEon+gmsHw8ncah69LBLqnznyKaL4j2Rt3AaLMPt0DXwI
Odk3tafjDvz5n2AkLpWkF0+DjaixbKf0wfnL0orjq/TlsFGa7ySsaaUPLcYAhA6l
zeaQsVyYcvR1ZCW4IuDTlbc71Qa6PLYUPTQOMtZDixjZPF1kLGUtBPFtIpUHNI1f
Uo6kKKIB7OamQ78oB3ZpNaxfQhyGFwh9WpsWdtQoabsIjmzvQvpVHf+Wlpyk39d7
Wy8jyfMb24APxk5I0pRE758Sfqr1/SqeuOwi39KjNlb4cFcDiZ/VDOHbAMWrlH7Z
2DBKQMnXbpaPXDMekSbRd+v8/MG7E4ndLBF8p5IxuUF8AQDDNQ/janlOStxnw/Cr
qSaPGOBDgy9erb62VJIJwFX7EXXlHVqwQFqJDj5tyH3lSO4bXGSgxPq8ynGHPT/X
jn3U7A7CZjAnbRkBeDIZXuuiO1b8bYA89m/Z16ldo927VfxMDHaQTHGq5Mq3G5Fk
ztKgJgMoHFgXLs+l1BhsTurEGGqcPp+hSW0sx/ifixVlJ2+6x7WXDl9geFIo2Hd4
C3Rn+Lg8ry5w71gEByxkfH8uMJIY1BR54UTky9eiWiFWOOqw/I+l5y4/tCypatXd
tifs4dY3Algeaxiww2jZwtjVmE23fPdaU1+pd4gOELKqIimKy6vVfDZECu8XcLcx
/UovuCTVKpQSDoHec9KGsdoKD5dladjCbHbh8r3TiLVn0QGphD6pl2gN9I/OTUoo
W2CsF0DkzXhIQLmdR2xHR/W5njW0A9HekpNmLFe7+7RbTNgZNKg1L8R5Rz6jTQDn
O6XskauENu3xTUnKCVHcPmAhkKzrA7YTjKRUclZ2moZmIRnLYCutz1DMpV6MpHyP
5Ie77vCv2nwbHmQHR6nOPRX21zRhzyOoPboyKCMO6jwXXX9qeS6f3CVOn2pY7Yqv
pJ0+LPvVMRVQtMTusLGDOqY0wNVla44FvKZSyibs26ZWFK9DOO0vZr40fbnKt7X2
8EfORvMrMcXLampSyZZIW4l9M4bWoxpieR7WOPlQAWbl9GgrF5rwSAhbaeFu6qhd
1x7EbWMjC7htopvCl7S75vGFXRZf0cA6Fh14cF4jmQXVLr/wBytln04l8caI7Ivv
wmSBiuABJpIUD65UQG0giUkrt+2AWHHd98x8zM0V7UvwUEv/7lURmPbb8IqaHz6e
FioWsvQ6CrRIpJXASL0qaZfDARi3Z8ouI9pi0kq7jsBdho1JSXhr/E/3qlJmwZ2p
3bYM77UKI2eHPmGqYTgf41Beketd/GgP22mpjwj+dIrjT/bwzBdsfdI6xrfNLurQ
2nG9HuNH19/IfftewfzsVS0lEh0x4Io2XyY/uM841UZS4YRol9qlXbwrvMLT2VS+
b01SrGzQQEMmi1GjH0IdVfPkiXeV5dIxioke6tmhj3YK54UX9vklA4zwvLMvoCcv
rFPSihfNLWH5Vx1Ckd+txShtdoFAb/lLwrz3BPht5JVmGuFbVDriFwgz/RJVsnJE
BVi5ypOAC4kuLn2fCDo7X9FxQnus/7IfzPIRVFlzav1sdwm+CQRHv49m8HSzV+x6
C5aYHV/ug/lDjW47lE2M4KAa025D3D2OR5vJ13+gyERpGPHJo1UGMrr+mE/0qnFW
eug57oBFpOnemhfAqUBVl34gi82KUIHBRPSXPog5/RXzzsSYL/TEv042RyFXrzpD
1kEdGYungzSWQBVtb6jo1N5YRvrKt+Yy3CyI51bDBg0LPbDM7OpqAmsG2p61iZTp
XLfPOLx5vGGBwGFDSg3N70rsOz/at2JaHi9KMIRMIjE5S2LPNjraaRznCjZTEESl
RlQDTNTDbKlcbMBTVV4Q2fV/2z1Wc+riBid9lpxtBf4pj87n72zbscZp/nv7OlUl
etyiox162+GelBhFymCY7AuKHan/zYL/aY2roMi+iLGorgyF037VWb6xBk+pLWjJ
uH3wvjyZtLI4bhxBh8ZLJ039d6FWVkobnVGeKIQ4Nox9uu/UU2d0bR1aRcSzAm4d
HRlSDrTjC0dG9zUrPTSmWlYtb/xt+LmzY5IRYftiLrqiNOX+feIYpplJDYRjAu5V
X4S13f2rMbztk8XDxq8Ijq0tHZNYIpp//+5kzC9CdPRCmxRT1Ytm2guBJaLjQ2ky
u3roveisUAHbwATtu7zA8UvCB2riPUE/NmKIhVaL9g4+ApkFW7S2SdYVF9S3acCz
saTg07ZBolb8d8C++IFTpcigwHZqoz2bXFxV3zwl1VimEltz0g2VaF1FicYp8I4W
IbaB1ALHu46/bIRat5OrOdB10sdFmjmo9s7HuBj8xPmwC8JLuup47Jo1ZF5BGzFp
8YpU9b0E8bf3v7pwokVNN3kHGsiDYe8v14yjkArsb/ORcBD6lNp2aW+NnpqEBLqv
g3jAZqzW1qZwYdjwydH0cHeV7Pzy0cW70KZzkTKanQCd5xnIul3nPRG/3viZUje9
y4QS1KTojy/H8FSaNLUMB63RQwYUAX98MX4FexU0IQolQWXu4nbFMLvSA8poGC0r
f7iktNdGgTgn/0MSz6WFbLmtQV4RdQ04cid7QC+Q5SINzXXTpBXSPztSW+c0PfR7
gF+LFdwKq1JRMIXD2EUXIm0+DtJLBTB8H91TseAJs7igf8BxUFhOO/ood/UlZeg8
ruqfcc6vHL1I38RTBGRoH3MHISxh9bXaNcNjaZb3myX2YBwdovXUKiMxxPRnJteH
84+JRMdvrbME94QSXvst4C+r4MJ/Av/5ibXqkKzjGTLHGikgShGwXF76pjmHyW95
zyVebObZlrHZi42/f1j4Di3CBdoOCWhSb3tq9qJVjhT44Hx9wfebp9GfwYNwPZY3
qzeTt4o4f6pa9mWyCANj+hWmZVsSFmsKwrtejJ82r9+tWpcVMP/gmgR2V60tlEmv
lnL4awlo6bRTlBLPLA2H892Pqlg4zaTY6LGyCDnhpse+xBPBQ7Po7etVN8VFLkSH
+enxe2uUoXlkssJj7SbvUs/kuJOTpfsOUMRDLm4OK2+6g7BaDbrhMxCEM6YWAy/9
1k99iAWS6a6Cq1caHf71gM4/v4zZocjr44Ed0fmkkaNbZvN/gbB5bBXUN6DCnO7N
4YDLHvQjzFPOkn03Fi5UcNlVtxhJIuHLChYw0U6xi2Vp53m0DpC1V2IW3jgQ2Q+z
uzp/8LesIMGKiXe90/khvw4RYsPr/WbbqZOOu2MVV4lZLo6XVdUTlOIlgrvXl3l1
HWN4cSwQjRm8SPFWOLMzxhf9BqNwGSKJ9PyhKuXIpBXWoNk7JVFMVyFyS39YP0ed
AJ9NnkTaYia2FbjCf1XjMjupl/NepZCdozZd8SaO84nrSUBp+d7CmS5I93soQOrS
sQwbwDfxfcK+A9XclkeeFZArSJ8ZhfJRB22WogBai3DEwKUMYbjp2Iw9dNQtdTYQ
sHUh8u+j+/uqZNJ41wkdvk4IVpNd+NsyM/FML4jj67CeCBsmYQDEU8Wcw2uYx+W9
EfHRFTxwBg/o8au2DMGiU0geRtLFrlompvHtdvOp7XYkiJJ/AZg83T6fJlnhb/Bv
arZG2i27ElyQzt9p9+ndv80sktPyGrwGKVoIXRHHTaps5+edtf/9VhA7Cv/eQXJv
kjkBE5A8oV7hd1fAzF5Cyaf6p/pMKGSzc8YIwucxwDROE4HqDEvejDclo0353/vj
wN6BFQYXEN6QOQv+xr0dficgzimDdQyCzXpwRKYDrmL2EgnEh5h/U+YpKZbjVoHm
FNsLbrDrcaaP7EG30a4F4MBXE2MT+qPKGzKPoEFoiIiNjCJD5/mLZapCX0eobdMd
VHAhrDXbDLJE4iC4YqHkVIR16xkw9a/PSPbmeLkVW71mdCxjQV99P3u5W4KGpPF6
cpWTlBYBB9RGWeKDCwCAId6It6KingN+HJiveOqQWc2RJhM984GZMt786yAX2WdS
Itfi28wAq85cLvwcHep7u5D+EpJPpvKzAMkWcbge2Z1XTzo90dUOwgxDFz0UtAl5
yWJznl7/6Yz1w75cSmJGHM35Um2ti5N6a2ToBJYxjjgTwVCPNiY9ZPBq4dDdDFF8
cLaovGm7BUjgfQVz5wbtLCFWn4LFbi9YKKOxhpO0jxgjFuhgjmyoUpjn9qEzYWfL
3n30YUNU80AD8teLw7QbjFxbTvtMRxOm8xEOI06YM/w7lyyM0GlazxAAdccj/nWN
MdMQ3tcIUBfJ02/iX5XAk9C8GrJR4DZ2ZGigpVBJuV09bDfHOm+9nlp6+X+Y4jGq
FqB7vhkt5x3BWTBd0dVVEqI/6TrsjffVv5TzcfStJR3dKtmsNkTgOSybxmoFV52e
V3e9onKB5Wn7RxCI2sWZcpXAsefjIJHyfsOaPVLc0JkUbXWLYwaLtEoQWb+XbK8i
zl+xuI2upxvam0N/u8Tsy8aSO9hSaDyFmUGjp/g8N4qDHOaIUKVxOuprqaq/ucGS
6OdVSHfCzUmEnffv4/d6qJhbSn05T3k+1yD1KjOP0IrdrjLAzCgdZ+1wkxMcwVmb
VJiFqsk0mZhPxfgqorVAe7GkviIbsTxknaQ04DFpFtoXbX2c7qvbvez8AuMwFLJA
8VlmJRV96auNmJES1qDETEa82BXO47HabYlwLwHkHEpbzaeXWApsAMzZEgqMSs89
zMNI3757YmdBAhWf3I2QzGcztGeufHasCjr6JmISm2XbOuJV5IYzOqi6LSCo4Bn9
JSlHwUa+jwrbpAy4TVmRKGCUMNFNisNJKoI64dziWL86sgvUWrKFlkTo+anakbIk
otG94xXvRc7wCx6Ouz8tpdlq69pZBEqFbt+QB1Lri/S/s2qdu13z4aMoSq/t+cq6
9QpxTKRfBJklwcwKaeLJfwGu/pUbT3M792qTh0FwME1/T2s3Qjma1shyWJNMXmXB
eCHCIxZRu3WLcHzowyN3F2Z8zn3wJDgWgHAtxOtOYfnkCqeP4XA4DKdTtCRtkJeD
8IDH/7BbDqRoX2m+UiuKA1WqU//h8Vc9A1KRbsLL0rg7ggwIp9xBg5vxHSlbF9YW
EBm4Ty4joV0xCDhP/irxH2Oeq+tBgL9KENUbmKzGpoB+WSq4Q6wJLPD5/Mlzef8M
4I1CTfMReovhsoux887BZrDCP/Yd8WRDRR076f1+9lNIpsHzuDr0vMieT5I6bA3U
IeeFqhQy0Q9ZyDgMFqvLeWf7teWg61QkkSlT2G53siXwnJ61kzP2NKEjE8DbLVSV
LsVr23kafbvncsJAMT7NLUkdZ6VVlzmad8lE0nmz52PKnBU7Q/kW99DvUc7Cc5bI
GU5jyta1Um/UJ9RxwMIO5LkavHhOIkTs00JFZLGn9u3UVJ+F/bO9hCzYD0XSjaz1
/ShUPShDiuQmwg37Aavs1iFPnSwypVphXsLR1qlKL3xlDLSVyvuKWvRrvWBfmhFT
eD5V/udEqIE7A6H1pv3rVsUgJa6TaNjo0wvK4cbjX0CNFsW+ASJHs/k3xqX/BYGh
yOXcQAlFrFXMFhueWutykeYj4mGAesQ1WOosD4O+cGq64ZoweOwljZBfhvupCoWa
Eb2DXk/bGs9tROYW5w+81adsVRbpnOGK/90BTfEU74H9e1C5RXjCiPB51IvcmJwZ
h4yk/TEPNhtxV253+rjX0WnQZHOAIEbA0SiHqNZsnpA3njfa6g9UI+uIGM0E3RDE
bA1cBpdouLGTxjZqv5Whk1SQZ4tzvFfHNBH8qOaAVwBdfz8XvuLDUKxY5m3MwcX8
YTxjQfXB1KTllfpEx4zP5TMgt1RcRxgUGinDpkOfK6q+xkMnyJv0KK25jcUPOu1J
Sl4M4C8sIBgm8XunlRcNAHqyUu8rrGen9FBCL3bWlCfxR+W3bXtda6gkqJJItReA
NfU6RMStetdmQK1tCUVEO+ES4Q2NrV1geW7l24uFnUCIp7b8KNAaEwwfPu+j3OCs
hBDnDSAcnfR/AihgM2cv2n1Jc1raQLRltutfvrDExL9CWy0xWVEdXh57Ejfp+M9G
RYf2/ROlrXIrgF0va24taaup19iJ7fwbCjm9ALDX2YF0PDd/+opPaKCJC5FkxGpP
4y2zmU0IQDPJgks/aJe8OFpK35wXOqO9vrhIcjPwxxDqkvaD89P1PnZ3lNaV8IGl
TUMeIrCXp60LZS9zS0j0kRznK49H9DCxrXkYOC3SHg313ZXkVb9oQdLsTa0DGRGb
KRJknIiPmQqoMCipKDqMN/ve5DHGkHF7ly59T2W37NkMqPeOeuVsyk0zLjWk2lDR
qW7L3eMdlR/s1IJAvzmSFdu/ZOzrAo1HTEWYDEY9pXEsjWiyNL3Criz5okprgmw6
OTh9dgXdiSdVasA6bCIJG6ZV1Bg7UUWlbPDilN8XPfk2OM8bvTffHM2I8XOOmpoM
KhnmxvHtNMgpogfxTfSNReAnsjTkDk+G4PyOIOxwTqSSdZwPZJkzJqTT6tAWWsrY
wXsCTWXkKdzmjJDbe7WHaPruz+gJhtyUYIgiQ+co+Fr2rOo7QYe5aRpVtJtL1cyR
6Uv5/dciLR1OaexMZBYtUFICldn5AIVhmKIh4sCkW5/HjoKfjCb3x9YdP2k8cm9S
ukGUgXKKq72AeksKlDlS8Fcao+Zv/MlbhtIfU+3/afWmLJuSqYmHJpb//Os1xsQQ
sLXmcdGFybA3K0mPX/GQm7lov5RnStKXjNnwLVHystMJ4DaFz87X0MfNArLzmaXy
YYg9lnamBGh06p/CJCgCsVTUJGEayGF5D+DT6Li2pxAaZ+Cs669OhhAL73PMRIXJ
M6ki34BNHzDtME4h3xvbOh4ObxNGTN/xRHmasUcIZI/lyDM++tmQfyy1eJjN9qsH
dV9G6BPIJwQxEO8nvfDVpSr+n5DMmfhjae1KhZlibw2yDnAFpib+edV8141j//8w
lhhcUGz86UqRbmeCdt8div4bKFrQ+6EJygxSYG8XCqwRkVb7wqytvTT3U6J4pAsM
Ia9JWTR8H4yyOqHQIdgFbIwnts2dHGjZOvih0AUboUSIQg4p9EsXKKSsBgdQ7sap
eMaL8fPDoouVhA6rGbct05lm1gnqQYgykpzvTdygR+hjj3sa1j4rXj5UkyxKFK09
F+f8LDrfG9Lg0tBw2H6EsRfJFeK9Yojl0hWkSnTU8FV7dH3ENk/2by4ZkREnSHj4
3n0JVojIuI20gXRNz3xR2GA3Uk9CG57WDGXUDF8TXv/t5sbc8OUXgdygrTJx9RK+
y2S3+xz1xATv5bBqpvJid0WdlEb9+hJevuwVlM8tXgFRk0YkrriDiMpj7o6HpFD7
XZAMr7IjdomXMd52qvtFcevzJAgv9IymMbWrQyvnvxZJiwuqQpeESLke0he43P3C
l8H1TYitAZu6MGGu+un3/j7yXqz7Hh0BjpsJ8lHTCPVvNvTgObOnXIMT0Lo223wr
dYQbeD5pu9AXOCNLaLk0ydscg60L7eM3V6Lc+D8jPe90WjHICHN17shkZBO/UgV7
7/rkblbjn+f0J5N7ocbY3DECpcXOzjFLzkjW2SVsIdTIjy3Lv2SCEZUaTUlVvO3T
3zL5uhh1yEyggjhIDgaXi3v6Mp8mSA5jUHlL3jms4mGHwL1+G21LEejK5axM+Sg7
XlqyhDEKxEsJunV3Rx7dvHImvVOGioBFM550MMR+/pZoXvXktqiQTm67jExuiXQz
4lknWZEF+o7M0uhniiso5nZlY+6p/CSaTqMhnkuNf5ufaexr9711b/yW8oQgW6QO
+ezrNUithPuZYVFXeBFxQFJyUcgzHbQP4LkU72OGgHDfTjDxPJaUzDF7jFiFS6ek
VyLe5nYTYPnsR3wSHsJjUDuRDMrS1CJWFgQIHnAlHM/RueYR0mEsQrAib4pdyZZU
KRq8V5Iui20E9H/PX6YrjiMd0C/fqjKVUCs/NuuiinE1H9e5EUBxxq5Kj+1Y+lbT
j6E3J4xElJKqIebNYB44MZyLCZcljWW3r9iEtDrzvSudXYxF4qk0+Xp3i/z7va7/
e4S2meotplzoYul967oabHi+A+HC7Vi7mrVOKMsk+BdymfBlGBau2oF5k4ISYZoA
feBA9+Hs6lnATKacpFEOlH7y6DEENptEJKr8SkZkpYFwqyeC3/zYgv97YD/zhKZZ
rUdo5gxtys9fc2j/Bo7DbRUyJOfCkYO50ojnAV24G3eobTKfTQfTYWrHc0JCeShi
dAnitJIs6/3QZIs/QHk+jJbGfFHaM9jlGD8DhUs1ZTjFw1cpVE99Lfe7Z+QQ3327
A1dpCoAwfX8vhSMKuGcK5cr2BQXY/5GwDhQrs10OFVVfheFT+yOo32oO5S2cV2TW
RoHd46UJqcyL8mmmZIDn+opn+akx25K6N3GXJqB5MeA9yrgpYGyiivZEvfD4CgX/
RsDg6hJ/iyKGGgng0T4PAd49T+aToO4oB/UXKOxTv7hD0v03TV7lYdZuMuc0Z2sm
CVmQiL8yyqlTnljZ9WVjfHVpiWDLLQX6L2EJRHHOA6ZCucF01IA8YZfGy2nNRLGE
n9Lgx4ANGfoCq1ejhYVsBmRrjKQcki673MqErkv7UcvHGuX8M9EmBUuHxmJKxEFq
QzEgemZqCuN9Oz7bpEOObltcv4o3Z+GCSSD4mVELHMgS/Qlkaa9ZAdgkGHcQLwYs
KfJZRIMAP5EuufH0pmsTEaHCANQChDR6/wFGUxaEcShI2iXxtsQpEWVAELIhLEHI
qS44upGJtNtuA8Ba1DZldkzpxV0tsyJl1800Z4iE1UUulzknrVeu1PIe5/RKVTOy
zKczS/1GnsYMkpG5x1oqejfDI+uTDKNpewgd82X/SjudPr4D/fN7z+4xi9DzAYnA
owoyaqCZsMIIEztOuE8DIzstvnqlrZYaRSuIAW60HBmHOqKM9T/TAUJWT6OQE4RM
RabKRyLSQDgDmo2xSjDgJsb+8IFnnR3DivwsyCti1d0Q/llYrTyHM4TrGRwd7nCv
vNj7ZavW8pwzUfb50hHWxAdS2O2Ey+6iaDJgOSh/SjdemM3S9O6u2NKjzTP40Fkz
hgj8pH7dVQwKwO7Q7ft+JU0V73YkYbqHcgkdXrfxr5MCMoRbkEwEeQygCjFYBzto
RifTIgn4csHXvz3v3xLf3oITYNq8lr5d3otC+DuJDCv8Qa7wiZsPE3LFNylpmGTw
qnS2hqK9Y0w1DHn+wJ9tuxA7N6ukK7cJhGswtN7QiJB9ICrYUwqNuib+nBrCLUD3
H+xQ/gNJcApmKNvYBaDT60vtsv5PG1sx1xmY2K0uYFJRwD7VhNHYcs/3aAgwbchS
tfMiIZ79RObwK02gBlKQa7InjGua1mGjHYvbfwxuqrnOVSIQxLf3f/zgho7j8kDE
AZjsfC9aq9k1Cxo1p9+VAxBiG2ekH+ONlH4R8K+QqxXXjzucenW28oE23oklbgNp
nPS6eoacayzTvROpZg6iuIQRBKAzcZG3oRO2NI7MtUOqk03ctx8rCF1RGeZayax9
mhsGAQbjX/shull97Run9B7hf3J3qmLST1ULAgN1FHxAe8NH5JReSrI2T8j2w6Fj
2tjrB65XR1oy6MBt5vQzK74+fWjTtITuy/j9LPfva0h/4fR9V/lfamcUy+8nj/vH
N4NSQpegsyKVXp5+sm57Nwm8ppvYHfan5/ZIXVbPg4OIf51gEN455k8eH5BkY4um
IOqm6h4jFtkKIL8TElmo2ooe+ChbXKK+2C9HqqXEsjew45YXyKgy+XGgU/dgjkPp
5wLvMzAaPW6t/EOrWUwP4CVY0V871nLqmbwB4CHG8TPrA0nTQIUTUsiGomeNtHPc
D0lbcZjsl+vF1JPsHSgOU2egaK3KHzPmJ9AMChV3GmAu900xWJ/2OCMorc2hTuy8
gOz4MMY0qTxgJ95TZ8MAQ6vT0mVFGfB7tMa/4wYhmIuJJq3nU2cMERB2SudEtVqE
xn3g2ySkbTXAVaKOu81KhY05hnEQ2Pxs/r2h8EiRHD2QIQMskJIAdamgX+Scs0bn
B4hnA6l3bqoU6lPdI6xJ7dHtK+FRVMB7NTK0HAescIX54znlv1j20ABoKeMJ6gg/
B+XIcIxned5F2U4LITEVEiBxYNebf4uC4Wq5bs9USRd/eQBVu0p4gFKtvHqvaZ9m
coX0ez8oEIh5Hn7ZJ46tzgZDkG56F5xY+VIuifz3ozqC4924Kv9q+8PDquxe3uLL
T9uIhUTVLfeT2ZXmaQx77ox6KILE7Jp8BpS6p0jWyg5HScPlxDPV4Vb1Tnp2nE9I
ejgkpE/PalEoNy1vk36aJ/U7/UYR9LfSSIRKQ9MfZEusIo2etOvrfhilGhDVQq+e
T2tMYklP5i4QKpIIvv6i25vXsaN8ipXN0gqUWbYD9hgQlMx6n00QoDygxohJ6Y0E
SLlWEE3Wj/jf9YzYebMQvgYziQUbSx0SS+snpZhrFP4uIfMSXXhUMSKw88gRGvLQ
wsMaD2kfvwypysvv1iJRNz8HOv0TQKV+kWhADQS4DaCqhjLgMIlZYuK9LKXjwFS5
mMdrkYUh2wFIO/bX9d+L7zbUQtPBQbmK0c3cTv9sgTZ25ZRddrcaT1yyQEi1sZiL
d1eS38sVj97PIZLDsFZRzn4d/oDzGl7LTnb5aA9g/reZHd3Dk5SNSpmXN6Qppdw9
02OcNduT2j/6xBxMoHhg6S10GmPTwZycCaHchocEb8u4z89W0GAirQS9BqCajABN
yh+d+PG1QuAF8gRIPWqERJ2E4sa5e400CJzai78GwXODDCDPXgkUDoYM/61lRhfs
/cjsu3kxcz1T52/xA+FX62GzIkT19ZMTl86bqIJHUC/KmUIMnw9vDSYmrmHKlRwk
fg6+H2pvJJRXGwECWwFXcQ2TaDiH8ZarCmp83jtQBT8kD0EsOGjraSm4enIoXijq
PsfkruZSjYDiriS7M8LelUvrL1U3C2uiGWxcqeFQi1mniYf4QYrhBEy9LeO2uFex
zcvYYsrYPeEXJ/nax0Qko00TCSt626gUJ25Gdh3nJnhlbUk8QGb/U9UI0+vKYAoh
cmXfpCsKj+KYzFJRP8fg5T8y4G6e6QN9uYZKIIvcITk8Oa6dl0+NQDEjXZjcTPLw
2Udx2fo/RMSVJvkO7YbhHeZ8g3KgZE/9aMtQT9DOF81amErghJd2eIYRBIhm3Nv4
XuCWl93oIhGWxIR4D6IcXTuf0D3gNxSLQLhUSDYTSQTcSEN5W0xVQYKfVXRaBWx/
eRcHQhUahoN5fzezu1hcw16acPI6lxF8jZN2B9gEPW/By5FyzuIqUDsKmn5Q63L5
B8MhB0dnIcPQLPatLASmf/EMKQvwLJ9RkCYNMU8VO5R34VfshWSpycaO7KhXdY+c
tMV2JRd0FtQNug0J+Ev2nnjgtpyHFRq3QFe3h1zNbO6UBpRLsbriR3QPCVAWKUGy
SREZlrE4e9nNRUspfUdYLkTbOPKHiiqBEorYTL/T0+0psZ2H9zR3x3MwQOvowYk2
sP00ZEr44p+OdIk7VRaZ9UsUYtGw9o1jNNa3Pv0jvPBuotBBCGvHykwgyUkSfc1n
OMyysnB/6cm+oD7v+mdU1ejazlV6i4LNuc7Ym9d9WbOqQZzbzuH48wY2OLje5xXQ
PyJ0mJeoQ6GBibdm6ZgwrB5rToFsBc3r+KlLvWUVf9/nqMGPODNd8GMl66CP9N+j
Vm3s5SWS4L1aAXs9WGHQG6GRaJRY6KB9NF7tmWhvV26nLmKyCf2ysfvNTt1CXFy+
TGVbWLkWhjA3LU2vT8OXNsYwWzOKCYdUdAt+PND1eqFRQ09FqUEvYkPpBTb3zfpC
Rz/0AmT37De+SYPkbhnQDzTMcEyHRDEt5KZHEqZmD9BKyrwDrX9wkN0vffhX5f+D
AlEyZF2tJ+/wbLN006QpGGqjJWN+67Yt5eGkVpBqAG5TxO1a/bN8+T78wfvDmrLk
IVbGTNsx9eqdkRLU/DJyq++N/GNf4MUxupBaHdMDa7QP9LejUJ4rBK/rmplh6JZq
zTSeSctypLgI7/QMQuPpkKROFwlES5YYoI9o43eivF/Q8q1N9zja5rL7FSO/iOUr
DDtVdVqp3Vntje9y22LfS4Qtb54EZtag+M9iUWj7bIcn63yqelqd4seqsiiAqfn2
bnJwM8NNZq8uPE0cKLOy+qwD8Y+sfUyKdHgw1MEcNUkHtWbWsnwJu7wSPpakmx3v
Y1v9xRqIoQ+r0VtHbLoq75iRM6wRqQj5Z4UIIXbZQ8LJMhXb6C3NBNTzLgBD8VVr
lrKyrZ5Vog4N7vXKERYydHKUPSartVso4mHWpION4QOlC7nYkyNdf8ZAskZWnWRG
obUnmDqsWyy7u9OYOVv0bwDw+rfVzkf93TAPmb37et0T5Okn1Us1q0N8FVreO7pU
N7PX2YYWYkYKYb9XrvsdprexUYvNXbhj9neYoFBsp468wK9H7YCNdEFqHKnBR8ss
ujlevQIZuuycPbVJOt4mvA7aI5w85MUOMEVTqdFmr8dj9OK43+kfekLYnJpMc3fp
saZvuwDgf5abcm5Qz/+YFd8E7BlE/5J+BT3bIRoAPG442DlrjqAzf9CX+ENtWDjX
yURCNSReImGCMgiRFA5sl13zFTOeIvq/nGRvul4C2ip5KUDq96002gTh/At5DrD8
fy1aXdKlG1IU/cp/OI+fcyzuUY1NXEKujKXEBOIj8VAVhVB1jf1ZaxF9MdVUSweY
1UDlA5tpchCcxTpuWHeNP4R/vPuKEBPUsHpzNjHFboO1zGGKx8FBFmJzo3xuwgcy
a0xepEKengDoml1zSwZ26VuW+NzCDBnu69BjnNaHsXxWPgVZ8MxLUqVZ8JL6uLHx
v6+oOQgxMV3XWEU611iA0rLrkJm6xt+HO9OHHK4Mx/w1FtFb1ngmo2q8aVOwFPkn
SrY+1yOMApUniX38fQ+UdAyKO0XUeOUHeEOVOr3O2n4n5DC4I2gR2VZcyjyHG67r
VzvJnTbowh1/aHnDWVKnu7eigzAUSIxw4OFCUOemF3EFtVVirGzdzA5VQS+daClr
BdOauzqyyNOh5qadFI1hJo+3F3J5q9J5AA5K3T6DLFkRqVveB7rh5POZKWz5USMo
2y3qzxd7Z2KL6rSJnCAWhpRui4FuCHA5yt4k9RLpf0nQzB5UbH64A8ZzihsLu81u
JkYXCtuJqxf+QNCfR/Q+BCqM3XhTqv/fKcbPJRAbAqLSmgPDm3Fk33uNmNlBBQE4
PdYAbSDzPxPI1zS1zXBq4Eny/SI4v8ydljikgk1U7aU88wX++6YLjsYntVlAXwrK
thsbl7dOCQ2mG1+4nZFtnRtmA0DZNrFeOp93NQcvtk1FdlYgJov3aeG3ftu0OK49
QaZN3qmr5VRAQGeWoIYnnPw6spsfTPBYmm/eZ4oEPXwGVIcEx8bRuvZZmGBs+LJG
YiE52rkhFEhKTxSAWGtn1BZBZfIXlbbGMtHhbc+Fr1/E10ZKHFNjFXz3x+IkkfsR
y0Y/i7iY6a3AzhYjb9oRrwQ8h4yftWrmfn3L6WHKxoLbjOgqY2EHBo2YLqD9P2t3
cPC9d+VJPow4BAAQmEspP7+LSLyr+xXg2+NkkimjTvS9QmjIMA5pzAdEQEboOrdW
7hV2HM8iK3hPsd4tPOvPt8hYMJdtAJUWjzWAZY1jfyEaRwFUH94Zho3qMj+72G2a
WMg1hUZ6+CUaLukGAZkS8AZUWgLPm1bwXbhhkG9ssKI33zfGyxTyP/zryWdKX3OR
CCNjZnXrlHlJ0PIOrLanYfMxvaMMnKl+hfhtQpy2nemxwJLZrSZxM9xomt9NuD7W
rdwCOcamjRfz8EoId4dotdb58ULX4nBWrwAK0H1SbfOtwEwPEyl+on1xXtFZGtwK
T/iNv2Qm98H26q1P3jMU7wcGhLt6ZWEiLr9+tWwnSCPijVAeVOWD/olUpNP4hvDb
N49pouOjQU36ptpvQsyrd+KO+kXRzi54+qVkwfCRH/0goILnu8BNM742FBzPLQ33
Q2sWtKwLZEBE4SxpvSVLJ9V+4KcxIMhy74urNT0alnOWwWXEICM80nZ/uvDl0iRC
lvH5qTc1eAcA2ZCfGgElWiwGa619Plcv5BcsBkSbI6l7oCfXpvv9lPuPKw5APeGw
vIzJM9uUBW0WUox4ZcQ2yS5aS7wMS6OWbCqamIXY2+IpEsoDxqA80hthabJU+VPB
PZKy40SECo3+UZwqSPiaKwOSZy5ZxAm8Fk66RHVr2lEJLI0GFasKx+lUIDGxysxw
huzHG+DgtnZZpbyMLL78gnSwoatIFjjkDftz3RoYF3OeX7VTEgfE/xdulaoVyxyS
zL9zHclceIx5hJcm3pjXRr2DyCb/reJzXg1PowM7UE5WPYt5hlVanDk+XrBPbvyA
bjRpZ5fg+hD2BxkIuyupWtWSBvepmNuVxgqFxn4jDfAUYc/u3+endjw/fAzctxIA
6z5UKsKdXTU6/Q+uSKkp6eKAvXito2vq9DvcNClnOYJ0M4Bw8zrFuXePnlInQwhd
b4vX2M0yMJyDeCTw/inDboKDnR//6crUAt35SOuumwef1vWsikRmFPIafxhC2nY6
Q8X0yii9KWENC8UzNXiPoD3rwfKvRFsaiP0E7Qimk1cSWIza+LBhp+GlqETe5GhY
SFj64PYuKueB8qC/AkTNiRf9C4ROby+m4Z3gzv6x8qxdgGRkBMCc0wuTXs27gL/p
4cgw87kS8KTpeVX9m+zAdG/BW+I5aN/826kU/U3e+XCqf0+D6tmQWA6WxYkyaFYu
Qlrtwbr7SGMvys9LVvEGdg4Xvugh7OsUb+1FEcCacYnTebAl+2vC+91afYpkV2bH
2sdXbC+dZP76JPBpqQ6rmesNgeK3fVnrqJAdmxoDp00I6yCipuOjHI1KRfNcgwn2
+XMvTSetwwMIPpzoV4kVSrqC59n+H5jrJrluFdvITPtczjJ/vxqaCQ19nHyTtolD
GYcOI+Tj3dBS87GUyCiW338Gdy5BGXfRryjaIkQZLCOUCbXtMxHFMd4n9L8fuusR
U+Vrt5OCSjc10iJIb2+F2GzhRPji1LYYo5O9iGqO6CbSDAmRnE5Jq9W7zFQlGQWt
TQNAUEcbDJIA9lG8vbZeLOMN90x9q9xaEhmiRKLErm+fqIoQd7l+ATnJeU+mJiKl
qvpNXLmmBksT/9+ogHfZNId1pPZvkB+CyhuEw4jS98tFFNkSjirEDMLyjEnJagBR
+pvDuC2mh+jUSg8C2OEvdrpO20KmRgvJcZ/Y64zvm2ftXGJpTWVdjavULgEzN3sy
ldww6yqZ/H+kdDWGnYIebQfQp93dnLiCY4NazxtUhBFs5MmzDwWbpAcZ1hLHRgdr
6Vl0czr9Z0GZBsDELfNmXdqzTkZZdnjUGpPMYJEMwQ9JW4LXD70QXmvtqQFdXEzr
OwhIuoTQlKRjxm7Vggi3PbclHVPfeWb8yT41hsXcAGd0IhiaDXZPK6mkWNq/cRcN
Lz8DcUAPrke4j62hpzycNqsZMcqehN7dHish7igqECVejrjtY1RSQ1SJAr4ZtU3k
MnaS8W7hoixw89g+oqbazvrOmhU50yHdN6z+KgtfhcoF03kce+XOFLGdmBx83uJl
vBQaowONaM9fI/WVu7j395r6lcB41Jhat07WflMH0eIP8SJsht+unSX4b8X2j4H7
TiI+0s5ybm2fYiTbjINNjjck4ulV9ZMkN6J9vU7maRDSK9gS9X0I2Zi66a9BM6wC
/akKHr/+nyEpS2NUkjzrmThsiQR2ZL8r6+nDDw4wOvsdlXZax3+FlRFSX4jDlmvj
pNmao15s9WQaCk/xoRHR41XFvO1KlAVgT+OmzBXyKu2olIQXpobKyX5oRKzHQZzx
gKbFlZp+BaJ2LSD5v/sYfyFHP7gyYO68YLD6XLzBe81/GufncQSsgyUj0RbfHgQX
/5mYM03K+XneXyYc+F1XdBtwZnDR+rCaG9YqWhmGJb0SBoYQFiKMINYhG4eeQ9XM
Kd4QwXckfpWbKRGbWNXanVmCHnGdyhEfoX6lmnoMFF5n/oiJkG4n7qsE0i7t6vTN
bKSI3yroUwWyhvLk6Iqbzcd1Feqd6mxz9AEhyVFqVd3O4tfEphUO9B8jnbeCWV5F
wu02Nc0zmYK0TNPAXf4YtGd4ZggIh89QGRVr+CcPPjaVi0A7cAZgVkku43Xe0B9R
zYfjFwy5RFpPHav+gP9vchY7ohkXDlpRSYwMKusv6dvmk0a4CgjI5nBNJMkLQDDb
IwAf+MmvtHyK2KK+VVvPKFsSxxeLo7mwpptkHloLWNuqL0UzqJr8yytcJuWwNRbg
h8JYry8lZK+qnzjw95jX6WqkspkXvatLJRDrZHczqSoodW/BhPfK8WG4NJIm5Wtq
nB5fjLP1awc5y10VMk8hufuSy/vndrLp3DgpX55GMaTxBsjhvQr8JZaIutspkVjC
GmKTsWtvy3BCz/Ku7JyJ5+izKl4FXL0WGkG9V2n+rTHYinJUWDYSxFN/iTDou1J9
Q4CsPW72KYmwryqzn2oZqBewBwywszxy4p9FS9g/CH6TxJgVn7CGoCU28kYiSo8l
0VzA/WcyQP0ooWwUHa41T4y+hIl5byTybDX3XeAV02Um/VghMdYSKPe6Gi01a+c4
TiIShXTfchq/d2LdMvVw24w8+5kirGV7xjo1+x0OSwgMbkbggN9YYQfTziWj+wj5
A+S2EVvQ9726WenDbutC5m7AuIejOBMLiF5U+qXaxmyrs9uSg3B+bUR5OET8i62m
ou0+mFWJXFnYOLZLRzjt0JUVXDyTCX4Lfe49VyGeiu1PbuKJWII7U5xvHfSprepF
7g3EboN5+9IOV2iRxko728bgaX+YFB8pHbBCL10wWUXq7xtn7DX4P/2lcKsm3Svq
K6dimR64Ap9KuOv7L5veGfFSVDOAQQ4Q6wPXx716nY/igCKhkIHyXSwpmHNWO3th
1WyAa7DdJBqhIGfAgGL39g7crxGPMnQxCvINe+VkIrwr/Zhlq7RSmX4tXMPRJfkF
a5g/r/hKd+cW0kocvKzKT8QlO33nri6Eec3/9FhJcCIFW+ZElAh2erO7K7bw2xnd
mWwVyizhvAYMWhiqWcCCIIDC2n0I6B3SfMEcrE//dorju8UPRio4G1UkAVVpbth8
qoEuvD3CGJl8wUQa1BvY7+KA7Kyv6jpJKdT6qfGMztjbFkQEEtIidPWLzz/pl5/f
5ADrrqJdpLW6OXG8Z5+YgeBHTYHQOmpwBlicTrwzqUdA7cPICu5IdmE78oLFLIVf
dduRC+B7el3YtXDz3hywNmxqmBSzOWjAZjBzMEd9OzLRhsekFwR/DcwP2D4YeM/5
06cdVYBqQTwWyaJ8/SmGgjNF7XtVQvWvn4JQB3Q/QKBv/VkB7NWNVeMHITbhkY6C
jh/quKEQkz0CEuZophEppRJ/SIakHlYtbF2gbOObU6Se2e7Gb0FPbrO9o+6gGns4
wPTvPa4B9U88MUwdTpmDJM8PsQAWC1wYwyvhr+lHFyY2z8RRstMwETFkhUZWiK0i
l1nIc/vqy5vT0UPE4NX3bSY+Q0wLk1zWtcaHNnEonBK6toHN/1/lsGNICAiwo/Kn
SFDd8ELQSgfsvpoN8z/N++TQHNvv0EmZ2DVy0S0voItdHdj8r9JvGNCbuAN8N+09
qOsIC4lML1+hxURtsasMFjiBgObopjWemLazRclYBmMQVVU2wepWHzTIo/ASz+Fh
rdAr1PJfkTFw0rGXCWcNy45IkHVxoFq+n/1jg0AG2cX0RuY9WsvQXgtn5FdB+5XY
HGGaSjeSKfkVKlaLa3lEukX1RHKfml1i702STMMZyY1naoraUMav+QfbtVjroJjF
rXlHaD+gaMhReMtnqyGthc+Q8ZjW3KRhatTzMnDoKaxNBjnNKBPKqdpce8HXNFER
uF9rWSy9eP5Vc1VtKsKtd+rcIkNv34Z+pmY/NzG2VGsJmUpQrpa3fd/SuQ9g+lsq
SuB3nKI8wivjcE60njt/YSgogZxbz6IjuYjOrU6Vooah1Yszj/DNnUgrKQsM8dD6
iY+7YBUfA1zP760ipXeuDH406n8ZyPemDWMFxoP3bi90UnAUzS+7Vh/6s+bUGNMw
u61829UqmfqYtzwiH+8i86cPPVoDXDXLfn0JJRceBeRbOj87qShTMpuKFk/a0hz/
VzLs1AXMWnccywXPu9VhzdEaa8HLRJd7AsOeeRDH7wacsltyiw+M4q1mQzNsgY5/
YhvX180UYjdoyVO8WBwnIS8P+K1JlmroP7ZEkoDXaYgfYwUBGLk7O7G1MQoH0VC2
iirdBV26iTD9yFz548xwoiCOn+DJAbz2HAmce2RjyYEL4MbZjkwF13Bgilo3jH8L
j/JVQ6f2jbirS1XXtItbz7hWYp4cpn2sdBZZKK3Z5WgtLrdLZrp1UbxsD18K6UGT
pc5QfbEXRuiH9eOmTqdpOFIoFgzwXOeZ3Yw4ZJgPHBaro8XIxufIbV4e+9HCGC9b
rC9YdMTeQZzg2JAj3+R4S7FMgk1yeQ0H6AZrshcFOV4kMqXPaDaqirCh4j3gGLay
oxuXTfCZhzs2c/VbA+BGT1xUamQFemm8CwxdqFQG71unemlJrJmEtnj0YBhkbsYr
U/DLz8tj8L4Zzf6QhBI8MeAxmoAYzJ5wKyhm17Qv+TJN2eC3TehpU7tIDbEUaJKR
u3dFm6YQj283X9uh/noJVF6zI5o5HtGfYg+7fPCR8UPZKcRlu/gZWMXgRkUUZyGi
HaU5V3KSt6O7XXoyme4oANe59kx17PJYvfPCuk5CYvexdiHAZ6XTwt4SXb7ctZh8
F1qYhJmIgU4CkxOqRsgm/el07Fd97CNrg89Mf48No4uRq8gVkR0zs79x3SQhouBi
0KiB2WwOtKs5GHp/sWD1+9eqHvq2o8+v4pBlJUAWysWYGBrAnMaZKO1FUgNbtQK0
v2gdzQhsD4OcA3PqZ+KQlIqHBrjuJmJtm+j4ZOEm38+hDvQCCH33PDIRCpGzs75u
y5bddvVDFPQgKzOCxgiX650IfX+vN5cSNm3cex53fDFuDTZXfEQMa8/u12xnAPEC
uPDIuUKq21XK6MNESmcarQVEJZXoZWMziosrMSKVNyc5hhIeg4QH5f40jAD9NxDY
jbRb04BqF4FWH3zoKr3JOaI/maxO9wiHgkfbgkr/QUuOIIl7ELfOz7z4IZYFJxDM
bW64GFu8Vv4drq7Jx1Uvq3husC5XkdYnwL1EPzQQHhJ2urtBKqeInlJ2YHggYNdo
OMHl1MU6XYK7yQ5X/gq1nC3TvbWtklln+KrLtYYRghXMOjJUxA3HKER7ppwoeuQF
LTSifXvSZnGq317QmuMRXUgQist4GKEOspmgCPTuoJa9y+jxc2Lu0CSA6D2+w91U
aJneTsVYlqjumpDc6prpYVUXIhswKlXb41wJtK88wp7VmpbrnWscCN1OWOco2hHl
Jd/BQkiW9833IMiuLQMF1jNSb5j7lvymwWIEcHkM6ue9Uq1RKFx0nR2ZQ3DdFhAu
l6vbWPCSQErHeEk7ylkK5acRsuQaJzdnMcHEFps0vqwDXPSyhRDiZR4/rPmkfEq9
YoIXU7J6XcGYyzI3zXIwheWHEeJENauUGsZPOeB2Jpx8hQyjE+BK2/mjet5LdcXW
Y9aAQNs7xD8mXwwyI/pqvXT2Z2QGUWmr8uxeAuDcK8WCbmgw+ciEWX83zBLKBQAK
W/b26lw5rEe0WR6cU9WKFKeIW8BidDJpnK6PN0aBkSxZ5ksBgdk1Kyjtwz9bjdyJ
F1mDYbD0uf+HLlmsJqb+L8JeRBSbbW53TNTPw1jNy5YTr7cv/q9xycN1fuPJZPI9
jqe8ucwKmKFXNl/9mdoSZIqMHoJ3gjtibEpwFM4JW3KpeDlgz6ftHrSsQ+F9vzaT
a7B/ZsQghIhGpDNQQrD8nfTGLGnk6cxiaTdWvRt+0Za4oxx+6oxE0uWOJrc3H2d7
sR1tcEfMG2RGdjQeWzTggWR8641dQpg6T3VHwC3Je38R7EwTQs53aF73HkzrMyRt
/V8xwpqHujgLU/FefyJ4Yr4l7dgcXmjv+lMxNWfsdkcOgROzhtgQb3VFGHx6wR3s
dl8Y/BgZ3g7wIGw4p1bz+klF61iBb8x2/FjCAlf/+Ze34zD56bgfN1yaommVN5vg
25uBwato2SjKRWiTnDETEPDh2T4JiXrAUxpXlsYiE9FmVsVREOFtd7wOSqQLvf90
n1N3rJIF3DumE8B341EfUZAqQ3mML4eGd2vkwrCCIg/vqSP5MGMZtvcITyZYLVSC
Vd1cfVgjGJaUEbcLtEDh3/XGdOjLDU/Ox9Yk20t4y9T+i0ST284SJaWrTW4/V1lS
1AvjcM5lo7XF4Mw8vT0Od/DkY5foEPDcs29pvhQKKem0AwJw8CiUiL5oddHALs4+
zA4X0XsHdbu+cFW5Cm5wBBP6HISYqOp66+xxpUEr36XUsmG+g+VjFGC4ZaoR/c7Z
twyWEqf0qZSaYvVSITC1iki0DbNmE7ho+Z4Tzj0Dl6e9oGyLMO501r/5FRyjp70y
MYvX0DUrEYaCoeeBdkcPjMccnwEVuRbwPR9lT0foVLtLjyclyXtwnPo5KoKjpRkj
FN4/3l8r0tAi5D4ez/1uBDYW4RaQmq+DLjkoKq27Yrega9q9cwqAJg295TaWRy3k
JwbuUa1gDEac3iHEkQi+jaNhLiwePpdnjrGACvtyDpoYNr5DVR7osm71RSkMCj69
NtpM7mFgYpkJ1CCL4QzSKkh1uteWHq9JxhrKxoqOnDek5SZqbjMsl7LQifVQFISr
0Gqf4e3NefzXscQheWeac2vSYZRltM/w1ojkMCCE7BQEvvcg41knRm0pRPTTMscN
qz3c8IOwJAKzYb5IV8/RwAdSgDvKD9PUaEaQTMTnSXSjmU8IIu2puTrtHCxY/uyH
/hD+klPfhfDUNj7PagjLZKxW8KZh8l/t2+VL3wjs+tQqcWqT0IGlyzl5EOlCqBo4
99kwFY7Wh3PwTKwY0nEt+v/JvbelC9vdSfMBr1WO8jq8XPxKzIEkBPJ9F/5pOd4i
8X4WwzJUdVwYjP8RVYNuCZyzcxbYiG6isPN1q5KjyEZeKOuUSLM0hkGPlQb3urNh
tMGDTjjxZIpp0NjN6k0mZfAnstUFZdgvqAT3r2d83UGakMKXzg7XwQwGhb8A8v2m
zPk+vaRR2OK1chNAk7YUuAbelw5XR/srGJC45i6mKTCvhgi9je7Y5JG4GI3DXY2h
pkozQMb8Lu5rgZwV/LjGTmv56n6N+IjCxLJpxptEOe4OVQPO/oWPyXJ/3r/FYwOw
W2D4oRtWe8ih5HiPH6x+6iERp7ip+Kjp/jPlq60wXHuPNKbWK4G7ge/1dp8vjpn3
y+5K35vP1dH9AgVd/keo0BTESeUp/qn5VlNpfj8i4JU0tJsaOQmnwo7LaGieOR37
jL/+MtZqQuffMNRzoJRIhT/8dbiSOJCHRBfkaKgKk+aTbCDyqtroN17mSBvYi6rh
W6jTzwXt2dr46+N8pa+E40iwqxZuWSmZd8Pw47GKI8QvNSfBUpE7zx/OpYJLH21P
hsvYsXubPpqGyQjkxIUbEWsVwvJ05acSnBoxNNXkBObvRnvXUrP73HmyDqjsnqaV
jPS4ozKML60rPklfcxFs3+It8ickeukBVKL2OteolKV7PvV7JeVvWfYHEjAr7+Jg
clv4dD9P/kwMhXQLtxrPbE/51uJ648EBkKjkjsHr6NHgKFC/aNRmkLCu4BZ9PSQx
+8DTAe7fKU5YJvcVyYcZJ2JBm8nZY+LBR8xV3R+/o097Ef8HOlyJpUekf0yb8AQ8
Ogzus8aOYLjxyczsayy8n+NK52nWdCV7Mup6US3cSyX9swDXPews81LTPUTODsgZ
EA4SOF0xbVfaGUxI1ktEpH5Hnfp6b/R7YNZvJH+y4fuiQ2s+5k2rCa5xcilShFpH
UJeBqqCeIGMDgc+LNcNyufQj7+sedw4M7rweDuNDJT7JX1QzBebjtt3YbgtYf+WC
a+BRc2ztLZ8rVvpdqrPsc2NLhBHJ8CEO86lnGbDDsTdlWqn/hOEhH2oNdYBdpZq9
0PjLp+En+QsHBbkNdxo8Z7vcypMV4kUwCfXEiFAnkoTvJhDQU5NryNtEemC3r7E5
Rfy8fG/3qJHUhuJG1b2klRV+pfrhvsT+dHTCG0eb0MVZvJDm4zHuveqfx3Sl/Jhy
+lV2K9B0ehRCc7EI9F/RYOW6lFtD8bSw3FWAWiZRJv+uVf6q8+gNejcp1jcj8f21
XXAaQy/zVZ7VdYRtGKZZwnvV4vFXRHAVyB7HbmV2BPGx/pEyyaU7qD1+ItqtSlG1
QzFXYhtMrufUWqNWMiyGoShbCruFSFsAqHH35y8C7hQwnofW02JqocmWr6p8aIrB
T3O4aZNgQ/VjPGEnu3pOfV1bqIJRKRx05SXW9ch4zNebJ4ss1FWdfoHwJu/dXKne
7fbdXwlK3TqGiPkPZfk/OYvVb1upD+LVaFO/doAHKJ8yX7b2ppnR+TygM6zaW1Pq
M4H6oeqKu89gFhSCRlSmGunaARurboBPzIldynW/vNrIJSlpFzO++A4MxWlJphkJ
As07ExeLbTu+TtKpguaKLH8TEEx1L9j3ID/Q65KsTtsPNNlbb3OArWP3L7f/Sdt7
K0YtSTieHhxplGoUMwP4iOduDoch5+vkCftWDsCPzF/G2xmRwIHedozOZ6fWztru
jX7alubHtr/N0xUyNXTFfgT+afiIV6TaZyaHop5Qh5rv349kDBQRdEM+p2CfNctt
+yR5pr2BdLJ7fzw1QFwMWmCPtm/pIpZ9Tn37awi9gUn/+L8PPEa6HYX0yWm704Ww
46MzIQCxuiae7ohpfPBtpAJcLWFgyd9t09usz3q5Pn18706NrYFWM6sOUincpXcD
h3y9ii58Y9Nlb1L23wEWajPM3sEvbdi2YA/UIn7jmq/5V/+g5QSP4LtvvxE+Qu0z
Fp/8RcpBleNoyGoWACYep7kv8+GgF1S5FRR4AmX18Pryvt52u8Lavpcp0mf08cZb
s+lM9HN92oUVCSIp6zcrusTTHfEEbOPbj702fdV8RbNuSqAx2UCkNU2Nx9xf5dYC
Flvx/5NQn6Z88Letki3yM9eD8cg0487B5IUcZJkmqXxSrlQfIF2y6/Ys98A0B7Nr
6vS03+j2/fiQcuK4t/tqICGIB4VxQzHpdcTi43RhuHtyGIxrID/mh2elKl0Id8va
5SPXqqOCZY9NrKM0uIeoiQF2usnvycWaEFsHStIk7/QQDddTGQMElYTzOnkcQ8QS
zAGSGihHhrdY2vjzO6xN6EZ/vZ4wr+EVFJPi54LEFY1OIAdkqsULjMV0zuMVdLYM
jwYE+Xz81LwgyZDSz62Zyrd1+V3sOLc8YskOvMVY6S53zzzSyNyUeQwpDlsWJmZ/
Jh1abCpN5litP8JqTGCeNKKAkYXmL+bEZmJrCcc4GwI6st8Hz5AmjZ7sbjWSOANt
VioAaipA7L4RkYZVF5GWLhGy8j+y32+lix8nRzIpex7D/2hUgSs3KeXcqwWO0RH+
o5pjln5AE207b/jPMDGjPuwX8E9KXlpscJA4+0Dkk+1K79UvxnzuiC6UHPX29JdZ
0kxPTpbZqVKeiwUfuWYoo2KHsXlf4RhyRT0NM+8byIgEVUkMxPrbQa5MasD/pSxd
UBV5PG92ji3iO5Du2mm3p40B/ZMC3XXBunoVm64OIj/RwJmT1isyjP7/4Wl7Mwad
a0kvyZpV27ToA666kDRhezSTGdftaPlPQ2L4VY8HEvgEefBCTk4XJTWt9JV0Q3dB
2aPzNTPWFGmqaN+ii89TglARCip1CeWAdvpRXADPJuxacgC8jQdtaqUjrf9Qxy5W
kYsjL5sqrhTVnmCEROXw51fKWfdljgNAewV729caMkvZRCuVEnPqI68WfvwQ7NAu
jmhmVnWLYSyTj0fPLYRi4yvLT1yFJVlZbnANAKMcZeuRtOWhCbHfmWYORsV9HXWq
2rG2M1OZgT7vZzJbGKFkdXGQeCHzdsFQcPIl+BYifi/GmIiPaj3hBfs6krGTgZI5
wq+5VdzC20vaKNCiKkrFHg74jc9pxfKyg7kxsAkxQU4mQJmqReSza3kWyz/FBvXl
+DFafVcL3tGOJ7pLK8crBnRKufxfFmgUuX3tnBbPLYk55hY/uPZR4D5nTNtOgRD7
aXiK+uepDRmU98aEy/lWOx8DgUUszLjJ2Pw2Nd9vP3sg4oJJcq7h8sgJwO79ScWj
5YrUzOEF/LCKig04YARuWDi8ufhTMGNWKEJmJ5WwNaWCHGLf+DEShhwkUnhZ+/9R
5Tv270AjBQWFM7Z8lmmEf+HXEvRB5zCMYFHjohUGepScXvKIiH/5jehB8hkw1aAa
rBNvJa5thdTnvKKfgXSvtCGBexuB1a0f5i/eGtGM2fnLLNBbuxNSrW7Zca9GofXa
3+nQhFZkUmC6BjQfnk4jEJG5d1lF+tenADjopZXInVB9MPEkuDjNeopwiRedZwiF
78rV0UEL5iINu/e2ZlI1qt7odYC96lGaHpdKsEchXRYGfJ0uOrCSuNkvECtrEzT+
RPwngkZ78gocAD+17pMUcmC4Pw8dNfcJ33wdyhGe41i5iWufz8iBIDlET8hu9BGI
ShJhP/pZj+833w45NNeO5MC1Rf16BdkmvB8l6vxU0ccy3LNODCrj4gNSvvgC6AH4
ib2XQk3MjpEDl/wTX0WaYRqWIXvg9u4bupgXzmjRl7eIv1fQ5bbgGqNv9/1BEsbE
Ihvlid0SzptRrBmnfvlhCUfQhxRaa24oaxoRn+KatYhy2xje1wAf8oFcx/uh/7m8
twI/DOKJorgVdM91WfnkxebRi44bhmqlgc+B7I0Pvd5DskGkv/w2iTmTaFpvMyNY
QWcBDhx0RLRaBy+xA1XyUz+ZAqXJvK9DZzdby674EBT/psaqW74+3oKZ8pMpT3zA
p9DZAI6u7zki0KH6Qfh/J/3KvQhy6N1gxxFEkDGghtYTn6eHn/VpOtKuRL1qHT7h
F67dDFLPiimgKaKNQ1SCbfKdGZJ55+lAhsr0a0YYMuEe87rkQyB8+Arqz8vBtEgu
nAuafmM2brdYaJtKGlOc0leokWT4Ojtn/B08uh29WrA9pwinMRxADbp8NEy4eq+r
f/xTvPghCq2ariw9mfnTbgSznir2jRYx1wsw2yWAl9ZDSqsGclvYl+noRwy6KMwf
lThKy/IEhQGgNxiL+EvE6iVeDezTvoQXjwtYiPihj/reE3kazNe2BS4ac0d38+a9
K9YMzpSKWIAw0vy4/Tdy/pPEnAJo6in7qjCXdo1VYkcHYgzO4xpDmo33O6l8Nwdt
sSSaTOw3fP4kiKsYJrayGtZbPkrj6RyAogvLjt4jDxMBoQKdZnlwxN4xQCMB3uIb
rQbx4u/2PZZcicAOu5AO0h/iJK3vjrc1jf2XE53BDQGY7YUMLcvNm4XyRBbiln83
dvhladxfyP7sQ2BAfH+Z2gt8TmkDqDoUvyVZCdT0uO0lfbZX4rStDHeA+vOA6Zk5
yNFRnKQHUwszLtcJAQ4xkOvFRjGCUGEsQliZzQ5KAyjNZOlljMJNic9Gg2nxkyq8
4t2qXYKFmhDwbOfDH7QVW5q2zmlKZeGw832baMbKuDXtzf53nZ5hTc/8Lv/mfZjx
AfiGG3C7JRM8NCwViuXe7b0OdbYnjC1TEiBH+Lr/uIYnWYmw2YFjGhuAvdbM7Fdn
9dpDQOrcDe1EFQJr7LaJtBEH1vkswLEUNFcgAgMP5iajJtjJUGMrZ75xepHESyzX
kn8VYZNh0qsQYoFK7fSNtitFS+ZEG4S8ebP6hTtsOkcXeBoAQ1lk2ueqrtjJZiKa
b9qN4c2bIXYA6HFG5vVmL8jCNaOhrQ9/fYBLo83jVGhzO3sBrCte1896AxAHKCW7
Zjzcf+4mZYqWNoDADUpmyA9Qw0TXHSAUXsk1T6dRlbbDXbt8wN1SJbSMZjUg67Lj
1Bm/LlYqItlRFQfffBjkR+vje8UdaBbgbD9m522suP7DNfeuI6viKu3pqYOHCwaY
J0UDTA3yvzBu5I1Kx52ZoyikmZ6Uwd36LWo6ncw2PBUm/wSdQgYZu+mdjIIj/Dth
dcsrTXjA1jCZtpgAITwqS7gwRgzCMTFTNVUZwjLyWvb1HtD5SmupWkwE5KbCnczs
6nV+QZg590lf5MmU5PoZdCforqpC/9PwY5LYh5KO3fiVZ3aNGOoV91yWi+3MkWUs
t3TlruQGc5DSGXYFs6trQiAVELp1A56YGcHGLBxo/IZczwJabQPrHBwXtUeip48P
gZGony+xWSOs+QGiP4L8fEm2ky+LrABM2ldN3gdbP/2SJPrLCb423GBR/Uqsas8H
d08n8+36S2L62KCrgQotwX75zHuHe4VrIrX+m18SZqKvKKbd6xExjBCnXH+UMaCd
WjjnB7Il9x/DCNp+V3CJ0aObsCV6VK1IqOcwYEhD+Af8o80FqZYB1hMQWcchdm2k
muEU7b8b6tHnxYsppb8suFB7rv51o4wKmfi8L9iJ/opNyIrIFGzHAIM6I89yYnMt
Q2JzZ7hmYNoQaMBvXmkWGFJisWJBk+ovg96+vEp4fAq1YHU7t0pIymTcBnSww4DS
/RjloZ2vvDh64Cl7FCGH1TD6ukta/Ala1RWIYop/MabySUXZTiyVc5y94HW0B8S5
8JwYrQLSmpJat8PVPQ9yk+8OGAY4bl59Ro1YDHbvSGsU1En8E8U8B6BxmWANU1zN
O2WX2H9du8mT27c63V+sJG1Y+YKuaH1p08UU8HU9nNGlB+vCuySHqdWGR/1xxk0D
k3YCZIEdFoz8gk3TV1KWelBdt9NhmoKYLCD6ANR25SKWOJ1ypUs9fU19zN/MWfaz
s0AtbIYjwlSNl5ekN0rZV4XHdO3Fo3j33Ki1Pqra3ec7NQG+v/w0HAaWH6Yuj1ST
Rlb/zD57/iDV9m35tI67ugGEAICZdbRruuRBLKdfy9xgJqWXAk7tqfWh7lyvNbrw
ARQymYsVZhY4DB0o0BjCa1Bg1w/y8NJLezzs0ZCexJ5UaK2u9jRknlGmeNlefcvI
Z3dJVdmK1MGBuf8U7b9DdsQtcwDuIylI8gbSk1VETAeKYmB1dboSlXQdKtfgPMA/
hSJuv81jAR36Pj1HC1SQT/9RlFxQAUshlYfflIhBgG56hnvfHU4iHCssZd5nYoFk
R8LV9M/xR1dhYj5GSkHTRGguXmIikV7X0+oTYuLPfIzKaKox6EeZvTeBt8MwbrYB
1M9SmqS/9NLwMJuNF047cY6jZJ+CI2cYnXGpu7ZjnuCMGfVY/OXFuVCHnt65xH1O
VE7YFwSurhHf22qO6M1HTeT6iD1LIEm1yYOBjUUuafivIitShxh4foQTJhYhexa7
ayY2QC9wnYbqFDIr/uB9ds1D+S96hT/QasXeDoBFewOXqV0w2lYFwwHKnUEEO1qQ
4qlAQ08y6KGdSO09yXV554WZ909IWS/bLEcsbK6O9y9QermG1k7UySiwQUc6urhX
EsRYq8pZfmxE1oQ/t+E9Zpm1VCcxytDXVtFoqSLS1dg4gY+xlCGDByv9jCxrM2d3
VXSp++PZ/Gj1XDv9cbwlZjG6/N4lAzL51zfrRNzYJs577Hz3soVlo232Zh5B5wfm
SvaBqaQDJj7osIdAO1KX0ti1tnwGq5Q0rmbB73i8xG9wtXvNiei5iAjx6K/nQfe7
VRm39uTbLDkWz6EYfHMDZxxMVT9BIL24y8cielNm78FJWq78i/8O9+354zlPG9Sr
s4bQnFXK94WRE03MZWNI/l39SkwxqAlksf3jB4BJDGQtksOfEWmARfd1TTE8QERM
mTcNOevqmy0nZOdUL4JTb026hLK03SyCycDZTxdhih06WkyyYsDfG5Rp8cUbKVmQ
PNqDLESPOxu0tMLiCKiL9JXE6/z3DRWJm1wwjEg7EHEHlnNwT7Z4ShowvNCWiaxd
1i/8pZrcpr0/8pNzHZZDnbJd9m6pPpToHliRBPxIcD+sVDndrhCj0Suy1qU6y2tc
jg60914gaKVZYsSznPRcNO2vchV28/WOe148Au2fDZ0WcPTBBYbRPqSg+BqiN6a2
qhAGRlSOwEQN3RHPHyqc+97GXibDTUrdNK6kzGWewPhTBxqXmROi4SxnuZ2xeafY
jWAnYaA38AeKy8QYcZXfmezmxe6M+GxZTVQwtPuoz5CLqByPQ6pG/u2TAVOHPX74
KCXX3HBp31Xi7BoscxUBdrivQDu4MyK7Yh1baKiOqVJj0U2Vz4rC7DB62cPZgHtQ
GOcpSE+z9v9gHPSuhjp0EcNKfyepWq8KCv4giuCPAJuqBoKasRaSGDKJ6744RkaN
/JNyvcru33pV9bK/vHEUSuMGClCogUm+QtlR+/0bzW550a/CkHE0NFmN5Qle6izA
Glr9+LTSe4WJOtRgQB+545C6lpPORTHbUjsmiWnaiGsLVpkt5o0kxjf40M4T+WdZ
a9GlQUFuc0rY2gECMyf7gOf182S++bQMn5QSRKVb+V7Al/3GPhCzbzVBwZKxOOBn
hg41DR3PxCGZBlF5OfzxCC4kJhUxuTIEDpCPeNWdr6lOzo8UdQfb6vIcs+pHwDbG
LVId9KV2gaP+xPfWmQKCY5/b19rydJgJv+rPP4plSEpV2YnNcb1dWNGtlxUo9pwK
VLRsyb/5n7l2wDdbQxv24bN+DuBBwvKAZgKIUv7Sn2JEce8eWUU2QFC81nqMv5kR
1UHuQidAZ+DWwTbjLK4VJo3gFRAcXD7hIeAhvEHpylXH95v3udLcLDn8KKLU5IEs
AfVXqpXVFxyb6WNqQRtCnqagKXKncrVHxAnwag6M7J5sOndJov9HAOkNAu6IBkJ7
iW5I0tvLvOGZ5km4kCP0iDt05HdYs9TABkXihQY/dMo5gdLC4pp0sxg/j8TJcpar
LGGFJz27t9u+OA6etfSwQLWQ4MPhrl69o3pORmXO9ATLlTGdsknGAtzzCT4kIOvn
ykwNZpyxUOF5o8iya0K2B2XZG8I1nkVzHj9qvHPiZfNKFzqA6FNiHFEg3Nt7gncp
Zw2sO4guKWIAgVGEr4D+8e5tcAaM4MSNMsNjtu8BX0cwESM4Q98BxCVoCQ/Ymp0e
Cj5JCoBQQG2eE5j5yjebWOl/opwAKJN0OcOn40b/reIH+pKGnQVo46yhy99EM7sq
Dpq0W8dxcAfc6GsI79Y5tHIhsQR1O1XiMpEzVTpdoA1TH0npQzQwEnTtHzfoN2OH
wBUKph6/5aTIMoNtlwAzEJRPbGKQS3TT8aIHrj1FH2SsFDV9IegyibX8Lbu0s3kf
6XpRHoHGvLGjAvpkf3yY7jYigABUoX7j8Y4lBs6KT6PJOE2bONotOXY2+hPECchX
PhjkEAnCEApxkz3/V6NJ3ts+58nR7/eY6l5Q3V5GLHCFJa9o3Mjyd7CqXWsRJQbq
yenOB+mkkyxwdDi1as23+Qp2eLagKIc1cpW1csrri/yOi9dV+bHOV/+Vmhy4hblR
7XCZsEokthSsdmL5HHU6ijEXgodV6H1Yi9OPKUx3Tq1mgGBA9QhZt0rz93g0XQAY
S7OIksJVrqrbLXbx2Bq7QF68sWW30zZZg/yJB+D2fahMRlrkDswoRHWsOI2PSrPl
5YtNE+TStFZd2ZgQiF2oVz52CGfW+K7aq8Ff500Y66vJPQBarRgDb/Uz8SQ2UmlV
ZXdWu0KYm01+h92jjVIvUS4weuMxZLckRlFzvIlnzdzf6aP9HZ7JSrfhAy4Y7DwL
xFtjLYARUVQOIATNT4w1U6nqmcAdfekIyTIKG31V4wIMwvwpgwH+P0ZYXmy75MJX
Xi2S7UfHGXKSOcuGkN8QOFIwMSidOhCvWZnF7K+QGQFjE7k0IIKtZq3gORpKF5RF
KAVpiLFO9VGMHu1x61+u/UHHshFCI1ObUkY7OfAgh/j/5cztcYnBKkj6LBIlAbe7
qVDb4ZIC8L/FIOLDdOwag3VfoqRfCxzGN0l/xGqwYosE6olx4Ta0L9oNk/7lbucO
QHS3eHD60ocTp0M2QF+/UtB0xP8LGcsTcczjCoXfYAnDX/jqwGDwC/uNA4ZN0RWB
806j5CJ0wn7wLXj4QCulUPGBD/4+SKAzfUBUMFnklVMp4G4HJ1NyCk1TCNaqeTP+
cUjaOsdShXcvmMqEBjXMUFHNVWKhnDevqnFgUKn3y7ety3l2xHwgX17w+FcHiF5b
3IKrJRXm2ocPeLgqu50utGzDZHp4YhmspA55KTWXl1aDpmVlTzamYgxGpvWOckH4
VwwjPvBH+oyxlSRwSwTT4nGbo2gxMZQPvN21NwPtKk7c+pARhxcxX5ixNXyYVPC/
l5o1CyZtY//6arWAdzMd4G6a+no4eHwb6qbLQiQetK8DpIDuyCJatJhhzQoNAtje
F/PoYhiS22J0x4UbAWiZs6vs/wJM0P+7RjyTwcT6v0V5n87KddfYC9nLVqEia6Lx
PLGjkb0jVj0BKWgVn1HxYfuiCcGjSaICxX2Swsl+4twGqUamDF8Li5hhB/th9RF9
NFexa2juKwaweC1xK9VINvchtyWpZxRxFVfhXOhg6ijPT75FFJmr6FYsJUo5ag3K
hJUIut1I3Vg6hRDZkuxD4HHPIHRm1LduITPPfKMSV8rhkrnCQhZk1HxuYw0Jq+bM
GcV9po3Vnh6mfEkyjnAozrDqSyYrvi4y/19bWFLC71XLzvfqt+ms5I55EPOm8Hiq
pX95BakdVezNTjHZVa91Zy2s3bgrTEZ8ITVRZU17F1guaPUimCjnOQ51TDmzXHl/
Lpv20rtrFgOzb0OXiIfhfbLGsDUKDXoxV2mysXLdbh+/B0zaf+/lK2YVRh796g10
9coECM91kQiQyQ+cdMEVK0+CjanMsRflAIqI26cgnIdX8gQPDS8qkUTrdswXbpJ4
5/0TR9Ec+Ra0+GNqK19LsKRM9G0u7gPysz425qdmWiBIRUT4oth6mm+DkkZfnz4v
cphBU+ewPVALodUHNCJCWuyQfi1j8CRNuLlhCcOUNKJNjOcajmB1aQJ7YIxX0xIx
dMhKTkRzlVG0rASZOxV76kuiin5Zsszu5XBFLcvHu7cmbu0Ck9ceulWvOWIjIAJ2
ljWmXYwtRQlLDRVb0V+lbJcwYO/FTqa10h3zddKzadJ2BnXEPoK1mwF0ZGZMkl/M
WBz1wFSQ+6HhJT0YbYXXvaPkCkIDiQZAmZqR3r60eF2fBwxAzVxFSVzxyOs30sMo
9qISXxZaguOvyopvppfv5DI9mkiCjlGg26VV3gos1eYT5lLpPxklQsZadheK2++G
yPP7Zf7IinrIC/uMQuzOmGs33uNUUbdRF56IBIJkWs6PJgnaLObr4BttE1MueUNo
rNNHoIK8V/ABD5lG+GdhzJGomomkYjuFtE0FmVmsZkP5yMU22dsJleLfW933COuN
qd21u37T8opQYw1vqCT6cGkXu7OCnSbnR9xQJAdeqRP+kOJm5JzkOQQbUj51ASXn
XvWyHtz3SYQMQQYPua7ktcEWu3MbBxaHiSASM3UJrfKjR4A/4DEh5fpiOrnnQL+r
ogcM0Ze/UCkLCjWjW8p6EPgqEXzNtMKgMPiOjLaDVBEmJqd+j5iE+sSz0ZU/R3xu
NOjn+8C1tVQtMp/jzDZ+sTfFnbpddkxEI2IO9jOnSEGYtEdI5KPVWrj3njTIruKS
rWG8gmLI5QjgsIaQ4nWTghF/ihFNq2j2uAynt5trJbL/4FB6kolDbUSXTdPPscKj
IPlsbdFD4VPnPRp34J4B5fI6soy/9BMtqFFa6Ynn40eStu93gtYUt0VhkcLyVr8b
16Rf+VgnQQVqnixmvWB/09dZEKHXTDSL4rONAqPbufhCc+cEXHwcBMLlmWgPnX8t
nf6qul8SHsbd2L68nll5Gsz+2xxu1UOz26FopAu/pQJNUFMsBtF7hM2Ls3Kz8/+z
x+Dtif7oC94kJIF62/LjDB+U7S+yXWXPuI3QuT3aiPTMIfd56mqSMLLR3SsicY6y
s3uOF/d8mzPznGkIJEcLMSH9PpFttCgVVhhF1A+Aa5PwIaTR2tWHGcRJp+s7a2d/
m2HDrC9/nEr3h8nbNYsrZAH6RygnMgbGj3yijbxQ9IRxbnse+racb7NkhNOtmO6W
GQOJ0qHl5SNRWxlcDj3vcsDmKp66z1Fdnmfls1eL1ebb6GiWg7HrmfsMLseDg731
mI4cHqVA+0sNipRE6lMmkBo/Pfi/WtdYAgzenHVDQzwLjTbzTGWVwnQoE6WJy3KM
Dp1ESzi0e5UXf6LTPyVVl/XPC9RIdr951gBG+zv5olMRnMB9KG9n5HDkZQ/jtol5
jSI7ZZIscwB1qdoC1BAgerr2pqZ/kYEekmpfFL4TC9iMz2T7fogPDUOTP17pr59P
N+qfoVbXu/wz88RkLR+PitU8my6sKmhDTF6FXaysEzvrmgrHMpo1+m4gVo0kFKE7
si7sE26NzC0xC/1ExR54/xycYFg1pAJS+gQ0F05zv0AmVYcq8JECLf7nd49oNdEz
J4h6p3H+jlgXNLf99xUwxtLoBr8AV7LHr+p6i3rsN+yVA/A3ePnatCRIOGaLqYXy
521+QFR/XVDbGotvzWaSjoGgWv77Yttn1PRznTR/0fLbLJE3U6zfmueC5ET70+3b
TktH1vXoLanowLlCqj+oi+k8Bxs2ezswZoM1253yOU7ZfC5O1Epl0f3bYxzkFL/m
o1+IX3hMWFUp56ydorW65GoANNJPxOX3CFwg1d1PUPrV8aUINqEkFdtIq5xymtLk
lY4dlMLhEZ7JN4eXDllqQbn4UTHXGlehnPU3m2G/Sa7hsq1K4/al2t/MnFPC3jzm
/FZ7FSbJXGspoxk4mgysWdy409tZLHhvPsPCR9RFcM/4UNFcWxAiRrYteZgqmMvW
BtXauMk5OnK573WXKqfqxOfIpWiSUUd4Plj0PuxafsQiM7PFSi74u6+AuKEUFZTv
vaRmnZ9l+ukzCORqyBWPi3ZTMoTGG3ZfZMP9bTkqg8yh09zm1nwwn9uabhQ9Pu/9
fOtdEingsuyvMvDd2g8yiyPWQacrVQCnEoowHjjNzLrcKJeDJx9qwwoTb8PKhYNe
L7qqza1MTft7Rh3UGQ/buP0fL+FLBg4yuPtz9drqkLfS7fKRoYl6CCkRN9WiGqFD
kt5chEwsss2qunlS/yLcuHhKOHgUKW2ZIas6HyD/fwdO3zlz/938ClxSyg8vtSYn
Hk2YZZl/5eXpQ+/weRipA0ATDmO/BwS6gYuAgkAXn8VDsm3T2k37YZWSBDZdf7rH
u6BTM08fio21sVK7W3n3+4UfF4pOXSqYsmp7qnPaRs3w6yYKpLgsiKsqn9QRu/i9
L5xt+hEuC8ZvHXTs6fQnC4yRv2sCe6Kp1cuPJ9fQpnY7xlWNVM9B+UlZbbsw699G
syfOTdq5+9HdvA7NFfJFEIPXNmrfMtUqUu6TOVSJwtFgpq0sMb4jYTAjqiH+XaZD
jxFiDbJtT1vN6WM4V8CbUyssCcXpc8ketiIY3CKr7qtRFkb9XCwe58Dz8c3Bk3jF
jaVymWo7LcCGtKEhkMahJk9+aRrJ5b0oY0ZCtPlPCcTN5ljiYhh416pYfoYotpr2
RJ9+0j5ZZhX+6gy7q9g9rGZ+BnE/C981bp+YBak+B5ox925wyMQpno3ofK7t9x/v
nBTWfPDXdos34xp0eEc/IM72QXf1XkjHw4pAYcdTc13ECaIOcLGUxcz0rHxoLtpV
1w6zPLORPXki8sv61ajMpTUbQUBUpUJk+H4bFPL63dslMpZEHWtWb4NwMoo0OnP2
b2oFV5/1laIKyyQD3UGfBG1hCBPwdMDthdyIlrwhhlipTQWikiKI+rPGhGrSYY8u
RWsmn5cUqzabQmt1ZAkShq5w1p9fI6fdatv15bJpxs379xLMF3por2PsOQaMgW1N
VF8sRs5Dv04j6GmqN+tpoNnehL841HRpcZhJBa6RFp88O4+WkPi+wxN1bRDZu+Fv
uZ7IVQME7o3UokRR/DATb3tbAuiJODk/TG9ZThNI2TAUzKKR91SK3oqA/V2/pY9d
qaKiqms9aot7+nVp04EfpVRZFvZn+izRUXGQCV0JzqDQewp8MKUrqQvFMwq5wqgG
Qzlht3p84Q+CKV2AVfnobz1fuhgeZR76QRp2Dt0UGo0YEt77FJjAvEOP/ycKqrnr
CQspzGQBxtoLpF/Nw/s4g4zoli47mCYnKAcD1xNipbeuyO4aIWT2Ix/jAaQQ5SmS
cBdLCwgV64Gaild3QxKV1skNqAXETPljLUbdeEsR0cGIXw4oApyyMr88LzO1BFcq
YGVfirv2RGEvjHEaYinXyFZYcJKWkreTWhDh89txEGm6EhOATKAfydl4smoRt/1R
8FzODuEOZO6vw4aNgNhPx4wLts76EZkWCe7QcxKizYjAjig4Oc4GXXwvO79VDakQ
bf7uAZKKS98nxqbdTBJ/8BUldtYCNrGG5PaMNECQEwBBw4NBo312RAiqPfDPFUw2
byNg5hAPPM8KC79NSb8W53AOIDh57RF/lTsnv3QeJ6ckfIALqv2MFfFaT8iW2mCc
754bNBWwzlGIfHTMCQ/H93fmn6Ep+FSQeagIJnyULG6Cjm6Ts1ODK1G2zuGdFNfx
Z9euS+QpRF0OC6/YuaGmrl5st+AE4Ix/YtTwBlagyW5DTg7mnQxUR61VqFmJ7d/m
O8lplNLzgrE65QK6xERi9Sh5Xzvaz3uu60XTsnBKXtM5h1P6sEllqiC9a4Dd1i0Z
qDkIUqsE/Ryl20R4HMwWdqn26qu2PGIVqTgFDBXDnpQMM82qcqHotFZPw/DUq31Z
1oanetjCrZuDu42WdmH/TP3LcZeez8Ye1f0LmZcl8hV/VJuFUTSo5uuAJPaObPoJ
hw17gdPHjysspfWxHv9vG8rzuqYa3ei0G8HOcjQ4xeo/0adaE578UreYDpPgmCiT
KZ2cbFEK8dbeej3GBbeaqL+omiUeiOCHdQMqkPuDsDogW84W6ARcdqMjumppvmdU
2CcWCzI0Bz5ABWfJtPIocz3od5BV+BUxFs3BLhT8EEY1ZBPWF4DrffV4JAuj4LcI
1zngQ2Rqze/HhEfxHtwlOwGJu+0D6AVjDYsuj0dp3w422SsSc34MAjalZZySFne2
78exgsvUSKbuYPaOfT6jpKBH4LNSHioM2PYcZ3o4c+g802oBGDC7b769yqd1lZHr
R3NuJTKGVwnjQuvBkzBKPGZPPNo+vwDrWY/8c6CN2iyv6bDNRcLy6duCnw1Fg7Qj
rVmFw8BD5rl7ilgRN0Z683zwdj7lGkUQVBj2efUG71ihdpxinFsEopP5r1WInHjy
HQEK7OGz1Bu3oYW3gWj8hGQUB155AwCUh8H15J+EdcrVxpj+2rIkFzcbZUJVuX5D
2ZYbCfhlagFf+GOHBfRP2NnwqB03wYAF23eBuayD5yZgCtlJgXHWwAKkGzTF9RAe
fxbh+9XlO/bmwBIDx9gRd8Sg30WmUU/s3ax2zNFh2R3mFXqJWmqpQQXCMj8lg7hz
CBO/yb8SLF4ejEtqv1tDSbGtPJd7MCEcu4zazKbkKvF97f7wnPy6qaYYAIHBoxHb
ELJxxbI/75XVWj/dJwVsc6BQhmJd7NLzaDAREbe2AxsVEkqACMsYdtCY22Cd5fJH
118AkyGNCrgKhsi8bzQNApVEhd0e5hi5s2SO7RlbcOlfJ/h6a73wSikTP+0pCQe2
eQ95JaOMUt1dDmGcgLghr9Yt9rwW7Yisqs2I2jNcQd4ILylMNQvg5x/1e9J/TCgi
GvQfsCzAO6OJNxSEeRKviUROySDmehm05oBkVCtqSqUhMlUVJ80VYYaa+xVHLgmc
287y5q0M1EYKTViPA5rDqK4qBugv8sb5x/rNnoZloTysZYEHe6TTmWtxsn7BcI7z
BseRV951X1UGbGhlHxJqPf8Q1mpjnzXLkks7sD1Nz1lPM/K93jqMRs84ee7cQzrI
g0ytEEMdisTJBmYCKumoxEPce/sk/b0SgLmxn0xVqI1RFM7oRbZORJz4Nt3kjRFl
4zCzpUljI5UjkSPrD7DGrO/ujvfOvEE/tr9QrHkn/c+NszUF29t1AAOlT+fMVyP6
5q9eAe+k9WbgJwnVlH4FMFOB6iLNRJGKUDvgWiKGRh9bZjR8b5T3Lo/K1t5co9iG
C82Tb6a0mhKWyojLkqHnmSapacvZplS69H2B+dEppAazX4QOWSQM96ppds97RKim
9Z3QGv+SF59HydhU6MhLwR2xor13i6PeIeiz1W7c/JbVyhEKqgNfVjMoJiES8E/n
F7fXo82JY5Y3MxbhnTKZAUuBVunbZtcn87QEDKIp1qZyHrrKbJKVoXohYHqjuPt9
zBbXbXgAAOiANakkR2OBwvTYDmvoex4J3NjipbcvHQb1EXF4o1W14K5Y81Mngwh4
jkR6M9lGQfTCndm0z8UeWAguWK97ar4wPDyb8dR4EiwicVaarakW4jX6QDi0mOoi
HinchNrEa52Oj83RwWjIq9vycTw59SYJi9VJ46wadKd8EsDLPo/dhf81VYqSUl0+
6uPzcfvIik1B9yQ20PeTTGjT20/nN/vrxqL83hRAQzgfQRwszWuN/56fCUWGtQLV
oLIwNz3jmqjxkNEUElEDVleuE9ZBPrRu6reGZR7RoKm6UjzDZ88qwRzF/LP1dM8y
8HhNzFEXC0XfSL9L8glne+9mI9Goz4szm0OA7Ar/QsT3JIGYRrYOeaS+rJlUP3YR
r1PqJzuzeNBtQ5RokcFFnHPWW2sm9LkWEufAKcnDBEw7zZHUFgHW/K2vSV9DU6hT
eyw3xQZpGrzQ5RSGD2pVPmveS+1376v4hPMkhdThZxB5eiUtfsNYYH+TBdVKgkDF
YlU3DgalwIfcfm15vuC+LljpamGENso8PJ1O1WrnW3/U1q+4yi7IjJQx0hXSh81i
g1XLQaPSY74P+Ntyuo3BY9stPth4unPufIWaZFDcUPr/0RMbaWTo0PDkFr+ywUxy
qPRd91B12r4+FHDLkif6FVYmiy3x4jgsMLXLiTBSbp1KeH0pE+d+SKqvphTRVuhP
CDpAW4ulhqyrzXUIytxokt7DPbL3qREFvoA/xqZ/ZSiLLNlSWlUASwh6EN+uxNvx
7ImojYIQCUQ3ryfW1L5Ly38X7t8K3I+IL3yzAGHE+tK8jF2FFiromc8Z6MFcPxnI
9nCECsI7i42WkSP5QUNpB5Q3IP/Z5FUbLOYmZm7Gay7KYRWt6OsDXJeIQp5s7d2E
HlVF5JZgTJhYuUhFfWhRWDNhadejtW9aDShlLEw7rgwdub84PCxACN4s8Qngggkf
YWX1pmZaUPTW9SQgctMihwmv5sQE3ARpsMyf/QAoizLVSYIE/0CjckSFxQcrIOgr
+9BDh9kRUEBX5iLgjuwsZDwiczf5/MxsiF0UrJfbf0OYtUlmplDtMGx13gzsWQz3
H2KeiHwMDVe3lrEdgMvfFMnyl93YLwhnxD6P9mTFtDF4djk8cAwEAZeZvqJ82yov
7IbsFbqESOMO3YEWMEi2V+6PEVCfHQEboQ9TpoWo3vD0d0N58QWWkFO5mXyJFAui
MogkeeUXsP3hKI44aoahzbYq/eJzOd85NGxcFUDmB4moEELjACDMR9OXaro7wu7B
EoR9l3aVxWSOnxS/Y4XBUGukal3VAbGK9b9HIQgi0di+PkepalZ18rMRtkB+7Qp1
cOrDkpZgoiWuXFhx+Zb4+QnuAt2HsRIXNC1FynVxCBthJWMUb7Sj9KApN8vZ/vsm
B+R172HVvRZeIoq+Hn9aP9HZxU0C+pTsGg66DwqDQ0g5bUdAh7BL+lA4clcVzL4f
VxXS4hqBJB9GdXf4A/ntOScur+5kLFarbtCtSC8LZBpxJZDuQ6pxZcAGUpo5G4HN
+kOGdX2xWk8arc2sh43GYlTDIVuBracs9Kh7l9R4vu5xFk5aUDKyJmWNnVQlAKyW
GS6qncJdlYcVZcFVGTjePAfP5LxJ5lepHoodlWQNtlyG71C559cW6Mt0lkYFXFnD
JaeywG2UJ474fbIWo/YzLdW5nKuOeviOIlRTV8tYLYp5H7LY3ewAPQv0zfa6Af0/
vMWRYbMNeKARVPzgrWXHlQz+4/PQdKroGZTCJNJNwWBhhsZrcrFvaTFqWuCArHRN
td9CpCAYiHF9+93+caaaGen8d3jh9USJ3TPPFd83m7p5ObOvltz8641a2DJCGIT+
JYbeBlUSjdcTSnEPro0lo1Sg4XCYDiqDKYwn19Rgha9mYfZbaYPrk0RnhyKmkwtO
WaixBqnsBx8d+9uBAhT1Uw9sB+lf8VxhsIvEkTzz3cmiHZk8x3kk3bM8yGD9OGMB
IPjUbFeF7EYEN02Ldqrhq88qO2O4BnYFpcn1xBGEQu3PVrkzP5oDVZIhsy4hRDlD
rVwePrMkHMyQB1dLHVR1urhm+xBRmNlLUK4v6nvd8p4Oxrlv+tK3HAfp2FbktZ1G
SsBF9/UMgowCilP6RJD5dunIBkUyDuVp99F9o+v9qUXka7keP7xLi/Gd8HS9jzQH
nsTaik9Y1G6pwlf9kVMl43wuOsl/UGD8CPY79GQRfcW8Bs3FjojHzV7h83oQYjDT
rNSxFo70eIl6LZfi2EF0/rE4xSRD0/hO6xMqQ1wbO6bUy5F0airAU3Ozkz3hiDSJ
NoF/on/Lq4jR9STY/BwnjUviPdoQiUeeEW2iFaigDbP+2V1KElptKIpLcbMC+ohu
Dv8syHCKNPfy32PQP0Wp2rmGfOFr6s/lj2rvZ5VH5GB3o6Yg4jbueO4uHQioCB3X
NlNInG+4Z4a1gWkSM1wJAXfI4rEH701tkQU7c4wqi0EcP5zmGZGTlPTUs6AHtE3V
XAEe9X383eOxoY69gqwK26DhVKbHLmbPNm+NYlcz/zvLAwbru+ItE7hfD9KNWKqL
Rjq1DgVf+lsQ3rgDY3Ezrilv0rzFPgspuNfRIITU+KupjEtehpq7LS1xGKP3K82b
5FZ/YUo9Chy47yA6XLZkTDCJ5xNnROew8a1tDFF4b0taQHEuj04NuqnzClUR7coU
tzoKmPvmc6QPHNqVDS1RFO+vuzTL94OAu4GkKRKO/dvA0RZwgmWUBqFBcdTV3yHw
NfDk3WxC3krUd1Bnr/1y60nAN0eHGLMzbNbC5932XcRm0OOwFsmGOwS9v7JzU5gU
qsHrGEn8Y9ViMR4X+Ef5Gf1dBmlAInczgC28MzXxg1ak5Jt8YKGPAHXc5tQmS/QO
bz0n93N5bofuydOqjA4bhO+hVqXuzcERjd1PROXbRNE//cd4+y94fFboxNPPxyqK
DyMqN+QWMWaxCGyY4Ul8p9qWdw4oM29TTJtRHOwfXd4V0ZufVJkvzk92GYCzi77C
xXQGvxE7ruxpcnF2V9G6qDRecXCyBtFbjby6LEYglXc4qhdfGy0TQUuvCL8fRnNs
DA1tY2W0NNGre4q/EWl7xSTKbwOSOSWkTOENDh980r/5AhxGIa/3M4I+xkIX6rCx
IAa9ih+zLPc4GYGEJ66jqU2CNyM3kNcBHpEZMnYNTCH6Bsp3mcnBdvZ1fVlQj1+H
ar7Tu/xPkhOWRZYh4rlLte8TbZPrDP+G8fiTFlL39PO0J1u4V+QWQmHdvHfMzjzZ
i6RZJquKPzjXE3EkF9fjv1aaFf7/U4hVmMgZ0zRIT88EaivhVkKcTF6L/kG8qdLF
UrJS8yjH5UN20TEiEoVHnC/MGdWz3j5lkJ+zcN2EU3QPKyGPd++xH6EaeKm95Bsw
H0fSCt4XYrfvhh4Bk1IVN+X83LXq+e1NTj+aB0mBfV5BHXQ4VK48f/p1YX6J8ZAV
2fQy5Qokw5hlD9D9K3mIipPgaPuWegDwHLM0wAdSDuwHw/+P1ILgAFNDIQ70SZGp
QK6wUfn+GL3X9eNoK47dKyJAFqCuHRdAnU/NvPlXWlMeUrV5ieOF/humTjpinFjZ
xRUWvDBC+0Ua2o8qY+ZpGW/oWdEBU3CHSW3rQGHhXaX14BVKM4OYoLrFGdI3TVBv
M+L9HgWCTvMg9xleKtA+gaRlvzxTD0f/Fnm9vXNxAAlMl8svUIOVUfFsc6hyaAwz
116OJwhrhZuXOZ3CIDDxTFIoT16MDodiZ5TPTk0tVthLgV8znCyppissSuFhVk5G
D1tvS/P6tCX0llTPTXZoT/004/ZYXce/CpezP9CT4HHkkdQ5ZU7KhIAUvJbZOM92
FErgLKSwkaa5GfSpE8Ycm6eqF4L2fqFHOkj4oDMVPbVAfGggm7NIlzMQc3a+vW4U
lRYy8sVA+yqByZ+RYTj54bCIhRoHnyTPkCDqW28bhLG4EmZrcQ2zRDSt5WPTLHhe
yV2r6P6focudj+ux3w7Tg3bVFKD9WQQfw0v3uMdyJFbb6QZkMLGSskuHcxTDB3ul
SCstHbYAdWg1h/oyWzSMd5hr85f7jYYMBkZKfjUl25WEFXj4zpC6zo7YvE0yKst0
2NJ1WFbk2O0gP1+5Hni8pSElHoyRr5JaWZUUYLuDCjj0zh22i1OBg2hACT5rG70O
NFmm52T99gRjIBFGxP9Bwgmgmv0FxseYqzwzZzKf946WsEV7N9/LadgBr/xmZwqc
u6hmi0ocDnRlcO4/PDl8ZOblRZ/HsxTJsSwIyb5ZnBFZIFDDyx8o7imnuEL+jPkc
kkCEnazaB0yBaISyfOztzU++pHMYMTcIWw+QD2UMHOONlqmG6u3nwkfG9EY2J946
QfYQv1aCBQGIkTKie9ME2uuN6jROAYDgEzDyJZHHI6yzirFS30oBjzNklNue98eZ
fyrQghTPw0Dq0e16yVWwmow7194ivQnJzABkPCPq2dGJ29vfCzrKE2RG1uHoZ8oO
7ww5oEkruY0v8IRlc3EvDggK9YBthhW+xOuPTbA66YTYeJdqcyvjPgYjFiiBbWpv
LTyCs+pVb9ghwYQ++HL7MvAcP2ldi4UvNm1uPSfoyAGt8IIYgwiKhUBl72kn1lMO
hjuJwOTCpLPYoUIbGdNcklv2fbRyqw1I9NVbyBCWBkr+YGxTvKa/nzKxI5dKO/dK
9+wF0SknALfuRn1o4JPsZFKdgveJHQmJIpkBS+8Q6lvlrkrkd5kzqktW8OBAA5mY
Tq1LVKMD7xSpIVytD4sbj4Q8l1LiUWLWhaYqsMtESHDbLF5wrD0G8Dvk+TzeT9G5
8a9g+08JSG7+XRTjArOyMc71p+cEBxBEETF7YkMAXWtFdMfrokizgm3x6hLVn/6Z
7PELWebaYl7gE5ihOkUU/aDy9+ukyuXGnEd9nUhcg7KwJyUVJFKsWSVG/iOTBDCW
L/j3Y3HKtbLAnb0WllJiUqVs34rtSKnV1ZIhFU7lZNkKzwxrQmn5q0qGjIKFYrM0
C6Nrqnc8gDpjmq7K436TJ0mmDhsbg2gJAArJsw72oJJIWbSlSQWHUPMtXa5o/2+Y
AvHHkQkj0S2TERNdrq7FhoQNlTl+yX9DrSRoyD5OBP5/vNegoBi+rWUx+4/UKvsD
ekFUAV4l+FMzMbYuo+190/75ZjYy87e1zosygdIM8quZHowvcS51t5v4uuRShP/Z
4swI+V6JWQvIfR9zcYMOiYw5iAiCx4O5BLQhqmHx4PC0Zf9v9pQ8qhvyc7zGjvl6
xjGqm8uF0nkqAXpAY2ggIitrWomc51N766/Ze2u/s7rVYRCWUd8PRZaCp9JB4tf7
vXMD3UDy++38QtpoWU5X20hvn2NMUFMlQERldxF/Eg33dlhGF4TX4Z6bXqfOhNhl
wu3ZZr60uN9yskHNMI5tJ7zOtSYjb4X9ZQRI6Hsnf0Me4EzPRDuLDPqKQR83WK0C
3EvS0spktlmseFpeFmvhoXZ5uhYbqqpXh++4MP6tHdzIVvkJA2vOVWaQgRkNRnXQ
ywM1vRFtA1Q0eDo1wBsZxLg/tsBeeZfeBJELzAADVzC2HGW/eSpCeigVUuKWM6LN
75Oi6F0+TrNzU2biIHdy1AsAY72dES2fEjj6yofTJbbDXbEGCxrSTaPWH4Md1BcD
/mIoBvO4Bf8mI/KGmeBOiCz0EFk2Ka0M3aD2foKZhv9KLBOLkwIDTB4FHd2r6K8C
CJBL/CzJxVU4ncMtFl2thN9dHmCPia5UhDrIiOAg2TW0F2ax+x0qWeNh2cSmJb/Y
CafVNzuyxAD7EYeAq9uayjq/6DqAk8Nu2N68/lvE5VT5K4I6GWs2zo99Wq9MGMpi
hxGs1e2+NhIrhjdsr+Gxq/KSD1VtQM+tyIkS09oshAMCeEmT210H9AkIq6QJzQvC
PL02vJQ5C91Y1y4stu8l2sG314+n6KWkXGXSxpFwqOynOO2Sjp0imIeHAJORbA9y
2flLN+PX/SjoWds2piKHSeOtGmbB/FhWboV9FocJh0NoBZ7vcy38fiUcTllwuos0
V6GxFiZ57J1k2XGQdzd3r/icC7Vkv/yZE38Q+gUcTheNU5uCY/k73DsOijp/ZeLN
LgHhBiznziDsnvpzT5otri+C9m24yGBHSkVfOAiaM4R0jNe8fPqDJ9YSCzZIJ1zO
CfVRmT79DnLKeeEM40OG7Rr5TsnP3XxOQN6EzgS2JFjJTH9sk3GqnYAWNV3sStD2
2AcFFavsIuB8tNQ2sJiJK1dCEAT9C0ziJ3pP29VoVY/3gyyY3/tGXUyc8pR3Wl6i
JCEm+iXxU3M2GNqrHGgb2lE+8BSYy+CHNiXMOnKAO+q7dHxFhTzl8UPCz3+yvZA/
7bq/BKyOG435v8A+kquvHnmA6Z5Cw767G3TIt8vMrObOBRuJBdawLFIQ2Sm8BWb6
RBhi9pGkam4EhWE8mXNCL4xdNFg4BCf3fw264PzQloxexn1bcVpRhWTbRqMwljWQ
lMH/qegjzSrD/41AzpjJywFueXx+wI6eKUdXZonpsYu4txJXEv6Ov44aWf5ByTrw
pegE48i/0JgexJDa6ttKl8X8I/eeEnPnWgbrSgAwtiqf+0/So3zvaruFChKkYubF
llMxJCP7HJbc1OdS9uqaU1WoCAt7BVb1EJdBH6xVnGDt1b3GdYgG9AQyobs5NJOm
sEUjPZus1M2o8K+5lmlmgpFb+Aml9BmJcLYS/WxtMXQc3d2g2LB4VNWGCatkn9e6
MOeIGZWpo8MtovA14X277OMMqSK65/86V/3Dcnz1h1xkyU/9LOJlTuuSKzhXDjmh
O9o9wqaHVDkXavCD6m+qS7mWD5GHjhQe65L9TRepRfLpd1e0GKoEn20i4Oy404gh
qlVfD6DfLSIVIrq2APnzbCuAxWjvfgKsDmDfiY1WqGFLvWhT/2UNDiwyQwg0Ky0O
xoB86MQe1bIUbLymBhaEsLS4K/AfI6t+TlTcPWfsBjXLqYxA+F7J7lKFXeMNxsMP
x+jx7o5pZBBcrb6KcChekD0nt/XlbYfNKb6JlJvxqI5JZED9m1xSvebDrR6v3SM/
gRAer3jMIvhemiSmuvvrft4zk8MNGycsd6VchJAgSULOT8s2KPJoA3HZirW8pQYl
yqFSpREmcyEIIQr6r+Vg+hcjblRUBn6eWPd/df59h24pEHcr2OnzH4ed3sxTMYph
kCR002443GQjAKmcmm6hvUnFFu35eBlO2fMsgfqw5S2bV3NodRhIoApcPGnz4suG
Bjv12u+9PeSqZDiqmdX/9iw6mGnI1XPyZeyedeFRTYJ+3zazss95W6ilnkCpfApw
e3c939Qgl0bn+7jXZQ/2VmcpK8SS0kPLkeTfaofFAm4rZDRGMDQJBTng8uj++7Dr
hQqCqfVyvSyZN3q5g+BZSJlJGtPXTj1Ofrt7HZMuldOxjryP6mhRpFIsSXmhxhkW
EaL/CeBbLOlgPtqkNIqcDql3QOeJog2MHKc2poq+eVPBUrDuwxDJyxGERJHXjilo
AMsLic9oOt0D+UxRh+XPi3OtiSmNNhlwYJH/iPr8BMTJh9L49yd2iEShJ/YuktZ1
8fsGvczbwjNIhz8X7r1qn54Ia3Hh5RaaOy4VuuDulzGr+Vz/yt4R/UfO0sXKd7R7
GyiPB/DDd+SOTDSrr0ZZ7xuUvkFq2Cvu8JkoKJhExk3tfKtfQPxSTv0k+K4iE4zO
p3/51Qe02wZADrMI6v4Kaf9NKHwR3P/F/oSNaNiSByGDN+7Jl2gl8PRRrKiiaP0G
ogmHvvP4j4GvOP6yoZDW2p8hVHyGqJKUUwV1adZKI8rLyEMC2jzlX6bYenmM9gGy
yJDFiq8y3JrA8fdcD2e6UOZTZhq2s0wHiISY7yGc+5OIml220IHUjhg5FeVIACt7
XkwXKUn47RZCLDBfwpcSo3cLDGzveCJUwAMo9pGgb4lp19W+6//FoK/xDDfqnaDQ
U++TB6wk48SYBcKVeQbA559BSh/USCBgOENQuK4Q6GOW76z6d6DBQRY+j/6k5Jmw
qD1hDCtpHg7kPV8YQWK2JFKOpwjRJrTENQWo1tMLqUi7eV8MGXTY5FWZGZe4o4yc
AHeb8hfi0yZDdXBpVmenF3yR44CpBRKMwzZFEHxwzx7EEqeBUI3BmhK7Yb20qOWQ
MMXFpCpcxL849eEOsUlRFHt9Kh+1fGbhLG/i20012dhLjVGf80lfXT6NCtXB6iHK
CaZS8ePzIiSGYz7Bw62UR5VUMGctg/VVPmIeBRo7H+v+vmr0Bb7QgOpkO/MppoKy
fX4jOsDNyZdc2WJPRmQqQsTNbwPghgd1xAr98kQT8nPiGqJ269d6Hy8ZPbV49fW1
7LfB3Upen6uz85nJekkGTOf0IiEbGfwD/n0iLJr56e3xsAKbA1iBRfEsfD4OGFUS
oUyundN6OiTaSHt3jKjrwR2DR4ZkkE8VZgR7TOkRIkGEKh2AkjbQsfLSn6NYz2tu
DJxx4gYPxixM5uB8IvV5eU5l6mdo3iP0J2w1/9HIsJ5S5Gp/s8RvPlbg7qJz3/Zr
h71R1u0rdwR+eS4VBeTgKcGT/fubKcbfltcJRY2DrOGvGrqnhlaKgjII35R3kRLm
cyELtiIPomYuhj4hnXf4RF8capuhK9yVp6N85y4GgC7NHFxhw3OjBp6wp6ZdE1uq
V7P7hnBKHXkPyd6bb+DvJTwsDqwIQ8YaXMdJaAYtL4OLnOKn6K8qwUuPYD4f3eh9
fCexfLGK02PbPQNCIT1saFowTbRgV0dyoexTLsF93pdQ8aX8wCOeN/58vL5ILeCW
voqQR7ZaaXQazNjz30ZgSJJm70QXwvGWzERdiNRCmD4=
`protect END_PROTECTED
