`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9EZ7RT442dJ7ScQrEPg/x2x1qh/nQ9n3zml0eYzORZZOY1RmVvzXoArlAj4MYyQz
bYqDfXhcJw6oXK6dlcrdK/g9vIJfkN9nQnGxWwvETWZCaHSmWArefSER/K2JOHoI
EleiVfefzvOXVblZn/ixtCXBrfVGwQ13qv1VrKWSo9wsanrXrloZbp1lkpjWRW8K
45t2Wl2k2ujVefSaEDRXRk6tlN0R5J0aLKu83G7ZgtSSmdBGu1MKKCWSgYXNjJLu
Rcyqfz5h+/ME9WR4Dm5EtHiagD3ze73YbFyXzNH11yuSrw2FnTZ1UsLv9V2dI94d
BJeas1Do9RDCJeU5G3PLJe54QTwYJvBnUZTtz2XGSVr0YolyNW4KSSjY5A41IJwl
Y93eKM8dYtTGCLRJEIU4aMDBS4q7Jqcx6kGWY7F4tu+MKmR9fqC7CEYFd17T/LN1
Nzw+i5jykE8O9UKXpl1lUokmRuwY47n0iZwygxPjB6xiPF/YyZzgdDC7Gno6GXLl
KxfTOceE19prp6dUrapg84thkPlrSzRQWb43sIBRx/PadjmAMp/ORdArsak/49EW
JW/KY924fS8jypFz4w7cL5jSD3+euF5AV8uub2eClBnEbqvEd/MnrcSVbZnSpcny
y/ptobXPmAzFepNwxgloMDdkGClpKmK35y9+kl26qZwA419e9fMjCkVopTMVydKH
fy8NkGe8QVnySF92ZrWlr6XUXF1Tz/HROQdhY7vQfxeqNhfvZdx6078+EQe+yK2l
Asnf+ArSXCBe5Iv2rahcPrJ4Qm9VO5qTuja0JmaS3Coq2VnUIw40FmKhnT2YTRe8
qfS/X1C79Bnc3FAYjoJ2atgjp5svIEcUyiOLiY3HMLW0/zc8xVSw2X8aDpo4tNFq
hReNDxgsA9w3Zf4BeFozf6w4iYzjnmX+7PvKN3NFcta0envmRiNIOyhKF+wnXXxU
nOnMQVLUw23WpB/aMhSF3Aa40XWRPS/7R8YOzIp2lyMlrPCIpKOJZl1N3Gkgnn7H
VWceNaN7LN1XPyAD72ksSePIyODUEdDUxJZmTa8OM1e4n7FZNSLqI031YIx7051l
aijB8YXXHjF2gCmnHV3gPkrzYs8JPcVp2d6rlcehH9h0cfzz2nqcPREvKjYKY+AZ
FpN+3VRAD8OtQ31MQzK7bBwaBdDh0q12P/58IFIhH+FCcRHeEKrrW3UxmPB47rP7
oswtTnnHXmea5oaDYCuI7aRQ8Ic4b6s8DmFwNqCrJEqudqD5F3YhfabEsMZwvNyM
D6/jnuT0L8I7F+ozykXATkZUDaZ2QcMHWuO251j30p06OYr2hBKqB5Gx/8wdrydA
xAN+1b/XmGg1lpRpjmVahsCQQmqY5MVdEIDGVz7Ds5DdBJ7evhdc4WZHv2ZA2HWd
S36tATsDBjMub4kRQW1qh/COPY2IpESy4MLAqcfaJnJkKG45sggoWUVSDYC2ofc6
5ILrC8quITbD/dvqwQZLsR9Wt8E3XemEuh0I4xrJbKqFczvq0v3b8zomf9pF38wF
vfTJENf5p/KD1om0lbQoGpM+Jm9dEiovmc8qbYItKIvMuuP67jG0APyUz7T6NRoC
escahNk8u2/ZhYlH/MlWkYyw2YOm0DKRR5RfaE9fNpaT4yf8WQ/1dzL91KoXtTVc
QOCjMRRvkptTFQ4J+ponZPMn/G56Pxg4JWOTkeMAZdDJlvf46NzNSU4sY4BojHbA
cmpOBncjDpdxWI29cNEAsDIAWIy24RQWnVdQhH77zPGeSzavHfCUEMfRpIlFFa3l
dRdC7L892P6fq/hUQY4MzGaL+b2//IO3nJvQ4kHOdmESAuYylYb00PAYOLtMzwP5
kw6XL3alI/rG0awnpqMwdNgDqugTG7r/yaVHtzMN7MdWsulmUtFflu5dlSGgtnJ/
Hce91EcaEMuUSu1twRUU7b/uD+KrkzFcCLGipXsB5hx1IqYgDOpE+cHNN1OdBgBY
N/t92WEsO4v7JLoPMDgWilao+l/HyP1TyBJWE1VkLNC7LXskgv7Ssa74boXJbJKI
Er9FdwaldaYG851JVgAOO/5Yuyx0Hy5NYDTp1uqLzLwmjojuOiehfwdRR/uMHap2
pKsK05jKNu25pt/uQDjfRJrwezCc0fygJFpwjPuEfWSqnC6vwHbEu+Qu+0KIbo9c
W+1kE7Uu/0YtlJi+dqew7/ABZ8OL7+wQgM+Nc5PZ5PlKN5Vo60/HKx2XctmlP+nf
8NDoh5AKbm1OY8QlaY0Q+Y5TDF5V9Xy3SWyvDqhqudIBvzvEBK9xBsMlAPuTuPtw
5PfyL/W0Xa6aKYdou5BxJzk9jsmQOMJdVw0ClSZwBmd1zYtp9oiYXBCcnYviKi8f
0ezdqUcFAJ2cg0TIVmJW9WJv0/RiiLShvXkNfEkVxvhahdHUO42lL5LUlApdXMim
jER4GJljneSIHrjDUyK9ZGP7HeLKubsBp7KmojqfxhL02dHfkX5/Lr/uzkuK9YMp
ms8nuKwZepcvLY7vvnrd1A571QDncstN+A6MXXZTHSk=
`protect END_PROTECTED
