`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pKtSKFh3AlqgDPrt6OSVjTb5altZB0dY35ZJCXuxMnGTH1hWKd4PyLpE7g0fczcS
NMa6Eh+EixeEC0B0IMOjqVPNgxznTtDsa7B+PbAMBwRo5vYxlcsrHjhhqBd6QDBR
UbE9KHkFVJznpjyQJgeo3O4kONwzsPefrrIZuiozrZWGGDtPiP+oyZX4tcspMjMh
M9A+MsoWu+r09dV/83u3pYPSXFiInWUQxNIoI775erZYmGrw4Yecr6kxcZ5pD75G
SZhsBkeLAyiVPec+6XyeH4w2H9OtuCAWDWAcKIOww/LGgZS2Xijq7o29Lsn9Q2RX
rLsUsTXSIsUCu4SDOUlBlwakf55nW/m6xhRMCMADPJ5T0DHHZCLWNaTG7s2KumPU
r2yhKtThKSSVsDOS/mDvaT7amK0NhmBjPV545HSUwLGMTPZu/zLUjeN3UTVclYAp
OzJl/72MZpvu9godLEP8xw98KeOIfS6qSSxbX652G5y0cvdRyjJF+4wQKLvON4b1
Ewx9h+1kpBvf76ljrsWFXqISnRtgzZYE6bqQd1Pk3LOIJ5A5pZCtuK20O9Sq8oE1
ezCHqo3rEL9A8L7l7u8myo/kTCUTmXFGWacRvITnmrj+166uFhAQSuMErmng7iok
Z+kPwFkZBIMAEmLFCp2wwVqJ0j+IRVPFOl2vve6Pv16Lj4KadnouCC0JuLZCN/k9
FhbGJSx8xxQ/WtA3rpXXBHTKTIRfamTPoe2Nd0gdPe1GSaWw1p6BIKOgjFP8f+lK
3VelO5N3HEpfXPm0SkqiSzdQ9+ESIRdnrMSD+ya5o5ODeJQC+O1LEv4UrIU5xa5I
NWlUFBG8Bj7fqcWUQqDDxcacjRJQFh0ep5NA4G0dC+NJhKwYCnwTdPBtMGKjZ14f
Uk22D6FnJZKeqJORq00SZNrphPZhH2Kew56uA/fAd60vQQhHfCz2LZKjCpVlaIcC
Q68hJ+ANUMD7TUicp3OmJ4HtQY4BmxW8Z/y5fKj5CW7+ZesJhyVx5ojqTk6Hi8J0
M9F8tU0QP5NjzBRWBcVQCDtWJIqYbeRwc8+F8B2C5CwUaU06Cpdi9vo+9t71TjHL
0f5U+91sGvgJKIXW2opPJ6i4jFoIEpvejnunV5eUYxdtZjd1bZJvumGAOZsYNUE9
0/jXddTcGJEtUwIb5Mp9pS4btqZITyoZIAir3J1vFcQ/kbGiXCgmXr5ZtsIwFd2v
MkdzQStq3SgJO2BI4xUnh9//8ZV7cp9/ugst5GU5P5ixxZeTRzBxNR1tPucW3Fai
h28nYwVPKqgrQ2vx66TxJZ1zRFeJa59gDFN7NzSp7pV01FI8ARh6wuMVmo+GsaHO
hIpFmugibFZsUb3IwRUyI8E6WTSI9RqjCPa/Ss8TMQGuM9EqmSTUb8xbS9364swj
p5I9frEzc3LIyQ/y2spXvOFb7Sd6b5pN8UEfupYuvqK1wwdSmNB/lJRfkKviOoDd
iSGxkreegPuwiCDiiNfdSbZOwNiWNYNd6DaE33K47qup+0/w6aS1NAZ3SBg7A2cq
UdmfIReyMdIu+Q2P0g6q8I/AOcOPEQJJ3IVKI1HADW6y7YdWbVyZq/KHUEDPSpTu
dbVUoJNSEKrQAUGndrar10webrlMeF+U5jD06XttlwmKU0++vL0X26jSjEXd/ly3
ajU7r40+2KH7f665lEXDCHmn4cS8xZIgaN3a2Qss1Xpn1Dpy1h5PIMWJYahdyi62
J3d4eAhoQumOYEBDWjDKZ6tvB4mm3L03Kc+uVFdd6vVfWi3/wK4N1oWO3TeQjUbs
0z47MCZWRuSMniYrlTDiUER/QsFDZyLH2qGkeVqpUPmFMw+BRYHurC7coFEBy5DM
cU7j7O1hwel4wQRfaZaUI3o2ip7lrGJtVqRID5OylNAqsN8gzefU771pXMoBEIrG
UROzjS/nCpAaqW1mpBqJAp/1vKJGI+7IqqKr5r6j6nEmyHV6iysavi2wIAHOYLHm
LuQ6/qOZUopWAZSKgvZ7KGKdXCjUqCcCHHEQvW06l4+duROHM1iNS0idSOCd3c7w
baHWvWMBRfxLRYLY9J/VZ7NNRTA2NZaBZEpvqaSxAxGEvdJb5qO6fNICjIk4c8HU
LyaCcaNnLV0/U7NyvUYDqqR+t5+a2SM1kTRaUMgnXq4N7/bibP8AzUi0+4S+Yeeu
NFL2avnKL+Xko5buEmjuBvUpE7vh1WS1l+ev0JCjoYgGX/bcaMVnwnhbWoyGnBP7
lkNnbIi4IhntYE3i7NkbRmx7RcNC+mExeRnHREkwWOKypHVlCCkEoE+ronKZEZkg
7eN5f8rHU4ttt1RodCXqpsBKXNmMTU7chms9yFSfsC44n6z1JK7o8ie2I+o4upO0
gaNV93JZM6pQ78d4/9JJUrvOO06wXf0h3NgVyyCesJFAC7SDO4PXuVItv2pCoW6Q
b5qiR7RW5VBTSCrjScmjCIPXWO97CL5d/ZXKlpKRdsKCcfxRh8c1PGCWgKPe7Pp0
wht2rY9zUXSeAzQC3J9Ef3vzLaPDKq4jfZWVbNxv/iXlUiQQiacGsqJFYtDYDI8L
y9L+T8Gr1oDfr9+wypm6op7en0PR9AIPBm705ex39yoU0/+lgt7x49mDWZ+a7bzQ
wulsBvubQ4YIYJX49o7zS7M3Akag5T0WC5HQUUiiL2rF5ZuyLCvCkoL90715arQA
iUUVnUyjx6OvA8ES5qheww==
`protect END_PROTECTED
