`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q0Xg7o6uRIFx19Qu3JpGGLqAsB95mPqJYD4XK0TKfsGk0nvFno62aa+oKVV/hDMr
BH7L9f+nHRv3iIevxT4W0acThp1WLzzshwMfydwGz5yQ/gDU1x5D3fxO9QpK6YhH
+DTcqRlUpRv+wlOqyXZBcZSVDT+wwd9jXGrazcWHZvkcK+6G5reH/WJYRq80weir
1FhKuWsuVId7xXav6v/C8CGvt+pcQ8yEci9tAK7HL7rzmXY8H4se+kZ9JpHRRGCK
CI65q1YQF6lpXfp4/SWKKWV23wH9Ln8Nrp0CSuIfn0YTvz+GI2cOkRsTVK1b3aH2
+E6qgZbJuSvK4ueQuVk2txZXXiOUd4q0aPHzIeEH1TqDZu+mfTqSLY2/dLdGzjvm
i4UlJq7a0gihQhuNfwUURNgMK4Yiw22oUkksTOEe5i5EBPBSfhazpIgo0D7Ldigv
F6VXC55IksnaOrLOWF6Dxd7yJGOHon5U5/OQITshIdv4kB18wOFulr4Sl7oRvp4T
ncQsxhOmmSlTuCcQeM/eYY0Vr8x5pOFlu8+2PyWwmrGvV7buAjCXfgcpAGo/rHIZ
JNdexXCdaXZOUVbu4qMgWzU3sPVhaNENoQRd3YfiPWfVs9rBFAgGVhRZs4lVtLxg
EkNNZZNSkbyRh5ZVjd901mLLOR80gABoujJtrWKXU3CJmS9nirZR05fM7I8Lm9T0
0kdlODKKDCbKvlFJpDplvTF2+uebNb2BwYtNIC9sYwVfC7n9Xt02CygTryyLjqMN
Fqv9Z9xxXIqrAC5TKN74wSjDYhbdW485tb9cnGpNs30cPaFazblDLgPb17ym7jQf
2ZdZ+thcpN2/nIFSFTNRDJEk+iWIr8LRkltoqutm/qETVJHVKXOCFlWfDgiymPeD
xIkOssArTJJ6tx4eN5OKjC1F5YU6qOMQmYeqXDyJaoeOhCN2Kv4TKcF9iaCD/bUB
dSDQPNvddg6fxIUbm0oiDs0OthSkheEXc4m6hLlZnhbt5Moii9sMbrImt8rBortq
A46ll7OG1dpFOrFc+QVpzpbPNaiH95hUS0Yil8yw1rRHny8tkisXN8xOmnVKdYyJ
+sP72p9/C5lhCjO7T1x3PPa0gcbpsdg7nxAgm9MFqLv84GMZOowlaClz60u3KHl0
r+xu1NKX8FazrWu5RGU6+i5/dXzQY/TzJTgxpq6PRtA8F1iXApyYMfeFOscF1BIK
iyT02GnL/Uw3u8YOx2IoTTnCK2QYJB5lP3rC5IyiseZbiUfxEewBeCUCEootIsNw
OkSq9sBYG+ExlPXKryvsfL9y0Iyp783wBMtR5ioh800og0uA2LyhknDGj2zDo4hh
`protect END_PROTECTED
