`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jhoMNkPk0WJo9WAGY63q6uqspUE9zovcAL0Ut0lqqNypPHkb4gG7MZj/OMDdbpUe
cQiZJele5Ib313sTZbkYJTzY05NhpneyuEbJc0EeqWSsWEgknFg09BOU+ihLCrJX
hfNXI5zPscZJmn6CJkDSnbKNyGXxHF1yUwIcGlB1U2joERuBcntl3QPSX6JrGxIV
XqeuaWZGRXuDQLs/OIOkAAtgkbvYPp3R1qKbZjENAmTtLB80B8p7vDY3ETSt4AAr
PYDM4yOeOyZZeoHkhM1njyFLz8HyHcVJ72Gjt/UAWwGsa07ATpQAb82YSF5GD3nw
A8Joub1pcFLV5iAPdAvVfm7bPWpntlKJVhcuSVO1uuwsN2dP3A8vkSeEkU7tskXr
Ygavb4iElisjvLsSM0zdDSPaKSwXQ+99X82Pp5JZRMBt0H4TMRmrNj4ZM9VfnRY/
8csTvjqVFlkP/if1arMmxkwUzeG3AvefSW9MzqH4NR0GsJA4GwTfVEx9hZ/BysIX
YkgbQ+IWvYKBZUHaj1vajocennFiSgYZAZoQQjhY0bRZVbVHaKRudTuSYUVO3Puz
ZytousuNwXgo0Zo3/VCnMqjz7NhnNPkI64koHnhK/DubTKmgm27UV+Ff26dwuPNx
JUuVTq48taSsqjEcDxQPvI7NoNlmVTKdeV1eFT7H42+pJcT/a3MiC+aKOubN93Ux
Kj+UQczEZRYfwC356fP+vdnGdqdjvBwLpzNAXvCflfOVg/yjdGw63nfLlIxis79F
RHz2U6b6lgMOhIML/Y3Zr56tj7oiDyD8iPTfmw9vIqoZTX+3MQ9lGCeH1xKInYV8
xRMkPBYyjSTNc2aHHJFJf1voeBbF0EATLNVs8y4VmS+p2xyFr/SPb9AIy0925GFb
U9MzXkqbjgj6yetUXlic8vak2BADd5lCeQceuEIky65zxjj4xB1+SoTk91CzSdzo
BgopQ+M5EwvaQEGWKZlW3hG9AzxvT8Cv6x8LQ6a+WkD2+rNBl6ZBvEY82pIqhX9s
Et84UFbVx7/SHWHJq/mqryORdA/9yoFh5wa5It/JuJS2ygiHAUyxL8qIDhALrYgs
6VSwjgOmycRmy9y81PbNR0VjgnDaXhF/ws1uZOutQ2u0QLngjA8aFaXN0lPbn+9g
CSQcdRGofrm6BvbkBMU8a8jQ4OOj1KpRyL6w14vG3wGqOkeDGmGVBDyrD0sCgLgT
0yMjcuf1aZhvDs18UIIb5xjS1tEBTGCj1JjhLfDl1LPK1fWv4zQF7W+Nhcb2eEhG
PmN0C8a5mHiag3L/eAyKNmG0VkDUKY12xKACBWplYataGJWGsbFTuPiu8D94X/jj
4sXaUzL2E0r6+MJAka7kTfMAyX4Jw9ES2B0wgHQuOgkxUM3J3XRxbNmEEKZRCrWC
pMqlRwpStaNPHsk2tdVibUqD5+0TdTMf5pV7Z6t3WL/9cyAkekdy8zucBWGArls5
WVWN7Kp++xs5LhIZ/o1sx9QqqqcyUOgSV5GeSTLkM78XQRyn2JFmwViD2Y/r0W6x
O09wLTlYCkP/EtseJXB2EmP7XDUHFxEAPullFgwSQwmuk4dfxac4tVgIKHSeIWVZ
VRBt9dQqDFxzi5TWsOxM4Q0um/MjUQ7w54CrB+BH/J38czmfKi1Pb7omqzSMWyXv
6bsbUxcvybhaX8+VO8jSYyPZTZ95o35AC4L+Dr0XE5Lua30KY8jJz8JT1DAFK8Sm
Ga13lPREL7b2SnSciYMU/B8+ACQr7MfrBzCJSsn1SmbcfVKm1fy9cOGeN371a6JG
gTkP7UV2ZJg+/dcH6+sw+vT24gi8QXtsFY1+4CXhEK69coViiWYg1FV2Qk10i/4b
6US2wSt3GU2eMnsEVwS44HNHynLMEFKhFL1MWE2C6EmqzEWJFqGD6/5r+w6dR0SW
CH46hoOit32izbM29IJz1aPSc6D8aXZX3gBQboV3JUccsNEQQwGStjCJkXUECtga
UycCrAJ9L9yvdYOHjrMwruh1rgpBty1FIVSRoD2Per5ZQ+Ie9u2hDNRHpWz0T+ro
g2r9WJng0pyVQuF33YKtkJ2cCbV84XbkLwDUtXjuXRLjYLHXQqPpbELRX/+IlHNQ
yfDG90U554KZdhXYO1jiePvrSdl8VuObEPxo85nZaDPLPA+uwC+hqz/RmtyiQKdl
7RqYKdRtjQOh7JEzSyTutoqXPKE1F4qEQUwrUARUxfxmxwx70RwIKwBYTWqtJVng
m8z4+WirCGiLaUEEJt0Hy9la+uvTy+Ygk5Fmvz4Nood8vBm67BdsuOpk2Ua0by/x
KxFO53np+yR3SK9CxG6aN4k1c7mo/lDyebm3h2PX2MIq7Af0Wn5eh4kIizkMJk7U
h7ui1La/btLubqyBGePqQNj71dyjpN5UtTN7gsbvIbuEgEED415EgONqJwzXNuMJ
e4dRIX+LbpDMpYy8iArT1nkaVDHNKFExbWvu0nnx6rDQP17RgQG2zA6l2qtcXgqL
96SOwKzV2o5x7pQArnbOL9XjKRbTGMqgOS0BX3YvgvLrlbmDtlCwRQFbxdv1xrwS
JjVmQGgWPeFX6mnNdE5LqidCLBG4WTlQeRrP0dUUnwHdU2m2Nz4aStwGreklytPM
qM0JSMqbRjocTO5UVky9WYolHnEW0v6o/WxpWzGAHRCtIsmIGWnp2v6vgZho0kag
bMhyHuMIpdXQZ9zy6Xfvy6F53G55c1TTkx2QV7zJJeaS7sxH8wlOH/Wqy1wzI85N
ayczl6WlKnwHMXeuU85vIyh9+rT0mzLdRHGaoht7oMw3Ufb1ABnfo93UYY3tvp6a
Ne4VZhsITsq0uVowfCPAEXHIM28Grifh8PQIQf81AdZ3tWmEWAxUNWzsZIWvpwDh
0gwIYH/r/HCAIxvKLIsFJJYG05fQKx6GTAPkiuO1xARrA0LKU6kh+8DtvPJfCrW9
ODPJZmp78DhPmKkpuf5QUQqxEc58BZIvDCcOfbLD4SkduXLfucSb6wmExXlV31go
afnCejp7IHeI6JR7+WuOVjX2AwueGj5ieSGIco5joAFtHO4qvQsJRcf6f4VhYxlF
MLiH2s6/H0QUbZA2M1yXXDNuiKfCvAM33WiUW0XE5ybiXzeWSayOCKXKiS0SYFFi
GxFmCdxz+Cc//7UpFQyCAoKAA0ZNnfu+o5cCGGF45OkAQPzPdyPDRleKBPtODZjH
H4iiHFZ0cJZHysG2CFtaYlfxF8jo9Rbfmt62IkJcZRZ5X9goqVuP/4q0YiW07IlA
mLWG2jHIkEiHmumnyjN7Bk6Vabmc3b1lE9Gid7gEmy0szYUUq4vnHsVeeUQHqAX5
DdXAMgHBY4KoKBWb8jITfT896y5Wzd2prNxHtzo+ptsIa2BpZ1XazqhprTC2IJdW
Unb/fT1x84cKkofrP3aRwzCJpy0aTNkw6YFwxkUEf/nPqnLOY2eO+5XiS0A02p/o
bET/Is5D04U8WrM52+QciNt/iXcaJygRtTG6YOuFOLrztjeQbDv8CCMvr+PDDEfv
8C4CEbcJoNPKIoHGkqOmE+yi22O+KtGpWpsoLKwtsOLd73dPkwxwqPh3rt+n1apu
XsbBL0nVYXoU/5FTzmHZTgFGFuX5jk+WS/Kgsxnfufm1WJXQQbrX3t9xit6tBs+1
VObxp51qdqs8VtJLummYfNlrWvqpdg523X7k7SK6kScu2dHhEsQjVBEmiTntRX/Z
m/MaVvv7vGkSTXtpAIRSpfVZBlCvEHQ+EKtxTmDuvBxE4xvdl7mjsPGkBgmDb98M
bfsRX5TDQn+De4JN7GygMOW41l3J+6LncjlVEgJqs1fEQYKOMnffSVa7VWEvOepI
C1q/ME6I9CmpJDk55BQVqTZf4SgwKme7V4ZJLXjUx+2iyHzNgK39wfe2KPn7h5mD
Xa0IHfv2V5dnSm8uANNHBTAuun71i0ZWDKMHOwqJV/MZqa4au1Sboo/Op13AZDk8
7u/S6w8uEYw6WWYCoO4ndqmxaUzhB07/vVy6a40lqNBrzwvlBuNchA2W6x75o9vM
stTuTAs0vgU5NjJNCKLj0YXYPX1SG/GLm5r0TzMAKXSs75HRCx6343p84wkuv2l6
SMLPw9qAMHAo4K+AAJrvoJYZSZ9kpASFa8rXrXdBhRDc705FRQyEM5Qt3YNFe2Q/
9AFVxMEsmXeUx/4P1cW5ENRErB36XI9IaZ5bk8JuPandVxmkSZoNYVIs8hJavjv3
SSpfdzIu3ByCjGCt7lNDjqcdvbIvq6FxAHChFatkLOG22Yx8Ecth2IxzJ/1HdnDD
hjO55oo42D8U2Sr+38hMahLCzPtKqW67vl/n93omC09HsU1AV3vY4pmU27zIq/so
fgLM63rXPQBihmVhyHUlbmLIGHjDiBaJm4gl82anY9zgsSssFDXt+FQoKWtiZ6Zb
u6NRtM//0C5b1cDL2xzH5OJBt+GI1R4TcFFadnG0MMyMq9hhN8F5BuT5LwMLa5B9
fi8qRnIUbcEzY134HGtBRqC2pMEwDZyM4EcNP+eXQ9yDUet4SSo/A2cI8oVVDSgM
C51LjlD9GAuxeTXXb5z0aF1T7Spgq/T/uVghnDYD2AbgAMAcrzI5w6BvAONtpBY2
UqWhl47jlXHr76VTsyPFm3SdjzyMz/GWjrIUif8YnfsBhXIISEwwwVW82BiwwhBL
ebVyeWUNg3ueb8AcdSszK8GvJx3x7n4sZFNFxDmg3GVrFKjKlv+OU743ih/2aQAt
yktAF6t7Iu9ehqtB2MR/bVWqrBkMf6ylepq2Ikq5GBehDrLLOeoIBT8JvPi3NoOQ
v/EKqabiRjPWWwLzyTkPrwfE1zUdunN2M9PtGkUo2MhZg0AVKM+HESy/NKskRGL+
BpRmFccTsuBY7fbguqEfzX7tpgYlEO2JpgeQfpMHyXJTxSsUNniMeyTunhVA9LHN
EbkrLxbs5/YIC/Ufg3nwOx1AK/1YNN40hi+K4tq8VV2rHmu+xvMZbwteSgYVy6wk
tTbE3nrxUG3rHpHYzP2Cv/vmZMRLMYPfl090S/lSoZrv9JzVGI9Jn47cu50IvuZp
uDI4TqzIYf5r+dAfECyKGQSUOxIPTgf+0/fuqKM1RTr92q8wB1CCoEodrGVq2U4l
wG7dCwkWzrZr3jshePmrZdZ0ZbpK41Zp+RZaushsV2C8obsS6rN8JxYo/8f8nPRr
0vah5zIRF8oyVCBQkIlk2dQBrEygEdxw42MUqHcdlNanJG92r0Urlsb9vu2dxRRs
ITiRuwKTHoBcvHC2AhxFIHES1ucYyNMO8tBoWjtDihwfybDZZgFi1TvyhQG4JGJ6
8qkAHU6nt2ULObDBQYVUXLzeUt9yzchzUs3xVgcUbNFzuQYM2LiIVGO6WVs1ulJV
3UgqrEAX7MzKfR4wHXxTC34DBt/p3seTLmI8af+0U6UbVH6uKSuDc7Ng/vaOYKCE
RjaEfbhX5isCN+CB9rD9Zj+x+99eDhb6FmT2zLbGLSZxN74JQtspK67MT8DKSg18
kK1V6vUGkKF4pPeRYUtQ0/nuLi8wChe0fXfEFAfau4FIgdvgFV08JX0FT41+m6/x
EyPXN9OPBpPdDluqZ2InP9CUKSsbTC2+nOUFnyU+Oy5JuWAlNmAi9bOLDm7DQmfO
`protect END_PROTECTED
