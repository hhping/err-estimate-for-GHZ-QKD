`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Cld+uEI39Zz7fVPF6iMMH6cA7kB8WAY/Rct6Xi7lIcPfIbYW66hZd1JYNhtj941
GhMZ4GJQS49o00mSchrHDJcQqYyTxSGtQdOVS/sxoPx9RJdepAjXmshpXk6FIcNO
Tun8eV+4wIxcj2ezTk2dmnUIm1KjD+/JnFAg81Czb5YAuzeTkF0reO5EeS7Zkjxx
sEngQRVV7Toqh+vWnu9HijeUxRi2Cg2odG2Q/lGN4FEXf8C/KquYONIMB73Gwvsp
A0tnJhVMgVc5laKYFT2W8ODomHzGD16siHeiA+yt1njehWYOEL8ZUFAAhbMgENAJ
HUmAZOQl8BWpTw7aZq9Wvl6aRB2tcx0Klyf75sF+0E7/5f9XTrqeGWbq7o5KcdR2
EgmGovHgbe+EVuz0+78icwOXFHkxh6b0I3/l/p+jYGe8lZvJVf5Sp1+HpxsFsvkW
m1DPTckNxUym7McUTFOG8Kmidwkqob8Ib3Dd52Ij3nQC7n41XLjEEam4pIe8SrOK
21bWcDuuTspXQ+X02JZ4z/jpEHAAYgzIF+jkxpJsk/ZjmedfN0dVTPCuXQwFXL2x
ddzqqObk8J/ay5qM9FcOtBRasj2CiG/xvYWKxs2gzO0mWnJZXbM3rUqaSuJbmgPP
lWcyd+WyMQq3YWEideh1/Nd4o2vtnDu1I8LnyYjrYdV2g9RyPM99tmPJlktIVa5o
Ce6eAGu6FpJfWD4KEBTlxnllWFFCNVuQ3Zuk5kRJooetZ5BnNG63M8JLk3mkcmDk
pHpZfgqwFPvHqCfiYN5KLmsSZApvGUQwhdAko5+RJAg8a5yMlbR5g3dAYqnHBPwA
Dt/wJ8qQoj2wYwPnn81V2Kq3qMQCDmK5hMKlJAEhLMFF5tFUYwoqsMSrL2b75tdT
+VZvej9c48cjWzjRM5bfAOABssuld/o5X4tgFeGoOfNOHTRractY/gofGAmtluM/
E9UdqCOEaa5K0kGLFH3R6UnO60zzYAht2RhvaZFKQNwuMZs+KOBhdzaVw/ev1XuV
fViyugMazXcyG08Er2yQg2KNz758AlXgpXgeVFfuvVHIjmnk5RPM0tRnN/EkH2zn
/weIm1Ci8ku1q5KFIpFKj/tQdPwdkE29I9vGAfvVI2bkrAV+aiw3iIIvEDa9+JTl
NVkX/vxW1dkJZCjzCvff2i7b1cN5j8Sg1kIfX3dzunY1agQH0SNUiECdoTtMG9Ul
8Fer6ZMlVnK1ViTYl3GdJb71rYNmr0d7ysMA4rLwngha3gCWlW9PQZW+JiUtEmCO
T7+hs7YFBO3FwtS/RT91koP4/kTzFdUbpp0GTx3lIBeY+1RrhRX3q+2PX8w0h+RD
1D+AN+4f36VS6GbzzA86qGWcY1G5h308DfXQnsNE/ZcMl2EGuJzGX0JQbKrqGWEQ
D2ZsyMjepZcXyYUs7igtNTLHUAaR6mENW9uvB06kXZC62tQ2k/VHcxMNz9PgYhYd
fvFqed+OjcSmITI3vPWPCp9HwOi6gmxYrJH+0kKVJ2Sp1KX799+axydU6n8pDY3C
urkqBo1qY61qRCOSBeZZRPMvqaMSEzkTN+BIRFUk02wFGyg1SiyUz5HGowcPCTrd
78Rsnf4FsNvcbpVeZtkOW0H8ASwVFELMANn/FHY7SGKH+NlTQyGcoaIpDu/xHlGL
h4W87GxcQ7nUH5ELRrFv+AcKnvGMqlhU22gleEAWZWDQRCLeCXTH0PaH5iH56t9z
7tZr6XsaKrwiA4GZNz4ulfdroBMs3j6mSTWKh5vn5ZIWAIR9vgzYCWF/ul37/QRi
D9Ib0GaT/M+IEaqvxqHqksxE9RPnezkP85DmwdwpJTAMvMoMQTeaI1BrYVfk+Kxs
aR0CvonFnANbDBKFi1ImHOJxsOIBuasQR87EFVGRGI8thChT3X1/DpIbxfz05SY1
XHeWtqETYaiOSgUAA/xMBVHww0mD6kZS6qR5nXGj3PaAXnIsmHWDJ8c8mlg1k63o
PteeQIw78ImgsPU5nlVShWPWGcl48ac3Ir/qiUbn3S/9g+2zlri9UYb1msvmMC9v
qgCEzlMGdzelKud3wAsOkd/W3xn/LNcZu11rpJY6RTpTWFV//eA5NO6vcBUTz5LU
SlYJAMxGlK8nUDhVwtKTpNaKXCjMOh3Yz5RGUl06Rx3DXlU3wyt80KCGJB8aaiDY
h1QP1dOTtwzznrdGYEiQCJxmcbXFL8gRHpPiW1UvuXQlF/Tj0aVCIx7AO2yMvee2
3+0j1LOJD/fjyxpHkunfgqDHPLUHnjG/+ddFW++h4TBfBX3uIas466lU2fc/yA1z
WPgaT+IKUS7PzWZaviIXyEwdt5oaDIfwTvoB0dBz9rIKQwAFwO//p+BFTBW7IsPm
LlIcCvUewUZivi1ETPUNySOZSJAB12r7Y65JnIZ69yrtbQHaKCzsMWRhq+B5ElP1
Q8QUBr9TCBtd9xcMDT+m3MXzhjRArZS9QQ9s3kZ9bVqYQvx3OzTFyG5/fuuLk3zs
O4BDKUHyc4C9BQnq9f8DGUQFRKrWTP41+JeHmlOiomuP6yMLKG74L3nNm0PcdZFF
BPqB0BfvqUupfIDh+LHCr5GQ5c9kRuEb33ojMuqrOQHPu94l2FB6OTYJaeMhxZ84
A3BmgtiP2QG77SoZMQgd6AB4Oxd6BgZWvYoGyLi2mRw2my3y05Aa3OEMvuWV6xTL
f0PsamtaWuQoct0xwQTk9t3FNZLZeffq3CgHEZN4b8LOEveiIoaM3ysrfwpYZb9x
WtTkW7Zb4Vsaacr28goNAo/FncQdXXtTqHwCjZiDG8Kq+g4fAzhNSgh/xqfe5Ft8
DCdPpAkbuV7x+7wYhX8wvXDRKsVmOei+r+a7hHf0azoDJWDOXPb+IjWJx5LvZqcA
gqr3Gy/VKlxNPlFmqb5vlv13KTxQO5U80aogTjGZ+s4GNfzJzqHMr6aWIsuO96Zx
tpk+7CaVi5lfPZ5s9Gvuz9ZX8HUR8b8X3PTk5ZYYnLivvElvY5AOSrFt9CsxDb8b
7oXBRWWUygZ4y2ztqlfTgP0DWQnnczYAlAx3/d45G9znI/i4mctC+gENSeSHgHXe
eXM+K9ZJn3TWtvvGsdJ1f/FH++DAzYNT93yFCqXOzVm4MynFHVO6rzX3U0ASwG84
8JxDiyK8ikpb/uftbhndcd5mqZAJgHD58+u0mVyM2tMaIlmKBg+jabSmZkzR4YB9
XqIqFflbHRO9cXfN+D5rCcPHarj6twnxlGruMUHPKHkXrBx8COrJWFnh9YS/9P4t
vPQ/4e7Q/YE7UiArvkW4bjMHd4KKtnSinWIDWVESBnZfKoFhbVrH4Sc5LeAXc/2q
Br24MCGIbn7ujhKwkqcPtvXnQn9G9r2GbToIJXXI5/FedL36Zrm8nq0qdv28FZul
9B5J6xHxXqQmyGi/w5LVcZGhNcBClpSBxo57ECR2A2xOTknrd4MW2otpNLdxIP0u
ABjhiJPYNLAXNs6UWujF/AG09dNtCA2pIeB7kqnLCTwcFFO3XSAqMXCmYJsRfy25
Pdsyyz15cYsr+5w0R67yyaC6zcYAvbP053maZqc7V8Mt44BhRO4xB3Nh4sBuOcf+
HOQZkOhmPD4CoH8dHIv3ZCJ70vrc5bIH51Zwxz1L44FHSkftWfcMul8ohQsYzkpd
adx1MroyODrNUs4lbMnG6vNs75+q8yPVvhZWHzAPBCSKlCYj2UI0kbT8Sb3Tek6Y
0kiFNqC5za0RO0VgiN9ILSkpqwXza+WHPCMQ8zbpq3fRN+28XVBZFRcWnlghLQaw
cspEyGZMh2I/VRiXsw5d3kTtnP7bSpuRcaokB4/SCEQnYYIQncvqoBa3L+B+3Osf
O2sJrc/mhhTo8DXd1O35Ky2jfVdfkuyt9MB/BEJ/m1kp2+rvoVku6JmYSjNysSZ5
+0blV3CRlPrj2VDZEaJnjUKrTv18A1eQ61F6TeaEuMziZpfoEi+8vQzPcob+pIQM
Pyj1zXCbYnEaML63k+EklVlaxX8md9OF8c5PbIz03ol1xpkolnieVfXNUT/DRZ8/
AFQL9uxjdeWQA+OldUbByB8ky68egcBozAafYOwrh1w/gohHzODbYVlV1ZeEKYm+
DdoFGG8y9fXvG7SB0gtEr3Cbk5G67cD/1aFM3zj9upfxji/qg/73YFcH6n2EwmcL
vNC3nQ1HrfDHh/VHYxPZ1GRUhJCvNieZLreKIwVsCgW1Xa1tRCnn23lHaZ9CPqfA
Ye1qShIAKYZzuTz1S5LnulZXNwgbL4ZlbakhKwGE3mxB4dw3I3y3XLdZtk/Oaxvm
Jb7mUJzii+W6XPR83abZeECVPmy7cYc6JlSik9jp+5PDZCJPSVB67T2R/n02+RJS
4zb4nUuPkYDUo80DlIKrQ48sfr07/LiFNWAnQsK2Eix/f+NXxAFb70n5k8tZp9Qf
WzdxJuHhyAccLRhUD8r2dFcGkeyi6AZawIyQMltWCTtjIz0SMs8YanY5sEgqFaMY
5Q2Kjysf9tHERB9s1ZmUfBt9uYAWQrTflLkzu5pn7BOE6M99LsbPaJJBcsJhu5x5
GEV21WALnC81r1ua2d836aos9kjzo8ByiT6L+pPsxJ6M8aeP3k+wGBNPpoDjWhFZ
Gmpcs+W5PORpb6IeTKPEG0X1k0olzLlk27CaAI47+Wxs7PCKPFY29cYVl3IX1QbL
55ZEdmHyzAu7oEkTHAy/fELsuFGnltCe5Mj0PoBIy8azjfsMGQ9jeHlTLbUChadM
bmjWtyYWYvtdo2Liw1ebcBPAZPPC2Mt+vDztCkBI1erHo+yR/AN5QLQutPAxLVD0
hczGFxRbILbBd2riMRfymQlEhd91pyFa+l9FTbqy71BlDVB45D5voe9wvlb7WwFN
gq0BSRwBtWjCsudHvMcw6p7YT+SCNxYpqEkUAkYQIaX08wCWt3Gu0ZnXqc85F3Ey
dqzZP35gRd5XBFABteupDrwb7ATbMBCaZZacCA4DWwn0C3BxGBm9ZOLg+dVl0KFA
Gyag9besH89kZBQD56xT56FS56pjpHAY1UG6lfWXgARvaLJiumH3i6B/bSLeH/PY
TRUbJVQ9EOQuoH0hJqMxU1mktJST5KOTwG+Ad0trEs8lDs+p87buIU/I++AYg6pl
1GTo7JbIiVyPa7NDjlHnpToCsxxjnxoGqZI27u+9d4OuG+3m5/KCpTRyd/x829eA
zwUlgT/jTGd2HkGDUvpJE8ra99SdAXJyVCz736qGWicTZ4TA0boKuKwMpXUotWOO
FGUUk5YXOyvZ4aR6vWUcQJIHCB3JCK/SkfbnQIdJWwWYxaEIW+SRgnkD3eEhc1zA
1IBoR5H+cY6AusqAvudB7VOPfr9njWTLzVhkooVpLKCDswTwVHBo9gwuQeCo1NPd
jO7yvV85wLoGpSr461USNFFO4gTll6TQw2399/pFxjiKy59ikg9NXVz6Vy8djsJ6
DaAaHIKof/nKCUe7uuQoxRQlmHinnXgHhAdScbbEB53ghzw8gHnfPPo/gZYoDFpB
mztsbyaYtwMeePSaNY2Y+jKD1mKauHqcUfEKsAV/hGYo0VscbjEvoaA+30WsnuFO
+TEabJpdyk2d9lVUzZFO+QzJFTCxUZSixY4qnyYQWa8uqNk2Tk6EwuV90haVcQxl
EhxtiaBXUIQ8waTMfrQV8cVck07glOevWsxiAL+ZQmD7V+tZFsUV9h8cYBD1uUXU
3f06d/fdvOBBmaCZFybMFZZmMo45s+oZ9CDxQwk9Iwu9d2pLvyYVCUIgUHUeMmui
evTubYZR87D+nF23/qWUwZYgl4U1EckDdpJja73MrAzRkqrVAdF+JZB+SuxwBqH3
2/bJc7VP0Fe8PTxxx9qisV67Tyjs89IxVX7/mF/WtbeE0rpi4XTJ55sBsqBtQ6YK
eXMCnuvscTQvkc7GMEc1hJiSB5ZCBK82FYSk2p2dCoDRj1LBcGoVpiE53dbyUnZV
RlhCJfzbH+WvLu9yFVCmA8vZG9+EwIS2kE41CMON7TTnPYRmigmFgnX01r7jZi6Z
7rIEvSGTL4yzrsm5zvpbG/6ORM8SegY5R5rY9AGy9nJqeOb95SFvEz7si26tez7m
YG8eCDemB/YEZBrPvk7Eizle86FrnJ5Uaj6O1Wxb6jHNOFQ/9fGGxyLSXcKBA6Mx
Ja1q8NDUsOb1wwtLKj6LzlL5Gr3RpCQl6cGz/XvntgG3bgoR9JqcrQ2N+EMcM9mR
a6RUCjf6mQRKEzzBhW4NpAepM5ts51Jq1Vh2hXPiY4gPGzp7uQM1MZdF1QsfSMM7
IBHuXqcWfUsHiNiGLENXjulpXUl9BV4mkayQbuDpOHo6Wm+rc8lGQajU0Ax7jQWf
vR+mag/tGqoOunCBQubiiX4xsVMs23ZjEVUQgHu5rgnj3/RTRAOIYqe7SUPYzhw9
ldP/5yX2JGcQu/QlR7h+c22T2vvJ+a2Ya9A6q0SfPe88cm7igLIMH1BHpsqxglw1
lIsSr5zsg5wg3m6D87PZr3EX7S/KZrqfaFZUzk54xbEIBF/eqWvX/sEIMBwPdzUo
ycJEDPfjsgG8IZP9jJSCc4FhsQo+eyMEBG5l7sUQm1mHtiTDCXAoqEGgSWmda0MC
2qXw2LUWUKLj7BcZ2rEMLbc9jgQf9lK12Bh825PyNqLedtRP6Cs76bfDpHqwgEf8
6BeRUdn9MiZG3QlRMOgCNIs8+IRB3jIMcyd47LZyHcnfFLL9iavUuMx9Q5upx3mR
7ge+o5EpFvpp8lcFQXtY3t/JV9kjgNqjo1xts2Vup7BDzg3HN+b6s2xP4Tq57/34
xIT+fqhkmdN6z4NJO9qn5qFZjuSqOZK4KCDoN/IU9T8zqVubWPV3MTPC2T2DE6EU
Eh9yBPEzntCUbLUr1TVcIDjZSy62Oi2ZkPvrQJh+2q3aly1/7jgUzQ/QHK6cm8np
2GoCH0U4Poi6u7jfkxoieUfr7yd9etSfIq7+BWp0L0Kd/Zwj/azgBDNIu3Wdwy0S
NsbvEhMS1o0kH3uU1jpaRhyOYsXl8GqEPOOtthBcK8h+pKBvqlpVbD+yJ/bCeNtE
FCx0hNJwafnHdtvV+QY6FE/y2BM3YJ8hvn8d3MwMdI5wpD1xqImDcpQUHB6aHyvT
F2bJiGm+CZuv5oQ0KCxJTDjY72i616K+GQ2AiOpHAzRKpfXDz7SqrqNGwzB16fwH
e4UjmORwVtZuBidHZybUVXEhF2n7tldIFPs5EsfrYkf5d+EsTPWD6GL8xyeOFUPG
Sheh9n8zXdhNIboM/APwRCTYa/XFXkpgddn5njNaHaJ2d4H/bCMzwa57qhzfr4Ev
JVmtYeDoxhB/d273K4Clgc1xgwaz9Fi7yfh53s1uaWEwN/oxgCLLtVg4NDDtU8GX
KaefIZLWJpft7XvtBOhidrJhInZbWBhSQAxUnPAejJBuPwxxoG91Iw32HZpMBoBT
wjAXqE9IBA+8GF9PNJy5B9IpjSoznSy1RpkhAFvkYIbrpjU4ti5cCJb4beKdmsBO
fzRn4sqg8FOQzkzXCmdKyM/yNCfOk7/p4rKl4bVum/2Fu40u9dxgKFDsMVvsBrME
LgkoWWabkZSFtNeaswE9ptPfOj6J8IcWZ6ek5TjamMOzD/kVyGKhKFDEEmVfz2k6
1mnLYhueL9F16uq7EUi+/loD5ixslnhptmmK9H63oqW+cLS0mNlC9Zv1uvKIfXhe
qwKtf7Ha6Y0e/yWuNZzH0FvEmN2tQWxgclxMeUrOJs6yfaT2VxZg8MO2Mwsr9h3V
tweMDcUDu7OcOmVQOpmwL3FcTbjCCmZUdiXX2bq08k9VLLotiECF4Lxhtqab5NQ0
C2jd3LnjXppiq6viytwxA1qsKR7+IGOv4ieaMtHNCWPdAkfbXUB2lh+qHcXij8Iq
Xuiy3RxMSa6AeBi9GzjIHFhMEee3UNMIZCdCfzA9+XRiFkG2faswRMESmW7B6Fjn
ixAKT9/yNIYfp92Kv/ccUIPndY6WP4DN+cGuzE0qyepZEYY3NUcAPv3KIvQwXHmQ
nUeR6d7L7olrqWV3vScFaE9JB0HwZJ0iajE+83pi5wEFxbTySibhFFK1Nx/qwtZU
Lsrm/ChCI4hQPdolP6qzqXo7Zvcc/dUGw9g5cuJo4M7OMgPpdzFrIa6SG2yOXBs4
weW8+mtz+996Pzu+a/lKwvYc7P1URNu1Bu70fX+0jiUPTLtCXlSKbDIUnSqvC6JE
/2lxWab+Ugz3yegzvjgQ8cfdoARIfDeCcly2GWC0/3hTl10Gp/7e9emRXUi/dcks
Zar0sZHUZgW6+PJ++/zoyfzkr8Jn9mbmUOcsROR/Mz4em3lJeaapgpDgr3IhP3xS
4uD9XsNvYVx9TPYSRHzsvJ/flERPM7ogMTWGUMFOd4cIPs3c//WOAVmaKs2qfGuO
pRqsXMDAk5BNHsvIZ+IF+EzlzsJ13Ecfia+3MLMEe8tujAYxpg4qwsyVIZgofALQ
AKhRBVR4nTBzO52fmwnsBGvxIXZYSbJIug1Rop4Em+Az5f19EYQPgp0zzBpiZsi1
uBGCH4o/3SUnz49i20nM6cyRfp7tf70o/oSHhaO4LjedzeONsrzh8XewCUrP2Og+
YtHG0BvL9u7ym9Aa0rrLibjUI4nkZ2vXsB0E7afYPuwCg+90TxeBQI8Bf1ra9sN+
Jq2sw23p2vNYm3QZpFc9WtrhAZUHlnd1DRPCW3ytLJUAB3s9+2sazgCJ7IgGrAjQ
filjhzKVYC1PR3p1OORxujwH4l52Or/rwPYnh8Vq9bXh2jziw/5Lp6Wn4qmOE24a
oqaJ6kTxQcXMvbbZF+qmL6CP5/Vpb0u8YOpNN7XMhN0=
`protect END_PROTECTED
