`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tDCCXpUjZX4EGHkQqTc+WRV0s38iyN5tiDR+FUNk0/4GQVl1EsEXAOMeaORlre6K
3bY59ZOM3ulRccaYZ6bWF2HrPyeRvJAeTuu0wEI9GdYK2hdpqklWu+zHJ056Wujc
NqiyAlkotgU70mT7FFJ12CNEoClxHOGElQV6S6kibKV6MI0DoVmyG8Rq0sxfvwzz
IefmUmFttAlpHpWA4T5MF7bhs+7QFE7elSelL/0jXf2IYTZzkPNJkaRk6vkmr7ZP
x+Q/oKjP84/XQCF37D6LMEtW1Ob3zvTKKyOQGgGBh95i9ESqG8sElcki054u8i69
qiCq5hsntDUhDoynq8Sk0hKar0cQEmQBLdGpTAlLL/NZBSdjR2eDbBR41CQOouiZ
wq3wc0gIyDGMlZk1nog2or1gb8mlBS/YGAJGOOQXEeA3UcqnvBZ1Qd5bFK58qkPp
E8umaNHqqYRHfUBdkund2FhEKgQvVlXl44fX90+iSmHt+Ma8j5uVtQo4/CBKJRRp
AkDta4wMYxUVO6Nj+ojizFyym5OT7u1JZk+i9Xqa5y5WhPfD4J7JvY4kyp2y5ADW
pLFIDG4dim0h6wiQc70+M/mwJuOiGXblpevI40hDV5OmHVdQKTNYqfF9ER0HBVp2
b84bbYsGPVC7mfLUBmVsFB4pYtvlhz+4/TJfTX8V7jvfbWyDSRzDcSDn787rrxFK
ViknucxZSw7bog7jSGEQyM2jMCnoJajA2dKS6asw/dDUUkwD+S8igZnNChuyJ3r/
u+k19NQmgJs8WoWR09SG+sOxnsdM+U4bG9/GVVo8Qu2ZU+XkG0cfLb+LydpYZ1mg
KG8h9I+RC8SJznWofMVay2bqYjaqbh7+RmzWiTVxC5Y2/L8xjZNGznAK2fhEKVF6
afB3Nb/gx/XUlYle9n3YWJYdVrspmxOgNMzDpPJxAbCGuhF/8b0CZKfMGpPaQN3A
yq2YAzZ7iCaGtj4Jfnp8XoWltsHX9iZU7gpw1rkl3fPlSXTQ1lg7POHpg0f0jkwq
gL1y4rzJzM1Pbq+Ev8a34rw5csd9qq/B1w+UpGG5DBRLyXRrdBGwSLWBisQU+D2I
HIjOey/pmqfY7tJSZw64mBvcHTlODtQDY8CSmdenLMAuKgmAd3Zi01r3BdDrutWB
dOIprXekYObuuUmKnQ+KHTFaNtcmu+uPMT/HFUVeF833KkKoyp+4Qb1vrQQUhxk2
95T3TbvomOSJ4b0J0U8PJoo6Z1Zor1dLLcMko5G+sp6TcySl7Yet/zQoRla5CdvE
7NBNiJ9rmM9T/Ub0IQB4vWdUWGQl4iOvTzQTqvqFf8zIjInSYPXAdd1HsHi+MGNt
Zl3ogbt98nqYh4QeN+of+1SY7Utsq4TlYnynBySxgYPBwvn4t8oQqjn7rkT9LnuF
4YsgV0KrqdAiziP2vVG/PKOJ6nkIDzHmVhQSVfWJctJk/6DNVzHnFjgN95g6QsEY
yEa8jM8IiA/PQrKu5bsecaITGqwQB+xZgvf3TwyzjeKAipoj2xex4ExtJw/d9fE4
R2mda0ykFjZ8bOr0aqGc3VB5JX7iOa8zL3t/b1AgL92X2H1rqm8OX5NQxUO1A8eb
1ydFadZYfEyh/RThtOjkjJ5iYlogkZNCgYH1+EOCOSU1uiqBPojomVFrKV3m0iJ/
ybYf5s+kam2CQiDoYCZpPdw62wrgBCiWofgnQNB1+otlj3lZ80N1R2lUnkE5pgrc
FC5qpmAUjqDj8f/3to5BBW1iCo0fZDKsoEEQw/UvVVDxmmUMkGbu4iskSqa1e5UL
w7nodq978M0PRJGWqoSwLTy9P6coVVbgjEq2vOUyVQiedXwJ/25sr6sAhLIHQq2v
b7XGPtkcsmXTcO0tPGT59yZvC0bdNBYUiiQLzicmbdZCf6kiz9RtM5uUE2R3eyR3
Tk9t1tO/IJBA9VO+JL2a1x0Bcj6qSgSuAV0BqTnHClvTYT3APu69ObX0Sjtj6X6S
0n9lrkWJFEo16LVZpO88xrX0OT5nBMJ6OW2XakxAL4xlLuTZj+3GBHeiCPi9Rudp
NdYzjX+zdpw5greo5X6AEWCmhrYB3isjxzkht0n63cjhuo3OXpCT78Hla6rHnXtU
/u3ML2n0rhqzXj620sDB0U0tqsCmrI0/eNbpFu9xzkOPPhTNvAMDCdPGVC5ffjUE
UCLaWUEQhrch2zCy2YQTHXyLjVMQC3ObqT7/n5cGgBHAIeu6VzqxwQXAaGP0CStO
At3urOJrf339S7RNlkDdrN+Er6Wc/yzIGCH0lOmlu8OvmHtZsmmHz1c/g0lGbKHd
JIGl+AnWGUQrZfzd/+shOSrgd9ZjhbHcPJ7XNZWOstRYPagvRgUDv3OukNdMEV5J
FNqkI7N8pAE0m9FAKZFr3i/O4n9AqdE2v9T6LFyEjwrOW/EoiIJl5jmCcTqkCIYa
IjqrFPVNe9NFV7CwOLTKzi2ydDMu3w/5BjhEc3uMNQGpwTaUvosO2fEZwiiKVn1Z
5yaiCFHIaNTshwySxy0Lckd6n9DqA5VQ2ZGPU4U0OU2VzuysNSDn20RMeXifqWUL
YorXlhRmkH6Y+XM3RzUwzqFog9VJT+tKvXnGgJHz+zBOU5gP+GL2FZFCrKwWuOEq
y48ayjNoxpfg4rC2DI3bXGD+gl6ZpAb3o8Yd/S6OOLfBPH2zvHIprtRjf0KLqSgr
0BORUgkZ2gYXGsU1/P3X405r4ZARWQhYR3r2dsdNuf8AxZ5yPzAkYeSnRO/F50dz
PNACld/K+aVV8craDne8Sf3RdE7lY3WE5cqay9Qc6/z4OKVuB9O/r9vg38/Y17m8
Ynbi9MHrUHXrymTcWDyJvO7qp3/w3s+Zaq09B8MfYXT0DClDkNDD7m3+agee8NVn
aKtwpsI61bBTwefeN/xULsJMIAITjhuFwtZtUpJDl0sqihuXnbvqlVbuWcTxdzD4
CoA1lOqHG5xPsix27Qb3Hx/Z/62H7f2XX1Bcq7siDRkJ3DaO/eVEbWCX//p4hwwv
o8CCEhw6IREUx5y2F/aMzRmDnCuaY3VFtk+yU5sr4aoOJ8Ds4ARwHaGmkz4KyYl8
A0xEatZZrH2pgu1OldQVUD7oPEMLR+8IMinpHZYtXHILs8+PHfJ4s7rtJU+KD7Hu
oLXdvVpRwCfDUnPowz0Ljo4ukjnl72qk/aq4RNQxjUVdYJp4VCYKxjZTV0TAJpcc
QeJvl5FtoMzMLmHBWIYkmUKCemNrycWMF8txNqcZGYC3fuOzLMb6HNioN0fV6Feh
0528WFXzPhVKX1kLhUcgvmKfOq9b6mnlL+obLW32eY9ovKF4orXRTuvNFOauqkDe
LimebNEmjq+a818eJ1Ssq9qukKnZKQiLkuaoYuYu0njYDIBbl3xN+MLnmyxkMOzK
kVwvql7fHTLwwFTAeUhqG2ZrIL60NSVADQpIQ4bV3w9gKuuDw4ZnUFoGN24u0FVd
+ur+SOOtep5XGz09Xq5Zl9OlGKum+qdQuHwUUu3bkkaqV4SgdKetqZFLag7iMYsv
cRtl/jAvHUtNrBiEBfnYGAsWXgH/HzUR3gWiA9x+UgM5c8OAKX8z0FvnbMaLyyrT
Y44lzC8u2O7kae2MgUETwI+sE766QoTMfOo0a9pzGEll8uUosBt4AQi3N2TTjwea
mB1svk1DQO1y/IP4IjRqqfBj2JIlg4uuuRUZQ18/RRSroi6n0UT+3EHaXyeaoy4j
Kw3ThFT5TfTBLGwLVa6CQRQPsr6Zq2TJZReXN4FBQCafoSlm5B3m/7bHK+jos3H4
gCcwaRyje/oqjYJtU9lurOdSD0hs3fH23pt0H6paaKCOUQ5AH0eVPOee2H+m4hrv
h0Ee2SAYCNmVNenNWIMGbxSKdaWDBYJTQqBQdTXeqFdarIDJjo66iyAaQ0jtDHy6
HYV8dqbBO2ZTyRqrDUTNswBvJbD0pI1M3i/6wmmLc1jFmB1yxa884HQUarQARFKI
F3uNJuvPH4iPXX9MY2ic31Y7ss7cE8pfcdU7cSMO+eAH/3be0gSeexWbGafjgF6c
8kPmaSEb5O0BPtDCGzwwwbKjxD/LtuEYZrZ6qRRVPmmb5v1tUcFKPGPzEYgYNeCg
Jr6SnIrqYg345ZSMPtZe6K7NM5Sb19jlf+yt7p/WiUJaKPBbjlxi2DOgajb28bFp
X/cXQENiZyUjX86Pc49Rcr+gKp3477Ouy24jPlcWTgFgVTKm7tfaNinZY3qE29d0
/MuT/O+3w3MJhn9Jd2bjIuzDqWcm9MSfmvHulA54ILMv5qYqGuU6Pu8JBbBOBOgM
18aTSiJm8vH3qTdstvnHRBoaBMOBuHI9z5EXlRoEMQdHSPM1zDgQZHv3rfLfFeiq
yJaUi5oEotwI6GHWc9mddQwMOzMqGoD5jr4Rf34rAu5NUr9ThcJjKJtjz2Mar1do
Ya4Y1sw/rBt4p5YBbGGILNRxbfwJc9yfJOFGWz08mHO+q3vMfdklOJbHE9uyaIEH
Ln8mnr2N+rqcA1HvsiyUcU7+h1kuwifFn2fWO13VSPZGl8tpfhhTUt0Ku52iaCdh
8jMiKMrTT3t9j+feX6RA7aD36reBpwUxIW1cq4IXlCIjwXvklCoG0Kkx6AtqY8Qm
kZ9Btc+wGzb6lr3MLLRUJrJykVIkoZjIfDeDHYuZ/fIrcz3gwZ4rpjGVyBvOjJqy
JLYpirjJT/ugN8LV1sc/zobo1KcZyejhbZ/unfgqnoYctme6NF3Ei84AhlJYLg8i
TzoU9timhovs/MrTpWUpvt3aijSnqaxfKobeclp9Y7HSvJ/iwO+Qjo2TgFwtv8vr
mB6BFr4XWit/DhSAVyQF3IxLxiZ/qB1p3v4UyNg40WQA4hmgf62FiiOBCXZjwovh
KkCIVGibyWuspRVhdhViaAC9iZ2lTCAd8SMKiw7Ggtol755lEaMrxAex9DBcN66B
USSg/6fJ21AME7C+otPlR41YzVUKJuBI8DfP8LBgWee3mviAJKqruV7XqGXrEi07
ikTgKrqvKQIBmuLD5Xob3jAQfHEid6QcAtnzvpG3ZzBg5H7X4lvdhX/TOz97fv23
WI/Irecm7YAJBsixFRutpy5G9+W39+Xx9gRIYfQmjxKOB2K4UQ0j3Y+/Kz4oMGep
gmF20o6uoXixUwU6+eGrns8ntOfJKlEOzZZPfpeAOVnuZnK4W31ILpo0ezrFBHdN
Cg8jK+/ZRiyyBTT3XETrQeOzbn/7VkFiFUtIWL/p8ERNxOFEudweYatxOp7a1X4e
Cj3KuwVl0YqQfHAdYixaOFn5o9x3Yh/E3JLsU4WdqYdszdLHzPg199zKNUa2vJHx
hZF04ncl/aELuSAbC9Zi9PxMLuCV7D2f51v+LGir9ueChRp7aU0fCzGFDyPnH2Aw
V9XaLltYw7F2/eG4OxA3hhVp9Mel/C3HsM9AQsXOM/D+66xNKgGJFVHkmqMZhhAO
KmFDg2/Qcvm0Ayg/AL+DoxSK+ZL59YMNLzVlECUUZcoBK2Wsl1dkfS2sFKL+t6Jr
pJ5vHsRDFwsvwUFsDYxkmytG7eTixFloKgWQ2SaxXpH9ULLXAaBxE7eWwYTxX/1d
0QknOnPgwyjA4dnjfBw+AyJqFvpXdUJCyCv5BI1Y51hE6gdaui8R90A4Ccd5fv13
ViwHoY3MDXwq0HaJmUBFix+U+JEfnFCYTpbC+mKrO7r8OeMV+D4jfCOHjlq4XVOO
5TkvSBCVaUjtsNkbbnm1uEJ/0pDpZOt7lbF3K2a+I4Wzp0meGg4yBHpKodrSXOoZ
e1VOuc/vrNSN7cLVVcpzYLmuFUUAZ5UwhhXAExt5QlDA2hDlhUvRLjRw4a7amVlk
A6r6F7JHTT5AjT94UvjvwPlnzhtsKjNeiHwrFXmHS5sVqPm8q8uJ4ezgnvmjmqPa
dcv9+YEPWgbTB4D9W0mLpp5SalbYoHhycas35PpRO3CTWW9SXnqlbXcBqI7yscbR
gzYPipuQd7FvqC1LZfEKS0xPghQiGi0ijE3qEgsLHDV7JjOSgf9221mxhyswgRmi
iXwhITb3kgt2gutHFWK7W0H7kRZw2XvbGebWWIdoC8wdGqSvyMrTCRVcIr8lFHzD
A8e70TyZ0+BmD4pP2VsqKH9gnhpoJ8VtBoQ9iyKFQPGlSors4hgpTNhqBM+yPXoG
AtesM8rFY51QYbrLuxzOkpnPFrohr3O0gvHowVvceHoZi6+/7VytJlvmXa449NUd
LNqgS/NLxD3mp9O5WiQcSXiqomLGi4pNoX9SHTTN0baUZbnDfREBWYi8E5ZHUYM1
DMn555BbyJYvC1zbaBGklTFSolfr2YswJiB2qY6rhupgIQ/KFarp935IenYGTCZk
30PELkb5JFnbr27NMzPqo05hy1N7s8DOTNRu30bMCjiFCH6wouLyJWKnuSosBxsn
lJRW9qrM39lMz6qWsr+YCj1L9ntrLY2vWClx2v1K7qMDgUQ1JYngEcWCMSgBJbBM
kYKBqD4cMwDDFyuxxUVv8yBZRI2ZZhnHZ/j5bPZkEXPbnS4epfXHKwNH2uop6+NM
/3Ic8ZiTO5xEClFcYbubbe8FY8xGZUcUuKDcAB6IZhF4TOs0huBnU+bBRQPIS1YW
5TXIsaxnF+8OK8SwMR4spDeqzPueHWW2cCtVZkJnV39r0BSyD85y2IYdnnta/Upq
dM4sAGtBKyaGp/YWxTePodUi1O5jbcrwVyES2ebjifilYzERdA2magrJxorFm5uq
HLpbHSJCFYjvJgVGXpoH2w==
`protect END_PROTECTED
