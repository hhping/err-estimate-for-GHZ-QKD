`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DNkdsi2EF7Dtlvhn9XX4g/NGClNFQrsOP/Leqswq2wPxpR6RDbrJAvp9ovIbLHkv
rSb3nZLIR4z0ViG8mLQRz5fJGIN4Iyv7GFyZu2jYnkiOhHU2QOPmQLfjkhINvHAC
3IXArL8cd61XqJYgrh/n8XS61/JISWwnf4hZgTewAe7zNFYO01OU17Kk7Ol9YU/y
ULkppRV7bLpK7dmvD39tRR3tH8Qoab8b7R4UkrhQWIHVW1FVpRImENESMmVgQJXo
tJamnhfvWmSm1RHM7qHUjPBgQ1+wWPju/xTayFxeK3qheshcFS4tKH98EOm//ISg
K6j0env1G/1OjdOGxFdXzE0u/SdS4Rud+T1W4B9TOKlOXPH2oqQkCx7Kt4S617LD
urgiqzQ0LEAL1cjUNUu2eonR87nTdepC44XsH+k64YVNjkZpZri7wLQEvqRXHOi7
O9LJDNx7vhjMrpBePpS7H7WpYzk2IJbS2YJ8EeGmlIjdAYThy3uZ4pNqlAKczNrc
KEhzcoiuRmrqSIbKvvMVsZfTLFrdwh5pHO/1TauLWPV9fHkktuVSaAAQCaJXGKj9
QYNOi5ImXEL/D3hP0CBrWOIW53Hatnsm/hsAFD5OwvM7mvKaZDmq2cK+/VziXXJl
Qw/5KKddp2tTDhKRCR2RVILBME+Mm6s8TarbAaoSq1PLrI4rJGKo/+qFSHwqPx3r
xiiGkUVETIve/2TE6GO8KxcI4xbtqrv0wxqRaSgQOXqTGkmSXOhzdxV9+TPH6Hy+
szqRNerANtvY1pyjpHz27g+Qtf7Dvhx2gUvCnkIDDG0kE7rngpI0P/lk/l9yJUCR
`protect END_PROTECTED
