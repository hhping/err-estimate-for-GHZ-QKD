`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tNhtaYlhzId71VHdAcPeHkr5wxryqWbo0EK34iJ9cqaA3BKBeubBHOu3bWhEfp1n
lvKUJdw3OFOyQyVJ94KumdRjESCmQbu1bbTnVdQftJMD9UrPVGuty0lRbyviqjaq
KRDIiJMftxaASdyQtVnDzEdbnz3u4RnC/VMW4rGxeFLaZ0UUlV9rvhaTqXLfF8Fs
GzqIYU6ElQ4ae74kT/oPX5Cmtx8cpEXZhFzu+U7itH7buT7te5MIX/XZI7IiOqkl
rXjJJBsvjDhCv7RmXVIgJZYL32HnyCFyZO9TzlbhQoXkdhZ/dP4b32KE2udg7xqJ
2LeYBiOmIu8HG9OBo2Ls5j5TAEFYgEWGs6prvoBN4nx9ms69vGSMnT9bR7Bz09LG
uA31RKXmGUysYasNkd50nniFR3yJQVEgFL/BdFBfSTcqNpGUZFxdsGVaDmtoMn51
`protect END_PROTECTED
