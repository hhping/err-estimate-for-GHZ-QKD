`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vj1Kpm0p+YlHztgJMYENtDZD4HbArVNpPglbLp0hOAXoAZ5cNEYa5aTieaAoeiZ9
IDcXWY6/vbnl8Hh3mnMjA27hESCvHupBmhsGPKHUj1+HKoEMN1kMNI533xm0Rbsz
5ii6ctTYBBZTnzCcZJNMkuEXB4m7WYc5xXzt/oFrQd2FSH+vhBgSP1cgd4Qk3l/u
AnerUmUFncs4Y7VYlndv9N+o/QyWrGHU2+6osa1yFjBBcIcMXSqvGiTJ69Ie3JoI
dSJaWXN2kKq/vZ7v9bULiBRZf6bJV9jVeeIXAoCTDkWJ2gZ3alRhkK2bKrvmxQFQ
RGtDOYUePu+sgz2k6NS56PTn6tcTgMUNWED6Gx9tdHH8rlcrT7cWxALzZSCjlTxJ
B5GpT0D//p5kGi/TJYe/97ASzbUw8xThg6U6/WJL6xc98KI9I9zA9JP0Si9yqQ9A
hLMeCsxIZu5qquGrjvpiLrPQB3gKD788qNUaslQUpMDgotQmTr0hREmxepC/S5Ln
pxsKBtb0gn51yW65NSU1TlPRyI3HSv73weFSYYOnE4Yk5EbMoRvXL82EDBGgYUvF
fRXx4ErD2HteXxikMg70VB8SjtQ+6t3sx9GtznNNT/eWGrX8NhDcy4KUvOkxu2bs
IJvAqsUAXE6mNEz97nLBM7kF6qBygnLnmwopcczJe/bTwPJu3aN1wdEhJFXe5sep
AkWHV1Wik/sR/1rX/SB+FKofrmsNftOWTmM+pBhXXkilo22efDqnXPIPhKn4Hrm/
5/5z5t74E3E6vMAaxg3DKb0xGNu311updsoaOjYzuEU=
`protect END_PROTECTED
