`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LjE7OB52ftsT026S+ROpEQ6vDACM4d6NXLLNBBJl5T1vaHgAgzhHTPhmJu40qyZg
jmCBs3x9gAhRed2pSw9DAxmYlvDiPCVpo4P0gNWU0nDlDtD3vJfO9out3pc5chlr
BY0Bkovd7yyn9KgRv/cu/+Q/d93cYpVPujqxlDYXFO4YFm0SAGTHna7Igmz2+zON
v6fASvNXrAZwfEZT0v9uNLIGy2Vm22YL794NtLhH35A4VTjEtrjjATPml/YHN9WL
8ECN1zxrSRBIyxCErHTDE2JMloZl29SOJOMxGXGsZuPuPZD/IU5S5tRqZoAGT8av
IDufWV4+Lx7bl4oJFx8sqK4HGEyzkIbyfsoEFiXXIcqqc5MBthBbzZMOtkzD1ZE3
pG88xD475CejpZQu+sttjHwZkcFsK6iYlqq2MFhoWxGqtGMDmM64QkkJq/T3WIX+
LyH2bAWCGbugrUY9KFpBazuN12CL92NF0VC8VwC+0YbNlcHZKPJqBTwAGlbevidy
7LSVJyFf+k99/Bx9Ri7PdRAlPinqqE61kgWP0fmRBivMx9wJbpjEvpKlUdqo7+wG
Ivf6XwPBMtiLGig5MKMANuHxvPYxBXDwh+Y3RL0K0Be62oXC6vBjOFMWuwOxjZHH
cq3JxouTbx6XAOpvdwCCp0rW7qfcFqkM9BfzRNgx07lRCl+RApDKHAPgyexSqNvQ
ctWDvYTEbjX6Io7fNczcPdtiAtkougWibjOH3qYbtKE3BRQT+V5t2mFuOl7zqqWe
c1LarMaUKfn1OuB6yKweNZGiwhJHgF/JEuSbpRWjB+th+OVeyX+aXVZZbzCnVDdZ
Ehlbsxxeu8vbpxaGPn32nYKC43EHaOhM7AoaIZ+cObestf2dfmGBrj5iQQP45q+O
r2WOFNKd66C1L4idFdfcFJEWoGwTCnYBF/uqafxjwbkOdush+fn1tA98UKfZVt7T
Q5fLo3GFOO9ztbU0jlKr4AXhwnQpXhPSQG0G6xGgbY+VZfpoUVkQu4uk6AFCn/m2
LxIq7PFCOBsTvMfJcLztsEDzvKiFVMnM4AB7AUWglNUK+HzXQXMlVrsnwKMWfK5+
D5AQEKiD7rTtErQd0FPQQwFW/EV6Q5Y+bkxguv6YDjloY9sdx2ZOZS0GdlgQ43Wc
M8YLdc8dES8TJHh1uQt/Vgl6F8ArTwFt5we2V4A22iOs03iK1Uey5/k3eY92JYLu
/qWcwx3z/QgD1qNtVwZDDsDSpdwSK8YOMCYmT9mofoWcnIJkAx0Sg0tfeb783UGz
8VFCjRC5oT7eaCrXkHVkqFO/33uhHfWWewqVGJdtQH/O6lXxCRoLs81fz1cF+ElV
MnT6hnEXPhV3e1OKuVgdXx8AUYIJmKSpDZ7AJyrGJB3wMUVvl+YICUM0X9yRYawH
HF4LbdlIDJF5keRcMl6/N1rVul/wV2LrjWjfDFuI9x/3iegFYkBARyRxD9miSywF
tqam1etydTmtgr3h159T18gMjJL0u+yBq8XFeyUDUgrZIDZDf3qTzkV5tzPrRpXZ
UJj7Pw0j7VEivrZ44c+e5VYFJbCnFnISs9wMCe02I6YztR+aTVIWa36UtvAg96xD
RpwzILrR27j0wYOTrByCRvHt8MvcqQkjge1RdyOr03lSHeIjkIGvalA5G/ydQ/oI
avlkfdyPf9rqV1LgqsPsXpo4ercuV4rxj9d0d+cQ34B58RG+/krqe9hzF/GqBaCS
lfcfQga4HOV4PBmuglR8sP9BmMXArDkK7tznhOYkQtshtdwTUSsIaJx4mJXWcNmf
UBzoXg10fdhSPIrkrB38HdtWrDAYWqK2+Le+r3Lu/qVax4IxmL+QlbScekQa2X/F
IJfT7o1ElpVOg/HK8bX0Skd8dWJilmNq8cBOJ8tWPLxvdwNnHsuKfD3f3jXhxssb
crYXs9Bp6WWjPlpBu+LEb15RGJvRQYscdzcuSaCFkbWHmaJBuv7wgsjrX6CoZ/MY
ijJKPqn4qPgDr/fN6fzif+8JikWiGs1GfuyRTklq9+MC9d/kClPGkGrcfEPsoPNv
E6zeBNhp6Csr5fejHAGoNR9XO0z8iMToDxi3Ki5Yt2uDIXIqDDWe7s8kMJdXXt2V
ShhkUoqR4HWDRXz+9XjRHXP6G8gaVKAyD2Ctzf8QgoCxZy8mp/xUuAB2V40O6iQq
aIQk2/8SZWYqgPMCYmQKV7rfS5a+LQCy7tEZeccyPvUHzFPVSCXWq5bQm6yea0Ni
f64GcfhxdUnLHoSnKdVEvMgIFB7cKpFiKatx36h/l04gnd/xlll2Pn1Ht5ZaOhpu
JOk/M+L9UofDsQwIhph/nesLNmDvMEBxp1EVJFwGzf6n9vxlbWQ+3b7o9n5pj9Yn
XKBz5sd9kmrUHkhgOMiZDlKbrgur7O+560xgIeTwntHIN85sWqHHPjb3tCBwmMGA
G1nxzDprCCrapfXc2A/PPm7aAI2iSD6kdGZOFq5DIGjdgiUmT7sLYyUVIljVGGHn
f5TLYThIQKVyJcfIHLxB8T7znmYe8+4qABlxOqz5ItnXjrbj/8ObsrkCGR0m1mj5
VsL12C/wHc/WW/JbaDJ10Z/DCHfuFj88702nR00NXMpap2d4FLFJjHjYtndRPNI5
kp1PsBexnQTrTmR0RZiePgBHeiMFKkEkZ+WRxPQxWV9PqHYagOje8mjwnZinaWL1
tZQLSDWrtybiD29NUpvBrig6mYIgVeysy8sP5N0Sha6UAyqiuLtv++uH1F42/kx9
QIMSsWWjV28rfKD1r32PjIzOpOXTFDlH1U3Fb8kKKtI2XGUawqbQdDlOlXx7e4uy
y0HMlB9G8V8VxxBIgBL5x5ebTfIVpY8GdiMr7dL5AVSmNwWzuGIQoGP2LXP14UUO
uFo914E51q4phZ1amZ5CzHcBhNwipA6I7OkOUwDovBo/Iqo89DcjtZgcWidOuR6c
1tLPDdYxn7aZfNs57i9ukB5U1Lxcs6dNA5sUfASdfF8Yg/IyBM7qsrGi3iybBKOe
NrAQlYgAFwaHUhsZGf4IX4bH6cD//jIDYNp2x2TIgxmm8uzxHF/nbiVbdo9HMWyf
vyVbK8v0CNMgcqXOvs0yYm0kaLLgs/VJ4LE3/eYk98sDi68N0QsyYgyZdEaydnW3
Nu1MTrXs+ZLp22YG+EwOTSIggphWmQ3ere7KhPbrCasYNyP2W3BgMt1bVY9wJlDe
16iqRoFG4AS7erfl+SpUMur0Jmd+Gi0E+j8lINJrCfBsSGeBfGxhGzc86uD5YDre
ALZJRGCfm+q7Ky0VV2kTcOV1Mu2UrSeKKEf/mLP0Cmz4m/PsmxWbaXZbfoNLd5cV
yDBId0DQ23wdMQAPD+X9eTws2Q0hHxEg3VxOHVkj5cslvrfxcOWsNKWanHTQsrVv
4WrlzZvt2537iwYAkL44spGID4PXD+2wPA+RpDd/W+EdDa8vU915YXRIUCerDvwp
i77X0cegpMvpWHCxlkudPWox3zrFih6hLolUNzW4V823nuvrF9nTjE086fakbswR
Ddxf/1D73qUaNKYlA6GP+22ycgJYlHMV0yky3qPHWffHsegucPnyOlPMiOUTH3jU
x9rKPJfgB/APv+4WTRr+FXRP6x4VMvlntsldkdwLOoFR+DtlQR5Yk8O5YqjJzH+9
hjf00a6ySA/jLX0S80/QLh+yhYXpSYJvnYr8tpYxzNNWjovVXmJGSbj6OFDGh1qK
8R50IPzvaGV1UNkhShjruTVHBO+Gu+iV9WcJYQ2Pds/iuq9QVMSt8i/PhbAoa/Ig
eBt8ZrOhCuRDS2jOiG3vMoh6D3Svba3kUHb1r7WhTG1FxBMuVk1Jlq6ZfgsN2yAY
pnOZ4e1JBBtjmFSnXBKQ3BAzaw0Lc2OATsPvIXxb9BApcw4c8Z0XJBOnkAZlyeo7
PPPPzzvKceWsjEmfcXIZBzewcOdsQ6Ff3CI4RhPMvYyKIB3cCZbUzV6VQsYjywnf
f3gZRr7PjeWv2HbcudwI+AcJ70mBPznptW9Zz69CJFhZ5y5x9RGYYavarHYQ6E/U
pQL8DIe3rV2Hrxy8skgx/N39seHEM1u0w4KG0ke71Sl7A4gdWk1lgjYeaSWAPbqH
a9a+k401lmYW3k+UFKEMAWRqXLB+iUBCV8fHLXwYU9KNXrvO0FMEBUIrgqLDb3zk
Rvzi43q4EjZ5+01hAJriQW8UXAs7q3D2I7wVC2od0RcuwQ3coPN5nG+o+RRlavxg
2r7+45DW/F1PZXZGO9qnJF5aIHJYs7vRgu9ndVqgJ72cUvd2/3vtWZSEaFKxp+lO
69eM2i2PjLl16VQewofzNFvNxlNUvLmRNM+yovA+6RPf8bNNnDsezCwZ/XHFC7ZD
UZCzW5gCZGWB2kn01MDfHw5zdfIh+hdjvYQ6+wCHoWA4XN4pXsFdAoq9bHsyhaWp
WUGMaA/k0vDJBMZUDZUlstQwZ+uVJO9bWgmdqH6xvIjYQ5xLlb+tagOhc1pHhtzv
JhmLmmff6m1f2cle5eQwlvlW7Lw3iNwSenDHjGfMYimPVW2+15Z7SuaHA8Mn5fzY
ENbq+ZiLkRekiG3/6sSDKH8LOTxiJG4eYTYNhD+0Nw9VWY2HiNdQ8HDB0Tt640bz
rzz0Ufc4WOp7IZSjwro7m5SE2+Vy/mnRAroRlTCf7gP+a/aGxsjkEha+Ih6NELNP
4KCKjiWi1TzXuYg9R+4rGULEQrSLRjreBmcSG3l2lskK+9Vb8kIGl4GzdnlGitFv
YOD0v+/WOoLTbDgjpVEKvnr9n6coNodYnaA+u6+VGoOwun0Zmm2biah6NuZgtmDw
QBWCWCAsdUu3XtPcDIOpNGAnKeZTGjMUr0pk6L/KMA5Gaz8kTNb/HOEJAqKW7Kt5
f4qX1WNZNtR0l4QlvZqL9WTgieWFMUiqcWne47SVfz4oGBI57xyJ3jkanTi0Prlm
Vo+y3SIAtG69X3m2BM4uJwZaYa6/ar1978VLzG131AsSLpMC1VsWMi9v20IC+URO
+j5skner/4XVqUL5DM3cuKctQb+aVCJE6e8xE+0JecZP0hECYQzhmQNntQmiQJXO
esA8YOX40V1po1ucDJa/Zl+3zcexh5v3W3qWiVic87er0NiNbftdYgGbqRbmTW9n
brllfCpipJOwP7k7MbUkVuoD9XjNwvqPpjyBuI4iuCcJDGNKFMk+3n78IPmswoS9
ojHoQJfgjcpkTphK+YteNx9UDzTfoaQyb/E7mYzct/7Jk00XnLCj0oExeQK41dHX
212mL07yLlrcNDrolDxBDULh7oQfZTrTnqTZZXMna7blcO9NVghz3+voj3bA5s3y
YNLzeOuQv7GByzlzX7KYDcIMopjOcJGj+dYZi6NYLS6bhqmSEjtL1geXZ/RlzhSD
4eteo4zQwjpUlYDn+AdxHB+iCcIi01UoBgLDBYhsH9WrV79iiTSCLR1PNIEt/EVF
pUvbGCICE3SsJ/AW7rCh25+UfYzQx+waKGlhUYN3sN3cy56SxeTm2EHiT0pSfY9T
gk4KinXiEUObXAKv4zfGBO/Kw2Sjd1jyRPCc9AvkqqTHkcc0VwXSyZIiUqp8At5v
1Wa2ArVrG81Ks0sRDalAc7Bx93NCRfojhxwqUSeV2KzJ6XWwSBFEHNoqGXnLKxZs
hc/3/YAvshbhXsuOncFccCdq+fSaDElCxPH8ar/rJQtjVU5uHS9aBQZcFcfkNxrP
IUKG00kjv7g1XbqdFkBwb15WcRbH14alRZw1ZcT+JanAtsfCWN5cPxSURc/H2Kp3
ZOpc4tuOWqeG+/qSOeMP97DFJLdq23WpNiaTW8BfD76u+Lz/uc/S0DaLTClO9Hz2
br0nL2R0dcaJjS0IdH98m7DTeubSiVQc2R3x087uH9CeRta0UFhFQ8xY+ycQabFw
ua0uTZVWBi7EJmLW9EaIVzFx5j6A3IPU/eSHnHbHS9GHfKuG0L6rCcBoO68Xq/Kb
AUn2569KdM4q+vugeTReSU0mW3NCrywVLd+4PQa12AtJlVKW/Yq59wXiVtIoGaUz
ikU1kHBIRbyIVXRpR0F4kWE/AocC62Ggr78cCi71SzO4hUJa1/LhihjTmWzNFtFH
38ifCz7cEnBlSx+p16/J/DgCSWiRUhAwrQaTJ7HTkhucX8nXPcUT0Pda2mW9Tqgt
kdyrwAxeRSMZZb87kJBn55EYLyv70EAipmKe/eg4GDWk24HNI2GrsRTCjHW+YzDb
fqzH11jafrVN4xrT4jMgzxbqrpGHHzlhMBl/Gr/tVYbT1D20SIi8essW0qVeLMei
7Ycok+uV1ey1lVUKhbv/yNLMY3C6EAH5AM+3GEfGx1R5Qchmf3VNZJTtWHkuSWIq
7U4he/yoY6rZfykUNt1RpsdJ/Y2sjxrFoomqNSLyX7NF+v1XzVxor0aDLDvel6Qz
dwoNHIfdYx/hbmUQYSP9WILpVJKzrl7tw5pufrvZhBsEpTYpajyoQo3XfHQ+M6uQ
dBxUxxmefW+5ZzLOCRpvd9wzpJtRWE3YhWJdO0NOvSW3nmdbTeN8qQBhVcqCt/qS
L5N6Re7FhRdUD5OqJqCvRDePW82+Kj6DYq0YvIpoI2xcE0Q9XtLosH6+HGEeBXGE
tz0y/KwBbj83XNxJtcOC8HB89Q3B/G52582LhnE9xyvdNZR83IhhRCGa65l+VN3L
sJ3WVZ016vDi60zEG17fA9gWYBtNcxNjsjx4tCRh54+FWtKJvRi3lyMBTZk8KPtO
gkru6hpzFTRi+0MxRz/3b8yQdFRucywrUXNRQ3O1PGeKB+I4CNRexhk3XFyzX4F3
fmNZHgGNA2v7na7hZijUvxSv1TKUtukUfvy4zAzQi+POfzxfRheF1wD7H4gGfHGx
btBbdw/3SjzPeUINDT2aq1BzbbtmznQspBz9BwFdLy7oDKt/BXixU4hsnvRMwlM2
jOjBOPxCn/SO+v7tZ0VyU5HFYhzL3Zry7y+EJEO1TR3n7XH3Umkgj4dOdNj4djpP
ERFYaPPTc7dKaeSldezy6iVBiGuAIJ1iLFI0T7DoOES8p4/GNkf12HOoW5/c9bmw
1/+vw/lrFDsJMVVo/RxjU01JvICdxcM/3OuHmpqb7DiAZiBeKPBjLYNlct1dIpoN
YtFjBEiQ0ircI2HuZsKvAKCVQzJWBIJgeUJXJvDYH9rWVWAeByxI5ibr3LUA+xwi
MxzyfacQRfQztGs9YkafNn6sqZpDsQ89tHnYrH5YHpsNBJkoIj+Wy549LU92L717
qGFvEZ628TwQNpiXY3OQzP013MlBLNA3hwXo8ZIdfv+B+W2DcMxA+AGtfrTqIPfy
Hbzjk6oC8iLtyfWGLcIXocRTGHLrRb44Cz5kMb4PyY42oQU8nvhxfmiGoxNDVLjG
NyioSgOTE4c0KI8CWP7CSd5rDHvf4Lg0W/zJrCLAuzxy2/RASvInfDNX/ioOIcQZ
L/bz6x7Pa4n9NLQDFN5FhfHlFrcdBDBs0oqU2eNdr8Tpp2ztcF5q6qbRqEaY44dA
dz8jGCzqELn3pz4EPNIo/JgYV+EcUHbhc42EZ3+lYd8pl+CgOy7g2fY8Bkiy7BUM
48S6deeS0wF6mpsn5TRT93obddRxb6dcC01bTTqTq18KUj94d2XrcHDoQ+jk+Mhk
dYrZ9635V4vNxfkXivAdo5PwQQYYgFlbyJfxY3TXHrwWROobtIL+TlUzwaEvLtaP
XsNa5MiUTB5vyzZEPtDAo7jibEdXOtWkVv4OJiIA4PddjdpVhxXasCX3lfHHQReJ
g0dWbb/Y/MSQsFvkWb860sJSJSwaEpcPW0BO7K0MpcsBnjATsE+T2YzkqSgxn5H+
EJerjqu8Mj9wAjwlj/XLFCN8q1O/YtWJkF51ZpveDWtEfWMaPR5bAWCrTCN9g3Mf
GoCy7Yfu03oY5C0GtnOioGEcVA70pZ/nJxnP5SnEClObmTeEYmhlBrkjjiuI4UV5
YvzWqRBt63IwHQy+9Ud2pCo3JQxtD/hdBytBDDzNx5hHU/VS18gNVP0j+Guv3tqv
ic0eB+8lvuqU5YSBwzagTHYSye+Dqvf0ghkvRwuBjaCBbdVzf728CmrBaMytSUj9
R/f8bID59Q86CabQ45JkIjxuG+SzFzSQZ/WUejB/YWnrts7ILJIWEQIhXI1LZfw9
BPNoFfmlLCVshdydSFVqQLw5RgS31bWngSMODL+GOI0FkDK/4weZl/tucWv9YCEh
3tYjMYOMyY/1deZi1OECcezfcme/yKkH3yvPXHR39/1mxDtQBQIWYAgwera39zeT
u/8ODHStDB/pK04a/liENmXQxmmCZ+EmlFegeQ8FXEwhOhzl/SMZX8NoyGoNLOkA
X1bf2bRZwb4BUQcvjupYl0IStd1JHVQ5knyi8PE/auOcLtMUL/WK1r2TnRqSKPeW
g4QLpVg+jhF/N5owkgUafMfo1Elu+s/2VTz6zbBdAvH3oV9Mt4DCVKWftwHj3Etc
rNFzJpupc1pDfXvMbvhuaBbduliYVQk3Z+wksylJPZuT6ejiRSaHoCKxpMTdgyNL
Xl6LAg3/Xwxroh8pN4sz9ofnOn2NmAvvzORY5VXw4TQAqu/cyx1l+xisRiJgZwkn
Kd8GQhzB/0+nEBPzf6UMWUBiHm6ViGIZr600xzPdd3LEKQpeUSrNH/a8gONG3993
FhzzZ3EEXHGCtrs+6iQmXExHrVojckRDeDvFRFzLd+oy50yd4GnEj9pHRPrbgeCK
FHC9PzSE845Os8NeMzrxZFXoDVyZA+MFz/2Bc3gA8/vM5AMx/hVLWBMIQqj/vxAo
/8h7z1RXa2VfPd7dUmYCY+q/rzlwB58tCpaafINP1WCwraA8zH2SVkcJSPS8Q+A+
vi88QQ6h0ZbHCmf3QHKAM3CCgojooSCRXF4GH4/aa7EQn/knw4UknlHoHuXJ6vDZ
ZueUH/wxc4weHcxV/wtpDh5xyq0dRT3n2++zK4fAWOAQ9xfz8gzz9xq93rLn7ZbH
iOkFQIcv/QcNodsZVxZGPhFvffwPESx5p/YYsUDGrN5JIq3wwBHoUs9/SudHsNp3
vDK3aS1ScYZbjUQF205fhDYF1nf6rYSquDfDpl2UWyYBo2SUXZp2SnRd+Z0CD1VZ
ly/+B6itmD7rmuHcOZqLgle25e7dUnqHzwfzS1occGcoOdRNqlEfGW+2xUyzvvIx
BCEZouhyzni3huCoTE3oXiZZ5OllJIPK60Zdowg/kHq7foVkejcSPfJX/DJ539tz
9zzV2GUoyIuQgkg+ddvZ+FsTOici2VZjNsX1v9KsX1qz0CTrXUZy0eFQg/Vau3lr
XobiWR97M+X0mhqvNF8y/PQObqwGFuxPpSXEAN/O+SY8ApMT1lKOhBW7tpbDiFnm
GckeyqpN8+7MtDDy3aL1pbWlzw/dFvNCn+TPc4oUrbHluAxWaEft84Es2R0l6H0A
QvvbTMjF2oVRGm1WOjNA2I+nAjxVdVJgoQ6bT8L2Ukpnctn1zq+2P8frPomMNfUQ
GCcSKo9FAeHAyzDsc09NAhS5n5e3eabCRIwJ6qtyS6ZjJD9zOlb5SIwha+F261Sk
xw28l9uVnlXyJ3ixyGlZZfi9PDvN15QgwnbQqTDUHx5+xI9TVR6Lp4ZHyBWgP7d1
L6k5wMBGRrYEgFMBTl64d3DxiYMcubUSngR4y7Yja/ChKpLtxxjvkKydrjhtaf4q
EQM8SxUSXrLsdbHdxzyIk1oXRkPWZr4HSHwjdRH2LjMFNoimH/1R1tPNJR6eD9s0
uF14WxwW4xmlB2uIJV74I8YJsqfhpE4gX+56r+4AGH7ejAJqXVCinNuW8NuSqFMw
LPzxgE64OhlxhsqXRSX/z7JfessK8Kt+lhrHWbMNm7pP72hR5F41/DwaJHjJvLZ2
337kGu1S+ijvizNeWwmsgVbnCJLXrluu5Zn71osipX9xshvvztnCtm2fKHdZh2q/
zQB2Oo1A+AqSatn6NOv3Z3epR2zpfpJ5/EZgpHcrLOnqPnV48DzPivniW7wnRfB8
/R4WfXjbKn65krv8Yfwc8jGTL+BBZVg9F+lJX04h8Aw9q6TfjbEEKBfcAR0IHNYm
e9E0PgN6aoFDKOuYhr4NtA6fjxFYXJxL4w4mCSbaqR3sFBQv1pveV3bqCQH1zigH
ZJ51L9AfYXYDlOU7GXAw4P/HiRKy7/zQXWDBnUCuOg4tnSmEWve6XzysH80++f81
VQfBH0bPXpgGAXVBh6P2VbwiPBEz4DY1KXYR9YTZ+6L4qd3qae5IGC3SiRNw8Tj4
V91XF9OqLQRr3EAAKzr7xHq5JsTx5WmU/k4FjUtInxtSfTs2ddogc9zc8QQbnCrN
MSFJ2Gieg4Mz3qYaEunuGdhxbpx8lzv/6j6gKr4PiiRAr1c2RdsAttKnWjW2yXqE
JUnZ0hTBfUPA2uTITm9Go3XJT1OTrO7iZd6AHk2un+8cwEENX7p4YFW8/pF0BAr3
Ngezj0iv1+Pal920fDTQlAyVctVHjA7TXZ5/5QRf5Gfzfly5m6aanS9OmOsWlqCW
7fsIHheh/2mr5tLB+3sL3RvcLUpu8IwYqzqs2HgiNccIH9gK+N9b8SoMzOBKFFPj
VV9Wq/doIHV2h43Feq+aQhLpEJR4eqycVMsHdfPQ4feKth+y4dL2q+SNv3uVo3Qs
n5GqxduCE1vqKPGK53hAkufg/XlhIYuOFomICVrii8SrRInRuvOVj6qgI9U/ohlX
8B5HNUoFnVRjhKWQ5KrmbDftpRSZZUfXKuIiyGuYaTOuTwCpT5QIAEMjzSfWj5+e
oPZkf1DM1Qpk/aToFAkcz0RTS0P3kwaRVXO5oBR6EDfc3tF6ZaizhBdxxxjmV6J1
ZSv0y9Xn8T8pc+pc6uztLzOfrHWVAggPSHLLR0rNvgDKjisLH/Rgj2yo7xnNnw1m
3HuEzh5RBXoRSWENmD2SSl+ItFnb0Yb3cJKUopD8Rnhm0l0FcACKPUx6UdZCJZ6E
mtFZFASH8bXgBtzzqLrFfoTqlaL+jCpHjMUuSRVD7mZD/TEh5uLg9y/TF9SwtvgL
bVKFOR13C++d1aGZxqeiDV/92Gmm+etjRBRbUfXzMgal2MEm5KiM4Edx3E/tVNf+
rCzy6Ho8UKlADtFTPH9bLslwb6lHwWWQK6tjlSrRJV4HpVyR3Tde0hU/1sQiqmBT
5855cdLZBi1fVuss9CJZK2Ya/0iSjeCHAI3kEXtPAbRoYgnkkHBUAu/79N8ajH8S
yBfaTfqDjwthqK0pg1glQiqf1P+5risIyezNnafhwZ7IH1QbciqvH17kqgbeXqsy
EHmRNt9ZWRdP43bUhEc1gwnezwMDJCzXRCbF1U55UadGuxKdzTPlWCGXJJLUHnPa
n3bXkzHo1cooSYZOliWwDggnEnqHwR5azzjtXahHmuBX6rXp4Upr32RBuchV6XWO
BadqaQDXX4uJX1vS+DWqrG1y1rijkk6OCQUYBMusB3TcArfWwQMoPdQscHJqdTCY
pbbNfIYtLgUVfmJkWjq1fp5IlPDBeLtwQE9KHgtKIhCxytYdbljeMisEfWH2ejlj
T5VPqVXRNopNIYeOPMzNxe0CxYD0UQv4z8XWUwIu31Svf0dLK2FgVPzfWkdcnOcq
Bb0ngLe7iDJz7heK+ex/HFSlqBXhn36dn+Ls8Kl/ivaoJkFlfoD/eeU4WuAjVREu
gA7sks31hPSmPGHfH0nw68pzfPWgl5hzbRH3rEOLpPzL68DC2DFXt5qTkH8p96Lh
fCDSHz9r2v9GJJDko6EfYKiNpw1ORuahjSCwSYMxkMedb59jqhrrPfmQ2xw20+63
3RQ8TLQdc897hIKQjflOMX08jC/70Z85ijpTB2YKEPu+loQlG5n1kviW+QZuhynQ
FLxUYFXEsvoF7kAgrhx32n7qaSlX/lSC7xqslFTV5CysUOBjIc/e27csD0u+3pYr
YenZuBEmkZRG06u4UvTloPSm352B7Qt1NZ+m5jti3NIo8F1rwoIqHWAiVeDxUr5r
5MeS4ErY/PXnAfbcBrRir5SNf/mFnInoqOxheGFqzQK3Qm+7do8SKj/gMktWNofe
x7MwCtsDSCyxkGO3fgW2pCYjgCRnH7mhgOxNazZg6Zht+dEoWWMALfAJHkEP9s0b
PyC9haJVRXS/hJ6TnLfo+mcKukfSgawIYe2hL3iM+PoAK544EU6R/SpIVlZS8P4/
O+ebtdcFh2X373IGutK7GUGYp/1CWFq2F9DdJMINGT0UNhuQCQoBfVvpp+uG9jyF
dgzhrWj8RF4MSlcTkgopi2tDdvnARb8TBHcaVCRfRbANtFyTFPn8bemZszktPyiC
1+31U1WGVdTOSrOkiQPGlXXHsyIB28EWovNLPQLqLE+gAT6VEx7bliUIMy13g+XD
KxUqmej/LweuGYYHclpOKQhKrSKpxBbSS8iQpGAi2aXPBj2vnVxYzF+b1h3MWbTs
Om6i5780OmziEDzNHxskpQ==
`protect END_PROTECTED
