`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lh0expDhy9m3cZiohRUlGtkYAp+5ezj03rPYQzKZhfE+mYCknD6WwiNifeJvWTDD
0LTTFzHAtxU/5lW9CvoicWTnFPTQ2aL+le+u/YkSrx1wGTEe3hzhyY+J09kOk6Es
Acfb3cW9Ki7nVB1yG3wnkTpv8QeohVfI5LL+Oqh5OHQ1Wjb8Jjd+iKkPmXSIIqeu
fyQME0JZqRa/YTTKcGhePfAQxu4QQ0A2NYKtoruHC67KWebDpxbv4RSVJx94j3Kt
6ChpSHoUzpnQXNStGBYJW47v33P/vC1+sOmM1rFAj1tLk1wK4JlM/Gj3PHHkuWnw
ES6JdyutajlAfc/RcODI9q3oI3ELPVjkJ7mFnQ3XKuX4K80c7jLUdFjhmHmY1CTZ
QOBXIiQo2d4ctI5hHw5gzSwK5T54x3Yn91o48vIk5yzbVuXL82/1Dt3/Sm3DPE0G
GH2fMn/CYOLk7TF/wuGNt0OpOk39k/fn7vXnnh7BSDTEg8n9oGTEsWc7X9V1RrJD
H04UrSma3L2RrGqop8T1CQLZ1GVyP02MfwUSjfziEYL3lEd871vD2lLO0Xv1qCB2
AY6lXmFsgUvobD0oCw1roJ73wO/mwOrldk7rC91ICj5gWkUXV963c3n+U7TEiP/T
LAFkWMuGFGkbqdqDr82ZYdqHc+1PUuUH8MQQkuyHI7bJpPyf9+v9xHfMmCghO0pg
/UPcJ9+rjiLsFtUjwk2BMA==
`protect END_PROTECTED
