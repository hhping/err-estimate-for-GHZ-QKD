`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TKqmwRpge+fZxRbosLxgFilqa2h87H/9CesynEpx4fsMMsaGTFqm5y80zfsHQxN9
7MaY7zjXn7UGjCzjoKs4aoh2XHKoGShZf/dE6BHhB42wpNOhUunBajZTe3sd0SCb
5RSWFZRb6IqkCWfq47RJFa8TaXizp35uc9vBbbnzAz1YWzGPx0VSl9zkF+SliZJ/
oSYs8JiKkLZyV7+a4XD6qbiEKBpCOR8O5hE3sYmAJYzkXTC1nCsCAkvVb75A3WcX
d78TvSu03tER/0HMcR4VMeUCj8pS4ZUd1GeB7Aq4ToFp6wBe5yZYM7bre2q22N5p
q59lSPe00WUKU9b+cfLDPuisptXVpeGDmr1rlMdLcERNxPMNsj9lef7wDJErS0r+
q5in5UYHmLkDS0nwGiqbZfUCWOTOPhQGZCbqu5ZqAG0Wz2vHVrr+rn4YdUXOzFwx
Ju2YvW+5d7Pk0LzQVZrduRe9pl6+kAMJEsIIV1p8IwtH+gZNGM5n8NgkmzRgGrmF
/irgc5HWqakrbjTQ7jcA0P0forht++V/TTQkDoNJDw4=
`protect END_PROTECTED
