`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DXQkVSzfEyWBYeHWsbjMcvqOA0dQ8xQSmCbEgjnbIqpd0gzj2BWOgOaL76nD+h3f
Dlr+BLlMZ+Ra4AtzS027Y9X3xqq/Z1K0Ponwy0k5hlOT/Gw/VMnC8BK2YqCJHezK
55mmUxCOXhRt8Bg2tcrl20Yk/NoMeL5Q0Rnxju+tMzSppLv3PL3TBF35rtJAgpqw
dwUPwyVXGuee3EeSHoTEHelM0zM8ZjxMjrqgKc8o4EqWeOnJHLmHWog5H6Apie7r
4h3fsKtMSdAU7YWpRCBwlMlqZiGKPB1k9Wr0ERysfB0TM0bp8suqHjhAK/9MvsS1
1CZZDoHdCxborgTEAfpaRkIeCH8LA1Fg1YEh8v4K/IJTPNjPwX0vt46HAHQ8/i/d
cNAxou6ZUXh1MeVXLSS+h9CH0g8fXkAdbDiN7uBpLXqGJRbRB0DytFLW+Fk4+voL
ScgX8qZbvVcFGkHo0eA8Ajm4c8xkoJiYx/eYDZbf+FRjAfE/5GU9mqS/BAsmXwAm
B7GB1IiKhgd8zA89Rw/WWNeXEpq3yv1HvkflR7zVn93own3eQ1Rgf/2YG58EcpLS
lW7PQA7KRQV5P8Z1rXBTyGonwx0vibeY+cj3VrLK78cYfTG3B8vDd8utDjG+Vtlw
nzru7wydwue4xXNXTNQH61vR0G6H9+pv8nWf+A9qp/g34EqSKEDi1ky0xLLy3AR3
GncXg2FrHHNZevdcsdU0/7TRviua147zshRy0fzt0TS9sSI9k2CJijJrI02fXCGc
RlofcZSwdNKHygUHkzyoCV0GVGY3uQkovY5iHyEg/p6DsEqa4JUIQPeQGkXt7PIg
9CcTUq90T/EHiuScLM+rJIFKJjnziLwiHaQx6fXiJbOS2NLvBOqrCOJ9HW3R8dZH
75wurA8fvjQ+gPuZ30xI1xev04YkcgQiPtsEOyAkb1oQR6tyBfDBRO6cCVK1xnNz
XOwxs1RH47f7HP4FpUadTLAlUIoY2DAcacGj7LZU9vbGsyedZJyTUO6goTeRoRPB
MS2asVwa/7TehxZ6prgon2R5BeU9VUlRW568fHMboqkVB/mxCq+Md0U/XKvjwmYe
vrYg+ul89iwWVHIFWKNPMYKZDuFxPm5d2SmXRsc8qZV4D+O+T6IgZo5jQLo3TGbE
LiZj//KJFaioj5+uz53x/dYare23g00h78G/+df9jPEs0VTKoSpdMieUP4Z81LMF
aV17sl6o1J73o50ajYvIw7k1Zypw6/px9KqktOxu+NPFWgkMlbo3Xlr22Tdf8O6I
7gjHizCqAxAzx9d2jKbqscf6lYr5m1rs9TdD6xOdQwHBPrtUyG1N7ThXkro8e4L+
KU77yESvacF5zsjw8mOj00h9/BUn4FL0N9fkcwSvwk5CEPWPqlaUdVNfNhE+QVT2
fa1JhW3mFGLtbc+L87UPf6h9wtoLNKW8bD7myq/Syz7L++QufDaGdg47YjhTPJXy
WpebNYbaAXLjYs7Enhgr7YB9cZQiqyVN3fxvhyx3n5omERMUnCZrwRUY1TWbj8xF
XkBazN5EN04tfcHCtZDDU6u0qSl4EQoh4HbO7VU84koIlwajCvLSWDWYG6avDI40
FXXAz4+favCbLFZhACeIAghZWHuHA5XTkWiX/p79xQHSFTu2Cw3nNUjKw/9gcQjq
sD9y6cjFZoR4eDS8qRmHIJsrAvRWViXAhObxZvEn2cpGLLgQ3+kjjAKG3nKvL+12
sQnyRPi2OtTqHJt/CFEfzuBpiLpzStvGOjG5ifqFRvtUgFLrsRS2NeW/Cdqur2aX
lh/y0Q207QA2L7t+r5sOGRhK3N+8EsOXjZXoA8MoxGE6Y/uuK5LRAkatoIRNpySR
6BY+rgGcCCphu9oW+yCpgn/PPHHrDKMI/vUZpWY/+xi5Gwdmox/gXKYTi2FWpx94
nSB0U6GZvzuNTm8SqBvXCvw8+ArJxQIjXH+TbuplFhmTm2BLytVNO54Y7oRLNkxR
J8zVmUDbM8+dbbS75zHNFMf9qFaQZSRIZv/JYD7ja3lETW9LsJzJ5UcjAg7UxQcg
OUGct0Vm8bhqAaMEgp1aRb7+YdoNggA3mw7hlxNI17sAiMemCO2iqqLCq/8+84AJ
Kp8aZ78FVEoz3v35eDJmlB1m1AzqMtQ5daaY79eogSdiH7d1dM2pT4kP7X3De0IZ
11JNS54i2/SeARZfA4Yjw3+vFJv0WBpoJs7EYMU4pE8PtvFbJPCprlquWrAw1MWn
oC4yLinP+nSiq/OZZMkiuLynm78q1Xekr6Xh9vr3mubgBSr3S78qqegni5P5rxZA
CL3QtLC7ki+E2xnz+LFPSO/Orr8OIFTIYAfhgLLPg/r7PZXV1crxx3wW0lj47LnJ
NxsnO+YeVhIu9bgbFH9M3EI+lptSlgU1ED+tqWFoNtVRQwauJ89shM9XdO5KzwBI
m/gEUEikaGCARbqWJRloEPwen+nivuF8mcE0coAaiYTev+U359d8u5G1xg9SENOY
Iu524nyZjxYmG9ftbxvReWafZR7oqZgK2ZY98vtuduC41TgjamMLhd/KhyFjb7Hx
rO0eZEgsjyQQs72H7+mKXf/s9Ghh5+P7xE2YyWKvF/USXjv90vzE+j1CwsT3/i9y
GBKfykNvq7U1lf2ChOFcbZEpXRC+h8CARfVqW0VV8zZ8+08G4VygLvYrsFp4mlqV
fKmuAgxTzax7kgS/X7tS7G8zc7PiLrqUE7uXPabD4skyaekThsFdn7Uhl62dWf7E
ERiEjwIJhQIlaLEeq0gOLozLMC/0rwZe0u/rrOjnGvTMGVouIjxKy+DVfy5STWqy
dI4lDyVOAYysVN+x6hYIylwa1Co0FW7P7bVZxpj3TZ9VgTVbEYDjBfDl95AmhFgc
rE+9QlN4vECG2e+6YY7POCMvITcKIpFrmvFLZ5sXYj9uKjGFEetAf+mHYWhcTzWQ
u5bMZ7B/05SHyOaYMRfkzdCdTaxcZutQ6D+Nr5BElwIi7LYVZIJUZ1XMCrvhUC0p
lAKqwfq02HMurllgZwHe8g5lQsZS8ES01ePAYQQ8xms8LxKdDPh+EmSLzL4JoCJE
moxpj8mpTKU8uddhe1+oEdozzsBkyjKx2fTNSRyAGXAA4IWEuqj9EM6EFyQmwRFh
ViJCpYsolGrC1censAmrygk8/64HYktYp0HQSLvrjuf5j51sPJ0gch89b7iyl/iF
ZStGA/E/Or+wazkU7aEYnRodWmdof0tdghxFwC3ijathCHq2H/zJiamFAYdnUcnK
q1PJaqrlqd+IlKbKifKYBiqf8zRMWe6MBdn+36efubPfcA66fFYEIa8couIHswrY
CqFHhlBVXWVoVrlwYtEUCj5E6RND3M8e0hkSnBPdI0SsltITdGn3GRVCi7CSNMJj
Q3bccqgt+kAYP5N1sShcOfPEU/wQ/9HYsMZ2VhvV/kTpHhQ7g2m543tCwaZtQ9Pq
uZr9McU20Y5VuFJSiOIaItaItyr+m5JC9sDIIrMWPxrFwrP3PheBWD8MM39ZBRXC
tXEJXLO2sFJLnlekf2rycSjmWDxpS8YOQnDPUgFy8MOY/WHrOOk5sGz16nuzr/Av
Ws6UZVuEEkoqpS6WGZzdr2EaaTCPOh52TihPwhH/gdP8M/5qLQipF5I0wMc5S5pS
H7itTkg3fThDoaaJsMmHXllXhLYOqnjYOX3US9h/+APJA704RAuIhaQJDDpz94Qv
88h7G/ylxNqQwUJWAvq1O9BG4O9k3e+c4mpWGCMYdGSuQnFzVPjYadyNdt9VTrv+
O5vk700L8Ew5H6oBUNbgRcIpwuqnni1TFFzhXM6Q3Dsd8j6W1Hk2y8mgD0Yx6U9E
0KPxTOJZ7PyoPLLL85X9xbU2riIG/p6sEWTZ3vBfYzpDeJr3ENrFGueSME/5q1UL
ajhICvItjkqF9YRT2VkGLibRq0V1XWANVKrPYCT98Fo6ay8JUTvX4ig6g92CeJE3
1+6R1N9TzmXzgFdBOAp6fYSoUGb0pVt4rYeXJe0dk/JFgNLWKfcnR5vYbxNF38JB
k8lVWHBXT8OqVjfIx8LkIcjGGoCzmOWc8S619mK4m4yMw2szR3FUj/8xejtifxg+
AC49AOFNlHISyc0fO7iHV2EUO0VuM/Y5eqIMwE9hbu4R0Cqo9VHcopUrGXqlU3Ko
x6sc4jIGZWut0vUA+/mdl/XGu/QP762xXGwwDod0aTqeeriKKOu4ROFzU8vjJZyZ
tArGO1AHSgPFevdbplgo7AMWMiM/GpHSWePX6OkI1n1OnLfhn8Omq/vbswAzkwsQ
iHgL8yBh7LVXELvHaLxEzLxiHMLF2JRGar2s02L9GGJj0kYmsgxqmR3w8mDfwbQX
e/EHis/t/EUVCf2Qy04WG1VwpvLTFqvazkBDAJZUBLtbSLDcAAX7g5fKkKfd/KiW
q2710sDZ+3binzRA+keTz+USSbn6x3NFcSgMpaOkFC4H8e5jD3wESz9P3x2St8vs
BE1QAwKAOfmhCrqMuTM9mmTWI7KvfE7z3Kmf5ZEPSk/+fdpcX7KP6CUCLGi4On1C
vElXFG04V5eguA9VC6Cy4cbwaO6YBM+44irZ7nP29WCr+VqBb3EbdKjBH7d2ju1M
Rg/I13YBf1GviO+vTGWMSguEWqvUEbHCBikDHjQGb2J+EAhXqidOOqOJLWKE3UtD
7kHGDsWLH379a3ikrTPoKWGw6mUMNUb899T9KUm9H+5lU2ykeeokvQRStEqBwVB0
ofmmmeA+QdJUk9FuFjTHimQiJxfqmPavn6R8g3IbVeK+jzsRy65smSmDQKQosqwy
YiSRCJf7WeNaWZ635rWTF5Oys/Gbns9XJX+F1GeGvKzCbX1hMUKg64zGgmg3afv4
YWZNf+9JdagoEO3dzRQkuVGGlgpLNZ+leIcerXGnzbEyEj5TCd2RbEH74rtzlGBA
KvTyNQKfoR7bM/nShx805JgcvE8EBNNA2nNBUJRjgAgjRKdF3tb+9W4gNfLhfqCK
cCd6mjC0aLg/sRVJhfTHZyAFbfyo1J94oHhjmBaD8rlGO5E6C1tR0rw5p21wXXOA
8YABnifu3MBAy9owReg82cJxHYII61WaaW/TGfZc9dt85roTwepspe/dPK+jQJgV
aEqfdty0LAZ7Qtd1x9GDEw+NvzdPbtVvTnsViz/cuYIf5nfiLXuDe3IiozrCM+9M
BnLCWMzgilUC3CYtTK6/kjoyatyfBWDQrGnX/IFfS9uXz5J7DOgnbGIv+fWxa1K3
sV0JdfSQ2wgtN4Cb7AP5YLntxaedzOKxjnfbzA/9uCNw7LOVLHBhixW56K/A6XTs
5UJdtWNlxEfA+VTmh0idppXujVR62pnxeRf7MJ3liyDx6sqNyPN170w4oIaRc4GJ
1VnxBxNaqlXpS1iSITfutHdYIRn35bBz+nGXh0W6kqzvWjxCtslkTG07//ti1QA2
By1qNXURPrCf78xM/Nj5fC25xd3wnrx9X0M3WutOChLU0Xaf3pZo7wnyYH052ObY
Tw5Cpu64XXDNPNMUptwpdfghZn3qFSZ9s/IzlYY81tG6GYb4ZMV68jz/tiYdpWQF
U14uzQ5xfpaJZ9SjNc9Z6SI3lrRr7c3Jb/4zDk6aCpkHRB6ceGYrVxEWWNIAzNRg
A4q3Al+GtlRthvaaJJDmGa6ZN3wXKf1yAOL7QsTJo9SsAyhYrFNnPbEwssKHltWG
4jrNrEUnBu0aKKJw2vjk74sStgX+s4fFU5jD07oKLZ4IZ1b0gJBGzaPxhgBT6HWD
7wy7qAKljCndm40tLnfrQxpIf4htmaQd+NJKtiItbY3O5ljdoeaaw1m885fI0/BT
Fz1u7eivA0r2uIe6yVFyMLuOPiVrvlQUiTKAPZ9cfzTF/gk1R5mo1ANkx8EdSm7K
oiMW8V+zGSuYeFya245kGCEzEXZuwe3V4lCWoTuQze3y+o/E+ybVwUACD1iU8Dok
pOyW4HMcMOPkN5DlOQduGiNuoPXNB4/Oe62M2+0VK4zW6pU+gmFfYWVyWF1+dKNU
GpgnKtJRjoy4o+VfT95xRAVLLR+m3k0+ou//J311KfrBqW68y6a3hh7k2se4pGGt
HGJj8yCR4MH1p7DabFMpG2GYMNqDvi4vV/uEG+Wwg0QIQ8rM/7lLqJvoKBDsp5WR
DWPRHcQoSeqC2jKwadhgU/8Z2+ZR+fdYI9YAQBIB1+NDHud10vgOfAb7camHS/dL
BNmKdmIBcMeQHhKeh6JxK2rRZfWfvd6GUQE+Ud2t7u6ppWCu7JAbgxhUzwzAoUxs
JkFRvzgwVRFF1u0mR1SUmbjWnn0/3TzI+FXxcIdzXRz7yNVOevYrLiCE2UF7lsfz
pAUIceaJaijYL+3lLzGRSCgiKJJRsGk5m838i2u8h8NwBXnSFojCtFhH3z7rB7+C
N+YdCnu+zb59BOZs5nWDXazL6R9S+DuGZ6x9ClSPzgcxxjh/tQEmUXfBZyM8DB6A
jFYTjqymffB45+NyULEKkUtiKpRkT+QSAN7pO7a8K0LvX53bXu8r5IBRw2lBC91d
eoxJAAFYaLLBDPpdFxqMjpU/HNX7zWW2oziJGjKJ8cijOW/YCH3xdcfnC0ojzPp7
4DlZmDRldGxtBRTDSivaRD344ihOZ1D/6m6aIGBqF3WCZ4EYOXrZNNRUq9Sn+FXT
SksnHhEx9UmYE5P0X+GYkFLzgv1ezJ1d7MnsliaQ/QN5uW+sBOiKAD2/1KH1pAG6
RwBWwROmdPm41aNsYehZ1XOcylfRxzciH3sSWjogfjmdNB6uqToelFh/hl2c/gzT
3LrVxl2FhCNiO75DV85mzX+/nlJkzrlCc47b3JKpdoJzUI/qV4FkUFDOcfUas2hr
bVj1+ZR4zgesJ9JXjbk5wjQIEwZZwC7+J9C9pmjqKYv0J59qqKun2/b3zJTpWMV4
W43t7UIEBX3kwPbeiHQOfJ1Vye7YeVrspYfyTZczUmYXKBUQj5d/osBW+UdOSX2s
KJVjzx93v45VGaA6/xjoRZXUtUayK6lqB1bFET5ZwJH6WlN/zPthlYvF9M5wxKFD
YinBMGZ9ImYxFGLcze6mTkvh9VTyAZpY3YOvZd7PIztHb82uJao3WHmzFYYvqqo/
o+adpYmQQr++Ii2uU2A2F6cutlTe9xP3wU283jvBK6FXGhNtXcjGcdQOmhEZytTF
Rc5V7lgSAYCKnrHtCzaTmrUb8ftY7CBZZ5PPPH+G4jq4fTSmcnxDjmOA/115KcZ3
Rt3nW5cxCzd8X3Uq1DowDCJWOuIfDkj6zRQPoyyAANaEMYhBwFwX0gk7Yaf4Ecoi
24w5xkWJEGeZY4MF9vvGK4HFMuSjrerLXpVQLMnvdSHtTX9Mv8MQgSRrDiUUDXnz
twsV7PkyBoDEMPrOyH79wekR9+T+08IuEknZthUGKJaICBAjNY4zHQd76SL6ef6M
tkRc0iMnwViXK3KJe27htl/dRqOzDHmklXNpKms8f7kVjz97doa/W1yo+YdTWCcr
hdNd0G0uW59+dRYyBunHjaPS7dNrzUTqanAgHiZfcacJPlA/9eJQ3JPOJZR0uxjj
ik9V5WcJIz9HVup9xSRgGtTEsQui8FDh2Ik0CDa/Y9PdkKeyYQ/eLcunhzz9Lemx
gPxr+/XXHd4E03l6VjIlWSZgQ/t6dW2u6bg11SdAphYtpkiBSex7FUEjMS3wc+7e
WUGEMeD8ZEg7LxM+h+PtF7ZxLQjDyDbxd0+sd+owmB+8xWWKC3I/SymClENCDd2g
o0cJb74OU3YBmp0lvNAoip0BKz9Go4AFmIxBNn0ZKVcaZZHmtI1hD1r5MsK13m0O
Jne8O+aU5ZdcgM8LZ3as76KASWML1uDxhp9J2EFCXNzEw8/HIq9Frd7aKGwq2NAB
kDEgWh5nxAFhIq/+5kovgZr78MZjZ0m6crvzC5fSnFi8tddf85HiTcWkNxKgTn/E
CQ2VcrvFrrgvwYRlVfGhzNJoGa3l2MlHurMnt38Rqsicppe7CFGx7V4RJ4d4Zmab
gPD7ZQ8rbBokM9tzwWmK5bqUuTnLFp5AiEuIgffF6VLpZznBri6hFFb1jZ9S3ioY
sTg3eEgOwcTwz5sJ0Uf55+6Yb5NwaKOBC0MfK6z5uBNQuYNUS6dWxeXtm2m7TlF7
iku3AJtoQqjufhPUKaF5oQcAGSkbqp/3u86ITwoUHE+mx/GjjDDdSEpYcRFRirDN
j2ch4hakqH6i+LLcWT6bEc/1YiIfWbZBtOrRvL8BIcVC2nfVnQYBukDAWGDOkFCF
QPpjlNfqQfasarTqs4pGzv6cSRsQbFPgaQTl9M/Fvl0H5GdxKYMoBA7tCxLclaV/
Xy2fQe7YT5rJzWuO0nu09hvacsbVIeO6mZLglSslFQdQcuMVMP1B+N2fvKI2Ucgw
n/M52wdgDPnjnG8IQlZ1W+AX/BVaDkvFT8bUdONcf6bdhSpP+/yTHE/qE+SCVFtP
3sO4tv+tRpaaAQoLmUJOIgOI8JRsYgGhZ6o8pc4jQp7TjbXDACWjN5NU92zuaxfK
oXJ9YBtDfPyw2oLTZwXxtlH2kz1NkX/ZiITC4KWBTfJLNjZeK/iyXUjng7/tNSzo
qGYbFdwaWvR+ldwLcsWZA+6iGwu/Ra+noboYFGz+qUk4Mc9ZJEd7ZAE3vfsQVSbs
Akik7wU2ZoKvtRmvu/sOOPaXgXh2nMnhcq82LPx1rECzhjsxCGcu54M+Q5DfAX5f
TlapjQBuaQc3y8hmZ8QoChh21VGHr5ARdcM9CyvLLJxQSzOV7HRS70X3wEYCQO2h
8auV2JZWTS1WtP0oLD4pdcldlSRPgCfbPark3fgPiygVhVwLYb/+DGc5ASU2eYtf
bYm/36fgOWZrBjwKFh0OIzqNJjvKQ/l9OF1P5kQHb58TUq7N+sMHb9d6fEpENtW2
XgsSXRUDqz129LtMKbLMh2eM/Z0iOCStf0komdb8dslF7BziH3FeYjUL704NkggO
Rg5OjDX+5gAQVx4yTQDh4fz+l5TJaR1sva9QODg6XH6AfeaeiVe4WkzO3HgHSLJe
PvuHgF6N0Ni/rHnAuqZjfWf0TQo2W6eaIa1hd2ZUQpgPVMsxRXO7LMoLCLB2qeIW
imX9CER2rscU80+dTqLY0Ae1/pTqEe06xSwxjvSVIi2D6zY3O3TzKKJxOo/mX5Mb
3R3RkCBsQh2NC//6pT4c6viLCVvtau4Va5RegyTI5JCnLM66fRpZnQudgRY408kB
alhCbP+I99hyAZ9s5Wk0yDl0dFtgdeHs1mVI/46lWs459vAJmvHKy96SIwh8GigQ
fqf+1n3CQEjLKk17lGwYCyZa2QrGYLpaYW0zZINdru9KXEyijtHK8rMLiXjWoyNZ
X9R84/tUDFLB6YDZS4eEqv8m0xwVu0ta3y5BP2WE1PD9zZbMPT8S3zF2VC9pY1Q3
rFi+mIpTrXyW4dgYKAtUtB900KOTgCPzw7+TPrUiAvflWB49vAYGpLlTCMS8U9om
dhYugLLFIlO37fNaZ69DU+UCuNgsvO5djvOC924kgx70cWw8h5qhPl5fVwP83XJi
ySwsAAwAT0ODu/7p3fwUPm0ZLgRtGBF/bp4SpCR6O86ckKigoXI6QV8KkyW54bK7
Ox7cSPICAuQNg3L/SK5gx+aQCOl7uxThRxN/449KGCOYjCheYE6nJGhpof7vqj7r
lQq1WqYgNs1PGpV1DsxYbLsAeIKx0Kv1RVUUFJbzGd5FMJ+abAup9xi4LntUtK1c
kIqfCLSNILXPbmZqBnI7p66CZpx8jv5V/mkuofQTQ8kC1VyXUIpNUI04oUMSbpXh
8cgYUmKRv/5DfzvE5AQGJyGH3cSvpi8z5w8ayOV71PcfkPH+9QWjkVHlGhw77RA6
K/vY8mhaPd04QAOLI89UZN3dr6OHhIwo8Qrx6XA8VGGuA0qFiAzyiaua/1HvtbbL
yw+2XZz7JjLfkAcuUrVFamDf55JPRkcN2rCT3ivHH85eG4rH32TI4KDw6zpksf5H
kfJ+U63hHDtrhw7A2GreBpOe3d6ZdX7FY6n6U3qyfCyi6Bh21eVN7fBu/ip7HAWf
pPENig3SZryGwQRunhbn6rmAYkVjB29TyO+p2PrxMCqX/zovCFJX3e88lEnpye5/
CbRR4/e4I2s8mGEkQghR+8QpeHr6YvULeOIzTZMGM1DPyeo6cHUL7quDbQo9mhvp
BSU5IJeXMukY6LqKsDuY8J03FUKbref2Z1aKN3Jn76/DipYpGlo6N0MVsCOuxLYR
YOsQhVergrAIgisaBcR+dAuEsmRYyO1swqlg8PPV+rWxb4+XsmtmAXfOX55KsV3Q
Hx5krm5ZZzwpVjm2k74FTEi/bYAJMymd7WhMxPPWGqRE39iyWWn9kv2SwnPgs+h0
aXYSdqXof7CPyzDuSDxABBN4NWtbxMyW8a1QuzaiOvSUm0jHOwgIAh6Vs3CpuT4D
Ok5kD4BFff3LYh6hbfJNxgfC2wdfUcA1dZtkxF5YuvX7fBiO6WjiByOZQF1eSdCP
jUB+ThZYw1ADAPdUliX3vhks4xYMpq/C/tWxcWVist+7J+Bwpsvgz/CLonwL1Nnm
BRJRZOOHcCNELNP7POGO0Ys6LK9Hu1OtRWeqGoaZis5dgOKT00jgKMRpXiMOlzQ2
nM8H/PS1uizu/Lk14yavunBR5UIQaHo+jc6TTDwWLZqd2o4TwcE7skZ6OQlhQi2M
WtIZPDSrQh7bmMjaUoNL1uKekzuOlF9Fv2qvnOVuWhJIfIQ9UtfgRlmb5ZhOhSCF
JIUT1rk00iqEEH7C52crHDcF/ERNpuHqv2vbo50QWfziQmUbSlbNurIhSjigmxWe
E3WtchrgN/BO62QwethGBxLE/6kWAApb9Kfil/zJy1yZ42+IjrqLPbjf+CeF/+0X
9UM4Vq8vLQ+gjwpdAnsvflVWs6IvLu6yVmxJHEegq/jfpE386qyWYOrxt1ehzpTB
XfO0/FD+pf2qZvN1LxzVC12MbwUDUkeRx8xA3gR/2163bVD/TFBzKal0KHr6QRFO
tuo6YIwC2vU/cMcfqfWOExoKp3rWXVkKiYHNJjT+bKNW1LyBSYdOIARsXxVN1TGH
Y3e1uux4p7GrsyE1g+YLpDixP62i1ZD1pY/w27kqmVyYUB1n3AVPOX8JBE1dusu6
X0qLhVSSypn8g4jwtR+eVQ9+MNsMchrWBz73xJ+pPwyOh+iduWG5FO+LFbO+yVYG
4UoTaeSigvd4CPfevaSMs4wkk1/29323jGBtFK2JB1YScknL1pR6XoAho9vLcnPi
PH7OY6/n0L+VUx0rZ7lKPVd7qh1lGe8wM2OQlcSSHDMQWQTXtC4VpCq8PmsXd30N
haWXrSr6v3Hk2hUaT81y6QzSiap3C92O9dngBGW4LHFz0iro3yiarompXQU2moN0
118vA8+LNn7mTeNYGqscaRNAmXyZJ/Q3bcua2Lw6pCbU7Fy8CV1GkMgKlI6zL79l
YHcckrusTaiWHbRSwjBIfIXNUvClLrhBsJ5a9m1pSmFUVQFz1ILZfjdDC+OAZ+o0
+Sol7zejOFn6gW+RalTWAForU6Rvv3pqHTwdJYFQYt25Zpqx3Ev0P6dgosM7rOmm
kZXEIrnE8CvF0ErcQzTybuyk15MnZLZvF2wwuYZIOl3D+D5rxtP+KOwi1sn8/L/A
ek5fyu6pzJJouxqlgAFm9j1tqlL98DGFPsyuabLvBAApHGHczuhZMDH3K7e16+aq
TWG8WVRJggZeVSF8RZMnI5/Yd+qZEf2+x7tNY96NOhYI5W5cfRUlO6zJm5D+Z33f
zyFxpYyshsGLhHWWqVd14+tt3OiscUe5/UC4olc08K6GZf9tW3F3W/Nya2jbifdD
+9zlfkx8buS4F3PTUgsToWaFvo9cZR4HuThop8KW4dPYIJWeeICMpL+4AhOwwFJT
ZdUC/z2DeSPSZN3jkdxaELAMSQfFp9bG3nFgazWWJUKeLG2DhZQcFg6Y5PtvLEnz
zZziuUrVUymBlC3dbdVmph71k/KlgMHG35kw2P1pMYewx5hgNAZiyV6CQubpqG5a
oYvcszwP3eXp+De1kE3B1iJuiTVx/w5eSOrAIjc+uRr/KcCPf4lu5mx3Cjg35WZX
cFwCy9pe1nzBclVjdc3Q2Gr/y7a2B1ORBzt0i2YFnbqS8md306SoQrT3Cv/5AlY/
tLumH2W2S/2JlPOeoFCEy0tIeRclrUMlpBo0V7h3dp/rOQfb9dBDG0vxvQF1Xo0E
Eq9UXZpbKfXRzpLXR+VMwkY1bwYPPm1SCWSg2Gdo6R3uhnTiH1kgCxp2YfH7HuSC
rxF4iXoN/NDD5GASXiQUXZfZPDTWWxfMU+1KqdDJ8fpOZT655VDcXtIHR6G8xKQt
nqwowpmAe5Gl7qFEySBjLQP79uwMD4W5hLPtMyi7cofTx/zAtShQbqtMJACgWox0
3At3GDYtU7vYAJb1bvVUPdBUz/VVqfwD60LRu5t+aBMXWd5ZaxaTT/jn+jg2pJw6
OwbcNrj83RbDNiaby3Mph2va/DxW8AkweYbEG7Ah8c1RMnPPNA6gxW7eZC/6Jzcm
pU0og/m30XywNV1EA4qkrfK80Ypo4E6kcEYqUctWuZQoHxJbLibys79D/wgKWbBg
gb2ofN3KEtiHg8H92h7A0cGQr1I6doVvbCWj7ZzJTyp+4KuoktNKIIslMbUPqXRi
Fgp/dNCMshj0zMGGKbIg2tVAUpPpafZuhgCjBqVTPXnMvzwYqH2K4ZjV9l+1KgPW
+wBkH1v9irbQsatjAkpy6pKZ9WMvnDK3QohXmuXChEodqYzzmPVSKHfhZyS9mig1
LkUfOWwNHXHncklgK+LUIg6RoLL3lhKhK80xUTlLs627rIyj4+Ie6PPYpt+DTzda
hr0ThzZbVFOz3mXb3sWx5ACPQFwa5aAUfUVuZb9LFz6k5YD5TL1rGjy/mp0skL2M
664vAOOrs6ryDvZqOBCvv7tiYLsuEGvbnbejmUAZzjbNZLzOCwdp+PY6hMKhgF7I
+2OY/tYiPbwk5MJfbbjm33cSAxPl0xPshlOchfPsg3IKTCp5zVwgnDf848b2hCce
emM6Hmc+dVCGxpI6gjngY4wtmJ5sn+QpmQLJjL4lBvM/NNkTtlwGR9etcN9dELxR
LnLKmWjakyUv2npnfyBV7FonXudPVtnA35f9i9Q7Jei1u3NvEQmQ2ItVXfESDTYr
d7TYt3vGTmW4IkQWcU+RQKIv2qSmp/OmWl4QgsK9TBx41ubeWNX7zSd1VVJFmaAk
AlKzRwhWlWoEKDu8GLpsjTBRt8e2Ql//NcaD6aIIhoVHw5SghRO30F2nLNBL7HeP
/14GZ4FqsyDvweNYuKiRfdEETX31bKRv4SfxGXs3Tk44zDS8MzvBGzYaTWefrNku
rwHB9VaNsuHbK8TlsvqHlTRhIDgWFbF37MZfywW9eGbjjdMem3l/0K+pBT/KC+XB
Eqnny9SE4W8nvPJyPAxy/sgKDLGy+93Spvp+8UeVd6LLBSUJtKVVtDzTs9v3cnzr
uTDV4QHocRPnEHqZL1U5dnTfTgv8RnjqHHuRL6SqtMcW86dfsQa11U2cg7UqRJHF
Iheq4/vxAnU0iigxlA9+BntskbugVrKlc6dXDt7Q4tkFCD+1RTkFPEk7DM34kF7S
FWN0R1Ogvney9HBf6LyDGVC1Z32fHW63fF/V8v721PwM5Py3gwOoftzvntG6KBPr
30S38SIvzzrdUjZUKYC103JiiRHmn+dX6h7NnaMZfP/gGNeBTcyn/wZ30/HcxjkJ
Z8qlwtahdHFaxJoctVT5GtVJvQKgSs+g2Q6NpOBI0brSLvl1MDwl87P4VZCWL8kC
uJ4FVYjaTH7kZ5kTCgQSaxGK0k/Evk91SFBU3FY/WHbzLX6ktP2Ws5ypmJ+HPiFD
MEF93psiJRW5qy/j4aU6/vMqtK7PFjhe1+xWOZhpUvdV2A23VNJf5BOEUP8ZIw8A
PWnha6kFheaOc4kU6NE0bMzWnh8zoeFTnmzowh/8kadXr3TTx/cnBELYfXBIHhVk
x6BFPmsuuhznVkKxEfi5hj16Gv7iuD7zmG1jzU3LYUbjzPPlEanxsSCUmwfJdI6o
rlO/e/WVrQhpVXNseUu5KooZn92ESy9NndWV2XrCPhx0SV58XL1nVbki8iyVWIQF
Ppca7FnwxTmQplgnCWYR63ECq7etPgBZ+AAqJr0/GVk9FYvvhx2QZ2qmzfZQ3lAl
dl/vtj/lFduO8YQJavI/1tRa3aHJo7/J1fCU+HIXRpsrTEv5daEpSU0Gz8ou3zgL
3FxruJgfn6GeCYkvvgUsxopXBzIMOufWnwvh20rfhmvEV2QYxlTqG3ExhCou543j
87XcZt5DFbedSz+GX+qTXnF+Iht10b/YOAm9FmoEWyIpV5uyilqUkfky0EBiNnKe
9xI6R5H2qcOtwmFEMd7yjhH0+GFrNGOP9ZQ5MQWmKHFsouvggqV2gJtrwKyqVB8z
SX9hC5luWklw9XE0PgR6/wAhOpyM5aJgm80B32w3OGZyqsCNDOLw76kFxJRWHDDo
bg6YiTNm/TVPqXCg8JIQTcb4AED5sDFLdkcogeCKMYW/1JCPyzMHtIbCxuzD/2/z
tWwniRVZ6UR2FEQMzDIwgO7vNHWYDH7I34yu+G6n6RVa8fcObTRu5GhGIBe7OSdV
8jQ1b0fqP2A8QwTvf36JmOX3JHXYdcCatFnWiDOyp51MydRRuX00npTZzF3FqnQc
uNnuRzD+PgPfqHhEELK63/Qm+MI5cbaW8TXmA/6gFrCH1fsFmKqNOXzWN7xz0XgZ
x4R1bDKPZjIATslqgdftDijuShvfRh6cT1X0nA6jp6dVQhcqAyjVrlQSyHJwAtR/
ja4rl1ZLqiNqLNncI5KmtPp8TTbcS31v13hPdoFu1sqBcgHfsdOBoY04d0bcmCe2
tdV/lL+twKzDGp4+Jk7hTR/8nGiDra3K0mLF6JvkK/fy/2RJr9KKJUe42KbUtJzL
uIp2J7k0jkvuMf+QPAkbe492aAMjMNNRRWeFfSJr1572vw/wrHePvQK1ZoSkptIt
7EjN3qDVHcf1td8JxP9peB/8eJfhaetLgn0/iGcE04q+ihQpRmo4NYdKFo2tvJjU
RPRgiGvsCm/ENlto3StVBfWuaTUZidNXyLFQUQGr1vaKIss6zs3fyAUzZ8IUH+P8
HPgQrx+AgyShTU4nwgA7RbeJLMcxen5QLJZqlJwkX6i/KSIqmyE/oudUAUfzdxGz
ftL8Fi4V3hSznq7+gtDwpdJsvmlJs5rV+ZJ9z0lFblCUMN+7faPqfoCHYiM50OwG
1JgAPrViu9ql7Ww586ksCisCPEZ7Troi65R2sZZoSZrYV67J80wiZYXQ15N99OgT
FUqN96RyBhQnoiJNoAGEkpMJdWK1LAlYDJ4jS1YnkQepvfYJORTbVOwki6eOmUNz
IFXMz+d161WOX9YWW3GHF67z0+c59QmI2SPsyzpzvTUAIA6R1B+GBDU8PK0aF+PR
F5P7i7GjtUyKfu0G/rAWA5BPbN2gW5wJ93bsVRcydVhJyFFYAcj9P4SOp+meLYXw
O6xxcg8OTQEDkj6AuHj7JYWQe8v8RjSdJ6Zn8uvRSSImAjRVxThAzPeJfIQWh7Kf
TOtuhEVx6Vu282qz3siFxLw+VseHi4Cm1cef9wihOwIL77PGuoAYgkXn6dE4Xw+q
5ynYjG7q59RQR/tTKjEMoLXlOQM/7EGuZiybs6XKa1c5TcrQ5Qv94SXeGcWh5ZXn
4uuCjXRwGbUBcW8OZoq1ZxN1G1yu6FB93Bq03VFGW5/vY+QGnXPZCgUpDLElD/ZJ
hVsFcV3BKGNJY1L0eAT8WkAvEOQrc4ZRlMirO3FpaQIpJJWf6+hXK1mfI31LLlcX
CofzD4DsNaNH0Gh1SSV2QGCzu7G7AexpV99V7rBz1E0IDe66407PBMGrMfYa2Oas
4uySYjEgkDd7DRumiBXpR6a9gDgdUxHNFoyPzleQsg/PQM4iq7009Rj5ssv57xiJ
aqQaV7iVoFsHPBNy3IEQ0GgsFI3pguB1qKHnbjFnJIM9QTIVDZr2bM3/sA09ZmVu
GysmHMp8TIwB95RC/6F1yo1LgUPoetcgZuj1GkCr5ulv+JqI4XMB0nrMEkH4CO0T
G4FdioeTp9F77Fzp94oaDhvd3ayZYPqx8+IZ7RTEzHiBJavqbmVViuk9x2K6A2wH
bLRI069inzFfYq7Aq1gXfn+r+l2QCdf8hBzCehbMPq5IYwq+VobJ04BxyF7PkRiP
xWuhBD5OmrUqxdtStJn29BYlb7YZkAJ35LtCCFgaHnfWOhV4B4mct3FB6axXL2GA
AV17SIC/TrcyEhpg2IrMlYz/Cs980FmgKioUAtRtSAP6cIhppZPM3LaVdphTKC+Q
JHqzybpFQBBZ1WCG/E316U5E/W3xx9i2QLUNXmgY50k20hZ/8WEX1NVquxulO5ys
8OgS32/erjq810pakiiW1HtYwdjSMizlHmpqVPOf4J0SLNWGlcXi+VO0PdgFWGhE
w3TqxOn/hGt5hiZMufFZ1nSV7YkQeHJJiyVLs78lmMi1Acu9+1Jz/yhqMSgT4yut
+N8e10iyHbo8Ux0vIOqQnO/Lz8xGktpi/0ZX057ID5Zo1/lMVZg4UvOvBgwPvms4
AmOxe43f/RCjJdudiIUhPbKwaYr81lUVGFcViIA/dYV72Kf3YnbkmsHGkOeBDAGn
zp6YhBceKblR4YonKTVCm4OAOAUegAZZHKjArmMf9vodFUB1/qXtWiIM93XuoNqw
zN0f596o29Bsjnj9cWUCajIuGN13wcmsupFSx2wy0U9DRULdLd7R12zPu8HcY47G
EG4E3HRSv+EZb5umS4KvQIjH1yuOknS7KjjkxVQ1bpXLUncfFRUGNs93VycV3Vk0
8BiN+LOIFnCDzAqPs4c+FdFIpb0XqZulezVGUNbOL3kQ2yD4DWgB6MM++tXrPE6K
83liu1/ta3k+IQULA0OhcFS+2VSqSohodUa6u3WIQs3YdF3cgzRvk7O2xEkwImZA
lcbKAAPDVu7R42+LccFlr9QloUsopV8jtKF0nNtt0E1UnftHLLjqBPrNgTL8ba4y
r+ayyEq2wbgLwOkCiubG+Q3PF5BTzd395Xiz9sKs39Holf2/vp0Id69BjWZd2jSM
qjLn5XLJ2Zp6ZyqPNsm7nKXY7t6iXTuN2XuNXE50J3NowPs8f8SDqqYWViOTRZIu
aFKOgSs6Kwf1zapj3tc+Ik6Xm6V6ztGnjk/0TEPW3zZ3hcn+iP5sZNVFT38WAenS
ae0u1Llxb8NNbIXgfEtjTRbD2zGKX3fUCAvegD0yXeoBtWtNvSYh7GYwtqDun6qa
HcAcK/OBxOu2DMpKIEkeQL2TByIS7r0eeILmQpuKpGJ+NrT7e0Ggq6K+7EcOGClM
mnuYv6D1tfi6EFHyEKA8XHRWomMpaEm2ITOFOO2xLMhoL3Qd8Q5TpbHOcBYE+jKY
0ICXW3rp8cCEnPiDmpn1ixx34rBhUlXX2Ro1IkH3smgVzWA9IJP01iqR6PfRrelt
ekBssaJ9tgZq4vIb+QWm827E3fSWpAFOP8F/Z+y6MixIU+eU6Nzp/fxSAEKk+4qH
Uggg6pAT/6KJa0Zg4Fo9AxJx4w2+TOgKK3GqGMHC7Q8sDGpcI2yWASUIB8yviNEH
oSES91LqkuEMcBjWY/qtkIuFFzIk0UctohN4E3UHTwHQSQhTGEbPk0f/j8CWKHRV
wI1ZtWSF4Ubui4Ij4QOdOhBIfHCGiTvw5u1D11OxnI63UFyyIlGCvjUDmjR3+vAe
sjdkREQuy/WiW+yLE9GGVL5rUsnfymK0/dPQIqIqfIR6j7Gnzv9AS553AM321Uf2
nhg+Dpp9/CXrlSfuDanbRsa8yNuUEH5ulT0UNg3L4Zd/JQSpss7GEc+zcYHOYdeJ
7IeSfBZwSapxSO2mICjSm0Yc4KJVgPACI17jIPhhkeEgT3Q/6G/rch6sGMIYzyyH
Eno1DigYIWRS/yaAjRwSz1O3YVrJVZmpeFgd6+Xu3BUWavNi+kPb1NA9AZwDTrzr
Y3sspsiPbnh+a+zAlLpIgDWRXocmH89F4icOQ2zKDvmfsL5Df+L+aN2PXfJUO/Hq
uRWtG9K4wAdWF0UHsILKHbrzjPhxDc/W5+IE/GHodz/utQmGfYQNHAuQrkohzreI
pmPTXCBjFo6VRv+eWR+E8aJVXE29cw7L2pMsWKjaBsdx4vzLXIOSF6nl7gtphWkl
yRyL8pYufZzkIbhMZhUwuxFt9gNWzTwbtUtzxvJLSv18BusXeKudHXGIHXyWdBhQ
jUGXenzw6RtGhdg8AU/eyyQwIE4ZEKKyKkH2wn1dTVrcrqhh0Ph8jKOSRRbT9JL6
txd0BT5SLQtk8L6guUuDAEQFQuBrS2UP0qNH5iGWTfJZ2bu0qZXlAz7vxtL2XgQQ
5Q3QEQl2ivoIkVS/1KAqa33sZ3ImlBr0wZqSXcFzUgyOT8dVKc7dufvHB8othoaA
FOW9vCUVc3aY1tWDdwt+2f4hzvpp0naZJwCrqlVOlUDYDsAt9PrLuhT4LdrnRhJU
7VGlZhywaFwqEWIvSxz5rsBc5/G+YvpTLMm2YrJF8Qa6xF2a84wsy2p9+vnT2oa2
sgYS/BskVD0c3ZvNCFObDoqrGW8kh+yMTOS5UZMx8DKJBlmTI8lGOCCq7VuluBEo
XF/EtNiYJzoEKNOqu+lmt+HqeoHiP2E8XUNq637wA/EE1gIbX0I+5p6LRHsl8Dt8
h79bVN+opSZvxwFfuoNIBMT/9ksiEu3w3C5JkClKNwY0ku2aMMwMOF4Updg6CHde
MboO35p2Tyj3g45ecYp5EpVCXSb9rGEGxDQEJgp5j9K+4EO9ZYWSN6RzieeBdtB8
WdBJM43ipiGTZdvyDW+f3reYRBW+1otP7v0HW8NSqLY0LehehttGnpRB7+84Ti60
UqePTrJoy44td6nI4p2VSpz/XvIFaJ4V9fAvEbTInUzehajrP19exQsTH1if/A/m
HDRcN/Ev37AHNDE+nIYoJn9CDilHxLNGqRLB/F5skzqjBIiLS7WB4r4ZR5DN/L4C
Uu4JU0GKCMTmbpy4702CIbBRDxngsIjzczKsffaseqLAUqdTtQDNKYkYl+yNGuUR
vlQcj/6QxZHN4ogctWmAGahMBB8WsESgl2WG76ZhCiHvpcL07EJT7w29somlVJtX
Wmy4Y7sQhflkQq5VmIkyOHTQnykcoMUO7KWvPmVB/ZTxE0T0W3AUrgiL0po9LhPe
bnOWv/utjJu9DY1BLvJ0aDvZf6+PZi6CD511DWB3UjC0K6utOZvTcflw/YTwNq8F
qqWn18X8aVRnxiHm/SMFXDRrnYS6tmozJHny9c2UM7wAZhuAfcKl8fYyY/IZzk34
5h9wkVib+qA0Gbat28VfgLZINfFgxhyemlHt7tzNGGNWybAuuPtLmpQjgrnRwSbA
d58rhkiAW7dfxZwq0iY2OvzvNEH9h2weXsehNVubSY8Do7ycsgQ867D53VdZF2QX
g+NRD4UhUqcIPBOGFVoER70aWff/mVdDqfFM4CMLzprDs5b7GR+LSdhY+Z4w9rpo
sQ77dXnJ6A9mIjm6xoveRH6+lnVkQCimYPlNXP9kAmSi9mPuADjrC6BNB6RLMN3k
PmSRUg1QHal4zMJLoDUe+FfDqlb2oIfoCZoB8ePxcDqN60+f5aLqvRiBK9CyPc/c
1lENrZWuek8WPGVvEnH7H1UzYwg4SIma9pQV0bAZSFNtrVtIxf+TK7ZJ+EGLp47n
kRwi+7QQztdinjVyLkP8oQ5ggiwGsFzmXm0+26bj5vKmlv6a8jNR4AA+78cFwiyn
/UenUdRw/PAFOpvTG9MgI39dz2Ht+9jPqXlbbLzyiQ4d9lBL8ufJdOg9PUrXEXT1
KZLT4SfctA76xjZF6JO/DT5z11i+kUqKs9CHosoKoB8pf1l+dufFzWbTz99FuGcf
USTjT9KqheJSM/drv0oVNgsPAVVaNH3KgUBno37cka/+z1VU9YR3/i+LFLPU4FmY
8ACPi+zvbhC9fGBPfUWllc6shk6CZUGWsaSzLOKA5DTm0+Qjkco5cLkqBdYp1gxt
jGNouGL7yPW2AjfAUjsTRV8DtWncJ6RcVBb4KAYgoLA6vt0Omt0/k7HRX5w9d/G/
TCUZxGx7+7RZq9ZEylX9oO7/zCBm8GRGA4Yjzun5o57IMjQltzh+/30OfLc4plPR
PMR6RRq1++R+a+hgnHJL3O5ru2PEsWP5MspLYyfgULD0bNkwxvhNJJwSWaUkey/1
LA9m2RWncfBIn/By93HbS9uiB906zFWSv4ZClda0UJRp5npFdSScLY5r74zK+z5N
ai/EvYxt6sp/zSXbtOTPEn8SprpkIJRqzXW6z46WyMNpjlzHz8itTaF4mjzZmVeK
3yaIxQuCSpszB73RXbcejvgfwC6exNA6NpV2+4+KMOr/AgturyU/X0+C47orSIW+
ieQ7CwiAHRg8dy8lSaDDMQxOCNHPI3GWA4kHQzBHO5c5f22Z0xeRG84OnKNG3QRs
`protect END_PROTECTED
