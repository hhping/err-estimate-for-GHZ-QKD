`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kPQi2r6jEtm5E/f8auI/1FY8EUnGXtsEYI6YU03NCvjKkBNr0P8w05F33Rh/NLmr
KomINmgMn0wlNruBuvc/Kh8+Cd0ZJEp4wX7WEpFtru4CRDyOW/ioeU7gJXol08j+
1j3/cOFvCYMvt5iCZXKA22M+xq5zs4ITRJVJ5TspCeGGfOczeA9hxIrYIxMS+JKU
buxEYHToRIDoXJmbTcPv4CNqC666wI6mYeeZ4gQLdMgsgBXTb8O9cc4A6OxjeMMT
xLA4sCv3yb1y2VQKcM19v+KW1NyfReceJfp30s8FRCanJ5zm+CYr2071TmQgI4PT
Q6jefDNCzKoeafqmpW3EXD/miEfLNamkAM636+7K5ijSTbkberN2ORq8G7rdiAl8
aALZ1ku15JpRB6my8/jwkpyQ4siTQLcdDgaFwUVP8tWHfm1LuMJQ1ZXM3+Okv2kD
2wa1ORsGw96ObxqK6rmShe8gXs72mkcXsOy0fqz2jOpmprjXohOO1/qVEgcEZuoI
kl9TklKyunyrbWhhZPNgu3ZZ0+Ev2grXjGFzru/dXAr0BofSnwtix5mAhdptrqsf
jmx7pHtRzGaHiaM+MCedtXQifwzDfq7Cpc70UsmPMkIRPOu/y7hCHZ7Pyn1dpYKA
PiJ0gjYUoq53SnfMhw5Scbg7qMdXvHAe4rMLFKMhz3Hxw9K0n5XcOYLG8oI1qpyi
eXpVCpFX9N+M+NNcCOuqIPI72XYFAz4vcqMyQzGyngqZfsSkAMKVedz1/nJBrqlp
DWDpeWMt6y/rsSsxNdPT6eKMXF/YQtVPu8PW3PCi32oeYUz+pkIcEZvsqqbdSoTB
wM6ZEvVk6fqIB6gsc1BkJoqrPHeIGqHNVkbHd+MuNgzaNyO0NpYV/c6tIAAhzdOo
OGaGkMxGy2ApknsFT6x8N1RhWIWjkS4Bx3Y+I2W6JvH+7ISoqGdohCHx7lmY42Qh
Ni/6446nK+v6Pa/R36P+CcYf7lf8NO/gl1JrQQOFTz6n+tFt+1gB/bpzUugFnPuh
l0rfXKW56eLRxbeFgdYcA3E73RBbxp1zaxObOdnrpk6fkkoI32IQCWeYRzDqMfdC
zJPfpBhDsv1GmzbRc+fD3E04Gwf5DPfCGXKjnOCfMwNmL1ql/CgDDOlI49bxnBtY
aQ+uLbcBvTVBmmUPwttWMW7fFqDX5PVj8xcgG6SS0hi6ApXYb8AggwIrQE41jdne
IR4cBgT7HtWktBQXmlI8+aKiPySRTIS1xem93QDhIc0HGAsrlRhniWZNZc9HbAj9
W3nC815o45gFXPJHZLrKC+UDSJWUf02zrq1Ydb02Tt0=
`protect END_PROTECTED
