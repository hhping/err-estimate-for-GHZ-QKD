`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PnkYh8RqradUuazJPXgnVVs5xmMw7C35NXoHRrQn8nme4Z2oRiL81AJgyBr5hG4A
/HQG6YhxMB+AXH/MS6z39Ik/r9i+ty3z+t1tevHbQDn90nyaFdIaeRt+CvwjMZnu
fCV0ST32urKGcO3MJNWVBBmp83DfuQxRvv4tOxyETaFkV36hY8ZRwgY3Dre3pGSB
mbBSosYoTqd1l+a0VJtc9rU/95PJcSuhZXvjhqUmdHBMm2Fzm0Laqd3GmXLdGzXs
NRaReuLkdw4vVOBU95EK8g4mZTRTOScuu4mR/EcFT3Dw9RscynsUEfAIP17MVhBc
gmEAIZxu6FCpZBNUfZuJ/WwxHTImGFtYqEEEPxCvwfx7501H08BdmF8SB2CKJlCK
YwrW3WbcSraVkcQdVljemnhW8PdyV/vQB1EwgWHsPezD6sBx51mzxErPNvF/WEdI
7a9Ci+OzZXXrmP8lBdXiYZCr93+PpqmvnE4zg+TrYS9rGFSDcxGID3I1OgPEkUv+
rdT/Diw5rZIEDBkrHE3pLnWDsgv6xyku/VW/AiUqA7c4VaD5kSyUuJ2my9LLa+Il
lzroTKDsg7itH4iUxM6grVrT/fiI42LVHRYQFLlxZsThjoYUpo3B06i1P1wT6nEq
YZI+mY8+my/vlaAA95WXwAl7guee/tlLJ5w6FFUK/V6vYca0UsR3OKOLftEQYNV1
3KC77DpZXlmPqBNKSSA1v96ll0rqhhXnZ3xL8eWVrhhOK6bm6X2hnvIQOQ8IzrV4
Py+TK0Q6mdPiul1O9NZ+0FF/G/cU+2TT9f7PBHA1DqcSNgXYhCHP8akJ7AollD3T
B0u9IpZvAa+wkcq3HS4v9NRO8x93vgFUhmaHSKw+fgMsxTaR3pFaVral90l5NQCI
U3O3rbo5BbDi0e0tf4Ujx+WA4CAuOOWagNVl8XYvJtWRnXNVbjUufnh/4RLH0a4y
XxJ9iTe1j1RRjnAIbgI2xR5IMWw+bZdooXyVPCayNi3O03m4sIdiEv23EAnoqrRJ
a+wFfhXsAl/NY6xFi7afnIeUG9tDi4idT5a38mtxP4CsH2j0X5Yy8jW7I1SbQmUU
Qbe4C0obzErlZSIxW3kzAjc7jR8wBGVl0y2v3Mxd6/uLeK4LSZj9nRpB16XIhEM9
u38jNFqY3AF43+NSJayJF0ATtDGmyUCAqQCe9jv4Cqp6UtvJxndmv/0yPGKozL0F
9qkLuMCTxl2pns7HhtgivqPKF+xJoSh8nRLuni8ssQZlnkKhsZbKNt4zqKDKUrqs
s3Jb9caQ8h/yMilkYbPPw9ygRcZy/BwEdg8zb+TuoWsNae9cs1b5Yv4lLXF05N5n
dHLKef3ciwOuAwq0mtJfXxTB6GYdjsHuXzbBg7Va9G07FBnIozM02v4+0b0+JUqx
gq9ZpaRznI5NRV1fvjoIw2LIMVoAIgA2o4XSLogkQwjSpozpm0Oh+zxy6V3KQOSS
EvPB+IYv4DngOYfuUKLOOxUsVhp43k0kRsPZBiMEbogNYkLerosP5KzorCxvjoeW
X/tk0w4IxzjH933cZxPDHiGAMlhkOePwBpY6Yb/TQ85949s9Q8QqxXFnsqqCcqza
2O525Z06ud9YMcqyqulOfiaaOU0Owg0AFmkegNKeA1I5zxq9sElK5NZXJpV97k+J
2DLjOC0K17OOv+iF0d02EBzx/Qx/wmC62gjRQzoGdCEU4fFT+Q5Xto0DBynPElJm
5Ssh+4SJDRQ5WPxl+DYAsfqgRFOak8X4+l1C61XsoKeVXAuWQvoWJg4L847uSDW6
k9hrK/BJjIEmtholLth1+xF7yO2n9LdwVmhevBpHpyRyi4ZQRGxffowVyioPZwIV
4UfT8NMDu50X9LwN2ggdQXTB0DLYYjf6+Ov+WqzHhjGvCTFxRygohv15hPqRiPYe
XZGdpgNG8cZ32yNT4mp+n8g0zclkeyajVGhXJ8NjON3vnsxV4pT03XlyQ+Jbx+pR
B9qXCvQNrPfIURFBmH7th3HR+rfK/w/SwK7tGXTYlQIkixa6BcT4eAqjgZG/gzI8
Gah+7td6GSCK6AdIswXzv7B1MPeTTnpsIyUU+JlPtvLCWSwF0heoiaUm06BWjPMB
UyYwLtW0jsOnf3sTA77f5JdW0AZA/O6Zn/Tnh7QRpfzrZ5pF6YThD+p9WLc5BcjF
he8Kh/m3GMXU2/6MVxtBaaWR9g3vwY7TawFYoMKLKxuXCNx3Au8ue92kWeOQ/daZ
/+4rVSeYP/49sOePQwlldXp3g7WhmlXVUkZOJHcJgAnYSpr48s2TJTr7dOeuiL+3
`protect END_PROTECTED
