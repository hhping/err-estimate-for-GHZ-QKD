`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9gHywlMPfxBd1x4Go0mBszwPr9o5rGRCYbzGOZ9nQthjpxArzGg1gCOQ7yFsFprC
1S92HY8ziezPdKfE7qXiEXGu1ndIgLvM7n8ZdouMl54HxsTm6vZGgU+mB1dn8IQx
/mOlP/S6swzww9B1lmgBiTSa4TD0cgEbb94vEF5ois0eH4Kdfp4q0Xs6QKRM0r3r
PLayfH3giU3rLNPmHaVHZz2xVAD80YM341L8A8lkpXjQiRuksdeX5vaYEbXgk4yn
aKor1/K8YK02uzkzgO65O87wtxt3M0KNzrTvxFKjMK2AhOL6eC08ZVjXLlcopKKU
aXIvg1RNUz58lEG6kC4hKtI74sg6ZqVETvr37qv5D3HsAsuY/TTvmXgxlPB+3/fh
hr77Ktc1rY2LGU4c6OWurggCEh44KUMANtMh57X09wphzOzYGb5Q48aEAVru/nO5
qFnRBZ5AWd89PJEn4k7oQO4uMnJ4gMIEhyURfVxQ6PgrPpsNXdcMMvsoBNJSj/II
BrX1avOajYVepl88FaNRvByaEhCovW09rJJ5p5gmIEME5JfjS/bMP2DD6+tYEoRM
rPqjIWPwV1NpHFwsNCPtOBV1sawrLX2KGzpRSN2vIURz+6Mgp6wMyBDyK0rWWAQy
Wx5oylrVN3gw15zNn9SxVQoXv8Lms0lW8/x4r/lKD30pc40cMa2qXaETCdUVDzZu
rs82P8WRJSA1BHXlBroV0tAGvZrFfsmAHRZ48eoAqVskemoSk2pjdtbHTkYhgxZs
ObjLdJ4iGyqv5sHGJx5xe2sUj6PVCKOCi3mDoDxJXW1TFFIuSlTW9gl3LmiRRpei
3z2fZnzM3uwGChPyAbqDvK7uL2mqFptSOnczzuLDsBH0rqnq7ARhYeDdxh5dD4a3
HQpPZBXsyzfoTp+L0faKFdXwWUja9VGlg1DP6XM6UmCtGuoUtKyizvgtg9IUkw16
BlJCZUm3zWxr5JRyXQnXSct3lP6UP8NUXxJkn11YEeSqhAg9XM614jnL5FCwOFeK
f5k0VpC00K/SeMYf0ezGy7CfcWeRH9DZGvOsgPPsmIFUVPzZ8VRK1M3tRUk69fuF
Mpa8MiM4rk56nYCYlTfxesgQ7/1j67BQ81WkKJUhBB3DieR56qVYuu/Gnc/g/b0B
ZxgpySvisAdWsbCfX6Y/fbPcCtq+LnFXy4tjTZAJWC3sMjPJbKj5zt1/a0Fiozv0
vG9kRg98FqfoLY7FsGE6IAUkyQrlCbXaT2dhhNWubgcJCb8KDwIooeHwpdmdmqLd
H38q/KT3uDoUWPMq28iZRyxHddJvxe4ZTwXOC2XPgZnECJ1/4kjZe/hr+Ee98m/D
dhZT2ppJk/lz7Qo7XW4TUetBHwFVtVCA+v6qCYxqficGYeVwoheKAPUcg4kH8dos
D/ClCUopVo6Wh/iBo6Ue0/Abi4ux4LMQSnbrGnWUG6XCvaqBtk43gzAMNPhyKsqF
55lcSlnoN+v4fSEvm1JpfWHj9Bpu8VZQFbVdlYPHt2RDsiUhLs9WbbJKsBA5EmOY
kXPnXpBA1UayXjYzuYJbuDsqqirlVtqwN+KwDkztdzWel/VwXMrRWdLme/YI+TGp
y4OdynPrv8QBQJhpgYE8Jcd2Ntn4PWGj/0I95dMDzhRWMZQIfFVpf/q6jDcrv3Gx
s4+k1uUnoU10qS1+E5lIkdCFaK9QA0F3L2AmRGWUyYB0qokIocsWrX2hdTbNcT+R
aqcXwkfIDbfuFUwtipbMitiaPDCzXZGvfSqAIbCnVLdidCQIxPQlbkUiGrgJbHOy
pNEMgVNL/X3j4xVpg/R/KW8A/dviOi8HqCYUZX7idWkQUwsDYX9R81pYCUct8wzM
4kIkuGqxwuM17KG/U7yyGG3b91nW1K56EaedRVqBLNQHgfI+0XxjiojSL7gtzVwt
9L/fci/0ajoQrTyw/Sfbx8QfeVnRmpSUEMiHZ+WSL9sj2re2MB7ULL22379fBBS5
jZ13vrUkRnm11Wr6A/IA3T2caDS5TkyGatgPGBu+D89Msw5D7I+Zu0zgRzaGmRFw
+59zfQu76Byw7Z+wxTr5tOVvWifjY7YT3ZbIJsh7+R+8q0nouQVcdnxiMnvSvLgT
7Jh7xBCMtlYoX9aQjHa40GFkb2CBIPa3OZxQiONmLjxgKGglAD0ot7oVhBrGYLzD
xUlX19M/IauWl8OItU//7Dpx2ip3LJFJVAZ5NOR9dagYS8pcqbVc5DUZIhCpequF
H5l9e/YfiAshBKAmr4CU6Q3fZHwGrKjm+9dTMeU3mIf5Ih9HZbXo/5FFsN11O/29
cy3RXhZnqbQAziLUSlCZryhVzozs4ySnT8VvSqMaKjdlHg0jfUKfx6t94caEkwL+
+YmNxx7uhjaZmM9N1CmU9KeT2Tv5PrNfE+5Ur0SqLR0rPZVj4cxG4qTiPnrrMnV8
Z1s2Vesgo93qnnbrguGaT6ZWV37jI+ZhGk5GO8IGAin23yTu7i5yoRA7KV/1kfla
s7NmS7dR66zK2OyKqIdvoBwMR7IGW8vu9auTCVTdXUOq/Dj1PQQofiaB/hKJL3fB
hZJqZhCCi+o0xj9Rs5dqZdoA8RIrPRd8GMJ1VcqrrovV0rmYC7puY/qDBMCXetKP
BJYV/onBFYWo1OeoJdkVoU5Pu2JEJZdrxoQtGQXPI/UhsTmwIV5NrNkoSXl9cdRo
ZTM6/BDn0/1NhVZlS3TL3Yh7goa4gklSuoOfp5h90o85Sd9/FvKRCejPkj2uULhX
yc7GQQtc3Y28qiJOBrA05X/YwdOU61NXONX/mN3pnwOo7ArTBS9kf0WVDuV/9U02
chlfndmD9R3Grd7IGwxxEHdyXpwBvGvM6IvUXEest1LUvL630go4eNKpLHBoQXvY
OiAj7A64zZ5oGUJ/znA8kJO58twa/FtSqdQnMv2QGQJYQqkKv4UOEpEOYf2nN6iH
o8rmB6IJAAVY8RX5wnBVruVkHlnH9atWDa2hkq4ftdov0dCGd0nnYAKo2AFFZg8H
apcAh4Q3ygT8q9FYahOyhejsNpBWWXbMXjhLjHcaInjtJu3tXve7KNKgNs0jprG2
1OwQBsDrTTuNQJuwWItCYGE/LZoIkRhbcl3ojJdNUOFawj7Jvu2SkXkbuBzsKngW
JFdfT8OmgLzp/tC/Od3se8UHtU9jtsrhHoPfo7v57r4xroRk+JIeqk0toqJUFr+b
215fZhYc0/pFCwAxR1tXY5qUPxx9S9H3e7rytmFeyB8WCzv0ccqfzIixjI0qVD2y
uBtzlkjfByhL+CO0geUApniMVgq/BcWFchq7++VAniuumxV4n1ONq6FMisSu/RzK
xBw9eOAmRsI0UBIrZ9hxIocU7gx+Fn1YzTRx2h8insK038wFSwiHBKrANIxvbiK/
/AozmYU+EFGlFGundDmQZy5A1U9UeLzTDg0Qub/eeKD6jIQ57/EDp+IwxawPUsZQ
ZBMRhKRtzVrCOgnwf5l39na/TMWU3eOPp/d+tdEEProgvbShblWgSflhCBYhSjqy
Uw+oV0DWHVtYsl8VJ1OyuH3lhVY3TLJ8m+newyngJKo/NTfZDeqo7e0KTJ7S2L9C
YYSxJ43dDt9jlnS3r4SXqzXunW/VC1UhvXWPtQjAkVsI7s8xJfJVk9joA2d1wPOa
ZUreYfh8iSnmcL+0gmNLPLQwni1OtnP4e74n2ByiA5elxzdZOx7yujGNGFr5YN6g
luRBCarmTR0+KImXqjSx3k1FS5X+FG6vNt4CwTQhX/BtxaWfPIMCz+/Nn4rAnk9P
Y3BooYTVo8tyiRZbefsqOKtvWe71nij7ITt0keU0u80r7Khb97k5COsbfROTTtVt
VOYvada7j+RbVAB1/LJd3gz5e1Zile81QNX7Ogb4flY3FMbG+IFjYkFBwptdDUdX
+KEigIM5wzKFHSjMPxacZeh/uHLXtRNhmHbdNRlO0SOsxditaWBV4FhjhpzqTqPj
ep60swc/mZpB6T4x6cVrqPNJB7JUhm+p8XMiAh0VF/4=
`protect END_PROTECTED
