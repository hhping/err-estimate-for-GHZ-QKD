`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SJh3QWZKh4Svu90WmzhLqvdFa2xk/cNsFbQi0hi7Sl9h6+PzV53mnE9pOfLL1toJ
VjLpwP0QmeylfjJOBpZ+H5exgXgLVNKZ4DYuKYdCZJE77rYvco0eYzj3ZS1uasxP
Lc6uO2Z7X9hizksFjmQTo6OSpwtXQbENj9l3HyY5gJ0xYVE8Dh/oazNbnkbnwr1Z
O8fg8WumxjF7pyWaiE3hmIfJmbTa+Y76Z12oo7gl/oinsKFsJCZHnY1DFYVffB+b
VMk/4zN37ak7Vualx17fi/t8wvb0SH4qZe5Co4VUeo/Ov2/LFDr8fOa9k900RBSK
z7irIXofxMVLEedDcD8DBzqVTvhNalhdi8/1m1KYA0bpB9e4MK8nAJ0DV5QiICGM
OnbCQ2yhodIaqHpSWJx+tTN00VZw5dmKjPvAJ9ZNqXGOe+1HuDCJS32oG3ke1v7/
/S+jJnGewXl9G5x1S8bypGLpKTrNJAQp9RqocQlkRQQsPyrlmQiBL3tH2QFGI8dp
4rs+eI3CLUvUDVT7rMUibVds3U1ngygIW3gZd3i9lPvfVCXM3b8emwwG5ojywdKE
qpnFmF3CrA7uy6Vg+upNv1JRs932H0XKnSLs7mbn5bpxIy9+uQVgc6EfyHsnoV+G
lYqd5GHE2waHE6PM8z3GAphEb1eBtfFwGpTltuUjGJ4J8iZI2CDeaqFDtcS+HbS2
87VDKoTh1EiKb/gXBDW6UWFeoMRxTOZD3HWebeBIVU8PW9+NCLqeKZ0cp6Us8/ZQ
lhQY4C69d/dk/cVgmram95UNXOOgzjhiDD/qzEX3jYGnZ09LR4x14vMFnuC5ZaZZ
XXFhRfxCpUd4CLlTUkcKXwEDkNEtwUibNJN22B3+C0meBcZ3PYSv6z1ninjTyyQl
mLHIErhBuGOfKP+Ru2L1SK/Yc2Rfsk/FjK8eivB6jizgabPdfU8pBXzR1Id4KfkE
SLx58u2cOdFIM2ySaoUXIm0ZUP4ZaeIVw4mz5Zua0VfCuxSTyuUZvYc+erwesTlE
Ju/ZBIxywMjF9cPysqcsj5Jn2qRMWk31J8Nbv63E+TMFMLpOqaL/uCqekW5TOhCl
rCqliHIq/ZMbjXDkOk1sestoCATuMW5p4yX2EhrqypARoui6zunDP1OHbhtOlJ5e
9L0ZiIJ2BNKEsl3IAm8lgdI+EvnqvoN05tcPNdbrfmPH2VcfzcMrO8BI9d/Jw0sb
wCXahc5aqnazOwF50amlPNr/ao4X37Qr/mXNl1Z4k6d0T2V+KursiotdjbJtz9+p
ne0iLGURv8tTosWLFmYWrDGF1dReOQSjCt6VvBlB6pZzoKrWx20edOl1Lhc6RQLn
FbOEVUQYjW9vRoOXCRdjI4/kPd7LJKulX/QrsrIBFUbMZYoJcaVK5MWci5jwUG+R
jd2pBP/a8M2aY+Rzyn69sd44wBHpAnkHjc9cVbJDNbrAdwcgkqtDQMJohRvhVux2
enZi44583T+x12bydYBISGrDz81dKBAZaCNlxxJMSUMCvhRIFr6eTFHOfadcqATD
HqNfiO7dg9QD5UcMMlf63dar/5a95YX6ohexCJl79qY8P2xgvH3Fp62CpSW/KMFC
h3Fr2MIuVcLETX4HeOTz7Im3EZL5NyPVT2kx+Nscam4LQ1eO+GAoKDOQz1HzfI1s
gBZ9POeQI3Ed2CCJoQIGb7xUi7WcUEmRVc3MDtqtUIMZnNrmLMxxfniLpgqf+ake
sYKvhgwDIKvFqNx+6GgTvtXkp/79ISR7epSOS3yKlfHueRUkIEiWkMXZqtLe/3l+
cXTG8psYDfVLBAFUg1aMjOK2oHV+Aeimv1K+6GJYP+jXFkki8EVXoJjJ8qHKkxm4
SnRLPIo/qhaf3VVx9BDL7RAp5jkGfdabSnC5bBiQWhdxEYvgFtGmstvP2/BAf3Gz
oQkmlRw/8fhLJ0fzbyq0vL1xBQ6w+Z2t4cgyQgqB9ZawLUZIE+GOSHMEIshGrzM2
K/vdn/i6KpzYRqYEEyPvEV2sk2bburCDzElwKtF8jNrsxta9BZo5oim4mGQG2G2M
xRQShjVAFh7BA+pjzDlyIA9mGLAFtiMtlh1yLS04pTY=
`protect END_PROTECTED
