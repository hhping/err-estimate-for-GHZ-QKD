`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f5MMbtvxpW5zWnrN65wtt3Jj+/wLbNKmC4HQ8zCQgd5RptdpCHFDa0xjW4VRvBYL
XBCMVtJFgNn/+nPwO9GhKfoqVOIZClxdpouf1eGDYcfm7dKmgYFImPYFs9mUxC6+
FWXa4slWrPLJllLk+tFmBgXRNfM4vkAFYQH2bjdwXsRtnQs7lO6oiZ1VwGwiRpNh
FVqh8/LDmmsfJMMXl+8567ZWavlExNqsChitJZul60iCtaAa3D5glBGir2zNb2ZB
VRWLTmH71uLKv8Wmr2cltsb18iG4TZSdhyLhQZPkMCyaSqYtF1guBWG+Y9SnXUMp
NefILEgVGSZtFenPnCZ8btlj+vSy6+bwsnbv4Qk3pXwhEn8cYLiaXipOKMVc+CDG
gQGZvVlLq51dzsB67ory8Cm+B70l+om3gZsbNb8GTFBEY6dICLMnB7F9UJLxbOoK
YFn56yYy0qiWc17rbCX7ceYtB//e/FYVN8QsTkhXw0A+wqxCeMSVlob+4uRzjB4t
Jez6Od4CKvLaIDtMCNhdVESxp7v8UnFTa5JHo76Jm2iuuxB9ruoKYZZFdK+NnuhH
QlF4IZ+5aYnQLn3zDpMpmb8gg5LWZfQNEitlf489OJE/1CSqz6XdPi16tVKsZHtL
Mid2LEMl3IffxxU1Z52SxGHq+pJpusICO+1PWjH7XQq/Sp9zNuJvYK/RJvD2t0Kq
CCZgtgvRFa0+zX3w7veoCXmPxg3pctWWzpbUCHjXSndiHO/XY90QFz+T3wxKkCTc
VrkBEq3MNFv2Avkz5ZCKB2VIMsZfo3/AW6G0/3725V/erNPO33hXKZ2JvWeYG8tv
YfWnHpBmCEsiOnM8SzcI+LRF+CEj3Kd/pkGvxqzOHvyrK1L3LTi+1OD3pQi28uiR
vk0jpwHTPIwBw2UdJavFE9NVQLqzOuyKsjrEQmcbH7NpHDPQxZVco8wwpjpnALgx
nOZO5hFnuH72qwsoIFZBI9wRbElJJwPt1Ip5Q1ugm1w=
`protect END_PROTECTED
