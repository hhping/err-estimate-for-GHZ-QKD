`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C8jlqHfemkBhhmda5actGeh5mIPZ82diO6E3kH2HR73oGKM7dxUz6fZAEmG6xjBt
V7IgawapWLOABQPOZ2pCAQg6wx16brPJkj7EUqynmXLE5WW5Gn+bdvNXyMOhISaQ
Mq6ybfy5UKuuKFgmtoei5pq//yHUXQ4bM1zocvtVm89bmYN2RHI5rWtws6Xj1zDy
XnoTFLkabtfp9ZjvIuHoNfy8vr8cINvivVYx5Px/twM5eJVaTn1NH4qBschnuNOP
4dk1scW5GRHBDjQdWwUb/AzBzclVdwaVxwbJZ+VsVtDDb0A4uHgD9WwCW+MttVBC
9HFXHVROKP6oUitJCkGntKZsW95X9n6nVO0B9wJuyJcU/+r7jVtHIEV7jsapCWFC
cert6jaZ+RZDjApvR2IT2aBIXCXASYI+F2KK89ygi8hj55I7rEEVZrC1iYQql6b2
R9evT8UZXXesNbSNR7dD+ldetFf+YZ/mXvcQL6ccq+L1pAwAU52SMwb8PBaIlIBe
ayHb4Cg9iODzEjSiJI5jKw/qBsWUeMyDPIoovG0pe1TI8amgevE3FT44EbcRtzkB
esj/D675Hc/7sRZZbgprFaHn0c/z+ZI+M4KeRWv9mNFuVJHy8CSeDZebRPFL5SWA
jluvCF5A0PiLKc51AyD0r7t4WuXZ9ZqrmNfPmtqfd711VWX+PowuuGGHDuUTGEpq
dahtdO12yxct5CJNW5oROeNj0Vh3/vyx/C6XcDsZ6YNlLOGw6wRYqseY3SNWp9Vu
Fg4Yag8i7kMFN7pOcV/ufCtUVvZX1YTRRPy5RalEQbM99kbtccxRkxckWTybScyP
jzwsy8RhsCKvu0coWJP4rHvNQ6GQNCu72xnDqk5CHHUjJQtqYVOMa6aN8oDxAwq4
bFpmATwLPjE6kZdDeCvOcYfQavPQcJUSDLIvHZvJCq+SSutIW+GQ45KY1N0xHQEw
F8DdNjAZYDZBcPjAPo3qBTRCNj8SndtVBbbloILBgMhRtyIW0tJ0P4Eyx8vQdA+S
AD82DTuWtBJQlS6ZE7giIJujMCAt17CYWmSNrqUCKtiTtpyddWHbAScgDjh/ircl
NbYacv6/Bq9jsjQa9Xy7IEeYbbK8C8HRRqLgcXotKsU7UMlLXa6dwar54UyuSQTF
RH3gKJky7Uy98o0QfHeW7xppGmkljbdjRIkDcjkvDbxx2U+R3PnrBP3zy/s34ikb
+w5H7xyPxPc60eXTVsGtDEsA5Ns9QtYRmkVm/nwFDQp+Lw5R5zytevx0DlSHoATB
tow0kLZEzOKHBdb7R3o45NM/abKZJCrH4jLSVXLqM2aMXT/fsOJt6erKrC5Qw6ZR
tHn6UvOxO2BvbHWycoGL6metiihkzewCEp8g7t1srMtsmJWLZpXVRyJhtNTJnCZ4
R0Wb6YkRTHNRY77MeyAH0GwelhmK7xmS4gI0awYzRLw6YjnwuhpNsRKxpXfMY3Py
r+4e8s57BtMroTEMb2n0RTPef0WRkjj3RjbJg5iP6o3tHsc8Pb8HMMyHdOSGQ+gq
WBg0cVia4pOAvlROs4SYLrskgjoGbfoG90LV83LpysttvV64zu6EHMXVO5tvdxaj
S7bEz+Q8iYlKWYOrT42z/uZYuk0Rgu6hUSNkAuyPjJAHVfHpTL1hpSmIx6FZ7HPq
hUd3CP58e7RTZr6v0KB+uclhylULYOqrFJ13lNub6UlmhazkYCfA49vw/YCn9wxU
tkHBF0j/fz4rykr0d9WdjvLhvexDk75G7Uy/L9l8pk3VFh7rsR/I7LpxMIY4llms
nY/ICD/qKwcN0j08MyeyuG8YbOm1DoofUjV+c1Lk1WXLYGRyA9Ka55deZmISftMJ
RWVQeWwzwJQaLvW8kocI3IVWYKS5WqbxYNbFMqh960eXsfj479CHsUWw2f7J6suG
mglALz0mfKAsACh4e0Gas1PO70DjIzPt9M+mfEsDvjNKEZltAzXmBt/j9VTw3ZZh
vdXZi3WAO+gZA9v0CJvSqYR2cA5C+iPt+pFb6p7evLZeA+dWFWhwFUJRmjfdOLZ2
N612v+8y64Yms2ZgRiwrelGWcpFB+RoaTMjliRdIXDCd5FtUWISsHn0e3KMbPtw1
zxAFHelRZOF2syF6II0oiKId/bygAChHUnHtv5borq1Q1KK/d3bMSx6rSrMv4WFK
ZqPOBV8vEJM6ZuFDhtYwlLuhoaQ86H6HV/gdANTgyCxz3zQMd0plED35UaV9Su4f
7Jm60GKr3+ioSAn8qgYOpGZQL5G2psf6xJPRuR6tIaPICncEYzRfJGaEo1vp7mFv
89HiNN9roKN8OgmnHI63W+9anYnEIbG7TJHfivUZkX2ikHlz8+BM+bwL9LhPz0YY
xOL5NkD4js8BT9QaysbtYEA5NaYKZxFMA3b0gcWjbtgUjqI5FoSgREJwYSv3tq0y
E21GMzkDx5xJufWtyvELxj8nlO0f4cT8qJjY2DpSdT9IUkG/SB6vuZlBzan7M6Ir
+NLls+qe0Ot1c7TG95NSFGdcltbGk0efgCNkIRv2xtTheabY/76CA+0V2WOYu7K3
ArLJyz9elwlHGfGOgkR88hVIG9pfZ12u+cSSlRImJDkinJmUv/dGIvIAzzYnjQD1
sf6UH9iBDrv7fgpimD6l2+FGjR6UihETVa6J4dmmGxhhR8L9jvK4VS5TYotBxlPF
7Lc/OhSUeDektJHnaUk2n2rGcGje76NkynrqQI3yIRP0VmBwsBnm0N8a/I7iACGO
FvlLvjo5qSAqSz+2xvpcM/AQdrpkXRs1oRYd/Fqj146lWW7QI6fL1QsZncLgINc4
0Zv1NcC+w7cThwX9nu2tDX9g0QbyYQs6geNZhXXgR7+6j3t9BNtcxfxyayzY8iXT
OoVHlkbA8lT/APbPYIxLtmQh2XERjXR4OYrK7oeftuah022cd6+6LL8lDhEYNXTG
sR0KF0hhW0yo+b23MXXssCxhsONFrFZ/YvOg9TfE68gWVvjSe+Seh4ntNwUVPGK3
dHIhQy6WQajRY/lfmACU6dSFAwkHxtF0H9MQoG/0Pe7mL/I1eOecXcj0yG5pdoSp
kTo9OY/xHdBC1DBFcegA7a65X/7XHww5XS8dywq6RUxJ6aqjBorztji9O8cXi9us
H8OGv2s7i+kZMnLFoOZiuL6oDqw2ENmyKqsm77XYhxrOu+otxOHN1prrthPoo/ec
hvK3kc0daCXBMiDw2fL6GXeO+sJQAHGVT27GePv+Z3zhwVh/MvSpxhmvrpE3ngOM
uO8skpqG/SBpUWtBiOlkjn25oYTDU7uKz5yLK1aHYJlwttFgNbkwbRSCNZAjizWC
6Tn0RadlLqHLR68nkaZFX2WhXWg8BerPvMBL/KH6pWuchNLkwFKpdZ7r1O4w8g3f
c7MNxNaZpch4HZUllqHNsvuxb7ryliYrojguCF3YX7Xs/Tf8MPaRbDsu/ZanowSO
QxSPLAXnkNZbvZfh3WckbStr/TNWhhCnxnq/VEGywTpakfvmJyaC8z80fyu2e4eg
Xvagq1HHGVw+uKlj7ZxZnepPLBIPA2Jzn9y8rh6Fhl7GF7gTelI6fa0O/VbtGu0u
b4cs2KuUx5x+5eRevaj7HqGoOJQSx4i1yl/AUGfON8yv1Dh61ee5IFDJm4LxM2pc
hJJyx9knKVYtfgAIqUAwyKTkYZ8F/E/FPETmW2Km7GBq0scIopR+vcsiqZxzNr7U
VH1K27Nwoef8S6EZGHdvxClQ0y9rhzmtawVX8jyBee9Yv52qxM9KTUK0vNcDcQfV
CyBxoJuMKYdOBjXA63eQQ66JOtiM8t+pnJPu542mAiQTR57sJ0Se3+HVXX+CWoa/
y2UVW37bTIxar98YlO3J8VWI6VHpeF1ske0T98T+R6WUe309DmwSteWO7TJh+/jJ
ragZoKrkRUX38EUOIhWhWqq42I/iF/Lz2nSX/9hNKCollbsFjabMOPft/c0YqgMt
oA4EujpYgZGAclMc2OjX7maEGwkP9/RPx4OA/ZSpMJFljZDVL0jFfbqvAyqMnkP1
AR2s937ljGMnpg+Si+BNh7cNGxKisqLtR3LIez2JR8uw63QI2onj0oPkHLugTlaY
Zjqv7Jti/18YEJPXcSSKb3glgwBzp/T32ceHOiJldRQ4L5cPNsRv1GFessqHW/ve
rxgNxGGoIsomD61tzIonCqvolZ9dxQbCbMXTLJ6+L/O5HCXfsNSKlKvbPrVgixXd
OfaZW3pBDg+cU8e2xRkbG/e96C31+dPUFmOIQYdO7HqJ9zNrXURKUK1o+Dt/rt42
MAfB+OZ+SSzQObhqNHHsigyWtCnrGpNiT6bCsyq2ogQlnEI6gdutpHZQN2WIRBYO
n83ls1hnRAQWfzPvnqM7+pGLVshriRH0lAEwiRQIOoTHrEq2N6SfqgFPtRfkEbu1
TH5PoB3CrXrfS1dUR7nR/crTL6HZNVuD9ccyLASMT3t2rlX8D1ZMTuCjQOiIKsoH
7pOS399gBKVyKnBKYma2hsfvHMJleys+J+mm09GWr7092UnYS2w15ZgONFdOR9sT
pPITpqPSuNt3b1kIZVWKE1j5cDTHrB2TQmuVRF+qSl3Z1uj2edmRdaVdI3YJiRwO
l/hp1cni1m0RRgL3YqleKsDsQcDmM3VxC63iBQbynktCIZxG5jUg7/8n+MI5Ocwz
Z0XzY9SWw/J1sWYLL3FSEsakEIqeJ5SEDRFNrzxMxxlHnXQHbD8W7P56UeBowiFH
dcr5tELeoHafleGJ3X0A0fllIv4FNJXf5M5sM/NKGvAX0agSfD704uHg5QU4iX3N
59Ll7tC+LAOHAyKb8F2UZFbJiLJb00QA/QCkFHy54a+YdMThu1ewrdYl9DFYY7OS
vGzYoLaYd4Vra796w6oyBSFAj/2lHKY3BiaG7AhfM4XXF7YsJ2Ey6xK5gJIulDDV
Um/dGus+/auRTJJY8PAfzRnLZ9OBxVSNHCgXf8RJm9wbWFnmz0m+D5B8ZCgzqG+N
+2boUkE6mLRoD9HSq07v3ItBpgiEOuLOID7OyGhu1ao5ZJZYpoPOHZfG0H5Y0Nkt
hjL7MU+PuKwCQYKNpk6h2FP5tmJn4SjMEA9qYCv0XyqprJd/P9DxlEnyO2P22Hz5
7lqNGfliVFJFJ4Mw6kd7yqCzoFEWRpvKA7LTw49XJDSB15WqDqF0k5EGhiM1HaI+
fVcTm/93r0EPu1dLr4JxRsOF29VJo8h7YjEau0XzT8tmTIOELdbqguuG4zl6bGcU
DyA1mw1YYjcpzAaTXbwg2WrEeAiDmIPlcoPqoQe7UaFcS1PuaC6g2LLryGLOvsQj
NDgcQ5+4jF0hSroWknlarOE2RaBTVULc+xrrvv7j4J9GMmoyI7W0NPboB7Rv3wC6
/0KuLg6TbCECDve5JHjCeTCwH+PEj10IJNlPGBJnylQCdgW9n3MRIidFVlJ0tuVH
`protect END_PROTECTED
