`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qmfyww72G+iyj+1pw1X9SeRxEbqwfDt9ZL7NuMv5TyJwOBpJF4BiwXC81pjr/b3C
NX1j60Oze4QRgYkK5PwQ2/1jEfZPp6fL5xHOBaazdg/4xK/RJeqWPlDNeBIf4WOy
fHG82RgE+RW9cCIv6bDUOdZzuUUNV1b3UBVtZdpcIZN+aE12pcug2SOFIs73/Zam
dPVa9Lc3nyg7zjS7jxH1d7ztYE4RM7tKtYieZ/oCSfA0qQR2kuIMaGml5mf5oPoL
wRiDQ8k3xMM6PGH6mwTsC8FPY7J/ZksyDxyW6dgq2RvQTwovNJ6w4pJWZ5I/fFKq
sGui/IkAjxuNWtI9CMqYBlzG3N7bBnCpgd33tXiKAhxENue2G9Aj/qWEusPB6nuU
w/BHq43U53lEjjGCYWj7JGzF12X6A3gv5GvxLgRQytWrnOBivBTMwvDBhNzxSmCT
TKVyulb3OQJ43b85q2iKVhSVgj/yt5pAzVpaeXO4lhpvC/WJdQKdvr4RwgQEbJXM
BOKkiImmKpd2dftzilekzg5rO/ezsTjE9yo2CIpc9kwJDBV4eoB7M9MAuHfYAZFa
tIHzR2c2Gy2vaDG/J7DeRtPSLbUHPsPwxRCDpAIvcTW0kQc+uQy66Cjv0S10r1PC
oEVucDhE8lg4+AyB/bm+BilLHxadD+a4u8Pf2CSgXIL5ghNY6nKiz30SsS5CxMrx
WKC/vqqnEj0BYvoGNVCK693xTvmArDB/ld51s7Fkaq1gsXF6t/uwNVlGPZRobnKi
wcuSwpwCVqaisWAtc660cUgMQzIEJRwafFsrpQXJk09OUXRryG9UL2uaXPQgo6Bs
mdFZ8vlPI4opYSo7gaKKaNxVaiHE2ruLP7Lng6TeIYfYh9mVxnFvKjegSGGFTSQw
/vQ2okGLYd2pOIuDPY1twytC+Sb0x2wkjUIRV6u0O9bxQ5wZ5Ad0+boVoEYsQjHe
hlLNDGQfhDfoCZ0+YU+7m37Upb96HG1gtTIyY0uSlYyYO6PLIUAyCKZEgtP+sTLR
oYb6G+23u0dyMm0rPp/8tdyyuzJOGDKvBYPSpLgsvIXqst0wYYamPmqMicgZCJwD
GBypouNCfwKir/C6CpHUs8AWC6ysbcJXIIbKg5gzPu6NxjfJK9lrii1shO35gxVM
cMousFy7SCqnqJaI0zEgwonidoaQE/GOnV6wMFcSkoJrXOVCD/1oWiy5Z2Q6elUN
u29vTGKd2FDuCfIU5fpPoVZItgl0NMMNhjjBV6BjnS9ixrYMJkTxgRmp2GR+ktyX
l/tuRXCuk8lwe1iiDN4wBnE39V/8GMYEYzUg2V91aBFppLXXUZlXxsamMu0QcA89
mSc4/K3H2AAqAo4xaZs0nlv4jHJMUeFf/Bt/RYhDLd4iZe5zcf764ysEXIT2LIbn
q85vzAeTOOAM268Z7KaBS4cYpjZkgskAo9lc+QciCf6zHXTNw/XTykd1joCW26Dw
G6gh+dRmAPYdZTFnycqE6imjSlkZ4EXLPTEPDq+rUWPBXs3RHRggP4FqDpoDPu1s
8kRDAVbfxjsgw2NYUgNbgNj1LkidJVdTQg4e2n0RgbDACeshbBodrUXU443MWyh2
0KDZwxrA/RoHcsrg/2DaZqDIOj7yDbRWKjei8nYNbGei7tSF7muPyL4VU+ZwfA+b
pHhe7C45ycymOEaO+6NJ3Iii5PBhMjqpDFiPOeCJHNxbeQQXgDVTCjp4XTH5L9S4
+mal4OIsy5tKEUYTCXfVAexVVI0TtKp2u1vF+ORRRbMMXHtJwLPykmuqs8PsHKZt
sNt3dADABQm9H4UWUsJpFpqnZXQp4oQLw58IA4aNktaCq84zMaQBBunFTa6v3z1r
F7yddJlhjKXYxklZlcqoc4nB0SBSqACUallqz6DG8TRcmB2WduiKxzCVu5kGM6Ym
iFns6Tlj7JnPNbRZV1mOq6vPHUq87eqPQRCycAjNrOES2coOHJ9/T5ph07ezECRa
l0DebizpIQPHJ6Pz5kL1v/PW9IW629pHQtj4IwGxBsmgiemS4AQH2iJJNVjHD+5j
Rmt9JPu5h2MxqANQlNusIFkCS96blNZw5qeJjYxYioXjhiX0rSchHUNdVR1PCAXu
PCVYuI/AUG/TNxXFPEjHChewaK02ra7j/HGk+nA8F43+yBlzKam7JSunk7KI1O5e
+VHIib10FGsNPhfkS+WMieIMPlkFwqXb4gQHZZbM8OFzlm0MRr+lhi04X9TPoEqQ
wXDE5x2DxhPii9ZQbrGGvEWvjcO8ohaT09H7sQ8zhuOn861/hN+GUGZvT94PzSMy
//w4qrdj+09GJMj+YGcoMmw5lcQnLQjTkYI8Kc9PO91ClaWsKd00gZtVpLv2m6Qd
iQJ56gON2PemQTLkvPFLCc/4JBu1/LG5MJNjdjWOVTiaNHdBepbWoRP2HyTXnGiy
VXM8kij1ORM7R4Tf2Bq8Zw03AHy/bo7gpOV3MNcX6Slyz1xl7I2Vt2Q3Tme1lEdh
qAzgdHKNG76cxUpiPAaZYt89e7lVS5frfKDPj/x9/9/AkJiMEzWe8cXZL92xXm33
qaSdrhlq4GKJ1qoUvUrx+NkDZMURxes+m3m1I4JqmKBOmvt1sGLBfu6LeObfLWWY
7LHgKN4pY30qgOEUG2dH+fN1LPlhZM6eUojezHYYNxbRNAl3KgVeN3U284woTZtu
KyRzZ8g1l1gPzSqBUyQn1S14JHJiqAMyDP+iFQQiQR3u9uWEvgwruQQHxxrZzGIK
C6RMqF31V/eMcP9dw6mOw01LqGL9/+6ldqhv+6EXavjyN6OrRS5Qul7itQ9PRQ4F
bvyP5c+pfXwRWp68M9kEjOdykxY8pan4GEPhKwL2BVDJUZ/n5y6psRSoZIm7qCsp
8hz33WmxcAQ86Eg3sYUiba8T53jXcjsdxuFcSmhVjrOOu4bERy9c5sgmiLdEg9Tx
yWnGT9r+rMg9RPqW7tiIVMTd0NkWG3p9/RHGbiqF761Ah9N434IhCyAJpsjHuwj9
arHwF2GYgvqllCfhvAxyfXiOkjSpd0cBrO8YHc2S2LoEDmiE5oWyM9xeYvcvZgvm
e8WJJnVnaK53JJYSLvaqImFQ78XZpZMQzZlFTGTG67VimhUSlDTby+mvG99/6TN/
Oe+s8Ie4RO3ZNJlYJNm+mQ==
`protect END_PROTECTED
