`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EwX9mCAJN3+gJrSkPwjenN+LlSVzaNV6G22SBwV0NBAz4+eMq51wfpu6tPnHE09A
0A/jCZyCXBBIJncUy2XFoqya2wEoGpAB3TcIPd2PGr5iNb1E70dslJiKOPEmpsMs
+qJwaw8yaeEVkUJmg4pSCNpA8BNZf08czW7E56Zv0kltnWtEzhwaKLKoT3LwUtqX
tCviDHidqGzguCR/ICH69PWS6LznstTB1kM5wATRecPcIyMrVF7ZqWFPXUxBmuYg
WDu9XEVty7gnHCmL3S+71/MdGmYQGpWQOVJK7igocIvgVytWOjowSpAvXTEue/Y6
IEJ2Xf23IhKRQng8DKn+84++m9+DLGqNydWpGb+43W/ZWwgc5XiSzP+/SKwtAexY
Nsdwj9bxq3bYYrh9ydNjSc8juIYE+NBnGRAw4IdRMl3e2A/3w0L+nZu7oS6dyhiN
l/Psr0xfd4JVyMqDXQ1MbA0K34hpJnVoG8vFgFs3Mt70tVLK4Lrop0hTjsPJnz60
tntsvNHxWS+wCJ+sGS/jrPWYhbkHAZkk1mPX8MXKvomvmxT66jrAUrfLoMQJhlKQ
EaxkWydzQ1TLswLfhdY/ac3onySI1Ui6bWfv/f36jDAjSPMLVurC6XsUM1wgqbTb
p7Jm0ptHYdJ+qpTrJ6E3ZLQxJ5VjLA/3GJ9nVWNsumzbCco/TXi5apNDBI2fRfuC
8M9i4jDc7oTP8OLRNutZidhX1MNIGVREgxihZmHgsEdfYmUfAtoCHkB5j2yrt4TQ
HPmFb99PeBUQRNhQlW6mLw0RPXTp6BakVw31QFt9bvlZLEydcqAyw4TeAQNsyFSj
2v4a1O9jUFbpaPOlsL/IRdJAXZTRhYTOTmEttDEQNmtyHB4SStoIjHYPFw8pT3t7
LQ3OfAYrRXoEJC0vyUrr1EWjD3Q0ay/LnbIJ1Ut14OIMxbBC1bsbBNjmb9tyukRc
`protect END_PROTECTED
