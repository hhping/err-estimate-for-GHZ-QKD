`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mzpUBhTsy4MJv3SFyluoyrHHkQu3udYjGPhANxb+e3FlBA3lNUQ/c4xR/+wi9DPi
WuQiPqJCtLUacLMs7qNTf/kYKF01flTMAiI8iG9n6+MMpBwYzPiLaTMv6K288y1S
XV0pfuw+3Z7hku81DXLmpPW9jJ8j/1hpLM/4s/TI2zHqJOcwIvmAw0kcJVyjla75
D+XgFxqQnt1S9oxvajZ9XqJvt6e562Xe81D5ygN24qinrnSOa9Bk3J6KadrITLgf
dM+oYbl+ZzDBCsFf0k+t7g6nzVd0v5nyvFDlkxZ75dxAMjQvRUmUp4LBY8tjXFPx
Pg8jh2iLoxBHLkNkQXzGRgZzSBGP3TIQ2oqfBSJGaCssel9OenHZMRx30d7urgoJ
DUl69PbzsWHZ3ktRrq89NQWFf7DczuqeC/kpvLaIlRUB1b67bh36dg/69i6rqLOH
wpoHu7mhaxUXmGiaXQQI+3iC1+B3WnQN3NUfShMrJUxTLxJCQzi78knAGZLFGKhw
cq5Z7jv4AXaK/eiaZc6ueDiKx5qbBywix7/eDnfJv4JZOuBmpPeO/66Mu2TJXY4p
zZq7eECFjOZv24AiunJ8tae4orIzwvCuKhT6iztSf/Y1SFXnewyM5ASomZIqjn7A
oNaBtb2+VbT1BEuKFrYvlEzXRFUPCFXAI8P8OpzUXEvKNMgnBottpzaSqoQ3idMJ
HXZUJq+NHWdXYRLWypG55DZXRYepvxAaufpuDP8eO4dumL4ZWR1NG5Y5xy15gMSA
WMZQtOi8q3Yve8KBSjavbzHurbQOG2LCkOqEeZLLxroiO9CINQ0wH1EFajnKX87s
jM1FmqQlyXg9ul0IntRDHQZBhBcEAXWGcqwzPejHKLN7H9iYsl0opNF4k3qEgvLj
YvaojApfEnIVsiHIhqPaZy0VU6p2PHnwfBO6aiFkwVo=
`protect END_PROTECTED
