`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HZ1MRwph4YJ0T/MNEoHi9yeYyIe2hk4gZwR86tl/ujTo4Sn5WXaeNzoaSdOuibxH
CqKT3hOIX8lnG9NT9DgsX+4MYOItX9xfmKOuU9lrrZaVAHFcYa4bKCNVg624u41Q
yWIn4Kva/qsWDOnvlq4WjZ6wZoxH8O8K7Dyui4EoA3ROUiaQ/s1Onn4chiMYEH6z
fAdqg+0/IL9CUvOBLncXWeTTgH+h56Pm6HlPn7ey1EsjHDRwZUYLob74aXtqoY8d
Ru5UWeTgbk++MSWxTEhHX2AL9sUPm+IvM2SphdGNvb2CI23u14NH0wW+/0QjAJ5V
/e0nFbBQwsfm36EuIH672TNR4KrWpHO1wvOUN8CM5B2e3SClRujPTafr30xv0h4m
lT6tSeZA46qMI1m09s2kcnGoTjLTHwRmB6eNAyz9OYZQ7OnzwAZMSmxFvjvuyzhy
VtBhoPy0qSfRFfMxmuar6Yan+fkPcrSCGCcYuMSzXRDjDHzPsmVpTRXRfxk+klaB
tNkp6Fa5x98rPYkJBNQs4pkGAjR9MmSWvE8WHtRHkLqk+BU+diu6ZQ7D/B3WMb0p
b36QIiIZKxtCJbof1F4hJPEaRqoDXFo21Xv5HjC3Oz6NRzwqyGZz03dBvoD1w61Z
A8mCqXZH/BqATWKUJ0TnwOm9ZB+IxNuuA4eyuwtTvlmg4VccZZDW7vf/t7T4HAMU
optNx+luUGGImZ0mSGfOn/DjSvZqhgsVN6YMWP0lu3FaurcydpKmMsHYXehhhKM4
dplxnY5uKsu/se+sTU8KFg==
`protect END_PROTECTED
