`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
15YEO3U/NxohM5+4ugPDZ4g+HpvfCOpyQ75luRXqPTFI0nxRYo6kYZTsU82z+skg
ZEaN+Tg+ioIQ1JJ2fZcOx9941vem5k2s+hXbHj0nHZII6k8R8bUW0AJzvOES9m37
lX7oyPf7AnYd8mtpXADFLvouz40KzWCWAEKYX/xrHra2LkCki/hf4OInmI9bqq06
GuC8OdcF2c6Z2C4V3xTwry0LzAk65TIAD99+0gX7tWq7p0bTxJAe2riBcVNC7Zsq
J9zotGYMwHMNMO3um7WE0o5w+b5X801BKkhPIRnemEMVWR2SUJWNMOSXMuytWGCS
+PSfvhZOI5GqyGTeW17zywsgaEC7wavL9rrThMoBrpmOJrHcNMxPd1FcdfT8kVG1
h9l+i41yXfE38LTbssO5Z1lQMokPQXCwNyWdhpPZJ72w2QDwgWfq580gcM1BU1GM
35/utqaJ83XLwoz053L9ujDaC35OuW7O2DhxwdTM82Z8TEy6Rklp2QmjInCxrkI4
o4BUeczMsJs4LWmFvG72an1SB0SU18Facc3A0YH4/WRzX8thCGH6se4MyYhNwFLs
W/ananVjl7C7R8CDcK0CstjsaBAog0N2qK8R8Y2lpGb4IsTA5xYzsN/zVxUawD9g
H+d6BAHCEisDeWI5YtVvCRySxHcx9leFsaQHqcwa4UEFRllAceck5Fzx7ks/0hp2
m/5qOU0Nrc7ULGT5wJ8xx25gIe63PBVv1Ax802DXvqZEpEAwqVwxqYJfhUcbXP8d
la88vx6dpI1unLCJouHUzuLSyPHWeF+dxWh0dZUdFAUvuFCRt7hQt9Dji2I6nTAN
NNAShF1nKBSgT7gGDcUoOvr+NsuhbR22l14ZIk/0p/ufWRnokwqc61JDKgOZcCFV
b+MLZ0Q8/Fe3rkD61px4qsEYs61zEGnY8C2mV646jp8dbgP8Z7z3f5+PERWQ8Ipd
jKmDUovZkmwB3P0bq7DrWKjhMCzIrEyUbSVJas31QSUC5fpN+Fi+1cC+o8ojf8Ha
37uChOWdbtUMVo1CE3MGVvPzAIO/1Ek2HcUbsMkt+2bRo79yepoNEJe0G42OjRaR
/awzyjMf/aPPDwwqKGpC7HzCvvP90bqn8qp6P6ZbuOORaLvUfAmI+CF7XYiMi1k0
Nvc686o/F9M0JkxKNGxWJtiPqEMpO0PMB343su8iSltKHfLfaClR8WP+2OoKzvGD
pDxDHrPOB+JOAqcLeSg+t4k1GZZimZQfSpS+PTDTG0PTzWYmqKk8fnDqX1cNuzv4
EAjxz3GzFeAsdH6fJDBSQwp9ms3TSdJ1by51S1K/5fI+YKXb46mT4Jt0CIu+YbAa
Shd68fKKroUQlf8IE6PpJK4ODemcmv+CulKUuJ3N5oGBa41JL5t9o7jN6KklDmXx
e++wvuiKg43mxnl9rU4ZAaV6JegFbMM0rZBxznLUqp7nW9HhG8SYmGt6GRx+rLN8
kHImI0elbiW5Ag+g6WmlVGEJ4bOBllvCFTDzqF8LyEQ=
`protect END_PROTECTED
