`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fc4Q5KIa/+WqscACp8E2u/XFpygyxPVTbYlrICezptx18iRmdQvVXbIayGHAMHYY
khFUBgTCY8XHWn5xRvxE/YcDBTyzBc6BxlFb+tIJHW2w+WA+EzqzSaOUBjEmpRdq
lzUCdViFE6Ft7j5F3EQ7lT/oMUSP64OkiEhLBkNASxFlk8wWzSGNdJki7k9iOvoA
BPbkf178pbhMWqVa+nhqsUD0175T1UqdYftcv2cNKLM2Qeu7xtooMfefx1Te6hCT
W2nDJsvMR/nKuEcwRZx24dAgtn/hCmZ3qheaTGufp0RGAlyfu78WdP0d7DUWltQF
kIeC042+hb8jW/8qNDXaa+ZY78uZCwzKknrTIcz0ijqlktT7GVlzhgD4e0g6BtME
LPOxW1hqIHs4rFAZ8stIPz2yFksLyfUG0uvKIqP9f//5oZmEa55XdRdYiPiGQdlB
BBWMMAL4elyEOP3WQPdUYSE3+C1QAttbDeCm6CSsgr4RyWH7mZPafXLS1qqyuOU4
Oo0dV+EHqtkLHZnOuRe23kUU6FVBL6D4fbYxcWitOD9d9+DJz3+0xPMo3LQ+l7oL
dSC0lAjo3xIhW6Llq80PCwTaeYWaysTvcLHa4Fcu5VGcUBebPuIG8WmEsLVruvKC
WJHViVDYa7TVCFz6pT4fwFbtImrLxFAGnWQfesIhqU6/17J/CpDNh9eR4fZ48UzU
9XvNpwHQMSEA9c05GPiGWLrmZ+IlpluL2IS4dSdkzKI=
`protect END_PROTECTED
