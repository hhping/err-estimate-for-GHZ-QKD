`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ud2gldI3CQxKHWUT6N0MTkfn12hkizH6NSeB0V4O51OpVjIxnpF2BknTpnzBP5mr
10QZjHISgZfcy8els6QOoh0rTwsP4iF27wkjiJLWOpCR8rxVmxbm22vfX1sTNuHI
WcIy5eVUpsS4PPZ2Db0nsyQ9SIMBGcybQJ7aaVDsgxvcwfmRIsY+UCL43OvXiuK6
cs6KGZri7XvCZ1k15isXVuKTLgaROHsJA20Eau73hUAOS3cCHQuCzDv7/JbX+2K1
SvqFIUTr303LJfH2FsuOl6fDEtQ7aczK4ntDirTfKMmP6a5V2QdBOszr81FjVitn
2MfPMXcQmqK9KREZxMUdcGgXz9MaB0A2JclvKmz2Ut1ch0DvO8pDJrbbv8weNSNW
Q0qWGl/crdCQrKklrDxEa3AhjlcHLflP9iyqJpfChLooF2BNufv84TRyVoqPR2QO
fHJaNXQSj8bvgwD88QhiEtDpA4L8q34EuJORgShAs794aP/wBzojzhRTp9HH1lEf
CZy912t5vLlM4v7XHpBuearsvxkqg/dJQzvNNzYcC8H3Tnl/bQfULzGHijZt7T3I
99CErUYjSI30cmG6hTtMm/jJbKjJGJhzpfeeY7sgYwgHlFqjyeBtmrbouXSlRkEu
sZKwwUa2MlLs38sOa509idVW1IJnhmOW5c/NHC8agsjuk6rOEjNK/f4gW5D20tEX
cFWAeny/jeG36blFd89JYagELuH3fn1XsldKR8DIE/ig6F3dAbD07W/v9ZP8HBst
6fkC7jDYZ4swqxctxoUMLBarZ+arjyyVoXsN9JbVILc8FPMbIHDlDWwv/pGA8/e/
HY/hwy12dkptJKDFpLJj3R2qazbk4c+K9NSrySolOCFylnDvquRtZaHsbOQBDsBG
b9YH5xZGku6nq0bg3V2/kLwu1ilwMFlF9txjJ92s6652Obl51j9p1+ADbMPDBZ3T
Q01NzAB4fbU/5OO50E5gsHdAqIOKrcLvqJsxbxGr+EXAXEfzOUcfdamg3cko2vu8
fXj5eVG5uM3iAALVO56UbA==
`protect END_PROTECTED
