`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6x7UyqFpx8fY3xFmqTgtA2L/XYsuYUIMGHJbzZFV8D2TUUzg9zgN1vvmVGV/4RkU
4khYaD8K0ltpq1cz1MvlPQ9Y4gPp/htDWNuO8cccAzydo+GIiUfEWS/c/g0ktR3s
FSScKxw9sMaB2sjvVF56vR6y66vPR2hKEzuhyTs84MIwvMTMiWNO2FRleo4FHdOQ
KaG4C6L54dv3lZTnKrDAdiBg0HOb7rwUnrznUGpaIJSnhL6b7v1JBL928IAnU1uD
uqZp9P83dXW4h1G7KXIqEF/mPDPs9d2kneiO8qv7gfInWR/hT4vIZu/skBc7pqmy
rQDCAYWRVtjxi2EF/yq3wtVdW4B53h4hp8pWWuBn0/EB/EB8O2o3Stau0FpOB6XK
eq9zIh8r3exEzSi4kXTw7HzM1kli1fcuishxQCpwJnH5M0KiRaTIRqFYQGQUveGd
21BSY3zlPZO46fN++RgNNVoGQDRbP/JLSxea8QtlLLbwFOYdc3N9MvwR4pui+RuM
RJUc4HPgMjpIgFPomXiObSgWo2RUfB4qpRJTKiXxd94=
`protect END_PROTECTED
