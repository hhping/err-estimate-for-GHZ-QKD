`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CmQ35uHCzQS5LvBU/Ki4rbNBNn7RE40kJAplUGHmpJ+7Kpu8+wBoOpGok91bYLzf
+qnTxjgpoWioy41M+AthDi5/POmRbpUpERMWG48FIbmRrvNh0wLJdScb4h2ByW75
0J63TucjNbsJrVQOqrZ0kzS56p2V/0Be7Ujv3+SmSdHvu9vSTv8n9O5tvz+JWrYx
ICH3n2I1yQaVXp3Jwahnd+u1RfLRaht4gD2iCLSU6X3HJ5d3wmO/IriCgKrt7W/x
IAuEeWZ90R2JHQAjxECQMpW+qjVkk49ZfhckEBWCc0ZFkkikdWDbU/7CbCkGVUiZ
3LG1sgYZSAxpuEnq/4LJ2zsHLW1gTsvb/m5dz+C6Tz3c3dFpCURDQdYzAtWHlHhc
GXxuf8mP9EaHQF+Wz/8a8r2LmTkYgbJmplosgYxn20vZ0lM3/+pVE6GMGcaeUrxd
`protect END_PROTECTED
