`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uHC5LB9vS00G2SFZEwMQYIqhH9E9kQterNejlhkxUGFEH8Ydk5/htalSpV/d9lB3
RI+uOSMU73Evvd+RBErzteQrj1rbRQB1O+CixU1fY6XTXw2S2u6bTNG6fUQOedKd
nzrG8tO8Mw+q8ETttlBC2jFM4C4vAYcDcnWn2ZzyQXMS3KEmuHnYdXp639AT81FS
hyKjdCRFfv5gDLTZwqCZ8qUGnoepfqk73zH8DlAhycvOfq1YwOrfm9QDcf9kptwC
rPtCwANbvyA8EP+gWdSCeWmCSGJWBalED0JZxkAdJYUJljt95IWyksoqFtwc7mmG
SniZvpC9D0/cAOnAIDGMGGpWLRjKtEb5RBxdI4rr/2tcEHK08UxlqMU1BoHj6YJM
m6+2i3kbWcS8KK4YwC2usOYbeM/NMQKBsjL65++JG4HLkeftSVZfnQLJrlQrJ8oN
CbD3633lCxWUsF15rfIQVW+2NC6CFOZHfv3czK24sg857Tg5FsNkI9Z7UFu3LI53
X2cKhE6hQ4NepP7mDcqq00GhrpGklYUo9SFNTUN3+IUOk5U+u6/BS4gu0inE2D7v
zH7NMawM2aTk6aT1C02YK8Hn7m6nZ7Y1dMukArrYAC2r2ddjpG9tZ/zxolD2zgM3
6UHmQP7IO4ItB2aBBrKeM4NogQDU5q4TIXjQ7tOwMLfhhq82aBdGlrX48w7hxzJO
T9+khOlUxbCAsYhtlvejba+8pNH2oIs3FsTTgGBmt4g=
`protect END_PROTECTED
