`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
93mE3Lfc7yfr6bdXEd9pOeaBrTBDsEoaqIIb4hOarnG1AxpDLRgswGQqFLdPJtXt
/L6U6MFDotRGPshcH5eEkGogYCdjG+9RDe/xVcE+xjuDuOF5tpcFHCotMSCW8e0O
AJiTIfcYm87P1P3uLBcIngGn0akZMHgQrfFLwgNiI9iZ8X5nn3CM+3PazKDXs1S7
aYQ7AEHO9M1i9lHced8TwqouN15uPRllHGgWFWdH9xcJg7bsvChs3zfRVTYwH3Ns
34PSZQI+WBm/vYgpq7k1ajke9oh3wtOUHjoRRN71Wc+aMn6FLcuFuGkBTEXxHqa9
o4JU35Yt52vTMf2IPgJ1EuU74846oyf40vC0X3WRVDpPoSqnn5d3Wqe/Trj+S//6
2sP1uC7BThxwQIZIBuiWFsOfZSrm3SuKHKGflM1671JBrnRQTvZCoZBoyIk0PbIi
pFjAFXz4hH2lO67asntutYcdXGspey0Iejyfxb8hExVmCY7vKO9Z6opt+m+Jxa/z
EFh/O5YfEToFh7zPJsOzcuhqjDaxz0JzsNTz9NerULTITRTCzYeuC/1ul6/MksMc
07EcU7HbVVoQKV+3gRbQpDtlsdzNgOXAsJLVRS93z7o1XRxUp7zhmmxZSih53hhw
B93xZBiwf+hU3Si/bWQFeKREJ8ccwr4MghtbEZLEFi9fdpnjPdp7H06PV2Iqz1A9
QbwqTtj45Bm9/sOPRGo9aFW282cs4V+d6vo27Lj+jM4=
`protect END_PROTECTED
