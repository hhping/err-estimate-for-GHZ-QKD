`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nEMYrYy5/vm1VrQU2eYLD4NXyjpoFtmh3J/Ksq17vRWj31W3xC/R3BJKbqyFxTf+
MRUwHrgan54Faxg26+Y0/HOajDxWWECeXH8BnR42PJ+nqzPDZ2zzxXdWROjgaB1L
XPomdGoBCuSYUp+qHOR0j8y+mBMtBeVD6BaGR/M3kzd4iMVt/StXjouxho2I8nrk
q5aYuNgyLd2l4up6g8MMwUYKflHnHXLHels4GZ6XauHzcHwOmwe93cOa5ENKJuWT
8rYRE7mNxOId3kHbns/fn+Win7Q+DMyOol1FUDZiWZzdO8APhWKPfmhlf73i/NZn
gQJEY5zEgqiAEwew/1AhqQes2/jeNf1jBS1qxrBvMPOhRaSFPVs8Dse8wkfW0Q5i
ic5+Do2SRa1+V0EqO4p1GwVA/HuBJ1b0XKUUVRRtRhO1JjwfbKxVngiJbB0A8PJY
tOu8F5uIhspps2Gp06PAQAclsbUoPiBKbI19QspOKQbvGDidesC4iP9YTs3AwpG0
YpzCJCsf65YJLlfZMn0txDGw2lNclXjfY3UYAwUilGI5sllYdOTg4vnySypGiyCc
n9dtzwCRQN0zbmx1xPS7XpjVtZamCHU0d4t2wRQrlqbjYPerU/3dy7zu25s0kwHm
4GMB1HQCR72FhxRY6bzjTbDaADeRwtBwOUsGlFwXBk9JqsIDl90lTWM4fGDobWTR
YSw6jDWbPH+w/iYEEoZEXLT8WlpAiLo1/MaUPF2ySUotDq7KDQItQkaGW4OtvWYj
kjo/3ZUjNG20tAocD9GcwXJw6uHaq6z0mSMWHBUQCM7qUA91FVcV7DzoN4dTvL6H
VpHIbvnW6nt0pja3pToDVcYA6Vn64sWjRwXF/DtffLiCM0sR3vUalxvatzx7DM23
kuMndUv5gJuqsTuHMVgQzbGA3PixhJaZme104iRZB/zhI4EMD1He2AYHUbomEvat
8EvU7dF4erEohHm/z+FJ9GA3I6pEwxz9Qq1yUBgaTP5kiwr2QJ1Fv80cCKv/ya0F
/yxBnpb+yu/uNlciTL1rRw==
`protect END_PROTECTED
