`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+Oa85Z/xC36vkuV2LA7GEeN1+vSBMfpLchhgBc6us46qEDSfsBEWiJ21Yh6KsAPh
0ef6yQMFl+5i+F8tGgtvReh5A5wpmfwpXdePEt4Wy8B9qj/3tfElA2mCZYYLl/yX
3RsDy2oxM9/T7UHX1QJGiCzhZS28HDqcMyPukiUoIl096znBwXo9j69JbqVpUWIN
EyBbm3AZyAQq3dIkZqruzxYU5onyx1C5Ny5h8pZ5rP3hqMuzSOTDXmCp2nwifYr/
XCf12hzrpdduW04lfdKhQ3UA1MEhlvm+eS5XKgZ4gLB2wyk5ew7+cbN85IOuHpcU
9NP1OiTxlUco3z903+Rm99HrpYYQlX1nN8x8vSdXBIQC+MwxNQVBUHQx4GUwRYtX
gg0A+FDs+mHdmY0PP22dnLUnMtHA8nh629CUKrjyzbqzcV0ajaJf7vQw768iuw+Q
CRgedVsA0wLodnMYbsNJakM/Z5AHrwxLbStSoMfjafX+CtAKaHewxk5mc0bMishQ
psZg2F27OUBPo+6qOrEFQWqPC4Jbe57whzrl1Z6A7ANBjOHxG1DQ44XISHBsrbPX
zH2wQ8xFvnWzmSuoJMAzyVf++anG98tu8QxFzjSOaRwJtW2pkU9wNNhcg103z3LV
58cE2I5vj7YhQZ1eIUpKOp0bvKvEGWBj9UhF3HoxaInZmYmFaWBijHsyAs3qbsVU
DeA0pWCSKeQKv6sHvlD0mg==
`protect END_PROTECTED
