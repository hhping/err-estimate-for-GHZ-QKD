`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TYqg8+ZNvTVlRXa8UBqFGbaF2vG3u/Zh/IC+wcgwVOY+nqJ+qbYxNdehQBUIOaEG
fgzkoARNoZSJrepTNKu9mXpiwV45FrBqw8Jn4CvKce2sXDrVQ2+qugIPC10eOIlt
XAh694wWvT2Hqbek2xfdgAHb61vMSJaiCcWAVAr8sYrQa9JZFSR1vjyXUCXKdhsH
stx1QRbk1VVY0EtD3jmgWZE57MBLqJASw98JwHS1vRdye5ML0D0mX1V6AuM6pbCf
KfhwsUj09moQYQ6KVtRFWVA85hVZcNGvptY93MhScunHVfLXHHAmU8eBCk8Nq+o9
PKM+bSf9qBhmdfmcgfWm2mYVBT8SSNfWyMhf5LXM8Ad2oNR4O5+1JUAj+QhDbK4c
hSrUo2BZY9viovZb6znWVIPk7NtM6MgYj1nwbS/mB13VY71s11KEq7S72OM1aODy
afW5/Kn/vM8IXF7s+Bo9DjafJEwKwjHq46YRGdBZxG6BncgcMxN+Q4oxAeyAsU8v
+bqLWaapYK1t4mOkz699TIBtRlkGoga+pl6DVjVN1HchEjaK1j+lbklbLLbJPk07
UxT5WzSDZkaAgT2+eilEar7IFjGNGcZWlgGxRKoj91pomwOqHvKcQp/o5ZiYqJ7y
DA9d4cSvfdSnyyOox+zqsXp0x6cRjqeWR/kMs+1EEx/cDTdNtKCAs5xnKLX2tslV
C0wf2L21yt48D5EzgG7BQ7FB/TAnt0Co8aCeBLPjrSpPHl6M2LWWIjtIzsuVA0MF
WljhIWLiIsE8yCUGEx0sVzQxsNdbuhqKojBvUOiQZsQM8c4loi5dFYyQf2gSxpiY
2OE+EnwnkNMTPdvMhzqU7GLYIMPsRw6KSLkyLl4dYceW9z4qGYt/R3GzuF2lIc4V
ObTsndWPA30383Ms4NOR2yT/YVRqtqOSXWNtnb/28IYRRrHw7Y6YzXgd95SJcsNw
H+mAbDbALxmAON/0LbJpPlo7biXz/87I604TyO6iNEKGtM6UJ2d8or9sQs8fln7f
tZ6IdWGlXqyuQsJSHEOq6oAwPowT2TNoXZlKYz0diivoxI7K+0njya/09LsvlRyB
wLob5p5VvYoP0Nq4FTXbouX7DY3+qc7Qcs9oyp0vU4FMo7Ydn7nigFo66Lp0G3kC
bLaZ9saI+i2KfCeDedVlIwxc3vqu0Ha6gbYq+YMQORYhtvO6tLF2nupurJ2P7S43
lLwmbsfAOZYJsH/ablHRJMcJmhNvM15ksQABRpjBEgY00neoHIvnTmLc6z6tlNzp
8Gih71uZXqyIlbRS8Ro9Yx4EsV8fpjHnlsxIwxlX6xnYMlN2Qgte7LWc79IK2FgC
uVSTjakjlJJPew+Cfp1o1V2wJj4ICZh+Ns41A4zLVfq0g1LMB+9c0LaLK1tiTQR0
sxOZrkwcv/BuMAURqyF74mMU6SeOLuSalAIG/u5ytIBqz8DJu/6/2RlUPE4IThuk
h+vBn3KXOUGOpGRaIxU9xDVxydoa6FTXLyqCMuBbkKJWOBaT1RWZKi9wbq3RT8Qv
p+/rAfx5+0G3UGflqDlVAktM6B/K+3ReOQJiCx8IG6Qv+84aMNNpnZFUzPO6dkuU
1JHoitP0hf/VPnvWHS33r9NSpa72HbieYdiCx+8ZVmaOx5MC4Iuh2eYSLv2Ga4Rh
bq5/cXFK4ul19vez4KG7+iXg5cowsLJuONcE3umdplWmMMyiJ99hBhlZgHUAieMN
aHgTUlhBR60LRzEPfvnntdejJGMjDrsNOZpRRe06PedqUwN06EiiTGuckLpmpfFR
VvGur9j4D1GIboHa8tSHUhmOQUHvRQJUwGazjamuk6tZ7nTEm1n44K03eAc3gHhe
j8vTGQnkEcXT8kPpvK7501q/kBTy9AKnvUiNJFnOo29y8jVfstj/HBrbWsqrFztZ
fVg1uB0//oMUr7/d/9j+iUyeQEOZUi+VKaVSjNemvwW4UFlRKW3Dh7gjzEdJXHKO
`protect END_PROTECTED
