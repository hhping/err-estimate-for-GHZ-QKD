`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FeTVJUQ+5gI+T9CRT99oCqgumve/gVNnSlLTS2kV8R2DA5bB8oPh2EqewPH38Xwk
eQjfw37NRe1Q3hLV+4tNXMDFNP8ewWTb1Ur3vGzt7gN9d8Uth/B4GPZCdiR0F5BN
WZswycQl0CgQPW8Gw0niiGNfK+x7T4hCH+mt+xVAhVXOhKxRAhcT3s2ch+DIICq1
XXkInIClQyn+Gpb8LspmH8yoOJr9NH9cfIP+xLNTWPeU6tfFZMYVOKob6TH1hZzX
JL/4+eQMwYcRmwfrHJP9bNSF8mJkLyf4es76z2JNgicHbt/XOy4bW/x/yRSlng7n
NbKiZ2uUO9NhsqJw42K2fxtWlhis3hf7ySq1a+F0aAxqhBtlT5VhmzcYSDLbtx+U
fCQ+Zup3RaddC2sbPzSToHS0NaDqrqCB9AuPmSRyyfC6gza2F0hKgiZHCzzPYApw
2KYyQxRB/DhfmR54RUsxV4YUvZwW/20Zp+YCEptimmdmuUHThY5KdjwR/9RKeu7e
mQu9ye6XL6kIkHUAj0fV8t/w2LJoeENrs9oizM6Aed6i+O9ItXFFeoK/osU91j2y
4/MANgUX5ti6EIMSvB0l1g0Fe3W7qP4CDIOFdSSi2fyfCTuLCAbPF9rwQei+D38M
H3mLgIVkbbdLjXlmAhjh0auRa6W7vMWVa6IzAXICpN9MRA3OIcw4UrrDPtuYKD/x
yQOodoC/y9SqbycqbI07IPOh2o575x3+x31gCkuANpUFoOl5b974NT6QeCHSjCfN
Il7gPVDsYDtULlZD7LqzHupgnPkdn35FojlA20ObIc2nVvLkPoFI180rxpef5sZX
/qviLPmnJEwoZmiH+M0pA7gkdhZCGZEq5MnO+yu5yRJMfCIzacq2etcR4agkIZaD
1zIxd6fnJMjP5vVCebCiaeQ3JlvHqt7j0OzNpg8fSd9PbJlvET7yjkGUfTl1wEhh
0Y/3fvdXutmEpzyDdMOVsFMOUFfKoVedU6aBl6iPYCe6E4VrN1C/PT3KJfDe8y8A
p4XUKI8LC9wrplLsnR67MniZpo+Vv4HlR4T9pldJPvBsmdyezVKyAd/ffdZbDneA
flm8X8zRKe/CElFrpHykA9no6A+lr1ozghpLbDC+Lzb0RJRIz2bkqcIh5+QIDz/3
CXxOH58cI+SahA9cqq9BsgSQr9eq5bROYKxpvJ1CkccIjA5Vc7mXt8Nh05VLK1xw
fndu85Do6GmZ2jSboufbhKotzty7RM33p65wDjFzWAwrJC/1zI6VhVkAYfrmh+61
M0TNbDTB4qgGVpz2I2Squp/w2YUZDrUkPBzLZloZxJfOzON3J/s3plwHiS16wxEO
HE/BKcukL8TUHuxlGu9d6i31gvXbPKn2Qhmnc1JQW69asdPShlkm8EgatEOC4UmQ
Jq0QucdwACMNq6jMFqh3VfBPVERhBiWWDXzNP9gZiDe8emnCNUbn2KYTv2mZdq5e
7sdT5ROwIysPdfvPrKNoPU6FFqhkc3lxKMsgbsG1l1/xMuekRs9WebT7GeXyQzZD
k2j2cduyUsztiO3QBaIOKqYUOvgTyGbJszD368EoMv2/S9t9skVMNJy6GAf1Bnxb
fMsfzfxdFXh9VngYd+poin9RXyTrmrnZd1+cYAv/fokMPLwNFEUOKG2UHzWBayMD
4vxjD2UBERW2L/I7Hr6DHiLTevFZvKHBPKd4VA3E1HjMkt9BKZz6rzLD72DIuY9r
ZsbM4I1JZgcvMc4Iok9QSYu1OWVElcJPsUOsA1mTBMl0gJ/eZpeohoccf/nebC8I
erfRkbHaA84/416eT1Ab2dmSRmt5bgGvBiAymx7sAF23My+NjZO+CIHJwE93tRwz
s847G9m2ZW73wJjgjpHqeW5UAqpmdei9I75W92+phm6FFQUtXQz5onlfKlBix5Bi
thMxDhdcicauROQ2oaHOMsata8901wTscIXAOO1YEoS5oKJK52jKXKrWV3YyBYm5
sysxTeViwsK117jsNsab1aInaKh8oNGpLS6o2lLd4fjR4SAi8rcA7BB61T+h+O68
hpBSPONJZ6/sUMolBKU5aa2gNwkw55Cu6sQluNSoE9N85FSKUcQ33zpRZL5f6LlC
Y9mg7dj6nq7b24cfBue1fz5o/FoWgHQJR/mOAKLc+MdoPg0h4r40j0PEZdpOABmW
eNlav9hI8ZRbcaMkD7+pX2h4JcihrNrtB6/ZTM9RhH3EAH5f1Jrz4EzE4iwG+7Dy
7dvj91fRPmNsL45UqJ5DgoH0/UQLo5xwexJ11A3IEn5Pc/kG859nXjfg55ZswhKo
1ObSYyuK8sFbgJqZZCa5j5Y0IIKdBYUu7OnUd7ONFF/FDvbWiXvZbEnr9oqZr+UY
zazfo9ESNAPwR1XjQpfnxe4fTtrCqKDzKH8ncaoAc1CgLJuHXgh/aTXuS9xVfPT3
ISccBghXqdIqXJHAybcD2g0/vU3m9rLtVBjezzBOW0/iyppQf76SRSOmtT82oeyS
wJi9IHej86kHfgl2ZhGfUybCWRGU7h1xbRz2U1m27rCZ8U6Gi4bT6Bv7E49qnsWZ
L2gihvmb6j4rdeXMdyn9eJeMxjUJakPXAc3ZTZ12vGqk3jBEhFTcB1dl4mmIHepc
L9Z+YB3njb6IZsPSxB+GTfookhiiJLpHFD9NDBddhZ3YrxaaYMoi22n2fwmkbgTT
FUEttK+y6j+FQy9Z2F5lq+vkH7MEOn4YLDlOrArBTadvILQFn1YJt9K+dmK33u8g
/OwwoHW54Bst1EcEfcFBwTdja1s/ZLokiFbYLCJppsHu7G6+SzlkIWaVDnva/ukv
/TAFHsodDETrnUBgJotxLq6yQS5sg5d7VvXTY+lrhNShMzF50jlJbTmAEJrFgJZA
58Mp56hjc/2yYRNOyO8xsx9p/3GpoX7rFVQ29+tXFiTvVLQ3rEi+d4C3HNH9JBaQ
vK5hYtdPnfXJEPcM/9ZBIk4NueIYce+q6oYlwMf+X5zHjOFUXskQREIEYGpCPF2H
nMyTgj/CwAPtEtMptcT88lQa0Iq17XIbfzCT5L9B6Fci3mT99bT2wkT2U21euP0H
Z7zSP5tf1RlYsVgnSaxlMRtztN+nLZq/kv7x2r+7jDg0yjBOGajSXb9/HU7hv0LP
kLee3jfrt9nML+e70yDjyyg1v/d39qiIoIgpa0G9UGHCTQMX9k9jyYNmUN/v239Q
MiCkBXq0EqQOeVLTTFR0kQ0KC4bb0c77T5QnOt1bPhKGcGS4omiHJMPTZBndZyHp
qfPo1L7iWFsZ3fl1fAscdg/5dzrhrjzTeN81RpVlUML6nD5TEp7zkAvW0GQ0ABLo
Ju3LsXxnryDBiHcIh1sDyiRJLMLz8LB/fpBSPSAWepat3VHa1nHytYHiA6mp7Dzw
L1b4aiGf/+mFNseBlErnCTjPMhzysUasm5G2l9oakEdWMPpN6r4RNRKR9h5XznFY
FwWkU14zExmMzC15mbo3W5cw7A5PsGLvdiy4NCnEQWKMb/8eMoqamKled5A/rJcr
RL+iOoQJMWtN+ObDO6q3ee8GsyEuV+qBvD8eyHVmpIr+iUqoLGG/2COlCGrgdEZy
Y6AiDwrM+KDKmHHM4zPmEs/W7zj5DnAPi/AaFZIQj04YitJvHyAZbQcgy+UB+3Be
1JahnYakIwxx0xEY0adGv964Jvh7aF79nj4ZoQ5AzaiOrdE5phIFB2djufQxkkOP
97Ehk7UD+KG0bnyDftRbT+YW1gJdZiDYN2cMIn9yD56r83K70kWAQyIE4RYDetTq
aEvfyXDic8NxeoQ3oMnMpJHsHqFVRPqR2jMhTcLYFGaqklWISUz79PLUiBuP2Lqx
TFGisS7DXw843CIokdNoTbO9xxpiDlhroADjC0dY5aTkrB4MqhK+YPIg+4oBIGAX
y6kMprcxj0UHA/rQXdq45YqhIJzItdvSgRpIAAQqUrzzD4o7gzD6uRKgNkpH0r2A
fEUckB59Ghklb24YlSW5R+74Sw15ZEtJbduFlPVDep17qA3u8uX7fpgSQM69GNWS
O1ATT8yJI360W+oyyhREjoA4+s/VV5TboK9wy+tNaUbfTJiDVQyZefLsDToEs7e6
HcVq5tOi+u4I/FML9GtcdAIBsrgnXPIlVFeIkMuvbqWYsHvs25ctp1VZH9+eyt5d
V9Y0X8zhpTssmNGEQRRdOKIs5tHtLoW7lgF3nOXSxutJM2LcB26/QXjkLkFWZT1G
ZJF2oTZTR8WAX8UdhiLjh0/1qt8P5RPQ/dnP05N9Gqmb+FKWW2fTNG7IPPh1wx2V
XPZReZnrewRfehpBHr2TwBYMzLSvYkDNK6/cg8sB4tMVLXfBbG00XgBCliB51l5m
oc2r+evdqBFGUA39f3XcZwg97ziBGwS8EpJgoRvgX43uuDdIjKuO08huayd6fxba
zbS7ckIpob1mALIEedclc9ZDMGj6W13S1roZ9PgMB4Yn192Bpy2A2CtpnpHIMDFl
CwFGXavsQhdBZ5q4lRL7qurEVHJpRklmJv0/yEMfuzf2fHJoS0g9Rj+mMwQAFsyP
92/9LdWHLI81vyskzUcjx0LM7xWduPwlRxzumiwbpAYXLQZkyIfZZg1Jxwom6jUn
UkPuaLCu/nlCQXB4m40n+9hY2gZYIMsz8nRFiNSnkDcp0tGXapr1QqMSV/GZBazY
0PicXLpvGuc5dCv9cQPFxWh0lcmpDrnSx7Isykq3czWZuZ7wRT6BJncPlyB88npQ
MWyvoZ2IKxVdzbjRDtVIZ7K5Cogkc8sDVq+Bkkt2bVEaddYD8tsB5Gis4axCnPa9
MGWdNfPB+ZIE9oa2poqRLlguqLvocbEvhx+q8sztz4ih+SqWBAYZVVcEdQ6wg+gM
RrA0VS/tn60F+4xqnKyY4yUuWJvd4PKHBq9Q5B+E703gWeznMmxRipZlHhqM150o
CsoIntxS7Z2H0HbiEMJTbuNSH4mJ/DVjfEsuMQl6RWLsyoc05JqD6XuG8AEWbYvt
TkozhulckAPrs4RByMgylRqxxNnySi344u9MoCKKUjeJNZq02N1A3vS8gwDicbIe
9HL5smbaaynVAQGFEb7PYwlcEp+phhSdEmV5py4JR5C4IkKqtXB3iWnBD6K3Ifpq
M4NKp80PS8/WK66psPKxnwrYWAAiKIUtZklCVh59Qw711PvnGmuXxyEF4aOKUOlk
7QXgxXPlGdRkUqxaMUtoXIVhP23yscEcdSiQ1ccl5rro+DvhmhYW/ULeAg3go0rH
7ltz2IKoTf7c0UVDY85TM+zUv24XQ/LwgWNswWcb4cS7tfRibfpKepgr4brNSgye
ix9WQkvBG5U6nP8NVAzfY+KssyVKJhkap1/el1F62d4r6DcNGNWz4cxXVZBxYAvk
oVUWqHAAi4z9teHAEFOoDwvwEZDHdwov1JMG5zMyTmGjdpSz7K9XL0m/fwoZLeiP
wfgIg7PaUlpuUO3UvK2WRv11Wt/xrlfclMDQo3uBrItoALJF2ZY8SAX06IBhEhy9
hIGkvgH1w839zQkPhTh+/7Fn43+HOXQyDHySh7RrcQps2n7EADL75+J/S5+6uyRR
uqk5Ws93UWpY4B5Gz3T3qKiu/WZja+42UYwToqPCXCejgA7Gi8BwKFRHzhvAAxrm
G3mMa025Hkbx1CyViSXNLQ3XL1XZT/GTskvDASt254kOyZm8GUj4Fs4ku4jDWxgj
VumDeX9vWsfAt0kTDMOV1Hvt1moDK0+OK5T/Xtp8s7JD/GFJUPBEYPukL2Y6xbaG
toG6gbjVwFDxMvPQo4v3y5EUNhlbqBZtXAArtQoVM//VykdVdpVZPR2NVqwkFeiV
KVrSQgMq0+EqYKV6fNUw9P1q6/bIyhDRyug9ZzpLtKpH0qVFxEy6AeNwFiJGj4XV
t4SxbQ6sTMDbf3jyrdFo96sPgRXLFapMcC4AfEAwXrVyrET1XOpy1WP5wNJ6VEWB
wufeby+1Jj5+zSCAxg/x+O5U1jhybOnOOfqyE9uez0HiQXueSNY8hdd4RQ/bRjet
1HczroTOHmLgxK53KSlNdtggtrwSsZxzTkKnurnhzHZnS0kMEmVtiNiLWxYBiXdB
rUisveS2gt0HAAxQef38NSIhp/l1y4rQYxbtLjgw5FW50QGmT9iiisUq6MZoYaR0
4mNLWz/Gro44fXFBNoTNv3omZWMWVEMIQjkHFUMiv09QKmTWpxGhmwZSdcB/NGP7
258zU2sGnB5J7S30MGsxMr4be/wUE1fkXulO93NldN8MSqj5smOxtICFNy84NNqE
8L32ynKr3XqvF4GM4ygSGalxqAhzP5nCH8t0EqUBh6RYm/QeXQhp2NP1/tNdkYWH
xc9QO/mFSiSM4/1BpXyynWPlyD03dF3vCU08vPQbW7yur5rPSYVgtyH871F3q8a0
in50W5o+ad2XTAuzbNquBKa3DNp3964OnrPxT+d7Oz3k+d7Wc1oQrTcyEITPF+ju
65RVjyktpKUYD7k0NBXfseKvajFdlOzT3ujk2rZfIZXy57owLOAaxq4XUNPwH+Hd
PLa1eZwLYtCrEvLdERcX0RN/1LbkQSgyXUxyTXLZij3vTz2OwFxSPFxcWjE1awCH
U34zjCgCQ2SyvfAMqICwixc2QVWopI31vfbRJAVnFcr0rMcFdL/rLmpRTnYGTEGw
ohRztqVhYSNkvKiD7z655cG/l/goNprWH0ECdhcMxeoph4z78KRTDyBYxjtGDYZ5
fWfCfD7Y8dD88EAhg1jbQyHaoUT8kqeqi1OuQyyOcRnjQUt1bijZhRmxmWwmpsUr
uouytu19PnCFPalJKfijNsVBXuLMcRCYPCl0k4wQMeH7lxLp1rbpqFxxK8B7MFs/
dlSa4ShOpMfM2KDkAKIqYtalmBCtx2mY+df4w6eXjs02fdJDf1hQ5uSBKKBWI0em
jPgzv3psjJDJSN2WscdLJVfdfoO9dPlOTWMaqVMSObn5En5QVKrSSQoVnxLuogPy
CjENthZKfA+Z8keDJ5/PHBoWxeuO8BWHeoGpzJVrZb0+YHmQoDi+jyDGhz5+8oN2
4yzidoPyEZXcPZ1rKKcVrusMElAtF+zXo/R63Yh/VYlmNKAW7U8+zLQrdQ4aUfZj
BTGb26gsou48dOfIl3wam1RDxzISjRGdz5WzH4QijtMxzPwHtvkTJEVTGRngW6Kz
KdymSdcUkOvYGB/fhgx9VlctLxF0P205K3dlnDZUe5GAcEslfeHDNbsgl5vTjWlt
moL/gE8eKW+oBKr7OlobU9oYBWiHouz+twe8UmEPvyFToNC8T/SoOxzO6+kchY1z
rX/E44+AiMOzALwu8z14m+JMLGxiCoUlJUdfQSKC2Yxtvr8GAfPWYfZa2p48N8/A
DmYjnuBJSoBY5pOCOsesEgls3T4f+6FXT78Kpy7dVx0n1xFJQiEWQvzZ5rEG/bMz
6nIIuTJb8cCpO4gqK+jAhhxujoYoT9AJbjRJwKawbod57Rwb69r3eYKWa9HiU6HF
ur6y41RHX3VWt5c6S4yPoV6ChWg8apiF1AFfqsRNLp1wgBgvkA/xDP5+e/77mxhO
dNvNSKOylFmyexgQWRiC85OXTuxVGynAImGiPNSdJXADjo84SSj7DJNi9PuApIIp
R1QSn98cVlmc3F+4FLsVkxu61spgRwrrh6bVNG5D+z5cLbQTJXbPbEBi3ifZ8pdV
LeGZkLp/zk+n97hhAzH4hT9JcQvTNuqDQUjoRpR5ybvh+/AoC4E5/zB9LIfIoLBu
DY9tYMimANErXSEO1yMkG2xM+aMYWK8dqrQyv2Y+jeqsvJ+lu9eQ21lc5IxcVrra
V2pJ8+Id9f1DkfrpeSRmG+PYQ/vO0IZQzNrxoAzRhO24i2xRglHykFmAOkcTqEn2
zpU31eKkaNG74QMUqDfAbsD2IIUXdUosFW9GprL+cEm9Nbuyg/HoVbgaU+TEPW1L
83pOswJpDBOoXyoAtIsARqYBboTdHV1l2D9hfC8n5L0TtKO/OSF629ouX4+foosd
oiQfne+EMbINbqflIanGGxHHaAwFvmDlHXimktsqhQ/J80iJ/+mdGLzSeDmM3qt4
tUe2Awz9pC79NkvU8GU+mq2l5ywQun7Gpe7YmKgZa0nwSzek0UyFRloamW8C40VH
rU2yMmvuSrdjQwLUz0UP4Gzr4UbWy0Qvet+vWp7IZaoyEKym7WB5nQSPmV+LvnfA
xqJy7yy+Qr3s2aHj1ecqGGLX3OE/45SXX0avCK8UlgXARQ9nqnuJGh5a0JARClo/
2T31l61g7tNxKkWN0YDfS/eLjqWHoLlU/S1zIvyW0Cuks9RpES3qna31znqkO+QA
CGXSm/+bF4YvONMqlJRbNzxZIvsBUA7WI7bqFSiUwWo1KFiS+8nsB9gyHLQoVb0w
Qr//69MhxZJx/PQQKEsI6Gc5sGiReMUTaYCS13eX4Z/MBKcugpfkaBtbORCeN0Sm
jIR50cxctUQLbcyAqHbpHwSyDPqOVCGYqj6y5GqoJld/5uu4dMwS852+5Nx4utXk
LuedxeTac9qsJ2f6A1YepH9yl0Hz0iuhD+nA9lpC2Ic7FIYaaMcwLXaZKCI4m+fx
AfsEJZmNN6fnHjb3XRTh/6JU2SLId2xvJIC+CjctatGLUQuuKOEFT+kFGqIXmgvo
CqTxVAdn6sZYczE0M1ZVtdoSjP8i8Cud0EmfB7NLlwJ/rhJ35s2GWUuhBv3neIBO
TqTz5M5/tNcF5wacuSykZ58Q3fi2rTdcNcQpyXbTHQMDpxMCMzzLED1+3DGXL6ZK
vgmwIQDCWAjUFfm3+03u9LTKrUhXGZNBnfzGskY+udC7INzs9BGKbzkgslDuY26m
4TP77h+mGwmXWwvShL0sjTJ9i0lMcuja9lxem15P01Zl7dIud9JppIQ8D/9sHOIj
yjINMxBW+HoWEIkVgpgsXm7O/RxquAVIt2OIL0GAP/Z2pwsN9KhgXwGU57r0RaI0
gBB0a5GjnK4AyOPFdoTcUj8/FYSIga5qBE8U3rlCcyh/l46AvNAN3Q5nUudoMsCS
D6RPJjONQh1TlwTZzbKUv8clYeKtg32Z7l/acE2diy+nfN3cFnul5GGFsa73jAwZ
36/K78ZIX+4SdciH87XDV4Jc5OznzxQGCu6K9JuxAyOFLMypKM+RBWgw2N4DRPBu
2sUFYqxuv2PNfXoXLVpfMlckNNsJdXHWOnrG0vrDVqAj22asLGCEaLvTcZ56sY/d
jXdUjljrrWsu1Z/wGJbv+7mLX1XrWC9kLmwOPd+CcR250wrQAYroxHjGS4VIHboc
rch/FI33TF7nqzh1soslf4b9V7BhuLvlLkUWKrBBuAurZm28Td+61B6vKYmm4prv
bj9VaWhhlwQPnjI1m+EJKHg72U3zX4a7sDQsLuobTVq5joCPcg1AezceVTdofRyE
6VazvU8PvNy/ig0cCy342jCEmlx4yFN4XExRYZkY+wKLxiCX5KSSEhOcr9S+nEgV
mkjs2g7qbcVozVF0nOj4jkRu0w1dwRja1LsACVIsT48AoJf8ztSH+t3kGxxlzD8s
b96p6lPEjX8yPv2fAa8RdvSF3eQqfR2eFhYmcjPiC07umIisCryBLPzvGOubuvr9
XSpL6+t2oWylz9a5JiMB6iIoWeM3X5os50KQ0F+oRLCoGXCbuu5Fks7sY5sKil2V
IZFPEUlq3WyovRZkXVsIolR8vXEL4N4P8veyG2Dywhj7t1uzDy+oHmeQRsLK27h5
7hnvrgrbXmtdX1KGM3EcJl/6dGy5XZJXSknDIxwxPLYi52uIjAvhrrZkajqhU/W3
X0DZhcVJrcDIb+trExQvVQOHx0kJMEqR5YyQ8YGDyGVpYcm4lKXW6huNmeotScNA
5oQ1zBwOU+Swur846KvvouSNFbQsQ2y7UlzXFY2Pcm740G0qCAarnrNMwenO9Nau
NwM6lKXaeFyUg2KQi8IFwzUdhV5/EPyxeSoRX6kiOgJFlwJQUcNFKKeXqL2gv//H
z0JQbhJaJfHftEgxkf0nnFk0jW6gmLfm6vJxneQGFP1v4wVHFgOD/sIsNBrBs42z
R964Os2teCPOV+8jDgUQiYvf1+ZQIqgp9KV4R8LSvtFiSg0GokTh0o+3dOVVlimp
/oDEMMQLm7FvWzQmLtRyOJhtRmwoxTyYf2Cn9tigWTtuzwIjNulPO3fIFdAzkSxu
7fN7LM7zeadAlTmhTyA0Mjyw2Aqvo61v5ikY6stOoazAXookuJ3B037UPKWxirE1
zcrxTqoQp4RinZ3KuB0CUP+Ipxgwl00Rj8aYyMoWhdYZSUo6TWN2zr85GV+rWKCa
BY8NXIZKgFdKi6O91PDoN6kKhyRhraDjy3aX+CPiJPxoTxNI2UMzGljSlOIQqBBP
VngpnbU9RDrmMUFem5NjgtqKyBnTv+4mZ5B0NlpuySXe/x2QyD84pVpxz1REku8O
K4e2AZ4QuzxcYh2OKpd+5G1RdtY6xR2gHV/wqzDev0Qdv5orV3YLE/7pT9b6MkaJ
uT17YEZ1cMpNjz/zBYpVQQCbq3aDUuVpIb7C9OJayQGc96Nb5xygeieBFYKY5yVk
IkmdUpwy+Htq3Nd0Pj3LaXCTKQxV8078OxNLDgmPb+ldbQAM0Ezikbc2F4ANK+qP
kSAZ6yQrx2l9gAfIidirdb/Kofe9fGnBphguEusTSVKeNEd2H6dFiyGAKAVEZr17
b0odJEcQOuv3YJ120i/NxhjXm2c/BxC/OaeZrqYcebwwApyiEENvEvUxFd312AhJ
YQbYJc1QD+mH1ij2wtqXQLq692OFtrQbyv8C3iY777KS5s7Fltl/Nrb93wuwFeZ6
5UUKX7BVxZg8nrqMwTqZTEmBsV48pnspUUK923XjdCnKtGt03EJ49EKd5lQisWgy
8fbBbCxMngYozEho7bq3DLNz/1PQpSlCK7BbYcNzA1nqEPJj3hylEtizT49/yyQo
rNvTJoC0zxfGmbvxoLFFrYOIEFOwvfEropBUJ9cgcPdKuqpe9H/OzFTLbkpROh7u
DJDlxrhjP4qUgDjVOUNLKfOZ8o0OZG8uGUwdF1Qb6G1GCovk/gzCHb2An2CQyyEg
D4anXnovjBaLXLJ3zYhHwSEPcycI2Pyerx4pId0t8MxH85Ym0tCsWTHkYX15aRrC
PyZuZZtlHKMG/Sopx92mlyTKz7cgSOcDeiNFtrubEODtq0eVQkP7QneOM9saFh9D
1eFBA59LD0Khbe1EYKhCIEzsOdxvfyC80tOIIYaBbEl7Q2i8P9X8nNksZhpN23Wp
RKLNg0u2zkOzWEKSVGR+/lyN87rQwRTqIFz8FHVgD9nvETloYS+HGDNQ+d5l1eac
VNE1HeYytmqQEQO7agvILGPsXD5Mw/05iqvS7oCEKnzmEmee1lpSlr2z4FtOVOlM
m2o6iExuSSDPEGjgPixp2TBMRh3OepawhxyNqkR1V+mgTBc2OZXlMBE1E+EnIBTx
j+qvAB1qQXhfk8weiQUCq2ql61AZnkD3jaeCdPlYd14t9/vaOzo7hzMalI6Tlz1E
g+JSp984csANN1GoqroWvVZ4zjP8WjKle31BO3vm1BH/ou+M2nT8a/FA8xEBJ6g6
frctPK6BX1hCFkTgcDoJ46uWXxcZATXWC1eFvy+IEM5Blj9BwC2IAxv6TQ+24pFL
uNDjKplS5naGXCpiKwotGrSsXIzBPs4L2H/P8lZfa7nvZbcgxqPK9D9SZviDG73F
MX8GclUlUPheP88ZdtTKJoanrpqGFzP6IIGPIRZVh0LFeTK0TYT+2oaI+C1GoCBA
o7bcEpVdNgbE7C4fNqA/BJq6tkQWDSiLxo0oDpWOYJcJ/yin5BsrpGBAR2fREr3l
al0uOIkCj2RjWAKSWQTM0yDVDgux65oAFbBwzsKT6U0OhrUKsDf9sJ0/9GaAqfAx
aShHHqDbgkNNE9DXXeTOfRHMu4Xvd/TfnMgcWLe0392w4AQME2HE58QP80m8u9la
KCB1+g4mPWOBZb2Z0CPvfKfPtWSpXA+6UfMF5d3QVkUXeZ4kJUN8GfNUC1zMWFka
gO8mkbIaDQhCT9RQHbhckPWCObRAV1y+oQc19KJw/d+jpMQcghZoSuzt+BERAoXP
2QGFK/STJR2xtdG1cp1m2n+/NtFZJy0UlvEmMD42jy8y+K0dBoZt6dzanUzITw3O
A4mkT5w2v2xFYCEVK//Ep70k+VX4Ul55pv9StPkyk/fuAb0GgnjJPCceg4IehBSZ
ED7GONL/nF/bW6UIT/0HbhRX5eYv1xdymKKbbu3jbAHPu4p2iLOKraxXDQFdNe/X
dUbYZp+hCvMABl1t9NZ0I0AkWBEUeG3o6MOTU1me1i71SrwKkHzpWVavUNKmsvbr
anWIruzNxNFPofkmuTZbedGBwNlzQketd8EpdKUA9Upc6bfBTbbq7DMso0ysGBlw
vXwssi0EmUiVtV7QeKoDXSPbiThOtRbuRPSOJcaNwRPAV8e3CtP4MrHkLBu/Vts8
lpZv3uQ8bm0Fm+ciIt4rfiT8jdByI2MZBAPW8CriLM8eE/Ql3x2zJVk0zQLz2BCm
66EIq+AGRkt/nZ5avoGOk1GCc1gZbGNN6pl7BiFIFN0vTR+sQHhO6L/NmeMO7RQc
pnyAjjAkMNZVKvIN/HIbBS2+1huJuvjqdmcOS8G6bIQqmggOJiTxb5KW52nW8ILe
Cczu8go/DCcL+FM3H7BkudHN0v/zB5UWOma7z4tWOIuF4VBP+I0n/PB3pMm1iLwO
nqZM05GiXGvsA8vtJ66wx4J9SN1yQXvz4NC2YQXxxcKFCyJrRsyIhxoSZ7z+vEno
5NNQdUHBuW4KABsCJy7PwrChstbE6sZhN7f8tmypc6srcz+f4665OBFhcpxqNskZ
jDYQaPvTMa/PXeOGs1UIOCjGlt1pEhixrepbI3ObQF3BgP1QS8+VTej29wS9VIKT
JVNDHRTc0EPShL05K/z1HXHUdcyatYpNx9k8ldCzlUyuJefB98siBGbfuLKtyLMT
IxJIe1jZY1BVu8c4XHmaHYHYjy8I3RVKxZSSV53LHPRxlFizZ7bLVxTAvru+WIh3
5FNEfB7rh3rmWGVa2+BNNLOIHfR7wnXiY1wmQCudQ5JCzUeI6Zbh/18FrkZ8Nrhm
pnuEXCYflDWzbLgdfXCPzi1Sva9XXOUKpyK3f5HEXksfBQ5u9icBvAxNZMPS0TMj
W962kxonReYPgjEROYNSti2xo8UteIs8SXsA/5jA9S6rPPiWhoG8Ajc/Vv1K+ocA
9z21Gdgx6Wv/Go2Um3QI0piTmjc/KjnVHYJalYf09x/v24NGZH0jMa3Vessslj4T
Qmcl/hq2mIyBoJn2ZHi1pm1knTSMJ0QQth6xHjhIjuplSv7mZbS3DlAceudg27mh
5IEd8zlzCZ7okVGklSX0TNDqlT7rjixZTPbOUo7zeNV/S/a9OF7bAnmomSllyn59
ohaEvbmLX7hqWlOTYrPf9/UluEOg62IKpPprGeCFAo7LwpAicJtnsjDvJM/1uKhF
aIsACon7HUlv08+ETzjrnuC+GS9dDJjVBwGHnIpMLNce5jbNxCBoOIChTnS1dQun
wCaBfROQ5xdA2+McsteEL2FmJylqosYuy9N4uzl8RyamYTljTCmGBensx5WLwtBS
4QIxhMGRaFcIbKUy9tRXp9QrqknXzLANY6mZIP8iu6mvtktd61HFLSAXeqKFqWfa
PIT+Bzw9jGJH/1HbRRO9xolWpFz+cd0wNlfzaa7IgvT7iZ7SVlq1Mn21vApjYd6W
6pSqzy2J5rc1eqE9t0aGZ2O79kH3B0x0q/m3q6EACbzgvDJUSb7XunylRYIq1AZe
VNC+ffk3xb017EODOpPHA/FH4ZEQTpl/DBXpK7W/hjePsEw2miCYxrtAki1Bj3aE
9vzyJoYye1SMR3DHlrbmnwd62/zlPfRwcstGda8nv/NVn68VIs0jKI70ivKHLbGU
YO8kLF52xuXVdMzeDOBP11c0OdE6dM81St25ll3DIViPG+pTQaxexgttJ7IJrdCB
xq7OxyvkSv/9VGPjWJIx20jV/AlSN/hFHrCL3ld4gnG/00G61x9FSMnSRbcXGXJb
RyBIFg3tbrmdF554AKR+GXzYzAiAYrft+4KqWSX/EfrWAQYPkKo5Rfn+PONcmNwU
+JFoLDkN3RqNryFYWlexTudxmeL7CMs+hNv+KEAO/OUSmWenMHhdMFLOHo6GSRB6
P/Fo7JP8xu5YYN6DGhrkXFQ39lPDJsqaBacwMpBGvZailnowCdF7pfNdA4NTD5BI
TC2WL5RVPFmaK1BtbID5yAFsBIYrhJZtErVL/Q3J0wLk7jnN+k3jdfk/BKfU+Pxl
LVxKTteZglAGwaBiqhZb/MLwYZDyhU/1DY4Yy0AR33y+XoYW44LPVosZUSy4fLsR
zStLAEsG7T5y0KDHo8r3Pv2O39ObYq/LdGl7Oo5j+nIi3jia5d0KM2aDK4uFraek
1nyeQj3zQxQQQ11oOkjB4sQGffmZbbdpXHejWCXFcXqHxzy/BR4lT8d/MvltN9O+
Kbx66PGJ7o5RqAi2qvOuZcaT5CQ7dg+mfwpYAWXzIksAV2s0PkdQGtlhzU/QxoU0
8b0Fnf7DvQa0zaveWAczuWckxPW6EAHBs0uT6KrZovyNa73ksHWpbS8ArXNs/avK
Ifup5ZFWrnSqlrR5PkAkqMVc2mbI9Eyc3uQglY50uL77EpP1pkvMx1wwwnDyP8VX
Xl5b7QDmJnq0dLhbx2g25f6tbVQfMpjAfrC5jnF9Yns8k19ELNwtT+EUt54LhgcQ
k/kL7xEalDG3V2KEJbWKyhSyxLWidenakVgPtTgafKsktbiEbW+NzJrkxfbl3QBn
iRhyZ4j3GNwDLsE/970TAU2hRe9maczYyqsoMndtGLVuUZVbgrTcZpc7HKXww3Ox
5AFljI8JATJYoTw+pZ2n9DYjx0ALNMOleswEGDUiNYidCjaW5A/NS6ldaW84nvz7
xSs/046aSDe2D4AEXl8JVkMyaOMilh1CP/+uQdWPvwBKDUVGBf/kQ79+ShKgUv7J
jUS0w0NreWGAgMHL781C2od+aMEIWNen7OFgDWn7aTu80FC6yWfayRJqZ6wpASCX
n/xlrDhlgiO6eeEsDs4y8h8MYSbj6oTfvvD4/XLPHwKav1Q6VFLFr3+hqzd+ADJp
aLPVTSs/5po3onKcGZOmRfDzkXq9qR+3V7usjJ9skH6jTAcuMhOfVgGYJs9wPy0N
VwQgB3FFC6RGbJNA+ZH+ggluxcHuOY2rv8lhlUCL9TrH6PIZQ8oC7HdLsey2A71Q
4c5tzp7wWAq/hgHvQTWzWiFkh4tjC+B67yk/WSC5L+rjjjFnxAB/lUpsnDCAeb10
7AYZBOhZA+IxwuAsTctpfUlgluttipTTiPZi764Hld0bE8GOun7GUalpRCsXKQWG
WDf/r33HipXUNUfzNmXKBz2CWWu/8wl060EBoFrx25vR7z7KjimqfblPG0kLPPjD
8SPbIP5DdgbjGuWUjZ9Kd/1mXKUJdAnYBY5lwr//du3pRRymr+UYCFvexKTCfpgO
z8Ib5txB00PIrHC9a+d1RFoPfBzvSmwWds6wbOfYfApC8DiRwQk8V2aZYL3XglZJ
6u9hEWf+yjYb0EucVVi3661CMZdQQQv06nLxUUToivLmtDNPnIgYqAwwLbgvh6W7
qMNaaotARtlcouGMwcMDSEkVvc7xF6xVIqyZfW9dzVQWu6V57f8HDCbwPJxxqWH0
J04SE45lzJGJqwDyW/flin9gYuffI0TA8oJdfsHHC6QZOFs2V9tGhVKB/YLIqjsJ
VDuLowcmxu0nym/MKRMksD7Rdmxa9XzeAwrFC7unhD+8GBfOyRZhrct34gUXi0qs
GnOkMcJ5AUisAdZh01JndR7cMyoxzb9HJKAtG4/S7E2XI2xpDLGbDhgjm0pCw0Hq
0T9h/mJ42iIqCvDiVCf0Ocxr9fXjs+mMRbTCj3X5BS/OMx6zLe9F0r322Xbphyp3
pW7EtGkmW6NW3NhE0ktfrxHVBRxxjo2VKtmmLq7xJRZDJ39/USoHMVSVG/ZTdaxs
6w9yBrUheMHSpyPIBr5pcSSoAoBpuw6ZZqa0n+WNa2icc0D1Mm04EVoVQ6zzEynF
QvKLiu2b5VFWZ7G4S1cBCaFlyKiiS53Zdw3UoQNkrDCXFNEPp2QE7UQZkScx93Ni
crOMYKmIBe5UiyaP6zvIi4FcPFokdtsk0apy5mKWA7m3U7wvFW9ZiGsp1kcROncH
dXUcJ/n7bcCUlChqZEXth96EtgjhrLX2rm5VDuU2yYJeGmbmHdJPhrc1aCVLd1j2
AqYYcGHUzdQL5/LQjbX2MCg9cQooSqEJ99G91TYpRrI0zgX1A6adQSoYOXZ+nJpY
dtJMdjrBsAaYW1K1NmCz1iVROrx3FZUwYAb0v7I9NjuOjg5XAN2vJJ8NsCMp6oDA
foAbGBzz74teXoqG86Q0+t7wgRvpe/aKBVbe5Jrr3CrcBcJ+ndlfJiTAQcE8mVh5
DYTXkjveUclIkLStRIuFPPFUKDNxXXY88i4DT69dGX5sXGayVX/cVvopqeSgftmb
cqRdy+uZ+68Uba3nfgtui9z45Qy95BHsmIfbwdTj0lykRS7nDgOYBlq+FQnbUsjJ
Qv/ZDG/8RKbB98xov+RcItkYhtLrUTxolM0ia1TmZSB79EHPSZHHRVCgJhbAuChn
FFQz0FBbSqz1taMhYpRu2PedB6rbMNjd7a61pOmzHao5OO2nmURgWr5+5bdfdj4r
vjQPNOuy6JAD5Y0jCtdnJ07COttjn6EjYc3iQZpWgHWvlg0Z3e20P87DK/xv1Ffn
yANp5vatNKROswuKgMsDbgms63mf5PsPBPOwU10esRmNkfmiRRBMUlsUtScC0NCz
Ye9CGw5yEADbVbP9inA1+92nYWSCfnwX7h0qJLsthJpHQYWKMbF798KDf7ZAyhFl
vhluvtRmcuQYczZuM/Bqyv60S1+WaEIacl+ieZRc1HB1eVMViSffnyIz9NKrjs4b
CIiCF4WYKCteeCyu8pnLX60yK98K3gya80zg+uOw4S5GdSy1Q6NYwCz/M/VqjdFr
wE98D4+73chHj34P7OLmwQC/lc1qr2kgIGl5YFNG0oCU4B3m2XRWLB9D7Wyq9w3D
Api9Xts3dVWtzuIW8WFlr4EQCg0S4XMRrGjpg/rdcuRHMunsgpoEttpFOMe9Gl/0
UwV9jwcPn3fRA9Swslg1/6C317iyAzOTYPRJOPgO9l8HxQKQ4FFD8JI3rkZAdCp6
1W56X1Ilcdr03F2j1usNsLWnutxHdzB21wP4k+L1ebnqjunkFTsoh7dLlYH7Gtx0
qD4eMSU/GPyBd785QLS4/VxOMmh5Lpw3Y9SpvtCy7n8qJcW+tdmjLU/iASN3IA28
Wtt4mRXbm7v8L28PU6B/UZgLHTq6bG/3TpH+KhvSgMT4bCRt6g5AnK4MIgIWzFHP
qCkAPq+hV0Au4QIIWm7tMJRZhWwXtmv26Hzfuh9f328OiSonXdkAwWNqfXqMUkoW
nZ/yK6RpL4hO9ZWfDdNlM29keTLnyq4K4j2SmNw8XVWNYi4xfNIQgMrpBai473Yu
riN/EoC6ZJVjc1Lz1b3T0Af+LHHBvryVJfmtRkjO7WVp2Xbrw9P+bh6yyun7BLZL
Nh2EGLbMjuJ32u1T5oboqg3lSsbIVsZFnkYVtIcSHj/JdgVDKoAjpgNW3UK2uCH/
4kO+zfRumhI0PFHKgQyKdVu9+6VR3N9iE58vVyh6KvVxtqIPx89MGwhOnwMhycMj
82LXUBNHP226a0o7JDjSlCh8/glgo4/dubKduBjkRzVNr5j9vEMPOIp6VzRFhX/1
hDBOvhWjalMmuFpiRY4cs7IU3vK9Nenl/OWiXjk2EEuGgbP7nPAWMW+VafaeVe/P
iUjiMdjuKYgt8PBOvZiQAxAYHo+HzR13rdZ0Er0ne6z6WY8wjddrOCohwZ0zRamA
/yfMzTBNIzmKlj/8u4ml6MrWzRxWajwxAjPjaNGifMMIgon/gxAFakfnjAmjMpDG
mtKRMJZizs1NFY2xwVZF7/7tD3IHWifPXvL3at4NgU26acYPtzxD9w+NJcnCxsVP
NwSWHCVIKU7FYkdLAQojCFPGe8ZlQq5tCIcryK1VE9DmsPABbV+gVV+MuHbruhJS
0bO+K2B+OBRHLfoVIhh12PxgJitYlhCELq83jV7QFkbdybcVWhWWppVw3vMopGPd
EGQM7ulTtCVHb6KCVKFp6bjhqHi46ByxO6l3frFHlsZ7k0+TnfsNSv7wTghz4WlB
xBz06z9cRhMCM6D51lHGe64N6mrbTGbgUGhqcgXuaCk2xGMqHrqgyGbpdbX2LNMg
sx1lbgTDYXp+IoL74eI4sW6B0oVHCtYeaMfF+cyUeDMa3ge7j+WCX592l5EisskP
HQAWO4oJYM9PQitui4HjYkFLfBvxEeIxDrGD5lu678eFrHwBvoXq9KulMGQWDqDN
MDDr/RPPUj5plAcYUKDIylwmCiIoPl7AubGP4/UuUuT0K0+lwRpIOw4TEu80z7hr
HXuDtyxSAfU+yiZd1ywQsMEmhatGVCxbVvagPO5SkEpPMtmujBwVQumTdHgqHSbz
oF0oHbprT6FZC8T3NXwQgNUVKr40Px/cQEsjToRLEj5qYr3vCeoFdAU6tybY91z/
TKHVVyjOzXKhDovM1sEl+ccmy+tdQIzI1IfyqCfs7JWWZqBtheC5ztYNkylH2Azx
58PuOMmWwfajkKnEpaaWBx7WsbJrqqtBRe/XRloLLNUFaPULQir0NeIn3IdE4LgX
z6OlVMtQ8kbYbJFzBGdkkWPTFvtpies9DFyu3GRZTv47jBQK6JQK5OUmVHVPYmrd
YIMJCqLBZkK7YMiVTxkRVgbax4NrlgdiEWbT1PGr+V32M5DWPlulKUoG01zoXVE6
4I23mlpp5CdpXLTl43HIIGDUf6utlqEwh9XFdD93s+BQ+7xQNEt0TRoYFCKWJmMC
w+geNWDU5zRYAHVEy5gGjw3N0cuf+nsIoQDA8+3sYl7exeSI+XbCyJUki7wGeAd/
bL3dyy84S3vqJE6DnMGV5PswQhrgoXwDlTJERAFE1e+xIW0XWhO2bkM3YjibkQIp
xD6Hg3W2e9JRF7bXtd30aIRWqkqrZM8aEeIHPXT2b9EFHhmZwEGEI5PZmiF9DcVT
xcLBmrv+QCf/qeaoEiY9/0J95kbhUSNVOtGIdo06TkB4XK1DrZx3h4NUGUF6JjBA
VmJE9ebqPmICc62U5LEIGzXL/OFgQwQ8Ej2RnYcUbEewwUR4YW4POYQmydsvsS8G
Fwa6KurKbqx+eCdnfMlSQ7LK9911XZZfTtqk4hP5VAo64+IubPgpzkUv/ivY4x+B
V4769zk2bzsFApRD7AvmC/WU1kykBJ3kvQA1/uvD+CsCstfBbK3MzvhYxPIQtjXU
RfbBWWdjMihY2K8CjgPAvXytX5Lr27+F+O7IrWqYzVezANOIM1DLpLw+bZQU2fWo
dAQGrMvDpum4Toh4U2FJM+Qfq/ISVaiXpvSyjusJMGd2MZjrm9ax1CBdOXFDOyIR
v1yvqHUbAQc+40sFyMt7+ziRvESUif44flw6qtA+cloBO9jevjcgqzJDsBk+PF20
zQaYgEjf5h98o3HxpSQx+zZ7BZUYc1VuFJ17FEOeDCo+e+qArtIASB01Xz8dIElc
/sDEX2L+Jvr8QBgURmnc2RiQ4MagyEUOIyGExu+Nr6HaSmSfW28WKliqo/A06Nge
LW1pMX95Bv+uhTeI4WyOLcq6Bwv+DCpTsIBVwEAGsvqkC0zkj4G047jWPAYsiQ2s
GyDLRHv0Dh0CVKdoD2XGSwUrPCP3sqIeKh2b0GWP6/7CiS2tibO/U1ndrI9n/TYn
3Zat2EEzVVU9S7/lbo+v/LT4ojF2Ik7i6FwFKLGjLLwPBG3SdrmhM5fSCGwY3dQ0
E0G04OB8Fgl8O7gUkru0xhJoGMia/9bph7H0a+Gj0dJpH4xfXmz4Nm+v49zK7WAD
FOIOBv6fiSeQ7hNfGVpO/U/9BQ6BrSibwMVc6+403dBNLa+Di3lgpmKANmJFUrcy
J33PK8ViIJHFkxKdYvsz6nXR5/vLZsFePwGgbxqwP+BsE4Vutp1HXuVfI1i0CrIJ
HYpnFMWE7422NR93WoPjP7/WG34i10ORX4h25lCohYTRwsC3vw56lXu36QWu1Jkx
6K4U+qwE7cwtG2xX3N6ODq/jijOfojomQ/eLH/bcKO9dqsCMfTLVjvUJjrYPP07M
7wXZImMpASaM+RPOiVO2UgLOndnJ8fQVRGZSu4Y/yIw+yYx+ohmJUmBsZaTizEt3
9QaO9kMrZo5teNSGt6lfO/72WZP0db5Mg8TTkA/RphmhGP/rlNYQkK327NyeMK0u
rdt1//7kchy6lZgMxTORSwb8HNWqWerJI4zIL7wNW6HVBKDHVmJh83+GxDCbNOsX
1Nv0x1QO/uWCG4Col+9jtPU2FibRuEGsXDENX/hfYeAZBjBlm9yFP0sfFz2cnXWa
YV/bNT729ds/M29AsXwp/4kdwH/pGQaIFvIYXutY7lEMRDQSLLVUI4MbHj6xlyep
HgxdYHvvMHuisrnpE7senmRR1s2V1tZBjyc7oVT0hfCEIba0hlJCzt6EdU9iq4Xj
03JETkU4W/mTZj5uY0pBqV2hF7sFzspkKA9O4OMfEjysF0Nhjci+1LpZW7FPThS/
3NW6MAdbnIctt4auEkKL3N/bvawE5aQSiKPR5tde1dxdJ/CWmgh2lgFDBURSbv5/
BDhy3N4IOytesnbImD5lPnLjpnsqTeALYmKKh2pRGz4XZOM/55jB2G1bNvhHhCEj
M6iBvReR0YIqFax1cMkWSca+fktNJH65+Vpag0uFVyjPZx/4YOF6GykE6YK6rjoo
UQkvn/OxwkZZ1SzTBOhfWtkSCfMXv8eCm86JkAE0Ss/yYNHovWhB5CXLCBMyhl5M
bTuD60LPBA0S6B1TsvEYDhWJJTc+DOhPE4QJVfJrfsOUHW+XQqY/+H0aiN7Or5nd
fR8YOpmzuAtFtt0zNxTwe7rphjOs9Bf0m213ZhvDwfxE5xT79LA4h3xEgmdt47Bq
SPgRv+pm7xhJ0pwX3NFoxTtqP4ry5DtA7dddC6vcEa2Y9uVjfscEpksCWDVV7Axw
vFwWbDDP3hQoW4UVRcCvfzarFimX/n+CvOF72NT6fGNd/uS8nqkU9GuF02pwfKV0
BgCH9R5Bn91FzOw0pKrZdYnxc7mzjaJ6rhEQRPA0Eq1tvb+HiqsmpmHORhPzc0mF
gLRkHZp7KlZLqh7GQO8SJcEsD096X3b9nVKJETb2w7x4cpNxfswfoIjOZs9lM74/
sDg3qzWS/InI8s183FXBVFM8dNrM0auMXQYnmdg324EK8NQonu4PFAtUjs2w4iqw
N8tq9pZvx81FOxBt1NRthzzaCdLtG9ErIhfpynFYtYCRzwQ/i/Vx6AENiqps/ayS
DJdqP/1Di6qmHPhsX33CKyrXriWAhyHq1mR3AoOe79gDjsqztVtxw/2CBLxEFrcD
JSM9I4yQyDDNczILK1nW6RPFFrEF/gbq5/NNXvCaioCwyC875X5+emptzC9QPKdS
sF/xuQ89h/pk+3SSN0bhy9LMlnTKMD6Qo1AN7YIMlBjamQzjw8KkaM527yFyXB22
nKE8NZCCo7rzPfF6X1Nl+skbL/R6mQGhquH50odvb7gOcev7JFuLoQN+GTHXLz1D
n/+7k9HNfML0w4rR7nE6Hf/buXB2LcajfUollgevUHyhJ6FTIU73ao3ThlnYu4uG
liWtqMr866qjNTdX2BaKwBMCUE23tAiuNVM0lIBKKpmH1OHtMl13u7ca2RjYY0zn
GyP4R3zT5vDwgzrddbzAOKfDxw5jos1SA4HR8utR40iWARnU8eWnaTEjWJDJTQsb
hJ9ZExRXd2mEYgeYbV5Z2cIQz6f8IDiNnhs7K2352q5L5thZhYVazoZMhnei28UI
p+2wdp74EKCLBApHmz0H9zHiyEFO16fMhsc/6kBhVbkdiewwLpKhu4GYyNzRQ/iz
yygwyg0vinsG83+DJMpid1y7ajOFmcaMWNBYIo+wttuL5dskKHv7xnbJRyBGqUEk
txITnIntxNyP4s1is13OOT1NiZvyd2OdMAxkUmMbhYe1/xaLzmW+WY62D8fGXTLK
4IRXv6gg545xEf8XGvUBiJ9jRy8jiH96gEPfoxLMlduML6Rom/6cZjGYk6A+9ZJx
6DCUg8POiWeCMSmE5cTLleFliB2FIvQHFhjpPKSs0QyjL+Tf6Cv0aV61E9XSiVyi
Yh+fAx58/POSHCMpWiZRLl/MGdTP1xMIohkJFCDOnfjm189mNgD4z2c/pFGprjTT
1fmpgb3f90+BVdtycKQ5kRIWIZ23QJSZJPVsZPs8eESQB0lWkAXWkQOj8cz7m8jR
P8KggbEfZYTqafpSi/NNQINCnIvuKUpr/Mmv8ZxcRHtiFdCQhIbiP6uvhdXjlceP
38gKN+BK0XZLEGyka3gcwVPoT+gZiPuuJW3T7Uz3COSE80qbkxxaqZKPvtJROOju
T4DG988Fs7BlXuruJxWpHqva8sxTvf2rL4H+pyjzsMxTvwrZXcroiMqH9YkZiY34
upslnsH1d8Sm/8mP/VlVZ2hXQlOoPYa9TfzeTce1hn0xMo+nAvSwwFIQgmpr8P4s
lxHrlaGrc0SlCXkJcrdA0ePKo+y3g+MXbmHTJDv678SFUOLo3UI8AlkfwEX3Mq1E
gsUcPg2uysmACXlr+Y58mNUuP2Mskvd9I0T9fVdjP3I9mtSQ42M3lfMIPJ/walic
/jGCW9Yn5IV7WsrkSdI79qOdylIhKFJafumkEj+Tl0+03Nkpf7PqXiJElgZ4YqPQ
l2SnZ6CyDjw6hAzDvdNqNLOi1xhcLJAM0U8CcV95r4KvRRywRXVrMqeN+BD5z0df
SUkYFlc1JAQ9F+dOXQ9G29UnJr8uMRkBEY7OS6utFPSI1VB0C4EzMOEdj6E740QJ
tlrK3H+97qYKNhAbL2//VShuI+IRgWRU8yd6sVrfsuNLyfI8pwQbgQBlBCMJ4F0t
G9gizW5mnfBLk1hgA3ogDQC9aU2sl5Td4RWZ6aGKE1b4Xk9TqMV47NlrIRZz8iB5
P0rvAAR42RlElfYuxcmv9IczLYFD7S94ipQ2bTgyKsU96CuL1Vk9Eotaq0ZoYdwI
1TZSBZDfPmAKar8vWBVi0oS6ARk5zxq326jJMumr4jpHkcXkxPOMU1GxqO7qKox0
LOBV+Yyp8ItVh+KB/XtE57gnGAJrsAUx75gsr0Ue+GcXUSQyKoq3cDqUByTu0Ilo
MxYGSqAg7D5eIqeu+pvMbsJyF4X+VtlO5NzOe8M0Qe3i82Xsaij7DFMKKB9YQLz3
ZFqLHJ1yN7mxW/c8PLYqNFFgvaCjL9kOb6jsjPTz0xAk0w+ddsB3Z+7T32Apf05w
pgqjlHyrJDxurr+IdFN1pDKAjd/FubAIgdnL5GfZAiXH17qFXcFvtlzWcyzHEv+J
dX+Sp2En0ghSVTMtgBdKv9lVrd+7nIziwcPCh9rRgM/C1uxXzUpiaQDSgf9AKOzL
lblNJSdPGVIrrcaI77yl6CfSRIgZPKyYv8Fyby1p3PdrCHY4lvZj5tg4TMGfmcG2
4tTYvqz2j8E/O2xRNgfYK8sRzD2D+mmnDGOIRYol3dk+c7cOweo26HNp4uSKwpq1
QuaCYiWdFpD7gSUKkmLWbxC7dqqC//AOstzKxSs8xMorwH0O1G7ceraHJ4yFfN0H
9W7ejlgXRiqxXkomSiasFHbLrWxgV+WMeTpiXhJgmTwl8PN7tsWQT4KuQpJMUSyw
8EMvVUuIzW9AuGJPGnYj+M7c1XuFoJO67VnZKUDKlbbwxs/CUK4GwV6JxcR5V9B+
cq/urxMAHiUUFCJ5vCSovR5fYedRIvwb3fzQxKNJmRsHZZvqJAwKu2YiDAhh3/V1
WU+/cNilqUGrHKc/JrakyHh/C8xjzcYz6z+OfOsKbUQt0hpXcfzz02P9/BehGTPp
4ehC7sP9V0zxYOWrc8cfIbFYcwT3NnSygIyLuBG+y4/DJT5BWe2axGY3JMucuA9p
mqdRp0Yjg8/NTZtcSG4hH+ZC575INVIpPqVidKoNdXghETPo1xY7UMIiejfoKVkk
menqtJUuiiX+pDGAl7Nx+6rXa53K1zshlJzDvf8qaHmSWFnCHyIxkbcm6IJ8sVLi
OpmBSsa8IrvkbS1+aYQHCO/bnwQkhXYR+stNvcgI6wm6IU6RBXCZV/AahK+rm/+W
YkHsfgrjPDHZL1RpT0lhFSURGHoStSYBGjWx/kbYbyDUTFxs1tJeyJEjtVAZmFzu
L3DZupUB5qiUQG7lJXZjDHzJdR4Ud4tN0F8gn4U371dd2YoGaE0JpUaJ3/SnBMjQ
a/xPonXkcp2D2IU+Z09Texj8SUJaCrNq6o+yOkpV0wdODUfSRtZWZnXH/Orl4jui
zx42ZAd9RX4BsbHDVYtZVKuiuFYDI+Ynt8wKWy10HUgwYTKpux9Lto4+HX559Im/
rYG570jZftmcCVc1qXUMaiSrMsI6FythpVFr60F9QjfvPnavmBWvZZl+3gyT6gu/
fjfk7fS/lLAU5bQEN4rzI4hc0efQZtjv2o3CkpL41gNF8+3iPqredMjTQKCyu290
pFBcgNdGLCBC2jvwPwqO/fn1RW2m/j2Qkn+dkwlv7vINy01f9CWYcO8dlzKAmFI6
Yx7ZOjufmEZ1E8oVR3IDpA7XcX3OLWvSjrJ5bRWgLB1SqaxE+Q7UtcH0jeLoNB7h
SRoLzix3T/AMjMZRoUrdfT8dcclAPsRTnL4Dkeseo3yf2TXzfvrh10gr3Odaexxi
hxty9jzsiw6ypfJffOd/nvMvbhQVg549fT3D2XnSQHrPdLTmctJ4izdKPKwcUty5
HwtRbhogSrbIGKnP0eIUqa8a8ZuF5+GIlOAk9onZ0cl+30VfHGf4/jZhcGdXRv7z
fY3cTefVIjFDhV6OTT+KN0pYZiHKLwKOzL0WxPm9oZEKBguql7xKk10LpjccM2CY
IFw0aJlW6ckOOFS3klxjfTnyw+l3dfRuxL581UHWw+loahwkoJzTf1cVnOv0Wezm
a7GwlR4BBj9/QzcqgbTtHsM9bojUL16Fas4jIz44wis3l9iu1kryZwpa8Yuq3AfT
X0SdbO7pGapSVSkFjF1Gb73uW7Eu2G6lYrERAtNA7OGMmecXTXFvMJO8JKRcQoKX
4GMWUjhvwlxIobHx4IXZmYCJvIeew92cjIWpEJEc4wlUgns4eLR/z1KGAiQBH6/P
WMkDJXq+R4mTUAFYvNHrxcmuFtNGkSp8istjjml3jBuXiWKCvmQmpbMt3epv1ZX9
FygK3LWXzTRrxfZMQ2JJoylB20IVYdEjf4N1t6sVRauKsqmStXdcDqF3gdQS9940
BM8QVMwKiZAxCMqt8dLqhFYCmdS4Pqwz4aMoULqGbMqdYHIM14DoTFKxbZhJ1x0n
E3Kne6oxNB/f+nMLC3ezNpFN8ggEJU7dZ19Kx2TbYGGXVmog30u4b7SnAte5s/Mp
NYDoJKV00835C7pPRXT4bf7K4Ibdx2HG6KKrAU73d4EJJgQdGlzDfLgZFi5D22/j
GhyRtdeN9UrpBeJc4lO/bje7mwTiaahH6TNQWQhd58yiHW5C0XBUuj1VbBDnpHoy
303Vg8KP1WgrvJqpQp9GS3C/NtobQhjF1zw4R9qXM0nHpJPnqoOIovM6o/IXFmSN
rie26Arb73Ml+7yZQDmz70YUBvFzr+J+UkNq7oLtb4RIB473BctIIksaTfQQvlXb
reJNPlEvEDANk4Fs+oO+MGZtOgQfW9hjdr4PZ+RR5IIAfwjwtkvwQWi52Ciz2Lhs
sOKvRqK9iMvz33+b5FYufTRgLDI5Dau/2P914yqJkai1Dq03zFzk7SnvDqVGCpdI
TCGHDdElp2FAnyH9e/gwbxUG5oxONvA2WCtU7XbATRSDMwuIbFeG9qucWnLzSpmf
ZdlDOvHEdcc6p9KjjtQzJTqcH+hrRC+B1+iavAVD7im7SMDQs/DmaURrvnVUGA/H
651xoM7aWBGY2xczoKQuIjEISNtCACyWzDSIVK00g59iUgX5D8MzxIrCoSrAkgXy
gnlPRWFsuSM6zFXlDvDp3y5zCdhBYxoseMS2qQagB5PWvXAn4M4/3ciPOEqbXQju
mtUfKY8cfWx9um6gyPsnUXo0ZPR8T/ePmUjBOgZ6fxLe3jG7rkgPuU5pCT9bVqL8
ZYX6hd2YLjgXZlut0LbdYUSB91CzCDznpB0y7vfddsudDxQ4X7/HGk25IMfP3ywL
jdlHKvr3NHhe5WdKdHzmTB20oX5RZSDHmTgJ3tMVg/WbWShIHL7pW4x1jtXxDkyq
e8l49H8ysPuBXXLjwtlmpj15d7uMzEp9Vfy3gXifHgW4XR5HFf+z01smXGKlZDfJ
Dqzk/rvw4+EhC/coD5/T//ZmK03+dMt5zhURjT56vajGTJXRiDg9vYM8XhDJlgOm
zZ2pSLyodSRbKRBEGz6A9wX8+q081RbxYaKb0in+delE/LuSvmfhm9pfBQJJT3Hs
xlb8lgA3HpWDaF9vDQxn1V9QvmXCYlsns7/7BnO4+d0yQL48+qvhuHuyb2aC/eVk
Ek/X7cLYCiRNkBRrT6DQUr5QLvc3FI+iAHrDEIc0SIDJHtMQT7RTGD9e8VJMhNKM
3Nc2TQCrtk0cv1bBNsewDHvLmcDdj6/6ku3C6j61H141v9I6+qdXk3N7rK5BG466
KecmZ3K5pSLNCBmMFpnP6j/W7jWfM+khJ/wDIAl5moC+cvctIDXZpea/IhuNwnNt
uqVC3y643XZpzQOUUQuBdTVUH7Xj3XUmseDVibz7DlBT19eH2K4tK9qJ62n0wXqi
m6g9uCTbjf1x/PpiXepmj4gtis7I5slG4AW5updV1cCu9Il4y0DA1pbl6+5XiYNS
t21e/yIIHrWuRp017fBrDlg1nG6MWH5Oc4uMPMK9rNpv6XWqMcPTC8FT4XRP3m5N
Kd5djucMkBSx0TYsD16K62VIUiJj8HpCMYAHqJZi4Pcgtim0ZbJp1mmPBMQl8JGR
UfsP6qnXXb2aEI4easMBlP7NP1GNYLIYdQOBUPCpgTqCRFTi/1lFxpJbJEv9z/zy
WyDeUDblUMhc96LEri8/94CBeGNd+alLWtdSIDx8FcVA5rT5wEAOTD0IMqxQA6RA
ZGzeoR3eyL70HvEArIcpA5tp5MOsRBqXVFEW2pXk6lrIUHpWZ/gJdc2STdFnB5/B
AhsUwldvRemon7gaVtYywL+r/xxeYgUiZ2HF7fR2En5ThhyDne83rJ4FPoUNyBZr
Q/v2F/Ldh+BJqtwvtan/xeVNiHbReNDfo3Z4fFqIRBJgnwbjbBUfs3p4XW/VlMj2
AsulUtDbxmod9Gj+HQZK5sSDyQxINeQg62uNGMhKVVaHnEme9ptClixm2aJJPs5R
RtntMHDWJs/tXAgg3YE5xlxJj7FqawwsqgTNnTCb8wJwO0yJeqPZsKe6i0bmM8eB
AzoF28po9JqTs/ssKUc2sppxf+lLmhDCDzxi+y8uw7lxjqDlQIiSY/cE0ao8LxQF
P49CT2tA5Gkh1OO6a6ABDya2NmBJmng8cMR7eJF38CpPQqsWoK4ou4CyKnahU8TY
r4Zwb8CaXV8os067hV4nwCVXi79l5chPvFplwL6DfQfPg6/neesFr2Lm2zHkX+ve
SFAEzVORZ4ieuWEIbMpQLNRLchjBNsHEggbRk+arwVHlhNe3Z/1gn+RgdB3kJftk
fBhUGI+zbq6k8fH4wvNd9FA71JDpjPTJXuqPW6QnzWbdVRa9OEBjBm3ohXZ28M7E
lpOnGK9lrW7qBnthfR5UbP6RI/ZKFNMqLypayzWZ8a3f8qE5iIrr6uxPG/Faa0wx
ooFxPlwq4riSff3/qjEACjh/Pk2dF2RaYIhwmNe6ZXEQ8BhMF3D0UR09l3RIobxr
6DuE24Jfbdb8Gv1VFxuPvz2YfOzycGQQ7rr6mgYnMRBsgLo/v3mHVGOtSphs6TcB
tOPGtMkSBOkPg3DdF8mgOQ16iGXpAu/6ly4Hg7OxsF3IwquR07yTRok5B/IQSQ6E
1oHVqsCU7PKQzL+3fks8YBTTs3Bxg0GSm1qm1wECocFrE30Yp0hgG7TtU0wcFVoZ
CgS/HSYPjGXYwlXEdJapxAv84M/MvmBnCU07DP9wIgBoJVO1Pzfgc8K3Yp6lr7l9
74BVmqrpgV5xYa+Kz34qDDhdskVkoXqaHfIydVa6sNwD4dHVyMbGKHGqPIcveGw2
UHGaak7egvwdvG646Okp/ubtBt7PuDXlrTOWf04Y0GV175sWv03Y0817dfs5FcGh
uioC6hJ2Xi7Vfq7cbdl6VjHEzgDrbmFaVOQ7VNBi3IpJwITztiF5kLQKy35zL5EE
iIvkWVUlR04akPKlnjAYcnXc6v9nZfva64DQgaJdwKE5Qmvxi/WAjJHSMkhpZEUI
zmf0t4CMnhI7hvlOw70C3399JtbTC6I09p3OU1wZnKxq0M7KqgJNWzMnOQMxNHhI
4ObP7mPuIy10xpqmw/WUX3gEMB/4T5YbGjD82Z+eC6k3pCwpeldfkjGmEOeOqhD7
W8gb56OSrNmiZFLBokYoiuN82fChsodi70IpAkEF6zChNrkKRtrteVkYJtm2ecvE
/NKIvcXtosHAH2B1YQZtcas1f77iCqI3iZ8ogKILFoth/0gTZKM510ouMFrn6I+k
N0EzpZoX4QpCtMRms4zhXdYyYa4Sf6N8BnOK13lya4W92geoT4fgG0aO/oR/L4MA
lyFNIGlxi46oEGU6Uin6a272g7zud9xbkONi03CKgJjKDcc4qVdfNlyzzL6oCF7/
3eMHj11h/xpKujuuEnQ879MDwoFXQUuiXu3zHd2UgFQYBN9W4zFxPsX9ywc3mZ5s
YK9fs5Jk5xgV7O+dcWkuPRJadtfian7CnH1BQKM1+gyvY1CqFpuvPggOdZNo00fP
8WVN96QRMPWF5bXsomI0Ll/gw4GfZQHeuLrop+HQAcMTpNV49xh8vbNFa6X/bSup
OJvqJMn32gfuzIrpoNFE5snAKXLSRxWiX8ubJ1BRmH0se1TXe2gGI00k1/TXi8uq
YEgfcZpEtfwjGvu+h0/wng2ykXo7Th38Ex5LWEyXQ+blODZkvYvAOdf1dcp3WbMj
yn9J3seRArV8WQL2F3HOH5U9P2dB8imcK6JhfpahOmHymJP9VCaK1/fFtHRab36P
KtWN95qswW2aU6qb1t3Mzyng1og6bDPw7ROJQeGkZY/7t9oL8TyCUTFZqLoLDJUu
VTSv7WU0HxFnmZkN6sjxK1G3X4kil+hMANCZor2u9pOVn84rIDKNt1dGSBQcQcy9
5phPfiQ9Qpfr+Pgkk98kVCOaOIMhuV0KwEqZacB9zJk89IoyoRz326K7XLj5AW4t
MD6ubp4xPLMNyrbM9sB4NWo9W8+9VaHr2jchYvpUhYTdc2+n7Xq6nZKtHm6zgGMn
R4yscc3fSGEW+dqTtnoBeEWO6EElhSK9tQZJXq3b0OX+DNT1iTqHd2pbpa3u5BzZ
CSO8LlpG5HqTGqZrt+krOfKChgEknKPdNW6xNLtnuaF4xPtJ7fTTr/WNP+4lk0GO
phu8EDmuBRD1lpDRbF0BRr4Li2BbQqGGY7KWvtW6LuUD7F7tIny61knseOlHk5zG
zZD9d2wVIPuhvYwugxaHUB5b3hF5LcSa1jNU6WjQ5qNW3WMR5LDKOZVFE+QXf47a
BwZW4+zRa3w6s6JFgTW8tgpj5YvnVFUfDCk2Btu6OP5N9E/xnkW9Tj7qMCtBtBx+
QLD3D7orckhBFgL75mpUMGqGTlKm/6l7Zj4DNhKjbLKYE5yfaWThF9JSLxyGaEIC
ZTzrOTu+mtvwLjshYfaJM1WO5mJEo27z+7Fg7uQY7SGC730Ay2ny6s8WeYMyVDV+
yrrhuye0dN+/1acKZKIrSPHyBxkVRjmHUxXc2AlPt7w0ncQdvcFO+l22UglKIM6i
1O0U2hdEqtARNg9J9H6vj5h/fWq1XmL0o5W+/X/ch+0jh7IV4MOrL2sUlVEO32Es
hLFTMVFV9BFcKlGDU3i1ZT1620fS7XD3kMoAT/K6Rgl7+4oiokm6qI3Fit6o4FtH
z27bAGQ/+ClS6YpdwrA9hEKtLrJn+n2hGD4EiKVdS7WznPItgoBeiURLS7fWIS4X
YUYzEMsuBtKz+WF/s3d+XLS8ed3aOAozOI6f2EsZBzUfW2iEaHCylNLtf8qHcLgB
sy8JbpIot113gMs2Oq7/90foeUgB1hYA56ft37cW4e9zWHeniAvfK8p2umnkOc18
sdkCPhAyxv2UNqLCah+9mUdCe0oxXC0zIB2mINVK4pAqRg3bkUq2v7LM+GjHkeBF
9gSjMOTihgTtbYCFCKOkUL7bQxAjyvCdAfj1wmTwnAlfL0fYiTmZvcK/Gqq6XgA/
E8I2V9XAtMZ9aAVG6nTeJ8tdnBr9q4ZHdFIricu47X277+v/mHaRxfvnbJ3dsao2
o5Hd4SREtAuxEJTH91NzNjfD00k19Ji72sSdFYTlnWOVlDKdVtWWulKd4zHm09gt
GG1iTkTE4JWJMTucoevlCtNcWBemvAla4q3vYcrgJwk/UvgEIlSWyuTThmWg5x13
k/l7r3QPF8Cyfb5AAvZtnJHVXg75Ypl4Hxme9Bt9VNXXgXcFgYSNcnS6LXlsXwe1
bIMq4qMAygJIWj6Q7H/eAg2K2XrQfAc9Hlgjd/GchXdxZvAVRqVwwCFZ4ZpEzqZm
1wzWfa3BX8PLjWp/i34mBbGGuc1vwaT/Jc59ObO4+YHTx737y3JfZE2UauZRfxR6
x1e++h3Asg9J/wg/l5S2zDStmFPEc/KLV3jt/9YinaMgGtSOGsMon3B7lU0gZ0xN
qe/8pUYbMxcTB1lfMfOlSQfogvSLFaKsfU+blAfADc+bfjYiI5ZNWvE+LlVy5mTR
FaPPgecxtAzPVPF9xoXa/R554zmwdMRW1VxNYipg4Nb86p7uPokpmfOnP1zZqx+H
akhLMjX96xLPkG9UUnj7IpZDWejY48Qo0PSvtf2tE3R2WwvuxHs/1pQXoJLioi/6
/0I9NwaEKKHpcRG/m8TVr3VZk59ckdgD1+BmH7bXpwMtpZJpP9uc+ln8d1C3k7Ba
DYRc78QshGguMorWG6ykr//v3/Ftw7G+NM9L84ewfhSuRnZ9v5+Dr56yonE38UZF
2E7E/jIx/Rx4d88i+0DQ0N4O8pLeVwGB0etKa+CGKJun2V1z5XSTabC28k2qcVVR
bKmD4O4Cj8FRv3jYS15+ua26N6U3GhLqoWHBjLhYg+k8WcRAeEjZbODiMsGYIQoG
Cz0LPVpgKtILg9l4q3m93UiGZwGufibdXz/pyFFCtprHGeAXhyuzgizMyq0CrU+Z
1/mgYi/LWXbHQkIidVKXDQdphzV4qCd/paWS7mlre5jsCD6qxxtOkqgZLE5Y/GRB
2WPD8JRLBzG6SvHWtRGAYC/jSJysTUVCngSWTdctL8BMMBZks/CXmhEVKnHVxnvA
CuGinQefegt4ZiMzSok2qmfztMF9fU9+k2dGM/pWKQKw7tqKcrmfhDATy9qIeFd2
82aza4Z+QzVSYt3gudmsO5oScTehW9YwgWjgrM0FfLGV53jMumzoF8Ht00cteXBe
AcXCzCq3kUGFc+CiY+2PbFBebGnX7RgVmGujfFGORsMGPOs+OMtY2m1uVJXzJnXk
Vu3IQtu73wqS6TLTa0/S9AvQWlWz1LU0DP+MAlvsPJstA4x9RWOFYwXtUgPkZbos
mAqxztg1Ti2yHx6BgKdoJR5oVGCoJrgBQwuTuDsPxDDTWUOpCjADKu/uCqFxxdiP
ArAT7MrqXedtecpxEgOXvFl62f0fxftGTnphZY5BIHMlTZth5c++CMCyumcDJT7p
nCv8waVM/vKJUvOHDcJxyr4vCj5iPPsVEiKcmlgxDienzHeH67QEUOVDf+dAvc81
U2FLLBoO4tBack6DJTmRo6ygGJrjgZ3DS+rGz9dhXu88Z2wq4YkA/dY9OGxrS6EP
UAgXHyhAosQwkDBpN9XGGYZFCuXCea73BGAFv1MAgdsqhrQNcn56fr8B74b0jqxW
Ek8WLjh58pNbY9O6oFyn5Z4oQ2p13tvG2vWPIyYFeRL/cyURFHf7aPS9qD2bIIQj
wyjZObWJMJ7TMCutP5AVpd2q84weD+5xxuFe0yJYbY7Wc160uzSQx7fHlUx2H3hd
Gr2dIWxouDBbUu7UvwUVZsudNE6CVVNxS1qFWrq3MbhpBcSWbKd8vq9Zd5dy78UM
/4Jw8eRS2SCLQ1posXw2XjsPaY1DYqzxwyxICk7RjPUMjv3wDvJZrD+ymsWcsqdJ
ehSLjcLFmOBUNzi7C/Fwwe+R+/zJskQM/k4UuygPdl3Yv7r9pyUGvtKX3GzGZ7fC
0OTylPfOku2Zk5OXiyKPcLqPLahyD+sQoabJ/BApArvYY7bKZ/RO3//V9Z2gdY7E
h74rNAlD3esF7sLQQLH+mjmP8TV+86R99P6gc/RhSIGVKHpL/BFS5O8Dv+U5etK2
U0MTYmqgF8o6vTwyv5wyDLMrYA1vcKPAmonxWL4kVnq8qHOFrvoBm7aunxoz6si9
68IOWmAOxALjD6ttYurjmpADrdD8cyInTeKOpF3IndzfX0Fh3ZUToIp/5J6heBbl
TCnihXZ3Vf8eXDaH30i74BNOGmlsjE4ci/C6IIjfhIcilzvaVN+CsysAs/6hOdxL
GLc37C8piBggequdE8UQA7JjJBobaBm77biWQ01eU5juq1V26rH+IHPaXPLW1Pgf
skdmBO9mmDb1fTtThNEdTd8/MTInp+pJ4mygEQfec1hnQnAHwpCw5j7KDMZGh0/A
Y/EapY7hhEV1aqoEtorE/sTcdsiAYWZtYsO0zVjRc5Eqi8KQ4N1D/KD5tWu9gGUv
hqHtl7U6xVHXkNu8EYU/LteV1aKOzouNx6QIPgUPvNIvIRcr+bg+4dPbx2QhM8ye
TRLbWoFVReYBjVZ7oOeyeoutYvTMoYOO9zOIyycPgS85KGuhgDaksp5P/BTAyv5r
u0HmO9ISXwzdLBkFzfy4sCzc/20YXT/PcDYDvFSsLekiHOSRfvUJ83TtKdWPE1Cl
xzjH81Kf+6DLm79SiLkJcRUdVG+ZtiMCyTSshyrB5HmQx4CAgaZ8CEB9HOvvt8o1
vfJDTWtegXjW4h2bVQ+7cN6/SSWI7/MA2Sa1D0MaLzruPrYt/IwHCfJ9uX7bjZKo
gpM4k77+haIA4LlyG+0gY7ENgAe+shbWqCQs7vzZjuNeW/4ZRkmFJBUfS8us4uEM
NzXlTFeDUoEMh8bSSsNZ4cR5iKDjWrynwi9W7Oe9/nfbZj+rHc/ZXDzNB0XOf2NP
LZFNQo0jGs1av7s8feI7SUmVerNSFYwmSibxrkAYncUYSaR5kO3t7fmsp7S/3Un/
RZar7mHs06cSgEyv8iX5SIHhR3F/lLbf7TwgnCMbJz0l8nM89ukSq4PJjXTjJFYl
Bi45Zgw7Myyl5JybC/quriphrHuzPbc10eYr6wOEywwQaF9o+bUmJjXWLPwL4vW0
GA+/XoR40aCI9Nh0krRgDuQpWJzFMnIVOtR0azYF954/nYSJeJbfm9sg7TesYISG
7TlXb6HMKbtm+CPycdvZz9A3Swjul8o2n6yAg/NQEsa++PaIwMROtm4r4SqWf5uC
sJfBNSRhv3dsoWBuh5ED+WjtnRWVm/LPni4697WmRGvBGbpAqkOr6cNRWSU59UIp
uGUZZ4tudiK5RoIAoyO0GMn6s/tOD/uyulWsPdxTXSgSiQwFxnZcAEWa2pbLmyk2
4vSkKVAaepY+/zkOylCUYRz7uV1XoOk7zLw1ret84zZdhwXxN06JHroBkpYIHUWL
M2XV9d5wMcD9oM1uJ4rZJTR9JDoxcYYep2kwFUr0rqtKsVuzMgPL+x5IY/6P2Y2n
RuoHar274bxWByIeGbF+IS6xG0Zav7N2K0nmPBlMHcCEFfkppiDGVOwPwk5peQ1d
gfFxa7aj/5jw7i+iygKxv4BupVc4gdImk1YOnVX4dqgXO2eiOggO5Oh/Ra9DKD4o
gQjrwWQs56b2ZC6naTUhUjZR6BBeTTKVWU0QEOz1dgRTXmhH59xuiI/ln1DQS+Ij
YbFfy7DEMH1RIpLRcesXgnsC8yc5G5AZy+EPSaodNwhAheeJJphcZn0XqL0R8Tjq
g/MXOEaY2RBTdCIjf+lFdWHOnWCf1wpyh2bIZ+azwY2nHNR3RaPjErPDDR3SaMie
SNIisPQgibWogoZvEaeOkTvcj32FdOZOLCUBgPVH0H4oTgt22KMQ5lxi9FMx3124
iQXlEHWPjNamWenw4M7CyhoiMq7UW0qevvsv7hDY2T7m2JQym5ZoQ1XiPWMm5fI5
za5N5xxetq1O8MTJbZoV2tLxqwZztEBotHUrcHnm54PYGfEDuSl9UtzU53NN/AqG
9rJH/eX7Xfwp51zLDLRckB+5yM+jDC6CR6rEak5GVkXrW6kSI3KJCCLtFMq1W6Zo
DTZcyZNuKgrX9aOMJTlvYzdvQIYQLEhFjcDbNTpmAbBURWdXEl+6rm4/PQ0P7X4f
S35NdITb32BVLOrgcH3pWBTW1X36o1CGJ0n5wEdB5jxTQdmlTYO5gc3koMXLb2eM
joV2fL9uXZgZ26tX3xRxmdF0StZibeBm5HVjdJMi5ojtTMMpnLb+/HfU/1Mx3hEB
o0Dz3z+ZCiGe7iuz4+ovm0ulSnr+Bah5VSgRyz6UKs9QFSVV6TaR8uHk9NqgV/6+
/yYqNAzVpfjoF3oek0IL8uw25H4j4W5+rSqq4yR+tANN/B0iWYlimJekFOLh4iw3
u8ywFgv7biRGGps4BEgTpUi7b8fGbw6MNSt1jO85Nj0EEtZz34UsOqRTSTnlMucf
t5ORUgGJrxzFJHCuSfs3oP/PCFFubFDsnsdD0xFa4G106MtUTLak5EBm1FEKGJAu
iNKHf2SZk3Ldivp4vM/s6Op5kZ3sGH7E1n5lCUHHSMpSJl/pUIgJdyJXyVcFS7XA
usHVwgu60uUgst7THx+HH5GzowZ4qFB7B2T0ifysHFhTXEMdXn8oI7QGpnD4+Oi7
+Iq179NhWH4pAOlDsGw6hC6mZjVpXqGCSO95Amp/kMiqi3RatCSxxLLx49Tft0Q/
VBQYHmQoulIqRk5HdU/4HVMAPp3VrYHYuCPixxS93SOzPzB3FwWeBH0XYeHrV01I
ttt+2dlYpC+ic4Pi3quyZ0ST2h7U4MF+DLnKLrSTjoI5ZZsZXj3dpMMoMMnX92ds
bRrsXh9YrGNM/l0upp8Vx8oglo6e/SqDJeYxbqfLbrFYqxPPA25SyMFCBUMPh223
EMAKi8HrrjhEiI/113wBD7O07imPDAouNWCKX36BcHsSVspjrjk4Q3o9M1R5c1S9
bD20Je/9NOxa9MrJwq6BKZq0TV078xXl73iy7IXRpCUIiS0oksYfmkyUSiGW5Cwg
/9KtsXGSCyLXc2JPlpUDo2m22xdIMGx2Fsc+oiDTKStT+SuXYlaXATOBG+sdIQGn
ZCP/Cma1gxV80SadxI5c4A7jBY959DisSXS+R+mnQ5sZVI+qADpmw7us2TrBlDHx
pPGSCxc8zKZL4hg9PdDM0VO1by7Gh7ewhOWl+vpF2egpxymhhJofrCP42miS4sHD
0EHUSdMD/16+jUkbA4ZYJfmSw0gGoOo0Vjh+JuvHdXZP1qJZmHBl8cbV+kJp3/rz
RlideVc5Vxvx0HtGSPtv4X3W6w77ks4aR6B8rpRKNJA1qr3WNrBSj6p6N+7q/cM9
pE84eutLqKWetNwOiV6XRnePYXhy+b2CjMLwwISfeMZ6nosp8/W5AEm3x4/psuhi
ei8puNo3/A+1unS/ES/vWInxHchEojCwm16lcVFubcOGS+RohEmbkhwZrvi7raHi
GFuQkoct4Osd+px/qGVMmgJp7bjA3qXSs3AX8UznzZlDOjgRKxOTyYXM/nNrEk9+
vOd6TeWFlGDcKy1pmsbdTQ9QDi/rpFzQKlQkiyyr3ess1at1yNIn3Q6RsItLRh5L
/d+NOGwLPvdkzFEHSjxpREr6n3SVlgxoNoUXUUhaHCYCnUpF/W+0ZXqAVPOEQV62
OyETTyz8jl/zHuEJk3WpCUaBNg86nI2pVXrqX7vmr9WsbUw//thoBhGjbAbbkpcU
AUOfVY/sEqMpOEiRq/QQZHX3uAmFBclqKFJSgg9Fh7oTmg1tX3kX6mMtA6X4HEDU
O2LiCuYnLLn8bfkRkQ0DBEMi7m85A0tw8oyiq5B2tYkTQnBmC2yHv51v0UyvoDGS
lexQzEOqSiZJitAvTWfLhDNqbqxuAprKivAG/moMnIrJxb8YMyfZBoicl+kkfUDR
MiGiyf9Zyr1gBVe+8IzTH0Lxb+DXy5hutXzPeORQ5/teKFbAnimD7E2h+Qa+ewOU
9I/J+zwXXu+Sibt+xy3DOMzEK4WW2+FR2vFXU8/cQhXSEtDKwVI9DVGKF5f1E0mt
XB66rHA5cPluMqsGFnN9lS8j9poYPzqjrJ+Z1R7ri8czWEolgt1JRvsCMN64SSdh
B7C4AevIO6r3X+kWzbyudMv2g3m2VzUQl8o5G1ZUyqpcxY3f9qILaUgrYU3+3rzb
aIHbg+RJWYmQZz3x6dAbl4WY7YL6rirM7zfmsun/YIIX6OyvYn0uAbpIdIfU5Y6l
O66AGaDxoGhSVpD/Iiuk97tFt9w5Pcz5s7QVgj4vGVwXsV86lsOvL9ou4ClfUZZz
+k+bOPJVmEC7FYPL/w2dgzIm/k4TghImYmne8QIEuNCWlYOMf/+n8LiyxP5Bnnek
k/fqwycHvTSnBEmYIJfxVYp0YZ0OJcTiZFDgVQP1gubEZTNP9Nh+O7B1DKC7MVjA
xaPn9lgCLwIJ9yHTgRqauVXVrOW+5P+/ouGKejMxb8kLZ5I/CXgp9nU1tRyhFHec
2Xln5I5K8vtpp58/PgAl9EDD/GnUzNZUVtzzuygys0lOLt4CtyXHfyWi6QYinacV
rFOZVuXH8b3H8emIIzYtpViZilJ+xlQZdA4jKy+bKCPYoL0PZrko0mrUCy9dGU62
PchpemblWikb1SsT1agoxyNxR593ORkIZv2g4DlIivf4JDHTWtGmpEiRHhU2EJ0n
7dVy2lOs6i1WRUHphgi3D9Z+n9ObYjjVeFf59/d/dcOd4WJST9uU2Btco3Em5kK+
pLx7FRl7xvszPQ0CSVooBkLB9+YWKGk9KtYoFqRrij3+fJxooV6Zt0y+BlLisn3f
z9qfCiCj80DAbjQYlfK3CexSINjqkCAqxPOu8rrKcxwM2AqGq8iD7Ipo8ryvgxFy
g0d+WBRSNIScIm2AxsTjMsU9w3SFfR/KL9VQYVnp4TsjX43nE5PVumaqtvgAmo7z
yS0P6GdVs3isWxohY8/Ayx6rNMPJPgqABM5rFEqCC2LlfosLsclUw7NgaL04pV2Z
FU9WmdXApUUGJlIspN0AvxJanwAG1rzjfiqP0TyIQ4XrxnXcVK4kt7u58WzWVnbo
oDQDuz6dyL5971k17H+px5bq/x6aMk+0KHXT1RfbIWn2o/5F+nB/RC5C+SgLAHfK
XeWhc80kEjDaRaBv/TN9MZh7Eq0x+1a6eleapN5NV8bgJZsPG1eBtZG62GEmwG4B
VyLTlsT9FneMczV/J703B73HCg4oej7+TLD0y6Am0ftmF4Kr2m4WQH2+9X4MDZhR
7STLvvPEtaslqeTOP3wUXuKKtuf6FF86XrYinN+q6dXePsDA1ES3NlvgpEu+qTsw
8xo5MdSIPAnILKbVJpOH1viFPhfzHaJQLzk/RxLLfGqXVdrty20u2Crt0roD6b38
am2hbTYy4bxwztNhocqN24uWSRAAnl319JAX/MN8NX7iqAzpPe5jrzqihNEt23TZ
tmUrsctQ0Jf1e+3oqpTi6OdYrriAi664kL2kpV9olOMOr4jkL9W7I/bNVZOhlwf7
tAhHuJsM7UxYkTEf8vAuIQd1xmTCXZAFz++eKiH9KoUiCx24ZTjFWIEStk3jM4/5
iXSIvkrrLi1F1XbTL5tGG439v/oZKOwcS7qnLLhdoRZdSL7x5vUqwWGEjC7PDxIP
JC5f2I2vRLMyQI4cS8RJUr2Ev785HthCPbvG5xB/wjVQWXpivWxK6KbGodSDfod0
LFxZ+QoovFPoOWZ13XJ/NsD1n5B6HcEVWbY29rc8okie3bzJxBAUOPzbcsu3kz2L
t7Cin9F4a6EqW/BZyGzsde+TpNXH+1lNn7mMHLM+llKr1oEODEQkkjifkHUTxmL3
ufKpDll5/zY4Ezd49tV0WvVBtVV7dOFeYgdO5lwDA96Urykr5NFB8nuM5KZM2Tur
sUpOJoz3wigiHE5d6MPc5SPM2Fa2qh54KOQuQ3zmOpXkPCgE4njWSRRP5tI4Tgar
kCCeWYD5kbAC190ucxXYJxuReTedFvU9hLhUz9WrgGif+ZddmAzMwWyZjJn48TTj
cz38AvvGDTQg7D5/ro5E6tuWf6rFAQ5RyaXSCi/97UR3RWTc+CGxx5y9fSLWCTBO
Qd8TM9Dx+5qC8R+1tWJQHdL8boQv9jlbu/30tR1Ll5kN/lE3bXLi27s1iua5Gyxs
InJggsgC2rmDQ6tl255BUamUNvJxWnxHdlta06wvdcODn9fLdhG/W1nYbEY/zeWu
sqwgNN/+8B1fzLXZqAmgVmF4IT7PYD3PPaQiLmIMy1Z0ovsTEFCWYPpf+sdXpDni
bQybf6QWXAG4uNnputnSvXDQnw1obMospNAZDDBPloQWaZX+QEx1DnwZN+0quMfv
L/TOvW2QAHu5G+5OKNpsgYC1JxXimUvFKDaouxvWxWm5EABOQ8tLtEN9XbufYm+I
tQWwTGx5GJzsckcDpAJ7cJ/iN0X0N7b0LLunnezntF1s9M9m/gMaQZiThpwiOrp0
qkU/gKuaPpKBEAye3BCZRVFKr0Z1oD9bvlVYxbtUYo4QNdsHNvY1A5TzG3rwGAPk
S9r/yO+j6uyCuiF5ONo46Msq7U1p73ZhdEz/trFpABhpZPDbah0eatOMwmWHidlW
/OTmH1hQn3aFoES9gZ5VHCcKVYxWjCzRfFQqZD/M8ivy0d7tbDijCcVTIub2CErj
beHrhIj7Ra2ajn2P/E645cXj3oE5BbEqEeby6J0+YMQEhJ8MJNsvH9tCqBdGRjoV
VZuxnbFwfJ8G/S/q8/k1gsgO6MbsdPQ5AnBl16b1ORdbiIlqGpbtiyuQAuqnTVt8
w+/laS2P0GLsKveHYFEdt/LOL84X/yXVexT6+mMfV1q9GzgvJfQfHFMEdZHIPtf+
N9SJYzaDmTdqVG6ENX0BE8CWFvD3tvRH8U9ZCw548VwKH3bVjakatq9pNhkW2F2l
E81C1vSnJn8E0gqaER//QutKAbBFW13BAjz3yBPlKgasU1/F22HX5nEmYOYgWE8y
TgEw+nyQHJ7+o7Dl/mZbA9l77chhKfPJkQ6Uo0YwxZ4XSb2cPqnfqaSbHCOGJG4t
cekuxlvWnFi6CxAdNEoHBEsub3+5XvYw0X/46iZEk/qQlZdIggxeREHqWO/D6qwY
YWTZ0zAm7SkBFSEWQ26ct7nEBiLxtdaRZO/G/qsGHrHZM8wvGIHv6D+vkmVFbAh5
+KBzIOrr0aofI2zICJZ+LSw2VhrUTSBEsjbEpNz3iQDSjZmShBQlvs+bx9GvX3vx
QJXGKvtSPH8R6I4f+/4Glz3WhCzvWMqhkAEZ+k5NIsT8l0vfRsGf80sEQYtpKCuq
7XqB/yUmCzby1r7Z4jjrYY0oh5TixrGfhSDyLQAvgnOKoj2KYBudeRE++AkQRbRa
99de6QpHlbW5hP6RCeKKlFJyZru+1ARYX7p2tua4dowQE3/1bQeU6vLkxLYZOPiL
hC9Q+qum3bpDeq5p69/qXLVwuVkYngVPwTjeHQBDzppT0fqtdoN9WtBFc8Cc64qK
vf1FuJRyse6b6bkhyasGAa/IjjIJOOBIBPkcWn4049kA8uHxnHTjiehS2aHulBca
+5PpjpiD+jMjZc8EUhiEFhfcnjCl6e0nXIzw9V3QSCPkLFHyxyM/fzuhPIb+99aJ
EpOYvy09SI+5cptBr69VJbxY40ADFzcnfw4/MIjBGJUtts3DCQ9uCXRk30v17qRI
pjAdFWLj1Pd3ZL92qAOFkLMEQ2t/LtyUIhilZkS+VLX7P4YHs5GGTj/slU8VHGjE
gQ2ix/g+1drs0vVoWi/SrryTZ4rGjiOgXQqE/9VQZOuQeoEBzip/zR9PzTH4uHzG
BW9GfJgYNfqBJyT35a3AtPyCQJ+Wjh12wVb6a2Rw4reY6eC8MHZCGJn6Yp+/x0dW
NBngSxWYfvrLz09Y10yWclRlUA2n5F7uZBotUV1DkMfgSqjna7oKbpuMhTx+f1TZ
j4M71DM/AJRk7uX6YS3bUBSEoWXR30NBMdFC2jntccZSK2RvIfTiGvEouFIl33hk
prBiBXLRB346mN0yseZAKHP++cinFW3yBF6uEd1ZLFHWRfPKs+oGNWZ1sC1RM5vc
a0ZD5HOOXb0yBCuXcI0D6wCBIgqq4/XLoJG1irhBMZrm483T1g2wV6TJJK6Cu1YM
OfIfkeLNx/aZbTmi19JoiEBA7Uqf1AFIXTQNxyuabzjXCVqYiNZ4Gf0jjyE4KE//
vmqUSzTKrewBPDkvrk3jN3iiDmcMsVlNYf/pOqVkRfuVazq0MCqlqslUa1IYPoCy
qhjVIZhA0oueZ3LeJppC7qb2L+0O2TAnntyxVyC6xRLh5GIZ7l87Jo5e+zcOuTwQ
TExnfGQfFz9VPNlNZiAEBITKb3EuiU6mhd8ArgbZVw2we1D88fac3vx9GxvSIYkM
T684DW8XP7C2hLt1lUhgtMICeLQXnlo9JzcYGXkRepjgu6VebL5M6+78G37XcW8T
n1dEJOT7ZnQcjWsSHHUp1hJfeKsJ2q4b7ZxH5xbQCIzkaEJ8q+pZGCaEQJwgN/k/
eeq1yTboHq8OY2YJ2GKzzlXYvb57DPtF9fKdBO6s6VzAgIYSmIozk0wDn6e0zZqh
CpWakvO8CYwFZZZMGU0I9kN76yg3aS3FkAXf0WqMnRWPLSGkmsvmmEwxLjk9kh/o
/n81RU1Ahnnmr0dvmBw2xH1X8dtIbI+DojpL1+JCFJMGy9nhobu4+gS1NxYFjkMp
C7Q+1vTeHsnYlqBm2K6osvMLD895wdWo/V/zkyPOElYBfho+w3KVqi9zbZoThw6J
LceKItuuzPF06J5AQnPLcNuhKiJ4Mx1Cc14L0LjUjYWoMvQ5HUVRXTqZGMeWMhlu
+MxgWswz1MxTy2/Nr2gFUM0WatU0FjpjTlsWE/r+d7e635M8bLTJcozev2G6/FMC
nSuIFoN+ogQEQ1Rfs8hHtXx9mdJnrpWV0BlC4H04UHNdsIpzyzYc4V2wEOT+kMwR
ICsSmKuyoptzbhv96cUtuEWUcpkZnWSOKL9RWde8M45F8g4ZRCGnYGclkbZs00sQ
cXYIdCRMe3rrS2I1l1SZhqxHeEl/VxNVBN3E/M55pQtMtipTklyx8/RbpoYQvRqn
vjV9XaEs8nh4JDK1PgZlmTcA82/12fLD5HObLVoJ83D9D8YI46of2/0zg4saIKNI
QwdUoNFXp3nBS/Dc7leXXXDaDYJPab9dDzez4sHzw7txnLBL0c8P4mhGVDtLCgRM
hwYTaAmJtItUF2NPnrjK4r7P8JkY5pf2ux9jH+OkvEvwDzw5ywsGZPckeUQxPIoB
wzafJ9H2/VtKWyUaXEF0JVAtd/TffTPhxTHgxGWENin/eFFPq+rm0eOKhki1Bm5w
plDvfOES4rFK+bCT7zzpBEVkwH9hp8xFdMuOqM+jWHVo9wU6yeJTZwuBo1o08piu
NnV7jhuI9YnvFUzd0l4/i3taFM00OLIhYvlg/F/Nju/VuAjFHwNYq/Lcz7sXhTbZ
khGmO+FqRIXHr54UNgZyDLZ12pwjGH9CuaqvHdKCFAawF1A186clBKkVade7S337
UW8YkNsGlMTp7YJNy/eqMasx/U/42wQ6GW2qlMxyAzVoW6H4eK6yCiRT9T4blaE8
ZuaHIKMEncSVCuQPuuompLBEa0r3VsiZreL1aXRLKN6JnLBsti4z1DTQQrkxZqAG
MyVda6UDgliMXkxc2TnOLbBa8nJriAfFAs6LBxguzDeIEceJChFztXV/J73CvicC
LHs5yW5HWwO9bgyO9RaBKur3f0Itm5enWobaccq8/zpwrTI+s8EI4Lo9OsO2CB0S
tFOik68V0Q2s/qBiI/fGNqyZw6KkDc8Kz6QasGmEdHF+LN7Px92v08vaT1p0N8qV
4ez+9FUxQSzgQQPxTuQmQ/4YIc1Xw9KSCwKVojU6r7yOJyEW16t9UQ73Zn7AkdEG
a94KS2VJ4nwaSLYXaGE3Gjje0QihnY1quWbt/CiYxxaXnlN1ZmhSDSwZEI0ZsZjZ
zAIyRyEiN3+PqCthB5hTizzTAJ5aPnmVtI/3thRvra4Y1R4PeGRVEyBulugqXKUa
MNnmg3ksTXj8KKAsQfPtTTBKRB1C7srzB4NxNYtXIGGgiO1ZN0tciIEfuHUUM96w
bMNDQR7yvA3QrGLl74EqBT6rnf+SFoOY8wayxZJC21S6U3K9bly/I9Qg+Oi+omDy
QvJQp3klgY8j2ry08YeJKrW48b0aNh2XW1CyxLdXeVBrhkweq69aSYgoJwYch8n/
jMoQlnQfb1hvNQ5vIOZTixDDN/YXwT10zU4IgnBd9o2h5mB7zF3ZqLsJNJMXR8A0
4UcXY6QYOhfE/F8uLnV/m1k9GHFNgUTOpxSpv1dBNLSE3nCoNVtJeu4fNyLtKtNM
eWkFvRB1DZdWcU5aDbgZsWG8Tm3i/6lnZrXozdM7u77XOcHRtWGkpSRecaueQ76W
1g4VDqnbaAif1B6HAyxcE0iLLCsgifE/XqfmbUo+wZulrKsqF5S33F/4HQvmJJyE
+ciBNtxj4LXgIPgtptmPbUopYEoMNs0+hNmKjnU85HJ29/rL0O9Undikx+UboLDA
4vg/mNFLsLgVbMfV7/iHwFWiFjvswixgY4XYCCsoZer08Tzf4FmuXP17wWmNZXs+
YkoErB17pV3uiKBvch1OwfTu+2W6n8UfeWQMJAObsiH7wnOIaABKpy2+zHb1PaP5
mrt8vO3LyyA2sD5/AyfhL9KEDcoicXQFm91EQFS/hTKDkZ+x0zcuJ87m9e7srQbZ
9HgERSOLEqj+7pQ+AWJUpgjJlGvnEncDhcPKSnO9AN/oviJUf1H/poTY5a7jWNTU
HRr1xW9YoikeL+hMsByGa9uyLEKisadEZIdvCRkKxXtidBvqG+Y+kumc7g6wtBe5
KogQR1+ebo+ftTLRO6HkqDbvwWvxtu1HdxHQboeM29bfZ2U0r/jbBAMvrZBAT+Vt
gP4/MVKc6oCPKSilSzUWYNyyvuBMSrfFL8OrSChd2YPM0Fu1DTCdnROebNklVnNm
zz2o00reHb2CKB7IpAPFcpbrqkPRgEd8T8bnD/5l0FapgKB0163aCRqnUTPEJV5j
rkinyc0Un5ERSWDCIGw2TNlWnhwnljmr3kWMRVRfQhk5k05nkEoEacMNu3IdcV+n
8Yrv71pYHMqDsPdoK9SQTcerymIZYJx6AqFRh3NIFBCSbrj5626fjAUh5VKT/0aW
AL4COHp0dUm3bBsi0etmKDQTsnLNoL3xyT9ntw57WJ0tHwYnWhmQWcf8dBQghGcp
sPVwUJIqODb0H/BMNHga0NbvCjRZxMKLt35Z8vmNfjOgbJ7etlWU7qsgIOJbAVUz
3n2ehXFxhVrVEvIYDEtO56U7/En9iBDSaYI1i55a7VMpKVLrNgpalZFD9kLEzUMN
B+HDHrLMhbsJ+zQAaNsFFisOaSkfj5IUknsrdOKjwKt3hhWC1UA/X1sPjaIUl0NX
agArcMK4j2eQnwssbVeXxNsOOP9HB+L+XRGiAo4AuQMbzg3QniUBL+lrt8pGn7H8
/AoK6LCovD1XmDCOs7B2CFPcupfs25a+LrRRukquT99Pn2OSt1z+QlOGA35qrHd9
SvUn01QwQJm/PvUTBHGsUSyhMw1dsz1wiAaHH6rTFb/nUghUbYdgznf/eIYyu6+E
hvaKxfpNUtRJ9aKJHn5/gHdz4xp7c5xA4tSJQ3SOpdGFe5yzfw+Nx2iGpfOggSjh
KhkuNlKP7CT0nqoTcOsXD48xCdnv0MN63FLXoST9Zvug1FLfb4JCdG2wVIk6Q5hW
c/eDZPx7RPTBpheLeFvGfESToziMQAOE/FWMuP7trF8OyLZL2WS8VM1rlyrbUUsI
kkpLfs4hg67THOBlvRMvkVpQKEDG6KPSTnCqDfXAR5qLL40RaaAxzs2NEqBXCylu
HX25NC9mtRPsg/KWCOw5PyR8RnuQuudKzekkgxi1A+43iSshUgtak+a5/2DJgmkX
CMLxnytFsvJTywDM/GpQudO2PCSyBxLG9ZHCxSFULpjoBEh1UaQd+Jc/E8XD+mpj
uMDgERSg7p/CS4vayh7/Jt3XlOFaOQuoYZukAdX5jVas6KwhCzhNiyy6XRfCfLxw
CgHVAiFbLuy4M5BjboM4lkU5xGmNoGviJZsyOj4GNEyc7hbSw1mOwwYHj2BuYGiM
qRT2pTlS1xsyUfLcdfMW4cW370H2+KPXFBQzTE1YtuJpSwt3XldZOBNU8U/0R+nR
qVDIc3/PRXPqi7ZkG6VJ7VWFgeRCXJoduiE/fycrSr34gY4j9uSJqSs+oE27DUzi
+1Bu2TZUuYbFDovJzuYEoDUquf0fHM3I+f9NtsgGXxCTV2+QgT61hDQN5pSPYb4u
lsGi7W0HqsUEzyxQgH1WF74H279A7ot2xhxGVe7IrgrRAvq0i8TSPNPImRqKcHmT
tspbiUpcce2c0ZbRTujCZTrsweOi/g1NYV13kQrIjYDv9mPEkvW1bZ8XbDeQ2bFX
hUXxbVBDojcdCe8FiSr1AI6qQ00Epy0lcYrxNcDuOEDprqSl/VYrp6AQI+aZ3k/F
U2iXEQQHY1bA1tSu64wdGWLwXxxk0GJZYDeJkBOYApctVKan0jcjMDAXkxKuDhhz
oB0fV4kI3kBFTHSxVei+CvngAeIb3LAJyBRCq9eA98vzZwXYG5cvvEgVczlLqAxh
vw7A8Zx3WW9EJuc+eGigQELnYXyGM+iOyeyNpaJNQ82lmWQedM1nlR4AbM8HzW4T
DM4JQsRsuX96tQ9/VmkQ/jqlF38f4e3OCG/pFdickg3RhFV/ftO/mfJbjLgi52i6
jgslH07wj9JnQGaBVhcsFwqA9x3+UCGgjvMTj6geJlOxLz/q0Ota8nSbqwbNR39K
VktN2X7rGCqgeThESsrEX9n5zX2FEPOaEeI8FSM7JO4oWE1XZVO3u/VKCM+/zpEq
Bl0RRxg1mFblSd9sx6TXOitjl1fR4Jps8uOwVxukshqVFIeY9BGqT20wVyCU2jwA
szmUaOTGs81xglYtIP4rPt/oNaLLftUW3X238YzFrGHEzVKb6GG3OTayWgrS+qzN
4S4n7j2qTktxjKU8uDUWzwkoZp26RxPF2i7OTeJgO0X+qjeeuUC+QFOMi4vwcAib
0cbe3Un241KygmgcPl9NGLsy9KW63PvFGWnbsubBZ9HJxMxsMqsbXv4Ad+2uK/Yw
MdcbiaZ5a/jOy6AubB2uWnDd0N4lw4umtIYf4P3a1Jfm6Wy7GzbnIoOTKnh+H9tR
PEpGhx9msPZvgG5nKqLjmQHkPm+fSu7qeOBw3HYtHbe+f0ikytM2pRevDOksU+0I
+yBdg4o8aXPpbmIN+5gORbByyAwGyAR4YRBxF1tXcdZoz6+6nyu3TurOnC02nFld
41/+o//95nsyuBfF/L07rLMry2r47CrAsCE06V+/e0tLV56qkh5b39C74w4r9Ftv
vQlVN2x6kfIOM4s6dDBnRMsemZ1zb+3Rnvu6nBTsx6C1ThwSxUuCKmHieP7DyyT/
CSDuMLH/EvTf8H8fAFXX7aqcpWwRys6Mw8wc5ZoI6d5s5P3YtRe1c3QXWbqHBn1x
HG7ecxrgRWEX8MvHWra1EX++4ouYvG3DAufTRCFWYRitHOzUeaXxvE5LGoqL5mT2
53B3eIyaN2BaeHxhaHtLCgjwBbxmzsBVhGRsYqGm6FGrPQCI46IVMRUICWPryjh9
axy+4SIP7S1FxtfqN5AKXPIigtg0+VVqo4q+iAeTbfoxZMKzRm1/AjXELA3sutas
rGpQGDve61aFZ9smeYFS0Yqn6UpNgLjEkpLSaklZcrexEwR7knNbVIT5KVqyYthZ
E/jkVpgn6Vpd7tC8CqCmLWBg5agRIXXcS5TCGdvlvwR2Sx+HVpucaCo8vh7sUNCL
ILEUA+seuMeG0K5Rn2N0IjaL+CG6nG2jzgG7hoel8xjgVogqwrV442iJ+K7VqgD5
rZTsCdOdhJ2VSbb/apvH3so2UfZS4tQMjbH/2XEAlFO220j1rqlfq4lMSjrEpj6D
LtUTBp+axsjA/QCLouCNK5I+2fjhN4V76lMsYGj92EsELMoKyYQN40f7v9s+Ak+R
f9kONN2m4RYM/pC6u9aeB2RXqPxEQJUPMe1FavmRc5j7+3KaMPnEW/Oymw7MsS7n
Ol6PwbU4FSqD5/lWENjWF4qx8yMgWY9GAvK92e4KntAxu0lEsqnPiHo/1PhpCsqb
F7QD4ZUYR7E1shvEJId+vDJygqTuRVJAFffjRe/aq+wj3HhgfUi7Hoax2npaj4c2
Fg+smfKyTampouW0dZ01y7lbsLweYQwhfI7oecT/0W40nnEjEljZaBfBMpqs063m
x1nYhe773Olxl84ixPoTnTMhCP9IvXx4ruP3ZPVSm5Qca4WEI9Nocw/fGksS17Y/
SgOzgKCvH0ENF3uAL9QphHvslZeZ4GssFtCzHRScxNNw/flqA9HQIpvSjN5HdKfh
BIJI8ZVlQbEwbWEHQCiR23lygwujrM8jNQ7eKYwowODk4c8P1bOd1Tr59LdrKG34
sJE+iOGwsXSgA3Zi9AT+tgHTdxyE0FoKckk7wOdjE7NSjKdbUZ35O7hqjZykJv9a
V9goGAFR1a0c6AFWq1vBMb+EScBGWzTuLBoxNDVGP7OP+VIREWTWp28MaP1V0GhE
0zxwGsby/civIys/5PFf6e9oYRo7sr//bS6StVIn0U7l4JwYlbJwSyinqRvSRsxX
770Iqg87H0ekdVVlNOZHrZ07yHKk50nFSwumKEDPbwPN2RLrjmB2QR+yPA4uqSQ5
BW+MouIhk9D7isOf2VdpJ0dVolt2eHAZBC9GUFDivCQYE/knMq4kwMAEZAYEXXVu
w2Ai7qH64KfYLJNr8D0jsqJPwT547pLnupWB9hOUDI/oPXh7aDb7jXSMm/iBYYh/
K9ffD6EdUqetqmul0/lSBm/cnv/kXD73nIxD2MdpBi7Haq922ceJtJYl7qGmk3zh
R1SaDuzWL0gQaYJnxlKunbE/o0mLyt0SKNgrqeLFf7etc8p8vaeaXx06pKs+BrMd
oRudo+Y00VELWAryEVXsUOBl6NqxDHGRCzE0bZCZXDTL77ZN0t2y8qwARC0BruQq
ih2oAH2igw8epQ3jId8XL8nhJeqC+/oBh6MZ0usEGntS77oFISFQKByiuJOtOXq2
sHrjMY3GdpJ17DEaHrmeh6AaIMhDtkbYicr6InMppgCaSqVyOEZ1Lj/UA4KDMy3D
EC7y8J0YhXb6Wz7ubd8UlVLSETlbyXsB4MrUdSUYUPM1YaYKQ2huqWP0lo5yVB9Y
K2F9NbbxAfxH91BoVq7d8USzNQolVLQuvtF1Pnh8JNRaOfbFhEsDNUKmQ3pJoIP7
R5WdastAqIiSUOiIIa53ej7q7DZ/o5paAfWyCfCNHj/SMEhWJ2+VxXlWfJUDXhLk
l19QaWm7qFAiEJ0vvooqxqKxXqiAWgYgwWKB2npSIx+uZHAgNHtA3McA9Zt4nBzM
A9Vuy8YK7qzLahlNVWuqOA9g2NyO5jmf3xs8Gqwat/NnLZdUh0y7X4HsX2l28ngQ
sym1+3mGqZwXiU+MXJoMPl++BkN5oeeTqzeGsYGosBkVeDWxt1WJXDUES+zRi5EL
eyHshqWAqJmORG/Xjv+wreeJF9ohmT+IxeZVrXMbY3WWUZpPg9OK7YnMyDHld+yx
6J2ybjM4jcHEgBLX23uv3pgeV4FxsLRLB+4vAKja/srwqZyDm2qYo1FWTGfSRkaJ
wwLcirOroofQbCSN3n4WAc1853FgWZeYsKYJ3OspeQmPjxJmLZaNcC6zr34rGFep
PyfMX6xHV0wiQaNU40kVzSxWAz94bAl1V/0eQbKsSF5o4CWCl6tg4DZwXD+aJLGL
4BEO2YeUfKpt2dA6DVpOdMRCS0FCRqwjJ7RnRhmgZ18Da00ZfguYfz73wt6Svbcn
HhrENt3eySMiwFfBYvquErd8L4oQjfRtTldSk41lFCvAT/CAl5vnE8QBh6Z5r97s
A+o0QcRbKYIdVkRsgtYIdeS4XOCq2HBRqN52Pt4e9A7Y0Bfa3UzJNi99/9AVbzC9
NgT7XK4+JhPARy4HgDBLQBS50QxdqAJLKKK+mz1ySl3+hcU7KfySb4njVfJKwHrf
OFQNO1swtgO0sma63nkqPZ2loQxqZu+d5C7NDHPM3kMyJMx6j6pbHhqQXNsTYJt8
1isWHaXiXcHaMwLbKHhOOyOOYbDFKPr4ALEes4NvY5XmRbYmzw0Ydy5ljXZl9clz
cAt6xJ8m1OjmoZO1ToCI9BUdxNaOg0VIYX8YQtHmRUgCUEb4dCR1WTUMPAr47ne6
VxBRy6RNkE66meEs1Vs2g7L8yyFFLL7OeDAr4OXth/OSyI2MRjCg6CIl90YTdndz
AjO+7yU/sTWwSegM3iqYy1dHuoOC8uWFkESxAL2b6tpjGIJLAwTxzK5pEyo359XB
1LbaRAqNTxVWzT/eWiSZ/L9HdZictsvDhixIEo2ShsIyQmvi8ZfLINzQgIAAWGBg
8J6UzBJwto7VPzX0VGvzwHa2wuwvMmIXWtoGuifFJmDUaH+AF0qpI+/A2OV4hXmq
YpWiRDyIKexJ/JfjoPRbXQbHJAMe1/KfX7HgJBWDtq+S/dG8bha3PrKN9oAFkFTZ
eWAzjMO+O8f2sv8r21JJwXiEjGj5hYyKmaR7JvCfBAebIXP2e+LSx/xnqjgPMy7T
ZN31m+sQi+5fCVwk1yvKZwLe27PcJWjUBvJ4uiESaV63AkT4DQAYMv0CV4SLuKHv
rv3g8th+PrvEeemtpsclE4ez6n9hcdSi66xNBS1ushj+stSFjgMHuEZfetjul1lq
axJL2WP/7SXY5oaduJtW3bjlkjsM7gVVXI+6FtxlKb4qcXIenH7J/sAqsD7F4tUJ
t1W9qEhQvC0EXl+Lusbd1YMHY9a113t5qeeQe3XhP23PL7XjJtPCxy9qLRot8ON4
Hzp4hYBEeq9YQ6kab+yGC8m4Jti4i6Hr/JZFJ3HNWzHa/a9TyPSOOapebY/OXBua
69/xWBRcXPxDlBVc+dphsfg+urUveNfVCuMfes8wUvpKVGMBXWfh9uzp/H3gkY5+
3lrS6zVRE8SkNDXBSjsn32Iyv8oGgZjyfAXvdwDO+mq8Ksbbvi2FogO1K7BsG7kI
q3+m49AQLcBE8+iDh3MhpxW+CA68Cs6U8FLr/hVpN70azYt6id8Wu23BIzzwpZuk
7h8hpTQvCeyL+xPGuWohh0rBYZTPlKKXqDusQFNbjiCLCmZF4SH5B6ZWPalAzSbm
vGQ0gFiGTSaMexxdQHRE/3oN8wFz+g0TAKFchpQAiRKTAOX93kIhpXZ2SmETjimF
vOIahr3CT6FSYZsGBvQs3kRxPjbnj3yLvv/rifnIvh/8RjG5AnkI9kBEkT7IdOmm
xJBiru67F3eWoEjEMRaA6mcEpbmyNjQNKSY5SeWpkC/1f4hLk7NOTL2vPeKLLZQL
g7pCWYP6efnwDenjNhRHd+563UmvWhFt8II0ji8055hErb+s3QjYc2On/tKV0JRt
htZVBATj5syXRNBlygRbJJY/9SD/cZyTcypWUsr1EEO/Mlu/ptVO5sQ+Td459StO
7xeK0qpmGRXd7LOVTMZS01yafuYKxfyanosmAJe3iWOXT6uDFgxwUUqJfb1zMe7K
90cxubk6N96mwwpRPMooT1YRvwY0IHM4IXeCmKFC4LEt+MVJ1AeugOFgduLJikxq
Tvv5bZpANUxlH9unkFHSpwrEvEmw4vb9iJ19oQYBKf7/t+6nv18IyBowSWU065ZT
lmoebgystxmGKmnXz2xUzNdrC4MwQIw0Dwn6TOYd6Du0vVa0CpizQdWgzbNJzPUE
Y06j6cBPZsNW3Du+3c+aMm9rqB8g4+FOy7eyKyC7f92nLcz9TtwDixDoMAhdufW8
d1rwwcXg2UgWAbH37b/VxchiEgscmv6rqOE2xkLBgR9RNAsx9vv/i/hoEdcf5t4D
ChcfnF/JT5/t9nbOsuPykD0wI2nLs95Bgs2nm/QgOGCDyrDmyne/REjq3ttKoeGt
5kEJ3UnZ46/boJHjFcI2YCoKUyLPI/URR4YEsT5zLqRLoJrfsYddko+7weM1Zkpz
emxOD5fKAOEDqJ6P8ThqrnMH7yJ3yfdR9kUer9ollrmzaFVYO3JQmanvB1McI8MR
Dj0wiyUEVd6cChmOpaWMVI21WEdSYjBhhuT8x/Fw0JjGuM2JfYEFPmk6gBdMtFTR
Oln2kvn1HULbZH9vRB2C9FzD9NZMaZ2K3Dzvjl8Dh3JhcVJUwCyk9A3fam+A02Fw
gQx4Awk5OZ56HWR+ovusE/uGDrwf2317q0G1gq1yxg82YmGFK9CH4InN9o+k42Pz
yPrwTuDuiYOhBo8Y2R2jicTP/6iBnPu73xGcqxgy/R0K/gtZQTE+5gaXAm8Fi4yj
72LtoPGDipzppDd3nAfXMY4VO+sJznpqtyYjc9xd+ExlOJo7Q80ptH48MdlM0+GM
JPAUxqoqZTv0GSqPAqPrx5t62lv+vRqfCXbACabePsiEvm9MbkH2LMGrT/la1YLE
O0Nh+EhTZIHFlT52usLKcVIrWStB77vLpKkO5jjIb7B69qlJp8FNFnWHqUNlOLpq
4w4tyo8AJQQ8hFsKNrKewctcrU/KA1r7nW9k/THLbkG1iKTmKnlOctRxRWsYHkee
TctS6eTM+3Jp610pSW2dlHTwqvM5So7EOu0SArArd6JTrhfLDDJ6fFeZaMoI9/Bk
pAZrak8UW1oTI1GV8C9I1lQ3+6ixc3vg3Dlw0ZrC6LMlJ4ldEgVl3CpCcQ96wITX
3/dL4izDLnUftgMqMCOtPxQ2dDO/JfHqyuaYQr69bnvj1d3f2C3+aV9/MC+qYjCP
bPRZ3QxRAJ0lKQyqDvnG3VfgBMzQe8+D0fYtYV/WUaKxS2VQXhWy1ECKusbI7Rdw
KQey4c7ex7AX1NISSe/MtoF5JX7bx9IqhJ2SVRjZqgeaPS7YIlxNg5kaUjZw+/r7
pJEbSW4xY82QFFhgem6CXuvPycGLzp1sUagRNNFbdz086RUfBjh1elY5AqKW9fe1
yNtPQmoWZ79tmqQc2jA6YYI0dywyDIdQdzxIonUNof3THXDpCvts92myKAtdw2aQ
P0S0OPu8gA6t4feFxRHCzD6jOMSMPlVE+Rg//KrB8piJ063CDNYlLQ6Sm+0X+LCz
oIWXSokXjxJIDTTD2rsA1PWCiVPmkjwed0xEBe/ddXixgyVScQLkVo1pljx/e6IC
tnKrWcOxbRuO8GksZv0+aMRIdfnRZR9vaJXWXD6KfMb7TpN1rlNiW1iG51Ax62Z+
7cTPi3uC+Rb6sISwet/l2eWLYC4G8f9YRl2HcDMMNmU5bRIR217X0+xVaXjgK2C8
EicRUQ32v4s8SwPLLNVK6zSRWKtrIo7HONORIGGQxt6Isj85JMvBagS3h0TeVBaZ
0XBSC7IcjZwk1jGcUf+v6f/G/llTqNC+ViqNcKEyoGhtJt3oIhil3iPiHi9RYIn9
Te5MhmAHLu0wl4OQT3mVGUkdEqt3pNv1XtG4843OfyXzoeSzXuoPGko4R2UQTz0z
DfB5mhIEwaROBF6CbcHUF8qSnTu6p2CDba+fyC7/JnnigrpvsAYBynwB3GKGVZqh
n3S/MD9I1X3JsvYC7s5Mt9iPYOv95moEesmcNjTMavCUCz39q5cwBaEnQdFaIuBy
BrzuRRDxhCpzttALUJqqn0x6vH/PHDaKa2aDPfo0wwt8KvSSaKoW88VycDbh6ZCE
kXl+Kni9ZVfLgA3yFGPpX43kkG1pmZEKaOD0cD6ai6/ANHvDnCkZHSmgvpA660le
CxaadlG1xg6TnzE64BRS0uToHzAXXNKbSHnDVJqw75ZK7TlaqIFn5sFIg0AsXJKm
6TXZrzsXaz77EQdRmWVyA8Dx2HXHpkylSo8luQlEu8KGh9qpinUpQ6KKNsudJEkK
JrxY1tpMxGgq2VSFvli5YfUrAyJkHAMw9T1ck9MZ9iJWZVaO4oKh4U2TYcRLIq9Q
FP19/UpRqjRp+WaY0NvV7ZKS9JyCdE3ozXHUVHd+t6+rEKUcCeJuPYwohe0pBfe/
hXATW4lAjKv+M7DHwFr90n0l0uQ9Jdlsib24OEKK7ezAkGC63mgNZmZ+x7GdJYnf
GNvm9CuVWwqDwvW1RT6bZQRT+/OczgwbUCLHncPy3JbCr98bQJDQpREhZMzQGige
Gce6B2UZu26Aj7XWtyJKy7G4km28bLMChnSWO5QEcA2isfQ2cxeUAt6PD8r1x0rJ
hqwcIEg+L+3zSDVg6jPwlulVdBVdKmi8XZSg3553F17BsbBpqoUa8Ib0PHZnOZUL
mpT3nf9H2gYXHaGqgjlkwrNANac+bSRZW5L1zB83CJpw52ItcRW/NAzWxzfAJYGt
2xcp186zZYPCYOSDCBFyxjld5nMJ9Oec36u61NE15BWJSNHmZfRwGPTtcWKSQGhK
yskl6on6DujicchU/+0t3lyhSDOTsb/N4/SfxvMxhJtuTPcSri3WAnbaKdVBtGKi
oSmAR7SnlienhukEf5ZmuOtZG89WLDihIA6SU5bgCRtUvDTnxStYe7hfF/WqXgUu
XXrsGOV4S4w7JZgD/UYTcP5wxF9baFzvPEe7wWfZtHUPzaazn3fa3x27fJ5tMVeQ
23Yq+8GXu/k1muZpa3JKkiOajLPuCVLrFpVMG0TCGXj1H4mJ53rCZqTVxpyQ19zR
ZuLCqtfffxdVRsfpi14ydQ44zB96VqysgLvp/vtyAStk5MkQyA6jSmoLUK/mUcjD
PsiLJSc7+XWj7XxfEQRsiywSnCTkZmnkwSwtOXW76TYzpCa1l52/V5bnE0TK24RL
GEvw9qRPH8q9LbD6dVmzEmb7xVvRieQEO2iovbf0C47C/kF5FsKmyjJNl9yv81ch
9x8DubBqJTLlHfKYO47RkY96VmDk6ebA9IUx3aROguiY/UgfViVHnjbR/fSVKi6J
i4Y1tgR7D79EsejGceXq934elFCSfgeVqpdtjb5CyYoUFNKisGi0dN087M9MliSU
djEC1q6LONlE846cr7zj3XbSktiyzhWTAqnOdtt+w+dLTvpBbPWobv9CX8tiCKQw
mNy4egJkQYu4hNYuB/1ahrLjTIfkbmQRAFT+4Kq7UT79vIuaUPloCdOcfEJsDT9Q
MP2FggJ5Z4GgmF2uqCXg6qusKfnLOhF9wCVbePHFDbhjLPyUR79d8ZjINz+js1Wt
V5ENJAn3HVt34tKFTepuH5ApmXdJRY8BIO1GeO5h0VUY9ABonydQxkA5Tb3tl24H
TCxYBwMS3WAK3mMC4yZosN+nY98P6gy3TAk9leeEy8y3b53riAIkC2AqBTvIRQhm
7oeKUAlZKLnkFKA9Wi1z1VdGawPD3qfE5Qhu3jym7KzCXXnop0JmtxF8daZ6uFCu
6QOphDGCdkmR73Cg56HEd8CVErt8GMS8pCPBDGc4hHxUn3iFms2xShVy9MQCrxeZ
KQVTe3dPgDyrgQIQ6Iud41I7BOiCqKMoIwJn/zwnsyIKWYVQCSZktos/rgMv/C+e
ufgD9M24owKjbA/eKp/mJ0gJ3smr8FfxfoQBezyg5Qm7YajRMsba8ES1HO1yr2xh
4cEheFhBZAaKE8A38GVE/OV7MIRzFL4lLStGh7YnDwM8rvlfqPlXTCDrqj1okTHM
cYuh4l3z+KO4k7UY3UOTFNKzzfILkQcp5pbrPMlGxAMcXg4BzHVmDbo4Lvc/oCDp
HS1LsB6EBMIudvGEeir0gVdCeIr38HbmEKS5CNEK8F99V/1Z3MMN+InKw997SejQ
rEvTnJbT4BfwmJlq/K7cuwmbEx0/TNH6MMPfLhi9wuSopd/aol5ELl2b+ev+egaS
dIAwEkr2lfMr51/6Z55BX9ilDEpM8d96CDZszMBsYftjrLp+RSLmMwG7PWrstmou
4KuUhfpFyfYIJ/NxZ7dIzXcJ5VN0wyYEcaaTtEyoeh/HcSadOcI6xSGBi0CeVKr3
DMRfA03iGHXfq0dngRclm4mFOnYFZ0QMfFtj6NxAwTEKbqO7zjPq89CKX5kwmaYD
lzrlUBkkOktW5pmz6MTrcMl38q8xFK/XxbqyQfMkPaEAD6XWCMLALntWXHu0892v
DwugbSPfsZKF35u6SNc5iN4XnURzdgt+XmpCbB/GRe6OI9WRAAe7iMCrZi4GH4vS
8VwldVs5FSnnzSBdSIDS1W7SAU9yHYS4kcuyY150FDx9NCTR69mobC7EP0enkLab
eaiObjNEQy057XOT4Kommp+soBFxqB6982tLiwbcJ1QcY9A/HQs/gbJvpAAMp4Ji
pvzjBbGbAjSztX6huAKYSvdA/3HG0tFrIZrbIv5Q14R/rW8j6YhmP6jSSglzHaKY
/yNbHCwXYNfmapyb5yZXCWjQlWErRVKjzlx6BOGDhqHJaEFGQYHAot4bLKwR1hVK
TfXum19DhGgEY8dWdPdsgvKjDg2BgxXOhDJ3ffxRCok+/dIqKym9DitmuVHUKvds
P6Aj/bgu4LnkGEARgG73DRbWWopo60lu6YkSLOqmBLdq9e6menJBuW1oUYge7lW8
lptwrrUHLGSdbHBOPFUpn+x12UH+Oi+ooVle4x7d9qu+zf4OkE5VVkCY1F7jVgP6
A+tYIhcQhh4AOCIz8PaRFhmueJl/o3d/96Bm1Yc0CAaoW4uSxOO25rCCRLndt0AP
fQcBHQlp9z2xDqzAYaXmb21S9BtsaiaaHkPUZC+Rco0MHR/WxI0okKJO7ihDB+IM
dz5zagbAgTWmgbQcMeodeMNawF4bWXgv2hOzCMlX60wSGe2NIfRSx9cPN7Fox5eM
3hE18SmqTA40TAtdHWXpET0xzizTCnV+I6CeLz1MYSxahy8mC9/EiyE8m0yB6b9b
Ywc15FimMGK2iKPA3usnm2DeGyMkAQCoVhSXnPJvLUnhDVh4dR/qNodJdVNG8uht
HtObAwargalbytp2GFF324UlffoQfSTjgpYuxu2FDEa6wAFYy5Xjl4r2ivfEEdA5
SgM8giHJcVU3nsVim1Rg/cnoquzF+8oQAlQivreLCWh0mK5ljqrFYnCod3kI+0K6
eZmd4T4NLhFPMubDoH8crBSlI+J0ngkEmSA70CRLBqjfOPoVpwkdBqHJtMo90eUK
hRqksamL/HoNQnE8Z7fw4wrQkEqJ8mqiw8BG+sIS8LYAaRVIR/UgxPXhLMKGmyL7
Icpmr4KqGwMnam9R/FehjqCRFz8/BMsN/jeNSYZ57w5ZDv5qXhim7qm8eAcRRfCB
5Zi2+GU2IygDyuMKvpAXN2D1LUITX2SNN84B8075uGhhkWenBaBT8FDk/sHgOG+3
bjjBdx21cXPtgGSl5Oyr51lYNnnj5GMVnJNNg+qxkHqoEDdAdHxtPMs+qMhYJCcK
yR+N2R+wRaOBfymeWPLokWps5zUSAwacsw0rkzbYv5q/HOXoWwwwYPherzYW4ftc
eKaKIguP6YTCbLOc/fjEwolL0hP7Ru+2ybDdRpf5LK1JOJzuFPJqfd9FiFYVuuRI
3i/LmGjUoXHx3GEA4aZrttBhzwIfh6IkM6u7s5chtNlk8ReEo5NwbhH5eaT/y7FM
5t04Rp6HeFc2/D1pkAg24reaMetBC2vjV89kZ/FXo1TrltxUKQgOqR0QvQvQeWm7
CNknqCvNQYKbv+l+sV4j8wFNuQi5vSpDVfF/ZT3QFlg2lnIgNib3TLszPfSnDl1s
Psm282VjBrxruf8isbRqdKjPhvUfNNsASNF+9TrZWOfKjgofiMhiCElJMrWM7Khb
z7QMSZ7nTLUJoTPeUQltxwUwk6Rab9VNA+T8O2ERaOP45cErvXGksSDNDQhM/D/Y
om6oyOmh9IH4fs/BrHMpckXl5EbGy4++6ZjoSQPPZXNK/Q4Jwt93V+J25CaGnTJ4
vDdzcgPvorevxFFwhSkVhemygi/naYxPlTEFjmMKJm4Ij4wfMKt5SMzMoOsp+KV7
u7TRPEVjhNbxppxC2RzUBY0Ycpui7c1qir/2L0ewLd5mS8+pdiBOAIhbMw35ohPq
2W7rAysXuPyeEeZNLt6sddZ4tVWyPJS6DWNQhiOqVpjR4HbhwN9hjvGRLNQzU7dY
lTpnkxbZzS+qz501t226dl1P2POwA7q0sI1GC5wDW1awhiE5726YmnjMDA9Lc8vw
PMinqI73bGiwa9nxfCL4IypYKQlWrzYzbV1/l6bJFZ72S2liNSPNgcy7P2SkLHsI
pO9//1o7y6UihlNN5lwaPsKB/2tFx1l6jb/Vi5Ii0uJKjtOwnjFjIJDIwAzEw59G
FFxFxvrouhJ6CSygbVu+TA4AzxgeW6vlgaxcxATfavhpnSCXKfyG2OjTqdy7PvjO
85ptE7z+eAcJDqIz//GWLpJ+CUwMFZRbBa0CcJAO/JDfL4zZ3dXCkOFZ9pVz19MX
Y4ra5UKS6HNHkDBnc8U8yxE7KRWdC+irM3adbb/HxDY7y8hu9js0Af3ZHtttlUKP
2peezZArpjkp3wDFLSfBEQCQMj7CbU3JmkHQfpbYKPYzMZMtLkBviFitNqtxRIQ1
9kcVV92ojMNxx7dAAUOoR5UQK+gwCLk8sfh/Z7iRIkWmcWnxAksSYwN+pU0Lk3Qc
PlhNkG4SMa4ERIcLIcKJ7DNOVNrZDPvT0a4Njt9Lb0YqQFartWU9Iy3RHHValnNB
711HQHhpfdFyn8j6ubIqWRn8Jp65hsNEBBUJDNAeFi2a/HDEKTGjDgOq3GNViCBH
ObWoVi2SEyN7VXGqSkk4s+NgbnWKEDVZvTK30M1ip7bJHfJ//O+vcpFrD1RzQbWY
Dn/EkgFeirgLXRsUUdtDu/AJjegqPWsJ88/VjavksulAEMLwkCPv4cODuNDqCvGa
78JVN0+lvh8HyTgYqzzVm+xAiWVFyDDFdBDtIedNMDNDRK8i0uJd8O/6WDFoTBWd
wgKL0VXhuyPhvYQTM6TfiD3a9gNwpw7w8pRy90KBccrEsLyfRMu7YSmd7mLCkk9r
Rny0DFikImuITLN5bbFnuM4d4jF/XyjbpJwpFQyJeM+oIWx32V6qSdhlxy27AY/1
rWkQ8ynyMdJ1xh9CvMwwM9Yv4rfhuBWE8D4ecuoiMy36QuHa11y33rXFB3cYUDo5
/V4vJswIa2xLb7jzZfPpEW+dP03feg3YCqRS/CMlUsSI+JFwDkC4kl+kpAp/Whcw
cBP2XDsrT+FUa0fAeG5Vx7qKSCLsH0L0w8ZhLYSnqYVp4zHartXv295FtpsPJh4q
VGr1vrEs8Vias9ZcEg77ptNnOquypM9eQ228+zXZIGdK1pSK4IBM9unntzXTAqdn
1NGr1iiOF4E8ZYjCkUF4xL8ZDicvt5k1eW8++iu+8DWOaCaob20KC499SCdbrfC4
S++zIFvIOxKhCy1NmaKVEK866T/FRfYuR/7GEQhcsmU/heNiH/VUZDg2DFP67Hnw
4q1S7EM3y6MHPFXz2KlC2zUfiNJDQWwpVY2+O2H40jtKx72q1cLuWWsN4VNHAaF3
jnSdvpnKkyL0xn4wDxj8sH41QlDIPtdCHzOQ/WLycY5XaaJrbfQsbwfFAaw2mCEb
PxXAZDkA3DaRZmkJGPXa4KCkz6Ccc/UWcvrAJMsj5DVnb7t2pIplm4iIv2wyc/y3
29m22C9gf8i79dRk2xLJn7Fd2tLUITYHVs7ecr98rQR9d0KoDPlJ4djSJWs0Q7w2
x3Fs6+VQv7GR5qKDOpG2zM3qRQK2BCelje1D0kpVQD6PxySjcjg1PpxuuqHljYYk
Wy4K7md3dOig0FHgO2vPWUF1LHHOwAZn8W5P6kBmsBh8/gWmY+q/7g0E93gkvTla
J5cLbXoe5chLU/vG7eIyYSp5V4u651/lL+MYzble8xYklcWyvG5Kvk23FPUSWWjr
EygHnBiOOXmF2Ugq5i0F33mQmaGH/y5Y5uLAWRDuLw0=
`protect END_PROTECTED
