`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YK9TVklY7+3Oeu6wiTGBawiEx2ILJZ2/6jy3OptxIh/OzdDzI1LMHqFQSBUPQ44z
eVOapOhHbGl2pTp+bc/8DG3vPa9CzOwcIydg/J1kU5ZgnFowAdEDn3VpQMHiBET3
oFbUOp/w1C5V55DVWXfcl4Ohj6YmQMB2/nipLgpo61tYoyRs6v1PPbtnMYekhd+A
KTE37vqKeBZaOXR1cup+MT8UEQUM0BfWguF5AZGo9tH9/G5rhEEBi6oLWLLZdBBG
y067NvSMhckNc+Km8xiosjgMqvjBZ3rVB1uSeFCpAr2+Bd/+PbgNqqCJ8rNjkob2
qEYdLwbzlz4Tz2mMvLJG4H0/kaE7Bkju2PHNOzPBMmJ7nYsJhjvP446aof4ld8v2
iLPODvP7/gP8DP0czg/FlMkvLsditmH+98bKtUGPOCY5J6OfNnDItlF3Gy6QdLLR
6gy/KdxFmXvE2KCLx7KcFfWKgp0r4fSFDBWBBMwyftGChvsA4H4IsrKY8lQEOmU1
D+TyCq1meBMqT8GHt2lhsqd4L6/XjFymzl5Pd35ChWx+XrSoTZjiPyLd8Q61YjsB
KQQBCE/yJkRCm4H4c28NKq7BVZBxVnZk5xlI4eDSbjiHvAGR7u964hQQWPlhtzoV
YTBs/TtQ/pT+LHPznCA3GlJiB457QmoD7aiVLlLAgWTBw+pIJcaqyXPlPKFoI2Ij
rwcKraYUtwlmMjm/CzxepE7V6e/y489neYG0M/mAx9X7TCT2ljjWe8foY46WXOWn
b7QgUCLTZdVnU99W625BWSsklwrQB3X8Rjkowwm28Kxmcwfz9kYkPr3IaXVuFbkl
IgpczKyrPq6J799l8YcQTkcYOnBZ+WDtNcASnbdmQ0A/ZB0pQWzGTz00nO0nn5Tb
p3UOLmiYXzHZQsze4fXNSUsTvITv4zO3j7C8EKOCqzPFcQ6Z5A/7bCXPKbIproni
C0skTx3hyeGr/NVhLvKeHok1m48LKnLZZ3n2qcvN/tFqUfixMOeEj1MecnbFdP+p
29Lfy6ASJrqPsLhG3hGfsvu7C6QU2s0jAvDU9et08gfphnF7jrcZrLMMruMcx8Zg
AzTma9nufuQwDEgVUWgqmqCbTft4nJbX6Ci0zPbWMl7hq6zs116duPaYzdyYal0+
kWScGuz0/TFMQshJa0aUnde8vc0TbC+tu1AAtV4WuNfaE/NlOq9rFE9juUDtyen0
Lripl+OLQC6NngNP1qLQ/I2nNLlBYsJeKWUgtDa06VI2f3+IDvM6USDih4Cu4dZy
kOJyavSi8ZTaWYxMOcotnh1gosPrWkq6rvuTSmNzCxnfLWkMOqrNZzNa+MNpV52J
Dh6D54oB8+22Kwak9n5IB0OTV2aWVaZ+9mdiNCFaX3hVOIVHlB506cYws2ectpRZ
/EkKZueURkEXM1QI2Yoa8b8nJ8AZajqDtywT5fdObECXHE/cHy76rAZpKkx7y/vM
U12pVF+R1vJCC9+QLrc2sN891Ct7kcSgv8XmNuwOhV8xKixouTYbHQxLO9A00ZxZ
vgqsVr4/VyTXMNKSmFvd4sa0snIUCMv/gHj70TdzGKRcQXv8I2SLpktvEprN50l6
N6+YvPpQgWMjhaxNGJUynkDLscgpWmM5qOMYgGwiWjcSZRS/rrXRQpF+cHp77xoH
tFP+nCuFRx0Ntq18yatNotLK7B4oyyFQfQxEZQ2KYE8apP0u3IpvjqwPvnQJmrrV
Ewg/C1G0rcGm2HtItFgvK6hieOHIFksgqcEX12mQLYpKjuK9NwPZvRj6F72UfGLv
H/f9LntEzYgn06YGOG9TVauOg9QqG8k6xumwrFHI+YYNVo7Nkz03kl2HmpqONzcS
B47iLo86jjCnB+lW/4sTlO9/mg9LGthUrI2be0XwqbwogHMLp3Z7h4+i5Wmuab/N
InfZ+M9T2YiIAspph5v/CKonN8TSOMMJae+D21idBd4Xv58w2e0iYTyRB/1/NkYd
uyPsc6WCbP/a8QnYp3RHVaFBSsjnc1X9QHz9ZY3Yo2EBnbt1iTdrh4EXb0W+XYJQ
DQ1rXA5eAP8Our0/kQZ+/dkBOzsDVd5SHg1AZmrm6CtUyC8OwMGY8dG9NiIBgJmb
Bl/A2EkVWYQ+LHq+dKvEuprZ7he/XtXxySzNHJnewpiw38qnI5l0vMIWu1xNKVKn
FqZJaeoTvymh5GfADXe1HA/S68eIWccfQEPb8oBiikM85CMD8ItHaz4rpPha+INT
nYlnkmA2eHhrHL5UG/ADqn8hUWgxSiKeLNSqiXVlRqjaCERGtt3fi7XNKIcTX8a2
pfxVKsYSnIHzRMmcGSwrlxFHcHR6cSZObAtZY04WdYJYdvqepDKK2GprE9rt3de/
zuBfXKWF0G9dzJkyCsbXwpVIaxwNkBQi8yv2ezjIfc/2iaAffA0JYDpRNIEgFEA2
6CfCTBuOFfWRsQuVFR0N/Zm7HmqtclogEsNij6zGt/4TDY4H11wMn1lGQkOJq+TE
XTjQ//tRnI+jIsLgUrpPNqD5U9+VPq0IBj10P1aU1jmINYELc6BmB0P4MP/Z6Bip
Lhaoh2AMN8v7xYrYtvxu0lm2adS7/7NL+y90xicqLTXCXW8AgRpH652LASXTGxcn
wDMYzlKo2Z/keFm7klu2w+Vt/FKLkfUdQhBGqY6aXUzTSq2OaldEisdchYwy4jd4
QMyWRGrW9vYIwRfkEcib5izY5kj+e21JL6UCbW6nx23miNKwrlA8b6cz+ortn9yK
oZLFmfZVRXQDfr+6yFvo1pM3pCtjDHV7/nc2oOIUZFdPDncYvJ4lKYKw54VW/7dq
TWtj8oCgQPkHKncRtzFrHy1LjK74VqABuqG59NMZDtANETVyNnz3ao8b+ugL1sPD
7iIilZU5NUUa1Adyk3GlhLcfcfVbZ5F5+k2baNkpLF/qg+UsLjBsRzNhFAOs6WTv
43d5SCGQU/3xSqF9A58Ft4NJQKXmVs5duo9JYKrY8QcqM9L/rl7Rv5D/vR8MbwWR
7/Z90gNWZOt+bUqCygZUL/6NBxJ8DbBQiEkNqWZlEcyjdDGe3Jn+7+yjYiFJhFbB
H8IAf9hjyRhHRi46caSvv/Rp07PSRYKa+QARa08Cqf1DABZg7PcsE3DI1xZ4NYIn
vaobHIYaT38BXqFQFb9Wmdq2nQjIiKNLdgeHbjpGDH4pRUAwvm4Q3VswLadr8zDt
`protect END_PROTECTED
