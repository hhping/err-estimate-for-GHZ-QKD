`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T5g6YS0f7nrOjjuJm83v2xKRTtbsk3NvMqfPEz1nxGcoZaYQY57jOs8LYVytLdH3
/LzUeLd/+98oIvFIpashGtNezTxsdcYBAhvhjq24Grry5FDkK8j6XrW7ELfIQUa9
DdoxWBov5XGl3aptbLl/nwXkojqCBDBlsXmwA5KB2y+UQ2uK9XqI1/pJsOrEiTUy
chUUmYznhEga1TPvukM/ksiQ+QG34Rg7ugTMmOSPFqLvByGNpFysOPTw7AYjNWuo
SacxufH50lm+IEBj43oS5ccfKkBKoQY3XErLRPc/qoTmMeulaJhz97F7cUj6G6zc
kR+NLQDmXzPEthbeYAug7VmmRs9xZu77rQ80YWH9e9WQGRqE4r+BczvXTgiEPD2l
3tojiAwBbf3gmOL5nem7vY8UpYNPOkonnejj9bc0KgSa3xE54/rAV5WFirt6Ylpq
1IJnpTZoL9refRx1oilmnUEyF7fQrSo+SQK+1B6CLdvFHL8XyAWddxEU1amG0hjn
My6v0mxJ/bmHrbiIxZkdeOs5fbeU6Vcn4tpqB0Fw5a/tbe23VEOZyBiGXN2ZvTSy
EzJsxvQcTh74kato/P6zGiCvyTwcPJNRs7U9FqBZdN+oLLztwUC+ii9WTo/GSe34
13X4r2HKRx7pc2L8g/pQFX0/aG33ZN0I11Mle+Ex3xxaGalMyvm1eGOcVUexGK/o
QtHxdjdnGFU00RKwAI+O9w==
`protect END_PROTECTED
