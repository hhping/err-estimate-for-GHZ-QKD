`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KweM4Bp351XF1g1ZkR06d+Hme0EpBwCQhzPcCV506DX2XzkEyOZiaKn1wDtxqaJ1
b6NqUu+NOs+WM50QnIcFLoYmOQw1yrg92StxqN/T9wNt4/bculh3RM4vQFloFlIB
h1ylsJiKrlP22WuTivnSLOGjTZFfNMsDn5BO6Z9MPorE/RSXRnD6FYJkvBPuuvkQ
sefHABoNDYJycsYuQw8H3BRYqYtfAexJeaOP/t0SH9yGEhsvzdgOrtramS8ciocY
P0GPNlN5YGnnqMK2L4VcigLrTkbtrejXGV+jhyEzN1kxZAjFvin38v29K5EiFfKY
MYFhBV0LJcgPFwxqkKhnUeESLCsovXptzpl5J4k4lDE7Sbm/BgFab1ABgCyIJg21
5QqOTHe9u6jCqm4hltI62YW/KXEtRvDu5cc3Mj2QrWJV4Fq2jARrBi5OAMcZ2fOm
OP1SZrYg8/L4U6t0tPM4bsdfzz9j3Vb+v8q+yTvXtLTU5QyVR7CA/KQl0G78KgiW
3evhBjoDsUqGpuAl6gnGd0Gmhw5ImkO3VRjlkHSx5Gf/QFvWzI+IVKh2QtrY4Vd2
1vY1d6V3ra1wmqIoiOYnJvpZSK7XXx2u+68jlrpv5SlIWN+uzx0i02EyDFQL74/Q
XAvdeRFmXcmRLk7tYolO7wKGqHfgj6ltw8K2ew5yXWqZF2Xr8hN1NEKdEK4zzWWI
vtFkIZJ+OrNByxoX00nlBpqnKreQvCVDYFwKtlguhtAhWYYfuNgowzrF9juah2nq
6bpjeiDEy3K8/gjaTUD3WM8YzE9nGLVCSczzW4i4Dsq9f4w5fRPIE6sgbDXhB/lY
IU4Go6gwbTTFUfgg4d6A9RRC4XdNMn9iuAAilwtL5IzdxTFs5D6oen+ya3e0oJvX
8w4NjT/925dG3q2X0qJDbKW3Ij4AVLBKCe+SO0xm5JhJ+DPzp2s3D9yPorNptZs/
w4vl2hUIqO+YjgJoeiODUo0tqx8SheU/wEYuO04wVTTkTwgU8Dnw7LlHZTsyusZP
CKDHXerVbDLxYQ9LfvalP2lqanC0a+7l3h7auBQztswVnsQxgkh7Of4cp8FUTOfE
9Yv8iC0glGWQgAG1sldcZ37MkdqvAGoVD9jqUvjymlPZBpcb9ZXBnb+J5SATP/yX
91Ju+JBUWIyVHbZqrltbKDJVl5mpo7JZsLrcyPl8wheM4Ks4LRS9gxSfDGTU2gvP
DLUXXr49LefnamqwYtgR6nANDFNxyjCU1FG5t8fUE3CkAxGIQhFkJfP9Hp3anzNv
aIOj1NrI3dfT6dF+eIJ5XO0aIOdyI98mBjdcpVMiwgKtnuLz/1PcY7u5faUib1Nr
/maYRPfQgH4mEUbD9L/LpR23SLdHdORnSMg+kuK966ZtpnJyubExhnC702ZXACT6
H1bVoRowKkNzO7EOxQP8yCwqlmNuqzv6OFnjYzDTUoN0bGjMOaaRn95vi1cUPSGH
3+JXI/SAcqXuzH0wGLZzz6F/G0zGBoKcxLRDct5hB9MFKKALyiuaRZLkWLGA5zla
NIt3iATVUHNGOAjDDUOdqISGnxFz8/SAgfEXijFgL6qkF8KKb95Iye4ai0JibVkP
jaUUI421F5Kowa+eYjoIndOAvx5ivmO0X4pMNUqQA/wVm+hwDKQI9NBnc21GvamR
ixTirVROfbqDinoicFCpIO752dfr+4E34Dfp2MpqGwyuJoIbNCmaUNg1C0aQgiZx
fWYYDtFS8FFoydQ8HlTGKS9dfgBG4e82lCutSJARnKQXh+hUdl7kR3qhgFrC4wqu
1n0hF+vsaCGVBxSSzgofQKlWJsvm98tkrVyRe9M8UYhMoDwXlkeMgo1nyFtYW47u
89AhQAMnfmayzk1S68+OGH6POqJj2fK/ZtgbAdCRbJYyEgfQuIV6qfxmqvVjqaIy
cMaZYu55W38yUEQgIXGyV1mJe1Km1NJlb4a+Ey8AcKYVxsemFbHQ1yWeM0BkMCcY
FvPQQ/6kFODtdVdoN9aT/WyIb5O2QJAETb4Ie8zELUsh+gMxxuge+8LIy+zzUogE
NsiR66TQ6R4fUTN09HI39RhN2j3xpthzukqcZhi7AFt3M5WHOuTyp5RsKqQmMdCC
Aw0fRRR89kUdb4RnFRgM+utTdtszVEGyR3e2vHsf5tb92RnOLCSBTt0ZxR2844AQ
/v9g9tP/rLt/xTg/3XK5NO97H4q0XCUQhKBcxQlOgcNfTU3Zah6l+8dFS6tFlD8Y
YmCW4BFtGtvBXKl8r8Ype4qONrjD/hKTklWSls4olW5fpoJ/fiBB3zgI5tufGnMg
sA52OEEyEBQpPi37AX1CL+N+wuWXFVz4Qg4QSGAWCTZpLMWFB3Cor59VamRIUGRA
NLLjRmnbmBjZg+334K6rFhvn+bKXW0F/wWGk5QKXPbwk1GZgKZuBrfpfYPYMzBod
WHVHUfABztZYKv5bRE/3jVxHZ1E5PRRSySeGHUdc4i0=
`protect END_PROTECTED
