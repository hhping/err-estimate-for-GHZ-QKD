`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Jd7b0PkXqK/zJoEZz8bo+GJIRs01/YydOTmUnSQO64YtnKaqc70CX3x+WpmJfGg
exDJZBRxmDYeBQTcTr+DyJQBtsRMEwH9LqtNuP5kqGi5k1eNWx/kkFaIJWxJt391
TyVMDzx0IHykya09cAEwLZDj8cfAPpy0tCFNw3MyAdvfKuajbabM2dRihY5DJFwf
qPAzooI+b3337Yjg799Q1YSrgMAWZzUrB1k6N4LWU03H/0yRv/hjw10/OfmCdNTQ
UjmwsGQtJE7OQ/zBiLnvEugAUmokLxM+seXHtA6JSAIQms7zwxh5NU88PxKjoYUG
ev7Kt7w3kRXkAfwQBHmf2KzIdYxGw8PwsZ7+dCVTuSbydAWXxFASAYE/5tohpjLO
vUBLGngGe6mXFJGUQs6km2ZnSMvfPB2TDFECNGLNEHo43FgabJ7vsR89GdrAd23t
EGz9o7MQ/zB1pU/EQ2ViVKdLkCMEyb94qImQ1XjYIMCDM4ZDzJKWS426vPY6wWau
HJ2bn90OnyvQIIxhciB2RMh0TLJGIcYiCjTYo2KpqCLd2c279mExRBMbkiuVw5ku
fonzdHZ/0LuVDhzMErGg+V271/UyWZHzCPT/o2Gwd2tnA017B+4wnIl3wZQrJEq2
Tpa3HVGiyJ+q4JHe+y4ngy1sMkiQExiXapIIy+6iX4+jRNPd0OyJKFLFGmtN8Xo3
9i3ws5ZTct/6pjRGQrGiIlZJkD4B3S7icMGfRucsJLy0LPDTRGnN1quxXkUus3B7
1TVOkmBqC+ulrs9O0mkYpTt/oGDZ6LBFymq3qsRarT1uvZI2CC+Jy0LKXcVYzERJ
QpMEx1N90slNvbo/Fk9tW0CIqCuzu9g5v62NvIEaVQzrb2cAqujjtULF/3YHSUGz
UWnhnL0Gs+XOCyjsNmCbNp4EItawjLiXPBtuTnkjZ2NoAi7Cx0mxhKKD6h3MgDUe
s6iXKYU6/AZRaETIV6cqLNZFO+nPILKCupqnk/xFLp8WbuHAzN2DpSNQz08djvTm
RMjB0HS2vue+LaApAYohvaI9NmZdJW+kLturX22wW3XMwlMRAszbUTaqsA0mZDX1
jq2vQbi0b1lPTI0NK8h+j7njsPPJl67LdGLbBE0E4tdTuVoN/o3sZnbDFah8pdu5
dK03075kc1knXhJn37BkyJP2GEjGKf2M+iN/aTANK36QrD+eRq/RelKeCkth9oFT
abrLPuyN+JfgHWMetkFLluUQRSDhKcXGVhfwFf7PZZ0ZLsMU9GGHugjdQJwe5WNP
TcJmMWibPhDaBxy7xo79OEXQn1iJ8ohW8lbExrx78ZSWdV/RUD9ke5cNjaNfeDn5
4cnmgQl8GWqXFXbvEIH5IaIOuO0e84X40IcPNvkvmdAj9YEKuy905GzX/lBx0gDc
ulPGo/54NtRt4ywbVhBPS/l2JGgJGiwluOYOrCV/vrk2PGORHdge0nOqgI5qR/aP
Q4i5c3U10oK3wd8cKOMFVubBV2J4hxoR0Eie3uqAwbnvwHN+CMtjcR2HrRA1EOGI
k/4AiaTQHd5sM5obTiXXnn2Nq4T5eVhHThQYGfcYAZxS2VQ0yCyUuhV9BD3s/PWN
r2mgvxo3tsKVlaNlDu+s9IMoeG0wNuFwO8dHuWVfbDhbQxlGePQ52/2RdU0XIDZk
5VhYGtDrHU5IbgaBgAf4ElUf9Ui46ak2z7W0D7nRXXZujIwOk1oSV98YYAGzpOPA
lPriAe/w1ZFs96LOK5gO+z8xGocQJ6k3DC0YiRJwq9hy0MMs/i6X/8Po2VOv8dxJ
J10R4ubgzwtjP5Hf3YgGuY1Ez8goXVeI6axbeHCR3Vme2TmNlqBDTt0KDS7nF6DS
SCCnO2b+l/si2aDBYD1UZdgWGZhz25HpzuPar+o8J3zs+AYX9mlbFAnP9CnttrlL
AUTKmrrD9Bbqtz4T7EisDV3427qPSo/ZTHnA+yVYcjeM+kHQiGymcY9prgqyNWnE
/k8C3YEuRiUXbPzKAsD2Rqcs5w9gVZZvC7lrjhrzLNVjMQPON7ag4aNW3iNwnjgb
e3DIEwUO88BRbQLDWIDMaFfnUyGU1S7U8Jggz87HaRJNRe9pXLqOXINWfI6AAv1L
cioAHeTVzhGeuPshcZ/Zrm0GhLSyQHB3FeuLDGr/lDCCTgOvYSgoR0BMFo2FWbtp
dOF44U5sAiCgOd05+YsWumapgnVTYgxPMFVihz9/fzla6BzWAa0hDHEDTKiGuB+Z
ewvxIzLrOVoDQK+filyOBlxL4xpw4HwpxJXr1GYwOOTDGZ4vCZzmcxg6dXxULFgX
vyR91qNanvIdwK6pTQ2XBb/18mvcLwk4ITcilvZo6ntkUFFZNN89tnhWmBevZts2
UIh2Dxxh0MfIsFsMH3XXpesFmAb0NRqb+dXyfSIA0rkyRRzHXULxx8HszqMnJmap
t4f0Ic1SzSvTSVJTqfltUYt/uXwET6IJ4cw3/+KwZe1+fyrteRGnLwhSDpNcqFtF
E8x5AcS2lDnZY0Vr9nWDN+EklnwT5AqfmfJwR2rn8Og=
`protect END_PROTECTED
