`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qsk1pFJhbFTjB3LSC4KXZnlyJ2H9q/SAEQ/ggWWqpSkFyK/umBU0Ftr/tSAhVInP
7jyRJnt55nuPLRWndTJAv8Q8Onslkms/VsZmbMvXhybppqb4apUxfWya4r3ddHjG
h9z7ybwUu3dynnuor81dhbZSDw+WWERyvCItJg/QSZLT+YfJfLcmdeOSXeBMrvjv
6UsbuipaLsWns34zM0TcVT9A6INtvsPgbsNRaQfLp7lzI2jwB+4WEniKl/wDuaFM
ZlipEBhxFKBeG/8hC9SDKtp3hvARKzF4OGsgO2wNyFFaoDH+Irxel2148F0LYZrx
+GyYKcE7lFmuVxzQmRq2H63MLmKvfJ7B064IXfw4zcYQ3NvUCJvHSPv8Sl9ZdsdM
mbHkuk6SxM2ZGxZUxcvBr+RZM0nvUdrDf/HEXeEoRNVLbWyEM/YipbsbgDd1NPWN
Tt7C1Kj/gYARrIQL4Cz43EQJqCGAaMnwfXZ8B8+oEb5EC6mBLr4rabeMy5LCNRaL
QOkWKpr0RxqVoRieuSW2ErgufKnCeKxRsa2HBRaaM57QiONwJgyVDFAXAkUztBif
5UMY11+M7RpaY58EwLFUAw==
`protect END_PROTECTED
