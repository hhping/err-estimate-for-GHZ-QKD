`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
au2vH0f1B6WeL8wVn5Ie2PU5wGr2xOodjmyloCjLpgZxnK4sv4LKgGVQUw6qLuzc
GEMoOGhxM9LNeUQbiLjQE7XILK8d/2Rz/GENpAyxojB6zHlP5EG2fCBZXW4NJV/T
6M5i/4kTzvP+0Lmkvv2OrmLobtL/YoMFK1N1peNHou3E4MVt4EbVrG/L+p4jWAcq
A3hUEQKEG90QxvOMqgAgAkPDyY5M8d08gZTNOLXO+swM+pKHLkTdYKvqYkZ5vjrp
v+GcI0XU+cLc40jErWcdfuVdnUkzMBqEJgLtFfRut/Lx0yVxjeUecuUey3uhACAK
1iT2T0dbn8gZ++5RdcWGAOwJ/TqGAf+X7SEhwqceNi3DCufjaqSR30JP4hod4FSe
yV5jLkH+wP3eUVuT69aWRHeZrUka0iyvJsHnoZOO7EyJMGFGS+eRT3mwn1NWzy/T
blEwJjKRcd1RWJ/EpREPmJXeJfZRRUio6v0A5wqHJO5HALwSvq8ACK8ptRZOB3u6
Zh7C/g8B5uEof+lE5iOifyzXAHwhR8hkmYhSCex5M2RMtJ3il2vbrPXPc2p32Nqx
6QYdmfKVI5udW+JcbJnkmA==
`protect END_PROTECTED
