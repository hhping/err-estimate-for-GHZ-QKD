`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
txOCrtebrpvT8ljUlSIJzacVJRsRTk3i8Y3ryNd+OfIRXaFV1zbzPpZN8+bq8OEe
zTE4nu5a/ptv/pof0REGYB+obyNB5qugc+Pe3txxdULVdLUnNiKRbG6bzu2OrY69
kog/ec07zEBbFKiJ0Ik0GKpj3SrMtNA0F4x1/WjXtufXkgLYhQcjS7rdYvzBuZ2g
lCEO7TLGhPj8wqf/EZNIzi/137X/rJp7+UirIQCgbYhGViijtnV815vYoJexakVB
4Vdv4ic89rxgf7bdusDNPgjVmgoqj0Wo1hGuJVT2IKx83JJVihy/JTcxMSw4LpqX
2YUXztpRsTPCPWuW1MqHW3yXoWgjvf1v7vGxbK7inEN0uyTlpcNHwTMwu9P+eeAx
bVTL2eQvRW+e+fjgfdajeueHCIcF3/aIhHTnEJXqiciR/Eli1PR8TpTo87AXzh/B
8syCgGseioGX/4i83fiscediBV/WnpmIpqOeTV0Nh3xq37hm3RjpqPdSwXPRAwOG
GKDEEpiFs/ZacvU6o6LV6TJl1sE58OmrvBM8rvspUVaHvOa4uh33OTpY7+JeEWB/
o1P2dQUTTj1abF8ihmKyjyrDiWlTzGCeCCwsz6iYGjKE5aTkZwaBdPGuP3ZwpLRk
QIqhaimcVbUqUFWPKnwZ+8dU4I0danfH5/yHkAnwAH60Qqsh61qLY04xmd+lkzzj
mftxVfw+Mdt6crto8rqciYaSW1QnJqaAHgYIlmWAVLo0WCzPd7iSzqxY2s4VV5g8
xBclcX9xYE9f3vG8yATDQeDI3/xRSY43Hylc/IdDNbgXTLtucyjWvb4YJkEDR3Tc
6mAXA76+bEFQb85VKAX/qIa3OW4ehKa3TCaJsrd89ZpgRUQj64tU4ylTG5NIERDa
gKIkgdP1MkdgrzKgFv7faU4EsLJr7Gbb+WmOD7GJsFlYPcMhEl2u449rnLswf7Bs
lwNn6oloC3tZRTX+uXzGt+6PAHCxIoCEiwQ3YNWavYHuD/6gkSFLpw6JZrf6FqD0
KdPzR9iGugMbHJLKDEYuhS6SJ2TtvLXLFf/e/j9ZL9X/Z8VtJLNPrdvVV9FFjrGD
tjO+jsx1ropmx/T4wNzYTQCdDtsVWVnwcTRuAHPbJ4d8d2eUo1qwAnILaeJY+pI8
S8VCsF8QSzpaZ90sjS+f0wRW0NoosOvKBUvlb+Pt45L7bbODW/Ml0NmH7kS2rExD
YpA2YJKGDtse8Ar4NrCPAdjDmuaESJ7FrC3/B8zNFLuzuJLRcts2AE22IZvyEeaL
K21UO/ugBb7vsS963/yhkXkwB226VfoFYzb8JPLJJB6IQrI+JGRnsX9aJC8UFoby
yZC6D9rzEOdcV6cWH+FCHxwviFhfa3HCuK5u0G7Ht9yaLSR+/llD8vi+tNPers7B
NGseux6Fygi3VpFItMX+DfORng5CUWMrkSHb1v+8OMPCE7YKWf2vu8ddrDDzV9jv
reXIaXQcZczj782989XbJnWt61r7Z3mw72pxKiRhs0n6FxTpyldZppT+mNfAkEqB
U5irqX82KawgmdPDx6yh1ABoehk4+tBWx9QHIGvuXSZ2NPjZYP2gbseYjOrGWqXZ
DqmGe9Wc2SKCh0n0lxU1qD8UO0ynGXNaPBKoP3FVL5Q6/BvHgZR1sEVEVMAcFo2t
3s+zYrpLz+w/p8Z9cHXajL+u8JLVN19uEe0lbhO7hqU=
`protect END_PROTECTED
