`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a11S5XYiZhnTwHPkTMHsAdjtGgEAbpM7p7c6Lkq5Z4Sqe16mbBB45laCcosd+blt
ktoeBWQfeEDZhu6cShUTcYCrzFsfvM6k+xwg1YFw1GId994JZObbtVnC0lGb91a0
HRjA2ygkDBbPoHryhKD7g8Ow575ykDCcYZaybMSRvCiU0hGUURs11Kcgu5l2d72j
wK3EvWeVC/7adtF/3bH1H5BDH3lKryK5jicPlgYIRTtAumauh/VaqAuB8as0UHZ8
1wtI+fr4ChVWnWU7IGR6EafswkIcpugsqROeMSOAOKXSa8lLhmzsSw3beVLenH5F
7tc25MkC9w6bc7GCKZzSP9PPnEDR6v/I3r5pu02PYgv2ci7Zk3LJuyWH6HnwwUek
k9G7rZpPeOA4TvoNKzK9Uwz8H6GD1bUGzHEENe6tM/qF4zAfPJ9epLfLnAp3DswJ
ttFSNG7zJMHraKF6zU6OReqZOFONd+ArRjE8Mtb7Nlk=
`protect END_PROTECTED
