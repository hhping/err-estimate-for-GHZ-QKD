`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zKW4LpcCFia+MICv82+McwAmfAc6cd6stQV0J79+rLEcd81DfY+J6YoB9Tki+o5k
71+0QFu8Morl8s1CixiqtrDQSNInrAVognVl/0subB7W65NjK53AdhCNvBEZujSM
SWig8lrobzU8RRMrpIkZSy0QNTlXvkqpjG5AmsiJnnI9yxE94oWZ4plvoBhqgRSM
zLsbhjqT//BWIk693bJ77xhuxORWyyqKHY3aFJXGaVgxxPztFoI5wG+j7Tu7bVEJ
pwsB1ny6DfYwlb3TG8Zwy6EgfCKABfvQF82dKPk192prbwbSKUxwkwlLLnm0nVf1
EA4BjVbUgMlqh5tfs/82JpO4JEDel93kXCTeafNAo8Uc8IHIMGiYdcvdE+nOjaCI
2wiuo5jOUUau7QtSuhCEwSNeCigmRHv8CIiAvPh5rnZoMqeeFMDDJIdhbCfDJ1O0
iYTNo+xu/DilTMA96FnFEcbaup3gRgJ+js2uTzWqbyQosHwFfhO6tTttPRYK3LP2
rHXd1oeONbEPAYkUZPG1R1sat02DgyVQuSKMRaEVLhaFUxy2sjlmxWWpr9ioH890
8PKV09mSeJEPaVZxfUGTZg==
`protect END_PROTECTED
