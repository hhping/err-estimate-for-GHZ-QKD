`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hvrFEdd074xYTSj7yCuFkXEJrWmf7dmHDe9D2ERYQLsjP1KwBn6oKWy3bg25LQMD
V1OnYNPfv4JVUlnGndbLDJPVV2Q2bJHSpoPdmc4CvnInAmgMkiVf3SCyurMXSdTl
Y8d3ImHW9Vsq/6oVrSUkpxyxBGrKLJ++UO8ZC/8zYQWpUeheNFYWlNymEk3bN0iJ
ObYQ8N/9iZDXCL9n1zZsA6/dHLbDDeyyCBJieeAZ8H4eHM0Bo2DuttEU9FvuLLGC
98EWo+S2y+E96XoSgI0j6dYPbfhPtiTWWywQLGlbtfUG180WM3263tzyvT7hqS+0
qIA2L+5kJ6gd061+uocr2ZmpdLuZG807e5Jrh5kc3E+Mm/yevmkvwEzk+MYXBsWf
2mGCDXgyCEwgZoHt2mlGkEJrvn/VCEEcyz5TkAZopSxAccViQfU/JuaqUNXVA4Wj
80GCrqDhVybcVLSe1KF2bt3T2uEh/LLid4a+JyFvt67QahTCu05jEn9IU9/LUSJC
0NZjM7hKd13Owktr8L88mpfDLz15RBGcp/ftXyDajhaqkxxUFBiTUlZQFxWROoRf
Jmv18h26Vs1q9BLzYBHd4k7tDFMjUJ+AZEYMYRwbI1MXWxIqO/2vm1/Fz1AiBgNk
x7/0X7Uu4tJH0e/n3t97+d0wnPAaBtwvhAWNbtlDvSFstfZ0cQUFdD+VjITt/t6R
J0UPmclIWkvPs7dxjyy50XQljznaWm72JgXstFirENtb0en9NDpIPllInZsAEkjt
oRaAqStFmWzBFdfefZZykEJMIUs6fXo5k8Mr1r/qrkyDn5xOL9XOCtJXAHqB+peD
d3y6lkGXiWXxxS2WGX4Wmc/8wWMm5kEiX0JrosBGkiuAUHKFEpGQBPTprhzzSYmE
E3RxhdEo+jhyX+VPAW4WI9dzv15uFNSDofxNkamP3VgSLR4u4NIj+qONFiwFFhjO
ej3ulJt5IBoORo16hcaGDfXvi8xjIF1qnbMiYBUHjqra8sihPtNTapRn09KQRagb
Kwca6Rq6Yc1Fg7rZoC0+KFKP80TyZJBDoTCxNg834e2StUi9WpBeq3FUH3wSSWY3
C3vxW/r9kw8MI2Aof2rTeqePVblU+3pLQVNFGVZqFhN7L+xsGk+eVbdQyx8f2CJE
OoLH3RAii8ksStuuEs9OOaZ7PnxBMktKTm3r6dhml8u7Kd1bNHI4C1y5BvXEKRkW
mWlMlgp0CxX4cBLNDa1pnfc6cKVS8xwUTnydgjpIKy5Ap5xrqW0M6XaJ+lWdPmdW
AEZZyqlRR5PThB2LhTXN0lVYe6ntXCO1YFU2TLQoQs/+RHfL9atiobvaJQmqnyY3
uUs5tHEy90X31EadOBaqH84R4VTVwpsjc88MJCfnSsokiwfcy0o3kk8owboWi8IT
o+BVvolrUcsfx+aVugJV5F5ckDy2fAcLQbHslfAWeFmwoGN5vqG7x49O7/Z9bzos
3UBZYioHIWOr89/Q9lrImCIByLECQNSWTm8QxYCq+7bvKiJJTUnZ4crEzuo9zoqM
HRIblz/CZ3blkisfGaEP55Tjq+ziZlXmBPuNxS5LI0vMnKEX36QxzGJG3fS37n5m
9g0LiSKEeWez7tXCFd620HW4q351IcFUEsJZ8mm8Y0c0QJooPhQzlno3k3eGZMAU
NWSTZuHrfXYitzl6Tw/V8KW7/41bHgVxLeDajZJlzmDpH46VPeEMckZwvvz2bkoL
M+cvZbCSI4j4NOp020knTpLeQTZ74BZFEl/RgtpdBf0PfZ4DOHy9EQMyiz8MJWS5
jmQf4I1GEXIi2JpA4ZFHVwAdrdv/LDSgKB0IgHy8B5wt66Ho17SgiWm7TD84zvBe
VVwbVML1QJvXU/6c4CWD/vPsyVu+L3hqTf/t2i8Ry7cUs8xBM/nZCBL8IXj4+bEG
ctcriJ7kqaw+AyxvKPieLi9QH1HFa8RiUzPijHswqaoKtixkMUD2ni7f/cSomFQB
G3Vi0hwl3fTnL9zSDZUvzuBBUji55A0oZp/V8x4Bz3BWj1KXcG2BBRMoktnx3kgp
ZvHL8v13bXyU5fAYB1orWh3XghMF6lw0SpLVHLeqUjwobOVS1wG7D8sUW5rpSeZd
y7p45lUT/nuXw1Nxx01hXxRlL9vNo1nQ5obuaW0IZH7EH/QWPnpaOTppWJoSqtM3
C9hn2Dv4lcKs4hiYPKHl8GOM7L3Rr1jedC+/8O84q7dkecRObqWI1eiEyga26+kx
a1deVIBq8/F9eV1u9LQhfcixjTApptSH5QvmJ4iEZw/LqL2BDVPRa0mgH2dYoZsA
CFXGXOFWmxwhz+HsX0Kfkq2EDdk/XIrUXciZ7Y9mZHU0wJXds8La/emuBGe6CXnh
WTNo/cLsLTsk4F8o9kheLT6LuKL1Bik4aw+7os7YTs/BfeWYhnJ3vgrfZ6EHVEfw
cGiMUtTre8LJOiCrSkGQaFd4ayqSn1Bzb1EEbqk/rCUXMXE2Hw+WMbdrxaCEinYM
bTUKtMVMVuN2AkzaKWyv8+BVUc1inZK9f2enIjtuinlm6SXY40Lx1qi2rVHTPRyN
3D5FrWkbjqsC3nBABL96YGg7NBodyLcpU1WY3VPAhlz20Iej2l6t37PGKeXgAJOr
Ix6HwRzjR65xAoiBUhlA+i89XeIO4A0jQk03wJPdpoYfo1STnSf7Sniw0ppWVGJY
Aho8VAXHdesxceY+itCL1VGuIjF8utlbNXCgpTYo8EKzjVFI8Te4MafYOXSbMRxg
gIGjOmX6B3m3XdTwoCCNL3N+QBNWMzmCduYRDRkV5fiZsklr11ZXSSORlTURjltK
+YqNqq2Q+IMwlYlrwTGR2VXYkOsgj/DLGOVezEiDL4zDhK1NBzwWIKaGmfCSBGdh
itxwsrjV3J7wkHiv+i3cHKy8qex+b5HuBywVyv6evMeXZrj2v9DKZ3TPe6NxZRYW
Iu4xuIEaxLEveUtp4rcU/bsyg/egzirgUGaIZr05fWhaclf6lOuLSvcOH3C52EN2
vzfmic02cn7yx77pWWrBAxAKN7VNIibk613x+HneFW7Kz7khkGI0lLNMQjzaWtdr
Y7MrCgpiYL2PIP+TpuQa1pQScqHQFZGhItx/5WEaIN+SAEDY+VO7ufOqJzPBPGWw
THuyZJAChkUcBAlvjpd64Z3W5jCeRJptfl3h3wqPDGhhPIzarQnuTQdK7krnVIqY
AyzG2oZWViLLwqRWh2sz8w==
`protect END_PROTECTED
