`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mmo3vXGmoDhGI0SR9oPOFfuaJBiU7iIbKafYGeBxMhUsjBuRYnExy7X7krOUtMjy
j8Tzr2PvCFAvRs70bV31MEnE/QDaclE+t4CC+vDpHT+cT0MumGbO+EhAHbuYgKWG
QqUH8wZV7nN7fD2xgvSIjNfYUgC0FBTFZZOG08qUtuFmBoaAdHyrrzZxHC1aiYCm
15aLdJFG/lTspgJIAtq7S+Qn3CkzUMKpujrqqe60PZdf+DkQimu7+xRz3NAfOshr
SkTXEusFXR2P2P/4D8PQ03lmJJePSQJiMyQ5uQfeZ8Qs3NR19uq+LJbYf2UEmeF3
X0lOkFFGRWr/nohTVrr8wi90VwZ+Zhptu7SP03cF1HyTJahSPI6ZDyEBkVz7+vSV
Zs+NU78X3Z7j9sdeC+jYt9DjdN0vopehjTzJrBZ+9EYD8aawuTzgPPzFToLQYHxG
GoqDX8gCXhthZZteSa02GIuwytgnhhcTpvQq5Ti3U48TK8KK7l9uyzYoFzx6jhdo
F6txZClj+3JxrBjZYZKmk3olHY9PbDdyxDCZsRCrdQGbCKE1ua5KOtyOFInaJgWX
Exx1daGRP1ma/LW8Tb5p9oFm6I9vEX/QRdcN7SGpkUYVlkWOGD1PHwsqPK+qIsBM
WoWgXuOfEyAqkp4xrEp11XgrOYtRaNnYVGjZ8KBaTz21LsWD6qR1ki7Qjsw+3mJ5
cM/BhB8hvCo20iXpUrvj6fqmKlwmMSVsKAYxH3mBBJzI8Z9Dj4dor3CJ5BzR3k75
R4e3LXy1o6RG+qtHlLuB5QrfMQRmkKikKWb+t85todLxc5PdeQqSSIl9CUd+hWyD
sE9Yo7DW7GPmTeJX5/keXmcJ7x80oYp8Zlhm0NOAHKQ/Iu1VS8xRbM6bRSqMAvn+
Y1awbIY0iDjKXBTZWj6qdCE70bz86FdmMcSEm22Fi1ZkrZsq5G+46MTF9SCQxQbd
DeVhmNvkdVqbGJwdvovTF7iPo90wNM9BqMO2ikp/DTSKmAfdGB86HwOHPGJ1rtIz
1BFM7KX7wtRARjqd2VBrBb+6HaFsgS2yYXXKogAQFZaHVvsd8VUZH1V1d1zvNzrR
0Z7vrJeJbVWtbmKbo/iGf+dbfstHkSjlaJDc+oS5KwmRormx8beXdhwUIe/GCyNF
mvdPjgAmkAIx521ThWcmSSzhcjB3ZZanFZvSfyZAFMTULogszeDb1Tr64ABsBok6
wTbsq5UhS6AnBdlBzzxpPYYpRQhBFltF/tPzc64a+PrLvF6LXV+9EW+bh8xA4KP2
m2L+10AQ0PYnmA+/URT8JG5EHlJ7QBZG1QhwElPSjcm4gPQL3eEbQb2Bv3jpnj/t
R8EJVh7q4oFGSiG6Z45BOi/FwSgObTDPGDvAwqMK3hJmY+q+J1Js9YRw/ez6FMCp
XPnru0SCsrWZdPKOEUYwQhB+tbU0IDfF0QJF9Vazk9lOz75gdy1gzYvMK0O40RBC
DqIiJXAbZuVo2GmTMwVu+xV17/8fXjiwIHqm/EK0KYOSm4wZ6gfLhq0YgCSxZLQc
92DwGuBCLLRTgY7EEyWBVXocLV7gWuBjHmq4HhcPV67UvZIwoRvzPdhBmfRSYmpA
Eztx0nN7UiqTRR4Gf2QshvGDoDhoZ2HxeP19g8LiEnNoTV7e/3EKY5srkxb3aHYT
NE1Q8ovJRfLSjw1snSCKabNi+z+KGl7o6sWlXgZ1tnDjwXhVs9kDhzO/Xzs4pggY
k/GxvnUF5GoWS2HLlTl3C5/0A0IPKmEQ8BEKOwhr6R9RxbeqtqfbklzrCQUOG/7c
lTcYpEIoHGZS5ex27vBVIdAcE5eD2M0mqK51c7rAVYCUP0WFXDp+nDlUKWa5fqAQ
UFyW4IGVdq771EWxE8dtQ0LcB6SZJaB88PS6oEPE/GyKrII6rQX7gZuVyw/XLe6u
EPnLo0wruXTZpbNlxHTGXFtHjH19C0RjRAtgIa6I6a9Cucd3EnakXL0BhAITP8kS
O2ERAiglbnUwVAUQJ4shCjYXMjV8ZqnMTpomAbuLDNgvtLLRlCfVNY2o5JgTXl+i
iKzMzrJ2yWc1TJd6y7Zsy9O6ejb06/cIYkqxyW+GPa1YkAefpZZsmIGFVjcYO8+2
AixihT8zKVaHz3hoG9OYgq3E0L4MTpbwne69y5ztSdZALl2T6v3rR/Sk+QorlYnp
aTG6AD9VuS4em1eLQQrb7JDgO/BuD/UPa9lOZMCvOk7hjDaY36G0VNWKAPv6PSK7
nl956pox6lXV+VTdiQOAgHmY+WcAKPt/O3A3ikUbK+e7V17JzHczdUuU2ClTh5u9
hcPks5xmz6Q1YgTXPteV6wGaT0tB1SjOu7O/II4RG/7/OkQZBFm7F5LOKXYdPVw6
wCYPsV0QdK82j/6MxXkypfOAK0+mlQ0Og5AEzXHp6VSYhhbSKxL51/19pCBMWF9l
45zbkggY6PkfF0e3LECtMJwY3jWXNimO2BfJW0plEnejSHUolIF6mjp/y+bLnVno
KTwGq4Idr+Xpg/SUxyo+e5Y/+9fjhYN0oL2hotiaGxaPCH5UUFZsKiHGPEBa0BF5
+GyUovFoH/WolE1/yKo/yXNm1cqwuyzCvmuxe3xyYALregEovAxsC4mBYSF+qxAw
OAgqdt0ccHdd/VfIhmA1L5TNEaRdgKZIO7gaaUe4nNMMoSvZ18siN20j0bdzcW6I
Im1MGY+PggNBoq6bSngKDmuTpIc0maVyP8AP7DMQ5YrXOwLcMkGSU5HRGavUZn1v
/80bvZBZM2IhoXznyQnI022/4hXjSnHeKoj0nDzJ8QoUKi+XzHnA0dAyrCozWDFA
y+qUgLjXDdztSSBSneVPIAE3jotC25ib9lhrwTGxv79PYDLP3tid/CEJM5T8KKuj
lG/jZvj/CJIw/WTUGliVJueDWKsP75f6pPequp8PANHVy06araN+0iad30SsKeBP
KvrGTvvxKnuQo+MoiEnM8XN66EcXhL/F0y3mXzwm7aZgcqw9cQqBPlYpcm2jN1OM
RyJq0w4Ds8Ytx4V7mYm/KAExfhxm2ue/r3togqKusHwhVay/LEjx7+JJaWVM4fdj
9W/myF1TJkho65Nay2OKXX1YE7DTVZ46LKrpK14Ff17O+CefNOl+fOa1H4lvbMVu
5PfkKd4z4sO4W5kjr5CtOv6otV3YZm/6AWunpWE9WXTq/7yFEE8uGY/Pm7575YyF
tZUJ12t018PomQABRCQ+3FIMiopVI1ig8+EvRcSo7aJojI0751QCqyubFXXW3oX8
E8jIW0lRbc+skXs7LtOJapDMNkPb8B0hKMFfTiPEtun8Sm0+9wscdCCbPBPqdybY
spnfkLLXaOjVJYsP2yNXMEQwcT5OAz5G+C/fDlRB6wVFQQVz2xIOxrR2OuCuSO9R
yQ/ZBebQxg+Lje09TMFz9gV1NRCGVy8kctfJDHlRV+hginBr/FTKiqlTEKcaYWgB
Jah+pqtQdxLJzEbkEin1XHziIyUycng0qsjk10/ZG65mDyjbrbvsEfBMJ1MrcEmL
vopnynrHROQPo2Xqe2g7cL2NC2dmwiyZZGbm2765xgJWsorMbclD5bj5RmuIQJYH
idGD/5tZxKbblhHHRXVHga0LPZLP0XiQD8PUmokKNW/6aJ30sUstXrJBSebjbYmC
t2VfB7Soc2QZOcotEwfUREWEphgLNjeTvOsvnGuorTMQ/KLJzbH2m8rN3fGhRn8G
1tQMEpuJgYbUu9xvXFFkIGybgO/nf4zqZUW9JAsw8cHJ8GmzyAQDg7AGrQGGhKaD
S5dcq2LBffbUXDIhr6fV+NAfUzxK8U9Dy+QvNx+kQAf8sTqct0bswkyq9apJjTBw
oTIGiHutZyNUfQHiYtUgxDLiJ3aqkdjLBJvvvrKDzgHIdTlsj2DVqnHcBDIhRNfp
0V/whGmhw5Uj5F3C1Kkkiaclygm3zYNUm9DRxk4aSMxOgf1ctZCSNcDQkCURLLfJ
sSQ0txEFisuxN0Yg7mDVhdClVNmQjxBA0NWYl3bRfxxXfWfPR2/Jx0+fgLsSyIN9
Fnrgod05hhDIql/kFxjM1EsZc0F0I4lR9e+PN2QU2Vg5nKipbhe5cf5nTkwfRO2R
ssEmh2c0gC4l4+gdAl9+CI3cPyMuUL5DgKgtzLVoPTQ=
`protect END_PROTECTED
