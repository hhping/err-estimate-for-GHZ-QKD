`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
emmcVU3Ac3tg0/tHgN7xUo54yhSDqvNQhehCjb0+AMCbI6KfVe8ZvEciudMLWH8U
ZJzwgvIZPXVtXO7KWxARV4eu1rCPFZd5xWpHDX2hFim7pbcWFEQokeway4kLWqyz
9p3e26jknWzubWa4AQolW/piP32QKNLXtcEziRFhPrp5AMeRCVZ58ZsgZBGS0jcV
3RupOBGeManME2M3M7N+h+H/5skbxd2mado8R/RLcwayuFHP9XejgMbRrY/fGn/L
CQKfpGlBpqKAN+17fZTutjeAuLwWgvM0PB5d/NlN+IFCsN4ZT/kM+crH1N9OBLzx
RywTwOBPhhse/qy4uQZVBRszLpwJzwgxCfzNcIugwboy7lNRVazwHCYLQopp4Yzx
pKeroVpzITvaUQ50tWGZyNBuRE7Tpi10ozQUFzUjFebBq3i+ivVPGX34leqP5a4v
TONlI48hpelDBShOMBlKL7+wlz0dBCUZKk6J/xxSNrANfUDr5k+NkPaM616AAgjA
ly4yvxXqceXjY7f1KIqom+zw6glbSXG2G/aSH8DvWTQiPZ4nHcbUC1UY3jsHsxGz
yA8p15isOb855hzs/5QNaDTwPZh5mD3v1ukAfibNB6u4D59IE/i2zPUDUcPON8Px
o8gRBKyWyD8F24PrS3GqaCb4BD51nYs8QR+s5JyHESOmcCD9W5jgR412JnpXcPQI
4kghIpWPTlf9xwddQ4hE44R47JDct/OuquczAiZihP8ZZCSb/MSdreArxE/mEAci
b5Iy3HJ/MzHCosjzL/uFZkgB/ZgzobBfqgFbK6CVNzAYDmCGmtd+KZJFfISN2KS6
Zl3/Ll8Gcn+uHRkaj8jTAME7fEc7Dsqcs+jV1z7oF3EBJDprEF2xxjajrQf6nvsS
LoM+b07q6mPYfuKzSvJp6WL/zdOJWqBS3PSKmE8qdF1HBt+fGdTFTJ4AMuA1buJI
njXt57eaIbNUdFr6YLGsJUYe3Swz/4qM9Vnyi/4rzjwaSuR6RIJ8beTNJbWTKwJh
tTp41AWDIxWY7R+oyJn18JGxfbL0PzLNKbocRQZzNt4b28uCvE/IBlrlhd6+xACQ
ENjdCOVtaiP1MXcZJbVLlOsB1TLHz/oK9zNgWJWcEl3Bcsm99jxiDxI4YTK8cCYd
MsInEzqR7NLANhoJMlvGF5gJxTLMMihKRW2dVpaRcTDjiff41sNNQ6Hw8s8aWlLE
YCCY7RPPNn2IZoDhA/oNUbFafQekmF8OyryhIXNOnO2xNRApphTY1rk78IXHego1
u3oY5akIXqu+yidKvQJFSIXvQZX0q95RaRVIN3SLZ4GuNYT+xIBXn1b1p9TPOxiw
KKLdkfObyoy4QPkJkp7boCF38BT243E5Vp7y1A+xZFa2hn8jb1P58mmSzddMm5h5
RAScvbkcfUogxkSPDGGiPDa0FNqH39gq/TwPiGbBjY9DHoC0+I/xx5GdIKlA8p0n
XYVxM4/8RfUpVDsmuNSYKKTiB0aNGeZ27ie54EooyVH34j6nlbqMu5lRLJcTpRhd
tc2tMM0hclTBwHK5VM0gLg==
`protect END_PROTECTED
