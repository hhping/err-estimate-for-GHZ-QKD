`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sHM1awUKpc+AEwWJ3GI9IRpopFJQQszWR6IIqH2wQP45CUZ3WOp/FiQ+DUA7QPxn
mqjesE6/UWjvubG4YGJMsoIi2Jrga0a2KysNsVWlsQg7x9l20cQH0kYY/KOB9y44
1ENjBVt+pRr+hPIN4kH4JmSm0GMqfqNOI9MMBgmGYk5XJ6RUIIgvBEMnMYdoi3bJ
knqKRQVDVw4FiWuzbC/6xNdfxLfBQuQ1u2nWzh6xcavVVhD0eQHOv88uyxBWmiQD
0C8QhUJEdCqZcUgyQyDk4PNQtWsKDKquhJWibQb2wW57Pj2D0mXGREAgOgK//2zl
wyo03Xf1DagFGbjk2rFg57KRnKm8Vp6q17kRrtcoQluM/yuBvFyfqOkb/4Mk9hTN
rCd+o/DiUhHkTmsnWvn9H17TPX96emnMh6m6G9yTO3ljqxZtcnTWVYRo3WeHCVrH
20XlP4FvttKXRg/UF3EVz8CaBemEXQ7xTABifAgzbpVbQ/QSUgHDcpUIaUSXp3ft
n/dtSq7WReTrQBGX2JNetdH1q62kDpT108hqMQdrmBWLL480EFU3ULiyrOciVxbB
uoDOFGPR1UbfTX3B1cQKdMueWN/16wTwVsIzYQB1e4aUF/umCN+2kFy9CXyzpkvN
xya85YiEFa6hLsBD8FZJVQ==
`protect END_PROTECTED
