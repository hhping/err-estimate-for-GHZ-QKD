`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IJ+TRBanclJYf15cP2nNotNRRA0Kk/eRIx0LjDbWpKj5cJyD52+gRqHK3K1Uw7Zl
/6V4vBSck1j2eglDMPv2EUwxoYy1Guk1XCI5WqzVWHDDJ4RHFiWLZGakverQYaoX
FkjlxwOxX+Y7SPh57ZlAGeug+aDjHVTz8o1UD/7A5kLcaBXCo5k3XMYy4VJEEJrB
nyt2+NIVOKSMbI4e50OBzJNl+KAHMWv84M22kruMQd/pT75gkovnCywZbKMOEwwq
cd5is7iygOQHUF1SI82divwc/GbNmAKl5koLUgdzcneFhbCtdgdDvK1w+v3K67Zg
bOxLoUR4wncJwl2skcBz1uarpsqTCDt0XVJbMVsdIzPUV3hNqfH1K38LXlj8iwhH
y5tQuLTAunlvDkiK6pblQYCBcuGp7m+Bsy8kFrPUebi2NGwh5lQXgPtg5kulQtrh
7GAtPMcKC4TDu014vAlEw5QyI5wUu3RJEzsZ4DuYny0JAmav0pHPA5JyI8vc2PHp
0lYRW0icJ4pTkIdujFcCmFova/+ywyuFqXJhTkpJSdey++iiv+fZkseMQ3PNRX2a
UDp4IRcBjPrseBnAIyTatLkQhDXoW4lleMjmQON2irGb1276STSNiH1mny3PgLDS
jeU+r4PdMTZHB8EiSRrJmPB9zmhKIMr07BPn/nHKwVDU0TopaswmjzqZDjDV6/Nv
eaORcQdhvPjE23X8ObOq0GZhMgSIb4sIMxQ3urepel40Kzpiyug5bulm/+17LH/K
WGQVHJJlA5ZkFL1fqipYpDo7hZKQ4hKmzUG4/nVl9bkF5K+7oiJfCe02rielf8Hv
fBgyXhnYpf7BYH85IDw8oAHkWVSMrvQEzfKZWPLjjY3cEhZ4WCpqtuDV5ERNhSQd
cZU1cHzL89pr+YQe3IOYQn3wtmWg8hooR8wesBj5uqyLl6uEDcvvl1mfecSxvAML
BhDXwfF22p4RG+0VQPEaV4ON32Me95qh4fHeGlUB49LKM9H6wKcFg4uIyb/erxSa
f1Jxr/wIHcTRulroIh+gO27R0sSzCMQthQHdyjrfoVSa1LgVR56b7KjgSIJul8X3
VDJ92BdSO/rTEI65USnwl0FBYSDlQYoD2EKsBoRCpQvVMql+7Ox8WvY62RbQIqI7
OPclxaIt3CiqmqshN95EdzQjpMNa6h6Mxav2CQHBH4FN0SMzTiMgfvE5tsXZeDiO
+NzNkueW/LjJnbvaEZSHaexc5tsuJzVgQ1HZSAO0fQ7LSM2meq7wu6qNUgJqi/n4
F8h8YHL1SnjM3sTywm7yxlYS7O0VRfQLdCAYMpl6OtRvvD/PUawgt4Vs7WKwYfB+
MX9s9y9O6LjNjrHPGGqKmS3secfR6rA3jQAUwfOacQ5Th30bTVk+6IpdjUe6Eph6
2EQ5V/GhTBDkw/RuPfCrRaZGIb/BG3BcqpIsIIBfvjHxKnCcNpmdtYF2HL8bSCGZ
vy/1vELTciE9Mlwjl5vrX+39CvHVGaTNTuRTcjyytbE3WXvErOx/Y06c4jHbI95D
fIY8Y8D7xR5Ri7j1lkhAbglqPLt4MMcJDexVgHzt/tg81jj2KKuC5GbmMA/W3pDn
sfj/j4jbU1PLLP0UGTrHm+dMrpfjwZEAqVeBGRqs5/dDLjT32ETzuUku9eE07MSZ
2Z5xXQuMXFEDBYSQh5tbYkA0p+N6zwGn30HNEsFk2ecsZz4GDFFoL0F39h1Zyxuk
0SfPiZ4Uv+X4Ppo2M4JKx3+HcM94fsW77UfaOYDt74uknHLmgERYvavqaGAkeiqh
jdB6DxPh60TxfmtOTzZTdwOa3oCFM6ZfnBuunr/k7i+QSNHL8+2KCZusTpT5mYTB
ADmyYjEdp8MVRXK3eXZyd+ziSE5NwVYPzyll/B0+3hMV9wRspJdwuhPo7M9H8e2t
W7zcvi2eWI7ptHZgga9wTNGUtWJZDg+EcURzyg3M4pFB1kHXcFS0IvWGg/ltcOUN
QJBB9VWIWFc/98hfswX0FWTpx0PGEUvHxaXMHwVjwAdzV9o7CH2hzyl+Ue9zEanQ
AY26oEiB+Lj4TvtD7Wp/5aRvlGmlnhH0HcCa5OqUj2ybU1S5JGoquPGO4p6f4ph+
H+qUr4YzCsluoIJ+FYFKJ5auXVReIYh3QOWjdfFEWLBhwT+r5P3eojcwJ83yF7we
`protect END_PROTECTED
