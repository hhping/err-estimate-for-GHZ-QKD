`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dW3UtgI8v4ewz0vT+XQtoEXjD7Gq/ncyZVedP26KUNt+AWXmo/2IUp+bRMFTbGyY
sp0WyF/xfdlYYuS0LOdl86w/SST5MjDYyeG56Sx1SXAfb7ohNh5FykzN+r7Py7MG
phpMCdYPEpuvP0uvhFGloS7n9VIIh65ZIJe91eA3tpcCXhdUxzjZ+pmLaU6vaRm3
L6tgRKRNdmmxjGRjPKob1rioobZoU1Yy4y7ZGN0b6dLOn6eqD6obo0IxPbgXLqNK
mSSoz8BZhJ+Y4leiN/7KrfcwM9s9Zp+jXP2Bg4V8ZZyEqbKFXOSyo123qBBN8ehx
nJYXW8rxBBMERdVWF72p5pvSQIlU0DUosLPwFFz4zXLNcYHiqHLvqBRmZEQibt9v
fro7WIIr0/GInUhFtOpbv9/QnB9Nw8opZh+dAPIB7+7oWjuYRodAasdNW/3NKKxG
4pim/ZV5L86WYUyWQE8Mig30BjRbcy8gavHaKdDK8KU8sbAPE/oDk4cH5+qgsLjW
dpErN9WpUjkLAOQmBoCIyTN8qAFJIIUryupZ+4Hyg+hOHEntSA5PWCn0xserVdFX
QCHkHHiUW1/kECI4jj1yTQU/JJ/xcs7PJtyvkvK/OYRRqWaf3K4RpE4YBuKmEURd
n6lcSMMftvqfoeMeEqxf1AixldLZzboOu02KhRnA/6XJOIHF8ios6zXet0jDVilW
PXaze3oX9qHKWyo1BmIV7g3FpOh8xy2xGQj4Uvo0NCgG8stw/wDyupmERkAmj3TK
3VjH8WdAqkSRRiSd9f/bxDORF6bITuxVQl4rxUtAGY6aHjtsVQ11D5Zlf/WBJNLQ
8WJTFviN1yNA9o4oUrFQ6rg65Oib9RDrjtdTlVOEXU5fXumDszKqI6r7uJj0Jxzj
D9N2td/87gGs+QDQEf62Ri44HtGHwZ58ZI7uP28/P49SpsHBzw5wpFqWg/xXmT0B
YDTNu/JeinJvCJW8l20rnzZX6E1D8C9qUXkj8dv3TC0t639Vh5DuY8vZAo6qhRCB
vpAx2xpY9t6CTcsyniOGvC5nqWks4ZaETIlgD5fYjfw5atS+7PNRhMc0FaiEjRpc
s/ldNt57TrwVoBE0msoM0tbTHjXVcbqN9MMmytzrCNNWuswIv58nvcJ7zLxfDK0G
Vs4O0Ep4pv+yZpSyT9vrhHiIcM/FRGG3RYQWe75Gk0EOAwwLKjTYMYNcf+Nc6zUM
WsQH2abgeoVfARaIC2AZaOVfrLVfwXXs/fdJXSfBvnnLCMsHOj3poZf+oW2OjFM3
WYnRl0bZRkWg5A7Y+I5TQq9qEZ/jLPIRhBMJCEy9Lrfy6VyecVkU6FE3JGIw+NPs
I+yF3L3lMhDaPcnhASXFEg0TjbK/nKvG8IElQIq1DWahAGOz4jcWVIlbjp+8oYAY
46v6c1oeUET19KE3ckxgszw39JW2sGNvfeAlZAUDupB5tRpjRhumICBJ+h0KLrkG
PimCOZEmrkLv44F7nvDvJlYeAIXZMxgaczLQaho3Cg+0jewj1VnWFVhYlygcR8wZ
VAKjyM9QkIR4Myl6kjS2HMUNot2gP6FHMZZKPOCnPLhhMnihOpVXOKks0hDU6jQT
KoxrgWhMOu4jNPCYAdgz4gjgNR+oCp6JXIcfgNd26/qLRgkLixoMShVwOUQWSRP6
CekGMnbCp93AIEDwngcqg7Jha1mOcwKupkaVCq4JTCBEy2jAcsiM4eazzYbLcoUp
AKjt8/513Oo3XpUb2LU0p0py7ksHkQknaHtWbwi0zY4fa97iH09cFGG5NpSESClv
600AQktvbbR3WjqdpVG/a3//euSaoEFiR+ClOTPvsTmGz9n/zysU6ikO1YT7S7yx
Z6GC5KzHtXT11CGRvRKW0bJ2fwQFvpAqpDJXgpXb7RwCg/XyN8VOA3Z/IpllB1Pk
vOyNRzfqB39gEBWDR1mUv2PWAwGAlPJ8QtORh0HHIk9Rp29tW8iRHk5HK8306//B
A7NoNX3iE6ygQC+jr8VQ3SPavTKOwZ0q9xYx9wsyrIdTe1UdjHBUuxR8nvTOdzwN
HUmBe71Xu+xGfZ+0dqQqehd7w1dxUIgj9Y9ZGf6R4f4an0Un2fmbyw1Y88L4oaRt
5EAPli+LVNf1rx2XyrP0mIYQFC22mLuzpK65zIOjtNMecoV0r4A49WYgT2vaZ6jt
pwl8V1tbbfzn2EPdkq5rjTWYBbqs9KX845PFgnNmN1qxnJEeRzdOf2/6Q/O6/Dg1
eRbECcD6dBVpPyWngeEZiX1FoYDzfYBV++0NXOnNEb2a/UA2lgP8GeA6CmeBIjrK
GXsDCdIjgbl9nTGR7cSOs0OV7z8IQ36rOFfaIIwduKK+YQVaBXHjkNVVRMDj4H8d
GM7qbPmA867ioeHhPJIfz1FyE6oMqOENKKuHXjeD9qjnP0FCu02cXYzhomPeyf0N
lV7h1hNu+H/SRpr7slY68X+3i6psvlxG6tWJe/m7ethimikraqGoi1FwL2R4LO4w
G4uw9wdc56j3qudXIbsPlxwQSA1S7KNkTqQAYZ7UqRhdJphKVuRlguVQ4FnCszPD
Nhbw6Tz5dfNUviG1qndug1dwpd8gaq2k2HY0idW9mA8dv482Hl8aIqO+Pf1MtoM1
ONaHAbGlzih4mwwNarBB69Sy3bO3ZXp8l47Y8/BsMJ39eiftya9/nHTQ+Tqdd6ga
R5YslMyMFyiCPCLajvYiHGvUWKlBXPB1xvYisKkQAeeobJaKB5yOF1wS1I0L5/DR
wAB0lLx/Z8sDPC/1SK4BlhxviGLA10HzRVdK7nuc66ENuQljAI2KU9OwM86BNx5b
C52jojfVGJ4oQaP6+t7TTQrpIk8zg7UBYj8B/PZl4JaUBRnmEp4cQ512ysQ6+nCe
qNuyRGvPX7h7e8hlPYMvHgmKol+YTKnW8PtLUcVqQvkseKo1HTy0PQ54T36FATH8
93n1NmjRHwaTjBgeFaUI62HuzmG5CWQCkOm6/2hWN1o72Z2mMWGxAAPdyAQ9pEyw
2zV4LYIzrKdfk4AKldrSlsDpP+bDmrEqfquPCR7O1MByOG/gVLEOlS1tfNQFrDkv
mI9NFms3H1MwkIKoizPDoejrjUOtzv/8PbBotze1UxAcM8Bf5xLjRHC4pXRGbr3I
wLMK7UWA3P+B+JN+L3n5w4NKFTv2R76LmPUfsAigYYcw+PTwoB7BsJR+jNCxCJGH
c2lwVUc0MRb4NxjmE10gdhXagtNjYQNYMZEsUwCE26XB+Q7F2SZuquU7MWqaK6xH
kcl+iblvakgBzJyjnvsJIRYkWLEXma9ZR8mMCdigWitiH1LquFMydwdy/O6wDLwd
3Obbuc2i4zSOGB7EAau/wOpDOqdY6jH4f585kuEoEIVX7pTICqYEWNQvxpdAIM9c
/pQl12rxIZIPqMM3fPcWNc1Wo74hEitEueRe0ba1BPoveCtzuyAV7rHnEoF/Y91M
W0gfSbTVprBXX9FkC5Wo5edhWWSbbfhWm8Wn+wY2U6qcpBVSKVXb7bID1yfNSysa
bw/zynFV+E8lYzSTdHk8hIFtRq36C0dVsbGHZw7Fs6KZjW3EOJT2ffezuaFT2n3X
pnMC2SGxWjiwgk9z2mg6uroGNBQSkm4WgniZ18ql4EVT4gNN1pfDIrFr1gFYHMTG
C+c7CfTeEgPSL5sQdbNupQwDV3I0sF3P6zBpF4ACEy72roScELXhuyoc15Qn6eEs
hD9Z1VdibTKEAT1HfLnfqiTLyCDd8kMfLO2XECb6rwILiNg6dcTXOPu4hx0pvyth
kUxfH1tbQ/5LYWZhuQuCisIuTEdIk74aruyJEFCNuUBYHPDGuPzLTGFJ49zn5eaU
WFaMlIyIKlDmpcHqM3FOuFbrH1w0FaGB/cADMIU5Z5frlH9cu6+DdDmpr//BxJKm
6u1LzOHSO+8qm3ye7xtLwY/wh9BTZRcYWNBY+IDN60HYdrG+ST8f3WqC2nb4tiix
NjL7ValUvQ4Tei516rpJz+oB1sa4rjqiLQ3Dp22OOzoyVFwpjQ4PvsABloPdkykN
RtXAQXXHUJ/j5Q+mUKg68Nm/W0d+rbu+4VqHmwJnJp7kuY/I7rh4b9cLvzJb2hrN
e5aHvwYmEZkmdkBNYTdSgmZhasat9wqWySPNnilm82GSo6Er7rRw3F9fVK68vsuJ
dVW+coSlIBcYK7Z1NSM3ZoxAPBPi9dVaTKnray1jn5K9DYP4xgbqziC1DGFzHRxF
rwClCAT+WHhD4Pqu40XFOG1Im6bTkGu0WO/y6GuOJO2Eg2OuVGDn35NUlLORZjH4
IDbiQyubknBc2snCLYLFBDXJgZH6MpRbprwZ1l2KOpgHtaQJZhcmfqbIz2CUQAmO
9kPoG79dXANnsMEeaoBLaomI99aErl2ipxJQnUXoy3ClpuxXRf/bNyIMTWZ7N95T
PeBU3NC8wTX/OpkVgQgAVTipUsI3WoexZ/dRWty5HGdyF4MzBZzVCaL+mIIhVGGB
lsJ+lNmrEzwsE8OzB/HFMJua2IPmJckbm1CVJ25hjIxF+X5aCdHiF6aUEmDAtx7J
SO0pEw3wgEW17gm+MshA9hfbbm86r2Ty9wJpFLHC+RgniIjUS1/bwrmsEGnYn39T
0ywDQjo+BoJD8DbGV4VfyE819YZjQG7Ncs+vuvD017m51x0rd6RLgdBPrQVWe57u
td/VowPWaYAFSVuqYvH04wd2R8bWIYjhg4f8Xxz+GX6IwHmatU9WhydsBieFsMqh
+2pIg0XqbrlH9Uxia9fCl6Pc9lAR0/df/GXi2vgULb9KDwXzxJfclQuYMrsD5DFU
/c3jKN6UV4nRDA/qHjcTD1Im9fh/FFqcmhstP8gtnvn5/n7uzy4cEq2z4LB9ILCE
A8opZLrbxzOUOk5kkgFMkb1+nQmrZSxiKSfhz/68tmZAua7CXeZNqlST+2yd3LhB
QdsrchC0ucvr9Kv0IMlFc6205NhjcQ2Q7/g5aKK2ZpDakVGPLUp1xAzjxovosfY/
KVsYalSYjjaJkDAv84FXc8qIV6b65bEIgcJmnX9lFnD9cCiNuyGRCaTT/R2c113s
+WsEDbUp/i1AnBKi1Keq52PUSz7KzWsonMzYGPtzDQ81jicUPpikWEaI7PifOZ7P
2+Qg0/jjRHlO6JN/319JK7IAGBwsVzlVCcGXm35sH6ijhQfFrTdVig/xT3Cze6QS
vpVwm/NF5mcW/ElqGvImVEf2+qJt7OFGGn77JG67VsViebRYebJE8sNtuH5LJOKN
gd694mO2jjgyieX2z/OufHrsAk9I6R01mC38KKjIm5cqJ2lcnJsp60Ajx9sYHz6I
NSzpn0l70Kys6rdpif07fJceVsiYLKo802ywxHMEKvEUk+RcTF7aBV1TGUio9Lkm
cKYApCWXYbgctL6VKLCzQ59zE0lzdmZ1KtlxUV7v84PEfo1gFqjes2D0vdFNS0RK
mgcWPPdQViGHy1j8/smLWXHkNHKzbwnlVfK0rUYR3M1bQ+6Owgu3sYgeToRzKhvQ
7p09LQSfePg+NLFVT254FrluNbWIDn9qmBacwselHvCDDxhA8dhNh1z+14BEj1Np
HQyl+YvX7dZGDD8XwvUsPDoWUhsWzNC/rZ7iLCQiyAEgeiPED1QC1lRyQq+/aOjI
5V9+cIXYZsyUP7UIEsL2hU8fSAKawTTcW7L6etjwIU7ehsQxacOWRF06rsIDxWz6
ZL/axsRjbS95Rnx5L+Ji17LJ5FVfa2PclqfbjOM684zCZB8E5BWrzu9hNZPKCMHq
OZehH8fA7a2d4zIt4l+G2KDp10vBf4j3VJqxCqOzBY7Ma74YGE1t7G9qAO610ISP
PGJ5dNuqL9AeE3Y5xxo1ChHpWBN9od65QnZ0v6SJg8pnCNONlYwAYe3D+60gNsHR
EAdQdQqn4iaAnJejfyMstRfuYoaNZhe/1eqCXjpiX92EC1Ynev31eIj66W6iDI5V
JNAuCpg6t4W5YYu7slCaL9knQgDznBMNJ97G1T7wscnOWhlKNhHCUW3AXKLnXNLw
XjLtYI+qtYx5gkybqfPXUppWmuD9d2hzYnzD9suXCnvWcAXUYsyRTmdPkt0VXyFH
X8ctJz7dFWORW/9sVW5egznUFS5n2jiFvLVBm0jmkueBt6SzucqCJM0VsZTRAILJ
s6TfoGJE/dQW+YuKel1WLg72kLcxEb57sFjdw5nPrLQSt6Bqq0cx7cXhLJOxTTGq
fv5vvO7hwyc84AGRy0J/4ONNx7rng5Tlc4N50PFfb2KAfa5O1T5Y+f1iFxVC8iFc
Gsyt1VLGj+zBGxNIOBAcUy98hwn3ajz7z4rOM9Zj5zMmVkNzvwYYVgD3eFRI/SQ6
kK8+j48g5pIFURCEWKro4bCTYcYM3LO6hLqpSvrDoMVEBi1wwdwhvnTXZHB1pz49
S9MMUdpObF3w1CVrQbV6YClIl8UUCjvfB3sLkCGl7/zwG5S6Q+TRP4/4owFMBSkU
JiMbgG6ktWIAb3XRoHeCgqNXzm943BOQrz9vSMkqHSfNrW6jEe/H1yKLCHx3x0JI
YT3WLdLcqTeWGPmEcGAnqdUieIF58j0TS9GArmvK2g6IFgBswqfHNCW77ofUrXHX
tYFpFC1982wgTboa6gnD+BJVaHMiFiUAmqHpA/ETjrDb6nHLWhbCND52YeBhAb0Q
Id/phld5OjE0JqbmTXaj3HNayvbhP2HZZmlXj3jO3/1ND/STUANiR9F9NGS67177
cBBIR3c09DQU2WisO065pOOv22YYwPEAYpeXqlsZHMe0JLJfX9bqDIZhqGN1FxaT
uRqyYIkx9HrGAf1m8t+BaNHC9iEtIzHOxCnCQzbLLlrJ4ZWTnrJvY+11/X8kb2+8
v+Fu6gGNH+wFcdjCT3X/QyM8j2Ac1XND59SHf/cqA1pe5mVzLEdmuUgIlGvLRKXw
qLrDC2zPawWQaif328hbEf1S/TbdhHsOH74WJ6wdWqnRuJOfG0HxGl9wnS7uOGNc
SaUk4ESftHHuuNtgmUOWIB+hG79yXejSVM3psgj3PenbTQsRJKe7Qdah0/0faMXn
QurSJlDTtYo9llwjQuxGBl2I9Nk8OS2PeMlaREaF08bX+51I9t3bGsBkhOFwPJxO
A+hqwvRSIxeF0+mvgrZsJ31QuK733s6kQ4Y/k3I3FRWD/MENk2v7kx9bfjshkGMR
MauA8FqKgIQTjXj0dU9i3SiG0nmmYwLR+Ev17PiViNonvN8+3yWkiMKZpi2iIspA
ypWOG2ykwn6VDdq2N9i38iE3U1IE9VZbucTQfOMYRDIwIk2mw8vXixjubJIU5qWQ
g0tuju8d0CG98C5vdargVOfdnC+VA5OWoCtb1EeFIcBXX+ewXAM6ukgUa23+HRIZ
xi3C4wRL6fDOlJO11Os0No/rtF3JxuZC7GKKHygHWf1IEb9gtJouh7QFrssIoa6a
0WSNnOzJ9KupRUVls9dI6HXY70SPfQKTiKrcZw08paHZSRpKEKuQbZBIF+BvBoN9
QHwfdcms7K6JdELf3i5bmjfSKjJgEAP5ilas/JE6ux7ZvGvM/JVjYqvcBOjpDYkf
jEJPa01x0kn+7ZGPOrXM1KESAfMVJwGpd/EUptdet2ECptqWN1rBwCb3typgaFCU
2LI9XZjD5IuFmfy4evUSVgexs0+cInv1ufLGWmcXXgkE54Bcfh0fM704vFkyrBdC
dPY/bVUyvrDZh3h7BADRFE5kBb3OccPdaocgzMBFsQ9V35xj1quAV928e6jITsOk
BC1tYSNTAaTPhxHucmyPdDqRkoWG6SWy2cGbZBzykxmDnOs+s9PnsN8zf/36oKoA
Z7NzO9G7qewA47c+NvI1KJqJoZh2SlYdwHzn0lI7hxz2gcjLlBlQryZN+nEM+7M2
dCh1O2Q7Fx90OV0Lq80nF22G1S1eDNQBBc6RhnDJiWW3EzccLpd7CqBMYA2wdIVn
7zrWoQuAqPsNkBzdeBnEXqn1JUBOCsXH5ryp3xf/uGLnKrCnovCXQqkrHYBCpBdu
CdJ+sMIPkVCfFTzP9bdCu8BUHbHYL5NoBswMVuptqHpFY2jFZ0zPPpskeHoIydiH
B5eNPBuDMdDcTfmnivcHUjP58J24CJgzOjOw4ITJJQ/OOqP/qBGxOWB7cO1b54AA
ZxN4EPJ0evgdme57n8mJRazMFliUH9ZP/TlKdhXB488zzlVNwPQOAnlwzbNS1trm
cvv6S7dx3w59mi7X9pMgbbEoEqlxuSj6Czr1XgTIKhqcTz0IwlHe/IzR+/fq0yRj
UtQYRvKCZbQXT7yqRMlqz5BQLt6HTRPFvsg5h9BL4hk+npNdBqfJhbcGT1CN4suL
3H111ePp0w5O5gx5rx2ZPZ3Eip2rsdPWe2V1E4oa6quUNPujiu5PQe0yGGUiYM2A
rkU5JYS1bmC9VTzdUbRTXf3DzGFResTwVhRQ8kvsS3ZIgFMlzE+ItHy/M+oKjMH+
TiBLufHmQPKoaI7eH9YnZK72MGbPKF1iuvwUMxvAn3NwMKxJwmwX6a4+waD5ZpWy
j49EtRPdHg2QOnMpmmJ2axxyJ/Txje0Oi3WWanStgP/pfAnlS4Nwy4pxFP2gZk5r
EBHtXRkG17UP6Kz+Cchf490U3ulpf1najv3O1Xg1/uEylIrA+3Dvk3wuoiwCiOcW
gJOmaV+kBzLh2xGXIuYLkfdnAP6QxTzNMwJPwBP3RZSFWqV64R+aLL5SJSd1su5g
MNOoXDAsOy9YlB/cSVFkJBV3N8ThKCFRTkVzkUi+SnuyV8GgWrJ7eL8OCcWc507K
7YRnwrulXE53lJSucjUEWBK8WtktQQz8EwhzIZGGma8hf8DmEG2qjZG9jcnn77tM
kKKyPLtXdIW3mmevVOnAJnQ36Z78g6Aq66SE092hlaDDc28eWsanRCXKS901NKYx
aYFY8BaCNLBlKXzT33QB8Hjzu8ZIcIxumWNOKmI4qwGGPvhTCTl+Ym+7aTv79IRv
PxBVDIsYXCDi0hjwUdgPqzWAVGofEgUc5WAGXoksL29MLyFltjeYvAib67mhMyUa
OmNvpFGO2ipeErtMiEZ2VU6SaX6FYTrsJRg8Znf47EE9lEpQW4TGh3TBGaMt0eAd
ThEk7j5Ug7QXaOignbEZ74Ii71NuQ3kFHEhoiWP3tEVvKxiUHFU5KAh4hkj+eLya
6+UtUXAj/J+AGERFcXVvh4XuNQJiyTRxfNdfQj6+rOb5sBGEsNC6PT1JOZ5Y6G78
zPcgQVh8HtEog32WaknUWbv627I+XkYW844wFouMk55GJ72D2iWYIapySUY4gi5F
OaHYcEttpIw6/042hYDDzadCMt8n/llsS4iEhDQdkBZ1NwaB/1l6Wo6M+wMH5U0X
o7Wht5ESQ5xquZluNgRxhlKJ40yM6aY1o3a8U0b7X+e9CqJ60r5IqobpIyyealpP
7tCnHA0bdPd+S8yUS/1rW6LTyRiaikLJz2OyHSRDEGkgEDZrWkcXz/bsE49Z5iC7
HGG1aIEB/vbBd+7/Db5yuFYOQ7lz0qjfGnzv/ryBnPvXj9UtB302banp0nmxrnf3
NSduHLIkoS9Py+1+kFoTg2GPNS7u5GKhsDSTYEGXKruhKCHu57yl7n5cY5MeNZqv
LqPNjwl1Nsy39KoAoDmmR7cEJ/MmvfAdVzGKCShBJrtupeL9dLQVnC63FVKj7t0F
8foLxE8O25naR+5SfajulvoVdo65B87DrJ8b7pofRS5yB48ez6vSKDVqTcRa0HN5
guibB/Zzewkls3NzX8tI/F4Drtjf97/NDDS8dMb4b+JKh4yIclndPwzIcDa+rROR
a8qcBf53YwdI2a3M0X81zRsT4Sw1hjlyj2g3Ohm5EFZ/WkjzTWaJY1KqziU1Z3fb
pUfVzb9vJOvOEyLpR/Rhk+BlDJRZ5WhACAsQNF5MMWuu3LjCxvelAW81DH6u7NfG
U4YT/3Qmn69BNb+vRPkJ0QGnlt99+Hkcq/zC1XqPq9OyR2LcLADrorI1xcCc0qOc
rRuqxpZLxWUX/Emtcu/QD6juf3Jc+jAvRArsr6OTsjhYtHe0K3vuwZHyax6/ZKma
6jmaYjkv6VpxGu9+Or+slOYk8WnNFSmMUaI5q4Flx3ldAouRYh5FKP9NffUjnFDU
0tymSOCtZbUrYnPYb5LrJNKcE9XsNzYiVVqk47Xjr0rJXvtkFfuRj9Ly3kAOMyZF
qwgdQKwjFbdpqgoW9mUzoLF8+1vfeWJJma+BP4Do+2I2RNe9XFJwCK5i/JVUQ5oe
smqxTMKdvR1PdgKCbdzy+fDh0XOWFEWK3IuvI6Spoe7bQo9BeHNjYFzoFdKgZrEm
+cy31PuOpvnTGLNci4S3cSKmAraPjlIM8w7FPTvP4MY37H/jgfcJwgnrUvIs5iZ/
iikYP+rasL8+ppth7of0cw6n/LmffiO1gEIrsmdDLC3S0s7WrreP/ezkOyQgXmQY
G1GG15l+PjRTV7R+PkL1CgbM5zgPDnRjfm1gAUsNQ54MYrJHY/6qXXSIhHN/fQ6D
CJMItTUy6Q7hMJdRKFumEGkozPBToCunngnYIjC3WvByA+1Xl5bS7aAw7Tbe2X3R
Nlf+joWBrQQH0o8oaNikUcBx/G1FBuJoncVQjXNmdWjiREqVQ1DqzhI/lYW49B2A
CNvZWbX4ybhKW7cX5akK8vlPAwFB33UGxQqAiM6VfYzijuG7q9IZuEdWSpwf/odp
6PXHL3tinuL+PWRW52imTOepSDTnEJPlluZKBETAevWQftocdth/8y/K4/ljUWA9
TLjkGoGt6MM19byB2VRkYyQlKbMCVvBGajI7ZZ49b1LGXY26NhV+k4pHESKxS1Ea
5e31L5fNW+39C6YPOtT5vK266t8uCK6AKsn98ZGElWudtkooawJNnWQf03faGMLW
4AwKLLUMimEjbw9eeimL8QiQpFafuopGGvuovggAmyCT0xFqpCtR9xMCJSx5PjJo
xHEWRBBvOqtuSXyOvVAAb6fQSwOWMovbhQIw3s61eAol7Jprtcr4g96tRQbBV98w
5QdkOjlKoYaenNaFkAZx9+wP4EKTH+jYrEJMJaKQFrBNedxLjpDQYM+pr+iVamzA
91BS5nYasIw1VRTXkEAvF14kZYb5RuhIQawIWa+ZP9F/oxEZFgH7o/0PvXVTPTEf
nE4oVRVJNmIa6JM9wrs9BXD1fEuL1Qzl6xb0DFJPfTrJ6hPeFxvWY2yGhqoFaop6
u1GazVjOAFcXoqZn48nBF/0mjH4BVtLk53DYIlXeD6PeW/WT0w9aa0eZuD4DYCMO
FzpmTUmAGCwa0bkFnq41TsV35S7uzwW9C203YRosa03fvdRul+qK50EQNOr4gsN8
getGip2bmmHD8Zrgh3WiztOElpfKIZhfo3e6Ca6BFe2Gp7KVVk41HfTLgT74O0PP
qbTMRwA8Yj02rI1j+hDcsoVwZEPie2Y7QgXaMt1KBqrBXbkED5MwFqds46M6qfYE
L9CM6gizByKpIQOAkS7S5BbuyKWrIJ5zk4NsJZ12DQYw/iywEQGqnH9QgUtR6xUT
uFSxX3xYAjH/7mXz3CN9CP0TeNcmETXbzxTCYV5xzpEUGdrYD9dqDGnkc92hrP1j
6a/SWg2U3HXxf+y/CcRvMcBikAr7Ep7UegMDRzY85kCmPxgOTxfGiAkye6MnJxKZ
0R7le9c/Uk8FWut3sHjJUIx3bM2AWVkrGI6x7tTEUKqQfH4dOembzr4wxV68O3CF
4YYF+/5EhwYPzr/Gaqf1mLxLW4Nka3FjuO+hkpaYnL4og3pNXadU7+NugDe4DyEO
qlhV6wQEaQRr7HaBuompdUtpp9UYkJKKFfMtnacLp+4P3Aa73zPrwtp3YdgE6BiP
Y6GT9rEoam8eFlht6+pgeDWB404ZtfFp7JjMb7RG9+EUnaWuMBohMQhCMn6X/Tn6
jsP65gu0u9PjM493SFWeJw1l/5iSfPdh5qROWxWlhG+jXWVZkexIpdnQJtFZC2ft
q1iUn+qKCvtoG6Nt9jVvYJjyaDD0Zu9mpISZ4EoJbs04BQygJgcOJk3eWkO5pZps
asLo557uvdGxJxKvzUaFI7Qn+KlZhXSgRPcr3e/RWelQFvEZ0Lu/rKnCJL0ZfSyu
+b++5euL2ouzmYIkJuu6vs0c/R/yFRC2+JUTjMy18V07wPtM9dN07AHI7ClZyLdc
MB+y0aculYrv3fckUX0Xnu/FCrx0/hHbPKCXo7YGQMfS4X7xnNW6moluebQXrj76
Gg6cvgbwbCBjZWh1VnE27hVmRvfaAkoRZh/wxG7668YczApzjgDqgjf3LVbOlRQH
Gudw2G/VqRVb2pgmhV13KD7GPJH5s+M6JaveYgGF7xMmhYoBnl+vNU6YioJhqeHF
hy4WiJSrO34MVg8zgw1jjWCZwE5W2O4YTomi69weZrHL65l3RfkBQQhIkpZsjn1I
a8vgIRkoBJhp8wSltMIu+HbatJwOfMJyJ/0ChcFLtJec3JWdSCuZd5+xHilSuqM4
RIYqCV+mvzG3k0wgMiIJ8mFgIVvp4WBtW8KET+7HjuQlAEwfFFBbmKc0kwmz3D/5
9h0//PIKbWtkCO4/2O7XDxzZvLSIR0/IbRnFYeNWjO5+rff3LEpGoU0wgsqU83kz
jUvH9D6SvlW3tBPIEoX8WU9sj0BffeJegQp7Cw8IGhj8gg3wjcBub7l9M9z48D+k
QrVUkzdMi3ikL/Mm4a5eIHoKoNy9G4VUoqAeC64hSBqtvWEC6ZYHZg/c1STNlJkN
wjfGa7PlW53vQx9u7AKEqCU86I8trqICLWuvx6U1cl0Sv7wtgEII6sy4uSGVm54X
nbnOdMC503pYTjbGIqgUAj1/7eyfJotLUzbBPMmNYIGFKXV95eJxzbP/gwcgm220
aw+X7yK4opM5yqrIAbj6Scy3yY26ydL48hd4nvYeeC9tZK3npIMxd4UortydElHs
d0RIQ1IwGXHEI6Mo/cirjdLY+j/ykuPZjTpn7KS3qvHyvIB/L9vlhG5U5UQxOVWA
BWB6eEVPZjxg0ouzIdA0lWZr8WfcX8CRa8OMTnbX/bzslC7BBOMg8mn3rOAf9qZl
8A8Ofg1l5qHw5NsswOOw3Fn31GBK3E+IBIEyeDVcQoFCWgCgoUfCTYVEDRf3t+mC
bGSgel1b0YJ7y1YpkQ3FPHXVwZf1gEt+kJnh8iuE7BUShrYO4q6DYbyQb3Z5qeVN
MV7oeL5RWEh3GIjU1y0J86ZJg3AsNhOJ95GbcDY9y9lBFAGThCiSkkAK9AkjfRi3
hjrhYA0M6BF52aL4wuWXocdOl4vNnrRv2A/NMDi+yAreuhvLEY8eyxc+EV4kK3IF
xYNCIMV0b6lZTMxK12WvbkIuXRBuoK4bxR3B3cPhdY1aJ9ohJwl0ck4oxVYOQOtz
MqCGEP9vLw/TMQVZg26I05OELB990NWgsIPWUNhkQZ9txSnC8HB4l5A39MvjfVz/
NhT20v6FG4BI8Jg8WtRV0l+7AiP1FjCtKB+Jv20kMoPn7Rg2rrjqEZdan1TwgnV2
tksuO+6fhZCivnoz6HmsuIammN1APEFGAtAV4a4C1MMlXeyfnMylZaWqbMXPBw4U
KKBYyVFYahsYMlncub7+cAB9u9U88NJgB+pmrDuz0uLNJ6ovr/0MUkKaJv567kFR
1r7Pwr/3dKMQpmDEq8fWwsahH06iULNDMUrplvfbLies2e1zFLwzbUGxF6T0ijPO
u27X3hpgd+U/JjSRMa1Q74lu+GmSLihU7KKz7QQwzwdKdmudmxaxlqQ2IGkbu8w4
G1WV4oBq5/SDESAi1LcB5CAw3xExAEbnNnYAhX5gjsAghEEA2VNbrGsX8a4eJ2QO
1G5i+okwvIKx7sKhqCVz5mJppmDhOEoor9y8wJYcKEQOu5hJEauUXo+nK7BJ+ehS
tRdwMI7xuIGuyAe8MCQTIZkm75ynDjkbNbw+Juy4QPGpmt/PzQMj7cm0/Wlh07RS
URbDbDrvGM3KicJaYBzTc5aaOOP3EgfFv7OMYapiE5WVmCWnStEcvcNPyM5ZQU0s
c9JBny+JXccCEbP4A1ee6fVH64tG9MOOr6egM0jqeKRevOS2SVKonIuFAn7w6SuQ
Zotd/ctcL30Rb5gEyXrHnzDaft+u7gQp9bhR+gkFUP8ELAYYwE/be0QHdecnoRj2
DcqRM6mtDmLUugPCNJAO7phziIaaVzYE9fuCBfy/dKR2CTtSG40h2rlBoHEuTOx8
siTrgm/nydPnSUcbXWMOBGhwUYG88N/S7RMwRiiWHMIzxQ1z21VwBRcwntBUdfSf
MBAOR+XGdjk6xS88SrZ+kBaBST4z7RiOJgbi+qI6mVxNOir0s6n/JB/StRGipynl
1cpP3a5OLJ3nSlEwf7PrNmy7E/Cz7FvoBAlt5kSyLN44TipiISS5G7AC4RA2PvEV
1tWFOl6wDMVjmut8zMP/tBXC2hM14ZQCpCwPPP2QCc9pl4v7BzErCFEpRe6n5qb7
iM61Re0HPbpQLQ7sGlwWa00XjpUMzYKLS9/pyhXwAr8Py1bA3QJf4D8VHspYdbmL
gyNcXA9kjE7DsfhNQTKR0lBuOMWukaEu2IMo5dLvybl4scItrLrK7VNnqyTbTehn
IjAYDx/xvedVMTHTzo/kNn4m4AEPU6tTfEuOpjq1Q4OYMHiyyFmaq+3R2LJ0HmJw
qPVbfyKUBPsIi+RS5VluSsJliZeTcKcozFNyimfTyE7DCDR95E4hXpuR+cgyDOl0
mqPt57PaV0SU2p8IVc+TOhJ0gTWKeWnaUH80UEbpiACrp3H2V5DYW8C1/YyPODhn
R6RncNqwCFPDePa6/EWoFpaAcc9NhFiDZO/FMozGWlAN5PoUP28BHOE02xwYtGHZ
VXZ+RxAsdax+Jpd1fjpod5Kp1m2B5EzPz/skSk7M+LqviMw7DD26l/udvE9UW7HL
28k00pkqHMA4eT5ET/wUIeBLR1XpCRNjBqOxLx9CyHnr96oh+lZmcg5hSWW2Seyn
8vFyQE6t1IwIn3yqEzLdqFuvvsTn2yFfHVWeg2PYjfUfiJ6+YmMCY81Bejn1E8Yp
+rp2HwPnOxUva9g7BdEUdgxiCb0QvHHTkGMgJWrxxCzunGWD+wtYrG7dJrsqPli+
43+hdsJCqGhsBAndOjB4sQ7OTEVd7r1tQ6/XRtIKI+xqiSCtJC9JtEU//fQTEviA
VyFe2lb6aW98ng2nmDK7KFkmaJuv2DGiUjVLlGv57B6oC56FmrzoZMuppn/v315B
+wjbJmccqf97C1KMsmeTFTK6UyIungUNxyIyzbqtNAhdMq9+bODpAYAMXq843C5+
TsLDO94ARjC4fl1p05A5oJ1CLLnsQih7N0nlBW1yPY2vvl3jFTzWchAjXJ9BQxqR
1umOu86B+rq03edjNocThRtyfaivCYuL+Qj7HABDPtZt3qgOlYlOfCOPrUCHT44X
+ekxbhObKXA1ggi83b0xuSDMComxrhioDnzSt/O2yYJoVhFnzRxiQazqNDN3rSAR
vt8QNOSWMMRplvcjrPUb8okGO6e4cFf6WbCJDV3QYNRvGA9ItcEHUfreWZzyeKvC
3SYo8M22VKnAu9RJaqqcpak5m1ZMAQOSqfJkhcJKvGfTYIbgAegxChhKGQepyGYd
6bE4m/+vHaew1UVAzWPdFmLHVOf+cCuy1ReTf5I08RLokEtpXP/7Mi5qGXWB36rz
2aGkil9fPhao0KbsGZ8Je8Tyc/2DGE6fCfqETXGrlnOnqF2jq0KHLuxfv2V21P0d
mrRyrjANz1gj78RdoPQ6HxMvfv7+xmXOzc2aFACuFQArjeTKxDFa61ul13vRqdV8
CqxWga4fGUiFYzPZG8f7gKAK9qhUoKqOi/7DJ1mTMdP3C5wOxElApHL1VNY+8Q4Z
EdHjE0fLk3rBMNsgZzivkUSIamQgY/37TYmI4JjGyZQTRVMJOgvMec8HgTIy9r2c
MWfx93npn3M/A6+rPhKLEG54m0/1KVIDlwBMdzt0I8r1l1VEEkQ0fn9vG2BkoMYZ
/H/Ceft3hTJrKfvytJ0eyg==
`protect END_PROTECTED
