`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uWkPzmYIcrCjTAOChMcr67zCwQYbw1g4Avesd6eGNn2efvpsFmECKIr+DG8j1gmz
8JBZNI8Iau+87/CdnCvofJYYWit1d3AXcQkR4OAYBhLy2Ve3qRCKELl3qPdfiEVV
HxZoHdku0qRsj0ys+nEri1tznSAVac4lVmXO+TDb0l+Fx+LDLgDXbAKJVqgmEU0I
QH/59m3T0A5d3IafWMqYrDdYl10idzw0F3kx2slQG6sX0msYOrtj8NDmCirJ/5r8
O1jE9ZrDKj3Ays62JCOM11ikBsq6jFTXxujTlqEumMhF3g2iClIEFKgklXU0UObN
O6cy2Qg+XD+stNO88cL1Ka7DCH2W3+qxKd/+QhY44HTFN1wKJjdhPME8wbx++q3y
GjmJYOIimJiHt5SC8cNWH1XW1tmyK5bt6zMMNljFo2a+dnFRueYgNN2EpBJCtjji
KUNvQS+iCw8uwdWsXEPGLFWorMCK2O+D5vA+PLjnG7RxKB4lvBaFcQoxNuN2MRWq
9JgZjfY2WXkdG6pPQenKn9Kj/FK5i0SF/1+6pL9i8hncEEs97o2MB63ISDBueQp3
oZSfZqAhxaUGO2/wWIjpuep90Ve7OgFCBh8w1gG+xkHfkjSBg5w8Y75ueqMxRuXk
EjzxtqrCfHN31WKw7hBdH0fjS5GUg79Bl9yu8ItRp2MwoyAb6WpOMmogya1682Te
/UbY7qTnzo1JDm6SZqagT9hURdEekXvrTtlAn4SYTa9QjrjxfQAPKyMUsZfXBY7G
EokfAUUrZVL8mvcEnPsUIzFA9YCJlS3eiDtpWVr6+KRC4KhgTD6jBiHX3bfoAkah
v2w9gstoXp/q8duT4AwfS/eUKSNjdO7CHm+vBLY+jpEBqNmPd4PJp243UtBVPLxU
whipWk+HMb+1nkJFYPiKHZPeQ0/bRHbPACwsiLkLWN+RlvgYvLX2uAaH0r5JUuEC
4IKihyC7C6d8cNq2KWcv8yJrLbs1cyJQuWDgkijrK57FGQAISmK1Mbbd+ZRfKNRJ
H+c2Oyzmp/YFU4T8b0IoemlGWN2Lbl/5Tu3wCVDY1TPXVdFjCBJ5Ey5buxSkgnet
/v3KsWpMpJ5/PsH12Ckf+Yno0H3Flc6tjW2rHC9N+U1bo7mduh5t+Bg/9AJ0e9A4
gFjXjLCtPlA7vheDA0JkxMo9RMljco5mcHV9O2MP29Y345Qjj0bwVR93O/Tz8Vpa
BSW4wz80jwGuRPA6WlX4pShhmTpG3Eg0hb3hKM6ZgF9/O5f+A1M1v0GIY2OD6To2
zOiNhsJI17IJalk319wKFBtg2ru/iXk16sRmP6KXK6wCiO+Tj/AmethzMgylbTRC
wA33sgbjLv2fOI+ox2kQbCDcNhESf3Wuu1ITc8qID48=
`protect END_PROTECTED
