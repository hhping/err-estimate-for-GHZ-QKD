`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RRT+wddGAf9/qEo5O5aLQUUKwXC3XMTAZIOhutHoeiLuj9u2JOTPCB4ygPt9l//7
VqgdIT+c7SiD5sI/8TosC72puB0VxP3+h8LCqK2bioI10zXYOT7KbN/OG/KxM2Nd
YNWtqfKq/9Rn+S6FQ8oN4wMWBVyzLVnrrWmzJ0xhvGw4BE/+Zfv5BUwUbp0cIRfo
JpTyqSsxropJlkOypfTemZ61v9pKWc0iROW+L4vK4keqZwkm6Qlyp1l+JoNtpmy7
xDzdtwsrQfSly3a4YzyCGjXSmETYOsQTkHDZYNnSZG8pfw6d2q767l3f0dTXnkFl
V7BRToX3J2uK8HigJ+wwhoJcPz4bob2ig1fy2U85D6eBtEO3ofIGR809ebPB4l6t
MwYOl9yOozpRieBm8UN2OiQCM8fOKD12rO334W19j6EEq3DBm6GVBmYPbqSZ2Q6s
eRVSCuin65CyAi/YU+5iJJ9TPrt8evgD4nXhbuuorBZquYVxX/FBHA/shEpIjd9z
XqZWBdoF+63Iml1YV0AaUeBPr367l4v0CEnwmag++QYYgC+6pF8fOCQs9hJpiKJ8
OLTLRJu3Z12lGvZgBKcxJLz//Peru4lWAjqsM5epMQrzZozOtww4LwMmGa9kpxVf
+qUmSEI8HZkXSvTxpv6zcGQ7+qWM56250FniZ4pwGRpQubjnDjZGsTe8/Kf8oZ/T
MjTYW/yTSITW4TNzCivu6k2Xq5J6N2nHY26FGkoj54rMLOnC63QNeCBXCjjt7m2J
MTbYkbx14s+d709oVY6b0jwHPzjj1wqigGN+iL02T/vEnPjavSuvZdwFXLgHxoY6
D0kKXVTv31LfyUld1cYLXv7fXP2g8rY661lyXG7QiBfj67x1gx1TIdkWRtzUkEK1
PQY3aMUKqTJJbmjfFNscund+VVj/10UoX2x+SxMEY9VX/CVlplcEn8YyUnFxJSl3
mf+Uk6Rk01ZAV/gnKCcStXYuq3s/VbDSJKiPekZci0B1uWA9HhkVLBzk0I8wtqFu
mSqiMKYy3wVyl6/UMDzSndiwGgpUBXMZDD2cLwoyRBBjXPE0ThOrAI1taVjE+EwN
yLmxh/DKzuU9A47C1/LqVcvKj8eZtez3Pt5ranI10gSCSbTPkyeP17hz0bbzWXoe
KuV9yu6ISPrWInnqTQpdWR4KVhK9GMkOgKMYvTLRWQcuhlAj9Pgrdoj5bJ+K8n4v
FNd+BoN60jkKbwvCsBME6VlzRH0NzZMCT7T/uv7Jbb6jX/SB/dbPF7NVprJG8SoR
2bNuq1pFLWhe19k0JQLIYTpsA78DXKhVlSAl8q8m0vgqvLVUzUTmqYt0U4uvoltX
sDVVw/sHO1Cze3j8l1NBew1vkYaRptADJE+2VfEegIWHuA2px0EwHmxbkGbeL0oi
UnH3vKt5w4jQ4CsLj9IthQhU74HPxeVKBvSrLixFVnhaZfWrIKj2HqTaxhRuWVhk
nZLQdainRHeqHj1ow1g6DHiP//s7q1RvUEino+Dup5lvHOinEgtvx7Stg3AtDHH7
an3RDLvqNZXIVYZE4I2K64fZGW8oCXbBz6fsrCuLtjVD4OCQ3wIWFSNNxSXGKt/Q
gEioW272zUYCPRjZxWajPw/QX/fLyeAE91D7lMr5rK/Ym5n3tbOOuLSYyUY9AZdo
8G73EtNVgVo8bPZj5Pg4FzMY2TTIMoalmDOdxpkG+vw=
`protect END_PROTECTED
