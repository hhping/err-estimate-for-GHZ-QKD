`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OeV0WAN+Y6yhGZo2UMyRHmoKF2euZos04sI4FSw9mu9/0huYXsUhMpezUAVRjGjR
IK595m2k81Ru5w6Dp0WyWmt5rlejJGgIvwd19bMP8K3XdK3+iU5LjzO5XeZYkgK1
X3TRriXbuMWIncofBdeUaGsPEfMBAw8AmI7hOZZu22idKnOJl3yc96V0FV030CJA
OkMrTgisMooMJUUH74I+x3+7KDN0FCwYBIViScM5oBgXpK12vmNEqV9Izbseo/6R
MGMQEYG3A26NjYhRBynfSxNzUUYm3eEzXo6FpMdyhYFGAL343zPe8C7ho19sAxu/
OOrg20LD7HONeU0gFgxHiqjN5AuK/laW80xkQbkhOjEAkaGsLwGIEEMu+eSncHOe
+01bhS4xcp9HAO5VEaRjmcyFTosayE2gubxgTmJfDEl0kVr/1DIyJ747VaclXeFj
T+PSsa5pQRocVc/Ov7P/2QYNa2mX7lkY8wxyaJJDQnhI76ztXkU8QVwPVKZhM6S/
pDodB6VK9VcnPV+b+LC46er2PkRRnFMDoGFESc8nUmIvQZrLL86mIN107YIqBJ/K
7ob6+upztAIwCij9G/EMiVKFzCS7MfYn4Q26/VPI25/WZRj+elQErBP07Q43N5xC
1f5ssyPbI42n9uDwLEFqREZDcTkFkPrQ7EvytsQiNqKRO7VeZbsnjuEdFs/mLQpK
rqoNrxQGj6uos2NNeVB3qrkcoT9GMnIzDThVG4Yd5So3v1c+PCAlmkv5vW6D4uSQ
bfz5JP7iAk+6plG5vgi+W0KeNEgJzy4aot285xuSNs/T/Iidb/f7qGJYZF5uWnUC
nlgOiAg3lNrZHCArzXMXc2eNND97bVRQJRtIA79RoGHVLUCHosl2mkYaRecwiExQ
YIG7wSws2FRT12+x3BaQDdwX4OmRSL+MkrclgChGLuer6lwT8E3qVKDcT1oqtWum
F3T5LQqdYLFsZlRirv+i6TgLP/pNLVyQ67gH/sq1yt/An7c52/ho1hDwKJVmk3nW
e/1kXH3xVzL6uqohJEMdoAS8esnTpBleMJ2GXqOfF6yrn3cVbm0dg+zYvgjR9870
akk3eW1zsHdoOv7a7n5KiuKq0lJIJoSHicGP3P+3gTkXNz9+lu7IxMJhPiZ1juze
PQ6A3S1FBUdCbSCif6yzIe+99PTswzs4BaY79nqi+fDDDLTjtV2aOuorPIzFUJEu
8wabmv1sp8Xm3DR668+rlE4oCRXT/mctkfdXlXWwY+Py/cTrYsfl2ImExR/yyiTG
+4hfIE5gnVjm8hn5Hs4sXdrVENJCEYmCN4oNCjEWIqpiVTN0vgP8ge8tI4YNsI8M
HtaGzFseO9Z00sdHSaGtsJ96dBW8v9ZiyUSekRGPe4NAQWB6LEyviu/i98OXyXYK
b9F7xxMvg2W5rV6QqwB5KZCIrcRdijP7LlKR0BhHs9Utvn9GFLgcJpjJvMI3TJB5
VN7ef8Ij09jficWo3e0+yNUDSMVSTvKU57Kdj6ekaQUWV9RCcGqnQQvtztl/aXmK
vDJNTsuwNcTGLcEWY4LVKPpWNUVSoeZG42Luyb2LeAabhMmAK2JUKjPixaaScayy
3Enxc7LjAhrsS7C25GGlk3akFMnmzqnlszwa9HPUNzfbfD7TZKMyCQfvplRn2wzC
bDa4+6E38Se5KRq+IggtdGqv2bkELuKR3RqqJOM3oCohUtIlwFM8yGX8hSF90+t7
bwBxLpUo381moGG7pkAHiXblWWgOJjqipOAOOFC0pMBNRLLphhljNjFlOhLoqqZW
Go6Jf5GXWSVJ5nm12mfQ+srv+uvTLUkltcqe6y3ez1rOFTgUQp5RAdcMWZowqEoW
byHEyUpk+LSKavPDYOu0+sCHHPBn4ZvE6D/g2BEqMw0GgZD8aSNgxG7kCbq4sIBa
QPKkpnbmgT86d+O7sF22q05JuZiRDfuElYAT+TrxzWtK2xNgWeZ1Fd76L5OOvjUN
ogk1XpPF3pvISghL0tk8qysJgmsNPKAtK55rMyqxDeA94Hqc1T39GWqgFuwvR9iM
eHvRAsQWfYkH+vKWpO/9oTAZtNntoHeDfkV+SgxAWLsC5JcrlaG5dHayVe+WyCC9
K42U+DVNJzwosumPRmXQlXPQf+AKmX4m5WH44EMQ3iMRZml9pCw9t491I0Jru8Rc
IfPF9kNM8pvrHqkWccu1qCMFWwnNQvz8HgMHve/FWCHSBhjHTA7JZLV6cuJAk9kq
LyqNDpeG3Zto0boIMxe0ZjO+xWnfj+L5mOieuEc+aFjZYx+eBnHl3Mk3m559pq//
kYBJeD3pbOikfoHpiigOeTjWw14lcFsSchZhvAJPYGq9XTVNQpN3TAK2X28o0C5l
/c7iUKtF2xyp7yvrbfgm0N4W2PTlbdRk0vNT/tNRRkL2AljbiB+PhK4ef8Iu9GTI
0l3akukSQslbsa6lAmpxH+5kvhMGFhTr9MOj3vRvY+xmJdeQs1mBEux6tY6wo+gG
c/BdW0p2nFA1ptb0isXjG2szHNX4Eh61sXA1EnO2Ep89M5vaz2cCx5dRyYCkILkd
XYi4z69ZyBrVQlH3U4/ruSPITBtqYwuC2REVJ6r7tiNs22ACSQItDZLh2Zu7UGO4
U5/djnDRBm3u03wzze0rSrJ5s8rRsgvnJ9wntWXeuHTf3Xkbg5Vnj4QBj9Pfi1rd
kgybQ1uxeqZCYqhiyec7uF+o7xvuCfuU9RAaQ6fn87yGGAUHujdx3mk/FeHfY53V
9uqD7Motrzucdb69n1uWx64jSbcRYixDdIpf9JlZGiZPp4fFjQa0QPy361rg/cNn
eg/ohFBzdQR7pQK1gkCk6BA0piReTwru1sbWanMYurOm04pT4U6KUgX6d9sgVUU1
WYu5P2TH9GpYSHiylu7fdpWrE/+3hCgwSiXdcFRnpug4EqSLBSg4F7/twY1pNc/i
stTbjy5Mnh0Knu+FHu2+iEe+LTyvbbr/ZrxmgA1DMLE7IUAu4jd+LK66gKbe+48A
ZCa9DR6g8+sdtf6yQa4jZ1MidLJz/8+eLMYRZsAqXycjsuaQmtt8dkxwe81OIbbo
KunsVaLIZZUoS8BBAngqq5myFJ5aWLZja2khKD2M+g588UD4f+376USTe5KWW/sb
qlevRy7jDrEYxsF/yc1ecvJrR4EQ8k/8A+zNwb4OF+cBaOODnADdf47rgS9GBonB
dcxk4XCgUM4g2RKxIWiry+c4GUfCA8+buGNWUKy8gZ+Dx4TgvJW50H7UyAJImIeM
QffiFIu/jaWfN1WnI6GEp7rj2t3P5EOzyPu/JbLeGD72UrzJhFr729y2Imz4Mkzq
btnp1oZpUco3E5sCWTEyjRh5gD69FPUGziMd7qBKWAImsiE0bbtbXQjsDbmk7ehs
WiOk4gBVakiEE1iySU6EZTfLGctK6Q7yctIpmvvuh5Ym6n6fDuYXA+xyhEFRqlT3
KASwrMI0N+5QxXHoV7jXAMPSY5aqFNs1on9ij5xZc+bXvhnzHezfZMxug41B2ofA
bP4WckcMzl9NmokczN4k9out38sA3qi4LWG87hCI+MBhyWfbuJ88zLQO12TXm30e
/EZLzBqrKn46TSB85bXZU/vKavDx3HYrinRxC8ocnuVd9KJfDdkdE6DASo7qanth
9WHYrxhEo39oRq0alIvtCXjkyawn0N4UfTbPperdqqtMHGjUReJQkZOnZKho7SIO
FYL52rxqmgZ60j+cqmd4cVYetyqE3RJoJTjGgBic7U6L5ZOOjIbxudfuvgz6q6x2
pophvy9OetQ5IktK0lbFWdI5C2XP8bBvoPi2FByjB7XH0InVs+L0vYxDIysRNZO+
uC11Z3TigeGuAgnmI9lSAkIFCiyqUJSols0FZ0AEY7B9XFRBruiou+jnvZmpNa0f
Fmje+on5gsxTWjXTwO7RoV6qc6NLHw4LCgjzl0/ZMgby4r58qQK0C7NWUtc8NPXm
YtnxOa+krboyDjM/0XMaaSzJWL1ly4LXrbdae/qC1YiCbb/t/VghUaCDcX7zFgTM
CLgYRR2N0ON7I9GHO+sigvURDi5n70S0cnyucZKz5Ob7VE7dcMWzmOPBhG104vBx
6IzkRzK1Nawx7hqFKNI/HIKeJxOc8Vg2eERo61fBjvhg7OVkRb+Yc5H3DxOwMdlf
KiGyKKIr1cQp1ttERyLFtej5TWghzLR+MpEqRsE6cES0tfPoJ+rbntcbbqRR907Z
sFhlJtPUA1DNv885Quh2g6PxVxEFnEzaW+GUkUtCRp/OK+mHK8gXo6qluQmZ5BBN
YNBGt1lwEB9Emt7dwPrrF1PjmTd0f+8pzeq/nfp4oIzloggyeHlTNfLLb07K2feb
NIAiqAf0rSh8RlhX7fc9vdnaNT5Ced08z+6aF2yBT/U76gCoZFp1iR6pRgUNjszO
73sJdUaVA5faONNp0C4GqplBrLW0tadhhOC44hmdezfTmIoB+cePGsv4M0LVsstP
3TcwY0/yXQmBpjYtvQzVDTo/H0Ew+c/vxoVR3LGadvqE53JCi9qbK7R32SCpkzOy
4Jqx6bFTEYX2aHQiF5H+H5sPb+Pxx/k2WlSEbTDb0Hzw0pXEJZCqbzGD27SrAwt3
GXGuJeoHQiRppS+2/x+RmSXQHMED1ztk2IhownFsej2QaspKLtuWrf4Hj8C8O2b2
tFz3N8V0bALRZGHWrhubohR4SyHlJnXZlavXA+wt41GyiJc9Hb2YoUlCIW1adS7e
jTgAea8UizxdPXbcQQOypo80GcFthLcWgabFMtr4KBAAXoyMdjmsXFF5NrCrerPx
MsNIDwBxE9/tcKb5Z60kF+aHexXJYwE+Kyced5FFVugqG83vvpiMcHUjuR/qtBsz
+XFZHLE9/jJw7s9gcr/4YcGxyXxCJ/WyB/lwGwtDwk9EoAuN6ThstSUUIyVSECSL
abVohCM1mtd81Y02UlTCvr2qfDYdLNh6IJpL1XBWJ38+W+5XlVOLJw94UdntLC4Q
hwBk6ho+bQvAtJOsqo6CXSb0oIkwsUGiI+HAPQJ19XeBTW/aFq5rCcozBgbxo5sx
a8XUiqc7rjOisMlVrzzKXxWqi6JLhvLiVAbwQgO+V1+fVyeACj1lGPbcP1LdL2VJ
w6BYa8S4Wz08RacThyjRVjJXa4BNSCl0Vg6Jr5bI4G0xw2BJq/mSvk3GanM01NXM
mFRL2H6lqILFcYHKkJwQsPa5pLDH4omyzmEe+3aXVLLA//tAtEj7kNKaKDxuFEi4
437kKYCOxWQIwvxsHY2grKOZ6sDpTLziNTj+athucWs1bo7lAJOTlFmZXCxCsiV6
rwJ1U029UWUwNe5REXxb0avr/2dtNi6uu0QxHrPszBsM6XYIKaPZDU9GcSMh+thp
i8uzefZg1zIiGjzvI6y0m0WK6w4oztqFfCyFst435caGygDzI1KJFKm3HPI802J/
rriebpBdKb6xifHBH3qtY5W+FGY57Mc9FuYMR73W9XCVCh+LASCiJbFj2Qfthl8a
m7EvXpBdWYIsjl/Z7wxcyr1n0bJEdRhvPjY7bL9cHO525/ul38EB0rJbMZNtYxM+
zMGZiXDC452s+Mgn7lx195SsJnI1Eup8LAuxqbdsGA564hZyKw2c9FwRmJnH1SvY
pcOb+FAuVst1MkA09rXpacMBVjqCmuYDQ3JmZKb2Gh2qrjOWDRe4Qi6bpfrOrH9K
kv8/NZBJGfBRKNxXcFNxhcMS9pfJdym6KHfBAiZecDh6c3EjCoDjbdKHnWsZlnd5
5HU1A/59o0T6o4xxWgFNx7PXYnUiiFmC1vOb4RRK8SHnpu5LcReK2UESg0gzLXtz
A7YvrU/g3Fp0Xzzi7r+IORBSy3Wyh9/7njaMwybYcLl6JafwVMhM7S7OnRUu1/HW
qHaLeyurYBtu1Qriv4fO0iJFllwOUV+RnC5BGM/vaJ4bQxurz2mcj/r+EpVXDLG8
oE0MG1ddxCg050vUAIQZEuR4qG1NwhwmvlX7KVUpSs+4fjn1Urx4j7hEYlZZQmNN
YGEKO3GTQU//yRh2r23ljLwTI1qgmUQxnGaRruPsdyIkpu24xU355To2/Uyh6Faf
/xA4GmCQSD/bhba28rXVxF0i5yP0QftSOBVskv48OfevQ8LCHWJUCrgncC7kvvFB
0b5hbrcWXPWgdW5yGBFjdUJPZclMcosZ0NX2Hb1tQsjDj5Juwzf3fviyUnZvc2cH
X0IrT+6duYCQ8+TZBvcnJKWI6JhnkwvyUcaUPJHR55Ph1vb5T/l7QePlKXXeuQus
f/0Breptcnzchvvc2qe/mm7Q4iyYfrCZTvUhnRr0dwva1IrEEqBaKYZdhAdoDGWi
0yLN6bPgql3mNTIUX9p5Y0XVWEQuAuIYPAzWWDRe+Uk8CelmJtvF9BLxx1uwBA/4
ViBlNFc2ttXF5K+pc+bTvWk5BOjZ2GBq10PpkVh3103nXi1kqakJucbch7xhHzug
egz+Cpw1/s1vkP+SSYh9xDzrSMQT86pYuw+MgHt9yFk8f4LSGBfLNtmljnUznt2d
wkVYmvMvlEgA7DTllHxbjaDoPDjg9Eej3PJYPpZ2Q6ShqRS2IpynqcLoAaspSgpY
UAp5v5LraE6r3VgSrl8oCrXByl/hKNe7g3tK/PuLeH0B78/jXJ7v4PkvpW+ZZ2zR
zZLPTr47h8r44QqWRQIEavyA7EyNfOp8BkK7MbPyd9vIDSQYtEREQ9eDql47N0An
H3eRBK2q9KtN2F9izGn584Ux5ZNh+RHz63VlHLxnnBV3f5cwoYTvdk7L7S7F5LNh
70V5gBxHXeOFa9v30aPSOkKJOOouE8WL/SsZBsZtTTGsfLHr5IdAvwMiSJGY2p5u
FAhJS5Q+GXjyhU9H7qa4Rg1wPK3+Fz2WsPsjKnhKsYfQd0+d54bcZbpenB4OirkQ
xjbpaz5iS6Jf2uzlisMdQ0XE76yYpi5WDrCXMBaJQumpC8DXlWfPAh+CipF5qa1H
ZzmC3SqTreUDdMvr5rsPMZAN0KIkB6/Z5wobUpVt7TeLMuXeeWFznTTp6BoyfQXz
2N7QYyusOLxfz6hKCzl4cUgZtRDkbCFkWGjY4EBrBY+ocPb+W8DGLS8IbmaiEM4I
H4r/boRO9/oUj/BZzXQss2Y4lSKmNn2PUEAuvMZAEK+t7b+W86tkUfjBBKtFlUlG
k/Z7a8n19L9B5ynQWaZVHMTHXQmZ1mSOrejmvQttmAV5JQ1rcWffIbEaATqzFG2y
WO51S4VCcfka+MtS00+c7SNxX+qNNy60cJNfAGwaUOV03qrD6y15todJQzNZXXHf
abnCCbRIbtNSSQuXs3s6Uwll54UyfV/zKoxVdNUprNuXveeG3wraJTWuv9GkC7L/
AEZWaKNGRXRfVWBEApCWnsspSz8Uc/P8fQCULgJVOW91u9MfsqvbDUI48PWAxqlv
7gXpE1U249/jXUgVxgUrAJaKzd8OJ69zAVOOuqBpuHlwamvLSwSp1IjekC67wyFh
RRKDBrp8qYRlV6PE5KNwU0Krb78ytyIFJekT2qh25AH9RyLmG5rdyL8fL8MfYdE8
CPbgLS9HMe3UFI0Wbnjc3cV0HHx3cCg6wTJoRq5J19HTHFD7sekjH6Va2fQ0cn+s
K/SvuK+yAhmoaUP5B+F+osqtW0IIinraDSdoW3uGAlTuosDEVdCURHjZwH+qTYuY
CF3qGU9ERnsmEmTWIRnATZj6E/xU/irvA2VnDNGfgoAgtawCFsYHFfQHYaM7VnQm
fyU+XbZdJB463y2fmHa64EOwbbQgTU7dURHPL+xHMlB+7RAOokwEg6B/K74IMR3f
JVbiWWdnXxgEyoepw5Uu6pO/js5zGBuMjqFfwcqv43fkwwuGyKhWrPh6ThLIcdo9
g9jYnbQPND3gcc0EaF6U0MVor/TjR20ZtUAwDCkLyWomClahXMUp51ekGvaXdIV7
chQlNCJi7FiNhALq7du2Cws1j0hQnXc83zY8DksYAiRoWdU+ZiBSJhxisyagwb/i
XPth4OCqFBMTwXrnpdpeSzRn/IRwpcocZRrfHcjWKBnNirAcefc1n0pBza5xI4l6
pCMVH+HJAAVOzXccQHhexA1yqSHu/v09vG3z5o1j9FceeT10QCMJRL9nwhF7Ixny
NVA7Adp1FwJlT34fFAlr7zEfUkJrS7IXZhIijYtloyE4sdyTzW67iCDCZTvMTsUI
c1sc5itvwOgMVUuVG2++I2E2f7yejspT3qgiuHcZh/rWRH9MnpeXeM8kDx1P6q7N
jbuLiOEBKh6OoAq3yYokmluQWQCj54o6YVS7JwO0tswhok3JYYZKe12lz0CuR/nZ
LmCoM1tA6ifFKx/dt2aEla0OOMpspVS6aTprOAgRoOjuuyX+cTWqM4Az//PvQxlA
+IAFsj/aNX7lWU24YLv3lPDKAVIy+4Z3F0Mae9ShshwAGzmjwoCfTzHWmS+Zxk1V
30SbhxxNGYgLlYjQbpgjAqt2cpinyG4NruGsS2xpJw71QiMhb2CSSPUPKrQPObLG
Qi53HQBoipXLy6ZkBWuuRjU+dzNejUqE/5fXvZyIqgRibhamkHRkwoMZ6YhMwKk4
U2yBfeOffNomX6CvoWJxuC6F7G8hO8DiHTF4akhVgFF2faLdsPgrmc7NqJ8qODwS
yiqUo21S8svs8l2efVsrJ96kAItebnULlAePs4knxDN7DGxZTva9aL1ZyY54jfJb
yOpsbmlCGGV7ruosPaf12EcGe9jjYXezcyO55n/eTz5SBv/G7ZG3qUnHIdsO6Ze0
sILotQXHdeJfTBIvsfYNp2UKLfY/GU8jAlvSVOcyYkHDVWsYm3Wsa5kkRT2CaRTU
alwMR8I0vfuxch2zzyaRdFsAfklPx7VXxyUNdwUhuXVS2scDd9P8M2e+RnbznXf/
lheWMACPNmE0im1hf4BlNPmZa3xxodyI3ZODtrq+aVK4Uzg7XfBGjypnnEJf6X2Z
YpWTcDgEweKM+wx3llNm42LneNm7WeCIgM7D+1anKFOC0UilsvqEOyQYa4xVVXkk
roPaaoLYffARYd7K6sRpz+gj2JYckUONeCrYWKcflDGLiRetOKD7Tl0IUQzwxik/
euTdMcXYq1lXeBHrbAve4gxEwQaDFqHPlngn53rQ1TApgxttFeyJQfLbLPMG8Jl7
iZKxGvKDJ1FUnFLCslepFm31i6dlXOEyJ+lY/uPZThMGaY7BHBmklz3rahqWloRX
4CiapgPNDjPGsNbow1ssRpyZDeb5m8nXCB02ZPXo64o1+9Z4o2/GA79kdN5yHlDn
59Z0kqM0UQNBvN7RIjxyL1L42VO4HODVsS+YvMY2gX0JDfjEvJgmY/UkAVuAiMvf
Ye5Clu1piw1+S2DpQ5w/Vqv7xoqJf+MQtMUwLNquOBBsZORNG9uMezmi2F1TxeJ1
UTp+16Y1kN79rjfv1Wi1Eo04heYDXlWcGP4P2JiIh5xUeJALPymb7JxeSYyUr6GH
3XeLwX4NrS5XXsLcLSAQLVBiu0gS1w8vWD+DabreLui/e5qnuF5pNFrZnzNvGGzM
CVRBX6sClCvTEDZaYbxoYT9wMjfKjWsXPdhH6xfTV5C3Dn56e0IIYZyTYRPhFI9H
CworulNNbiCyOiD07VuL0ZmYuqXqtLAWsApxPIgk/AYZKSARutBgP/q4eHkvK5fX
uDJfP/9SNV0JKOGL3nmgN10b4FzhV3N/FszLwpizH+DrASB1tltk6tz98WNBxvPn
0t2T0yCScP4xLte0o03HLypoH6i6s50in82FLhqyaZ98j2wq8OTpd2UVmvSMNDnA
UKrEhgPrvpCt9vkLg+P5dNo3qtG/hmiC4Ozkdigy8LuMpeGa1K6fyXyMmGUJlnrB
uzRFzq3dMavxeDR1BCIlVEyYX0NUSRRXLQpcnU0roV1Ti4z/SJzDLEtS5ITnZ4k0
rRk8LF27p9BwLkcazf8+NrbWKEtjKY47yRX33WNAtxcQ7EqLyWL8Tly0R/eYWgIM
AmRI+vvttogGGk3SgL/etNDlSK9wRlCSlNPoiweSe2AhlDqarv+lBBloq5p9qNb2
pssvzmdwRbZSnswSlvAWEZcZS4JC2hKCb6ZIi/n+Y77WRwCuUE1SVnQrPhnXAxS1
tZw/r8FcEnbW0RtVuv0ipOT+rMaLvPqoqUEt3viTu3RqrdC512n3xBNuPqMqTXu4
HnWEK8Cm42gvHw4YNjA/4uHhf1qGWP4Mzo0U4hHaDkLINgWD1Tp8O7y4+f0nB3TI
GceC29gaR8tamgwrvnBHr6+GPSH6s4SLxwVxcA12hAZwltXMZmZEwaDchG64j/wI
VglBRabeqJzp9SVYcxeVpEar0DIFZy7BP887UX3hh3wtPjSm5zfieldflUe2Xpnu
ceySnH94+W9VZY5/JxjLGgJ4rTtkLE0SItw3UfZWz1BI+1QHGSEnYzB//3+vio5J
0acW/u7YvG8iL7dQM0H8nXrbYvHHZbF5lsXyL4i54cW762O00/u90j3qMEHaalFc
917pw34D/VbMa0b5JeUDeEsqRk0FdUU0aZvX7NglVebP2YUHfPDppdkb4G3XBlLe
JMc9+0XFXHeS/lkf3iCd20RYgk3pvbUvQoVB3OpInr6wG5bf5yslUBf8LPmchvHI
txI6JAUHGtxrQ25g+3PNrwwguT9KzzIbw2fUQnzNESqV6QdQxeqPyub/GPAqJ3DH
1qzwbRxsFlzlIac8J4yQWIAuF9rW2z7zrKbUBcbE7ZhOsJnB7+JRMdoHLjz551tt
F41LV9LcuGz2nn1jjpJzV7a7eTBjlTvc/kMhU/odXOy5/Pr/D2RiDb8Z8+MXtBLm
RVgiV6CV1G40f9L+a1pR/x1/RxWUduDEcaZ4y9Bs8s0DmR5w8qsHp13993unwVnW
l+kuRMjMPwE0ENBBq+VdFEiACG4tJoucNal8OxivXpp9EB6PeM8QSJ2dJJLEJM6h
qx8Fuh4Ae+28Qm1Lt1jPQuGCMo1p1GRBSpYP1th5brkhRHJOc7Pmkb+hzygx/ryO
+aSulugKkPgpQTO4vKjohPGIn6mhP9PlJGPC7Mh56IibxFvlLFZvinKR5+d9Ab0Y
anh8VFLTJyAJD4WN/jBlj2kxMBSPi7xyxogMxMiD50K9shIjoiyt2U75WCT94cy6
pGoChYyrjDTxUzvP5NXXHO4RxKB27xdTPoJpurTREu1sc+bICEdLC3QKjOw8Gl8H
csPB72qfkhd19V4SMJGhLgX70i2uKhRv+0B9UkTp8oOFIJ9EUP/IWmzEbePwtfcA
utIwxBjNjCcqOK1jfxVJA3efn5OQwILkhfsJCz6YaYRnW2xj4eM5zuSZvozLVqFw
AccUXZ32oM62T4bvQznwuKuSPTRaZskXSaUtJ9JWwFrqSfIWbc9UkVR+hR72RUhv
3CvpgqTMgaVUWe5kXPEeCUjzz2haPkyn4UuX1NtyCqbQxofLUpG882ks64Oe3nP6
HGxlTLzDrifU3NUO7ykbbQKxwf0M+l2RwyP434VoXcmtOFxdKBkt1D/THRrXDB8X
XzlwSaqPdSpsH+Eirm5uUX8eQZINAM/AKsesfvPvycY5jWiUL+A4j1tFMmUlOrDf
LhD6eoONI1r6ysLWzmEQpGoQPI2wyE9NjsPXTd+h6Ohx6sC9MMgmMYtZO9HL99yN
SpaGYbIliJMPwu3u0ekXT7uoOcttNyEWjpHEpgpfq3qaPMgpuEQ8Np8c32hcFCrN
8g4SWs7bfnjCI3cnLTzInDH2G23+UPt6GZrhm9ZBZenLZJQ0+5KOKQz4XYqkKW2V
NGoNy4SXR5brC9sXR3gO9rFe2KPp1JDS1mcBqyfChyLG7012YOq62wzY1CxU6KEE
eAWiFfigiDHusFtFHGG6yGLmkNNE1Vo6ZYFRwuS3YtQP2JwSfgM19RWYq3qR56Xj
Nci/Pwfuuw5tPsU+qrmgefZkslvvnqSP8rJlcuAasJge5ItV/scnwNC6pAqf+AWL
TZKeA5Yb68+Lp+rch8UVYh+SJSigDiVpQBIxV7cKEu+n/7JflejiWi0+UBaBUG01
8kA/YpEpcJ0TMw+2tq83Jx0ePciS6MTDNFWBZgyBSTPvCIFnyTYAzWQQ1NLO7oL4
6uaWjGPIldjWkl9/lz85TlJa3mo8XKH+o79qRjx0y0/kJgLozD7YtG4c5mLBKHTd
W1r/dXSeHEmY9HvcfdTQUdjV2Jaln7brwEzouTHq59jGN+ipAIe4R6b3MWiG/6kA
mnwfJ/bc9hkpP6j1Acw7zFIEQD7YJU1dgjAUfzKQ/aYSlD9uTooR8gn6oUGV2CZR
V0VWgwtGod3qX+dnh2OSYe66KHc753GbtR01fHpuPy3QgjY/Ue4P3z8w0nBinP0n
BO40UisxACI5apOaMDAvRt51BawB5vMe3k7C30rKMYradnyQSbqelauYwQ+TmZnZ
othXLto5UKFynVWSDy5ENMAohgg+enMTxTKApG+Tly4vJw8LSw2BYK/jFCtl6czy
pjlBPeenfq3JLLk70rU5S0c1TnW67W/QosqgadBnRBEGH4Ect8avhd6MiTImlFaV
01NhmrUcroowrAulsj73gaT5yeHxwDvMSv8rFGk2BKxb+aC5Gb8g8+/0mhs9RMkx
iVIR0t4bi2cpIg/j1uuZFL/0Ei44RrJV4U4oF/BZ+ZWVWlJLhIFZghj+tnY6IWtp
KpOlDO0Q7r2Xl8uFJsORZS07jx3zV3xxmqsoBllKaXFaMC8enMXg8KZnv7JkdeIt
KA+4DDf5rJ160KiXCpWkQjUbjI/M9JmnjttJUQxqnCznJWYKuiCMMNaQIZOpJXS8
2BuYGvoVsTBEzoHGLnxs7ZvNzxuKvrotbZdpjz76hZXu0yJeVWnH+uug4gx0e4pN
hvK1gxECk4MYomoGeP+rKpmPF4r3Z65tkUNsG1Cd8PA8W4tI5dRiJQS4T9QLQJbV
0ovSC8uJeXp89Uw+i/rplvE71CN/r8Mq/WHRGTsY1fwuZLklXjzpqcCNXiN0c42V
+fCR/vP3vwDwxlYQqf62SKqsDTyYgnhcEovqz1hjJyxOp+kkv412JLXJvuEsG5/S
b0RoB1ppAR5iin5EVCqDgYkP1Uv/3y7xhy8eGmFQUPqK5+X1E8ZgAuDWS2JYIsp4
jJOfDw9BXcL/bxEWwODGU9YsxBV45UvVgixBTF+bABK9IAR/SRJ2PywtE4FUJYwi
xY2tWu/mq4Mur8btYKJUCrE+fkR8ny0mawkzm22FHBS5j5G5VQwqOvloinDcT9x5
C3m43Mk6FgRa4CzzA9jbi5toRFPBjpzglLkEU8EkFGet4U9gNJeQsIj59GBbAGXC
fRHchjY0uLnyPpR2xhsgZ8eOst9qiqhZaMuxmIjtVjKxkJKSY1MjGnImsZ8WdZ9e
8XX9V5fWnTkuF5cDjVOpiFQZvzClPVKEPIlvjkneJVOUm2gf4EfY1/NappILgfdA
8eVt1dvCjmp8taitAI7HWdoLGk0oqDOCzvQfL/63/yDXIToCHx4fJSzJZlWBwK28
QMrGvdKG8DChfgYcJMgwVJYg9B2KnzcucysGMepJ7ZIX6R1BPQwydaG+dk3M5Ft/
rcqVX2P2lOiwVSDjb8VzLwCM/6RnUwhvJeEXKjEPzQU/IECtoGhYdYy+wJ3Pq/M2
vdknfCShWEW+IT4SQiWQn2RP/OrJcEfe97zrBiVdA52Fnj4+yLy9PPV62mXR6+s7
unbVU5qTm7btJevKRVNLjoTUXTPLvBlo1MQCmfsTnNxoRg8FqYapTiiwS2QI0Tp7
HCkwzLwLR2/bYYn2hfgHSTpXwe42p2LQ4MUlJQigPp/dh8c+Ibz8Dcxb0ck3dnR1
U21RW4PKt1AekjWa5ZNfVdplodjeGRvlnjG6ohA+oATZJdPqMq4sHAGMBQ5mKhJk
1NRuX9RERsutdl3QRHOFmVUvufg6024PQPRySS4dFDcSOXANYe/KIgzUd6YBZgSN
UYqnJyBqkGJXb/uUSplqNTBxhuroAJPf4PCAN8xPmTnyDaH23LA6T7EhBcPXd4qy
Gk72+d70W87/GMMnD12H+aHR9o255+4n9kTR+2ok1ZxRup/EvMkTDqIEG2EhjqBe
bV0i4eCYSuRPagXCPZMVrcxGpX9q2GZmzsrhuTeI4Mzdsansir/WLa6PIrWGk0ty
uMs2bd3cmBv8yfsVhndrcPGXp3vVW/ArQdLup9pcLs20DWBbAFVAKbinoee3igUN
T6dk3ScfuAIdZtTL7nlhz8IyqPmH2JQc7SrMQLLDbNSpB/S6RErYk8XVjkDv2gbO
u4TAbSkyw5zJPEz1BVArYTPYGfvZwgmOjXb34ErfxvlHiDU50bfKoh8HKiHYkcon
4N2wkzveXSIDrTLi+bjiLJPzufPd0dn01jyLilrLmi7kAO9ZatYTuben2iH+JnTV
sBOBYrHiuhujRbXrDCNu3BTMdtSQZco1CsNuu/99nH4GJtd2S1VS+xi8Vfs9n/wW
cAs5XTE5CV6Wr6CX49Av8ThSGa4/Rm4Ju71qGVAVLDKuhmVqzP7q/K1wHoORNabf
oO+kYf1G62vleQIRHj9PWM8yiH3WUerIldqeE+MjlEM/n0evOgDKCQEt9YWgcy2M
+bt6PPb4SoOLqpoo0UPtlSxNjZMGf5esU191kw5VFaM9YfIb/MxELFhawjSnMF6R
uUaU5zIEZaPml8wXLUivrFs3G1x+7xNVV9MTUVTqJ/gCszqShMyRb/VtSS4bDayZ
TgYnO8iJmUre+uk0Az2SybjKOKENa+6IhXDKBIMbrDTN5Ym9wKd6q74498JQTfxP
1k+OEJW8pYt0gC728afuoUqDenupxGs7OiLmJqKmL0NHuekHW6VwnkKKgcSTu6KT
JvlobSMcNQeb5xbFxE/j3dxYqU2At28Zd58kQHdrOiX9kEPag9yeJigmuZm5hEr0
/9j9EypfkoGxmD/kCQmdbBqRcyx06gQQdcE2kOgUVWVAuECo8xMcjSvdXWD39YjU
5+byPKGfys+NoFCJvAPdChKeiI9iw1019+aTNeLlL5PRkp+Q/TqBtZ94fckmI8qc
Y+dkDW/jV4ZnYocmHS1WaQU6lCTz3NeTDNMTX/wxy29WNP4Ym++O8ri2lX2lGfOz
xFoshLLfRbZ5i5PVqxfsexK4zz1bq6DVCr4xNzNu5W/Tsn5K14ixRQld2Q/PxeIf
/sMtwnhttX+qOCCuCWmZhTIsO5NEk5UBLLMjp8xQKm6ZtUBwehN27j2czAGNnhGE
H1sFtrEE8Es618zIF9cqM8UgyfYsvLKdGSuXZwd5dXjkEGQYBbak9tTyA0K+5eah
IlRjx944UmsCEYh1RaqiXYCT3NUNb9p0KCwCU3r3Bx94WTTX1Icl4Ev1TO1iajXE
EB0xOm8kManIHD0Jn4t4KlyF5vBWolTjihc3SXGJ5iQSlSSNQK2SpPEkKgzeCBnM
MilrqxgGeUpfxxRxb2YWBSNCGDS2U31F5o1r3oraGK8LNZUReppOH1kLePoeiHYJ
HQAdJ70sIx7xtBycbNRWIhtc71qWKke85rsxxmyh5sS8qvf41JCcktgCzVobDRcu
O29/SO6azgYVwz+NPUo/I3yB4EmfZiGW+VuxkC4mhS7gFZxM7iyRLwLDP1+wIGN5
fXIhD7dnyJEW1WL3npmG1xQjOGqqWwHz4e80wkIMrFih0n5ja4H/51vhB7RAsCjR
dNxDTF/m/IapuuZrusiICHRTKHMfx7r9BGRFpDzjXDhXYGTt601grp2ozftlwR2F
Zl7prgLVV2M1W3g57+j18neZg8tGCEQ3y72QmE9B2WRPIxWGeEC6PanDi+Ep95v9
lqtlKfutBQMga6DLKUe6zhIsJ4WcH9fZf2ANRLzXQrVQCOPdOvFbNdabrxiU1aGZ
xC/bsfvAcvwQXonm9JmUSazlNWBRkClLzSCeB0yGk0mPk/FG+TkYuDD0q22C/vn7
X5M6WozUvbmoSmNmXWWBFquQcEf9y2sK9me+tu6G/D/78RvxhHYJEcTcZlbk01D+
9OyD//YcvcicfkYRzOQG3CPd7MVmItNGLso9jC9oeX+kcrevOWL7B+SCL7KQX44Y
NGJz2rTreibMxo/oVCZvtKXIq+Pz6Zvmyo8gI3E7OMh5SZSVjjmcDcGrS476Nrk1
oaapvU/r1M8LcJWxejNu0wMoJtqP78hBc4DvOGqfNW47iPnfQQvpL5FGkAx+owVW
plfkbJPXPXSIR84VTdV7MVkKjB+1YBxJ/P+zS3nnEZEcOjVTgN51Tp9Kf7ZB9kYg
Ui23tGuBApHHnFtqqYZxbjuIng17ImgfFUDGrg/rUNyH4hKZbY4QKduRNpS1GZnh
jVHnHRjNysJKNZUda1RkPU4NcE8v8L9/kf2PmAi2C5+gj0lmbY8WTzCULdRZfg7b
B/Sy5fJg895twLhO9+J3DrCinogtHy2zbhmJx4KMrmrcp4AqMkh0/QZY1SWauSfx
ZnVRkzuCS2xSWZtQ3QIQQ1DRukGms1vByAPUt/ZQ91dA6KbLRQKiR7MP3yUwklHW
ZIu5j9Vo0vdnVlGHkAa/PG8am580ffSCkAk9EvfMY6GYcB42n9Xr5WcEBwX3DmZp
dLmR7lKopqsk6C8dzqHNAEGjDMSZbpP2PQJT8e2Zjs81sh4Q5zy5v4xPLC8TkS4I
uN4oKVJsuua8HDj3vJ2bmaLoetDlqeJWETKaLp/Tox05I+2SBsQ8rv1i1i936rtv
bTH8azMV02JEkIuZo6KhAdU0ant9z1qlG0pYsPwFRiWqSGJKRGIZr9THnu7TYp9P
XGQnDBSr7NMjsHHV2Ys3QUMnLIUQnfjJdvJh2XbhxbMM6c3q54gohj8i6c2LHKkS
iCfLOI4kb5sT/RjIud2Nl8zVVZxgzMme19sm0SMpI3ykqZvwBossEDvA5U6q4SRc
M6xNqJXkh8n7VbfnGT8vScXXGAq1kg0NI1A6ayVnwKRsDm+WuZUJO0+4+IiFeIEq
WPJipGNO8nSfRHwbA3xLgq2nsOm0hpQMfPVUh/bEI1E9lBGohwAwySD2o/YGgQn2
E2Ccs29CGzZL9nID2T4uNj4KoxaHlXkt8tj2lJyKDxtRLE/gqorcHMUrnUH7yVRZ
68cqqcw989X03BCl0eeYcPbjPdjmwBLK5U+w3yom9PKy7X+nryIGzPPcXYKHR1CV
Z0VnmZqMA6O65N8euOu8g8PrqttYN942xyAuBeHK15Ed/ylrINZXw0NtJWDEBBur
jRyAB1t5MRtoajgNXu0xFI1Hi/a33FEIz1f0HQqMZOXEjtAVs1AndbspthuDfeMz
AG8gA6b4gone2MRaUNDTl8aVxh2tbFXeeLU6FGPCqoRzI7wZvsvR9ugOkwtJjfxg
8wmVrZzRc2Gr0udEdJRPQwV6soEPQukDE8tJFjVFcDpyGv7PUQicQHJCcFnLUEq7
kc0vO4FW4VXg1flAZS+ed+lHUGbm4vIMGDUu1k3/j3hPB2dlZszcP7XDuniRBK2a
R0J2D3Q6QvqJFNS0BMUWiadF5Zuc01is75PdeIBYtsqS+1SWk7Apu60RGd7v8BKL
cE9US4tY17aHdkvmCAK53Cp4Nyq+nkVrqQO4UvIO3wZg3Zz/l1Q20wMDkmSYeN0I
9zWiz0fhSgj94e2aBKdbvYteqNeGpYDHWcVCASujN49c6nou6e9yHib/21jS6mbU
sHHjRvL1HaN63CJH5vTc8Xk/pasXATdFE3Sd0YuwPhFtlEhTqVWmazPyD6wlMspC
KI9bCJmt7frGgDTCFcBj6+HzvJeWnHCSOeWm50jIg8e0XMVrfVfLKyrF9ESE2KPs
8BT+LOsvEXQTkNufBsGGseXT8erQarqwOJ6bDiw2g+om7oaHQN134hg7kMz8nJv7
a0lgim6TF58+qY03rOYg0scpwLaxH0uMJ+H0hlBWAmCRhv+8eBKmdb6soPp9p9g/
F5UKtxamWcW9vVoWKKB6Vq3RpyWZtL581BuCT5xne8kZOLmxilcOagpay0g2ykVA
noxzTqb3U3QrW39VqQOcOOuMH5G1b+aKXgCCQYHD+2+izXxZRW079IIBZhp3IkQw
R4464d4lZiQqOZ634IFuPvJLDHzzk8K+ARAaluqB+QY9HBmZJxrD/+NSPKVEdz4W
slHhL1CYUVzrZBw9qPvzo41DXr43wbCffX90WBegyTgpn57IFvxPcg37xRUC20st
uiT8s7lt5AHBgN9Xbqo9lLwryDNxAJg6XqKv3KtQDfQrniIroj96r0oc51sDm0Fj
Ut6hTU10HOX+sV9T21AWi6Smg16bwoS8SSqeJ0QtnGp9vDo6LwqdlYIrE8xMyL8t
GF3+ddNaH6BEZxACiK3XsQqn077/U6w7MjpA6TlbaeGpbOVzWLqK0DEBZQF+Z5v8
ljPygI3Fk78c4Tai4AvoKG/ko9wlDw70Td43SqFclKwUzOCsUB0ByVYSvvxmlGL5
XWglNtYJLy9ku+ept60FjrgBR7XS/3G5NhEujIc+RWbYRL2alc+cS0eMtjp3NqZ8
JeYr6Xztj4Oduod8o1UVHk2Th/nRJ3VA7VxWd2xpDFtPhelcdWFDgGbcGwdQ1H5i
eXanmNwyGc/riCYFsKfpXut7GQmNkpqWOsOteYzy7jw1h4kSZ5aPbiZm6s2S7nQt
BqEdtWFAMrBCF2QklgznIyPy9AWGEhztd17lFfg+jWNcWyS3X0UOLxsC+6iPdqS5
WoIOd1RFt4bRjneM9FkAchcEIvLe9+jI4I5a15rTjnp4y7a5M1Sugi48vhUGLiQQ
KpcBOkRBZ+fc32G5XjunPxeLOVmlxXPxVBvqibmspoNuGHDguBKu0Ur8Q1z20YpN
KqySJ431Y26sC0pQYrnb09fdkBbtg0BOlUVCl96BuxG7fxpPCxxgiHxHltZVUGNO
kJNvzv9h0LXI9BRiT45wlEX1IXqhY10uMEBZ9nazKKwT9GMhr66EnAbyg/npvoa8
BCgywcFHtJ8kiLqGw6DNeV0MBCfqITF74noR4bXjuRjeFbFY3wiSG0nbHlkrQqRy
3COUYMqZ+dkdAPRDKjbdUFfYiv4Xl7vym7qSsrY4B6V7FpX9oJM9lox0NiufU/OZ
mTGlM9wgEhJyY2SP0YHkuzQq6BF0jXqo/OgyhgzQL7OSC+QjUDsbx1WAeksuUNIc
oH9t/XkDnLlYD/J7pC+UOJvGym5ICNY3oNwI/A+PRU9G9T6oXpC1xGA+nQnfTwBa
ML5GnjQXs/GNlX6XxH9fPzE/IHv6tHJVDux4J/Lou4T2iuBd0ljbD/RE6qKtHZbd
sDBoher6k+yRt4rmJZahwNb8gcdwE1teUCbhKBY7Xak8hYog2b/0utri/e0jPSMc
MOf9GZi+oIqosh8z3uoDiSd2CMb5xQ2nriykfSHruv4Rovp0RRp20ueA0EKi9YTo
k/PNLqZBqOe1YhbI2LhhGGUeS4Yt6F2ixv9vUO4JZpno5V7MVVScTNRvU5345IeV
lZOX7mNgPaKIHEcMAgvlPs0eGyTtze904jWn3Cxf1VvLcGbg3JaJruVUzxU/Ev/U
5Nm6XyDek4UsridJDDr6FyP+alSt+3ILXrJe0T05KAiysW3XHMGcjkEeN3RS42ep
txFgrpwVNCbY1IVHfU5r8OMSuur8+mZL90GubocI9xT9X2NGsAhSLNN7e7FBetLO
EDlNppK8rRk9XMYrIFCEv70+E+hbrXVXD0QXFOjChlXXdnzyb+Gu5KpbV+L8Eozy
2S+sHTpFFhT+2um1Kb806be0pvHjo6iHfu2FBp8MIXFZaHlFcT23d5ynYVHtK76f
ZvSV8pjGSqtvaMUsoALFB7vkeCF/8nHH0qgfOUk1X+Cypvz7Y1VYcvIiNhr1V73+
p5LSHvn2CRi3NRggXygKSCJ+5gfccGoH/WKyvCbinMKnkO2AJ46HJVGbHk8ygVIY
5gPIv7a67PdKZCx2hnZlEjWNLip08K811GXhzlS48CuGzHP86hXNuaeokxF1R2y9
U/H+kUVe8oCIPrUNyW6dMVppHUzQ8esJbnhP2staY6qz8NhgT0V0E0Cts8nZRNqe
eROXTbMMFDD/v/54qhPGYKeVoAa9VE+eEtrX72ppnwBA/JBlOnEO5JoWm8OaOUhp
B9NuGOZ/fjJujEv7GEXCG5FJAL8kNjj8cHa//OIRKKmiTgu9a9f1/q02lCuY+4//
ahAaCGCQaWkpwTweYKxoTPewOPLG5eJCurOH4CU4E8bCCBWXCGXECcVVMmLOPSmb
SLErQ5cNrblOalOVI55LInPnLFmMEqp5VfkOOriRCliS70YMnkShq2bNkN88limM
xU9MTR+RprkY6FTN5vYMSPyxakfOvNL8TzF11/iJ1eURYQUsSPOpurV3Jv+cEs0Y
g06s4tZyNrHCnSeaKd94I4cByKo/hi17R7PG0Oxwbo61l11HWtSB+/vPbdvpRzxr
Ma5CfdhC/WMJXefF3Z7ZImPu3GHC7AmvotPkhjVSGug7RRTsB+UCXu04w4/2mBNc
LZnAX0jNMvBYHro1o8zAU/M+0GE3ifh0f7elGVSrGckXmze66LXgw1ndW2Z0htjB
q4c0fFpll2LrmluaJDCT0tgmpUY8I0KmAXMXtsN1Mdfz4mJY+Pg+Y0s1IPbAb5Dz
E84rbepLf2Y3bqWR49RMUl0sQR2jRXo/n+ukEBsTpfnW+uGVugHE9c+wgr+ppTi/
6rhpYKc/gO+FgOH3FB17UXQ9JJ6apFb69Y8GZusTnbcQMwnQyoIBZPbEniyOzNB3
CTpVQZgjCFNchrwcwYtEB8fhlytgZZIXHbjXaD4ydyFe5V0bdVKc61G+wUXNDR9A
nXx2UuiaSXEvD0+MRGU4SjdhXk/gFwwVjzkmAw27Pnx5YjdiiPnd8StieKTm2fZ5
pNVHJXzNtVV8dPoIoDQwgCcaJFGrBSTh1+3yFd6G9Q+QzqqVX65LLmW6usBSOdPt
2Mg2M96yOAySzQiKQvpb+pAChpaAT/knTzINLqVEc+zSkvzpA1wKzBOqQPK83DF5
ciYY5YbKaJjkYidg9qeRapt7dH99oCOMpFDfA1QG/5D0fbWxEMLXVV8FaTymbcR3
yZfGQVFmDZt5zob1U9oDzQGaLIKSLxBQee14yrnZZmJXX/zuKr1QiudJOHlRN7bv
s0hTWVE9grQyrcIIoJLTT6PXigA/LdN++ebWPZRbKPFsttm+6X73fKKNraY8Rxcu
qzjtVPkZ+2PLynZTGZ0xaRYJzxjNYavNrQrKy3A6ucI6JOGgW3LfeutLDfM7r5Gi
uSQCPOpbTnuYxv1Smvq4u6R0ZnJfoYFzrQueXS6+s+Hmtu86aTj5QNIkQiIkTalN
ssqKv8UageH40EbpNme7widJdXm3AbS8cnZo/dU7uiJevVLf8dw0Djcd8F4U7J0o
mhuWNodBjvmVjnAW4V6mX1KyEeCJ/SClSAFRyF3HgXi4lZh750HFUQKlaWf3otGp
9JTyCzFctDT/2NlEBi6v3wNeQk50MC1H+SilwkQQtEVwbDVNh/b408Ohzo0xYtz7
oFHIzxey8RDj0Qop8pmvpCCm/3gRjm0PoYzoMXwWZ90rkgFollxApYZwlMjCk7yB
MIpP0VL5MmCLrBna27K4JyPH9/X9d28CpftkH/kXKKE0yjKobmsQdRhfMI7MgXpQ
R2YKNqL2zBzxzZuVIws0hJsXjXcIQrXeKLD1FRA22wSK88Q/rl8A/2rQrpH+NyCS
7dkNgp/ssCsyLipy71FGvQHeqgkquGTWJ1qAVHEwqu0MlU94iZ5lR1AJL6wLmcMN
LuEeHFUkPPkX8XIQEjzjYMB0sq1n6MBpEyphRsxOCD3QyeUDCcoD2Xev2VetLnEq
HfXRAJ3JANgYOUld2RhlI52CuEDFMf2YJUMz98PFdJ0UR3FDezeKzqjPX05lBJtK
+PoyfyqYXle5fMNklYTttl2qLXHhhPQtcPdpePZp6Zli41syzD79uk/uAKP+RoJq
WD+hFi/0kcxFmzAMxLuYM007aSIkqGAyTg7g7nb0yFv1Zm77wG/Q5EfNxJ6rKpri
PL3DvSf6BrAMbOoPEcFwboT2GRt3hSqI8owPBafy4EP8U/IyLXeLZiyJ715w24kZ
GQhJ5tsJPENqSXUrerD1GDqwAZ6cSg6noVNNLi2trUSOmn2NpXwhXGTQsZA+kvug
L35GdizuVr1WCwWJohfSzgJohpGDBCYQZO1hSOa471xpNE6R/kq75b7LPwkJxCpc
9OKqedNhXG/zn8M97A0QDCkegHqYrtk8kfNDT338ox7F5Y3CKxDSDy5D5pVjWjfK
3sbskdQN81nWXPCeBERyu5U6eLlGWVYBh/Bb4FzDjWmfIH9Z+H7bx+Rz7HgiRnzk
BkxOZjaukZ7lknmO5iLZVKJ5i3iV33a643IVhAiW4nXRGJVjGUKeDnuk97nED8Kq
aBPDYQuT9+EfjfAql8yJUE4agYjWzdklFwKRsdkK01OOftMfC+Vxyh7B3U6FeLv1
ObfLH/6CD87jVlG57oWjqoTqpXoflnQp047QI5AX8AYQvvggXQe/Yzeg273y2PxL
RkAKVt8Dw8SLfBIXcByGSeizbTjTWkViRayfMq8TnEklCuRzllHhbbuV840iZGn6
z0wWpEwpwNDcg0HNblMha6Mg9pa5mPmZ7PZhy9RQirFoR4bKWxMFyIFaosOI8jke
zXBLXi7hjIO9pGcHJUghwb7PBpWSV5XMsNPx+oC4yMw4fBuNh2i1s/OcfHK5ocBP
TZmIO9MY7p7id4VbQvIuCORr5Y9MbPc1firaIqffIT0bAPNVVeFpTfJMUd2rTTkc
ML/yQuRTMR+JWLuyj9X4oPWd1FanJx4bAp0VyFQhUYFxXFqX+z8G0q1ZmMWKUwUI
q8RjkwH0ABfYePFp89kqV6Rg9Yf0frJzghwaqrKmuzXHOHp06rlgcSk7A6gHGMwj
u9ie78VumkH4CKoS+BuOAmGo6uMS4A/wRkSbRHnZ2RNdOf/w7RplpWOCfcfgVwqe
wgweHdOLYEgRBGx04lKEr8ynLcUWoJM2n4vufHo5e6GVxlwqrqFWwLHVIAkmuLXi
ZtCLp9dStlcyXFQvZE4H9pTC8iZH5cM0EAKjPhys7nw8OfhvRVooEc8uB/tFMtou
fKQKRYRbSYvZFBF0aaWtVEsNgm7laFjzJsLL239TWhLNDKoZNyTf82gNpeN+L+Lg
dqj6C3x3XbQX87FeFrBmCmUo1HsMBC/4XEr7AZC6kX21mC1KnKfs7aJDK8JeCRED
7KCu+c1fvDPDVjYBCOS9oO1CjiNKZ1hEP2vY0wx0LSeQu/55NE4gJjCmQnyUfttu
YApZBa0Cf7yhgydCcC5iVkDZFG1GjXxHr7w3Ydaovstat3AyfZQ/mbh68Q6VTtv/
j/yOunFqDGxstCSnzY82U1k5Sk5SNZM2S/EMeYW10sKc/sba+DeDoymh+/fQ093U
4CJGPc1p9xtuftF6y500gB+a63CISI29ukq7xQMOu0CqaVJUm8oCHpGrUAm41/pA
thNZ9lOR2R712grT0tgKrFgk5H6u11WjR6zwAE2YwFaLJm9wVFU0k2EcLM6sWzfh
pqxWozEnR08aRu9aXaVxeBZrGQq0+me2npLyuuIS20twefJLQ2/6GPH5UiCQFHlp
OXNNjgQ+DRi50UKetkGf65cFfGsehLgQY+1AhoeeOWwZzGA0+5dXMgl28VC9am3w
/UsCFlRyV6B2gZMvveG+ZVh13wOxOtt7SZM1yYMoQDa4p9avWr50ljmMyWGIiTYN
sfwc8ZDXVSWBhEqgHR55yXSaG4/qTUCoDNXLQsNAdRGG8XSxd/nCOILdQsMzhAXm
Vy8Rtie4llFnfcv5p9Q3Nwb//S7reQOr4WKFdp5dc/LvyUByZ0y/U1htwNaoiqGt
lWoag1juO42yO+XdZ9SbX7Jx6gQU+JK5fDICC8NPMY+/zh5gQmIMgXU93fXg8lL7
xFq+ie6KD50IuacQLM+8p/kFqc5B7NA4rxZy1icOp3OoORdoP5bDck3K4uKgxrA5
bl/OcG98Qe/tv+N0yuh4yPZrv4YjA885v0G2c8Ci63mRjDu2QVJcKv5faE+1Q11w
d/5fJ342G9HW5SkIk7wsKo5Ycq5wIEErdylMntzhfs25uNfYljc9SKcMvfoR4e2s
C6yzBpz/OHMawUKPAyQC6R3yR3Ymtr+fCa9Sz2/pkfExUzIEzhm7oqBsX1jy/mBG
45wvUgPrYBFFlqG7aP8FHxtLYPQ7v/n6qnJdX0zzZ9jsza/ZyQbgjnsis4YYulgT
S/5NdRCWRiAXzXHHyYUmq+fAD5mSIevV/Xc7k3XT1cYgeEHsriaKsscfp9OvpJfI
qVyh10ptHQeQEsHqTRfB3MWGS+d7uivsxAp8bXA+9DQyvcVX1cVglTomWeO8Yy3A
Zky2A06N2sfNEwlP6xKtxfPHAViYLrYXTl3CZGuB+A4wi5T8tyM1+LD7IjmjIqRj
15CMIrRrQzyagHEuwXaSqjpnjl//YYKM/FkcGBSOV1PqU7is+8N0IxrzU4hk/z6v
WUvsncZPZpgkHclJj1PbSGEUkk6iXNoKoC6CJ7kBlwQT1f7sYekuZ3yiYLDpY1fZ
gloYALzoKGj5vkNPNL2I6rFYmV1epSk953Z2QIyHlBePqWvZ5o8ZeV390AcK3dQH
AXTtMtNknJtGbMXMGLLYK1blRKogtFTbS71tYb0gey2EeAQ1+4Jxw+kYRkcABVzu
xsTk2Ug3pZ1ku8ZML7y7pM9Z6PgjUDlbC+zn94z8eHllcH9tuQIXNExCaHxjMlHY
KxIeG//wnSaRgc0DIn002Mw93ekki2Ygfl1uI06arGpXQs64U0F4HHFAsEUAZKXF
Wgl+MHTdhewA2DqKct0Vkvb2VMMASpBQF4YDcAGL+mtO/ZmnbI54xeDv/+CYefvN
Y6PSYp95QKsxw7BW/5eOm6d3MqTQZPnB6x5CvkWxbNrreN9mFMju+iEoTf293Guy
CgdNlE10Ltc84m0lIcj1vhxejC9aBXkHQnxloMjUckGem4/rCbbbDQWYUnf04FOf
0Vcd9BH3dS1y0GpMMLgS7TdGLesoI0QjKz2j5q0D+1RjeGyJCa0+bpSv2sFwUtSs
elGU9NPed/Y2Na3rybgjf61VgK01ZPMSNQhYUAGXbKIeQO/8zAqeTSf/jDQg6wHg
2DePNc6B0fhSTXYaJVYagO1mNOQRjz9thD4SwyER/99a23gLkxJA5DXF/wCxQYrH
P5wdL064ApCan0X0pogPCJxfqbDwndiEOoS1FVjzJ0qTDEpQbv7te53HvTxN2cE3
pkN19mS0+QEb9o897/DlsXZotnkuqIV24HUINgDONrZgLwMfNFnLGA39x5Ks6hzH
SDHDc2z0J5vaDEk/4GmMyphhi/oRxy1ArV+1vssaI1fjxWjEcZE/uqNOpFUq2vTE
Fm6yHCCXlLXE1OnKAmkJ2QHkr88TmVShOtBJVxYOGeTl/+4Hp4y8B5YfnDUtMyfC
ZlabHA+FNwo7gWZ6tPR3clqd+7hVKMh3B9MFE4AAExVzUFAVLoVTbOFqboTuYSFf
n4s+jFmUt09VQwsS58DoMaypsP2cnPYP9XGFBDk3+D/36ZI/ZND+dCcN6qATHmW3
Ew/1og+1LaFI05rbQB8pC8rVD+TdbLkHMHvhi46gFUgSwqpX5WevRPrJAcynxUcJ
NZBJhmw866Qm1ghS2h3Tx2FqpN1gT0dZvSwo0z4nKO/Nh1h36/FfqsMj+7iXjyJk
PMLNr9xZpEbzqj3qE6kJCyMZNrJ4V4oFqtpxF56/fVMTPwvDDf2Hd9dUTDAvAjzS
uttZ5Jl5+hhvcTDZ4EHfy4jFjiJnAa78irq688KAZBs4QEoqdMeJWp07XuJGgLIR
bWMkTT7vLH2VUAt38P6mCVnqdmqfNvrCSa/kxsjBpv/7F5RWjtZQxTqntOnKCfrG
XHdCTNRCdJXHhiwCvXkUzr3tLGZ0t0Svo5hy5n2uizRsUKl1D3mVl0CAiNC2Lbxk
00Uv3rumI93Y9WGq/aMWBBqJcS0QUy4d3D9gXeA2udixxWnPgWtBp2mxR0rPKB1q
aqCAz8UgUhKVJJI1yaRpxkFZtOkNBAh0kYXawWWK3Ch4yyKpAuFoTLRvzuiDLUjC
ttg1zaF5jQO9MKUs9krf47FrlYdin2tccU0+Pcjv2eEU4VaSZmFBBZHxYwADkS7p
MRPvkzaW45Kf9PN4MpsfT+wE/nbmWmgUMwxTrIdAeNllIqxV+TNlCnc8SemY4Omx
VV3w/NPjdx0gD3GxdnG/5bysJ64ncybCOV/1sQgWMEsIAfv662wFSTEvm9Cv+sNV
RZA8XOvwFqjVekI1Gp1aEfzJyIuLfecOjl2LRSGrjRRviL6BdKcbxjN6NObMvAYD
7ZWnV7IzfjM+e0oRl0Fqlyf3nbG7iM1wMEV4YOpUFb7qrGeuS+1R81alC9GK5fFK
UgB6t4/rz61UiMAhfiKhhZNZmrcU8XKxx2tWyCu1H1PlTUzqcNBiiSWwYJkDmOFZ
ie4EeW72n1S7y43Ild7QOcIWWWTvo95vELWodAQH3kVics/0W+511uq1MDLSoqzU
xw/fnrk1EKsNqgTeljbUPPCJDaVeN14TJynWersCOjIFrMswpi7cjge5qafpBdpg
NOHiz70JBPcI6V7TNC0wXnZZ10viPy16n4qeAN9Ay3xARNyp/agzp08pHI9XoK99
oLZlrbtNwYVUaBi31O4LRtx6Yhwna0XbEsDEZ2Ls2g3sbfyGgDvScL464B7FFEEv
lu1n4AoA78WxNYnd4nO4WIRDRI/agJv/TroePyRUodkNFzNkrQFv/cnIUkxADjHO
pszky7NRgKt4yCkcC0NLXSgOLNkiMT2nI5icMTMQ0UVug8avG8ODrcyZGCihtf+5
2tj/JBgWE+7taoUNTHN+fbFNGmrp71RUvADGjkxPrMODOuBObgqd09jtoJUqKfwF
FYA0BvGYd1BD9N78Y4eeYcckJiZIC0MMquYMvMbHRN4v2gsXNLEq9Vaf63QW/063
27XiHFuQcJI13CrZ5SBwwHifpywX3hHRWE3EnAgW9O4jKrzlkDbddOiaiUoWUuYf
l4P6wnvW7BrgTvPTBdPJDPR3xJ8It1EJqnz1RiES/88JFbrFHije1dvHgq/lk0VK
KebQy4oboVb2bwlJFAU71/jfiTt3zDGaIPW+9LX6tzuy6KMrdQWOE9ijtfNjkzhd
kRmaIk5NVP+9AkO9r40hE1shQuiKfZlEtFYEThqsBsWD1PT9aZ2dkzGzN9I2ZfrY
Yp3RbdEe4aAf8mnaK+vi8an0B5ecc1k7xUd4SeRFCWh1Uan3J2XnElvd321AnpNq
9paRQ8Efl6XnrfgGKZxuoPcxhOKO1AugQepn5+pCbFtH3Iw29K6/quGJnMTejE2a
l0CQv9KR4TBExiApMAgCpv3RaVmVODDS0eSfo/6Pn15hDfC33KJV2grBTzFM/00R
VFphSawMimq7hjGHmwLLASpTsi+c8uY4F8GNI4dnztBjIUKf5gp8jDtwa6dZkqFF
4O9w02g9d8DQVSJRJ1vntwI/OyODvGjSnEETcNLLMDgM0HgxODW/62TDXT3IeZEc
BQamlzworofAbjpnP/A9c5xjjkXcquzMnPtRshn9W1dmeTSOmcOmuxXe5162F+ic
Aosg0P5Yf1HZjkowOSARK549tuoW5C7qviSIBt/WoTBqtjncBg88WpXkjsrAFxLO
cR5IfPXmwnu0Fvn/56JVJLECEdK2kXpQ5G4pbtbPYiOdoO+kyTrHIKwAAnXWGktg
GMVh11KioVqS/TT4OWbUJBi6xJDcKUAAK6jiKcBPJQt0dGR39yN98VKhvNpDaDab
1dcYDDNlNygRxwI1L9M3oLX0QkBoClqqjXtzUKj2V9FKqx/14I7xbEztg0zv2uSn
VTaIZEOYiF89IdPq4sIsd87EWfARSQedjbSaweaxsnYY07SryYAokDKDTzrJQBTm
xxMhbTVXibaWWdv7ZXXUq6fuVMDlY0DYRTS4bmjGIIDCyfaVOOby6N+K436dp8xI
JYxbuxaRWqmoniU/CVHJLankUCD9KKfF6mMvNaBfFANBOg/mIm+YfrivdKZo/XbR
O0srBPDfrIRMxN6BPkUxEwnh4R+SKQwKuWz3bZVASljdQKRSJ8h2N1Mmpo4PtPKs
1cVO2EXLbP2FS5jF1ao0T0ZOdjAsAC+hsInra+4Rqz6lNBIzySYO+Z+pXpVszBqP
uDD48NaTqmMretoFRh7ONyy8vlwGruyYRsvGkcAvI6SFY6rlwRgphI0I/jCpr6Jk
DOqpo1h6HgD96E/4XoMYyOZ0ibinn95sRcQMMjul9g5Fo5xPBMUJuzdBm/0bhYfD
oRqJcoT82hRhs/U2QnBn5/9F0FL8KfaC6/P13amjzwgU3qlfe16e3agfyA65XQiL
tzV/GoQ2bFski9Xu+qNzcT6E7ZjlnimiaAn2LehnQByjgEFA2y4gfy6gUEhauBnC
qa70RmLckVqFYjM+fRuWNXcl0UwvJUu0/4X6+KuxVRrjUPT4zO9sbuhHOvzfSj/t
3b6ngJpo+Pq+505pZVTtPz/H5lYs2GloHyPAnlYWima9WiRJpXZbEJeL0AHxIS1U
8HOIpEk7LRfM8q6dwfm8nOvownYlvBJcxA2ANvJhGfaVSG7/lYAdnX96mLcX8M38
C0z2s08mtmeNIqbBe3/+HUsr7EmcbPrBcExl51r6VKCBEhYTu/J2GdIUc3/k+zH1
bF4dCHogpBovZreBnyJsBiWLJcgIQ5fN/n0pukUI7Zla58f5CUsz0PExd0eIuimr
EFZQ/mRdxRZUiaP/R7NUL5O/B7Uqznj2atZRM2cV06FNofMkdNEmK9olDp+JRrKl
3eR8wb2HiAMFXrATzPrxwEaXZa9A0EdAqk5LDbtYkMUjRWvdYFpryWRPDkMAo992
nxiPRBE+LCZueTJgoB5IlH33wEzVZZmd4wnmLSVjQfZjFJ9IJCNz0aJcwSPg3pKg
sv2jBwMqa1lJMN/v4b2dSWdg418zh3i8HOV2dI14nzoDTTcHOT5JuZ1sa4HNEa8c
mWw8S36bTngciigaVXIvNuUcIM+e2uyCbOOdEIE6oAW+kXnX1QMLT8yuIjF3ZHbS
uqaqV53bajLclHCt4vYmnkJuJYxvtfjvUzFjZQswBuEsQzp7lAo/t6BRTLEvDvHg
8Oii4aeZBtAqHT+Q2KLCvyDFVPfKBrvrE+fujlBLw7hvbPZ/T/xnGbQoRIXyhsf8
DgilelY/YpKW4vi96n2BhIG4VfdbO+u+Zz3oscoKQAu5d9bd466sABmgj7LCUTc1
mQHQBTcQqbxkHrZUAJZ6rvLukyvOhTmU8ylACgakpq1q1l+T1+/RVZjSMnLM+FTB
e8x+ZsWmMaBmcLDTSTT2q6LP256UtOQrIdN8JzXA4RcV7eJ2i9ortHn1HcNiiJPU
ZR68Q7pTyl8lr22E/G2TmxExSaIjG+P+459rZs2E+MqgDoImXhBKR/ykdln28GUe
V0aV5ectoNAfrFte6UQkj0ulBZL/Fi5DuMpXaVnBzedqvr+nXqBDaRZjuskIdkp+
PxsmM0xMInI2CnaWZ4PRZmAajmEcKML4ADqpzGFVsL1iiiFRRbgKQPMZqyyH6wMF
FPWpUcIRppWbyPapZExP0NrmuIYdEFylqRxQYjn2UW3UxSlrFVWIjOWZw/xIlfhi
I4gDhIO8lbnSJGmk03jAmRkCj9cqwINkiIx8u7EnKUMKwWhmEuJMnBzEdE6Vg6T5
2OHCxbAYK5W0lbfDhZAfHU8RBWRI7uPa0VJBVeI1vGbYa56wW1VwtH8wXKDgvubm
+ws5NIcdDYGCK4uOwcGldEVb9T9mnih1fYDNVByIElC6aCOfx0/2xL26v5CQ6oyd
eYYLdptvjGM6ezKW9xrKR5QbqLCneMNNUH7ou9/rSZZz/hsoMn5HQn+yfcHUtZSj
3v5X/xY3ejbebgp0FP+GIvYd+s8KVYC+7cvuHUqiEgTa11cYOvCQKPGFw9HSuIyg
OY+PQCYSAYj5gfz86Bl4TeKpY7RA4PVHlvW0CdqXbtbmbskHNqL8Lj7DjGv6qNpH
/WLZtsXBsj+RZ0vVab9iWs+jiQU+jHe6tN17LykAAFtjkuoEpnbwAeN4MdKC8iIu
vYSDL5HKp4zBx42Aoj2nSD6iDYBLefEfDxzMjSPdmf2V8fbdNmxzpBHxP93aAS5X
WzoREDb7MgO+IywMXkWccKwo0GsIqIo1edu85W0pIePfRJYbpVKDXqzxfQ5J6Voy
46edRnb52dEgUZRX+/7jmnCFgR/OTJRCkX2X/KX8Bs8HDhx5qWH1T7ZJC76OiJ/H
29B7OqW0B0cZHdTYQar/D3FaFT1HKUOHgF7u7k/Hxp0DrMCWsfGC53BHqw8uNr6w
MBzIGSN8d/gFGgCXwOAuGBBlOj6r4iNl2OdgqbqgsD77HWyH7jncoenw2M3CQGxt
z8Gi76uAuLhOFIme78s0KvBdt84vU/ulAV5MfBjWPVnaw6AuZAktV2eRByw4kpEP
yeRaidGx1uDNJhswpnkVzo6rbkgqdBLqSuXKoBl5WDLBILaEoHCuvitzLZ7sp+cF
f8Fud1/PNzRC5sssvbSkxK8L9fxk460yoFjzm7H6eoHRJLLCnALQKWHwjtZ0rRMV
6EHne22/or4kQXfoyJ4CIzVbIaoGaLWTvMo8VwBiXmPYdGO449mghS38jNYfEdId
Skc25+ZutqdanbR5m82D9IJ6869yCP4s2yxMLFXdsDzUm+FcrPD574Lq3OZVWBwD
X28NKp8UE2tYm4yzHkDNhKA+n59vW0bp9RW8BTpk8SuOwP/vp/PUP6JtM3JjVxdP
WC75zzgEcDFAs4DXD8R/N+QZPQsZoi1guSXrlzZDFBn3SuQ6R0/0uxtoPmMjey7r
g9imXSODIlBrEey6iJTuvmpS0sHxeFk8SyobsDBe+PjiLAzf4llsrOuiN6AWu7WC
k9pJOiKHvom6AtZs3J3c9aJtKVCAS4fpbW0Hqovwy4PTw6vBWtLfMIxCKnPKWF6k
d9aN1j70R4KCsWdFKPeGsmxWMOufxOZcKJVEkTJvMc2SmuD9FfH2VdAAcBsf7Lwa
Tzh07J1eQYSim+BRJW3MUDa80t2brS8qM9X3FRB7WFE90QUPebO7ejdeCHI57n2B
WqipnssVmGz15TSjzhaAF2vL7ueThqg/TERREo3whdCr+26c2WyEQGTTvcyzIy+a
xD+e3y4l68J1+sWdY2DvAYKAiWcgZc1IdYsAmjpIzQLWguxMmIJuUBvmqjio2AGH
v8dBhL4kBX89E1aU4uCFX4Ohq286jhSxWz/Glhp21Q1fEG1+wnSCOGOx0VCiF/jx
Rt3+FZr4NwxeTveRTdBmqsLofsMQxuRTlZPaRK8NORPWbnCNq/G0w1f0Wd86huSf
aV+nIFRAMW78tEa3/PU6w+/Mx726Hn1+2FWMq0rfKTmUpq3C6R6kuSZigiBG8/5g
AIc56ihzeD+kn3E0+EGCh2ThpWULHsWnbA3BcV9RNM1ePUT0A0STTFVZbXx8aU2X
swkhT3IWtufjpC2veeDXxPRwxZh5+N63GVHuIj+xdEuDAuCm0xBsLVIGWAv3NRSk
80NnBH3NvYN+y2rLl+56CVZw12I7jSuaKi3nKpFs6JhGqSvOUZjYlcjqZHWmBZQP
k6Ezx7/h6bDaWckKves7sS4HcIOvZSKYqb/x0ijSIVkSJvTEObRJHZMsCtnoKdKZ
tBmLnbgshy3pSffV3kyfR1ZMTid+ZorKfn3OB8Ax+fY0pp1l0s9qeVsZZzUzQp9L
LpztkLtqnSQ2d8jBK7jpBCUWttXitk+WuyhyS2xafEieGqoTJlkcDsf0BgHsJD5E
AUBvApMR80srqAbVBkQXi+1KKVjS+4fro8/io93Xe0D0nM0Sn/ZSZPCVLofIsFLa
Gyl4Tji68ZMpktaQXOKXGwkmems8bKrUK/Qi/ZxqSE74Q9q+S7Lggh59LheJlkqf
r/fQUVTLrB+t3PaeB3UA82ar/oQTjHgcLSV3HC+WOzc6McwanLGTjpMNUGEOKOcd
dOF0yA6PPw5iiA80ZpgQ4afXgth7H5rTr8MWS3q5b60KeEb6wKENtnIJM9P8PG31
ZP2vhnOELlQnjOI8mrm6mxc/OArzutdln7V1cc+h6qgP9R4LvsJa6keYqsWanH/I
M4Xc7yioVdAGO01kIN6X2BPnmCj4yIP3zl8PRW6DgwwkcMyfuH92ozu0RSTyQ2EV
H7OElwqN8jFYjAIshGnjubf0bCyE/Yyfhm+uj0Ag3Ug91+rIHDYRcJ9AhDIfFYyP
ZHDQmSXJs0IEfYTK3R/LrlO9l6BEH5ojcpLOK/m+KqtHG4r7Kg8F0M4tDXW6wO/f
p03mx9cufLYt0Lv2V5Lv4LIDpOjLEl4teiA1Z12peJs1cpmG1UayFTch6bcxWEn2
xuHlMwcoJAu+p8oDtVmNKsSoFRe9XEuwwbtJuwipJsFi90l6WJc6l97TqKwWyqm4
ORnzf3J48yFAo63+ZBzd8XQMPCqC2LLQ4cy+03XDYVXEyOW9nWujF0ejTQwugT38
lYhDaIqGsQr5q9uBSqyPO2CP4jGM198C0dXpoYkqrYnpfmgGeoXQftRMr0nn4bNL
B3xbp3NMyZQi33W8cmjTXf2M3u9ID5cDbekXJ8Brm1dGEIqwnkHNytvqXMF7q/Bt
YopYX8GukejMVFZmis7OgNgF/meo6viVE7y1ycrf7uuvpz0KcjLE3qefuQ6xCGBT
MsQ6h6EEQmoseEU+2Ci4cH3ZMbnAx5IvfylA42QNV0+neVyolGTWVG1ibor7VQll
UDmg1VbAg4U28cMSEjXrFlJky/9Luu//aK527mYDrk2wc8ZfpozwXyWBddvFGo+n
qAULjuwDGGaSKh88JsnmiIjcArKiUrsEljHKBSd3/yYqIRxCJMNrp2DRfC9mCDgm
2EA70nat+bPIkEFM99G8W9msgQgnov23vMMSnBSzwLDmKu21qQOfXLsLYPtYNbCt
PdUN+MHrZLs89xI4pC1zLSt7uJmeN1TEfYdVy21DRW3i5CBr5yyezcBmR4sqpnBy
i4h1yu6IiCY6jNdoAZj1ZUQG8GM+34e0Fz7FzLpDT9/BtAAATSqZVlKGevBeP4ED
vGdzh+0Hmb4Pc8jdcR7NCQJiL52I985S8YVx4YlerktVnMEVFzjItN9zHWzauX7R
oQbpn4wcqiI2wQkriaHP8V2WTVAI54TyphNQzaYt3BhB5HVLJ+qucGZXtPOpqy3M
/bIZJ/eP7ZHe1pgv1hH+aD4XDor2EVxYq0k/G15zzzOzz6vsWFhp/6uSsO95f1QT
Tr/sLjYp0xG82Ur/JDN1zd2xZKoLc1Lq/3/YEI9c34dJ2xMuwueidr06JRW/z/Dl
YndkOXHWPoGPCoFwARG53qrPDJ92LbF/TjzNW5x9Q8R1+XfA5ddLgdRCI1FxAYdV
DBScOi+rj8KLOjCrxYrHVSZBsIsOL6tGLFHlsT2Swt2JK60/dvJ3EQqegVYYL312
eV7P0pyw12HSZHzd8ddPpT+fYJiBVvXvvlFmvaUyUPO/Ch7fGigPnz+xZzUa3SB0
yQ0ae+FNSb8MsRrzvX/DLBqo9S/0I56VEnu2CsCwUidMv+XRz+8gbs5uT+ZWqUo5
+ohgd5VTDEl3dqESkebCsPMEQ4iSFLGkufd2AB6Vgp8HBAEomH91Rvmw8bQAnE8C
1ADc6Q52qBGHWOIdLFSO+lMrri+q4+ATF5p/QoNIamzPhW4lhmV4HwHJefQ0dyOQ
8Ancd9W8XDiC0HFgi1APHeYWIfMXUTlVVOm0Ol7KDdF95jZ62eyPaecZTYeHF4yT
C5cVf9q4jDmA0v++j6eXqDm8u9WZj2IqyEhgPMrIZpyXN1x6d82tuSvMrkUqOfFU
R45XgFcfukWrIc8GKlWco6GS6VU/l71fb+FNcTnQvKUWmu5Kklxb2M7JKESE7gCs
c3FgNQc2jDkAOoF1U5xEj1IuqStYtAinOdx8/ZWnTolSSXUAcCXsSY4lkWh5gUkS
N2SwfeqJ1G6YwDFI4v+Jkoq/yJMvW2PVLqOyNEeTsn5vKe2OKFUE283kMwcRlfKi
dbTlkl79AgwmeF5sEhKPei8r8wfddL9EKfG0X+EyHrSuN7YrvRVh7sjezc4A+ZkH
OqsXNWzF9KPSfZCRzIlNjBpeJI1iAQIPJJiZ6GTBBVj2iryRLMKbLnY0YN5UXjAO
5RvA2TpQPgS8hCR+lt5AuO9EGPy8FahENUVle7dF2/Db1bH2anQ6vMmx1jiBecae
j8TaejMv3GPrz7RLVKNQby9T3bl9vMF7SruzBjbOjer11Jlnxr8pNrv1MVV6wOsR
26AjgvASNfY/YffJcl4/hJLme2VpNxolrX81m0yBdv9Pb4nmM0yFBMn6DqR2/OFM
Xrh3W/PAMaVoDdtg9M3qpkrNLLg/rv38rTTOBmev4Hd84VGzNcAO7f9La0A9QG8E
X3Sx+cPtZNBn8L7rEUXqYR3q2bmkmZ9HZwhU1tFI1Gf5FzJFKBzhTWhB7vBkcesI
6W+nIZa7RdJWJZKHjA+hp236TtjzDI1gPcq7qIAn1hQ/yqM1/HvhnMzu6SlZzMBf
2rMtSicYQp6vkOd+INZLcc25sy7MKiJfGoOpkWV2lCdcBJ74le4lCSQlms+cYf+c
OYW9sGBGLk/FyaRrOxmvWE5nLWD3rWYI/HODPArbbm4R1sdVoMChXjrj2dwvj8ln
DpzV815BXZEf3PlwGrDuBh0xEK4pJYw09Eanc50uGOhkqURajuNJiW0VOUxPIt3T
y4QXRTEIL5/HEhN0sxo+cjdUqUTcOVpOX2yRczMn0J4hCsXgMOL5fHf2vl/UWSJP
2IGVJkSOAL78bh6riApmUgHLvuDOxTOsQP3Zc8MVLfA8e6ubxvHK/59tda4JPsCa
NlkHGrYAUJJgOi4XEgUmLbVliUzoODCKZKbQM24GvX1NRqUVaDwheMcbQ6/ePuvR
Sh7vs4Ok0Iu6m8MT15OJeQnA9Q0b6N2rQXP99c6jnXYJoaOMdBfOdzBZ2oYLDG1b
EBhOiQReP6Mk3PzLD7MgaGqeplI6q02AkWbAajJWi/ipjfZ+yP+pUIhdAJZj4rqy
SYgI2PsS2KSl3iN7JW4pJdjrG139OVFm17/59BcIA9XxokiHdHkW54mLFqzzfAc0
CbrrWSUfCXLKXNq5afqeqyq2ob/BDn1elRu17mdwxzzEM4Jg9U4F4rwZ/YyHPPPy
El80KaSNOZ3/ChhPlTqyFRcXoSf5Vy9+ksQmcqhnRNUxLxga8pEwTyf1My7Lbq3k
6c7XFBHslONvoGicUX1xjIAsHuAkiVzvEqbQMiNhM9edOmKvqCJ62QR9yZFpNDO7
WzNLwRC9oltWxNzfBr9CD3BCp1bnTsTvY3fVkNjTpIOk19O0bWgCIPrHChnq4o8g
6uPyjIlcC5Uk61PtxD6kLo3yywawDTuzjaFkbx5cz93sXV2TAHY2Eg4yK7/D+zRs
wERJYOgbGx+Qlz5TRduLzpyUW7oHOm3/HgNz5Z2FSg9jyCYxtQDBWSXii8Fe2T1p
Q/4DhUqZTy+6bo8d4rs8XEbxVHMSmOLY5b6LLNrG3SZCIVb5yGkPhcRgm9y8DhJ5
HZSJMQQKaLi/U7+FGv4cvS7z5Mo8u3tNawMNnYmYuOGGdDEFHQ6kOENANM/XMb06
qXiMGZWXDZdIaFeiDL3ArQNFUgSPV23m+2Uyg4yGkYITaGAc57+swHS+iHfZCU9M
viltxjT/QWBksysCfLafIvmfNn0xSBckG4gZQsJt/7nfKJrDyUUFIAcXF0e+YXjo
f7wugZecwryk7CygVkC2xKgKkEOSbc7yicMBayrDmFwevZ/oreVAhsIdu1Qm0Mis
vqDTFLNflVYUl0MmX23Ha4knawbK5Rd0uicZI+sx+etpG/enA1GPwPcwCULxs1oa
lhHjT8HBLgdN4Tro5zM8nmoIOPeX4Akk9o8u5wTg8blQ3lhabdoW2aTq1tDfGO9E
OlQth/CafQVTuGwrLS85kL8emONRVYM0HnIwBlqv61rsTyWSHVkQFXBHxtm5tlDu
dIGQlE92nR/Z0hMnGVHLel6ljYzKSjRz4IIz/4l6jEOOaEfbYcZ1qF8ImXUfFAaP
ZnttNBZMu3hajgrVHF3AZVUuuEOZowPbrUtWFBMUj2eR1GjE9oAg5NTHscn2h8M5
npJGj8CsdcRjk1+04jbdYQb1thLhLiArxhI5t1DYoUsAJ3UZ+b0OkJubOybhKhPq
8pTihzBlPxL9yjI0RxJUV4KPbTuo+QyyxcOVTmh3uoQo/alCpaWKLW3W6q+ote8A
nJk3/ZSZtYeTpMAFchRjScsSO3B+CX7pfmeBq7yaX+r0tHos9wwUGCPh5NDBPw1M
uQbmcJ4dG6kU7+atGo559ItJ0qyGIZB9JLm+ffpSMsGWcmZMpewinfqoUqO9NyD1
JEm41kcNTHy9YNN1zTZOU2mQZWv0IYCKAWfQ3S7uwltM5S8TjukvDpOY9tiSjwMy
1SOxxb1NhMDN527EDdna1WX/5O/ilvkebzogpFeT4oStz0xKjZkaGfmN6qd0/KtT
5RUTF14d5MDQxGS1yhhzPCT/EjaCh8ZhJyLrzUBtA/iXMh3T9n4/ZWXJgBbMDCFy
yVtBs7WIKki9P7VrZEUVxMwtkDoV5N0j8G+Dv7/knfdECDgBvY0UUb+GGi45cB7f
W77PSC8aCvWvNDsDZrCC7F2TeGYbUsTvdbNkBHld+OAa/uvD+0OxZ9fTj59LFHrA
ww8cFSW4FvQ5FjaaD4vgBVvWiHEu9k1JusCn00pqsNHWp+jJGGRzC6DL6qLWuG0o
b054jUQ3DyUn89deJUbPcGpFaTVMGSoht9WESWyvnWx2BrO6SmvAV7PM9Rnk7Axz
R/qTbbs6TusOpT/Lq+zjqtfIE6dnvLIKwPf/nqs23U5HHSwezrBsG7BKregdoQ96
p1tUZ/eUsuqXoC5yPurW0TrzGbEi4hJoSytOOedP2eHsI7vVx4Np1EwcwlsJeYoO
6/2crzmn2lvkstoy5Hs7qXDqt0h98J5bBgEj1G+ohjozz+Bjd6hViLMZEMD1uq9V
g7zire18D5e6ERlxQYP2HR0ac1AmQoIt0e0mUP4nb0BdiB+qHPUDd+pjdif+jbKb
qJyQ5iKrP0kwLqLOpRsWPAcg+V9djRLz7liANWUZMYKB8Sva0rup6Kh960ael4wz
v8uYyvD0oaYwCdLCuBsg4QNtp3smJnV84uULZKasJgjmqP4E4Txr9NUMM6DenShu
i2rP+3SaS67+GMBo/+UHBzpI+6aU0SYIKDk9KkUYzIo8wQjQ7c3YWTKsR1D+54p8
2h45OOJaUe2KwrjEPB7C7EhpV1aGRjjLbs1bpufe+q6dTm6Ol56HA3ONPpmYgysF
e9wc+pPu49NnsYnrQvBqPfXrVRgn1AOl18cFwPqH8QjbXGkKlP/1p/x4yKieDNIQ
mPLbiWhykYY0xcwTSnEhw9A//hSNNbesWaoOmtsi55qFchiuKK0K+P+rFa8C496w
heu36E+p6fUAwAmh4GSVl2+gH6vDwBESwTOxuRqoUA2snkPxOv4f/Ru4G/Gi6imn
+tIeCxxSsanaGpeQ8jklWbKN2TTRh4V/vkU9T0OOP6TLKyKk2Ei0HlROSBcQEio1
FW6D3qfITae8Kp4n9WpNvNC1sVbez+dJNtr8w5GIpvzY2vrjdkUcW3TvdjkGU+Jr
tygoewmo13DF+9ubeyM5DIqinPwdPFfGhowrorqKRYl56urpkuN04VEzY5HJuxSJ
KkN6gj7TTUcn+3LrHXFWCZyrmTxTTyNtO89m5Qe8mjli6Gl1yyrq5ddR8fIVCFNo
gpUR6Nqv5HbjV2c3vbFq1JYqI0FLzOGCK+bU3epEdsW7p7dfrsuSiBVf9YrBlCmY
IcRZz4nMqzfvt1Fk5C0Cy/q8FRve4ByXkm/+ZetolakJnLwmB2yUc3DDqMGPmiXk
O1/pGiYJn7oXbjraQ7J6doqeN5BIkfg9H07sscjcL3n2QBSJaJTcLCMXxKV61Jcu
2O9+Qz6uWk5YO9fsTeGtkWQprmMimAW2gPvndXe9WSwMJgcAqbyu7DKVNQcw7e9+
IpTaGVX5Gh1gfPuLHcfLokfhN7554PSt42NaVQharRbwyHgjauZU3Yg5ZhzwUMqH
MkVGFsgCnRuiqOSY7btbf4h5XSabN133044D/8LGLEfREL/CKUO6aKWcelpiWmDC
729MXrBEehSnnD/Y9dP5Nn472iWPfVz091BwImq/RSRQGJQLd7LKun4jk53/b1uj
k3MoJyncL0RCBvudfazrIHhyd0EcEzPYTAe7v5A7DU0jYIgxbsQ8ErBj71GYkkwt
kxsYj1OCFYD8dP79t2fkZhLtDbrKvhHvG8s9G6busD+NTkmJKHvUHDqVADJMopI4
rA02Gt4XYeZ0eokx/w2gSzSy0iX19nJ8e5xqe8BYK49qa7B83WJLFePW+SjlbMcu
fRhm72LocOqTk7hq0Xliv+oDEKIdN8emtSL68D99us5xOTqmYFIEcnufvSmf1dZ+
AVyz2RKwFUZs7H4oK5g3IPrCeNqGoxvzyNNt+l9zhMGH4Rmk9ULG6qdAZI3d7G65
l6rpbkV5c5KRSyYf3biM/6BVgLwhrAgIe0ZjALCWy1Fy/hSYSjV0QFCQM4ALq3BL
MlDdYomMfNUmkl1dsxdlDCBACHTNNheoNu3Lmj3trlSfPNdS8BGQ/h6qylZ8BDnr
ggba0KJg1/Cls9zII/RDPj51VPn6JcEf1jxALWQZDVSnXSOqDrUD+iecz0X2TXj9
YNhzp3FSMzi4P9dZyLfu8JIuMEHYdeiTRaycmPzj7RCINTW/JpmKzlCenzsfFoGo
lDe8Z1OsxdRMal66c0cdZJXMrhLnfsI+2guSEy1qoSHiTJJhP2HLsAZLFR39q8UF
Tnb27mlwXkJoCRYDqL2MG+AV1vtvDvqSab10JNDl1qCzJmmCxcTmhiazE6NWDM+b
kivcr5UV07z9nvHpx/KXFruFQSv7x3xe5qG1kNVdEhAfNJLnTFkPJ8y0ortEhI7v
hNScEt8DgwLOWEDYtVIpnLMxL4ZQ23N9XFZ89hIcTzJD6aaJcnEW4PvDpskp76dh
8d7furt3BelY2snZ7+yH3Bj1kOGf44RpqyHTLxDYTIgAH3kO9hplolE9cLbWU1OA
uGqitT8nRXihHJ+c4VWXYQvbnmbPxECSg1uLcvS17bHbNsljek1Veza4tZYR4x33
Ct4TNILlX4QgmF8YkYD+kGRbVMdlnrWpUBRgUtc1jRPIgD9poKGcYX1yduMk7zpD
zAhT+IxXzRWMjtVUrV0lcnzV7V5Bks4WMAAIgMG6GkMTBrGUm4cdTRStzFcoAo6J
vFctJ/YtLjGKLfHYCVR6eowklccLqmScViaeu5CXVySjKjxQVAPxc2rABcKl8iGA
4DSR3XK3d27Fv/aQOEalFYK6z0JTHGbz/6j0LbkYrnpcwMzf72N0Qqk1i2Cuvknp
cpXHTUQB8q37qrtFAQYhTVWkNJKIx49HI5qJDuyVRdvX2o2XEgJK3mMMxOoGhYvn
aguRLQLUL/HQ1vEdQPo2wRoWKr44JO3QzHDBlim5CLKzgySIZtYnX346ZtpzZeyE
8GEARqxntpkHO2BoTyFIAUPLS8g1vxFQfEd4sh5d8TNaHzZ5HFSHPzbAeua34QMJ
Y5qkvqf8zqarmPLauxi0SuapCOFB3O4rNS4GcTPzmGY3zIQwGrMSXAt6To99VY/E
Iswqx2B3CpXvNum5oopk01iQK5VcL9kXvVnQ4NFYrG6KJT+ObjxN7BEQ4TAZI738
lZ4pJjbkZX+3f+SHjD5opkQbgw/pxzzDiSqA8qa6Wa0qDhNIzUqWuHBXazaszic6
ptR8qnBBXb04NY+MGWnUMJxlPt3OZnW32FxkXU2Fvbh1XHfRLLjm5a/RgbtaPmlO
Mw2TDtEBPjROwy+TduxCUbxqTZeC3slL4tUg4MHLnwQobdWcCx5pGwtWZtBt3t5I
g6AlDveNvvWH/bscz5IjBdbBeLAvsRf+8b3RBwXq1nkS4/DaWHoL9bdMqqMVFaDC
J1++yqCKOwnn3aW7t2jCKBcJc5UEGtxNLWjjGyE7Fw5HDY+s0oqen4ybHFSYlYnR
K/PIDFFEFirz0wS0Q/tmWTHRtMeVUuprHi6gpgRDfDo5shkO3XDn2Fc5qDNAZXYt
Rw2p0O564VM7xGkP6KDcrNJr+4fo9VRtzIc8rP76cxgsV1NnL4j+7qf1OpTROWod
M3ThROcdFw6diMR7hD2FynLpfQh6SdUgDVVPIBH97yWg9s23TuRwwfrg/129s+yO
1yH3xTjvrh/xFxHfgn7P+CeC8XFJbr34thPfQneqVV83D+KLyWnMGyfJB4HgWo0L
Gty2haea0UOm7yjAkmj41n/hYIwmvk13bkb+CbEMA3tjiedH9PtDZQ7lvXwCV62v
ZPvbGB0oNe9iZb827X3I+dK2Cz8xQdt1uU2+DnasTyPPaQiRU9wWuubjfl2vbShl
HfDxql+MCfBNk15FermUoXK1GDFDPmWEy84cYasemSFwx+RZKzXLvwJBlBLuCRP/
aLBtXnpRzl8BbY1dXOzoxhz8RJKj0MlndV2dVjjlsjovZoxAPDET8d5zNUnuMBuk
9SUdxTgCmi5iH2x7Zzy8YDLctuC1B80EJ7qv6G/Qsqp8RCVxIOWC9zhwORzgVFC6
y9/jELPN9yfl6Xqe4kE7TaHObEN6iXSqYQuVuh9stbequIivfaJ8UeO/iCid2MTj
WaBXR1jZ44+PdOJOmpqmZEZJPtOWMJ/CglRAHwJplc1CTHBXKn+yXDAWPPMNkJG0
XZhzV95j7wfZLCxEeerdSkQ0plUMT9l/5xhoqVhnbiWwd82Fd/KYxUEujXFiu20y
rnBMRieWrhwt7vvS28aVTKPHFqJ81DNtvcXtWlBJzIoPU3lclkrkhaOL7I16IEmd
IdehmGOF5s4L1XAlX2Jv/91LKtLuVi4LLS3570njtKd9c1Qe1/ZXs3/D/h00wki5
qEGBydMGgGBSCsy5tkCeXSz3/HrbFCPbhw92w1x0e9I7+o9YeNFHQu7VIbtXMhVh
sk9Nqe0x+XQp542HfitNxGxkf7XKYV6K4e8QHQxkW8zmV0GhPk2lxdX/YIwMmM3s
MEtcjKb78Jdi84ABpyEAG1zO0kigEC4jhtPomc43FMscxaY2uwnrvHgJoEFadRLj
z8JPus1a2Q5rz+u1CIXpSfT3pJn+dz+8GbXx1j90S8eRvHvvKFlxt0N2HtjPoQup
OlzRQ2T+Jq5XWqT1krYVB9MbJkhaUvok/9CBisDnMFCw9qo2a4tq2VDeMrGnFhCa
FWsqXa4A4qsXgkU2hl+r/sENzsH6mk1NxvNWZvB45oW5d33AW0P/TqHlIOAtOUvK
HHJXBt6yspPnlOgPnssbYYXSkUGN/l0hdPcfo7GZVJgNyrFYVB/Be40LsCTJCFcH
kk6GAJ6VhEej2V0126Scr7fuasT1nrcVP5XZceEYMWdMY8B2IpyWxS8E2bBCt5Ky
KY9nrGnIuFNYKkO2YW9BscaQthaJe1gD4uoZMwGhs1TUuPZQ8UcqCaaZzv/k4Q4b
0HRTP6qItcIgtB8fTFq3GIenvxnjIEtToobPqPXN0OTEwGgJw7X83bBToQf6wWo5
ytYQ7GzVXqyJezLOP8u5OSPXEcbLxveK0ehPInrkOKHdWt1KAN4JAPSSYce0DHQi
lGb2RbfM0wzRVojZMt9anvBJW0tnHk50mC/7Ch8KIX0c8ZHufLy3+Selmt/ISWix
IpTw0CqPQqMMobrM1lleWphF+1kh06YdNNWfXzRMAWd0ukL8wmskBMmYn5pVnQwo
qfeumOMGT/0ZEN/80k1f0KI+MVe6eLP2CVfJmj8LbqToenF+pOf0W9JDc40TEcd+
P+FdvsAcOqeFVhH5mJE+wGJKoNPgCOY19sxroxva8S1m9l0UTe1Ofaprf4V5MjCA
ee7swzabCjej5LguCp2Bp+yptvhkPv/JOfjKMlrklXYAPL4HskjcMywwmWdmoiat
xUu5su3pPdAsubyyIuOLx/FA3PL6EnF7GwsP4AHHp86uXSMfQM25+ui5g9hKU3JY
jELhp8CWg2Y/meOi7ZTiKgednGSd+//zHTlHsyfSzsktmv4pAY6RnnoP4e9VVeBO
ILSmTeBE9mj/XfsBQ5uUxis/p474t3Ra7ypX4quR2brbZ7tNukK/R6TOBcscsPWU
1s1LlkqxRQ7WkDYtM4vivkLU3fi8XvTvXp+dig300gufulVq8rKyvTyjV8nuenJW
BKILwowo2IzJW+t/8y1ZAu5b34lJPTd7w+ZwB6SMBAyIkdVPl54u6kCoXvsHG8J9
VAwgBe8pmYmklEBzPYFxiH0zY9IZpOZ0uY+UAO04MUzjpTSH044yMVJtXtaqil5s
uGRRbrHBq+vrPpiWp2C8nRXprtL/E4flqTPBpCP9BFXhUHTb7h3KxBQmKB+8BQs2
3bfkccd8X1DBhgZ3Jxy0OwU0JlnTNFG2U3tBg8P9x7oN/bWxAWBxNBGcusPdZhN0
EGN2sRJDNH1+5w2zKSufBRnDjcXtVwjOGAi2zOBslscBxNcQUP5OtqvjaYH+oIF7
kXI0mxpQcSJx0cJvrIU/VUaeKEjjl9MsJkZJaSmR8JJ7pXT0kY+zEMsFJURLXvQH
LXuUja3KkQIdjn8In64VmVkC4k4Q4LRe15L8CX0Pf0N9Z6MsrvKJ6xf8M67T4mR0
9MpJ4On/wqOV7vPSrDZ2gylvl3aU6Wzcu9in7v0EzcdPhzs2HiNZmeuGMoLot5AK
adTwjZxBsKty/m5PzjwuDTjqMG8c7KWkJjFFbxXxqiitWzyARXC4IqlILHKVVL0D
dkz/mGA1j+hIVgQnDi36vW6FFvw/o6FFNeOB/qwzBw/h5g0gp5aCtlwOYvyli28c
I+1E/xbd3LUfzYqg5iRQmJNxCYwtd7mNVVMaX9LF0vkTAhLhgKC7RpUeSnzCT4tI
Knhc2IBae5/A4ap4UaJ3EQ3VxJN8IqU4DiqKQ9r/uEZH+TW9COS3CDfs12WykTrj
mw88/TdZlf6fbH12Yy/IC7N+eem+a09x4nXX1v8Z9JyCSlg6/5VvTDJZ5RQNF7iL
z+QqSNHf3kOd8WIdCKaWoezb24DEMq4Y58jKcGVg/fKYSb775ZZ6EFQpy5ntjedD
2TXNvkmZ/Ofo/dVaQDCVESchYdWt2qLZTwsINXEZj0nWLEWnDpqJuhdZn4FPtkQv
zgRAXbTvqKb4iypv/XX1QfNtN7MWUYk75WlB1Hpq5hS0/GJMYF7e/9WBSH0iJdLl
WNP/eTJU81MZ2DZxOXlStw0IGSc/hObeoXvdy4hcKBJ/8Edp2SDkKu2bd9RfERbe
Jii5nPo+MJc7Jmtifs2wtzs4F6hr6GUaC0c4nLUWhTfqpSCax9OOzyi7RpFt7MIt
wxObdAdtKm4CgCFecaLNJylxxbHnvJQBYnAbMwf+WXU4MaNsMg3OHzdmqkeKFZYg
NcP9KWbPCcrKPS5hb9scCQxRl9bDIBzfubGNcvvm1/Gjv1V6cnHUB7cXfc+xsLxy
3IWsHloz16CzYpfL47wNKLUkMKjQKXeIrBYgDj9lcaM3SlWJ6Kmz6xtdG4sPT5Lu
1d3Ba8lhTpgiQYZhcNY2ULWWYekkQ2iUpmuDREeHUlYepnCsS2sCHFdfw3Lybfqu
98aP52RprIhZLxiaFkgShP7bxNcFFPeLAOuAi/XRK8ne8pOxvwcUdJaqWwqQE7zE
Iwy1HUk5LWFbjfQDIBVdJMghf2i9AOKaY7+0n6SGiZK5mXfSKD3+qjlB28pCfsWy
+ljla+Q+rAiIyECr28Gt6d9AFNHILlo49kqkKBesFEsFHL/77gX+HJFUoNGo7RAv
PvBQ0Fh2Xyf4gCCf5ODYl55YRY7vPTT38nSBfxshY59BtTIEglDeDvLtlhwbC8vd
mnVoRgH4pxqZD2mQKxoCBgYpORy9BnoZQh2abdn2Z5+IEJLDl6SHLZIGE+kYn2Id
3PRN5CIEc1rV5jWmCq6faNU/rKZj7tiPhGNav9R6aaghntg0noGOGbGwkZVSu5LZ
eb/UF3DlKZSlgrSqYaEZCpgItCLUJvhKwrbTwlBi9oDJU5ytjTIahawFvSWCl+m7
e7mA/tB0SsBjZuvbtiQw1nRRIzK8Dol9m8dIzmFpJ7CMO30Dry54+8OC8MxGBRtQ
rQqmzCXBqAAKHTvcm7piSHSzGEWEifSCw/paTNyzrdD2uOev0oTwyxuCDkXWPCAg
6IBf8F9YvLflsVCHAf76Fw9edjizXAQSG0XP8ByIJGkO2kaL589APqi5lIBYn3dc
VFO1vEVOsZQC75c3SpzNmLxUf5UVpEDB1xa/OvWUqQxEwtiQzFenfBGQepeXmp0X
xBHxEwZiv9MeKqm+ucF6Brdwj9hMJSg8pMDitgJUy3HqDtChcoMJyP5NWOkP1Fb8
8pW1siX4aeA1ZOudT5gG1c9H2II86d1Lm+4rwpF633vqcT74ud2ds8pwGJgZm7DO
ML9TUPuvx7GCOpxv0oui+TQgv8rjpG5/3AcCkmFc8Eh3wDQIH4ExFpm+S1mGxDun
1uf3MLx5cV5LU9QbUi9WORkA6oWCglavaAfnZ2OFWoOXuCKZy3o6TNvCj/HPNOrg
lWSh71SBazMrviPonZQ3PmqhXO710BfrQLyCI5Yg4uScHzcnt23jUVszPkHRyoNS
O1JAKJaDXZtWCDk7RhPq4ijpydXkSGosULsZ3RRInk72/XiVQOatQudVfkrBuXXX
gM33z6+bnljPoE3tVTPDUeWYh9TwL8DR4sluWMGL9wZKwIvTe4ZN1yoaeZ/c/zBw
WA5Mmaxcu9VticXxSKE5CgZ6jiiLdc7QSYX+NjGbpb8yDr4R/UrJDRV2hlTRrhc4
BRAFihBxjWEXjjnIlQWHUCwX34XgH3z0FuqxnisF72yg1I1P6TpbwuqwlzUccpVG
a2FNNt07Gvm6byvdjqcrQxxhF5q82eIlty5y1eI4GoTutDRuHZ+5UIUKqaAX1fwU
MVTalbz7a72qoM/N93iyqqP240DATsyqlHKM5SNMU2Onj0LSLtxnHW3xqJp+QJsf
P4kFHGQ0i18GZQwNlEl4ZiogRIIiKwPVmJcY/+WzBWM73BlyWEYBPMGPh2J/AjBo
DCIyHIEpyi3MXQW7mKpfBblRsONKbwUeWtF9to2Xk4nrUl3qWepwusYNRT19Jzhu
wIn/FISNy5AR6DGxzIMTgfyifMdevy6od6F4DUzDRT0ouDWo+uRCRqKA6MrTqN9A
FauCbBie+PMQzwqdiN9vtQYq9qaLjEv5wyyMg9mnCPFdp1ToxugY3jbkCut2w9nN
6QsdCqHIuqEL7PtPkQ1AMpU2utbLBu3+lhoElWDsHlO+kgeusQorpKHRmd7sHoxr
n/5RWBIPrLsrn98QBUciFwDeDw7u2lmxaDrL0xf2eY2ETvjx7Y1Or/1cKy0hGo1H
iXn5xvM1u9SKM+KjoTx0SSzkNW26q/DZO3O4KJevubYP5IG6FchR7LsdVomMsMyX
VQaevUgsqfqaOQoqzjwqEdr/J04Ins2ifYMMiHqSnrBWwVu4eMiZ6NYsKyHZQTQY
bF2vES03RR06DesTVL4fjxtwnhYoV5R4yGTSrh0897+uwPn8QkBY5r60XpEnwYRc
nBNqhKadV0XTy8S80/nA2perZYa606dRdxFFbDQ6VMotD/lkFf5S2pPBnn2wvdi7
tQMsjb9uK7XFZYgc020E480DKm+k0d2qsgyyzEzUhKXcl2itwjQh2PlNyMGtdzkp
emdzLwqYuMsCdr4jf2dHZmU/3aEFl9944/7YVWzFAfXE8rCV1CaAzpF9XFGD71NM
wed/DEEGW7Nobsmvy+Bl2cnunSr1iHJIheASsTfqQDZCB20Ct9wYgnw5Hy//uCgJ
KX7IxtkV3qWXnSiUanWcYmyZIwJiSNZ9960n0IuJ0B+lHymxTkHhf2pvfB32rRUz
7xAsWfSmDZ/r5A9LJEsc4HuT1Bz+BkiCiaymBKGA6BAFjxsfAFOMeOdMGod71ogX
s11fZzSwUl3Km6XcNYxVbpkQnpfDylVdv2BOJR/fRxyndHHXAnRP8JqBC/ncy/mA
nsMxnquUhwHrtklJ/rcXFVIpT/dB+iX3ml9NImL9JzClfngeoGqtJ5GDo0HxMBKF
cXSItpnmrXU9mgjY+kRBpDowvtKEweDLC7OXhBWbnTIq/0+q/3mEzpOY9OP/c+F2
9FZuVeZ9s9qXQqd1Vx/VLpG66yZyxUlp+ltoW7JeY0BiI7dqNWBDh7J8J3+eNdmZ
oKHA/tdFlwNObzIsa1CZWj7EP3vlV8NBD3jhvaCF19wZmw3MllkDY0AIB03s3PNo
WOvdomJkZl1fA5ywpp3bhLB8Dwisu8xBUkEzgRZBWJNnYkAYX+92JJvp5/GcPhJ+
da+4fCKFB2JkpxXzj9XfpS+7NwLAiML996anebass/Ma+TnSa+B3WAF1zlrR110p
4hqmalDLtqhVW1sXdD4NqbjJQQPR7AMhLAgX70ZHKUFy32aFBNfJMbfFBqW2nBH4
j18B/GCAAt8anMdeV473ntXvuMBrrzoJOdCIjCyKZRybcy/3r6fnKEM1qNhIgLgA
+puT0GU2Ay6/8WMmravEOgBGJWwcAVLaJQRkNKFA1QHpnUkryogs7tr95OY26lYA
oP/FJz7Ko/IG/8ln0h7Kw9gtFohw9/5ZrxYhs3AMsuAbms2W7t58xJQqTW+IRYdN
J0rFygtf+VpXaqqjhkGPaEj9HWALiotxUhcvnI+aXXR4N3z31n+oungSaQXOCN1L
MKstJjsAKGPZG8xRFGQZjPMIvNO43IvhT2grfjCd8T/t5IjB139jAyrS+CZiUzkk
mMHPg7MwyT4EcPKoBrdqUQrP9D0mxdb/cGUIH0YeHT6tS6vU4sHh90spKgikpxUX
akI9c85cNmIjWeddo4r1pAZWVgJNrAjhXJxYmcF2EFNmbho3geeJ3XDpHuMrshQR
NXU9nJPXU4Rvq6IHoooj3IpUdvF/ShDbrRc5MrahpH78r3+uuHjt9OEdIDhWzXQP
9kh2CAXtir1xUQpHBMeepYEVTnlo74qDZoxKyAGm4nvGmFVIGVEBmSKciX8nNUrp
7y1kArdj+dq7ANBvarU224X5zsH5JIBRGvcsqIR44tWKkS9s55gH57et3k5ZQomS
D07m7y1umM2qhOBcaNnffjDtBSqhvGd4AmYuOhU8r0cGgwEGwwWmHzoNZXgBWBBA
nkuBYXYsnv9cpGh7DEV9HbMGkeLEGqB0E4KzEl2+hKg/KSZdC63eTGA9E1ta2Epi
fIoGszA/UUHKF3JAjJIgFsluq3SpCtghX6erHiK2AsYw+XscQ/KSu5o3aqKfqK6I
4gDMYGBZe7DymzKoJyR/0mqNG4D+MroJDwwRpPyo5xAijUVpO5SgJxg+uKZOdLPZ
0cpTztkMELJXmKLD76Ruo0YeZeYSvYcHTI+pzTj5LyjOReERtAeFjI2FnffVyzUi
kqO6wKJDtnNM84iW/6CyXHUGCsMAeOun/m/FGx3y8VMD4tJiJIJpX/mGGxyU0kpV
vlWDhVV+TQ/d45iRUNOdrz28DALcgwh5htlocSMMLe/T7I/pgTxwP9T8sfECC0Mv
l+rmp65j7K9YT7dHodtw/4cUdvmFWHjD7RrfoiNUwsuzoXUBrN2ouBOhH6N3g7Nj
8gASv0i655QEJgNTirUNgJO0WHIeBK0bSVlHlXDCGWO7O6U1o5uY9A2iQWhx8MYh
c67mIRKFBZg8ofiXuphyniGLb+nd8HnJfE4wP3UYvzfMjpxxuvNBjHjb2dcGEage
Y5qU0M1duX+5cvxSeioP2xjOx/cWo0V5GdXn7tziuEgkg0MjSjK249GqIZNczzcH
SYezesnUQ/LOcYnPP6sTG5r4UqWICvqq964d/cGqwQM2ENH3HDeZeRI8BPQc7oAA
2mxpdUJTQhRyxJtYmy+3W1DYcgwf2hflKZvSUzjxJ5K6ADsijx7F1V8z7iInnDts
tACeb+nLmm6BlUd1ls+KdiTOwY+wHqhC3yvuYuKiiRHFEz1iyFJTFTu3HkJ1t5Ye
KvNCT2Bl6O3QWnIVn6WJ7dtX0FqGK5ruEYp868hZQi1GzLVcZDQFXuJ3e6Ulk6PG
xUKpoHLm9Ea2BrhDlzFOxZoqQIDFIetu9evwG/hfpkyLoqIwItVF1bE51jxJfqp+
F4Ka9GZJGKXFZ9qgdhLil7nsDvWZ+FKgevaoVkPu8x+qrvccGy4eUghI/KV9yBxk
pth1X2fu67C/534e0XFIK8RMA7hHpio4XfZ0UkVUrMOXZrzJrP1CdaQxyvVdvLgJ
OfwydRNCpVaPbg2kiy1dauKjRXrrzNzwoGBe3iFn1mie3es+1u8fHaA7kP3YU//Z
RsDgT/wzX7ebMEtGBbomLRNi0e1RbAyH5WZf2k9qtjc38gZ33FUNHiOydek8GHhE
b/AidAimNWVoiI5NYJ9haZWFNU6WmypV0TiEFZkDkcCOAfYSkPwo51H9A2cTGIXi
gFTL2C4EU+F7OjgnJf0tctHlxLyhpSJJO75c4P74ixJuFJy/A7lB3/xlejQfqCcV
uwEImVaOAPUzillw0ut2iHvBOh51o3A0UZyOV8vXHjgiPPMAP0wynrflMlaJymEc
bvPUm8ChmS1qTT4lcpKe2YIlqgy1AsiIuaOgwEw+3hyxqESD5+s8JvEZvamti3BV
lPD763qxCxDs4xUtZnZYTf9XDkaPzjFGCOMi8kx7x/hBlFCNUfS2kLmBPovU5WZc
8DxrwDV99oEXuYH6D3jp0AMxZv1qF2lKaWDjy50jE+lF8lJ/QJxYK+7f/Rtmye2F
zy6Aj5UFGyM9tHn1Xta5Kgrbc24Z2qXYh4xLYgTZpAIW2NpTkY6Fc3iNL6jTYA1h
8NDCVBORtklnLr4ZZQwGicEGTOAS3lwO6mz8Qhst1ePsvTDenV4hPSIYshQMXgob
NeFLLTyf59K93PXSl3bs3TmkFs4Qoc13Ak/q7id/Ve99jH8N0pBYsAdZVIa6nWOc
zw88I9mEHlhemS2Er95XhUlJQYRhF8Q7YwruTVaCeN7AGfLFYixbakyNG3NMB+AA
fq3NolPUW6FSmnpJ7CEcN4kNMkWjFm8V2+aOkrlt7hWS4E7H0VFWHPFcL6IkzCLT
INJZF0Ngxfpsj0u8UB3PgE23I9F2LLcSs+bJ8xfVEtF3FGDaWcbdixKl5KAo9d+k
BxmNBp8OlFvXdUmQ1g6EUGtBYFZkrgk3rd0ndp/lsbkrJ25Vgw1ajld8hiWpJK/Q
fyYKj/R48qT2mNWytSoLUWgl9tec6E5sClUHNlrk3wwbT3+mrn8bnojO6R89D0a2
D2PrZh7CGL5oOycOlF2jrVC8itgFYIFLrXqpahza75z6boCKZGsWG5iUZ0F02Uj7
jBan3ODocInIbrUDWw8gbQ34zu1Iob/CO7PoJNt+7z10etDg5SBKHHgL50MjbF3h
gWd/o2C02q78rB1L2jb0NnL0f9aA2OIHtK+eBHG0sHHT2/jsLB4EprmV9rTRcewE
gUkvSWsqNRBcYiHhnWgIAZQI7wbdfMXy+Impo8KQfNjawQQp0hCt6h6XC4XZ8Dmy
mekfIBP8xJ5qjqbLau7c+WPD1XCIkTr20fsBAjSJNvGHrUX9oYglrpo2p7jVk+KG
4aREhi+fbbVrcVDXjIN9Lt73RVah4ZnXbj7Zr4CQEYpzo63NxArvXsXGii8YnrJY
1FPmBPtQ1boouXmmc2tZemwnJhwMxX0t3u50ngTB/KUJv2mxRnyES8epBczvr6kW
Qyhprq19ahaz/bISvbS2CXI8EnzJlNoNdBHaYncrS88uoB7Ez4g3BgS/LSA8zFKZ
8XfVsIxUKfkn1Bce1gcMyCrQgAfW1CGdlVr9Xe8L70o9a4nyHAptzRLq0TVnH+Bl
kppEy2FY07uxc1GVYq+/snUkygRSPgRjJH++4jbZxoQkIOIm7G3zLzr5MVSFfanb
huKqfmWR24ZBQu0pNQr2VyTC8Nquw9Q4E8y21UEia2cFpGoYuYzIBKF+QXxnF2oi
47Y2sdt10QB/SrCmfM7cQljXLZ2JrSKPaiL97WuIVjqofGBnrt+ZyliL2o8i1ckx
E4V9sqGkmG/maxb6Sq0x1vsKYksJc3USlGl0pqlOwt5rqf5m/YSsm5LDXvNs0Tst
wuUtseGhDDvdsDh1WPRhg5DEjG0pYvS65hVJOcXjTK0xkKvhcybF3foja6uHBUGq
ZnIyDyW+rXk8895v2OJtNWu/tD+J2H9dmJgWI6MerEcB8ZDtEao21U+THOYpSe+w
4mFtXlGcn5OFX92E03gIA/gqIHWHY4MKG0Rizg8DuK6GRvZvK7xnenBGc2lEqU/g
uIuRrYMb5H+6129xG9ku7tVZjfR4vRUSfJUvjuPq+kcx1Yp7oepEVGeT9KCKJJBp
Mbu2ISgGzIaOsj1RU8PuIcbjqIkDla4d+QLNPottuB9WGDO4A0tzDNQTvENjkJyg
h8VbbLk5eRtn4t++CD7KzxW6ilwlTi03hQv4PilSVGeqrshbNqn8jniEfe9TRn97
GueZs68e6PJfi9XM2HaxoeVyR7sMmY57Q1jT7kT8dgZZnEUwF4CA2KjqeJkkGkk7
Jnqk2meTSkz7d5QejZE+LG8do6aVYzSNG/13D51q3YEb0SJ1KwG4eo1u8BwEhbq2
xkLuH+EXkU8JVcUs5LwoZIORYW+eE1MOcvzD5RSDf1gyV/g0lEb9a4r31r/Ftuva
BPdIuWxeknGKqBif2FFm0pKNfNQQfyyeprpGn8LrbL7dE9qrQMwC2pCNAST5L29N
Coyxwy/dU/GA7S5phJC283wTFG98ZHwSyKTbFiKoTrrBcJU6LLDt4tDxjTRpine5
31dvh2M+AnhSXbCuaZTtONvf3vD/gFR1Wb8JFetlEcFJUy8NPCl2vN0BYt7HLPZY
n00F2XPlJAT1oOxS86vZJI+/DyrDVX4eDzSWh3I3R/rEsfExTllb3aOvhvZoGVBN
JVHTb2pBqE3j3Jf507pIMssCVCPcr805BJHhcv8WktT1lpAvvWQ9X7ZLJdJcDZAK
nMncnhywhZrkpyTi4GLC3qHi5IfW/YIjzSsUF6Kxv9JK4AtmprGggKjNNvqaOUZi
860dxGpxn728Qqx2bGxX3mpNQH5plVmCgh8iXzlLNrt82oD9UWLJT5XTqKy5fnr7
hM5obpr5PwwS8flX7DmH9XyOedFTJvOIZgr5lUIJCQw1OFlbz6qqCgnBeAnKdqtv
25giJqvnYBl1xFTZgiji7mRjTZeBB4JWWXXVbaZZ0sVDTXuVlraeDFPCFzWkQ1sG
dGp3HvOP3eVkGw5rPGcD2bKOCTvnashLNdmmP8QIeZv0ATiKdgVn034wjpY+EIVF
yPvPhJlakKGqnrWF9evIb/H0DTun6bH0jl+qGaaIAF7ngDepVYThVW3JkV0ghk2a
48CkIhuDnlGm86OfVJrpjVfia+4w/lgMgjN+cgs2z7/GfbZWBjGptdiGxsAdO0eP
OK9+6Lf4Ke8dty9qJJpiN1qdZXrhyvT69RrkhvROahsXuUNIkHqaD2Fov0imXtiz
PEzQ3Ncn1PjB0epfkDU60YIfD1ux4UYrmyo3w0S+k5USUTnlO8rdIakPXK0U+O+F
gNe9scYZqAabISUKHz+cjSnee5TOi0cJBmc7NXHRtZ1XRM+DUE1UfyaSJKsr7EvJ
dghHGocrdUXpwbZq/OS5mZfzZvgn9st1fuLjJjNNZRxzEdjPXcenTYzikvKBKwsO
JVUrHlzjlucoV36eJk20f3yDQQNlb3+rqaTsDIXCTLT6TJ0qODQzhrFcjlWMXmM1
jGiEd/9yuEz+SEwyr8QlzGBEUwcIoQaop9UqYBg3989KFRNQJYYtEZBQKP+MEJ7a
+OPQgO65hxBDZr82s/1UlQR6hpta/PBEp+ZwVTMXnikwD+ACVpvcl7Jic+axr4uM
Ax4iudaKbiUBIUYU+FTWI7rkmCx0z64ajbY/qV9EsSvyKOVBluiKR3mi1gcB9XY1
Wk1G3+pvaIIrfq07pysiRZEk9/rhztYM/ZP5g9C0lPregIlLxEXEuB///Nt2CBlA
lXxgZZYq6vEMmYC4IP8/Dxt4K+cutXtVh2sLk88JEK3AIZsfrVuAiyvFr9OW5Dl9
+nzLChMJdzNtRU8ik1sQGLtAVATFwlhZSl8BkjDUqXaHegAxp4FK6qj7Q9eO9VsL
hA8WioO6dga5B9MC70XzDtzbh1U7KCDdXPPopFlM6oMduc/5eOIuWPETGlhIByxG
yF2uDbU32ghisnVwtt5rBL/PFzqemyrgYV7xznqxsVk3aV/OnZlPD9F92kqBNC8o
gMF56o79cY5aggmRZhkJXDvyBcLSAjr4B7SstpAe1DN5Q/gE/ybjRa1NSh0WCzX+
JronDmMxDdxRHJfR8pCixklznYT8SyZjQ7c0B6Kpj8tXx+BPTk2qzFxTJ9XWQuJa
yvX9E3oLHJ6EcQF58PJZrPYa3pCjf80PgTtdQ14RWl2WasAi+PExFV0WiL973VWe
mlAGl94hz8KLoT+9eZh9zkgZnJpBk4KhvZt0bcqt8wd769hj9fwzw8ez5HrItXET
BgLjetpBrkVeQgvj40f8XmspW5fvRCyg9kCSNSNyxM+XpTPLjTYE4vnXN6T1PwTZ
qx0dDyVHe+jT1fEnyqIcu3/nae2NjimqldYvfN75RmPzcFCpj376CCU8Jgw4xE5V
fTVECRhiNsCqld6iiilERM1wJtR86s7o57UTVKiJDpo5N1HmET+axQgF7LVLxMoP
p+NzF75iIvojrno1o6ZJXfKTJBC76c1IOysObykGrzbB+HFq49ZF+nOv1/lXJuf4
zDYi19xDKzhHMpcUezzV3imoz3NVYWDMyAsJkTKUn91ajj3P2bE1AIjeyRU1SfKk
PF0IAFKQnRTj5ldLWd+8oLiBYg5ug+FXZu1eNJdolIgrlQXvOeteCDW7haVU43h5
OrYPaM0dd7qyoIkUUN/6etiKp7rnAmly6zBmicLy2d2rPVbulUFz19Y63na9T4F/
RGtdmN+FySxXdxR71pyP7LBivcbpkFv+6v1bIDrdaM/FuFtfQL+nrizE+/RQ63MU
pLCPmVwBijtUKOBdKnJ1p9Ga4ZA2QadyAoBDWVNX0khQ0QKFIKgXIh1RubW80T9h
t9ze8bkXzw3ygGxzRcKtGDisab9H8+cqZYnWB6mlhoxDxXk8O9+WtIswRw1QNQVn
DIqP12d/JFMMdBWZA4Ls2gDZ6xEEAQ5kJSImpDOr1ettT2M1BEhzH88TeC9Us8vs
ciq/2rl2ouWYFyXXkasbNO3pnXrexXV/EqZFuyiw/wQRU7XCBLkOwH/90OLQUryS
AlkXAyAn1QTgrWdf/84LyauidWAPrAR2cqE7b85bHeEHcCjmVelvADKzNRMTk2DA
zlPKkAsMeXMXicc2IQhAP3AETkP7KlOHUwSM/ufLxaGMeTvGvC5AO1ImQ/bdNse4
tTvtoAIoWsR0IleLjm1R15+53ONgam/A8TWa7nmEFAfl5Lx8kTKmDTMFR89kLJGw
OjbXxk56/T7kzYLBfRjGtIbwag5Elji7LXYfZxjJqQvWulB6Nd1/cwnAlviNLY7j
FHN3NwApM+/Z8QpJ9+rzwg8IsuNeuJY0cBrj+5FgPnJI3gPBwFlremJfwLeeljZM
K4Jp5bwLAidando2h+WD+qOuEEq1Ha228CVhkXTIxrJdbr5NQB0QfAlX4Vgm49kk
n02XfOC74BsvBLL3u7A9XRSvPtbJuyiUsyqhgBAuy214fHmIsfZGKUOFEWQI67h0
7RRH30PpmyHtWuiXNtsL4XlNYcLTJrcz4xJPq+paEPR/RYwxRvAsFYrEJRn8oJ5B
hqVl9IMQbS3ZYmZY3ecpIssjgo+lNqjEoqrQ2zknmL66Y3fKaMtCXLH7pjC1Hbrk
kCyGdS71iQhjWKbV+J8s0AK5f5jT14bBP0NKGm0hjqzi6Ph1GTIn2jVtyLuwOTir
Ly9itnmuNUifnneeAQcp+adG1FEUa+xra31mFo111kk+EK2RoyhQrWuV1JqhJ6S3
GYF9zxzr0HTeyBauirJtqy+pow2DWvRgusxAzjS9mnS8BrhzfKPjF6PbnbGsw+Kz
s0wVrkuLxTyN3c6oQbYggpcRemh1qCrKWnjT2hAEtkvRUJKftO0027xcr8fsuiAl
Zw/jBaCd8FCi+63Zs0Pj6OYYh9stMPnvHVS5uJC1kJ0seDihII1dUNo9pbgrqPKt
Idg8cC0EM5+6PRtqaxpyjXwkVmrzvzBPXFkPba97+wuOXOwFVwnZAjSfzHHeDrjU
AZmkE1HRG7e3LpH4e42F238bMsw2lVI+7jEjmAECe9AKeiyezfXwLpoczKmfL9mJ
eJ9ubA6y1Web0824Bjm5TN4NNQDDjjx+WVQYT5WvPlFcpbkxfEfe8EwVA8J2giiY
R2MpgEdoGOXf9FnPGtfq9hTmnCNZYp07QTxHjPTxZoJcwBhOZVWL2x/dS4YC3NZd
0t7tarOXFqC0kFB8dYObBI7zonwhil3r/7mKkB1SOBrmkClBqJnfvmKj4o2iGu6h
ZzgQKlJwpM3lZpCx7OG1O6sbw1MrstKGfXqy3jVG3ibCn6lqRHvMKS++8DVwyGT8
uf2EOxpz8tSlz7es5oo+rMYpZxc9KnWOe/WcFjyqwSjsz+TJ4TKIW0GfAOYqXeeE
C6Rww2vSbDei45r+01jisB3WR73Boxye5VEdN81NOnNdrTTG645tI9e6K+2GvrsH
eeB/wVvSu92+U2YR+qUa8ItsZeqyU0PD6dsoJZDAt9pQ+2KeKsxkjComUVDrb1PM
SVaAsmC4kJ8E8zT1i5g1oEVtR0S8EeAE6UkL5vyOKIypG0iO4wlQfuhdyRu2huwA
gM7vQ1/Gfzp+3IqJU+/3ls0SuKiVj/rf2rNs+7rgIMnrRPWLgZO4M/l3+Od8XQEm
ejmC+zBgUA+vi3qk0yjzA769L9jZwciZpDpiDptpD0AYRVyZPiEDMLZ/LvYBXvjn
qfI0TldjzSTWS6Qz6H9iNCbL0GLkEckJ0PJjrncwqTZ0qqNp16DBQBpks/O1IdWA
pxcB3Vl7cvIBvIGxA3XgJZ3rg+Qxe07RPlH1uQV2xT9VIb6zfrrFOUpQP8gmlKS3
F117EYbiT+RFOv5pSzFq8O5JcjqjAPuGdJgzYOgxkHUMbfoQ4axZLu7ImjsfM0Bx
WZ71oSJiHij4yWEd8vz8WDu/Svocwt138wZGkFOvGWJDRbiSNAJQZ5Ypw1zjTD/Z
vpJ4N5SJ4n0PPFDAHnwxN2psizJKQl9xxfn1y2VZuRKUbBADL5dBvBn4mXEBzJDc
Fz7cfoa87aHz/6/10UIvnE4nMSzjut1MAyOnk5pjXiq92ZL/oaJ4Y1cJcDke8+E8
4p3yJHAiK3HINsa89D3lC7+kH/w4DBqb4urgMjmyalOIeclFHTCt/NYv6P9vAUKZ
+IIWE1/MYhXTOxWgI/LTGk3lR2ekKRiiCi4FEIazEIk3w9V+/p0gLQVGH2wYkZlz
V62MY7lC5go2xEzm+ZzaKfyC5ld5fPwGBon36k41cEtqgOodLAbPDNQ7yTwGtBDU
uN/+t4gcDSjhfnsBi0r5dJ3H1WAT6/SWmDqXDpHJxKAVpxUM2H/WTAV2pcrrOwka
0cbXtWfaLF88asgqN+Xauvfj+qOTURHQ49+48m1i+hBZobGFKuvrBpiy8w4WKURW
hDDImNxvJGIP0Vb/Z1Z8PLSnugKcGaYQRbekJjdZwR1/ftKl/uoxSogTkqGNyxHD
Gqbf+kW9nhiCharE4LhQ01FWkUBubf6+FM/kFpdNNgONn5WSX+1vINK2kYe9Cgr5
mK5lKC0k/SSb/MXaxSiLqBRDfiI9IK/d/MhDUz81DGEg+684RM6b9u3LDlLRDw+f
HpT+6hxeIqXleGzNfG+toueY6aoZyb0wZr/WQXyjbR872/SEtNOWoPkW4Dc7gcsl
o5eGfBHeMSfJE1ftmRJpg0APG76PdQlskVNq2/M29lPWdYR28qgHkQmp0Tm6epPB
obS0+phdVEbOv7GUjw+xbygLqkyGdY9obMANHIwvYTsJDaq4/ILq4vT0kjsveE06
rDfPShlEn6JUGa82bg3Rle9xvSduC5YrPeVNafuzAjQAmXN3K57+AdYixlei8GAC
pv+zc6o7QFCENhr3nvJ4XZz5rDi0wxWEYBcWCt6cK5f7k+YwV6Dyo14uaZAqE8zm
/vkTaPkdVIvTzqFpS9B97JIycP4t0xwQRtbZYedC4CmW2PBg1uHrH3S9SThOZiA9
UJqceF1n8AyriH79tv1ijCbNrV47yR8GWUjlNVuUKcMmcQ9DwTzPODqiH+EGUKSq
67ExO3s/F2VJQkaB3cKQ89mtsZVK8UoUacKr+QT5O6CagD5TDQLFNfAxbBp/pB8T
OzaA/mvxY+C28dlb6+byoPJvrzt6qFi8HPja/G/pph8+/SiOCjrQFyzxU+nEHqhj
uPgcXgNzcVJjBsebDLAWrmUWrFaxrEf699L6jak5KvLjbqCCiDjRkRdeEbR4T5tk
AK0Vsbu7n9Zaq8P8ywiSPsRDadBSi/uKM9RKT0AcjoTygR+SSeaZRCYVXvx0huyM
hPa/y7Cp03DltxLIfFXTJOktrqqFl1bWjnKvB8F7L8eXS1Uoi8Aechd15+eKyvjM
7Sklu0Eqr98+lHmIdjds9ER+1bHWEHBruW1VlM47tUO0+aKCiNJ98LHHXCBOFacm
PLpEHMUf/oWI38Y5nnzKgbOAEKZUdsOgDe7vPLRm1ahRLfb/hzPCvmL/JtHPyAKw
zkPOsX00ArR0DnU8g2piFIZtJLf5gTsB4+/mh7tfyCYlmPo3TIjToPxvD1zT8P0X
Hk/zaXOvZHnZKh+4VzJ4PwonEsZZTDmqtmy1JRSb0MJtE93kFN3QeEn2avSw6vUk
O41muEY9DHClYAKnlOeuzgwhWncuRF+THwnom8/vVmoLwfPfQEOPxDs8pgn9pmI4
4sH5KdC9tPb3unkjiqVrMux84vzt+TYE3ab6vKvJWwmSVr73NvJzoIas3QwSyGCg
gO/lTi6VTOC1FFREfrXunEmkdUIScKNm3oDCbwiXkQVIPAsDjgAhGxeEnfohLUDt
Zwl7P+nIOGiAvyrZjfU8cZsPTXe4Or+8kAFPWu8yFQANB3IX/6qw56rDgmutNjFa
zxjhMTrBHk8DWnGFDyf2PMJ9gO2RM3u3tdB8byL9MdLlqHhZuFkePXdJrQ5uXTKd
5yzfvizoNdVm8QgkV04esdg/MgpqD+aENdt3NfIg1oE=
`protect END_PROTECTED
