`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yQp4D01j7OPUM2Lcdf71AjR4AR8elCKHImNvVswE+0avIMHcEGXDLUBwbqgKL5W6
BGRpvgPaNyGZlSHKBDtDNkXqFSOAWDw++lbPS6M8137RFpyV0XW2qAftw67NYuXM
5Lt/q+b/NCWWDlCv8cDrWcVA+LO+PvFyGgn2Zw0U8WmFjmcfemnaOkRaIHDMYtg/
T1Gi5eBSJc889zj0YlURCdaI3gmu8CiUBkZWafnDfYdQE3zhO/H/5SaU8BRExwaK
cQJzaqpq9w57Kup0evzbUakOIRrL9EEC4HBkVrpQBwSVImBckIxrF/Xv6qhsd+bI
kvcpaJoOjVIK+NzsDcEg24OVQ/9RA3IkE8IF0EGOijSeNKtLlNP1f//XPM7W/5km
71vvTQQIRqcFyN5Ubv1So/bwaMBb8YLPTgR4G+DwBokqIZhjTW6+tvgdcBvB5Peq
iPPkgScOmjMqw56ORN+gBc7BlXFYLl3605iHEDSu6msN7tjPKf5t0DboafEabu+v
hUXkgiEll+lqckE7HY8wLmiHsQfuMQJielNhfszhJ0a3jRQGjJMjQdzlTxHKjf2+
s+0mZeLw751OmQTIyGT5qtvK5UOkFkyQB2KOw8D7TkBAZR/zrvEWoikqfqUOejcj
Ylexfq0oZGMtrwogPKNbqaafoAhDd3iKiPWGTDDu3DwFuLu4jv1K91S/G4cEmBNL
7uns79a07eErUv3DbmB/DImt1T20N+a9ov9wUsTojCk=
`protect END_PROTECTED
