`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HbvmkaKGvXfaD3HXzGgU1aDfYVRy4BDm29nUaIAHMrRB3dfr8Fw2AJbVtlXALvk+
Rzj7QJGmSQqePRMsjvYDyrg1FCV0NXVzItzjWE3qwC1h7V2uhF9ywoZWjKzvRT1B
tJSswRHOePG9OScFUqu56StAHfOXEXNHzvH0hxMbhhVmatv+r7IyN3BUnHxsstBO
fFpbIFh58BI47CdtbUx6qRK7r0Lr6Gn9E1AoJ1vgOL68+38ERHRngP+Wl3JbbWqF
kclKPMAKn/YXlr93nPDTsF7njvBFaGlnhf6eU1tOmRq3/pRcyhn+GLBK5N2YiljZ
UHVzQKa2M4YZm0eryD0ojXhajH3ow8E2j19QiehBlo0ZKLAqtUkexuuPJK34/Ztl
WSfHy4/ZCigxEK+g6zy3Cn5ZNABibNwdacMoC4/I8lXw3mwlk/LZ5thL58nbl13B
3UvXs/RUs0HemHfozxEM9Au4Xsc/YgvR27WirjVpSzZccF56jIWRmfJbp4X5UfoO
+vQ5F0q5x2vRK4EnNeuAyxN0UEY9TRIi5QdY/fE6rfFL/+wbY41JG180SfGfHbjC
s7hisrScKz/NgCeS2eaLV3Smv9oC9dQm42WWSSvWwb6FLAzNKYugRrWzza7Mug70
8wERGQ7OkOXq11t8cI/+f/BTCDY2rS130osL4CcTrGhD2m6cy+ZzrtNmbEChBk2R
NL09I4bsdBy9VP3Yfv2K3Z5d9Wm9wWuHitBlvelKYc3lyIxw64iTLk4tGcgtoOFO
ZLuapENzplnpEsQ7Dj9bylqkP8m40t87Tpmcm8YkdzROWLMmemuqGUqXt0Y+iizD
sQrBWr8PG6cFO9tBkw9Dp6P2hP6Zy5M6PhKfUqPaCcLc9l2CtU9pFrDtaHRmxvWW
9BrAAOn+slF4LnPzUMcYQrMBI/GX4W6LR3zUxTTWcW+Aput+Q0I5auFjXH6G/1iT
Oh9m4V2xIagpfuZ5MgKN9CZwhUviH5fng56pHu+JC0bKn8lc2UE5hxuNuFI62zUe
tKl+6YOOZ8ysZ1R+Ixl/Ym0udz9fC3SUx30qnJAgyLgUELX+2n+sLNBYl03cAa/C
RshtTerHZOoM5Qxrm3DcKAQodF4CDxlc300d7lew+EybGRwZbQKugVbo3wQc5ImR
/lGMODKAVzOEDWDQexRW/ElDE8Tkmu5iWwnCDTw0mFVn+X+3y75Nl5I48Xq872Aj
K9xdQqcq+5TYvnYR+lgCuewdCr3mHWfhEXaQZFUadCJyPl9riwfODM3Lveh9yx60
ET8yt+N9NKeYGBFDo5TF0xEfLyduoV5P92l6sYjtlxCvzGYBeyF8xGq6BBLlHldh
ZKQOfOUSbbNuRdFUzObrLfaXZadlsk+0v+znjiMYkAhM+syaMZ6+GKt70H4/4Px+
3YqmoI8PG3V10PSdA02/rMhuK4y2hqveg9lWje4P8uFyQNxAJ8ed9vYN1WNnohIx
ni1mdcv6kvQJRn8ThvxQRUUNTeSrPidtFEumkPFLuNU8OfiPuEJlFe2DQopv1Kna
UYqNbgWlJ25Kui9z8y07D65u91qZ3ISSciyS+YwYKuJFjyLJ2DCft0b5dNoZJQgY
Bg2cS8FBEgt65gxaeNb13R53N/IsO1SYxzSfXGBVO1fL9442LPvQa4vSTJaXg968
tdE0o9XuOBHr/GOgweFFLud8gq/SZD8x5hLo6rIzzUSFBuGsx3AQM1TwEXUA7Lav
TMUSqK5bIrHhcdH0Idyk1/7zMmmOO15SXJHeyuc7T9qsmRvk3tOB9gwMVRBwrQVm
/BYaKYBjERof2F2QmMRvHjdHyKjnoNfF4/WbioU2EqSyH0Dv6MoVE6wi+1PH08IX
CF7xMG3R0WZK6irz250TGJmVuxGWgvHtYd7q2iywf23xTjRUuEpbaQuR3GrHsYLg
21nxCs1omu+KsR2GCanamJoYPm3Q7wJvARdlGvA/Th2JPc+cmHy6pA0fsdLA054D
Mh+e5XLP0dF34sUPT6CPxA4JfhGOhkOBJXEADPpCeIwm62fHbXCdXiL0Pv9x0R+S
3uJ+ZICMLB/oFa1Fq0Y/kx0RmXDFIdKg8To2wyNb2yIjnB+Oufi9yc3Ovl8yNaHT
A3UKlk+CMVctr4uqHNGOQmb7Uz3GvihpqBsRIiCQ1qRUmpnTbH+6ac9aY522Et/W
UXmunTNWYx4hHwxpfZU3H4rR+VIubZkFDoAcHrkXA1K5AbDYLCyOksSpQV+i2n5b
FQNKVZUonOrJZvcYLfXeEyPgWppdg3YnNuLXNDpR3h2nqlKZswPELeMb1STzXsKt
aWibiRNWbGdrIVzEFZaQrTPzKAMXcwutIqHkdiRBz11YBfpZQ5FNWh3VTw1aDSRz
HwjJfBJs9q68cbN1w0YGLWDuZhl+bXxNn+ZiPD+SP4NEYYijsoytI3tmVRxfHEFh
eQ1xDBX0Eia6Ol4o1pK37upv/x0GAYHWJ26qhN8zvLprLmxJVrGHwu4phAWSIl+d
VWXL4kdcVWGYPe8jtR1jXDMcLmHHQ2SmRTOs5PriRhquWS6l4Mcht9WumQUb8U3O
h0gRZLFtVnRVErtJNK57zAKdXFwCxJYja+CN+u9Fxo8=
`protect END_PROTECTED
