`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DN+oOdgHp/7tNOG80G3BsyWXjtElYrbq3RJCSbqBFAOAyCvFGxe9ACF1mtMDbe/w
LtUNrxkmdO1Oz5PGHehJfZ13JoeQBb0Yy6MV16MSQEvucUyahDTUNbnY/o/4EKbs
PtRrqWtju1mOPxcxH77rWn6g9zuApoeSED6qjkNsHDDv6nTxTslBdQpzBQ3w3n0m
LP7Ts4K2K+RQ+oW7wKUzX73MsgdqESt7BHAdS6pATPGZPEXeuSzK0yHile/LBHZ7
IsL+5Q2eoLKjtmJoC3mo79UufLFnbRcV2J0Vg3KPiklyt5JlHjE6J76kmPPcL/Af
cBbOvIiV5iNBG+L3JVKHG7SkqiWU2Jw9Zg16Y2Yspx5DwegmyznMtTPROwodCLxW
Sif1nmFodjsXUh34LovJr0BWWpcY+FZ6fOlAuP4UR1Si24Vcym8o6O7kUtFs6w4N
QHWd+LR531K9PKoDPhivwE+Ac5fYeCywTKNKgVCBScLp0GIKVUmbW+iUGfAPFpCy
E38dlXNqb+ruEOFoIkonNmLkv/gETrllZje9MhwROj8ycR0pd0ITmmAdZ0OJG2RT
laFOYKc6+jJ6bjnXCdYJD1JNcLQl4/vIDvxlHOnPrOrqefVWUJnqlfwScyJwT14N
cU766pMdfnUfaf9l7NNJQu5ciS2wK8yKDXsw4pg8M3m+PgZ3MlyV2jJdX4y+xdKk
wGSwXREGFHVNfkHECcXxlTIHUUW/lxVwOEfNXJQZAGtjTuBqkRvuBar/v55D8jrS
TudijSbKkb/VDNEoIYdX4sXvXbHk0B3L+d+jq1QV/KVp93Tb1eI5Uk4jexxXCrSX
W652sSOi7ZNKSW2yDTlC8La28yoK9nX8tfV8W9cIVNugkiOrz+rL56prByTnP/gs
mCztIwClb/6bQtfjWZEO40ksiAEaBu8df7Qm83ssvphcocCfM2T8E5VvNf8w8cqO
NybV0GsPDWndW+SzQy+QT4LsIpKNCKUIuHrVjVgTQULxSZ6nSN/1NpzLAsmoE3WW
UZzhzND8czgUOVz7prWRO/cWeRHkQd4sNFnT0/FLerf2hR2mY1kBlM4GFApSGssD
kaZ6qxrnmyLx6ukzhrlZaMC1t4hQ+756CLo8WUjdkWc85Ibdk73U1vNW7AD8Gh4+
ki33bNBVhysYUltYOUh9FlBtJSyfSPfvM9Ls7BypbaKc0KNROfHg/kPT1khCbSeM
D4GaCdIBhsMBFhxrtAGDw6L/eZfBX4bLC+pzahxhSK1xuNiigTN4wu84y1liY/KP
hqBQ2flDmBBMsLvK1TkjBn/2I+4ruVzcilkCd7A7VJy3noRV3XD2IJSY+DS05REc
d7LGht7xdVmI37c1r1krru9PmQvTeF9HLKn9D59SfzA2Ku/ECzkMhPlNdR3CRDRu
moLikwRApzk++wRe4NtDkSG+ZPSrmIKZgSkgBJRIjO6Og3HzzUXsIYYv8cHKdkZl
RmZ8aRpMSk7Afr+GO2q0IjdwqqtTdTtvpcl/vJ4c4Tlby/x75DpiZ4Lq0Q7ifwJX
FXC8xBOzNraWahJfFV47aCgnIRF/VjaCUHO6ketH1jB4OaQ9xAL+/vjEduGV9izL
JVUl5mhm+2Wgazd6SfUiS/ESCYMGDorukgT8N98bsB+uW/H62PX4/WN2TXSdmyUB
2Alrx9eHJiwFtyk06YG12G8sRilejXhGHZ/DQi1nHE/R2i2erq9xTAUtjUoB6WLW
9Yo8kkyNKisEqprLwYn0xyBOuOOCCCWsXYM0dLTCiuw68ZYDmwewOCCu0dJYlds+
aouBrDzMnpSAmGkmqMTmMyt6BaCmcNRM1yVZKNeSoA4XUyFEgvAEM/4BPKVBBuKI
okHMFGFssfoJE+puf9rxiLu/bdJgHywjhA1Hc83axGT/91Y3zbQM2LFxskRW5HK/
HCSK2KXKgE4Wl6oTImXMPL8wgDLMLfGvl6wgRT3E4LtbqGcJ/sK770ftE8ne2Sct
iuy22OIoDK/WNl4gjvaphpAu3t5N7QbEsSMkv+zpsZ3sueibejaciyp7bHlgOy70
tqRArKCHqtOmqGvYh9xEpGJrYenxQNX8sVWQ+v7N2uhPT4pYWj4TccxyQ8kWTyVl
AYGluzN0imz3Zk3jQNOOdJRT3jZS93nTCcCImUHWGtMRTlzrRzbtqwl716xQyZ/n
t2teHj4FUGuesdS21qeQ0MGB+PPNhx2NuC7b/Jf76u/lXsfTZiP+ptW6XA28Ygoy
xb2FmJXB2WzqitQdJu2ADttigt/y+Mg8LpITS/WgTSJ0YYWdz/iPoSoAtyxK6lyc
vENAcUboCZZ4eopapF4hY0si3WxOFAFuBe/55g4Km+0T5AICQok9WrpepP5O6wVR
FMVQFzP5mJsgpPq4pqInW89WCXImESM2BM+da73Zl7tAkwBZz4RG1jkB0Qel6BCB
ReFNxc1kjMcZ32l5LR4r7qINdzO2BHwZ9YmEIp4bbTLpW1VzhQ4GgfytxZ2yjo7R
rHuJIzjHQ5H1YdSkmUCj6MbjG8Iawzpw9uw4Alu3XwkBlowtSwCNhWXDdQiD2r49
2+yBjN6qr2rD65qDG96sGIFowH4ruxu6mtjyQYqzUfmqsKxyDlXGVlbqpnNLFaMv
dJPcNZ6I0VV3me3eg9VdDVdi0uDADvdPAWh/BOYuGVLJEEc0gp/B91a5vLB6ybEy
EKEvrjADFgYnrV48oU3WOAJlQo8cYOirBLTxjWd/BBu7kfaWgVpVGSi0Pym6C6TW
ASSPBGnCMk2uq0FIFCenbXtVY3liwP2uEvjywTPCCaXGhcGAy5qyGsZpkLx4P3b4
4c3CMfr985rkuFEZMbOlqusEQkE1TgrSYjBqjFd/4BMhAd/k/bg90u/FzyZwUGPr
`protect END_PROTECTED
