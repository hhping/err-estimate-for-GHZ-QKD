`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bSYGOAmxNwaw/sVJobs+SaJAxuKTv+L4hBn1nWU19kUr2DV3ZiEPZk5un80DmFLR
io9fTNJWxAwzXVWe5ng0zv4ONuv/sERajul5qenK6712ExZH4nFRbJfnSg0WvWwn
m1ak9zVEURGPYXqx50Gt4fWy/j2C6TyZIiMqmp4MqtUXgJ1SxHXaeOZYcZI+Z+sJ
69T3/JKLQUWidpIPsao1X6v6Yra5Y55soXBi1RrT1ZLBcZemJQoVOO8Qs/rMv/ZQ
5h+biDAakiHZR3lOfNULlw8cNfFny8vtorZ5o1PtrESQmpE78+3rSm0tNKBFAIFV
ZQV5/kzQ3qEK706CmNia7mvE0i9Tm5nPfs+Gc8xQpqidtDVmSwzE8xFUtg5q0LZ6
tVIfVom9g+JEGWmnGXyNhs9ynf+jv2EtBe2N1GV5ak2E6pSOsX3ith8UFietI/R6
XtN8WYCO7Zyz/Dcd6dkBRifLGeeSS45aAvLyD0Ap8L6VSsAYAdIUda4i/G2ByjsH
aJUINzhqIh/RxzCRceo1g6gt6Nwih1i9vP8yuwRUQjpTSMufFOWu6hef3mW+Z5/m
WSqzJfO4Jdt0EPLWqwe7896U5x266kKyXisrAoYNn2Ieew9yCiQRN+2KdqsFZp1C
voIV3RGq4UPjJrcDl52GQtzGvz9dpBV2irMoQRaAMccocGta16diFY1bH4JNiWH7
4/q3O0l7o9yPNsDyboxWFWlgObV8oFHkX1hrsNGfzscyB5g0Wu0/Lao9ju1QuKEI
+Ag94sk2uLwNWYh7AcRzV0ro8/8biQER3To9+FPaIVBlYcVsW9zQWgv3HI5yX5OE
9ZgC2b/SNrB7TiJ6FqBvFp1wuXZzV5mim0mBpItI5y5SnUz0tCDMPKJ79tqg1G4G
SxFpghqKvLlj/b+WPYXTIcxzAg68I2gf+ylmOwIFWB77qSqN/nRwaKEkqQ92z1DP
8r5OW2XNhDeHm2r1qlfOsMZi/gsz5exKTuDMVBNwZSKz3Sa7lHO9NhL8bhPQaiFh
Nist7JRl6mAzvXYCh3duIjC11i+5ItoTdA0Di9CN+nbukuQs9VjvrqDtpalMv2TQ
hffFFkTTCihcWxe1Q29ev7tBUgOB0eRs8dCjzXrvbiibksqZwpSjGEvMDtYHVwwR
i+SCMhWIddjwSjC65/SZE2tZKS9gS4Duo8OJmA/IIU/U9GImevb2RfWpxe/RqjWc
YZ5E/pHSt4Jfeyc0u7YZH5jPwTH92a9HbDRCXmgQgRx6FTvELjWL5NSVOG0bUh8m
FTrL6NecpRMaCOELk5lMle9gOaK5ZrGF7/75q44RK9QlvObNhrLKQoJP1EKoa/9j
Kr2Fb1jng2D9V7VK/Uvhkft6KvLwgUUfCb8SyH2Q8W9LB9OoymrELDS0ZaMBLKpo
nIIsw5UdRk6B9PHkj7emxMbrJA6PxXTz89l1h+5a6t7eYLSVmjjr+a3AWQOHgBXG
NPPFr5OYOZx7Z3PkCRRsbJLzQadm3yfqViCWfu21WHZQxbfDh7LyKxZtA2BXee40
ufPS9oiWBPIAL4eZcT9B0wi2IrRKZdhdmrtWRi+HfD9ThqHeLhfcFaXAFqpPZ3WW
Px41tUEJ1YVLqPw98pyRECxfIRAThpUFxSXeQbFOtSqNinyNflts1EmWv+lrsHgl
NEsxmUr3+G1AfqEi4vgnmqupCPOa5XCk1ZZ9fMLX3j7CmL67Vp2TIMnpg5RVJfOK
WG3F1IFOubQqIr4KzsnS0Q==
`protect END_PROTECTED
