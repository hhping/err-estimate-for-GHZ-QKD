`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U64D+iJDcUhyqS1MfTAI/M5VuhLqk4nd43pUgXb8DwxWSp5OeVqVc8JOF5TyH1en
Gp8DE8+U2joqEnO8ePcAz4SxPJ0FoxY3jniwnlE+fsRN22GBsYqeT7xzMzCXiDKM
Z5WXST0yolTmbpE73H3T1Bl7tT1ncUM7v5yWxe9SmEu9gWmO3eZteErHgjt4KZse
bZBoLevtnSyF933DaQJjm4M5S/CPY97tr+ZmuoZi0Qeg78NfL6CSV0DL6m5Ym8sB
46iS3M/yZ6041GpZZsyuO85Le+4sXrpZ6sjar7J3UMEydFp+/cIu+x9/g0qr9tKi
8EGTG19LTt4hK6DZNZgXrCgYcdQl+qHp9czR77ski3PwOzfNrIgG3zZwyZLUWJlK
be/ugBGnwBQIZuKHqdv+XQ8boITnrgbNTywvJCwD2hFey27jHW1VsrNPqooU6ssV
VyZev3sg+fyeTprWfJgq41BTx8wIBTsncvk5ZcuLMMd/Tc801P5IPvKN1XNrfQOX
nlLmcKVe6a1zC0zxUSK8nezozG4XiqSsavNEXOFhVwszPQ8+jXFlYRQBxJy1kg/h
4f5zlW4dreiRlLoQXurkzYpHy7A+ZBEa9G/lAX9UTWfhpyFOBwIF30T/e4kk22Xu
eYccZH3yUuk7DvCXmjkKV30yu+vxnvw4d78P5dr3hyJyH9hehtTmEvONCAjkUxiP
M+fqCk5j7o6eOKYb1cQKGKGgg0rFaZOyIs7icR5MzDxM+dCg0A79UXsPcwujtaZL
`protect END_PROTECTED
