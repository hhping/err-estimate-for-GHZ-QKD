`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FkWpoOchQvj7Uq2D1BB+O0YYgNxitjVDhkZoFyEeW1pJ1sLdwx4NvzmrVPh74zXk
0/iBtzHqAP0CFaV+tLlU5bS15olORU9e7gpuHUim3lHxpRQDe0USyyY1/j+k8H0X
JZ102wxGDjh7afN4uM8G/Xj4OcL7GRNbIwSCjoERvAn2iFfVTZZctXuW9emLpRDh
IVEK/PTjy8iEBvOApinYj1S+wPiGjJgp+d3+ocx6WNQ2fNYe0jgqiTU+O6uT/ybv
fDGU8CnWcCXTeiAU07G/W5yXfhiqemB3x5q7CJFmZrsTB2kDsHIkJJFdGWCuFGux
Kor8kHYdAHc8dp11rOtXeJ7Y123GEf8O+BkYuri+Z9IG3BGoMTBoW0nMb6AgJlnl
boq7Y7KonXe/5rULHpA2UOrZc9AkTSIVGVETNpfEQt65EPQS/aZ+5lTDrFBkZsBF
NvvS2SYPtbmf6GxygtAuqWWUZzmFVtXdNQ51J0Umrrz13ZWxpfTn/DFrESvQh8og
mY6D3Fzi0/6JTMbe/NJyuDVGhFuzC5VKC5uTfFYQDfZxwHVV5QW1SOYSmJSHUx7W
g0q7LpwKZDSOGFBYNSolFf3mX6UriEFeWbNk36cqmYMU81WIbms0LuTm3ZG5MbGd
64ezFyBovNeO+c8Pi4VMae1MTP5YKvgNZZ7qrBiIHHEocuZ9S0mts27mUAg4D9OQ
xEOw4RkApDfhfAwOvGr10LVtq6CPWxYf5HsQ3786EHSIgVD6KOpDDL6PAigQ52YW
mtitBIKx/dHD4qFCcacOkbz5Nf/YiAKLmPNlK8mnNfknZ15zQHF23p5noJPGGdX3
hH+wNhf+51GcRYDRpKsC5XdgXm+anYuzu0gkgDbtaW/IdOEPQmZMQ3aWJHVNbw1e
pvtXKXy/XqQBlSrUCKk+ouC+H9Y+w1PW9qBsiZ3A60L80vZw0Pjq8hbeAZqSn0Bs
kUap6rJsRn1TyhK0I6TGBuW83T9fPQ7TCKjkQ07041MckkZkx+RgCBNd3mIMSnGO
8U4HPWsOxPAeP2E9LF7JLxmBr42sHEPmy4+5J/iz/j/NenYJg8kGMp+WVHeq27q2
Tewhpfh2AjVYXpgdF0TtqZG+2eTLfzInZW+MOgH+Zv86N/p8XvVYQhBue3746kwp
W2Ry62A4vX1e6K13J8eUb/v2hpOqwyfra2p6JHJHDeAg8950YHWsZYEfrE7sQNNH
YNRkzAnySSFNEW7aWPUGqlqrDPZvKIZYQLBbSbZFUKnOhNa0XEkCtopoKhT1frEc
7ISnYGnPQlM4RfBLN8664VYbmUPjabqIb4A+oF8ZfTybI3BfuDkmsnmTzhEUlagI
CSKBtgV5N/vn7SIV/uQYf6jG0Gi+7kE0HyqCqXDnoL2/n19Y7f4b8fkkyHVkSHS8
7JHEwRCQs+dcH43OyghsnIDvxf10ou9ZMxoKWKVQ1oTj2oWtjM2NsFdfH1PcDLn9
oK9XikA+ayA4oJU/yBzN+nfk6Wk/7gG0aYZ827Kf1hjTl3W0ZFV7hDMGyN6m/kch
+zSsq619q9Q+eu4jBt4If+wctcxRv97baK6JEuYjCg73ah8R3eLzhLRR9mIBxg4Y
SbipndAoGbeulsMQt0RQ3OMkK3ARHiNustCYqzyl+2VoUqEn77PbIaQhFEDNvqe9
Owbq4td2FU7qPCQjVMI2g3hWZG5MJ3lP10lTuYj8wme699FDAVwfbDYcPSSKvCPS
vIJxLMPDqyoarHhP/hRwyuAN0pzUE9flUndqU/qLDjyKJvNvAcO1U5GOmBej/Bnd
G4VIPwZflPXZbjWLdI0L2BfbCSxRZGn9gQkFTOJStcRoEYmTeTnW1z+gIMSKoDpE
Y1oaYmZN/i7UPrsytuDKxQuOqska2eY64waHMrdj5WcLWWuBSVKMFI5uqxjgrbGw
E081MRcW4VvTVrv+PXXSfmoHSvnqj4S+/9p4CaThLtTVRuIAnxz8+4itZdjOYWb+
J5t89iagXPrV0IXXdga0N8/BBpgXv9/48cYFrhLYO4ZlYQiC2NjsL+jznfxYmKP8
/G8/OnrPJyeeZ4bG/qL/LAieRYn3ylfLhMQDpTo64PlJhdYoD3XlQq3/n5ipF4q2
j1Kybc+HMxaNGjivhO5icuIDqhhLZhR1gEEBhT3w42Xu5yHXoMnjNOhLiwt+x3/4
qnaDUYyrKnWpgnTjo9zb+BzyhK9XAKpKUXdVWpVmZzyIe+JAK2sa3562J2DwBfgl
RczEhnFCH3WjfnQid51xLQBpVrQU1hOPZzBOtnTmxJVb9xSaYZ+eCZkbv1T9zLj8
ykxwxy6fcZP0e3XWsXVKu354oRZV8o2ZPW/OT4gEP4pGwazk7vWLq9HgBF5QbJpK
N1PVKF6aor+KsK2xqiep/SzdLeNHCplSYH6eSJFn6Xn9xcy/hx8MAiiSoscqVGn3
GRvZ+T912+mQS0Un/YuLMBVcYxmujFvoynXzC3P3pxeu20Tg17m+npKkikSynLph
lxH7T35xHM9yfa/1Z4I/bUnwmboYi25Ne21Ij/ZhheXs7+1g0OJ7Ppwdzt6j7HxS
sSrcIn/q3GyuVEyArAw94YsvFdz76Xq18RKP4qtBrD7w+TEpIF/TODOB2xsoL4DA
WQW8NoNvW8xt88pA/FrFnalkdz99ZQoffB1rI9Y85388NCqeNdLDonk6j/iwBx0H
gP3utWBCIfqJ84atdIg1B5aHa37NuPAG2bZdVuXtwCpZDqdWw5EDyYiUJIGbt6+F
uF03waqbDGqHtVlCHNAKrJqvmlLUvCSJHU9raVpCy71RYIgNVjvuW1O6ROaRa1I8
OYNDZCqZhnNg6hY37QYOrHSv8jQP7Hyw/e1gm1zZrFryXJpKbblx+HYaRgXR/0+T
qJdazFSXnrlp6cBD4vY9yQweYlhyyjm6h08rw0bLiVSv/P//K3b1Zn5M7YOEtzkv
xPlGskvFQKxWKiT7qlGJLMWg3Rv7r9hR/esBCFuYeKKsajxt2XsSgTkZozMF0y2h
A406Lrq9YKd/jEMzYQY5c0zG52lhAl8OLfaRzzXAMMKa6Ewnd8EGiJMCiEoom49v
/fOQ3nky8zazPU/E0f85VtzXVovE2N+k47Cdv3Ziq6scaWuorlpDR5PxfBr9ssWC
sJIz46T0RLJ+xkc88noPec0szEiyMLiV4AdDOHZkCGbdzg+RbbcvUCn7uAQRCa9Q
rZD8mstfgc9y4lyE1VkO4NHnOtyFAcp/raUhRs+46vukdGpwot/pjSab+eiYnToH
UuL0uA4hOjCpTuu+N8O6ZGIS/xYoYZs4Loes6i/ghMJ7jnFILV7U7z1QHkSD0uxC
LeNlHkK36uzNxY0AmySkRbn4ybSmpK9qY1mW/wcvYD4rDAh1sAvmd153ENcS8/oq
f0gn7y1s1IcgDfKLK4TUhF+A6PqJQ+4tk6ch4P5EGpvYKk4HI1gqZsjWQV6Lf/lT
tm6vsHJt6sxXAetLt0UC7mNqwFZ84hN7VB0pOb/2uqCwnQcuB8+ilaw2lN4lxSsG
zMM4dvmvUyyO0MT6YEFzy1L8+iuD1h1Eodf/ixXBYsEwbjrVnUd/FRTgp43ZH8cV
2GZ23wE3LghU/m5tGaKn0uvppFg6Ou+oG6Oua8WQT9akOVolhBwA5u/0cQPbguaS
HOHiu9wmBIzeFoWgReNzSWEMVeTFROZs7nw4JE+Qp7fJQY4tDG17G6gVr8KJosFH
UFh3tLwpkpCeU1G3GC+j608gnZAYfN/OpMEzBlv5wD1kRP09humbzsyinj3kbU6J
0k6RRV0treX/Sbjs2yc0qypM6nSdLUZssVWzL4FZVm4SnyhN8CbEQVz1G8Kpy/pF
Vnv+QjJkFRCytbunC3h6yfPRb8sjItuChYctjJ1XW7IlT7FcHMMwP0Qsp6F3Yv3m
eGnX19T56JyqoGVyGoDsmvwXlUPknnZbt1DcyhGApt+lchst1nTtQiKFKDxMvEPH
TBrIraJm9GtQgewDDRsW0zVVkwn6BMV5Lwpy//aGRr5RcHQJMr8GdbbFlhrth8Vx
XjSQy0RYfLtXp3zpWStbrrL6rell5VAQK7xrmfo+NL0FDBd0NBUttRmZzsf6YDY8
lWNrW3A/j/vY/ZOpOEtYSlTTIoipJ8w+b+mwN8aGzbk/Jzrn/JLanVBlPtHKkAwc
cO7LeFDN/OR/7uYNFvviT8jI6fhbjGGkKszuhqnY4ygrHK8fCq0O0zK7XKjpRJLZ
5CHEBtoSL2aUwpDeq7c3BlP3VFSLtt/gKAPDVXJr1N4RtXr48BEiGOpZRrhF4uhU
C9Lekckn3S47bieRIb6CTJbhGziHwXelYyC82IWWBTk6cpOyvFwoJgt+R6vTG/gm
4PgF7HqXdLT38PxwSMsJALDDlGG9KXoyZLEL+bzm4unyLD0Ac5itQ9LyI1QxewJs
VHF9keCBAkxtHanCe82pDEPhnaj5rOuWC3lB4G+Lq9X/4c4At6qaZoUGxJZko1QS
AOY77JjNQb6IhkhyD3RX6CTp0RRYFVbm/nST/6/xz/LLoSebrxyTnQPGn6KcqIZG
QS+9jhqqcX3FUSvB45UdUuQmlKFlA/0R59/JS4FTx+THb5h0nBq6oa9eizrpVcke
iJNUIKXpy0ipX//CrA+4pGc9yujBKgytS256eqjvySIL1J75/ytNFCoLDXL6/jbv
4nVT4Y9xIxx3S8MLzylMxOX64Hi6JIOKkhgeNauIEXRUxPwqtXgV6YMNSocGZ2Tu
SlQVXGVIVJyQg/ZzxYCXecgYh/4/STTpPCqF9GRJyhEoEBiMN+cdzA/pOETMRwuP
z4z38ao/ch9hzxIKkBzxbb5mmAxmbPbWaLKzdcdmZ8dYfisKMxzuUEY9flJa9LuL
i+dB1taSzqieR0dzHAc+m4YdRiRStW1OfagA1QmGgT49SrCS3DpoL4G4ySy+/MW5
QkXMHxENxDNVuPrEvd27nya4sLrDAFExLVdOr6g+DWuMNsJtQK5cekejPo0Ca7Dc
OD/Uh5EK6pae8JAAVrA3wqPb4ITronxYqrIrrNTcBNLiIIyXmrOUIG3Hxyg660gi
CHAhwW5TQO2rCQ6ZAkN14bReno+Vlee32x7RVlTxC7fC/69qNuZHJJWoa6yayPv9
+5V+pUIG2J/f984MerEOFUJ9p495/Km/4jscckTiK5BvPzlJ8bnHO+whjHVJ2sZf
twHgnP339pz5ISe0qSXAkM04tKsdrbwQ8HYaMcnhCigPXo7MvEGpbtH9YY//0rQh
t5GW4LVDaOymOT2/VpK1dKBcL+zyvnBX4N/5ASAoT59gobyiSJuqtB9xrQwCP6JC
Mw7xkHDnyoJswgrokEwi+KbOfBgpcGEsjhGyxLoJKhS70IgyZhQ8DquzSJZk1sjX
SevTUaC7+Y/J5urKp6IDkVu702nykYi0syPJ+XEQn6oByO+/ztPY/AoNQZ+Cua5d
sYZaiuWujCqZHPWsVK37w15Ul2CXAnog6q7ffCPWRwQlS4O81tykctr67TsC1oQE
R0qZVXaTaDHA4YsiF7xUPbKT+PimQczYjWZHNRZ4zS6H29eHIOrsWz05BjkZnz7L
S67nmQgy6cAWGpTQ4AyTYtrStY/lqrWqEok21DN4LQyNslxxkc1bGRI0IjP1qi9P
8cKF2jrBKi5cUW/6+VF4293hYjlM+7TFjQydJAjhKK6F9Boa6e7ohjNQsXbskLAT
ixJojgPGX9F49IjfVKdoNRMO2YCDi9WHa6acVVa2SEhSLlOFZAnJbDd8JjvzOJe2
KQLbnxs5j87pMgX7yQ9uFeEeXjXe0jta5IirgdQhuYVMYoc7UmKP6HQqhk6Rn6bd
m1mpCKSpx3xG9mgVrKnBjXlhTT+FEgfqXGVd62zhqsFMJieR03D/Ghrd/vFmoyAF
/QH0P12B02sibelitY0jjFsbIdkBQbIVt9mEO11EvBDYPLmNk7V+qVPIRX2C9xty
4AsjvfzpbVH6gc2VzerHN3b1xz9bAKGiafwuosWZ+UvITPOImKyuY3cLkbr1xxid
7j3LIVlOk/VNvm1ulLxL6HFQJfKm4mow+fJLtV8hyCrEx4fPLI1Fw4NGPbE/fmuu
gfD0pgTXWmbrPkfWlDyMCP8kvRLU2yGyv0OuRzd3LqS3AYH2qoQMgdcCkd8ovyOp
cdS9lw6coqnaqjRizxic73epp6FPfF0ZNBswdQSDmjmHawUaeDVQYcaDW2mBhDHF
1GGI6yOEcdGJKH9o9n3KHQCHU7tbPy5BMg75lL8iRXstEbKD/Sj3INc6klPZK7Jf
uYRKb4itnFCLayIkTcZc8IwzWkbH3eFHligC7FNpWmJ5nzxidU0AzVrtDwSDLbnb
FD081O5eOREiHFjCP595eBZY55Td5NqGT+MD24hebl8N/cSwgh8HkJq3fCc+ofSN
LbTH2uzS2xSA5Qnazh4HRvMvd8bIvr4mL+jyi7M53F85isBhEJBtuzwTaoGga4Ic
YtO3IfiwY/oSRuqEi9atMtPvTjiTQZbKOrTt9cP57Nx81UuKjsCrl0o+x+D9+mCO
PJ/mMtJ7HpPYKqKVfKpkdB/yccjfKRTpmhNM4M15OT9Ks1bvD80FTqCGhwflpYUe
crgjQhLo26/Y/fIDlV1n8QTJe1CMDmJ+vZglbQocQlkHuJBHVpEIiRqhwfpZ1T6n
ZSW5FsaEz4ZWEjhhfO5PlZsZzWwNiW5fw1ECqqJym4vH7C8MmPNx5G3pp3H5oFyq
Z28CMsoEQfelodpizbjCdvNnWzAljAjwMEfcr99fOOyb1zPskGbOcYzkcVtWVxiM
Gva/VLDuoUKMwJDnK04sqewAuhWsJ56n9xBHODQYyJTp6ftmVfZR3VplzSq5rm+M
q2euvx4hF4Hm81Tq3VKjgigDxg6a4Apdt/zDdMB5E4REQHQFBWd1EIRkjMZFolvO
bdrvFB2/g4ObWVmGBzyJGzFHo8XtsbLF51MtBhROW8TCb+Wq7R7KRev9KgRI1sWS
AeH3gSRz+s4TE3gRSuNaYkHeGfpJa1Cym2f5qZRvgRaED3PU7hojt7+w9qHP3g2W
2/KKrBWzDs0tXi1xe51YGEMXzjvsBk6vkqvyaEQZHtkAzJHHgaHPlZZexDXVL2Va
Pz66Mpn1jEAi2ZyjTpbUQw==
`protect END_PROTECTED
