`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JQ7H98b9c9+S8Kl9srvx3nuKf7w5BjeJGYzJ+0nPyawDZ32od6TZskj4UpgDZQxa
SvAqXS7HO2BDr6L8McbzzoEY59xu8Q0SZPUeHM36ecXjiROipOp0y2f1Qjtfn4CV
UckbeoATW46Hd520xTqW1Jn2pwZsQ/3Nsdd/Hp/I31jmMQtAVX5VXEcPVcEXhjON
4VxDPBeSMwDb4WElO+yLGwsurdgZVXJ1ws34LIx8MnvcdT0iLPLLpRlyrT93p/RD
p3lr6RvDuGKnG9xu8Av9lDcjlxAKfu5BALUc3bOBQUg=
`protect END_PROTECTED
