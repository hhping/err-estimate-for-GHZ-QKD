`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WMy0zWCCB9pGcv1lyMQqyEXUW0b/gYZeQtaaF5bW/h8Vf81w39ybPQW5OPzuTSCC
9L71X6UH2Ue/wJ0lixgbnvfKKJ31FOQ1ujQbRbwy6j9eMBBx7/EgrIPGVy9TZ4qo
SDnxY+RIJsWDp2d9PmjKA/ZHURGY4Reg/Grl6dKy5v9NdpJZWgr0Z9e61NQaLICr
HFT62CWBvNeUR5tuXYXgi5VYEJueyidYQtbswlKSi7T74/b0RVqrny9m3LUlM/yN
E91oARGieUxdZEjnvzSPwy8+160RpFNG8L/Gb+XfWhwZl/BXYbkhZz3tn4Pstpt9
G7i5914KNSiM9Eyf2akKxSrRcyz7KNafFFY+4ID4rN0Zm4sOIguJ4FWdkfP9Ozkb
4Xu3Fm3QgZOPtH1AntOaPTswc+knfX5NwpG3Ir0I1ehmzi5yGEfcK7ojHQ848MDU
h1WE3VSzFe6dNnOopy3pv0JgaFnVhvmdWKKdBAfoeYvEKKUtajGox+xQGXio1UdA
YMUra1LjlQy21nn72VGPkNi0ooaXTfAC4Nc/HCmyAmjnjKHeNLnvHII5sdGKqTFN
kd7T1Nix3S8lQ7nmy0dG2Sah11oYAlxf9udL+1j8qSwMjhVDOYT3ci1GyNaszE6F
eFZcQKrvu6yER1nM589A6x0vxxdkqG68So0FTlPDOeCgdCfNtrF8megfuPNsFwWd
OmEPXrVxJanJrg56j52UAm1ea+dkwnzCjq7RMyQHQ/Xt6XQiwZgYqbeQS08gse2h
uuuy1IgJX0GNHWhIrx0xahyAUgc4fP9v2am8SoJ+eAYhmEFmZ8fHvHEHFGjywzXp
bP7Y8cTs1MwG2xnHKM9pkrQV3ZLLeoVpGAnJm6qY4kepnmc5o1+vX6BnwFk5/LJU
yKF6wJ7x+Z7+d4d4RRm+MWr21m1uvJtGINY5c89jW+q2a4AZr1TxDATHzedkXqv5
4QRcIqXN0fLJknLlh06xqM3oZ0H1MGr/mbunYwc4ISbp15M2UDsKrahIqWp0Lrst
qk3+ejRBqzlMybHLaJIa17/sWLQJNxO3tkh57yUBHMCIV7XRNVwV06GBazgukFH2
bO75t8kO9PeP9gPbfGVkAUuHKHOZOOtvOrQVLQum7v1fhd7sI2TCdVe7fFCYJQKx
re3fqVqxIB530lMmNqbGxPa+GOOaYDXMWvwFvwsry8cqrM8tuPNAVKO3R8Irfa+v
hTCh43Mk2BqiuPtV27wPO63bLfJIXmMdhllrzPwQBMYa/4J9k5+u4aTGVwKXdQWj
HiKVZQB+7TXbRUu5aGGXy3l6QXAVUyexhEpcrcP+d2SKZmxg80Sh0sdsQi2LQeEO
1773HJv3JwqLNsVJCp8W+XFu6Hc0+IzJrqoqa9JVNLqucgQik1/faDJ6VhqCd+6v
GguV2UoggSbcVeML63IOBi6+Ud8Gn0yyrawnKWX+1bEEr+gyZcvF4oacXtvHQEMU
yRUXdDJvGgjbRo5gy8EKQzcqKCF42PR0ONpzqZP3M/OhMDFt82JtGqin5dhilN/f
FnjhsPA5VKAEdDphZE1ueIWzftZ/Y/dCIh3fMWlAEKFTimbBXEhnsqkvY8pIKrjj
d3ryM59NfJ/BXwHV0j2d7Jngv7FsdlBhOCr6iZGA6NQuIhu9dHyZ9baDJbu+k/6N
nGmbNg7kmedoMKHtKxOT0+Ae4Nn22BlFzA6jg0elzqEcXPKi6y2g4azM0Auj8+t8
s2bH2KMv3YmNyUQOBRV8uTYTHrbImn0dxj5ofewSMHYZe4IPem9mMv+ZsZsHMKqW
om7tPkcig8wxh4WskZe2WG+mGI+J63cVehZ/6nLlhgM2JkOh14FvwNOwRVAZSAnm
sZpIoEHAQU/3LIGpn3PLNVPSGk947XO+50AF1lZ6oLUia1gssy9uJz8H0q0ttUoG
oEgodx1UR/ylzWxU7tsWKDaaD4gs+f5lcErkqc4VGdyy6IvxEpKJHhecqLJrdXYF
gY/nYvWLfo1qKAVPA5kI/dTrspRImVLJF9MSkdRgPnJmJu/EIQy6O/hCHIBJPLAn
PRPOIcCfWFLZB9hHGCwwVGI/a/4kQDZuZch3JMhzj8O1QOwBgv+y8YiKa8iaTqTc
C5Yvk2JASXLF1u+sCw2V+zEXh+tSk7nqaDb1Fz0WCi7cG2mnSyEyETT9r2EbHpZl
lRbgm6CKo4XtLxNZhko2oQ0wC13wQ1KJztgCgQSlN1vPy2E/VSrPpnQxIC37ivTY
MHymsXknY3X2RbXtKMdPU2itfA7PZU5RcAXLutLTIhwTm17HUrJQ27ik5cz2tee3
j/ffNmoIqJGoyZSKlIUyBrCyIA0DIqvljeURxZ/4Vm9XJmgW9xuY23WVFIzS5qww
BiYmpizRAy96MU695j/KNVtqmQ3JSCeEajKpQjG613WD1AraoKhznnYT2UllglVe
ASfVKdJO6U8VyvYsalU93I5OHU64XZpnxBsFY9F4YDl2IuAo64dcadKgH1xphkCt
n9E2fhrrmqcOid1yh3k9Oui2lKYv6DbJ3EUZw+Rj1OZKTlJDgp7t0jQh6MCNecZq
eXOat17R98zeKnPjCEVRfK0E82V90i+5nEy4WcgHG1SIfiaXUnSq5kHNH/S1EXjC
W1+Nx8I3nl3+2cC0uKWH8lDmLH47pPHtVwHCzT9I6YgYXNz3EHUXVfAQYISQSVRO
jmm+9424puzAQPZfIvvlfBWJ3DNUuyACR3p9DH3lsTRkJbKk8L26qXWltMG919pC
X2Nf1X8Iufn/DzWyBLmC0KpggnFgPat5mRbwXteSy7c2cJ6DEBA8YzKnt1byI/64
ei3DrcBzAicjU7pavbQ1trFomHBIaacoaC2uVIOu+2beorJwXChQq1189UlEet/m
uB5CrnjEJOZu7R6NKE/OH534KL8oDQSLArkKp3Kw1shZzCZSQRttOZw4cAZuxv4e
7QDMLdwOqcz1kSSswf1C7/cS1nf9mzgOFPwWVaQe1ap5LqMGN/M2XWqgu7lMkygZ
ycAglRDyQKOLEMYMTpP1M3dPKBBeso6oo+7n217wfp2lBrtmpik7eQeHj+w6F+js
K7zpo8wcGVw6MjReDO/dHs9N1RQ6/IJWGV2W4zvyBKWbEeJg39NxA4Q5iuHAtOhb
ywHR7SObewohYFzrxfB8/aUHJUF2BXslBCbuFODzdqZYfS+MgZWCFDD8IC/GrbWd
vW/kNaFZKET5P/8DRkkio49Q0vxSFiIPeKkUDSkS/XlP6cNc6XRgWSbZwGgVIKZ+
9zA/hAtUfFWqA2PsWe5EMyD8gl2nCK4xNhlfGjqfcSV8lNLjyJdSGwYBhau4xqGx
jaQSG8RznXTlHT0B6H/Pq3ae2TJAudVn3Zukw5tmDC6sLmyPDZ+9kfrsl+qkniw4
h8XVIU4D5gkBLkUdXBmV3BkbBaN+8MCuwKREFjZ1AjrQjZmBRcrBdb7LPMbkFof1
aGyQT+fN1EwWXL/9QvvO49FHOq+32ZlF4xLWU85zODzcEATVAOiXKV/SdW/U2FHM
ApP0Aq4E5elUL0Fl7mpQPhiREDeeUKfK0ApbFZk8jV0nulEiT3KPMqUQaDqJvGpL
JLQZkUN4HDbDzDY/bFpU4nirjLrr0nvTI1YcKLOK7t2bYU5nnPFdCl1ltCF2j/qF
Zam4T5Y1rOePd6Yx/kIY0E167dk1iWrS3mPG1Kygt0cKfMzcJAyZwzWkbWAFwyrJ
H0PYEOQ2e5MsP7RekzQoVz9atIOF11cwUEiO9duMZi4N97Nz+SLs7GDELYmhIvSB
A35i7FXb8zWAyqRANOxPxwlJyZD6a7uqOvQ4O/jbxwDPw9ufWuDmCMNQBeq//Yy5
C3W0wL+9Mt2tFFqG/KrxovrTBySbYRsr6bdd0pAvNkBpEnKRmml8/3BrY8ryJMEl
GgD5IV+XVLxSnedVtujvolJ07XTZrm1by5uI1CGIwtVmjvhJtzOZTcoMXrYCQSJJ
UcErcolkdkMUZEvMOpDUKs82/tNImY1gu0S0xYPL3nGGnV0apoWq7rzgVJlheGZV
R0XXX2fPRQa36LYhNN86JTL02Ry32ZajwTfTtuIgeFQnXLsLh2JugIhVNgS9jNgF
Ya+45EyRjunLrZXzBi/yGra1iJVY+c18vqmmPeDdclc5TKofxSM++fKPTtzSb9K3
lyLuubsg8Jpzpw84/CnipImiUOZaLXG/cMcnDa7d8tZz52K+i0m/MvFsehvIzemd
O+l8l3mJbkrIHZkj+wG1H8l1nuytuLcDw4E9u41TiD1lZFCKrYzsa0gARpm1UcCM
B+rPZwVaNsRmd+tLeoTEUDAU5PWcpMqMJtj1R9s2KSf6ziDRtmlbInhfURqdJIbb
CN92cec0A9+t3qhyJsJr17Uouip8nZCpkcoEXY68Wr0Cr8sY+Avd3SwZSCn+enMl
BGPe0NdCGaVuBqh4TGAu5E//Brn1UnHsZYSFdmz2esS1Ee/WxC0XWRPal+d+n2ZB
2mHy/lv0A01mmv4qkyBVDbhF/QQ2YdCRH2djU+Oh2s7W2oYwa1wadm4DXvqfmxK5
FI1pF8X28Qi3y6p6c3+l+EAphA6kDUSDUjuTXC7h6vz2J6jSA63LlyUfK6fEU7dX
kqKZI03aOMID6+xfUusR4ad5WiZ6qMnZDjEJIBYLGSG7Ds23GDkN4Ur5N1junCVT
PREXCFtVEME0wgQoBSczi5tQbx9OVtYemL0TCSltxGwFkigkJnhYCdVnAFI273Nl
ZTuQHXc9dK20Z1vsSMapFdH92SrGl9k692PmO3Mbr7K56h0PE89+zmlUuWsDIrgK
wGC9LE1SrIbT6t+Dcr+awu6vEKVpzyMfeGtBkjkJoKCx6usYIs15A7XSJ9Keu82G
0cUIblWRwH1VJMbjpvHNYbJnR9EOqO6SL6n6IBwQI0tYuXjjKSzWfHcFZa60izEw
+KT49100B1IvNZYS2cvKQrlKD+tgzfwOioMvmD2Uxl2ncXJn+AeVPnu+KBmimJi8
BdHwEPZQWgU/TGsAwszaqYivqImXfL1q1By9E97VqTfNLdtIlT5XlSxKBbfi44n0
YVWG9R319H1Jn/l3QCiSZvN5jouxwoz83d+PB++vhC+cg9K7m2qWaEE6eGYL7V/8
e0z+wwWkEhTQPJPeNIQyn2j0Li5zZ7Mo4bo76ZpNDuCe03qskWJkkOgrHR4pxIc+
KYFNCdM+9FcwvW23z/FDCbdegHAOX1CeG3L4xNcSp9M7xjQlAGu5gyOyXHIg4SLL
j+yoxZV9/ituxkCzXoRanXTBi4QjjYJqlOkImS+Kxsi6hcb9Ofi+6TwTdbKXNQZE
KFN/crFJcue6/zqaPV8Pja3F5ZVvXiIPBdat3MWSqzAlUSVTLQqq4ZQUocIxHwgf
iXTrW3YiAsqGdt5IacDvh3E+6ViBiwkjT5wR7qFghDGN8BhKO3eJQtPD9XcNgFpd
dZpadYdAeWGwbEH0U6pmtIKOU6jS8NfoYaUR+0XAknQ+akRuvQywVEOocpgDS47J
N/9x2CEEYKKzxKI0SeQlQSNlPb1ijXfe0drWglsRZL/uHz9XsSxGPc1ZbW34cwbw
tAAkyzGNfxV78CPk9fBYd2x1gmArzMU+qvzpr+VU8aJYB5910lINNCN0QCPDG7KH
OPNtf7v6voQSjsF/kLLWkeI3b2YgVXZWwLvubNJ/+HdQNdfzAnYzdE9ba6gVYvCm
IoEFYyhVNkvA447TtONzNCHdovukmG3eQvZ40bpkOMGGObPaDqfPILDK746hwL5t
2Rfgat1IerIsuIgYK20KGwiTJjsnRAW0p8pMSZdqWMudCPxpJ3I+ef7jsePcUHeb
3a6cHSR3W+9Qftqxgd7wcvKi2aUr42zwghhfaQICDuEizcwM6q2+2/vUUjgGQY+n
o5XeIOstsEIznDzV8BCdvuDPylJdukfF5GWnTmQAjD0I7p99HhwS1V302XVVU81g
d4wxNq+zVlnN4vMJ9uYjfwORO9GFiQ6IvfGV5JTaT0v9gUZihf4cnlWxrbdojUbA
7otarwQ0PMhDvIo1vFetelxpysqBnHSMEfZGxwNMwGn9CJfiIwrUXs3nL2QFQZxU
pvt4ipH92qh6FkvpC2J0n9pqH7TihhKnFYxm7Ug2U5oiHlrC6bW+5/1xas/PZpVm
WSbv/PhJHUuljZWFRhtQtq8islYD1oXkInF4p3kSZinXUClPwrB2ayZ/QkTV0DUU
5rNXXwB0Rc9YFAG5BzxzwzZLwt2zCfIxm4kZXypnVEDMLkuys7RjidiuVddTNPaP
V3auoBuNi+F9w8S/BzM/VOLZRp8E9rnYkHSwEtDNAR1EOQqPBjPB0oDtMqWHcXxV
p4DLxvof0M0S0X9FFfVcpgrZVNm3yOiWlFmnIS3u05UAlKkIiUTT8e6nhLvUqLYx
J4KpfkZmku6Gt9BOLkptzufmMIU4uL83+F9MeRErgQygehVIhOSvcuDDmm220YwB
bNHUCYTGLIYCpDYBkasrNedwCkNhEVCvZAPaMkYJmCa6Y0jEN+NVts3wNVh+gsGQ
hah7aD0etNhXHharpcEilY6GamwJfFACxhhata99B1eE1LVnH1JMmzfy/ERyUlkq
5NUkoucResrhObkkxB8yHacAr48HllSmmIZaV2JtMFe7BPcmgFflot4UIoWAl4ep
QZQjWBw86bG0wJ56HltV879rm8NHQcDEEJHLyiNnJZPd6xKvVbvOGuX3XsSnVNsN
jkFwg0w8qpTnIiVwUTKN22zluPBvCkgN5DTKRqaR1XQjA6zztsOPjjkT8h/jbz3w
Xw6/h+oENzs3RoUJDLfgiuvgYtuYV4Kqk8N6lF8szqpNbU3w31Ft2X6FaVrk8QBv
7zRicd22HmkIWLUTGLCBy4sUfQW6843fU9Ig0AiU/RkCVDqwHsKAqyB0YUnU0Och
P82pXxmaAqRT0u0JqQSBCwUaOQI+pCjah4D4/gEOmX17qtiZy7sKxVP1+gNEXNAW
ee8pSA25bJAGR2596W6g87pikOMhDYJ7JDAJBzuwtRu5OmqFJAp1duNfugcTZJkQ
Doc7qR8CoupOOPVKNDjhBXUKLhmqxmX4v9FxaY07wRDmqzDF4jy7hNX9eQwoU2KC
IZ5iRwhhJK21WC9h614VlWWyPmLwLZ0wpv+1RxMoCz+gQkfCc6or5jglk2x6RJsu
Y5pfDWSGn1ECy8RQoTWyDG9oPlEiefj/Zl4AgS9eXumyof0RCYUiua/R7HdpkAfL
MVeBHxanqcmu3/3N04sOWUFZUBra3T3Ghh1ECJkcLBjaBMdX8X3Fy0PPpMAgG5Es
kAjKXvj535W7cyiSgef2oEQFOekfr8v8lCtvq2nWnZTWOMuX8nLsxvTnXmFNS8+5
E8USdou3+Bq6cK8XNfNzc7ctAfDCflWFQXEKDEQ/Rvf0zepZyX66LExlfcmsM5Tb
iBKKlNvz20J0PoLyEPn73v1bQ4MjAeV57wrUNS9pnME2Qn47js1j29tCwgcaiPeF
NWQIM9W2++7ZZf5eBB72yB3XbF3arXWQYF3K7dBFWhGhkhfP/qZCASEW3dtNb6Ui
+ciZPlLmbEzYGB5ShPWdaPPmJPWBmfsydx3o5FTofUTUbaXiixHz3LHUVOcP+HFf
r3DP2PqnqFFHdMyUkSVGEa5mv/CTccQsVyiD/AIDjFlXkajBL5GJVqXWkYYhSCxs
FStVuMx8tKB2SddMgkycSXyMV3mVZ3FVcdXBFP/uDZfTfB2Q9KUouulo+U1wpk4y
jnQdObT3S3uytXZS/9dpjPZNsLdPaazLt7ZM6Ro4ixf7IBDnp+8sZqsRVw8cmdPL
0I+TFZfTZMLD+zKAE2kmGBNKGvzH8lgIDbQ8FgPZEqmIh76NmMabNHDKI+jz8n21
YVmpXWMjVVi2j0Xs7bsVKmRjQabnlq9LsRJ/tjuim6RgqIF+1HA6zP3kcN1TqWf7
HIoeAaEGlafRcZnjXYJYp6aTG3b3T5sxbAd7DwZX2BvblgQGdpBGZxeGy6nnuXs+
zbkfNNtyo5odB4DGBjp6095ONagAJ9k/wZCy4hLpW2hku65MFg0NfD3soD/lQ2/5
tzDROGjbRkHjdDSP4DKjJA6VZMgydIQMtn0F1lQV4tgqSvd0Vdg8ra2xX407s8un
7Z/eY6ZU8oRDvkF6jkh1yovIKvtIDVA0PX149PO5X6fK+cdFxBY8FAFEtyVl8S6s
l+n0yoRQQbkaGw6nK+A23OGHhVSjXlOcr/5s8/hCIJHMD+gQ0MtQnIJGUVIK0IpI
HF9QEnjzPutUrJzABVEygT5Up8e9iD3TF7k9tzQrnv4tsntWIcOWsJl4BV6+txh5
bfjJqX/ZnVqF6RiF9W2md0ddAFMMt2MCy7vamhIVFzDjn32NVmkn52mLGEmRpN+9
wsvZuDbxEOUTtw1YsB1JfPZgRf35LrVOJ961MSlS0WgfUFdlli+h+bFX9fgm1LA8
IemoOmLplmOr5WzkF0Fhxf4Y2fpRd8nPEdaNQNzzXbCQ7b+ng/hdA7kknqWysa3f
khMrp1rxXjP8L5jmaIRrewhBwaaVwhDiKQIIQCMZcCfnds0Az+7EeHm8gTfItsU8
Bd8wkIDKcSrpAgPLKm/FbjoX1IE3m+QDn5HSRFTIlOXgjT4lgU0NGxXToQIrd3Bw
J3izLn9ewkvUEa4HZiizjQVrYux9INSRpvNvmumRjJcfuaawqW81/8MITx7kNUO9
cIAge+ZWSq22AxRNwO4+oEoMcYePuaBmqrRDCF1KRIdzylpaJXnXSGNBopBZo9kT
wsUF+ot3qUsfH5JmRnI++DWysVQAuBnCNr7Yc4BNMsWwoHFER4uAsyJAcT2sOQQ5
qXNUzCOEgHLSGkfHA9pQ+GJ/yxRcL1zPKOYp/12L4xxufhwSqSJ9NCPT5D8FJw5M
iriqKJnEt9dRl0SRqfHBEaaB3w7V0qHUSq8a+aSLu9P8tYqCmo03RqSto85G9AdJ
HkiSNbzS1QX3qLTL94OP5wkHzWXBoZpCCgthfByC4jOW2vGVBVxeUiUll90SefoG
92yy+7S+hVxVdI5fHMPZog/567kQSWfYKQWkPAqmY5w77HpObxZFtN6niiXP3wcw
olqgcEyQUZ9deGp4gKnm++50r2qujNfrfS9xHUQniY8vMEbShEqmyYlV0NMnUbj2
gT1316LlyN7J5qM5XaHVf96XUFaJszZGRCSuSEzoWVjKZ/THNvm9l9n19zKVebZw
lvDj5PFz6u/vrmzcm1b+fJp0VKHyad39O3EI4BA0Gt8EBP7FoLqZu9XvlA3S9sIN
csVMKG4K3dR7B4P/k+NwwQ3rdLU2ZNs5MFvihsjFJf7+EkZFq5ml8u1HxPpclHfq
VCl/P8IjN1c+LwdGq36hFv5mpXyWABXvAJ+Zm4QScu7vra6tuAwa3XppDCbONMSU
UmP/bTCQCMzagWR0oZOpWQ1jcvVsuuy5SdS08BW+nYAPQXfxHw/sfTMETBE7MxmX
wglzrJIPfrZUFyzvfAaHsh1yq6aEq6SIaHRM2GzoPuyO1CNkT49rz3cPHlnL8T74
i9ApknCSBMYQoZ6H2bV++qbXr3wGGHND2nLwpyXGFBs1XCypQKaKf/ZaQYWCpCBS
u2KBTQ2qW2xic/+BUHDjGxWLs6vqrVonzksWeAXABU6qYK7d2vYcBW7ODiWeqYe6
T4Cu8p1IFXBc81mQ8WCPXGrAa3jgcdn4nBzk+k9yp24GqT63rzcvZ98Jz73FjoWI
DjbvQS4cZSzVVdDli4+W1IhErOR6uN7bkcBpRbGOMcoT9ntFctHu49uiqwTs+K5Q
D9cGL6AP9ya4JKaPuRywzBOk/vH9UROPafteA9RicBLNFgs5C4nHRDKhAzXmvM7k
3oXhrD8nABnOgO4rFC+POysLHgvvtxwQJANQCJ7D8/xZGIMDS0p0esBPf5mLbcl3
iQIjBqate2yvzhPd7xfyf8bY22HLjmtxvvm8p8fvvzq7IyLFM2yRJVkhTNM0rtlb
8xIJi9d7x4Q/1PjQgaPAPOLIrg697UmV0R3KD9dl9yWtHGrjQ0DQCnAgKifebSIc
sqsWjhlrKd0zx2n/iJm590EZkdgTShmR7O3/b/EhVreFaxcF1meESXRP/QYRk+bS
k6ioKuCXd+Heu3YKs3I8s2+kf1YFyGzLQZlFgHduKorrsnNprcehHh6mvdnNlWDd
Sk8f+kC65o9W3LvZPsF+Q4Kkrmr4cFw8/DEwz4ZLd7UqJcGW0WF6Y9Zm7uFJSu8h
IP3EhUaBXNC0CpqmnU42Kc9/uqIf3bKqioMhEWirQzlqkXsvaFaSvlcNVQlJyKnc
MtxpXMta4yr9e/MfntOZd2P5fULf0X/0zJsYl2/1HcH52+oX9kiFUyURgIi1rkdz
POCEAVRxT9qMVGY6jfTHOK+POb7IqtySMLhJrkHmUwlCZej+YWaGLeEb9L14fm9Y
+9CxiD/DwBiYiH1J6ptm4suiSxj6tf6YC9GMibDAr2kzV9Sc4yTn//RJdwTuZD3r
EHrvelG6+iVXjf+10a12aMibAMnaGzVsZFp7P1NyyyThwtqbhCNkSztSQzv+Vu/Y
CtEAiWVAGj3aUCAu2+k969XO38nea26/MUAs+yjV54SPxeBYxBn622uFApKHdEys
D/EKq42CH+MTqjncEP2peE3JcQRSQNyv5HImD65bKWoVN2OJFo3NQi3gKZnIGhQP
oKkNVNVv06HqgrtRQbUgA85A0MYHxt7lvO0cmMgG1gvj/huv4BBP2mzF5wfgdNof
PuPdQxo2W8kGaxxATfElork0i9FP8TavltDepxq/jTdpK9ZnQnRgWdQIphXEaDJ9
gNm3gkCjHVIB2e6JGpqr4sfg7SiL90emkUZAkYkL8DpirqO3IzDpKyindz21jTUN
Jm75qped1fQEDhRXJN8hXoCLZZ9gZGBKoem1gjhrxfBN3UyztfxoFxW2dZIxC2v1
ocMr2mVfFoL+3BKiA7luFJuxx2uyyBvWiWpGpL8mQU3zWLcJQGbRkcKwec95loOL
/eBU+JFedapwEm7Igb2RC68Ujd2SpPt96L3DC20v0TIrc4KWUScIrSkrH8jOz7Wh
zanWAf0KULpC6jhb4usmgIgGDdKEFxHUb7kSu9bd6L6B+fX0eyA0WG5MnVBlGOVM
ssGwSErFknORA5ThhbdFPXn2pB5aFnCYDXNLN65LgxjnqfN3o1MNHXod/sFuF5QM
XAe1nkiHYc/hRj8YF2gKDwKL+QfviDcghs5t986c7TArl8m1TDUu6B1w4v94KOPg
RxPsYk7SJZwVkbKU/u+Zw9k1+TFUz1+bNwLD6umPv3CvE9rAK1wjd/ENmM8sg9bS
kk0OiD1V0j6b5+8RdSqIzW56sVyrvW/dgloMzoQUZBQ7wPPUj0BsOdc9nBioWeu+
xMbBGqt6KqqmGIlOevCwe7buYogTVxjsxu+C66C3sDhm/ZLkklJ3WSQzJ0Dff55F
dfS/Yru04MYj5PBrP/L4smzJgNc9bhq7xtVRjme9ige5vz4r8dBpmQlmzBr0z0xC
BSU7+/oB7aQHVSBsE6lHfu+SHpT2c0J7gxKhCM9gP3PP2VAejSA5PUus4rz4qeCr
HdkBgeKF+wgt3snDkO8KSmI+Sk0/q7aEKdu6be121h2yYQ2i6NNpDkjU+XKjJb5m
a3IBl0WXwka3hNRAlx8/PpTxhaq8sME+atEDQF0tsac4Lk867mhIRK0oGxTxcwzh
0wPiygEjTZkzJX7FD/G+SZ22laFj9mVIfmF8io8qbNw+pRbu3DyYFLCXVtVcCIFM
4h92VA4ocajiX5kdxlAoMGC12l/eUrK5vkitWoPu1grlQwg5CWa9VEhxWPp1Bouu
g1zd1OmDD0PNsOBCcy5e9uiYXLoA9sKX+wTuR+8/8soYtKbFAKUFXVY0pOBZFc+2
JK8Xno1sbKvLIlgN7JJAVMHwsI7/58Hb1+DZCqoA44j7Kuk1wWVqRgAuYVhdMaik
rWePuxqRrBFnYDGwOUqnNBFou0DjL+PGCM+cZpHnlfC9yuXXIGZ9JqQBDi7CeeJf
w3mgi8ShQRhIVz7Fw+BbBqZufbzBPX5rSYsXaxRoZpGrWG/gzeb1dMdybVS8lXkE
2AIaCsx1B6foJM87ABH2gnNFiI4WGd49h8Sd9dCES5LLA93hwi/piWeVjoFG+PeC
/+WKp2wzmtU4M7QGeA6OGoivkMr2wFRkomFNDMaZBG4Jz13CZIdBTO0jdNm2GJnv
Sp46CSrxo8AkrCH4V7G1kccl8TF/QaoWk8B2XE4KXq73jZxEtm7YDYoTkkJ1oh94
yhSnTRq3bfqVH4sse0wz/+TjZAeLiGhQNToAOzvlpkhUudmAfqu/A79oWIBPinhI
MExGgSgoyjdbKa0HPB9UUi+JZK1wKppl9eX8SBptptNtHGDj4NPJW0fNJjRsvCP1
eBw8YhDizgM0y2XOGlngZDJ4afuOEgX2FkBxiCJPwKFLBhR4giD8ibaTqoxFE1Na
84OawhKo2dpq081Fs+OzM3lN+D9ZLVy9GkhgQGRu6+ZQE4d86Wn0tXMQWhOGP7dm
j3UnXyCgBCyrNMTSWOjdqU3EUP1ntq3YPPlbaTUeWyx2VEygECcJeAlZwsAxki14
tV4SBLmQt0z4H+xvxEZtd845Y7amV6H0P5pLsm2zM3mQr/1fUc1NaoYipY2c1vq2
yJLdPB+P0imDxE9lFlnD3U9UhdMDe1IB4TmmRtShJkaoPVKdjFU9eD/uxzdizx9N
bjbVjkcQU2evPDsD8yx9HDvZGckZXqubpRuzxLyApublC/3BrLBOJLH7M94PWoSW
ZUaHSMYCDBfwazDiNRLrOq0S2uYU22fXxMrBbdG8NRuzJoQKp/HY982+aGcG8+po
UHfQrKvbGcUgY0pFq3KdrcIL06zlyoOJgQotDm8zKGSV8KkHPUFv9QpLjrQN7ibB
9ktqgnADmWeiT+KgAH3Q47zqPNN4X+3dwTAEkaM9xV2t4aDe0ZGT6qtrWIYgK/44
v811Sb7fEfAJsodlHQ3M+JA0ep7M28f25Z+U2Dk9JQ4YbIZI2j5G1r9AccNo2nxO
yQlxia7GK2n9nj6Hq+mZTm5/tOk6UDUw5m1ngp2U5SNzoLVeAJZ6LgCuYQjqy/1o
oh3S4ya65jLde7kfgbquN4kcaLMWZBNDuyjLiOBa8jP5BVDX7Np08jx3uBgzFqDD
H+Yv7in0A+Hwm3cVcVBmB+o8jdwiclral7qf/OduOHQsaxz9Hq0rN4A+P9bcL0Rs
z2hfURbBV/hSTpE6erwpOeaJVWJvPaK+pOwzW6cLpFMHmDfZ7R9Io5DsjJzSoKqA
p5f2by5zD/uGpFa4SFtAYLKrGFOOXr8XZ0ZSaioai4S3DHvW3xGHVnzqeDButimN
NUnOJSpJjzqNIqiUVbp0HrLJpe9Trpc886FpNjHlyY7v2Ur7zV8Va8pFXlksb4vg
MlHFAFTOv7CN60d35Q20AS0noGtcO2tdMqLAykTDc/yvcjWRNt68KRM+pZHcJoRK
Fq5fyr3wRe+e2cNj9tfo0mtJDMgqLerHo4QbY+7fU8SwtmaRFfowHOsuXZYEFpUN
IgNtOcHi9yS9jiSgCk6SvljL5OVr4oeEIMgRZMe1C2cJl5HR3f/Bmuku84LFlLe+
j1iUrsSD7N0SscpijmuVxal+WAZ12B3eilLc34m92k4Y24j7iZ7Sl+YP96bsbEL/
NPQlhxBuAErfE1lSjmnc3ltcvjgUqI3LKa+s/MufZn3vAji+5GmjfrIO1YIiQLun
+HKBDlsEAf6WHd7DoyuWJGFfQrnRuhLa8dTmoYBmIK8Gaz/Y2XZ67Z4W9prwip+0
`protect END_PROTECTED
