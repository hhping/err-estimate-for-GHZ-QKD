`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
72AYnR2/qYQymjOdebZG+3HlhmWM7hYVHThtF3X5pI/bTKuvTzlt7f5ApmELkYLj
U+zPoKhkePUFZgXJSgtoIDq0495VTtlmSgBGcDUfkK2I+Tqu0qp/wAWRUQRr/4Aw
O/6ihtIIakaRiYg6osiPy+cO8+HoZXXTo7GhiyGGh6lZVfyFZfUejIv/OvchxDDT
i7P/epula5U0yb4/buMi0PdhNNARffV6gfGriW1Ul7V7BgRC3j7AHWo5ERcJkagj
YYHT9gduW2Ud3Mt3xroI8lzZYy/5/mBAtMA81EhA3FOYuw+wh+6O4GRO9tMz+jFQ
g6HrKxl0rbzBU4IYWs9L2RNCJe8SVgiviUXPN+MxpToyPXNGqgpxTbxeVn1FDjAK
u73bwTbl6BBJA3sBFGX212tpv0P2eRVsRhQ0Yjib0nfpIVz9Ub8EbKy7W0y5+Aec
p4/lD9nKE55jBdb0hAXXDwWdXCOEO0GjhX6jOviCaUO0Idge/rcbfe5705qQwCdm
OIqy+w1ZYBtk0FT7hqJUI2vDpmDMWl55kCO1teFDRR4XCJXy6x8Pz/5lThhsnNO2
xI37jfdzd8qORi4Z93WvyBatNqi6k/CTK4ceykdcvi+n+vXhcmgtPu9ooGdXqfPI
453u6LI40wdYkEZTGZ/w+5vgmR+5rJeD0JgjMJfWY1HvraBSMmAkx2CRmXIZKEXR
OvCONC3h7vnwvy1xGUuZ87Sg1bI91E/5y0cktm2uaZgtMlN3CexEycGX8yPCd0aO
D55gN8CbWGhVM9LDLV1urI8k1kzBfCmPpQqh5MvF2Qr2Nh/tzuXCVwM3XZx5Y5Xy
iVGzY+VkdIly4gcuIHekWg==
`protect END_PROTECTED
