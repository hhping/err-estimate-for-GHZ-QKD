`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rpq+4bmlfD20LYqtKc1knyLMBbQ55A6Tr741CmOYPS4fOtrSHW5/5TLLMri2+8OW
bUAWDsE+8bE6qqSOySUwjaUWnTSGZn14xdKyN7y3MM01QTzVhM1z8D0ktqIyJ26O
ZAL/HDrni0s6oSI3vHIDZjHWQT1RVduzAgSA0dHs00RuhqKbGosEW58zL+bt2m3E
M5Zl5xFu5SQnmGDLXzT72rBohJSz1vER5gQzkutOWQgy3utW7C+y1DPSD7Iq4mw6
o92H7O8a35+WRsPuWXvMg60rK6RGXeHW/v30eZNAON2GMK/W+RiQDTUT2dvkjr8V
y3uEwTkMddLKdoetaGn9Go03Gd/+Ibf04WaIY+3NFreDxeNjDqLg1LZ+3YlTmcqF
HrzoG0iRFlsNFd75VqcIsTdlZvzaGHE+bfmovxj5EsnZvHQh0XFM6Md1rE0hamRG
Pz87tEDKvmVg0re8himHa/qpYBD3nrdWmJrSME/4As8CWKe82qAMo3n1O9POTMOF
D0ZZAniL0bQv6hmegZIw6yc+oPTGjRgoFSvrGItlpFhJDrMsizMddaN0SPhcG2c1
HXc86SzwPaQvtEzRyeW+4dOw8yMVvgiUh7Mg49okLWgE/4js+FtxBepoZ+a/lLgM
2turAWUQsnZoYMCPxyQF+znYGpeI9ACV47ajrHSs7YaFfP+IoD8/BcXvU8fNWHUP
58fHSREKRa+aeBv5MWsaA6w3GdkLsEWYz2ZpqwfSgJPC6+NfZ7tQE6Y8fn9f3MNK
fmZvLnit55yiepcMwrVmUxFhwJwvDKO3gXE736eQSZwfTvLh3wsF9yvdqhOd72gs
`protect END_PROTECTED
