`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rB3prNrOZlPg9bFm6tZjBAxFdQKSP7k9T3RcfXnLWNfboK6nZ4pnAIVhQO6ied/w
CVIOvMn2nxDW0tIwtgDkJrJj5dEA4M0cgtOy5SIqKCaGjMcg9wA3J2gr5TobsW7H
TV2VJG2zw6OByAB1WP7WAH0c00Sd21OCSZzsOPUFFXXWqb00JcLOOWyx/WByunNb
96GmuIo8oa7SAye4QFAn/CzJoa/vx9xLt56gNKEREIg5I6iIKjvhWKIqShqaBIkF
KzRW8eUlxFEJ6OK5wukMQML9pO72pCZ1yunAa6pgrBfGJ3LEIKv29lMXS1zplOVA
hiZASTg+yYD8/p4UYsRFBnLlofLheemRay2SyYB47cQVFTlfqGv9jYSULmiXnlIL
WMjI2ojrtLrk8R5zYbrnNg==
`protect END_PROTECTED
