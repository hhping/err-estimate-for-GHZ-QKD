`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/aZ7Vjm1OEZxkRC3GcTby6aZPd7+aX1d0sq2S+Kd/g3Rt9Wssdl+Z4Iya/avqkWc
gloPa0K3O2enQpm7R/CLigphivHH0N7PAcjMo5dDP4QdtcLhnmKgVdm8aS7HetiW
r/L4XlI9l1tkrmnflC6FDZTb0JLDqRwxWDO1xEtjed/7KDYuint3q8ho/pMv5lQe
JWJfoq9yhDQoeA0vxYL68pDTF2Mz4VGBEMIXYWOav/Hz1AEs2mwQHeyoGMgCyTSf
d0LcsjoRX+XwhTOh1zFqEPcfeeW2b4efaqwZncR9Fd5jfuuUtSpqxkIPj/zRNokA
Er/GVoN9AEWM6QaUqAscN4gBoN2Fu8QXSqxa3sNwYEW6p90G4ep8M9xNerIRNo81
eOYtLTZa8rA1szQ25C061I/4TYObEOOptrjE8yNPLDwyjDB+x99F86YMVhdmNaD2
eWVSIe+BMb1/dHkTQ4nW0sTR2uPW5VkvuMqMX1hHVYBr/enmaTA7ZZkR0RITXQuf
qWOmGtI9eFcqSLlS5dmtXB3C20cB83yTzsMienW7ZmcDt3rkzvpK6xXVmc5hNkJs
auFuNYNTYIimqF4In4munk6dxbF8wcOHDVKyUVlhviaxVYEYulwNMMo+EBEkmGTU
hJZtdzomgTt4zmzanlf7/1048fK/4EB/fsLIvoBqL/eM9KvFBaQZtLo3KQCaGuud
6zgTRNAr56fEAaCviBZ/akoKS5XdjBalJS41Ij1KOQiDG88+Rn8w0u8LB9ASlKwo
z8F/iBp/V2iqRjPh9xe0kwywm7mpY8UaoEZRStoZpbzlPhvNoVEy4EiKP9y4snKC
OqyxVFF/dlUDPfTOaTtkRbM/rVxIAV0UbKQkbPFkV5GyrSmmicDPVIq/snfeHJVp
xIbHBiJj0xGf0JH/CHoduNr8LoubY8ZbmISYqoqNpFhcs3ajLU/ZqoeStphLvWFN
fWCVR3N2wi098v+l/tOzzg==
`protect END_PROTECTED
