`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aOF/RrbqtzUnrY5anxWIvRrLsstlA/npg+/GQC5AH4tRWfFNu2p8Kh/tAVfYIBKa
cjMeZ9RI4EQ8pbhEmiNjY9csdGXIPHqITUfWKm4P3lo4ssrklyv9EgYGvhP5JYlu
5/j47FFPTyXUcn1xB84hOlE1G64s8sUYuCwA+M/Y2NaFSP9xbMdXUMlN+cKgxKEs
/wqhB/ReatUEL64zh+dXZR0GzKob8qzHloOlswzIukNTgenFU/Pbolr0q/s2w3Q/
+0x9joxXPc3BmpCk1MldW35sKpqLrMzkMkiA8WWUZ4QAAOvv5Z89v73+/UX3eR5Z
C8nt9rsPXOVYrpzhOZX74+ubeVImEwuIp8t64EPEmnabOk6tjgXxOD5B3fzmQe9E
wAIZrfic3DQIE9jIwl6SKcdxFsQS8WH1uGRyWDvmUg4385zd4pscZHyqdzuTKm1a
yPUh+mtJ2zLklNpGN2osH28hg9A6fQCoMv+0x+GHqnrUq/rwklP7FL8HCN3HFSFO
xcc6yDpff0eIASESSxq3Dp6qbiwivKsglQ5bzDGjO2wfGLAuzeQrwdNNwbULDMpm
kzZyyxFkVr37mJpF2sE+vhBMnuij3fOlKB1LYcrDlc9KfXwbpJyMy+pXM/bjZbA9
HBS/oqBkEvrh8yxMTcVs43wtkQpHzWIAzeMKWtpaZZ1Ou5r+/xUJ5KFBZiFbCfeN
/qaH7cZvMbX1VFlUrPK8B1O3smgpm6Nrcpqaa7mzPzMOZp+mK1SHjJbEqdKhl0k2
p4hgESmhEFVV32ba19UJAGfob8yHBDI5PRuDIcs9M0zHFtFml3BNZPR4/ZnP4yvx
ylhzwXQyQuq2P8CJFYGcgFsiyA6+qDTOqU5ro9n1o9RSoO+H+cFInvuxPuEulzWt
ApejFGlb8faE1zFq9++b2gP1t348uryh4/RXqDxH30KnkH5EyhdZq9n6/+lLhwX8
xmaHE94XcDIexEyFB2IzloEdV6VIV5FM3NefS6jcQ2cXKPWIpyHi5QL1W7aHKOeO
NtCkThO/2WULDd/RFSR+yD4WbxUotghTgcUMRmR+w109f7cj1ENXWA0z9byKD1Dg
GG9xU+HpqijTsnAFY5CtYeLNN60TzoorMzKNX0CeI+Ecev8VccxPsnD9h1nNIvsI
7XfYz1FxhOiBA947NBPMZNVSCSW/rw/pfshpHLXO7NDFG0G8RhnGsCaC7BzSWZzQ
C28jGYiB0YZ5kbQkYlHEu0wDUFl/zzvs0H3txdRscNsBMju7FBEAsU8CjfOFci5W
UVskH4Q0fDXVRteeXl4LfyPmsoJksCINNh7e1oCt3wLg8AczOGO3qxmQynLyKD1T
4z0wrHoUlsic1ZIYM5nbS4Vz0zlR6LHXC8VO4DJImwMe26T8vEuapmmGeYxhmHTd
y1ciJQLsRAW7N1gXBdFJJlTWx3y+LgPFuT8OxmZFzdw2MsNTls8ep0CEj1aLbXwj
ZUkP0dsirCvQAKxE7a0yobefdEzcRy61aYokWNNhE5LJe2itwmxMTawH7PmITGaQ
OqL6/XRGi6HNXLsfnpCTsghff3HBHkafvrpEqa4JLNV3daC8fbFsfZnj4PMZ97OX
e5+bsYKLeKg66rT3mrLiZvEqNtiu1xBOpLo2LNLPNnJZV/zB5uK8K9enYQ9rOuTz
KssFHcor4fWa6IZstLJvUuYDfzxex80eG8P/QlFglps2yPb+Uw7IY+bfHDH14oq1
JXSzEjSuznuqTn6aqHaDkuyWbClTtlFr/paUB2vyfzDkN7psnsIIn3Gy7Yo0Qa34
ENSBcyose/Iqf0q12SpznOhRQizxdThhB9bcbGwGYce7CxIDfO4IDSEj8HUSFgpU
+GK28EhECDzRAf6vi7DjwlbzWq8plfN5JKwrEmo0urD10yBnCq8HxVWJMR8w34Nd
B2Kc+8n635St2O2qtBjrzsLyfqxvcYIBp90Q18UhEjvooh4ril1zaVzI6KI1NLwG
eB1k863XF8FpvsNGH9hBIHTqm9heq9Mdm/4FBn8QryCUT1mow8YH8IJYwQFugz/I
zvBaw/5IIg3wLic/GCTuudfsFPlrjp0u6pWjwm+H0v7S6QSVZt3XW1sz7CQ4y1El
csCPdtZ2cuknRN4KH2KcMfJCnZ6xUQmg+KrcnPY4J6vJ638JTk3UGKO/sl5cKryH
a6N2QZCr97LfXZMHmA8htn9UMkm0jxh7JR08i2SHX+7sah2xrz5Ex7qE2b1BI8XN
7ZKPKikpnvxw1El5K1UzMxVsctL4Q/g6B9seelsluVb+K6vozjtaPwjmSF+ZHNAi
f619BlvtavwZnYMvD+jwbwvJLc/9v3nvfMSIzhv0WC60a2thDyqlaNM/QR+TOLu0
yUSQexb3lonbyQ3/WQeiOCtwiYq6HqTcfqW4ON3TaA9GOhtdQ6SGBuxOP75kRnWL
q0CmRkPowmmr/tNwvUpOqcLASaoZfSDuJuuQbcxGAyD4tpSKVguKqPcZe21kQe4r
cCi8JH9UrldyoCZrHOnjIyK3DRGj1Pn+ZNjgE5ySA/XElbyS0nff9oPAL94AFqgO
Fwdbgx/69Oiy+81L58hLDh/Q5OZbt6EHOKfO75qJ/EVGNXzk4YWtuFVZoaSE7URo
VaLyuBrWfpawxmjVbIjBSeJ4tb77c7CVXAxDaM0KYK93h1O4/K3aYz2mlOP75Pvy
gpovAp8HbXbyzp90nzWGslU5I1Tzt8pgoFFyjRi/knpka9qpoxoTllSBG7k1+Hyf
VgJ2hQBz7XcfUmL/og//CEoUjzbw5ElwiXmwgoAaZIdSxNx2NI03jXQTR58R8tdx
Ml4m33bnK3Uas3A0v1QINlGAVUGzvtZ/ESul7n44HuSMseFGHYQxGDBsC0Xt0hIm
ulj94eNhK0fQHq4HS1xJxfonTsWGoQCZiJDEzwRz8ok4w941h7HirQcW4JiZPOf7
B/HFbAtvoG37ARsxBAqM9x3FD3AzL2RnZRnDQ0MA72rp49K0eVtpfuf3uUrtMW3z
mv9rG8stuME+LBV/dIA/JjeYwivY9lpto2I3T/gmf9Is+YWXf/RMtSm3yheVrFfc
za4uV4iDBK9vUlYQqL94XgtkvH8ilNBNc3GNgOW466rwlyQrWmcXzRwjTu6Dzju6
V799h5fRO8MJ1GZrwInMuuxZhuiziFZfYM9LNjP9lD0Pjszz5myMeSDwWFgXHA/E
2SWfj5JAEfi25Aux1gCFpZilDuj512NigzBz7bHLKgenuZ8bq5RH7ssNDFNVpIS0
iWL/eZ6q0kfohv+gStB5iLh8lmG6EjAY4VApsDez4BKBMt9SdIBJ0IfbJ8x0JTLy
+R/MPjHYpmovwTw/TxwhvM1SnQ4yqRI/uKlmIZqFacWZKQgz3TtsC6Uhyqpi3bV2
TqzDv0zD1o1Dr8RJFvFOFX41VCT90ateZder8EpYVuf54YZHuT82XQTTTsgIrwt2
W6hZmzF+3aE+g8KSOaj8JVl80T7pU0hyF+bEVLcKS+31eIOJQIFairxmtgo2jKbp
tcFpchiDTWBetYL9WiKrwIBO2ccfguTcX9nmF/XZXx5phQVYHnGrmABoyYHE/BJR
dX8LGnVKPLyVMDQn5znJMx0jzyJFYKONTS0rDCzgV9cVDSX28X9t6g+gD7JKYU0p
Mi4Asdcq5AOD7i1cI5JiAyTC/weKra0De0BvjN5Pd8/zRLInJ0guDMHzcyMi9TJM
fBYT5LrtclRQFDuVJB5L5VQRht4gBMVNgCScWMtloA4KSHYwoVuyuA7aCJyhsS0u
AUGxGKauJj73ktlFkolgwizcC9bmtxCzr+WKy5WI+ucq+4N7qzFsRkDrSgLGYmU9
dxlWhB/lVO0+oNnWmVUn2s3gNN3XeQFdOyw1FJzdRj+qIZSFd1uqHt+eWWl5D7jj
BeqNrlPcj77WJW+2lUvYuyfAPX0Yl7F70p96nbNEXR2quPRemhfxJB60tz73VYPE
O3gSIW2ELQl4ueB5m/QNoNMMZ6XrSxITGnbXZ4qESsmYMw7AC9HWT+OUInBTssx7
IaIEn3m5A2GqXYmTccKbY+hyUd5a+4TrnmR9R3Nq7bo8O2/wPCtjsf3P13nu6fa/
pM7nt1SUWfTt/SYQq2a/TYiLW2pYbHk128AL989/EaHYCw+QYGiqNqnw9vpxbMGe
9djeI6IL3RCcsbrx7Ms5MiDME2NrT4lfq8zmYnS1LK33557O8b/qjUJmByRDv6yc
VOvzvCPFV3qcc/2GpMdlz10vxvfcJgpiTZwOs95u/vroC62AcVFIQv/CPSMr6+uC
pp3e2uCSwleLE8SzPhiB5roCAgOTHl+NAOgka0GiY8iUbdB+n0muYrJbtQjYIqwJ
cTydDR3oJ0wvxT7lBf/n5joklwVOAKRq/6L59iyxy8Sfx0BKKQ0tatQ0NimNeEl9
G/nYA0gCFeiDoAPQjmdpR8wroguDNjSP9hGDWktZRaHxxKIqH4BsVce038C6XD81
HVQofhBnK9c2mSiLpG+4WQTXijWbyhs2HFe/A9rCg1l5TDOpU59niVhpf0H+CTbb
voGyunU2tm0FNPOHtWbhkXDl1rspnJykkHrLtt5xnAfQuxgrtwOxypPj+NToIyyW
KjPsJtUlBQnrSZI4OGj2moislP3++Toq2s2J/uG/lsKv3Tshqx7yuwgnFTMF1wer
AcPC8DKwuaQOIPM5P2SbalrAqghYmZlsCAX4OO0mwcYbSQzNsWFgHkqHPCU7grtJ
4q3XMnivlEeeK6Cr3fTb7YW59QAFZ/1pNu0cNbnk2dGgyO7T3BNcVlNkrp7cmdAy
YDCPnn1D6fOUGtXAz5hsl7QkX8ZKqpjgOpY7YQpxKXv+/xerk4tIz+jDEqZ3q0dv
qAn0wya054lPNyGxVUz47vV2AEyw7oSMdC8rAxMgBdiWWANW3PYG+rJoyEIYS4R7
AsoHPvkHqC+/REDAXGsQP9VQDj0Rba8frJfK+pghTlHs4u05NsDkaC6AJN5eDvpS
OLg9twpBLKooKpjZk2B90LpEHywTwPIVfz4Ox3ze9gW9rei9q2Pb8dsSiqDUrfJi
53QZbkgzQ1S59o+0p+jF4zJYNlndqzxiFh0gZDs/JWl1OEEgNegF38fxaKOStb6u
7/IK9R03Xuicn6LsHnf94m7jk2kBsdJ2lz821bfDdVVOCZd0L5ESn/SKI/Q5UFqm
B/KQZFqEbi1jdc8KCBtiY37u4nanHFMIzaLCtgwod1Wvw0YIxF7TxSmy9vNSaNyF
Q8J5DKiw0NkcqO+t3QLGKXXD4qrr+L6x2Q3J2bO1NmM=
`protect END_PROTECTED
