`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gXCmtZx7tYMPa2dQGAwmDysCoAtssGXrTLuu9IBmm1tqhv+QydyCVS39XkxakaZm
TytUdAxTriqaDvDRWGdA1lCUnY4QisBZ0FQVr3wkCY1kS/W32T+nTmbbQKK6XdPs
1Ei5g5OmJ6XvBdHD944MIaCqOlT4WlPJ/2jbGkjCbLNuzSA10UB2PmTChGpekRL+
8lwbstp9nCQGsGifiD9VNTZwu9C+BcnlkjirKu+4ryywzaeCi9eZwNbpCBOHBDnJ
0FzMyMTC0xbVq4rHO3RjXcgPi01y4casDU68JqnYS0NZRE6JyfvDjipfJyzKZDc9
QKW+BgL5STjfePMXeP5YpvkFHon/LZlr8GnsMLJ5f2UAl6RPqD45hFk3lgbjdjY2
Au0eKLHZiu0eRE42KvIEWRug8+E2kELs51Uji0ZjtZi6WC7cALo0K911KsXHtsBR
Jwwpf/qFWf9nBuIey5PXuwdGSNIoAci03uw0ExEIH4fmnXrtJAXs6Ke6pvIe5PWX
Nxt7T7vzlgJhDIVBoaZdEtanq3thjEvyhHzukBwdvE/7dXQeyLprqZ1tNSOlup40
Fc+J23QknyuxxqhV4HtTzRiUEidSOWkR1r0MpsU93MjEv0OF1N7d42bBocf9y7El
Wtnp1+8+kI1GdxnKxZoa5jQ5GId2ZS6iwCI8D4o74tqIlRDgg8SZFes9rg6N6oFe
kEf9P6HTo621pYNMv6m3CiahJ7+y8K2APiKVcQcT4n2+rbENVNQQ1Mfhc/5czwJD
P/ygo6V4KRuEB+/aD9GtaqLpJnxmMoU/mIetgKnc2nMZa4YhOTOEiY37bYg4d4nu
f2K3Q9HyoakI0er0EuZzmAbTeTXktcFgORLqwiV4u4y08CEnkYRfz8GToLUqXRao
tS8NXTmZQkh6HQYGNpZlZD89ZsYVwdGUs9HPT4ZZI14ceTAdlUnZFPze8AxV2/H+
qg08XncBFmF6GFn4edJgfYh8BHVUtjbudVi06didfirtYbVeRHKqqSl1oJCkiyxm
lrBFzVeb6FLFJ+VY4m0ocw+5ZQPvC1+yRE3//Y2hLndBfgIu1WZFScVfniDE351H
S2itkCaPkaUM9BAa/M3x/Q8Bd9TILQBeQbkZorZmpyCHJxJYI1Sr7/nPph2JUvtK
bPs4OBYzTCZI1DPSlMkatSTIKbzriLWIg484NKKgqe2Y6883DnWjD5Dhp61UqdbU
Lbn0DAp6qdAOSbEkTV2pY63tGYrlXc1McdeZ4Yj+eo9264IZ3+biEEXb1VhP+blW
rvcufYj45gOszGGoiUvWdaYtjZGuPoUbMXAz4eQl02jenZqBUtWbFwwGBqcY/MW7
h6vwcuxS04R7u5sb09ZsH02Z1EVrZs1dgHP1K56QLDpXpFkbR5ctQnE5NP0zTcoB
7qW76oMnQoci9BKr3zLBGw3UJfwAfnsKZLUparlfL+7qOT05hCuGRFvi3Yam1TbT
Jqaqc66rQ4Dcx2WBu60rsBV3D+6HCZBHBeHluCNuMd3qWgyBNfJNtrYUZsYNpOXr
xAMG9fYkuYo4nTWvwASkMw1pp3w3cmjjOdx+RP2BAOlnBa3wAvQ/d1iORyOiBkvr
FCw95/F6O7K7wWYyj2oYGiGK62fwWOtmQJIqGrZJr6HiJgvjl7yTYU2uGO9OA+3F
XOLt5e3OQXEj8m/XSaFzRnJ1Mo0fN3A2Gq2sJzJg2NlunF56FJTqgbBEQQ/VSCV9
bnMnIXn9/lZa4tCK9RCXNvQDUvbJ67c8LvNWu2t/DV/sJw4XIPZ56KFwVONPDNSY
ponEF6f0wu7ppsr6KaaAgey/B36w2BCoNEUPGozfPxB0JQkaW2Su4qZ8G+Msyxi5
A4S2U7URld3Z7AnKwiHsG1oENdSBJBUwGo0zJvgev6imsTxqmhvyeCqxYNULNxqo
n2tman0AbLMC/DCKiJAgXC4s9Lodfk4YAH/z/D1Gv8qQawB7ubzpHKw0ItF7pn4N
a/O4s5td6RstL4+TTmv+mKBKWd/HyypPv9pY6qLVcCd7C65Hki5hH1nsQ1M3X/8G
m3rjNJ7MxOVuMQ+mLqdm0OZa8pEMhwp41Nr5cy9g4EbeJgnBsyl8lSFzH5Mid55/
hvQyt4LdlXpKDQ5nESCTmF2d72F6L3K3FUZWm80NohlcAwayYhhxOkpqQzZEo7RY
IsC2cJ8gQWIXQyw7POuaViSXi2urVhwkCttYELzxSwRfoewDk7oaedc78DNS1Dah
9KpB5eX7MVujaOzhBhPjT9RG/kmNXktZb4pRnATWFVH4Gp10dnbnb6/vbZzCLyRq
XwNc/Z2Izpa6MYxYn2fJvjPPTRX0f9jf6VIwHkxB+F82NtweYvZn/svvurXKvJkw
jclb17xB7WxzYT1fNIZO8JtghAnrCTB9leYWrqHIk/lR3xH8duRfvN5hsZ07tJQ7
k1WBFnFu/thzIgR90nW5JRAKRaa2G59toYelJCLRkKPnUC7YbjLCE0fkMUo7hy/R
QHfGNPhpa81EWzonAfwV20mWRppG3V4rJXVJT9YobqEHIV0FQF0CzkT8q+g3ieaa
fVctfgmHLwMn8nYuThQO+HJZrxuaE18qy4RLpMbVhCWHPZNNMuuTxk2kqheTrCHl
ztQNPfyMLKRYn9dL2/f/Zw/3A3tmQOa4rrmHzxcWJ5S+VJfa+y+0s+uJEnCJBNst
xkPad0b7KAoyaA4ZhI7VriGz5aAQr2gSxUTkaHbmLCteSgXLQy5bFrWkSeSAedBi
h6jYf7MKVJYco3TUEvwdjZNCHql7N6aDUSJGz5gU+oGNrNUdZ0zND2g1t49TgM5E
mmugVKorIvQ56unwiHrpJriLqsBBuasG5BkyWEzJ+ZKKM4smeG78UtROERdRJOYN
WfaR27FJEi97Z8xVAOnNryP8558rnQ/HZkW6YsOLCG5QPR2UM1PVdZFX5JEf1Txd
ADvVvrq2ZdOwTUuwfRtNKpKvqHAhp/DNU69ehkMu9W/rkkFUtRBxNNWbLhwn8O1Q
Ox6BwiU3XyVY9ldvDNEAMom9Xc+MSxRZlA5H6pUrHbnKqCuNpWXzOLpI6IZqcPLN
PwmN9AE5yBkyZWc8h4z+fwdQG+ycs1HEMV7Ww3o1pOqbD24Iso5dSsPuOhsCkTsl
DihtzEwKuGFDpIAA3OKOBjmNWFEZruM9axq7OpwxaxFWdehG+Y+pam8WTkgO9+0R
0k4ji8zupUi+vvSQPvTpMtLWdCGsvdhmf/+SVzI+AlzJuIy3tp/oQvzW84HLmD3F
K6qGTPFQO/paPlkVBQ55Ok78L7ZTKUXb00jWU9GnD6EtO2z2Ho2rtZztCw4tMDaC
pchnkU1geN1eZyFU2aeQ05xHH0Pcag1ol1F+7vVhW5dridI2yXeXKkjXm4xuF14x
AzEvLz6X2KCZ2v7rkPvjq3rCaXqca6v86SC/7ArZbveA+E/Zw7HBvURs7J/UXDmo
tiNJxLUgjr1fl9w/th7iRTU+gOap+FaBgadaJgj+eUKrGUai08htKWwTu+a7tEz9
wdir6+GomKtoH18biZTjztDHBLrQEEF2EkV/UoPrxHfd9JB+fifd3U8xuAhoA4xM
KyU8zANrie09r3UBxra05ZkFjbB6UnXi33UARvHBWfsle3EqmubjNWWmADYcfwiN
pTH7g30z2UmCM0YXJ/NJjpc/hi446hMa3c7CxoiCwFJUzkbXuRKe+PRuvvmeQ1sT
gDkSosRDMArbEix1QIqtdOqgl6ueHaDJI8U451AYjEIgMs3TyEuUklErGlrM9Hbh
9MTkRQjndhsNobsuFIJM3MpeEO/Nuxjtl/tv9Tsk/n6dBiYoCiWyCThVTtzzvLIv
Bkmsa9lGiqzC5VmBvD4zmYH8gsk1NG9GFo4wVH4xLmTHsOgVuHsz8z3xUuqWmOOK
kRqAufxvHTfsEVWRbT3W15wCbr+dz6WrvAiIuaaEvWi2SvrDCgzavR7cS+FCFg7f
o3q9zGtcMDWfkXHNhZVTY14CCqNqhhYCkcCWMxXIBHGVKIHtOapP95ofVNstPw3L
ynbH+Mxek9VRBgATwOWlhpsToU21jF3tXFmPYrBSSxC174tE0ZjzS3hxA0x5HOO9
7y3lKhFE6JdrxZIvCkb6l+b19fxBI9wTCG+fHvGBHssXABjz7GItghld6DfO6xLA
shsBj3RNRiW2JDXhXBOKOuecsPRNMCH++QZ+zWPahlNHd4GiHiGcRzaF9o4txebx
h+xfm4MeW7sDaTiqAOc4vuwOUlKcz9iGcwgqtguQZ7deOdLL/gYso2C/0zpGa17c
mTSXOrVNtTOvfDqUcgj8Bd9FzwaWUyBLqtbYd0hPtmhPjakFGYSdSr9Xxj8o9FWv
Cf2ZRc5yqHqxox62SlxRQld47xK1mYgHqLwFADszkv4oC+vrS3N9expZgp6/uhTY
w3hTJtsDofdn5Lk07zXZos/gsomBi1RFdxHht5yUxhPejQJc1Y9QNZ1ATXRPjq5Q
uHmw0FFz8iopkIBpqEpvc3K/X8KuQlenvRO5DjDciLnE7sHCkvUlLc5erSX3Gl9l
j3dqil2zX01lPuBy8TMN0/22IKPKO+E8FN302j2U/39gR5VdpWvtRlwPSISPIUc7
2O3PSCohih7gtqHbBO94mSWrVOorycBAcnGA0UemS7eVwBLJZCP/srEccULQiV0m
gFXsUn9uQur2vz5DByvn6Ber3keyS7Eo/j8EEaDQGhW7SlKwCw9D44C0bjaCmIT+
6ITsqdZzbf9hEm9U6M4KkYQQ+3crS6g2wHXNqB2IQmKNeIt0uuInVAHoY+30WTKR
SeBHTFRkk1RjPiJ/h/DV2d43GIs0ELdqhUfSwEFjoJOBKA+oPPfVFg+Vr6etoFjd
eUqreN3ke0WaxvZARBKnk6wppkGPIEleTuvSbrb9gvOXBzWA+Eu/vvcsWlBzkU9w
sONxgylJxJDBSZVWDhte5vbg0aUTGxpBUVR7Qcz6DazxjH3NkdTNoGX6dTEw1KBx
SHPcf7LvGmwECn8wQz20qZYG9fPShNBzPmiqAvQSyY9sbyU9S7GZQEJJr7cvoQ1V
bbWqvLGHCeTCINTgelwn3MNUo4i0sIS/n0Q9dtNOlvY48LCDiYVWglcWqnuhYcWQ
YbVX7SqflsVzeYAH4CyLAe7lUkaHj42wQUYj+hPmGca2S9SLCrco397eVH3gnLsr
K9HqIJwbLlxgipVUQmrHApNwo/tPhm/Q5iNLkO1vKqC7VRtQ5jVjPgJTwx8GyEHn
ecJcpD1NFc9xQ9zPknM1KmVTKjGvZUa8KOll6QYQl0/zr8Fp47hEv0jqY+K35o+n
hJ4DPhFztJ45hM25IDgNeP3ZRD24UoXmIRLyQ33StabeklC5G5g1qf4kCdt05oWj
ggDsTc6UK3dd8sxK0L17FZbsCFXlp+uAM5vCaFF9CSGU4VG2FYAh3t1R61YXZnpa
DIohIbCzxk2ItKuocPxAlIyo8zjrIFnVUqTOTzzgKAn9/Luv2XYmu8iVwaWj/gEY
WRoO+P9PBFDEa+8EkwA8IbFG6AEQOptK3I+LGZx3Rr67N5HZmXt6h9ofC97O6nAI
6OhT0o0OTcEzKjJjvvmMr9ixvWB3WkpZz6GNU6q8FjCGnn8t7ZnJ0Bi6k2jPA22I
Ah1wbuXX19syYtqzR1oY+NP2ONTf9BWO62Gw8FKcMD+1b1vE/t2tFYXo5HysMmZP
aSRjwuwOQgp1Y8bpMc3YPDNgLJ8DTF1mjDBfy+Za+1vu0BU09eGhKmyMMV57KMfR
/yKKg+UfNIPvJ36S1/RDZ6iGmyvpVau3F85hOnqeTB4ecvISYnqFvlftAlAjdh7l
+KuwAtMPYWsurL8azm0uCtjE0m7iVoywZtUi2/KTu4B0Hl58M9fhMZ2xsIaq97lT
B9jGHHt59EabXOU5Hefn8GPoJbdkz+8/W0gGGaRdZRCrXEoOXldsuKTuIqSvXZDb
y79jmOMKltSDma63BCf6BVyjYURYdYFFImFIr/3je+eg2/2gMsr9FnIjpxe1bCf5
PlGLbcQ4d+rbjShLK3P3iLJXCo5XHQX307oYI/4AQfq4dYbbPClVLYlDU77Yw6v5
5kKJyOFPdAZzz4sFXfW1RCczqC6dXKeJ99L3wj7dc6o29OMxV3++WYJQh3Agadb5
8rX33b+dCsXOyvlZEtvbhWqtjkRvjHBRH1Qe6rzzwWmTZVKr5Q61ky/HE5ncdi1t
2UeP7oUie+6wOxUzuQtLDnZOHO3ldpBVMHLsF7KMDA/Zja+E7pDklxFwmW7x+lfD
ccZDhilcSiBEL1SEQIq/IC82pk0DKepfbC16exUm4VjJAypxOfWBVzMWMGXJN2iw
hFQy3BnYvzdLzaH6RqIr4N8ujZikGh49aWoNikSgxVATzjt69hEwD/WLzUfjNrNf
KwXROgtVq/YoB7YhlCNVuxPBZuFDDng07MnSxHaScGxxS6iTyCXKgGE/+k5LjT8u
Gx1zDBYf/NOO3g4dMqDezyEzIbcSkBTyCoAKIp7L1ZnvUMZl6oX01/4H2KdIjHmk
Ax0CkFKqFR4jKZrfgffNBZpBlJcmYyH8b9iGYZNi7ekUasE8dY0ioMIuaCl5soAI
rltzHdrNfnksf+08zhInmWzi1mj85/VuOLClv209sZW7+PJBFcE7zcJnj762ty28
7ZrzoloI0Evdpe+OTLaW+afHNjYEKl5nrT5fXw8vh5z/t/hfszLPrOs4+5jRmMGR
R6VEzLkTkDCyDm+ccedTFM5HkM7TUz/SKkq5/r4UxscxgcSeij/5buJv5Jr9994k
++UrHgQYOTKPW1ynJd9iZL0wxTOpNAEwfRL65VhZxJkDq5mv69jIYC2tOeWhOluZ
MrMnMxDWQizLve0qcaiaW8bBnsvN2mxY9sV8GHL3n/wD9OAhZczUUt2ALN76ilLW
Xy3TVVWulDDxYDHDu2Wf72F8R217eUbxoDOX49i7gKfveAaYrx+TAK3B53gRcbjT
kfYQmOvXAczF3+86DFQj8ze/DxPmZjSiGKmgBXRnq3EzgbTmZ7t95Y27QDZmvPOf
vfvvTag2gPRJj+/GURcU+N3Q2Nn69n5nKj6SNMGEZxlxQoZF/Lp9PiUnFEyAtBIs
RpNsXr74A1GVrvVH1MX4+R5eJwwMwquGGeb5wKxk9MbLm0wXav5edcn1xJjDEXz3
1HfPpwsp3WSIksO5A4WCnoR9YUnuGoGd3s6GgSvCTFZXpoi5Rwn9Tp6KHCbinVLk
LcrgYV/vkAucqyWdka3NQwrmEp55ifIrvGUTqaE52luyiUv9ZY/DR4ZsAGypWe86
XiXvhITFzeYMSqptLJoLzZh9UZb0FuoH1p8bPL4ACxrnDu6b04OSUFjmPdCQNoqI
zW9ONSDmwC0UDx4ArKOlLKoRM8G5IkfKStvKNJtQkFJzCd9N4/enQYOIMcWpzBkv
n3Ck+02ow/xgAUv2Jhxlr63CyWsOaeJIKYmKUYX8SrRZvMaGIlE2GVlOp2dUJrlk
zENvzzkFQoNfXE73H+BdVTNddfGCf7hxIgVMmPZnCNF0PJLfMNQ/18HxLVkvXX/s
ZvCZP6VppogjQ/xhN8uXgZHLBHMOqLJIcIIRIKyBJq1Wf00QOg05eJ5c0t0b8Dek
aGrtC04Dj8t2jORufa05jidNnBXCMNIBorxfsAPf+3M8th/w61z2TeZixz4GQZ2k
mYsZ1zh932pFp/LOO7Mm4cnO80k4oEmfbmBLP1GdL282hiIcstF1W7oPrY6vq086
coe1TVlHVATCtzni/MR6Oufcrk9SNM8/Xw/usrZ4gsq2Tb7NBEg1MKludv1c5XSN
TyzwUtNKYqmWu2fdGxDnAQz5i+2QTNu80t9qvu3hJcr0u4X37J3dnbGyZj1CREfd
raHpgqbQsMtzsAB8U+stTMAF30/b9yx8LPpGJttTf3ETM3Waum1Rr+JIHQ+UT2dn
tXDSSmgQof9QDy8a4TdsM/GzI9uTVegyUlzIV4fXKy0LxcwULi5B9lNhACJi7+Gl
oOIROI8wsS/7dWmlF9OxgFoOzf/3oM6oKaC4Nb6HJZdlgdsGhP+tH0nqxmYywykX
WBZNxmVBFWfro8Im0vl1BE/MkDR0Cwah8q2WXj56wZSklIDeFoUnVgkTV6P/baBP
Dx6NlgEXlPxPluBMGR+rkLA9bWzNrYb5XnT9Byu8MQVLxfRiAy8TxaTHZlOlenZL
0bB8U/mnV+TRKlw9l6oTqVVCqSLrSSyBC6FaYknaY2wxRM1vhDyIIUv6kQEeydv5
U4DUPLByUesU6hC1MqlxMWh6DIFkQQtFn1LQBTVON9itidpqxLh+T2/oF2aLSF0x
epMM6BNZ8d9nMiNr3NRhhRTgmYEHwPwEczYk/rP7AF6m4Ycowq/mZHN2AjQ/9jsZ
6FfmDvvLpZZmoZc2CMVcVdk99Bu06gNrDXEgEflVeN0ut6iUzyQqUruWp2V64bg8
G2BqSQsJD9tA+u87SoPFxeBAymzKSf7TllMWXj+ZHBOwofAxqW/vqxJ7CNDlwa8p
L74+/U6dFxX/ftyPyNzIVqFaYMEASit8HHUXQXzy3SR3Zdsmzi1V1/5gdFbjQKlW
cLCWr/rVrgI90CTrLNrg2Ct/ju++CKfMHXiJLRTnPTN4kk86B5GQ3ZpOfUn1Augt
fzMJ7h+ewj7giDY8FeT6gm2ThOZMcb9U5JZsQHhMj2VU+MV4IUY+/FdUS7/3nAbz
8tTCPD235FW/bvq1yDBedWwk1OgbVhgqQwSBHkxu1MRTd0fiJsTd/JG+vAJO7ITY
oFnvlecK7xv86rOo+dtL1/LAU9YwlwWBdZoKnQzb8SxVJENRbap5j0HGVLc+sZ6n
jxFCKdbdF6gzRrETdX9P1XcAkG4QXP6F4ZAhwHtegOjACuwoGQk7fZW4AKyKqH2E
WwsXKxXa2YJBUU+K4hQ6mu2zoJJcxjsSG9xSJGKcGMa3hCnjOgUgpOwjYhosXFF5
Hl1s7Naj9C3R54yjRp9Q6uZUkoUX3y+116Tui0c1qRP+ytYSVug/7blrBtMAGqzX
9+v85ExrQEpfTVz9Tx/QowbSSEJwqda8wc5iIUM2ajz5xliU8OhXghMKZzNYZ9ah
m9YFgnRNWM2dIDTbRlJbYl6PvlLFDzp3W0ZEM6aA9lGGk6+l42NdFh9wvDaQTpjJ
kvq3NF5WkhHlsxLQOg3xAVjiPXZpZGh4T1KlrOzTaoF1mWc8vdsPZjkuYTkOjfmh
QBemp/yzv8Tm0DKcU7ldg+wmzJz6tvvV7KkhFwcYO0lvE0l6och3NxlYs5TYmSh8
zh2aCPoRatIFB/xmGno7YQu/KMhNU7YdG7MLdPYjS0ohcTqEpOafUhUl/beWirD7
VDWh03y1+leJbZMDMlGyTPzThkMfFX3X0dH2bz2y+tHUTfmJNqraugDuFb8J/rSx
DZHDtgMjzdCtgHC74Lh7cgHDRaVZGPyEHPhCmvf2Nif4GcOPv+HN0a9co2+ZVTWm
LqzA8Iksvx0nWVY5EuaWSAdifPOC87Vlp/4PxKgwFt+mN+cyWpSAcaysZeZQ5R4k
LQnklc4SZS+3r94u3SP9Z/JISBRKGUyJ4A0f89lZBQagJO0UQrkRS7VOxYdJAeXZ
Ph1Q7aCKMBlOCpj6NgJSnNSM+dqkBl0iorZ11lyasn3vsRXXAIQPydyzTGXnDkXG
1ZmTIZcNKOscVFs/GlJhrt3CIcZvuSRVWTyn+1KT9vxnrjfrmxYbgBAsuVoxcFUS
QZjtOXAUOvkWqfLOE5cQ9Ii0f6THrgT7J7KTaOihe8FqZRuE2kp3pE/w45JWPk/D
16teeUsOjg0jZY8J6Txtz8V/y1M09XfHC04BiTiZLDAICEurGkyvKg4sB1u/GW63
lZAabpJWiXmrctf2NwRzQ0Au/ggt4KQe6qSKnTY2tpArEYIj2YbsohS6rUZtsU9i
+d1yfARdeWY6iuB8fXlloQ/BqaF2EgYAXGXwMidCfQvuPxkLl0kDzNgb8OMAR8kc
9caCQ/oWaQ9XKWfFcY9w/JOVDTsn44UzEFFCUWb9L8opSN3rcJCftpYQ339NvOgH
vapC2Lf7bwZWcrrzEziWuYnhqEvtndVd5xotfMh/JxvDimzeiodxmxVQSrGJYyPT
zDQ0YOHeEVMuwF4XYG/NmK8E9Qu4peL8oiddH+8/dldCqY+xitrlwOIQIMuKN42j
OSencb4M5GjR8gvMx7RqD3vPEi7QJ5MDnruYLXtittUqJg6FFm2fNJkyfsvXMSUg
eBDy+fYq8SZ+3NN0b5WkE6yPbfcx6l9+KneaKMjZTnSfMfXjN8YauunSGvAo8RiY
avWKhvRJxHazFPD6VTEeaD58TiocNCuVH/MOCE3J84sWlZl7eszPkYs2l9IkkSj5
z4m3EEHnkCvWxEcet0eyNNsWATSkjHCZnssBSynKEJCJtrIWNB4y6W+j0n4LmxUH
iDJbU2JfxA+oi3pswd9LH11W0GVowPIn8vLnQmyKeXey5fS6D8cpmNOyLRTkOeYF
dTQz/KWUk4dJWGEAHqUpdsUmL5LyNKwLicUQOikXDS20IaRhdo4K1tOUM12yrlZJ
egC6f5O0a1hU8BlO6xzuScpERqrdUSbsyip8bcLZJ/aVhaXLAbQOn1KgYkj/DKtZ
kusYBrmD9hzd6trZbQwzTkpGZDJM2DGFaL1vSpoGa3ddfk5gAShKNG7wW37beiNA
K8XZv3Cx9ZxOtrpoDv+VGI6tycLsYYfzVjTq17GPEXh09I1si9rEwEHZ8BAB32AD
wMaowneF7wlB15LnQ94b1a9nBb+vRB+S0MTGmkq5wx2jwfSrFfz2CzGZLekICt5b
9egn6P+3rC7yHc3d2cnlbpjXF3Keoisbh80q6bfwpzPm2Pjg3KOfm59P8zztP+iA
CJweqJKr1pR6mXwsvDBS6Daz/WJBXMsXh0f9pqAbCK9RpWEqK30w4pDdeF9GBzJz
T55Q2aLftpsWcAfyuKM36WNqRfIC5KzVDQkqHUr9MWHeHPxNoiKiXe9u+xM0HIGg
gZFqJz2BY1Y1Fhnhq+oLghkD/7s+K1lM2Q/hIQLmJ0P3cPTn7C+V4x8Z0+w7RmVk
bf/1Lap/P4QmNjbbVzpTx2h0EsiUX3+289250GrsWGKOwbXVAW5/qDxgiw2DHphl
rvsmBvzHBsCFNnk/evlzO4+xDXw0UAKDLt2cl3uslYLVsLHf+8pLmfCqwEYVB1EE
3/9/4id38WN7e1TD5Vqe1yDbdAM3AKoPiDj3gle5DcZLdJ4eA7UYNaxiDjTWYF8D
4RdoK0zVkAVyiuUrhCtOKoX5TjinZ/xbwzTcnH14rC1mMZw8S0ZZHJs8Cbb9xeAr
F7ZOBo6Pc8F/aHRP+OIXE/0c/EMG4HzaUZi5Yyp+IpeA6qTb1j80+2/OwS+Ad32b
gfdaLiTPno0n2C6MEleu7oxEQRuJpOHB62rrhJnCxpLRWQz9FXRANty4Y8abYvLU
up5FWtl5UOlfxcNKgx5S8Dy5fK4u1G3lyqNeOrmS+xpkfGjHuma2jM8Szt7lrOqq
Cfm/eBwXCGCNFb59tEFlbPwE50c4OgeCu8gTKCVqm7NnCYHpuH4OwuAiDx5+aDaU
0lSEUaMo6Y9sVdt+rHAViZYiPlHKREy7mU3ogZp9Rzc+5bIys/Dy32Z1D2UL59fi
xYz63PvXyc6CBdquOe+0znlWdnFh3zMkp3s1EMmC6JX0e/Xn2wCRwqwJ2Jr267QE
RVMQCH2PUwc7X5SJFAcCloxxZg19zS+boCJjh7XXtKdvIL7j7JK9jQckUqa0zAwu
JoGXyWXX0RXiCgEw2g8FWGEu/fU0MvksSG8/GKuYK4wJyh0TfgZzDJFoAlTgoz3a
zxZ8I2LKXvxk505M0u8nikQH2JoqfNRoDEzsy3bWheQnfsOb1m8KI8iewansdMd4
MmYdXpSDznTJ1TTepqzRxf5eaR0euIjiFHJGgCJhQBWsr30zww/CHlja5i2lyVfl
PMuc4TDsN/KKuKiXHWkFT5mS+/0SfuD6YWbEXRCXzNFVlxdnOqLNa9uFThZB4hfR
Hi9eoEBGUJz0FNxZCgJGjCn34He1fAaEdA20DlJZpfI9pVNGMLXHQaQQMEaDCTbw
X1KfOTLtSpEN4gL0kFVT2gGocPiQlVsny06JsoR1+zV/sEWEFusOFuAUpjlFvmZZ
Yt6OmMjBuPvHWHXywAU2kO+zNb8C2js0fk3KlSSmK+vvykOG+SZjFn51lvrKveQL
5CP+9FQ1HxqYPHudZKS9Wtum/pxDQNOX+O/WcwxZ5F6IXFJsdQJ+xqECRjSsoAln
rTfxXw7686A7+q0FkXqYnYcr2Me3Cm6+obKHoIa3GRkx5QT/p6EGm42+QtnKggx7
Po1UdX25reaTnY8V9jZI8JDQxNBYIZAnKh/u6wyOWVMU74+7c8rJCfULyxOHl0ca
3bh2ZX4BuhoBk/nXlpdMGAU57xNdxWQhOP786mpv0wBgsI+Lrqu/bjJ3NOnVy0EF
+r7EvWGbRWVi/acbjHxNWJlFS+nl6+xCIpBbjJQbMM5ZTM4IRq7eAtO58K+xijUj
L4D0O0yWtRiMVqGgDF3+YmE01OYXR75EST1qwIoPG8947TK00ELBbKHcf4/xCa6b
p/FhP+KvsEDqRGiv/ccqQNKidkwpTPUeD9FFHHndvQBD2z1+TLiebpcWzKcgKw0Y
hamZ2oPNIJ6IUjhkuDLVYTyScX8wPnUl0lDjGQEguDhTXoZkQa+AC/koZjZ5EAQM
nUWgjzlswTXqPrqGjKqFbXDvrp4A4ZUrUKoQKNyr0+TNy7L2rasSS1F4pKpL1tKJ
QG/qpt2Swf3OVlUgVxJ8mM0CZMnUO7ea1rLmkda2ZKzRmAHxOVIGC8dBkukTZ/KH
SugHkIecj3EBd5FPHeWn+TEJ8OkyEqxjYzpNJ68uqHx5TxYxxbZR695hrcbhtVwv
6DTsSM7aj3r+1Hk0ECcLsfyiRBiSuD9kZr1TgaHlS4sYFAC3dmbx71p8iOxxqmKY
n847ZWk0Ajn+bcyvdx0mDJ2lC7q88wERNBVqPQ4ox9TarnLjiJXZfzSHiNjxL9Cz
FABGG6N+uTUoSh3Sf7KHpf/DVPepMn7xqp9XnzBSsKFbdX5eS2DREA5S0mh60sUE
tnnqLrTrOLhspEuISMgPtxH7lKfmk0EPluWspNNQ0WajLCpu7f7KyCi2MqwB3mlU
9OFtWaCdzSopKj9AVxSIVsvV6CPlN2tGXsx+xF6K46X2Su2R+R2imoc48oPY3VAP
66B9+Rh6qVyp0YciAz8VVQmdDNakmmUaVm+kWIj2x238UMSd4zu+Bi4t11UjjOtY
QyS5bfuSqTDFXSW3G5VuvroOBfws3TWIEUeTvMJ4F2OsheXky1yD1eeVoZYMnPZs
GogK5vQYkAOZWQe8eCCmYps9fG6e2/DNo6mGN5DBbciCM+S888TXJl3BUWv1FIsu
/EtPtAYPW8h6nzy/Ktr5nic4v4Y55ht3JPSpxNcgGvAH0sYev8WqKb9kH56RwYeR
9zerFeTaQuxnXwu6xlz3mMxUih94f2QIpcEmhDjB7aUlDENyaVmo6xzguzgu+wHH
feU79x+w84EI7sLYlhiOsJDaTLPJEGoMrJAh/gWi2xtEfErZK2ZG1A+zobSDT7CC
bu84JtnDStN3lUA81urDtxDTV0s7BF5wCXLcoOKPcxPLd3FYiPaO4P3YbszNyZeH
59l7nDePsBSVUtwcPmaNzJXAvufe7sq6EIFC8roD0BpTx8+iVIL1nKiPbqXZJ0aZ
D6j06EwjP0PaxqIRFd9RbfwIg1Q45vSVHO9N0CleKqW7b4TIbqIAr1LkQZxfuwS1
XRlFGOPI/fvrtzrnxTifMd8U3tiepEj4Q4CEt6+ccvlCM/vtVWD0RKYReGd5HZB1
1phApVQl1JUuLlBUqHkpU6w3dkBLjjDUYEbaoecPSpx+g/tZD/saQ/O3ly7OAq6W
03aCsl75RGHhcd/zfiDdzdj15v6KQH7H9ZyLP/MKZDP0UhJuI/axeluFUWxXWVoQ
yaxiFz1LB1YQ8GTR98N8zxdede/2E7STnA45onkiAC6SAwC04ZcU/SCZe8nAvEqA
5XG/BAbGKjrBZVo1QMLPX5aj9kCLnTE+IM8nVALqgRiaCjlrPUaPrUfxpQP9ByLg
ODEh1n0cT5NfxY1ul+nxtQkodt9YkAaxyS6jZPSIUrtH8RFk3DJewbqzH3x2z7uL
9fVgorjIyELTvbUxjQs0fyjoYDFeGQsv+exDXbGkGU6VEih1TuuqQbOBaFefbBtj
TeC3i5kT682BV2Iul8MiicIrFOcoZZKSn7Nu+vWXxElrfxOv/R4dspKQkQXXyrGa
G00tCuZ1URoyvBxmiZ6w2sUMXU4DTIRysrKMBSTip5Iz6GWXccY2SM7wB9HE6CbO
eL8bxoVnYOhHMdb6JGXvKKjmzAw9pzV5/RVfuGBxNRCkR03R3ofCWY5bHnxlBDKx
QvtirEW/iEBx6YYmgryabS2Yr0mqtLMEYDsbosCW+bMVkzRsG6Zd0X+WwDYU5Mqv
ZvPnegC0yOgtUg5x2e3n3Q9oruB0COjcZ/nrCzMG9hUurgVaAQvGCsLGI32rzWrX
q9o2I4Tb9BnMGI9tIyRkLoHxY1XNSxxIyvOm0fFCcXMjZ26ZbBQ8vHlFmYVUryKb
PAKcs74ExGaqt7HyaKkDrfJtzGw2JAXARuei0ACNEdl1jC+FAxAOXKqj3ZR+nkqI
JoGSpakfi4dyEVNrsP2qpErRJtvoifxcVLs18MIQH/MPq8nQs+/q2P75g67eXUGS
N4kjRFArbqjlVcl47phPEP924iRvte4QsdZTYE5X6D6UF/LkWoQqAHRNL/b9uq4C
g9/ZULolNOXrCUlw/65xBoRi2dnQ1eOspcnNJBB+oV1TNp+p7FEIx3dtYcO8KhYD
/g/lS09FixFBD22Kc2ltdTqslaBAW/tDyhmn+xmH7UtIxUgjL8ne4F1vFMGuIl9S
FnJinF20pU54+Yt2x9NHF4T5ZJG6U0NXTnA1Tj35grBkkEQeIQWcYjGTKYWw/YQD
G+Mt8tyPFILl8jiIoiOf7O/BpxxPriugTmHnrWGCkV6Gcy4OiMFowWktSVfuIldj
QR+1BZMW0WdPT+7XtpAGd4HJOPmurWJvL0K2oAHG4y36OSiA880tMWux346dYUMw
pha9EBWBTRcxjAmHk9tYS+AnYwZDSC+GNFX3MbMxsGJkQS4NDmNu5t4ronQhDlJa
oLAYej9t72KrLT72Lj+FlQd65aL1IBD7I1qfTNhll7DKFV0nOAs/9eajzV6IjO4e
3b4w7CCb+MsQn8uCqSG9Zo3jWsKZhOteToWNQKY/dPVkkf7CzT9UK5H0/h81mc5y
iD7hJhz2pTgViC7csG27zJzvnqtSGWFzRbPyZ8ToBnbWL3Yn3N7sXrt6ponNjumA
UHG8jVnd0NLrEdY7oSlljsBeDJZZfWsVR/LEPui40YhSp8pTF1zJhe4ePdTV33Sr
lNHg8rZbLQ+3J6UnKaBbV/n93+dT5OXH05pfqlBxD8b/33uYF1HObDa9c0/2St9I
Y+ASmJ1FJGPPpfPB03xKV9Xd4iUNiO8jMGUIn+e0ZF0g+8QQy/3Gw5rPQP3cmaEq
4yFj/9b6j+2WvXEl4bhByZWAt+2Sw1pmEzYpgAwPnSi2AIXh/Z6GbQ940A/1AT5V
5BdzILOL5eF9xlCmiU6anJiu4J3XVygIdBclbQFchRptdqdlVJBSH91FxjXZ+yVN
MTvb5sY38r0LKvdV6LUvtC/IMpLN9nkYjZP8vklc6t16gBfoNzlKxvoUKSMlKt0I
aJWhioqJWY74qWs9S68quo5vqqBZ1DRz+12DgMb68AHS+LudBCjfBw/RPy91DWHn
6QNb6hF6vrCd1p2YcE1sj6w0dFjMX2ynVwRjoj1I5Tt5q9ytBFqnVeUMCYbjO5yd
UUjalvTA0LZuaZCD2qLQeqMqQAYUc8d3BcPy+/cgTsvJ+6roZWOJp7GtUm56r0zh
IvguQkMxLMo3oNyRfIeNn4fIh6D/VmlHVRKgkw0cDuvm87Yz4OsJdYfPbpcfC4sJ
HKOJZC9jHEwhmCe3sdCIEgAuCFYdZkXhkUYTXq6pK5fJjclN5sYTqQeinhBo5FHt
uHWtMJpySR9LE540wrdvc0Lfhz4JzC30PqZ+7pRz6oiQ1uKZmT0lPBlq9xIH/nzM
ptOHhCDgY/7ZxiKCI8O62cc7NKmuKdKJG9Z3Uqz79+jdgxcJT+qYz3MQ1Ugy0qAi
rJkUkfa2AQPXPv/R5lz1SpJ+oKEdHZCbVkCJtJ78ME77pYKk+o8SctGrLhcPl4mo
tDIhvxo9Bgiw4dbwB4kdmB8XrU638XLBPo4hsejFXyMPDcmhS7DIUhRCim37DXIy
q8Wcqklbbboiz9UHXe/nu6XHiRL9ayeRUT0gpYxny3ff9+uZTwTL9O1KAz/0+YnD
XhIcuHrrcsI0Iz9Quu/ad8ckAjzDm4W0fKZNyQgTIj3wOUMbVWbOpk+Rpdyl5Ogj
f/3XfvSxJh0U/UQCSPDlFOia74V03GhVjCsPsSS6lxq+cDN0Hll8hpZDl/QXnn88
BC3gcP0041ynAJpjDSyQOp+SP6RbuR8W+23MxrRMOhAwm4Cok+QVYneJVEfKrlHP
JLyAzL/zA4rvzGRaavYN87Z7HhY5b3o5D88tftQ+PBISydUJWmxEj9LBc6AvOZqg
jaMTQDbwPneEB4a2TyloR525uZJr1dMs/wYyXeqdSrn+vZRJSRc7m5Hi8C8+j3xT
/NGDL2fL3NsmTV9hkcNXhOsrbNvkDttTGqIPKJGtvYXFo+8PQepOK4X1xImQ9HuG
SVJLVwgoKA/Od6elRbnyTF+fJtZ2yEWvu+raiW3HkuKkBxQs2FSPcloUoHyKVVH5
V0/h3qq1pcJWQYjm38GEgHmGXZgGTD/CDj4ipJA9bsmysqnXTz3+A9pFpj+aT9Cx
aOJEPlnhLwRE47s+NcYgBDCqQU61z/n12Twbw93/gKym+SBOvm7+AxhuxcaG8dF/
3IbZ3uwTu4PtjHhmp3LXwh0Hvj1bMCgrlxsmOTxhsyll5RyGP6TUk/e8slS+pHGj
lMLAy/hFhZwPmrb7U8xHGtupMnuql+GOe0o2jufaGhcb4OIyau+xhT7re7Um+2KK
/uWGe0kD2o+BYvQvM4QzCeLTpEC9KU0XVSHLhHyGFvVc9aoWGIgBcymipuGsVRpw
mGDB9zEdBJgpqP+7MNJVBP+eJHxxoJ31cPpZqmBzt2bjP6YwqTWOwXh/tZQGcM6e
osO7uJHhDyw9uViG2MFNZANiiMBF6ybc+3GxSrTvkiHHtuQth+SOYRRN0sY6gwHY
z5wa9EXmmvzIQA3xPY3y/NidhctuUqsY7zbs8C2WnsyR2x1uNm8j2saAuZPsPxnH
N4KV2MkZXKJPn4vjQMj44viTsE0pelh2TGhxvmXuQ9tz2zfy9/f0wgN1lSy4pGD2
99TP5TlhHg71Fedf853UFPcd9dHhdmPwfJtFUnpc3HQei5+0zQFlW3v9jSQmcsb5
vT9M7O3jzK7uXyCOtBAlzriBeDxj7geysH0ucoijz9nzJ5UiF6kdA3jYQQ2HhopW
vI/2JCKrULrQjK3XBeNUDy+wwoadJ6chU/+XWa/MQqpr+L1CjKigJEi4KdEkFMdO
Y0CQ4QXo4preV1PLOqi7bwwTxA0FB5jIVvL1TEsewjVU5owjC7v0WMaVZJold6FE
EFaiXVc+27Hv13jtCSbewWy9vVUJjEr/1iNfFsTQmK5UVNb9YPqFOSyv+q7Lmm1h
q52rlrwJYqoq8SwqQ2K5Ai4U1sei/FhQ9l1WXM4KE/JaPBH/0SkkrYQhRHh4TD6r
RrzaVrFldsC6dxveIMCPW4JQxL7VFiwi5iMQk/BmNtltZpaGCmpQ1x3gfJMPBzMs
kv8zsgjJ23r+bjiH4ZZ6Uz14PpirQWiya5ONzcHwEdh2nTbyi66HXJDrjgZoT666
V3aZiAac0Vlm8CKlI0x1OLhkA4aeKtjE4lWOV/bXCeIdhC5q5nCMnsnGJHWEK54H
k+HOTeiEPmUwCv3iSzhYqfcbQbPDPhlkUD1mu44z9vCRQHQ7YVBiyl7fmhT9EoEG
11rRGXX+htdz2oGk4YpoYhauPLTtHG+ky63QKzh/phLroQyb9M1F8wagkMKfAzhA
nf2FzulwJtiwB7ge9l+/ufREvr8PGku93lk17sKRGGlCc0sUaAI7tEFDb9s/vNFc
sTGXNrwto19hbUtjGCoJX5CHqhgs62FL8ToNCmFwmBETOoP7nxlISZCrsSffH8AE
KSf+IqksfP3R0ODb0zpVuzEfxdjaMKB3ZAHgXhFPOo5EvUGx4ZvSrqhvhhaVimMy
KRPmka4bkJRNOVIxsFtbhwBjmYsPHv0cuH2Ji8eQbwOxeBA99S6ebtt7sYt3VFWi
bmVjN39tJTeqyPYJ2NxTWw9A1upRhTerWIHbS6KpiPzSchwIAAnEGt/pnNt8ZLbQ
rfEtElh4k6np5DtIGdPgdiZJI5uD4ncRqD6n3UCoa6psVlQqk6+cGfjFxYokLT3G
K64wxIICpiquEHhAG8T9rRDOISGhQwQaVqxDTTvsKHD4TzM433aLlnbEkgHctRZQ
8A9ssEcsIdSox1PJ039eJsbcPIuK0iHkIyGS7F25+8eeH7cFe8fGEv6VfwHERYCT
KbinwJEmHDPkkvhDpEMLSFWi6gp861bCcIE6i8ID69bYb9dd2W6khA1tG1t1tAmB
b4y2tXIz0QRRTg7zzyjdUY8XoSvzcmclWNYfTlgxfv2NX1v8qVs2syy+/6A2cqqG
DVoV4RNLrmxoqSI8z/WsaAwAsK+0S0HGoDkRkiPZmCk7xd2WinX4ITqNfn5U2hme
kn76G9F70/BjGEGeHrAevzsFivQU6XqwsbBk+iz272OogHzq36MYzx4QVdhEuRd8
B2Ka6kqODuDK7kqKi4TggeRv/ATHXzHbpS+IhKd4yzrdaAPJjeSe9KlRb9FycD1E
C2sE3yNrgRqLSDQuBp0CzCcFLHDgmLVogFC0CBGEcfOxAhWC4X93MoBG5c96rpeW
9cs73c8E9J6GFFoeSVV6aCc3hKdX6DcfTRLlgNOYI0oyWWSM1LUI1uMCaQamq1Ly
G1d9TigQ1ruq7Ydu5V4jejRD3lsMTXxphgohFlOvHVdjjzRyEWOFBSzRTCCr60eh
tkfVHAhHbZxBFRq7eGomA+A7aFPFDhjFH8ezSj46gvKJFPavMTx1h+uaLViISDDw
wuJQNQt/kKh3jRbhAhArQaTuS5VSfuxx/1u92TNuXEJc7mp5ctbLWMG7niuzRg+F
30oLUXT5in/puVR79lOoXtnW9EZP9pcQB+d4SNPep+i3SWWmCxZT2G+twStE8g1R
eQziQ7I2B9wUgTWWW95/qZwLy9iqGSxrzhGWRJswMAxE+5+BcsRPgYNttFFRtD4z
znb9JKkBcu6rIYvNNMEnOnCDJHkeulAlYQdTeKeezMRoK/H652xgdhfyH2wDWWYg
GFYuHlISIIS2tyf4jRxNgwGEvh6601O0MyowVwlgnvcNvEw9uPtquCrTlWJJ/BSB
Af2jsFDzGF3ATqYdp69Don6l/1ngRWdBm1KIhiNwWumby7Ty0VekO4Z2Dq4WBvdQ
dxaVnqKl76krvUw2Ekoz/SObbiEkjdRXU7e7C11iAQMEp4pQ8wN2dLYzl1veVpqL
WmzdtpkNIg5mtcm2AoQpZsl3b0QAEeLtCLW5M0R3kA9RCuKNKd230brxu42MUXdW
gF3SxnL8jX9LGIYOdey0n5DAmZ43kr2EkDODe5gcHtvbjvxiwmERsjs0pvkM/a1I
Jjgu6Ya1u5RQugf64Scgs6vVmtliQ8VlGhqlWejEKIkwldkh8nmGNEoPKpNFi2Hd
5zpBVeMFJBMYqsAU4EoefhqYdbyUVr3+krc9S+LohEIfOzfNdCfMNCDac1ovZzEM
ZovuFpNnSsHgiwJfFf6O0fk0sGtLnyvUNn9HflTflkWQyEq9O0opPCGyREzeHR9Z
1e4IJg17NhPe0LiVedI0p9xPFYuATnIRkg+ClvpMM7anEr7LBfcAoNi9ym62RHCJ
58ua9IM5Z3W/0rTpnt1vCVZTs3rVv2VnzRX/tPNuXAWMgbABobQz2lcY6ft5pCx2
o/Ha2dXrTS/0mzl89BR080zWp7yqo9iKgppQxijqqna3xQD3H4Bhj3RLh8RkDgux
kyK9ilgvgirinCZProaHrQ5M2GXHF4x/IbSoyXTIL4ybqy2g5T/8x/adNTvCtBw4
H+XRsmCSu94pvFRBHIy/vH/2gVeYSnFjGn9vYOGuT+d0xk537unaOWqFFo2bCe/+
6V7lSHFl1n1aMPMQrojB1baTGwwEjUnNgDm7NYi3uVROWqW8R50aMT5SITjw+APQ
dx725XWit5sz8gnhOW/ECZ2MDow7CeB6btEaCfUBHcFLe8ZPhYmuaMsUdzqOv6Pn
ET1PM5w5b3W7R9BJYs1rYpOHFmdHiZPLrNEHeZAkIfTJQUZQ2iDtUyu+oBMOadqC
UQsqJuoIdQbiKevHjzrkUEllcPkatdFDdP/oazZUK75R9cgHEqUlSosgWpWfZ4bE
b7frd80uR2yLsmFk3X0vZdLg9ew0sbucbYsZbUklawkCtmPA7uRA2xTDG11bWhJm
WrsnFNWZFSEe+TU9DWkqfszzm7tE4+HOkKgB5Kuzs7M3eMQxwj1oSEDJf8l3IV+n
zXAV1k2/v7XtHHX4qwoufEdQ34JhLA1ZsK+16SoCghvzmYeedxV8RMznCcxm5H4n
l7AIdjo9nGlb6cjCQAsbyjlMfKbQWMNA26IL8fjF0SZnSZ4b2pQeOFgU8YtA7qJR
MZlusKQ2zRspLh1RPbYpyvYcU6bnUVR5gES7vP5qqXN0+mYvx7mXwvupe0mEOhoi
BDRgRlY/E70h8lutgMFVhbaqLHQE5CBvuugKb33eDyxGBlBbtY83yiU2e2xH5WZ3
8EaOBLCIcNQMvrp0pZLYn7OyPceuclLxygQmg/AwxJhvr9qCxkoRuiSAnVfNOCms
KvS+BHBDrp0ud/xCK/cDYv4nbrzePhMeORsNylZWbThwJSmRIaittiDTKnmfhPV1
hWkEpt4UW5j6D/dnGBonPCpubF9zFGvlxVdd/MbOI4/pdK6n9u7zoJXbsCLI+ZTw
RIy/4SGMEXvt6MRcFvkkOMFdZg1ZFC3Q4Nbc95B5k3jIzLqkBv9sb48nXZ/L9+dm
PDsK2GLN58ZBp5Z8YGQS/u7uwYdZDBbMMI3U4KAstPeJiSJ2gqZ6Ff0DtjGEGZRx
heLj/GcXmt1QUZwW43lnQYjrrJ4unPK3qjTETTER5hIRfBWROMLarHtd2P96cyf1
axVwwq+vYhTuJMT8NuiSsDsxiMgW2z7D7NjJSUSJEErD3MjYzC8l3jt9XbPmBsFe
A4iAiCGwnCf13zzh62Ei+cqqTChD1U+fX7Mr3gAajMgigEkVA9HFD/T7NDWt6Trk
xP7MjAhB1ouZEEakjv47tyetXxhXg713hWtEW933XQFnrsWeX2UDZ7TPqj73nh4f
EnLZibSNRcHl6UdX38px04BpwPjjf96jcPJkydo1cv33a1rfnSejnEUWdKGUmtQi
UH2Svjtj4N2gwbVPfovXSo1W5KR4SB0dmJ0Ine2ivDzisH5HyDOhA9bmDpt/fmou
9L35AUAGDTMEZpdqWVAPA5v47Dp16Ew2n3ey17CwJZcVrIRN0TDX4J6xtaWT899R
jgNdRvC9teQLQkQeiBopAak2U0yg+arPr6ve/BKc+MSSJw3p0mettKAJev1Ql8ny
bQF6JWaR+aBiUliKucKnmFRf7iH+lCp0Y1L2SEDnAgmj9WuN8y/+gmUh/xdm9XpH
4Rhag1F10lFBoxfadHTEnaYDawd8yFdKp0UySFICoBv5nx6ZObOckXYv6btEoWD0
cZPSWrDpm2wqpsVSfDHQFZhjPU9scXZLJQxIlsQXzfwHQ4EmZXXsMG31Jl9Je+4z
IEDbHbK7fakSMTg5glg6fXseiuDk26+dgzrxm3KkNMggZfuqBIrxxXLXAUA2RS5n
Qfeqvn8r00Ph8s49C/sr9uSa7moFSVMp6q2SwJC6L0rcsdI18ruow2yHR4+eCDEc
Mx4qyA6rEiua17nK7a3I53QSl/EbatzJwTBGe7W2pPzgWYCRSy3YszCLh1FU22ea
9kzCBXF7P2304sDtHuuGct0X0mxeYtAJhYxE/et8zRS860w33K+1x3VSH2xfh49Q
047mlCWVj2kqLjDIbK0UyTCNuXtC2/RgdRbMiRSybTKx/zqVgPNOPPFnmTXiDvZl
k9E2EwL3s5zxX+/QqLGfPy5KQIvII79m/yvlta0tx/mhb4C0NZOzGvht4dftCjJK
KVzJGl70UxCQpAOW7qkcVRz/I6/tyzwzkP727mrsKnb+m8TnvGktQgbI+UvFDixi
nJSttNO34O7sQrfSE3JWj1mGfQmG4qKABp8MaRttNoFY4QoQUFVA3aTamQDkU/ZC
oXehkkRSdZcy7rOkm6w/9h0c4i9YjrvVmIAJF0yMwGexy+P6jebDXD1gdxk3RLEl
yS3llu7MGiZAFL3NNKPkggMmGpCE6DA6EkZ2KjLYDxzwGLiq2LQy6xvy80+f7x1q
a5hXzIWlfzDV3znfz1Y6DjOGlGKByBt8EnaSUSrmD4crLKp369h7/DvsUYqN9/ut
U9VgyIkd6HM6ODllkBA17xeIYvbPsArpwbeFeOGIxuaNHQmunyRyjIiyej2q1Eqx
WJG8HN8VhPFkgvc5n8OGeV1BukQLHcDaakoJR+iae3nmaR4pk0tFqZdBx0sbg+v6
00x/CdhaKzrX6dp2HJ9k/NsRFyx2j6UmcwMr/4H+TutBNRyjq1focN+nMuknl9kJ
2CJFBZVMfrnwse0RAFWzuCjTKaBRhLkEMajEp+X0pRwVrvQNeDIjALv6WrhMh/BB
XPQG7NulpjKa+nSf9+E2He3jCWK97Q1fiiQT7pzX79E6M6cw3EwNLejshSFqVXID
10dPCJvGvzytnBM+pZAeltKjtsS+8SJufWa9DAUQIvGXIiegfL79C6ADd/dTFE0g
4+9OD/x1vVv00FsTYtuRS0BYHdoZ2n0hlRMFK7jF7H9axVZbd3bi8PJr5mSarV3i
Ded/lkFVk9UT5pLKA/GqoucxlpZ4SLOPQkV6askuXQHKD7+sSVsdmZ07aTsyb1Gr
B+ftrYWL+yQJMrmWUQWIewdN79Ytg1wduO61kgguY/gx899Jw+poeQwNXliluzZE
VI9FiklkcRFn79oPsGnNmSWFMP7P2gGs7OS/aBu4Vf28Cqa7juG14KwQWtbgrTGo
oXnyRuQ0Ln1Z1Z5MjYYIq2/vLWnjg9Z66DfbhYsadzlbbw7HTICCrVu25fwV/g65
QUBrlTLYZrWbE54qTJdTc0Nu1jVQhA7hb8nvclf7Oyw8cO/1uO8yAQ1t1D+VUyu6
cNVC/MBtDDARP+5zRxfBNjy256XKsWJV+ccIIvTj8/AkRsALW7fAw+WxLdMLB0vQ
phtt+EGPES7z8p8m6b9CZpNKl+zdfOoRYI8fznk5yrBXqbjJERV0mwK6XjRUMa2L
IwM00oRUmlJEeBoKibe5NFHoUvwpjB/HOfCXA5oLqSxItKwhF3SnXyoOl2novGxu
ZvotO+E1BMG71akgtI6X/viQXBZoq5sSRFeoK6A41soL9jMDI81W1RS0sVcGOTDE
VuLU6AbHz/htyRwasK0VK0NmIXKbhG0v1/Whh8B6AYkaCSIRxSA5Lyj+OVOy3V6a
FQDJ+4d5DsSWvTia32eYd6jYe+95BGQvpWmMTAvqSwiLdWgNmScM7QHSbLpzcOX3
s/y52NfQjL5KsZbWEN49cgk8yDPifQEuHzHVy5l3wMrcnEnIlfvJTKZOxw6URNha
XazGkU3ZWuvqYtB0jp23hII9AE4HKILd7tL/fVoeaU6LMoV9jjuhNZZ9Y+OjyvLE
kfiXfp++ZnLRgNEb1Ap1rtAPjh3kUg/JaW/4oNsV2qtums5Yb3l67+sHWYt6pqGW
DR70+EBhcjMKS8GKq99aju2QzSk1x67FV1rGCvhiRv2P09ju4Z6UvNPCdM2EmEJF
GR+ko8cadnYztrXT6gfWflPD4bLq53ziY1SXMuARoqFu4fA0tCjgvwEbijua/c89
DYcGCWdw8qETIpw6pdeeWCrJ8UDzQtwKEuTcl7wac6KNG2Q1QugAXsFzZWKrASbx
ad9nQ16Pnd3ZUT5myRU0r66GfFarcprxTQ0P5wBwMjltCrQ92KYHwKqClJjOkXGy
cdCmru5FgdXpQLUDIIamTCTo4WanJl7kswXvI+V4n81zGsppYf+IkDMZOUusjYKe
oOq0U8v+SyuW7Paz0GmqqTBpHv6eygOOrgJA4frtxz4PoIA1ErmyszuYCRg2223b
sOGzEC6h7hQFCB97zcAGVJOTygLNaVPvJJ9TEgnmT5k3GvZWTf8kEg6lQ8OQLqvS
xl8bKibi0go5xcy/UCSjATx5tu+JOVXaBDVcIcg5u2Woy8ELSbCUzG4IyebZHmkU
gBzio93JnlhLYP0gosaLKlC2X59cQPZpXObb58WG1jbPACHJg32WjNP7bkIhKfqG
+Cjw80XkdpYLuLuWTTyLFSzi3EWIfW0VtoCGJ+hxBsDs9ou8Rz6yXSNwo4tOjtie
+Zd8CW+gTpPOidnc3OT2qqZeWGcE9gHJaLBEnXAxpNC3oqebNzviU3FrVekQg2Kz
MvO1EvE8eQyhEiwZwak57uAsqj7AGNbPF/LQxXMLxIMyIsb6xQxD6hHoXHgf8QcI
5rRZ+ATidyF9Qms6xV+eeoq23yvLsZ/KJ/AUzapjtuujJ59wY/gdzajxTwz6shkd
whKwRyhx/VVJMLLyVHe5zUD78bsPVxlZXWzMUFX0fLI4zdbpYj1RPN9a/lsD5J4g
60RlbJ7aQ8ZYkdFbQXv1PBxs7GJ6jp+Vh6XOiO5KWM0L27yq94D94XMk0EiXHgmN
Lg0rQKnu0nnrkxsSr7gA6pyzvtkIRmsUtVZ6w2qSY5HrmcPS53nYV8mO/m2Q0I64
nHqX9NiuVmJGZHtqTnEG/KR1t40Du9wskkCbyVTNHFt+aeLlLuAPFPp0ky7M/7Tv
8zIMEr1dPEFgMr2Ydq341x2umOSTTso9OrSi8WaQ3G1yjHBuIcWGTXKqwT9KHcA1
YTIU9WdsIAW2RbnQeGxabR6OtrSFBgokDRPCicYwAq1wdBUJtlHodG4urXTlKzjV
x6fJ4lxNXUtQX04U/HhvGEzu7NJiUCA9xf2Hbbf1abcSkm2+cqJsuRZa2fpfBH37
USzXciL5c1XAe3Sq6K9dpvzBLjKseqb4ih8+O/HWWjg0q9igr+okBj5fkbBygVvO
xz8eRp5cyzsRuoE8CHWYT3qms9dCMGTgcUEOTEVzaceF1XnhFg8/1lcLHS7t5QwE
9xV9ReuZYsSn24sVuwBc2bzFZqQwMsOcVpLNFlxR1vfpvGNYfgwzAUAQvqsg1ZdL
hg1WJD+cmvzkIVEgwbz9WG6eKjdKIq35kxaXOoIH/ZVmrqMOwTRTmavFI+Z42ihr
Z0o7naHMV8FyhbELUP9XxKz7rkAVrFnihmn3GfcFLcWWA3e/rhf5wzXHE2gYDWJq
Iu+vySYOot97+JVxcENRpjOyt0ZtQkqLauHyghjOca28kelJnct3aveX1JcqqufR
/oRz8Tmq23SFArKtDjAGyGRwMEZEk+j8+DaQqCi8/yAvfl9CunjAZxVH59ytamMb
D+evP7jYK5r0pyMZmM5CPkG4B1DNzfCeWdNxBNxYEwxct0FR+rBu93IMV3CNDZ9F
PMvBxucFSU08B7ZPKcrpYQzaJLyElQk1Qv74Einwi4CVvjAVfCo2/F4m4+cmZUFy
K0Mmqf/ECsTon34UaftzoTtAHmycJ2cSaj7Ci+xaXOPizRMWBuZop5ZjejIwUJNB
otxOJ14QQxRlHAUQqk6RBaBVz3sCDxD2/f8Q3FbZP1PRVyd0B5XeyyOaC5bCY3aG
qfk+qH3Xa8GrL+RxE/br3e3mQSBZkemu+dAEiTLQTYUDj9z/i1rg4tS8Sy94uYm8
CVnsyeGI+eDZSkCXlVXkORCyKEaaSpqpno4VPV200twy4qLTzrnHLCdyzKeGi/j2
z9vBE9HSnnW3GLmyKC7E77npT2xeXoImrTd36ESl7ke8c/HJ/ItPx6zShmp46jGf
rvQOM3rpwU1xGvxmjQvFISjnme9dAgGqBeAdLxkd69BMCrvOLEd2JWUzabqun9ey
uTEhNhnA/32SsS8CFziKDNz62ds7C6ImLXJRIgfZDA7kiwVc9CAKxDKHpQy+g4eQ
U30j2+CZrY3UMeon6NIHmQZ2Tjj/LZSd2l8tv3gUCaA2QBTNNDGs041XDfuH5zty
LDIpdRFPuNzPcclwHUHu5LQJX8GHU00zpcZ+Fp4/LeUh01IDf/SYnjaa0Vhbv9hN
79V++DP/l9nPrCbxE+h814B0Nm2y728Ae6ZmLcUGljvb4v83/QiS2ekwVtUd6PIC
Vit/QE/dNZJvTIPUnrdkWyeLvLJ07dHUa9NP5+di5f6xTHmjWi/B21q/4rp8aFDg
d4cFhBf3PVSlwHEJ3xmtYTZ9EV7ezntz474rRqentqR2d+1NMp9lY7PQtLp0Pwm6
4sc5m3Bx6NDmR9sDTxLBEF6Gbm4Fhn6aQ77RbRSwrf/BDK4pokZrZ4+g3UEvXt1H
cAEwBBQoP1KrJBQYf3aL/iwnqy96IB8Hf6eDCaaFLzk414mFmdVkGrX+YM0JqxQO
SqNXeIkRHGs+8HvPDYaj5eZIC/eO1ysqCC8PgxTgnW6sjxuN6BhZMe3xXdtjfboA
w0fKKXqr0o1xhIXBi273TCP7yd1wz5pYLDrhnrspltYSJ25jNOTHaK7TqSMILYu+
6/U0OlX55+sU2uWLAWRIIfo/OI1ERLwhB6XSPFObOKu+Unanl/2Wh0CHFW9Cy5UM
bx80QXGqUfVgIotjeO37LDyGdpZ/DEADI426VOI88Mkr7koLuU97wqMZ7N+GuwxZ
RTGuz5au+/dt/Bmzpe0uN9v7EYG3p5iEzSX8Lq+8ADDYHcBTsRtg116o5WmbTiXQ
iY4+rTtvQr8tT2ERNz+oeXH6qSg3XGyLI03gX4RlWwAQJckd2uuapSXYiQItaPlV
LqquMRGNpc8mFn6qyeKNrzNahSAsFns8/xOYHwONLfgt5fhnUroeqjTIUkZHYdH+
BAvGVeGcOGVV8Lu+sl1h2ZfdLtigSiBJ/M0H5TtPa54L72wrQKD67I46VuNG2WWh
v/LUVg3y5XGqB6WEEpV16sHdXD7JK8ViLuJU7E5Qete3kRnWNjnDItRnY7eNXNNL
S7tl8HHU3lTvAOmAzIobto9TSN9BLD34t2nz9TIoMUyXk/Rlq+nNUrw5LCAPp2Gi
9rL+341E5krJg+5mhYUPELiUCZPzBRCdmbfiCX0eAh60BJDTjX6P+Tz/rWjJM465
6O0bEtR1SbjFqQVd9mdtHWsgucaShU66HpzgUPuHtC+84jEeGEjJoMAGN0eqESUN
LTK97gRDWQPK1GJlwthoD7H5Xjg5VdpdAXambx4n6Bl7CUy/vaJqaUiNvVK68IQ6
gxn5X1wPydHWNQ5CeWM5YigiJX4ASJsxaohisZBw8r7JMYU7lDrCz41njqhSt19Y
YSOMzj54OXHXJgHEElEtP6xAnFfyKy9qjlTm/BDjknLuaptLfravmm5ewQm6M0zx
7RR2MXgqJpm8gZsLwYuv69mI/zAExBGAnACeqscbyTau9OdSMmCGokk94zX6t/zE
cAV+kMVCO2l+kw7HZiqir3FpLqYwCXhiAzwjC1PtaTH9luxWEO6RXBEawW3UmR3i
agoFsOCsVewT6WuQGzIjHGOPmrO6w0FIXsZKkYIuBRTlYG7x4zCZLakkwlt6OzNA
bKqwsDYHBbEP4OKNXtNxi6Ekbhnj5ahZUevDWIrXDViNtZOWsr0SIICck/6kDHEW
1UY/I9+zCI77oIr6QB3WpTlWz93wLu7HbctpmDsTUdc0uODfLBilg/h0x3y14FBi
9xTXgjaGKW91avnHNvTjN+OZInyMdYznlVnhpo9LTy4binjh//k7p5Rw1/Dsb6n9
hZWhnupHgarJvlJfuDF6vs4CrQdnL8P5QLJZQ/58WBHyr/vRsYkVy2VkFde+ue2d
8/dtVbJJ744G82RLrx3/m2mk5XUQaZ26FeJdyOS/BBhoUECNMipytYReorNM1E/e
GMBQ8GCEjUOVDLR85d/ef0SrTGH1NJJiJJP04KLOpELJgsat8mz31QZxIUW3EDX5
m8euVcwGaQpDxeMFMNW0gIYbAbzDrAI84c0urIdmcej0taF8mwRNhx4jVuqps45Y
dewXSBqqHVFyPKps44bOH61dmSztHxCLj/kcyfameskuH4a9OrS8IstbHgNEKoC6
fbXladA1JOrs5S86C5A2qRBl2FSLbnqtsRGjSS+cTg//4HkyZaMun1R+9FPaQeHO
2/1ekizdPt4TwkwqGvYNUR5RcJVjC8KRK7t4j2o6irg/peXnDVXvLvt/e6PopEs5
4MHLgHGjPZu5lffn4wzpVJbRCrFJAOdrXflefT+UWCQ6FhWo5i2mtKKG5dk66X1W
3Nfgz7HUlMU2ysDeV20VBlnn1SNpRLcm0WN4WV426oONoYZy3gZ4Op/jfUVWSvW0
29yU6VN++j6NPNvz4IBMzmNLRBOBSJnXk55HwR1i1OlJW/1iOcaUvMpvk+jLZIYk
z8Kllre47erQzYS0gqM8Ru8vDvIDdhBuDzXr9DDLU8Af96tO1z77F/wc3GQbv7Ff
VeSLOcGVQcNoJ/ImblayRFtHIRYbOHrRhIFkNmGRXs8qcrqmtBc8S3aV1dHttAth
oWs4mJED+dcodDInCpri3z7LiWYzVHNkC5dCR3aFQQK18sgal4i15KHKxECjs9pB
deJb0zj1ZFpDdo3Hpg6DrC2osvT7NW9qe0IgwnqnOo4NA//XRUg580QFxbPYa3Sz
LnZl4qs5UvSKLgRCPA93vd05qBA/zu+JF3LA20a6MAqLMpa1bORaFOoN6JuAqGa2
U9JnjHWZmH4ysCO5n9tTwfWPt7bQLSrQiUQdhX4PWpU0ZpAFDV59P1CvwRGPnhFI
6wkBeZ41ygZX1heaTTZYk2WpF5VZteLN5rx+FndoR+6BU8Ww+2N0AIzP0CL9N4U+
jJOxGeJ9mx19MoagBt0iOKPZqmkB8eT1oZgVA/bul18easf3uhfyVuuRsYx/ZgRa
LAfR3j0B82wypvCMCxIPv95j62cRWG9iMHOsfJcmiyjMlBS/H0yRZ1pZkW0JfyGo
ZH8jFX3HoX938r1/Utu+w5oUrAJGGJk+8zYTUYo10rGs2DUY77V6okqFmMm84Tya
z+mdowfgab5ebZBZ51VvlVkqm0grdLrMIpzmZfS2jaZOUOX1X5CSydQFxIsG7SdX
6VWjMB9iuX9K3bDXIHpHOPniTIrUPC3+ErBjjA+3JVUgyrcqwDCyHAMFkeKPNiKB
MGN/qQ4swgM0Cz4C+BWEHc+0djNGK13aZCQMds2ziSYw+92FysQ+4hVv6m7klaDw
W+cL71aQ/2S4dgSFoVGf6E9Yj1JLssPIRLGeoXAY56c3vlPaUg/BmBHphrmjjygU
MunUhnIVGeiyyUhDdx564nHiEH34uZYSGpY283Q6Ld4RPw6Mwcqk0OBBLrQy7TqY
KDw+ruOORTkw67m1uLk8lCgZ5FQwDwLFp7GP3wFff3/8bWtoHzlD/Ht0Nb7pKvci
qnmAY0PMkhH3oudmIjQpX3dVSKMlRu2wC9Oe8q1j5o4E7TcLGYfjMp6EzGKp8qzw
Mc34PfmF1lUyb6IFLa6BERgDwMLY2dDaa18FZ9rXFMYdC3Y94Xx17KEf23WIHrgn
jjB9DvNVtdL9JNnb+s5KBUK8X2IEZ8yisPb9PRnY6uQukiq1avZqtG+jQLXE+/jt
AJN0yU8SjMlfwu66DWcaKvC0vJBgxVk9DPqvf9q4CpvKMHcF8vlnPjjfY6nKgq2u
01EEtt7e2P5/5u8l7cvs5Gga+KeHJZxV4/5dzd12APU52os2HrZHbsfjG5HOEjl1
y17/B+fQfNFM8DcCV8u9DLYKXdVhn+LrOjUNv2WmAXo9+jMGOfAjWNMEYDTmFf5J
/0haSVvr1EXLGSqi2yLD4nZRjin4ifbhuinUO3t7qCZCkWgcLLi0c4HdQwS0JpQW
KLJ+n4tAdi/Nni7YtJuW1F6IC3XGEqiuts/AjThmduFq7Z13QirgYMmgNCgDDxnn
55ubbU8VFfdCiVdQfEbm0dPvKn+SP1svUH+UAbKl19ygtICs+GplAPnNwIcMfDJI
mzzfZZ39mMIbLbXtX3MGNg36jllsgx6n0uSc96y3mge+jT1xnUfFfxd0sQ+uVKkh
XMC8+lG65rweQHuHjdrxGZvq8YbC4IY3wIrf4I+hWJ2jJdkxSFt7VQJVKSB7FxtS
obhsZdoSX2VOlG35xQPG0sCgCxWFojmYCD24PfC20r5c8JjZo8G2t4g95ge8s1ao
/HsDinoGn67J18jEi9z4OnU19kKCZqKut7B88WCrVSH+5akgj3jELYX1BVOEWXKX
DmjnIXgVaiwP4jTyaTYFLtzuE5Y6qy050ks2LXtbNeTEh+Zhe3/OauRUVXvo5x6x
7b0HyX4+iSm2C1GbodP+vJ26QAt3LY9oi7M+QcpNodempSaSGlUC+XhN70kTjxHW
P/QG891q6ea+2LNONqHDRoiyaYbJ3/TZbj7fi5savJ1pKK82spOHn3x0YucWb82l
5ntvwwIzWh0JnEy4uVN2OiD5165nGOMQ0JPX6UkDOexZZYSWwfyJBFOC/hSc8mNQ
sWZJXt4bXIa/Zr5ssCXLNPOTYAo+Uf8A5BaVN4n5qo9rRG+CmZyN5826/Fp0ERf0
uPqeDEgwgqsg5QBcT7YLPExzk0QkDwj2nh2zOIyuC/Ypf6uwauFO53ezRrS0/E/C
scacyTccTXVnlwaKy8klc5GvNA/f0As1yKKCEOUvqt0zN9UsdxWct3tjZl46rEBe
meqL/BRxbp/dtzbPdpggASooS2Rf1pqiBxByMkXLkOCOr9bXIQq435LPiGA0AZAT
j90HUcDU6yZAYSGq+d2j8n/AtlzJjb7zYT3tw+k1Iua/SCjIrFnGGJpu9Cr0D9oW
beL+j5ay5qkYWgdjR3GuwMh8QfoYXM4UljWNXVWBZ5AAY4W4ZKMFVj+WDszZc8Av
UT2NDtzBfrXPLfhpTjInCbIr6Q5ZL/kKuZW+I97BQtol57mO6F6fHAjpN1N9DCvh
+74tWb2m/3RVeG2k96UCt3qhffjyo35f/8yAGRxqryv+j0OUbaYctBqST/B7sS+9
iVxJzlL9Y9Y8QDndrtK5g2CRHb2ml5rtk/aFu/Xip8TerLLOdX0n6AGFtqpIeazc
Jj9ZSZ796OuqSBpQCSIxCw/dY2FsQIrjWV+IVbgJg7i2V6SjyIYHJ1MixcIn94ph
MAVb282diEG2Ol0jm93au0jtF8g46HPltqQLjBX4SUzzGBbl86UNbueEgQWEzSve
xQ7am77BKWqYUuKVyDYyllsyKAQM2h8QmoNoY16h3QGMcPu5Lsegiw+k5/IZr9mP
BGY9kyDLLPaoj+LmjHXKZeaYR2XJ0PCvq6zfJzMjJrxT8RPMlISyA+LOJBjPbf9f
hSREjbe6DFv5UY6OBnuKaRv09ak7Ld08/hxY/jZOgvrf7KbRDfjMsl46fhmoCfAL
Ij1onF1Ru2UWZE2aqYFlcio3Q2GTcK2FJc30Dn8F6xkZp5je/9eAoS71D20v9DqM
GvQwjuUaebNsTGiNk+VcQtlG3NOLnyiSx1Fi/fZO4LB36p+S31FeEseBcHo/qJw5
mU1XPuk3egDQbZ5P/boFlAj9nue1F/epV9TPfRcwV20x1/WcbLkN7lzKo5Ic8/Z0
/kYhGtT8k5Wb5DhMxXPyGXvwfjNjpp6yW6vJS5KS1cgY+1clbWR8P4Ny7Iov+WBU
yWYtplJJVn7DAco6aVdSmpXKrbSL5XqgcDTQK5+JeTYeykdwzX1Fo0dSHc/B4WU3
tPCzFkNBW3BPtBBzEf83ayzAgom0BjmQCea0Oh1SEwT7sL38cajgfxZRhuJPhI+1
sPYU5Vx4+g6dH+5QSlUcI/2DZw5WN5DPjEyFC7RxSYXcWfvTI8mT9ko/oz5K9X/h
OHSLCFeZhB3MtIq5E4sF8t0xAYxORzpfgd49op/uY5uZFfB3e2QaCWfKEnxTJ7BG
Qu/EM+EoA/k9VrPsiGl71lgNDJKwwpfvqNkzi+JHQ4hTA7QunroqgvBPKqdrb3Gs
PGyXiLuN0bOB5s9VgiWXqVV/UXay+CFcUzlSq+zBxTkMoz9BR2WUjs2Us1x+II6K
xjROJTovrTiexcTzMxZdxisGMTyDvBqojyD6fz4amt9/Qtio3KaNt2fK4jPzm6D+
Fill7WqLSqr6zSJuQ8u2A3JvjUbEeJ3JkLZpk6tXWCq0V+OVyIEr+zED98XTC1Nd
v1yVPHIbMzZkKEEZ5P50rULCmbxRwPQJMG3xvjYd+HO8Kl8bpGag+jxDDxTawTQM
3+EmmgU6gDpjr2Tyiw/lrtv/dFha2u92wdb7gaNptXBvVpDMkrHAmhUdLkbwIpBn
ve2sjuW8pjMpQIxUuj9vCmzpkAP6sfxPjoC9/aSRK+epHX0nwIzmBcGjQrHHN8ZT
nbSiih9HCEwvIK3n+ckDw2D5Z3BtvmOCKwk5sBmcypzmd1cRkP93s+yw2kSWLAv4
qXQslGFU161UzJfl0mMdL/UJngL7dVIphSiGBbvIJaRfIEJuY1yDhURtDtma2dCQ
eVWvgw0A7gHcb2LsxGM35I/xD4+M4/XHQZOvom10pI/IgyixOZXK9skABK3kUp6E
x9C0aa/TiULUzTQUTQBoPHqltAhnUG7jRzVvT/CJtHLBmIEeBvVK1nlsjnQQvsTG
zklZ6t1YlR6XJfPG1UFlYAoL1Kwsz8tRXlaU0Rn6uwMdyOrJW1X2977+sv1yT1RC
hUKYP4/DZ/1DV8Ye4o6UoIScm+ZxQamj0MYAmXjPCED5P8/+OC6/5PaYcDanOtAl
ZPzIB/PuxMzVQhBIkFNaej/sYBoKGe68RDKXCO1SAfJFVDDbZCjWsRZ0/EZ7aq8j
SVHNIibjXAJlAFUyhXzOeaTR/fYusz1Q9wJnDhH4dLzYqXDryBgcIoRBt357U8mB
4rvM40DEd+ICyV1wd1acNKTCrObbbGMdnyBLAIkJQZWcMjlVRYHSi6FYskzJLF5m
wfBKPK0VMeEeTUGnb8XW4oMpFXbst0b0xmbjIcCWJsBXBpmenzDYbbSEyGxvHsyY
7uIirxVWUcl9mCWCBTof+QZPq+jDSi4JM7ZDK1F+A4QotSqLSXjhP5gyaEPEVqbE
Njd1Ol2yNEXRE//uhTkle7HEodEprVbpEqqUIMri3VS4hoe5cUDfGyWXwBwmewA+
tRu2VwiEGDg4IQBPLTenJxpn+jPES9LJfBIN51gkm1DuRGnToM6iA6HfgD/rcOtw
NJ1wEK2rwuY+QxmC+R0q9BTMlHASdB40PK32+dPSk43+Qwafcgqseuh6lrwlolyP
BCMo80h+pktVWzpKd0u72Ttp7K/Tg+laaRp4OuGHItxw9Ktynr+TE/C110EdBmKu
xJ9pyVQHAuWiaWaf2aL/QNuco5zUJC4ebsVytFVmnIuekAiujBfER2eUMFdk14Ni
UWa5URWDx0s4RgvrJYY2RqLe94VsCmaHTG+5+ohwS2n8jR/OlHPHRX6gS0AtlyoD
FrW2QJWv3fwbih/PWZtKBHuv4TWehgK2BYnzL1nObM9Z9H4dkHWe3UpPCp686XM0
e2XERIaLjAHF9Ez3c5ipbJAX0vuE+GeH2HlU2K6fXWIBKANgBfASy/eXXdBQf7Ce
2xjk0iKv2lDRhVDVY9xY4itugHI7otNEAW49h2fP3UgNox7rN77Oia3qILJJZKMs
4WUiGR/I82mq9jYTc+arvwxVoYuOS4w9dMFWNPOpL2Bv4EzZDVPpnUPHYd2aiWjx
uDBCq1x9IfeGjfbePZnNgF3IjNMnRWzoUio0LipAKAvFvdNF71zsN3UuZJ0/ILgV
OizmEp1oi4avfmkCBKgOdl/tvB7LZJTLyJKPCQSFN+l3i2LMNIZd4JeW/X1M4ikh
nOhD1NsMMB35YyCQA9pPH0Mfa+y25fcH+XMfscQ7x7Ao365owyoxgMKSqRNGQEoX
NyDxhjdPdwFn9+36cOu9A4pkzRCQeELYYZoo0yKfDGuco6Z3MFnoVXm5G3Ls0FId
rTpwq8h/eq0NLzYXZNc16cKDrR7UaYSdeAmrWTFWrkIvxr65ivtNRQNV7Qhla9gu
pUezLmWyr+7Zz8++V8/I53AhoW8YDuIivR5V/Srf3MTc9hTjEZVfAd6MtAAZLru8
Xz7L+sezuyIoWgteKhgVy072Hkz63phj0RQhdq8RQbXNr04BENi5IS9DJ/3FpLE3
2pKcmNkDfBUTjcfD81hQnJ1HVYSWjoUwNuFbU4zKw5SB9061Xvq2sy7GnrhtC4Hu
T+Yr4xpdNOYS4kO04vpCCP+LhADu5KnAwh819ijQkJPc+/rwHMrScGYJQWPn1nQk
I9Ijjabeoilla2BV+i/hBOMx7kXy54MO80BDnjcqfMq2EmdMNNuSTq0bHnNUKRFp
CTAZ7eLjaETp9CIeUPAlEWWybIP7p+TeYodGeT+D+FtA3mVmwxeNnkvd2AYy3ccd
oLVUkvf0u+O0G1mOwwh0ZM6fXssVv1g0C+5yC9YKnSCETSLq8zXOGhXzmiOyvNrx
MjYBJ7fF1FuBILdr+nT9mS6BPogMp0k2gGthHly3vB4jQdQYsU2YrMfjWPnTQvo5
9cJ8HO5I/59YPpmyrTq/KOkXnHuNtVIL25shr6zZluIgcbaUry+ppxhS8TgqF6ty
4D/uPWD7DeOI9Z/uvq5KTqREwqUQqiGGV1ita+o3FE6z4FDDnognBko2Y4wFIPZO
ZXpGwkfnbT213yIDIv8MaSREPVu1w9JkvxgdaMo9fOzCQhKXBR1L4iFpR4HRUIDc
gmYC2tB/bOgRvGx8fFeesMn5cY2+c5IeCZefhnTB6iyUek4GBiNiw2Jc5j8xTvRz
lMcpyFcxFnixcsqCw+Ll5GWj50jFOIy383VNqEBQPUAPAiVvoSpJZHkZnYUp73Xi
XB20DSsTCp27a3vBs4S9E735WDZZp1zIfE43wtFPDCs8/TSKoaUb2AoZwmJPM76o
ztzqDmtZEBT1MZTu5a3Z1B2Lq1olTbpE4N2eh//lKPU8cRGL1iizmQrQrRSFh6mP
L9+nXUC1GaDcXx2rcLam0q3ftzv5ezO/zZg4sO4dIbOCsS8j/UhLurH65UrFvij+
Bfh4q6fWnqKJC2Vp+fIGZeaic6wEdFFOUGu3lVy5vNWgiuTkH4nHwfY4Fv+ySbkC
HObMVfLfKkRGzECiKhh9HVsTjC2t/RpGuGx+yTECzG5HA8/1keUikwr09NgQLprf
XSw8lTbehNFlvXV1ugCpWxPSrYw/MlH3rIKa0xIswtHcZTBcuq+/vn1s4dVXJpid
ESMYx4G9IYvRAdtQvVEPJxDEdIFuzgd8JhMkDG4SgNMXffDp7gHh//OhYsqvEAuh
J66WsCJsUnjI8UAIqrKXzwe+UqvWPVuPF7icPYePx2w2FsN6m5ISYx9toak30dfo
TVtW6p8dYV8tE7ajVIZvENtbZfgQu4UFb5T2enSVP+fTC+nic/sD3WkAizFxBkTG
GVE8pOEv78SznoPJQoJIGB9m56upT+KCFSR+5RSeUJwAgXkMCrpGKW+hlVu9JajH
zyjPAWugi/KNx+CcVDcQvbXu7SMEyC0daZyIj786QCAtWrW5L5YNK+EYSGTjfQKv
H0lzykeU1L+bGPpgaywTSqHKcFULoQZM3/u19mtr7V9vWJFV28+ndXXoKS3735qV
zu4+UQaD6jBI0cxbAcoAR+Hz+7ItADsLp8R4TgCXJAy88n4g70MK6SeVblrHkpTn
lVr8f8utaM8hTuQz6QpOsHJqQ9gHwEgf89HP1uaCEn+Y794+0KceEnJqZPej/0a3
nGiFY1qkCWV9dy/NZFzhUnn1M60sdNUPmeYc8dQ5FRejh95JafErsLo6blUalXwt
zyLh2dWbBOl5J14MD6S9kib9fi08V0dAuA+uHcwPoQjjbC23t/U6Gmm+5Usb0Gsd
aSUFBoR/mGpP8YAuB+axYtAwRI1Z5xkHtt5Bn1Y9d46+/VkvS82tNjJZ+C+FNQvF
Pur3omMqVphZ8NxrJZ1+ZIflhudk61WxZdQQ640GbLH63UnGGskq6KEmb7bQCSnU
yNZWrc94UdgVRqtzXwDJVT8ZjxBdsBQ7hUxs/UeLqxSNmfkwaAH9yT8xh9T4K16y
zJ9uBIjnzHpGrZ0ofoVY7VdKAMkUKIBcV3JkuOFiTTHnfnBXGdPlbw6fRZXltAPP
7hBGok/4sqUExOh2W3VVmirhpJo9ODihLnjAR3bw0Sn+PHSHvy0rQQYzxgV8TCOC
nbiXZ1S9o4Bn1TGALJefTYywgFMCdvM9S2x6ToR0uwnhfD79SKx9hYYYYLVCUmzq
Noo/U50qYUQD1TzBjnyU4v7bOzJOPYzAefJV5n/hD+wXjQURFAij83hamgGDXWoz
aOqMtg29Nlv7ORYObYV/rIt/Jh/ry0tWngV4peWiDQMGB+/AEFKW2m76j0PxRDRS
PrPkt3ccqs2RUDt/TMaO+Z1s36w/6+QaueJuMHttZjfCrueu9VFDzdneuWfzw08C
5kbkiNldQxMvYe/k2AkL1HBR8ZLMI3PtziAOqjNHtzHzg8F0FNnV4k767KmYcykZ
pTwMavO+U2XNgH7TL5JjI49kC2TIc9ML5aI8gn1r3bXp5bZQYpjkTb3glWNqrpTl
0vtlPKdJ4cRes4lvTac5KLFHd9xTQZcIGBERNJooCzN6d7YqzN1NkSLrcxCunyic
E22BHvDgsbW2UiFRaY0Bx2QndfZaZAfVscxhk81KPO9x88VVjbmC0yKqnINr1cPo
PTpXlL54PxgPx6hedq72itJ5+e2zScUDqQabimHme+segXjh58lw7/+3kPN7DTSI
PT//CYlud+GSPxhlcPfowZNGGuEtFwwmrtVJScJ8hlfXLPQVlKt5y5eT125w2bWQ
WfrCXlzRwipJ1Q3ldXAVJjoROSztUvNopbTNU8K2OKagUlZVZm0vpbXvpZzhIMsT
evFFsZBT2/2uww07bsUGY/+u0eGvKiQ2n/tyslkRe3CH/9vd3wF1wzbMGHwJ+vsd
H/XYDL81YSyRw7RWx8axYZWsVsRTHWnUsQJYF16F8ZDiRc88jvlq63l99r2vrefJ
7Cm86pWW6xntOyWE+jeoyf+hdombCZ4+uttrDyhGCkExYbWJvngC/1WAtgp4HPTL
ALCdS007WRsmUmtyXVfwJKCg2RVOXF5/0OijSNmClwKVGo9RAkRaI1+It1LCcwZ6
K4Y+HWE681O2Z1EeHGih+4WCV0LcF40gLis0UTFaPjXD0LTsl8b2ypaJpLuD13EK
4df+h8MBIVV+voa78jb7ZoZK9gEUhkqDoFaVGyQ/jiD/F4DBbdW4WE7ml3yxyvwh
Tpz7XjiqZGjLdF+MqMIYJ5Bsqs05NucfNQnhndzahrS3pA8fEj4C7mxOSC9Ov/fQ
umTasyTeyZUOhglaq0fdSeJBWp7CNbNwD8eday7Y8A2Ptj+DfmUiFdbC9h/IhzA4
fTrUmxzGmOkOdwx/p+ZiYO4KdNyKbTLHoHtwr6BTjRUCOKvchiMhfXSIZg7OyRvS
Oen2M0WMPUQkNjwFvXcDekE+TSb1zLq3kHC3mOw4Y7+J4HjBI0cElfisNlhX46vd
OUaNDXiRY9FajX0ZovlQYVhpZ3YMTPKYOWexvJhZXwzm17xhKgxlheKRiESeeaVu
36CZb35QunHY+sv6Vh03iHYvBpbm4T/Otgiiy/Wh90zyi+ms4XWyaH8MYzIJUOOb
fpxhwjxMPeS85pnJimyLxTarc//18Nd+Aj4jRlwRWkMO23TKQyGFTBUr0ebBR7n5
3MlmizQR7dDoTEQXD5seOtzos2RNGCKXMt7Hylso3KFD3baE9jigtdbjOiTRxtrf
h9MFngBK88qqCBPLKbNusj57uw/fT+YzXFrE0rLWu6iCsnjjDFFLWY07pC1H5Nvo
gAQwtOOhxvNbTAw11zW686eFozJyunFDHC+lO87aIuzDmtgUzZqudr6uxf+UDD40
t0O7kaljk/bf/5IHFfTa9PJlDm9BhO3DaIkF01Obrnsa9RxdFzM12iUt/UNYtTOO
1hoAQzUzz6iURfcsiQesG6bqYkDJ0ORe8zp7/F2brD4nOX/7VTBJdjXYekT3HfJx
YHsswZ6qDZCy/is5hOj6OoEdrnTUzyzp5mQesNVnDBql63aORtLZP2IgrF8a9IRX
JP9dPe5UGCIXidkOk8F3lmnD9vKJSeYybByd83qGXQtB3fxHubiGsHkOohj9lL00
I89Nu4ARJ/OrRH4zd6FzKiMk0BIQS01UYHAXrHHs8qw0+MVAucw0mczKSsqCWMVj
RzOVCklZ+X8lbhG8+tOOg5vi62xXr4sGqyUe+loAS3a0XUdkfhYHUYX0/C9zXhHj
GJsfGk77hk1clhL0VS1QGoUo0CcTT+hDFTT9Q8rt7mvrZAcCOrHC1Tuh2nAb9MVb
DVfKdSR9YR5fUrnDxwe4Zt7s3WIYJYbo8FGriLh1s3SpUnzGYxzcQciAHsfKR2nL
n56gDhFBeQWQbEhaokA3Ad1a3fJU9jT25Bu9FoozUeOv3ibvW1yE+jb6OXMu3MxI
awmvC03yD0KXQMpSzoMw0A9CYNmx8Vfy69ywaoLTQ8EXasxx4GzN/UqdtWZDc3pk
dw2x5tfgnIk0+lX6aOOY1Qgh8ad0/eL2o1PKym1AJ0MzMfKrIHMba+9GNykr45zE
CunrU8Y1v8lUsYkxY4dH/CdN9UgX9F3qN9UNDU4MEHrzaGIJgaZmYOXTwjNMnf+5
wHWFGLII5wfvjplWFL0VED/kP8ILbEahvy4OKj8iS19A7JdGDdHnp9+V3KLHrfQu
vnjjoFOYU2enJOngjirNe7q4VRuPzpw/lTvyXtw4rrtWdK4zxDrMWm+OKNfhQmgD
TEOTnVdySAwN8RtEs4n6g/mPBQgMW9rdT+LplGdPy07tYj6is/Y/ykCz6/ctUQ4c
FKdsQeB1n9nY7AsQF6npyXm4dNQ4yh//Yr2w57kvo8L1br443ARDLxQpAQ5RD89S
jbr+mv5jsXIuUzIE5anLa1r+ZHFN3bXb1anRHhbfVCb3U9WHGG3y4ljJ8BYP8FLC
AQirWoXQmLEO0J04ZvnTV+yASQWuyOW6bqy7Kpdb9Dm4xvnRMLD8rp3ETeKW8Mr9
kG5W6q2J99GbLkb13YmXWgX7d6IO4tKFn9H6bprWEFLV6iEqGxKgFCsNo6mwnpaF
jagbT5m+/+k8DwZsJLx0QvrYaXxoFQvvKSJlo5ZKj6WEWYbyVqvt6DSYWqB5F1jU
DO5NUHbWicB1f/3KhVzsWbC6t/XQ50joIiFzL+qO2f8Ih8SN+3PYMDvzSalYdZSH
P06IIthfMKfa/OIUA5L+do/8qfCZZb5mg3FAOqiHm/ajDN4pHYVhQkdVkjRctaRH
3x0NeXe9Nl4ykwEQCN1X5NA+FuiKseDE20zWWdeVDWxD3ftK5XhX0ap6vyBczz1n
H8Ysx4kcfn2Y/I6N1HVtqJIe65lWNiAuoIhMkAa7Xt3sUrp5nA0uXQC5udEkBLQI
zIe8GtQosAcXWd7b53i0lwoyH8+ou2ZgVgvYJh4yOgchHoCwopcseAN3TVOWMeCR
6IZ+G7Wx5QZdGP2BAxKypzoytoi+4e3nSZFKU3+oy5n1XuEeKFM8aM3BRqJbY/5t
drQVFJYpzN9ItXTmmFzGuLeg5F+pe8J7k4eecOVKSbzQzmZvqLDmVUmFLuF0ij+a
rbTxa66YS4R/KbS35QdnLyHwcE24u8dyTOf8rA2LK+DBE5seiLIQOOekzYj64vy9
+rtrCE1C7ZJ9q9W13yNrQZh76YCEuLZLg0OLGKb1ghFm+2TVluObxQclvj2GKrEu
5qd27K0WbndfuXv2yHAJRZ6Nsi2Aw6mFoSVUIS3HEqfpVFIqempFfpwuS2/sJYkB
DZ8u1Yq10OQn3BRWiTLnd0H1EvscLOfxfwYU/HTQnqQWplg+OtKg2t/BX6OJ8X6P
SAJlfbmt5a86+aLqomERb0E0SfwyhI5/59n2ASQxp3UfgnK1VUGaKb41owJ62nOg
J4c5YltlXP0Jku0SY5ZLDT+7qS1EYVJiGC0QvQ52WfGT61559u/q9++3um/WNzGA
9IhQbSx72+GAEijpPNRWCRjqmy/p6x3yyO7L1OiteQxRFP+K6XvVrm3xzgb3ZYsG
GdjJ9NUQil6UAScTVpcfw994TfJY9PI7IY9Qiyir2e4qhDmBkAnvllAf0xTbTka8
zBhGpG/jsEcBy5sbJzJCztUBeHXgDqVHvdV3Oo2Zof3ZiE6ovi+2E0QBsed+4tV2
DfMdfZcyf+K5168FT5laGZAEzh9I5k4x55q/vyLBHWfKGdwx0Vhj77PgFVfDiECN
4Y6maUwzHlflD0M/xWGpEpzv9onVUJMeyGOX9hy5WMNbV117XSlxmvJmuR65yMB5
UkvL4sFDpFSoe6LXop8ANL6HTGjXlSOh+3Tu++sydKHXrKqzogUFZfnCEJXGRlbb
5r9y2MYZSOsghifPc1exxx9BTJUVG7mzB0KFMGMrLaa0C9Fu1I0G64xRBIZ+9353
nGV+f7MpYRAbLKy1qiIFrKDZK3ZI8mgx2LylDqo47WxOC/ubfrICWFaf5nNp0r+Z
OnC95/0oJzNWFLLjzerdWa5Xv5k2pzqovQ/03ODLZVuUrOS0ztaBRKVSCDzIRJFG
7xilw2kj5uPIxFIolgbdutgk+TkTWmKlYmL2LGiGPVD4NwKHcN6X5BL3RFpbF5Ea
2CorM//wICTt6FDd1GIB65tVRomBydSHQcSvcYz1b9WKS1ifHckjJ0fUEz0q8eLw
/lIGMBcGHXhszMk+XLaAEk2LZpAoxxHu9e+++Uov5yn4OmfzzDOGt7HD8Z+brVHn
4ptmTxTIi1Dl0HTucnVXe0n1SD/ZGS/HJlRXD1Hb51e3X/+ra39TGx5I6+OpIwiS
legZTwoAnTS6Dmy1Qjy9OhwagjsTnIIWTyXYuBIAl19KuIOeVVW1tyDCWqh3hMRr
8rS8F2lEQ8PpbKIaXP4bFgijSVQPdw8tGA6pwan5TZGrmsWT8vTG3M4TiMI2KBG9
h0m8Fa/XhlTpGxaptD0yOuYuhE1kynGdj9vQfT00wlCS7XM/7K4aFGh006vxI2nN
5NAjyDTguNM56KabEi7OlVvHoiuGHwmLs0SP1tEcKfQPZfXKFHvrH3GVCz45Rlwk
JboDLtorsiSE8nPY6pi7OADdxXeSn/j6vElr0aJUEboMz0ronZXuN+wXzx+1c6iL
6ZBp9f4bdLTHPaaixX3Bri4Pwb2T424mwMpL9RVOOeRnNWub6URgnTWXKabgjOPf
ChCWoEUYa9zwijv2Rvbe/+R30JK31T7MCkR1bRGByVYTjyG1XZbsaRUXRnhozdUU
/9O8dh3MPq58ZIz0Rx6dsHLuGAza9daW8B1iEfHr+eHlGLiw04g/c1j+9FlHsxG6
zd/bzbMnDfeA0ClHB84LVSlDvSxGKQAI0XhStLNhdEDs5QnH/I4NgJuPIdKOkJGm
ral2/bRLHdmbX8w4Uz5y8wJsvsHPwfp1Z4NMO2IpjloZpbbhSuV2CurxX1E6npWB
k4IO5+Y/4r8kCju+entZl371xs6bXy41gzq3qkV/2wD3MPLzoG6ZEIMECCHb/L57
9j+CIgTuD1U8IYOmhvoqpwp/Q0rypRZSX1gtBMJy3tQF3/YtaV+tdpBnUQyULUx7
Mf86iBj6BJXai4kvqnowGXWrH9urvWloNX3ImAwk7u/pphZZoWSEC0vrUnE1kX8c
rjr+Afh35wXMxl84vHHfFVFHksvUNn3W94jCDDiqHlGhP84FSXvFkh0K78GhPf8t
KW4DRyKiAsBuV0VDwyiMidlybnwd2GqTsmCiUkCfCmtRDpP3RGkFk7VfRobbSio7
cZ5luCcGqPN5+b4s0cDhekRs4ybhQA5ahqiT6YCq0ftL05PpRuACAbuaY3bfR7pm
8ZKfpfxYhP58eV8H+fHMo+d9Qk3vVHA1dXbhdghxPnYi5kaqrT+GUbS13UYF8ObN
eie6cRdSJkk2Zxp8zrvxAh6e+mU7iYzXrG/tubqUS0/93UpDdv8zmrpv7TVSNVig
wtNQ753PtkXkK4m1vS6MWS3sJpB2jyX1zV5Iowyz1uCxvHPNai2HHTPjgrCim5pE
bmsmitzlXJo+v9DcfMlXcwU5/t0ivLFoXtmfQ4HTI8GABWzIiNWPUj082pOI6K2i
hEYGxEJMOA/U/6D8PZMq+vo8RiWIKSoZitaV3Snay0mp+7/4KJir+9l55XgJSeeN
xx+3bJT+oJZkOg4rxsw7kiTP2uST/TGzPPKOziv7YqIJ1vf9M16zUCFirhToKPX7
denbtGXSclSSt4N2DImd7Wi4zQxX7aDHXLSl5BolDLrJsXkMme/9nD5wWaU9Wm+g
xnegCvNxev6EZ+lK77YZCg2aw+uPlfA91fciVzNbcOGb5kJS7MUpt+72GhBdqWbg
wIFSMWpjV2U8XInwX1n1mjWMzHyv/PeVa5+JkxTI/SYPcEWqH4z/OGu/nRROeaTY
HCYFQg2IxYXTSQVwyGetaPI7Ar+F6p9hDOoGStkrKQuJgkHEDfm1KBHlRVW5cMv3
MzPgq2jJrOiid49VC1Hn7z+CQEt6huk6dylU7L3NYlZhYtwuFhKyvmJ71evaeWTj
KrMKY9BtbXGNspPe2DoG9FpTU8EeXo7v+auspzN5vUlxuDICZTtVrbY06gGVviHg
0Od0YBKQd+cxiQoztcgnFf2ITipMMe76WoEHgxHfwOwDzdqpJsAVOVKCKDRMHA6W
TkSd8mdDlfcJfAmHJ3uv8ju2YaEboi5mtgfeP8k0ZPm+RdxklYpaETU15uw6mqUe
zjsawSVeIxFKNSynSjrPdFprEgWE0SEs2tuMEXlAilAIAZGKDGJZkpa09HeKxqn4
INrmGvKHLGzyoxyna6H1rUsgsj68e8P+De0a/49DGPWc/wi2Qfq2jgFro+zdfy4E
JPyQNcJWgP1rgVxUSFBeDV3+kD9dVGrG21wvYMHEUjJaiCImmeYPtVHGa8x3UJBS
BRaiP81Yl+KP1JxmFQCCQWtIvRf2CkNQyiJ5dxZiVprE3fkxZjotT/YYXbYPJDRA
7+jL1G2Uijaxd+jp5dG5wucHYa1NYYWPn9HUlum13nihkfEMXbbfiWVHUDe8CQII
ixKU77caxEm2kS+UCI3qAaNGjsxTXpT3xrVw8JlPLf9UKAbd20B2TZgIrGoSrTfK
ea660+minPJibjfpePVIBAz56u3jSoHUX9mLkU0/3fsq2l/7fD/0AQ06xQQ0Cwia
JaXlkzyI7hNU3RXUV4sO7793B654s3mGXdUac5I9Ld1av+PBlBkacAOuD2G7iVZR
YfRKkqSWxGnfkcCUvgf+ln/5qjqe4QIdp/lT86TyvmmEDbhVsPIX5lWEmYRBY61v
O77Pg8CEdOCedYThE9Ik+rnmbbnQBA7wYUbVgysv0k19DWsTaAqqtMvjP2PYKln/
7lDBtJ6R0xMU7pbFunSXLcm3QYtx31G5BmvO01xDyxErupUY6S2sbDc2Dn3oQF6/
P/9g3mUZDyNBBjTCbsRSX3kZL6ZlN/20U5b2Qo5xK8CYRw1gQpiLUO6+gkAgnlpj
Op8WDQneYayAsiomwFsNghd2MNdpO7uce+OI5k7ji3QNyJlwBvi3rWQxQwBPFvVA
qfjDm30SLb2wM6ogfnqBRQHAnbzFLDLu+ks8C+4we9Z03WCAqv0vVdFbcE9z1Xmg
wv2gk7Z5V+Tu2fDA6vEospX7DDC84jYpSmlDfOaVbDZY0bJ7eIQRzG9uPoMFz8zz
zihA6Qg+zhNy+gd4lL71ddpMdMEs2GNsdfgIZic+K2vMPFPzeDylO6hGp56Rjyrb
99rAUdF0OS590uxzk0qdtFXsoZoz19wCqub1K4ODNuJSaRi/gkKD+CYV83k6QL1E
KNx4xikilMZA0G/+urqublOojhyt0jlOsnSDS2wRE1ye6fUOlrM3DuhxL3yPpfkR
IhTRuKmWPTFKk+faGuZmWvxwk1ya++eCIR4TF+4EiPBBZgfx3B5muvKltN5ptWeB
EIfKXAXCaLJbOfjdZbuFAz8I9z/ChUQMvMZUX6YVlXkMeNaSQAf9qOWSKsTSCPAb
BnIA0m9ZDT6lkeqSL4pkq5SQYGQ/Vomed4XFHMzXwISieaw4krktgzTbpmrIAnv4
5mUWuamgzdwXy+7sNaB96n4iAHZhgDzs03EWOczLqywKXoDPF0neVe7nUzeku8et
Nwby30YvieI/6RzKNWsk0qUp5ZFpuYE1AXdWVVvSNsB0lKbMoCn52aMEokrlXtN0
YA8gu/qs0oPUrl/xj4NjOizUs8qVVx5jOIohu63ckrt4deRq6OjZkGQnrn80BZSc
L+q8mD9LvLDg9dRbK5HjMPL241PpHbfJxHvg6FAlqxIF4ONXW27ntz8rpJ+46Vk8
U/wnhKwfd9iNHKG+jQtBDpFgj722I8KdcXNnrXBD0nXlOZcSgrExABY5Hh43Js5s
8PlxkGvUqffCybDWxQG40tcIXMHKkXKCrM8HjYomzFaGL8K8LINaVkefc7oNVQty
1ixqQOYV7WHodvFJ62pJNJoDTrxYJCfpHBXBbDxnLGsMGm4bVgY8uzYU9whrlwsG
weIX9M4JuuqAJvjiLhX3XArqf1jc4h6bmRlGbrBVriT6IJ45RlU9wUNWWtAMDGB0
Xc4cqK3nDnivAoArvV0YDoSzboQCN+d9NCSj9QU+k7m+sKcFpmevXn+FQZ+Ed1uX
5BuYJezfS0g4Mtxyf+fV3ADujDbCIf+j23p0LYpv0McwKO9UlLdfRAa/tOVjmEnY
nUdqxOz/5Yp77lFI3ZuqgDyHflZgET325pWN7QzlnFBXQ3WdKs7lgYVztaKtpaRr
QcdDdnRAa1DHannC9k+kyXsnRNaDJ78w79J8iOuCTpcgp9YikGI8h/rerrV0S5Qc
Ohf6hQAq4v7EKSCEo6RLsJQOZ3j8fnd87kgCMkHpybNoYtBAe3oesClpiebrpMgt
IXxI4crU9gi6KpXngfiqZBKDakttfRZq7xUuZC+Rs4FXJzJb47VmQmpWojGnW97A
CnbFBFiI+nPRkNb8XQOs6yYl0dCJv3i41QuiIrqZUCR0skBCKPjzUCctQrz86Zp/
BKNqsi1khZ82OuDY/qE3RnkOpmJnC53XyulswBknA93Vx/x4ELXR+ygTCymkmqvZ
MCJTEGL7vwwqAUks26nNP4L/n7W9YDtarhuo0mwb6jzKed8Ts6wkRPvoskYIYXoh
Jf8DX8jxy0hh9M1I/CI8s6yl2d2Rltdg2WhireqQAPExLby0bbcdOS07RNdiX7Sx
lc+4pTS/TViZRrPgMWvnMNFS2bAaa05B678cYpJpDiAOASpJklUh76Yd9aM4OOVX
cmhdsDOp4/KUdluEgwizf4ZGk21NGwaX7feOkrkW20RpcMVHE+drKXmmtR9bsIQb
n5fZcyXTH407PzN3lAjPlmQe5ekpxHiRiVDy/5aq27h0BOyVPmOFeFFVMAHNIj7W
fLLH/OXKaAuzxrF2NlqfiFm3lQJI5BEHHr7nZ9XPydleS7sGWhv6rADa1lq057EN
BZji1Ieeca7Il2J/TkAiJ3DJB5dL+ak2WQNFib3DnTKeZCmWLz4QtxqSqCZoLMRf
7Xr3OaKCvAVSYm8lgRDWhnJIRNo1fxddtxSRTYFsQuOuB4LPZRSsha1uReuL/ntV
9BQ5O7K8gqPEV46dad91KU82mxa3RNkkClx9bMAF3IFlQ+hV8XApGyZnyqGzXZx0
RC/D91Mks4LBh9i0QIRdGybDo5S9hHXRAdibxdpGHlZWkK5kADQa6eGeShFVcQZK
CCModQb2d1801UOJVJi79OHbLJY459eq+YoBS2HSDgJGO4r9v7gzmtqU84hIml1A
6cjUQou7aT9a7R/rxZJcXs1W3Fqkk51bfF+i1JC5YfbngVfRXvIv6uV9+HUOgLqq
6o4Im2ZkS+gL4OhzuWL9aXxBL0G3dV9f1QFVpqOnWKMR1rv6JJ87vB68Fro8VVDa
0mwBIarCdi0wXYF42nA0qHsno4b5/A90PX3mZMurnidiiFRM76Wk4M44IC/uLC7s
+9aDwEKMcbOu6qCeTRH5bulz3qxx+sBD3s3vCDNxuuwAXu/9xHYF8K+CVyB2ks+w
+UTS22Nes3hivrEGVCpxbArufPIiGu0/wnRE/lpKcUC7Ca+61AvMZzBx3hgEmnAq
84jWCScu20is59b24HrRnF0wyqjrsM58xqfWARdVSzt+lcGqFtDlSoXK35Zrm7br
VVthLP+CfkqzuGHA9Pca1NGmk7q5EmMTqmIPGCzxTzBOTm+DXEadrVV8rWe/HIet
WzZaUfJ4f/XrED0EEYmVvePxaU/FawIGsptQTG0ApH7T3Snb6Ue72+Kc7y3+D4Ol
w9MOZGY1ExS+K3oRakW8eQCuiJwi8pOLExp31RjfOl1DZUS14mXBmDPFBVITytOc
gHezLTfZu7HYIUvaIUPd2ZGTyxfGwf5bceJGVqxyD3OgGJKKGGnnpvHqP+kUKVsP
wyOQmXn7sEVvt90cdQGtLJ5BktG8ujcK8E6pTAl9Ru/J/+tYIEinrFSpaKfm/don
7QmqBYtbVhYKNS/R5zWs7nczarJGGXiF3V8hmPCCsCeD/+ORfZc+oq+Cdsz/alG6
sB7b0mDpq/yQXvlkjmmvXT12ICKnY5N2cc/mOXEFmqys2Lsw6woekhwmFvzKlKxo
GuQQA3CEx7cmtTGi/o9PFT4QqodJxBKuEU+Hlb4AwX21qQ4R5sdpyCBZYx+Xlb9I
y6M7/Js/KqdKkNIAqutGO/YlincpNiV9R3/+sTiz5wJCYfMfFafHzK6u8kcZKghr
rTaxxvwoZz6qLdujUmXSS1sAFk2ClMOM9XerRiebG+4wPyVtcH75zC1weQms4pvl
xUlFz8qbBTTOW6rPk5Ig7IY5LaPzrpDieqh3CmYBDAJWYkV94dWdlp1hEQNKALhl
avxvrvcNBy9KfqVU1rjHYCHc7O0vDidAY1GMAKAvgBfgFKFdQi1fXphnUWB21uks
4/+E61LIEw3RjKa4bVExvssxPWjxBl2Xf8ohzMCowqPNeruh7k/5zh5SY2nh4ZOh
+VXvnBnIZUtlkUww6nVJ25VHQs7ztasN+ZnGKut4g1u53uOoJMuan+yA6uyZvKjd
QlVUJ5kXOZutwwVFEt/MF608EERxUwIAES63huiLIJMfLGzjdH5qD99Npm6Suok1
AOzm83TSfr3oliD0KdlpCS82OKuDDLwnzURNy7pJGOqNpg89J+ca3foP/35lZpLh
NlY5/klhpDxoM8QNstqoZ+K7KFExsBpy82LV6Xl/60Kx4OODWXpITD0je355nTG5
Q6dDnURF6YXCn3NbBrRdiIH+m42dW3cZmhL3n/1MT16RpQUpInVYDfgHyEvOIQwB
z3XcYm9mIwxkQKqxKoAGO3uv8j8FG+201xKgu00PDgZnGWZoQ9NcG6CY+zMy5wB5
hkEyP1Ss5Jph51uFAqRsBn6NBt66TcLgAPSSpT+Z2PYp0nKmiTABQoSrPWZa18/G
9FV0xPa8NYq10eibeACeCwTzxhQ9Kl7Eqc7AR/aFIB7O6lqpCTJO4ewVWN25L+Dh
8bT4nrEE7Vi8Ua8k4wfIiQxHZgzH3HbY2QJbMUmmAG9tNIIdhLc0jGfW2Yll2K/v
eCihINF7gMoE36qYs1sMKyVcPz+ZQzeKZWWpgF9Q/8qPL9xQ6YKVCdPRFzG189OX
JsWoFtowHXw/QEQOlWcone3hbDnHoKLYmwXa6xJ4qhlawwdDjNJDb2VE4b4VM/+f
3WjTWhVEKnX8P5rpWQ7uUWgknJU3nOFB1WUz/GGFIcFrcgVm1HY2xL4pGrhA3xav
AvQWn6xinXVZRmI5osQTaAS/R/RvEZJASVplWMOlt2exqqaiA770kRD6550lCZWz
sxShJq+nQQur/8Hx/yb+z1PHSaD0/fAn7ChErVNEh1cz6lTFAfoHa26y+fLwDVc0
F651NXoM/9Lm/u3LqxndOr3/2ivWpjSP4Y/tX6MKbb+aLD0VpEynwd0dtQsr9uHG
ZAT5RTrC5M0f7+RNH4IEXqlu/ildMkId4EFUQkCjzMillKA9pgs1y4L4gnnFBHXr
QvMkQZHGjADAp03aHCZ9p5HPCv0Tr+hGUCOC9pGNJVL4DaiKpEm0nfLswup05RkL
6DUYtCyITE6et1w7vZ9diAqa5JEF/Vtw4rOoUHVygKCyYaL4eJam8Fmn+kH498De
uMkR6D7gFR2TZR2CDQg6X7/peAFhAw4kG0aV5IHzhrNvH23z4XKNPlfwskza5Up4
jECPXbXDgp0gelGYCzCB1rxbK3Xh2IXdMHHgYLMDsfyF7mhnIA3fxrPQHBc47MgG
2SWSpRzt96Uw9QeYc5tW3Fi8+mB/3nhK4LbCgDY7M/kGd340DFFYXzzdRXH5GVxu
V4KCMKkQdx7XLdXfsvERcmV9SmrB+5d+LN3rCWBmV3AUWB4yN3zX1MlA0dd3VIi/
8CsEpsFYAWhH2S8N/COl83IpkDrnNwPUHW3/5HcKDlUTuP8fLOo2QamLfvtdWI3w
1uM+/wgN5BKLgIimTuIB0Xy1UVj/usIGXMztSlCWIxPQK4fPUyZQumwaczsIDUq1
BQt2fIycKDi/X41xKeV7P8SAUqJfHJUQXtw+CrY8d1JoIaap0LUjpiJve15yDXaM
eyIvJwFKcGbHk6BeB1ShYCiWvvKepgep6pqT7pgQh8gO1q889rkmJrms/yRtKAVU
wfGoYXZpJQ2q4NfG14NXXsBpZGWCCagV27cgweEr9t4kYLDJzJkclQBijJwXK1yD
4RNr5XaHWdBwDb//ibpxG9xpMeCQbfjhpt4Gj8IYXlBZSrFWBUeeHNvBtJq9OBI/
uJkTj1hn1fkm0bI/Wl1DLbT9DpUcrKnh+mPcmJt6BLYe76mBFk0+Pk/KwLK+tsYp
wU/aR+1j5pXvLzF/dS2Rdh7hVbHqZd0EqCZydy02u7VxfddFCY/gKYe7+usY8Dw9
DRQrESG6HGj5zSDUziBITPCBiGlKpsBdYzBd5PrVV93zWP0c7E2QRawBc6qpDRVu
ZRiOtcTgmuhiADn0v/QNIsBMBf+Ot5vqgjid+yRPuJecQdIdByGLzt9aLRh9GHSj
r2TM4o1VK3aZnMZWhGi7mFxbAn92A5jZPyP0ST61O+TqP5kRLzkG+KFAUUC3mOeZ
ZybxDJIYDvc0NXFb95xQdW+X/ZbqL1vTKbyJJdx+zvVGuqDpIxdGwexdsmAAUN5u
VWweUOsC4rJ/mSWC9jjMOzQw4Oxet0KzvnRGAZyevmBnuLiuknBFGT3XxJAi5R4B
+D/yzr8cafBAuiivkCDZ6F8QngDU/E1G0+mLgF+17FSc+CPcdBxNJsQlfrL0QSlh
fGj6MbvcCxnjOlfuC/MOYgz+Bnny7zPqYsyx3AaVHvCWUFxssNxjF18yy5WrLRXd
bnuH4wfz852UnBGMTYAQB+aytwIk0qd42Ym4nz1+VzAfZn5dexOV3BAhmVHDZlU4
dNG4V2kWSEJrPHl/dWkFPjT0oj3VJYYknHiEbg/hpsgJG1d5S9cmF3HVGMHgzKKr
PCrGCxHqmP+b1HrPRAE/OlBpIO3suSTkHDQ+aytH+pYa52Ko7dyEJ5KCBlF762ig
hoOuQzhyV/wQRQ9oKo7hHPxEeiunsxbRJbkbMCDoR+vRdh4i7QqxvxAkSCZQGt4B
Xe2IMRcaRViwY2fjspqVI8P+T8mVLBk3IUU/yGNIY7KqacoBQYfpTKkfaIl58MzW
p74LoG1h3RjTRTsKlbJ3U74jV8lfVBvb86vZkyLuB3oYM6hRZrd7ZclwAWbhENLS
/64OLMtpL/q2cnHp4csqrLhgY+bQSPrkiCaA86oPBROg/H/cJa57HhOmGRuHDjdY
X0UQ4UNBhHqHAVDu1hGlsgOeFgL8oUFQVnBiuZ/P/qIIDD1innDxhZqxCQwHNxoA
YnfeiNn/pjmqSz+GnpW05ftgyR+IKZcBhwAJCb2hcjgQ+kb80wmhfZvyaQcbj78x
k7rQ1c0U6u+kas5sw8DUDXsa0KzDMDrPPTg2+7on9kP8LRtooUR9f103IGHpMARi
vP5rE2OIbktTv3CK3Bv+YCQSnk+YUaRqNFTECNhpAYxs4iKIJ8DGtA66FGdvxa4m
+BIxafX6XRon64sFdu3RPnrvA4qn7fwP+DDyVp2LZFXsdxAOmy+z/nTjEbu1mbE6
lQ8m9Y6NKhJUYV820ylgpUzgllWe6BvJSU7WcaCPVbm/3sbw/SQ6JPfev3ItHbpe
wR64W6U/7pT1LVvz3DDSIzpOh02R0OLuqj+DisLok4m/w2Q8hZy8RbzuY/hEtJaf
uF7w470CMJJUIFhaG906vqMzVo/5oBSpVjTtrmfGldwqjk+mtxkrQUxVUUoveuOI
48V7dMXNvUtH5NW8nBCgKnW+Kso0lfTCwrgd5tEUgq1zsJJrmIKOlPmHvDLDioMl
eHOh41URefXjgBB6GR/LC8RBkJF4oDaWbfBA4wR1bIURRLDITsnrA71D5dHzd5HY
/d3BcaxgU2b+2eYSTdvKJTXNq6uIbM8XpOjGinEe0l2qUBXbuE7vJDNri+JCc3Z9
YhVot2eoF2o+cEBxCzYI67G3d/bCrOVeqBcM2pD5toKHsJRcidGyBo27k9Z9PtFC
hP3+XvvIZHMefkVyGn+yIpuHa0PgcAldcuyK/k6SBsjwV4X4IGlB00TD7A/h8XBG
OAUzLqw9YMMxf5ll5JM4BNAfWoBBlUK4Unk2V6jwsAA0pYGv60NTMhI6rXOvO+L5
dzMCEK2YsThApwYC6C00icLifn8DYoVvPQl13Xp4yPHO/la2LgbAfSr3NJcyny8f
NRr/bhdmv2nT69zGStYUtJKzj9uM5Iu1cZXddReyn7siyKGOfBUTDsRafifbHT11
V7okBpBYuE21SH5iYKA9RvawhKTQzR6X2rXjE8XwsDf4jVAhInLy5lEKwUqNTQZO
TmJ3XZypmliACIJqa5sqaZpR6kdtSb/3+w1vLXttX/RHvhpuQAjod1AngCr+wjjX
KuBOYTcvOfxyM36v+XFCsQoVfgtXnqSj2jW6GwEOfzf6IiK45JSxVMGshT8uEggl
BdKEduxgIwBQyau3ke+gZk7PVhZ2K5Q/OPSZnZkDZN3BEXlVD+LOEhjPMFtiEo34
6HeYmuFZB7ZfPyY2P5eI9cmOuyxSeP3owMeDHYBR/+Eu5Ud2/zFYPcNGZuxzuWpF
oLsV4Pxlm/rEIr36JadVYUZ9W58+c6WFKGehzOmDxjCADHDPbZ/FJ49EH/t8P4Zt
romjNIIMrXTrwApxPjIOMteSpXxx8zA0keU2ZIX6I/Wbz6+IjeTrBBa0D3EK/8PL
ejA+ROgAOtZVpVoM+N6+0AW2dOAsTa/0SLVUpz6KAdByKmV2E1R42DHgmyxJiuc7
pUWpjKIMYfGh07mCKWuIKJqto3h+K8qu1qXXDb9iy64orjPQ0Svm+liA9Hqqrydn
QSzmAEGlQo97xEvx+iIRAdgwGS5gr7PBh69QbNy3nM2QRVzQGbTee0nconjkUrJZ
0GBpgZqz+fSPJ6HqI6aqO4u0VWc1DNaAtvfpFyLThAKV67q83ZuasoSl6ghzPLiu
k+W77YkBQqtu2JdiNE/ZdQLY7nh8nAkycSsHZGxB8yJHGWD+M2TkiycZBxkUULY6
YTibLpbrnzxniSdXcI2juz17ABaLl4GNrFMWL7TJRjhlvXhG7nRp51wa+JswrZ4Z
K0uUjlkgfj2MTXRTX8aty9wt9T8WpHqXq/qnzd60oyMo7xhtWYVmzW53DcHiF5Hb
Lq+uOFcLCPjG/qPR5fxpVC0rcGQur7fhM0wtuQIYOzCe7S2VxdSFT5mzcsGbBFae
BFUleMXz7XavpOrVCBwnGW4sgW5ooPQ60UYbJf6KdgmPj0KApGWWZECEGSZbfHBN
TbcsOU24mvZIjvY8CdWrjU4d4HuIOJaZ8SXvjQWAqUkHpoPDaxi/t0CNnKXYzEYT
swcPQdwEGzgD0Wor/2S2UzxnApPbOi3gNv6+aW4vWFPA8jP1Jk3ZUtwmEyinlsF1
AinJxVDxP6+tvEL7Bg40BaoJmRrJLR4BhXrpFAQIlUWxoIgLte++cXSxqjWKLQwv
Ryw4+x/swf/BC0CN35iK3vq/Eg9lddYVVXWzITWK94kyNmyz84FoYENEpGgLlJxs
NUs02eIoyU+nk4JL0gcRTWlOZxYbYJCS2ZPaIjY9HV40fZ7jmx5nf2VcwPkKLsRV
rmSehdxsEwoRvmsTJzmbRIraqqdd9SQpIbfmnownfgJmPYsFIrzDiA70gD+FQ/2E
eydSpSa4nTsSrtUxHHCBlCou0qLidz0jrUkOPFTta4aZJhFe2K6Ur0wiaTYIBONS
njeO2ccjn6P3c3ARQn71OxQqGCrR+GFy+UhRoB9b//p1Qa12qBjkpR5UXmoZdR5t
XEF0TvIxq063BrkYAES277r+G4oi/No90eXQCfv/qq5OG4wVaBCnM6WlKnA5XgBb
UE5ebfrRTYv10MH063snQGEHD2Q0kL/n1Ar3U+ASdtSRPV+DLeEanUoj2x4Nwyzt
QzZJKlDldMse8oEnZaZn2SpugJUauNi3CU11uMJYu1dgyrYHn0eKfpDZt4nxZkP6
nUvSIGvhLV/bQAv+tUVh9SCei2+yWjtL9zXpLX7VAYwoxW13SWLTnBuTHXcy3Icg
62FkZtvBjnuOM5mjf9Dw2v2YYmDje3l/YZj8qazZ3zRW+5u6DftiM+3FMqfZIJtF
pHxfD3FfItqhXCOLxyWSePbQA3QB85UelC0qSA1LQSyqH3DSE2EceDIEJ8+yIQwe
e0aFKU0rfhMQseUPqqSD7unraa2NWa0XrMZgTlbcxrCgL3bjWncPslzFjajYDKi4
CaS0+p1mMd/gB8Pm+BbvXvd11wTS3NIzqC1fdIW2NGyaaKVUW6jEKnDudyNlYvBI
XGec/j8HcBTJGIQFutDq0S3AKRIQkacthZCtJKAiuJKwcP2dGt0xsJKLz+Yt6/p7
yUngxP9HRXzRQisf6Ry2D17PgWIW4bovPpk7HiC4Is3CnGzUMqeltcYBqWoNG+77
woOvxQKrwQU19XpSX2vB7PfkaOpFSx6hqCHBdIzx7Yxtcz86JkHT6JAbHRcc+Lvc
rghyrCr2J9He9XL51I9gfYmdK7jTLw4k7zDtDxwYHbIffP5wiU2I8s5n1yne/Lxx
kNEvtTkPuNO4Wk1eElY85NXWodG8yOdAOMZiJVIdnZ3AjY5s7JhH6K3FX9vF3g4k
p6tI69kHIhRQiRHa9g6A92s05jN8EWb0PNhRCg0+80eNYdtwL0gNyL4tlrnyk0iX
Pxy6KwpsCcmGwXwd98UIP0fMTb+R6Nvq2tBinL1xlA3eF2asJCvq7V5vyDgW9uCj
scJ7NzSvRCxcSYwl2Pkwf5u0wzTBsqRfh+52u3cPcvKWkMTx9b61Pa9fX6YnLvHi
l1gS9A0FzKIXFehuWiyCysK1NlA272d2F7sxfOy6jTNTCDkwsdHnKKacoC5dUsPB
lgqYcolmM/e2gFEruzb7Oi5tY7GPoPeAU6VsCJ6wM8N7RNmCSGfDmW3Ylo68LaLh
yijhU2LDNiL50GgQvlzV9u+whem7y2xAiitRADw2e+pgn14U7VtS8RJ2TT4kq7rs
90n4RRkQppeG466tZ/LR69IevgDQ9xxhBBfSUYOMHUJAQE3AAS16J+tD28sEoKd5
l9d8BkpXIzgqO86XpDjsqEEHlKKr2QD/HDisN4g0WJRzuO4VQ4cqZBVkeQG/dDqT
M0WGXU2OFL14N2Ioj/bCKw2JxJcmsaui2bDXBK5GXm9DGlHOXJJN3hWUUXOnndOu
vk0bWDEId9jNsmNHL8gOfNSEVPG6B5TRLG/PonmMgI+/U2/PLs7rmdHGlr5T8r2M
GkHDV8WDvbrZME0wt8eqhXoKGnkNlqAXPDpnPW0y3AvJU+UEM24vj1sF1PzgomGd
oD1QAhbMhF6wyeZcJb4SUDSQnu7pkCq2TI6/XklUY5T8HryhR3G2HtiP8pAwA+VT
BE4iyxG5TN4NMMzNt+ZkC6Y3vdsDX/O5tGVnKgb567spXIIY1aGa1M4qdDJ+ONcK
YRnbIe/jZmx/fhiWVfPR/gRc7Y2J/IgW81+Nx8k306gaNyAJ8z8h7k7UQerxDKja
A0X2O/LOUsiS/q8SNjdxfu1pKIs8HelWD/0PKh1COfa3P9pToGZp1S/l1pX/fDgW
k4xqThqT1YhcsAcRFuMACuu+SI2zwH9sB28oMb29arNvZG24lzP6BJiftvCYMrYh
RLIlGxPNEpHRkE0b9JhXCdA12eY4+309kTXvUHahd7MWK17mWrHX5P7DZHzh27as
eIEhRN6is+PP3SjhCODZVnv09zh7P1GZy+0rk48RHb9uk7i8WASrWSc+MNeJSH5h
V6AcmmyeWgkkYpc9Xy+4y/ejG+ZH65gZT2UGYv1qqPZ48+cRgvgwymwD5wLcsGLt
+GCroC9nPIXdCt3phPMmWOC+quP16NqaPdzH86HxfutMCmMjOGaENTO3ogAAhFGL
mh+7JDrNe6B0bpyEOuOlNen7AqNFbOI2hqscWbrl5jhMXKTE1GN6trRgj2hgzfXj
gzuDw4iBJGYTe+magDKL5u06+LDYh18mbrZQ1EMqRpQeMNRBhcVXgzBNQ6iiYjKy
5QHc7zOP+3B/5UsFo99mZSWP9b+VFFhFn25yhEpyfBpu/yTTB/uq/sI+B2rwS/Te
gP/+32yJWGZyrUU65iugHoiXUH6et5z8vvlZHezRgGt4ZRI2Ek78CLiWBz/hy6aX
5ykHsPQO0HWdk7lAD/ryoDNey541Uk2WeRbtCPsJ3WqJHaq4AoG2wsxlbBJzIHTm
iXoMs79hKRyikYDRDIBrdcy2SLpGvD9RlgwX2GtpV3qZxrGwEQ8Jp17pGdUZm8vm
Ksr0hzPwGEzdxUK5+G52Mt1UPJG8qV3y5Ry6om9Jpq+WEa9+qPdZUg9ZfPgkIThQ
Zacck13fqRmNq6+4yucKYA38/BlW7hIkMQMZULl76+WHU1x+4+hPLQt0lS8Ji53f
ZJ22IyUUZDm70FjyZ1nP3FQBGC/oqC6bdVOmvLkI3BWultCw9lxvHLBmczQZ0gEs
RfGwKLGp6dg8sB+FZPnJvvEAGxxlrP8wSBe9723OqrzsOh64ShzF1m1wKkl8S3vk
TpdkbNlJammgkEg6WKm1rmSijXuBus51HGfVgsuKS4+OByYVNyOWMCdMBcNhNqqt
tuH+PoR0UqtDWYptzsH8hJ21er5mpkh/wceZnSnsIzcul6TaTBdqTBi95+lFFAw+
9x0cWwF6nmZBVXizpx8jns36i2FwyPx1fuE7u2GrSiuvxmvOo4hVeJo1mxCtuL4w
zXOHp2/ec8HMpcno8DKg+xcwRfcgE9hxemBBEzDJUmp54YjZA8U96oV0x8PpjtR/
bnJi60uPbfhNSr9p7u20ZtY8mzlga4bs/brFdERXKkoxFh5cYQnMhVvWlY/dMCYQ
iOBhcv45jDj+Zc93ylxwPnDjqBjQm9L9xPJLr7g0MkYk8fysaJUWiD+KnVpjvMwx
IHvj2OOJGBDyKcuryQSIxjNd8Pkr1oj22xqz7KUEfKKrDzip8Qs6j24eLgv+kEcj
4tVzDXOfB/sQIzAIyk5Y63bizFdrtMy/Tju8QkH6yWQArOCbZZWyWNXtpKHS38u+
Dd/QDrJhcy2Tnc92mKZHKhCUfb0fZDP2eUEbZaPIg7wha+S+Fx9N2+aUkXlR2HU7
Livr48c/J1qZjUT//w343J28j4OEnAaUUH2lafRRU3CU5ZDtoYahpL7L4B4+a60H
npUZ735H4dnC/IrJM0HKn4CT8pliLfjiogu1xQlgO8b/VUKqjZZk9cRKqGgRBmzJ
KYDyKX+Oq6u4ZNWcEbhI5A2/qxtGCjHR4bO/kvfjyC6fj6az2Y6CKRwBsmQIMcP5
K0Er3Q4AS0LfncwAnRJPMMRwTnl52AX8U6OehZljnKTU+DXWhi4OfsHqcLwDUJAT
GrdnSGXkXznzajnblwgtd97XfRMDeGx6HzT/yN48ttIsg+OcxwQ8VkiXr/5HSkQS
0gQlx1mBcxMIoWb2oA63K3JkXws7NyiNg+sjzJB0pm3HnuSGi0A/TJPF6nC/obeY
JS9iQv0vm1Mc1jvX8GTlGquvUVKWlHGqA6eJChH2aQkzMxUHAMa+IQENl7zO0DBz
+8dWIXuQVgTbiQZKWn70fHbHWIJQMEAQ2dQKzlWYHDEyjgMp5teBOEFH3aKDt6v8
zsu1thlL9k6SQDtSjn8+T9w0D6Ca9wMLbqJU7BrcE31S89CtpZ91MW0k9Ih8cKpE
O7H+PUo8tiF/FgB4P/smRRmEbfifdeWL00V4g7meygrkZcWbo/J//UF1J4OZDjUS
csSvEHWSjwEvXMCnamsNjYi1Y7Dx7bkcdYIGgUlFzesCi4PyafDTC52K6rwh6f92
/a2qG9kAyNEzjtA8uvotLhNLaNTJAwslUg/pgZYxu20mr1wD4fqC4RsukuUY3k3j
ws2FpsLHYZNRI8EUg2Xrv/bGXE4m4HuqQnHTeKDj0nTzkmvi56oOAgX8Vmpc2VTK
kOMo2H4I4Cy/r4n4/LD3IX3qypGe8195UqoKmiEOFaZukVRhs1bcR6aIdxoEEXzZ
K5x33TDoki6bsQdZrL0ijOaPlOzEyMEsIHRu2ViKjM+FKHLtDnFSTUuQw2NOcA2D
bqy60SeBVKhHmbdp8zl/24ubG4g4GwHbKmkk+OdB9/jNlj66FcnzBGWZS9SWEY5+
TKVuHH+Njf9abaL0/K/Ck83+85QttcHjOddPhLYeaccoZDd7yq7NUtbwfQzczlYz
BrH1jg8SljOzRAuCY53X7LUSJwK2xBQqLC5w1WbKD03lGQX8gi3hZ+DA1jKHBw64
R3bLuOzaC+ELRNZH1mKoVeu3kII8t5hbWHk0m+uURUyDnsQrzQ3i3RTyWXJ1xfwx
wxiTEID+2UitsIhFQzzAV1WnhSInd+hWsvik/7SXxvHvUGYu73XL54U1UmD1xJcv
ENuyPALuiK+47rkkuaeUgnKdqU5viFQpn91MKdEnK562n1gAS9ThCB9bDY68qB4U
cjRJG2Y5l/3lnIgeyBX7cdZiNGO387o+smlfosnm7UQ2p79Kr4MGPoMKv0kMCGde
QxXw+lOf9giqvFQvv+et2D5YM6Kp7VRDUi8I/6+IJLb/z68ni52XB+APaBVOhQDW
fyXj1zQiVdblVS5hrrVOZ2EIYDALq31I/RJwoT2r4VAUOdY65QYLeK7qxT7xdKZ/
c+CtmkdxF5HLgI1l1JdMHR3lgscdQZgZT6S4Fr5MSzbFumU8FYdJBj84mj1vaAFF
4mho3GPCH4DXvucD4B6SvpvBX8UOVKZys2fuqEV/aP/7I7DTScCyuC2Pl4uj+BOS
pjWRCV3smpYePUm47PZt06mUEEB7wbtumQSaSZElxY/Hqw87KQoRGcMG3PDHAk+L
9y15VOzqjxRV3mbhmbh2bjzoiwQINHaNkNvCyJPrAnfaqQdKmEDuE3UY4oLf/BkL
eLeTaeLkeKIaeKtNDzE7AIJ2J1wbeB02akMnyIfZgt8INEn3uDD28rcgxftMs51E
TIj9BJuPfZ6Bx/6Xl+ooQrT1Rb2In7IbQxxY66QBtOaSED3lEEaxtAPgxLP7uuGd
S6Yz5atdf1+90a0GNt61BFkTVWPxhQMIMBld7sM+HRKUoIB7g6zuu8oH4hMa2Rj7
MMqCA+xlS5GrC/lCh4I2CA==
`protect END_PROTECTED
