`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KsXu6eePHWXArhGcjrv3x7IylLPJL1LIIiG2c1wuhiG7Zi2FqcvkBr/Sgsy+GqQI
gpmJUfcnRBS6cBklXclLl1H0KDBHTP9bWs8EWYCl9Taepc1dyNjZxnPILmCux42A
Qaf2CtX7sjz6xelL24haJoho0GsM15RCG3ohk1qfic1F3tLi1TfwgwqIRmPZRAPJ
7KnqtxruLsCYPxPPomtqBBjCf7e19WE5vXmaUVPGgSkRnF7QZy83bHzcp38yI+jv
FGf1nvWULQItPcUk7WW7iH+RaNM5wQ5i13ZB+PJ+GwExUmS14/0RN1LRt5GGbuut
9psRLX4v2JFb20GJirpf2CpMq96j9lrfa2CXBDLtnRgyfe4400vsM7fN4QNBD+4p
HgXDXs5yGNPeCSn7GWAaKLW1lrmpQWN7mIplk5zqo1Jh/2XJWCS1UUWkmv0Cfz1O
PxHSf9NP3MlVWeiJFJuwd6yoCLPeaJbsT/jkJyJT/n/58rZHNgFgO6Xu4S3I/qCH
6/NPBUPmU6LklFktTh8+sP/6PFRwmkgbY2ydsBFQzZ3bRv9kEvihaQHY+ZYjqVm4
H1YEBRyUJEAOpViOoIR+EWQqjOm4EmNVvaa2YJgnyB9nZtz7fOrGubwpipUdhd5R
GmupS0B2ovU8scrItE+RSbZkjqUhuQSzpvmFJjF+X68fBKPFmA1/MJ/SuXWe6Htg
hVhbvtBlmNBXhmk8KamogbCA4iYtAY+v1qGDVsF7NGXJDa3Tc4kAXrhv+gJseQwt
bvD3oyUoZrPG+ilZokIXFIgtkhfdCsmUR07JOHcSsaFYBjpb+QR0Xue6/cR7iGKY
vNSfSr7S01qq+oNH8wcE0u/7c1Ti8PFD+Cpa0gEz+CnE7UqFULE4AllIFl+pE+h9
lewjfpl+BnQj2ZP4+xJiJvokbRXdw9XH3B/q0DtVqbqsYY+NWfkFrmZR+BlEbx+W
y/WzjzGR+vunL70ZBgCE7rKKgKroG0qJf+6EA/OOD2B9xNFX9dRYKrET1RlOK7nc
L/z6rBY9t7sTz091UvEtQwk5Tz0CD0MMY+RhNR1SuePtDQGnyfTYr1lqRjNaMQZJ
Z2/9VUx4QQpNz+HExxBQfx4Rs21PKX3E/xwr75kWZbeUc1UBi1ugjf581c/096ZC
4h6D0GnrJhi4uLKeHP+TRTsDr6f30rcF89DilHSFLYk=
`protect END_PROTECTED
