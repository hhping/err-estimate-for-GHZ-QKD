`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uFJ32MyyZ3xW/WNd8iARriTQM30LRGEdJk0JM0fXwsfhnXY3dB9zMEXcHuvtU5t5
N+6hPUT1fmGMfk+AUFtwvcyA9Ne8zKmqOJdpg4AApgFcGjBE2Q78Ohzri8BTnvWX
XjOyUjmuqqG61kakl7v1dKaqcvNdb/1JSqp6/gG13RWgV/fMcRmSUicQyeZdCyt7
gbA7zIvnAtZRsOIqijD7NCxdn4NlDp+J9bj+BOCH4ibbBJbc86XdFRrnd6Ho6pHO
3wxp4ZPw3vxLRdzGdyzJdCHvzJZfdR0NWZUYyJH46nmV5MI7ODFQsRiI8TdOZhLt
N4dFsCykMZXDi4Krb3FEvqz9gk+T5jy7IkKb51Kj02zDQd3RAkYfojeqyd7JpDKJ
75MQ18JhNJ5mAT0BV3Uf6/UUmM9L6BC4WW1+nqqjkcp42wRjN/dgdsd6891rNI+Z
Ll/dRExVoiFvcWpdN45CDPEv4myjvycNUsJTkTfOdVV+2PKbXIdN5gqPlx6TjZ3S
G/gDJRSc2WVizdVBc5nqEM1nFp/bMabzshe7jbRTW5v07ptObb262rLJp+UrZO9I
tODVB4nmLunDW6UL/XQCAEabpN+jrx/pQ2uYx3qgqL2H47RwQsIFFyL2fuAbAYiX
e6JE5KyMtqouWthC2Owwmg==
`protect END_PROTECTED
