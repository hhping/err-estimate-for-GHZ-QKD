`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HrL9KknyFu7n34a8nrbTv7YEsUhSqIewmIxTJT5Kdfvge2jLLlvzCpEiuJU7s8Ki
tOxQhN90Nob6/RZd59FGAkN1LnxJdcInQeYQfxdv0VuRvc6ewFKMtDin1v1i0m9H
kbkMOQptOaK7lIHMmNfebwctH7w/TgPlLFyKKoVgK8G4KOlMvhC+VlN/mlYkMR4J
/rbbr7v5yGiZG0SU+YgTdLPHeyApnObUJiFObEElhonyhxyGeUkLJbYntI2YdqZv
HgpGX2or5GgOo62pF0K9maPJqL+B7IgWkEJnA4pnSJ6diPMYotFL/Ych1zJGcHT8
jc+gC1h+JrFynVcNQebulqfXyI6N5Z1uGYFJOYW9GupEPEFHtDrRsawLImLiC5HF
RRty2r3yvASS3SvDmgyP5oCuLxWLPHyxFtuW4dHAQLOWZJct98a3R8klc/strExf
2zzI+wnJptdvcMjS95Pc3oOF2dN330G9SVfzkAo+gV6XkEnIRXrcFpdj0rlwZsfJ
YmsJ4v8aLOVLl7Rqc12QaqvJ0kWf7nc16Dy+zZTaA5FP92GdWzI3TbuVVbXRRujf
erXKNBUD1knHhgiQkOs6g5b/p4g4lcn+1EyHr6hgKpMNudilvqjd2zCbb8Yy21MB
j36DXaMSwu5XBYZ5Enh7F4vnrXBGkTkGwgDJ7DNGUfFe/s2nzpwGcXDGCKfwdT8m
eGak2BVp//wLo2pxizFF+RZW2ipIm1wC7JoJ/U7FxRfSbwi5sEyExogUFdrTJvs4
27M9euAMFhhFecotVpGIoFBWdReDuboGZ62JDAzxD4YEL5EBOU9yoES/TWyKAHXL
eJtN88fTlzAc1jLgeaO34mo4KyhAkHcndeRC+UfjX9QWT2VihoVRoU3KofZ6UM4F
wgeh2GHfrNI5gYbhmvl4ljimR8PtRukGoF11n/I+hS/UJgkGL+zBycHZkJnSUhc9
9YzxpBDRRtgek4FDovMSc8SY3/wCKgWUgoqcd1yrSVv4DEgUHrg4dy/++7zV1W4v
XRM5mLwnGlldNmruzaQfuIfPbYGMDm3fzUq3jZG7StAAtS8P9dVqbIKP1MTIP42p
xfn++392fRDScWcfBmX53YW5XUJfwYf44khB4au/dwrhmMyHw2AhnL1RWpPSnEES
YsqT7sRAshdJgutPYwkRrrY/AeBWIGh4+7IlJwnlymMJIlUE5lK+//fLVvkqMApq
CKxudUMDFDlikR6tEtEeyMWhS8s608sNbH1HWFHjt5XzB2GULKijLuQKWk4s0s/o
K8xzwAOVCzhy2wEjb3sb8KXVifC6v+HEgmS4U97ANEEBYQmuCbhJP03mKu1VEh41
lLsf4LMIWxcAzuJSsy9rEgGg715TAw5db/sCT0In5uamqWQLGJMmKPOT7xJ6it3i
Dtgj0AMAIn/vZ151S8c16HF1jsYMHZvtcszqoHSuQ5EiBTayxQb/ttU6gYpakqvY
pHxFGQAKBN6EeUJc7rJA4NQ7ITl4LFv1IhPBUS3EjS+Ap63Mv4Fxe9rvgP/ADWJY
3poM5wtH1iza7tc2L54UNrxtyfhOM/9B/hmArTuvxUOvaGy0rYqytiI/wM52kkUv
IkmMWqazQyRmXw/vdlSiosOdOG1CwA8sejKjxScnZ7a1PXxBYCK5BoIpIagVFXNs
gtQmaLZWdAsmCXvceYBsPxzZTt1m/E9NXx5Hc2RL76FFsm8uogihOIFCLKjA8Xmo
CeNfRJghyHAL7ShlHgowsmtI7LVdVNBQe6XFG/ui7qecHJtH7GM3c23FV0En468j
/Xs6WivkfHAlVryxIEA2z/9YQgDssupjq6qcbz5DCGreufox+t/9QdKtu3+RehkN
96nQyAJVmvNVla9cTb+54M3IQaDl616P/OPQgBdo1VyiZSFl9LxntBbo9vLX5xrf
K5OTt4Irg8kmnnbIUYhajMLN9Plofnn+gOPFNBM3fGvfjCiW4VSadSlLYWh3eXi8
p5CsL4+Q9ydQWCQXwgyqlQ==
`protect END_PROTECTED
