`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Aw2MWdo+Y6GSx0ZuvAbOmvr9pnHu+J709lcm3kdtI/jl+0dHU2YQEsQOvNFCdlIz
3t1TDeJ7LS+5LXCJgKlmJbIkMiiC/M+o2OqCWCkHr3krREfBV//rOZpnh+9c/KrQ
M9YJ5KUnxy53ozmiUP3rKg1NVjeZ8fGtvcuaqLMTcK5CDqfnUpX2gb6YVV9nT622
j73H6z8RVJzNjB3BN7bm3CqHA7nMU1hPI6hUVXKSmSmsMLeEkOII4mNMWJAjD20k
OV8Ssuns38uNa5ibjEfIcWObUY3P8FI5t0Ea8EPJMpz6mzQerXArRWSCi1WQtW4m
hv19Fjb4mLeUj4JTp6+UZ38Ha48MFXMKOzNanlDfh1cCeSefxUHv312QPkyY124O
zD82skp2F1B2M2i6EP/YFJmiKArkksSQtZEp5qMFstnjZ+4avUGn+RknJrVz832g
5RUILWSgOjfpgCBM9JiffLXaPID9UMMM+0B6/GgGrsWoYiNzx7zFjBFE/TmtwxEV
F0nktQZbn8Z7mP/bqkDDQqQG9fI+kVwDCxN45BMGmgo=
`protect END_PROTECTED
