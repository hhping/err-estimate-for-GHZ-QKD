`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X0WXWTJleZb8dfPnFZHXt5Df5BFZh0VNpjfeYCjewYxDuPUT5uPlJ3qwOto+mg18
rLpvW/dDYnoUOxrAwMwoU3hr3/AEiZQ+o8uQ1WYIY7ItuwQbYXXUNPzi9b2QJeon
EEC0fXNXXGOmOfhY5l5Es44cqDHi3fSgeVjTWv5jpXFkbgVTc8hv9+csj5yGhWib
PsN8zO2P3/KD/FWA3E74frMK6AyQgZTfuLp8EANrCXkO2jJhLtGQs9JamiS79fyH
OioY9dsjfroqDjhBR0a7278yjZRolpkMn0MGq6Ro4MnqZrARvaWVL7Act7xkr0fT
1gPYIAjuj6z1cBNn8a0pAFDHW8PZnUP2B0C135TOqD8jNJ9UJHZkrtlDfB8iUooN
MsK3/KlLDbOmJFy4l4THpAlo2mGqNM0cfQbNXKSe7kbB5LdGJvSjOg12YgqMK7sV
/TgEciKt4UEBCERxQVQtM3aY5AEAnXtat47od17yiSYVoOO8mtwjVo3ysj9utfh1
YC4R16PB89iKmsmNX5qUNHCLyHxof5EXj2/fLU/eJa3OuO/IWss3AQmiisjM71D6
dIXKt3e0keaAd+9fRTWhvWV84STfJ83dT0itsHwES7XFrxAGNS16hHY2qNdgBaXK
16ElAJSoIInAwhBNfMK8WjI14O1g+M3jAEqC35EpsuB3I6pQpEutt+ipHSzFxaaT
utFN0qxlp6wHekUZgUnXV4Arhb5JMo8EmKiKFY0q7/CkaAxcrqej9OnBpf9Wioav
PVlX95oPQHcc5TE6jBemVg==
`protect END_PROTECTED
