`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mhWipYMOoz8FbunPC6L7lButY4p66+fK+pXkxKIK7CarnTvFc4jgMNxSPzj4oBPq
6HRjOJzNXBJpVTGrs15M/piwd6D3vb7TBuPSZ6fGFuiS3wweeudWQ8TQXN97JCEC
JBI4evQdRZfSuzeqSobvO6+eRrChp62mZZiw9VQ3x9JG/BjBijxVaU749qIHFh/h
oAGa3SZVtYZKIytsZaPyrIwdd8ri8LBRu9I4lvqpCT3aMWBdi3Pnc6mHF6dncCZS
jh7BFryJJcXF2odLF2xOVp6cTvvrWKNXf8h6SBdsry7FaV6IzmfDMfAhqMsOhih/
FeuLRRwC8YY+mSyEfps0TdT9RCLTVErtq3A4dEe+jKYZklhKn1nPX7pHa1LX3s4B
2GcqWLyCJQUUcZBC9j5Bs25TX+kGDwfsRvqv3M9+Oc8dEf9AfZLxEO1y1kpCCAzL
HVero1csdy4HIj5h2i2SBCOydktBqkJnodF10Ibt6iJLiF0lW8nh9igeL+aWh7NI
WuCf6eKGKuUCDIcuZhHYkL1dN9ObhBSg9vyeif9CDAM2oHMMt2pu4RcymS084GUm
HR8TMNpqaOsAvxeFD8H+ABPQqdwCeYGANdzt97kBiXpwyIepfoDW9yrspTC2LXIP
bnxigSVha4pyqoN09HGI+9w4p/X+cXizOIyPb8kzzLOcxLRAEuiRJO/NYgnGeSH+
yBUOZNnkS3LoEJ/SL7so+qED7N6f7sWtsI1Glvakzqj8YwPzA0quZ7KFhVZHw1JG
mDsouBWHbRsEqbRygvK4/acG9Vgp0leeDYSs6dGBvX2lh5cv9QiBkE5y5fKwRoET
7ys5uwo8D08PKqc7qj7fukhZfz9S+jLIhDdby2DVMNNPSD5Z8ojoKCpfmFZImmEc
ygxK8++EAB9F5TUVBXH8Ukbtw83Ilhpr2dBjc98rrFZIMlb7fiuT341aa/mWAyfI
loJUsGTbeosI/2TD18RQ/g68Kv5GTA3xUGopwvfyHDpGDfjPurlK+Pezg72bIvWl
5NNxIMbFjeIXuRem+PkyzBBnmMFM8QPhNemFfv44oQjKovPMrynDLi/yzhy0OI8U
C4lm7M1dpr2Oc3TPMDkOusL7vyza3cEO/OemZwPw8W6N7s6I8Uc2t7aHQnIizzTK
GyGRiGdwLU3H6tpoo2vGIuQ5SevkPfbYBnifee7Ab4UwchZ+3HAxO0I3j3bhgKVA
4qTMrzAzL0pgLehGnVOUhBOe+QKb9GYMJj6kDK2yCL6JV6HIgVrg8zRZi8JA4qkM
EPA2fCjd1T/i8qPymf9Ax8qaM2o4OOKb9wSOlsGQYSAmc4XpnUCgT/DkhWpGR2wd
6H8tuq1wPltQl5V0qIj18POl9STKWkqREf2GqvB7MvGc/vTIv39ViGZUQb/fiUqX
hQnkESoeTm+or6Kg+/9+leo30BGNwUuMGFhDQ7Pce6AOSyXG5C7frvvBRaalSbHJ
JtKavOY8xXq67M4Q7eHFSuYykcNL+zO92S4todJn52l16/UwYxf/uTvfpwKneHz9
7jrOqpsTgBOs5eqIOeoTzg6xmyd+TzG36SXBPwoXEEMo5LmvWhyw3tRwERv0miHh
sfIoUuikYqGx2v3V9TPMkTDmy9yn/KwwsAaxfpGSFs+g/J4qaY/Kp31UZADxjuot
0ZbFeYgzWn7Pe/eXdVf+od7wkIyVFGn314ndSXipVzBWL30sDebwYAZa0CS2WTpX
IEzQSzuEJ9SwejiWMeAJBULEUBaDLxB83Xukzv+ziInJO3l2b6rP6mrpZXAsl1Bl
7PS1TxiTHNBCRh+nmO7wvkJOEaD56lFqujyiaGOaZRHO4Sn2w5V6A60Qe7shI1Ao
QoAGwW3MRtMED0gUlCSIroN98B1aYcP0VHlC2kPn68twt1qiA49EDH2uGBDCN0j4
O7uRtLbaNLQjN36kKmTH+5pGfAA34PpzPsu5vrTpnuQywNevCS2S6Uv8FeQdxphh
TNRqOI+lheys2ytmOYAp4I92hULKbOVyfZzkqzVBvwhNGO1g+CaCn32I10lhhNCq
El7HBxcNenuQ1w+9cnbq2rmtdJ1O/TacSD8lOvEKI/e8Picai5KwA8c6waJj9Dow
JlGv3OkYORTm/LWlEtqLG+B1dNeifoQzUgNbu4ZHi3QvNAtPDwwmevYLETB767zU
TgmiohTMSAczBkL7I8HIactlHeQsAWaQmqnikObRkShCSr0C+Zc+dVhkPKWpbgzM
uhDNzgt/xSG6yRptGHHUEZEUuG5OcVCQX5XjE3VhG15Rw8/0mD24KwKFPLp4fmwE
9Ehp6G5Wl1bg97pKygLkTyzQ6oTjR2jyoquVTlno+jx5WaSjMGW2ItlsN0dLbRSu
`protect END_PROTECTED
