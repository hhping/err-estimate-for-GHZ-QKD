`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
92MoTn0uoRzgcO0FAHHuGfIFmokL2Cl0hDPVBZDS0FqfnTqygJ4M4vsan37FyIJM
JF4rmZgTPII5+OxeUaGMMCdMcA0t2jnC/qP9GJz/gyqyUbyTSA9aPDHstzN64EWU
cGXAeH6MZZzMIP88Hmy21Xq4PI2QdQwsLW7mFfxewbds2g2W2urESqmlxpfLjyvs
uaOQRzvh08rUQKCf2/evImYwCVrB2US9lWN01oP91/floRboh37aY8GUDneJOigV
dhmwS4aEsf7jeEir3+76N22m+Seep/pWyXYcCVSJz8GjPAtPd+aTKhLoAJZaHDIM
EDi5Cq666f8PEi6b71Vm8KVZoyDS3p7F0AtqGMnY1BJt7unSWQJeK9rFqCm57N2C
kxY/zEQUQ+UTqFG3VCQHCbCr29PXcyjtdNskRklOVyhPyLU64W1GxIxv/VenX0Ld
dypKtER9uTRfsbrWyWnOL4RB+H9mFyTCOAHkXzvnCc7u1DS3te/qkn7sAd7rC2xB
0Fi7dqfk/A3SG/U9Vtz7Ogxjj0cAypWW8A2dxe16iicOGRTZc3Catzum4i0sq3ey
aL7lS41anW0ndeSmvlm7JoCxrKysrYhvlbG4rM2Sc4cxusCn+4bIyBjvGT2A5tyg
PiK6RvQcu7g16fIA2CcTsBL8jjEHz3AjgFKDK+ijZMnvf8zYHwXruWbcvvwnlsrI
NGduVnRlaM+4vGNsshWmKwtE3rcsltoanrX+E+8mv6gheKqK4+SJGESzFWyqGJTR
klYgxsC8Xe2cbqZ73x0tBd1joxFa2WVNHoQyjaPakOmiIyEc6sZKAu07EJ/9BmdE
LTBQvFOv0Iax0yfGw8DySFyP8cjnQ1w3PEBxwPfJO4qPTFGIpy667qe6s2rypmwi
QE+pQZPJ372rp3f3g7bu+FohQgnlQItmMW0AGp9WBAzpa7knb8olFljW+SEoSiR4
h6F33tNcYT7IFQAH42dwE4mmz2yzPsmOOPd1JEkIhA22caos85Z4lR+b3Wr3QSIH
6Wqc50VhDbNgPsIGpkJ761ET1OwBIHLm1GcIw+8B1vbhIHF6MkWtNRmNAYAObj6D
eDIyKGa2sOWR5qUIbpSkveRZaLEARWtmtqZfw2TA4QtbROLRGIy+xvrc4TwQoXvn
rsiGpBFFEZX+hEmz6adW4En+HOmM1aQvzuuW8rZ+eIGUpThssBRxx0mCfYL/qJ0s
EWDWoeV9BvIvb9PPgCymIS4//H+eyz/cBJa8bnshaRUiMscHZFoNE3j2ptDPI0cQ
OpyITRdHd/x+BDfIhCpKORbSXUo+35YGb1ngh+SV4JHmojj1IlW41lF6nay6DNVg
ike2K2OmzCcWlEz0hbXrqpj4KG/U1N365cHROk5keGVNrsCrdToAmYHSAI+B54Ye
Kj2w7bxYgHBkRYHwjy/es/xZYGe/+3xb++ESTzv1p7E0wO/oo/SmrXbFXrlQg4uV
BfNW8ySdEghKTebA6CUARn6MBVWFSJW1Ld5Ni7tvP6HOklKFXltoV3zkQGpX3KYq
24Hm48Cn8c+xx6ZiiVjilUPCp1EduX15Cdj2JoNWQiXpu8Ju/OJTn9dqzu0pCkaq
ed3EjjlgdbZ5IvGyIsbFd11OQP9h0WdRqbSmt2TZMRXxncu/y/ScvaJ/5Zw3mw66
XS48cXHmhTWUxdKDDfmaZ3hNByZzpnNgqa7pzz1r5hXrwL8RoBw6Ly1nI+QQscQF
X7hoDvEsSVJG18R4JgUaksYorTYyXG0RP2MF5lgIB4Y+/CHMumYfwbbw+eb+6335
ENurOQZmE09Mx+GyJREPO+4/ghBlABEBtEyYLoOqtRtcvFKnetBMuyp8uMDTW6gn
+daJEzzqEqR3vUIY7VAjO43Y0q6O3Dgui1peA/KL6XuQ2uIAeSBL6KSZjSJG9Kvk
FBaO2bAG6gwO05s3pMcZCZ2g+CM+VtYGrpv0su2fDHjJxf6MH/JoCsXw/H6MLCnO
Rij8ahdJ5VadGDGmfpkucmGmiPTcJLJTdwWLq/o/r3SDDiUF127nl1aDS+LAsxy+
9a40KDVBofBA48AA/MMCAFM0ZoF9uJr8aLJvulMy5oG/1v25qHlOKW9vQDuuO5Of
OzGlNOYU1MCN7juXNMhrwsxe5MoFH8Q+sUbR8gd79ZLu5vziZy+QxsepgL6rxzPu
5rlYB3eV/Lq32xiPWT0eu1XeelsZqdwZwk46vGrzUXlemly5dSYl5NxjB/kmJ3ox
2PqthQVZ8ldJwv7rV4wjkCKkLuNEA1NDp5SfGJT5vLI8x5i7BHdjJ5IXM4wV+aEV
gx8fG7dC3/JQHAQ7e8KIyj2MC74yZn/4DVIlg78QDhoRo+WgbkTTU9ZCOI3WKPaE
pEnsQmUAhKb1x5etRvbiVz4lfIOWLSP6q52qFpBBwQRpzVFHZJrSwyIbDVzZ2JCg
z0qdp3Fhpbd17d2hyGbcoVBBzDvvUO3asPrQ56552BYfPgobbV9937vcFgwdjeit
PVbj8/7xZeWC9BojcUQkGkYtawrxfztIrJhHDt47xtBSYSTCAdx/7cPWbG/lPKVz
7kC8SRsDmYqwtxtQlUqYCvtKwHhv/3dT2CssYPO3MQA5m+TPjKyrPS7QC3tgAGhV
8bzzLFyXwIXvKz4MzMuRbqWXzIdB5hR9FZmnhcdr0WQFg7fZ8DLSflM2I2qcPlFh
EPW2nfLmitx/DElmrTxj7KMODIiK9lztCYvZ+ZD0laMrwla9tRs05Gnr5QkGZNR6
6hAZh3C77V52HBclzCIZ9SE3qG7Ken+Mc4l45XC6DDsCNpoSGaUVr9dgNxxL4skH
NaSr70/Q0cMa/91dzfuU7QPxbqI3UbD6pQIALVjPjUFJ23OOOV45ei4ql1yAaK+R
+LM+YFR9a3sd7Rus3ixo26xt5hHYXMX/UPADT/KnSPDyQsjRgcQTxjN5tbAj+byc
+nTy6FK/yMWwfst+OtyszcFVMFW4rxpY1Hr7dr/NLtDjRYRsY1SHKyy3bttizRFH
qRs7K3JabNdct251Kvl+tQJT+bdqZY8idClfM+XjBjjpgTcOE3WYpvX67KVKZ9Y/
5Rn+mYK6GEhJ9HM3zfmy2HjviYM5kk6UUbSoorxWNP6+4kyMHXfDHXyUKFXLRp4T
tNyfoM4UE7dCbAiMlJNb3MZt0LEuOsuu5B5IWBcaHl9h5NaqPeJVziIojvfLiZMC
E6ea/g4zlHvIUcrFVo/YQ4uNY0U+1oom/LmxvvF0vsTLfpiA0fC/QpIGTbBizIzO
zB6e9uWhevI2DyD+mD8kfoimjRD97lDdAKyc4xw3RwZOHOPPXWre5mJ/UWUWPKi2
hhC99tqRHsJ33i8RhIGtgt5QKBT47fgMAFN8lS8N3Rygk2r1HA2Bdl6Y2q/7rtgJ
6iYBrINr0oYANmIDuuUMuIq7lObzZn0fXMLfZL5DYxpC7x8HwBS8uZacxr2djEQS
1wK/U6ytC31OpygreS3f6rnNynO+MWT4HY7868CeTHqi9BZRI1vg42bDeRt7vp12
Fz05BkgY5Ly7sV9+0zb3BB0zJq/sAPlm032dUrNRtL/kfXS3BzOixCa5xYge533C
B9FpWz2W4Kb64ESMU7KBtz4hsZIpAZ8NwOT2UbcmBN93JGZM0aiVZ0QeC24QPzVf
v2zy4PT3iPOxXmFVu5n0LnVBosCpQ3pAKuYaDKt+gA9EdbCgvGvUgToz95YDP/cu
AbGUUJDmOPxMytjTI/OdnG8B+xXWho4wEv2uctQYpgIN5B5sEzMo/jL1sikLwhkN
n+DEAxl1fT3JF4klLxxKBzHGfd8lODKzZE+jlNjTPVm2hKhRUsMRncqBDk4Pt/un
oq8EYbwNgJxVUSQL0NSv+2aPoW8A1KQNWDQ6/uwF2D7wWUnDvQBlTs9QMehDuUgc
DidnEX/8/bwzFAs6ddjdHXiunOOid7yApYNywigR/YnzXVnsq78yx/JoeDCCpwYG
oO8WtNpEMsUOXIZuy2in7vXNbib0ODt0hIlqJpYb+exKllqjBys4GyeYtTqwBpfh
T4NJ/BXtE+puE3zgj62LYodawvWavEre8ejRPOZ0S+ldA+/+/FqAMGgC9zpTDQdf
x74x6LD22r7j4aR5tifFDg==
`protect END_PROTECTED
