`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
31Iwfp6l4QKTbvdi+muvW19knGM0LTgmYVkpLM2NdQC/Jt+R8K1+zwRfElFGm8rV
+9iN48sGk1ttiLiXXBan3816vUhq81onp4WYxzf4UCTl8kpBiuXBClbXZd2+Tu3K
JUDRhsvBK159hZk/iCSNkKpssCpsY1zgTTIqzNQKqWOU3vwXcsuhmEEPiTorehdi
e/7pb0iryMD+wGJ8k+8CMldeOHM/RPB0SqfXyatD/RQwtYVWkDfo+iq5n9D1+mm3
gA349ALmYeV3I9S8e68j3DVr+g6mlMRS4ee7tH7M+lf57DzvRC3RtPoQk5xy4QdL
79B31FC+XVepF+N4/G0DN3rlIFIcSVWeC7e+MMJNTkx//O3oI6k/ptKnM5OYhySq
WgxUOQP2SfY+idmcJXNtXL7eCXMbxBNmrFOgXjOI4Wnt2OhOSa+SIftfQNU6K/uQ
MjQ3ePwROg3LGa4RfOVj2ZDMbOcIlMgbKDnPMfPERbqasX+5yrwvZhCJkZrImBOk
fzfKCxqVv08APtYLiAr4iXdLKyABDcqA+DZrgW3Z6udSjRnqKqhtKZMdmAaSQVpE
RSHihmcR+ZT3d/kGgNgj5rGVVok5SBaKV2CJyMwq+HV6eGUIXWtTwnlxq6HyJZ00
xkXZKn+3RoxHKg5NepuHhYNTUEYjmF6ob7XCfH8yCF6bjyiL9t+wkcKU0xE7zMlO
b7lqwm74tH7/K83S3CpD3vsBZsYdw+V7u+x5pJ6Xvj3N6GoLJ7yk9gP2KtGs9kqt
z6fwsEAv9AxLlSC/TCskvmqJ9Nze7C99fmFTf+kTPZWWVYrXVbFPgdBVgT+0xZhw
jgSOVuLxE4f2Eeat1OY5Ah1VVJJK0bElbxcWwjhD1Tv1Eabe93VasQ6wkg7DFQf2
W/7mercVYASkjN/8chXOY+kM4ImvPcJVk/Gp6D+Z6452w9CKId5ktT4aE5W6vX42
KfZKYLxSVU3rGhudo5USXR3SN+iD/t7kwpk/K1fmm4zZlvPfc/UC7TpKpVaVs6CP
wqIVRyebc0RGW1v1qmMf+zZ57SE9q/mHd5duM5pMN3ChA7PJISQxtb1zU5eg9D5y
E3CuUVJhwN64wLP9nKpxrONZ0mbpvUrH3wGsyqORn1a1KO2yyIgrQA/xGJaNBnyd
nlatbKpgMfKkVGJWznAVrjXpF85HiikdTwbwmAe6g44hMw6bs5fKEN9IHFTNIjYO
a1IBACmM0ZfU3CiK2R17CyXvE9dv/zcUhkHjxevHyWFWJD5FNLhNPOA13F9KU0Qr
VR56Femt96Ws74pZEh1i8+qP2cyDGzwVKIG1QwvTXqyC0sUSVk+wfJppPvwaY+/3
qGZkF6b3aQA0kkPnJAa6NyQiy7LjLMTPE9zt3VhHCJ5cFJXTgnoc1ZqGvr8n5vBy
rTujY5aSmtln9ZuoZubelYHwHnAgXU6PS4/v9D/7FOAEsK7WHYXr6brfVO/sr35X
ADb1MG3WVBPSA+9d6Dkremt11OW9nt1v4ISHMtthoMArwh2INouGH4OdrENdvDzN
NY2aApcasmQ/hMGEXKfrCuXUr1bYUZgUNEJJw+ggl4sdcciSldJ1jwUTuYDv9EIV
TkTOKuV95mjgrWHF5mSx7oHeNKTyXUXkdbnVtIrIuws2WHHKqqkOncoRv6jVMI1v
ebbJoZELocN+ELeudHpcNRViof5QevqQy8Sx2IDBlNtDRGhP3U/wsrcsY34X2a/l
YmvgRTNADpJ8iNhaLV5Px00Zn5CTjzo1oGJh6zuuC2vH0f9EYXkgOious3Q85p91
qDPSH0wJP7/qsiY83TEtRquw2wbPA01kQ1Qff0DtFPeNaCrTFdWHGMmkG5Nl8bVO
OCVeSNlxXov+NsyUY4ZspQZ+eq6O1/dFRg8f0VuHEePSglH0r2PJahz8UvPORxM8
DekyZ5t5fgl6JtToIu4Wpl6GBxAvtvbgtDViJPifsWGoirYoqdKV9HR+iAKRa5v7
UrnoAxCDBWnX6kv1vHQn0FUHy0IAzBHCiepTE8Rhj7qoKhLseuhK1X4sD22s12vC
uTre8Qu4bmaMvuzRowdT1C0sSxowPeKt+VGgbSh5309mOtMUYO6r+lUvDUHo/fWD
skbJWBwD7iZETrPg175EbhRQugAc0/huV57tTyUr4HkJhBlz0FPVjdFUo3Qc/srF
43lXtKf+SJohRCmUclEjmct+vwp4lHgFw5+gFXq2eUYmPe8oe8yMHCQ6gw/ogWrE
IezhBs3HpeZFNGAulmE7t2zxiKIRAegXP1Fk9bc86Y2LqdL3VaMe8RSNhR4Tkw4Z
VM9gJdyqaGq4kU2gxj7NnMslQ8FwNr0fKC45BWv8oE4PHW2mrunc+t+4CsL2nhZ3
8q1aWOqyI4bUGVyVtPI4wBYl5Uxga7McKYyQnfxcr8CLSwITLg6kUhToumd/gBBc
rP6+gan+Xqa1HPf1A0ZSctzrTNf/fmzCBPMvz/zVG2YN5Y8Dw9pJT+ewTuJPQ31j
xjRxMkegHbrf5oD3AAREV7tesrtpe8EaePPMpMA3/3NWqORKFaHi9TM2q7DeNIys
pJXsLNwoWFsgOEggmid0u7YHEKQQy0suNVR8EjenqoXjWFxKyfJ5yInSbmFJWpKX
r7bVdTz0+ENwgdmQ/3F0twXKadUve6tMlmOf4+RJKR/CS9YFJJrOdwxGneASs65K
pZjSsGZxs9gMrBFoHoIMNQ/zg3421I2hni+9AsIlpFZ2sazFq5zjwHu371xq6vq1
VuRDVSkpf0utCn0kDIQ9v8rEclIzoV0oyuVDkZmTYh68WJ9ZMIQ7FPGE9TNFTGIT
cVEoK2r1t1Hb3kvhomFNEAH0VzKwOtRywSPFtrTPEEe+9gtS5rR8b86hqAeO3fs4
wu+K0xSzqU0UK6vXR42KyjOdr5N8Rp2wJ+mk6aO/zIO2CzOAUHjjoWRZ7IQM6bM6
OBBx9wdlWZf2eVjKjeMqft9XsxAjQSvKA/bMAkwE+TPyzzfdb6iGLkc0f0RukZnC
wLloH0pVtQWdQQI8sCMaft4MTICyflXHZ5BrONSqKtrR8d/CPRm1U8IH4Iw9HFS3
6pnFJBWAXoXSlkxWLuyiv0Q15JFKX1k8+GBJOMIWZyk0FMrwO7hJS8+DqWgAxuvC
bFO49Pwbj03KGlg2NrJSSyEbHvX5mFU/YTFIK2+UBfKOAPYQM/sP+t4Q0nFj9kjj
knDwElvyu3pEgfTFQxO6ZElyyaczgGCltnZF5mCyYfGgWGpJONciuDqzEx2wDXmz
CNSxdRT9hGorOEjVeIyjdidH/ljWx36FsJBRZ/Hs4qmyiR9OgOdhk2GSDtcCIOux
AKsUd9EeUyn/fwIQxmnc+9Nx03GsVT9W2OtQLS8Op6HDKn2ZTdH9Hrq9oBx9lKZV
HXDtfny6gKHxYSNqxqS66p33U792NpZTys6n5GcvAsNAXZkq1uHQv6DgODzofrLC
O0CyMxuX8vHr1BliNxQaDUFSRzqPadKDj/NmiEYeOje7gY2rRsRT1xKRqIhLLjho
bvHFJ4PUQ0CYreMLI4lXPDNZtvvVDmE0SJtly6i7tCobmzZpIaAxGydqHRzOqUaZ
kIEyKHMiKky2XFLWtUhunzWQvoZLkfcnkA8xhKcYlmJ8odQP4ElaZF1D6oR4v+SX
0KmYXJNb0gl7ohIxBgVqVxRkA2R7T1j6rBhQzhWpKP+jZP3+u0X237xklDPo65bH
3md6x0LvA1qKoAsu7MYmYXIiXN/G71USnV9maCjc9feATRE/Tlaw/9fucD1xCNjy
7Ti6DBEzFJF1l+4DUctDumlyNtM73GObrCLsTOo3FchjZ28xQNN4po7kwto60qOr
w7OlUmmWiVGXGSgCqjluDq+RVOOSt1M6DrYuMd9bEjLW1n0pZBqzx22nZF0+KZfW
zpFausJG5zAl7EPnk7H7MMCgYz3vjOxsH1Ffap8cV6KEo3o6DecghjF49d5HSvD6
TNy/jHMRYWRlUzQlGPUUl5vmJ5e74b4yjo2iTu0mCAQu71Qwy+pYDCPkEHxyB26g
EwSt2ZZk/kY5LApQvXCoiEd9z9NQQvzVso+qq72x/BivJ2V24hj2vFtZdQ3tYiUm
3qXwFYNiDbMYzSwTSCUPtZzwLXKjJeaxRm5fw4Ybw0y9pdPwScGtUWqgrZWScw4G
VWYU5Ka0FOn8Bj96gENBBdZf6KwfT0d6Do7jhQQzGkEIg5VjUP/txFl5KzZLJhUv
GZ3YENxNyHP7Krs40chRReIinN0S7RcDKdZPtmguM3eENmvL6EW0QI/UlmApbgrr
jfRFLxGf3oGwU06OHBtlQf6/0G9LVf5CEs7uzDzToLf45DU+6qjUJSQthXMvZb6S
Uds0itQ4r3f0Un/jrGlX7BijVkuEtQ0FGfLf4AORSInXoR9yj78yWWTfYTHrBrsM
86cR5u8wAXFvRfaQcRZC3A7xG3oEm+L85HT40IJVDBsu7XfQwUBcN19UzJJIPeXU
90QABg9ewipGTT7qndbKXtKIxcjG6CVKzJ/X+ZYdaeSHfoz7ITuc8hiKmkPOPSs2
pzY+uYpkjekdtKu0IZL757zA7Fs8dy1T5q5OaNwjYO0VLGXeBzwndEjw9lFdDNUJ
Eo1JNZwoC4tXd4vJdASvitP2Wc2SC5MGI1DKvUUVp3f3MSZ9Jn3EtYOCOFk2xzSB
YYK17is0lJPnF+lY6+Uzm/WD4eInQsVCgpYsOh8CtvZoTMdJ8rLvFWO6uTOJVIaU
OVmRafjQdLAgQotXMzgF8TlpQSjIhyvcHi9OONZL839nlJRAxOFUFFwgVubPgIw7
ma10NimGn9gdap975lhA/lFIPiAtvPkoHTfJ82mrWWOlyzTA8TEQLHpBFFe7Z6+m
LfaXll67bTCfc+rYXa0e1XGzZLTE3v53/rIu6du1rLwgHtL0THSqj/GVN/+yfvx4
mBpk+lUzm864JHYWA0EXWvhZYJSZHjjf+w0GcjbbLN3CCWFGPBSNmqj4r+V1z2jv
Ge6xNMAz24ozX2w3OGRkS+ieLcR51gfbpsscmXxH9r0HAWmTfeWJ9eUpf5F9rxnS
qFl6K2K1pwQT0y4U3og3Y7iczMAVsbJ9Ji6XdBXLwiS2S/DR7Tuj3bYldxpKreAw
48EKaoxzg+j1hNhMGwT7By9lKNFzLlfAUUt6XKxojRWC0grUx9wL29c8Mybw5ngt
BEK9wscIDbeAlB9p/qk7VF7XLRDZ3iRjur25ql4Gd/5I5rG2lmYdkht0cN61NCae
Wm80X1hetu+6bkq4wQMXrPe78HBLkPCIQiJ1HZBTwg3JUQQKFHhqFrcpu3HWUbfi
+FFFlj3+SkiXv3n/93pnWVGELoeZfIG/kCOuXo8Qw59IcUADcfzf5PDVXQJipGgD
dp8S9/RODflTWGpl6ygJocO04c1q6zKRxlCOyQ48ImPlKVUwWb1XyuCrOIjtUybL
Hx7HOOTh04gxREKjnx95vl+T7e/0p31LT0RprVIt8rd0kKJz4nCqV6Eu5Z+IhJya
NYowNM4n5wuURn4fRImg9/pxVg5opJzNca41waV20nRZ+XlbHbL5X8+wjcMZOBuA
OTKsq4O5/Qz5e1W+cvqzgp9UQBa+W1n2o2c/XbGTlQmAQTQnvfww2rg4GYZkKdLF
XV+TzaLPF40iv+GaxlD/L0hknmZtKZk14BCBxUBd4Olb3QHG5uaQpi20tJ9w1C1r
1CoosCMBUCk5hjFiZ2h0038wOEaVJ1/4jYXVE3m5J1v0Ly4OCvsWjk6pj1r+r1QI
CZW2S5Cu5m5Mt/pewAsy6RcUMqzdk3eWW+y/QhBuiZpxbxh78JBDpfoIFCWz5y3T
J2aGK8yuEj2JM84w/AWNhA==
`protect END_PROTECTED
