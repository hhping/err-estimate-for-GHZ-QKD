`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+xP0KQ+X4iIEH4YoVZGd6wDPn3IVFIJNkHqmhVFoKxPge+KgyXyi13z7pfdOdeD6
UWGz0tqaeDTh7hVieqHm57PdtvrvWu1Zwor4pWYATb4R4zL3OPDai0aGeVqBv6eb
g1c/BA8wIglgL5lHyjp9I+gF6HhkPeM2SPVkQGPQ3/dIDQq+Yb/uGrTInpDcrglU
NutjfsgGJ11uVZeyY1kgRfFbVuGCgP96vPKQNjqvP1tvsC26IqlccXvZY8H0YuH9
TA7WBXfeZA17TaVz/ULI2EoHrpMPWj+8QcIgrg1vyyq0vUayOR+HLBLbAng6iTTU
VWsUroNeD1zzAvTTEI6ymCknhr15nwn3GdvI3Sj+BTIkOZrS84BjjyYwyzx9LuD0
AbgGum1ZL9oIH/97DoyWK8TSVdbFYB6r9byenXqYlr1GM8MesCWEBe5Gquro63eP
j/Vrej+YaPA1UJulV1723xBZIuyax7zDgmk+oOiZzSHsdcEU2a+f6QmR4kFdpeDX
DILxM5V6a7VQmtB4zmHzn70ibx0RecnGh0wezlNxLMAQgKCyIJWCAUYTJQAl4N0k
gc+3BsFsgRRiN1I8BF1yTCeBjQHH1t7nmlxQ6p3IYKSfoNRl16sRFGZ+vgKZXT6C
AXBYXpLvsbMavcBQsM0MF13YwpyKLDqmDDQdltrEHaUjGF5R8HIZ277OicZ5itOP
gLcbAw+imOxeMkTZxXbXMJwI10lhpYABP63VzslZ0EDzVlid0G8TF39aUtI8ruh5
Q5BrC0/4OUimxBUNcMNF4CXvnVYFqeAGXB3V16XI8a4nbWbJdpRxp0dM/oj3BllR
jxOlf+DDC70Ljc2TcOv9uy9tO74jc13Di5Nq1tqboYKVANDcyrLe7yq6kV2YbGhv
7zMO2HkuctRlASfWNXHGuK5JACcF5ZYQ7MNpQ54S1hCt30VtzfWTXfqmN1ojXbJ4
FRfAg+enk/X4owUjSiUNBwLOL36mVBJP6aZ4K6pFzcb7DMil1vI23zMATvdF1wlV
m9h7CZoD9WTZgE9aAmTKHpZSu7PXKGhdhKuS5xw5RQJULSTxmljMeP7m2qLQ83f5
zu5C+sCBoKA4IQ5I3wMsqOwgbqpSyH4bvvWgIJ4O7eoXyhqFpR46ANfid+VIHyjG
wjEXt84jd7J3xUXk9Btcjz5vyS3C4XBsdt/jA/UepCiTNril7VdS/ia2mj3WGN1v
Itx2khWIH1f67Bv6c9i8Gc0HdyDwhGEW/QyOe2h+Ttt+b4APw1M+Gm0GAr57sSL5
RZ09SM6yFi/cjz8XU9158WEJIwOHsp1+sbp3rswbW8F+kLGeCkzQcJMXN4H7swgp
+RwtNV3xaHsnSdVr/YI4qt4sD39cMi2YUFD3PXFZoJ4wSnYhMhLcEG06/JZcfdjd
X4LhLRfyB/e1EgpFPXMUbtq9sh8Nlr0wsEd8+uBQ+iGSLR8qvNUf1GZ7SoohYp5I
fJv5Rd6/EElh/nmA/HgreE7eAn0X3y0G+mPsuR7HKVcfdgvdAcjT331o4PUf6fXf
nDpq7Zzfv/o6YJ30xHlhnhci33HnDR5xlIYbOSrNH14=
`protect END_PROTECTED
