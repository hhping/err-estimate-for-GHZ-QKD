`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
parJFt9bRffdvCmC0mdZSDpjSHz/nbCgDIRSHPg9bhY0qsmtII5bnQ05PGDOWNgo
eGCLKuuPiQKOBrGgE4IUQXglTt+nJAefkOxVzwactiXFB8HiAoiLE49omBfeWGAR
V8nBkvzkD9RTlXGcEjjAL2lU648Vj9JKVAXRhTmgBHV61lP/RRZDI/CDEkdpkuN1
I9UxN9aeTvUBjEULOLoyNIjevMYPIZBW4YdPcoJWqtNxjp67PtmiFeFAIkfBVQzW
gDDNiqwK1cLkZHJy9S6EZf1U9q1y+p7ERHvklddVtQ3+KUdMJbDcgt6FXmk3B+mQ
3iJqR/FZRy2UH0k8fekuG9/TTZGz6KCgXvtBH22reW6mg1d3YMzi6QRaJ3haXvDj
g+PtV8yZzr5uxXfW7U0HeE33JeeuHYbo0QZb63Nyx2xUgY5ZF4biFdQGdwqYgdfR
crW8wiVuEH06HMF9EfpY9bxAuBN1Ly+QvujkvkAQHdk+rcGVuQNI+nP9BPCqYDMg
TiUv+oQ5+oW7gTmp/vbJqV46lVVYfFxtUOrN9knQdX0QLNLRMOBarPwNF3iU2PXF
zXl3KaC1AKLeE6QuRL1FPAOvAmoxbPFZdzSWB1mWSiAoENIBPU1M2BUpiXo/pVuN
`protect END_PROTECTED
