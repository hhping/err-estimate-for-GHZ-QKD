`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
poqazRNIwEMCiJ/LXYc7VvhRYhf14fXFquMC9hrvHGzKnpzaOL1opQ+2Ia2ksbin
MV+3Uc0S7dw4XzdBWQ1l7aF0HcMoN2Cih5HvzKyN+4CmRqKJ5jrVDklF+ySvjBmT
GgIOMNekkA0oldGvtInaimBZx428nxgY5YxK09AhSivvP0yKRjrag9lReG3DbWhE
+zfalk4wGB9vWWmGbl56liHC4KVbFAXJWrbph12w22pE42TMJ7DP4C9uOVapA4U1
D79auavzS+JMHuKZ4JGNGdT1b9FTiJenHSCEoXiL2WRU6TM0TAAwPVFhy3H0Dj4W
08EYTPlMOWvsMxB90abiBRsS6TGAPLnXNQuWtczcexzqE1830kSuNJ7DxYmo6s/Y
H3b9DzQXRmtiIFMmpdBtCpMGPrFXCO2UyFfOwfPpdHUnoK3yZeuuwlHVAIq1lR4+
VEGhGubfVycpl/VdZCrcv9PvjL1o/oQF0DTOAPq5H9f/8LwEoknUwy6Fuoab0hdf
UXQzWK8Vm09pMim0vfqeCQw6zAaTYJUbpSUlEkRFZkbDYYtQ4AZxbNXe4xRFpF5g
MjA6f5W+BShiYv+2iDnazN68T8y8WESaJrd+z3lR1FfpPXn0W2mxRYNDilCnz8ps
0fMPQeB+cUz9pxSuqa/uPMHZetFtRxceWYSkLBbb/5KHkFwMwkqg4UKwk1uLARJe
apX7BUJrhuk9grJ58CT/YKYnOhcHRBoYp10tuUap1Dk+e2enw4GkeHa3TsSiNFLv
4/NYmNDxRgVcU9yAMn34bhk2pClWIqothw7vS/7mmGFRWU0J9OByDsrGxAxrKSBX
hA1vlEU7jEJUXUXPfiCcA0VzHQh/P0lXIK2YzDMfnkfflOVqDT5tZravRwA5thpl
XSOJGvi4BqlqwzcFq3Qtc6lpNRYWpbz6QWz3SqBk7Nl6i46BQjTjnc44vuA3lHUj
1G3zGqYPpZvogLmQVUdzOXejFCiunan9MzjE7We1omVpX67/JHNE8XBiKSO0kMJH
ongWj79ycqwU+jg9QhXQcDIxMZWHvPAjWoA49CB9fylxRIvVHqnXjJawNEjMhfo8
u9Q6NUAoiWwxA0pGPMr5HGURzth+XUkWO2B/in0iTOOe80+4fABPHRBUHWyl6Htr
7k1R1aaXTQjBmtMK5pMkxlU6e6J+BdL1ZsuTfmHDC2xMra23mqPD6kQa7IkMJRfP
u3pawFPLYgMboXcwuEm1zwv0Fi3NMigEBTcKRuCyqG/DzHbUdNv15+/hvxrDEBg1
vMz2oEhfxrDOjJ/LOeix2yI9zvVAMnX4LnDlCxNd7nuqVM1OjRHrjzdoXMe5tik5
Y5YTt78Xe2vgKf5DEcO+/txwiHWZWOTEAdHwSNNsVxHrwb229sRCnJLGn5wHmuI0
MR9Qy6TBoEd6LqnkAVcLc1uht+14XbPBj0ClVlQ8QnHfmMtYmpKzIy5g4XlcWzgy
AfCcK4KBP48vx1KmdrXU9G0NYNnURQMYv31qFwx0peD1VeCbJjQLOVKRys9lukir
+B3R4vXglxBeov+oIAgv3GlWXdVyd0u29JLd+NFZ0GnOSRVp4sftxIJSXuGDk4FA
/8Va3FQ0yNacpF2hkDllJWWBuZKJxqCz1lidDr9iI+fyAbkKmAEdsfsHchRXsN3m
trdNeMXJprl6QxKNlDi6yQOW9jYP49h/ENTfUqv05ZxK9qeMfxXhj8sD/rlURwfY
JRD6w/i0jP6v3JpGukH2Vr3ZZfFa7C6X+W4y3z2jN6Gz1DNztR3MAIQOmm9IfOMr
wHIvPPMshr4Kj+chhsxtyyrX7w2zgG+jsLd9v7kEzORwc1gEiQ+0h0ckcy4r4MAu
OXytMQVgv/C+cH4rwNT75/aSOGS/dtropeiBu8h4mYTlXdOsmXoiE5VA+kQ7lc7W
akPIpDDNBsJnZryAigHFnwZvc5vaBJ/1FR9rbm+2PKPFNsnuRvyRq2nIyY5VuqZl
Oa8fuDWsPY05S4FDQ2eB5BIhRjMMoMDPjXA/yDjyEaIyMLgA+WDyCnPjNx+XtLDr
zdEFeXd98wLtzb2EeCRU8FKqPRAwgtk51HcIajKGB4C3+ZonBkg1qPOjTY/z3gfD
01lwznUV/C2CtCozpg+zu2klyttE/C91zxW8SIUyQHT6cVxyvEIHaXeCgCSIke/a
OBawWe6+3XCnmsSTG6oa2thpl1BM2cTUQ6KWMYWfDngeWsn+LOWb4rMZsnVFGRC4
pSVwUPNo1S/dZ7cLkJLlRA0L3wg/AF4n6SmLSTq4adY=
`protect END_PROTECTED
