`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8oKa3Ks5DUGi4euw3jQu5pfqDBz26+vmsSrwOxYkyXFM+tMQhQ9LSmPZznTQXxT1
+C489yYPRM0S4rBkQfamJzEQKa3RLS6SlLr51Kw4ld1Y7u/hemF5WJjhs5w7EDSi
AlH9dDL6s576NeIVWNiGx0R5wf18nA6exMhRQC9wwajhwL86WbRSX0pAqcE8FG+z
yqs7sF1ix2UH+44dZe9LLclGEBqmLmCRvtonBvzggZnzEK6W1e6myoXRQe/yvIEZ
jvu6yxlyoMqCRUoMY5wESVCEbYcLXr5dl1Cy4sn3KlD+Vy//avWBT4W5tofw2z6A
MV4JQAa9NKfyMPjGSUaie2mpQbPHzsiRzQKmljjERgbhQlPOzdv4b8czEjXIJyQw
qAtDGH3ZqLjGpcPBgx7ecj9yWlAzUJEHhvN/k7V60aVNppgZU+nuB6QpHQNBAZMA
79VuUjxtNt4Q51/XlBLGGBqreW3GIXIxwrXbWlbXj37nZWk/KKBD73UqkYC7jqSE
tH/G15MvEbYcVnT+ZSF3cXiau1mH+bt9hdjD1W8xNHEf7qB/dqhLAr75MNnzfUS1
YMj1s/MMAZFbPNvut4RQTcqUnxIWVO7JfMWgP9/RLJeYmamkOY3xNVxADwyoGoTA
sesFSAFAovfvh7MPMjQMWGFuwoIlJsSlu6uEfx4Vf8JXzAQbpzoH+EAxfEpjieoV
Ji4jLDfgW96BDjdRi/mo7cy2M6yJa8qnLZVQ1ZUaDZPbkkfuiRdJrQ9MCm8Cji4e
wGW2c/BP0pCInNsyzhhU6BprwOrGAQPMcp5J+7GZd6n7roNpYejQsNhKdF8bLYCh
ervFxkoDNvvJMAn1x/O9KAYkXZOzhOZM6NuS1d+zI+O32YkEHun6AfK95UQxpT+E
7h/+VCnWwWtFqTJ6YoC35QC+CWbJ4hGPwpfbhEBKsBpsxxPveXLaDM3EjpOEhKAa
V/mdDzklXfF5aptxhktj4DCk6tGOUusQIpjRe8k9Vn3dcj8K+CkkEJR1g7p6lDDz
XVhvhSdKgYqdXTPQKEITWc3Cx/Rc8E2xX7RylVkFpF0t0/XOMvw+4W2W4bA71ECl
ZPzx9mZ7PsiK4AhqmouLDCvFTGrzmgFMDQ74Vq4waDB9JcHsEp8C7rTBkUCJVyGx
qgvFPCAC3Xdcuv0DIedNxEMUx2nkmwPldvvYf4zpbMJ1wF2NqVCLkhzjXPjzXOe6
uHl9EEF7aKyWDrY2Gbj+eY7ZK4/bX7N7eqkEUfjZ7CuKKdhOYfOmPa/Oe9MVGegG
k+aMl/Y3HVfVH/EWZ+CsNoyRSYdLqUdJvhqLZXUal+f4NKFrXF5fIfrbdNWaTkhb
95phLGZLpOlWhOC5ke8QzM8dZSPnJbRdPlr2AVHFz7Bor1DFpc+OqK9h4hd9YgI+
YCGxsBC3S+ZgNep7vIjG9Ckf/eai9l8FpcszbTo5prVgMfJ/3/2GnzRJEPU3h2Rt
7Yr6zt3n4JfPr/c5mXhUj073ekMJsIYSU7yxiHdmKfGzT56RtgQ47ViL3E1FPv50
jUBJpKuzm4Cv/LU3goapIONK0mvJdpR3FdY4XKJxYNilcl8XlUg9WBb3b3V312bz
8zat/SRQZkBW0FkyBo4MtBJkZzut1zjc1OvCx1FbdaElYCCRcln/tQNuDG7M/ra8
GVCbEQV34h/yvDQd+fXpXXgpa3Z1xyrvsa6eKwfA6ZHAX4+Ej4ekDnmNwe9epZv5
gMBpH2s/pjcx1Pfgt1J6e2aBR6sYbkJB4WqMTWSU8VSJXPz8TQdTC7tttDTdvrZq
Ac4boP242SXoT5heouXuEBFJzdXdFvey42Jg5S1FrCAf3l2VgTJGABaT1rQ7zmDM
qj2Hcv3fW8N7WRfH+LHaaHEtn9PPoa4l8c+B2attoHr/2er2+QEg7e6PD6EWWPTi
pMy+7REn8KPsAZxZ41Gzpb7hae9W1XdRykjC1RYdmtQekP8fpSG75w7ssrvKjlPI
5npqAqEuvbZGdp2xI6qJYkidkdODUDGhtU3pTLPFWxyHDWibhT47VxVU8l/15eYK
AQ+3jZnDofRBCKkuPxSqn776SFHjnWAryLkJZRIu3p1ZG4jfl4CeXmjpSWyfcySd
Osembdk7ptHqmhza6pcYG6mxKAqhg7/hHKFmzVsWR5RFH+qXl5/Nrx/egrY+/5n7
quGsRiDc+wS65r5tOOChgYojgTU889kg0KmhVFxZx0Xr5IkaZ6LctD/OHA7aRyb4
0ZMA9QePt2tZaHVWKDhdjCQhSwg+l0MUMuBS5CXvvBUOeHSCimse8/Ultkw+KAC0
RWfJrwXuGXX/uoIoFp3X5vXdrQuwmyn9p+yi+c4Ju/kXGPCQCRi2gTBxgnnw77kk
Xd1dsGGGzGXL/kLHHfqVMm6wVhYxCaGWLgrql4h0kAmBrXaOskS1QvlF9icYk5fm
9sVqmC661Y7YpB831pCTJj077pMHUeFr4wPcYnYmo5PAVhIFCBJqgvY8Vns7bM8d
o9VXFONuaN3QhZM4qinu/b5RgmXJkhHUv7pHkZedwa7+e3vamuBOfd1vkmwbQZ48
F35gLxKJ2lGHCW1pGxGOePQFCB632hI73/CVONltIVKIh0UwuKR2tCzEu/wNqkKo
YAZ1ziN4VYNDuCWP3MvdrickGeVIysEkPppccBbfNKya1THYPaIRaF40U1ltv+0p
xWqkFKaU7NEmVMxpcom1X8D95IrgJ+0f1bTzeqz2Iuq4NvtqPiQRr7Kxr3bHO2Fb
UdJrgBqeT7vtIrR7Y2azFSYE3V5UPTxxxDj1T04RO8osTE1lkPT6aRcL7knP+4sk
5RqCl4oeeO6nVItNdFluOlYP5fEp46Sbc+mmtHvyFhEslDDUx7UtqoUpdqQrEFO/
oAQWRujfVXZQDY7AVjbAvWAEKmoMI5VmdEoEn5e3J5oCO0hO4xhs5PDENxP8yr16
94gBQbGq123tWkUMj7gnmvONLKLskSMaTRUr+mys62fZKeTFxbDLZPH19eNA1p4w
muFj94GjZjYvIz8jI8tfMlu3BaJOhMIRJasVKJDV8X4WotIdwywGrHLfIY5UbExE
1p1RRqwoi13ta5WdV221iTUs+fX8IMb4t5YgeXSzWy+TJ+VOKHYEBeoWXhOybGe1
V309SNiXnoqQUIRIi3QqsVqFFSvpwBYWJ/o1uzVVxV3YrVuVobZpxfPEyrq83qD4
nE+ZDSuY5QXutCfat185204llx8rOmt7O3V+JhzcusFzT5Xel2ir0qXB5hJV/UJB
x3SwuzYkdIi7Vqug0hasxz85C26TW8Sl/CYnBmD0QLD8f6a22YmtrJIyfmDK29Nf
B6Ze3wWJ3nv0J+y1Z0zcisC5ZS+cQ1/4JQqZ+GaZzdlTpurNJHOCXW07mQMPY1LZ
6nxbgT9sepdIZDqOZTtRH1JhvHaOi6wU/D8uHjnX12B++NBL6MNks7fbnhhdiSZA
Fj2RUoA7U5ie4JRdM4LXeFfflg1kyqm7gRhue+zs4E7DlcNduxBr+McMXoxaE6Hu
Um99jsUYOUF9F/QDEPKVAAYM6J97TvhZb9A5LMj6bfgPXStalVZAHyqCKLD1GJf9
oFrurJRrUj0TpJKe9R9O0ziNAuZEmaA2SyRm5nIH5DV3ucg+zXjYwbFB7kQMqg0R
MooRS/hDYv30hICduggTSpXER33kzQbmiDMpj1DQCYwv1HkScW+Sn+idYAgUCX8c
XZuXiiuPCQlA4djcUttQqK77FMEe13ilAQVFrLTOBIz9UwLKMhSDo/dYqHhnfjr6
GNLpZngQhQAE0qHRsYLLHplnbf2kzZARBB3G/Hl3pjcIuMzlDiZDG7BJs0LS7Cwz
mVUVCy4h8k7MFsX8cfbkIbxfL0rabqh7UGr2+hFo4vInhFrKOS87Vp2jl3/YC2TE
O6vvNLqWY888fGmvjAgui8qDNL9oJ51KHyjGTF5xHx+0yMcB/jOuTWr5TDb6J3qT
yR1CYUyFYRmwsqaesPXkJcG6iSdRSvi8LNtKwSJ7hoo+8x7oW08mb8OMJukwp9by
vaLoZzD1Be9cRsEEHnswKNVWjSWXIwof0aqae6jVlX30hsI3YODmVOwZM96/Zdnv
IjE08wT1+VsnBRxgSUmLn6B0UcLw6FN0u7Zfc0UnExAU2RAyuAqeOUfeUbjJsjh0
P6AhBVIm/oUUlJ2k4Jzlz372IJHVDcRX/2G8n8KT+3ukiF1PptnNU71fBhuuGdmb
Z/OTrFpPmAVYsdXildIYWf/QwgOn4y5qBSAa5MFxdNVNKyOGzJ/Y7/LSvGfSTrXp
2SRp6NHS5w/Tw5+kFg2VHwjhCKqo1yOMIlKBIGSsYuSeznAyYKt8swn29OaGb1Ul
TZX+ZY33q8kcbulRR/nVgMGD9hABxQzAboKMpyBM36Pv9/QixkPawp5yYHaeeEaV
lKw7YsJ7pDHvPrKeRmxTRTe++2G0FpNKXR7RC+5DnOc0Zrl8OO80YLlg7odiadFC
nE2ilmpNup9VgPWqr5nw/+CoADIh4NRwzxJhRIdTr5DxsOYMT31ENg+Rv46pu1pL
b0f5F2yaR2kTR3DT/HauvgaGFqaA6N7XmMQxhd2LlB1Rlaj6lx0qwd08UKU4FUXo
2fT3w+wbtCYebLWjXy/5UvfsTe4ViVjCZCbX3513aoEAHBKdQ+kW4H3EimH7g47V
WjycDoCU/RMrfwUpYjBe1k1+Sub8Hl8iZcAY3CiI2St/1KXMflOZJgC76Yahuipj
8/Y1NGMCzVu4Os9dy9DoLWGFfcrzR38cNUQ9FzhUKPtZ7nK9lsMscvO+S3D3yxl3
5Tktdy50MbaEfhckHukxtrknHP1WrnQMSzyPVyoP0sZYYQjETA2/Fj0uCHcifH2r
1rnH8ur2Vomuaw3fPO60g2MT247cesIszKsviC4G8gZoC8G1+iS1qo5YP7yE0ad8
BdHOTVLJVMikV/U4R3KsOlrwRs/Uuv5kzqQdEoZxA/X+5qMC8md0pVONAgAORyDy
W+oL4d9B91VNW+cItJjbwGtWerYdkIPnvh+jY3baV+4VoZW4p8maIZ5SW0CSmdd+
lsvpa3LHeUX+jCrrkCfjF1ax4qgW4fgD7JQH0JR/WJQEsAa2ae0h+mwk4X1leodH
1qogQEfobcZFxLX0PL0XdggisJLXk3tZCaw0FHgptzx4b6Ad5m48/nJeSw7RANhx
UPClrm9nXKSHby5ZouIdoNFTMpaFSmSR0dYPsPf58s5HjInTaA6z5FITHvUXOkeH
bxX2B6Zd+PsTSN5dmynpQhwC6bhj8srGRstiPcQtsvBPOX/h0h4MtVpEszzM7Fsm
cNbJdEfPlHMzDYZ0EvT5mlrEDdY9rJ9JRxSfNcfWJaETqwcNqQWhEHbz3LN1YK7U
JFcBa4SzYK5WlfcAecdQCpOh1/7vlVm0KgxbYLFC8/xOpMjgq7sVjP7xpnFgQqqh
q1Rdv6zFQxqU94MbWWBlfE7imxUh5560yG9c69Ua+ZVsDB5xqUpM6kTHkNLQOqne
yk406AYBiy1m82d4p+zdWdJjWCmyqVj1URnGRg7pwjd6FIrggO/hzhKHALNxH9ci
44o4FVx34T1YOU76FYUFPRpJ+zYcx8rYp8wuD5LfIlcmFCaLgNi8RAg1khhgfayq
yDpxHp4vBuf5n2XRwIGPIvQvijyIgkgNloJf3us9MpuAO3Ytf2I22wrdHCaBHFu0
PoqJNBdS2MF1hFdjUizj4M6hPbH5MraHdj33Dj975gg3iI9GOD45geZ0LL35BdCZ
Xyb6fY3d419WtiZ4sreXrGlCIg/OuMTVRSdtTcrkdPTL6J9+kV/+1TswDym9wJhZ
+W9YN1NiI9HIJnTqLprQY44BmhZyYh3sC9ib3l+3VzW5lKF+4fK+YheRUXBJCoob
pXVC4Z1oSmZQiQAjIoTOYyJaxmfB63MqQX9wFnnJuI7f/aDe2RHeFwfW/y/VKKaG
zJqtdzlh9yZRcwIVd97bVapyG6p1Q2UdcqVtqLkGJv1h2hechXr7aehvPSSZMRNi
4PHi0lRlHqUYdAcQcUcA6DHPhgnwuU0BwCtQyq2nNMhJkcap/WN1YsuhBq5nsCJT
UUx8Q4O2/tJnJ5i4W7htm7nN9QbmbYqqrXI92FyIXa+lp1XDcI4jqbrgbIXQwkgm
j8wzADydaaHp3tOONXGsYY2G1xZdc6WwgxJro/gdb54M0EISLv8t2P1pRM1MEA3H
3PK3kTBe46hWsy+opOoL8GsQTPDySsNP9Rv0VxU2Yrzxs6TIzvtnFmpb96tUkA5w
Q5ABW4H45eSnm5LXLCMVLA3D7cTprzJuPAeAZkgRB5mbQGGqyG5nKDZMuEQ+YGYm
6yD+g96Kq311vXgvx4YJblOta8SyuOM4cJlVtH31AjLGkDqWS8pdsyTrt/A+M4Qp
eAIzkFgkHA+AQhtrsH4iVnf3O/YkB4BCseoi/DeVms5qMlnVCEp/nUw878QpUMe4
N4cx/69OUZ5lAHAHs5ETQwPn5EDCjvvYDE/5Q5vugBBWEherVJoRf13iyEaRrsGC
eFUVZhiYa9E1v3dmEYt4W5SW6MOSMrwWkR7O28kQgsMwBLFlnNnTkcs+psNiVu4+
z0ofeAYfaDZ950GE7h5Fo2p2+Be8RR8/Yf5wdwWoEmiXApbK+OWbauW+gmJ5o1ql
XBWFoFu6E2awDpCaDqT2ElUKLcWLyUoM2a2/LRzrYhNIWjDSLotZhu6M/p5Ced/U
8ryuIO0bhJdgwIbjLrZgqfLWtiIl+N7uzr8uAEgXyqu46YwnUx+TgTQgCGhIQWQy
Mwx0etoexy2fg+t4WRTKP02CC3gJOsQuFDsEqU0hBTrfvvFQ/5q6YTn2sAjswWla
Xu7aBWyAnS9ZoHVI2P6l7J91SUB2Ff0dL29kYiSGEzyeC9oXotlOkPH571ovn9uj
gBVckpfNICfcnSaL/HqwD6W2NVhCTfIgs1s8PVB0feRDVrZuPeSzcUMqhAd6P0TJ
wWItAMz1mXo2oX0ON6RYZqdMRjZVzIPrX0Yy3bhOz7GeJv5FCSkS5Xcd9+jUenYE
aNVZaTEdhwmSpeHMGFWv2oV4u68+OUnfhRaYkZnpKUXsiC0rV/VVRjMXPsEQzv02
P0pPkw8Y1MkIAAsVb7/Z8J5kXt1505ktuo3SXdNxLK14QWEirkLYwZtATWlaMYw8
7Mr6tWhLIa6RCm1L2ONkz1P0Uj3DzWQmg12bLuvxxu2Nnxsrmy9s+4Clo4KMo2QS
WKNhZXG5Bojiv70gQkkY+3W3nNup5Ewwe2D5CzrFtKT5P2pN4BdDsthJk5Y7Tpof
boiQ25YnNMD3IFe4HoxW1GHR06c35PwnMZibNmLcCeQ/yoxCJR5qxkMW8nufjbuW
KTptAFZGLtWAK/o76W3fyVpPAhR0Gb7zf8H81WhTdYrsfuVvD4mPVtr0Yj73emFh
1nSZlZISxf/YQql8ZIdjJmkPZoMuK9lYZhQS4XBIaCXs5Jp6UEV5m+ZD5/Fvry5r
AYqL6G5hGVg4qBeEameuio2WyPM0ChNfWG5q1y6dhHCc0PBZ2g4VOYofsSVRA8Hu
2oGWY5gtj4VLYqHZtyPcsS5ilxur1xJmQeaTVxqqN4vyIz4+EpgJJ+HTByIkpnf1
Zc9Ql+IPIsHXN6qhRgwAAMqi1CNwBYrVJiNOGoIyf2p9PjivPEPh/knfOazS5Ab9
iAdvJr64KDlJm/8FqBrAb8ajxxztXFzLxPprAPS7wws3QyDN/ZPL43E7AG9z41at
AcQJGlfEKHphykEzU4pxE8foYcRjLtejCXnm3UO89HovbSN47iPKNogmDX3Wz4Mc
6B18s4Rhc8JRftEOEMLRYudBPC9eliteDTLkBXGj2Xw7Z0shjeI7obm13/9S4sYu
MuNwqJuaI5jxB4cgSeeanWxO8mZBi6T1mxOSRaHa7zD+mkQeFeKwS+l/W6p38l7O
IlIhsFT3F1L2ovJZHUopZHYSs/9QSemIssWKiWQFYT80JGDepO9xJ6KztCK2gwnG
xeG9v88SPMea+8u2bT2s7KzUZkQbsLqdKY+9/DN4RKC764CTGSFa+deK2ZkqvPfM
1TlPzprnfuxmPn4MiguIXK8m7AjSpbmTdWYO/dvAw4uvXVbjfaPxwE++ah2G/ocz
voc64bVmZCRahmwyvMeZGUpdEaJYLcLrroL3qER0Ptxahs/UM9Gv01YLiQFmvpnL
uYtRIQGfVtoelS3hSplvbZ+2a4iygubscXNoMCls5sE9FoQlGE2iyL0fgsZtDGK9
0JbmGoLO3er4afqpB6aunt5aclrqxNBULfm/ADhjUPG6C1noELeatcG+0fEsG7GA
FwkXTiduTNJ/ayXOp5Wpor3wlezj0ApYRmGs1V1Jl3MfKEVa+RI0RemAA025dqMZ
69FEh7oXNpfuXpe8P7+sC4cEKWFiHI7i62ayxY4tHr80R5yLjvmXdW1bdiAx5HuL
8HIJNgXJiCpUmnuwxK4OUfGZ4wRStsKntlgPZTyVxSWMbs7dN1u3RSxatMLWDdpB
65ZgglIxNBnpypFrhpTjRqFcBvCrlAmqw0bLZZucm/J6cFMRPxH7U1ciXw/D4lWS
SZqd1ww80F/JYirXJPGhwAH6CVstjWcHx4hPgzVxFPI5n0gS9kx+4tHE51iA4FoX
3JpnaOf+mWlzTP5X7pt8Od6NbH8vr56W3f6MbVk9UkAQZj1aIMxduhOtleyV5u1x
uPdCqNdDFssO2ggNxNxJ/fcy+u0wyCPIcWYc0IDxXzMVzZX8XKkf13CyZ4UoWibz
Asi/2DX1GWIPyr5nHKW8eWizmUzpEMUbZKQlnevu7bAHFXyDp46b3SjGiSvP4cgU
I41dwZOLrnLn6Fy/F3KMe+NmEXu4MypUngrscWcCqHOmFneN2LVxIsLqIf/adQ0+
zn7s3I/BwM+BqCiv8X6MNJx2D1vU1wKIdGdK8v6gJFX3E031EQUMI+uJC/SMIvim
Ee34dq1/FwYKGqUcEIKQ8wYS5E/fsHEZ2DVhSebw07H/KD7SKLuWNPrxFgTGcL+b
sTsxgY48tpXTMl1IzMCMCQ==
`protect END_PROTECTED
