`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nFY+2fVUZfecjYH6mKP7/rIW4Ye7PlkEbgOFjFKq5McNtrQLT5yEwp+5gNefIPEe
6bx98YGHlbM2wpeNobsuHeqTfOdwakRuy7z9O+ZvZAp+oxAugCwHaG3Ucfc4AlSg
cc1xAtcmkfKxOwzjsi5tdMeDYy1/oW5ufCXC2telQYKTqZYj3bPZglf4ORXdee9S
/d2LZoTOQmLESb9yq0TQUAg/cD0ANzy/CDIPkaSbnpLlmezfRC0MF1DLGfFUCmiW
GQnK109Dc1kNe6mWjmU0bnMqg88YuzKKT+Cb6Z43hgAD8+DSFX1+8IkRaT2OtZYh
h6JJMVX5XhR0L6I33+AcjSgM8DzFzWsPzZGw8LghANWnWqCr0sBsVwh1YsZs6nPQ
9bluWd3nMg/djbJBrQPOmVLbBc2df9Ur4eGae6yD4bR9tYJYIPu7Z8fhyTgimaIL
2clb+4lE0I/wCErsZxjXd2m3hnKPJz4I8tRlfY58foRtmeQFE+J+cQvsFTGOkN4s
UdXZFPBfycNpFeHDFhxS/+H54lDDd9B90IixSpPHkNLJZggnT9XKqX60chwQ74cS
Ar7fg2LecZSfiANzC6XGgK79cRNiZnBtIu7KiRFddo+Pl09I6Kyi4cPJ0bV+o9GN
Xy4gTeYgPrkSetawm5BaqZei8UAll/suqKfrlvGKszIRjBpO34WJgpH/+0T0qWoq
PBJzD/+//h8I5PzuUChYM9dmpoke0q6kBIkSqF92JdGd9nvR946TWZV5yxNz4970
5l/J3StP6MyoaQTpklgjCftlu4sfknhK1L/WMQqPjXwr1iR0F9shjq/tLxU/z6hf
5eXdy3b6Gqn4WCE4NV6f0KHuAlk1o6uqfae32QaeSBTeSRQ/clwtpwn/9y0h384f
H1plt1O2FqPkhPfhv9U8CNM/iCM7wUSitFiO512gaoA2Se1IzlRMOzHgj8iOTJqn
aqirmmLtBuvEAMegwnrBna+CNhYbYaZHdW65gHbe94YktoL/Url70bjGYJM+yZri
1KhYhEY5tCsyjh+OZXOWEk8AvVXsZi/hRiaZ3+bF8eUSbnWt47h2p2ltb84vJdXv
2gOVVsk//fAqbaVVu1aXXFu8tizgt/xKVZQbmFcPXiag0/ZRCl0inAswWz04lQvW
ELosfCTQUjpmAeDZHtgA0csJ+xjiqD+jdYVEm79Mhrccdzu4ON+FsRP19hLftY0v
94tOaxq6ZAhoS65E1f6W0a4EVW4nsDcOd/hpzSw2/yPtT3ZiICDt/DAECFA7YJAy
ubae0g/uNAIVcaoxPnRrhifcnqIL8Lppy870Rjb6GQZX9+QV/ERIBwuhcl2pgCo7
I5E4julciuOVAeOfTnMENVf+BdxfNHtgKR1xR7fRYDe6IMSrbfjvRkzdLjMecmAm
CfL1QDwQqTa4VWdt2zJf230xA+CLgsR8dMKJULbTMBBkeUjp0ozvPl1otywTvJW2
FyQj6BZUMZ1g3FHL/XJnhOl3O7aYGqHzWFh6BZI47HPMPvRfJf7QcTIBz87BaXoB
+Tkd/kd5/Ih3NEPbnWgMPy8OE80wcquvCq/U2DdnO4mLjLAFQ1c19Z4/XIgQQ/kx
WeOmvex4Gg1K4VKvBINSPg4kgKFmWT7CtjdjN+tianVVExBYLS5CNT/YxaJgc7NL
lMSEGEDOr0QeENf0yUYH3gvDB4jgOk8be6rwiQPuu7XwGU01ohQnrdJbSom+gC0D
HsqZq9ZYXWVtyJSy9OZhLAnVIePeJIWDrwZkaMEnzjElDG7htoQLqUKRl6YC8Bh0
ZDDb/5kblcFJbvwlmUW6aR9FH0vHwxESSNTYrm1W8pQlLqt38YVXzkTdu9naDATk
GAEyWZH75BPFvc0eVFjLUlXJS4nWduZBDiO1uw4a4ruApk1KsZDfQ0cl3mvi7dEG
xpfUDPSzp0De8+J2dZvtMGmLA22F9dkutvrnZZqUxEEiUVZi6Vy+V5JZv5zgHvjs
LDdiFSQWkzl2F8zeXJOor/hEntgvsIaXpdKjTMeTt39eKvjqmLIFyvIwwWP1W/M1
HHHdl3QbcCfd3La9KixEzPDFnUbtgU6/NcIITJHjg7E8Jr9G0TYAe4hP4WTI0qiA
p2S1nnOzAxOuAmdikHUAZUrJGE9hzS7KM6mMbPC2ZBcztTzvIWfCPK2IzmxtQmvm
tTWrrlkry8Eg4gxksuhV1PfDhsuaEANY1g4JyJgCqb5bmjbEMXvmNl/WQu3O5Ajo
gBZNflSIRiCbjFQR9SiTMXwX4iH4jHcFPlUdOEc8obI5gCgTb31XHsmHCJtRr+M5
hpLtnERt5AheG3S+06FMa9Kkb8l+ilh39GUISlzYbIpqxhHMURb4FLEAYndvMSGA
bMa82iH8aQc4vUTEkdFo7CjywdiVmZ85SR+srhCB8vyvjsiwhF3aa1M/hR/oRT5h
NW7i6JlaPFSRhifrT2gEg3PEDgRtctZl5WxcmUMYO29EcNVnHNYh0Da2uxidHmLT
nUZeANbOH7SUZsUdO6MYbe889fcVinijsqvGni4MqsY/vcmonTa13OWPHaWR4iMf
qEkqncSxZQX7V2oVcYKdJwjbej6REwp/XkNmV1arhIz+lj7oAZq3wFugDGjUA9XO
rmZzpwWLZGhqnsneKnmkFWdDhK0OteyVKR80nl1yFnupApxQSG0CyA5jIJuxgO5+
ImbONQ3UKsYdgzoGhXOrytYn7/Glz1DUJ026L41rnMbPXG/qt49OOTAJCdd43nwr
8Mts9vj/qJ7Q/jv6//2Tv5G6OMYUE9ynkHIqJ121HVyN2XEz+qSdoPgM/amwmzQK
bgxG0W9EXLiVfbxEPya1J1gGjwLNJp6kRnk4fEbpVtWI77BX+Y9pV72falXR/kI2
pf43ZhHHS8DVNAv9uLOCvfcGmnQERWC6KOX1bH71D/LqLexfPHHFFI+NyDbRNusM
D0XhRXfwHZrS9Vn0GuayjM4g00a+b9PV6ysc+9b/zzLstKajuYAgJw/GOmRwDuEF
l8RpfziM4U4F8Se37jTV8PvSoGzmgHbbN7fJFuyWFkY7B5Y+jLCir3ASCM/U9iOq
zoU3SopedU6nWMF132FMdcQaKEoOh8jq6bfchkojE+C4tWDBxblaeUAbtAlV4eiP
MOAAKf5MXqJS5DfC8WR1fIamLjKfPhICh60WbNEulbjgZrtKJnbCY56Vh2nsgyky
wQw3dGMn9YiDwqSPqarUQHX60fA7UJc766Jldb+U/yfa2OKkusmJrzieB8sqXH/j
ay8VkBYndTmjLeWJDsBu2NDF7NnnpxL+TYvG9j+zhl/700edvO6HSTpv3EAJB94g
xUWIj6CbQe4q54YmO8o9//8Gsik6k8yPYXJAFi8gCux1nApecoSeUh69EeXPGIpj
gpLhf/W4QXjM6N0AejUVsdaHOebGAoaDRqAp9GFr3KLzMuk1rnwpFuSL2S8oBX6L
rNq6VXr7tpsBJwmjyWKvNmnz+64zKPYHkzCFagsZDknZaWC3hnDU7ZRWEtw/4kyc
8wTvTWUV1c+MSZY6Axm7Eu0DIUvwZlODuBU5qlfL4dLaJ7hC8vcQiI+RspUKuKbh
ENU8ajKTci6dO1/13UbOcbW1YYljazvFS+sB/SZ0q3+78GuXCKhbEOflUhHVsQD0
OIqp1e6de1tQG3Dqdfzi2oSOwBMztB+nYAZKpHBiAOj2n8toRNWo0clNIijRPzrr
cQTxtwuNrqFVaugyGfpRmQdipHy9wANmEgJOL6swU0cF+ZcC8f3LWUZ+pSQwdA2o
5275aM32LM2qe1J8Btaowq5s1d85j7X6/rMwebvdi52jtjHDWgw1a3ifP5W8H93l
Nn/kfPzc1s2koiozAlQhvXn9NuC0XzKBLOhUX3HAsfGoOzhXVnX2KUw4VNpyI/qM
yScmbyL6HjTMI7eG3fEq3h8PNwYpzG5VF9Xsuf2+ZEYs2N6B+0E2GIUEdJ2Qyh/u
L/lm7VV6ZO22bSjqauwkVfAr3WFV5tHm8MnvWrWx0Z0PXjbC1gnjzFDcVbkEXsPy
qs0A2bwczkk3iE1lS+VqiWm5jw1xLDNZ+duYZyL02GTUXMRyp+ODuGxkJCxCSePt
VQScIXT18EkAduLFf6eqWTilokcP25iy5QO1uAifFbq5BQjHahfOqCIb4xbj2rnF
W37Y+nuOPFqbqpQPIPfCO04Keyg/Bpsz31sQBOBq8nlMRH/uisNJ2buK4NLqYr6o
Ym0iUVFMl1iP3nOcQqOMjrVwJpJPrLOJo8MemED4xIXHWiaqqLgS6ccPtBUA5mwp
rXjup7V5F9KXehR8f9bF613AFuhzOhjJffA/jjlZf2HeU3PqgndhAb85X5zXjmR2
pz5PQ7zX10MysLh/VEWhJtn+cm2KBqafglMH0nYGjRpy3y1C6BrxO3OcGLVZbpNi
ftHkY082BBLV/dR4MlNAtqLj11tog5M/Yen1BpJV8SUsBqlTs63D4+V+gqy8rN7y
cE/VvSR4tXykrz+YY8udBtaWhaFprJebTatQUmmOEj8Cj+d/7LwU3p+NxoPxJMv2
5NtrT29qhrtiQKni6sYwX+irezfmLvYVnwlS5I+KE8fi+GMyXcodrTObYb0JO1Rb
3H/XPyPiB0BHxVcHE4/6hFyy2QUpVwqsg0K21BKoQaeSSg7frYWBSpU3fMBGaRBx
1HyA+YMh+9cocos1Bviem6bldjIkYkbmb1sasYohLzbLqYmD4tI/+afYgObHtR2y
cNGQFalyjEd9sFNJS7FQFcvLw5XaOBjAb3jY357XrY/bf3tOfCDzOGCY5gGK0myp
DnV8c1HAHvbCXy97xq02E2x+z8upcwKWrvOSHZY5ZawsUvBp4ZiROyXMh5d2mEG5
945NDHHPGX9AY8apfKKstWwhhj84ZN+OOWRaU2V/evlrTF6te2uTfKvgA3xhSY/T
NcehJjRgBzkkgDC8EdFXH1jQ0e3ExbhMqrqoHcBz5CrIuqE9sr5LpWk7DWswbD7h
QjgzeloSbnEYKNqjPIhK9MrH5vAdubo3u/lNky8Ubl7/UNihKeRjK1NwiXmRSiQb
qdKazeQD+Mq8EZ6MGPbmz4f2UFiM/wgyQxjDjtmUXmtBELmDtAtrbC+5UVcLUZdG
Etj4q+tjcaTaTY2FMZmp4hJ5z9oa72+x9rz3Fmz6fjx2jwqJvhFASzOVhGLQQU88
KO1DEIQcmW2VW82Aa5wSGHr3k4oyZfkwY5n6ENPxG6rm1ZoXni2Y4RNrC+yM46Nd
woMhqv3LxotIL/M4dFxR8Lu89+u7aiWshuOi+LSCp24zaf4zgjTOqK64BwS7sbCh
KSkalX0ZpbmSthTZ0uymsD/2H2O0Ttw+1+rF5GojH8HfsHlVmRyoWsbovWyQ2GRH
qa5Z2oMAyg5vF1K0ZBC4mJcuUAWIdi1ZjbvorxLl659qYg4Wz+/pXcdYK7Z0j1Lm
juB5S+m5YIrEOb7DByemCNB7sJYNhFRZ54STUNHR7dLK8GBLfiBrojA7OvuOVp01
/G/gTkIRMU+fKP5pdc7ETTMqWdacFwWHJv6WaX6gFsLBrBBBYbXH+lMdg9pFNPyd
FKFQLz1nuNUT9iTqM11pAGRqxXgx1vyXBjvtJ4QzI1UsQh1TNBrJn869+rhlKOJs
YS0NnF+P2IMyycX7SdxGkHnttuVKBnKf1QTLxw68egtWntGQm+oUaik0nB8/jnL/
fzSp0aejuqF4gdF8s86IK/bRg+k/FIN+baFrp1VdWrXKWFPARqJi4qkH4qzx6Zdb
4qHiHlVMKSEOM+Kl1y3xCcMQ9HNp+fMi+rgft5DHCAUkzqHdCD+DEFUB30XR//ZJ
omjhjxbsUJafBfEjaQdGxLGdRmsbkkJTCrEN16PPc2t8vsiiC/hLq5Na47XUypFq
gEeTTwP7stENNSGLa/biRPeOU5uBGrl1fMvLs4fBRwXykcZCI8s0QNlSQBO84NtH
eE/s4sYKED5dSSgRhI/RdOzWmVgYXGo8gsuD7/bXXCg6HTBJQ07XA8sBUVuc+IIG
vBq2U/j0crULy+CXbapnq+LMP3JgwdBbl744vgC4dQjMnkFgbtTJMWBm1B8VpVUa
vlwni7FiNm2TR43SUqyoOk9F03FaTMnLs35lpMmQx/7RXMDIJ+3d50KjKdVuGGzf
xpzuswn2aBopKPFhUiX+7BswLw1gAcPDJHyasOdkDBtuavvsYbfRubA8lHhGcIY7
ffSGCVgVVROSVQdWyoA3ApHPG1if38Qu7QE8lXoInPAI0fOQel+8HQdXPIbploBm
so5x8+qXn2co1b9iuwnBc6F2l2X0xWtkRLxaJgJ6W1CmcuqFd2AVvG1VBPuNGaYw
zfI7L8QxoE3sdwGoTcdIGpzw3bUTAWGyZXior658VlY5zRKO+2iV9ZTPrZyD6FCc
Qx3F5+1Wb518TH9d7697yvzbXGDUENDadQ9MeNzztgoy2oKXv3hfBPpdHQ18HQRG
YNwz+G10HYMIXIqPXCViuJWPnkEqHZ6hYhwGd4IIB3UIrVc+lnweizFd3NTwBmYu
mz8Qqv5pTe60X/yP5gLJZgdtCdQmsPL/e9C1B8GOIITeLjyjZ4PYG192TUA0eeQD
9icXfiVssKwAovzDuq72ihM4DsvNKCmUBl4wUp+Y2D96wwaTQCbZfW1+Kk4eLzuv
j5938DhZOn7YNNImBOSg7NVkG836WNfG0II8e3GRQwDBOFkAtBXgk3r5NGhu2apx
MwH1sbyyCPsxfNeldvR+39VUznmlDagplJR5C0rm4Hwd9oMsXFyuLuEzLW+oaoHc
O+WHa+0U+QDKoPG7hP3tmhjdfCH0MPYWmK1saCmYxnbS/jHFZq3rFBBw+ROxCyth
He51mpz9MdXDwkaXZJ49zdniKJxPdQVfxRnGeH5Vh8gth09zcgnEgj9UVNfVKX6M
ZUyPpPEttSyFMo3Nb5VoqUdDtR7YU/7Dhw+2b0rQtzkoiAe2MEzLM6QaRN4sVnzT
EnDdSoscFOWc+3Uotj1xDGLme2abeGKQROpH03mQdTGtwI2jfHDlFv5jt6fIbhPo
8G1jpsosmjwQtK0GkFOMIQdR8CDgGTkfGq/whs7nGVBnecid/6oUVUY+dylBS3iT
KjfvGE88LXAQdeTA2NbPM8SMwaQP/MoGWFIWmHyrp/DMJcEte7MxjTaVCOyYWZN5
/eWSNeq0DDENrTFWdSt1yHybAn+PDhCqWhvzwffebduA4ek1cQNlJ9IVELgTpW4R
sPpE/JPbXiSyBrsYC/xF+BxvwWxSA6r7KNAoJ0N4L0OMHLQSjCY5W7kDwgYPVrzg
PqgZO7rONoqop25+pg6ah5bCxAv+xOE+X5Ez+eo/IoMQIBL9DNolJk8DfKcDXpkq
LalaMrbWHh0KaBT8FdqdRy8ccV8oyddjY17wzCZX1CvV0GEQdUtBwasxNZ+SJlPL
LkMLj+0/zBtpHe0au+wZuUPBn3iY14dOHK4/7WTlmo5SI/G4lgDF3jzRLliKUWPR
32Nd39gyL42C65kvBpuZIRcNfzsKliXUeqaXtMrvAHri+n4qjzQCX/wpn5nRtiyM
z1JVULNQumTrOoJtbVPaeeac28X59S8/W3EQkhSzCg+7SA4thw3TZsPujKIv4pUw
ew4FkwQFFH7bFMiM5Q4EYU9lbCevnkLu6AwyqGyHdrIgjzEiAwdkVzZ/ArxWiU7W
qjqDiIfF3b1OueSKWgbqFMK48ARhLJCXet2qsbQECfRQJsSJ4T0oeOEVzAoM62oM
bSW3ljg48fudElyBcJ/CWcFvsgJFpelGXHAx9hQnc0TdkeCpGI7JtEGAVR65Prjv
mLSRsYAn792PUxtC3wVADm5U9wBBTPmwhXqzAy1IYJysieygcUmxQPNiMx+nroBO
W3UqtWBQObCupXjf2ohHv7uHMEzQ1V64d9cfpbytEPtj5e/xg45l9IRc+9VkkZr3
4NW00dhU+7GibfXVI0Plqn6quzY7Rs1ABtFgD/QMhGwk6XclGLxVy9J5MuVU34vg
fAsNhFm2EwaWYAm/QyLc2eHPR/eujlb/MM2HTTowBuuuVpjTMAI5L7eTJOxqQdZF
Uvde6qFYPdBBxYps+KLLhzz8ju2KcR0nPZHtqysNjsb5GKsHjZbmBabYo3SB31rU
TDUXW3nlPqZbsuonTfC615gA7nE9nhaoQymGj41XdaHi+8fre/EQcSIDA1Ibp55i
5lbxkTipf+ijKB0iCVJaERyBFOd0910tQ37mRuBk+siUOyoUU5ixTEWR2IAK91as
hu2zxmy8bzFf0OamUqAUReu3rcpnqBOawXL5XRJ8TO7iot9Nkbkb2D1QKxqArUUY
ITpymYxVeoAFY1dP7x9MZCzHzG9xU4Zs6YV+kYjlzSSdScuduunPpZKBJ8BaCnOP
5y5rg7AcmC1gNyigpIgMguWciAI8bPpz24tOBfvXzPOAGWc2SLNpne5PTmxCzlmg
w4pWtPY4Aw7G4RZBRbwMlOuJcKvnnMaJ9KM+SIb1mjtwyaJehdJt90CTA0tQY6VO
CbSSLtjAi5R0zIrCG3lUJC/+MzWj0i1eqHmJA8XlzssnDGV1jbcFNW2u0pZmT8u1
PuPmbnmsXeOBP6zzv4D7xXXCh9RXo6B3xPPzczDl5j7U8K2sRvmbc0bSYztQMKub
6eVsGdiPgB3UIj9vCJmTuUMnVR8yJter3hMY1qYAhzeZvFneddcHVBWmXfpCGF4e
5A5JU2FZJ7RDcdVndjZ8AxDxJRSqmaJu+PRJpJdeZqvdi2L6x3Hu8y4BKNe+q8NG
yITVrzzmLMOfhsWxFW/QxI8dAio1zQZiYwIX/pQfz8bfWDG0JHx23P1EprBZuv6v
WfOmanO+fOPu8SBZjU3Z3TKsa10+5yOfjNEwcgKMC1ljhJVCpTxwWtxrw4zovyuC
PC6np7XkCatHl0RTHHNeZyrEx7nFiunb/LiEeVybvkuCMu0HGtG+1uuE9BGeHjCm
uEJrQESRqLSxIh85lfsD/PbArGs5/TFuWckn82IpcLlCUoNTO1nbuJa0ypjFnDGF
U+Rb/8jfU6dAG2e6YUeCigmynqd1ooJvg8sESHbIJM8IV70GcwKmNgoW2jHs//Xd
L3YAigl1kUWTV2QWnVDkczV79xpfFUXd9+7GQGIlBCtaldQ00i4/UgMFBL6a0y4X
GdSS3CzWxwf/e/w8XweQi0gzD7gGR0IqoSToosj2aYTLSxFzZPNGWZY0Xb2sRFbm
nPEtc5esBFyZ7rBnsPOdvPAWmyZ3ka9+90ieNcv9IbyL2uiq1cBKdXdToM1BPTtG
oBeyePRHrhrMad9puhndbAEBT6N9k/St5TIWwLxI+KILglzGfdq8s9ZhRz3YFLHa
dcvQEYIzBVihwxl91PvUJx34YN2XIafN+35j+QdF22o0c7pN3RiZMgUGwDUKlklH
p/EFUcEbqyyn2rZTkdPy80O2++Dn13zJ0x3DhWXjugsrm+EjxRNNATnv9lkGnxc/
sVqODk6Y2zlMXvFuwbE/S1CBSYvSrJnd8xWDCgmz5qnrTs4keZuN8iKikhwFW94E
HRTQnJlEQ65BuYSxPbbSDH7KdIAvMuGxeCT2ey96fspGisVh22qy6/3XVCU9ZfxK
1ljsV9InV7+QVs6nlgJ5BYj+bgLIu1UZyGo6ZH8GqLWgb6DhyJQoeLnvIkrgjc/L
UQK0yW5yHQhPDMm7I4wzzhfQ4QtKL+s8Dj24rM2WYCd/48o64yb4tGpbRPGS2liB
C0sCrypclBpBjAn957J8Sg2D0ltMnzp8/jlbN7jZpAmwZDJSF0+of9stRi0ZwkG2
fdVOuaw+xs/tZmIppRxcjzDbtOA8tpFPhvXyZhY7Gu9BEbHp4TR2EPsB3dg5JNDI
wPaDyfCmZ1o7+ZxNKobEiLY/fSBiDq/Xj97Co4O4Pa/MQHyuQAyge7zWpBE4RuHE
qXMaJ35h0r35dxGcSLPfcJ5kdCKf0Y3jwJ19DtJ3WFkEEm5EvYUH5e0g0ti1e7gf
sE5uZ41DCFHAGSHZYTBzaIAi2+reO/NeMhAENjKGihMFZCU3v+EK9pUIFbh7b4VN
zJB/pFCFUdumAXeIzoG8vQTtSSNuUcz5BsFTAlV6lOoadM3SSyTPqd16aL7yuLOY
6i/gKToVdiFff8H41oKiA36F6g2aBU6K/gAQvXggD2oT/lpcEHUg/Mx9PPax4gSE
OC/8laiVPNEbECKIyviAU7BM+vj5BNPVCDdpzW21sQvoQH4CEWIwVMMWLDxng3Bl
KZO0kd8t/f80lxrSl/39eZ4jxAjXNj9OitOu1MoLg2kqBrLH4EGXHfMpGIBQBawa
6rBhho+KAbVQdsl4njuv9y0B04oulP04qTE9IWeeXqyzYp6ZIMQsJtsosoSN+j8C
/G+ylR3JrrRFDZTXCNvBHt4GUTePlp/sQl7ubNqtdURjPuDNQBkPFFbh6afMPYMM
BUaZRTcOnd1gqn6/KbezKMWb5jflct3nMX0uH/rZ25az36Xptjjo/D1cudiRpHAt
NMoaK3yynYVNO1qAeO85NFmRlK7jkUUO/ek3uam7z1ekTB4rBkE40VAx1t/BtRWb
zLDuQ9kscx1GPjIFq1fnt+Frpgn0y9AJK0p1ljTDGkAW1yvihTJD3Pg5nF3wwpub
EGsNXr/ASXvBercCNOtwRNcyl4jw6OZtoaHbNdG5+Gy0ZbnecDIDCksQKFwBSqRu
JUdiuE+YjmPiiNTZXRg27RKiUb7YM/hJW6UpcTNJvvATFq3TjJpUDD/PKHn72atl
NfMZ5M3vfN6Pjt33KGZbrHA+W6CyIDYSAwqQZtqV+RUARDSzcCRNdAQ/SyF2fPS6
0QywX2tCWjjV90n/ju8wc+Mo3GAzB6mnZD95xRvMi76yHH3bCQjZuDSvO65crahJ
fdX8EcEgj9hJkgwGIPGrSdKwCtn9XieObuzWJdm5tEN/+r8B0b6qii3ZMWTdu66k
0cqNKPw8ISn8AETdzFzhJpZcmCS4OkuetS8TDAvknbsGo3bVWD9+1/5Abc0rgjRW
heGPS1/93zZNgJofbYi3Vf+XntFnuuLz6ocb1AF3pxG4KiaaEJdYUjJuuRj4VOEu
GqPt/aVmMfB7AR89NKKHD/NjlDFlBAJDcmKWrz5XV9Ig6nlDRpTWAREs3GW8FpbK
DOtevrgjLNXMzE2aERdubQjAYgaGy5AJA6b5BfMTXICMwISluyB8GtoXDWjV/wXB
ZubPXneR6j8WL99KhZieoYmI3DDn5KtGAAcCPX+ltb+sNNG21r/zda1PlQv5ZmLM
2LGBS3itp5E0IvLcenYlYEN8t+ELkHH4dzJP96IM1Jhwh77eoim1om0RKkzsIqXf
c8ViodJsSKV948aj/Snjb5XDtECwaMUJYi6ECY/vCO9910xFdOAsNtyK+OTODRh5
F8W9BKdCB8k+KvrYNw8gConDV4KiyNaZcehuFYBCeLMW6mKHhpTr5rrFfej5kdtd
qJH5RxiUfPQb7ppMUOLZqH9qoenB6J4QWaEoOtORpUfsPKhRTkZte8UF7POuR/tq
UMORehOJHzy0HkO0qViz91UBKB1RKtJKnBOkPo9HcZRAMSrM4pfyCmHcKW1JmN88
DJLQwkzDKxOQhKG3M46LdD9ByPSDDxxQ/PtkNQBhI3rqejnCYr/n4utpuNqGR0dH
axIVmxsRv6/9ZrNc4DKkyPT1yzIUo1MFYmfk8C5iGXet0hCnJ0AHcIlUigT+q5+v
gOVVKTUPA1I8jaW4T4AbePM867eI+KXD/qtzdAMzTd/DkdMSH5OCWsJh9cBm6XoH
o1966OLaC8LSCGU/oBM5l7foacNtK4trdv0MFspgtPAu3Orv0DV6iav+pw43DQYf
JV2kMv6qMtam43b4zFIUnmDqJgyWxaOLdR8Xl6iO1lUUkwybnoecoRhmRU4jBtvF
RXFcmT9Tk4t3vo2r0fI6QD9h3O2W6LmdJ9YOSbWbXZWCDNxYWc5ZhebD7CMg9szd
niywnAtcOvk/qH02ijlaMbv5Q/OxbWea/XeMtIE1H6KAuTiPeWpSB7sodN/lHPkw
g4WTL+gqM9GgMVulKldLDLEsT2BpIZjqXWWdvio1xSFBwRLE+CxLV/fG3hsUaPCs
+VswivSb/qLtHjHqPxroMTUPFmcJKWmjFXI9PCoBmv6dqw01KF320WgtuO0h48DL
+gviQ6nNJGjmoEODLQsfls7afsGDnvQxNJw2FJ1nU53FfCd+sN7SORRI1+6FgrQR
L9R8GcaFfHVuX41OyzlGmTO9+A33+zhU0RqEa7iw7rPSpmSZ0Hzlw8ViAXUYepXk
p8X/ghX/RYHE6+NHkaRrp3cuZiJo57oir9oljIz3A222KkWHVE3jVSLTK1eYCpgC
LGKLPCJgZywsirKprL13tB5T+CbDeW7oEaB5lRrjJeA0n2Hv9Zgrx0s3Ss5bI8k0
H/TIaOGxzUYffqWsR6x02giJkByvob750T+sP9Jx4AYD2VD6Jbcsil953PDDHCMx
Xxc41Pa+f85lq+a1mtWAo8gDbZxROg4wdjmwpVIXnBheu+fLkAaJxjfghd/0UlzC
vaRaJXTf5RB8VRM4AjNtpUz4GFKENzp9rC8kmWB3TgVzJYuPz2QGxGpPW5Lqd9fa
6jSmZwjOOGJ+jI8RaieFEP8z34WTxQHxW6fenthsKTFe6Q437SAZVPDj6/5f1tR9
UOuuolIzBg6LxqK0PccDkKiPJvQl7tTZ35OgJwHAPjAMFDvFXkzFt0TPeiHYAtvJ
/yf7j8D0nm5+XqKWkPrBXaigELEXqbsIUZZMbEZajbugsvACpnZQVoqBTd0HrEeN
iHifW1YDcJ+DEr4jU2+p18fQAlLO2lFEYGpu3mrYiXm4fnwl5ds3eQYbU44LXFJV
8Sh8cix8lCbQkj5/HWHCrTCNuBKr8X6Ep1YWgESWlE9GqMkxBRGqaDWAcr/Ahbv6
7J0MVJfcndLWe8njrwG8Jnc01811g1/fzgp3am5+FAc6P5toab+KCr3crtq/8NK3
e3aVbpdLJtSAgwem73CWDVqf4yGta6kVt+8H6+kSe8Nehi5touLaKqar3INy+acL
jUmiA5yPhEMEimHwsRw1aAKFSoTuri7gNzg9aCIDdUaAyQ1K3oRf0bl1MYXlIg8s
IqlMhHyNhurIoiLjuxWE2UjhBVPG5CyypeUko6NXZTjlH4HHu5hGyiJPxTE3g/p8
223R14r9CVwUTbg4qoFXpXLwFvBRz7Y+PjppqCCDrifdbZfU8yQ4XZM2D4itsUVE
ULaz0ZUDXt1XPYFFyxpHORsNz55vEZoyn0MkUj+0L0Yf3WNAAbvfy8NY3U8ZfEJh
Q7nyythWBvlAH63Y+WHI9WzWbpWrBfxZiNYCZDxTxov3m69Thij6O5xCpNWYVlJH
0Mduht+/hQQejqPmOIaIEftesx9Tn0xom1jVNPO0hhAx/Gwl6vzISFeIcj9JIOn/
X4FmvzZNeRgv/F2emJvDgK2OOAIDcES7bEC/NhSTHsHRCvMFg736sJ96PnpX07ez
mGMZdQOy4L+OVrTUvQV3gJvc4QSJLUedjmM/DJxWtflF5hvpp4qZnBDs8b4oFTf+
BT9Tsfb7s4zM1wCfyU/KJTxqTYb8AkS5AoxPoHdjxTg4vYd9DRzIO3z0A3c6QWjl
YQl67VecPoQYyyKYPuN4sBLl8opZR7ljmg40xHoEY/skbdE8a/bNQfV9ScDHXYGH
rbaFk5AjedVw8MhsBmX22XhJdEOn/j8dwRpAuMfo5K/NEZ9Jupk2bveZtriRaoP8
EptGYp5PwCgFN2jABgL0hT/mp/FORh44lcuzs+eJimcxDLN6alFyROVESiqLzxQr
+VS2mbhumJs+ZKqur2HGwGf38Ob5QUxvPLF8eponjfp90rKTOlH4LFS/jk1IigzW
GpRPyyIKia7T9+H4rI1Nx0lYmQGCR9gKpfDG6Az4RHRGFf+oGod1RuSNu6pLGZhL
j5dNnwkZYYjOjin2CBXize3lcBhIT+y1OIj8MTPobl8PEVTrUiV1XFi4E3YoTGXN
jQHZwhyHN1JXGjn5SazNLACtmQKXS65SR+y4bGcABEOFH/1QdVts+qXyO7MKXwN/
ZuD0+cxsUVlFJGOLQex1fWBZZS7VFuDdIcRxw3oDEq068pK8fmxJ/de/fX+LC2OR
u95T0DTcMjwXb7lbBSL5dgugXgKjz1xh1WHFt4NIFdEAYKaUwL8YoCn5clQUxBWz
4fVVBAMXHVowjSd/nJwynhwMtJxaa0GXm6EfDOb9KB1gQiQv3IIqf6C9Yk+bPDjM
W5IR+rnT7C6CbgHb2EY6jKJlFBD4halPuMNAhk0oJTq/kOy6Kunkt+sMfAsE4Wqc
Y/lEynVLFUbmjfCLAS4iRR1OFMvdgffnmZOBorB4smIvx/2vr2xhhFymeC32VsAt
aPfipLzxgKi5/w0HoaLUAgviHOwHfd/jgeXNGBAGaFmGDO22+wsVQi6WIPAymxpc
k3TlY8ucVo6mdJNvL6Sn9GSSx62RpeG195wdiJsKX2LWv+gYnZX8vWjIB7KCFf9I
lD7zQJDcQeu+6Mkem05Ni7xTMJZfpiuzJrTFtDRfGp4DMzUsmKFmDR54OK7MV+S/
q0BK+3PwF8AW0oxulzA4qfadQPc6BynLy/kOZVllxIez56euWqHYqHQySDmYBuKq
4r/3THL1O/0CzwTLfzMDskufm3DSlUAdD/R4seyldxwOazkMv3zYfmogjMPXgEDx
d/+tNTPVVFX9GIykHJJuCuXAKAwfqvt2G/yrp+mey3JevcFjH1piLxVjJQVGDhdx
FswNg+ki64SCf2kU2rHIkIm2X83ioduU+iK1oTNYf5thayLatQ7UT93UlYDc6ptF
Z8dTNaJmuVxcZVVaBKLb0hckwYY6aOuqO4VGF1Jfdd/QB6O8394yyoRi3v/MZiS0
aWlLu54cT38YT8lszSKt7f6hdybJUVRS2Cayr0XKy2kV24pwdND00rc27G8QM1DB
vVszZfb66GeFMsVvgQwuhAb/4fy/U2l2pbOwPzRb29BFRbhY4tANzI05NTCAFim+
jSTDbxBydsPX8N6sBOV+XeIzmY4HP/Dfvt1KZn1XmnNQcuAk3OmQyV71URz+ZCLa
mVUv2GpW8PYMiUpMLUL4fQNIRdmqrmBGE7pnOPdbtwzCEQPqKZIWyK3s4ug3YbVF
CLPH+3WfCUUQKk8dDz7zTsTv8XYoBKAl4DmrTlSu8znSfbbYuQrokL0gvvGh6uVF
s4iXLAeJq41kKDOQ4oXJ1YfQ3+le2ICj2znEDvgUy0qb871OjIyXNZB8HN/f7Bv6
LqHquNAlDTTIL3E9vRvwmZHKCFQtT63LhAagUcOWYwJcFRscP2d0o16ukapl7tJ2
HeORoYlbnwXKnM7Iimq/np/t04Gtf0ak6FC2+zeoZ858tv4h2BQDBQfkjGFhwWP5
4WwYJizv/4RcqjZoVM3s3qKKkHhiwFdEY5Nfiuwzz3a8g4BJAA99bkl/nyfY0oRW
4q4whL8umlSC56ZxfycK8eZJJZKlOavXMvfiC/ivdYg9Tj8Bsc+U6zYVMMGiL/n/
6FQtERlsZGd6Jh8lqf5af+Rhne32sWGYQ5+m/a5Yx13wRwX8F0RFuYEOUNb/UERo
PlbzhmR9PZx48Q8areWHADjaZ2tC5cXyJWHAiUKMgsgT39DYZT7tmNmoAjWdmCDC
ZIFwdgFbIOr9vqG8hVX/UhTz28a9z233y0oU4w4liTqgHNOzLQbxK5AqLVc5eArm
m58Z2eSdqSY8MIHshDYpl1k0q38juUwxIcl1iEcYJyaQgQHX9mYDSEJBZp5XwK9J
7xI4sDJhxs61MTAK1NFuHWweFlG0kIjUBNj1efNdfKX6CxDl58WBtjCafevf2kor
bL2SPOUcaA8dXrVSRA4DfInIlemJsqcOIqmGVbZ9tPmkBxaiDvNNJVrph/Uq7W50
DqBpxS4NyZcn2RyWzpRzY8y4N7UIbkk0tKtYGIcEPsOTO+TjvLfZHvHsR2YQGfGT
/rcqOUBVQ+lKOAbvx0an40hTfETAZbqYn5hevpYw4k6PcYKS+8u1FxOf5bf72Oxu
6rZytC9TAiwP7Pe0OL+uTU/r+fK0FfrUGctejzHQAWAe36DGHwsbiao5SJt8I+RE
b/h8qE8wCtcQHGId6aNc5mrsQEgTmV7SGzxmRrGF6TZRilb+fOMYJf+acocgJCfr
WcgcJ/Y0+99zAzQhxy+oL3zY0mxDmrBk/nf+Uo/Qwo0pdo2GwK7aKB4rVdbr5a1N
dyjHGg/a1h7BHv/hOdN+eL7X9J3Xkpzpkc7ODW3RdYBzNuCb0acy/Vpj9axzUx7S
cOox+Fg6INmJtrs/YAj+zQtk9IlaYLAHiI0A6k4wi0rN+U4WEz0PTWc2wz7TTJWM
zm8L+GBwd6fitub288mLYp9z7OYb6sCDUDsQIv6V0VS+kHFJlSTRknC9d3TJ6u5a
HEPKS643WkUvpPQmxTcdfR12mUjC75lMb7DqgQmegFouPCBbEIlFnka43H3QVNOV
jZqUctJ4PJOKHAyQwi7mg0M2t6WGbLrBtvFE/VyyjHW99mItHn7YlIbKaIMPC1Ug
wnV4df/miVHfN8S2MHATikeHZeEjU9bl51eKEbOEIX0whm73GuaD+ccRVyK0nZ6N
JETLA52kQ8m//QRMfVs5mSZSPOQ3t3K0Gb01uUWAxkRW2EmQzwsJ0UVW5XvTWY2I
Hbdq9v2k6Mr+3juuz/RP4SItJmdSzk9337VE28oDbvFkwU0TFzV1cWBggXpeEvp/
AOes3uAr66qwWk/Uzxb9bgAcK1y8hfC1CdG3O3nQmcLQEFONO73DKN5H10finzsI
8T3i8z3fcrB+kGrrYcO6fO6VVHEaCopwM29eIC8ehmB+TRBUqzBnyc6on7A/BMex
NnoGG/S9KlgS23LxE0AkjnGqt+gdfd+GgVli+oQOwlQy5EggR5E7A8iCuiMOPHAL
xYU9lnvxUtVdY64594VYtksKSPDrmOKkqjurZZLfKbhzLjPVMc+vyeTFZzS4zGQ4
WCHu2ifyIAY0h4Gj27Aq0QlM7qFzc5P94x/N0QpNEathDppwUKEEiWgJweSN3LlM
9z+/ipflVxVcD9KImwUPNWEHBa24+WuPPNCXuYZhonkTQoAWVBH1a6qNfDBL0cOk
isny7Uyl/2FFfGi0JtlOTqZ0FPXbp5jqxI4Aij50rNiuaq2xNPb1q3CC0axkcNLF
70mfC2yuVCo5ew+8J7k9E9K7Byq3XyXBgvxQVLpRBbvIo16Hi7me6X0AXDdBEyeL
JBK7SeJrFhZsysRjVUkuknIOFOKMzivJz9mlrQVrLmRqEC2xArnSuRAgRjwqHJt3
U6UJDf6IjfIte3fvVahj8ZQgIV/j6KdwhFfNx5EQdH6hc+Y8BtIPcPcxHpmMwKpP
u+GCQeDhzdGllOpzwLy8qcfmstIZLM2afTG8vOwR6xfFCKmWNxQ8gb8yLwBw3V6f
274Ncv2tkl2UWav8DBjEs9ryD+F+YQrPPmVPp16XB3/7wO1lr+xraSYh9E8EFI7B
rOlkPir6+eN7Hkdx+uTyf7MJU9b0Wb5e61X2kuZIKkeiojuoA0lAJFTBDeutL1wk
IVhrh7RSJlzt+OQIpPl7lxM/h3V6Tgm7Nm28qyGKdmpxuxLJQMtqkCWy+DCIQMn/
pTmBnxT0/YNHUE4HS8GAGzTjYTJ/SIaDkDgxsUBTNVToyVSAXxfQWymajJzX2B1a
x2tMem0DU5ZrtHgdWoO9WbuV5Ny5TQJmK96Eyeuf90t8tQQ3s4WKkUX2bVNY3QfW
rjGJ/9PU1Sj77ws4aAqkoR2DxjRnNYunVfpJeuSFpzm3vr5byXTIn2zctJl028Zv
L4mxBNGvzieGv2ppWjTevfDbZy6eY95iP6+8Z0SetixfJSAQcRIHh4YNM9yZCg+N
ey2qmlIF4Tbvn1L3ZoIkNyrOe9KrfIl1NTV4au/eE1NGPqs8ZGRSJgz8+nOoEIgB
NLOpQaElCaaEb23QC2Wr/nD2VVgU5185foFLFsb9NS0Zv15ES2WNW0TtCmutvhS4
CsMmj1UxwUiJVGOvZ9dQSbHNiGnujp/6IizkRAAHzuIkPlDQkC+5snXibj0rUN4H
QKv58/6BvCwNNXbaylK/oX8QQ4xDB/jWB1D9vMh4BCLW5hHw13/Ts70kARY+uum5
JTk1fF/bTpT2g/bOJ+hhQEXKp6rdDBeNLtrWoFD7SAhnQRrjvK8M3NamLTryqtyu
3oiLrzwWVjmPBlQR0wjsj8gG3VTUk8vA2yt0smKqG1vuEi4tFMQFEuJZrxRg4bbp
ikQ99KR53LK8dVvEEe2iVqKXSLTZUFT3PdPo90smoilGpJ6dVow5UT4o4NK27OK1
uu86OAMBhGT4OWE/DeOfLyYdRgJFnO5/f0IeurNQsR4ZesDW8NBkBLDu4fgBLlJD
w4B1vnidiPhj0/4QKfF/4rKCgGNM+56TE23L8hRdNcABBEU9kxLB9RyfN0zjKYmS
/kXe8Gw7By5OtdnS4jJXVbNAh2BGvdwx3KL4HcIGQMl9W/6GOk8PKn2vbor84XBP
tv4gTiTt4jEyRu746xXChQ42M71boZ9R12irtCdWdRd+PXIPsWU74zaEeVu5BIdz
+38/1S5oaEy2Lwta9zVq2f9oetP9RqDeu4WgWZGrdl7I0XR2UPYLhB+sqOvihD6y
W09aGxPPpAumZIZ6/8ooN5PqoS5MYWNZ8N9tWZsl5zTp9cvwEHsf532mf+fuShw+
4QMrxlHLDDIXPbYl2FNAhzB3zNO6GLVUletl2rAADNxk+09gbdSampv4rV1Z4Y0y
P/Ydp/Xgc9HCC/wYb1wQWpSo6OHT8TiWmh7UFyyEPDt+RN3ve9pyf6WL07zne9KT
0VfcAhtPmrBtRYVfZ1+SA/z+n+v2hwLsRIZqmU68FIxdvZNjtlaeAomNoevuzQvl
5ltUwSM+C0UIZP9C8jRpFFICa7J9UGngOGYuMWdrEUU4/9A1WDOopcYyRE9x6LAT
JSjVjgkFuKgGdkJ0sHs4AM85HYYDHYFv4SgacH8SzkGcRm7ywjuhcf+BDN8y11O+
YZfu6jjCmOPjBfkuKnZSxpD3eodebYXs1RXu1NOByUNn/ITmzomzSLdS+nhrPtgE
yoYgo8Ds9qJUVtjnv/Ob9Xqlo6whFw3JB6HqZZjzKvsEyhPTUnNqN8Ywem9zOLAo
ziaCh1GmOPO31AxtF6j7Op/iEpkslE2ufd+qUIPg01jUIE3UbDYK8aDHhAdrEkH/
pxG43WtF1oSEzaOuWXdXB2vqq+VRwPbChdldZLBYi1uosHc3KqwLyYCBKE8P5zDj
x9f+zgNtDhnC/qBTWtJAjeXh+PvbJ/qJ37vcEdiZtfldMWfwPO6bocfqummU2nXm
wZ60g+Z6uUGppD6XsVJs6hw1BkpGJjN5fw5TzbuGo7MavncdbZ7rGHRmqvoLhfBz
Jt7umsQRDfOOCHTe1JE526uQVfiRTcuW/iS9QBdt2A9OqvoGtJwHCn+BGobRW9xg
5zXu+QTf/x4xYWJxGwh5S3SKZ4kQexPm2FXKHIr8Xzio0sTI1L7/Cat7/vKj2Hbk
Hj0/KgsHTFaMu+FML0yhdEbWtrW5njTZ4NzEFOTR7TOBx9w0enwHG9xrTO53gBbe
vHXYHblzU4a1d4IiYfpK3vgXVwIJ1xNFL10F+U84ezuywYXiM3wKtv3kg+eu26zF
rmfw3rlA2T203xQsF6gppBVI9ZRmChaSF+ddhgc+ysx57c15Nz8pdmCDtB+ebQJR
pyM1ySbGbhZyKPHD3KkZyko/qwDZmzs4qlyBllbnD4sKCbIBPDtp9DKMRSkNCz74
lUvpmirQH4Q2QsdM28OvYQf2RkaBbsDfRhKecrlwTZoEI8bni+Bjo+3olBz/afJF
Hy/sPZcfIqPMbL8ATASqJs1DvKxxtrK4pO1UQi7+4W9cPcP0Fht4ejyylx1JeeOz
upE4vygwIKsYFMsiy9kgaJTRjoheaDb7wn8XTkwh7Gfo14Osjdbjo9Qpj+dgJ12n
+mu7TjKO3/dbXu7Xot3mVHP+zyBwfdne+0E7XwskCZswunXKjEx8SuDRMQIa+BFA
ZGwD6YXB3kMwzY8IsKDlrr+iFNRJMdC1+ZmTj4eUo2FvRXSLEho/orOuXl7ZH7kb
hpt30o0/6ylRDxmIR8mBk9RGb4u/xafa40wW53f0NvukrTljzMTrF4CWUzBmC4Eq
jQ+6SssW1nZtnZHZLPy2W9Te+Gs/4bNyCZwRzpstDUN+We2fM8lECQDwqsLjx5+Q
Z8x4jmwSpXC1he//RsnBcFFC2wFpmECofZ+pbK2vt02Sv0XU1SoR9X01jFmNdwET
f8Bk8+IIrodAOq5H0DBXh8wcSvlKI9Damp3f6xhOIcyrUn3Uesn0cDPlC/nCVqf1
S92l3pD2hi8vzinTBwN+UrSxFwtRiFdEyAxrbq+b0EmmyzZODZcPSaFyJhk5OWRq
llCtipzz/ZfzufywTcrVJA1cRGWDhk/1TKTbhkBaAidOsaAgve0N19CrkaKIGZx2
66nNHfRw8SYE35Yl+iFC4YhKmnekZchBLF91Mxs2OQtp1urtr2xVmPT7ITMXNDAZ
xkrSwOyMnyx3nUKV2nyiYtReeGys/2cdPGOT7/+QbedfUXo4BmgLjkZ287hYhKIf
+Gl9CZFh9wKnvCbFqE+im7dYK+ZgrU5ziCsf89uwLF8PyoePQ8kzKbbfu2U7uzZX
6dJMmwJpi+hiEhJOHBvgnl/1Jwvk90JGYVmxUSips5yKMplsxj0bTQktePeiJy33
NarxTqm+3CinSceL9bDVNKE5KJUoPMH44HBjKUNqKSNrL+Stu0p/E1o3KFR8P/lE
1JMGDT95Cqd4sOLGk4XNiaIFe9fZ2XbaAb/HT1MET0mFuS5oIA1tN2LINfuQq96W
onp3ripxnVDxNYYZm6z7L4LiLtTZbOSnbz1Mmsj5TYsT0N4HZsHBWzUL/J2Gc4b+
ZDIMKHlw/9tigM1qLcV9MZJa7vO5V9+jBlmme9DYBdfhJ0jHjvSvyKWOK1GTEeHg
BXk/mfP6YSas+UttJ1m1QuWZpZ4+yKVS2WG4gPS5LbSIpNLY7jiF+4MY2eJPOT1K
i2Culc0R9p1iktIkdQ0x6cgc9foR/eKILgQYN+sbEn63gisdN5qksUFASl85JnU3
Y8dHRu83+3aShHlYdrEHDit8lqvJCEhJVGnu1IK13pUtbGRyPGqRGokl1yarRPtU
dupo7wyAPkjQhToa82ZDj8WrsXMD/T0+3u8a+FaNVU+pVJh/Vlj8BPKl+T59oBqQ
LhYQ01dC684InloOWN0gA3WiysTEmPcuDdbZZRajwQyXoi0Wwc2oqqdrwLSwxpUN
suIm9xi6F1BvADI82ngj4JZugO48SFtwnnHU4htbxlkm+/WkY7ulHI1B7+4xyF90
hTs2OsAffOHHqt1VfYtEIeJjjddB71sGEbkYAtYfeu5g9sJqIVBZiIOaXN61OBYv
+Q4yih8i+TR2yD7DOJCi0xL0IK2SDBfb6VzAO6S/0GvMbKysbaRQHi8s0tksBEQL
9zZPahg4x+VxYsL9esbx/wcMWFTlWwWVBvGOMwMbsmALwwWj4xQzAA5v5S0/8aXX
aZg/JD3/H94YFkbakXy7dPYiPpgwa9o6u2P4ohs0Uu4OhobzCdPlHbS26NCpq8ic
EKt8j94lSNRhuq+/c7ey9LDr3iVl66oUnfYZIciuaoLRnGO8IPLHFHuX5jo7b4YR
RAJhWELGYIkmJaQZpuREfjw9JBtgYmbWsoTZVG0WVrgvZbDoRG/TbEXPi3eOgcS3
eWmQ29lzzoUgAqiGJ6AnswQYXB4vOOAb+aNrgwB1xhljRCLS9LRTUbBZJ71gBcOq
dTnK5JbDoO1n06oD66Feq2p2gWUBBAuD0YRwlguXRCa91/3m4oqraiLQvYjXxJd2
UopPZhRhhE/kjkYrWCBH0COyC4UANJGVj0aE9FLeaWw0g+X+GnGKaUx6ao2eo/5y
zW4a5pf6H8GUT+v1aG3RRow5S/oL1MprvNya33TjpiqU7P1TyJIzQBYZWItSP+E8
I/s6DVDk4e6fpXu6NitEXIF3YdAYrfPRs4f2tkNjLkSAJ4uhUYsJqN8LOUbaBR1A
hFX4rjH7Q8cmO+iZU4Eua2poJEQwhqWZYebUeGvhalyiHJgM3HZkTqwzwge4jiSj
ooysN0MFs/+a3VQdybqqFWPJVo3icYaG960GW8fMo9bj7g38IfjaLal7B5FNxWci
6v6XEMYycWGOekwbyuVZ/cVRw+piohOqpAXNHFWXYhIwW+4HNbfEOYPXQdRK+WnG
AEQh0ms+adT/VL4XRSOI6wZ/N54j8k3tp9cXArbhAuRYduJLtHUqi7GuV4/XgL1t
R7NojuA0g43GN5StB2NIW0G/dEaCnmGe5v75A1glJGWgiPEpQ7JXKrZRHKddANFi
dp3NOOO8d9r5Err6I+2XHovpzLev2X7MsFnCTL3AumUuOBva+KF4UgBc4CxyrlKW
HuDRVmlnA8nAcn3ZlbHaZaMx/L87BLyWzAfg+3pUEqeA5YzfEYQZmOhq1OlZogf+
DpZWvzXZ19xWJmcOCF3O/eabUULnc0jq1Ng75e30tH1CmpiSZfpS3Xh5lBIBLwNT
rnDqR4RDR8SC9Cn3Iy/EcZHDYFxcJQ3Kem46g/2sokuDcmP4skuYpioUjqh0Ie/V
V/trkkr2uNdbRsCjmuPpp6BfD4/wu7jqbB5qjRO8hR7ud93X5XlB3rqUqq8sCKxl
3qd0farQYl2yX2v0eQEdM+NyXYApB5leXQBM+XfFTgCrdmdZiQfLiV7lPEeUh4Wy
X6RUmxXH8IrYbVZRETayP5GElL5wugdF34KF86VY3sFitkZl9UbxpduR9wBjjDl3
C9YWi1WOiRGgrRRIlu+OLIJhTGdxqX6WmuLNCu0ZdCAsjxsVE9J5BV5uZknCAcHB
wHAYf5CaE23+kUToSDoJk199wTl8w4rv8wa+SDz+YXgRDPvYdLooi6We/9UlcdCV
m8d7j4pD3D1UkFZKX47Ci09MJBP03Gx3i/oDO5vYEr3rPc+lyXcKEITslz7hnrbW
Ed1fodNEb8DAh4Pqs/mSrNqo693V8Jddad4nzhlAHA/7Y4eq4bcPPYFVQWO66vCS
lTRTbUBW3irLMQP6xkex8be2c46oGoD1TQXv9noXiZsyddINdqfMsBlvjfZIAgFA
7NYneFVLkTjT1lSKjh2O4MnxFpmLZQdSu2NlHDZL8q0CBoo09Zot9aW2YS2mCNNJ
3KuU+HxbktTuVsHYjD8epbDDok23XBw3pgnpUE97XKFPyhJckrOCv5UPwAkARTIF
I1YbQahygetdH0a+wQf/rz1BdCP6H0yi5s5FyMah1kyfXL6FvbB0XaDMone91ofz
/YXrGbTKLa3ohXxi+B+08ilUWuWU+zgXxqP+5WrktanywSK9+q/7vXZvGxyD1+Xd
5AwBXJnDhYnLHIq/6aQMgbxGBpad7w5/inV9raWvnSqaY1TJdWCe+RbfrvIVsudK
5pu4xPNxdw7oEu4jU68YZeLC7TO2JTlGfkcFpUODnhYD29aT4vJ5q2rYwbOwZu9P
mh4RA1YvXapFr7G9/zICeKzNO6PiW4r8PTIKWsn8pt4EYVuARPyQKhA6YAMMhtHd
q2vSKC2NHA9qnqhxnnYtmzbmFId4IZzbAnc0IcESHXd/mXQ8TTkBnlbKaazOHYUc
BbSqtWb+e7Jqdj3R8VbB+xSCzkwJds5MOE5eZxUcFIgnXRinOnYGGIZchZaRhFyY
VkaNijfratlu/w/W3rg2yebyl5hrHcwY7WZY6cETOzj6Uqnc8v6YrrEPmWogMBqP
UeMDAU6ukiTYvc7j1dXbKZj4kSMmaI+RInhXEc6MgDSHZdIWcKG6ALqbBGkY6Fw2
R9uOHNkVfr3bpjA4DW/jFUYJaTabvDr++b8zPw8lXUWrqmekpZ8Qiugfao6INhdm
XO8A9jzi5HeKXdi43tKkfL/6jeqd2ixwPfzDyI1oervIliialhCSPL9F4MC0mzeF
q4eLP+vc5n40U9J6A+gPsXBts4wAcWHGaudgiJ4xp0+hW0zKc5GLbEcwpsH68YUV
mMD/lYB1VN8rqqcFs9yMt3D2GKjVTdd6jmQV4ba0C/vFwsJM5+COdhf1rq/rgKG1
Wm2t5XsBQ/CfA5foCNAA1fBumHM5ircWkr8X8OdPRhKzd6SDni4fKPHKAOc1o93a
bI0v71J3DSvHaOgFlbDqadGuEd6pfyrLFa1Hdxvs4Mmp8Jh19xKYL0mxHyzE8YP/
p2BTl5W4In5RVQ6+tqTHW14+1gpJC1yXggydx6H4r68U8RhGFNDEa3wkjQWbVROH
i33yMdhnVuTdhTWsCe8IFMs/wsjc4ahGOq+c5LnuaQkfD8y1r3fi5dw+tMZbfYbR
dSHtyGkfGLkYUKZ7GiMfBYaYPCe9BpXsr0BWi4OorV4xzJMANEbinsxtX2UGXeq4
2lp0KuV+vF1xl5p7d/PPl1kfwrfrrXbG1NB/u8YByqpE32Be7sUHjvizQq5Uc+gB
K2r/Y0+c2jtqATvpf0k8r6r6IXtG/rZPAFtqvPU89H1xTNEXjdbzNH8UCDH5zJig
ZhDG4f1zz97HGr0ztiwOo9VPaOhz/5q4Z0BvdU83HALPXSpV8s/BXJhB3DfJzJsx
6SLENDd5BbojuKNqqGJWDzHae5YWXR5WFdklw1R93DvPx3IIAAV9RkTrb8dxkahn
9aebfIFznYdlruRePM7wqV0ACapGczE3jhpK/LxbIrsd7rSeSjzfA9pyo2ZzUNdF
89brGIjO1317FkS5TkXniM5uEgcy1pXPUa720HK35lei13QEB7ckV8bgFOf26iNz
pUcuY5LAbBU/leSwvm7qLnfj0aH3+mNshEqMFVTdRFysLQoaazzgbTyvxHgxVZAN
2JpYpl6JjzR3CL4TuabNZgJ8CRAt2Q6BN82cCzO39lOIK/TnXyihNeG8vFhC7Xym
5HY1X8zPcZpGwwvPEOWJcLDCFrg3fbnyJ8GbvrYdXihYfjsyUetUag3Uljza92mH
7H7io/ikjY4kwrPSNUKwetWfCbaLocDo7rRH1YOy5kDPuh7Xpw125uogPjf5CRqa
GShgHeZd0/2+JpQhiOCMIogX1QXSnzTRHX0XTsInSSwUXnpENPBr9Hbv34edD1sO
wgxnTnGN0NZb4fNrl3lzIAB1t8N3Q3Dw8r4RYjZi6RnPV1Mo8f3NXtkismT1n9aK
BoGdaoxTjsWOBwKTB58u6DdAnA9pXnys9uJCHMTEK8xGF49G4qvwWaqZR8IGEbxI
9OEi2B1onqd5lk+cZUGxAcmIX/KSd/Q762QQKGIGoG2uV9E7Wy89wJdsusgXVImo
b0NM+4QrF2nDjVyZGbuQJdovkVnOr4h3HTQ6ny/YdcJlHTuPfWzCYfKM7HFsSNfp
KvnobUfq1Vk0crkIWW1tFJI08hta7s0fklxWE5bBWSxXMLzLl9EHSE7qUI7iEVh4
x1Ev+kC+x+uqgDhklQ5sgdjlTunt3aLX7k4Y9OyxkKY889nVK3BTvnxqZoqwP7Sp
+QsozMu6VY1h98ZD/L1lMPS2sz/zp4xotfNKKneIC7lmVzlYFhHSxEeTPliCxJlz
CvFa59RUR60N2D7epC338TnWtTdDjGYnAUx+Y2i9sjtcZkLwMdIu149OocrB74yS
P6XKuAQXanNf4r2hUr5L79m1fh2U6N5A0L+zHgAmyUHRvwRfUaFA3BQbYuSIcvRC
GZg01eu3HoTz69e/JlE1NHqk3ga/8yqrOA56A+oo59ViIfQaEjjzwiByLRVfdwR5
F8sBrintkMbfNlH/Zp5v2+5+IxAOOApxY1eonjNQmKTvkn2pLbytIgjLyQw6d5NB
5l6QnV9l4Cypy0F46KBrFqT2/Jk7IdJiXkx+CQ99tyQmIpSTj9MmDA+u6e2HepVY
joAALEBEUGspAF/6HZllUm22mb9RE9Hk/PiLWZMEeAlU1/TUmb2HHgWhwWNTdCNy
3wHaHhZmkCtmss8bQAzKNhqgd0AW7U6iOL+cLQ5LHSFLY5CLjITGswrrRS0TFkqM
+S5TzMn60pug8GhQlegK2256YriTWHXtIpqaLw3ayzv+XXh8Rqq3dOa9Zfyab4V9
Hp9e9kiakOkkLV0MGSF/cdXyALeXT6xtj3Xu/SI6+CqZSX3c/ah1k/Ldv8Ka8TEI
0SxpDnq10NkDN2Y8EpyGVbBmovMadh9yRAyFaNtNDnm2+zkhZM/JR7efBK+9lQ+6
q+SNmK7Wec6aAPCxf6ACFyMIvP/vMSmJ2Jmdv4VffxWwmh9DExynr+zPX24gwhNT
ajqssXhoEwW1cOWUU/Ly/B7yR4ipQB+O7g+4U7m8VtlPKlZWUxZ9Sx7M/B3PtDBb
89O1FBxciyZF5ita0RqbMII+TrgSMYC/mUjYl8RiivjfJROE/RnXzmzQkboU6OI7
8z6T4RShoq/5VpY23eCNNAWFPzFVfuL+aY5yi+tquy4ykhih0Uxw8DnIQnUB/g9O
F5MFIXF0z1KdBwo0D4fW+I49xRxwcV+0mFo8yvwqJB9sqCP9/EFDwlvdc9ynr4XP
GtGtJL8bl96Bif+ua4pOXSZFzVw+PWUkwV691C/4a8dO4kj138d/YT9YdvxG09ZO
/2WFbEqvVathIbnyrDDvAoFO/DB91W5qXt9SRjL3R/VtIgDF5KAeoOIIT0QAWs/U
eKtxtT0cPLd+6lysYZEXIxcU1NGNuLocWJdI5oXT6iepfQefq+yDVadTgpf+Hbu/
PE5sMiRnj0JVeJY4trppxHrWtJj8F2OcuXx7IDMBoug58rqHi2h6eR9GOTIM/G2t
4hmwsWek+hun540ZoTXGeoGam2Xg2Ouw1gvrcOoiuhN9D75bEQh4ZNjKIiJp/4DL
l0wZYbfjw4KX5MKafInI11K9zvo9pW94LSJWD+PXJiXVWz9yVRwBGKPCcy8gmeVM
ZXLayMXOO0VaUNGkxy6s5XbiyEV07AUwqs4xwXf513utyeVrLL3hH37V+Ii2jyji
olMfwcw9tBejC3MH5gVrVBlp4deU4L+iN5HNuZclf6+nqC+GV0GXt9sMXRiESTcJ
eCTcB0deMfAdWLh94EDLVwCbluxA9pFXzJF1YS0NO+SQra5EfR9k/m8Z0obPJcW0
tcJc8WwhpevoOJO1+wbJcM7l/ns+r2vAM5sw/oZic4B7h1SPecDyxzIhABWkPIja
v4eEn2DNfq2F4ugt7j4Eina/TSBDYbu+xFva5MdU1dcwFiA1gdTIs6LcSLZYPLsR
rFImva1VP7ZNAU0vbih+nFdrJHLh7gaT1G5KoI6qeG8yHiRJ5c4fNoLq7pkeK2Ba
l5WfzLaKdOVmZxmH4zGUCgvFJvfh4owMV9CN5aiPEw56gXM2hP4mTBujp4Hf7RXC
8D5xXnDs+6trHlJt7f8R2LE7ML77RrKeEMw78EHIQXWrpq/IfObiva/MZgjh/v1n
KZwuvl+QKMnj9NZuAiyzlAtps9+JvtTf7jVZdERBIsL9JbM+xWvtht0l5S03iSnB
9T/jGC6m2uOQYfiA75G5PKylUOfLYaDKazuqKxmvRyXfBXK9ApbFB+VhdUgQEje0
yx/CoEGPKTfrS2jUtdrSUJvi6E4275oOYA6rxp1budLSusx70h3rtorcd2XN2Fhw
W6UM+gzHUzGk4hbW5IY2G7tv/3nzoZkEgtH4vb6nochB41v6+UeCrF3ybwyzBvaM
TUmkJKyc3XBt5LIVB/Wa75mPcQeqK//9/tBEeezXZSrkgem6lpePI48DOXuxZY/l
T0iVY3q0WHLRDu/VBGp8Yhps0311cEQszd+FEP5DvAGrwmPRG0yfWJtZrneagXmX
ikHN3vwYlLOJ0w7GPQU8dzKx86YMpMrwkQCSwox0uKvK0r/ra/+V2Ty0iHP1Q4RG
I5Q07AAR1isMajVft7mXk6j5BxGyXnIujclbhLezdkEDDp/g/TisKDupoE+mXIjm
iffXpicLiW+C/uV+wxacV4kIoITi24bRGpx881EIxrRV8pwT7QnfrQtAMUOAg0S3
4YhfZC4zxB74gGWxTWHeDCb3a+ZoDuo0/43C7HkYfhB2+ti3ak6HiD+RxPjm9e36
xS1gukHfZ+gecPOFbS/YocvkpYydcBvSAlajPrFq5Vcp9XarfOQeyHWlWCe2pb4f
n7eoidiwURGIoQ8OCGqSM9HsoxcsBRjerqC8GSnzKixFlhA9fb8gjKxHZrXi1uch
zy6FN0ffphkmx0mwwGAVz2cPpVZ/yhhiTeMTLs3qgm9+RTLsvw4Dfflj5iNNjecl
fwiZ4gNnqf9YKW4NFq6vB1ocPIqUxJQtlrTmlLPeCNAeKWmND9EaAC2A7/etzNY1
twgkYgThRsACi5b7EDnIkOPr7aG9yI1aMTn9I/JrOxSBtMab/aVOax9rxb1gkqnw
LUI6LGgJ49Me5UD/HaKA3dO200AgVqLvkK/3PR+WTr4LXgJTHoDRaJkAi9AzcrQI
1IUlaLEb07+joNfE3eXbSAvIVzbFcKZCVCUViwjPm7DBC4tcNWm6HycI7kVmcjQL
dvn+lAxHYNpi5Sw/2htnmrqFNQG2W0I7o403BNkSNxjQTBCMDW5CFqjSNcHmcUd1
cXHKppgQREDquNxd9cbJjC3MEWgNcEweeYPO9ls5xFe44qkmNXRHsZ3HSGiDF/Om
teQnTrDmvGxWmfZ27ABhCTtONgEhtRBVtoTPGo8wAJyFzpWNnZjkhXJwvwK6h7bf
xmE853Ou671n+JGbFYirOBDHjjlpUnLhbT7frOOBPYw9JXFR/CYd2jZ2meth3+8C
tjqSRUJPD8bIqRUGIpgVGxiUmEG9Ff8FTOZWVuV4eYtZFXeoO/R+tEfQYXKy+ul2
qrzH6RPh2VTJIK6VTGsSoUDMB4hbVsXgVDYNYM7G9z9cgjvqtnhU9X2OWb1Ilndd
3kqN42tIzpW7ji55qYknYCwZVHN25wJwYomSfwTe5ibZMoQHT8lZ2Zd+mpbRJ5Xp
pJwpH60rSohandmXLJAYTbxzS2bNxN5T0uNwMQwWiYQxL5u3FYdgjDU0RzKv1nUp
u5Fr+y++dcCC+8paSx5o8d+gPSCM1+Mqvu9o51yPvPuf7t1Hgaqv0nvYj+mqIBEO
ORWdL9kGO3K85BfBIyLF62GCKoP8WY3VmZjAb5F8n/pPH7vYzGGr7cV+IG9Ucfth
5tVukcxpGyl3Fg0JIo+oK3MuIko1if5H1zSuOtrHvahYV3gyThN9m53TLt/F9jXo
d/H6rR9x0TpqYiyB3qQPSakm4wyC8PBNxh3AuBmXYvJnM2tlobG4LE/0c5TOLc83
1Jy6sbww3LzCBRHhnGz71Iwwv84Q2UugaKHDqNuVtZb7JuSxm6aZFkMcM7OzX9LV
l9lSVxuuWiwX4IdCYdtirTf4Aga7brU0NbnnyDLddr00ybmgOIz8DlP3Q2peqpK4
51G2Auvde1+WOzNfrCacG1Hyhxgp/lQX34xVvCJAawU+ujfXB57vraZOfPbqmswB
7lzbA3yM/YlhgGRLFmKhjLFm1yqseh5OWubqr1laS6hQFAx5Ah07TEHd8PWKgmzx
69kjRQtdR8ptU28HKulow8t9tTSSqKDRLuksQZ1wW+EcI8bLXL9rgUHnYC0czpY8
oSCnLDs6DVXEMtPw31cZivWP7nsH2cgJiAIsnPZpwSCAbSdfEa6J5Vk6FVUNTGTc
wtDMXNPNU7ORvfZ7k2lJk1SH/xKGPXmU6S7GOdlwztZ+mtneg3fW28w9o59gXgr0
eRMKhwZ+Q0W6zBwgSPsNg0ykfkoEH1M5JM+L0bqBqCd7VrMlAp2iyvR2Qhq1/7G9
iGdDJm1+8zy2bDNhaXVzXJ7teEju8jaE3ozT3QQ9lc54/Y9fiFHg2HhLFmNUVSwi
vrx+iXYQmMBot3b3Mo7zXopJsoU7f4Tcjt+OTLY0oKnLTVplS1z965HiruJJTMc8
Lg7cwsloN4OV7n7ZbA0z/fVQBGmb18fI2IAk6ZlbffLX29rNvsxNPuwXmG6MmIKt
buRFmb8a1k3+ZwKRp7nIqp5bj9dbFpr9sPB3z6lfod2IfBqNacBVcdhaY1e7fW9Z
Xshy1tvqjcXnLqDrUgIV4PynwZ5W3XpPyhPAgBiEZkwoY0XmI2PsCEsMlD/xYuTS
nzB6hcs+Rot4RepgXRgBeZVY/kL0nOraIFNtsN+9D3AMVy81bBygRsHF9qnxD3pU
2rWaTHyCE0G+tYukk6Ec0HJ9tlo0SyjHLPNFQJsrpbX50o2nNJSqKAHFxmkncBV9
oUW8CRMmCQWHKM5KLE4fcO+2hQQJmWyuuPBr+7eSk/0qwkJqIwucWIeJnp2+eC81
mhiVm601qJ4Y0a8e3nD3ds5J3nMbClwNw/OWnUBfch13vfmFcJhkSoorpVk80U92
ySiuHlUnr+HT5s/yvdhu7sOcZuxfMQmXg66NUktZwjd1zGhd8zt4iXlI3Ca+ewJe
2kKUS+1zEGiATuLhhJd9LhQDECXvssWtv1q0VBoaNdTGo+7otOqpuq/nzY1dvfoz
1pRI0I8cNEcmh6uRDjUtRbE1AQIQqDCzKZLbMkuvfgju7EFS5fKztmWf4JwFCVOS
DRQ7G409wm6ZKH3ufFThYTE9bGNOLhDW0OkEIAwlNMseHt6gAhgTlmvDCDTTc6VQ
S5cBuDg/J7lHceYUflYPK8mOFXb+IoOrnximNFKftv24Ks0li7rzaOmwODRVJg1D
LVO0vMR3Glxa8IsllY5LZ/6xiV0A2bJw9Nkp9jm82xIlcuwv4p4sxikL59PwPItF
WJ6dEKeyyz9/Gn0WZCAchER7HzbrMiqFnfjnDtK+PBlZx8tlensYNh1A8Dq09TyW
4mO8JYULBp2ERoOsADVJGGDQNWN0ezAx3Uy8EkUMFBcdS8scckvsGYa9rjqHFSfP
8vX8BikbLSYBQo9+Dir3EoJV9xNM9YJAMipV+Ni+Hy7Ul0CjeYwRMEyIoi82k4EP
GD/mHMD2bWphVg8D41iuTZ7LSQvnF0n2cCD8Vll+g7ylZbbKx57SoUFod84Gu0S9
fM10KlyywbUZD+RMa6FQ8yCuUxorZHJT4sUx4dnQvLCTyG33hmVhxbfa8iKxZeFC
WB6I3g2QUrR5/WlCtZcXPjznLNsmQNMSe9pEjUZF4DVHBuPimdpM27bLIna0IIhp
lEfkVphFmUzkWinPKEjQs4VDJDFhAEZ7l0nBYv0TNxpqAVFUF0oAttag7oPskZi5
KHQgJo4wVHmxyPA3upNb+qI8RiiM6s86wOpzcIagDabbvUBntycbm9bHPSEJ6GHa
Fv3N0AWzWFyAW1C+yBL961C7MHoEh7xsPSWq59vf9dA5Wy8yrnx4++HxTyFtXXq/
Vv8ClEOmi0/o+jU8ZyVjnLx1yFc2WYBAndCqp0FoK0oBRS6IDhf6X3FaBCJG5cj8
Nyy1ENyzuSo5vLoV15INZqeJuO6iu1cTJ7qPVxIuhT3H0hihEzjYOwITVha2yNav
nlZETA/rDdfR1Q/U3QhE/OSgLt/uMMsmJR2m7+jURIDshUMs6OS/HYEDDmpbl7hQ
M1NqEZZEFyGOZxHh6MeUMVdPN06MrZHtNR2Ds2NlfO3y2tzcn3vKImBBxSikgee4
VOrHYDDgSrobEAohTOVNGrqj1iUrZwyGC+cAkA+bdchmKh4ACC3GnNEfvFsJ3E87
QBya4dCMdANxltv98fjx5FoVblEIM2mO7rg4ataUjcuPLJE7zMsNKdYu8ZJoQzaS
GmF0wiStP10X5ee8JHGYXpcHMtNJVXBQNfATJg9FWIxpBdpLIqvBIMef36zmWe67
ZyEksSR23X0SlbFe7WOBPnDOdQxZ9/EPmHipgUCr/NMcAF7rj9pWc8vkZJGZhg9V
SgfuWKAu7qgRVac5yfXVEIpgsze8+fux51+FQmdPWB/yW0c+/yHGg7kiZnRxcQgd
pJY3+lwvjHqEFsL8P4JEoFPaCsChvmqLBG2kQeaqGWpDpLyUR10hO9U3qGpV45Ql
A9dNYzQEys/FvSQo3QVh63hlTY8TlzvWVyDmSGl3NfrLQhi3WaAmaQwpJoZ2cgnB
UtYJh/Vz1o7fhLcc98dROd2DhT2ejd2+04xM08+V2cf8QQDOokKWJGBP3Xh+q9B+
xIhw12rpFgs5QkFcLk1iZoWrpgn35njkEDfWAimrFwERDrcowe53kTqjTTe0tBTr
4Oo0KZLSwZXI7aSqHCB5mJdZz4hbM0Fj27RTviTCJzOhR9wEv8NH98vYCjRvo1Ds
+FePhyR6ICk+gwSqXsbr4sQMmS/ymZ4gIy2fWXpg1VEFJ4+7Tb8fLUldFUAXrU7+
yE/eVfX1A0sLzoNsWMJtPWH3MQKE2dQZaTQn6LoovpyFaeqmABAGAq9NFnF7qwzC
wTFfCRVOEzZRw0vHNX2IrWe5nkbIeJLTWSfAeGouY0wPTmvf8flFVWe4jVJBExcq
yXXlsEBslSjINMKfUSvGFJj44GKzaLKqN3xrAtzZsTI9fH2CIFAusAZ9mHSGxQlz
sF4ok9kGD9R9QnXGjJwRueJh9no6JC1i2CVrsOyt1FuJcVKQSvDJzuCdROOTQCVh
clX7/D4anzQmpgo5ed/FyMa6Qc5OL2oOmpVi1zTUT40qMC29BkdM7H/u5k3dmjpF
fQDDPwi6sw3X/bxzTFSOWEgMM5Rt3k0ZrOorfGgG5svXxQWSCy8NnBgVNCIrGNXa
/6tnJmhsobbPJGHBMPpyPS889cNU8ZYlqK/YGWtAE4L8Eep+3xVhqabfzbmWJV5N
Rd4kElmnWeDvoXXbnqMAWaYMm6bxsjjjyj8DIwo9fnZjYrthAZAbI9Eb40GhkXwW
r0EwSeeNQoa+8HFcCbK+6T9kCzWNu2HCIn4ioCoavra7ouVwXvAsPNDBfq+nE+R/
+ajm4VsO3YxS0+sHH/Se7Yre+rYEA0axRGExDIykAW12KuMDMsZSRUeMbwqeO0d1
Lnu4ITwPuKPy07WuAgv2JT6s5ge7LnsBhgh0pvRZVPunv3MsxsYhQTT0qK6tnjRe
4+cFwiPSMeJjNKBtkofynmNQS1xWzQUeROilxLUGQetV0/w3CfWbj3UEaxQBmoyH
39y+OezGmXzAzOHSetysb3MxDpJknZENMFHf2gHyilc43i4K514OKOlEIlIlffKo
U8ikbuDTEyBogwmTIcmfanF5G0b66QluiuYEOUWDVbbc2VlgdvHe9t1ir86BnrjP
cmUeY/tvH1cJb7auWxjg38GRpGwh+invkbgB1H+n3C9BNT9jMuSWzmUMczOL6Het
5l6C/HHuoOR7LXfy8j/PxLUCutEINL17huABUC+EiPrXtwJIrPX9SrYRJsc+OuyK
p6Je3M0MyDEp+hpZ/HvYpk6oku/s3cz9Zrgh0FQK3sy2eOn0YwMBIRH1pK7dHa60
IHTDLYTAc692EZ5jklFbHyMrawfDL8zxwy73OkuyXc1KExL7uxyZsL8Y1g02mJtQ
Og6mT7I8r+/TtsyLaWPyCU+lywDBTsEu3OCbmq0f7CUQznEAA/9HiWR/DmMn2usU
56IKOZ+ICmjR0S5rlDIn5hesBPncwagyU4kplizeSC1+u8hdV3br++fr/3Z+45Jm
v0/vTSdh6BVTMHEG20H2PUS6vI0kcsl41LRfZ5Hth0RhqLHXWO1xCt8i83TY0ytM
WZrRofcy8upV7apqXHrRg/0BRXnIYFzf12a1lfzdwnvTjPdGVL7uphr3a1VCslYz
rKRc1IGz5ACLs6OkyTxegtMOjN7VM3pH07+OheB9SpllSR+USJ8Xh4BSCZuOp6EW
E2A5kzOl7IJS4w3ZWX8hP+nxAGP3FVrtK3kYZFWQx9YOyY1vcduaujo1+WyEF0W+
JRkAPJO9e82y21KFRv4dNFQhPmBzEO5vu4ItGjSY6mR3itD7Lk+D13AalhD6tmGI
IvPRDcmYe8hMN9VKVld4/8EVf5fZTu04yishB3trQ6gm+WKkYRZGimLhU81OuFQH
AIRN8HLjHUCTqse4mG+XfDaOnwFANQ0So2E+C/00FkiUeaaVtjYVvZmDTObHBAgB
TxNq3zAWbobzQmSLld4hy0S3XDgzohEeFf/FdyxlA9ZjoIiDpHxx04vmV5nWS+iG
4kaPGZsQmWBRX0WbUSwrOIc2uQ+BY1JNbKj1rV4MApi9+X5+Bob9hc7erfXzW+VX
rJFN/GTHgO4NJpzL9zh0A1mJga7SRBosWjT2N5b2Bq+6iiCr8nfQqDL0cIO/9hA8
yHLHZJAaZ+VFlO+gyirBivZ9KDNs5hj9tf4Kfd/RitTsVEqX5XCKVL4YcbiPxiv9
X92yNDj4djVkpyEJsTas0sjSe9eYLGz1aaJU3lIJXMq1nXKC5/4ota5xUP6qbRPH
/kDQujOP5x05gnfs4dFrOqqMF4xpJW696QtZcm+8EY3YI4hTRDkgo0q7W7koCf7p
km0Crgz8wpk3ExNy+120+HSzH0499Ra1Ww9zX6Psd2W6aThqSnTmKCWo48kk5CWv
mLS0jogiyzQS3iBIRArsO1yKsIVnYyGmmW/DNhsYL2WXIen9w5NPP6v6Lfmf+8SR
vSkOSZCc7eyfdRXjpCrFVcLhlJKrDM/h9qtwBVe6SSJDTeO1q/tCfyRI/KaPPAFv
kDJ+yyHs+IdDvJiE1A8yRlfcdW18AvkUMu5ehfMDnMV3WmUdk9Ubzqtql6j0FIFa
sa3UvGHur0T3JairGu+jD79JhIyS3UfsEmnNGfGgLen1bykTds9Ia4/gePwY5dcH
DZrilZ6ORjrEn7EM+6hoF04Md1ZTNAg301qBLwfW9gjWLQ3KwdpSq9kZoKd+26md
wWB3XL0mT2gopi+zaWnuSXCFcs4cX2VIuTgFOVoUptr3t3UKHkONhqG/6VYC2f2r
//IWGhU2iuiDpGERAPNYWfj5/kBOvK8PIxqI1a1KwggBjEKXK1tZitDObpa8ALYa
0+UFLDl4B/4vEi3rN8MfwIqBvya3ZOFkNlJUejYUJUg4kkSoua4yLEnzN0uzPXSi
W/ws6cq3EVqvMovpsjmfZKtRR3fmu5EWso6KyIUNLojcrYGA5R1V1ptJB4Yp/lJW
R5kOHp6DhEoJDtlMpxUP70/7W2Z/LhGwse7wpLRR0fBMGw/tbOp0FeZZjfIx9rho
bIbyJbnBdlm92jjk2U0/4VWT5dsRyUjJR+kTDMbQTZn4JUD4zR/pCclmcjnh8Pvs
Qm+d2B/VA7xHuvcCT3c409qIvopVLvNGTdfliJN/iQuROcjDQUqI8kXqY4nXhxCL
hFKHDaAjD3wvifO37k66EodeMNqsD6zeMv1UBTDocmG76D8yh0FMxkBNtzrJGy4z
+/5jqLRVC2vELQ2sN4pnLbtFqPgudbWHpYHpGBULYWd85RKPl/WG/ypvWTXxtlY+
Z4jOMH7WlI00BpnyKwf2CWQNIOUXSQAq32D18YTd3QYoE97Yya8YQ3YlPm0U0AdW
PMQFLdIkHwE4GRZ/hRdwnnIoU3KaS91LuQeafoV77uU+q5FiSI9OGxwfQRii6N6s
BcUcnXCWrsjPOZx+52VSyspIsByVQ8Wp0MtRkpASTvYDYRl3IgJ0R9Rs/yLWVd8F
5cSM77pZi6AGRFjeJuI/K6ZM7e0i1VfBpeQ++UHxYuirDHGH/EcMOv1aKYpc8taX
4odZL8FzQYAsgjQf0XilPjYDGE/oRGciixj94zuzfqXaJfrS7I2Mtf+w5RunuLkk
qEr75B3D6plWyHs6Sz+Vrr7jRtQ3VoEeTjdDHQJ6xoLctUPg7TsdJduuLpKDv8X9
J89FrmDBt9qBSiD8Yigb3ES4id71hqz3HcccYSJOrL16asGupVXbhO85kziHQO/Y
Yx/WDeT/fQdYiQ5sc6NhnjFJDztyJdvqFM5ynzpdst1+2S7D4DFk8N87MlGIfcGm
iSqAAK8ceFlopt4TWF82SOZOCS41PzMSkArUtUDIY/gU+0eK4fR+Mx+h+HvS1WIz
knLYrT5cmzhwed7o9FUd64VuHrzpvENiwVbhpSA86lt5ZFlcPg8FbNPSU262Wa/Y
mILEXZUGQkrKJdtqlPbG0YnfaaZqZxTdnQD+TQxq49Jf4H8WENRWkcNMSikJWUmo
Mf/ov4d4e+ZdKKnz37c3qtrKF1jiIM7m5a0ywMA+TZJDNsPNYI69UZ1I3JPQhGkY
akjDnj9fOspLpTntamBbJdLYSiTAH8r/BNiYD8uxJJESUSTD8U3BIfgr5xl+Ipih
bDdWoVuhPbDO0/BusTz9bx9cCiiIBjIEAfNxVyTbpCw5zOE9IiKC1KqOJ2YstvYa
sZPisjHppLMUbXaUqQ49qGnXv7Zf1wsPiDjHQeDE0Rj1j2UFmTCBGLgxY2BukOZ+
Ge5jT0IRDQFLlJuGX4wOQeASPdUxjgsDBfxwwfm7XWkjntCw9s3dwdTs5+aZOxKg
09izP+S1wsb5cOCg47ocFIQA4CXH84sg638z+y35rnneLAqwXGYmu6e5mKVHTtdt
bbLzOMhl3II1CGj1j1NYm6qxbSCokyEa6SA08AuhiUkRYA2D/FJ9v2T+ltsfMQcE
NbtgDPKQPT7J1xeYMosEuLSxkngvUFY9yUWgJEsnPPPpsXhv5B0oSFhBJVNqGpkr
2ul6go86klvVedSyiQfCpPTpArx8wSq+1qF6L0yU63SzfQh4TmZ309uacVtT931q
MWfddKkaegspwfXWzerK+xm0CM13m8BkmrJXli/FEaof+PE826s7NosJPjr04nIH
pfSfIRvYPcNHOPFAtd2et208p6PuobjHelXtE24AZ2Fka9gZjhfxsoNKhaMvX041
mDPr2/BWGCfIauKUJFZtDureZslr94DqrfJZq9YaSDCju3UNwlVlk4t8NclKWnqo
cayAva2lef8XY+8tEo7Sv9CdJajbmDXf0JQght7Jqtqm3k+ZIkLuxY0LALDoyXNI
ThERE0XDV/spngkC+bEtRrqawxM9QTPD9eBJ2DueeuS3kRBTbKJVKVOtbMzkR68q
hymj2kO+ip/YSkZVR1JD/EHyrhQnyozsjp4kVQp0p8YHzIsDKnOlZRvrXh8wjXM9
blXd7Y54O429lpxbwAzs8BNIzqi9IcRr+oRedPdPfQT692l70/tlJYfzgED/c8H8
IJMSHtyugxkv7yPT5ezZSoStecGSBEum1h77bm9PdK05fQM84ml9c5W4rt6/gxgf
NUAWQuGzDIRi3ggkzULwVFvWkJ8BK9Y+noR+GMG8jqwswuQp0uLN0PYSSm9I+vWz
y8+7CsZqWoRTpZWMAKRGohYBIAJmsV4Ljjb3HqNGvUx8LDdTojjte8+lA+PC8jmx
NbTzwB3DMPe4ZESH55VfUUX7XqoKpUqTydbgKsU/l2Aan8ndp1rApC2kNv9FmdK2
PFUW+Jsy+J9RQoqXysLZSaSLKgBsTpzqnqdN5YM8hp4n0afqox46v0A225a92J0C
aL8nFoVOTRtek8xAfYAqWDQwWzTlf9rt4I5HhcesU6oyKqYo1ncjkv0LbAYEBGP3
08/lHO/tKPd7KVpiPdkXFvwcCavKX+EdRE6ym/VZgXSmBVLAGtnPUyxeISX1sIhA
pr5h1GpdQHe+q5jgUO5ONyaTJh61QgaCbHResMGCKGWy3GP9K4bXt6x4nF7WDs2e
IQhuSQR1tYFkuXsv2uEQWMHN7kZEiJ1znGldurJGZ5lvXOWtbijxK443ZkuETVGD
poVvKRYunxUtYBZKBhpNYh4Izhnu/7VcCuz4uTBxz0+1UPXO+lsf7TnXMG2ySewL
JVk21b8P/dvAhzOMPvOHIDZsbkmIKUyH7f6p4cozuSxFGHdULEehv+bhP58dzki9
hG3wias2sDFxs4mdkHIhUJfgWur6JbZQ2Go3WNbw1PcF0j98f8/YIj0W5Q7qgdSX
MdNQSGEgg4TokaEUfmMChfg6XtDJFnaZQW1ft5FngcYkPGgkXzvBjF3v8P+K5y9t
2wWb0uW64+77xcTXR4TGD9h4VmJ6W0b+gFUO0OqRTfHz0uCalrfSCes4zJt2yjNv
HtUo7hiDhsS1MsD1ADRySju+c93fZTIs2fQFFX+1hVkJ8V0uSfjW9wFurhvCsoCy
PY1c3pLaabWPLdulbtf4XrtUX7C3WbsV0gnwbNvAVx5KgNXm88O1f/5+dGsSHxCc
r8R+6wjakkbdhY/v0JlWw4KGurHAxCez1SbXdMAThEC9DXMqMhR49ke6FkKRjmWc
NHVAMdTb8GE++jN94Kk3ApTt+DfOThbCyXG2VtgVQXsNfZMxC9bvYFJVnFbXz8rB
kC380RZWQFxSNmvuVH7lIQkrVqvxctxdvBaGbUIzigY9QFcfSM12lq02hdSaPvd8
6sZkJfu0/xsOGuwBiekfDGV4S4ejEMIGFwjxFVRV5v1B5G2HR4Jt0+t3SPS1bJX7
dq/sh0GX4bnjDvYBJMduqbpLNlwMNqdfBsKHfT1jpeNCq+Ytgr3NpWBKDBnT7677
oTsjue6pgO1d2Uk76+sx79htHP8h+0MeQIv9ama3HdMkmVhOxBEkN5aVMZKaJm9y
IloeGY4VrAZ9hSbr2KUHBZ/++Bbal7d1Nsy7uyevKGazbykvaD7uzFRnU2JVFLLb
1A1i5RYrj22zR+k+7rEyz6oH3KBNdCrI5O1fBcug/qrOU9kK1/EcFjRGrP3rt5i7
1hvx2c4DjFf/Diu2PfqaEAti+sEH37SOdIzpkCUAths3UHm+8cTXFdo4z6MEsaJS
5cmpJl5rm7aDsFgTsq2C3tO4U9WSb0w+GeZYw/yGBONmN72Q7WUJSwvcKvKosQLc
yQwbcaO1YsYTN/chmOQCvRxsSC86ZbPhTdYfDbkyBMIU0JxmgAwTEviceKm/xkfs
8ra9UMv77hYMH9gNhrx7Vzcz9N9qG1f5niK4NdnjhMYty5TLcACAT91cFwYJDMrZ
4OzRNN91AbRQZwZWWLTA/ErUsFUdoZfKxmOA3/rVDteYo5D7KTKGODR59JgFyKBP
a3CPodU7/42qUV9PjQtdXs94YJCT06wPa+ar8FIJONapR3c9SYjCM2hwO8d9NHFl
qqTlPQwUtMX93STmBDs1vLNS2WkbrLP6oXxxzPuRmc9AoqB3kuHvPPWxuD+FsUps
67HUME0qVJPj+SNQ8gbUSX/E5zrjCGOQtiXR/4SrOXOPXbqx+XwWV/mbKmeX4yLe
cn1JKQ7ci6gdpaeWLYdrlevi8z1f3sC+Jj0o3aK3nhh2O/jk5X5W2Lbey9Tuq7Zj
onc7IoVa64eJ98F1QBmRB2umHeROpA0qS5/LZSvkiFZjme5ID/P8S69XiVifuNA1
4X8wW4AkyPkASXCQzASZajpBJGDoHaEXefMKbDXdL0EIGjU8JMEMbj4IGSIPS75l
WB6eHqioBUqyuBGH3tCJ2f9O0dHlWN3sHKuPgbHDrtstlg7bl76+P6ckKvX5pX9L
bR1ewQrvX5c34IfpFpnsYJFc8kSYWcMX5xjDplirjcmW/PkzTvi0IZGMqNKHJx26
0X9wXQkA+b+39a0AJiRkslpDNWyYQxZwxgw/qWfo7gvdfXBv/h/PiulkXwiy2Ksr
oqA+feuxv6jd4Bgr006GErK7OcJ+qCjb7SzOVKJgoiL1o40xX3+geGNCsnELDRig
1plxSn6uoa5fzZeEhskAOE+GRGD9Xd+GKfkqzp/fFRr+20mZV0rqaJNJ1eP+ouBQ
W3yMIhcfRpPtbSFdwyBNbqOOw6ZAn4Owb2D1H/pIdA3Dxgg4qOFDTaEHMCJZ5Pse
MxE1T/wrtT4j/jo8ZuorL4dyYNzS+Iq5D/5nUARaNQ5tQbo+C/N49DURLvZ55dHg
dbud/lyVOATtjzvFKus3T7uVcxyIgpuZ3YEtyOJFrCJ3rk3ml+ZcdUVQEaP57Sfp
EMwtOd4O001NFRX9Ldq0r2RVHDaOzBOHyKTT6J/dOQQO7zP9rkoTBu3c8MALlx6i
6ASp3lCBgzqYwGzfc0KQzLKVshRrKFsHMQskI+FTqzarVZXo0hurcSySKBHlQxvN
v3BlGX3ccfiL5AOsbshULTGIujLMRdr/N4Pj84b4pqi+A9vWvkZkHWNjL5p46VBb
IMTE4EW2wwtKdUFP22tLmVSqFuNOv6sDv5FccjCaFD5s+DFxp2tnl9F87e65gb9m
hdI6Y3IrSjTM/THExlZnHFHa+KM3hbNs5QwYBBH8fCvOq5cn5zTKdZ+keIELUlnp
qbMIyBl4prIjdP8T4YoJKaDMvk/78boLqu1Igym+YkFYipBFryrwr/aiK1lsZ6zd
w9zsVORgSDFdgIPFEQKX5NtavnZglaZ6r5eAOQ5WNmDBnzZZyLLAqHZKH4RO2yKF
qDgA0U8ZTz+wMc242OuMd5e7z5u3JOd4FX2J5KZZCHDd3ho9V9KuDFqkQY/2an0C
3koKQBvJ91oUvZoAl2oWW9oNNw+DIRjEB7ZuTNmeCeupCJClvkGlCgYG0EXq6PU4
8Gu1d43hOqnSmyhI3TXIduMmYMB1rdnwdjUU+6XY/9lE2U1Uqdizc2JtxbpAQZw/
+awmhw/7ToCRgTCkBILCN+kuL8peXUJFjNjMbGOJdwNp5Dp7ltHY5p7zf2wQOAME
Q+P0F4DyzBz4icZ0z9nUw3PytgYDJOKyfckqK1CbKQWMAsNMPVle19Q2B5SxBaw2
Jha8s/28TBzXRVAIWY/ftaXvvrGOL9wwj4CB3lC57FzgzOSkX0P9EcFj2JFDLoKb
4z6epKpTKssi8TmKggXkdaJ5AvDw4gOp4OZJypCKD96G9QsJ5UjAKYuc9TTzAEbV
jqz3Bx+8RLRKYD0avMDla0QFDmWM/THp5bqEd4PJPk/wV4X4yD0cYYSZBYd9ZN7M
D/6SMzPSgu1raVtd70xIzaYyXekPM5tO9wmjUKHNiu09SPU0Vjvzvt1lpiYHkGxz
fzsZ7VdpAjN5Q8WybHPQfRavNeE0T93cq92qfUvE0tPVvn7lHUAdPmgBnp2RAoRA
X6Tqs52ZcSTxIMLHWKYYBv5OXfO3L3iJ7W0i8V9nue4pj8p7O4EcvtLLOspzE8as
kRpz9ijGWUiTndC65HnvlR8nZAyWH7hmfkl8tAtkvODJLplhxUfofSyrtl8r6rrf
72K2MoGI8nD3if+sZQ3JCAyRdg2fZkhY/xcgZdlnE4kzNCa+75vjH2m6bcULsn8Y
bYOZCZYWQMoO0UuW0kg5S8EpcHQrtyNWVXopRQtvzG72wBDZGjiR9Llxoxb+NxmX
T1/tGeqANboc0NFIDQ6eu+vluVJ+rliZT5Z9vnXMlR9Ip+nhQZAe1VZsPCTUsYAw
3sEM6EvFHgdqyShY4jawpW9tNDxyJNZ7/A04rxFHMide39KhZObzGKnMJWbA4TsY
DbJ8AoDAkN41T99VLTy95+wPtA5k9hvTFScqpVxNTo1ZBz/T8MSvnEPWqQ/XBasu
IQrdBsbjczy80fd90cFqvTVe9X2x4HSLj5RjxFRBPgB1yFLHcVgX1s1x9ojmHhMX
ZQ0rVpSWGdJJocFjEkC7cJagoAgwUTDYhkeCdD1fftjNvqIDvRVvNY4UVNbI4pm4
4HY/8pxUqs9AkFaLqBatxWeyvwqqkE/BUBRNPpEYKZf1MfiVraHNeBoyFBg+XaBc
19wWc3lEsWuYXwHePa0tbW95lXSfSsTT72hdqI4U5R4+lnM5ehP0drBEDAoLecbv
da2hpltzMBzKopAZegxwUDjdXK/zN4iwYykret1BRnVwoG8HJItgHnsP5iv023k+
BH1RFzXTUXLHaloAVY/rdSpc8NkBCKPqANASGZIdhRsMzyndJFTZOSW0vXqgyc3l
qITtuzxBlzaOXbC9iyqELw3lt4208PaK1L5oTvStK4Sbcmd1NlY915OGtD3cJzgr
mZ8r57aArMm6hqkXs/r6SdwbFOdoXyvJPjqd5evbSUphqxjEQ5qv8Smg5tND48Na
81fQElAQvxPMgeANmT/m1EYcb6JEqrxmb2fFi2w+8Fvh9lGArOs4061wvTCE+pGs
SoXKFn9ge7NLLIlJThbkxOi7uaVEULETwJ5YJgl2ggqMdhrT7nOHE+PcqOO+4Ip+
gKnkxEZiLxFUtQkii/A2QKx3mkGRj2iDVPARITSARJXm2ERI7Jzksu8PBXhjCJfa
BRDK1r7/jmWwPyLUz9o9jBXIn8U+Js2QKDtGZS874h3dVwxpCOBzTflCgkQVb/cB
8h3ok+ZGR0rx+gC6XJhlzwL1/GtNzXiQuG+E26ZdqXtylVm2YoH0OM16h9jaWUo6
QYuACO6JG/ExvWxXNd0q4jcVjJvDzTR3hQ13ma80HDFICqrOfdkMxarvro+rmC6l
2S5sxeZVt+6frBb5r22qy29Le7JLlNNrV+2WoCwlnaysgQv9/mKmlsF+MBC1GzxZ
tEzDHzCXoQR+C19AhDWw95QPXUPNKgMcNtLHyE6F25vcit8UHL55aNvRwgGyrfG3
0TKZk27L6DWIC1RwT9WOiUEvCeAJvdVq16q9KwEFDN4KUTF/rM5Al0pvdq8Yl61q
c3xUVcdNbAn3qrV3x7haqUfCS2sSHzu3fiCZpWJgeAHJ9UyNCVRwKcMErXSJ9tBr
JLXt9LryzwDtdAEHtxFpfUWOb2VlqzrWCqXZHjCSj2E+N0wTxiKlmu/uDbzkWMP1
prGkNWPp7pojdWPf7unyXzGFADu+WNxQuYT4zZTyG79ZE2+u2vMowpC5oMHHKb0f
wgzhTmpLq6RxZw15tzMuca+r/ZnvTbmO4Uf+eMVwZLIveyUvfHFq20A/MkD/ORV0
+UJTBvdF4r/S8CE0dYOzlc8RIvlPgILF7lzNYbDcRIYxTcv/wByiDtRMYZjfWdGI
V4u19CQN6hs4Mrl6H3nhZ1QZfgF0qz3+fcpoTlLFj7iGX+YgbieL7jL2gphTsceY
A22s6IVg9V7q/6ywKdapTlBHyeY/Rs9h911HWL9zdLPVJp4+JKQj+FEBxAJ7S+bq
cvPJQxUU0b26zF8gRIH1ZBMnhCD3HrgoOq90Heh93SMry3RGdyrLacg051LX3Gs+
BN7EbOsO3DWPf82iGHHs4ucnpVtOqJth6fr9L9hayK3tKERWJNTyXU5zJHtyEity
jYjB8n9zmG9LI4gYnj8vRBvG3MRgkHaGdXVt/gYYgymGaa8g7BxHHC2wyGdkvpA3
7FIBJcxo+cnF8bNOOaE/IFgU4fc4a/kHxklPMsZPONS/kFTbPyD4ECcqS2Y+lzyP
2Gp7adJs8v9TyJVYXjPfo0fxe7orlDLC+98burAjGyXSFoNuWa8d0lOsRA4F1GHA
1tTtoM74jtD+5AOxCGKEaEOKwuGAmxctJN121FJnBysVLrIV+H9eFdLJm28CjqB6
y2veQQHMCvfuSClrSvkV9JLG7J8RKfR3hcDDJ33tW19/ToSbBWLLt6OvruYFUVMH
EYyIA+F8Sj7KLhQ2UNGIVrZCI3Zgol0nb0hdB8OagwibrXZnhQ42vcLZU8yFVLx9
Owo3i4rrJhIozY/5xgUAtqJKkia71RJpbbL5+5PhUFCIIlbUbn4z5Eey+fEcnBfe
U7LLXGikcARvsoYqdaR64CWVy82SY3iHOK141sWwH4Z+69RMml1ANwzVOqNEP/sR
Lnxyj/akY9sIaHZ/rfQPMhs27FOx2FolvKxZKFe1a1GIpUxcnrCF5uRHHH5jOolQ
E66fIXjEgeb1mk399ioM7OAq+Z9PFAl9S/QdSfcM1q9UozakrVD+YPFZpalpuCFE
yfqUOK7b1/Fs1bc7lWlVHJQbYCRV8/p3fitA0fAtdRX2G0vQnwHrHfGRig/vuTYB
iFQzP+RhoRj2neYpwur/gR3mqKhWHHflNfAefli78MouzqAGM+CYJbIRtrkVOed0
/km6dvZ49XLFeLoYl4HU8Bip37SGlEicjidx8cAaCLtVDLSUSucoDEwgp3EL5SYf
fG/Fl2m/CQc8/vtxsuk8Klm+Qi2lPhXiZ5mJsgvJQbQtPNtJLmwtSsCv8yFFtc0+
sfZSMFhMXWlpB3GEVj1UkazdbUGwiEnX0MV9mBFuGO1bcsCC9OPvppIDM4diVGdU
GBsA/3YLSRquzLzLRfch6sNYuDt6yvRRIrE0suZKWnI2vn98STNwMaJFQcJGDUse
/uuff4ZeW3tP1TO64J6gOcIkQI+nUZG03b4poPfKhHT7J0DieXr+VQCZchLzxCma
jqMK47coxl9GBijp/485bY25tLwfVpYmh/rV9seneaviUdeLVCAGspDRweNbETd+
WyH9OSyXi1VaT4y3yh8bSfzs/R23Hw1YwIES0DVDQMqLSVlSd5XoqD65W/4xQQ7P
phkXf+j+jAygjT9dIldhC5WIxW4wm6jFwNPjwP2j/yMivopfwzOwLNU/tv1BJkZK
CtF+rNUXIsRGn+GOMTPVBJO26A3vr3iMlPjBaUWp2GucUrexWcwApYNcIO4bnUoA
W9OesIOsbTJeRTQg9WAO15hOPDmQw6wN5Sig1GvV5UmzlAsCVlAA3qJin5mtAYSb
KC86OSxiODOoDcmlI4Zf4PubtqHRN701Os929RFS7lWRuAtnmARDSZm3h4qBN2KF
TDmYggpyTJ5q0DCEPtVIF5ozptpmhSWjjK1jkQujzMyOc8LYI+LO8iZYm7VnuurV
xSMVe+NmNoG6PGc0RB+FLArPtadq/o3bYGkRapgyiEFvxRqfriFWEuKgI2EVdXAm
6buHuiJfTpS+jJXG+4BrYBFYvBCRKQD3EUTnxeQgX35vbZ0x9uTSGYl6APBwwGII
TeBgbBMmL5LNzynKxKRai7fYQpggRcWFcUPNQqMcyBfzXYiXYVqH6IW8mw/7T2qw
aioGJYUVgNMu4H4w2FRkXLziIAQx1aEjE9egplygomG2e9avRid6VuLKd5weWZMl
G/4q/Yy+ZtC+tHawOaPHfBf5dYr65TQyCkOuAMHBVko7TmVp6XB4TW+O2SRoHqrZ
Kn+Df5SV2DSmUEyJUqqvwie7mQJjPwvthSchDOA/nqfCcAkUFnA3Qo2uQL3AgQ/V
hBdjjAmDbAbLVTSwS30jLuqoEat43dsuAw7LeZ2goHeN5myGg1LVcNqLLig94G43
4ZuL1Gi67scVsYEcn7AJag5XlOVjmJ3g2TpBF6aXjiWUWZAKFjlx61qSEwTDJdBX
b3YYF+1QBGVPv/QQAP9mtQNx1E3Qp3nD2jD98bM9fnYQm96zVGfbx97HtwdIXEBk
sIzW+KC1oMS9oAundnOeubtSBlQfmGHRh3Wyrs/oFVD5tMG9BnwpQOzy6iysB/7s
7zheFqXPDUQqYWcTA/SoFs9pAv8zfvi7iCAVZPvZIj+Jb8xRBhbHH03B09lYGJn5
zKKmI5T9en/Mb6N08BK+SBDJG7o/495/NHPjdt0uJb+fzcPoKBfqw3Ryx5fgo/sf
owGzg0vz9/eIR1VSwjDmGMmkBQj7GKb9gKOc3Uf0rxEg3ylIycoapuJN5JOhLl6Q
g180bWwkNdM4Gt8O2jvlLhDRIDWg5QPPu9W+S+Ho4+jDUqkMPa9UaK2qATmnAdY2
cOMS5sX+mmuEsGf4/Jfr3UUXKRKE41AIXGVL4mi4cqwkQmfe4uhedhBwOEIEb/1m
zOKGkGR1TdTehqjCZOkLXlAYgp1qpRa4DmhShv3ABG1DX6OolPb6q1/6XwhQgAWZ
ub18+CiFOw/VJSJNW8N7XhPSfxboT/PYWPiILwttWmdX0+Fuj3a5uNsqnfRfpdQx
ujeZ95AY6RtRz37v0Iltpt1HIshTfSw35/VVr8dW5O2cvKhjJDtvBa1RE1Gpho9X
kaXaj7yTeFMDbE+54ffedzauNjFy8VckVd/gXvTQzSEsmYcYzuEJq9Ej1bBJem7G
APuV4GDq+2DY81xlTSfA1N+jybRsy1nHJ4+1Qw5o0Hf/CnffnAc0vdb3KuAzZx/p
4FeBaQ0J4o7mIzFdehwzhaPYpHaFmdJwmzh3WZw6tIoZ1772uL9GFuold/uMH1DO
ezBjjfC+zyBH2gDh864hZqEOFYuXTiaFoVcS1rbb2Q2feZn7eTz5YHQWMUTA54UB
3BkSMDfHfl38Tpydv3d7E33Nx/WvlR589YDQfUHDMgEH9NRWt++CVpc6HMN/Io/f
tG0f1BJLsLBWNcIDrCltianlozTWOXiwAaqUEmmOd8PwAWJyyYGPIuruoox7q21Y
cNQf7s6+ftXGhyeW3PdWMFj5owCDV69/I2Sw6OLYSPmh7Ux2PkdmfePK4WoQmVql
jDyr+Y52aKqGCm+uWu8bLlLLVN1zmWytiIeslTEp16ennJCjFsmnL6VybqXjQ9EB
wtFzBx+jlFH9eZSFVeZe5CIAkATGXWOJAcfHFnv7IpELkniKgZ7aN0VxZJu7csmU
OJCSZVqn5DTnBhALaZ5U2zU5eUqTm4LqoH8bNQo0R4VkciCcMR7EF6LYpwWKb/C9
jcGtQyBCH8yeC95zwjfvK7sW8p84o0BCuqYHISmoIRnRwwf632BxOsgMmf2VJieo
x/XPIgtbqoKAU0kDBOo7FZy6qIsVpQm2wMJwwucCMmRInrnRP7oUOThrxwd9nslZ
Pl2L7Md7WQwo2TIBnkGi+DPyEsvoFRw2ZSGq4FoEgl/EdojtkcRdT4RdaTK3BjzH
KPjW+DwzRY0WT1U9onFcY3d0kf5XCrxJSf4lJcvSADQyR+v/5PfvWGmQ8kKNMKLC
lvFB3Q7TUxiQ3yxc1Q06rUG9TOr5lhriI6hu/t6eQPYS+kVChegfw21Aqvre1H2U
hDM10PcF9LtnH1g4rYsw3o1RobTDna3+TAqiD2t996bYjPvvNdM4NSdjJ/aJYt0o
b+62VHmrcF8+nnPxSP/v7NkQQOaRbeRM7l5mXWtpqrwzT96bQPKGO8VYImCuFQLp
PH6vSKvYp7gLkw0AXxicSG7VXndl2wQRHzJLiQZpDruiAo/fL0WHCNhCtQsReiey
4p3vvhz3ReW2Of7cTAN6kVnvgIeO0MJgLiiB8jShxaLcOauha8SK/tzpoCB1wvEY
qnjwU3qDgxPgVn8b2IJTPDcaqeJuIouinr8vkU40guA+HQ8SYhBr4TFy8bsNbJAl
ElfZ7dj+ZFk6KiyQzu3+EkgyNh5bUd/Y5aIsG6rlcFa/V/HXItDjhoF7ak8+Id/F
xU0pNS7LBVSvJeNqXJ6xqAXUfYuhVpqBQgXNSEG7fSQaWi9TfnNFhQ3+zN7+9ZFq
YAB5OBzJCpV05Po8CYSICdzpBfeJhCnV74obxGzPh3g5eBvoffANwF/GY+syGxQf
AIaBq6iMf2QDwkc/4e84QXMP4e37NgScXA1fv4CoIKihhLwffm4loSvxwT03LQeU
h+lqZNxe+kgwoP0lmR+i3wh8sxlF9xNkqyjDh+AZCqUa7D0bRKsBfN/JlWjKNRSb
Z3Joteqro0ySRuU9o7LBfOXHBsSimxS4Xc1vGULUlFfb1FFJHOCUfR5Acxt5a6F2
gnQmozWhcveUI2um4aIqEH3kNLwjKVleV0WhnXd1V3TwN04cJYbtsOunFfjzjJ21
2OFvfPwDUTL11Ucx72kJ3vwwSgrAhat85bZ7RqkYIRU7lE748odOmAuPKLkTBXpY
Xb4+DAvGqux6iYfjQ3wXLdZhxPXglm+sIIhgcBAHnzm/dKodO7JS4DFQ/nyz5teU
SgUprqOeq1wzlRCmFDkNMObO8lQ4iamTSs2HvoEE/P67gI7g5FQTJfOgSqUA8nJ2
o/pUj/DrPz1MzrTr7SwYDR63xvw5dacX6a1jwx3CP9eRy5lVE5sEt7uWsdfoafbK
yKdS6wx+7C0MoP/DzKvSmaXIGR4tgeWNiHFnjRMZT7ECm9Kbqa5nJjkagxAj0T1m
rDMp0f8paYLvYvrU8JLxODDLDz2HKxdqNzsDcjp3OKk/1ayaClMnse5DE/j1WzqO
HMmR5RI6ZF7rcsxc320vLuUr13c2t6ddbdZ7lQE+V5gAKdJA9SRlSuOJQbDQu4Xm
KKJgaTEtKShbWw/NF8/3UMRg6VmicNT8MXiVtDrf1x0ayo7tM6siHEbaCwXyJqY6
cgMwIHUNbKjzdjQ4O4o5H6hqtgl0Ln2KXhZ/PtXnlfjWmIoP2weS7kN4KLSM2sVD
+MtubHcHeipPnc96y0b9W9Jlmn6DpdOe4sx53QVba5mc4qJCXGASMfnShBKPAsdg
Ilc2YB7ukA4irycMfjBv+P5n8pBT+Bluj4F42msLRYnsKU+mG0v8WXTEGLRVEDMJ
4ELmfNvJYtQ0M0W8R65mUDF1m8kCCceBHJLdzuSMZxJOmQsz9FSguNHrFUop9hQe
UhQ9+8r1F2fN45MUx+am6ciaXz6j5VnqcBhUxQRe4ZurXmo3WoRLA+EpseG9x5CC
3B1i8VRfgIHDmWbqhj4AwgYS92CcXJwUAJHPND852bDaihTNOAZ98GmaWGLz/njS
52E5C1t4/7R7umV1s3A1X+l6VnehPvodUxXBm0o2BEg/u8LYrl/26RRHwMb9kJID
l6//HW6Y7m1fdO3b06iOphsLL4+o/y5yQbUq7r01OHwmT8WHKrCHfPxJSATnBFfU
l/zVuU1mOgnPmtuS4pXfhpCxcRyP28M7ZDHPBnNzM0+inVvK5ETZ7Tgc0lKDqdsG
bWS3Ya+/wl8nSc3GqcD+J3zrRmQwRce+Mp0l8zBEltfax4MnZq4Q5hWwEI/pG/Sy
pvdeMcaEjLIU8kQuSqKPskGMKz6pCGg+WHg6kHUmyG7ayjOlUjN69t2puWoVckYU
WZs7wA9oyURp+Byw70FmetrDPy8lemH/OF5GrYvhXosZQV2tiY6iPFGcJwKdI+ys
91YwBGvWfijrc+dGknBuZ7tRa6ixkTVmBHqAzHhOq+XV5F/w67FjsjzkrZbmqk4Y
Ts97/7FtNzN0UPAEW4kin49WLZJpKjrajXLzHGYGj1R4m8RmE6Yczjc1B/4j/7HV
uzBrfgJQeTMnidr/3p/m5PrmTayTdErSLbjoUmDf+O4mjetOBbV0Z4/pahZ37ojC
VqbJsCxHZcSuTfEzVM5gzZQ+Pa/SJaTtWerVuYa5wRfjwBnBrn3/SDYWbVvnOMoW
ooFhMy75VvO0YGQyIlj6G0IBUaWsHaYlm38DUF7FPXA3cVw/crQK7yKwJrWbfx5F
XiDBVtMirndY6i6mN3fyXNX5cJ3A7d4azg5ECRxBXZRSSTzXE3FCFAzSvyKPpTHj
BO8/dSbO7/lk1nVCm2RDUYZ9L/X/l0LssHVtyUmZxoaR5XNS5ojMiG4c13EXUhPA
gGLutgCRtqgPWa2QmrMK9STsg/6TtE9XIsq0w31rVeq1RWRqyHMpSTayA5E7NTej
xHVm5G2S/0jmVrL+YddDLB0WP+9HHWOUIIHAZo1rVMmoKNWckqFb22ENTVS8Jq2T
W3s72kUZS3GctOux+3LmeIIkzL+3N2ckEI46hE7iwUVhlJ5nAUxb4fTkRqgPTc1B
6qdxyi2W92rlIE4CNn3K1ApsJ++E2Yc7DceIgK2/d7S+9BPHnyqOG5gmkMma8Pzf
SduDIwPgtRNtOrfbSZ90BvqHu5h8em9hUZSnMEp0qUrR5xoSZfNXBT8guosHlBWV
pxjoU4AZiRWmVGL4qGYHzC19aUUPMZHYVbamCznZHtYUjdahVI3Ocpml7w2gjxsB
xa8BGVtyCweyA1QlnIf7nCsUGLRnHeYQN+8qn6k3wXo53T9bhHewXhkDQc35usa8
gAaX/tsHFS+FFHSWBiYupVxXJ2kD8ollRvcpqqP0vt+maZvlxK+bwEWxV5npXywJ
88FkTDx2ip+L332B1NKL4NIU1OwuiWylbIkAn+lBws1ZRheqHhYLfLG3KU7Bl3/q
ORVQv4ZsEkaah1j/JtmvKegTTJT9e32AbcaaJZGC8S71CA0nQEkIJL3+6yMfYd+F
yKDQcQ3uwdSQwJs/0AApZhEKJ85JiMxevrkmtpI1KH/6LbhVc6QAwx1OEy0Uca8e
k00xPPU+xBvRab2qdcGZvIY0P1toIdhU53sRC9vUmT5pQkTHGPshBUmgQ8h+9Mlc
uG1b3KRIBRAoN7GL4pRW9E2Bez6upSvxh+WjkDf7CCouq2j9MpoDubiLnG7vsE09
BwGH//eYu2QSQiRJRhLqxTrCkQbxoiw+9OcyZpdk+1swo+AiSQyucMOCEa+ONEAw
FaKYvctsQAG9aGLXohsRG7ErMM16F4cvNyo5YHwdXrIHdiC+9zMKrv9NKWEOBIzD
8s693RXMSTXN6mJhkI81ib64FIUDkLN5uRFvKhRPpApYwpkTl3MZj144bWzPV3un
A+u+PZeQV4LTblfYSVU0EmjvDq4+Cp70bbl9wFjxfZ+q1ZNLt8tFBdH/IlhGniRA
gjbh6OXNeEblbtUMfFvYX18YHw5ApkqXkeYZnbadd6gWtKZ2F7NuurACom3sEKd7
6UkbM3/tKmaRH1NqjGH63/2IyAofdWqsdx9f3mwMMpltYVniHY/CI48qSKPu5Rwh
kYitymdAONxBBm23ZVVP4xeE7MyK66C5kvBQUi8+yb5tH8VWHGZhuPGB/PtXQniR
1zBS4sZIuBfsIKimUugka92Fb2RjGdWXK3M55W+vEdoltiBqI/NOJbsxHxToQ8ls
xURhdg0/XjoA9bgUStGLSnz9Ku6bpg+3HGicI/bJtJxRW6mj4zRjd9i31wCmbdmv
ESf+e8oa98YjB9WNF5R/pD8SuNAgLsc5/F/fSr9G41NqrPVXYt8Z1DyaKAQEYVVB
swQJ3zwjczIvvbjq3AHqGhRLU6FtM/itVUhzf1E6kL0lJ2NwsndLbmYewy0jNnrB
UvicM2rP7kLvCLajvg4ka0a3maoKhpoELl2gQnrafclNPPT4fmIBTZ/NcuzJmNLD
t4gSukU9lh/E4jnjfvGPIeOSiVc/lsr99FEFSNK0EmZnknQHbJhjuXqU0QEFRVQA
qeEfd11VZpCqafzUf3BqgAEDOXTxj+ftUfFlRHXXwD2/JazIzidp85BV6jUZB6da
aoNZ36hUgb+zsES2sa6b1xhRENnDK4l91jCemKvyzr9i5J5GhbnO2sKF7yz4NXwq
2PiWp1IN5FqCP+un5D/oVCIsffLa0fuXehwcNIMKGajXztmO40Yu1cn31Hk44ksw
edNunyMXIvNVoZ2HALRnWTHuJ886L+mVD6HYk5CQWMyGtGZvVA1Jtvc0iQ2gsSuc
qHw/Zu0sjs/kxtzT+ucvJKFk5eIOe2so49W23VFgoxUKHBMrNwlum4o/cSktpClX
3lvUnOwkdRHm3RRfzeBCuIedu2A2jva5x9wzSofvCqhHQ33bZxVhbSIcwthz9yQE
XVRZIUj5jZUNhj3XnkYpN7ZCC9VOxdmqy9VPsHwzxQfumxDZ4hCAvQBw7fjsIbTb
SeVD45HoYp95JL0Fxvrgc1r3eEqfEiayiRnrGuvFjVMuRjDk5JoDp8VLd9C6W8fZ
7C78I4RVE5Ac0wj2zJasAxFU3Ahy18in4ODAIEsduUC71bUoqzDrcpO42TsSXT4F
4kNMcUkVnYBIrtMbHsMCMFA46BxdV20tFRKEzYzhuRwJLKuIbHfyscJswcgeglqG
7z2csJA+B2Xt9RGZ6BS5OQ6rFcWypgRtM0zydKeuAVaEEXRwIJssVP9FNrxOJ1ZZ
x/KykiMQ4TgQKswMPv+gH0TWujrOjRu/1pSAqELvvsONW49lsxgnzejGn7qHgigG
PCapFWv/jn8hPESakEq42gtOGT95vtVjrepGvGcQmXeAlafzUly151NLg2O3qhsy
sy9rEdbRCzELbI3HbVV/9DORD4eAKtUpJIzcxmZzG9T159TPCunoat0juMCW9QCO
W7OJIjkZCQe+8EmwPWluSF023a9CKQG8VNhGHMabFjK6prhEWsuikUkOUyIirLJi
r58kvRx6OZyhP8UV5Q6e52NmOK735qsMTGDDkSMYTLd2BSGIiRN0oGgjLSet3m9G
47h+wPejrBlmBTviyVucqCaQYmL64XGIH+pv+D2FX4htDhK/EkQxsVW93FtvueAo
vTFMVz0fT8PZfrW9qq+5eD8IavLLgAFKmvlZ6WDrcd/so1IhZ8Pp2PNiMswyuUbx
MrDlFkhECCgtwZ+OdzjqBsog5vrJuq7HkmQisXorFbRoUNE7B3fF3rTFi7Gkxz/u
E/CI4/vKNG8duUL9F9gbKcjGQuhapGxhxlTh5nM2QEyf+bqvJwIkrgkUpDP8/gYO
nqVKGzmqu1LktMN/37l1PaPRW81737FFCr6vRMVSbGGBwdLUTCf/Ia2zzqjiek8Q
8rFpp83CNSPay5GMTOxtkf4d8ZyaUD8cua2HY6mjMdfUQ303vqMvIshB57F1PmKr
KXiFxDivUqMAO2UOdnIST3HUztzvEuSHLT1N7D8D2ZPgDm2tc5O4M6FL0dVB9XeQ
HU3bAmdrBDb+HMi2VvzV/XrENPF/OmoQOrNM1CrOzX3UoJEH19MpABbrAF2KKQlO
Prp2ekpFuhfGVF+sewbeeQXXmyETxEwgLvX+zyGvYNZUz4goDxJAFmNv6YU5A7zS
AVYwdNDlFzRzznrsgB/umyas817ubwu7/+evoU1hgTC0bbu9QcPc7t2+4HCah2FO
xuCfCGIqVxhmxxLQopAftt6yG7HAWDmMKk6OqEGHnNFIAbD+E31fi0CX/m+9miae
vptHjTb37PJr0CczYu8shwnn8Pc8rM7vmO9EYhlfYYCiyb2bVWqzKVD58STuujBq
iKz22GtAzJUOVXUPQVaAo6rcwHS9sNnKLe4RAZ1+9URrlQ4nFfq9AyIBIAiZ5HEG
e1+LZ3Pbx/lG9MfeMj9VBx5e9OtOUZcL5YeP6hpAlolwY2yU2vDCZuyet5SxXbI1
2scE8pEYeKW4ZDDqtCD1UejGi03LEGHapyq/cnLS5TxrB7bMIEImfB5eYvkTFOlJ
fB0tWca4E0T9l1aNJdc29udlDj5PjA4SaZLQMs4ElRziVvi2J7BL3C4ONPLsKun5
meu/2b6l6wb8bu40ELoKoK/ThlBUy04WAmSDhnXo3ih37U8plhLKlA0miu/APMAR
HNEn72Ucy1tGWGsT0cBBCQTAMk/wYn5iYML0Fqg4RauQdmHk8WtCAZi68VAKM35W
UFDwNn3cJukoRmXgvMtToQqEsxj1n1fGSszHrEYWRYRDfKNZqWVEx7+DR0L0MP+a
yPRLCQsnMs4786bgCFPBQmS4RiwRw0MiEqr2MqnSgzdyzzDS/v1veqFEg/FtgTuP
rBZkaU/faZ0ecqW2f2gd6s3WXhFFOGMMSDibynlSdvPOdQc1iUmeCKNA/H2ugrXE
A9ORBRU5DhTrvHoTLbxFRd3MjxdzDVE8JedMN7Man2aFt2vduaH0/TfXiUdLc3wk
p/+nLumfZNCbWToU+9x+cOSyFyNbe9QZcOfe6DLU6/oLTGB9uABvJMKKLJT56eTq
vJsYrT+Z1S+JTcFphdyvGRz+S+8/6oCgEgZlBdBw9XW2E80mJqFVghADHYAVnVCX
U58oLkCMJJEWMjC55l/c70itz2DvL4n1OxXOQohaa/A4JTek+XKNvFj1NCfG6c0k
OQfogy3d0lh5NxG0cQ5DbumPrarbdNJIDjZtqvikAXP1+1tpTD8pzNRBrZFA+0xW
V9o0Rz1N1lJszHx2KlKLE75xz9COCjzaL6HvfuWQCJm10JdcE0iVKqrLt7K2A3XE
h2mxZgy/WGOLNCTnas89K0+Tm2xgLihqd8jVcchJRx2mKbpwVWM858Z6DO353fb2
dEBA2xbaB2LavdbdBlj4pS3GTkQcDX76hJwV+F+PVZws+1DTeFA22wK3GCpnYpKI
C+hDCWFD2I4rtERaxAtdpOkr5B7Wjs82hbcsb7KXjwixSMIs5XCU6KO2Z5OEDKfd
DhThwfz0Edwc9FP6p1dzToBZiNK0buOOurUmXQo0udUPcfZqPZxMNZZRSSURWDIA
Uj6IC+pCJ/DWt4yur4xD9NffA8H1kibvZowvejQR3CvQdx6cVdgfwJ0rszrX+imq
14No5X6MBPiP22GwjM4Xu2V7QJpmFuOS6DUUUhc6WNetL6tswkzchPQ6asqFAdn8
oAQqeHLG46P7U86t8/h2K4imh5JSNTPR4ECHpqBDCMKQ45CRWLFkan7vW/drBk+W
J/Ea+lU+0Q+632pHtf76xKW2tMzCN6p91cen9iXets+CFd4tI5BmAf9hwkiE6yVD
bvJKrnwwelZ1upTnBeR4phQZhiOrOPZK7YOa0948o5kX5jOM/Yj7szsYKpAfDaVy
Je75ks92yMNzryJFT9Weo4+KH+oncOqujFhI+AV8K9y7FZ3N77f6iSCrFEQaBbOV
iuNKsgWJ6CwThbwW+pADMWxHYGtQYZfOtiI98vBNGaO9Edec51SosHVziMZh+csx
rfL19nkaKFV9rSGkiPv/eX6j0fBJLNoancTJ7yOaaV6Z7rmRmhWDdGZxvokmnDYM
zqQQd433/J1PiV7sZNd+Hq2d69BVJKW1JT0wDsX0pUbqHol96crsByhpPOH22NQH
wB7X9ySNvwkoOuH30iEU0O4yw8QwIpF9AwfVLqIQREQ+ksVMUhwG+b5rNnbePiAX
GNYjSRhrvAO09OCyLB5TrlkE1xidIxWOENcx64BJigigHgBhP18w68H98mm/pr+o
kNyyrwPMAae+StbZtvv5k+rbtf/NvJnfkzawvwFOXfvIk7Xje5bmW1wy3wW1R1jJ
kZa8hdWyupi2u0Ny0vL6tw5AFVx41eBjuEGxJkPf5oMgFzPhVGkAk6jQw4Frq8e1
QXmw9xb+fFgxXOpWPp3lZlbngQBPi1hfrTOOfibidAj0QZJuMYnlZ6uaEWfEV1UJ
d5tHrIq80sKFsI4ml9+tba1TOuuSg79cRUzmesb8UU31Pu9im9H+STat87qHY+Cj
zlg5LAWmRq0aAmtdI2D2ibKm1pHoGgqrYHxzhV2zskMxI2UYsiK3tzykm2RNk/j2
Rw7OWFk8IYvTFMUrBZTJmSUz+jArxdCkyEn66Xa+eF5bpP+LanMNSrE+Ox3AaAjV
eIoRscYJbqwpcmfnkgHydhjRR23sNW8+6VlyVyxht9k/ff26Rp83IEsVrN22yv77
t330YDWZL827IXmElVJGclARuaiacW3uEduGRO9to9rvumi3QT+ZOVDKZ7ZHc7L2
ph5/TKZpYqkdvG+s4jP1v3mV1djRjokRydY0LKFn2m4H8rgZ6BsOC6fpbhjYlCSu
9MK33W9EzQYCFhdSokk/3tbak1cweHxZUGZiKQyMeNmx5d5IoY/zPdumdA86kcLz
jMQvE9lofQgqDPUAnk17qNXFNgiiAhMaOgw8740MAaZp2odn5uHhH7KqyWjCRpSS
g2krpB1qPI6y9HV7/ASYLSm1z2rn2ThsC1qcjeoZHdzg8GnqGTELMJCYS1zfJs7C
6SZxPVdBkCDS6iGS5T67/mYmW2WlcrBPun1ixU2YQVgNCT/BStwUEVZHyzbzzcNl
XbjP1TarvvGgzDyDa4yRv4c4MmViUVOzTnNzf+day9q91WSEEhLFSJ51WxpYDr3m
IyfaP7Fe9VFjwoDeLFvxrb47ucxJgvQpR1fAPo0e/CXSQ9mt2eZX2nDarlJu5kG9
s1qzHDRxxtMhEfkYVEl2eIXa112luOX0ZE+kxEfHuDPrw3sgyU9nZywJoqPQG4T3
bVQZprW2OaFauGKqXV/VCjasdNcIldEN6SltCa+gVYdpRHU2wZbuZu/OzgElfypx
d7Lo5yMFNvKfnZB7P2Q2KCQ2leaBxBdo6CS2LFttXXwn60ybOHpxZBlNn9sjECoE
DmUSbtNyEcFvXJvFRgPsQa0NBKQwQRpc0GBfdcgq+PDw7IgUIQJad2XxG8wYLgDw
xcbUkej8v73b40BfNKYAoBCZdgH+z2cUK+UuADPtFy+h7lIiXIDxLxM7FPBtEGUF
7tcN45cDa1V17swmLDUWvWPLRiav5UHAijuzvogKgyBQl8pdSPMflrzA7k+ngE0J
RfdWp93XnGSC6acAg0QH0iJNlgiUQynsa1VO/NL0teFmCGn5LcL0Q/o/OMBu4va8
194kniATriq2H9dg99d4Amnw2fmG/BakYSJacKil7OQd5+O+NbxQWiy2eHr3Okl8
2Yeu53ILkBIPCOG49j5lFKGDTtFjgYzluecrutDLtBmGcFc3fw7dJG0WnnyVSt6Z
2Jm0FIbPsP+opUi8Uqj8lict186GJF2Vr6nYKeOT4AW8Wzvy479w8nhziuWN5ZER
Zg8K7b8Il7DLFWSrQKaj6bklHung3/Wx6sOuWiP207Atr2HDQlsHBWgIAxHyoMGe
g+V0b+2+EnB4mDSuUCPHcMS+IuXjBRnjOuE0YhgNrIBT20U9ll41X/LzdlpmSKER
5Hv9qo4Zz1cy/8KgsljPES0vJuCxZrqpCdQgdyXEBrniXF6NqhDuob25O4zwVs19
ljLcKkIBnBLlG6Kmzh9XUgiqZL4LTzcjzrHEnV0ZCN0E8c/ViOe+T22KC+A9+naf
BgxUA121hW9ZBSbSnhUEO6U6uPwMBsmq0p6yStKTBJjcRzT7etpH++h0afoJH0os
KFLhNMsX7hJo6rxjSOu5kNj57QDtGctOJgIrqaQsHkwt8f2J8a6ah42er/lipKMo
K3yVhDYKYju4EWjob8IYG4sCrNvxEI39Drmj/vqVO+0Viu72e6xou81XgBinQAdN
ax2xIDGvt7R6M+9Q8pn+yHm6cykm4+LAa5T4vjtI9W93/C+qe1DRtayhA/E4IfS7
Jy1FVdWl8z4gTNR2GI8F9Y+KEThhdSQS6Tnp8npW5CGIEdKHBjIqKEG1FLasIZhu
lrzyg3MRm2hBndwVMOCBxVzqktfuNJeH1KhyzXx9chhMeI8Y6m03En9KjTXFRVVr
9D/9UVwhjmDRQYo1c3axcIDT9f8mYXUiUrDWkVv/qfnqi4smOdaYdUdtPVVcYE8Z
MNDuiEv/S9dPSlOiIikXVfJnOpECs0jTqbRBW0LnJ1aB3g5VmEmpHim5tjnnv033
ynjKLG18HI4568M/b1o2OjFyb18JE32plf031yCGYMB4DWOZe/ar51TPjxg0qKBI
S/SbC163ZxVBLB7oWU+X2pik2o6b+KN/GIJOk8aFfxaBaV86Dc41to1mBsBGv98q
/OWG3j0galHWWN48btVCjk08oQw5f3n1FWjxgkDaSmxIdEGWsouL01Qygg9eQVMH
xOMfKSMtgzognOteDU1NdJssRFUrlFykc4UFodNxoD4hHFlBK1u2/vnR7lciJRTi
+UpzoZsLao1No4e8Z+YS3g==
`protect END_PROTECTED
