`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M/uiaeEgX77o568K0bMVDx2aFI46fGu5TAXM9C3aQDur03f7FpPh+tdlfTBE45fX
NNliB4P1Ww/eoblRWHyyLrnvixw6fHZV1XiySFDFiD0Rw5Z0T+qA3u3c5wMGJdd3
IosyybJhSHaaOrAQMWMGRNkHjd9XZoTYHogYdAldgnjl/Zw/0APOsX+n/IJWxk38
XBVW6wP2+GKeW2ZxM1h61paFB2TyreAfv+aqBdeAO0OctglS01iziwUuSmvZsps4
/YooMT5bRipGyDtAhwoTA3iXz13sV+MHYOSLMuBxdn+usDFW0Ek9cvCkRxVaqmSZ
+61vAW1IGMLWVCUvOv7iV4gV4LJAMt3lkr0x+OksZYFEUzBbtE5aT4QSOOS015y4
BwThWGVNgZuUB2eGkJDqU6DqaUrqI6YFijVm/5Z8J3gZuLqf/fsqqYCX+ZadCYr5
hp7H09pLpKWDRbw4n/1yAcVv5weG0jB3AdQRS0EfVeBY35nclQuTIwUICOOfWi15
GSMegnz4N93pHZeAtFnoffA/Z367FujhEtI9N06+iWWvCdyTC0aaBPAsVEjpA506
djlbULW2b6/i9dV3QuRISlMHAHZS/0WayO9F6C+IMeIXt2Ooos2f+a9EMlpl9IzU
sl586fsvTV05WtuVYW50SHY8/UfhFE8zdnZp3ybU1GTEc4OJz+KC65iUVyPBtdU6
apYWpfzgyF7Nb2b9DsolzZcFp8FzN9vgJBreYuASRS5klgrG8NhQrp1AoBFdD6MR
JuvEjvGMP0197RjTTzu2R6GpEuJOiiSMO+KD9owtMxiXVm200DYfUCBAo84mG6su
ATFXHrqkuicqdjNmL42UwMPUt8Ww8y9GyOoVg/gL0i0fZcMpI2d8IyYAGYBqht3A
G8Rv5z3CpiuJhJux7BUo8pHs9EEN+wTguG5UQIELYD3rbaNMpJHDQRRqVWGcXjCV
ToIv3L/Yn0kE6NBeHJM1+WQsueik3/tSy9d5mAxIJwS9upiIy900aA+Gxo7tjt1u
HN3o6ConqDG64BhvANoNIb5+zFoaGIc/k4R6PbTvvqgINE0gFtypRUpoF7olB+Ia
u9xR0qvYFP+aN6OZ39xt+M8nzpA9GxMcPT5dNsURKalq7cGdYZNv4ddTksBdvM8j
bSy9gdU73INAhvRjp8ypv44JPuZ4gNAlG2VMN6Em30TT3ZULm+03PGyjDxa/kclQ
vyVY9KpJjKqnsXqK6x0X8jNDUMqOf0V1FM4dSmDx1ZBaErtmCd1NPvwIaRKvctGC
QEqzpTOkv9Ey5Pl+o1UoyH/vH922Ph1imqhvxowalaDa9ohPa9+Ly7wPQGiq8+jj
6s4lTZ0HY/lgGDxc/2TWRRjfTp/p2jQdxcK1wxTogr+zSE31jjpY/R8eTS4Rj3tE
bEVcAff6EnJctVtS29k1f3U9PhVgPKt65QRQuYw0eHY=
`protect END_PROTECTED
