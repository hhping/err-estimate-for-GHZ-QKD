`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5LbQn1mewl63MjAiIll2c4eU0IbamQTxDQSywoo6miXzBJSx9TvRAUxMM8InM+Ym
0ierPcfBmqG6pGfrJan9EW1+LxZ/YxeUJVfNHFZ6qIVP43FacGkBsCXv/MVRowG5
aP+HohD2F/Q1W6hk5ujANlCRfjDSJB1Q+semE4WAZqLNbyxC2uWKB7DWI4jiBo/Y
oA6qDncfT3+P42Quj7fDn4a1M5ZcNbZSSXvBih0gco8Ngh7K59E+bMNJpjzk0IIW
i2bovX8qUVlFzP6pFhICrlEfQxIYcihjoScTKlo25fx/lSjZw4VWRiAwnu/TFQcl
TQ/NCW9jIFxjRKiMZ68e5lSvocn3jxReNlY6+Cjr4qgCEMQBk6giCDLUc9NNpQoY
sJRVWtkX6IUbhQ6BjvZsY62zTud96sH2kIgoS0GttS9HqsxkF7LGeIVEy74DOQ2i
ouYBM2W9a3akmQj4xRPkked61v/oc5HHzhghguwY4oBuwWz/Jxm5BlqrCfOQ15dD
I0oF1xV5QMUTdiJPaWNgPy3W4Rh6181sgJdjGdrxYZ05x24xpcRnFkh0oqrFMQbH
g0veiNxzNBzLZo9yTR/MLstpwhb/qJiQRJcyyzfuLBhlKCIPryJy+kWldxsjQram
05aBBbbN1yS8H0+/YTWl6QUihljmWauP9MD9fymUaApwP5tRCwqnUKyRirdczPLj
NTruPld25yndarDqArCI8xmbd8vROvqVInp3LSkXh8cbMjT1vEDZJZza8ah7HzPy
Wn51aw9PCm2K2x9wMEQ9Z/grDhL5gk1kgOcKs4ouBlxJ2ffnR1oW0WCXE4lJOAgE
GPod3W03p7n5OfP3LyuWs9biLD33qCKw01/Jsyg4ckacryw5FTV9XvyDZV2sJ60y
Up///Fg61gXimFAV2LvEW+pVuDbzF90ITfMDZVZej4q0V/goQdZmFMtD90Ccxy+u
PSOsGjTqyjzq/mOdaEycSRLrSy1L4FXXR0PgsLyOVdKL+UeXibjm8zgPHjVZXzCl
2L4pGgvPZZuKEs2FxLuh5CHFgyHv0pxFLPG258RRnhUVRqvmBxTuqZ4JYmja41I+
mPIyOvYRLr4QkiJDdQMxhXzyxP2i+EUvbmXOQqP9W1xhfnMtW3h0mikxyEYrmvnu
N7V5YlLQN1o32R3zB10bqPdyi2ZFXh+fIvsIgpk7Zr2JMnxXeKbVl42Srm7ipO1a
bzGeJwOEdst+ljttNMeBnudWgiIFC4Hseb8duTFUuNfKVEXvHBjvRUZhEcGsp8O0
ATS++llgOyHzu0E3nA2fof6yCsqwgR18Et898cj5A4n4BVhOaei0khIMEdLmgyxN
ow6OAhx/IAYJp7RpnMvC55nYSxbb8d78xpEYsWlhqb8x6DSpwk4xbg9kUagZsswB
R2eaqVM8CNtA6zJmMXO4spVHfF9cqlmW1y70FW8gHqpglfBG8UdqqbNfoH6H45zl
PLVN4shg17VCpBAK8XR2PuzDK/11gvCVPlRP3UK1PT2g6iRQJk4Atmo2neVriVqr
5UDW7uE8Fr6KiSJXA1Yvk7aU5KlBvIPiG9In9zOlsHyWbDHiviFvJYEB5RpJIqxY
rCzd3yhdZtOH+ZmoL4ZgHFLCtLJCAvsMhfDMs5P9nUWbTVFAa8Q/8leLfPb4u6Hl
MLfKEOwEp0woBExTycwWhAoNIalTgLENEimo2/05g/JJWy6y1dB0cLcKmre3gJdQ
`protect END_PROTECTED
