`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RTDfk+27M7bTJHszAwMfhdnY25xxuDdFOs9x90pR7dQTf+gXpblp45NmMZbG38GZ
+fFL4EUH1dprehwBpzxTx+SMtdHDHym61aP7+3iKRe1NFA09g2GQRjMe+gwhqNuz
Pil4gWo0M35kNRSZuQn2+WChk0S+V4Gr7R4i/G5a/DozKx8fpUUk8in7O/7OCFqj
jn5TIyNwYjZPG+ghPaoIvYpTUxPFhV2Rh2JQifSa7xeHMfRFXf1/xJgCwWWD9SLy
1NBuEUOGvUwQtVBzxGUtTfYhv7f2ZrAVctaqLm5jOJW3ElmHBshoerpp3CDpVok3
Lr2pPSjs3lwqYP4SLsvSTWE64uS6a/AbpzrG9DaDpUgc5G/17JSPqKE5BAWB3QTX
rxniDYZgwRwEzR7OP5sbt/DYzJGAXw7husfChskojbkeQanD3JZm4ibbdi2AUxZp
zwcgUc7/tQlXyS5+dvKeVQI1dlSgNazAKwfcKQknH8zcH+bGYi4vheJMCSqUyCPr
Bc+NBzTmpZUCpafvTGI4kNuwIwLg6Pcy7VwoXOh3volkSjYeCx2POuXnod8Q5xWA
BSRkXQ3jSzTtMinNr5mDDlG7zCwgTOmD4xdDxgPsyuJZzK7pk2zpUo24hdNSLhPx
9aM9/RboAMOMHTkKGJv2GmLbwLD5v2SxLwpztp+NkpTtU7jdDPElW0/T6dqBG8Jl
xHYrnwQOs8vOslkp0e+aEkv16Jisv0ukFGkr8MstYETXu0Tvxtk8D+cFHQar5G3A
hLX0cLozSxFt/XZrE0ymnrvNigBAbMYvb4QjsYZuIo+xRmXqMXXAEphx8XWuvXdJ
3EqDDRRWginBm8A15rpVNYTXhSSUFwLTksXUkHjO6NirvVtDjwGkM5Q7+A1OqDzN
n7vvz51OT7seuBfJCpyXs7rn7qwIuBmJM7UsJOm6uC8g4ume2rdkjAZhiM+bdQaj
`protect END_PROTECTED
