`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T4ZV4wu2Y59mCGgvRKel6Uj5Ed6uGebC2r+PbWWyusyuJvy9BzQ0RSawIDW3tc0s
+1JJjG02Va+Q0cInvppm1MrJwY9eLIUZhOq+bo+LNLDOMqOir3/bC3xlhyCM0BUW
jMTG4PzcP9S31jhoLng0amzSENOn0sHQy1DNhd357FDlOeic8hsDAjrivEha7akU
JQVBVzpTTMAduF03D2zTw9NUSRQjMcis4EDtna1+WG1+M5wgpVkJKnSwdEhgwgq3
Yn88CqLG1MI8tXFCdmLNXNqz2cRxjy3WqxVAQ6TUceixtqsZ0169w+EwkJJjnCKT
1Nye+zzU5fSe6HSKM/Gzh8rbPetcfhaE8kcOPPLin//tIowu7DbUCNklYImd7zsR
u5g+i9MKiCvvHR483hAbEBDQ2tc6Rn8XULRiV3Kr6A6zoVQZHN17+xPQpDQC1Tln
oP49rt21hoUunDswX1fASph78XYg5brqe5dfAX+SFmlecMcXU8q2wnl7yQaMX1sS
JKAUWVbuxEwZxmJMVS/sV6o1RdjcfUeXvILJ6kkJv0uH5BxTRFg5SA6kb4E/Lxvf
u4hyH7RayIojAXFLgBZtP2EVS4HZfw7ektFQYJKAmXkDbtGlJKHHzoO/RruIgflS
y7PR7kNV1sxz+oiTFWPYEVzfLjc36Y/IPxI1oX+204bsDDoxES2IxumQ1HPNluSz
+BX8IPsRb0Pd8/BLLixSIEFNEDdejEBL3W8ruRDIF+FkeFNy3hpPuBxfva/+yTqP
GeCCfKLo8kZ1F2826MpOYD52tZFpx+23VTRZIHpugPDNg1btzADu4Ny/om/U/dr3
KNQaHstIUgg07UL64NEO8EPzBT3tiWrv35e3GYA+TSF/PHCtPLFJ5OH4eYMH6SrK
r+7kdyWf4YSWqkA7qPIv1+BTPI2DFlzQGmdjygVAG+Bm783Dyt2VgAq4dyTdkN8I
VC0Vr+dG7ODr0zkA0Rdf1oA+/9/dtpsaswAOlMNfenXsj2SYySb+myp/tHBtuD0a
baHA5ZhT98BS+s5pqnBo3WEvy++fD5YyVGzW+IoHLMd0mjRuniu5Dh5xtSAwPLbB
LjYQE7xIlqeuP7gskbWOnoIZudPQ2hdRWMHYefI0+xDgWCRKHkEwG2qGT9i+RHBg
SFKyJo5ALI74EmJw1egikUyXytSA3SpPznl8vRLKNk1k9Rjn2ycaH2QGIDgbOCTQ
vk9V+pkl3qfsSa/LEmYKIe780D8d8ABcz2sqSJ7UxiM41beqESJrXVisWZ2CxPlg
vwfJDml6WSXuc5uV1QnmYj/PWLcsLD1zu0TAYcq00ZGNqvqPiJVxYbdkH+EHQkJj
+Ap+nbCm+xAvKTI547r5Ei6Wb2bRS5s9FTLLC2GuFJ0IMv2NNi3vji04YILyoTlb
OqprQkrrtai8l0Xj55VAF1m+ssgTQpf5jhWLEkRnHssExwvVwHqlrX4tZYBoKBM0
TC68HmcJ0JV1rGhyLsWh4b45FwyIaIN4n9Pwj0OvGAKuvs14kxaBsYQFtE1Iwyij
BxscJ3gcqmctB1zejTxDT84YWQJOxHxKkZl8ddYeDKIdIZL77Qg+zX3UiEGuiZ3i
rIw7wd+2eOaJTSGBsdeYAN9AcR5oxAABReUa9TqVQufOG4PbffW5zeIQmKdZAl2H
HsiFAlybrYfchgg0ZAddHz1gd407b/spTvtj5VUoYw6/64NIvlkXm/KJ2o4Afcpl
wYVDYJ7fFPg4RSWygUQvgkAywQNmgofVHDWpT3e5b84VezqKf63X7BkOdNS/MP+T
fOzuHog3QVZfmdPie4JlbBYd0zdF65VeFxwI1rpYO76Pow+/RoUGaqW4441FjBvZ
ZfiZfphGgLteUz3DISMvclSlI/gbR6JHxSaW0BeuG7y+/0v6OqPB93oVVjqQJaUC
filLYLk7Ka1fj73vURuiwkGhetpJqQhyv/116AXBfMyQKO/Fmp60gP6FwBAw7AZk
cN3SIS2O78W4gnkxgTjvLmS6yz9X0kh2BFeGgeBk+t2BzPTgcqo1K1QNg/Mrmkub
0PDXuy8dSt1xgrDFb57lTOdkBjPjJ9UB/z6bwWRWZ9+8YmYcEeLdNIMpUqeXle1I
c/qDqCPSZp13U8P9SfkiqDOhcayfnBKo667gp7UPn9mOWfwGJ854UML4vsdj6/tb
3vdJCp3j2QkToJuM/cEvyr1tS6c4fDkwHv0pSrSvBrHhZi/ZJ1rGegq46JDonsy7
7/82SjXpW/UasEQPxJU2I0wmG6LuJqF9XGRvZPYw31KUZUfxkiuJx6fZqtCMPoVN
wqJ/LkPx7gM1ytNXs8mCX3BL4pqX+o31kO9Gx1nG2ZKmFxwPkhJsrmwQU51SEjfm
vECqZFD8qCbJgIzjoZFryhGIOhDYNrhq8IGZZw3xAiq0OxCv1pOLHGFF+NtuFyHG
oI26VeD7zdng755MoyGLSAUu4dLCFz2rwAN1/juaJli8HWf4bAD5CrN9kFHiMeiS
D9pX+s8mta1AgsAIsAQv8wUz8M8cxFMVMUYm77CpahIP+FrNKgtn7pFHRJgouYcn
kOrx7z3iXqLMgS98HVJolxxoucShaZ1h7csF3krbjjs08/327J3BUKuASfkZHH7x
mH71DiYhvb8vGqtukEuuqTcwIKnf96l4ZaG6NJMPlPoFAKGwbSk7dcOLqUQ37RqN
Uldfc2OEdJ1ridHM1BLlOdol+o5a9Nr+moFLApay7LiZl46LscTFgkd0DoU81ZB6
4ZzKFm7Ih/D+FIKDn/CsG4ZE1FWzgk1ViK6VRIITNSbRbzmEVqlMvdNnkX2GX/WU
v/s2ipkYU3OwkgARrJBb+UTDmmYEQcLDVrPThswAGOsczGQ2tzzA4PLd71eNDFcB
7RCrO2tpMIlXw8A3Lgv27BRP87UDXhNN1Bd4symNmORQ+Z5Gf6xYEJ5N7mV2iDWv
mQf29pyXRjmx/D3pLgkrgqbSiSLu8konokBUjO4W3XDuR2JWm19TXXufOfTthlIX
G9GAd959NQ24dETNYOJyDJmkZ5sV98vSKY6C0QgfQnI=
`protect END_PROTECTED
