`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2PMCgZgTKAru45TddhE4fg4nJzAtIug1Ze1x0iZxSMZc3yC5eM5fqhgvf38OaAzP
a/sKd1jFSfC1whTt8eqRfFY3kwIlnHP9cp/R0h3dJNYymCQ61Aw1f9HSaEc8DWMr
9lAvqjFS7tF2/wT/yFg1Z2ecSVF1Bkkc4vogWfCHMoE0KmnfiZxCaDofAjzSce15
9AsJxMt0Lu0ylecboa3T3EJJKg7R/Wm7GLT/A7sKrOCWvhfG0yVYhO7JijtsBfHy
fkWYx9v5SEEg9cRcHZaPXEVXIUTpW8+juy01p7RccwYE+RuO29k3Pd4z+ClNEVLb
41/mPf0c2fdhWkQHMuAMxMHzM88qMJ1MGtoV6A+g3p3MFgZt375GJTU/qyP3i6q0
9yaGaC3vUyhSIME1RA8Kgfh6kAtCXripvkcdz2zeoq4Z6nknZs9jgfRQbSWTmrlE
Udv7glLRQSX6aWl3oAO9yZPvmxoEnRX+CvDxDox5mOHVokDNofK9emhHsEMGZ+r7
rD1wBDZzBxA/ZVFa11wWCsNsBF9q4ydu+rjscCook9ig3WZrOwqyFIiIZ/JPXZtC
4RkeIzKiVA1e21b8mgMRYvViP1nK7e8Zi3JH3bbYG4pa1XCuO40DsRI4ksUG38Ag
TnALXGOpj7kz9U8exv8Npmd9jIq8WLI8vcaViaCqUZ/dqrrw9Lt4xTw8mdWIOG+r
Hy2a3/lQplvSEThWkAwmI5oDr5fyfH4oVwlqa/C/5BM/LMHzMqdM7+TjMecmgK6K
U+U9YDHU4ZvBamYxUnYEqIQ5dtMZg5cQ4vL6mikLDULLFPEBr1hppMdFSNih7iB2
IMHPkGhWTXiVY0oqFNIk0umzz6JBPIkgKQRqSQbyr0TF5xUvFrL99+hN/7Ye2Mvp
y6rweCd7XqVOVJvn2hrEH4DDfkonm6FYu9A262fmarLaamHOMTNN6HYst59YE6kj
oDH+JjByn1R0I/lbbEmyPDFNkOLNgOKwn7k8CWKV03CTAtBDYy4ERdUJ/Drcu6v6
kX62vWKMV8XM/cPmvNIAojzpQLP4qwoVRcBtHu2sNyQ4rukVyn93vjsVVO8eT1Bq
FO6F+vZH0DkEk0j0Y5kPgHD/M42jBs9piVbdVzXqS4kiWZ6eNW+G7eamVVdJ4QcG
CXPIlnk1156he0U3tHfipQM9roOcdRRJjHNECAM4k3eeatG5aTnkclWZuyeoVwL2
RUJtNIp8IoF7h0IPG9PVrpgLEZY0LYNiA7VGhSm2Ikulzvx0xoRW4ZUqt4qKoki5
1+cyD05TMnECRwIwsWv0+NH3jIqoV39t1RdaiWFeoXE5sVteeOgxytrWCaGEd+lR
9affrhmnxukaiz884LpVXqLfRiKbr9QRTMwOjKN2TUefBZyuE0ZYvIYy7pDJQbDL
hQtoCkiu61XRp2Q/bYLURkqZBaGFxsh9gQ3CpJOYQLK958ke2MJg6M2InwGQW6yH
wQm3bmVEatKrVpHFAo6y+wml6MaaxvwUzqyJQLWAnYSaKyXIzCN8bT+7K2oD/Gn5
aQ163tpl6sCx+JBXV6Jr70xjvlDgV3FI+La0todNu62ytCCvstfkQpLW4tRHLbbW
cCMAW1QQmzw1xQf3qdUuUiAuVfYe/j0MQZaX820Y3hK2VXhausxvJ9QxfQR1hEN1
R3Xc4ekGsHyUBXEJxKsF+DGL21H8IQ8spiR20fBcmdVjsJANUdWR5DKZzxAup3SR
2332exoydiFIpymO+sTuLmVocQ99Zk2fGSD30zJzSURB3OohAXLpPOtvuxgqMMBj
uhCm+dlRsQeTNYfC4+C7DEJcQmzzNME87ScaimubpKCzeH72KCt84zbA5+lulJy8
TZ/3DOmI6EWPWlkj6LnLY1s084jWhRItdGpBzOkzNB5iH/WzXABMI5LW7SsZEmiK
PSYPj7GWOwfT0Y+8lW/hCxUIVCIdnWBYQELdRCwG31OnFIxVKPKtJ63yvVb+fP9b
4eUuHAuViCphoTUPFbTCSvcZa+05LBsGGZebQIAQGZG9tDvOn/1BFUNe9B5v7RGD
7VnWN8CwnTSbABJ87uSmu88Z2EbH0zuViNntbkNVtJ4qk/dNskTtNeA0hxpIxfh8
HGOkQg/r1mbojbutKFXvXXNAbCgDnHSdE+lgEcAavCuHAF1NKwEcdNsN5ZjUFfUn
kMYzibm7ZDE+VxWB/JTEKUkgdubqTWqVVNxasZLSlvbPHqtIAyIZ5xLFcxvnJkSE
1WZMcXGlBoL7Qcv5pzprDtQ7XiSH+QCnnzCWEm6w9x0IRxqGH0cRZRXea+GcR2ps
Nh4I1kM07GXJFfzLvSI3UV93XdKY6n7lhghN1GqjQompYsT6M74gK5YEB94MbA9b
M3eLdjZkyoYcidYwwX1VeYgawJXZw3jup5dmc+ZmGyt9iLNw0K3OV+NOh/MktLdF
NGUTeZ8wjHt6WurA8Exdd2tj//ktL6BDiYk9ViLtT/jo/MVhytyeBhWXGAI9z/Li
WJPp6nbDxHfvHlOQyJdO4r0XN10ercFce50ZKJ8Vjc+Jfz5uEXKfEY0ZdrqTtqvy
4nUDHumoYG2NcaxekNHoDe814fn/qBXZYQ+5jeHn0vucHW49l3GnIYQ5DoQYqR33
ZJFzku4zhoCwpO7fE+ptmYk5diRCmKsOiHHeX8xrCgr1C6dPc4lN7NWGqeYDpcQd
pXpZ64kJVnmMFLNvS5EAy2nP2rRf7qa8QnVLJgq6bW62fTH3HxEvQ8NsSLbmDFSR
UlqAb653n4qmgGeP9mZDk9R9lzPWYaMoBa5V5tlwFgtMNyTR1VNJYp6Eog+EGSEk
tyVc7CyyGRC1cydr+Ay4mfsxORjukORLiRt6SOOneyxAAO4Lf4Fzl94tFQxV6I5S
e72EI2+jpzHADVsvy8eZ9uvPXXd3XNp0V0eooRaA7QvPpi0cCopfy0nZ9OchtJfr
tbd2V+OBr5Rvv2PFdOTuhw==
`protect END_PROTECTED
