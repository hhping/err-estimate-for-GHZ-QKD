`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sINknF97dKNAzupArHRtYHBsYQALydeWGu+cYZqzAJL+8Qt0OUWAyfOjpT4I8hlE
9S7vYH7E0zQKmuPxCBxR77u/uQ4oVUCrJPaP2/LAcoyMeZSDis/9f4Ij9HTVgDfX
Wh+JiUHi/gw99JQtGMAJtjUB8WSiT+q3p925fpCrraOSp7iwUxDRAX9MRMYbQyX4
H0HJMlRXiiWhstpCprHvuHQ9C1JwYPccm01aze3A9Chb5wGXOrLCYD8g4PPd+Hw3
yo8sTNzJWzyI7iIZNRfzhPttLCfvF7YfxG7EiZloZBPo9BNFppR1RdAz5oDaP9pP
8YMookos4JSeW7yz0BLs5OD3P3PcbQdxkbvNA87M2FOs+f7gFjqh55+9ETvSP2qw
L5tter+NqJaPozDcHjPNM0Ajo41di3G5VlbFWrLEn6gKQ8gbGFf5n2Zuj3qTWfvE
FDfiPCRYbTesM/Oeom0wEP8xVSM3nGWaaac9UGgFned6iHKPufTVWpASXx528+XP
n8etGAj3TWNi/DdPkr3LRS6jy+DqfQKRs1j3mDtGpy1tTrHRBwW+1qZpuLDnSMcG
8a8+fll/ZhY0+7+7hN9HhxyR1mwPbc+s81edJlB7gSjf/m+EG/KeY4+onYg6j/pq
LXSCmqZnY7Z3yrxXNRric9+mbLEPJA/kvRZzDTP4Wshgq4KDQLwDISNkJAuDr+UT
2OW+VY0+mNWLfwvhtW3LsqlHaYp9vEXxx9L3w/MunGjLv1mipcSL92lKA4AEhRvh
PtqEgELAR5N3aaw/UQACEdUSlhmrhAoyAZtdgCzJdQSb9AR88SJOREZdCUlRZfIC
NJYYh4znTwukuQLzvpdU+6VfqN0V2U4oL4TzQUaFDRrE8H8rBhBVaI1V8nly3ZN9
EMlZIRo0mWjgk7EJWuCzZ/VrpsFB28iqtHmxaK/2ge5Oip0f1AXZ4QW79Rgxj88B
zXftehJ0hLe82/XBXZBtSIAryRA1igRjJgvRJm+MBnSlfzcrf83J4SENiVgdCYJp
Au6tGuQio+KsxKXSxYsaaO8HEUrMsKLrYacvl+hyTNJhDeqpRAHhaqygnslGGAin
ES0lVUMyeodIciDmrpjznEL5h3CUzhSq12IanBe7lEX2R1Db2LydbE4SLJOoF1fI
eSJRrmCHV8qwfwtqfMmfooJq+KgBAv1JP2XDTK0KTxWnvUx57w26PPPebDvIGcPk
+gdUcbHRzK2KsUC9H9hJuSQ7T2yE/vli2g18ztwsHPdmrANW5EFDr12rFYW8BeBc
WqWRTmtWn73WDPLiDBSXsw==
`protect END_PROTECTED
