`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wXR5RBe7oPq5ljemrRP2afAkZTHVJSyYkDhOLza7pZemKlrO6SyG6Q+bMnN69wK8
tIpd7dSKlvqT1eJMq0oI0/c9rLAFeWGer+l1OzYqSoyJVe3C4Jj51JpJTNgwmYjw
/zrGQkTMunA/FsXl3uMGL5MLAnKaJV+efP+vAMiBwqT75xHC77T6LriOfKzvBSLL
v59l5PNe38a86xOQnizPpoIz9IofXW0lf6hMqAzUamgd40k+RKjxhJc0bZRaiyMN
C/Jy69siOdvF3XNccRxt1U7un+olFNGiGERyQdgcknIdhlUC6NZuyPqUtQop2U+F
kpKA7A1gpOICXe+uBV3KH72lQVAlCTZNb3KssOiKdejagXM/U09SoKG3lh6Qzjuk
THxQcZAe36d31Op2HEiOgioHy4klCzEtpOreOiIuTqOoHaNTwpPKy0/GR/oD9hMX
aeXDX+BxZtMiQEttzrqWJ2/TZqSGByMO1iOuHSoXbXjvvoGLbvjHMFINAvkyn2Hr
XjP6pZ/o70hQ/8S5qFzpfWOBZ+pt/mnAMZZYho2Vd7FHOr3zPt4tkBrY3GynDBsD
XO/ozvIR3x0od9fxm+IuaQ==
`protect END_PROTECTED
