`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M4JEBwQkW496fkgAaiA53UeQSTsb63zs6oLqKMnhV0XEaowx4vajLzFrOgXe0JHi
prSucC82FdJ3IZEKeZewQEf4sbM6fRo4q6gn+Q+RYoIIbX+a2UpuUajwyCdw6oNx
Axk9ptwvliEMsaCqSC6hrg/6K16YsUvWv7gh7I3FJqk9a6eqCu0z5ivnPBVTJx+e
3Iwfgvl2R6F2CzAz2+joFiHWZ4l3LxV0NTak9ki4IAn/4KmAk80g8S2/5LjR0KVb
yBZNEzqJWVJoM02TWPu2b3dAx/vRNhat8DD7POFqAvT+I1+5UotHP51Lcl3KcDVf
0k6bwxpbaCx+lvnRKwJCD2dDeypk2TFZ/ybhby1HKt+E7niryLdxa1L9sxieY6AU
kYhiMKbwld/GwGvPvgqdd3iria8zfgirte/w6+NOvxDqKAb3GJzCQjMoFO2TFc8h
AdzudWbCo6/GYAxf5plWfcprGvGn2p793VefD46MoFRaXXPyTU7MDhyucajaAYm7
NhhYhtHjU8Jo5Ci4FH3xqcHFcw7dEVhns/mG4K/tQ1hBRDIdRR84NU03lPy2KUCh
R0ZumAec5lad2avHP7Bp28q06N9+uqsIH8K8GECh7Jzcz/2XpEqve5N6GFCeDwAW
gHRrbJSZjKXq2CQPDcAy/xNFDlhMnf7pW81OhgDhdtCsmCVBNEGB1EZwbKg9YDu2
`protect END_PROTECTED
