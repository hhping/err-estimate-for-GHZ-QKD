`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sjkwmvGTHULYGYtEd46Mf39Omfg+56mgtFmG0GnMZZ6CsTJky2Hw8Bx53KTQhX13
r0L4g0VPRwPmNxrJbJr3EWGONAuG8BVE5LY7u8OScA51PZpbpbGODWLRIcN+kTyI
Oao+e1gN2jd9dMdyTDEgtcDVgz7T2NJnlfdUVvR5fPBO1XAZEipASB/wtQ70jGur
VK/kExuMQAOLAwPFyl5HrioPGGZVOguQ8YI16shU6RpNTV8EOWg8Ip/3pTcMd3z6
3n7DWXS5PGqxp8g5touFgVmbnIHOJboSbQtuH0hevD4w5N3rHPW67z2Whx0nrPS9
BInaBUvMq11e0hIKNoLhJfteY3W5V7JHL4s7ZLd0HQ/buaqnZuHSpR8eFb9A/UgR
AGsDDDsRbMeFTbKrbDfIiS4MVVhRtzW15N0MSQXMlASZ4DrPP7MFogp9DLhuHVxN
4t+WI9dxbiasn1E86T1wQr9hG5QOUt86j5lAHAXsR71X5ZE5fyxH+P/HYBz2wJ78
9sjKF8wjodrogdkKAodCaUgaCIQ6rxOJmCR23zmUJD7cWNqSCTgjBZdVj7d64Fwv
L89aiEYm/9QYhVrUwrXJ6c8+ykCbmpHG59YAFzyXG592/tKdu6N0mkaaBUsU0fzP
n4qSxn5vTNSovKC/H68i28dj9gpu6Tfm87KoEs3cE5HqZ089vi0Srg9aU9/MQsOb
7PrywiXe/DgJR+6vMQHPRn/VWgDhtfaDtIjVGot90fe00vgOcQ2vFIpUsky+yFCo
NwaLmPQkVyNQE2JNdgUgZ9sTzEOi2d1eMCSaZ/dOqLk=
`protect END_PROTECTED
