`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MuI6McZ6mqsymoEnxXWK2Jcl6/P2DeHSLZCHw+rlcSLnp+pHQg50+vzjjqzzbJgc
N/JJ4yLV3bw8ECDnNL8MhIyAilCnPR/leAV3eL11M2Y1RFo3X+cBTgniAzjk2MnP
rXowrtDrD62ydaT7IrxSUxeGkm3DzY1MhFJN6ws68qv1PuMjYYc+OdHx+A0fSh2L
JdP458T6ENfPYBFDQ22thLk83eoo8MxGZ69bhsncRNqDISb84aC1wu2Q2TJQRYGy
jbWME/u6osErZbNQiYhvglmYYSg+EgAK1rki3jqCVqL0misiOsqy8eG/LB0jK0ol
lWJIXRR0btFwOTS+fyDoCPFtYZyH1+bE8Zx01mvxl1S41d8MbwsIRrTp5ooNCLce
ejiWJbqseoifyYs52+LKf3X6173ELgwbxi0DnF8a//5rltdkgVDmV4ZgBDuxOCuo
aDbVe3IxA4zE3tNyvHhPd+bqn5ZTmRQ6TWg9BLExr5DYPCcMQX8CatSAOsO4AQRH
sFkp+HzJESPvgD7jQwE+ITujCTo1afqnQcoVQFSPXN1goN5k0RTsDMCbH/Fl9ACp
d2Ymf5WxOaEeEm/xgOyFvPosDQnxpECy+XHBhDgbaIk7U+eg83lEX0mVo795enI5
zL2PRxKYowkDSmv2FTuq6xjzKbepla9z9U316PxqMwFdub2vDn0uHyhTAUjBBdOW
tO35c/no1mXGFzqnWKw/LBlimXpiLk/uwWAvQkH0E8LFlbGrvtwXGMBLE5L03Jt7
KGw7D9l6OhVstmDizsVIm+ntyZLa2apo5CPZfMwXqM89MB0xwEePmLFLy/t1HDDY
uI+/ukfT2AMonSsRE/oAsDp2R7Cc0U4uiuKeh5xqn2cUYUYpNN5JG6CEtKcFvFSr
SHIPWgM4ushHzC0MI55Kint15CBONlYLhJbPj1CHXwzPmOMrea6Pg/RZnLqSzZXh
uzyuEnODf/caR1h2yYHtHg5eOuzQjfP/xGVHJCphnvsMBvPhWWibLTIBRLlxU17G
s16InOijfEsVmaDp8/ZBH0jp1WtF66nV2b7+YtjxdVIfLiytag7Y1BnbrzERk8/t
isrHLJIU2Ay1Ltx0xO9L7lfqaACqFgAJHH9LGTpprUidZ/qImKST+9SmpIIHLhyV
J3lq1zuz7av7UG/Kk1j0i0RpIbD7nbHUbw9ypfdY/l3+yRTZ6ep78KKs7RkpGLE7
rmnOxrKs4QOJClGQ//BgTF8omRWs9mpSJWoSwcQhHJ4lw4G/QHecYfM5afKauOK3
CE96qzLqWjNpXACiDrpijF2PwMfu+g3xQnfT72wUHb7sMw3FXun477Pv7EOMluh4
UNNK3jq6/naYUywEMUd5p0nM1hr9AXC5yKZ5nVEAIDkPUrRaWEZbh2GkxHHTh/oi
bIfqsJK4LJnAdYsfWc+WI+WYJpTsTD5U+thicVFSIfZilpvxSBdiFuB8ezoSqUGO
uzmGRPPQkB98qqoZHIKlGSfmCoLNm/3ecWiBnsclYV8pT62gD4QKWtPEKBsYl2ea
1eqvttj7rxexATEV6cCndeRDhKm9UcyEmNov+YkHt2+K/96J5fC8O9/NNqDJhvQk
BVx/uaGA3w3Ujdyof3aixPn4Fn4YJd1sYAEvJPFTo96RBqDCVsJe7RAdWleFeRJc
E+GMO5LRPkLogb1Mnfjy7BkbRHC7CWiR+Wnr/YieOUYMjcGjxO4ch2QDH8viSeni
Vfg0GdSe1qeN1Qg23xxbqEXiI30d6TGSK4gET+351b0+oP+ZGsNRL4TIVvmCsa/t
Di/dcUY3OZqNI3IGJtDkudKtn7rTNC4UqblSptnHw6aCiHCFVvFgF/Io6mogCMXK
6JAU6zAS+/Z5U9C1QSPDdKytl+92/RPA3TPpD6QaJjEZGVNc7vle0aDfnSfdDETf
gmgEJ2Cu9g0AY7ARks+bOdCu6OYbi9CUA2VzP3dIctKTb5XdQQf1ShJd5tm/X/3k
lbBzJV5PkR7L7XVcV6C7KfMiRjvPiMxHF1RymcjoOa9Xuy9/miB8R4SQ5YPrvHnO
2NyDM/uX25FC/DgeKYDls1+ty/1h2swbiipameBLTPJO7rRWj+Gcbipl1byIwRkU
JThPA5ELeFMDzqiCXEvElgARo7BP2WDGbUcdk/UDzzkL38g6XvpcDIwD7gD7JM84
5FS/DMeTVHnGWR2lMO0LKTriCfEogSfDz0p5z5C/ZeELPFBxqA2PD4ezorsAzstl
nEJYWDwNZy4PfKzLRIPpBinJuHVf/1qt0LEI+4vG6SV6NS/yeYoiShgr15mqq4cW
HKH9XgVuay25yS1oc530Cx1vIS0W7m6So21uVRAVWlHTRu7gYl40/DwgiDdOBO3E
ZxqdPF10bSnFlQ8SAbrrB5tL1xZSPeLkWh11Pl542NW25ifhyo8sv6E/0VUh3+AA
Hec1eqpEh6LUNYZvWpBDb0LyBYKDdg0nEN89kFatsSKwxNpOQtZKW0rYwGdlWTvH
RyE2hRAxOl3IECqpSGOR0l1Q6qEO1ONdD/TJF9kKMEfmHfwX2YXBcP8uXEeBBVmi
BdSqbg8udS3EiugFcXtmF78aCrhTNdTY2Q16FOMXLvXGAvdoV2QDMAowrUZ6E9vH
WX/IfHaxUy1NPzmn2OAUPTByU9C1t5FVyykZgpz8RL5K44IrjtWZdHW5X6UQQ8FQ
7h8mkO80EmEZtt9IV1qtcV6AialYy2r4NrLxlHkAY5+sJ5A237OMgguGQBNeUFxE
aNyLga8Nc/2NFW2zuTPCJ4u/Nf8+UYm+YCWzLftD1Iyw4HyRCtO4iwiIAHH2QcdJ
yP27LoWD+cahxcmXHZButEDtNJGLYIwaiVsYWxtrcu2NSmjg6O9oR3FkzKpJr/G6
yL9mtPvqiizbA+mq1QBBvQcQuu11U5cIonmCdXxjR5IzoCx8aWqukwUhuOcknnuO
EWeO8yKAgDJf8JpVxFbAP5JBrT1Kw9V4QR+hLQOcZvv5qY/uFA/XJH7JE/Jkzbyh
SuKCvFAll4ZNPfkMkRqidwtj73QLp9CU3AV/aYVZ7js9rspw6hxCpKZoE4PS9FrK
/E8/HoDucUL5LNAoIFa16dfcNRHkADodmZYOl5fqiH8KRLD2tS0pRIF10/FGZ/A/
C41gkRa1uwCQ8ET+EFvu/2Y8mN/gG6f9ywKdRu8OQAc2HCI4I/rtjCWVR5WRJHuE
0I4Ibq6HfkbH1eFm191Ka9+5yFPCRGOvkj9ubJXycneOT4TZQ54VtoXXKCM187e+
UcBrSLfo6WX6m64WnbskiXyZEQu4IRSvAbwW3QaPcCiOjuKDn0b3T8VXwJJAzBE2
/uvti3ITIyK36I2ID6CM1zf0CZ7CdHLIcGPx4VqILv50Fn/2+ZZHitUp7ChwdKx0
5Rk3J1EGl7Y/pfKzinpKaCbJ7YaxSV/jOD5GA7zCejNooXGWeZpREoPyOJtioQs8
iNSzOG6RIkxc2XsXG5YxNCoo9g4tlMEnEexgbokRyDZs58nWKkLLODnIrjexU2mo
wILN5dGy2WxhwyYXJ49kpT9/7weHod44FWP5XfVgB6HJe0YFTD1ua2pK7WuAuK4Y
4TL/jzwQr/1cFVY5Uj+kUHj7iDDkkqaYGB5KT5/KDt3bG3TP022IA/92BjOpw3ct
h8sXpRghoUOEeXMgCxLEOsssaIwVxqfDPnlj/0oF93vEV5Q2vMfYlNypWrFxP8Qz
1/0sYTb5pNmK32z4HuzUz74d7KcUWX/RVN8/YbjS5uqOcC0pfzrSnawJVBiAZm/p
aGb/cfJzmwQNSS0SELPyCVxjlB10uNf2ws+XxTq1zMAtrI2IM1PJhNGj74fWgM3b
Fep0TwD4WAR6Jc40RqZGSz2o3b2lBiVsI+oyo8VE62dJ0Nca83LBqYqyXXuxCtOH
lV7KuPOkiI20dVF1ytz10/d/0jBFosmzTpBVq+FmDs+hMj557Wowr/SH9nYn35zz
1OHaO5cceKXYmvUeJBYZdGBF6liBNPoMJ756imR6NCC3lLtnsVoQ/M4OZN4qIrLi
uQPUeWsn/gjJYnZwCmqqhkS7wHDsjRY8wNS67tuqjKGVVqNgJgVCWKXBRSUkqybl
Tnh+s45uOgwYzMsOJ7YJhmMBQAHv25cgE4V2H/KEWiDVAQIb5xl97rMxM5Jyjw0L
DZfWzbl62/CHRMqH2HR4pWlzdjaNwHoz59HTOm9lqh/F8uWloK5xZHvwEz5Rb1WW
O/tqDzRTf8Lqw0txptnNTb6PV315qPGClkdBbc6NIbz5KpK/GLNAj80iiVYL9tSS
YqYvCTc98hrUXk492GMUf6staAYO3kFXkPiyGSFTYQs59tSgz26ICMUmBAMgR70k
FkWGEzhkjPwPPIhVnKMvor3u62nnNkxUYFTLnK1y3ZPtcdD/NodVwWH2WoypfReq
0vq/FERofR/b1teotJy2lg4fKAemh4lJ5S4E4kzpnWeq89v+n3b3BtY6hcR1EJ0a
NnyO9c13mFaQPzdMwwFls/44151TurmiCcz1GCdcNAUiLKLxfrRl4n4og+FNKAOf
n5TsFFRBuogg7uGV9P4mWPXh4620BgxWYaWSrOxfkGVGJzRhUFaOCYVfdV2966KR
GqdpZoecUbiqQ5/BS9a19KV89SB8jlPa3McJDIDGOt/0YKvSAUBGUfz9xTlsvAdJ
/Mhr7+3l+qHaNJ9Vssd3xUnbVlBVcSsx9Mrc1/bZ4nplSRB55Gd3M9FGX0paFcaF
0NtKMoDBTbqMgX/U3lDd5tDet+36Ldy6+26BQnitEW3N7IfxbMb1XZ5Ra6Vo9WMR
pqdE2M+CWhYFznrDqgU0UCtrI1zGnFmtkYIf7rlWyCiain+/dQ8TlcAMLvlq5tKZ
mbzdR8QubLXJzv06WR7niWqkDvZWsNUzThb1dc0ZIrmUbKjgKagnHvm046vPRp+D
sKKEjqnWhu/CDgyBggd7HXQpHx2TuNx7HKl3QeTliPBwQVB3O2c+JSjY5wGF4/nM
MvbZTF84cI3fhsi8s86t4kExaacHwfJAPHczXq8GK5ZlU8gMgcCorod2XKewl9NK
OKiRG58FibGbMsNGfqniETdXU6veFi9SL/zapPZGkPqgds/JQTXtD4FowllI9ECO
fysx3u/6UBlIlKcF77AzkvWCn/tD1F7ea71WpL6e+Xk4ONJTBxemGQhLY0hIUXtS
Q6ORUWa764rnPbvxlJU+Z+/rEZJDwn4p+MsG/4lusJHjuCQXrufATfJIx/q2iSRz
fiRaeaggb2Mj9KLKOg+a1LkUxqLqqWFaPtgTPfHTVWEwPj08znHLaFQ4p3y9lHrc
jsER9aEpY/gCAP3KF+84TAfzF7uFcZyldS35BqdRFxQJNqdqATlg+BAetiuG8y2F
quUa8TJg17WUGEXBqzzR84yhp8xoEotM03vKuc84FpeJYVmC7YAHiNOkap2i4jId
14d7c8eq+o5y6YdPEj6x2vlbZNF3E0Upo/QLGxtXBNKZykTqGBsJL5/+kbghcdkA
fYV2Pxy9J5pqEvUs7vDUaHh5sjVBuhMKhoZPM6xhQT8kJmb9qjdBVhDBpkU2dInv
bm29Hw2YAGFSwEFya5/4ay48waSeNpYwT3J8O0EE49bM86EUhdVCwHri1yqDgSE/
zD20cqwKtvh7Or6GTdqoxdJ3intMsDQ2MO7uV16SH3+ZF/9/RtrmF/P+jju5R56c
sZBiyTEOKEqT+/DjFq4AejKNQaDzv6X9nnmruxzt4lNlWEuCMLuFzCFWuBgbc0yA
h3dWSkAofTt/yrWwn1EI7Zi0vQdNxdzhldqQYHiZgPdCBZlSDrVM7QvRzRPglUrR
Me6ej21S1Zjdk1mk4gRjalmOFr0bJOjUbKy7zLo8k+WZfptw4s0NBR2XVTJcvwI5
x4iStfd2DWu9fNh0ibanLnf0h9Xe+xvn/VIAnVLK/cYLcpJDTW3OCoLWpsm4cL2F
2YOI9ChNJhBqhvnWlyuw1Z8p0z87uOlHRALyD1xHFBeB5m/PJYddSjYzUhu1EoPr
XKBSBRNM/5l2lxbf5IowkVb1Owx6+Rz/a4OKzaFgVSe+FIEO79fUVUGalrwX0/Rj
hgyc7bo03MnnJqVdbXFxhXUO1iiZBPSaAeDjeYCOD5ID7KTDq0F+1PiuuDeiZtb9
utLYN6NykCTvhAbV7RflbyMBxvzKYWmnS0V2jsPZXuKH7A8+zqrq39YlPKT4gIaX
QbcjPOCBeUgHlyoBVN7fAUgudC30+N4SVBoPsa36DoD8tlZtkkOO5TFTqqtWSHID
3PXnQFBadvTQXspWk8Ft7/0NnBAtSH2ersy5F+yLGHenePoC588rpGA81yBqdlR7
zKW4b9YPYe6CYRFLBka/H3FVrcsIKqSGxFqQGH/C/lvHs4OlCraNBP7rfWYWbnCu
0ehyXmlK5gVsxGBk84drKA3NBi+IrKsGdYpeaqNBAHF2LDNV7t73f2OQA4nQ+P5F
EEkOQ7kOq0lMG4v0gI0LcPSWnIGJKHWAaJUglQY9D5DgjCdmjhj53v5Qo6VllybB
2dSpBmMagcmpeJRzjPdLTBKMvXRlFLPuYKPALAwZQ98xiClDkNaZXM2y218dS59X
5PLezWmZG6syaLZvQHYyi57YLQ7Fmv7XZcYQNDNz+LX4TTsIMUcUuYdK4e/z326Z
VeJm7eM0mSduf/VqNHV5SqLTtYOsb3z8GdYKnrp9HG0CjZfa/dx0+eQX3DEiw+CS
vDVElSlBmctdnXVYHIXD0bL/wGbALbmFOTkinG8fDJNDOysW1ubT8vT2uYwqGBxU
I8Fb8qBqi2gg/BqJQViUt/GpaKvkHKbqCzDywU/xR9trSUuWq9N1igFdZzNIQYpj
CLWVtrU356N5szfdPh3r+6juPfzy40CkrRydlq9JC4tGn176hMsEFVviQbmFvT5T
PON36CFYwpxDnWlm2vfo+HeZ0pULrl8G156OH6yZlxYlCL7x9m/zjmRZA+hzZ/Ix
mbbMw02uJ0E+kuBjwh8UPHYHJzMoXLeObCu3LkUFZ7muB89Fmr6rpjw0eDeEoS41
cSnPzfGO/X6p8d2c/BMN8H6Vy6D2DxJO8u3uda8vFehNqnZE5nA5hPrXt54sRKeU
X96Q8ZSf6Z4B9iN/XIYpbGuBEFDLY8ZJIwPHDiLVurppOy0Lf5L8Xa1dhvwCs8kq
5NFYbtKEM8IaL9GkQJ0qNyFhkUmfZnfqDMVab/UHWepSw5eNJojm01ZpqBeogcGr
qXdiuMIhcm97JObiQGt1W1aYMbCVyxyV7HGrUhCi1EH/Z++kVAwbeY8NqJjZGzaH
aWySknTO6buQVto3z6Oer1M18GWG3eY3XlGxVWXHplhIoEKTbkqQW1bCjxbi0Gjk
VEupaqxackBcTuulc3zAg7ioiFKzkP68ZLBFmv6LWaHK4bGj9paA2djxN13TCNKT
uxcXbbdxi8wu5o7o0/rc3rTyUbQ0IefXTLIYsSHsqq+DwXO1HA0FjZ3k6tYVJl+m
F79Vi/y6rt8HB5iUH0ZMUm+BEOhnCvRE3mGHfxIwJM7/Fg1a7Jv1S5fYB+P43JNv
b861/8Ly3Ev6R5SQ1he4JimEXmIq9DXhXcs0VvCIE+wAupaysL7B3rRp4euAFMJf
fiJzkkL2s5gTqpfVq2CSGEhvX+SPnFQUGY/1xZg5Fp2vPRHjaZ8oucIN1FL/jdy+
X6QRI5hiolKZxVAI8vX6ysYB5DcBxF7GcwqBIEESqjrPa61RGSYuUMe/mALz8wPH
dd2mQt8aRknqD+usrOrQBX1NXIpNXU/8paxRthslq1r5gjVsbX4DRj1COfne17kG
r2sQ/pcmaQkKiBb4ak64Ot8Iw59FJFHfwyrk/ctM8DAlZ2Qd5sUafXgRrYdrnU8V
q4ilJJnm7Lfl/hvoxjrvx08Vk/7d3zUHkRxg5QKmsRSOfRoLf4Mkjj8Mt/noQcT/
MQZLokSkjRLCJvZuD64mnbo2rSioYgK5nfkrCBbCoMcVVOEB5N8Nw3dfdwUkCzh4
Z/OhiXKxnSQjlcjHcT1b9eSp2fOsx90nlPehVdlOXhJ7QMHSj0ijsYX8P9/5J7YA
ixOg8KiIMLSFxpuYYj/LFqm2rXy7GPmZUXARwi912sxeQ3VuHtDL1qTfw24Oz4c6
x0e8e0g+imPpm6Bu5DUgqjcGwYrAC5RESqRow+ToEAipDGNWXmdEACXQIQ/bFC2G
hZzpysstYzddKsbbLrISJLaWgFghhDsJzsx1TyelVJ8DGrkaXSLpwvXRWP2RV1rk
l3ibvVxUbYGo3eMoXCLKEXYedTiQoNYRZwcB0yUVaxF0CZXVIcNwSxMXxWobFIQ4
iDHodYziPNEsxCftn/rPyem6v5T8LcVX1M73ZPVuXwPLkujkWGTP0znwipi00SZZ
YanNYF6kVkXt8z15H+Ur7GreD+K7ODZip0mhcE8zo8Cb4PGJdGqpW6GImbKwg5xn
RdfjRuFo4suItCNGBqKZAKKM9zqvkeP0gq7rswe563rEIoB7tO3NP+kf/L8IJ/o3
f1wHNs71hNhP7SHzqeAIhTFR40TitpH6GDaaJc6D6eXGH3mQn93c04hMyw5xOuBw
gpG1fGI80Fm7omDeZoilliQjJvSH6yff51fw10PGLTzQXZSkTiEbleI9mO/kvFLy
MefihTxqp0dOhiqMxwbh1BIWKWGuUBfhEKbCBvE1RZE+xFqs0Vj2ukvMIuB+zosx
DjxcLSaDpit0D+xA9RgafikY1RiubDfHN7gWZGYYkDKgVBhQwHldU+r8nRHw13fw
n+vqtcevpoDbPuyX504XnSYHQt5D5YBHkCWfwfWSV9pxswN5YY6xluDXoDUQy0tT
emwCB9jabL1hrSshznhs3JgZBqqbEdL9VTLRsYYDSOLNRQmuTudM3GBWamPOzt3d
/JsBDyvqicEXmDU6dAFZYw==
`protect END_PROTECTED
