`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QJK7SNz/P/fa+uEoxSHnT0ByAgAHcl2mLbLmCXI+JkoIEg+X2s6F4FtHI8Ih7eiU
BaG6c3SvbfFc7tk5L3GgiOBmR9UoMh5zzHqOoDtq1cUGTiTQgapLKpYIwbJgU7lZ
hMl/vKeGi+6TY/gD55xyZ7dxoGllau5fSCvo5vGIuQ9PiamlTNRkdmmvG91vcMq7
PquFDMiWndy5P5+MOEX3Y4XuHei5oV5AV9jyWrB8io8bBWWsFXlYk239zMoS+HjL
yn1BNWKb2ANGU0eS/fqkehVFWndX37F5b5KLlWMzv2wrwCnm/OLH/5KK2bRqkpmT
4hd/+lpXMPc2/WGVk3YCNTJ/gmGzrnZNM12sIKzXkPWEz0LVlc7yJpBJxZFAnFO8
U+mYxwZesJ6uGQ4XeW9O3nkqsXVchi72ZzbmwnXp/tS3GQ16Jg1mB/eN8Ksa8Gcs
X9yhZdPIT1tz/SW+d5mp3z0eorxIteQAJfDLrIdkScI8YNZEVbdbH+6tfa8l3+Zj
c7fQmx/1BpXjbMAm+1gfyykarUocnqUlFd33ax82RTNnQbPrRr3Uaoz6ZXJE1fZf
ZaJnBVnj4awD/pSJ7MvAjQ==
`protect END_PROTECTED
