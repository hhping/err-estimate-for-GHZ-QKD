`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jxt4m+9x9zAaqZcjHwU6YLXWU/GPzAIq+gUxoxhMrPKl7P2hAlYhFKg8tBIm9tqc
6AaRgDV1w5K2QPK8LbcIgpnE+ppHDfvD1W7/16GBg1TrBitFM5+3rt2MWMSSkLfm
cZgRbZesbKKy3j3VZIaeRFEE0ViaNltF4nbslkf+KhRucBDNIh7MHd/INvKziU2d
ud4vjRomjsIISNqjvvpoczx7ujjTcTSag9t/ObC4dsMQkpXRI52hy+wzlnrjkBYI
/IcPzByVPHZSPVWL11V3DqIx5xhht0Zb0Tq8TuRfneLtx+bdg0bkqS2/RcKFjIP7
`protect END_PROTECTED
