`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zqpmO8ALKE3iC4IMcOg3dvgnpYYpMY+HNhG/6NEwZal5Qp6m0qtWAGXAThWa4J+Z
r/N9lrBZEg6V9aifhUEu7p3MQvvjiopYWMyJa7Be+RMlbSx4aFMhrK+pIS8xvcrs
KSgyrvjlqsedzZurSmH0J1JLeeAFcEPef7bItQo5e+esJK31Fu4KQDpakKLuXrwE
xye2f81bQ6jWpXJ8SWEEVq2WsG6nu6t7IP8ec2hiZ3SB+07N1Tcid5mdDa8HuIWx
TNh3Dd2ycpGuxSzaVOAKWWRjfi8EbzlLTTdNHelUYEM3kQEt1I2IROW/036gm9nS
uNlxZ+hGgbQm7chpBbxQbwQ1n2GQJem+wVuj1FAC0tf8pFDAFNljX+Z4RrT64E2f
Z3HGyMGswalAmvJc7Zq/bQ==
`protect END_PROTECTED
