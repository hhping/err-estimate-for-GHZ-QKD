`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PunNDzwUMgRvrWV51vd9nlaaj+G4iiTQB+yexk/PWDCQS61Cle35aeKBYNyt9TVw
wwiKEtDqgtR3UKUVZpxmKeWi0ewChN1cxND75RwF6DN+ncMzUzWcNinav26WtZEE
4ChDFYDJXtsLzBlskalqhTftVE6tnXbTSUfA+Nais6hXXtXkuH1/lA/DOO0/ZKyC
za7J40JziVuCUlR92MHfkLacirVpIUfBGYI/JJAjEDdVgW1FcwjGZepNBf5byklJ
kXR//PfxCp0EUaNIrWlUmg0HN/aV4yChjwui0TZq884i0TO6RP6rlP0Epxf7SiOu
Q+OjeyzsgtDV5Uf33UyarIWfQsub40w9vek2x74q04Rj/tMUr3aLaI5Iuioy1EPy
wGbw7MihZWy7+mJHzxSR+JSystiQsR7yQqFTe4PlmKhPsbFF0GumjOidWiiMRzHf
g/AbsQ0YSFjfsbS5+X4F7ZZDaAUI587z53ypr2R8X3TxAaFrVxGd98bOml3habx5
lpl64wmbGLrv7XcXnm+ut3chPrKWys8Leq5pM7f4AbqB6m/fmiu3ZuvZRl9dq28J
aob7OqQ1BmqGmUnijeXwcEh3x/WVjvrHUE/UGYgizHqRJCnTPHZ9yz4ye3mUva4d
Cl/0w/yw78N5LKqdvGeW8Z7cbaFU+WIeqtp8295W0gWkqVWOY+8q1ngpvYzATbNp
Mbz77JgEODLiFlzIkcOBg1Bi+iB8SPkPpg6PEf+900dB57YINKzhwb3OmU2etkrz
BX4pBKmIJTHfmeCRsxK5LclgcGUG6Jp4jM29WMu5+h9A9ZpUUTb9TbNdsbue3ZCE
`protect END_PROTECTED
