`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4wVXKkZbK4rZ70h3dbJ7g2ezLNoGRBUUnWLFxeKKbk7Y2r90prKQurUXVA+fK0+H
HoZJn2hB+yR4W6bdnVyHWatsXYQ+xsfsbe0zskrLWYTfRYG98Xxr3GRRsqHSihoN
pis1zU+odLuE120AqJmC+pUDVdD5ZgUfKNAfySw2MXjMajhrZO5XVaHakKmuwwUw
IOTCJ5LRdK/+WjrjTel/NhAeibjE+5ZZaVGwmoZdTjsIzhPwtHMJi8n5Eme0PLbW
EDL1ZGdHavcA2yxIxWBDvO48+c8HFgt+1c+vGJ1fE0wRULfbj2QWPCKDcVRqScSW
t/41H6RBboDGvKTp49fwljRXInjkUzlSQvN41DW6klRV6cruUUcbUzdvZ3UbTO87
6TlkJW3xFs8U5trSWwovnqwwD+2WlUGmS+ZW9bed+7bOpOPvqqz6bDPfNPaI8ot2
HJNDtC/XOx2HpL+hj9mXzj2EXpuCWlwhDu+GSJfHCFwzl5rqaGalEI4EvL5hsmGb
XKKmgqwVKr31IxbNdfY6GNmTgVAMP/1fx/i+DMp2a3ayznVH+iYSul9ue3gxxh56
JYp9oV2Ft3sAbWcfcyGLnRKYNQ0DZNR/dmBr29A9QDT11ehFanyNiId70pLn/xCQ
oJ6uMpog7WNM4bURHLs0gQx+hKAOMPDYQSINiFfGqc/Mbwzvjy6sdNsA/tkw4i9h
aASxvj6cRxgWHePvPybyyAydSSIP9kS/LuW88oSMCRcLhl1jtW5GpLiNXb25s/MZ
mMj+h2gZ2LM8GTAq9TQ+qowyeYmkxIrvP+zInvsbzk6PB5z+ChyojgQz5zJDIQ83
1xBkXucPz1qhUPIfQubOxQPh7CyeVNf4AgLoESs2Q+GozZZxVjuKzwWC1PKNkRef
E4csw4Qwu8lQafM1BROw2mELST2D1RjQZVZp9htsctGhP75h4I6jDU/PXc5Gsqyn
q7ynjXtLAPi8AtMclHyweAwnAN8dlBYKt6ZNiVc9XcdlulHX5fryzYa7AT2YFQ+P
NFut6rHd9fj+9nBxqAZcERNon//N2MN/MrTXit0g2qKmfofWJuCBBji0TQD5nhTP
cpkwImPXZ+ACgH7v4IA7xQql2qFS2RZvxt26H4LlpdhtX0Z2kDz7t/qP6YW57r4l
F+EwQ+uuP6zpYfT9DJdgG34/G6JSZ45M36ZH+ifrW80NRPWOEh47eaKrmp+46rxS
i6iclsgf86SbzUtqvsNZX++Z/rPVa0kUQd9rmm868D/uS160noFUl9thaoP4MAl+
CBxurTUBQniRjskAvbdUzu9dwImw9hFG4mgAeq7mSTeUgD7ztJvZkOkSBiOvXwtq
mmM0Gt89axdf8qXPVuXIx9TiUHYEqDoQpMhTQk6gxwnvdpasRT5CDUFYAilZkrUn
7nUda0oyvN3224sJ21ZuylDEwcsK93mtmZ9HhrpnR3ZkNGtAEg54anDyvEVLlIWh
8sEHpR65QpWUVqGzNZrFGD/QI0MzPUslER+xzQMQMoyF3xq/UIIz02PNNkR+dZ64
piaRgEJHMjRjzAyThdYddw8MduDDKnqgnx1u6Dwxmh88oe/qpZ4aSouvxhy9+zt/
neImBQPQLP3wXDaETEn6TuT9o8zE1oPqRczXB709NAjgdV083aOShoGBUvhB0FPR
Pnxs+2IYesidcUGZ3QD+7WDPfSiasCpep8ESgzjE8qvXJOdWPiO0kKYfunojyDxe
mE/wqM0GiimxzU8drCsqEnZ2VJ6k1D2DeLu5kuUEfwpiUIRuLSaRTma4Bbs+B82v
7ZvdyYiSLEm7gH5CuLarn6TBQD7gYUEdENi05U0iw7Sujfs77UNOqaKahvb3CczH
y8DmXu8CQqdJjv74DGTSSvPWEbKmPBOzjc28rWf3JFeaisAWJNQTZ8wb01QrJ4Qz
+D3cBHOAGhQX8UGfRRfT13s8UBZqSbq89CwB/ukS6cJr4veIsIS1sV3rTPxpjb88
YkhOuct6LevvA/X6nt0lU4p6LuNLAIdR6KcoIqT8g3W18tajT6OU5eDwlrNQHhzQ
kde6jw734CiXvWR6X9dto8r+AqmMTm+LjBIz8oMuUABYQEhTE5dW1xuJR63/vta9
1RF2A+Vto41MTJyT/nhGFi7fni+tT6euyM90veYSt8SW4RMLYRiN8GKPq6gIH2aZ
8v5QDuVM0irnR9Y9f4IK2MYwnN6NcJ53RN+zQakJvvtKsN4bb1UHyRsu1Qzw7qhn
5KA8Plbiy28hBbKZlSAgRdbg1kz0EjEj1TQuruzioRclwwmmx9xB9lDHgBtLp1dJ
aRb29uy/kV7bJIMCYhKPSjQqCaSxkV/SPaX5X+juAbpASVK8zk7tX4aA18jaf0yT
7Q0lTDKH471HP0E8nhovWWAYcxE7GC1wyA1kDjzTyhULaDXYzajD1euMWPy5BMah
XtIqz7fHvyqegXAZxR5uXE561cfjOhw7vritZhsWzmmnB+eBiWlM/7nOxBDGnGO/
XjJ1NTnHWeu1G9bW1itgCEtBl9fscVI3LQPS6cf5uLuqoui6onRRjEhvwFSD2Qu0
7BllzU7fiquCsqFASyencCEPcVDyNlwgrOKoK1+zOSC35JaH57ptaN5RX+2b0nNF
U8asE9Shkkz/TCyavn6Klc2qpB25XkYonHxqW6oD6DcMT61TTS5Ng5fbj/CjY9BY
sC+b4c+urTTkbWjhtMgvSIGKPAZC1M5r+H14knfOAI4NCHOjJqn0KXQiwZtB8qBk
SH0E37G7ah4FHnXCpo3Aw3z808s8bvNmvWsd8eLrgtRZeMmBHtgGZZQtpGOPm3+s
ZPhoW/h8PYnW/GO0QQTaeYmtBH2v057aiM9CfTWF+bLJij7We3UJS/dOSQvhoWFd
ItdvlUDwNKL5t6zN+g9WI6GPDqc+oTyB7fzN4SL0iQS0h/n2sYRFwlyoXIVAQa/G
d2oae2U75+1touuw+p+iKhcE9iVoW0nUFsanjgNMEltOdxmRfVF9OV2wwuvLSghu
mw586bX71QyzUcVx3yS1HxFlJ81nJZqJFiz5StIEHJ4nSzhh2Yi5QbUyvPyMrE0u
YDE29v3zNSWEN3esWYcpUgg99mBvsT7T/J/TzSuGTKVIkwLTqmUeL6u5KqFdy67p
y65Zf2SqA9iQ3SvpnqnE1NtCuRRWWQNC6jBlDxeF1ncxq804z6c6/hnaJBJ8GS6a
Vmq7PBdhjzhL1U/traliA9XfbuWf0lDAulAMIHgnsKTsCroosSJIKxYcCcx9j9N2
gr4D4jvDk3jXi8Evwic08yBfUeRHUXP9C3yZKkWWWdmY03MlgXyvRlGy6DXWRKkO
1zaU3znKOYGf1EWoRDMb2pRG94o7CLos5uT4fjfHvNZcJH7BZu5X4sBnCGbQ680W
w04kqOIbLAHNvNbsuscSmQEYgsS+s7Mamx/TTLwhxbkQLLSH/V89gHM+IUz6nfmd
eC6MErsCgvCHf6enu6djR0ZPiErMUnjhszkHraqgThTT14ia29CbVZUME3Ezf0zF
zt+lrR9afMR1zc7mjw4ZyUY7Id4n7bcQ1jKpP0QvUsh2aP0qLhceDOvTV7bgNviV
lM6h/XVY7A/rFS+g5Jtmfe+xE8d+QoNmI2is3Wj4JzGftauH8StZWBgS9Clj2ai2
rbiC6KoFvtOJ5uJu26lgX2a8432IHMrTPBPUluxfKtb3wI++HekgkprkyLy10B27
tae9GMEAUHpN+BgOJAqCb0ZE4Mcm+pmg9c2yDY8ryxBHcIhEvC2o8e0yickzT+Ph
Tqz7pt/0UBKlHsDeJEzDU2TM9hboI9OhHtrJlBq5NrVgNqmys364V9GNkfZqXZHj
i+xZaun4bNVNSQhMA6pFdEMBNXKwnw/+qE2TBlgRie+fHQrMilFF0Uh4857Y1XKF
0P/TKJo4tw4D/1aKAQ+V2sC8ek9WfmDoLP/5VT3uEmyO4fkcsCg71L55Yyli7Bvc
uhaibz4H5YelOru/zPRp3GjOpUjn7ba+1ZF9y3DKysxfT7kGS7oFonEAv3TImU4n
Va4coCnvH8ZT0EnzudRQcZGqix2ZVUAcL/34AHbUqaVcVHamtfQOq2QLNFIP0SYW
BW5y3hgMqCFNjKPpVVT3ymr+1ig2OHFyVzBqRQ76nD6b2Oe+3yQwjeOhxpVJpLYN
FSfwPEW7DEwcRfhjAgxZQcLeaQf+fjBn8rvssfsazU0vR4Sbi00Fg5YHOR1i75h/
ShYl6paUOzCfNkt9l2idtNIRIGUpL6O7ISnj36a8PsXJ6ZW2OOb4PWmddixXw6hO
pzEz+z+0nDZm52CM6mHWkohgtPovexZ9BNyzRpYSDr1nPAUUIFZTqrBqDNJ9RyOM
Yb3EpS3gI5Y6FILPojqDoft9lIQE4Ae3V/7y+wj8RfxQFRnuYgXE4/kKfqOeye3N
lExHX3CNVJ3p+PE/UXmS3m/ptsXnvyTfa3Q1Lyq3XwKMej6sVxX8jsD3IHIHBvUW
jH6zaIQ1cBUYdqGlPdcjU/mQYwtRCVUx3FXM7LLEzZdoL3D7ANeORhVSIWqgz+YP
KZVsig5EeIWn5dwMUqYNB5riV4SbHE4dfeGwuNjtR32DgDdHt2C2ArGBztV7WUlK
18uQMAuz8YgmUeT8A8FLDmvZ0AUpRXIf8Wa0lgJkrXbnig3D8GT2YT7cdayJCFfC
mrxfGiXxDsYveRuXiUppl+jIUgMtBpen8R/DAjn/aV6N5tEDQEOSX3MFavVajrmi
dge+jPV81eBw5dqVx2cxCOPmqQPA87JJT3PDzPe4fPM5lrCHRVi2exH0fHMY7RG1
PHGdTObKYytXM4R/UhL6S+7DLEHvr9k6Oxwq+xxF+vGPmU97t4Vx6GlJZ3+WwUE8
8Gpd09JYZgnO86vTTxYzZEGKHNNF36mChR8G3rCwB39tNfDH23ZYTjYpX+6zGinQ
8PNjE7wZjW1f0J++yzsgdPx4zzx+TmWKqyMhIA/XmAa/nuI5zOzMydLxaknk5xrP
Q9boYANqigVk5JYRfP2kW/6enHORqYzEYvHwTJAgp/uITfI+PvHsxiqbif/95ZQO
lTibhZsqtW5P1xzr0osclOrJ9cYYPIyoyCeswTZmcFH0hRv2PJEPkeC/w7TcY3mE
GFY5/PFBNyPUCebcVVDQW8QbvLVVFSH/3rU3eIyS2ADchV59e483kkA0MdUnetL3
CHVWIStSyczyXmajrMgM6RtaB543d/rrvOHbn45hXlDEbZxzKz7T4XJUi+G+QnP0
dMDup+KDwcjm+3HGy63vZ/KmG7R7ymemGnaR6GAneU8iIgknf/SuOEfIs45JT552
UL+5a3umMBf6JKox/eTG5jln7rLzNGmJyGXivQGP2n2JRORfoM7WHH2ll54qffdc
z2n4Fc+dLvWL/YroFHp6Z9tO25523aMvIId3dUWd8Pl6WkDy0s2zdnRNDbXBwDeB
Bkt+RxhEYTi4Y300YOXewW+YqE5e1/gcPTQunvkOS/JCHoSzydSszStNR4KpQcFy
GN+2w+sUsNy3TyRsh82eg/CuOkrVuoibVXWd+7sr8Y692Js9zHfxR2jsgELgp47z
7uAPxLQyzkAXfk8yds3GMMnGlzgfkL/lfX9vNkqSmhtVvAfepE+MFh2nTxtgeGZj
v79iT4mTmTpL4S5np2mtbOqhvACqiasQVeCiXoxcw8hxwUAzrKpxhvvoRfRFZeTs
SyO7fNf64V4BtHwaY5LiP54qAAcJfsQg5/xIx5qWlsCD4DsBSeh5lYN0zrUrIpWA
JDp1PBA0ZKt24ayyqkTFmkdynju2LjZvd4llzrCTwSjX4VhwqabxBzmizVLL6Jvy
9UWlw2WOLCfHa9QVj53ICsx7ZGWxuAVqQ4MxjKGtID20uNVzqVMjFgHJl1RDiGCh
sYUXBW7eytvWzBOjCwI2KkS2JM46dosivEKELq3oDOAuAERxzL9UQWubyck4nQdh
igJsRoGXAow6NS+mNrYW86MDMn7aHdVQp0Xzr650jrAcLdyplHoyHkmIshjV/uRD
b6OpjA+0gLY4zqmzbtTn97dDVaPCOBVShve3dytSGBh1bMGUcwMHsj2HChKaFTcG
k3EbvwfQ5M2DItcw66ZRuUX46GOvnQBfrIxg7AM0r3tvqyKp7C5GOpGVEepCCYJ8
9A8N77RofFZjyY97HLp4TDOh74Urp1BkKr1LfW+Uv+165ird5iCHX0l14uVlW0uJ
oojlZ5qofle3heoVS95DNrJ7XyHVJ1gEZ4X88ELfjnmrfd8MIMKqRBT4XOIzlLu9
LtgOOmRHHRnJMp43M3snM8yWrUM3SAUQcKi8OwhBmyAt0A8Gh6K91xHzXRWo31+q
UeMrlEAtycwaKQOPmS42QpMo+ilqVh7WeOtWkNyjnKtHzH2cuqj+HfooI16o4IHs
zg0uBmXox7Dil3FpbXzY4PtlRGu8yTQHtxkrX/w7yW2bmHrqBCkIzjJPyd/cQhga
gD8oQbW+qEGavJjWisLv1+IhRgfk7h7DCEJXN70H6QR2NmgWAlmAHIGI6cwxLsZB
P2/QbOvP3kZtRZMVJ30Cm16PX5OYDFuyKp7bGTvyg1uWcF82ym7TuQsFYc2XbIcu
yfDk6Tn8h1SFksP5OJxlqyjV1HwYWqh/S3/nroVh+Lp1t05nA4gpspbbhSUTreC8
Kh4FuNMslLC39lepZF/EW3MF60hGMIBrPooRgI4cd9F6mxK6EvKdfs1inj7Tg8GF
lkRWVPe1tauS/1BQNvDMy3NNPmi0Y3iFcja0FpulvRAbjsFatsk9e02ynyziGh2r
UGSEZLqlpRB/8doww/Z90y1jQSzpce6rW/cblKQYLSXEMiqt2RvjkGat3V319dS0
0OwnIpZFyIvS9fm1G/igYXclpXxTS20DJgrhGI2YWzEv0un0eIU2RlXORTLbqf8v
KJoUXTuyfAl3tLw0keW/6w639mji5xKTboCVJNy82W5QFYXfLv+muPU1ps3KFnSf
Gvvpid0+H2nmAZagOM2206i0xjjI4xpRTBtJ6B3kAKzDlsBB0FgpR3neO1ag+n/J
we2Amn9SDTq5lqtwReXhsFmdz04+tflTTtHSgVhXi0z+/kQ1soWC0NgSPXkone7x
AbXdHy1mxSd8GtygPQWhF0C8G15CT4cUwZXZ885VI+Q7WgHDLCXT9/JLZ1FYcZBr
j0FuOTxqcTjxTHt4VBg/l35/sDS2gkN1tmnDmhltm0og6G8ufzL+r+Z5madzSOPo
AdKq72pwTQNHNSdpAWfqnsXSMqqszwPEciuogWpMw6edQRh1pjKqY98e9OBOu0ty
dRDm9jWeTueaw0KY62D+II+P66BuM8H/T/uUMNl1A08+L3h+6kVZIOfPnLrLE0Ok
85oq88Sonyc82eLJZXj+DebUwXcfHfmpAf9fkCP8NxjvvBo7xoBYNphQOf+UJQjj
zsvGvjov4DYJaPaR6P5HEev0Q3GqI9Wl0yeUEty9++7y9ZsnDczfGOgZ7bWm3aEw
74OCLpre29kSnB2rBWymcCTiKtC24ZOsHypWINYQuuFT/+1Y8nBe35jkffXdvbeZ
rrJT/DBrvwWOwzXie1MLdiop7kalFf+/ug7FFMIYISN+8Ym/lhwHFeRaN+Mbgbzz
ljDzU4Aucvf2jG/Vh0KhKodp2QcGocSD07DsAB/OUpE+A7HvSpM46f0gOLVtn+/M
chHIojhiewQ+dsfcyHN9smxk2eDjq1BtwYcw4m1MtKiWCdgKT5grmYlxNvvC0C2w
FYFDE2xSAnPHPqTaFFJt4coCs/T0nMSRkQDJWFd4Mt1C/6gGBasTccjBm4sy7Mm1
HoyuRS4cR8b9iY4meQNmuSzWnYEsOuigLNIKC9YDYhDbO4HyDPPJ0+HXg5H8fQZu
IlzBOg66std6wkFgFZGjSSx4g4t604PByd/19gZ/CSMqURQ03xh074TaiItze0JT
i3pqT0mPUc2T6mlm5+Y4xfbnfd5ggtS70lr+ixt8je7ugSjkUTs4iv0xzOk5/R0u
NYaWiI+uoBWGY3ayZ4ncBhI1VG3Je+flndq28AfYW1Ksc92q5lAIWO8AuicX2xMy
huq24p8Y+03I/AOalntL1GKBWpYq2rWkEwLBXu2EaUV4btQZz9VmE5DFNVEj6tKu
QSp7mEaKgTZUDAgC3TaIlfeymxJ3bXFuch+JqsmhVb6g8i9lIX0YauhQ+m8bD/TD
TjufI3Xrj1cbr7Q71j0koKQ2adMo4YxwPjAL/EbsSgJ6pa03ltFFTa+ESEdAd0aV
pW8i2eK+Fm9+iqr3hZZhutfPRAdQzyso678WnnCbU/67WqhrfCwfukzGZ8mMB5UZ
jneJZ8lAGcZWZya4csZfF5EnGtevJsDpa0UF56XU7YkP8FgAUrcLQcjpeMGMdqDK
KrWUgLw4EMkHkdEySYCMSZoi0DzLguHBSDgFpfsFAFNhs+EuEuQqJjrM4Qxne0DE
agcwnNLWZWidsnbXwE0RjpswpseoeiVa3jYOrQr8+Vzg8od8zGrWq0MSbiCPx4UX
fx9zZb0GjTDD9GIsIjnrbooLf7hIGccxDlWrARc3PPgLBPVg9eYB4nzU6inma+wm
BZ9pt4iMC5+KbbKW7UbJwAoxxqS8mRgUjPUNdLZ0EBubCMfphUCuCD9yiSgkVIXy
kryfYFnjRIXnHNzyJyIgO/QGy6lneXTE5IDjsqH4XxVDOJg4ok88l95Tck8IzUfm
c5/fs3JyeSGf+QY9c9L9PzClQks0J/eJLnrjYS4lkXbFPRYbgXkMrK5/Y1M4TkGT
ZUCsROgCM3OWrqr/j5uO1mo2V7XCNgbDndb/JE+encpKgCg7X8pvuB2UTjQv1CZm
qCRaNCPxfXR3IoMIqYVHoqD1y1ZeYfnVSyfkiZl5IrUZrhVcZyP0Ly7bfP9VsncH
UL6l9i5Sn4CmUddVKyNHhq+7d/LTj3gzK4mxOxyMDEOJNwLAV4mgeGUll6u1f9U9
tiPrMt3GaJ1MyOB9YIdI/+nzC2YgCC00urhLjnUYqofEtyhsHv7DgJjwBZpT5msW
allZIwY9xmXrfTesTWX8tQ==
`protect END_PROTECTED
