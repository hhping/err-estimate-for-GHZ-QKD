`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
al9Pr4inTeI1hhM3PwiatCLf/YbvlB/XzW69MrArI33iqAc1ZPFpU2Rc4BvFkc0E
m9WRKFZ17bztwcYKJqVrobTRhStz1WGmqSUKXJS31qXVNwZ9NCRod05cnrdG41oh
pPiaxfd4E3SjzWUTQ5CYuhNEHy+8Qh00bBeehP1pZc3lgFki6GsqKdNIcwi93WE5
pxfkRjXmCIsgoG2jCHZjb4yfqZr6yhRe2G869v5jvrwq1VLK7y2fZqgo3UFEhUU9
yMS8YsJjnECNjmVtv29931dXEiVKadh7WM7YtxIS4+GY3D+Yyc+yFXpXqItpJ1DL
8NtutH7X78cDZL8MROg4voCBPnUGON0q3rImAOUG50lS+gxa4x776p8lvbgnlWSR
Swik72fcdto6ugNo50CEZ9SkZhRGWFk9ZBUHucGh3HtjFAxXI9MvSbg842/odkv5
r2wjFqPiEnWUdMDqFBSokYJV4b9eCnr6CVgmfG1ZQaMoxIlvgH0HZyrroVbt6AT5
F06ZZk66CxK6guB3uYNlAVSTjEUF+3CjK9iRcfZjwPtzcsgXfl5V6a0CzeRG7KwL
RFcuj8yOUEbxLouKydGCZKlFtGqoswndHFy7IMAdXdBGhUUfX3PCDudTEUWrjOXF
14tFiGAVvnYUb5Xmf2b2S4ABCkUiqOrUz09yrqLRkIlwNM+0G3KQk7LpUeqCNy1A
nPm5/P0vCcACb3ah1mZ7sUWptjlLVfUOJrrBSmFfqXZg+75lVgnzgvoBDvN7HybB
`protect END_PROTECTED
