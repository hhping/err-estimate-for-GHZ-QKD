`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wWN4fr6apWzKMPd3k5vjnYiom/cciKu9vL/7xOpPwdwwvjbsFXAZqOD+wmGoGLjY
BXE1ZwjV595INbmiOgvpAlNDI6c+MDkHHt812FHdSEMKp6JmX1Pub+kZAeXe2m7G
3YcvSThMfxxhv86fk226weXFKb1eqDsBxBnVcBlePFNPYVbaTcACcLlHQle1BZFM
HGleLVZxtAxKEVoxT4mRgeZNPvKEZfN9JYEQY+tj2G41eo0Rz3eSYWqouGc3dC4h
HcTPYCzk1fZKYol758SfzD4K/dussRxeNLpPdjtyBXJeWg8wRy2k4ErI9ifHiqsa
jut4E8geEp1KeEoXvgObtNtkKKeM1rllGd2WlB7k2rZOMwjCc0yVrr2oz4WXG68p
tckUz++AhjKcsOZ+GIrYz0ogc8Ua8wga4XZWmPoilrrUUyI4PE7Y91na0ctTWz8e
H2ldtMLyueCOP2i+9aN2/Fig+5xX3HLRBOI5b4HF9p76lJLNic5vDpMpQeBTBEIj
nuFCAbZndxhqEDYvV4DADgwT3uPoPQ7oSgbkinBmcTQ=
`protect END_PROTECTED
