`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vVXjJlplS80t+l6v4UXzgOOtQC1ekuAv+Emsliy6ZTbF4uUyMFNFYYK9Nma9LXK8
CJQyAZbZBk3NyL6TB+1spSXxaGKZryol3pPT9EtQR4Er0pWMS3qM+u6cw32A4tne
fgSPca2XJ24rxxbpBxkcgjDQOZD8PIrdkEoY87kqjWh/p/BL7LSqsf0Sr/a0nCeE
0xR43RhFKMYYT7h16/TU8SGhnFGvIdNFDGxQeq3OujtUI8KtDAKkxBZ5IlgRxKkb
TyzaB0GsDn5CfeoXC1KYXDDiNYnVNqCPTid3hzCA0vP3mGFAuYDQxXSjIAZgn94y
hQ3EMMuTnsSilVRNK4KZAC9TaXaJztkoFYnz95PrlOkrXedOPhy8WAjQU4LiApMp
XbQlfv4XGRIabJTyNrzaC3pWB8nLEM0fWmrS0qZs97sa1vQMqRzkH840KmBkUS1D
rvZfqObNmryfS9gEG+nET8avu+1sbUA/itmU3vdBCk55kvbzs2DNoQyUEZ8uDw7C
dDQRXLmG7NO3RAE52n8USsg/zzc1T0Qb579p/WfvLRJNYlJJqzH5T5HvGzWRwZkV
JFvsJUsfkYq3zcyg7tXzCjmXUfDK+s8GNSE5LDQci8thsR4+Sm7lP3tS0WVEBqmo
SpEA5+uvbDrtc9V/jxOLAuXtgv1pAOadkKPkv76wq3au+kquiVLbyCHtwgK9Q35b
f+/EvaKu6LpZA9d1Rn8SqXAQ5V2PbeUbkTOgPvZ81YWu21yU818ilLdrItQbIj/Y
+QrmTNtOSSD9aFvIghoxm62IYvX0yN8eLtYYaa2eqxckdA+E1a6WgeHAsSJSXKVd
3LgnsxyOu/lStYOQL3LSsr2AUlrjLPHZ7Eya76kBmzOyTtNfJ0gkNooOg5LyDz2K
erNrAnSdGm1jQfO16YmLv2MuM2/LgVIbhBxjBN2tnE8ClXvh/zSq5Z1sJA5ipgiB
X9lRpYT6RpHys+Hvodbzv3dK2tMvCVjufgOU4lHxj9p1SKTICBcFm+t6nVw0246l
lsX9+AJ8TRIh9PML3adbkYuq39blyHo3TI6JlVIB0jYWaBAshuH/VW+DACGU+t9y
vzI0eupoXhPq8EgZr0j0k4Z8whnXX5kKOPCVv/9pFN9chsU+Fo+L2IWGVqdHJfj4
9++/yZFITUqGYXHHUWQxEFPuUbp2ot9TonVyF6GMoJxsx5HsUYQ2EQnhdQN4cM4D
dSiWXK9OZuZhkoTWp5IbBBrYTtezdAi1cAt3pBGZFWrQyBBkFZim4kCCN3UOYuNp
bxg/4zcoNcFF+e2A+v3pmcUSr4C2cDJ8udf8fnGuyAs=
`protect END_PROTECTED
