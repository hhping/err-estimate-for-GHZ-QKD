`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mKLWaUK7j/jgwl03tWauePYfFcHzGuundZH+DehZNzdwMwt1/sVZzXscYUje3OWv
kRrjwx7/Df62/M0Y3FowBT4tOXtsKbXWbj5hnLYg4ApXJ5yzYyRuZ0SKxFldvIub
FMfKo58tGK3ggSGX48nIi8Ty8G0OVGX1DFCwL5OSrk2AOcP5OWPCOweO/vYTJX71
7i/vT+gMYVPZlUJ3aWIhhZKkAdNvmbHCzsre6CEDSyoO7E892IxqBVUxvE5lDGtZ
nJgM5YBTaQOdM2/vOh8USboiyQ0NvCO+w1NKySGriwc6ZsJySHFFZbSnJhlM44hN
+Y3OvKMiyl4VJvRvNj3Wn2b73/VTVPLQFx5E6NBiSF6D57x9k5X4js6p71MHwCNx
mUS/rqLnx7G5NvOva/eKheyT+R70AA0i9f13O0Hj2EgfLUXRaQTXTF+2CAntUPne
toTqiYal3SC6nS4oaRUm8+hqzgef6PbsS1o+ZQFwIL0oR+0U5pc+Ndu9WEKXnSxP
KgCL1uSipTZI2WVfES/rWJFbwsj+gqpB3khY4j3HBtYnvOxe15Q+AXVdZboeG4E/
0Fw5yiJoSfJXPIJLcz4cDKAQJGm8OsD4IY/Ny+NR2ShaVYzX+TUiQjLNzZpBpBB2
zyY1/hckmNWhUzXb3WvjDieFxSAUQ7i+bEE8uTRZZXXWnp+IE2OnPopqY4lMpnW4
TLbkOK3iq8vR+i2yJLaEdmqqIyT3cjKuhJq1p1BPZwDpAvx0TSTp+9Y5KSVZkJfY
+2q30aniFkCBCP4gQjeIg6040qsjiYjPIgNkLym4Fl3+b1r4A20oJmKXsGs78LK6
D/ccyUj8GUygwN2onecMgfCByuZVHjNwrH+neMMFCQhvIoSUtv5HSDa/axgnYI+d
XQxV1xoo65DhcpavWH0YxdrYi25DB7Vwc8JT+XYuCjWZBjx3zMq/kCOEYjbN2SDR
y5lNNoeDEX2jChsuxSKTXPUDqqGoQjK38R4uyWOQkpuzR3aP5Qy5xxbo0f3HnnZH
xQcb68Mv9eHNBEzf3hxxFNEvEXht5teENjEGj4c45ETCQisCg3meK7NHlZXNIKNa
FNlNHzeFYQBoD/d5rIpmUVPgNNvEC/hkhs9Pm44eNePKthDaQfWGgHzx4MIGOsWj
+5eBh2C3rI5TAbDdwLVS7ipQvwFMI/48jGWzEaDd2HJGylqa7wkrRQmmIdtXB4Px
3rg2/GjK5rPBUMtpH1QcIqhkbevq3gCwYrPeekb2psmJSOhkYqcXhYr1uwtv01aO
N0GMu6xiW0yrARKli59kIY15LLeJgozupPsAMyk2sw7hFRFzkYsk/I+oCXUpaLkn
LXT/A6D6qd2rfvhsXH24CjVMzu9MlLb14nkq8AbceZPMMzOZJfS6EtH/TVsuIOrh
rVDAdU9iLZJ5tJL+mjclJLBgIdiWBKM9OmnVzrXUaii+incF7BF0URqZO3+Z1FLn
ptJ7eH2hVuiHE4Rm65ElmFiTyxNlJGmTOavidR2WwrIQthiSCx9GxlAKp+KbCe9w
N8riFBzEewfKAn1289lz3jpFuWLB1k7ny//fijGvxWcUdsY1Tt4Cnwz4NdtgufLF
49nnep5AycIEX42jWGFoGI4IL6lDAbQks9npZmlY7RE1Tdb9gPeFptZ7AxopUe7c
2fPmBcmspFWebcyYoE3P8TrUFb+5wf5cClhvGytNtS4S2nU4saWU1ybVavPNPfWw
S+zhowJ/REldzqfwY54lyY3aSaSVuXq0gdAW8j2DkmNe8NOVq4HEqwdG8nV6pR4E
gv7osRT99Gko4nYUyp7dyHHmbAhqF/iwMgVvYJqIt3n1/m2LSlCbjogatR1yZ/rs
kof0aJ7xoqrbf2MdSJMe2DmS0VvOJ6QkLQXMNqHVI0TmmYIcYDnIx1iT8CrSH1e2
YNcMpqCvN/gNoNcr0lC4spq6H/CjLZ/5s0F45ODq3FL2/MRJSWapVI1xOf/ekI4X
k0l2PDgw63N3nkQNG8agLkdalHLnbAtos/2AQIk19tqLVz9S+lFrxK9L0nJuh0sy
CQKao7YgKR4M1pXQQ5V/0p4QJyvtCdNpT/JpKMNVYEFEOwC/bxVrSUf5Hl/ZaM34
9OqnIr8C+kgTZJnbpd5tHjU6eEjh75hCe8qvY/6W0AljEau9TM3iMDkTcaqJ0Il7
a4qLowyffiWH3o6bHmOZCZIvWtRp5MFpTtfuoHRW9DQP3sxyt7aNmxYtGcNRFIVJ
R4kWLhJC37s58QYrj85esegK+TrNBH6XuZharD4bpP4TcVd1gntZAH0GfCutYxDl
r9hNTGYFHTIkz4QQE2jVgto05fn+sb0aQAdHmZ+DlHh+DR3A48IbjGKkvnIJV/6f
IATxHd/r/KjUTHcVg7qybao5w/Ntsn8ia1xkWVV4Y8w6JrvFDJYzszJ+uU2fZdBt
ujUXALn1SuyQ0sOXW5Pj9g3dcDwilB1uGgGhVw7cKRwKWXKPUJnnjt7DCEJCAIHl
eB4OSvv9xPIRbw/26FVPTuAS+sNgZBn6f2fnO2LJIN7zeA91w+m4CoqX6baL8Fys
mwVy9QjtOmwNYNurhUDvPozPp06VueAaBuUR5XPbAsN8OcwqflES6TMk72AzrUL3
ABdEQSF9agcTEIEDdwfKWqgeKRa8m4CC7cYam4NXQHWweyXqT2TyGIdpWA6Q6cqB
A0IuMeysjLU4rHbzOFvaurZhaF+LABKXyzAVijnKkBruHKkd6NtrvGwXPQiCwyhT
iWKGUwAtzJugYYiGqSdc/SkZQETGW+1QsPw4oVoVqFaIGmbhliNG9UU1DHlgI7AJ
605mV/Fvs2TRX1BOsPxPBizMrg8enI+m9Q4zG/72gZhDEONv8hi0wxGXBEndvNLV
nQV8v+Ombfq169CfKGtq/dyxXv05M7IFLeocODmVXLf96lZsu3lMSS+2n2SH+jg4
Q355RmCtfi0bEtwaPm3cvM9b5w6g83uOr1mjXOKd4KWq9bS3/Pne31GzLzwcX/Yk
R54iZEeWiN4nhCqhXqmUm2xTwsuv6VTlhDgRtcN4yiVvtSkZPlGseWPVCWf1LOmD
GqONzEez4mJ5gh6fiki7T5R2U5KQ1cObbvx+rsf6TrAZhqMhi9Kji33iPnExoNnD
uAhHWpZQRpPOc8k690IBWh5ai/dSAdR+qZTqSxcIUOYwNsOCgeKqG8LX+XCs56R/
TvVnwB5vFjmWE8LDChHV0G3XsyuDxbCrBwbbDmyN+gMHnll+RMZd4gvMKBM8tKBY
rODDqg7dA8+WMUzOb88KpS3Q9gmpYsevfjiWdSZODPlrNzrnJbzdujj4biTVilEJ
/4Kjc0wK6yu7MBRAnGum1umCcDIU5uWHglwAbi7qHgRnwsGaLGb0o6pjSAcMCaSU
stD2JMDYig7tibd4DxD9uNViYCY4zg3euV1/Rsq/5LKa+boyOAlN34TnpIUR9/S7
U3e51lT7Vuc8FM1SGN37Kuvz87K/il2r0OV9znaTsfyAHqe8+uTuNE7jwI6LTSqE
APfldHsg14K0Tzp3RSBTv5WK/l5a9toCxS0Eor+b8H/aq2Bkw2G+cSLM2RgnT3V2
rYXPEPPb90gVAgjvcDDS2m0gAzH2r3OO1xLI6PXEts9VU6yyJnCcryrq3S24ZhYZ
GndogzLU30CJONwtlblILqnyd8fJPXAUxiEtdWTGXPYMmc4JTn/2UvylHVwjx1Q6
IAlM6LXH01K1nPW4LoVtgc46AMCKciOsh6FXMwUuefMyaDGzJ6Flw+0DR5xf83cX
JIt4fSyx+09MGa3X/584YsXV/ZLb+a+4paT+KFRA8NK+raNW5GzFpLcHryi5t4iI
a69sTsOzjT/T2oaENkPm8LBUQa9ti93X2KmWYCt/6X8xs+rKPKCMns5+QrEdPKnV
6h8FPMFq8HmsEi87P19juar1cpquoR8/4nQTn0CgMMf/VIoPOMux80+tzMSa11Zb
FZt6GFrUPbqf+0hXDjCZ20Xq4sXadN03liQaHTRflytwyLRE4oqOZDcKkFuex1rb
TDQ0DjQh2ub5tJII+d17Yzy0tZFFMTw6Aar7O99L2STvUpfh+jdn9Fon1zd3cngh
K9TA+qUVIY9mNUJT8yMYmskn6Kf4gslr7ENXiMSppyB2gt1gr4jBQz4/vizNuoJw
pNeJMd1eYijxp3StCmpLMs4mL/GXNF7MIr7E+3OfPVxAqxLzKyo5Aj5P7P2gY9y/
u7cgXTZV2WpjxnCaLGjW3tHZBqxgYSah7WSbKUkYzkg7RJf3C5jg8qrQsyqtHvbL
MB7mY5ogGlSLJDziDJPu5NZ8+ESeYgkiWiKYcqanV/5VyYcBcmP7w5jNle+H5JrY
IxLuLqCYAVZK2ahCzaqbUvvsx4oCY27aUAqkb6KbClOWfn5ddqriGK3HHj3cXHNI
l6bWgDCaABX21VPBI+G1NWs1GDMvCus1PJPXTWce3G+ogK1zochG3keAqOUtH03y
b7p/iHDI6NNVLJ4W6btYqWA4TvOqK0G5tY0+rL1H+gk=
`protect END_PROTECTED
