`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YmZMTnSpRxcMbzq/xrJ6pNqz3MLEHYCp6K3vP4SNsrtTZ9ipPso6UtdNyw8pib4P
MEiYlM3s6sXAM1tuboIWgz8BbucLZLW4lBa4o7yXl5R23x9AmJRCUZo/g52SBQ9c
vn9KByNecvCRwGXA1IvjdnRG7rwHUKO/dsID2tTyFSu7NQ2q0LpOpWfaC8EjNsl8
/moUEMil7eamgKR+V/80ndZ1v3OqjSYvFog/kNP3jQ3XJYoAhpoC48wJx9PUvybL
i/wTBQFavrKaORCQxu4mvW3ToyLLGd55+fbkD+CvAbFp98GLLjmDpPgufzPrZ0za
EQdBIAxO50XnzdA8fjspVOfm+akQB6/bqNpyyqcwotetycm3ZW6ObD6nD/4f2d02
/yygkEnn3BWn2/EeVSZ4nSqqyJhcDj4hd+ylIotpjhCzhDGy5Zh/26gkS/rr1eUK
cSp55uVttgByvOo0GrkebzMC8WWhow7NjcWnBz8eEqNVVephqjWBQF9r3Jbpe8+S
NpFDbrQKfmylDMUDcecrFMD/35ICj0jil1z5uoTnjDgOLaXB2IgOFMNjk7XA4x+q
X7aa0jxDT6fD4c7y9UBd1eF+wXK/MOpz28v+MxfWiAJrVBKarETplB4Qq4kH2PRP
Ze0wRuSMVHeb7wZUyvgHjACJLo/YsT1RU1OTGtse0dg8HozWD0ScE82HrYy61ZDS
pTfKczAkLeM2qeUr/a7v+ev40iakK4UuZ9fOimDobQIcAQjO1+p8FTdA4pqJfXes
AZ0fBlxePpFInquZAY7iGcHSWtOX0FPRgeJMXvkCnJ75ALXsoYedsTtqqw0GIUg2
YCoD9T6kk82uAKZhUwT8LK+PhwGmum065deoBrDpfM0Y5735RVXvu1HZe3Fs6fue
HzTB56+Bbkocv2+R0/viCqvvl2Ecx3H40W+H+ZBjve+pTh7XEUeTNiUD8EOgPLor
kqSipON/rNc+IIqH4cFoWX4CF6uoaCG3WGe7CJxqVE3WFa6CaekgnZCGg4dRNrJO
iRQqmOB/btiULeGC9kAeDoLqfziqwCvuQdUNwOrdZGdNa4/IO/g16OeAyYf6SzxM
1QYOcqQTxAbNd10sBnt+z9vjouaIb7f62Tqzne9kMk0xZaxe0Vcl59H2Q+DfOU/u
B9vynwRZ0zqyXrSzgcxCleVWR2E5VVDWN0yz7437o0HtfOwMnown89J8ta0p/eB4
F/Rzp6Lqsd3qXnqogcbPtEossDOnX8kUzyOc6hRMHyU/hR0zAaKuCG6Ims5pKUAt
GyIDvcYtnUZxEJRMTdrRvpun8SbBbxf/sWrwykS3wflsvMqm/6IVxGgQ6tgTD+QU
jboR1im6Gh3tJ3oepSSnxeDXntrvQQSHNmCeRQDYdx4vrGggTyiGVN2Ljqo+h6SA
s3nHD4p7d35uKb7TYR91bulN+9qvMjmaPncMOgG5OLaZdkWNa9oCMIv/GREqtAUL
oVOIwwYTDqQm3KRNidRM7Oo0gHtn2e9ADBVMEOBUXzmOUj1xPGYLrrkNWXR3MZgh
aA9ToPPs9euzM8qQKDS1/bYkHcjsilC6czhSjPqsoSnyHbC+u5TmNk/LzT10PP8i
j/Yr+dmkAcr4TPqPDr5OmyC1dfn6LBe+yV4y/3wHYETyN7mkQ6qiS7DaWSTs308H
coSskjFFmFh+COJjzbXEotUYbTOfkRJOqfS5AB28DsCcxNV8EVT7PzkpOjWvXIpb
o5Al3YoWV+pWRiJSfRSn1m5x8+cO0mto6AMFHjSitVEmhDEKZ8DRvYkMVyah0CMM
WM/tI+kfyn0Jmcy3OTW1y8BMaq6scJxgGz3zLNEsq0Nj0PmYHGCIJ3OYxmzNenyt
6CAaIeg+svnboFMx1vtSqb9OvaFMeJb78IbHmRdzbZevqLde+dyGVapc4h9xdrZS
2oa1VVLB57NPDGkldMqM+xI2WJwIo7JU0j119M2JOoLRnQpUESTCQfRLN8vAAptC
NXbp/u0aDd+WZA81xhxQXVzguBxIJEycwxGCmj8yGAOb4kjIwWldl+rMxktKElEA
CC/3t2Cia1/dzpDyaNxNxEy7G3acvsLhQI6Zrk2cb6JXxqagPgn5rPhlY/CnyRD1
st3q9ny/BV94J+Zt29bQITvCT2aHLV8W7VT91O1e1ogKoXr7/yLCw8xHxvwnmHc/
9uMjh4uVzCH/pyQsAA7DPD1Ym1Qr6zHkSEtNFb8N8qjFfDj3deWEn3JgHtjTFBKB
C0f/zT0twcpe1okfu/c6YwMcURBXtgC10yQjuDSDQBYnl+aT00nWJA7cZTTCk8aR
Kn1Og4jbkVje+Ck0/KP047vc3V8Il/vE4tIghzU3S7isJUAwFBgbQBh3xnFcmAdX
k4uQbZ6OEDOT/Ee/Z1Vt5PCGagzxAqHMcHv0c9rXbVNwYtvEplm3CTxB3og0QuV5
dYOXc/8Oq89nj0Hf1CGiyE1Oeo00JX6UI62W8WVLnnWpMgc5AVb3gg7Nms29dNda
DRBC0H2rdJ31I0PtZcp/R5Zl0UcyGTp3qh7BuyiKopr8qjRJveQWoIIJ76P4rLeQ
pLeCqCtzDBWEpQCVLdBPdTqrp3hQReu+W/mUfmnQbdG4oR66xN5b6/G40eDAngAk
G+1sb0hrXYlNiW7t/XAlINcvVSxrsOBvkQJeMl9RdbyMBP27qxJ1YiHA37xBdflo
4zUpiQOQzniww0UgKwuJHrw6GZ59wPR25xUunQlkhq3Ae6paOqRoaSirlcc8d+MJ
7FdyxZnFspZW5QnOfD8yVRRHxA85VPmRFUROr4dczOiMnYr2JDnhhJ5NYhn+P9S2
eOo44S569VGRFBFPh1+Frn+K2vVIRiCrQRGt3Dij+qoUPqrSlgGUv/GEZAwK1LsJ
2OesrkyFf06HcepJvZbKo0aP6TEilgTkWNYDPvQIqJMvzvmNia33JyvoP6gZIRi/
KOo/0o4Fxf1lyCwXMc7YObLjiH4GNt3ECeCYWpEOoQDs82UvYrtqcji8NIua34+k
wDvAw55myCkW9jxmE/Z5ovMMkmwjH8U3N86Z4jgeAPoLBXCSB/3G5fSWUa2LhTfr
unF/AWLMwWaFYpYNOM7Ck306e6h0ClF1vGk502kk5G6a37zBhfIZnLYemkx2VmsG
d6GPq/G/ZT41pNYc0kQ/Ebs72cSJjVrRswKe8rppTkxgBV25vK40sq2xcmEkiUXS
2ipztkg7wksU6n/DP2lcjL5prvQHQZ793FyFLe6M//med4+eiGI3zbhdwcYJDSRB
71NnLV7rfZ1LJDHZTXPkdUIfcUPwCp9dGhylPJTiOfAE1NUhOwhFliNPmys9SoUG
5qVEc+AOnPbalwtcGUHunR5MVwqNIMm7R8DgvmCf4oB+7yA5WYhOOHEKKEK4O8Tp
zL1tA65zER1pHxpfIi3cs9vRQJ2VlF3gpXTEWelA+mO7A8RsON0cRa6yZzhKSClA
ddDLR6LfqysRA1mWQcOMgwGDLRcCaXN2VqRLAhR2rHk7S+CVu15Y6+fPS9u3SbRN
ILXAhW3Lw+ub9Xxktppuhx+nohdffDILFvMqTFMcSt+gbSIe4MpupdQ9jhL5CV18
zv11TMkJOMfEQDQNBcJQT5vcyzGPnUPLteJ6TBVLx13oEmzM7n/Yfh/HbOC39qxf
ZsJin8Iy/4ByiUulKTeEbyiyopbHpNyura3SgM3YB3lJMb1k8B38HIEqpRVewQ+O
cq1zxEurdz/UN1GZjZrDnGdQoUQWdvTKXUCXOY7JoFA+LRC7XO5iaC6nNenPTj+c
Hye45XZPDOs49vwtooERERGsDRKfGyZxxnQGdj+34LL2X1LztXTQVVUrnLb39Zm9
PHzAhePaVk/MhfSR4uT3R1B9wcbKLJc1oDRoWKSk25DD60wH4w6+msdMUsiNs/MT
tr1xB+YZg/+99JDl/d2U9MIcodR6mV418PzlH8jiGkRYnk1VJitybZLpa2CRb2Mr
IEkzVfyrF+1efvEWZVJqOZ1wdp5cP3BUax9FfcLP15WhTfxyqUda6D7a5qavIzl1
7s38VwG3+ZVGg2bZvz/blB8lUxLU4+WAymg6/WKQ2jy8WFy0hDoHpedBeg+WzdDz
+nTsewKY31roh6QaGGaRScyG8DsLOEqC4BcWUQrNIpCL22zGo/8K4cEYQnu9sQik
ou9rsfDuwXBpNURIRmbqTHI4ZtSFOfSrUHeHhO4ISqlgW4u+Bx8Lb1aDWl242eFf
dpTW9Ns23NYMO3LP2UfuwaeMQJapp//vTY6uS9fLbpsuHmABi5rohsXrJV8sgZh8
kSIn4N2hKCOL7Pe226gZJ0yZ8X5+lu4A1OeEolLdY//BDGRMSMSaUQT/KErW6I64
Ao6QEOGYj2U5FZ55z9qDccmiKBavcXpKpmmsGI9wVce0RbG29AmIYff82BMcs5Nw
cvJS9SeZVqZvvc2BaBDhLYFy+nEDo3bg+4LSZNsAABxMwlL+VZu8IwnatwzzIIUl
3JKjiLZT2KtTnnnuGTiyuel1iNglGhqbAHIpDUrnJ7WmFXJyFyB35u6mY8RrkbhH
ArDiSYKbfxK5hp66gd/zyLk+s6uV1whlNz6229vWltAjak/jtum/+6Lp39S/4In2
RPYhJaq2hAn647fYRfrur6P41kUWZNfvvfUjVtzy3d9whA4mBVw3htXoYBvFKw1X
QxWEvaIqamqtwra06tRC/zxv2kvTw0tQrgzoQdxjD5amwMtz3zieUc/bh02lslAK
1IkU1yY1mvWJSmCZKlg1+RyBx3qgiVb8C8CpCuaXXwld90bgRcW3lt3o/kKoTYWX
agMfjGuHlLq0EaMiFwG8MW8fULwW+L4Jkdq18pxEaKceRbMNPr93AMC55MJ6kzvZ
ioZJkONyGLOR9RejZVcYaJ0bUAvxwTap4FCLOEUwXKNcHqhmM7EKy43Z2G7B/vA1
Nz/OFdbgDX+YDUSKkXHMu6TSnRkWFOCNDnxftwEYf75a5D3+RrQKrceRe3tlpi4F
P1oTRPSCH+p64kAb0zwxW8YS/cFrLHRciMePOPlqua6/ocIBGdtOWgcmqZea+56j
967+nkd999OpC9WRo8nJryeo672abzor67nbIsmn/Vj76RRjxLIhiI76muCQXVed
AkyFFzpxrSe+Ur7Nv8U0ETLju2cla1RWHRaoaC5vCjYRmz/TsrLeszt3oNrGpogA
PsTr06dE/52wTlOOQjbylGKVHyCpjLXRXIv5TQ+lTRnGPKZmadLtuhs7Bbm+BIxq
M4VjL/m8+gqbl58H5uetS8MkX8Ri5Qykae5iv6k0uuc8Va5Q1Tps89zGiZDuqt82
mx8632Y5ruukJtQ1BqdpYdda1kYkhXVxechofkeDseqxJS27xVCBE6Y69Snmqr5I
5EyX3x3pjIVyYhn3SeoTCOSQcoPxJbAVqBqkap28exzSeWAjrs5V3x/Cm8MDKWLQ
zOfuEwLz4hx/1+z3AURyjXG1TV5P2oaHRB599NlEWcHLsyTbK2T9xM2SKo+2+HQR
TdynZW5MkoiDQOI4fQVhL00lZeMYviqWPip8bFGh/gGXH5shz+/Okxz8qCelTYyn
uVb8tdHjvuxp9A2/EnI6oWPRZXLPNMjv3bYNk1rZqQu37b4SRfKa02/P792xFftt
CcfedsLaxIXPoY+sgI10C1dD0eI59GHp/eezz40Ulc1VKKVSqQYnXj4C6qW+djkf
2QYmC/WXhXcao7HvkEvbS8m1J4MOEkzyxGjN1K57heIv+e8xJC92l1WNI2L+04Yf
XAFY6LA5N8xcIV15W0keZDnFeBijZsr00Tx6DmT5DFBXaDG3eDd2ImQAnTbERhBT
eTrmrWqjCn8gB6DQgSK+qp76tdh9citlicsEc2k8/RM7PlxA4cGfjPYXn1T8CO7C
gpCVFEsNmhzLPebs5+514xy8DOD6HONsNihUP1oYtNQVKJFIbmIpQtRZGSmnwPbG
nNwysO1Wwb8YJPX8/uuoLeqWMUbmfbbUfVsR4IvF+uyfJ3BNwfY+n5gwUHh5Hrt2
F4L9a4HpWmMW3tmbZWY1Arbru7D2lZyJ51yhVQOBVMRzmgIdIACmUeu2X4093gBg
Tf1ic7WhEoHfLTF7dpHQ46qZ3VuKBzF/OVUWTdmRgLQTccfRi6LDVn4II6i0vQn1
88z2HM518SitAMq4+3pkjx/XD/ozPGWAq2xVjEDIxqXFvK9ArX/ccb0lFZrjNrs7
j72TjVsTkbDr7AmEEh5dty8kCstpT/QkOrwX5zqzNubvwSU/P6Rw7IJ/gXHhmdJ0
YJi40nnTfvH+INsV/nNGaNnRxdxYoy3PseQaoyx/iiy3h4E9vQoMepHckXqBGDm2
wlHOd7eQiE7RmqDY4fDsT/5mzG8V/54P9QDbxbKOsymurIArzIsCYjR1mVCZqzD+
NxYBO8ZNh4vjNjc8vYqGMYT1+bPFbcXg7X2YqpF/EFObKn7NzEDU1MAU+PC2UU7t
o3t3inQ1HOxekTVFc0y6YnHREYw4htwW79bgTeHawR8ZudfG2yvkrYQ1/tmEXRO6
LA9Kd6UX6CphVwgLcpGercxj56AOu8lb+Gjq1jwOB5d1C7psSVVj2/gVVBmAd1N4
Gya1lXYodWPixkdT1SGVDojRdhblwhavmfm6C2CGO+nse5fPbSXO0L3nbyzdkWER
sUayDSSPWCnjGM57WHU0oIxKhdBAHMaM/tMnRfye5D2dIkF/XKBmcJUffJl0kowG
btqETeOyQYl2pfcQB21XZc31E2RuNTCPHheE4zaacUgy5cr07DP+1zO4N3MEiyPY
avjxBGQoGPgZMOBcc1t3xMZUi5SA4O9xQxBTRVMNLLcybMJ3apJVJqXKZh/oZGtM
mQfQvrpLrSDIucvE4QVoxGWpkA46LktvA3ZLsuG0ZL8qoZx1JdmrhB9dmhssQYva
UrlQ3lP1tw1S50OlB/pf9+JRNpqZjmoYH9oXKVERMAO8DJzwqVEpjqSjygdFblVq
D6L8ZA++CfrkxfR8TNcZKUNjpoCEzjdD3opAwR0phP0V6DUCUedkmIWOBpXWOsQn
rNf1Fi/cDPihT72wqVGovGfI37+I1WE7vPfcxVE1NzguRObxBTNTQuL1GHMDMlJ+
JBdPxMoOHRMYbfbKXD32us6ImmitTD1li6DCc78B9Tws0vyvKlvMiTaDJ4oydoU5
aPflSNEsBoV1ATBjYhvxubMKhMg5cc+qxjtHD9TqpiibL6fwlSMQmW6FSE5AWSta
jKGNGzAF2420RkwCDPwcI2ocvPuwHXt5t15zwpO+OfbSA/EPFJlkByWCS79Cpzk2
Eb0GW7CwBHOPaE8F0G96PwqeXucAtsOa2MKksBJqv+EQfcIRhRAIFqGdB1MwlrxE
rDZg9Yq2czxbFQ9cTPfnWLJRqvB0Zh8rj5Rbl5p+hiAj8fUyJg/drjcY1slRkA2y
XKXqiv5zgZxIvaekSYnOaHVbeskwG+RHfrRWIDqjNfSVFNp1wNeI2X6Tjp+0o0yO
z+19ph23Zzv8fOddzEAqJykvycIz3jZCGZBvZICgatMrMTjgEiuXI+s3io0S4WTi
UZ+WEjG7WPJE5Ur5GCepjDW0F/zXxiT3p7l83KERZKIVSc87X1cZ/Yrf/TEf0S1e
RX/wvl3a0PEjqKL/XemMlAV7DT3O1egVZP348E4EDhXbz/ii1/z0zvPDxboLgUoT
pkBh2VB910BcBAoL2LYzqqQpqgdj/B8aHqS12BHItOvTRtbDlCs2ps2RCxAUWqnr
BA75bB1Tyc0HyKwt+zE3VEo6g9kgyYuJuQZBF3tICYjfgKRDY6YgZLqVsv8G/+Jw
kQ5ie5SrfUDqnT4eJjJY7p3mVyJ2gTic5LeTzbodMYrq5Bc63wn4WYD60khgXM6J
5kNLSJmUEgJQsOKPPsMQ4LVfMW/i9Ocqw0HTbeq1LgFqifbq7L/ggutrjTkGrPet
8I3e3gO9VU3fhD/48810k3Zs7JEdbLfTzxMeYR+MJg5haHe2XmqU2xcwTYRx5GcM
rtGKwKoJNVy0YMy/J8EDgaMG6BzPEnsPlsMpNNUkEu3oBPQVULxV1O8kQh/JdXou
dmV7OhY3LNPQKqXeDf4PI5sjYn4xH3n01gZDnK0StumDjOCy0yek0omOALl1CKoV
B9MaYAknPIDxXbtzMWWGM69PTkjt6rbHVnG4/ChbUskaKx6zRjpcA7kYlL1V2aXn
bhyrOZFoTIMvd4hoUYTIjpT9wYeUoU+MrXOqNzf0h3SE+j8YeGkWjxCb399e3Tlb
rIb97rDDGC79W0I15jw+pNaPRx56fIOmnOs7Xq/iA4z9GRBvhIrRrqGF/Nmr49R2
VssXOdqlGTnXllVc/Fk3DrQwqd1C0S2M2HY2DVh2qBOhuxVtc2Fade9NGmpAUPuR
rhXpQHpeznmBEpRvvGx5ECT5cRL+SGB0xEqYa+YOT3cGZ1yqx9jxBbdzSDkdyVN0
6cWAqerhDO2DalWhETK2DgLamDczIgX+BLn7dzgVATHDgMpG6vLbKFNmsi4G62UH
8k4zrtYzJV8XWSj+zNtA8uRzzSZGWag4Jdl5Y1yAoj6UXm717bTd2ohPVbh57+cZ
rs1fIkxmW6pCbcSRucpdNixANJDt4UMrkRfrUa/7Cl4AhE6EX7vxNRsMH/R+NbVN
Pp6xb0KOHRtgIwH+S8z24hFJu0pd31lK2PAivjudnyXULJ5zZidiXul/h5klTVl/
DHVyAJxwC2ZNgN4FBiqMdlF3GkFpTkqdlAO3k5JB/0/QbFL5JFryZI2DTBC1Kr4s
QW/i8+h82gwefMnxkIYWLwS/kOoD6PkSPgQW3y16Vs435VzYttJZfd+1kl/qO1fP
bSsZp974fpc1f7w4Zw7JxIanaw8zDYDZ55AIJvmczrAi8WIxyfPKhYdytUKOKOT8
chtIiH90bkOaHmPEm6jXgiYKOO5xBkcAJ9tFhluMKKuylFljJBtZR8s95nuTdYGr
sCkP5h+UeibeVXgLdBKcsUDEJaGujQrHukUj2WQbRthz0KZj1crI6zL3/T8GbD2z
Htsg8i0FYzh1aACebRGu81y/+U5Ls34o1eQMx0gEIa7BHZOB6cRvbMIETJwKZO3g
HvzuZ1xedYRS70wxny3MFAqWKwXN1TNIXC4ronVYgnNApf0TcMyLzF8mzpMSs++j
OUSsXWZg5hg5s0FshvQRTRCWVp5Rg/KMAWQDmZm7ap0/uhjAOq1BZczPS4S7Ew85
U2UXfnHnipsyCIxTR4cB7YM2EGpR9Hekzz2SKGrX5FCgu3e4HqWC1Pq15PAb+KSm
su6AQPM9KbnLpYPvayZQmIclGF2euWlmYbTG5Ekj5aHagho2O/lFelk/3v1qBLa1
pysKHkTtCo8fOM/xaU0rNpxiZX2+wYo0yR8HOKcnwqWe99nlFKQ8B/WykyX65w+2
9v8kIUf5+UvoZLHhS6G4sS6IZy671eaCMbrlUdJ6ptbc4VvQNNNSGKX2xmSBVTVU
xvQ1sBC/VGQ5j0SP1LjrEL3pha3PZESCrWoH+QH054FuiPkgG9fjvY1NisFbhLfx
tFK9THUWVPOsulWSirxeyHbLiElQX8M5h4bid286kUoI0ZupNRS0Wfz8QnsgzjzF
BMN5SwEIweoZDmYJGbF/vmcb8hu0T4DKGKuEQjZtIK2VHGcWC0vEgfMZTxFDEMWT
PZkYC8luuNcQslgqhRUJ08FFgNXeZRCew/QyyNLmtSHY/jXhuQo99xg2Hkc9j2op
CCENh+pyc1m6FRkUykzenZX9avVIXsnMCSZPNyRd9/Jt8ErfFIBcbhdKbq/cpklm
Z7ZWmo+RpNdXFhcSWCBPddlS1JYUb3tQF4Hlm0YVt93EBYSSfL8zLhRALh39DPaM
CjL88cBF02nmdxPW0Kz7/3JNGSaLIBBu3/esGe+7ENOK+uOfMEKveiZIzFTrAQ1d
gwQ2hTXcglMRb9ddcydZJU4aQVwHXyV2U0EKB+X4mHdooBLdqlwL4lHpHf0i9RyO
ySbTwbeErJxn1AS4nMxEoyfyBZBpMx8TG6iZqZghzoKVGchtp+Vro6/JMHWwnEHH
peA9kwFJRG529cSPRouqvPB2G/NhzsS2S1F7eoLpsfAIjldgawdneZ+SILttlyRD
0Syt36AjLj0qHsIFKm0RFByfjd2I0h/d/0dohsBB84sx278ZewsTJ60mWTipkShA
sEI3axl7gRHa6Bd20fHSsGbVwS1q0w50Tb4JsMiH3xUg9tY62Or4qt2EZ8jXTbvD
o9HJDCq5BswAGTqocKYmGkcxDgtQ6wJ9fjfdqH9Ipxun+y8JFn1xb3uvd/ZVXsx2
UwKSQammQapryUrqBamyFp4kK1wAL/JiIQmInNwy9jgfRxC7G+hYQNFUnJWVoRun
21IsGb5MlFp+rbAEAMgMe6aUnkjQ9TtDtj6zbyCNFL1IsAERO996jPPPw2fRfqT5
t8/wrynBmNKBw3VWNCvLqNm4A5W1u3o21iCy/QTYfCFDDVejk6PpA6pu3EUnC08U
5pMMx3vXXb4CgXryw+BRYe/l1ahkPaCNvpN8hxfOqfvv1N774ubmCRvDYV3k+DC6
sSWOZHoVYdQqHuZ6Q4UqXrGMbepVAy+fdYy2A/tmRCZB7BSXsTHYp4A2ni4NNb+W
CFDONZKyScdqWruoxZ1atusa/Tb8GU/Qd0/BswDmq+9zTcht2xrjTlSl4v2Dm3ja
S2vxxil1623vtwvtSdQ6QmAz5CLcTgsyR/VBKFYDB1UHU8xtE2bobcqSpYGknAI2
qBDtH0mAm31vB6IQlopXVeaMPF4PPRss3s6WzT48vMUkKrhlmu5iUhWj/xAv0UB+
EhErMiSYFsHImh9iUxOSO6BVRHtou9SiLlpTFfPCX9iM+6lk8r+LjFALB5job/Rb
azB+CCPeZdHc7iw0l2QOT/etEpKuqjKDuUotxarcGPRMa2lZs5bzSAW80z5t4SD0
ZnUXSb6pZxICCTFxkmpYBsb9tri3scVx7gXqu42w31GWTejJQSsv7jwKofSwCD5R
Ff/AaWVhp4kqmbcF1bFs4uvzBXhX3Svh7ovHo+C2xkrSGfooJKd8fjLM1KayOD/p
pZRp1c3YyYl49s4Ey+ApghO5PrsuJQIw3ftX0FoJkTBWcGvq+lkkPPvVnpweHeTZ
J6ZqKRSw+9MIaZoCpq7Snbbe+k+hsJ7CCg9opAWaUK9ry9DiBbu9RmqMLMxPKPu7
NsfHek7AV3kKzs0gXgKAHPLtL4JpeM5BHInRQP2S7IrlP7klkhNfO14nlAJSf3PX
FV6GuMKACZzGFX9YnzkGXgf+N+OiA9FLDTfjNM5BOU5xZQMrUwQKKk8AA8Vv4E7I
mdYtTE1JmWLgVGKPCDpkeLl6wpt6N3zmmFsiw76fmjZM/gnmfl5PNUbHFaDTe2EU
WaueGo1p0Eqfe2tcr/TrwXi25wPgokJVwfeRHc1Pa5rojry73FoCFfGjOgJI3GUI
CUi7jD+BDfgp1HuuUj49nDPD4gGzlzS3fXsn1j7rmQR6DGnT5bfNhoaDziO2zyPZ
rfJ7d0eUpk5InqIAWxMw6NrXn0wdLNAFodBfZAVHjF+hjO1kl7dWXeEv5oNn81bn
H2B0mFYTL5uzhFo2FJ4t0J0Q/YmY7cL3Ms3S/i7qiavTxk+cbRpiK3BhAckGao6X
7I6V5C7i7J9umGIpRpAX+LW0yLZbqxpVUvPy5PKWMgAA7/TyuQVKKzK+prYYbMAV
60Y+WT2y0i65bk74jrdrcIBS7/JDSQCCE9waQ2vILai7+zYRQlhvpHm0H0MCG75i
JQ2G+AjfztyWjd1PaJtoTfv3EJ5eURdlRYsmRMcGD1q6UG6CGsvFfpkMPo3lvTAP
Xm+zvLFKx/od5S6Tq2mWLBo0+lH8cNF8coLlP4/BxhoBlfiUljqSx7FH1xD6zNKZ
nBlvdwPxb2jw08owHETTVzhlN6GStpm6eLAwz5slfDUcpE4aF8M/Nt/dPw4g7Neq
VdLRb1WpX5jECWwP8gdJ7z2jlGDCwOxTFUSZ86oZPyQ8UmP6Zjw+MAUHF1Bh/COD
5vRbWiFmbtKHqzQFc4I9zV40Jb+XHdJcdadtPldAIEB3F18rs0qWRFpDegEKxRrq
t9TM/XVX/YtBRQe6FkSN6o73jIq7T/grq2cCH/MfYAXXoLg7T6V3Aujly2PN72CH
K8Ys5N9wsIKqQAnqsnN7Q45qN0SheeF+aB/kf2M9KOYA+JrBfKStTEQ5JXJa0T91
QWrGvNufGO6LO5vp+j98fwm9Gjiv0P3rkzcF4uLey76xPaLQDJwMcf4f+/iH8+Ky
YOkLU6/XxFUjEAsPeQL0nt7xfuPehWdBYNoZhgJ306idfNRSXFyf7oICvCK0rGer
PXt4m1KFvt94TE9ov3EqKTAN0hk3pb+d3ix7UcGJkirVVMUEyb9Fq/7EtEFG/TcY
3LomgVX4ufrvsaaAcKKQimggHswbKNgBYNCFC13RovisJVC6aKarUdJcxtBSP53z
MsUSq7IA9LEmTW0NL9osXPZ1mJNTmmPHEVr1tkPuVcOF4Idz9AlTfgyfhmeePlVj
P6GPUfbI9/aNDy8lk5E2hpPV72svmUkIZkEdXd+FCb5Sc72LMCLuJANuoCNbvu/A
3kd19RA3DGNu5WvAdPpIxgMb6aIirUXvT+PADHoWu8E0z206496VAw4iMINRLXav
juQ4wnY15CyKg9RqPmNwaxjMGBt6PLzxwoRwlrR8WUkiDK1IJ2Ny6vusYmNXAuQm
3DUXC5GQZzSYedzUp2gHDJTKP/UTSepOGs4/68PyWyRTajnduMdCPRsgtxrJrsEE
80T/4tSiByRaEV7R0tkAMxGjz8A/fjJ9m785O9bncdulgNKmzBRCJjca3fbgEML3
rJbGZIG8y1Un59ffuZi7ndApnsKYs4ygoIVNp1gUjv/0ZtZH1y40f41CvkYhHA04
yoRTRT5O6BPK5yva5+zHD+GHUsMeEcLGK1d6ViLepVQQqqfwt1Ysqv2bWvO9Lvze
ZNjmf2R0F+V3eqtSuRcMBM2DKbTW4fCo6hJVPi49MGwW/z487YMRWgTvTMMso+CP
VuzHMlJ/VnLLhudZ+rAeS72dVNZGGhIDVngVSNyp4yVAT3xorHd8QaZNVtwHB0HN
vMRywMhODth4cjUdwwtzzE3wWJlZO+nvc8p9Ua+LjjSiT7+MPwqw8d6xiz6jE3L5
p/rcxYjA688dIbu10ApUaQneFCjfDpKTj/nebEQu1LYY+wbhZSjgRMIlbuMV2lKs
Daxu13dp9fuetM9LcW5uxvKblHtydi7kZX3eNRnUE5zIiVA3OW8gN2+NDsAg1ZrS
1qdtPR5LOQcgrQz/UYJbEbQ7JAXuVX2A0M8NYmxa2WARekAf3/djJeuHbjOIdHtx
kZnqsHPy7q/ebSocaJgOKJ88+lm5uIjwoMfzETPvJ8y1JcV5wfej0riNy8I+1ag8
6hPIwnh+8piGJ+/sS9XmeFu4lOwSctSLiSRI2vB9qGbsTYNiYhhOVyFdS3kd+lqk
5NSJT1TSb0xhTnH2vCM036QnVhgd5It5zIWpgbRFIyytAeBmP9dcUXmhb+8GEnJL
Z+oDlLKZg+yV9gcRIxM4o03Rp7c5jhFg2TGznemrSMrfyoMYFhvbWlBsPII4nTr+
XzyXI8Gco9bimzLdyjQzHlz/yM1Hz0Wa4vTPOaL+KGPIoRqfpIS5dKnOwyAtZzLy
cbgFPjmuECY7CGSwco1m9AVIEBFiwlC0tbBKsnJr8MLozBElN9eXidym2mWqGEJ7
NJJPcc81zXkQc3mcR3pLORUnqEExTY/V53M4TOdqEiS7HqTOjYLfQLHxVogy6Emn
b5ZO2ckNL29HtagsEqnGdbboSxbufHhtBfy80U25WCIn3J4xuxGSk+8cU7kTvtNB
5rsXL40/WnK22FnakNTpsOFtruXa+c6G1JNJp4S5qC9YutOSOsBdwQAfepFt4bGd
BcyzbIrUd5nsnpgNaDilBGnStcmxfEb2wScpCu/mj0U4AMTys5IcXLNeqrU4xKVt
HDCfXqNDBQRd92CUlB6ekxHQjUCxuv683+P0n/akl0gZWAon1jWVQ1N/bB4seEkb
9aML7BaY+88XRqd6nZEUCAXbIXNSQAh6TkWxV3GLI7MbPAfiuMBPXl7FflWQnirH
8L9UWE5995coNgHN/JAXO3oXNzoQqCeh9OOXrQc9WBtHrT9ktxskKktH/74R1JUb
KYgxQVMuT1ie2noE0HRrBPWleNTpezYrZtTxrPUrpi1uho3AIm9AglX/psPaQTvo
OB20iIwHau8D6ucL8lkPNMK+WTlrjXAh7IuI+gDEsko9gANR4OhNC5RcDsXqgFYQ
iD5p9hgsnzsJc+35v/u4hNC10bbQmtBMzcUG5Vet7UynJO5/6/gFkh/NQdY67Rl0
CsYIzvW//cjIy6DggD9SJpARRaW+o9GmM++/dWaOsMD9UnHklK3mb6DGzmdfqYZz
FeC1E4o1O7GbSro3MxkE8sRZ4Dyz26D1XS/eG7twwqhAbYm2zchqqxbsVvrp1aQ+
6UBrqHi9aE1/vgnR2gI4U7QONU5Tzpogc9ZPx0UU7S/Fu0n/EVl+h7M1uW8U+kvr
4krPl0U4D1fCbwIeOiPZ055KGUfvXUoE2bg2DaOEzeRXpXNfIDlZCEaFXPu/SQQ9
beAX9Mfro0osD/JmrheWeCbH7pJyYJUVczhUnfG/TEYWQFG2FZSheLOrPq1XrY60
Af7QZuBXpHRdPqKJyWgd3zM9knzwpkT+zUnTvaRxQ/8Ar3+/b0fjQjCjJC+kWAFo
hJ4K8HWn7UA6QWHDBYq0tg+LFJ56/WNZS/LfcOJ8C7YJJs7nvEzh9crq/+6c5BEb
bDyGnvZolyE+k8JxJFt+vwHK582oTVS1v1DZr1G0adRDzrFXINAKjjEcDsOrMUkk
dX35yVDaFhqjolDbARd1DnR3umP+llGWvpJEVgtRMRr6wiA1atOOkxKVJbMmFvGh
qwJzkc2YOAHSUAO4noHkwi+uU5bM1kfuOybgVqG0rPivNmNYIBT8bRa/ovJteKTs
QwVRrCtj7ZLy6lj44kL1WkBaBhb8I1ZjWCQ35SK/4s0RDLUcve9z9AsypsDJ6+Ev
Y4nWtUw9R/BuXIbQ+7nKg2GlcmPcyHqEMoUPjfKuAsAh5iIj/bpv6/JnHY++cUZk
ZST+xzfBNsgzOEyiAf45J1yMWqlPWvMg/fMr4GWKoKKAvUbVKqaO2p0iqbRKhs+A
zmlwI6L5yfbhMQh2wa99uw8xQqIscJMbkjzUF7gb9Mmjb/t7e3ZX3mh+BoCKf8xV
s9moS/UE5zHBMTYGbwJWEQMrY+544btgWzdFQ6uMFYYKsTUA4I125P37OTsztFpw
ZPFMGNiq1SWGyeTvoTP4LQSDuap/Vvs67Fz2gXazS8mbEyC81fM2CcxbzGV/HTsE
E6floCFR05c0N5FQZsiawFGu+RX0Wdd3JWHQ1RriX7YFO6K+b0BRsvrnbmgibuyu
QvxkfyeHECC/BZwMnXNbxm+W6NZ2eZ2LvaHHoI1DVca+QI3n7obdo+sSUEYcLaB5
3/xijy5t/mwotuzk0dM9hhE2K0WYwus8pfL0dF4CMoPTHQPxSMZX0Mh7YrwHG3pr
sCWiEUJNyohMffOuWmTMVW6/y3NViaDhQIPH4CO8ANYTXmrhM2G2i0/jFA1pmkHu
XMFtfq561IuLuNZuNw7kdY39QRV12EBZ1ucma5D5Dv7g+RkyZvzFVF2tzFExac+h
2Q5PVrYHSbYlz5c4xe6hW2hxNjMi3kP94YLTDq17Xzq13EtpwezsJTBVIFOVH73w
Ufz5Nck+flUnskXS3R/rRKUMnNCIx64HP1nViJV2aw+m9NiwoMEKW7rhH8KOhfzf
5jPrC+YPQB9BUI8NShFQ2Aatmt6AbKM92ovfpv/UfR6ZyDaHZymOokvJ8ZeaFdry
K42dUw08aOCpfggJ+S2N5WLqWQ0gZf/YRTzt0Bmo2J01ARhVNTuN5q43V/Rtdnn9
h2P92qJjqoiuglN2Pi7L0cXXqhr9daWbj02m8Ain+7giWWA+LDqKiJ0KjTl+/gGQ
4Xr9IXW2DEjueed+D2YmOnGW1Y2qW3pDmJFbKuVSi9xmc5bkPPXr39hDw7pas24h
AmwNDlBVAOJHZb3v/0f9ivIX/X0g1OgaDsjGa0bEM9+DIkvfSLvkiE/LiI8wXSkU
lzNCQzCN3Bbp6z8dC2uHGPJWjFFjbKA/bqDmX7IN+0gJlKPVOsElLhp2LdwyZ9GE
oBNqq3wYxKeBOSkKKczXC1YUjfE74YrMxpdBPoNCGgjTDhrlFzmTBnzegaEGuZH0
uo6UGFy0dgsGcU/gC7Pv+5hnmRoEEvB7Vyc1te3NEdGYHemadt81MbFxOqZVO5Dz
53GxasS0LcNlG+Tsa6wwqLdz9p1ksBZoUVDIh75UNDpyiKiIgLv3rbOHwHjUqa80
Z26Oa4caLpiKULVY09O2dGjcfxsi79tczEXU86Ak2YPx2aknglrHPfuwbOb5Z/+f
+kdQcs9MCimQOutg9DWsY6GKFLLZj4GWqaMjyFp/s2baIbyikid2HGK1kF4nB80X
Y25FlSXCbMUXSOvP9ooKDS9oKtRHauxHPAeQCMz1dNzNMBCqN1K804eV2aw8Ra+9
zZwlOJ4V+MyMWG4yZaIdeQn/wEMUcJGnrTT29n+18ceJbxjbJx+zQ7Jk9UlS5Wxv
BKFDt/vnkVLDkeMe4HrJrN/XBd7Vwbb4HNoJLSSIEIdiGxDdw1YAv07yOmhbhuiN
Dg7QkrI8QwmDzFn/doKFFPVEknmqXeDmhXhObiCUZMF90r7iP8s4MDEUSGRkx/ZL
VcfUR2aJ0BMOvIDW+j/MPppek9yhX/OENUuP2U8xB3wty6SmyNVHp+X0nsTBpGuq
yBn0u6/6gAMw1+6YVdDUi+RG3s1/cCQRlcm33WvpBU4RiE+m40Af108u3y+AGEqy
MQaO4rui0+/zsLYdxyCXZ/GwQx17vhhUy/XJ1a7m+TRAIxMhG3WRdsv2lCCxqFCE
ZI0YKsMGT0eBqK6hK2JSJ6lXHCga1eY2m8z90vMVr4vcWDVILJbbmnOXNPQaFxHP
URnh6/qCEupQ2PRJ9+2kahFugBsprb0mutSjt+4bDzdtN7Z5iAdSshkumxbDhkUC
mUozLcCp7dajEzPw8vYGCYQPF6A4mnZ+QVjZYr4s+Cg7gDvQ2mpCt5UXzt8ldb5i
yyuAQRiKuHzFkyHjbWwEOgxQrqDp1kzI8OuKBr8HatQSrOP1XvQiA6beMI2e23TP
THOfzZu8+l2bGTkfX65suT6hU+u0DThCROmIaWql5u2tkXxwO4BnkQTuP2g4zSoi
e8w2VFilfRNv+pWtzyKVw0TFUF7IwgfKNkNmvQF9CT9/Ugfs37E2IJQL8k9ILTu6
DK9+b+FfB/+YTwOkUfvDVMZwekXrOlv6o7yYMtZcd74tXHiB78aUgAnHfiOnE4Sx
pn1O0zLK09dMm8ubB/BiOZo6xmY1y1KW6tG5RcskgKVUBFi6RITneTSpJxjQg4FL
EQ98H3wcmiF0wJYPrza8dykYeABgn2zwcJB6o8c/aBIaxEe1UIAzRtJ97GH+dCe9
Q1rtpHZ3C8fNI9tsrJRaohl50QL1YfXDMzV5cq0CbpsIokxMa7mqGXlJ4hkx6SsL
m5o9rC4NEdF7/aiie+IKPPgJ+zZA1CJ8rKxg7ZULYHHzhi5BnlUeW8l2B55IO4rZ
hTISF1oOuemtsH+VtaSUv/nL7zWTbuasMPUjlLN2bVEDoo6wWfKOHnn0MHVVtqzQ
qgl4iE2MQx04xpi7k1LsRKYMc4m17ZvmMhWHC3F5w6dosojO+vFzq8IuMsoeAbBt
WvgW3R9ZPOvCfdprB5xloo8ob1vtbNwre/GBZ/xcn9E/qclM9+oUSWorCKHiNf2t
xiVX2bC2Jvr1PYlLfGahnyfXtpl62zDYIlOvxfoss9jUE8lPA99nrXA/KYupJFH1
efTzs7jGd99Xcm81g4rBb/Xllf47Y5wn2at5/Q9lD444uQpO8IDaRoA/6nHfSinr
NpL5syBcq9ecTrbQMTJlUTsaFRYcqBhcP3b2P0K9gIkhbjQ+FkfK84C+e2O4rt8Q
nZJuhduORFjkaxlUPdW5OYeB31a+6kWXc89IsaUX02ciocGUB7E6ikn0lQNgIS/m
KfWqveABrpU4wft+gSDSMVayncvq/DWG9mql6gRKeJH++CyNJeVem9rlTd2wz1GF
ONLvUB0O3ECShKADSEurZk/gFOM91/ahudrn/B9ej4ou6CdzpUzJtI3M6/VceNLN
fedSeMlOJA3SHL2BMKGjkP8KDbb9NOciVFY2XDi1odlNFOKsKxxliTjNcRwH0egU
ElUHvKQx3mRQ0KcGWFN/OR7h7/mpLxjumepL9xDxUgIUOpEdMfl0fq+5W258jhu1
KQzSbz0o/jD3VJMSKvtBnrOz7frYdrBnCRUtrtjbbmVxxl/sC5CkRA26oNBxukrc
VXzQnRbC3lVXFttzoq9a1hrvwXSW8W6HQtCdGeoVgwoKKhANepo+2PqiCwVl1Scw
8wlC6FeLjHyrt7Q+hPX2MTMGMxU0q5w73bb9jroGXvCcjXjEYuw68gNJsN9jibGZ
D8qsgjissqaQ+FbmLvcbHUq94eOOM13BAUr18G3PVW4TZnZj5onvApZVQFrs7kdj
RGIRjh3C5EKdQim53Xti34O9AbxXev/5lx1jbrSgERDpB440HVqulSZe/0exHxc4
sZ8PeeUFuwFW81SRKqKt0/v2sZMUyOo1dO06HHSyjCIMs6HkUwCi6UFRAnViB8mQ
OTvZITisJAN6O/7gxNR4nuItj4bcGU+o0D+rwpjSk2U5ILPIFxg+UWPUZqgcg3fe
odKLlcU2saSBdcZeSqtUi6q/TfOlhJ6TAfMoYmrvTEg89uhvquxSH/O9Rgk3YWvR
0esr6KmE9zkYC5p30BFvOWcr/F3E8vGbNq2K+n0QsDTR37js7ecToasBekiE1Fn2
nvHvm8qYeZGqo6wNdIF6qU4jGhMuXlJJH7vv/L/9peclqarjze8AO6dMG+h2CSM5
QijXyKEswPhMPg44Rn+lDmBdoh4I+FMyjmMVMf5OtWun0TSNrAwZ20v2bD9KhOZz
RRL/C4tI1JPdedN5cP3PPyyQNen/Hkx54rHp685hguN6yzPBT37vnLSa0clheAF5
UgabunlWdFwab/AyMUxrXy6Kh1/UxTzYQ8JsD5HOjMQebizBWZtNfBrwnHi5kyzd
SLUGyMw0OCRQftieVfMs8lEATfj1DxPXTlg4tlscTnnklhMwGkZTRb5NOM2GoqoC
6eXBR/vyU1Kv3f6BHZk3AwxgxqiAeJiKozCurJrayLD/M1G/3ehpaUe+oJscxu8L
/Ze0ObkL7WmG0BdzavqrFUJcVk1PS5Zlh5Y+aZIuYPQFnZotKPAEAXLMDxGU6m7L
F4k3TeN6S7jHCSTSw0eBVEufySYCht+d3nIo8XgS8nFH/OZgF5t02qm1y1zhG3R3
+q9Kt8tCwNl05RQJVn9akSsCB7J70HgwSj+7rm14OpD0DSqJErau595eKfl6KH4C
PMSUKAlt2+OVSFHwHGkBCBR+HDpvMwrMGy1LqbmFJByqzLTN0IdgiHRthSUP3x7F
+xqVpf2h/FU6htAacK1HpconIv6B7R//2SqxhLYKEaZv9Kv9Ii85e9Zkxv4/sa10
DrzEgD6sToHvlReP2bV0D6E3gSUKH7S478W/kG0p0ThUWsgBBqqedyWSOiTNcjH4
ePIkD1FsEXP/fK25HQgdgxSyMylPxiPQga1j3CnKqGIQw2PRRbUZx5zizUQqHoKP
FkK/0VZcZos02rjVM5pX59O5VBreyPG7G8QDTlU/pufZHtYKJroi47obwMQ5Vweg
tSQ/5y97jyeGBQFmHLKQBTzuVnwWIHDyBCyd5PXVBQMg0Qe1V9scMgw+LMSL9UfY
/YwPC3YHz7SA99h9IGAOpCCk7pFD3KUDPTP1VgDWQNkl3NqP6/aV5eP5x1irunDv
WKW+Ol8pGqkPasr4wKmKqJHiHXMHLOI/fzPHLPc9nWVtZRHQbnCTC8bvXHhU3LCt
kwDvu88SZaPjWsC9aFg3fM91UuSvZgMhcpxlDVEzMJhphHSZUmQKIPtGraS6wQWW
K0ihFyXFwS/dxyzAKP+pMSCO/erFOv60IXyNwp9kwbVSbdlqfmeBaRybN14ngfxR
4ajYU6SqHnwpn/u/z2klG6gNgej/0c04hWjJnGO/b1/NMEW/5BUloh2Qw/IGqmqX
d3l5mxHD3jzTUTsKBeEYfA66L1XlS/IYFf7mFHOF8C3tl4R960usWmDKPxRlOg+P
X6mRKvgJI3E+JSd/2tedO+EF14V4ejbYuDVBhjsE6QtJ6rxm0qVzcZcGNHCF9noU
FBNRwtmovG077wKQkEKmTKnWxIXkxAH+c9YLQlcQOlrR71PzXF1UXomaZwDiEXg+
f2FBM1jRF2heDMBpjXJpCpt0MJWGAc4ZPr1RbzqC0lokKcBzG9chITRdGBdk1YGa
mi3gW91YiqwsDZROinMgyTteFjJ0iDO7JwYnC7c8mYePfIuEd88Pip6NmziRac+g
svTJ+kkfofgBGXE/F2g4sHh+7Gi2ryqZgkCTG8lCvR6UeQEvc2sU8nDHSD3JyrX4
sQ40SfCT6ZoBgSNEPTV8sepm5YBV0RaBkqjzuyO1DWkzuChI8BwuxM4l+Qo6hR1I
c/BHT8BlUFTOTD36v2wMfcIFH3grxqra/GB1NXiA80KIEHEdAaV7/YOSbky/yX64
Yhe4oJfX+Tt8Zh9/33T2PomwpW+tcrnBGxmrgMznEX4OOJBEvSU8cXlss41JQvtT
dPZzhQ8Aqfv9WgfN/tTnCZHMuDKDVSRrlt+HTpOPdMz9t2zlj7WwNeXfssbdLLOc
Ha3rMEEwRkjeDyj4hUQbeo2P1I8SgXJATCA3qImYbPbyQbEltzfUr23oQhrTzZHV
vsV1cOkcV8VqhALkouwyXtYxMO9XRsyhZyUndJDwJ9NBztGU+NHFSCbHtBLvJLbV
hojv3Z2KWBjJ44PPb5HAEanpqpxcbEx8moBQArnu1Pcu0vUmHgukLZOerRgVwnVx
MEgScy0mm13RFuo0ey7xsBYRMkP/RKrvTv2Lisz2sMp8hg8rgtRNK+gHFouxQK8b
ioFJp67Gei2JHqarKIKu809nsPZLe0si+yXHDEGJ3z5E2LBKKgD/kfHuUE+GTIpX
O4B/ZEFJAkgIDbeS5qI8Mr/IDsPiRBLVETMkPfvVOJR29iYFv6mcEZPV0+7Mroby
6366TkLNw4f7rCNVJK5CP1eUiTrUh0bWaxoF4upn+Bc0C6kUYm0W63s59GRMH1n1
8hKVRnN8l1ArlWN4Hi1j0jUBeQ+FesuAHFKg+ovmqBQLWxEzbu/8v0Pydl5DbZod
OgRdD4Fa/FBk2iM8C79XJwIy7YFqtdueScUN5Z9k+2xbZ/BVCwKfWWbVbd7azwOm
/gT7k5L++oMiLZwChuRv+IVe8/Q5KqhRCAsqB3Vnr5VvbJI7WIwxtUW1if3GhgNM
DYdEAr4LkwiiqVAp+mgfkJL7w8U2V5ApQeW0Llv8MePKMJW8MRPo52izwrXB3XgX
2k2a/bHP9vF+1wA7K0MWG6IpXkqthNf6DIUe8F9v/c2bhk+1Y/Ci+4yRf+17EITE
LsvxhGtmsx9ZAmrWOLweHoFBBUmAyUMLcO5Uwx5mgiChuNGzGhD/57bPbkZdvZYz
znNlzf0tR5+5BcoJeMYptSCnWzNE0CiM/p2ghkAQvNa1rGkNAZl+2DyOlI6C2waN
QeNIVNb5ulA/lSo0uHRNenKwR9+4cu9KR6yUj7F9lHeXoVheZ4AFGkaNh1uc6hvr
/dTf2oV6eRHSts3mzs2YAXsKDXzrAHMHnnPX7V6KQwFHaYcWe+vF4G0BA4AIgdcB
UFFOL9aJM6uzTNbVqFueac/zJLXKcdMslUWQFCCrBQUM42il4BuAgiOdrZWbTYu5
B+b7hvNSUN+TfiZLrRfKa2qeK1FioZO0bECDqDCS145HA0imqaYe/BjOPYl+CERj
wHoYbhcBj7vVc29lqltXUyJIZi/Qsri13xokdIsJVU9zyW7MyG8bpDOMbKWLAYNO
sY/XjLZTFyDzuFxA77wPhyebXXvbY3loLyg6fFEnqDxpMJgyM2ndrIHRJlKuOeyD
2/QrmleI7vD4g3LHpOrYYKHlMHgZ9s8i1uo8g9dpIOc2EvOb9Q3U5py2XKXNN2G+
W6d3hJQ/QfbNJtHw66Oa9DaU7RirWBjfn5GuuiB3x5mIyWKv+nOpTTsc8+MnZDJH
8BwC4/TaPNM8DCpM9/OSmRwJ9B4I4j8jFqhRfFzDdXvWtbTBbyf+8pbrq4CoTi4X
j0GRLjSoAb3iAuQ0q2/OSyxrd06M75EsC0+huOT7N6sqPJ3qSqlRqEAVAB66Rkzw
yk4UKtB22OnASRLaQB31lAujOcz5OOseIViZhHS1js8u1o32FxQGoXt4/4ZIfaVB
pULxwfNae6AaZpI1/2LJVCEZELxIiQBIKvH/sstdifpZwOrjv+HqYepdpaXnxt+3
7HA0T+S/bjMVGfSN6CWx8rPyjm6/96B4sEs2wxLfdob4TeByEa8C7IaEdv2WKOua
CaRKqL9HpIFbm/5tzYi6n6u+zFoUroGb7q4rE/BWlSEE8DjoIsYKpHZYmiKtbruG
iJjZ91hmzhZ0qN5d/piPSYSieWmtaMXyKQeBT0oZSRyrUO8ihkDYsE4OSrCHT/fQ
7GbereITU+mM4cGK+evaAaJJULALPG7Rey6wcqeawTxzccZhv0iXcADqS9DRmDgt
HyQaYX/4DSV0En1NcGvQ7aot/JxgeWy7mBL66cYjWG2lTqo4bsWfe3Db6TH1BigA
od79FiTlM4/1GPw1KnpfaLfYhKki5Uk0T8RTC92d5/zgiK000TWeZULYURA/e//M
5Vf7LjBfygvFXYkcgkQFb5NnlFwxSp6+GVLtOgfWy5KNBE1bVB+Z4f5ellmkTKzp
TeM6517jwtpKPAUmDp5VXY5gacozDNaJohBKBqL5XTdEfNfcMs9EyHmdIPWRL7XS
+p+ctt8JGI7vq7KFd0mZWf1jRwVsP32BSxkXNzX+qrifSVNRfdeVBS5xZ+bJAN31
fzFxvXFIMSeCUFFzO6kM+uhUXnmclHCrxy1wPOKMHYM5Qw1VRcLLh85vPaLUQ1GJ
UgPzXxChPqCY8VLwlEjTob64VsI3i6Ky1UE0MpIOsn7Qyxu/c87e/XsnbWg3IUSw
nfuETED4N8hvqyeWcfcBZXyn+TB9P7DnwjAv/ettpdDAYnv3jQgRtjC9YrozMDqg
XPbetHPb5gLeUw60S89HAOB4c5xKnqexeJCXwH4YwOs92q485YT1FOBUK0Jc1HRb
vMLTleYm9UBB9AFQH8e6DDiR44qh2bqTJGMizdS+aHkovr5YPYluuOPsNOxq6ltP
YzqBDNlJjvDkWyCvh+Lw5TcJIbc0Bip9Q5jKnF5ZgDAOsnXwzMCBrF3i3VzIVACt
BcKh7X+fZyB/UL1FkBIPWpDW0gR+K0hwQRLDPW0SGWTnROkeEJsgIPuG2uEJ3y0j
Zrxrs1nt6Ww2Ch5694gyDiAFnA19O+O0r+h4B0XLx+vqlCaUNVGPbERW+jEqaAte
mtT6DtI2TG0OFlSvSEC95wJcerjOn4rfUkHygL0/VaDcbrNGbYtF1+Ek2POuf4Tk
ZSM0/zl/IE0+byit5q0AJ1yarrMNQq8stQz2F3cO376LXC9+cLWslvncIBZidOSl
bY/Q+gKSjMiGhGmXNfIMytYhRywER9g48hBiZAzhugURAyTX0dGW/b5qGskgL41+
AkJzEQ93vBs6vy1QVgrvTg4RxXkK5G7lAZCtkauUvAty0wOMFd1PvQ3e+fLN1gKE
wY8+5WiAJDHXPjcpOhnfesan2dfBfhNz4/zJoaNgWTfpG73Pnr1evVi6ZBK7aqXs
Be9ogxYI1qPKqjem4Kp1/4rmdris6c1YgDGPHnhd+8tg+HAmBV6tkQOiMOQuEi09
SjrQ08f7kCVulXido4O2an35UYL1pJN+zcfK48ZuHZ8p+ExI7mfgL9eOIbqm7oNO
6O7jEXhYYMHx2bHQqiKVA4GTeiT+7fXQ5AmsIVfqJ4J8DDQgd+fmhj+9BIvdy5+T
8WZKSaJD5/lzFbzjcPLsIV/DlgXs49DWTZmROjnJdVM2nD+65T/QQOCtO2OHT/SU
eiDj0fgYbyfersBRW69/1uB0bOm08bNS6/LPlcVg2MGEMN+n02paFrv3qtzYZ/+c
ZPpnRyYS0Gos3noHdrPElmgziYrW4qVzKQRznbIjErbKtbylYQ8XMT7enzv4YanR
m1cYfvx4/JroCDs0gHgICHV7Soi8LU2aFAyhz9JSikxi0wLCi3lYuW//sxUnCL4j
dCyzniB2kGmcHYrBk0cAi7uh9CXZWDM4BQ/57PKsU1kcHmY5RribJjVWo2Dw9FTd
N2XTQia+s8IDn9RMhtwLFZC3Cm9GQNqVNbSem+Unp3uMPW9eZS++zniTfxyPBi+m
i9X+ryyAyjv/ra4WjEbFGLv8lBtlHc44gAZ2CfZzs9OcsSfuEb/S7WuEv6ZMrTYW
uoJFsuNpex/0W+wwmq5khfqL7u2HTWjqrmfgFkhnEYade59F4d7RinfSS80VxGR1
+kTABDWWU3jwDCC6+VIJuXdF5iETZkl3AHzhDWS+zfb/6CNw7Df1umzl+QfYXmo0
JkrET7TlBY/hWpltns25zMCOCwPHZcAibZC6V3w2D+4AIxypMPq3rw96tiSi/HKm
HTr/KZmpG4x5OPaUbXsUU8TzXWSsPg6E7p5/PsnDcc+Fd02pwCuVLmNqQw8g1fof
EgUoVgIsTlJV8GXh+KYUC0y82qJ6MZhzUGknIYBLpNlpNvBeXiw/ran4Lyrq7OkB
ZO63LR4L9vuUT2M8GyQLIYSFlkMVo/5QB0dUgOWWIrfDf6lD9OQoUCrg3ffrygvH
1nEyBjdHDcstwkX+0LrtKjG4OyaIDMKOIGTjb0En/St2cEh9b0fb06D9ogTlj+bX
ThUZs1AS6c2FzEhDMMNXmqR/YV5Uc72FYV0ZRZrOuRMSmJsBstaaPcdbqT4dPlnb
mqwM/Dx1RFI66ltDKQ7a3bKFcU//Igyy5kfPW5U9z3XUYOZmP5p6RUSAuH7A7nsi
Bcsa+B+D1udpta6HpW/RYuPiGt89jE/yfVKWm0aqTcrtS+hZgAU+O40GBHxbh689
yoyr0BmHFQLKKGlC/DSDoF9ZcIK3qs9i3BlSageuWHYliXpjhmvfRpua5GbnzS3q
OlMZdO5ktgDym6syL9Xl6fxBqqwWI6ZvZ53we1UXbQl7oRJNl2tT9nMNS593/h49
qTQLxyOBfNVTx2wh+wys0rPb8anzjZduwCRDoQ6iTUcR0Np6erNI6n37H6bWYaPS
MCnfy7ARHvRCRd1wOWce7ta9IOLaESmhqksmV7ZQKpyXQGgna6W9LexX5ze+M9hb
TpFQYg7I8vqUMBkrJ2v3Jza9RV/TXZuBW0iFHxLAM4UR4glZmH3z0mcxre3Ligt5
E0luvDKdEEc0J0KiT8Qo5gbbctv3CdaRFx5wtZdrmEk5g/KgA8NfwKrEZo4LdKVv
nZ8T91/Yw65H3RDGiMiQhFJObV/tzA+WHIY87Cldn175FG1M0tXBK6zWgnCtxZMu
pKpDJXjLNVIXtWWZbQCpS9nB9+buIXtKkpP0O63OdwLW57I8H9eLd6WBxeF3Kelp
FpC/DWFYWNTzHFZIzm3f7zHffawtPKwCJAY716Bi5swgfpk8lQL1YcJT16sBgywY
CA2DxLe8JisPtuAngLjQhJ04Iq7VL6Yjyvid90abKsqD4weP5Fw67cwlfBXVRkLV
Q0yULu6sBbkp0xXAe2J91fSVvS5Aw1/aPVmhdbG8QFCh+A2pAFRMgXpSDdlCXlXG
psvdkPOa36/x4XyxTi689eg/xVKAU4kBkSzUzV3UouLz/5akoh+/F24N0NcTNm7y
N4udiHgKbMWzzrXe/XgZxagXJLbqPNn3+kD6BcolQbzImIhmjf4mEpyjEwnStDiW
ku2SwSQ6AobTQn/gHCEbEXqsowCkOapnWDu6IppQTRBnwTOa+DQmSVxhhfIYAXaP
JWK59kKBOp9T4q7EpzWC6WE3D3S4gazIH52LOQwKbWsrBPgR/vYtTZfEO1qDxlT8
wH7oG8zFTqSQiec8xby1i/tzW+VenBqVfBhJDhKVs15Zadqpq28iHRUzP3lW59OX
vhquFu6unvdPj/3v70NNodouHInZDOsnKiV8cusaUbtiEgTlbMJcZd1KQAQ+jXgr
gFcdCijOZbwfQkJK/au2wWPP+FUam7kTNCi8E73qw1PrWljHEt/VNrfzZc+HakBW
3igRNBprfez2tt56Ds85PeXtpKfyRNgsaO87lr6HkIJTk5qWNoNESisi3nNghpZJ
OPGBPE1xgWz0fR+dG4IdBNnihi1EZ2EK/pL490HzvgqKBfz0orwOW1U6oMRHqbLS
hwaFdijfxiOWxlG3/MB1bwnp7akbWj+VHSclW9EN+592SLXPY7P5JsMyX9QFmwRF
+LRwPAPLapDBvvw0TJZiPCXRNlFEkHp7+vUbBbw6ZTNjlxrJPCPJN8Z5Qy1MlL9F
2qZhgCAjIyvepeE+yBZj2tEwK4YWH1Q36miuXkVvQP7HNniIBTM0Bjc4KQLSyBnm
BTt+pRksBEnMxk/yZcncXbtHbulpMwYGOFXqqsqMvgX+Ly1WCYteRR8ViHUtSL17
zF7YVdNl1uWBJ7MgQheKBWixuXiFgoVmmu660Q9zuLO2EbmMpqkJjOX3ByDA3bbS
BPllne0aul395m6BQnINsLsE1JLf7ZljvQZEzJi+urtxkGfvHZ6rp8VFEJMFNJnd
FgzkOyIiUkq56W6yPyaY39RNc9nWoyFwtfs86JgVlzmzqlP3Xw0MmkgKbhSRpTWg
TRYesdK01bVbIP8OObOWBqms85gr1HtTUV4syr0/EqL4gnYrVc0O9oo4ctJxURh2
cq+uUkRyf8bRU8065foESrzBCfz6M3Ri1ZttyAR+260W+ang85w8umiYeKbXnm2m
c79mPkrtbG6QN1Gbz/tMuihO9kYWvts6e6DrBwtvo3pebuaeudKdbIl/Dj3aBat2
JvwJ7vGCoinCV3FR6KRFA1sBm/hWN2rVNjK3RNnVcgtDfSykqacXH4keo2xT7oZT
xk9+4ff6yu8rWdiUat5/KqLgv0pBhpgR6V4LSFNAsYCz/mCS7EZQSGG7rcva49Vg
oW2Eqs4w/uJzVMEB9iVI8Nniw6p3GCOzFD+t48jWlqFh0K9Ugq/MKJRz8c121zrh
6IhRX++nm8VSDxYHHw2h57AFTIdd21uUx0bxvN8Nwmr74xwCOL2ZIWRCamzvfORJ
FjDy8HsMckF04Tj1O4E0Vfoxsor930Lxv2SYArVDbR9oPt12YoGStQ0Zdzx8fDGZ
xb//0pG/e9flhTTaAW+n5hHZOIcaJsMfyaRud2U7TYoI+LM/zNNMzX1vNzBkuH9K
+3aP8e+Nkx/mnXlrvImcvzNgfIcjtcQ85XvVDQNYrwMVtoPsi13/wFVUTKxH7lx4
BNq4y2NiuEoXjCsDLhdvdcgoiYPXckkWTkedAEGuIXbekyipCoxV+Dv2FPIJU4y0
auX5XckxihBHdRfTX+O5e6xlIlfDBl8Jd4mNgqIo4j0Ih3cG3FbRTxzHYpmcwgFD
VW+5IW/i90AF9nMRoAYBnStaDAaatT8iT63u72EzOMOlftKp3Npnau8mBIf0dZ78
Rfb59fDdVRr4706aBiqrefrsn+DG7DOke5bb1ulWmZTEwILCZWJhQdL0YYROtGT7
eV1jGomd4rfAmfvTuduxD3Mi7ynmIgdMIXchWnZ3nfmtpuITnUbvo+xmJNfwOJ87
osUcQEYV/TCSau2Xe0mVu9XUAc7EjSANl4SC4Zkumv+xriCe7WCt5m2tvjqYacj8
kWyPjt/FsED0wBZ857D3fDAgZ9+Gldw4kBrFG9o+oLtZRBrlUjM5TBZv9DOTNvVH
JDCUEEIjJUDI5SNilh6DJArka1KtCRVoNOwH9a3pOIfxZE7Hkj3ctHkqFchEzdmD
Xupe1SG6D7KJVMcKTxSy68WzuB8h7cUpPln3tKJSpwS/w+jQpFMi5Tx0qi1FuNHS
OlZaUkqZB0i/ZHUg57cw9APB98+lVxnH5Sy4qllqNorUK9Ki1v+KHTEWoBfG9W5p
f5cl3m5tcoaGCnQ/zxkWhIndKJiWrtkeR/a2Y5GGJwTmkDgTnze4PULBTVhQIlGE
gIF3yLO2heBwGC6K21qGs2FvmX+fjF77wzv8bzevxIdhmldp8BY3an8EeYBC3mhm
cCrB3Y8Y3/pGdCFoDwFuN2+0TqYBOcobBr/ZM5XYoK7qQqfR6By9ByySW+cDKliv
6b3BHB/NHJXL2DBj9N+WOSTNDSOjgccg2t4juHP5GRekpv+H2TpHKnTV9i5rYL/h
4NzTfMYD2NvwbSaYgpfMFDqlWtlrVSFGm2loBB0VHqRDiFe12QXOBxffy7ZWn4fN
Wgny912XQ7O40uBwS83Lr3fM82P//NpTuzcMD5vkHW/MvUSxnyNAkiIBMzz3DJN0
vMo8e1s6CVsSo1emF1ocH1E8H9XTqT+qnFhsvMEdLU2aHe75MoxyFr+N0POQfe+M
NNrIeqd78VMm2CcFM49ndG/8goYz/Lr2wAkDd2iy25cUgZFYxrzqTH+KdYnRiNnP
HEyUoj+OltFv1IaslDlRH7Pw+21cYF0qOz5MT3T3xwVwZZJ6eenwDxhW4I5O2Qk+
0nebBt+ki8HYzigqw2QZ076nr48beBFRWKjzUKgxF38iMjUGEIymOVwO7612hPAy
408Q4/gNmudf5aM1HLynXz8RsaORDrHRi2k7ZB5TWM+hiwfMSwgwLPBUz2d6rqGh
umEpf6xdtgX/trW/DQRDZJEXu1ewczfEh+xNpbyQgzvVTVvohuG4/JI40oBGFwy8
T7dTIQxAdJm5sF3apKGs21sx3gxy5UcvnLKQz1Xxxua1vHJIJ3wb3Q9xcrVtq6kP
/cNMqvV9v4imB38vCzlsiLqFTMpRO3pShX5YoIGum6H7PMVQNRFmZTzUkQajEuVy
vzNNtj+5dGWrHdaxEIKARo3Y3H78fLjQoVwWZOa/YbgQUjyAPn/nzmvow3VUqLyx
fDMSp4JABscI31+T6Um4T0pEJtK2dQ9aYvpOSUAb2qUt8jyjPtPpr6aYI7yrK7zS
6o81Ipkfkr47BuhhtF3xYT5OzhQ/ZxC7xtqc8wK5EutO3qWHm8QbkPScDFKIkPyl
ZNvTImCw8/d49zxGHT9YQYO9cGlwaKH/1QvwFIZKeY/YNDwqhfJcucRjUzvhePRz
P9ojUCYKzajOFl0W1r8qp4uljnu3qCFo5nkJRA5mwmrCFBobeaPmwoQULmF2NAji
uHUphyXnhumSy4Zx1xKn3HcZrX7K0B2yLNwEWozDartGhm1P7EhPQj4xEWpJGnY8
sUOFy53re8zW4PIzademukbgV+BQhTKtyvIzy4eohfr1DtZW9g5gwTahMEW+sSGi
rlH2zD//BuyAy+kZEH5gK1O0wT2IdN1mAWLb3uqmR5lDusG179P7sVw2pE/YIkbq
VEw+mwWmEQFhZ8rcpDbtWaiuwDmwYobKgz3dcStVvgBUNAddUci1swaNEbl6gU1y
5PVziaA80KCQ5cDKhvtvmoPOLe4csAl1xBmzxQnb5wXd/ySwd9vFbTPUdoJjdshi
YAMRlCOdoRlxGNDK0sDWLJKvaeEsX6HAg+HN1M33uxLjaHpZ9VuYRhTpejoFBCnE
XIl2lVex+YKhNNPPnlt3db8YCSNpRe8b/tqSA0z7X7ZlB5i6F6wvG4yNdeAj73Lx
zohECicETYItdy80v4wxuSSP0liHZ/KAjiDePICy6VYpARfaypvcHn/9XB4RB39d
g8iZNmqYn0TMIlrIeUECvRIvO4zVNIgB4jgwTaFcaqEf6g4lfasN5elqCixtdshe
RyP7SxAnxEepbs3G/L9AXHDsQElmRvvi2CP6TTfFC3Pw1YPd/VPLwCvjlClDt8kN
IXl0x+e4zq04I6VH0Bx9mI9a0ZoeEZhHxnEz5kLL6e5YaWImE9trTWTxRI3XUGDl
B2AE7UTQx4qI3yMS23pkvrjCAFDKFQ84BNxuj7KOXQq/GSSzgan5d8SYQnjU48oT
58WJCUxezd93iqqsuoqcctlTYwJO6POy9dN6Z3UCgCGELrehgFznAjoEKCA3m+f8
zNUkqplv4Eb9ePNhwbeF2LvWk3P08OItggN4WgYOgRHbIgaYXxXnscs9kzZhs+gK
9Gxxs1RPHy7bN/wePZhT258XP8D0/FMMm45VGYQKtkZtfYrXtwFZ97sibj1o++n1
5Af8S5u0QCo8NZmu1vduo/zzS5MXEF8an6Br4MYrNe6vYMoERPT+nZoHE7rZWBws
0xh2xp2KtzzODFAhyf91xyZoDaLv8zgJwdRL+MPm35lVEnvEUphER7jJy4GcFHdM
smhAbN1uGLetvYvladselxNj2H5HENWImVuQPeL/cMVj44OzAYpvjlYU2O1Gyswf
8qWRo+2PfI0B9jpja63vl8s+4AehwyGJyneu//q6WMdzcaauBsSyYGTNfORewvsD
w1fIDA5KO1GlwfIzT5nP3RHikgzP+1VuKh9HRBtIpFkkc3hdsK5Ph1fEBcVbRUo9
f3CJEfRezYkyarHjiJ+CG+YEb7DR0OOEaiNB1Y9N9gPzneV7VFwiA7wegjL3sc6E
ujzxdlvfzTNz12XY5m5fdKu4feiqURylhVYZhZpLFmMuTRUSRCB1E+9KKg8Cbi9l
721JCQmD1nWjHkBjbdru0dOVN2iP8n3S2XzWm4nL3CyhLHOnZ0x/16tuvfQVr5Hs
YX5qZUULJ7U4RAHLOc4JP32lKgLVgHmR5Unle8oZQwe1me/8qrqvHm2yXCO/LCFe
mdBre424J4gptOKnt5MqnBnR0cJuvf9GUlJaet53T+aJcCyQ0m/RLmopRHG92MQr
Bu8kDxwMtIc07QEO0w3YD3a/12tGLVQVXuPsT3N5ripzoGn/olbhxj2WnJzqZ8sG
mdM7y/wP3Yy+AIpI7aDvs9nVS6EDWz1em4nOX13qATRCM5vlwU/oFMii2Wt2xCWh
Djcw93KihMXY8y5jm/yOwapi55/6dhqYaOI7jKQ6LceKHljcqdc/JV0+qB0Ld9my
jT3PSmurHaika5cEn6D6Q+NYgurgzNFJKHkFGagOcyEukf39OVfNtSb+3mDRyj0Y
bjILpfVJtny1adD0LrCNZEXMISGeayK9R0ck5GCoJSe9GdcoQ8VXAIJUjFb3l2YE
xEVhPBg7S1aaAJ0ahdvAQI1vedvyHpHBO005xviaRwvBgu2gECDtIDavI6XjTvXi
1G4Yt2zIyEzjdDzaVE51ZMWsOt1AJqQOKU9vLyQptoMsSZrgo6WQFnAuBahygcdZ
E+EVSXE1fWIU542EbGExXZIADvulRgD1QbGiXeddGRjggBYQkboFyYoa/XsvNoF3
FNaYxNvFUhzm0ta9yAg18HEd7k44RgHtEJ2es35xwtJy097Ujqk7+wT98vDwd5OH
Dw+ap9r01z1uvT/j23v7fTPL48SYQehLCCvyzhgp7VVcsXY/56xh0Xp6U41HLzRZ
RKBKf+D1QCfthW6MAeloqX2x0GFcIYi+CeLkKAiVOeRqSYx8vE+vebD1/Lkt9D6i
L1Xdj+MxDZVmkXvS2vD5U8wI1KTKD2xJfg9zBGvk+A8DFoQyet8wdj7Jbfm1TveI
SPIH6xoPzOixbb/MEEUjuPX9Y3+YsXTenySFBAGNJl3Fy2sPTAUyttV2PfqjnW63
DjyhOpp3xGVy+oQ0EN28T+Vyg6zJhDzqWSK9mY23Bl5F6WB32pzKst+IoDPkt+Xo
bD4LH9PQDjorrZ/lZ+O1ThfomB/3VVci97LwmTGdFHuIoqR8hclrKtI+t4o7NiV8
2VbS0b2niSU3afJUVV4XLGp6C0PiLlB+CXa/Vg5kqVtaZ72sAk1+Kf2mprTwIKrE
JkHyu0Dt2A3PunHRGT14EBEpUN4o6TSS+dK3DpiBhp7wJADNoPG4RuDDHMkYI2B+
YNpIKT06uhqoYSmb8p6kiF5Fy3ALlGm3lUnjBJ9rOGL7x4ifGwHinPymqZTe8ct0
1eD6O1nPVqO959yMekcNxByjzBh07prnJNn4v5SiTsfU5ibI2LqY+1PSoorNVzXq
IfcvnQaBy1V3jctASomfud7WpAiL9rJpcdZ1Pm+fJSY1EQ5BuV+0gIc4hAKTxyeF
PujWDbuaMx71CzPuqR4MqBS+LsRhGUkNrp1mWv4bXgZiRcyG90JYYvDpumpyLdx8
GROwxDJCxrvqitFV/sFxNOOivrpm5r/ey8dPQ3eQnhl3dYFMHcAru9vuHtYYiaUU
bM7UboskOwQpdJ8/TxkJK4wkJdMVUdSx/6hkEEuGRMmCe4rK89h7oQN0HqMqsxPL
gTqimR9bQveWRm4Lghjf83cvnSWKifuZU3hDIQCsREsq+eho7aDIQNIavRvsFvXR
oE/WjnSv6mAhB5hWDvhaBo9Z2zyQd21y2ENOmYbHRneQRLZYYa1zp+eJsvojebR0
1P1Jy+nLeGnOLjv8NfxVKKSg7lqOfcgvKh0yqWDYr5VGZUqjW/IJwjzzeEOENJyd
sv9D471SdZPrTTmRtlcqGgHMK46YQPf8cLmYJNJxaz/JpJ9MPljtX6YI6oodnFWX
w9BCElRqNS1p6GGh8XKVhd820wRKPnGCqPyJR14XEzDExwjI0mqiPEkhpgVPbg0l
gXxehH6KILN3OpPCOKJfNZURsypICkCArp5r8MUh78maWkdTwbsrhr47tEpW2ePe
CTxvnrmOUHGDI+Xx3KB5HAE5tL+ZrBC8lQZZ4eXHjyziaDplo7dFtHo/3Sj6a3J8
v774OuOPu2Q+51fyQMkZdU8hWh0FLbW3I9cnhlu9UPWQcau5OcPLur6Q7suYtIJz
sJ0ZeqS2KIMSTA/628X6AdUtLEJkWLW/2uL5qmIfVAFSNMF1Ggc527naXsgVVEFa
5Zpju4GM9OhAT2dnP32tf/1TkmbfKQHWfTMWsKllaUqfa9nHaISUtU1SttUni1P3
VhUIt+Kj82NJsgdb9G1tfNK1tYRNrqcS+KiUEVXhGviDqlZjP7Cq445HwITU8zxz
5hvp02ECUpLp5hb8k7F+Svrqio2HSi/+Ij/OWiACw0d0eIeW9Octapoofs4Ct8mx
E7/C5phsPeh4Mt4CC3ajj2e9s/oX+nk9SGCE94u0NhRA9/a4+ArvmQNCmajJyI/e
VoRcHvWk2xftfK1gENPUWGz2wpuGIOOk4a1kPVwA+AZpVKV8p2Rp6jUz7tL05F05
GHhgENgxdCdWKniMUA3vq3kLoDHFxSH5Xd6Zbr+XQ1vJrkESv8qmPv6XP025/zzD
X4wqpESOEWgU7qvtxXlTr4v57WTMUrrVcT3JHGTnYN1mSVvXQOIxiBwJhI5yVx0g
67kgqHcndpaLj5tyoluPrfgY9Pok0j8u1rxFMutLqoyq9tVEiaDIVGxDaRHxKfng
DV1pyJJVyaOpZzBJhROvjC6KtWIILN6IpbUvs7nsZystxFk2cBd0PlJFib8Mb/d0
erE3/6iCJMj19+1P+Mus4N4h/CVZxE2wDfviMj5MCHv+sAKfy7OWy7oHzfrZmAUz
urHBrdrayuakxr9cukuetoaLJp5SA9UEZQ35urHAvplQ+tiC20myMpot+Ip6j1U0
ewB48TL24YNMZ5H7Pd2aLz6QNeEql2rI4s8Ouy72ddVKFfIcz2FO0w1Mn4PcVibA
uBIleXgL8QDeFLO4cG0XlCIpX0qBekm57wBcX0L2SgEEx+nN0PDy0b+ZkIlE7Dpc
AAllPrS65tYyKcyAl4a/xvhPvgHoJZCRk1uB64DBXCRrd3KTEstLZwU+hjBbsph6
v19n5uWg/QeFSPYvFGqmPSPIbUMh/hi8YeNV6J3AsulzsHvAfDH7QMD91I13Q1BK
QAiuDYiMuIXjjKnQ5PcwRBs/TBYM1px7u9w9bhUoaExxmr7sJL/h0Abfj9+Igfdf
Fegm3W5/Uhfvy7MsFP2tpxhoKqMZOnLTdhhwt00PZRhUOGjnq4Zenjw9eJ3gj0Zv
K3fEm93lJPyDAQI7XuK0fmLjG3M5f2XXxMifkbUUVj5YElVDh7Zf6YCuNSL8mtIv
M6orY8qgHsodDVN+NG7WUsV4Ybeui+eEGoZybsYBxHGFIFFxwHxGBFYeCxV3v5WC
Rji5X9KgZNqTuB5gvvlxB2iWDz+p1Od2PWQVrldgHUqh0ECxNP2htis57JS0La5D
HOyqvuCA67+wHoRojWt1BfNShM4HO5dvxEHYS7cUvTFQVkp92nVGD97IJYRIrjBg
g/UgR8HDSReqT1Byr/J8hj+fYcfiicpvZ4NRxqtDVYyxuUd+dv5FL7AmDuk+9zF2
oa4AdOg2z8K8rVsg5v0Q574mk+Alywp6qETRkOEj9+eMezc8XhhEG1/FLtOMg193
ioU92nq3KyKx3XYpWdX/qNvFcZZdwGz3tZB2Pt50Rcps7Jnxkp7m+9+3neRvWsDq
KoKS+//kz+mfW69awfJfl5cPX8F7iVF7UCxE0HhF1QOi5stBO0vzZgdmsJkoNgsk
7XXAhKuSq/hFJb7xQykTbXAdo0uCAgYztv0ltF6WlRcZHm85yyHE314OMgx/fEC9
m+yzXL5CmvZr5xF6aokRBb0JKt7DqpOlUIDqjoxbQVrvxg4UAoGRUPJu8xPvVt9F
AoIi0fh0yhLR8z2cSvejcIqcLziOBLgOtk/u7K6XMN+/fCBskQfTKSRDKLAV38ml
ZnuVBCJix/2zg5Sulbxz5PsnI3/lZ88rH334mM8MdRsA0JJc1TzZNUIsBA/Lx7iD
tzLxvRYXzPA/sjE3T3Fe63JZH+Aqa/Sx05JxjlzKj/Mw7bOgPh7lT4WNTHE1xL9i
jUnWJIkpFNkegKrTuN1+obMrCHhJHWSCgOz1X/mNc29n27lfIQfUAn2Z/APrp6us
PEb+8lHRooEnmNcDFNKYFkwH4A3fRXgw5bIbfpv7U6oqPmsY7d36RWTIbx1e9P7o
Bb8jW6Uqs2kD+A1BfEyRgiCKPAZJ9evs+tD19+ujADqVwwTsdAP9EMf1Y//es8SD
pnA99qHfswsvfib8AsoRFgbpOFGT+cCCixYskSLRSOv9xVJm8p1Y4Azm/ZPhfPCw
Ovw34thW+GJAYKfSD27nt3aY+OqbNyoQlrodIUNSKV4LJsNB00X7I6kOSbgveL7x
yTPaQt4Wys4z5B0+vXAS+qae4du/0si+oUKP8jxTcMWrhzNrSTmqkk2fF24ppjAP
/owsGaaIC8aKNddMlU0wiTStWovjzY481kQgE2o3dMJxDkKTBWCiHKEse/r2+Ig1
7AUOduw9O6GPe6N+MBbv9uYYpzgOBPfXys9Rwd3eH7obs6kPrWrmsK24ScrjK5fk
RMuNesN7oN9JiCJ9SbBCLH/O4xoAi+CRtFo81EG2j5AYcRzMBkpcMLDjm9IOYDuO
ZmjyabaY/c9aUt/Qac4VRMravl/B320TGcqEZOwTULbMaS4TDSvU+iJCrwiprpK0
fT/8D5srf21eR92844whT5h+QAOAPvD+bt5lqpYC9BT4PNDqeFtpkZpDxG4EzB3J
q6OjsR1xlOfI93XtjG/QagucFh6/uBgijHoTJkB3LtwB6sidtO4ZmaMHQYZA0wwD
pJaKlZjGfDYHNebMkAyaitG/+Mi+D6XeYVT6YK3BoWAUxx3Hi8qyujOVh/YjtqLj
u0lGV2oxC2OYZrrLKMRnuHQ+780xz4Er01or8IVkvpWGUYO/bkjmDUmZQ/kGqWsk
nNz/KEk0v2s6qNj2323CbIweVFsILYW+QXVfJi5rrv2J6f4S+Wg1ed/toHSgosvA
XcedkDznKbrPWUve3TkQpWRCKRkYn/oQ5VFFXx/EhMmOV7wCdR82qMrpZsKTRIdc
1Jc/CIxVl/xi0Pv+noNUuZxbBJtkR0DWeYcR9IcOBgIo/tmErMvbqCxUvspXgV+q
9z0gK9B+dwJl5ACU+jNjruULWUq8HwCnCyCGM8cD6hu6o315eAT34QqqVzgJ7Pxl
uiAI+EnqHmJNBdFkTOEm0GGENnN5sVP/clGj63pqY6jQs8ONQNewl3QL9/79/duY
oU7QkLTOUC5q9vd8lai8UjtR3irrJd/RsLDjdK+BVpuCf/erbZdwG9/ysBbQIyAx
hbHrG5ewLe9LufkheO7FJeaCBGEeQKAoO798fJrPAo8JNgHEz2JQf74cOgCCC7Ox
aLAazqAeQl4RG9pm70XzsBPJKKXwoCqHTuKV9AsX3nMnIKo6RhqiCmEUwy2RGPQP
Rtw2svd9A7+tk1uPYQDd0tbt/f4npYF4V7GDMCZ+mTPINlY0BPiO4J1VjGEXgeee
8vereMsucIrP1WH4j3iHpHGkxzpEG7B6yrwf15tVb8meJnDp/BW1Vkqs1Kaush9k
MoxVqjwVMSbPUFNX5OPAG2irTKCR423Pzpu5vSDNFS6YokER3yhXGPrSEhvmrBWn
hELTcCGJWlwiV+m/Wae6Snn6mHAswLrg3RERWtMruySAHpNiFTFnu7LplB0E36h5
Icn1F2gqUKbCIaZzOaYCZshxRsx20YKMlp8IcGz3Nh2UKVcemvu7DYDeQanKMrTC
kOVhot/fIEZXsxEUjmII3Uf0j8gMoL7SEYl/DxLW6aNqqWgfkY74UaBxCMx4AkdS
v782zQzod9RSY6rLh+3iCLHvjz01iI0C5rP728IiIAE6oj7QHgef/BtrazkIA/6d
lEibQHAQt5GepFEiNGKJioHlFbG99iJMXuNvTvO0eot0rwWH/4R4DrgQ+q6JS4vK
4r0vC75BGqzT3RbP8ldaJGKg4CcewptcLaUcO0vFxANLy7UMSrM7TWbkaeh6of/Z
lTHC9WyEVsk78cCDzlkJrj5h+5EcePzxDHsyDJHvO4wtuu4h6vRGGZtnW32ndDR0
spc5pezU7gzTUHEbTzcg/hP8vfj91CA2Vh8zM0CwdJfr7h+g5xQ+qVDuM+2I8u0o
fnre8W0PyCoyqI6ow678jdNBsdc57ra9SXWgx7ZPfp8+DOKXYm3Q/mj+C6sV7OvX
BU/2hw8YhYSRfj1a3t9YE3tC/M5zg36dTeOE35qMsV6xzjzws16UVpvGcc8+6UMK
gfcj08puIGN/E2yYy1ortCG4NhXNQ11ecEZDoaIt00TGLS40x04Cza3PeIDMpZBH
QFBmYP5YDKhH/z1mNH+PSg6AeH8X8gjscKicw2n1KLjzS1ifmR07nT1ydG6+A7fm
Fyi8fREDO5Y138TOOhL9P5QYNNy6Ezjh1njnBDHobfglBj74b5xQWXYo8emQM/Jw
4S616Q7bzRT97+GunbNzLxfFnB9RBLgC0e6lyuh1wvMTnA1kGcEJV6t2yaCcLJ1+
9QQAPTxxtMfGQ4TIG1yxmLMBZ/a6dbuXNwMxFUT9EwqNXkdS6+edtBYwJhAeXLO+
CCy+seO+4VDJPmc8qwmK1DDqDYhvzYr4N07jfbjQwHaAPRz2K38nWaLpwZcdlanI
jxl5FtDTHm79iynXeYtpz7vrc3MgGN2auiw+iyFN7fWH1HiNBQhNf+f8IwqYRi39
5COD+h4j0xK/BWVVWQg/4g7CvMj+DLyA7F5TcsZJ1W3FoQfZgrObi4EnHkReO19l
vhQKVj1XirvAtfTZQOmT3CT7N8k3HCY0ST6s1jwiSCJe99bUa0ONs9eS47uuCjCQ
5uqS0yebprXRd9Nklb/VHnSntzEzMXWX84oYocSECXKyo7Ff9fJpSDxWOC/aGXCT
YrDb8x4aWCPdvfZqaggpzHijYpg97rSZIYj9xCmDb4D3yEYHnm7yo7FKWQ3itPPr
hl6+aMUNSyMYHl4/VO5THNA/iSXQtbKcihdXrfx6Ib4ku8Dd/izE7OKdOHsft0J4
AqskjRGDeRoNBQSxkzF33NQfitrfignAgEYUpnP4AtfrvCkWMUQwz7wfQXJAoAMi
D/rTz6ohezEDoT39SYg3KwR1ZgQT+g+1mIMOROcM9o3eMV2HDreGyrEafJH11kqp
1vdb1+6H6yaFXPaiHtJOIbXWxHHE3Vex8HCD8VbQzC8Boq+PnhBYWy5xyMR3sgoX
V1Btw1E8FFALps/BSIajqfgLVkquDWIwq3w1rto4K4Beo00dMFgR0RA/1R+kguRr
oJuJVnGdHCvs2zwuqBUAfdioaomBfE1qj/ryId80/ANO6GWBNXn7SJnMf3tndIax
xBcZqooBnPdFAjvcYDX2ljG1qVgkph+s1/XF+nSNqS0A6P+bnq4iTKIlmm/Ri/wY
Qw4xy3P8JCmKbQfLoXjmygqhKOzh3VrmrPPoitdQq9CVR1mCNsOixjH6jFfMPQvS
KLwHb49SUuO5QydAJMMX1isJxd/HFG5umqS/s6oi1gaZYejIx9bzhdgn7ouB+rHb
oIIaflm7rkal+jfxDxBCskizVhKLugikz4PyG2BXp83qtyyRmhjQ6RD3auhK+SNl
dD8c2FASjzW5Cah96ZIitsqC5EgVBtABa1bCA4d9v3f0IPGCAuB9YKFAkFe79kTg
S7P76+vMZkGcOi5FlIA0uHeIcCzLd8qgpQRhwun5S8W8ReXqwcDOeF+OJOnDFkCV
IYL4tJCRC8TejUhpxmmN63FkYnM5cx9329+COwprbptjAqbyu2EKTT8KlUCRHmBy
pyPh+4S5JQYvBQxtuwfVUvH0z4WQAJHHVdEC6CkCGsZGdT1li/fj4t7j1QmmiMyV
OvsX0HDZYPXpLxNXC/EqGh4wp/ECvvobMuanS2wvr9zCn6781vh3v5P9oysKorwd
wYmA6iu/EYvPQCoRgKV6O52N7KG36MeXleg9Aua3sGqT8U8AXnETsAwke7kt5SCB
Xe6kjtGe3lZ/M9E8u7PgJLMNMff/UzL+TeyYPira7uI9S1pgIOhMRQHz2/We1Cot
TRdOliKMusd/zQ/L87EnfBkd5nSDmBCLlIhTTsp/+LO+eWj4mSRC3hmhO5sgx03B
qzRTvqYVqGPHvXkR+HezaU2zWcEqKrUxbZjSKDcpIgB18pzcbR9Wd9B9L879PPdp
Z1Plq/t+iqzR3PpdVWtU6dG/Lt4gTRsBxpDHp7aUvAQGZ+o00k+egr6/aCcMjOxr
Fk4gfC3u2nXVVubv1Ify1+7zA6pNcIm1FAz3i3TLzVGuNlnMBba64ye4INyzwGMb
HmhE6+xCTyAGDpHoQiwboxN1egQwmPJ3JfkHaveMj0t32f50zZAuG1Od7YqoIioC
b/a5YeFdd/LNw2voKS5GA+MahG1aPBvLq0jg2IZTp5ISs+lxhAvhCx4sosEHRg+x
jC4OJpJG0F8oEuaA9YYT5kMcGeG6pnnEb+vpEd4aB0uIbteCQ8hsvBM/X1i5yncI
m00hk/nHE7R93TqcYxAWGO77j3cGxeRG+7Q77Hru0+Mg2cOi0GKZlGi0oJqTwdWL
AvkJVlSGq4NTQsIiAjzj+NYpOUG4kEVqMH9j1o6mngNEvw2FHRtyfs6U0aBuhDq6
lbL1JQZXfLr2RZd9c9xHWffZtkL9x606QfI8yNRyHRZcDsMUqj+KUjjU6EBYZeF3
gg+OJ6suxkLZGC2dKSi1wZyeQb6lsqRDoD0W6US2n7zCNRBQpIUgTDfdM39fRJZw
C/ivUionvNVVJEjiuqzjs+QDNg77whRI2MxYIfDle28GgUD81h/4XeI9EB0Ck6zs
RR3XqwZ4mfLk4MBFa1bhnbku+GreM32c9iBb5KjETZ/S1KBvLqfe7PS5YlW7rjoD
IdaxytGRmIw4XyPcwi/adYGi/CVd9K7v0TEaT3ShnXeUWYokE8dnfjAifQ+ysKi5
WYeLh7GcJdP7+dhEY3ie/DcPhG8eby2xPEuxokitqjzihY8WcpBXhhG+CQrfYOAn
ucYXEJFYg2VxvPLA3jCQOotXlhff/QaY3Frm38a76qyiMilfK42mzSfWIzlZtjDD
JyU4pIbXNO0moi1cneRLX+NlK9giDTpdsmtr5C2RFLzRCvoORdWVY0IpITrff0oV
96iYvU01jN73pKbmW3TZF3FWmcphAgsXwOpyAzOeplTZI+GOCL0nOsdo7sqSiFHv
hAPExXzl8RglI0417fTZ6MIqyjfEn930B+I3tqYlVUFiLRsY/0nFgmlxtRYSalsV
H2wHyiboyroytEHh1AqPBhVpOKuuSW0dweja2Ll+9va/UsBPh4WV8PpjWWlCk5Lq
aMkeD1LB8n9BCzXoVuZJ/GHcVr2VF3RW8UPy2dq+GAdCdLgIG3VqT5vyacN0CKke
2IYc6KZmDUselLESyeB2CBt6kFI8RZtFLjtB7BMKFAXwLAopVsLGasNKyCF3tDwm
Se3+cYzR05xDzWijjcpBz04yZRli2b58/HMXlF133s8OIGmbmiimf1AUmKPz8WRo
aPhoQSvvflxWV6KM4072OBKgJrLms7DNmagtuMxZjbZPpyyVCUsD9GXX+Vhxxn7s
S/eaRP83fQeg9sIPfG/OEAhp8UrwM8yFhiVRKoDdqa6qupxsd/ZuJpRoDdSfayj2
YxcCvGVNrjTzHoX6H8Zb0KJdn1Hc5hvnHed4T9HQVhhMvb2bjQBCCDjRy3n2PlwD
iSlpK/Aw1c4jfAjeleZMIyGnOQAn4iZTkhjI7P3OESV6VDX/ttIvDmAh1y3gKxEv
s0hVz2XVjwmKJJzNdNBDpQAvWuL0n/+xL9KJKoiU/owNBbWPLh8T+i3qsEdLiHT3
Z8tSj1OydLEU/9Fq8anXZO7Ls54yH0urleRGkuO+0dUdHOB6M4sfmuKZrSPag7lc
hbx0Wk+Qpn8P6XirUdlXVixonuPFN5F8EOxtEqVGtx6AKL+HzwfVWBgBYxJ1Hct1
AxbLp8lZbmk188a2q6uo3PGlKtYM/wKQPnHdsWcvZutItQIJMSfFK3fKcY5LBeqt
yzAQ5d6Inf97McIVTpuUonIw6cfDKjyYi/Qkt3E8bX2z4xuznzD4T5fQCCZEj14C
pxSypygNo4m62An1/GRb6yYe0jHnR2/t0BuKrzvj/kqF8az2JzL/l8gVeOPeVmKU
cw7uZENdnG87rdUDizfY8ucIJf6ufrDjFr1FdjkwCrQ/yovt0P2x6nbo2QI3BeAJ
DM8kTE8FKUY+MMfWlrU/YlkW5oVjGt3aZ1c+6voJd69J+0LdCOjM5KCCOpaFrlz0
GVu/3X7zA0w2eJs2iWdHgf1fihKoBx3sDxSvCX29BP7CdgtwJ22gImLVmEXtSO/B
vY7Ncur9Nt+fmOt5Fgr+d7E5J5NNQcZsA3dqPTZs+TfE9Vh9Gjwq8QL8P25onmN3
2nh7srZrvCKdShy/LXbL47QKnLz3lyJJXl5UOqHZarZgQ2cxj1T8GX80E7LQUHal
ff0G0hqhVaNzRil3y3FtOmsuRXMtwd9ccrz8v48+VvP+GrhaIoiq8bloc82DgqaL
hbo+KpnWTkOu7bVQB7OljENHccvMknfwrxtIBnpt7omDRkpPJHWIMpGiLxafJhDI
TRxyAwWJLQVwRdLUCp0iLjHoIFrfUgewaWslp1qgupKoJf3bNwlNTtWTqjUHM1Kw
bGXMpxxMEYeKLMFv2GOO9RoHlM1drG7SN9ZOYdcIO43PkfdEkmOekXwhG9D5DjDj
0Ugrm9aFd+SpovW4Ek91Nm0y/1H6jQCuseJlCfHUcGr0lna9zt/wTOQ2tKTxD9Ka
RUoQrq6BRxdvPSgBEQxCe04HBwrs55KEIxi4ms9GeAv7wqd8ZCGqYIkD41zAhskf
tYeLHKuvDRqahLodQxTpe9ROzzbI9Rt67GR32zN56uXDxvRx+40mtET9dYPcO5Yf
ytNOt+Sc6JlDFDItuCqj1so9E+oew1EQqETfPnjbQ1F/eKRi4kx2y5IdcKL8hcjP
3geUKvmjkrC8oszqdQsB9mUWgInPZIQYKuV6PcVXWl8XUPHT6EY6wAJLvXgARuVe
32ZibQlnfC3/8iWowprFejVK2squHxDxWXo898OARGi7hATPVXVS4CcjFhkzZHIG
MgvzmyBqpvLbxRShQd6tbWKdcAZf6nMrguBUJFP/dGnmCdtR0A4tLir1mYMV/3+I
nC7npmRHDqTeheJUdmIrtJ5cs3ilcuVqsWq7TxuXdQC5seoi5Jr3cLqMb4Zvtkz5
eBWV6jzif4d/SgyXxhZESfClWp20jfEaOdqXUcrJi9rjHGAbWorxljsVR1b2Y2jE
0YGLhSaxCb5UnZT+rIierly01V8bXudyyRaKG4ya8Xq8FxsuHyhwZIgXfshUZI4H
ECFZ8BSvN2IsbtJFzkBbxos/8ZbrL6X5VvvP+kjJG45vIMsCvTelGdh7i2h52N7x
eXtW1uOt8+S5+7sshC/YIB/IiBGqWTAMe+0hWV7KSkxHXWUloKdZS1aQa49+lEae
wuxhqlMju06DOiUqlYIbJymXhBS+m2R0F/Sh/29N+l/vT7qgGVmwFBDjdxle+wtY
BRJDuLyzY8N+FrIGCP9ICRzJqrl8lWi6Y/sbebvySq88I685YOFJrgXGWrSioQQ+
b1dbmhQNuiTCS0jrDtzwFQhdtLuAHJx8zAXQb+u8o86BDMC0eoX2u3fWvVvR/htQ
Fso/WFBs4XaCbybqN22YHPAeXHE+8JPcOtoi23/bsYu49ZYLoH2CdDLNnFj+Lflr
5qTjhI09NR90b1sXAGNvGPe86nhAe35xXZA3szP5p/jUWEE30UG6aXKa3IdJTr+9
sKAyaDimJgg56IaqkN5lA30tdrm5tOd4eyDQpjYFnKXfnJAbId/GOi/Ig+sdg5Ft
ZMytiOUEXhDlaXs5Zbje6JhJf9hAYIaT8PralvJDq0FCs+fJmF8WukeFiyOLtG+G
7evhK8YG5NCk0D8HYyvqIe9C5GHrz9GqrpdGTbvzZ602FAMom3rvphzhBWHOzV3I
GyMJD5m+LHUqbdLciREEVdepmdRWvPEaBuvIAgmazST+bIIl+0iYb87sJCu+cyVa
Mq7zZ8msgYsaUz8VnsyWvqDy24l0Ov3S8HiARVvH/qpMdydRUjjHR3pgTEvo/UnW
1pP16vpNsvQaeCtLykPlRBylZQNmk7hKD3IQR5Mkuj4xCjDA/rYzQH2vsLe7CqIn
8nW9dDfc3pic50LiITaVsmgUdn6Pdni0HRPevnJaNOlvj6Zo6BCOYLOzKZC+HPe3
PHUg5cUpYXExkNA170txIEcKFJkd2r0inDsGxGQeLuoNbrNcnvwbIG7RWXHBWsmv
zUfDSIcJXEVugfSYpMQ9WpcLcnbPfexqsoXNg3erBoPuQnNjLrk1kG28Py7iZ2KL
quRd1BLsaH9d10pcTy1487cJ84rVynMnKa4pe8tUxizHYfTqoyrZEaPRkaDVgaq1
cNDBMLoIq2eaxxYcdbZhvpyqQ39P5+Eu3zlmD0p4JgtoIDMvpIfRGKfSGbtGtdyt
LZdkF+f4eAaz5dAM2MMOVqvuxDC969cYErh8h+aJI197uwZ71dApjopsEExZgnxF
0XIP4JoWJ/0WGhhASuVLpk/3LzK6RKr6Nwo0Ipy7Tz46uAmQ+oqgqIWAkxCOLBgn
zCb61sY+gAU/uFCM9mvxFRpu0aFq006mZnicCnDNJkSWJYsEB5HInsG8zKEzwaTp
jT5oL07TU19X9OogLYqyHUGklwvBaAXcMmdkhZ+BcVXjOVSsJeDbfBFuUCp4v7bU
1qPg/vABzxpiwuUSFagOZpRdMpqxgnHSH3GnuLr8ON92DvhVjd+PzLaS2tm7yDpo
9Q2W9IKT59nKJsFUr+jG/fCVFWMkGMsf2KGdOXfoxKw/Fr4G586WNQuluF0Dack8
B2MCzB8VlOJoSA5CofUjb1BAHfWnxj4QArzNHYTpKdqtZeAkshjALkJHxmS+Bd1t
65etsmth/5QLRWZ1TgtVYr0gTaf/XhrHcxdQf1YSiGqbl1jy4zWc8XthHTOnBBS6
RooIIX4gIqeHQ9qj82e52hETqpC4Qe/zbuDqX7Dfkz0IGei5Z+BMGjlpQ9nqwjY6
or+DvFXmj927QrOtAHEGB6xEgD2cbdXiSuNqCdYDiB4N16vPhl4Jvi5JOexK/W4q
fwjfHTQvkEvTR3M0/5pf2jFSoJbwVu81ECo3LaZ5opF8TMCGvZcu6EvEcbefimqO
0UFws2hxrmZpCscrlZJfpcqdO6aQwFwT8fMFMYy+1gkK/7LDNFMr41NITLhPm/wB
dkOAiceq5ErUUg6poYFzG5P/EHJ32f7wymRQCDWWMUCiGEnfTa6DppoFxAjkVpB7
oDOfhmvQzCT+8TEBgOxs7FG8So6qoyzAYOCXVfjEdIFMoOYxZ796hGdxmn0tIpZo
76qjUccwPLWVrDvNwHOKAxdmMZOqWiHXYFuEKK05LRZb+wdGRQvv8iL+uX4L2jvt
qQSoIurwz+LR/wFmTJBG+kgrfZyyOteS4o863xAp8jth7xQkMAE5xw6uHyEUwELb
qa5mLQjsDVeqtYTuNQu89upxyzusN3vPeziSB9HqwNKsMO3gXggi/75B2MMRXzNi
spFOu15gxz8U5Sk0eaEXvwsLGEOt0btBsNLu4k3vWrLnYWtyGxT5J9RS3bHd2/qb
TnOuDRAmpHiNie+XwFMTCGHD/Y406DUnzHvA6FLn1PRFMS+cfUC9NX6cdZiFsMja
J6xZt3U+ZoCHmHGrbiJGz8WQuBfV9R6/BiYV6NV+zMXn+cr0AyibFIR/ejtiWPTR
UpJja4+O9NzK7jYmtB+JE6/IAomk9OkkEk/nzkuqgqySFEQd3t/kCmo87Zjy8wcJ
Fik/FW1Q6AT0dOMtslxYO3/16poF3jEAz6MnOR0a3I9McpA24DR6QvmwiHR8KIgz
L7bUX5Z6k1Vjn8KOBXbFC8lKBe2PpSd+97Yt1osbCAZHqvExz5/8oQNI4XLsIoxb
U5bkdnvAme9LWkDMF8fKUIbdjiqqZ0f9+fiegOy/w9aqVn3grhNIborl69XvvkEe
L2teMCCwUGLA4fsgyybw+969lwgEtdoGSC+Q3arTCnKONq0Vv5e7y5OS/ceTTBmh
sd/TRfxeanjVUKHFeqYemwFuh5cVnuCwX30Ob+MZ84u49JRFOL+lR67+QpZAvGy+
v9AIOgHzYTlbtgA9CL5hAWWNVQpbr5jrUazWCvhwh3jfaawcmdUNmrjYDMBXYmPu
v0rNeLro0nAVFZYuvvHwF6XgNnDIb70vlw8zh9Qg3HmGUK+tOeBKpbKRHPtCCOHG
PV5bJ0+p7b17yaHIMvShfNckMTjxNypcu14oQ4MxydQVGcMQbc/DWSKwu0GClTwO
ZdlvOZAV/qxeCmG14sAMjsrrWlfryf6InCL5n40+vf53FFIcmx4SCkvib6nNLZUb
ublx4neja9DuRDCZ75eKygh2y+oKNTN+bm+b0/x2ziqjOyEEg1FRbnXMgKFXF2bg
+AzNnnLtGlHy6rgbf0IObBBTq0pDlQArc2eHVhkzVR9Hv1wmls3Bmnr5WZixnkXo
JoPDm9ua2NsXW0HSmISR7oBUi8XnMbYl7ED4IASMS9cXSRtda9P+EGajwW4v40WG
VypnVoWaFf9dT2XnK+3YKUUOfLZj+mpdw7pqFUuw/rdTmUuAWgjvSnjtUrmMmh6W
fJLwOxdDO3Ya0QnVpk0yBMfzYFAcKfVJDqdY1kPozIjZYVzCFl6aW11LGU4j5YaT
ZJLGaS9mlTkeOwceXtTexAzedBf2uXGYyb4dDTGtE9NcjL05FR3/9Bz/13GrXYEz
Ci0L3SMC/1SUqdbg9+2OhAiltrnyGfyzHj+4MxDygEM4QF7BrrL2zBaXP7q2tuhr
Iv8Tj5ve9FRJ4eZUnHsqUJYvU/sX9+ynQCNukPFFzDFnIeDQxX3keFNSzUasDYzT
QnLCBiNK6JXc4AyloAxdmXX9F5eg5QYaMGPNkfAPufB5JYNOJy7fsPaPoxOubFQc
tPVh0D9lhdmTFlZepq+L3ZaT3h3Ep9/4+6AMy0a6uZXxDoHF2EgVLrCY8hViE6oT
5lovmMZfGnOGO3g3PTRa5Fk2HaJlHcH2VShrWU6zHQu7U44nstVxgjxbQifPZJIN
BjsxPmgsHt91DI5YBm+h1x5il3YTH/wmDDgafNcg7NQDYBOJboXLjZDSBO8ryB7y
Z5Gwwg030IFAVcaVvWSr8EoS4Mtr+lmivjHXzPM8soHAkUr49peMMBaJdD2RWAPU
BDA+eWGXv85vjRSGJjMrLWxdiHfrBH2yMsJbuCzLA8OPy1ZVm2qXHdPQOdKTvcly
x+kj+wjQdhN4oq34gssGh2pWqk3mzJwsq9ZSlEy19YXy8Z+KLVAw2B+WtRB7fN/Y
6PUn2ggdP0QbCIG/K0DARTepREWTNgPmEWLHc3gqEo07PN4eyzXBG+hvz9m0Lot8
kn/KOg3RULfxDyUZO6V4WhSRAaBR6xO5GqtCMbAjQEbwGZL+D1Q5cQLzsvknDz+W
ADk9YSwBRUtjsVa1WafbwsMuEooj8V+AnXf6LcGVsH5vdz9tgj+zDA2HHO81Qz3e
wH9DKdJtKBgAo0apkp0WV8AHghUbNliAq6Z9KjU0q59qP7U+99NS8EaJr+KPnvAQ
AMeqUoZ7IObPOQAt6e69E1guVeKLIMBhoZ1oUMAt6Gq4px3MIyjnBozPV1ZvYrMJ
eJYpC5ijZM1mysLnVgLE6twTv1x5x7bplphT93aIYLCA4I4D8/q9D8QSE3k9eY8b
DwpJTdFl9uHTwRJsw8k46vDxmzfxqCquuAhE1oo0XaVTA3IC/0ogMK9tSxRmlBMO
LfyFXjNG1GEVpsK4FIuam2VHkU79f8uT+oc7SWoJtH+wHIZfM//wIkVe+XQPc4C/
UJ1vY0q89CxsOZuUIio9grdJTTvbk4KAVSCXy+HakxSmxYTUgWGq2nCxoMim1eTj
K4js5b5+MsrDHRxv6ZbSvMqKaHuqxBy7F0AM/hfbSDIZ3UzVa2DoxXS/paJJRwjA
xbzi/+FJhAbU/rkO6XU3TPlRRYdmj+PorvEL1j7nZ3WPJknZwiQI43yi4JnY9Tu6
yaihtZHykcpCNT/NobnGT4PqLJN05SIvl6itwo4blh2W3phO+oPgf5rB5os6Jgc+
ayRmRyi09J+bhc6U1jMtvl1PBA3homM2lxEiyn0p9pFse+ml535kfMPWHWLTArM9
14saFzyyist2FnNWMbnODAocanG/Djaq5EMOuW4qXUrv4Bz+I4JTmr1qbFH22xyE
QR91NZNodF4IKOUwQqsr08ybS8DoNWy+LrxdqZQ1zs/FYOgipq9JoqqtCmggT3na
AURMGJhCLPF8oxker5+qIQdpgSREqhsdKQ+Ldd0b6b0V3L648ZYMXfeCRHhB905u
GuCtO+1H00RznZFgwxHF3cL9NPwpGjG0pKWMhkxo9zpFWR/1iCYd66QWvmkgfF2X
GJzUTkGRPvlO1Cyv4z7UV2EHBzdgBWo/mH+GKqTdfb1Jip2AzpJGjSE7QIPWLYOb
9dF9QK8EQ1Fn/uZ5wV2LK6m9emDNhq9yIV26BB7MW/lTrnhst/KmbbAjbFeL9WbA
fQPYW+uq3QbC3zuoHNgpAMCoYGPE9n7DUbAVNvz76wpkwO29abDFjAwvWyB7Rjso
FZVm2y3kRuY7lCCUs/t6Ou8AfFytvgO4isJj0j4vGnBHpf4r++wHu+/a4aVAOn58
WG18VDw2Kh3Nzef0v9xb4nL00xXN9xkL6Sfw9YL3mttBkw7FZGoJB8/C4DPJJjut
7r7z8x5a8HSUbHZrFju3ZJz+ga6HtwNGgWRSJ76zz0WLz/z4JZUdwisWs2XJsEbD
FoGkdiTFzdXtd7iwtPjZLXlXUtQ57kOM8NEr3HGITLWs/xOcQOavIM55RufASqTQ
ASkGU+yzgj2/WSz3VFLgRwID8nD2BkBvT7sGJe8IR7WwZlCO/e5/APdt6cMFucgx
J7DUAciWvaCCH/p6cquTBEgwCrDAMtOhcQfXQfRqzFA92eLahO+XW0sJJrXoISfM
rdOkSZfuS2HeNkArwBbSvmo7ICOK4PU80bd+vRs3pDe0WeykMAnEZE7En5YM5a1i
gs9hOneNX8X4Acdh4/IVTAC6Dy7eKhD4R1JWSmfDvuNCJs4/ffZOOnUzIhqLnPWv
BmCzc7F+6+YXA9NM8+jHod8RjpVWsXhq/nI+b1DVZmLUoZtslhKtmh7Sv7RQHOrI
RdBl4Lp8+5RkvN/uEoR9v18TWdMcAHN3RomC2UlS5GD1Y2MgGPtbHSiAbO4ctwQB
eOHF+pj1KI8q5h0D+jXPIBAxdE1qe+oq6dNQTuqE8gIAjA/vP0Srz9XHQipKo8sa
04uT9Pa09phMENenkOzn7TaYDRhxxAWxqECms5e3AZZd5vpdkW9BNAyDQypvdxHj
BGF9lJgv1s+Y/IM9/HiZUFC0+6PJ6OQ11iwZofJKVVdPIqpsnROE/agQNXURSnDE
ixpV8jOiDW59wJzTXKl7rWpCbN5XYXU+txd+Yn8hC7uItd4xg2Hh2IgQlN3I+EO7
L5tLJjT25+QK3aIt4skajO8JMc43W94s6r6+FBUK7LSCpEf6FPjYFC+77pIQhYrK
ippotpDAlxVhmAbyGXYnxFHvWUxqcjKJjhibF7ciXx3pWCIinFGbKktwI3r4Mq9E
Mc8BpvtjIB8fgg9wCB+TDwrjE/kiYG0z357GPO+PCkeiDjKaTcLSX9NYgDNPkaTj
A4Pd6Mae7DU/1C++AnpjeVsZSGTORDsr6uJnYJsTEj3lfpZjXAp0Nsi7g8w68LOW
wqp7klUks0984XtQyV9ZQ90SX5D9d+2fcHRGJAwNfUHQLujPjkVH2WbAWZuZyrWw
nNi8MPUeY8OoZlJ4o7pfh8p801og4bToCe9BOjW1xGZws4p88sQA5hyK/9V9hftv
cyRW3VikG1RPT7znMJmh2ABXB5xEe9m9p2oNHSxleH/MnGHRoORq8fc6OllYbJYs
ZZAC5/zT6DR5ApIyWCA4J9W+4e9Sqj0maPF21j8RzcTez6bkzW5CgqLBhag+oYQx
NXeEW8IZe6fShOk5c7unZLtU/tB/Ci2ZFYfZVUai8acEaFbmUQcsQvE68crIOsDy
Xqv9EPCUuawLcJo9YRXP/LGo5Z5Gpms79pAa8z5CkN5JJ6x0rJuOX3eOxQU1n8fB
PAH2Nqude6z22d+1FxwPXNPFv9iRNTpfJ+ZyYSbTxYmFGdwBMf0LZJfjIhkRugru
fSI6lfpWSJ+6hb7DR5OQ6nchwgGadUbGFjDAmyhlWgWJuysS1P8Pj+KSnMsex5xl
bIe3ZdNjZB2P7a8o96Yqf2V/qw/kTZrSw+YEvWBJLF48ZOZDVaKvsHnZO4iu+U9V
niT1p/MDgYDw69hkCp0dfmAmr18qyjhH/fRodhitJb4fOWJ1GlJj4AcXZkZGrscb
AL4bmG4E8mCe18WcGY+oU0s0GIwEpMvTMmf6QtY0PSDXq+oWyi7VliB4illdphJq
7cLZfFIpgIzRyMwkuhirvXscq6eCNhc+jFMAwrdtYzQltELu0oZY4Yo7suVMEsua
L+3LraQbpA+uJ70gMPRh1DIYsz2dD0qFOcPP2idSpjeLV9Dys0XfCP59jDUNmIBJ
uV93R/mrd4ZYvt3Em2wfY9CJX+f2lGetepfm19oISOKlTBm88l3RR6//MnuIR3Mt
XgnvndGkcoCTLKGBCfGcHAVSdMW26NxbhtF67Fr0XDehxGicBvFozOO3gf32sXoY
71hwvLfncc4pkrHpi5AK9lhCmNY5LJjhn4aKmbUVJIgtkKCJRIZSljAr/2JxBB1b
Q5WRfgQYLUO8G4xOL+0p0C57KZxfzNmUTUcTmLSMrGnF76sT45k7URibJLKT9Smf
gxIw8Y0XQbr18JDjV1cubMDmRp4bcPYmoo+TA4tZ6adx1sj+GsLeqHqjfxb+5JdS
LrABqYr7yrj0cg/unJcv1BTBi+JfLWjNvNnv3idw4C+DfngHHuDakeHUlnuuBAsV
irq3eb+Vt8sCNDovSGZTaZWxIOcad9UgXVUqBT3veXVgUywaN5pdqcGAsXWiGQxV
skyvT4K+cpkA5I4zziVPgGROXcqmr/JuuuKqUIHTs/g9emO4GrGSSPFudm1h9g3K
dQHO41/IAJOEs27RCpgkYpmZ0E2v0pXS9q+I5xjp48yWkOywaEm+zXBX1iDxZW8P
NS9SHBUnf9ucrX6PJnJNjjm7Lyv92XpNKfKa9/AvsFSi87xBAhZWiTHtRinT75SA
xqyf9ww/c527tZKAsJtRh7zJg6qMkP2wOjnjRnDG+mhwKo8qEde79sPiA5/Ky/7f
E5ClkRc5CAJhJ8cGQMBOjJR6SDhHLJKMbgy/pEYR2hDJHQkSxu85iSGlQf/m+dtd
tdDWINvgKf+j8bh6C1xOEXtmOkMlv96G+NrWf5KDQnG5PYoCcc2Mvj5POi+mns57
U13tIqrXl93FKBJ5ZZ/JcxE8lIyljDGbyBgcBuwACk/DBRZb3jERxZQvkGr6buJk
A5t+JcpeAgRV7lQvqe5IfSWCLV/zvITaQo7uFgPHRpklCuvdD5QXyL2qiJIUcCjR
qFK5XFmjxrwM/xwBOK+FiWMvDIsxYl+3plOOCOHEDje3Yw+tRIrehI7ttA4X6Ai9
E44ajKQQ2d13HnQaBTrjK7CWkh1ot46i0AZftRRdqXMnSMsjTPc0Kmu6SOex0jzv
CBkxJ3Dvu2YgZvrdCjKm6EXblgUgNjUFJC53nEfFqHhOgLNBzjiXBjH+XNKA+c4/
JJAB27RoOrLDbKvoswslOR/Cixyjb4BIL1V2tVb+2lGOsGSFxo0AsQaDIwMvtrmJ
fDJsIGKztD7txwGJkm8dN8jsbYHFOfRnlMF1bNxgfUQRqTx/1DMb9HueqyMfPMCs
JdTWQzJXpbSZ7vsr0Rt7cwmJu2CeavM3SZXcDHcFuC6z6jpBtOPwc20bYrmip0o7
x8GoHRlJGmCjliKkzcLhDjs8eXiDSArPQii8DCujh6HmLFoOadfZT2Q/9h+MNaby
1bM3oD3unJa/3L7S33PuoMj3z9DSgGY5kiW9E4YFEytHk2aQFBQGO+6WuQqdzFLo
uDIJv/pglZFj8oteR+RgQh7Fl26+x47xk7jDzhn25YwKqksqrhNZtHLilx9o7wy+
5kfnOLMcRlj21JCH4QYPGFD/RbFl/sSjCFMdAu6NGeFKyuAG97kFwY7lbklC+Nfv
hV1/QNa7+y2C/Ki2AOJD+qKpIMYoGSN45UZ6tFSsIUcjIl3a1i6OdyrGNK4zSvRX
8PGkPiRN8CwEvy2dRTfBHHtgFt7qDXCpPO7a+Kuey8cRVfyu115YAB4qoRBD6MKx
zzuJQSoQdJFIsS9m3n5XoTogoqTa16RISXGnAvwU3O3WR9OS/UyUhSX22nwY8LSX
C8UYPb/+SC25xVEq7qDSPZ1aly5R4AGIDkFSDRPyEOoT9+B6ybcEFheMF3GhPUts
MYUmB1eqcNCnApd+4vaKaLO6W9oqaWnmVmIJdZIUsFB4nhOj/nsgd02kVZQ3iz30
o58hGCmk66y50dJR9DBVw6pyUELf+eaSYM0BerGkaTUrp611dVpQ5SWL9wzOpwkb
/NHdxKo9pjsBPQi4dDmNW9hjV0FvI54Sc2Jpbu0tqSZIUvDcNVuejKF1mQdVXId4
qxozA8qiRC32k3a+zOdDrRnWso1h31z9lqavmNQK3eboe9ceBw1i9pWKFUZyUn45
snBdsIp3FNi1WyAa7yh3Elp83ur9vgBBeCBqWg+CeTKin0N1UmwHUqR3azaSrmRC
ziFg4jjZIhqdi71VDdSC1nQxe/7LN7Um9ZD6Z9NPVyBhOEQVipAs7fYmdJ8w62nF
e0KUzGZLh4NKGyXp7Yj2XV2A5v/cjwZF0WMGz3wDvLWOX8DkeCThsdcgJgyUHvK3
jCIiz36J0/XA82PMe+RLOwsVzAwwRshIq0zdzQYHGO1R7rg6afYF1Xh5I5K5reAg
bbpbP0ASq5KFoy8KFX/NhGmrjomQwu+HT7Apic9xkpEIFcOwpvEDtCplyd8wqTOX
GJKNy6RsKKjtKuqil1MF9HSIIm4AojVvhk8+4khR2SgPqTbyTRGLVXwb7XDSsfVG
kRSCC9nYA2uH7XefnzuBB4If+IVLUI2kKSB+tS0Jo6Qugvw/6dma51ZnmJqimYeS
iihGeDYy/mLiNtNHFfMGTVvHoemAHEy3itpC7RUbRgkEyOKG9v9ueaQ0UHar4Izm
tUBZgIbKuXr2VXF6aV858M0HJDCNKZJbjmgG4imJ60S6zQ4UBNVP8Ozfq+sHZLwX
ojkeeRNV99fp2iMVBW3ns0uJAxKBDbWHR0Ha2VHODVhEvHaySBtuAr5xxTAr5EKz
WnAEIEk00tI4/rOVozmlNDZUvIgqfRarh9QE91mJ8WimNEM0qq4u8nw+cXK/FdxX
mETQ2RV92ugmqMP754bYQr0SZZECknUsTwarAQfn8eVFTfloikxeNs3oN2Nbxqjx
6jm5iws/q39tOizNdkQhPvs9aHt/R1ahl4jj5ufP1ZgkLNExjkI1nbGhWFLFcufC
mrwUbbnmGy5whxo+2KCXZ1htjKx1oRCJ/qQOuOSis5PYhJ1d0hSkGmG0T0JXkf55
/Z241koU8jnDX51rL1L9JYWl4WNYrwYlmtsPlmGE1NYLT3Mz2zoNgVL3NdAYOKsp
0lwq+SI+PB9AordAA6cYxcpHANjR/wpKRECQRPseR7j0q9hgw3OeFlOaFVFoLi3F
ip3hkoWujHE0bsYJYbr4xiuQf3Q6KRqV2/XlusBJmydkq2/kD+1AXeUG9it6/lEw
VPgCFmxr7RwnZAVcRi85iJdvsBZk6B66LRV6gRkN640K7vW6k4u4IbU8m3hVqaB4
nRf2kMavtrZMbx01XYXLLths0VgewgFNIvooQxxBWJyIdqbfCcLMPz8KCnLvVuNP
9225a4VqUCajRFvbyjAF/P9Xn9HmnKZNAtjo4tdvbeIGTt7u0gH+rlopeTQv6klJ
/FMTGsZD4GUelHm3jU1svUUH4pXQ1YZNweBL4Mr+qBbiECijdcWRlRmU+56eQYj2
3o1/JGBfHf0SK71iVnOCNIzJ+tfn99t1yppMpvVfla6QNLAvFrm814bWDXH8nZWK
V/uqdLMch/3cocJSDUBmzOJ0XtN67f0LlIKkiv0r9Iz8ZLGxjooD905PFFKLiVG2
qdoF3tEpkoxqJjwWes9NVTFwdO5ST6Qp4h2tS8RLS6wD5o0eeH3S4RhXfqgK0Zkl
Y06OOFLZ4mR5yYCbyFrs03MsxGZmeCI0/xPOh0/B5/HpXKQb4pFpfF7gCNrDxIjf
xPmRy2V8AaV51yMCbk/h8sAHEDYHsgP8Tt0FetQWETTGRU3W/ceyQFZgfBfXjlk1
015J8GQDbW6ahgSgObFz2oocOQRXbkGxq+6xLipy3XTJzMVnvcqtE3YRztpJgx8N
EXp0nWU4Jd1boHpkcaph6aNwxQtxsascrWnwwWod3txWdkuGYrRKMCvB2GuNlO33
h7vi2Znx+0Wuand4b+BSywFEF+9VrXM/JxYzpRrwkXb0Wm9cZIDx9C3XQaqYajLR
rsypOt47myCV1OHPHBRhw4h3AX9pG7+nLMd8QRZEZQaCBy9l/smUTeVtFavpxZGo
+0n0YrsT61DS2AzG9ZHrn99jAMb4kd323ztcq/IYL3UMa5pAMw4+Vrivz5aLWP2L
w6uFWtKtSXtQlkucLqJ8EBVFj9uabLULW8aRnQ7S+0WJtOE2VU/5O76uIys9BDlC
sGYaMRPGDYAG5KqEmpLQmp0xBU65RwlN/b8DN7mda3PZxmfVVRVgdHNaWIpraWLi
Zu5tRfU3vSfOXmEtoD10gk2L78sJ2JVsJ2bv084oeRm23+XJxb58wBOOqaLUsI8F
ORWWNYUWnXnPV+xbLs2220lZAXnGq/NNcbvSW2jn9goBWMOVGeFXoSgcKkAX457U
FkQdFmV6v3DWNfbqhnZaKKjsS3y87GkkV8utkZQovtf+2Hy0+ZyIjKG21UjYiJcF
ggcBpYvXW2xkYk6SFHa7scFFgHxUjyqE7G75EdH4krb//kD7QttJmP3FoDOA6BuB
bxfGOhA7MzGa0BLqu+vDHaPLLnxZbsB+JZcAmMZZD5JBOm8FAUhg3TZnwszh8RNs
Fp+y5KNFN6DiLMSzBx+MUY84/sfC4IzK7tYrW/DSz1rMCqKHSQX4Q7sgdfMLZ0He
KpQW4UfEuqLBabO38s6INivUzIB9AOm7tvfn2HnwwhSTFwQuvJ9yuEt1aOTEgubv
C+6B08RwXJst23tzNeikBuPAB1OSdpv9FbExe/5dMAKYj5694T80NafM1x13AhB9
wTbfM2dPLHixokEjURfDyRT0XLmTaXI65oRhM7HspZCE9G8ZwJaqexT5g33r/+Jb
5SWgb4nuONdNb9q+T6n9XsljDEOnAZ/QGOUx7NXvo7Jtr5NvYJUGSl21KI4e8Tyd
Fp5M2x/rXYH4HvtWwB8HdaXzwPfD4f21ZBSJ7HvNHtagjGLg4fs4Ze8sEp8/A6ve
ASZBXqjkQO5Aa7xMWQtBfEuOcR2Jd1f6dDlTiqpTwo5k1CWAeAZtlYavpAvcMVae
8SIz5h3R86PEFk5Vfrc1KI7R+O6Bm/H6U2/1W7fSDVJcD2HBUHV5vOigDgg2Ht+j
VW58US11rIi7Pgl4bWtfs81F31dzxJlIOHTfgMscY7MIt5YVu+5pBSIFumnRU9Hb
eYOd/k1Bgn7p5A8vTCs8sGnvTO0WZfBLnhRNoJ4bdnndO8ww/sSeEaaXRftgfVFf
Y8+XR3gCVmt7C9sP47NvfzD/jBh3oiqlobI6SMJnmIjJPqDTzsNRqZUINqmXDKEz
3x+3oBJXm2ZKFWmJSOSkIgoOfOzK/f6aJVFeEF5xZDAL/BrWFk0EyjH0noXGj3xP
H/JHRzlzrG+9N75bQyfCuqbaD0Y+R3Yrv9sBEabxOITBZlC2c74ZeLUkF2dGo/+W
NqKHD6AR3Zos3s1N9MD6m/h04CgYLogHM//e6rFDq0L956Ce3+lFFWQNfI/TxHF6
3wznMIztxNy8bleNPzqfnIcyg2da0rjjO1V7PpgITAen0jQp88CfQcZyRcs0Rq85
kXxmFrFWnJYtZebqw+Jm/SUl+BqkTegSVoHmF6NQnGCFrylDZnimwSzM3gZFxxoR
AU4vFXYTvz8ojGj4K3AzgtEOd2LQdJo9YaRV/X8SX90vdUtNHjhExkQAuxQKGHmR
JBTcqek5goyMXEpU8N6ij2FzwfOyR4RWr3Qog8UmD6k4Jcv6+67uOWXJvDhOnNTM
IR1mV+BrCI+ITI/+Y43Yp1oODVkerRCvTLd3P1oIlScZbYcuQ6lDO7vr3oTXCWDQ
wryL2n+CjBa2KhGFfW7Po0J3XKBg1/EDGSMbtptKUmb4dCbj2vsm7E/VTFwZRy5D
+C7O95IatXZdNGfh6tZq/GD5FFzcnOaAfr0aYvEI2SLAcwwNl0a7g3f6b98/LSZu
CTIXaWAZMA92yQ/UX5/UU+Ucd8CSTfowQi5eU3sKaOfjlIbC13T9fE38z7cb4Lx0
fm8hQZjKMPMUBz054+Aj8yHmDhIeDCzK/3SsR30Bk5K8aD4gxyLcRuM0LtmmkIdL
PvzxId9TAAuQR67mZ37HDirWHhMK+WhKUHJqF174ZQMAC9mc2oVOouCkU+CQlWWv
tJAhpB0XdXO4j8kM/pWh/yJU/A2xAPoaN4SDB31jzFgd/OdoLPDrMXpKpIaN3liO
QPam1qYSAxyIQ+U+02JfwJGoyfoWAIpmnAfL5lUZj2ksV+sDRa5EJlYP7Z0wkZh+
TvYF+OY94etCguI5FKneCajdnJf7/Fo4i+oWXn7RmvNZFW4Z3Tu4a4g3O8dgTE9w
VYeOajF7nug6UnSYjAm2epTgJ9c5tUxRHwBio9J19CTir8EiZz8cA+TqVbqSSmDN
Zi5xNGfX2oJLlqdfXht1C2tj6deJvhF4BsqL/nmCNSdWiKi8zm7qshrUBJiCfazi
OSAXJyjsbSe6huvL6IbVTReHCIPtY0Mseczh80zfs8UnMolSP6xfOY3QCBAJeRfv
VOtW63//V/7uKBkUYh8Tgv9y9+r7Wgxy9PN1NRDRDdmfxK/goKD66I7liGGSOh3i
zXEHZg620BIeniMB0+kYVXxH2wTQusfr6WNC/FcdFXBJnzzyejMxCufoQCzwbMuM
66VyJfJNvbc4uulfeAMUhPUwXv+GNSEfMZ5/xmowqyh25LffENzSLDB5+MBIs59w
CFkOe9wZrSmQofMQEO0jsMp+bJ6LeyfX4uL/8EIJWA7Pg+pQOcMdpA3QWHUgc2l0
+OMQMtnWOUkQMeh/M752sRuicTj5OqlULyhaoQ2jxfZnH9L6/22IbhRX0fL0j4JV
puBc2YJrQJkFyYXRkK3ONiIWedzgrozrQVbe7F5F2j47Lmx0yOf3ecAuQyzVdzO9
IzPMxcLAjgkP8o7JMAxTuGiAnjMxTUZQh021sHaN/m0WjbbO/L7EpbhMJ6Rjm8ij
bXsxv7dcRcltp/PSWmISxO5B3H5mmOb7z0H7LTyvSEouJKE2pP47Romxz5TQmf9F
+YhJSFr+a14TmjP1XwOIY+ViiFgU0bQKlyXoaQbBO+KcOsHSuBd+OKTselMkcEpX
W/NqtwDOPlfPA9Z77RK0VWN5PSyXB356vndPAH9VbAMdiUotMGU37Na6gZPvGTaW
brVBXqBCsocXWhWLThn78D9V5xB/MqIdKoYNkTpB1M0MP4+uXhLdlEnv0J3YBljs
E0njJUiU18KSU26lAPm6mwfIUZlq54LAG0/dvNakaCQqeCXtj70iyeYOaXQ/+1pe
et+IKBj0zmqoipHtgpADCrLwfCSFkbUCJI/MW64SNE4379epxHqxCUU0CfID1ZAk
exRr57y60fNVqMmY6TWGemYXRUVqhNWlxAeACGyEfdSmunhcLRdWD/8l49M+fx1j
MT9pdqsbzUuye5+Y+Ftfq+UHiVPFD5yZ2Ggj/l6lzFVGUkLlzldcW3Zz1RQNljaP
P/lKCdaWp5BfKx28pjNaUbKaUly9yzjYLKQ08E53pVzq6z2UVpm1zvnWbg4UCDCq
wYb+R7OBIVjafWeP1zgr5dIdVyTTrc0ObTP/0fat+CSCD0pXceCCvLwYAOX6BTfr
WENT0wZjakaSQeP2rgEaCx3UrvR6YBBEL9BZ7u1MUDb5XRl06BUVdvKxsDqzDn1z
xzk8+owtevqykJhgvaYfFAlIroW0ttdYTIck/Izod6w9eHjIt7rmpgmQzDrgx1UJ
t93G24mXKPAoK53DfLzL71gyDBJTRJDuwiPEHS9IwsIfBFwYAtzEFYhTr67F8sKJ
5ph/7o6oSvXZjdYEsmx+p+BFuKt1t0Rkct0UUvWrETNBlpenUxbt9FVNB49PzJ+Z
FwO7kC523c8l8pne7CllU9xwjVnQr7ObU/uGTBHEcjHqRVOZkTUcEJ+W7uDkhuEk
TaFLeXYsYNmSdmPZlP0wilIv3gsrBhFe6/xHKLGD0yQcy0HrvYnxaT/xaTWDhjnp
kuxzDHaUsBeXMKxGsN+6k2SqINzVU4U8yml5jzc9L0cTOFp6lDCrcUz5W24UVyF4
mJG03pMWn5YXNA+vTxOkY78np9DUQvQH067rG3+PzVWrKIUo7VnrBqWjmDkpUMmk
CqDrOloeOsKydaorxzzSV7qhOtzwIoBGMG/nSWCmeUKj77PhpZywlrkrT7S9cLwX
a8roTuJTPk/1qOI3FEkpzmxmRjjMBPU3MvzH8AZJ1re7KxeOYFW9PkErtz5JsJBl
kJdabcio33AjE7jliIhk7pI9APAYf94d4O6Wn8vFHHDoYMgJj/3a3qfgE5EXU+0P
5iGy8+wgenGiUF7aGJXz/YXyT0VNgga5zlZ9UJ/k7KVosYPH5pPuqQ6x37RKLGK5
HLSd8mUxbmvMQeirlNnWehWdlMROf03enxECgwuKRXGpqA9YoRNbUUh3qYOfw/aB
cSQ9AgPjy+p2UVkqHXii9xlxQDCSDXHo+yBsBnrNzabNOr3iiEIdITwoP3vBjWhm
Nj3Inm6Iz1D7Ld0BHKIRg6HV5OL43SG1xOnGxfTmNyB865NHWuX4ySwwBK/ebLjK
uqYqxFd413pMguH4HkDx2Q==
`protect END_PROTECTED
