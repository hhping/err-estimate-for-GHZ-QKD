`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fHrodhYEC0hGDhrF2wMsrwH1R5+rxYatOzU1CrrQe44+RyKeSvG6XZYkNa7Mvim1
eMklFCw58NxwhMelmwTg2gclhJOVfFSci5OeytNc5Bv/ss/6YRfI7/rZpapCPuWi
f6yvsIfkeACjVPy+MSRqaD8Zv7SWu41qZr5wkXaWqERzgeRLeVyBzfXlL1mWPHNh
9wAsqCTxZX5axOPFsMeB6Vz80VSNPahvf78sK02C5V9ThKg9ChZakCVsQhD3JUQk
MksI4Da1ix2+yDg+rHClLvJVksHtlmcPtjxaDH1gYBpJq3PaSVzvV40qsa+QSDTP
Dvb/zU4pjLflUgf33jMBiA08d42Rp2feD1u2yoLGqDDSGlhB0yt3lgQBD67DlciJ
oGZ/6i0/Gqn59sGtpjGLdm6u5ULs85OtZkc1xANfe7Z4HqQ5TylHLZAFFaYDvlye
3tDDIngiYFoB8TItruG1L/QJkJQhr7HRRxa0s1yvlNPaKEU5LdNOYePD0tpb8w2C
8NOxLZQMFVkrxLdwcsJxSv/1BxwGlmoWE5gAc3E9OaJP+mWdGTWe8KogWIw8x+PL
lr5z5bt3kY6BGML9NGQ98yUPJ+1gxeEFEBhu2+zt9sDMUT/99+Bs2JO0xI/bcLJE
LnCjnFWoMX4aCCgFvvCTaMOV41/JKnxHp6OladPy4wurFS8ptbnOacWW/OxZ/42z
nS7cd7jIP/dVo0xqmJThN3HQetfnasiuExU/BYzS0ew=
`protect END_PROTECTED
