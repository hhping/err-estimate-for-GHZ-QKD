`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kxYYBJKglFP8O4sWWCUty/hoSZxlbk/bm2v0PMhA3DyrDXObRGTgpCfgsqc2fpgq
GBHwYh05FSZfm3P9pKq1MXc71PKxyjTqL8fr05zc+deWeI+IryoXepqvoG/oX5ys
REVd+WyZ4E9bUeV5+OcOt1WGWLcqa28yU17zHxl7PPwN+76SK0XTIvHM8kR5Aw9f
OK5CaRCa/cB2jgGcxdtuRWwRFhH4YClj6JwKKWzDnEEX8640HhpusGs/tPYJxzdI
xdgKMrqtcoRmwAFGUgijM2HmwZ7AQr78RrKcROYtQ6nBNlLnMLgJ0B4Yy3WewWSR
TO4uf8ULSf99QKnIbYyeS9jBJsHeqa4H8jmnBec4DYakdBqYI6iWB2A62NXxFKLK
YswYIAaSf8g+QV4rH58oySWxYLnFhiWAnBQxK3Svv2KgCUh77TrjpjP+SOST+9aO
2tBr0MreaNhBs4RfhUdvQ4GRiLp3mWrxIMxNNEOn+TWyiQoDoeOjDYhA66EYRfcB
u5dMRKleDcuge8yPhWSa30IMDKW91vpieEF9+V18hAYysKh4FaL9oyL1Fa7/+PvD
L3xi73fRRzedKGuRYVvEQEzwA3nPg1hJQ/JGEJzyv2WRLhoJDGL3dnjk4AAVE1eW
QLcKGLlVPw4fcFNBeIGli/7OvWa3V6frRWKyuMTBvKQi0FVi1JEaMaFBN1uvj3Gk
tql9YBs9oHb8Iehmp3/HhQ3Qzy5qWwWwDXSeSpV/FRECLUzXYIiDAIsTqTiswWXm
fSifrX+MDv2EXEVDEZr2j49BojRqr/1vsqwRsBxrJt1tbx9MM54uG4f3fit6DEmy
ptoiYwkfuQzvl4c2I1yjcXwBNHN7kkrKnKWlBrbhMiQRdRB3BH0in7EERndK6lCI
`protect END_PROTECTED
