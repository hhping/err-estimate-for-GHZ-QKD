`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LY4+t76rjRrNNokINy3EiMKEwKqvxyK6ZuYx9w0lKvMGMwRUmjKanKZnztetEOC5
tt4iXq0KLWFdY1ZmVC/fg9+xgcFQfkPeQ7Kx5D+TadnBzwDrFmLfZcFPbt2Yqbjc
5NCcdvgZaEgORK1J4ojABmAVg/79FePSlpHTIicZe26A2Jnj8XwVLdgnNRFrKntt
EkcBroVwj3NrJX0e5KH/9CODQdSWIR2/2aL6lHzYgL2p40uoyC+PtiqJZum+XchH
tmo/0WYml1CZ4rWyPZ+wQwFwplsaT9O6yaUe2jwr60oX/c7vjukR0Xc2X0hy0pBj
k3OYY+GsbH9xE130FZvDZ6zhNC+xUWmbPWj1JO1PVJCIqsUzD1UQHXS2wIN3u11B
VsWZ7aNJDe++aXDKYgf6GDqlf3vjDDmg4luF99dot6bVRwcDooLEXvU1ORumk/s4
tgzn52Gz99i5AfJwUylVHQ==
`protect END_PROTECTED
