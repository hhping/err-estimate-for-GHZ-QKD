`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
knAk3R94pPlQHcERL98WOLFmcXf9ePXmeUL7DgJ0EFKIclcRyiZURhz8lEiwb20q
iZoC7SBl/5n5y6/8g6N2aXu8K0zSCalc3yqBKL0yvqntSyvSbTBbukw8YubNmq+5
b6XeA4ydXTouXF70ClZJUabXH+7y6+AAxIkXOa82Z0qtzTRrAg/Vvv4v3Nh4oH3i
qaDIBuy6+5rX65KymoYUJftW8/tvjIE2+XrJe7YuFSUwzoVjTiQ/vO7rdUDJSlVx
TsmpH2Cp7A0ZBUuHh1mPspv+95KC+Hun6T01nlu32SHrfIZyD/Zgf6aWyIxqf+g9
CLuf01DyTmYsOp1INyQZr3eYFKa3xDOsI7YmGq8Ebla+TqJplwgK01kPrkV77lwx
+G4djzabES6q5VyrEXy+UUg252mFbJTzjCb4hdyslgn1E1sqiHcT7fG6YsSyvz2k
7QyNbNYgZJ7Mx9tpPHfI9eSnnvo4cmR1RwO1AovxNqpSoG/DThu4ZoJL3K+iizxe
/eQWwHsKN2EUQR+LBl1MH55G+9d7TrfLhhGj3knw++R5EFQ+g5mMwLa6eJvNjxNf
d8yFa6YF923h/Q1+0YW8AJvtIKnsy+G8oVGG/FdidmOo1jyJz9HGULygfMFQqLSh
Qems+MY9tc1nv+EhXYGlTtLMZ84iaCTZa03qyZZ6loOGNiMwcWxzxsDJnEqr/ntg
AoVt1xCopZPE7wSFfVkxRzq5oM0/6cNtnOnS6NF4KvxI1wbhJfJa75vV3tHc4J01
rEEHxJooak4Iza9UDHNPkFzKZ6V2a2dUyvJ/ngd3NdPH8eVqgN00YnJXgETdbKJw
7u8RtpELQRAdNYAIleaqoic0DG4leW2fZ6Df0oaTx1IFkakeFWwUpXOzzoLxG+JZ
VTcSacPSptA14IocIAPGztlENW/VwK1pqfcZbEklmYSPK/XuYHdSSS9PVsK0O2rz
9WMsd6dUPQ/UYpx7gjfyHc7NCtQp+cjGN5nEHrmX4KpL1wNpZU4n4hWeDOH0PaC/
1o1wo0orm+e8sC2cqUDgCQ9x62W70mY/7hNFNefPE4M=
`protect END_PROTECTED
