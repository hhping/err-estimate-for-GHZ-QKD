`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cbq4/0a0Xxo2KCGIgB3cMdi9RBAIC/XLA1mZVJ40Bl2T+dHYxH/ne97gz+Mat3po
YKZA3i6G1M4ovTrs4ogkUn8zBo0qJoqfn7hN7N057IOk4qLaioRvpXdz/UlMTExw
S0hQ6ZJpPh93LBPyc2Pyy2BUeifKGAWH08Jr/VeTLdvBALpN5OBBPBPpUI6tNKVf
XeaoRjS6i/lPJ3/w7JXDrHvC1nZhC1S6jGH/VJA5kGaVjYgLAQXHvkThsqQQN6tm
rrgHN3XOTx6LUBlofqk7py5MX/pjS/rfesYj/B26l987jmGMiY7cKNfedeLk8PRg
m7dAyRaqYkt/NDuZz+HlQLk9RaPpjjxsdaq4b/rVYRY8UbkAv++KZjoLaQpu8Da3
JwneWqRIOcSTGkdXU8sPtsVYgeMw2ao2sPwVpEVnvp1BB41YMrwa4Cj/HERFIXG0
lgfB6+s4Jf01aDn8lrIOExvqcOFqNZJG6eufsIwwBI55/BoKPy6ptEEtXySTLO3U
tW89KVCIIivHyOvW5FAtugxD4iCylyysaBA33Qf7iMl1y1xPhQET++mOsWwmlmY/
`protect END_PROTECTED
