`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nDuWVYcMNw4bCK8GKqVGoWiCUUz7SqPv2bGcwpEfnSBwDa3gsFiTCFaBmVP5YnM4
iB6xZ1rOyvXSkhhuD/h4ze1dBBOmWTkrRD4/aQk0CnY0Orem6tEGf67SLq+8VUvv
0zOPVn2o1cLJhDhZp+ULgAmyC98fNlc4N7YVdy3jlixKq46jBTtEjzLw7QLIPHSW
tyGCEykyyur8OZECr774Ck0eHNRj7cpRFKv8jHrkPYEoo7kYJG9CcG9fPSYrPpe4
KVQbpQvp7WP5ISNDzh8rJwhf28hdadwMQlDSZ+IIoQMjJ4bI1JjRrODtbkdy56IN
cKgjPz8xOrnoae0Zr3j2bOWkXHpxtQWx9bIRWgJjpQjgXq+GZX7cH+jK0PeIcYV2
+cGaPklqyG7lMj13AJurUfkjcp2BIq7bV7ORqknDuKKWaV9CLjk2FiM34RVlliDW
4o4UsgMw/4Ij7q1vBegSd/BNqxXktqSeHo6zV7fxfsnxCInPE6pwIL+yDPYC5Z0q
jk454tnV6HqbHS8Q9YbGLMcigiSuCGcrtmmMdlIzGZaI+Cwz/mLPrGHqPP6oW1Fm
Np7thKiTbhRoRdhK9/rgs7DAvrkozpN7qadxYppg/PKw7fwxsuUFaQjRmLAipRgi
VS+SXFhs5IIemeB3FmiDqfceKlVJSFYXmK+JhSfftzi7oeG0JUb+RuAVCY1Ci14u
NQULUNN/vh0zuT81bAzVKS65FEclQA9D1MZ2QCFxi874ozaf0iTzQBISUgTWfTaL
zxkjAJhpxuSxKA76DRylZnh7AQFAiSzfxvSaMixImpQnvJ+5gn/cx+LiO02X2hIM
jPYBQLMlK48P70g6yqy37ND4KlG4kMxB3UFX4+Bs23+xDtOYRtZnLEVy31K734Fy
pVXjRuuUHAp9H7C1xK8y9qZIpXFNhwF0TXWjfgig5VEUCn6MWI+pa/VH+Q0vA3+r
w7VPxRgtftI6dcEgDXciUU9WSajfbTyuhrZfdZnYocDF/5+OtkNJRIuUFr4yYz0r
vJQl3yNDcesA8ypEX7J0jpmtX6OL/g91nscDOLmMr96DRUa+DL2sA3sL2N2RYUV7
lMcg2FDuDx5C+539SX5TsQLGlp12X9DZUw3UM6nzD5uzqqGKQ+iNZjJW7fcHondW
rpt/08HGV8XDsF+O8MexT7goE1U0gA3uVRF2kCerhLTIDkI3o7+XVPJREPLGtKk8
+TCSs8PgmIpUvomC2VTK8s+QGH98zZZC8wQYqIic8Je5gnKnrfk1yaeb2HItvVSf
pTqf478yFJPA0b98VcvrFA4iWIH0IF6aflJt0v6o7NsrPBcmrrQonEeIpp+1JM1x
EoEEX8EtvWUfcORn8iUkxUtFUh+fitz0uDwyqp0u5pe/vTPSoVQfW4n8FutiZUZV
32nULekV4I+5/tXemYBRJoLE6lZRQTHeOgnSu6fAudrY48Pf/LDat0Qdgj47GOy0
xBT8Adfjmr3opCfcVpVcpc5SuMtzdnTr7uNrMIcURQuxxZk4STruSZqe5Z6LFucz
xhczE+C16Y2P6Nqf8pBdIkcViSXLLiNKsqvt8w0xz89SgkZAVRmCaf/ohv4rIJIC
MGs0WCR6Od5yscWv7TSZH84ZddeYrkAEzym7cqF8912h2L1sPGCDtHigAC/uHsbd
REE2la7TItn9n1qiCbaIFI8PNtrx4RmSXjV7ohjaPg3IavVUrfNIs3OZoOkUjuCq
pUp/lUpCTgwmXKLWxTi86N51jxu4S6QkjORka8WRMYvz58dsB4UErjKf/V3K9GXC
4QdNJx027pWLPemr8rqjbibRcTyXIU6XxlIc72oyWNK5b+HqFkztub69K47P+8oN
bSCL2tC53uUBvEmBNzG98gzNSwvNYvYCmHrwoMGCB4UQuS3trYubFNpcPS02h+jm
wa0AD9u02RckE69D4f9CfMyINilnjw5Jsn+LGLZvJqwDhf7fBJeS6xAFbxn5wStQ
hrPS2yJ7RlNzn2Ye0vRdUcDU+JTJ1kgAzqII+7Zlu+i47oMcB3STtblugG4ZIJgA
KimnLR9bnogxJLnLyhc4iNzo0icLxTrEzFY4CYBmwMK/uTCR8+Lz9UNBOPs5r9SF
f8EK3tBXILc1kpODuvB5UUZF/wdT2rFPn6OJPdtOUmuDw+K/nQurXyHy1mOpKLbA
Yed5ZMfhWx2Lxt9zd9BNPowpKpWW5M2rJLMYGvt0l4y/olkgEEh4qNFRx5hKMQxK
+jule5V2tpOh3mOJ8GHAqEXM74hureUDkcZ5TH0sfyGygC3OI66F0vxeC8SvkdXN
h0YDboVg3X1DbHU78ihxx4dcCrrroaHYcvdjLDbDujl2c2ccsteM3QuJcxG6e7+L
pAgP1evoWQ6eNZfY2TE1thsCDBErwmA1W31EH8MpAXowgivoNCOwDkzBnZs+e3r3
9vphrupHXROOOFWmIJHCKCUv+t/1sFf7+T6Nuw46k9NeaWoWgK2VvfoYk9Gw714f
Z0ChlRUGh32AQ+IxD9SigLr6JGsKI1NHEDXq43TJT0ICKaolpLFVHhv+QXmZ8tDf
SZHPDN5emtHr6T175wOWC6YvQ6PV4sLpTc/aDz84NRDmkGtirMmTU3+nn4PhOJzC
Mqg4qC5ZIX0JLeJR1cQUZYT6l04pDXu8RQyZHGTaIaDCHr2M5QMB0d6nfI5pf1mT
8DYL/ruEthaVrTtvciPZ2CrwSCkWDctSl2PMtsvu/+kNyVoQdO7By1WUtkPLc6+7
wMI6yV7HoUzV6JF9Y+uD3gQYMhEPXX6pMyLjJydc1cefYT1tY4u7i5khM2XtzY3A
uI1W8Rf5Ls4ZzYX1iD2//vRZ3uHN/OQQJzzzW9K5IZSMt9FoMWKaORDwdJNtjrRk
SFkAZOPsTLlXbMmqnc1c599Fwbp3mt/Q4/VgNkR4HDg4gq/HQGaPLzicmsRtH6zs
Lc36EifAvyc3PiZjo79ECQMdSQHoYNyJMrdrGJEK5s2EXDpnMZX4t1sfdVu5yArU
KOfgEGBwV5zHG+lITiuU2TH12f5Wlpdfw6mMK5XEDR3TH1p+hUYqbB4MDDWvbbrS
TAEvPZ0rMKI9gq6lN9UGVFpIUzQYx2hoi4pNMfMuwFYV/IFWvbHNIPTBI1fA5jfG
2bH3ZHS216k83+mPOtjsMHmW39CZXqrQy/E2AkDuYQc9XEC7TNpkq7C8Jps/0mgP
VUbVgT+YsLWlCRe428Li2D+AgaFfSWlgnSIBEsr+RpwicPlgSkJIWhhigqJeCWEJ
urO9ewvHQjs5VGQdRqbRyzkevOLbvClD/aEPdD3yH5S038tGmWftfU2mFRZWQYpO
wxRrIUvk4C9LHpokr8dtlYN9ZJ4aMuBY0Rb2ouoj7u8=
`protect END_PROTECTED
