`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xmHrd6ogqC/o2MpvruUIjkhPFOh2Tefrv/XViILANmLc5ee1ZWCAMd3r6OIh5Bdc
ljqWE4jjT+xpdcDlUyYRP3JLlZCXVPuxCYtDWBeXmgw9JqA7vMhbMeI/IS5/vujn
QoGXO08XXye/2BLY1kfBP2mEgIAWRL3c91JD22LdI+YDgLIvjD7hhnTFk/XZ4udx
eFH/Qe6QQ81cUl4hdocFaBOkQnLf60ysP1VXWEDqxxYA9Ori1wY02LcqT6toNbDd
gWM1anwq3XKD5uwoMwC2D/4xGIpqOZwAJ+MFbMiqzZw77y9WYyi62dWM61Ad7xfQ
Shtd9gEBaiF9696MWgNCXZoDtkywPxsnY5qPWvXn5yBmKJxyZCuaC4FW73PQRCyn
wFZIpXc57TaJCuOl1xu8GhleLq6ZqNoPothFYi3HDH0dSekJRetbRMxZbytDEaqW
/bbD7gbp8Y0JLf3ezsVu6nT5HakUEOSrLrhvFsqiIOzVcMUjLwA/8l3GL8BgoHv1
LoMTI1LJxvy9E+r4dz86FlBNRT87PeiXlyBh08D8BBWhRSX1J9GLRwdpB0Y6Rb2u
Z7Dg5o4Jq2haR8aZILphT0ZEMLnXumMtgF7qTQCS4ZLLc0CVib+QD5N9n15Gn94t
xQZFsSuiiS8Ygg4cKx0TnfuslyMFsZVh4pvTrO1hYya28yTV9lsLwq98QRlLTbMF
6m9RLfWUFbPz6IRPHp1zulT1JlxqMhzYdz1KMT6OIVnXlVaNn6x1bDTsz4p0kMbd
8hwPGe/WbBc5+zj1Mb8PrVoOy9qGhGVmZyAwoPfzKeF9XV9PbrdQBOwqSoLmdRci
QeIpn7Q7Uk+05OX2Mv8Qj0oaFzptCspKnu8gzA1rwUKMZOOp5bgAdrl2TstCowzx
ty7B3rJpKqayKGkdCylPFNjedFofkEMurKGHjxvKsSLuQ7ghH6i9Yxo67XL/2tVA
ssWibIudOxeWtv2FKzJifGGBDhYRcIMDKIsuiA8mXLQqo17WtB465Rp465f7tP2A
0r+qeYVEUM05W8pNsa/N6I642IxbnBY7pE3XOkER/xYKNLfKL5De0EH//aKpeEPn
zYOzgAJboPiUfSqTp8hP3YyE6ypI4KP73kmW5srF72wWtDmsm+0m1r/RTdNm9ss8
Vl9bYLKnaMe/KxxCMVv4E3HOBMQr9gh3E7/jvrIKwyGHCZa0OSIu7gy2fAy7r+8J
zIgSq6I3su5NIF2VKToXS4i08xLN2g8Wr4pB6ULqDqsHOX7Vz2fm3z9xDCKR1IfV
PchMfPY1PrSXPwsxiXrJB4GvQZ2C+sxSPjnXkAnu4SCA8h6DAer+EKpckQqxw4lM
eOinsMecp8VF18r4qtZwE2LHiZLAd3v1kDlVadpBJpXC8A+R+HhxLJh5TIYSGyzV
qzKy/cSSuFo/xE5bzJaosp8SRntZiwPH940DnXC9vh2ICOZdDtXwHs8r62B7e2k0
YQWFZkF7g4nOvpNguiuen6K4vWSbDtRyYEBHGzl5ZIisP2wi8hIB0pg88oGhsn8g
HSXjN947MSlkS5avIZsoEB1LZys3KrzEgCoi28WQP7eO//7tm2TrVO7SQIQOrRDm
JmDLFLp5UFr4DjadQZinZ3xP/4dcpbbPd8DB8dw2CVrh/FJHhat3bxxutJrgixll
r+BPHVL6tpG5/O4unLZqeBPqg2luEo5TV+FlvoIqdit6FceRcmaWfUhj4UktoXYs
1B0SBJzrKAtaXoceQdUWELZD5FROJ6ZLv2af2iO1iETgP+ldYoslBVfYsYiNdhXa
XYbiVA18OHak7HpoIIxVC1JtEKYFEAbepidIvFqpcblURnywDcRNAeOBkdH/oDN9
wMNizuXMnJqlfnMfCgNHUlI4L6U/nRCIjcVEgO/IWNp1RSSLIXcHesIAA2LowbDr
7l4nnZqBVA7yeulCauu1xHTyT7lyeRFVmItcSq7s8CGNlQbhFlcEOjimiDCWJVZ1
poxXQx7UhA759G4xkG1iweMlI58qRAFOoACcfit25Srh1v6Jkk0kzS59T/342+Ga
v4vFTCIgwXS/2sTOhu44P36aEhJHVagE7LS2E2ff+c4R/zRkxN4tFaxkrIC/F052
32bCQOL1AKJC8Lq7HFX5fuMi62hmhDCHV/pxCQS77Jo83sehzhfZ/gFefZY2vgiX
ommV3xtbIIfJXujv/nQLFEdGMtnsi9bYKmvBZ7QecEJ4HUXFHgKgwbxZR+QsLiV1
d4EPXsXq4JQMKoROIWRlvYYklrQoE1MQ5efrDU316zH82U1tD4lTkGA/5KdkGeEg
I1a5h4nehjh9N6YWNUIFNgfYXKBZqxhhoj/6MOhrszd4SQ5feKYm8bvrnPl3r5PF
rJuPMV1IdJ4l9dotlW3lES85fDOLmvAezT82jaj4GK1RJPfWrYlJaWFdr7BNaLYG
1VLccNKsf+f8+/lnnEKM396mli6qF3U4lOqZdVyCFUnsTE24yRydBb2d1tZ0QAKf
nSqd4B6RrNRmSaB8gcyM5YLKroZGlxd6/zWQRUe8gIbQa00JcB3+VEmmMusZkTM1
AIggAXF+1CCTJThdnWfqqQAjIEPgwBYtO9kWef1/Am2bFcVcNt7AvaqZ+GvXkwHE
F+M6qpIU2/SszhzGSk6mZ/8PJ0dl8lLKF7l+TpMpI6Cz1gf6CaiznnvR0obkB0k+
G/K791dOvyC5N6a7mTb6/SK8LlD4sHyedNHEakzKRpEeUFdKawX2Rnx42TzpDlZg
xsnajGYtir7WfWCwNhXhqk5mmlyNWCRgmAZSjfOHYZ8LeZ0xkpMYtl4/0vRUtXTy
HiQet9TqhvB19Vsa/JbbQgIIR/YindqwwWwF5tYBzIjgXRox6RvV+vecyIDZghLD
jbS+R+JC/FGBARmqSxR70YIMySx9xjB4PvKHrlxRjpNK1ASjvTBPWEWtrce0sshQ
6t1aoLzlqy/N+RJaunmGPjj/FHOJLZ0UFx6AMRLVEnf+6Nq10Qd1T24Mm8J0H8jb
5T9Tm3hX1XOo0u3d67x+yenSvMh9c3r+iW1foddp05CRdOYAmM4alnXHMsNDFZd3
BMx9djmfXklkCfLrp4Zd5APkCUjLg7/yedYYAOxOF2jFvo1B0FvVJnKmT1eGwwE5
D0IvOjOTFv6E/DTZiW5ILYujEUVDmaPvtz4NvJlLVvPODAgxEloWnA8Ub4tToEfR
heE189/HJRyrN3u7Vcy1FTM6AnrIHMhGT/k+S1axR62yrNUV3ubYAj5hxz0nBekk
mSWgwC7Ak+rqUO+CMTSquDzURGD9pU9EyY5WVQQxkP5ZPxjSX9EO6+O59poFlwvw
4C+qsA4DbrKBoX83vYC3fWh3vK8OIsqILT9MQRAFMPUjKXel4TJSkDZdIrXu6026
VH9zt6TSSpTWsrzvABC4VzT4OEz/RrAPbG5JHjBoE1cvyBNWmblp1PqkvcknrAd2
cwwgW1NqxENEwhe9+zigCHGSuju5Totcvu3pYg4MXxIfGTnxJbleB16wkhjK933/
jyZyyZ6QqlXPjh5RWnQSjL8we6m30BIpP5ILothVJSXZT0XY/MTTepYDw5uoM+/W
2wA695n4pBBS1sLFgGB7LwVvB09Wrm0uaGGJvTdbuo/QFHfL9ChBeBKQS0lhMorl
mC9n7fSjo9UKiLQXlTLHr7pNx44SWcu0quNRnbHnFvG31OwQiYLysZhSD25f62YH
ckXpWtpC4xvxXUolqXDv8N1qvOb2Sr8zCajOrRaL7w39Q7oY20SxIbyuRd7gCQIY
`protect END_PROTECTED
