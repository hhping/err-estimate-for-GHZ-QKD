`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KmrxRE+UTVWT4U4M4paeJRombrbOjBFoOroD0tPWsHL0PiK71AC9auoelAzi8Wh6
QWZhrEDGbHCC13jqxaiPWdGHRXnjsyZuu20sG8U/CeMZvr+Tf1uvPl34a3E59rLw
2lh45E1F3zP8OPMmY9iZr6orgkiYo1to5yoGkYQVRygKVYu5VcaPEglphccJo6/q
REICxz24KstRa2e+yMZg4pnUhugxR4bZPM/1cpR2wHeuUyyaABPB3Zm8GANZDsjU
Yms1Ipm+h2gTwOGF4azZhHmUEGlialNRjxAi9DcV7IpxTf6RVrUfeCvUag2Qr9+E
jtAEN6NpkAF8ZNSTovdAFVvlMdElSSEI9ett8RWQEkSY+gZ/EuHqYmd1Sm9XlNnR
PlcNBwPJzvXb1COibScwpHOzJxB6KoEyN2PazQPY92MOdETq/CoTvNYDhG2bleBl
3ZYt7wdJlc8Om0ne78S8l1tjQwwXVaxxZDvWGyXCjHA0KJ+UgLp2uzjEHD3YFCbt
/mOU1jaPuYMuU0QYG09Ci5OPA334Kg4HV84K5w9pidaErYeR12mXZSKXX/ZXY9ys
WfjWvvkTjGaBYA7r7t2c+8AxI/B2Uj/tFdA4jU6oaG+mkn4yLwwgfR6f5cnotJ8T
X5AWPsKHxkkYGe4OtYpumwY8GzN0oTa09ghY/bBLN/0t2AHGpLxceLb4pMmdgui6
PJk0plUTN+DeiJP5+As7QJtl2OUOSVLHjksgK6PD9EMNcHxG/AkEeE1Q7t0eTTNh
glTD8sM865lK3ZAVjBIFlEEoGwU7Wue6eE9bfHdOovOHZ/aPTM9PO1740M+DKWyV
uzBks1reBezqVg3nV/DPL3opzqdL89qkI5+7hYZv97OckYnuz8pHBrOf/YRFQDG0
ONak2p9qaWhT9Jgi7jdzGdiqM5zhdzm9HPTu1PKRNHgILWi5Oo8OEgldMa1/Ny1e
5lgxA1b4j1lhYln6Qi0d8qphMJA0Gq2B3cflNGFawNv0TFiAPxEM0cEACenVgmJS
TZ0nUGymqIt/gCnSHfcYXg==
`protect END_PROTECTED
