`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ei2jWWOzc3Dp4LF5Pii/4+PfCxL/SIZ/7ixCir8a9WVb4DgBdm60tw+sdtp1wf9w
YquiRnsx/jMlQ6gs3SMyeP41r/32ubJCk0EuoULlP/SftUi2kxGgUn838Mju510F
UTcOfwRhfB/oPVyreZ2J4fRKYubDgHtqe9ByQgNVfW6p+8FcyQ55enTCupfL2+1y
8ZyiJpXnbm64dVdKhsjzZeTdrhLLSQRYEEUndO5jtKWAh61vBxDB/lKuISTdXNHG
WRHGMQI4vVl/i/MsTSWEDuD4yLr00+bd5uXoAt/OBgsY3qKJa6H/N2oF+mOWEph+
t4abKbwbB5U27tDNseBBzwHju12E+vrJChcR0C+88rsJgLcA3Bx8HvzSgvi/bekL
tG0nHaZopJUiiS3NpAXOsfF/coPpKtqJUZ5zf3PCTN6pIEliPYRSNeznvPf/GsmA
7+yTVqOn7D3rrZfVFT8raxZIJxS/L3+LVRyk5FhHEMwSDfX9pauawskjf54wGXzK
V/59lnKOJOfqgCuZ4uCDawJVOfTNLzouJO+mbZ9LIZFYoYXXiY4lRjqdYVuAVp7g
Z7xq8xMsTzNpWLINJxU4ZsXYGMg4tp0MMAHbEtluyBsAE+mjON1nVk31lYELoMFf
wd3hsMSAHPt8ssqM7GOtPJCJQQHnarJARw2AntXKxDnpRhizVIK+QKmhVjaTj9zI
CQ9OFOWV10/U5JjzDx24xDJLPgjBj+XMJyL000w8W4OYR3+6I3js0xbANCB+hiip
2HKNnjbaL6t/MU3MUtk5KN+Y2Z+Np0PVWL1yF6MVz0Jqu9WcsqZFN5OIqt1rswbm
4codjO2sdk9zcu0JfGL8pU3/eZDvMxwhL1MTR+gG5xTkGD8mujbXmLBT58XkFomX
HeR+AR9l80CaXek/IaNLHmFLy4EpNJljVpqEC09zZ0JEvohBS+yJ6PMOvQnXyMgj
M90uBHrl26RB1Pp6AjVrBwBjLToJymD3iok8QB1AZE2WrQ3YrchjQ/cGu9vsotaC
RpA4MlokNfKgSemBU7wUOtsz49AvY8ZgOsUwdSM3HbXupLShcYFUAb7FQJxUGu1B
EUgO2TDVaPvGLinOXTUB+AelWXFc6res+h/OEpjj7STwtvqUvAjRkv8LrjjBlV+S
9rlDdQzymzQNN37GjDTK6dvcXPjUXuxXkpo6pw7r9QRkld5Bq0rhzPFksMws82mh
xcnc1lqyvXUdA4z1CvbecLnTACgLWHCXfeTkGm0H5dOU0MstaoQnbrvKsPTLj87h
2c36yUPWneH24zGgeH3/1XupRz7DoW665ThOHaRl/fKZiH6pRupxSTs0kwqq3luC
k9mB+qng/QTl0xQn2JN2d9PIQ14MGWk23xakYxrUZEPfY2+z+7lgx936kNIcNxRO
IbLggSV3FjwTosFcCv2Cxb26R20/1FkybxSJMNJ80MF5I/xdbznWjerK/mmZDehl
SafezurSc4VbwCSQz7w7nQJa9NnA+SDcnRPaMRZSrRdE4/8TJpei+VIeRgUNpmmk
g1h94ufvmPtZ7KKD7Lpp/rTg0lq+/0ESVQTSchhwyjuLxwTGFEmccKWIgrXv1RK4
SVMuUa/P8RQr3x2oisYg7eC3h501XUGDi6Han9cPlrO0uxwv4koyYX3aTvhCCouu
OyXM39S5cnk0xJi6CebSUd9v1VkGYfinpK5fC8NeqnU6/MA8SqpUg2PwMpwHWgk8
QZRfCOwIgPUDglZefamYi578oy4urRZGNHV6Cy/jkWUbXu8OAyk+bS7mxesAjiJk
mbx4Xl3pA4HcNnoVgpmqk5sDymonb8gkzeVa1QzCWDFPKxzP1qqSqJs7My8BZXw2
Ou/bgPM2ZA0mTzX6yk7N7wJY//W97bV8zoo3tXBro4BuIm7fRXtGPh2ELQEvlR9v
INjkX+E3tyzH9NJc5ozx7xkLrHb2YBlz280xw6d09Su51G23Hhd3t0ODr/m2+nkp
VSNqqnhg6r0No0Nv+9GXUQk/lFqN91f4AWqF0mrLqGggI7//GFyGJV1xJLWeTNje
vq9baiR1emzgDz7hb05zie0LBjvj6hqYGyTzG4LvkKiLEt2bMXbUX3fMMVXaa7ry
FnmEhjFcORXSYFUH/cCYwjAlLddEZILYIX4ChvI7DSqMH9qQzVvUXjOvyVgiH9lf
dkEw4/mpqlpfvhtr3862UtFB4IXb6ed/JkAskuQpvN2lPmbVFYjKc/pVVcnfVanC
3xVxxrZaKIl1HmddbyfuZn8ib7PzutacdmIXVjJnbsNWXAYkRmCkwMwUR+XcECsJ
Po4333b6rbLLSB9wXqfGlxIEPVC7frFdc1dzeSNz67Vnhzco9VVaYE7NvXBxZUzM
Gp36X12Za8Hjm7GDmXRUwYI4dEG1IZBwoPwccBHz6pTu3kEFDNKfa33455Kh8k+f
ps2o8va6UK+7zHZrZV8VOlE5J75zTpF+UBWujSKfR1xRrFTGzAAMycXKzSGhb2as
jvfot/dhT0PSgD4lu7Tufp2kw8KJuEc8NvmGzrDpXTQ=
`protect END_PROTECTED
