`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hm8SRoBisc/ssBZiDm7YhrmKDEGkn3Glhc+Zin6ZSrA9mzFXteqM0huNZKuSHMRb
oBcd0eKHOVlHbBbjz6TyLN4PEkmbYW6BD/jip/1Ow8WAXTYIfPI9Yo8CutV6v07d
g3wh9NQz9xR8ajyZuRAuOMor2J+PYMZXyFvy8P+hj9t3Z2L6uNheR256u/C9hBqM
6qam7LqgQIPDHnHNbuzhoeifLKyvtOV0dVNjsZOcsjGXHOzrSM7/5U6aZktErJ31
2dvIhiElmU1zvI/AFvvmzYtCGsiaTLU9v6XcpDFnjBScA7XwHrTmF8H3dif6tndd
9D5pRMNkiXCsu8uV8Z7SdwEiMFMPDZ+KtKxSey5JV2xR7Ja1cKBd1J1uCSdnyyIp
SFI/LVTpZm8E5blEHkABloEg/FJjuQrdCb8aSk69zzjLEMQQMFuUlUpa0nMI6ztb
7PTjZWr5hPalbXBmGaS0kwKoM8e0a1VFBX16HECJ+R+LxGsZq/6a9iw22ZjhTZfJ
`protect END_PROTECTED
