`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hgsqahNNY2zCvUEYO6sogaw0sE8QkrYxoTXb1tnVihD8bbw+qo4LNGq07vQ066jq
L8Ut+AiYDaQOIBOD3Q+xRMi0hax0I6H7O+fdp180DCTFtqvniVBFN/yGXuma5Ylp
KWTv5Efyy4TcXie63Q7OUY+dAb1+vl518eyAQiT8YWJLOmZnfaFB3i6RAQfKUfQ9
7FFjRTO3tIl4yxJdUJ3UxhZG7G6LQTzEKgKhSsbdQPXyss63D+ORr7IaZ1jM6mbi
jzaTbfm8Tpkr9vB6jODCS4GpnF05+tVgVRhUOn/0+PWj+5U/KLGy1pZEFMsYBeJ5
7dYiJsqBQfS0GxWhLcEKV9J03ETkj1hunpyXNHYeV/pLi+kCMWCqkgeITumAMAys
c9evvGpCTmcMXvnvCZ880xZM7uGu36nfN47ymWcGiHUNeybvoCrDTyp7lRmaMqK3
YrjQHBqJAJP9pcW6d+Fgq4XBPoWpliO8DftjFJ6IqZhI+nDV7SWShJC4Kbt/h6gS
kPms3nd/TQsBm56ZR2FptmduQeo2YAgz+SwZPGLhv6AaNj7tPvWWYnpZp78RNLyU
QiGP4a9b60ZFji/6BZTAJg4LszmMOf0WvS6G48RPqufBt/ccgy7ghOo5MjvtwXeA
d1DnJULkI1FXDwraf7K45FbppzxoCoX4diW1eZdF4W8CKgGAiP8CGFgtb95shiHZ
9a9ORkNpzB9J109oMrU9vJ3MHYi/ZpsTvFlYN42Z1AY=
`protect END_PROTECTED
