`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X87AtYdH1IGiep+mkPieOoYTp/7OqqhFAohnnLEVW+6vmiYKrTOU4vJ/ZTIHwv02
TNtwKMtY3z2+7nySFNoaDrh5j+r4RUhv2oeQu3sNgvslI0z+ZsVEGWbruSVCgDY7
Nv4WUqEGKCOGajonwi5ts5/RKTXqIy2/q1zpqRo0N+qIZJVDLfsWR7FpnEPjeQrO
eJnykMg84HVwNM3MkQBRo7Ksom/aa3qyrJNySNMkR7CBA4N2949jFFic6by7iV6n
o6rNt+X5c/2XYeevxGe/7Zo+Rnc+ZQslDUOqb2BZeKHvSlLdqSHKBOE/rUH2yZFH
QvQIqO4F/NU0QA0rHFFczNjOxc7IK+GthkBktEQejt/71pqBwIfHHOT5v73qr7UH
x3faPJ8T4D+j4ogRKGEjsin4WiZCTfrCnYLBho799hl4iEcCErCKlMXER85ZStv8
RvDFI3uf+oIuycooe1hkPhCTsenBKKmbmxWV/gWdqRLhVGAS+23NHMIvzHW9vCtq
kWXztBj2sp4AZOKI+gJZTbCukGT8D90y6s0vhP5E+AJ4+1zFcbs7wbzDyA0w0LCc
2cjBEgoLXNMhK11uhW6QWNNIWUqsLAHf5a5bVBn7+pcFEHCiBHwlrPsvBq8HBb3a
nqtJmj+qWWHZkhnMFOHyoPy6dNU6JTOPhYFPgWqgGue2CP1awpD+WsasEZCrfU0V
s7+RIX0O3Lifv6izXceaAY1DSGMQh8vC4u0Zq7/73vaswDlYmoiuj+pRzs7n2Qg2
H758H0ayyihpWLzzTzqZc/9P+WqP0cYIgM4b+W4Z/LGy2LrS6QWF2EPkDC2nX9db
SXer5HQhsQi7oTGVqIaDbPBAHqUCYCh+21T95iSvR12CUf0kZFko0HM6sZ/w6J+s
ejyXKIp+GjStLy+UgfaP+evW2Lg5ZwiwXXhw8dZKg2s0was6a9SX4oJLe8yAgmMR
pfDNH13jHO2WSSUf++FEcxemjKXH5AwJry8PzjcWyVat+X9DbsP0iPrgm6cNeJT1
/dyihHpiJJCMPuFgpalBdEqT+AQozyoBhnW7c3C14nf1yBqn4bsmA4hn9Fp4NW5e
DBakyESaJY+SgnMQT/gn4g6tYXQck/H3tvTX+4uf57YpecxglI6Km/AxI4wcs9wu
su1chO1/rOjBUT3TOz0sa20KjAphIxba9iFCU9162uzzRQbTpoNkCO5KmpuC9XOw
pP9opxGLlGbcWTgbC+zh61WxwfOdUqi2MyKNx3yJHHRXEImdTGqHoLcFB3Z0zb5J
gytH7iUJ7CKrxIA20PrwNXu6tCzK6ibIKROLk8ATWJMUBxvgWgBhKLfofJNpT8+T
nc5+lpEDAD1ZMAqvY7h0404b1dsvSVGAEVz5VOIb/i7JImnCu5Yxb0Xf67Mi0gyy
0SHPtw6zmcX6WHUhu1FyorMnYr0EsXyz+uPL+wcU0ar0CkBJpoU6uGYCbEiSZKI6
/MOeoHk4wPyEVLpjU0BqmZ3EWi7hepFEozBfJ9ftMKw181ZX5z8GqGqgmj0qBgUD
UbylNLiCPklUk3t+zgDmuiaK9LY1Rhv93Gd0lrxIvXz707x/9KSiuTfyQoX+v9Qp
cpYsfJyxX2BgFQdCbMMYZPZ8wsJSVACVKu/0RbcQ39qXvmXE9/h4vZwUjT921unt
M/Khw2Uk+U3ssey4RyXG7zs7gk0myhMSNE/pF+feSVsYauWhDOcoiFDx2QDJ9+DI
+nAVzKw2ZEGEO94gsQGaVCyWbSLr3xwb9K455JiH942efzYiaJQQyURJUqx4Ls3o
bW2fO8vnh3wMUGWwcK6D/YjuMp6EDXGFEoBZ3nwnE3Vl1KNRuGSR9AVDV0zEKY3P
TIUw3/y/EmDrwky/a2ij4MO3miRP23sBlbeRLvH+95RcPCIYqxoapOPL4ph3LYSw
vogTsLPhWzTErxC9mZXCIcYjoKg7c8eUHXLLQlyLrN16mgQ+14AQUSB3rmYjZb1J
Mw/PkxZxdW0/2nU2wn+swbR/M5uf9W19/oGDHEEU1tiASI208yR6RTF4szfCB+9Q
ntkj9GrB3OYaEhwqC4/QkNKP4L8bJVtjsCKiDuSUiGzTgulAQsIjkOfb5BKxMn1L
2Y1bD0s1inZKkvddyjLY0qolu4uaKHrCxj8TdKEe2DnweIkoF/uOLRyoYh/Pf8GA
48rSGOXk5o3McHHRvEyX6wVbfGNMcXKnTQhDZn5QpVRZVUnBfjT4YK1SSH2G4BpI
VaMReZLi5kK46UukWKn4LSdxFijuysxHvp+MOrGWsebB/kT5AWrCGysNQx3K1Tz/
H10JQK2hsKJgZ0aqhwn4AXsoleXPQNAzE1s7NuGb9v3dir2sr9jE/ineWQFd/wVI
A0xsOVJ4DI5BQL6Zcx2f4aU6h6hrpa9nicisDhirwfCcXW0YhvqsYDrQhxHXUn45
u/VYc2IVe5nj98eHMYQo4vOLd1Zhjfdtm0NUWhW+YRyiwkdmIek9+UMhXubQacvx
Y3EIQ5WzpOUieDRcuSw+hA+gs/me4oI4krTrQ1XvINnTu/Wap9WSpm1RDFfqL/gm
6ryLFCGlcnO0USNKxKMiYOOAWkOySTLUgHd9GDzhcjLVCaF9lzPpRY9ugOoNuIDl
p+Fwrw2wE2LGOrhYZsJfnG6YMGld9T3mWUOx5D6Qaj+xYc57brEx8Y8NkmmmmXYp
Tp1pNjepKmo2x8u/AGD6sNnOsHP+/6AlnTS4sU9jaKRwQPhBxpwe8eiGIQC/vb26
RrVmUli1VZQrMEWgR4Engz5Gs3Yujgoirv/yVUlQrELgBkjlw5bL442eQGLfI9eI
OIimIBeAbmQ3KdrOUlsnTfioEOZa1gCmDXsk1DO3o9hccYSQvATbSzG3TilL5qSK
b0dLszpnA/zn3lOvFpQBVNi6w8djmkF3GTs2zg/q0+OY+e6G271z6tB4otD19k2k
zEWyt26y7hSJyAsWlchnrgL1Av4jSOJ08XhrbzedbF9yqE9G2kq8Acn2bU04IKrs
Y9rMZOaO+YFMXCh1u1OMTpAPrLZFuVlpHDJVpB05izu31iD5oN780qxmqoZ+Lnj0
kuQS0Bk7TRKEHiCmIF1On8TQbp7jRz/2abOyZgWCDI1O3Jxe/3v8LvxqRKy/qVwF
PJ+Y8Zlq6CyEUu+7ulNR750LUGEtnBprR46U7ZscfTL5M2CMmJ9ukmnR4WipeQbb
ePvz+Pm+CQqdizkXoHDBLQ==
`protect END_PROTECTED
