`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
It8ciM+1rICv7DZKQ6FXnXFioiSnqr+2QVPPuy8WPSSwKwiB/1Wp1z+wHTWj3C40
h1/N7lT8MhrI8rKoS0nd9NvVGH/g9pCBX1zxoJ6txzZkcwvkjlqeJzs63BmnSN0+
1E2aU0OKWYcvGmtm4UK7Iu8B/6vyQ5pSRD5FMVZ+AvIOeHUWQhsTeL6aNY+BZJsJ
JYKQ9hvTUrQEAX602FeQ3TIMQ63vfeQNs2EGJ5w4AyQa8sV0on5huuZ+XzO3GaG3
3VAOGMSFowW6xwcRPtVqnmTB2i3n1ri/0h8lTAmzi6fxSNZYXHn6LPXjrPyrD98P
RiOQ0ZOmR4yxOG+uccpZudMppK1rbgsi4ytalrjZlaV20IYmvvMDEVLl6s1u7thU
zvUSc5HJLLZvtENVAaYViOv4rTRM3dL1h10H0H6ZEAuB9WecipEuDyuzd2lY2Rxc
Ov5tjKc+zwZRU6P94k/jUVm0prptDvnpB1wTVRxlZfDLet1Xr0OnsNEFei4LyD1/
vcneSX5MQ0ws+bKRiqCw3+NHGKVoosrYyIAYpbBXnmGSPBcQ9ZZIoJPGMQqGOMNU
I4S+Bcv5peFksx/SIYyK5u6nkGmfySr+k0xiH8knAVhmVBQOr142phqwpAs1V0yc
7NtYTcyVNPcsFjH5/K0QIze8wJj6+HtPDGgLGTylVArbnu8IyUVk36QrZcmW1oFU
QhnMMXOnjcN/rkQ96qqTUNQukSzqM8DxGDDTU/RFUncFwMIoDtcKzwXfM/mTryi5
tqxtr5Z/Sz6NxvsZ65jiXGiCNOqRRgtJaAS3qlMiC/ekS/CneXHu/lV1kNp3OhKr
rmUBgolo2lGAPXRUvtiF56SfnBoEJTu/c35zY2fgEJmXio7TSKtcTmSy6yjZBi6E
hUdZkVbmjY/629pcHzH6hlSePwRCW7RPMhpS8qOUszpsJ9jwDma2yN0B015NKfXY
AWdUnsBN51gq/9M21VQAL5jcc9yMQibzyNRMtBQgPDY+CaEEW62b0UCWCttw5hqc
QAcUSljWooBMTupbaWxwA3F03U3vcSrsFPswbTEpRcNC44gWv4jpFmCy470HSIdg
kIFU6J4NxGJnCM72QA5srLL9zck60CmfDZDuaAarWZia/pNWrMkjxNLot/fBD+d/
8ZQ3s9hFlbMi73a5bgIl0w==
`protect END_PROTECTED
