`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ME9Gm0wa5OTINqd1cCIDBemPgJHJEHO1LowgP9Uv3TPGfNcmU1XQ8lfFU7OOoRt4
1DQbxauiJpA0razuyBSPrj4tbYJwojMPL3EW66Nt+cTzsGY8FBZ2bhdzoh4fk+xx
Kl9gCau/2NBSXSdHlLsAplIaPTHQsQwchX5/Y649HX/Hv7scHvs4lsxslNVEtWeQ
G4NFKE78lFNMcvvCpqdSrGWAIEcwijS0dhMdUZTw3nhR+or24H/d/OeyEEiEV8cP
qzxwQpWvTXV9uY8Be8kkqPdNM70o1MoyhwTtca1m/gi7ILdfTOv/vypw2zOmF/Lt
dFFWATtL/POeIDCvgFFRTF0W2K5uvXViL26xy3I1eq0ZK7HVCJyapDaK7ZMQ69KM
bp8VlWzNoCmqNLKgLnlGQH4tUZWTsAr+/bBXnKWhYTWCpB6I1Dd7UR9eJ1uJt2Le
FOODGxmsH5Op44cxAZhoJJqDsHca9peuTmepJkurK8HWv/lGQPr+zlQtR6aHEehH
+BGOYrNKM4RlZaphGjAFmukjvUccQT6sn7Zdp6NLZ/bHNYAiG1ofsnWo5X38lEN4
ob0zy09F4QmiB7as30CZTgTbD4vh7MQ1fpmZ/Hx0lDCzfC7mt2h5Ijur9K+JLr+q
jzT4TxjD9MFhcmbSzEt+7X4MY7367L353BmEmtPUogLRVvw9ZCZf+sJ4XEbJrJHo
J+apzD+QIuSpO4ttxs19nFn5NzsxVrnh53HxMfttsu6yRU9dzpqVIC/wylpVOK7/
jujm11sgW5CVdqiTbcY7JJEKymAgoTdpfoFnCaCewvY3erXcM0P01tmPGZPjgfVf
b4HuQqE5FEX+cS/B4YC5AOtA563sBx1jBzx+/i6O4roPD1YHIFyr87ln17eSZ6wH
irzbhNc2FD2rYeuFs8MbEALd+08V5PCvsP3mqMtu1G4DOi0V5BC1QycnxgozU1Yc
zYHQXxj24faHBEPPL/5Yq4Y9G7AXmtS4doksvC84GGmdbaaafDArv1UfSgDMtQd1
Sz86vr7W7FO8aCNKExSwswv7pzS8QqQyVTw88SDEqIlxXUOtgV91i0E/+slrpHpC
sXN29k+puynXmktM1wQIeQE9EV4E26FSTxBvhoE52Ox6WQN9k/Dtk6PqDFDAjFhT
8zHTUf8lGPN9yuKI2j8PraSQqXdFBMqX9ZRDPN2ANshdKMAkYSgR5IIUon7rsSYG
0JZrcRsj1GhIa3z5xH6DamWeyKYZFzXnzJUfz4guyw/UV62WUdF0U0DSMnWehd7P
2jhMJsJl0tZOzAgPVGIEzEtNIns2IXyhZyAmZYw/gy0rEoO99pJjgGo9G4SzhWQ8
TYYPm4T6Ly7SgBGC+TPlrcAt2zx59NB2xFeynkgDf2y8cnEvIRJ1nZ2NnsjGblWM
NT/lAsySO6K/HfJiSucBuATGMTXZnd41v3yU2yk8tqilB//63ivS8WyCvmnwkNT2
DGCeohWCYaz48Gfo1lDn403cDZt1zJVSkr+emO6lZxebemDB7Hg/6cQV3fWZ+SNU
1CnLT15w2V/LtRyi8V4WUcJy1y/3ho8VOH2Y6+YjXSdNxAHdApfMAETPndh+u1k3
or2mkWUuQzB3uTtud2ODFg9kbBN87U02sWXnqTZDjHAc6Qt+DG6XiV7WMngTmc+f
LAlfPTLs4DElPhil6wprmivg7UGhGA16w8dd/JIfpUcmaj62zJ+JrW5dWe+Y1qGT
2IStf+cYKh/iw2QtttQ8tuuE4nqVgccwH0Rqh7q1jhoqyqKV44PNdULlcx8kOKja
DMIE9LgxEnR8Pz/BlfLJUA==
`protect END_PROTECTED
