`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
09OQNnNZs4dyk1xPe/w1iptA5zWHBTD47fSkAQa0/KL3BjNf80IilfvlsdSsRK2H
UBaNCCsd22/YeZf6OkmdAFiJfHM7Qz2ey7g3HwG7SNEPIZ3pBSPjGELUcJIuKn64
NxHCagWWDBakYTJDVJ8XT1iGfjTA1V3bj9TCvVBdGvRAKE/xPziomm8xutNRNjKn
B5imw2q+Ab+ePpgK11VgZKWCIofS/0sCmtKjP7NJwF1mP/DDS8cHCKcNAMUFnERA
wzQBGIfs+eXMSPtMoH0piDK5phch1zWWtuScxNA7jr62SkBd2R/o3bvRuyonBcSE
kKAjSaMQxwC3+l9lcxkv+hyrdOg5kZt9DcO2BzX2jY7XMXAm183lkdmAVw6glTln
+ibnZkRKvXfGbiMXMkf99D9kRax5FH9lrdyWA4bWlnUENmz70O/oWxUi9+R5J46U
0P0aA8NXdftkHyzujvmbmAGpxO2zwwQMhljqW2ULSGGty0YVEJPuJe2D+EkbWhYv
nzMLcMl2jNIkNfgbZBqg7A==
`protect END_PROTECTED
