`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hS2j2yTRZzVvbK0Q7pZaLDli6hNxQdOXQV26obPSZQ6SYDRUo5F+Jx1RGFj8oHi2
4bkFsTxWMvF8O6UCpTBnsUjVzDyhGLjDRKo0aaLBd3JUJX4VBQvZzy/OeUJ57PRi
wE+claGKJW+1PhCRUkmqninII24C0ZFH9SsPZnsMfkkiwUtkoQZhT0QpPwrtumFB
Y2FFKgeWmWOD2of1YemAAZQB91VxBamTU2oiMWvgpG/yFexDtdiLvmrY8sOS7F5a
g6vkbw7LspuDPczaOg0eYAzN5G1kWE6ORwVFMJb7qcyHVi3h8ZXzTkUAqNsiyOfg
DHA80GIzoLy8z0MtKksTsNro283vypFYu/+oMPgIbBjPrQ/ogYb5Yis2O9hZ9m98
eoQFLsq0FfFUEpvDklZhrjOcTz9OXmNikp2/i/Fac1eRIvKjD/9TNN5G4la4rg1V
kVXNPdVg3JuKtMXcm6I3BBjw8H/37tR070Q5ZPn1OeiDT+2ygXt1KEBvZ1XKT8o7
rFgX4+8y5Y1Ke6XQG9OagU9bMLmqQw8nfAatiTGilrLUCJk5Jqtt5UB1LIffDiWA
oxpZuoDBKnikCWGLxJYHSWPQ3JLPP50YTxVIp71t022Ah9+tlvQ9f/yliGkGiJpZ
g2ArfVssLYl+zr1KP5p60Gdj34syKD6tIypIrZH+EEqhwjH7e0ZMj3siV0XPIhE5
5utAewp6oxEpW1MJyCs9xvce1I6KPD0MpMeB+6sYJpw=
`protect END_PROTECTED
