`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bQN9f/SanrFWFllcCzYockRVPIUptcMoEThG78kWPhQ/5yNdatQnt2RN3UEatH/z
/Tx8UlypbaE1ny2OWTAZlzBodBbFTxYZKcZ2I241TNRKHZl5UagR5spRQhZf5Q7t
vb3hIS4qSIpbCRX08yjU3JXwZ7RhccR/3pO/WaGKPS6DjZ5MLD2TZQ9mlVKF5VlW
UujN5YQ2gH+0W0NIN0FRfczTe5+oSlagXMIuJK2EkhZ3qRKr/uPFghfIRmhxYv7n
QDcujlQTxX9vOlrZx93wWjIH9C6Hd43PN0Z1sSYXF9gMyeQul9z11LD3CoTvshIF
WgC9XzuX96MjGM9i3aCy8So84Ioyh2q39YthgovuIbWSt5svyXzMrx+9REx6SCCh
If+udCWeMPFeB1gQ16aDq+bDLt33hqvG63UKwc0wmV2iQZud4cH1XReDx7xZmnVM
0hwc7ZIOkWyFcz3HXhb0LHAAQ4kQ6omXF9JbPibUV+Du5HW1BjjEUwpCZWMu2gV4
lJzngEz59jxgTYGx6TzZWkPZCelswNHDjTujfzhyIjF9vYqBYvV5zsHjnhc2k7Er
f5fOM3JgcHQuIKcNB65F4V1pGjHi0xH9XBFHiMKobYT+LHIP9sOdUMPdK4IuRxIg
AiW47rONIqakJYp8K6PcmZbUpPhB+goNfut6LmwiZFUMiWw43gySxSFHzPu4zVmZ
8bKY/+8Xj5KZH05w/+ERelCkEzmBpUIEytXPhftZsdgrKOSqBM8K0jm+ISMmVl9r
b9oHhTlMKaCwkyqC1NwH5nNXtaV002F8I7BzDcT5MhtiOUgRkMkmh202XNoJcao1
SLYUFfLJhj5o1pEtgwql4a4YZoKQ7iFfgpTvNrfpWJAwAZeikpCFjMoxzh6iujQb
Lj08st6SsUxn390cT4b4LE8nqk1x8V1AEPuAz/NXJKQ=
`protect END_PROTECTED
