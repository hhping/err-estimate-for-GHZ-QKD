`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
prb+5gRK4Pcs/QRZKdOWIq6bIi0lWW+5/LkOkcf+vYaz2wDWOqfCmU5dtb1T57Bp
9y3eFaXj3Rsf6I/3/2WxsbsV+KsOmegd7qUmHU8Z26fYaRmWITOTD+6vHobb0Piu
IlKOSr1qnIbiXWzO611gee5KE1jNfp+OEvC+4ATq6E2kvgWQWmW7uiEtlRu3vML3
E2fH1IkEkA8m4tn5vw7I3B/YFM5Q61IrGuTR73DzToEPpTrDOsJ7URdlstUNAbHr
IIZCskIb7oyUltF6ZHwhy9O3w7JA2Tr7PyfRafBzWdBHWgK/lSRthRN8LQ2gm+N7
0bPAXFT6ehtYjEN9st6/Yjr35bmktyCboVK4PuzPsO4zgGbz/CkbILfDTVOwkO88
AdvAJjs9HxEVJ3NHuVTNe+8tNCPLlPs2J2342HFXVdSnazmyaw1u0wRQaV4Giq+s
wXWb8MgCqALJQcn9P1b48eMT2pzXPa52KqyUgAmbvSDwB1Gc2NtqzRTtj0WjdDsk
gpCjmCzV+NGcF9jEdOdyaQ/qvBYCCXA1en9f4x3HdZ8f6D5M0qn72PEG+Q8pP1ul
lWIHFpGM3OZLRzm6uuU9hUUsSwMrwaf71L5aHKAZDjWvnbQApM7WAhBhqiEvnJl5
zIajSVjRc05jkffv17Nedk0TDchZcShhyyPOoLGIFDuqNucYPUh0eVtk8Kr96uKe
8bPsKy8PXxgx/WDIBnNNW/K5pWLteuHS/aby2Y90fM4=
`protect END_PROTECTED
