`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QmOtP7yJ7AbhZBqazNTqNKn2ptnKLASfnJNR8AGcefSpZhWums07cTSmsVg8yPAC
6r1FdWZCEJ+ELZRu3OEU9Ch/0SEqroKwTfwySXI2Z6+UGNr4FVjcrsOoDgF2Jeqa
y2ItgeJXo+8XnyDLQaBk1Cx0bmEhdbNqKpBaTG4jWpYQ0EhKdjIUpu2ON0PPxCWR
NrcNgFXQ55AFDhITBFQK1+53dnRii6pm/xG5xQsG4ofljIsYXhSI+fn/BJqyxUkk
LworoV7b20h+KPzhMKGjqbzcHbTXsiGUaNsL5fFp1FOy7eoyFWtOUo4D/ugd/YY0
xXNMyLT9fd+qAgEELF//d4fm1tDdYPuEngQ75cayfT+SWQZjUINAOsZw2x8Ghrcz
yL0frPAAw4X31a27J8mDjppP9rm7HnuXoPQIQN8X1S237Ueixa8ILHqQfTCfyir9
qetfqgyPSmiHIJ2vi2pUjhcZrm5nDExQDXooojxeGClCY47PQlNlTiU75b7YRfhj
EXghxisEiv/8D1270R/IG3WfsHIpF8wHKl4+R34H5nHNg1YmfCrWoQio90bn4SDr
0MEu386lu7Efh62MCVzksXM11hxVXH2BlQp24rVeHKSFHolFEZ+4RUDzFweQietD
ei0CGYpVsv1u58B4zOwuev9G/hmJj2IiKUhTqgrnU2U=
`protect END_PROTECTED
