`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xm8NQpwJNSe410CMBToRFLw+NkVbuvR3WBQeq5blDRuDIsXkPVvgKOV01697Y5vS
GzxUL+YHKfkF6o18igVatWHrRkyy8OD0qSBMmCqwhandNWx5qs2NeWw5OF+gDlR9
VjaPvvSbekL5fH0TP+VTNxABD2Ja6sepMEA9imZLft4+c7fxSMm884fFuILnu14C
ZvcxRnxvJV4y8c6PKzs8rtpR7fw/Aikz1zbWWWpsrpIJDOEKsG61OOgD5s182ZJd
L7/uoVEMcehFxFitJ5ErslTZ1Vh0lg6DZa8GYLA/W1Enx2LDBJPlDWe0kGIPem6q
V8s513ed0ypvCNaQzXSxkXHNsNersApu5wNlklgGf0p+QD7qDofRJFnFJABaZo59
dCvxPvQ1YruG+gko5bhN9IUaEHclIjpxtUeOgP6HndbOuS6/3FTCZNOqCfs9AEjX
H0iZPqA+yLhyNogCR2MP+qLfpCo5yjb2y82BLgJWOiMv66+fnrJdoRcADYqZck8q
xg3SxDeO9yn2cXtuvw0zzugSdC7qNZ9g3lPKy9ZGjDEQnnUopMkm608rJq57EiEr
CFb8ifavVijydfaeTnZ6BdYzQCzeC/WPtpAMi8icH13zuO1sXHxuqSXp7XCP7zEh
sMYnsleuxGkv6bPsokTUB7I8EE9mWJ4oE1MQnbjwOuJZ/aEgbDMLa3bzrNeNeYtF
g+c1xJcFUb5SY8WJwsknmJD4sqm29nZLYS3WHawWQxn+43b1uvlStpBJC0wyGxIY
1vzXSMxs2YBKw2oerLDHtoT0/6SoBzEXl6uR4cn/bdND1Pq7k1gGmdfqkoXDtTFi
E7x/9gcBx/RzY6pQpLx5MI18ZdNoendxsMfWf8KqjsbAKfdDrZEyO07+VzWWue6a
3ZUhv7HSSzcT7ddt9uLdtaB14zhgYPnZ87A9LvDiRP012dINcD0vqd/AZh24/Y+R
bVcVFDPdXW6C73qQ81yARA+8wHCndTrza5W41dl/R4YB73o1VKrRjvj5IAVhDJ8X
i/I6Qp42JkFr/8dHlNrDq7KWqDlds/aiaovXX4wH555Tq8ymbW36lD9dpAzN2sie
4Lw39THWu5SkmVCn8fiMiGCoUZQ6ZG7iQLCeGjClPSqgSeTvNMOIU5/sdmAbWTn3
AwXb3xTxHUfW47G6EkC9yzwNnmkuQNo2ews2Vz8BKrAPFR8iOeD1CYNI/Aw5mP2H
l7U52s5tvrrXy1vq2KakVXbCzX/gCqDGSN9ILf8GLcyhgNvsDykhFNlizNQLlKYf
acm1O13iSEtFYudGNEFHbxVCQjJDr9sEGQPyj2sSOw8UoBRPMgT6NAHrIZlGAiah
5hvjYCKM/CBGe4wM+C4Cvod8OmJtU6pM4YKvs0YkSqVOFnO9Cq1LPlCEJFICbAkU
KxxHXLQj9IxE2fbvGQDu9gVNMpLeiJ8gUye8T/t8vkh2bnQVcFdyJoRxN32vSM/Z
MYHip+FzrJus3gcUC+qbUZQ+J5Z/6uEG9PbkztRFqKXI++H2d1+BTUBz/kP28R11
dSjDzUTNOVxkEyRrHKkNWnOFdjTH+INiouupVbBOsUs0BZgQ9DxTfuOpWqxXUVK4
jE9uvWLdaaUK5FiTd6JuSNXgcaZpUMgnOWF+4bBPOt9FbMGPzck5j6XYNiUPVQIl
AcmKZfViHcUUOsqER2px4aupK4b9wIYNU2Sa20endigsEEQNPU5emvMbDH5Vrixp
2ZU8NehlpTqQ01VXOqMU9wa1wsKohOF4Y5EB8o1yZRX4rMyhso0ykzFcIqwwB6Wg
H50GB5TrPPaMtYK93wZIrasDjgXLuxqlkY19cHYdsztDNIhPYY/m/YXkc9QiuJ5B
dwW7hGq18XV6+CHkLwEPpld8PCBVYfBdoyOUZ6qFODqDLYIHRSjGDasIlCtVuzQY
EgEFPZKboEZOH3xuyj61usu53MQtcji5hrdmUQhAyyK1UmstrWdWiAgtd4fx4l6c
rV9Ah2SvnzqmFS3yUEOfb7JzjueFpkjggDvh56WZtWxQcNxxF+ezzYoGTdPvOoTJ
SNF47NOTqdZNsv8UNh+kg4UvHTRiWPrGpX9xC/qYHOUzYiukEqhoMvJC/bbaTKC9
T4kQU15TqDkkGq+rPH068FakpQSMIIuC9dCIdNyeHhKH1rxI1WbeFp5YQkm6eWbi
VbUs/bBfYethpQDk01g2konm+TcjBQAkBxmE5OxXa/VjOysqiOtUBVN8rRz3cDAM
qrAPBaouvQzuojAlqzlQ/8eEVIgKUrZ66TEWibLp3clgqOZQRlHiJBJOmV3yvBAq
/e3p+qxLJtQ9XCRUMg0cgjD4lbCt/eWqOcDwEDSayJNfo2yYIPg+3PSn8sP15u0n
g+gwhJKJpua0e0/k0L0Rr1JIWckGZLT5XhxT2ne+KRAYKUauLW4ztQYnYNd0sFWd
Jk24DEeTte8rwcbOyFFXWZp/kS8ke+V2HZauqgBGVXwLX/4QOSoA0V1pbcZvvMZM
CPiQjV31XrDfOkHlBtMkow==
`protect END_PROTECTED
