`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KX5a4M7/65QH5Z/HXvAKRtlnKKtKv+58Xia+sl2pBwBAhtylTlTTiRDYRChO8NVk
Ip34p9EGGimW9drXEcO9aQfjMQJG+pcbbITsRFn228OkWBgtNHFSYe7SYIDt+ASX
0H4N0T8AP01j+uZlWIr9oUpVJSnzZQ1BKGfox7W4/rGQDlW40U2KGabJR90oz5/9
vgpSW8f6C9U0bPPXf/49rJolzk2avxa95pkB7Jt1klmKZkImlQU8Q5a+EEhpxO9P
a7YrEqKQDOMfNnyxn5kpUTaaSlHTIcLt8ZoJ+KB0ms+4UigaS+SIeRnU40wH7RcT
EQSxTXc/y+jZUFSdX3sc+7PCx+MSa9s8UiId6UEqCFoSssdaIB49yafdM+zB7aqi
9df9CmFNVee2lI0dum2Iqs+jdoxcn8W708QT+yd9A9wFkVvMBjDrRpO72zqG0Xk0
GZ0PUCE3ChkkJVHC5bU/cHogbdo46pn+oiOXCGyC6mWFM8OHmYn4gKZhaoaSM0Ym
SPMfwUhnwyLcFSigeJgrC5GH7qkF8JmP7N1bOpLU7AT1mtz11TF8NGX0i5CFTgyt
DX3t8zJ/jZjzXPsc9nR/MeDe1sJNgYt6oluf50TGGeJclrkx2c9VOZ5YvyzuoX76
llH10UNpxxWLQ7oZNfvUYA48qWwLY4ManWZNMJNTrH/Hl9lC/zqjqpncHGc5g+Ka
W1qoX4I7g/KhulW8S/c9Tj89L8gnJP0PqpeuK0Cb7lM0AMpqgS7JZtRsvYoD3qCM
nGYaPIZNljusYtPnczZAJwfiteEFBN2gkMaI2pMTHg/RaPKwUTw8n2FHmqov+Q/u
36sNSYDFDVYj8l/FxKybREObOT09gu5VgW9YfNn+GUNskeCCDVj67KTtlGcKycgQ
OI4FFy3lO7yO282JfrLeZL5LFoMQ/Ohj1BPaEwzXW/TADoSW2Y5Dv9Gcg9shzNVh
zpWdLm8dKv5LwX+UpVTgBO1fI4abSiP8vRLu/oid91widMI/x6H/8PY0vdk2jWwG
zlntGQsWDsT2ThOFEPxHh6BOT+Ld9tR2xJgW71Q4tl14APSPWYGLrV5SKEGm+0mn
WK65FEaDnMOFT/pD7BFe6r9mbtq3lUjxWpWUkLz9Pv6qD0drhOA30qK1HxCArY0B
bqJwsPE1GhjXO+YySB5ve2rPts86BGejq06G80qd5NtFFjdbhL9jxEqp4rlx9agz
NC8Qgp8wi6z0UhCLcWo5eg5smZ8ZMbGfIM9rV+djFtehAHbOYvDKhNIm6XMb+6hu
//wFTuQzcU9nBnzEMb0zBibs7ws1tX9VIi7FMD9gi4eT/X2ZS1BKB9dwb2Smf1lH
D/7jtKhDOjoeBIJaPU76huKnYFbHsaYvs5krVOykh4aaVWqURkWVWcvTt8AVIuHs
TBGv612nfZlTGMFXr9rrqq/I4YcWBr/bKrze/OUSMxB3DOQReBG9D6xlz+iZN+M6
xIy7zY3fNR+YoY+yQm+7I1EgVfxIxyJDI0P/GPIOuEmGaQwHvl+Ls28NJ6bNUbwA
Xs111a3zdXhPeEwedb/YzGXZKIWfI6vjGzvV7+ny9IJyR8qkBryopMwAhHvBU/ZF
bZvzowyav/OEG+djX0hWIoV0sOp7op4ov0uVuG3fG2vGB2o0lI1/dzepRjhkqRmD
bWz6FaBkYK48Bwld81DzWsomR/Ct/b+Dx4nm6qLea3GyFLyRLQJkNEoxVaArYamp
e3H6jPfG60+eUZSTSTUMt4hbM0eNcBqdt8Y05E0yIY2aAQ6IejQq3WwPCJxmrt9G
PO9gR9fgqjsLJXKr/9isQgN4ittEDBikMQbBVYoefRKJMjiAhkYuenI5PyckYBeL
qQ87cvz39GtVkqI6xrHfl/LOTrUxOmbOtB3VyY0gqHTii+FXLah16Ba52qpu7t6u
U22BigqVOvhmr8qkxBsJNW9Nkq8PKVEi3j78gQVMqmcjO5ecjEs+dzRuJcqP7+UX
44BjSuW9pE1kuNIcqseaLpzq5uMwXG/mLyac1rLiZ9gVO7O++4ZYIPUetp9T7nJt
iX70S74yUNX2CTZARrMKnIgj1q38Mo2ezi82uKQkVl/BNVHMHm1s9GgxxPOoepvq
SAUZvDzrqXCOmckI6D4LbFGKZLcNK4mVqcd1VISWKmLpGWEjv/+ONfbqEUgy/tXt
MZPWQV6oQYfP6LUgg9ExspzNdlR8hkvML5uc+/BwKMYfuA1b5SDY4vX1b733Lq86
fQQhXSx8O1OF/9wJSlutPAWDYnfgIQNaPaWupS+DQvEFBAs2ho75FwKBd8UnaA6q
sV0rcRoWQC+9bMsRofO53GrBlqLbUIdLMg1EAp2MJkmlqFl6GupqZHgLMiM6kkYf
ydoFs40eIsdd1/2KbYYf1SeJs3ec8xMaB+NlpqYjj/4LVG2a8VJOlApkJjDC5oY3
Gykdu4HhxFWYz2p7V8gaJbsJRXVuLq08N3QYbrIbfdAHRoNL0MFvSzpDQNGetPIo
vwiuMtW/STmfCxjIR83FhMDEPrQV68OQwQ8Tc7wSBsxpSZAGnib23czOiblKMs6A
oQ0rEfjMaJYUxJYFAoO+ohTjBQ9iEk7trIlO4tqfWZCniRErBoDpp6B7gME5Xeb9
RwP08ODDSxG62zhqBrZVAUK3JD71buCmaKNe0Tj6Edb37uPdRZUh7ZmASF2HjDfc
5BDnqo15HuXoF2DORgeWgP+fiRE504u81j6fSOmBk2ZAbNrCvpVRvPH623dBvQaS
HpZDGQyUFmQRl56U1kheXdtjZjnA6v7J4U8xrZzDVWFkuPcpyQhtYspxyODpHjEp
xpYzUsDMd9NQix+XpvxNUO2PwayV6oF2DlCchLfd3vVfzQXCf4zeBxvW7FRs6ARG
W0KEHZJ5XqO/UizdnlMh3t1IHkDo5TgO+K6yKlfrIasoy439XHGLTOFfbdbCyzuP
IJPb17pEyaH5kIIBjSP32NZzivuUhJozv1q3v/ZuKEGcQzWBBBx3IWgy2dxicHAK
6KopOpuIlVCLeuBfkDzwHlnjlobFZU6HWzfMDdWodwHFw+DbulvBG3ca/i41Q/jS
izb64i/PuNX+hl8ye/T6sAJVAil4TbZrjEUza9Me2jhMmm0rWupWoz1fNFxBVX3E
YQzDn8lCnbdYai42/nbQxY+im7Pj8wyYgF1RCtQFkgisA8T2fVLosNTUH2N7kEAd
33942yMFoAD6i7/s2OeHsd6eRiAi383IKH8d+u2KH/fkX5pgFA6pLKj7ayD5YO6h
r/YlfU10gq6DhldHMJrA3rVk4HTH3Zj05Ltte6Eqi/pUoFNnzFLlqXSXPBxiBmy6
2eC3+zuzDlZafHteiA7ZT2U1BG1DECUpx7QkBRJu7P5weSoBBRgnI8wVxayySH53
5VFE6KaFazVthdBgqdBsBLnZtfNuEhaANFIiRXPX1GzoWxVmSZ31Tr2cbRTrjfat
AKn5ojBqDk1ttWcyMhV7zo9R8qZlHZ6AlGGZckwzeYnSexJwnCL4hoARm09sNaSz
H9Aeq9ZLYNBr16u4TRfOoWDjKwGcppyERYkMx8224f1t26XZ6YBKmu6UrW0Zm7nh
9mHI1vdA5dY0wBYS5E95u1n2QyhXRRyhPkEYq7mQOsUHoMWs8dRHQZYjCa25FUdB
c2VcJGOXBA0WpiTHjYScFF/+GuaOlkdpPLmiFnE0wP99BdSu2gc0/upLZgNr/hF2
9/IkXvsTYR3Kw2icBqoaarfhcoIdtHVgBpfunaj8/qUDgCPfZjCuX2cBnoiTA8YG
JlrhDVtjbyt5hPVIUKn7+AhZN5brP06Z6gmltI2d67uFMwoJgQVruHQ1en6/2MRK
pq0cjgdRZhGWtnOG/GMAzV+CkGZa7PE4SvknZHYRI3hpjpvNJEshohHRdgHNaaxL
wi5pP5dAc8u/OayfZlB/wk/EXgtJ2KaNtym0kc1LykDE7qhkdyqkdE2wn6nb0kyo
37xpKs2HqiqaOLTimHRLFSQQZ5hEG8g6ZUILKgviqRcpgg4i2VAMlX8WHzaccb1Q
iVOvbna7gx0ZfZCYNFUAcmZVvwQ6IZbjolv3o4/LFGNDRsQ36affDQ10s5EO6wlx
4yHrlJ8EuR4hoxCDyM/Cc0x7NE36eQd2bC+7b14UpbMcTn0dj5PR6a3JfZ/Uyqbg
ETUq02RNGr2oqUgRx+hmas94Rko+S66NX3fzITr2d5/QB48bqxSleDbOx36Jq2FC
OlW4rPrPE30EMIovx+3/5rKKIB6zSE8kq+tLLM5ohm4BV5UPQJdY0xBc2CjPb80s
/um0Z47dOJQnwUu3MmmK+qk/0HhxMrnHbE+CDOrDtjgN4HluLlItFpkbyZuowNPf
kDR+60P8zJIvh+J1Z23BFHGvEcGjmn+Z1GqzHi1iWHyqz331BIfNKLrbooAsUTRB
S0m5mZ6bHzw03EFgjpInMzYwbdBp4BQBLN6eYXbNnL+h1sUO4+qGVF7AoMTF9Cgw
28FHDk6kRkfMe5yv/dpF3CUUv8hFsB5HAO7XeIO80RYTwQ0e771BG3AptkoFPh1j
U8YatmiHxRlj7qbaud0/sf+/FFuAwgSBlFjyvPN1/SY8zyLT3ppbM5/4n5qZBQ5/
uEOWiDNjUkOLkGTduJYBbKEMrL+13f3VSDR9+MQKbpZlInj0BzYYjg3M9B5yZZRZ
r/8ncp3DMqK+ZU6AD7vK4FMls7zF0onjJmKwFK162RPS4uZ2ILmAjFOjneOcbqvr
cO1LqQZoV8dwmwnTqmPFdZL+mfSEtCdQ5KNf0gim1aJjPNPvSNduDlXj3shFb8cy
joRXHp4/w55E4VU0oU63AhRXLpAmUOmSXJH6XAYgCYFn49q+KfcEs8XYF0L6LfZg
nhDbLYToiXxGAL1rStDggvlmMk+OJnsUv5RCgepFCNq+d/IQGhOdRz4ZsfgcPVOR
ea5IC5lTSGd8G3/yAWASBlTafzcASn9YH7ZSLoY1G1T/pYX6UeuPhqt68ugvW8oJ
aD8ycXdhJS6gvOuce9BD4jvvncZRisTTtaqjUu92iSuzsEmq/N80ioQ4Rh5Wz+Ir
qBaHdfSwb7BnXpApgpC9BTR/bXto8gyqgdEC7m74uchZsSkDTP0CulNuKhzeDKh2
P4DcZirGDaTHESzM4AMdFx9CIrWhhirB98WW0QC00mJK4fy9NqutH3EkJu4o7V0d
sRUuzp25wUaogbI72u1G6/5z9ElyhRaAHQPfAlH7biRrGhsxz8SoKPjXNILSPDkt
6SC8fq5q3fh3CUJGaL+mgYHqe7f+8wcXP4PAnFKHAZd2mIKJjtdfcwTBVL7GE+E7
UAoqWrGA+gD4GnCfLzcnCd2X7a3Cbrrcunk9Pt9gWwCkOPx3h6L3cXyxYsCoF4j9
z67Miic0SXQqXhJ00AApe/YDB+UBG2jC7rElIyyt+pgWIjsAcyjcZPNM4DY2ouq7
aV5ZP8+J53nNuYRd1U2qMoWTrT/BEmhz/od3vk1e9mXMVY4upnMOfD1+987UjxHp
35eomTa85UhZwbB+ttE60MHLSI3uYX4upHMiCyil/EtRDRx9hfvApfm4GD5f3Gaq
KIhOCKulI2rCD2a+XUq3UeJrG+CMbXP4ZuAfgcjxSxZqK/Qc3YRRP/nmQEhkLFwR
/ND1BjDpddgkz2xg2BoB19xReyA4rYBOeceH7ENw6KakMfLPXW2w0qG53frIMHuR
L+5FcEBY6Aj5auC2x3ffsvOLvgFtBTOzpj18U0QFSZkhWos0Fio+uD7Y9wfUjEpx
RDyE8YwgekOUAReEmhH2/V2yhwmRVLkWj8d8+22F1qr/m8x65hrwZ76I2jBgGRc+
7M/iDGJE45zG1ifnk4p92+BB6N8/BitPsB2IjhcAN/f8zy88s/r9OAJKnFDftbuU
iyd3K6AKmkXyJ5pEDQogAH8nakCib0+T1nt6TN5+O1DBJ1vakGFu97R6j4CZZGVv
1YUg16gw0zmaiWSYsTACSvG0zIlUWX8aKhqh518eVnwNy9Y13kOjqAr5LgRo1lb8
SFp4ciMBpqwLXtHah09FeSaf04KO96NFmqU8bz8tn3ytbYkrZz6vOvttjT8SWirW
Gv7Xn14loE7/pFJfvnBGJx0qJaTJaBk14ZuW4ZmQk/I1Gvf5Ddda4WXrHxLjCYW+
FbVn2q6QfbKT7XPLSLL1av7kk5XY4T2WL1WBHLdoHcUsCCIlMsmWQYR0fvX4yFBO
rx3+xqzhLn06REr69wHRRw26R4Jwft0RoWsGTPHVzNTgN/+x2YbhtGePbV4b5EWD
Cd5JMT7ibLnETq5XCgfprTW9xqk9qn+v1L1rnGAIA62TyxEItw85d267vAl/L+Iw
dONRG38ajJZw92RzKstmX0wCZK9oPZ8jn6W/wW3xmqrxMAY+mI5xJXaGG/KLG9tT
vQrbkOZEfCcTLdfJeyAZTNUzrYiFS6M8uUdUxdaJcwlqcnCW/0iIiByqqf9XWUSG
L+52k2F0zQNkDaf+A58MSoGTS2GOuQMrFf4RZj6C0ncLKpJZZS/hGJ8M7AvVCxFL
iDufoQoMHZoLTr6aGvRTc8LXItFYMnzGNqbXo7nAxzVi70PCyssSRPxRqMG4imJt
CvZDCpsmDBIMAfUpDE6kyi8g63q6O4I5XFqPpOmM7Oz/qL32OHgYn/WmIi1V0tQL
gVxlBm4Q7Odc5eIM3S4kufviNvasRE2RuqL5eve56s3cKy3EyxsuG4Am5fx1JChx
XWdQhWEUZcF11I4zUwnRwBVFkc7v32wyPKZEd8G0/DWQ30hEniZbALoHBRJgFni5
9n16K7o4I+V+SzI56a1APX1rBzV2ZsDvVOATqf8FhS3R2/JTvJW+WrSwLD22dskA
8jPHRBfEpyMiE9XwJiW1oZqUppUlsGrZAIMzzLK5ZnQkHA2qMZ+j40nrcKR0bUK/
QyiKlTkNpWHcNjHMOzSOW8Umx1QdEF6ZWsFIuQf+SNfIoPOD9AZc8gsy2cu+ZGYr
xIC20//ahXNTOKExOHcqqegWm4/WBRCvHb6W4SbF6t4aTIWKS6r4wDbh1epEbrfL
+3NDuG5Ko5n4glcpEy6Bj+Qs4KZrzk8x1MLJa8p9r8jw02vuxhVpNpWNvV14Xr4f
7RWlAKTFJ1poZF1x6s5n29j2zycRfgZzkAgiTUhMfloa553wkwA+PeCn88KFPWWn
nICszwIBHuk9ABJLOfhF6PsKGvpxVNpjOrSvZZ2HSnNN+VGmyCBqNSpVvCjR6yhP
Jy3YHCRLRKEMliJ4ioQNl9MDGOGhNIOz2FP43EnuPEDQBv+RibcXnPEuMxi+ofCv
NmM9Peoj6Wgj0S3pVELEEenqPq/wMVnbCj8vSSl3Yf4bRCP49TMwW+b2EOHxL4gG
BPxI3uI2Yeko5SRKxCxleAlZuMc24i+qPB6JXHRvy77g72Gu/SqZoCj+S2Y8r0Tp
mha18mQmWjw/G+4WVm1pu+4Fpjq21iG4YYMKOPNlLCR2drZdC+ePIc5UNN0G+9B4
VNONcNlnlrTxNXuvbRS4I9J462g5Q+MMuhR2AIQrVW/IpfZwdIcigslnimsIgLjN
f5CNngzkDih1PpR5XnyRnZxTz8bj12EiF31Way3R+Q+lN7WfCDNFvRC2q8HKT/ry
lSorcwz+Z3LYzW+rMCjv3vjBQLzZVGUpjOHNbAazPiLfjV4TdM8HQryYLIOocUAm
VUpmQy95TU+CNDulrbLjDjyzIUhUabK7I5sMEDhRkK+RSCWtb/Y+EQIdfy78ov90
yocnngB3DNZRdIdF0j8094ufJaquVYC1l2MFSgcQf9ZvnOYzXaRCgKVYPSsG31tq
BfdOhigYAfdkkneI7H4WYm1d0n6LN9xen9Q1J8MP9wNCwSmniRfFIVr8opn45qXR
cqSLIKTbqdOx0+kLoknDH7k1WMiczlL0kyijvIL9B3ZOLuFLtmq51hF+cwfkAI/8
ztffBYKlZKaUsnBKCcF0xcYeBocJKUDWnrm9MoI9xWHjeon/vRs7dtRoZww06XjF
UhSGjmcvUQrDrcfnA2cOwKEuhlhayHDMa/6ESa2wy/cfTai81pAYq1Cm8PSGfBVT
Uht2UdcpUOOsTMzchclvZ7P/mIfeCJDs80U4teyRkizmOZj2YnZ2e295DRkZYJdj
aAfJ+Gu+mkd+zq32rAZAjcaDI8+ladkMADcaSmkMHE81jqVEt3ngt57YSjp3ob6c
/u8uog2aErfpfmU+RLG8j3FMtRzTgqGpUnk0Do9HLEg5g3wTUuOR4fwbC1OeVdHZ
2ezICaWrjvrI2pobKLUul5yeq5qI7W+Laf1gOrYulJwpIDqU5S0K4xeLnCAl/kL0
du2JhFuuEZsAJIox6REOdoWpphOUiToX6JAyhNPAAQmZQO4Sg5nZ8j8hyiMSL0GI
+QRGZEy1FfP1HirgnnoHYGJx7dusC2c+UpgCtw3bc5G9C0StstQ8WBGgBd8eGVv7
tDR2ohIDQDMi6lEyf6c7cW6y+SbmbJpLSIYEYF7zUt3vTaGKZ8cFgmKBRPCWBruQ
1wqQFH2Y7FR1unyv3UAWqjWJvKMPYNANRFK8jBTe3P0QZWW7lhukfubL2kATcxRD
Yt59TTlkEzm2SvH+frmi+dnNuGDtPv3dADEpBe8Bf1KJ2a+mwP0zoWQUO9T3468j
Cr8PZXOsgJdhjFtBcJgUK45yFJCVQaWIiqUnRfXboa3Br+elIYlxlUBAKe5Lf0Cl
sBcurGivvqWv/pDNI6u2HrzJZR13k93rRJDt1BMX/SiUIGdkVTRtrTNICeZdsobH
JMWBp5+TaQpY4R4fK6lJx+YKaPAQYo9g4IGxBjQsx4eW/Oq4qhW9SPbcFqQnjJ9I
bQCAABLnYLxDF+8DlXv5tmLH7YUwTpH7ABFNiyWNjHblX06e1svf43gpBVUSyf1f
cLcB+FA63KAQov/D3JGr+aY2ktLI61MNvd5+rnZXThpSs874iO714fTbfB1v2D/Y
to2AlvOWoGCZk2jqUDy3lj1BylEWfPyMHWjPPlFfuMyJT15iL9GlFkMWO0P9PIxY
HqF8FpKqm66I/Sn3rYcV3GYQxGM28aQefPNGKx6ecp/3gt8M86Yh8IFfM4FsKza8
u3UPQ7upb6YIkdI1ixFevllDBPP/Go9fBfpt6scw25bAb7ZEx4eiChF+Jt2Vt1v2
YV14LyOEmo73cU+qfsfcXnjZxFuKCOqiTVVf35ERD5TPeTI+V8/1PiUHSBbw1+V9
nBjlva+xOMj8CEooLuAnXK8Me0q9XdHNyGLehDhlGvKqn3DED6gtNUUr2UW6Qwy0
fARCO36qgBJVu4/KSPBm+gBt0ZKBrfGhxkoZ3AcMZNDii5DhOqFwqet9upLS2PsQ
Yh3GTM8iNHHlX6nt6hJt4a67vPfnjJMDq6Lh6kNX2EH7cNyu/kGAcxqnffPRD4Nt
PNArPmzKs6T4MTE4eLzIt8ADtzumtka18dQRAuannp1Qb1lh/RwZMTIU0M28NlZp
Aj59jCH6G7NHWClyOzSR4vB3G3lrJv6bQq7mRRUKnrWPQ+TtijiipAHE3JaH651M
wF86Bh1F8q2W/H6hb/11z6k8WkTy0ZOsixcBnn2IRNEOpgH/P8Et+Uiyt+U8DLDp
GC3kt18HOHsDi/pNVMfizzadPmW5RvLy6EKYwMe9ilA7UzMiCWeXIaULX1svSctZ
N98dwEPoSVN3SxWDBwt/p/vYVpk8tE+e1hURbfmoKI2vtCIQYlxXYqK0WP85YkdQ
28BPNbob+f3Mi+y99te7I4vIbNcs0BCrk10MPXS6gLfzr7xuRa1XzaUkh+0q1tG7
vaoVSVpRn+ygA3/lK0ylCiUjkrY5w9G27FYayDnjyamsKU3yYTF5UUUkSeqSk44u
Wd1O7J+P+XUtCl6b0NrY/s08Om8V9roarUxGAwZJJPuYe4E+EIrlOzO7jYqGLSgC
Q33Qj/bXMgiMD7ajg331FYQT+7R+7uBsAS8rzcVyLwKJsBL5H/0ly3RdY+8v5T/i
tJlUl5nILgU3bDxgfEnT51Q+RE/MB6gyt70Kp+sficeFz/XwIA3NPim3i0GsFt0p
sW1FdciHC9BiajayQM38R4WHy3vJXGLrd7L60xN7LhgZhtCXlnegsL+ETHLPoTNb
l6VgMXS+8ajq8yEONxuGVHvuJEjVcdeF/2AlG334D5VT01ULrvr/nvwxu4/Vj0fh
luzeAvm6sSUVUKMl9a24KfMIQew8d/1uZBdewc3dhuk/v/egv7QyETsXRpoRZvY+
6/U/Ncj1OZ/A77Ntxe1qSAQVrVOKnKJXyKAQt3e0p2IVJqEP0YGTT2PxPY6i7I6H
J8k8kTWRv6T3EbXwsKVD6GcUpyPSxsp/N4Xz6FHyEqa7rlWA78vVxjpi1CdmjN6c
n/G8PdJPY3ijY1j/WAnXL7aa+/TN1wtsq1oRoH6U8A0DUuA2nLLUuM8BAj/6PS/8
X604uqcSMe6zMkWEfi9rhfHYlve197JXozPhgmbB5JnJ7+Y24XTafeND/RAL1zQA
EWBkLYXCArC0y7unUR48TpqaUN0a0ldI2+Kysw+VRxc3/G2BBpLv4GqzWhQOJfpe
TW2Ui0D0xOzUyxX51yY6iFGVFiBNNDBecvKllsHm5mcsRS9WbbDWi/nn5chTb2vo
hQZ/l3nXzv0m7+kPEV7WYKj1iDr/GqysaZVtSV5Y1mT46cTFYTSvigWXO6GjfSFV
bd1e/nbRZpd7wWvlGmn2dgN0TDogWML36eTrJu78EiWExQRObudXfqdlv4TscflZ
opfzFexDKEVL092vYt/aR/o2Odr6N5CODcZwHkJHwq7Tpyq1lQkiA7KDSUztws5H
Rli4wapoVqD/P4isDnbMmaVapaHh7ApY/celruoQVq5jPIy8P1cmAn4CZFgB91J4
4CJvUt22i2aAi0DFHTFW06dvoTBrE+LVOfYt6gk6ZMiXtC6mrxUesg6ELwEqrCbT
HBkLkzA+62h7Sd24NWKyKBGW20J1qOWVqRmuYH3HrpEy9BlrUhCjp6zwxxJkaoZh
0xQvCUhWdtdig6iV7TFBB7e8ERb+Xx5gKYh0nvb0JeBPuL40zFo6uAtCEAftdUj9
Exma3dICRHbONdPqSK6Z6mMNhrn3hYVQ+sfIS5jqN2y2BMMpTn23r3CT9N2g6Aji
Ib/Pux5KAk0vQkoHw21ZQ5yjKfWdHFZCtRwlBpL1TCvkXXWHjSoDYeTsQ5shPJmx
UXlDiYoQTqKxYSmxx4sD2Zz+P/zZniPgfOPjPgL9C4Mr9d+AMFWYprAFqUoOzjsc
Eamax/SiJsP/cj4SVTtQ0a7fyLoJWBm3TRb7WjYs4n87BszjKLMNlBmDrauJM66v
149n2Zsfxaxg5MuQgvi7a/c+Z8oKzm3/cSbd0hJnaMRDjxYSM1rrSMS1+5BbsQlN
xZOpchkBkE2yAETQ6UG73tm5DbuGw1733SQY9RIJRVtJ3OfVrVVPKSbbaD2TxKuo
DU7C5DH1mQyvnM+ITg2mp1SBKYxmna3SIexIFWX3Fph8ugZLEyzT5JXwf+aWCuok
7PYnMJYmmmRdUcADALetkJ1LyUWarFVWA1FPC/CHynDB7f/N7mOqY/HqfmzZTIaI
QN08BXF9+/71hiTFMHHU2yGv8xtD1LFCi7ieDFGodqF8QCtwS5xOyqx/Eb44+5rH
dNWTnHlxR33oTd4Bs+iwpGLklSVQ5Kw7ctMNxee5RmOfLnUEzJzCFlvpGEmLaLYf
K1nwC3NGw7o77oWe0/xlprG/1vrWryrujv76JDimivK6EOk20SVRpA+FNoT2iRSV
/bXFeQEvxM2XQ7HwsSmbGaWmQRntq4lhWDyC9NPQoGJpWC4srTad3X6F1uScSOAB
+FC6lG0N3wse8SnaMy6rT5tAwfYl4ttriWpTuSn8jnGw97Q+p852Ta+N6G/IEA6+
CG2tqVn49J85xonpCPmOT+7PTZRU81qIdYWpnfSC+eu8g51PO3SfvNYuZ1MzvDVY
8HCBfEeOYsw3o9GeShcN0hCrtSUBdCctJiSH0a4gzqiBqduNs9aVzdo7ydHHTYUA
y2sJHhHX+nL7Yv/3MtI7ooLNKTFPT4dGxnm4IIYT8JviwFqa8tJ0kRg8MLmeh97j
KwCBTYT5H4yh8XCBu7RqPfCHxha9ydT5422MVFx1gGR/iPbW920O+rDBc4yraHah
m65dqEv201Guf0+LXl9+Hs2M1UebvKsj+6RWjqfsFt/JU1R9nI6+5MrBOMsSq96G
y7mMX0REId5xVQPTDONzkoTDt5pJVlXMjJW7PcZOEDf09AHvp8QAtOYgQ7+86nzL
eQvKmHVafdoGyTSzxP3XQOwhmauu1sQBhzGOzu86cwoCOP19XDiGXi1ic0pQd5Tf
gqoGB2UvLu3GKubqHC35Qpq8AgDq7XCsm6eDA/J5KLSxLq3gM03ai4JjVyT4r6y6
E+ln13AgRA+DVOMe//glcA9FVqX2cYMfmtG8MklNIF+e6RabQ2+iAQtyPD8moLlC
zMx9VXaFD8jitzxZzOttEzGF84YEOPSCefkBCVg5WcBb/kdCwhWcK0w+X7Oj7wNM
pHtdqqdS+UAD2EkgLXhFWiNTXbUyWDeOsOQTyD8qlX9tZfnNyT5JAf6sgOFOmX97
weNyLk5yE+0uhbyLxH2miIsn5K6c04OaXuQ316RNo15WUQN42DXiGvMkaq6cN9Iq
8H7FB/tDCiBtURqyXIIB4JyPPwpO5ae6cyDHt8q7sZK63R9BRjxfBM+SkASsLrVu
6hbuLyZk4WH5J59CGxeM+3eeoIV6NUR32X8bB3WH9fokmftlTzYjPFac9U/jcn1K
XPt0VZp233HNgRTJje7ZzVMkBclBtdXkUm8f67MuVLmrvjyzC25hxiTiieclw2FD
fovfo2/YIit8WkR1rfy8DdcFacQMxh9+5klE/AIe8Z0HBDXTzAE46vbwlNikOHUh
sOT46oEEXiIbiz6nujNxuLnxeqmyz/AJkuQCBmlkLquQ0fx5rtpJrp+x76Etfxs9
Nkc99xGM0UXO591witGAxkBRkvU8QTSrbMgILHx0oQ6Y29uRMlb73UtvXJB4hkr+
6NhPrgBBwF5j424+8phVBvtDzEnM/sTPMqVGwAbnaSvPa77ymUjOnoIznzEmEQ9s
pNvXqAeRdJGq3oyI4RAxXOV4RlEC/m2SafK5n4QVnJxnxXD1q/DTEMqdJakMxMcS
fpoIqmQiNg6MtoAt9h9uTi01mItvXOJMkXo/U++Y7CrDIIxo4qeesdRY3+mdIAw0
4ZKtsknntEabE7fWC2czIlBTVOn43if9yvcvNlHAbgfdutTJzUkQeg2ElNKq/iul
yhrK1BVZ4snTE7jSclKvvHgWUrU+L78pHJV2zO0W9m/mPZazPM/QebwDYOPIt2X9
1FBMvxEK08QeCJJiRexfpMvpfGQYg3jXImKgckizxfc+G9lXWLvgw+2xPiivEhBp
jblEA/CuLpFzT6Abpmdoxpt9qG4+cS00x6BrUFf0EGXMXoBaOeVS1ew8U+mZWNp8
ac7sb9vUlBmuWbWD4XZJUmdZVHETOhMLotsaQE8NobTbkgCXoupG85S2pK60/sFB
fAEVV3zfhdqGBgMrxSSTg0YGeKEutHEVPLwZYPpp8Wo6MBYkJmpXcPFk6rm9m56q
DdGNsDMfv7FdaR5Gy5hZhYzl2ozV52bozzD+zPk5QSVzAMD6hXtVbH1aB8q+A2IR
+KzrD4FuxFMyUs9WAzJ7VTT+56E2/mVSs7bDhJID9ogYfti4EmQgpF7dUSTJ4hpv
zRlQ8rkZYl7VIk/ZSTVQamECXsuIBceDlJXbUEmYRaJrH8O4KlkJg4LyjFAsP7VC
RbB2meHnS1SyPhiokIuobYk1r1DpveR3ShC9n5t4iRbyV8EfBkuG6D1aDXNv+r55
91iHNwIF0ATI1IvOAy8d+lv4IIINwq5VR54hUD+YH7y40oD92wPpctT0aQklmMOc
guCyK6rqdf4gEupH6bjulrvZLRMHgsfhDmmAUZ+OtHNfdo23Wq1IoUqvJ53zhlt6
mmxGpANHmljoH3/uej7GuqD/T9OrtN0ae7O943tczHL8PDlmw6P2CMqZGBpy3Ybg
I0bsnef3x4iOme71CwFBhxXgL7YYw3ic1ZywvoEfW3Iv5FQy3eMhqrY/68JEFeh5
8NMgjpXsoZ/OzDx09eX3OTkU1f/tyJ0HvvTUAJCaHbC058+ReevDDHfGBZdtImVC
x1C1iSsE+szkCx+RoU6/4XuqwhYeyNIOwY3m8uwuKpcD8/0NmEBonc3o7W+ClbxN
bvo3KtZ0H03c20uL0CsruqT2wjcZ3JxJTszsB4HEWIWolKNcyai2pxjLV/WYNO3f
gFkDuuXzbXItWASsk1sUxog4tF24yaKrJvyJy02bvK+pH/5gRfHUrRkox5fuskya
MLc2uNSKKoEsh0SP1zesZywoQrBZXOeam5oZmmT7nDeDxh3eMfDPMt3zo8CZ6V1j
OiNxq/sBNuxOAoc1FY0pTS05PemiGpEnIeu5wXYFRbxEYLraKziwClX23s/A2KNh
dGODe6NpTKJ1vXKjCFqz/2+UcQT2mf9sdhApECTFm3L0bACnefyoqjGFP1x9ScPv
3QuF5JomK6boNrAebAL/w2qIWpdisXX2HCnz+Faqgahdl9DnVEUf4wjMsPqpDjlZ
aI2N4ZMlRVizRS+uejQ5OizoxT7TFX6h2MbooF267+mbzQqinHIvBSYHtwqHdNOx
5wwxFry13ruS5wAYEglIdTwQ1whv+FqINrkEE0/dGclREYqprC2fbAasfc3B5riJ
jaZE8SlhuPiOkW6GefE22g6kL4mDjRMa7AMbrySUldWOIFTMB3DnqlOkLpgyMTHO
M1o26h4DhSY/vA3W2YVpjuTVq3hUt564bYSDxx0DOTh/wEnoXWw3Gjci0T/jJf7J
Foqv+g/tRMxG71CqK5ahsZtbfk4Wsi9Gvh4c2gL1d+NKsYKjr+f7jzJUM+T2RavG
ZeM6HV2I3w8yFkPmsuMrImG/8/Ozgf/8PsFHqDsJnv0Jlv/nR4Sf7fKnsOYnG84r
iWZuNWn0kkwLMIVnBX8AtAJl5SqDbyNu5vr4tYB6qI+VWdyNsp/E8gnLdbWpXGQ6
kvEHSrkUDcjGLw7JWAG16kInbgC8dtUCMh9MRFT0GseAGJdj+1tpH1mXzvwoSDtF
VWr4DhPUXPJMNbe1u4PQndCpBbHc5c1PBACjmCvBHCqyV9I8fYxepXMIsCKRNcbx
CX/9fekSfYJ3av2ypWwlNqCIdRp3CVegFtfid8sOlu1hsG3z7UwdvsaPvaEho9fI
aHADkWhUEZojhxIBNA0OneY4nid97bGg+8PFt3dFc59FLqt88rn7hXgg01Y6piZ2
4c5f71nvFDjjQlmTwDP+SyPg4UH7K01ln/E0qYLLEkrOP0tRfGMXTqEV0Zy7avVG
jwod51NVx3zdm1qLHFHyjIeAD2gYg13qFearKac0NlboxBsAMmsy4gzGjB9hNwW7
AmwOpYzcshR+DEkX1whIm3QWr9XQo89G+hnvUfeUHGg3HwbziBp/yVTGMS2kvmQ4
yk/YkQv7DSHfcZrIBqdYCq3qBW+PCneAy/YSMPNQroHwbiaTSwyWf0ykIZYPRXle
jCT8VZJ8NJX9XrupRbuI7L2SQoZxgk0CZLdYAPjUdKhFME5BQEq0M8sWmCmXY7zX
525z5DaEfnIZjCbjsM9/PuSftMTMuHW+anMSg709jhPAInwNj05hUEIqHMlboAK8
6ZBnHFsy8J1w/lCB0jBIVhR5k0t890+fXoMSCvg8egpvPOochwmwUxaFj4UYfbR9
pk5TKeplJ40A6dDjI4g00/Wy4etf7sHWu60P1P4uZMoT+Ebk7l1YOjaUV2yAioBB
Z1WsKlS1a5GEgYgaTBZg+7WdU0OIe1ItRL33So32rBigDSmF4L+U0q5b/j2sgTrM
Ng72y2SSsF84Hc0ykbH/9KbzngwnVutiyHBGDhZ8u6J8rpNYWchHFdV6r8Xqf2St
ehdrlPRGp445Yc5y3YY9/TtHiJTKBIusH6JRRQ5hTyODLmAzsWymeXUlWi+vz7Sp
/SlA1U7kYYSKBbN3apCncVDrUrAIY8X6qapTgdsr3oPo7u2MU6lhkrY1SWKq0VxK
G1W6crnQW2MN5xL2UdZJg2vjhzaNvkp2kvRPQsQsDL7pmBjj/BhWja1+RsSM/1a2
i3BFWJAdMTYsO1ncsjAh0Pmzl90PAubkVvoQJzMiZzrJUYUYu4cyIz8B1mcIKVue
+MWMr6wLBu94lnAxiaMdmvI9vJ70gsx4QvWw1neDZlJaW4XCaIFDnS028FJIPumL
98AJqk6jZ4uhOHR/43tOHn9P0ZU/Ngvi/atC9RIIZr2TTChqFZHLcdWMCYio7pbL
rv0BHc/b8W23DV8p98SCjztbtNva5VoBVcMTu9hRge7Y0+OEOMz3tHw2xvrvpa2i
KpavFsH/QQh+fXHfLlMj7RBsQbK7aDtsH1ABg4NVJVrkMD1stK5FZn0NEEJyuh0v
C1GK2t3IYhn0/RDRxeYIvdJTcA+5lT3YDuLl9Bc543d7WpNiSRLPTG/qUdus4qYv
Df4jouAEwErIXKYieFKm+ivP1FsgLWSLEvpcdkv5QUTt4MRXy41g0UBys7l3n2O2
3zJJauEhAtHmYuwhBqkKsVPFX5OsBicqJe+FINxyqSl2t9kP00zirmznh2VceeEi
kQ1re+j3a5XwuLnNbb0cU19R8bQx2Fhe8HEE7M3Z5JwZZ3VF4Hq3xykiGNwbHRfQ
TQA7kmE75ed/9fqSZc5vG/HDTKToO8Nvtv/zi8UzrIQeOp5lwQ4Q+4r9+YX8a9TO
GxVEkschZPhYU4YQt+2M8t4Eb3pfO63dqBEWFFDYc7YFu8JkzfSIEgvYc9mCVoGQ
TAbVOEfDdr6XfseSyWYePrW/EvhSwcfHP2fq6rjjLp/MwiK1rFj7llQ4wuJFLdpL
Fq6vcYqasC0gBllCvEyrigrBgnFI5XFofFgvcHeNAZzO2sUL7yAZeavz4XkBBYEd
+3x/twZyVBMT4IMBWTwfG5HPovBJDnTi7e5h0TgW/QbZlHKxiJSRgRrmUTCSPNmv
W62xhi/hrnhdBuam+3GfkNTuNttMfA2D7jlXuX+fSK/0dRrdax3Dscs1FfQKr0Zl
hjXuf0JV7txuEdJPwP6RGS8OhJ8OxDx50UBjyTzb0uC6Yuwau8y51R58eiRC0jov
mrwkGyEvWaHHbqzKGuNl97KOyrWbq3QFpVfUIZCPB3KuXVQv30IiajlqSI6t1Q9f
qOW99wGaFk38UPJ/gLGdvW9sBp2f2UgKknkm76hTOmrRiA4cipeiA+UW/bd00Cr7
CuCT9IpfkN6BIhy0/o9a3rnspucKP/LHi9e5qeKvnWci3ncpehosGo0wT9YqhO1/
m9PR0OHyL0wbncxhK0jWWj6zWwmH5BL0tPe3ugFwG6sZ6YYKHiT6Goh2tHSlXixP
X+qOsjm3aaHsr9LQF44EtnMaPwSI+KrWcAK8SOMbPXF/FhfqAaSFCEv2JijVxLXL
YsZvpKcDnKIzTan9D8aLE1n6KYwCm11UcE8qwezjyAwLGwizk/8Mz3LtfK3heSfm
EVJOWOR2drxnJGrD7c0CQvuNEQP9ysUPsWK1VBBjzfB8J/CgzGbqH5cXdrNMkAZw
j9gIDAV671GvadlI+GbVIPzR9LX8F/GWbKa2CGPo6iy9i7cJ+9dCK1fkjj6g3yvk
j3h71W7M5/sO4OFY1nofjKl+eGbCwbV591Feg77ODwUnjPY9b6CkvCrxuihZS77n
7D2MYYOkxtjQn7/TG+z9JU2d0Gbs6OooTX4aB9ND+PWmBBACO7sRcmLtzlyARk9p
rOOJ1siI8D4KpLaFYxt1pxZrpjuaqm9PfnRPxhLsfcyzdWvMx8M/xA/R7jtv5hwB
6sKyKjURDextV8rZMV2Gn0ykoCt3vY5WKK7ynWOhvuIQZz8OowbLc7HVjwILWIEp
2swrybEYezrH1CoRvzGfYK+EMnw4rKQwJzz3Hm2jhYIIXYdutFLVC7BbOqx6+FUv
v5P6ct9iSIa7hRmc9qe2UL/MkDgiZ8cbUO0K3riLCYEXMAo9/N69PwTDPkWL0GJo
rEnsmjOeiBbIupxSxfmUCjHAiXF+KZAVCPJGJblj5fupiqSqH0jGwKPK1SjWS31Z
IBLCOhLZH9CE6WLKLbudhmOTF2yW5JHT0ahgoBRnMntw3rZ9QlfIPgbaOH9gYvBx
QgySR5Lzm9IiqBU45eulL5Vheg3XP7ogEn6ed7Om/XeOesdJwCUuUTbUTqvs4vTc
Jm7uJf7Yphnu23ojrtdWYXQkBy2s0HGjY7BvbOoV07I1ypNQhZzIuvDwnuxFNOgA
M5xQeeYZfJe+tnmgDlZqU2W0ZHoAN2KhEc07OtJenn13sjKaVdYkKxVJ00oy25eA
/6moxbFqsy2hxbm2aelg4Qo8fj9TC45egFbryc36bVcAfbnEc2dGW1DUNTUuOGaJ
4phHLQzm5brAQ09C5CPAYwsKuF/kFzMyB2XEHhD8BS62WgXjvxtIbNwWj1ECFu2x
fBS82YI7gev6gGY8wltfv5RLLpLY+t6g+BFbgF7m3s180R0YwknfMPU6D/FoO/b5
iRrDPy9TcprWK5fwXDr+O0obiWHp+kIsMmoKdE9JpUCTBQZb0eJ7vRJ4WMb3Wf22
kbSwHN/jwa/hn2/wRHpQt2JHVAQ8s8vCI3aUOuRjHw0Jr95NYhF1vzs58flAZ2AX
lu096MGzjrMFtt1Lv+6kHwZ9XYuBBPJljJAq6E1emvmDMQtK1UV1Mgng5aDLEvvF
F7IQZf4iK1JSlVU/BQE/LF0wytuNNQH8HngMky9r91tuhELGLmoQt2rm/Lewwxbv
wyX6gb1AkpJNlDmvXWZi8FwgjOxsuAjwiwnt6Q9BYID1UWViVNQrluYSiJcJLC/j
4B4FbcehGTbzOMI3uJVVb3uWUEJ+VdMsIuBz9SB3UOI5rcOQSpvw23c0Y7nNpXFY
aIpwOE5P2PKxD0ubXNriH5a61bbuBImH3/snQ/4LQKFR0raqJV7Hda5rMAcQGFP+
2p6fpW5mxBt6L++xeiD4uvbtZchnuCIc1y3pzYz+/59kzLlSxnIW90JP2mvYibet
/eYYd1tPdUiamtxsnx2iWzcxg1WXu50xKYeBevyouLzoVIxS1Z9aS1BO4RCF9OGz
0y/KTa+uZ6D0mo85EA82hI69SL9NmIIgAmkH2WzrFcs0iMLy/TUO2w2aZP73aycO
tZXr8kW0rC11JSb6P6AGNEJCKNgFXzfu+ZjexDwnIqeM0rfFKCEOBhtPwRiWwJ2z
mMdj821qU0smDh5S4oIBjbsBn2VpebCM74N0AchNRkLejpO7AeCBgY94a8gMJS6J
KdJdavUzUnKp9t3AzfZ4Qr5VVOkV66DNzoaawlsC1SPqCD4EFhiykMGY6F+MkxHA
g5STRq8ccWEczwTf/ryEMjq8ocjQ2fdXW99IFbTZ1zRiuVqXb7m20gUSe4Y3FwFW
iXkSeGQvR7HFfcW/Uh+cdS+Aa3GuSEb78ykbi60XG8XZvGH5zbrqymEY0mr6cQwB
+LX/6/sfnfANacVErDkhyv5ohKVszBLUAznJA6eZcJObQqxUz9qyhV+HCV+Sj5Ov
gngweexHVygqeQHdMDppM+kbYt4UM68/UoJGg0mbaublwXFtf+Ur+czYJGi1VwdI
wFN6Kyi4vBXMsEJ5RM3fCxz6aiKa/6+RTinSywsaYX+0M4X4WVktykf9lZUmSZhK
o4YJlZmW0w8zrJO0AJfrFQMYO8eDPcK6TqbwaTBCeW6NhYnzRC60BErg8EQLfmNF
FRIKKGuiStQharp+AGUCDQi2x7tHhGNjK88Avwc/KTdx6qTtc5OJeZnZqXv/qKwV
KzpzpGZcdlygtylOVTALluQ/EU5fZS0uBbilBm1O6pQn23HrjkKUkfLZ3FbW/RZm
4d4ZZwSTJvAOgtbvdeVdpu7FBq4NepM1qOOUycfxN3bsCvnpUzx3TC9JZpGf4k7a
OOaVo9CV5tfWtxWNCHcncvGFrvJx03f1NbubPj/noVzV8NAZX0BK/B9bLyBkeTmj
rSWAaAqLnoh4UPCANbTD00DQ1X266VqaOIcB0WhBfgfwB7DrJtxTe3lpV5dn9GFd
scrKOsajXrZ3XijuIVl52fqCbGn2bGYpMlzov/uTsZVegHblZtCl76QB22r0mdsL
qN2gSKRydCZyOPLBpgsnBKqU8r690OG4UwHGonlA5zLZf38Fl51UUXd56gsc//ob
7w6vcIT3WFnf/RW/0lB0FGl8ChLUajRMZzr39l4UwNYXiKKm2Kq3uLUtn71NzRe0
awh0tiAJ4xfrky4X2L+GgPRHXzFyOm1JuzI4XiHAYvGbh4ByChJtlg+fhuleEXAx
Ve8Mbmng/BTs+aol8iNuWV9o+HuOPkNBhcJIAtLONt3ReVVBjJ0vt+27P7F8p/83
yzGUMlQIGgPbg7FY+9/H5k5HCJ3xsTDw8cBOAC/jnk2tUn8tMP/o4KB/w+m7VmY7
a9Nky4Qo0VBkAUdLQICdJ8b2/YjUdbsLxR5Kr5wtKWoQDDuhBlk1bBcf5giGvb2N
3/DyNdVrTHe/jXUKIPsVh8K7Q2qebEF38pu/jQlCPv1s27sWvaRoFRpB9lMUJKkp
B/yKuJHKOV5GuU9vKrfiyqW6mWTmrr+NSIWlKIHlv2eBV2yJsEbloVCptHUA/clm
oBbQ+QnnWGgZiAjn2x92Zf3CHfvpMx4jZxGmmqAdLgz7F5nKao4t0/edaLEuxjJ1
qSHUoSIETqIVvLG8IUxSGJjrTdWVK5GYfeAMlnbfqseUQ/KQdCwWR3zjZMZthFb6
ntnB0I3eaGftGdRhRObD7ry2um1+N71l2dZ6QyaaMiK0f4WOK0xnAMzKBDBpgxnG
8Gn0Iw036QXRXO69R+t8oYmFrZruP+9XAlNVfX/P/MwgrLkuToFpF9rbPIntS548
d6kCy/QlEPHiQBE5vZ6vpY7ZjsVVZujPcvFojBCh0qtL63QzAaIHgkzavxPbob0z
FKC8pBVC2FllTG+FC8C0SA5vE9s1nAmWcYTLyNhbEfJjMcdcBRtdKk6xYBudngSl
wn2KDxpAc50YsxY4wVNkpSNvSzeMbXLv8M1LxIFfdQs4XVaLsZW0ect3T6oj6Eeg
yMjDHaC1AlRRDNCLa7ciIIRSO9+p+D/MN9JALJbxTX0bGBsMMhzDtELJJyQrQfwX
wREqjFbfsli69j5CyeSko4YM2J3muBk+qqL111oz3o5oO8Tn3ifoPNve0/EmoRrr
lAVQlt5XVaS0E0xLJCHpCdWZPcMF3Ia6I5wYQAsp3iEe90mJ7kKgpI2M+pAMKcbB
NSUzz5IQzAEjMElAcRB+zusqdrWnbV607/NKhjPkcU32j6SPare1pcyd9R02WSvw
8qOpvQx2UGwUjGzbxN96op10iaw6077fshP0R1D80FlPxBPWFWo3sBtVMwJqK6s2
aYW0V2H3VTF9ox6babni0rILGUlcUp5kLs+INYwwa3HiQgPVHXfq2CBsFiUlI8gB
viY++lL45HyCnnudfZOWKhbEMM0ipT6Wtqj9tOcaC0gz/98cDqV+yeY8hiDvhqBs
gHxbZ0QYpRDMH2XSvlmSDtnBd3xVuD2wXna05WC3YAgLO96Vqb7RsmBEOGP+7g3i
H2UZlzkX+kjMlZ4Hm2ZHn+2sEwopFHwb9EyaHxjbUDwUvp9VmyUBcTYmQkk0dLBU
Y/iM858QXCwylIiFrTLH0BiPpRMT8VUH3kEn6ETCigpkZvYMOlg3E4bw/crHi3KG
RlN5tTEM3/m8hFm8CbtA8M1WMcJNoBtMjMFQqQBrfWvR+A5tGDNiLvELSvMX4o1g
ySCtkkLao2hZRQCBYegmk7gyDCNo/64TUpH08J/8yTPdA5qD3Xzl/1g8+zlAS6/K
toMeKqkOdwd2Ft89afxiUFjTmWxiOSzUrhhlsd/WRP6ZXOTQflN57/eotrAClx1R
5CagpMkO7qDxuNBS5sVYf5YEfO7SmLA35e3KEHjmom+K4BQ7RZdtlemPFrL2ZdCb
/KoH2fx5RN4x8e9p0t+hL4W8e8LTr2a9ng6ygDMOpheYUuGRKCVD+90MqjWdKvWH
hGyVpzJvunK2RDaX/AHXWsqp0f7zb1+2KCKwmLarVwNi8CGEiETUm1iLyaUi/5z6
SVBlQxRm9Oa34xcTOPORSd0tZ8bhwHlblGPIsUOh8fK3mZRF4iTgP2lt8vz6gqaA
Ojp+h1/3C2Y/aPNs/vsSZGAjpEzyd50Vtw5jNboTHc4ssMfcntiigRoDg/F5gk7B
wCRjoViX3GfMztBsYpm1cb6uPhQMEoSjjTw01QFIRepZWqWDFRZ7nSZjBC2rlrkp
hkAw5/54D8KPPPMIK9/jzoH1Cz+kdyHqEV83SewnyxM3Ce9TW/EneWNjgbk1Y+r/
E1qO5Hiu/qkqtuSMl+kV9XUkX458Vun5igWlaVYvaePKF+BxBpjpGAIrOVkF+89h
0Mf3wE5xnbejdQDFgHx5G1Luz0iqdiysRCUCg5s/7h/TQtA3FouOoy3zsGLuxBfs
BDuGUIkZJi2iLW0AQXefQaRyOGxGDWbToHhW6EpI24JovVhLIhO67hYB3CaMIHJe
tj/25izF+BwDHtU5y3xJyc/n4+IpB2fbZdbdcym29LNVuC6SwbbXOb7kEAlw2rUh
agmP6dk1EE6Ju/eVYSL5V1p0ZwfYyTBtJWxq28ettcvMOx7gewhFdtLdaM+Y/75X
EUd+j6gmve/71ZKZzxBLUof9cAwnUAfuxnaitGsUTfzOn1DFcA2ZQKcitONND41z
vhq8MX1Hr9KO+UTgE7wgpZ50F6kSNM3CB0az6jE0tGDNvyPkn4ziJBqcAL6XITsO
9GaRq1nLP4s7WcGIhrusyIMX0lF82tTYlw/8ACYUNcYWWwCEqepViIjTpa5jBrm7
YEISg29nbS6VxvWKcp5anE94n8MertuZQxMxII65BmWVAIHkHsDGt1BkwQgbwxke
NKrE+yuT+b86vDL3C+FpHabXv7exXd3BvXNaJFzNxzODsTF2OkAI/b9Zi672Sbx3
myWrj+qz+HaDCqOhM8tIM08dt+c/DMRNa8GAVWN676IN3YzN18VlSfFxZD8QkxbB
MuFjHnszjJG8GYPPi1ZNd4LcC1gvrVWMseD/OpJdTO437nNYqE47N2s8Nm2ebhFz
gXcJnmYNkHk71F8vejb2O1MJu6NIEd7iK7qyn56hxKEaQbSK2bGUKGYcnUvK88Iu
tKXEo/MwzrZ4Dq/q5oHlC9j/DDSWoso+Scyc50YbsLub5Z5GucwTpcwwmsaaXdfV
CLzsPFh2m/tftAgfa1jBr/zDr0L8ONyszhXR7EX1bI3dHfSM3ocrN8J32YIe+eye
ZK+iK72uegR717jnTrHQbtznTuP/By5ZmL/E/rdoM2h1ITuzuLnBE0BbBh990R37
VXfXrNcKtzE8ZA3tGdT61vsOZccUC9IhF7uJDDoS28ULn0iBLLdD6nhzYrEAqY0V
86TIk7utjcwxSPLn7AoM817vr01AhH8EMzzJ9fZb3GCvPvjFT0qi8/JYS69Xnx8L
Vsu2oPiUHLYcI6niPwh7p7yCtYudhnXe1TsUFCRWllLuaJADLtv4Vb8cj6xgeA8q
4BqcJOCGtdHhcenPPF5qi+l9hdeNcj8SApkULIQZTDGfCcifJkW/DWLoPK5Mi5R4
nC13YCNUqx/IdL+MBR0ITqzTJ8e0sZNLohhQIBbCWYZ681pW8xGmTdi5klvEApYR
Xq3BrV5G8WviKLk3It4jE7LUA8OFAvqNRJuwRIpZyjhXb7Qi612ld2PMkcujxszJ
5EtjXYpUApUutAz+Pd0VkJl6PVEM3ClY/vIndZMgOUBMiBxJyljOkB1qQAFubZKx
GZ2Leg08qd6/7sr+7Hh2ZEP3fW5F2dlr9wshHfErWipTsIsWijrEGIJkOQeBnpcq
pFxOsS4VWiMNB4tXaK4eZCEJZXI8Es3sxuEkTrkT3SNwKYvN3+/l8z8vOcDLILMc
Of5j6XOs6dM3iMx90myBuQKHDgIe0hIrHQvDfBsz1nn2UbhrNc8EulwzvnDDngOJ
mJ7MGMD+OWZRN8UFA2Etydnj918y+5tPJxMNHaNnlcyosmyTS1j7tMpE34bl/Yb6
EpHWdDusgDUvzQombSTD3FQBIuOXfjKKolnfusmb9oWE19q2EIWSCOu3OjHAyWnK
Vnvuif/UQnSC/Db/028S+q5jBEdLJ6Z3y5de0Gk6Yjnuriv/lq/5H0c1GcQ5tLNX
6Qk8EpiyElQGjy0zePmwZ72nb36h1OLMTC/kO4/lP1PMHGiDOXYM0LaSY6cJUrT8
wzGz8NKv8M+tps2eD1XYRNuxJFheuIedVorSSGyvpQaFKRpeuwlVpV4kLAtYyVCF
Pge9Vma6aMeGMp18UWoGJwNpxuEjyia1bH7IFFRbuWpavmjnhsSylfHSKlIUl+/E
ZoQYjOa/gmRkTj1QHDUPmWBaEUlqkz6l+NYzip8hRIgM+U3p3cijNE8KSE7blQN3
w4zACQbMqDfOhGKr/j4QLBWfV8+lyas4HnQIN5trur3aokTRxVVOF5pPdP/02TVJ
/p7+mM2xwMF+AMpjzAIM6SDZ6tcqcpsAl+tE5CNQaeme7IHNjOVP1+0WXMYl3x7v
ompe5uFBabKMBmPdSh+j9AFfVAFFLCZ0pIGZpIb/uwi3Imtp3SXqmqMkOFMrqwNY
JDCahm530na3kAvlZWuJR57JssDIInA+PLcCTeRgCPyUUDv5G1hDyF8b+Pybveuq
Vkg3GjOCEwL1Bkm0WOt7Az9yL/hsBehdMsetC4/SBPciSVv/zD8QycufYxNfi72K
Z6ZBCRO1KkbSJ+u1swoWZ8sXkWC7JUlGgGjXUAr6EQ/oUlu2t36kP/9VeNSWMm4x
BsgOinS3qrRanA2EPIOX7rKj0p99m9MN4GcfFFSI/fpSMkivh8Qzn8MZiMWgmP0j
QQp8/JUosiBGpC2aJ9Uf8oWYPOiRiCdCXHsCCrMQs9txqF8YySNppVBgxeJutwAY
aIV7z41cjkpl78e2pE3jyKM1vYgN9/zZrN2Ilghhy/KCeU+LfwBcgxJUagntCF0t
MuXBjubroxcYZY0FeqI86hdy0obFFWDCN1/62f1AjH+3VuA8mpHfCx5Y47jfJy8w
pvDW7IIehKDInUwbTqVsDHGiGCtF7uOUD13mutxr7I/K5P9+4u0FfTFdl1EBdmZD
M2ZiIn9HaLneNj5Z8J/vjci4BB/T3fBJOhqfOX+J5tnp+WKYKvnmcg6e5F4YWWmp
SRCJJhY1NPXF7yWToEQXkrfNkdXGUXm16Z+eEvAdSppbH85uvqSaHsGkn/ZA/EMV
xjWzYtEQbPi5W7Z/25oorGzPqkph0N1AaFgrlR27KgS7hLaUhQ1DYFH/0mEtFohH
4irAJS+tuEYxkqa+bHR8csjKy+7l0dR85ALPvnds//XypBfccTNM3aEG4Gsw9+DW
fgL3T7vRvHMhVJtX+f3Xwdx3R+13NJIj1tSet7IdD+DDUtpEGwdHJQF73s2pJYO+
kWm0TwlQ8P+Hlaup9LD8a7pPokogVyfXdqpXuN3gV7HbquGVIHlo1aFYMytEmaM+
M2JtYGu1r50+SD3lSkVTMFxIYVbZCMlGONXzmis0Lllyzqym8OAftVJLl7gnqMmx
PxWTPmH84nZ9SRIJRRdRIzPu7xewCdqlWFSfiiyqbMJAPdZ88TMHBZrV3yHl5BwN
hoD4pbQJk3HO1HaO5w3pdvqzFVtXyge79ZAuJ+eMeiLhJeZMSIdBwcLR7HQ4dnq5
Kr5zzK77gp4/P3WT1694X7vZVIr5jaRbdtdC/3JidzptDR5UO/wwoIVGRSp1SDQL
p7BwiyqRr+y5DaEbsJRRwyEI3E4Xr3Ri0j9VVmXr7h73vqrNrzRUELhs0CasPVBj
jO5O18uj9RMVZgEZC52NpZmPh9+KsuqMag+X2WO1NeQe46vM0PUAI7vhxWE9mOTZ
iJqxUwpqzgGSrkwRCj9ciULWIsRJj8ZoAPLEotn/3P6qNf8KcH+Kq6HSCnxqzukA
7XiKHpIA4MBOw44y/j3nmugY0Yv+gWE8+w6FXXHB1gs5YouuKNxpVfNEmMlcJ3sa
8h8/ZrJeHiueLRPr1tFA9cZeM0lUjgIyDaAO2CVaYHL5SknzU1a003dxRJioSz5F
tLBBjzRUrAMYjtJL8nhSkCZO68hdEpooDfD2Fwz6GXbtqe7ArwztsZIwjREARYae
3R0/0Y9+L34kkQlvyGJ2rugCp81CGV65/IX9RYOS85HT+mxjNC7Eyk0qhmgdaUQi
NBt1lOBll253wYUS8IJlyKo9OBn/yXa66netOGrIZ6RInejcDZP7+RL49OCA3xe7
JJp8dHY2SyVtQ4ZqEAb8R2NYlp8xvLIdsnZ4H6P6lsJRfMekOlSjy41cas91CXT5
qwHnrhSKqIqtoQEOcKU8iFwcTV6uFnPf0AIG3UooYxAKHp+7DPNDfH3QoB62YmHg
BCUHJjaOdeHe8jbZchbSvd6fE0F0Gr31jeNj8bMzaAihrK82JP1drPaFerzxVToH
gabg1oFh7wwBHLCefbheVHRxZ/fqchQ39N50lYWQ2HQRrmwRPdDezYFn55+OafTL
J/N9e1tU+3058puSKGwGPdwaxcWMjpdCICP+ThRKIsi7f9YygRZGA8KuF8VMYjdL
QLHwtP1Ay0fmVl5bJiL3F2bBH78EH9t13Se9hOUR645H0Tcif81uUihl7Jg2YKTR
tsaAkH5C8QzscOgGSZlWkOw/U+LnjTtSyNri15/ebEIN22IMt2pA4m+NYX4pvOu/
H3HNdywmVPYa8kVRq9tNDTwm2+MfiBHVKb+ytbUTJmv3EiVa1kKKxQ3bR70r28tO
XsQEY6dEHtD0AIq5SI5cgBlCgsGJ10hrc7jQwpsaMMq7cU4C1oA2irR0nS7mXj7F
j73dBBG6LZ/NZpTlRriq9yw8MWs2OMVdhr4O0GVJ+brInB86lpT6MYXbh7FFnmr6
8YLNsQIOMh5MxT6el2fgiRzq2FdccoSGsBz53AyhlhFSnvRjiWCfa7tKlNTJiUSK
elmabjDNGp/NNKdyJL+KFpm9iPUW8z1F7LxucdPWi0DdrO5JW8YTdU+J8zBK7Mo1
j/5ItSrfJ/F7jHn5tv9hDcBSJbLXXS/75FUKLzKh0eLPwipE4TAuWztmN4eAuoIk
NY9QpgqGZCbNWzgs6Cuf1Jlqh/EAYF7sD/yMo1JC1Rnxgd3qV0Gmpt4s//8x7xbi
wNRmvoK4KyRj56K0RSW38HuWVLGo3udF7h4sB3BJqKnA+hCr+Id/kpQ2Co1peZfA
ePqLrkLsz4CHIt1Pa7h60fwwbuZmWNOLhJXM5aMKozGRtuhSbZkIBUdueop92AMw
2IGr2UawMvzg4HOZIn57BMjj/vNzMpD9h80fzMwI9hTTG2+ffh1Tg7PigtlYzquC
C19ZKFRtJc53gFKt8fyaXN+ic1vtghrATKnkMVXHpG56wceDCxRqIflj8S3yBBN+
zq5rHLYeFy58VQDKL9b+dsicTkH/KSwruJOvLNo5i03XUYPlqZZlHIAb0ro9fYUR
ypUi0sGXLAingt1aths/bTGH8LlwShADpf4kz2dYFIFFlU/g1o6l2gELVB17w7P5
4CFay+ooHoiZ+amSSFAiwPm5huA5Z53jxNmXWXQ0mczBuRaJlNmeXy1A3UeOZl1s
XDoPZniYmlKlnnE1hcWruN/dEXog0h2w3VhXxclaxQ6+JYkGbxjqSkAtLsTT0bca
Ig2PeBqdLmyZTLSUrRMRI01rOkBEBupFt4lZUZrzq7aT93Jy5fxkKbS6TzBhmw12
GHnXTcqEim3Z6fpaJnwvho83H53YqcOyBJk+3Ok/fX3n0YnFm9P6uqdeB2rDbznG
ZZMsz7ZxDAjU/ynFzKeJDppePC1gudkSvZ3Np/nYfQUPlTMj9ObxFhlqO+Pz76Pa
GY9sx32FdaBViwGornrUMLR9hTqFsjYUxFZIJEejXbDf88KgNki2gxLY4QGFGZ1R
c2KcWhpdSQDIyPcmKHSkvnkVbdd6ymvEC7ull3mmlS+a+uWuSKmiXTJAkVh3L08X
1FQDKYZ+WFsTpgZnDlzNINoRhej97Zfog3df32kZo8d026s9uZP6OwIIq8090LSb
c9geh8JgDG052XIJBU82zJ/OUZqIiP2n3sKt1mG33tZfGpki3r5geO9jTwNnb5K1
qrGtgTs7JiWq9AjSO/NXZUty38GrbM9DmOvsf9uql/5sx0PfbTc2zugA9v48J2j/
IayfqofK+pAjEr31j+plL3uausV0SWmt5rHvr0c30EWU3KrCGo++Y857FH/tD+Km
Ay+DkdzBC5ApFBt6T77192wDaHFT0Gmbcj0vaAMRc3vn2VV8ml0n28GGkCBrVyRE
Ks/Huz2GOhRLHMb6TgJpEQq/DqcxB/cDhCy+vxb+BcTn3RAtA8ZUz1bGApwY2N/o
jZtAEmd1I/7ZCNf2eGRpE4WH0CzcRvA5XJECk1Dm8GM9gfx12p2jGnjs+vGhOoka
83d8f/TzaIHobyWkgI4Rww8YFQs37LcF1Ve8CgX1f9rcPBSKYvJdqVLgTpj6nbJg
eqUazUtuCevc6Ori/Gk8c+agMrfGGbOnR2V5BXCTDqwVrQ8mDAb+paL29WdA+eea
lC47mD0Nh4E5p/nXqbGpB/MxLzPtScBgPmgT1A+YCv0CZLFV88KDACf49y28d769
MXBjcSaj0qbpuQTjANbSFXh9yxgIj9lSoWTRSpRc8UGtYjBbZaNrrHmm4NjaZsrd
ctW/ePLcxekYO2QXSgRKlc+BfSUdPWCGcUD4Vqx37I5AYytu/hwtcuovt0ukXsHI
cT7zUBfpPy1Ml0zbztZF1faYD2IlONck4gObSli2v+mv9gh9B8JlV46pkknHJGRP
zyjaTXm8+iyI3sUmdRoF5xG/D6ZApbxQtr8q4IPA9pFYTETQvdH8epF77gHYjyib
C2c3gRsC0Jvfs3fZEGW+95VrlViKwV2MAwLQTRIV3+O80adXq9lT4tY2DUHpdCeL
+bokRBcKnvNpSXvLEd410UMnZI9dvZuNKOJPyi6OwXM+XEg1ZkH+7Q/hXV6v0CIe
XG5N3wjohrQFfmyFaybkBbri4EGzJt7bH+Q44NFu834BPTmao7yfc242WCme2LsZ
2M3aucm8BdARQ2EVSwGxnjT90qvQjNbmYSPCRgEsGK4eGSge2eEAX/0vT/fwMrph
Fm/K3RPGv7Ct35keRDi6L3o6AkFwRsL3Ybpa9XPU4e73yepVCY5YgSt8xsYHN7Z9
uojYC5XWSFWpz3Pre6zM+nDV/msNOdBLD3a/yuvdkQAujwiW+QuwTlG1Hs1s2ZdM
/dK+zts6P1wgXT50d7hKNElsrwvv61WnjyavSkCBPE40KgSpG11WqlM7URisLcGG
zg5gHwnawzdM8Y2/LB6z5IzHxA/IaFUSd9UY38BPgPzO7cfNDKAY1kZGkc66f8uG
XkohLPL9K8yyJoXy2R6WdQRT5G5E9BDAGvNF8mDVd+V2Z3Qi50LYY5MlCouf2sOO
UibsEF/7jU0eSd0qk7WoLoNlzxTIy2Xvu9vwCPXB4MAOzZ+1HdZfDNQwHRnV5LhL
CYEgEHkzz8bhV6uA857CPjquEFiQvqfWDnGfSECYPn+N5DYr3yx4WC8nrbCK17/U
CUkNQlAhw4sXtLv7FOS0uohYCijmF0+qAM13frVnMnO0oVz20YgUavi2uxYz0oZb
XfF3v26366Dqcr6HFtIn+W7TF1wLC3spNan5+D8DIT4F7eZcG5X1vNweobWjwe6P
hldflzfymE7zvuBHnkUDg2U6aGQlTkO5fBXHOf+UAwTSgwW9wBACOtJDaq7oRFdg
eey8Ex9ovuNFQqpHwMCR79ABgMVQT0090aP5na9hKnPfj47Pc0iWBN3ApqFHORLa
DA4VzWk2RG8v7cRT4fEPmhdXRVWq/0GCF9FcSnvLfhaQUSwjmXMcMaA1TPkU2T1b
l2qfnUh1VlnQZsWpJKisSEyeCjIffNC1D8BZteS99Byqi6DcfQE5rziaDGMGqwvv
mvkk4SZ8h1AAPo1CawUWE6GZ8XRy4PJTpSygBxg0XBkTfqWtM0ZbNGz95gRqCITw
2uHZ2rClbNJRWx9nGksXTab2r4XkmmwqFBBewkKMjeKPsuln2DKb/ZN8WKB+W5NJ
BNB2OPfGWGiyawfo7tgeeD1Wxk0Bt9o5nmO4T83MiPa7odvu9n/L1a7mW0Dxct9w
DpX+OgvG+tAurcRUgTR/WMw82jCKnV8mfdyHoCwOkVhPbFvURxVoO1QbxWKG/dHL
j5Dwcu1fOBH5JaQ2DDtDttdwIKYEo6PHfmo0OkRhw8Vrz1kK6oIyD9eF+P1EPana
Bl8pnmcWvi3S+cyedsg4RshJBAF4EpEx+w7LrpxzXvlbLyif4no33QqKYpfp/wUk
36J8Sd2TP0glGbo1mKWfrKj+Y3knykkYVhE0f2l05jI0qa27vGn+d428HAJQJsNZ
B7AVRHLqJ5LVtl0osBY+7UfqGPpR5F0M8TIvlHfXUPIjZ7+dk4cOWMKjKYjY/98I
DTK5inhLAlXWBhY7wfJqq6he0+sJXOaiys3wqXHF+A8Ki2xLEH/I4Bhmtdhcedc1
fwFRWkrOA0NNYheuazxmtp+VrQ2QdJewE7aDAFTsNAbTn80v/A/Wb/CHlNfi5xzW
xpvOGJLjNbQlrsK00rkWTkjaJ0kDOhvUjuPhfTybDa2RkI4MRQ//4ol5fFSaDFCo
NsTeRpWCjiNTv7L1LXVkrjjXhgWF1/yn3DLItvouh4WfxJ1ES5CSOzMbnR1q3iZX
F0pgan9mQ1VPB6HtvD6hY8zM3MarJ9ZtAtGAnQ+X28l6ho5i0mYdBf5SF8686NGu
ulFwWzx0l376WWexBqwcHWA0n2WCAUDFlx6cwOozVn/S+hgAGahWhnTvwGSYFyR6
cL8gZrNA8eMdx/npaI/ZfiKuTvt5uDdme2We+9yaZYEAAvUJKhb+nk/rVNjTw40x
9pt7Kjkk597ImRrXafHIG2dzoBxPggpZO7JWjibV7LrrjqCTTV36gCoLedcndgkh
vQeWpHcjjgdZfRWzXpe7DoBcUSoN8YULKQfDQ+FWaNWfB80w9Nn2/yEP7UCLtL2g
5b9piaZ5c7ItmPzE/B4s7Eh1k3S3zkihrl23HB0oR97Qn0PHYnySSBe3OIMBlITU
0O55CmyW5NHPC/fhfIOYBdhoj2N9VuES143AYifFe+zIVc3cvSD5vTlGyRdQ9hbH
Ias9Wwnbp6eHA1+rwLH3ALIqUpnQgXPsSTgeqe1BkHBIhzSJpA/82DF/p0pwbkr7
JdjXV6MxAPXJGmuSTtRkNaxapSVHqTvvoqMgsUF5wzcBF2noh1fsz1h3xPUXuhdv
WqNq7mN6yWds1XXLysMwPShTnLvAMRn7j432EgHU+O8yboWxM7LN2R42J3RFj7WT
aFPDy6WhX2faPbxo0o1VG2u7i4ugMSvvaYK0asrp4iFPZtIDKh6arG6QkJY2kezl
cxTuAornehxx3UOU/YFqvuKfZfGpM9dI3JIXS7SOiLE4XUZ11ynszMAgVdG/xv82
fGQQXmTaM1dTZawGsB4hzTZRdNdwG2FoAMxxka9NzeUhlv/JQp3NOUxAqqcXFBKW
L0vupNo1ePWqVOPJ7h1yNqaMwl5eYymN9JfYAXBoDxauP8T4OpzuibcUKYz1cYlt
CB5uov6t6n8UbmJPnRWC4BbqpgyU9VTMMDId6gpZXm8o7Mi5pqD5AckkEjTuHEjD
YCaP/4JzxZwsLOOCZXoHNnMBak2FyM47IuJ1ANfwdiwNYcpKvuGUQd9zdw/a5xTf
GyyH/jTC/gov92LuHZR4o9ZDB4b+beYhaST5CauZ/qubJz/pMZ8RF4XK8CkWNU0+
oa0NuNIkGQfyaLzJaSjIfwLLGXSWj25KW0jIlHd3F8KxHoz0Ht/QAah8OMLpMsXf
/1VnagiCSCvEI8AbktVbJVoKLpvn1Xs8LKEA91RAs1IafX41FtEvgjuyykGxw/2F
OpgPGJhmEqxs0syKWrf69JZvh8zqtsufR8x/PQHY1w97ykFd6SIaOW0RojByDA5T
ujrtaBeN2He/gAR6L3/WbsmSbz3XyZUGYxMun/Hboxqc8FpprwIRuZrmVx7uBwaU
sLVSfgqQ00hDxYoMhcgOv8oSF5skCvflUclB58jv8PQvgUtM1j8ClAH8uH+P9l4w
7LhxShPeQ111njQCSGReBQT6jEZQ8RV2FMpRQkLM8IboARteeY4NAxdcGvShc96H
73+7nMgbF6+nRie7Ddg/r6vnddor8eHstSYX0FdlFmMlPrKWhr5W3Dq9H6Re6YaB
OIutQQFbKCf9oZkXFbm8KMsTPW/h2DNLNCVl2+aTHagE4q64Jetys7lCuLCW8N14
cGzLvdEBq0Z3xMRW/bSohMJITdcVU4H2HgB4jphB3WcGlrYxenj2mRP2z1ivZZt+
maLE9QoqruH9B/M0+q0KRj/ra3b7psO43tWkA0XwlMo+EbOhp4ACa3wUpwsiSroP
+420UdCFfjnn2L7NfzPQDVm3tqYNB/g1dXZtjFGLgJQtBZ1i2ErYkFRGDx3YjlWC
NviNl9WIFrWIVrpfoDqFUwcmcjOQe/lvXwbyxhop5sbGVw388O4BxLDeVQLYNBM8
x/Ko5BOSmQXn2sf56gBd74/aCeE+G4cwyUHC3tnrXBPSRnSp28jb4Pc8loZ7PIVm
a+XPbub4/WcA/SjKffHw9e/DkYPJLTAh2qv9woInD1QpFJ6FDhJ3fETRcUeRLCVH
PA/bllnxOppquaVejKrbCuCkkY1cx2IjaYwlCU8DKOQvkvOhxoxCjBZugd83Si/P
3CvqXi6n19frFkigkxaYveb4m5qYqKCJyV+XkVvBYqO+XfMND/HA/UeUNcrJyk7l
43c/U8I/cxnRl7uFJA+D44dIuEcGyXL1Blk5VefO4Uc2kHKtfoxyQMGf9ZFbtPjd
juhcq02FeidFT7eYGpJY4zSq9tw9JAt0EnmwYlYwBvKMvwMMTGMX06/vAcFjzi3k
WUNoSw8aqALr7EjX94r359IHDeewDYyMIUHvxOJr5fmrZzVkgLdqps4F1fVqYfw7
2p6AJSSAtS6bsOt8p20VOfgBqRWIbBH+Kqr5IMonKnxCmWY9jk28AVMn7AeoDpc2
MlJe/skB6HLbbevEVTHQFIFYEeEMQv2Q7bQgdmVQYZPLJAcK4liMs5/uCJTRno+l
u1WqkrBJ2EHyGzUIls/FkGAOPJNZ+v+YdneCtwCg6L3UiaQtq6QAaeytFYURuPC9
mGKVz3UQ85Y50DaxXx7gC3wEPnnjAuCkZ3rkbVVQMy8ZKo96LnzeVC5gpORR9/Ll
vjGyDFYWA2I3FNn1NkQwk+jBm+BvCNvc00awyZvARYV6YjtDvj0VI68x8k1heiMD
f6AHpQumiyzDIB9EKf/FJwFucdmDNKv00aSk1W9Dx0ErEdDFSzTHb6tp0MsHlph7
/HlJFR7TXl8ARkXPFJm7k1DidMT6RtTdAllsimFLsJvmh0iKt5oZnEo+ggIE4L+t
dZBljKYdYBvAgiQVtrKfIUGIZny1sQTxykmPo+PN1JNNxq79uVW//3kiZnWIF27y
oww1ItFVL7PgTH0lJrlozz+QI9dExg0UTBYuB3SXB2vPOWUDtDDuktGjOlq5Xn1K
Al0s34+38DoUr2TPd4/waetsPWqkTHepmoZI+0IpKLVVf1TjQrI4TSvNFDBEfviY
WOnZgR2HI6mS78z4ULGTO7vQ5nZLDHRIImLO/AItbB7JoFMtFqq1ShjvncPwkEp4
GpuVIT+lbuw4aJtBm2zt7Vjw54VNutlDGDgsovEc978IsmrPHL3vB5bpYQTzVXhq
0VsIw2WzxHRP6RYwQkbK6ohMJQtyQNub8w0S2hl39gULmSmi6l4DbQmazptV8Lqt
rJ5HIvynxVpdbQ92WmFWcpPqzD6V/Wu6VUKJpi8knU2zpCBNRy4nsN6f1GxvcJeR
DQU9LKE4d+tN2N7W+SVJJhCS79ygUbfcm5TCNzh10mTQHU1EfqNpPbuAyz2gdrZY
b2olbXu5kNy/HqVjdLkK98in+nWeH/gf0jYAuNMwKW55EvX+Pzu5jI/1UGdftzs3
tKPfINwnzXjxcZL8FPPc6dCt0cuODP9Sf1sts3xtADfk2wPFvBw3T5tuO5x8M/UU
NfQrl+CHEoV6VMRViyv8I/18nlIq9xcUlrKr42lPOqw3caTY2ZMcfRcM9Utq7RiF
AX+iTSZ6RYDI8Q6YU+ChdjtTWk5jiSw0nn8lx8pJRsn3TFranAG1TMVxQ8N3Pq5a
Ut23M8xnM8dHBG/+KTzb1xFTcxkCITLLKL098mTmbpnreeU1Os61UUXeXsen2wiC
oMupdjkJIkv/39QDPC8Ea6oFaFUZ+v/8KAniyQL4GVhgL1nmz3XIEa0g9SrIX8du
8zJ0SYtM2TNAPF00LK8iSmntFUR+Q1OVHMFkE/AzqAnWdsZYRPoEm/f+RdYg0+W3
LovkngsAeOTNvLwsGVGofrIkZ0wyc/v7I74tFEu+0/TZfz9MO5U/C+T6aeqetQxy
g5xdkXO3vhjF6Itdawc4joqdg30/HhEhj6cYZjJrE72oO5u6/ptbSQhLhV241tf3
6aZnp5j/0s3x6OyxVYI+bwQU0Hia9iWGn6Y0HZXGvs8h4dnVZ20nnVZkBXbQLKqj
PayTJaku1s2NIxm9I8DZQQVmjoPUyolxlls5ju6S9OeuuLuVItynNLyuz3Io403d
eEYZlFq7lxKz5eQ2OnxRyVS3fvOxTmY62GqZXmwtogilEpDs4L8oLWyzyHZPu32d
l+hk1bexYQlm+PK72g+khE5daV0qlGTHvsrdv3BaNjVFgrIsrT9tEEuDQp8fA4JE
qpd3+AjU/LsLfiZM39Dv0bjA2PWF4rTDqiGs6PWvdOHPld/sLJQ4y9LLNCFRslWn
fNvpeZjeMjJkgNLPxIuh3079A+GgrUUudgKvDCGi4YU57uhMyCNQaWsVTaZV/qsm
WngjIG3Tavv6Vb+yfmv0Y9wyYIYxFphWV3drKH9OS6kTGMEy8Y2ujGC7q43WxPWB
HCmveDBDJksoLuaUkG2W+pT3X3om2MTpCQUqpQNqSvI6OIuBe6to5NYeWiBBv0bK
dJUzGXn1JIcDicFRMnEnROPYa/IW+xT1IGWWaMeNVn28EB8TLvV6ezN8RLFoG4Yp
rliuHO/2vqGMu5WpNDutNGiL40qPkNpGy8bRH7HTijdW4PRxHcvedUyh+V2soKAv
ZLAAAmFMYD3cbqSVoIb2n4auIGhR90KzVOnvG07wbgjTQh/4OrW3kHTmSgmymkz6
/Z93pDAoBms6MAaCBsnhqe0j1tujqU6h5a96lPhQw6VgTungFD6t0XRr92Hokkiz
OMp11ngxDtN9NHZAoIVhdO/iQ2RZX49WixC4qS3PegCPZSc6PC+maniss7Hf0OU1
k7wvDBYH8NYZ6i+bfGbvILCBr1Mjn3yezBbAcDFii1vFo66uoGhNuCGfaecAUMCK
OJVc/Ag6RP8GpWR5HgWGco6FDPHlB5viv/V4b+b09JDmMRhnWVMd+4+ikZSLEh7c
yVhTzaDElcKVvkXq1rAyEwhv/Sj8CHIscsUYhKBMsnkWrHFBg1qwrp/HDMlipvZ+
XC3yLCZOGChQLln2tMz/obrvYBVJBUt+/9aJnJ36651KLrFsS6gVYSLXI9adJGoe
oW5y1tmVPNWGlGKHZ/KoqDHPxUzfO5zHmGHKbqDGzi7mEh9NMlATqIYDPAdN979B
QNBFTKnZsff6XIpw+Ztmd1kgvZd5sPNncSY9xiplb1qusI+MpLjBQeXm2WDZqn+V
OxW5WD96zg/qmhgoItXdZ9ETVLaU9IX/pXqzzx/P70P7Z9D3O0KtMZ5cK8VfacrB
sbnEV4Tl85O53RVErFjPBE92hmpBLpZpyE27QE8N5PC0eUsGIOnEkhuU7RODa5mT
Gxue1EIN/vWQpItZ2jnrWYyOhHc9gtyigWPy+7O15c4hurbefw9Pho3TPScHngOs
I605uA4qQ1ukpXrP3QibkfdTyXLverrQOzjIJp/AxGIjkitoraw6v3SYjQzhBhW0
gHLAkiEw+p/Vvdf8hchN9Ts7+be1C8BdL2PlJUjF3YktQZHAkHmIbc21qRYJV4n+
5XqYJiVhg7kon0hM6QrA9z16M+g9mZJ84RghmFL/rkAP2QdnKX0pzqyKu+2PgAxQ
tQV+CsytM7TBpNtBPNNZ+zOfICdeQl7BOr6w48aZZVOpNIydqsDCfv62vs8rRy9h
9/MIYvRHRkFZdWRxrDGMJDaEnxm1lGCxOk6LPVHyfjoue5rxAJiMfkosCHSzpSEh
uvJsMLqL65y9OUDs0NQZHeyQoRpHay9bjNIvgN6uD06Y4iXk2dbBI057aB7aBtlb
f8NtIxPiZ2vUKCe9VuiFWLRWrLWTrALURXZOG0yKBFOffu44Ra/0VmZNHFKw1Cv7
BAnG8NubOEAhBvR0FtrUseI2r59QQwrkFG5B22TZoDzNKr15GG+S3t32kjlzOW32
XrvGZkwtKK2lVG+uqVg71165WwrLrzs8oZGQIwBPzbp5c8QkO0L4TJnph2G7MCMt
7kFwHyu6fCea+bXt2W7Y7eDZdQaq19mjU9mWVEt10OPsEPJt0+2JE4Kcj/4TMpk6
7MdENp0m09zTfbNpnHyI3fRsCUq7l5gJ+FBVAB8sJSU2S2LKzi6vhW2D0Jz1nu9w
i16IQdKfus+xKMtkbfDu4OzG02lQ9xlzihxvba5ryqHAn70Z5d+tQ1gT5xN8iK2d
/8ssvP8YU9U/RgvJtOEyOv2T5Y1HBO2OKHVjD0I3vWvKlNG89e5CBZyxcBCsLRRp
zsGEiWx+a5SWL51jtvPQpMszUzbOS9Cxfqv7d18aVCOf9xGIt+c6P7U/PXVBo/tl
yZngPaM5yHGhynHtT94YX7uFAVoWceD4NtP3Wf7sTk++0iWD4/QHWOp/SqzP1AVK
4qzcEI75IeIjkx8bDURXDf4Iqvnp//0l4/FSwf6fusDDzsFjdPfxuhh5DoxTYeQ1
fzdSngshTWMW+Prssekw2q5/FqKH0tZp0x4Z7/2IAdCfcuI4xh1tLibCFIZR7YIb
6VFYgeQsi9Gb2js4WbdrMj78p6lMP/1p6J+8zEGmPZKn/BQnRUXhVjjBbsbDHify
QVtFOJonacmWz8K9EmCdeYfu9/CAot0uHjPEvs9V4+GcdoKsfeCH5rtc/tNEsEIp
rBZ3FR233OSxIm1qls07evyueyijQn9UG9Lclbaad6xTM/oI6z3LETIFMsK6AkpS
d4GxM7nmZwfonNgy+egzVuj7g1+oy1REmFGFLnRImdp6ZFyQiF0eVCVGdfDPr9bE
sqy/fYsoqvJ/8p1y9sUbDWrqPTvrFB+XJe08w+pjURduEw5mrh/HFjvuuvh6UeRh
dztVJqa6FT5XHMyUROWcltSzsUY4TOnL/ed1QJ0ZGzJUvv91KUWLSQeKLrSCqVzG
wT9BPAlUx9cigP/Qw/8efnqcPrx3bSwlsAQ4JjWUC3PdnUv9ErffQMOv16QQx9E5
HtV3l9mR8KTPdItqo0h2RyYmJo7Hon/asuR+pAsE7YN2OzZ0pOJoRB1PYBNyhZis
r/WGjDvvsodQ47KuXZj5SLOtFjv0CTy0NM+gdvYBA/5eGbgTAy4FI8gou5+ER8Se
+QETp7gqBdgdhaT0YPYdPPqqXudlZtzYXgHeo8IS29mhxJsDMjVuvWhNmIxP9PMP
ZLHm8+n1SHayDx2LBweT++LW8Th70qGxNg/1VTtC5vxNAD1fzdMP3R/AErPY3xzA
RlLx7vDucn0ZgaUBZTHUGszYPCL/CiVphY0BC6oef+2iv4IW7LZJ60UtcU76/GnI
to7UOoBoQ5MrQr0ewEcCsMd4dlNrli/iIaYRW+vSs0FRxXMd8Vm4ZG6CaqPaKrE9
B6SCc032gkGpRTxrtwkfAKUyM3n8s1j2MLqcTr1ov+4oxTGbLtOvwJCpWMC/jCcm
EQ9fPsJzJVP43tFKFcCukB9vd29cAZaJCDAXc+hInjqzjVSi3KbL6FysorTdJprS
EDjUmj13D+HO68J9AFr9qXk34zjnjm4IrnjJ8l3A0aImIHBhqRRePRUwlmlKxVJM
PwT+xxvg3IJfnVfinb+2nV8oMYA4kUfUAPlSGEFOJL2holwcMkpLCEFUuLYhvzWJ
a98+hjeZTIPnaoKyX6bi2xntHg9B6hUv/26Ce8TUIQvnOJiwgw5laZpl194Q7T9t
RHXoh2hCK5iDrizohhjd2h0HqaZ45811H29a2nb0q/pplZL61iKJX1CijkQO7YAf
etSMDQSgU23MKi6+kzmN7b1V1PvO1/02VHSvqf0RVxUtXRBlFc8zjg309VvtRZBH
anpihUNlaNDU3BNuRgCJeegZwrZDVVI2AHZ4x0IirldqvXKNusMEaZFYfKZzgYRr
DuP/m59CyKMvgFWfeLow2OdmmbYiGJPpSUJVlr7BMdxreozpgnUMlQf0a/wJ8l2F
L88vIPKZJFTRctqrvKipAR8XnClaZkMJOGF+/TmfE7Y/EkoEbirrVxnq4fv1Rh6d
1czbfDBpeSp4fFB0Phyw7HuJM1yeWl/bGDoRWf0/BHIQTy/QPZYSPuZchdh1S+o0
d4hQPukuX58/u7PP87ZswzIeCktIe0SCyXtQ6mtMNZrwHl9QmKV0WV7JhJ7hVbdo
eleCnJw13QoUso6D5aspWInxj04x0ShS71kN1dwM0YLMzq0lkCARb3u0wdbjmMWd
EiHJkiTzct2d1XPiuDJxTzymh6F57c8NkeEQFTbZqzm+TwzW7a/tuf23I/m6bYSb
nvSO0yyJPMyxf1Mg7IA8/bG/ptKIZlYg7nunne/vsDr1/D2wIeQHjdz39kqIbRT4
7xSTS5r6vN+R8sVBWRF7/ZdbG6f6cEVUKsVKBaYgsL43HRH3bAnSruOMPveNiJgL
B7TGEnQl9tlhqEIdEegbBGegsiLtzSul63xxXkDlLj3wHhcySr8KuZLHvITps4mc
tHKbH0/MbbM2Nw2/3M3OqM33nvIvC2tq7JZpMemD/Z54+3BMIJCc8zc8qR1XbmVF
3ZylhXJ2AzbZU8e75mM1Vew1tq3dRmZnAFVXStHhV9L1ahPP+hO1ZlUi36A3oQdK
BoKs0ncr626uc9PtQcduzaVJLlIXInwQG75vo3O00NdyZNA0p465JoYRjkFVnx+A
XU0/OSJ/3ghnW72CjWe8lmK2ukjDJxWTUemmMLV9I1ZUqN++TeM75eLVqSLGHsi5
X1hSP4gXWabhD2+P93m6S0QEhl/gxGCYFaGgM8uVa8AUc1ESkkXMzfKjzYGbU8et
5GKHJfH69jiR2bsYcUNKbZaWwa2SORWzxGpdeGQG5fGbphj0V+rlMxBCifOaiotz
c53TQYgV8JxGGqSEaUSQ4HPqsxDyKO39DRDEEiHDADXnq53OgUIPd8HwA9gP/tSK
JFLsIqcIV/HvMhJyaizPpwZZn2jMxp5MiPqfL94Ri5Zy7/CZYgkOZt4lmUiQZ+c0
I6HcKiYHKRmQJGcesA7vHS2VZHQPN9sCTK9giCD4FKsBWFYspq0hdhxZ2HQm/kwl
cBzYu0P+PW1h+hRWaXZAfFeZy1Z+vjAoSHCpuXl6quJMXnaGCJkC4tyY3mb6gb4k
CECE49XEF1hnpOc53lf9exzEpi+SNq0c5Ctc/DXUq1DbAnnk/jkw4CJiV2fr1HID
WNg2a9SIu4xdny7aet9AWSf8QOS2aw8uit3qShN63UDbOoMwT5+YhiYdernSvK1f
tB9ggEgC7B4GoPP5ig37WuPcg7jKIqlr/5ZBaOt/BZ+RQkXfUL/xvALoOSRuKDbE
TYYtTXzHcoqH/JHyRXSxw4AwT8Yhun0BXk8vKzmv8HUlM8norYZ9sGFHa6qrwb3w
/nNv0eUWwGLyXST6WmFDmEwIhriKCIkh0LNs5djy1q/LHd9mQFH5HKwXq2L8xAU/
rAAuOhliCuwPgbcdSgP6eWK4h6fBRB5YTE5Z0KqopJIiBlqtfzolrXiToCwxY1Xz
0eAkIcErwNFmCzLF8/35htBmRqVIQv25dsQbkuZ0SAvvba6IZOkvJrguVDLcv6QF
QijsHoy2sS3KuVRU/e83e1eupjrR7m2XXzoN5gPv7pKZy/3zT5ezgBzgXbkdYypf
z0cEqkjGf68/9QItDlx1xVOqiJIVRgaDt0Yc8JCCskotCxCz+0JJd3OZ1Fc6+3Yu
7dYX7ylVdz4FnSc6tadGFN8sG9nf9eOU4PRR/AlSkXtsQoXEe413MHX3b/TLOuJt
7TZD01ISuTtCiiL/bPDz3CSM83h0Lw0Btb8S+p2MCb4V452IddygwwShgQvk1rcT
egzmf8I/rhHJ/4VY4F97LGEdnZoTyfRvlEbsFD1zGmrwCmREgXK1/KubSeYEg8ly
oHLGTmIcwFqfFkljrIh07v952u0c5rTF3ag00FTop4RTpcTiiL/V++vRk/ZAoT7D
/PUwjv+ZmcS59ctjszzKhK1eW+/bYVHXdDlXiyZxnfE95FOLdH570M8GqLd0HaB2
Rw1GHaRRMYaJvUsO/6+7F8AjpcVvnCQkhhjdvE7DegWrQMMeb/G5KGglki5PLAVc
0BlFasHRtFA4Uchq4QLoRof7JXO5emoZ0tVH8Wi0WhDtKMsSFRNVe7L0clkUWQ0+
gbqRuNMGwArk2z/tNvO++CGvb4ldb668bagHp9/WqJDaS/DKGlYwDOjQa/GIlRiX
nE2GGCulxqx7R/rvsgjGZToXGYszuiVeBpjflbAsdbECJYioYkb6VjlwPE66fuAe
zGmy3vf7xKuwTbEO7ZkIwOpti1eQWiKdOeH8HUjfoIHQsLh7FMEu99k086u9Ibe/
M8UZiFc7N9FEpnuiIAqJyNMKaQjFa09nyuqttk48K1KrEZzyuOO9ETtajNeIsBRa
WlJXcFdeGePQ4Yp5k+P6Th/k/c5mZyND07SZYxv2kYYiyNqG+G8p6L60ecDoQWnn
x3TN5LrmmSQpnurUYv3mr9pHv8lo5Q4X/X4YM9psS87orIj3I7GwN/5kJjQGF3t+
4WRNRzP6Sp5RlZMtZy5VcpmRYJk8h5z1z/Z0ogWlSMLdpvmUkvaQKEn8dS+PN0K4
vKd8o4HT4AhL7+RQv+Vpx7IyyjRoQR1lvqeGNAB5OsBlYn7eVLfdpGIWldv0+Sb9
q9N9BgcFIDts1DAH3Jqd167bAaSXc7Ay+Z3So2n/CBJuIMG7RPPz5JXQm7M0f1jQ
Fg1/W1L9yQU1TLGQ77noyfyTgxvRtY4jUUpXnw2q3RVwL0VZCXs3iNBz+5gCvfVM
BcVxVf9v+/hc9q0p3rLA6Mg8a5UERpnSQm3oh5+0k9cawV/dphnpfO3h92cPkFU2
B2NrwzEgDBvZDRQWAVTZk3yJnC6nKIm1AAnRiCDhxKoZcECZOndvyZ+WFxwjf+lS
vmHcTuI+cTHbA/MdrmpnAT21TiL+OEoaTE7mvWySGX9+8q2w4pn01lk/5kM3YuQv
9Lzd0Ae9JDKUwfU/CJr7YhwoXYf/ECXti21WxwQ8URZ57TCG6SKwcpAxNWRzXzFn
hcSVupg9pRl2k3AoflJniVeGA73ql3BH0Dh0bXyk4JDtablPTcIN6Dfbd9TOLbWB
chKU0Hp0lJt1UwWPTGeVCl7aGoxYQx5niY4pdaJdGUAZtliVPeLtN8xUPfzlHA/v
NPsqNJDgdfbaS86WOWdiYGe9SB4MJ8JrOpE2wLqPKDwpivAGQLipi2hLnCKh7omR
Ywz8w27hRn7DveS7IS5oxmLkKdB3XYxoRk8INusPD7+0qwZohjL2xLnOoJH+It8x
2vxIkkBvK6W17G96/3DtjKnNwN2TZzcHYWcGagtLtI27wfID0DO/SDf7wt12LcF2
yIn2fPJc9M3JdUOG8JepdxqfJQ2veBkMNd6rEO4lQz9JmAyu6yiqHZu514ToPL3r
8us9leafBHW7UNcADvms64Cs37OYrA1O3y+OZnUp5YKFIyTk2rzeYfAxhE1tRh1g
BNTH2MOGenHhOljhHxlpVH2KX80ZTIrtnEWV+E9L3C4ZPSKj8n9GWITm/yQx0xGy
4e+thbWrgCb/kpQJiMe7fKbVQwqKejCexjg7MBOX4KsQ1PYwFO+6zkdUdQ0qa+Np
BUdnFFk5E680rttOvSmaaQOeeu8zT+ybJ8H/khBCwb/TKi8Mkijhax5WqoLaCCFt
IDTSc067QKkOeqmzH8fAcpBb0Gk7HfXohGUVcjThBNz9Yigr0MAMgITaO5yjAHPg
U9ZqqtlY2fSD2Kapl5PVcrwud53aV6mpUDdsHsg64zC2zAF0l/6rWatX/DIrCCuw
9X9j7y+3YQTXMIHuCe+Ilz+Cz9IXODfXGyokwjqT9lat/6bklwaeKP7mBOKbcuBA
OVgXuTIG30rQY8/RaOxVllKSZg5WDYVPUllhFrUjb87W3IDC9hsWyyAidLt5b7R7
QPIp/APZkNdqKUr9SDgJpD0hGtgSjyvfkvEIUryttQlv5RmhnCKrKUsVnElXIX5W
1p8q7unkMZ7ew+99ptOvXr4mS4Kyf+jALCcERe0P96aZ23QVKGrJTw5F4/juEOUH
BM8GyTnwgUM157EYnGwidwe4MkUa5tfNIhbTM/6RNZJfPPZyHe/9g5ekXwAKH5mY
XEwYaR2cBxeDhAZ0fVVjpbltgeYydTZu46A+ceTDhdtvP/qRYGGMujiX7O553gv3
ZOMfNdz73d3UCGTQdsi9/XE51y8PMOTj25ouWPFVqseoi7jAWQbxlfr6nMA4X+pd
c8X+YqFyKGurVFlJHVIIaGT9770Dp3k+yKmwN5VOvMja/51/ccjLBlSgFLJue0jf
Ovnls0BCfIzgt5H4t3aNjKQazEiVddRhhThMFVmS3u6sU4X4ZwWNs4r8JSYidBph
yGt7pEFH5dP1m4ZulCsvHWaMUNKs9iH5uZRPRh6sYII+GIClgb6+r6VIDtmRkzoK
D1D7l7SzDs6pob2oARDnROTrARZET/0xQQHUnNiIipViX1joLIo3Ko3mpAVPpgrx
xOW1SGzHhlQPuOq/bkChkGrkSL/dAc8IcEDd7GwbNPUGpAov09nOg8jvP5b8ie8Y
kH24X5LYALp/2eje3eAe+ulNTZ51qi+NRrqyRf6Dgvh7R89bLAoSELSQme+VKyKf
DCkNLyDJ8U1LVUNkccBIAzWp0Y6csOMXbfybDglnDB0TywTSjhu6Zb1izJah5w4X
RqPquMH8PCS7+6Hy/J3hyxTM4+4n/H/GAZ/vultLw7StnUreiElzDOKW5bysrJnM
PMrcP5oJ3ZXM1I6/80RGsp+jNb2K7n+4RpgwczoVHrEfNIrNDllGqqU/qGJesAk1
MaECVusWuGTKUx1UCy4C18oNJbgT2dR9+E3ZYrbVbAUPHX9TRdYr25qmT6L85QCC
PJ8xw+aUmnlXyeqGHxUyDpW9rEpNVCk4RxLhZQVOz2FpM4rSK4WKMlsqefChC1h9
zZj80J4snUcInRdz1dUCMFgjCCA7bfP3nnOxYt33SkiNn9SxZDRKtCno7QGyyWix
nQ1Kcz+luBAoA13WMjdBB7Yji06MzcaOqHUSgwkqoLO1B6CGkw0aCQShBPUC3+6t
GrE81YCGMDXYt2EhZu9LX+CioUCUeI16qL+qPh2jlFs5e1TASq61mw5Q1Tas3G1J
GeGOxPrX4yFoXgMDkzKDr+un2fdMiq/H+VZkpbLqA08gsgAUOH2HtDnkCHDZnC8H
8XuDIwHy+OaQ6WmG4dF2T73KCuXByhODJ+Os7O/lHZlXWWD8fIUNrsiXiJyaZBHc
QFmcVkz3+djf58gAURTYXm7bU8URlEwXdiS3RF7DpUo20ZbFsbjjjmeEbccZLcf2
/1ewf0r2wMzxuuEz72ipI0PsUqQF/6rSVK5lCTE3OToKE2K4/49HSe6wYEz5KMEH
NQoTHWTOkP1PwJZhDhvbvcdq8Rd1fjyxALEa/qNaM7vZnGNQD3FKt0YJPztnGXBe
WnAZgeMibJaLHSorVZj+UqwWW6KD2om1WPkDZ4oRdvUxklP3MW1BhBUPjby5DpLM
Zh+yt+xJH8+TpoI5peixdJhnjNXu/N5Ybxvp0eX7mQwXmZHbNroiXUvDGh7wLbeR
E+JHc4Avwp72efxQsw4OebIuG+WaDdrY+Jw+pHcnJ7fEh5LBFhGY57NCFPpRymJF
GjGPXxTegIH/2Riel+K7PB6cP6wPIIQVLZvHC1edGf+tdhxDygmC8Hax47JcpMzr
AWL1SYC/KzH48VR4xGPtdfiaz+dzfqWUU2IrL/9GMpHT6xJCek/CrIOYnwzH8qG4
2e+guIuhW5LtqZ+bQTY4HgCio2yVIvbwWj6AYPtI4Y70V1IqcW0ZGppzhLjK9OhQ
UQv+pqrhTN5IS4cBekTRILi3DcA1raymiLFCYmpbhnUoa7Bx9/KiGP3IPzgCgMiv
WxG/iOrT5J6ZdYiPSu0AXnhT4v9/nKN+nvOY2Lu7ZL+UJosfodEKSMVs9pG45rIt
BMJKMP8Kz3ES/X+jy3hxHTATgFUJYYGtRJlEgtmjDbhLUhNEYZUSZbohPUYqXD/7
012XurYURcPGU7BB1FPm6icnhd6mo/+89/UXIlNwI5BCSnUCWHBJYFL2/L5xPtNy
keS/n2wgeF/mwXNzdo10Q/yk4wrKLcwiSC1c44TrekZMSUBdWZqSoWTHhBahaG5O
E7FNZ7H2IpHAuirb1zFsAFAwNKo5U1LMk7KblXH52Cz8QSD83+VGFFoHg0Mw3Xq+
1jsD0fcYApyyDL+09Qg89UtY/9600/HCizCucjNEYdWumESxdnOPS8HtsUOp064C
ltJUU6kId2pXsFgdqkLOHlcFEiRZPlMCyeYvSK37U8xCkNqlZ72+SCxnC6lsW50/
A/oz+cO+VGoiI0Sh5m8XSMXx9nAtdTuuckQHieptLjPDaJCapnM8+R7AklalNz1p
rx0HXZMTdPPYt3/oWuJ1KDG82pTC16jd1FTWaAT8BwewLu4jQUpi64c1MiaEnWn+
0etmRaNEzPTp3dBFQBALH1OFdWI4UTgWFYE36kbnduD+e15v5mPcxYdEJfbZ5wPc
GuNvJyjhJXuCUVu45A8k2VkBcmBiplqbOwYkeJcJzyw6HGtLCLrOXqEPnhm9hHGa
xzfYP4DczNT3p5yeTQML2xGhiSkVBwGVS66cTdoOo6SogAa3MKVvvGDfEzU0dZ3C
kAjbEzwZetOJJh/ul/rRIi9FRKOWmmHkm4Jet5DkGybu70mXnUla1PJe0ADLkT+u
3tljwAtZapiz2hL/H1ppusVL+80Hial5cbCsZ9mvNS011iX0ZtieMdTIKF4KEQWI
7/VPGfjEB2e5m1/g4IRUVt1pckz8tzAY5hOdtSIEFMn19LmS1jin+jFIb6CI+BLu
NNhdBmuutiU9F0YFWrQKujTu1HTHDoMnIfvO1BodRw+5we9b1fahGYKA7AfhgXP6
ObJQhM2C4Aa/1LodgBfekz7pLzTsK+ma7Bi3op+86YR1SX/+7TD6Y7j0JD5smnfT
Wnmai3gqB8voNjmeCDeCmQ5au12VQ/ysTSHypYZAy1OJ78x1kPFOf5PXgLfUQPSq
qrH33wcJwuupXbxeNV6Za9GiUoYnE+7/qFUsYjDI0sRyhl9MNsemosZwol873SfN
Tsk8M3c6PmKN05aBR19rV6j5M4EheFReUadyQ/LZ8v2Alwf+SLpVnNFzE/Agoo+f
dxAqI4//tj+jcl6sBU8VyNissKJAoA2pPBz9k/+zsE440MyurYUJDkiolBn5IsOI
mnxkdg06+hcbIHrK2Ns20nIAJ+YN7gHhYqC2/y0ypUWwv7jFCKYsAU/iwkDBUMBM
f4k6VCn1Hm/cZBye1MexRd5m4kxOdJiavrzyemjTd079DDJEPPaR7NhwX8gN4aKO
qWRgVPcT2QoD+K5O7WkCiGilZbkHjO6M7hqLZZWFgqo/xDZ8l48q482W6naWrDaz
nNZ0UGk6xvYOOUvtjsDTYIZwX34Qe0nqfqpqeiHFxxmXNy9yw4cHfo4mlGVK6Al/
v3EBBNfGczv0q1UZPaNuyILx648MGJkzRxYsQby7DPGnOlB64vwQH/ayCQ5xVngk
6NEBmwdq2Wz6HuCqvvkeKMXUQJWIilasNcDMe4ZIGz9vBuALTFWV8AOzFN2mzCfg
cjCUHk2xAHuItLqrSrUtu5tnHzyS6esoudhW8s8gFy6Hz369um6i4FU7QlsJDUtq
/jkDnp8qEG4sxzUnft4tJAdLIqlvf9Vh6iOyP6xxW3FKraoO2LeAQJ6T865abeS5
THmZIJ83vE4zQU5tLZwHOvUlOxOkWHbpnVnm59z8AtMjTRPlhi8+bEWo40So9DT4
pt+pKpKP97RY1ISknK2yhnaZTrbP7higetS/dR71+sI7CfWFUN0onBHrD6cwEU3r
wXa9S9vVNvSwvNifOLzyHJQYzXFm3oPqAPkTVJCuHMjYymopxHY52KAZS9J1tzt7
O28fA4BE1AsJxti5ib9ccoCPpGG7qtVtEXZeTQR8nQL5YqS+bYcZieP747pCndnt
y40EnVcUCVU7WgqyBis5za2eCXVJTPKy8OYbAU+ChXjTHZ2wbCUc7I9cY1+ysQVv
T+fIY6z7ol92la4hugMJgVWgAtXFEocceZHG2T/VOiTCM6pGzKzfOUG4GYczkdBO
ahq7VtPiYvQBr9Me5EBoD3uIkSmFaDiH8aLmq3Xa1CrjKrXods8e3pVp32mqds24
Qcf0CwpdyVW2+Dx5yyvzF9STdACCAyub2vbhNjDafOjzAQRQ5LiVxwXPq9Q2eziW
HGWrcJDnJKB/syi7ItTMWCF4UUg3I0AA4R5eAj4Q/+w94dg1kCArKg8RItthLglT
kMWfI3f6Sx/d/ba+1XAJJq54ooHhNev2bRVQOJ4keutpSXAk2bJA0Z/5BgDWPlg7
9cDpB2dXv+TmXjbKXvlOVJyKJ1kW65NahhAdVq79yA3izetJBAYb3Zrswfik+RU3
0VLA44bIimKtCaz24HXPkaQlXTuWr1+Uztn+jjyQ5FsJU7uGN/cu6ZCIkN4BSCQ4
cXAOwOyLXICGKHPtXUDAyTsqF9jq18aTQZR62RlhInWYaJaSShvekMspzvPj+Uni
zuaX+qnTZtY0y60pYARqk6hZdjveWuuSlyhc8Lq3xl/C4LyLe2WXjtjo2qfjOtj0
WqRBvShqgr847kYl3pL5yuq5Ad8AkHXoz3+Ss6Z89Nb+jD5N7uFENhlBhKI4vE8H
OMFywXYMQzaxgbd8YYkP4hTREHJN5odYc7x5bc0E4dcONcrFj9Ya7+pNf91fDGuZ
e5WJOf0GYVwcPTRI8hbYq2+N+/FbPCWXTGtGK7zaU83jEARjdE41wIAmTeDkSclc
iyVpCvj8grzOMjh/A6g3Eo5MYGbE2OR6i+9nvIs7zEEiT1joT1NooLCOqM/dK1dG
XKPzzaBPhiANEfG4fTnUsuQqIA08t4yHETmzvBtvT1Chvof0i+KtTC3eiVL3oepG
k2U5ReFqFjkzTDXlEqedVaTHVCZFS97yKix5NHfLrkOIiU6YRDvNO+ZiGjszos4N
o5sd202YW0ryMWcj+IbK/+BF0h6f6b6M/NH5UchrNZTDJBnhGIotRj2kQOwniBcs
EBiY0VMHhmT3/0hJOu0TWl6kGc5Wl5oGmleqmdU2eZKZBSJneD8/ZVCH9V+HGtmh
DlYDeHcjBMnMzm5eybjLkB56FK1A8AQ5QvF4PnNZIyYNbJG/g6pPeyetMDLrb8Xq
MVhJh2D1wPqGV6Z7Ma4yHGf0GVuBWGT91cHm2GSq0uqOenfCf2CprGjWwfp46l7b
k6RU0VDR+vkPvN8t+l7wo5iJfqoeaCdks35toVjGIgil1FIwL+u/ennW/dchcASY
+DT7SVVA7X6BFup3SYgLRq+2YDiVje4Ry/CMr/PGB6Q+6R79Iyj7icUy6lAxNyg5
fuq2clGSvz3sItoAkseAdw4HZBV8F4/nGCmFR/DsHyR+305RRddy2tIuFMW0xc3f
HSCYUooqwc7hPLHTe7R2W8iAP8BWDG+OQ4LlM1kCBLjoKSdPciZcxBd+iFUDQnmv
6AFyCgm9lQr1RCFxUiW015TNsiuLpl9nQ3YSFiVB3GwxWGs7Wl8Fhfqxiwcp3Aw3
4Tqjuj2v42p0hk7sXW50Rqv5wpYfsQjum702pSHKQyTHM3BKrK2HGNZFd3Ze0l10
pnV7jD33RJLtySxhbbSV4iHRPe7SPwAavlj3MnWsLrGFU5+2Dpg3BY8jB7aOCLlc
pSBfsKEye6IWL5vvATtUs66dTfl7bB8WVu+wcBATexOKc9gwXVcEAPB+sfKt+Ao0
2lAjbPKdDJTgQxhjTRrH0l4vM0EkLlYkFeeLxYO/VW69W9xP5lRWwlR0d8bbZwC8
LY8k9I41+sEUIg6ZfO6wPBxwQsl95ArnumXByXuMClHmXaY8kh1Kt9e9DVoJNT54
dxH4zrQ/IqEpQRmJTH47ZqIRp7JfSFm/50HRkVtkjKPeznC8JA3NLTe9J+xLOHgr
EevGwdV5cHISvAxRZsRDwx8DGck2zJAHz+6G++OLydrH4ePRWoHU1ZpmUw1on1zt
bcWpmlUoKwTnTFlnVjtxGXy6UOvoReS8tGfqiF6CFlk/Guo+DRvcMsCT7guRb9sQ
WkI1ZNl7ioBMndkWhYgHUDsWKF+mCnBKD10TJXuKcbULxKpfZuzlGtjRQaADb+r1
5IHt3V9vNWM0+qORXDbggaafG4X8mIGFTxtXdrD4eDvXrlDHW9QByr5g6DMFr9tr
fLJOOXpHknrabyyUefEyJtfgQV6sBkRZjdis+i2/J8xuL/aJR+oZHFf03JiymnUi
4luky7z47hvq87pwMzIdUeM6rIQTfte03LMBNK/OBD2bx5kViRxXxanJJXUcGN1l
80cGBUGQDpv7L4URwAwGEAV7317ScU7CWNMssHKVeX2qcqsaVFg7JNIAhCMY/e40
hMGMPvwBk5+3vhS5nfswei6hb5VoHe9/LzHCtO2lnpOb+p/zk1fLWBnLX82YiiXX
wTCm5tkO7i+V6OIyQZQtkzE/kdSN6bX9FzdtlSQvJdJKmYKVT9YAYBeHwBkxyl7c
2nhIz7l/b6gZS2nmGrJcz/X+ATPPE1ZHVCsbjbYXOTeV5gTzA0GLccf5CmkWvzKv
0I6NCl8P9sMIiNoTsBauRa5szfsUJJ5IC4Z0s60ZauLg8foxuLz5fVoJ2RoVVC2A
qxlz186m01E1p0hvxACewBe/QvNHBq95B21mXWKHFw/a/THuO2ODTko0TG1KavqK
o+5uCDNngXL0yEwz4xPD3nQPUGnj6OlEyVCSw+5KJYLSYW5wb257MctGY4Nahci6
NXaNLdx21RVH38MmcGD3C8su9U2dekYxtPWrUzXK7GpHy+LxqSAsCZE0flF0ViGn
mQnWJyaAwrVAwacsO32M1BwhxC0siQPjsjjJGaxiWACkC6z+4O1Zt0RY8J9wQb/F
ycjTzdghMBSMWL10MBEeukOavjv7QZrxel5tKKO+/242hIzw3S9/fJIpAG5rCMws
7Gr0eLQLm/Is36W3BBwcXgklWQUmXHNl2y/mzZe7vXnQONao+3h93zC+gIy3poZv
wwwB+9YfUw9U4kNVCe6+XO0zrd3ODK/x8abRS6fdRWY6MYhLUHzL3aOgXdn67nLb
I4Jsm35hKB2jLDZ++u/ZuxhMUTCt1wxdSG/7SmLurmXNE3mT02JRXEYxQDpLYIWr
qxxKV66l5yFMUEmZ640cA21ChglgF1YIVxGW9PgAnnZY4QXoWGbJdirN7alrs6XX
rzCz9H8MjEQFbb+dsAq00Et5/+Lq123r4onQsrz1F+9isM+LaMQaFXsVBUuY9Pii
T7UjqJeXQR+SS0sfaz6CGjTQrJWh+FvUch9GRc9ybaG9UwHM+iDVRHjfBRzzwqhX
wphfJvT1re0hxD9ZnT/FghDldVcW//filOfrUj2IeSdMgUzz2vKTY/KVqaQNDi3X
9u8o3GBRCk2nUHyofFcm8AuJcqGVxve4cE6QoXe5VMfiF1vXBX1k+lcYe1K8wz10
uZSKAiYRXqgauK1/xo+mhewYVD4YUC1itoFwKZZfP9pjlfwNW7yo8/7hN0OCdq1h
Gvm7SFGHeW+HM8tc8cBOL6Iny3AnKyxNkl3anLpTxUZiglgZONGz7YsfceigSD4L
bcQdnBwlV8pOItzXHK+CfVrrz26LFizvV1zs6Z5tJO9aeMdyXwJ8gYCfHd/YQ4rQ
DpDnJxULmLkvfqiW78WclcLjbAX/1SNYyuFAcrvq7ANGyQ5RZtAgRBdC952e36K6
P2vdkxH0r/KSxNuoC9WawlkUy10xCW+RgxMZgbGoSajHw8Z2lGc24cSsORhlSTCP
JYPBl+BvhfPeFaAIQ4smYvV/Tlks9nN/umsePOukMLaJu8HEqhT7HwiDD0okzflj
f1Z6u0bHKUVCdeOTIH69NaozXVGHrz9lFTsXOXgsGtf0j35S8ITZc3joh+Rp9lwK
p2myOe8HNURshH/CNcyXEko0XS9v05FDgpH0W8+crq6bTyaH5vQpxd6Tv2OvGBnm
yk3PBDU3FFBsOoZmbYCRBRQYdwdgnKWVvCkjPzkyaUWak3yWSIt9QdFiT6srktS4
29r9Xk0oJoaFHCZw0jNIN5nz39lJhmwotYRSn1WKEEnfGWP/mDCr9uZdhp/OY7TW
gkYWLtFWALIkB6DO/iILiXpgpO69/JRuGObOIWwAEMZNzFNFCcSXU/u2KLdKqvt8
8oPLifK5W/jN8LGwKI7fv4+OFvic25IQQjdf12e1lAxzR1VxrQB0Nvm4kn6bPAWL
ZN+LSK+t9AYbalGlCRfPo4AaX4OkleXuVCFPuptdq+24egme2sYpdEHNAOeE9JBb
PSyNYonRkXoIFjYyDkPy4cK5okAo/j4ley+0NTmAwWi6MkH7gvnQmrGIxxhxe6nD
/1UJwOOGsBSPA8EsPWslXJgiHbif71ndxiBnmP1glCbrjMvjh84OsXt0La0BYp7N
ho8z8gAa0xSvHu3lpNAMCPYWS68IRVxrXZi78B8+IYlkM6bHLAZSZHxpGXCuYY+d
Tafk0CrQ/Csgl6ILa12T6zdBTK77Y+R6LIWA14K6+ZtFad88u6pplcav39LxKeyA
+08Hw6mI4D/o7Ha+MIW3PuHjzLirlaR1pCPRbCT/62UTlhr/8/D4g2q9VRjlc+Tv
hiNye8xZ8fXAarePGPi/pMYX9jKPH/uLJbTdlSBPOGgBQkeW7HrOx1Is2tF6f/fH
Ye08esa60AtFcbbdAPTXvkKJSAVf3qKE7vFetjvitmO09Wid57AngH6pNdfVaS0l
oWuqxOb5JluvRrRxXXlulI8trrLavhj7bOwRYqMb+4f0g54jbWDC9RxPJecaKKa4
fnjsul2dMeNcH4TnCbIQrBnlQNyTQaylmtLNaDcT+IzzWEtfRyiSKi+jRgZDOUUs
fO2cqwKpdtSwWilXep8vUqEVUbQcTI0U1h395qJtiXhj897TRJTpHIL8Ch/TmvGv
re6hYWUIVdSyTooR30RD7dJvx8+/ZMdpBD4InBc+G1/6lcot9Pe+fOPeJ+r29BQP
A8pp12S6+GVRrS4JT+fdf+DBlUJfLg87TSaBqQ/msi4pZjoVg6oAQautSOWvhSuB
dWyp9KyuVS2xtmO51EgKkpC/nPnU6+79YEkFwRojgHLzeMgc0cT0SEEAr0tX7tk4
kCv35GeYriasgc+F3RBLQM9GJFzdDk2yPPM+OmdWcdR6yqbTQrpEUZQxB+nTruPC
eeDPy9S0TydVwLhjgiG/mks+PnA1mYJs2bYcKsprmTAxzsjrQVFpLRVOUtc8SjOn
oyMe4uaPqqvw17Zt63stXcDEx1ThT9G/lElXglxUeJ7Iad5tYem3v6qvabnE2elQ
A6Nn45SdiFZHFXcGP8yBoR0b1SkXUsDNLnbvJ0NsoY5UVV+totFRRZzHz5+SM43o
cKvzf7GzRFtMENxiPTjspFVznQwlhXZo+Jy8+89zztpetwMq2QRrohNW5+ncDL0j
9CvMHpkCEnU3EFDwHsVoh/23j+tw07Wp52G/4jbplRMh5iyKWUTODbdR8F0aMJCh
kP4XWghGcgZNO+aVxO8nrkYykOIc5YnI8yCy1DxJ8a/WvlkWUgDlPUlnxJziJEEy
+kW4W4r+MZ9LHgQBF2Jk6fLLlfi4GIkwwb1Yubo2YiSE+ptEOcWbMEcrXe32Lckz
BpRYLPYw9ne4TqeheilGx/UMlAlN5imiu7S7G55AOiKxItJagefl5mb00nPPZ62g
bvKbTgU022AL6TV7FqNGN5oiSAF+FcvTiuuC8N3qG8+mZ/a30h0B3EkQNuJnLzFH
fDbnsccQ/3pMrUR/1SnadcuSATw1rCOrmzOQeOmxpgcQSs1tCVUVZuF3hl/gK938
w/B4zN6wVK96qjcKLHUiyjg1CQb5F5kLgV91LuE3TYUHbl2+zgj+nHhcJ6WDqjEW
qA40kegevq6xNCicUNmOyFq4oVjghEzPN9af9Zm3JgPL+WFSpHAdSTKRJ0Ye+voT
+z4fK/IfHUn7+TmnK3DpdNzlFV7jeBLCgpgQvInNT1ZXdggAPhK+4UUITN4ucW46
fDJFeYyCVBrIOBuoBfJgdeZCRl58r8ToeF3S3U/hyOMieHnh/FusaS6Bh9CcdIfC
eC8F+hXuoJjERmtOoUJVEXR3v0JkF5/VFNsYLSerTyC1u7JQRowWAE7XAJxI6Mm/
DCtLSG/kOfUcpd8M5zX6qOJybmSJKE6K6qrN2hmR+7nD9q8hklYuafaXRc/Ogw02
zXtrp8HHEofKeDcB2y0g6SUgdK4SJs3MJway1euxyLCIpV5DXbH9eB3b4xsEguzG
QeDd4ReaPSMRSzJ9YFRWh/HwHSnxXxA5PbecUAvxaE0mpkMU6r42sy32Ick9qlM/
lnoj/pdWZNb9Vwxeg/rZaubIQWUtXNsMu20F5x13rVMMz9Bj9XmlEKtmNQOyzYED
f01ixrKN2M2Z4PnAAqFWjQz44+HknN9di5EwXgDvSObEtnhujEH9jkzkBOV2DoGR
Im/v8VPg31C+YsRpGCBjn1nUkZ+6k73TyOYcqGBYsHdAi2yvQj3QtvXk9pYPRGpn
nx5pxeWFyX5M7oV4aWK+u293i+3es0pQsUFLPeF6Fe0Ov8zM+tpb3fvuyBsZaw/P
4lbTh09/2izsrPj5wCAcdMh87o+WoYEuei0Rlat7SFopKI0dk0v6dQKqT37HuV66
MkUtl5/WM5N49E6XNCJDEmIR6h+M6WnM2w4Qw6cLnXo9wz53FfU61u9IoBD3+KYM
pq+NULnOIgPUYi/b7fF3+wRiXCQcI+aE3PLgg0GWddLa+ECRtBiteuxFw7x0EI1M
ytqJMya88zJ/rml7c1VsxoxZt5f0sYnjnbviAF99rxqdifJBwMmb1AsLO/htWngP
c7VBAKY1N0xZaSQqTB/LJ5PDbreJ3SjMm8rhTaJ0HSkyIJoA6YmcFZurMoN1pBrg
PTa+3uikEeMojjz8WUhv2pxqeJrs7BS6lopMg3AHCR/DEzbbaPuFQcPQBu697M8V
7fu2eefIhQkV4gknqR4YSpXbSzwSticmMSa/d+YYjJmfKllSpfkq9Zqte9LbsnZ+
v56uchQe7RrvFXbBbM2SMwV3b3z5ucfH+/63LKuGRqgMWRWfvJWM0RSpBsm3pdVx
224HwtkvidIR7hOhWxn428wo2FXdu2Bn5zEEoGzvjiQpuW6lrX+sbG5kKXDH2/72
Nt2AkNn/W7ZYVhzsZM30I++eEPstfc0D/9YXi6MYOckIxev6Mhp/CpMhIIBg2eJM
nNUhVy6wlmV8GG2z1UiaVCv3xIX69B5KAz7FdObKkQc3p4Qv+/YtYlKtTb//vh9t
0qwnsMF97of1OQR9xb7c4NPIqwqAa1YjNpso/JKa0b4wk6omPSWPrtsP4S6gVY06
CJlkKltCp8PbNwaw5UbBjGOwqupwlE/7OXFzJ1evCnFMlp1Emw/3ukM31KrTYJMS
qx3BYlT6ATZ3teafZGkiv9oNOM1jntGlX9XjYfvUhyvpZ3AyuTct678p4t/Wyo5Q
mW6ysHBOOsjAisUgNTlNTsMHII/9H4ByYDhlFMdAGp23JdinTmvxZRKfoH3fzaQ6
QjP34puiyK5zZ0n1mXfX3A3xJkgYQnZDH0jQPgXvmZLrCagrREN58aHg6LGFfRqW
yk3roEwV429MN3CwCau613b70BlVEg54gMdhDgUSW8HDbDujSxbeME3ebvzJL0zC
K4bSYbk7/r/i9B4rKbOG8kHUKbyWbLuO0zDbXlDPys4/80UK3clr6TCi5P/vACx4
Qt86UQwueuuY1zz8w94S/y9a82PX52lvM8uSMJX8Awl92dfKxOZhmV4wzR7eCHu6
f9lNOhmriQzk513m02DpLag5nMSpB40oHfraDaKAmOIuW0NjEfTyOaWP6e6nSiY1
K3BpW5VoVQP/MON7zrbJ+kkz8eP8aLbqnOtZi0APk9LxNXfv6ZGx8HMQMyWZ8oy9
//iupRvd/TdqEehBGPdOJlJjRC37L7AgFjOeELflssszngPfAhcXoMvxf76TU74Q
P1WdoN2Kc50WwZ42jZ26EPQp53pE9c6y+5QVn7cO4ai/9fCVvE0+BBz3jX2Tizr7
QwzdVKSGQeNZ5CoDnUNdzKgji1vj2dwZ+py7d0reeKL/AohuyUeXhBGWn194CtKt
Mb5pnfHIZMRzazK5BoyYlLQexCqsMKTj7VUTgnMizov9bvJ2JCC+4HeBqxtXoVL9
waVrEI3Sxa914PKVvZ0ppLheELbfVMDYvVKBdiapSXXdkNRDPnkc/Cd/qCbTg/Ho
tt99LlFV0FZOFDccl0DdNa1Jf2vZb1Ec2JRzsnKvmYMGB3A55QOLaTlcwU3rF5Zg
mHqLGoTCPTf7bIgxRBuw99LcbJ5d0jTqX9mAGx39+osbscF4OpYbV25uEaqbFv/v
CU1S4kqdYv0YIJBa6eMQFnDzp7O7k4BvCVsMvbJ6Hcw+I20p1AP2oSCCZzJcorOY
deDsf0uqfw3vKPhA61p/FdJCJSQDNttbtLObrpv4p6TCMDhvTZGolTjxuwAkY2nK
3V4Qhj6Hp017uJ8KKgHru8MDqdfWcyIy4Q1QWfthCTSMQFM5h/Q0j7TkQVqeKafX
TqBRLl/on/z2eB3DFThkMBFAr6YRMhxzXWNmaZ4iQje152GvnOQfLblf+2ZUjTx4
0pgnIf0Vlvve4gMagh9c7zbqhLFNnjuNY2YBh10R4r3ZxDTOmZHhOx+5XuHjRVd9
Qt6Kx/o5OCmlQtwGiNjEJrv+aLFg8ya5/UKDVA4loKPvlgt9/izSKiCxX2Ibx/3p
1QYfS9Nm1cb3pANX4aUPXvWo0OHJ4OK/NQTeU7lK/Hs8AxgiUB++qn4DKfewUzFi
Rj33jB49Uy5ArRV1b1Ci5hHuQ6JcQb8HW3rsUyNBgttLz2av1awZzJxyCs25SBNE
GbNSXur1MQVWC+jbqtdkRI/mfiXqT06hAl4y+agy2P4M3Cwnt7rmuJ9WomU6TJFV
grggznCNOYW8PWZV8gFw1pXJn40GYITy2X24KxM6HxjcgYLb6m//JTx1wsRIWP2D
7x55ve8bvrDCHRhhNzdKS0j0ufkxX5wCXSgBdVlRqSgR4s1rhaUo954LfYMDwOuv
LjQ3KCdUJhufugc33914kD3EsJzTOVugBnEyKpQFl0TLbhoDF+chIjUrlhGsWbZx
rhtwdA5Aqbnt+BeRriiFBQD82PQMJso7lGBHCmA75rJbnUWIHWPAlpCbVZo+mHaq
4nWAUxjp5Xo8qf/LjrTXtyYZM9rKBSYAGDUbHDFca6xwHsXYwu2UBwPNSN/Zx/98
bSJoNHmlqZzlcuH94peokagm00z+buOu4FYJkUZssiUkkS5VC8b+eg7oUAFDzavc
NZJjbCBSe7qd8Ak5VA4ilyIlKE5cOIGKCF/Sk7xfQ+9sDXRocr217gSc1ju7+qDL
Emj/DwUx8Z5KDGrEfZdwH77RzPEEDTg9yC6z6XWYEYcaa9XcfCrXC5mzBIeO70UF
i3+kQ3g2vvRo/990tMKeB1L5ahb3/t4uf6Cj72n9LEkWFpmdemNaOn+k/uhUSEJs
uGX3ZczKbC12OedcqKChobmUTRJ05CIlvW4iffDeIoOmQ2JqihRviaAPvq4g9fAF
cJyA4zKMIQoGtY025FdNI3NxWymWl6ioQcxRwa9Q1GlDkrTXc+JNZQnB36DYgjMG
RZcm11U5pppYNPgTzRZnWEzT9e2s1fnJIPXoMgQxRWMXWLjIr7VHUeJ22ZECFHvl
4LCPwxhfBb9n+4CDFQ05GCtLsLjL0Ra9v+dli8mlJWb5YNBWhWqdGbh32UsOoHCI
xaxUi1rAMEM/hqAbHmmcEyPwGQHMxXxGtDdtzglpsvMcuRX90t2vJYdIviSqjAcC
vAu5Oe/YduVS0GAcDf58ss5GDsfCmPgmgcuilHNqde+1exUR6BIQ4cdYuDQBkVUU
51Cl19ZlhMtKF7IerhBg3i7449FBwMVhVJktMQ/nGxyBGvVemd9n0PIpUf6D8h9z
G45A5X9fCmt5oJjXefBX8EP0NbBFv4FI8wM9Dree1cfB3Jrkdqy/oCt/jE7knfxU
SOtb2oKWzLZDW0xfkl89svA0hkHFie8VL/STw0/HvnNMejxQRdk3HASa5TSrec2t
KV/FZTou7PaFIzvDv94RPXDpk29SYQ+HP4H1HW824l9cul9fNEdhiSX7ZaYRxDpL
fl6VufcVjWiNwRyC9qCHLezu9Q7sEkrIxwDUkgu0lRrWUg1Fl3IXe5/iOkBZCaYh
KXHacAugmdQbjLw0rE1mVxTkaZYk5GyeNkrLK0WGi0q1hUR0wanxA8hmojImV27A
0MgnE4JJ3MpyiYdeOjiujqQ48lbHvhdbwEEeaTNyspn6KKm6+9ODIFVRw89R0FRC
4VBWk3Q+Dzaotvqb49N3/Dp0OShz5PcOOYecReSQFOfLF7jGBNfPb2LmJOZaRQx3
GirZdgVJ0AUVCvxUSS63S8IG8RQ3eT3fyH/pl6wP9MKOQYW2KHOF9vvayBrotAgh
9HMExwE5l9DW55yxhelMpg/jKOAGmnEx4LO4jBpdpMI/sqir8faXq3LmDpjXWyu9
6lOXcJrQbmkAx/dry2Erdej8o2ZKfjWwwhuRiPxGUegDh6IdhW9lMjaVI6rdkG7Q
w9h6LP2s3MbGGttFtB6wmYPWzoO1rJsz+hlYmFk79iOjLm2epsoWF4Z/xNy1qBc1
nEfJkCF0oAERzl6xZVJduosyZoT9yNMq3/SrSRI0xsDK4dPO8gbp7LT7OHTrPHOi
GyFt++uiJHHHI1b2s+D4IjMU1xEBYUlfJP9m+gfRYrQEokAr/JPNirwCJEyij7ur
BQ7D1m1P5rlN/WnNdpRb80FLQk6q0v/AhNXoDV3L91jt+4+y+iFAqurKae5sY020
YdIxCpcrC6Np0a8IBPijVUpwrnOa8i0ovnJ9jsU3wdWoTuLwt8TxYKhegZTlHSf2
Ze0ujgxvLHIsCfcGGLnbEMB0fpoXHqmdq2K0OIK4PXSFcd42+IKpZrFQlVYK6BNe
8n9BbGEjEW5rNphlQ7ng3KPZSarmxMdCVB+jVsGm8tIEmjp3me3K4tze7MKz3sP/
35Krym5S7BdzDfgUSchKHbc6HZo8s3YHAn7BEaqB5iwFJVoGaDgkH8+l7aSeZRnD
c6pwy3e8P1K9d1l0ebLQjVB1tlYfHu4S7EFspPAfDWhmcMFVB4VYVjH6UiKFtcES
5IiFb+ZYH0qWIZ20Ga+ly6LDYdiTGAQyxMVOsMAJVF8re9ZGQ0Kl0fNUXDgGLtj1
1sPr2kMeqkTG6bSvAAa8dVT2ASUnGqpR8GFqSDN0pAKj/Ws6Z14atL8iM+vg1WFK
vegA6n2zDpZ0Pj7xlNrDkB8rT3RCOV9j/DROxgawOQAs4IXJaWkr96XBcJcQYBj+
ZmZcKTCj3fpjcnUH39Z1SJImn1wdpG4eSsOHCAL4V8BY0vb3JfVqrWcVTuE4bbA9
zwNzLjp3oQ17dlicSWlSGprQFDVx1AgnMfdVPA3eCK6D6fmfUShds6664iX9TmLh
D0axg4QsiFNoLbSmCcytnVOZrgiLhq02vDG9/1MgNA3crAXjvjdGKUXr/NGO9Cgi
4+AjobnCnpip7hMC4fKywtP4F/jpN7C30l9v/29frOfLxSVo4/7TVvpz5NmKcmAl
Og+rN93hUS0N1N679qWsF/liC2F1fbK4e1DKzrZVqeb459RSgtO7zNLm5jyWb/kN
VXbuIAw6GJeSgvGUIct0lEG6AE27NXlLTrvsw1J5qEFYSLjuMAiNcxlmrB6ogPMS
9ufbWcr4f+3T2rhq7M0qg2XBuX6SEi9p23iuMR4K+McZFT0noB57iK3FRkHntfyN
9qPgFFcIYHjFQUzX+QxrUUSX8NRG8TMssLmiRF/NaEYTz2CEoNqIZJ9CTdvFw/K2
h4FF4Q7QQOs4eXGxREjzv/f9StLbJJQ5+UjHye3nXopZ2sPMXEwcSLmSr4HkQsjl
YVPSjnOXzReSexkDarbvfiRRzekfLp8VMo+8yP8M3oZXHx0/kwvi1J/F0nU5mCJi
IOCV84JfMs2uvWyUbO4qX49CV3mKR3y15VC4GMFhIevr4LC1TfT1qLNzNVAGNcXC
OdW9smOq3LqkpWbuDwKCjq4GVcHkflEcdoxp28Lzlcdokhey+8scqldFcmgSoflF
nZ0CdB41XgFv7fGya2SF2fVkSDOkNcR6dKpmhqQRuRqxX/dJmZ3GJ0UF07ad8cRf
CXq8gV0ByaprEGdBPPE9fqrC2CrgixCDCEc0wPttWOlDgnkbxUG7kmuLhK8E4eeN
PTtwS8JIXYxwp+KWRjc/5UPjoZhj5b275rrnvtND4PePPw9hZJ9+ZNd8xgtu/IMD
c2gZn30tn+gswK6wo4iI+e/9QgFBVsuwKkd8wZIv7jbWM1G3ZRVT2QrPXn6Umu8/
jx97+q6PdoI5mcRgDEocWQPjjyRJaC/5qxJN/pR1pR7IKtowllMypfS9ShzbaotS
1mF3oXRBArH+auI3dpgwefSrB+qgXesLCULUZNcPWcowRrekEpEqWiPTekbbKY4H
KfBxx1cLJVxlxZYATIiz2WV73HHMfuAvVSEX8hVdzTEMG9mRTg6Im1692z0fh+LB
0s0rC+j320kf2W/OuQKQJfPKbYIhSjWvCis88XOkP1eN/htJ7j0sDdLRyVFK+6B7
2qClAc6tcdrvp3c62gZnJCTROxtaTj1JigxuMJAwM33XhTcH9bJBUyrzihxmbg09
ula2fsKqONvqSE9K6s2pzSYnxSaWIZBLz6I5VRg+nXaEvPBGgQVheInOeTQAqFZ5
cezPA/p74HAegVEOS9l1PYWq0mj029dN5wUwcR4Zl3d9udv4CnJT8KLEBrGJ7Ghd
V9ptp81q4YtUNd97VYv71XdgY9mSqv6UjfPdoARJ82NqBNEMQEZggrIpaCyGUw4l
4Kd78MjzA2Ls2BP3xeEBlmw1ilIyinU+37b+gOTuYLORPA0JEnbaTozVWGDoCXtn
s+B4riyT0XEerZc307cqCYAcM7P/qo6csDjJ2dyIv4X2xGLd8NlYrSR/8rCG8+EV
EBwb10mBmbFxzbpB9Ph0snCGExyxkzMnDomZ8Z7sD6EqWqVcMyELa9r6NceHgpVu
sSOYF3lDKxzxuTBVQtNqo40LkslKjlIEYzJORojmnojdyLj+90J+I+wfczwa81lj
HrkIqI/U4qjKuZ0YYXgOj+rC2WUpmRT4Cj91sMb7YQNIaGijJmUcuovpw+JKRj5k
4HrBRa2DuMgX4v+l7OwcrS/AL1BnBZf8aI0KRNoINI5hEhA2MvLrEPAF/Rt7Tm0K
p8TkK9YlLIx93PPYniwQXIAQX9b0Fhgmedj7pCXHGYrv62VJTDifjpZ3NruUBqN+
XGOHQEpVxQLYcMenhuoDu7LfrERGhJPDZbD+kyLHjeoOmyGJi7zPewtjRxeLOUo6
MkF9LIGB0wvgLZbJvbanslYuKSj1NDvUQQY28bPbv2UfjvfBofiHiyfykpzguz3V
ILM/UwphoxdHsY+qDABgevYnkiXoMJIee76XT6kw3C9JyxF2daDnRjTQ5/+vB7gy
tXXBcUKM9gFmqwovendxUXA7UmFh3TMgUYf9rlqrfu754fvNH0lBzcovRhNU2QAA
KXMp48U9Es9UqYPYXiQd599T80y1r5QFOT5qcb/DWL0dE4OPzmXTtPGXvPMrnfKB
nUZEGEz/qjY8PEXUJFJoJItU3Nu/C47BN1Rtg9lpB15TKy+IrbSq3eS46lfSijg1
s/cLOWZ6waaOeH67eGqlO3yQNugXPuDt5f4/MbYapEN6QwKNYzLoVU8LHf+xt14W
IYOuwMbaNZN4L4SNe8/oqbkfbPCNHTrcqZZD95O6bx7U/8818YhGV5zywwZsGX4m
XeKGOgL0MveWTBqZQk1Twz8YqU2AnzqCEbjH8sdL3pUsOlxNY7AkbyNoOb9I4vFB
ltAreMfLUJQ2IPwcBNOzalYHK34d4TCtNztr1tMONsLBe9aK1Hev+FyHZxX1oQN6
0gDiKYK377IMHzvFd0Tn+E4MAbaH+JEkw+t3i83TsiqhVV6TxQwHmVrPjDJmeMKA
peQFwOtETwzgvJHK3dDzzqRj+Icibq+uu2hyvgdELoRlYWtgdYXxmNhWIy5L/Ntz
5Gz/pzVt3S/USSr8QW13sZyVBzB3rpPe9DpQOJyKq0DL19VXdfd8y8+MBUbcau4r
UIvZ37a214x9CP4W5s+iJpWqyPnOvvYL0AFoX0w2vscS2yhUvQS7u8CzCtyk3Uhn
Uu+ZNnB66Jdw1mo1dz+9ojMRab31Sd8aXryO+Xqs+02PVPS0EIRFhpZuTomySNZ1
f1SW8EtA58YxiCWUw6HhJHaXgRVZty0IsGxSbFN83Y5xsLnsgx1zts0Y64qQrdTs
uWZ/dffxfTzCwhGc6hn5/kXbl076gL/Jn2YwsoJPfb2HzX0pOyYzpr8VrbFfJUzS
yJ2GrJ6o6yTZaxM6Yd5xmibGv9WZb5LeloUrFyw7lTq+WSVhPp2zChzFny7Lobk8
NacxW9kmcQkHdU/MAXy/CjwjPPCgA7wNIHSi4QJ51YOsvDA/Y8ST32v5su1nf3+s
Ij/0K6Q86ZDkNKgtE76hCU40Qtv4BFUZLmVPn/tE8l7NCzfXztq/WQUmUs/T2bRJ
j+6zZ0Fry2ml1XKmki78x7JFA73374RNHGbwCOmtdy2zowhlu/6aqQlFZzwrR7Nw
RKngarxzoJ/clgZjSS+iU/Wv3arPSjKnbUkqon4IaHZNSmIq4gjKxTErmIdi16MM
m58ElclIvxMKrAHkaApbllbtuECRxngrZEpfM/kvd2A4TVz5SmrMOSq01lRqGEIy
iWlDZClxFIqKUIalDWV0tlM6SFGt4alP4TSuZH2K6a2UFmCija6ag3Yu9BbeVKj1
oDR+VMGQC6IzTJOarlnlDJOgDoLnQDJgHfqUbsW48xdX3x0c7cs1HN1zIm3Gskbw
AJw93N/w1ro9w3GGwFQFpMGer9s5Lq0HtZeqfMiSQhYaCoWNoOtsqmZt2zxKczat
l/nr5qW1+4/0VsYk+RtA31cWaCU16SOgpGKHyQR8DMiDm+p24Bclad4SVgXDPu0L
BNJDNmaottI+RoLUwBXXrbuTli1USaRod8Sn+PMC4qyCwneRqBSPruGUv5R0U3ME
ythPSELfo7j8JgAN9x6MA4OZJYGh0veNiqVZcllIrH0hLxQ0Aumbm6ml1xyxtWbu
N/aGsDDbNhG6O5H6QLsthbsxKANXO+HxvQm7u12HQSozt1wb2LEcp5YaAKXm7wWn
PDVeFJBMy57JRiSi8GDVkQdBiEbBsZPuYPeXHmbPm/togyUtOLZU2vN9SbxUJk7P
dxy4ZCMP3PDRKXU6hj0vRXd/HinbGEYh4gZhHn3QICwZOhcL3Vw+S8KEnh1UXFpN
TMiUPKhyyQnOyqQSYNj5fNap4mlDgVS9RC8+oWncvdeHXgSjksmnIf7hr8JQDRry
MrDNP/DmEU2Bxy1PfGlOt9YFVhhtpq4EE6SZh8Yj49Jc+Ej+vjh8RHXn0Wgryd9V
rn+vWwEXeeTtrzUEl02JRCGdBYudBys7FxQ11xEEW8rumf7cX2HaKnBgkH7QEGXP
inoJb/5CMkSs3loyfM0J9clMBcMAprVRXYQgvTYnudzmUnSgjgXi0jFVesm/jAYd
Xn924jjQNIlhRMrGhBqwhRd6HQpgPyc2t8AtVVMGlKx6xIQNkFTe4uHciBth7o84
F5nHtOsxlMltBUgIEULmJREvnKW4kJ+Nu1bobT9WK0ndxSyWjGg3XaQEhzB1/HiP
OR5K6+rpUROIreVKh7DyPmr9Dds874M6Xtxr1swLCq0r2ytmsnger/1/TNp86bu9
Kl+cLC6jbTGg+iELoGqaSmJQj+NWuIMfq/YfHN981RhpxrOWqbDxRDlaVNvcyw2O
02YX3/FOMXl2/HkFbbsFxy8r3/zY5ZL8wIW4DqOfPtglZuS5DROkpfiyJt+COsTc
EVU4lRsk1uwrmiQUJSY8tYZaY+G3G4Fmz0la1oxnZl5sgvB6OrpKmSkWIF8rPxlV
uGQ6t+CcRVjRCBpjvWQhmenTWx7DiO0ubvWHTHF8XD23Z4pBIHW3bMHMUSslRE5g
C8lLAb0/nqGkBchMfMOe46IGcluuAOyXYV2aBfgvBqk4lr/cpgIWacE7tefJtl63
4NKm20COXNsXfVHwRZSHIblVWdFIr8YYMTSspYoHkEqVBRtafmKkZ82sMXHPUczV
yrTBbsf+szIAYUJIkR7N+mgJybuCmlvoR/SLwqZDEbk4dCLIQHn9B/yZUiGgUi1B
xQKUzxoO4EEqV+tCzRQxrs3mQsggteJqhDMJQq5r4QyiCmeAdDF4dL8yxUY9fCmF
ghamw+97JieAtPSpkaYkh+eoEgcbBgJK7qe1UC7VfsiKLkU2pCe034eK+uq8J2Li
6KNkGZbyUxzeaw2EB9Kf/bjbCo/IMWCgxxE86fDOqMOvbgL65ePF2ftXSz2aIBls
K5TMJCvNFWkb1xpa8Ohh47GST6vTOyDpPSGgXkt0dR3AAHtmR23hPolXA/epigN4
fPKALFWy0YaLjfwQWKxlEtEUORkyDbWWrMQURAjXqa1q0/I16HDeoOYtvEx3g1hV
CV9SpYli0NDXNTiz3RRyFddvXAL1qPAYFuBF58UoWqOHur8Edtmq7ZpD1SpN96zw
/HPPxH2kf2Utaezf6TWidcTT8W8CofwCIJKeNaSNLiquNapATnCpwb1R74guxvNr
hijydfgwnYoT+MMnRVeMtFgQ4Fup496GoLOvagatLNSVM/eXhdhxImj3uGLJEiqI
XjYH3T1OpGtBXDj0NfaS8RatdN8u8aaVpe09zT6XEa6eoRuNaUgqvwvlmH87bemX
QTOgynOT4qSbw9sYSSJsDKr3KwJc37n3dbchs7Cm7MN+W8OsFIUqXJExb2/ywcev
1Tv1IuJyDL+sKp62fHvxvkLPbLzk+Js1LYiwRMK5z47qv4ivMJZmMkzNGNITFIOM
Pb32pavRgHh9lyCz23YpfQBw5xN9PAMjT0H6NNMVvKg3HjQExyFOFGOY6FuG++ef
m7ITAn6OtSj7x/lp8D3FNP46DRpPSbcTUMp8twTCmr5M/5el9v87NaAvqBBL8WsA
8AsBJev7A3h5kB0D+BSz0sTdPSLDc5GqVH+tk+gB9ph8GufpPa9bKglkRGgBZqKq
QMXEsCqjAFesEvSMrBXOPJJhP9mjvGp+pXMgLJElJdjxROhknyQjc8p2tlLLadBQ
B+Hv9kMWcasu4Lz9nNUh2dCya8k5BdVvwgO+QbbLg5eg+HejP34eknrPMn6yNv2j
81UWz7sLrnm3Asb7xEGMPku/OPl+xRqj8Bm+RSEEilq/R7iOu5sM2DRCjjG3pG/F
IUyWKOJHwKdI49wJMDR3NHlDXfX855pK5EKp9XZeL7l0MX4IdkPaXUNmgSnakK+v
Fnut0yBkNtnpcIH7tMPnGrOwi0dt0evz1Vv3zGv4F29qMaGG/1JEKdYmNcuEprCL
bb9yZGVV0ZOIz3CpV2g6qWnJumidyxSEkMP7OJWF57khSParX2UBTJvnivSq/asZ
zL20gY7cr9QudhyMUAn6sQTKVeiaQRKPcWelU1NgXWd76pOREbVnvmD8nLvRI94p
EfMhNVQNM+RV8p4bAQvec0fQmWW2+y/LDr8ZpbT9G0UKelPDpJpW1ChKKc1L18xg
RixKHjWGy1zzvToOf+Dz3w==
`protect END_PROTECTED
