`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H3yElgWlEs0fKJptYT0g+OobIuJEKvtynw8i/jIx3UVeh21AVacDTor3m50835sk
vMzeTn7tZF2m5glfajFgxTJvSzaaT+HadWwvQDqPE9tHHSITgbmnYKBPZbRBkJPA
Tci2+2RLcL8+30USw9fF4ZGtQL51lpT5BMrLZ+tdje4lFkBonbJ9DqbsuVxdxHNN
oprjcl80mYFVdrzQaMNjU2gSJG3XOOIXQb/Ssqh1mOTO1WU4w5HCty6OqwPeCggH
erL009ZeGorp8c5UmHT6nb21O9Pp7X9m8hoYQJF1k+h7NrMgkKDkq5XqCn6yzHFi
ktk0YTjWKPwmyiIZ1Vj1UjCGm5pFtBYuXYp0FI8gxlXck4JqoLS46kCRzWJDc4RB
wutk6ku4uYS2GFGeCzmzMV4IKLBD+YK+fZmhtERUu7kOrmMhYQMyFwCs10egld8h
I6tO19GjxV1GEf5VhGbDrOlqYglEFpy6A/we2RLVksszHL+QRu+9LUuY3DyVaDEn
svoV4nn5fOK2cp2ClkN10Ztvd317xxwAQqJ8FY6S47Pm6nVda/vE8t7p3ZQ3iC1p
jhbkKkzjFeCYnQFL4ruF5A1XA0n/k0jYjwBXKw1tDEoEYnmstnJXgCZ+S6sUwgna
Qrn/3GExw7qw7JonznhU4rUqRXMQOeLQ5afJ1hp06JOJnfU3mc1DepGtVdzSARwb
NOdH98XL6SWI0UGSI8CYFKmCKLHGR9ejEnsvfAhNDQvXKq/inzpbNq2ZPm1st/YQ
0Se3qmPqYhiflIhRnU2LwL+fVREp9Olb8TXtp6or96iPh34TScpul/YSysdRjqxX
ID7Mrz42UmjCQqzC5XSAO5GB+yCG6Ca/f6VeI1AyOQhJTVXYenfFervXGdFjPktR
/NOm56lqMidx3hkQbua0+Np0BEwMrs5J3yeDpBr5OXJRDaSsKYX8ccLMSWOkLBWd
0oxrzYfvmv5pX/FoOn22hJni+Q1TxfS2Nj8r+UfKplRkwlmvDjwis7ztDweACGCe
GCAMaS1eNlxFGltyeMqtfTCC6sRjMd7VheNhWP4NOhkjBqxk3L5ZstVpKVcYV4Gw
Zs23SDCz/g2b94sq9x435ZA6WoMqRLFmmiRNLdIYIrCAe7esja6SFAd9r7wPVgaQ
upYgx1FGcQrWtRqemi5JG4h9exnbNd+7h/9GScxW1WyLQyQwSjX+bpJvIhZNVuW3
7dzhXnoTden7LALUqHgJlfVxTY4qhCMekpIPAoIasFIQLTCmq3ihbgaC1IPlTi9s
unVwnh5epz9XWrJ0VfdDySe3+a4KRvpLOSgIBd998y2GjBFfyditm25PraxdyYNe
AVKaxEcanNW+yklcwC7QwhIE/UgfifFSebGoEFBv6lJNJL+MbeZq6GP22KXw3iTx
zDJQ+Q1w8SQ/NzVlJdqX61ic796Jn22arWXP3cPIDGwGnJkkGg/R4Tk8d9NZR/qG
cw5cnCEiSfBq4u+x0nTRFrmto9r1TisBAsQl5DXp66MW0K8DUqTdovUtQtErdi1S
HsQ0yX5VfFT9aFRY3C+YMeOem9+WDLwYeT0R/7p6ei4=
`protect END_PROTECTED
