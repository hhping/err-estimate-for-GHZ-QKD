`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vkUR9hY6l7z9wr1kAsFX2Yftzodb/ssxCN57OpUEPxXUikwJKnsFgjMnmMxc/urs
0vdwNaFv3g3zuk8hz0lWvPUW7HpWOIYsZprMVNdLEQfAse9vwqYNVLqROMOewdrm
G88xHS9ddW8aIF8vEXojryhsRkAiG5CcxwSDTucFV24F73kepncZa2a7evvp6bCS
oD0v5j2pvD3aiAkB3GieXTJaiUnBU6i3de4RusJ0UwxTzq3IEkGhaKjuC7syPASU
QcimAQ6OWyjS9ivuFb/2Ru9tgYPmW7VqHkZsbDver66fSFsKqYoONb3SHpPVOjle
O+0gPfRUasAwctjXjbO+7SeHNODWmI8/3Fuwep0qJRCPQRxwsMrrs+kokU2VRxAU
G0pU3/Apme1IPfVwxpuHdUrOC082UfpNjIrKB0OZPdQ=
`protect END_PROTECTED
