`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5ihal/OUBmnMncIp3MNUPjP18b6d9ST3AnkYERLWdH6crmk3VDLKmjQcc2yQpPGx
0pv+zWTUDMq5lpQc3x4ORStw47MPaOGFz8tEfJAkHkkCRfx6njBmIThrYN5XUBfx
Z/p9KlpGPr+t4O73WwlU55Pu5RK+zz2R1G3lFcXN6aXCgEiNZRm6ml9fCf4bGwyP
Mz0jw9b86jZlHymYpP+x/igfCsIZgP9npd6pRjC1NdQhjbZPwgp1F1Wk3UP6Ngiv
29d1s6i/1Wtjero5s80olv5ikuCy1C3YJNtaVA3ilrUEbmSJYQ1wV9Du3TFF1KQ/
4CzAgt/K4dYUQ2wKbB4D2CPuvM+aNK0ELPm+8PDjknE2pdg0nO4iRXKF/mbQvgAT
gfyxZvGuGqqfkqSgnWuAUiANl7hibWqW1wtTZ2MZRMfTy1OuOy900U2ZwgXm7aq3
f2yR8pj/qkL8DVWSK8ki12MtSjOOK4kzSnXSUCCpmjnsqv7ysw2v2KR87Qvm2iy7
8O7iDMSBPMDB+Lb5as1iqcaPauzjFuWG7SC/mckreXNNzB1rO54QBAHNxL3ePqui
SQxybnLE1rSY3sZD2MT6w8/WVM5UR/q7ifsI3+EY8qSpwslAATjPSa+I6Vu+v8E2
2wlW7mkisVZg7DuDhZWX865xT0XoE7mJNYLCjnY7aqXP1OzturjFLhQtWQf4uB42
fvIl+eFg3a1HCxIAlqYolrvOGfBicJTX+eyJq88PN/Af9KqyzLLcLanGnQ4gFpMG
EhoBPhpIR6T3x4UIqNprMEl8ei08qKi0s+v3ZxaaxAoyyNbrLLkcjKABmAb/5aJx
EVfb0ulH4DAF6ctxJeuInjD2ltr5FLG4hE9GwwnW/xeV19iddl/ctsW3xYQ2GXiJ
J1GPHHHIhQktDYlrwofeQgZWu3OrePrF2HT6NvMBw9DYWvinWZI7VRsdzaolZw/j
FlWiWxksgd8rta2OmRa6bh5NUtjk/zERDK1j+bCNdoSmqGy9jpJ5axENuqbPXaUw
1I/aPSbtRNCVCk7QTMCu9xcx9KxnVjLVUtsRnvT5gZUIm6fMOpAODc3C43YPC0kc
AeQu+NhJOQOBl0PUMz0wKE1ual+AvKjcOTac8QpqaPK6RxJKBlHIlZ7qYCJY66M0
LhmEa4B6u6RtygBno3p+6TbyAcBzXa6a+ZkbQD1cayIIWcpYnDDacKKgvh0a+KC3
zqotDEGMW1q+Eksif/uRZuLE8Jro71eAcl9V6VyE90hKxDZ1ZblW0sX1DqRSxZc5
PxD71zAGVwgX395rnrt5u1AS75SFv6xZdIMmTq1X8F32hHUUwQV0fLQj+5EYnzTy
Vc+rVNdZ/RYT5aEg3ibP6pyyri0exKegCRGpbTIR1RUZRYU+FXtoOXloR9o+vVS5
xgsIjU+j4dW1QydRbT0cNyLi1PS9rMvp8QnUPcRzabaJpdA2FpCPDZZOzuw6hsXe
+Ccug9AYWqAe/X4fYenId7lHImglsyYD7Dy56kLATsjvWeGkUNTgw8Zd9Z9AVBAE
GMqIaS/UgFL7SN7qQPpqLPSSX8nVUS1gGEdPeCMv+NSbrmRpwKVtotLzl5flj8aT
s2N9F1XWchg/1oi2W1I0T3WJY1KR9qTgtidXUvD9qghMAdSOfIpRMQe0B8q1B23A
X4xW+E1pDs1kIf3/bzFW05iC5ZE6gRmVFwWHGXm+sq6QZOXMOMfBUvrcAMdAF16M
/9E+MF1q2aKI9fpDzxnn1R/ymc9MH4Ewf48gNKFjJIWTrOtAbXhyjgppWOhUN+G9
DDhJuDu2tihCgj+8wuWVVsnnyF5QH9f5DAPneizbTxrba8rQkyH/wqMkCOxhzmI2
IZj+PRT8kCrvY5CKLK8HH7ZQHcmiU0OVBzicc3LLh1sgwFu1n60LlXUF7NYUMxFW
4R9yEbexekU6+vCaFg12+IzfCLKWfRdSGqmIaE/aBC2LEnfGARDia9cZszr0R+Xc
lLjXoe2XDvlgsD4+V8kJCiJMEAx1zzwhUd3uhFeGbDcw5KozhAzO4flsngyggc3v
1UeHFIFxgGNRnjS9uF73FIcQ75oMjv1JJdCVHQHGHDbFO/labZ2HAMTymLNIgPA6
`protect END_PROTECTED
