`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OcU58A7fm7W47VuGk6d8YtHfQiwzBOx4Nw4h3lX63QkpOfnkqCRHkDvaHakTKQJc
+W17K4XEY4XXaT+vTHDsSvabHFX5ggmVLtKjoSQmTjacxS8X6w45WV+Guvsj8KY+
BWP0hhcbXe9lqYXsx8pDp2v+jhx+dYHGSFLOmKsXFdy07QyypvHQ6Sx3OpOnncCd
6f4kXApo41d9OyqcIgz/wSC3tk+XgOqzoEXXJ+QPOGQiFPd2aGYfIYIZNDXKm4Si
Q4kM7E3CIevOb0weZGIo1ZhqlgWdJdlM9JjHeO2KI4Nd4MLHZaERPfoIMhE/Hag+
d5GEgyAB55YWFB06NeNxnpJBBmZX0Htn8zTgHtEdNc8Yb+du1ILJ+MdQ9qgoEFG3
CIajj6RCeMFFZajGFsaP0Mu6IkgXGO/a2wQ2fQlAYB+97iQ2Jn21P0W8i7pRqgR4
1Uj2hBIJJNZ04/7d/yfwk1ITcNjc/QUV+phXZoCTpqzxm4Qka3gSZ3OtxLYXEpdy
cw4LNtb9yguCnINEO3pswyYQlHe/2HdOW4p9CYXa9sbfM+RzpWXOYQHB0FAJwXvj
aWjRE3ecSnzfNFVV2lAxv1HbjZtcHyL5fDOaTumsx0eBx7oUpN2EUsPvD4jRw3ph
hrW9JKY58no/JUJMugXarA==
`protect END_PROTECTED
