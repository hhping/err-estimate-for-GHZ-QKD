`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R9Art0ZvbBLEfIKSjWXza+pK0IHVZ1miA0qWhFN2dld024JhNO685kigED/lET23
7gYeL2SK5BzXLMKtlfiKgjzK1wohCE7qDM/bkqC0L3cInngILrEV1lspXA1X1lnh
xwbj5QQ0Z/0+4HTTxY1pp3/2PW8gSrsbm4nfprpPDioPmaJjMDg1DvXl11QuNoR1
OqID92J9SHpqmfPOoemzZnHylz63xy69COgObA+HnWbRrc2fpoeEepyvzchK80in
AX2673B27HUyrCrYR4tQrV9UPcXj/Y6VEz1JyAVUiKty5xjWKAZD9jp+49aLzwad
1VaMZxQkyy8KYITVM11/TI8SMHzPURtlzUJFAtqz7aUmODmZur0tqKAigp/0wUOz
sKWG6WYfQq8iBvP6OWf3bg==
`protect END_PROTECTED
