`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4gvCUi0vkc17MDIJEEE3fgFQkWO77ru7Fyiib/qW0nqQr2g7J461Yd8sNo/I8cFW
4g+wsiDu28yER+ncF10GCedT1SsTGXBGcN9Ny5zLxH9Q1WhP5hRWUD/74Q6y3y0b
QEhbT2anjzAFWIePG8oP+1vWThwCx8EhoCl6U+60iiV/qkrh7X3mG0li8kXf2SYn
Cn0Q0GKLmdvoN0+FnRosNxJBD53t24879lHI5pJeAKV+/KtFVf0SwBqvmaGO+Bl1
K/A3dNnKilmEWx9JhDhjpNNIb1U1hOMGaz2OukKaszcOD6hTzU+74cVYUQsMBnk2
hZFVZLw/whsgRN0uFCQ0N/BJfJ5YIKweniLy7RZTs9Jq0I5+5+KGcDys2Ns8CVH+
+CYxckJyDmxkOoIo1Yjw4+EX2sxRsiz3ti4DacyBmilEWGwhQzyc65t4VwggwxlF
WG9i2Myf2RFAW+UoYfLizKB3r7w0t5hmM1qiDQ3YrMVZUO9g9USzDxLJ1+ecjYAs
CaPDNFu59KHAWXPGUtBp7yaZJ1YnCibF4TsXJ1ng2dFMizyarJOhGNni9tu+azfx
5Q9zTIqI0QI0x7Nr7qN5mYpDCYKYQ/GtjQsAq1jqt+KIZHBRiSu8NH/Xy8CpNjcS
QXtP5gel1bveVdW2OP3etQ==
`protect END_PROTECTED
