`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HwkcTvrnxXceTrS45RTidQxLixapO/tJGeT2jiEckI8Gj/nkFZklwmuDYx4rxBTz
XTA00mKfKjV66a1wSi/7E1uUyYzD6rF8AlvAhUeXWwgXb/gTddiMbOWaynjYX4hm
cp1+paE+RTSz2fTilg4eFKMDD5/Cjtu+eO5UNBDCjnNp+P6jolHySFTbxZP8OJHi
VHrbKpobZFwiGw0AsIeweAyUQ3QPEhHECtbeTaiMsAakNqAjjn+4KrlCk0t1UBd2
C2UetHOZ1gLcrsC73d/kkHgVfRbekTKHv8sxDCFFoeKFFdJjZxr7U08XyHRFuCGk
jwiRUAJ83d/EhvTmRHSlryriFQAGj3dm9eganj3phEgNc4roGFbBTNW4MMYD/Kdx
kEG2SAuSv1XtgoGedfa4wwB7yISfLUd9w3CmniKPVRTt2iJNjCihMH0PlkF2dmyd
DXUeYqUi6A29/AUv3NCqzqNWkvOH09jaZ5dhDAv2kyqbd25+dyP+mE1Ekr2cHM9Y
gkS3vUQUfB2LXnZ0b3q+kA==
`protect END_PROTECTED
