`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AB7w2Rh0/TrFT3OwNkGMpTFeZb657VW6EVbCH1ilVgtzZovHe/+H+K1KGsv+YPAv
wrsAsEWujPV3WdE29ubqwZTcA5HfggQPtGSwvL3Fs6IB4pQQReelgPbOgkWFx4rf
FpqTg7mMrkHF0VPhEAvYRdNQevnPSP1+jUvxO0wYOcCspJ1EhfwvNGBXgjeZ2YUJ
ibpNxOKXmALIYd/OxHltOASMoDDnQZAadlPKjD8y+1DDN+hf26767JY/nzSVuA+5
EWN9FLD29v7UuW9P18cApZL2DbQSzNw++y6ayOk2S9JrLS/epsbnEj9MWbyrJjP1
rDOP6n1zLyDGeF5Vo30IxaTXIGQWJtMgJK0BMibPgeRVN+rH/isDHve3yV9m27pP
jadXQCFOiKkgMU18VMeaN+JVTgU27bUqsDWLundXvG0I1LS61hQgHZdRRJ63AFE1
EJ+WuBJrDeF/eNKfCabxVILEl1mDGIXfkHB2Fh/2xvk=
`protect END_PROTECTED
