`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/tDxoZuwMYe6jiK3ZZAZh0rCtKIg19Ez1ampps4ehnWa2W9yWyPclQoadgkx6R//
us4d8D99IxS1lPstemG0GjamJHRF9z4yGojzK3JdIfSefRi23t0uwNf4VlDf3h3l
mXi38q5TlpOMmvR3bfiSh6HCbk0w4DGPQ5q7YbNNgRHW68qyFMsnaS25mmpfOiqZ
1bvYO+7Pq9JRTA3jPYg7Z9W3Brw6zmRnuVNNZ3qpXETyM50q3hfT7N6UsgtYUSGg
UxhLFw3DRjk5F+gO0mL6CaT5KQZFi0dGyiu1vkM0gzrJhmWNe32K98cedGzhplF0
Fe/jAtn2RA69eEOvjXVyUhg1eGldmvw8dODJCDxk7DEyd/xRFXW83cS3JFwb5Sve
rYG3lJ/N78kdPehUua3Ed98N8HqMsSO4HZV3FAANWYPXAQ9SUk8vGfOHGkaaBc+6
cHRomut79DWdyMxnwOs4RhxLxn0s/S4Jzy9a98S4n0X4Q6UwlLqjXzWLNiGnXUbR
`protect END_PROTECTED
