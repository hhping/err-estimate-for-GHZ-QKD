`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J4t5NSMI+UqMJ9+Zp6N1g18iKSYMKO021lujQI5UbvxK2sqAmAfgSjB6v7zAq8L7
Fa4MhlkRsaNq2Py8HZRX6E+tn6gCHo5He32dVSJ6lMhOaOINpKplzWuOmNL2z+uH
uiPhK1Ga4DYL+ceLrCUi/Je8LOPSEV8JSc+TvA7h6VxOqfT74lbFKelpU54x9doM
3rdb94dgRITd5F+KJ3cqC63i5vv31SabAmHbRvnuNFbIk1JPnvFt8lLd0Wqv/NRX
lfOTO/0iWuXRHZjOqRMgo5PIT+GB1UF7vAy5Y/yPTPdsk40qIfo36IfBuQbIra4B
zswbzMIgP2j9lVdJlWbJ50Su4sFuB2s3ndMOwi7KiDAGUZAllN+pE4Pzm+B/10Wl
D+pRoKdg+2a1XS7/TMJZGnOwkAT3Y2rhPVvyzIJMVYK5eGaRHz++UE3X16tdBspE
Ho8ziDdcUbEhO7nHVFsbYvEKB/g0pJ0ks6GDylCOs8MCvS5A3PeZA4OJzrXtwuZc
UrQg6ebQ7HsML6h3xu5lcozdbLvYuzKFeAKCdZB1O9IOxz/OUCKBD60h6Lu7qyTO
tTfe9v215FiRg26PAbc9qwNV3NQAPsnenwbft0eX2n7rtdls2qe4PGkZ8/guQFht
Cnn8t/i4K7J/+NDGAB2kEZOyowZ8qQDYaUZwCLmosPXiHw3zayUIX5jM2iBzelY+
dBjeiQsSUSg2rQYrd/w1rU7Tmht5X6Z6kQsBAudT5qWVWOU9KXo/of2yyaBdZX1i
OZX91qwOW2zGagMUQtOXQ5qkx8OAQzC8y1ex2GHd8mQiNmCeGTGACkfJMnZOx/ab
2mhlm3d12w55Y5gwJPAcoyTuKXGWQx9Yx1VbpXiPsMn6Deoryehi7ls3MsIqJF9T
hhvSML7GtyJYy26cbLgKy4qH++ZLImxYVshnvvMNWAnBPHsF44Sa3K5FizivNHRx
oZ3jUj+Z2qDr6yp2C4KSGKq0FGWnZKxKw9BJU6/sJ/0NyhL4r9vnzcOjSF1rpSM6
Ea0OWFRzmze7jhNjNJ7/2WKntCro3aNdAS4r/rLCYWVLirEyxRV53GL7YzHqjST8
5HLJAd2/r9SjF3Yz3dJNb9BYteBruPy0+EPTfBb9jd5U67qI9ijbkSL1A+mO4BwO
rzQWGQ3eQHgKWSMW3i43ZHG2of3JJV+kVGjJfpLIFkSp4p5QiEs63g/9+5xHJKB/
QJhA4fz6oSM3a9TFwFMR7O0hoRgx+coIQZ76gYPOe/b8oVzMgnLPwm8CUwpmAa0W
bSnEvjq0XjnZUWYnM/YarkTbbayU7YMyV2KBZ9O991jT6E9Z8udgmE2pxGcdeqt+
lk4kAa8st9dcGiltaoAJfNQtzVjJEpsrI+tgMuH3Z0zgds6gMmvtqjI7nGvI2gr0
CiSXjZwXZohqcwSEDExK+b2LQsCADZahAf8qnvD3aHFi9ZIHjebiAoTzx6tkRDDi
WKwt+PSnrY+thR17jXulJJ3k6uPi0fh+LK+rkr9BhMSPpNNq4mWSBEcSxfiw+vNJ
vws4GTuYXJ9zA6uf+j33mBUFiNHZFwUGXSwecrFC3npo7EklJXiCMHq9FZnYNWez
Gub+pHa+qPaXpalnP/wBHJBybyss7ghSiWRVBtlMGs6x0odqEGkhFxZtrfbPLCom
NzEQ+kpr00t3SDC1bi1hN2NXVa1hm5dOEfUNMyBctNiSUPDm2vgk8VX0cAAFCLLI
Iaq7SDPvWWj6Eco8yxAEKgMkFu9CTgy4cYsNR9EFEzO6KcizZCcwhwsvbRuUmlb3
zVr6yKWBRQy7yOCSmbsWHALff4LVa3Dtm8ZHKYZuGGeF/YdMBloWgKwxlQf9mhJq
9IlMyCX0Iy6uXquWKE9xrFy0QJk8C0ZW6xIa6zmI4Bvh4NbuyKvyqLy9NVcj+h2s
ad2JuCW4qAWNJ4bQEo0yRAGeOB6DYRfRZ0Oeaqr9efBUt/NLc8FzErOXo/s7rk8m
9cYqaAWGEMif5SBhaksCeirYG1vgivVH923dkI8Mu70TbZNNeD3CEjmod5t1cX52
w5hBRZfDOKK83MfZM0zqBlMAmqwfS8VPBuap/spA1Mb7Yl1ayjfhL+BbseL5I7lx
umN/Y/9T4dSCRm0AjxQVkX0O12dsrzKQGslLbcex0HQBFaSkpo2BkloBVi7wwAIo
HJWkZvcof3rwsUL60WdToG9z9RqdVeVPChWHoaHlotOK08tAhszK92vXJ8etNO9F
z8SaVpCXyrldfNM9fk+KZqlYvIM8NROav1SyNSVGtAm4MK8hn5ep9YNEKvMFAzJO
42NZynXQeMWOCVNtPFor0abxFtuCkKC5QMLsyC+6bX72cQU2Sg7nUzZb4D5m+P3p
V36TvWgVaIySuPCPEIYA29bdOOxA3r+KztextajI2JAkD8rjprSIkq/MHhbuWR7s
YBKHfTL93dI8Xg6voTCKtuq7uUetk1nxC3rC/IxTlg5wTj6paihQfTAAkU8Cso5B
/D6jyROAPhHowt3IkCH/k6Mtmfp1JqpQTIuLjG5NevfjkljzU/v0NmLwfzzz3jBq
U9d+YqlhByki8IGpQTnpEixHhjhZFmbHo43J4KwSQpG1tXgwMyTIF+e78MtGhXNJ
yk4BkX/O7vCigV6v+a7wLK2cdOVmHbgd/noMGJ7Xabvl42iDsAe8r8AlJy+NVbR4
IL1iZ045l0KyY+rI5BoM6BvEuPKnMNPtYrOxXAV7YN77OKV8v+gTF1oPpZKomVLg
CExwIO4qVb0DNpfOXWoJGDaWc4HnUeRkr+r6SuBnIU5Q8TUpB0nfKZLoH2j5Yzd7
agjdh3d97gS1QhOo+LtjvOjxCnNbVMS+IMl6ToJXSaKdSfpPjBzr4Slz7Ei7orQq
oJvKueALSNqNJCJLtrnpEmH/x29mjnRZcdrIIw7MBClkVyDOL5eDD3rhc/pExb7L
3UxfKLckz6mkMFDo9H/9kIqCi+1s7NoYuZAcWYiuIPUOxdfYI4Y2xodf3ZkPXrG2
C5BLc9LiJgcAwSyCIgY90ItM43Nb1240605CyPBfqnOcT/H2L3SlzXBmzkVRMbgQ
GlDKZZN3Rjtic7WN0GAe7vXMxxjeI/mx8IXl8sRCEowEeUngxptG9xZee8MTbCNM
nmAdJ7LoHLxN7/Oga++iFf3EqjTdQ2MzwUgCKDCLm30=
`protect END_PROTECTED
