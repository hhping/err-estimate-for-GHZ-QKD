`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6msJGrYLov+uxtU14jtodbcYNXZLbqSPBBGCqMEuQ+RfA0QDF0kPdzxAQp5lVdS7
FpiLvn1WikXb2PCfLoMTbsOHNpmYln6hByVIaEa9bZzsboeB9rS2T/lIQP8yqsq9
GLXGF+UTyHTViu2F6EZQuIXWZA9Mi5sQW6ikgBafsPVVhcV3Q9K+HPtRO41PUa5+
70UO1/+TaOvve8Iki6SWCYb1eniYStypzqKNTMML6FxXntMkCdaL9nvZTEuNmYGh
eWuvayAsXH0Ibo0DpNGuDQXW9xzodY0diZFo/BNM6WP4KUghY0T7++nRKwYgf7PS
xbmUX4sgVL0qSuqpJFL+DD+yM85u3DqILEO9Cs/ZBre7ZDYTO1lKxQA12+r+U0Pf
ryzMm8eRBg2tWh+g8jm8QtG6Zi0Mko9rsLrkh45wSgXsW+9OfMJthiIsSibSnVsq
YtLJIIi8f4aO5cobyJo5SzJVSJRbYY6i0g6kRaRDqK8X7UGMC041hqff1XaUWxDY
qneyJacyXCJzi22Mn1XLv7igWpjI5VHa+2TKS2NBZ6jkH+oyeYx/3+hR3qqXgND4
d0yHMolkVX5u1RJIOSSMb2dX0JEuDiZVNNul7yJ1A/pjFwPHwUVU6W7AOPeZ3V/2
w3ATMI3ye1pR11svTiSSKq0gJiWsbb/5dYD880D8JV//VcbuVEp8S0LlDY02r5WQ
fKhXPeUzytpCc3kxr9njWgBFhD1VSotw3KTeiE2gcbiR93Ij9XyUnjkuRt2H4oMF
90R8OS7d8yKCurt58OwUoT/7ve9DKJN93801a/8IynJ+bF4FzA6PhOtliAv5bGil
NjrZhhiJFhMllpH49G3IzXWcx3KOugg7rkcd1jmCMxmam0AoqaOlT94+ol/Uz+DT
fWgHnfqAXKhbrRMnAgfHNraYRV1dmr/iwtxyQ84a39dYyDDDGTxrABt5jcl1Jzkn
Pohki3ANqZIj3yVCeiKTADsA8cKxxbqHan2Twt3opvx+r/6m0JwJ9bqWSph8Eq5J
m/4YD0OtJ9xoE/96Yx2F2V57UMvPKVll6wRSaYjJcsoqPWIjU918zWjY2im4j9iQ
cglPaHmVbfBcDsNOdG6ciqTnBgXIMdGckGQMB4wOQjQUxgJ2NyxB/irTnqOc72Pr
PrE7h/GomLlglqZKC8g6tDS4vdVZOgoSD3JCk9ZiKbAFFPszJifxjPkrP4bzU2EH
awkUIg0i3PHJw4MaG7vyA369FZz4v/GnRICqG+Z47+HJlG5C9nQIVvz2mG3Xdzfg
0MN9dJiPaUq6br4+C2mrsP37iRw2tszOw0Vj7QJ+JnXNT2xXWDVSpjt3ymh6Hjbp
7a6hwCwC66/in2RtUrjrYkeGdGVEJTSCe3jntezwqyZtIgVM6sif0w47R0mfUcyt
PZYaFDk3ghxM+6RpMOvhaxIRFn1ThX0XbCmjuCnmS05Hw4eXMA/msAXE6QcrH9CC
ByvTL4KY/80R0RJCRk4CQ9uwEcwdwgzIQDT37OvEPpOGogbB7Fjd51rSoEhdudQr
v9j0JZ2tvK2a/Fx+V0SNcupgNZE0Y58BvDHVdQGeUrA=
`protect END_PROTECTED
