`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S/q70CUqyX8ecliB9BnWRm4tjBldTr/IZbbAH+XT2Y1SoBrV0J7512+APKxBX+kR
i800803ymJS1ICl2wlUvs/oNM68lCuKYXdZzFgkd55/CCLFujORh1bEKm8o3t+of
vfT7Sz7sdzgr9H7YxXOoeFxVlqGpsnRxrcCX3mAzZI1EdkPhvi6J3HQX0W2KlzAN
b9IeHDP37XGKHUz7+hY4+Ew7wH0Rass0sXJiYzQV5ZyricmXNntmMVF3qeNGD5Nz
sJTaAcbHGfq8jzvTuQqreZCkB6LtOZ+7ICBkRg9bmaJIzOthOu9NFgAGQNt1GFKg
KAcVFYzEdNPrAMh47B1VErCPKNzb5UjyMnXH1w1FrULLxV7AmvvrEBui2cI1NyjN
kcRHP2jOE8Tx3YM1secK8cWwOMGrI7bRCZDUqyjoMyMAHKtii0HCusZvvGHNngBY
c03WAFg1KE5cXKTZN/wI1miVK4apU2CuOBrItPvFJUtVwGxyya9+ATgVa5SFxLgC
MCArPIxDfQHCeB2dniYCVU4IqV+oIgMgNbRrDJYq9D/G0SD12TTSFf4FrOspRoiA
`protect END_PROTECTED
