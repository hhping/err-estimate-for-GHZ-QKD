`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QtwwenNL5+rwqaQMPyjM6YSZqIDdTZ9LaGiewtzXcMKnPxPY2Ygf9xzAnlydJUip
/60/Q5Z/NzF/6GNbr61tfXU6TXtl1hTlci+vzOTgtwThUyRmRxPr/xtx7bxrv++L
U/+cnQ17LqrwZYEbD5FGuIZRGXbc6X2iKubR730PXOALhrRtDqOB9EzmfD+zLJRt
vpwvOkw+UzlsmKGJii79ZhmB4IzlcmxGUUzdZUWeEDofTJcall08IEPWC4PP6o1W
Vqb4meSO028aSi9jbr7wmFxlpH+a0CffIM2H4y0qic4HufXj1BhDSQrJ8nEHMqSE
9kZYKBBQcdnJW08q98+4jVypdRVuYYvptMMUskrHOEWk3WO6cAiZagQsB/H/uNPP
CEb5gUmazdRD48BlbdablEMd++gxKhamU/A976hKycJUq2zKXucSioIlkovm9EML
JT6j7NnYdsJCweisdpjLYRGu8h1uBZBM5BuwF1OsJwVmq2JTBf2knv5cHcTP1L+o
Pdm6usuyclAXF2Lq7xoz3eC/2+qUyA96Tt65p+tynh8v7VbegIetPdgnuHofsUuy
Y1GV0+CpeSv3rfNgDz9IB5I8NuH08Mt2D4hDwoo8pGzyvhi0wHMLetiHlrFbZ8bC
IXR3nM9vO1bz016x1/oPAzDHoXlcrCSJZZ96+wlw8EvU1b9opaKjfvXC2Ci2PO71
tVmHx2tIj6+WtkUAN9eHL0HvgnVV6PL4r7bGS6Ug+XI3tMeOcc/5uDRzi7ZENd8Y
6DYghjydlUR8u6Y7LHewN6bmLe6X6znen1cOU/992yZqOlLU695jAdsy5ZtSIQfK
XgscErcvDQu4A+f01c8nr0aPtJ6RMD45ZH9VEG9zCDjjbb75m1tyQy8t6DjCFq44
QQbj7WVWqA3z76pYk4Dk+uAq0mkbHoiFjTa47Z/Z9p32twmR9BT8mglkJ78D2jNw
lG8hQFkuI8T6olZyjuY/9J8mwcv90n72d6oT+io5ZSusYXJc0SlHsA8l8DZ6OsIF
tTYTmaKYIroN96iErqKl7WahcImhK0CoBohl69xJ3a07X13C0s7rENTO0MtiYwYx
Zq1z9MpWUS6fWhITgrUI4EoaJouHBoT16f4dS7z6waxhiYFHKTH0bPZBuba2Bv69
wRA04JIPkUVGXnc9yb2HK7sn31qBVs2EF3MZi/TuBMo51bGlSoWigLiDA5l4IDjk
iGHfEJ6K2WgBCBddGTNsfO/Ic9zrxNAcQuHSA5/vuRnva9R1ON9ggGlfRhj16yEE
a5KXehF1+KAg6qHABc7TQJjUVHfFXd0JBxdk5/K54k4=
`protect END_PROTECTED
