`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lgrR+5Rl+eTQs9WSSkGk2XOAjDytpWpl7Rexd6yl9ughnTJ8qlxKIOT52C/BI1a2
M2pEugItKoTaxImV8V/PxX/4JTb6e+SoPX8IHt2DPF8r5RRBwv6qS3Ttg0Nunwv7
kH69awNbINidf5NkIzSw5eqEI0tIMTrzWt6n3SikO6tZyWEYMHq8HMLnH+1rPxxY
t8nxVA9IBqcqpOP6gu8Z0lCOLEczhI/p9RpusApqnOGJwRGNOeVvXBBqmsP33QMf
/YEC635krUo2JKkvx9vlIjmTo3bVL+MG/7WlSRQ19m+Ka5ybleuvN8dKiKmETRla
8taNI3UI0Bk9eomvAT+xOZwg8sQ3KK8mLb/2UvvlVcv94t7ELMHJv7yB2sukmDsO
BxK25GJvcOfqU7zCfjy8JOnZVIoxGIWU/CrQmMy8bYmI/7aSsdroA5QCQ6JPsif+
k6pv5aBsL9/Ka8Jh+bn9KPeypdWda/rsz25dNxG2PCERvTPUbcXrCDcP0uPmkgOu
chjP3z8Mxq5BishEHRpzQ6EZYpscnCiLgAjNDIUy/5dJiVqrKkkkx3TvWVONxEz+
konwN+usb+zabYzDTvJrxoaO2ZawIvUBaK0KRjiSrzZUWJPzwTsGLjZraOqjcDZQ
PU2q6PMD6cik1gjlvEkiQ6mUjC8gXI5n3d5QSqOZE54hAtHv2F99N4mwtQCLQAUT
bvYtopk3IfpKrcFhXchFHxWx40t+hLGFCH8nnYtM6qq1YAQFh8cyHIMMIElieTrz
`protect END_PROTECTED
