`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GEGvYnrqw8Fr019lsYgZI8VG8BoiN/rOy7VCxO1pJzTBS6qTZfWBjffB3NRCt3h+
moy0e9N/FekHeWapv7MMsn5NCKqtH+olmjjTZwahMsjiDxmJAKO++5mvaF1YoLCe
1iaD7ItXQJWiaS6ud73D3ckr6wN4aQUhSBS8bTrGnlQLZGDYOx7Dkk5F5LV8NEdI
LSkJWUUr40cZr4Gz4IKhsKLivkvgG/quw378lBOmpeFDmgCM8AoE9jRsCGTF7clu
opmqDzwuyt4uSSzeYgQCQ7SSZpgmeqix4wozk9gMr2gKx5RTxmZdb0IL3EUsmG3Y
401ypUkwCqphBmySXZ1cLsHUE3/ltwrzTA9kvJN7uEUJE9fIVX8FYEj7VwIbpVzg
aNqxzjln7yclIGt5tqbawzGKiU8U90iwLk1Y0xkJFjT3rCalhVq21PsS4xQO5CfN
kFoR/2PBV+oPDGDnTMVsIUYnHjTaTOAHeG2v/APWR57TAzeK8tE+IGF0QVk7lOOP
92zfIl++bmj3zU9YGA76pH9VdhfPPdK87oDBq/QPFQIzGf1TTEVRsdfMgXURu0B2
KWSoqo+69LfrrT0IrTmFIfLLtjg+qD8JMTPKr/YJGH+jRVjmfFi1TDEFevqJJkT4
U57j1ILXlf0K/e2EU/d+k4t6p8Ss1dIPyeDs0dT3VxdB/VqMf7Z8sM0MM3qtwY1R
5vfC95fHERcKDvDUhkDMxxmo6au75wd5f2MZrmEB1VUkm5L0fQCfsyUUtXyT3qiX
S5GrjTqRKi9veRiqeR3auV9tJMmn1tSpCl6ndeNV4SXWthWVyYzCAd/azvvKHePt
wR8NXiRndR6fT8JKltwDyJ5g+jsAI7VhYXGPicbcdzANkKkxGMRG1NFr3MC9Tna5
ujix/KYx5h4kMezbE+C9ZaErbpsXMmpChSgR7jBJf8zir9qCFQEOa1bJ4I9GQ6vf
teZAk0Mm7T4rQRZk1h+NooW0+hGDqJTnC3cjnQFkc0RD24fKXEp2Zjuwuu5FI1oy
tCOFhtwCW5JjA0aKiVM70Sqh2ZgaMw/5HU96z1xOpFxK5cY/UmK2LHiymeO4Abkl
o+sZLEeaq66SQY/kDW2uU5fnKhjy3o1qoQ2EOpwpyvKDv49oVBg4anrRqsSfrSvX
BO5dfQkvVePsnAFlZOqcZhwC+3MI2UuyBZmjd6gI62X1SPm31WJzRKW5tCo4XqTP
fSaLgwuCwC3qq2aZJ3kDrTS/TQ2GV4sez0kuaOap3K31A0h1AA6zVsHG7YnbrnTa
xpgaaNC3H7UQC/P4W0ch1g==
`protect END_PROTECTED
