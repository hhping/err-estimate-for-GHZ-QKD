`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FVUHhIQIiYS63/RnE23+LB5QsveiPDWDb8Ju06s5uyb5sLD4TK9nppnRAItoKCp8
rptfHHprnQGg+CNKPeoMxNf6jz6rgMgxJ1YgoAkAKk3xXyc2kr2caT6PBK+edSnb
dEX/VNUvr9YSNb2GrZXKcyW2A/6tO3D/p69h3+TSmBUjuBtyqbt9RztIl6OEM/2p
lRYgy8HAjo2TLhfLy3P1kJM6CWCrokzGkL26VYOChSgoiiPoHod1faw1WznbDShM
GhVbE75myS9ik2bFkgB4g1vcDJEuHusGAz4JFtJ1SUhBzEtZb25qS2TV0ZieX6rT
wlix/Jp5Hj+zV9tc0NvZBkjvhqx+hWIiD3ZTbPaLXkWavz69j/X0BKflk6v1x81P
uwShhbXOqeMq4b+JxeMmXE0UNQZA00F7a3UPBJ/GCLFeFWM8CbZ3m0HyRdK+M3jq
+CpSoPLz1pakiBrotlF4E71um7RWFFqtWitwldqBbQhqWMWVWO0SISpiA4aDFtqF
2x2GorXlRc0H0Ukdcz0kaUYof1F5q7vosNp0XNHbuQZObpVjBZhtfR6WhUwWVXUT
LaMrW4UUqyIc0L8Rfci8MO136+C1I2JeQ/YQ+MiRvuRbQrSe56Lzt9W5mRDBVvOg
2LsoYRRp1apFD5cR6L+lV1LY8JUCrr8EiBFhhiw7fO563ghgQu4xp0b1J2/EB0iU
8m1RqoctaQKpNDuizTfCTa4sJ7LjqnlBfHsHZPQ8tG5nO0RAWC5OkRoHcFLOavQR
NGswB1iPT+pOA8DU6QlX2YvGRPBHOVk7vujaA4H/+m0yUmo76mf418GkwPzR76EF
sxwPleSyXITMH6po8NLq6O96AyzxNlyIIUCgwqLbDCC0wfxz4KjJb4lRbLBcVlf0
JmhVTe1Ukq8kK6JXcxaM1QM4uPsWtphkQPhtlUbfvmBP4Z5ktze4jYKJG1jBiJK5
Xn4QZ40yiq9iRDrHK9RZD2RVGJwK9U+7Nbbegji8yRisjB3ZtxvixvL4qOZ6fqRx
FM8UQTs/faFBVplgkJBnIeqGOp47cFdlSa2HEaJhaXMPyzaA1HWnWuid1oAld7J3
tuUFdag8zMy+PdPw6Lh3dgC8ozCzdsHtERQG9VGnORKKqtBU07GJ+hfWu+x18XB+
zwJ3uDxK5tmnTLeH3VmvQ9LNA6kdBmf+ZLalRyLQTcan/TIz3BwfbhnLNVfwPa5Q
Y6+9I0EMygLbJLVsENMvEiLfPUn8ytncsipVlMXfQSGO9P9fCwj8te0SJ+pgMhp9
7rwHwr+FAw34IHiw4lIJrIK0fp+0/QOVxO7xKRIJ+rQqbEpkkaKLizWioDdaBTdw
9a7M8yuMd1IB7X3MbkOKh3ZDBfEX76nRcrSVo6ml0Y9TWAabuvVIhbcs6vE4cTI1
DCZxil2Xy02PbJcsEd7Sg5OuNDwJVI7rPq+aGac+BIJZCX4k4Z44+idB6yhgZrYL
qCqH9ZbPDey1Ih8aszZijqqcmC4JNaFDaBZzpJP2n/m3nKQNEE8jDJ0xVQpwcM3B
b7r2PErhmuI2VZu2a3mASnha8YOK55V/FGkzci0JEam2NKR4a556uDaNarJdQZaT
nXYsvwkm/YIqusHL148RoPRH13CaZZyCLGQbBB1JCfVAe6MpY/iycRfhxY0+EzEl
Pty9S4KkEROVN+lsU4Miv1Qw43u7RROjfiUtDstwiuqW5twtxu3FGJXofv7m2kPC
yq58cMlFHu9d1QpA0Pt3WMQ/tjY8POOS3RlXVqbaZPW3KWs3QVnmBxX4VJ4Q8YZp
3wUQuVCeCjZuOtg8eb0JkVcoyc/qlKN58wsPtXzntAU=
`protect END_PROTECTED
