`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qQBTzuJyQ0eHSna+Hk4IFkqJquLK7N/tA7RoA2rTSOZy9dl+E8kQfrSXE+UIFhmd
EYXyTDc7kvYEMW3kZAPA0ChDGsbfdKtrZxArx3Nms3KXJONrg+p2n3esLf7vPXHu
sACeY/MLq6/zd9VRm6/fc/agw4O2D9hh+9OMf27weDzqxAbnRVpxf1miBG1armHv
jYwILkgRl9KrBXgvSSDxExjMCclyEN7dsCBmIq7T1Mz8RYnBMkQ1t5JsYfUWeywp
1L1h+X6f36DS2wTTWU3GAnKBVf6fzCeBFM4qboYP4+0bz0c1KM1k5In/xzYg/dlE
Bkwzpi7vGSGfvzzPUHU52AAGiZvWBEGdv32tsdZQOyPPSazHzHilG5hj/J34XfH3
p61a8t40w6KaFlNqYahhG3dWVyWg1HRac/79qfzkTtICtygxs02LrxCHcYAmHbdE
Vv28fV89Feg1sgBwupWeA2TPBkAKL6He2tyMVWEw6HVxw4KOaEeKI9HFvjmBFRCF
Mgs5VI5bxfCdUKhKgPxB3q81G+H1aCWeeWg0y6zBGz5BwDKcDa+qt6Ld3uaM+EON
yMrPVWv4R1VpEBTVCrH6VvSvAwuVONLqq98u8p0DdUrkU4LGknDZm5DY9dFvkkMR
Daw74Tyb86UEHwvVwGYl2WA658BtxfhMSGR4is3kxlAIx1/E7XgsOjcpB/wLwJhn
b96wzxyAAwTscGHadN21XjWKNgf42hfdHwXTCoqTA86hz2GUrCJm15KxLKyuCZLn
/awgOsy+KGFiBp3F772fglbmY4OcIK2b0suVyuLiyWbs2tyxaCJmytlkhpoidcSG
8FmqbQv22VLUHT34kAWmVjt4+nEQZ0G9+a5XXoTbdhWJ5zPVy0SX8XqEF/8ExDBH
F7y5ysyooBNh3VTZCesco6Zjw1NjvXTD/aS3E+a4H3fYn7OBaTq3p3mmJ4dVPKQt
2eUmoKUJknwLm8+MhiK9zuS0BPDT+VsR/C345zYXXrrAKAMh3zPtTr/c5fKRqSSa
rhFrHdIqUGFgjx8xnn4abb9BNnGToaQOkM6ne3wZyaSNQM0Qts1QvPjM8NS/Rjym
S9smmpvZQIsXgrpVIZ0y9cqOXu/FXcSuQGWwTj3Idj+tg6PuxHaaNQQgoXAvkHwj
ihxqdozGPIO0z59ywghpXTor3g/I3ldGHvqLKmRmjo/GCjR2e80S5wLoS6YEJX04
iq0Ddsy+dcV+M72xTOuqBbge61kleMmrpAnvvK/FMauW+4okFFkQUNseR/aebVvG
F0UdmlcI+BiTVb4+DkMK6AZeXidqWJjpNH/4nrRoLZ8XFDpYKAnhYa93Ushl0k36
qlyPnobV3LpQ8dqTozTeajqPqG+uc6xSK7g4C371XZs+S5wU5kPtuX/CT2mrRut3
878pSHStfUzIJ0EjsrLZ8Fqu8pKrVDmGAT8bH94klsjgM9GYQo6977g5vPbtl/Nb
P0iXShQYmriv3c7ogrCqV+notve5vzBukL4vzLJr+ctg7rC9tMTwCn0VqXfWdS59
FXmaFOEiEuZ9cE5i7tXyU+QFm/gM1iwF6K33NbIX6GUGYJJ3LA1hCp9M3oXv9XOt
zkJmhcmRGsdJ3y0gl9FKzznrd6YU4odfcuyzz3xtVIe7SX94ZMenocR9cDe4tJzo
+IamLrUjL24TYpYKFx76VN44g0eT6wEnQWz73P170oMiIMOnQQdJdMRs6AikXgiM
1V7PjyPI0H7JHFi2Zikqa+c4m7n7q6ctFgcb3hu3CWFwKmvf7NXsmVSfAWiZwZX5
DicZeZHLm7BJcREYKHP2PM0TUKoEIVfSBHhVP3mWMzOaAnDzT7ZFYHlQG3jK1nXP
orWbXp/fLVVURcA+rK0/m4Y7XN5IpM0uJpGIcyGEr5MtdhxGyTML07Oikrwts+tS
`protect END_PROTECTED
