`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
evYdyFE3Rx9sGQWBIRw/td8jy4GcSyGEIX5DODNKGaMCXHghzj99eyXl6pt7rRB1
rHq4MfmPykr1rbP4L3M/GsMydVrbPxU/5Xx+LgSgLFhhWW2ODgC/wuHPsNQWPsRH
DTgMQnbnGBzi/Y/LM2oRf4x1NjINhAiPy7CWVtVmH8NVzzaPJHD/NfIaUIsycgMl
iANxPcJtuD6pjZFtDOwfRjnXKB82rhoqvo0yhKbiloU1Oc0ZXcYQa5ZVwI0SYcX9
haipQaV2vnmmNYI3jcwiS2WGQVpmxT9I0K7G7t6hqci9iYSF6RUKdyrMXUKDGojz
Npe8bjJancg7P10YoCs+xT1k5BAM+EjMy0e8HsPh8EIhimZu+KtyuGiGYtJxMhDU
JluCAxrSAtpI/G+QzHPY0gDhBPxrBInm7+GOPTDdxmQ/WERRit0Kts+dkrqFVls+
m87TIoNQWtMVTLyWjuiWlLe/ohMgtnI/g7Shg5awjWeVxfTTYn8OHrJTOqaszYA5
oYPPmw4jirTmheIR6Z3aVzKMDCq5AkL//127ebWTj5lFexeiDxBQlPVpcNHuDpSC
`protect END_PROTECTED
