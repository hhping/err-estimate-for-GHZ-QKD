`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cqowqvNPbg9D3yqB4zePkz95BO/hK255bDa5baPhVfxOj1hSdU/QTSq7Wq3n0iuG
RS/zkhm+YHvMgHsd28dL/IBjpJl3vjXlYgH3FU17VXCDzRDhTvjFScfFZLNtZxBP
WiPfQIFkI0XEGa9x5iHldRaREDw2KzSOT9B/vy/YEdi5IHGQcrOCFMl48oCVkU1D
bfENya1SalyWxwGcXWfa9C6cP26D8bKQuP3Hgl+vgWV+6o6C6LgioudSvtwl68Jq
gM6ZqLTDTcBratuXRLqaKre9YybBEbk3FSPtvR0QXOmAFSaTLKenfJdAfxgJ9OgC
v4LPrNYErDgxyf4Nze+Xs8DJwt0Xiy6SD6U+LQ94j461il/24Gpmb0td/w/uiYlr
Xl/hkXP8Hhbcbqie3UQxGKLeZSqKLsSFw8oRFm1aczZpQtCJQ7ZxOZffsU03RPtT
kV+WszzcVD5/vEOA3icOXYTVjXmHfXMPC20/SD8j4ai3ATimGNzT+tEADtbFnMYr
mOetd2/RXAPAErKGGuOGQ/PPxlhn3csqfm6lPXxc96UFM+jd2IcKVGlPxwd8hOId
U9uy0a7d5G6obEEgsPXi6CiZ+tsdaVoc2VHXUV6YfpHNBOQ/noM/ZoMqQk25zIMA
LI19//ifrPVXpGnRcHHw5q93DUcfG5ZXy2QLOa+ETakfwcYfCsx4AK5EWHYRYbiu
SCuxThJyq+GHjo/T9QucdRJkb3x5Hi2ljK7TXv7ChCKGZdn4mWB1SM9ADFF4KQCE
uLHLCXTx9ZrB/QSbDcTFp7CFcwrYPaHRBRivfc084agYlKNGO90A+1MzAsaqOFY5
v33uywCJGBck27J48nllHMin4BT109E769PjWpsNBT51o0xLncErE+G/JnTwgHs1
rN2T5OExpSgUx3TBm598W2wdJtgUb8iBLLb+TZs/wljXJGt47H1Tb93brj/5jLrj
YHHOKwc2H2Mib6BoJ1qjBTBewxPkBEcp8ojhHtTQIJ8qhDynNH8Qngk59ql/BR9G
l8x/qS73WjBf3qXff1DssJbRhmOhjQYZWbijzosggJVktUqK/77wunjr3KDs96s+
NkkJhpXIP0l6GRcpyV/ZRO0Qcm+Z+ZWw7boeY3G7c0P3FxKXsP8GCJ1a3ym+nWTt
12OrazMjP0HOxhvEFubQq+X10F8VeWvJCCE/kYRHjoDiV3T1WTIhqe8LpJYjjL5A
UYS5dQV5p5AvQ4UOTkdMWT4Nrnij6mAG+w+hYmWQCXrv4d54k2G+FuEeYT9FsjwM
PjLQcxpA1zWlWrNwH54m62K8WP01Hg2H6rd9ajexsyDdHBSysZT6BMWP27YRYJc1
/PhLI5wE5UHUdiuCzsmwv137CKW1QoQfMGMGY/fhAJbLxA6i5W0sx6QZmjJ3JkgJ
tj9bybIhxzfBTav14AX07HbJpZ9d8oZhiAxH6Ocx97/ss6KTWq5CYXrwKTvRg3BL
Z8bvtIYtUpdEzncuKXH6Q6FlaKOSBDvSM9tAfuskct5TgUUBsnWsiSfUYjioG82W
z9GdpmYt/CXLzgQkFSWQalg0kdjmD4FYI1z5iA+NAa9ou7BECOTGFMJsvGYepd0e
0CpCRavGyahlVLqjYE4ewuxjYvclEfUx+BOVGawb8lzNC+AkgD5vfdLN6oCh8qe2
WBtLz+yIbR8nB1ZR9H/aCHoahQZoKYbzv/gy66kCwslqM92Zdu/zkPJcuprfLmCs
l+24sbPKF5Fjhm+7GJvXe0cD4HNGrIvSAodu9LXMltZfK1D1mtlQ6OEV7aYLsqKE
hnG+L6uJd40GfsLy3qwMOxafXllJEum8JnWpwCK8185xUO0ELrUM3B2vioIbD08n
NJKTFaIpOIuDd6fB7h9giv3QxVBsdCtFK47k7YUZmwckvAMPoZxKYHhuoKuw2kGx
tDZuLafFC7K5MTMXRAJoDo2btufZ/VglsJcDT6zxOyJxKM7TDpmEgxX8e3WSXPz/
c8lVj9OmQe9JSpqpqbTIJhsbODLO7/tBk5/Vu+kx/Rh2U8S46bDyNXUOfbRDF0EO
WV+HXvVMeB165wUZ81BC5G+IDzJrA8nRk2GfxqQgtGWHRwj3NvybO03tD4IkPMdS
QLSiwHG85A7UrHz++O6aC7mfz4Io1sCdMVn4ZJ/7uZXMj9gxXhaIxUTBxopLqwEy
nqphiVPO/WLZ3yD56ji97qJm8vBKM5nx/pMM4p9c/EU7icbGDT9P3YAXagqpqiMQ
5a15ssNhVmEzrTFsuRhBV6hFHBdCrO9mbHxa8SivJ9Fw2FbYR19gahj2GnLMduOp
mdmbtOVck9iy8tshOOw2l2RGfE9Q2ZyVtAiOL/LblKyWfvR5MVfjVAQ8He9YKE7U
cfWUWCQvgUmY9bSm146boMcWaaoSQNsYYldd35/d9R2r9GI0CxkAmshVmroQG4TC
HX+QYTM+JggppSPfnJQEvIZVB3UxLrgQDZ0s1qXPYcBBTRNBBXN+dNn7gqkp+ALG
+jFC/JkvX8sPlerSZQLUw/hpg8fzMaTmZuQgfkHhd+nkOGivv/84GdjObXnSLSBz
hPjGmf6yl8GyqXVOPr0bcN5izzKIBEr900beHiyF92L/SKPwgNyONrto4qVjSzA5
ys1QV3gd8b/8D3c++g1j7Ei3DDCygd1Imsj+i7NBt0xy+z9SKcmNMgjRR2iz2QHQ
FX7MdNfU54MeZPaY24oBQjDFkWe5SrAX3rMjXwWuwj71pe5eU8D8lpuXQaS1m0jC
M3reWrOIV7t8nq2yugCg2Q687v2yCnfi1SAwLF8msuDkvw3IkeU9CXKv2AoJxWls
+tkzMn8T9R8Owa0C0vNa4YjSMcA53szy0Zve24fZWfCc2yQFk8SWhoiRXlMxZ3dD
bDWeo+eOe/NTtUreLCZNofTKTf1p/Qn2UVdERiCe2Gnqhc2FoWZzDVC+l0OlNi6C
/VwdchLHmfXlg/GuytLofNr4sMPicX0awoszm27OIq5tcg2sRCBm2tlBfVMXUVxH
AL1ponBsuLigKMbyAyIj6bBBnKrPQIx3GSjRUM44z30uHAYvqXMNDpMBPAEUsXgg
65M7SOCzAkO9ojJyrn1AErdsz7sPrGJn+1hR+jyE9e22hUZQ7nNJDUrRbiJc1Ket
V1VSB75O9K2xQ0xD66pvGRVrjK78fK0CkMTcDbcaMkTDEH5Aay52R02dcng4bqWP
kDVMYzeppZkgl7dwzYEu//IrsurI6AJ0MiI/nfetDQkbvczkqI/Q5gUlWFXde9kG
L1Z2fIgX6oK5gIhIy75p5tNkCHW8uHSoLV39eRTogycTFH1WYF0BfFVQ05V9eDyV
d3D/33qkcIxVFG7qcYrXFl8nUWuW5HfpTnENZSuIUmq+wdnX0EzZYYRqvpg+rJ+e
aahCu0Q+Tf+WgqEDGcuOiErOI+GcyJlpUgqZ0gL2+TAeZAGhG4NtcNp/mO3VOyda
nvP6hjHhvvie8Kup8MDnz6mnpO/1mJ+A7BzFS3T13jphMw6VyEzQ9zVTF8E2cuZ4
XKyTHV0fTcduSY786Fsbkk6p6yrzQDm/YRXByQHp/AtGif8L4dksv6EEHyEyBCrf
a8a3UDRzlCBC41xsmUaHBp1+6sXrtD7jOvrHGESa4H8NlIBFWbd5duXGiYZ8tQ0S
n2Pl6CvLvQGg0h7BFeZsOr1GukryEcKMwv0oXQaPjFJpnR/ExEdHSQIyleFN5I2E
J8Noc6vtyKul2bFvZkAbYpde7kFzlRmSxYV5K7QB8hMvWTG0+SK9qLlKEEL8g1qZ
OaecNfEfoSoTF15yCPtNyANcarf0aw3/HtVc3/muxGK/XqrsP9aH2NbHzIYWU3Gd
IB0xzZDh6SSbZVEV/gilnabSte5OoMishMM8sMyClZSyB3aDSQyTBW1eb/Ann9v8
cbso/Dyv55qrE8HnXiutdfV878oGRjR99DSVKKkGQk3w0JpKujF71aex8rfwARyC
IGAHBgwi3kyRN8j+x55zbGzFd7Jb4DPR3oaFqU23zHYSlCMr0Y5K5YC/fyGV1LjW
ADbocGBIYNcdDJMB2c139CyuqSYJGn9xhjkxgiNWLTRBx6UFe3xU+27nZc20GBI+
zN/ueTDE9T2FJPy75VzKMsmI3EQ/OELmrUyHHI7MQqV5rH3mpp3DYHgSgHlE7peR
Wr+XCTmYr+3qofFcwXDwxNLC1zcfMOC/HyoOW3zMiDeGmNuwk6gWbB9IxpTgZQam
gU9dkRfD4QOJTAcz81LonBHtdSVIpc+bObtYULwJQHNSmTlh0ireiqkMM//oHkoT
Xy3/vD97eYbnWVU3CL/YnCKvzircJWtdvuQ0h4nmzsu5zwW8ySH0wCpyMi4zMDFk
FwUQ6qXQzl7tW+YoBWfjr7gt2v6cKk8DgqnXZznZ8TDmryT+1e8FqLLy5gqq1OWl
TouZoLACuHZ/ViSHcrDoG37y0Lq9fjXHOEJ4T7l9niaKLk4A+fAeHyGaFqIuqHjj
qvN4XYCmohMGBEiIbrMKoF8OGD/KMKFhMzydycf9dPe1Y6YIcoGrFtZMWD27ASr9
Bx7rIY1+VGOFh0Sge9z0s8BnKTumSELkAh8+tiSzjVBh9It/oG1mQrPFYbI4BjRv
R6bu2b8csfg457yEVXSHxN44PJF8BMAnHfPn4ri3FDqdfxtK9qS20TN8fWZT7/6U
ZUYyENUn3pbniwCNMqBqmobOlwmc2A9XFBPr1fPDb8aYagCCSPtm4d+ON6nvHib6
SIegM2Ud3GHz29RHUjX6Aof2SzYTlNVwt8juQmzm0PIipnLd9+62B/+fdHoOSX8X
W4Zgdw3X1wJCGFCcd8QYWUDW25FGU3cERrjXKAq+me1ZxsH0VEZg5Az4+qh2E8WV
+hef8GTLyY/noTIu0iTv3XzwHMu+vsG7XLRtU37/otM501sKGzf078TkslPaqPIH
FkMwjAwNxWnivlSY5ebMWQobxmB+unDPY1zHdSLDF95ptScrhGxvNyUxLOkfrvRn
lC6nVyoJtz4c+82bm3tl+J1tEu5Q07OWIvBLET/NWR0AwI87NHoO1FG53NTlO0gc
CY4WUOzAIOoNFcS+JFMWL0C1B+c7AJg0mu8RJsHy7TmgTIEo6fg15HjmSSaiicTG
vkhApRt0lAWDJX0WcoGA6bW3iusmiKsFq/AQJlSYRVBDLRskW7gHgggFCqCEBN0O
ycUK2V/WDp5lGXNXfhiyEit5fDOApkt6oSXhljRiwPk1XCHma6xXXjqhZPCqwEh3
WDIxtJX/u4pug0yiRRi8DByt3FAdjEw283i5XyMqlb4sLn0BW1JksqctunoMJGzc
u8t3t2MEYmdHUpb9haNwNVqvBrQ4PXM8V1HD5AxXXLgBIIbDnKIS3PJUTyHUwZJe
7dc2JsQbTq6dzvrQtcBl1gLIycOcDMHbSzZXVIdRAzg8cFGrosLOZ3Ckp+mBfZRx
LthxF65UyYHrLBqQIdjQRrEoRnjnn4Rl0YXRw9ToYbmqjQuLVox69Dg0QOd3ED53
ysIPEqOM2KikpvJpSAiCGipsrbNupTE7vO7RaoaVpmAhzEgXKtPQCF8Q6Iaa+PnQ
WCQScD4CCMr5eJKk6itR0qXP4YKqRXcJ5kABfZnMRm1mGjgy2kN03MQPEYKomudz
IUrKCCa1f2lL7suTo4j8NRh3mfxpFM6gP7G2NA1ZMOJjG4lHJl4l+kIOxo/NdGYl
16vqBuQDuc4xAcLL+vLoUlaN7VNgVCnY3M724qzmrWUSlsySd9OqBOYRJvVzvNNV
3W0nGAGaCbGGBXyxpfHT6w76ygi1aBXbMK4U48frmPnAjHaxdl/6+pnmheuEI0jH
xzfnt0+1fIyGmiZJUL3A/lVNXhDlA623tBcs7KeuSOgLeJPrdFKwzo9D34pH7/Cc
uU78msH+LeIIgTzBezEoDXu3SkBKAl/gt9cO9HE+Ek01ipgFf829tnxSpRhgG25o
++TwB0Kr4dg4VEvxDTDJiwHWBjgYg5fxjIAa98lyiMiPdP1zADOii+hCFe4z5F1X
+QGEj5FDHTTbLzlEyWjLj55xDjsets4cKV4OPM7kbnkkou5fHd4KuFe2BqTKRIYO
pHuw001XIZM5pUm6pYxr7EiNNtyQWeqSK6SvlAabvbfP2wIlCpARG2T7cxr0O6p+
7a5PsRtseXAJqwFHURbn+tbJ3uqGjZV8kWGxfNTLg5t3VmfrspkfRPKkKC3lgWbb
TgQkkiU0eTzmv3YD47NmvM28X+myOPFpVK07Zh7AllU8hR6TdSO7dYL8ef644pin
o4YvTlsHfr48YWL4j3qAxzKvaXVx+Go+clDJRc/grJQb5DHvKjynI9qV5McFvI+q
8ctTWdcUyoOmXxG5vzT4jYvPLEhVF+Tig2fnX9rmvW83J/lJk8vmWhYp1KCWWtfk
lO+gsBKGOPETvHG2igCRWdi3DJgdMxiKwU9pRcjEuEwD/KAmNTSUDMQ47BfoKJp2
0ANXymy8OHU3yhx+XqdWVpoJmI/GXTKIb6InJOpvaMFXo3qC83daHWhLPAypt13c
mPB0kLo5T6wkUL/oxfcHX1f0PrbAGilCPKavheudiIsquA+n0EHctXlaYch1VS5L
c4nBdb9SgW2pSfa+FdoFKGVWfvwdjvAM/o8WGdMbjYRrGmY6Huw2k88Oe6O582bo
YYqpkWExYFW9oESPBobN6yTbq8VE0mchW6iO6YFcjUOCWyzSvoBJ/aWPsauK7f0s
VNlWNYUNTLuFQCx9KZBNfXPyL2DqG7zBm/ErYwrY3cq8GX96836ShwDaKqqOVhUz
/Q2CKSGCEHJIsM2JPsfsWM/jXU2142p8vSOEFKW/lysDCXXCpk9nRUFa4p0rKjNw
PuVdQYmLRROSUgB0NXWjwf3IckrHJh4tL5erUXSCsVhVD8Q349PcJr+8FcFVND+g
cmsjCCE8Vcd42ykxUv5JjF3cK4kgpb74gcy0dzcnu4g8gHllj3t9s0wEzHoXRMda
NHGLtTApkcb6IBNsOGhvfl4cAbaej27dwOTRbx6odPiu020fAwDSeSgg0CGBWkyT
Kv5nt0R9oVV4RuCoCSM2silCJ4DF0U19Hzf+QImHt2rDRQzfWTH/MNnkh87N+YiL
WR9s8MMx6JBYs8IQsRip2wn8j+eAWbjIWknT8qALcb1TCCOZ3k7YFZopyU5ZklyG
7Ddc6PxFdxE+34tlJzxv8QhN9oyq9hHR/MIMN/42FE2WWOjCVL3bTOReNvEVWvhE
sEV7kErUH1obevB5N1RnKocMcLGzvnL+2z7YB6YOxFPj/I6VVJjZYnzF3QcUKOIi
g4OIGP+Xn4286YWx5aIx0KO5IXYmIpx1V9u3TCGOQDyQdjye23sgAU/L+fJoJ6sa
LxTdSKU9DfmEmCOIdQIFrlupn8vdYy3DzS2m1aBw2AwQk2+trERJ5Nzu7BSW/e8y
hYOljuEm3BQ6Sr/Ql3TsBiXz1VLJmSkjtn6WaTMradvjNdKR9FHi3ewhoJyIDsAH
jklq0qn5egEq/gJlmvAB5aBE5QIcrfH/kVvChDhmpJU8dpIYaAgYjyEegjtxfnyx
th08Rcuqy+8YHUo1r137ADdbxOSjdzpJ1QFClNlV1dRy6Gca8FPZLkECC4XRCeDY
J2y4YAhpDzvoJyDui5xo5gzZbFChLbGuRUVj5AtfYxBfK751kt8506pjVPWWkImN
xirjL3Trude0PwPDiaOq0LqvWYK8+BgBr/jtSfX8IR7Bm8gISHxK2Xl30qkJtoGO
XhK+1O/zppkRWmkWMo/RDqs5VTBKAvl7eF8uyxd9RyQWCDCd4hI5hisJRFiyiCuH
SKshj9QAtfqCrKy+NfdTjUCw4PpN/KCMPe94LFEEpM3rZIqsc3cS6GbCIoBTXdwJ
vee0pKhzDkysC5JMO0VtrzFljz4BL4pctBFd9lcnqgfmMzhnbBbaNPSXls3UKNSn
/ZG1ciLIpR/D+8UF04qkaSaITpk048/QqyvoyHJFPDi5f0mBqgpcLWMVBQPAo+31
qJLpnAFu6K5GIs3a2D/1NoSnmcLNxkAe17sbwshw7rJE9wwV436L5GJn9wAZH8Yl
S4NjOnMOTswI6ux7FrHnvtcWZ29Fjmr6MhALpMDCwR6ka0iQWiwwDopVGBKX3nXG
Pb0Ph+ETZofYUzZm16k0QKPNy+7LRr1hrX5ikzdEU9FzM4LIgtdbmY0cu9cuS8lc
RfMu+dMGoMlfmKaDV0kaYvNBkSE/d1idC0y+/oDd0qwzF7cZleQ9pXs7dhe7RaOB
RgOiudSQi+7nTTU1IVwefj/w3+5to84meyeuzfJE3VzfBGXLTi6mIjTC4NerQgMe
v1ZU9rJ0gTBCY98T5L1HCx3o1jvgdRie88e72pKZ5GZVTzQQkhylJa4O+oS79Vmu
rftciG6QAvrhrq1zZOPLTwVDpOQVhBQTWVC6tRIgNMdB5TFIowAcSBcU33disjHf
RYKnSsNLGUBoZGuyXdWMfH2IrX+SUOk8oURDKH15D8m04VX+D54ES9uXfd4SoGzz
BwUVEiHyBszqJcDlwTjpCM1Vz7xVWMTluTG4Em9xlU/A7J/QYKTRvwdIg7uafrrq
hEpE4kXOO7nVpbyZUzzYkTltO8EOQo6/sOEcsS4kwOV9lz0zFZeLyERTitJa4/4R
Vftt5dKXgZ+Di1W8sVy6BHAsTZnUGrZUHsU3bjy9Rjy534kwbv7Wo3wY++o+CVJg
Rx3/00cZoFrvaV1aSrb3BFL4Rm9urWCuedKI2OHQFwz10mqBDiDZmMgqiYEFxGla
Mr7eSLoCFpcHjdFCowMF6vQEM/pszPlh/lXkLx78pNajgzdUsyzf8QHnLDHLMulv
WJmEPHGHlRqHlKV55RQwn1APvlzY+RebYAA9dDZx8DEJfLwpjutnc+MKcmyFXpPn
CD9vFLglHWDtG/Un8zPgrvi3EPEE/cQO+ytqH+URlQz+fIr/BDwdYsq2UlYIa3lO
fWm3gGHHjDwE8HjAgEbhdk9OpBTVxu3VktGfuOPmx3905rD0ze9wuMp5hyaU3lAr
scezNg6uQ1bZzi22eEhc+HNqsGlT33DsnVV0FK2LC7VF4gyQIkhBT8Gn0L6t/ODV
kUlZemOHKzq7mBE9zCBtsme+EfwwhAixeOdkJCj9FMjM1BMM/+R9gOlznlRWFARN
NPbVZEjmAP7MKcug9S5msYZrnyvZJ2teyalxBAMxp3GzvLqlLwUNQ6VCqo59uvB5
3DfGALBCr03WNPkcBwyYpFL/X73jQfKDdjuzxzljmEW7qumyz54786SdZJysVl/h
JfaE3+bkiisJr7rmk0iXPGQOKh2r8WheChgUpif6QOpjlg/9Lj1aKOn1Tltietjo
BhzppZB6zTxohjzeOZVL/TU21ff7hG/P5bw0LK5efw8HIkngHeZ4qU19rBZBxmAA
SAYryx71rGNCdhEqAlAPiv5M+psOxJGm97hzPg4R09uOGRzUeRxUJK852Up8AsAB
t13pbas7DXPE4sE++nzpxsk1R4sTuRoGCfqpTyTsNz0SuHKKASRvjjvlEe9qRsCa
V27LZIC+scQARMLlzHZA/Ww9FD1W/Y7EZmu7kHRCb5LO7h+usgIclDrKmhz3Egr7
y0oz9n+PWlFLm1m8bsaxr1GEf5ckU5WJUqkNxUhBPW9n+w3lI9AQdyruwJfjytxg
TdFvSEEIL1ZjhAG3kWHZLCvFVs4CO+oR1SP82rRwIQqUsw7v3vK8SHx5XwzSirWE
XSNzanQT1y+mlbpnSBZDwY1RFT62m46bfZyaJ/DqEYl3ZQEKnS/FGcQekjD49hjM
G1X5sOtuRiDgugiHRnoUjIk5T1FIGNV2m1bUmsIaWnK9IuXFcdd5i9b2mBL8b9H6
2KtHOfYBBcSkhKxusazyXkfDLWp0VVnwQNpgxzGIbIa9vtzioq662j4PA808OVu2
slIOkjwrTj53cRbPHb/msT3lHXkZLOitc74K+hdc4H5iINOn1mJJz7WdApuOid8h
3cn0RzePl1T1WPaTSYqG/el9wDKF0Jbuj85zfMA+u5fwcKns1Tz9uZIdLE+wuDPQ
YswFZm2qNUjPNyiDaFcE5CdzQ18wP+w43jyr1IUn7V1CAPgN/3WeFGWgra2rOT2y
QScgv0vRj1Teh94ANQVRvAS18JqczjhGjYgv/Ugcdiv8DFoab+kXbYccJRrkm9/7
guyvDdJBmVe4qQ0J0kwFEHIag0NF53AnRReGKYIPT4yLwpeZtBf+EuDuOdifGIRB
K9SVhGfcX45xjy35NOycRSXH2EjNE4lmi06ajbHXZJJasI16Gsi2c0k6KOM2QwmX
RSYU6blyv8+lbf/pg+yItAYPUbXTJfgj9Tap6tMLtANhdiqNqnccG9Iqxj3sPxcW
sPVYb2s6o6+wRWQqWaI4pkmzZhZorWyr/Xg9dCzsZ/js0VQTWapuK85QH3Y1qn6a
Dk+FcaWZWs0jt9UgHUdjUfDgr81DwjrQw4Xj7EINHXqktfvWsrqX5esbt5R6uGmX
54wTQura+yztbquBbWs0fUO1m8Gf2DfYVBkxRIYEc30fQu78y5oOJN1lwNLLn3Iu
2yPBpl4en7bxS7oCh7ob2VqBCJOcSTLrQUmRd4Rv8SfMw1028xZCa3pmGRNrnacC
bTkHVA767/9ifJI2Wng/ERPmj2oEZu5c7Wc0j74S98C7V6Sb4NR8rB8UZn3CodXT
cNix1rkmK7hwBHBzaq2ryMJae/D1QumozfyaiFw1l70uFh6uNv6HxiGZfK9trDfZ
CL1DaXSei6NeRi/bbXWgRZmr6DUhCXF3M1+ozCH6SB2VcF0IgBOiYtyCkrCFTM7O
kjh5zfw0BYvWUUa5DVTM63c3Uca8DBaVYBa728gQrRQOje4zfV8DHxP7zVHs1evy
FyD/KERKLrsJwg5E6cEfVEret2AZQrvqJeCx1KhCsNKPLTfK9zXOPI+9gWx68+DQ
tfh2MQeCRYdpp4YvIXYMtYpFrWEQDT1MtYuBDDwiWWivzphBKyZ0dCPBbQdNFdu5
rfbocFIRH3RrzrC9Kji5KtVniWKnNPwiQ62cwW0LFjYaFG+4iCMPzhzqAOWlVWIj
fHj1EnXXWL/xF4/FB4d++aPaZZMvSZ9yiyjRxGCv+GElIjiitMonLgA89SeTgi4T
NZIERZQsxf2eqozaZRJFa4RnEo0CufZYBq9CunUutKOzIbcMbZzyzfnnS7Bs0I0z
SsHIN1Ag3ZI1BppO/aa++15/GBvnGJgjnnLSfG2VfuaQZ5Kr5h3BzA3ZUTxxT5kN
sKori/4AxPVAHSe6WXUGO7QqWGIBV/nuVOM39ZQAJ5LpAI2wGnoA3JcCikUkMGsd
hvQdZpx8Bm5RuJnpzJ+0ibMsuPGT8SaLUZpNmwsynp2pDKCoct39DURj1ijCT4ll
xzKnxLpBUwjADLKMy2xleRqsuSCeubUmR1dkIzEQQS9tDIvvHhXYieJhFmkHENuA
K8xsYGVXlIZRk6waWuRLyTDyH7UIxgEAHCt127gDR7bOa/bEg/8j7y5iFwWKsqp6
ZJQ0SvStxk3vrzde/mb+KGE9tIE0z+TKX/ZHLsFhXQt4qA7k3HEIdPHMU1Jc/mDi
RKDhnzPNmTKifO1F3fIN0Azt9ScwfLH9GO5Ts3EB6sw6LX5p99hjXSYWpiwwjjTM
sxH+TO5hNUsUDflXWUvBeddqS4QLZWS5kwYE4ZiRVdKStNOSPYbusvuvwJowhgwS
wtKrePL6gjNeSUFyEiMKz2o9o1Fu6WcOkceSeaviCG3/iTlhpqnj4jTZwp3XqrSD
BnDJQFuCb6quXfzJqF3H1yf0zqaKynvQfPGeDMg5Ig0b8eYpNkkHcQIEeGG24X1U
oN+7RnPjxz+QbfeCXT68GcklF/GuxpplV0WWtEZkSi7wgC8Y+WoLevYfbRYstRQr
k6Yr7ozBzh+o0uYW9UIkFsGuNUe856GFzdJ9S/W5xeIBLdNimJpQ3x841ygFemo9
K8w9r7mp23HWOo3VAcD1K18f50yJAdVJEuyhmAtBOWt9TDEylpQ4vw9bFkZfibro
26v+berQ1tCm+agKFEJ1Z9PmRDEzHEWFy41/1wRsdPvBu+x8fvUClQfDec69zy3p
/5wxjPIomY8w4ae8TDC97HVptSlH5yWhQIEcxPKtR2+fk0sgh7RJYKdBd6VBfu10
WDDggcA0GQiAph7j7R9YY173AA5WGJjs8IlnbrCaTOQaXEYwl2Q5VKqQWFnFQ8Hb
T5MZezLbgPTjT1LQ2UfN+f4FF+4VpmDt+PJItRCcxfLBrFdRT+AIiTPZWhWiY5nL
aI5mRs+NRavyogyS2WUk/CmxcguAPFiTfqjf7jeXmySWESXoeGiMNxZtXqIuhSev
YamuPvqMuRFwId5AJI1HXsQNOlV60696wn4K51etQLhoasD3r6auRVO6/kEEXVU/
eq9pfXmywzZajJL88+fJ+DBlFlfjrU+wSSSTYPcyuzijbYjRX7XBnMrprk1DjGdO
YcYxRhZ2+UJKHumGtsn/OXCJgZcYngxXmLjKGCtiVNXpj8TA+QJDTRtngerGC6ZN
7DVXD5/by45ytLBA2Lzzz4qq0Z/eT5EkxmXEpqUx7IgG/uh1VX5Jj4MUnunaEcVw
G1VzouUinoEl3sF+EdSVe00i0luuZuKLMK63DJ3SLTGVb/Vz5429XRicZavJwpxX
DohLGqTFGdKNcGhPOa8HxYw22XweWXazxeynZXftQgKZgQntJY6jvW/l0iGMjyj8
b5B1nDK+IftkVadVomqXyHV0qSSHbNkF9yEbfIEEy0vAyO2snkEv1+GFcGzjpZ3l
i9txFq596oK4wuIhXuehjce0OSgk8VVbRf8NQA40AEGo7hLthWA7hIu/zxTwFk+c
DyAyQ8/etCq9EWOSsM4mx1NuZySSuQ6tTLgYqVv0JlNY9rFAw6eN6y1FtWHV7Ba6
siFlx1Ck63IMledmK/ZFUxUg/rdbrKPXQusFfoqhBW3lk5mbvxXSJBETXFHt3sAk
pfhN9u/zr68iPIOhWMrvKJ1Sxi0SpJhjuliH74bAoe8FYtKVvlb7x2bkcdM5mo2A
jUW+MnEcHMHcivjsqlYD6IOG5/RoahduSHs35TaCe5wstt6lBIJxxhxwUp6Gj5Xb
kaeUpHrlupyjaIl7on9+wofqvWQ3nsC41uPcwY8wSnjz9nEa+5BOt1Ammvyz0r9g
UYuqN/2QRtmUzy/FgJgt8dpgFojsfLuy3oLKG4XgiemxTz4nirX0LGy8EABkWUgj
TvJFJ0WqlD5DWkY6G1FlB3c1dr06YSZmM1bJkuskts6B/gUlyZYyVjejR2AuTJl6
LvIg7DDcsG1zplJJ+qkVp4bwTTIjSl1n2FWl1lUHO5wuGRkuYg5A1pqFS3Xs6t2y
AKcjf+gu8cicCuQ7RVQsPhcl7/DwDXrz7AZ7X8OhN5ePqXL19OVIc89UUdOilmQF
ysFKvHSvmnlSAOsdEzPWewWsolqFaU/91Qk37YYxSWukMQgWqluzonuPc5ekYMkf
EqmMbOQVk7uzJfP13yMCtVcXHAnVupyX10LbHva28+nW5h1a0tVue1tLxxUft67z
DOIAlnKs7YGFUxQS3T9vHegVmEyuPySqpWcO+w9RcnBbWMmVR6QwLIz0J9ba+qHe
HdtZ/uXi4dJheaDRv0ShEYPH2Xja5s9Fw64sisFRxxbh9POe/BwRiZ1/j9a68YNK
Au37rhAKGFqE26bNOA3YhK82GpiYIcT5aLEN40QrH7eoSgqTvp6bPyCqpObWbifb
7HWZIpqDeQaoEfwKiVLEy+NGba79Xlwg3VsH30KmjLgeozGFs3gdnY0d4POSwoBD
9F1+9WwTqTFFYcmEVinFeUisGiC6iNoALxk1YtEOc4LAyACNjq15c6Tl8k0tdgOV
uJXbBtYuCQU7shFzAWxs28BYW5zPfACuow1nLQkbAPOg8zMZCRqiej7Kxt0iwCXZ
KGjTFGjpR0+nzFJr+iLgA4JLP//Pbz5XEgCFmKp5rCb4cB8FZkCKPfvP5Vgrj/ro
kyzN856AJoMG7dF90MddZlbmi18ivo42MdxN8FxmxEs1qzVkuxspA/ryMNCt/tg3
D0usE4r1SbREqyaefatblbBafKvtcYr7x/XGLY3Lcp4ICfow4kzpVP1Sv1v47fE+
lOqR7H6+C4tDqSHtRZLrPJl49MuNaHP+L0xE3UeHUy5cki5YUzGXO+bVGdk8m5x+
e/T/sxSDBco+dugrEBI2QfGVoA+RJNKFk0TItTQ1TfYc57t18lEbixRvhzRN2gl+
nand0xZLzdipQg6ovyZjjSmhhLMFKUbm0kbipC4KpCk8BEFYNlr2B8MZsWkGJAR2
/7bFZHMLGILN0fP9WRPfVU0eJj4SFg0VZA+HU6M3hNXH5eGleDW62Vqko0mRhOfi
QMVdg3njPW8tUpvTiDh/hC+yMNlp1+HEYJr93ZLNHc3B5lbhq3P9p3ggHfdcLiTr
KeiFqr6ElLSsiRExGeXAYFaxj+DcLUxSn7bElui/UbMw+1tUAAvuDCfguEpshpHe
3o7PaaFtKQN5jbavyfpg5D9DTi9asLIZheh2DKfA03wj9eklMTlgdq/BfUymAmGt
ZshWzSRXZIfyb+Tg10oD/2wbE0CxQ631i3Ti5KfWrY1oHWmwW49WWSXsEJUORvqN
zUiBS1x9y8H6QZI+Mhhjx3FtNvVQmcFMy6nMSeh/0of35JccnAoEIuCO8kR6nnX+
E7AwBJ9TmskiU3LtCf4MxcQYAkg10gwjKdS2QDhu0Wed7c5Hlqp5lilzRJwM88Ug
y74wexAs5gwIO+UTE1azmE8dQcYkwzPqWeLCfopoks5mT6CkQA8r/YbOagse7rCf
sDSHPIELKlr7WUB6I+cQ+46Cob/1V0beuhDcQcbNzY6sET1iQV+b0iwHtQ6najiE
dLDr57F4jEmjy3OgHB7gxre5v4c8O1UlKqV+tpXXQyF1dg3PepqaXk/LwKk5r7/a
J9i0wv9ghcyJvmxVacBLzcj+FzBGbhKzqYsJFeeosUePSPJrJ85RBPdsXvia5ZDZ
I4hRHBEpXFNMq8lIC+zcZNAworFKeU948jXuU7co5EGnENnV4dkAN/R0KorpdHEd
ou4EoDRLDnF4FSBr8M9IZzpGEkXxuPdRZkCrJ4yOOy97eIEK940DwGvQtDKPlA5A
jwbkVM6/ZvjmAQ7TsNfKyTPNdJb3Fwhc82zgwkVU8f/82dF8eS3taIFS7yGBStEU
0pTZEzHgP1wuEaCTGyfk1xcHTMdz++vGIav4qOGQpX/eIy8hY5aENyUZefEt6PG1
G/85BatqqSj2KspbCIKhOk1sSI9d4pQmI4Hu0knxI1rckfO7cyinoapQC4xIwV7e
Xl8JvKGkKKW6/VGULpy205UScLMULu1Ou5LpYFMVEi9DsztqqhMnTElrH4XBWIFC
duKCbcMdkxrUurVRIwcWN1q7W+Ti8a17vaqBQqrStsnM1pJTY2onIpVo14i3ql4X
2os+uZK0rEpe1GJzAZCjnUM4dTvlfzl0Nii3c3L9+z4C3SGhMZAbII7uaCwqzHTO
uIC3XDvCMaKR2aOS69KwH/2ma/wfC9lqUzeZ8PDHdnfRWRqA7bvi4QhxV8PCU7cD
pPehfQONa68a+k1Rcg2F+Dho+lCtdGCcAvXj96wtLKfh/ZObkJxK0lmfpFVdDBqN
9WN8P/B09eEcVRXiYOmB0i5rgZEWKfV3+Bi2bfFsO46BASJkmytc3fXsudzkti0+
4Erp6N5ekfUZkBBUZISpondbHQk0PYVE2dybdjs8EuV1lLvsFbCcTasczQB1eZrF
ieC81nNIRDMDLG1Wy/kpFv2BbRDxd6nPQf/b2SeAQYY/dJZNgoNYCrxbu9Xw8Ieg
2iPFxQgi9/s9Ter53Zwdq1jh3S/yIg2fTOlyGtbp7Hx3K53uyeTYXDIqPeOF5N6A
C3EfvrBaBLX/5hiFxBitu6jw7tn5enhmDoGJ1XQxBI0XCKpd5/c/qt03KlNXyQ0h
oVcPHPMSeHn9TmRlnO85NeoSzto+pHiyxAwuszbvaEz0XSyKxN5MAszgHekHOIjZ
JlmGmRlHhJZQoGNVMLkPEYdb+eYpCjb3qjfVEATH/AGC4WpvM5itWrsz8cvxAK/Y
gUG/Flw8+71cABGYMhBrrjjEdrE867L+djaI3xJIh4zKCzgsnXJt5KvIvJ+aEW4G
225B56MRbSrdesC1CeqgeGYgQ7fK4bC7ZxdpUFVVoJq9QsYQlmhoMJgdPgK0WLtX
9PYUJOVMNCPBoG9IsG0kFQoqnM3B522eEsIBdzpjDriwJAxqt1S+wz2xj+4Fc0ng
PmkV8NRtllOgdLqIt98zmi4JDaO0C7TaoCUMZhSobc0JUsvM1LtezOMhk8S6hL+V
WsbCX4x2D0FRfix7PpQTiIuz+VWZBsuf4S36FUt6jNr5yZGXlLXnKpSKWe23WFJg
j07hph/2ljdKWd15G7NIWHPfLHeVnzzIfhAS0myg6oh7Vbi/LqTL+hrbidHLo9qj
HqNEruE8/Jzd6ZS6EZQA6ST09pe5ZnspDVJ8YCjBEFzrTlLhN5NMLZlqC6Cv0SQ8
UjIcx0xvsNvk5uihvHPmiJMEOyX3ZaY+oaGFarEgJqMGE4ekmoPDBY2d+BHj6Lhp
2UrFZ/7IwVW2ruYWzWVES04OHNE42LuwMj5HeS5o9QQs8zSoSJFVPXi8h0wSnXJX
jTULUsSGs1i5cB/w7xl1b3TDUYsdHpH7PP6mkWBcgaMm7y5nEnu5zi44fTJBdPfz
qOLoRDOJwdwnuNyHsvq5jXgSORSGPSoP3wATPFlVzT7YyXIXyTKub++W41BOQAbx
3G8I/ADzUnfcu4NHcVI/BgrNFQyPADxHRKA7LleiMTmqWG3G45GvlGBQIA5ajTQC
1BMR6OLRAIfRotgS9X4wShiKuETYcMjc8InH8Bf1hpoYjHjn8QKDOI+iuqVwOOPJ
zlKTyYT2HartXHgb9TquSI2QS02H2+HbYc4zgChMhAVoCWbA/MFBnQqeVnkTCmLy
47kqs27IW/7OC/fSnmUh8Yjpbm+IVao8XGPYz/lsPH954gOUYPuG4d1+OgHUjRvN
8ALDdn4hmLGIsOODZRKF3+tchx31/xEwORzirvX/Wfl1tLX99JzW65z7KgvrjPrb
6x0M7ohHqoFLW8KEURDeWWpr62d6zxctaWP+iTmmCouAxxynasmuMJ5DU3mQ8TRJ
Q+KTHjSxa3ahnGUX4aooreIGEX/yx5SztmRz+SijMHSL/XKJvJKPrE6jXzjTb+9V
NfbdkV3aYYi8aXyyQt7xKI8tJJ083OoerxpJhwvPf1kisVQACNAGjgV9ru3i+LZQ
CiXPbvjPlmWQD5EHsy+cJNwpPM2FGj0zNoTbfABPMmFt6bhUEiRmGb8h3Yr+9xBw
WkOlRM/G3ywoQLonDAWj/p67WlPsuQiYFfdOeG5UYDZ90fid8P7qMH1NZREcJBAZ
XGRFPWX3YmqGcWAUtNGXyTsxk/ti+O1VjK1baeiSZ0t+vByHpxylgeL7DqExCGbu
Uv5JYZa3qfxRgVn6Rd8l/0b254fVSBHg9Ui4YG5bBhgSPFaMwYjd+YNeE2R2pIDY
S9xfDfphI41hEzQk4e2vV52cTsZYEF4hvPQ/jCxB+xwDiK9dZlBWEbxfV7Vi4LNs
Tgsb2D6mL8S1HR+pUYzOCUhY3aDTZ9yD+VO7SOroh/vuSAF5e2Ti4qjO8aGhw8D6
MBpbMntVPAc997z/8L31SSLrqiWy3hx/O67xxZ0tvQ4Zcsc37DTxbF1g3fgIgSdN
lXdx4Ez9JzJdODi+FI6trlGvefeQLaaMbB3MvsIUn2NvPS75IiVzWR1CH+P4xhFf
MtBYolTUtinPjHSIe4Olzutxz5l7OUkRdfwqRFc82WfwpQdBolu8o2P/pCdLLzJt
MGCd1StWWA9XYTECHPe4MQFLnH3OrMjkma44yBYIZF9xpaIt1jNDPCXq9U9dUDIi
0wlzEAkVHFNSie2pdakMjoo/8a6ZlAU8HISMK2dqUl0gW4lKybM120nvfc8CpZrn
Q+I/NBaW39rBl9bb9cZ2+R6yk4YX9VIPPCouEhZkxugyaZNd+xr0/qwUdhphB5VD
0OfrcDrB5S8OHqGEjPna8eznjE47KcoqncHs4yoRAfrAY908HkMzKt5ILecK8Yac
McKgsJ2Ix6Ve4ol3+p3hnG87qibo7GTnW4XussaJ9232kORV9Mmd58RAuQsNha7b
RQiJ2K9e2UTZIa52hNJjxxdqbXAF48c1Ix1/APG+CuhYxODqKlQw8hBrMEyo7Fe1
SOfRDYynEEYgxAnJv1kUy/UQgyXm+nbg4d7LTewOVXkKvUQO66AnOERnJZED/qAu
8XZ1iY1bC4qKeRWoqSc8AXRp2XdRjf7LdI+qyrBDWhdLgCQ1j6sYp5VOyxjdpP/g
c85HIz+xvvEWPARLf9SoZZvJ7gQDpu8SlkfnwT4ayrIXVEQxLTSZ0lSD0mbCMMfR
4/YjsYE8GxqwN+LITjj/lAzMg00dPCJzZn9ugbk5Y6RCovQbCx94x3+zaM0yN1MS
PeJoT5v+PUjLZdxARbyLVZWh4foIMpOQX1SKLDUKzjX+iCZX6HR6UZRrAV2yyMvE
HfGGlF97o6wnwdjtgl2TB9dgCp2dcukSWENd1AmSEkeQPwXEKOfhaVHdvPPhchY4
R1r4zVZAehEaQcrPV8MgIwJyMmwTOaZMxdhTa1Loj5E+ZUSbVxkyFxAQXUtOS9Fh
TFIUpvEUMwmhsPd1CFWGT3WVpq7Jo0yEoTkMpVuJm5AM9yLPK2A6L58UGcG8a/Je
G2KrvQmOpdefY/di7tvrXIf1E8kYD8sWFne4afrVNoYxjc8ON0R4rUYBNZF2XxI8
m2JZHXdhEL6LoFyVOv+vVbcEd4+c18vXvKS9WSxmiZoj3pnOBaVX93k6zMe7rDD7
UcszTvJ0ihjtdJM1Kvj88CBZek1i2v2MzF/yuT6OXduqkzwEUKN18P0qEIKswUxa
wMrzf9rvyW8DOgncIxvADyfxujjO9xBaWr7T1n4w6GsQlwRkvuKzXP6mgSlzlkkx
Ctm8ZboVpPQDzNekU1dRGMUIShgI6tbbvBt3TkLY21rYDC/Q8xKp+32nWj6M8Ekj
97eAEKi/tBPAAywlHRsdHafuHc4a8nZh4jMPpBFkLJXxFSa0R0JmcbVywSZovHXh
KKwBF6y28HzI/Hhb3ZwTY7jaBxHV4HmrLbdTBHzd7tt8wa0yrAhqNMdkf7ABk6yd
oNu21rvc+H4H15WK+vmqOCk+Jzf8xZqBNVuARfLyyOcopfIR+wWvkQaGfjD4zopr
h4j9YK4iGlk3P82Mek4mnkBKZ8/sRhpp2vDgMJRTL0gF7HordFZPz9esuWTFDcih
vZYsBEkBypQ+GvN2y1m2otqqO/ZGSX97g4LMVDtGmh5yVtSaSFP5BoioZtloD04K
7HZnL8BWSftjaiHVW/lpxVAgEr3eHu3cZbiJGXGnwqyc8VVd6I8jX7IZsOq7BOI9
5T5RFfh7luD1921BU/PRxEUo0aVtGHMpkesV1mSP/zAKyojQ4+rI/ybKy7om0X35
7vfhR7KfF84ij2glWKOcU6VqGz0+YUl7e6iaDqoKQc1ElAzqcKSbXTmnrsHqCbvz
QpyQ/rrt8y1KxWZA+8AJAGbFa/5sez1OgqrbumAa17MPS1qXYZMFX0QZuM6p5O0w
pJjvofH/JlJd6sJQJqJhEO6JR5K1yF6GCiRiJ2+K5H7e+iAFUNeeMouI80ALQZRC
gGtr6o5PY49ObhhtK7FIgDbyn2XC34+Lk0f8oMIttNR9fc9ogmXypXr0i0mQ+FGY
a3xW4fRTnJyecYfMmuSsmvSz0T7qocUP0bnxXQDLzpHwY9tWQvF94kA+XGDCmoBz
mQk/7NOEog0VCtxEi0xAI02uMGPgzXyLSyJsJxy+UFppiyq1JhTTOUNsIjlEDbQy
tL5Dq/8ayXuluheCxeq2bwZDiGvJ+GWIpT3wAhGorIqECkgBLUCy3RMy6gp5918N
Z/hwa87V+n3gj46jVJA1G9yCb4C/3mEeHchz9o9CGpCZuS7UkuNA6T7ooDvJ61MX
4DhAt1CAPMrliqngOKMSNVbS+fZGt2q/xLcxNhzCyjGVxVqUe1o2+RdAyiR6G6bH
R7g2aASViH77J0Om702UXgJpW8UfO7dCr6hCxzcdiEMzgpro7TJ0AizZQbRHihJl
jscpYPQyfJdVwulF/6GC+i3SEBIf/EiByXwrDJczobN8KS5+xEPO0jzg0GCu5PSI
0Qs+6hXuH8GlB59KJ4rgQouRVvDj5Ml6b6qFPwVdA/H/0CUeOxJXmcEc65leylMg
c/NKIgqQwLsZjnDRLyU6MxtIhYRLKN4LokzSYbwW9ADNzVd2pNFqounJc4ma3ZNX
CqM+bXkfi4Sdl4dOon9+H1R+tqYzDdkLF47NHFMi3YaGRIXnGlvTn1rZYoorMFuS
HXD2r0w3DB3V5uRqsO8YhwyAc8q/hs9K/akDtyInz8Ir0u1TZ7+gpOseeSGggiUE
AJvS3uykL8Wi9z0xJ6DlCfO4ibCyD5TMXA1tVzyRnYGijjX/q0X22HIWg7WHqa5z
2Qc5dh+Jzc2zktSOlM104AkFjsI9hMCiYf2dwiWcvC3k3pIcI8O7KTXw3zvbKPR0
8BlzWMXeoCE87UhMeONzGs9a4wGiv99AOljIxGij1ycQvqi7rBhkdQ1YrlxPk+re
sTyH1B7/EBJ9QE/30DsZyR4icHNv/2tp/yAeakmijTLkfn4AYVk/ocCTYrMNa9P1
tCYOdZU3G3edr/NpA8HNTMWqBOrRmB2R5cVPLWmOg+eLwsfdY/vcTcLo4xaUDoQc
NxkG6SfjuGgxGa/Y3X5jmCJN7A9lkJcxgS7XMbu+6IXaHgSUXQtL3czV06Xp73su
uFVaYDmBrdO55xWuy13qcaSIF7iV4Nhd0AifaImFm13uPa1JretRvIyv0J3WeKi5
VoYeafz/SHEd6ge5lRjFgX5UAc9tbUei4i9U6Q02U9nB2yJJ6EQrgLLeSAaW7SYe
EKkNsHzxiUId1uodOXldj3/mzPpsdsNZ/JqjK35eIM/FCFWuHgGFM6RsOoY/3iFw
R9xFo6kl2a6uvTmKNNz5+NnNXga/Tqc4eLQPAHyxooA/cGG20R+f9UT3IA/LFKVl
iF3dTBK+ulRV1ZPMa1CguOO8K5NzexLtzikkoN2AuUsyRD6H8MkoPN2vd9gmNHzq
7QrQJp8hOxngoPR0/2dN/h1OADKLy/WNbR3NCHvRFgX8d9eBzbvzvWDK1zghtW1A
WOuvrVgOobe4/HHP2JzJ9l7uoexDngzjd5HgL2a+PYxh/9tBryi3nOgX49J6ULyl
xOrgO8870dL9/tGS1YeGJoOdE96iQiYdYivJApLg8hiXqzy9ay1oi/IwVc5hmDX+
2rpr3/rtl9th15h2VC/IrG/uVFbj91PQ76kf89iXtpDvTTx4aYHsj2xdYsOfdkk+
cfDMtJrZywR/W5EFWGSTTQcTrHbMilLJbs+9RrBfARWSnd0kV+cLGW6pbfJywe2G
nO3XTRgEPBnci19BzLJrKthmpA1bYqVwy9ci32d0ekUswhNSzobg9HH/qyLgy2va
n3RUfNMYz0zeOPUYvVnPgJoEiQz04yUhX6b4cfjfZ/s7OqAp22bv31u+4uhNiRLf
yTkolL+1w6jHZM8IwyLYOx/hWtJmauDquvTHTvWcRKoBmtZCgdg+xNEs0gE/jW3y
QC6cuHlcuEbQ9aiUGRrjkhYM9jaJiUXq8yb29tDZwo5srszZnGlIsy7MFyc3fbeP
7nbIIP+L545rGNxV4GPPL1UrmQFyeuCdSX0QfazEOQVHFp01BERXqfwd0mUddSBM
sdI9vyBnZRaplCenprQbhv4SDIkZhq4ezZwN71dIqGKyUw7d7QKN67ucqlUEE+lP
k+I3zh1NFr/zGMJUlBQdzWS6zXF6V3b6leB4t0m1josmicKI9kOutLHUttttn5Gz
GLdrZTgmjsuwEjB6Rd2CCwb0o0/ZRkYjAvGMuJ2CISJyULqEb54KEw+ADAz/BDr/
yJW1XJ2Rye1gNkuooPcdBnSro86aZAxQBuclbvNaAzrkAVYJ14CadQLeJvkZIgoR
F26OGz96g9UgKl203UJG73tY0uMM9hDcvjHqV+OlByAVriLNHzUnrcK72nD4hCDR
RS8htFyExEwGOZslZBhv982jZ+TJxPpuolI6j2EV+mRAO4TmDjmeVsta0kYC38ol
saWHqNr21v5iwnWLR20opUpVdUd17sTLBIlwCXpJcTSlRDgnnOv7EciGjFc3ki1T
+yOLVj9a9IXCzwGnmKpPWA1uyfRLAbkhH1z58TONuV/+jFD8fX0AmNr4l9N7I6Mu
eI7NzREJNsqz25d7A8N2aKl2dCaDqHI/PF6NVweTjaqwh2IOCBFWFXehnhpoppQC
1/FWWRu6+ijvm94YwRbst3v2ImjO3HuiWJGRpJ0xj+e84/n6PI/j/demE0AyTUCv
F5MIMoGw0p0ZmACQrOR5l7UrWjFAJbQwDRXXe8IwUS+rSh3LbSHFvzeSjBb1gCY4
qRaaFMuQg0SSeQZ7C88d2BrE7zTk3Jy+/RoVnHXl1ixu148SFt6Z2dd9Ou/1+zGS
+6kPPlUP5hebxNvdZtfS9vZKJVlyvJIZiEsq+KM5ISiHwmFCcjpyGosNUROPEGWQ
hcklPLeBjKJ7ius8+TbpmUuE/OnhVdJG8AtXGRdupZJ1yBND3KZ5VP6L+Pda+MZc
q285kxKHbBPDTQd2okkO9CeDnb5/TBVLg/vkvakLxEMbwvt52FCUGv48L7WqegRD
1FhbSZ8QB4V9DHoLNPAExOgQYy6Zx49+wx5cRB2PHlw/eTxN/an/42l0oo5N/LVf
oDvUyU4Z/L8FpbcUP+onVTIgqLk4KZZLxNn64bZAPhR+mZud0EomO3HMyiGEYC2u
20CtUtwwwp/QIvlyYnMu7Rxj13yNrP3kKopHKeJi73ymvzKBv4x/9ikqVv9gOsFo
q561Sn3SMLVhH5ya+F66//+fhETR+RnQtYzOD0hGm+7maxBFN23CQWzK7cEbZ0cm
7fJC4qYCE0MO3RDtlABfW2AQovuLgD+vS8SNNeA73QEES7PLEZ2iKGfHnDeffKLN
sM1dwwWYKXLeZixsJccpyfXBq19Kq7kDww6lzQmmDrLsU3ycrWWw6DA+qQAm2EEx
9CUxPiaMgwJFMHwBu+8m5VT5Qn7JZeeG2iFRJU8NDPngaaLMcTtW/ieQG9zggQ24
Tm9SvDjeLfV5qwIBwhW63FLPgsNiNxiTIT0Ai2ZgBQEpSScr6lP28qauzuUZv7mx
bJ8Sr/VPq/g8D/Jp5okvh9t86LL8zQHs75L2ax9buSkdZX+sErZUi4oiE67M4htU
Y0tA3qbcp3KIAMaWsbhoPMB9q6Jysf6obByjmGfCRhlcmd8CQvKu6V/VHPGVqdFB
T07HSBgHHimUEzsd224NtM8dSqre2+WPe34ltlxPMDdnP8wMwcFnTgFK93ZKIEPp
5FYyEiHVgCUAM2KDROZ+8cNR3qi58yLkqJfKYoE9GCjjwB2f0o8kILmLf6toWbTi
KjJm7HRUxThxITMe3XY6fjQ7h6sK+Bt8Y6BWUASDnvHB2S9mtMs/kMlBj/wTINfJ
zPLP8MxBbKyjg5MCxpxxdo6EY+I2iwYQdd5qaaB6CUitcxiesU39swyzn9biws5p
GdqyJ48M4eWKm5IrsSP6djoSVLHsei2aa+Zjz4gJPhIncorKLpFDnw0uME8Pjb8b
bIATCKuNnXLmGIqcMTVuSZiHboa5JHcYDwDWcCYQIhfii/DHRczMtsqEJyrs50bc
edSOwnWNgLCOcc8V5n/NFr0tQnWZhp2M0AfwiTliBwhcoRcyx79zSTBUDxs5LOIV
0cg4uWxw98uz0ylbksrc4w2j9C5fMTQK4lcn5XB9+HCffAENSxiC2OY71rDeoOC/
+JkdvDOtbcxw3kTED750NkY7CpEPcRtAVV02XKyUhHnpYTAqKKOQXHVhzWfIJJMK
0N5ZIdQLcOjgB42lG/zoFNczUKaHvws2ZXKsLtuWaGBmVNeSzASsMoD/7Vkl6xqT
OnwfgjW25ztKr+v7Zec1AQZpiwUB94rKBU66CXXxzOALr9UphSSqpLJ7ebOogFUR
CSgHUvGAe5XwcKLNf19ulV/cUPZselb7Z8mfPXplFsxOPJXuXyZ8i0NSTjAV0D/h
5yg6g1qeCfaGH/RJzkrEvVVAhI13LO1NNJ3GfsYTuc1P8LBgCPDjJeRKMb7wzYAM
r2e+54MyLPqoe3LNm44uBZGMAvkE23ew4vxNEaqO9PIYr6Z4jTQVm7ocouVa4Kq2
NmTcn84H0NPt0yxDBgq+8rhi5+5IozZ52LaIHAzTUJ5wL8hfPdXXNUNqiYrn84WC
hZyAEK2Ot4lbbyl5klCzAxZsDSpmrr9BSx0lC2FfmYZQjM+ErtuR1pZIMuZf7/gZ
jDKhvnCHMVRSKUC7pVVWIGNaeWCHofVvUnWDfwBtm4qxcj6lp4Z7jxQpiWIiPGW2
4EwQ5rDGOTUMTJb6pDcNgr3WkMiRWTGNkhM/x5evLlQuIkUi9Ildd82JxqjKAxQo
08L0xbb7bxY0EKwgB68ZoBJ70m5DCaXJ1uMkyshnEwXnBJQ5G7UVrUaH6747oHCh
a+veeebSiRIg24HI1S5cpUxSl9LpayLwpHHz6bj8kdWf0agVoeJSlDj0o2iBm2Zp
ie8PTI+FJ6ohZ2IyWxv3/Zs6FmdlhRMFXp5VNCWQGXOlQ63edZW4Y1SB15aRtoNP
ATErkgZNqMkXB8sgA3VGwVsw6PjXp8lBG6fIgfIH3ys1yvaHjjjv5TftDN76Prfc
9pdwK3h2QenAcjMcvq9k4XOhctvUrOI2dH6qYQXHXBzNEHWYjZClajxeUsbtOX/J
nVrt5o9HNqPxUx41SuwKkuVFD/5R71tTa3VdrAItpnAzO4lkNIw8H0v7V9nxdnx8
Ugyyb+kLVD37con6M9uN9yC+VISHRZAMs1u+p/b+n5pso+TGyGrRfXUgLCs7hYhs
gvXE6mJRPzKD6VdxeGCMuW/TmX44QPJCCHVNgXTd9HlHrBG/HP147cqAXxg2f0Wq
l8j7rZk0n+GBncfGLN1oTCnbS+HinfypTNGHkNPyZyIzpEyeuXoaqHI28wnQOxCs
RWDjdfNqIGJZxSVEUcABWp6DDED8ogdMjlkA2QMmygro1c+XpxXOG+Elo/uAsRaz
4IIWPfTRd1hU4AzPG7R50MckSgnjTCq7Xci3Y0QNGg9FrMmu0LA0kysXxu1TQ07M
qdg2hdDkiQNBI07PzxW/TTXaZKGUEhA0uw2PB+K8UZkI5mLjpuJ+vFeZKmtxR/e6
QjcAs3SyZJh04e/mylSICjjR6XG/ypFjHLzWYW3q1NDhiPDmN9yaGT5as+HmyIPY
AHbQIuM6ywxkLQzdUlgEoU3utUujccBYgcRSYVj293iO73gGCECicKy7eXuZ7F/D
Z37BeTQ87Lns0kxp0m1l6dGi5G65C3DLux/1HO/l2k3TI5nrvlSXeRYOsMYyHcky
kfA68Ex1juAFargmtOlfM1cIb7bzU9dsabTZkD6BD/xNB2MAp6EsHHQV/9An6G6C
JxnD80QS1fbrT9H+5/JXKetmCHREPTGkuEVVl/08UzF5r7GbF9Da+2cN5qdccwkU
eujI+KdyxFNPhpFG+NLEVe5VW9CMFQ7Dc+OMUl5RDWI/en+S60N0y3IriyjNrnAq
bIVD2lW7F47AGkdReMLcV57XLacEKQfDV7r51mH/5riYkLcklgw7UO401hDYqjUK
niwRU++qrfg2J8lIsOWrTSVABliguOIqpkB+F3oJ5WNL/9/T9ASrC6tpBZTazghs
pFsMpEX58F3DueK5/abNxsuRM2CGpsnLTXzuzq3VBOQ0LF/RA5kybAkirWRY1bFX
YT04Jf3pVXZxljH8ZcNHhyLHgbLIVFVfwBqJg24vK+BK8AvT0mv3Py76+DjAzXaN
TM/jecuIBDk2l0UMooPjmqtVeGK7lrCexF7XmZB0iceQEywcWkGkS2K6Gy095OfR
YeHaiqCILW+XVG70ed1u8y9ecE2TH2tvV0giiTlNqwB5eJegQ+AWadwzR1aQT0cB
lZ0vGvSZfXCRk3Q1lbVM68eNfhBBhQWRr6u2IF4ohCMKro7plh4Sg9UoX9c3zMuE
U7SwHikXuOhKTY40ww+QaY2DkO2bPMsTiJtPQfao4id+JcGNPZiavVocoWRjM5Xp
QwUyFA8IqAzygOo1LxbJn47XV96xng3a9Mr6R1FrWNh3Orh3HyP+buCVVx5dTu77
eVeRYIhWCatsp3SiYdaZ4fR0M85R62qzUfOPGfo6obMjjZVtXL3X55lxQ15NM3Ew
yXcxetAU7Kl9Oka6tGFMdzGjFdvB8dDLRHE8UpnlP6sCRLA0LQdf7k0AjRGP3LvU
lI0SFyQ7hrIuBIi6/Hd8cNrWZRq+Ed6kANUMfp66JpLhOkekrhm/YRBDe1/0Alro
SdFEMhkXjpvGh2PrDa1FvHLyqOvia9miX4mWuiEFOE9yWqvNNHqiXpjSXCVL0NyE
qq0I7xcnafqiGyhdQxwm0fsW86tiPDj81LKJDPUnVCHEOshE2Xmi4dOT6YldoBpH
R/o2Wck4irvYz0f7pYXJ354hjn7x+5MXAIdMc3Cn4/p/iwpBtzzYmwOG2LjplK2T
1eycRL5oA7Vasm4xC73CM49LhnVbPr49q+dyt3qcYtpPUcLf3VCnprrB4Q2eB6ST
ET1iUBYyQOPEQoyC7UyMvsDoRpgwJgH3G6YcO9CDRZTnqBF7ga1wYP0uR/f674dC
O4Yq17vA/+YJqSzUUHf09Dtur2iy0P/r7naPFV39ipUuqcLwxzu516D4NnhBLKhY
vrweSLaiCD6KyUgQU0GV4ZXNW4MyyWafRwKMXIqs+bI4b6A6SZMpn/nXxxS8yo13
1GiX77TwZ22rfsQp7ck7WWdNuGB8q05pekBZZEcn3vumL2p0HV+8T289yr+HfpRM
OEQ+MvTvkp+8VfiJfiqzh1Z5odJ6g7Za+b0mYwtZlAQDVdpvrJXKpmrHFug4it9Q
624muMkB5I5RYcYck+1zePyq2xCzlNY/uDqwYUidRJTsOdlJKJPCDweF1TohpGxI
qGz2fGH/18VdYhEPQ7GpLT/pL/0gLggOQri6i7+s4VY6L6eXnmMea6l2wl7KjDKp
MGEuzmjrK/iJPPXDxwoNByN7rhDSSTTUPCPJFQazZomVQivC2NmtSd2so8kXIv0Q
lRPBDCq3aYfE9fZEHUyxDHoEgHbXNWBiG9njBmECJiLb/N+DRUq7NK1zhNqUVLQ6
1BjkoDtxlUlvJ4hPtILWjYiLhGZsvxviJCIGwGH3bq+1DeIQzm0JZNO20ujbe/1P
QB3h6dRMZdlgp01TiVoyckUBmIk1eu/gza7Xxy79+7cciBppRQTvxMiFFzBp/ydL
RwCsy0oONqcHFdiHgMvJY/hvoL06sE3bdeLeoe+eSKgbkgAvR8hgplVMxN+WTnJQ
+oF3ur5eMl6ndpKdTGatbiZj2XRNMmtE4emup4+G+FWWnxAGr3XjcN2iuE+4yBhH
VfEeGcoHa2DCGxQA03nOaTg3mk9HXdiZy1AJLzUHifI4cmvu7QolwGgl0m5XgGZg
nvewkF22Q17cX0pQkN6K9J9Hgs1TJpRMrVJXRY0M9y8F01A+kYQv9WZaFoUFpbZx
vwzL9Pesg1xb9hcN+LAujfXVIynokfx66dvbrUhsKVvyjOgfcEpH/DihxtiwDPC4
49i2yVQbYMphh8g8rNEEV6X9U+SriwN7yJ+y2Hm/G31TLFbPfNearRh2pa+VMMec
f8KsMblwryEjLmks7fK60Xt9X1oKhFas3vCdsc9GC7DygdPJTwkY3WeWUq0VK/QR
+S1x8Ebwx9bGRb1TE4wSXXSFpaT0Kpc1CDldaQDoCoTywcCgWWZragB8uV0A1eKX
KCR6pBkJKv61zi1y+Hv7OKOF3GHU90AsfKeFli98Wnj211X5U1YY/1KQSllw4XDj
rljXpreiUDloQ5Ou3dEKqZ7KdWttU9bMfu79XAbjjkrdfV9yxpcneLXQca8InxPO
8I8Cf762BU7c7UUDKwgudRSoka50mTy4hOYbJAQuMTC4JFTt8LUqnSsaLW6+ecyX
Za3Fxs49oZgmn9z2Jkh9nfvBZw0Nv82PmNAXWQSWVmyStZi4BdsVlh3XEHTbbDv0
NumQN7Bvs7GtweGH9ou1n3VPDNS1wvboK+GcXTN81rUtChN6xnievdrx8CMXPt5T
gmbVIGZjxR1r7PZdgDeopp4c3E4UsSRVnhhKZF0KjolJJGV9Wp5Z+8oERsuQEn/P
ecJkkSG/hPhpjEDeoTMWagIfa6l1acu3hvVfDOG/d3JCtJrOYXDTK+VF/rH36Jlt
VPgfS7j5NVaGsBNrLpoptPqK6LEQWPktO1uYBLTIfSDF4BaDtVEf+v3G3infZinx
SgNk4IDwXaCsFGAjc6AnFGFlTsuFfzRqFny5NKxDX3+74jlQSAkxs8GwNi95dk5Y
T9rPD/upi1E4gGebJAGoCerKV1gxl8XKUw5EtSDHD0h4Z1PxCNVcs+CSEwdVgz1G
SGWQ3JXif8DL/2/a4dCsn/pd7SmQiRHhBg3VYGaTIXcYBpIvpGdTCkJk44z3p7Vj
5O8LRg94kjp7ilv98GkwYhHmOKUsNDdRIcprlEQZxCTAb1qldInyeTlALjXUX7MC
BSuTcJUxn+YXuEsXS6xDfns+cifEXQb7Z+/y4wsZh0wsn2Ckpj0leoNGa90Wzpm+
vnm4QCPz3+bxBnYYCS6nBLZ5P3h8M7M7NPiNoDjAyE9ofhF06otnZHKZkJ97P9rS
+DkUV+F+NMI4yTaY19COD3tw9kKpA4nXX/EiB0cMlBg0WaI6uMoRs5DbznNZ29IE
1Igr/WfBQYQS9LJZIhESYDv6gVuXtQWdFDygM/BeWFebuZgkQWhWUO6n35PQeELz
9bXTfvsO8Bf4q0xE0BzYOmtxJG2Hh5kn+4KXHgzTYjVMPrxSSxmLT8RfBsVyeQy2
25e/lZgH/ppsMMWeRgNzPYVE2JvOUS8rNH1sROL5XRIUga9ynxuFN+XO9H4GY5oo
822hXfYWbjdYUXD4iiN93nfaPZc4Ng4Uc1PN0kB/k+ZioMEyY0K7qW/CvRvjpT4C
5yvE1Fpu27RV84xEjj+kBrbhTiNYpnyzC3GNnRkBwK6qY59Uqv0YAkCvmmNM5XgH
+e0L/7xt5AEALxEKp+eUjyvd8RmaaSDCd49p53TIy6vYRm5ZN84F7X3q8tevkUj6
B/R9QglTmB3ZvIaWzq61TQeZG0mN36gXN+nzwlmHVk2diJW1wjtFAg+eFIDv9yhM
ldSrUFPDAXZb6tuA5rpj5nCfUpBmiDvg3xF73kguiKQn9Tl1yfSRgaiuelpX2x1f
yQXkGoVGyIxBbrt1M2ckBUlGuBWEXjWL6W/J5vOxKdnly38gQS+Fu2v9iu1028tm
Zsp8seIPHqRsxrGXnn44fJ9+CfIEk9AO8B4UJM1HuevlSnMn62n3XC4iW95gkBSp
eTrst0a8YyEyxqA6FVf5S8lVSRG1sP+SOSTqkINpgEgAdmacwwrlQkReI+kg3nAD
HrR1N//OVK7XeGIRzBdm7gq+CrLB/bJD1qT2eO5Y90tWdY65UIhbOUjjEiD3md00
9OwC7VazcGupfXlLRAsMxtgUnUSn8kNALixqkt204dbYzZOKt0m4Oil088kybLsV
KFbzWj05jz1S3FrTGxlQj03d0jE/sfG18a+GtweTabwM13+RX/Uj+Nx8H2zrhUVw
u4TXg5gsECZdKkiPCnf+tc5sa44jZC5eFNJOFrgzS69nXivuaFkwRQx0h7SFggGf
VVh1D5ww7v3Vj/Salg4Qp4wHki///JGOqEtQsqm6XTcYM2qXENmRkUbzi7mc+bZB
ljc6jIi3EXyMeO7CMnypmlwGFv2glcp2hEH9XBXRXNhVEMTRv941N9QQq7qhUFUb
B81UkyR4xqwasSJFycWITjiHQCL07zTJDeIYh0ZrxNZuONoNFSho+Ljx+z87GOBD
sbTk88avAFo1ZSS4UyM63QilkwoXr0gdvaWaCHnR3tCDj0OlejDpauW21vnuGyrs
AczTmiCgkkWrKoNJXtpcN4a1M2bZf+Pqqx9LzKqHXcgRrtKJp9UW06LpswqJFoKC
bsWvdbsFXjS1M9fq3ji3jdOoEEJy6kNWTPS323TNJnZ4xtSm6Ci65vPMrYCwPKVx
TaHSKjflpKGs9XeN1HmlUwgkV4YHGtkOeKTRoUKVEyuFQhmYAO9TvmOnIs+YiatB
61DJoMQe6ugafyJAx4DbN6exQcMRmskAImrNqdshCmh92mEZTgfdmFihy7PMvH8L
Jr1vYkklXEGFaTo70S+6tpmzNcywrQLGLbN/oTKxmTdruKjGNrV3oeiax5EPnvt6
eSHLrxWB7Ko2+8XY7J9HVagK3oYTEFmMbJydZe+glodGv1WQbBb5zexI6pcIAm9e
KfB9TlaptJF7qNlQj6uvv/nIHpgtPJMO8mpWWcfM0v4AzdguRDle3KbxSGfRqHHA
SM+Y2Jj0KEVXlLcDPTKxVGV7b8ioq/4HeIBJAnjxjlR/H7TJcF2gQMnVWt4Clcye
XMZeV/qcBiKxM70el36eUtz9mwN9Qo5VkbW6dTESR1rQ//Rzuh3XM81aA627WTj3
PUuJ9NSkLFyjMdkK+xd6dC1E1K0BVUyO2LYiAf+97uGBR3h6rV7hVbRUcrZOlQ6m
OCilvS1qga92GCQ1dj7S1oQZS/HU0EA2hjCLC4GcTSFRTdHjmfm+0Zx/lwUSfQj1
bhi4umGVPXHZGvxlbxlXvOOWlUa5uRAEAEzmhxCxLcOqI1gUr3A0UZ0obmug8S3z
yIBWLX+MIcciyMxQMHl1KNLi1M5AeKnJnYhxuNQnCEI+/mLGAOtl8AeIeuSCCe3C
aFtOkQ3E7z9KZAafr6Ax71Wi4G7PuWQfYFaN7dNFg7C2V03N8h8guKVbeJNrCiSZ
KdCzzZeyBXGKXiSY/gS49MqjCEKD2LKDBHzhN0SNh/QHGQpbgaKr1FB1I0ibC7Xe
EB1RYIq1kOkp8azMcbouZj21XPogForToZxBJ0p5KyBmuTObpDsz7lXbO3e3Y+CN
NSFtZgfGy1FKYo4fskPSozMMOibl98iYbAbbVJG0oMpVeOVohQK8VWBOcGzI2LFB
S4hj+a7lhbYRAb3vsUkIAffLUHUophyqyG5VN2Md/CSIZVADw9OC9zERykKJ3EmO
xzGwGJqffrn9nWTVT4o+aijRdMypiGAgUYm8Mx+cv3bFo5hWrelpZwkBxNLUzbnc
9rVY9Cpz6NYO0uGg4N2+qjFn1Gw1ABL5w2o3cW2ropYnkwiKtKp8i4G0qNqW3qNM
ZAnQbK5TDlllD/6rqVa34l5rWy2M8Ap4Wb6/0KU/TmRJLXw+QrCoBqAa12AMDPVR
1ZQyCAAid0Pg2r+DwbsnVCzyG8yQVHhdGlVjohP71v78Y7Y8Wjo0p7HCWCLMi+QZ
CqsWLY7KRwErwdYDcoKTBFbYWTcDfzWCkDKA0fjDn6w+SWTX1ZrPmMo+KlBGmgaM
iJ+u4H3LMwsjwYoAeQVn+jw3i/qhlbTHTig1aTyiTzMLe+hnRhZROEzz6JuLL0X0
Fl7A8IWXVcXI7PJakBp/F+xRA7wvbSy/gRkgGADTcYy9Cpq9qCFvQCT4sJbH9nRw
dZkTJ5tO2v6GDMJTMSqyqMqf3Egiw4iQWBYs7xCeEVuiQ81KkUehsT2YyiJofCI7
1SQYcRm9s+5IKz0mqeuzn7W7QLIRIQEyewAHf2H/n2qHFgtICgJX9sqn7uHj9Nft
aQ7uvEoocRZQlnl0ID56y9s6koZX2bJdL902C8G8BqnzASq6sbnlP8vUWCdvoktl
vxD7ahUiAF7BSgY5uFsjFoQTvInrLUbLByH6PVr/3AObaqsQAk5ix2Ed3WvH5xHv
jwD63PgMwUTfz+IQsCdqC3SjnTCazpNsyQiVu9BMuhIlcyI6S02yIJDh7H1SzQo0
viysPo2uifj494su7vEQUBHdx2QRo59fFzDv7ZxJ3jx5KfwB0knv0we1ACi7fVoj
ptyBzE/vtrfFnzzUPTG8e3XuqBqPF47cIHpVBMsLTOOCpzat8o6nwrsDRat8QPBe
K1+CsgDqEQ5L8dLv9xoKjptjZxiDiVcL+bATLtVvEYK/aok0h/Ar908HiS7umfzE
wvcGtuUhRGeVU3Ia214qP3DK2a/Jx8XwvKeeSQ+ZAvRk1Ozkd11+ETdd17LurhWs
t597XlrRTi+bDLOz8itYro0wHdYu+RqpoSH2tnQ8N47sl/tL9weoGAlyjhFm5RgE
9r4eLVmwLdRNqEvM3NL5/EqVV1qs9aDNTVy2zdPvgs8z6AWmwvExCRmk2sFOMEMV
LbnMYb5gVed9Xseuqah0HOURfHUhbklp4+VD5AewabYBtF0ktGOi8WZ8bCYWWl9n
JPZ35kD7IZWZ4s2XtZEDM2zHy969uySL6VVARYhHCctP2D4k/5efMveYYntG37X1
8lnPFfs7uNvdaAkauxgaagpkIstdVAPDw80A98adsx0ocyvF50NUEicn/c9rZ/Ip
dADkPbC6zO52C3TlLSVhyHXD/b0IyYdBg8DMWa8vwdkL/V8YZ9bOoWT6V+uQ9S1t
GR4UOyohzEth+x4q0avgk8ocHs1pKXfGswRWmMgi7oDIU4rTfpfpS0MiKN9PxDXA
P4Xhuk9wRUujZcIM0Qbp9oKs7li1NeW9PIgULWK/4GPXlKIC+GkCXSxNYqLiNlSA
1eOqgy2OAEF01dJK3pHhE+ptwPpdjnm4ycikdncqz4QhHH0C7+282Fa/HYCCKqDM
nRexB0DShG4dmhc5zQruJrIRmQlTUPlaeO9vydY93pIUmX4LwD8gMFERHoyw8uZt
fWYhrCpeZ63tKj7OwmbQijqLu6DzGPOVxmdNQlLAguJCWB7BgZT3DQpRX0SqBszB
2V1PEigkHWLJyPccjHwfDiRfn7Wde4lgBn303hs02IuE5cMBgCqL80kMNMTOoMA8
IZojr3jh9tSO6/GCZ621dINygINXJggpbEwCBlUp13ldmfK1grea+npm0mHtJqq7
3jnHIIh7Lr1riKMHYSOQAq9e8XRwtg3LOE14cMdvAkPtr6csfZcXKR7ynh/coM6Y
7xRF+Uwea8rUO8mtIFFEN6V5eirY59vUZF53jOmwcDWCUp7PUWdpiRsOayRHncES
Pjb/AVHcG0KfX0jI/mP1oyyJw25SbBqogfU17cxkfE3a9fGkqgoIIb86fci13DLA
iSpmkJNY1B8xYx29XPTAt48S7s2dVAR92yJoEET6EISmXe5E0PqHrfZt2VrLQUG4
pom10OJJ/AJRmKSaFkqskJWYtttwWwpZdHFr1axT3WfrManCnNLZYVR7bXw5WPRk
m4aY54t5MZ9AhFF9w+OI4b8JirOaZFoEXIi02FWAFxlyM6e/5Za4H8kVuN+AggxY
6EN4D5Api98stAJ9F84VcylyylTwVJ6jriHuaT8uNwHPaKLZn6Y3UnzgVpPr0Ri3
npLAZMQCRWu7SOdjwuih6POyTZd9jxLQrfVDPooJuvtGurBbpxaewA0aYVj0bOJQ
HyXQGu1j1Qc8L9vmjFalJ6Ew/d4LBE0G9br5i6SAW49exkNujPbiTDSrSR8OWVgI
4ctCbu2Kxkz7WJbVmjcsjCreylmm2QlDWW1fAvmoDpgHzglmycGVAcjZaGiBCjxc
ts3HyEhGVPpsf7vqsCIM+w+w1f9bqWrF8ikBZpsvN9gOaff+Tdu3hZFmvqHPvqjR
eMxzWjtirqepInSwLVcQECcIJkJTZap01WaSEzgtpNlkw3D7gvVhkAJcq0bke601
+lqayFfH/lwI+1ReClLlqKMWbKRXz5bTfOsq53PqnPb1XIyBFuQLUqpPGcIWETT/
J9kX5jPvt21Lg4mSx0zyl8Gf9JLr16DPpHosv+OJX1r7NLwtO5GGtS9tzMmzAmY9
A3yb53tc5EccmP//kzZu8mLjYJvKW8SSxkTqfmGmdzdoi5UJQgbSBubdAFdQnGB5
lyNMTL4D0M9r/lkQ5gp2cVEvr0rOuVGrEbxpKGCXpKXMEgsec+wEHkVYUd0wy/kF
FDYUoE6lLFfWB4BsZmVqX7vNUcfdudKpaSlmzRgmvmbJown+4J09IRdNkJ7bbNhS
PahZtFWW3L+a4bYScKZACSjFnrA7vx0kmOnlZ4S9hdEPzo9lG0PiqURCRed99gi+
KDcMvvmM3R9FOzf+eott62bHNGMH7sethCSQEEf/8KUl89u2cssCyF4U5tMeYs3a
fjxB7Her5hNmPnVHwQZwaXj2sCiO42gPj71FVW9sO/3qrD6izaQ0dB9MYoAH+YZD
M6Z5Vm+ZG/tpnUEkV0SfQFt/VRi27XN5S4aIk95fd5skXdPIsaJy88F1U0dVgGFd
H+qhA27/L+5cCwiFfULJiNkOkryHeyLRNzwGav571d5bAYQ5MS28zCR8v0vNRaKt
g49TQWTjtPOLixcHu67IMdXvCIYMisa3dgx7bCwIRqZqWNi6GHa0l2+RVKT8Sxkr
A+wNaj55ga7zg+2bVdCkTKP+n2Rtg3H1tMTeL08PxPW8oD1+Qt1C0LOVESMknBIz
fUZ3t+KM3gg5HWZ7TGZOyEoj22JJbuvSsQvszXL0vuP+IebO0udjus+bIXkQP4b0
eGpuPYE7ZAkqHK+CzucgmWnCDkz8san7rrzwYJCJ6qyqRg1ArqHwZybIebMtXpfk
tqh6xiMBO2FswiRkunY0pQ0Q/IipQdV1rA8gPtqiL9vlz7S9VTgGJmFKJTfis42f
p3Q79pHteFnYUAW2aUncCBtTWtgOfiLzk3YhhONukGCjbBMYtLQDgAGjQMTibkU9
ZZVohdpmw+ipEEk73EMjyMzRsSF0oMZBLTd8KZ34gQF8Q15ps10Kf/bo18SneX/4
0qZMKt90KaAcKNlK7T3kBiATLceHJ+fB9caWvEiJLuz0lw/JggRwkM31x7bZ0UOu
6LhpqoPYY8v9TSisW6rCdxp/Gc01htSyRPFdDJC/9W2wl+iTxgNfX8du5zkJa1Mv
bZkVgZ3MmBf9MRHjNOPB8A55ZaQZJApQbqO2OgPNOn99y5NwYYPzzdS6nfQRwz4S
flQ0T3OLAbZwChdQ2wCnWOCfV8IZxTL5j4M0imFjOA4r2VNQJQxRrGtkZyHCirqa
wfrdenN+tWPB1nfNRNffqjxuHz5yIeWm0N4m+p5NO3X5OxgkNZWkNSpLpJLPK5o/
duxbcVkWqBaYv/KrHTZoh9i627SQEZATjwrYNLw0/WOAShdo8WdBzuAhiQ/b/K75
qrNeHRuLwRZIHBUp2EJkBROv4E68zUByNbSfOEA+XcvI8gRDEKvzQmJZCrdLrZ4r
Wx4RICHVr0tAuGVXh9B/UKlLBVPXDrZywEzbWla8+PHCcR/T+MuCEwr33KLCcbqz
mc6CELEZQxcZOEODJ2eISPcPhtrzOdxfYKBlr/xj/xZkpPTg+KGxko7C5B28CfJi
0NQbAKoHud2sXRezTstJhuL1vGqAxwcwgNPBZVL3fWyN6dM4j/4SrEmVbj5B6xhc
wsFHeOKUe/0yQ1F2KPC8UI5VJjlvumY+k3zRZ9cUiQjwFPZ9BbDb1gULBIxGDafh
3wfXqCeXEDHNHAPPB07DTIx9zhgM6uJDFCRFtB09n1NoWYhFDvz+jQxN0JUCWsl0
zFcxgJeYAoNAwoe6tkytTVv0YTJv/L4kbc+0VBn/6sJ0m+56WPzVBPzuSgNPuTVJ
iIOWSHa9LvTYBNa2Lk3OS/yc8EThDbbxv2BIS9eyyVUY27ho16O1Xc70byknuyrh
8UyihDXaQdWQcltHqs2Xt+SrRfbQiodlY+lmN0V7ypyknuTIc8ir4xVHTDGS2gzP
3Nok+PI826HSegvuO1It1XFkhx/2+WrByJdSjJUwK2A3HXeth9yl8ChTbqZ/fA+v
QJuNJ/9wXIdd6Rqb+MwRTrefj4gm4C0S6TRu6MFHRIUhlJWX4Q+/HhLjIDPsENiW
w1cS1MPzqRsnr34ETPS35q4hptX6bajL/l7fkZuRjz1aCGQM28V2//TSrYg6RjVL
/dkuZtny5q5XrBW1idXsY2jvSMxcgmDtWx4sJim+Ra/c35/+A7NCzi4Ncvz8p1uw
/ePU35eSXl6vHkItdExwieDERj2MDrbigLPOkw0TLX1tL7BztBWREm1jU1Y3Gt1P
oY8W7n//jw29cHG4if875NPOHRfkOe8i3tqki+/fC2poZo7G/7KlYSFC0wLKRw8I
3Cdq9bEVxFoTM3PcxLGiG22vryJdCejwkdfrVivpLnS/91GvIekbU/UmkuFsbhGF
AHl+htkyA/aX+Zn8+ykkssC5zsJ20J48oeI+xpms+ACJkwF3+V2q8S1vahP8ADpi
iSvxeiG6I/X33zCz3tv5C++CIEsWQl+AkNirVeSrpzGsPgj/NUApFZu5XK9QrgrV
G2Zvda6zu8c7Zy5oWzPhAkDqsSeg7Z0c0foggg1Bm/VEt4VrBLlf9/z2HpNd2e22
T4vvFlCVpRI1X85F1zQx0BDQ2IiNjLvriBedqzHP19JM1+B5lWE1wkWT+Ow3eTt5
MoiAb83GeByXRR634zPGqa1gRsiQ3zVgOABKghdw5CChrRkhP/LFgV+rhsRJJCuw
w6z+CNDGjy1Z8hcrOLCoJeoklNWB0OhpNQ3HconhJNL6ou3Iy1cWviUHLVaJWAcB
ltTgC5fXAmJixPc/El2O+y4Vch6G83XdNsbf+dIn5wZvYfcrCvtfJ8x4lmRGiztf
Qx4SkZY21h5KhLiPbUa+yArq1oaXU/igD5oE012lvEWJpudYtn1umYRp5i4ZsVwo
k2baKiUurnpExTQfghzwqsv2kD29A4EwRs5dH84nkKfHUhLUd5nOOhEnbPROmSYF
koFzHD+u+0eF2s+T69v30tAdfm30g65ggc27LHnhn5P+MCMsYjBIvSo2fELTWvhw
GtoIXG4seD2ImctyHbGZYljyH11kTDZ43P5MxO0vUtXZeKidzC7CLhXifKvIrE8A
id6LwBzVij1cvlA9sv5VWOq7dR+3SzI8lRu5lpxMmpLzWN68+/cMieLuEjzFDWUJ
R2e6xsfStEMrHwEQw1hfB5MVNaj9ZKWoeOSy9P8Hj/i3bg6fyZS9IGiLIADT+iLy
OQlzbtU/7bWyfqvMCV2ZPdR5litNxbhHGP2Y7IobPV4rzIeTbB5SZJXAMB8Ip0Yv
pBA3UdDo8Lurq/WVkh/aYTXquiombfo5ANtqJcfYf7p2OLiYuGAD4p/JHFpjgOtj
mVRhsL1oswUJYYQY/watyep8fK/hTsv33yJhnH+gs7KScqZkxQ2ki+xOiIXBtksR
w52wqIIm2AvmtwRNEFSKLHvgRd7qIjt+ZoYq5WE/1Ubk+5Epqh+oml1PFdyCI/IV
aw4TbsgKAMwbzzCcmyO93XHgGTULzqgLkvq+DpVyulJHjIH8PX6yF63XdwdzH1yO
+i6sAnTKPS7ysr7TlkqmjiisDPoj15TtA6Z7g/WFn710BL0NeZITPgksuPXzalPb
SkKWdNE5XCAYdyXx9TtCWy6ZmwUf6pCQNE97kZDuQ6SYA+sC1b0IeeNnAYCFV9+E
40RrihhOyp9ner9j45LTU2gDWB0SY4mSK+EBWYW9+eV0xf0AlnELdN2Fo0HHCK47
IK5rL7BEihPCexvBsa3T1Q4cNOJapD0vKuRYOoNqwH0rEpjcYhA9y4l2aXylPVBH
lO91Yg9AB7cO1mjWL9d+WkkdIFmoSqQqU+FAA09rpkRs/iXAwJxIepksGjsyN81o
zTV0xFTw7o+iM85br638P7rM/FV6Ml21kIG7W1qAb3+7O3OGxwMXJjA0exGgdTpC
OplcmTtoRnXtkIGF1GXVkZthLvv6Vt/qh1NuKacXDiy2G8ecmUGwA0UAU62RtgTs
CpNiWv/bKsvlKSdd/s23MFvML+6DCOaYF8cNxrdVs8iRBEv7xe9v5K5itOScYKQs
yN+FESWeLB4RHmm6v4YTJoIBYtYK7xTrKPcastO7M2i8QSYpTCPzW3cqvCtoIJvR
R62LbGWRLvZxJOt7Aae5Vq6AbfE8Te2znbnn5QHJiTp65Xp79rNP37vCGhW5naMG
ozITMtrfBQufspzfTeqsEzE8wscLnIFAT2UV6pvnBbUvu9Id0BrLBg6MQXX7KP1e
J25Du+srCe7LicjPG3M0wm/HktNIC3NEE1tCpHrM/1IM/uS84n9NV9HdydBVOELO
d81uVIIeUQ1SYEM6jmQylTxEFW77wRTIaN1bgTydCTFjMdt7bvV+TKl6Wv96jCzj
1DgYtgHUb14O/kNxkWk+UTOERlGlU/fzljpWSroGuvzdC/rT0m4cAgVAMAMdlu3Z
D6V4HcK9attupcoPbDdWLFMD6R+u29VH7skf7G8GAgGSLgT6EVAw6kOxJJEdY/8d
FxmncVPNX1cFwTvPFC/q5Wa0lQtV9WAyq5gR37xRMoLLoIRx/QMfGothB2JomQow
8aWcOxax0l6KYsDxzW/XH9erjvalVcKF7VISzE3o7ECb+CrI1Wf8ubjBYc+ffDvk
bMRIu5yQVTsXCY+AhR9S7Md6hynsblat+XY2TnM7zRf+hYi7p7DHy/QXqgxQJrTm
chFa63ITvTBvl+8IuHKYUZ6iPhQv1e3CU2hL0z6k1eu4A3MYjGtl4K5WNl3Uk8rV
kmBVmTmfuTWuTe96n+zAC5eaFMaXWflGS0Xd5xDsO1/e9KKMgDPgTbuS1X0HNN25
//9tktfWgi20E82uXvsQRSntDhQtCtNxWrvn5fNEa+mBY/liLePG9AG1zl8bV6ux
sTQAFWgzgvmJYHGOX3S+zEVoUR2zomS0ry8x/ul4177LDm+H3nHMo2DkLYtXy7+I
wHdAhKNkFxhM3Iue+K6uP6EJcKmhJoV8MCk1qZOvUphR7hfxLaM7Gn5NBSEfrMZL
91CSTNuVko9uBqx2svKYGeGk9tVWVzg6hwR/9mYWBf/Wq6lv5OpHPombNdR2Y8Xw
9ltuor5GNTYSw3kfWxkoc7nQG1C9dQYKcbUnvt1XrJ9SovcJPwGOq+i+jxylzJ1S
bgRQ+4SQO8EXVrdDUu9ODD23g0KElIQyuDtgo0006Mcg9XV0J9HD7K62Bar2O6qY
Sp7RvkWwTL4ieZ2/ozw0ChXtaYfa4ePu4Tzdxg/eiuQbWTykEzQKMy3igWhVJK/6
oSOJZ/lNrjTGxNAMtkG+dW/r99nUpOgA0VAQ3dj383F5HZPuplqQ++ZSUx/5adJj
hHyO5STTwWNfiLtzWPehz4gFf4ZKyrjuYY8XURUKhQcETHOc7qmHPuiw2hheL+Sk
ieOhaR0f584EhQBo+9+yO5yVt/c7w+ZvZvwl0f6a0z15NdYy4IBRKHvWDUoNVo+c
0ESV+eVSW3ky8RHAFrm9WDQ2yIbmd902NQdyBCGxLeHap7dOjrBgc7Sj4tVRnJWt
tvwgdE67oA9Blp58UmWGZcOkRnZjwjGxeMd+2kkg6xvKXB5f77hHUKsQ9UAihKQm
Vee0iujuXIa8FvsHXUMr4u5utoz15w6tB6P6+rsLCFjgIsNYKAB7lj5qGOSAnsko
h/68fS/7QHumG1uwj3v/7b/0n+Ffj94qOuGaOsR8ABo8peH6Z9eQS5ijkK1ASl9/
LsrRU2Jjh4L4jZ5L0KonGxC3O5IEUOZyTGcEPmLiyE/Ij8McdRDCM+IHPM5jQNMq
Mzbp8tD43fEKu/Z5ipTbrQrxTg+dZtfLg8sunKFemCWilbiS6pjAkUJn3EOsdUbp
0tjDSFdmAM8+Dh14Qune6XSkbpBdEIq2/+GaH5v5Hla0hpAK8zpIrfCHgR6eaWRE
CETaHm4eLzS+jhOGV5nzcGRj1lQfzTs4i5UgC2sDYPdlapA8I1/zOPmQeDxImcPO
i67fi3LPLrO20nFnq7Aq3OM0kZ5mRM+eRT2FjNGX6cYX1rjiTYvrWMFioAo1Np6E
SjjoPtljnoiA03xfpD7T5gamBdukt98xj7bnTgZFJiBe4wgPA4czyceNUkokPaSE
75pjg3TKBTMlzO65PPTJ1tptyga9hQMKZU4Pg3Pe2WKt35I2SAR52rCLC++FaVOw
XmQplWRwxG+t20dEyvXobl6e8y4mzMrIqwaeWvBkXec7Hd3guRhcLoLfhDRNe4QZ
lzZp5gQUFOh2C0jlwcpA/6RgUFRxhxO0/kxvAUkvHWpalDyTi7ne02HruGeNn1Oh
FTK18K3UmquExw/kMPQIWUAvvMVv80w++GZ0BfKdwWE7GS4MVZegVYPtb52B6Yz0
Z+p5erpoZjqAPj/Zen6Ii/NzL0fJx/GcmP+R45ha6fk7snx8FdFNhIDBaiDL0wP8
hNMYuU+qQYZi7iEvh0y3r6OmEmxvoA/BodcTM0e9kg2k6L0HhIwD7DsCexLtfB4U
e2w1Amtf4AEAK+ugg9dk0ydUjWB22EH6V00cXPyvGxdtrC0oHEux8Vq+sldMKOQt
56nzqaNbPgTXh1cZSdIuox5xFDfsKsxJomEuMeQspExJfgFgFilqBq5e+GRBBFLT
mbAmNfeyCRRz19sYBjEllYF8yZrUzXILGuuBmW53XW+0su3mxX41EUJ/nJB9Izbd
8OINIf12myYibwRQp/gvhoLrdFmwaFsquXWjfh1heIzg3+3O2CU4DMZtiLlSWgB3
MqDqiAhvTBnqC6YKYDqeasVIB74MdItXuaGC6ultF9tnPDY2E20Ed/EjddzjwsLw
sqfsPiLpdVh/qiwRdK4FaGOn1ADvP/7NKjV+Ry0RGX4nqXt2LdTOSuatyR992NoB
5I4a5x/txWy+d1b6hmf7M1rc8SOzT6AQ7vRBqr2ArMEvcXiphP5hb4kpvZSC0RCj
btW9oymvbp4uQk5BpsrCgb8ivqacR82G6nMczPscHqwKfIgTTXwI2rmJxeDnlbZU
qTtHNOM6QQxTSr7uzLBL4MOQjkto3coA6l+EnXckJpuBrOJrpVKvM0YSu5pq3Ugs
n+ds9WPwC+qtX+mSWJVSyzxFODMgg6y71RsnjYpdwvTeJ5AENW2X5AD4M26a3D3i
29saio9FjRpE9Ie4umv7ccpTBQJT0K1nY3Ezl5KVUVfUt7QjApAa7AKtnm3dcWQ2
Cp5A4z+cDsTJKDTuHUwYsPPUP0/SRyDCzAVARKQS4ocYqH+lvI0GyHopoZd3fXXs
rsO9O8BX+66b9YLlx001980PL+D6A/qohgZS4K+72lJgolDnWGjqnEZL0yemNd9N
zxS9ycHy9gjpzojIAparSijqsv1ROzVJImzDbGw7danNdCeZjCoDak9feoLhJseT
YoQCOQVuasSWp2f8DwB6EEPxznF/S7macL+6SKW5198fvjiYidAJtFt3KmdiImLk
Frhk221brgEDuLqymQhkm0FfqxiE8tMOndGZfXXRMWBiK7/cnlX/yPxuJ3/km1uG
aPxdq9cQkTFNGcGw4OpPq5zPct/SSZBbEsY2uaY4X+wZwsxzpWCqem2fVUNkk4h6
q+icPo3bNum07Dap+GuW5tNXTVvXmjEAa+Jd7mqWC5jrK9rGHFTxxlQdqckder4n
1tuL88qsEn/29QvKgKelbqo6bnqxR3YEL1QSX4EcrmMDArF13HMoJ/dAhQ27C0E4
1/RNXVTybp+S+muWLUEhWW8yAHqeJ6jAf3DVsTAtEhIDaFa1SX6mj4IFdQ1gJwlO
IkmksOjwDQeXEvKaGFchaKFbmW3LbBJ1o5rrQas4Q8YNjOPYNtsQ8sTutmDOhTmC
B/UhChRO2t3/8+DvZia+WisuZYY/FUd+5C/9xgrbXGMlonH16jukQVW1HbA4zudR
1UvgzsDpBW/v7+VUlmLUPpqKVM6CD+WgBJ6QWDe4XmscDGOipE1nwmIsczLg8ftN
p6sS8SmktlRgWdo6GMUbNLjZmjVpy8uenDLsnvEeVSUWJqyAObsclzUDVqhG6rYM
iuVAqQg8oFX984USCZWno+OEoNmbG2D9JYuzMgTYtpa+haEbWgLS2EkESQ8ZU+LO
ahYvhnNCq9suf1OEQRqYe0eL/8Gs3imBpU1/0v0qZdrtDT65aNEdW69Fx3QjsRTW
yjbASau3EUiKOv+BeuhYT/P1fZY+N8DK254bAOv6QquGc9bo8kpMEZ/XnJBYP0Fz
4DLiYsgMk2U/aOOA745TS3nrdQsiNvaNdomjaiUdVZwIaofgIDxb0dbJcnBVgEGD
XNxV5SpgYGL8ij6/wzNzH9dPYoHZSLH4kLCRCRkDl06Glx0Uziq1cmRShOqBSCSr
scSfs/+27ingEzzHimEcBZCgGe2oJKjXd5O77vzYW95xs0weozd/pzhLZ5QDRfRv
WQK1tB6K1Rx7rJRtrw5FrHQ4xnyRvgfKEFe1msXYPbjwOrSN0pP3uZay0G4x6Qzx
7JfCkt8NHnF6T9iffBEY/cV0Wiho3B9c2iQjSwpFMVrAs6nGS/hZsiNqYktAuI/5
SFEoeoa5IpqlNE2UkEbKtHNwbmYMxndTAtFsit5cXV0zJW6tE30Lnho+VqBQVAMA
oFfV0kh++FHd9nEhrYheFJD1L0Uzge+GUpH6+nh6CNwG8qGMHEbFGEG1nbzHylqJ
gxAq7LowYmqckuTCym8g9sdy/9SBh0OB+u90L/SGJVXybDlWJGXnxsVsaKXrjAMe
A8WvmgOX7zsWIPukvAc5Wt9lGxaWkNXe3RJEJMqByYMGgV75dwcp8I1o0O5m9IpI
ATKbs5EHOu8qGsDFmzf+P3BFa5fnN5ty3oN0OcTdV0Z/Qf0BcjcjBIVSqtdgS2QY
qGXarNw1yNZOGHCd71qyk3I6Gvl/lG5S5qjaZrI2RS1wLFLWg8e2kaGntOC1aug3
uh2+42S06uCqdDJeVqCh2cqR8n5IYa4V65QrcX7IOMsWlb86Mz5mt9evn6Ndnxmg
0FB06v/wzNC1GBa2o4VT0wHycTBnRhNtTKzPLN9UDVT5jnIHwrrxQPCdMMmXqX/F
YIU1yc7M/uoPGL+72lpdwCBIw7u+daIa7rPJqlpoAwGFGAOJZgyncbnmSQp23pqz
nmPwzPfGZfaiFoVsra6fb7OCFiI5mNYM497QXj8Bd11kOYK7VtBfuuRTYouMEm4O
pn518ZQ/cCcwcMrhifstEZgQ+TIEiQ0tlsTdFs2ZBy18fSXZ07dBVeXYAUZ9BpoU
iIgdPY/IMmr48eNK6oSf26nk2Dl8OBD2Qfon+SW9kR3GmGwYK7oyTEWo6kTTvF99
zbdaGLOCoXIraDZF9evL7/5swhGzK5MwtN0z95N9fs5zY4Uz7TpO19wYFDyM7T6w
oasSjA75qaxEXPBpAObpkStzN6SD5is+hiGOtpwQ6s4bsIxzp0CwMSs4q5Bh/qd7
Ornh9NAnsU0vDLlBNXoDzYAUzZ9giU0yjeahWHnU4nLg+Exn1k8hzDFUSseMPlnQ
QQatSoNa4iavobE65j2BWBRpRPFc0pgWzxUUzhIcmVcARokOInemKjMZ8oFJKAuS
YcH61TXQaHfz0zEuX6QSt2hDPMHNZXW20WE29QNjHXqJHGZb3uvFreUbX/UoTxbF
ci0uXOb8jW+qXX9/hnAjIFGVLa2KXYT+lYkPfOivsKZGpG+JT/hd4OHJEhSaoFku
BXs7aIiCdJIxqXpDv7K8actSK+t9os5KF2WlW8JXcleVDiK8qi8WNwn4olijBnuQ
5bfiBpwciQO1aHMLEd3YpjabHqYfsrYjnPIVRmY3qHqXbKFox2+qpu0O22uqn9B9
LFeu+8cMWoftpVK/1yyZPzz1oa99z/8DoyEx5jkCVRZ13Z06vTRRQB1kout9Xjm0
8g2WwT2po0L4Ft6jNz85e9v+hkMXCvlX+qNeZ3Qqia4UDs7kBmieVKWT13zqjMqL
ahHzzqrxQF3tj4xc0W44V7LcDMsKbEUfY1ZPIGV+bLHPPxR8FZjLsqcKNRa1TEMI
+XT0eBzRPIdkxYg8is5zwN0OG58+d1ne4fwVq1U6PG0jTHtoYh1ALtLhdZ1ciBI+
Ez7zy8SXN8Hy7bfcss1znkkdbSX+afuoRCW+aaZy93Hb3RRTYVpnSaVE5vvo5E/0
XrJU1gB9qDCU2WRUKYEJLDWNKFdOr140fhPxn2jX/rdPw/mTXSB8JLqjL38R+xMX
WTUDJHWO9pjokrjhU7gby7NunC0hmZuQxKOiRqMPIaQfpPeNRLvp15+/HSWNizHk
zlDJA84oEOdp8Jtsh5Ds5MgJqBzULX+Ma1DdgjCixCxpnfTpL2kQyMi4Tw4l9cxY
YG5B7sCaAs5m/z4hO0OLVMRUqQe3HK0dXF9WwisqxCB2v2zzqtoCu5fgGqqt04Vt
83JXHOrDzM8w6ibTGb/rGDxmnbUua6XxO4CoxXPxEmnJtY9H5rCoqv4WL8PUAG7n
vwl5XzH2/ndqVp0qipzeZ9865zqDtlkVt/CR3d6S7gjuEpvlA86GJABWdZoZz/45
OWHWSU1yVyjjRQ0xocsKrjYz6PYwcyAxjwBCzIYTeO3ruAmya17coPDpyWX1z6zC
M/7iuNx69g7XjB2noKhM1mJ/PmrYtOMXycOChZ4TF1/NF4A115jRReShMxn172Wc
lUPlFOTXXHwFUJ4BA3lxp+mhVmIJAmJF2jAtwZ/C30elcmnnlrhoM1KTsilDlLbx
1I5MnQHddQzU/d5WIb3kBIAwrfOhThvFS60+AXvpOkX4vQHr76NhGNwkPTNlocO8
PbkNrZldBdJU7wGGnF22HqKn+JeZ5qpQA21QZvMRF1x4ZqubobajPUGogxHzdZ2o
0W6ygFkIeClfZ5BowHi6wzYzEhnyiVszBNA2unGKNFm9jJj8CPkN6q8/pJiu3lAS
Aljmbd7DPHeNUgGRGSZdDQl4hfkgzyPUqoTTBuG1kZ13n7cyZGf+uLM8Q2wzswYn
nJRuoNZhHt4l7M60Tb0b6Aagz70L+KCZ2/KtpeLjA/cC8QA62ijeKGoOvkErhrln
g29YHfVJwOzBjkzWJaz2YHRjUYQQvBB+s+QMnZgk8GqUrYSOyyddXuK5rzolD9jn
PPIlxqWRW6WYwdLyjjgwm6oVe2bh3xI11Jn+wis6BMovsqi3ARAV0DXus9hj2G4o
s2Hdm23FJdcK4+JZd8dogQshBBUpWJviOh7JfCGL1I7LEeeuSs48khEbTPKYdoDq
rBiXdnRmNfEGjJiGeJtjGaXHpBhWAWyHqQT1Jj3KpBdTxAADLzkOeZEBLusqUtVx
XegIlwpNr+9pKmbTlRqqwuTNW72rn+LQYGfz17HvS9cmsuBRQkJnMYvm8ImCKDqk
PkepRMZR8UfXV77v7FLMphmHJo7JaARDO41fH2gRAbMnxUp3x1zy3WlYS4lA/VHV
66d3uwgq0IUhHjLjcow3/NFzqSkiulauZKq1chnt2XKTXKly3H5lKb95rlUxmgcf
ZmeRMXQsg5/Td7RL784TUevbAfe59Kxi029tAA6pPZVG2TRjcBijvT7hujzPyea2
kbeT9lwjPTu4Mq+GgWybi2hkbFJAdzVTkK2OSTSqPKhFrGCrUaZV3UdXctSqzFWO
fxmVw27PHYg8G0qKN3XDypseyK2HCslHhgs1OlCXzPLWx+MtCHpus5VKB3iQNIlk
ZPi5nOtqrvqnEqEn0i7sDiFzhJmmXHTpsBn+H04XJkMaJ5us7Yi8E3n6qe8LrV+X
kPWOcSCYXWIbX8Ru5cReXhh1SPTIG/k6LrENOvNpeC7tGDkyihgrarQbInvV1Mud
Uxuj3J6Y2mKrlicdSEjnv2OyflUpYTk8czy7X7mqmsBvpnhg0kPTulni94bLwYSH
AJ9liNmxlq9rU5FHFl28xKGnAg3BqQeYSMUl6BPOXfU+8SSfQyyNnPJjzN/5CfEc
FjZLPbi2iOQKMmCbkRjTA9GbE0Oby4iEkY90eRUQLmFAJWsjiy4nfvTrIdvHu5U+
pbQyYv2nGbPWth5UTw09HeIZ4x147bkgLAb5iHIygnfv6yNY2XOR3sdCUv8B/lNG
AuBaT8zOVdqDhoEmraRd7YpOMP1LajbeVhxK/n6/p7V+ZGc30k6q4LSm7+aGZmGF
uRKtl+AbnHrYWtRjiYHu5Lnln1vyresahbi+ZzoA2kNMFIbLIok/dGSBOvdXQexm
sdskodT5TJ9cZ8jQlmVRk0VEKNotSQoWvy2y/xD0An8B5joCtcRP1cW890+D+ZQc
ul+2S4y0F7K6w+xwGNaHneVJVYpu8Oc21vqyY0EiO4zVIdPQnzSpSShRm/FhjFHb
DauUPqevtYvjiTRCvlJwcU97EN/T4ENri0V9W4OMPUGsKA3vaj0e8g07xiSH/jq+
r5aClJvrrW7MEBntCnOIsGIGCLYHqSkLnPxFs9DPO6LgBQLBo5uIg0WFepJDkWt4
1bJF+9OrUwiFnmWbRUKBt6LHK/0X1XlTeBLD7a50rKYe8yNUSOSzsvpkH371vCsX
bQubjaRtHH0TQfv+MtpO5g7k2S/C5FLBbMWdhGDVgI8fD+lsAj68yGCQKmllJWih
XqQXvFDzaZOgrOLAGeKLKpdAtUC4jC1onLJHisq/UdbA8y4uvsFYZMW7EMxMw8wF
+kwCn75LTgBfKoVc3YQgffEW3niXuAVQqZzJF6OL7qqCkbFaWSA0QFkXRaQCxzxe
P+pePVUp0Rrc1jsoitlCoxlcl3E5SkN+zpFVctsDOz3gN7tENnKAJfBSiXWhj4Nz
//ZQvRoFQkwFpAfLsa8iuAbdY6pjxDW5JjdbZq+tzi/eb2sstrk8lD7MaSn/lT6F
Ze5TQ7hPkUH58fLfT0h8F1sw5xGFGcN4avEdB/shWbvORkJ9BYpWJjeR8zHaXIRq
yWSOTrNId33L468wENkO6D6yZ4YLgng7sw4iMud2JS9QHX1Oh38RTpjTzbW3QOzu
AjfVV4KlO9ID8fimT6MAVSprMrr63UXHrrDla/Q8De0XU3wwYE6DOPCinFgBhdGG
jDscGDAE9pahlIYIqZAJn3aARbBejc2lTVFxR+SluoSAR+2/w5OcvrEgUiyVwSAI
eWSNMsGE7B4zIW7JOAvDxd/Gwz9nuq0gkyp9aD0ajCBKKHEIvclclcCUdhqnlDQ+
Xm+2Cwyv3ldWFO94zdbnqpl82rkceuf/meLq7y0QACTq+vuKXYFOThDYvhlQbFHX
+VtJ2GJRfWbZvFEhYjbRvWgqYVLLXtKE3UIy3c1OBpHMVhVmNV2kC8v4+PLd/bMQ
V1NHwnmTqdZlxifSesqdwumyMQWIDosavkDPYjFaZMEkqKX5JTB/b63xaYvYu3pW
g/GewdU00cMqHH+T06McpMzMsL5tE4TmKp5W51hPJQDeG/QIUhViwrJheRwfFzzm
u2A3b19tAjEkbxX54vk9Z3SB0hiUwqFBqIfK/tLv+Hkv5TuuMZoPALFGXbgEVG8a
K0EqEWt3I3mmrq86akVPpUkEtCjZwgAgNPEHGa2aVsQv7QnVZjG7DJo6FhG4KO/O
SGWn4Ajnhd2IYQH27X8F/UI7ZEoUDYY1V3MxATzBozD6Yy0V33xZNtEJFsJTg9X5
iO3dOfkWO7NN/GnDB6VGfE0R6Sq9zZyBJLvaZkpAJZtAHkoStOjMTtun2yJzHmNA
0egIAstSFKB90fPLJ35daTfs2bvstP8ZFkdqDy8d5IO/knHmm+UOoCq5EGpkoNKk
FpqvvrwYHr9a/PRpQwMng+5ORDC5zc5QfalqXg0dlsRKbFhOu90zs/fy4N1RaXzO
+lzx4LpowtW7vkxhpWCAj4j/pf2JlUJC9UhTclrU/yCF5VJIghexrJ0O2YW7UwaE
AKMJv9YUZ616Np0MzmqHJkNERmUvptKDmw9nk/xjiV2v9AGtMEHRgZ7xkdlshgXM
keyioODtEmNew/+kbri44Keyg88mdmcDYCNnhnp3uSA+OQH1nszQereY3DhW5y5S
zCnPc/8y1mWg/bg9hrZIZPU0bzbxkys1gTzden2W4BqA7HmzeD+qKbN7ry7jzpoc
VoufG/R71KwO2y2Lq6VRi+0Zosl2COIEx62BA69iu2v7/QcrziQhKqKUg05FPxJh
KYZ7HZ0GUKCReeUfgGJyEcC5g6Ldad1UjzlJgQiKQK4rqP8YsVmDTQYSN+lg9ITF
Ujk0tlJn95Z1DpFcQsygC/10iDHxZImOQSzFrob4HZUS6TnUPlNjGSNOxF54DrJd
IXPfzJTYb0yd35/8ChzWKMDOFILuMn6JOJ9MEt6CXZiir74KXN1nqHdMw0V0sLct
ICpv4aduJHcJw5csrslOl81CDKe+yVcullhQDTjJ9xwIJyNand9NTy0AFnno7KyT
LATyqe0CrDlnxI8TD0DEM3RQbgU7Lj8Th4GNQO+WHMpK6M33WFC1utqTSIjWgeoQ
bPSPMuldGWQdwH44yMBsXp9HB4pplOVC+xoSjc7UfNXOCM4BjX9bfzQp54uhOPIN
sgn4Wd5haCOBZ6hYQSvKyNmPNKxj9bv6BTYutSvwhMdC99phEs2kjjhZvENK0oQM
bkz0nsC1jlQWRFhRHmAUsND8iXkRIovolkYtE50Z1TE+PEnfWUOUXettaQH8qwzJ
gkDXie8ZOF1tXh/ts8hz/hrbKVLTTowwew6GfKZobqG8326h3eh4q3+3EWwSfG62
B1QZxEdvo30L7imRh0XnMGQBUW+b5QGt3OYGxHETULz/j92OuSBhhCJKwmRk8gy0
opZ6dXJzUo7yzJE8kFupS6WG5+uYZFGQtQrBIt0bRNT9+xf53FER+bC6+FgMolyB
xuMY1fP8YN55vMXPGh1m/Sh+xKZHeWB23nuOhjSiKdYLgzYITb0bVjydetlgGpQJ
v7FN4LkGVicFJDtC3Rh3ubUNWkeL36q4KtEp/hZXiI845NNYS232i69k4OH7UMSX
d1/W9gWn5u2mioIFY4ZNxiVARHObRDNNFfGVe+LP5Pxk6Uj1NOaY5Nh+XZAYEEc0
QxrtprEat/4mhi8R4U1Ck/x3vzB+AKwpZPtmIWt/OZ3LrJp5oeNCvwDXawV4UFBe
fgId3IVuNcr+4e7R/Hyn98mK579UrRlYpPd+ZhxG91dlyvc8fPvBYWsUY04K0A81
dA0CsfmVe0QpreepLpBby/7j9JzFSvoMeBglNOKR0TFmN0xN1VmF9Y8nSGYzFOld
YQl3UoyEsf5aEMrnrgeEu/DHeIchK83FIcJeJY7a3Q0JUdQwSb0beBaNrjl4gL7W
CVlg15RFx2Gptov3dXZlmN3nxk2wwNrPPlJoW/edzNz0btjn8bQVVBApo351AIxK
rvnCV5oJwZbyYnTN+ad6GvWXOymDT50MfaJf4OfESD2dwOhnHPfRdSN0DXPmBrph
eYC9QYC6QjHXI2lKc1J6ZuqkvswmDmw9aB7CD8mSREhpJM9KZXmNfq3blts4E4E0
AxERm9QeCS8MBcSQeDBrbog9QT3aAgZMR1OnDJ0XXJ8mopiez/fNtrgdv5jvK4FW
Rjd5L8dhSpxwmTz87+8M02vDzW36kOaKzx/fjV9WMwGD+R6bJn1rVarQQ3HLfeDw
fVxq3smaujJblpHkr6ej89Jx6YQ5lOCUgeLwSjrecmgtSFiUUyYW+e4dJ1rRa1AZ
vCXRWxeFBRHDf0hn5Mro2Q8yGLSw17jpocbC/0EBm7sZx+/XdYDnZTAFMi5/oq/W
weyiPLUYRbbDZ/be+8Fx4Q40HRm54cR3bENKn4p4o7r2CFYAHf2c5TRzgd2mPUTJ
iUsktfnnrgtljLbGq9eZxi9aAeDBkqZOxFk69isJzs+cn9WMtpvFdIOLBkrW5JJ/
XcRRyE2cgXJalRcZ/lFRTpm2z589BXI1gKwH7ay3Oh0+kP/f7B8o3wkkc4v4aOUy
AV0COneLVOSIV9ecypSIeB2VYafMVXN5ZSRZiDtUCNYsjvnSP2+VBnrG/UAmDeb3
uWkCq3eufHH0v2Gnz49F4V595h8x1cOKv5Y42V9XrTOwtpYAUJbPUQCPwsaPNmct
WR3JG3EjQd4pkZbBYiMQsyP9n87la9FcFDfUl9Pv/amZXd8Ti1wyaDJE1hLLh+Aa
TRaN4o2ct3+4Elpau+G9iJjcD7pNKr+uOpjTGRXmzRtxXwA/GtvJJxPUif+Gu1MA
nqUo7Fz/BYloi00OE38tdlQvvX96cys/S11PCiSYDj1Qoh3NI7cf3uCxX6Ff7R78
J4rHDarS7lUEsF6l/O7zIcDL8JnbcGPP8Qqvb9vYoC2Dzkd3Iz10mcHeLrGMWSKI
25/5KiEUTAGx5KhF1BtXKROo4zTBMtfzzY79cb+FKBjxKSjXRyfpdiWTlPnbYwEl
xsjsyxm/Y/Ufv4qxMAj40psODG/SQnoeommRJjOgHb6ZxDmCO3LXQVk6vg+2EIqx
Kvkq4uvHCiMcj7qiqeNLj6oyqK3VkkyjogVZ8oAB5jCUkQWlFCrk3aKXS/wpBiUc
8BWOb+/rK5Hx+/41LYQscdCSxAlczkK9CN1zhxN2SGa5hwANU898jyqJDjjLhHd0
c1GgcIB9DCpyWDopbSY4Q06MXFmeibDQVIGxtxIF69YnzoQr5KCn2aFFm7OI56Ec
VHz8OAZt0Z3Yh3ChQx1xU9/MConnaZkGM5fuPnTqNt5ejwh3AegJa3FpDpdG6rNQ
4Cezm9RLxo1cADMLrY9DRPrttqBsoS5Ir69NK4B/hIPrTgThE06THchY+/KsWmDP
iwVIQpeJ+UOx8L4B1hAxoGzbN8mQMkj4WciSpNgczlTJlr+LLo3JUW+Qh5XMpUMx
5VmZoqdHOZBjq2yMhreK3Hn8LRhzdJYNAGqycSODWZx1n/hxwAQ2eKDeuqs5svzA
ghdAkHv5KfDQdyjcpkiTtAiQi1/ddSfiiQoPf2LtJLgKc+Sw+k2wcWBGnr5q15w2
13vzDh+1XNN8a6GdIq/aV0424xWzP/zGDHPp8+LTf1lN9Y/thQXJBNbcvfNZqXfg
BDjazTnVbTo3WUxKIqnnM9+IiDPeNkeQmeQ+0MNZHuWU2HXzghMVe8IysbOiqaqJ
/RRyVBTLzej3c7wAtYk5etyEypWfUTXp2ULxU5m/rcq5xYpeIp8zrj2KJ9dRP9fB
PINRrMc/fQt2GAx6mVolaMZ5zkDfW1o3C8wEcoLqTN8x6QjDTl14gxv/G8HKgZ5f
jHuPp42jq8qAb1jordjUXdyFgJh9d1Fj6+R/wRjrFMOY3NEzGtizpm6cMrS1gcXq
ambWvNE93B3/ft0rF9jcCOTg+llqW3tFmmJ5/dDFpxPMDaO1J0CrAonkJ1U44N3H
fDc8adRp8Z+gtkj6ZnAd1h3TpVNQG3wzAQyC0R0M2tkevzRd8prXPZZvaZ/u3DMb
eSyY/xWPjlT5Qps4lYNaIVE53uHfE2Gyerv9JReZmBBZf1NHdIm7DHi3qcSUPQjq
9B/J/woVEg9h5Pq635rNGcy4vNSTGPtV1V+euQdgIbPYAr+/f8sGor58250nQHWa
iu1DEYEfJDP+gkD4UuddErkrFhA1WXJlIwaw0Q2PTmouJ/0Fr1bBkF2MInDXhVgv
pcRMbNna/Nh+k18463OcKDrak/IF/AKIWOswjIAc87UTQFR46IFic6Tejk9sNeHT
lZ9IR3tJyEy9H/6iXddfqavxD10zvXdR9Wv+dU8Lw2U4aETLYMjBUbso/zZ5d4nr
880Y3xTXJBBG8M8PNKN2NtK2ae3tu1rKCIDCudcIcyRWnIIUliIVHW6/TQlDY28W
/G+RwL2pAnLi0yRncRa464wVTKNHnMO1FKGuV+h5x1C00CWDxnLesFSIuVAH7vWN
Rqf+sAflYu7Rm9cUTaffNhlYIXvun+lQjOb1nxxkE/KZ5XWZRC+PqN1SOOU8kBco
Mj1n17JKibJ0XcVTn0e8CfI9oOxf7agWYiVCirkmL8VgwBo3fPZimAHCLIqn193o
QDGY3D7fXOeMmNxL4fr3CF42QRR0IThRupBR5rs0/1PvtoEhGfyVElUWSQPki1/T
XQ6C5YHTRtU0BNY9LcOll1vCO7dlQpuwbjqLlzTHA5b1aFfbQaZ8uJG4GKGlHx7D
e4k2xL1Ne/MHt0l3nhXlsI9/cvVpjk/pqD++8/LG3J70ccaS2KSHfChYF7PweWt0
47ckClb1RuYIQCZtTaTUL907pkq+kFnaCW77tLhySW2zVpkIGmrvKGNoGuygSjk+
+9InogGepjFsTAEwiYiGbwSJG4KW03VuQPb0viwemPu1ufveaSD7FT2Gkt6EY/fI
c62wzALnFfurUM/nvfGBqOKeDgLuyjlDLrPL9MYJPHpVvmb8cbvsJ65PxLPzcWq6
9ddSglHwlAm7rhKMWpdsL4E9aXWTo3PzcvyyotDLr7cRHuQIzCmBsRf/9oL/PbXI
sQ3itNGEbO/Fv5Jx3siI97W5DuXuDpLgymWsk5BzwbjDrbN4J99FxUbc9sfDhJqj
MjpCKTHmh+RTpgcJns1bEIMSyZb0Zwpm0KSwusc/EPvC6qXCehtDJJmj/PMSaoUs
Ea8ghr5IwjjZXgxekS6OsEYBfzj9muV7lK3vRKyAsqA7MHeFYhR7Xi2xfotjjUvj
HT6/eq7vaiNhOs0saG7GTX7SyLP08NuIcQX4CI3Flny8BsymLpaa59bdwPej5BjU
KB5IVo97meTMltYWMxaDKTnquwEBRgg0bBFuQTwwJvCetHOEIG6F7dTrZkelmLQa
OYyvbSkW3He8/KDmzqnphgvxUm6nh97+HLH+Lnk2ZlqCSFYNR9D4gurijZK6eTKe
Tl1LpJpWzyrnqj5pjkOMrEJ6v9XA3LfHmaS+tlYxTpNs0vP1+G0kulY8EeRiPQ3F
ILXcGCLWJqywlS0O0P5XTyR/5CHHjxANUPefz1MVbttJ5p5VT1iImvGrK8m9rODD
WkuzA9Cst8nEUR++lWZyjV5O5lYZ7lO0n/YXpRS62E1alfQxD5BUYZpeE64zRvSO
uT4JLKkXZnmcHsy49GHSDK5DbZuK32stdeSTzYJLjnzrAGCL/H9/X51Fh3H7ErON
fhnfv75DqY0QrQrj/G+Yn0wArgKoKLmJjB2GaHfTZg8e1kd6UOXs74hOJQ9MkHdl
o4ixbdY0mbaLZCUXQa9Ja8vQvK54I3j5SWId1Xtm03AbzQBSocHyT+FAUsf5mMEu
eesLoNd2R7mbtobY8O8CsvkpWyHA4fv5daZr4Fd8Hyqt1PRw9nc9OxscrHyJvlbq
6j/82D82ddiHbEtFPQH9fdcd14vskbHZAVYAVNtiDR+v0ZT1d1iMtjoS1qBqhjLe
Zyi/w4w+0O8trrOHyuKBl/BNo1jPwGorHhSkoRmlrQx2F8IM4FtcPXUdJLI0i31B
6Z1ClN7y3eVgaQtwANCwYFbPaXPFPLgTjqgzIaDQwuR2ecX1+/Qb9CqnR8nvIssg
a3cIO8ks4A+juuuLzfMsrjeZCNBARUCh49UOc7wblu8oE2BLXAYmjG0ahz/Gxkwh
5sEX+U/XlvfrS43k8tmsb2KEEwyidJdClOfrbE5NGRjHJfAjOI+/f5TrjMoe1ipk
e+tqXiqw3fWhCYCU+6T9UQjUDmGqeE982QA9IwXDO4UH+aI+TjjrA/tWH4rHAQO6
x70hjqelQBtEgaNPV4R3EzDqKd2NHVJU0mcKrQFw2xPzAqHNXn0D1DOePOwb8eHw
fJDfyEaX24w7vnEJpycRIz7KStujt1+nSHhGTuxbQ7RdkjBD1BZZ+wQHSDNcDN7f
5/5nh+gAG5R2+9mBBM0iNOKhZH+pkh1z2B62lsRt9/M053EUpgs0qiukOnHxQvsT
0lEPDTdMTwvprlNlfsAsZlIuDachWXos4BC/vYGhI4VbT26gYV6RDNDGgqnsG580
VgdSkrCHIFmmq2Aw8ClUR0zAh3JzoeP7ieAbosCZXNX2R/D8KdHtds06VxQkFtxo
V9Kf2UE+c8lFWUy6DeH7TJHzIRB3hZKwW6nZgKUwqwJ85WYvPD7NO9/S/tgrydr1
w3Z2bE/kiu2aPjnTWStkaSYOBnbF4uI4V0ZWQp0r/GRpymCg5jFV1o4d9r2hFOvN
gBpTy0Tnv9qMYXG0Zo1Q04oL9nghmW0OyRGlmvklPTmn4ZE3rTYRVOPsJ4FHm7YP
gr33gJdF3N/VpU3ERazizLYnNFZctqXlL+QD2F9ky05DaTiLExd4AxFwYjuS0T/Z
niNWnQU7wgp/XR3RvOj/VDE4Gl1RwfosnasU1tTGElE3Eg4jMpb8yE9IGv/S3zVU
vKOLvWATjeuNFaDuAHVG2qx9NCxwAl+qUtrywyeLbvxXsOdmuxvFsRfg7+7CQjEf
Vx/OOOxof1pqxIKRwh2MGG7b0gTgIMvsFF9Wi/p27iJv366uDrEJEgDWultXCU6E
N9ZMiRAXorbADNTxJf3wQAjNRMB1b8AUYTiTvWDs1TSeAuuCskug67vcshzOLD/h
q7fSMpER2dYoNNg0MyxqlpmSufSjmWvVFNMWT486ssnbtpGcOnkIGNYX+cYyOWqy
0ym7/5f58DUAWKBjPjEnrzzmTHV9jAiIEqDKPPO/SVLMiTKthMQOI/oZ2p60cAF1
ltr8wFCRUy1QRMNpfWhp/0/P4sKAlNKQps+HaV4cRPlR0k8/FY3sKXYjs9+RVtkC
j2KVorUFOSOZ28W7QAhSRB9v1xiCG7ju2yBiSPO6uxw7nb/vO7dPPrFZUwm9KTUF
JLlreCJNX8amwVn7FIun7p20IKIDKSekJkJGRTMmLfZUcy1exz3uLZnNKpGgo6Dx
Ci2LAKqZbgZfxHdZ6i5M1ZxwUCe+IlL4tSR3qAa6OwO0dbMTQoqHTcc7gx3Jy3vS
y9N29QG/7Utnt2CQY8lzXjHxE0rlO++E/HJPXxQnv/9VkkCuAYPZ9ZP2xDtn73Aj
MVB0pOD7Hs+kR/DwnwZcoYRILcGo3GKBRfu2RHG3hiUdx7AIbIylZRP9Q1LBF1/o
puS0qX2GhxAVaKQCxqZTZO4L/0TUXyRtPRMI7mbiO1e1+Ah0XtgXTVrbCCClboFp
0DhKKRLShQ1DTBxZFSH8K+ts6Ztvsg2WkGUPrzpDNVf8fUD8Ej1Zcj5lrKOrCzFH
TnpxP/jKIdGQCXKVBoGQZFeb47b+qrfX6JTEUH+/UsmbscVwYvpb1t4WZbY10Alh
RSKisH+dq8+cdbMnp9tG1fRsVSJoM8gdiSJcHm/8dCYrcizhn5Xt3qwXLr4DoBuV
5lf2GH50PApQ556zXOIlwLCF6WziXs2IeIhA24qIOxeewpaLLiFhf+dn3eLH/8sp
TxUtlCm5Y9GCl3c85alEQ1IZMQyww/EkG9n0uYMWRo1srNkpUwtY2o77vR5JxDMo
2XpF3psvJGZY0QuDuPiDjcIocycy+4Hx7+e3YY6fXWvr+pE5mg/GT+nphTkibVaj
WBn2W/pc1XRpFBlSd1PGBkq1TVqNVuEl554rq7Q151ilJzyRnokpTtIYpjulB40Z
CNuE9nwGGTll4uBHar5GCUaCuupfaU9tFGUXr3hwkuhDE194rvfBWMkR8Pcd8Sy6
lGQ+5tKtsAY7P384U6qCc063q2rY3+dqbGLdPZJvI8XGWREDNz2/eWITwGiWKfv7
3ozmYq6Y53jNoxGNNUpD3dDaUTF26hs5d6+560w6wHTJdECcsiICjvbsx9PT3A/y
pp7G1GlWkxxrEuCMjL67vYj3wfwDVouFD8BKiNuievasQTcbSwl3d4trfRU2w7qL
USBkI7o9SYKCqRPB3xqvH3FXctBIWIaZybm5AllljpPKbQl4THZTpIjXztMn5I7v
zu/jqxd8nvHBSz0eIadV3g8V3+XwQIZy8S0d+/9kiqcnZMkONmazuG30YiMaBeZn
0yCYYk4iIn6RFtwpvuUyJIF4+fq4Eo8qgtsQu1SYcpd6IN3/BNi6efXfvAfboES3
Uw23VDgowsXNqVXJVZJW9SMZClIaJVfKVvk1Xd/kFUvUQWE6OrIK4Gov5Y5eMU8T
N2q6tsTWDqaxDijwIWNFNPlWUJA9jCLO15p3Bw7DYbg9Geonyozwrr7h+KsQ2aYU
uQvj1AT+qne7q6vjfoJJIJUXvgosXYS04RHWgFjpaSnA692WJbZbjwOaU4BYoxmT
mZaFUN5fUFtzJabyMqmYrKnuI04rLzBK1XB9iwa1icOVnqI297IVC8sVYtFb6uU2
b0lS+YXNi0nhfgFA9TeH391/PtCsmRTU79fHqtGVsbOfqw2MdrZ9JhkPSatVR4sG
m0ZO6FVdmUWutd9haaqh2U2PX74bPuah4EAKBUqsMcLM0XubdH6VaB+qXKyEZLsb
/UllPfhG7PiFrw/uK+Mi/+zRl1ONEiDwI0pLYnKxHfHLhwHXytR8srNOK/3pLg6C
RnbbTW0ubVi6mkkbZjBwaHBKvlMa7OxmkCuqCU+l0EQKxkJlrZBweBqTABheSf8d
o+YHHH5PHFgMoDgpxymGpMGSIQzHk2oM7AwyoNunmIZImbYwI1SGe83w+BfY1lm2
7Y39y17dxMJyHeJmoD2ayurgWUZEwl8IJnybi54zCxTSJsrQV4ZjxiI8ZKxXxrk8
Br+k38aINzh8mVsRzN/lqfgBMw89XVpTMAmpuy4qOP82ODaXhUacjgmfyjoiecP/
yWZGbSQnnYdBytRL6BQrLEe1bna91Y5mBg/QCg/1kf+mNxaVwxinMcM0UUObRs+L
N47yoiQVT4yaRp8ra4tY+8tS3Og+djyI02ttAehrOFIIp5iC3JcX9fKMv0bGGy7l
fBqoHmJGCCAi37heRPtUmVQoBIVwhC7MCS+FIe1ZoyK2p6dsUe/SzyJry5DLMjOV
YCBErso3aJsOKLoX1rWLN9MxdKeRhWXrrEILQxfS8qEkJPCvQRj4sGjCruynHd2y
qccxfikooF6B51FyY4N81gZYe2vZbFKw6FseUfA2670D7ogmG8PNV1oR5/cGGxB7
gc9067PJiC6vmTTt95sjde5uuIUws+fTjUADqmBdCz4D5+ZdhY7XTDHj3tP0MM+d
K7QqCjkdzDextlN96ZJ3tT52a7LWHXvgjlczv4dSHoIwOfCQZSP7lJgbQ1ikOkT+
yAM9dSAPzAdM3UHemaj4tVly/mn+Ji6LBxV/jhpMHECvx1oKWa88l5uL7NhjYwUj
urXjW2YTIiAXjk1VRH3ZxIrymjDDO0XCL2FOl7SzzDakKqI7K7EEO1Z8Ddi47A6+
T07gQbuJB31QgEgOZVeVi7O5K/jgN+KcThsUvjSYGhYUrnFdePwWsddnc1VDMTko
rE7ZhM1YzRwYFWjBj8Mfx+cj8mLBmkmE3LgT7d7L5ie9nLpzgSycUNKBgKlkNRDl
wOVoz1ibTweWLm9ZD82vl71ly/Egtwwmd6VrmlO4TY9eYUGjZ7ktij7h8zT1lMHk
IW8bWEOcWvq2ejEArgLlT1NebUP9OunCb7zvb/Ctu9WrfwnG14/pEBUALdHO2CXo
4VJD8GDdyp6fcG10zekbXiM0n/VOs12z6dRXYHiMGYjXg6tjdmit/21iQZUTttck
BVBZejhH8M4ITmLeny7x0VZicmjEa3kYxgafNtKPN1uIMBy++gyxljcVLIGW1pjI
RBlIWi8xkJtTdLUZc3k4ZWPD+xW/yjnQ2T/w5vJkCRDtVo5p12aGqLEDXAFwbspD
F8q3wGyXQkbMlNw6f7Ghl7KHC6MpWsnWzVMp7JJffB2hs5XkUS1PEhBB4N6toyT+
3feHl4p9MA1ZhIcTFw50MY6ZUUYAFHTqAnITwx5jh0KJqqYT4lint7Az4Z8BxCd/
QKr1wIv7SLHjql4YacbGLUv/rbOkZPsVBPOK7Td+LSprqksM5v6ypR3+oxOBbhLD
Xjuwi8jgXGq9TpDv2k3BiQnuceWuEVQBW3RdjI/GX23NbK1oiLUu53GqT/rCdy8V
qixz4rswiARP5kMTfF9bgfUrraaFJc5pqkZGgQSwTdoVXOexSvh1LH5wWKiZraUt
GLvs/Gq37MqNZWshV0pzrrzrpnfzfaqznroXIAgNWGiIGc+9aoRH8/V90kCXVR+s
5vDA55aM0nnxIc7zQJKau/XvUtC2kVTV2yKSoexY0GiEUcpFTH6LLC+KgbzeF2WT
1Y9f+ZfWQsI6KvtC015daRnMTrSRhXLs0d7brG+eigdyj+aXUSypy2/a+helpm2l
83KoQg7O9uyY642PO0nkdKGX3r/ZwX1SHYHZ543rOk5R2Y48e9Gh/nJgt67cptIp
KE5aujgsxF5KCgsVWvZsha6nXb7a8LVjzmmslcgyxJESBo3k0s/Nb1tdvjnM3GGC
OabseIu1e0EfC9nBsjTtaOYgtLZ6blc89H2sGKGEqr0pweaX3rajrf/Z6cuE43NO
R2uedJDp+d4jc0ijVJuMhJMQiwohxNmOaLYzQ7ttGCOJTnzJ5mkjs/Pf2HUCYTM0
+dV02i6xcqkCRvB/WmqeHGcVU9jk+SONKUkUKz/ooPLVLG1gbKPmoIIrmQo8i2JZ
DeQ0or5GuRaRVsdNoZoIGJcNcCe6s3LCqpWdHZhXc9Pdc9tZ0f5Hy0Elua+o5Yer
mcu67FeJsVSCREQ2eH+V7YoC2mUyb0fEtANWcY0hpPLVgB+JI2qFJiXcjUOAH2nL
pKCXWLqrCHIWzNl2w/YK9jodCHOjA4iZiHFCciU7zX4/DFwf/M1qt1UOrB7js6I2
xb5oy/SmBU2Adbs5eQlK4ZtR/ncl9ZEoS3jrxBcbpNj+duPYS/jP1D9FOyFUh0C6
I8dj5EsBN78B4dYTmR2/+Yhm+Req3K2N7gbeUzwG+3oRtrWq6l6+hrGOSIfczV9L
S7y2NoGRXMsKN8+SDAvDRbUuEOZ164xHUD+t8mCeS0KDX2U5ilps6683ZDRjG78N
hRCkFuOmwsIPqfP0zDNUqqGR4j5z8OqzLBw8Ap+fmLfKW42lJvhg1UZjv/HN1iNJ
s00dbNrgIWV7mgX4z8udnblk9ShnvESRryB39qm9SmImhT/qqWmKQOUHhQd3/NHD
d0bxdhrO8NCOf2dnyKxMJDmbBjyxmHL3ItP0pOV+mypdbcPlwnR7jM+WIfZFgc5X
O5rbh8DAjPlZgZ5hCnG7iLUA6BGPsmf+iZt58PD3kuOh5EuY76s0tVbsCCiP9XKM
zKpU9GeKydCFROyIQRCxOHpnVVYvRVBFsIBrRHw9IIg8H0BuMzIxc0Cy8FiqqIEN
6P+Rsjkg0NWmg73BQrUOab8OuCEeqF/zYSertcksYuNn4FTuZKgdQL89Ijll1ptZ
53WBAXObtYQN0ebL3+xRP1+KiVT9MZhOXp8BNGH016TVq8FEo312XYxqdvsZGvKH
RBXtfbr0973Jq1iQDiseqgErK9EI283+SW+zYrn5obAIq+qIZnIwWjX50O56O5/F
SLDJO70jPad3QioATwM3IXWXYTf78e2l+DPbizFVQIxJ3kpYHPzMCeNEUFlb1Vz/
4EUCZVGpNyh43hGHZ9jFAySvMdeIqI8PFSOyuJ1yczxFJAK7ay4yl5elRlszSGHf
1rT8dxPBlXAAEFoPd9F53Guy3bGegyxZsgwGYTNuMaCnY0mVQcIT2UGCo7nds2qk
dnAt5eyKVrIxlwQulnc+ajxsb2cQl8ysYaJs3r6XBm3AniziUhIWfQ8jIAfLWkkD
JJQwtqgsdLmOWVzF69/zrLzOXsuA8elyfFrRNI+AtK/zzl8ScoPjfV2vfqmCAiUs
BtyvlH5Kb+GILoK3Y7Eu7/32ZVqdJqRTjdO/iNcR+PtB3z0CPPJhFV5REjID1/6N
PY57+fa4FARgWiyfzggZ76q6WloGTDPqcZiKJ5spKGfzfhDLcbD4BL6PT8GsyqPn
mf/DREuLjpwEp2Urmss4/vffbNVJKsEQK634cU92Zt/4Ndr8DLscWXUO9YN4Re5M
NaRHDA1FrmC9NhuiGTuAZFcE1dtVqGujQ8juvv5OWAiH6uvn/ZXJDh/lr0/wIC8P
A34231h97qdX0lZ5jAdP6pevHoI4gv99htG3z9wPx4vH0Q42kgv8jnHS9R2NtsEf
enOnUPaAIIOFPzt40BTzC/obtRyxsBzffTTS4Zvjsoi9CrcFW9+GRoz7QueVJ8sV
gz/Htpk5NJnN0NVDGCSpRTC5W9WxeXBWyIwDE8HJEor5QrCw6GQQipWoxVrYFNGR
Djbr1J3fgzm/9nQGCtLr4BKSGqSJ1eM84vOCPQt9ToQjd/i8oubfXoRURmKdCXM7
l58zqim+OB1iW/X6pMlkKKBtcHax8NFWi6+FWaeUjCVDf7oH4+wuPa09tzOVeG6C
mU+v86UW8OFqyy4Df9bQVXthQ4q8TRgh2oXbqMnMC9JTxiGg9Ng5tyODJKC630xh
RU4FhHp5lbf/WNEBjhiyQy2ODmAHwfn5r5YDxCx9i+soSVj3lzj11odDuascQWwF
6vzvX6J48q8Eh/58TPI0rd4QMYaFcQ3comZ+tQZ9oUuKB0tFKwOWsnQXY2RKwwzW
AlTQXVEmZx8VoWhpfpWEaC7IYSEJ50yl7DTGCSGbhfgb5ATGjS4lLva8b/AvJy36
zq9PSVgotq4rGXHzuWN2GJB7QtfnWtYBAKTBxFyNgj+0nBcxMh+yS/b1/oYdTL8r
sGIfptBl9Eti+0PRT4viCUcmojympZc8T0sjTualllU=
`protect END_PROTECTED
