`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nrAyXL7EXIstylOrjpaQ2KAHmXeNc3vGzqPtzCvVqii3CfTkYnCf5Nz1t5PIo2F/
YS72Ofv5y+pko0LDo8U5+BBqnyp9618HHgygjApdJzo8lKJ4C9retbZgku5NLHog
/BWbv2cYp6baKm94aOkH/LrB/4oPvctzsRBKJbu8TQYkCh5BXosn2Zj2rmvOhIa5
Eu8OeUZI0M6W2BBzb76MH9P1X6GllMiDEjxFDBsxY2JHY3H3c+m2uYnkqJKgWd/Q
2R2fzyDUwKUU9SZ7yxrovP9CIUa8gg1qTLdHzMvT2HweT2pXuZFSfLdywW4TOwaE
BMQPYX2j019PR3SIgmow4e3FHNGwaVnEUYWfCCIhIECgU21KXZCf3yPC7dqQyh8t
J/ccsXx4cOIfIJulMf4w/VuA2qKKXRccXvNvc1nwRoYuMYo8rCNJFKorADOzHcEu
FXSKfoq6VZLTlR6l7UDAK1FPdCfq/V975F4dxCwPv4F6oTAqE52s460P3oud637+
TauL0YoMs/XHX7EjMKlUqIkEiMyOz85uf3osCJ4f6XQYChgEfVSMxJecC2XLc5zJ
6b2Zfmj/TFhWTKfjMQ/zey7CVnpaK88ZTK6M6zt6kk3y2QpG/MXhabaBdeNWVbpx
9bmG5QHLav759oFPpcmtM4Ej5aAs2Nlr9YbJnOZXu9m7KBF3doeBBIvEMD89Gl44
sRbsdXfiJS+6ffeXq0/uHexwunQtevtJG//Pml5wG84/79Hd0FmwEC53lPxaU7Bg
`protect END_PROTECTED
