`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+iJgMjXl/ujqDuDBRxcAqr427l2L7/QyGX80xk9kRXlgxOKjvCupVdkIGi6LlFzS
AOWMVUMiyxkRJuH1uTGbu2eeaLDUxIvoTXH2rYW+g0V5jiCuaMAtwV+s/aCMz9/I
jj/xkzCh3y0LXWCo7rELKyGr6Ksw04NkccEs1XG+8Le8DnlduTRezL7eKpg8DuSI
nhT4Uk3It50MEzjWp1CeB8py9apGLkc4oWiNDt+ZyOwK/sPL1RJcy8ibf85++hnm
VsJFzn3aGnq2osPR3E1bL1k+BG3KV9Prw3OxPRlwPUgsV7cuJ0JiHn9Uke53f7KT
5axXGPFvharklCxWGDFQ9okLl08R601qzIVg0KeqBctqy2Udwf8nnP9xcF2fmiXl
aXYLLMNQpDk/mn4PnL5lsKDaRlRUGXSxOxdA7wcTCCaYSnTn/wSuqe8SNmzDlbkl
PnWOzHnv3XqBki3YVZDbVJ4l/EGACIIIoAj6tG9AUQiRA2LWdtMUU0nXJmWaqQrJ
s2FXN94YLiGEd/Bqz6ABlH41c31m2DOdWt0HfTjfnTOEyqkcJwUqBhR/3uz96i2e
jHaiFzBYF9x24ldKMrYxTxDhNqAmCETeqNxg5O62kGz/XmyU28ZjRnPxcXZLa4zT
v4TkPU6NU6HPfpILv9K4ZLnCeLG6h5jiHL1AV2HZpRO7COMiYqpWqYbi8yCzUPQN
+pfLrnvo+ERXBh6IbpQALaarPoI90pdCJVgWqGHgclK6u5YJm9iO3QpPwKsCoYft
qpc/XizVcSnLZfgLJNSaI0sL3BM3uo5ZvViEzr0nEc3x116eHSavHDxEFiL4wmZ3
CxMEpdQcyyPPtvRnXjrqceGm0cOk4Lq0U915iVATHscKSv6xJ5QzGyG3JsQo1CqT
fmob86YXVGELNdLiWd0PmFt+dfVtsLRVZ/dPpeOv030NkQM3x77woPULZgGxH7Hs
swSctK3AK6thjbZT6ny6IOEeUchnxSyyu4plkYlaroLaWJHp6Anq4L5uNiotAxbz
qvCyCR8SLvRf1/t63dQGTF9JUOHAseHovS17ar1nV1tL4gZ0HG/68vMqqp5KnoRZ
pMYXg1+brZbcIqsfe08OL/fViGY5o3S94BUWfonmf7ImNFoFajb0EV6gF08iGZD+
CJwb5uYQvv8lK1KE15KHBf3ICSlPZUKuuE6OaFTdBKnb4c9TXrqmpUgTNOXGCFNq
B/w7brx3fXPOCcP1Nf2uqDKWgEfEuY8vsOpg7Pn8/4aSKZFQl7KhFHs4h5Bq4U6V
7D3vHavC7HHMwkjJ2WPHYi1e8abaqHwl6eDtWNdKLx0yOFJHiVM97REP11K6dMqu
4kSjPxJn4SOlh88SUoX8CniwdXaaB/F4RLtDoeTAQZPWDej5HEg8ABRs/lfhYokQ
cxmZty97qNRCz+5buKKJilQIxpdB/sZjzUlETIZVB8HNZWKxT+11ILk/zHMvJcyz
DcgSezEXDqXEt6c3d1yFqRn2jlqy7uHbZ0nJFa+zUV8CHQHTDPhFZDjrXz7+GwRq
ps5cBxTdW3XwFjcgpTKBWW01k3LNLCRSXIh9/B7eCHco7QlppGQjXxAC/vM2oJKG
U17i+J4GnqbCVdv0I57D2icqAbweoAmtwBLi59HixJZKX+emEH6F842B7bK1YbML
uXlpGD+BfJlbGlnsXTEBl7FCt1zjWFtqyO6G3x6TlABdEzVOnyV8dbSfQx77shF3
tTJhE6vJMIM3TcbelulaC30lkc600ainhw9PHTOfhsETRx+vUbJFfQAsEIlf+PHv
HUtaUpoOGjzCGZq3WTSJzfnhVaqGNU/2mpwnGwQYWQEI8QHt5tkmcyQVWJAV4ogg
uRRIznS1Uf0ZCDZjDGHQUWdD2Z9wSMJOyX9WQau+rx7c4JWwCUYbcKQfDxXaiZx8
2egQv1RamEIJwKFXznkLfYK9vdNQoY5Cv+mEZ93dqIe7rt0CCRWBwr0dYUAs9zDn
zWU+4hGyf4Q+gUJpF1DIlrX6Y18/opEJboRl7uDKrGlr/9FAFdJUNmlVRVgBpR9d
MUKPBiXUllDN9TGq5bnMkieZyYuA1/vbyPImeXxXSj8lUz2lNGpyijc3CCEs7YKx
vNCSaZPJkzrabHmmbuOC01pPPXZLNz1XlBqpN4u3kboA7ExeKeBi+3zNmoE+5rO2
XB+X5Whb7QEEEng/Ud3EWxFEGQ6aZdAGbccEJfBX2Vo8wNNwWZ92pq8sXX6CPh2y
v5p9Ia1p3ABJAb30itWj34Q+jtIF1OX8VxH7ukh0npGUDtFLEs64BcC7xr1GfhXF
kO7Bsq6CjIO4u1M41N9AIScBGMwhqdjZDvphRQNA+gyZV/Qyk60td4zSsXuRdpks
MzrAO+BQU3kblW8bNxOvHPtdDFk+4C1Da4KkkrGBFDm/nS0sc6+vrzRe0xGav7tW
IMSuvndqIVifHLIqFO9tKKTXGmCrvYzpPzI9tylj4oCNY7txwL9T8FLgfkyDUkjq
Bd9l3ngzltJcS0QdYnyuV8lRaeEE+Dho0OU8jccQuW3hKme/9CoiEl2mn6hqAUy+
`protect END_PROTECTED
