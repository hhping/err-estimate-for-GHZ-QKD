`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ivzdLNpIwcdJJBRJ5lPEqqtPD1rc4cNb+yYSPlL7tvQ6so16yyV5n6yp5Zh3Icgz
UdeohQCfCNBOzyw+1nWI6uSwFvUcHs36qOeRp1r5cIsb8IBc1eHK+dNtGNsCfNMm
dMEIEyTHz6dAm6hFNO3wVNXarfIZrPMg7yLWc6QE7l63B9khUC1ULJhQR66Xuvpt
HdaZXgP2Vjj0OySCep2Syh+8rZC/3gVQxKIY0UDzXX4hy4U98v6m5bXYUH+hSUgW
LoW1zN+cyj3ELSBrkXDDfrYx+IOeFDV5vJ5wRINcLY4lBiC7BMicER5EGsGKgWbj
OrOigNak8aW+sNjn5Kd0d2PJU1rM4zglFs0U1qF+xNFoiow5Gs1dKdGAfs9hGjFd
wmZIbOD7wgUIMtCJKt0LpWlPoObLdZGts0FeJk7mQbFJaCLVVTgXlumA8836oTsy
f/1ZYOnVvM2mQp5KBKlaqotDegqEoRu6r8/22Gbdr5lznDKBPygoSmc8BUIk6b6X
qi1HIc/fQibmKyNZHL05sNPbrVHmJfgM84xBJWCzxn3R9HqU2eLzUtrbI/otTDpH
2AbkOSAZgT1PostklYE/3kk2wIjMoqqp4LmTCgZsv6wMT1ORTW9dQC1lf6SDMOC4
/uiCcx8yRgvFGPO75SLBHluFLeCeRkV7okdTjXQsB+ZJgAy1371uYUn97ysV1ILT
nWOLMR8dOM//NuPkxI1yL/LO6UvQVqBM72fXmnqIxM5c+AhCaG85J5A3hYIIBfaV
`protect END_PROTECTED
