`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
snDNJFVbGe+VprjhzAMMs7BKZub6ILO53Tsi4+vl244J4xHIMjG0XKdj+YO0T71W
0NotLZ1gqHiAgy9xAtt7tatvV/YcFHKso53QlbL9Kkk0KuIit90XlZ02UvzWKx5O
VfAxk5kFkvkP2D56WyRnQjq4VubK+kzc1KlPCvsYtyl5SzNXpbS8+bxt1fgzlnzn
+YxsGqBWw3bxxxfZkSIgVRnIQ6/YnazrJwrYu/Gta6q5E1NvzzULdD2elVwiqCEj
ncbhi22lGAFuzOp7JRAYEHnVI50PV014pOcYOn0G5/C97B5n0NaasB4rK3qLJyQm
blC//dktR051qPafEqVBBi1lAomhIz/boKq67AmCzMEsWpJFbaWr2/t/T2jY4aR6
xZIA9sKAklXLWVuBBUoRN/isO6QPfnYp9NyJ3EcoFbuNDrEFCxKE0fV6NgHqhuee
Ld2qmM2SuD7MKt1R/eSqY50fRmXjnK9gnCGdd/tuGKYySDkwtzcoXr8ABvTYw9nj
yQ+C4F5UaS5hQTnW4ekVK+b3eX3iyH5bJ3mXpXTogv1LBUYcZZ6AO4jfwL4FhBwT
q3nI/tNzbJuDeGiMEpk2/6ASl7kWnQDlf1RZXtgLnV8ymKrhiglxxKdOaGIBINgs
35PxGNchtAGn6Kw23F+ANhzyz8OGqvMywHiPJQ0wnPX6qshmMyJybcAyxC+Orm2b
91vK6tERzcKH5f+SLs7k0iZBWxsgtAlvOfKPJpeRg8KzFW/aR4SORIwxmajjtTOv
GKltTMNd/GexmK7TYostKaueYBdtpHmlypdP+qB1EZF04Mt8FJYY7ua+AElhXijZ
RFKihiGPAaG+u4VjzLzP2O70JtGQ2ERXD0bPTBWO8OWy1qFBZ3sEk1w98nn/nE85
Vqi8hWpeqir3QGmuvO7pqSyhLeLRbHx2I7HKCAEodN4kPVHsqXVKVCg3BUzpUTlT
bTL1M8Vsek8K1rpOqMjSnp15fyOFz2DIoGxWk74ned5xgEkuZMIvguh09sYeYwT0
zx/pxjYu6k1xgZwKaOy5qzznRD20n6kB5nHD6jq2AsLf5CL7rQsm05l60w37V1wL
BbplLh4Guw7eV5yNdo153ADz1rCX4VUnzcs0PGT5lBOW16pwE8fjgADMVzkKV108
7fF2oMMAhFF2GAp4/KQy+SRQf3z0Z83BMAIwoPbFixoe1vjGK7y1snVMlqruGzR8
yw4SdrGpW6Eqs9Ceh0a/8nzTRR3gKpGkPwQjadccUvxoDDbHry146J7HN+94kMtX
AU6Ajb5OycNqOz15IitUr5ZKsbpF0uspC3UqkrRfIEJAFnkb21zMOvqWRsv6hxe9
WJwHbfIwdoplmVboTr3XMCtFRjpbVPsrpRk1yGqLJkQoei6rEYV6o38f4LPQupev
AsdkFZOPCZP+eA1gahvryYgVUGDFewxsF/FS4QdOw8qmcVsYJIXzuLQehAttmqVz
dZP5iW690VydztY53A2p0D8rpT4PWj64TNmqRCMqtpQc2CSinfTRnKJZUdH6y/kH
WFGhJ/AopWgGeIcaCulbNv3kEqz3DwFK75tTWIEzWcexRGHmtpRRR+LF5G0z93pa
lm0fPjMDXs1QikB1A4tmyN9YyCsxB6zCrXcWCohvGSQTjHXmCrcZ81eYAkaYZG7o
aKFMQk95a8HTDO26U7KVMVGD4+yY8kNNG3X1rH4IXOESK1KE/NMzvRy0I0zmtL9R
Kt6wXrXDtjmXkFTVjEDh3RH1gPnZ8ZML5V+xCoNVfU9GZt2ISgeAHFlXcgVIXMJn
qtry2zoXHXY6+l6b9tQ490rqnZMNpBq7T07ycPlJ7oiZCKT2ruO99QHTe58avWpO
Gl1oWYUG50jONxs0taslA3uAQOCQk/f5wFGqRBOPo68YQ5bcLnL0/PqLcOk4z7dX
NT/FBAW0roZQKkuPcpgzUdHgJzQQLj/xbTsieMDa4Ayvaexee0ER0OuJpI0iD4ui
WJOlspiocRYIW/a07t/M8/dGFi3+omZFivPxKDP0uaGKDdwCnbBq9qpEtP9dM5sK
cnzvRLInIV9vuRQu3zzCqbTQJQiH3SgP/iKfNjfqvuEeBo0U+LLlpqtGE3kde0eR
rTE4ISKKyvETcCjCLlzI6+j4U58JMuFN9dTsJ5JW9vONrzm/3qFe9rnaiy/PiVNQ
O+DYJEp4iGi9IYiWg7gaoqZJVe2KQItZsR50nJHRuzd7+BPrYHZGdRsiw23vJcnU
rIFRCtSXebvgjVbAiq5CJk9aCau9XGV/D+SBxmc3rZmOzDw0IclwTxsMgaDclOg9
WdJTsP2KtAUxgBKw8QtIMGrejnP+VoVE37d+TYxIpU1Jhq0hZf4w/A+D5Cb+s6+z
9qgh50XL6Po1v7Kuc2hLvbPRqxHIJtOgANpDSfGqKElfuC1WCiBfoUC5eftavRUt
lxJyjQGwmWQXhGGNS6g/3w9QKKaCHzd3ligwd/LKkggpLUM/Pl7/PGw/ZaPthAYB
jcgRjgFaksvTr9XNGAHMJJQRA6X5iwH4Zm2SY7+YzMCex7p/QOtyQH2O+lrTb7ua
MH1/kYpDHhF2wPLZ1htHyYZhmGeGzpYLWz0onvn9w0VhM/+lXuU80/nnrYs19ctM
QO+nUj86WbBMMDeSeXeYHklJG+NwMpwQ+xvEQh7X71NIXa5zLl+ceEyJeEEDjBkO
Fa3VlCfCfEFMY3Yt81+QbN5qmUSOpG59mQYZvRW8ZmDY2FMflxuLlMF/RomAZtJY
Q5kFjI7CMpLWMiPTgc5aFrhSfC4hHw1VHAGiuDNK6OC5bmjDnKHq9skpGKDz8hxD
G5hpl/8b/9LVX7ReAyNFa8KaMU/8b+8jpPV10nzeokE15OsodjpmPOpDNlvpj1Sn
BCYCpxU1pJkx76KEDazbWiz/CRdq3PqhpnPINkqdoxU=
`protect END_PROTECTED
