`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MrGjXDVnt4nu5SexXezG4T3z7osN3HyENIJmLg6/EYzkdgAAf2Asjdv0j7MqFRHa
aPp/Qv8DAFso0Z/LIBamADpXxQDnu6B49Ivf3/bITVAqv8054W/G8gVHeTdNtfRO
mMVHBbWLlmcYXmNFLGlEV5NwhHwExBCFsiLDyg/7Dysz9PTmSymp+kRSb0HHm9Me
so2blWy538g3TCUtYZ5l8pZbQwYaioaavtA/aZ64SWRIAVPWygni5pg8wFvX+0dA
KMAnj9dmPTpigopPjIo+KOTlef3LGFEMEihAm0AsuLFxzlTLR5lD8JsoZZEEw1QW
FYV7xwbOrSifMuKYvzgjSs3eP66CrnAyDvo/JTxULbMPjRZrOfA2ukRGM1qwjHvz
AetTbv/TEBhscFElI/UDF6pUEA3G2BlS8gznJ3OGdxKCZzk++CFxDWkg1Pe+NPAw
Q/NdkdtkvvR5eRBE9pNuP5frIZhkSe2RtrZNyI7bqbZGAMLCI0jDRuM3FIG/4X2R
cpWMqrGByAr6uwzFGGejCu6npaZa2Jb6jmgch98IbY0Xcv2T0RVvvyc2B86dPR+v
AxXr9X/kZv3sm6bCW8+LRRpBPyZLzOrxK/KNhERK7a60uxyQpNhLqRWwjkcAVj1F
USz2KgO5pZS8SAbjxtaSyxnTmXy/kaLWHodzTHhh6Tri7QzTJNlkaoPs4eClX5uC
8R4F8sYYGCUcSaxwtEEQmQdxqDm/2eKEC9VNLVDCM4Hiq2EQH0YQSbmIPML5boHW
ma3LhhBtHNizqJWQH/GFDmDhu3OI4w4Tsx4KiaETP0MVWjrIeCAE/7BcDjJ2nmeX
MGnrOksAGwoc6/+YekK6SIRyUEFMBJ92BbyL+lkVmRI59lwCpGxUOmf+gG/RwCmm
jEzPA8AOzA3d2iIQnYSwduFpcMGYjknxMR4tYaTut3SVM4ifyp3XmJkSb8diLCTT
zm7z16ZoGPeVi2MN78PuF09Oi7jPe1jeeojo14JKG3SSx86OZCvUwv3jz1pQVRtm
ZEZKpL02Bz/70ZWQSO4/IDspp1I24/ZcrnGbvjNrm7ErR6rE7MyM3XyoOYsfTp0P
O6sqoBR23C9FcXGbGS6juCrlYg45YjXWZdE51IFf+UMnBKpl6VwdfYU8sUycIhxR
jyYHFhcBd3iNFAxzr+WIwfGnPBBF4COjv2mkNfHtE/cWP9MN1iHBvLf6noQHr4L+
81Pddwv56DvOmaaMBq/O2PIS4ZEcYU056/DNvZk2+KlsgR1y6OkKMXeU+36W/HS0
WzsNT6B+KBOpbaULVm3jNKOXQzv2WccMlt+kJsRkPcsBsoerfoMEL4ICIqF8wfSV
ZZfJTUChw39DyFbxVxCYGzhfdN7jgqTnUOWs9HMngLAZh2MYaiVrOlL6qcPu83K8
ZCaRhlfFxHrYCbN4yvhVh3Toaos8KbZJX65NtbVU/Do4wO6EMD+A6qdsxWUoySvk
gzLcTnSWzDIEsfzPzruicj08pxlKDNfZNY97oPN+5zxcMn6c8V2eQrJ/MpBQpSkD
/7bbT8ym4nNzdqqAp1s8fDYLy/8YSm9EQZTx65XaKhttAGJSbO0zioqg8jGyBU8w
ndZIpilKhX486P5GHk7Q69rAKQV06KEzn6p9yUsC/GQiZjP+SLpL7+yecvfKtZeC
Pt3IWdoxjC2l9iOeS4GcVOoPjJSO53Y5t2r9e31EaJbjJUlq6ZOlbOvK2/C5+0Xf
wJv6otx9tgoL/NPy5bKlQY4WbqyUztA6pChksV+OzJb5LuOKflU4ytzB8j6UiIt6
haVQEHzi83TRba4go716y0/F2Fy+gVGCxI0f2X0XQhdD+cLxzg/g4zz5IA460hRQ
+hBn37F0L18fPZJvcen1uKTxjwlIigNW5uikOiw5ISxZdzPrgdyQuown9HDr/MwC
u9LY+nXqE9C+tleQnaUh5+mIhkuTQCZON+LeUhXL/oOMZgFeA0m6Jh5j5Au7poC4
iG7zV23l+wq2tXDB6ASQIf3H8ETCExWCr4dYJkbYMYrlAALBvb2PMXgpI5+mrMIC
9GkNsnKxJO7UnCiLNqKrQcsEoIuyRfBlNzczZQmb8g78LDY5W93rxivE6c9VbBMW
oxV5exvtR6xSimmU1Y5Thf8ZYWOtNGJpUb5wueZfo8WFBNl530Oo6GSxQGkmd9FP
DIUcIsw3m6PCAhskDN8sHSrocexYrEWzwYy2jpq2UaRfeiGiFxQSQ9X6lJ4p0fSe
vpg4UDLCMwmW0/7+lXfSiLGnmQyKsCHo5vUcDT2vprgY+kRC+6rcmNQqNl9FtNw3
WyFh1uHZjuInce78BUhVqQjJkoHo+uP1BhLa/Ew4Nf2p3ha7Zcly+7451Qa9VNfg
lVCLhHR4BR4j3NPpf+I2BNHoxVJDN8FOoSFmVryEEMhVMPpiKEtnlHAHLffU1ixS
vYa/jsqAm29f5ci/aGLAjx3jrQ6bsWpP5oFRarORkd1/i/juUNRfZ+V1IbR7Bt+N
lvDGHvtMw26SuLgjsreWzTbORm83nBqkPtEXlt6l0KeEHwDJvWdc7lY+XLSUSTbn
ZHMz/Kql2OXeD7xeGnoZTdVT1xsMrgbZFT64sBtVUtJ7KTBYxxzAWdttBKT/DDuJ
ngdwax26qkiv/JiZjoG+QlGMWFv2U5rLuCwW5pSFkPFFFq1T83eiFLKrhHw3qcZi
Pq8m1JB8p58AyAE4BjJrLaf/RPujqXGWWDK8fwbPfK/1oHj4wMomqg6IiVQU/ISN
FIM0oRvLO7syAxQlMNKEHaDeVSK+SiES1UQmRLI4zW96JDljbmUeW65dh6Mk0T4q
kSt61vvYnyj9vZ3LdPVHwYbjlBzTF0797D0Y16rfwigCRzu5Yg9SC4j+Kipgclub
usVIkfBfwLBLfwn4cHthHFVD89A2rFo5WXcsNg+AAjBbnEQ3P67zIdfa7Yd1u+D+
/2TS4QFhJ4QLGMeAn5tEU7R95t/4Gfb7Vm2HX/hPYRg4xL+lGJP7lXxphRBggnB/
u4jAoCdESGNu9xsrYJM5BPmOgmlP+v9H5WwKJyjhUi89Sn4AA6iCvhrKLmUNEqHI
83DN/BR4c90f8cSXNPp/NjuYuAOQIyGNb6sc1HchDX/asacnWko63jd1D9cUrzQC
YUz8cEtLG3SSX4Vj1dBSwLtTUJsj2Saw80y934GqvZ2sbBjovesB2DSYT90kJDM9
IrI2CxYaqD8LI3YQSscN5Xk0Q0XzEN2L9XyEm7ixLfGBpMm97nuJLM1/fszbsS3Y
TDq77CNx0aMlrBvbin+LsWrsftwdcs4iweaCsaIJughP0IdWJSmy6YI0+89Cj32W
3JPEvAh1g+lKYO52TB9eEiZaZAw2euXAjQNnx7hqjjzG4fsGEJvwJjITVjQZBmwO
6iHV5yc/PM6ZEE+M4ykBslkPIEzprZ7EVHWq01RuXOtEUobJUhoYKw0DGH1pJtO5
WMYKiT/EHyBkJ1D2Dp7GjAY8QL3Qga+8aLHruXfpd4NuqJhOK0FLexkajuxHJc1a
Cp3YauRCpvPiDCnbGqYaAMUokf3xSz7bOkej20QnCTzXdlDjpj6ZaMOlHS8hDxZ8
jAGaeMQ35ADvdYpGfL3+T9syF+1T/xSKv1QQy47UdkmAvm4VXqAqnQpvoBUexBOZ
i1dNT2Qw9BZ6a03zuLrDPPFc1W6Vr9V/LPifnCdPeVUjeL+jLXChYONVP6q6apeg
+hE7O+cxJfIQ+CNqpohDiusvKIN/4yEUQTYh7hDh2HevzvJiu3DGej+STORIy1Qd
uJxt1eDiVts1mbIn6xOWBw==
`protect END_PROTECTED
