`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
frjy5+pb7zfkmT3pjHXk52I11Rb9IsbHAvqNlqAex0saAYNMfBP6Bo8jFxkgeCRS
i2lHE9JfsBb4Nl83hnURTbfTGwOH/xfhf+tlIuFA61N/dF1UmtBDjfCHeUmCGtHg
Pt5bjwp4pq8fanOVJwyd5RAWb29QCBiIROezwt9Ed1nkbE6R+VpZkWYVZJeJYcBU
v/eygM7YersueEzCm+xfdQwh+Iy8ObEe3ounrrOf3s/ZHanVRPXG3qlzpKJcX/if
4OraOdAzX8aaeAD6DdyPiqE6AePgDTjlMfhU1vuzPxeR97lULmF4ScMLSc8xZ0PX
vQ2WznTw5tSPNuHjAXt7Wqjz+G0WD5e1Vnz5i9vg7dxzzHtOGz6G+/1Z/552zriU
1OLXL8JHimvV9wPH+OACj+/zUamw/EkF7exwmgdyN+pHPjTOlWKT4NDjgh9Gp3WF
0YnJ5QcUqIa2ktupp74rVW4CnzDgLExq42EuFcsxVyT3klBDXPYaa2YLJW9M167L
+iVOSCUYotM3jAqtSYJsHdBRF6AEyfzV74xgwdoGMrZjrZlAc7Stxkt2Ms9JjzCt
VQpBf8Vp/oTjenCQDWySwD2AgDY2dkKzmel6VkAjuktt4VorQsuSrN5NbKXJavWl
rZUhueOhJFlfMS7YGGvHORV9cTzNHyWS2zOPZQp+bWbYo8NDvE4w//XMbTMHImPN
YNILnmBzTKEu8WWY889WbJbeOZDjB7/FU/3SOM5CPBUk9tAu5YGlqlzdsiWkb1DK
dqgebHB4F2HXbv4+bdLXSPHokmLiakuHMtR/jjzQKs9chj2bwtSsjQIHhKvCiU6X
my25e3qSOV1D9A9d6dYP6zq8KdeZ9U0zJtKjS7O7BXLUt6RPkNMwRw9Fb10sIjm9
eKb08hpdvMq77tQzrXoj2MfX1iXRecqSKyHpqvv7+f0+J60C/0dpt3ck/SIkfRMb
sX3MAwEbWbEa+YmN7d12GRPLk7FIbSA8HNQ6zVa7CWV44liE9ptEITmDTlb90ECe
iXs89GHhmrU8bkCbPCU4IT1d4RvzvsVXcJCl23SFz+dhTtYb43RIgrTESn9PNbUC
XgBuIc/K783dgbHiUBNbzwNHHfAP8d4elr+zf0j1S/s8EFqPaSsDfiA5nF1bfk75
OEDpxvn8rM2ZtqqrjeQxO82m1DOI43/5EWQRH8tW1SbDNhzPDMBat6H3k61N3e6P
Xg+PKSfuAxLg8GmMaGSwbwTnRxxBKWWD96pSF1A1qfI56pWojDsdv42yy9BWTyDL
tMQBUGaoZuyXjB/5S/fYjx93hPcFTQOL9fRcI6pTM416T1qRDVla8iXrGyarXYQv
wU0N0Yp5utvtuL3KDT7UNLiX6GHHpXgvy46zRKVBnuNbIvRqPPbE0CQ4ykd9k3sC
Cppb0AHpDBqqvr2slW2J0tCXFdpjtMx/1HTrsQarTod6HiQ7m3MTYbQyKJIOCG2F
nubGx2N8yQ9G0giAvvWpiv4a3lYrKJXoqdGdoE+UK2QjTW1kOkam9QM24C1hmIoc
7iAPcNfCwuVmZyEOnDTCMdvLdCgr0Tf5WIHicIcn9AvqDMy8NE6NIqvojqpUaAwo
8iGEGuCeWnWBCI2+eyep7Zs3YgNYfDuzvLYXChDZ25t32Ekbf5UT46OD271lnr1d
pMIlisBV90JnAnEVlXo1418WRPou+wtvuck4n49LVbRPUYjrgEJnD+QBFOE/Qd8+
Dwl5/HFZ3ICCCj0/+YlejCm3jGElQB1f1ouBQby0jADlwxBiuyMv2pZ05qm/pZPX
aNZAPAkZC8jWiHQmVEonOgM2PPv2tBhzt7JrwSpittN0JcnqdJ0Jp6nyg/S2yA+e
7HQJNCChAen0HINIoWzo5frKLdVa9tSLowiGpVU6uToATfaM6fzYVdfMJ/KltYcp
hoeiOG8OAlKnDTzTxPGwhIcihEf8cROEuNg/YIN8UyxY8uHq58prYAXVFDlcD24o
vKXshBy5F5s/8xqMv4i3sIsnTCPqHhNTiElaSosgZRy3e23aWQ558XNrfO3MJsHp
sf/l9EazBiVrsFjfUKa6CxrzRjHQ7LgJvtaeHNfzdUB3S8bszKPuvuN2NrWovAXH
xxwUbmFEfqd5liYUxZI8WiH1atbcb27mkNpDA2La186+AdVcu3bSfOmxBXcJ0Vyk
7LLim8HhfHA1iKdsQlM+IRI2rtHO6pbLyKKURIzR2LPLGFaPSS1Vj9IGwTVxqgEY
j6w2GXrdssyg0gpzfZ0Tuqusb0dqAGqGIBb+SbrE2WdzHyiDObzRUC+t0L7RnuHZ
Z/L4lyQk3rtPkKC7sfs5nCoh9/2OEvMTLguQhCxf43EpfaMb6L0QrP6G/ieo+24O
zdiqXMYaZl/PLV8cCp090v1w1S5ke0wPBWHA7RQEd2fjLr14YNF6T5KyRxrbPKtI
qNVXqmIxGn5Em63NIPDEaw1r7NnevzYDvHK2r4AnihyerbzAtAcuErdK3OD4pPOf
6j2kfDx7ohi+/Xpsg50aNffQuKEAYuOif+RCPryYWZFcTHcSQRCXXa0MHM6+Mk0J
zHvMh40F+EV38aHuE6AImzM973svH/QfJ59cHlciS/uCnvd69PF4Okayx+9aMR3o
EYtq4SjSeWLZd07v9gkkcSX9En6HW08fSd4eZJRacDlCscuNWMwIpcE2BJlfU8JO
CsRvvIlrvaCH0zpqIxVgcfwxAZq37Mq5sRchNPqhQVt2HJuHPOzQCxviYai27w5C
Qi5xx8PgBE79ut5T6asZ6rpLfz4fpmv6EGBo79Xm5PDbJvKawHjyd+GylKCjsfst
chGgFO8XSu/BEC+J20Hqj5BUcH1FHKIMzMbMluvM35mw1b28DdJd/7TeqmzFgF2s
QyjameYrGW5zOkvLtAJn7+vL6Kmhj1LYSH9a28yJmz2kxKaMPI766/qKpoy+e6gz
ZoehdP6P0o+S0O7HK0mxwrJp2D2ynnrk15o8ntummeUBJhLKABHqKjYA2GDq7FrQ
kPktNqVqXQa19XN5M7G2YCOs4Hod4ZNsZ/xMHeIaxsKK2+bhKm2AlSVCr5bXHC5U
FUqGT9ZS4Ot83tNqaYviPQ==
`protect END_PROTECTED
