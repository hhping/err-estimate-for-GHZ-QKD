`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jm21cLIXY+9CGNSW6vZ9mmQ/tl407dU8XiiWYKW4NGUbT6TBSKYBmmKd3eTLhi5b
TCTHfpEDNR696UlUnJgvEaHJX7SGEXFKm9QbiH2J561bAtBt18vGGYSDJ/mU5gDu
m1GL7G0016dXeJWQnRXGNGwFnA4EFJwwH0g/ElkVfKLvNir+7dlXCYpTJH1M/pQH
eSsXi9DECkibPlrXCPVc53j8Mm/z4w7DQ8KZFvdT535n4uTN3YxBCnDMU2ow6yPJ
h2ev4NPhxiTSz0WfcLuoQ4R4xD9IlzKNxLkGfpUepGm4oDHxhIBBjh8VkPd1dqmn
zcyvFeKl8dhcSrVW8uxr0BomezpP2Fz3Q4bq+2K3IPZfYbo58g9KBtjnc5r/f81a
VUfTz7w9mCafiahCbkW9zFvrwHhbSuYxOnRvyMxQofmaiuczfdwXArtsyEWkGr8A
LxLXumR7wTWEQ5il3WWVMHOU6zA6ugbTuy+OQ5CnHetjsNHCDquQEADqnNZO58V+
34SCEg73o7g5wiHN3zeZ0qKuBI3jmJzBgQGZF4lbofBp/6Sn9S9QebsbViN2dcJQ
oj82pzfSSkK502mzy8JBuWIjmnwkTjkq/SYWHsMOsKuy961ybFyVgSsGj1yKrcGn
b3EVaM0acXibXhNDHmDTzeBE2FUB6wxtWvDyA3qZpLh6NIzeG1qGb7kil0CANz5y
IS6T9iuLe4c5Zm7RntrbZhyOhi8febwxLyhhNOtr3s4abbGfbY/GCk+7yboBABeP
K50ff8TM8moyccqV3DiW0LhWn8vL5fMI1GYEzxMoeGMfjAD4xWBN8mJmOg3vb4HO
ffqyW2xLqVOPBaIwAnlsTP9eQDSjsaDDwySubzvspMf3voy+LetpMmilC/PAP7aj
QSPi9f1kfqilcpEQ18aIvVlEtCL49/JMLqRrq7xN247LpLUtB8R09GCrvbx02/NN
Z1vmxfPxdJBZNnn/iMEbhQ8Vb3d+oat+3DGTOdxli5qxdGcfow88Omk3AeVWwrLF
pp1GhUvNrrEwtvEwszUkw+8HVo8xwizAgvdQchPe/n/r/FcHSGe5ZyU+LmAYZf/e
D1jRBzDn49F4VxefYT445+xmPY3y/f8FXYI5qtcmL8zNDiQkudo7soyfwqDHIRGi
6ysu5vxPCIu9Fm69UW+MJRdctuBCFM/Ded+/5A9CoPxdmjIK3vOf/YySWSzWiigL
bKpZsyxDYe6cdt7m69x2tUkIGmQdFQL0Mx0RRcYnqutRGteZ9XcP0LsA+tlxfYvI
3oXpB0s3ceuft1mGtzEjuBIEwtBsRVGFwX+nmUfqu3OjoPz3X1K18BF5ZQ8kjZyw
AadW04/qWbi2qR/ikVU7q5jpcF+TngoUsPMjD/AmEixtqYuP4KVu7SitBssmA/kL
dMjvn75JDtcHuI/a7thsRCDmV4U45HLnfA4Z7lO8x4xQzD7VF3dGYOTERAhTf0J6
2O2HnMzbOQHg/vv+R2eZ8mnny7cwIoXV7RSmA85cv+ED9DJ8IKnEbLag3eu+PZc+
Gtx9045NRCN+mGglvgYfJYQ3P36R7TZwiR3shFKYlgCHFcH1vL0VrsoWTaI2IDcG
3G5noLx8FAC9DWAzArxJaKJGJIH3y4cx1bXojNa/NsEA8rB7p+yEfdVXYLfJb64V
2tFD4aRGEmY8EHa/ExDXBZhQ1N5Y178SwzvK2T5uzCl2J0UwzU1DlLYRa3rwkQNQ
+NJgWfjcDwxSvnxSvC9VE5CgCg3w2eIP7TBZYGUIy724PXIjxA8eQWGw2nwIETIx
ILeugFTY+ngosmDxu0+6+Y7YbZcMxAIaLmi/k959Tbvtl/pWoil7uN9HwZ3QbxQP
BatRNMeQHhuoG3ZjLRKT0uw4QjlUJ25lYYzAY62V+VnVO3hTfoekMnX5mSIaF6KW
sXiiBdePhSAJxCLxejatSHpEXVvAApjQ5L8CBWrZk5haaswNb/m1CNtClhvTD1Y4
3zwxiqtyinQ18Rbg0ABChR9g2Fol/PamLOQ7alYnJt4+hENNwGHtoK4xWgtZ/ct2
iFhYem0EBZCH/o/XpL01Wo/PoGJ47xCyDBp4dNyRZdY4toEOpeRPNFku/Tk+mgrj
NGslS0QLW5GuqdZLF3IzPjNQ6oqfjclXtQAc+kq/ze8DfggthUophwHDMPE79O0Q
ACAW6QMTKRgOZVzhGw4+xwjAl1wEqv1eNVYY3ehJdU8fvq0ybA0YqoQ3VoktE/vm
E0x97tkl5E8T6Kd7QRQPDKWp5SQKQl9qoQGs+JPAv+fW8Eb9AuoPRGTACAQKm+Fn
wfsCzJNrSia6KGd/LQwP+qXCfLaEYxxnYZcvgexLswoJTw4yB9rM90kZDapv9/mK
Uud19qOZOt+cWIUH0DODABAGVmDd7YT4cDbjVh+Z+5PRGvL4gE/9cGC/qd/DsRWs
+rtt4nlHRxtYfP89a9pvEhwPmWMcLL1AGp2gfYIXQFnvzNOchnA3zZX2K+VJkXzw
Fkqb8ZnqaY0l8OtmIMXE4VJLvkaqpDGBLuemjROsGqDVBWoJJRHCCHreT0sh74L1
0eKqSMN4aGMOaiIRSfjRCDNVwGcyoLOnLSht0GD9BMYeJ4DTJzwS17xWy5MDGVbS
/6ywnH7o6hJp0MVrmrErIZ9sc5mdqzK8MXBMYW/nhaM/yzldV5RqurXPNF//UEJF
4KHZRCVvUToQOLWDbJHK55WsaJd7eEL8KJMTfv0tqdZE+/MpOoHlTyS1XJ+Q90ou
kmSmqJXArYDZQvUCJ51ATyhGGyhc2f0SWMgnJR1WsGKrcWm9ry8CsqKB7uWxKdg7
Jn9fSxkDFVGIIR4wVwlbFPFJo0RLazTRzNgDAxBDRNwn4KhciOD82qLxHAbMM1PK
591nKVmEVHf+lW8yZroSVhC7VkfWg8WduafKH0jr069pvIdovBnJnwsjzEPS4WUL
vhk99+UjHcUux01Y1tsgsIrqRPEjYVq9tzI35ySw16q9wIKULXJUGUoEiz07iMKh
duQodfuAchSPZBcJvMl6Ci6Ixju4pkyR9suPtQOF3GvWQx456yVUOyd5XrtdryJ9
Yb2X0RqJ06AZK0WdiyCPGHpBfNSh+0PLtMDqEFHPSqFvmIDHgLzfTBZgZAWwktWw
pBXcQsHxI9UKX3qBhq4F1ljs8z4VW9xCa9CnJjFrbpBaQfGkhvmMGaimY/zNtUgH
hnsWxukzqx+yDmi6Y/j0I4DN2Uwj0Ww+OfkpE2pZ5LQixAcq3BY5rXKKGsnzOk3q
m26hDpVF/OpCJ3yUbO5RsGAWPKuQwL5v6sL2uXvDd3bsH7KUmmrWWIvmlNz5uDeM
cRawuyB1kzyiq3UcMMHCAWb/Ddc8nt6Zu8vLyqHvncBGf1btTqaJ5qHMdTcgfsa8
yuID/qRO/ZSJkDUfcVTY4sbwo+j2Q20lfibS5SQxm8rouL8sD5hc74dGoJ2BVzsz
8TDIDC6f4xhKf3staNAFqvS8i/xlOmfz8qtwLca4vIpSYYiq+CyawSrsankl7HWJ
ho73kjHY1+CL+WRx6OUR3VXCjYHvMPK89lbvc9yQzzMy7niz+8QlMpmlPabNef/O
yVf/g7qHoqI/zQ5dpVc29NaRyA8dOlrM3TRWbBTUtzKDzlxflzmKGNCaPWTpm/or
mUU92SvMt5YjhyvXOCtiH2YHEETsJAJBGroSyQk1P55nNbnzb6bp6fDfBeMDmjMs
U/kK+iYVARBPb4TEuPM9f/eaP6fqu/wvX8J/W+tcd27vfOYHwmF5c2FYJtW1z+Tt
J77HN5BlO+9W9i2wheB2spfxpNFS9XBN2h7QxffMRD/73ZN2rn4sM0WO2hlUWnu5
4k9F4jQQxuEQ8kKtDt4cfHYhF/hk3sVSM+fsNZT+H9ClvK02YhrbGMuvAHaJoRVZ
H9n/mJRjXV2u3l+V9nIDifO1PuIXKsAf4FFI5XbGXRTy0oN9iFvZb3n3Ls0Jt3Bp
NNQlYfcras1BV5UIcVRkUK+ay9p064yzpDtOnyhlL0HCiTV2B3pB17OJBMrHStL0
SBCJFZPZp1R42eEW1cHjFEXSHgPgRhpveJC14VEyhcSpo6VYbNadlJxph0AFqIUp
jz5T+UXDIFvtmDSu99NPFmol5M9tnmAqKF4G4QS4LDhkPDR5cFU8EtzCh7/SIPwc
yZewDPzJUZTe1hGWNTPquc4ITveiSMF82GRIGId4GUAWmBfn19wZUqJerQQYzdSu
/zJK6WRDO5PthTMYH2jPVXcW6HfYr3IhladDrY8LBJkZCq1coZ1pN6n1IocMM0hF
BtTEhJwf6L7DgQcNkYwTxNZiRvAQx08q8opZojX5lZqN6JzZY/iqs33uxHF1WRm1
xuFysjHJHddyHTgSNVcFG4nslurd9ixDqJaG1V3y22ZZy4/m9rvd+cMaMKVT/zRM
YPMS5slMmLfzPp18U0S7tcrvQF7/01HstuYFKccMcVEDNFiPRk4+XK2PsHFfW5H+
HUxe1dD9GkYA2lZQo6e1+5gNFzMqxQMwhg3JEmB4iUtEAZbnBASU47fCqdgNbFco
1BvsRHK/MKLOXvvbDvWzygMhhMJbxLuoGb8ze4YgYg7S8BznP19HvGJQNXWncsNw
JBv+GHdncxHvKFF/jgre5rLj/La+UYOxquA332bbJhO2CNu324Eflk8kie/7PvDt
nVu/zsYQZiCDQQ2gSx8oqBAMR0eowVZlTvZ3BdMdwLv9JNdLGFjB4wyxIoKuJTgi
dtoSHOHK9Bm3V5BmXozHsYuaZlSa4iWxc/d+yg/IpD9O82BUWwXEJ7+KKXPMpiVH
b0kpCBUuoF/ZsSeCr5za89ZtAzSYSqqHFMI8SdRuM54GDqk2f5XZ5q9MddHprU5T
RWitXzxha3rqkmLmNumZbrzdcPpW8rvvAgS2blV/uZwaIUIGuh+cc6xzhxLE2SDL
BZ207AJ0bszx2hicuJnVmuz+0Mr4+KXgX31fDNGpinQg2m3wEmfJmWqrfP3xLLe8
9HRjr6mAZIy7MTh4s7LFbyR9cRpYJsb3XBd34vkaKT46+4gcx8ezQmGnifPu1ii/
VweiuIe8esdlTX2oZXL93j2jzAzPEqwaEUrgXbw/rufZNr3imdssrUvs9DZQoTTi
Jtj/RqURZIafmXDKW8agVC8SBCw4x4OMAWQvgtyyCB1HBuHPPXpzj+sTS26sRIqv
YInQ/6oYdG4ojcTBjYCjINV5SEHlnfq6iu1Tnr6uLoZyyZY0Vqg6q+i7GYqbQrJD
TPa1bEDWxVbxnomIAJYdInw+72A88CeqZCQZXw7JaiQE0JxZ46RV59QpBdtR/c57
8a+jpDw/AtSb+osdbpbI3KBydkJUU7Xj0elfXzOEvSUDxxH5CC41UALylGVX2WCn
vjBru1epwK5LKCKr09yUc7tT93ogvXUQhrQWwbEhUsOXMA7XVelMkBuFwg8xLlvw
sbv3/yM8BMX7q0pMWdsoWjJ3KjUjXuZJkDFQvYVXSQ1JPDEDfG8O5wQqvtOuGKMu
XLKmYOpIwyUG/N3zXiChpjSP2ZuvjifWDN8A+BzRf7CvkxLraXFt7QE4Q528pVQ2
LYT0Fk7R7POvAvkrm9973s+lSVMoXwE0sL4oQfAlO7dOr7o2gx74F8ZQSgXq0i8R
/kJqvXTCFiCNw5Bp3GMOaikt7PpskLYXc9FpQGY8Is08DoFjV3A5eT5p9of5YxEG
TyA8ZuFWrABdA7bsKhmAgTudg1+oUJg1+uL52uNK26oYvdZip/puHiPAeRQh0AAP
If2DhCGtC7TwATb7+cUDkQQrB3WOgiDQjwk25FtJ5MuT8RyvlDyHC72iIVJjSYZW
sSixJJSrgH2E1CKrNK+RBVt5tLtDg2jNtm/9YK9uHdgzzPxmwjxWXATL+hNdHzOi
VCoLGqY8iFMnsuLXKcJjLjDcoe6UGE+73isQu/TZgsbeh+Tc83NOXgJbWTVK12Ki
7J/wprjOvtG35Lg0x4lHfqCDadBY/OiPWIjPPzgRvIuGOzsZuDgseoDEDi9NZMaU
Ggy2Hi1zqJrveSvxDqe34Vd+I0pqAXjGU4WLiKpynUQjWmsprpyPWhQZQiCIWykh
PKhMlm9otuhWk9b4Lu1chgAddWVAJqXUqboaK2GrMQzxP4PXO2mnzdrY+7S21Ic3
+zF5LewEgRTKeAGHlLIKVT6ujsTnkJo/pazNxLw5G0fg/aKrJQkX0gHVoNSFAatx
b+EPvcoKmqOBmJ09b+B4Rl7VmBFvhYYBuJBGpy74Uy4zn0wf515ZAREwEI+zGq2q
3vGvN2W0Rr/G1aJWniDvN0VDbfbxCexVaGwkoeiLiAD5SErotqZ17fQRgG8IX7Vh
9CI2ObANeOU4CQAJmnen0AS9VscL4fWPfHJKjboAwveD1r91bqcKR9OHiaOKLsO5
CdMOsP8OFVBSQYdZ+iSHOfJpiz2TVH2GDYKgifwFKuYQJoFwzN3uEuWt6auxLMey
KdRcovLsjZsKFNhFm2CGiredv3gguVB5+cBrMixbpMJY2l49p8QsGtid6jYHjRJ1
2FGo6yJAX9rXj0Maej3PnuBMVJEbOTCXHMk5xIwV2152yHNVNLUbVmccItE3jztc
7qyVz3sGJHEfmgOI3MB+Cohjdjo0wDet5SmpPGeKkBu4H0axZIA0myajWMdTnldA
H/+0h7pD+/d7YywngxiUSgz8PPe0JdO569HNZeIAd1XBRi8JMo4BnmOQdP6LjNjq
ukiTlbuQx4ZqpNV4jUFN5dC4KINvEV/rMpffV/ndT7ZwhX6P8JQm38+/QXY3KgCw
2AW4x4YLHjzsHouk5ooonJEEG6ff/bLg/1EOgs32pCxRLO3MLcqxIYyRT5RE3JEi
jmFn14O0imjkxSzMmowXL33VCE6WhxB6CRg82eJ0aFYE4b2FL7Q9zyc9JXMxyWRq
5SKS/X2MqM9mHiKbi1LWRBRbuoGQl14GG0a3YT7UEaYBxIZvUWa4a9tmF14E2QSO
Wl5B9sXud8VdGthC7SPMPaQUZiQXzD6RyNbO1RLC71F3NOrcLjA36m1aC6X7N5Ji
qTBuyS6lb+z0y65t9Kc9DwS+Fj1+Zbavv7yw3p2Vkrub7W1DRLdcsqA064Skn5GP
4P+LPZ/7pHQZDA13/spQv5bwj+gWfJGnkRayBMkT58ydQcWG092DWx76X9rNq0sj
R/aYW4ha+xw77Vj/g3KgtaP3GbKAWvzn3dzyOmbYZebFckuNO3WWTIC/oZHuJOrs
JYV5GzlIvjowN9g5s1wHTfkmlQiEPpqgLWoXT7RbYZe40QnEy6+reJ8Q+cTFW58D
d/X/9mvE1OvDKJH2Kn+qrvWVLbjDJLa3V++mNp4TTWb2BXzMSp9/O9h5dp1j3A8l
YnogCi30dgUzceNqD6rDxycQi0fz6VBf6kQFbLwxUUwTzU22gysiiBkt+FKfgcKC
DZHN/wma+0dAHr88Y83CuAXCvMHMB0/x4e7usHXQlldYcrvf3rb+aoVxTv0bMjCf
+DqAtwifu+Q1V3dloozmoj9cDVCAv0gO6m5pj4IQ88iZ9PGAnHpBISelWRJZFu1R
Zs8e7VALxhcpdhLCl4cX7HsoG9KoueycDgeNz5wSvlN6F+hDe0G5XPvsB8Ju4pG2
2VOXtF4g5lMC/9tpngZJKI09zipi7gaFrDFQaO+E5AmAlza0a3tWdUlyHaMmPoso
UO6nCMXyMa0TV5PLtmbEIGYzUB4sl2C2scwk7htSCFVVLN4Q3SJaTuOeoJUZQbEG
M3SSZQpiqxheDXcSoipYJbHF4DaUV6o5JWLFTDBWiw29P1mCT2ARtaspZKk5G88k
cc7u3l5YrokWCOe0CauhkSb7hTNlhZgDIoGUH5yWRFj/UtBvMzSooleoJVQq9qV4
8jBUOpHiYHYnIsT8e4yQ+XsekXo5AEzdKVyV4XlIhhdQADInFWhj0DeujpIznryH
aJzjr2uwOMCZPbx64MHnznvzr0VqqIkfo0THsMwlpSiig3YIkBrFWrAwkzZr7shZ
wwsxBtSEbo9Zsx6lXw0sNvboGL0STnIEVnaRdT3+qEu8a4fGCe7xrRHfaPJGc4so
GhcK6Rf+QUrFbC0Zv9kP/ABNDb7juDIV+xc14SlGSeAEwE2re094ouvxJfn6enGZ
50/yXcFVaAOuTbJM1ritkznrn4U3wdW57cLgXEuelMuDS0bC9pc3vIzU1suF5vgk
GD9OWuvA91L/uRza2J5g/CtCemksSKkZxGSqbTcnwrBprRUPI6U56JiOfvWDOf1a
iQnKw4edLunm/u96T/B3gIpN3LUNcFVlBl+6T8BntEo/X2QzOwoN0yWRe8n1QGUS
LDv6sI7brtOAq8/fZzpefkDsCGRnzNrVdFk4RKT2Qz6BmSiggU3W/WL2pMZctzTK
jhm8QOEUNvt/AJRi+tBGi6gpB6VufHYvcGga3JDvEtLTxtSqtItRLDy0vcwizOS6
liGsjLX2GNz/xk/K8rC3d3f3AF0f+D6M4tPeg2lKryMJ0Jfm4Vr7xCV6k4cPWWLm
K/ZDQuBVkeIbz1jk/qOdbcWu5qxnImhk7n14Fbq3ZoYzSzamSFWaUaoumZfRXqa6
TQjV+S5GKUCrDjOBGS5DHX7EcfHkSRivl8AsktkLihKV6pRvNqwVtjuSdUkiKawd
RiSiTi1tg9UyRhj5WYoUHY1iK6QILe/BzNiNY4hYWhM4i7/I4sP+x0775R+2st2V
SXTm2M2Hyr7jBhN0tBgrq2swI1V+ikLbo82zSpiDPPNeQVYzuTYojhvdLG1e/UVT
yAcUwXyw0SbVVof2FGeKT24WNtp/wbRdCrLGcgwYbMP6aRP1zH72hFwroyzo0t7D
81Ss/AfNG2QeT4bC0LDYbgmnR2r2di+2VGEjGudZ/FJXTnJaClIypn0LYt3DnqCz
UZDETi/NtOKH1hlK0UTbSfZo3Si3+2Gyt+a9qNjecTJnMO4yndDH55cWsSsKXR7D
jDrFVZmjqzqr2M5jtveLa2muVxpCltoIu3bkPZj+88C5EcvA/ZRGhOMhCFUGRDfq
mvA9w3QzNJIfo6zouaqV1rjKXggkukOZQ3AxEaDu24Dr+vt/GrhxbJxORH7LCvyh
nOfHkaYRfpcOBr/TSsAav6qjzCMxUt0L9Kv9XQkJyZtJvpr9MhKC/HSNsoXuYocU
Iw8aJbItWXT+HD3m0PLX+5EfGZC+KI8g7a8LTKvjiCRZTvZX14mbbDRZ8YorR3SZ
HGbP1/cXo4mwTKOosF5bHvIWALUecmL0/LLk5fgH5O5PtV5CJm5tV27Ne+pIIQ0y
FbGotJ5g/rxDXD2GlFWetOIMhWFjZlvjbNHMEie6sqtz6XcWbcTHvYMb3H7MrbJb
om7CZwCWxj+nLI4pYcLHnNqHCGTJxBTuzTk7OV1MOQ1lviyvd4a69b/uqOUpNe2k
7dGZhLBsQEO71oxuGa+rlIa3cEt1pZTWeotaMoYBIsIDsRNCs4UyqpbAt9G+2SHP
+yBr00bPVgFJVlfZb4vOqyX5WsLC+KOE+tcqM6G9/2cM7JgmlOUsj9lvhehF/BAU
8UpRVCqZHXu/HPBtbrKa45dJTgQtDXisuClN7xj8M4CUa6OOh1SU6ogrRo09ELVT
ocOj46qyZ8bUjFspTi3YlkaBLLYr7IOupdMqULSoHtErwNsZkIpXODQMQWFc6cF+
dIt5/LgpBa/9w+i8R+nQzdB6Ndrdm8kLPHzZ2V8ig23y+tBDV3ETz93mm2RbC7Mx
tHeVjEW8DGt+LBc83iHuXDYPcoW+/M3r1CjkdN7y7yUQijojDBfdT1VzeMeY51cB
9dlH8cIylQPFHjhtIYxuGqhl01SHWV7JFLJ78mm4bjhqOIiYYP/TNDXANe9hj+QO
fJBETyGMu/i0xClYX2c/ASzt3Ot32TFGKlFfeLIDQMvfTDUNigY9akiVKR5HeO1T
lJkbO7IEz86p/o+VqavwVk+UI/TgJxRHoMiNNHrSWOkvSXEEHe2p+bsx/krdZfvO
0/7ZIphx50bj63toK7xwPdGSJ/DhaAUcMBaXpMgxTL/z7uR/Oe9J92tjACJj8km6
MQtQ/YUgXfducALsfrtYNGD4mMG79Uij2kZMHXkcWOjhmyS+gbGgvSLJeZE5ShaL
0NDjns8NqatMLjg5aOJ0KBde8JSVrp05fFnnDsI8xHSjA/NaZAUdZIeKB3Pymgh7
EMsBqRr1ihyygST3ZKwhLmTPYqqZP7ut8ZDnuE0EM5jxbJ2tCn7WcyTUjcK3eOvK
+T/QVyPzXwRQmcF71VrFCSk8dyPmn9cXm8aSTaiZUx46kLs6ejfmqeAr1LUOfhfH
d6XZkyZfr3dHCdVo59w/oBXwM7z2wyAi12D90BGQ0i/cDlp3PSFF1oOtZUOlmt+0
II6TOAE/iF9FLqSPDTL4kvOnCiGPVZ+b/nyCO9TRYR10lA6XhWGrlEq6FH6NhsoG
L6Dl7wEt7X3cQjatlrR00PPNVhB7ahZSCP/sANrzuH4+AKsP8VY9Y6LRESU247J3
zlHC9PXpI/1w+q7dTO4S69uSCo4fpNJBRsItapdXo0XgUJEvm6Y+sVDqBXHN0NrF
6ZHfzxw6PAZ7+eo06xJNq+V6W1cDPO1msMvPuj9T147nPjN8D9rb0epY776RLNJv
RCrBIJQbYbr7zvnVsgqw7+H6lA1i6NCSnUFMCGHikySDwc6Lnxq7shH487jHjkCY
t+l4cbMh+dJLiN/bqZpVyzp+VYHfr9GQ88GSsiyyV0cfa+68CyUm+oyTt2hB6Vqr
wPCrQak6uwaFDtlfF+fO14DNQ15UQ/U9qu+yP8fbeB618fPwwG6d2beGY+4cYKPP
a8FDxQmiO++2C6bq0ZQmo5Jhg7OCeEcet1pZ77joH8Axfn8pqhCNrfnrm8nybIu4
f2EbfB93o63Zu7y0mOW0emcws1TPyAjlef81wcf7exlj0+mtzIX6lXEL2TLfMAqZ
SzARnCLuqpTGCbhg/AwLQx+ZBUWrABz+cP+32Zzd5V9NpoDG7Wsv+NV6bPTtX2ov
VGWcBOz4YUiOWvQFNohls7TUoL4SCtW29WZsYnlw8kUyaoerUDGq0j8aGzqx7VNf
pzPf/h7x/lQMNm3KUC0vPGicw99JUhNrFg764tgGeSflFIU+yD8yaP6LvibZ7KEU
5JLGPYDi42ZYT7MjpUSjCa9tbHvylVAGOg8le2KGchamLH1MPRPi6PoEsrLa41mG
2KSDW/CMgN2xNchiFXtoHP1wunpZFvYaT6a74vhtsOUB81gNkBkmTdXmqh9cawZo
kofrqWRGFasrrzMnA40+FL1e0UCqKCHoFzzNE0NZWoQfvD50xpZdVJq7HSdFjBq2
aaHX0bSyODW6qwNgQvQvxLDxbaKT8HLdidvohvxPwkICjwyjnHN7go1K2Qe0PiLp
otxCGtMZu9cgrtRXRcw4mpCcC6X16dq04TdHmnmUSbHIg4GuYGd3jU7vrIKBYzjS
ARfHiNO8Q9OJzkv784AT4R/KFhzaQE8sRF0ABVe8dugU403+JRgAD4ls+TibZU8U
DHj+3DFn9TdzjQygG8U3CmlX7Gb9Jt/iEPgETno4R/Fc5f05HkuB+Pk73KkSszH1
LFwvMAQy8kRbCYEK1az2YYS76wbxWHrdUIbBUGApS8AxIyMwMlXEEVJgFC7t+ifQ
JAXnLy25qY1LUwss40eoVYfwLGiYn2qaYvsDDWfGP7HOFfnFuhwgd6EwwZqfTcyA
+Lnp6QhUgcssvbZpXqYctv3n6xmqgjT2kvIuUkID+ZP0EvI3IQm766inJZ6xhiNC
Fq7YHtaP1o94gLB+1fJtGrUcFcK8MD7GYwUKUYt804XKX5h5axxf3zofgTBXzilu
kMu8LR3LmR842jeEg3Ap+hwVpQOg9vUuOhT6OnsPOyi29EUhSUUjBAdmbPBOls+B
HUYVLuQi1IPNKrkguH7KzrwEQ/frV5kJdkmLZ7Mn/5G8xCgNl5sdy5F78xKJd5Ub
/KBOJ1njESAnv1fsyNFN3Cc58BQ7idcJ4c/kFJjdv58d2SnUueyl2oTQz08ao0xb
yoJl5uy2CqfSM2i08FxhNpsh0ULoiVScafoieKrL3k7GZTrtLOQcvqh8tkktOQEy
LHoeu10Y1LJl/eUB/eqmLLjljkzghOtK1CD0tK53uDN2wBrL/JGN8jmIq8ao3k2W
Waix6E+U1GuWoPYds7emHyCNvIffFL1VDLJwTwesYomPmiCZ5tzA7Wz3orsXT3DX
Sj5hUbOBV6qf0FA40UcNlJFydI6jbO9MizeUT3FObOgKkTmcpfh8lCsZO1QUHONk
4L8XgKoj4aJxnHon8A7G+lol4sw3fzzElz+L6lRk4MoICEW7VDaRI8w3HJsCxlLK
O2Stvq1Jx9lXre0lAKUaEPF7TCyQdS+W7LUMqv4JqWoC7u4WgGgkwsiw9Oopm9Oy
K5xnW2+43ULvvD4ro9T0BAat0Or25Dvo6eykrwrjWz29uza2rCm7PyslWk3WHner
uvxD+1Hl5Grjusn1rKsgKo7La0XXtRk4E+F37c6dQXobnpDNVw/v+WHH/LuZctbO
pIR5usMWx4L0hLHEmRPb7wHZJb2q/Er3lQ7I7CkPjAfmHf+gOTFF2CkGu0g7fKNV
5HOILK5Kg0h3GJHrv8Unq2OYytWZDbha93zdK+kM8N6AbUFrCfQnJyiKo1ZU/11g
A2hKQYz8HjIl5f2n0JmklbF50+sRImO1HUcbl2lV+52XV/zPvXf/1lC+/DNfgq6o
Ud9TdjNw/HTZR4H01CgTAJ5tLEct562F1uMU5mtctmdeW31UxMZUB7p5J0f3pnpW
SGh3aFYtNrHGuvqlgfLEedjW22wIFSLaQJet09yOpJVfIQhwPKhPM2bMIqL/Lnaf
UZ9+5DnWQc9vRakb4XT9ytRWZ8bqh9JgkYakAC9vVmVlAaOHRohCatXkv1ycTOLG
54IHJkLwcMc9XHbxnQ48C8F+SbBPToEUlZ1PagSSQlGnhJn+9e0rakAJHThQgKgu
BLXmsKoYdx8pdnMxgVlsqGk6ytHf5k8PcVxVgLzroAQk10hjQ+XFwJD03E1BVB7h
GEsUpJ1/yA0RO74IK3opYQLXGeTbq91o3BbpV7bL7NgmTqpU8pnVyCRCyGYGvG1v
XxzC9j1/9ngte5St67iVUbJYryGr//npUgQXtnb9bI2qzVufFOdGQ8k/SMkJUS7Y
1/12Wo/mfsCFt9twchVV8QhDwY2HAIhIJnnCfSykUh/sKK/gKImgycQIzKMOCPFM
7rxAD2iGqc2loQRPyzdcVd+n7u35hh5sPq688FoHlx6sjdzWfpqOCOnZya9mk2B8
BxOhuxDo2tcuiIv39N222ZGsuE5mLyNnbqaPGU7W+lilQvPancCtJ+7e/XnaJT5H
Hj9BFT+mvvbgXTEfSEOT4IbH26qrnTjzY3ALpYA1svKK7PdCLhWWl0yI8UrGVHbp
cxhaAyxUzvatyxh4clTBNm7BJ3X6MYQv4i5JmoxEYqV1y+X8/qJH3dw/CwxdcXTb
iVmybruZXkkBQ2PF9eG93IoNJ+e4uzV10Ewor8RYd7KqtkBgDDk+h7zteftQvjYU
VbSGvVTRjYyu/ImMk1wiiF2D99quxNx5vM+3qmcUm9gyK4cR+wYwCd5bnmEoncKM
6oHQDz+rmjCD+HHBvjiRterYMmTU85Oq4lc0wmNtVHO5APNKKK7q3Py3Yq2yRQvR
pZLM4OLZAbM5DmdIvbb7U5ULR0E2reMFDhM4LjE7k7bX68kVZMpD2Rr9AZGdrrso
2g0gVrguYg7DeyYM6ZbY7AOrPxJv8aEOF+drpyngHC4Xm0+eLeZI6CQuv2RVq2XB
cgk4fw4RzvDsL0uyS8zFpYUppsPu+vLV1pVAwbyWNvZJI4IUzYQ0nOC4eEEEa+Mj
CxO6gC1QKk8N7DdMzbkHsQk5q6iv7EQnOCym2yUOSC/IE1PoiTMvC7ejK4lctMTS
XpfSPYRuhVl5BAtDIBlgtYzQ4hb9nvzyD/EyBy0iycC2BvnZi3FqJT+TN2rCypVx
l727S/3vScCYjzyEI4nDFuD5Y7BFb24ZoYmhs1iYKdBRlRGWygRieqCoXySZb9Ip
0rfXYX0RrMVZ+fAjhDRV5R1lyWXpHcw1G1vbdT6IjIaMU9J6pR/W+BoQg7aE5xly
1tkXExNbhJ0tUAx26yXv2mh1wHDBh/5EdQgtIZ7C60DKD00PmDZAPD8Ege857fyM
O/nFG/79YcT5UUjCL2MeEHeI5hSS+LMB/oXQifYXplx2CUgFqhD497c4Tco14dXa
bI4w+kL8M9iYSwAo2ngtSQ+DzE1x4qn8U/sioAuqcw29cHxq5y+RzI6NQLMYcilb
NtiOG5sYLq2pO+GxClnhfZ8E6zWsiNx9IACKrRCym1QhZWSnJ1eW8ZImPzoAb9ev
5PpxCTpVypjLt1a93ZaFxOu3wogg1EpsfScVK2JlYKMGrQdtQMgc/EfJSaZaLVWV
TWANNdH+Fbaz/P40XhRQTylXyM76ODKX5ey6W13w2sHHZ1ui0DJTTWlx0sDbI66W
ZvJf+ojTt8BnEhxSl3CWLJ90BWvP33gaFR59i8rFXNoi24C81eYTVESuwmNVXAWM
PBd16Pb/gxQuAtrxk/JnCzJQREqEDy7Zjd4UZUVgxhnHyX2+lyTOmeM7Stic1sQ6
5EffVzIphBNXQGa7RhYmOVRbB2Uhj4h/eTZmux3ZfRAiKYQfZw9AV6+6xOcz59Wx
YlCa6oiNtH7mcbXkDlUFXDCTHd6DhPzQrRGLtNLiswStSL0fsYyl70uDIcP2UMl8
nixxj/JVxl4ockehSuLW1nFxL5nlE3ZaG+qSTt/g5K5owGLwRoNxyl6Bn6CgqGqU
oGCYJr/bdj038jk2choSritCspUuBC/Mn4HNPTMDgLARjV6AXkgMy0dTuS5uByLb
ZsRBWw7LzB/Kz/5apbjqG4UMV3OKKHvu/kaZ/cNyHGh4phszFlWW6I2U1orJxNyR
0d7aiLSjUUHh3XejasRVW8wr68+63gs2Yo3PCOgIIBvbwOWyAi6XRChWSHpVLCtb
lwBF66lJbosC9NgQD3Xha0CgGf0Wd9g/wxkiFAs5kO8zBc5kiUjDrXTzpBZlxTew
dZ1Qp5YSNkuRfnnT8NaddaF5Tye9at8yG68QP/13UWRZSJySb9JNw34PimYBXetq
/BVHp7afQFS4P7+RIwLmuYEXBHzCqUynJkgarjfMnzivIQE/FONOIFe2GfLtdcey
CnvjWeVDs6XTS7tIBUt8wWYDfZCtapT/a8j9LO2tPP4KOU0MxcBVj/QB6h0ZiiQ4
brV81iO1lnuJlMDBS8MMj7gyrTiJO9Ixr07l+eIaewqQGn/gxr1WyDt0WQWbrhm3
Dvs/3eAar6Tw+bX6RvYSEp9E+k1wDiiuMY+U6ZoWmoJ0U8QC0vQDAfyfnqClgDU7
1tLMcNaFkROSmWU1FycfMGw6EIwWCSCXGJc1ZrJCN21+4uHAM07ABZiVoJbPPXzW
2HMsp9vsZ7V1cW9bKHbfRT4K68sar7u02MTm4xHM80ChJMKPP/M8t6EaHA0QWQqo
OkZadfQuig07zKj0y+foV8fKVn6qtZLmjcUEWKCM1QwzksEGFIrmRqdEz6GVyx5K
7t0fGXp3EwJfaHE2NI8+U1lO6zVLgCOibfMvH4KJ10hhDq3H0ezcf6Hplz1so9dx
grlJJsxd9NLe1JwvOHWOhcLej5tOQq7GQSXS2AsMGc4eLIJalO8+eAyi1j4bNhfP
CtZonPQsecQcDSIOrTAHexDFV94mvGhWy+Qlmc1nnlbs0OmKlD536G2at1hklGPM
4g58F4LNtLAXh4elzlHncyM6QC4be0h3M2mMvTLE8IjFGaxct4U0K7fmO7JzDhkB
DxSj2exZAr0IeTWdZdRuBTmtaXFpb8/IkiVHTahO6AxsdWGT6Bda6X+2DvSS8FWF
GUJcBLlORhP22Resp727JOmcmEwstdMfTIb3O9DFQz+XfnQosRJzUgGluIpTc+W3
Q3OqRk6L8AfHFvBMW7UGm5e4SjcefG6xcxO2rpdkmPCsrvEiMB5Cl1+VveKmqdu2
13QmnjBlLKe1IE755M3fvMVSMG6LDgbmiK1RRbFhu0LiOxdiYjnJZCJsQGobrLnV
ky0v3vSsRERy2xZWpp1aEIM9NfFWOMEBCEgPs5qxsnMdCNS7n5/D/8j8/gRui/HM
kpld8yvKGvItO+4ovQHdfwKU8RAM36ulySgfUhrpMU/KXssUv1vu7ApFUKM7p0cv
qSE3x2no0t83h9i8YaeIHVR6nunfN4N39Mr404yZI2bKmMBJGawP3MRp2sPoXDXk
z8BJ7vkBFpb8Jn/2EqKR8VsONusa9W4sGZuV02yuhuxt34EwenJ9mgBYZj2GuIeH
2fiMKSlSptZzVtrXQKPG5DNrdrRRlrNXE6G0rRRYTckMVhFds0qkoaAlBAwtAgu+
OET/U2kdfiI4rByFhPFHzFCFA+UZbCp7iyFhhAXPLV2aGNQ8+yp6vAFIp6FSmITE
eUSp3CXZU5kfYrUU0lRkg90BJtNBAMaQ8LLGhk+SdCSfZc0kOwAbfUBGp9kdEW9i
k8F/YjWj2dktaIU7PqjxYfhtb+2PRId596hMVjdEdGuU2030q3MZ44Fp4tHrhyjq
XlKVZlfBJ3g7mmI6///z1KwaPJckL7CV1CfAO2HfK2sVxWidFuZdpUV/1fo3PPfF
5d3hH7wjlJ65saNbr4Vx2pIRb+mnZVKPfDyLZzhzgbv3Pkgxwqv972QKuOVtlo1I
8IiMyN4ifucINZTDEztS/0kTJiuvdzsBtiEHwLxmJosEp+fh38i6rQltPHr3Y5CM
mT3MDqUBC11E/EMhyH4cuIpvaIYeSab+eTTWbXLpwzwS/Lzq/iZA1m3Vnvgrgh+3
ttHaKOtc+xMJGjLxza05JHO577zeHbZsxWU0sqNuMJWGTFPsPz/MZaxuDwgibKX/
o8UPK62Zfgyi6r2w1ojdlXVA3Vj+OOzUD55dTnFDGXGmrQN81efv4qGktHqfDyQJ
c/BWdE5Zx/vOv4Ze3cGCmgx9iaC9ckblCMLBQApHcs69VOFCh7c5gwpvfFGi1mUu
7K4hQy1YBC/pBFqvKP1E9C31Rvdk6ctL0ZDthu4qggNt/BIN7b5TiSguWOISC2+/
voUiidHRfu/hVUb3eb3xMVAvH5wb9+5X3ijQvRvcU2VxLTBhC5SQDpX318J3y8BF
ZYkMClXIIljbkNdgnpzw5n0yGiqC84zj2zUiK3J0rTHDdIo5bUkpcrlDXQcVbDWH
SYOTqJ50T0gb+JzJp9hnq7xl6lOI2I+qc2lNX/FjVazMM6V5XWixwMTZ4J3jiLr8
OABwcqg+FDc4GXqmzcLsvQ0zld4sNfiMhQ3QH+cqfWkNrpDfG4d+Y39pljGZTixG
nSB93Lt8gWLUeApVle3I75XeGGayOkqjwMRrLI8BN4jljYBcl78LQmGyhYHDq/fl
nvvZrNgsf6wkD7eiEqmdhzD/dRnXocDVRGmWPlOdIHA6H7ojaebyx+EfFcmquqH2
ZEBd2T64Cm7eykogxrFU0OHwgoKbsxdHJMs0xYwE/6GmpgXlAc9XJdJPMArVrzJO
+6Pqrr6Cjqr1cRnmv/S8sjOFj/8GWUmZ+fbL3Chwmk6NV4nJc5KzPXNkDaOW6LRk
LXDeQoPZ6k8SYAq9JGZi017pOHnQ7V6wE7Wg2qc1llCBN7ktAZqJAcRqmhfALpsH
t/+mUJPKIhwzQgD+M9IJxqsEfjTst5Dvr+FakAmy9mwPLsL21w5fUIhaxmlO88RI
S2+n/EHxSuBozZheJ+przR5hszWL8l54HUWMDu7BsZsnSkmWaXQZsYXFrVgvn8bv
cXoaIp5BnPIT5tEKSAl79daZV8DjlHmLluFV3kJrUti1bBKC5pmryvN94WEH+bRi
cQtnMGZ58K2wKguSw+ugO0hyIWbKPO10NCZF/0O3vRVXhOnTJX+bznjKZRMg+sKK
jRJojxA98HH9PLCTWdorCXyH8eB1bqMn8Fmii33N4112EA/DQ6KkF8nUQ0AhmtNL
Xs7jEhGbxhrEc8VC47oZcYTNolwJPrfAfW5cmgIYJT/i/4Y2uWyKtPntqzCnI3EJ
qYIsaZXKzebUpm1u4Np9yT/Do90YckusQxj3chrx3JJWGKiiyd0k2LgHPZ5GjSsb
6BGmXtFjTkC/RoPdLY98gSQ7aBShLkxp5pNO7uVJBTX6JAYf2FvurmvTw00eSYZ4
SWXoeMMRmBVW9LhLrxYey20E5x3wuOYVedpMOe0HxYtjuEWlVWwdhHa72rKMjJlk
16X1K00xU7vlc8Iixs09y9/87Tyd2AhmHX1R1z5qNKK/laiY9yNnvnk0BcdRdSYd
4yMD8Fifo9+K8PhkJig02puQVMvlx6ORcodHUnQJDmplAFobgemCQgjoFOYvGCaS
GtudeOWzHoFG5bqUhQSQy1nb/UL4s5nDh/+zzxtQXcV/5k+zxPjR9JVdlOngJMnY
U2c1ZitNm0ijUG6yphbIHoE+Q78EBfFW/G+9DAr2rqGMBU00eOOIFe7+aJWtHueE
9A9SMAtyJF3DUcJJ3PVeLsdt9l/T4bKLkTMxVDRL/eB9XpRr6DxRGqeJOcdM7fQd
2GdJmMh1EoIqLlCxmju0EnKuatesRKy7AjOxfucb4g777vZLuY18e7gzW4gWpTjT
TbOmuUioQOFtwsauissctiPLAuhmB4jcVeF2O8MLh7m/DChK9uqOHMk8lWLGtIDz
EhDvaHzvEhAfG8oeZGF+cJdTjkHGzums3nVr7zZxFMcdQuAuLdoa2R0jIY6tKc9T
jadaiQF5qRE7X4ZSgWODee1LQ184bCAQQupfYFiP030fcfdfVcc+sM5O16yblDjA
xH2fJ5UeYM0IN2UnQWfTg3VqXD8seRIibzRhMNZFLjfmFFD6Vx5xuzBtfuOGXftY
FY2831DmF8hLT0o3NVTMpQSzTVd24vHGMGte7DqTO952GqflHCAI6e1hNT6puZBr
R0lYaJ5MAjQITqHG+YtTj16NJ3qfTcUwjsXvsCpJIcnv9SvTdY2jZa4htSHk4zvs
2GlDwUNApmNb9mG6+26ZWxYcF8fCjB7QOYTREhP/Ecey4eEMYd9PMYNQqXGukqVx
dhT1ZCRjy+mt1L6Loc1Q+rUhhG0IvYiJqDDM2xo2I3ec8V6ZkQcHjCizQaSb/UUB
IxpPjAzyonl6jnT5EvUYa5E46YDg4sky/ymKqtKzYcxF8NOWpclX9IihokAao5Sr
5Ub3j9VnJn2iLXtdL6WqvTVTqviqR6aEGRs54RPRP+KIYbGh113nI/sOROMpNsWC
V73vzseaMSWmLm0KKpJPXwFX7aSpbFm+qybb3/OhnNC2jClqgLfPOYqgCvUZnNfb
QxsMlxn5+MIo8sxqLsm02VLAM7kumEZez3Xl3SRCT27WFFDqVv24NPziNeEuAZ37
ALdFHxVnX8vLn0B3q4GPvOyuySD9vC45KROxh6WaWAVXDJcOD1FyJgqxvlbhMvLn
2Daseh8QtXaMQ8OcgH/UgUjTh9Sw9F1ezG1lRLQMySt+CargFjkQip+18GJg7HKG
uDCxZvVTRR3WsKavEdBCH0W6fKrGkYDV2Na/17gaBngOEsoRIZY+QOBTedVTXpGc
b+38PgwYAhikpfCYHEacvNH6iSk8h5WOe+IbfuDTzr/rszY3fihtRSmbkmwTKlfF
tbLSHbSlm1mUuOk50T9WSAD6pDjSSbsM8ZfYeoSPFdofKUuAaap5f0uf4soAn1Kh
QbiWx+6NrSsXkojYocJS3YqwLgsLd4qubjXyTamUk8P0JYlUaW12xjpI+6oL1Qg2
D3nGeA5f+h55QSRQpcwUMz5E9O41KH5h3lzLYsWUebpswIKCr8mdWy2owJ70ZYZh
Q2FIXRcDCyz3DXQznCS51qar8Lg5fgE+zfOmGn7gR70Uv3WSCkcRxTyxHdFPQoVS
V/HLY/LaKg7pArB8RTzg0muBonkkvmbwibGPIQic6NJ+icxjEneeIpV2uRX/7dtu
rCH6upSRfDog7TpD4BOXfQv5zMltBVsaR5ojt0z7XkXqjh5m0BrdE4EUUJQ8qnza
GHlSyt9PHUPq/dFym8f7S76p3RtcmR7USmWxNhIOISJ5UVMMar13yrWi4jWFW13E
W1RFeCbxgDRYdf8SMcY/vxQVtA6jrc2ypVuu+8ahCjVyQHowGH6cg2/7BPz6kEsz
cIf2cFsPo7hqzy1eN1QRM5+DtqcrsMn6fKbCi4ebCi8Xfp/91CKxDTiRIOMsYZuf
MfRfPHGjgKyBPZ5YlEJj0JDvBh98DNETEPlyoZJFPsyIBuSXtUlTDnLUWBoeWv/m
KlI1CBNKiXCmeefeunlqOdyAjQ9aHiK3UkUYU4I/MShLqX8R6Js4TTMsGJhbknEm
aY1JiIjaXpjCRO2w5cs/6sd4XHkiO6aA79a0xxbP9iXrDmt/BuVpcHHiYV6xPURm
y0D9N7gYocUgyNCBqooU63zGrO8JmSTF/n7BbrDet73OPjw4RHbCJ6OlFrhvzc1/
lv4WVfuIGTtJrR490MpeV2dcM1nJX4Y44doUwe4dcHFphk7qmhUYXvW9WeA9bcts
sUoe2+gLwxECduvbSxBONoWKH7brsqhQ2EfaK7cOMYoDbUVYg2llwVxCrWC2r9ta
xyG9prJXFyxr/6Itxf7rJY2V4PH4xgMvBLw4sG+nPydNIR2PYzc5ZifqjFWmW05e
LFGz2cNdjwcs4tRJhN3V1V+0LFTX2TlTVWwyadSdhH/+/a4sM/bvYJFw05V+GeVK
3QrNdCrcuRsKlER+qLLJvKOVQ2OfQlA+Ga6c20NolJMfTE8BISGVq4jv7kzcf7Bn
pQkA3+Rjvuy+dDCNzmSfEBAAMm8eEQ0zY5MgB24RqOcVhLlplR59fFhgw8P4EB1E
Fh0Rx02a60jVXvF7oEzz7YQVflFRWXV/v96YsHym5HF0pZYut2Sq8152hS2XsPAe
e51jP488cu+/zh4lYzIvmNX75ukG6pe0tU3o/86/L/GQAU+IOURds3wgzs4Fr/rU
d5Vde6vI7QjR8TlCW8pUpbUK3anLs99ckPPejuVZS3M2faT5Rnhu76QTWbtgNKFD
94DXaSWgkwZKLRu3adFO1DXxqLThOrom1lBiZugP5m9sC39qYOdgefBH0LizHYcZ
jbXJrrpBtxABeUDNVblE7JNMgv290MW5UYtmyjVrz6hXYHdnVKAZq7Ell00M+1IA
/PyyLMT5QEWDPZS2LDutdM7Klgbm0Glx0J6TWk8S39hij0uvVZUb1MwOoZ3mXi99
J14YP2K6xiWfROrTITLIsD4061TuwDAvgjk6Z5YkMmJdhZEuOTaI6QewkSCCygD9
EnEtSt5Tyw8H70yZkpHo9SV3dGu6moo6cvG+sTpCqR+WPMwIPru6FjnIdCbgBFzV
+q9jL89dyJzTf3Xfisq3G25sGNJm87ZB1lXufS/g+m/QzTrkX7YI86tPb5h5z7Sy
93+TqqpI4xGHRhiKAsvDQ1OzgzasvNbNxF3RxHUPPHtV8Onp+8h1aKtxH0+3ZzYE
/Ey9RCYrSkhVEp+Hw4KakpEYuutdr23bRfZgJ5f/x+B9L6eydDymMCGD4yGhmBxW
io73XKIrh0lkWnRlPtRaSmt+a0tyRJwl+11797TExxEQnQvvQl1aHIFTGEFsIS8x
iyhu/QLDmzigRCBVqFrosKUt84Pa3an/Eq/d/SKtZPpiosD5KnVs7GoqjyphgwTE
3cirBN1Zu1X2UNwZjrQdQdS+0ySuLVmcIXGg4wd+DbE3BgqZk3ALQDgpyJ1QrLJ0
Tq2pVxkesTgoDuCh5gd/rq8QK27/XXx84ed2awcEYHjD1X7B7c6YYCBqiuK4Mk3q
xFWRKATn5CFRgRJxbhJ8r1jdhqe3pC3HefV+Ml+ZRJG7I0jccIwXJHUuYsGjQeGd
c/lm4lEfxPahWJIfUVSixVbFF1MjvWshpWvhwFB+aZ259eZHDFFtVoH+c4iSRb2i
q8RzQBJTOkBz9iS8YIVtbV7Nv2dc4TjexaFWCzcp/NPweSFnSVfxV69nZih9KAYi
/oq+GMPnbkMKWt00dZrjnNIGTpK+D/2eyYerroSX/MlNOKQhQIYnA3mDmflZ8M+s
e/AOvfVOu8uVhzeQyhm5toKFWcrPn5nMLb61OOK99PmtORiA4KFmruGNn38wIaVJ
b4PkumhIxtQjAdRcRj3+DY08eP5anJK48e4DunWXl3tHBCGNH7jRgGjn00ZE9Nv3
RzoJCPiOF7dLDqzjVzgoWI2b+UI26LP/VFvTXle1KgsaAURcgWpkSahySi4T0B7h
FXDX0WSnY4B2dIH3jAYFnvpZQJtuDsnvMMDz56Y8ClezzaFTAFfBrZurTSReNC+Y
Sdzh6q3RQSc2I+OhKq7bjUw2fxwIkPtiuvI9bqzqhfxxdI5fbQVy4XNcTIBH/b2H
UMs2fyouNu/52X+UPiK+lHBBuXC4BAPp89NxPINIPI7BJFqrqRRULyXl/eRd5RVX
zai580VC15CcGZFfBBwzQhS55LvSIlqt8ZusGBc/IR2j1Z9CvGlaR5D/+i9/bOpP
hDx3rins5RJird/MrYIYaxUEwqcLV1ZxXdSaQB8uAPF3FAgDXWiU5djxbL44jpZD
9KCPB6c2DoeNTRBD3oOmUaLXemnZQ1BYfcmuct50mxnQb0ZUVw9OuI9NaAWzmkly
qtNiWwg5emttZ0Mqtp0gkKLF+PG8hpglqGOFDVlEFjPWpUMls+t0tsnhShNVLINm
fmki2XRaTHd3xvAB7ZugsA++4xFN8fwTyku3jRiPrjLNk/9m6Y5QRMOzYXi3ehVr
b7sP/uSDNVC4pGIqLlllU9AGu0Nz0Fz+2qSoL8SkGZi5twXH9kKERvSHkQ+RRalG
3iwEBXuhSKzeZpEP+uUmy0Aig+xwZ6n4oOo0uoVxkwTjFRtv0aoU5BY4dyId3F5N
HHB/PBUOXWb+p664fkfOZtwNyfxs9Y9PlxlE66oRn7fnJ1e/IaHMphhzFaIXAyH4
5Glw3iZ4Hdwlgsgsqm+f+D40M9rRfubAn7U+fOp0th9UKIi9vWSiuxN6KDXLcvEd
C8gPUIlL9xwa66ytMz2Kl/X0G+QkeKbb1/pGtmKQTWczDAMwlqzC9ScNfBDQGvAr
IeNT2Jnoj07adEgem2bHn1zhDDpJZnOo7IXMWe+Xn2QwE0H2+LBX3A3W7O5Ss/tL
DbxZrt5e4EUAMOepj3MtXnfFTaPRCJuAmApan6bg7P9eslO0liUN6ZbV0KcnUFN1
1HXZ2JeuqHQkkh4zaq0//O+9tuQbSmnaKk6fiT3EQNsm/JAVOAz0tkElgoKUOZgA
/83FEk3brCqugKC9y38W2WkzWSmr4ggiyUGUiXRoMBdY+u6AKnposF5AUBHnVVWs
89MG6IwGXoJXEYKuGxlBes+f1oMzVXuqdtquDypXTtpfbadEhNnENgu5DVSV3UXG
yTs5KLovnjLkiAqLZZaU7vw2K7I6pjylJ9/lydRSEyZc3Mz2KzgfnRZKTKTFKABO
L3yanuTkL8+i0a9i4ltuw1mOx3ZertAZe0Qd569N9DtAALYpEo0a7aO3TV+T58Rt
wwWBRk/6On5owvJsd999F95zj1NOPdp1LK2uXciUu+epSwLZwD8wwXNV/5RRpcQv
qk9y0zT7QrqbNNLWJzehEqTP/kwXg6fsBw9m8W6O7Z3QO62PmHe+7TNB85Rvz31/
Sx8mM/6USPCWEznE8l4REW1t/oPkUIcJpkOlNkG8NjmdPQND1DK8ZdpGp97eaz3b
l84H0RPn4klEQdVTsDyB0PG9sOYzEgM1h8ty821TeqB3ayzrMOJOCqwdFP5SAVvB
6kCcD4r6CF3jM3WvMXeIZI2qc2uEjRbGeo3NRzn+bLrZwgO2z4zVQX5v+JHjSdDg
GwDrQbz3QR+K1ewGp1YO5BtocdfLB2Zv+SJlp9PggsaoLbhnEQsWjqNDLKXJeR18
BWwcZWOGAYwmy5ZbnvuEMryeCw1SIvmLMLgLTIWzb2H57IX7AwMwWcvc1d9LwwT3
nSe0mdta7u/m56boI/8/3SRV+cwrMm8W0XJZw9hcFLX3rP0gAq/SXUMIcQSigiZX
3eK8WsIfkrbNdd4Jx38Soz3oPaUrU2NbnCbzlDhnwmp5mmibjMlWTllDW+Oa0bkz
FkdOOFzzBUTHlRPYY8tHrwUYIjqQhVDyWhMMqtaa20AXXD1drHUAsXt4uSeamUmF
6Tw387ajCJgk3GytAOdKx0IsxgkTwNLewUZdgfazbb5wu4J/BJClZdwoGGqyxwrs
1gLq5gpFdOY4h6bqNrD1I3+dpxExKcygL3awaldlvnWQt5H7zIqcA6B1eXLvubZH
HteFZvCwaU/ZV3Ft0lzoSgah+TCRI+0HczxYTJdKD0R0hs59sU7Izy0P2CR0GZYP
3Z29cFvTHov9qctjqbwwIZZQ3azwPYbq4vRrqg5dn1ZrqAiijiK4f5HTTqal3OeK
0TJMMqIMsWXF4HTAskHNSAAJ5x0qnOHRIwPj29iej1j5QVhvSvIm9/eeqVkuPLvh
j0SwJNGaSTdZdEDnlIcWE7DNX0eYiEmGeVc7Hrc8Z2fUswLJY9yNzSeaPYtZCQSj
bLe8z2xIHUnl5bdTrYMgC/CmV0WsWk+oCUjBD6HyylglBXjm3H7ZIF4yylnbM6jy
EZQgFaRGteA/EFRz0YCVt4+lyKz5DHc1/eb86r+0940pWNpudC4ilruwDWvcKRf9
sz8lLMdsC8Sp5Q1wL/c5GzWBVwICHYcz+T+H+wdrtvGAVbUO7PPcvIzX80fKnqBs
gmzXagfLDYpEyf9DHcy8cIZOfljnrjopbDdHAltKGq08SQEM/ul3KtT0bNQdVb8p
KSy+Q2TuwWki/6t7nCFTvyzS7J/cW/w1um0JepqU5OG4RNu0nnOeVLto4nfQ+Mj6
BYOSk+2I3Fptvk9xd2IP1qELuwNbCAIu49TMBRLFLX5LxvKL46PVKcfVhQZounyO
OuiKLZIIjimrIUarU2RgYmPmYStD7qEd+GiKT/yMXeAtmP9r4+/JfCQsYEQkKIz3
dzKfpDiZ+ufSQoVEehjAKKvi/MzGL450Vouao+2HK69jZCx6R4jv0VEwcztW/bjx
LuGUogIpTvkwrTWPQUNix5uywvznafjR+FnQz2WBJbaEgk/QDYQIJcrlRw2pGHB4
+qDg5EFbL/smt67Sl9dchZuiF/1WM0gh+yEe4YPlS779Nia4Jhs8nbXy1CNYE9YO
IgZcA3k7H4N4rDaC/eQOZ+xFZBMJLHFuh6oFuf8b428B42wGyfwTeTWmokXxJuV9
uKBJRyYjITdJxZqBNi5jEsmuSwpXf44P7roKanBZC5+iZaIiifyEPu+8aJXe98wx
+lZZMFjWhpZdo7iUxD7Sg/dWFlcRVssgFbaz7MLOgnxeCTSe87AFDWEHxyA7prkx
fkrIth4eM63KdgwldrnCbGmVzFC3oPhFKawbRcaw4CQlBuOrtgRHJq/JaN5U2R4F
KKvQFq4s9JO/0Lc4nVDtBIo0F6KflwHyK+9pdzDIJCCIJJyk2VJTIAFL/c2wwfoB
+YB/6k23KalhxQUz0kSIcrvwKoDKDC7JcEvgeSnlGZaxAk52u2MSCY6A0izsVs2f
575UHzMsFhcL+xv+00FNV0iRvp7BhNrLCX2YxNGUH/quG2FrJcSFamI0om0Z8ClP
OuDVKad+Bx+knaHA1jz+Xzgo1DR9dAdYkqLXBvG4SDQknb3PPLZIkGAIe50ddWM6
VO4qMeEH/bwB31H3mSCUpuppN8FRRQkfvcqeBOgo7LVjEGZNKg68HI78si9awyuq
UNrmtcYUx9GPU/mz7q+pCPZDnztR+yO7/RbFWuoJ8VOYYPiF/qrYrc7SIom7nLR3
LYXitClQ3BhvsUS4EO+CpLwdKCutvZ4EjNakVdud+SXQGXPmUlVarH0e4j7M/1/o
E9xGfLtW5wVsx9hug6FkFbIo17Fwfk8/nl1DsJPdYiI78MRtTuUv6U3E24W/BuG0
KRwDVwEqKdKdogyqswXLC+XTThPNE8fo7v84iMKInJVU/+xTx3mfTAIFgb3ki1lm
C4dS+3zMASaEaq0UvEYX1heMb+ccaErF/Ae2YasBhXj6kfyAo+0It3QqLe/YYcmt
m82wFn8BM4LVTz5mZ/T/eftboGQR7kugnVpgliE+iaOtpYwbvkWlfvvitqnRLjE8
4pkR1q+XHwT9HYnBfbxRh8vvox8bazOxc7k/osGhvBrcgO21G2caaXWBvctv4gWy
cL9aSxEWB/QOY3nBDq9MKqlftKCoY2nqwFgJz9fzPJtuQP8LUfwoS+eBlReK0CGR
p9w2hahfbNhD8LR7F/pLLZzUgUMqRd7Boz4t27FSViLYiAFCgVA2R7XnZ5h9Dzz0
P5FXQaOu99xg01EmUtffHRnH1whhfaPj4rE3IGIoPFKYA0KkFCX/NixmGwPe3Czq
/RYcpe7bpFqkFmn9bJUdF+pHVYeL0VSRRzF6M3Wn14mwCEvVJt/NIwOy25IOb76D
QVdwwfA34XQBi3jgpy3EJwlmEKdLB0n/WtvXI0VmKxn3zAPrNqq0E5TrNAmqvQVA
Dxutvh3kwkAbUEo21j2ngudwwtvRVqMw1dYgKLusf7g2Z+m1gKQqgDrb/OpBvy3l
NHuGh2dq31JuFl656DQzSnozC7YzYhM40QzhAm9LW3n2JomYz3DiRfQXYmofSMXE
T23R7IXI+dhPTVpPAfc42zrbI1eSKaoV2Oe8ZrwYfySV93JbUjyzcwfbbjGNqxh/
XYdAz7c0cpC7zCmHvebO2xKB3OHRFRiCHUXVYH9TX68V5i3veXgyzYBH9/ke2Ffg
cTsAkEcAJLMQgsDndr8NAwBGw9znwgKvGP11MlrlIIvL7OaPmGYFYNjUeWRg1x0I
sNsJ+XKTbXcDIeKZ5do1ZlgE01Hak/upayCDzpREWmjHfsU017eNKgV7F2NYBFkB
Vg0Wnq5BGGpOTycHIPEcqvRbu2KmDWz5Uw596Xc2gYrMXQ0H1cFw+KwzqH8iCakH
iAvU8gGjVAQUxbZmwPfEEIBdcbDeZHEQzRqff+q5o3KLGeBDQrHhz5WTK5Ehkv9T
UzyvlDCarNP4xV9Qq+90D3OnG2TZXpl2MUgpkM3hcIUoSPdBnoWlfgeCc6uNCft0
71nZ6qu6PC60qxxUywHpPI5R9VyNEN5jA7g6e4npgc8Ztg3M1RALRP6GmsDFa5bh
fKSF8T/ResdF281Gy0cf2kQBfRnMOPH1fzoZuif1mj4w86bWMPqzi9wAQHjmMFi5
YMoseC0lmScoSsZOyaWUmn+datO5qZvzttaz6FPqLQhy5Ss6duger04xLGEbr7tK
Wp+PcDtEwBdk3ypRx1XzDZdNQbXcXIUJHht+IxVUSNGMJRt5/+RiwfXe7Troi1gU
ycIV2eQ8W6Hde/LQHq8a5ygicn0U8Cwf9LfW1xQ6G6xGXoN9VU/cWpxe/S609kkM
xDWwKzEBPlPfwQTxJSpKinP74ChCufNjDUhX5+Ob4QUKwOxl4H9Ji8f9Dl3nRKEG
rY1xyecfX0C5pOPu1OkA8rV7AR+0QTbes5BXkYgN/5xloQPVfl3Yrc+8vmeurdp0
5gyS0r304GbKnORvIiK/LfKb75j+j4IY1PbKPi485dBKMKygUQRyKoJGeXVhpple
hm58U/foxMcHnZBlPMNAP4PpgUJgNb/py+dgS+KgW2t5aou9XLjP3s2idkBj98tJ
pvPoBtotbCvLZJOkp6RShDSxc6QW6+3iJ7OZZODT6hg3wEy3iLxTzpbXXYAHhpjF
ncrwTpbYm9dqrZScOd59ItLNTufe5wV9/Re2Hv/T7/J7u99WWoQiZ/lb5dqD2pwt
m1fl78WscvqZHjHtApz0aTX1ZCJv+Tw5Hij9J+zA3hu2DiqRYAdNRJQ/vLZwqAJX
4nvo/M8Q4US1XUF+/gc41AeRVLb/Wtm/kaFp/44JN39UZqO2NL9eLK2KJ4wQ2jIe
hax7AP5qL3i5WRb2g3orihPgFh4pBIhNkxDL6IJQJFh5i4nT1Y4ApxV9EjQpOgm6
1HQzwGPgEGxI4rTMbEW+oUE4/z1Ze9Zp+kujK49zzYdwZveRFV5eXmwBvUrSR94p
fOPONkHzS6WYkmmwBbv3q38wB+oz/Ja4pnfH4xBZPSf0rZy/0WJidwgsmW+8fL+p
5sjJhr8dxIVLEh0kkmVLPpxe6gjhCplqpsnXXektew5/2y8RXBXZwW2L7gchaD0S
XXBRcDbpJGwWlYI3Ha7Wg5cN6Y7upb3lFJTDVOcBxxmDal7nYBgaUkZ34g6zGg1o
GRLLrtBt941eyqik/HZVjXylLosmMUDmf5MaGQGIIq4LtlVR8PBdiB37nCEpBK6Q
NORsXTKaHMtf9SsYneplo5LDLO4Ha5BQPlenJ4wHEy0nEzWIibqWxI4zsrVFdjFS
xGU7hKt/aYh7sPLN7RRwvt4pKQ9x33KB+CAQs3kIzwkqsHFTpcIf4YPTjayXcHLz
8cpTmgac7W7SjlKVEWcsQU/iq1WkwBxzkbWFPxrwXPzkKN9lQOWrHJj1Q/fovjTO
Cc9hHskL9wB7GEGIVbCGudOnyagV5fWfaXdg2ByRyq1veUqU0c6MlDTeEXlBBf9w
zncDY4f63oNS1H/Innp/OjT9XiJYcFk4PgBFS2o0aVyNdBtPgz/9gc8DvUZTL2qq
iEhNicOSuj08SyTWP8954PC+0rQ7iB0tQHrQd9p62YmuN7bP4lnbr1nkwxP0p6WO
kaTfsA2kuLsba3C57CAbHqKDh51YfirgFMpJcj2FJG4biuY8rvoPhSPCzzKjx/nY
b1V60CqfO0eIM7g0CL06jSpGXH9KHeqtlbzKrgRjs8KNUTewE9rZbOBDyCBUAg6X
rtkwAZsI1QlaxO2OlwsfjH3NDl2qGQb4xAtxesDALK/1Ar0dVTXY4sIZyqt2P8R5
ASE6Gjj0/h2gPCZvjgGlmHJMiXF4gRANmPhSGHl6aG6lv8Shu9IS+IKNBPaSdlay
wzOWMUL892UDRQNLZPOhocrVG7D5GbBro2CHrHacIsx4k+P4cAktt3NV4oBL6PSr
dy5WMDFiIoF0LrUOqAJDwRl9uV+8bUgFPH9lflNezFqS8/mZKgW6nk3eESXuRyw1
nvI0eYUsf5CDF2c3AOjuFQ3yTUhbNFu00iYyI6MHRbEFRS3pl0Pa6nsxiEAvQZ68
XJJzvbOeWyCfhE/sfO6MFgAwHXyAmDLfI/I5vyRuiEgAAEX669ff44Me0/55LT/T
HB7aiyT5/+b7zhcJaDklVltsEsYQ8/0giXHXK2JcquCSyuHzQa8ZyjAC95arH+GA
hwp1tZ4j3vWXhjDZH0DCncJ62wzITutHCbIVFOV/5v/BCK9tMjAVP0FLu5C7bflH
tcMvqWvtIyL98Z8ZPX1ThXgUWGQnjfcrFWsYZsjurhivS3z9PLUNRjIMF9S+jdiL
xIr4B36CCnbQQgAeze9kGER0yCcQ4QHm+TBzD5OP+TvEK7dXJuiiEZ5TjBOnPGPu
YfA9Q0GfP7Yb/l4ub6KTu8knOqR76d/wkNzmypd2m1no2lVJ3JpDNZc0aT45IeQZ
R+TI6bsRGumNF1OhYXp7AbX+hS1l2IvTl0FVq1I3tAfSuNDmlOfpT7tVlveAjtKG
d+lpOCYR+X9d3G6OGBzObggsbV5jubzcYexDqfx9cwWWDAgstUjDvBkjbxLTdtLk
ZhFRyK2dwjb0UeTQhC5Fz4epnwiZoUBkcjNqSxUHKS88jGODUb9+AWysbWFLMCPu
5S4wzGd474Tc2w29XHErheR1xdJUwLOyqnBfB+aI4sQNBcByFyWiPa2Mspoc0yur
s2msj5gIl0nrpQrdyj/blbKAQi5/wdju1ArOLGVoB9F3qTwKfKHkxn+godEg4zib
8pgX1Td6PCZmXVZNoueIzG1hA1jgAW0lp7u6n5rLJ8Tfg4PN/BIvWAkla0sOmcne
18NC21+lYtA/XYPk+9FUjFeFr8odtOtI1eQjKOcHTl/SbH17WCMyoJIZ5Mkk4L8q
Y+NS55wOpJH8oHQXppyOpyqL5EilvK19icCgn2A5Kn/+NMwXbUxzqUAkzaTjFVd+
JwXHVIilSgjQm2xWWTIGyqyRQN49QoAVBQ2q4eWXEb2MlBgLVLALXQC9+NBREERa
t9m/hAxMvqt/+vsvau1wYvskBZKLaXwhLRsRKrRf9PWSL//uLn0LqPbsltom7XYJ
PY02UjPjTTI0mBLgginGsQPDmjIOIaHsFg2UZUbCvEuXo1AEUwYDmf6mZ3qgmXHR
V1uvMwSwRl+ZWTuhX0fskFkuJ90B8a0Hv4AyjqdISiK8UK51OV2Tif/WduocvMOL
L60ayCAgrWDh/66kBGlDE9UtCUVUUtAWP1YM5n7zodgOE4FqgscMipnUOziXl933
YV6rCKxnJ7bh77zn6v+F6ahtpcQ+xecOTg/cO67KSOUTcwwT5eXfmIWfrXpdxujL
Po5PiVVX6GkYy9fRJxR0Wqj0ZVUGKNhZsV7409EuHa+pc/dr18Z4B/GSPMhyypYf
RFDY7FLcDYOVbo9irsI1nZ2AzK0oRFcBMOjKLGE6+e+sdguXqmETXo18IGvUsL/F
eJ+TYejUKa8GFi2olcxBn5ZGw4sIwp5oMJy5f9fKGFU9kQrrchv4wY5cjiBlKajZ
qH+cU38LTmLGhT9sfi5U3MmGVXDA9G6eVMrb/3JozxYX6IOEEVH3PzR0MOJblJ1E
J1H3XZRF58jw+QkiasGHtD8YufYMRAkT5Nf9Xw7QNRgzfqfwQTespaEliQj0nRjb
hFmToAEvCQyckSShCjQjpGGQJXIWa/Juoxaxj9SOxWbDx7z0qfxnxjOJvUOv2due
ayoc1PRQ0brKPEnrbU5XLHJ67RPWJvIfRGupYtEfMUwybJ4w8DctXco7KBqWMS23
tGzpq6DTM/oAjx86iruu9Pi6gMVe6BzzakGFfB1I8SdJ98tLk/lEjVOU/Ird4JII
4ovRfthss0qTwBVevcBxUL1NP6dwpeaHAmfKTxVTwjVSmWUf5y9PXNtXFMqZSmHM
qqvTXtaNo30NslB6779GwXvXWAnfDzYRQ2ClgSJcgfscs3zFSnupU2c4JK0zhWIE
IyaFl8d5Dp0NtLb6D4fiQbESPVL5zusEaty8FR1Dga0NXeUQ/KKcLVkTeMMNtQI2
XgSKJ1MADtqYp7LJnaz7C3DzBWlisAY2hc5z3ddpeGlzKhWU8Qy7IcVywCKEa4SU
TKuot4epME6xPd46B66xGHTzc1FzP2Nm5tCnbPaeHo/d78XGH6w9M4g9xBypIDHx
jSQo8y9+aw/v42+G2nUmy+d/u1iVVueTB98P+h6BhJZqysp/5gGnak2BiuBA6lt8
SWiarxx+7tREHQJYxjLlVWl7E83hipf0T6QY8boG8EeWPX6EeeYzUunQoKnnmQhx
QGF/76vFMD4AWh7lSQuPC5xXzRShWnfddaabFOR8NBhDOVAc87O63wbCOODMI+9z
v9B6ma4lMm/I5JmK8xIOgBdtBnXXvgqEKKiB9q5dT/09b+mreRPg2Ny5oOl8yBka
ezfZ91+ERO/bKu0snxJc/c0OIxIpobI/obYtm+stgbtAPgVh3ple3JM7LXX0ggYe
MiLBtsDFR+sKWOLe4OPhINdIRTuBJdXZm3Z1ZhPSzD5CuSEAdGlnaCD7qAt2ozTh
aCCWyBCpciP471p9yqYD6N65KZnkUOJvZFyw1kk6mm9xd0cKBFUzt9HM9D6qrpXE
XpWjNbJNCz7hGdmTmI5b3K08NsWMsXaEbvlU0Uffzwlry1+qq8aKHnBTTSHST1HI
7exvXmrLUpGQfRWLKBIRbohzItP8UKYz3PcwMAXKEJXosdqrJh0JXb57xzt1/F70
cuC27ARPoJ48xq31LNJLUSZvBOykeIPs7ga6yFK2XHLLsQXIYPiLRJOd743XK9B8
AJEp83HMZdWSPgkiH4Gy/uvfv3VnR/oslCWUrHpBsTcemfOzp42c6bgyl5kZmdJI
yBQ18WfAJyW3A4hku6NkslhqsrjxGFG8DlLVF5464INXGmlE9eq8RKNjMVAqeRXM
Z2JU6CcTt1IUCLqmL9UpIbYUTUcRogWhbEifOcPYHq1Xu95dTFo2F+V5BHQNaqCT
WK6d7L9DnUIBNqyAX0A2f1LIp7N+a5V3IwMTPlJp1B8EhinTVNJXI4Hi1QDni1y+
y4pZ1DdvEh+fSppbXko/ViXJg3y9ZRnbD/9lWkWwnh561/d2iwJvwT8OpgtW/fnI
lkeNEJvnpXqpw3bUL9Jh/LF6HJJ3r1YBt7nLC8RT+MnFZBT7smSbbN1yA/U0x4iX
15yIDS2u77l4cjlSEMoK4TjuoG2E25umiN10VKrdVDp09dG/1p1X+OxRw9ALchP6
eEyx2+Y+ZxFRFLuQ77hLj5UBtct3ZaJCXWFFnWu1BgyH2eiqWclo+pQZt4LkQwxe
2aGaadn4rcbQu0Kq/ae+rmAaVXt0d2gglD69M/DqHg9Ms2BVLYamNiJuDUhG2EEC
WHbd/xNfVmXzrPdOiVzP8jaiJZr9qzXmANwejZAO7AP/VbOAb3/K5Lpy3BF2B8Q+
0GOia3CM9/yr6EfL7pqkim7T/J/k5AKWX/Tzau+kchsQnN5Vtd5MSlyzgJARCgzK
MtGdsF7ueX/cHnbEh2FlQenUk191s59lKR787MRGCWfhN8Q+F4dbZPlk0euV+O78
VQu5k8nT8iKcBr6YXceCmmp+ePXO20GBVxIT2RN6Em64WtMakeqBNWjTwVkVbBf1
C9yXCyKD3VPDcSwH3dj5C0KRVE6UkuSL7y0UYf1ZKv1SFuZfXRHpTItC4DmpyKE/
PzsPSJIlazjMIjZAUjoXbWTXtZfomX5fjk8mFn8/8G9IczJx6uunD9BPNRCM767c
m6WBXP6JsMqJ9qMvKaJnUUMDR7BV82ll+TmgxCWPDb6dv6IMMuprx6msRgeBhwJT
e+7zMwGKvec8ykCCznsj+n06Ikic/Hj+VVM3I3fQpFcgDRdew+WTYBZrH1rZxNZg
Vw5Sdlul+JhokZ7rToiGQ4R0vs5yacLMMzHsIL6KSA/VW3Yd6PvBvYSJqYjYNOzw
gpsjY+AisHuAz2b994MaRmMPJqQuQmv4vH5HdMfo0g2RDbYtuRg8RmgqE+z6nnou
kjYhSjf7YYz19rA986FeJuwAzqG/QPNNmADWOnzHWaX6VuPYVpI3pEd7EImJjkcn
Y41fb7KkKqIK/yE6MYv7zT4nd3TwR5mIU1DNCul+HOV7pCglFMOyqFC6N0bTfxXE
Ynxb6wT5cE12zRVseSaIZ5DDvd5Ks5l2EqNeTBMchthuhhlE4xOeLnaXc38ga7dV
jCgIK9CFdWyFhdeafiLWTEd4DpPP/hjzvop44D4lH9Ypxz9977NL+Qkh1b49NGZX
fYHMFd5wkVpzWhHPsQ+iXXWH6nsknXaetgNmeF8Dr3BYsbMcVLWLwH6h1w0Guq/v
h4sdqMjMl4HeFZuSThfLPfcOByq17jf4i1vs23Lz0WYN+orNxeLnyh9iZQ4gMcsm
8Tp7IPGeuQWd3ClpDsKJYn8oZodPyds6Si6/EapQVNnxRLWXBpOjupOsov83jupp
yfxTp73uIMSChn29MTkxWKT8kgzCqqlO/8YNXAxSbP2TfvtaTkPBQDYA8sXdcGHB
Za4UgLMF+RaxfldYFXo6BHaojIjzev+nAc0uQzzNAKXtNhxD8L1DZm2QDMd8xLU+
ByRLh05tuTfii/dYiL6HzzzewgFCcyouf7F+48poFk9qXLDXNHUYqzVCbivN6SQF
FGDpEP/6/Ly4tVA9XOvzuq3HMbaoY4WF4aPmpTOP1cxMpa/KDOnm4Q77VjLFCAcf
qcOQ0i8moDC2s7xplJ3QAmxZBQ6sGvCRICoYWRnP4VMX1BWYerqxJWdgypcfIf06
O29r28bolRc58TYhg41N2QonV5qCIhPAVAWjlx0Ww7zLs5OZ31f3fC/lj72r2Ngd
i2+HrDAwLnenQA8COOnyvmcCHyEWjpYf9y2is3h+2uAlrRpWxFBAbqy3Cj3bDwPK
IguIULXEA2KYRctJ8WWOzte0IRVIEoi+ai4S/vMA5XXDN6lm0ikxbHqL+yMShPnu
Q6hBwRK1DeVn6bWvy4Sqo7bTrAg+86hR9klRvHFHEAazk7ZaIM7vomCmSyvcVb8x
u/tF051DLnyYGkjvX5kBK/8Ouzvot9G75hoflI2Lz4yQNeYLzTTK3+u6Z54ByTA2
fUAEqYaZq/+GwV6y60AnIetITXGEnUMyifsweuqfBPrL9QEe5Uqzba1Oxgm0aBmJ
41ZRdcIOeXBFh2Lu7kTXzX9fZ5/WYfDsYJ/XmKfOBQtSMymQM/371OGsm9QlmXdP
m0NL/s3CjVbWKmzaFXn6K2QMkVAw2ggEhHjyrd7nZ2E+65VQFHyeBrF9ik7TLAHv
Ccdhv984uvXenCu3AQgFbrFyNcfQ9MAdGs7GWzWVvsrhWnif2xBqkfNjm6bqRtgn
oei4AARBtF8UYd9ffbZ+BrmcWHZth/V0lSGPlWA/xLxsIzAHhO64qkHEeGFmCPGd
+bUi/s5Wd2BenvwWngQ52UUEmkA8ubfhOVDSfRx8DQjLrHikYWoYnx8915w5jPKo
+FAHNINOmqONam0ObVrpj5x6UF2xrC3RRwfSiAU6PHmxKxB+e2yvr5qWe7DGByvM
EX/P9O+jkFkatwv+r/EcqHPlyNlQudoUPtIc+kzVtW1EKLXuVM3xN1YA+Bv55v40
e5e9AXVY2YwZbs7PrgKQAF4TjgA8SdEWTdokmRqWzhaF4l1WNKIZkzQYHX+NgHIZ
OKdlmknLEYlNcWyz/QzQW9PdIz3EgZslano4AzBZzkOEXNA/t4sxR6eGIwqadgHO
66o15x2YOWKDy2768zteAJne66JnN8kKd3lZ3XGsjf7yeaS6SQjesfNOMVk9+DKB
uN7fp1wY3/rPJB4En5jzeE++PEuxO1H9eVMfKOegCqrlugkCrFhoBCyMUN7djDMq
S8afPsjZudYwa0eWismB5xmrdsBJz/c0mKajP9M4YYTk7V1RmLRo597rUATNcFAQ
cFSVT8HXTy4PoGEb4rJK4bmezr06mKZHIlh+QfN14uVRxWB3d20pYvHrJE3+Z+R5
W6dDN2qSo2M/DaKjWMKGsk7iLuJ8C+yu0a+hkS161kzUnpdM/NmlIp4zXxi7sFVp
PFsci+fxKwTEcdzGxGqZZGXFpL7d7Xmr6lKNocnmh9wO9e3iV2UW8MqZGWBpci1f
j86kC1NAq0+AAgEPsILHEHTM/OIfGCzS+CPoEBb7CV7Wg+KOBktWBbkY6NEUqguu
kqyZT19cwKKX063GJXaKR9B23M1IGvZXm7fIZvLmBPerOEFDKhzOIGELDSMOW6H5
S1gWwvrYGK1bnTkuQ5pve70l0ikLzrU8rlmEjGeLFzCkD/xv5gzhGFob+zYXMyRy
wH+mxtuc07b7cjJyRyGqvX/FG3tg1KTbB3+yJQDRNjEX+uNN3AM/oENgn+rt7xfm
ul+HKkXpTkL4/K8+HOl8ccpTyLcRD6QTqdgOzRiHnTLsqt5hfjE6jDC4OGa9sFuY
DBvbxzDB2K+eBnVcoKk45RzTWdy6USTbFXf3rhc95T5XP6JsF+ix6Rzna+myITHf
YpfUPfZYUfEH9ugW44cd9E/B3mzSH73O/owF/zXH998KhpJvNSk2xmfoCCsBnclD
mNmT3hT7sxaa8QZHqkLVT51EEhnDlfm5hE3BjVczb81hTFZbT22W7PAxdcOmenG+
eOKyIDJ5WLJFOy+IgWDHcrTtl3orViwYY0uhcc3lLMhP3Hhj32vImLt9imTAy7r1
aIJWGH/EckpBYcwgI2yzCxEdAasV3S3O/tXirVr0HSQdmj0YUIfL2wqiPvDYkFWd
8feUoKwEBfrgUFktPQsZwik/2rbG5S6ZAtnpe2C+FqwQep3ZDwH4JE1ypMa/2Evd
XZ7UAeGIRRZZjkgCx/dnEB/2FzqMofchVNC2ZCljLUx7mGnGddHRMwwTEuTHWLHW
OPyVcwhDydUsAZhKWAEhzQWhn2mm82ghvC2X4CPBEH2g4TLfMlRs6GF96vzkMxKY
vb0DLUpZvS1UwA3bNXBZ3ZZ21ejRiyzh7uNvuFIcsjgkXJBSxCWVxny5zBu5EAPC
jswNq8uCA5eZwZNdwbAcx2fUlTl8vut1WEvFoQQ2c2+Hogy/b0zYUNWZy66XhBSh
WoYjwFJKpF8ULool24QJiYynGje/4c/sHrMorSgjmy483aUKh1rkKSFqdrb3FBCA
JNYGSIQBfWo2SdcKWJ+VRehepCzJ9TGmaHevDYfjbEwEj6fcOhnTzB853zMTecFo
Ufpv7advS8I7peiCWBwk9+aeVB2vi7JrCE1s2D8rW1sjmCkvZHsiQnYfWegiAQ1s
iOaBXBdbUt503mzkgKEMTU2ifMpcTUJAqQTBCiSDZ/ggZTQ+SLs+cOCHgRqy2u0X
tCjCsClXcf5rTWPxKRnAoJr8u+s15Ty7kLh2DpjKOz2QaHrvzU34Pnf95Dv475mo
xSRgw83dPnslj5ctgyRlb0EjoMfRWSljLPc5zhj4VajU8KgEP0Gk6Hpl1EBvOtD0
+r42x+HHXsoEPrYoNX0sc0yu0ZKOOD4mzrlA+3h4tmp/T8O5MSI+BXX3A3vaRNdz
0hPzdYQ+PgJ1QmLC/XBBKb8xTqXquRX06198rHgN687esXlM0Z9XGNTyupBqO18J
oely/w9B0rrm8ODBKf0G+qMdch4ADwMO3hccnMEGmybsseNVusJm8sKP3c3VSLIg
yFqKan2YZnVg9Z2O3voQJVcdmXJAiZqnE45FcjBaLESixgvzSrIilYxyQmyl7WYe
/EZIZCcJFsroASC5emv6wlhPF8mHrmU9+D/GOZLyWFLUOf4RtjVv90zsPWMUftWL
GTPn+1hueaNxMgZQyPlW4d6YSVRqE/Sb1az1X6VJZuo8ZKZ4PXjzp9e0q2c8eK1i
Kcq7OhBvLWScwkidgdPx0oPyhgOkxWxfXC63GE4cVpuXIjN6e7VqD0MrrseT09L9
1+ptAKs8SFbab4yw6+Q4ABD1mwxhnJgxRzF2oqog3SpKZB7xg6w9ziDbElMwfXo1
TjY5e48sJcH/HkP8R5pLPgpwVBrk4lNNu892slYNI1n3EDPKKD6VRqv39Ng1QspD
wjQHx0dLEQHuQA/ovwqtqv0FfG2Fm5exm0DeC5T/VGJAuQkNprSPpTdVxtMkdB3w
bYSlMPPxmFP9SKwkfwlhElNUUdy7nMCrudJFtyjJktj26l0cntmcd0k9i0s2z/6r
lGnYhwTu5JYakW1fI3LA8HWLgQxy7eDu1fSqWY0tzljnfIFWdfBm/oLHGGD0aFpW
eBVWydjWwICt/jYn8EnxUdKqSrUeXkKJxB5/oWJ2kB05IZhowqjuI4Jct9vC0WX5
FdkRdeSQUpjB0+rb7xQ8Oo20S49VLAtEb9yqzqPBZajI3tbOlJLbmsmayG1ewoGz
OE5nIws2DNmExTeu04djNuBvVNgOKGi6zOjGv2QRNJWo7220OgsvyMRGQ9UbxYED
0vzcb7p5BIWpnBHNNqCIv6z838hrTkFPAcGDjZ8pH+CEkn7Hi0Qkild6Pi/LTH35
1dTKvY4drJo/v7ddEjoLlYUQflCXCsQPS4E6PcGs1RSxkPUb8kAs+l7CFG/fqXJ3
DueccU1mEmmROb5wtDCvqsAjrjhl8uyVbx2SnzCIBgxZ3vKrWSDIUTSwXwmMblHh
vMdXbiyKSUmn6iadpzCMFuIoX9NJtiHVx6PugBYCt1YmRo9WtQpf2bBC6q13w3uE
+tUIVvTTK1f18aTWylIy6zAae79fZ4j9ntNqKGP0Uzzjef3im0+gyRWcAex0Xq2x
C+wT/361zXVSxwP8qMbOeOYpzFCM2aLGNsPjfJCUt5yiMd6aH/mESj8XCt1K9ZIe
teePneEt3pxppq9JWtVIi01cIDG6tM7LfQFQP/6WeFbJJe7Vdo9eN2iVoMvjxFW6
KsXoTE0QittJUMZzbldIBtC1fAeURs0ISUTp6dUeERKB9TdeHkHcFQV3X7CYldPb
cHOR5c67/8OVvrn39l53F6++TE+YtScqTLFmtd1vwF0usMPANgeZ9LwYPEv8/EgU
VTcQMyBoW9XHg2sM6LPHA98fRO3DgRCf1JfwJTgMiIqzcyVd9DsKq4JTayOrdnvm
zHNl6zTxfRt+bNRBRb6hvW6m2IfixybX/t2ePhCevT36WPe+4dTa393sS46kvXvk
0gry1kR0UNHzbDGR/HKse714PWsRXpIQISVkZ82z/44j9efVQB7JTH4zdlfmCazi
d9ejF91vZclvuu8KdLlqUa3XHQ+5/nRgycYcwRu/Fw/ztoOSCnAdNveXPyrcX0CY
Wi/4j86l7WwhxrpiWd+obyTr0yG6lMRAgo1ZT/CUE4xgHfrF+oQw++mzpB1l122r
9Len6sTF9nQLwYOfse4j4hl01f8LUC/eJFNJ2/GUmjYyBU4hZ2L3V8NBq/50r5yG
yrO+BdrQR9l7MraJF8bIk7MsbDr/kkEWjO6oL52ash5tOUN/3J+wVlAIeIZP5eE2
q6udVXqOZ+yD/EtIcj/t0RrnSl+TJCr0nh7wcWBgHZ6diyBHHdBLCaaW+RzkhVrn
Ndf6aOOYdNaU1+zqe3o5zzsc8hsqQoT83IkmIyZsl81ALH17CTlKQ1LM/eiSAy0K
yDOnG/LFrqu6B/fKM2urUfIW3O3/8KHrg3bfEPzPL4XzDXZjsUoQA9og0+7/gX6R
ZG6PWeVynWrVW0tIGs8USlhky7OJnc8CqXuRhRbLga84QzAg+8txtpvI+5DDcnP1
2HGNQaimTN6rjF6hjBbD8dJ9zWwEWeWAx2qk4V0/F+S6tSwX05qlAHyil94/qsbd
HNcJWopT97dhmglg7cDsWQAQ9WuUDqB9wre+zBOaw2j9QXygVDxuAr0uo/v1wwP6
jWFZVFlRrmEfiBXEp3OGa0oYpkLlT9tF473rzr0u8tvIFLeI6Eii7KxSvPZn69t1
fWDTe9AApIptFCfY9o9EdMyF4gYdyiPNvopex9fxTNgVqlPnPDLDaqsMU9P3wlrk
IzaOEo2MlFpyY8aYjrZIam09/fp0YK+PAJ49wBeOwv6npLpNBdzRpu/XYjCO+Ck4
238gBKfgKS60eCp8zum8/tu8mSeK5zbX3zKbYCFeDj8EITJiUmV6IX/nTi+UdL7c
t62OXUpo+a93jiEjX0mKmpQUXw+Iz4cjYtxdH76kDefvZUWyGTA3UAaKijcSAqEx
AmBdFECEBDU+z1c2Tho/E6uvj93+Cn8fnuAYvOO1MKjNSKmbEkxCnCkilF/XXhll
A8j6dLOiXPOe6XYFcjIpeuEco4Ya6fXe7+6EV0ovaUdkv/pe+eVyqbe2QjQOx9jj
rzBOaua2Zhee/DLiLZDSsM3WyxXEd4vUa8pMaP3FMDaozggn/m+cRjpyfjsY4b6h
Qqh0dpuaJbZ4QIbZUaK110KXwoazSr1aT0LV3YINSVg6lLu6PDp1vXrZ+M0LDkKV
GExE+Ho23Ixpx3ZAsXXfCKJWUH7wJTyeJz633UYmTISMBT97GrnWv6A61TAC3Ndc
OGaei4uDmfDOrJ0wuBqxBf4Bu3fsxMLzVb0WPnIUYiZFH6sVqsqvdAY9bg+0qv5v
3bfzOq0Lv+cJYZtkL+LzEKtFieycPUPOXar5kB/BEYu3d+fFU/TXVpDQ1PYTmfyF
o3xjVs0McZUmWTbwQuRjLAD77iv8jw88Fl20VFHZcS+SWNfP7SXx0k3JESebWamH
Yj5hKSsNwbAzBaNtxj3IoxJwXsdXA8rEIbCJPhVgeFR6x5yr3qNShW2YGPprtGm8
wN3UKA4j38UhX5M7YAH14JximkH70xC3gceSALLeK3sw/ojx16C0fnnPit8gf34k
m48rqP5mEI6XwqkX8+2pfLIpU+evv0JKyISCfrPIEcMmirX8L1w8hJTtxyvBhNys
l3Uoa43X702Atyt/5/bcfk7e4mIjLiWqAZc9Ke7+ttmpsBeTKhTm/mhXsfYidxpR
Var7LYlLyQextyFwYt2EWcXJRzq9S64E5bDqEXrEBMAQiabVpEw5U62dzenmZSLQ
ivHSwLoEuO1Y+ipXs9nf+NnUqnarNUZhF+jdOOVRxSBiGYS6MJlXPOrin8sTTbiW
luDQQMuxj5buAjAK9v+UX7B46/H91Jyzpp7nSGHE6WrLMWAk6tduMg5xwAsvJaMt
sLLNizBAgglcKAIuglEJWf/+zxj8i20hA/Q6H+7PDfvzBJTLH5o2LA1PxTF8p+Hl
fWokVBx+uDWDmE9RlowG33cvmZ5aomKsQb4ie8gKblC+NnTWxCO1YehPmwVentNx
wBrxcR73kBe4+xnj1Yf3ejcJw2xh2+sURgllTZlq5lc8uV+vQ5GOXn2ScpH7UfOc
TZzKzBDtcb3odkfOnJ3VHYSoDmzBifVZSikhVkOjrksPAVYoDvfQg2kcDxiGF8mG
D/gRDjgMukR6VhwWTG5KbclEK2L5Y1KPuUg+6AIvgs40ok2FgFolrHTJiAdPr67r
Y628STT42ITR1ey3o2TKOvaRU0w6maUjhW1QG0gTPC2brh9/K5mbHTr/BiIw0t4g
doC0SmJh7B36FkRb2gMFPT+OFbwu261VvQU4I9gyQWFbSm76/6W9JuVTgTRdQW2u
KftJJCPZIZsziMuXLseQ1fPXQaVriQM2SoYzGbk7WnsgfBkPJF/tFkbzPh5bHEdG
xXZZ7tLVoxzTm2EJvUgrAqE7hCcAsQhKYF0lX7H8hlgeZJjqm4X47D9ZPVQ+Hi9u
3otPjG5Ddot196DciiX2Ij6sBjfedBWn8PlMZOjL5n/lKipBhGrecx0sttMOxT8X
RK7w+iY5YxMTm6Z/hd79LvAY2vHf/95NPiBtK4JvzaNu7LnxpkPi8c/mgrZCQfB5
OUVV+d15hCL6rnoSvHXyDm96G/WLW2zdBNZKdxmH/coZYOvdBvpTJk4LITCZfs9Q
9r8fAAMa/X5Hi3fwZksB3yK61naD46jXQ8ONktwR2Mdm0Uie0f16/HJk7nlYLrrh
PoNVCIIVd1o9VSzFdtIYKBb/nktVUCmTxNnf9q26Fxn2ORWisN0cV2SbXmMfs1/t
5URu931SJnKjXE7kCZ/XhcyadZSmTyPnU50EqfmK9tcHazvItsjJmAFWC0taNc86
nZYu+ah4dBlm07qo9qEv7T3QsIzcSM4w66NK3cysctXwfltSBbibYcLLeruykwPV
exELSiwt/6EGl0DiHRehDk1kGgCJkO9VgB0GEpCC+eZSSaPBMxCinD/LadM+GLdw
0YpfIXkB7oSUV7VzIo8lKhIWMhXRVHyqFPEKgKmzULKNUbdJpYe4h9D+phi94Df1
sftdBqNE+HcKLtb2FA2CP+FF8Crg1DsOm5t7ZZa+7XA/CCljvP2JH80QCwR3w189
0hZ7vq8lJMrb4dupsHRk9zD/dBXGtbaPWdgkxGnw4OQoRpZtL6+17VjUO+xZWrL8
QbRS1JW4XF670ftaGlFFBueZbqHYL7L8l46+urCXcEle2N1greqjiy9aUCAHeT5Z
Go5KWirfjiZelZmPRteQj5vvsPLhLEXyA4+u56i2e1SQj6eUN1fEi5gW+4gJbbg7
T/BOT2dDWwKWtbV4VmYLHHNpEoqUq51Fq5Ivde6N4ACCsUq9qzFfMScBIQxG7OVN
LUXMQm3USNvhUeyQodsH3MRIA+f+fVxOOmkhDg0fd7wZarUSkqyImRnX8BwD4AKb
yoUbxdl26WnDNlsCT7DF1OQEdOxxYzJB1Jyxj2UW0ZyTNpI1aBBVT1zxofpuDxCQ
3Wqs7djITmAXf8yI8DowQZv4c9UlaKJyVHrzbfoihT/Z8CouSnmLpD7cBO49Gg29
0gb8k5VFxGkAQtCccjLfYT1STINmSQ2o1OG8J60k1p7uUyAXSPUdE4/XKesT7Jo+
gg3r1/J6QkDsW2ogtwFllaLJAwFhmlbpXauDBspbpTJmmPqfpf0lHRDOdIFZL+qi
Q+NnE6xl13WTTVDWR9qQ8oZ0X4UXD3ORiMRx5NN0hvZpCCn3JuKDk3oa3M3v4Blx
kjSev88T79dmrJtQmJvlMTov0gxFSHhd8cvzkuN8YZRP2rx0eZD2Ap/iWsukCOlC
7oix+NBTPFlGnROOnVKgrYIgs2Mf3zvFhlKzRc3CulYxp6bjUhu4IkksQcM1NnaV
06yhse1qNULdLS75fibAS+nTyEKiuc8oXd1R+tlv7YJ42A59xcqSyH1omV/VYFJO
7kPD/+INvxC3+CuGRAUT+ka3UcttmGy/lk9kfxetPg8iHMhHD55+rEf1kgP6ysHP
cTWFpjjU+kU8SGa9gKRxvKDot819z6lrEXZ+Tc/ctBv79/udMkpBmTOCV1y4Wuur
ODgX4t4/dxiQbs/yhxomx8GJvayDgoq6bWAhtdYl8zaalL0s+4lW8PClCnDrwG0I
WtC8qYaKoJXk1Y7voO6X2tJ2iOTVbkIyFueQDSc3xiO5/pKym82wUVkVNg3szxm6
ahIwW/qm7jVzo7Iga2GeleKKnsKQeAtGBuXhYmfnjhvhm1031XOSiv9iE7qZ0eEh
plu2pbn/PWD1VRWygWOpvJIbzv6jg45XLSNlyzleSrRhYjXqXeih4cu1ezlf2/eY
oAgqV9lumB73AeEsS4c08Kwt5IQj4FYCY9DDHvGIlSpjNPHTQKULx7/AkHN+lnpw
Z33XJ0I+V6KQhrCFyCPyZCD+XcAsj2n9Jv7lnLlCD8ennqtLEiUulZGD3rNIlHuG
w2yr5qkI4D5covsjVIUr5+WMN/N/kGgHliHDFIRQc9ZwsqFdE9k1FfCTEXin/3tu
UBzoj+NjW0IRruBaKsKHsjP7AHOMwUOLZ/SwtRPDh3S58VDbCVtSOSpBBfd4j2yI
9/iJY5PkPsrHGvSncFXmhB7LYxOmNixiXRnb4KLxIhT3h5qQtY1K65YXXZP9KHRa
mGyMRRb38Mj5mtrs+MIMnMEa/U/vTWB+puCkl5D0id/aMAjXBVEF10QAjtHScO/O
D7M0S30QMKSRs3XfJd7rgaPt69KPAKHhXVghyO9VJ64J0D3Ln8qtAwp1k/h//x+l
OnYSu+8drfGLHh4fFAZPshVwGV5UFshgEGkNe0jqPvVvjljowHPA9F5BlT8446IN
OdL93FBiaEKPd5I869H6C8ljoZTWKNqeBS1xDtgcVp5IWBkkEAQd8FDA66Zn3QWt
8rbYv11aHDxwk4LXctJ5vVW0C+ggWgSBb7b8Ty2iOrYGnAsIjNqOccGIAVrfz6Eo
iMEJNOKNEujYCcArkaUUAOEHiEqc8WCkvqkY+UYRuq3tclawyYUH/DvrOV0v2kFq
HxbhKeehXcf5ZJ49VHVjOzYSyN1QuliQ5RCgno/UfIoN32rMOnjp/FmAjzclgDd4
qgzhRp/artmWbIBeexDOc6l83OmCbhh+oBDRcn0XgFrhtsDOk1nd6C9E4kPPPtlx
ryPSNdueMXMmOm99ALf3y1hLPLWgD/i8xcmbZgQqHcJaNz83RH932bxzR+pa8J19
uUgYMDiFqWKx5KxZ4q4GlAqmEs0VktW9WtPye4IKKuG/ZkjzvBrhK++7Xp5aT6o2
Sf848JAJjAG1bJH4XPaui1/9UZM16rgYgtPWyUGEaekYb9Abd/hrLTAVAxmSWiGR
c5/KUu+qij/22kou62JujI90XkezLTmEZAYNf2xcPMTx0O8cME3CM+6tCTFW2Cnp
vkMdzuwMgD8VhWCREMibu5RpqhniXTxl0xBKXxsZpQjaLIF8sYAMntxrCPlBiWU1
gz4G9E6JJn4+5cUHB8BDuZGz3Z3twsO9wxD1tjxccXzVHpzmCRBGJrGFX3vuvOGt
LX60qmYKf4wcCZ3mTiCvlsZiFSy1ArPsyb4aRzKDA2+ZjOHLbZhOWjSJBO96eScQ
RJCMaq9UCrUKNTebUkJWr4jBqfdI1gMxH2RFN0XFZKZTghsJp9G6m9QbGQM0evkI
x/UmrBgvxGKI8DKRbbs307GbTASaqph7bqeK/GUvFktFg+jN7CGaz+/Sv/99++3P
v8HAeuEEZiaf5+CI4Pi6HgngOKYlnJ5z7UsyqYjvwB7s41N9ZAhfdiHLjq65XsMZ
XdHSp8hvz30WLPz/qDWRckE58kUFf/NEmU95T8yHDEvS213WGPYi2y3yBmdVeMRr
jYYC6cDSH5yhVr+9tg+NKUXphVOufR7+684zMfIq5CSL7Wj5yGNX50dphphHhYRQ
VFW26uv6h9YYM3aqMerBrPrCykyuKUDXU/HlETuRb08FCItyh/nnzwi/JGI+rQU5
vO1m+GRT9y982LsaZ8wHy4S3gnIKtJz4S1y3j25mOmO9tm/YQWvEFrIu5srebB2Y
ZMgdJj1I6NWsxLNdClGDswb/hAVImXyibW1rAKZvYpM8xEq7N1NIdL/7YtdD6/11
PjSOgGojLaM14kjWOHIFLwCwr7KtO9nfyngxC7s/ogIa8Wq+UI1dFV00FjpwFg5Z
uxHQM+15/Q995DniMKt42FUE3LSTW2goZ7w9vR7eQM4OvTSzu6bBfIazVl6e2mNQ
L/pnocF/kGZUGkSxm3ueutWL2AUv6jF0ylvartnhcoDGne/acmRRyy7uVJBL64Uy
EHhftHwi8GEvkOTts+SzcKKzerlvkkntMh86OLVNWM8sUSqf+ZeoPdZYK2oE0D1p
8PiuXA1Du2BfbVxG7SZD1yhWZB8OGUOI6ndRlrbZb7y9UlFHk2o3Uj1j5HsF3q7a
Jv42ECtEs9YqqEeIkbkgk+76wFSsv37AoGA9xVI6KJTir6oAY841UrE1M4Fcq5aF
uSEwPXG1RZ/0JVhFWVBeC8vbAaQmQYhUYE09HHf5fhW2cCgyGspuaUNEqecZMba1
YGokn7d5RaAU8SKbw9gte3NafyH4D58R4hAmgH5v+jdPzFLaexvl2y4421mcyPPH
hhYvVRYJTl9BVhmurAgWQPyhXLHWqHwBxrKiyJpyCCepoT6CITv+gDIXb9z7q7mX
I1FcPZcSEG58G1OYcM01ZILcDYe60Vpl8DoIzmqKzABBR6/qnxoRrrlwQFIfdQyd
aU0Cx8cZilBAc+Uat+pgBGNonM2qkbZ6B8cCIgmkCJnjJc8KGp11UGTKOy3kZZND
HxMzWPR71/Wgiif8ibeWWwTapO/LqCN/jglMauy+3K98QDUt8R+Y/vWKZifR5ypH
+P1oMV4bmM8RGRsW+5XTDvlBJ0PBLtVEpYJjMI1N0AgetuTbnAMrrizJM6uQm/Yd
bW+ov4Kpv05ZRyjISM+8uZqDE4f1Monuj99NGGmPOvTLXxunGPdI3JcWPZ7JaFo5
5Svs4tE9NqyU3P/yTLfIEj3l6epf3xFzzuimR11ucuSb5OlxQrdZMe4SE7yOQaDB
Unf71sNC24mwjbeiUrOEROnPcd4hDvktmXadbFoTw4AdVJ7Ew6TgFiX6+d2nE0Ch
mnBuQrt45CSaKgHFFXxDNOYLB5oImI9aujz5h7G0kuk2+O86u6gZNhJ2tVHLRB39
gukgrZh5Hxmlbyxsu9veTwtYy8IGwRhvcEQkjV1b68X1LCayuQPL3nYngFWk57tu
qqBZwAur16+ZfQ9qC8euMSBKHEWqMopivFkF1LC1erAZJ/ria77ZfhVXNzgvN2Um
ceTYDsxOzQuF2mYk6ikjbicQ/gitCnXYkBVvS/PItsBB2OXllhFWrMESj1d6JIH2
HlRubPkn3E0rfy+Ld17IOiTurmIkteKX1y6SrezEKKOzUurjWxe1m/O4z+UsX86b
NW/N0qjZN+X3Ypao4o6L7zLANrupR92YribNhJhvYsZxRlp9tpgPbFNDllmTxO4a
6aaV49DmZu8xSQe3xghIcF+9HPDFoZoiQZch1tsaHTf44W1neD64dMhR2yPEFmpM
c4V15ccjBRbnr5kAgMtcXpzIN5S55iDypbj9845pgKD4QaVIH68gjJ6+RZ5p0/Am
p81v1QTTbMm7IETT17UOOt8TWUZ5M7p3cCUsBGwKMJJjU02v9aVNddc2t+Lc2n+U
wIb6BgLpE5LLXcmbH+DLlgrJiwLGJJnf8WcHGPP4ehVVTVIN4DsKbLvES3zjNaMN
2D8KzTU/Sef/N/PIVhhJQ0qzIH8GbIl2gF58yJD5rBQ6LILQIVqk4U6+HK7WqEmN
oy6Nwo/0oAU64du/EdHoOavgjlPDTXBqNiVSq/CPrR1HO3/fLXAG4rHVsDAopZhD
CcZQYJpMUtMObL5cUhT+TGhYGQghuDGoPHkDRLhGnpBWqi9Zcaf7ccr1VpP3x7ls
RzB5tOqLqvOSuadswOPVOKEmloOjB3Is52/pcpvUA5WyEnrciuelX/ylLDxp5mvX
GEknedZXv3mogxJ1JGuXKJt9DXNEXwrKJPvR6fduy4GbaHosSVHSALG3+VEsYivm
1PG6HzL+NXH+I2godpSGsvpaadeAsQuJzcfZ/LbPAVrt4NdnU+Bd3Ipgc6HSjkZ1
Ozy6OgYpCoSUUREs7XXjov+a50hL+2pbnYCxDbRVRQs00iNvLFKfO2LqX45uQrL6
HyQ2J4b1+4VvIbvRPo9cj4qYUMXyxGR8zUabvqsbMidS7uCFOAqdMk4kf0YgWMqc
JW1/R334z1u2aIqtZfjMTYuiQbXQDP+vA3mSmbBR3qdKhNIATAbvA3QamWbQTG4h
JtYAneSFf7uuEP8bv/8QvWVlTsfSiGdxfZ9VBct1k5hDGEU5BkoFU2IdghJpSE2i
Aci0AMgkDwOZnJUHlbUiuvzh/8VhBkbKDQ9gtJTakMgm8gbaV1DdbZHMOXmH8iFQ
GGRVbqW15PHZjTzQfYCtqGSGleS9MbQ/C8IgPP5663vti033zrdU4k7v2/SdSRx5
SIVL7QVK7Tunwc/mqgdtj5L4KJJdGPHew+cujIz8VLo1fGm0STT5rnIOBHcCehcK
cFQFmVsBpcPhx79sbSrkEvVLllZDZ8Ab4KEXVjUsEIg4oO7DPoWscqTl+RRckXPy
+tS3+F3Ro32Bkm/pWwBYaeJ6DCVH7Xp7E1vCC3ethTT/2QCM4rh83vKI7we7Cjkc
0ZzU2ozOpqhNlmPq0a5l5KpMXwhSZRYVHuHxM63y2tCz9Ir6n+zy2XwNrpobzNdj
m/uA0YS88GDScpmvGSfjB/rVVBLHRabxG0U/0Yg9iaVNOkmKdtH9OWOx/Ido7LGP
N4OPGfg4vZRvMitPH0U3oo5bN0DkM/nYi/ZvnkzOrS93cy1qI5tP9BsqxMgs20VY
jHK8IQS6XWtGSeEvLCfePnnr4WfXmWmQgVqDcwES/Ss1yA1PFhU4ipr+RBuQyJbQ
r4nJqA+O+acLB1UPhwPu2LVJsuLw2ktNo9FT7laTOZNewp77Vt+o8nrH/SEhYDVx
TF76GU+A6qILTEtrMyr4DoJn0GDo9dmr4x1pc0yct6PDttGFMyR0vVeBmhXdqI2D
vUJklrarI+KNZhVSK7Q69vPpNjXmqgJfMYAZuGLg6wd92IoipoxrHUJ3WOfeNuw5
blYzCl94n/+dGn60MQl/mSho189FrkXw3gMzud/GWMLd26EyU1+SawrG1XlDVu07
POZX1ShHjp659fRlEzU9LMauVVWB50doygRv/TKXDjatn2CeDqlyPjifietCnSi1
tzSJVComZlTeRiwy/4cTqLLMNZOv+N6Hz1wMkppVYMISU1S5oynjUOiES0r8RZs1
LjScziQg331SGAk5GW6YwaYVxiMuQHrC/lrOV/DPrsiMxc3B33LyUOcz6/gKC3/e
u5NyS31vwg3dG12+GPPP9dB+yhD+HNF4R29ZrDY9JN5CUKf0ylq7E4wXhNKkjZsW
VBJ2WJ2RtVVzmP69+WHMwDrdIotTXVluPDA7LzLCjPOulS6pT4jM+mMV7t6GBsKv
6NhPp6raQHpfBcuAwfnNC2CnKqAWiHinM9tO3VD2Z+O+ZnxC+HAB8/cnMt2uwNMx
SwaODZlktO9l6Cxh2Vj/9PwFf6LjSOH/TcEGxyafhCNx2ccQ5W9aTIwvjheYaM5N
kewtbCxW7UEkMI8DPhdYpJEQJPJBzowVb8kdY63xMpFno5Ov2IwP7qIGgayLhsUd
QC6ev9jCCjgzZCrowAhDfKByZHM5hxfKU//IRRjNi25oKDchnHD112F0sIinsKg2
CBmB79jvYEnCSAvrNkjT9NQrGX2tqQfayRx8NvjNOZAIXJlDwJ7DttwvAbGEaE93
EoTuBjn8UsNLxVdA4TwI2fmBfYsx8KcnAssKToZVOXsvHYPSjWL7nFgLDtwqLV7g
Hbm7NiXtD9O5P6tKWI3L1kv9yF4VUOZ0MWaiLjc1adCV1mvoNrHAa8QbqLiRe0yo
m2JP9t6pYhuPC+QPEWi/zYmdiA5wdL1qYtDW//JBe2IE2P68qa3qrje8yEqUUJAk
pN4S/BKamA+5yVXvtP5FPfZE3vLBEA7IQXaCTyWyszT7QLuNbDsIX7wvV7B9QGzf
jfAADI4z0nxzPL7inKecd6oXoqVVTqb6uyF6ExyvnEtZkWToymfkUPFeaoRnTAsE
jx3GqdgWO10P3VIzvZJ2xMHRF6m5VA+hgJAPmiPELvO+JsZlejnZSCs0imIo46EZ
aP2Nk1YgRhFEETIDor9Tg9eRURsbPVtfHxUCbbqKIuG02WCUzAe0bRXJ67af1IT5
nAzNNjzxj4nXCN3f5yjoG9DpSSaWQuHuPI/4kL7zj/sGqWXMarRmnKXeJUcf2Dn2
wy1qeot00Fj+E3NFy9+viXzOUROau5WOsgmtnwmgdYnZHo8X6MGGDG+L+C4GgStR
QUujzITQxruyAW/LKRb5iCYHh+G2fOlKdyY7JYg4U2IiCqi4yLeiGaotaGJuf1To
jMBm1PJutWnhNYwO+XbpXKl/r/cFCTB2r+Cf1ebl/ijzjdWkRs6zTVoLeaXzUfJC
31L/NOKxSOgZ9wuGmpnfdX1gru3k+DRdqwuppkopP3Qby7rImq+RMvFpUHqQ+v8h
LKnBz7TYgpipjTKPewQp9WXIhQBSkftYYtCP4+btehUR3Y2yu716Utwnc2sgfZXA
AOfIDH2JpJu0u+kI7mdh87NpHIZMvug42taES87lT6BLPFjg7/oB9zFBnuAKvXcM
Ph1ADNHNhugpCDIWZM3JnOzjnTvb+u1/Fru8INhlVsXCvf3mKxh1JRCbPUoblsfS
thkp7aIjew3JTNm2aPeN6gk3piAsqB3G6KuM0FvM8LiwVYyswZwiKdavXtgayKRk
au5VcYPH1BZyXL9zMp3hKZZffgyKci0myjF+Qnc5V1cxWCnQ7Lz6awBvQAFcaXZd
KBCSMrrz9YM1MwY01AJZ3YTNi6uLuMFRbPfX1BoM9IubYewm6f8887uyd6Ei0ljD
L8fC4bhwdTdZ/+2LJ6S4TBf6Rg6KBzJsNqxCi/Lnp4Q4ho0cyWLQQuL05mj0GESt
PTA5KaOaQ+Ny668hDLnvqeK04UAI2LZkhG1YL4DrFwonPylWPyZcak4Cr6MTPkUq
S+QX1zgHZyjcwatumGkndGql5AcCsbJsZxk4zTIhZMjcbQC1yfjT37qK1F4tgxGH
aZHXstLnt0W0m7DI0zqDuRjHIlP8JsNHHX4R1DaQucRPPjtsZvlCul6x4nJxqVt+
uudUoL7RKpWA4ePvL4y/LrJs362jg9Ntsirx23+gv7f8SZotjGUpAYKl+1CqIu7e
qfB/603Zg5vELqS51kuXqX1X+X8FaX0N2Mc60Rbom3vohb6LK28/WZ+jbmcL6eZz
lmtJx8tKDkPR8A2sktXFF0XTXXwqJ3s+3XJ5mS8ZhMO0/9PYittkKUCPxRjGFI9Z
IO4WLlejp+p9xG9sBoZjkSEFp02BNr5SYlwuZI6VyG39IHgGv5gRnpf5ydwukvAT
yxyYq+rSql8nYvSFJNUKGWpA2VfWJUeg5wJl9XF1ZqQOx4WaeLFsdD8bcU2aj47/
QijoLJWrNg2AererGqG2UNYUgbAAsd32qeZKLjhAb96HRSOxaM+C0zUKbPAcn29j
Izi2gLV4vQ4Q7frkobp13lAM52mIpTKLeiRO8k5oGjftVvcdit9wzOy9GdW5ADc+
kiPSpR9k2mfNHfMjyd7wvWSb45qfywFjtvKaE4yWyMtp3zwZs9hl3168iVxY+ygD
KWIHewBL/t1/iijgSxLXmMU2Rl2QKh9aiA5XLsleoG2VYWYPIlKiSDs3r3+nBgLB
M1eUo+PLDPg19wHySmnxENbRLm5fq4dCK8ECg9XZaFO0HWP1LfqCzS/PQ2hhUB3d
Bh6QoSEM58i2B4kzOMiyht5elZsrbkCqndytojqkKq2TOuZkcdTk2uNphjPfXiE6
0yioEebAJInH9DhfJU+NiM76FsH5yevx7lbYyEfbxw2e9bd+x2Wk+EARzsfGRknb
jJOxJydDsEKFvgO6t49vgavb4N9osD71rObD4O9tu9CRTywv0G9x7ESP02rMWvSc
ZsAHAsJIyF6RRBbPwRXg1t++ikLZJWS/LuNEZF1uOTgwBK0mbqYaBn2kVhAz1efh
vT8/l06zA1fO5Y09AVzlz8flSvWRWD0/EoQxzJbo+hZxs+fxXCeweGFu2TfIb/Mh
3LcV6Fa/Z7r57xb52uWFgcRjDrdwneGbHAbN8hpnAO4TjkX7QrbrhVhgNggWcTGc
wMRSg56yis7Ek+5roEhWwvYdyZvE7dnHwbqAijicIwNQk54wCrju0WWc5Cae//ps
0VWHuTMfOcvpcnyyYKvbXpus2McJ53iicoHPWcqmupWnyX/bmB2E2quFqYZcj6xO
5UVGzmT190Lf4bYaCGMVjCJhc4f/TZ/QBTn82L1zAR7xMZtrvPNOxSX1fNa9NAeQ
09Pmn6HjoGo634DnqWnJkrax1fBESIaYxEbetJBtXUoPp28VtZVNHHXLBKxo7rFX
0+I0YpoR8a0RmRQcprs8jMyTmy2jUt+bdjwwUV5PHtahTSZT08jT7Gb69VwxjMAs
zBaT3Nvq/Ebizj0Kl6yqMof76aLfBXztRgaDIE7XuYZPGwdBRoNgRFszudlvE3b6
EMO0GTozOxNBqotSh9rQZEPvmQpj2GutTz9zqjrRWwexUzeZ628dfwgQ1fRyK1I7
Cb454H3dwRQbCuazPR1CWPv9/wXfETpFwFKctQ3/j/01pXMLzGWsw7PZAnXHKbyp
e17f2k+84cZ4g+aCRxFEWJCJw8rizxwMfVx9/SHWThl7F23P/im9xL3ODp7SLTGJ
j44v4FN3jayuLZglRdIbxQL78t3YC1h+d9KcFqX73VBQdVqVpEOeR947667jHCjK
gNAQegbMSt8jNRiG2s0BQFx8+fqWeQuF1Z9CWrdnFBf/xVkqJHKsMpYGNVl7ojQ+
8mpTAHXooHf6FP87O1On4oFQMTjLXYhXk9+8aZcho6aZnk+4Sb/HhaDIVuu4FXtu
y8sLbIZpS7z22cBtQapJZzwMKkW5dgvEp1ZNWYGBJw5BDmLykvrZ9jIMrwBtAx8c
naYK55RImg7HUSKtTZ35OdJpI3+2UEHZOkx5Dtj1tBAiOvuX3zCZrp1UErnfNPIo
T5duPSl6scI6Ktf0JfJWsM5sh6GAsBnYyhhxULvF4GzBLevCi4ETXwSo9RwZBI6b
8mX3+bUPBpiZx53A8FVnbwxGz137efQ3KwnEgQuoWQwNQGhXb6T5/9uhD0Vbv1tr
33DXZM+DfmbLVVWUw+kbUUp2Mul2fX9Xs4Z3s8r/tiYBuAcOe2BWcByiZ1j6p5t8
m3eQKFwCIAlRx50n2tD55bngQmUrekiRGPLRWxTjXhcl4PKX3QMnITw3faJR45gg
HpKrB9Zm16Rpi57xBuajYF6uJrRQVtR2HkNXmtqYYgrGC5zf/yNaiwYLoEPaXFGu
qVyHVg1HljDyrM2MXZaodiEvl9xJ1xcyOIZ7S9CpKFSlBuZrj5htBgKP0Dym43G1
ttdKIwb2lto632jFg3mXobSj7DEH63siVNEqmSCbBTwV6RC5PYjFdB1P7wAgS6Iy
ViR2NvIAyOp41ReEf+1x6AFuOCQXqn6qnmCuJjQun47eYxT/MckxTPUjlfVBd3l6
t2zvOFFiF2oPA32/i4BDR7sVc8Iz82/7BjWt5hJRDTdYcxCvYyYNgYu9i7bQ7TMZ
l33hm5scrsbvtqMlgkr/kJ7dLZ/0YCEn0lTVEbr63DpXW0o3AhrqfmCW6hdnBtIZ
Ss5twufkNq1aBJSmDTOf7FXujfEw9fbt96V4j6gVquqgVuqhzoAykJia0CiRpsjm
SZtXPWwrBLnzVMhS379w/mlUEDcvWJMXIg1koOm2/ZCtnexn9iQeDtbKogUOPB4q
cZ8t2x/Y1CwDk2HvSE1vF7pmuFh1tSc3E8nJOeVANUufUcSDhrQJsHNRpn8vEY4T
8iUKuo3SAXFuqCJDUUlCyh1lGDCfsg/ZfMkXNJAiY2+f6Kcz8B09hAgEf1K+9X3E
IuCupXaIgh0jYzbHWihd0cIMZCasaRVWs8wEJaTjQED0BAIUjPngYqov3e2DVwRT
G2bk55bIC+bkVeslWCplwXNJP//qVqTATV8OAGCydJ6V9k66cnwbOlvj2QBAeeZy
C5SX+9B+rTfLGumY5q536qZQS2xo8UT8vn8SYaj733urHlQOfaxYUKqP52GJPF3l
IH3GgbtP2/Dpk0RXH7nFjyZQcee3cOx/G+TkPtalK4AkDdxoRoLUTKZY8vumgDny
LpieSEAUZPYL9QoJh4bEAi67X0gjsTk0w96YIGx/Ztk3b9NWMDgjy2jY43hLt33i
wkbkhoOUTtn6F64iXs5NDpQ3WQAx2Uswku4lJlswQt1Td0v6Sait7EHFFACoVvyw
8A0UjB6IdQ1kCYfODhXaa9xMet6/yKkqlqtE3CzKm7QigFctt0fDkFmIG53+bMgs
PpEvG8xLACMdeTa9UAQTzz0CliMJrVMg0VkFeGOAwgRTy9GZq4j7d7+r9n5Qbvmx
DoY7Kg1H5ly+BFWLMiAinVdNsedSoNeeJXycJ3SFUZKxXs8Y13NpJFcrVvGsjtaT
VcmM4AfOZDhX4hdmZlhycBoqnLW4oKUPFxyuikXrmwIMuipuJs7AUJVPHBxp3Vf1
p3VoyBZLKneJQtTvcU8gD28/psYz6AshUx5Fy5ug/JNA+WEAeY1ABMfbK3P2BTI+
lbuRWkfQNzYEyO4WfuTyVcbBQ9Ymnwo4eJKAMYIgsaWrOiLs3nLXwcgT6K9oab9Y
Hi3vEUQRInZEZFBsLRyHG5Is1LFai/fTGjx3TRVhjmLl6qJpIDR3iiuxYQHex8ke
O1e/l8tXUUbDzMGSnoXrNl9KZF4ql2TVMibEiHLxxjVtMLfIWol+HSLO0LL6wgys
KhImyepVBQvKXrtx6s8nChTSXQrSsGwPMrozjvyMbpsDDh+L6MeiyUm67iOE1CaP
x1/sOwQlOTSzgeO3XlghQrbT39e00ZGF/wH93swhbRsZMU1fAo2uxNVLsATwkQ/i
deq9ZIsZdKsGOcsAJpzmPDuSLZ3kJd0Pdxpt3dIvlWvfEaDSRP1ThXZCWtRt003b
qb+D3ibaN3bMUhwS+vr6IjY9mS9Q73Ny1x28kPTeDi1KT9K1U/y34tbpQg5c5ypT
qaqubh9OibihF30KNIE82yg+th7lnYy3nUhmstEUymONXvgwsqV68X4e0MfmKmpT
UI5vXIeWLQOSMBep2KYA4ZGUGbe8PH+m0ko5NgWf505glI/AhtbH31mIvwnAgdIM
DWhV0VYaugGzCPFZaYDHsg7iDYvnELVDW7VPI3+pOmi4kW7bcTgQ7F4wigitPPN3
8oiEnz+3FMc/zmNUtbIhUNsghgScWntO2WQYAfe2lB++QU7EJ43QQtF1ZJAvu6y3
Y55NwSMDCKCM3pV5l6tRIakeCFWS5WJnPu9uCOoyNRKh5ObVaVIohPXoSTmJOyFS
DBViLRZKSp0FJ+f1+cYpgFBTvHCTcLlYxxVR08WjuRMp2jeSG1eDMCfih7SWj1s+
q/Z8xZG77+057cmjy3JMPtR+CwFT388wLpwWKtAeftkaEkzSne2bvlzFsvgc0fnb
ryp6nRlg6sagKVp5TSVM8BGj4FtOyWUSKv4tpguPTCsiv2WlPOtAnjZQEnk2Aqdd
l+M1xRImJcuoBH/rr6h/kuUlPfzZ8lwVbdO0su1CCSotpRgq+80AZohM6nu1hnNR
8dEf4BwF5Rkt1cagdiTfgINsiWCiwgBkuy/fsL4vSFr34oLgWyuUd8/UBNq/C5J7
RIere66fTqanDu2G83JKTsV8K6rVRoWzsivzjphBxNKT/w14ydzZ8HDGLJ6ehhqv
kxGuj1n0D01PFNSHenACUsQVVMElOpW8dKsScHelcAby5bYHPqw9LZYCRP1P8xxT
fKLFd77uuaYJYUdbb6+az24EsaEg0Kmik6qS/xZVezhViPho4MTbcbwc7Jy/TiYl
+poFF1Oe/O0W06AX4RurCev55hrOR23Uq4cNzBggggY7YM+pu9TppY8Zpyb1MVXI
sIfw33R4QmpP4mhg5icfVj916PnLWf3wi1hwhVFHOC5suGTIdNv9/nbI8+2x3UGY
TcRoOE/+vQ6Tclzq60X9mOZ3QiEGZcqUwMTLOEzF5Bmvwv0ZmE4O4wjHjFiHprb5
oL5GEbbwAPG5pEacth1knC4nb4rbDWXMOQshHsRBj2FK+zUkgUiswxpMXzNUDz8m
Lsk27e7em8p1sd6AN/tIhFmVPQ3tFxTnT5jyciWyEWjZWS5mzLgxFJMA3t+f6iwF
FkyiXp4alnpV8YOpHJfGdCU8YfYI2KDvOcKSJe2JhVFDacAiixIKdYLrMFH2svns
71QJbUF2JuBxeLuYF90UlIW2ZxuPDvMxSEg4hV3bRZcQbLWZidGIjcNFuNOBPQns
8SRfDnBRgDpAkaQQBddftb9qYN7TEgDdNinlfYTTc94x4Pu742moNzT3WhvfVoaz
XKrxVGAwjn3lFt980fKQE9Urvn5aJ+G5Cz7Dnj8pf/Zb+9BwfFy4bfEn9SkLgdyG
BqkUDlEC7dfg13ZTeRLMU1mYZGWKBNwhsYdnkMZK4yAe8C1CFg5OtwnrjVAiqcNk
K7rGa2NGfCaOVu5JIszwkeBdzjYxSY1/tBPFzBxC5bM4ttTbhQBQ9N+FlnkNGgrj
IhFiC0UWYv5ZuLLWU2DxFdpL9hAehh5YsJoiSoITJn7cmAsar5bW7zTktG/toMWh
FPEHCKGYNjF9mX6UUjnyHgAcuXS22OPYFLZJN0sQ2wfWX79e1+E9k8AaA2HNZa0E
tO1Pc2MCxty8Fu4urti8Ucma7RLpY1JgoDJluvAtB14jWcOQ2Id79ETMU28ufumF
DocovTpqXx8BxECaDmwe7lMcK/+p/D6qRKM25rz1NZrdAQ9YqoolTsJ+wvRmM2zt
iIUfPZ/tIBtgmOc1raFp1LKZ0OF+dxydFeXmlZ1DfrCJJmnoAUNAAzOmshkwTfjR
Yn1pN3mCMnXn/jOTRj/Zbt6fuKi60ezL446x+h/I+LtDkaVzujVNRTwckzIQ2dSc
YpGE9+RYUK7ncuTBCZEne5wYACJ14ZaLx8XhmOn3lGZPBFXFZfOVAych7mD/+kGG
407GGhcOQhAbxkG5L6jKDD3VMtmqNx9QOdg0ir0+VM6cXMVDUQxqebKZjAzNrtlK
Jf0K0FnYu1hiPDXxPP/8r99kLbt8VZyhzCaXz/25vQd5KWB7FkN8QPOKBsrypXAy
SJ9tEy2WeGqtcmgHQ9vNBDOHmcY3IZUdR+7G/KJgSt5oboBaUizNQPEveEOKWFe4
Tao4+d2CwELmjPeDLOV0V2lXl0RjCzT7MS9rGKXYDHMQFT684s4V+VW9DbHZHi/+
yiB4kdkojaIt8Y6N+KfOPAqYcocGKmezF/Bxbho07isIKjEVHPgsVXYOFHRLz+6z
zSmAoEWg56Y8J/1/cozPF8IbeuYHfEOMAf02VV3aaPlJm2OuIWId94+mZ0eo5uyW
N1TatCfxSs3nUJdMmTFCx6RUMCR13IUUyEY7yz9lhaJV5MFdE2P0x2RX6gfZUEQS
HUXjDEyGAYdX3EqIKcWznUJI87qdSgPbhXEtfpoi+d0T/qRIh7iaBDpyBm7IQhbJ
FynHdcBVu4IOeyeHQOIc35i+PJZ3dxt5UurE7qSA1MWOLpP1PPORdMvQRko/dSvJ
5hP+4S/GHQvmW4NJzRePmof9n6DpKa9HvfYUXZeDn8w9EFjiLQtU7u5VMbyZCwmV
7KI0kd2KauhKqCxlgt1fOeeknj9skcAGkiQcC5eg2xhR/tiC0PCeMTahrgayjlti
i1rbLrdDPzrhratde2T5l/eJbkNC2Xr5mbsGbyyjYkZfmwbyDVpXAdadcAGVXMPT
X+sYhjoLAjFPc1DZaTs5eGWDggg12ehrhBK85l5wcm6qml/20aLX9VF8UQWEsnNd
YdxVzMcKx+gd00NDKoAzaH/+c5zSV2iRqwJQoaCCohYt4x1SY1MpC93xpZ/BA5dF
qyVo2jHqxMzSns54fdL+5d2BLfJKFxcjP7meOwryC4Z2VpbFNI8C7DSgdJ1dDLNe
1Lulp05D8piG8jeDPOtDD3UQwsYU41REZoK6E0LolaN33Jm0S9WbPLUHZjIcrQUz
8W8K/D0g6eqhSkFh9msy2bMkn5pYqT0M4+JIPEVq9T8vmUtoX8XsCJW9+07PTmSY
RBjpciv+9n6I0nXiJ1wcNRzK0lVhHrdSc5ldKV+7DnQAQ6QH9cK1SYgpne690oLY
AnGY0R/V0/k+OlGQEgN/E1W6I+nh8ccC64yI6tCC961d6slCYcIuM5JC/VxENGqW
S69M60rdDMWWiihTflTRrztbR5MKPV2RYb7ZNWDyjyRO9G+RoqTBPsqiiPe9bUmW
GgWLobcr0RGS9rAGzdarbR3DJB6YKSjzudT+7ENbMA+wsas3WVwJcSEy4R6KYf2I
nfbDPhg/qtymdJY/IIh2dyGiYfYZdVgWXEcHgeBtTOS/5v9ajN5ut8jLntFOd60j
HNu5aWkVZsj7/KCLxwHv7SrEDuDJUAoscI2mxz8i6j4vHxh0Jn2WBM9fF3CzNx17
aQApOid4PjbaMQ2uS7xsNn4G8NLx0j17BqHo0J9ny2zxxYVcIrG1ZNMja8P+WrXr
PKBtLMiacIG4O3ZDUNXiRx0MlRUCD0WjIMjhkO5xyV6NwFm7rUaVEkwGhCFOK8V8
aejZUsa8pT59TLFcHyhtGJLt4WXm0Ms0kNFHGuN7vnWSa83z904rjwFG5Euw17YZ
rNZ5YtuipkBeDYWRLfRbuYFIK/k5dJ1tChKS9iE9Op6vv3emH7Yu+qDiSqnSFLTA
UFl1UmW1ouxFquAh8Wwwni9wmZuwoPr64sje7kWY8aQ=
`protect END_PROTECTED
