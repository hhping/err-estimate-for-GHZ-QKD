`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z4VGbWm/zBrcfyQct+9pIrtWYfXibKMFzJ7djZVSY775IeNgkuukGma5PjZxaMFE
7hvT+eMgtK/OGQyC1wsi8LH58FkPtP2NivzHZbEb4I+8e7O0wJZflAhdOqCITrz/
ZjcxQ4pCEXd3UPxNpf7as196Nc3bgXzRiYhAEnm1J1+V6Arf2CuFGDbYfCDNEhxL
9I7aVCmqAgT4ebkOCl5yC0A6k+p2hDJL0TKCwbFn+cmZxVGTf4iASqwNTpFk2nmy
5gSzGV9V5afbXgA/6JDLhOfZb3tmeQyPaFAF6uf4QjNnw96/4mJC9+ofLAz6kukN
67//2CCCzMz8XwyBO35DSN/ywktDA3qFOBZ6lHEUL+viVgUet1hNzV2ro8mCiXrF
87T2UNpSE6JjrHhcD8U4ZZxqRMLJGDy8Z44d+QSJz8Yg51XvI6YKu1exryRoDNWl
XYJnXvdLnfecoofo1ec8BNriT+duVRkYRHHtcL270cVninaonSn0naEfPZkSapPN
uojpnTvjLDiiSJitHAiNXRF9WuQvSUxulLZiMNd6qR+LqhWMoxtDUq9TR1ymwSXY
FX/7bt4OlWA+jBpJMcUvVHw78lM/5dwfsNNWwwsmGqyLKo7NhkysegRiSyUUzoZG
/tcxtzu6Mo9yBNzSKLhLXVHxnINYpgkMOdphpIqE6/SpoqdriFEBYTPYXjZiQkfr
e4NBpgth3nWhzVms45uadNJ83rXt//aFy6EnrZPmd3CZN6ujCk2g38s82l6Ix8hJ
ij2jRIEjtmrPn5bMdzjmSOoP7cedU89OjCXWqg6Qo+Yf+Nz91dXNfl+EsLek0s3p
imlHevjJyG5gwjMLkOqM7oXqLEw/XAFerD3j4skIQngrRpvonagXFmaZi/4oL5Iu
X4zeb5iMB3TUwvxiWkDs4qJ4BrLEpr8Rgz3bWfbYqtbUAGWMYaFk01HkW8JRcafq
GLgeqMvy88YoP639vBgumNy+Chcaq3GkSZf3r4fsJwfK1xyi1UCs7nUN/AozNd2C
DuiE6fNg3O9V3ZIXdhqO5KBGkP4JnM7wGh1w/w+9ZTnsc3ughPIypSMyqs7J5emB
S3aY/u+oLabEu1yAYXVNuO2JRDWhmfT6wO9fmia9Tlzw0Wcj/hroCI/78DRGtdKC
wG4ItJ6faHILNab+BccoqlBILs/th/mB6X00cBv3+qiHlwiV3bPHQbkElUWM6ovr
OqHw6cK3/xvLqOXnJToA8oKT6rtji9cJFIYJ/m2EjcGxT6JOk3wuB+Rippk8XARh
`protect END_PROTECTED
