`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zQtwb8VOfFqxKcVWXmrA6yZ7SUFDEgW9f5+Zki/nP7gZCQhgOaIxbzScAVCwTaL3
GY68Hgm2UqD6hqnktr4SCINzKc5jJtxrbXDDk6FNVphgWN+MWbGTVGl8OhUazMyZ
iIOFqF4PFaMDjXkLnQfgMzjOor9tTfWu+nNmkzz/lPncEUXjh1nAbKUNPlz7dQNm
1vlPySdiDURTGTAPrCGY9qLJdmt0r448+jYzj+TwcjvFDEVXT/8Y3obdhTiHpGse
N/30RmhPZlX66Oyb/Z86gVxSTY7st4icnizc6kP5XrEOFJGHrKhnI8MVbXVHNUvi
NEzVWY/JcK6bNFhfZk9pBh33pNVawrOIcUR1a2Q80bhOzzEuUYenvZdpIb7DfMz3
iF8StBwoaK4z5PUUxC2ZYLHy0mCquB/suk5bLHllvSM23so5dvYY7MlE09+opRIS
01+U8GZOquAvGIEvJ1xapQ+wOYQDwQfNKcsP1y26mdvhYrM31FZvpbq4/h12fcWb
FmMb6eQ2fDDDP4RKMQ3RaVH/d3InnGqb9wK4vZCSaSDecAQ1mrQw+WOePkVNg/Pz
pTlsZ3Cwug45hXXGs1H+75oZYsnkA7yGyNhpRiW0nC8Wh2vPfFHM3QesOfhOIP58
muEvl9xFo0dEMCSwwtmCds6zhRL+bgsCK7jSC2UbU0DR60jZHYf2ziEyl9QD3QUx
Hf5Csv1Bcd0tQlaOzDNK3B1ISwMRvreJATEVoNEALkCKnu4CZPZWd7EvKtI1OOH6
+OIHbRH/f/vTwGXJRg5j19Ee4w091yiSZmeXOCfhrBi8JyzggUonuGorE+9tEipl
Ml48BHQ5rfnVb5WBCUg55baadhkZkwlJDe76LU9kB93ql01d2pdi+1kz1Ic2ROvY
BZUbOBBdsfvkhqpGxnB6oY26LFwA0yAtDBWli3BlGp0=
`protect END_PROTECTED
