`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wGaq78oTJXlTIaz/PBulPLt2OLiRflt0HCOyRyZFi1QfJu/oy3hQRiv7+U1z2J95
oJi55B2c1pYsmIvlw18CEITQI29frv4TLBHJpMKKHzAGAgD772k+7lxU16MZ183U
p+io3IIBhkIrQVemo/NE8MLQwsLxN6csSizShVUTS/K0TDS8Cuajfsp8qemrXdl/
Kq9zMYiNtnd0YzYDPi6xxSYg2iWnHgQEnGTmtEbkFEuI5slmBu+7Gl6EPBkgVZWL
WtrOIn5y0wfH1aYmAqZ6+QEYF0aU37bRIpYKvUJSXnklNvrFarFTENtYQGSEpIXM
IQEGyFpiRTGEajFvJfDl8s7DkcpzbN8y8gbFdn+uPBT6Wf+wLZBzu5/GYFdRro3N
hWJUMiUx3NcfS0jaijuJvgg/d2xgA1iQSHT0fGue9c0NBq+sXNkt5awAd+WTpyd5
M0PEr6D1lnlrQGIBj+Quk6WZKk0tCfEdqDx5iVRmHnONXQ4XPvI2kbGqv4hgP/Gx
1NiNK88GvVUHzXx692oy8FWxIkOu16G33G1Ej0N7zpI901XeCg68iXgnPdc7Coi6
h/8+NKdAZdvPGq9XkJ9dKMxoIfQIQw57SChmXomRbZ3oRD0JCtOnmAsdOdqhNpwu
Q0z4tCpGbTFfg0aK2bKPsKP8UvW+Q15qCSsZhkYcpFb/3q2mKGSw7vOEr/RVrmy/
SYjussyKTBBjEFSp/kESMeFZWKM7FhhVydmR9NpdtLxywzB9scB+E2igPD5HOz2f
Dg8AzLs0IUEBAaZJK2C0tA/3m1tfGxPG5IkggmyyI3y3ew/bEVaIx4aW8Bt+Hhqt
ynuRY08PjFFgkxHOMQKtbzm++5uXG6w27ZjXXp5+gSj4IAtE+RlPms73BBW2xAQY
uezik0C/x9y4M8FuVgLvFWQ9KxxTsqHHCpEj1ZpzdiuNtiys2kzHLuLWezkI8HkP
6Kk5dj6X6u4M4BGQoJNPH6bv98MalgWwwMTg6Wzy89Po5Wl3O+ga8SFn40dmKhtE
mtdtgeV7AX7bh+Yg81HgMGM8il+NzZaEGH2PyPNMhf5q9B92GNySB4qAQFlkyIeT
K3HMQ32K5234k9syCBdw/L5Wk5pfEC9B4r/ijXurWZKinZGRvdY4v8NYz8V5Lc8s
dmmiwd66C91LicqNuFKiPsAp+ommj4PrSuLZXEfrk24a5O2T02Xt0SAp9vd+/Fs1
ZxuWYnuC8lRm9tmdXwM/t7UrsqhPmaq+XuzMeueDtn7xS1dik9C0mv4/vkM7C9d5
5m8n8BslnMSR/BkeoFPSVjA6BmtREq1HC22361Q1U9D+dW7XlcCYTo7/vogO4Lmu
rDUBQ9+ErcqcamP9x5rj+ZA4uUq5cWu8ugqGqHg3YVjL+CBPYIne0FWDoEclJmjQ
vhtXrMeTIKTvogudt4WkKrvM9sdBDd515zcHHlAs1BA+52Nbt3CH7i8JHb4MXOoX
gnVwmtjsJmCUXpzVPU3vL6phb6wiBOg0aDeGwhC5InT4cHGJPGzKE9duz+Eu6gEs
na0voeEdYkQhtyd2g5gqtD2wkFPwWG6Il2vNUwdJrRiiwceSkdIC0JOSoO0fjydA
w8Z4dpRHUBiQRWtSjh4Q3aVP0pK6EGcP3BSzOSbRRmiIABYFx/5WFmPmdOZ9Bynh
gSErsqfnbEbABo7HOimR57CvObRzlLJ1N1GpukZIV9eJu9qOIxJyN1qzCacFIGHC
38DGvaqmsmst89vYgNKlQfDzW3L2yeghPHgxYDKolw5Ons9HjGwqZMu41hfSYs3u
TVY+TnDDheV51YtnqKqx7rfdS0otTbUG/d6Jx+2v65cFpzmkQgrzTSKi3oJwPbdU
GIUB1vCto53m8PDU+h6jk0cgShxqDfRDh3WLrIDSzj1yIHWAi6NWksGa/i6LAUpm
p81jIQ4J8O4pxB00FV1sVFxkDh7S2n5X/9YHrtWDtCdndmOO9FjblufFSQO+rAMn
QEINOmsucjHuEjbDu5qvHIrozH1AciaE4TJx7puT2aThDvA0yooem3pSrTZUYwCK
jYMUOnUfkhz12ULDY6IFClGLRM181eRIlCtmba/CXnY=
`protect END_PROTECTED
