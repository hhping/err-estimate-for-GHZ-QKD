`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nhMpNM4UqoRPxADgPOFtaK+V6rt8x5YdMbIZ88jBXkO+oeqo/s7YxVvQrNpaThPQ
bzoLOtXQLZuhUqHLeS3asCvf2GVttb6DQpkL2b8iC5hAaxfEvtW+h8m3DRAXK5B6
qjk30psGWCZ7w63DGqeZIoj3YvRX4S4yuYtGrXHf9LOIDZDREmKogClvWjs5W1HR
9Qb4ltBrPPEfzswiFbw+fwCjE4pX28nTwCuYAPNzuup3FHA3LVQGsxnhpd/KXuai
vMa97nCLdD846Ue12VniaRlEaOrKQplXvAHeOUTLUsMWZFBrmQc9dk0g0PqcCUZI
dHshxd/Tr2i0b76SmntPz2hOals1x6WXLDdJELjbR+7XmqEEIx0F1ovHUAW8DDlo
ORlHekzqSH5Ge7Bg9r9e4936TX/1io0mbUdYZBHEW32imUUlI71ceQszagt1bjDP
jnSclp1f3Lj/CcneeZehQkSInmBGq226hKAjTyUKi79QdpYxThIchNfL7OPp1Jbv
cFaNZP3CmLn/Q2sSgV9cKdOBMhm4kEAIwBBi5Q5E+IfoPkGg5ZuTSEIh6lKSLbY4
QgI/LApgMIOluQMxkb8S71T0PLKKibP1BaDA7OR2f/Zuf+Yq/2C47KR2p/wMiPh7
q/84On9RlE8tfwfzGJBVlstnZ+W1oCuSvQOKTbM4KSE=
`protect END_PROTECTED
