`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yuXc8+uqZ0pjotIXfhdt5Pd4YbNDCupCN8Kx/v8FGxjOBPv7hygNYuJ6PS0mao6N
uuF74PH/CPizQe5TmgY49JnvXl2diAkVi7CS7Ab5IJq7atNTd+yexwjqZPd/9KOG
jSCX5LGPDJu1zamIUKbkhKeyXsXCyuJyy5fz9Mk6Ara6JKlrysARVQfws5fnIXK1
SumRbmkRGPw77LkPX4xtJQpDXLlj2RJJMCdSImpxbvkWeEArVFbHz9vEU1XL+16J
rKHbqEjp49d1jmjcJcHLuU4oz/hTaTbRGL5CbkX9uauCaIytAuRVw22V/7fEVc+L
smeeR6zMNuY2UbxgiNym8R3EQ65mtpSwuzYcbS7m+dgyeTHY6Q+GrbipAbr3u6mm
ioLxdEpkWyP3DWHGP1mxi3sNgW8OgMvGLNtgg+XtNd5xroKxc5vLvR3G2Vrl2WVP
Uu6dOAc9Kowqx5aKbJQkJveCwMkEACzLMFctNKxADtyL9RXJ5Pkf7AqDj3a5CidP
oj0ifhMgwwXMmDEGRsFMo8gtQIEgLpUj8vZRU9v1OzyoIjtp8571P2SC9088+F+l
oAUKJMEQQi+BZsZLsxoc0PXkxAZN3URE4T9U3XTfNrY2Q8aLGfTTu6WBGUosSgm4
Za5xW8LXq9olWjGhscB8v6RRv2EQ4uo5YS+KJZTw73YI0sv6IwamKGaKW5CDG3L6
IIUIz2cZNcCb4TThcsMGjHSKwzv/PW08PGvXHRssrn9utzJiWnn/8uMPEmPsk1m5
557H9mLCh5f12H9CWu+VaKRQfYPxa38lpQsOo3A8T/4P1u73Nr7+q62NySRNf7wg
cmsxzI/TisA0q1liXtNV52of73cR43lpTTVnE/eHQWVu7djbfvfeHoa9Ncjzlr7n
nX0YpOxpT7cOWFKU6XhQP/FgMTOFw0Ax95a6gnLI1DvPX0zUnSdGIA4redpolc5O
UyneuOBbrd1Kz55lQkLgSSbreengENotWPOEHJ5+bIp8txuCtJUGCHanpcvteJ1i
O9UVVlXYSEJMQ/ZwYTr/sMLkLrLnk8PbsORSiwXAWpnzlZ8BGr3UC5+84JR45ZFv
A2lVxwXZYF4I/gga8ar2ne+ElIES5T8ALZALvKRiaUZkHP3DvrFdE6B8bNijt418
4+xzvS0z++6e63/x4SC3AWgmfRjLXoNCchU7Rey86Zz7xuBWzBAqpwlcJNaDPou7
XtEencUqhS9QEUXxwxtGu6LoUrw3AglwQZ3/qiLYQWDNqY20g31f4MBRiAqMZZP2
cYN8ZHmBjHfHbMg7lDUgfyyEDwDIxEEHLSgeKgdQXlLDbuH0OPefcQDqJR/c980D
gOpPeANAJC+HMiuPpgETj1oCT8YZ0kH6Qc+nZkFINpJrG9jE/l4DNV0incCoz3Wl
MJJln9uPY3D2D2prfoMw8R/XTKYlkgtDUdPEmwgnVtJ5M+wcXhKCDLZSagBPxyXe
7X1HR4lyhkWBbVdiEVIsEiWd07Kl0exsLvimtvpScbUmTL/FrRa8YdifmxVk9I7u
O1VLdssoVRm+CjCMm/zZlPipYTNp+U/91NVjWcFTGes=
`protect END_PROTECTED
