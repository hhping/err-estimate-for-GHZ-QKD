`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o6rlvAEvB/YRSLv8u5PWVmiPeVGDfjVQAFd2FA2FlXnZRKHWSlHBnf2UdoGaV2NV
716byO9BtyEx7ArWOW41j1eA/F7tbe1LZ4ar6V43d/6EiqJrg5Xnq7mQ32i4mTy/
ZkvfYAUfB3v0FrXO8Gs5Gf1z3zRbmHL4NGWfmoBP0N+7VFsLw85VoD56lghD38Ij
xbQklZpvMCXI2wzZNtPWgHiiZHPp4W1jjT08pCIkgcQmfQFsv3ssNgpJoVhjSPRs
rOJuvseBVTIgUBIeB2hov2WIGdsn96PhN2ijgss9cVDE+abokcmPUX+w3dG+bu1l
4GiOZp1+pIW51QqLgIxtEKy+N8ThlgbwrEVPemmy8V3M05rnWp2ZRMMl9ayLljFD
N3Qi1e/AxWAgAwV5xHpxNLLPnJdPZGATAOLlkoTp0vQ2CavKgwvT6KRIyOAkGnKO
RJF7w74nK3Y72C3d4PH12L9t5emhvOS05cGiAIm8LGjMVXgS4Yh/YeyDyEr7of/T
2FNXzLvtneZ8CvG/t8ZJhorSMHYa+ZUSdNLQOgZ8fFW4ATWFe9oLxmHnFd/Dehwa
+uslnx0SLRBRluFxkHdovvSZdV0G+hZDSWg0MoZRpiRSqm15Y4e22CDkZJnTmFJo
G3pf9BmEVxJXp3BgNKmC0hZ+5VefIgG4d0wZZkcggO7OrfTyN4w13RLSHYXaBCNa
PfP9NllY02rgcFlZ26Hwk9usoAah7BdN2sWvKIKfEp0RF2DwmmiZ7XnGu03FLH5p
QsTpYVM9kwe0i7rDFHVJLe+Ixxedi5kbsL2WEPxp4wOtLvGxVC0eewpoAyMRV11I
9RikOQxQUSdAQcG6ssoVyIitJMALMXthYKnyz+YvwsGKPblhC/CVJQfeKZwqdQma
i+d82w6pSDauE8qmYNgWbL8Rl+jofSBy8h9i2FGAv3/ogLDk4KAYHfYSI52HhOjy
nIul9hhb+w9EiXv2cZccCTHiF5/mAalbJAVK6BFYbuopAO6D5dd6Zsz+AF6QjSRz
sgyvcARCUiaLafQRGbEMzl1RbvSKxORTr8W5Oe/YGgte/RHgyNr+esDXbxEQ2eRC
ovdv4iFSJxgcxbTYIRVGuU/kKYo+fY/xrkDc2BUKwhrCfGr9lc0spkonKBq4PaBL
`protect END_PROTECTED
