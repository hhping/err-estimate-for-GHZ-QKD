`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0hPEQNjE+z2PvjN31hex4PGt8eDhxAV6t+nRkUXnLgP4sBHWkWb6n1NrpKVatliA
14Sx5fb11AAVFss/5wicFE/EMbxeZAvr0bKiOUjeoroaxHuc9E0kFG7HmMo4bKp8
HXGOo3zKENwLKT5qIUw5MeDrs9ONU90pqtp6HrHWUQNOJjhOO803lLhBM936Cerl
qp5Naeg46O8cfbycYRWlYdIPs71EExGiQR8BNqhnYAQAm8EbAg2FLl/8T/OEYb12
ZMG4mZT9U4be6IIgR11mCb2REnWTvXf8I0qqdReNZOKtFZXQYRZB4Hz2xM2n+Yq2
5I5gPjQeQ0291g/dzuXMQt9a/8DonoblWmEm43I3kwQ459joI5cPPohGOHmN+h1q
uxLkQ7rzp9RzaaNWyRkYCZ3ojrrQJ0qEmWepkTcIRrProj5phyaADE7FUBbhou1V
g0e6OxeRT8tv7pm5H1h2OpeTkqjpii2VE9Yy3pqS5fCePR0o8BnxK6HhWAa3h/IS
F+eUgK8ebhMO1wXp4FD9j9sgDFcocDN+C2de4XKaZb7pbfHNDh7UIDf67y7fr5vi
vvLdt6GOjlxhoZmgBsZ9iA==
`protect END_PROTECTED
