`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MuzZ+hBgIIzJCehjVypLScdrLzTHSzn07uA5HU9I24NpKk38B2deFCPYgPpi5fsO
XDVSrAHgnuVeQOiTHGZnA50F9+GLSwjj14Nl41S5qqHZClYyipk9HUe3p6xAEFwT
RC5aH0XjSfnZFHiJCjQLZrkwpqC7lauMwUQ9zfmeQgJPtbn8OpBIAg1yCwHJ9u2o
j89LGknZZWiCH8eIj8XanpsTZZadg320I5nj4oqMRWehiMFic53CUIL0DZ8Emf7Z
bTcnYUF34vncLlGjRQoB18odkN4lIT+bVA2mV9myCBruJGq+9xFFbZO967AYU1EH
XOGXdDCA97ui4ym0M5PCwe/Ign2puzJC5h+Kow+E3UXQG+wALEJWzzxsYykZOC5m
wStmTrNQHpxb092IEH90ZJ6WY+qfc3E6FrRNuqg8OhHPBPXO1TyY3VYQCROPuIeB
utFviUs3cI9uC7I/AYEK+EVOGNsdx2QO0qayMXMQI+dOu7mY/lCUbj4TnYVyMzBs
fVmo1q7m0Ol/sLq5VJF//JSSgjL1lSV75v2qhA8KbSJwG/QOXcw7CD+vGsdSuwY7
04HRhQu7xoI/XgWe7MCVmx4d1B6f76UGRk2ckgHBZ8IWXnVCRWxYgVc0vCQVnQEz
BWuXjsMq6Hrn0GU1IuFBAB82rW6bMK6op6c/A74V4tHlVN+XsLQnm3HEuyrKomYa
wfSwHXGxsZwsPFUwNIpHhBq59uT40ecgwFVpz/Uqyo/s6iRkf74EiaXug9xM/xD/
uU4LUtwmt60nEtGtC/JmAY16VZtCIe16RlMZsWeuccmVRYRi9Yhl6anAzox3xubv
Zb3BFCEJyYn6k9sWp+X6r6I+jvyAYedbMExYQxyrbmzGxdcI7AV/NjIReSuTxpkR
daNVdlGfzRy8jN3FSFvUogsPGvKM9iEdQ8K0dNG3p9sYgsvSRJvMUos921yO5WXB
yYatc3fNUm960YnMYLtjgLp5WZjpXNR/dD6VeW7TRcgnEetQ1lOxfr8vVNSMbl+m
QrjPNz41ivN4bBXtD4bZneJtv/JjwBdT+u4th1KttyxJd9wXsb8IBR6o6p7V4aZn
sZ7s7FBeyEFZfbRZZ2GyyA==
`protect END_PROTECTED
