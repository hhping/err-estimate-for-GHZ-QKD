`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qamhDHyXROcm9IXq+Sgc4RG5k6mskmLM/cCWa1Oehgv9KsZCKGHwoELEPHw4qQj0
b3ykjv7fbPkDO6d8EadPeU+cf5/icvm7DrwjpYBTmiX5/Dcqy4Nv204GkPpI8x7r
gBXtD0g4LGREfyyYH6dvFDHyJM49/bzwEPiOpLSqckd4es8cV3l5CkLnSlVvWH59
r9+jeSQHWhTdaOw5LW4WnELMILfsjQyxZdnZUv1XkAcxtsErTOL9snylQbWAj8oH
JQ0fJUrQgsUH2SOnDWrjJYGj2Jz3r+U3GJonO9yEMoIjD9Ql4tDZZo72w6UrZUxn
RYn9hin6j4ia5U0ePnHz3HFiNewjGqiJdyMJCa+N7gMActzCr4w0JWRc5AmCBaMd
ERFSI24AP2b6mtTRFU4sgupuOb83+tATTrY/UWeGdzei2lAhchVBM1mZLk4nK38X
Ti8cb4rpvPEEswF1Tth7OuIrjwBddKzzcFlxR966vGI=
`protect END_PROTECTED
