`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fBpK6qZ/YTQOlvHxus4w58lheDkeTCFTQYPUij6LwpK0xROWho6otwvhBbS6Fchs
OYtMf3v7LIqMW+CUxnJB1g88dYkWtA300SB4/RIleAWK/cxjMjim1eZecSQf5/wb
VkNqscVMEDebARZ5895R0i7UeoK1GA54rE9Pk+zEhX84kk0f6fxGPY5cU7W1n9j3
SkAGdUkCWiP/GUxDr3zMI6Cpv6K4mNNuoOYU1Lln9DNLkJ78H9UekKK/+c/DU/Qw
awNKecI2MYDClMFQ37hfeIx1Ljy6661ru8KM5E9xZ093FoLpH68QZjtZuzMEsd/l
APYfO1SgAwEd4L0OxwqLDOy+bWvnZptnPSAPEUWHFrV3Ez4zNt114jjdkL+2/XV8
Io/YZuBs4x3gK8wyGzLwEUMQNBC+qe88MoO7Ium48HPPOxfyvlJz2bULxk3VLD3q
+uiKAoYf9gBP2ZGHyLCruRCH3hxstEBPdvrRmCw7RrWP69ICwblKb5sR1yzeo/FF
AQJZr8Se7yUZhxB5HlHhxxf9RMct0iBTZzkhUJcqAGgeX+hPWuqIDboBi3X+CUNE
FTxIG79qJRR97XjTlcX28ugJu28aOW/fBM8FXO2cnzSwhnPmphTfU/PHMHfq7L0e
qqrjBxjdfDZxA7RFdSs+0w==
`protect END_PROTECTED
