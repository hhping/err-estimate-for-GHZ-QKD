`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OQitzPfOl+CoeWE0VOl3mCoe5xomiADAP0wmzCrbo7kLHPOGMtonROna2hamdLYa
m9hl0+GgMZur79FLNVa3ndAq5RnosDkAVykUn36Nhs5gdm3LH6EA5KXYbi8p0D3p
rjLTHwM+EQX7aujo7IJCBF5uf+s2pc8oWp9/9C4JUwovlPbL8ZOxnz9G02VFhX5E
lI4cw3ShbI73/o+s0YF6BUdiwuDPsPYY7ILu4X9omSp+yv4DQ3AleS/k8IA48d4V
9EiMYmDDZHPiIe5tghOhRnhpgrALVlhW8RbZHhreKVoLsxo9GwpUKEHrIYVMy2bn
4ddwI636HGtOnwfLtceEjjATSNM6gpq6gxG0l7BIXl2lfoTsl7n13v5bgSp7QhaY
e4e/oCvO06QATF/SeeG40NbVyBVk5Bwh3W0fy/kwBlLODABxvoIdvmQa30AQ3RhH
uCe6bkTOkHIdTfEK4+77fgd5VNRcac8c3QXIkqe/JPpeHxU9sASPe8oh67FhQV8j
As1SPi8N4EElPS57Tzmbgmj7NLf0m4R7kM7lxwcgtItceWPmEN2FI+1U6o/Pu055
DwipGnGk+tX/iGeecJsOAaK7cHDD9SDEq3bl+d2lMpaMLuMyOjVm/nekQNSB7oqm
dSdRMuA9KNw7+qPjOAYunM0V0Gz3G4W1vZXg+aCxINi7BQsV4jZIDSXCos/C4PGp
NDDl6KDPY11WGHJAIL5BY64YiHjrxosRr3HKvhnUoRh19VxN3W2R65qH47XndHpe
0/30LG5Vbks4Na8Nelbs2nS2e4KbXrfEOhRJl66EIm75AgdXZUtGlIqf2Dk63qHy
8oYl1/n1RVxt6Z1eK9nRvLmt2yfTZT6sHMEmFqTozLdqZbRpL2CFj6pt7EfGd1Qh
n9GKisIMzZOU/uJ79n+HWtHALr0a5lBX6fwz7jGDiy+Yy1perp1ZdwMtHOrOWw8k
8KioRRJyWMT+3uEJkUbBFvJT1Z/Ptj4Romu60A2fW4eTkNtJlSMzYsUHDPOUeRCr
`protect END_PROTECTED
