`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SrSgysj2U4qGPV4of/eyD1+TXa95/DL1wD66pOXLFbwIiBINkVaVEu3uTWwUkS3Z
IKAn9/kOBXWTFgwhNrCpERuzoASXIOpxE3AIgPGmD8EWfnbhaFLz27O/nqNtyTR0
py4codp7mmS5VF/WAeBTHALxFwKmOGV1nwbJFYgVyj6X0eNIUgD+kvfJiDE2a1ZB
WySZMayD30xVGlCGUla8DuLm9KxZDCOtg7XvVkKkluOx1iN2EfatK8IIhbuOmrey
gRASdXcbrplFmqVZb2U1V4yb4TaM0/yJjuPUFSoH9hrhs7oMKsQRkE89YGA0Q57M
uLjPHFg4pv+uGVnnJV5E27AEfqZvOviKIkYh2bcmRUIeunchnz75OAhPVrzXiKZP
D7MAPMc/RS0E5IC3Dmjt5TYWIBy2xSAb67fQ2tpipEHrDrR1snTM+vqitgxALRlD
wNRbVOIDbm2kIUiXU3TnJ3Nxn2ZV4S5wIFJjcB7syLx6df5P2WcCJGyiZs0f9sBw
tpMbpl1RC9aPt60Tlhw1AAtWolRLqQr6HqPTOV1CokKarh5+4X8oSOmvZzxbYbb/
cPBo8C2tCy5QqfY6wb1R+RV1uaw+ayScW2EDoEjOsmcoT0/b1btVo1FWfk9i5876
jUxjJSvJIcP5kKQgxFUuRh0L6oPugGrs0AwSuhRgWDQuJHTXQKOieV1CRklUAGNG
yiMOQzxzLtZQQeI7s8VaM7l12o/loocaL4bALaqROtidffTxfNCqRv8f1k/BAYNk
h4RR4fnqrEQ7+PouDlhSxFb5bkPma9fx1KNwaoEf6qml4EWXBa6A4T9wZfridjUf
`protect END_PROTECTED
