`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NiHyR/0A8ThPmh2wfaxrsDA4pt6tfr2aiBUuQ9q5GVT/R2Og1PKWpVMlJHs5cr1e
o882SFKKJxDauzO9yAKC/j6mX0IlJLsPjxfleDd+3cUfB0bX4rPjvmn7CWU6++A+
GyBTanBYTSKfK+KP+pzwOTY5TxgiIUaKgEJqNGZUTxv2VftKVyq6Tvwf4/DlAs1Z
k0Mc3d/jJWEeL/Cawq+nXib7VcIGNurcK66ySfP3gnX79vnjv16rwH48UDfmTdEh
AQ8Cr1kUvVUPwboIGVxMHCVvAxtvFKo9wylxG0ZDkRNhMPt033ZLJPlR0F5Jn+AE
9J3i5bQeq9PFomK2Ew5gQRblAMOrydyiq+53lxhF9VxBL3/0Tka3m3D+E5oKRpai
ncXejv4614k03d8hZvlTiYKnGtuekK704FsZXTv9TS4jRVqkQyonL+cAJGpnrIRo
IFSrwsHpsKCpGKCjhSE7L5rH4XwrTxXgDPiwjQucWLp4NKp5uyqFmHYiubCig9Wn
oIR572BisPbukk5+gJ+XI5KAbylnYgzuK+ZUYk8jgnqR+7X7vikqjm8SYlyx0zLB
OX5YLG7vRD7g1miGgZDyZU+CcMNJ3l/xWxisv5iZ0TtJLTgk193T4VEClqamr4t3
uHtL2qtN6FosvTxVVL+rK6CLJj9iEkx+VD1LJJQWKASD+j0MhfuOaWp2dXwwysyW
fJkt5zOIjZHsBM7fR4AZleOYHpPgdBaZ9nH7Gn8mg+oqi5yBCODTMQhBgrPk/BkH
uxM/n25jaNU5oF7waOHqi4SZFVZvX1nXwSyu/q4iGD7AXbIvxq3+x730MF43YKCg
kxvq6aBRZYLXjPxrKwbmH0u5YARZAUi/IsP3Jt3uimaLLGBrgoSI+NZKmVGtIwNQ
WVs0pPbCAt/NZBb43awjGnfibpDz1eWjdcxc3J021Da1d3NOjd+CEt9MX45rsoyf
CxvGCkyQJN/9WDV71BIbyXj9Cnu8YfYAOQkbkXU9qS+jHf/O3Asj7uMiG60AXmze
WF7vfQNB9tErDGTcgugS+2DpypadU5xSIjqzhepPQgW6xOOiUnFaBv5LiVt6aIzb
D/9PWTEydEWFA3hFSK4CD8VSMAi1vtkP0GkxdEK6i+Bn38vEHWnA4Jlv0JI5SsUK
ptTugkuF8QAQXl9zq5LexauV2lS3hTctvMsyf7ve08ukSJpjIT82WejoskENPyFQ
J4AHWW+6a/2rB4/MYJCyolJq/O+kwU5D8ovuCJAf/W/HbKCkSX7U0zSWBkr3ddWL
KJ1jnVWDNJL9/SZABRSCrqVRrwc3TTNjQR3Y0HNifXmVwpCkCULrSPlSIbGJWl8Q
8ZDbzuitgjBPyoLqHRaCMEVuK2bcMBfjtAR9EdRjBCfLt963EO2/tClEdvPSNmzc
iEj/tk+7+DRDp1t0GVvP8XCMpJFanWl0uaMW9omifmzyThk2cgsTyFw21+G4jcbT
UrB8X+1fdFnxRRLvOxwLq9Ud03JDQ60h3UDwYZGgS0Ufkt3EtKHBOa6XuJJiqClJ
cbYkRCtCsu8A0/uIWMA9gH1XQh87SXhDrjZdRRKn+KYEU4Uxm6zBCSQXDpaDxPf3
fUH0ijutJsNmf+PV6boSM/yiFZX+9EJyIbVlbpR/Ii6+cMtxIuzkbvTDrjAfU1W+
TH/UHqLByaNrdH4f94ysitxLkoJMRTo5Hw6VJeMU+bfF1Iawxbj2cvOpcuK4Q2Q9
C1URY0LApeIDBcJMiwlFUud8JalM9miY5912MeOPK0SdcZC06SJFFukM2fwseOdo
DjYNSvws5QliNKuN7uBRTUx06dyBTBFGavySkWN3z/My0z41+X//zIdnx1xxFS/G
pCw5SG4tS3UXFphy/GfEcBe6BTBGXN1El+GwjKrss2+NuP8Cih28Wok3n2i0a6Tf
TbXvnbpUFGH/tWVmjNOS66cBAbzbtVLPD37CEVNP71qA6bjMB9iS3wM7IRkMiyOV
I2AlzcPghoOhfUAwePt2cfhn2tFbNaK8YOHO1uGg8H5IZac5UXyNpbnCORJ3JgY0
ppveR8N1mSqBgtFHrHzAuRd74dEQWfS3ct6y2JjKeyAt7syUCQcPdE5zYNjgRVD7
KTcXgaqupUn0yCQvWeQjrBJNz4ySG5+gBx6Kfg7M4z8GbHs2w6FeSYJBpW3TpQY0
lCfAn5tT09vRnjAhMV2Po5gRaUw1se3aySA7tb8j1BtSvezVqz7sr+ebulo8AFo7
BUBosMwhwNxSdcQuMXtxhysI4Fpo2G+cdxLAHSckgRqGBfdZlINbssAYgn1D5l7b
ayTCMxRrP4vyq97Ivm2fq5VAR5IT6OZm5NClDQqkhdw/ar3ZbuhFmeY2cBdd8XKV
3NIytsamLYTq60ouGljRS58ohwwlu2SUPP+AZFa89AHm4tD7SaX6X9WGgdKBPxSG
b4DIwraYzTujZSU8NJdsWFFFoxz6XKRM5BEEu9mN5N0hOaHXZ76nFB1zMGIjHFaV
LcSB1b192CqdYv3E52p0hogmxqPlOmOw4CAsB1UupHEYRyNYtablS6LFkjskqE9W
WpasLoqNSH5BCfOM4/z7ZA/3Vi2LnbVcbn0NoSJKZJ/tTPxZRTQlFP0PhCZ39+Fo
02tKinMWv4IhHz21JNMrDHCIc7r55OtGzseJgIe8u6J70Zzj+7hElyQ9ArqwPfW1
MikkXHU9LXiJjMum5LDefEmx51adZslLrkXDZHMLCm/EfOQI18Qoih+aG3Z3siKG
Du0rTxQwwmoPXtOPGPM9Y7n82zCW+MG+kTLjh7TlMlPfq8cvoO4bFJQSAzVXCUaD
BoJmvgUJ7swg4XiePPJo0RbXzjIx4sRzDbLgLFw+YTuDyVtSL9GTGZQpy6I0fIVp
BmS7XRzTqf0/IbEGwAiueKVgYCNfYIGYCNaurn+rG/L0a3gaKWfQ2e5ZdqDzRHnu
HQyi1BBLrEs2rYLa0h7P08e4HKGUcB8UREWg9OM6u7Itk7prZ0QS3SdIelEI5v6v
4b9v+lCOpq9OEiuJ9114M00wvW1cTkkvmxKy6U5IxVHcOE/mqq1whrZGBCwKsBey
5Wx/BuwYQAH1KhaQZ/+mkHxeSvgh+mAdN/axiEUw8ep0zA1jXmAheOsfodBOb6nI
weCA/l6eJkTOvFFksbr88P8jmrVCWlE+u8OYoW4rALiIeD5cThvlc7JUXuBDW2/N
RPwKJgbNMESCVXl0APWCXZcVLEFQPMQ6tfE1vwd0SkyIP3i31IIhC8Ci5bUS5c5d
6m1UUMHSdQHBw3UtQZ+i5OMPcuBNe/9Ra042H/G6AbwQhDrcMVUbqBAcPw/41giY
uq1EsqDzcHYIqZv2XVtz6Jzt5VpP/R0KYdBK03EGNPEpTVREx9eY82KBs/gHlS1Q
jqW/WUhQEvmFJBesg76lAmsxWOJy2mZarIejgHouSPE0y5ftbAb+CdVuykH2KhTc
bZv7crznleLqVMOe3RSGbQOFNVcUnWg7MvZEzz7dDtH8X5NmAfopYPZ0c9cR6TrX
4vrJb9p2ccwb5BLFAKjE2qVZcke5t8168SCZZZRpMsDXnZd/mrAzwDkJNdGRAq9X
a308gwtdbv8ZnlHHRYDxHZmBSIEbJFFa5h7SzOdWt6DiogWZa7AaPvEYpmRMXvV0
EKCZJjx6kAcXlS5uGZjyXwOfJtzMPIojIJXLksgrxIT2VI+DWNOFQyFN+T0Jt7eV
M8b2KDGfbNWVLYAm622kfQkmuxWHsDMQVlQ08Jv+gNXNALANt/dfGdXdPH5ze6ve
JD4/szs+v5dLFDQkGsgmm+pHNLARhIvvqX3wIUBuu/6PRQYlmH2v3Be1PDTYkR++
L2sIPGkBk3La9Ej32Mp1ZW2P9/qz1SJL9DjSouFfg3sSseVJ1Vde/DWnx1pdQwXO
gqAxQRqJ5FhwUNN2og4YqrMdLnTFM8jxuVThKVX6de64zm1Qh+pXbXe3+NbJyRGd
HbZ6JeSlLLrVtyP6zClo587/3MH5aPZT5LJhq5MZg/bbg0U2Fd6MLQteV4hVdIFq
xCmL5PC7sp9EjIrzcTTjV26UgDIlJUosU+hAFaNFd5PS8Cm0Bv5Z1L8XPKmNRfuF
Oakhm7U5lXPByeoi36eyInDV/ef505esGGoyJ2AlchVcrunWWPZ1Q0ZhX/UkOLQo
S3jF8/+UXSeuMBqjKZl2sd3mfned5k+RZY+sIDi+WRbgPAgvCU8ZD2CPQWp4Utqx
YTxzqJB0GuLmyeL9tY3bJQtyumpIB5XdC5R+jwJSsCzMmNB3poFIME3M+KRQeKdN
HkcA5GgqVHPZusiSLZmj1Jbbq30CwsuVUmoBUPmnZak9rhtUTLJXpAzJJhi25FlN
rhEeCoK3jbWOCi3g4ZCastOuNwgvs00lAuOZUXmMmLJ1AEgg0rduqB52EVBvWGNE
l1SgqIQOh//MMhzQBDhdPSdMQjW2QRuNdKNqkLB2F2A1CQpJMLJBX7A23FeXkK0z
EOzfMkQq8Kknmvls0C9+cnSPhEQTLiXbAOKbZ3W5IyoJujVg/D82AmVd3mP9W05E
Wr60OJ0C1CXWVhrKIIz4O+W98AufL04Ya9hg49ZEUHGV0+TVF/rkNh2YXvjoNHfA
g6hPpAZe8FcIT9dpQUkLU2VPdn4HGBnrU8uVLsT5McDx9zGigb8Zg565ue7uznQB
PJDBDXdbgDego42jwvyaVSPoDh/yqMS75cgRzY2dfeY1hEF4T6+dF7CQPURn+y9d
Be2YrNorcfVSazAVALIqyqwE0hw4agW6bU4jObIyZXFlfi+y/MLGTZ9ijEJdvGyN
BiRpiFDPBFu6IhcXFRuJC59CZBvbBKCpFnCyB0EL/MdFFKTm2pXgTW73NqwXUSDb
S6YQk46BP98Nlc+yo3kWxk6WRM5CBlx8t5HJ4/YfleQDWXk8lFDAm1i+7apr9B4K
zHrOAJE8S693tI48LHTEHC6C0J348+BiwyhTK7YUrMPdGe1gC0SKn1ubuh5QZRbH
5yfCVTma6F4fptoM9RErwVPBefZkR+P7Vn+Y7Pvy5z9/jMnCCD04vy6/dzjMrUla
4ViEn2edCijiZwaAkHi1u6aQvdozQYw54zQGIt64ljNpSelkkTHUDtoKd37plLAG
hkz7jKnhAAoCjfIwQfPaxqTKtvsic6YdLk39S1CfLJLPjr8NJPGbJtYZe75Pzs7F
suO6BQtEheVsjifByTAD9YLTtGG7sFUG1V9rPwH+TdeJhQzEhw6vXz6qwYS0+tMu
U7YsxceMZgXGGmCKw+mchCmxvY8NSWg1MoReUHXlys9B7iOUHOzcZlXKfpfhDiDE
xDOi52AdFNZxyksj3iCkCoPw70nq5mcbzC++SSVnCMendE2v1f2R4HPRUiNp1Iln
OkUin6YIrRx0ql7ogHtoIiB3+PiYVHTmCVnBs2p2x0vQ6jlM1Uq5ADZaKhyKh55U
fbJiNuz9JMB020T1AcdqDa1wWYgW2KQxcqLgeslcZPD2MTH2U5uEt8pMfEe93r//
iet7WFXeL1egqGIx/NX5rLlISwScfyWIFbYyJJPND0ydntU7b0VkdH8VXjTptPHa
w3orknwB5hMNNyIBdlx0jWjOuyFVPb5tLh58nhn8KzxkuMwia35flVFzvRwNMswy
D4Q46ZynbAxTqu2b6RbglPLQWxDqAGzuVLKW1L5VqrglNyfV43g0efSmKI4/QfoP
dWJRg0RUR4NRq3Nv6K7xgeLdCfDeeitawMW/BzPh2ckQpYz/DRclhbGpjDP2UcHU
lNzQwGYibE0iwFCMJ+6+zfmSx/KgIwNSbiyf1zuhg6eLIMbgoT4L6V4Oe4S+ibw2
lcEUZj5i3fPKOGphCkjwtWbJPKSD6anWpilncm9Vr1vlukZ38p0OhKtBaHszjnL+
oIa9XIoYKW+OWNMlgRJbDpQyHzVX5wCwWFEMbTGVZwL46Jgzv2Mdvyst4iVLHtOF
iXvMjU1I65k2qFQM2dlrBppLMoBLscFS3ZdDvZMRDKhyPUo/imzksx53P3ugKHaP
qVgVZEHLtfdF7zxuAwTfipG+jCPOYScGDam5SZ/sgb/wHoS8eCuonTdyWMXVatNb
OYha+YuWREott/3xXSXR9VPVOTvS6w0NIVIhVANh2M0/0ciHDxp6WZhXj1Hw9ZIF
Bc8EiQF8q4L/4hG12UHPBPtVqMcRWAELXtHPe+vj44+++WBuU3hepItWLHF+zaYL
gOzbbtmPdOjb0akUspGEY0QEc/VEL+Top59bbPL9YsNDh7mPTELg5mZ0U3E7qHv4
J8sshMC4qH2IaTL9TjUHVYyBBe/LLgw8qs3poPY2EKyADz0AlGnpo15BvlIbYpjJ
8VPSHHkm749V5f2HpkRDW4xiP7AA5xEBYIRynYmbEgFDkx1Z7jGsUqyjYDcTrV48
wZ4jA1g8Rqk5hQPVAeQCqgxXxFmtkwXinzXtRERJiKIpuSlkR1IFJKF+Det1TG9O
wGYHFLM2u9ceGEUPVkjQlaEumthh/0dE46oCgUOtsr64/OrNSnRRaGC4L/Ff77Y/
gI2QN3fT+TWSLXL81rYKHZt+vn/xZqJLs5wNDQPbcGD00wr/yz85Akt1CTzkRwgS
k1uHAnQSQ7bEujOHovv5+bUuZuXYpNBmocfROs6MGsWuIJEpxuoh6FNAVZFq0hEQ
VGgCViSs+iKRPAFDcVymL6ZjTR9+UOnG4HA/xEbAggqdeyUeBAP3Q9g5fBUC8217
Gb28uiCIc6iGg3R6tAnYIkO7mAF9I3vyTsF2npjavJYKzwh/dM2rCG9EccSHNEie
+aMc6B8yGPpfszcfe7tpr3NR1QCfcfO6e5N/uJ89sxBbEFDyavAdbWecF3LUdk5i
3l4ofoG6qjwUjhXtBdT5fy8kkbg7Xia89LhRkzcgt0LlTZE3YhWzP0yCIvhk4Vk7
ydpmNxRAuhQCCtof5hcvxvux1WTJCqp4RYkaSAapVnLeBfMX+1u4YiehpwHnIlt6
CFa8mBhMvMHkGQr1HIKJzwaEchiFypv+8i5QYqWM9br1UvGyh1JVshtPWv44F4rX
hgCQqwSYEZVKwz/FRJBO7k4XLNaFLYGZ8vcYHznr+Tkz5RUKW0fGjW4qYBiHWAti
dfVPz6TuzApydKb0APuBx6OCm0lcz8AybNKIGKZsHYUqZC3fvmPHiAe1d3bKyqhC
1f6v2sVTl/lvOr6UjlSbFmoKm8DVIyGyL094hWyrQWznrAZb5IuqgIxUVUlP8tVe
YdD8MrothRwTUuE0MXaVF2DB9B0DO6MyZyarhqnKCxi7PG+50XJnuu5nV09zStcX
AMMaix0BlbG/oJJkN3WQjb1PG9tqc05C9Hz1W0Il1almqs6JY0GradNRVsZwV+LM
c517Q2aNlAREpbor2DZTtFB4PK7pTo7eSuqySBAYcZTxFCpdnzoJTuVnav31n28p
+EouK2eeVa9vmP+US3aKxnaXqymaPjzeeDSD77gSvrYOJhf+QxuPyJAHjbQs5UCc
n2zhDUO6SyDH1c+nO4PHcG8AgKf6s0tRqD+ci0pVIHgjZ34y7+FiW48wEhw6udG1
PpfjsYA7OHQbhCR8RWfajzG3MuhystYIwVKSj88mb928zFRlo4MIGZRf/il5up+f
E+YLPkCiBCbG4rhCTpTyU/C7B/Mhtec9R+/FCj8LFQtOK58lyjZnUKOivpMvjRT3
urHiNrZwsrZSoC0UL+5Ufbw/XqRM0MMBypqVMRY2FAZKBeu85qFE/Hl5ddrSRrpK
om+noQqAPUNQfDXSuOZl8o4pialf/8zEcXt5IEgtNlWJQSWCsRhCVFTzNdZP3LKn
8BsoKCSdLhuFJBLxf1k3+/Yx8yho1WM/NlS1h7wzm6Ab0oI1f220M4uk1HGSatAf
7z/qWXpX4X0ElrV8YX0TfE1tzPljcguTQGvUvnC0MdyWMS4cNjw597n4/11508Gq
CTZ4AfUvmS3Ag50yvJUCvFfD+EAlMK7EZjCg+W/WCy67ZQJY/vU1HNRRUYCLo1pM
84srJaU9mYzGx5yt0ffMi5Kd3eT/D80EAEb2HqWlSmXkxb6qA/Rqj+67VHNqUaId
wWSc+H+QQ5bopUU6yorDvjcCC4KE0bVBwYmO36xPaiuld4nlBCkeBIGx9OqHeIFw
52bDIvLfOGSGL1uQaZaiIEX5xsppDFGsxaswqdHBonKmEhI4xUSnAaa4xP0DrJj/
wf6jWixuUcbxNWzHdhKoUnj/UIBMxOGTYMq71HGgLz+MW7WXoD+b96bt/kiB9QlV
9wgfkW2LhyvR1DUBo9LiRUhhUvBXrL6lTL5evnMDhLRcPjhataTR+yGSC2biIztQ
n/RZyQtktn9PZb+Ld4Ilq4ogdcdX6OOGaUK2XeVgaNJdjrlUrOi+ZO9FzNdL7ROQ
h/Nxy1pJLIsmhXPJZkZK+rDQrgcieRgFxprnEqbaQExmmhJuY97BwRF3dxs/2NN9
kmn4xDkTOaaEhJCvA8GGOKss2cntf5fc21FNVWYbel74qN+xVtHtBQXlm4DuoMed
Xwo6yd4j8zJLa9Br7qSl9K9kvb4mZtbqPV0GZVsOnRjKsD3tkQFTGX8MmgaECqiZ
UHD81iemZVTtChFX4kG4PxqPQqJoiY+bf+0nuxPjxlAi+BADypRxcA0mZX3tCUQb
tjBVm5WXfstp7x6djfE4BSe1KUR1rxOQR3GTiBSyfUHdFtOOi/cjJHxDnr1dVxa/
lY+p8GeTDKKLtwJPa6Twk19mrtnaszIz6Rqb5I5Qm6f5fexKE/+jwaobP1ydfDU9
bQ7okUp1VuwzhSbZiA7a6JW9J2iG9z2RRswp7hK5UhaT9/j/CbOhUzQAZrFSR4Pl
rGiOoDSzmfUuHZ42lyEVUao7FQyNDCBjJoq9Q3SMs9Dzn7t0nhhwyDYiCXSzsL8d
gjNEkbScCJCuP7cphgAPUfFmcLckgMcqTUK9HUmXOW8Z1VFc0HeAuEZaW8ozUU4D
9/7S1sRjAeVBW5pi33Wgn6gaZNpeLf1X2lQz89lcK+zyfZkMsnxHFdG7LQcwaH2/
LgpKabHcZ7pvBkWnaZRX+G+Q7tb8MOdrR/R95/0bQqpda8uozSkPHIvybi7QUNkg
/wOB23dJi6PzS66RDwFV7B9ITiDrffHu3Sxd6HBoo/wkKCjWa7sX9y1mNIvMGbC2
cZp5Kg3JDYpcULYqxaqunEL6Mktf6s3i1D5BBGGdedTk/A+GTv5e7dI5b7+/Y7sl
2Cd+ogwZ1kxLu+tIgg2S23B01bPDkYtVQY/4teyt+/D/BzGXtsYbNQthvU+BOOF+
cXXKX8Kvgvqni0vz6D1UiQg6eNTjKsUZQb+HG57TFLnQcgzJjBKIP2UjtOaHz9lj
+pKS4ec16U4XE+p3r9WJh3wu7siXYRavyEM7ziP6aT8u+Tgk6PQE4dXk6b6r5ikb
LAs0mLlctOdvCpiQBQwVAY+x/e6nmQJ4LVwoCWpsEuVs5D/aQaXeT7QfADOeF9MQ
cTb7OyQsAV3RG+dr2vSMQGpHbkAgchUAm4qEs3ebyfmLEz49kydfbKfMBo+2451k
q2gbrhPFpa4BCXeBak4giimzJh6nueWFUkf9Yicz3tcrX1/F3MaWckIq/L5D5YI5
q7BAvAnLbu0kKZzTAocE2BBMy0vCfD+ZRtcBcYMTOocvCVGCyuocTlDULwGfIqr4
W3IlDe8M+0mIIlqpQw1OYa2oTDnKEAkh+99EsNtthSFQ91z6ddMrcA+hry8RTDKN
R9LWuwhmWpa+Cu0kmBiDvIuu144ByxkELDC0BD08tI3vexHMClUd/eAWa3MQlt87
VNt77b+HFI6ZipoGgXTs0ZzHaaICTZ7+U7FgsdU0uUag/odY2JoNlCp2tXN51gfA
66Kw+JuZJirs8nnbiP2zkrmVIkbsNIShTifuIu5wWo9j7Kx5YI7l/UrX+ZI0BDW0
kBNb2pzY48hH72c2icMSp3/gISzmWREV/WV7Ura5RwEV5IQ6F+ZFGyZ/QpjnuB5B
CtnKFf6/J0JuK6KMMuvPrEd9/jsslSYq4mBzPMTeN9mRxtYpGEXMdf7Ps7aSp8HS
yMJimN0Ha7MmZNw87d6W5ts9wFZB/7Kg79/dJq+y1UfY6VZ0geoM4hOF7YYj4ou/
wurttpLQEp8ypgSLYhNlEeSHvesYWcuC6EETqysDvPZgByR9/A5wFZTLuMK0mSyK
aDODqxjXUsPV5pa7ZjJfJpSxzmt0Y6/Dd+ZkzY7wnZ1/w+a7ST+9cFkApw/wndXr
x6I550WpNeUqwd66X1Nmfs5NOsQndFTQg8X4FpGU8wq1RTfGMqZRvtJvNZXYyvF2
2b9Rs5kSIyThbHMDdvEkiJ/cBqxwXHLKCPUdicT6VBM8rPmWyuLQ+ck39iIbzv8F
F506EOGt1NN4IJdSYAhe5zQUikTsJtrQsjfQqYOYVhbuF1UAeqofdE2eYdZVjtgO
21Iaht7wniTqvCEFwnOaDYvMUG+uUHHei5NhuLuWCvQKxROg5/ZtqhMCjNx0WzCC
KKlrkZHr+nQetTeuETneZ+CyelbPQtecFHxoPs6/yz/v0WkRqL2bIQfVf27mXBvp
euPFSz8sNIZ6AkhcXorBCIrRAa/AlJDJ4U0jrjtPvUM0Th+kWKuaKerpVKWpB68D
jcJkiYZ4ZGlpOjwpYQyYV67hKnB9OFam3rx1YQgD9fL3UgUOWP678+6kkk6K0O/T
ljDwbNHa68W3QtI+zFyDI+7jS8uUg7Wi7HGMnnuOXxa5b1UijevwP+YlHaafbNEC
rp85ZW7jKjOL1ZWMO2jbndnv6qK1Cj+aZbu0/skI2cuyTWy7zmz9ywz3REVTB+QQ
54NLU3uhbLfcJoBKlckvpzZxeTfVvjUyXMejKgZHU05bViIhhaopgUBpjekROPlA
BQtYw8ug3IZ4Uc/WsKcUUPYDjgpDja1k8JXOHpFgS6hDySgy2TMhoxeG8aS87/Qp
gDzeyq0onTYnK4l5ew0guB1rBkk+HaQRanBHpGVTM56e6Elc0ppaokOxt2CLbj6h
strM2fbC7x4Wjwz5P6/evtQZqNjF0KiCOS7kiQr3CaQfMX0G6z78hyJDVnJw9qZy
WhXD7DN0h4hhINgMNxLZTNZmjxDTOTiovuUXZbohYHRXahPQJq0P9HD6saJot4ZA
OELnt+2wx2AGL+hUG2GEsM8RK6P8Ep93pHOx+OR2hjY=
`protect END_PROTECTED
