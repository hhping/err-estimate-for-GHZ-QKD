`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qmszOK0t437m/GMcs1z7suZDS1jP9iTc+GGQEsE7a+1ZSUujw+W3+sVAOgVyvkYK
bDv6feDGJVmWaC/K71C5IgzWJZmfmDF5DNzS3B+GIL9z7N9jkdlTdX/ChzB/zeOG
XOaDV5bpldgSVq9dFpBWctXwc/IamTUe9kEu5p/b+ybV1q1MAZ8I6vthfDQa6lIb
pv9rckq5fjx6D3W9mv6o239kSicuKHPfUrz9yEKUACWloAe5u5PvgqejZm8fr4PP
jrwQ2xIQO3tBfFUu10/F2j6wTvjP5ofYbVL7JU/+Iy6UwBIp5VB4tNaVpoNbUF3G
B3SP+D9+3/8Cm3FY5MSZJ+F/UP3P31ycZ3Zfsxy6wmNACwXJ7d7HWXKstMuzadnc
96+4wEV8/iFkDZ0foHEJf8zpqVOE7YCGrTdTqQ+oNANxlBgafbPl03otoKWNJvXB
hSxfX20qG3tBMOgfzzg8zHKWeQQYzZxA468swewjeeVOu+TIERL0/7CZBkLSHTwf
3YFRX4k5MW4fk7D8zrnJLA==
`protect END_PROTECTED
