`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yC0si/Bg9+ya8pQAuu+JHmiyofqXRxWmU7dM5MM0/2ahpIzhT5Uz2JU9ZGn3OA4X
4YtIrrcsp7v4E+utqHz42Cr22w+NUvEUwC03IOd8ibVarZp+KrDpZIuSBp9B78ZD
fXsaoPERFxG0wI2B0F/PUroMF6xVbflKrAPZgUsIweh57xuD8ZYMRt4uQJaCjG9H
220k/1/9HxW10T5A1wYzmr2dSEGeTBlWD1HYBjCgDAA5/dXa8oXtMc8LVdufgLpR
3h5nBfvZ7VHsJ8XS9cim7wMjWF/0ZHkl9EHwlgiDnlQvqVK6nmrfAbfc+jLzYAV1
lw+zp28Tt+mRRHuIu0sreUUR6oI/iTQmI4CM6GTZW2zYMwY0GX7SfN5JmQau+g5T
tSSrJceXBgCgoSk5Z437Sw==
`protect END_PROTECTED
