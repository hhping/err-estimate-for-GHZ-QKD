`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JH7XHY4hsBPY0cooSX9rzIyswQWPqrx4a2Vzor2GtZnCKRKL44jZ8eb+0lVtZqIu
41lB3FkBmyB4SfwVRD55jNDuaLOai3EFjuio7HzKce9ntoImG5vfd188t4sKvsgw
rIqmsY/OA1GMc1Wx1lyXxloMqBjAOP05vkrmh1mN5Jdl5UmpeGLURrFR+g5r/Vap
fwFJb9cUnqDKb78wTPOO6XLn6MzyxOgiZMqP+pHvPCsRN6Z16mlpZRajv93HIw86
cdJmA8gYwthpfDg4ZF7/M0G5gseterpceJfPpllS6yxKYklrbYbxqSaxXo174riA
B69OiniE+o9GaTIqgyI2SUvDIkQIFQfd7EMOS1WstYP0d6pRqEtRxHbflznSJqo8
RL5wrWfJZxqn3c9Zxdfbyv0PaqnvB01iGO/kPmmMmw+gt6I8xMCe6rEtCAxdqsOu
1/cVDyuGCF+YDLxcuh1DFMmJwu/ma8A0EvCzBhBoPP9VBu9Fb6Vh0yVQJdVFEkuO
6lei7ma4wFw14JTP0/YkIvaJ4jcs5ENQEqQ9XNeECtJbncOBKyVnXRiCMrrW4utC
QOj5Bf9Uy1/9H9yvRyuvkxv08bXC5iEknJHNaO0rEKyGnOvb54kqXyMfP+rBqxD3
zoTd3Q7gt4lTG22gOa5/p+zE7Zij9VkY48veArvkVOyW3DWjnzwYEcJjueaFWNfH
/AK2f6/rw48s+3pYQ/8svW1iM6e/9Wkh+JZvHtAEh/78N0ikKZza0YbuagYJ5NgK
wIr4h5z3GujiOpZDivY0w464/1/TIB0LMmwjcE9noY4vyVrkSf5HNlkwFcde3zwJ
zoCIwczwrHzG3msFOsrSiFhLimpwtxtOdaX+jf5U2AQjxsRR6eCg4AhHovaH9X6L
vTrLVXoy/25sOFl64aQcr6JrGER6cBRNVOjIMOvj8AXYmZpQqXw7d21iQWaHKTMw
RUECqHFxMIpPVdnD8O7+Ab8A6Yz5+JifIPH9onJ5NqGTrTAuP7axnYi3+KHnE40H
UP4qgBkge/840fYCqYVq+ElW4dG+tAJMuKgV1heoedVA9VS5SwUMmWxtcEtQZXjf
3kzLkFQiCr4wZa2vTgPhsHWpzVBc7VQlvFLfczJ6tuQzpR4L8SotflrYKDo7Kd0A
vCgZWdKnpaGo1rrsgBM+mMtNsr3P5vekRh2V44sqG3hamxCiqSkrkshbWvgMP9q8
U23tBvF1mVb79+U44TW8L9qoZtY14WYtQmBtmEzKnDorCfPcFGsye9U1Kg94Crk8
Ay5OS44erJ7FIfLQ0Wyp2ITV1boM38RncJ+6u66l9p8oPlLvMZiH0O9Gt8oPA+Nm
LCvqzx2o+KYARnU73bvtBmdy737oDlhDptMpLeo/ytzzDTkA/z6xU8Q5DD+toJip
gDGJhFnuSAypFPL5NFgi2hsmLP4aa5MzSsvf7BP/t/xYLAoaeA411Hi0epCjIOee
gcg5G5xh4npIR/aZdl4aN4M5X6G8ElOI8TTnIwux7rWv5nuLhw99W8l13wWv8+hf
CZgTBTJ7ky0JUcUfKkpA1H2enKkvXbvo6RkAONkPfplYmlppJW5nAUaIIBxwIA5S
r+HPxLK5jebFqT10YAyMQRlPGZEAyvdzjim4jcWndeWV52inlZmGi4emIS0G3kvU
t6w+/35YX4p/915re5u3ClV5kP6FEsy+GtwNV3nZPca3UfekMoFjFqHTYjh6fhIU
GpT3C7xVax3W/ih9cPD4IQFkw4sqNhHhN8Dr21jqySzrd31F7yapdQxVRT9IZD/1
vfwOQwRU6jw6QoMB0NUP2ljXzPaDPplJWOreI2WsDceaupAMkdZNsrLHHX6Md+VC
X21b8H8LRXJK+VEWCVhhWXuVh7tkojQpT//BTRiwKSEgwTapJ78GWdOJJcIp97Oe
Mwn5/ZquQARZyKWjNqoNCPmiRaZyAtNpLzznV5yVflKnc0C2GU09L/UZo0MrARL4
EkeSd8fQF8XrStgwnghvMAFKxq74em6dQ6tSAAor2lLJjdJfUlMhua5q04j3Vl1Y
VzTdgWhI3YYajEkUu44atYgp6MjQJqUxOSPZOKpqsNyqQujpH9tT0kHQs7wM/X21
+y6d9HZ7DHfWwmKR0KzY1sTCi6EXKpYSJ/jxU05eJz18y9W5RvI2nG92wKIq/+31
FX7m+i0WKC4Ob095h2lyUZ6xGGIAgqhIpoGhu7qjr2/RjR4szSYeIQLcpsCl+aAS
PqSt5E5s2KeSd8BK0h5Ypi/eDRfBu5gq1vGHYT71q9F7CYibXwkwMQ84c7iW3T5j
WqrWypa26w2bHRf7Olaro0VxguRwEJIFRffO2ZIACXIdGBVcRyVORSEYYALd7YQ3
YjylDT7BeLFBw//FkJ1xRcdPRhLKn/TjpmInMVO2e7sliTA6YaPOZqj/cOYuU1Pw
RQx67GsdGGjV5fKhWgVGdACqoJapkO3538abk/Hr09fvILx830UwkCJwhGjp4f00
aTr3obou8mpXcOCctCL8fbdPbeU1FM27gBR/OjYOrupd+4+W9eaj03+Uih5Iog/c
PKNaMBO1UiCRe8QuWfl2pzz+jHUa3hzK0X/pSrgiCxI9GIm7qWbrFIftkqeAkGUi
imvkgLu0qP+oEU8CZQ4VST8lhP+spRJoVb4VA8nO86yLzzsx17FTO8eabpCS38Gm
KlDOHBtJzLzJP+wmNR34GB1Z5L6iqbMg/BykEnRG93UZJLm+/pmshHHdq0Z/3AuN
Zzzm4ajzVbi75iurc3N0V2K08FbVxFzYX6UYxWSSH8UUZJ76A0VhwXmQXwb3pzkM
rVkLR1YrAaZqY7h+67YXU0ekkQ6/915o2Oljt+n7o+I7sm9eAes0V3c/DDFxWfRE
cUcHQabbX9egNeAAwWWRl/Le0cDHL276/qYoJLOx5ogtsSfjIGBOIWTcWwLNitKK
IhJE5I/bYknMCFrIq/EaU1coWFtzOUxHKBbub0323EBNkaTQ/ck8iB2EqHlNRswB
nNPhfnu45p404IazW4Dxo5Y5TPgTdD2IzyYAVAtp/8whYpIHAf5R/IE44+lFkavE
ChXCG7G1fDFrJDhiHcr9SPT6vXuAb09O+9202io71J3Q+ovgRWwLXEdtJaMNj4Df
JXrLgwyLTL+Srus3gc/sjGAPMup+A/mNvLWO/iJRBnOWNcZdZRW+VHeGOq8cgELx
YQa+2yH9hRVqBp7eAzUswprhTxzbGCbN2lHeKBBYUXTaaUtAmx06SvJobx5IgB+6
ITGIZSiZJ2F03se+OSzoPE5El4yQdrWA5c7/7d2grKQ=
`protect END_PROTECTED
