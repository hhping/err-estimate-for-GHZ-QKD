`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SBPhjTG0b85Y0XoRwML9CFrEH0yREb+YdMLcFdeeKKBGufOdyHn+fAGk/KMCHArm
1ufHJnx0WSP5V8SesaGhv9+AgcB7469mW3ucP1sGMV6OQvXsRRW34UxvF+EiLFPn
IewzNGg1Sz15pSk83M7XRWUcXOCx0Vr4w4ZX7FhPSzzTopKKM7z+jFrxGeQXOgwn
8ynQTZjL1Ga3tvzGYSfJDIQVCeIqrsWmjU59VgaCBqjP5//hxm0kCqplCFUko5U4
Mg1PGuuEtLvaCmNfwpV7q3NY7P+1m7k4s5lX7RVqpdDMNIS3UadKHvTXmkVirVl3
mCUiW6P+Othy4T+Wqtf+4ic/HTmjmWmGzWCO5QCRc8yiE5/mPi7G+BCY9OOZGwmZ
5o8gw0MLMVaid4qBuLJATpIGfWgpTUqCrRP+BiwV04ko+8LhPNOVhL4ODDUDeFGR
euzHyhIRmhd0Jt8BPw1Cu2J3rjZ+zYub/wKRn0OIHy69m9DetvKOwzn/aTcTJmY3
d/TcT3KwUzBuyAq6EfZwOO+NdKCsWnj/CN3spm1nUdicCrdHIHRaQCsXS11tZnUI
FkSBuJ+roW/R+EnhIpOV5/9VxF1LzR4ONKgwFME99UAzDBiT2PYCiO7+R7pR+jXa
nI+9W2qklz3OlbOqFNtAKSYsRfCL1Om3QowowRKPwYA0N0EKBXUMbDxl6LluDRIf
VWrCE2yQ+NAftZWFqWvgToDbeg0IPtTt/m+lECV5LLk=
`protect END_PROTECTED
