`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IxPmk4ZKSkBqzIYGQQbB6cEpLAPPZMzovrz7cCDotQP2ohgYGJA4/oLiRx7+hsGP
g72DheXnO6gSpYqoXQzY/NOB/5bYD/RohZqoimlSOAHt7iq9SdDRWOAJjchfLAwG
scfKkPjC65Qs36G/XhUFfFpkxb2+IUEcYKcsqUKJFxcnKilj+Po2jxNTsg/OD8hV
zXqqKKKuNvByxrOKjafVt+/nOlelDKvDzsaS5+c5BpUgEs6vMZAF8nx9DwpQIyXH
h2zgGFZVbdCrmPJPRwi70ysMs3LmdhC9haeNQvwf3VRegxbtq8Igfm61tjh49hPS
vcmQPhbYtI2mpimFdmKep4dVpwziN1bf/fYvTc/cw2sAnpSVb0D4GejzolrdNY9G
W3csonmTsoIMfaHmtCLqgyq/oKF46cPw8THFscT7GQZqeEuOrYpKLKMGrzX0Y/7P
UkcUof3X5czgh+5FAsnDr2O0s1IqB8ljJhwe42720SVy1vm/qDOnjAbjEfjPBpUM
DfpY8DSWnKGK2GolUXzeClQSpp+R36T8NTnbn2W01vyFlsnOxmzNSoJM+o7Xwhfo
TkZ0bs/Be+EtuTdLTBMpVKEmns0rFDiIAXOqfXB4miScWMYy+5NTeRu06Ju4qOV3
/zwXKpSUd944Gs+mA/PNuUy87QLVbMEgwWJDBaWlxaE=
`protect END_PROTECTED
