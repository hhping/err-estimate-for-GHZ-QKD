`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xr23FWtY/LSElqqcQMUHc8hL4Q3ljT+QYTOsX0TmkoyXnF3bZGB4DyLshteLULKs
WrobwJPRi/2A9ZEZ+oH0UKFUS0kVKsVRGAuO5rz6FnTuJN5PtL3QPWDyJa/2D1AZ
aQcR2i0R30PzOCreJ1S7mmwGXIfnl67cufJFmpuSnljiH4NZd6+E4BpQcHf9OQ0F
W1qS8ppVQy2JcCjfFfQn99UTj1DpTqlnN0OALwqPif7/l49QeOSsvA4lECiDwoDl
VfIyztwG/9eYc/H/Aq3tO+d9rV99Eljm8DpJTydPGQJim6lAh/l9nYfquzzBEIB7
/zvcuN9YZhBoOhvWFWgwKOjd6uGESPLOnQpdZLp2Gi7n8oIIBKQ6xw2GAEgf4jno
p2M7HRDsiabJNSIYghZcOEGdu1kTwgGNo7Q/tA8aA6Nt85sHYAra58bEzB0dfOLY
g0RyaFZU3bpqTpdk7/0Z/na2SNUElJ/4rV0ARivuYB4cLt92BaAiUVuoVtmkWWR5
zhstV//7PsEDYzd6SgHCkTb+QhtpcQOzb+mXy6jk2Dls4E8NiKMNZM9sCH7Tb3Jo
MLsbMA9jMKH2TpUZBXDvow+FgqEtLNL7b7EC6dmCQMs1IV1A+ITDBQP8QV/Kpr25
BFHD1nTFIwLoZ+b7ka96Hd+fWxQszFVwfcD/NSbmTheELwcMCJAES1+Y1DP694x6
q+myVo05vmkokreOGOEaNfQ4dRAX17TvWpa5qrPlDA+kRetulNn6q7+IVRQpz7R9
LgEeAnNJ/VcoEer4tBD5WF16icLxr9nbDh2x2J8uw3yHcfKQ25MQyxRuoZ9ZMHZp
gxDcHK2aOZi0LR3iztfYWhQ120xNWcLCmRaZRXLngYl3YAdfGtNpGnQ5ci210GPU
SAicq6z/2QQrYFiRSZQTV0QCuTt5Vsm7qt4Nn98yZKjnBJh6VLBVlqcnMMKvqr5W
SAD3vd6BfbanEzr4nlBwVLYkBbmjfcfhMNnvmmnvHg6ha2Lv6GwvQTufXzrzTceb
+s0qCAG6+jbO1GdEmG/qA8PtErSqDWd4qNOoE3QzW42t4KfKc49zmAcQ2mkYHJW3
MuFF60R11pQmwMoQwPSW/rdetV+kzu2oFB9MjuPPgpLVGyoD9V9kETOSBeHHHi6d
wEznaQMjJJQiiGTYZCYQ00zT8FcprclyLcFAeVZEinJwoxuo6XP46xxhKXOBGkj8
BasXaUMQ9bibm1ELxdMmuH5TOeJkTeTqse9jRFjdCYWcoQ4v4SnbdJD8lolnegUD
dDLZQdRe7izg1rNh8+oJMCICSeu6EQWIZxAJ04XyoS4KcbXXi7gtdrIix/4jeVMv
lrqEbObeP3rEd0N3UBrHfBdYPQfJ4ONLsmVE6qBw9rkLta9wgaZ8Q0gZlfwEras+
Rml6CIzPt3lMK1JzB6bJuYETNRBbEOpAaOV4LVQCSJaQ/CsuYaTAA9Bw9dqagfnW
LmojWOTw9y8nB3H9CrKfbcNfLk/VNpA7vufCtOa8U4XL6Q2rH51Ra2tW3DIe2KMU
3yOgqrYZgBvJp24i7w+mAm6Pb62FcFL6FuirkYJPs+F9Kug8aTAoO/h71rTGQifX
zn7uL/EKePNLJwLe7YbZz/XPxj8bjNyJcLLVQFPtV9hAezUL+gi2OCocouU2y+iw
mNAlgOEJEDtpPKHEU2ULuEGmKyLVIgukbLNtZQmv8Yu73mdiF1FvbqFXJWiiriW2
/goSJLmx9kdSGR33QMGzKfHSU/Jf+cQ3sZtNehKYFtTma32arDiL01YTWIh1uIIU
CwQxLQEiKxgYwnajGUdjLbmX6kWfbPA+i5rZuNLXCwoBYy+uZGDn96/R9pF35cRK
cEFXICLUjNkUaUWCbsiB8Vd8YdZYWQSdJPadY87HjCkphRqa4OYDeSFZySZM79rx
PiXG5MCeZgM0lCtdfaeLP6eypqhuUJOgBcrUf82QQ6BaMlwfcvbDp2RzaGNnKUWC
+x5qtmm4RNoIlh1h/q3gPWvtqQjF9q9euGRjHcQ2k8YxzupLYmizHNo7PNKWKUGn
3gSY0fagLBj337/k8wB8Vb7/IKTdgONwaCWF8RTvofxPZwtbzcGv2uklEex2dUBI
lYljCL8su71PIi8/Mpj+CNWG74damSQRmz/ElZx4ajov6GhC//WCXnEkXDt6sqlJ
ll9JvpRbDcprBDrzRYsamV2ooysgXQOXK/NTzezUY1ldHsFiODmIvWT1F7RmGp34
KeVKmPq8WRmf99cQ4optp7ufYxEpZOp1UociIxTIJ6EoK8w8LKjCnmPkyrcFkj4m
YRHHb4hdlzVcTNWzIXNAXP4INZYQ9/mID1HcMKDy0tYzz9p3KjFFGZqKunFuPdUu
OfJRNHE3Ifbiqth2PikzX3iOxSgcOFf/O+bjxV0bLPKlO3QNYtERqKbh3eOqoa8d
VzGXhWwQoFUV/2w9F+DcRjeLiIQ0boYCMAG2C5BT+GMx89UEUrzdLHr2SppgvR3V
ZVzquBiznPXB1ckIyN+YlwYrjKjFO2jOMOU9a+juKoATd3e1QDAvWITTPD8seOZr
HYeZotqeR0I7sKBRY9oTykVLUzDW/wFkm8jdmHHoj6R6wxYhqb8Ti1b0txkkipud
+unEd3rrNcIH9VKA+DJ+yFUfD+MC0i0IE+piPu16wMeAUrVPXID05Fv1uvd9ElNt
fRmPFD/zsEjpZD7P1y962yzT9/KbC0fODRXBPoMXVAjd6cEyEeuzPfKgFDa3SU+M
ADOKVm2Vay3LO4iY7yipfUsPSckyOkQOzWWFtR3NDt2xUmaA5XiHzbKZMv3Qe+SZ
Dh00+HQwe9IPX17X5VRhyMUfu9Iuj+5ZNjSPn/ABgg/gkd59fqu1tirJJEHwdQux
deYVv+C6l/mZPJv8NIAgYB7+DLIvhGvXsHpB8AEdjZ4m1qLpfIR+Fo/nAS2cUEvq
aqAbGAgV2xfPZfH6GkrJBk0hu7pNXuMniDrsHeQ/6MqTEH5ag4V0UKtUQKOC+5DP
zEr/0RnaBXkm1chqXyn5nwQtJzQCW2Ah+u4Pq1eu2YMqfYwRpuXgr9mVc9mgxI/o
R+6jC2AVj7Jb/DHG5yDFQT1MtaufP6Sf9whvzq83p6j81t9RwPTbcfZ8Xx8BnSCI
3/nES3shhvLJE00arhUHg6yGydF6qp20tHiE4P3X6GlXfeFTLf0jGDMmO5cHttyN
7/MIEpz825SB8qaUzPcvPhTQ9uwLvU5FnpEiU6RIrRZvQXqXE2cQv+2Fxgr6y+0P
xzJdm0dEjmZTy+aw+gkYLl53B/fH7mEmqc/J6gKdS6H4dKn9zHDnIXJE8fpRV3qf
SFr8XdLsV4vgiN1cLNVUVqrs2NAmmXY1qqMCL+Fc+8gMUlWuQFrS0MR2QBu8wfNy
5A52iANNjsIKz4tbvBx2IsTrEH0QZVkZIQGIpoQYHYlUVDCBmqbYEWKTUgddaNqn
UU/u/eKX4KkqZrn/h/c3+AiWMZvQQeVuuIfQEkw3NpWowxwufocRbrpBQmJFxe6Z
NJY6uUPBO9PQkJgPMREJl8v5NnglM4eBnffVAtzxwLjvqkeJ9RBCV8bq0oxSZylW
0kRS1IMEoVAHh4IEyULCFQYh7tJ1t9oB7t1ugz+Wym9sJ1wcb2dCdVRNSVkVaf5r
h8V1UyMJNcsYAI77VCGhCtbYU3VvI6q2D5yeASopiSWrwrt1g5cmmdKVUQdEn8jJ
3RtIWy1KTsiPCkFXgnueeYNDVip+8lFyxdMtWGpigR983hYA+9FSfEotblSrDFkg
XxtReX23xt91E8CkhAfVlz94RfuUJ24qnmWZ9UtL5hLVPuxx8XN6Hp/mfDYKQrgY
gNQcCcKgtvL2GMA70ZwzFrd13yORt5pFxfvOzcWrn03QrHT47oa24N1LWBKYYJTK
liLqFJt/BxvAJAFxD5KYji8T369CslfiWvC7UistfDfAF5RuXwBSzQcqI7LWFAjn
y8D95arY+oack+0hovxLx/bJTkSKKsoDknFeb/TqjzSnoLZGpKN0kGYrVT5Bls5X
B0hN8wZwatT85i+MPJ8EQa/e/prd6o2LKF80tNjndDRiZ1AsqVuz4kXL0ptcVUNF
brXNV2O29BXSXD6uE9ktTYFVdjXh3lDjFKMW2w/tAI/t9BDvKy1ZAjNdwB89jYIu
7TF0Ui0f7Jg4ofxGxB9AEHFJqRO8wZuIWdKNHE7aYFFH0Z/ZjnZXBEef84n06FCg
rVDO//404tLO8b8qGUV95uMGPPx89t7T8MgdTft790iS/aL7y85lsn4M0MApAxG9
0LTTOUtn7tv65aVZAN5cyQeIwqp95sl9uNZwy1Isu58bfWcARD8NlVgsto0TxhCL
++53hIMqooxBR8dQRbFH5GImTbuVwesDAH6gR+esPfcjewnUgPAmtXld0FiJogx/
M2uxe2/Y7/lfzkFLj9JJZof/DrvbGQig0vaw6aDJUAIy9Rvzf+XI36HPf5arDI7m
+0hp2epSbZ3u3hht+0rWd6MDST4kIGgqvLjybkL+HE8QtUXg/KR7ZRl3lw9Q1C3l
DHEU2/yWfIgR3H9ArBOmy2VuA9uYbJ25q/3EyFryF98KHQk0RE3BS3up+gLsINi9
Bk6gtG3oUKnV7Bpk4wXVa1Cp8Rakg9gB3pjwj50Ur7ChD1lq4YZSiJtHC+LiPdW4
eBkVKfdejsljpm8/eOy6y1DGKFJEdOYZFneuWf8OQTkwzrVlVCsk62u8KUIGEmtg
CgenDw30E+0fe+djDACvgAZCt9l+sKWPfmXhLpmtxOkEwS7KT4OL/2s/wsCZeVQD
JIGsq2BECn1ySBDyThh/LN91R7je1TcF3NlbTHi7S422WsgYwvrZNntGLRKe/afc
sA+q8vOuq9e6udpyIFGE3prRzrwDFmhTm2MCesXjCBjQxbO1gQit/zAhHV8IOBVs
vT1EzhkiUdcllPYT7sPzJj4o91JOdAqDB7uYjPFtZc3RkjaYcqnbP5wctJzGnrCG
6n0ba53BOHNoXYMfmMpCIyQ5Mz6ZIjxi8rOljswBdVsMqcLe0qOnS9VvAeKKGdgp
LidMcgzO3n6YIHJCkbEq799dq+tAT6WqXwYAuwF76IH+XiNKo44gnfDMDYfxMZo4
fB9hhYtwcRpQ/u2eQWbhSeDy/kuG9czHeVxtCYEh2GZcqy1TsIE0K/I/IDDBcrTp
HwouvdcLuF5b4QRsSMdY/hO8quMySbGA5Zv3YCOm9rPeUhTprLMBK/NNBN1tWuky
0hqo85hUWTQyP0WDnxvomA==
`protect END_PROTECTED
