`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OFLa95+nj5nvfp5nEOAW5Tf7cU3rS/WAdxnlntb99RBSOV+VQXVNUuhjp/16OUng
LXfNUbQkkHInesBl1XtSGCXWidGNc/Y90nxs3Fd4mtATqwcLCqUPN/KLXq5r2a97
uvFMa+/jvhblpw2EIApwMo+Qek+s0ZAmvEdQHyGYMmxe+rH31Ljmv9QfqXmr/Zh7
rrC96BQrkNfytY9wjI1dT2NXvhln2g1mhXtK3lm38BDKSnFLM0jmr06h3JdF3ik/
4bWpAkpsdvjzTEDBAc6heJK9DfL+Tqt3YiUCsiRs5SjIS4q220xMs7WEuVBwz6CZ
omJWralc6Chequ7Zal/cLirWpaq+Bv5jvsmttycWjpUwJN+fOxurUTWbq42HhgXu
oZadMNp6VI+FiZdOvkqRs1cYM6Kgut9drNcgufUEwxM18/lklPOuv8Lfy+xs2SGM
oGXcAqBTOhr8kf/m+09dOfkLRM/NXAgbAdqHIW/j18EdF/mXi1RWKbBDM6folhLp
SYL7mgGIVYTFlOSoBZVIQXCnZSXY9FK0yc4MeJSf27Hi8ZKdwRdxLFT+E+s22P6B
NohnTB88d3wj5vTv5mGG09Zd4ciOzDG9amqgtgWHPLWCdYZzBtg+qfwlG+5e05nB
3ndfrt7cOwDFCFDxquoEfjpgPruMaTAkEy+827I1GcADuGL0aZidbR4CoMxVljUA
SF2sGTn3Jap+wuTRlh4EeWINFe/7z2OtZSFbjvCd0hKJGqDXGgqhLnI4nRwtNg7n
yCp87O/gtjE3mOG/oNl2oGyOgxcOCQ96w4Slg7JJGyl+duVSC0tCpYJbRK0PD160
7VdEMD+4dZ75re5U4RXR/FEVVwiFtqpUm4bkxM2XzWWdnLTZRacYKFYDby3fQHNf
UWWJqCS600n6WRsiLpIDqF703QHuqottDCQFxc1ujK2EyQ8BRWMr6fnad76lpdqQ
DPgLgq4pzp7scqrvp5yYV1Q878mf+rPuqxyRtZytW75vs12YRD3l4dYVxZjzm4dA
8SYm1ZOPVY20St4W1Q8k0vJVClY0p1t6rzSeHWiN5FZ2ys4IhPZCTQpmAVRs23CE
VS0j+yM28FwiiGOgHXmkPLAuVHt7jRg2PL+F5iKIeLUxZo3Jc1i4nupHdx/6BRs6
DeTmVQCEkWFchK45tott5EiB+elkHA+GFhWx+NdUZ/LSu5q/1MyNXC7nOyoLY7fT
eo806EmVe/Z9XXnF5Ou45982aJBQADHRoCtgmNBzGixNhxXATyWLWXN8VmBMQbhc
PG/NuJhM+4DPJ5WCF00cq4eajY3eVxsmVdJu09BDjuCdbp6atK3hWs3claN3iLzN
XlIKD624gWg3TQMHIzCrmGdyRr5DDC0RbV3tpEm476fwPpbuVlHqaUllRm4prtA7
1g4fpFBaCqVpGFVPNXnIAInxLl+dpMRg/ZnjJ+82eZ+oso49wGtnAwC6+5GKhbTE
Nh3+DeXqhDATDyqEYH+FYZM6U8EmZu7cvmU3l1F+npIoR0a/WvW0DIHIZHvMn8R2
64Nt+rEQh3hKGG1bZBYWM2qMxLm9dsXjbz1QSFGL/0MPY8ab2D3hUDQOdkJpBQlZ
uKzgkjuJIP17T5oyqG3kGirDf6UbtOtoMab5BH4JS+6cA/tIwI3z6LScEHOTZktT
DhsE/OmvUXaSEoWsYZhjUkh78VcIcCDefjPzRDPYwR1zeBcvevhfrxO4UUoBbZCP
kzJsWNT4XW558eyH/Sm1gHlnPfO9FD9lhTFaH94lAEYYbPJHeX5G1NWqUwR72KhJ
iEU4lRn33Ua6rmcBSJGPZT5r/joye9cf2Kgp8ux7QTichIMRI1tgWZ4PWHj+zV8y
+BZyTmvBVQ8fkePouPYzci04Rl+853wa3buATUv5L+jzAAkdpccXNR/AxO9kNUVm
lIcXWwo0Kr3WAucvI6O2sSA/ClrFsA8Q/umvb9DvbNCoyplkciZTO1x2RsvOMZHe
Jq1dp4+UvXWywy9iymat2qbmM4AyYbjhnVrE/OC9D4SLzQmdluUaedel5DM8fEug
n9FBNSdwppiSWuRpnnZ9bVKTVCjKp4QKIqF1ihdf4cJ7RV86ahILnIARl/W8ZT8f
xUNcXdd6evMJ0MutS+tLeY/x1fZ3QpzDMNJqLs4xd5sMkLzBLdF30leo88nlZmbh
`protect END_PROTECTED
