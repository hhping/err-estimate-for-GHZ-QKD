`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JBlUioW4zq8WdJ61UmeVPSpzrrx7wFyQAdi40VjryGEJ4vs8Ti2wBncK8HuG1P3r
6qrlzs1a8ztiI3eBck5x1oyrzUYouvUOXsvkjqwlq6sveukjSmm0IjWPAO2Ce5Os
/J8PdWJdykokF5FtJNHlrovqVCOhgYE5BCmsH1g7bhA4XqpqKNCbHpLsYF90Ja6R
o4s6Hl6cttoNPEvCmlel4s52KrG6000AhUYMeKUGUnpud73QPgUnZmIUH1Qa0K4J
NHOsFVogCjhce31+Ya3S94ytbuXx59dAXWD9rviEOSIKMLWTz9HvihNb8JRrMJja
THqtsH/R2qbxos0LCg2DAw+OrbhZ03r9fV1qs+54d3hpBxkmqzP4i3T4QwCe7TKl
EWtCPUQAmn6DeS8UUruVt0bgnb0jw/UWOUxZcd9G2mjFfzP2vcTPjOn1jIVpRFHt
VHqcCbznk9BQXY+JQWozpQOesCY6NZhYYALdqauXeQE61N5UVxqaySiPQRIy8pZi
JxpXg60ou8EXOQvXdSUEmx26/PkZv+kvlf7MwQKKey4mGq8ryDoEuRIzBhyNVx3Q
sEafl7hW888BAXeffx5EU9msqPnMGrFKJNYR/DSqRg0uDlXVcl+iNH9UVNEHrcWT
ZDs9eUbT4OWgdyiQYK5zOmxTIkrRHeZDRz0JDOIfU7QsNH3Ovho16WmD79yxodwO
W2gcg435l8vtrO6vnNEKbrYw+DTX8eRbNgHJInR/yx1Aworec/7oZpx9SyALQPsp
H9parPicPhwm49/6TB5R7FMZdTMlqSbz8rLAh+b/ZjpaaAnbMmWa/nTdfJaXsmR8
`protect END_PROTECTED
