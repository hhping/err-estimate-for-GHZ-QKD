`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZuUx8o65T9zw4+xFPjv6bQw9duRuD9aYnF8OVBO2XQ6HI+J0m82MmkZyqq2wFGGf
64G3/29zdqTI5CfsuL8Ipv1+C858GZ9OSmoxsDIiBCAqqiHgk/DLJdHR3eta5zdc
snWvD/nsp2aC6RCr7u77HWT26yWe2AeTFD6eznYUcr2MGMzAF0eOHmMlrPpHVZVz
CnV3rlgSq1gFzVHnmWXwnDE9gCPGrWLKMcmU2YslZRDzNEOmmG+yst9awrtDraGH
AMVTnrXOb1tXiR/0NagSncu3hQOVLwQE4yPL+67pZb91tEkEQ/84t9h84YvH/Qh4
vEJ6BV0WMpooFVKADy1Ea7V74EX/V1prRspAhRYoLmRHWT7Gyp3IKIy5YxNxr5C0
Xz1EsFPZkdF7hjg2/lfqz/jwl18jMXQnYF5Cr82x5LrM4kdUzEJlH4U8HiIcByl3
diEJuUYtCAygqpJbRAYtk6CdovPgQt/webOlznpaf1+XhFZuVxNpREdP6QTmgQgh
queJz34WnXZp2jIbAQuRMMm4Vqj4vdyxz8rnzhR5X+K344K46kdqs+JQ52EhRFJN
SqVtW/kEE9IVr96zjBPe6atu49sAAHdsBAEvSO2CYU234aQe/wnWvw4WBJTKh8Qh
ZhsLyrKlw4xtX7YC5RyxHszfnr60+6lnsImcJYvyWWVnqvsIf6FoulKOVt/OWoVV
lw/8EgK88pf9rHTIFIWgprEKv2uKkfcXIhKgWGpPAkpYKAhnLZomxTXbHCZvGb+l
VMu9zgl52s5KEfvv5HhMYoqb9NHoLvd3Oifi9Yi9nbMoRVYV3Y7hw3whs5iWR/aY
caQyJ/ThOd3CsFTZqaYHLU6Wep0NeAV6M7PLd5hQADwzXlED9spGcO5dvv9QTT0A
BzDmL1BkGAQB4G5qLBLxq3aRzysBqjEmFFX82da6QoSiO9m8b/c3l5pc4B2HiBFb
ggSQQJtfy0aOmaW01LRRvjbv/5VeVVb9/oZUjTNUcgw1R08we5rjFQjf7XtbZRgc
AhNDmXDi3HF3zg7w+SLRQT4OgUjsERFvyjz4YHBuoNUJTnY7yWFGATp2foPXELPF
om2et+dDVBcB8qwsSj04iRM/bZ4sv6Ftqd+RrQiY/hKQU8IwYHd8If7X+XnyColA
xdErvjTRcIoP2wTAPhdy/7f/9HVnH0awajIgSepvnK+7xF9wBUDC07ebjz+eHD/5
W3qpbyVkPHr1o5sVLRLKw7zZDfEo03L/DJ+OkrHEKR/ZSjFak+RgWCxEaZeIwZjI
SpAS5SmH4NUCsTdFZFLNMrws5SRQtzYuHLHWLNzOjzL0nm1+Ys/0ltNcvqOfXC+3
jvxwMH9eQYnEVGAA5ZeHp9ZN7oSIjJSAZtluBPREBj/thCjZo12Vd73NbkuskaW6
R9yll+VYFNR8eOL/trYVWg4+N8nIxA5nMuDUcYSarNCDlYnNHIoY3ZMm3rqVImDN
aI1w/mQb0dP2BBPHFa3Rt991ypWW0rLTyqY6ZBCqwOshqQ32hZl6tvRlj6SbbJBq
ome619KE1+iWTXnZ8jYnbj3tms1FEJSLlHtWS5f0kMIA6GFAycsLWx9mnnzO6Yey
W8IkXF2xgbOKY0Js+nWsF8Qdn2HqhIJZlJT2d63zp3yjjxwT/HJJNQSKTPOEkVp8
jXwPSda3DhDZCoSez+bvbRkkcM9Ur3RJ6uWixgy8wnyVtN8jgxz/jjh0UtpbIsOw
1PiPkKxIEjH4YE4/hwM9M6lHNYD87eHk5P8mcjqpGCJ54tGWAp3zUjbvIqSfTOqP
`protect END_PROTECTED
