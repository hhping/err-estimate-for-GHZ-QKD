`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ynGrk8Yj0Rp717KFOvNE3F0oDZwxkfXSlCugRJhZAptdxuH50zIa/BfYulD+iiI9
rJ5l1W5h5oIxd0TlvyKz7t4TbUTgud1/tHc25BZzHBF2YUuBhLHuQoAjMwsCBoU9
iE4GqTHAqMFPabkhpL0TJWjqWXHpebljOd642dWaB4NzywB2KnN6v9DgosQd+ydn
gqZQndtOMbHicqX1Oi+4aKEyrP69uHa1iW+xlJP8MLXrUVsqmko/PoamOKMExiOf
BLGs8ocPNnJ/Wjc97i42CyZbUcxFvsGUOsqXLL+kTWT4XGnPXmVoejUgFLpMBrV8
QUwz/Ncvleig2s4v9KqZB8s0fi0Keey/hqyWusfz/2MSya+NxZ/UxZ9BK2GFHxkr
JFWqHK4ywKRheMu1tUA4JNz94XbbVcMvhB8aGSdmB0uddzGSXaat0KstcGbdW94L
Abzk3qLj5q9D8xulSssbePxZvrIg+XlJaeRdix3bVkFE4WyyCAR3kFOpA9N3RJgx
Gxbsv4EnbilN87/3s5zjQr3q2oCmSQc73H4y5sn+GSqU1t8KmruIDAbwvEG8RXhR
ZanOiAfoAGTqE4TdmZsyR9qG/aq8LqGkvi9ujzBPi/mBU5dm+oMJlYHyluB0Mma/
UnH4oUkV+lori8YHiOy6KnViyasTxQ1DI046tiFDgP286yEWQqAWW6tGx2w+fS7Q
EU9DrUq66eESLXLHCLVjB51Uze8oecKos3q/tYPWMUwRql86DqXIabPxE+BWNM8s
wN1L7MwneWH7HOMESGaVl5qigyt5WeC7yMbZcuiHQQ7dEltO4YJpK5HoSHN+Yn7m
vll0NwhKJHKNP7xlbUjzqtk+DUn0oNc9qUogsg1gT30Ukf1tW+UjOFBQVScwxU4f
tBOi6tlm/YlVy5IyK9QbMGnog5V3M7iFtzRWESiDw7keO4KjY+o0c8hPCYDeesKk
0/8nSH5dF9O0XmUPKB6ChGtDPxauvbVPDxwLPstxaKgacaDtphzy7zHgN9Qkjrn2
/bRlQRFaiOe8+fy+TX1SBBq1citV+4gF2KthukA38NeuL+V4KCM/SjEB9/80nUfN
UdwqAPN6eM+7V3xX00dP5Ybt/y2n3Gf/WfRz4adwbmIAsTtrJd3vE98c1YiBobwU
zhqhGeO6m+DBCTXfxlTsoV4DQ8W2KP0N5inJLYPCkDqnvrpEj86NUyRiJDa0ZstP
18MmgV0UVwcxvI/4ehx65VMCHxPTwLMBnHYEJxNy0rqdJgJUfED/CwDJexd1eoOH
EVxBT45Q+pPf99su61KUKwir6DkFMSjNUdW0d+UW6lzWwqKsU2TfT53PoSKXHwsH
DQ82JzD6/DS5Zj+Jh172ZJ0Ui2SnG6X4/36Zz6SEv+RnTUUjPZ7SOrWtfpr5KYHG
0EALYBZEXHQWXRN4f8K+lXVy+gQMQ9WWp4ASQxL+IAJn5ULq9pdnh3KUqiKEsXgd
e1zZvDKnFErRUteMueAcPcQ26H2VrLNfEE4sOI5EC57ABom36CrqhvVc4LpvQU7h
vPkFDPP0HoM31hwq9n7L2fgv1oFdjJOfRZf1NslOtj6X7IpusXTATUlfQ8GwNnCq
rqjm42DFMqX/eH4jad01dZUAUWMbxviZBjr0IfjA+0CC8kDgOV4Gj0xwPcX/51wZ
yAVu2WjM0psrXSZu1FalVj510Yq4SNeXuloOiEb1J3RXLkeQwNha4wTLJay6UR74
vbrzjaU3zw7+DrBt5nXlfKcBSCGzDsiYy5pFXixmXr/B9zKptzhH9ZkUP4X8gCA5
ooWOJ0rtFj6iFcWD8sCOJsmR9a4ni8ouShWmwel+p9BOLoF7LhGEiRVtssJCn1gI
zFdxJ32pOjLwQfg1Detn1HJnYLO363flS/Q19KXHg+epCTDKx16IAxYcuKN7ulw3
96unYUnlmfW/Qssp9xQJLYlHkiPbaucojbJkH6ROPeSFZNykZvWXn/ilqgYZyW7W
VoTpwXz/d72iZ62TEJ/5v87JIcD5iu8iE+/xtHjto/mAXuI7G4wILW4BCRU9+MOQ
BJU6ac+TWGFWvr5kel5AnNMxkprTJFVQDFUl1WdqZebfsOya+LGvWqRhHbVsz+CC
WLIc8qcIrMgtCB09nSGvGojkx0Ixtyjhsgdq05TzlduZwUnT8zF76+0I7JEYuMj8
68mrA8nqlnkVhAiKHpv+Nb3PLcuBqo+MAkzdONXOmWByv+43g0n8KiOjTxvSOQKg
yqU7E7rIFdDPFy0GlFPkwN6d0N0C1vKotpK5tI89cR614OWOOHq2W5NF5Bm8KT5R
m6AyKlkVQjklVKwjDAhz5QpUGz2SRezujAW4UtcePgEv2Jz63cdRagjE4CEjmLN7
VUTVF7Ru47Sj3OSgSH4GHK/eDqKuZSwRziWacYka5hqAixOKFqDWaKydAbq4DMK+
Szw5RLuHuk1nnNz/KimvApXfZHKE9Mqg9UEEgE0orOhstrmEV+qJwbusqs0wrKBy
kUolVW8WsvBdHLxMfKn9XcnnyrAWdLgzA8HJg9zjm/uYlnSMCwVfRqUPgL97Emau
poRBU2CCL8uw5p9zTU4Uwj9dIRuC06mAB0w6I3BY3chdWOQYowRlCtQOW6HCaDxs
AtTz1nwNQlCGtQx56ZbvoGo4GZJEYkI8kWFZWY75jqdQt2iD9EsV9JMdd4rhp9Sp
Wm093KtN6+1lK9rsZTZKrszpwMKFTRyjNoBHrz55Mr73SWnI5TlND+YCYkBpe4mb
85Fffb/v3hVxnG4/XvGWdzHaru2IaekJ2XqXACEdOqzGfPKumUVW5i206ZXOkID9
DmeA8iKvJ6Cq9ZYaGGd+V6v5S0h9CbrgFDnyUIcv9yLO908eqaEUJmT9aAoq2p1/
`protect END_PROTECTED
