`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mYDZo72vrR29PPNYJchKtZofBYEAKalUHlhrni3MrelJQeQhdWnFJwmc53Z+BD0i
MiCfTvOYAa2hDECUAkwjDq3nlZiRDPVWpVk8zs2z0572t5UxxUWLm2H501mriaM6
j67ZPQztrrVJNUAg8QMLMlWSz65Zs7oBQeDT7hVOkkzs0S/p/I/VxwfcvjYmbg70
HN7Zq4IZLU2UEQacLMh86c37143U48PJ02oTL0Yf4myPph2FQi/UgtxEy0AHq87B
tyTA0FqK0bnYY4l/mI2WZR5hd2ervY2bP+tW0MrxVvWIjBW5g4r8jEQpEwvPYx8D
J2+O389OANH6FTD7q2i7e6RHlcD7QpFPcA+dEcm7yxE17bEgXHD874APYcsT3bgV
+3TgdEfOTyGr3xaenjHN6Vmf0orgnsWVLRawHYGeDNpY6T7ZMGedrkmBnzkKLOA9
nH+ON9a4Luhe4a/zh1c7Q1sMxAf6nWspYj4yMyCeIzcr5DmyXHoGpSUWoS522Tf9
U9MTc5NtWvmEiG03aZdSVS+gG60A6maClaS3PWHiJctxklElJVq69bfwPbZxae0s
l6OtjUfEKBRlMxvwXCPXRJh3dL2MDkx+3CtxPI26Rv0Go1zvBRCz9HVRpA3bDChI
Dkuv3u/xKpf4SIU1h4n0/K556/cuVCqdTngS3Wofz50S6G7Q912mTmOOONBh58vE
5OC1k6BsRMdWkDjrcPz6WkMhsUhJ8FZUx5rMDGTQidvbiyHqFcMbtDVfNGoVmVhx
46aBE7OCo9T1vFViFDM3AmLUgvy+yyFxeOT0TpHhGWgF3uzIrYBjlf2ChkxlW+z9
DxKqdfsgbOkhlpNNLJYzoDOcP59/24O44xonFBTUddp2qMT1K8OcbpNpwxjYdqxK
`protect END_PROTECTED
