`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zYRbYi/StsYGLjx3kd4tP2KrjXaqMz5OZjXgkEzUbfXhcVWhEpTkiTd+KHIfJo9B
L75lhSiL53tw2oBIPDr1OGwtu+LZVMEGFf/aZR2lbTERVJkswGy7D/DmKv/xQwk/
XoUb5nMU/zHQBbzSXLsMVEyyd4kLWvXTua9jHZADuoISKHDc0pvzzZs7HjHrpEQs
/BO47toyDmw+t4976+WXMJpm/fYdiSiun8dhPnjYXP1B/6XkT6uVLX5PyzMF6RbZ
acbQrQWof9uF1+mAqNghxNrt8LPk7jDPg0DbOeE8zUSa+nHGzwrEkvLQn+7scjaT
unC809o9MP0sanlkVRpBzlJbtSO3cMRcsbtB5SrWfL4d3L2Jd0hn3Sq7XSAN10PT
egdb7zC1ypOovgPmtSPfrO5KzBLes5x1cwZGP03SPL44EmOZuQ8bYhebLdk13xnA
/RkqBS72WWPaXFcFVPmt3RrF/d1lID3LlaOtq7GZs97OT2pzdfb5bqi7HQxYopXf
m48L5N9Rr025MotZDVAeYnuozTeIQOwROUSuvKeONieu12UBwDhyY1SA09yKgZlO
h5NMCa3Qvdq7Ct1EkJQDykffl5H9LcOx2NC0Q70NsNdKy0qk487pKhUvwiAskUZZ
tNj1OcbARt54TJjd9gVkrVL4VNE+43Jv1OhuwpgBiB2qlgjfGxCTu6esaRfurEkN
A6rKFEMfqm24jTFW5H9PEHfLIuT6ZGr1ZK1WI94xEX4YWLuSYUX030n7yr/wWjVi
DykIswsIOoJ01nZ7UjOoErsd/rcg99dEs+yh/70UcULapnSa+wa0mz1l3qdU7AYe
y/Fhbde+QEGDJ9RwJg/el92hYoBT8OQM9HxlZ8giht0/zOyvhxdTBLo/APB/wsW+
z0b2n5t2Y0DShp9ZaCr1agVrmYCmjuFxwmPaTTLw7p8SzTpN/vbDp/+JY1NKoZ0S
`protect END_PROTECTED
