`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xJNS9L4pOJVmxIzDlM2OnodkUiCIW35/DLCQg7yKvCYUvDNeBR4oOieNYJcoaxDh
2L+J7Wklrrmo39oQlnlxl0QvVZGInZ5pvNo0T+EBb3OpK4eddHhlB2gq8VHtS912
5Bxd48uK4KmPycU/Vy/nYBfHwmsfh4iuKM7JoKj+4suq2ovTuYlGvDtIMS9vZJ5h
GNZJB67erQNgqF+qfGZv3VpFDuCC1W5kNDNWjsZbn8Zjb47IQYK1kFWcbVz6S4ip
ytcRuQhDVMWupQrqfPeu0swkTFTCqJxQ+rFDWazzkHyxiWRvyDeSmDAqjqLqRgCk
w+hDTYUPuFQXanSvcFzA+NIOjmHJJ1CgTyruqUITr01vRD79wqaPih2PAK+n1Bku
9aFiTSjHhARh1scQjYLV52oruf3m5Ffyx7fcJAfXw9a+2FAQ8A3Ui5jWhc6CVKSB
d+l/XOOTO7rYOGzOtyEIa/rGVtH5ief7eu766etdZ3Ca/+L0HxPWhj8ibYuAU/5/
SD7BjumwkD1iEO1+W2zK6TDE8AmgjEzzlJAAn74SISwvfuIV3ESkDV3NxcmIPCSY
TBGTONs2QgfUJqdoUXYZWQANlpFfn5ykqACU5Z84c0ijw2mxxuwlDwAdaEsaKBBP
i458UAgYddCHk8j6hzMzqHNwUBVHR6O/rpCUCJ0U+QHRSgg8oWJNDyNP29XooOLr
8vfLQMXgG/ziJAZB7LUFcnkLY4Gov06GErnX1cjk0AQZOprbyd/23pJxw2FpevDE
4Jtd1TWMn30VXo2TJwHaDUyleu7p3rMu/jBrhRWdnzbjGzONryyX7Kk9hjbHaakD
9EoNJl2x+/xOfNqCvj5btobADeFSGSU+74vuJxmDCZXbbeM3wZGdoqSaNS00CooB
1Vl4RsyHsu1Lz783XvlqFhZskArDH4CzBRE0yJd7r8j2hhBWn5OWCEEYf/nyMzNH
EWrCoOpdCRb3l1nMZVlumOPCEARv7ad3wjk0ZeM8y/R+Lj5YXolah/0Zx0LrIhR2
auDvzfWzXLtPokfwxyxUnmRR+FDocP20ylDzejukDxuwbbP/qEHwPpzzJaUek2Gv
qGZtLboVjqD86tzzocQZljVzQcSv43m3k/QCLEkcTz2OtCV5i4a0XNUKScGauMb5
Tm5Ery/RrsHk4IoLCJrFjHcAFcA0h0PM174aPb1Ll9o7io0L4ZZq83kf3mtbD6vi
xdGffvD5XkbOGfDsQCQtA1VE7u1DpLCSBO1usC3G4K1CS4pgG3vXM+19IXAsM2JQ
C1i2WlgJZjNbZDLAX09+2amr40qoK7ac6e3cVvgkugFl/wxqQn7R9VJl7lo6YeX/
fQDDOUbh57ilwwFPIyjXnA7DLYIz2EcF+XyA0y5g39t2RZ2dIa1sp6hfMoKNLmUg
SlUQwvyiiOAiYoqafvUs+NBASJJtIrFvSMmd3qNs24Em6859uRQwJ1acWf5WDvue
pRYgUupAh8ai3TAa/xvheJdYECLC7qkG8zQkLZyU5oQ=
`protect END_PROTECTED
