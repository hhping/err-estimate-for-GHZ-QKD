`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ucB3OW6ekuS4jP5uh80sV20UWg0a9KdojRCFDR4uTgmNAK2+e9UbHNrqREp87+9K
ohW88y0jRUdw2lIDwNvdodQFqZI4J2osOP7pXYIYWISYVhLuLLBtsoxE4PopFTTV
zDxy33MXQzULswnEq7n+S7aYERO4DXRUL0dV+GXMMzBDUp8plFaJLivK26agJyWp
qYDl7dKbrCAg02YU+Z4srlXQVWqpw6zYI6uIif5NFz7rOiqyv4ImgHhpyfDE38rk
6vg8j+KA4eBWiXvW1yGnXh95FWUxGgDlMdtoKHg4O9jk+afIQ7+FxS+8vGC3bR/f
xGmUhp4zWT8o1DxF6fnkh0YMJefNVQcVmEgAwZX7bu6QTMoiws6eECIhFN3sq4+l
AyFPYeIvMkd284qutC5f93K5ufnJ4DoSu2Qez9f0eDzmQVxhRO5wy/p/jSSPVDRW
lj8j9jOFnxJ2XLfNzDTF9r01aFC8Gupa0IwKNjgyOz9oOL81gx8zwl+/5shtEAoU
l80ZcxLhEosVQfLDuBuv5EMYYQZKOhhts6E4WomOvhjPX2P6k21LSyxvXcHm59bC
LwhsIpWuhWYdDL4kgHdHSYoCAqwzKp0sko6O30XXy6VxIoWMeYNhuSVGRXDRGl1z
+KrMSyL6UURw4CWIW1hV0nN4KHsUwtHNpo/3UMCJaV/wIbO6vxBUHYTHCV5qtxJ3
7KAsoY6XRJVmapb8P0cs32onN5q5k3tKHu/VB95FNUnya2NoXlx4yGXP8vUwvGcC
dO/xzP90WrSwwYiZx3L03pwu9vpzhsS4p/JLliTB6MmWmBpcEHvygcOKZ7zTBp1k
wa5R3PAWtL40/0rr4v7KqZjVP2Ioowcbuq4jz//vF2i63X0m65aNZ8pP7komo9u6
d5jqY04KsEyW06omJWJyZmZt7ivXkHCncsN9kcXniw2R8CyHZeLdj4NipDnpF02I
WK2Midi/Jf3UDzD8MQ8Sim5RP1uOUXFO2FxcpA//RGYId6z1WMlvZRQ2OL2gZC7G
dEH0KjpA5AOV7XZunF4QvXdn9HMxZBt75YOM0WOzTt49est942xIzedl864nymSW
MWjawbKYvPXJpSLR+raSUH7evXZsPzIMdoWHFl6a/VBHT191AHKOziVcaah3MhHH
ZaqON1kOw0/EH5pqP7jQkbE6Sa5c6z/KfSQbeXRbl5ra6QLn1t2/MsHT7QMQWdV4
ikr5PVj5aj6/4aCBXkxtNpbIgDyNpa7scypWCDWTep3jT4p+CSZURBgJ4zVbemwN
scgPjAaF3Pm1P7dUGa3JTxuBnJ2UWMm45yNQ0pWFDqfZQDlU8IadeoMpgcXnYkxr
qBu+LWOJO5AYmCUszS0/Ir7f60OpO1EZwFK8LmfzFE7FrddPGNT3YQjXwP/Hn2W0
5QHnWgH1OP3UWtrwhYf9NTdjLiIb0vRj4Cf6O2V1S3AL1moA/tl9Xo7OBnwl08Wg
nPRjAKLtt10oRIARlS0QQ4MWq0Nr3TL1pkr3pi0QuTZ8FfNhZSVEhwK+5fH7KY38
isQ5utgvBetBKvdBLlzcx6PxCVH8j1RIhmPXe639Hd0lrpHMQJPPc3FeKMbNw97K
Co6LEkN45ZcOcOohjRkXhOwVzisfoxPojOG/2ii3DubUG1I+g6Nx/X+2p9KBGZ/R
7zQYMStKYneMcuFaJDQAEFQHUmNBH35ryI+Nu+6VgvRPmE6FTPS31YSg3vHX8Pq2
1TXKLfeyzj23Vit82Dnj2Sk9VbUxzOmUENNlVU33MWAACw/IrFso5KecPGllje56
+tamLocJsrnm7Qz8CKTMecp4P37W97WOuKLmjnS3yFbwGu+CzziEFNEblZyOcrM9
vkKc1Wf5hZbIqQ0cPRdCB6YF0QIJftMZ2k1lD7wfmfqD+SpJjJRGGKfP3s99Xi57
4//XGyol6/LCIwHv3D4tvvoXjmMzTZzgQ6B+wDT6LOdc4ApUCDvZuZ4H2IO3oMke
CNEjfZd6t99Nr8OZC3WXCtW60NdG7vex1vCYpvCyNnYsJGyTTTBCqIj1Hkv2Ynf6
Fn3tOc1qh+jptFrPnpyfX6WFdN2ZpuBcSihFtlu9J+Oydh1WxD9xsY5T2WdowMy9
RdmnWuGw7LLOIg0d0aT2n4zf4Pq4QEY4T9pLduohZDnbPJpSB2KoGCI5QD2YuB4g
DAXV/EHXvzQG7X3fUXDmu13uw4gqFxqpNqBO3Mie4Ehkd9ZOfw1DnJBB7jffuVOT
0YW2EZnX/uiWb+xZSDbrJ5lXdbVvPp9W6H+P1X2u9bgIeepTWYjpAKzK7yKpHre5
ic4fxi6YAYUsNqXgdnby3iuLfhnLiKlA4/WZ94BngPZNg3KVAEHfxjGtmWLDDSP9
EYbxsDpsOsKDBL+F0YVhulw9iiZAxAK0ZVTMZB2rvOFjDxvynAWagqWQK0DZ+j0p
yU+dBpYyV7JcfimdI6n1Nb398NW2A/9M0FYZy7TwEhA6I6Zrpm/iZtdD/NKeWiXM
n2DwkyTIYGyb+S2g3BtaR7Qh2gX82vvfEXFgQ//lcQftaUpr3FbFrBriSyYYTOYX
azqNqBjDh4n+MoOGhTuBKWANhytkP0LCCMvPzLB+GKyD46x761H7ZpqGTuEARzka
jwBrX+64/EyboUkdq8HXqOOV5T2uv6TDdk2GAw/krjQPqhS3wtZ0GKbYe5avbS6U
DEnhT+wRPUOIdh/iOdDsWw==
`protect END_PROTECTED
