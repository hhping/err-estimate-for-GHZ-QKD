`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jTwvDd1FblkwQW/M1xPTAcU1nyMvtwmW0+342dkki1bEPQYXlpE1QKPFk8tNukA/
aOfqYcZU0inTiOjJ+2PnPl0czUX9cw4XN/Fj3foBPRo+5lYPWVYpl3vYB8H+vBjs
AJqbAvzUwxAfVl1rTjnnlchaXSUB56OTEa+tque5vEE6yymfIBV/9ijh3YxK63y4
cIVOHr2XIalyF4ecIesjXKokpte2BhQiWUK9lLbB6a6JED2twGCPQspGe0Sb4wvF
VQXDeLCy3fPwjzsR6Tbx/oMIOqwWmH8LrrpnZB8I+3J9GIJRZVfH7bh9R8YgRmcN
tYjeThkfmh39p8mXyydgmUTH/xUBtRzrz0UxumobiIhCzltHgQk7mrU3dqjTNV7m
FeTC7kV/k3/f7J4iklUPA7Z5eMi316xi/VGM3idAmA6D1GdWNB1r0TFfRLItyG/u
a59j8LEirz4n4VnFz4gUkCzxH0gJfax5WtDSui50j/cbvZzlZTmgu52EjStxAMMQ
Teem1IqVJucYyMzbS3345ZKg3npOHno4cedZT6qccWk/mxAZjJ1QWk3+7DDNwn2E
9YW4996LU8XYpxaERuMzS6MAxDpEI0i+lWWIn8teYs4keKGv6uLNCHXWpNKtzrMj
6cxYrQVlMZZk8+y1h75oppbeGJPL99QF5LuSu/oMH1NVgRBUYVl/GdAQA4+n64Fw
9Zh9TABlYqnp5kBCtMfvWAaqOBD2002BlyD+FlhpBLWVm8TEBxGX/0ozk8dwCO7i
hxAo3sK9kbY0Ulh9k48Yn4ucyYBHvyCK74hXIcpbYXzbXC7uAc70QGg2/XE/qD3M
xAU9O1eIWSXEQWNwU3IpO0MjcFMgEZ0XYgj0g1ec3ZuT/ghszpF4yjJfzRsoI6Ki
`protect END_PROTECTED
