`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fF0OhEbmuOQWQLuf3H+FkGWw+mgvoT+UwDFgvsRcSPuXRX7KXN7A1SGpCZ61Tyuf
qsbigYOA9MRZibqfY2g3VHZX9+TWjeCYQeDOvjvk166BkzSGmuCjwh0cX2TZXMxQ
Jz3/oU+QSUcinMRznbF5Uap1tx8POCiSytUBoUup2vize3bXd0wgG55qU4xCFrjr
hwzGqT4CpdzJT2GcBHUstYYUjfdMFmbER8vir9OT5K2dOukSSc+zQbavO7NcvFUf
Ht9L4v0xG99zGigDqeJd32cFmkn/XSXe1c/UaUgd2QIh3iZk0T2CV+NI7fny2pS4
xXhS9N1AGhRgwXtcGGEfRtZbETSBOcHrZ1PPfAguJgVyP1cKDESZ2RL3M9LepfjX
WUvBCNfC6Ah1YvqofKFuIy7V9NWi6HF1d7L6dAzoGqvFxdRf9sFT+lYXtCbfJbZm
auTfQVEIAyjfvPmpyBNoilzMYs3A8nTNzNra5eMCX0wB4XheDyRRpMnoc6YZT/Uv
iZAfDEIlD/b2a2/oRISxlb4/ksnJt/9wZ2O6pI+s/gYZ6HwLbdRpSYP9mhFNkLJz
BGjXR0iaGulmJyfhVqldvL2ivL+AdjrvbuqN2ar19+ZlJWyDcCknpP8IInCMgKph
ZZJ4+o1Yz+m4+7RnyqkVBcKgLOvU1xS5HuewvIxp3tRXbr5pHzfBOzlDCFjuXnUN
Hd1iRMfzdFUzso5azfgHlIH/nxDkVdnYkSMKt6i7LAm1Z9qLhudajvlYU1ea+u5t
/Z2AuR+sKwhdDgfix0L4QRx2FxQA2z/haRxRyvkAa3d7P98rqpRMbrkMxYeKjlv1
q0bguYrFitPi8FhsDoI9sZUh/5kMbsovFc2PaQUDeiuYNgic6u3xTznMxa1QR/vV
PoF58nO7XwtOnZAYbdw/iBDcxlW5CTe6t9+Den/8YrDO0MPx7r0kwVnuM/3Sr9ZE
mGav4JGTlwtV7yU2R0R++T3ox7m4MiR5tOdVbonzRTWiCDSFOM4LScPCHd5Gwu93
CFVhHjMHNyNqlp87q7uzO1TRIDAoCEjySPDHMrUAMGTVw1LVpehiWQGlxUuyJQvL
ZiEj8mWeXDfUl2oJlL7eUsNGKSXEXvP1tkRF+s4fzQmQMYlC50EH5B7FiMjWWddJ
JbcEHW0ZkEHgdOhozt7ADmQ8+61MVCNrPKZ7iE730aYa71yyYdMwMVJmv/mm/C2x
FlbIPXIVGRjQYN43LQEgYvr6PZdUy1xx27gJ4DJZBM0p5klq/cuyqypYCb7hebDH
LPj/P4AnGWmo3R+Bt8rgB8MYqzaxQRBd2FZvereBnE+BC6OZoW+1I7O0SQ486Ial
FQnfkoCruIj5oKsj6cXW5AdcAQzhEKUxzIMk0EwNuOb+p4ENVflKsEaVDjR4B/M6
uK2p6JE05Jyv0WV32pTFFmg21cl0ZO/75YJLBwVfkTIYhRwUdfqQ9CslkzUUNc7Q
a7IHl+EGKsxownhMQ+8LtlQamZGvOsbfQDTmJU7T1Imne7X7f93PIBrMoY9fm7+E
JPo8T/uNdyy4kyF/TUg5jpvj3JOY9+XBsBOUpgFBC+QcsWeZrEM5f/vORLaxUa4W
V3gXeOfyQbiezZYOwesW+Q6D37hP/rNGr4R5q8CxZ1EqvIP6qeO+74m2QXOWU3hK
srCA0JS5yvC2m/mTftE0pdhNgOnS81EFgz6QyM8tYF0O6lRSzOoviD63xc/zXCvJ
V58B6WXBGERT/QFhxVtA6yEV7EuuwNqt16yFXLHO+t14pgriUDjjJQhXmuqWuPPx
rKSuj2QzuEvBMarjgiryUoWBWZZLa1+k7ANedS6G+a+VDSpWo5NALlFdtJaXMxTV
ONKX+32pLtA61Z26EHci4/cs19a4pS0rjk8RMkCq/nuuiQtNSvxyebWxv9IaHINp
zkzJlpB5/oK3PW9+fOqysAIdc0VBfetTcLfsYy+VYenZMy5vMlAtFfDl49ojUNC7
1BTD6rRHc6155xO3ZnlDOlxdJxBMhReNJRuMegjRuHrH8oy27SqxgFjXTL3VYld9
vVtfDTV7OZ2vVqZMgTOqCsu/0zfnK2EZUtQqmmpaRmh/pnb4q/SXdq9r+8SQN3SJ
/VXH9NS9Yl6sf8k70KpSU7Rst50qHAthGCoo3gMg/gy1RmU0aL8vPr3ubukoTFuq
+vN4daUVD/t8xFCprU5rxYVP7biaEyQbWyAAUQ88TcTr5ADRsi82I6zK9RnsLiRX
m5nSGv8l648NYUz7jQMrQJtDS32VboCLyLJB0dNbbiqV+q8YH00ch935GBys14Eo
9r0xjexlfONLtyCSi5NS2rNdUeA5stapM7vozi5NF6OPV3MNF9hyFCGtIHrX91AS
00ysqKL+T9zRUSjMukXufvxKThIN/MlHQwNT5Cw1xp/fiJF2TttI0eIhygfHm4Ji
5kUfbjfMXugqn56YX/K77AaHpFZ3rEW8fsvjT/iN/dNdKzg19Z5NemCx3VDI6oZx
78vPLAb8RCEiXnwbKu+iv0RzTMD86bLmPR9DOXEFtJSxi41jQv0Db215w1gTXFrk
RFNtu4aXoPDcuu2Vf4d19/ijKtcyiuzZXjsKiyQBrrGE28ERDJ0JHbTd1koOdOnZ
4/xa/wrY34YKYOI3budegitlrUBVtQNMIhPpc92nxM6GtcxciMfHPJAZiKhHknvc
C55AvStiUPTojRTcvcDuCeHaQk3w3QAFi3mKZuBJdrYTvGJuvDQrPyjzbLd+0wgK
wXbXXOwZCfrcpuT57G4VSZW0/Vv+Qd3vF64uP3XNnXBpIjOE/u0T1En+l8Q+zyaO
bI3+4XFgdtpFd62xpCWqqZUmMqtIMomebjnSuF98O7tRDFliQ79cdxrPSbdK50M7
RCRiNOtOJJtuxP35gxlDjbpRKT8XF6nlYqxPbfE7RY6MCMsQTPU/CjGCMVVIcefD
FHJ5u/BMMIa0iulbg6ii92PMCoE8LM0eeRIdbt/AJZLOrGg3HH/FzN//Sdk3QCmU
/dzQ8HQwK/ABdDwZrI+NzYs+632G5cMv8TqfP5vX2LYAV2UuDxmJpsg2qtsMBlZH
j4HM3qy/ccIooYPShyU4Fait+hCmLPzmCwjJHpM2ZEYt5Pp88btLVYbw6ARKLj23
MzJEQwHQs5uatk05EtQgf5BE/opVCC8kRt2Y3Og4MnpuhPaXNtpQlnXoXfL1Wz5c
tZoczNfFbLgBYlUbsQdUwqb8srJvctmcB2p62/R6wMSJaCJw3pkr9nShvE2v1fIG
YWUYDpezSgwpH3oDDbpInu4R4yfHMQfILMfwQLloGuK8mrn+gertHg6gu+/H4lv8
P3HHXreIeXzKfh7jAFtGaLxP0t1WLT/7LqOUnr88c1wljSh/5ybXL31i3TC+96h5
SHI4mfE3W5swat36H01j9m+bcg2UD47Xn1IovrXj12/dyGbFhgBUe/knoB1BL4vZ
C7eojn898aTNdUcCI3mhipuMDJAgiiKRdM5ixmVuEDJg5/yEjfGo6ThS7iE6DzGS
SXpl7a978fnBfiC3lm467hq0/ZSYh4SLYWDURyw9axT+Ny0zQwcradeIzFBUWPz5
E5NUR/TKWQHlB81YPkPJpQUjSiLFIfre5M/nt5AtBKvYlHCF6YqPsdjoK+1o9VmO
8hlBwaLtz6UsAcNU4H54wfSYK2ruL2w3fbkYVqu+Y21pGTv8taUjoJVF+dGOMDRD
9wpiJwzCp1dVFoGyx9NwkGXS2TQwmEX7YU9ECOwnfW2PbRdE3Bo9xTevg7hWIL53
IRo31rJFr2BztZA8OpqK8QoGjo8mdhwF/0+OY+IA7LHK+TlDw0QEItwv+4K4t87o
/d3FUAxeQfAi09XDOWmKjXgNyG5JXyL4bEfKRNb4qfX6w/tc0y95wUxkSH/JGBaj
dwY8cgX6PQaE67Eq02ydIxHLxvNDp+kXw+KymKp2Dto01xqvjr01GsJ3T37IpAyD
DjE+YfgnnILSPSgg7dTfGKsmxZJ4Jq9hTms74QXQGfkULROTKzabyg79SnFVwfmV
qoqjYdEgpjxhlzMTBiGp/8+MQu36wKgOKmZKMII8PvBRuMQOrGvpmzQz9Lw+OVlq
u0ZvEBcLcwkSfRHMz7/tD87cpu4g+JfYvX3tiEfq3LmJsfo6YZj4yVwop7CoWWzr
YjsED9XJT89fMeeNZ6X/A8pTED3DjLgvX7BmM+3sTAKEHiF95vPnKclyWFC037XT
BjkrXAx3Mo+xfiY8L79GhqTWikUlou2Hzmkesor6EQox+U5dRHYhhAMiddrrlYGW
2kxVCWPXLMfs3AyU3pxsjmW1tK2qE0qLZL5vrrIpGFba5ssvEzKvFxNEyjhOaoUw
Unl85ve/OZJG0ece2hNYKXUspOO0KjFP44MR70gTXZ61n/k9BvqsrckzzCAsjmLv
8mrWwkK+3GA7o0CUmM3ix/EFDNr/zb+/8OJ9BqWkFfGFc6f3Cw1l8qh5Ve1cazWe
iGWJSFtk6Nv7d/P8FLkW7FPJJjUbeMpV5q641mEdjIIp1hBoGOvg4Xwi14UOLO4V
L7tgUPVL2hQhNkzVgtga3EQWfSBf+v41zGKyWmRXwBuISxE9I6hgo14XzuySWc6N
9C51oCU7/Kw6+vKxNLiv0SL3gvAljX+SGC32YdWS81PAquWA+Ig+z6BkC4JAVGi4
ryqh4MQuN3WunuCZ4rNSkJEiui1K1rxTtIem3CQ//xGMR3/t4yIf2sbGn+78l95a
iNrpafFSk1ww4u/8JUPHNJ3lZOvRi8lcrCHtOJEFrjvGFBhEZLWZBWKNGc1vFuQf
SOCk5s4ZQfBVXEPTRvA8i9LsQ5hrzBNhTAmhpAF6G3IsbHklkdoaQ/lyfiCxRmvJ
K0M9XcqP2qnQWp63XXcvh42rj28fL0C5ULVcOjZRXpo9EwEW/tXxyzh7FVdXMhhE
ya07yk7YmF0YJ8E8Dd+zFCASxFuJXnrznLjAo25usH3Cixyx7bKwka4+ZbJfUtPw
NN9RLYJPOUYz7kG6GIpIbP2vD2Aq9HOWxiWa6Rflf4U+NuRJrqprlAjFeUfhbs3l
o+9VhKl9EHq6U0Q9Osu3pW3TMUUnGcpiK0XrwNnUhhFGyYwyoQen7X45T+zP7tgM
1VmJOBPYYkHrcSn1nP+ldTeOwp4EH67IczvTSEh0e1NMyslkiddyJMzoKSNOTDDD
cxCXnaWod1gy+xnFfgAC12V0oCuQj36SgBphkDcsKQctT4aCLZpZHopNUujtLIN3
jE7RMO9JXt8hbHfnTeSizmoyMJy1KguYhiKhYnOppf6Lk9AE+g73gJfwErhoDz92
Zlkwi2cHf7b8Wm0a1r+A85VXTVTfNTic93ADzDIzVJpL91ImDVCC6AbR79m0T7p8
debeX7hoy/2W08ab+RXKwOZ4pK6HJYRin42fWi5ahl5QecAStvdGd71y+aMhcJYV
RVzOrizzduER56LKWlpk+PK5IlE3h4fZMXfis9qaZ2rwyv6dPUt1k9GpiMzHSneX
fpK0i/KpHdMWidiS0RX3Rj9QY6gkRix86zAxsGlrgGXg1FLAwB9T9mM7sGitT/uQ
ick8Z0i4afa8B7gMvY20EXdS0AeU3xUygVJw46ftTvttXTmV7WpOuXL82QjVY8ib
IOkG5yX4OlsCs93G3QtKH/lvcHP0PltWs9txTWgR1NVjh+lhft8607+aHr5TJZM6
hO8O3TeG18pMllwdBZPFus8RZvDYdIwstGqx/tPiyrxGGyjks/aijccHBNH151DJ
q3wNncw3nUj22ixPpzsp5b4/uPmvi6wGaoXeBSe8uv1Z8DEL6OXmqIpozm+rqElU
0xSs6uQinPPwxJh7jX0OpZ3VJ65Kz1vLSydaJQbot12yI6vBKjSzv8tDM71TL/7V
BGrN5+mpRNKIHaoY6GBffQ6pjkyg1bF5uT+JtXPpT8Z+PBREpcZnWiE3dj/GiFko
NFMjYr4enZ7s3J4PozYazDvEj+gOv1jWXC4ghtXtIlXtSa4OgtI7KDBuXABAlxLV
i0Nh/Ovtyhvrrvfjk2tgfV/SqShyRc4AjTIfGt8QSgMpMzIb0LgQPvkd0gQkoQZ9
ha5zsjlUhHy6fwFJxICIqsfuM6lnKYlCBe+7NdEvxrBCynnTqw2mAdS4zbnS67SX
wp4IuIta6XEJnmtyViH9MkYs/SDY1m/wRKyYVDrQnhW05SkAJuV5u5oj239+/38X
w16sJ5hrpLv/FS86jJDuQ+kB0L9Ipop0nyGzhJeSSwhPSjLCPUyGfNx9mO7U5HPW
9niDWN1wkVz+cHknAw0GPXlB2swrXFdzLyYhE1m6lOmkRM/6rnklpgcftIwWrNZZ
nBzKORmOWcI2IY6M0A/mitS8neBkp1lkQsYZxHQEeD5BR+l5KbqTQRSUUWQHjLQ6
l+EOwD/UDI13K2vdDx3gFg==
`protect END_PROTECTED
