`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m2e6DqCzDRzIHSiusMsDz89vud9jUdXQXCTTqwnLDIxJcA2xw0UpqX5YECsIwBCy
DfSgSQ9PQ8F8xulj0GeGeO97Y3kh7hOZcxHoVrA2jnt0i+cqqRpXFIbVToR5zr/g
SFDOiii92AbA27DESfGSItlSUPSgP+HhjTBLd7BH8Q3XB8U+BfOALxiAstx0jhJ4
nNWInZP8vzj4GZIMhYpIWyqEUx+v6Alygn9cph7GRBD4lGaclaCD4BtO+Gnqr2E3
OmB+kLQ0j5ZoZkjPOABDhNiYJtmsRjtdOqbEm26yRRBrIpez8Mk0ic1M3PsAyAQ/
8Lam145g/Fkxc1hJbcwCMRMBmavzJQmR7boQclIJ8Ed+gMwcP8B74r41Y+QM/XgD
PWI47tVbjVEJ8+970QNEpVb10eMF7ZeIb1InvPaNv8Qh+nhD+9aJZMUL4zjmaikv
HpW+qC4jOe3Mi9/6C0WLh+uDP9Mf18YYb5ddEMOTGD6+OxwsIWp62KN0lHt544nb
m59fMWBeuZd2nMZPGxtrZ3ynBYEmr0gTfGtX/HFsAl0VbpwmMfzzsxesGHqG2epO
do+zW6eWCEkZuQgdy0pctJnFOaxgT3Rpp96SdZISvaaTAgHbpQorAW0nxbhY/Deu
drSZLavaxh+Gm181054081U3o1Jb662505s6ZqXB5J9aC5czrIjXhLw9utpIsOZD
Q16F5orSABp4iwbauxpPpByDD3oR2eEO+fMqo1orelMJq1ccyh+UEJFjinQxMOL0
hu3iZwRoH8u8Iqxr2yEnEk85Q93eG/yDIvl6LKGGNl4/gH0BCvhvtQ4WkZ7FD2H7
LrhF2BKs3DO+3OKzcF9TORuWaeWAeMqP0JaMVseWrDVj/FKQ0IPypLz11pW6+y2s
nNA0z1eqdkKvMiZTgIC6eLkvoaBwY5eFBjq8Zxx4pxiPSRuyfyFUX7EpUbfwBsRC
UEHlYPfpzkgjrUk2w0TI1GYMG99dUSUadyg0eq/oJk5J0J/0AaoNfBAwxiDU6iNV
Ft0H9osRVQjkhvbJpTVrO5fAgjJL5n+hPFudYmxKJjHl4TA2lws22WTFHbvYSe7n
RoV9soM7wCEj/jbmMbJy42ccvjtXv2niLmOC66HFVCbnY7UIjOE2c6Ub4gmJijBH
iqLabMNZOhdDOpkjOtkdcZfrIWannGf5K1ZtJ9RwPD34AY3trAtH6hxLeABEZx2/
TGWDlKpinklvzA6vcq1HfsvEJW17DL+NVusT13+zBIb9dxxuyuY5oA/faULYb5fz
9J6TgoQhHCedaqxTlG3w1KW+pAJczkuJ25szIVKDPjn1JBITDRQCd0+tf+Urmzu8
opNr+86o6maSGCIEAqfh37hQmKfBqXaFNYHc0tJPDGVSOfQgf4kJ3yM4ei7PRyip
VmhGm/b5R+QXlngX4sC52JVdCBbaQQ1ipF0lguOm5Erj0n+2spTEo8lJOOTJNyxY
pyS3UpCE+AWHIv1QY8hMY+7xW/HV71RClTQI87lqTgw38NXdp4329p7pxms1rgAH
2SMdPu0iIaDO1MVvq28PiBUQxEhhy7ICzbHhZrxJA+kgg0h8wgaABWuTu0Cwr2hb
hyCzIEC1jTT99RyCz7AQcEAolsJLgNCVn8cmbD6i7P6w5xognSIsB/ZYpaNzZ0HT
6HxsjxI/l7bD3RzJY27XomJ950e3o01s8Za3Bkcd3jBDNkFWNPoaI60f8EJf4bZa
WAvVn42ftNzlV+mh0TSd+PqCVjpl2BpKWDpeH3U2xWrod7K9T4oA7k2B8N3Hnpq5
CvdJ47YTLQmrAqXFkiwfph2v5v+rL65Q8MAqPeVErlMr5AY9E6eG+j6Q/x1WMlEe
1GRe1R/gFDWOgt3quhvfVWiKI+g+ajZ9p7Z3+pzBwgO2EBlWuH9d9Bb9ToueCuua
5f8C9scervbePx/l9sYd+QFp48LS0ugq+mttfpZZ0rfD4T1eZ2JI6HJZsvOyyzp0
jADYo1dbWyFQD+QpYQJZhvVyr1Rb8gfeNOUWXIfOFCIEi6mgl7OLzNjBZj68+u9C
c+ojeDmmdqEQjrFHxbLPEWFB8Mm2ymrFdb9Y5zq44Mb01/5yg9Hs9fy2dvAxRvA4
kja0Nwasoje8mxH4dmKIy5Xj3SEdfGQJc2LcZPiA39TZJmia+nEqu3JBPBahhqh4
6AZLSD2lHNmWCwgsda7k85IPyHs7CWZJhTuoM7+smP5oM7eV0W9U1kvrtDHddck4
lz9+C9jmDhmQFOQsO0AkhFdYO3Bksy7kfiKcOCeeFrIl7Ec1PdxOFL5uVXRWdQN3
yvSfKSSzDHso//FiWArnacOHsvFHS0oHzQQvA4tqGi9hLFwGKQ3WeOObmP+PC/WV
Qpl5UlqmgoNE0DbEJuGMu+8JvSndpR4WuQ2KG2PCgzg/70j3SIre/uPHWMlJ0gu8
fj3P/5chQe5/gEOrAbXl3H7UnX7lx1xAp88SFlznQUHVaX9+JyqvYMJ6Ls0MeeYh
GUWdgqqO8OkL4Mu+YwdwwlFx1DCKKViT+ASo5V2KjOwC5ns0bjjZ8znWtQJcLhJr
ci45F4RlIj1O/qlJ3+zGfpKYsPU0t644rtWFtpFMxig77dFyTLAGX2RkpqKSwaVB
aONepswWM+4EY7T6wsaLUbwheo1wqdsQKcACDSZHxPqJdkoiaC4hSjD1okMehjdW
GwNPXcuij/9MuBOPdGLqzTSVMhg4E3+m8DwRAjZVr5uM772hEXJauEMTdhrqHIQg
JHk73KMIOPGwPxhT/EKvory4nQkEsKi7SBdfHPoU6p3apbpW+SJmMkc3d99x/7r1
D8kHYulkMkhxxSdhCXmgnssI+bQsMvN8Ihu2NaciYS4athpGnO0OTzYZx0y9lVZ6
8/ePFJDF2N1MNciqq4Obwd+omFGvETWQv69gykIr+FHVoy+sbNxOIIlB7qbWbgjc
sy+YyxgHFxI6LGqNGtRE7do5mSr26fOGEIb+PtK0aW0=
`protect END_PROTECTED
