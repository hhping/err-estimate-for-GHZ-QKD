`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ckLaCe4/2mOKGT3wlQUNC9LACV8d6YD94UaJFAlwzI0BI8uKSXlDIozkIpFwVUn3
LUV2/ajsDDsu1pWUrtzgTDmAtHxMIcXR2g/GQYJZOFDOXcrVPFWCG23BvBDyj6A1
1L9ih+4yM0jLcO5dbtuiEWmHGiW+1QmQA8TkDZq9ihMFRnfmiUgsASm79I26mV+V
uwib3J+TCpt22ceObVZ1N3Tdwqc4jCmKcCNfWIongT+dderPd22/robP5uh/aI8I
+JgTowmdzPcqXZucTOcXhgymcGtW5oNtFQZ/0IETFWNjSwcayVA3LlXZEdtTvUOP
Q/uMYC05ymf8yk2d/Bko3U1jbFNI8KZDjPwh8rWX/PvyyZYCBtCBqUhzPgt9n4tL
ZpG24ekTbMcREZ7E4fYK8OCohRaY1ePAJkP9fCp87IRIxJG4UX7GMUEk9pP4eZty
fRsdZYpaxbpnFYMjDKkd/13+hA47ZkflIseGceNPXNY4bOMsw4gytXI5ASnC3ydv
5WYzXXcXkZjRdCS2MNNMbVOVA55/3ClLnxo8qIqpzJRSSxJsWHcEqtUuF3Zzh80Z
6yzgfItbvHtH/xbZPa1v0BD+TMCnof0ShQgKosGy2LKM5yewax01RsSH7WL60Cnl
vvy/ciUak7of3aQFCK/RgLuCMvPYGuT8CFKjacMkt1mhtiFa9XBjSjxoBtXKh1e7
3r4XqRYQjCKikVrcEWqPNKXh8Zb8rwXo3p/eq198eXYjROz4p5aTL0ez1XigZO9I
BHTlpVmsNEtHo0IPzhmrhLvHnq36ERmUSkXsDmH4Nz2cYpWmFuWhwI5Fmqy0Q8L5
tzGURMQMhc6nvbtAKchKI487WdSgAMSlYeoAvIaPNQClZMSC2vo/GvTIxDAuuffZ
EYP6ssizVevsZhGegGudxUngE3N8akiqgAxcNEumOPYJzfGb9GOckIyMrbA8t1C1
VnksAIXh0dB6NcdUzWj6EbbGmyfTQUKj4csaeYW/L8KA9RE5LWEifBseQo/p0VxB
RxAJg84Y66fOMqae4rtLDw==
`protect END_PROTECTED
