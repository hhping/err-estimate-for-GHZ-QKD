`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L4T6WmYVF/Uw2AkGQsPfMJrqDviHcriko47frDjCvZV2WnbcdvrElc83JvLZjaXp
qV/bVAqt07JZdR09rfPB1t3OG7XiA2hxj6bGWas0Q8Y9Jv00gjGYYncff9vIOYzr
n9UGKYf02SPFfB8LuFHGtSX7ZolfE/U5hmGBNwxKJF09i9jnlW+To5usmbGLjy5s
+bH5EqpKD8F0LuFgG+wJIAbvqhxYOtZeZdqF4ZLHcbpPwZI6av974UbSwjaRyxIB
nrx/rc65X+VWAOLw9yw4HrGheg6htCzLMQbQjZBnCYX0clwRLfIu8x54iQ8qSZa2
V8W4buem+UGUA98O6lyWOXR4dJZvnaFVu8NP2eBUO8vXkwF3enjCNe/NG0HDmtxP
dl2lNRLw02oH7K7mca18Qo0jrb2/gQ0VdUxJxj6U56ughGG3Y9bUQVB0vQn2cFbk
MRXf74Qpt2LOvLJ4O38hrUBb9RJMc6mybSWcW4Md40BQglLyN+AGL8HLo+jmEIF9
h/hyDmFO32kVItsIN9LBWjlsEFwwIgay9jIPgWVFg0R0TLxs8JpBggM+YLqUHaCX
NVpAT+7vuXdaIGm81IbeKkqu49mmYxo4FZAWxYRZDZze7qjpaLzLtl5i2BENRcaT
X3PvFxFQhWX4JCh+B5BwSgvjpSdJybqaYbyVMDtEIoyblLBsJzUHviHI9wUxEjeK
O0LW4LXhyRAqvx5QHlrDINdawTsOi5EjiRpEQND5leLhIpFkE0aqe8JC7doVc1Xi
pe6CB/Qd0c7QolRHN+/xPV27TB7TaEMmB3Yw1y6xuBIS5eDqcsbvHWAf+qzql9M6
l+fG/yufy8V4cw/XjlypH7JWikYpuT4P4E8BmsedpiyySn0K/OfEDCSPGPF9dR9c
s/rrMZyrQMZK7DKGmCdWSQAGrpOcu/2eXrrFPRgGsVS4sfind2qOGWP26M0h1nVn
K5V1WGDb0wFcIJfVIOtb4bHweLO9MDRxnOi9vlelgsDNqgyvxcmK8VCAGE+BP0mZ
VSaqKIqnT288kxr6W4alQqmiEwvBuQmFk6x0mDVtmpbDPwjZeeO8tWy9VuufQzhe
hDcTQjvU0gGkeZaXPbZJVxllJrMfnAqdjExKO5mKnLrntIV/jxRzUgnXZVvndKdK
eRd0CpgaxoC+NlhOfq5vdsFr29oyJgV5ggab5B6Llnk+Ba5bPL6faeaNZfGGsMqk
hHH+/7+HsP7w3KGoUXxkNA==
`protect END_PROTECTED
