`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1OREBpdsgOITDsQL3UWl5Rxfgyqn/gaLVHFrjLYuo6/TkixaHrQ7rOurq+5o7Ajn
6YQlTsBfE5ZENsIH2moX5ZJ54eZShrVJp8MeIvrvlMNl+kxyl/LQErFEzA21ckCY
24fu1Wfa7g10Ths3E3SWka5VyHYKyd7g2RI+jhHF8CLFUHtQ/yq/wQ0dzKW7zHJi
vkjm2sFM+z7bHewx69XEdU3OrIicFEUzSANSCAqCK3X9EiWYqoCbeKVDRUr+LP6w
AFE6cZQ9ipI4soTcjruCmxOz2Sb6vurwas3OiyYPCHSbzEUuysWvM/lnNrDoPBnY
bf0+0yTJI2dZ1HURjF4S8mhIwtTdempn/UncInvDp5mTH1vEgtRnmCvk0ayTH8KV
4vnmqcuGsJwAQ9GCC0vKjIgWYW1RSN71LNd9ZfF94gvW76XfbeNCONK6Tp8DN/9d
YqpD3LtZt5kI2k7LBwfVwNaGK1vIsJFkO9sRtuVllDQGwaVqIzfWXPA83lfEUs/Q
9TdC0r6JnCbPW3kiC+RqYmqLtaSL94n0KV/Jxo8BBGiN3/dkgHdni5luTGYkES/K
ULvvNcVeafCeD0xU/kwKwK8PY2UlnNrzT5tl9gdu5yOurmYu8w9sWGW+QU40SqIA
JBmqcJjsjsoLg22IEsvpE9QW8GqK6n6mNs5wfkGVAcHCj+vjRmF5nP3hWiJBxEY7
8g5s6/ZFXihoDmoMLlzVB0gAjjn4y0xV63uryc3+wMdCiht9VRRlS+ZZazCl5bqn
sCWGRnn4pSQkouQ+tR0AJk5UyIE9tPYuuHQn6ZwaEU0GHYmroxWSxCFr+7ZqBXHc
Sn3WevdE81ZkEXLCucCxNYmXzaFriqIvbXkkFLRqpQckf/hAHR2MeQZcuJQvG8Fz
c2ISyaLEXRTelVhjrM+PK1UuwBzfpzLsrVW+rn6bcmAk85I0MCLwAfS8R0SEZSfV
hHZst4JXmDjR5hjRWjUX/WOAo+LXNnkTCjOJK4FgI8COr/FoZYQaFoiNZ3C69jg3
j1GyCcgspvCQSJpcsw2TnGVeb8SG/Q9pub3PN0TnQl4JWxbW9sYsmcjjWUdXa6Af
MsSSqk8kr/MxLU1azO2r/OzJ5loIKHeAL8QI0uwncvwNV5UFbnjWaasdplPp7oqv
837eJVhho4zjsTFShmLYSzrhvF6It1DnvCknUO/0wkQv+EOiKMiPspO00Dg8VlhX
kvGQe1JhT3hBKaCubss5vTu5HBNl5nwMmvdPa/hrbitu0h/zBQdJ1EZZRTxUi/GP
v2QghrqjXfCoTwGb6X+TXePuTXBXNCP19zTF8+O2t3kyALnG4GOLowGb9F55lbBI
PPulE//I+yk3GgkqabWrJk0Vqd+lxynw/BX5m2AomXfY0HkjbgCpTbi/SnlP8v20
Y6nntbMS6yuBwFX5sNKcSHr6RUXZqx1fd8RYb2SyjN7VQ1yCU7h+HcLqMVJIylB5
fqE8+iIwoJEqLtYmfSc8wuAt6zIACDcmynh8koICfLJ8GjB7OkgHGK96niEXY2Wi
f/IgPrAj1sZs8GE90MBeM35evN6jK8pt+5zPhgc3LPVdaOjz0Fc/RU+kUaQnNlnr
O3TTEiKFlPYVx+0qZtNIbF+Qzm160lAbuD759bUe2wPgVrK4/FpuQNMBo36w/ZCX
0MBiCEkXTB1LmkPAXin2II+oryGj16O76nw9UR7TriIt9lYo5R73RU100MQSWOMO
UFrZoRTeKbFf6rk+S0+gbhDV1eqZpQgfy5rVqalfcIrMZ5pZ694XbuzYkXsbbOyV
sY/3O+uhssHmX/Fg05ScspT5ArHrJYpLe4np1+IMwyNt5iSlrHSy6ZvRq7YjjtGZ
f5idYoza5wZP/f4bvr8cwf6H7kQBr1Q2lYsZvCJnUdkZ7JSe8hIR3X8lM1hLwGiA
fNbxY8hT1Mpqagb8ODvAcAu3PGdI2xSX2ZeNLtY3iB6eVCDv/AlDAAdcUTDzZOgP
VKmh7FFE2rhPhDpZ1IxZPwaDmV17/WvWRaxQbquTJPpRIUgCQsEOs2sbAbwPwD8V
Gobj1XcFWPLLOHdQ1VxOjs0DOae9ZcwCDswnHIykMRExT970kdf5ycHr0mmi/Tuh
AoLSgZZpK0ViGngguuX9GYHCuIDN5fE8Jpy/fuP/khTmbMjoPP0Kl9icew80Nbug
JubMlU1zdkwayALHpW2EAKfNy2De272/Agt0+ZHBjEz/qBgHGOZC3mC/ZJQXR02B
zx0k0Bvi46FgsLwxnr75F7aZ/liaeTOjCzXSmiur3M7hwiy2/mV7yrZym1GBawx5
IS2nq5Ht11Vd7bMTk4sDWiki6NiP9KKsEWLMDmpvRCxLThT1g1w0soFB6go70RjO
/XQi1zCTh/Qa24nqU9wOKQUsJmGS6zSwBrCNfe1j+jFHxYI6eljoC1eRNspcxXAT
PctQINW6fjLkeY4oUWfvDB6SEzqxKAgUXjcnOm8JLmKva6FwzkLAr1xlwZ2/O9Go
DGb52gtuN7DxJLDpIzKyC0gznvYej2IyKStAYizGZ/cAHTT3ypkcChuyBm/p5Oer
24kva07O5wEfgfa21eUw/yQDgNrA2KV3ezpJXnW8SYKthOrntOaNJHWIoS2Ej8De
nT4BDN8EtjsQ5458DP5Far2wEx5LYo3lGU3zNsSkZp8JY5CetJLLFquZuJoPk8/B
bX6YafgFigYStMRvUL4aHzQlQoVKBb42MdmQSHLnEr6fhJ6oTdniHwZqwcxpVM5U
DKS+T2v/fS3hvguzVGipDYkJsZNF3cueba5d4H6jyIS9UfKghJhaGZpPBenMikJZ
P6W7Z7/3wcYTDl3QLkqwaRfbmRuJpIi9EjYNIMaR/aCuSZVxiKya9PkrK71RPm2n
chpkwWu3pF24KzMJ4sUGUlcALeBv6Xmdm2gakn1eTL4=
`protect END_PROTECTED
