`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gt/DzFbeR4d/zfeCb9WFuTxHuNLOZjXyelkR/USN615mSVLxNUX6zo/DGl/EL/MI
UpS1PtZMK61uSYPI4VWZ8MaDxoHi2Fk/NIU0Ah+5p8S8m2UQKwhdU0R/BaJAA0dl
pNkmOW5ysH0/lgG/gaSXPJwQXmLg0cmfaGfUWKzezSyh6kMvEEjoui5U7zepcDW/
5baKe3JlpfwWfUZUi5m/IzI+zOxbs9Imza3rqwmKp98Zc2ynXxYtgbraXDDDxrla
7Zt/BaQqKqErcNjwJI4IzwNhHWlSJIhaW4EKjHunTFxaUDmriDl7gUK1t/LjXmIb
XU1mS7wDb948Zejpww8pceL5cUkj85/cJix00eXcKLPWx7EXEPe2CbYz9akIBgft
5bZMvBk0nxQOM3VfljR+ceSlqcsMFu1h+rTIn81APP9GmCkYJ1iZAukbDhZx481i
PwQayh21K7VAJT0MQVog0r9xpNzHS0syZ2ZVmtwWzHveYV/pMets4+VjFFXSxMzG
E/D9toVf+4nMRVcgCPTqzYuFuehSJHlA7136GWT2ODBX3EQV2ppMREo8E2o+R78n
Gn0sjLgnrqA3NC5ouATkjTVaDBlYKKI+z4E6MC6rlziKeX1V+ro+F9gqm7OXLmq+
FGD+mbPNR/6ueIs5+eoA1hBg5/2132j+4auAo7EUoimfmNmEp3c3VqBhITXXUeFj
MX5/Ss+/CBC8X3+DX1w2W6omYR7k4RtfJA6lUlSkNv6YHnW1R0G5jOnhpHhjGVxp
i9OFjaPCXE96k961UPVi8/qz2sCfBXtwYt+YUUBU4XTxJWBxaOfzKyOHQqPJs+XY
VWc2evDfuPKsgydpfDVdkMfpu7krcAY+tRfAe4fc+qQVtuneJWOKt3y9ot1zTkut
Ig7vRzkU+B5CpdOXlzsLYtj6xGCl9XLrMG4W+Amc2Cytfm8/YPiKADd37YlqUvpt
OexfpjjCKa3yrFmjr3Xaue5hJuo/5XlfFKHuoDSvUCsVQ5sU5NGWmbeDKtoNotUD
daV889Yl1jeaQoEEEalxgUcE+exHRW0T2XQ7UMOeLlJ7/2zMGEoe2G04FU29rqbv
+JhjYjDArDha5s0QPplhtiM59Kp0mR6QsIzP3RzqkAv1lLyaQTgBC+gR+SI3Hs0k
eA6dcie98kY93EmUdSJkQ0gZ1e2Bf/6Da6mxOw+n93zBlcN8j/WP2VEJkem7DiMj
D9Fq5NIEYJukOPWHtiaHBfqfBER3xswFYqFUZfypgSSWp/5rMA9ZNiJcxnF3cJCn
bh2cb1GUsLnFWM+e5aN/olBtgVnpoGocn9eB4uQAnEtMWa51bv9/hhI6rAlmNSCK
+EpV2JN4c2eS0JJqPi464cJeEFr9jsOe6hAKaGz3XbP1O8aQk1vWGk6clCMoUWpv
GLr98Nm4WGtXBoeBZbcTGd4/944qDXxrXPY6goxb21oHBdEzN0LymYvbOhpubyI1
xAxNK7NJRSda5ymSOVkXNovS2OD3yOZOehzBlrFK/awb/SiD7u+IzP6VX/OEUJ4J
MS9AARuskNDv3X6IG3t7CePsSKKKQbQip7/5Mx92xzBxlQsYqrUyr5FqN9gVptCA
cLGOf/pJJNVKYi1nX0sZZhBU/F3LGQ093O80GG6AEbBTnFy9IwPOBVUi9szw+L4y
vTcDQS13U73FtgsuFStOkkEnNSzBiyBn18ocRNAiehr93WSAiRHdZ0S+O4AjrTJO
be0fzA4mMtmi/ZmizuaxhJZWavG6/q2ffuw5yMT6VWJQzJ+hjtSAsDwqRbHzbgzl
mmrhV83T4JxDTd8dRBmJB6xe8OacHVROBNbyJPr7ms9SMinXEFqjKwGjNz2FkMqj
5et+ZWcwdG6zo6vaxiQ2ontnQWgsAGHbOYdFTt55vDGiL2+hgUCEKZe/zDcznsiK
NT8fuxbHa3V6ZWCxNJFaJlEFsdWyAbA1vY11XUo9ElAgVA1pcPBbMNkxaM6elL6j
GS80CptkxNwmSC/OWRDBLx8e3oNBrdeAOMlOvfxCVfo=
`protect END_PROTECTED
