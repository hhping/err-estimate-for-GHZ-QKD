`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/uBiJJYHCqpUHf0d53gHOVQAHASawisq7ATnYa7WkbvXMSklWkSECMp8STKpNxRU
IvoJx2pemn+HQEiXIGyhM0F2dPWutJuNzqVTd7S+gOuGkXsF9EJFpQZb0BHXdbd0
PCq5TgxL0Gir8ZDNIrMc1z6YvMhSpFLPbhfcuC1P+B1BfrJhcDxXcueNVGONau/v
apCOa2B9Oi0/GuHbrgqNdBR+cS7355O+5xDTcwGqLy8gIMAPlPk93SAptuPkm6BA
wfoZb9WX1UpO6+z/hO/rY77io1RLGzfAaFjm2XeKbW4GfoPLP/4Xl8XY/SxhAVz8
D1AqnVxnV/IijRSRIYsRa/ujL4yABK4HzIFWrWylzSKEd+lboj/IOye09UVbG/Sy
Py6bSG0SXulLkcUN4YtsBYR3g17MdjfwyAETtHueIC3AhahOS9cFWnk87IZAqsiY
nC7C4/O9iOcPFrDuQte2dyKXJgVzpaOhTgjqU+QjEZXsvQBFQUsjKgu1ExCuG0ew
C37DyYHLkk8qgS1XA0grNTTTxxdB5CUNNr4difWg239d9KCOrg2GehfWV4SqaKoY
cYwdE0BXK7xXSocwXJ+VE++y6MPL+9Cqrc95D7cUmFitdyctogTtQZyCHLjMhco1
SN36+kiSX7xIF5ijF5ZvShWlWhaFlrj3v4MHwHifVzwHL3+MoSu0QapWHYIaiyGf
6nkHLZaW0Mu0Cu+g8ImnoJSzvgSLvERtE/fBSKocDdznOH9Fj8kJSuMz0CQ1/9Rp
nG/9XF2eESjHdICCmb7rJhHL0j/7qURC6i74r1q/arQOigpssoIpFpMDiwWYRP8y
iKL6w/jwNZbaRYgnlKJ6+dZ0QZMKq1BvjEC3EGuhvCJTexJqzlN0lI3+MjrmA0go
MZ/pax7YPo7JvIuzeivUmixEJH22suOjxwTrWFywUpuYKR3dGdRNqFUBWP5TLPXD
7E828Dy0YBgT9fT4eHQflasGCu3r95QAykxRESFzRgWEnMXmi3q9dnLy1KZYfx4W
PP2ekELbUU/y/8Y3BDMXK52kGeTRrXV6pUyUFIPtKMA0tM3k00LZYww3dRpErBC1
LDzu1wz0E/YE04ALaVCsQZH6uMjtYk5ZKKdseNWkzgww5qJquWTjmXKEiS5ZD+TK
j+SXit676QcQCp6k73xudczMUXFL6x1kZ1CDIL6vO+Pp1QK9QvMLLY7BLPmGzY9T
gvyY8hFFMQTKJZPEEF/tX3lq3IKOoLgSIzI/5YdTJkNx/bot6vi97Lt9KVPutRDM
L2nRSXXM4CMd0uTMyBwe7aq4Z1LEewlj2F/z/gDtIJD26jYNGgYoWifgq8ZKfjnR
kZntaR7JXtzpXLRwgzzBg9EQlJopdWVcyfQos475MR6ejZbeIRnJVGHvnnJh8DYl
2o57uRihOZCWGUsCssL+ili2rt1e7bTbYpfHk7lQx/EcRLOi3YkYFo2LtE0Wk/cR
u9+XEvkDt3qVUA/WYwSP4UOEhMVPGCKvATxdXHP5R2anQFwe5AHmfkNf6MBO7cWl
AK9B6ESTBKZVHSPwOAOfi2AEIkLakMb5shfVS9bnqoqPlIa9phHmPytJr9RjEFIT
tZsXt9mls1g7FpHsh8yoe68stFRm+6RidNoj0bTNnJoSizA+20ZhZmW+3s7zQNOd
u+JYstvCLzDFm0FeDGVPpF7+mJl4loTF6OdEZarKBX6Ll0rE/ejei74rZ/MCyeO9
p79XXv6fo+bljxGWr+7JIhadrznw8vHfwhXkcfD6ZHyDKDpJ6MQAar/isG6SwHjy
koRZEbxAQgO+CETyEcWFYF0kEDb7v6KyVzjNed8ULTlj62H4JsyWpvkhlw+On701
QcrBndMfwmAohEIvZhYUAT02DBBvtsVhb1VKJjIF1NDBZlRbmzjGcTvmGouZ0DtS
oLU8YcuZnd0IkjryOVS7JC9WvCsTpNXsn/0U9rcvnjrE+yGCrQsNEa+GORvMd4za
m2VnrtNMI9t6nSYa2XksWsoqSHEYX7UACKV7N0FIUJRwMD5Vv2x7DuTrVS58J2M7
rq1WTj/Duta97qZ99IzAGOUQfOHxz/KN8fP2mr9ysDvg36HSR/N3Xs04EoX3k0V4
05Iw2YAiYZXPaamNYQ11q58YHa3v9P4l8r/Hrwp5sm5k6nPEhUkLrz3vpCoIuBbV
HHryduNI/Ef1Fnzk1YpQbeH2ruEOr3nSQQz6+PqkdenBX2BkUcu7NwU0mpM2Pt82
WUdSiS5xCBlHaack+vKHAJjr77ltU9F4tvoTViHIFKWYuLxU+CH7nLo1kxwLEdbP
GZfIidb/Oa0wTfUMFGK7oM2jwft9MROHlkBxJ30jnroq3hqMi2AP347e72tiLFB8
o9ZS9aZG3jddmHWttg24fqEtpSYsTDsV8BbXqlR/LzA=
`protect END_PROTECTED
