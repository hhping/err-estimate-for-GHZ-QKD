`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
og8oSUxcJBJfRJwyMhu+XtBG0MYe+zRbQtBgJSqNEwgKgcEUVNkf0UMghndUWH5T
dn2/ihRjItP2NbkpI2akpBSbE9fThOZQdJwnW8QBbX8LYbX0Zj9zDYKV0V0V34gz
1J5fYWuGuszAGNDRKfhFDDPKxAITBL8DljI0qBP4INaM1Lh8/CfENOSD61rIoqU7
hnI00lmu2x/f/JCNU7FF2tGcQOgUikzS+U6uF2zWHqWlVpoG58LNyMOQAVtxEJJX
T3C6AF38jUUcg7vpm4sQQ1Jyi3kUQLcTJyN+/VuDggG+U6FQVS2MtGpEe0dX2Noy
4Lr9fvVEUyxpaaVOqNJywrw5YkGDDT0jpQASzeJH7w1SnUKPGlEAducUgJ8Kg0ft
I3kGzBQ5txAJ+enM1gYULg==
`protect END_PROTECTED
