`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DeFHRteXCGu5N4o8TjZHCahwD5sYh2G8Mz5Tq1NoJJzRd2ErBjk50lfvq3C2daZX
MeknMSjPodi39gIO/JZ9/ru0CpKRxNcOAae3Hn8gqmFGaqsujW5yiaP7l9GXCNFQ
XZXGz0CwceJN76z+rmrR1gFnhv5TON5qPSRldZVrds42QLOkI6ukxzVKGjlJKwet
2DLZnFVeRzVryozQmyTNKWEQIYgPv3Agb67UcENjRGxV590jZhruOiIkCJwH8dWg
SFRUFkiZTapvJVYrL5uxU05osdmQjKsG1LLyR8z3O+8KO1qJBbVdJVfhboj1zPWv
iSxffLDEGj5JARv1UTJPm4Lp9L2SZqbY0B3jkqI9/BlePVEvfQb13dLK5lZWu/y+
ceC7StAXzGC0jF7hQRbtlJ5exMIYvzEvoTHio3+j/gLgO+K/epcVu0z7CIqBf+Zr
wNAnEDfNvpxJ4MM7m2s8afr8lhQfWy9UoX2ndS5W6Xwjp9kPL4DL+dwqGmK+sRkM
SuC+D2GXQ+zbjUPm/KRX+z7RXsiqgbyiQHF3wrjG7CD5CgWrQ+Ty4A7L3nuytoSF
w6qomHN9K2a5NY/sgI1VAp6vngDU04Jy8yxyEy5Aamsdg2JamCQb2ZIutGRTZH+g
Ap6aTYBtSKZ2JtieKU/z8BymQsXnL/2CKH+Sh0XE8euMvn7DhaN3PDcDO8m25ut9
elhRyvW0HgOOlHbYRPlw5ZpuY2PejFuHpPq+DYaD+3cQi9RL4Xi9neDfibVuIFDz
NjZmJY4xuCQ6TMsh4zUDBUtq2pgKFQ0zvrYwq7HaaoTGFxKO+9wBxS+bJNJFliKa
Hxd+RBEbDdKK69CswoOywT3uWhH7GdtCxe3vkpjUpw0ScS0Jppp6QOwRVx4z2p96
eI3pknupRxZtGsT8xhcM3Btycy7wnKxdpqXySiXP98uBAxZUGeWUzlj9gwZYPSzo
y70gMRe0ry4lrdf42Ivj4e+SmX7F9HUX3A4g/wiF11fVUKyt8VwAQ7phXU4Jlb7c
hR/QCB3cpzauJ1mdTzRCmeS82G81AAYbVfcSUl4P42DDzVi9/EQ7qYhw9GUIL2+S
4yFEDLqLH0yPnoNGTnm3+NBDdJZpedL05WXMoSIRkgoVAZAf3UMZ+t1pWoX1CCkg
AG1VkWRcaMaXCgri9ot0cFEwB4owVUOHFR3tQmHaD/0=
`protect END_PROTECTED
