`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0aguwSN6sd94JRQzmiXzXoDbmv4r04jrh2LDUAX9I8oczctlly0m3EVcf97rOQef
uL2ioCv1saSLbgnf5T3NM7Z3Q19ue4Mz+iGlEayspSyBkjVhMIgzV17u1HzDknl8
uwwGXN2obWILrzcd4Td/W5x9ECcKhDCat5OofM7BtLCJbGK4SpB2LlAn2GQXEgSy
k+9aJx0F5xHFNfx16Bd7z8PE7C6HDIRrgK9Ames3yhHQh4bEDfj3XPnWrs7j3Z4s
tB1im04/3B/exUgatKG6I5eH0cwQW7kVhkWNLxIJaVtLQCq/EtBb2i29u56NRxNO
lvfv4bdrMhvKz1WNvyQExLu139V1MioUCP4qIyTOu0EGmCsHt4dNvlRZJtfjSqME
O4fcc0k+hYB93timh+xCFy4qex9eIKNOfFqceuX8dn+1zmF00Em1pSLNSn6Z4nuu
Zs/Coq1OdfaWnfFRhu+DAN9VcvLDo2ht05fUVgUGVdj9r0J2oB+B+4Es+Ts6N8j+
rtN09i4/NiKoghHWmweSdx944+jCn0UoAQfUrdfyXWhFY+2MoZ54eCElwMxE/caN
N2JeHeYhY17oRYdbF97oAWlV+ON2V5zK7lxgU4kF7Wu/LUhc608Jd5wsplIp0cCI
N9NLgcTCaIqhLeavfU8mMMH1x7CP6mVQRGGrJFuf6bUcgL7c/29IAI0HTDfrzrJn
`protect END_PROTECTED
