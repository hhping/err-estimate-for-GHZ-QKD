`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rMywG5F/bJ7wDCDPov5rtljIFPRLkKpIFFWp4BfnLXzPi4vgQSAPAQCZEwcV8NTY
3fmGh+qk5lFDNzvOD/gfULC7UKPwb2nQwwXZIJn49YaavSoDahIteisgqwd7v1ZJ
C1uhJHHvFYjRej+fKhnw0xvdgvTf2/r3TbvIFnwmb89kmPt/DeEkBvnBySqImDaT
PjhCzNzkB2FrcCacMocJ0OhfckupJmvabPauOwoI+KXOGa6T6br6xxoW1paY07TF
LXuHzE6NlRFueaJ+BaXac1Kmu8SpN9hEnSJIchg7uobAd/DkWNna/09K+1WqwdaW
4RPmbegl0AkQJvmcCtvOn2x7zqKPM79wHKmS+ZALfNJiPceXbQNDLRZDpAjuISi+
EZEPfnKP5Yi8WIcYaGqyy+iT9fueChVOvAef2BGq/UKchm/15L0U7x+oSgo+/AM+
FqSKpdtBvp+s/rbQGr4XXZpUmvjuWwPWbWTJi6kQo2a8sybkDZ8CIeI0uslFAu4T
iVhfiZrZN8dfwUCEtJxw4cz3Px+ZzeLvKLbI0CVLtEydjE6TG+Xsu4+0gfhwXxFe
0NszD/imyGYi25d9OT9aMMvLyMn4wJA7QFzdXTT9Az1X9mJYIYY6kX80wIuoI/Dv
/9D9b66Ga2+qpvJ33XQd4Y9XiaC21hcaFwFJUsmUcR5d/avlngQeopigPJwPA0ip
CfZ+BqTdqZu7t8/EDSYoXvrJo0duhF/Q9nu43PjXUV4TWtHAWCoK/F2rD2lWLVJd
/dzP5o8+lctnSu2oeQJaR6rPCqhdR3ekQzlpQeiPKsH4QIqQvVc0lGym6F0WfukO
E5hKzww3pR69c1mVrxcW9i47mwhPMBDVpTrMowwjFtDycwu9pBFZ9+ug7ttuWlvn
Bgzl1wtEq8gdf+7nYmGz8474hhV069KSYrW4Un5OKUUyJQpnDkI1jBY7v8lmMRT/
yp+FpWJRI2OrX6zxqd6RHYhVCD3Jiq8COrhZx2GeJBgtu3CrG78o+PwyuX5PuKMJ
ys+m47eJlkKAF1Pll7CGVm1enTs3/IgStAdw90b99xJP+DQHvqVMUkaXqlXvoJIm
LJ3gOaRB8KU1yAS7NBNuGMMEoZ+Qc6YUTujx6GWOJ+Na2SHy6o6fzBm4As5DeOjW
LIB8vsFT2p/oy914TPp7MvIFrTjN8aAH/5BvHIAycwayfgRHIg1R/9ek364bba+5
JQPUkkbCNtFZ33YqepR78OLmxDQ71d6ZxbqL/uOWeA84ZsKGAjPqsQ2RCp2C3Dyw
r6qKO1HwWpiBVLO+KsRduGkmHEQqboW07ajR6o4saGnWfapJP/7rxKoWa01yIKsq
2kYBZNv+ZtLKumbQVkRN/pJ/sUHO9ZO2i/c54lFhYeyI/+1dsiylJ94QVsGEnjxh
ZSTe/hkUGG5z97oLqJSU5QCDLJouc8DBohmtPIR6I0rirqwALOzUgsZjEX9JxpqM
`protect END_PROTECTED
