`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kXBWRmADKT+rTAdpKGZ8ijb2JpfCwJh7I6iZCgMN7ByP3NRW/qcSWl1nr9yhBNWX
J8oNVRz0BoRK78W6rGOB+cs1j/V3Vm8fPvolqNx9Ir7MJ84YY0oOFbYwjdN3vsS2
aM/q3SbyPzbSEqqsqV99up5d1Wnuf19WCKR0ddf+yvpUEScK9wuMn39M075aQWV+
o0n0Su70zRa10LarOYaF4S4aSWjW83ABwfTwi62kQR9OpT5d1g2KcwMieNwh4yRx
0YDMjks5A356gnoLliBtJWFWnUSgd4iQXNBft59lcvdy9a4ZT2i5Wmi95gnRx0/O
Vhb2Un7IrH0Kl9WnXT2gHrbUEKBBo5cRwQCbaqCeIgd533Wrq2CRH0lEKb5+/DyG
V7OQnCC+oVBMh3a1GScMLEmEFXyK+YMqt8hwWD7WaUy6dPjAx+WRVIxJlA9CpGnJ
YndQ6jnH9DmbQYNTF1v9BV6fWA34AcDWfSZCm4MRoOxjiytBvtiY+UmJ/ni2ZaYJ
qf6tb3SmryTZh6QazIqEM0Yip8z6EzpLevwuy20gnHrgg4lGrQ0mf3ddQhIFn1t8
ySsnRzNZv6YT9iPhRec9u0+d/3+Ieiwb+G2PScZ49MCbXnlot/2yM9/2cbUSA/iJ
lc0MGeVEv7l8VBTtE4ySjXdE3gaXYiMvkph5aUpcOr/HBMhFBZfbcuaOnBbMQktr
FgytgzZX6HAXVT5q5q3gb3M9zu/NA6Rw/d9pHqXxJlPOXUynxvEbJny80LJINfo3
qUmAGe/mciDS7WzoWGQJIMT3QRMBGhj/A/DQSGDXhyzHxxAULrximJ5y2Shd47Hz
5mbRwLxPTme4bnaFHT6rYv1kCNnaV4TZEtTla1EUeb0GTNxU7uFTUzFX/uzwwwze
2OnXkVq158TSMYFGIdmVT50DgAvarRMJWn8066WuAYu+EdrwKIKJBtzkFm96Exm/
bst3C61VOuab7YlHiHMYPXbU6NsGFYmRqggtTyhYRNGHQ0CY+05IKlw88p2IYXOY
9HKD24Nm7EoT1kF4RWegRvLTER+yra5pLKFhbbkvvXMiePfFLJXd1scOjsu0vFM/
4sWalamAnt4w5/ncBuRkXb7sv5mrREMnLCEPTbhl1fQlT7udAdf0BOYmVgmlmXKq
6Je/m1BqKKjit376sIDtWUWZRYMDLBHyrnhiMGx2UGi7tt/Sgd2eV8S+0WfVdpLW
lVIcoaemMfreqNpbgKWY/H4IYe8pzIX0doEqf7uqjm1OmmxFRrYGCAdl3Y5tDkHY
H7W+ZGEUS0ImlvjBtfC6PRAPISHr0bCgxP4hQaSoPx/VzG/ZWFRb+TawYIkeWoRJ
C20WminQNylkJ+vwPtVTxqNV7EimsqpfGIMlk+yStxzFds8ZBkq94nqCU/QW3L2Y
lMa+Jz+w+KO2eHSfjo9NsQYFb9vOKzrnHwI8/r1HaKo3enITxxNVwhuY5fwVU5Xp
+MxY/SzfRRICZzpskkcoBo96FraBEGL4lvutuF/Y2OxbajZWhp+LQQ5o4dTzLW7W
MWK3h1BUZpDtx0yyIGgKatG0Ry5fLiHwMijaIN0JAocp+Fa8Nzr5mmEX9nwCI3tw
mJAswiJ7fIShw02GAbTCp3Jg2mHOZAl84gcIt9qOxTLPOC96OOhRxkFTlR7p8EFR
GPNu8tWhIX4glvz3wEkbiLArjQPSZLJP7vNhSaTlQX8xMvepYvR0Zl860hb6WdDq
kYit0VzrX14V4oPQVW2cTGfjLWTscVmDXk6WBG5RdTEg8EgiqsoQjCbF4zN3t2wq
jFkF02z4ZNgvv44YqYXPaMa8cd+B9qLAZbdIRmopCRuU+eaoWReaOM/OfQ6LbvZo
HE04JoZhEUXYmQ6dYvF6CnourXyYHgUWd8yZNPpwvwCN42LwKglKpFCobhBj0Iiq
uWc0zYjjwEfrGwA0GtsvWej9s0bsdxFG64odlshJvs+FVbcsoK3PwuNgms3yEwL3
HQr2qQFCY2ZZW8daW7ohgVxoe8hTpVbV5qzBNWuF/8KDjqtvh/LNbA8n+uBpElQL
PpiL6hEyCuZPehF41b2wXso1onqMQMpPcX1dyG/5SmSY+lPlBluydtwSVJJH5e1w
P2meMh8r2N8i5F/m9d/WLHsvD1NhJE3s/TFwNMY2w+KHVha2v3iYWRntr0lVoj+u
6/mmM+mkNWMIm/hQjNgU3XnL9jWNbTVs4Tvp/1Ss4iEdVYbiWREDYG2QxEguoTkp
fP5nN8HOjbKR/KrIxSTDAZ4edwl69kzHjdAVX8BaK2KaIN6+xRl39003c1K263dx
f+1o9qoROgLk+skBV3ES3bYiUOVQv6YPiTgUG3/uv6wY3Q7diYQgzmwXBnRj2G6j
UXnSIafeLSDseEqkXbF/AApA5CvyVOYaA2o23ylcvawpoEqRl60QJWwn4gFpYU1C
Uh3EPvY5bRn70Axc3ytlRu/0i2wFXIDVJVMDqzY+R0ntjOSO04UHrArTdIrdOah4
ulrPW8LIH5klsO0AkJEYcmglC2qdv7KymHcbabCWSU3wuEGoer0wIn6rhurPmJLq
Ubwf8Eg8fPgBfN3MyhfAK6+D4W/2GkMOCBbiIGyfrF36R/6spUYub56jJLAFjs6M
jcUMgHwbOMv35hvRDghTOgSLFHLREIG1rZSpgSgr4Oao3IiEzIr7XIRPLwXtiYpu
pc1QrAgWdCBgzSoS40SZ5zpxHV4piAUYKnz9eeXOQJcWpv1h0HlxjGwbaBvcATPH
Gf9H0TBTHWIYM/5TaoQQQcWRTqdSxCBjFExvxXMevluUbMC8udZBD+Ar5U6SRgmv
spuFz1yxaABuFqbFYuLznG05bBG8IqVcQNDur62L8OBXqNfKcuINzYzX3w8STnJ0
5m0pMja38WQTgVABz33/HvRPwqN+aSvi91xj6iBmGmxKXXzBrXqdyvsHRq4dN6+C
Nx6IL4uNHlaQ8hj8Mo6yC8pxESa40DAyh/Jac/Rm4el2EG7upb3soXiDrRVzoCcv
hgXejGm2fLInZnCioTNHn+6LkVka2QLcgw4Y5vtikQ5lY+4c9H0Cl8ylRj3+yhHp
rCTnhnUN4xkDKUjeK5Gz8NE56ZgNeP0yK6UvmvjX+e8ZoV84PU7vj3IvbgEXuCoJ
81kccIM9mOXgzYYahpHe7fbYZt2Xv3sweXQSqhvt6avfozlgXFmlXjxAkDAK8kTV
GPlsuHXm4vNJDJj3FAtfuwpnWOKmUsQBZAzq4Iz6MFa3luGqz7D5BIkJgHvCntnd
fPOObWCvkKURLMUuDwfYDn1Ks0bbQmIZgljtJcyD7uhKRG9IZvOKR7TaiaTAL8PG
DOSx7nsFR1u1jpSjhFbu8AOCqAWCimF3Gy5C00JQ1RCSzC2hrI/eoYhi2hWcWllM
LkfdkFvu5+y/oH7CxfQgr8sH2uO1WYIXst9u94lde0+4GUuNrGBdGRMbDEMRv6/h
k6UWxmj7PQ7c0YKiJ8uSKsnD3yBLzAf6EqD7h5hQu++K9g/buybaTo3qfHtp0prF
MWn3nM4oIZrr39Egg+XOkeZcjugvTi5AM/tj2cTJy68mcYZg2fLwnm/zFPg03XTe
hQm30efV520CzsllWN+4xCkzcEujfev89FH957CX1QWFT8xORcldxWdMG0hgg1mp
JrEH/7YrqM41iAdMlkvpmiIkU0ESKU+feuF35JnEKjU0mRwKmzAqWxSrowZZKUGO
Cj2kf3XwoKrhtk1Pt2YHoiOwvIrs2xdl4+s9kIlbEYc25Kuz+VlYPbKJoXQdkUaM
YkIXw+1yUnMcI7zWdawtFQIbU1vMa63dUk1rcnfHH1PEYYjz0XxB2dNRwr5sqFJh
KmGKkqBYprswJ60GU+TCImJEkutmHZ8glsIGItXiPVrxL6wiNzt1FR/DyrDO4810
bhTWhbsrxOljsAWqeF+QA4TITAULG29r+Ppr6q5D1EUue3pi+6M/KvFxz5s7ORdz
P8LIHQjt3/YoFSCNm2UiYavU6o6GH33RLEE4W87c613C9qP01SsrBUBNSi4mEnwu
2hNYzUDEPPUgdEzy9tkwGPTBaAuKWqDp7toVXtbU0cdffCjIo/TzcnId6k+nPaOT
J9MTnKgxnhKdi/4NUNFzC9SwYauo0cu38XppX9EnIfLAP5ZA0BocLVyTd2bS91M8
as5lb+qDHB1JPi8Lf1LQJczbefjOgV8vObA65wP5BUBYJwWawTvwxwbb3WtQGFjv
33YOkYRcrxXF2+x23jZg23CQ3nP2SZx/XXvg4jS/1hMvT0n6Vyg5h5nrjr0tBqEM
5ISm/5Lybkw1qFr3/l4SrG5tGykQBs6bJ63XZCkzzp8dlomH7K2G1eyxK9YdWV7c
YEPavnOdcy4uaWh8F7utjD/sSMXoBe/w/N9jtTNbo/7B2zc4P+ogxRz2uW12nDCP
4ITYUAXmHtMhhyt7daOS3dUj/UcyjWhx+rVh9xdu+rMKv3I9O0dN2OCnHCLUIpE+
A23XsoHbfwoDqyaXM8uwSybgFWIFuKVBGRBMqZyo6b8iNCNGl92zzbhL7KFG2ChE
q+dtRGtRxDqntZb6O6ZuzNausqYWc/DVi7D82uk8ZZXU1SqXTDc0maGtkYwamOeB
x3PAoUAh+LMITVMlpWmH+enM1vdjApZyDOjnud/3zm8YQWnGrMPIj/jGcrG2/Q+f
1gh3CJiDIl+2wuLIncvbOuxKJ43mB/ZLSBFCD+EBVBUr/sGDKAtWtNqlZ5D40Z42
iQ05xK9sUy4wCzScsJEylb217TZhOKQgVdsq5+no2Lyzfq+pV3ublP8X0ssT3uO5
dKzIxjR4gYEF0o2Vr4P/06203I9KBnOSQO6cTAB1MYy0BdnBxUl0h/yaT3SuGB5O
hhDSt+RZIvbTnzH+rvYHxBvfL+LpiMxGY0uBf/ATi/qpd9pKUEpDwJm7izr9AVmF
gcvZz9NqclqqiXkhD4kjUbxpoIQRCoxn3qffQgmrD4RCPUw+75mflKuaEqAI4OAI
73lAokbgDoe1qqmvTKfnzE2icSyY4+2SpwPEKKem31d0RhN7kAep4+8wC5d3XI1u
fhwPTFS6OGywulTaF/9Rqe49/6gG3wa3YX+dzfAkn0zhWFSdB32NTpzaMlbhc12p
6lC+TTBWo8UBqRKrfu8Cmh2DbIC7/o2zOqU1F5++ZWTLIZvlfBoGFP2eP7dCSk0S
YGCGQTVzCju/VFG9EAk5HsNhn8mU1b6hU6pPtYQ97NzL0cqfRoGEg87mYt0MXUbs
T0fnTEdlNWzxDCQsZVJVQHSevtdJHQJzoVH/cryhKBCS/e2O1LKt8hsat3C2ae7Y
PHKKgTwksx8SisL+h+29LOwccGCox0uiUDWOr1hgfHyAFD0mvSmK77LyUJC8NO3e
DCz0034eqJLUsHhTGaD4dfCaU+QJmSrkfZFq9WSXcsr4S6XXbRcrIH3S/4QE/MPt
C267Gw3YqZ8lqv3zYg/x2+g4FZhe+OCiCBhMDTiisGqXcNZucOyjrVLkKnWELCYV
ULqSnOmYqxzXjujEQ9mcE/QPyCWUJdOK8Peqo6Fyf1XSDuZ+Nakc7ZzoleUBwyUq
jAxSXts8+s9xnjX5i41o/7srXR6mY7jZ7Y+FtNNmrrx7B764Z7LpFTbZNYmzBpUt
L4rX8rxnvz31x9vEUmU/Vwx2HQIBWLWqkYMR4cS3JIKAor447bUGTc/gNe5VpyKn
2y/JOCEFB0L6pdvp3SNT7+SB9sgV9VklUwGb6z4DBoY5J6aUeCMyzK70SLlQ0mI7
x4Stc30oxfi6JzPUSNrkXsHDSKLqoTz7XDlT7TJsDhtbmLeHrYRdwWRnArJkbgr7
/JbWlZNt091KEl6wGZzWj9qqbEspn/TJ87tQ8KcFe2rKjTZN+rsz20grV2k2cBLj
Be1oQdqc/9xTZrhbhXkiNocIc4dvxoJ+LS1Xjl6SJ2xpS6HbCrOX6nBqMSO2uYVP
xVedXQi+h2Kbda0cfqasc8s6ZvtwDvyQeZ9q1TRahN8PjuCGfxV0c+dqtNi9Ftnx
GkN+DdJhi6w0UX7PvXQWsdEDEMgASFB6AljHMJxurHv7UJ97c3A56cTpCm0G6uiz
Amsb8wGdaC+M4aNXPxvN+JZS/cZAm8LqKqHjfcFSYL/o9vUBEz1SV9kR3pt32m2y
mEsVDa5DKw+ZC5U4Zk6bJCPtuSXQeC1WgwEhOJYIs9bY2vgoZgdY+U3I6vtTQF+V
3Cgt9fEuFSRqtA9/gcp/TCnD1wlpfZUWbpHnD6yCADOjQTFYKB4X+7XJeAON/8rk
FU9pZtq2pgBfDr+vOXqIYXDibvUo7kKO81Sf214AMVjfSZfwDyKBLYJr17mBH8tt
fPZnQBMkWwbl/c0H4SN96nFHFFEZrm+MRTwQAqIowhL1Q/otj/VT1yIVBTil9Jha
T87pl0ZzZFjBYBjT4bx2ENSsW2nhB2VLlWQtGQr5CI++7rxDt7Ojcp9LNnsvE0m/
uuRP+Gnc4NSCbn6sLup22n74IwDxLZwP8d91aFGe+L53SItCLVDThTRAY89bJKRy
uHcKFUCS/iEx0EvXe5AYgoTVPmZQgatoJhlyLDOiWG1/2GyZOHxS/TJzJlSouZBI
9nKXRv/K/4KitUY9cDThuvDifu3lhuYPeg9dnKly9PBXZniB9sJhwx7ZeVH95Wx7
nYAGdzdXerAzHG0JHr7a1xAn+P5TDfYk8c0wwMhiEWVQJBqdGS4+Ah8oRpYvLOGf
wU4h/mAWyGFOiwXnE/pB3p+u0S0R6Pre6I9OiLuTlN5T9lFkpKH+Y2ob2MdqxkSK
UObX9pX3BSsaljU+p0VMH1nah4t7rRS6GFNbCJe26AbuMYSJv05n53Ih7dQgxB77
yohn3QlOrXvuwkctU+RlvkNjS2dVhEmorHF+C9ZFeFBfDhhGvU6S3KLV/vhWCQ+h
nteqTgX/+hyUSD02WNJqglGzHRsU0hiv2kcA+EATF+HRcQGI7zQv3zecNip1x+Wk
l8B8PnFLy1+TrsbIJFcnfaQkEYyPfZnlNjxBn29WD3627jeILC2biA2+B3smuipw
cVTX3gBA7XXcOkrsbnm408HQspXJRd5pYVbutvfnFXcYZhPdd7s+kVuKvMw65TJh
SwdxGc75YEXIt726uaOVN5l0ALGpm9DkOBkDj9wh/QxNt2HqN4PfRs8BM4y7um4t
2knjW19JxjtaP7FOBpxCtOp/0nUqpxGlswzbkkyW6fp+AIXE8En6KVKQE+/+CQ7D
KwjoFTwwGA/ffCiTsjkHa0v1o7Ebm8bmRMaP4N9vckLme+St3QRZq27ynyAnlzKN
I9+EjvG3J8MoeEBdMunOkmFcHnvSdY0vHVh1cxd1aNoAmj4fGTM1LuOsSLq8pSbb
bX5Z2YxEjBLRi2wQoEfcYWr08lX1tgZWUBHWoIsixFgE4JpnZuzjpk0TdPrd01zN
YhWmeUFcCKEwshXC96O8MvGLrXetOl5zppu0zqBikr04bQe2DdrQDpdQ7qxt0HwC
uc5U/lQo5lGsLZvzwk+pEks3GrG+rPLoFAKc41nOt5BbM9CcXgYAuQ6XRj0rzIvE
ymi+gVuknh3OfWzefX5OE4gHsg1pfD8AhjyjzGtLD1ZQwYHBVBmuiG07sL9ASZyk
ub83Q09Cw2eXhWK0oaEYnqtivmX7nD1GYuXZv8gQLgxR/Fixz7LASe/7aO+p8i5h
FaDr0kndsuim7YwfzVbzx8AW/i1gNGYE1IYLrnWraO+MipJl7n9IbMX8aHCuYqla
fqkp9cLZDV2Z7Lj9NmjBtHbXIeCQkDGt34b4IYjw5TI46kjtWrragSwg399KwOBJ
4ZZQCeIJgPIqbQpWmxP19l3E0dI5+4cvm8uBNlyw5OfYMXAuKmFvFdMceQL6V+Qk
gwKZIkMRionUvyIzelMW/sYOtr1ktUtUl4mKv7HjFlPaGpmL+AIJxe6viTdM7j0t
xq0fRE0J1c5srKzbS9cmImk1+gYE6waG3QyGdN5699acjdCt49OTajrzhU9SAhlt
p/3dCB/XaWbZW8tcESj0wIBB4OeqcwIVxt1e8KwtGMc45V3rtvdg7XcbZxgC/o9s
ld0FnKT3w1ZNCiS3DeBhrB8wxp+iWv4Hwlfv5zrO+S3G9of1APD9RmF4cxYRlbEF
rWWbjmFhw8umHlcAonhWhFbIlmi6nA1g8JHI/UzogD5vC5xDerzFIRruAQHWrR76
NzH6YsTWJdxwbN5LsCjH45Z56tmEUczE9f+Dac06tSmRonNV/g+VE9RdbGe3loxc
ANkFAKXGyLgBVYs9UQq4rhe2Roj8S4LnENXfp5BFxVCgt33j18FZDQ6yckr4WRxa
lkh21IJAZDFizxrX2aFG3TveMMtym0uietT7U3O/W89wWslzhIeJCb7gfoH66ne9
wFKY+U3mapgOnaCksrim2Da/7P4w7FXvClhSnFoYhoeQV70kmsz1WnUuGeNrO67d
ApdT4Bamoa2+lf0mnu7Y2OL0IbS1Zj6cH7HY2mEpP22LtO13edaeT6EM8edEhQsQ
b53NKnK8BlQEJUzwgySjPNzqH73wZXkVrVJFIZdXIw2gynW1HAyMUcoOlcnLS+X+
elJ7YDC+/CEND7Dk954nSgKG+3JwCtWCIft9X8TtjWyZj+3TmhugTeGW/Y8Qt6s9
Srmln5qiiVwkxG0QszuN0gABmkGmvJ0/Ur3gPrkicltvpIKeGf3jAltPifK7rCX8
yaarf2fRmeYqWVJzFtfuaOFfC7ZIpTRu8Xf0z2hq1xhGlB1IgP6rrqMsVTTPVh/Z
qPLAWYtsEHRdMSRSrYiFXrOt7q9CRvw2iebtMu/fbQgxVRHYEdvWLLsvlkMokytw
m7G5y42YXChv9fYhsLmCWmfiVUBsFPeBvbR7D/6Yg8qdWGXVP08EOLoSQEYpTasc
3whejsesdYURqAaZw3qObQ85DtXgFq/qsi4q6+1iaNhR6MVNqJNKCWma+TrGPYtQ
+OdymqdJpLXeqhnk8vvat/MCO1YqPKMAtZE5FoiHj4U5ColZ7K1Y+8B2E757W8kl
0n4TeJu8egaeh2zW22fSumKmr646fcpJYN5q/bP1MAzw5llQRuyRgljuVZPADiKZ
EOHUDrD0tnMP7htyEZR7dA5PuevVZeAhF/+i/EiqkIpjINbGcHpXLmWDGVSAYHf7
/k/EHB6bjAy6JY1nRfhbdNHVkCeCi/pD/7B7lGt7LH9Z+tpZEDmye3GziQEU++QY
GhcaDYPMVFTn/08gd0tciPvTCRTghCfcO4ef+jIUBksJ7xtDnvn7Nkv53BXDiq2l
DPHqCCuXP58MzQg78eWgw6kliWDPx8clb582wP7bYTf6AOr4zgVSHWqhhxRg/E1I
ArqdhB6afInmp6jbdLahihkD7xGrmW/2SEWzDJ68pLUMHHhp2ASTzsliitz6O1Fa
P5PepWLW4HR8wXEcl8285SGwV0UqsJV1MgN1UC56Kpp2CkT8jtGlYm69H8X5UovS
tfUVY5FpvzNOqw/VarWhjJY2CP/lr2a4zo0DE3pVHbev8LEncByR9YxZhBjjDFyK
Qxi+1Hx3Sgcxi68kS2EYRkwEWb+CjQN/KXkizsAO6YGsk0VBQWnwrto9ol69yoTt
PNLOl80FaxduH7ejdwUve861RvDNWmREXtVOB5NrLaDiN/0cubLupSHVmRftrzPy
S6NDHndJkO937qwpvd1amVfIRWNdRhErgh6aSJ5fospAztQSR/qoBJdunPt4wm1E
+F7zvHxE+nGde24HBYPjr60aumJF/0/Q+vWwxUbd+gUmljxf3AsXTQ+JMTZeo6V9
b6ZdcdG7VtUJccXO5YtzfH05rCz2Tv7+QMwNFc7dTVS5M7N7yh41iEqLmS2jCWIl
1qyDo245ZJS0klGP/tlFp+q6LnNLOxeoau7NGnyKjTU+jMhm6XKNlbEIMpPUyGHd
8R7p3d6kDLfa3STlQyPNwS/kDqMSdZPe9fJ7gfxEnzG0zzQr2guR24+JkOgKI3iM
6rb1xYgP4K0JWOZoR+dDYgeSI/8r9BD4y5G1qkzjYQf8U6WMbaGaJ3+yVlIncvZd
ibhiZKxCNFcHSMndvyc7O5KP48D1qPeEj/awaNR4b2qF3Y205TrALlPT+F5Ey7Rs
17qfWqX1hf2kWGb033wGc+6ZaM/9JiOBSN/D7JJTcB7vqXRrPIgxMFxyFhZBr+om
L9c4pNuilZ7nMR3Apeex5CdJuDY5Oh7oKkB3sXosV/mA6oLJ6yWM7lyH7tIsvei8
2EJk3WRriynp5TDXC5jPuwPJ4+P0hPgnUXsctK+X8AF89TfXN7C4IcgPnN8+hV9A
WLVWbdVhlrEUqGo73rBOWxqnmc7Zrh+b0Xte0/1dQxqwWz8W5yPQJdI/QHFhiweH
NqsNdjj9SvJ6zD5VxnFps2Yn8oZjN4KrHibtWJFnase6BXrBA6J+C182iHsEU4M4
aHWUlFJ4lJLHt4d/p67L4AL1AK+MxskDX+6JujRCtEBJ0rrsVl4L3KkRN8a3UUBC
lBaZ9m+GXBA9FJlQ7MUhLWws/nkrJrHWLOl+KXO6p1144FiD4sUKH+wuETvZvkss
zB0iv/LG/WJUmmXL6gqX+a/xgoD57OxodO52GAfNIIEw8WwPKmLTyuWEuGrvhV/i
9AChjwW779wU2s9KHyWWKYQ5co2iBYfKTJD/ekhHS4fJiE6O6ZMX3k1fDvqo+FJA
KoPKKZ+7iBV6JlOz3SdeI55MeTDfYJ4Cc/pHV7rcnTSPmDX/1VMbYuuUIUuC7aA4
LWkVkUU4Ml0KVw3GR8R5Emq05yzkJaLT6ea3XRExDB7bObe61iXz5KWLHvkaw1QM
k3JgGTYR9Iqiq19fzfMKHikie0iMvYgUwF08VQ0bj/WpfnYq/HaVBQ7jtvm4zJtC
91+U7wQP2gLO4SGpYGn3c040ilbEIFkc8JXdJSgo/gDD1aVDrz0jfJs45nTF0HTT
d0jvW6iciV/rSv0bksrBH34IjLC1WCee83m1mE3JkZtD2HDHdwFjENsjafctY9rQ
176UYWzhzHtSrsDcUs8XRoXP78vuFmfJpy9/9o4AbyRNNS0x/FPIiRZCJd6RtZsI
YjiOyFj3BDSfknX+s6BC2uPHeV/Fz8JKoxF/WkNbhC9y3Z/ZsguqS5A6UOMVjmsG
Vr4NEepOECaPphyEBKEqCZhtD98XZDzr89SCWlGiKc7NUk/Bp+2IAp2lR+kwzBTA
w8lQ0tnkBbPOZhCecmgNFc/o003l4vs2QQfZTxpTpEMRudZa3QiRwvvGVJjLkJ97
pEPnPyCQDviD5lqUGZ2VYHj/tEXeXPxxv3++hOdpiAUoTepd30YlHv1e3XAqbMnM
zkFod9jmZiFqCVU5EY/iwRF7yXhPasb8RfSvcpinHabZPfCVHqN+/DWYExrUstFW
MOKh2wEd5/Eb0yA1lAwLun+azOcuu+OnU/R3jqAE1XyJJK5W/3v/kFd9zSwF3YpZ
YpdIGWixZtPWP/MZZ6qkyVwMZB6WSVu72mqowtoojmbtG6XleTYtYl32dfHxBo0C
uI8r9J/Vb9tSp3IMwuCST4c28q1qwaOl/4jOmE5YhbpJU7AnSEEPvS/DHADQ+hAL
apTQrlwzFRvx+qnG7UPXQ+0WBXAFldwize4tbm6uJ/R4Ej0uAD4Vw+Y57POtybHE
ym8qfvWUho2DVhIBfZ+bBXwY2InBD5ZlB0IyF+L/V4bbYS4UaTZgZP9Xz1Qv18OD
VNr3pFXKAcdKX2mxB1ynpkSlJQ2yRIoXkE40vbqSGZ59AuLHhWaCGKNB8xmdNxTU
VfTC70kJaYHcnG/x6hFT08Nu8qNJPVtk5x/aRFxNBs8/l0009GVrF3Fhrk8OjG16
mp0AkSXm71O/q8KFKPv2hMU/Uu7naMjD+YdyvHSB5wGz+CQQSEHmznVISDiOB2i4
zsuOLzRQ+TC0GtLqZFm8OB06tYN4FX7jY+udNQvD9B6gGoyRLVQty/GMFGzEnw2c
jMRi5pfgU0QPKsdZ0H6so5AhMihk5nfrKaPNwlr5d6euo/YTapzkJuySbkfnrMWI
Vp8/RARi8GhRrSxDHuCmIgi/e1MkgmctDny4N7UZ9J4BcvX0ItsMkEI2yjvZtEGt
yKZE3hPtwj3C/9d4JvIwzgfQbViHkgroVLFOQmY7RfEVXUMm0zmV4l+mmIvBnuaT
f5DyM4lTLsGRy3/JC3SEx2PKxJCGmbCOXkO2JRmdfMig4Q2EZ8qFQc+MRbeg/qK6
s3VyFYfYb933SsnQ6aYs9+EQtkwZbAbbQo2DlfhBCbMwnrhAJWMNxD6+XBb/s9Tw
JLzkHBpiorl7pqoUQmd1xbhGvWX9xZ5cTQdT2/E8mUqWYZ8VKpTIxTssXj0f/K0P
8fJaJM1iq6waJgVmxFUYfoueKUeHXh2YCvDy0qHCRmEEeCkMktQ581hLnzsm+vxa
+A2zV9Rk7I91Bm83BOSyWE82O6rtt4kri5beAKsRsuxp9U40UUHj3+rQK5hnp616
qgU/G7NA/aokhsCuU3bnOU/CEbmVMg5dMJHMJWLAl74I9fv13ZJcq8lY2iVVrEkL
dtyWa9TBJ5PJ9e8KqNENb9AdOCw45hnTg8veKHR0A+rv8CwxSzbfczQVCDl4/qN+
onuTixwZrwpwuri3PKhZ20/WPPR0wjhjMlmkHTP1ncMYckl9HGmk/9wF+YaM1aZA
1M6J4ed0iDjqXOONRWGuXcsZUbdGR2SSrPqYt3wxClJ9pqm0QluLQdpxeB7GDDmA
+vduo9AHCrQJ/Xv4Tzd0u6Rtbfpnug9rpASCJ+5OfJIzL5NEXfGKFRuNPtjJpEqX
NqjoqH739Xx7O9+5UiSzSYbgQg1HRAuUFKvVdWK2QwF5kSIV/Er68nLNz9Vs0Egu
9lSrc1d5UTYW85MHhEywF7HbmvacZN+UProS1s2kEH+IFJZj/wAjp2GThVD1sLnX
0nVrB3/DVwDclldXNB/QHG0kOrjeWB/02qhU0GjaPIZli+sKDJycWsLIGjAtGDvv
RQpv3j3CMBmR5ebcbGm/eSMfN66UT+oEHZYbX/sgqhGejxTMTUYNtzD1ZINtVW9B
jz/DFi0apobY+PMyCZIw1ZZS8pzb51em0wXsLHqYVdJu6toeovvDrk6F0Tn/H3/2
XCXSNKjvZcDmzH/7GUxbVYhZmez5Ja729Vswc2OJ8QQTr1vMFGqoYdRMCtTh47Sg
e5d6KKBjmUAqXfS3cVHLwFKWlIPZwjnxuWNbwZYGiuyDgOxO1oKNlkN3BmQOLpQH
z26hYR+7DkZxrsgPHEwdQac3Qn22o5OfX1whssWV1kgsWPrnKZy4bBgWm6dlJr+b
MQ3TPs/gJ9BC+u1+bNt7CrgURfQaUwI8m9q86Spx86LT6r/p4aUQ6zEslQZkd/0D
PBBRyq3o/dp44ot7uxApfHyLIxu72c/+uZqVrozEtLcpmDnw04EejyWp5WdE6zaj
Q73Xcd8jBRNvV8/GGx3fc0ZIRlBUxzkBN/d/3AyX9OTOi32h/BVO5Bk6pLJfvvGk
Nrk/t8JR+akPEL4x06bCbPhSS5Q/BCDvG09jK+0xQHvMy+t53b8c+U5O5zRRyfg3
8bVLtCWqJ8+tGhOgfkWW6nsU3L6vv9pEDrC91lKwSOOtV/Zcm4kA8S2QzsPRfl+p
a+gyWK2yH0ts7BgxCocxNEJD4bOrjtWDlinvUFb3RAejPq8Qtzlhf7Nk4jvRPM3H
pbQM8jS0yD60kicXyo3u5qRrCvrM3J5WsakrMWtwFUoAL6ax7B6UENv6O8q+Qffw
i+gTXrqhzCOekP6njMttzyE+4Rd1QE5ch2l5xsHcK8sPU8Lp60btsO2nVOBt1gTS
9eTXJ3/893/mUTmhnvIRsw1xYS6bYVQqIFDb+p4Ye4zz1RcJ5pknk3gQVRRL4XT7
4KYa3p9oraV6aMaE9zpMIx4lFNLe/PGgivYfYE7HO2Ty527Km4DdfGxzh4sl/CA8
/nwk66/eWv6eMDeW0Ao0a7aQW0ZEzqQbAvfp1fLyyzIrcMlb1mYqzkx5Hqza8MoH
fGBWzMPv8PeXRKo8cok+J8FjJObKb/T3Tg7nuYulZSKBVKxDMVCM32REOOzz2cro
Xne7pMAMrQaMrikC5spr298p1QxYPuT9BX2o85Xo+cAclpXpDsx0TwfWVbVygyct
Eqfc1xEidr+NlIl5SQb5keogQEmzlm6KxnhGGuycVM4HBVmhYzOr+hJyMA5A/ZrZ
PdSQeLiPrYgKYngJU79qQ607jIZKjestesaMs1fDzYslshnaDAUfZ9vuHCPcg+Ya
3oUWqrsEi6oRW3ZVRBaqAUvpuE1YCR3NcQUS/vYHjVNtH4b1i7TMbdA5FxyOtqu5
8anMyybYq48YZhiQ7yNA9WL2q8yV1LfwtZ1k+n62MiIoMmBFpZrZotGbhopb92Af
v9QmGwlS/ExOVPF723yaaBjh/t/8EXy8M8bB70nh20eYooQ5+ey7WoKYF0jYa6JX
wr0so9Ogg9vFOt9jjavAxYLRan6J9PThrJsYzTU5jK229hPDuL/pb50NGDC6n+K1
GfnC2S+Z/iE6FvYVNJiyrRRIDhvau2FbgJxINghcHOYjJQU0DAgyuN5zY3qIexUg
VCODw+WgTu/uuTx4oBKo7lAhRzMFokVMSOrYhgUjqzAUOyDlfWgZMBIjMgRaldF/
CLRdaCO6f4xGDjPQ0nxwirrGhfB8Yls8KOIVu1ja1g1rWZ7zrA7LamkX8vaF0Iu1
ngJNfYjSDUh+vRRVLtmpvzrabtmmDJe5JkQYLRL7zBakJPKoGBtNlNz9iBJuEN5J
kIK3cwmSL6y9bOsk6Tk/CdYnSTf5oQDW9Lt4RwNFJ4sK88Y7aGWVBTHx2MxXqQDb
RoARhbT9+YiOk6AFd4dUBodT3oub4nTcyKDR8rn0tc9T7NSUX9qJ1ge8oL4dYDaJ
gIkQT9BzMn7zW9LEbSrurY3l8DoMddnpcZzLwmCYOI4nAF+5Wr8U5M7kwnK57Idy
A0wWxzFbPLppvYPh+kEAYwhYZK6mdmownLb6xs735RvJJCfIxiwNXjKC84PmBxOE
4c3JOuBZGmijl7GZSBsnNYASePX9NkfM6h/LebWVKeSSQ9gZMb/6cGmuIvrIIWZM
nbBugxJ2swlKOfBeV8jKI/GtPm77qsC4vKoIIEdjdKqz0gafTF66qTmeYo5nqM6w
wFulkF78rFtCkXv3sctG0rlHT58iB6ygZsJaXA1xc0Lx91EJ5JUiwPgDLmSa84p7
SOLTRYz412IkZzKxON5rDqWsr71d5weiJVX1PitP6A8lFm+6f/d7iCIetFo+/NAo
z2mlK2+CNky8USRkyED4T+EsLTx1XRvYHU8HBkPd8WxUAS0ZWuU7LNpsz3VKqKZ1
7Xf970ykuLj6EqGWvewFrAMi/t8vyDgVLLNYhFpA8kXrRVSwsk3527zWpZMPPhmP
Ag9mn2OjmBESG9wrY5zIVsjsj7ho90LuyFmyygKiXbWzMXrPyV9prl6uM61JJ4UE
T/AWoZhm+BN9QrJk20kC4x56UAN0KOhjczfjiIW2OgunIhiFFTvLVc2D23izEsNp
v25sPTlvuxbkxH+jzf4XvUEWfALOvcmMjpjNmulFwb3nN0XMk5giJaTgnTD8SB7w
NAyES0OsJUda67FxWh0oBpjFz5oxdFRxYagnL75PNaj6wAcGTrjkwnySbWupIW5W
raLrP2JvMdxoRoH4yf+fmq7JVPeOCwSpyXOQs4mEMF6O/UcKF4E6gOqWl95zb54U
5wQbMqzNruDi+KbUODzP5qkWtghHRSlzZx/DTKW/6L7O3apW06H6Gv9ou5zccVAB
Ds0OCvITWBOUuNdgSmVOfCESiNc4zvXR8q6sUR4/nzunnrOExpQk0j6X+yAX4hZj
Et6tu8k7IWi8HBXvoDgx3IxZUNO9YnsdLbAMtj/0RaW3vv8wm5Y16r+ofq9Ea5He
vv6fhJidx9aNtoHk7Iifg7xf8iktuc83gj7tPn6WeRkKvPf0kPOCrzjg8iDZjAr+
bX9Fu4l04eXbbwfdQMNp3kj7uel7F87z2KohIUX6b/44Zh7IS9v1CmIu2HMvRZ8s
qtCGh+jo07CszBMpDfvMnbGdTf7Bk36kRyUwJAKuTthvwh/TNob4oBoU4ob2HOzo
l9MDYLxyB1FVbbdCKM7n1q/2Vl4JjLxp1MlTvWRU1sQI5lr+ZnDHPymjH1c+zGNR
2SIdhOb9qDxnMN3RjJGYgQyakEQ+WrSw1h12e3UkiCLodBpErt0432xkOqiyYdbe
7Wo5F8Mv9zX4hpX0hZrnq1WhkysLTRNU8msXwlzX2mQPxzpjKAAA2WGVBbRTcabT
SYExOpb6+SsmS9XFOyOkxLOOOYnMlo5zyNkyxw4ClzKtFDVKmipGAYAF4iMmEeam
CJI4MOKLTLD5F3PzONp5veAnigk6Cp6jh/ILsA5f1DEvgxsdc8i/ZHO9Ccj9pXyN
nfXhi+CZbnZUlupA/UJ4rqcyGIIj8rHZX5KPLUSVQ8OpW4AgJ2hoI8cv2QmMkx8Q
ulsDRb7jjhjsb5ruu9iikVpdvsXJnjxDills4PGfbqUZwn7e6Fgu+nS64/gn3U7h
nhS6fPmZnbcOFMg70LYLVtUee9xCewbDKZCXYxelRfccOqwywM54riSAQ2rZPlK9
FZ+5RMH0vIHoT5d5kN9DLwyA8O5+nKPtKG7KUhOnAqVN7PFY4CyyNWE6+N87WO3t
7JlId03RCxJuSmYPWGArjdcPbZDKtSzR5jmwQKDyngRSS7baYiBkneaQ/Bo40w5y
DgcnfkKL48eyQgLRbwICbTpvVsI0S9XRrEhA8RqeieQzxOr5IqWZhUhoAQNJv597
CoWoHxS2WGJEiTV8JGkwuY2DEJaiGwwCsGt5SQBbgx8vc5ray/tzv4hL8bnbLOvX
tB/lrnRbIMDwO667OzvpWpeiWElcM3vd0XUhIYw18T776MzntRDTUWm4I6L4ZPwt
n9Sau9L7jx1SJhhocqlW+Pka9vLIK8isU7YhpR/6LpDAgg52e4jaIedh4yBq65oI
qaBsUJAM9/ZOmpd650lHPE7Dfdmj+Xk08S9PU1KBSRl4dv7YI4jFtTXYBMa7lOUH
aJkYWYIcoqb6pyMNj+7CQgqkyFJ0m3HzRS0PB6GYW7saRifCnUeVR5MNsFEh7oql
LsxNyzBXqgSJM+/IaL+00wsBzzTtjv/57r4saHOOGw6/E9Nx+0hchtq8fdBMlhEE
71yfsCr+IJs6br40awGMgfXYgWXYU4DRkhSUOrQzgd3ggScIjEnjIwtqrJsHhCgt
QhcKhW4SASED53jsaOU08XiaJgbDNc8AOmDLYLmT/K5T2JDDTy9euRLSwtGc/gE+
45+jTId/uP1yrNPVUb7Xc6/creX+A8dmCAFselaOLKUEIcel/1RMmFZr2HCQO90+
HKSyJ6a04gEvxCLZyQ5RBZS1+GMsTW/1osjj7lBqzvlcak+9MdB7QZC3urRzy6ko
Q/mVyFWX4k0Q5aLOIM50xj0rgL4o/nn7sv6zdHXsxjX1yVMN0Vsj7JjYJbteFvk4
20LwxP61lSwxjJfm/04GDeE+m73YREph0eDM8L7ysRFqov83JBkqDh9NoIvtspY3
/1DtpcZlRu/dXguKgP20irO3F1sIdhua8OZKlhYM9JqD2PKOg6Z1/iuf8QBftxs6
xLXTxYMBqlvuqFlCvgg041ptOjVIEycXI4bunGAVDSv+3YocbU7HEoybcLl392P7
6dim/kMp3ve8+Ph8QgblTjYPooCFa9FMXQ3oukjOY+sZL8/7Kv3E0H1FNxv4SEkO
xrQNjQDTmT55OLGmhKXbYom+Xy71X+tyOHGL+ayHDMaRLwiEirBsmKdl3XfLwm1V
Ebf45aZNhjIkyFsw2TH+2FFiN65DkdrHCC5g9tmjR8rOO4jBImS3/qz8GNsgOGl2
hp81pGE0Lmx6HWzDv7/wVL2fmNISgWBOGvpYT9cI3uVKGo29RApuvBMXpjDh+KHg
wo1bwfXRVm9ovNLY5d/rzHfZ4bbOHfrKcV16nN2pNTxcDIdDqYytumlTqUwzBZzv
2t0qhO8Y0/m5OxdL9jElkvs+YsAB6+N7/elDVZDxQ2sXo/Y1gNkU0vzqY/DelMWH
onaP16o0LFAgeFBJKjpbRivb+zqMYKD/25PkzQwNxT4IBfFAo10w/35qVPF8fj8B
UZF5TD/VVLpQodF87PC7dPIJuoTIaVgJY8HoPU72+iArXBwjYQA5Q3RYfEpQpkuz
bKWBN2spi+0WUS1MntsHNiTv2e6OWPJQ9RsCY8lrZlboKm0pDjTXkvyz65pPcVSI
/+MltHjpIlPMsNsye21vzQVN6JBbTrs4lck/4bLoYPQCp9ugznuN77Z1SvuWtnf7
3FHM510E+5mPOqb8N3D6s2foKeyHXT7eSp+kcwdvMuV6idbxB+tJyZ4mQFGfsshq
tuEwX6o32yYxUuv9GZvHrKNgJAmFuted58u88DNqmq0VLamC9YGJdUVA/JDi9r0b
rXMeGTWkelsHSarIQPOFAOB17VdCa2twks1TIuMCdPOKmM6DCG++UmEBIi+Zb/XN
+5rlR7I1SIUxcuwLXctIk0bR7cUtC1NNbSZ843ZLSiJUYcOPrPZ2cgO0GiSsMvL7
hM8VPQGGuOaK9JTYOwLz3ljHm7TTIAHxRfZE7gzwQUYdGXwP512cmJICIWRk0OS2
W4vV9nYHBYx3BZfEflflXREcfcHQGtBJWhD9fFzid6Uhk6sL5avHIkyY3wiuzx4q
uWD08QOaiDH3qKSNGwdVf7NHTsYK2o0KPa7KaGHUubMsXj8hJlcdjaYX/c5tsLKA
Edcxvip0AsdCPaMVJvvJxMCvcUANFecg0TXeL1XPTVGIOVnWuVwCJXQJTS+lUvEg
bnyg13JDgsow+znWcvImpkNTg9rVFfvXjRKcyYYJOH6iMTgpY1nCtD4aJVO5NMyq
TN9mii+xPY/K8JQ/r4sWIPYWdSB4pNJZRqgppLcLXaxuBySq8+lH8s3APGvGout/
aDMnbvNS9PvoqGKE5LxZGYAnFafnE1cH1OMYvqQzTrUP0pyzVq7DhbZcvK3wzVTi
tak2dzJpbGx+XDhTsnmQzexx3dzhNpqJxy1bHgy3mixQGPl8xnrt3/TawmlSHbiE
f4PWTkjU1Zf9tljTZgghhRLhtlvQTUJ1e4adr6HToZrcDkA6qV3CyRFrdsopC2i+
tH1wlaz9XEEGSUyvA4Wk0+dd7ilxcjGwa5aM4j6jz5+2vPDD5W+4h2STGRXuI/el
MOz7Muv8uZy7Hk2OMXe462S2lfZOVv+QcZf2yyef1aqI51kSViYGTNoEc4m3T9Kl
R2419T6NMIFS9ftJDjfKZHZHd0S7vduKRaeR6/j0goKiqF2SvrpZjTQkrSG8lM7Y
Ld2JY62G/sqJHwRWyqZ7CwGYFxh3hAOGCFHqYg1OYOQXt72BMQUtKBR6mccVfM57
RymGM8JXPCbEdcnZuM02DZ8g5APSoTMLdAPislVEw8bighpmXWJpzSwU4RMUS1iQ
RUQvtEt7NupxU4TL0bM3rZTEssBHQQgdBshfvTQ0HL+L57Qeke6cms5IE4VlPO+g
l9t4X/0bdvlY+YLfo/9X5GmfD0zQYD3NZdN38zdnFDJAglGO9Fp9sYyyG3O5NA7l
W+MqeRHvU1GxkETK6v5RsFCdtFqxy48MqSbMzrtmDAI09rDvY33tAKjM2mLxKluO
fS8hZzI3fPjv4u6MYG4t58XJRffmDBCqSPHRrwlR9WGC+GIlniKfdxBqh7tNURPc
Hfx7he+i86MBxD/e2OwmhdQ2NHWfHVZFC65j4q5R+Fe88fiUokhRVvtftaUDmVzr
v073plzrQ3+MunkOWOMyMdC80Jl7OknnKmQVsJwdf7fWQ7a68bDunCbVg7aIPFez
l7A8gdE/LJuvWxzJkJN6dO24paMcaPoRzLb3WT/7Yws+dIK+w+24wsvBIz26Lxk1
TDgSoUIptFUQc+7BTxHYvanEQHLaM07ZH7NgkK92LNw18NksI0p6gXy7RuYf3e42
SgbD3Txh2lbv6JkdoPSrWL1UcXIwz+FK7uHpkG9GkmfbsYiS5q4+Zc44+i3PIAR0
YBjv3Ne6rjxPCruWIVFX/YRCxg6xWlciAH4fbFnWRE7roQJ45U6vBM93NwH9spKf
FJG5kiYPhRXFC2f91I3CX/Ng3zrdxKf2i0D1zvQUGJvhMdH3QeYztG61vw1by7bX
bW3YFZlkBakPjs8tUgAjyuTUqkvxvL+9Pdk4+ymSPt4MfOtIQ8SoV2ctVG0yySDj
r4wEYajYkGKqJ2OgZxyBFCjBfFgBf24SpTWgHSpkvDwUMlWGwrulgelLPxCHpO+u
Pt5AoVYvTXzRSxzRCrx2ItTz9w3pkbDd5/LYfYMebTUeYpGwleScM3g0DXLWL8yM
0u8Q4LyicNtN63IYuAz+k96V0uQvyCJGWExOqgnxM4y3QMBt81rTGt6/iNpCfnhD
vxGQrlPSPugoTuUkcP+zjBCkaWYkGA/BEF7Azo0sWsyNRFWscmpcYeaznWL4VKzX
Xw720xeNOaEaMhabI4cT+nleNN+tXScarLIKIhPZTE8cbUgRyLfGSklmImzMkr0L
POvWALXzLLU9lhRFeW8Ee/l1GK/rTUWg5mClpXvNrOgGoeWXtbsiVWuodIOBqTIm
rYDvVEG1X5yQjrRtN4Q2pz4NwIQ6HUHsjLWe8RjzekyZc/GaiczBEGHJwvHmf/6C
2BrE6gggbAXtyFiQWdhdArAFCVCUOfgoxtJSpmRGQBT5JhEPWOGU6VlKNSE1806p
UsyH8g5P2wTsrGNLhqdtONWBLHBHkFMsoxQyyCVtWAsqk2d3IFH+Y9UjqFkxa2IR
YxE7g0Z1xkMPnmPd4F5P9AVCNoUFtxaT4w5FOm9g6Arko1CNa0SaaZC6Yiu3hZeP
oTbjP/lhBoYAMPR3Bai4c91/rckj/fGztHuZGNSC8SBncdeCB0ZcD4jY26g+Zueh
EKMXahzkXwDA22tZUKaejW603O/7NSAg7ufFYIGZmajF3t75Lke9Ax4hbuv0vUTF
8C56VssLiq9MKmB2JOycvNhOp9TfIkFMEV/BNP63IxED8gx6fuueDZdS2cWpZR1D
jLQnPpjnYy7qeojKJNT35qjEOeOt8SPWtg89i13prXs1BNi5575NIffId9A6HxxZ
0tq9yPNri68L1P67QtYvAEx61dsY8m5nyG0mdetp8WEcjUKiCSGrx5twRm4mPpXz
8RBT5/zZmBn0Oh0mniyHIWi2td0gnQS3YfScx96PsytOsYmqoZ8WCpUqxklSVEQa
IU2aDSUBunuCyw8W253XSvxd5kZAxkk3W8NiTuQFAjBlYlp2SkeFoviJfQOd4F48
Oey1aPaR8ht2L75amYw4IuUzuYHGspO0mq7lC4TZ9VdYteDCel0Z5eWlQId3gAvb
vm+1HcIyx47OXrkCjNLwCqB46hhgfxN50/YARg86M9OMPiJdfLjhFXggbwfrO+zz
6twDZlubW/oe7iJRR2nOSsgneVIq7fjJknmy8Ls3lOmN4o71bmGLzZSYSX5avmiG
lAdqG4HxIvEgHlZhlx2bgH+xatpwoZDlTbAxru0vFolS36bBUMgpyhNEZYtU5axR
0rWKkfBnqpMFlIkVWRSTemtxBO44BcqqMYdW/ozPOyIky4xH7m3HXmQuBdl+bc/y
OQHg4K7Vr4mB521SfQGiOAqq6OYWhPoFQlQsXPmOseqfzMrZjQd6PT6lhAY3KQ8r
XttcTlBhJW2R2Ko0/Qkupizm3o3h49cvudndDwsIQv9jpGd1nlYl3PoWOKdfs1gQ
hO90Yk2otpRl6mEAcSYwcVJhXgLNx1yhbCy1RGwujvmPAo48/n8pM0xDpuKJ6XUV
KVRtb4NuIiaE8TGO0u1dZu7ZRZ2+o5rIGHsdX/Dta9dHy9zDXvI90hRJBJIfX/US
JoeNumu1Ee2q2TZoYGSzeqQByUohVVFzGZlGA4z3f8W33kOJroDty+clRFxrFUUK
e+UsrSFQMLXbRLtGwFVRZH6KLgllrcImm8AaDL1aQOEzlbbZowHl8yvnrrPeUDYn
7duI20aOuB3/LbOhc88/A3RsvajBm7aB7sShGRGDl0FJ9GkBiJwpwg6VD/iEt8xB
8KBBlWvTRiSGqgBtS6b0kvREOekrpFVnGyPp28Yl+cl0jJO/QgL6IGUFcDkCzPvg
lofwcLKp5gXWFVYzy47QtrRpiqk7S7voYTnk+wtC2qetOVfHvv3DPcrP6hplAoXB
BaSJhe08eFuEJKVo8l399c4b++YF3D3c5lR2FdxZ4oY/hWUx2xCjfmCzqdee0tVV
5JcruH5loHVOlNbO0Hr45KB3zVIWuUATYQV+bAbNxEZkpDiVH2l9LhEiR26plk/o
lSnnYDM2OPlPrFPxpm+ua+XyY5udKiEe5JqBng5WTQdnRYgRwWlWwFhVESFATMWl
Q4JofVA3+tIvPHM2DSI43yRnFKmg+dyeWg4Hi+jjTRO8DHTA6WS5tyI9tVLaCEVC
5KYem9Jt+slFQfk4O1J2Ob498JUuKsefBvr5fe1NGfHYaG3n+7aU8JWABHrhLsXn
AdDQj+SfJzwyKZ2ZYZ3nbqdcixtm5Mi5kn+yRjZoo9QZtHsE3K30AmkgXjsceq+s
szOQhuKLas998qTe1ZjmYGW07/Q6APjARb4n5ZTPYLHdAKWMzsZ5vHQ6SiNYzwos
+/ICcxzCsP2E0i+draAaM0WV6CX3pkcCIaHQ0VBU4ID5DQJabeEQvYhMHDCIpA+v
bYB0dO8v/0OmRfA1Ct6IBOnk88bQyWGSy3vLGyMkbQK4BO2ZrZsFp4bm8xMO4LWl
Ok1r2CctJGmlqw2aTa3LXDLe9CXyEIntJoQJT7adUDDiPSoumfjSVMdsYfP/6o1m
ZkVQhA+TZ+ecvBum6HzuagXMUH4Q+W+BYDJeXup+1iDYcs5TnPQTLOXhy+OumFh1
8bS9nRPahgK65DctoeoFteGnQ0nb/3VfNbDMxOiW82HMbpm9/DjoB3r9uAQUNyX6
lAENHc3HvZbUzs5csJLadCvBZWpTj5SxwmhVRgTVN8Wyg49XwWtEtpdRmeAqe3b+
nAvGVhhihsdDGNIQM9yrjFbc60mOcsk2WXcdbAws6nDwLwLVCi0WMGjjaoLdjEN2
qauf8Orp870ZRpbWSPQDTiCQOh77B3Vf+1up+PO4hImD5Nju0/hPZ/hYlyKYsJBJ
RP1LlAEthbjt0NdglEsl8evOazD79bUELfHeuPHiggYVQ4kPU7H7JneStKoZwjxt
pZWaDCSfWGZIAB+uNrCQ0YN82J7+GmaTIOQO6jJgdoK8zVsbHRpF+n0YN7yf6p82
GWYrunt3MHMqA78xAURhTe9HXGHnhJK81QA8mFTcbsHHY+RSlJNXaUyRlStcnFZA
spB049qR/n/OXgEr/jLsCav83/osl6R4+g3AV4wfANmj8Z90M+f4OrwjTZLT+0HP
BjovAJrwrCJoZoYyi8eEpc2NIb6k7YVWb7eqW6u9xdcLfzcUovAHDDI9MF4fWdAE
/Sh059NymYqw9gt5dIgKGSEyNi6FCuPNlaxd8+qLEfSqnSus61upgAtRtBCFGw8g
J2MwtyrNSlR6lDIrowXOPzFyVzNW1+UvvHtbBTaPxDLCy+IsZfvxT7FhWggfyr3l
0RzKyRpSuzzv4QHjE0LEodpCLLP0gapem9lUoROSVylOJohB/IxkxdZB+vB+0K6l
afSkHlzOYHiuutHoA1bKyiLLNbArnCfe3zBz81vmqXC6MrpnBNzoVmHUywWpk/ra
7F/9W9FbgFenlHAQTrulwoMbpiX2UwIPcLe7U+rDyj1D/nbNUtiwm4RmoIdpp+Hr
hnBJ0K7g2tblJ5JIbk17WjxwozIaQQgHkOFlI43LLcq8W3tG5FUczKVr/3tec2/c
KrmS6ol+6sHZkLN+29Nr2O3iYg63fB+ErU2SUF2OsS2iE5xIhuX8WBvbPSfpX29K
fr8/6iVUYRtDAeoaNVEVVMM0HLVBvg3Eeu2hrHj3q+WsVYlZmBp7dKG8csRNYZL1
619g0lHEXmxOXJ9Dv5GBfPwgdgYU/ZpaRKVZIosUnvhRylogeZaSUTsVyh0T+yYx
qK7R+LLF8dkfZgEjJCtCSmPa80zJo0o7zN9Qo3tMzq+T4aKLPKz8Hz5rUxzLfoLJ
4WC4k7qaUvFxW10gv/o7P+P4TXwm8mRUHQSVXd7Ex/LG7XezGzzXeyZzKLbhCSAw
xLsM+PgCql1j4R8ilJ3oZmG4sKDBXHjMwMnit8xhnzbr1ioAcWKq2dLaiBRlUPWN
XoKk+ClLtxAXhVyEaa2hFkhZc5pVB7emxTDAZfiVBoHs03niDEq3hlXdkZsTLaYw
x0F7UYdA927sRI/wzNCcXvEj/gyDQj7vtFhtcMGikbv9QyD4pzrRTTUGGWge1pZZ
RsIDUl598eExDBZuGwDsjO1EiqAD6fvmGDby2VG074425ag34KjfoxFO8fVWaF0u
yHApHd/hwrMHf78M6CHXgyPKnXC3L38eUKJ7LR0QWJetKOL33tshVF433o8O+G7P
YBZ+RkJ5LXqmSJ3Xs7UdJ3MlPEsuQRYjX2np2rwyPgpm+H1WL16lCtr/ldMYdukx
uD8UUOSm36ULvAPoGsdWpHaJHYku8koKrPCUmUsfojJ9pYE3Ssvg++gHpSZdQ6eb
iragx/jU5ZoTmJr3piZ29GzFOB6q3z1eiEh5XIc9f1xQYf2P6qthPdhKJuDyC8uZ
6eERmfnL8TvoDKnA0JflxzyXUvspaMhuG7KqcfchI3cLr4ux2i/NmsazedSpV9rm
FBMVqqbrUWQgjaBPySeEFPOPvImVTlTJdun4N/X2zrX/E7tkLkUyRGKY8g3QBObe
THl7mN9iLv6rTgdyOYh2fgocgkD7vU2UaCOz9WeYUqypkz0QismG+9dVDYym7ShM
xlsvdaIJ0m8kIvoO91u9iAS33jTHacFYUREWo5dOPixzcWgb5+XclPkxY/hpsqwe
fcmP7oaPjxtjtLikrJbVJER2XvRoFBHq+0IV81DyiirkxN4gv4PBHEIm/DgoANqW
s9smSx1ZPQtUmTuOciw6BX8NeCb0i9OszfwiABo2Wp/1h1tU2Bsdm0G0cunIR6gm
HfXTylrrtmbk+fUXarniFRyzi+gedhjik/kkcYM3vYvx5Js46SDvi+IyKX3KO3od
mPmuOiFytSVHEWHkkOtZSNS26pLR1DDggIpZbZuimOfWcujWyEzE1ATYww2p8Uvd
oTW0Nr54TZC5kDx67JzrKNnAi8o0zwWG/I4Ed/0hxtIZ/IOVX2kbBhyJzgr4eQ5e
Tg0viWCAi1qkOgnjFEQNmzltIWZBgFS+3W7KaMwx1/bXpwGqgkuAN+UB62U3vf2A
lqQtKsGI7cMLg0ZshV78ePx3vgu61/UsxQoWsYlDegGdCDENbhl+qOks/+j0i/Wi
RiRMURouVKpQRzhfWDnmZ2MSY0IWsXLAc3eluu3rkk105JMW8F5mfewIFDoyF8u5
b+RBPkcZEwNg5ZWntQMuWHl5F8UsJnMdyer8OBYiWNjnVCbw7vWDBs8RmH1d1IdZ
TfzDcnKcN2RSm7mY1wC6RJ/WNxjCYCt70ZcSEacDWxfja3law7o25ct/zgnscjfB
5PFBBuvjr3y7N/FR7Oyos5QFw9o7t9WPlwDKBpD80khsI1g24ApHupVuA1o06+oT
hUJm2io+pURdhzHmf/hR2mKS62bUuVFjWlyGtz63WiQiNTP1zckYpduaV05gug2r
aXFiKnnRcEx5x9WGbPJbc997i8c892drmnxfHPS/I2IzteZ4n1jZx+4xXZiXG3yS
J1DRAcMNTmXJyb+Tg9UVCgyNYgLii1LVtEBQluK/Aacfm9hAbc9huhNl3wK6y4eA
gh+0oY0WP81iiCjq6b4HrGZn5xl8dx8hojyITjPcViN6Ns6ak1Bwm2MAoc4OPi/v
eXgoqaUjG/rpyT/eh34ISY+NlD4hb3icHr1XkDEl5hGUWouSLlQf8IFDsYFLoy9r
4HNxkj0LUF1SdBTQEarkvf0xhraeZVC+3v5G8QSUm5RjjiPkDua67m4UaLrjrUR4
kfNE8KNHFhRpzKLGqrhGcOaWFSLZ23W3PP4Eq6TMTGkJEk/89nqfNKTuB8KBtpGK
U9tn12i0nZK8KCEcKwJkU6fLq9qfagmjQRdSKsbOHK0TQNm/U6pUTYQyy0qylJMX
Wj8wYDU3JWy+czXnxYnCfcIbIzNQVsRgelkssLHXLED0NFePdxddTanMdeqV4Fn5
CgAWlongVUGVhT7fLNjK867hVuBpNWCkqcT9eo4JZJtj85VyjwJz87BOLgWjXTZv
0cT6QlomF16r5jZa7bV1yKuV+opnvL+Bpdu6aKI4+zAu0b2Ttzwd3wYFFDkUQDIg
row4z4sAkJQFswK8qcS993SqxxRYIMJ74CJADuAKSzyOFNupvRCl+uB7SuWeWWb6
AWY/IBEIgJJBsjynzb2QmBpMq1TALL8gl8D0jGSwiUeWXumIMo0FwpnsJMnI9kR6
lWRLifpr8KlAYE1HjtiwVREn7qaK3knrr/JKd/y/PH+w1I9yjU0HoZ3HdxlPpnz4
DR6mYz3ZLP0bHinadqPjKa5T0KcCL+4fXZ0iPAfbvdREEqeglPRY5enWyUESUBoO
wi5aXpj7W+BkUxnTVj7jZm0o1bx7+4qxBbcoeQ7Hn8Bvh4lkQ8jUJAhvOSigHvZa
0DWhFNi4Ba4EK0MztTKEwzAiHQojoc2EHdSqoSzcAbB+LPSRfoCWGsposH8610bN
3dUbWv0CcYDdoj0OsvRy6815JwvsXK1H960vd+r3ylwfsG1cB3vUYPXL1xwGx/zt
1SZTvfBKIhH5EBblqi0o4KLOIXajT2Csc1+kyiUR//6MKzVxNxbYRFFyRDQjumhp
pRjwu46Q77Sp0BkQhic0JPtDPOzYAXjMDZxMdtT0xWM2RwtKda+DaObstCvA90ni
wF+roVqkh/udubDeVhrh1aBH2mtIilBHmGTPpKklO3hwlxCythgZpYaFFJqahcWH
YSy8Kd2S/SkskqyZhSUrc/3i+9R3xCBsvyqOxPgou0vaFKPulWpws0IjZBgF2qeB
eiYmCsA8r7KZzE2YYlJuV01cOneCGJY2msAfRey8+JTeVroWITLmj606Nd2ZDdlS
F7udSN7UN/U75WBc+YFbRzG9TiiZPd1kxIM1TvUa9nOny1v3D6ColeQmO/6fwIeW
XA32xA3BQCYojv2KcnlweQaKJhvL+eDaDYTkJPhbKRoK+TR9x2ysTwPFUrkcN3bM
YwPDkfPVsFPxjpJN+QmDdTi7TtW3tI0yg3iFDS0sjwo9YgIGbzaXweRI42dg/qNN
D3i23MqABNXQaa7p7QUO4qAJ/XTbrT/5cRzB6yaq7jvFM5OQYgKfywXSrcMKKSHW
hn78FRfUqyi8WZK+gOP/D2YRNH3M+LQcIQ+MBQII256hALUa6NFMWNTvfxrmcb3d
UXIjNLmmGXe9QfdYPbpajiMaUVa3dDnbqeKYxiAWRXCepJZEQCMCOGR7JpDq0hAF
L67mO6pDQcaPfR4MwaqJr8FoAqA2DbIqe4KTwOo4S32urrm1XMhe7R7+oFOsHK3e
FYtIIuEjO81GVHMNty/Or19Zgik4WmuZBkzr2Br/KuXAFcrJa8+Hbl4V8LQMkFs1
/9nlWd4UelPB//VB2SKy+bEyRZRtXdVcInRa4hZSRg9rmHDmEAg9rvdCEbIExhQK
e+Bbg58bzmiDRtG56vaOl16tvOlYzgE+eRrMle7xJRBrtjveCTBEPZ8jMAvZKfvK
9zpH5u0Fjh0xceCscgBMYxIwdlPwgiDzFsMfCKrq8gr7T707qigM8+s2JpkoEh5A
A0lb8yhBcGx6LX8K91QhWbpAMlvsj3DY7r2UsFDMKQH0D+bZm3FT7gx2I6a7YJn+
Vvt+Of80hCLEFFtauvEU5vvvChY9t+SFV2dx5lNRX1gWykyQhc9XXwFKLSmOShS9
0emKIYZFkH1qxucqoJEysRqcW6B06YU058TEzhGSG6NzQVhBDa0lqT7arYAwebRf
SA07+UT0/PSEGii+CM23F5b7EKLbXg1MWoPLJ3eYV00feeeI9X51RhwuQG+Z6mtG
+H7gtD/wO3D1H1cu3tbE7YpGJW+Rgm4XHXzhhinAh4n7CX4lzaJL7DfPFFbLdYCe
3DVLls0XmxpWW9FHWMzVh5WvPlxOoMEOEJz4BU7duZ4Ub8rStOFHhfUlyJINDZUs
f0GDmHneEomlBVs4BS/UNeRbgfxh4ju4FeUjow0tbXMRQ6zVnmU1CD+AfHO5ICfh
5gNi5QJPMzF+tlSercY4XqUG4PriaNTUpRlrPaPMj1VOMbvtMUGLcxK5OEHVziHT
I2RQtPdfah+0TXCK7CTcMlFi3TJa+Xcd0VKxw/nRtyl4bVavKdD0Mh24S59zb9Wg
3YVTpvGKBojEfx6wZvguU3aguHFKWpto/H68Y+lcZeThqeLoMwGO2A1Do12wDo0g
HNc9v2jfIIDNX0ybSlnzIaT3ZMGMOeRt2VKAWE2WSbHqZeCTss3+HzIWU+nbMXt2
o5jWhKVLBd0LM76LNyTT6PjnelEogRv09gURDbR6/McC3NLmWcZUrdgwcz65DqkB
zRqfx3VssP7C1QsrLfg+NIIu0+ZvC1Y8CfrwGe7SU8KHz+PNjcsLtEbKLy9z2I7J
1c6ZV/zQv+vFMaFbzP1CyjbYTD+oUEqvBCqenHz697gSX6IFkkmWSnxfZWSazSAX
9ienblcvbPzKXLITQDfyHuDp0/OTZ8VNG7G8978m5Ovt9AbYBRLyhv5s3aFrTwlC
JXEi9gWVNp19c2Gdeas6UHgLH9cc2FMn7ruCiAlrKOi4FnrrgKUbAFx9mws5G3rW
gZhQTiQKNC/lzA1wcQRWYw9nxZNPfm6yZ+ImxOB+fTW5fVnd8uYwmld79cZD3Imn
fKCFmajVA//LpubAgFls/Ubl5Z0zpLPWwjbLcwT3vaTqLUrt8MR/ttBZSoaPqqmR
ZUVas4OPUvL7p3DpdXPKsse6ELH+7QrG+Bo4vMM1X6Hzm0rFP9MXFHnNQtkgA8No
j/0dxqgqOKdUd41yJiTGrOIg7teRU5LKaLoqZW0cdJdz0Q3OeTWkRdJUxV4UnZnn
2tQJOFBJX1J8/JAOyrTedPa3Glqco7/pQZpECm6CYKM4I9IdLklAb8+viI0YlFkU
fVz1cgh+gBDHHw0agshmgYb8iAKFMhdRQPGSWFIXSoviqQtCq4yP1AS0aNJQkR2w
L+PQboYlTONdpnCfPV9wTxBXzNx1M8pQ2G1VZVe5wSuPmgXGuxeKN1aiEfTX0iae
YiT1BsTcM0yk06bFA0IWEzmsM+eE4Oq0K6ObivHLG9S4CIeKRbYq7q0OaYKn7x05
W7UT7nTurEvu+yHrffKOVNUh8g9XCZ5Vc9IFqx2qUHN7Sln0pcqwQBIqyXKBj004
gx38Sh1B8jMRvvXv8EBJkhfobkWGiZKk1u9ST26vYsW2s52q6r6Qjy83HAUXAjOA
MCHyOHj7uTz4/PvAElhKQYKiZQcc2PRJL7w2I72yxXNW8RXJwMV4X2ll0OwcMHug
H/EQShvProPB4DLPJE7ZWIPkH0yQg21+eSU3Pb2KN1BJm38QSkS6g7o+2Ct5naSz
JlQuzrJZcLJozgCmmH8Wdi33tq+S74AWrwPrKUuFVqObpWA0njyaYYwb55xWiPPV
bguYREs/FuAEopdW1FfIa0QRvAqxFDypCSZPx07d9XgfERhHK/xE6vIP4D2MOoVd
CuvM1ppHyuShttjG3IVGnYCZ4YOYN8464zZTulRO+YFSDywPWsSNVoLdYBRSBa7m
EXAU4U8fig6EbC1fDrcKEWfn9JNFvyAwiE2BICjkevZVBtJAGNDSX07uRbQYXMty
x7xgLiIlcvLsnvUfzCa9tdQrHUfymklrgvpG685sUqdFlGODyZruObPEPVG4PTWM
1c9WP0hZ0cGTU/REF/rXtkeO0WmWnJjDNUAJTWrk+NT9md0NkYh9uzoSEfTiJJd3
aoQ8HV934ytlkgXsNCd5oyb74x6X2gOKvWKNcEBDFeFAYTR4cUVdEDS2kfxJvd+d
+JaKZ5Zdlw4+w50XbgK/SypZrtvatbWUf/tgqGAoRBlhzvKLMRKvveAEAMepuDSO
z5mXJlFzJ4mztYRZvNda+eMsZP9mgXRgRIbayFpUdLLfJUkz3RtXiQOLSdcs87kG
4L6R9ZRr5Y1TwURkAek8Th1yu/o7Eq+Ql75UuLyvR2r8kf7Yxkq0jRUVrpwAOGYt
8cfIr8iUTWp/gnCDoEw/NrH/euZHig+Z+WPl5cTL4zVGL1GQiLKzB4lkRFA3arDP
CyOsZK6aTTwkLVLFx8VW9dN3YYaW0kxxcUf4wsey8HBVpPG6k7CiDV1MHANdP3NS
18/1FoqdLqoCoXs1rDiLa9Xr3gmt/HaR3TheTSguAXhhCctf0dPWifuPkaGEWrzF
wj4nGDHNyj8owR8nbWpigDBGHYJrhanmfCaLDnUVNiV428Jc/XQfbMMnmmbGJXa1
ViptbqPEAvIHOy21yY34iWFbguJOIWKmkYEHqd1yr+bIbCY21OzOMBsLGgUCNNfL
t3pXLobGuOEmyQTebiPb3xVo3eD1ZErgOeXHSIJpXCAwmfyEFLFvFmRcyroUa7Zx
BWB/F3eS32/ILYXQFxNOjfazyqy3+vIxMYdoaS/8ZD3z3TNNtR+s5fzb7MgR/tK9
TzLYeUCSRMleBSZQWZKA6rFVLQyK3nqYeWUDI5c6UdD1FxE+pUJ0zNPYIl63qNFR
0m/iSO7javALFXXwkyoBSQMXGVZuCPA3MXdIzvq1ijJ0luRHRNr+p2M5Y/MYyQ0f
5kdNAy4GON/BhFRBfbLmZvyPWv/xXaWh91xqRi3J8zZWfDo6rGhr/FEtUOVEF/Zr
Ngjt0F8ENrKi/orJ3UJgo8zKG+SR7VbUf8bSZIBKEYJmA5eZDNc6adPnLEvvbnsK
Lj2hrYbwzWj8kCOyg6StAgSvMDQykbMPD+AR69J+o3F9vVJWakt7k6Ja/SKVfHuv
WOAkF2KaqCAfG6FW+MQHNEBB9lh7ISKQ+1yV6C+lzic/hfFVDXn9Dbw+KDKo9txJ
uUhgFgckfsU2obkiBfi1wrA/y/f4z7FakD7sNfc4QHkUTCusBTWTYTR7uGFb8QBO
ig7I1ZJf5u7cC34bRU+r6aZckuT+Wh18LxnsiVM2SXSxrfBS4O9rYLucenu2+KR3
YTQya9gWgibo3n8dwr0tnJTMrpfYuChMP38A0vadX3IpHPRgWPVq6RBuJvN3FzZa
8ueBrOT7MOC5MpAeGqYxwQIGTF+oJoyugjLNmuI1oq4KyzuIuz+52TOHXKIsKFnf
iedkrYkye1sCThsNJj0bA81NKV1S3aC+t0Sv9n2shpcTio9cDOTB1/lq+EjQDia1
u/PKIoPzyXk9/DcTnOrugMT9gwHjKAlOM2KEl9j77MxldOx2gi4lpXIn+rrL9dnC
q3JGBf9482n+0NWBAOUpux0E7is9oT+fExccT4tR8BJQTRddIWqiI4kmuMJYrS77
CQJ8HiBwQvCMgg0H7f/wF3iP+5ug8ePbPegZZwoI68aeOw7StRigKQNvU7kjANlp
Nikw25KHdneeU/fceDmN9vb2BJtpARPJgg1uRy0tik87pn2XKdYrpO6E+Z6HaOG1
pvUjDFZIOuNI88q1+OxV5bT+FbNmHOOdBXSUCpty4+nV9/afyURWFs8XaN4Hoywu
wE6kaSdA3/OHGSLiici+qThz6svp8pkST714ngt4heOKy0o8FhJRrBqyM94Ytkq7
caeoxoislsFOKNSujII2F4bntClUiEpSk/F6xeCzPStHTfcofUjN+Nmz7fRP/8kV
Lq1u8RfCd56+uS4ct6gF76uGuEe0/WpmGqUH0t8ulSoqRZOFp9Kq+QD9YDoo3FDd
aUUAnenwR7Dex1gX4cVZRqDRSELH9fLM82wkoGFpOB9tQRxJdzyXzkSRaGc8LQ2Q
nGTMsDAtCS//o+RGh40tcpdWTpHGNpaI+7PqeLkT87GAT6QmgH7fEd5CeF++EG6T
iuF5mDr74QjjDsrItw6h8rTN3lVVwKZtsrSoIRDH/ycwbus7cqPzTOwQge8/N0ce
MwincMwQQUIrsxCGvsKlao3f4XCEmG0d03sBuKLPzQRx3pVdIrzC9nBgxsNF1BP+
2EgCjcK3uFXlt2vYif4+z+kZmAnQ07tsr+qhxIa0mWF3S1l91bH1GPYAaH5sEdYb
wpQTdt3n1hIrAIMcd4CjzJkMnTU1hs8ObmcY9DMSMsZZMqbcgwGb/6/3uDd23zUW
1+ruD9RT+o3CeeoIRKC3eYKj38sB2GVMQfxLV96nQERUF0+fJS/483+3WBDGoJdN
FH9SOm7PF0JOoqyltKcPBN5oCE8n9S6sshVykDoe3/RoYdfZDKWwTWpablCX9KOF
ANcZdRUM2HoUjuh5s6wSCS2JAFT7veSyOc0YKKu2sQjN43K5nFc9UxKmJueICXzF
rZrXCUMyMqLifFrU/Y9+96ZKUKEFkwPiNWy5TAz09SGqdtFu4+MYyWiQD8mtzZ0P
QLNPRtPg0gGIzEgZWsXqMgPcOIZhO1Zreyl5QG4aWJykGzrHQzUD61t1QOe6Y1yM
2l0YSou0E5JaZIbaThaQsS6HAr0lt5bbxhIze+/NG/wkUXsWTf5btGU8aRifYB8Y
VGuk6UfOUTkw/bR9Iutbcf2qaUS7XTCkm0Y/wrEiuXiTSXKRQpKWpckuzJfSkGlC
y5vNilqBzyIBsAC7h302kc+uapxfEL5WLW//YFUAWne8lBPuT/r21ZgTk5M3yByc
LZy/PttXFwsJojKm8lA/M5plxgcKp8ihJwiRxOOP6rV6fsTtM0VcAotM4f1v7WR6
/WqhBwlTNfc52UA6PbOC/dn89Dd+7QALdkO/3RVUyNKcflV1iA366+NBHbel87lc
N8wYPwUFKkZc6CT2jW21o5ZQi69HYqmUhzzPoAklin/s7LYK6WJSJIcboJ5ceLqU
GJvutKNd7RHJ+2+jet8yffiEv5JwSxOv5nFZDsgzbCj4mneIQ3F/y2+oXrZ8sfzZ
guEXk0hv2uTECg2f7BgmVTGtz6FMCHQEeHMkBJTbaWotgnFa3N+ekNmO3x5GKsr9
vhnWzzN8YPEZo5BZbY9ZPdfwUxCqZxRHl70nwdI4xeTMm76g8dxgWuDpx4yNu0hu
5ug6BY2eEHT0zrikqaT2LcUQcuvlURQjGI5jVcBgM33mVEgStT7nOH0qzxMCFUu7
LtjXekbM4ooxTSJTgOzTfUggAkZ6SzRvZMhDbgQOfPIutjFSLtXAt8ivQ+Qeg1Ad
EsYg3P7DYIarTyvxIoQ+zr6pgptzZWLVH72yjkmVCYsKQSVG0NuYX+JKA4Hcatvl
f7phgYbq8HynNKNuT7MY78+sInyVq5BfEFV7uHmIWtrT+qT9iYl3wWo/Q/JZFPxB
oH+VhH+EUSOxqzRSe/qU17aCsNsZKzaae+frL6mnzAEVVBo/hDFhdzCj2JmzbHLq
HUhoVPEYVBfUh4an4LgshDmHL0f45p3ymhsKYSjYp4RMrI3TsOHYgOH6SQNI3REi
s5sLUr5K5w78rMVzECjPnCFujKTcWQjsB198BHRX4T2lU2z4ESh3N3KxeJitpF2R
N8D51NiUZpi0lSuKcusft68YRgtXtJwMlPfg6mpRtX9lzoHLnICX8QfKuP5LI/kl
cSukKMeMERLouLiRqJU44696/Gias/AHYKcDqNHelxoSO+XhyeWhwSTzuHtQ+9uJ
B5GMx83pFjWbnW19z9Qlse+HJYD9iShmhM0IgIQNYEFl/X3SbJT69H2YGVMf+Jca
zlZppdJ644GuPmUxfBKBM7e26yvbmaX9KRPDBq8dNb7lM3hYhgZH1OFH0LyNXSGv
uIbqW4QmD10oYo5dnhYe3sdRMF68epP4pDRqgdvdHpBaMBMQaMqKGJteFPfxnia3
XglrM7MGPC7a21jVKWQR3v2m4HgJm3zzUOcPmf32S3V9Zi/ZRuqo+m4xqvkBTnil
7Hqwl7aPXWiOp81bo294D71gFATOXV8S2Kjc6qYmF91E0WXKEuC/Sif7KXBldnJm
29iAZgYmDw8UsDKbL/B44wcVHmlFbXgjSD+VnONxamgf8CiTNfq4WJfBhw2OkB9L
jmHQ1hIPDp7YzU4+WMrQiET866MgrSCz60zGac5Wv6iU9U/R3ngqZWLgvfrJyYZb
BpUOsUfNYrCF9WZBhghHMbIeNplbA8uikFLc7o849KkHPmXHRLyUP4+g3kPGBCFW
YTC71b2N914IO0d/ZD46Xr+hYD4yDMqiRVLgDH9ch2d71bMci1xWoyicsNK1oNZC
JT3w2kX45c3j3cgLQ8rs+8E8a/qRUsFBdL5nW0GRTsJWw85g1RfzlguMjTYoQngO
GMNHsmoe7UbkrV1izYRmCSZiGvG0zEefbPjQQkLf/w/Q7ABy4ldPVvw0ad3/SF7v
zcz+OKqCHPb66U06vCxgDa10dO3llafxHuhLCU7qxdwJ0DUmP9TZM+MXDrjBnmU/
A9lkKkq1rWUbc376FC1WpcoH55nxMLyYRBAGeBCTCvyxSuM9V67zcv+VXML74g0t
b/EOM654Wm9fZ3OIUrv385txc9NNV8wE54T36YpZ3CZjTObyr8qIJwmO44vXgZjU
Tm/uuSsC01aILDnSFnOWpr+PLb3eiGbGmw6YFgWLb4SxeXQpwvYtWH9ANpV8y+CD
YHr8E9pc4xuVaG7s5hnSwDcyTGkTrxm6Mgx8oHPhZSNJGHD5f4khhMCZFZc5eb1u
QycYbtwO6yvdH+rgvt6RznLy9+QDZ8mcHQTunizCdrRaVQYzpDMeB1XMcW39FiLu
PHdr0zgdI7neOA6rSPXK9TmIo7ZLA4O+aTOPayqIAJ8viH2Q+iJ4HYS9RwYMoL//
VONGSGtAyumGZtEWnt837wDf7qlo0nBc9Uv+iCTUNM7qzIlH60UfGzI89eKCZBni
Y7/7saq8fFuPYjKIaJavT8QhIM5LOqU8tkwqodeLFG5l6RzN161pzjXBsTFmpDEA
UNQar88bCXPLOlIgbQFsN8G0L/YSfHWkgcbcJmjwhY29yGGrsodJVgkmpzjfVbcx
ZTIs8PNpKxWk7YafZrnFw+cA0RUMJH/ne4xcpGsTjd1BJu0x2ynjXBs+TWuO4i2n
l36rIIH3BKMIa/Kxsf/lPZs4/I65MQeLDRDfIjWCv7Wdc/7DHcLNovvsx7O9AX2B
iw0H3RKxyWg16/8Wt2fKNuwEe3Cml5naUECx5R+WGQFLZFJVGJo3cGOSEGI6AD4B
VALIyyev1ZwDot4TJ2XjDB4vSQj9WJ0TfxuBXVCw/PM+T0HJ5Orea2mMKw6iAFOm
obM0FQ2RwEhuVpcGcNFuIj++8nawKJWA76fXpSy9YZ2RaYuYB6yBGSUSoFAEK6pH
1BMRcL0G5GjaYYPmIlrdkSZPmwHxWueUN5BO8MDH4TGpCDUpU2e8fDFK1Tdb/9mm
mC1r+HxBVRCYk8JQQ0LqC5iZK0E/NO/dFlx7hIRiHkzNXNZZuVA5tywKF9y9vZxe
dloGuWeeP25J4YzTKRP45xMP8o7bCL4xi8sEmqn3CPPeAEed81egR5uNTMnWlHP/
WCReZCGoN/5CCmtZnCHqohWVfDz2gxGN8lvyThRNrOrCarUaNsxHaoAqXnhP44WX
gX8hDBLES3NJF1bhIZruvNb3MtuuhfYxAsLJew1DMV/eckwTa65OnUEMpjp/lgxN
1IhYJxfhHa63+oGQ2pLDqcfiZwBvQFenBM1EFeTkmTJ136gBxhvV9jfp9SF8N1yM
ZcjqYe2QvRB2stHcdlACJSkDdPVZH1kQ/48OvqYEGheEpWnyAOR9cs2H3gVRnY1X
W7cIsK+qjIyyJTj36ii645YVOXsESZ6C7+zoLl1ujINgil5NrxbwqHqnublBqGWP
cqQDkLbQWNHnoD+Zac474hERF31ioBNr2PAhoHUFqU/TO326JmBhZUNzZ0gegiq+
H/5rG29Td6wf8r0ANrMFQGv+G9/gzaw8Zxr0LYjBrKYxJJhpXV4ZmIrsgt9WRd2o
cDE5Wxp1a7pmdDZKzW9r6dms6E5+0eNecYk0HTztlkm5CwGPtci/494i+qU/TH20
kGqZ01/YWqDMkpEhk0NgUNH38UBUxZLXJp93ULyvibpaHZJf04sK5fxwoeNzImwh
Ry7H1DpmrgmekQpQZcoFbm9Bk4gEZ3WuOQUDMupAfjBQ6+1T7SVgsdIHkzy8BV+M
oql5lr+Nk29J+ZZr6g7HnaNUs6oo+TalCTI0Hk+ZAIT0iXBGweFcjJ7i/6kKLQf9
nb0J6d9cD/Cm845k1wjecZobYo5OlLdx06fxJHatNRRlCBEGm8S0aX8xg5MPMpOl
83fJsOAMH62PJQ9DapWsjlLdO/poMbjSwh6qFfttst+/NTyHXti7WtPDH1X02aKS
0nV1vjqMWli8MUpdioM+KQcBt05woi9giVU5JTHPTywFm7Ez9Rh1jrECuA8X+hL3
+lAN9CIZ/GFfs9CgmF/esxJJaUI3GZ2WDkXF5zNpgehNU84MLTqGP0SdlmUqGLmK
NgHbvZGzmsAHqxnzqxF7oBKhISXe8PPeRRhExXVKfa6Ejgvr/HaXLohSOAiVvkqB
1DGxgZXCjeYc+GHR/NZp6fyi19/wXRpoPzaxj3e1If0D6BpczbrKNxN6VdHaVC+n
xyLpPGHc4J2Tx1Fr3cXn/0hppvCcRE1eZxeDSbOwzS1W/OG7qDKE7f2X5DL6mfWu
+A147+PYMhET0kS2OF69i7Rxy/30Iy97j06uMuYkpTqM3aimTKw/TAmkjLxhR+vE
yBVpH/Q4cTNJW5xXy8YUc75pdn3bmoUwN83PyH/jAUuSGdcLBacbMJ5m/4HotMkA
H7IfOFdc41hgScJyLc1zSuczd0M+of6quEiOvgeoyDtoKAqvkzIFbawC8tXSQGCj
lpHr+uhxAqav3mbOyd3GAoB/SOc6ol2tdWUriZ5UCI1NJOsd0LzEqFbJbz406vQ8
8/kvLsN6BBzqodlqkcHa6jSOyOa5bUKFRsjv0Q2G69yG13Gif0nF2ImFgsyt5y48
mVvgpQuWp2HSS/I7KwlUk9nHjOVZcxUF4dKw/kYaYqMgrDJ5fyF7nnfDMzRLthyW
A2WxW6D0gst+c3r0YjFqAtM4MIdj1iF8FkPXwVvsRx1Fy6iXXXanO0/09lw0/q6s
kFPdRL0oZRs2A0TPKW/gHDrAYshzqzREojSdGmsMQ+JHb3LU63NUfpvfsXzThY9T
/LN7uNNiPlcsaKHV5UIraLY80wL8/BVU7VF5AOBmLkFgy3LWtv5BTZuRA/tp1f5d
fTjZmwvYP0K3j5WZWbO/q444ukzQ6Ugd9e9+2nImc5hqpJOMqu6SuYrpBQznCFut
MKn693Y+Nebja91pUsoql1fite5/rxa7vgtpf2WXH570yFExgzbokBdlYMiWGuyZ
+gKQ3SvGtwWwtFoRYICDy0gpeJuYO5gb/+cm7TByy6j9YWRWg0JnXApbjPLvZnMy
oPWIuACbHTx0BVm/Ii5+e+D6zCs7HODb2B8PDlhs+PD7uy5xUbcgC2Q6VUWfj9hb
Duy3kQUkbtQ4wU64+VMqEi1O5hs3DumPSRWEzNV/3ZR3hR/xjFlKQWmRYjzSa2sQ
86M7v/HwIVhbV7dldNB4bgilFV+tTaUTGm4CnMwv1+8U5ESH9ragVX4j43GFkA1Z
c/b84OJIaBJIi71hHDzgmh75hCcVwTSjXPG+kARlFdoeFdwnKvEFynN4+W/pjs+L
buL1zVPMzMWlHqgSSaavVzoeNqbvdqOceeF4yX4HVETx7eA5GMOeJKZmqCrAIXaI
fA+ha1fGqpFCLFXOwaNSDh3H3UAGls05OaZ3bQiKRHFPH9XSbdKJXlTwabMYPOzE
DHo3yA/z6VUlR2kBBlmCh9M9Ue5LLjoaPrHwWLm0O33NemPxe46V41u5jfxjkrUf
dBSCY4HUiptFRs470A+9T6TsvUbDZOvI1Tgngo79qxnMYWq7n2VoANDgufITcn8G
SLWROJTdyrCZA9E/KGleayIQII9qAC6t4us7sYEGKSbdXRBpijyZ8kyPlO4ceCd7
+TyNWVn9LXKTanD28mMh56zwRXJ+nb+rugf9aF/i3+nqqL7QTSmSKhyubHOyY31V
ku1aLWbB9/tk3UJBriDYCrU61wTRSFQyPjkQdhqYZ/3Ejm3RwKqtKda9GZfzDa2Q
hUhPWAo3J9VHwZSHkJGDFPBYABBrBPiqDXi1J+M3/4I8BXFnvo5UrXqOnpM0LuWF
KpL6Pzi2sbC+y1Zi3FU1zBcEJS9xS7xIp+VY2ePySZWEsdl5Ly2eXTXNw7pYFXtl
BWIQoFEResbWnqZi6PoF0F5t4VOE6XeTkX+QwUbGORXrI2Vi+1TMSjqKPiXeMZ7j
bc3GVw4LwVWJCEI3ZcH22oCU9q6354cdN+TV69SWNwrjeCMflWOja4eMFxHFNi+l
FE7dZDfWuI3mca/OrJqyqZs5e0uzCBTAkeYoR9XVcpK5TQD9gFcr1e08rYlDfoxD
5E4nYyIhKk23BJX5GgGcs08wYvdz513me7tzw9Co6seiX76TIwrNr7wO7gWudEPX
kTga+VnoHqzupDr+FLtOZRPJgSg7pPBId63dlulceOP3q5GS3CgIQhe0pyOMT9Vv
lth5YChQh/3zYp5mpMug9bvA3EqJp6C5y5qD7Tqa5QXA9qrCGa4iIS+VoIE92hZc
/Ja0nK/TUSITL0ZdZSTgHn3DWjSpJmXt0cyCDK04t+asK3non7jHQDiU362YVzES
mIqlgVj6b4SD7kS4K330FcL/ZGJH88lVjfM69ejQ7F2u6BtfGWmqCdP9EpFmE8Ns
3r8Hpq9NnR864XoKhkPXcDWo08aEa/q1kvGWOXi5ZsDZlZw6Yrs9eh3q5HGmEWsh
QIQpLGVYbNtYj50YmZZchOLtn6zFqEDMOgUizmozG+sHmn3rWpg5Rb0SKxZ3qUgE
ZbSztl3MKG9SCqPbLLCCtLBMJhi138vPKwx5UAHIJOQ2kCgxm0qkOU5SwvF+CQU1
ADoSxXlysx5ToM8s9x0+NWyS0QRS9EGKs+pKgLsTXwn6tQX5EVCuMnJ8u3xzPms+
bd6lDdJtMBgkyL42lUrIDcI8pN9iPMUxXdOmeNYqRUcWSdsK9wItgv7T768tDYGD
IWwD2pggz+YM+AtO8RKCostnyzWKlsORXvngIp0P5emmrYHCfwbmWcPf8roTE1fQ
FlxNAd0qPqvIVJn9nJrBcHWWcfsVpdhVFfa+LrF8dPW3yLcFMvt5HA8qn6IlOXWZ
XqNUxM/fk7J8P2CYgmmKwi/+JOciMAhoyZQpU4LHmIQDyTYfE3IkyreCzv3Fwumc
XcHchf6AB24GwwO7g4dYgsHhKKr0eArUQiaPt7oQ9f7uB756IgeTWujyatfThtuo
VOZWwlxC1a9jnW2DARH/7Y3hWRmG1bbMfNLZOXpzZtGLwCYNHGQbuFoOprkwmDGI
I6ASdUBtBUBxg0dwP24jT5Rym79t+u4EpSxqMv2po1JCauNMQ2kHmUMBQ7gU1sgl
GZURvnuCWfbcpVEK2T8rMs6wAaF9N+cwFAIYqyC3cSqySjzmIo+fEisiNQlhjZzk
pgpfEf2QIzB+klKu3WZHVlwZ/PKQX7e645OB4xCgyVo9EOz1WKxW0x6UC+t7uVro
nDxOaSC1a7/2ta2GAbQYm6dYL0pQAHEiX+EYQn0tsNOZRkvI3P0pAYwKg/oVq2VW
zkhQNr5UdM859M358LN4+GKQwu4+jyXcKr3DZIhi4eJvZYynrxKiaDJa92V4NrFQ
/il8IKbPItnisZ7phIsGcg63CeRkeYEntOKMOog3Zuv7TZYYedBqqTNpzH5OvAcB
3aFkw3OrK56xLlyzQulrwookQR80EeMT5Zj/Q/CPpw5K8vSnxTjtHRBSmosJEknP
ahqmCCoBvyq9nWQtNkYAx1W7Ei72A7e7UVmKqvBqxY+fNegYMUmAZMK5ouvv4U3d
WruwYWYsNzC8GeH3AJ3RdbbbLjwNE0dZfBZfzx9I2lwyJtJiP2VWXHcR+ByObj99
qkr5vKEYFPYbQoZKLVRYWtDAE7UGHRvy9Zdb0OV/e5wkfEV0NKPQWc1a+dO+u1uf
+1imbtW0sVa9M1i6cFwq5IyIQxIoigVi4o1j4i2FIbahstpto9fYpa77vjJd+1Sz
sXKD70s60WO9AAbwSwiksyNGdQ+C6niqtD5hbIJ0U3pMOpGQFALrngS1ySWfKPhT
net637kic8bYJK7WkilV13idyi3/jMt/bLa9uM/SY03fUXrFuy06/UrpdskBt5vF
R3qLTaQfJFmxcRZEIwE9nUnWJtXY6IEMSsZetidcDSDwTDwC358oTsbv+ziknMyA
cS8Bbzzg1I+qbU81PL7NuJO9HZ+rqFBVc/gjjSIeyvoG3Ud/LSH0eebtRuYPhQSD
Z0NmxdQ7yEq441t25eOgVi/cvPYTk9oXGhTQWBgnRJFgZMO5Nmlh3EaYQIRn2K4U
EeOMmPPLwQR6JdgAQyPvfrEJ5NLYr9afaUemq12pFrwjOkFHBup2MPyiUKCq+E2M
GX6aqW6c3i5yy9ANBSUD2Hx64HtT+3r23UPufK1stV/3ztB8YCVBjH21dEYXOQKR
YkjjGe+m6JkJhre0TcXDtRRoGArMiMUBFYB/wEeiEcIyha11hVBRkGWuNJExtiW9
vYa32mK5u/1xGUA8vKcgpUI4iR+Iu/r1Tecg8Y8rNTjpbg4A2MWD7mX9Wh6dpZgV
vTeTS3XVA6toCH/Uvxo3sngzkYE7DmSYsK/dbYvIwI/D+BjNBUlr5ddOqms9WqpL
4ScFGcEVrvQy9KItTtv3YjKKZPo/48zxFDuTDK38MjQqhVf5HAVa6FgP7RcdENQO
ZkophyGwLamRBakPo6sh+D2gcT648T0NicHeYhAXm0ZyEff8Z6rFdYXwir5NT5MM
LdTBaHWc51yA2kbV0gKOCpTYCP7d/gaqhpIMbz3QwmSSxxJ3SCzpiYPDQbQz5IeL
IX8LOMnK0PJRzO3PRoWt0t7rhnsVcKVn0B//jZEPwp+nl3P0fR58Y05GO0qUNp2B
1bAtUgipxn7bE2OgvfWKHJcGWGVI6yzt1/oKoD2xtb1yR2/vC9Kyr8g1o8087zyZ
P8AqEZSK93ytKiiPsqOF4FgPDpevqhRezEJYK6ai5jdpU5KzFJEfaRVyowAPUq3q
UkE+mYwXfo29nyBnQyzpCfp2d5cCSAWOowB8i1zAwlSMmfbSr4zC9kKais8apJgV
+7uoHrhhsvX/8NHWkuv3Ts63JZC9pgKL5We9ymLO5I37J+XKOwiKYroZnfMM4nBC
39UC4ipIlRx4FlVrIknfIGtwSmkPMDDX3sDRrKfyc2Ys8BhbmL6i/isaV1vWReeX
kv9GaxgIySNpFn+2YvGzJLSGinl66lozfOvAn72ItWGRfCuXteOg6x2NQE7heQpL
RmI3aKKffpOXI1pwgVRrskFbzldi/R4VYyeEoylYuDi4sc7mOs9XAVf/YZ7SdsNc
CPf+gWV+wPmJ2o4VbLYXRAXzIxaOJeuWnJcmTdC7gXXoStN7cwTWTMKAWOjyVI08
ek2zxM8/y9bzqOs/oBHb5lBZvR6mKwKhlh+0i6HzkBSpU17It9ITsShw8CpSvuWj
4nNt0IjFGovPEymlst834hDqNcW2EPjV1FvQunR1NA57VIw60LIHRsd+Q1adeQLR
l1O32ND2kl/WmWCApytzfM4r5B2SVJO5gxSwQ/az7mqofRo9ttNf2SeOmKDrM4hz
N4+Pdurk5jo0/oNlKyLAcscwsys4YEzNhUA1njAMp9tTqKdiRHL+FyXKFCUAeMlf
rRBB+xNrF6qDE74c6wzJ9MaNW1uaqbbE45rfLlRIu2Bw58d/WL0swYx8YMiY1yH7
g+Nv2FtzuLr/X3Bm5B76xX4aU4lTpSw7fYjrWAu4w27PTozwEItQoNkIUmEIIhTl
2myagmBbF+WAXVuSIAcoztbQ8/o+J1RtyfXda95DvyPIX+LkjYEIsDOdr2iOGFXF
ln+qNCjj5YMtyPrLQmgaJgLtO8ROLcxFk67Xq64B4butohDqR0OxOjtmQCTBWxsw
er6h1B98zlDtfUqEkcjVb4LiIiJiZKCc4BdgdFQZTV19JiQnCEgArhw9NZ0RwEfr
vYNscinPkoFFEtQv10EzTuCIdB6dhKeKFuDLN4k+zBR50kly2dDeXIwLqHkZOddZ
x0gbWJhXBnnfSkTLKbZAVY/RMR3uw9Qe77dUCEXe7cU1bPa3HTFDLuTEhOZ9fQU9
qcC5EKhGjCD1E5S1WS5I9Wf+ChBRrt0SUdu0A8+n+8vCxFMArtjixC7ZyD+r0DkX
HSKiSzxKkN+GoJj53Q20HQI12b3BowUasAICRzhKCQLa5gUsq7xzu+KTIL7amHaC
jKdIOAh6rUuKLtpTujJXNXiD7+STfMOzjSnnbHjlCLhe9z9ZUquGm/3Avpd8GROq
1jrBJ2zVhFJdbcQYmeN7K0yhFGwY9UXu8IZMP88PvTqpIIderxVhERDO1sYS316X
FmB8P+LYwKSEBcCXgU0b5yYqY/8Akyvw3l+WvERW6PUXqp49f5F2mwqK1Tx5ZKc0
xOa11NIbjF9VVMvgQFe7/qOs4vR/FX67TT+lYior3kWO3gsUahT37MD5dzFFfroW
zjZTTfC5KocRLMfs7bxZP0IXjpWNIY3aWK5N0HdIlUSGvMX7lpeYsejAA9MJ2WMn
WKLaKqkYX3OHGUv0ki6Rmpthc6SfGm+lr5laOgViRFzL2xEUb41Dpd05ujmzmX+t
q9igPbrqIgy6m3dNFtpmn8P46sbdni5vKlhXyevdn9zdZtBFCGU/inxxNQZnXKwl
62tcUa4LZC6Gq8z9STl7IGYzAI74gIc3vAnF4SluIAlZKxDufltzAEAXty5ErTbD
fDoFvGUAR2R/7CzEOrjEJqQqUvbCJP8hQJW5qpfz7bATxolIXHbTCZIRnhXhj0Oq
u+/BTslezyg+gdmNjK2zKd6xL8pElu2V2mQjpumWShI8qCebL+jv4YvBGMG9jw7x
fvHLPR/xx5sO5ANJTWbTFM7e28gpzjctyQlIzMBDeRaybazHDD+zni04FVJWfhQy
wDe+luxH31B2RxgaDKzFpO8hO72ddsMQgFfzhngK66V4sKOHO/ckmoagDbCiTUDy
ldBx55r6C+HZxFEiDHqTir0c38LLrnfLsLwsBmuWNLd8pf+kO5LyBe/jkFuCzlsL
/ET3fiFL+Z3eVOeNReDIUfzI345JvvInh6eu1UFoxLsHpUr60hkqtfaDKPxJ4Fwh
0+whkdm5Qxky+aztycrp7/qPNItrItV1xgxfRKdtTanu5vcPFh3tXO6tLYYhfqMD
jD3ln/pu2PecUolqlNNBc1rLsekvIiS6redWKOn+10Gw3vKXFmr22xFdeoOygZHB
kf+BKmYAY7/mZhwJCrDZhxl/kic04O2rjlM1NFDgJ9XkCY2km42E+iEtfIsmL8Dz
7eLzI4DWDL3xwtVt57wwCxemlYxdWCHGwF2rIWTjtcCQ/q8HeMO9+dm1xRWaagy+
CBD4A33JiuDQB0lA0wfh0IfNyDSKF8nHINDMN18iUj8WvHR3yKQQUtsXwNYMlr/j
rZJCe/QQ5haEtScylWVePS1HU1hq6nGh2qSD3uBCrBnZJ8bspz+acvjf8B6u6CIq
PAXq1ttkvvAQVMc8Cndik5JVctNTMo8jskShbubvxAmAoqPj6ZKbaxoHwKbCUNZG
x1G0lbbJD0LyHNnRrCGtKk/Vs+wwcvbsDDblharb1Dw+bTJwoi+pLHGoCOvBWaum
A3icUfIYNjusPsO87aHi1PLNHZvReL8bUZ4JmScdicfkQ6c9Ourk6dFrdD11e/aN
JoukijGWpQb6zOH/OdMDOiW4VCdO7pOjM/oyc5qr6axxaZenNO+GUamk6r01SJkL
Lg1SwaSuGapJsRWEXhODAtf3XAnvSKFkZrtJnpyNs6r7OOZ40QK9hhc+hlEZ29hu
w6yCHouPIP8a6T8pXfNUSuSreGFTCR0NM6VZtBXaCmPNB1gkgLXwNGGTKcMJMPFb
dS/2Dca9wJSjfWSi4LjUSNrf10fjaWOYNaSFLqfW06IP5swJS8gXYFOfG3Wt/VyA
OyLgL6B15Q0BVpECOcpvSejbcqMVnUTwwhSZ7g/8q+6o/kWzRVmfXm3hT7yVyj3l
H30yAR+c8Kvx8/yqU3XaYMih2gUWhHriW31940kwF3mC4KejIn9DW0eWgAwT6mL8
DCtKmQNSmmFoNfG7crE2P14VMPi+CRj5lYpnqCQDR69MeZM3b+8XK+bDLcutThGo
scWq/LJnRsfSUW1wH8Kee/xW8qHiTmINDjtd5rpU5ApmjN8BtPPmF43xJ0fEL3dq
bjr10Jflos2UI4LCmE1XW+gduPOxT4hl2uAZPjsGRUlduppAyzJP7FAJqBnueK1W
7NySlSE/J7SyGnaiCmA5HSdFveoJpSRBdskE+QOJUYxWEY8aHPAFPHI7JoBejlbK
k5RLhu0WrOpZ6ivy/NzpCdwoXVWE2E4XrV4DKC+Mr8WrW388ZSUolXsoBXgQdtNI
MdM1w20MuH7Na8cjewcmTMGdbDEpPHYPm/n76seCTguSZHUJvdaRHhonHdjoT6xb
LGTyDPF1A1SToFnSOEfHcGRbejPZE6ppq80qe0Zc9Ha7XEOyrCKYecrvoBbamlmH
N8ogB4MoyWmXLovmbEXjbdZvc7Dc+zmTaofnsDhB7hgxaNqeQ4Qx+R5rStuKfSLs
8xOVue6nKZRBryCpBRk2oqbTyOPPZHB1yrLDFnpEa0/dgDkz+aTK0x7CN/XiWUzP
CZ37uqYrCwZHd57nhZxFFvduPB9GgOlrMC4ynccwRdvIgfhUlq/QyuZTICl3REL+
lr8w/9r5tvfLjfjh/rpKBr9hQMpAhMmzUCeei67aWWb0H7iMaim1b83/Nlq1gOLH
QDQFwZMqCIfPAgaHaSZUt5zXHcvkTMu1fCoxyhxNHQFrcHa27g3UoU2fsEO4toH0
9yo/m8OchJ8CsKo6w7V+c0gkfA/S/DQzsOtpmkNTMRNlMEkdZRaUV6iDh+se7mkK
tQvtBuoEThFiGsLkSu2VEBwRqFrHBX58H97DQ2ECTb6Rz0oxRY/RPHdAts+m6Eok
bcsrgkfZCpPZjTksRZqAMCRHyjQdwFY6gpp3JDznyFGQqtgHcKBpuBrg93hTUkQV
vUvFvErO0UTkrOpSFKte9P8gPSRW3yFsq4cJ+qcdOT7VhhFmsp1AY3ESls8UD6kf
+PD6ZdD36hKeKYQiLoHl3cqpUCWmnWTpDgUq5BznS/ILieGV3dPF0LA06vHLrd2U
83dmM6L8a5ZodaipDLGpMBxSid8rnri0Tcdo60R91RTUVAzE/NOTZUBrLVTi6NwB
g/tr3xpi2DBRe42DrIq1gq34joIAXPVfo0ayOBwr72z8gZp3tQxNEK6aAGvlW8AC
A+3oPnPBeOru5Q4VP4Zitfnz6hLUvfUsh88u8QcOxPGLvjDiZF8Tuz6S65Mw58jN
vFrmhIh+aGEi55LV9mVRHvTXje/GHqBwXMeduGyIXDtDtNAJDv9Y90f1t7wX+YE4
btbHM7MQt0PjwoU9/QuUJaOZtttv2QZlNZZIkGq2Ex9dxwo7qsd9ROePCdVQyyR4
SHpogEjl9bcvFJIIEg01boZ1orwF4vyY8c5jH+sse7Sy/0WItgKcgbI8Cs9xbZF2
YMJIb/b2ckMbILz8wIjzReeNlLi+iapV5cM8SiSGu3HaIEs1boPCB5A4dVEuYDei
i5Yj3yVmslxpdUdBMvvMjazoISoNnTsMfLSC1laIustqCwk6SBKFdPIFUjI9kM9l
j8Sg34vgllPvDmQSTiniG07Odbylr8r+8GqTu3dU3u2WyKKV2HuoB0dJIfn+Bs5r
uOafj1WCvpIe5qNSb/XLrQs94MZJfWSF3DqJVhupIergbm7X77/RdrHg8neiyh5v
aZhYOSP5RVFbaIFYqLR2czcEGb4jWPZiFAu0OE4SzdwNdEnC0jPKoeiJwX1GjCLP
glgoUjgSf372+gGwQFNT0Nv/OD7XmWkYjIonGkZU2gT/l06mWKJATNf/XeAGIrMS
gJ8ACCOpsvBkPkShHVQfJUckFv2yKbiZ26irpMZ3TnxadlJ5pUIo/6pBga/mhDcV
Gwh+z/al/7Tani9MUZJRWMy9iwly28S7K/KgtGblASbzRGpBZk4yIjznPvoFt5/H
5O1p3/yER/JmghPx9e4s3a5BBi1t50KVWMcvw3CLhNswuJihC4aOH/TEVA4QMJHt
jP6oawMpTiqgWPpW5q/GYDknmGcWDMKQ+K7nGUXF+4hygnLs70+9BBvJpdAu1Ig3
xCr4hbaqVg940bTFf8TRAYBgvGK7nfC6TTPKQ37G1ErpBVdN2BY0rXE5C07u8GWj
hPBeuyXi4LXLN4SekK7CMdu7oeVT6k6t5l5wffWKd1u3nleFE5Q/6bPAk+qyp2KZ
H3WRots15KPm8/J1yAIupgGojUKoLZU/l9bapjdNi5ym8GV942oAzdKxpLCslRTi
tIpFzm+wYSBJtdPrbomciGLhSduIPqruilrTVFWm2CKkvCxNZSSe6CogoQoIuFnR
iLN0qbzwQFUddg4CsKI4AzyRYJTYV9I19wkRoP4Ukyh9EqGRDQjNOwDRZKHcLi+5
U96mqIguOAb+k3XJY6C/7yF4iq5TooBj0ZZ5zGilweumsKkaiEqjxNy5nrf+dUel
jKYT1cC06SXOrdXdZlDukOD4gWIf5xgnc3Bcxi2BRfsrr+UDtOZ46WXJH9evRfDR
gmrq9zO2o2df30yQ/TZoyg7ONLGKBpP3Lo1enpL9HAxjrvvejUiAqqgxTfThiAny
hvJOK13PKg9F7AcGVOTdcc9zCD8EBn+PvSOOXmwOOCo3JAJjkr0dnSiFUR5G5Sl+
QY4NktD6sALRLLZlpSbtXUIKQoq3stRnINhjEo+QPDYCo7GuHxdE9/fUR0PbTlh6
0Fj1HqwmYB6NKNjcTqwmk5DI47HBEY8vDUvJrZ+YSx2WJgg+b4/xYQta6kQevItG
y854wPsVeu4RaFVGj7poIB4x5TUPOMj4Yd4EgtD5L6BeRQhXzkwi/vpt8W7VyLOG
3tPeKiHCjTldyygTTt9LTOIZ0CouIjWRgYQqRAGFxapaZS6ugd+j6xroaTIpV4Ot
G4TigNB9n7v4MOumurM+fJNEc4x+03P5WdwOKPjqfQPj7XJkcZYLKVv458RAeZr+
GRM3foucbYg4bBmXQF/uUA+cUT7HFjfhtVq5lzgEjeM84fSqGMSE2BPpGiLFbsvZ
YNwiKOIxpg8L0b4uE4MwH4JzzvA4LNVa8p+F7qeo6t5XIf+j23vJVRhA+74dyJDC
RWwBb4gIRpCKKSZ/ND4V1sBTa/XgCBk4ev4PpiYZ+f4nBLkwWdCfaP3fX4pzuXgh
tZKcUewPXd4xQRoRQuY9v38ydR3K0XYwDTTM5IJLhWmfKa4r6/hl/2Mpd49EE08z
V0RhqEz1T3bwJPdVc5bfQJ+0cHVZA8Ffblt1kxAhaEW8oQUcvsf9jUxMFLDa8IdY
4AiL7rVD3ABSVL3yP0ReLJw4X56UiqNb0iV5/e77VR7t7oxdnO1eoB0RRdjhTXS0
edQIyYGAanKNQzAmp0jF0rw8KvT3LFaO8eMLl9POUnR/PHVY+Q7SKGoj7acjfhP3
cvRRfHE/SfqbZFbS3qJoBvt+iVJ33Q61H/rHfWUToFdbzEVmM4V/WdJ4SJtnVzSP
mbibfn4OvLazdHx55Wo/iVsoZomrIGlq64+L/DtUk87VvCzxK43oXXxACVpqn+qk
xN3iqPPjJq/2wy4FZnGwabgj149bnWSPXy/URf6C5k7SnrSTgSgR/9v9J8MxD/Ls
xgjP1xioRvU+I6DA3661BGrep0I9w9Tfg+LhE95eqvUKAqtik0/lbewJXmIAz+9V
Kd1XOnZos3jvkS/tDM+di17DeUegPwrGGy8XQWb7MIljB0npn+adthEx+bq1OKxj
mrpZVLODfbZBKgptdjRPH5PeUV2c45qpguZtS3ba/OkLLWrb8ycDjW/Z2f3/DaAb
IEd3wurpIIgmQ1v5PEm/DvfONxgb93vh1ie+Gs71X7Zss+t17M0ATeDZbqW37+5G
Fn7TENSDyUX5Sk/jl7ChrO8iGr2esYR+TwAbi7p9QnTPxZ/Quj8j61ZOMnNztrb9
y1CinGCj9+arn6Qg65UP+Z4E0KBk5fU6O8jTHc/LUqINdGCM3kvUbGM9SD6jlF8O
3GSRXfiW36e1thQKCWl6zvPhvy+96m9FytJnNRp8TqaWFArnlT1OTXWrQmlnaDgR
o48dl5n6D03G1K8HZ+MWE8Nj/goI6SP0+yJH6SWjkp/Z3YYtFWIlY/W1ZHSK9UvO
WgEFueRSHSvJ6vKlT/ezBCirDtLwtiYeSXnk/kl9mFRGog1Lw80Vuv2V3mZLLa+J
euBK4/+Nbv7v0B15PYzcpz3dY9wFVJrMVuxY4cjOUBcy8EDdqQgqqTHNIT1q0ZMB
l5P6n9HaKTONa9Bl+C9ncOvnQrJ4dY6mo6WuBPSTG3QAplFQnoyNESGo5JGjwf+a
lRa1ExCeTjuWk2SiBICPOuMNzc8vxrIvtmSrYRdCUmivnf3yJa3z7hEF7CvXQXFg
xfcUsdMIITpdljYKuNANFWpJ+jDMrSBXgYi+2srZ5sQfWbh/LsgwUZqKiopZ8IRt
DWUedQZ0X0upJIhIzYtQhEAJ1Tz8f1J5BPe+fkxqMhoTE27Be+aDYB7MvMY0A+Pz
8fQ1PjUKjj7BNofMevvQ0SyCz+aA0tiTcdvNoupsIc7W4pVktV2wEdIzT7tL6ACS
85H0hYub1nB9EkGuzNIqy4nN+5vp5pWXY9B8kKYyiG3ucmdK+SdlagD5Ml1Q8Wga
SxNO8GNVwZwGwACsnh2pYRmX/MPzcxKb8qgH5j0Zr74OZIQCZqx221Ykp/0rE0be
WotM1otMHYLo7j1loNsBKB0OucgzsrM+dM0H1komoUU6gRMjynzXWv1JMauJP0Bq
Mqt/4/e8yfC28nQjpTngkxLIo8wpHwhqPDwaNv760bpQ/JEZ7iQrTE6fypLg2UW5
yG2kAb1DSpDti09KlaOkmoOzMJKy8TWlYZOIDe9Mf1Ij0XcXPaqGTG4ORORYc6OQ
aYgX77XwnTB1JmKdEsqE6+wE53qjCdf3KSVfmrchC/tmoqhTD4aAmveznjT8H0N1
EEJHihf0KwUq6RROofltOmdKL+UcW5cmA9Flt23KD9qFSmsJDIePK+sRegtVm64k
S4krrur46j1FG3Z5dOn9HngX1YiHuh1Xof9fEHwZWxJJE3JPJTTON/OlxPSVLBoX
zPAJwuPjUYKfuGBL5VdI98f8eArcu3T0DA48FC4vBxPVCuZHXap5gY1Be6n8RDNM
IIZll0UZeGm8lp6NRdkcICP9+W/YhjETAFb0kuNJYKgzSipdqpZjhokrX0UeoyB9
qinXY3ii6iLEABOgQnLgkt84emtqSDYl/bw7w1gnW9O7vM3PtvXQ0KamFQAkrVdU
QFnzQpJCnp0bplW4KteU1c1LqR10Zn2K96iNRaz++uaCmzRdwtaO1PK0f5oyjTF3
37EQzqywIjC1fh1fDRKVKw58H15800AXY00eiAD6RFe8rOMOQtT9XSC4HQ4wMYcu
7luFjXQxraI3iS8KzFgkVuAH9GNDKoUQjBQNGXHVyUf+Ekn4S7PFmYD0+m/KKAJD
c3XJ30yQbiFyBRrvnyZ10NHaANSWQpoaOcNsTafYyjwy5sWYTIoQA+cYbjewxBjM
/P9vgIrNCrh+EVFD2/Fa2W/3fY4HaTnpCKBKjO65pdA/5TtqXAdYbxdD+RLSYj4W
9wclcZJNZWuGqCjDIAmgHEQYfh94DZcO07Vh1w/bpxXTubkANVwKuniZPCs1AXsa
WyjV2MdVHQ32/9cp9Ztgn2pDrxGQXPKnASnWPdQcS+HzU5BBgncukZ1ZWWE6nWzp
S84nNl1CL0oGp7X1Q5EuPSEwpVP+PaCUIuuhWUZsLCRgCae+nnV4VxyVREuIeS2/
2+KQBFROsgk3UI2OOCuQLVuZpHOniLBuZVvqFlCgDIskUWoBxvD30YuTyhPfrNsT
5S/fRL/bp8a22aWyuqZC0utnv6n3UKpYpzeR5FWjofX8nwzcix3uhqJR34rJWEDs
qVsJMIZ3n+22HrxDQIGVzY1FItel3s3LGi+O0BMXKROpOfjOHO5tw7YZVVBD/zP7
aYqVbAqM6HTOGP9Pn1KT1jJ5fYsOaAzKe2c3kpH9zWCT5fJT6lQMp+nwhCDcaABp
Umg/j7KCE/KSVTItzSqdxqLUdzzJOiSLD3QNk8q+w2PVg3A5kUph/NAwzaf3Kv9a
QLUPBPgMVAOfNi7rMCaYR/IHKP36Tv4DYFudDzKiOOi1OoB6PxBdNqSSi73htSJQ
hVX4qS7vLsbtmnnzoPVK60PKr2gtcI7stPzDCBec095ofVolWCDJbJudVHyp2RAZ
Q0ZV4JZMk/39oVk+0PgsPBzoYK5DP7UGCXa9w69c6J4l9TKlVCaIi8Y1e2rAtq4V
oWEtwpVW6DJHLTvcus/2Dd9uAhO8ygmdMJxDPM9hcxM5XzMweMo/XD5dOLl8EyTU
AUPCPvMqVE37FVCBt4yHJnPVHhoCc2GgcpSkduTLWZXi0cCJ/+ijlCh/TLXaHiYp
xaPQvJS+97stN3joX0WV08FX344w16LZuy6jjuOAOvra7rCCLkaC3qpsNEQsFjmq
hZC68VefWyUXFNWZMolf4xA5g5MjPaLGYpuTs1rdtBqeb7ouVxNfqt9yYv7ndMyA
97aAVwTFrq3dfgHsXsMkkM9EGq7O+1KVFNgkUYO54ADPpB8pLgd7QlWrI5ieZVcQ
xRoCOMRl68hwM1L+VwWHrHRzdKAqGTDUR0V/Fw4xWY8cGfzZifPH5IjBx0sDBYBR
QUkB18zbMqOdHyG59qd5qzFi2WkR8UC338E3KYtqieo7InNhfyO5FycltMg8GBib
+6X1kI241zSvu/zgPkvlAH1pRt3RgSDDZ+cykC1F5r/IewLuToTvCPyleYBBhrLO
5kfiHKrBeTZ5f23R0eLoEV6Ahx81wptXnnSVukH7ZR9e8rEYh58cJCeekd4NLuvD
pDRIYDOZL/d5eTXnBnh7atMenVPPLjdT87o5z8FhGr18dy+jznHH6tMbINoGhOvh
CoRXtlk9Z+LKqwBXMIQc+DZ6vaX6IWmG5SktgRaPjWgLMERs3CVsN33HjzBOcfWz
6GjAzCyn+ED0JdCDj8w9DwezAfWZ18ja7prXPGhZgMDZsJ+7VPLQSDCwgOUK879R
lcS1CeBlCtHGjax7bSFbpPCDs8gn5kKHynSd+lvFvJQ1Y2k3jYtrs1C8lnKRYROu
inHynqgUXvVQoc2tkpODrSuFdBYHqh5o0tvKesBTAPJI4WUW+MR4PpbRQlsCIatM
JyPsVQ5F0/JZiUX/jrVdhLt/heS12om0JOJI4NyLJbo8H9tr8LsxaEdeCkGm7KBd
adKm+itsgq6SXBbOi2WnGVzl3YBFBlNUejsoz/cOBszYm4cjRN0L6bTYB1BZv0UH
3LjJng/YnwOhE8bo7w5aJOLwmNdAnHonLXEKIIfRsGGDywxIepfm/oO3k6En72it
xlyqFzrUIB/hUs+yuF72vCxMepQTp/GVt3H31g+I17++U1+l9EUooQfehp35CYdj
vxB1T+C1Bm1Rw7HuKmGFOdXOHnHQ4jmIxmok0rpFTvW2iLF9W6U5tiNjs2WcC9AD
kdQGOzJpcaBkAm0Lmxet2V6OtAL9q4nc1h0emFP14zMX3aYtGiciSA4lY5jBwaq2
3MCb1eaLM1J1MByEHT40sWPXj4ozp6jOctxbDJINhiEn/+AkNPHbb0t+ojM4DMWh
Nis0k7PoFoaHLpv+aTpys3VwRRDE/0ml/b8feuzQUCgWi71EZ5Z10Lw5yaZTnzNN
7m20iWqbIOywrP6yt+HV8MgEhs+Ogr7uAo4ZyKmo2FKG0cUG4cbK0EZOoPllXOhM
RcE74enp4gf/p8hMQfF03wjAP59Lh90MUSFJkatlscoz/63y3a606OOAHZcN/+gB
eLRc7/z9RzYOp+mdr+gegrcai4eHzZzN5YMhoMHKe5w7CSXNGyqle1I+cCpSghH2
utHjZXlCbfILWxXBdrUcDYenWkrW121SJXRLjl2AmVTrzYLVlYJk19eTWV/xmKxv
k013Ku00o+UgCFX4l55N6zmtNqu+rZJ26L+8iuHAyFsHbfEiHYrWwzuNmnqz5N2l
VbL7YGnShWEuHoc6MFymzC8k8cr1+pr8lN9h4P1lZR+sarGUGYyOf6ZnedrzecyZ
nf9KbMBg3tyKd9bgHaVXOWKhZWcTb2JICzLlTpz9cDuhuXxXs218z2+QAK2VKK5J
e1WleZv/90Gq8zlz6s/TQ5odWt+L0ScK+mysk2xEv/W3z+ThomLcqKdILNInMTKB
dEz41ZetHkJxhf/0eBIYjTu9x4pMCqESDk605AGg+mr78fvWTELPTAb1+l0RcqRE
qdb6TSBRCdZ3jKwI+21dNn0FfyWbY9MtscY+sTYUkXinUHRwzUToGJ6glLHMpCTZ
pd8XCTUdBvFYYitxnBgGJrtUtNY4xoy4T3LYtfkhz4fLR4MXztHWYVxEM5rhF5lc
rQVvqw0PYym1+E6bZ9SthZuKB1lPflinM5ZY2Me+J0LnD8v1rWwtzuydXmsieMOx
YcE4XJkIal/UJ/capkq9t9zcj49PYwCY8Iflh73wBAryg/JltRDMyT8k0psvCElj
7vd46j14QwusUQJ05JdWdP+t5LWrebQ4MKE2hJznM0m/5mWXm0UucM/CgPc5WrDr
IFoHAt51CKQnQH6GxoKuCYA+DtqE7vnyFOPcwUyJ77ZPUGxfJhGFXRMmpphZo39a
iUoZyVw/HavdAhDA5BvvGAD/J1WiWmPGW42kRmSx4xoYA1jxC0r/tDgELw26fWbo
weupgyFFUT4fWhq1l+f22ePS6iCoV00UXFKGt+fMcWlK8/y1MYpxLIJk/6K9wxHA
0tcxflpWOKPSMKnXv7UrReqk3QlapY8V+Dm56i7LNtuv7BlJWqZ8O4OItZBQVv6I
QCrtQLm2Gl2xewEa0OSxjj9dqTSsT0l0c7oBDAcXiJPBKKFFRv5fzxCxB+spLcs7
c5NUcRjPjOVuOWGMaFxZ9V3VvhZbSuX2Oh/lCGIVufXCQzDAC9+6r+lBqj0mHdo8
e/SH9LiJ7KJ3fJzL343lMKgvzH4sggLdZUzjkQgKYo2hIskBTKn3UnF7QLLjxhIl
FdDY910WCkeppooBoN1SW9UwmMaYWAIpRi0Ze9OBwLuEMg2COjlhmosg2SdtNkw9
OUi4cH7wAuVwk+HyySxlEEDY9FRxsmzLSnMu4Nde1j08GaX8WSPtvzpu5WJjlTeG
4V1EKo1KJFGQ/WjiH6i9NjQGzhJzyEleEcnTZmMPIa291goXwbkA1NrWpzMnMOx+
EyHFiWivdI9ya0fplGAChjy4MU8CwZv3ReKj8RAGiS4tUoXhnKaebAnt6WGMrDQ2
lLU2QNHeV7eAW8GGOsdL8t8uzSg3S3uUNY+4j3n8/M6+xSrdb7ysU4+bsuKeIzw5
vsMVa96cqbGI9cHAusiAfWGGGJBqOCZjp0E9GPXPhjURRjPlMj4EO6pmU7adZfta
lyiGeHv5LhwhnimY6waH34bkogtZv7aTD7oWEy1obj77lZRXajPQICPAvY8wv63l
ZrpQ3EelgjqazTZE737N5S06jmAZedIXGPXSuot5Lipgxff4JJk27UZWHierD3O7
frndwi4szsQn88fXLetBGOYWBew4+q28VaAUssDWVF51zlYyFRWAsULS0qYSChaf
RQISoVu9tiOTEO4nYxRhp66O4uxzaYF9mYaTynOkvfuq8n7QQD7HPqJzKYAeOKiZ
2Brihu9EUP+xz42LCyHdg/s0nxJgVTmLaGmr06QYMY5MK5zmpoZVj0ZXxt0z50Xs
PetUq6a4bdFNjo694zByaoOL5yR0IWDdCxp2DSnZgwB3HmVfBPesIWu3ZK73EHG6
zOfEd6iVYnLnmvq0dBpmHm4UxRCnGlj8aYaTEdoSqAyY9Bn/Zdrmm1kdqhliRsrO
LNHV1uf7buxzTdIESDfEZPr9GZhX9Khp9Si9Z81ZFY9qEx+fxJGljYbkgiWjs/UL
06KEvecclzoKomPmVbvVmiNwK51la6HF9hCGZ99e7QZfTGuycfgmNsMy0+t5C29/
rrDBdl2ydPtL3N3GrQQvfSkoDX++paTuA4fwNo8Wp9GdSzgAmQLGhdP10dMWHmcC
NByFHbcQ8WFE0iKKg0RdhU3+gtAK6uAbZKSkVAnoAgZaz5tvlhhb6iw3YyxKv2Ee
2C6jv/HNZ8ZotW/sfZalOqMOkQDNlD7Ro1mZqjrRJO0xW50ERCWeeT5rBNW5om37
6yRdq1Kfi8L3PNhwU6G1eYPqoj3tT71gnti/0+IPC3F4JsZ4E7gcgFT30+dsSW7/
YjlL9xS73b+bX1nkr9/2g1cE9n4znw6ojKzGU8w79w509v7PmSi71K1sjmInl7G/
zejevD34VfR/bGgHLwNJpi7H46Wv8UFpF6UJGgMJMZYTvYh+VikRFL854OBiOp4z
xC8xaEwsiUALCb8aB5D5+VL41WUTsEozXLLVHA63ev7PHh/aB7bybi26Lc1/sObb
GYbLoRPuMHNfdaKa529fpWsK6zW/lFYDx+uhpffRrLs2aHq7G0sn2gOPxVxFcoqB
aqi2ilXUeug5pDi1d8zYftv3AI6epUw32vGMw8YPFAjXyKAhVCFc9k0R2UHBLtou
JGA4DLTNsXXx9g6sXkqTq1CMuk3zsZXxpfF5nQg0kGn80pZZSR8awMxrGHBaMG/X
2k9ZvQI916JqE7fy4ZUHFZ4r7vc4HRYUUse91WaDaue4M2TByXzFcnK7d2jg/W1z
aQtskO57c248bs6xFnof/dKFI9NCB6KQpyI9d1F79Chw1qXoGwvQM7hGwI6hlffx
aShb/lobA/gNJ67owuoXBraGcBzxD+cv7hjvb63PB+lCy7SRDIbKDBzaWoM/ip8V
AtT1y5UZzMI2bL/SeIBi1Hh2m2RQwY/3iVWYqTxHNtOe+K82E9YUPqYycHJrAGO4
KN5ijD2uU5X5XjDSBNiNDzaX/kRuKzrcPUMd5HUw46Nk0OPa6Gw1GzdzlVc8oTp8
o9dJxM65R5K5vqBUUlSLZpPJUenX2CmLKHdjodxpH3DIqAJWokBX31RblN/DVPXV
rs9ExIyczocj+Y+zpIJE5Cn49YTLPAZ9tCbnXPKvVwyue9X4wqnXYf1ZRkLvlgw5
uB39XS3mzwFzWucVVMf6QJEmS9ApJCfYIW02k/8K5KR3+ysunfINJORgWbhvOb6Y
xMvTgHtGVOn+bmklY38WC6S73pxmz83/t2wAOLlqTBo0BGvPFYKlpRR6juy/aL1o
RsPkHxjSHyfc1xrQvOOY3M9f+TiskECrmDJhEJi/ClVh4NQWlqlThD20PzQSf26a
zi/efHQxZx0uiN3oFrVF6Cbz27l+P74BjG89Vs1TJ+xCB35aMlg4rry7WNxrHEL/
6JeO0jfQNryc6bux28lr9BCS9NbY7co0EIoUBh7W0a4T0oQuMhP4+zmD/C8zjBxV
t123w4RWOe4fLOVmiyqMluZ6juEHD/XUY2slVRaqq3IAjZbyTcxxtZRynSEFKFwE
VHSsBjoTY46qx6tmRhh8Froxny3zJB0F89ipMBFHyVswK5QaZhKLhscsB7WDJGeg
yS/zSNQi0cwmUh/TzmCvqICLijcsLdxJ3M2u2GQ9TiNxk7obWt+q80JkarYpvFa6
s40P0T4FD3dwlsLG6b2o6ptYXNnGxGTceAFdyqhS68dAgnbslS0H9RfVs8Eg1NlQ
HBypBdQ939Po/rjJ7vYlTzWL4W6VPR5S03WXaiaCNK5uoQeAfcuffs7IhzfJcMdR
S6vYc7lXA5brQ75HpKsjE+o6nM6jdh7iRDsVTgGmKzDwbpYp6pemdF19as9bGWUH
YDcygRfQtmBBC3HfAAARTM5HF0kVQu1a3ac7PxHrD3XoI4HewRS1r1Bb4T1Gbxzj
8hUeriJJyDCsyAHh6SKztQK/pH5eDVCxnMbpmJPlpdbSR614nQnNAVDs2oesBRK8
0mPOl+ZikMbvSsN2LIjE9u/oYx7Sybaxjr3alua0BMahkPl6HSvPdfQTx5/FJ+fg
rYxODRQJ77I+BUxl9TBLUJrI4LAUHJk2iVBGWCdSnbKlEsDC9ZzWZVww4U0k2BrT
tImQ5EOtwZ9X/rsxvgGDU3CY/aZRoOVr5wekosmYJ2dTwdFUl2AHaa+vbsMZaa3u
Ix08qFGKsMxVIkNffBzGDxbewVY7AHCetn8eIu//ApV33ZRn9g6KWLocgJBNMplr
E6i15B58k3Mj7PnnNkiOA9ryAAEEjBIkEGBZx4r6F1JftxfCsoaUv8Rude+diNh9
Wh4kQ/8ZpZ8Tlzdl6AT551gAbYn4xdGPLVvV79MTl/fmHVQ/1/5l6ynUFUxVzHi2
TdoyrbH5iabWT9CRe4r9N+euODkDTQ7daD5r8oDJ5jnIPGvMhn+Kc4vwM4hl/Isf
2+z+IWajUy21q260nds+6Ys/dgtOK5gZh2bGWIjw2gFNRR9NEpqYIAsdt1qQA3qj
fxs/l2bilyFnUuQ8keKsxziaqxRwb4Z6GsgbcXzSD1xwObE7R8Dub7F1EMzjElvS
8MTfyLDNFZSU0lhAR5eH4/VS9DoaID+K8upneLFQgIatEMJdkaAJg5PlUNo8doOW
2yDAu6NUWbxmdfLxNRaSJfC97aI5weqQE9m40sJRtooWgt2cA10SZ4Tw15p/6VG6
0dPwhdKMoxQolhTrTBFcwT8Tp7V2h5UQi+ONseq3ULKhMSRf4ZPgUgxaPzuwZnC/
q9NW9xw9DkKegfjpc/vi6vjMLhaDwUUB0vx/+nWDZIGt/DJu56HbHmWZZ1YfJfDz
SAxfd7jpvub1+jfj73Tbz/mBVM1bP1zcQrT+j71SKwO7/5jNOPue+59X5oVho+Hp
B57I4J+Mzvlkm8budt1n2rf6WpuKbA2ZXTHvzJ+AX4+KzC/G9kJW7097paQaCSBy
9eEo4MKrRLrh4b1XKJmgbh0A5pUvylaCf8Zwan+rnB5+bSCGMh5j6iVDrfttRSK1
iM0cN8r8TqhdyuWyzZw247ID6eu4gnCtK+dN9uVQnPLjdl+hsTyt7ynKdwu6IvSI
7UkdiOK8cPKLJg1t/PKy9fcPpTnSZa4aQ52o+kkjG2poCMgCGRUi11TF84PAMsl/
gGXF3iT4uMyyPKOgkkvuMgGeLcmwMVMQl9ooSIcMqKwSLYYKiCk4vTSwLd9RqETr
E5/vbL5lSE7vhtHHUNf5CriqVWFsihGqS5jmvccUNhVGq6WQyIs55uQD3ssStodX
MCL1YjqWQ8DUnNc3eTaqaHMKvkzcMXNYBC4WRAMoP6blcmEyOvDawgkLDB6XgTW7
vgtLuod5yHFUudADZoHkmHAO6XRLVO0NqpQZ/wNU50Lub3Eipb3xNiFtMf3uTsdi
H47v95mAtC9cExiJKQTFqKREySOhucFuZQ91U05VbC92Xegr7hY4m4VIUSF1oQ9x
dfYptnXsp33bPmPKZzlFzGjcG2KaaBWgoBvbPWuv8B09cEXGXfphPbBEajqh+mHB
pwSlCDR/zPL0IcXePTzecHoBeMJqXA/B4aWQpuvIumYxcOuerBWdGfB7B6B39PrZ
XYuKUbHiKQAh1HnscJb9rmnr9gf+xMU4e4dEN1kxDYTvndQ5j5K8hZYrkHcAuGLm
LfQ92znqwKLlyz/qZkpJGFCJTd62CQ2MQhJrqxMQCh7W4D6Zy2vMIDDG6Pe2QeHi
k8lEEBPW7HoiMre0la2AEMg4rhphkNy6faSWeZZ7RR6McY5B7Fb+1VJ4q43Qpx4M
FyqCadsqqmfvnCpODLeLf6l0QRHDMPoqkXHbrm6yTbtgNjjVuZ3EK8Q2ZFWKJ3j4
LoKMtcJwGodkr9fsJ30L10/6JL3fgPYDwTKtMycd2+W9cCHb1kOOc+dbDjXoWUuU
ODtq0lne8VYgYkHfRcN9B+FjM1pUdy+5KZ1xyUAdeDZlA+MliBbTNTCsNYDyKti9
SxfMGmRnwpB9RrOwIy0gjs2RkYonoH3rH0hcO7dD9LmcR4Jq1wgaDWwPkYxiUaG2
No7h1LTesy0pZSnbAWCpjrThSTdSnKikZKCTsnQzZZk7vXLEb1f0ACFpnCa40UNX
NN+iK3juJTpi8GziKOrQA87f7oGEJKvR9m3+TATVA2rsa6J+VUQjUB2xqnpZj8YU
6m6ejw2YrmRmyZh8cYzRDg==
`protect END_PROTECTED
