`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o1yBJmd5Jel+R2KEgMhnO/FyFfpvnbnBouvF5feG7VOY4c75UeTGtmkbIsojcxTz
njLGuKa5I+mvvk1bALo2LvjLGOWzZG8INKFW3lotbbicBheqHThvgQPWosXz5z/e
sr9tL1Sv82RLyzQgpfroKBgJ65bUilrNvQCun6GxnmP6YKn3hOrYSStCW98NYwiD
a7SxHxSLqUwKpKf62hEONUpiU+wSPyX7uWGHGiaHmRpKZlR9VOjvZpofSzo1skK0
PkFsI+EnU4q7DdNGgmCG5Zh5+i8lwRTKhZrLDzPwJSk=
`protect END_PROTECTED
