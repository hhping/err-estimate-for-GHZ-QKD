`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VoLpkEvjPVEHoB9Gq/NDQCNmNWrsydx/HklfBfUp34B36HMLtJIqcS+EinWKBBmq
N/TS9jhn4tC36tPaGGBdQt2ruazM063BBghlTVdHeoNOvpJ3RWEPLO0Kv4Qnq6/K
KOIRrmc4edDvaQQPIC+bY8D+HfRi0Za38gYtQUzJqCp5eRYxXdzz7seG1nt26vxC
8X35nGrnEgVXs79is7S5dSAUAq5eo3HoukKtFcXMgDe+Sc+w7GRbcq60n9jmmiOA
7aQJZGb3eDrl1FPQPH+x/TlVo4PUTnv52A0JDJEqvlCPae2gwcXNHYD5QW3O0Vln
kOG4wr+lwgmHq3lmWMGKachVGnblTUMbL1dP5IEuxx1sOUBaVw0DzO0imXEb0bR4
7wEBvMs8s6vsyqN6cC2FDwpl6+jx03+L97J6WAxfDHbEr234e+Q+mpdYqhkuDHLs
S/XKM0AbVzfZPZcVomVzzU5jNwjdomiVTGixPs0vDi+hOQyI93qPBtWMpSol4eM1
loQZ/REHtqyGC3EJaWaPK5d5XicsO+b+JlDWrDwYk+QxrmnAHUFgryPtKxTc8Txk
CtmxEa/E/qmOmVOz8y7yojCT6biy24qWMPh2X1nQinVI4RL2sMbkWHUVNF0PrXFF
g1q+paa3nz+EcbfXPNSL8z7dVEPHPW4BAFRIX0K9Y9KLttNkOU7aUCtV36mf/gaz
FT57Lnlre38HfeL5iU5/XbrU/oBIJ9FfS2O8j4OsFQ0C2yPiLhmzUwbBdNWgAOZb
xYxc1mIOQQQtyn5wxE/U4Ny9AdWp6nqPl4pJ3MkrECOKn+FS35NaLEtnI/iI917u
loTkLhWGJllA37Lce35jAHAVN5fxtqyV0zkVRcTS1YpGl/eeIxAifW/8L4lXWrdE
A8iqZgiKD1UK3XZcHO+VG62MaufufuCbEAvq4lkAHt6J5t4lcACCfdIXcxiYyaoR
LhhOgkj6l1QrY/I08dkSiL4NJJw0g9V5NMQueDM5HMjSRNJKolQW8O3XoHrRRtW1
p/RXMXo6SCb7Egs8Qesj/g==
`protect END_PROTECTED
