`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PPajmzqWooDUUTJG1KJmIjgKmjz4bwyBrHDcqxXAXJwm6aBw9F1tDlN3IZHE1Fpn
55kNmRUNUwUPY0k3BvQrJBgiRnuql4wTZO3c8KV1HGZJlQZFxn5NOb6RwI1nIeNV
+pRwb54XLc3q6aY0bx0wNvNK+SanCLdpVY/gYvRRQQu0qzrFBfUOSgtC3SbbEcdO
EiAnHXUn4Dk711IigahTpLu18sfkhr5pGQMVLKOVg0IRmAHnl0hfywyM7ezf9e71
LZJwXn//VqZVt76a6Uv5B4pCSmXjhLB0scHHM3oZhEa/OV63AFHa3vfFRBM9Z2Ml
fCJww3CW5haR4r7MyYZjBO2frUha2oLkhhWyxzZOt0Y1sGzPFkfs3+ZOzbZL29hJ
fO2TdVqcL8LSgt4bHTrxqcmuui5Od6vqhHZACvKd9eSt2y4cike05woG9GZcl7OB
ireyyXOVzKToW18b8kDpUxME7rsjI6UJlfBR7PJydPC9jLLzPqyDiRHpHqUUxuzL
ao/qT0V6auqM1dJEaUzsCnqgEsDbxC9SohfwDEAJBXAKK36do72RYBu2wWoKKj1e
nlL4bjmCUJerKp9oFJsAI2f390EcX5PYTyokbOj2eryCZYvv5lmyjqMpXM29/0xg
OOjvuf1Mhs9WNQ6gE+t9H+rsHf69rx54r5Uj/wZRVejCp18n4J8FPvjuwJ9C+OX/
murSA/qi7I1giCNcfXVirN194jxcY/CIxHICsst79/BaL7xdV+CtQKuqLn9g7HLB
aXG8I594sfX3E7HH9NItcTzDIU8j9WtSprGCyFTZxPYLN55MTqevl1t7yvNfcb20
aFaeAGCW3+rdxJe71d4eTZo8EW81JjcEj/cz5Q6mTVmkTwEuI0u2UUvhkUsdOpzw
11w16PfYvDlSkffNch7vD6iSnMnrYuwUZnOb4nzYFQ0IJeQsHjweJsrgsUQlICQb
GjvyLyCkVkx1mIRuCb6sgwjwqCMUwemAAjcId3tnzTnPoU0CUjlisdlvrn1w6XHq
r3jOSB/g1CJw0zLXAbaMqbFng8kzoMroiNm+F29hk581+DUPOVyETT46pD+uc3Gs
Uv+LNh4crEkbSnWpMA/RhO1IYvmAHmcXH5QgPCmc9D5AVJKQjlyJnOVQ/+8dkl/d
JWX+O+sM3CeFp0mHXjq7VqXoru3LK30O89HbJ0oRzQkkQoGjw7eX6BFBe2ZejnCj
xvppEBQs2O3ECAu+J/pNhDzQshX/f0O1Qeo9pAM41Glbdlq59t6QZ6gOMT8LITfO
Oa8B8PyQPdvR6FoHcWqjHi/fRsHJlWzYs7FS/j1DkBHNq6ckYnoSKUXqBVoHcA+x
yjrcsayCVXgg9tQzBW8I1aRrBDIwaEs2ieJALNDlgmsx0jQ35SgPPSRBMO3NOtUB
ajIIe0GGNlxqVXLnEc0prA==
`protect END_PROTECTED
