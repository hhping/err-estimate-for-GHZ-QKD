`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tr3OMOq4fgUnEOlwKCflAHOwok/6jUagJr8qiac/M5/VFyQCCqs78VW6NXENDoRY
Jresifa/o56P+wXEH9JFWYF9jmj/8gQh9ULX8l91u8Ce5Zd529hgOcaKITyGDGgr
Sp98WtwRsD9Hmp3ADxHmzJ+BFMKKk33QRwHgNmqIZkVtv2/SsqlYVK864XCxguLM
0+sAw+g3iSppOocLqERqnhr2/om1FGaClY2PDWCu43HIUrv/nDD0jyp+Eh2Vwb6R
/FUjNh/BNcfU1aI0YE8+P0qAA7eaxPCrXQEL04fRpksbkBuecu2lrZ1UPW3bL8VO
MsFDrKLA22sAEVpeMrY/lwhoSULGjUrRuBS0VMaQPYtJd2YcSekPc3JJKGp+N0vI
f8jh1fji0b21nyFGtYOO4ltH6DHIfDP47vh4Cjkvf+CiHWU+4PEckzf8SnKy0hqE
9Wda1er928FWzjLUNcLrvXZrQTCEFOeQ68ZK9zY1jOurctWWKcJoyokJ9XYYyH6t
VBiFl9AwTMehxbClXTfpuAqlgvnCOKkMhjZGTVM/YZeqNvPeCYfm8vqtT2FT1o49
BII4b/9kx4nqHuPA9VYwMoSAaU2uLBNFJ1xSDu7tRaw+l6VyD6OD3+uVts1jX3Au
FBVuZUY61ypCWnxWMdOu8DwobchViqfJi5SehxlDUbIZruczpJfq66chytoorjfz
sNamsjY3PxaZKJYb6q/oMO/vfB0ynXFmtMCy4XraJ5qkMZXAuirOGi+0qbS2pXXD
zVEutvM+DmjMWb7c0kcT825GFneR+PM+5i1P9FQX4j727Xn9elmMAqMkc4ggKBiN
/zlij4XSowLgPoukjjn9YTpk51RB1UQiAnEwu4X0aWd1BVkIVv88/YQC4+HDwfi1
9bwoBcwUCUhwjBlGWPPrbnxkEqiUfpqISrFDARgo7Xs702LH7hwT8Bem37Pt27NN
/j5UjKrVKbZrYg9US0zhrDJdBROwo5pWTmHunzHfUmE/+F95DncRdt80Pmt15fAJ
eNawaDsaJKFO3qkQXM6dGcPMIcOG2YDak1+dcfw+5g+dPlWGkfvOhn0qBlkPHOQe
pEjHOGP9VKAwriYxqqxQ0TDyAKYFsmrbpPpRn7+zQXYjtPbPTii0siNkhb+n9OYZ
Fc0p0xgQT9erH/a6+qDfJtO/+lDwx43e/wvmiiPo0lm73UmXYMPIMlYf2ooz9DNC
V3nhUZKBNymKC361tCh7v0wTthQOe4f1MeLtj0RTbv/jkEj7p/NsIvL1+F8pGFfm
djnphNakLfrrhMmnOAIJDzfyviYJOe4lMd0QVsxXgXoGFPV0lz2n9X/YuxEJfMg/
/nJwGdBHBGTftdRlXZoJKMvm5ljCHbEiUtSYlk7R6j+FAIKYjgbP4TrHn/adhVq8
c8TSfLy3jUhsiejoVl8q8HlKQ41BCNnLEXuJM83sSfMLY2OJwagSI/uK+eYDbVbN
8jZ0F0PVET435yCyEnRDzflB9hAQdd8gKxC/O/AzmZx/rhuCHDQvCsSoH4n1JloW
XzRNfYrTkjxdqKOmhFKi6MXM8z2I5mret/1jZwHg29kWA3023bBbYP1OpUScF2KI
FdCn+xMglbG+a/TX8E5ktWxHmyG8fn53fs1dC6l4+lyvV1ec8cDtlXyaXsdNYUEC
w30MTvi/RbfcrysFsxcR0cQDWGDWAuxxjK6pr4cBnT/et9ZfQgtMhxlm+iTDkA+g
azgs+FSedpRjUecmD2pHhvE31/JQs3pH2SF3cV9Ica13QgVuiHBcve90IBoyxZRN
ejlVQDsFKBiMT+3HFg6RXOGeubbDkVhaG5RvDs39/uy1AYpEcgbq3jRH9kx9vRas
kagqQVb9D7U14uuQRcd3dUth+eXYnVpvHeV7kuH0VJMATwnlyfjMcBkP1zpoYH65
2ArmOcEM90quZOnJ+qGfhHIYdDogsfuOYC1TTmMx/ukNm3m5uaXPhLpb6Aim8Xaw
bT5bREJWsR3CGaI4qOXkXjTL92JVYZogIUUMPmXKKIYe7TeP85urD9fXK+geNMJt
uEsIdcn6eQQ54tvDLkurIcJkoX2Mk2ykmNlNsv9Kccq0BWf7xvMFvR2j81Yr4bVo
XiiQV5785a1oDxBzViy105reP28uzSUIq2LPDvRo5V/9E0O/kst3AHD11Kuq5u/L
79BFXYnrb+1YkSuq1+0Gl7GNqbOMC874Ny+Kirr9VCIx+sgIh+00oeeHqSzHI2M8
rD0RWuZ4ihWp3LK7X8oqxUl8E678QjxpXImOIGLqAT5OYaOkVgN/M8wq00ft85Gx
61IURtYxYtKKDPlDxROBK1XH3frnUM2bm5fpO9qHzqUAWLYKNjjdRw/v7vVoj2tk
fkS4R99IWfvR/CzzrlxOc2UmxCdRwF1uirvyw9O0zzz87FU9PEeSoi1ERFUhqBl2
jSEEAwS3f9yX7F5zfk5EhtG60v6BYTEWhquz5rcdxEszG2DPrxuez2yePt4juaPk
vSyFgJPapNt5J4PPKqWCl6z6HryNfm3YMwRB3TtoK+dQlJuoZ+3M919yhI7NRdBm
iKGn+yKDGGYlhgsQgAqa6AjUf0L4PeousTiGauk5J9L0il4s6pcJY+1PjrJOS31V
RF3CggAnJ74xWtdh3pjSDrSDTVNeo3ha8WgVMs+XVRVrC/iBy7vV61dBNiOFikJ+
CuZBCzhOAAtwPLt7rR4elRDRRqsdhU5wd+r7YQixVyASbgUMIXzX/CoJz2PkC6xg
kh90HOb2QHbV8gaD+HrHHpt3o7+HbGW8t4cLcIr1YVVMI8ptbKSVLYU5cqUaom6u
lp+3jcaPyfy/eL06JbeNoZS2CpKeyccuRdXVKPOW+vCM/t6L4heHD+C5hDk08KZA
d9Dc3TKdwl7XZqWFqMNyYF0D0v4rwK/cTgBN92R/VFBvxGNBGRkh6iWH4dkTBclp
KeX98Jah9Oi/oFOtDxKd1xkvp/lrRgF4UjDHGG5NAMfPpc+9yLAYDHRgPMc+OmD4
hgpXmcMQQxiCfdalI/4sNLwlB48b9MTVKNamYUJxwMTGAQuqxrnsXoHwpvhs6pK3
8jWNrwOwkaswmQM7kI5qJZ5o2uu17VQGWbo3YhLrqta5vUag8xmRWZkfTZsApn8o
9S1VxEptfvYCqiNi2j0Grf7oHGZ/57Xkmt1NRJcZlL8UVgwSy3BVaQbYlWsl02Bw
qnrVAdr2whtMuTsCcJLsXk733QH4gdba0vNuWtZKkdK3UWMKt4pI1ClHjlycfh1J
LWqCm4YbkUDcSie/kmdqALtjORhgSQJu7Xx7zi6ad9Y3rKEpY0sp8BpeJ7D6oT+l
/v3RuHT52p5eFJGwnwMZQ/asYeJdvXQxykallwDbwmwTJamwArfYpicPjZ6H6xcp
bmVIxjSaE/elez61deX5iR0bT9k+lRVmt5SGm7bJwGEvm9WpRcjZKsdld8yuy87H
TOu4h9QhrL0E5s2QDxh9E9NH5ldLVjmqfTGUWiKF4hKrGw7aE6A75VVRnD6FFsOF
3z1V8RpupNXI0L5gnFJMAlvx4w6WdSqRKWGHIgUQNDgEagCvGkFGAuVsBWLXvEdp
aFgRJFqCfZEedNTOfn8YjHr6UBvdnSSoSzMuPqFzYpusGdRBpWka2Vs2Cl68krYT
Yx2bxsomwCM4csVdGqshR9IdfYCgKsfXAIDR/JcUztHUAPZRH3mgfiC7cxdWcUgS
vM8UCyfX6PpAIuxsrH8DTKbROVFqCGGs0CMw+8KDVXp1YMHw1+5eG89U6AYJt4vC
LTOgFYVRkaRE4jKK8uc36o7HkkUMaTeedu+3W0qXJtxsvCWyYDLDT70mbQg4Mnrl
DVVUp3q86xbWKo2HWosBZk7Yh0j0btpo2x36lbOwIQRDNr9EX0JKpSVi+XOU7RtE
h7aLDmFycJ9U+EWFVAeSgDrGxnbfNRlvIoQmZJqUbIsoE2uuscC+xDxywpmbZBJb
oKqMclH85zSPSnr7ElAy7okur+WZd72E6SO/eWMwyV6gnoN0Q0G8/CkFt/KXfDVf
G8xGAVvuRpwqDJniq6ixIdtzVLCl2CJAT0OgNbyQK4c9e/CgF1VMN3gVcdEKq8W8
cRTxD5BQC18CN91qfnBjDdYzJOCQzZP3nIVfeN9wcgcGM7BeXx6+BqEVsc6kFF+m
9ubui4oFcnvqW/cm5pAtCcFihnVTj1mO3Odg0rh5R0ltgsA6Dbpd5FjqJCc3Fj8B
pATE+gunJFnmxTTbp+6qLCqRRjQkoRXdp3j6OAl0cSeR2HPRGF32KNk/S9foHDC1
OaDuva8oVFJQSp7vVEqmK3ObOlLyQtoiJYyUu1kDAu7t945d0iQ9/Q7eTGNfRuyb
QZ3TuMevd/kqa9Xy8r7a1GfF449fgcBSnV1EaqSGoPM9A6YuAtf+y9dCMZJ7+uTg
7LGAnFBBxSJXUOOoYnHvOMu5pir3e3j7W9pdUgsnezeGOe70cvZdnVWjRdW7PlyB
BDaVdy9LNLrFUS3tUQPcJ5K2Tn2is+BQctk6+pUQqsOKjwpJWYBW2+yY93HaB1vA
sXTyxdpRKAaAeteVy9TZrmbOj5hxvl3jKp09CnM3V+7hmn9vRvffPSNcVy9oGihW
p1z9x1gMqKKJP769TJZhvgqJTzivDb3e0gG8s+wQ5UGw+ogPOD6PWsiKra7So5Hg
goP4Ay15/OC9TY/n2wXMKl6i50aRLiVX5il9AbixHuTqynub3cGao+A46OFrsd0V
KmN50VXw76Jh83vQDGbQFq5p0bl1+uwx2xYiU7IIPYny/XZUVgBkuSZk53UvkyVt
lH+ErQ+rZFmcn+7YAZD9RC7G0+Jr7XU5zvj9BC8tL9Oq94Id/oOYHkGx3W5ZYDIx
PmiRZhIsVqy1m0u2DbGoBQyyW+Xa9cRlCWmTvtSXe3Xto7XseE8jNj1K7degF8tq
M69duuDzY5o0ulofJSecKrGUsOXPSdVR+eYEzHlYQK4Jx7ERz30BEcvMSN1BEl2S
mmoynXth9NnyI2KWOvW5yJUSI1uYz2nKpc2bhGROoUHGE/3Tr7j97rmGVqdyeRGP
9AypJyJpg0LzzgEn4qKZ5i2Mp+dVnwgT7UlNIP808zdomYLCAOfHJEAW02pdGaNH
8T3PgQsBuB23JIptTUkrVN6QzsybIEASPT3ecXs2gbefE60vV7PNoCX8xZWrDZn1
Tx8peTUJ2OfhEH2EmOKCg7xZNz3/sxIZov/e6yFTTM98KXAL4xtJcvn9HpAKpzUF
zdlK7y5E7eLuhQU+rX77gksXL/APVrc92wkTA35L6Vb8GLmkix3pT26yl3F16c1w
VsWSzjeVm25CVw1sY9FnR6ET6vaePSHfZlViS075fOl8Ekuhzj43uHpPyA2SebiZ
nMTMtl+ac8q81hYaYK/CRqFZ3Zsr1vGE0HV/7TtRVH0SI3YMM60q/bLCdPbKy2AO
zbufznZF1zjyxGcwjBTb70NA5r62AsQVe7z1JI4hVejynHhW6cU2UsQIxwBr3p/S
HzM6v12b1j1Swm9S955zrpA1vPHlfpqAptreongx1AQASCwB8cOq6xojZOp+vC17
iuWyuViKSfDRLJIxHizRgkKOsN+iog2Jlf06FwZHDK85xlkd7W7Q6JZPv33N1x6k
dC0XoGmv+2PL7/ZCuQghlKdwDJkklYX+BMfL9NA2YMN2I3gnPwc6rdlpEED9T2V5
/9ghX5+EUl6EA3LSBoYrBsCe9YXhIk58Xp96RVskdK/c3o/+aFvvHLzbdq7LV/uz
Uz8hvhUrInnynDQbp7DUxY1Vdadmo3Qls/3lHoCb9QESfnQ8FO1XLawM7GA/8EoS
BrkLtYdCb3TlREAPU0QzXJta+atUq5m0wVg6Vp31aVP5r3guILX8oIU1aKAB4sj+
oQsVbWbshdgboUEJgfeCDIsHUpNaYpGbPuroourayJxiMxEk4II2W88hNIvBrBPJ
Kmxpo9wigVipMxEJIBFRn92BiQUU/sWRr7gkSaEPArRVjf20VMrNdKw4aTpwbg0U
Q5PoGYgFaU5MMLiZIUP5+32RhTEtXm2sBvRcjDUXd5PcdJQ+1W00DpVgFJr5FEKw
r4G5p8mOIrh4ebwOC7tBAnqlIZ8N0C4Eho2DLB0+8Hq6DbZfgqyg5jp4KDWe98ZM
0Qi1dK+4folenkCdX9x2dnmwqJjj6Ta3hqRfET89KpvbYULgAku+qKyKHzxUukde
w9yNOLqlwgaUlMWCWvEGKVkwxlZLEgqrAPtfx8vKy3rAFFgDSMJyCTDl/SgLVMUn
Me58n2Lda7sW/4482XBqfu5rDs6G6rOOgHPpeTbMMHAKMBiIV9krX1I3SxLAy5c1
bizbtCNLnb/eE2A5DEiFQxBu9QgUKKU6VeQEwV/vwwpKS0BzB56k+xX/EE0R2PRW
H98QqivI7RtZ+S8bsEfMjjiegyRIPOO8WDWTIyj4brPCAM4I6DvHCN7RHNd7L73k
FVdfLCdfK8jsMaXjIxsXB3JvDpVCgJIBKzi/zFh2jR1WCuwRPb1f6oBd0uKwd+GG
rFw79GZ49f3OjnWSK3DRh6b+9zQSKtapZf0NqPefHfoR3SGhvax+JDz5FNARSfoq
lW+2wJLk9V4Mwac6Z0Zlmzvey6MNi8203U9BuZnsszDzkfBOtv4T1Rpq5arnpXYX
Nj8ub4X9C34eWZR4kWBBjxi7ATbHnBy7lkOyVjY0Om19u+7QY6ttpQjFjDjIHTmY
R1t58XnSSWrMnleow/I9Oousakes7ElTFmZO3FT4aSritEIh8BlIj/MDQxlR9h5n
pLgE1rdc4dyf8R50rS4toPWzJrMBcVWDUzrlSBNA7wdvSKq8yn8oBNld7uB0Rxat
Bz13aP0tVT+4vvJvt3K9n1aknaSuwMDhk/hYKyGNFGVk/mOy391bjziirXEzRNw5
tUOrw85ukY3j+JvQ4IqI6pIhhSsiZdI4DpbZv93euaAL4j8OfpjUdgnjMJ+9eWX6
/+9Mwv4mKBrkOuTYalKt5fAjHvkivFlYrNvsJiUgiDxFLcu5zDmmZYsnNSFaNzQj
Yh7zOYUYyNkLNkDFhiC4xn7vZvWRsCM/UGC85M1VDX1SS1qT22g8qN9EEbDsyTzI
8QnnmNOKumkE5OPJIYM3Xtdkvw8nWxE0qvcGFc0fUPRUq72o8FTXIkDM4QogrQu2
VN6wcp5o/lxS+C2cR3Mn9S5gajjNw7PZ1uSUbLdds0AaenIv1z24T3V6Jw5eq63F
dxry3eR/gsfBnBIH3NryNfJcfql8GHsnEWtsqT4QjzwvqjyvbZRImr/QZnp78pWY
LxeBnyaaNy3GWhgLTdjfLzJAnYj5DaBUr4AtCx2JWPPSYNWstwr+c3gv+1ATlRRI
jeB7+Y2lip+tDTbfIyQTrSiseyWg1CGoHrAt/ro1oPyluStPDYuwLqnM3Vm+565A
Sacy2RWLOuVw5ypeqkPYYyg5H5GTBNBj4kQst0qqwK3ibAnQPTizYcnx/W8AIYB9
fcfiilGqsBBiedeEfThWSKchGWPnQioltPOgoZQ/cPrf6Fkbodj1EsxnU4XL6NSw
7aCyEFLmMR+5teMrDvM/H9WR5QpLQsr4YgWzTm7nxnWf36SEDdbfHC+IP72MnJDu
/twBhvhykXYfOgd08x2jtMqU4Lo0QsIKdJx72S+OMBa7FmR0Px/tAs4O+okX3xNJ
ts95bMjJLEdvoMPo7rRK5DfcKede6btzBHfnMW3wDc6FI6mmcZ9AKXyxA7uQJjGK
alZpuvrEwzVs4ES9ZTm88BhZswrdGDRTh6PtMGLaaF3ANMdhYG5PJYqBRI51haaQ
Qov4akLZawc3uun2UmdOURVsGXNi1cmYpHxumt9oPr/JzgY3zEWNBUJgLxsCl/Zr
ZHC5M/W6KUQbb5VxEgdn5P1vTV5twaG51d3MpYpVWsgkti3O11KqWJZAJV+N+476
M00FTo8F6K22J0P3IUmP8j6oBWTsywWtn/yvP/gPm60Y+eaNn/aFCMCoVAdoItN8
VDCsqeK8qHfgpeiJR6VG99MvnGLiTMcEi+wCCsntBOVMnAyTN2CYtJ8PbF8MwCbc
paUpEZ/Hp4SIT24pGiqfMSzBhENiQ45DGbdJlX3ToJaxqcKjw9l+ldwVjxTqNukN
NwxoZpnHPdoIz6RdhA2j7Im3ZceaQH1HhunwQRnY/sWDOBDOiJ8K3CkLZZBLqUgw
HTRc/j8qAYrDSDrw+3o7um1LfXdcjXKmShv1VRsxTD3OwjAQ90RmBN7mxCnQzVRG
HYbrko/4G+OETPJlj4Xi17tBrTmHdIcF3T2XjGFByu6kSKY0fZicXZmsX1bwrd2k
nXAmlGH2Kx+ePE5MoSg1972gUTb1sUvKYypRXjd+KeiU2Z236px37aJqBFGaPcjM
tGzPPXRa75BAkNat/gFACl6J8iV0YPnuqhNFkRy0DXIuW0WbpDX0wqbHpeqiaLqe
7J3GKzSnznk2hTp7Rpb/MMHX24vPduGzcyavmBi32cSFyf8bvQ6rWiFM6k3HJxce
8MrvuFKJxQxdfTFsKgkIULN8N2XdS6s/mSUfjefvChl3z/4BeqSfeqwklZw+qFae
ZvPe2nRRWe3u1ncZyLQg9ZTvkOSvqC18qAdp3F3+DPBACg0TBoZnlCWq/QnBdSbY
R7jUdFkj8ZG8YzQnk6/aFWgqVtdr3XPUeGmr5vSzKUT99FTvry978wazuQTRT2zm
npZtwyUESgB3sxc1LrIjbhQZIo6Gf2Y/D4NRSIUQ98+GySni+WtFry3PKOpzZOYh
rlgKeuXov1+R7bb0SXKmkA40DdQ5zxU8qvmyeMFK32tiKi2MCb6nD5BXo3pfBvaw
/yQGJAkmzeWcpP5j+rlaF1qUq35Oyt+uDBtDsiU1NtPo1FoqQoQRkJJDqYS66hF1
4GpwPuf5/wyzIyN2xzAHK0YKgDXD36r0lPNHWw+Ufmtria23Pnji3yTt/O0H1E1N
cvyjyfcsvmtnmcAxD5ju38NQ9OAMolAHysBEoeNArrzy5GEfD0IiIV3GlC0mPvwv
dY3RFEAWClxFuodJuzhWZgjnvKBsEAFTKCH++th3f3LMkoZ9o+/ZGDZoJPMg7+/B
yxAaedmXLZnIf4MgLZzw6Qi8/1oAJJutO0dNVUgiASY5//4I/M9FgcMzMo4oTjI0
JKHDcRelp34isIdO06Ebh0bUHbiybcwJfHSKFNlzqR40/J80XDtAYcxLj2KjzwNU
pwoQvsyvojYGzapySQ1F2mpj78jLqpfw8Uc8RCigQ3pWtMIV2mY2A60ZK0XPxkim
`protect END_PROTECTED
