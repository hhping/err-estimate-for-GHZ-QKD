`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q97x5rRMSt9kG9m+waIB0Wzl9sY559pX/8tynmIW4bJfVXbuU4p4B46dy+Wj7Jn/
Ea1ZKfsfhNNad8qwXekchtCbBazrqfbyyvgIGOmURZ8U4exbe3RfzNxLU3WdTWUz
DNDTABcYRFQ1WDCjZTTAff54jy2WdwfEX01KDcHhcUKYBeTBTUxGRxHJ4XaWJK3B
Oc11lkkbplFfP6stLksQVaWk/e5tvCXHnQ+i+5T2vvK/ySZ7qvQ53qslqljru054
Mky1EbbcEJG3ebVouxdn7bprDtrvSHgUAtUyQvCQMm88tgO7Df7TwUm00W4TZwL9
HpuaO5AA8bcigAdQL7q4hs6bfIu6aWY7A4CCMmcK6Mx1SR2af4bbXgmgxrwYR4ht
5Yrn5+8q0o9vd5OtxFvWP8G7ZHlTxWSmX61DG7S+te7SGTJCyC1bp/IJzv1sWtIO
UUiAnNkFUwMMFWAJ633fLCpphLrqHtaekRo/0DgGEakF8cFEfN+BfgNFWvmtU0RF
U2k2paIwbG76m7Gapss387w7k55gKvMfIwq+ETGhatH68bWa63eFOLLKRTA9MnBf
YrifefkWbGpfvxwD125fGhsM4amu3gjEazEedDCB3WOM3sWkxEN3b1HD6GWYxz9z
9oI1bbTpyhRkC8TrZGotqOJS9j6xo55lilrGLEK/KNOzqhhFWxiwP8al5aXVOhu1
pAyhFpat/+mzRGVcGx7FR/Yclo79rjsFqLM8dAS/CAVMherlxrKln90QyEJb5T+J
aI/BBvLbWTLPpCE9wp8q/+WdsTdf0B9X2uzAJi+Ki1MGsst4vTbgcLc+iykyctk7
sfPG6Mkky0tw9329EO0yqMWyeC1Gyp9Gjzwqv6KWL7lhnPmHm/bCIJ1A7hgeEjKE
rstBubfbLINJ0yrkU2FoqCfY+pJF2wZ33Fv4Nqj17aTCTHpeitXI7UyYhZUt6Zmt
1iu9Kn7Y4BvE1qAlL1vaBkZ9nurvrtqqMQitRLljyoHyD5HEEnFuu+vKSiM6FnX4
U6H+seDzKMYPQ3gtpBQmiYdU0C0MCJPA2X3v8VV5oysnSX5Uwn7y/aDx4D9L1dyN
Gwu5Qd++4kAACKOSejMRQKWBu6+HtLEFLe/dHHw69l+Dvi/6c1ekxlDUN7PlScpo
ZRkb2DUHVPIWOVlEqSUG1uYrxznSbM2wC/g9UqSp24BJon99quLfDFDW+iq913r5
HOMBj1Mx6qGaRPELXBtxAUUuWUNifQe8LdQI+bWquKNhJS6uRL82HLBPK64Pux8g
9i0diapXEUZFDSf6RiUoNdAq+MLBZ2a+xW02ELl1eRyCB2oQX7IXTO3aSD5SEA+k
7g5Jz8GvrFe/8Jgz6MxOo/squqRua1j/JoJJNmak3C7kHvNVneF0bLr+5KUoxrUC
evMpqbtr1OM5h8p6rJCAf8mn/ZsxGf+L5E1K1zHtH8iAVai0uOlbicW1iUasPLfL
aYsheFSmHfAaYTee0KRUS6APd+SAmJJvX2nBRrIhgsEP2dZxFbuINjhhoSZgo4ZF
WsqZJiUPMApkUyEqHGcddBQaNcUlyRVjqU2ZelYqEaSZLK7XhROERLzIyJSuL+MP
AR/voVqWp+sdAdAc8B9K1HLEurXqGeEXH92LW33ZNSN2LLzjwqRnO7MMpTNWf7SK
TNfZbKbLeTyq51zlQnUIYB/Mcn4D+9s/pqjvvtrD9QlCN78UBAxAShullJJutPDE
6QRjPeODb2uFdUYlWsm/lTiaRMsXHMAVKjO8zAPGBtOgHKm1mCq4oF+y8m2UcNp3
WW/bpL9p0TRkBlBn2yjmtGhsnFjGp/Ez872emOyy7TihZs6G37yJiSd3uBRkLj9J
0AwP1sUILfwEJVhXXCRiw3AheQ2Pw4vmUfCdHJAmwtlXiYNMSj9DGBxEtlsY9lnk
5fVryqd1VMbw6M3awxpHP3fhf/LqCM7Iramkm6MqeDXZRehHKZ/D28tiw62Q8XyQ
822XaJnxjhehe8Jy4EEo+pbMgnW2i2RJQbYkfjVZSV3lUzBMcqXKoayPcEjM593C
8FZExKiBpri+kpWfAW7+f3EUbFCD3ZALW1EVhTLn0Fyv0foeCrbPoL8+TYT8kvuO
mYe3xjCN7czFgBmhgRdxbd142hFZTo5pHh6SMRUoLIBnTCHvC5Apua3QY8+3e80z
ZcC98VavNJ1p5jJ9Q4uAFJWr1XzQmrkUsYPW8ZPSyOrHluN3rE1/PaBl+bn/hlQY
9Aj0ON+5CViAfjx4vqmPZbXMOu4jCDxKYTp1xfEsq2C4kzWZSe5qZ5rHcH67dKM4
OI4C2bVCrG4deXKjbPaGcFYqP9uFBTIwLc5OloQt2RHV9zPkOE9nr2JC7lKNcr0S
IBjzhNlb8I6ygaMwrs5vQ1AewI2qb7C+rQgqsuuT/CfzNFge30SeRiquvaFQ1vEo
wJa7RiStRmx2X90LZ0EBCRb66FjSeUBjIYR5ehFgRciRsyktPiKggyFhDTwS/Dgx
mOVCqzn5QVBuwRc8AkN+MnlGI9k0BAXyh369Wp1YDAAQtfEok07BWkpv5jpMUOTQ
JHThXQDS5uPO5icCeu/tluv4dZFjmV6n0nVXodwF80DDNY8Juw3KBBWaemFNuGKi
4rf0Rx6ums5dToq3WhE6aiS5HFIfw9Iy+DhvhLLydEbeyQ1OwtMNF8n5V8uOqsvA
RFQXYce7V4G02u4X1wAe+XGlgyjLqfsB0b+XfNTHqE4aRfyXFIt+Nc/ow9MsstCm
zxSx5oBXm7fu/6kERCxb7WzdFYHqje8/I+UDanB+tEu2cjhDTnsMlwXlUrFYiySV
L7WUlCq/Z+OLR2OvGJshd0gs9wrK7XAGbnSh+sgUMEpNFxKthHkiT6sRyI5dGqp1
LwE0sR8f5oee8G49DGlvbfvY+IoscNUOuqiyERF2ybAfhKMgMa9XWb+BmJW5Yk6v
6Qh15760cpQbHa+mSAK0Z39BHGegpKdxv96SnbHDvzs/xuUIDQVO/jedWOKibyjA
amQq9I+ZsGYnE2xBatmJw6zPt6RqxBYa7wpFGEl51IeftxuOglJi8VqHHf7jc5KT
/ZJ+saezAkEaZpFIblGRgTzGcIphL0I4mFcpphuPXsYJuvsbSj/4AYRsJKe6/lAO
tx/Us12zN05+CzujPzt3UKNc6mueg51BLvr6e/84P1bchhhoIlXUifAje8VXkMOy
L4/HcjRB10iUjzWlR+5me+0Hnv6y5Q8vXpzV3MYKWZGOIDIc0VOD4Dvv2QGH7qb4
OEnFhGNypMoZBtIxQZrJ8UHszeQnxIlWwg/sGQx9Uvnse2aElShDIQPE6ufJkM7W
hlXXGvxSdo2Gaqpa6e40V+H9NBdt4JI4zQE/5FDfigG63yK2V5Vj8NwkUdHIeYTU
YtAqXmwnpYaL8GfnkTgHx5zYZGJV8nVtpxExdU5EzlrGQT291UidHCBuGQtRjFHp
8Cn9MG+n371kxr0NiYrrPDnnznRNeC/SBAVkwH+nAoIuVtcAVRGB9OkyT3oK129H
57YeJ3hvu+efaL6fcwPNoyNgD0j3UdoTgoCCwF0owp+DGFzHXWy5uS7+4X4tFEfB
j8T6FBQRUQklQJWjOSiyVgiAjyd2HY7BtZexZyx9G5+gCJQ3cF+MIy4Zd3NpZowk
emUOnZQKZLzuQ0Y/pXZ6jykAEQtown1SeL7QEZdb2HgVrD7/Z+gRy1Vh0vVMH1YQ
ce58NPVVequ5WvuHz9XTMHJnWleeVT/ZM1gDSRRsJjJZYnE62+0SoOG7kcVbsu9u
L/n/3NRKY96ON69FitQwTTXdIdgkZgK7OE2leoR772r8DjZpqTzVnR0v4AajuIIk
tO5e73MVZmooKgZ3XQZ1xl793p4I+GbuJIxfONg3sQYXpNojzktRmg3OPAcMOa8m
jblqZZix6TbSbnnvIPvg53/7n7D2wi4vbm5zZBNWqrT0BjtNUkFXek4xmtkr3ea+
q6azFGWffX6DMDdWWkAvUpEzXzE3he6Yzy0lhRd3xr4PcvLthOBkUnDgOl1l+L8o
InxrpnSK8lOczWJZYXVAWq5x3wdlKLbwcsLg1MV8F2l0pvXGblP2XYIFgm36HiVD
PedOvHbxdTew8qp1HUWQjXvHjMHL78VwRHBCq6qW2MKGDYCRLGMVmV6dyAxtutgM
zzx+6wBnZaXvpRdcgu5RaomMZ+nvd7YCbj8LSKrXyvq/F1H7zT99Li6ctQUTaIGq
9Np3gdezwn8mNjUDNeBmhnL41WIAF39fPA7Cfy/V74q/7FkYWgJPL4olcJzzO3nO
h59AZWBGMtcrq3TrIJUOKdXQ7dbZ2dzQ99GEnKw5/Gpl8TYJrLyMJnIeMeqA9Uav
Bm+kGEYDiK1ktQBZRpZpnptjVktz9Lz0iloJ4Q3AbALeEMaqUGo9aiu7D4y0BwAM
AcjmGEs6nmOanXW5o45No6fX441lf5H6G8EwokzLZbyvEWNTSgbjSlQvAeTAE5qb
onZQlLEZTSh9wLZm866LoaX7o3mI5gUDusXM3oDu5JFj2HiEBOK0rks+CB34ZX/Z
LzqH9v6V3Z1YPe3WgzyrUVH/5jAZJGqPMmKczfFHjQDL3bZEi+tR5AudRhb6FJWv
f8Xur/IFY7Z2PCaE9vpbZaFlRthw78d8cfRf2StAqtL2Ika66dbRPt89RwGzvk3t
DMgm6R2CBWN/0Z9iFJrWWTaF2UYVr8Jy8M0k6ZftrG9oHZztSlc/vOiozGWVOmw/
38Svnx843N+zQTtMIrvEMgTh9vOTlSJYvqysGdbvrTQJvPBiggP2RO7wKG16EBCr
NhWipIhKCsSTZyz8mXyUeEwH8VcP5g09hxhd2g0T/o2GAv+cymi7VEqCAewXNNw9
0AybQW01IwUOSSYo0m9Wp7EUUAnRh6j4ZiDmyBx14uz9Z+q+HyHGUqIdUjgsBWRn
wgPabJzcWSvzoM0n3vgWsrDPvt/Ev5C+PoItyOynsLLwK3vfpimD1kxiVz+Nu2po
Rm2K1iOlkOiGKXmz+TJvHuqQwPqwf5cmTnkcaAyWZrRmgwP1fJUJClOryXbevEpD
8gWqDTc4TmZdz+bKRhC5IKhleApij8yjERYDs8lY3KEDpSO33+OPrFsigmWWqLei
P++SdFmOQ6UoiBckRjBNaV/ZUJnSjXurIwS1whOwDammUBIthhp0W/4LEDcT34/s
TEQYvwEM0V163hje4SqdirzPjbgQksRA+7XQ55eBK9GEJMFHhIUpb14HzuQAycB0
a5lxF5ObXPT5yKZvAspYDlDCDaqclwZMxvdZcGGqY/JEvksjMVE+ClkqLjHkSm8Z
ygISgb3eQMJu/uf2iEZWW7LSC+K6rJ65UnIO24sh6UkC+mp9WIJVnKhH1IRnEhay
SzK9cl0MzTo1uqp6Mam8XRVfqvJvayi4hk78kR1qNn1noCrhH3APoZlGDCdlTIQp
WvkpEKQW2Hve+HhVh8Js7SrUgOftQvtiTRALeSzF7W8VulSH9cjOjaIUbPYaI/3m
YTSeKm2j08ix/vANyMXRxrH0MqTbdOtEJjrS4qhUwpM2Uqb4REgs/h/nm9Eg4sIs
NkA6RjgRAzaPkge50MVidBWm2SoBzNyExlTURq8FZrl3HDr9Cim7Lo7f/MnfbfO0
YIM/AGYHojmA0+u1F0TfMN2V3ZR3aO8mPhZCUArA00ARemceTeigeyzQSeRghUe+
kkEmGb9e574fdhdyMjp7DjAqpTcPn9agU93A4AIcWHnWmR6RdEPgTWTA63CcbDzo
6DVhSKtJqKmx85KtJaSoVRzGmuv8a4mW5RQstncXkJ99a9FmQRyV2iRFT/MjlXPY
xD7r/iuJ+XGHowpfjG538TXg7oDZ5rzvBX8sPW5ljyvF83bQ6Ey7XCtOu+3uWQNG
NJppsFQBQGkG+SO6y7vVno4ryDKi5j2t/SSs+HsYIuct8TOnwJ3zW7Ek6seDFsa+
02q6WNNF7MQJpz22A0u7eZyD9yQjBfAcBntAK/u/wnijJtv4gcfodgI3QzeQ5/h3
CTrGeugKwYssPiKq6i8VBCjAOM8rOSTSXfKqV0EAAFtWADnSqHfB7/VBybaKem0m
/gDoztprdh/oNG0ChJPn0BQKEmMrFsjNWxIWTc5EzjTagvWzfOLT5rziqtqDzmME
f6s353atcEAKxV9PiRu7sm/8cDfJ1K7WT8mcI2ZjeurcqswJEDi2bgsroiCm48rM
za85tgsGDI1xxBWyucVPW/zMj6gB2D7ud+G/g7gg7Tm8fM2KekA5YpnlhGUyf8KI
CFUVz4yvnN28kFpREZMqCcPas75vGunyhElf00RADeJ1SZSOSYacymrgWSHqMNgi
hN74wvH7b0d1qDYe9PbNjGdsRmcw+2stbD+J7+N77LuCCuxS+BltXiI0CfChQBuP
YevxbhEdIMQS562dlfaemw05Ctgk0ToWgByhJCjF9ydK5Oev4VgJg+KW4HCk88/F
6TYdOL8qFg1GSeS/NwUC59u+EAs5B0T2RAHvO5jxlB6aQVBudO2lpC/dZEX96lDl
5U5wAM7B0c2VnjsCOE3OcanNkpDrzFSJHIN5U74XwwhuhfjhFlFOrzeDTB0QoO2M
3cKL+ycVjcLLqXEX6ejGMNGwSJ8gCGKBuYgjhHcEv/OdoylV5aqD9/C7z27Dx6ci
MrsiXeluDWlfyZ9DAez5F83TJYW9H2xryT2FCYt3hSY+cYgSXPwbREtxk72iSoOa
iwoBgt1QeMA935aMIHWGXhS2OfpsaeznRhKa7hv8gXO9OSA13H1UfUCDtKgHDPyN
U8umFM/Gr3xI76eyK1fehBUDvmFCWJiUnVMViTio/YMqzLdTZfxMa9yGipTq8zbR
zhxz7/8VoJIUDqyeDwIWr+jUF8Z3qhW7yqE1Wk2/v6QXddNPVhpPip+SgV07Dq1Z
NkyL94xXTEUBcYa1CyOvnLWgcpK5kxzf7588Q/CkDmcaf0dh8BWnrgO7JrOnr4Ib
Nu35NWSXNjQx3VdDyMWvwNdApHd4IkexDARAvbD1EQ+EcLvFwSDt25FTBCwhPQv8
V/dMkbUzF9s7biHVK78Tsi0Wy/Yj6fu2xuVA792khT/GXWjvOYqnkkzBHS9qt4Bm
ihlzN8YBYQ9pYZD/2LnIK8ov6fVhPhCybuld6dkiyzbcquXNofd4SSFM7HPovufW
cTr9BKuHCrQx6xAMFVhVCVxNc4IxQJFkPM1lHEUee2OdP26m4QdK00ITV9X+yvYA
P07LAJlMn/78wb1gmeTWWXeLcs4B1+9PNvsF85yGJokXqx829wi9op6xzLkIfgDD
L31MyUmpXoQTZkU1ACp8CDPHQ7SILEy2NiThoij+UQEJX6MqScJDjAYG/NdO6zDE
kmULKsGt2ovtQYjFqMo+plXdNzpStHsEO9fGOgpi6RDLQdZ1v2qh+Hlk6A0Rh+Ks
tErh2SH0BnJ4d+6RW6b9E2Vxonj7zPIATaRj1A0ruj2cAY0U/SJAKpoxDrp183yB
G81hGQjskQrytHy/dTzwi3TMSYGENqx7a3bdWf9Z5KQLyCxF/Qisg7Q4F02lEL14
laE03TWnpMoOHBoVBF+1IEkktBBiTbeQSx4xm20bXdTkvcLSFviUAcnCKzKNi0oc
nyasBuPkTNZsW2fP66gOO0To9x11djhYkxpVJTk07RT+CvCGQOjTahl8XfUoX/3M
mwZYig1RUL1p1yqDGFicU5CWN+lBlWhSN6N75uj9lCP711985usxlvCwmemoDqCz
q/gNx1CMahVHCIEZmarOqLrkl6TWUuQs0sGq9YN4JeGLL/r1FFiiualfCD3dT4+o
pyyT4ZTFDy10PdAUpkWlG0DOPZjX2sS7HHUzk4tnDIhiPGGx/faYRutvfEfS8iFG
ZblmkWtLUL43F2HDUzuvkQjnX1DzW0nCM4AVEjrsLs6LUmfL4dX4hAnhuXeV3Gc7
xEDd8kq386x/Edv+fvyRzu9KpKAUor+MB3N13MbONx8QeJBrNLUrra/yVhv+PE3z
1+skQRGzkJWPi69gd4ciEdB6ZEFsaLJxKHJbTulD6s+mlBT2s2hBFiuZuWtnsYk1
9LDylL2jGQBlEKlUgCHf5gUA9xZomOoGnW2KD2BXwVPCu0suVouoPa4Iqqf5g0vf
ggpCjvaSQruoCupEb7o9ujP3bEFGg4EuYQWIPADNMyg5lB4puHugE+CqjMsQu1HO
fuIzF8MDbRfReJSeWyaPNybRAwJuvKMWjVbj9rqdM+HOBy2hqJk2NgQQ1OJAh/xD
pe/88dqw/Tfcx1vhO6Ll+gXYEz6V30f+AzubNb8uPgwTRjQproDjJjR3/EGxInFV
GYQYY4Noz+eMy1GJPLstePEwK+J29FdW+z3mQ/13/+GwjzcP6bjbvZkwf7HVpcXw
R5Yja2imO8QcZHYv9dOJJc+9CT52SkMPjblq0s0TTLkRTZEgSojeklMpTo5ywVaE
OkOVIdr56AQVyd6sm6mhi75Ohd4HEjLxO0lluZVAAjAwJlp1YWCjdvYGiicUTwFB
C3H2o3Fq9nm/AZQo3OZQ7BOoq7ZM0dAEY/Wv2OuBTvtiXRs3AFc6zk+FIvgU6EI1
LH0i804YcNdEWgOdwn5//bUSPfJw/nxLeImAlp5NZHd+zeVyVEx2Xqih18W+Mevm
jkZUIoho0xfAn0vx6FAu67J21ZCDd2+N3EqhrwXOoX8i9PIqTydNKecABlU2MUPr
xQ+3yjpnIez3v2cV09DPu/T9wMgcA7wu5jJc7N/WM8rmj0/iZ0JMqfafmXSW9ugr
Fu8Nzm/NgMh/CmJoeL6jGBz5gyolnA6e04XNeL8IO8C3zzDjb+XEj3ghIz11q7nW
PaFyZiy8vo688767qi6JcFCWmuI6jYAWFwibcnyXP495dyR+ddbPWBUuPhFqvAxf
6kqSr9zzfEwXe8t0cLi/medi0T0N2g7iejbmPZ0QvVaSquE5t0juXiK2RINvV8zE
INMxRVtX+QayINdaOYputE7Kg2IMgbiipREYknWxnyskj+uGWpkpUSmOsWJ7iFeD
zklbzb5d40Bym3slwk5/ySYTs8e2d5abajsTzCet5PaX2mXApLHlsnTEBipW+NHH
7o2bQQ5zKyJ/KP2dRWJc1hfpGSU87ZQuXRKC3LB7dEPI4n7cvwVl3sIvCWoTZnFt
0iSPruujLCmjO9SQg2kBcEJSnJ9S/lauK3/s8Y30X17BiB4nhQ0ce9jogKs9xWNH
OQye/mjFiBWtP+Lv8Brw+B7b+ksHKRA7Uj6JKfG8PlNZBAgVu/2g2WZT+xtdLqHc
CPIFgN3D5suoWpRXAGNhT//RqxLFJmgF4ZONoXTY/5WJ5VXpdY0ADTLa5kwtWxSW
RnAjKTeWO68DStzj9Hz0NpKtPxSZ9TTtIHGGCQlUg6BicKRlLBHSepbI1QqT/Hd0
Qh48NJnbDbQOhh7AB23ewQk4KeedjkzLGgDrOA+ILjfXUknHtY4rLNs6ZJev0ciT
+mxkgse3BjWNIlKbVuYnQP9YaGJY7TnTx1yEzBkcb9F4enHBJNybLllQzjKwoNW+
L3pr5Wu/pYe/vx5VVdpR79FMDsCE3i1g6gQY02WmRBM78/v09p25zbDIjD29rMgd
XzKGnDfG4o+TOUBNpBXrEHj8BJbxQcIToDiP0TMcktCrTKJJhRw6Lm1VG3jwrs18
xuLWHO/lKYfZ6n/rq2NP/la65vsKBJ6FDbl6vXbVjjXL2MPa+ybH/qiHaEstZzKC
piPXyDozKrBxR7S7LAXKdZ0NuaiJCQm51dzRxUu9hL7xMXUrDOaAh5Gt167Ha+0T
ncbEpPchs/r11wRRvhHwf3yGmi3an6/YWaRWg2JzTWLuoe8cVLRL3S2iv8mX99fJ
VOH3Ybuj+PtR8+bryaTT8/+JxPsmUwW2RtLzFjEl1gqqb2DtDC+DjuDF3deSQXA1
xsbXiH4mdbAaoTWNNFSsEyu95ub2hywaa2CS3jIOPZDsRWJ9++gVTK36j0Zuazts
pD+mOMF9Q9S+pR9+Og9nUCY5ZIMfLAJbrRWDSA2xWPOBfSi1HSjFpqPebeHbSh/2
195c0R9P1Sb+sLYC5KnDDW4F4mJE8sHaHP6l7AeuJRyBQ7wROLp3VnJwSY5GkfOX
SF1F9Q6icS3e0qLQvJbhzMcfT7tQSdAaZk64wxrh+cPwKWAOTNGC8h5f7AzzSVKT
uyhnDbNSaLDGKjkjiGoavq7/pFzwEVhHSWJjuadMAPA699hX8N8XkGshW/MacYd4
DR4KL+Bn6F2vYe+W50/RhR9tMzAUGg/m0QdQhD52VkiWqrLiQKwrMXuoJdeO3KJt
TdBfZjxiQF4RH160ch5pX8gCP6x9E1Z1bJpqiVDUXJH99UyKWfPlx4TaUowBcWIA
Kr/u0au0tuEYpODXHecJ3vMfIWM2GiGuU0Ggxjt5OvcpOZSk+wAj7vtARunLuzfH
lYHC6RuxKizz+mNNIdLn74eNjwU6YBOLCC/HKonDmEuvwUFfzxKaJggPAipIvxxq
d2Z4K9ozksbWeVrNhXpxqKw1oYXxJIjzqL224tZLi8KrBDAO3B88hruggutMTpOP
IhMIRgDkRec+3FLy3UxWt5J5da70J6b5agBL4gTO0twfdB996r/UDOAR6bKRT9lc
CO2xbDiflRqaeYBpt93eF6Oo2wUGyU1WD2fHLtA3PbCmmHd99dfbiQJ6LvlPfSd2
xFuY4MP2mw9QgXCrRWsYsAD1h5+ay35MvCH/rXqrZHrtXGKiytVPLRgN07AetI5t
d9dPVyE82Hx7k/A/pel/knaMVxGK83bMn6v7jJ6eMEgzDtGIKE6gqYzD1497zGls
oQSVYinhIS/i0cP7TCSnKHQFPPzTCfePnWrYTIBs0kFNOaVX/PwkXJIhn0sUPJHj
dpaEu0FM1rZ93dTeElGHV9xywURl388seiWsrKwk4NfttRpj9i/mq13TDprKMKYk
dfnajpVCNFo1Apnyo/BEgmxXaVHEiTy+eC+xs5+c/uvUjqPmHeqIWsnSR2A8EOhE
M3fGXtpFEu7GJIKfaX5XfngFCsKAJqZSPQ/ZNloJrMlCOWAaHFXm1DTWVg2bGUFX
X7//zkf6fNpDg66/QfnlqNYjgUMLUGdnh6bIE4hEMTlw9K6j+iyqxI+ySiYMaYi2
XCZg3QyLMQGiD97UslW7WqwSHF/PjWouSIxgDshI0QLmQWaFdC53kVY8CBe3tD6L
FOG/FJCC2fch0Hb4q87buIYX382Bv7/v6zjwzVWhX1/tsuM/l2s9nXcpZznmensz
banM9px6kHWP1gOyqFf/rBpn3BF4jGS41ye45rBU4lK2ZB8QR7sDxFtdBJm/+Edd
DddaJ7XRltsFGNuPaZCJHk3NuzgViNVcUEUtobEUXJ0+4wn+uRR7vNJ3O6ZFXtDc
vSzC6tvhnSzuzwdMVzI0mfFvip3hObvAUoFRVOcY4jVq+tuQOdZBi4JWK0QhQSi1
S5XqdanJE+pfCQL8OYBLigSt1A6J+CbjNYHPBftRp2B1U7KvloyrAb+afejC2cPe
szAFmcnsSm1mILokKwkecRqP4t1+mwrnv/SFtMZ8rLaJ9wsQS+tISRJ3P4keDIOB
EwSdYeTFS/penpUklF6TOlkXcJnf8YjgX6jsV+kyAxYbZwSAQzJ9UV2ZO314tmUU
sIPSmAPNU/cGBSCZKyg79fiO9SgQnQkJcBFESoTG8wvpDWlb3igjQg7+dFAWw7E2
01C0UPtlqOY7cLXxneTJtrxFHEOUFxVjKjQBNs9yPvftO9Y9Qvat/GzYCgjlw2K2
65RnX239DXtG619KJh4PycKBpl89HLW7qzdoPp+GdhSZogZoSWCLOX0G5o3pPWsg
W6bL6Sl+O62QHxJt4cPnTuqZnECU7gVa+OECwduPHA9Kh6TCaCvXRfHSafOJKU8w
ZwSwkJ01BhSA8fvqoGH/oE5jIHQKFMuoNAtQ9JraloJbO6s0TJqYIFKDqbMFujDK
/2Qpi+ZwRVjDGKpMKw/aYLgnWq2YlCOzbFiIXTGEMrvvXNwrMrejvNMqNLlhdCNA
A/Vt11ufhNiZy8W+0TD4OLCf+05aDGjGkxYrPASWFojilbqBMjp8GGPZ5lDterqT
AaHqSINBcom3A1XtKXcm1WLjj27V19lZFeEnZeTUrhPeE2Kkzk7SKHjEhSWgpEK/
Pp95YlE4YdW6gzKZqzxA0Ydm6uR27QUuomCgJqPBUaHvm5Qm4FUZQLOTjEIR0+6b
yj5qjRInzA2j+BdpwYbvjMBgEoVnT30BK3YZyl6uB8/fhPWV1Rik4g/bEKAkfbm0
kGvFUniy7EQtY+ND2uQvLwexnJI8YIxoofHwEw7ezFDsQwmkzkkKo2p9iDgUA2h7
wSdwfx95w85KDGJysoZs3jz61XxJyqU6c1DPJwnu67IxSuDHN27NIBxL5z5I+lXJ
OSCC8nM3hD5mrr9iSuH50Pjzp0ZF/NqcVe8kFlTBM6J69Go3vVtzRTXL4Q5IAE+a
9YhQa+/PebX9MG1+E/Wr4ioNPr2Y/30VzXdOFwFA2KkX7k20yo0tRicBo1nBABMy
BNILtpZ8BpRmEBcrQ1DVaCxJSYL/fG5nB/525qU5yr2MxedUUBdy8Mrw3zoYcR42
k3SuUMnFowT2BHTlDSMiP8IVRAx00RNZOLIBrKB5Ey3wvrV7UJX0VtJwfmIyhzTv
5q9rFwUQP7mbMWhbmWwMUnqr/WT8bFmhapQjMTXBSsflPhYuqAlLTP0XuMKNkWmn
MtLIYwZpBO5fzwP2WQ1MTgjZoUE9Cp5BrqAL38C4+g7MlAg64zeLnjHJ6NNHmkGn
vPyOoxv7BDXsPl0UyAVh3xQyhH98l9pJzfOxobbp26UbnRUNVV1TFIAqOrL4+LU8
ErKkGMU1aPeitos5dI2h84hcTV+zsWlO7rMyyDWlxxk0XdG+w41Pq8KuiNTSrwej
dv7ltsf3LJVJelKjqO7FjhSCtYe1p0DjQLTb11O6MIWbuax3KFDuYkg7uHJv9gxG
PgVQCfElntPrwKsDRRxJN4WhlXgOOOng1AoAepQWbT+bkBmQBOdXIhmXFfehvq/4
yF59YlZrAqsgoNPLYUyCIDc/Xcm8smQnHbHoIE184iJtwEa0LGUJDPLXlYEzhe3S
4OvYN/crUIcOdaSGqJFibiPsBk9ArUe6TEmsIQiTXV6e87TcrXKRAEDLEbiX7yYP
HLbQwOyGHWl4ie00EZ0zcE2rcyOvSGg11FjYNfB5RXgHK8Li4AQl/EXwOTyATuAR
UjEw3hnQF2TMFK4tyy0UQGWVLV6m3Brr7V0aonvr/TKmyX6H51Awdi/Rgt3PTt8h
k1XNLDniWJTM2yW2vGr03MBf8DwWl20PVDlrcOdNIgvVSuLoVmqgtajGYGafQW09
qCJ8Vs+lm4A6bYE+xm7yV7smfm+IG8an4dVVndMdgWX+P3AKm8r8SW05BtOgpnd+
TYkZy1DgDRHLK2eDpagCFC+xZYDAY2F9cbdPPwWxRjpscR8RA0Rns5084nmGcKms
h4YJJ8ZXQnCIzzSlOWE9U9/MOtVhRB0CfPc//r1ll0+1noDBiPoOs6MZvLI2cgIt
aFggbehcYJS/20loBeV4chvweEIzTQYEBWqbJsE352c9lrJAl4xgOcoqz7b3FPUU
9xzPsci0FbLnVuw632oeKE7Xkd9n4CC0CPGGJkSul2xpS5r60gU8+DwwerRk26vw
luYvCRuUPtAGsaegQrbyoxZquaG2oLBx4H0SdfPfoy8+cU7DkENrlNTN5rffSQZv
kd1pr6CcR1fway2vB67Rk+36w6qqylb0FRT67120SRlRQRTKJ8B3wLyreJnwyUPf
DooXlmSNzcnIukkrPYswyAoukmD8ocLVMnGeUNBNR/tmCegtQeOd1LqAZN3GPvsM
H4ypTTF9myOoMlTK7jboCpBOrcbTNkHVPh1FW3T+PU2jZkk9+9CWlzYnheooqL6X
wPHSHqZ1Tp5L6zZ7YJrbgx4u8R0OYkzM6tkcbY/ytmz6Gw+wUVDFARwtxWfe4UiY
YNliGhqwVOfmKbVE7i5FJ+CWQWNKB5yL9trMPlNpFNLiDd945W8r26Pt9uaH3RtT
onGA32rqvJvBr6eQDTefQl6BQW4+9wb5C6w6TSMjxSNueiacTPkWAQR6+Ymzq19g
EiPRPuydWX5jxiBdMG2nTe+mVTGDRa2FeXBMfVuk92LGbGn8oO0d6Ck0e+fc/Pt1
/qn+YZAOkjJvHVtsSuosqe71ccf4tc/IZh7eIE1Wpes3D5IxwqgcDzw8WiKJDijR
76ZIUgt8EDErCgiyHSw3nvflGCV5rbVEO7wVNdngNXGC8Qm0Di3cx9unCEU7i8Au
obQ0728s+0TDZGgxfDrnsUKjYkLZ8eeArVFMF4JwKX3NjvcgO89wlMLQ1YX4VV4B
qrpy7zEDSidkOyL8G0+h/qM4CdOZStTIyad4EArC1i4VnNMeSrytkhzzDLwURZX9
w65Ulqj0ro79Gw+1bUYb96g18YIXhwaRnk4qhyXCbgIIDBWx3thDZrJsLBDt6cnb
MG0BK1XOqLUiy0XaOXtDKcsmUDHm0Leh6RmSkik5qlqWIwmqhWkrZNJMmOChAy16
W0Li/g/zE/coNHU9uMFklUlWb2Ur5Umtg480w142UiSH9BJAwt8C0X0C/LnOZXlF
XiycWnA9BdGIHa55zDTh4Hovn76bZDX+Xy7btZ2O050Le0PVjjv151fR0SdOftf8
xpmzCg/ag1LFzHpA4VoFqSw9nDx26EX6yukol6wRlhbRDMNXZRlTVjjJ0LLybsho
OGPjR7L1v4E76gIr6PYDQ+91IO5aKfsXUeTMy5MQCbirNUVTuYDVg1auC8FalMck
W4XUdzxTlknHMAyX8pjfKI1cWT65kRKqh6Vt9U1B/uPjxRA9EnbveZ3p78RFA7mp
lM5pTHG3wgz3+W4rrFWLeQYZLqwoKw7Bz6PQzTUDwcv368wyU07d0uL1RrNnFHEx
QRCKqsf0yLJvJLR3LOT+FWokprf9b3C2wmmSiojMXYUvnvpNbcyGj9jDtqYYTJEt
E0wokXNo/L8XzRMYTB0quf1gc4xgrf6WYJi+WWSNwvteC3rIumxqgKEtOF/i2oMm
6WLx7PCw+RfrGZ9ecC2Q9VWcFGoqmoG1A6A/OJ3n2HTctLPIutvRwPUiiE0eNO8A
dKcKHsj98M4w359djtrgqFsO2Xz8eW1wbGkiKw6xEov8As1xHWbhGzX+9JSAYZl1
uXg1RRvb+WXvIpRpWm9yjz9oJQ1c+w6hN/681vM91D3uy7vHjNlQSF08N+D7/+Kp
oXjlb76M4PjJdXR7HSZ31GZkCYIzTur5BgSWD90F6X37O4Rmp5ND4MIpFF838f+o
kwHMCArZBmN4ArK+hx8hqRQPmmWWsrhOxqRh3g4tLGtq3TMn5K+jX4263RQ/u4+B
tqqZ/kRCasM7CjnwZO/ges5D3fhYpiFIZCxufGXWBkVJxImVphD7QDpBkeFtshNq
QWoV3au1gbpqo6v9H9EY4IGebuWGtBGh1cPLN9sxga2w97NAJ7ruHgUj5Ad6mZeO
e4hdxa0TLqhtOCduPs98Dzl3ss/PI42uojh9KTT3neO0yy7FUe+wJwBs4nu4B6Y3
tJ03p4qaAQMobpcCgoQR0Hku8ppSddBu0XRWMP+J8RNofIYVmH9fF2U4S4miPmzm
lYiZTIznU5B8Gix7WaHc10PUN0gX3dz/IjhqIg9SQxZr6pmvHe8UD6hSYS+iCqa0
6N3VRTkLHmpacv6RHZYxNj/13T7+jo6+iPLVGWJDPwf7wLYyIUY51TlOPCbB97W4
KTzPsotTZQvoP1Nyckl91Edtp2APu53IOd+i4je0Mx4x2OrA/F8VfQ43F0YQFugH
lVXfC/pE8AcGoBE/jC3LEQRAMUwm8bSJGhmSKB0KDLO4LcqQ7wqvtwZ+duV1p7Hu
0RLmhs9Gp0Sn12cO1/lZcZmarK8aL8JYqwv2Xm85c4ieeRYW+7yx/FvAPv13i/xF
dKagSw2fSOZS1TRepgWMUmdTjPFuJ+ABkJJTPFXw2pYEQpoMoT/dZ0ZJzkF/L/H7
0nbGhHMmWITFR546SI+qex0nNetqQUt+sCQfnyxy6nd08crzJp9JkfP4XcxHK+gx
kDIY0dOKHph/ErqM9v0cn9xqrFHnqyp6PySPHxTzaN3cYLpYGgCGDAVv0oTjNnKX
LMGG36Ft1/n8v9hv26RMBqsAx52m2Na/b7wjzijvO5KY+WVBFDWMG1YHompC3gyf
XDezCfHIJ/U379qcPtHbE34Ma83UuOZITxptZeEjSJE=
`protect END_PROTECTED
