`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DaGs0oP8o81L1mdXrw+QWUL2ZR6YMYpxYfxYBFELz8tNCd82EAPSehogsnpgKd3k
+ctNhn5/WRdqpKs5QsRk0PgfBWNB72Y3msMJwlZ7/jAWYauy2HFXgronrhrww/UW
SNj/JnBNy0h2SsXJTPqy2QES4QfxBcl+8wmLtWT3+SA2P76bh0gK/0FEVRVo100+
//wWrV4tHPLwNvXetJYMFwxajn3W9O1iZgeYvTeYJ45Zxdvlo/OggnPr4IHA38ba
7Pw6fQNXEW7D9Qa/jbsQtqbmhcSs/s4DoslzfGFjCNJfGg7hrVveJkNYtYBlhNHS
xC76qBSuahTeByfeX1PQh6cZSrAGEVNmgXyBHPnVGd4okZ8xsjq21NkCIpy8t/Dw
V01OU4hptPE3kTNKp8PrPEZFluFGutuCLcP95unHt+wlZr817XSi+g29jTbLLf12
S40gVORLyn6ESBbeMOeLCRBh/qMCNEk8fGMAxQM+tf28ScIi7o6Ar8XGOwZ12Qqy
fYZBFkzNM/C1YLvU6F9VPphqKGCtNh+h3g81PCNPndq3xsFXwAXgoeHEkeMjGn3E
+tRXrvljWjgsjcYc29wFfjSxtu8OelRUG/gNbDwC4SQSozzflXRHpQmF90KplIzO
l8RS78fNtNuK/BnVavyyDssH4vCOHN9UZFZHvI/EihwvgRWv1stolBolX3PEAepF
zh5sJZVWkr+K6BR4TVqVp32F36b41nRoOLLxNuZQWsUXvzS/2YnhJWqgy2DIeYdX
vB7e2Do4zF59WlhRCdljuy0riX2H232cJZoulIiMo6hZkLbtNjYzf191biPn7syi
Q55/2gqOpuNJ+exjOveDzqMQTtEEr7eC15ZeQf3Q7t3na3h+Rtn7gJOw7mF7z7Ur
Oe0sPGY9VsFR2oEmRicUC4ongmfGJc9WO2kUowN2sRBmiaaDkJGJLjSHFxi29Yvq
U5wEdWyO0E2RjA/btYPBgG0bnanoiVGgNy8gSJCC9FWUKyrSDLIA74tYQ7peni3r
lFA3vFQOmZgt2uk1ksaYd//qii60A9EgWx33NsKh1sWTE6RH7KmLSeVSDHKEGKTm
BBPyx9/rgJHdmyD8BbCJtBKRtK3cCBZhrv7YXm4uz0Lhzjl6kJgrHV+JVRPrA4Sh
LeYjPTmBMB6eXDEBYvKXBoGs0nVXFppVAPNZKEQ1ACEqsh7PWgRPlEuDAMT0WWbw
X4+V/plEmK74e6kY5yGiCaFjByuTWNhy9Gvpx0tdthTNK8iBOjRKve9HBecqQury
bTwajnyqti8xA6cpDOWQO4NCtF6vLMFFkG/ekwISVfzZORM+fFZNi1xy9RzTYiDl
cUN13xTaUmWFm12YuBI2gvzVnGn26l6xXV4DsHJo7kQUU2BBw46LHiwnla1+XVIq
yYSFJpNInP8shWLB0qJxdD+fCkkPboiUWwOArJ3+v6FtWeIS1n2mbVobsmXjiCzs
hY90umVXuKzF/szYj7+grPBYlitj0pBPgAEArSMinIAwFFC5nyYnf07e0arest6r
aDOpVVAQsc9X/AwMlRBzWGGfoKevjYHwxyuEcA0w2QeaqLRbir6hCBgzV//vWsao
6z2P9OXjYaP+9P5mF2BAe2g9OcF5jTddrDfsfb3mR8rmnhhl2688hj6wQX9IfcRG
57h50aeTv9rSIrsxDIRRM5FprRnDby9pRoODHDEGn8g7+s9Hn+4lv69mYShKHD3P
PGyndARZVbc1xhow1r9IdJXzCpCcvg8X4Z1sU0Qpq8xAiSYoOaaG++yKHQo9OGfw
KLQxZk0ZHkXs5vOzXfqjc7T8MmYYx2jpzThPDmIuQWmQHxuAACb3XNx9yXiFNoqI
WsFhvq7SvwYHK4wiV2eGggqB73QH4h+EA9Eqa9qlJQ1KmIM5CLiCMBsDBZc+Y7y6
+PGr/fOdkRm+hpFpSGZ524MuptV642xiCApXyKezl6UkmqzYBVw+woRhLhnHkdaD
U6geWyPtLNV36MNIQ6Q0+aaSzAx81tnk5gw2qoMqC0h318+4W5ZVUc0gNxpKzX+7
4h/4S8t+yHHaERyghhTzeNtXjQUuLU8R/wJSb2HCyVTmQEq+vvg5XcJecTuqEZRq
24/GR3FXAeeIfOzuugvRuBN80UopR2Ny3dZSEsvfZlRVTJ5czU5sS5Khp0Ic0yMU
kBBuqcCXj/1aZV3wH5d2j39Rbhsk9WXZ2wfiraLXdLDaa6eqGmL6L8wC/NdqpmMX
Rpy9Wnx8i+xDg2fV1Vj8ib7NNy+8a4mS6Gh+nedZhLa6x5KqBPIlmRmKj6kHf3fu
uNY9tKBhZddpvNHmmjZRvPKn7VOYmVw30nfJDOn1R1pZMTOPS1NsCSXL8ljZkaVB
tbqC/bHUHDg1BCCaZgnA4pM8IO4c1090Dlonnza0W/cIBJyAogBhaJdxRZ+Ex8Lk
1VDz6w0SAeCbaLCE/gU2nft7+IW53sO4bPFgamjaab7a6HAUOuZeFX8/LktBf8si
vDHpsV3sm0eUNG3UXaqPl/+qgdh9uvgHJAhr7F6XVztOmkMrU0vG/ahrdd9Dd68A
LQoxKG5D9W5qRlYZ7KAnnTqNHQbErv/DWz2sEwg0tyx6Uc7fT2c/U6V05iPj9kKQ
gHkYvwNqPZi4h4yn+X1nPNnq2OCrbw5DwOUFpj1SkAUr6p+gX4DArNbqFozK5l2m
6eDUZQbVR3kDBaREH+IKK/t22id4De5X63AK014akrFuYFp3lqCid3reRlyGmMhl
N64epW1szz0qhGUqsnUcPn89hDwqudRPMsQBcAWly02dwm3lA3GIBg5Ll7tQ8P2t
lzBkGhYSV48aq53vcAjOGV1XWXeggx8wm1GmfhhUaI9rdh45C3gOXoZRo1ZTXuIy
vyxlNR09ZYlYy7yZcbQJ4hjN5shH35SUlBZ2Cy92KPaRAt3uTb+JaFQ2QKZZ9OM0
VD/KAerrY9M9GhVA6eMxs37Kj9WkZs3qOjfoTyqpF5Wch8R0AilDXn+KQodrMR5O
CSGc1tHfP/yYp+t8Ze68sp9CtbqIcQ4xCjz8+20mn2RR//smxzM45Zx2gHEdSyBp
hth/neozK5B6W3GhzyuG34pXUpvnxsIjDtehHmowP5oZpYTKoO7SWdbt4HWpToy7
uvN8aGP4sGWVdT6xZLMUUjjKWHB04id9U5dRYdFMAqzPAcKRpNi21M7VbmcI8yEw
QScOozCJ1LuL2BHkqn+l3Q9Y/kh/RtV4QJ4za6NAlAdVqtWVj2GB4ilU6bTDuQaT
ewURcK5l+sOhmqjnx/Lu7jVp0GP/W13HtH8oDkoPGFljcXyPzrLreGMEO8oXFA7V
imStey203/5rnDXWCiHtREZv0wmKuBaJtlpos8suc25U5CDZlKDI6TUIs1M80CTy
a4eYT6CeTXejT/j/qttKNQ==
`protect END_PROTECTED
