`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3LULefbN4FBX3TaPxvE9AcohVXxfjZe/ji0OBFXyt9UM+gx9Yfu9zMR0pbPnK1iR
uuJHDiZwOJepDY1cIiRfHvKY4SKegDQiTX3xNlusG5BjLc3AP4UwD7lqvBt8iGQO
zoMUIAHAUpHK9nOY9gjPVxplKggfLCAhiJy7SgE4fd0tiuxvcQeSOmVkAir/J3FK
R5ja9jTrUsFNibBWfxBD1WzFosdsT9n+xSAPUkzKxADMf4Gakjfl7NI/6rI7qrAv
IJzUyafYfNboI+l1E9lssdYZ3LTRwThonDuRuU1ZWikskIzye0ff21grLmGhWnd4
ErjE3h7AkOGZnwFzX4TheFzOLfwqTRTONUywpkLP70nDJ6RAGQHXXKCTQm1qqxyj
0Npt6UHRd12i8lw2cV7VJM7aIyHRWu2yCcJQjb6OkNty9WrMzShH5YB3lAiyYUXE
HQb/mzgXE7qM+m0CZgQOlA==
`protect END_PROTECTED
