`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9H8EDktPUfcpA5SI2nq/9YTjspIIHQCW1xG5lNT4VphBFAc0k+6u10OAgicPchy7
SDvu3oBc6OfIXDkqg3/bEsB/a/+uq2/H83nHFC0YS69uPRoN4aWD5eLIp8epD46K
/Yn7pOJCxYbz5qHA0H4xpTyUwpOYkFFP8YZ+ry2AGREizA94HJ4Yk18Tbpoy/tM1
0XTZtRk4jkF5cuZCUCJbc5K3sKHQn/Q/O2BOZD3ISCNn8Rdgcrr4t12m5mmftgua
eLdBOEYAXDQDtmVDUQODX0pDD9K/6bhHnTcfhtT9QpnAExV4qApaK4se7zwO0/xd
4oMm7+g6MG9jKVFSOeYJS5/C9HcBnbLXJ5LPkjrSo+9bb0Tu7v2ozTeLdty+bDvY
c8JDknSpMzQU0tIb1KMaOw6ad+vCtgh+y+bhkqM7ZuQha4W9+NL5XHTi6cQw4Ynf
/1nw7hx/U+NVgRBXMP5NU0ff4dO8cEtvNEQeglc0hwlWwVAOGuJlOdyRpqSCl/mQ
TE40RN50MWq4wmoAs2c25p7gEOwNwP/p3gTKNvfUz130WCuswpKTkubUZnibHKbv
Jtptrbq2lIoqRS1fF6eFFWUqwj8AS+eUAdSnHFfHJgBYttXdUk2+gBOFJDBW3sOL
Lln852bz/ykY4umXf9udLS2+oMFmHhERfr4ghD9j1EoVpCMX8haP1nS/it72Tx/B
lKJZ4Zi/AN7GD6SYVxUbtMnEGAzIltRXG0fp2/HEJrlYnLC4mFLEQlDrAECqEhoh
`protect END_PROTECTED
