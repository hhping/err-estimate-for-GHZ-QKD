`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Yv+QHznfhXL+8y4I8Xnr9Ma9hO3NmCMzfkNzBP0vidTFtnMFS6W/Tz04DWeke7O
gTLZCp8njLBYntmBcHBPv9J8FHx2OeIw6/E+gavx/zJdI0lYQ2550sMQtvX6pPnc
7rH29ZYQ8R09dylebI1G9nX7nxa8FGlG0T9WfaVIMEnIOJsJt5yCT1VESA0bvdkR
4FlnebdUq6GYOiTQl/j01Hu8fWfRcaB1Zw916zJQsOrTF3q7DEkRb990WO5ByW4b
xZopBiAHJsuusT+C+chziSHjpf07nyun0aczfCwXLf2Fr0SP2dn+XHsYoovuuAF3
GuHlhi1akFv2G2T2fmeC7Waz5OXr81PukI1aVSpyxh+WVwc85j4OOGT2YVAUSgkF
HbvUe78MCAuQpauJ7CM6ZdPTzd8ELih3Djyc86dVIrT7oKI1f2FVwlQYQj20Xoul
sctUSV5GE0zHabi2jqtpP0GO+JN9lhIiww10j3knA//m8a694i+ZutXutUpTCxFe
x4qzYOTmp4b5b2ObDhP5TfA7sCDgBK4uA5WBVUyWCp/x3SZbPOYyZYyjAVVCLMCr
DAFoB5RcCAilHkNi/1dVCBetFNm85HuGFpu3xKeBkAd4YeYANSSSlmars6UO0Eou
hME8IQvLB0x8Z7aCtZDFm6WgxWkl9lcZlE7dTOtrYhGriRB80u6vz58fgzB4YZkF
B+OO2pwjRP1IimJYjROQm6z2BIhBcvP1wDgo+hu3X5Xu9vKLgidWuJusedtjKDNj
dyC36fxyN5ViOnHDIckjg1FudW/6sWo4HfarNIf0cBhjEid9Lfcz2/gVsULnvW8r
UGpSYT0VAApFHhW748gyScRelGacof5RqYLRkNhRypr9QqCwYG24PuUWhhQDsvLd
iM9r3OTgUf1b8ulm/1nfI8qbMEMyg2qX5k1O+ypL6DqQ10t9ddq76L187UZ3Iuoc
ZMp9k/YJdBFs5yerXyidY2/soBnVPN/X+CY2AV4E1ppNO6UFBghkD9Mjcew6qOfQ
uF+IOmf2iiXHpIwrJmdb4lUAQo8LcS0cYOPmFMQy3yqf5DMDj3jkJ2GcSoKbVXY3
nHBJXeGnql3d9VVJlAvvT/SoP4V3ur328AERTDjrfUFLUrnjSOM6fp0PcSSZg3ah
knHni48frGZ/YCzoHavL456Q8dGr6Jphbsq0YEtDyyPfxkDOn64qtlgT9put+7LR
V+6VECJtKft8RP+/YLOmbo39h1EwZr1WauCq1HhOcdoOIdUDK77q8nZiHIxkkum5
`protect END_PROTECTED
