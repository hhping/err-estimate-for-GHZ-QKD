`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CLQ4dIHIrm39hKfoKwswhDlMx2EaaCwSMAlsX+EYBNQXHuksp1XuQwcJ3KwoxaHw
b+1NTw8QRsjfXVuzBBuKwhoPU+9xIhbKHNcRt5yGQzzzme9HoHLlB0J6Np+2O+eX
CZ7S8iQ9R/RwGjAi5/7HwijSqajBh03fZ96230EsBvv594lmgHgqKslt8GynTekR
1Q6ZYoGa3EQOV0U8l9f9QN6FuQkVvTh1iKbSShPQAaCc4fKlkX9+dweeCvTdFt+T
6pywsgmSTWvM0GzrW+MwPAwslypZ7CtLKrE2LdqauZKeyidAB39fzM480j1n1IgL
bEe94fv8uVDNnCbdf/AcLmFqDdI4zLt20bYUPTYFjnsoVLnOOuUw+aJqODdirhQD
pG+TCydbLh+qky7aMZX1Bw==
`protect END_PROTECTED
