`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hTTNr8ebFFi7w7k4gL9FTI4t5VNzgrEfZkCdb0YsTPGhZORz0CVf6qTr2GYPSWZa
IcDnB+Ged9RpyJO+oZ0xPLd70hBvV9JD4FMc74X0q+1Ak1pcSmiHPC/iZWqwpIjH
FRp7sn/MFcc2aPqXteiTVgSJX0CREFLTcKpPWl5DoVFVnnTjhnyFxFATW/Teocas
7qoc7dfQMhNKZM0wmI1QGNY3op4ua0mAGzMqihMlRTYhkfqFdfneD131QpGTm+4o
1bmrLcAnjvCNP3459rPinUCeLKlg+iC9GFCOeHI1tCoZ8W0BItLmTNxmM2L3lM4v
Z+FswVrg2UJsvuliKxVItjTDyPyNvX2ZoMJHm+87yGukC3P7kpLoaO2eI8OU6YOs
GGAvW/jJ12jxT2BL3urug17uGZwdgFt+1YtAO7oL9J/VZw+Y2xeCwm+edVggDA/2
u6hT4eCEbMpo3OQvrK6Boqw35vEgzd7EvP4WCTKbnEPGSyp8WnrCQMDULNBFJ0sJ
YXk4pqm5cpKwB5R2QVGhs71QsTjqDKAbKfnxhVhnMUUNeeRt3u0T4nIIuLVm0WTu
lL/cu31MYbOChLS0P2oxOgNzDMMzMBSSQn5/xb0ZNApKGKZzsZKI4dXqyGRquRx5
Bv/W9u1B6qOw1JO6zYANDh+eFXfaMrl4ab7eU0pdP7zCGL7M8hiiyY++mY1xA71T
`protect END_PROTECTED
