`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SJUU87CbuJmVYdeIeFojzXOJJUbldUw6uIXzhkH4IQbFn3GGEccGCxGKmavZxoLY
GoBaDiCUsvf5k1UTQQE/QzDxJcdZlpDJ1dyL30bkfC4BmubADTFpui2PhPwQjXCO
4gI6sGsK4ReJBsIlNIDlrhdKmJTUDWJHWM9tjDcYH0KMrOCuQNp+EpwRzz2nlfjp
K6AIV/ZxCWPspnlOqusXPe3YyXVwtTc8pnNMpqt3xpdds1aXHQjmE381FgQ523tr
5kbXSBIWXlOmbGeXNkS2sCUfTdPLkhz1m9J1pNqn+lru3HZbhz/0LY9WlpvlP1cQ
Fu5eG9IFv+Xsgaq/Tq81duT8h9T4sQGJAZ5bDDWHKF/WC9Mly1rMKwOb0CCKZm/d
H0NS6i/13/WONZP8Ro7P4vmHPl5budWuRlsOVBI/smMDSZJtxP74W0NYyReOgypK
4LZjY7CBERaEZjwaThskOzCPQT3yLPh4BBOa75+lD9PrKyN2emkuR/zL/izZVNFZ
75p8H4cksTwv95TO6yyAG1A5iar16e5+N2XvNVGSHWuiB0YgZwQ7dy4Y+eI2xsMs
hrccSTB7RRlAKKHjIuCOLrY/vYomCH+0wm0ypMN2dLz9nZPp7ewJ8FyShyPi5XCM
k79K+iu8lccuQayXX23EwnIVt5bgn3Z3FR7DvFkUIp8FNPxusN66V1bfNXRzx93c
+s+r4wnftcTDiEiJHSz6Yo/akpx2UQEbX12DESdYSXbPr9dlmPax7DU7qoV8Y/Af
X479QyVLIkmEMvfcPn8bOkmxPIS7sDiyI4+NbvP3X4Wd6kbqTJvX8GB/kfo0u9d9
9pwjp+TFLKMpTfm/X6VAnnAzkaRHs8O5cZWQOfSc/yEP8pcs9VUrRSEUdrkFoUN2
ZqDZsuhmHQq7OnRL0cGFtgb0vBmA5tlWx/BqAYL4cFdMCe+SOC35TYUaZzSvZ6Fb
`protect END_PROTECTED
