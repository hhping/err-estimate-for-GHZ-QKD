`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tCXUORG9O6kYa7conFHmOpfQ8v7PCP1N5Uqj6pU0cNe5r9uEKDRrXoubJfyi7uzS
yURh65F6+p/MkWO6hYrXiP2vTIYTE40e5bZhu4ZCGX9mFVHH3ZH1SadaN148142L
lV3ImXXYLUs+AXlfQU4kYG+QnLlfRgRnxeQYVKGtlRxe/miDmaIuLDyWadXNRrYY
Z0108C86gKbf2eOEjNMWz+wxstRo1n0wtpqB6lp+FDloa1RmTxNdB58IRDcX3pA6
GxcxedvQbsYTUQVU+7/ZPjNrKRly5kfSo78lbgwT7ctW9aPs0jAETn2efoAvtxKY
QDDlUh494J+K8CEbbh/emhoT6l5857Ju0XsYkVQpN72q+gGQVAohTs3WJOiypD+n
ZWVMqmYpJy8UVthoIotERFasHmb36K60eYc/Ye6BRtIsXIvNHminSmohxQpXIdSB
XiJ+tETMEL2v30R2+hj7rCBHG5LlZLeTGCZvXDbTqxv1Hk2Gj1y2Kivs4CedPeic
utTmAKdSvAkhws/ex5FCfFHlJ8uEDkBHtvVky/BSbohppMJgcZNQdl4VMohhyWOd
lHKVy4XU0rgdI6dgvnGv73GOZcB8ilHxD7gwYVoc/teHgJvDvLjgUea7jqXcne2Q
NaxcvA2/1tpINzhMEyCESFJ76MBsUoQjVqt4JkuGCrgBfKyxks6w+IiuO102vdJ7
hAOQwdyt7dgUBl6xbtlKDkwVjdKwJ5CKIwsMzaXkJ6EIN2bqTUya51sPdDw2WTYZ
Pn2Q0o9qJbt6/sAftadsiko5d7/MbTZ9zjN2q0GRBDMQngA5LrFcCtboqJF7l+ag
agqJz9d6supvgvnoStVa5kDPh8GzcEZ/BZG0/78Md95CE0Tz6ASeqE/oX83oFCcA
18e2Eb65BuLutfltTRgJeLJrqM/6YoHi690zJaZ9VzseYq1azHNsDi6kKUBIk2Bi
jmo9SS8iNPW2+7lGczeXbv4IcK+gVTfLCwf/l7Ooyzlr7H5+8TdXybiAWVu9YmHZ
KeWa9SG49BnOzhzmIqrfgydR7+JgrlDeGqwrkVKFALGxkI6n0KSYb2TKZmfCq+xc
eEl2t7SwpIlHPOrrCEkDfLkzc83ia0oZgfTfwdGhziVEsuPl3KNc5amal5ioPigB
DeAdsLi6IuCvWkxm6F8JWzn3fyK93lbZmLUW+TA14CYMK/k3YQ1U56d54M2ETU4n
da5x+0IWPAUnJ3d3WvYG+UJkOboh6EGzw5vVWPVmmW43v+b0LhXWbj/IPsCuWeRZ
xIZQnPbJ78MdPmhGAPLjuBpl6ZCW5yaLsuNKAwEpJBAnVa8uvOaufTWX3Egl17sw
u2UEM+FTmQ01oJBtIPJzbAx0BXXUFQJw1ITjOXcY52l8vk8B0VlZbCzMMu1kbnLt
AjJr+jjO4lTy+004YjaX7dVLOv0LS1B7OmiGknzYcADRQ7BJ2WbryiH2+YfLEaDT
CYqiGWGcA9gvm33uxvlgqMvqVBdt5ND7hrEhec9gt/pHo4D6KPt9AlIyJ1ZdaJ/p
zWcnOaSEHHVOj56mOZNy3E6moFTiZyYk0pqVNovaAnysux+d+/g8g5yuxDa5ngkH
GRsM9nLkZIG2qkA5nqzdkwV2pfl4CYdFAvdibI0p84bMbGFfzcGumCdCTDDmCKXX
F13mKEvYLtsvmoVAykQjrYc/pvuEySOebsONs6WcFelcQaMvMUcT/FphqnOJuV8t
jceioBzO8yhfNPqdBs9fu9pEBZNju3fVvmpflP75CLoLCIi+u0hUfaCyu/RAgdyh
AkxRSlKCkYfS1YUoDtJQWyaXXADy5obfl8NknKPs6jWZ+R9s9JdSCSmOmYlckaYn
eot+EVGIMeBOk/wbAgsnhTszwGexM5PKBIwupBDf7GQugQy5FoD8/j7CM8qJspuu
D+mLI/Y6TfISi5WWNrQMrjEJPVOshJA6fALaw1tEmi18IE4+LBg9orOX2QsLioFd
M95XadEu5HnOarqCyAungys/XVHQLoIaJTdiPuGK518YVGmfNrhYWbyTjhTvieU0
4HVSYiQoOYZxSFhxGrad5OIvlNsEHpW8hvRIT/Nu5cuFNgciMblqbOgxEfv3gUIi
Vc38Pb0uxH8iD8nyNwI4kZZ7Z1vq9sbpAwSvr2nabrzosiQDzQB+ZhX/eMbUg4qD
+2z9jPUTjUuo3mUnXGwesAweR04iW8Ua1Bxh6pkhk3qa+Ez5+V6JVqf+A1BGaKih
Nj21KNkDoUZ1mkgfGWKBMRNLsyFfbOx2U9YuqWHaFd8/lZsQYXKmjOyygoTLHx35
vcR/rsS3UgF6nR5wbUPYLi+91sSRQs1EynqxK4vOtHm/jCpePd0lKR4LXDl+ohIt
UFwpdp+JE/lRfmTeKtMolV/4cPoXKcj3uyAXGI54V61EH9+5q8ZMfAS0I8zsS+Fm
2vWDNS+EiH/pezeuagsnt6hYcpyZRoQRQY8/2XorwHU7sUw0Cgze/BFUkjUKyvmm
Bl3Bi6JW86kgKfBOYkvT5q9fSxTMzb6S2Rx91vdVa5M3rKq3/LCgvXyzWKerufCR
qdBRyA97aQmdR1n8qZsOAMtLwZ3hpESyP+hQu1V2wpMgWLFIZqNBKKGsQgazitaN
Rb1CLILmxEdwoPPvJ7d8yURdWtBYt82xDTTzAV4X92Kr+0RlQJ9b9U1YxNXkALxC
cmRHeoHOe4wQ811WXLJp0b5AxcBeW2WVX7y4rNHz9jmc5roGMhSEGdOsP07FrAuY
x5SfnOJ/5AxQq9IhSFoOnSum51DrcMVPyGxkEXDZqmHftpmxQS6MOLgVaieUg2r1
HPHH8ZHSQVkURwL4lfVwnMBh7lPzPG/glPMr+CI8/iA1+7C+UR0Iq4UoEIdX6FSX
SHZnRa8a3/TB9yQM1AFwK35MKDvX9nkLjnSUik4/nHzyFj4vyI4VrKdEbokeZOuq
878kbCTG4wP++Elc0/ShBCvMWTDLagOAjhUv79CSP7d90mkP+9b5R2T4x5lSE3FN
WB1sX+7dazMfwXPmLAlrdlBLUx1inRqPoX9mIg34GzpFee0g2EesW6abPChXVdeK
9Ic/tDcNt/tBcRRCDVSS/fYombseeb91HmGQ7xBu/0j8KW03PYKW3+dfY1Qchc1A
YL3tqNzM5TD2c3vY92lkcZ2CMvygW6czbRvLhthI6aY=
`protect END_PROTECTED
