`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aaeC/OwC5v5qiqeHL9S4P3CG8RrHp06UOY+lI8L3avWcIeQkvnJt0+5HCpAi4vX6
rwVL5JS+qXHflADaqZ5If5NVqhm/bBDTUyEUbA2tGVWoD541RG7FH6OtptHZ40ri
AvsyMrq8kSVzazN2EoAZt8uqiikFtidTFKiCiseYbOWxTkcAlCysF0LIbsRO/PL1
aqyrPaZtgVPQ0frVv568ATWeMCejoNUGNYv9ieYSH+EYEnOhbvFj7Y1HBoGY6Iqo
ijJsrVwjDhiIsUkje1xGNGaVDL0lVzEu9tDY4LF+FusUY3UyE6MYv0EyQCqqhHzW
YBg+FowdavzgBVnAboT5BCDLKgw1JtHpIsW1Jws27o37h4oo1B6UXxdcNaOkXE7m
jwseUXHuNfTQPyr1uwl98OIwWJOun/zo6oRu3s902VRHAP37i/RPTHQ+6pvwYLdI
TiaTLulTQf/gvnp2tVaaKKVGJVh5S+IeQDvke9BK7TDaRTa8HFtDq6GOUxF7GwYF
bjvMu9Hzn5asGFjfLpFKDe9KlTu1MGl5edBXVX7tZ6hzTPKhMf4lEYfiTpcXnziD
`protect END_PROTECTED
