`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IcvpU4fAeowhm8YrWdL9tporqhDfvyQf71TWLD7EE1TlpZJ0D6xwXk1yUJbuYhkw
Y8pv/DDN4x9yj7r/+5q550y2OQ/30NVrNH0gF/6gzGuxWcJIP+79/lnvNzJR5sHS
POVU8WzMfrtgvdzz+wO6FkmbDpdOHVZEQ+bxLCHIpFB8EC6Cg+15YgVAhZHi1SJf
XT4aGbOip5bSq2dLMtr88TJjVPFpe+AaIGhgGueR53q/6q4qCEL6AonXqpRh7Z26
mE+rHD38GuBQu6ay9KKpNwGFzJy4F3WEueHBPp2jNn0Ku4ZJn43Gy0dEJK07HMLu
wrOQz3M9XqZ7+P71QmKKWySq2vRilDnIheC+B7zh3wATi9joXcMmtU4pcEStLurB
+BChwg/62W9F+2BsQuMVl8us4qj8y7v7MDb/DdGgxno9ZVHliCjDDNb7q+SSQoB1
nwCLyitPec395j2iA+lx/cw7GZH7tDpkwDK/7bVaQR43fDGCF/U+58L6Io0jEYJM
JQ0QAQu8+0rPXc55nLAQZxkI1KWs6gi/1+WZVL7C3UXip9JFszj1TMzk9ZL2nAZ8
4VHKm5w/mMhpv1kMoXkObQD5jXDplSFCwSMHKTSGb6RCk/YRGBK/LlCnOblP/jdU
0jdWIj2DXSmwM9efFNyW/YRDnH/ZGKdttbpAkS7YxnBS49kPdRMuUT3ZzeshqQrl
KhD8Kd8p1LkR3dHTasVB/Bz/bcUdZ56N0h6gAD13bxe+7cb6mrw1QTpCOLviEuIk
AsICwWD3qqRln++NrYRQLddOpYVN2ThdHWj7t7CsiuamI88DHDPf7zWHmRsQJn+j
GXA073lrYUI3t0KyW8gsRKjGXLSg7dNsdImgasbMPxPxw/zyYyclo3xBfzbPqND7
OswU0tdl49rjd23qoSJ8fZdZkXGgKq/M6rHzwPCwwrx0Im2TspUEFLTeTm7lc4FK
3jYfcvnGQ5bZTYt6+RWQboIlVgR9EDnrSiQj9L3w7a2muKfu8dyxEYkd452uBA2c
evxZRHKJfBwx9p9vykNKpLKzLENQRnq/KeFrlJHQ9D6L9kiLOFC8Z5MQJx9BTUsk
eCZ54uIz2gMfoLfWFuF419f/Y0JWLq0KrZ7y7ugpd9C7WulUsZWWaqNDxxvDNDv+
TnZDI4Fgyeatke7jnyw07PZlFbQoLFJ/eUwQoquoUHC0fJ8awz8kE7kbmcIO6+xy
TL2spwhadv6BYxeEI24GjWMmGXYHkbwGQa5hMOEPHME7w/aqKvTVOsvXb7dKALUT
uUIStK/ddRBphitJZVo5pAIoZVLcOlpeZR0ThzSHpjU24lxeHuosciRHKJCUcpu8
Hpd4b/2WWdTGOpaxam7ztnt7IzWaHr+iBEqtdAmvD5VWGWlcF5lCNmaSgKh6+PTP
Z5maLS3umwlmcLfwoS/P3mI/SauO0RIQoEMRyqAKB0fZ7D+t39ieSnXk30N2m/Mt
PGsFwnuLhnMsnqrlE8ISXtgTX3MB/PKZ+f0LOZ+6Q4zw37qkgqGW5PYyi+0M8EX/
OXuV9J9bO5qWt0qXGf0oG+sP6w3TBfcTSkmOphhuqCqjBZIg6SrganyZiZOPS4Uc
nMGFA5EIpZHfbmBhk5hO8cO+EjQhRMBxU8dh/rYlZrF7xPxIYxYW+1CO1cpX6Knn
PhwNmtfngIP3Ba5poSh89HOuSRM6n51mhdfSCIWZ123AhezkW3aGJ4pNnYG8zkax
oiREjTLII9tmT6NUoxeWwPBXLV6d9jvbRC/LXIBV2B3EjAmVHlUM7l91geRz6cav
u1bMAtA9vsob5AmoGHV1K0ZLy6ry8/McGJTa5mebO4jv4z6NIWlKyvrPPFu+KPGh
UMBCAqhm7zvJVDpTEDTgmtzmSw9I/LMnJh+1JRf/fywDx8XvwpI2kHs0SW1s6K2P
etKCUAiegIwjdcPsVZH/6q7VD+/rkmjCVl8VIrqRVdVtcI7tZD+/t2dPkLbUiDyC
1BfMb1GD6hThEml+stf3POB87rjUF6rx7kYdit0VE2O03MpubMKWKxT8X4AWNwFR
uKCyNS96wt3IrfywyIlpB0Vfvnyn/be7Ck/slvwBUJU2a4MSiJ21BZ3GU9cUSWse
777qayl5Bamf8wE5fRF7Ary9NuN02fLoOVJGZ/fwRzImgTSBW9jtX+ElLtR6Sc+v
KPaKQ38qikpt7euMTOoXhInlThedSQdPI9SV4zkkBO3UyrMq18vuFPUmBMWVIgHA
Zkt1lpwqzAE+Ea18Bn2KovnoyWUdP3/T+jlCNS5JJHkJjYzSVPDK2ssKfOZ+tbzt
hPS5oII8V3XHogqsBPHnRymyAj9jeeABtnAe45+YTQfOmxt/Osh+QhzySsGlc/KW
osGZG259FwBwZAOBE5bKsYnvYm844Bz7TQ86118Avs7DWuJJUQocZupUAYxcUsbk
WTOLtE9mKLYMBhh0LA9DME3GHG1iu1BmUbt7tGi0glUrC6YBz/O5CRJUlPXBEo0g
RIvtxSUSJYyYruYhJX+vmZIPT+whQnbxueGOniSqRl/DOPpzmvOGwb8FLJimgcgA
/7MUH8i2ic053kINuvjAeZw+lkGaluuD14VOJazf6kkA1Bqdj9/5kJ3161OsYO/q
JQPWsDLJObxydJKSiDY/lYuovWO87GnqfBMpmxIpAJ7ff32z0DDtAdi2eUYtBIGR
B6lL9sCzhdLK6uqdyhZBkde75FM+MtVsmLj3NGvkD4vg1gkStG8ePm/B5XIFOgpG
0twNrZg+ANsnj/xhOnTdcI04Rb2YIuVj1Vh7Ah/9U2hiqXUw3naW946qtQ9v9PRG
`protect END_PROTECTED
