`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/xlr20Z2c5GIIghhEL/oGPSBXMzXH/lidPAfholphzYRw6ZucsZnaS/PgMVca1gj
xt0R+DNaMZVPOrR6KqAePlmpSv18+D6raS1X8oqvdNwDonctoXAW8FXyW5Leae9E
y8T2K2E4akQftiN4/ecduuaFjhsYlXaielu5Tsz74GS1nns/UTZYeLSt7MoA+SEh
+/8bSVBhrxXWso1j2UQ72ewLtZxaRekFvelymAM8uyQINb1CbPwgccw9JOVYaldh
m65I74h3pII/KrMOHDCB8E/dUYOZ+eVFTqPB25BcVqi3dG8cOsLXKeCwirO0Qh/7
IHIAut19BoDzBHYyeDrPHWh+mEouvyojfn5T7HeqtQUwfd51GFv+rmfSYepbUHGZ
N5vnKzDmKrMKD7A3peNOFL9Pu3u9xzODwtYXcBD1Aj5p31JLt7MqWtdqkxOhhcKc
ysmULQpCukQklJdxSCNRz500r39R/HGwLQVEkOUWEv3XnVCg57ma/vIyBtDNyKvU
eMKFuYoemnOGZuBfB+ofCLIv0BjI4u+GNuVnHXHdArsy3rQZF9FoMPAn8zxUp3H3
exP7+/XDFBbeDRdr9U9dnGBOL3V77DYXVGJ9THDlw7G3BQf1bMxaXis2J2QaF305
RTc2vjoZLEW0LBgGFbU5GGryP/FNp9yEHQAAvbkt8PztDvbYg3R+2a5OLIxmfm3k
I58lXtoNH8S9qZKmKA/VUtr1nAKMqJdLWKWv8/A+QbcYQOE/2XjEdj2WM0G3v2KJ
eom0O7I7p+7MTpnM63BqLxarWv2U0zmOGSbEr3Jl4kbxJIuBfCJ+wCRP7WcWU3aJ
QKmEemt5YEvAkVkJQKtPrutxoQ4vGWeucyyUqPJOUkHZ5fCyUp/QVKVrEMkQMC8u
6iVfSw3u0vJ4CcyNexbT8g==
`protect END_PROTECTED
