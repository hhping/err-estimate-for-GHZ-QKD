`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
49TTyCEIfbX6uaRZJGZZp5d/YpikLY5je3O5BfYXJ6bi3v921nZdPCYYzQoSYD37
RK3lB7BfGjXJRt+S0DZwJ1/7tZrWlriyHBnSvty2nfify3kdFpQgElYJQBLBEW3z
Q4mqQB1+T5fXKx1/u0W6Fn1D0ad3HD/Y6fz8fH5vTEGNFn8jQ+K4rPpvsDoiUFLc
/5vJPIQFuPWx1iY/i/5UxUoYWNfT+/A1DhKpgf6851LirkuRp1oqecpoDCDUg5z9
0y0xaT/rBVYhRrbya+ktl4QoRbPdP7qnaXgkMdJV/jJwQRmZ2mki3g0Grob1b2v2
2aUCOJSw2PG/jq2TMeLWTQQHjKijioP41Nqe66n/71X7OwpUDuRT+/NCvX0yXVjB
sz456kRVsdJqr8NIWxun9EQ00upxaWQRsxCy949zogq+VLXS9IqF4xlD8wGkHb1X
VlU8HYKeFwA2MsSSesGd03dVjf8fFfTqeBoJZYQegaxyaEcqnZQXnxf5Z8YrIGik
AZvcHpn5v7Ia82x/PKEWq6bAvwaC/N4jErEZdon7OSzD4emdxLGk3RqWtVNDTk/8
pEN7Z+3fGTvER31shkdcr6QSus6wsDpJjCHyX2vW10TO8V3alyfUimBn6DAgf9wi
fb/WxwzV4EgY2uESYxtygtcnnWSnc9K/dWLZpzA79yMK51bZsCpjkvlsUDbZHYq2
DliWjMad4e1KkyJYbNstt30FtuRf6wrO8HRjS8wpcq2UNHaBXqzxmjH8LjJ+s17s
y4yaEZh86kXMXPB0r/PqL0bpsVBHfT+VFowi4Vlx0rcBYQgoZqV2z07xwDiqKnqF
2KvR36CrFrCBVIS39w8NnKAeTCotaaKrLGwKyB6Q4mD2b75f6cr7T1qdz/hpIYsi
9+cSxoEYHwtbAqr4amCTPvOqrJ8F9FVqLhzyJN1QHqFpnazFjF0zqTEFEP7pyccM
DE1jZH6KTDWFAvJ2QSy7JVl2vPEV/LLK50wFvtaT8/zcSwBK+VAGorrjw/qCApYF
3FkOUgbGLlcoJUw4lkuQ/MjE0JdvfevhBUeEV0v9s/7aFvVk1za+Hl1dl0YwTc4g
n8pcwkPbUaoHV1W/uRqiUCQT12kS9yI9o2gV2dq/pgAGJG75gRPbEMhNrADNMJgY
LClBn9w3Sc/qssiSuLlLPgnPfqT5V8uMH1IZKBBYT2g1hRIe4kmzhOT0vKG6Hz2H
B/TGHac+xFGTHVSLIaK5aXSGkDgBvvziNI897BWPyaaURYQfUHKLrBOniTSEDDkb
Tb5y1biYyNnAz0HYZF0M1In1D1SxHKHUM7ENN8n6g2iY/8tatKwXUjlRtSew7J2m
o9AIu4Cn/Op9CEMWo3O7RSiEN9GfmFsm25Nl64xnAh0qsGRqOKiwYeunVVLTTyze
HRkIUGbf0N0P+nk5W36Rom3wEp/n3OsWEZuibV1zGwNYAM5R6ZDCdYTlZ8HDUHe4
0+0ysR7JfnMsBK/muF9xUIXr/r/9ROMtf37MvIPxxEVAb4FWcHhOh8CuQdgAJn1h
KlkykRJ5XVWMjsTKIV8/ofojbps7jSwhlmYbWF7U4i/tE+UEyxlACXPWHa09UhXx
dpNFgDpe2fQUAS/AFTHmXtbxDazAiAVUPqJciKo1VsVvVnLcTKDC4QVX0SHr2Yl2
bu8sVzro2IgqSaJ9IXIqxKaLKc+AEBb7CY3+9cKK4nK/Lp/cV3YXUfKd3yVQQmcH
MqXuOpfePFDh17gSF6LOb5DLRNrXBKSLhgsDz0ZGVL3ezcR393nx3pfz5Q0YMbUS
qPG5PMbHyf8t70RQQcXeFljByD2xNKeVbb3eVR+rVFz8Eo7Otwyj0zXkXeA2VrpU
0djM/6xOWo2Z6okwaUppe43rPlmMs4IsDuyXGMySqHBwYy5as3vNTYADhKXoLWY8
+ijQXURgWsd0FvnK+MrA1a0KSxyUN3a4YdARmC0BjO6AHph9KGX12B3KuLL9W5FR
u3nvwcfO+k/ZSueqS4ejCK8dRSSv2r+lxHYjUKLuos8KlqZef3FJhaPq3cvOQH/d
cugDL+iCBXcjx+q+1WbSslHmowb4QapVt7drKBLbKFMzBAeuPoTYvpoYzAnyzGCU
FBDl8c1Gv0boCaMa+Wi2gAdjJVZ/HgX2TpHpoEHm+wG0CFaW7J2bYrPtKFYuzA21
y4xF751V3qWV349MRQuORftMy68mZT9GbU8EJRJQ27G4SCNiSB86CQyZGzY/w1lx
oC+gOH4TIkpR6MPBorcgorBtmxblJELVqyBGqDu1Z5e6Uioh7nZPtLOYMF+AMRNP
jqoNNauy/O+qsMS2Cl1tvM2t6W2KiWRomnjh2eF7f2tROqQOhNi06xSg6DPGSHNd
0K1bWBi76vsElmOCrWksFmB/SCQ2ZO81mQpSe+Ee1vzLPl9mYX2gYeZ7Upj/tO48
GJAXlQBzK4gkIx97ENz2S6uqIbZfIDgOajcJIHyvtTxbYTEzi0RU2eX0hTMLs32j
wkOFlEDVU+1rnYRiQEZm92S8KTO6VyypT8MXtumpPCl7GKaP07IxB9rgLEE/vUmp
mr7mACJ7z3IY/YDVjZ3HCsQb2luhrGnHOx57852smvihPSvQwoQZS1eBQGR2Txe6
u+hJtudMZEDm5KsUO+/dFSOjUCqfQ414eW+D80wtKiqoYTdQBNvPE/7ai0xMDbSh
zbRx2t3keXLMjCCQBhgb+eJ4aSp7E7usIwSVB66bGYvn7UsE7DrVPWA7NVTbjmMX
P7hxEjbpZAYMOwKppoWhmpIPVOWnPct/LF2bDtI1yyET57RiWdnzG3tysAbZ/dZF
IdWNEXm/qmVUEwjeFAZTFloOysP0VdUn5/N5AzA0teqjCFDjJ/JBiA5+fDLzz7ri
8tOo8jjbctYl3SVeKkJb+2uj6ZcyDy1KGeQ7xR/+KTh3IT0ehWlQrBAWZI9h2qnj
vCr+iWIVCP+0PbBsGP6iAna3GlSnOPF4UQva0UzKRyJRdSStw4JASX4UqcYGOOEZ
5s7Iw1Ns/RsUAIDzLmp5SQoFhz1QBwEDF1lLEznmJuc/eK6evhW/6Wg5Pkpq4UqW
h5M/POx8567ySYJ5gP6ZRK3cI68jPTVNfArjRdf8DVJGf9XXrY+V/90CCmRVwSjM
eRusszkrbpeHBykJk7hcvq49nC7lbelpWOAdywzT612p2RnhOhk22giaHo6m8eJS
Qck9lx114KNWkFImU7tUfuD4KcFTY7OJK4olMUU+1jkMkpf9Vu59fLGKvrm9Scnz
TCwWNGI5jS1UKooSr0bIsN0VhrDJdeMqE1RHO6q6JURfaXUnSZVok9TAUISyRhnL
pddJSRLPyFtL/WQakR2HWVZAVLmnyboWhY6pU98REpnvP3mHolHWi2phkkL+3RFb
kOk+7LuCLjbdh/vw/9nANq5GP+Qnnw+Xg0BQAQZTtJAS7nEG3XL7j+t6+Uqc3q/y
+URAl5TW7SQSUsJSqyIsCT+pExN6kVJ76bEf8AhOqGZ+maqhU3V1jKxYfHtwj4Ot
6aCIzbSHPyaR6ewDvWiXkGW62CbwXXAZqPEhCLV5jMU5hE0lZ6yrS4ujEIXG7s8g
fVGTjq8NKMyIj2LqDz8EuLWprLqBj8gbeSwJIatOVootAP4dgLf8iRCTmQzLwQja
VV2107uj/Zi5rdlpAzl2/Vtt4ILK3tDslQ9OgKm0RfW27xDZaVWRVn7f5bLde6oP
JjrLC7WGRlOm/uDaPUYTJOdfSG9ObChIaawoNr0ufBkagqVbNpONBV1lq9S+DZPS
w/FhCMulaIKYj3xuDR7pHH1B/BUlTSFGu+oFiczuNYFlZzoecZH8BXa2p9DT/gP/
+GHcD5B0pmr9xHD9oho/rgZSqLC24nezwmQMaX38SRNMmyMZ/CsFJfeFu32UAAr2
JALzWCKiQPV3aYU03YOpa7PZ9U/AQmF1PWgWvN7X+sNxFSeOW6f8OoMzUXFQXi6m
4FR0jRtuyECm++k7U663YfRQbHrER8B8QrgOi7HmF5tfXzx6h2Lpu1fwI8lo5fuM
6hqZIsvPCWqTcQhTRQGktOjZXu9W1v5By2X182Bb50qlmtEJCMvDbK0OsaMa4y0b
/eTJk4i9ktmsZMnKw+t7wGA67P4yXo/5YFXR7/2qnAMAKm8lvVVUBptiIEqADqE9
xXYcH5Rhd4bWnlYJ5ucnBLpgeQ4xEjX20Dg+XjgMhJpswIHiASS0aWzuUj4azL1O
UPqXLjOHSQFH7YvYlFT1kMyz6gUNHukPeY9APR2JFH9D1dQiVIRNCj8ZKijGlhYb
OoXyVPaifAzMvV81XjpMKhnvArMdU1S5vD0TifOAoWHOyXXJzxRFurcXcWMWD8Zs
mBjEQVWg9uboMihQLPKn7f9cnAcS4dckmBCSrnh1SW5EpxB2MO61xg1nvzJyaJXQ
T5+ri7hISbMu/HD1/0HaLz9gCuq2xUMEorNhnaoGQRaT9iOtehaHeI7wZ4owWe85
tCgHMlCSssaevVmYSXosuVSBN9OiqG8zq3GHF/aoLLngqxcWGz4UBHoRgU1TVh/a
uoK6SjhTs5y1R2h+D00UTjCRBjfCgZHk9fM4txlXG5vqJFF/3/0LDEbnXa31fjY0
v8/SPqPqV0QqbWT9Mb8UELTNP/RLcAaTVRTiIfW1QOKZTiGg+tr/LbVN/NULdNYf
WyzxIjT17AdOVpTFqegVjpHueS7LhjiLkxTc4zYzTh8saa1zy+7AjEPX0QVm6Yxy
zJR1nf3qvCu3xyZ/9J/n64gteFFBnaLXfQZm0fjETUtxFSybVtlZplfhz9hG03X6
LSMDL+/z+Gf2HLDnxWjCZqPGnBsdXh1JYPvnnY6JTKL+eO/aZhUdre9skxfj5aQF
rEK8stHZURtYtr/AhJToBUv60xGBtQgvJLolOTVj1XnlZ7rOI3SHdvFYNz1j9l3q
PZo7ezZ583pz7NNDob+32At3POwqQPQ68I6TNmGz3aXSIrNH32vyFUR0UrC7pfps
da27+dZK27nqHDTg7Xq13sXUcnkVNdQez0jhgOi5omElhL11NjWpOG8XyXPCqfVS
9994OactRiy7071sOFp4u6f8MvJK32Z2K1yPHXfCTvLDKTm9YHXQsVHJxAcPmI7B
rCfmTeC63Ld4IIhLaPLrXHcMhPBb/bLBDFFrARxjVNzZ18DXZNgwhOSqmDucZZz/
SQlovtOSPcKzjGZ8BDUZn+4tvmfc8R+YDjmRxsRbBwcT01evZp/DjA0shUWiNJXc
tEoWC823qkqQhTmYEt27xgOBQguI69V1S8LqBMqJAb5l+MGBpOL9JYa2WDBG8qto
LY6wghBuD0DgLuss5xeMCTNLf53kUvy/lHNJsEhjTuXzbZtIQzXS0/RUzsNy6Cyo
xehIu2YxyUJwsRID3ou80IyQWoPbZ6MF/ZjKCMgQD5zOvkaG1Qd4U7JQ/2vaOW7o
W/kjM+GxEfiOKKdw8AHKW9lqTx/DNC84gXedglivKcKHitikdZHh35f0r0J2zOTY
Aykr1jOCgiZDvxgQ9t5skCY96oBxszrXdF9Y6RPV1lp4vT2patV74pvgLFLnaPZy
l5LJzIDbcdx+Rjtn7gtFMFmelNx+ev3bvzWS3CURFO2PY8e1R6L3Wa7Bc1k8kCYo
CwlfXnPUhr7O1nyI2jMVkRWORk1pWqQsOmtEBrey6dXOtWwm6AU0tHHc50RIYgBS
q1zmbgyvQFpUTEZcDcSoIuiZ5WJfNhKchtqFcAG7/Rv45BhqpGgz0aMiZpCrgqya
GdFgoR9126XaqsdDlvygYG+8pQeAtSRmyXdFLCCMrnhwELcQd08JoP1xggXyKlf3
ajj8MQxvGFl92uyrElnnOposVh5ISasPwdAdIBSEBbQvgOXYSCfejESb7sJp2e+g
5diOWzZavb2U3RlQrbLorItu3MbXlsasq1WPWC99gjTtPXnIJaLrYA+5IVJZHYuA
dSIMqZFX/MJddK43gP3vk2MijVQRw8uewz/fey8cZvgTJnOnWnlpVw5cD/lZJh8j
mXTqJ252OJ5ttvVjtrMWsGbTYnCwoX9U9LFmNeOzKKm6JUzF1dD8/2ggE/H5omaw
QDb3o8fawDnOWzV98X/4/n0iykW+zYyHflcEDWARwpnqEdWWpFn2pju3RbIHO8/l
h3sl+bKq/FGO0cbndETWkylPsQgkFutvelFqjg+ROD9P3jQlG3q1P4dg6gWso6ln
pGPNXLgge16VByp0ZPDpHjX4LYEFxg0pwEqh2AkbTafLNCwr+aiyoPujHexZeoKX
S6q3Jxm5NrkTjVmCeaktAh0JIKSKxrUZWm883gnMqb/pYIdLD2JWoX3yAkxETiVk
ZqJJov8uK+OCcA46+tdPn9ikYAdqCWCgTJSV2g++MhbP44V936iEBAtZsm1g402X
GGwTlgC9MfpJqVXgmpsMRujT+gMLrBsi1KkHKSoNUHqXmUhn4rCjbN+1VAEtNrFV
ffAIetnCIrHMejk7TRovBVKvpJNr6WMLBkIHEXx91Xymtmg+IEiZHoaleVwz0DFO
YU6gVInToTjdG893obBjbCYtedofyYRigSV6uJBG+79KC/AMr4b/qwgvV9PvjfIl
dyddkdHW5vZEv9n65vbX3RzQQcapEvfWk1nErDbx603XSSCWgvkNmsWhxj9mrOyN
jqR5Czga40Vl+MDSlkg2GdTwQV0P+z/OBMwJcijUqRL1N8Nd9woUvjsuOAhCFuOX
b74lpNas55+tsa4SU+Lprz1GY4xud/sm/2A0rohJN/I1Qb/E/SmA+iZaW/nYoS6i
H64H8sEsDwqcgxcqvHJCUVXlk1TlW+h99jxuyDcXT2X5XBKxARBEXnw+3le42Gar
kwDOokjfNGGmw5r9umPl2KFtcSMi326Pc6uW/zMDf62xgPSshkQlB+NMNLPKGyyM
z9/9X+wjDdjgVj1FgYJM7psOc70y1mkDpeAPQ3QNs7xt2SXFZNDBOV5NBUF0c8VQ
GEgfknvWKpA6PpObwZuJa50i5NyDGZVwANvhxV9ZD0BDEVebI2cfEe6vXDml09rx
DYRLfJeajIcwoIv8I4mAbj4bmxJEL1mHJHvTnaim4me4ZMfrv1EjgJbaRagfcIFP
sZVkL1jNJPrRbbuxueMQC5maXU1CMiDXuFUAJYYugs70qAgeJgsRxRoUu3zuAAvv
+9GklTG8BxVu0pJCGlwet0BOY7iunEaurEWinOsgIgCRnAbT1zxYau2YjlWZPHBU
+0wOLxX7h8vkljx8xtWuKf/SfY5HnA57gK59SfFP6tpuXlCc+w5RnHILPCe3FZyO
JO56vcnk/N8bWZfPQXqDI2qUjx76/DqaAG2zx1Wtqo8/Woz/mYOsfeGafK8u25WY
XTztrR2yDbjKVLjOIWwv9eaFjDXesw013jsN12Jy/lAoYbbFo2tJl4w5GLm/bvt7
Ut0AiPJELPnCNHkeA0sPBHFWRK1C73INJkSvshCiEkGz0+z82LVkloNE3TvHKFdY
wOl+qcqUlFEa0hrZECf6XdGyn8x/oZqQPYdbM135FQb06w92IJ5GEU+SfVjl5vIU
XdXNJLtStLf2Q+Unjpa4Ntg/mLfIHeBcG2ca73ZlGHVpmWEbg5i4STczkIZYnhd7
upS3bseYUYqJPKR/w2xRv0LnrrAepcIy1JAZg2v36apXgG5cq1UkAb0FngI1ZX+8
vz9hW/Uj8jgrtbTNm5oqpeMpPp7I1yE92sPVV79+Px9Aep/ZhlCnvkYAF1FKi6LN
oO8R4Idca0FmGhliwb15x2YzAtHn9VLKsJ1n9xRTkxOJx0eMn0XlrJ/y9UxXlvUT
55qBjB3NMEOLz3LPHev17tovkTuUwScd9c3gOBcPHMiWzruvnQbfJdZ9AcU2Qrqg
v4MjLA78tQaJn/svDWry9p3giIU22uTdpO6i7T4TagvGjkbAgiwryjM6OTiNQIoc
nxXnMNuRygVLYVE90vTi3VxDFr70Rf8PoBneko1IMSCanmWyLIt3ozTccnpdMFfy
Gj/yNcP2fQqqfGgwVOZKnucieqDwqd13Vbe6w5MAvCw4ej3woWPD1XcyBwU6Q7Ow
wQ2xqJUNrELvSbu2aJXSqqC4vgJ+BEmiA61J0vA5XlfhfMWgxCnJ4wNthPQ1LG/i
SoUANapPxRGElGCwb05BGRndxtk6mbHtH1wo7DS2MY9quXebzln8/WWn8FMrUbHz
nyd1ScWGWqWYqqWo5jq0bVEG7jErg3QOKNH3HcaQs9sDY7nzMiuKv97AkacK2BXA
sCpmLpgRlPVfZj5ROe9bIrFwqAFR59T+Ki6WauL/p1HR+EObeWAQoFiH0p/bLmR+
In6jNtiQIZhCQyIy0spEEVK8zAUHmbsCt9Uin2jK8a+O4zEuKTLmU0C7p+5Ik4q6
YF2b9xM1dP0rlTMpevsMVtIYChRIH1d6/dBMl9nXNSpYriosA3YUXWNmNy4GKj3a
cel8Kgr1wCusfT5WfAu+bd2UDyEBNdUpVZt6Gs7xg49R2INWRl1d+ZOw24FRGu8j
E/7Y1a9CHro1BiWgUT6kh+uDbOOceSYrb+L5QXQaG7uAMDlEFewzlCFR9pAziBYe
V44GFwyFO5lB8aQqgnvs75TUKTW8bJxSY0wGwz75WpDwTJOlRpaDTQeCxcc+RB3l
YtdVbec8ot9IQYC98/qy7Wytf93K/S1LCAjGYcoG0HUiZI5AtkTrDIctKYN8rM5v
KzZWR38RvxjUK+eIZTBkgOR+tqvfFKo29d33LvtKQD1WLSNSOA0VOYW2jYEG56cn
1GpxCJ4/TVwst+UlnpxeUtHwUUZKQHKiPOqppzET/pEs7//qHi1XbzxYUHOIGzzL
cAMDez/3zaWDME+1l9MZw6jpqcYTTUj9cB5ZsFvnjay0Az2EREZwt602+hj8VBX1
42Qhph8TQRe//0bfCuRbi1hNLggv0gQwoQiCbKjH5XOvSexBhCzrNbwIl9pGaGBv
C2cIeAjQdc67tLcrr99BHJN2sy8ktiUT4l5IY5aqYmmRlFPLSKY787jkS8H9dc7k
p4bcQdXGNHNoFqmAc8+VIvKEyk9u4+gnI3Vlxn26/30oFu6YqAyOKwbBhrzKXfCT
QriLceXUHKqbnHHlvvE67118GDiJVk28kmaM4m5aZpVQU360c6dXpY7Z4z0T5oPo
NlYaHzCGJFKbFSEZtwL37wOLLhcFJ+sYYl3tY7ZnICREMIKMK7Bm5W9X058TzF04
T3fpqyZ8wPkBJpa5P9CCsw+gmfkg3MNI1SpqAWMS/6K2JMZdAAF+nTcCsPR6CXG1
ljlNdTaMC+B6CInZdxeTp+zkMiEluKPu6HiTCVUlQlO9lNqKXmph4z/cWlllPR9X
aJus8UvFc0D6ecbALdLitHCEIHZfynGiVo2Ctj4SAm8lAvn0z4pkqiXCb/qkWibH
W+KIaB7vkgQMRp0zyWihgpH0sEHIoTYwRVLbgPv6UmosYl1uACZDT4mziGBQN1DQ
TmV3kdiBLZhzH2I1hX4HbROTw7W5AAmbO9Fz37dKnifeKIbGQHfIVF0VcNaBO/Gd
smDSRq1Fi/Gz7GWO+H5cBrj2wGn1XRHkaz9duhaCdRx4Vwh+Eg4ibkobcRxLuoaI
j8E6l/1WIW9Fui2eUknp6Q5wnrL1Oj1xR2ttYQmzTLvY9j8sTORLmvzbBYX4CRRQ
DX9fnSxCH0/YL3HZsH8rr5s6HI9+xRhwF17+C6cWUHMo677w+j+d7Iz6/ECAX6nB
sblCPFNvg01pBwZXZ0UOAyRfv8LeW43UgfwS5E/QlrOaUqb8i2UWm/79jPWJqBkW
tnBZ4cXURJVRt2BYq8d7puTcw8gqdhfuJJhl7BmkW7phMMqmTPAaxWGeRKMZjoDV
3zH+JWSXu22RIVtmbkPgF4097X3kTbxrwAG39LH6s6CdiZN4U7724aVfospJXets
ZI/XjfuXIxUj862A86jJKFzHfcZtN0ZyYGo++YZD3nX5MF8zZquaMdTxZEb6tk9x
I+PBIYGuwPAk8ueF12qW9k1TjelOxVUJSgLJiR+AfxzsRA7pnQ1ExpeS8gxacWid
Nq9QP7WhXHLj8bQ0BvsBLQtY5FhzEJwQlc5xM7jCMWkmrukKDEoJcPXcLrHV2JM3
i9NvEIii1oVkSTCF+Hdcv60qH3oxac953U+Z+2BeHnlRxYbIaRoy4hSzf01RLUJH
q5dOmMs64xuRpDYPnG1fY8mp9yMjOhUqv70QPT3r4P1j5puHt6vywkaJBdOtEaKL
DW9b49B54B4rr1tmRWl+5ACj8ZdePADmOJDFdsS+S8kPBm8NfqmXfdBt+/RetRwl
1uzEm8uUYx90HnhwB+W8EdmNBQuw5pYbKVf+4nh1PBr2rm0JWsAdY9rkDrJXxtGk
Kzxv8jrkJP9BKZgwhThwXtHJNqy0gLkmeQ5j4zghhjYrn55oUU6yKgQzDylnenR5
plK6KLItHmOdHrkz+D5JUyQU8Adwr+n4XSsg+whTvOVcOSwRhjWhEore5l2/VhP8
3YJv1tdRU/gYkjiUnleNJuF+Vr6DmVkiYQijXt7eFNMcfXCH1SOy2aZ0gbSMeB6d
YkA6tSN+IFr9IvPvt/mjY9LJl23eI5bdz+8HuC3/j1RyJFIz+8S9fUAd+QpmdcAR
Ws+OuFxrSjLrWmd6UcMAAmL5IS1fw6R4nxWLzzX/JOep/3sEp/TQ0FH2UdhE3J4l
U6EgxME9+MPHkfvffpFHa/qSPquCNx0LSOhcCkuESDGc3OsCSNQgMvFGpTglKPCu
dGKcw3opmTrJRYPvX/QRR1O462BP+cBjwoGLhIXmiIBWT5dY2dKhEmJiTxS/NHnC
ICjJi7xTKerNKhAuCp27PAJnh5dMjZ8bncVnSByLYd9mSUpAseNquJPwfr3ILKAG
/rZKbKB5HIN0+pu4VSe5TCHOFCioJ8aIMZ1JCVQNLY+xs2CtypYItQrrUqquoByw
6J2BrnB1rvvM0z2iksbosnrsEA4DhazZ9H6YqW8HQeC1n/iJbi2e5fJE2IsHBwuL
UprByRxEWLqFh73V/U2EqvMRnqQdw+S7WoSX7MlwOZCf1Xi6PaIqNfVys/rpJuCE
+PlaOKqasu8bpDLo/zSWK5ysMvIiQeSwnGEklEAxcZMeFeGtYOI5IAIIwgLOInbR
mTjduCAvuReCpV6dqwTT3s5JfZN7yYRqGYwtnrkdwRWGl1H/DtWSfqOXpMKyaDts
8rwDk8w8D2rI1sEaizQMyFeqT8O8qBryvm/T208LAMNgBSAkxoWMEXTCJjCuT02j
G/tgV534dw065cRVWW3Yjh2gfABc3//VOzsd6McCooTWKOMroiwppJjGZYPGe4OT
cs5ymu9d0mx/9+fW/M2rXVzlYuePm8Zcr2j4aSWhPJ0esff8ZLLPr57Whf0Bz0G5
BioVe9mj6kprW6T31ypXpPGc8gICw6o2Hn/OmNyccX1S0eHoFs3zvKbZWUOwwokf
kjRPFUCyC0NhoMZXWmdqVVtsaKGo8ffYAY1pWzO7I1IbJV5jcuAF34Pk//gfhMGu
Nb7GMYGWzQjkOw2n3hMfkq3aPY5B4AQm50TxrDqx4Wf0R0OmRpFESlsMgc2ptVMj
4DwZlELZXVn3ROC4z+qB/lkdQEOGX3Mvi3xXBjMllcyR/6BI9rd86Z2ohUHgHUIy
yNZ4T3lNcblP6nf7SIrR65blUCaehUmNF0f7sZYL1eNRr5CkpNVbAM+aANdi3ckJ
2rA61Uzebx1y62EAgwPgNQyNoj5lDWAoZ8FPBuIWzu4ngYXJilBF7fswDIm1x3sR
UAroab+Y5kNjRR9RNTdoUu4AtmEQAfzypX3h8VW+5nvEGHm1YLRj0ulZPnP+TUvb
nQhigizGcfrtWiLkdRNA+0oHODRuR/mmszReg48IGKALu1VZMfnHMxKAZovW75S1
QJZkfh35S1kDcqnjdfv+53g0HWAIE5a7ogfDsG+Po/rgtWok+HW3nGAn0jRPkus8
ZXoVDoa/sy2ZCLOK9cRvPm1vaZkMru5J+5lRY4k3rin2MucxDPIkpv8xP54OOJTV
Tm0L8ckWOlwAdlRPWUpPxwqKRUF3FlOhYvS8XGam3f1VPozldOAdijWOaN1xQ9JB
GML6cg6yRnCCfkmdrXq6RenoY/8MRbsdDBPbEhBS+jTMrx980ageGSAGKG+hgkiI
k2I8pfM38Q1XOO1+e5cUdoG/5Cg2RmrUcQKV/G3Y85jnXIMJhqezm9hlFxHj+CwJ
keojuO5f6MRUE3fvn2k9klQvYJmL5iFq66391rSNWYxWD4xD0PIQK5GcXlsElSZA
4XEobdv+1Rt9R5JZWEfL3fwIRH5yLMolbiVHTnFPIa/p9NJIf/ln8m4dg4I/8axV
xBPLPrPqmSviCqV2QGs/LKRy3pZlWUodz4KZZh6IBvEhZmPJlzqAhra+mbkiB9Ur
SmvaV/a6438VgIMnaQfEgsEcLyxZJA/U9zKyZ0fqv/a35mZBQQwYTAuRxxsnMT8P
6lZy0GyOCwnaJXGJwPvehb0Z1B0pXZl5mxwwIatiMpgt0wAD6OKj9iSKWjZ8si6a
E+Tk3h7BAL8If0OfxMegaqlNsdzP4NDLxwvBWTtluocG1iQTAz4V4nM9vN/lZX91
AL76acrY8FfPC7uwfLacaV2Cslk1F389u2PtuZ1LZ3VJW59EboOmbcaeen/YHbeu
hekiCBxXP2z9uzkIh2Q+KVNLiYZoH4oStR/vtZugJefk0x0+TnbEwJaDWRGxzuw4
Xc10udIpOwpvm/X61T40RVA21N2Q9LEBOLoDKxxyUJK8jyOsi4Af2+vLmrlcAdq0
HDZ5EJq/mksgmvNH0lmOEtuZ2mPi0MRU/ov+hIcsXtMzICngBsQ3cMm/KVtcaC0v
sFPvk3LLz8Wk+tYQcAYusi7p9wUIOn4n2sEdN+YvKUdeU9llYdWUk1CKvE80BhOg
bfsLBA2B4YpLAYIp0EJlq1iEKujpcMvcF+s3EWa2K0cLY5mCLZggDywj4jtvj+Hd
hXANcDmcd8kGT9bKY2W6B6N8mVKaS4GVU+iyfT21eAeg8j1/FavliVVeR1Vk0lDB
Z4rdiEwUrVLCUbwqOO/Ct5p+fxTX69sN+Hgd5qfDKdu8CoWqtTnGCE+GZZbgmax6
PT5pGMEekHWjwnzCDq4KoVQMbpRBD9Ez/BRbJprm/jXihcULcr78clUipXYnctOT
xCLwGsuyYLNDb/LzSV1j/f5/hwjO67KSGsy/IDFVmKTcjVMPOL8WzNmky2eeFz2k
5dcb5BYJgMtBXJDJhygB9Ns0ZEGPFuBmAMmrMwP+WMP5KgHPOaVwQxSFUTtmnVCN
azQQOGoCRE2GSl2dujXRAIGov2G/IOHAdrLlDg5MkOdN3Fl6Vj3o9DAH7qcVJsnf
isZXo2f4TvuY/rZPVs2UIzVZZAUWt+V081m3nc+TZ9PmUBCsyY6Hh7DZs3N1wXpK
Lfp+y6pogCsp8GgWLof68Y0Zz3aXOn+8g8btvz7YEc22qz7E1i3ReuCz/8K+RgqC
fo7RcHw++EHjpDcVaUFgLK8CAK1MUaloV9Y0fV1yeXtW9duhgCEBhFMFGE6Kmjct
sREIcBnXPSuDwo4hhcvmWuIni0MSZ83YqX5g4nIsAdK1vz4IRcL2J0RXlgBFqGmB
ol+xuGlHGZdFhIAsLcybzetn2nFvkyh6rEyexKJJs1uCtVEo6uU0XHtAUbJMHQgk
tjIttL7jFZvyoNpAvN3nAu+96tHs1/Y1DrUvAHOZ82LZqLP0surc/Tbk/Ai9a4yj
WkmwlapEwvJbdtBONAJa4TB5mBlt4n+GSzSnUG5Ur4M3rpbiRijTh+tictrONr22
jBGHqag6CSfbGuIPo2z69UtTyd0g1fmTdPx6WLblXj21WTutpyqXLpXY3HVoKnvy
76sCAzosJ33AT23bnawU4x8sankVcTNSU8vmO3L+ZYtqrjLJ1+OMSyYZvwtnAf0x
enuNMlzsZcwAgi8zQnf8QtnVgggg35urPEEVRVLD2qLsqdT9Rbs5+joUjZVwDaJH
uJk444UT2V1FSkVve3VifSLhqPTx+r+f+v7pT9S1cRMffDCdmUziyV0tE0nJFBv1
6PKSWYrjQBJqRYi1BQfzqLXzi/tyxQPgSOqoCLyrz1kR6jDO4ZOx1cB21VO71GoN
e3AkPCPu7PLj/KEmpunK8yhTWjuehti72zoG3Dpzw2lNbA/YjP/156RspAGP1DXO
mKBxgUOfsoo9U9sl8u3jVD9xMl65Cbxcocq+cimAcCg6wiUnSA+7cz8Hji681y0K
vnt/uy8Bzdt+lR/iGQMCe5Dow4WP2VJXTUx4iV+kzol6IN3jPDQwJDciGCbOoGpY
DlZotNUhrIAUSZ7beFO2VF8biheeNhIAA1p7BVZyI2QgGMJ78lfF23ncJF1N11Yq
S5/IYg/4CeOE0dbk3oG7G/v5EnjtYwG93ncbdmmLq5wBaJhk3JL88jXjD7FCLj37
e4yEqWpqD0+BnQ2lohsofbvy3ZRlu6/pk02yBu77ovNkRBlaHlWXK2kXZElkM7MS
TPS72p1F16mRYNJT6J52enGVVT7F4ReZ1x4cFlRCN/npPhESQFVFIIECp5kndxXR
lmbna61ppMCHcOB/C/3LQio5MocSgTq8TfQhLNVs0VQPs9mrvaKC/DD+Mry82GGG
Y8YH0QtT3yJNY68LNs5/aRHfznwTaWhVtdTfyHLIK4aOBxFQCdeyA+L8n8AU86kK
eKZNQsv6jjNQXKBB6QUJ72+BHULo2xYq8gjofmX3Xs9XSbP5X7BVyx/1lJgNflRh
Ck/lIGaQnFUySW+/y636z/h14XtJ7rEUGiAoXq2FNLYc8TSY6WeBTtdsJxBWr1LY
WtsKenTTj8CVdt8cR3n753uPkjarE4/lWR5wlEy0+F2G4lXbSdW5inECH00zs4nI
3UkaQWgLLLUp3TC5OqfaYfJ8qq/xYfrUlSPH6vOjDZLj2E1qpAlqLeQZluLCjhEz
yScsoSoGycbBnGMgkeB+I0TF0yHemHDaB3MjRars3LqoqOLcHLn8wgfofmOwdgoK
3Bd+V1GaY5fv39XDtbEy+7tntL7ZtCAWv0tE4rBoOwCKtNUDvOhxl/obgfrkOYGx
JLgUbrNlVYDhzzCxWKsLo0YMvQ9g/CiKWHB+NNlEh1FmfXtK05URGKGHgfq9Nb36
9NnZ5TX002f78jwexrDb05A1UGqoyL9HdKMRKIer8hakIUF2uwQ8LuQsG2wWuasY
4NyjgRaIHBpfNRwSt8nptue9AsozatV7xzr7rGzLs1rmqU7iOrS6ychoef3J+RQh
qBypuX1qPSiCDdTaw8FUgeGSXXe1UeyPJqaFavChsYU8q/+F+1MEuIYms00moUsH
jcD/bQkVlE9xU+AfMGcgtuIIubFaNJTkEUMCQvzaoIdE9sprLrEHLDp6oTeN+nMi
46rnwB8dOvSUldE496VViZ4Ofo9+lTzZHf3l8xABU43KlwqA8MeQQuIEiYnRksBi
GXfI1xYv3hPDEGB49OPr573w+FOV6aWl4nDKHFnGZelOkZXM6b2EcOxxP4zX9Pgl
AHqxxLgsLZDRmyAOPNmlboV2tq1E7LM5L0ijjIm3ZUozZTumcnviBa3Ppjrzifc3
p6nqoHk0g/U53A/43idovJePJagX5S5BXRTxLsPIBfxkph4mQMM15PQ8NJiveeG6
W+AjZ5C6F+vQyTzB8NS3FnR2c+4tycWbLKusqwuG7MPNPNBuoMrzPRaO98cMNfPM
Q7g/WopCGhFhA0wqPG95TUlF84yK5Yju1f9jE2hHKI4HPQ/zEhnlMXJ/EIZ+dhYm
cwWLF+a/m2aKVj81L4guvBslcat6ZQzNHgBJaJBYexCG7Bg6dTHwzyoRUA4G4xl8
e3TvMsp3ctAOHE1m49x8oB4jYSA7qXo7rhFs7X3tBfanleXXgz4E2DvfsBYU4ZSo
dCu1jdsPz70KtMj4W78d3OpFdqTedK2sWaTTMfcyXOG8UdU5b9IMNTfdTfdjWdX+
dvf3yJEuuWHm+WtqmYmcYM+gJ4gxb7sAUo97AI7TE5ML+uGNud+4srSY3Gs9p2rD
SL7qsASIWD0dFyJHYuKt5sEaOX3IwQl5lvAyN8XYLKQwnYLLcKyRcpHJ8OTmrK4x
rjrzOt3A5EjUPOMY0X9C/SP/1+Zl3CCQjWmjG/iuAE5oT7iZrdrj6QclhRQQcYv5
Ktm9RkU39TLD5DJP5SX3NSy1q7WAkqYHGJbQ/j5FgkZnOeTVB15wsYmMOqR76PQg
e04d+zXRWyLrSIykAL7Q98r4aNkGLHtBGpw0w83h/WenQLIdDXGWm33KJPfuZSDH
YtjPnWpiB3GYRsKqypAnCrxjbN1yji/jDq14Dj67Dz70+kNZ91KYEgCZnUuaeRAs
WzD+pqqMo5LMKQrmEec5OvcjObUlGYy8QvrA2SIXWp3YAm58A7nkYEPGuXOTuApQ
x5CdJGgMqH96BNNJ3x0kPdunDZX7nns6JOg4ZB5Ud71CBjKrDUYc4D8GHauA7h8w
//Mmgeduwuavp7Lm6wNzvJNS+/4A7QHtCSTen6dHoOfSYv32SU2x/i9bp7aOgUsI
cDFdKju3f7LX6eDLQYsuAsuMGtjJYpjoDnluFWOgXWKqUlYiWzsQYKZfdxzoQmZ8
VfxC9ZTMVaO75oVlWEKXG1DMdhkbMPsmyttg43b9oNreegOFywSRFsDofWKQezVQ
P50MNsIwCJOA6y20F2GFNO7SnhbBS3uR6SlEIcK7MwFUY/s/GPQ/sOf9wBmlVuWo
aYgiOErKjae6DI4/6MmmHH2ZJdh/LTmgyOqmfNGpFKXrgTf4uaAhznFuonIfwxWC
If5TtOY/gPHpfGc7Nk55OHKvrK//uq2tzLxlH4mqT65cS+FoOwNPV/+6z1UFHuw2
m/f5t40ncHzDatkddc7pOfwNJH5NsXXkfjt7VhkEmgxVSnSztvSD78VTIBfNtFY4
qEzeMylZ1yddNtztZLrpEuGTXqDiB7dItm5XS04TTRyF4WJakS6hoCgCwmJJtcHo
2d5A1AZUWE4PWela05bqaooMlrPObblYlP5LX89YtrQ/Je/L7AQMX/TVQxBOgpii
sgLKwyqgmptj/1skEIUOKVrGd4a7nOAmE6kqd/bL3nMtoKVG5+0QfcFEUOWCGdvs
nAUd6oB1ffRzQJJaZBqsDuj5rH6ULURwLroEGPeCSzosRKyFYq1wNyaq5c0B8Jsg
+UflEa0zLA9AY0Xuwr1E4tk/SN1IN6NgdFZ2gEWmcEh72brwS650PYvjNCZjou80
5E9N+RhqNBD7IAUhRGa3cU/v3S4vP4XNjPlpqmncZGALMpbpbHVCozNrm6nc/qWr
N67zH3Sh/FQz3YBrtEuB+rtbpbs30vZFLezIKC4bOEQWk+Tyt771JDwaBIgf8lfW
ZlIw/VLwU0REGtaJ2ENmgBXbiNz7TDlriXxt10jiNtoEdb5IBFLbHDpdHB9o4AGk
YEZ11H08cSH8Im2pMcVo50MSrdRfGoGr4wmBcqBYIkvQL6xLHz9aywe1ESKuzKNb
Jako39+70/NGIoRKcVzX/s5FGtvJXG5kN94GnqdjND//zCUJbw5WIpz6z3g48fh5
F62iFl+qtBr+A2AyKCHGCOEfYyfPf0LVwMkyZ5WCYV4k4Gl16PnERahJWxwsA05r
uXrxVYqSB5pBdWMWrIG86WHhEUwsUesXDG4ZyhVYo5OYkCeu5gAJcoVbjeVciZw1
WOv78Mdi2Ntxe554WwopheNsAtczwgYV+Lua7NyLrEAYnTEtTyfrJRu2KF8vMSJk
iiTzPy1IWARgIWKWkMSDwpUIQHZIAjjJmTuz6ZKNzTVjttSP7GhT25yPeUzJap3O
VIggiyzajjPx+ad0P+ith/cVqDKynWbBRF2cMShp1ozkLzkEzJrEq40kTqxnPJVl
KSxuGhpy7Q6rl0TDbxgQckhV9Hjz2rFKMMgI6ocuDLkl/5S77ObwODRqmx48kHhg
5I/MgLilyN3Nwce9Fvnilosvqvr4J1jURupN546rW8+C2yKicsQZYjge6f1mum8U
TSDX//pQRKWgcvgoP5m0OfO49dQNL/od//2pY892/G4YmEO9zLbuPU5BbeE0CsJh
sbP3UvN04juUJFNaO84n/KEINhDzLqkgauAuWA+aG991Xb1g/FFGo/QXxX6lbu1R
rjsQnutTCdMI6LS+/ft2WaJI1MgbHqMW5d7yQ/rurXz3g6Th7quB8QCgdDnlD54a
d4coVSESqYJBHppEATQ2cE84PM4rYj26ct+4h7E/rCTIhNT0pDfxYAVkJirZ85HX
zbHmPDNpQTwHv02NVp/sq4E+V/EromyPpVRAOOUl/TgFglE3SkKQSsovyUjx5ibP
LkliXFE1E5Y+eznFkPwnDDrOsmrbtCPzG+Ltkjp38vcArfXCscni6rMl3nRVf7n6
79ddEErEoldQMz4Zom5ruIY97U/MA30Ds9LLcz1wl5AYOaiLKFLDKfXHhosegrFW
HGNtkJD7IuGLZr9O8OnFa1KwG3I+WyY3vSrZ/guWgs5b0Ha0QiuRgLBuun7hZiHH
jF11R88GCAtaZOpNKdz8eZa8IxfY5wCoye6B6QXULrhtXgducbCBd1z67jkX755P
gfSHfK3OHO2qK2f35R9GPInXAAC9LOHABis69eWCiDhiwHpJfv7iaAwLHWglp+0n
hzbqfy0oRWwYNcL2uF2t11XMcjuOow4y1y4NxrN/eYAO7f2vL7Fk3EOMeeP1UCtU
HQ+F4v2PvOp7vBYKB/LUcw466+FI5BO5ALUlgaqW5HWXjBypmfPYGY9SYWtU3PI+
xlSS1NE2PUrDofq5WP7YEVm962F1L/O3JVLfREQd8YHiDz9s+UACVMLsyCR5trB6
Itba5PnJNs1Bj3Tw7lk/5+5HbVH3B8lIITvGmOXMlBNrxOPHj1rWdKGDdkVEOCLC
eJBwYEZXAqaTmsQ7FzkG9zHEBZDpPJkE5qa3MRQ5tzvmaA8GSSsa9DxgX6t4If1L
1KyHT+fZrpExGXX6Vrq/rFdZNu5uljS4bpffmoDAdNzugrDJDPQJZ9bmzI1lBoMc
hSb5EgGEpOiP0TW5HpttwJhl3v16M5auUT/VbiOUwoYsB1T0im3idL2n6UMEZxPf
jlqTOww13Pyvswyzou4tAgjTK5rv8Xqi36K/ORu72YxVGJo80FUBxeV7BhkkJX/v
2yFlfUuaTRqSMZYW0AbsRSj6cWnVb6BJ7zGPgUgawJg8XedRUc0SV0aFwU9vjn8L
v4fhw3sFIsG+hXCohq0r3jMjizyFO6NkidMU105pH2HycWAu1+IXr5X3RgXa0uL7
Mipd+xzx0Fo6RSdTvgdiscf8chK+Ku7xAgIEaOmQBcrDeE5CCB61nYLKO9ZXV2pv
ABk5JhWg6fczjLpuEqfYi/Gdivs+kc4j+Jqt2EUF+mrDvK1atU6WdfH8zxFY7w8U
dO6QERZw4gXn0LvYCzXDWLp9SSdYBtHihOMMK9pwlNxcpN4RRxcECSbl6Fr43R1J
FlilAg0JRS6ufA1A2qnJVUyvQA3w0LsCTBDSRDZxbkCF+cSrHYeO21u2IsRWCSJL
5/IoK86VNsqENu2+PimnJxPBLrNUK8noyP44lKyhHq180QrZT2XK79Ia0Yz5V0Qn
9Y28+a5QWUR7xraYrUHRDlv9On11nzMFjfkJcNLSWdtI3RiiDGICwkDoEqw+DPJD
7SoB6XXi+RupCF5bVZRqvw12bDU6buMcfyt+aSR34ka2ByGqzri07cByIMLzRQ4Z
Z8t3Hk5n9ov4UCYu79Mw+Fg5OAbt0uPpKpBe/9+zAQFOESPLmYLDqS6ypHrcYmNg
8olACo1Kf23CDUu0RAaZkqgJjFBIV9IXJ6k6xNoc3681QisATjk/hY3oKIxBaCYv
yYB82W2WRiUshNF/KWAZaNoZmFVJuBfQiwJlfTTeWKSgTnIlc+EIDCVcqhB9fAb+
n5buKMjnVQp7zU2PB8SXXFn7pChjNcrFIG3bDjBJBruVSTohqxIbCZTJbWZygowo
2UWK5ZhHN1AYf42HjeDfbGyrISLSWBKYZduCYxnf3tytCfO0mLgfuuUGa1gEGKmk
C8/7uV0ANqlEJxlWz3bvLldr2EopXjPKipJ3CXZ4HmywBf+lLSOCIL0D8Zz9qS/f
enOfanBR2wXfhk7BKbHWI+0FUcdF7anT7ViG6ul7oX+ili54oRAdL0Zdr1y1lpPH
5sdB/LD5/334LlBhS/tesNBz0US44ttyz1YsnBsKSj9ZQkAhPSiCvQ2dhdwJdOWx
6mUqfC6oMR5CcKCRVnq61TMofQcPbcCZ2rPEtjMmlCE5uEQvppMJmgw6ANs362n6
LEcpCRj8OowCf5c46C19YxGRR25Er0Sqyqhfs0VtPy8vQifJfFP0EGqw2DGZG/mS
GH89oUELSMlF8IP7ZceNNS6OU3/rX5nWQBlAg+GbaTEnxh2xq9D55kkFUObOpCbD
p++z2aWXz8BgsXQLLXfi3imG8sauIxbJ0RYFTq6rp8yGuMwTmx02tzZTtSnyZuAK
CB14sFuYvPb2hugyoCuaq7X8ijqYQf7ruhnSJJ0N9S/GRh7kNhM8Gdifs+SCaADe
EKG9KhNGkHbGiBLqIweKDzOZ8QcoBHwaD8xB2oAXmz42n3kFupS4ShqrLU6OM9Gj
9HppM+lGGctCSop379RAae4RM5rgetWBllIdyIK/uS3k1ZVfmgEIARB6l4krqvfl
wrdz3ULKUpOfx0bpGae8LlMsZmd8r5YsQty6KY2Ba5Kykgg8HKaeom5RVdsZJxox
7lrdMjlNGsUAw40UE9vFzcl/sMKvDADKBO8ZMSgHl86GM/pYfq84/7g5cfZ7SRhV
BCCeuR+AGKpBzJjyTzdIyuhrwSaQPaWmny0mNMenYgbe/fKFVt43i0SN2C26ACMJ
HMJHIty12sGw8l40z/A7zPhaEH6XHrQerSecKcgh+Zy/2RY5c+NmGRqq0AKisPJp
uyakd4WFMjI8IN7nJgJD2IdjRbdayrerz5gcrbgvROK0KqSMkVamKiq8u+f4AycU
qe/WPCUXBrwxlQ9WJpZhAj079NWFxp3JQxJ6GJhWZ+5+jQqQ6KAOzpirMK0SVMeP
841ySmd52/oTL/UjkXWt2GfxTaZntzZh0XumSGvHR4lngZdqUVpHN13O1rkCANp+
gSD1RD/l5a2rEsoDw4ATH+KF8A5fR71lyPH6ALEk/vyJCD5p130m965VUDztNcGe
PDwTz7bt8ddkl3Fwp0El+lwd2eSd93vwYInn+ii0zuZDlN4hk6/lk9YSrPPw2QJn
ZuxollLSTxNUJ3xBUeuAlkjJViOAYt+GaIL1IL3bKsCj63L047F8H9aBu6zm8ljk
/d6eKZ3V/+POZ9VColI1KqzjgKgi+1eBRN4V/u8fdl0EcXg02efnMKX0xa8WsjXP
7hG6HkfP3LCNFamNOMcrV7n7XhbhSd1HnbxyGzzRar976I7nBpG7vAEwp+DAAeep
gj7Wtehq368BqKFha3e30W1BZ54S/EdDhKTPgLZ/aYLBWdon7nIgRk8coESUy3qX
PQRyKNouw9uFlQJM9JwJ89R4e/ShvWnJMgXshlFWbkL5SAICrs9K7M3XXKhc/sZ7
m9FeYYCLkvZ/c01R1/17O6bmYN7s9Q7XRMOqbbUD3Q4cqiV3m5zzp7ebMU1zViSz
DQmcwh9NqlmAHxALvznC2r6amUg1XoLGhZzWn3Uz6/hd/m/bIEKE4YNsev9E+2hF
1hzuriQw/Ik0rUCMJNySl8xnrGU/OjaIotWLql5Edo9C7k2vOM8H+bTORJ9wZqR6
QsMSOIfyewP48+aX6RQtx4JkpMXFqWjRrMUJZn+ip2K4MgLy/nQ0yJpkEVvoDnzc
dj1cE+EU5oUodfkRYorirbj9y6YF7JLpeHuevkNAk4NXXo6akmR2x4kmAYSQikh0
Y2BZ4c8GFvmeLvakQf4IiuXuevrjYsw2UWt/Wl/rHKKsHzVk1/UTVr0szLGsr5a3
UyK8uYXuBi9IHIFyAyOZJmvFTE65QEYrRRfFfb/uYOeRDidqnz8Ml4Hn2tjPFiGm
uDJZI5vq7/crHi3wm0jeIYB3fvfytlnY5MkfOhcIVGoqjn5ptMrdN8L7gDkbQKIF
OdmjJlOyBRViLKTuErIGnEMFJY6IoiAn/nKnA2GWA3US+cL8IjYYrhA1I/BrZzKo
IrvU9j/3Q/4Ptefpyo6ezTwSCflD3eaFUwsoDQYG/SZo967wM53ZDBn0IdC37OHo
RQLVmuk8egc/XO5UWZ+124sJMIkOdLkfl84ESTtiezHwDDe0v9qV11ggRNPGqLXh
pkd5FoAYk3qs5LuK6P7nrySTISzLMromnyNDRbruFqbGrH4m/2QqYei7erh9XCL6
8G5NSN4M2QBQQ4UYZXpEJxSHD39AYwuk1Q2Vv908kCG9p4k5xT91uNONL8aOfHfN
UDw41OoGdw2cBjr0TGcIylHVxX7kmja8pDcPg3PMhBXSDaB7R+OgTuGrHlIk8lEE
1abQriofgUx/jm7H+2a/NTvsZ11XdXh8BvfCAzO/37c57YB4Qh/hVU/JGPlOzqHW
WjxFHg9rcXg9Gy0oPnySWX5YwlZf1LsLTBPnFeK3nj8mCU8vS//7549/AToLXu3N
/Eo+cBXVKJbCtyI+Jp9GDMCiqI76q+2kK4wcctpfbY10b9RWCkZpJS0B/nypTOlu
v06ZxtzGQfdAL/xXNCdqLq93xqovF5ek9q1KPPVylDISiI0xBYi92W9U7JoF8/TZ
quyTYuUh3gWR+amEYQKcpEZvrKqQbWeZEJ8Y8TGw3sTEBQrSh/paiFrq9uS1Xzo4
/87YyraA3/RnpaI+8Mi8YgP5SQO4HtJt3MlFL+zgnVeAkxfg35JX9glf71qryoRD
AvXuUvp49NMHv1tvwWjLtIfDwfHH5XoRFcioIeEqeNBnvRxx4OwLKoaWeWJsEMys
Y6lFESKwT/6PORrlSwvrzefwIeoqeQKm+Bw7XZLQS2K/ea+nFTPBtN8PlMood07H
fDwSepAKBTfcjHebTP+r7Q07qpKXCqvv3zgA5VUji0UJhg5QcYxQedl72mxgNknt
YF/U2ZBDw7y+Vo3ArkXnrWlfEd3c0kWUfM5vckBUE7+JX9Cvk10wDuPwHxfCigD5
JHbYmy5POCY0pbV6ijaTA50W1JXKnwmsUH5fywodtmVKudCawq97GdY8qL1vgyxR
NLy1ChmIFD+ivN+fXZoiK6NFBTGWtda936mOzAUQHthUwvy19OxzzI204v2W+IYs
K0F75Yup1/Ng2zAUm46nddheFdZHzcSUu+n9AcO2rw1+BbPmliKMkkFAxCspRNLl
I7jkyj590vBnyIde/SblFsE+O3mOeizr4WFTT5JM2WLvRnaN/u70v1TJJCS40Vqv
5Mc4NntGFzkBrgoAZu8brCDS3MJbfJAWS606h20Zk+xUtJidjIraxxD/3DdkB/93
t0VorgFHz0NaPMrLuYQxQSzerIP7LcGmkOBzni6PRxV14XoCWuN4BBi2DjP4Tauz
93NZORPeH3S17y+Rg+XG+fXyY6gb6huopV1s9vuz6IiSKJAsUD/KA/ohxgbCtINa
GWcUtbWxrpvZtMkjJ0ZESyR6qBHuIY+4uLEKS//BeH582wjQpxVZP3YwWthb1qQv
83ChU0ntw1oN26ab511YdnTwKGfOtf6EhFqpV7s+e4xkuHRV1QaThMEbcCoAS3Z7
J+t0amvcV7avl+gqYq0eEnOXOms1d4kQO9hAa/fBVYFmqxYTJVN8BUW9rR7UcOF3
zAdKNrf0xcSJAS/vDJ9Klf1OmouadKXPgkThkvndGFxZhfVJxMdvC7Hr/FmwxFfo
Z8aHf7pjgDp8sVqwHKdXOejgpKkB1ajtj/KjkdaPN5G7zYyQ6AyP/4gja0ZgEJgI
C0q4xItx197VRsaSjrHz/nq8G8Mr/20MVRSF9Nzv1d2p7zDo3FBVL88zR3McNXS+
emyy3/izbpYzlIx13TXClKNVyRqA0eBkKfZv/xo7SCjjxcupSwj8Yajf1NuygwmH
wWU4L90CigAEn1U+EJNhHzRGSmvJv1t+tcWgUnbV9MdV8+AR5rFOUmyzwsv+yhrp
Z9InZsCdvy/YXR97vT35MvDkiggh1rZIEv1bQTa6KPCaadobIc0mLgO/3rD/2tgb
7nBhKMQZ8dxJO2US3//P+fmrSG4jwVMKJAWGIddrFudC8HyRAjcgwkwCvQuwU1s9
BXgH0E3m6QDarPp2QR3VxMa3iQ8HbGSpwEv/6ToFN8UUucCUIQTc50D5WANzEakE
apJdema/NP0vHWyZpzK8qE0fd0NkXhWv6BkHP9adCDl0YpRxrQlX4HWND1ZLR8k2
PCGJh/B6rx9HZeZf0FhcBr+qIPe+OmUjXaNTpORu7QsohnX7Gm38F6IgrMBtibbQ
tv2xSaldDWQFoOCH7k4odF8zYVvr65JhpE1twiiRwRqk82H+CZGjRlMaG3SUuT8M
vNBzB/+LBgN8Mzx9MLNioqaq3iVMcsmOhPpqyT2gAqHrCNQXpUKVTwgzs1uxeHiy
uc/bZN4Pgv/HyUaCo51gUA2mLPFuwj2ubXX6QvTpQaTx3S3AM+V05R9hLseh/IxX
853KKcmSZMkgd8oXQ9M04fz98pcDVOUgzA+0hQUNGN2a49MfbuuhYX6dXOVUSbPx
L3yUphg6ic9TerLjPW+E+OyIMjuCHSyZ10g9rQ2p8fML+jdmkMRI94D5ok2YoKLA
S/R9aC0jYbSTZQ3m/UvOWk5U0mC8nHN2Y0f3aozQ6AZ27jfZYOPS9JVuJZq+NoXA
HuylIHKABGM6FgjNjOQPrLYtMB0g+/DxHSAgD/dV88fwLqxMat9n3aC4fFyRkJ9U
l+EuJH115N8WiKq4TInE4QdHAPa2WSKQa5p5z5PvYb64sQAJHLaVqwENkN1vIfkg
UPRtR71kzMLeGlUCHueIPTu/UxqVLrcijXAviuCjXjC6gJRQB13kYv+ZP4BbtnUQ
pS611HECp55WhYE4bUS4vlFcFHWJFYrlXuICHCRR4tEvMWppJq0hjng8HCc6iMRX
JlYFgLCOupP0Q/XkiKb0gwHOEU29H5sVvZTDMLOBpTP9yjztUVCJGjUiS0oSkN4Y
xLEmB9BuO62193LrfRbnb5ptCdI8Tq9puxcJWyrdjFp3QNsTvSlHCmvGCps7djH/
9WLLuWpKW9hv7D/smw4F/bj+/LOTS/xkT7LxPkAJoo7Pe1L6ViKp7kp8ARxJmTVe
MPXU9xDKT+de6ZUyGKEz0s3z/lLIXPHh3Yu5gRNBqcM8UHmJvchH51UStFCim/Wd
BE15aPUSjm+xvRxNeushMbQnFDUNnWnM+oYUSY6yzeUekTkp4T3dtVVv9kaTpaw7
4nHVMs4vup9q0Q2gLQwbt0Hbvqup1sgFSQ/k1LLiHeLKbr78c9c4E3lOw3oWj0IU
vWCxFvP0QRRe3UhBXYXNmWWy53UX02ceG6RF+SLiUe/MrxBnQQGaS9AB1j1l5vqR
CBoz7oE00W0bAEEBQVDOztdMkgQ42n/1Nim73jWIQoiBXnK1cKET4upWDOxiTlek
Crkdn2OlWG0rloUyf5tycGeLlVocwDvPQggZ1mpbKBSu3BDOP/fdQvoTZ6cSGEdu
cvQjPjGBg9Aqvxrc3OSUCjWNpodBrY3bld39rZ/b8GduSD1oC533a5gNkqaKHbe1
Fsxauy/RJN1hSAhidh9kQOaBCcm39qkas/raXA9nayPJZQflz55fAHjCiVhDsvLr
BHB9nXMak1rw/09nFNuCAnLu+iShRXNukeMXCU4EZKdSATeDdcscqERsyzUNhsap
8VAHVZEQvd2GaocW6Ejj/uMKW2zN5y9j8j1ZLLMPuTJxTZ1iOELRTx7smq8lLWny
BU2kx0+liw7ppMh0t7xTFGkT68mAXPCRcjJ9cT6ZSLbbM0x7cGpwRAy/SQiDvAxK
O0ufFWcCXDqv0u4SyjXbj0w/Id9OO1+EeRYnMW8zqMTk23RuL2DS1MSMxCm0gn4s
iIYitpgIjE3hOr+c7A7a1vVwGIXVnCGrlu+yCKt/7a02rcGbj5bvtWZPXdocw6Hc
iTeFp4F1veLYAAlWOg7dy8kHwVV9pkFfCJ0Y1Dq8rZ6wBHqJQhjhpT0K1DZRYi1y
mr5qg8xbHfaFTbquXqgEDXoV9aCcuRVzQ6t59hpbt9l2wT7ZjbMrYPoO4yNiM9dO
o1RcC3Sbkie0rekQsgbDRYJ9CtCH9Iph7RWo8VM8K0LW8CI3AgwUc6rjc+e+TTAg
7kXEYLBA1WqUllQZLJ7QOEYOoSRUReHoYuyqxvlKcpmJ1ZX5w5iILO2e4DiIB/A/
6ZiSHTn5kns068pKXePznQevY3WAKWiuxN5XnJqHgpWMQJpABvHftTBIX81zzvjS
aAsI2Q5TBIdZaV7OAW8Mvk5l4zyqwc4QVxsG+twXCvyP8HVoDsWxZcahwI2kcOiL
lpiBCa/4T38kgO2gLEyFFtSwme4enoliuWM0dwuA5z7UKpvr4L/Vxw7wyocRJx4l
CkFOIGHfScM77QIqlzIjjuRgPIN8BA/T5abFh79g96swEF/JWTCOKBhQ/+bZfbb2
6Ua1B0y0Uvu8ySuRqd05dHehPS7XJCscO0TiwtRed84hDaoSQY8514sVTu0XHfTP
gPxlhA2EZGS/ejS6UJpk5v6iGZXmVgsPFPQrmw85Wf/9C+cbTAFMnRhyjAEmIHOU
OmS/8fbCVQPqCIPPESjk63IYlH+mnhuy36PGgbvUoqeT61QSMrsrrW92Fe6QRE27
LswcDbKk/f0opLfv68leumKRi8JMIwF0ui/02/oP6h8v/vc7P/wIRfCyKBD8gJNN
afQ7sezzdx18hAsN3pi42e9H1jdO4exPXt6NcSAyxYDXTzhquaIG0iIvl6z/Wg2Z
7O1A87DDPWuKChtet4VyYjV8yzen4YuqDBGUJOaBQYMRkg9SRW1EP+gqj6fU/yiH
l6kquOuNvtxsYSwnxRWJe9rDQLyZAUdUIe5NXmGP31Ifr7MCC3xYpW3ZgcjH0oEV
0GTBHK2IQmE6ggc5/JuCF6exWJk2Ly0l0CLp+ipy5R0KTzRhXZtoFPwaCfmpSOvU
+99hWf3IWPTogRL1K7wVs5aCAyrgYRkMjRcx0csX/uIJzICQcJTmMvbDhl4V2MbK
VY8WOOxdrLXjSd2yuruAMtFYYqT/uTAExC7Q/AAre+NuBzyG8Z8z1J0zx4v4/1pp
zPfg4lZQsiE03x0OnB5ixRp109j3zh4+p3f6vkqdUsC/0h08onEEXR7TeShZtgCk
11nYjF3z+/z9ebUXmbKZkmjVU8p+4ZhMnlIQlom9NUSiW4HrxoB8k0RXGB1fCHXD
NKY5N4STkXYPy7F+wQh5e+K7JWE7qN8/xx9ocZLtunhsS0ykQObv0D5Qzy5+t0qe
EJ/NOOAtY3XqmDoPe1M/n4vYWxkhFKUyuaP0be9a7axoO9V+AmgY1pFN/YaPOzug
Ib+tYfTo1u3SasqKAY84HPn39dNDYeWaRucSD0sJ5iDcrdb/mboWJKbGwrAe3and
4Hi5shWMFUGirsMjGVeL6kUT2ZwwwE6/RB22RHB2CgObXfMktVSJoUGUl4t51PFy
MoRJkbTpYZGBiz4ugH6QXzfoIrlDSPlUu8342SnwgoW950kitwKq0zZXgmLxAn/W
JUrAzCCwXiuZxYqh0jVZtMW8n+zoQ/BnY1LNbwrNUuFhFiaV0j38k9bdh/D7PPSs
FlxBcWkWPQ+k7rhVlpiyLrHfSos9JjTLyTgpP6vAciDr/0/oqnry8z97oHTo0NHG
gHMxTx6v0+v851o5OtLB0Pp0FlW1A//ccz5npkM0Tx+GbNY5PQJAAGCemXybzEH6
K8LIq6d8DesYrl6JO7ke1qfHzY4pT9MWiEkHHwehs+ynxcYbKgapbNapbBVYf4D0
4YGkvyxp3cxKoTjCNTbhXj4qLTUQFUg9oyTQgnga7c2LOQaG7pyLF3yoA5Bbhrl4
nlbvMZxJWSbyNO3+bg3D72GASzZ2s4G5PkxCNhOqMjBAQG77itVgwmXOlOWwBlCB
VHOu1R8laQwB+xk+H96pr4e3hM5adVbW3ypwbtBBuwwI+P9rcQVvLYZvWzOUcP2q
yRPuJ9Tmxk4R/E3qiFM5DZ8AVPv8Co07GS0INWu3IV9hGWwg2u1QoJw+g+FDdUKL
UBBQH2KJhQuu0dZrclTkNOwz9fbHEvl83dUL36VHRP+UbhIlGWdmBCkbXRL9hjg1
cgDsOPnKz7fiSbg0a8h16xf4atRaBY7xxy4cSzqdh6NGHuOGGtUjuslY2rBalOfS
/7nXUl0ztPrUrFHJ4mKLq6G4A757sSqPmCuv9qyk+gOXv4pArPCsUc7bZ2U/K9Vt
OPnvq+6vtemz4kV6ju2SS0PBTuGG/w0lkTv/+qHzhertYBHEgD+w+Get4CZHmxR9
IwPOr7Qt1z0ZaFxQt+9iLY1eI5eQgJJJv9M+ZfW7oYAffsqf8GjDdALuR476umf8
dz3CZAjbpy9YfimdbMwC/TEmd9P/qhCKZHnIoHUa6OQa9RkOJmSFqnWV5ih+OsyC
+B7GCgqUcPLGmA07+BL/Pq/K5YB8bx/6F00TgPhPp2w7zvAaAig4SPrH3CcDl8pu
bamgqN7Lg3bFyC84lNtDF1DsPNnU2hp8hawGVHSsqBY4S5Jj/gMELOnFeUovVnDS
Hh3opFvjYMqASbO+X77ks3umlSbHeqXUhTvZWAnaBx6cb9o4vHDtHDRstDDdg0sY
FlbQF7pMrLDj3D4QW+rfljQnKTjZWshNsJdW5UYq2+GRmxzneuPmbVUXoRoIBd8R
y7jG0WdrJFLf+kTsZ7RSz4CkoKRRAsmyINTYkl2gYYwDJfQFA1oCNWNirAMHQpR7
i6rBtNohrRgyp9wGvuEGCQu5utvYkGwrBwQeh51v1xl1K+N1s3QuV18uSrYENtvF
I8XXzyvUl4pjuWe3TAcTw+J4EGVyMO26SMIHnXPhGa7TlwtDvJoABWnJ6FPPgYP7
YYc035K8ulvprqoJQgVTUzPiSpRkLt2/wDZdvyDCGgAM2295ijJ50VwTWDdBW0E4
b8zqk/3Q11TZj+LxJngkXzFtNApf1v/K3sIGE/LM8c6ZG8fgJ25VU45UgGWOZcC/
Z9uFB8e3rgL0OSBbVLkybuIsvs4z1TeMDxPYFcIEiZwdF62at1wmkaPDcseU6ELE
+0C4jyJ8M+1bb2dd5Td5tLlqYyJG6MYa9d/RgSKaas1IKZO+hGybFV45PovvOhQU
zWQon+7jYiJYaytSDNdKp7p+3NgiufZTe4dVGM4OoF7YiM2CmAYEcbPDPeKUFeaw
dUTBO6vjfEuimM6eZ26Trtwu9pj70fYUtYmgb8hb5kya7elCgluliBN8dYiJIQvD
xs2XnMzn8il/Ed9L0cXkLGtQSpyuI71AqY7VIGLPL9uxruuxJ0di72xsYgXfwhAj
UMx7aG17yaqJG1rtjNn8JbHdCZK/OIL4bA/85veNzo3Xgs8uwahODMRwr8mQ/gZ3
SbUeGN6xFaM3SbLTC+qYQeRQaCTvlVwM/7gZ5vEeomQjxhU9uQpaZfBMdTWqpZOr
njGd5L4TgUWgWfPS41cbiWe1GJaVTMHRd1CdIxiQ3b+VC7L0nNzr8M1HqNeuwbSl
9gD067h7GpmZ4JtCbPgid9Rvo0d3buq+CxUL5sM9fMGQ0cQtn5raIRWOa6S6v6Z7
wdHUPrvMX2JkvhfhLn1QcfVv/bT18H3RiOhhFrYgUt9kRsibNr/uqImytytGPSv4
oWmJOItGQ6voA7zlYSIM0lFoc9cC4JU88/hVZsMgHJnA6fYHt5uhRv1Nxyx1fA0D
6h5VsyDz3R60ARC/TkRSDliIMbb++wSbWRAEUOJWUjcbglf6KY6v6zs0I3V+sJeN
NfgzT4kiZZH/Dz6OAm3aUFmH8fjOyvVuCgNdFVqscvo894iVFj2zJDoT3EGSjenE
ErdpWcJLIdPHWFrvsOAC8QROUK7kZRtExp2qTS3Uef/ujJC2UEb6TwmqgAkFwY1s
75/+Z8WWtXPAIuEJgnHC5wgd0eIUcq1FdQsiCvu8SnLXg1jIFhetQRjiUFKWb8rd
9estz2ogfKCd+Un0lgnY5TRtUgUMEfPbTGYbrOFX3amknCuEFzZFjW0RaCAy4Pe7
S2NKZNZ4Qg2hCbPBNRrDi0zmQHWWQ0jvndYS0TZwHFiSMSPjSYhygBaYrcB0387C
ZrJgRkz0mWw0pj7tIPyqR2jbsTdLD7t4cI1Zgr/uPPutxQdlfvqG2Z2fwYQprciI
HvkNQR/36CWgNYzpRSqss6XNJBLTUturpiRaIX2bfSHzvEsDXb8YbxTo55egRnBD
O+4I61UdT7UxwCxgQUpbPIHseV3yePF1eun0VE8SVbsYzfLtxpDDey4+xyHaUmby
GPjr1D31PlLdOGvV7mnvZ6QFle7HwCmQuBnBhmct+0bOoBaDFP/tfOWQXDYIH734
juzVZvjUvjLKhKLIl85NRNWsD1ungTwS97zpyRZIB5U4vPRB0RHb3ojN3JoR0aQq
BMHxgZDLSaGx0FKqfmLpIBqAfXjHBO/rsoHqwKvF5HhH/c9iuJ9wB1y1uG+LlU+W
+bGPDGCsJegZ2STJWPytpYhcr5hqYFzz+9MaiEpARKb+MW/3LUyrF7l4RUzZgXKh
fd0rm/B7ULlxS5jbalvz0KLrQtQ09EFqzQX0ehcWXyYHmbOaPUYAgxvDy6kC8rhq
Ngou+bvEfWzhs5EYMtV5jGDs8/rHIIpDuPvyhg71jX5XJBVBM4KP502mr57Bo3U0
xOfSBCpqfGm+QZ8adQBFqisMfF5q5+riuRnFh9z+z4y28xLyd584o9VTcsyz6LZz
sNXZmP0uDaBMOz2kSSkb18U/njpQbDGT+emYoTOqO9HDVJAk5qygcM/NR15q7RnK
rvD+X/bMLkFAZL+cP0Et9GM0yIvqRFPmByMisW6y9QsnL5AHPMv0yGFWK2WkL2hy
aBv+QPqsX30lsyU+plOOlz57bjZ1nDKn7f2dmJouOfONF1herJQaCwxMd5QpuKt1
QICbRAsIx67z9zPGrGKViEQj+FGr6D+PsaTZAiyBL9JwGZPKXI9TsZxYhqyS7wSO
3C9iK9DJJtJE8SxFat97JEpwrrIMhL2I3NRjQLvzFlQgFlFIgMI7/o2zeola2xSy
Iqi22qCCA9M/NoPEAI09Ejqn57J//aOCn7FqmA/FQzGNCaxGG/PsqzphfAPqlogO
q8rho26n104NRDvaqnZTAQfmT35hIFBg9UpMHmal3WMrRbFMVIfprJvH531k8IXI
XopQdLQdGxFcnjJw9l/MOaQXr3qVppUGEm4bTSbeZr0D98YADtys4hWw38UFDtg2
ED0LX6H1+nHQ9sU7d8mV1ySQYoRAcSWcJedGHj+uPpkGXiuXnpWh/xi+V5xOiQuG
lOS03m0fIy2ryN+dm1FCbafZBZqolbJs07SzhgihYKR9iqjW42KE4XsKemmxHhzQ
4tyMxgH8YQrLOJ5OJWuJOGXsgUuqHky2oDnyeQYOziRzejESH483bUuCKJsc8fOI
wux1KRUnhiQsgObwQBPbbJpd3pvgcTTW4lfrSkS986ayhB/knEReU7tsFs2d6f4u
VRAh6iYnCVGSbX/syNFh8hIue2FsLZEuWQemRxUzqgHz50Ho20qvqd1JnhHweBhN
Iu5NQ2VfVFsIbTsX8t9iq0TUcxRaEZvrJAvmPLF2gb0KqkI5v6LVBoGWbUar5Da/
gwuMWnndpSxu7pyqtcQxuzszIZwpCCsyb2iUB4tnckfSMJ54fpr5x6jzXUvfBmnG
6hlG3QgDa0rRrzlgCVmruHYYx8gkYmNSdR7M1sugYd7530m2hxvhV16VSpV8dm1+
YYSeyRztppeNrK25fczhwjJdgX+/oABJDX/ky4SykT08WIZUMSYWopQm/jeLHmWl
hgGPbPUfS7cODdTjsp9jTy+KOEIXX3o3/a6SwFFkpyOdaN+OGGEo1rvo+oRTnATH
eNZCRWmrUkDUUG1kWp0Q73ttHunr2atW+WoiIt3SCnO7A/WcxV3il8JsZD1p4u0F
ioH1JqpzAqrbzSmJxIp4+nnLlHnRCPVRiugG/JsnurI6LFzS2mLstZGFS3cG5/rW
SMCpI82+8JVsT0bvsosAlSNrr1OOZOyiUHcTuJdsEk+Nr3GltKo2x7GTD/9KueUU
YWZ7NvFF8AuSqtLv8oxz/RN4woTyq5bgiXqzFV8/kznzWsl6L17w2De+27iG8hTH
xY8Um81h1JbgjQU5/Y8xz986yc7ogMk5kfJuftLv1emrfwEuygzEdd0NbJXBwtKX
wk49p07Ks3aKCWW4YG8VPb3A7zfGUlqriFUZZuWjRdjk9nunNM0dSxyl419OOkY1
58jpRxv5M+Nh0g4tTzwtqkgjlQIatX298trtmKI3/5G+Y9uJT7uozGJGR/QEGTOC
61o1KpjNlF0eF+mIR8Q2Oc/RJGX+Xl+TialqoH6+QQsGxC3LpeeTNkD5n+Bo3VHs
mi19ZJ8XhqD41Cqi7yiVZM/ZL9BHs+tVlbD/fkX+mnvCUBikwWvdlXKqBp0dNdlf
i7KxYBYrWXtaGQHuxyTKlKKMOKOhYgwCr5qlRkoMC4OjxFzBrS3JgFiZ6U6b7tM8
Rt+bx+MrN0IyfU5rXHK98qL7TKrWjZsg156dzXlrat7Py22sogEeZ03YslSRPeuc
wDrQ7yOtSxdHOCXe1nUO+7TfsmA0zE1AqPJDdHngLeBhFK96/OOhGqophibdzkbt
bmopau+glow/picZootHVWPtyRJ1xMM9yf4B1x5S8S1zsX2CYkglO/rPmVk/GAjy
qYyQR0qq2PWcGg/syIGA0vdRnlySmp43I5o6GK6JFHwp3BhsAuUmpWDdgvl/I8DW
6TSDrhgJJyNoDBsxzcfJX+FNfbUbwph7R1b2OxWwjj65/H1JOZfLvCx5X+sWvgDm
n2PoBOKuEboemf9RoYLXADOg64sKuCzThQjZ5zNaKvGX8iQRcG2X2I+E+qLgwKym
6rmbwlt5vGjdMZ0E48GlSYbD0EOjdz+5KOFYvItwnB80cnVbP37+/DvH1ZQm2zgM
LZzWGNgctdyCLvIJA6+1cd3XNIiavBYArHp/yliYLbbiGTXSXnPF5SFQFEwPydE8
hpqt8o3j3/7uf9RJitsab+a+VSJy/PqrC22NmA/pTHVTYQTNvp3yPLFwzOTijdxU
l1O/GnZXVBJs9TtRH+e0VaxOP7ggr9JD7kVhovLwfkJU957jS6bbCG61DHXBTr0/
wEVja14MEnz3nnxqoT1/Tu+ziZ6DhSdJ5BFDWvBkcXccOBZ8w7K8y5Kwe4vlPWya
W5ujHFOd2bDjytdaPlNjUAabYtRlAS1y9dff8ih8Q2oZ9G01whPIml0S6pBumuNP
F7lkatpTWP32MK4OqoeDxv4mzSo4hKQnStQaBIhJWaaNezHtBgQzSNp4GPVD35YX
yuYyqHL/5ntOMoA2S81nz6U1XdAzRmP2t16sbjVial6tHj9K9djsyl3GQWzA5NPy
bOq7TmMr992JlK8s9bZ5ilEMboPtRBJ4sWxxqyhPCSm5p0Ah5pRwKgk16TI3djvN
f/huRZY0bi22F0TJ6p3KZ/uhYnsu8gT3UKK0FzLV2h/Vl9dW9vj7rzJKXgbxyG0q
cPnIyusYfCEgMOtQftowdlSBQObaLIbuJ+ZbHw5R8YptInVo3mIps0LyQL1y/ACM
XVi3wSedFSTcDIGY+V6GWek/89NUyxj/r1dbXvi5S2SzEnXOuyPyapOrpiUBCo6s
HQxewjabRKH6kRxWETTMqZX7yD8CFRU4pmH3/dLyRbb2lvrNRL4SCH2XSSF9aqpm
GV442oZIcmaZpDWF6qEn2pCU8XyVfn0/KcBuK5lkcbjjDgz0JIoaJMO8Kro/1YB0
ogVt1JVbKkMEu3CR6BQjC1iP7OdM9vre5Vt2oUGz8RVdvdKm2kvbGAR1VhXq5km/
BjAyaKus7Ch0FPP6fnvaEnM2C6HC+g/L0MiL4qEalzkvGiAT1gVkIQBNkZPqDgua
oMtmELF1OLtApDSMF9tsKzQQIoQm+g78HDC54fGf4cLeaf3UJRQtXzEfUEqbg33O
9c1p1fYUaGRQmI7Fq3tVlY9ZOoUz/oR+W5q0p5pR66IoifJ7TFF2w5CQ4A/1gxWi
Mf8v0ky3MmRCrs2h9I46F2pfkR0z5ePToXqGuTyJCSYh+As8YDlWJ8YmGNlaS1i/
UaWWtLCQNWAgAkFULv6HJv9uXk/7h9pKTMVTh/oMFvevI75lsB/0Wzux3rtwwYmZ
OsEmw/ITwDwrQbdz7LrNnWOJWbA87HNCgebGTuSDt8TT3mWn3q7SZxeICFGn2LNw
6V1gTHpSfCnOgqEziftuBauun2aBkBxnTlq4Hg7HkKOG2Zbk/c+Gl322EVONxAnT
F04FBy8t4COVHa4gbHTVpihnb+gNmuQb8G/hjwrgeX4h2B/qizcWA2ixykcjfWLs
hNN8XegCPMMqcjOiVXmiCVw6oTkpMBwBi7qbtH6/z1Apu5W/uXiXigXLQ40gvvBn
M/PorY3s5ffm2RDVpS3XQPeqQ27tvbidE3HzKsruSn3raIUI+MDvdg/WsFpkWxTj
Oxm0AKRDVrRrdD9NzTRxWxwdB9TkVAMTiWjZiTZp90DBxet+V2wa4LN1yShKV9CJ
2+wsbiKy+BSWkyG88RM4rAu81a7yk3lBw/MNkEho5WOVZSm8x3ZHODpXrUMpinzQ
N25WD23MBW9xg/xQo0mVqI37pTa4IbbNMwuuVBCmp7QdNyQIdsHszieHwVmyP4xA
IU5WOMl78ZorDehHah2Xo8sNWnBiijt9Vv3KdPSFGcHpULuQj7vfvH/4Vo3HatWQ
ALGVKPonI2Re5bARn4DBoJ7iAbpI7eD5QDVaNv0yUpWM83Jm0odYQv4LvhmiuKeX
9WJx1bA+I+fgbOIixvQ0KFeZEUfH5mAfZWMiMHeKcbJL/Qd4R2Xq3c0ylPDEuOGV
/5Rh8ZJPXI933B35KmE4KsZInblQntCW6MiQQrtNjsRnP/EQxMIxhrXKuVxSM+qA
a+8dK7AIIVxK8/5cKVVgWdmD7A6U4Rh/KX8Zg0dhDhuYTsYFyuzzXOSCfBJtkekf
duDBv26HJuRIA7l/qODNwGerW5jqOwwvJFx0pCVxEG1S9obz2AAgmWgB6Jf9Qpwj
TMFif4FIWEPGxkM+zl3s46IuKq6Na0bULHplkwveTwIbfoY6SP+icY3I9MEQRzcp
O3idF+vUvTsNNRBvRueTeCHmKx6KrvTdNQnHcbwE9A22pPwzajAOCpmaT6oDxnls
UCdqbW6EcIAbce+8fe9R/v+QA/ILFtH0linFBoriT8gt5e5M7FEZMpzMHkxlTtXY
LMaRARwrBoaMh+44hix8ITFF/2ASiUGw+kAslghoG9VIhlnMOmNxv9djv5Oxhai3
Y8LAfch0if/D5ivAUMDHF+RpwlQEmik6y2XsHOT7EhHOPJBeC7jErlkq8E2l9GM+
5MdZKThl3cz1kmZ3KtNS2Ep1j6QEobfKXrdvF7U78t/XUYlE3FnTTcAFd74IG/wc
8kYHLVONmDrlkZQ6hADwe3FPy/d46RyVWH56u1RY6kJq+07Ta5Pjno8UN1h3MHLH
BHe/GqV3tsb9b+Xp/4O9AisuH/bNvjXQungRZkwjsjARM3abxpQMaCq2LZlTGeTH
FIDxodgo+gorrYn1PQL4gDRJtwmnOmUMDybTlWYlKBa4epQBxYgfh9Ga08Cat9pO
KEzKWmUba4BiMoQyv2B/aspac5yN2uECAwuJaVtu3I/1ss3SB2tnGvo3VuyS8INO
gxCGh5e31MtejsvQZKfJ7lOfXpsvtaGrlIw2j80gzJ3aeGvkGxM3+1HUfi/dYdca
Bg2pzPyKZ/pspJGnHFmkvAcWHIgYb0NaZ6pKCe2w3RC/RffZzyVtIGCnAIFaqbFo
N2kUcuSj0KnJlf7VaCw7Wa7eB6SOoeAe1NZc1ebp27zRqL/X+jwsBF2U3/5lPsdT
ZnUrCz1j6GpyUrypzV2STWwXUnJeC8FlHI8sumZ7sXB3//s+0UCnSlzdpHEayt0R
oPHabOtO6yGDLB+B+wRKdMGqfJtrmr/grQnlL4ZGBHUT85L965kGjI9MVnczSpDD
34rOjjSWb3OQ7u3dp6jlpZmHayy2kH5kEQ6tbLKrTwL442i22h3Ek2gh1ypJI7+y
GGcKYAglbHnTPhS3Ddx28B4UVbz8/HEtNYRYWezV/5HvRx9voRCI/uQmz0mVpTpR
XZKk7ZmAtDbrcCuHSjsKq0uj2zF7Ft8+McKST02MNMGjxHGBknZtxG/mZit5gSna
RQOfZjPmYKilh3KhXFSkYD6QX0M3mcz9I13wJQyWWbm9syDg1wc9wkNWzbsBrcEN
/T7w49/fvW3iU3VvgnJc8onVql/WzqWYdXIVn4OCUWsEcwSJuR/f/tmAH1HTpTGK
RnzHFSVTX5uZzTnrRwBFvQxNHg1zL/t3ZLFNzRDaNlz3+6FcU50XCbAYygrhzz8N
hNDO9mP998Co69XmpG1Z86bnH9xwfZh8UJLBdD0o63AiKXbDkgsuAzmG6w5nrAe+
dG8+W9tOcGTlx7IEyykCdvu2zPenzOIM8L7gp14JA0ZlsoW8vpc0MNZ4kBtGIuNl
QTm1ab/6+Vaajko9P1k0OY1AWtjHPYc4AukCKbGzWFDW7wkhde5cBaiq2KFtdaRY
gighomEAkSKlVSfPW7NYGxlgdDcGwAlHGaxnHiAn55AZCR4Sw/97ZOUGcC38lFqA
3TaYXfkVM3AumkNZCxVEUhAxeOfOo6FxGxfU63hxer3Q1G1gEZXo5DvhnU25hDA4
4V3sj88Qijv+1p8u4m/Y0LeFDV5972CEUuPR46ZA2oSRkLQMU+RYH8xL1YjSlbEJ
vH6WW0gScSAe5jMYgKEQmY2eaNmiF+9ho+e+z/X9eRkLd8xypl7JI1KVw8dtZEfM
WZiEslH3O1SLz2MOnBDP3wM+uuSnRCAlL5uGKKTw5yNMEtGJqCddIXr41eexpA89
IHwnmWb9q+9wKgz8hf572v3Lff1Ws3xEaNDWojiTcATH2uIvAucOBKFfDSfkt8D4
2wmlR7TqQ2Q+8bsHZk0fGkXKOu4JOrlGCuIsDH6mJGLCVr3MU7tdSPRGNll7Eplv
ulfMLHpKO6DWiHx/YqjlG1lqLeGkgWEYxlhmKYk8NBg5jq55jOSFfsfBM7fgHkme
3T4xKcIzvFlWDCGcAhWt18DBlEChDeooSLPj9iQg7dL8yQGVAaRLETGs047nGCgt
/IMTs6CwFllWAehKj7LbBYztHfrVjtOInC/fdjYdayriBE3GRaojdC4T6qdKQI5D
UIuEiAL/D2gcxpE+XvDbkhiIP1Drm/42B0FOmeOwi1wSL492C0gNk/Srydt9GbjU
DmPkCDAsyNliD20PnG3hhORgzC01kssHLVesiYQ8KSnfDn3fLvKpKg/BbLwj59Hy
Yb7HNR9lsmZdZjFtOH/GjI5b1YLzZH/Lwo1Ac5GpfzsxuIcond6Rv+bpQeBBhpxH
O4uxNRMHP+jwCXDdnrXTVhDGsiV8ujzxXQZlGREhcmAe0G74Z7Bz7vdOr7BkBURi
eZGE3dam/bjX8VYSIWTt++edLdwVRIpmebJrmd/4E36Z8eD75L8vzuqC2+D6znn6
OsuJwWuR8GqNbp8FMoRNdmW4D2O7Vhg73HEnP3bWkyUvzL9KkFKi4rEdCbsHltKx
NAQUwxJUh2H9SQjcujX8HVQQo5SyYzuBmS+Qo1hnS1+knPv6kuAIVKnlUXQ3BPfd
m1lZYVnACLkao31F0OfeV92wEw8O0zf22Zt8iLPZr7RAHdxn+Qcpabd4yTMD0H8p
d+WbHRkiOSxczMO4+IG4uTnwzoQywhXK+al7HCUOpggfNA6/dYwPWW612X2NPZ95
fUxPRkz5ZA44teBX2jdAoFjipRAMIEc2iNfAPaiaFYqOvn4GQdQgQvy8F9p304BT
/Zu9YwwW7tkUcLdtZzM2F9Erzf0Rek8DcF6XTlBD3psdjM5NxMNPCVSXqihfUlnW
4at6WdA9dXrm/r4ZC6qceU1KCqo7g4W3b4xtdnfO0abtPrdejx9BRHRm+ZHMHS8z
LdwhvKpFGlPK21Onxfk2FwQmpPO9Eu6evigH/t4t4L2u755tRS/lYDqdbgIpuxg7
SJzH3JU2nvm69QqKWq7ec2Eut8trRVEZZ0rTQqhd0CqttzUK8TlFfLJnrfbr/tfO
2wR0d34ll6K90w9WcLVIaU4GFcupS849jNiKctpNc7Y1Fd0XDYif9Tv/zVw2wJgU
sSoZvL/H4Eugbs2YvBDeKHEhXUV6BlNrTj8IQ/0+1rEvRjeodGDdgLeNUGU7+mYj
nGG2OfdjgklArbkPq6kS33btC2t5hv6CoZE4jye4GO+uVQPie+UrIrkcLUjnsL2S
1nPMjD9CtJhl98f1ec4EbKNA3QnKtx7yiIdGvWE5Od8W2XRXtqfEPXvpH5cwliFf
I6KQ4YFaoRYMcdhjqUWaQxC3672ylYHyU+D0o4Jx7NPMo6oQ+rV7p3uZ8jbHDTFh
rxrJXtTkAxLctUNnyQ5JstXrzPltpkvK3xfsRFJ/+Gfx1d23am/05YQFJd3FO8nz
/Z5DrcHU5ECvL0SjX3P3k6IOQKypF3CG696u4D54D69O3bQtMZHa0OGSEadNO8gK
ioRL0GxxiBfTyqvp7RF2iLjCnfPWLgo9jmIwEbCmLYfjQY4xHmuKnPkPAlpBXR6c
Toviu9kPxv8IAAStvDG/QIDLAGOcIeVV8lIXu/uARr/Oslp8CVovcJqUt08VWO2Z
bHyADdwuOifKH0jLztImpZAWumdk1ILHgZu8wnYi+YYe50QvEWwFuddAUKf3Zbpg
1g2gdAiMbmYGdiWv2IHicCOG+eK2GcTa/gsQrez0CUTnFy43mprIu5N0WZA2QnSl
7XtQQCxWU/XRRqL+Vi6e+KQ0qS+alKbwvb/cSm7vKu8FkLLSY0yLF5+tuyiztAk9
PcXlYTDjuTlH3wv7ScRnz4jjI8NvKFxafk/gLkYn0NlPbOiiOh4rcvcW/Rv0OeGq
KwPkOv1sbqDcTiJhA5O0cCiAo9Kw8hodcMWWOODew+rXkCmhybpLKwRuWqOH29xZ
WwpuX11egM53OfJ+I/P/chBtkigfAoYNFRDeOzqnr/Rcrz0hk9+DIrzTAEcxXn5h
ph6WF5XE7sa0UW5Z0kqe8sN8FMZ8YJMXg3BxKb3N8zYfmQqMMto+/xUyIqaF/Po5
/8XF+CcMihrYUFzfjppw7KFq5c93egnrraFFoBsmI8MuXLGWjaVhbBc53SI2i0tW
xe3nGoMT2pBv9OfgeLBCU92GY7KAVYy9jyZ2ZYgc1NjjGqHqe5qt9cxImu1dqdXo
3mDqApKMfxXvztgt9kGmud4JkwIPJ5ElU4T3Rbjc4K28axL8k47TwuPKcqM2U7+R
ZqlpJW27nbys4v2jrLBWRnTO4C6Mu6A7pdYwAYAWvmQjuNDPrVoo9y0VZ+/xnVtj
kLrzOowUmAIbHBGMcnnkYnL9LcT7ud3XahM5VgKJhSvyh65h5oQ5HmT0YiFluBw8
qZvCrujvDyYiYtX0EmqGloJ9jSLzINwVa7F0hQIP3DNGVbdgJiu6dqbbppc6o1xi
Fd67AlczA09tTJ1wydiVz2p14pEQPRHX5Gw9z2qenHzpb33z/aMMpZhYQg9QKmaP
87/EjnKHE30m5WNRlP0KpaasWRjJ8tEgErg53eBqe+RMoD70+QcfPKYjcrG+1r0w
saWXkG+BqNd30XVF6wdBU3ZNzCXZGziHKGlX34rOr8+lQ/QbB1Eh/boVnsrxTPGS
gHiUigNdvHN3gSQTfm6mSp4bxcvXaAKJ2Xq94jdtRoLgHiLMIeHHuHw3GuiGVTYV
J/9AGpOP0lMfSamwDaLwGLYR3dF1dKEWHyTRMZck2lEZZ4zPZNp6jENCVaYY44/R
6oiepe35iYgravJa7WEEs26e6lwh1FWRKBSYFgI9NVyDug1CpwsE2SRb8HjdiBRX
rVdVXdBZfI36hmRBWR7/aZMwVwUF1pqmLlmpl7cm41Q8x3I3l62RU8B7/yf5QMSu
krOZCzmQVYxz0FxbEKYHDjmZVg3oggar2/mBBMaHvw+QQghp7eSRtH0rA5aRRO/Q
e7O7IKj+4QTv4W4uxhrwWyAdBAAnvqD3cp1QwdS5imhsYIlMLEjKiAdTO3zSWXeN
N+K4gGOxg6EAGW55GrwfSses9T1soTbxVmXRbjfMDcjggdUTzx5Is5/ann47W8I9
LO3MH2ADb8A+HMZRYfMFOWGhe1mh/O/6vDYKTD3WSiRwvkbHQxpqh5Z4a2ijmpn+
QLIQJ8aqWpxYqJXjPBfI+P3ZawmMFXMT93h/P1yRBPlkuefA0ShqACJrWVmBa/AX
bBq4+SMZkeoowirxGFWxxWiOgNWXneBd0TYz5fqYTUit7JGVlGneaaN4cHL1opL5
krOXaLqLfsypP615RMcHUetxEULu6OEwye+rBGOHZljUgfv0wLf0X3HqSqghqFn8
U0wWsOQfVXvDznx6QcbroOgfbVrK2trGp4ssGLG44r4bGi9Ul0h5mC4m8dYG1MNU
yjN+S2iprW5DkJIM0ClMeKIjR5bb5sfbsr4Xwricydl4BqLsdjWjMxkXMQWI0n7W
K30NSNcvQmams3CVa5WSu3B9tGLMxZti3eZKqlLIKXj8QIwYErOlky7Njf3XFIdg
KY5qcIcFKiKKYc11cFc6rx7zIfFqBUc+IVgsAtQDOMThQo0hnc9ht+jwzCZrErQV
XeicMABA/pV3eayfgXDOriSCbvbuYEHf1xFppVw052kYY+uA03eHLJeYz5sevRCM
4uHocUkmDWGnoZnqGQBGvFHcby3ZxYKfUxiWgI6LOCzERNWDJzzClHAZMJlXaDs7
pzQjUo7hE0s4Cerwz/PQCQyq73wGFTh3DiAdrig4qqJu2yxfGossyfIqcUMldNmF
aYBEZhefU8DbYXDhN4jZgq74An/Xycl/hEHFoXuXyrgfgC+9BpQ0OwNSq8GMQmRx
HTzvz9deO5mFU7NAcBqgARAfHl8TC3m80ts4OmHGj5XYqQsnDaW9FgZ8TClgztJW
8a5q6DBBsnwsds2laSkF8w2m9T/z9jrOKIQtwT21fxR7mZ4jl4FOIEaeMJokn0z8
nPmRYLYlGQmwIjyQeyA6uEYmrHhSYDxH4d4DMvvwzJQhGtF4sTN5vCtNVs7tui83
ySYyubVLb4vCmclLJs+FRt502e2RK1VcH3wtNy/Gm2+D1Y+zmzzAFmO2Flms86IP
7jxbUOR6hGm1tgTiEHaaSmTYYMMNIfMRgIm0PLf9ZjuVk75eNYeWWSeysfOSDgd/
qgDJtMCykeLSzBI35HMvbOmnsNvijsJDuOcGvC9zGQhyf1c2VIwnQ4xAanbZi7N0
mB3Pb330DbZq701QaN0UW8kSC1XZYhxArDTblLkEv8ICiUWzQkTqPdN/Nzko2PPw
xHxrbTF/sCghXeOK8LUA7qWsQfYwV7Ggf4ZijMaL5aE8KwbVoVURUwmgn5wsdyRF
/b8/sLAKSUUMY4rlb3fqj/l7HT9KmxOn8VK5YybTYejJShRb82Ih7q4nJmZ1Zx/Q
NAJvo/hhar+gmRpt7BHJVOFx1oK4GFeDz/mKiT/R8+DnBTbz4aZMJr8LP+c39ITX
6a99hVidw2dI3NIfCxY9cunMFAMTElgW1HEpJWHH4B8U/GPzZvnPEq/Pl7B6LGDv
BKoHE4WrdbBpAsxkbQWMWgexEJUxrWSma/060hwEkANBPn12XzgWURalbBKaC7bp
r1qHkzcaN0uHTCX35cwppIvfGsKU2p9xgGuT7qB29w7BPzaUamjrfo1iXlWAiJAc
3YvZ3W5j/DIRwQXKHuxGDEuTPLr7MCWSYzCMZ2R389AnKXU4wq1Ia0vv83YYbPNE
2MZ8byrXk6rEv0dwCs56uhRcQ+mm7ErGQ9YLVO33pg5iTJV+l2xZHJsxzD+k+Kxe
Zed1xfZGCgyit5Ql3LrdjXbU769piy9Jc/8GL78FquUnO2FNnND1w+XMHJ51vpfG
P5vudaGyVVVKaT2UGZLhz2DaT6gBZy/YEUluwKi8ZddP/apgxUvfvFoXsdIHGTYc
a8pcbKAIAxB0vJumIQH/TkDcrR+iZN7oKn7aa49ODycPZ8dqTJFoynvjqo7pWsPT
WCGoQ/95dtH/1n+JiuJsKKhb1Vo5sNsVa3gn1MUavficuXyNyur8abx8CJUSxYxm
pyM2T6lpHDaTxTFKBHDlvb8L9IwEvb3ZMY1N+yIfNgrsjTNojXqxMwSMtf1dg8dX
D7Ayn3wD5CeVD1bHnGaeJiKBDk7DYLrfUsCt1vfaUsXdEIt27xGbvIKx/yCO4Lo4
ASuCV61rTe1brhwTrU/SIJ9bJd+2pb9dSbRsCW4bZ4Nv53EkHQjtGveUR/28eF85
whkSTsL0xcxF/8G2DdUYAg3lfJfljjGMrKNlYWGREQ1kcmgMR+mBCpK2bHdC/RmI
/mz/3M6KxtKyms0oRQ9+lVM4THGIWjsrs8ZddZRnsCmZvyJ8gcG2/4Ii/DaJtH7w
Igwn47jaIe0DHFRJfLr8sdaUaEIE7LsbM1JgDzShkayR5tZ5VkjsGW8jBjPXbh+g
zghJQpxUI6GfEpmi+TSQO9uNF7hgD4dnzQyVB1l5gNZwv1oJxg+z05s3Iaczvrg5
jIyooGQMdXN2n8nEgj0BNRKDZdBrcRioVnbtpEbblH/Tv0FdYyDPdhF449vlPird
fLG6x2JD46uHvOwUlEI84y/2A4izAwNS0CpNZz4DEqxWuAXjBLNYNobjbOY94spQ
ZE3jzhYAv+DQ3vLV+CEJ+hRR68nBvBr8+A+xsqtIaG8trBy49x7iIC8AwiSTsDK+
EO49tgT+aX4agpjHGU8ooLkqjTNJ4m3DY7oXwz9Rr/LdBKUKe885i8DZgrQgSnHx
COIBLELGpJkwPDyoZLqqB3wlvrWQdGZ1IaPY9veNOpcPsvAYkcu/SK2a15RUAqiJ
CHPxS8mQP+mEIb8UNXKcAuhY6wRdkfLSyqiAFsOM2/eIgqvUDXAFKzDsbbygU46t
F1QnVGUlup5s7YFCAjedxRN1JX6T2wga/Cq007GJlKxiW8Aoy5xuxa+dFnWO50m1
curPGtQfcdB3dSQropFZL7/jtm9KWBO9ps1jTu8H6cQErskAeJzamE/rZWjyemY/
OIWzxDv6rSeDsHXtpek1/hDMNp4xp7JogdkLMqCggNpenM3k2MyfUR70EV7iH7om
Q5OfdDzOmlHnZEbLfPaQ//V1FeAERBfYPziyLSh0X1sT/pGrOTCNG5jN4EHln6gy
9NqK2f9+lyfEsXa6L70XM+MnSoFm3132+DptFvqB+8uXIXSXJdmUubxixoHcSHkV
Zv3h5mL1DqOv9IRyPNJsIuEdh6STEvGpvaPfFWkXsCsCekT+YyaCrJm0CidvdmZn
wAwIgCulvEL4pL60BG/4ZTXNIgMjEVvfkTrdHi0k7+rmFlzpB1Ah7Zrp6Io9E2mp
V+C4mt1nmPdyp1j4+da4+dVJGTQFm/9THlyYWDvsKQmQ3X8meWXDmKW/mIWBj458
1k7kVGIwQ+Gne6th97/H8JhFxlIqfOtkO72rTaIooFg/pF35GoE1s5Q8FN51yfNt
mnhcuRQo0ue6blRZ2yjTcMFvltxAKw8ECT+1wnntU8+Ew8G1pc6WkJmR9TA3T42t
b2IvH+f12OQfShJG8cb4jGNpw9Qx1T6f/qtVNmVT45FsUsJiW15kjfqxXq3RpxkE
82coPUUF7VYr5olSiBFb07ehxSBpbwLtrDp6BcBgU2A4dPrglcXua6tVVYZTR70a
GUixHcbbOe5KVnLirI1fhbpn/wyMQXb9mX6CvplOeVrRHNeZhkAe0+d3O4Afpt7S
2G7nEuRwuwOCa9HRORk8peVB5RaPN2nGrLhbV6VShEDqXU8dM1T8c9Vr4kcx/QBR
cZH81chTh02wlous9sX5pR9Xz2Z8rtGMRbfdb+2jmjYPb3RrDPD5Hnqj+X0ncT0L
mNf6ClrnDAcdMIF+pZK3zGdhdyQZvJCFGvFTHC4fyiP/YauS+JyaUuZgaeaFnDDA
rVH7i+6Ms05Gn7dtxVKmrm17k1puvJH3mGZGxg+UF7b3ka25VUgIZH1zMTG56jfI
NqAJ/gvCDneBZV9qiH/wS7rXq7SztOIAfn2h8G6wLwGBsCGaAttsCXeCGf2gSjhB
3+qABFizrEyG6802uUIiYCuL0k9DvMF7Nr7SAcZxePuT4oX05srDSK/RD5pWKj84
cRvHJurhuRVz1v1Dfonfy0UhI7pT4UlFwFxtIjddMCmp1BoerwmwQNHu1Ae0h6AR
ce/lxtYgCefbaziFez7jtRoWv/geEDr3lE9+o13jt2joXe/M3Gukq3uDn2qRWMDx
ySBqHc0SX3Ihk/pa+MF7H+GtynNI9Prm7TRrKD/EwGdLI1bNIvFmQz0Y5+Rx/EKU
QNbcmbGNYItkaqUO7gz6JyrkZHwA1HqPeO08//zR/+zBDHGfP62USRRJM3prCvpx
aaY5HCtuENnq34K/Nf8Yurjh1OsGJekjG+QBv0++WrD3NhK3g+VaFQD/T036oYX8
zJ+7ta0xLH8SBm0TT866sibhzod5N+cS2Br+BBwUziWFrvDMjnYoWo4lAGsYZIwJ
xAWcw5GbMRiP5a0FI7NZK4PyMSAMEo8daaKKZ8A7Obyd1m8mM7n0I/XFq7WK8RHu
cNfHSviMLrp9TtJtJBmvWtCugS9GeatuKe2h35H1bGw2ljSwK/p7uHoZ83DbTu5t
S4LQ2KfZAtic6kA8Wsx2lFYrX/9dJZpeqBFXPmlfx8Bxtqb60nwLq+j5UYZXlqqa
PMVrXJlmJYAF8K+dLC2qJwLm1k8suwh2ocMP1HxIbSbS5Hkj+thlv8SL2q4ikOqv
pae2xiQnHKVcUEoGu48DqxT/GNsQ3xBwZgbUXGDI8/cnum5R6bey9Kh2dwtyZpr7
HkfxxiDS73MeGw9DvqLY+zbKYyMTseI23FGlAhrIv06h0uuKO9Z3xKpln07K3F+P
v9ogf/3h44oVPkTvYiVWo+DqijAfEw+JHkuCt3YYZ6TGMWUFd+4OliRc57v+daFY
pLL0WcI3adOaKe2lyUKPDtG56s680xSyF0IS7bn/CW4VmkfuWA4joMPFA0qKVrJR
P7P5e+Mjq+sBhVwt49JJgXBQaB0wMsBke8WajmqCMQ0I/OjQBGgeHk7lA8wVsRHs
4/jQkKEQlqsk1YlkOYEgek4mcj9ApoCK1vkeuGDm57WyJ7YNYGTKl2XSa4zj8ffc
QsbOODYVigUvCMM9jFGanOzLpnlLrbZL3Ek1F1zb8YgwMnBYPCc9hSS+rp/A59a1
ZhdznbEI1dNmpHUjHFeCxxyMebNb8E++PYEShjbEP5UX6Wbf3nBITYEUa1/auOlt
Ml2/zfVTxcclUs+tz0goDUWZT4p3Z6c/jL1BABE2HFxqhefSeAmoGUrM5D5S2f+h
T2dfeQRZhs47fjFgFx4deWlk1tKrdetjj5pA0xjKwo5bY8XyYGbcfDgH3PZY/JJq
zmn+MeoUlPYJrusnnzlZimS5OajccWMuzkvO/APpsqaMKKDJvMxY+1mqHk2/I6IP
zagWMFo7ZxXaIC15yzQ+t6/9UtCiOkEaBo6iQLCu7mUsqtTYQ8JTIZ3eH1MnhWZe
bDzPdvqGW5VCXzasQ7VCXua9wMYnukvP9sctFd3l8aIS71rcsdHY03i3zApWwpcS
7eJ4A877chZsGtyfYJ94mf6iHYcoxgTlBLwKISVZzbFmg5w+krqIMzdYGhs+k03G
XKf994zwoZ5RFarS535G1JSRpwSQINWjp87cmRbcxEsSpHdh5l/Gj+H9eEf610ZT
+Gh3ylGP7aWXxHV1lDcbn2/QG2nXSzarCJDGrSaQxSJY7Z75yj+HYVD7+TGAfH1Q
z+rdFqVxqJYnkCJT0GYkhu1b0IyPphiY0j8LNNEUIbj8LPJUPhR1a0qiQkrM4yIz
61btW0ncSi9a/3JBt16H4X5xnrbOmGddungKFOe7SSJe16OzlMJEnc9uFvNsRJR3
MGpnsYEemFweelEcgVFhjKP8/2ElaxcMehlfQVcBCJ6xfSfWHBUBRAiDFtRt7WFK
e/qLR2wnT7LgRMFMC8GjBoJlBDN85+UR1qazQpSrNxSf5W9+AIRnteUnrzX23uaE
1JeGF1O6KyXSOE2T2RYtp5ONW0PeIVU/e98QYmbGZI9FikE5W+IyYW38Nq+5vaKr
qra4MOWQmryW8cz9CBvJzhwaGbAMjOGwvC8mFPpeuHoGQTdfYc4IUHoufghCY2iI
pSRK31I2ZMLpYEQTKLVT+SLN+jhrZVEpG2Iej510nupv/ff96+qMd/ZnJ+ikHYeE
AO+jx45TQGdgJ7bKu+ujNiXE0gDyKgaI9iwW9Py52XlMRevFWL6hPUvq1S2Mt3a9
93EV51MgEhdHjFqlQc2CnamycoAwCW3F6RGSfyJyeGXw4MDeL0Y+MuzzP/+aDw4n
h1RXgZAWfgLTtLLqSQ+LNFnSQeEv1f78/JnGQod2huBKDGcjEXtAFZiASTiE9u9o
h6C9Mfdxp+glkUKHnWxebn0T7urGkAymk1e6ERiQ0UyNQOtMd54TYqcOp/939Va7
UUjBY4jjRSeZDXF4Dxt+33KCK04K5sXp4vD3krqNLUD1P+32zfcUXyUGo0z6mYTN
eySdUNc0WXV6mytJNBSXNJZ+J20A6De7FmIyWhN0dJ75GnsHMxkEQClvis0Izx+2
CT5bRuxnF6LwF/t7j58blfexqwk210yDd0cOjv2Qx+Pxe/cIl7MmJXE/urUiIB0Y
iPkucJJSsxFcREkSJHBv3bMErP0TaxrE4zuxukmAs1a6B+GTF5cLwKIqsQmYG5MR
lNWT6+BIuNzDG6mvWurELb+PVxP6OaqE2EYlPsFaLTuc2mj8SokIB29znc9Ed/Eq
cDl6Vo9Q6TY6q2OHge9ib6zsHRebf2oDBrn81PgVLeF1ohaT+TBMOk1Jix7evVEe
yaTCPN2qq5vIU0hl/VN4Guvrsf/R9uopTsIB2eWLyUCIfZFJG+XzJ7mmSuvoFbWN
CKz9w0JYrXmlQzYRVwz45mE/QkliAiLQivOkIrXb2h9fT3zMMow+RW7MTH9SfXZK
alRYQGJ9xk3XIisKzXPZeRg+JmHUqIckwLhBr1EYJK7H2rd5baz7NoVhKxAy7bih
VJyNnu4j53q3pWe7mocRIDEL5rRMQ5CiRGdKFTh+cA35BEZLsr0dimKEW2/MbQMR
0B4qyN/oUa+buztVxcJAxd+3oN9egkIGMiW06rPslxo/qTgfPtf8+auPf99zMyRD
+VZ54VUCRUJ0pyqYQfuAQfQ7GDHHF1fpttzzPCBCLemfb6WBqqxO7suh2xKNtnEN
PCkhQ6/h3jGRp7TPuFDDJK0LPu0ylcurgKDDzwkywwxNjozGJrZpsP2VwdArjZyB
n9QEgJTtyhg5td1SF4FBtT6m7Xr8wFJ+IdhGazuvQvTx7xKYSJog9IXaLmrC+8Ab
SPs9VZMLu9FDLFoPrQnbt0apQjKjLLRMxOPKlDtofYpUrQGHLf7F8UXLLJ8JXQS7
jyFJA3HtQV9bIqeX+iq+QuB3wfHqGBzFgrt+wnRlLROE89AymoBsO+FhOj5ebJSR
kBb5/y6Ck66kla8JUkhbSNt3hKJR+ZIWpC3qlHV4XTQ+mHy45CDyjuFYUN7G/9GB
t7Ki6YikEOHunddqQ5/VZkw2QbAa4KhPkiySwEPhc0w4SW6XWBzE6FYQV/D95N8g
n7GcBr1/xxD6+haO7Qv0IBljCM1sJK5MBxTSaU5UC9SvmvJl45HRrJNsLRD7nxB9
RLjLjjirFfYInP/g+TFPbron6fyeVTD9X/gGcDY6ZPxgAZAXKI2uCgzCI86xnsBT
pNJEGDWreI8o0njP/oXRCFYxjZxoKHdxPQMIO/RC2j16k1uT5TwmQs/b5QDiDRYB
9K7Gz9tS3htyucxYEEUjHwfQvjhU7FE/RAuv5B6Z342lrQ0NYbWv8qGTaadZxDMD
hj/lbUIqQwKX9oJIslf2yuhgD68HNfRDzDWKBBpE4Oww1huIKhlYCl+SyP/0sX3t
npLq410GlzTsUlbSmcl9aO0TOrY7JUEhvVHarL+HvHg9WR33TS/HTpSdMwluHxsi
B9Hpal0E2ijSDm3UZuoyCDnlzDkuHYNh+APOkknT3kOElqgzhGEE8Vd3PhaQNX+W
4fV5MGcQkRrQn1NUaecdx4KPruclfwprh2kleyE9QedzIgK3r30k4QWKe3KC2kcI
NjTRkJiB0l5jmzu5TGpAG00a38ywpkjfYX0hXCbTSLmJ0N8yMq4sW4CgtFeVkjgf
Lrk2Bsf47I0zyoAj9WPYm2Ue88zJoOI92/SDrAv2yDzMFObeIRE3FcgktdtJbWhg
udlxF13vBXgZEJqw4qixxPq1JmXgeeZO/SPNflmna9KJnZt/TcuJ/KR1AHGJCKvT
udGuXnQiwXbSjTZRiumbV67SbjD/oVoiHFNPfvXQdvq3YpbiAJWn3hVn5MQ106Q2
HDqWOd4cYBs6dXk70PzkYxG/1yJ+CXUaHKaqffIVh20D7F6hXf9bTQBQpW0eyscl
ewlluR1i/wuxkHr2TktsbvnFCSU+MVzVnYPgPj5IX98SaaQIrDWN2Riasiejv7Ud
39fGcGdcHscek6dW5yGfML0wELU5pAUF96txUV+0MZ6OeXyjLw+61d4ZJ2Fn094u
HT7Oz3Gm1cwOwFROeljPZKtGJzaUeI6GHL54qhKSKWSjxIpc/RTPNMAtkdFaly5d
6xmQQHMCl/eacAYnlBPGi75p5WD4ncSRt1vJXAD/Zj5pOxfpJtTMLIGiBxpl4dl8
+rzTFiJoQlzG+Zqj9V7uAN/RdbyChQEQYoYKXtH95Cf+7B4W6rtghlvtW+brgDR1
V8tUO9A4AT5W5EveUn9uxKpJBTM9HrzdNo5HW4G1bVnBhjVAvsahT3F+HS9oUO8U
nvy8z4ci3c2o+Jxr0dZuPKm8yre0PyNBeTQs6YrgnEMuOQFQrCWpKnZLzV1/mLOq
wUhydfIe0effHqTHjVlivgNj7ypz1EXBc8HgWQLjZTizqYkAlvxj0eDE9Q+4oGcr
aDO1+SHdi86uXkfQBPh65wjwXyyMJrsREPkTdP80LNotVIDuiuk/C+idN5igk/yq
4SSevfozJcEoKy8NTm8232tMvN1BHcYvGG2nlxejq3NCuPMtCUWS3/sEvwqDBAFu
xzn1ECTWNpYKRneZsyogRq9a3s6oGCg/aZc+OyIyKd6MQ43jiihXuWX7+eo91sgo
rFUs5XO6893wRHSDEpPscu8RLlGu5EKLtNlb82386z5OToXMeBejqaA1PGMHYV4c
a+M+SzJSOFFf1sS8BgYRkic0RAsLtqIMSrf89KwyX9KgIZk8VJ/yj1mNKkJnUquA
KDvv0ZAjORfTp/28A9YylwsYBCiBnmwl8JcwNOe5FZQjxrpVkyXOXdUoDpM3Fjzz
qx022pECj5s1DHirk8PChcNfpfFr2oHahG/260eRA9RgliYrey9lUYHL5XOkRPs8
jbtdKsNSNbS/XpzIv5yhFFiTNmp9eB8NcRdUfMb5pH9MHX/h17GSA63FEIeXb0Z9
RGc8k3q36yJJZn3bUyvgqLiYV2eNdJ1WYhlfm6prJf2+AZaUdvGi+YHDEb+S6WGZ
5qYDGMwVX6g9Pv+iTneSR71LcHnliiOn9mMT/x9AuVbPEOe20grgvXee+kQ8r0Va
jBCPxkoTlrTu5Sa4gtjt3e0f3/b+D3yK4UcCrytQADZFF6pAt+hdBzW79qFz4ikv
EMTd8WGVtyVHBtKCg2fQB5svWTLhncr+9dbwwwH1nEOUkbrt6ZxuR3DhbCJ+ELPI
UGSJYd8K3z5znzjE0KTgveA1lgGco95VJ1zReOfxPDnVaUQxpEMeqAx0lee0DOOW
MsI2p0CHJlegSSf+NCjSqBFbs4lc/fIy5RBiDxAUN660q3WwOvOjQIKq6KBzxXVL
ceUdwdn7lYYneySXchBg196tuZjxDDjoowHuTP+2EjEmYBJXNRV/JQOqVnnaXu1l
dlg23OUusQg2MrDiINPCXGhivHha2Whu23t1M7qDtpGAjEk3gTIeuVRkZCMmy4yJ
RhAuWGpxK6WPUv6Sgr1m8/n8wlOi09ei6JHc+616gB4DplwUcewMDW+nBX8H5deC
mRBTNZoHHlSmJEV4oiKnpZa+SD7Yzi1oO9TwvmQ7Ztq0U/UbLkYKbO70i35kS9tp
uV52ShIQBW73PhvxjxTrG6AtdbCD2BPDcA/qTH//UCliR5MtgEYujoDc21skrVh7
Z5EwhCVtfi8DxVpnRzRE69zDJcN8A6BcrjT9+GPDFIAdC+fOF6RqnyiHF1P2h1cF
zSYZlyC4J+QREAE5LMWf7R/5rMxcWVQg2+jIXO1n7FSHKRw6hlUgXQ+CYXT0RhHY
D6IgKoGjug1XdFGxUxqlfDFGgm8pe9Vt5aSBw3Uw/uGp6ryj5g5ip9WIQcorK5PB
43YTHzyFJmZaJ6wya95R3UbBDF0NoHbFZYlcYgv9KAS00fPbFzAvliCW31AtDdRJ
D7t5a2SSr87JiAbwYtsbJm/6X4pWuh+hBOyTcEpWL52Rfu3wKMDszFeNKMCY2nuP
QEWT6LWYiW0po8WbSLNTxcEtk1qa2q9j1TTwyXVBdHP4OCLcWxAyttCDwj+kp8O9
Ov96emhHbNQJi27cF22CKj/xE9uDLuFpW64A5FlzBo7+nWHDAtNS9iYfjU43Grib
LYi+WFYDeqA7cHCwFcv3ya1jklTsRnVyuxCfAQWfz0BcJd1oGzeLEUxLes+V4grq
ry/7JFhrsnYbSKF1f1VeBwoxa6sR8pPKIC8lsnUoik4bhEfdYFIbKmZhgbugAMNT
q8P0GOIINwkXNOTJkkkvom4JTAKsqNUP00yVU5FHDKYIdqmUGU3FSeuMBWzHjnow
+yfGkbAHhrLDhYLZYSJxghqGsYyqGnAF3glnk9ilV6FAaehEtPJjtGPx+YvNcPRU
QT2sQ4OQsre1AQwe7aCS30qBXhgXC25dyTapz+K7qnauX/DimD0vzw0068yBGFS6
Yb/GpyQcn5cs3BWrAhmyMAPEYNxg1PgvzRNOoDhCPbWGzowodw33XyijOz/WLloV
SH8MsW9/4usbJuooCkgiNYEutxIf7BC9ZBBMlVnXjb1KVrlLcsbNOEZHAfV2LHkB
H9Mlc5QC0dlvQc2tjdz8JRD/v7gPTv7ZlHhrd9prqEjfkAClRlNUBZAFGuqa8Fkg
gyk2v7kbdbAxrZ9LmlVUibRn5JBhVEq6v+w0oFjs0ynRqaRKMTVImVQtNrJ7LVKW
MENy0Oil/DUEa98HotjOY+9gScdZyCSxh8k+8gN4T+XCkoMwADNiCx+lYp9eafyw
+uLAp1m0ZZ3xWd+5NG6lJv4xkujTgmkldZx3DrU7zqJTw85R6n+o5FntqUEHgcJp
fpZEKumXrdNnpb83A9PmuccvnoRVChfL3wbxXJf3HrPpZ38d4u1rHyGnWfzZMdds
+OAVT/yCh2aPhVgIxC9YxG4CEm244HxpFYrQn5wooBG1fTeIgg/UmhEXAZmtni7m
JHTb7UpXp1zTIg9otbOJ4DKdzra9IPGRARQV+pdn5U7Zgl+myd+csHS6BKJ5hHWD
TXuGI1T3YXm6cRt3A0Nk7e0nZK5swL1/w8bmpOKri6Lsn4BVmDXcK50aAOCNd78w
ZPW+5AaRRbAP0VL1L8P/jtJkgVn8XTcORu1peSI4uahzxlNlKtyNgfgahe+8fsWt
tmZ3prSddXLfR4LrJ2omwlUg0nBYSueOItB9zH+akf10+JfO6RrSInjJvSJjw+98
A1oHno5PnYETwqZpEpnB9OQaGbcFehggFJHHJrcU4cIErPmf/YK12D2GjmE+N/WT
hrvPtwPQtVmti9827ZI5nOKFdHPTlgLM5GlFWwBKD3NikcoGQiwMVUWrFIXBwsst
AnZZ/7otqzJ/EOX44RLfBw==
`protect END_PROTECTED
