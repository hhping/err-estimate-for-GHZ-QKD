`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1dnJy23KRCQkstOjJygTs3HffBO67b7tHm9Wa1cywlC5lk5v4PelCT9L+50maxLz
KuDh7zAlASP9hikRQIKSrgZoZtNhOSfePRDALdnkn2UlsJkPK2oWVyRWT5qboAUX
DxQLUL0gRofCiWM1qJATWmbPpcSPyKD4LosU6DJN0s5iF+QBWfH2B+oI07QuRJ3i
J6CQZR39t9BTXiu4NDQ6VrzwipsvGsxC4ztcOXU8kGfERb0ntkeI6zgxvLYlxxhR
Rl+1ykLh5K1+oPa2YJ39SwdtfOaAI+QY/pO7A8uelDhGQgXeMR475/0bCMavBz98
I0yobyqzqR9Ek/q19Ejobuf757HmPjlrPHziv7qBhYiuMdFNDFjIsuC5+Dl+Wkpu
hMzWHufIpumVYNSm+2rq9P22npw1FJKHYL2agK/92ajasYofmJ3yJf1Bi55LnBGC
QUrh9nNMDJOXVTA3dzUNt7ddeXpyEO09tmERJb5IeE1m6Gnhek1C0s/M465Ap7DN
1d0JcWopve+Mxo4qtems6636vN22NeMNzkLMjh8k7tFISJN7angwtVISbParnAZS
WWnlSDasZn0GS9MpjuU/U98xD8ZyP/V+djdtdmT19GvvbdHL1l8wu70MXNE7B5oi
ZdJNoboSFghiMlqxkT77SlQ2dMBUUBn3CYAOGGOgwcEfbjn5r4HcCid9ScTWgT43
YAv5yIXgZZ5LDoeOMfoYmwNTa8IH9N97HGNnOPEo1nFu85cCaW3dD3hUPr9tJ1ch
ecPXVFmHJH3Q/pFBbTy3UFrWy5aBFm4FcnB4qRG47QhKePJsaB1B4eMSZhXV/NnV
7b3ACQIewiX6DbdTLLIWBURmbbedNloANegZNHxzVEhvaT8eKChXMoR9+9eH+sHI
07nJ+kkEgNnQvGCfim05sqQeNtscOTFUxb+ck2HevxqQvdQcmmPPKJkAWh6q/gXj
D+BY/F5ONJJysl0mrRJ8L4F+4kMCVIUmVEMUOdwjy51jcK4zS7QbEkoHBurMHq7U
P0qYXDEat8GjkYal3m+pgVGM4Jayao7mNv1Mh8Q58su0ohMh/RkxM9iNAtSOjb9z
EIH4yaCQs+CHmaRnxo21eKoZe63mBXjHoQS7FNWwnGiB4TAOmF8Bl+fz1q2SWeW3
dcIDvsCUxmPiXD2DsouiREO29HPi6JQqQ4sewoeExEnP1xHoiBlq8M1fL4T0Ficn
d1mKvAxT79kQLk6MXcPrPrtlGVmndentGgXJQrJs9tTQrfhwCgibyQRffPx4ZmU3
CFS3F5C/D1w7puOt6TspF2weLi8DTW07o6NDRH73Zrfa3BLzd/7m6eRjFDlVow1d
GhoOrGetGhC9C5dk5O6d4vzYGq2veUWzOr7Ds0bguLVOUUS2UMsyeavqFOrYYLWQ
gj2u9T37Q+Y6y9PajeM0fnyH6dTvOVY4ImCVp6cqYPx4r+lguznlB2AC2YQn4akK
992CR2wKEyQW8xJnIhZeL8TqvDL32H78mLR+rkYGeq0OvQR1kxkCWPoYd3Wm6JKy
iwV9XR+PynGJ8/zex9qJDM9zDuOBFmHc9f+azfZvHEilwFUIE8UBwhR7iUc/bCXy
pdsTkKbe1Iv+F56ceiv7bssJ+qZg3nEdLvhlzshTWMAUMSwE+VwNADlQOC30YjYR
aFX0pagF9uWipEvarOhoGiv//SLP8J4VX6IG+JXehU0RhRWLJYpPOSrT2G8Z3yTE
UzyJwmWX3XzuaZcUOoGupUwm+9N0VFiyfsPQBcPqT27Jsf5bm3CPyQL7qhxlrisM
v7XZo/6CyacjF/q/FFla+Gvg36MYyqZpyXJua9kA5BI1G9gqDTsWe4VRLpzR12Fs
sqTFKfEg7BMjBVmEz4yPy1P/fWBPDY3fIwImog+tFEJL0ZmuxTudxn9N0pFJ0Nwt
uWtZhyYCr/Cnhu8uAUa3za4Axyu4zBFKUDkDV0ceUwvBlj2mHjqt2sGkQEvTAu+T
FDb5McAGt+eqWy/hc14FXe/PWzh1UNfUCA1zlkSs5E1a1D2CxnOQa1KZUAjP80Ws
ONPmVl4secw7WrXA+jFLeBL4GQgudHc2A86vxDlE9tfnds/5MbIMSlnM3ELu9xcS
+ySUvUY4oeXsVJZZ1/PioWm0LCepmZWeTz0+OqWWmJStg6XP0M8Bj2DYDjVCGMTq
wSXgAeN3zkCzRO5759bQVLGtK6+lrpTRQjmMprMZ/6172SS2Mfiwntb3q4UzBXY+
NVh5HwGgLwvhl62WQhQ1ri5h/nYwTrBxcEJaht/m/TZY5HB5tCgQbNPvxEwcqPSJ
ERAUP5gE+Z49d+lC2bdVE6DvDjK+Lea8whCpfj+W9u/Tqibtv8/hRg5UIt8tTshT
F72iEJuughNMmuVveazEixivEHpsLsDsv5YOgm+8q8LFGbkWdIZdQBehXjtj5XPg
+KfT64F7F4yggN+5USSRAOLCEVBSyIBBZ53fNUK52ArGxr3G+rxcovf01k9MG/I9
2Mh+FvDywVdUtCiEdKayGws7jPfvlXtrFRXTAU9QH+nXsZIngS/gmby+P64yq5kZ
khlUAbueXy4DOkPBO9RUuJtRBxH6bFMcWzhtwdZ3Pi4fI5f926N+jO7QVJzDv/nb
IxEwjmHvM9veVeOdJWBlImsSbpZtBKsAyr8tes7RwOQUAkC/2qBWGDtVm7VTffRs
DviBUBBZHTWMHElx4IaUxlg3Ly8AuJBbOILnQOo9sjIuxSPVSJNE8hhFHfutbrGP
l9EySE01AIWO2TBAkiNmjT89mIVm0BhA2VmYLLqX5oC6WrQAB5n9IoM5zI9kcSSm
mzNk2tMgR88J1Rk2rxjbCYQsBlIC+NQVVGgDPgn0BnfOvK/QUN93+52M5AVymqVP
2ZSc9pnkcD22yMY30mKm2Sb4ZAbqcNnUzFtk+2r8HGbzO0xaTtjunK+69pS3YyAR
ItmayIu6Z6vQX6PF21qqg9NcZfuFegC+7Vkg8kn1/TlxS32eyORYsuBUyKUPOAWo
KUzx6rSjlqe1NCxFs+J6yM83ly4f0jj0zXXdltTFEcSxIcOmvl0zyVkkHcamnxTi
9/+VQjYeD9cnokYFjJbGU6JBidYUkSBpuov3nkp4Vw3uerd9jRpVE97IbhknKOO9
1ngvS+DrT1WSuOkyllf37jlLLouAOdkwCK/GQuYR4XGtJzhwDZS58zBwkg8rZIWg
OIYYRY1U5xhCZFqmK75TpDk8q30wQrvuEqEkIjPxaLMhwbPs8v+hRDVWv5StLi5V
IaF8gREYa8h6ChbMh4wbYM6R8oWut72QyYDKGLQm0X9HumOfqIA0wMtLslAoOvTj
Zp77xtTY8TbzV5ilsmW2AW8vV60gkNOobtnf+o7t2EeMo69LEBX4hEv5BqynM93O
VUNDp3L1TpX6CoiedEUjyNEnono+uG0/uERxkRxn7e1fdKJEGmXZ3XGQCEFNW9FJ
2doLPCG5ivIoxgnWonegs72LtwV+qZR73Czp45ZA7BC1nu7LvDQiDsYIj/xt2K80
cTIfV2QwAgPX1PsSbdC5U616eTiRwpx9c6jWSvcMc2F5cLK+p4ueHeYW6dVdu552
XaGGJlVmhAVTXCfOEh4aYfL5tjhPlxuT5cECE6wPOObfTHBTA6KJjl3pvkrXtiLK
LuoeRM/UpzXEv1JjhEZPkVT3YJCgfxLzvxY4dvXBsgpyUO6RLZoZZU0WYvr2AGwN
28/+PBZhw8+2w5yEs8VucQzwwK/x1rxhh3tZfArRSYa63QHRPzKqLylM6VEVKjoH
m2K+fF6LT1JHwKvXqnMZlhz4y28T2nyEOOCi6pewM4Nk6MmVCMZP7jQN2n4UBBv1
bSBP4Y7w5sCRsF7iktYUzULn1zgGj76BU5yVj0Abu7BlfHdpW/t4iBBn+/EFjmyx
979wP1cgoBXiE28VakOA9BRal7RGpVUYLqXEMMBjrHJeoGTXfE/kTqk3z9JZubWD
fHwW+90zDrfilebi4ffk8wpheDFxaKKqQtZYvkGNMv3ohTyYcA76yuQ6OXDEO7Tv
Yq250xxWZTt7sRMrt3Dh/R8RYLXvx5WbRY72LXgesB6ve85ldRliL0CsfPLg20iM
7USo6YiRKjkYGG07IZmLV0t06cY0+039HCvPIys1RA9aPILplmDYPGbzNs7M5IvQ
BghkrU5i+8v+1jz9m9H+BaqM2RMwgpb2GWuED5WxNGLljeXl1o41GQ2s1kfmDRpS
lSOXzD8twJYFrU3GUABXhjJMyVXkJCNUScP13kWeFjPgnT2DIBAFNEW3BwNdVhvj
HzT3P5V1RawvY3G2UmOhX7EoAAtCGG3wnn9Z9DE437E+lSs5IbaWo8eLzBqXm//w
JBkEEyU+1dCwyDox4VZ1odGpFLEwWkRv/xfUQ4hGBpnMvaoUtecwQpMCBWX+TnVu
WAvlNFZnta6Dmn0g2mrrgk2AuEua/fmTJprbOK7GzQ9EQqwNE8B29a64+UWmlXj8
B2MHhWG1QuB/t5zuwmvXUvFQ2stKSB3lsO6nZPLbc3tvsfr3kf5mtd8zFl7i8HGo
Y+tTdBlEfAuXHCkcA9zxff7/NMe9UCzKu1HWpgmk0ej3ajWfexp9/mKh7IcengdZ
uaKCEkGH8wcOs4cJ8ICdERkhi4iou96zZLMB6iGLVWbZ77tSXIOcr1O7u6CZswsN
KIIPDTBFCqRz5fU/rzaOXrb2Rscja2wZEHR9A36FCp+AvnPgmG1oCvbaI4zciAn2
b2O9v1mfzXmfxYGIZDua2Yji0Kc/Hf9bFK1BpDwSResZpYMZZwVuaNSxEvLQNphe
zbItBHSQmF+qGdvszSPxd1Eiz94sX4BI0gCxA0gLW8T8Om63yvZVeLBJr4NshCEy
Yt75YzdkY6hYY4mZ1F5IuQXegAxXhg9hD0WYvsKZi48JViUQUeSuWJyrbLLiwtKk
f+Sf84jbmFQsnhfPddn5JxkeK+1lCjuFsYfzLzIqgcUIRWAS7JMuD4+QGr7lqjqg
PaIe7XE52Giqbvc8rIoSbjl7btvzsdABoX81rh34kuMNmlk31urYmhJmd8r1YLCb
Nvlo2OtCS/4j+4aK3m0njnl9HwoqoeRDGCb1RvCWPQ0VpOkX1+2xTWYMq4RKY+Ms
6EX07es+jKPT9eIQDWq/2Il2GeaoGXEFTvyAd58N/Z9PjZkUYncZEwW9N51V7C1a
EsSLxTMWfmIZyMJcImAwPwFJTsVdyWjm3kGyL0KmhwvFPm1mw4d61Wtj1ZCP/3Y0
ZHrAVl4dIvWll74DeU96JgtiBWgOysGQ28LRHxN9AxIJpuVvbhvjURVL+JgUhQLU
TEzZQTug2AfxT0RshAfwo4Fmy3qZ8s83N7P5FFzBDWmqHw7Udi9Up2Ko9ltUWhRn
lVkllm+spLrnsZ1KWvqIitulN0s+slrbEbc1h4RPoiSwSWIO5glO/4rlNkzv72FB
zwEc8RMPCV88RPmHwl6J0733BoHBtkV+WdDAws6FpH/s2Nj4aUJ77fHVcVRv/rBI
4Rz0t3DNs1dV/bV+H1c3envY6IU/XaGpwqhG+HdRR5nryAMY0F6Q+b1s2b1+5jqQ
CIUqouA5OoK+ph7F6NDLx++01lKuGUkS8M3AfsIrigTX3L0zMGNEmWvN24TOnJqG
Vz8KN0SK14hs9+BG5U11zzmAYA5/sxfOLZRRwERNT7tRbH2E6PC3hhIyZBODX0a3
jpm/62ndSmZAU4zEmkKY+7DvfBFmeX/eJY9VJdwfcri8uGEXF0gbxqew9cneJYJ7
iOB+36PS3iyzAnPMYrQuFDKPfuR6hYidt43xUPUlj9jqG7UWB5HAOkYs49ktyURK
/mqDgdYN7K0xx6Mr2Mgsh6DuBg3vmEGZTTgHEM38CFxOc164uddBrcI12BhFuZB9
WFVpDQ3zWzbLSxh0ep2/lHCbE2oYkLBy1ykP8rstOOnEcZ7qBYKPN02K1xE3L/6P
Hp0cUePLJJAi1xHj5/i/PKoI932DbESBSPzX4Njj8PO33I7w75oPzRvvo8T8VErF
Vg1jEbU8Eddy5a81j44biDa9B6qppgbmZkmVMgvqDwqfuRZ5cmd4UnbN09DjAIMG
qAuNNDgsoZKHcZokffRpVYmQwdWsP1e1DoV859o8cZ+0+xcbA+wJ7W0oAnNmK3qB
jD3zzryVDdZlJ/LXkcMQZz9UnqKhDL9ZLRaAM/f5povgKg906rsBty7VsMqbvBFe
j6UFaoTXJK3R9GJux/DeEPwJ78+XZY9iUtRPsgfZP2QkiM9NWv/BvXN6W4qFUX4k
FIwrigZpcqbSH4gygaCsBV12YlG1LmI8hPb1XBKR2FVYkhPmMFtpDsS3Qk79kx6S
IDQTti0gtAIocKsnlR0ZEWB6GUn7fa1R6FAlePL+UJrsnhij8FMdae6myfRX/3BH
4IBwM0ClDXFE6tYMzZ4wMX7OQ/trrTA8cob2eorlm0EeSD/pGiK/EeEUtOhOK895
t0v4U79Zwjx0jmOIyzb27LAkBGNdsUQu83B9vBR4toOaFOaQO/sUMYbU+PWApfOl
wQKa1MVYHXjXDegQFwwXyTixnRXRBU1DoSfUrJ6wPPQnH7n/hcKc3+CqpYTtSTV3
I7Jqb1TZihh8570K6MYCUBXN+maEHOjhZjYZXyzYQVZSgvIbuTBlYVQ03jIKaESO
ydkkDQjhvwtSqlecAwOr1J6u37mc/hQ0/H2W1hIe9/KTXkDH+PtknDzHs31MG4kP
ZHmP0OaWiRSjXOirczR19/aJFGJwGL5+hpRPVLIt9iYIj4zThUv4MPKW8kbPnsNR
hyGnYPVTWW4ip2RJ//8ZFMw5+3bzHGKms2pw0lUQ3sT4GKHMNEH3pu1GMRX66wOq
MLTil+F0ZSrnyglxZQa9TuiwBlPcaf2y9CXsz8v/W3XeRB43LomCSi/A8XndwgNR
WBQZYPrtoaC9CO3QB1/heM6fZTPRjbPOQB9HGF454RaQV4hXYF/MiU+RvVGP0iuD
gRo2/40YjMp05yHzoWAWDeZE88iguJ1lHgfNfFe2udoerIir+G+UzwT12xLMfeL7
HoiUalr5If0cul/MpTilLwOtRgJC5gPXLi174TvtkoHh3UzWAgHTgUl/r8W7rFMN
8j2IkxovPmgO+neh9prAMiQB+5lxumIfd2M+o4bODazkK7wHpFKZfU2ItJy4/O9e
ReN3nU+svYzxWy9LUnAGUDjO42OFQBwfs0IqjveXpAuLpwmZWWeKKJ3JU8tKWHNM
NVPxntRTb7xLlmbD0clVKTxPgBQx1vZ/PXxl3O913SlVcUHnFPWIhMRS3nUELHo6
p/yex7nB8gmyeGDwSzTEnIvwyaDoIwpxNG+P32KuBUC74ydzyTYQOb45lnv8ioEN
rS41u3ye9d4oS/7jssiqyv+mrMGMyW/tbD5GgH2Ei4IPn4xjnhGl+aWMcUlI5JK1
h9gfBjlfHPjihJwHY+LATLlTjMOYTnHMZZInrp9Uj4jXcQ5sM1PpuQvw9aY62l52
wBllPKYFoQ2c+tYj9Q1s/pgmTnhLKFlVUXmdOKZ7oOLVB9rWvleuDoMqW+WDrp9C
mGmA4HlPGRaaP7Wtwi6rHMuZSlPTjBlmgzMcx/1u4YgWtCvSiuUa3TBaeU3sgjy2
ZgJA82soq8gbyg0672h+JGZDWOUrXcyQjLW9ZYOH0okwOnURM/bcGswg9TvkWJ7D
EeNip7f1d1jogQqeb8lvB/rSWt2bsAKgZDShtjMhLg75Kku3JAg22/wAgRSTCqih
CoJsItSyPXtX6TPyEi2ZYbbwWl2LF9CxyxLBPANdUEWFBqTde0QEef6ekgbdHni1
fD/kUenoe4eXIvmWOS22RPacMr56pQGyDWSkIhUAx1BjzxZPqPbkmQFW/b39fgBB
6fLa+oA0RB9xasg4j6LyQQMWLQ4w/WekSRjAWTGllxQe103n/fJ2RtHzlTEX+d8p
2DinQu0pOw9cddTcBtEAQVDloBP0hLynAEcdLj3HMvZ++RccgmoTkPynvFjHUAB4
b0xPp/D9tof+HXn8nchvH4IA5XP1bF8Npvj1ndZVnxDHwvlBpCaSbQwrWUTa3TCT
vSBQLGzziJ67z1YF5R9a5sSA2u0w553yG8xt8egkHsjPVvEOsOaQWvhu5GIqZunw
lS3GZWS1Au6wTUXj1gwXZCBxo1ZnRueBRm4h+qXBaYg7C3/aK/B7ybog1xRT5ZQ+
8jtVYATCx5CNKpYOgJ99x6WRH8VL0IxtyhBkXMhaew8egxiKjEen5cjMLfpzQxxm
bQeguqjOzw5qaxagkX+pBeMqXteTuz90mxpxjuWnzcmwOzqY7UPuQoFqHIPPlD5J
Km7A3B43Iq65jXxGG+zt9zb2ETpRHyRkJJdr8N3vmZX+poUcLYcemMvNRCFf6yGC
sspdPnWmsW0dRp4O0E6KM03NWzb3/UA6qQ/tpsMJtwoY3ep2aA2NyK5z+WU2skcj
JjqOfT3I03jmfq2CPNiuqWbuhttr5igSFeVp0wAaT24AK9K/0O83JxoKnwTzf5ml
fG8mVpGMx5XeVy+mzt8xCpx3MNpD2jykcJyxVvPBKoAfLzr5UDidIw9JZBeeTHUd
yQIJBG+b5P/WRAyKatNDMeh9gM8E3Ca45AqCON36XxxJSP+6JYWPSQLrj7nK4HfW
QHeFGhR4ftzwDK2oHoY6SocKlrvDJBGXKnjpeOtG7bI=
`protect END_PROTECTED
