`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fPiGZ/V9WLHe0UgM9+ucbIbPI0DEXWeUVWgt6gqTkg6e09sjYs8if5FqIOZthpz4
PfvZ3DYq1vubwtGu1iGQt2D9awjPOkAHxduNs/xsNJyvY7pOJ1hWRviSaPgpV0Hv
iGrCgGMG1pKAESNEjZvFTicmx1IGBZCnBr+VZ7lR/44OjIC82Mgun9jjOItOcWAl
eeAS4xlt2VziaeFTDATxn4uVni+YMS0v+CxGGwT71HWFiiwY3h4n4zwY/oH8JTi0
gp1WKED0GQ4Cd7Xi2uETwrIBASZT8lFQlIhNK2pqCmQ9HxKoB28iRuEoW+8gacVD
eDvsDCkMH2aC4syf1P8FrtsQbwZrCp21VCPOqM67wHGpIW7sO2t9H5lXrTJN/xuw
QQoSt1200Vl6jy6xSJbEB/AjjpHE9batJjtTm2/kAt2MM2k2eIyJezr6PoKMoaYr
1G1ySGHXHlYyOYmUvW2hAjalGSEWZ+aASNKGFmLkuaUKgUjit9tLjkkrPOu9V3ry
dEEMWmwWaiq7MQHPZyAGq0fH2eAMW8Qw7obgup+091uvTBTLOQk5Wo/BlYJJc3hh
OqZf9nuWt9F5/Be8nvXYvQ==
`protect END_PROTECTED
