`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0x2g52LGMs8HY1Y36wurqmidHcv708z//IP+qU5dA7D7DhfgV6CroZFlNE/3xENe
WYZraFlg05Q0ORRJQEabIam627xmEaWvQUTKWNFTl4MXa9PkymTYYAQCmuxv9K9D
eXx6nNUOv+Zurbr6f1loDXS0+mF7yfuH+2w6YSgTgokbomwQRGGnU06BP9L1N97y
ubSkXfereiW7b2xnybW+OiIfZ3tpiuBLKScnZY6dM3IF7vSWNr/sg4P+gKYVmQg+
Jlqj2NDfH8QbUYbpmE/f9vlAnchmIci3Qed0KEhkFabRefx2zb4jS7VVPyhwXlZ3
QZvUV7w6FCrqBgR1tEGroITXhjMEx5fDZ227Cw7/cljNlEquy6UM3Snu9e9aFkyp
7sfCZNtml8sBzZC1l0QSLtDwghFTQuJDip4oLZ5YYGoR1dYCb6lhNXJiFhLr9CGI
TfzQvvTQoiA0OOcXin0XPYqufqY8aaBJqKy4yZMXb0g7laA1Lk1UyuklvhTcpEpQ
MRV1LaUAGwLcqz8A557qHEMmF0GnH+G3P2zGXtG6qJOrH8BcbyqHsuSkg1Qms93M
cq7+XmyxtynSSzra90/hiTQ3/jMRie+i9nmaPFZZP06W53IUnjklTa0n6I9fizcj
V8xWaUNmmKnPwxu6JciPy22a8CgQMyKa0l+bsb/PABg3Yp2v1TmmcCSc1LmrHsPh
sO1fn2TSlpdz/4lxjO9/QhunXqRGYZdNe/nPypNVOqsnaxH4keURaiKoELi65SnQ
/gvPwxSHpMpavs+4CJ2gT5eT/R7NslaV3MLhWOE0b2LPLuyfvZBSddXUQYP4vumh
DqPVy1nVNG3B7b06HUP0lz0qqi8aPBcxwN1/QlZKXFpBPm7ajP3CoOAgSBFikdC1
amKceRrq7lYDnGV7LRUw1dnztvL9QtDI6ST6VnH+fWr0DYmX20sKXaL2IkmPkHw7
zrnCo7hc+HGXE2IoyqBuWJpLSSOxUtCzjCBciOl1ntjNF0ccMkkdrASdaB0wnp4w
52g+/tLd1NpkpOD/xOxOtH9OYDUzLswL3VhOa1czsCpuJDWEAI9m9CL5sFXQJ+JM
5fTY5JLdWh5SfjV01KuyzK5hQ/tPac4HeYxmNmP9uYLFm/QGPIJ7p6JfSrM3g9Ne
opyTP+Ot2YVnGot62wwrFvzJSSV1P9gCs0z78iJVZcN/V6y2T0KmoAWkFH3BKYuS
rEe+HHOs8rlzwyxghFXjuQy9pg8jz+CnE0dULydP0Emz/kZA8r1Aq+ZZWtnKFYTh
D0zfdI4extWDiOvCFfZ673LfeJUB3HSXIA5yVWe6uKOJjdp6AgdteO9UtzZyQQFt
ZVkMNKRug8bjKxM+ECzpxg==
`protect END_PROTECTED
