`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
swEQGlsNASUaExEcJo5aSZXoONzxaKNqBgcYwZDBNiWpvJLbll9Xi9d7HNQhe8JO
SfKat4oLEIMfD9EdJsfOv7wX9NiUXFp0G18n2HnFsH0vzUqAGAiS+rJ2P2JnLtxD
Hm8vaIjdrB20w+0XBFpc1tM4B5lDtBwhOBRjds6P4xrkNf37lNNwcyhpu8uwGJ9Y
bhucFmK0uKNyAzMxq2yYWWpQWZPon1PnigvSNBkuKEAru6ExT3BKRDeIZ4PHkp2H
qK/rAJu9BAAwVyUiv0LTd3Q4bBPsenlxZzdPDCHP/LfbYwHDRjy+LoVXMaB8A8Lg
6f5Ky8hEST3uSPI71v1M1YpYFHgaf6kWmdtP01xiSnvsHRxZVQh748HaAIQr3kKS
72A3+e1E5B294CExazD5tNbKcEHbrwg1QNjZw2C0wACV1nkw28Q9ELtaL4mRJ0Io
kOrR4AYmI6lB0AZZAP2C0hh+O8wRsR/JCrOycojoxWMpsfk69YnVAkJceMDby5eI
pXxbSljLTk1Je5XNEW8k6q38k19sFZBRtXA7iwXLjxDLTikmiFDmgBewfGJXIb4e
CLF5RzGsrJvZndkuwH3bmUK0v6NkJqMrGjP/JTddOWsDCtbWqoGizyjFKaLjap3f
XCsBkmIOMHUemAntHhD9l6YoVKLtz1A3UHtGQyQ78NoTrWFWu96k6nWTWGLdkFaM
c19ZlybXVZ9iKfQcTx0sAkg/PTH9//d8eVyAAjAJLrYDpcodXFxgrm/M3lFBbEYI
zHgxoc7a/47qKwGIRupjQhZHZlmur0Rqk0LMy+FyrzS4wgOx+33ZfbzvvVZcxCdn
aKcFf3dSYmRGqK8dUtRzuBBAVbZYaXkoyuc/fB3xksZbqaykjGbeQ8qFtBOl3NCO
G7xlOiFU8CWdE3xFP/KzmU0IL0NcCoFzJ94ZU+hC16moA4wNMVadSch6D+ybYz5A
WLw2NJZvrE+X6uqv/pity5BJ2raR5i35F1b6f69Xs0P3WovgAOoxG4LEpQK2GV05
zsncYI4sEW5d3LrIUelqVFH3nhub03F61VB1Na73pOr2l01WciRO2VjFqWXCd7yO
utdLbA/lFBjtUDWQLuuJ3QXAD3HlICwWT2jHk2rqlYbJRDRavFJvZQRslt7Xzywy
A7N8Sl0qUgZdTr4HHrSu3h2nqcoedz0NayF8fzYwoqpSFZBUc/ohql6ID17Zjo3N
M8tCaPhH1Ig0AVwSrg3/5MyynyaZ9fswweBcaIWQcheyIZyn5Ut2Lfg3/8VWad/4
u8yQQ9kMXnJugDOklSaV5bCkKSZYqzaXnbt+Ge5sOv89D+oNo4vN70PCvV2XdwUI
nEACcCUv2GZvWn/t1IPO0nr+4luWItstbDR+UJPu3MawUrJFNUhKAX6Pj3BmW4AU
MSv3HFkUbseRUURDE7Y9jkY5aDgzw2naU/E43Gb9KWHyW7kpSYLEYPTaODkcRrNq
vdvjoCOiN1NCEAhOd5o9MD8S0HugYr1cCkYHqzY42+g=
`protect END_PROTECTED
