`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v+a2x5G53L3lRKyKyKsHi5zNVJvdCFV0mM5kVaBcL6eOivwtNedp1XT70wgzmM/h
JA7GB9VZZj5KlqXyRK/a7TgpWahZ81N4DQ12ZzojE+s7Ygd60QwOMo4tcUEoTflS
gOAcJQd6/90qbxd2aubAiZ0LDwXW6AFX1OFyC+MWh+vAHWkYgwZ1rH1gCjIVTONM
urH54UL0ZvH40F82uJjEczLteIVZsYe2oGsqDCix5c+rb7yiRK51l8s7ED3ldZLj
ZhqxWkvGFvdzqOz8/fpUGA7f3WRc7NYCuyRkQf3vrLCephqKFnLoPjyI+yLKQkFl
hBU3Ndljxafbv54XUTh+DnjFsavTgYX0/0PTuCCQV4uSlOBEKjOXzewxFWQ+8D67
ft2NSJ3LdVev20wzP/J0saOzMA/tO6W/IK6lwEPvqHFHiuFCjwAiEVnOwd/l6Yjh
S7bILTYSTND/Pj9kuVEdq1jzft4M25RfEpbjXbOEFpB4ECl6eoG/L7JFaZBLqv9P
`protect END_PROTECTED
