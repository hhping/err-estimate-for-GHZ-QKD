`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hAjn82tv1g2kJNRwsvi7U6xdy/bl69iEr90flxC3rc6aBspwkK1ssRREelBi8p2S
CEnN8lFnrCDrfYtVgX/4L9vQA7zmB0zMKTj3LdGkUQvBJzDENGxSLPhEtrTxA361
bcUq4B5xJ5OMytnXYeDan9/e/syw0aABHwZomCHu7jv20LgJ6h0GPxoETSSMawjo
rKMSM7knAjS6C6AgG+osqFZS95V6154tUUR6P5ewbV3UW2AE4edYaMKC9ENq0eCX
4vwmiSc71wnmP8qU+8kV3BGuAam9XP8kxOo6izEEBNYmvGQFKi2sPPYBTB7GV2uS
ypx6ntxH5+7knTRPPThHdmWC1DK2vxHamlX+kTS1iNoz4SDDJzXSHGu3fa4OqGe6
lHA+RjdmtGkvUv00zMoQRMooTwtrsqMW01+2S7DtGjv2qx70S/QmyLFqebcUpWbX
qZUj+g8gF1vO3BPRP1W/ymHSJ5r6sZpwhDzmnDkTMt/pSoYB8uiizs6WvWxa2+FM
7yrctgY7I9hBdnbT9UXRTBpMoQ/Uo4jxvVCg6darN/U/+hm7nez2FO53nMPAQ0CW
+jwNXNZ2ceqVwar4gKxFhcjgGOEsnZzOrpC+9j9NP/+I5APrbv1OJUO+BfRvswoP
3yrz92rNMb2qNnYim4G9XtulT+h7SUfWHtmlzgfr5Ff9HodVin2UeZa7ccwEYSsw
wOEBXxctEUiCYtD5HRU/SlJTACzMAeGl1pXwOBG4GomevoTO7ztUj3tbBmlrsseR
fXoJbjd+FBHpOXn1FbJkdv1aEZdnOjur9ntgtnGnKPG1AGIp8pXroAmTaL5H3WUx
6cNixTltD76VEF1pLgYsP2nRFPRgCmjAS/UxMypQRQRXVEGM2lMHWJ5RGraxPvtx
5m1j2t9fKAhYK9kpEfrHaG1+cR5TcQKmAo+JL3DaB1iW2dgOF+XsRNa1dz421dA7
vPGApmgLzVhvMA8BIvqUdNERPFQJOGFFY5tF0Qs3FItrlGKIAP/Bdp+TYY3rjQ9i
BAgHuDJ4OwITybaKQG8Y1IH9V7vhqex3tUblf8DZXKb5ayZt2JF9ouDnClFzvkbI
kjU/g3aMfNDAKc/WqL+2FO0kfe7PMgm1B7xclmAcMiX5lYHJpcC24QRYpRIrvjFK
ixVgTCw6RH+6EgQuFlolCAu9NvJ2L2wdedAoeuxh70SYrka06MSxLw7Q9UBw+GM5
I/W21B4iz5mLoSbTv8MhXfvPtuGmcoujxQxvXxzPeQKgZdw0/2WZSI5utFl6XlzO
kqkN0LCXzDNMRFaucQnZVUI3NqPHwkCAWKBsJcpH9y0wyqewTBB/kYIUTK5PiDM9
udOL/4o7HYQWgbOyBYHT+nMeBk2d3Udy9j//vbRQ8POBskqaeRp8+Li+Q2ysKhYh
haKXX50wggjXZXhmAUdh9YPCciA+M0cqiuHCjIbisNc7PnVeKkIQhlBU9+pVJOZ9
g0ESuKAsPArjdh2Y02NoP7nmHiFM466sHd1irIar7Sw8JKnK4gArkd5xckBbl2v3
P+ItC94s9LYgDV03VIkvhU0XiNleFfyTlQ9OPWN6KE8Y4T4PPYrEm4g7TBximFw9
NBmKGBDRSbJGZxXBmemWruCkihDlnP6GdKxvQZpaECssTlXnL6akq4DhKfsUYT85
ZS+bo8o5AocbJSAB350hOuwiRH5XzZouBUMlwxphpTKbIxm78cdj80TmRpLCXGw0
9wH8wJ9P3tQlUHXbx4eCT/ICuupV/IDgsQf5DdpoXKGpAXzWVavUwVMUqJhRhnA5
kS2oRM4XOP/aKWB4tqMw80g6vfEqa9H/OnKo4XyyNDHY9vL4Pc4CxRL2vuIodVMq
V1AF1/9RJ4dezR6WtUzW4KHnkCDekIOgZBmwdxq9sfwqx9n2wVnTTeL/tsmuc6DP
AjUbvmOHDx5b9hawJ+BRUG6ZjY0UScHXhv0j3/H4M3zC2tMeT0Lq0KDPqdm5Y/NL
WvjkEv4mKw2tKpv3Bt+G1uAw8gW2Rz5EpFSiWFzo1sxMHOTx/WwsibVfLxXzRk9U
0djnHVsq2/5bsWGW2Dzdw41upaRoVro+AIYlzI5Fn/EMcVFO+QHozOcBDhia9Dpc
k1w3nZS3Vme3pgTT6HNFnD486tNSObt1nK3WNRwnNKR17TpR2NQZlDLCJDIDiH3R
dfLVltNU4tNEiibOyUJY10wgwalGvvcTHRjW1XoIIW0T94y3AjHtmQEkAk2e2Q9+
0u+cShjYuzgUDn1az/0q7EDby6rF/bzBk2vpu0YiYBaqa6YIaZ2zhKzakgQA+P6o
QnBKu05PSDRIh1/jFF8CsvB9rGUaxSTVdYhB4plwlygYuhzIMy7AQ+ZAnFlxeLzq
aJgybxnQWDVFhy6gdqjFD0mrJpopR8vbLIuXsyXx+po8JIm0XP4i7nxPnJgBIc/C
KUxuZ6BVYFeggx9AqUznYAlfTdtZgOWfDaH8B3B5LrPQbnl2JjjyqCHq6XnRPjOp
34Ly1WsQUCM/AZesa3nGdToSFomnxtT0vta4eyyhIBwuGeZDEHYBMxX/eJBh34xs
zh3DeZ6ZsjXfjnzyosYFPmq1qTZIsqQGPjSEdQ/XhvGWoTPE/T0L2O0lyAn7o8x+
aC6CeZXfbR+jZOpOOvrWBrtpiLv/EfZBP/qfg4AG057H5Z9GwUTEQstqCddo0fh4
StF8R1t+IDDxOmZ323qozHkjEfO23/gQRFpbzK7nISJbuvFk2CZ41egIccL9p2WH
1z6X5kkBHhUFRBX98TQE02K+d61yg74geonTqVIK9Xz/szCIotJFwkZDipRbHseO
7+8+6GOTlyH+bwo8GvXHHx+XkXaBxmM2rprfI1Oq/tUOlU6kitObhpTJYjIKMWdT
6tTvgOz9lJqrzhtzS7snyevrbuD6qffUdhnDzr8cn6Yk88WADQCX6x90l+1v0fN6
F1hxnaQPysQjYDpCr4nXueF6ecvtTmA78wzlroT53OI=
`protect END_PROTECTED
