`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o/Y8/3ZIoCrxGU5Su2hh28xz0bDSX9PGDnAaX3FgHVC3DsomzuMWBTzsOa3Y5ADg
xCl3wdwEfLdjn5jmp99LXV4GzfTaDL3u9Gzu6IXwnT5j4/ZdfYy2gZ7AhwFkzmGa
bWI1Z6gcKdJ3P5wi9eF6+4HaCNvEiBPEhp4970ROlymFt+efKMfJXs0pD1ZLUG2y
S2Cz6iR11Rv+Rs++gFYMHlFHlQe+nrLC0I1KXhkoroNTnxAB4jfgjDY7HUUomCyh
drdUOwSYyRavj1B6JxWifxW/B7hXe232yNm+jurTco7aplkV9TUHeYopvUlC1eoa
RI1QefIrtaKvgDl0vpftRbmxnlMLsa6/5MpAh4b4F4UjyeULd56EG760PVKJwUmy
+EzO18UOWKobWU1QW1AU2dHIAUI4tKjgFRO6AMjUftTwnAkk7DExKkElIBQtPsYS
oxqzPqq7A7WKefWQOTEpCVQ9Uz/1CQNFYMSBzCZjExh8aVynaSCktmBIZ22oLAlr
pA14I1g7ixveXFQqoz7iQ8wpGYXeyWXqOLGe/arJXyPWkheTxs9incrKf/t3xBHR
cqJP/GfhOdFDtj1pHSyYW7vwtx994sFdZ+khkvlvBnKuG57KcLRzo8xXdak8CyyP
YpU29XblVwxJ4IYtv9vPK5YpryaA2fp5q80K3uhS1cGsYnBqL1n5KxoRLDTee+GU
+TS9/xzrHR2DI/jIGQHhWM6xIsgcS/sZ6MtUXV07FcMX5+iWXgL03uVeiJJ5UioG
dSB0nqVwqtRro5z6WLLfLvJoX1+oeW8hicexcCSfRoeUESoVYbLjuF7IadlgVOlx
A0+85Wm/BYAY64CaEBIb/kw3jf6U8y+NRlttPe+MVkkABHyJMvNpA0Crd6wwmMVG
fPJX5dTJo+HYfr0HCyMNSCP8DuBwaCKds0Rxxmd5EAxNnd16Xz14eRHxe00OEKS4
BIIY1zGZsFTyQdzGKZTSWLlZTb3+ZrAnAhkPRa3rnclHV500ZeIqAmD5v61wcoZQ
oVpEE/PaacDhXzYm+0njX9pBt8De+KRg2kw226VoPDy9b+CaS9MdXBs9gPkT24kv
B71Fo3rTODEOp1AQ3iCyYQwdo4/HyW2Ym7edZbaIBqetpjPi8LAusCShcawqda5I
P5jMYgSDTzVMqv5IdKGBEgUBow71Pp0O5kVwjYekc56+XRXcEomqj0+48LdvE/l4
a8VSY6L44VZ215lHMXwKRCDEo+Su3MhVlwW/kxG0wWp7o+93pABxNEhcOz1aZ/YH
YV3fkh5/2wpp5gqroZ7q9to0Xkd5Xz0Yxl0YvVTfCgFSrBQAvjBa+WgpVPEd3nSJ
aCn5KdV5h4YjTRbljc5WZArY9UD37AMePxANkOhDOjZpG1yTtpmslGKpJtqTUvVS
9BWDR2pv1gTtFL2zvgRl2e26Idd1QyHSDPUpCcDvIjJwsnlZUHdRpNe8MA5TUMqI
fSixsGM2K7KOMLdZBcD1oIeFrkpLUa1ERknvmmH4lWc7F0sSyXrcH01F7/cVj4aP
DfVPf0z0aq/x0ih44D+LhtLlyymuOHK+hqjrJ2avsb8aUf1jry303Mg12NEr8eEL
K5fABmLYYTVTv8xwvkRD/YzIxZljAgasSJLX3TuiLmq/l3Fb7u3h+TNlKWtWgl2S
wqXLzJ9xUHpYLCN4pCOp8d3df3FvU/16t3nXr4A/YvLpzuo+Nl1SE0h4QDb9Rlrr
n71J8M6Jc9+pVq+wWG2tg+Y8QhcXStRH78uBqdnkloRtAQzJdfHcO/m1UgNE2Xng
J9zO+6tCxBRaMlxA8aO4Tkyznw/7FwTnSFCVsCzusmruAJgn8n/g6t+UC1HeZ9SF
6hmJI6klBUAVjJN/ZEhEGxNHLZAe/8LwHm863KI5u2UpXSDMHFkCbugsuw7z5Dfm
bRK2gTnJkrJtVl/SIKFNvOCMnCxzJc9Vr3VR7s/uJF4oEI/XmWIEISdHjGHSHZpP
F2xyV1t9gUvfFmGEfDr+dI5+HERRysvN/9X4YbN86EApmLTir/ImCN6kiDsOCzjn
exwmaAUDmk5mdYODz4llDdipWJN3MrevVcZr1H1G48har2mjEksIWpDnx7ZQhMMN
/lsF/DEEDp1M+SwHj0LxW61E8uD+pwsZBEA20ynmq80UyppSv7CvPt0mZc9anrzY
7zl9orSHapCfPqul42BOZmbb03cDpyOXf5DTfPgnBSB+kzKRq85hLa2hhienOjp5
orPlK+O4oYEoPqCq3Sm83WAD9PbJlFEmR8QDWhaaEGYaQqi+hH1JYwNqLcF0c2XG
gAmpvRrJbGDDqkWNJHYdx/O2uhNqdFpOHH/qzrXmNRXK4jrMrsa3oG6TJaKYPov+
symDEOf/86yPFcRRa8hVv7l5UVB27aIwyf5PTROpoqIVPGx2jZD7TyQqHiKDQWGM
d+n341Vs/db1X0ZwSgkWpVJfTGAmV0ErfJS99PgIegitMOQc95g2MQeBcGERx3Ek
7VI59CdA2pZw2ubOp+diH8fa0tBDfQWdxKwmUxCMTxXsfVZezh31XiUg7/ysAqHs
2jQ4QMDRHYBpih08VRlrYtIcCv8YMQBmWZLvdK02sRxw4FLove86jJ1/ksm5+4as
03HaWaBqvSlgjoUa/8cfuTiu2JW3aMzzfQZPcWaYT0N4YT3nqasnOOlkwXqpbm2z
fAD1QNAhPQczL2Xtd8jX2ShfSI5P9rNg0usNtghXrlMKV8szFVK8B5zXOGiCpPPh
TNLgJez891pbP1BxT/tO+SomjeUbBzko/LL9Tsu0te7PAUwyczSD92og4zn3zurR
m7SwaKd3gZgzriA6jD//h5R8GvyX84vyMzn1FPAwkrv3Bjt/T6brk2tlL5tiNRMW
VPFcRDylFyMZ8dNErHxxlSdS+mfVAa4tSNxDNCAXfXYdbIkfH4dY7bQPElwCBeHA
NmIREjBX0/lG2u6GW1qbjNn1tLvxC61MOBnw4MEo+qjTlSzWbjmO/uYjqvKzB1rz
FruoJg9AdkEeeByMTcQxFFDbMumRS6XRYUs4WSbUSvBnAgBiUF20ObGWEolPi8fy
61MK6lix6wAfNuzd1pjg9X2J0F+Ojqcb3YAnregro0vE1ztIjWMmXMxLYe2aAi+J
vutW4aPlt+3Ml/2RS5jzQe3NTkuPD6W/6WQfge+v6ehI+4FAp8kJLGMt0j7wWYnd
N1JTN8p2dUiLn4R4J7shlOGXcCZlhNnlMRP+MinR6N44bkKDzZl/5jZeAjqUG2JC
y5VIXS97/1TRWfJkj+NTV9KhqM6JlqlRtBc6NNv1ZFTbVDqYkf39cGeOtVfM8O8/
2o1iHt9kDDFqAkdFdznwrcUOHnHc3gAywXPmFHQ8IFR0p+4TCCjA5PtA1EMaa/k9
WF/bJQdQc43+J+O6De2IbkeEjF6S554lgJajC7WSJCPw+5rm+N6z+7glDNh2FvXm
1B8g1P/OelhHPssawCAQNTdqXgGp/l96WWEEgGsXP5JbCgrcNO13XAhdLu1UXu1l
U/puR8dUWd7x/zsoLaKma7nm9mnLfCRNwLDGiIk9cyKkDlv3IKqoojNdzTs4EkBm
TLp4kpYRoB2xSEU0UpY9hNU46bTRLcFV6sjF/lxw/zPirdh9SPUxN5RBvOq6HsGM
8r7QLHQ52V61d8e8kvp+5mvcSOT5nq0SduxmaY+vIwcawmLaLwW4Bsc9YDafgR/M
eKcjlq5w08aS55sD57R4YVkhCuSByGfNeBS8OyO25AanpJBAnrNpIIMLgmE4DEeU
wpSZoP/sfINVK1ZUGh7uLnHCIXZ4k6cC2/BvMCVjnnNw0r62d9HVlBKRvgFojwVo
aZYbGNlPM6ovR6kazs/Z9cIKnkVPq4ie4GUwIoWwNMToS4cmHml+NBjS0k5y3vi/
8W9pBiGj3M/WMHoh6DO55uko7VPoK0C80KnEpnA4CXWkjQ9n7F26/k7h7n0hV2ye
fG5lqowyCTsv67E4dho+LGqxedi4F7Ioc5mLxwn/npbSfLjzdrOvF+sycpygZmwq
qDqvnszlS5SJEX7Eu0Bu9qWxospIc4gTCsqz3tr9lbNArrCsKLzNEAZ+h6rnuK91
ol/eEDFCzbn0A5Ty3A+a1mZYt1FQt+xY13MMOHzRdQPC8po8iiRJh8yjlpHGuK1I
wrqZE9vfi66LXZ1YC5e58LctHHXq6+FMjnp5HcT7jxzZVXkI+k9gtDSTagfubk69
3zv5A/RpO+WD/2Alq096hJOsMDjrxECgf4svLYzk67QuHBl8Azz3yzOaKs0V8EgO
rMbDw337DC8NvuMqgxb4WwYDf7+RjMLA55CAAvqdjTnO/XHayFK/oUhIJttVzyVs
m+FMmQMT7VrhaX/UVIw1ohwpnIklNyXtlLOG11UBlxAKOyZIEiymU/IJHZi32/fv
bgxGrijGa1qJVphWBq1rOe4GEYhq1zj/06N2xNgu4IQpFSvB8/Jovrv0smKILlBr
5UMbXAFPzsVaBESC62OwsQb3y8B7NKP09H20pXPxkVHPfZTBBOGmRRIwiied3+Ye
0S9ujOglbcQnkFIUn4xmYRh1Gin6l68p79y7ilme+0crEKDhmXAivS9jfLH4G9yO
p5WJWoKTVLbDuGwKFxCXY93s74YrisPubP7KJbsKNxo7af3p3ORs/2M8J1OhZlSy
gkDumhZpZHp4AmU3sns579jUS7m5+4h2ySnLMKwMlIubpWM+jqpwC+yc8ruKOXxF
gUnRI4//04zaoH0yuUj8VUIhj+BPqhZ/B7/O/EfxsKNvhb7u2e7hlEyoLjOoM45j
WR3k/uwA6KKFuPINb5x/VqQHLeyA6crjf8zKcF8cV7WLgURpQfxborBGe6VrmCpi
LR2IgZTIVw0sH88STnauD8b8UsJMNdjeME4ZJmPBzLeedW2wEpn9pZBHXEu7a63T
hVjTCisBQxbHUZdvu6Fkhrmo3lFAUW8FeZlDzy7NX/pa4qrJJrkkd2vb2GmXJDVh
+QwDPd/kiVtSTM1rih8KxD5TwqJMaeiNrtF99B+TRcmoXctOFyriEqGbEtwpuExg
8y9rI82Lf3RZvGKrZZ6XNogHECGnoCkZeaF5pD+oYXH2PCXsQC65PsLlVidD81Vh
QqwuRjcuBcNtr6vqtjlwIqvIbHyiauGzXjxWj+xC1bRq929qU0Jh6YM6XvT/HdqD
3d9oHcJMAP36ezN2bTmEtl9Xj44bjRRV9LgK/xMvsQYJbN6zJo3zDskLr6/bDOwQ
gWVvjGKbGsPAqqBYbTb2nuNQ8DR23r+I00oBhEXsIX4=
`protect END_PROTECTED
