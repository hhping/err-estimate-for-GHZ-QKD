`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
urqEUiteKtDT2AReiZCu3l3axL8cr0mI9QAzneWg29lI6U97cBRV2jJLJfqQc1sn
f6PovSMouVQIcBxZgh9DEs99ID8UK3rNURln0ZSbwXrbpSmkN9TrQu7DAR2gS2/e
lMWIYqHhuD0wV+SYKJmQkTn1mLGZkX5CnI2NxRYXoCvN+CVb4zBulX+G0IRkkk/d
OGbM/HqOVZFyZHEJVzGtLcom9gRbYOulPN9dDcRh42o5x9tbAAqUSnAywYOLqWO3
zwa216FTk0f9ZIdKJmU3KpBCfmJ5NyjZUzy4KG6MmZMyUyMKomzU8zMzC7x+2iKJ
dv0PMXqroIX6QGK9GJr/3ij5dncq868S/2EAlWyxFTU7zl2hw1+qd8a1MpbrBI/u
cqlYPX1cZgxhoEGnDyekqKdRaf8Qg/TJe7IjevEOJL62lwBgw/z0Qmv+grbBl9dB
vuntVMeq1Raxy+iBVMGfwRKadxCbwC6qkhtwgbFvpsvm2nEHrVvtGr+3bmhS0XVx
nhaeNRpgdoQ91JSQCybGHKsCc2vtW/uDbFIz3vAh7jiGUazeASAglkhefnl39ngk
L9rR/y4G2rwY/FePyiiqJJ5mANkPx8tNFnSRc+VxUiX6gMFO86oWY4nlbXFrvkOA
DIwY4l2HxEj8vGgpLVl56rOlzmdeXNLCwZjxYtNnFeJArA3hX1UYQN+kS9mFDo4f
54O9688TlYBYWXZCwf4owv710TUaGm1zXSO7nWTQW5bHGV26uvxEXX5PyQvY8uLs
HSwmtirF38S42T3i71LyPAcigibUL49m5Lt7i/RFfujA0nNKIdg64Hf4eV7Zv+Ah
PjUTltePN7ndYV3FtvwVYGMyTbVCqVYjVC7MxvivCqFoCTKU0m1RL4c6SZKUXeIu
6H5AHFlWT1VGxnkU/+FeVYDTiMPtQw74DPm00glBUQwRPX0Bx1EK3twiFYaO+haI
7qch6AjsCgiZV5DWV/TEMw9OEgZJULFRlEYKxJmy2HcDqi2o/87pIURl/m+AxA1K
urRSv8MX30fcmXUWX2BZWvJ3Iwcq9Y/8TS3+0iOJP+g0FY8VdgFgoNy5tbaworMl
Sz3A+AZZLoWaOn440FOUYVGZIsCfRC6bDKgC4dUoVX5NK5+r0ikMSsicJZT2Bzyf
1z/0EXxJyIDloMIUYSx6PqOmwUfktJ+Vfj6+6bNcU+9MjqPdSRvT77VCeMd5ChKK
wtqyhomOC+UFHDPcHUt6+0h85zsxiqSjCxRSys3yW2C4KSx5FwiKbwTgHwTCatfD
pcpRwVTdJaulFhKzCZCGpnEPpm8WuF9FnKLnJwkKB1HalIao+BUugW1WcLWXuYFn
TBUQXu8ynwkwEroAb9UYTg==
`protect END_PROTECTED
