`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9HNgXYudxwYOd8HKZdd9yJjyn0krUMdktv0QS6uHsMzVkEeCFVjFB2dCNybg5xEf
JcMUa9Z9tXJAnP+qrU0z4klXBbrI64bXE88/7Wvak7TIAjzsFjKgua6kCZt6AZX/
qQZHDGLOQTVSiNuzERxm5seg+33uDkNV7JwPHkySm0m5V9JJNYGWS+bzg+cNJP0e
PaOzCm3qhwRSE9O7SNFCpfAdNbwr7qhRiwTPJe7QuXq3QaoyBQkcJqEXKbfIelo5
Sb4whf0nZtrYHNFjHjgKmMFuxhVccGvmG53wFSCiOqcmtJnYmngvKzoB9LjzjC5x
XUp5tX4V6FLl/hjs+QHDbgKynEM5UTA9ZXIjGk4D8+Fw+xx2O1v3bqTYwabA080X
pipVMMmTsCsLsE2CEb6jND0hHOnC3hHeTRhE56pN0FvIHlYNfg+iFcevzNawAzz0
ScEjgg16IYxUHQTUy9uRLJhGZxh3Ryz7D9phMqM2DyzLWllJL63NxhZU75iDD1Pv
XQeI/dinurbBAu4kyTiLju0dIZ2F6CgnjgvmrS6Yrq4kHhEyPvkKGWYLr0NypIWx
cOBEaivfo2uuWj17TOGDE4QNrlFEuPQUI8ThEVDpy0XhqrG6VOi6hFmYJXAL6oa3
jXFSPVii3f87VsxHGSMqy+TP6pjOGGGuqA9wFb7LdW6KZgkaZrKECur/Ysm0SfFc
VtSYhbNMwdMKbPmeMmeUuHghi5ryZXL9J5goc1t8oPzMhWYDgCLnBxX1+DG+xhRe
RnSg6kevSuul9H/i7iEE/fLyUVPdh6GDn43yvaxhq7oGxgBG8domXEigpSI49rBI
h3UqBrHUy1Fo6MNVL8YqI/D1NE0jFRC9nwgbWdWAqUxH5+tc6xc3YgewTtzXHZC7
43frfuDQJEzDFA52zx4Y43jICmBo72xAJviXvNW76mc+LxFH0M9AWhfCXxw/Vrm1
u8nWlAmIp0ds1bHUEXkI3REeQYlCLQYDQoJgm4amNXxo/he51riCuwjWNwQBI52d
/4nax2MQoIog9NqQ5e868Wkta74RfIJaVY4RVnr1kj0V3+RVvu0uYYZlx/v02o2V
psFNFnjx3cCT+gRHFmrmVxZLfLshTo7SRg7x13xgcSnqsM2AmgOmxkyVMLT+6ipH
cLE0ZO5vMZ874KwkiTF4uc5xjBJkXesZESFS5wvkLAP1vxBMtUDhtZaR4Ri46kMD
S8Sq+/q2dbwAxzKcDpuMW3TGpwcZcmgui31f6g6ueW1RTBL1nYpszDmVwNCiv3PC
Vp8GNcBqoflfo4GzDRt+6iNkFKh6cx/oWC6aXO7dLg+HgOt+69Wjpzos+cF48TEw
6hL7E9Tbf5uxhZfNBUR5SvoZuD40ltmTSH0+HdrNjXXQ+1Hj4NMKTRl7wzHNhq1H
ywrQMmkOA6CbLkGI/eugOUrOy04pimZ6P1F22htf2G5RQXKgE6QyW+qRvBZ8hbF1
kf8b74phSUP7YmOhLbMfk0FFe00nyZPM3feOMH86IuZw4VmhL9xdizMQiUfTRTWm
T/F5glF4RQ1XNR7E192wj8Og7kJRWrQEX/jwp6V9OvrODH6HVYgSXVBdTl+qscTE
YP8aj0OAYLXbb1pAajyJH1Z2PnNd3xgyAhbevDB7LpGpdxSyXTHL6jn0z+1H9w+6
7rtfhhWBOTTv/8yd0JWk0H/ISpDOWQIUD+9K6Jqcgul6GLlUSqrhxMv196gfjex9
WShV7JadXtH94GlxVN94b69Ogf1QICzRsipUPoUqqDL8hDpJPNmf+LznNKJY4L3L
Ji1i4n+OQCd//8n/v/2wt9GoyE+XY9pxgq/lN86gW45zr6I6DMdAF1iEWiJXH9Vm
qfadg23gVhvwRM46UzWjJqlBvqI68SvYw/uG3ypYKV9yDyCFVi7LZhc2+Wfx2Atr
NINzj5EO12poZo7yAI5FsWgyaTPb3BhJsemyLnTqpIWTAwdOitOfKbUuUTJM1I9t
bF/hHPcld5QOyh9gG64t7R6MOXgH93AOVWSv7tsbSiSfCd/UeOx2s6Vx1wyvkFnF
+8Bku69xMvMcPbUyO2y2JdZ1FgaQMzt1guRIElVeDCGMkrbfwQttHl6stxOjXvDE
NZI8O0wG7r1wXgKso4Kmv4e6YA4K9C3Wrf5PS6BfdNkl3yC8sXxjRb/dY2P6S+Hz
M3ZoVb6L14LhcI8DSehX+KAzO0FBWf3mH29R3zWAi9tF/g8HsyWbp4R8nYDbxtZu
4vrE+4UYr8+4CpcFMvMEEWmw6PcRVPyJuiDBiGkmNfDhzb3LX+Asfd0EZYcXotqb
TgI81FHHM8765uDU5SqroFWYCbb/3HKrWiMpMSO2u/8wfsn8mGEJBVoOpOsTEoXp
lTAQ28evBTDt9U3nPpJVwI1zCCcFPBOpvDAhTxGUj37blAxKT8M4uqIg6KHfoq+8
6CMNIHX5gPPK0Cmly3qtbN8WO6faAGchw48LiMpzKLxiYHX0fmQYO/Ce7ld8y2Lc
zacBGSqmlSRPkFldxFfGZ1Lm255wkGRsPBo3/f7qO8osLEZcYIjxYOvJsbVB9H4E
7MsRuaOijGe7PJO4I6urB5tnIXrI6basBhCBc9KcrfUYOVBP7PwEBWOVMM/p8I6J
zdG3ZTsy7pv49dzUK+Bm/H5lrzcPG9LggHeShFv9diRn/9VP332OeTtbbvuHHWwN
cDkUJ1ld271BXHGZ4yDcC0yKptGI+OtX0UJE2RlUdC7+AySAAs+fjZwopWVZTIn5
teaBP3eer2AdPUdk81m33MxsQLYehuRie6IDE75mYTIYppaSK9smayEkjBkRiAbz
QRFNlrHHxjdS9ppJsuehvNJxMGK1dUF4ceEsvi4v3b8al5WMbe3477fLtxvtiKdY
6XUDKe8UAL5udWl2IOLmwEsI1T2LJ/mYkIYOWBpassrawfc2R/NFE6myQgZd6cha
KTGVYRDyeQCGCFxY4WSo5iZGmItiUrl6m+Me416UGNBxkewTFjYHVHQo4yiU3AGC
sd9j9AHOFhUMKpZKSTVSojpUucqIw/h4t+2JBjOXmx0vJj8ChmIuKub0cq/cQDI0
vja+ciFR9M27qMk+ee/PQoFKQgfbOHFCizaceXw0AZvILoRt1FxiPgDH0bNHYqvc
wqA1VDwOcF0X4R3bBidrz93lc5lmFUkksjbAbMRqdne+jrH6Sq1b8LQ5leE7fBeO
aK3Y1jvhrXNF9dgvQG2tdUgptyyRajUUgr5XckHg/4ugdvRdai+zq8ILGMgg5JfS
hGKonWoWUTHJP/keqW8cC3yKmSCOoSUGR+W34lok/5eIpoJwB3PlmCdz3Fk+fuUO
XouSBMZe99booh0CQHO0zdo0F2eaM8VaiOFiAEfL3GnNZdm49g26Lj6tBKhbCtmc
1CgfHluEWYHeVvx8fDj1vj1T1/v6FZPsJCflLPlWfUIIqFJ6WpKE0g+UY7BEh+Yn
O1w0Xy+xlBSYnaNsVM3u1je+7cBYjjEiOtbtaUSVlu3eOkRpLfdnW+CPoCYl44Q/
lKfPnmhKgdvIIaG1J20l/HhzzyYo6RhEJtKEhwLVXtwXL9+ZyHc4r702C3McibX8
5EqfXNYFy+MACKX836fLl1D6vqmLhy6p/GxMvWuagtvmACwe8Iw1QpZvRH+MgvK4
C3PcIX1p2wfA1UvEICOoDN7WaRhFvLRbj5EZ8ikZSj0gk+VEqEVsaFrYtIRWQ/dn
yTwYJan35LSOCS8xVysUafUZytBOpdYN70SilXfwN93gdB/FA+6Hbmm1A2l51HCR
KHhQUVuPB5IeWJMfHpWzKUhMbu5DS+/KZr0wPtViN9wWLrrV72FH4v+hOBlsDC9F
kXcGPKwKKGOxaTGSJzNsGIdMtAqoW8AqpAUm/q20Y2NGCrDGGbxZ8vD0HVVV3D9A
4rvM0e4vHgfObXf6zjHsoJSN1lcKrABzbBd/329RT8MjOUqIxdyWueV2l03qiBuH
VWfhUG003oGsmNY9raARpnoK23hACAuvxA989q7/WrVMP5YE1OyMgh4+cUjOskh3
zcnObvTdVI+56QA3b5bKO9OAQ4WRNyY66ArY1T3a06KbSZuZp0fPtLj5rAbjPVdH
wICjjTrrpHeRBL1a+pfLeyAXPjsNvH7jB3MzbPJmelNtZNoyUvoAQ97aRMOkZ5NA
G5zElg6Gl/9vLU0m0f+Z400+P/+fCwSviLLVDfVEGoJWPw+kwkgCMDktaJ6CJvMM
Dyc4pF9RtI17QcZtANilvnztF881s9XSg2kMSc5RRBdgD8Kyt6V/MrgeTd9geDvv
0H3DmTgENYSwAMz3wVnpGjM/YCcFvhAON5jDROXboll204HRi0ACohR0NG1MnoKJ
RPRyAKu6IUQbTqumLZ7Z3qNySP0sb0BnXGRN9bN0KjKANsEsHbr7DjRJnBmZ0ehJ
TuOiCQIDOy1BUCha7e6Wmae36Zkn4G1ocfCOHieDXgHFD+qDrjbKMBK20qt22aDO
l801Hq1fBI2ezElWtghjF1zY1xbnT7SulzdQQcVG1Bhvzv1Yt8rd0JNWKG+MIedL
3h9pRf0IQwtcAr8qAvy7IJlK8iVETpKKiXnXtpiBeM1RdxgtHDrsxqugN7uUk3Ri
qxHyz/q7ietUccu+twZF1vPy5x/Ol0/NI2Itt/AmI9HPRfsJBXCZ4Q/7TszaIhPa
QfhFTpratRmVoMjei4E63LidMW4Hj6gqypyeKmVwAzKhr7JU9YTXRO+BtYJ/4onr
odHj6gNfRw2g7xeaDd+WydqQi2p1CFiUbISnG3ipTAjJqbtYcyty47J1Hf7yuwlz
EXUjRVRE4f0FZB+RycXcasYc1rtHP93mso9xoTq4RY/5/ljUaMtwn7zWM8jBNpTF
iMPAsp0fX0jJle9vgzLI+84jh2HJCEaXr6YPA5nWYWS16jsGgUo88p2dOPqKq/cu
sC+UW8RMQcJ7UowbSGA8H9diw0268MNBg1l1u+TTzqr7AkhthbXk7Vdwg1sdFlZ2
rOoxiSxo3a2Kc7EfPkC07kIuKaBDvZtSx+nS0ar2g8kNvNWJm2hyW4omdIP32uMQ
d0Vb+lyj6RvSg6IO7l/Ny1pnY3Ho1XXAiUof38+8ygj0n1fmtASgJDS46GQO/ASP
kcnfCYD6bQQtnxZFcaqt30go99mDdnahdEgVgpQXkLE12+bDZhzGyM+s7nKSjIaw
v+6mJG3j9d/VB026Y2OPzHWeEx1LawvQOmi7aRPNN822KUWjzA32A/AOR1cgVqrf
g7zcApHrpKo/FybqeVUGua2rfJWnAE+4TmY1UXmllU5FOIAWTDiXid1Oz6g96Rfr
neBc/wejwJF31dj/vdpra9lZlO+LkQi1ni+MIapRK5/JAyM5ywfMQ9ijRflDFIXE
jg4YdHvgB2hnTS0PNbA++T5/xywF7Z7KOhdTxArXPcp8meb1d3obObf2+cW+8+kM
Cbo2Db6dKSzq1ZlUf4zr7oFm5IjhnYLq8fXwHyYMdBcbhU5657xpAQObgd6seSzW
633TcyYc8cEmd0gShqo/1/QlJ4EDGTzUZtp4/VIjrrQpZt1bDvjPUv8IzPT+3Jvv
5VqEyfVqf7sTAIM3z8zmcGStusSZBb91u2Qu/hlvmii2aOebcvX2m7CA916p1sdI
/NNQ2uI8ftfSMSilbKQjRD6y/jrJOb416BRXigp72TDT0Opy6iVpia0oWYypuZmy
0CK0an6lqyZzzl8CD4oXBgzorkxqF6PNbQMOE5FSQkHb214JMcNRyRVkkHx5bgbU
xtFxduT3qgajgowRWTaloivuq2UOhLbRF7EMbtjCxz9ctPA5fQizxeBGiTrLJshi
1Y6hg9D27pCWIYt1oVm+xZ6GKyxmBzDP+/ByuNli/JC3XIuuU3fuO2bAax2b42/R
wKtfuizcV6geP25e+X0pC+E/rbyv9ldYOXV2pURiTBsaG4ESbDg6oh2yK4mRmS9+
rWgsFPtazXtf56OYITLGfldn1QJaBFamWDY5WOPVXdzq7y0+Jgxp36AMEoL7N24S
fPLHKaE86t2tKRPwbscn2Sj04+anBHnaodRVoLsEFyp4oDcUkjFk1BZ4wceaRCIy
BNWNKrKsCHhwpowxTJ2cJgw9dkmbDeONtw4ZCQT+wkQJf090IwpLQGr5ulTHnVG7
fcwJNLktD1dP1cJ1hOr+I/DKaRfU9l2ZrA9bOFfyWVFMOrQmwT+tSqhDKs9+4Ksy
v4wWSAg8hmBIEmcMmnwghTHUp4mclTWd9le1saP0Zw5CeAApHhATuWefR1eRmnCc
/AblMN5r0E7Xhjfpx/m2Vot39SlA+Upz+Bbmyx5Rk1aKTnv+SKKMByAIcYxGRo91
xCdHXZO4CeF/FT+7J7bidD9rsBA80bBjBO3mDPl2mWtg1SnzNcN7te4oDuVAyaCP
ihgALbL6iyVmi2/8fY5f1YZXUYmFlKE/mczvOpLf3DmpIvxtlQnfCzfu2ActpOtA
KHaWi05XtdaLhmupqeOhKrcDFyL6BFqDdmvVp5nqm/rang5bQn9ua/hBto3gecAY
cN2If9HOPha8fUm4UsiwaUld1vyXzR8zrHZmlNKqOi4a7nAqAe8QetRUvj1QQFEI
tyTi3Bj7Bm8ni3G6IrI5s2JwqysSJzSAW2ybsRnuvA9TkTCPCloI8331kyjK7dXN
zeQmq8A4Jc374AOeAiALxWfUz8S8dLanXS8GWKJDbMnbN5N2IRdRNLq2wSft7bAf
PKNKW6z/wsrrob6C7ZPRw6CgJ9QCf//b48nTtjfBhAnRwOW3zaqDCtgAc6kpDXFp
U5hKvxO2djOzMZ3dKYBFwHh9S1j8EtDdbHVSP0VE1g+8mH189qEG6/EDM/HvUtIY
WYLOypKQM8U9CWiJRSeYU98Oni8nzBam8cBCb1FVsopwLnHclycGfqW7YJr2zxkn
MWLgWEuoISOvVAFdQkT3siINMA+gG5Y86r/TOcWzByY9+zBhRZVVwlickqGtO3zW
M3uy7s/k/Efqdz/cMNNxKJhOpMd4DM3uENwhCfxfgTpLdxU6LwAgtXDYN9xYwl5L
wM5CtrQML3LkkW0VNSYRyUYzw05mCGe9vgBEZDFU+QSgqiC+N40PcFyBx2GOfqm4
8EJzwZzZGqw+L490oFsLHDzKBTrHjWl58ErLYgX13G3XjRP0HmzZXiCqAWSCyBSQ
ZS3rb8MDlNZUbuQHbWalDSInchoswVg7svc3RkhzSOu/RAHl3Q+K0ja4Ubd4XrHQ
vO8+U7lMb1A/5DLKBefu53j+lOSR/OfDS8N8RK2DhrpIzvuX2zlv/K86zNzjISGB
SppsG968iXrpprDpRCXXIeWevErzOwXAqVR1FERDBrQ1CCfpjCbFyhTqYdRn6Cuf
h/kkRb1Dq2qIPiKsZUUZJjmc727HPOWEbFpSROO0oRsvQ73BoTikjyoPGZWK1fdx
HUiTjn59hSdexpiNXEhdYVbaSKKDtPeI+ZUoEI2GiqYIH2BetNPUCSfjtBqHaxF+
IUXK7dR+zjDeZrpoip5IG3/+AsbMekdQIg4zdkh9Z9PEh1dBeo3+fmcpOoyFOqO4
nK7z5tcNE3LhaiIpc5ncK4DQCikl0ZF1bLz5004N078WGaydtscWCCkdG93W3a5d
hiizoanzkwNaFIuPnei5EfhpYJYNAIRExcSU7o9n4cBRrY4hqXJ9mP/cIDTRM7Qh
Hk1uhI4IDHHKc/Of94h+vrzxayBRZG9Qhy+kWPI510iHPcv6buub/d1IpCJAdKKU
2JBo9snt6oueftr3SOaqTD0opB2Ub93HpNKLGY1WVX+DNfv9cVeP3yp0ktOqME+4
xGpnyQn8V7EQo9/olGAE/hBS5nA6/NBScv4M0cjxjOJiXbQDSppqf4VCWlltZUws
2r3DGpUh2ddN2MQqI7xs9h2+xccY//yCbPjyHmmtbWeOzl6EgPAk1mDMHkRQuJki
JVkBUNJ923gZH1i5EVIRp4/H+9mT0ph5gyLNNs+BsSBqBBHZp9ZSbXpwYZe5j13m
FaE/mIKuOIAdtCGZIrZeju/puDwHFvB65/W61WTUEPz2/3sfdneDPkklNjlpLr04
SWeEZVVxIIuU8dis+4jz8urgvvQzzLLcp28S0wzoHA4DHBZcyT38VhmgBRAEpvee
TlK9goyugFFUg9haDpyZC8dER/wwrhVOE4O+cE4B71/ohzJ3NxdyJT+TedX9J0kW
Yf/npBuhXva7z6jQ8Q0WomeB5I2rIq83eR8Uz0heAaheuvmbDmCjotZmJOcse78P
oz2x8eUPqsWTDQku4lo5qlO7yMhIbKeqx8ezDm8mQ2ZX0XybLIpeV2mr4p3TdeH8
ltbPeQMRS4YVJU1OpEV4+b7DJbQjwfBeaKH19sdog8slAtxGZF4yDrkxPKeASNZa
/PuQ0Ads2XO2MEUcAG0oqA6D7ksa1gFpqXO66UsjgmxPZlu7cYl6qor2rLRf/vFC
eZ/9d/zyPYR1/AQv0Ob6JgYi4ngjzU6sQ0xe1DPQuFgDY7IzS8SlUioaMXA0fWat
LZNgIu9q6bOAzLdrCQKYs6aqPnFqMHX1uhOE6qQHY5PAVeoE+fYFl3OSEc6gXZDq
nyxZ7iJZBFGtBXJMW187iZg9/O6kjAXZM5VVfbrPG3WNsCX9Vnx8ltn4eKHhO2ym
i6+/gJBtyNmDq/eJc1mRUAElY3Wy/VEWH6oo+sKar3RsW1G75c+1kpVeahaSFK7/
NLNL0bdXeY+LjSaWBqjJlnrmd/c+cacMN14Dq3U7ZK6wqFhy2aUn1tIuk2AFkuLt
9DyQpkgp/CxEbwFMw4gpRwytqO6Rg20jmixDSR3kqEnGR9Xc5Qxn8IZDLlU9scZH
ezIz6jvGi+IswxOvXIfT0zTfiQiNPDwHn3/KUdy/1Da1dtSCumv6EbYjiNChzYX8
Km4P93xkvDSQfZyIaO18/Sd181hnwKWnADgBSDG3kDrvc/85b7B3luQOMv+3k1EL
2DF/qxRrNmhPXoxueFxBMi8noTaa35Ns/Qg07Wa1YTwxj5vakzkgVHyjY39wg5bl
PiW4fQikbCn/seyKuatEmP3A8fCGz5Jt37nTxb3Dm6QElSZlrscR4mKAjUb+czmr
hFWPxIfvFmcNUXokSSuQ6hX5rCoQSZyoH++NjAoCwdoWmm2fH88+jcWU+yRjsv5R
bqYftbw1yxZZVemfkXv73CMJ80Cw+PmaaDn+Xrtx3P2xL+kIMFAyWf78shGZA2uX
qkZfBHeC1quwWkormgiUBGSVd08827zaiT3j6RnOqdh0gsrme78pjCyXLnTaOJQ/
OczcmezxEn4O65gw+XXuUXutheqEoFO8lJTy0e9n3NX59K1uzYRBZhH1e0T/15YA
ENWQckHtQvXWxn17GPWBA7LX1CjLP2uNFXev1kyG3GzhZYw+M4BI/uklAOPuMa53
7+8VYoWDR81ZNfle1SbexZkb/ToaiAc+9f13B5H6RiR8M/xqyPtKFd34pfx7KeY5
/CmGRSHxa8oW+dLfIb9auRRP0m21sxALYTjf14Jogb+LnuZOz9iI2X1B8rpBVVaR
gnPCDpuVShEQ20XRjnhr1nE5lFHUeNjuM87tnAAvB4dN8oako2qHI1n4t4dDzzX1
ssG1pgkegUL10oFVk7s3zar/iBub1y921nm8l/uJPI2MfNq0eUhlnk4G+H07csrM
GmgyP279EOhqIj6bj6DPytLz82l/I9zj3ffMeGC3AhaggpYCGbi9KIbuJdaTeRfe
ewZT+djGxzTX16zDCleGc5Ky0A1/w0LTgPk6eT2NoLcCQS8g2e2p/C0pJW4wtjs4
QkuWkq+YmLa+biRKQN9dh8loJ7zAc/cureVZw+Mcce3lHLYtCuLdI6Dz4GSHUsFr
5sAqG/t+XlNiXXDY1FWrpnjaqQ7obV16kOVLmDkMqDqDIkj8Y+iDl0JOpS+1IR0t
EGTL0ARm0PXkdNoW56yt4g2kSQl5TolV1oE0nJHnKmO7P4G1DUecY7R1U1T5h01N
bWssRKQJMpW7RKMELq3ehfJJYM95e6fZZLIviS6fAAzXxRFYKCGqfGFW4YmnkQ9H
6/yAFiVUzGeRQR4zYyqDYRBdjGWD2XxUnpqsIVqYz4Tcl40qyERlP05elnECZ730
XJ/qJuJBZCwBig4CwRuw0Utn7xyMlH6SGfEsmrxfAf++dXrJ6EYJww0M4ufmqx1s
rZfg+2KFBqk9Is4RauLfnVc3RncHRmm0c8C7s5ZvUSB2LjSHJJsGn41NHMj9JGqt
w4duu//6v1aNZD2cepjNKvw7glTC1Nlr79WqM8PINAJdlG7TH/k54ZROSdPsHYLu
mCS67CWgq6f79hdagSXAchvW1hq2ZEo/0HlymsxrJRfJE1+c8gTbEvGZYvof5Bbw
Vccy872f1WzKBU3m1Zx41XraATzTAVod6oZtgU+FGUEh+C0FFbK7IGWAcxwpncnu
GtFIOJv1rsqvIQ8zT+5pPfg7PvIQ83w94Et4mWAXYWJlwb7OvmN4YGFPF3v90xcR
G+kYL91IE1qmi29T3YzG1ZTiH92iTVINGptt3DDM4AwOi8E20DAXFR/gYtZV+I//
J/nixsvHjPXLqLDz/rr5VUmBgyHis3EvTLWNqqeJ9OD8TFI3vBbnWlKL4GmV2SmV
OSuBG9RHZlRYDVH3PlIUgHhYOtdgFkcX48RanUrtoYdgYlP60rrx/SFZdFBT/Dhp
5ovncTcB8apOG7Kie8ebwvGreoHYfktU1F1nyClvz8hczlzbUeTgk5SdgmuIKWP+
NvIOdclHt0mktKQ4bvaTQG1r4n5n6JgBQQFuhxMYxePkJxq8X668CpX+lMe+IV0n
pEQhWrNClA9lDrYtGaZJgMZ4e7ed9GqIizafmL/PKt76+mA/DCwtiYNtoHHRe//m
FoX1B4akGJ3U/6O5WfEJAfVw8W1WPa0jGyZ3aTRO2yOwyvux6gBxAsRMIzndyGkr
ROpP3AgjwW1RI2qz2waBMWfXzd6KKvp068L/X6r9GeofVp3ushDQ8XBLrs9wRyET
VjumIZXfgG5IA6Meap1+QsKyotg3RM8kkn558wmBmT/RlMT2tWaITq6pgi+1yNm2
3/c38DWX/7vSnrpj+qmNyCqPG4yh6ghfQQbOZ5Us49kHyAYnxvwJcNwBXTN/BDr/
auj56tbItdSI5UIq4Fn7KpHGfvnYYZHqt7ycGQEhGFMxcOPfLm8q/YRssG8nzcgX
lqIBSAAkO4i/nWNq7rcK+NRO2l+ILC9rjEWQvdbMJ2FeU66q2AFzfGfL17HJ+XPw
qTj5AJw79klfr5hW79BPAx5+w+NYj2MiE8lk2QEHlo99qVumV4sstM/igxxgCv5k
t4W4lHjJwiVIf0p0cD77d7OhHS7mlm3sSCqwdjWVkGZh3FoQKKdOD/3FZKN5Ltjj
c8TIN8oKWZFZYH2JSnI6nNkmIwPwUYo0hvOYCI141L5adOIFcdrK7W43kIpL3PO5
eO4onFE1SzUxgxVx88rkJrBPgZQNmOWDjZdo4w/G7eR85y5EnQgzOMMaSlwH8NCO
J3z8rfHH03De7ACxVEgRfhWH+IoeY5mRgC94NFdmJy60HbDiVPFKLnvallW/gDnp
sgEArDVxg1i+sB2a26wVMejJ+OoxOEAdodYPpfBZ3ZqUeEwUa+nZwfjtrYCSiFLM
yKDesYJ+Xzp7lO1w1lRQbvF6zVnjcU+7u9+FxrKf0acrkxXzAz9weLoCkLB2JxhL
VeOuY3M1/x4KlEfxpausHtavEUrsHnwBgTbRltj8TSWISl37Dg1uHIe/sgRUBqT6
w1i2Fi2zrDrSdyWqZjudzH9Fud+p+5VGqA1OjK7+qqtleonJcmmnqCutdulGPRhD
bICAuoHU7AB8WS5kS3s08hBH2J7LUMzbN/20XAsh0Ybv4wFvZ1/FuEndNBtAJphn
PHZbqoXQFh7pn1x2iFoHFsu0ElINwY87AZMsyj2m4m/ES6gpi3uZWKnCtWK8dXe6
GOtAcSjJMpINVBkdzfdF6dr/WlIZT7bigTdMg8ATes4GfwolP1LhLOn+sig9CMdG
xHSCLFYZ/z0kQaBYQgmuYQ5O3sLJj3bwQ0SKUlRqDBUSegN83/huoVPrVD+Dr87G
21JFYcBJ/ONIbN8PJEusEayWPFgDKVtX2mEd2dQyFKTboBF7ptdEiirvzGKyvWeJ
2E4/qyrXbvbkAq5q4alC0CDmQdxK3dqO/15w3bZyN3vvKp+GdqBabiy0nMQnZG56
/AKBL97NK27MHDmmncdrDQJYlKFdd8zRlUk3EJBkJ8rnnAAx968CIWQLCPmkXcm7
VY8wKM+eea9sFB4qtql7gTjEpmoP1IOw6P8EGYV599gwgZ0ovXYF1xnNgNvbV37g
nzf1XlxN2QV0+iQup3CCr7mEhW0Kt9sTzw25isUwOXxAhEA+nU2qM7xgTTgD71Bs
qceOHgn7ywQr9M1FhSPBANO84wO6TzXd+qZFHIlbfzt1og3VS445TaE2fDyXwFUB
AZ6A1btrLCKJkyUfUtbBcfhKOsG/Bguz5lE2olE9Xok+UzOhfhkgRyh7cWNJUlWT
KeTbQo6U9qIF5MF5KLKAdIEVIZWqM5pwHgsrHt+Yy+uAuTUo/zfRmWJMYgzFNVXz
hfkXC65HulcIcByKCiW+KE2xsGKDp7Mose5KKe3lSdD8fnYYgRv/8K/FAvBfQVvz
eHCsCxdXfxF09tO3VsDAmhyeWn3COoLZTcbS/ggAtG5SDBddBfAwjpilK7Iynk7b
24MtoFBnMWpTNlYgD9K9r57dZ8LwqQUPCbtj+yhdsa+JGaOdzS0M+8OzH4B42/bX
0us6d/RRkTDx93HlvbLimb5lpa0WObMXixR4EHK97B3WvorPfv4Am40kyH+zlVTi
jQEj4fPBmVzqNsuBdOTjHD430Iwl6W12RsBaJvttgG0puzeXyAfVaXivFiQq8/xm
yvJcjAUZ9r76/q5pMhdNDtPQ2oCvuZ8TutJNIJlEZRLObfX1nwm+u6cMPQTJwrIU
/j16uJrgvzVuo1tbaJMSWPYRRcKhfeYux6JpJ0TkPHZGX1aNEnh+lZMKjG6ZY3g+
XIBktfnhnjYskOLogC7dUNFmbHMMF/dDsHNKknRu42t9xTFFJg7oeHP6cn+SgxNN
QxO5TDbZrdxEIBvAqezXyR2jCo8UdehC1TY8O/PdQSLlITSLXZg4R5CmXaFal4jj
dUvoQqE3fljzUWBnQppchphp3pL2OwXZhs7hCy/nnXeJ+eX34cvvTBPZOTJRllBH
5e1J2TUFQLjCo5T12HlVjP5N0DAXKW4u21qFJUa+DdpEXHCq2jb2A8cBpx2HLFA3
sDZKHBFXyLD228RrLVbLlsxau4xaKtMcgCBPWP824TcBTRX+qeIfS9NQgheSDvv1
riAgGgyAjSWcYa47nLUMCeobMRedxGd8DoaDWTsELZR/CYaSliChCgAYqrdbmFiv
a0qvTtRx3VYHMayc8TtKGrRJ5v17aLdjYTMlA9B1gDg7Acfq0ZTQJmUpuqqkXXMP
0uDcHal+P6UqkrYDlB1M3qkgYijbfq/W3Gk2LKqF8teftcIXxINePQS0tsRdXc1z
XEtSgN1jF6R5kfrtoMLdBd2QGgicr68SdWEqRW7xIE1ZJgifhkzJuDf/SuBDgtxA
ZPrwEVWip5RdQcVACQR/Eouv57WWDfWsgn60Pk6MeQ0ppQdpAWeAFkKbPDBIwRYw
t8svGqwYBYTSabPUvzLMvGA0aWe6bpik9TG9BQbItCVyKn9jhzHruO43lxRUt5yp
IQ0IwLaMSWQV2ANXJhbL1/RXQ7uJRt7jXlIcqAOFf0S/YQm+c3yVJF6Vt6SO6w6x
A+IIWZcHCgGlLwaq5+GicZivGNtfV4gpAqrB+GxLwh79fySEw9dfcnbxm91diIMA
B2g217IizCKojTglYdaLWIxyxyUOBe3HMklcM2eZdZv+B3nL0fe5oz8ZRR2IPB+Q
TUbZ3s7cotxAnAZVAodMYE/hCvHIMkGWPkAo/EoS6VUvrvkJzkGnTtG/xbVqk7oc
DYaImzr6xxSqVDpLlND3A6//nm0jNIIBmG8dVavlstCG6X41dK5e050sXOkQw1eQ
mvA5c+PUCigH8dKx9gzaRaDdu4CAlCL5hEZ5D/4w90ZAi8n34jHTyVUWJJnhSWWw
upJGrr+CzjRxFo7JKErm3V29RzqaR5vh3a7EQv9DU93gW5QiFGptFz92dgW+1soF
eQTun3LyHTjpyYkVy/WxwsEX/1meKrHPBfAUkHAak8RGsO1zwjbNf0s/mBPnxN7w
o4rHKe86/s1C1bXlzU8Yd1Q9CXxf5XTDujO7DbZK/XI0uej6y70itX6+no+p1JdF
MAa6Chc7mahR1EhuayjK5fNeQ29I3gDAMPc28Xd4nQ0xAV+7BL5LOMZ4C9gF2Qfk
hb/N8z7NrH/mEmwDHPeCAVC4wzpfUKZXStg6MdFVpfNeOd6JykR09EWVkigoeoQt
ZMINTku6FB368zRNdBpXR5M/9O28CdvvcFMOXR6p2KGvUTRjIdJf8R/PZaus9K1P
yvWD9ebPzlrrlBlCumoyb5gTDNUVNBYMI62Zzaf7QwzlIUtnniWT5Q28HzV8Sznb
JjwIEDqu7cm4CRMFc0HxeUsYhCCo0/TXfXi2Q9zoH3CltIK3lKobkTan0y/S1G96
pWrTi4RwYSlwiC/aq9gibG/+6/Oq+4rRBo/5fPMSy1sAAH5jvFsdWnIaq34UXfUE
kV9E2sU8E6ohYxmAw+ax9YwPgUS4ifSeH05VJwCAG5fJqWhDZxVSERli7ziTwNnN
ALeDEZoSj2YSHparpIaVZ5Q20xGg0/0u6ui5TIVa+48Mp75Ir2/Vk5jWzCJNDo4e
bRqWimYvz9fyDi0jv7LOO6aNKoKowxWU0YXmZHudtT6tbgVHeK+fR17DSEaCCt2D
+QXVzU2fxxlmXf5+3/mqpp40Upf7K+5fQXxuOy6W2n568G7L5puEC9ag21sn04/Y
itNwkFlmXts88ByKIos0P5+HiJ4GaURv2lw26fgc8gEyPkmEmy0/ccaqEaLFNvvW
2Ks47kKwsi9TXCkrnU0ECX/h9H/gFpg4NjHqsb6JGN42NjhQ46Lt/CMWqb3Q20sc
Bbg5MK4QfwEB8vXbQBVnj0sx0mCjdl+hNPZMdayEfGc7xRjAoG94PZSIqQJnYyk/
aak9+pzSNoQdinYY538nGLAPnsmH3EHRrR1a2/Xyhj4PlF6uz7XoZuboaJA+ukuJ
hp8rRtpcM/EGgzdkncj71epitcta9ODO7beO3rbiZmxIcDALao7zbTgDov18TmKV
2b+eRvJL8WH8Pv+ZHSeIKh2uJLAalRz7FVpjFsiCbffSN83TSEiPmBOS4AeGGWlz
iiwg5yzZnTz/BJzECSLG/wFgfb8+g6altrdZeiPVE/aji5s6ymTzpP0UsFkF0LQG
ah/IvBOUh4AfjMR0pIIIfH8cCl33JHiBv8D67O//Ppw0oRthcPQAzrySOoY53UEX
TP+GncExHnCvippA1F9Zn4OJTYV711s6OE2My22Sk/zUm1Kh+cm1cKqDiOuzvZ1M
dUjD01TvmVOOJIpjcMiJeN/LVsTIFSdHIqHQkKUTsQ5mLHEP2e4JukoK7qUSbay/
JBpZRjzFkp7hOgg2u8btyuz6wtLFplEQAsBxpnzbUZzScBI2lu0GbTjOpLrl0NLB
rur5GSzliE9VbIhfXc30P5P7Cd6NnakxNxUn4njAki6WXTFyDUTOypNysWuQXpm2
cdppV4uUGuHQsMDbuxpAxWloXT5tHj06oVTdM6sHdr2Y0P34LeVncHT+rTR/4vEa
B9hFKKPyeubKjfowNJFT9j9DwwDuYpXIma+4HyaRCcPCA00EzGdxnrYAoAZUt6sl
+QsppZUaP7UjBfSaLDP2RVFikkjGSdBX8F9r+9xbd0weB1YoUZibj2saRxrFJcWm
jFftt67pWY7+wN2hVI0gZ6o+K4OtwRApHWXzKaFh5KtRf61xTy0olOGbiZgqAFGp
G99ZalfYx0KNZ9ZxljzGYFSq8xrXTrBNfYwoPINyrUeGWM/YXfpLjzCYORDLUdDs
N9FfQx17i91Mk+22rnlUFR9P7okwrzcRwfLMsJOUZ35ft+4NZKlQoMifl6lqPRWp
D7v+FrYYoJp1wF5+ZTZtf3L/aXHyOYveUjYOn0BFg9o4VWJ0v/vxCySj0CJ9fD5A
ngWqZLcIBMVw27masneMYcTVzWRlZipywy0fYkTbe4TcKKlrI9iz+1+48y8KFiEe
EJCmAIpqNA/3Bd4NQLe9EJJfYoIb+pJPqfMUkPminuoTDqF4Gx1hF0AQd1hoqQI/
gzS0YrAsmg0tb0w2JjIKVnBJ4eGJ9pjSPERFwYvfHV7zfyTWJbOwWdKnkmRwG/pZ
aJiTEUeCAypotXsDkFo3Xlf04bZzmjv5piUDuLtFj2rALpM66W2umbI3dVy+hrSe
df0AB+5IBOUXFhZQooRuUACRHpttPvxXJMnDfOgXWL8GwYpx12VxssJhQtXszeEJ
4Dnr79qO07Mvk5LrPAvrUZ8ztmvqapm3oSU5gIOJwbxL+N+mTgJDzv37QMUZjPe2
zNagii09xNU9YdFM94jeH4Nrpx8duBKjWQmoMhyvV74RroKxL7ImMkkUa/b5wUP+
bIIKopkNAEtrMggXW+1sZCr6jBRbuIdoSSNfeVxpopYDWKdB3WEKkcj19ZJ/lQpE
ydrhZ1qxKCWdJgWv8n7rEmnL9PPvKKakrJQaOSvUB1B5PchanhBuGAYagOjd0kD3
oU0rztBc2VR3vVkEfLT4+xRMOpsH3hrkWnIY5CDHdzwbgXU8um2ZE3EUfcPEB7Ta
KeozC5nENhuuDTE/kyErObU5EYdmvBVLePQFNFopO1sWtWNNJaZnWxYQ/GJBwDx7
zx3SdP/f70DAp33HPoZ9os5sDtm8dr7UzVkPzvkYh0eP4qlwaaRcqspep0qoeeYj
NQqNxzmJSnTQTUvezlqGcYO90n7QTpaBg1c5vyUfcnfqCFj/AT6VJXA9cFn5Pf6S
0Ct+PqY1eqh7juFxGpYKjoODy5AHTMONCPhMyP9gjWMQ2t391PtaQRM1o82kO7oT
sjMB6WzEhOq7usOgd3ILTuPZeftTNTQDwqAmnzDZEj+16BVhcy121S6sPK/rSpvP
Uffpzi1bwP3FGiyPb87sww0+pYibS4tycNPLK3getDQuJnJoVTKLoD520Zmls0fg
1BfoC0ZdrJFlQgudXTzYKuRJ/wiHYbI3AzDsm95wqZpAJWtld2aruh7xxEuFsG5d
y6HGk42C6BvdSOYo5Mjkkg1hljwWuBPjhoXweMkVQTgUg6p6LyR4/kbzZx/Fxrgk
UkJRFathubQzY/yWLQ2J0MepfGRYFOGFz0N9d6xZ+A9g0SPrPukS2wFhTnlVocxB
rvtXWB/LDFRdacy5Jt9vgyzH4MU5OvtOujJV/gCFlBi054OPXXb3937VdfqxCdrh
d7gGnsxunLzwmyeGAzW5LWnHmhRfOKffPVkl7ww3CkHyIFYh+LrXdRQEy8UNifJX
JXlIQQ/fSA4KgnBqyCYyzCm5iR5dPd00LlCF2kB7EWaw1kUespHEn1YiaUrVyLPg
LTjhsXnqknfuLFQHsONRLHDr9yXLsE2iWla5UU/OhDccBFkb466K/bvLkzREPYnf
Jm+uBA/rbZC1u1AYmdRG9QXEIvML69vx0yvZWV8dd4ulGajKO05X9uEKFVR+ymdv
eIt6gLEpNIF5YYodiLURezNfLtkHJ7vGUuQVpsZA1p1sGp5ET3dpjtrPqWkFQL3Z
YyIs1Krrg67CijxUpLer4wF/ZUoqi0o1Xp4HvDer9Wy7wAGpVSohdtgFWSykax/X
SHnRO9gjvAo0Pr+1+LzawMUB0uxqR+fbqpuZDZsYVKPTyiiUjeDQR/1VFvZOFbj3
A/fL838Og3DCDNiEqZFIrRJdnxE0FIJAN2HTUsjlADy9uhoSUT4KzPralWMt2GC6
1d+j/BWkUIaE/2btc4IRrzcyW+dBZARArU6bABWsi+Mes7wO6v3A417M/tiGejUi
SsV5jCc8zhfjkInxPkniy1Mezqbgk8BznV0pyObBAwC4TJ3v2CVR/Ekr1JWQX+wK
8Z13LHZOuF/ZnqeA9SoOIrzi3cHy+yHP91BmkB3V78BvJAle3qAspKWCe2DIBL75
NqMtroQiI597u0bvekgifkK0ZmsIEcu/LaWkq17JmLikPQzhx7gbgm2/D4B72wYl
7QwXxiKSYY5IHdGTpOtfQdIzsJQRIBRWc04depG0vSmxXva/3bI1OKwOEVV8cq89
N6jaSAJy4JRpy5jeSbuguOwkeT1lNwKcDRY0XhIgiIr87z6UTOpvvYTJkev1cyZI
PxNmdGM4xdloAn0oTJLGL/gQm6Yrm+di3ECJcmCEy1CJsake61AwSUN7YT174G3l
TY2GXnsjfYamaU98Eu89vPAZy1Tb+aQfAGat9kyQSjBbfRcIbJXClRWeac5zrrSH
6rACL+8FQtCDutVb989JH6RhvokuPe9rlUq7IH/IcLVSGIWNtn7A/a8E3MSq3vWV
7ZGhTG/wmrZX2xf8ZHRWcjK3Ah10bc3ta9XG3Bs71YetnwyqJUmvjeErlYFQZUN7
pkThRRwVhjTE4zSPEDKvUUl6EOkPzkWdbu4CN0pme2cuAzUT/Fx7seW/QiuPuxRh
hJG4oJ4CkOg45Dc4huTA6m2AsB141ge6cEPuzO482bRKdUCRvcSnVyyEyP4cd92V
IWj4vDcrBkYEqhY2F5Got0SWAoVPnGc9nXkH6U4FdRfJ5t6EASNoTdSO+OjAZnTX
4d1/uhqF9QOuR5msc3bPk65z+FTZBqQ4yGT2f8SlQ8kGm5IJVoWagWLagnxra9UK
LTT1UZoRAU7hPqRj5hTvIPaKiNXk4pIOF73UWNi/95BWhK5boI18Cw34Tjbcv7XR
zrLRuc+7yyK7Kkr1IRgbHbCv/lCo8cGqNS7xhSBncr4uCdZuRo+/0/5oOR0cJXXZ
gPpj6Cy0R5FbNJMj0KHGi1ATYF01SijNbFS9G492cW9/F4Yp5mOLsdhnnQVv06jX
KmaHWepomvWw237lpweDWW85ivDG1dMRxCTNAyu1vjG5sLcwEK4pQQYUOhHo5vYr
F8E7FbzBEfWxSaFcWozPXoMntvxZn7M7XgK27lVuu1GRhriepGRxWxx85+znhIyD
Hhm90cGx4FpyXNnAJ9mx6AfkSZ60gZL6KoUmEH3QmwgLg1+ZSwduGOhhWGvHWJ+z
BWsnVonFBPuEBSZwtVdOn6z7Bym5iZfob7iY7sU//OaNENdWg1gypIQAtbW0vXkV
JvUW+Go4aKSJ4HBQB0PIC4Eaj4nr/+2HPJ0IRlSAGVPfy7ZgYIANOHv2TlSMuw9J
zx8erVisRgY45AgSNH0JFSQem3um+Z3ZeBWZdxat55I+2SaCTLQXj3KKMCovDBhm
HcqkoYiwjhNvI7egtHuvV/hMFmecGOBddxVK2ZDDFkQtlp9IX4EfpxLdHVrZyXue
gVwav5R1KR1hlDMqWVVKIUNyAwIatPWkVu+lf9S6TNxD5yu7XM6ewLVfwkmzUvNU
9sciwA6z2vH3XuTkQEtEgRN3is20qD81RXOOdjJMu6V4PySoFcyQJPs/nd1dlfvq
JZw7c1lGECQcRAiZBaSrkM9HRb1LTwq7efjUuBc8qVNtplK5AvORB3yXfTyQZUPD
Fwe9L30o1MxVZJr/54QOa+8L0IGjsS4txsd1pQ84/Wgj/f8bN8wPuTOE/TVvKxQ9
kF46XdIE2Whum27DeQNDdnja99avjN64tCLsSFO0fNCCxIvIEzAd8IoaZV+PA7e/
ObxxmGGDh9MtvtW54595Hx2MhJi4fxxTB6AwARqKBNgjEBoekkhxZez+EUxOGWsd
PGW3dAY+h8+oGKj7adiuMntPkiHi8GaitgYfKxM9TSCuhmaJ8OhzX7hBQ0+QX/c3
7JETdUwnvjsSyfId6iUPhPFbuqRkPbvr4MxjwW4djxuLiB11iSaFiXkZvyL1Iqzp
wJvyfqQ63m67oa3lwkbFmyNqeEb9cUJ/yR+CLCO4IqmykR/we8LkzyOj/8nnibLy
Llu8gPaR7PtYVbATI14ttC+Dmh4kQo9YyD4PMEWNKs7s6p13zD0sIurzzZwpy3H0
YYS5OLg3VaxSnyyYFTvkd0gyxO2NqK/gB2fvyktZmfev0Emi93kda4OzCge4pBqP
A6M3iDjGQocZ7wmiyC3Rmzz8c9XmFIaeTHe9G4dLF/+v8UpUCFiT7WRUWLpLKEyT
loxMxCjkZ22idsnCOR4uOMnibTCjaj3wjrX79RTSAjy5UMGldrVxwLfn22frDcSn
3C0W8S/FXguy7qeP+Af9zEfaVTrKRPbHcsrlDAiCidiWQmweVNj1jdjabm+8ANT4
Au5tfrc9tdaJqW4+hfwscfRjpzpZ/DaGp1HZAEDn1wBy/awSXgxGql06WnnQMwMs
OApsF01qDvTIlfrEWkshdpBxaQeHLtmScGNoI60H7Isq80MYwS3q3qI2GcH47mEd
l/qKZgkaopw/Cv6DSRJNJDmJ77RQqhHnYdukTRJXTsEai2RkoHJVEIY+M09P76DN
vFNQhPqKfBxTsP35HHsOwa5HYEIgLvap5yXc52DPy5Q1tKydkIgu6kKawU5Q1DYJ
c3yPc3jMz0IHYUH/qkWT8OoxjHaf48UKmKJnCcX8vDThFU3CL2GnsbrKxVSh9cuR
QSDBaMUKsWMFkTDPPg25ReMlQLA/KMAsC8vUFgfgN4Y+CFnTAyFU+WR1CEUi4v6o
fWfaDrZvPvOslcHIjlFT+jVnDArzd61luhbRAqoF9C0hhonJOCTHe9qrq/EsfL7Z
7gZOHlW7qZiJHPehwICf1MI3LL1rY9b0E7IG+t4mYdDGbky879Fk5RgmuSJ4e87G
JMDs3BAFbBjnoRFGlB1YKbOHJdItgIx5fWx9BIDRst/pOcHYedmwA4P47MpF3/4Y
3qWUksyXP2I2AzA9DtHDSGjd4KH5WOVOdUmrTS8HrZnVUHvNIJ1qnP21/Ei5ocnI
WL+dE1lnM51aiNpLZsRlh5+oz9UG28pHLA5SokYUvV3JYW4oSN7kiA75cJv3eHeP
0we22kWPfV+dOTZZW0kjvVwhOMbw5LCqZD2p0OpJJ4mxhnKAi2rr4oIYGPoPbA86
QIVniDKCfn8lpdQPwGxZlyDeBae+6UZ7AwAWtLCSDaLLng3xeVPk0iiK3SE7d5ZW
clZF+mfwSAxJv58eyPkwLQmJhqVYVRjkViHIoYhhw5iItSTt/NC3Jhm6T2YdCLCL
ggOdwWx9Ozo9C8NW1kk8TO86O+IIirzPtfId5Yagy3+qEw9G/6ullpkpqPhH0YhW
N5aO1B3Cjadt+odc5msIDLv6FCRgB7OJhfPp2e5LCY4ybX+I43OMGvXam/UZZ/+i
IAre8zunB6qoCBGWNdFcNA6l0DjgCY6naXxAXJ/WKa8dPsgHiEym4JhuwwEEpGl0
z9UBY7p0kOh1g1F9lxUKjn4FjYf0ZAOQ2XokSNo8sJ78tj4rQJkF3NY3oIBRyypO
GhtILCIupj1JSW/ATaDsuerSdSJRBfP4wEdF2+ovubk9Z1u5LkyPEjoy2ju+WfdS
cFO2bOjrtmKPmv2yXIJ1TjLoe4J2o6hKkrfYzhbd3KQQ9L81sYmhrCgNwORrJROE
l6vPwK3qx7FFTaWW9/Hzpuupl+0D0S3pIyM9xXLyoo7JCoYQoriGAqnjP1RVhBTh
Ux6lIVBRHHxY0agT1E0Jsv60EOLAb+C2p2yNnVe5ObRWOp8ZEQ84HUqe6cdxtI0C
4QQac2Z6MK9gZWd5YiUZ4m6Afe5MEfuZJQoYDlax9kigoJ7zrRmbxPqOd7NSiLCN
QN3bLEgKXaGjDAlvmE6AMszltCTPUTBi8HFNjthCTwCQJnVeS2QrnIeT82DF26hK
iNY+erIUpOyWHfSuZDmM5Sbk3uvzq4YTlCCQIbrB0ANeWQmAkS0eT8cFHf/HN37I
Ve078DSIxEmL+vHArOvl6TS7jLOgYYVPYbyiNeJdxirl84g0ZtkyPXHh//bwaa81
2CmMQIUuNv/xvLejGnwnYkGn1+ALaywSdm4sVjWEOZlGNk6q9/RT/E+Yz7zEfFuF
mr4IOkipRe5z9Bp464fijApePUyKjGgGDTbivtOZEtBNQ1rnDXJaMrKVGhr5dAL9
BP2ebxHVfga1/l3PYS7tVU691vr3KtTRIERrvconpo87t25ccRS8UfwwIoeG5/pj
6HNLTa8jVYD+kB4/VHshWGYX9gAQXlMCgOUjUWJZI8sQKZ5I2PtNqqZ01bzx1KIh
//mFCHf/hMPtkwQQm3eoDi85eAEp1WoqMHJbDsjbNmT4ioL6+NXrKrTT5Jhdf064
55wuvj+UJfk0KVFI75LhRV5UTiYocY0k9NN2kIoAsYnn8U1ArddYc/Tcu7jpA/me
IyWUu7i7bf9x+MZf9cpr1Rm3QEBff7JXnrJB+XhCmJjuyzdYrn3u+P3oSFUGhSy+
e1NzOftPlg72VzLvMErRitCJssmpQRuBr4E5fTsI8gIWRxVLRo5eViab2bPX+kiw
zm1Xs6UcX/RXXpDCQSdR+onMCI+BjR0pU7xJ2/YSgqzb1pn39AjVxe5hJVQ+QpA2
i7G0NGLk4wnPgva/4VJphs0gIPZGiwNmh85ZsHvEBz0mn/6TzV79ux/D0zwLejed
lCyvOdhzmT8Hn9vx3WPVoYpu++7P1H6XtERfJ7IMqATSr+us7gl6AxzacrGh3hYA
k/3jeG70Av3f7OBpMP4j/GHGYNQqwfBtVC0qQj5K3eHiHsPjMx3a3edaroQYtNxq
FtNGB1oy2QYYyzWIUMAwgEqFQm8sXunBsPQ5NK5qxxumaSFfZ7mJBwspuw1bmifw
+bkV0BY62uw0A653o+1u14B7moNFGqrwqYJPPXE3jbmpRcQcIxVFqqU7mTFlHJcs
npZ5j+9BaRRKmfC3M2aQN/s1WvSrigw1AobxFBjJxAlMz3dP9YUDM6bInQ+zSmAt
QlANmGTF48q5L+o/OhmOg/cR4S7wD56LA1TWciwUN2BT07CC8OUAXYNXbYxvmboA
yo4K3g7b+kO5mrLMWvJaJ9ScswabQOwMNJOkD7yLbMhOGqRuPGD/sw8RKarHgWDV
GtttgSZoNbF0QxsKY/3JHxLD8qEqMBYOrq9QJPFfh6zaWl0GuzicVwTo5XdFQJQz
w2O1RayLxMXlHeMPbl+UFWwJBoqk8mWPTk7AgFC5+OOU3pIpOSZTl9GsM0xIwGpQ
TussJj1vSE10KxAQFGeLc+2KX61XCLBmLmzo1Vm3zxnykciHcI9K4CwjUKi9EL7o
8sUC2UX16BfCFz5dXBHBueDpesAVeih/3m71930cg7XchiYYwK16HYf4RLjwXXaJ
0VnTljSAGO5WIM5tvY6mHQ/HKvSngL5WRvvYrZchQQs+iExJZ6eqS177pol2NHrR
YiRwJJHNULIpqMhXXyHReF2vSWQ6R37Rg82b25OzPDVkvSt4p0RaMJKZbdsQg/w4
m9jAZ69Z9LdlNVFwGv5hLX784wrkbylT/thgCT2bZujfINYgh9HE1SQVVIheSxcR
Jh3dpdhx3tDWslsh3zoF/oFuWorhrArtYi1A5864W9Of6xPOutVHmiIsN0EDmkqu
ClDSNPjOrFCodO/iIDI9uCDr8rAM4KytlQHmma0beXCq/GGvrG9oUSboV5swQoIM
Qlm4/gpaWE8tYDIgCe+YoxruPsrmhFCFEZvSNS0gV4x/BIhd2xOI9BMQ9szB+vSz
sLQapejyZ4kACx4W03ZWTdS8Khkza1n+7PczxM2YvMdv4Wn8XT6Ya5b2NCghERnp
PB5PvP0AcbPaNX20oVoIL1juogT8xeJXbQs7/sEKarbTcnobGtFpU6LSQE1eVojr
AGQoHxpspL9y6aYQueCK6BFFNTgyc5mbQ4Wmwcn4Rw2yACnR4egJnmpE1FnREiPP
095cP8r/ZieH/Grv471U6x8K5xCY75U26d2aqmsu2FdLrNMu79jB42dL8rj5wQVf
Kzk9yW18ONAGbupBxoPr6TP4UOgx+Jq4ZdP+irLGMlPpnBFRM+os3bzgDZCBWqIY
oQdhtfSqa0Az+FcydZaUEow9D6UoBcZdQuPULdbz5KZg5olS11B+6b8hkIPSzeKd
6gABVlIpcrPPUx2HHM1kWK9p9Yel7iq190LxJUt11fRPvM2sPun+oCyvls9NfZof
xMYK27F9HaPCfIxxbtHEflejZ2inek/7Et29qR5+G72xjBU52TvUPY0wo7IZmo5X
LuHP2D3QYY35LA1iqbEIW6ZwsdTlvf3fiH+BKm5UwnmAdyrGj4TWzCK5+nI4eZvZ
7gIfakMYq3nE2hjbB5H2Fzll4Ko9Ynj9Do9IlysrdvvQYOcOBpIpkT4xPoWZjN20
KsOleWl6UOVDRKg1UkzW7ulCMMvN2bFmoBEqrzkxbVAo4zS2jmJPhMB9vxZQVJ7r
9wb10VQfehm05vPNXIsOXNAmEfJNHLkPnAzkpANWIGEnrZ/2y17Z4tZMJ0mb0gl2
LewSpAVHCVHCkaks4toQBJqpPvJ+P28VAYK+PYQmtoLKKhu+EGpk0qv56kYIUo6V
L5hUHtfh9D1twNjNj0b6wtmugo/RWcP4E3EW90lp499tPwJTYE7jWU3cC3reg8wU
8H1yu2sUynrhibnvnhXS79KNtS/J/EYFzH3mAWP72FwrHzzj0dLE2gfjeUS1PW78
nwGcUwKhfTNNUalUxFrN528FtFD3+BpterWhyrlBX4Bc9iD+/t86ygTLMSOpjkwh
M3TTLfcznN56NPDgtU8Vs7hj8UEVIFIdx39M3tcT9D1NPPgL20d9d3q23SRo8wJB
Ct6wNzZysON79o2uY3ZLHio7PJotX+R8tCO/JIQEOcF41bgSgnkF6d1AEmnrPptv
HYPht2lFJTpuvmMkt2ocYULrzdEJLV2o1x5ACqZWDUEAucwKv3Fwqo9g2jpZHc4C
M2IbwLnr9dpi+TNfuaNgwTzVKIYbb7ICM8SNla/b+j8kfWQtIMFQtBfjzrApgJ+2
TCofRUUfHC2muIvE3YIB+hZo3iHzJlZbVddbOvnMeeP3vZi5FCz9DCMe7nrPZzGu
n4DibBaPSR6oVfe0SSMSKLZEtUCJxOvIliSQnAh3gGNLelKZCpR/yoBJjylCcJ+U
y9XahdU5Mb7CL4DIXO9UL3Fk+qj6gxR0Y0RbSPx5VC9LOMnv6UlA3JNrNaf6BKDI
UAp8fsv11ZbkVdZeQLG7qO7i3m6/WQMlU2DildQuU0Ph8ECHXIUDyB4zKZuQH5rR
4scfQslwUfDquKRyik9mP1sr6hO1fu2XHb4tyTXHTVM6fyj70uT+2VwgFuUAzOUB
dgf+nCChMdVSVIa7ToMIEjhYM0qz+R/oWrrhNzV8x4RMFUJG61sjlx3Kn4asUe+/
1+QsZMx/czSIsvHZQTXUTKwZZ4yTHbIJqq0ZlqQ9oHUj2vIDoHVe3PYFi1MK3+xS
J3VvE3LXCjkpaqZ7VDA/tEsJvTy0BIYdTRXbcZWF+w54eieQAZHRWyeOZCiqJxxK
/i+3R7ZKIzu6api3wbMJEr7gS/0wrOzq6hryF1ImJVnLRhp34L1yFyCLCSojDrHg
43wV7eMZ/iTDKUuLvXhmkJG6Xjwb9RB3hNnOw5/LunWERojewIpHwWKwlk7xDmqg
0u4gxS629x4opypbnYLzf/HrTbjkpjzEQUy9KBdqfEnHml3nqhLyHGyqtvxNgkBn
Wns3MzmHr+3KKdOCyOY1jE7deVpCpM6dFYiz9l+pIId2Dbl7nzp0uEWhYAytNeAj
chWv0cY5JvlKbbJXNFMrTUjGaAUj1Jy8921u5u3/MPbiqWrZWEQE1TyJUUZW1t20
9KqmukYYKjveByLbvMkCoOWyvOsbygBkktAy/iXil442P3O76keUkuA4ebcyrTXO
IW7pvx+Xg3bv8VT4mWlimJuGK2fOft0M7lAmIqKef2449B/6OLjr27UdWfIzQ29L
xiroe45Y6ZCf4H15HKLmpfmPPUl6Zc55hwQ+jEYIP5ixCdLItvOBrjHNqJgPO8SY
EXz3QSRBgHadpuhU7gP3D1SdYzWh/CckAhJtBRy5/Vg7S7rOh5rhfW6q9L9jvVy/
7MJit2Lr/HFsCkqfOrCnpCL/SFpPuzgPd2WQsLzrUVqWDkCgzG6I4teT3X6/iYz3
ML7B8LYITZ+riMELDt5QDdKWCcQox0/y4DVpQrQ8sbWYWbRRHRNKIGI5dmUwoC/V
7AShPMGUbCNF/H9v5pNiRInFVdOMczn4REQ/EJY1b4nXzpbk12ky19clZRO04eCO
HleaUOtdQBimm0xHHZ7VOUh3aUUhEdJ/DH+9EZb+jhivjmwizs2wcP/6K0LjXLO5
26pg9carZPm3thWS4gvddKdVjRrGUL0r2o9jzxp5fqOQD8HjJZ8XFjuqtyGw7eOI
kaFL6S0MJptDoilctoQB9ylJQXwyaOrHO1sgbrjYg7ZLd2uLNrDVs+GFFwgJWsIE
azI5MpIUj9m3vWmEX9eteNaj9xs8unLTE9tA5IimetQoUPpb9xqLLVOD/cOXd6zC
AjInO648/Is7iQJjzNDKQWKzsZgQvxqWmKq3xH/U2Lmw+LeP2JFA8yTbfh+a7wO9
QBiLAMHUeJGFSxoiblCs+CckXPxQQ3DGiK/5r8U+PxKl9RcXCGdvpuO0tVVqRbtB
IYXKFb3QptKrLWqgm1TDJ1DfExnOx4IG/bhhudHARljZjC1NErPUMqy9XSN8HoOB
NVsGms1vh1plhMWNIFqKXrl6YnvYwlCZlUCUOTOQ8oBy2vKbWQSXL8L7ehh2YU8k
CyhpWT/19NIFuhPcsYflLRs7WW2uWPKIRnTWfTtGLWVIkxfdPedQ5hcMuuQhZ+qP
SDJyQ+AlzDJlu36uz4nIyyn+yUWTjDISsFTpikpWz+Sv3l64ndMW35eNixq8pXJN
xW3HQ7RHOt6eT/hNRNkQqm4ohqRB67NOeLsHuIrD4tlt7Qi15EqyixyqX63pvNcd
ldn/kdRmX4ckEWOfHKk8LeXb3HtjSlAtnwYrq7CI/MJVbBz69qs0Bx6nALcnERVw
snPxrKRWwSEYPPNBa7RmUcG3aCTgyVrgNJAVEMjl2TwnCftvjfYgDDOcKzaI1ZGp
avWYsdpro+Mz2n8QsYk6HUROrSv1oUduqevtKAGCarLus8z6SWK/IBj5Aqlfh2EM
u8tdzPQwIdDCSjcX5/caMMJlOMEO6k64YGCYZlSJ57MgqdXxjTAs2qsFlHlwTRh4
Q/gO36E77HZmZ+tLuhoHo6DGMQ9MQnZK5PCfBC8UBkxTsbS9wdmYtvOq2gEWIqB3
hdp6b8t+W6aVluGL4/goXaJACJsvSrWDZe00zDp5JzUFwRZbZJBBxVabKGP89hKn
aNNfhdwbUGsaJbbNxKUZmEArW+PQmPlpReiwzF7icnoUq8C9vkIerkHL7O8HumXJ
TdWiwLLIxRcIbBLlQgNwdsfJhT/zuln2RCzGLQuj0MWkEeiBSzA1CMc9I9gb/vxq
9O55TcuMsZmMAzOH2zW1zw+5CrqC9BFnyHKH9V4J8sH6NCLwwdrBkytFPHRFqCo3
RdN3NQ1uDNl9KiqX+ycRntRML6Zw2zYFn6m/TQ4ngg3u4isFWd6KzCjweJNOAG2L
xQ6EFkpHF+UbaON4w1VhuJYq4ulEZ1IFDOh/Qz50SIZBuHg9tuHK78SeV9zSPRwK
lxrq+KtzzRw03PDrKvjC+2mB6xa3ni/x8ebhWPSSvjNfRf5Q4Sj1gNaFPJNCedoc
O3c9B+2YfGmEE7jyR0TGT85rKNw47ogDeRJ/n8HFotYu5ZoVlpjoFeIVBMhms7jH
wpyaDbrfRr3xDAbZPChfRPSjzPPrVIkPWstLdhJpQUU2zh6eYp7pFX1wdLQVFux4
oACDALqN0Tn0Lm8jC01zy1EB8OuCR1mvhVnK8t+riDa48QIDUyZdgtK8gTGK41hb
1f3ffwdXgx9fZ88E4wlDm2OtPidZOg2laEkaYwGEHcT+RVD3oY9fqoXWi/Ta1PnB
iFzQGRe0FsY3aBIYZzV96Q24aZ7UbnBmLViaNVRjRTfJjPj8rN90JMaYNLaaVoYQ
yBwZUxwgA/f23E8VUEvG1CCUD8KHUYphtaMXqGUWh7OI2nRy4bJafXZ4nEpUMM9O
eyujSPE/LFxJ4qFkd9rEqD0FSD72NlvOQ3iyqdvdw32Br2bPPP/j71uZYt134kQb
P8j1KQsAtcnUc/TDRPQBTq/D2swU4z8F9fNWtQhooIbz0EWtI2joaHo8J6nWO4oS
xft9g+FYkelnglaeYvfKWpDq8bOol44qBXRHm1bPF5V3PvaCUDp7GMpP8d2VoHy1
Ks2pwYqZnbDjyNCbSDRnn3bP+Ghv7F8ghUqKVmMV5G45y77zWsEHsHF80ySUj43f
bjeDxP5ZtKIOpyRZeTr5kcY5bShri4ADp6jmsaNxLM30Gc8wNZ/qDNSbrcGznFaX
1CAw1IIeA9qHLmO8b1+DeNJSX6QmVvO5komZXneDyOkQ0LVgZ4NKH+1ZygpPQblZ
j6o3pXdvO8vh6kbxWXo3/Kzpz/YEJ5ZH6qt88u4vW5VJSOzEWg3TWdyfFZe0nu5q
pO+lvZV7gefnNV4nvtCr9yaws5OV85Dd3kmHAWR/9+EHhn3HxJGrunh+6QXpML04
S0thTAAyVD7Jc+Go4tyo5280ot0k7AYjiX1hcRGJqSL+9a612cvQUx7Rl42vS6FS
+0W2niZ2cqQFmglZlOY5ULx63o/lORsiZ9k6G4eNKwtsFgDDawDLLc56npH6LT5e
d5+I5nq76dPqTKx8Mj5ZSiIXUx0SJkD3vtiX0hGoifWn/6sQFEYWY6NSIyJGwcbh
T3QRkHL5a3p76EdWTPRTAWHiJJ1ic7qSkAhKs63L/11Rx4CS5DKnoIb7GsB6qCp9
3fNzqTQIl/xyXvOgw+gXL4uoNomF5xE11GIHpgS9GwEio5MqLb8OrFmqiuK+yTQl
8nkh3sOVBq46C0Ny+hqIneZVphcZGlaPTGXjXVyCbFnpw/nO/U2ojSN+PINR54IP
3K+mxCJFynggEr0xcLWRl6fP/kDaGa67EYjv4lN/7OjSqXBiixRNDoEe8FxwkRfK
eKtAkp/UeG4aF7k/1eDRT/tD5yGEysMwkWQdMNbU4uM7RtHQS2CwX6oGsr7IWDz6
CTV5ny36NGHubrRCPlAnZ1NUj6oWCa3MU2V35geHWpUDTZULWrVEghYdpFYV+N75
VF8texkoL4c/x7UJszcx6JyGixWRmCC0UNxIL7j1qwv41RKrjYgIpDSi+01BAe5t
Xg0GymEAn/XI6l6PmfjkQTdAcU1ZXAY6EksNUNB7Zyqyv1BBCneJ1SWExYmm2Bvg
G88qFmwxXtxCEv9xgR3jWdJD4n7lolDYkH2WSxXIhVpwocwA1RqCbKt9F/LQmd46
Fea0LhDyp3/Mu8mKNuRA7BYfubCHPJfUjW6VOAaQM70nCtQIQ5dJVW5gbDFS6YHn
dNmxGoU7TX5q+iBuVFER9v7lZNGMF1sBd78Zs9msOL0AQ/ip0FDB9kQPgN0LBevC
WK1xjtqg2j8Iv4OKK+1a9oMyQcV+5KRqMKt1AW1Jze7kR07smBUxjIz7Ug877JEC
hYhlfVteJnHV+ayfbWNXFELw+7frwf9yOd7zQK/k9JHTAm8ieBIRwN88BQy4K5WN
VNEL7Y0AMDtHYCRsx7sN3hKjeOlWGEV1OMrhMqfy37PkgLMLB5d2wZpV3bIl3LM7
QyB80OIaZNxcj38DT4afDpejnBGT8hjzPgRjpZrR8EkyigYup8+KquBtb5u024lp
x/ldCoINOr0u7mUpg0wbkziMldpx7Vd0pdqdKaAxtn3QMj2p93tUw1DO8GNhc/oF
8Eh6L58YnWvBPpPQFeMU5DFZxwpF1kSPuQRf7UFoTE/qEhVpWOODhuLhCCy8bcD5
KHn1Mw8L2+hEtHUMIiBhzLsIB3Zx5womC6xAzyHglJkFMxE3pycnoIW1TGiBcXbi
F6BaB7H858jTNdLhOANoI0EieDmrL4rLzMfqRPvtIVWYb/cno4nAMmCk6rIkOCn4
64Z++LpqGl38LhVdarNbccjz2fmGSVVVJDaFrX6PLIIpOxfSXGypi6Qe/p3jB3Mv
Auc7vnsmzB38ZaOrhKXkE+K5j4sY9yZM/59KAObFFYmC4TYmqPg2FWyTIFb0qN52
NBkQA1bey7nD7XGJfiqPXKWK88vjnUyAEKMPLYdCXGds/1rnamaqC+n1zN6Q/P9e
WZCLeO/Dh7sZZM6nDZZWaILU/UehH8F3UxOLTNUPvnjzhg2o/dtmju4TLpWZ4zsq
FjRyL1fRSmlUrRFCYWEDAnPvT52nY51bsPv/yQedIW/Fx1vIuqPhk2ZqrjvHnDFI
TyRQ7sxdAPMES4q85pYEcxSTZHRNog7aM9w2QGXX/RPt6Tt2uvE0zEJf2YqFA4pl
Rb0i59V6QBPNAPn47802dgpuSj3KV8LDuSyhplmyFByna1EfXCm5E/93tL/gJ2xY
RBt7fRBjkEvLjgBdUEjnA2l5kMjcbVKnkJ5VJPG/MuCJ/ndJIHjXfZ773Ji4psEr
LejKko/hjReV7jcBUGmWIQXKiXz2/zLFzSypJUmwUJqp7nYvIRhiJD8yToQSoq0A
NysjhVv2bzA75v/zzN5weZRujxfxA8KJ8hnHBIx4A+A2/7ESb+l/yDwA8obemN3D
0QIln/bDkbLU7okjK+6391U7cA1fBFOLy0uH4HCetUFAw3l9jdtB6ncMyv/tUI93
Kpv+5c7GYRxm/VGJazFRDu/DSro+BSJMVDLqf9EMEtwWklX77CBC7CUSIOYT26mH
BEQRLgIpf5JZOohcsclSQeTZ2rrQqOVufJmO0+Gdowu5K6HM6n0JDwonL4HBpd9m
NkNPzQb7+EZsY1jaHMaTQ65YDx1rZLHS9RlSVIVyaoQQqdavGjDPp1JFeBVimY1C
CUubJGZBHbNLh5FdnIY2ofJhLupOGiXu0fCeVsJuyhP8jCmTMND3z6rxgKPWzKTx
acqq9JoxhOKr1VqENOFy04FD6ojwueSX5aoSxYY4BBwmURGkqyrxD6aHUTRy4LEJ
9nOwepEbV/2azZL3add5zMwWX+EBFIgl1YTAmKWISL2oGVBr3iOg5EF73WT04W43
wS7XY7O2iwgt3nUN0ECX7QUonrhCfzYbkt6IaiVpQ02Gtz5Q5A2N3WqX/OAzL1wi
17u66F35B4ILm7wE7b8n80YjUDc1ZEUZ4lKlCnTZXSAuvQu8TPzF98gjJ81st93y
A+FuhZipwbB55GwiP41pDRY8h8L8yk8J/qsgvBwn3LlVsxWlZRCO8YQRIHoPtHcH
RkF89ideFgtDLLWzp6l3KojcoxXrEeuOO4YztQ4VMou7NLI6YSpOcX97q1uyTRRf
Go9Cf54+eNH7V2d/mw+m4vCjEMhDmGuCWeFjijOAAAYuy1m/nYAJO2EV5iCXrIye
oR6CeNxyEu91c2DzXsIZC+XqzB/YSUVTjSuuiseWbmFTiNvXjNkS3LH3OykUVSMl
qktATFtuC1cBiHxRi59Qq8o7/llDw9FF3PweM6gpTaoU3ksO95vIUld7HcneEfWk
OcRe7xtgtSi/qoZ6lVcsWhTyorKLDi/GfWC5dM1/ZoQNZUTUSag6FXBt210c6T1L
L169Nm2D5Us4TS2VLQKXhYkNcuQNW20b7t53HoFTb9Co0Ef+tfRoE3krjCgw9Zmi
rC2/Qedl7JeRTGZfXwpMR+1DVQMPdGnRpxuvbAibxJPEhXciwVI5TCSFA3rr8wzE
1fgqG0EfloNvgSdE2NP1Ps/9y5ikA8tdGgb071lX2lJeez0A09Zb4hhLQXWI5R61
IF4RYnZHd3tgWa4Na9I1ldA5rxtyg9fMEF1gjHtUcIV/QFuIeCyj0xwjRTQGNHgf
iPHhRfXdXEqimclzB6C233C/00t8YznTShuGVgoU1hl1YLMLB0wDk2fCw/4yit4I
lKiB2f6r9hK1SNRAr5PlygikA++OUdujCN+iLD8tlkqLuLpFFNIR+2KoddINQZss
iQamY45tqpjxle8psb8kwk3BE4HLl86iM9ZX1T1hPY4s6RE4bz3RoXTbyRVsHlto
bi8ru7ldTtpwkpTnMQhy8jAwslg/kCvGIwbrA/7bmXbErwdcx5klqMjo+KDk2MCH
DG9K04dXZ4zZwC/JFahDWtP1ubLBUCWB5gHyK1TC6jXT/lEnvOIHgpHzR+uailUE
YAeO/TYYF7IBIVZ4qpkjALsXxVrSiEvtFOrdHLuvTAE5DSPcZUl1VlhXQZKqNX5M
Epc+kujoIVfhe8PNuKa3vucPmn+HFU4ZqIoIGILLmAQsppL5ge+mikY+YFLL7nkS
g9scJo9Svou2HT5zUNK73gN/0X1PRndR6gtk/ul8RL85Gw4wrp5+Ll0/XjaDUpsG
zfh1kJ+/QG3r2vWqGc3p62mMI2Vayn4xHhKYVoXxkWeSye1IcJq51loeg+mppW8S
9HGYMl2fxY7Zl6OLvr/VfV1cB8leNGNuy5WfFlE33eHkfyL1CDmU0XMcjJMKNOFn
bUf9ydLumbF0JdT+Cem6oDsJw9B5Xoxu5gIJkobBeNNNVM/6rUrZMXHHNV7KlecG
JG6No/TCPDtFpLoqeJGKqzheVm2QcTwihDACx1zhUTSkZeEfC78shzIP94+sH1Xk
oFhUJUXIPpkn5jeyZAagXvAqFs/g8vxCg4pd2aZNkrPoo9Mnqldl//1bIhNviod0
5OZiA3dV1T2Ld9R8QMZptbOFW5T7WZSL4jLHdihUQKGUD8+DV7gRi2YykNpCjsga
nMAmL+b53Rqjizhv5KnDzlO4uolLZ0S93SZ5NbnTlr2JwW6rL/gzQmg0pU4Zarc8
sYkIcvxN95Gv7hbANiR1GBJ6OEf/pHDAvkqcVqUaXlqeJstnbltHSyV8s3U/rkyD
Gmq+cBSMJn2vuY8xoHe0zSxdTKNANQ/6vK9mEkbdm6w/P7kV72iH5Ry6Fh4NzUYs
uF5qqKgt2zpPk29GCoICI3deiLjIETdjayaAQcgSS4OqjyxgRJRPguCcHYsF9Sv9
Y9E7K8UIhb7UBiCcgfsS8wRBfxSWOZfZh6VBw0Dl4DiN1WfvDirzWZeNDZYPNUmJ
ND8zAC8OY5Di+tyyLik5GZnIULWMcWagmk9g9ZdE2654Icgdz4XuYgG6aX7wbPLF
EtaRhYOlZP8yHGYLEVXP0r4K0e3pmn0rl/sc0fDm/OIVLePk+67QSx01Nsj/NoQU
wREEhuPRSQOq/uFd2+KyuFnskZIGWYBWG5Lps0rfJSQlwTikOzfq7YMq3iLJWGmL
ugIUMaKd5KbfhKmzP6bXFBFLjaA9FFb2fV4Dq7ajrkryNdt/nIG3LbrvW1LeDTzp
B02ZpojK5dpfTjYGl8opcPq1BkfMYSPw8D9//u9Be47q7gh4UjUUXGU2gjBY6waT
QUSHZnv8xiAjuYomMSxP7qspa8OfkJU+Uyo7ra24+0s9KoEQ8WCiwpKfy+lrm4jz
zjKhkxacvGF4oEa65bFXXOtWDyCh1UiP4/z/g4LrEiILmt2rW5NdztkYFs0VKcXM
q3LGZ/m10tW6XWxZgzlQExYwI4DfSRNdLOFYIGZSad/dKGvWeqB7pSOJfplqbxHn
e+9GnkyUekep2lMH3SkOutoYAK5wg0acgVtub4Cy+8HCL7lWwlCykcBeZ9JJZIb+
Nu/dqLoeocqoJOw8TGKA05E2mr7vl9IxazRPNkCkz4ha3qK/puaZPbuHJsj6Epvz
ZLPNUUlA8rCA5rxA+UKPBRenJLec0SRRX1S9EFia4krOmvC76Aea9/Z6Rs3H0+Ba
zBcxfGyBhpTANJn7wdsXmmfRo5JVhWNTLWYGjvROV+3ysMYC1Wb/qJKHlT9ZohKG
M/dKHp2C8lIcZGk1bQQgmeF8LmQCsAsJF22M8AusqAL/tHV3jbglI+fnD2xPU9ZS
20c2ktKxWlVdJeKB0tTHAq00sj2M150zr620FXj+aNsVAJp21lM4SMVHpjSnyu1G
QLrMFgdKRyhy0HAJGGxz8OvVxf/9KwyiurOtNq8hVd8NI+GDlPRCU+G2Lss2mD8n
nMUxl5j4obkrGAXOFdlin66uhIKyG9s2A0MBjESlDtFHCnqgh86MhnkqtZdPdbh8
6rejZrsqN5Rg2yRv1g2ouRKq2NcViswVM3Bf/RiR5Q0gH9c/CVmaFdym5F4FvCUE
XbhUeIoQDcpLPw0VCrdXDcpwGFMURIxRlDdpewHvvLQYAe83qIt02EZJaAjm9gr8
6P782mWQheAL4F3KIRAK56YRzUbHwoDHPv6asuLvpvvpUQ5uCdDmDzxQ5hH/BTMk
8fEXKC2rV1FaYupagwwWp9jXmx4GEZyOPoxQkZDT8GUKK3PVpjoblIFOLAU1hU4e
va/rGsSHAT3R7Jj2FIXHutByyjgqoqZ18ii4mPB8opeDh61JMid75evbxixuEp2Z
DVpEEkpRJNPJKyFDDT7457wiIkpBkum+ebVtvKHqEzGO5PG6DQxhTLArMLA/Chs8
9nUiOEDjFUe3qpsmxIVDex201DQ/PoF+x8ANCa+Ye995oKjMOrK17UCjkdMp3rr/
9zriYVspJ2t9FapOPqMarW4268Q1r3t32BzXO8ehXj9LfGJEKS+kXgNVaFMe+xOG
zSM0DtX3It9ocmNj/kd/7oUz2Np+E4Gy8VO6XjzTO1TsShc93MTb7ANj8u3+IKRs
r7yo33JErfgLwhp596o/A8Ea9jW9JTaLEiDk+LpQbiAzVd5uKCKQewyR8fsYQRun
E+S42nUK/AWI85yGUJU61TXwxKyb4S9DvhfE4d/vCnPAL1TWtqH3yCWJFSnSCQig
cixdtGT7jXYgFqQGJxy5WCEHEx0a/j9gG6vrMJfESSQjdcNZUZf771RVV8dvolsB
aP9Kg92ICf8891cvb9mihf0bYEYIM+FbsqWfGMwtrEjdau7XrA+NSwtMfhP4ay+V
NXAWQSVzU+WIhT/DD1ZWXWO9Gz2uuSaF4AHapPQd/nIuNcz6j2zMTbASDG5++ox5
2MgJ052PoFOx4Jk+iYh+NiK10Jp0GIOIrwo/z/kBHxqjZfYKwAURR8jeT/cXvy0M
J04/qNI4W4YTbnVr5rdgkwDKOM794FVQJ2i9g1WtSl9N5nrD3AT7ns5mua43k7Cw
6cwEkpIMNLcmlnfl+U7pkCbDx4308d5bavmClqtI6LPWtvPhrdxNKwHGQNRcqhyg
bh2GHqT4MIqdUhiJUU2LpEOnmWuzcyCBkhX4wv3tRtnRDv/XIlbLtYL10jbWc/wa
Ad4s2yFdWEcV0KwKqtK9O0p2XPWTEcOwggWmlRomCB6SHSHYxXW2UMu3tH7u3ggJ
Z0YOwh6qXyFUQ0/WsugMZE96WoJ5BR0m6MgIkLVNGf461/dn6lKEWVn50/cN9pM0
aftiH+htYRS035K4sdFo+tiTThBRMYZkf3LkDk7RnPk9G5L55HUV8SXZILboghiF
ZaxOmfr8h5KOrA2fECckvUMhpvBJeWcCcBfLtTiAaPaybD6PkZ6M1frNlqLb+TzU
nn9SkFQzGP/amNoidHNqoiUW1dzd7/Z+P/vwUlGsd5JRG22rGrK2lFaoWRAUqMsp
U7E8zrNK7wQtZUJQqqcCccW+h0yxJ7hor5u1LHQACzkOD1A1K5obBXv6goRB5rd6
B052O5yBMRSLbpaTOjoUU8PgrI1RhGDJTbLpk30j2hH6LXUVLq+OWZYdnp9zQD4H
GIbn5WTcFLvL5HCQQ/9uyjugNj+dbQGz0N3I76tTF+2NTM2UR+lC7KpoXeeSNIG/
qKutSMyER0htMRAEURzFPdV2fPrrf1+Nnj29lQyyabIVEYwWsf1ycQEzhJPnF0ZJ
Q2+dIVgcwwlysT5aFJD8HMZ031EopIJyMTGHXEYMHPq9/xHO1+n237qu6izpsux5
aXQ/9qm0+kM8c8Pe/CtlYGctzbRkIg/OgqtTthWIcGEeYVb24krXwGoOrUTmAaj7
312SWngVs+67Pvj3/5IW95K01tJ5Z/7AMousdOLlx00sFgi2NTrzXRKqUX+huivn
0l/yXb7eIQsrVJ1K6T35Wfw+aCCorZxGyaCNnwkZ/T9sTKqISL3y2PsSmvAOd1XT
k/I8Swa7+CNkcXDqsJhbbfLel7IrFmpG31SE1qJhU/3jRMN0TE1QsruRdkKHVvCb
bpxDKjX0GQFD008g5fB8SCIj53916PSbxX5BS5eTbT9Ht/nPCFviBpxDcM1NbGn4
zpd1h/QiqXLFoCz9A9DkiZMsAgmnvs4EjZ1JmoDEwHtwIkn99VKbw11HDw2LfC6J
akNv2AcXAgV4ctGUhGldrEZbofScMfNxN+G8ANK9cgoZtyXz+ic521xi26xLz6/T
itsE0BkdWPComB/DmZwhcgnKEs+m8+r+dcw1o0i+cNAr1uhu+6M05XwEC9P4ppLP
vI//ztuBv75k3XgElXhvfwMTBdHse00wC/XdeXzUjLYKddqStEMVls5TNsHyAlYj
VQSYN2rkTpoNVbcgNdL8RL7qIx57OiquPRI5GLgbNWBASoJqWXLR4emV1jeicLzt
oUkYDNJus+fcGAIiXxuP4PD6gN5CyknvdNS6pdEfYk/4Dsbn0KstXURdYkbDnboq
twqK4BA6Zsm1DggEWJqvMSyDjtVvG5l4UlQL5XvohFkpWUzQJGpRp21Ror7BySVs
wHR907taXMEcHDjk/2CP6S8RW7cHKGzKl8oY6VAIJFrLtFrwkPgWXhAnLA2qoZp1
M5AsbqXW+lzAzGjxNAPnuo+XfX90nqWx9yTd8W7Ahc4mvMhcckTFFpLbH2X1o3Tm
+hhkeunZcWeZw9VH4AZW6iVGEQt5raH3OgHmvLBoyq+/kVqV8jJryuf6UaWs9JRI
aXJ7+xkfIA+tQSZC9Odys5UZ1mY8KKxHyNSByI6vb0zXV/dRDTIjT6h9kzVE2YkR
HGIAand4swdjYr39lVQU1gtv0mCzzaTyDC0aIIxz+TZ78WgGRRsjbt4ZZFgx//jX
mAVpDSfxulGaJkikzMlkw5ncbV1Eli3qRB8e/QqaiUagFfHIzaqMICxlwkVxk1ZI
B8supH4ZSVHSBvLnz2vSq3sMbH0WKnZmFwvKI0so6XURBpyGBwEqfrY8qpvVYc4L
wTtSkCFXCY1ryfnabi3n3N81EfmCbk8QFf/Fjgi8zzrAu1jcx4T4LAlqUk0/AyWZ
wrurXTarf8Q2veOq2YsePlO21h8GbqzehFEyTkzaDOoQR6IKJm/bxmSphmeSISah
xepwveg5B5gVOTR7Co02fJ0gRk7NjfYHqtwpoRCkcxUP6NWkVth2axMUeTASvUYV
hOIPeD1l5dMzOfeC8atrax/jl75Hbdp+aDCRU/DXNlaCvpHPXL4CRnDZZBIxpl06
NyidddPEaDBrMzbIsqQGdT+jLLsiLd1UhDualGNU85K3V50TfER3hflabtKQQe8I
s8cLTaSxDcE09mQ+e/LxrOZnln8KUP1i+uGs0qO6fPqCcXDS8l256XMlh6PM1MVB
y+B9Nt1oZe8ZBTt64xijDLmybatZ1j01K2An+5gbq+/H4R5XyvtOKNLd0cpD5+CO
Mj2SUNyndvPT5o0WS05+B2VK2tbwVCUU+Ranwyrs5AxzUdv3q4hX78NGVEVHLMWy
ZLn304mpj5gOwmt8hVTbylDGfvw78tcX2xVmC/xU+aJMCcGmMuTR+CKIr806aVhL
+2JeBagpKVFmoOM7Wfcarv2nKCOhS6nKpDHR4iBpsqoTxEt5sPY9nzYHPqKk3uju
Tzp1bmww14wKXg8ctcs3If+oxsMmJTcq+tMLiCG5z2kbEwCmy2P0BlfyRb77TIR0
40vfLMLAZC3vJZ+PHMzC31FabBqsYA1UiwV9PrcE0mDIb5kyOx2SXatqBLfBpMWm
N56JKpgWQdPUx7+vESCqkagaho70fImCARRviIO+jehytw45e0NRQI+HupfD4pof
fvO6Wd4kWC0Zeepw08llmImAungDZ946xRKuc0Hrml2IsstHPE6tryZA7Qcodz5Q
IQTuPHtsoZkgKKWOqDShMj0QD0qi6tYu6bs8NIEUDX91t5Xtu/lrbPrbfLi1daa9
G6d6mQKk81LzW1g1Bb5CPtE7G4CJAgatQRhlT+yVZZUPAu1g/7WN9McJ5EpG5YYu
1ipWh82z5AlHXPrkfgv4OvmxnZWCY6OnxM8Jfz3gaLZWzNf1mc8t4MEfYqJpL8ni
ll62pQK9uzhpmz/3/waFXMV0J8dEuZBVCCCepPAPIhjU5GSVPdUJZ9n5ZOSdhMFu
GPU0vFBM50l5dUh87KtG4pHXSSyX2yyyLUNsgebZzJvrq11oUoZBgFs9MofQalQG
ePYntDdAfUhyiQtAegtYkU4+D1WC34ZOAZk+XCBhb1m9VrrmqzAwylYfxcuo3Wy/
6jt29684jeA/8br/eniyjqsmMIbiIWN9z897AD5B4A0YJNXrF/fjMPO7QL1dQA2q
mLo1No6us+f+xWpu78wvWxfAVh/+adCsC40YMpT4a0gzouJqNbK5EZDiIWRVSL5B
/XC1k7oW/SADhsBqPd2FsN+ZA3dOMSsPo/I8UGXF2RZc8QoT8wI3w7QEd1rEwof0
ba7E9PouRoLAR1jE6XD6clfO7a7WfgedKwz07yxLmaLWu/LnVoX0UGUp4bMpBmF+
kT7GtfHF8PgQpQnjeu5BZOKxCjbTZ42WrO38inyvbLAQy/JKcN+IgwG63946BxNQ
b3+kV899vEh2v8Zg/mZfiPQfSK6SqWUzs+MLOX+m7UJgjoMRXcnAvfeRW4Q5wuRY
GRE6pkloAac9Z0oL3oWnKb3CeErq1KqrKXtN/iaT6WpQ1TrmWJ43k7dbIL1QAIx2
4BHd+0mELRtadzffkgZKizi4vQlDfub9tZecL4EyFqeKqyOIfIdVfZFF2edVMyWw
H+68ivpOxyi4W/5odMJvwomDrqJIrBlArnyg8FaXV2efcyXhpaMhigxDbxEPhhCM
fwFuKH/eR8nEqsvJ91weMLTxIVONWpUnNG+kfO65gGZTZiPU6GEw+dATBsjCExDW
R+A3Wg4bGL6lDXC6+0y4BK4s94QuSZTA9mAF2w564Lz1++idcVTD0IKtF1tmABby
z9lrccI2zSSc504FPZikKWea25Vbhcv27+mcg91pbn6pVEKrt4bre6UyzZ4GRIGC
Ok2b0N9w7ZpgD6PHcpkAIO8EKNMAuGNvzxpFxwD106+iuAlL/PZYpmc/tpccioF1
XkglLgc4R8aP05MziVnNnTGVwBytIyd7Mrsl5D+87JW3wbYWMoHtPEboUUjL86CO
+V16v9jEmbTfEoT7/Z1q5pR8j94UEDkm2UoI0ZQR18Ds+y/RQGZLWZP2FiuFgxCt
hMCChhN9piq8dXoSHclOUopL2uqZf6P7UNwkQGO2tXyhTyv5q+w1OPDU4sW83prt
GrxDb5DHyFEiDA2vxgf+SrGqqqg7tFa+Gt2amuNYxShVSdrqUbuPc0rq4FnrA8sm
BM7sGnKHKlnLaGDyIQmWeUBVfhLnAHv1rhhBYMCDK6iqRkmKZVoghK7O3XYmjch2
a00uI+PVao8KjWMcYxTuQKT3iOaUOeVUrmmCKcdxAdNz59mgwPKr9jyjbUtDpHcv
O7uws2LBb6azOc6Ia2nCFqUWAJ4nyTeFKYywtW9bnXDgIAZW40kSk+qIiZlK7V8e
9kNzSykBIhZOP4Gn0PaYyBgRBuIP0c6H+zQencBDbWateapHs71+U2eY4O8vikRX
/3BW0sMDjw2qCw9QNbVNP0a/dgUYImIkRRr9sWkAWRIRM72tBdkt2fEcXPe04q7g
pXfYpUO8aDtmLlGIx2WmildS7UMt+KodMUMGbJtHa5Ux1jX0x2U1wQWljqQvNmF+
UIWEjp/XncRbWxPwn2bBdMcqKisAwQ4497gChg+6PV/yuvI0E/gsksb+JeOZujXq
SNjc5TZ9h/J+LC26XP9M5gdMKC6quK8lqJbk+PCVCbv4OeMi9C/xhJfR0voE+c0u
DAvKjPqiIXgpyFPVhrehogPKczs4mvfIAUJKpik74XiaRTCwQMF66EDfmx7V1Z9H
q7Uh5SevLGtqrFJSpOb1b0uiC7yAfMsSfHGHayCCYElj2+4q+eLAb0nnOJXk4TZI
blFQhVw2WvjQJOrVtkl+YWObJNradPMT1dQ9lNoPB/HLj+93LlfkfQD607SAahK+
JYJLaB4KT5RQlwZaypI9GHOF29D54RYWSiV2gO2vArotQuYkWsqGkOWmy4cc9ypR
IB2h1Gq+6L5AvL4XugR0gP4lwjVH3RiaspmUNAkP8nA/4cxZZkjWO+2RN4WKhUZZ
N5XLJMDen5BnzSTYA7XB5Xa0SGdV8tK8wDF8FciZtBP6tIAw3qWmd93snqeovLcJ
LzetO+KXKgXHfEOPVu0NoVyz91kcy5PozJCN9V5NQZ6yf4sB+6SvCzoGwL8PsRUb
LgSpOLe2ApUsu5kC8a9eyp6o2sGAaFnVCqZhL6Os/w4Iro4i95KCCKtDouqqcY7f
Iki+QsBtfLTi7loWKdnMibiw11UzR4B8mJB7JqP/s5MAHGZNGyZOBH1TuhF9jZJ4
8qFMTahAdRGu/LZglpItcq+JwvBm5pi4EWEyyx/Una+NJL2ASHIadPw4PgAQZsYU
zBUlrgWEitzBeCx3atnAvwddw1yFVGChXimBFZbDoEtbM8QVdq+pf6lHoOKfHmGn
08HtUleNkiiEE74TzLH2BMVwqWy4aBW/9KwJ0ymbxgTDIiWIduwK7ylyOSVVZg+8
6SukdKogi5QMD2AjfvsXh2+85ckEIzWv+qRiXQ/bWddyn9lNuYlqSmY1eKFLkMp9
vSSzzY8LTmD6uXJuN1vRU4jTGjS9s0vRJ/DFYDvDLvVSLzV9aQXPXE6A8sE9sfl6
TqldGoPYsAqSsK6DN0ryHeFHSH2OX6UwYKElImTfTKCenPt6mkQv8ePHK1BI56Ix
W0VyFM1RrfJntajNPPCA51EumBSURTCr62KZAy6XJhX1BwE9Ewjrhp7T6Dhc2T99
fw+x6nhSKvEOKzpqkWZiqX/kb2v7nQh1Pg45gg5HOadGQd6TNzDUKzkHqxUKIsTP
CiX9IECw9G+Kf2Lc+UzRiDqB1Zn+zYDJdqTXiZIH5MMT8wq/OjTmehPlrGlHxShD
vg8Fk8XCDQgZBJWP5JwhA3b0BVjzteogERbmP7aQVwRCv973qMI3hpWiaZfaK25S
w9LgeDDnCI+Do1awDPkq+t+Zo4TEM2k3mTqgOtZwb+aZG6pYW3oNq7YFrcyBH412
KkGlwHi3YwTRd0ar3u+lGYA0R3MU5uNjZDL1xzAvyJYXW1X2i0rgUV5xxyWJ6zLS
9Loj5U8XGyaceV73Sjatb9Ao9QfBdAKO5OglvTVUZGCRr3mF6YcPuU87vP9V34B8
fy6uBUgI/mjGipofIaa/zXMrlx+IPsgRjU6Op9mQIOBiskgDqXaARKoxWjVcrK+F
TN/wqcpD7orSfk0n/gPKsXKL6E8xwhNZbzqSnSrs231DS6Hz4BuGJmFn0CLYwBV4
RNn91Hw0UDOh4CqdcNHjN5uMmad41W965GX99rL86JL5WAVK5mRgr+aNzHI1VvMc
r56f1jLh3I04A3scgsG8mxtt7VgAioVD99AhDtaOIcDobLkKKafZzp7+xdn2P5Hv
ZSGizPGRkY408/L4vbInCPPEZ1J8vL0l+FEJOUdJot3FZkdgyG10VMsNFtjeIy/E
EDVcv7tTRWAkkJteeO3y71YD+QI2UP0o4rumO4mQVj8DDhHb+WJsViS5t3btL8kk
SykW5An32vyvrxaVebCgLZAlYGCNmeLovXLq7X73VZiNbwP1AesLteB9n60SH2YH
84korsZ15ST+JlIK3tWFZlvhGv2M9dcfl+xEKT7eZyj5vs8pvXMM2EunNjwPOa9G
uP8LhZ1CBpVrGWM5JX5wY4ILb+n+CnjdetnBW5QnLd9clS2N7vrrZnde1nchFQec
f8Ki6M2drdw9Q9pp29bU+4R0f9wrFIB9x5brTotmMMPcIOgqtAvIf453zKgOnpW5
nhJDpFnLu/cMDcMPoEjxFc6rc5TOdYz3labsfImzHlyQnM/oX0I33171nigaoKk6
UE3TYrIMqJU8w0NGtid9ewyP79xIjp7l9jMLauYE/6QQpOeEqqUXEFLBTKkwqq/8
vQWKGU2e+IPmxCJ6d4PBA1ANsp7p4WpTxLAPvtlXSg7t++5WCPhNfbmduBm9QaXB
7KHLaYig1jngrsj4mMR0+3pLDw1G5y+sQ2lEYlGxLGX5a5NWzQySv3qqmU5uvqnn
Tzd+2Ch5L84UiATc7ZdewfVKKZbWT8BXJ5eLRK4oBIpv3PUqDdHHE0Qkq5yNZLRb
jpGFyQigTVPQAowI0Rkvee8WvgT6/WKea/FbuwFbM6EYJX4o14C+d3NxKB4Ep0p0
7ldVbxRo+J1pl9Zl9uXka+g6MXSAxtZN7iQAPvhbh5xiQSxgfZgtvUjq5E77Gijj
S1T0dRlwR3G+yaI359AxCNaiRkcDSS1USXejuJBJjMdjznDEXFtSsG5mLbhOsN0B
8fkDzCsqmOwhWADWFAbiv9rBie30tJdg8TmK9bk8AYFO4jzHOetUhA/zdhxXyGYt
AY+SVJPMyszZhFX4XWWDFlef71kLGFB3HOwRdkC9S6jvgpRT/v0wjchmd6lgTr5f
+xeLn5eyV1y0B6KPo5KOE0aSKZs4U3A9pbuJtlYpJu3fa+06tlrw35PQLGAWgDx5
0aQorHO8w4prrWqW5KkbGgMJ8APJ8XiZ/HqYWHm2j9Ug9KAwlp/+bHHy3iv1tsmC
nGkGoU8X1d5deXjZQ/cGbDYXHSc8hzkKDlQw8Sw9nIRPZAmbPc8H+oX777nvPNn2
JH6cS9tUUvc3fD1B57wA4PMG7I7AYU/GVRjwUcjR6aPgf8zlOlVOco9dB56ZIYuL
u6LlNt0hy5IfEh3i1CTChZwvsUMrvzN7aOFUOEZJHrZ9z10nnxT4GnHID5P+7TMy
gCGTTkJg+W9KKusySmHkzyB6BvTBhoYES2Lj+txTolcSxRKpCqKNQ9/TmYNd6yXz
bpAwFjULdXt0cE60T9R0Ypie8BsXg44kErC62FLzeV6AkQ14Np/uZfDUVD0UFgLb
fdPj/en/shzmRCLXW8sTa+NhfUJpnA96GHupeh/cP/lcKGRPcCUfggwZHddul1xR
j7+HnAsvQ1TbBNoP0VfUaULFI46+xfRopgZsgDkYIE3iIIp7EhEeCQsImiiuBiQf
xhOP/0Cnwy/2cxBXSEV7Qrc1MKPMAYVzUdYw/ut0GDC8IlL7equswgZPVa9yd72h
lIQ+0W8Nx6fz0RHqO3MP+0w2kBaaaFKZyOGivEl21nxDYW+ndpSu38t12aLU+zqc
LHv0SQYQtk+R8EhETxO3eTmW5qqZ7Bko8vFDe09hxDYO46T9e7B9c3ZgZhEP6vKa
F567ddygMfj9bN8NHG1NKdZjbbUU3zUeI2m+2EEomVppEopKwCAtuZDr0Gvy1R08
gu14OQLNkXCKqagALRALtJOaExoEf4RGhLn324rhLs6RE4kyNBUYezUCRfj9CsqT
2fO3eVj3rQIFo4sy8Mao+glw5BYybMXTH+Ur5AlhnC8Wetgdotq7KuGGxMLe507H
qdUuwHvrs66Ci3buzP46BLOihrLgyU5Aak4rg5fEHPyfEFILFFJFIkTYYGj26XTN
NZjTtmYYKRyCnpwvZPDwDM+CJWqi2eyHzaNok5NtuBzxfsew0eN4HZKb2DDOvzFD
uzBSRI8kRxxfUGPU5pO0Fz+MyqMKjBFbwtI7Im6SRPq3S592KLrOdc7esDlUVDuW
pq+wfEQx7OLdmPO8bQe7+eBe1SDMizf8X+DCTZ2f11jrBCa1Px4iwS+R+4spSggu
6T+62lE+lZKWVa4TcBTavkKOYI3Fd9oqFgMUzpPR9eS+CJoq5tCThCTHV/pZq30Y
fVb+bd6jKD5CtODnHOCTUCP3GhoiUXQ0pMrvPU6Mxz1e4lDTM9KMM1ONwnrT2GF/
GrdXwuevibsR3o5J4qkMii186+DsqO5lVG82Xj31Hc2VXo2OWuL7J/w90Mj1MtKR
XEb6HXsFywUpNlI/Dyr4QjQ4gyFErPAKJ32NtIWMlf0ifqq5cW+JXzvKLBWgipX8
mwyTY+flVbpBTIxkf5j8i90zLIMDDW6Ag7iU2Gqlqhj3dobnRvS17+goutWTZNnG
sXm4RWxmHO7sdd9UAsBnLLq1pe6R0oxQErxOhbKBom/znn0ULU5dMUEZT0V8jKMQ
sWaRwYcUfNfqtSCCX9+fcwqBbNXw88K3/mCNgG4S0QqP6wMvUkrTj+51VQOjtREp
rjByo+27FzplBSe6Jla2mqIMg4hCdAMrSbLhJHzoU03T+VYqIOeKza/MTfw3BHe1
DXFmU8MKETzcblH+VvFGHkq572gAuPLR78y4XGFFrpYJ4poDY8SsaneQau0GP2ZE
Hl7+1UxS9FpdJvhie7LBY47qRbvEj9YTas5R99J/fpZeTWYYgD8Xhin8u2B4aduN
yJf7wFTvs05fJDYiRkZdj0I2wi/jReiG3kqFwTZDs1LVjA+BdMgMEPg7tmrTCtfT
xiwgJX/K36l0fftMQKJoJHb0D7QOT44SR/EyrEgr77Z8HV7RsXwuGtFIDSASiH6w
JaBa1YRwidcmjSdU3x1Q/XA+QFjL0IR4A3c4VK8ApN8DryWI10G01P7gTiMk40l5
AOJu8zWvFvpzOrMOmb6OSy18GZHwcnkZ2XhSvn0u6dEguqv9epnhZN8ShlThz62L
24hHAfBuhX7y5VF1iXAw+RoZsMTI8Cep28Cu1TCiewDZSmbTrCCxYscF7SN5T5W7
KoGwMznvYzBKExbRky2SLkOlKFohSoUEY60seadr/X8nQC5HIpL9qB+y43bM8Mml
BzHxtgtYIkTJreKtBRqZEOr9UKY8BhF4rvNVbn4Fxgr2iQvuWYGn9ZmGrKhIkU7h
UweIsXQzhvaEOA1w1IJKd8Zm93ZjMgRYhmV2SVeC4mEpXLPddBQ7p+a87W0rld83
jsyMkzG57Ij937sPjAxXM5AutCEMOkzW2WtM78RG3UbDuKdWSUaZ1RZJugqm5gyF
hgDhNaUpFv0zAIhtA12TMrKW5d9kyjfi0lYFamam13x7bFCSezk+sedMfetl3vMH
nJFcQDVgyyUwr/44T2qtFrQWFWgUTBXz5Kr/aI63rTAj3UQ0V9l/7l78FAuH+BEP
LFXEm+HwDLGgChxKmNW0czEQiqSYRmJscIuiKcxj6sCPJ6jZ2Kl4Hcg4HR3zGv0e
R2klCdfGUFSDqThsU/RE4bQKbjnlERlDdNFnSqkgraSGw0lUPEmOEy0H8f2f1M7R
RlJSSDlAQ7A8PoEWn7zdWmff/546bN0uphnODNLCeWZsy0BY6GS8kYS++bVH4UM7
1QdcfC38d0PeSZ4lEAQJXXNs4IUgs5UKzh7TSwgmU1hQCIdnNVAMYwTQdJ7k3Rgh
zXIKaj/nlVwlhkBkt0Fz3sqNTjz0EMYb1tVlJvB8UhfA/mDS2twhITqOWWOYBE5r
B13B8/kEMnVEbU4VrzSoiKfFpY7z+OYcE467vjz5/ESLpkkv1yxAniISyB38WZan
P/tA1b/+f9ubu8Kr+t7zdzNl1bMy0TsWZn/UkMjCI+Uf47wP2wP9/17oSEuAoyRN
xGE/ga9l7FQbnA9u/LUdLZivsQvCSPtZ1XOAMW/uAyHlsHVyG1ISmMC+QzKLNUEr
xr3n3Ypu6tgR7ag5bI62E2JDn/693tTEmahMIiA6ftq+n5isDOX82V/kqsydTTMR
TGG8gg50ZgLx4pi/68GRdIBQj1X0Xc6ZusefGdAwiZ/lyCvxQSA3iCdueHmWd2Ej
HUUri3r/cb+BnNopXJxc4gdm7JHgVlf3P0eXi5SjG7KMV+6uh8yKFnc7t2wgiQC4
9XokL8rSbPlQNORwNcxgRWOxcgBbTbsiLVBheQ34rYbhHX+V/tUTcNpSMfpFT5SK
rQ2pnCaIyxrqaVzeOqMz7ujAiLr2hBflzJxN4dHwKRBLDI1RfJ980ci2cThoqPHT
JB6lD6VJlVv9a2/O9Rmrhe8vJNjcfsdjV4HoegdMD2FmQsf6hFCgzpb0DqjFXujf
2BUvs3j8/hmgK0IoV0+wAOsB03qn3csiKDMfl/FYOJtZFXN2u+1p6UZZGPL7WAIR
JAXRmkJrVKn2KxBvXZqoKC8Euwdllbh7jqKJ0fWRmaLdTaQ0vgSliiQENkizX3IB
LkfOuRNdA7oJmSlFgTa3BX4PDcjtr8J8DPlzS75hwDyPw0cuPdH3EK5Nvuxof/vR
K2uB9qJCnyiWCUj7J59Gth4AC9oJT5PB1YQmW0KB10LojbnhAsuMAR1ZJ2/KIkjz
ywOfvKzycr6KdW3T9R/zdVvdebfEEFEd66LppHt2qgBTAH8SmRhsAmXGJlPZw9YM
W7BLLLRtxG+IDELpiwc4izlAtOVQhlX8C63GpE2BgRwtz7XVO5u3Akp2hSPUfoM4
SWQaa97EI/ODZYGOqtc7ul9cYdX8UsjtXvPbrQJJdWTAJUTMkFqM3yk8iMhb7iZM
yjdj7kjHQkMiwKsF4azscLVmXxbUv7nx5IQiTpTHwhRc2OjGjw8SynaEAVj5FrXV
Xq7VBxKM0LwDR5kbMYb0WRgeBbzb/B5vpGOmprroUzkxvs576U+6GgR3fGZKSPcl
90fKLOLXG1dw7Y0FjPDFMgS2Bk5AQgMK/RO7Xuuxf8+WnlgSlt2I85xbt39zAuQL
KwMwuwIhIldp2rDmMptIvKMgkQ2plvtApF0Ubft5IKwgXREDtyhMaB8iOGAqTebb
N5b2hQUJr/OcUZDhhvGa8+IPMTv3JfHYaA7nMUYyE4GHwF+n8mFqSr0ANXnNhl25
qxu2zf2qEmwRI+/+git2raL3wk+PtZyATfQ3IDLhhWDH5YWu6Gwi5UqTSYBwPflW
SxKh4IfRMYkiPBqSskP8C5kn16qHT84HAvcQ9DdltnsqewwWyc4Qa08elSn3WTs5
Dqmz7+outslDVA1c2LNH1VVhrYpDynXUIGvkMpL4v+rDbPzXTc6ouuWxkhTbf9lt
iFs1vXAouHEKzA6V1BYukep8tS30Lzm2KMI1o5eniHyT67ctB0ND4VgNZWIyZ84J
gwWo6uDmIQ0IQMDd7Op/vvCei76rLj0rBk5SluJFi/sfrPTPbLcl/nDcxhWbxogO
y/HrC6RHlBKWZTnRwC3/PXrnWGgQ6qcoMioFs9MiEBtFXlKgPMcpXBQpBy0h/srm
N12vKsuiW2EzZCdg7vCdicYuf5BmuThj/xOb3UUBEvwhSdxoe6UOuoox6MZvVrRO
ChrNzhNUDuueh43NeWrxK/8Zsd0J052ZXxeXbfJS2FnibHoM3zy9v/GDdT3h3po2
ArcCAW66kRhn8wMjBMAzXWKCdRL8pItQ6sNBUJUp+XSnNlkL+mVF9z4MnYWLaxvO
XGVP2lRHGPX9QZrQedQrz3jSHJwuGz3Vi8oO6654Kjts1e+xRL/5cSDgPtUj0qck
ebi/puw4VIcXu7CCMmxVM2sknWdMKGmaFCEgNc0uokH45F7xKDJRGodSlnBtcLwE
KWDIBsIEE1UbneNcX0JZLJwnf70L1h0IoYLFMUKdUYaThX8sge9dd0A0mr8giXN9
wxAAsEiUEr299PXY62wEmthDkBc1gvUGBcOzWBV6o2x1FnyzZ5oWRl7c0QfqiwdR
WUZ2DFuN+mz6gwyJAMm5TQCqAZdhLMUg7UDYzF6GnFItus2EyeSek2wxi2P6Te8L
WicBnpGQVLc7DfxYdjVH2yc3RzOxa8HQOdPVoG+fnE5uAdMz06ha19V5DUAB1MEY
1ncGTeQfCloQjytX+4o+eIfZNieYi8FBT6c/o9ARWbItPSND5RgORoSNqOwHMmIS
ycZ0y7rLlP0BTkAHJIrAhgn5QdmYy68uyWbyL3l2NgeY9uR1/FQw0WWGWkQS1z5K
1qNewXRn7ddVJlT49G5y0JY+KiuBL12Ez8kWrz2Pv8fHHAjVCJftie8xhDdflZ1z
1rVPsY58EVgkmHLbg3TRbVcR3l9pNMeaScKKjUxOM9Rb7hn9GEv+8wIeRIqwXX+C
0AdRiWtP11KTQDZBecGcSiyIT2IGQfD7NdNc1Zk6yN4KLyPqdq2Xcq98Aw6SdE2Y
HHdZu82iW3rn8DNpSFtif/PB2rIAvUYlN/EQA4P7vJ1RrWRv0Zt4KuasgjIgNZGh
+2iCxbXSW5XvsZePyEWjNjog5RTkt9wxaaWbjycWts/y0jscy3Z3ChWkpk+AN3nX
xud/fcvo7GZA91ebb3nKeQDSWQrsmaRpxBFyU84YCxK2ydOT9Wx+Ji7VhB/haH6t
L8k7oA9bQId1slIf0IgWkq/jmcUDoWHcwEAkN70Qr6TliySAwTWABSAmVrnGWpgL
AUzOd3+7CvDkAIpQKfDbIx9dffWdDA3ggeTN3g7hSIZykhnEi2fp+EMAEXN8P0ts
Dfkc2OH5cOdlwpbaaxcD4hs8BFBuW/gYCz+85dih1WOdBQOB/+AWoU+LD+bTXUjf
MfgiEgyQrQT4E1lmKHePqeJMNmlRi1Jm8hyevXDfpim6I0ilCNeQq1UpChpHyfMf
bSfiZ6DQj3A6ZVbSeuzSLoC0bYUw5im63CpNzKo8Yd/3pZ8YlYd1o0oBkBgZRS7h
QAgZT2MOqx+nvlpyl7GM4KZY05vQHK7dUTdQn0B33bQkn0wWgLWXa+fJkncXr6Ov
tB/H7Ldya/UerlvVrVEaWQABKQBtjOM6VfYhPPQ9wxYIYveC3ivp3AlyvN7bxnoz
h/RfbyTuEwlnhVinYsnEOs6xZQVTRAhUfMxyi5HPDk1MIN33+t+cX1XW0yq/IAwV
fnMPYGCRPpoqO9SM4kNXtQTCtQuLhp/94+NNXWPO2mvxQP88U27sAh4J6cOjG7GU
CoQ2ASjCKMiQ3uEsfjHzcUOGMd4HIA1F0WYV54vRlB1D96tKc7w4SWgDkKNp5GHr
n4bKNOED/JWpY3mOpkOeOQ86pjNJO8lIZAjE+7smiKVGoazRHmA8JnQAPwZ2YpHb
1+EsC6VVaQSIeaaguv+8PsMtD4E58/rqKN7rbXE6ThMgb3c76qVjp2TRciI18tTF
3SKrFYUFxNLih/7AZI7FXMZldnR173Az62tIFVj2SM8DFlwv5lB8N6zq96aL2Avn
S2AV+8SuYvE0ZpPvbnz0Wu28OhRswYDQcY36aQSgVpn/Z513bnBxZ0jJ65BhppCU
GMmqJy6J/LADswLPwNW2SU8Asuu9G5VJWa2kHxDog2yd9cxjNAfxLf+8CzgCkvtL
xlPw/BDxZWbQ0Jrv4uwUMNmQ0max9cGcZHW7m85wYyTWobCxNBJSAcTdkBl7JKpe
6K2VSryEEE/6L8nldCdKfDRvSDhbCfbAt0NuyNe2Q562vJDzWDblQ7eloHjPPd1+
LFAEU7ZbBWmR92BJKYADCFwSgXBVC3vdwAR7aBbp4nw5Gr02VJsQR0iLkWn5yDCS
P4ikjE/JYfp+AH1/k6wNcRcPMiaZ69tyW233ORh7CsdCo2d7znqx+47HgMNCOcOC
FLEUWgbxNlibSoTyWwcVsOsXWEwlBWU697qjDzdEiAHc6PcvXz71rZu7bRAwnvxp
agE+kXtFroYCKfPzc20SBOEfWiLgn5ZikhE5t6US8+5NeoyubUjmx2Q5p1B/dwhE
r4v1ZIuUYVs33JMJGXlfvtEUIOAnqww/xEaD9PoHj/iIdKzcXNPVl89PNPNcBXaX
JbbSkwvfBcOc6YwZWmGMYCt7ZjetERqKOTeXnf23NL4R/Am1YbU+BwNNdU8I/c5Y
z2eRP10lvlhPrHdCP4ddMsudJI3VBGsxlA+pXM/rxvCkLOBpfuJTlB1+g0TzVVx7
ETXesh48pg9rdEhkrYRlIY5hkH1eZF4vmUnz2HHVGTof/otJ3E2s63/ol8PLkc4k
Xj6ehoX5Wrv7I28EZmM9LTJlVI0iuqNROghmQXORIw2iKSiXGQV4mnu33pG8OdIo
MoXzx7Qt780X0v54yp8yAAtDtFmZdi3nKjPhvvB4lSoJ8hVWtVRAZYtps4RMAJeg
xoEFnC6FYo1h34RmWPZLGvG3sAIER4T0OfeJrlCarM6Gb+audkUJTvs6frpt1kQO
7ahLqcsY5zKAw7gxvwC/9B3mbQ4btZPGImfH2IRcknWv1QhEWYyQD/zSECT57Tyv
Ua7nsMEB7smkHoEwPiKGyYlNi8KnxQ39DbItNk4eV0VmalKNqBkBIKgjWHx+D5sV
wQCpR/VAtheyzDlLSmK21P4KSFTO1BAq3Q1/ajlS7+77v/wfU1KKKWQ22ZaKP0Zf
aLLHu/205NCIijRrZx/0OnCmbN7bp4fo307eXgRz3qkWA0noANACC/LllPQjcEw1
SwDHZZPOEpf6McfXrnOCeI+AdU50F4IawbkmSbi4TujTCgKBF7miZvZ9UNx/hYs6
yQhbOjAGiOQiq38LOHboHsQEmSYL+AcVUll18plK3N1Zrz21m+DVzs64CZGLCK2G
UcaCxjr6EIOTpBA0IA07Bj6+YccG8FvUUZtxbrButWjGYpOecYOI/AdZqpaGlu12
NAIAES7Sgs57NXW9hbY2OTand1wFomUjJq2EBH+e5t4okCpzKLxEdvWmBGPKeD9w
eaYDlKxXyLjTmE7K/czBq2pj5Hh+VQwD93er1GU6cmwHvkZpTXV+9QOpivE86iEw
Cxqh9loDbMOoK7NDMFh3GnFg2/NieR76b7MFrik/qzqs2dqmIZrzs5ToI+4oIKip
7ckkVPG1hz15PA5GzVAxKTGmgyrLdCcMnusHIM9ZGSQEEIbWzj1EzJum8pVIrqpS
0MoJnlG/6LqX/oTTcViFJbHy/eEDLEEAsf9GdkAzW5ZeTZhGqwP6qMQXsoL42XBt
M/I3vB8bkG0CyEhJIEJmC+EeviV2TinG0ChpGvnEjhVdXIn7UvYspgU8AhqUIFM6
Z0mwqkhzEXMkP6rsrEKwzX2JIgntUjb2ZBlIVn/Qj/6LfVxU3uovkTLmmY8feDbw
A2zT3W+/Yzxmv73b3lV47q6MUX6fGVWu4a0sD/bO3j+NpmdWpzFsCPegDsOUQYVD
3QdQB/9YLiQcJALN7PbTM/CizM3mMliAnh8q7GdaqIkhuwlI9huTiz+sZyaUf3sG
SIRio16uq9h1S3m6CjdaYeY8L070iwcrm2/ZOCGWTVzv7gU8pT7LwIAbFZZXA4g8
UQv6sYlRnYOrOeaA/9FtwGwe5WSbdw/KpUvCiedrdXVWligVPGJGPgdKhW3j8U+i
9gejEZUltYla5PQquiLAso/BRzCIPaqUuS4FQVP9Rxtlk4OyzgzguUMFG+rdqsrl
1FNL2RkTqAZj2FXTRB9qb2xbdrYcSz1mCNuXIalPJI4/FcV5FmuNh/9LyyZJp55O
Fw+2rOiHMth+5ZN5AH86RUFFv6Fh/Re2Abozsz/EWpGQgMP9XWd3jY4ZXORhdeP7
zP3J8niFa/r4Arl7f+KhODT3rsJ0lo8bkDMekuaUTXGsCMN2wMmagsEGAeIRUWcu
8zvE8kLEwcDSuM0e6TLZbBXQ2ITzBUhH++Ie6fF8RmgpX5vcDtEMC3kBJNMmzAAw
Sl0S++JPpb1NirX8y60iP6ieD+LApa/dqDt4sT6h2pqvqB+vRS3aEz+yBrxFzg57
nG8UwQsP8IrwpV4Txo+B6FbzBbQsPXbJwNaabiain3hnerRMfHshgwNsJUW93fYo
sJDHc+BZ6rx/J3dTrfjGlHU9pnk1jRLjX8dAtCtYnL7PqfP++B0figQBGzK3ie4R
oeReK6YexcQHSxCtQmfuCybCWTMLQ9b5neQH+6SWf6/ag/59XNtzZjONLDSiNsCT
WfGtCPWh4VlTf8j/EyrHCe4DXMTDavXs4GJixL9GA/99v9VBxRUi/S6qSfCmCC0U
9Ti8jz+3x0I08otj7raXbq31LKbjFCUMprQe59LQL/V/HBcFK/Ppd73tSEQhiati
cI3qig2I1dRNUI/UMMAxraffOWc7bh8obgXwyr5U+tIqY18Nc4AICP++fzV7f/SM
DqgiCRFvKovRr5h045/GtsMsSfG8kn91zVdEg+cQSUU00p3K7DfVm3jNRyArbnsV
KJsSfYBEI4oL3wlJFbk2beEVmc494y86N3VFsSYwizk9oEVyGOLyQaY0PuX1leQB
ERcNgPUnjpvLF5Z+OLyKqF+DLTQeD42hosRxU6TfkbVNlsmnnkfO4TOkBwYnDgFr
nWwS+rRAVhdXepUIU0dPxR4D6As3QwcjCSUK6EjDnpb74DQSX+o7hRnAI7iK0PuJ
1+jB7W7sKXakaTd3I9l4nxLnMwpvGnEt+GnnNAu7+eyVPrC4EzJt+Jpvrn4Nseu3
DXafdDkvAoSqD4yw+EI/F/j7INGS6p+LiEecRpEcnqETqP7vOy5nYcC4a9R+Y9ZO
bkhenhaliOzR5hTPSdFmehNR1gmHGGFJilbyqVfKAXRsQwYb4i6VVpbP57GFaHMG
/lEzPnqs+sRk1SuZVuZpYRWcc/ZyvYdjlnyLDNx3twCHIEnYHGfTU/i7vYJRM8Zr
Sa744UhvInO4dumLrC0SYcAELZKfNAnKCO4wvjINPEvKJbfV/graX0UkTPdwNGQa
hmdp3bRDrGp6tln5opw6Nmr1+Owwx5mrPWVU3WJMsYsgEkdzcdw50DYqJQ+or837
90GX86n1Jukl8xq96xiLhFrqQ6qYpr/vJ7EhXAUQy+9NE/BDytW1I+t5kHpnQuDV
43mkGhbFlEoa98laTy84hC6J5dGymyyCwQs2sNeK9lXM5y+NoFqU6U8l+y+JHWml
+47Ev7ncJbasJ4nOcR7XinlTcKtOeBHUEB5WknOjIoaJARCBDzu0CMG24QcX8w9+
ShcpANHw3eu1zeaXnPVu3vfOkRNpYc2+bN5sdeFT7IDQu5HGRJ75ZRUVRifXKNtP
wVWs3LUF49w+S7Y6nGpmYsPe+gcFGKopDDl3suzlGX6n4HKFNnggRNdUtfyZ4vdw
PtV8RKnIqyiH8revvg+ewsY/lnPw3LdX+/zEaJC8E9+CZ7jk+9YIqaxZEAA01VmS
07etXJ0Bt78ltGw2GYR/KLtmGlyz9EI8vTlSoWP7A/HkCHI3GRlualkZJLfqb5PW
h6rFRa/zD8ygdcb6Jp+xVmsNXG7Bk9mXOZd4DUhd8v6lSVpXULU8q7F8Zoed/NGD
BE9e0gXY8wa1IWxXufP2UE337q5oyBo9ZVSIbUjq8CWH38OI9YOrLK9KUcnNAlQp
AcKJCRJOWFQVXeklZDfp3fBZNxxjA421nxH3exMfvD4futGxtFXck7/qB6nBBV3y
Q+LTRZ+I4xQ+PyNftPQcZWYzOvxBsiIaxvLwlOWTHFLHvFep78uJRDa+OnaDPya6
V2Jln5pcZuBe6T8vt0fP5gN1mA5OltxNE6pP3kXQG0qNLoItfE+4boS7plAeoW+o
UtgnGfqHkx+f/lW+2xREQ+1MfIYiXkafRcE7tYoQD2Q57qqwSJoZR5jETWq8ASUy
2egOWsZcn4nlhL7lZorkTMrVVGZPwEJ8RCdlN4NYDI1OzD5is4EUap1+yFduHWeQ
mzWC29iZeaBsp6WAaP0iiI3eUQGc+iGgt+V44yC4iy/JDMPyVn8dqKgJvEUb0aov
6KjnoC65CL3Tk2jHakbdzrWLMgBZTNeh5yB3XXJJ7qnC6O4Ai/G2pd2yMz/2D4J8
CjRomDly3AQJOmWxy1+CZWilU3ANLSGxudLqLw+jA5b/lZ/zf87pDWDZqgXLE5bd
V5J1UYvUFicXi3Mm6/hC+0TTydSWZkNXI5XROsBB4NiWy6EJWBPU3RSi9OfGwcGj
Yu9AISvD/8ZZFBw1ZvzST5sN0nj+AUuCT8KqrdwAV6kGBOUQV1ywfbwye1lleQK/
jyAmVd5IDveZk/eTfgiYG5ZMAJM9gRTJXKs4/6+RswEYvLdNigt2KF/NKZwbIfiw
qTIawGuJVwdsfz2VurfxqDg9/jKhOyfDxsUWveENHcCCbgJokK7Les0aB7mlBIjY
D0ifLIKZvKkX5SZxFc9VK/dDulzdNWjbwyDRlQM8u61nyuMz6PcFORzS/CAQIH+r
LhmwRt1kAYDwCmOPgVB+caiQILiO/aH99oI6ZvRNgmpn7PUZMM/MIzzSC+SiJWpQ
/9AENQlxLAgSiLdjR+8XO0q/+FRnRVNa28wPZ0ykvpbNmN0ZDO5Ku1dyOyz5QrL2
hiBPDkMyiTko9EFLtGnMFh3VGXMYUe/AdDWT7a73HKSUdZOxOwj+E2b99buQKx/j
uzTpVCYHGSztNIRNiuazPK4bu2ll9igqRjXcW5aEEI0xb64vvunfHCJ0UnPHUHpa
AmYYST97h3crkBu/4uY08rYwOSX0TRtkfuNYVh9KP/zE6WTHAmhk7rW57evuSHbT
z5/UTqjZisKJbdQHFE3STp2W9goyZszYa2ngeaRLISeSft5jwn2hZjjLAEVH/nfM
QuzCqSy4+adGc65UFQYurccl27M0TpcwjfC3+cgvnq3e3Rxrb4XBLT+wTfHPR5NU
cAcu2spTqBsmm3XKc4ef0eaNQ7KlNFVrWOrXzjyz1+lkouJbBOf3OUE+raYXBLvB
rjCZhmAhcfZubuVHoS5bZ4DrLKr6a2rFmyfILcGXjgLaLYTQslbp7K/e+bs+QLL9
ZL3W0117Zlt/yhylM7l2hw0s6if/KmVP69+qBfBehWPb5mdTEPvLNOdrLe9WncN9
l0EaTaf6BWFVCHHyRmTh/2BOcX594wMrtYlCGbLxQq9rjjzT8mvsM2efkSqdzbjn
IhWvXdUqLBrZB/rwfske2NmKOqeVrAqHp6MYt2/FP9IZ51SvLxMY9jICWaPTxRvP
f2rOLZq1kiDe1SK/qG6LfLpjVqRgd/jXLfkSOHh2cxM4hkI/H5Rr2pC/HCH+iWi4
J5GMWLNEh+Mtmpd4BMVcE9nF3Al4JpbADtxyC1xF3zo4J6XjpwUviKUwasSa1lLW
ljh12lP4xaJOvzk5XJ6r71sEGorxpzfGqXysp0QZOZXqlNO/pVq1joGlsTxVmLda
k4E5jYLlx/PmNNrHLg4k+WpJqu9b/DLbqLhgIzaRWjWn1m+6r0XcuANUvCwNbW8h
eRZkrveUVGGPajcRRkA86WA1nhb6shPtZGurGGRBskw+IQPHdKy2MEWNcWY613P+
Bn4B5CKD97x05p00KnPs/NUHny0eOtYdWky6qBuFFWQ8eBgk2chEA44YTV3gjsdh
Eez8Iw9PUmYRWNxKJSq3RGEUS1746D9Z6ylSSq+wvDM1gQn+pNrR6J/dSpWyQQUE
pFmffVBXQCqxgPCBDqEk5xQ7ax8ov/pENinlbJHmvRI4a3gpMHIg7347o8TldyBr
k1f9TpdgZU+DogLajoSy3vLMqzI43DWAudyudpNkdQv6fjESFLrQtTjXlp9BTwti
roX6wGLKBX77v/UG8lFfM8rQuap3jDoBvaAWrRmAKgDX1VDCXXaZ2QMybTq6ihgy
PM0Y8xB6ZOXGrmp2sSro9trWPIOisavpjEhDCu1j9lfZ2iJsFirjI1sdzMWAuUGS
wGxd9OjHubWgce11wiUg84UqgJcgcwSMj+Fp4SsHt/DUEz3xMMlj2hclJEKALO7W
qylrFCA9FwSwiNNzywSLCUly62fQIJx2f/6wTkOXR7IkJn6eAmAq3DhN5R+OirCJ
KRAauWYZ4QtsgKJsPOWR81GW5/6J9irvXQcsmWfGqBlbjEHUkE8KLN1AXfqgseRM
qcPRRBIrghACZEclAN2cU4/BPqRbcxB0J0Rpz67TSyTgewQvNuvdduCDIfF8+nN4
AbkibyJFv+QpGUbEMWEzsJ718b7C1qDn3hrDjmpx+ULqgoAjUp2kUlR8ruI3aaMK
qNydzocTqSU6BgdPe4N+RGQJOmKlhsmBwN7v5Wpm1ZGIs72gpKdNjHTVNMk4uyI7
D7HWhvG1XQPsLp/SuvlAGQueL4Z01fBhSokpcFMtvCEGYAqq36pziI7xYFn+YxkK
X7GGRADiZVcJD/9rh75ungjsCZWIvpPhdodct0dj/7r4C61nTDUlfOD0UWDghss+
zFBOGS7XA9Yk1IJ5+u8EleTweYKH9UpYPCrAzTOPae4OwOiceTGsj9poZkrmL+/X
E6aYw10QMqzT8dk3P/wMvwoV9muAGwjIEe966e9wmFF2uz0+akFLRu/JI8OaxgZR
2f6HiA51kTzCJDK0rA8HSpjreEHapZeVyed31VY0NfZrydit5m3D9OYKOQnrQOyB
nhVPf2sCipbCBypUZJWZHlFrEqoq41S6GFn6xEK48FXsnWnAbQLJxSDTL+e4N9vG
n6zaq5Tj08GCBi3pIIjqc3OwhQcNTJWUhSJ14wah6FQvk9houhn8PwkD/WyaTpe+
MYReMxmEyym41bs+Cv9DSEWXkKKf8NH0igaN6rXwE8PYS+J+JBobhM9cGiP4zFcL
wOauGVpgTkQuKQYqHJqAFEre4vBUh0EYTE8o1eAzKQ1iWpT7YwQr+1/wFhnK82hK
VTEJ+R0HkK+5FKXPTF3Ab+wauTL8vauvUc86v9IYTOqO/P5ioWdBVEAOJ4qNtxwc
XHiXSjr7FkyMd3gEzMjoZcFx0Ryaesiq7tl9FvSuE1vISfP3w+bSz3cTdmQk9Cv0
EhwjUspPgQNZ6T0Mu6f+s3bNmtWjR1SAn9l3SF1bSVQ8YgGW7L+aaguzAUBg0sZS
G8W0/xllt6zN1ykkCEBE0nLhlt4RaIiuLQlSllyb0HmV7IfjkesDDCCtTBAKIsaL
zZwGUkTC1gAF5bvqHB7i0lAq77bLpUzZtvzNEjM9Y2cyezKW2SwUCMHIfceQ8l8+
KsbWrR0KGEP/OFdFH2X+lQ60AkF7sb/skz+PpSy6CzFL0zegn/MJeYKZ26CoIYhQ
HaFU+H2Hp4CODiZ6jM+Dju7hVAC55saIBG0E5CyIS0bZD3lTqGmjuzT+aq0ocNKg
IP9AhQhPNayDvpg4az5GNNA5ywchX2wKh/YJBDOQFlrV7uBFcktW7wbUxH/IotY4
J1ON7GpBT1bNDkJLFbMjoxrIBqXj3jko0lXZytv8MmKmrpsY3foNzycaeUEP4sHz
3mudDCsVMsPuAvYCDyByDpSM0z6HPVg/BCdpNSZf/IHeU8MHWwrZJ1habfbNhCzh
5jCJHb3ino2Jp/Z8YrqMR3bKJzJC9lX5iC5Eab/h3K+/8gmkRKzsEvyADAiiapn8
vaP1fwjsPjzwqPnNjm+jW9KXxf3d7fh7xG/AuZuzVRHbvy/5/uw+8ziwiZB7nedG
r/foxlApxnalenH/JN7yxoLNuLF4Uz+4x/g1EOgLc8TC0oRNIVzIILrDCz279VDX
PUFroQVGxAPp81O7rre12Y3tJ95vKGDohG6Uodei21clC/vj4ehX57EyUPQFCKuh
dxU0T241baoJt5/5ppx341On5EDA+oRVQSmukFx7JaeqHewvyNbB45KPnxSl84Sq
tAx1aOJJs+E0LZzDWf31weV8tINjvckXqx54F0LkEKIqLYHy59jpwxmvLxgaO/dX
kJbbtGM3ME4FwCUrFjVYHmY2QeBv8hOogvw1RQ04FABJo5RZijhQaYGxHT4usbws
8jp2H581lb7eCofWf5dKOO1BlvIf5Q9MxWLBTvNzMyOA6B0jvuYfTYD4KykrZwIM
MsVljH0Ytt6QZG2qIgULtl2EeptV6aQYOU6JlRPOmqdeaT729GcMOmzw7hVGLIJX
0hMx4SqKNNMhs17a0bDorIGFRGTEIWkIcjMYoxwbs0CDXvZAfr6nk3EJjQw1YNzP
nsHSRUlmOPkdi/hIKfQ0wvzqy+5ViMqoyL2RF+BZzJE5oY7WOquJmzmwbZw/faeS
B1KaCtVqpytjpR2Ulz34Q7nAksmKDu4aiyO30g2O9aSdppU/3CdwsVo5RiDUb/cI
hchrVNL95DWByWIJVFe384RShQLrOXFwv2XfsouBvGO6SE/PEVXsK3ye+aaIQVD5
8sgVzn/iijiDTi4aP6jn40aBa3y4yRqUCBjDjazN7cPhIfrjsM2x6+fOqJy0MqJt
PNQ9675T+BsiwD9vETCaypWyXQ6NV1oZfv+FKSW5boDBQbAeEwgp1/x14rr+ThZp
7As3N4cs2gjl9u4s5XcuteavuhyAJ+XB4mYXi/7at2LHhI5OEh4xVKqRBc4fA2pl
FwLteNcmgNEPwjjCaLbzBh89C4QhCJld+rrY6w0xdQeHEiHFA9jTkEVb0+F/Encb
4uAEG5AHCBdFCifKbWLEagv4nkbqG17NSekC22H57Ik1EGnRMLlIOuGzKnhRdJnS
E/JSCxfxPCrguM2OD7bMtOZxZjRV3+U82uzEghXKSDZ/mjsvSeDCGnYiW4JfdDfx
Az+RM56/7S7iL/f/glEdoVPTsk4xoVyBEWxhYCUZKsdwWWWIuxpEpq+Sij+/vwRo
WCP0TSsn4oU373cFw4m+yHrixT8C/lmxnm7UR/MpzlpAvYCF4Vwxj+XTuIjHf54f
PP9/7iwUU2xPp4FwjCviGg+ShZwbC+QTAMaf5Jn4659ek28KykOG6EfFW5cOfglS
bMQ1fe5HDZhpYhWBnkK+PsMbZ7djmlTls4Rm8RVrTBgNxb/bTRYYImJ7ZjwRJMww
UQpoTYQsdQLg0veSrdgB/TmZrligIs0gE7ry6VTKCKZCA56HXE0W+Bidr3pst8FF
HJdTlwDyxKyDgRxjvk9HWpFTZWHZTVqkIhovkpT8u0gsxFzCCVWx7pmyKumvZFQ6
BjplGdUOzgYM+3n4q5eeJHRtKUDtuM7aIH7OWIhIFa+Dx9tf9um6mkqBj9Zs6D0V
BVeeBb/9duhIVaIgmY33SfeamypBk/t9ARNxxcvZhGGprG/lLIX7C0Gzmn97n2Yr
71Hv8b7G4r6tQ8v3P6gZY+G2SIibekxV9vBWbBGNAEiuImWEbYCbfFe9goyZp2sR
R5H1vVfrucE4KfzCaX6BUKTYc+6OWMRCTcK1g0qJcAVVwXCo4Jzj7pbyKAPzdOHp
8XCo6xWToRZNjcTBfW4Sw+HumJHGgccAXppt3DpBzy/WTxF/Vn83QhrqEcmXuwVQ
sPu/HmP2lEf2Pp8fZTetroZy1mDqb8RBGAJKnqp4iOes7XjIsUYYYr9ZFccmmaiS
v9WidJbiDwB4d5ZqXMh0Hf6mw7owobkoU3yG+JdzKiPHIHcj9cMol1mTrIR49WoF
Bk1M6rWeAM7VDcPuLwMYtkXNhesQMYd2j43ucfRyuSo6I0+siQ2ITrVgp6liE5oW
KHBMOJp/D2JG1yXv64oN9cTFDxepQqCF35XUCiBpZ1BKwT4t4wQ3Y5iS2cosu8sW
xCtGdU/mxYlebPLH4DBBylDrcBX824iD3VrVuR2XaRxk5Dgv1zha2eJIUCjkw+cq
MAOC4IhsyIBpnIBiNN2pScsF9a5KMHW4pDYoA7lPr3S/nEtSYdPkPSm4loy4mYgW
L+VnevIU+G456cGyZ5qiZOTVc1At9N+++uSCDUVqQjNcG0NaeJzpVlONX2kkVjfy
FV4WQ2jxToPzJvzos4M73Lv/OyQp35u57dR0PA3OTy9UHuBhEwzwZrf3qAbGcPpT
tmumEk2Fzwi2Y6eXc5dsWD6Zex5frTVMKo5A7W9Iqp6/hCJ+GpwrwVow4wscqvk+
KvQZ/bGx/wmqN4bjSo9Y9T5aItzg1IbYknCMrcYxoZzMkfOTDsTxgwXQz1TPYx/e
/7Vori+IO/JdRlIXjoYw9taFNokGWkI2+iRgO6NheuYo47gLDHh11omnmMk2FgPs
CLoWnnnU8BHeVctdExJhCk65vYB1gcYRgrfPzOKjV5ySiKSQVBWRqix3h8BFdtz6
Mni0VXSFAx0hO7VU7rvEGOrT4QvhWVTGaXCtuWl3es3f7bGzmDd9nyrMkkDe3ixi
SK7b+VWvhn/9QwAUopR+EeZxLSGKZorkOO0bpQVeMyJXMDOmy6l9Aj5I8buV9puC
yh7kDD6HnayU2eynbRtEKnxKYmTFaR1OwTtG2owr4ZPIgi3mUtpB+lhG+xlvgIls
SLxu7kRQKGAg9NR9+NiP5CLW9CuSvsB82yMQVqYAddo+woNTjdC9L/3KrKnlXDxz
RrnmMnId1xgLI1x9pF4gxE9CLnuIGFiWmx8OKBkz0klSYEqwgBN6MccVf2u+t1Ni
dN6RWLsiRRO1PntqEnJnHQ+C8L2tnaz92HVEhzOsDrmWZEi0eL9i8WN64QeeFY45
+UAH8mgdoUHfnpj5gcrpki//KufRiNStRE60AHqjrcwD3k40MmNvOdFm4LPkRbvb
dHVUcYfKB9771nG1kMZBLbA2Qnbm3SpPI46FchvbOySG+ZRZIGZYiCZoEOPfGm7e
ZqIfZ51YX4zE5ws4D2j4lUVm+MDwLs7YeQVDX05YdbM1LpkFR/xil7TRP9EPEUtA
SUHSTLk0BgmmOILWFc3N6tMzLRT4o4ysaIIsVjLS7wyuXkqMUCCkaedXmB6hKb5Q
v2Lka1eg1yU+3JmN8ZBj8a+XJBRyh1X/tHCKD2254Q0HDFlI2oqAkAN2Z6w40vJ8
+4RPcrxyXfA0m6Yao8EJvNJ5TTJEp7HQa7MksfY9yI5DK02cTnNlvJoruBmZa0gB
4KlLD2cK41wVGCht47PoIivZqpVo8Z+GPyJqee4XQNZC2nhudIYmAv89ippKl+9c
BgPOzK6IRqyYTalDlHVFQBPCQTQgMBWBMIJnn97aG1JbnySz/JlRVRlopGR87AuD
ZOMrn48KtrklMCRQIqvB3XYFdWDgwkUTllWoIkX2TNnxVR0cgyB2eao5g10K8a2I
zShBQRnkVr8wvP2oaTJdPX7HmA53wFXe7d2Uzg7jCjQUEeGDY9sLWQncBWvXqOJF
Ie/MuHwAJp8o5WaDK0hZ8j6tWYFMxNQHPhx37ticKwziLgcJ0JQ8od/9yGAtjq2x
Q6nFfNL7Rx6ncx22CXLHS8q6jbIgH0iMy9aOw8F7Jpw97n7ZXD8aC9DydgihfPJs
9o8QofeKn0vopPkXq6UwGbO9VRmUx3/97hco55bmDj6UmDkMwOMeGGiRqtkejGeG
cQPJu/sB+HuND+L0j0JNR0mrT4mzZo3nhyTcE0yWUFj6AZ6sIgKiXB4dgFm7/B/l
qETORWjXfsxAjyXNWyz+0ItayOZncnbRfSgUlchwq0rDckp8/alFt7DoLoniCQh/
ZWMQ0Nr91Ujavysar34W2W+P5ABxO6pVebuAgtHlfXX72TgBscPs6Ygi4dOB17oy
d+eAOfIGFR82X3S+/5b8b3nzqa8nq78LrD8lR2tdU2SGEIdSfLqzgyD5O5Z9bDMy
Ajqwr/J3pP637MONSeRlhzQPEy7WkuRmmqFTaLBLvOPMsUvDBRuLcSxq9vq5VLHJ
8QfPTi+digMSVEDf/LqoXNwiYbtjBVQZqCCubV9lqwG74afhyhtLkBN444gAfCgI
jZTsdAQTcpmrzven6qfMyn6oDtOR6MDF+NmrayOn9Gf8noLztOVVNTia7Bs+o0M3
BqEaiXtKtjigH7AMXmBFBs7StVf341q1gm+BR7FaYRFbN5zoK6q7GSVHsvaDL9PT
tLkhWDjhrjK1aJ66WC2IFRVxc4KvCmCDfDJzc1+NmzRCcsmPl1oyMmDOZdmNjOUm
pUVs8XviyrjnfwUywFPENcMWfPb2sBZ1/zakkfTodconu/twjlN41RqmkmD5Vdig
AmtRktw4lHVxN9hRvCm1CZZxOWmF3Kr+cXHGRYkCyDc7EuTlug8o0aio/LF21zD4
qkgNmaXaexLgXMORzpsOOEtrgJUCsTm8cCk9vnPp8WBEH40Q+Upgs38Nwe9uFkIG
GWalgzbw965PQZntXkHhCoVKXxpAglpo/dO0THT/cj+j4NdZnaznT+tT+h7bPhjT
dIYeIA0uaJuKz+PSkjaMNxd7LisYcPVMRiYLOQstW01X/Oq3irccBgHNJO+gs0qs
JGY+IAzT38sl0NOszsGnjCoTRafDIwORbTfKivNMLyMkqsXES2pxcm/46P0IvGEY
n8YxRK21yRc2xeGLAP5yvJ1+hRn9R3zHmTEuR2+01kA//FgoxLtwPpHBTI+5z15R
T6uMnSSkf8kj/aGoA0L/ucf4hj11M9ZSqJAuHUA3sEg4CSFHC1hdp8ma1IrpFS2T
Mg8vyistI62oou5o13eT/V/ZPd9qLBlJZbF8MBvOrv1EKNYzFBts2CpHmv3X/BD0
J4vAhNaysRvfqppOEsCQtIUTuhfTTzmHoKHUnHm59DwarVX17L0m4xtR9g03Lyyf
bAkwr7DFa7vDyphpon9X2pmJ6bm82kNHqi67KffYzmWavwfKA6lrjp8cpe52VNfP
lUrLIIZbst0/VgHXWm9v7pTPWtbTjUpCLXYlMojiQgMaFAOS8mulnm7atMxFw3PR
k/rSym8Y+5o+wKtbiIAWdzSTfPGygQeLYIw07mAhXbEGvUQ0fA7ihkxzcGeEtZB8
aYEWILcCAy/bVNyXc049ECJXONfgV3A97+DRlgoFfJGyNqH7pxwXix1OIf9OIA0b
6K9s4zi1YfDu3GueJ7qR3i8Ayoka91+biyKdzGvUv2sSO1NdR1b49MDB8D6wGG5S
njbWKTAoPAqwNxSnQ9f7315TEd3NTrIPFVgqIWOG/p3BNssnCLgF3OeO8o8Hnjct
F3F50hMiBVr+P1WsZmmMOfPEyS0QGkHb1u+cgwitszHkE3em/FoAQdPHKmPYHXSK
O4lF3qivFOrff6te6tGRyPsi7sCyLAROMuT7MwNosKVHa44Oxaam/wCOSEMSMB14
4UIYzNXCrCkisHTlhzThrtvoian8exeljvBNESzzFIourjLMyGOUyYTAiu63NjAD
d3E+wxCMfsfhAjyAfopR69jMxQ6G3wzysJUcBVVZbbLly4bo4BriluDtCpwisvOA
kYQRoQxlvXDG9B0WxO1DsYwcz/d+/396jOzFmANm7RMmwnWdHNMRcham9p+JIFdw
yDQ0dd9WQrcebkhsCWYuaSF9pzyoDxUX7V3wwoDFaF8V5nPxVM7Y7BgT5G3Y74BG
MIn6wkkpoXP6M9wQSgEevN49OLCscfdXGaGzASexnh3XyUKxAmfLYx1c/Dycbg5t
RNWhQ9FzyGmMdEquAzvd/6p36J6PAjYQIgFaY4r/XBmL+YIs/aWFaULpd9LeVzKx
iQirDiBbU38yEt/y2D2o4X7zTeXNARZTA9kLx/Mjj2A7QM1qhWJegTltSIN13GrO
2Z6Qfhjk6uXh9fSN4tH1U+Sb7JPEvh2sqLFV9+6frcS8F1htkzwTXlw8Sbao1GyW
o7782l0Q2PAuO9Tnh00lu6fX5VOYGn/PqSHgJa/KTGIeaDvvk98isxIitrCq5/KV
owsGjyM/tQKFTuoQfR3642zy+yOLHy7xguUNvqVQ3hn3z+K0CE+HiVWfayRjm/sk
empujrFy+/MT9w0naH94n1CgauuugJat1rj0/Io7V4nq1kAZWAPH5g0s4G1swhFf
09kDIut4aBXCoog6bYa2DIK97Ut+U0c6ozwvm+JyMU0oU9QfS3c2cgCXOKwAxEP8
OwTpkr851qrpXoQxw2e8RxTPS8E56WHDtTo7YVZ0IQm6qM/c35ZA7rBbUt6rF9K/
kDSjj0WEj7pAflpWWSoyb09TrXPs3WnuyzqDkK6FD7nqeXePVS4QoKkdwx9Ic2ze
8JCHAJ+DmynGUPKOkccaXjBUws3iIZ2s2K4NFY9Nh3uYZhucOHIaRi7eGOIcRNDG
`protect END_PROTECTED
