`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kNqMn2MrmczM2dW3kWZKcUlsbLwGdQocRlpm6dvQ7tstLMhAhWjl/Bm6jmw8/4tg
qovetQltxIKrykq2bIGo7WBWpAn/QcSOhYvKR2qp/SDOmBWrqY5Nqj6knn9/tEDN
NHdzV4Mz7cw0H4+4T7VcjzDsFrqLsuCIImOBaOQ2/v3+OWwLS3DOnjzMfRQ5KZMg
YSZwM6MhL+YDk51/eoIa9U/2XvlTOGwclRzT61YOgz/yv29zEXlaORzhy62ZnRYL
O4WPGUgDToKWJkm1nhRlRPljC/MHvCqiRI8uXua2CkHbR5HGH8lEyReMOfekvmCi
eVACuKZb4KhEcq45mpjsR7qywGci9+evHkdhk4gPX7ujJb6SBnTsnK2IxCsH+lpn
Xrbdkr/90wGz2t7Z2oJfj9CtfelcL7503fP+B/ulzuXR/X1LoTLquPl8yBUvtaRo
`protect END_PROTECTED
