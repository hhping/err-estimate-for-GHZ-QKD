`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n7kf6zwL/6gLYeVIMpdmNFQ6iBRWPthKALS8b1bCMN+wHB8vZPpnpz9w5T4WZk7k
5oQQmvKob0vDauIhdhDywjGHCwbZoN3cYTyMNo1+R1pxwuSC/V9Yx5A463AzpTz4
WelW9MkU5AJAmAowh5sD7F/CSjfV2wjnQQvfPI6d5X3yilN3tOPrdt+Wkyp/emch
/qq2CINi8EPlbkbypfHMFkTF1L9OuAB1NgcQGoeUq5O031tHTZJhwltZHItUxSLW
FLPAu0me6BN02XESUu4mzzDsYTd1r7wtjdCNZ0V63VoFeY1w2R6ekc5ptu4dIQ7B
r69+CM5SUdK0+wZ7I4EPJNGbcN1942zGwSRFRXwOdmAyrFKixz5QO68gqLKVTG0U
Q8LYMXKeYAaua0iNo48Ux8Dn1gT+j7ti5jvJV3/xLNaH6x8LtFzRBCUmfZNAxJSj
m81DodYdd8kNk6fZvq9N0JvlZKdMGlrs6QwfaWrqLRIbi4vfw+v2dQhQnZejt64i
`protect END_PROTECTED
