`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t4sYT70UY0eQpfSmLDZBJ0DEZ/rbMTJQHStaE0p3y2kox/qeDU+AS2ZL3LNbPVSG
WKXAVX384VOJIAxrHLkV5WOT5JrYUW4Uj8hVcEy7lE3w0sW7fbVXaVUPzdtPSgeC
CXSLncI0Ad1J3cmMZLY9ZMicVd+FFMUAooDFf6rv9S6Nv25APASUYXtaWHqbyZq2
7UN6dgCJNPL3nMS0A1EgACJt+R4VIOG8SIkCZAm+9AX88loAvoly5K39/oDT0xc9
HDEdB6pJ6HERmTAS0X9OBe9B1un8rA3nveXLCn3/y/nDcKhBMQVV11MujMSJdT5a
Kko/onjqLXLGuolakblfb+hAbJdArTBhr4Hnm8/ZAqDJFvZPmSTYTOCsSrDzpZbl
NKWcG2XdHQlhYakYxYCTOv917zDsxGYx84PjGYIhtlnQ8YFfDw3bEGXEc2fjSj9O
+6By2hezEhSCujVBqd9E73ydsUcgTnIvxXSOzMWNatM=
`protect END_PROTECTED
