`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EpDFgBVuTB1RBSQKRWMa8B19o+8TGaJw8ybQicnu9IGE6IOoIYDpVmUYmkTpYIB+
+cv6lriIJ5biUkGyQjgHHtxPyb3DbFtvBxYum+DfStUll68jDMg+O2Qqqj+yAXVg
MhQeYcsGssqkNrQsuz8keCzknkw7uWShuPUzAQewVMUP2X+WclBymgFpQmxtJUWQ
BsI5fnrZPV86en5R3iZKHjByhWL8rtMeRQ3QX0dBodRfa9+InQbIIbaB8A2xhJ+6
0Zy+gqp/CI4RSvO+1iV61JhL7WUo/mo16mRAQzlf6KIWSqldiy5Wr6zUiAYdA6Eb
TASJUjja9Ucbysd1OvayU18U7wbfhnDXGhjaXJog/S1KgfOD1DkxP5rW9aKIn+H5
EuLuVn56o5gN9JJ3kN2GOFug24NN/f2wsUyeoIVCBaRvvmf4sjufleh6LgfzK1Ph
hBYRbeiS/70J+RkaOroov4bN8wV+JcbLvQxzzLy+ZPXYIa335ZlSiieCg5RNz0tr
QI5OolTGQ23q5e1jCOQAZhnYF3Ox1ibfsWcvTtip7lguA6jgZCfMtISb4oG2b4W7
7AwPpR62mz/jpMjV4f2TvwSD+aYkiF4MgSwmc/XZ2eS5Xjv71s8FNpw9j+GmefUm
PXxnVPKRhfTDn1CYqP64bCxPUXQ6ZBiQniILbWj5hVsMIem+rCKcd3tMW4uKHacO
`protect END_PROTECTED
