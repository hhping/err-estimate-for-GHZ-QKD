`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gBHKGuHnwhjJvIW3gmyEF1KWHa8NRb0kjSSITpb3CjKDtUIT1dD8ldXR1b25UWu8
VEBIh8ZNAQsrvCjNgtkAbpoUriD+UZGjz+gBqOyQqJ7OEthoiKrDXCIMZxIBGHau
0wlE6IxFpWBOL9HZqdfH01t6cq8xaDPkkUzhOIdL13dCnfGjXv30xZoxUw1g+BNB
fe3jVZ25H6pZJ+ZxsHO6o23Bm6Nb09Cv3NpVDZnroKmNxx0NDXmEezpFvLInu97H
jOUARROEBXMtnX8vXYYoaLZZEKk04/j0VdFzy/S8e+d0jyN+B2M8akcLNPsOd3Zf
zgZqqcgywW7GAOz+U5ydr59MZWvSwDkYDP3bXJv0plmTDSpz6yG7t9boUlt8HBTU
5V1TxdhH1Q9GM3EslICUGfg5ncxAh+fe53OaVQjdMBupjinda3xszAGyHCpXvjty
rzFM48DFGLuL+60MlKPmLRLaCGKhAR9vhImWHWkcHvvdLTYRlRZRB0v0rMBUyDJ6
NbTNxKtOMP3CCN4yBDe/tZ0iPrNwJLhfPVkGHbW5V3ezrK3tnXtoxfzPXblR0mNr
2FDdvU0dZ6tX4sW1KjwQyGSB51+m4ekIk2aDrSF89G8IhGFlMwQny/jQYa5yEbig
x0D292kKMbd1Ips2yYj96MJOQOWVvqq7avT4n+0VWcxfWpWmiScQRVORaiLagVTT
kbKMMoQEmWL8BZJNTuFwIzFnIW+Sl+UHkmY53UgwUCp/oS6rc40m86d8oCspsTfP
PvwSUB1sw95RER/Pez/rj828QJz++8wuN364sIC0iSy7Zngxw06+P4sZmLr5eqDv
wWVWCtKxHs+amWVue1zHJFMqXbhF/WChzbVuaLvi5OkYa7OrjdH+wSI4GmaLFC1x
7tEV+UBQzRzTJVPfig639ecNPsKNnBoDseyZ7e4EY4a23YILYyfluovKDwU/nmdR
TmfGUBEJDBQiqkunahMrYGlCg5INt+HA0Q4q9asi9ZHpzx6Pt6/2/pt7eqnGv7yL
+yEb2IZorwhqBuJntRZtzfTqp1HhA2UdfTNd7RFm4wv7HVUU2HrjoAdlFvcQiV9t
aX56U9anareMaVJrt57CTt49A2Gvl5ZDk58JP634aEr9ogACTOJvGJO10a723RPT
2Cs5xiMAkUT11xpm9XuHvfiTQTclV5os1Seij2tfNc663M2lobu44Lq7n1QGztKc
RZ1iee5PCudx0w8Un6EkGvPk+gM/6aRBwl8qzxnGXoGWIgRCr6mX0aso4gAHwtGM
GaA0/WE/6EjhlXJaIfiKEQY4JRFOMPyTCeu8naWmYpmuI/up/r0jYPeB/crD4hdO
r2T9YfIbwMZgw2KmUrmtoEh2sJ6ZalDgrT2nN6MoU0lpBMJRoZfpxYDMFBLqEpWu
8S7YkHcXv4bJjdzhzN7ngysQPIhKn7ihxPnNh9czr4SWOpVWmph2VtCsTuYd2bC1
97FoIqZFOdsIwqkvs/Ry+OYSWvFgBqxL9qP1xHwEPhiCmEQ9WQvUgo3/Tq45dl8s
/2Iy5SDf4fgDqtOQPVPxVLNKBxl3c8T1UnwR/9HUfbQTKFPCGMB5bcuRbZh0Jc1t
QMF0wupOUFcF7gn694CgPrxfH29qCJk7tSXy3BFr5/off+m6GtWbDACKh2HgQFWH
5EJQyOB15PpgXWVpqjB26Ii+x0Bv9k8Kcg+b7wkzPJJ387oCyVYepsl/5r5SzVC3
YopPNCO++uxdKID8w+rp+ZtjtLpZwCsPRBgeDuKxy6OMq25QJe4xU8pEGnsn4ysq
YvwqCD/J3MCAnQ8uAg9vlDXJNZDublgwtrf20ISXKoSTwzOKjuLALRFFOHbVxjsp
a6AkwEGADmqg40rx6OL9y4It7x9xrJe3gK4/VAeWOSpISnWKbvObmpDdPrpCxWJi
rUNOt8KTlh6UDYkvNayxfM1mEJzzHGyIenajsga3kfCyel+DNtyPhOuQKSTMG/US
/OLJra5tyvRCMGnN/hZQbnq/MBxrnMJ1ZbZZvtc/gQe379mT/uvK47Nn36X+SBEx
oa/v+nKwQ/5PiTUH0Sbbid6WyMHJBseE7g8qlWL5QcSx0nC0J3D18p7YZ0vX2cls
1PrmJXqgqWP1+Z7ypL/AhEOOrH5EPm1wfTmcUzFCEJtLh+1eevfNnAxKzImVl5aS
2JkSVPKaQhfpYxArO3gE1YEm7HiA1UhszCbv5M6J5eLTTIR7RZU718kg45eWuJ5K
LMzrWX+EfcSae6+8A6GJ1fO7cNSSuZOroyelRdwVDsKjpRuSwpl09biQPQfiEnSC
QzzUTzgsGyChCyrcJzDa8ukdNH8hnVdWI/cerAz+Mb2TsrRQEItTDa9JLTqAZyNa
RXjiCKPb/voCCOtEEfVK6tiFanvmuc8fim1wOM4u/c15hFlkSUhoVYko/HOZ3qi5
q6KZbcq+9A19qa8rGmvMTQJ6C9bsGVsDdfLHRyeVzdy0PSKR65IKKoC0ZFij4uxw
KyT9DnKYVll9w5j9qy9SLKehNQ+FJ9c0aJPAdJ7wGWYEMSGmlvAIs2RKrWZjLoIB
m9T9kZjsgLgHtIGYSrBDf33lMAC5AKlWwsfIkmwpXut6/XIx7fdmgjSQTej/JUE1
bS2A0MOo8+hH6vlOis7wJg3Zh+Xq9fkqMmkSo5f3k4cSC6/LSnLMGnoQSFi7Iib/
cvJdZ8W6f+7DVjqipZcyhtP/BWyJjhChjeF0/qkiDdWPmc0+WOz7pTSQR3W9w17b
FYNU2UsN3bLILWxTPdNk07ezHZ6JlwAOaHlS0K+ls9TcWT4+dKjAGvfyGX01IAbx
qyh+ro71w4nFVlOTce8w7h+fdjtOXiIDXccQ4VmndyIeaM+i/yh/rEzWEtxzW7E1
FQh37GZSR8kkYpwyhOFanPj5InWajsUW3AhlF5zBCqQJxrhhoM8/PYAw4VNhYs5o
NN0M3oFcA+cUs/ig/qvxJfFlmAMvijWslY23wYoegWOM9IZRIjwTY4/WPCp0kg94
HmQOxKri9BwJWGdKBeqvSZEhLlhgYlD3XTfGklDbAaHCL+QSvh7Sv7a1hnuWu0SG
0lkhqzQnUwW9MGW+EXCGR6aZRjEoEA6REsweyMJrGhG6uhXAPJvFA6ZmXh0aObmd
8Yyjn2jDIc233hcpEFWU8piZGjFht8TOOQdzOWuMGRmpFBybqNnD0fKh/x9qn0dX
P1CR6zYqNlqGmlJ+eKJhrs+x6AbwHPjB9jMXaXqfDG995JiCnH742GuPXi36555h
HEhxt08ejWdLA9WDJ4/z4+nVYDw4wrKGBdLkgAe6yw8xcLZMWByt6YKYlBhiE88W
dlh0NpCEW1ERBlTvGb5nPLP7D5KQmGvU39Qto9fv2diQ5XYGSCQ0n/wCeJlMRi75
tujTbqajRtn7vUMjZjWmyb4D2dOfqFL0CK285O7g6QjpQeuvtDECFM3A+qHAOqGq
TZubQ7/GlP0Vjxxro9nIAJcKWvQffdEyxFHHx++4nhAjdSSKowiWsQthmF6vROjW
F2jCUy0Fz57UCfk0nrIkqIsU4WPgCQW00v6zSIPU1bw2jOHywQDrX/5gk713rx/t
hF0DoLX6RbpBFydnVl993P3qej3REHOE63dghSGZYzrk10CJQ562d7tEjseSbzhX
/daffnDcqdlaX21WPDmrLFYn7eibLX6CGZcxImHSjx8sC1KoKF8S3wNpsNtAGOzB
7i0zPjwxgmCRvX6+VeEex3TZpwUfPpsVicsbZGWIXkbS7JsugWxR2hW+R0NC6qGy
HhOZxs2VkwY6V+UnQ1xtbp+h2huSIJVu4PGC1Jhf98MemxhIkxuffQIVXpJAsRmD
+6UM6Gs8OAXe7NnLLOOBLrTKesIdEyTM8dso/XjlpVhS0LpLlfEvlkZkijtqyC8h
URhHwlwn3vONxlsEQXMfda5j8Wpc7WBzWu7iykuZd5lr6o2Zg+3ZS+iMCJzDKEyI
gnsnQIt0XGPw1H+BsYDuSZbBzmLbK39ZZlCOpZ4pSOK23AOT3DQ0V09GLfjU1A5x
ljvXggCsHjxedeGAbUDBImpyhEnF3UPehYqXpAldiydhUp0RVGuw6HxEMpi744r2
bWgFFlSw2apxEhYVf5ZM8MsipVLSY5jujDVo5THwM0mFBQmD+Kds6wx92H/shull
cgLANHEr1iH64JhbQdtONgz9DK7UcYiPFQlqZrs+MFlGg813phC0yQqvNdCPSLRG
EKX6TktIXTRVD/b52LkL2ROY9vVActWETE2s7jbRMTTNT5W57DQQXCA+g9DUfxBe
P24gT2QIDh8mwQFyZTLq1HNkjoSU5nz3rjOD3Hg1oyBhoSH+y0q6Rna83TmwkBa0
LsAyvBdeTbNZzXapDq227wHaeUCw6vSmt6mQ89wM3NkTuN5rmYqJLNzEEp8bH0/G
hRYQfiGtiooMXrzobe9Ln8YnMi8eHlWslI+6nrH/vFCaTQAcAx9bZfpHlv4Shd71
8HaBevTF1EsYiidwjbcbW0Cubv1y4ejwJsMbA+xzYllAcFGCY8gCfHMC151q9Lpk
WiRtNkXBcmpXLaABwhajIFdfniA5o3CLR/wj4ThA8YLdciJpDClCxUALMohBf110
Yb338vbQdTUW1WWJ0PyXuweUYPzkODsGYw8D3ar4Tk3+Ljfys/HBvfa52LnKSQhr
qWfcgAdNGt4XyGjV5PbTgfbJr+W9HoKv1OC0oj5Rr4hO14gZyahtOqjFeSdY2QCl
xmi+FUHJAGSaohO+m3yGQ/bZq82hjrwilCydG1YSVpoyFhy1CSSbZ8P6k4/8FmlU
csDJ3yOQCjkxiohJu29usBJndWv3m2yX9hUzBM0iXrn2pzP2fizsy1ocIP92K/Q0
ompP1mp/k7lwE8wL4AI+yq/bO+GwTNi9H2BknqhUEpweMrnro35fXS3m9saxS3J+
gr85RlGKXuf7oGQ2OoJCBgmyrmZy2RHW/4Gdx2Te3M1W/NlOJzD7GdmFeJZiVjZu
O8XmaGFgk85Q9fUqE16mhaY5SDFMnqptlwXVCrRHwZNDoRlhPA3bjrRha0USfe2d
XyGwGcJLsjU00L6rQ26tZ+kxxXpiwcZ1gaJsTa2d+JXGasrgwfslfZNGRUcl9Hpz
S111OuZGfaRQnLQFB/EyC0Nn6OH4mdz/YUEWcost+0ljMj/DfyCoFi0oyMC7D3HK
VXbhbJh7PoURBrq5wrjnQAbGti29SWkqTbRzzNCLFEkPPHE+XLBkzfUig0AZncmB
FGnxHIm36ueCeIDe6sAZAPM9Gwv4pIJPya/gWIZue4v5EgbDkbcIPF9d4699q3e7
YWxThIPohb1G1CCcahhmOpyysKdcSteVjeXtccf7Pc1Kh/QnznbpfJuoJmycjAuL
p7CzkYJn8Upu36Mpwk2r9h0DVe9Ah4PtQ6NnE2Ldhxj8l24E2qeirOkSK6hGQr5H
nlaiEwuF9rd6JeKflSeGfmnN908bNq2MVK2MUQ8kjU0tyZO/I44AbXmCyyWpa+SU
uTCHh0fiYY5sb0UjjRJ840b81rjfWub9u8JrTG1UOdCn0enN2Gz/vGiDnrZ/7Scc
bErc/X0VxcAzQpvoTXy/0AETYA/FFKzN5wyjdA/tqAZF3yOJ9bq7jcB6gMv/E0xg
yPDg0EObiHNbDQ+YCWQswp/omUBbiiCEoNnL9tU9/LX22LxTlDcNvYhzcSC7gtb9
kIgZFf0Ys1HzqOtk1qN6LGnTPLiujP5mYrj4WF+daL5IKb5soIBrijrHua1wEPfl
tXMjOm8SdTRTOnS/zB9QiITNsDc31HvqopKnhILbgtaDfWmt8d/8rUPXwvo/SaiR
J1g6nwMQYAw7EZTxdQpoQ/FTepYbGvMLB0wU1hwUa+KgZoaSSE7qW3QJg65Yx9rY
qb6UpGsSjOaZEWbmRl1dxY63ikBBCRUm7ue2rRcNLd8AC+wymouxrM+c/RT/UgyJ
mx8gspF0z4AyJxFlJVQ29wzQQUsAlSgF5xQEODaLxU7UxIcSxlTBCWzBa70kcABi
zMjsJP8d2UKEQ0cpvOm7OI20BwI+w3mSeWlrmxtYeZTL54ANVM0VgTsSFPBb+/zR
O97lSdFzN+H3H/6AjQ1mMCBOt11BOzJz43HGOkuxn8WZpS3FqMt3xw9jU3CZlvkv
GiNleaE5CCskju24cX7lwhBGMxMSPSCCHNmUunZeJj6buLZKpzMzVw2Z+13bDMFH
mDvLbyvEUpe6soQ3EupMg2skBTjOG056MzAIXViGeEU7E1WvA6xPwsghCSOncfoo
eNNmlHKsl3QXOCzwuG1ken3vTarWDuqbKJe7+/3jvMU52kN5b+LuuOWoHtBECAeV
Ui/bBcXyrO8HtSvKsxHYyMWAVqFAhVjrOcecwkirm3vPjs6aecRRKd81QyEh/nZ+
NfjmUruZSAEkyrNaYgLoz03BPO62083XIEXaH4nkOfAE0LdYupdDSbNjU6zRx46X
JKoaNAwpQEGNyjjXLcxsDq8+NkSJaoa1kPzHbE5h2t4N37HXlSrBKFSqE/bVR4ux
PfuiMWB09eM9lcd6GQlNjaxgdjQSaMX+crqATVN09m9aG2t5oQf+8IsjzK5iFHnI
KdGig6dsI2zlk0Y3uhCnT4ak3Q8qOh1g55pwBFtKI8nZzrdXvChwFcpcgzkQz5Vo
wE1/1f3Uw15FxfWjoj699ISuxo3YWZcUcVzC4lEviqCxeoOsyUanBtuFA5eTdPCU
NK69b6RI1IgecK0qkPatCvWI1+ESng2qk7h7T8ABQ55lwHc274OUugA98mIqh4mm
MjFcRqb346eNOmoxrPn1n6FcHnNE3d308nJBdGv/6N1uQ3rXuj+xgS9FKo4RskJj
2uvRKkS5CIEPJZRVvLaHdsPOCLXfhnZ4uSnabSj0ljU84rehx4nzW+jIuOLHonpZ
KLYidlGx9cy92HcIdZ7ItqrQMyVmgHhlAEM8soSIQRr/5ibKzvBUaJJI0ueqn0zA
TfQw4DKQYllY8Z1iDC9UKahDPlmmj+ETx1shKnz7NA9gwzXBl1b4VpH8w51SFkPm
C/f8aS8ldYb3kb6mkTDgTITagjXR9H0qTOLu8D22oJ+xTxryfS5cooJPriI7USkv
OYVI4dyaNmuDFg2M3uFtoUbDlevuEkIJhrlS8l+jPHxAhFkSrC5b5poJBBGfLyQR
VGq0NwTZNbztHulX9C8SQ03k7beCC0ddYAyaGwOoO/AlnIuYI1m88Cnvz/yR9ATR
E8YwKlRj5m2xZXD3d57CbLSxTJRJhmMpirou0eSMEepnPFgGCc8jz7fmWMAe4hwn
FCHJtOt90lC43KosedLUMRSALFz8PFicKkrHaeKOFlecukivpKbl4OZeNBUGt3Jo
hvD/ExP+/SQfFttht+3e/Wopo9NyqcR0S7ldR4t6SH1H3uhhjvRmPYV+HL0CPKQE
+vlRrjMmIpmt5msvhbEE9TjKEAVZiwn2xllLPfymkWGYNhPswNPL+5QnVaSQ6+FS
ocs5u53dfASy87/J3cQ/9nrbNlKvjdCBumvEis4Ch38eQegt1vki+3xAllOU2uG+
FUanz4O3frB/Gup+91MchBKbkFCH/36RDjx845kmt9NspbmQ9s0TY9RwyF/uE034
1s+HKR4NtGtn1cAzl8AisigSEKz+xZFyDD3LBFjdtKkVYIYi7kbDf4jIyqRbSCVp
GByNee42+/HBHLrLJlKx8w1S3CcAHjQfsX5W61BT3+C5uo1RlrOv/EsbWikFU8Sf
qgG09wHZlEMXkJP4woP9nYSkNgptjvT3MW6yYBMNxeSfnf45gkNGMYLlPLsaYU8J
CuTG95XEPGQcJKHZ+JQdxFm+4wYlPDj8ZcdAy+XlkUELT4cjgbZ59It8OQO8zGpg
U43SvOJVWLrvw+B9vBFZ8jslbiK2dFE/IfR+s3KrRtMwiRPQhOOFF22xwKLi2/nP
d0Yav+x4CYoNcKP8Nvu6HekL16Xh0qVjZUtqnpMIjew0STOH1TJbyqZMhlSgOf8u
7e8WBB/2nuAvCToa4mEeDYwrHlV9LXyb42uDyHL+Oey9xpM0KREfLoXmU/rDco6q
v5yagvGouDJQHQn3Y+S7U+1cg+tQjw2gSFp1l9aD7sxYmLKynDnOR+48T3sGPBGS
wvyR/2kyZMQyapaVyaMiSiV/5VyzfUVnUq+8jMIobVNfEya82cKz3GX//1exnDOE
Y8AimZ/ta9u3dvDq6NNGvG+q6O+MDFiLIPNnev8pqUu1739n2eQTwOBcUstGSJ3c
cOnJOLvSes/ezeE6hi0eSASthRLLiNthYKaHEL4Bx6XtkaTt/05gOeYa0PAn8WKA
Bk+pXpmH2ulLapHZYTnU67BVaz0qYXh5C1CIYTPdk5W97w0eGjfQdlH6395CiX9A
OwCzArIXQh3P7oDftlDnubBJR8PSsXSFNj3Y9Q1G8K8BdRT3uCztzm5SUeeLhih9
CTC0aKn0xqFDSu0NkLTh07ytxf8LivPjoWpdRQ4DLUM+XmjNIB/FqYGtgkOIrMYK
xXhWK7KDNFXLUv+SWzpldBoJAPaSQ8kqsGWkgSPFr9FG5odGVibrBbxYwGt8Llc/
BkCuMunjejcwNcyMn2mHH83kA9nQAmtZJQmi8QLjdzmOumakV/YyJnBnnxgMlMwW
IdzKEgYeKCocZVunmFfFJOdFj+0UeOz1glSRM2XgEbH0af7Gqftl8tnsyEVjHP8g
xBmfEhb1p9tn5WQ0gjgP/sy01EjAAzAY2X/W6GFJigBz4r2QtXwsqe2Vphe3v5WA
TWtszczo3X9QOdeYfe2/Eesq3gz+nasJn2q/qD6LN1gIHv6+c8MBuGi0zOfm2tOC
kFGkFEEUQsjaGFmKE5jTyIn5l5ZjFfvkZn6M8oaFcEQdn/mCQdPmTM5kgturASJB
7IIwyXY/Nm/U3G+aPdP7by6CrDzQqzw+rPFVG3n56wwHgIt2evoN3nQ8aI564S4F
yxUAEbQCJmoZV1RENaXKOtbnVbZmKcLpDxWmgcbHxinNofF8lSM+MkrqIVJHOydb
P660m/YVCvSFfh916C3anZVBheGCYsEV87LPrSeRODUHu91gwTEk4Me7EcfU77d4
Hmp2BDDJoCwk71d8lmF1ttipjZjvftsjFdru1QoVvyJ34LSW5pihFkoB4MXFIfKc
zR50fhQRne7zlMOR6LaK2lyh0u21tosTe0aSzzA2QBkrvz7We2mNVNMaUDivLflU
9SXv0ImnkDU7Q7F6bRe6AT2Iy3DWjr55VbqkmdXiDtowzHOp7gFvXdCQWguHikni
tTx7OkW1dXX/H5HZpgfl4NKPCqkQw9WAsD5a759Duf0ZvQcOZr1b0C9cbs1y9Qkc
FexHsfJ5lQbSyRLdMxdfL5LS+fzKiAf+w3oXkyCdWjHEcLnYnda9X9In4XifBTVw
VceQF8Plh07bgKrrfJ9dmyZ0G+iNT3nnKzQ3dTw3XZdFlju/AnOm9OqAKqg3szDi
B+/gp3bcNRAYN/AOJFyNyA2stWt6GJWKGumuUt3mFZUlBbzSkSpSgnJkPVa8td5p
Wp7UcChXtvBsJceJ+vZydQqqnX/NmPNPlp2rdFtz6pchpk72vd4l+svb4E4uH+N2
Yy3Xm8qEai9A2VjUHRwNLFyQ9JS1tu05AhLqnmv+VwqJkZcAqQ1OyLZL4nn0CKrP
/beewIsRMhQ4z5GMa4xdl7b0jCAp9Y2wl3rurB8iTqHdigkTJzQcOahwjXVVs8Sk
5tvw570hAVThFYfCDBYCN12W9eooc3GOipxd0SZEZksUR99bXv1l+2xg2ym+dams
jtBLybgR1KXnSAQUd1v4ZSx4vnFy2HnGxC7y/eYsFd92fivmSe7z6dt10RV8l6Hx
uKW1sLfLf2ocAvschn9F9kuW9eoQnJIdPULTvaGviV3xFEQFy5Uydz7nddZqGa3J
H/ZpcjitFp4sOfxIVz6LiGolcIn3eySpCW6JUOiqOWwGwQMQ6Xb0e9y6+CQD96Pj
UJNEApsAhbYL7pnX8t98LvncIHgqOlnUCSWuO8NfEiFhJVgUakJxfSArktEynH+i
aqPiOlnxOg2PsXBhWBOeo0PM3goPw5/9U/SaJLeMrPQs1L8q0o97bLF3tEx1vXA0
Zkhkuj5nbmx/BCz5Ms9dBCisW/SWbtOmq5oPDhrSWh1FU+eDWjSQRCZhRZeJBEwc
txizsoAuldysLpm8A9N7pfFldYiYDKoj3zeXoYWGe2j9q1cEmKbUp5VOulE74gVp
VLl7vYsyhpPw/xhaclGJNb6BAJ2H2zXi+tF07PYd/z3Cw+5wu2ialCW+k5C2vYwF
aZXcpOoGm4IgssXmSQO9VFInltzVyVo8oZPckuFlu7S57Lxs5kygncOwbdrWfu1f
P8UYUW5UqpGYxKARzCB0s1LsNGIoLluvofVidI0xKZdZLxquUo0UZ97n2CauENXu
pVG6GdNRNN6lW3re4OyiLkrv9ejfmW0hSwimyfvj/UMYIrssayrk0jlp12rFexqT
QiVah3hqx49mn2KMWoq3gki6qM+99DLHFNpBJE5OOa5WNZQw1JguzXoydxKEGFZA
uDtfSUPWq/sXEcIUzKUoqwtTxZVtj2U+R9pcL5yGr+HzXp3HGMUdOj1GAUOiRXV6
xBf68Ghcm1mMViwU/++WyeXnh9W1Zzz0IViz4gUa3oMpGZsPSr5Fjqv268Gd8qku
lfRCbS5YOzMwHjzZjc7BNpclx7CNVjbOQWBPMhlNMGVcBrabDUOtmqZx/g5+euVK
FxFd6yNUFgnPYw/BCaTWF0AY8NsK9a5KDign2a1KzrcaUAVTCJYAydxWQP8pogqr
HuzfKaB+zoABj5GRY210JQ49UudIYdp5y/FDPmCkGoMs8tOy+LKEFJynxmNmEGcE
XXu5VC5196LSLbHLqKpvm6LidVqUvWY4JA1s/9sf39v4nIkf3c276xJRvMFW2xkD
9qrKljyiK2lYuiqgNOx7QeEg7d04z0jbcKVVkTZ7Io94Pod2pY/1EvWOBwRJxuVg
RCmMXz5PbGo9XxsfHo3uC3Ds94apTVp5AZOsuHKMdMixMjgAOZFi7dQoyaSDndyY
cLwIsF2NfNxWQV32nIvWIiZ8hZYRhAhSbjTXnIdNVbBz8J1tkccU03FC9H7+38As
epOFScEe3KhtR+9ckdCP0BtABbq0UEI6pGcyuN34vj0kRixXBHC7zC+YhgmUI/SB
qMs9Z3Echw1Dl7EC/x9EjyAOeY7wMQ78FRcG/E/ji62gran4riajlSmPv4zzZk+D
nEDT+v/CmblpEQdix+eRXLIqcNT7SU29HkyjvMIRdvIPEa4rMPIKWF9nAOMCK8FM
Rl+4b6Qf875topg8Zj52Sfax3vjBj+On3QQezQc86bBsYxBswKqdLeoBZPmDTTrY
lueyYkHsqRQutwISdDlLQOsI/LGsKUpVEgytMZgBP8OTdOREfwv9jJfHmu4aovkb
45kQelkYZIvFckRy/CoUC/FqRxSfNakOKJkfz1/o0hxMofY6MnZbNmJzmymsZdmc
d43eAK0GNDbiJcDmMq6weCkE/XTUxY92G7poYQLF+bXOo7xlL5XOGecjPH2DxVH7
QTFPq/7Ei8AYaNiidNjq39S8PZsHgX5k65C1YVyIRaaq1iVptB0mqhlJvqerZDc3
rUUe/2eoXBmYx4B5QeM61/14Zcpz1DOC6Bzoxze2o6ohX+7C822p/A0/0EOK3LBW
Ib156fZ2BVFCZRVwSFIFq1+p1KToizcgCbmc68F6GPNRqECyHPUfmYh2PsnH/Z/u
ULF254mWXdlphyQV/dv5T5X9ZamjE6JOJYmRGXrYdqILnSfQk5n0mJUAZb2vWYgD
TdlhBz/xU/0XaA9sCEvNEmccvBDkMTImV3N/QIKUIHaAiG6oDNBRamUqrhmQqMJw
+9QQfPgo1XxoUn3gThchYlryz2x82edaPbW7clLlcfz9ZIidfQw7WT7wNCY/uGIv
B6tvug7ThI0kVFxbiR39oxY48dC8m9q7q9kDnw1QcurTanl80XkDbJ+slRj4WbU7
wbkSn6TUG4zKL/FfpV2vPhrSfk3kDlCwx5xU+ragrjQRkmfUXvLF6pRKQiO1dZue
IQ8P3o3IUKMGQ9fSKDM/Hxnou76FDdtz5RU5dTdHo+9wEQffuWwG6NtyIpFgl8rL
Gkqhj2RBS0hmkuBvZZD550txLcR51KGYJKMcDxCHpGAC1/8BXarMTsxQf2e+PFBq
c3Vt8Cp9KHmznRmIrPLLEBkzyUxsmVvGNwbYHPft/piQ93wX+jrz6euHSofYwvTo
pbe4FyDXMJSASLqIiLFnsjPXNkLeUIgx/W69e6KlINma5nz4QdG0vB0dHeeKTK6k
m6phKl4rPsKlPvVu5QcUyRndR2JuoFRtc49YYeZAti9Cn69aC8nkcz+PN6q8+lil
ZDLGAF9gdBlcon2rHHutucj0FA/gDgGxYo7JfsyoeTFEk8wyaoO6+3m1gFMbld0R
QFxsAU68weBqF738BqAnVzD75BgqiKXt1iS5LHEBLUb8iDKIZPr2zjKnhLOm0suC
QfAPbHHao2SBjzQN9RgDIoEIYSah2eXPeLrr5iYR+fB1OxVdFY2zajJ8TYk/H49u
WWxcnYJbKHa7zIADMmSuXuu1au3v++EzHBu/T48dcV7+XwPsXIm9Das3TTG2OaEv
7PhqMnYVj6jQCZZ/MnQtZ5Rdml+tyWBtEq3ULrr5/aN9b7wc8g0h4NrUP7OF4KcO
jcF7eyUOEeCREaLLrXCvWNtflzizqEWjPdLp7QvAlsgYtQoerA0IZboTtaIDAkT9
T0NumJkDlr02X0eLBHdQBMsYReHEQVMuoerRQz1ouRf250YA5x3qZegDnY5ii1V2
a7yTKMHvzj3P5CQKaoge1Bkd2SM52y44klXqpiwmLvXUReUV5CNG3CCkdO9Y7dWm
JfFzA/P98Q/hF1h2tmo0MrXEl9zq1nDB+j9Notw1ORiAE02+S7LxDCnFWyG3dTdI
+FkUxAyndwp4JWgO81QGzchDmlqvuYqZKUxawySahd3AI0JGDtjp0BRXxqCjyGDF
0+b1cZu+nlGbvBXwphJ2bTIh3cqFg96UH6WIgS6ADNxh7FpxTO+rwAzwb8DnI+wu
OWCE2NznAK32AxXXfSdP5HTtXDQeMX6WwsEALWb36wxB5sOYCXWKwdKFhJ20flPb
SuoSsRobj0DNaKRLVl+tDJDXK3RRXZP2DCt89V8Mo7iErETbFCxVfSwRrn060Ixm
KpqNtxC14F8GnoBfn7DKrK0eTSMdqK/p3chogzXksq6zstEDdHT4hROrH2ehtluA
nvbkAhjUIgctb0d0QSNHmEwyqwEJmB2N9mJ5apsJN2TY3YP5/c5AKaI3t7wYzQTH
gSmDVB6jaCE/CWriinMP/xy3MVWl01+rIvOchjLy52nS94uBxbfpPFjfWO3ebt+D
Tsj0S/0hGdodH3lUN2y4AHkDk64XG37TGcCcl/RaCINbAU+SHJgjNdkHD0JqGP2I
Y+PqCtX0DZpUHZv1RPEsr3CzXs81FHEURTqdqcMhetsiXDpNOahIYhU2Z7gm7SV4
7DKtjD0UcHj0oXFnypwXTa6Lu6BKrzfl+jXPFyYMHZMnlL6IBzb/a7C3SbluKyjA
xvJ3V9Kx5dV3o8R7MwQPqChHpcnbfAYOpfL1Hka9B/rm119k0C+bYgLvWJxL3vun
Ebmt/h9MW1AY6xlqENAIvfQRbCnKxlmWSl6QBJ95uNkFKGkQheuIcQy+G7XKYkQ6
CkbYk+9X/EqdtIfFPoXxhnMtK3ihiPgxu7U4XEwXZxYZ1gpza2QoV/cQfKujmk7c
DTtvVWb3SxQ40/PWmnK4pHhHjBfcBR89OKkb+1VRGRSNRfmSmg0OA3XFed0Vt5JR
eLDU9a9EERs/FB0XnplfDQEWtgxtLjauSHGTsx+crRP31443Ql9rdgRYllLetCWd
GaInMHL6Nt+9vEqo+3hHHmMOt1kpS/3rWlpVJYwR79vKv5DFVAQfjex4fDGbiLI4
XE7XzI6ERBwG7SZe8sObA/KPvw2JTP2HIP7HawlZRKXZ7wez377bPFrzKjGKEVBc
/keqsKWo615VgcbVb/8jCuv2BsW3KWp9rKRe+exxwDPQEyU6hV2DdD70hxLwssv2
Ht5/zLpTGAbc5kE/5GMZTncObf2l5oguRq2sPOmtvRV7nnt4NTd/5YNsnZuCatOM
CGzQJXYVGMG9r4hNBSYoLF0Bp4rSZ8AsybjaIMq3y8VSsem/k7OWOJEBN2qdg+IZ
EKKIRxOOO2j02/zKIyiP87SFOwv7cK5eaYEugJ+fkfQQQiMyVY1i5GUwBb/VJXtY
zY7VXo6zIJaxMv28kwRrM4PpdKqHll6VqcIbKIg1XUoI14liupfxvlbHoliKVbK8
3yLCYKg163XEAKAc421dQ0i9UXakmtcaccskF0/C7U7iYSHITZ1SpvHduHg/2wzB
XTTbdnbIvnhWSE3ShzbMo2ZS/yjJYxH2Z0z+xP74wWDWJERYGSKuYU9bwvi6TAf2
OJf5hMKCYEvNfkI/7B0lO90HJAFrr0RVkh4p+AwrfI13K9vGjUo8qh1XrmPgTYVv
JRtUdtSel/DNFDfww6g+jp+fNL38aHwJFVZ09BljxrIPHwR9gwMDc6dAIojJ2W9s
iaa1sjehO7GbCWPqi/C2Xxqdi+oQAcR3vwUCIMBolBRvYYAgaioj+1Zl4rUn+zVV
5ng0wMgnnaS6XWhn8H/FmTXQizlWpOAqhC6LyYzWkT0hzSrEBrb8nNVF6agh8/05
re/hOcRwcZorqhXZ61ONLTH5wO0mzV+HP48HLQTlLiA6+VhXbDttsRYlYECfDgKg
FwJtDc/OYNJ9da8WKcsf5mMm+wXiz7xoxXsH+Wbp3j0dWUjbBLqlE72tJ9PcpoRw
r+0c0aqNHYGxFd8JzBvmISQJlTg2wiHKWs6wEepwzZ4L5Pzt2YuFUjDURMIbytVl
cxJcE8aT56S54/SvkeldY24G9IS07s0lIXVfrqB2TGJqbKbaTgX4ta4I/DWpNpHn
9ExoxP8cTQHxXJxfEkmVsOcZArIhKxvmaw19vlzbMHSQkx1hrsILUDeHP3kOtNqc
YtXXrtoZHeseSGHOlzIBo1CmFIMBMpSfA2q0zdUeTR+c3l3klN6F0ZxaFnvIe+U2
il816Mx/46otKV/s6TN0dtI204XMMNGRpsfWT2S/0cXfcmqfmlDbBvx5cj87ONrb
JlnjtlOdy+YSIcfuhxmL/AvIOvFBcsy5GbDJq7oWjMF+CDxBkRu2DvrVqecXXSBC
9SNvDozucyJFdGcTS6a/y5tIENor6jlD91zu1xKbx2MHCYc+/6zEL48ZVptqju25
qEjSbIzfAsnYI+/AxRjDbg3KgiOKGN9smTtdyDOwCUrCE8mTFn/b2L+jIBlk6NUP
gduwB9JeUyYRu2w70Ie6x7Y9m/EDpzmrbJ4QT9L3ADIgpmmiz34YFsSDtsJWF9CS
A8nDLwmasYR+e6ZBnym+Ejxs3zA+P+B1spo2r0qNqKwKnXfBs5ZUns6rQ2pTjKLM
8V1ODRb0t352vrphXjsUC1lTFvVW6p6Wvl35CeMg/ai62riK7VUJ932qnPCoHjHr
m3alBc+wLljU7yXp213J7wN2jWcqZOvUfgYBdGxPPb8IDosGuqgB4fVDtiVRBwxs
4BX6JUM7fR6C9CjaJ8RN6aND891GhgA+t/jFKQIHzaGYxUaCb2/EDpmiiWhxqD7r
Zbkp7AxydJRSgPpB88Mr+iPXBD8nomhOnDIis5NeLmGCODT04EazA5Atrco0DHUK
P8HvoixlKYVOiQxoA2p2vfNg9tBpg1dEJ8y2UjPpywj1RYGczRXZ2WJzrxbtvsB7
uFHb84gOnk0DwMtk76WDgcTYZwTNkJr4My+c8kc93wVtc11wpSK9GDKu5qi1+3gT
WAsAV5CBUxZmPUHpxP/QZcOGzQco3apse/GCxl9R1ryQv6MR4tzJfgjmUjtLbEf5
GyILRYhsYPi9vleJecMzwpprr0B28t9xCBxH5/z2hkvtqESt0KIqdwn0FqK6bW9d
N9WLfdl5Mn/pdTsT38rQwH46QcPmG9MFbu885CK2hvRadzC2rxs7xQKg3AVdYb6A
sO0A8OQuR3g0w1CqOWDMcLZqucL4TEphCJd6FBFpuwiidpJ2BidTFK23DMY8xjap
6Lm03Cme/gkKqTP8DBWPeG/qxqht8xoNc/rc4k+aVLH0Xdy2tamzlyVEerFH3c2i
oJWzzbhZ3wkR/UX0X7CvVLtickuZJN+5pBCOBe0c8JB/oYvQwDzdpiaSNesTKeD2
Fd/Q2x0GrTH9aQEA7mNFyiJV14SO6s9oElpDQCxk7kjm90vPj12sV5lmnrY94WIe
FbmD/kJXrOy2u4DjgwjGMhgPAKZ0Lb+ZyyK33a3DagoEwo6mFrJN28nk/8PfoV0K
Sf5CmjuakAQrdBOCUOAuSHN0+qSTmInlts9FZMpw6RNsS7r9z3lE8+T1h4lSKbo0
+i76nt1jp9it7jh2xJuFLohbCCXqiaqkLO7GmemjGv/9DmEPVMfuAnfj2xXsGemk
kpTrt0xtHnPuFC5f1yhhewBtyrRZNc8n7ujXo2OeEk4FWnLea1CRUcKPCMx8+SmF
g1n+8vDdaTGuTEgkjSYDV7B8CCNn9JiouPXf6IqecULRNx3LKfGcfrdBh8EKKF+t
yXYTw8aNjjWnyaMVBdTa47GAI+fU0CjUEWBcm2/wqmTfjicJa0zdWMTpAFlUtAub
jY3bVOJ1bJezUvMY1mzXCeecS/safZNQwAg9JbFCJiNGXc43SNFpbtDldYlK0Gw5
TGJaiBxvjNxtQzL4FyYVe3qTBzimzkJBddWbGf+Le6lyY1UKeM8ZkG8Txpxo3q0K
pl1Zz4SmjriFVgvNkNT8NrfVO7UUPiTg0FVlj/jEK7wE9jWHGsPMHgxzRquVrdwB
pVwGcYgznvkL+WHwMbNMgtOxk0ABicBktM1LriDzL1RmEzu9d0ki5eagATZOxKP0
DgPFrdSiImGweKg6Quo1Ay7BzBXVo2ZEJwiT3lRqH+zLEodrosq+3hfv5O6iYLpB
fikbyiPEPsk86dbdoKnuKlobzvpFPrdNzjaWjF0JlvXky8wvJjLKH5Ra1NMnpjri
/aDemP57suEesrFKesA7xSHwX0w8pgCeQGj6Lm8hmAoOr6Dq+/0Ywj24ZNBVR7id
2s2vGxCVKFVi8/hJoyNXUwOM2hx/RmMcf+uV5a4snlxcidw50LpJg9JRYJnyhx87
ua+/3YPn0YCMvRxgPK00jydLqx0C6enNl7BDv3XYZgugTRDZ47KTrFoD6O3FTRTA
I94d34HOBk3tppFD7fwemc16QMd/l7hhdSMcGEWw3pXOP/wHAYJZDKrOphCPWmA5
4OdwhjpGl0gQlGShLY8ISsA5+q9iIRclt/FaJW+Eeyl3WzswEGrYcDWKjN+Y7FxW
vPZ4hvbtpU8/M3BtgqQDOdFNac+l/2g3Ec20t+O30jYjZBzc98Dfn7W33iIooNhk
hFYvcmcfox9z++fOc5kQyGo346pognhx2RiNf10DgtcDqtuupBb4VaMaocu/1oqu
0+AhjCgM1RodCyV4diqdQWE+phHJeNGiImA8Xi3/HMWiLRVeJzR0NcpIF3SWbUUk
Y9OkQqa7hTAT6i0AjlqyVdCP3sEOpV4ysjCvKNzT9JIhd18TnjgLPZHiZ4syseUp
S9OuWduZEMjBklKBiwcrzhQ8t5CKD1tLxBnkWnEm/wr9rv2Hcy2be6uI07Yx+8Rn
f//oJJFSZwPF57xv79xqkG8JA1eqaIx4c3ccrgQXxHMlgRPmxO8AxgTiHm4fSVkr
XRwbnlc0Th4DdjxTYAsI2Mb/VqtqT128vgTM8mz+3EI1ydYykUUhrg5HBFQmXPm6
eMrIYAi5Jr33LSBPpcK51rFtDz5RizLoOVJAstFyRSJKx/Z1+Jq1tDkhTWGLmJy+
tAKa20ZaU6tUpPG+dUWFCdoXXrF4jHCEA5pPihy3ztmnfOhOFTxewYC7S2oAFXjE
MLRy4lXzZeTZu1LSyoRZAGYAVwzHW9gnUYDi1kjDUst+N9CsooVS/+/c/hDQQONG
PIFpn5Hr4KmdxL3Mxg6TkAg2lbVrcHtkA95skW/XWTA672ohaag5Z/zxbyAPICOQ
uY7bebfL4F/HMjkvYMTdY0h++tq+7RwvjIzUT+sn/f9ouYbdYLQQBxLe0nSDOLVJ
wMbe9PKm/QhhGDkfEBYwHJVJUatgMUWJgdW5UtDqJZR4Fkw4kAiXczGQ3ulH73Je
CkBly49JNmpFX8V806Yjojbcc28+PJ9ppLTP/BwPsvlydoQzJgmFEqMvvb0RaMW6
wae+XhfflWC87nTAzlrGJRsUKlv4RL6Sg0STL/Y4wLS2FEFkoqDH1VojcSOS6c/1
m0NJLcm6saL1z/rV7eB1+7LViR3OIBD+0vYX22WukwatA65Gw1go3tRyxFV4rcEx
TdaabsEoKD6CkpJmBXt9Yhf7fAbeYDekSRwUuC2kaSp94DOyPb+XvNJJGFtIwY/W
LqbjR00kRvwGHT7SJj3Ju57kw+0zSO5Z3Upu2uvS29luPgMJjEPZE8/URRDBtcYK
r5nV5R357ZOloukFu/iwArzYGMcBhbcs16dZUCrqnM4AJhfWKkEDFNn7GfoQDjfX
kAVaBbD/nx+1+xp8KIqiWjVBwGh6BVYWQf6gcpmY0ud1IL6cOx6bJVtbtgI3nZpl
dMER73IOJaLnjw+Ajj1pmB54E+8uSnDq0cMmjmXdr1Z1rHV9MGjOn6r30cLm7WW5
+QSmBdyHUoiiYKO4QATJpYt4IZLFvWWV1wWcKUBHm6ok92k0dHIPI1wa8wqY7M1S
HE5tQG/PVW1sEWsCYVLNQ2wrW+B/O2OsPxa76Bow0z6zAbv/6oauv2YjTtErVOWO
9zA2XVmCwSQDy9GwAkFRjWL5EfFZpbtxTVxiCeL6SzIHiOOjiaWHtyGN1NqjXJEg
EACQQHYvUPBoZm8HSmm62+HXxJt3Yohhnu4xbSLVgQo/g7hL+7sRpif/RRAMY/dI
36h28+k8sVT2KsmItYWap355dwceE3HY2gOhCVC46cHNGdnURmz4zxwRoymegzth
a8NMpopAOXBcIVAY8HydXhjKZ/eXJxOKO4yd5WSKp0Jiu+tNU5xaxjmC/jcBNUrJ
j0GotK84n0uFL0iOLXIzMtfO+k+qXnUbl/aN8dJHhxdsoxFstr8deE+/ml2tnwf0
Xtjw9eUiUf4i9PvDPH7CKpJvaWZ/g9rqE6BVoU7qHFmk4ED2kI8mqnjy6KtyEW6+
Afxn3M95WdDhqjNbtfFxPGi3thmm9fIRuMyvYKnMhoy8Eujm+cCJi93Vw4LBCjjc
nV7LQoCJsOMLqBU5IZs9B7wE+j9xklUF8gjGSD2mtGtbJi5q66mpIrp+nGQCGaJT
dY8cDx8r+BJ294o5nN4mQKQ+Xn+1KMhRLprDwyJnOk0DyMbNcnNmsmBFXh3XUBml
IlhLtDPZHhrYR/yNTCopTjp2QJ++qgN40oiLV9mM7/1F01Zu8YFpXTBrh91VB3d2
E/afCS2+R/+yaKaEqgg37KI8dS7Ks3J5HT6Cuv67MvbJahnCoDe2KeT43FR1+qTg
iXrAgRHN+eOMazKpsPGrYCCyidBno2N38BTyiDNzlbJ31YM2cA+2JsLAkermr16A
K4Pje0jIjKRJBeLqFXxmL4PCSMhk3dUK+W4riAEMGywbC9h9LfafEGYNdo7TS6o5
FnCVvYfIdy1bopq8k+ZbjA7Vlfd+7O19mLqgPeUC9znautD/ltlyb6jPTl4uhoRf
8NjHSBqsNLK8iHMtmT8RIOiVctrDGVqD8LAfLXC0TsnR0BtaijvqCZsxTm8ETusa
lQswuRLwExnZUYc1ehsL60brpY4YDrttRHUExOf6kOjpU6S4IPYajGVitjBQWCxT
/U/UteqoAZ5BKLJ7PEWgoKFBnRU65++nlKc0VAopaI2r+5LrQbgur/WONyIs7j2I
JNZAw/SkHgEQPEf3kuMgxDYzd2CSZgHbKidWPaMs6fdfmv5/tDi0Vm1172mKuFOQ
JTOpAVUKYeT3igyhapmb+XwufIT4Fv15XTGonsxGl8CDCCd4RPy8jEQnFTz7ndsx
A7D+3e0ZXpOO7MvKTS7OAPsb4XULVPluDrqVrmyRbf5kcumiCMl+KgLSJhmpH5zK
22envCGEdRuQOH9gzM3arrOucxpgIzMMYcVSCLedddOhXqdpPpW3WaC+cXB9fXjl
IlxKuqpI0wRePBCE7q+zTlzcxYOoUeddKXfzjoWevAvhinQiJhIzwRUQGuTCZU8/
ZTRj6VeWbulXELL6xAp2jUy8+S5nyoATj9mH33EzKUaz2IPMSI68CAHjDpfgmpC/
aoeuZ/n4M74J6q40FiCHKIO25ddUdLt/zjKtkd1pmmpn3e6hMka2fT5NlYPaQUlj
/02updJzg+dNhda6UWMEdg0S3T6oguGhFXuW9Y09duJviYIs9lSLtYOZLRoKolj/
c6Tcak12dOR53zdl590nYeja3s/34lXHMpGMTx6If0bQ5IoUpsDgjJNpJVh1Hbd3
ifWvLImQlhm1uCVgwcpwt8vn6os1TAOsllRPT+xiQspDoLEStPYK1895WLhINXjA
dVB5Jekn8VBRKs3hgKfNmsKR57gvieXI5XEYJBlw9RyWbqg/8mpfuJW2+UaNnGHa
MExWQrstLvYJjFPK44yT8/TtSZykvKvsQKeQyzonA2+unPdcBNu5wN8lU7atu8zJ
ss/px6XxR5VxneLj04nBJyRID/lpqG6rcbmqiGjWe6lCSMjmaMDmTKZAGn0zs0gD
52pYiglpk+1eJMpT3l2sAFT0YfrM+BkrcKZN2NZlIbMzGPbd7bB4N5r2+LP7sqWr
8usut0oMy5AHepdwyZ4JVGOvv4e6bhS15vKpFF9GPG1KGp3+QhVMxdKGUt04/bon
h8XeQRvuyikKzTQx2p2tYSIhMkaufw9QbieM40P5R0ReWv4VfbXa2EuGUKfEpNNc
8fdC82e/0YmtdF2mNfNaHoYRhC3yefajRZORIT9GqMSIZejkCv0fLPijJjf9tfoh
75SqJVFygJch8GDhYvm403wI53Sk3IC6Jq6xTLjpsrN3wZNx7xpS/JdpmUyDGj+T
0jScwb7yx1IYKPqYXkzLJHj93KmsdrGWxA1RApa4rCn6owQXrSDkd6SGg7JISddy
VyGfUlUUkBonavAY0BSqxjFHx2W+pQVBGtvsjXPnnmIQdgKa2JXHVcLwbvoaCGKA
yuKUBvor+Gz3j9KAwg3HX2hDIJ26PQ/W1Sh2PtMrbUDeTtYXGGbQQiniLAaIMWlQ
LR9QLfyH8wrCwMAhD8jIDBRrD4n2XEoOG0x7N6R4ZMnjuoJETbYjPrEw1Yw0NSyz
Aq4jsuonM15tNmuIeE7uejH9BFOPSaVKwAnk54VggTPBsyFAc8P52qV+EyA+4A3C
VKEIDNOJCw5QXf9FMEw8FC0Q0EYmGqwFRkwSM3kRLUa+uasZxwWrzIoAdPhNbu58
566cSsXyghFo7bNhr6p6VVN2Mhy5iBT3VWYlAX9pPkLbzI/5oOd62dYib3Kl1TXT
4pq9YjTFw0t6UNfM8Dn0mHLCZ74y7z/sC05zymz7plt0aWs9MsffblrEzFlydvaM
NbTX6nuUHcho52Za4kAPEru9EDR6CghcXpGTJnURjLJU3HowrH1A1Q/FLROdtphW
VlwpUk9jBZGz+H52q3Lhamjn1bL/IYEHwbbnCh1KWRhzPGuXYBobQhzozoCBLPDG
CiYnLRh9QZI4AIssMuGfyCbzjViIgQeKIvmYpsBiZxmaiyVupmiAXk9D23LJP7lf
cPzIQvWPkjLgAo/TjY2pFxKqTPONS29+MF7k0kkMFX4OuZqQwKp1NnpSv0g4hO/8
OhCfBFD0+QI/vXtM6uMRrOV6PCqPv0IJdHb+STE0oxyKTc9Z1mV+mTtKdLzXi4z9
p3Vm4UeHgX+/coqNhrIGeaIQ2dZka+QEMoOxQWeN3tqIeJoP7VHW2E8bBNCl9iaN
yFAStRCfbqETeiIOreK4vAAu6sy09JRYnxGNlkKWa+CFVNNwftvuuH/nNYXwaKhf
+472Okcol4xR4QVeXmC5Q6+CuSucL5GCdhb75H2rzfrhJKGF0jxwCS8g/m1IpCpG
7A0508/5OlPOfjfT6vJ0JCbR5MlTag6rzoDfYhJfmFiLRqTcq5LZGIJ9WBXpvZFz
xbttCZXlIvj5oKO/S4cJmG53aeIoeLne2xw0OtBLVFyVTtY7OFd6sVuYo0Ny6VOH
X3AC7g0Ta81caL8PporMwAWjfVjOhBw0wN2ZhxywDIOceBpe67ZDEPcRJRIx8qYG
P0PeX/dbKP9MuKNE+drie3ALkFbFHC/6pcuMCMoMm413n3rpXk1Oixlf8qLbP0D7
zAui43D06GRT+VJtNvaTw3iIcpMpeNh1M5iJkI3LlmvCgvJHCRrgVfoKoaBDERfr
5j/MC66IDFCu6NrjQzJMY/SroJEyJKpeLIUy+F9/eX4Jyydu+mDrWiRarixgPsRa
hzEGxEQEhdISqCp8C3WeujlLn5lfABZRfweA+bCXO0C0ct+BzEm9SUjEs1xhmC12
A0ZPqEE/JNV+VodpznNvtBi3BqUTAD/rzWrMJntb1h/SLbl75LoDPsdBTzjP+iiH
lveTvZM9blawSdUvHnohQZu4fYDrfwA/8+OZY5+pDinF1u1OgqLvowxhgn2opWLm
viH1Lm06R9Rnl3/aKaccieqZv0XGpveTXI/pf5j8B1hllPgDi/LR3NAlwj2iff7F
iQLWcAGbVrsslXR80sEazTh0p/aDJpcjq2DcqFffODsgkX99MJWaQKAjNPDyjf0H
MBLaonsutq6DToohrHFZdYc9LNOIcVbN8ylUY18emGaAzOKGkXUgmKGco4JSesuB
QtAAEWVbS+bQIdkDgNqQlxLayTlf8LlCfEEkaugCGGLkOj7PtyFJweast7USbAhC
SJMFgDAVfuJtJNnpGRHyUixk/QiU2Ykve67/6oAg9gBHw7Il7nUQIUk7DmMyIPO/
zYryvMtGiwc85Tf4KQNHZcjwnLX2UN4p1Z3uMM+NIbjq7r+kdzMmGMWGucAkoO/Z
TiQjwn98HpaWnUgFhwN431piMoqC6eJBDi0vGErsfUfXLYp6zdBxE1nNvnuPmf7I
gnqDGgVI/6zsPOCHFar+TYIBKVz7E3GrSEiBbFtrjsZTjFt25/YnJ6DlLoiFh5cK
wfec+fBWi6RdWMagHyLbzSi1L74omnhNtxPMuDvzXv0eFsDE8oqBzEnypRLv7dMo
mZzwPAZCksk9wazUhQAi7m1CeizukR9JmrA/nDmxIoPZkmntpLmupME5jEx7RYOu
04IchtUtkMGE+LwsC29aM8Uhg+K2Dn81d23gsJsEAGcwWVGRKxkRXKxw8UGVR4a2
2ujkr1ZC1I7xLSMSmSUZ4Ee9CTSgNjRsIVhejnJ1jUxpE8IKXQvmvrK0TfPgCtbg
T+W8vM1XMQxZIHHbTLp/1YXeK3nCh7WBwo5HN5aYRKbLqEpFu4lBW+vD5/j6DDci
WotpTl7H49HxGorvAzPVOcfW7FO9cwbgCjUrxc0D7j000ubNifA5Svh1YF5lQoq6
2cW/g8UY+uy7wpGivYsgv/2e8yNe0ipCpuTZqucHTfUfu4i8dQfv4A+JC+JcZw4/
bbPXcfndiRfHAR2tiYTgEcyd5Y0sCa4le/etvVceNS1QXA0o09gtazLK5Fa73239
5FODBFVst6r5EtXQ2RaOOwHQzAOhffbV3+ySczLfNWsPS8zzO0sC3r/slzzKTeC1
yKq8XKMJe5TAAU8CaTwKoj4qy3CprWNUHUFD/uBMVHNcuNDEuH9FspMhHT6IiDq8
JCVVSMosTUhqfAWCa4jdrBFD70gBYgpHz5boowJA0wc/AIKRAX1hdpZKRrnW0w/S
cuEqlNgsfG2/wwpuntllUTPinNMZ3bEq8qFp8M+3lh/NakQIZGMNsTqqiHzaxLX1
flGpk8KCLi3wZOFjpJ0ayDrTTNPlfw4qKlqMP2xlKuhyEWv7XLhHMmAhA0UKho0d
c+RA/f7acFG7DVG5xnTyiXUCZqcd3S+GFZ72C/Sa1lnT/dlpQExwovG/oQQGGHjo
tc2HmKfQ5puzX4anF7SG7e+bNurOIsY8ADF0TPTdbUknIBOGxUhw96xjznAp3uto
bkHTBJLkA1lNomcBcljEyPl+EsKIkBw6FLFNa7Po2wwMBizhmdJ6E+hm2meWIb7m
4Y10ejXHPbqJ7sU5wTGue+E50sgKNwEeqQAgKtOE0WMDO557PUoMo/WUzYvGdOhk
tUxCB1C20xND3ny8l7nDVbiNbEzA1QeUCxWdwGhY6Xytrh6xq9ZiIHR7Cez11euE
OnBGOzxQXLzJM4MivGAsmEMorjBOTNFmz2XbT4tLPxijbraQ+JoY5DNM+FD1Oiq2
hvKUOxPQtPBa3SEwGY4YdcPwMqUdyTe9kMIB8I+DZ/01SGJRvpGrfnMQBo/74+4u
iZj+vH8kvlGlNnKj9oLo6PwPBcQuLGjCJPJxVkVIX0/+FpsK469WyLLANbqWHNQJ
7BKLYBcMtf6nVKtLNChrwMDxXvn6KVDD0C+DXDB/qp05m7rchFzWMSWEVgr8EYLh
tjimzQpJ79Lb5e9zVcTOOrIn1NshcMAuozGIBtkXQ3sIeUjSLIK9bCmLS6kERnIe
4upLU9teh95HmA+/B7FH5IzSn1jHRbPM9CNaWVj/yesAwUraoDm0lnXUuuGVHpGR
4+L4qgTNcKxeJLMpzIKqPExwsxgId7E+wx3v9vOohT8QQTZjeHYZPjXQQN4duVWe
1WlUcAucJKKYlfBu+fLGdfKbiFtzE1deQjKa2Ys0Dy3QfO4u3a/emxRPm8Ugfoc0
F+GGdeChBzkJQdyVaSROTuqN5tSnbDHGANf4Hwp4Cc2u6wyHIBojoA2onx5N5QL2
Lz3cCklwyC2MIatDN7Yu/zeY002t1GEm44jGZHC6MXFsP1tstZmhAAVPWgfov16d
/yw0G5Ht18JB8PSuz8ZK/XCbyi9VzndtbrIiBwHJv/+xBj2s1YbtkIBhfeWH9crU
/gfNj6cxAqdcYLCeiU0+scRn0oVg4nn8Su8pTo2+soX763yn0RTGvkDPcW8IKVZ4
Bg+jaySY5+G+HpchT3cZdJH70P+0jzmm3Ga6VGl43iGJf+60YhuVxp6CQLLtehlJ
rFgaz/J1lmB6wqYvN3WCPljeGWpx4gcwaB1KubpNoo7mw5O5dBW3OaRKAafns1aK
QNGfpPsCe+iwjQmMaR4QeUFvGYjcOQyN/LKRRKCfJZzvColM6dqgWmQO9qYVnj9d
Z3viktpyBU2pMPtsH0Kkcrr6A2sZk4EAE9EDFy2JscaJjZG7KfyZWDprEhM/7eWc
sw9aj+H6v4gGIFPit/VGxMdprbyFR+k0wAipA4ojXQ7ropgiRfxTkqYEm8/+Rxu7
XBlzQAwImZQz1zOuZk8ELo0ptCjSmoHECGBd5KdYwXTrMJHcWpICpROybDg/2k/y
OYI6OhsUDX4EXxOUM0ja/q9a02f9EwuCWBpO0XS79qzopLKy3MyOa6dNDgzntyf0
7VMVOSyz2jOnNu5udTE6OymGqsf2jf92+6nFvUXc51lfuieixZZzMk5wb8Gmv7PU
mfwOdQhRUu0yAJ1kqCR94WB/HiGfT1kpraGwFxjH0Z63NtK4fJC0zazycLj+yu/W
u0KVhAn8OzCw8sBB4bHejH9o9qyswzSqfVEtx+hHpbpl1SBl94u7JTCRvFYC5n6D
jaYA3tLWOkBy7gObDUI7QXcQrofmTIS/d3S5phVq82lciVXMzdD9VoegjCljMjlt
shDqhRkqF27xGfUlzNwyzhzrYwNwoUV/adJQm2dcDNINUokcc8/zWGI+ntM+Q9/7
Kq20iHdcbM0cugQjWW0kSyP3nhhNhFSoNbm25f2VKGZoVw4XoLFjmf8OAqJI5DMe
Nlw8yI+ou7KE5c5tQzcJ5V/rs8+4OWelSMypiFRA9N07Z8aHwf0YwVGg1/5W5OG3
pLEkjfgFuQf6aIGG4qsZQGmgUAT1K4y2LoF1/B5P8CL+bP7kphv4CLT/IpcC5qr4
gbq46cEiapptXcLDRaP/RKOdHwWPVGCnoOSlcKsaCEPadFvRg2HIShhql6AeyQFg
g93mkhZ4cQXYmO4Q9xb4JrmrQNIaTMXDD6KIoFKbXJHFX+ZxG1pGgFMgEygojOUP
OmW685WdmwsJMxjpw5FL+/zb8vX8zzJb8okkr5MRt4f5b/yYtLrJdguJ5iexzub/
PoOc1rIk2U2PHz0A5ALMQ08HKRa1M70INmHBy9oliBLh9iOyr+wJdEnuJ/+FZPfo
EVFG8hHD3yEhnLRsx4j2DYF7fDlTCSXo/CqJEXPNsSdcEoV2s6ZALxASrA81fYMM
uIs4CbH+5yC8wMgmh9+nPRG+CCojqmjyg+99CuGPfqrIOwJKL4J/l9ZMUHLcyIwD
WkjssFhV6jFjoxdbWrIxuum3DrIKkvrIynnGYauDPuzMPwxGYFT5RdwrL9S0qv6C
e39Bk7W5C7qCALA/sIB/26HHrNRRit5wqlu3Kr2wUCL0swwrTWTwuKWM7RN9QhbT
Wfp6+hqIKJ9xGFYvBVZ/W4F3hhxedqS9DyhSzNccJjLCdQ3OI99ZwuEZWwEsk3BV
1ze8Sj8I73/tgts6UMWiip+JEcR9VzmMkTBAKCGnAlbOTJiYuqI5MkHNoJ1Oh/8u
O8irCqHJSy4zwnUOy6TZ2g9abQTdrUrXf9/tqLwZ5T/epiok0q15uGTX6p1z9FaO
Pt4NRRvG0CAAVFJ3RT0rS4Tr5nsqgtvvgZgaowrvjmrKcC4Z/hWSbomxF1Xzi0YP
isr9OO1JxrIsjP9yiFH6EjgsbW3Hz8qwyEVcvK+QudfLZnG7sd5epG2ek3h1oAf9
7BVUTQL9tA0kjGcCD1qqtQR/UXEu72PUgc20Oo/EsOM6Yhdx2EF+nwAvAPhCjA/x
K+JFdyzg+IdaAFBs4GonDp/65EDQ2l/T1Oj7dGAGYFvPwwg1UwtIcvNn8s7fKEAw
idUjD4KHI+kawalexFG+3i4dZwBboC2qc6K8MjtHc72ui2jUrKEupbFNmV2ASJ75
qfZGf6E7PFvemJXLFuNFRbNPtTXe/i8PH+JsadLy9/ZdvYDU1Lm2ZD+9SdCVYm03
Zp3WF67jnRXsmCiQrybmCkLulptGL+M3M6WKCx2uhDHIwguWNpuj7n288tdoIPE8
Bvrxnjt8SxQzi/1tmifIUWKi/GuH+mdBSph5kWrjRNTISyncNxwOp4ia06U1jOiC
XDWp73Bz5Wcgk/nP9ErYkILnoWiRoU/vnhmjHXpjAx3ITp0qN9LWt5UugebGfnXI
DrDCwgfzK0VMmadKvdjV8UH1L1KLZrtbJMUdkTnJXBan73DArZbN8fUlCgu+Fc8Q
oEzgpd7mAtw2MppZXzmt5ON3peQkRP5D+K3vPSLTkePltoL1HHzTaI9+UI1ikzFP
lTKU3/kiqeSUrgdC/gSMpL0vU7xMiHO76WWaYvqgOJMr3Nr6WhzIEKfh2ppjQ1+O
BMJB23K/DxHNbXxH0PWJYOCA48z14dYzQU9uxRiGwyP7zXdrL3b34w3DpKkL5J1c
2g43twmhxG5TBatAvjP8v5VDI7NxJhFYYdSM+UU3NTVvjGb+DDq6Ob1JPhG/uAhT
4BByJR4kmN9R2nsC+1zOV48TLqWe/v8ABmuC2fIxGKHoVytfzfF9+0PP/DihAV9X
1iQvYEHipi8cT0kP0FjXI1Hna3AkTl62FCZ6JZZmZ3UZUmlBebSQJxOL+kx7+OC4
71iwyUKa/iNDfaU7nT2Pr36lx3VCgCfStu728DLUv4328tHe/FI+CqVpJ89ocEmL
2GI4BmmlRu40elLNp1PBAEUtZpL7kGICyPLI/epuV16PGErtlRHWTJ4NntQ6CF4O
7pjgzrn+MFtMfBQAMYPdEt1rc5lzeY4yD6AGHoqANgSVq1xDRVlhG/PKlDiasB9V
2DWljmU6/oj3nmjbWw+/kO8Zk16zG2568CnBqaDHIvNOg2t1/0hjGLh4xc1oYrUI
Q+esCIdRLV3nHERgNcDfwV+/j7nrt9ol4fg/nzzjQRt2WX1oLu4H63YxDhTZk+3N
OScWVMz9mlYG7yRzkl5G2uz3cWsPg4xVI8bI/eceq1Hei6SRcopQJZMqf/bcVPnD
h2IT3x0JU8qLuON1BTI+pHKJKaleR0LaU93jh27iY4HSCwbb5jXTF2B4Y+b8au20
WTiRRA1lQbrGHTydn+Zyag9ff+NBfF7/fY/Dy4IEP6t16AC9MI54ZfZVnliUVEpA
QCoHEVMDqjVpB3zPElKStU8t+ZLU0A0bZ0ZmUqN4avK4fpVhLKpcYLbr3uyegi8p
mtNhHkF/SjVw3hotjBMP2KCmougylV3LSOF+IJOqi99WzXEu/5TCkk9Ow4K4J5Rg
o2SlRac7ML4xG4U96cJStFeFLPlIbdRWXsjaNZcRZkF5xZiXyX9iXTWmg9JHNmVf
PBxPRdQxaMt/MAtbJOvoCcAIc0Qec7FsZZ8AG8Q2YfKt5HfDiSIzVRcx2gW65d7n
a9u8MvfAo5zT9UxxJW9a/2JUWqwMR5M/K/clPtfqktXj+iHFD0X6rQfVJKOHL2d3
QXFtsvA5Hs/KEkrD+ZL32qyBHh7Zf6uXbadtWQfkviMuRvdJ4Nc3VhTIZ83Z48ZB
sXeS46fOnEG4mlSFxadjYBzeH0eiDEiIZL7oeFZtAj+TXp3CuILjbKdXWoDtcRYg
P0I3CeVOAyNUmXkNgDIkI1qXcIGZlYevEJNDiYsPbRQgjEN6Pd8JLk4FNwNhSu3c
FzNOZyolKRbSQxfs1owxHvdDf9APBaGfAfxVaugN2m9+M7mFLWfAaJ3PZ76yleOP
LFM5vSaKmyDGZ/1BDqCf9eom0YxwKzrT228LS+DMjXhgDUIKRTQTdBatgeobG55W
y1dUGPD+8g5zCvQ4OkRQYsxzfXfu4YMsXfiktyxcpCXY+vxin2JBTM1K35eiMY1a
tBHAC89NoXzcpgt/AqnPU4SnVlVL085AvkU4mzCCPyMZjnBT//5aPmeofk3JMMiA
vDhMd8LB2/n5p2E9xU3It0kWTqPYikAYjYIP7hVp3ZkgCmZVvohbdUiMWknW5l2K
HTZa6jzpJqh4LnCemVTJ/Rg+9VWtVgoamuT0MBM6gGvOIySuriU7R2+UiHrg/gH/
+oKA0XVMQcTEDkJjYnVQfs1y8tsSjDui9mne3A/kKSyjrIRxnpzi1CDOWtzqioq/
UKiHg9hMDcyb3a2xEy6Y5FZZYRh4Dyz+sJ7jB4fmtA1CKtSF7t8HtZX3ba8x22Df
P04KjzlqHDDnCtZwsX1scuo2xxpYOBXqDXvAAO4/qgd4XGDNQItSZ/piTuBGwNWN
mPxHIDrjGG1Cnj9TBdfy1lnlZCI4+DNVkXZXpv0eqh4SQrm3GqvZ+ZNiTZuAIUNf
PXySOmrzVUw7zlRsZ9A1bCmFdcdovF1pLag6Hy+K6etaR2v0WEl4ceDbRYbXimqj
F4Y/6f7Jc8igdYC6ilgIGwDd2WFolWaGeMuNja2P4DDb/Qp03r5ZRM3z59GLqLjD
jPmu/9wU/+OsFOEzf+Y6gPdrfgbhMElnuEzx6gLVvMpuRFEaJAbk3K46tu1uCdYT
ObbQRsCXJ8qgwJvpVVg3PKUfXk88KrnC35xM8dLyb20tWX4khzkL2dhheJaUydiE
MkLjZPyBXv/SIkWdKViPaDVA8qWatYkrhnzJ3w/jZXdSgBtPU68DpHOUHY+D3m1v
6X1na8O6Wt6epR0/vCP4xd2DhkDE4f9i1G8+zNYHs/y8VZOvB2JVP23nXrFliaM0
m0HB2He+e9YvQmGCVM1yfLKiNfwnWt0ECCoXENGq0QOJFiCfJaqyBacvJ/7f/8a9
tvipam4xKFvAZoC8eSMZKO9TlDn3zeDeu18yeg0IKwB6vw48gHc3+SpmOlry60Eu
5s6v8PIReADbk4F9zU8JysSRpobiPtDcIM8B/wFZ/gORUR6oI9bFg4Cipnxsh9bt
k1oZO275cI3F5Br75LNqmGd+uZVFydAQwjypiKlUZF/E/G1sHpF3Jj9BXo8SBOyb
mjizzezLEdM9h0KYCczioYISnumtygOHWbGYFKcAD7DhSYmzxFYiJTfvGiZcuLAv
toQJFBmCLFgdJNKbBQMp2EkJ79iRSDSwW0Kl1L1mFPoFXBuWw47TN4+MrF/Ao7y9
mJ3Q5j/0y3xG++OGUU7TM4E8JP26inJtkgbbYP/aDUWxv4p/qRd4fUizxZS5kKLu
5lAQOq+HPzmMbFnNFeGQGWhmyu+KPPMpR72RlvZAskGv1fUaZQ88NGfv1Rt+YkpS
UixUgDu0lkxmzmodIN1095ZXJk7EtMdru3k0MP0syVCyTIyd9txe89tEHXo1EgtA
Bz/OZGL6oi+z2/krPplOEIsRDFhQsKsGqMnDJNDMB5DYlvHEM9j0POqZjtBE/8Wn
gkXOFqXISJ3UX25sk+CgayfdM1SS9eBiv16esOkPNkFnBM/0ACeGXp7QHedKuGhi
nNq5khn8FrmylGuhfLPKLTn+MNvCpYREeXu4MXBjsPIINUGjwgZ+KWBZt9uidHSM
lNiqNdsGJ60UHaBTBhLIlTOYvxd7WpySqapFlDzwdH0175U6ukR1UmMzYZrneesU
uL5BEkla8TKwPInRbpc2/wiXoeQmqRAAB1265pwIHkCSQXuHVJbGH4VSp1g6FCom
n7CJNSWPHb75szfyirEo5e1PD+H7Fpb0Rgoys60IepZqCC0R6EbrBqDzDZ/u0RzM
tlV/hgaSM1CcofUZNI19W0EWPl16C4BjSGC5lfMQbGqhrPH8AgMVMuxYAKyeyswa
TzLjkd86VWZEObuwh6BbOULiKmPwnk1Pk4IxEa1fNBT6GfYqSrF5xDPgcN7wPqkb
0mbv5+uPNtLl2Y8+zMMwUJSAvpwiDLxdF4/Gzfb5+ROi8egMzgXsh2eQ3Zk3/yOC
h+XSDFhncQsmhnpiMfM4y6ViVpeSNQ1F/IXJ4l0hkECelYbuhqBoV8udfg0Y4uzl
yoryZqcUPokoZkAgINRVlC6Xl0EX1xOAES3krG+e1EZSu+GBY5YwwWRsCFzKG2Mi
EdP7ImbTT3dElnaHLf4dpV2ZHG7x2dbEdFk3eo7a/QzrPEXL5zuq+G80x/bMLQmG
kKl+IBkx96N8sf3NqbLnxp5xon2ObdKR6kxgS5lIH/lFpxPJMIrhrygZ/N2m7Y39
26unj1mAW7qA7Oy4gZRkPLwV/B9fWc5aLc/6sHayxiSPS+4JCQ/6LwSMEJi2QUvp
GNuHUV2D13Tc6mz2c7iA5hFYMHhS3f8O/dGagzhNFXaQiRme5vnvS4LNkbO0zMlk
XcckMIACGXRZ19H+e1OOm1Z1k+iEbGo1eaZiasb5Ve1JKnMteC+mkEgnusuS76RG
i1zABK9qNFcNQC2rs6CzPX01dxtf4LVHmDk9c0bjw/tSZ3RMAVnLcL3r5dE43yuD
Pd+hocARjgW4UXZERy2b8WFUXYW35mD/LNZYYho2PKr8RJtEgDGImLnRY//rCWP1
zOke1jrz3gxYMMDDCFikhVGhfqqPMEj274c+kfXPpuEyJSozJ5WOj//RrmkMFiro
u/XpTfGy60zQyOlIxrkcY9fPwEB2zXof2mqC8bUctWwouB4Nc111TKULO59T4xq0
IySTrjKkgkZsoP43q0qsWTJ1KeAXcXhLRBkvdSFwXAX6Mt1ojU0jQtMdtGgFn1ty
8fG/WM+JxxdGoxrTXT7uFJ6Y5fGk0Q5zjd82VSkEIMzuGtuFNug7+T6bo5sLtTHE
kIGSeAY218XLPpNISJnxsQbb63GKKNMFlPgRrx2tUtIuSb0kN0H724zcNRIbYqWO
JdgouskLO0F6GJ1LEL29rtpp1mIc8VlJuE3i/SHKnlCPYTyXFnVdPINDPpgEuUoq
FMF+jNZb/1CEhBE19rlHDK6scUq6sePxhqHgNj4esPLJ8tBl1nGpe4xoz75+gyVF
gfgjg9Y9nJORBCw20TvKrXgFh/+0NpswzSNJmDgwIe6FKi4CbSTflPm3rvHMRVXG
/3Q10KXjQkJO5dEqp3bK1GHgPIx/tnU8SalG1dokBApZ2TV1uADcFAQYEUOnoKoD
5KjdAsr75419ZWSt9+NM5zZCNrJSyK+31uGX/qGkV+Yjb4UBrb8e/Ng+Ns/pnzcJ
4Hcd32oFXtaI5gGuaDvg0fnMxJoudWx4Y9S0u31NM0iMoQkxHKxYPxNPWIB6hxX1
1I+/hqbOs70wvA89Oj/cfGCGrN9ucryekpLRhZCrMAjVSX5MrUDTGsWlVKaw29e6
oyKcpBwDw2CVlqMFnXz1E66nb+/+iGPo3fxC/SWYS2yLU5m5ymRwdCeQteGMJyBS
MwBFsWXN+z4EyO9AY3zSsG0H1TB1Ft9dYZRI9Y3zvd6MdBXjh18kPsfWUY+Q6GnQ
hGYE7va5/54JBoG+x0aw+tdMjwUqrEdyVbmXbbZaDzhpGtDMcdFgmQHRZzN6O+nO
UT3RhzRTaU97+Sk+UEP4QS/7g1JLnr/IVsRdf6ee37/sT7BWRa5Q/Ki1E9Zj3XtN
tcvjwcAzHJss75dR9+Zmj20t5GcidaAjT86SGCQBGY8Os3K0TPBY8yV+JGmqc6S6
CYV3HJiQ6BalDZTSJWrStsgRiHcYhnXXSmvaZKMAKY2VKiZKihZiWHd0HRf5NHcR
aSVwPzmfS6x4YhuSrRMnP0GeltTQmWyMkakDJ2UrP9JQLq2lXAI9tXkH9yM1+MuO
VOi/rQ5hofZxFCBCjkIeATaSF0KxHQrXDH0YXCsgTldRI0/aRnSIqAa4GlJM5wKb
3+ZRViyVqwkTLJ+riq+mfnX+OA6UFlRhg3nI/ZGYzL46M/QPW6B2dwx9NIDuUm6M
bW4BEUrzbo4wVezyUKok/kKDZJvXrTcy/Cw97tI8Ve4FvBhC95Zzaedb+nEcpIAn
1siURnc+NKO5O+42KPPUzBq82x2xJtut5lBm0UExDsE0tYcET8yLWo98QTQ+zuw3
E9eY0C6Y+ucuqQqgPBSFk3VA1UHm4N1vJaCDF7jR+0SFUwX23y1TRlA13s/uK7v7
FAhsLeRfG0oHdmCA7OlOyvOmekUUMMOcXuV1qBGzfZsqIvYY7gTpDKRz2W76LRmv
2sOKXIpZ1N22o9hpsGXcbvdkHZgCcn4xjVEf6gS1WJktLzBG5DIYtkLP4nP02JUu
nYQD+WxUqj5HZAheO2bAqoKnGfpW003ChngBgwToCv7XyL7hsLNquGSIr+DoUhRo
t2w3bP61f6v+UuTHhJZiGp+Tx4qXbh9KlOELQIrbUfQcx/tAi+Mpbo/RBectMvnO
9I7EHhiXm+WieyTII0JTfmOqaW39NWWMXsHGIkLMOpmsM3CBf1uGSsPTN1zMdsUt
EyZevqdayeH/gmLuRrTjV78xs4vEW2o5XKPTa41GsSfouCg9A5lF1IyZMLXRjQcU
F6bjbuvEwRBLbqnEJwga480WznT94PHv5vaQTmOjxRAHYIMNrCD4cRtLUik/XIfn
EXaixdKbICpUlENcy4Ic9nzgny1HMufFT2NxGpV7qvfY5DbIgOkKxM8rgZUY30nX
3HGqk/AcW+GgQTUUeEHAgfQwjcjVY2kzvI5jI6sp4CopB3pqUu948X5H5WVh7H80
kiQPCB5MaCCzzObwVtV+0h+UOo1bXgrmfD8mN7DZMwiqPKAq3BGqlrL2I69fDioC
Fk8dcMUkUdl/2BsxS8+7q3U+S+JZT+eFibtbthDAoRSx6+MZxyNiGX8nuBulcD9T
Uyr0FlQRUykqrrZTXJ26MthBW/VH3R3O3VF5IATcP0VdixYcak/xLeCcGictFRT4
3BB5ek60nCEgIjZ6nOPIY/LFR/qLWKQZ6Lup56Izf9xEZD+KjBn7+AONN2h0Te2l
ezj8Wx41BDuwF5jNwHbeRwz3JgwwqdRb3OCFj46xP209gZos+45rewFaQP38XKBB
jA2US0Cfn2rRpg+GCiVJjZs6utivF7eyo7A3rM4NNKNU7KJkfIxOSWbwKPq9jOgi
jjBQETDDp2XSVV9A4WD7w1Ng/OSjm6Bf8RjNDcjqoNVVnQhhQB5kQ94bEIJK4clH
k9m9k4NxvcSQxnnadcYH7htk+WE+aX1wsr/bd3yGAssb2l9IU7Dqirl9mE8P/bEd
EiYseP9ll4/sRE+MyVJxbGX85w3ZrC7m2KB9tldLuGZKMkglBmfIkKJH0GCwtGvS
o3XcQUfXzuvwGgoAlhDhlKLY81PrvnFpymX3wa7DUzkOpX4RMLPWvBI6GR4sXkgM
l5Xdf+NB8bhdDTK+oI3ImOO/tpHzFO0c2Z2K/csLluhpNVP6E6Wm/owht27VFOo9
s4xJFRXeMvKCEHh/4H2h0D/L06inGPUalYnjk8de5WGDydpNLx27bfdszzsaxH0f
Kf1zFpOmhd3TBhvnzY41aGeRMeHm90InZ5RdrJ5EHKpFB+Sq9+PbGnfTADZwMdDr
nEDY2BS/rQJZIyXHSRd51v8vhvcsPahQO5Fjhtb4+p5DEpOLNon3styhc0o+zTyL
qiFLVbbgc0/EbZjDK/H/IhBweE92soIZK6lmMOvJV/T1jsM7gGzHSPBwCdFfzmc6
pMqoWuxrodl9tGlwoNLTcoKsLK4B3muOxBfQava6GbFeRlEPbVPYES5nFpUK9QwE
FzOcBd9SjYgF/kHeXzQ8z4LxXMlkFqWFbSb6Mzns7i4/pGRhu/iZe5/MZVNeNS8k
OVtOacFRzvAx85cP5cbo6XCT3beuCkNzBcs21Q53Mx9+Ih32vshacoiPBgGtQSB3
VdrDRHItLAT5XtYp4GdQIZbClC9uGcnKHiEX9vL2PNwKySix/VFlUavQiOaTy9R0
jbSoE6dwfDOERJZNNeouvZud2wnNQj0XU+kGxU4cIAdONmLPEqFAjgzG3HtfveUV
yYv/tRSPf8H3pEUQLxg6x8tVZDvht6vjE9as1/RYA5e/95UEzPLYl5dXnBMJ5byk
1/fU6lSP6OrouMndQw+y/boP93vQ73DZZnlMkokFRQ09y4AkqWbq3crtAi8bTXHM
k/gbw8Kl411W5ZArdp7ooqy4uF9G6EaWgaYiR0MxwPl5OJNC97gSMjjXhRfvycim
2pcnByScB1LGmizUfrwmRigrGIbfYSRlDgH9eR5vK1Zs0tnLFrflV21i1VIjD51y
RaA/nMyh/QEhsVYwb2Udq6HJfdVzfotdXXksGr2AnkjHpDEBCAxqs5NTBxIN0oJo
G09EV0q8P/BXixuZyf2+wXefbsvqSB5fAQClsgqz6IbiV8Axn3uSlngAk13usCEV
KOJTtrJInZ3r1vqU6V9Hb1DzdjTijUFWg/+mGNN30/Y6apZRKs16lidlKY7l/ISq
urI7IpLD2PbTjRWN6TFt9AIEkj+ZWga+HjfrC/wrrrSXoF2GGrpnhQEw1MaAi7vd
Q0x45kVGSA6hf2EwnqMft0fjaEFa76n7U+BHLZ9xFd7MKSqF722sOd8QDlQ3Asd6
UnEvhpXIyJUeOvPTBvgN2+N4OFmOfAM6K0wBoVqJG0YqIK/cIy9rMi2UU4iWoKUx
MDSZmSpRvjkEjmi40NzcvP3RTAhNRZyDv+EV9+vQc81xKlsmqiMVRJiquhv7txqE
AHHSGHYDF75wYn/NuLGWsLeb2XCwT1O+NYHJ63IRCKNFkG9330XCRmwCBcVNRoqU
CWtCq77Q5cYHtJQBTYCelKVfCHsyk22ZPnrqhDabbum4A5TdXNZNYz1xC2/OF4Ze
4E65o4733P7uBQ71uhmJEveZNxqVHdwll5/BS02TXgpEwenKUmGO9SFnDYjSl/L9
6Ekt/+62Xc+URM4a6ZxPuX+WI+XsBAEDJh5xTCYIQ6GN8glVLghPusv0//ZT0hZQ
96MOFgSGXk+2gAvrgXaoe19Fn9L0T79pGWV5QIRs87COKD0ea3AFpg+t7ipSio/k
SeFwATMcQi3I0/J1rn+ntPw3YMFI+VpAP6roODhND7rnsWpsi85O+69/rC/ltwk8
8bS3EdAK7Yme0/ZT/uQ3d5HEa1P4UAajFJfbQxtZc19f+Aj2L8zb8o+oPMLeOh0b
bbJujrYWgGRo+Ym1ZlFp1Jx0njVN1zZxJm6nVOhlMOO7FLFpv8ZMd76oHWIqo0qS
tF68YnhcWU8g6DOfdXo9PVJ+k9Q5CCocWFotPYpLurGrzvsXaD/OE6IpVxJ+uBJp
6JQkUWrSjkFem/b4E9QR720Rf6045yady8H+dByEQMxSqFLQZAF4KxwXt5fdqvX4
sngfbWYWTcaxp6khlw3IunSzw+BGuUVnAvGRaNr9Y6+VTCh3brapjxmczbJi38tq
SwIomtgrf+TgGkvuN6kTDCqIExRNGBjnIPhdYk1QB1kIpYKZd8/4qELH9xvrkANs
BkJsTKqmuTZ3yao/On1HOZZCEy1KxKV22Q2KDPZXW4UIDpghe2ggNxVDG+hFPrx4
4kbT/u3B3x79DNBd/yvZjyK9pcqL3oeEttGlskPxVF/qbDDvkYo7Y3M02wPGfDBi
IXXPEe2D3f2AAFBWBEg4XDQ0aSkXl6B4o2b1y9WrXjlsEVTFkKaoD6Bjse/RZQL1
rve7yLl2XDAtt75elfqnTiitgikZR7DdG0PgVp7wnqPLugaWC/MqmKD+srPvy/z8
hd7z08A702eGMAyRK/7xwN655TD0ItKWSXC7lCk/n8ZGKc1hbUAlgTd1LD1TB3th
kt5gP55vmfguQ37dcHbIr3dlrAKYkHiP52JnElYyNiH1fucaG1sGzbKrK/xUvnpe
ht6sXVMSNgMhSQzBTMOEBqhhvRuhvGw6mIx0XWMAvKayNMVSXkCyoAmrJzBuyCvB
k0eTS3b8MCOO1OwLWXPfLrGl5+HJ6HdyAix7XJPTry8paieGJ8iW65/ProNmyOQK
39o8nZU8iHdZhuP//FhiWUEN99GkqZ/zF5MkdYdWbk966LJXzAU2Uc1VYGbdU4Do
VyVrciV/Z3lfFq+hPN+p+ja7aaTaQ5bOepfGe3GeFAP/qoXA8r+xn3ai03UA+CbG
r7Cn74wnwAno5uT2zzGUEORUFlE+3UWMpzxEgmeDMlYR3JFlVKP8h/7XHE8J9onl
taDurh7oE6QVpMMmoyNAaf6vT5mN+pRPS/tEBHDBRjdYUf5NX5H6qUJIPn+eQGtM
Q87eK+E7nDYIkElsQ3PGW6fJoKQfvmnPJfqfwSnm5Jq4tMALM8C2WrVd8lwr8qPz
VM0PN/JkIYoghUUAW796M9IW0Aj66v724yaNIY/AkR0pT8DHE9p2vCR//g/ELrnl
IF/rEC4s1W4dxvvmiIFbCtvoloQDSnPoWiY/6RaGkg1rGrUcdNP7gRpy8JZQ8LfT
b3GwWDuyXy2l0tYaVyuxjEBAY52tfN5Udowlh8ChXMKjyfiziYIJ8qBvPQf703Ex
C3FuVGIHBORXdNYQAYm5jAb1WusKqYh/p4OFTD1kFNcHcLyc0I7V0IpV1qgUHAyw
/j8hS2KiK8fLlTQ+0sS8+Vlwvwbcc5zi7Xj//OcYEsQsS22jhnXSmwuq6oU3Gb0w
GpELHvcNUWUY1pqxYxj8x6PPmYYgdqgF8dSDta/4UMCmSud9iwO95zuY8/U7YHsE
UQ3RT+sKrrJEQGyZyZOfaqsDS02VZ87Lao6eRaEOAyaL5+ynFo5+ebidZDshSraR
lslFj4PsZ4P0/fktnWSEoMh0H+SkiUoFRPgdLtrzy4sD4929Zm5bnj6L4SnahH9S
xd1Y08yg9uHEHwWVdVih1fjKYCEHvaih+FLpo552HY17XmcMjfkQ5Fax3wKCma5w
Cx4uqkIC+rno2mhTv7o2fae36tqpGH/r9qcLXvLCqdTmzo0+iHjm+l47vgeWLagj
Pu06dw87a44EjJyLy0UOLCJISbIQqfKrLscXGX8grMqXdURTx7KIokoQXXQ49MkF
92bgnCfMhxftmogqCeAHpeqoTqH6MItH6gh8clpxcVjVz2xjgaCVUNUcDR6Wt+/3
DkjY7LBFMO8po5UezVoXya2yelBsElczZ8qs4+tGotQEtSZaJ5oGx7VLnISUdHne
fbg4iVki4TkcD9VvARdlNc3q1Iip50YU2+RFOOkIUWH8eGdXNKGy3yeqFo4JHiu8
alP7tvg27eQEAJpVmXHvBiELudLWV1s9hGE8gxq7Hci+P6s8Cw7kZ6cQ/bf9hYRB
rvtc90OeaVvlg14jrbqvqXZG1ZwEAIihIUDB47S7gaNqabBDIpcEhrQrKoIRVDmT
BoipjRHSVPlVlY3jitDCi5x2zPUcYJjC2/6frGDf4YM/9Ixc9XPnswhfoO5HVmx4
yzNM7bcP8+nztiQyYk+HJllRN5c43w7Gubd3Ey4bwKmE5gUfRroAy/60oppezsKU
/b29Ibkj/znepa80UTSQfidRXSrsgTCbrMsA9oqL4KhLWu+JBvNlZI26tRd81PAJ
DO76GU9Cuduc+5M3QkfycWbspX2Aazgcc4XYfS6D5Zikxdz1qyUp1GGzw8S5OXp3
mbh6AHbixd9jpEYljuj4Fcr9ftUSya613wDnb/Nc8OGpEvOEpdkLdNCawn++IwFm
DNfBnZnp7/XOxlZB6ZufT6o2QbGrNjpC+75AdhevzRxv7Y1XMnxJX+m90Dxcyt6c
4QhSmeCsftdsAayRdv2Uhi0OYEjDV9NA0kPPNSpBtN/3uLxsWKwAlstR1S6okcEp
83aqN/oxWoOyJLNxomaevtTyF0pVU0pkywM0TO048Nw/kI+rgpOKuoeFY4kN6J9y
tqRbuDYevNBX5DgGUaU9SrgdoHQbky7u4xlxyaJi5NrzIMhzO5Fl6q13jm/7wIIx
AlmHfP+wLbGgrJ3AEmNy5sgRPN6Sp4Z0dhWN2OS0QmfW+8ggZbmD6zWyHkgY3hr8
WOBe84e3LSCWJUeVT37blmFlbmgnjjOUTaLViPOxkiFFShxniLid6qHXmZHcdbqJ
zgNKCst1TBX5hGSVNzi2YLnuhSyIF+U7iz83BQ4eNAyLszPmd126LTvp4WdGkkEH
7PQkZvoUhCCjrstld1NCIVDb1rnNx0/ULD+Fw368Y/YLqJz7LUFCmKcK5mhKDMXe
UBUS8AGC3AS5EmNy+T14dU/AK91ULCkRxkFFvEREPy23SjIVBZf1AdiNX9kApqq7
imQDVfsI6JLSkbpHsQA3YH/7luWokBIUuta2VnMdbtzHKgq/YVkbPGX0Dnyz31QS
RN3+lKAeQ1LaxgFwDiYjSSxM68+kFuNsP8q7l1C0aV1fbzaxwHYNA/qsEYe3V/OT
jVlnizLs8xxdYlHRvRfsgZOhlIv3Vn16msZcZTPjM2OC3jvJdkVRI3a5OZkai+Dm
I4HodS4j2JLOnLyfrb6WrhIxjuot9SBQiFTMPprx9Oqv3ACvOJsjBcZoJGvO+a+p
JzmqJ0RJMLLRsekqP4jWn3kBuFgz+XOyrqlRKL8BczKHvlYfuRShTCQHnnrqz8W2
GMDwW7lrZBWYMk2RBLU11hCu3tCj3Uzdombg8rX+29+R89iE9i2lPNPS2XKdHyFI
vtluqNjvWMBeGh0f9rEa7548rZx2IOR5OBPoPJl4f96N/+jSBebqtYsryix3xCdX
KvyjF+U4VOImypZ50rgpz6IaunQevXQeBs296eVYhh5SCmhqhM6gCxG1UxxNOXsB
F6tAnDgy0NzPeIIs8uvGGBbyH3Emjl7xftpLwHv/S8KQiosZPqjaf/dphL7t9UZw
mbekEMnmJT9jLGcDizcHFrlRAT/W2ELE9wWNXax9b9F+0+/4I0NClas/ipU55W3f
beHMMnYcYSRJdMSl5hLAs5gmj/WZhugYblQkNZ+X2iHZjzyMXbg7jef+IFfTW+55
ZGDAxE/7fmelOMuahPEm6vyF9DvmREc9aaDbnsFyuKN1ErboL/443HwwwzlXQOKq
HR0kXlimRkDaWqxNFHyhXLtbn7S3frHSjzVqqvobFjHyYvUABa8yK+1y3IFgdY8n
X9o6vJ9d9oDwuxa05uGNw31+x5YH1+Aad4hUEEKxrOwqa0tnBIrk5tuy7+oqhT2Z
GNRAW986smOUrl9XrhlE4Zw247xy3RvxvGEhXWCvku8BVNcMeOAvW4bz5mOvtwvu
Fph+7ygjks4z9kpKj8G8GKRD9ROFL4vava/d+FjFljROcd57rOoDgRCgR84RuBwL
LoNRW5fDsgv9lSf5iaC3M+52oKkAZadw6pOxr2BcvYr7Xn1+NMnIUJN9KOXcH2OD
mw9VCeJ17VrGx/YSOk3PfZFJKS3jKBseRzu2NnxmsSc2ghE5TtPl269qubX8tc/H
5G3D/89+X76oA2N9jBJjn6q2zLGbSI54g3can+5ca1n0CXrz2aytJD6KiZPS8S+8
3fYU7d8wnz9bnqkLmgxfXlUAW/yXwcej8rKoVLYe6eu4XWk2Gti11/eNYYTURQCA
IksGcVDMOqNIbV30wVqCO56cf2vWdKyAmuufHz91EiSIMk8VJe/KzTfTDnDfHkva
Adw37Pvqr2/pQ72mBShKKr2qxW0ILbJFl8C6h6I8bLffzT+J5t8KVsEPOQNTvSsC
Ry0QG8R7Fc3UiWvh/lEGAQpmiIEiXIftlKjO5z3/MShG4LFy5ZpzwEZXxSJqPZ/Y
KNNbjzbyXXmLmm0JHGRmw3APUXjjigZPoP13mQUi6RYh5WOmjou3TSU6KrT2eN6f
ZivIoT4qH+juu+3wtI1NXrArXOhdTNaC5sfzntUkIWJEX99jN4xdwBCXZZNDxjZL
fjzVeYyAPok2nyWlP7w5XHJGPSCsZhAJfPHdIBbPAjObyPnP4r+VQkd5nOk9SLzX
ROq9ygTqSmCGAjSQBcOhRiIJNn3L/LcGy4imuBZytEOR4D/Cbhjn4yR+qo7VsSOB
+rlyP2YXilpFD9XLuHOIxM3fGZGL0dXXkwNhkP2O9GUSXWy5gBSmUqNLIoJ8aFhY
xZ5eBOduQwk8bq8ZGIXnzzg40ApZQTdCxz4kxw5IPbFJTYdkU94SxnACQ3HYBGht
+1AsxywHftQAWX4lsK27JiW0GkClieTYTWl9I2dV765Mr9W61ecaZ7q50XJoP8bD
ROa4YpA52GxOKebtlW9UMRTTsvIZiGoUeZD1R1398l2PwrR8GiBURnlT6WF0E8bK
UKbMI6eSP9rg5OU3j9E0VvNdqmwnAH4+fDCqWRrSf/deJF/Euq7i+j00vIa/sDu5
s34g0ZcWGu+O3q9oGfYSGWTRUEezSb3Dwl9fk+181cI9K4t73pTLmq4SDvWYBVWl
0rBwFrSUdPMYz76PwzB3wwUVmZbx7tlyfBdGFJzOM0aTyPMvXQaIvlvC6+dTKRgo
zrjtvnI6S+FqUv8s/51vUpKwuvq/bWbYYExO3qk5VFbkux0sdqMhCSzPNfiG6CjB
COaslx0x7t8RgmBbSSZCNu9PPaaRCkQCh6MFD4Q3wmbDl6dpY9kVYUxUvBQUxN/L
Wp0B/Jx7yMjdBmZnYiUbF78HjphIoi0DcGOFq8s/zu6WLrDAS7Gjf/xBb2cPjABt
uIXMYX2WYzLIgEgaB5/SQzSqFG3p+za+hUjB/0gZZeapf7LoQIGVsphH1xq2dUX1
Hqbkqa5Oc0aTJKx3TPNyuMObpEk397lw1fsBtusBogysoBTNbHdmnTxQiaEf5hzM
YP/KAkFZa4c09N7a8Hu8QIYYTaV+v0q6zeCBPyh1Gs7crP0DSh1ZRo1A3WHEXLAF
P8VCXmQp5hqpjuVSMdacFQK/ivai9Ui0SNIthDOu7VCW3G6OlZv/TpYUHdiLOZvX
GBvvww63udzspBvhfIsylWCznSypznptSNPCvC/mpWogQO+JBhM02r2v/9Bfo4XS
1Tkxp8Ahwv7W2QVio84sGGcF81qZ68I6dyXSaVc2cQzEu+JjSLLhuoUV+LHQUP8J
gmBakcWCLXJK2GALd9TcFtSKH4BRC7R1CcCeL6FELVQ3aDapqdzu1kwaUBhQmS5M
TeB6NPv86it/JoQUwOn9Yg+5mgl66xEy8WtwQNEumc117bZK8pdhIeB/Ttfp5vyo
LYuBa88CCgrR+59mujHrWVEsn1VrS8VJxmDqrE42DpvgmtGCy77pmafD7oSxoYst
E1Hws3DjjW19EFCWIHJBTOo1VjGHhm7tJ7nsh1RGlTGpGZdcUiXCu5BO54Sj5lNU
UNU1ps+9q3BvHyMZe1jikGDzoo0vGvj4SqzzdOaEkJiCGxltF/8p9+cW8tZ91WyD
Z6WrPrF0JaSy69U2sUAA4LjUdTyVVane/1v6RedEQJC06it7yXxf3KcSCZ4BWpSI
lHID8e3kgyJy8FW03UGGyf4+ntariUx5+PAGIgfVKmbsiRPcYmDyWcJBu9h4s2EP
lHns+egO50Ey7ofNs7El4OeC1IEzvliyqyIG2C85l+e5AiC74I8fanpneHqbupZh
XGWdv0L/98QkqwLMxw/2T3Y7g5i1T9jBmRKm2xANm4xJy5x3P+TLv4zeo9KzpaRZ
UoqCEv2le0G0XwduPlAfIhSOFxszTZryJ/cYmaOuvNzm6JMT2ZIliJy/y0C5KerA
j/fi8VmDEy5WUT9hegjRkvCBDTnoddBivU7Ih3stVYOHsHSgUdqeZDKBeq5dMyus
URdyNjsNuR5dFvJssKxu/W1/sD7wQvUYHfsBj3GQhHaYbNoFY2XXF9DFWqSNWV4X
4V6jYUcBMCYIn2sFbmIwQ5oJzA3k8fUjZnxULxfeO9lzaAlFikeYiR/E5Pup0D5K
44u3qdGZiORGh2bB1Clc/XAMiMZFlsXYLOTFZc1ghZETQgz6ejRgCad8aFWSzW/o
9/XRgRa+q89QbNjQtJ1Euw5WZRTIvzV1kMf/DfFZgX+wXPcePy+Fb9aEvvBLiih8
RrsZjWYGAk/VptvnRU7o5btaTo6sKcOUk/mLlk5/ol6GkjYNnao187/+iMR49wfj
84FvrET1oGOKOD88CPyyAkHIFWTgxjy8rEjXa2Aq9HEY72+98XwzwqGvwep8nHl3
AnkjKKHhIlrx7EuEmJKUqV80MNAA2K7hRDNCNIRh6hRvvMs5i/xTZmd9ygTOZ58/
dtZJoFMxKrkrRJMM+piZLIXdL+5b1iTgXuom7lgSQfwYVS+ND661U7mD6EH6KUmW
imh/tIl+1s504I4oBdHpAxCYRTNNO57/miD8Oq5GeyyvbDJRBEHRwa/Cf+BW978W
d0c45hhfjEeh+a4Gd6qqeDqMpWr3KcKylYuUJANrAAIcsRIhdrn8gQ1H4YDeFSUF
4DQ4wvyKJHEjaEnzVEV+z9fe/KYQrYHmF5QCQ6Un2cBlenj9VlDPnugkbq14Z2Me
/U4bV5xSNhCQJ7tgzAWfM0abS1DttdopYGU1i5BivNVtDkUWlDdptB8DIeAA2Gvf
AhxqtCOJD6M0jd+xyvurNTrIz4P5//tj63lzQ9oR5hN5uTMq/aO1YLIExa43RVgX
c0baBFUXkXZEMArFBLy6lh0w6zQzd6ysdjlisiVprz8ShgwbHCxA2POf3kvn7cre
lYYr2y26lMd0a4/2X3yUSU8UdG65XUYO6SSXgrAyFe41ZGWjtw/M12FwyzzTJoLx
NdENoMdnw6btCgz0KWivLpNtJLLN3l/Kvq+X4LK6xLqsYkWdL9waLYEUXUCrUEU/
WiwurcDloGDW+6Q1MZj7Evm+YQnDHdcd33FglGUqOzxeGPO88OvUgOnjliuw75rl
wF1PNXD5cR2UMQERQASgAEJhyWdqrxu9shPKr/lLaQeXMKgYU/ThvSmiiGqLKjCf
Hi6v62J9Q+/Z6hgjeBI+zkf7ygZ9cGnIcAV0wT3JYeDS+TVQr5pYG4XfyC9CkC7C
TFwMH3rWQfWA04EzKzIDzyflQtNfoV92UfuHjw9n0PQalkntIxQfKpvKH+1EQl/G
lF5qQeZi9Xr1kOBmaDs+wqKp7cpUYdjRZHKaEpdxlLROCPL4oz9+5FRSs86aKygL
4pepyBVWQWDNLuYGkjOKJwBVlcbcew/+LTbT5Va7m14GYpUVKPza+btUNqlwgk+V
4zjiPJKPrAJZtWiS5P4wg/g6NhSzkRxRJNBK2vKTzF/KjqoIxdbCbpshGYPmPgey
n5yQz9lehUqMgpcjeDqUKaaZfKmOTE+CT3qRMbPNXMhdHC3gStQz6wNEiNC/xHUG
+AnIsrY2fK1iMlTcQLnEg0XSfNVmEbvzVouwqGn8gpmeHG3vlSi0wzVNB/grzi90
S7IoXfgAMLkQs+GjfFQWuS2/LMEbYU5QXipbMoI2OK15ApyfxEN5iSQN89GyK/0T
w/azK4SygQOu/SFnRgaDyCb8kDpzVBdskqgi2U1ZWP3G3/wlFvA0VbjRH8ozymed
jUmXGH7KENuAQON6Ti6BUpRbtf47Jb1zg7cfo1hmU6l7tO24cA3zBxxvdeudMdw5
ozRzDWdkwhN6mTfAtgrj7C3LbdPQBm9tMDUtsVUP5GR5VxGZuDYfA/1Qt243PcrV
AJbifvxPGylLsGMNG3Nw0EjNmpfS8o+3EfNfnnf9kEARkHeXbZRj0INR8ZqggLvl
XLzJkJajdiRd06us5X0mi0dBg4FxTGQ99YuMA3JZ0WYjKfGwDFwH1SuH42hUmBkw
tLjYOVtcj28eRPvSkq0RD6KJiT4XZrOFpjVQoLN6h8yp6/3w8iCPRd07MOSXOZum
2f4NNnerdrQO6SQASbgvwRx8DSrSH9Uaro5KupJzCvYnef6vpVt8gHZjPL6wmSKD
PmChQ5D0qp3fCVnfW/GkGD99ym3zkp5i1zl163HIBeyV4YEHOksncMEargk18VC4
cMA6qHuJQ+jLzNZofRH5eQSa55C8xYxCMXuON17k3qKgjZb18HuavSAKw3/IGXKG
Rcr/JYVSO0orObDAHIYwHBsRDsm6fMDYE+3IiFeUR/Z9v6xX/rM3Do/8U5sVhZN7
6ZugLYCOnqVgOFDCGVvCDONRgjFbshkN84tGbBJej7WDmY/hRx0XTH1/Ubh2jRKD
fZoe437QNTrSjHiQ48I4Z4AzSTUI0ChJsshZRMvb1ej8/Xgg010LZcQrVLzSOHYW
HoqnwvCusc0STVrtCb26jNJ0DAun96fIQ2feRV5j/Cl3T2L8QuQpZoPW5HN+mFFO
8qNZiWAlHzdGpvWOdTFyrMkUGhmszrxNKU/AijMPwgUvX99xd5cUjngN+HHx6NXo
9xGWl+CvszsqjjWoTypu8BRU8zQVC9BVasnQYXdKEHIp23eVe1cEpWzqL6cktlM8
HT7crlQ0Z9h+uHP/ruLUXjVMq2CXoF7MvLiK6bTZSz/DVTe+BbDDOxv8YP+D9YhO
wlkbiCsF9FHNa2UDPZ/HriHYiHth2A8z9Ul7sP9/cOt9hc+rM67VHG5Ifm0RkLFB
RCRmPCrKYGL/SiDI+EYyenExsYsWsHCfY+jOpHc9iWtKczVpjWMCIOSb6AlcKD8D
2KGNA7M1OJHbJ+V5XpUWwCMPGzPdb9/ojm7R/QYJoZXnzKgPmz7ajga2JjyfnqAf
3Kagne9Tv4jpSWKd9ENH4pwllaOXcJZdOarZtFgGkYTYzbByOsLDShT5Lb8uvP0d
3IgKilq+bQ1AZAYzaxdhieZXn4KXvNzal90bDAbv/C4yxHOdmr2hm3am4wGh2QOB
WsQqXZ5xqnOhSZICnIRXXRjs4teonwlDuJqkJtOS+iS1Z2HMXVt3p9877QRa4mbq
QEpXDgKQSNaehvvI1b09Hw3/tkiBbGud1o2eS4OHww7XnN6Ab0eatm4L/1S3eZJb
4B+pUQiz76H1kRYlA3vszrI3qjjN1DKUdn+XzbXTefntcmHpWyjY9od7o+XZH/02
WhJL+rvsYVuc0izJ0TvSsge0glIu78zM62mta2dwz2QUOOAUO/6JOSWEubjNMFMb
TZix2PNL+fzd7BzuRietbTjWy2y+VLw90FJsH5F69cZiJit66JR3ygHRAF/aX3PE
IPWd3U87B8xQLPe21vnAIuyilaLmzTv/jIxNppm61uauuMLazyw0jTzKqWIuEd9/
k2zJSDMMqjrTuDq1+Y1VYmvilUToengVVnUfh8yj2z9ceWjJ5nGISIA0Zos0c0Gn
auDm6yCnMcyo7LIHqMqdmWZXNYJl6ihq3E3ZEdaoS974pz2nUPKlQ8cR/RfjsiqU
ZaVLZFY4m9WuBMUaszz4wKyFOEIBEm+CwM7SKVD5Db7jEkWy5+USsTnqByFVfU07
4/aPg6H5jb7fxhUSWGXaYB5g/MFQ7NARL3+E8moX90VfjPU0803Hdq+vM5qC2Gcm
B2OK4VjbKAPQ+oI2wK+Fro02IMKjiHF3v5eLmb6X5mmhupg9Qtmw8WRpWiQA1rXn
7X5+FvuzE/OLC8wZSs6t80zt9PConqtO+xzZQqq1nvkPCrxv88jp3wEiPEQJKbf6
0avF7jv9FWDM+RdRM7R7i5z+oAQHINMnqZ/i0jdD+VHWio8Ombajgb6//KDn/Iv4
vNQKuIgOwIoWD9/sPOkRYYJxQFjHRR5CwZjluS4IFojqS/OjcYzN3Viy9CcN6bSH
FZX/qmdeltzVzE+YWqwdKJDS9Vk3bGlpxvnR2APXXZsmJjnhHnLxvSbB29b1kUD5
nFlVXldKDFaeZUzFu8AEVt3dABsiRDJ3KakXkXDHiL5r3ai1uYxXx05v89OUaGFv
HHXdh5D18mOk13kGyhonXKFM8uWsTqjxudEqEuBCutYdh1PC+IO/TrgnNFwPScsN
Oq7q4/2+ki6tuLjz5t9G1WPJMgmvazSdbiywvuyk0r+fwjWelSnjYaal4nJtoM89
ofuWWLqOXtWmK91Mrv9iDY2lbIDmQY6q980yw1LtRESQjszxXuA6xF4VfX7ifqmL
xlHVHnbJPCe4FUWS5Es066YsnsbHbyWFtNlSuynf4QJLdsYc4zKDAOInuyfy811o
xzPg6TWzRPaiROjtjQdNIj4LIWoY2NrWym9nVqs+7rEnPcbhVqLZsSx6PJbXfZLC
ZeJsC+V9TQgiyt6PvoLbs/2++125i1AR2RYMZPN27i4mFMfdPvpfhfYR6RQE5SVy
90n3IHjK6ipRocg7sTewgRFzyxW50+m4uANsLPR4r/49biLW6ijQpXH01C3AJ5Qi
R85VVpKNrmVPLC9mPpyj80G6KN+6Ect90EPl7vle7mfcc6xzpy09ZdakLO/fdRDB
iTvytQIuvLWz9r/oxIhqTQn3o3SfulN0buXdcyNlQHpsgmUygXM/IUA65xG3yR4O
d9VRySfEmnrNxDwemoawP8GAmX+bHl8yegiL+fZ/9W5SA/f5umA2qgER4mUBYz12
EFIFBvJTRkx44e9qz6oZ0lZ1le81yJwbefUay3FuzECSYItS1lk40/dhtM0j+xM9
FhNzuqKs98mQcFeC9oOhHsct1LM87OQ5fexXQOC/uRJ8pgCRj7MlDZW13l0zT8Rt
yGeHh0EUig/998KHA+ToTup7GsOvkiNo1ELrNkhuAjjJkPoG45Zg+vRqR7a0R4LY
lnI8VnMFzolZqaq0AnEHE8Ua7QNzueRQ24+dwoSkVltgYu/Cjdls12c4BnRgDbU4
Ci0rdOx8xG8X7zOkLqU1MgqzZpo/jVedUvASHTsMy18QCe0g9nlE8JKvx+x3d26l
SBoxU2hjbF1bfy5L835YX+NTPCMeGgP6V2zzfd9I7qihCVNOegkWFUaQvNbiklxQ
UXYzJtgMx9XvOFlNMc6zYfgSMTn1kfb6WoUOg58gEeHU1rMCwLfu67O3C3ox/Hvx
77myCn2Fov0Vh1PnLt4m9MX3TEatKwEnhEiQxJ3B9iQVle5ZTsQuaId5wn7ncgc0
4nEVeTUFQj0Wl9HhRLHTJx++trhQpqZYK1yHHnWanbDYRc2+UbT+hOtxS8nbuE0P
qMPBxoepb5W5vyBAJCDF6PxVTsMxyDIcrkayawx+CSxjFMjIlcGLDOEN8YKBRTFJ
oaW0vMPZ3MOHj5SrPCGTH8LGHqFutT8bBnZpPEsHiUolW2UsDNMOsq85M+eX5XJL
wbWUvCDOXOLuAnqEBtwvdyQ1ASKKdDRey0463BQT0hMefi8wmuaLZo11tsC/Kh7g
qJNnU8YydalKXj4EAG+0UhBaawQgsghVnTwSFEC+ALe8FPFYfd7vAWvQvFIJd1VY
TZjxuDAh20oTnnYji4IORIYd17OZDds+xXEVxJZ1I/qea3xiTJDQazB6YM1pCA8u
pa9YHKu3QwH0h6j5yXzQ55xy3nlOfZU54u6YMEVuYHJL8rEvxKKZ/vgw+m7IK8q9
XVrfGYfq3d1PLUH688bTZHX/Q+4lwHqkn9sE+17xs+ROyCa2r35DZ1ZRuei2zI+/
bvroE9BMb11OMj/UdxLbbJrGFH4XYhzQqJjjfycpWheYFVj6Iv5puKyf1MkpzQ9E
3liD2fn90EVtUtF2WsQ3brZgN+Lu6H0oEf66HqeaHpiZh0rc9w6wiJnwxi2NDJs5
kqBzEQU7yd0XAkGr/D7t1W85NYoLLBDR7SrmsuIb9xk9jq6t4ILzook+gT4mqNZP
/Q1p0dYl1QZKzh4kpeb4KesD3BMvQNEEMIe28d8op4AfiaGjrJpeD8mnqup+5TJV
PE4SXpVtwWa41nN6/Bli78UJdVBE8SKBszyf9BXRIEdZMv68jUe19zD4n1ZkS4en
NreYXOxuRzetM9d/SgJa7p+RETeotE6p7okbnBgMdx7k2xExE4RwEg6UJgD9A9KY
Vz+h8XPU0sXyBkfs7DSegVes6/Kv+/UMGmk/Ix7aSqbpwJjPGF1ys9IvVDb6da5O
CO7zfLcPE9KfqYkkyLnQBwwuf/mk634Ok5bF9TCqsw+G9c7s5qATdCvD8IwfyUm2
haI6FEp+RrL0W3e8Pw3t2/7UNaHyeifVEHKCmdyxXmBs5yFWgsQFcCEtuueybSh0
AHpVFlrbskoVOMZwYWkzn4iV5sbj7tiZ2FDg4tM1sXKGX3/8YxTDZNIFGUDZu/+t
k4hjE54/sZ9bgQSbJzvyPbk/84V43D+u5f4rFzAopRt89s30VTVxpbJpTTpDBd7X
OhC0hSCvWSjF+JJgp8Poj14JRAyOhJvFq6Xn9OV3pbquCGC2H3oDS6bzT+ETgBeV
0onztkGrA553+eWlPz4X+yqhPTCm/xhtEOEJwOsBFvaEbIiU9WSC5zH/QjvtS1Rm
Et910cUCoslNzJKykdp19ZjlNOWNBYhO1zgKQ2rHsnntOdX1olI5TxDSBL2xU+44
GUkJgdT/9/vnV5bx+vOh9eXUNC+pMFrh4Yd2k1Pz32XggLFyHUNV1Hdq5TVDKgR0
yk/GozEHVLbKFj2UYAELq3FxQNNEwBeiuSSyEk6L9uAPV4iDxRPLwdx/vhpAjS9P
RIE0fUUvNSe20qz8jT3ePhUlxrJ6Kr3NLE1sMn2mJdQcuoxm5xRHuElSEinODY3w
rxORjiQMh9lgEwAJoJ8J1XOMRHQ+mHDa+nEyasSWheuIRVXQOZmTUuFF8148jSyX
0yOUn1wbFTWnAernCA0LlI9MDGVm+C67jZ1i8PYkVaKHXQptBei6K+XA9AAqpkbK
0OdbkysxKxFXuzFLPNmVUtRGHL4ADSzs0hRemroFXydA7ialKJxGj2DdfVP78uyw
9qZiV6kFV8N0z/9up/cqQflU2p+iQWvonKeJy2Qmm2h7yDSorAdjkP8CJvpKqDvK
T6wo+aM5tpCF2eggTAeNVp/Z35oGA+dl8tSY/BayEUhdXjVlDSwfYh036vp+R65a
PObQTnTTOjz3tvtzv/Q6pD1M9G7kqrh7JLX4dOBn6B/5fBRQbw2bQ6ep/tP7fjqS
tOlmqnZYoDVqM0mRaVb0IGKzQzNZxgHwyCXKUeiMYKKCAqDVYxqj0LmlG4Vfb1SN
rrRREHtvvhmla2MIVsomKfJmxIjTT4pqr5qjFa8qJ1YNq+EB2ojHq9pZ4M1MQUko
QYCuHaLSnLWL8uPMvs51YOD2ogm4G7K81TPt2eGF+vuGp+pRt+I2Yo+mZWNqea44
LJGDjXbdfTjIDUfb5We9klNCytaXvPjOL8eZmkU+ozH26VDSGzr5t0b97NBQl77V
Lhdmha7HEpFH+y7M9wcRqH4QyUnuYh+H1WwSA9jEsSRL6NOqa8qTnF4ffQ6VSgel
J4l+M3ru2w28nzGNeOHGtSks1xxupd4vFQaTi/Z79vUhJZVonPViTVLrZMYBVuk1
1bCbUsKkNA/ZhjM86Fjxycd56NPmexKKAdlik+si9X3FO+OMHUxriNPSgXNPpDXz
uX0oXNHbdhInyGttadZGcAo8lKEZnSZXOhAGqH/9p+FY7blhjHrwrgd8GOQo2oSz
ZuCN3HqtKuKl4U6sn0mfAaWHNvvlbHnEzUAMzkD0nc29Y5/5ezYrpT/x/0RXnbOP
rpwzKhzvQr9T5vYU6fCkbexCQxy2eEiQ+kxxs0gcCzzc0rbW3mNEJ16Mz3Dk0z6w
mM2YiNdCnWNar/f/QpkMbeM4tn8/Mk8OBsSI8IF0HdBGAsf9+VydTXq5hHRF3yuF
P2cTCMnnxZvYm5CoaxsHWmSIAqyp0QU6PxLaZT1GY3aksxQG2EmPKVvtQiVPy3U/
vjxT7cgrHaK5wHqS+sO1+eJLM6yZt/oUgH+pfE01x1yXgQ9rY4482J5muDykbsWt
kAgZYlfVwXKJep7wFRDLj4PaZcxW/Czh1vztkt9LOx3sKxoW9qAHwXPK1EqHc4tm
aZ4N7QRB8MJsDH2RzGe2sR6p9ZG7j2sqhR+njAkxmAwsV+u3zTudeC3nH9vEU3q1
kT5WEi4vBPkzbWO62maamIycSirXKy7PbycBhJs1MWcwnJWT2RlrqojXm+LjLhxJ
w2s11VkJRvl98X7FuRXTLOEHbAJlTzXRSAbkP+HSZ9FF9hlzKuyLDFFUBr4wjSsc
GD0tXt+CXrszyMpgk/2skja/Z+OAMMYyun+yIxkdEdLk0waPuWUTT2PQuUhYgvtR
3cmrWZgD6+YTyBxs52JO8LVK1bTFg6zXDIYF8J8wd38rF8daM6EZp56sOC3mn681
v0CZn94hiru/GB5/wNjItCbyHIORYJ4OqfpyTXGkaPKYVNvv84n7yusLjp3k+BKo
KQY4TD71tu2bIiZmvPjH2C+fiXhwPBQpnKnvlILAXExWkTLGhqDEOPci21IjzNZN
UqCJA40I1VPMLhXh3bFrjVefXXGv9MWmZNrlOYIWH268fa5BLz45OE49ZTj0kFiL
Y3OV6Qv9Id8ObWjDYeZDFNN7KLmx2yxmp3CobDPon3Ez/CUlnBUG+D+R771Tt7BY
+c7LUoe5VX4YOmBPCLZTy21rlq9AYecu1830p8uapITSZai4GAYs46LIPNBpq+oH
K3VbXXdmT6KdACsUsnEaxCeR/63H4dg9HbOxg1kedLUK4RRjPcXlf+V4ODF4G9vN
ORGNt6jz3CUcPhXjG4kaoIfSPD+8q13DbYe+MlxacpbBf5ZMhCPnBaQYDR4q3u9U
HkwYNOPhb6XK8ZSbEZ1SAEi+GWOBsHO/Yck7DGfaYXcbH/lYomb+YJ43TzrbkTDH
0GWIz3f8+De1ly7q0C5OXFtCBUONfU3zQdnxa4cnmOPD/VMqdh0gQNNrpKRIBVlI
Lh6bYA+Q0xk4aqtn3c8ttis7c2svvZtWfRJ6BiDiDUEFgTl7YOyozrWCEIgS22sG
RwiW0GyTH5HDOEWfrBclY5kJkCij9cwa7e+kARus4KCVjlIH37Pz0oLsbl33/UO+
kdfoqFt1oMOR6qk2cv/AnLyp5BW+etPDOqgAJGJSt+79OSdeCYes2651yU5mu6Kc
eo63eAaCo8MsGe+gP2R/nNTEMp7U4Qp7Nj9u0bAUZDvO6vwO2rDQlUF1gWvYn9g1
8yPkAPAfDHdNgOCblAqwlXp+0qg6MDBX6GhCG6/3Nl6fpIQZU5rqrKEWY6KPNtcx
GAqqpOd4hJc6d6iSrfjBOYsYkmV4USotwTCdJuqxuIG3EOXBqEnw6QgNskfF9HmR
EjZez6SznGydJh6Qlh/V8syKuazNZ581UhgOo1XXxdDzy6f4WadFgRzvNa5Yd4XR
koOfSDEbQk51iYJNKjsMDbh1JgBHY5yB67HtmulqZlUMn5yaTGaWaXUq6pbFJQKz
7sauaZgHeCqhLlE6tlLUvlFy/9EWXT+o/U7FT5S0be2WzGiLeN4dhQB0JdLyYd5W
K5eCQAbp4pznwMgECTSOcmkjcn3c9bVxV/ewmXytTnsnIWFJElSSfahAP7UbnSCK
ItYbPaVlwWXHQBZfGyRvx54rWMjAhZTebsURftYv7yaQvbh9l6U+qAPfwZFmDIg8
fJIuXNOxLOLVtXPT/otMPODn/cDzON+p3GV1l9Bul4rey1nOgryZgB/nMARC4det
U91jphwQpKEl3Z6tLzGfsIoeiUpSvgh32EuErk+d+tvLmQm4/uVE3wBLJNIPnSq6
6tLUtsACC6jFVeW7FrWHtYEJVml2vivXfkQ4aTQHa74FRxNQNcKRfWyyJXXhfbCl
nxYWkXDoBTvt7l/uK8fomn1oxqJSoOvs8XXfL1utuXSpM12SPtZpvhD9fXrIC0FF
VKGkcAHzfXB3TPle3JWC2wuixMtJNcReHVq9rOT4vuA4lfbuR7OrxtYR2delp1LA
tmR2qfyCDZ4or7JfLvmWIv/+UDY5puynBToPR8t/v192waEutAHM1+rh6x2QTR1j
G3GX7dnJblHrv0NhOcDKJSO/KKsc5jDAiTz6hjF5eq7P8YHr2y++/OhgQ/7yge+L
zGYZirK95D6dpKFyijQKlL1p62rk53sDetcCuoZcmXEFKssE+LeMF8cicklbhD9Z
4PrhOPBobKyaeisMahUKfhzpMU6qGAIBWpbKn2wuZmUmmHbY/ll+gJqT3H5SKvtF
kYjs8z4LAtfmWn7P3DxCjeznf/eAVB7eDbm/OzSjL9yvtPBAB4ZkP/uDCJ/0/xzH
PDLsrY5mJ6xnJVBM1Sz8y+FzPjHxNn/+6MXp8+Zsv0/DJA2/sLkYBdjHT5Mc4Aha
viJ3auBg5kZf3xt6qX3HV/Ibw22qJ74KYBY8LnXrWSO01zPFL8LBsH3hXtZQkESF
Jm2gvcLn3ZL7Gkf236Hji9HCDcd4ll/H6Do39yne1zFHsQWvDDzCG1Erql0zTiB5
CRUjLBV6lizNU8Mn+iDctI76sPX1AwiOVl5ZSD4ZO9Wiz+9OLqESQnf5GmNhTUbH
BXDfMs1vPoWMdCwjzgQL5cab4NvbtZvh3NE304xsuGO5l/fO2W3kImDYP5WqHRYY
P/ovbkDyXbm77EG5bshMuNlkPc7B3WFi7cPGzqGQVbH6TJugwjyeGjUfBGFFp3gn
ctmx1Ft9bhN8kB+Lt72AzwlTKpsVv1fq55XeOeTipMBOu64+7XPGkpleXMOUBy9o
6g6U28vv7d8bBaPuJTPCUy8KOXKOURY7BYLURSZoUN4G0p5SvjcuK8rnzHpl1G8D
UiOZxNo6qghNFiwaDgqyCa61yotmICv/HQ7pg2i4+kAy8X09jIWGtYr2zzfLlCon
s4LghtyMW3LDN8omH6du6gY8e7AN5zjmhdttltLVGe4geiDUyi+scepDuLtWLfK1
joVwZQMcCR5JMWhoOqnilV0oE++yjkHEh2iX4EF+04IFn5DhRYKmqy6n00tJ3Ozp
o4YnObyj1+8Ish+u9dLW0hJH1FZeqfG0sKMvZ/pqnmjVx1y3AjIi1Kbnup85MjsA
Trq730g36htCjRIntLC0q8YHlrkyfnQ1CIyS/0caMAhGfszMUVw2JlRbjNFMm0WF
D5HGXfGHn5IKIOK2wSEKrc7TCBv7v47+z1XU4aHEQpnMi08F4OFOMfXd0jG9drKL
HDv8bSLkvSVJNKbJnWilJ3DBVvIvKWmX1qjv4OXVWjOIyLYpC74lgl3Ne2JkRRH/
PdBJK39bFhcarzs3qVOp+Li+fhNwdbmp7DQdKgx4iRjKSEdO68IDLDb4PVSrsabC
l1+IEju0Z7gGRLEYWBaPlGdgyIaXEDMcpDcIoyUpcSkS8yWH/iefxc8EaEZhBCdU
02MRZkTiIwxzOJItGjpdmCr+IoR6GriAJuzWQR9x68syRGIQ+UfvUIEke6gVsp0d
C66AbTk4CNDEJ8WhjtPlx28ndifay5KrFps8HBgQbpBA8pxLe8jKk1/Qk4xnZUzJ
Z8uhtwlld1MHCXsUN9BeoT+ahgLWZ8j1syNWef8fo9nGTSt7t+tLk8k2ljKjalPI
ysb1IklAFD3GMHmdIvYjVyZouXEVPHGFeUT4ccACSmRn8RTP60ODtmxit+ZRqw7U
JkhKKSS2ad1KOEKMAeGpcaEvkjEfF0v/9DKNHxfSfnYhYga9hcoYUNUMgnJuXYa6
ORQfC6t1BBWwzD9UlFmu8wAREfIjc33m3VnnL6qEhJUZSnI0Djxa97Tm2tGQeOTd
YyIhySGwD2rAVbfiR+xRcr4GnlIj9cM40dO2Lr62Ot4iv1vIxfaauYOnzaGVRYB3
wUi6cyPk8nIO7e7OwMWuCkv6/m06NYXwzhHdX9Ghxyj01OkRt/wBNQFqE9iAECXX
sMUhvQGh7SCWYaULU3Tanf8jDHYZlAjJPmGYaKt9EMX3A00hAnJRCzsHKtDmkTkz
GewH++AC3PVIcBB7PgFh6m+9qEX4sy7pvwlaA92rJJWR4FxsunBR/vtUjQHn9xAT
mAwg2ig3ccfjkJoPT73LG5xZ0xoYTt3PLHKWaljutLlty80GXuScgW5rcpUapbJ6
Z7+lu3C7bZ9BgCezI3YLLI7ufBSidZi5pla0zHbcEM588yQdXkBfZMk6RP+w4KWO
9soJJlntayQ9ArHVUux8nzrv8MtYzUo4THpLDJxuub8u8ultG9XpuH1UtRMUmkuy
sSScFGn0xEjDg3h6g3CVwZGkW4KSmRsEIcVZIeoiAUh76zv1uNSkwd9+w/KuLgv1
ILne91zUMqhUkH6GSGwguEQxtlW/ezXGaLZhfGR2UabYChxXnGI73VzFDhM4ed6W
s/s3AzuGvYc47huxsugLD4dIE+1w3WBEC1sSXdSdn++MPhM+YpAy1Aw0vZrRkBIj
O+M9peEVVYxxevdCTZ5HF/SZq1Ku5iiRwmsdIGL0sM25Le3xGfF4cVEGifZO3Yol
K/+3eFIlKEkMJRhNz8fNtSAE5QU8Q/VAKAFaA5387YpJwJxhiQVdTNgGQPQg/G5N
zxr0tYktkAYLBBRJDS1PRPA/L4FMX+inn7RAII5uJl9Ck8iI4jEODma6RFComVgd
AqKyRu+I23/v+QW+nSXllun3TTUGwK9xAF15HEToj7jtEInXGk4xbBPhW5YydMum
SoH2defZfsaBEEqDzb3LXb/mibHsgHF8jGoEJiXwCY0CP+v+eqBE6bAE8Bd8e7UT
BtmhFigu5fqkzmm2AHqrmBV6gs4QmW/XriOUf/cKb/U+hSuSsBAg2PsQhyQ7ukSV
QZN7cxUtYEq3eQ4ScBTRYO4XLdpr4G0v1V7dDz9P2FvHDKTGfyX1UWB8vJeKyGHE
MWD5X7A+YjJR5mkfm7g2clGJliHqSMdaccW7zK3RcQM4/odkjAUN14JVK7sRw+MX
GCcTvTRRT/rk3HvOCH/6o+qcNWqvBDsdFkbkCTarULR5/nlLf6bGhhlBNgJS5g6m
76hoUMQLcg2VOAGdwqKPWr2BXBOeqRJlZngTNKjNTI1TjCZE+ibPyCSgOO2WHiOR
O/X7KxGJ9kiijocr4/zZQREWAlrM5gWm4qd4bLsnp0XyjYFd3n2xAApFLo0+mK/w
OzHY7BVjBdfIN+pt+IvYorePUt0z/ipoAEPYlsER7FSh8or92saD6BNgcyCeZY8I
94Nq+3uAQ1Me8zG1/9OPEtxx6NUC+i1dapJzAIyzohM+FPtmA6Te/uTbxnSvhug1
zAUUdV67C/IY8biPc+N5hlWiptQveoUDmzMho94PYKH3MjER+Vc3snQTdLVP0P5+
fQDim8q49lUSE/TXKbwpUD6t0Z5u8NQkh3pTmxaeiCC5PkVqwkhReECUFjIlRg3J
ngM/LHCO+D+ao9yeDXhpoBnhI8Warar/+fkP7sgnFLSXbUmNFrBQMY3+ceWXCTQw
i3GHZDySVtdlx+s1rmJd6DrHo4ZWQmjLp64Pp62AYP7Ntz1KokBuBqDehOdq8yWG
trVCKhuJkMLVmkMnhEjCAJISmohqYvw5Brs4oFcKFSXKY8cFlVufTsxrMb/QGAVO
Nr9tv68pNO2VUN+7mbYVD9BJGK0rb5t5vSDHInKPdq7V0+3N0F4HUrnbrOSbLHQg
i/+XqAA/LabhySo1qbSHjwJEVlrQ44CSCrzcAgHA/hj7Fh8g+o/CBIYAJNROIQyf
1bRtt93JQ4UY4vvA2Um2W4ymvIwhQA22dOt7oxg9vnrym9WC8jdAKjVXsTKZ9WcX
7symKUDZEpedCHI4XXdI7gr9s6w5tEcj+Bx4/O/ySGhiq9nSH1cdYKT0hg23wvCg
ogJT2dimXEq5JJKYuO+BDa1I/ex3iTss2L8guqHhsUZretN7BmB33PXLpr7MGDG5
trDzcqGOHuEp+1WS30jdHo1nqXsjPA+xiud9aTbNpQuK175a0aansPrxiUlkdyI/
3afSWpsb7QhLWXoeU/jgdpXRPlqb9qjQlNsiHFqP6bZq5bEUsfWd2llvjIbQ0ajo
leZxMkETuCoegQUiZzLNSp1+/GwJZCgRvrNXFE/qC8aNoVSq7/DRON8BlRM9weVT
ZQ9iiRf93yZa9fBX5dy/0dTcHJp3WAV33mve1EFAKU5L4f44BfKQSO7htb5mrEfG
XbBvVQ5tPYNAFSBvwZ1WOxp4ajWpwWeFBZqFFIb/PLr0wMpB/dhYxA75B6VGC8Mo
gFiVjGBzWbtT43xlBSPN+lfzXtIPSBvmyXKOzkrgkzWNG02EpaciDe5a0km9hWZz
UjqGTHVcBycPaqlKySnmikgJ3SjujdUxW8XoFBA/ls6WfAEOLwdgdxVnlpLo4Wd8
ilIQazpp4werVnpyA2IRcXdmx6WOhz7r+n3UOyOygjeIQrWgCswZQB62vB2NpRhy
CN4TwMzGWT4KNjVfOJNsUNPcwirFKl0Z6zqRgNye6NP6LPh9BnF6g5VyP9p/NzHm
0L97PL+gm+SHNFpraVxzqVqZNUQe1dTW7BII8OVOz3Ie7GYI1cQKV3PXb+r2tNhL
uiGJeCIvcsVOrqqUqPtL+MGMobBBbFEYcUtoA/1rXfPmrbWK8Y+XaocfQo0pdZzj
2mZjM+s3Oii47OMigNox3+WA6FKmLcSprM7wYB0MgZxvUnmvZm2Q74u4QYWAktoi
xh9tgb+L95zxtmYqiW2FLS6wFf3Afl4y7DVjue7BxqTTkRzBi84+NFv/IT7K423w
PlqtLuNCasdRH/hiIBX3qdameq+0guYdvlc+733vXWlmWIDQnjj+nfrW4RpU9bf5
X0/QFgfYukoAU0nrFAxbC36FJDy/hg6rpqWvCLDGpg3CV21TmV6NN2fwD+LbL4dP
DteS8doK2BIvfY44sU+VRraTIAFWJaN2mhPVvDSIgB5EmxXE9VpvwEyf45BCJKpH
XAM4nCanXJctnqUsAN2inFdwRFiDgJE2JyTuhu1yoGYAwqdEtEKAxpqo/wPfQVrY
vppf9UY+Wd6r6HJbJDU3A4pfZpuagxMpJci/9IbRQF6OaNldJ/5Rbvf2wmE1Ugaj
OGgG6gj3iQI7CfZYuDahTemElcwGtpBYmqafCN4EwAWbysmOpB/E3zCvZ9jy36Le
C3fAVSQ/9qSjAclSmqFHFqhhbPVG1Vr9UzNI6wVkUJPBBc2ftVINoJBfw5EGulVK
RG17WU3JOi+o5K3+Edjobs9HBF/j2yPex+JSWCJICEVWO5TfVdvuMwMLCsliCP+V
dfr2P4S5yXWQWFS12nwP8frh4UrQaK9JtmEk+FQJMX68/5Ny4V1zA5l3y8Tx4/W2
p4Xy1zEhojN8vCKN1Lcy2Dm+/69Ohtg2Sz2G7tkTGfvSM2suK/QuvqmUKXk9H68o
BSLRldo7ARDv/Kx5g98b4hTGllkEY06BuArT/TRM0M04ojWEqtbmv8cwRpuSRmnI
IFd0xf1l378kk/3mRySWWJDud0n+c1uwecQgFbKog8/5ipD+UWEZskR283SYgd4X
p+PP/xjWEZ7n7hPwCSNBfuz3EMjTWvRIBPILW+y8C3eHogo7pgiq9/eXkA+BXiKM
fQMdPiWvczaDlCZb8xlTbEPok68PNoeGAcJde+BrlrspQYt3O2IVq5RzMDdheNaa
DSROp6Y63dkKLNqOrAawVYFur3Zg2v7x2SHvABDwMQV4m88+Tf2T7Of+pVbl4sMn
7QRlx/Z7utgyaXc1XM4GF0FNmYc7/MuAd5wGdz9IXN0yHo5vVvtKx6SooOd2UIky
XwOQs5fI60z22HJeW6P6CLsLNBk2H3s2Uy/G6zqMemN3/rnIiDF4IhWfOW9tLwgP
jDYhi9Ur+SYjxUjarYDIoTukorS4Ah0lGp+KTUiSsZ29CXM7uAQPjdpAXVssFiwj
wtO2z26zVUR46bbKEnYDew9GlmsdqzhCMghyolJus1bsbxU6SasHn4rfoXOqO6OG
nFqk6UhhMtiRpBhnbeKnPncnQHEfuormkwZI0bKGmN6u9iP9O515k0zXUCGGvUek
RxK92U0MqrYnKm6zsCvGVMvzg3x8Fr7k81qNqDOd40IVxFh61btUuTtSmmCTg2H2
HHJSTcTFepmzCWeBgTfjEab7YuxaWxoR3MjYYaHtTnBEKZSr2XtuaoHQjNR8UsK2
f4uiXGfG6LkvAithOxkH8sKiBMhIWj+yGnmADRguw7JyoXqSqkpglx61hA3+Bbfr
t0iPkrjbGi5e6I1PVv9ppE+o+krYLbI4/tweDjkTX/TLasJ7eSoawQFJsmhv9cG5
8ic8v99NE5DvTkYjUtl4O6VBJI+WBBTw/6o6npV24lVuA0X+3A6Q+4+L3/60DQD7
cTm5+knz5UIZoRwo0UoIlX8MoVMP5avo02+7CSb/XyFoLoZEiFs8o92moi8JWh8C
NjWaUVLUQS99LGJcerwj9FCOiFUdI01rszsee75AXKXoOSjhWGVZTIREJ+wB2ymp
YX2Dpd98Jq3pywWre0drzm4Goj/OL00sqKjmu4S2XQzgcMCkX+KrEi0fqMla5fb1
l/ohAwEzldrf2ScY/pJuMr0pu61PlBYdBcZ7UnGmEA0995gAtOvdVtRgwhVnOrXp
kHTod1h/Bp91z+zQ/fJpsszMLlz2sAmQP9Y9iXxP4DAzNNuBCiGh6jOYdxct6G7z
lDZD60GvMIwAWNksyWA6rx17nLtfuEwJrTXtFhB/br4i/kx2cXIxeXRdYK4bBpXd
NzDeye3Sr3OR+cwf86LyzYXcWVRfq71CVui4E4c3FyAeER6F8jb5gugMdXRVkIad
ILl2Q+mgFJGV1qKn5esOL5O1tPaptmthsfodidEuPrSQ1TmKcqUDqpkIyIqYWCgq
5QuqTuPeC8PRlIQyonOYYPzNk657OjHcmIcTVK3Kr04YZvXN+PWk1hAIUcx54tf6
lmeeCIAZ6CMKiDoDaiXl8LwFe4TowLj/BT1TG6xTQAXduhatsWrVNQbFPNe9aGYf
EFDG2QjLj3T4VpNihZXbDr964Vz8HWY+VEpLXiyDGyqiUr8ZS+5VJ0aP97nbG10I
pW2e6R1suIlwRZVy7mOzNOMufw0yQVH0Yt1z2GBdQkUscSXL1yVxXSQhuHx6clhb
FSG8Dt7r3Y0Ia2QW+tGMGwbLb6fN82uIkFIeIBH0l1eiwFYJmgdNuD+12K5NkSYu
GkgmclNTtP4HqY42zNEL5Z2ZhB2ojYgCjhR9uPExm/eFPyD3AYWlQHnQ3KK8dLoz
cOtpzGVAzkKB5s96KUkONDbj1VMnO6ZLHqpxLCB0MhX4Nc9klrrUmjw8IPSeg7nR
AZH0dUlj3icIO1ykh83WjxOV9cACWSG1FTxR9ysS5gugVOO5RJzkavC+YC6G7DtC
0kaYaGEoOflxr+NUi+YI2cKfipZ6Rx4h9xzW4NifIEi6BoMrXMVbER2GsurHPZgb
Pvlwmoho2QrEHGbZuCToKYQDjXEO/2BT43pk1Beeudtmdig17Yye+uTNiHwV8+/9
ZtGQn+hbtUOuMYRG8ShGFLMSLjIra/zHQ9WpH92eTB4n0wbJ9gTyoZVWpl88TuSY
xZGQF6uY1wuHMat3aiEQVmw57MIchsKeznqsClMRzfQKRmF+lCiP1DPOdJqG8hhz
XNlW6tC0v9TnobZzHdeQFlcVJNdzPZrotVSB5+6WOy/WpEb4FI51Ua2RIKdHgRiQ
jRT0RMPIb4IDlZ2qySIIH8Y+1LsXrTU4zDn6qgo63OcdElIvL7HGrZKu9KSgpSvP
j2swrGtQ/WOeQHvmnZIv59oXNWLW27n8uNJ+3M7yX20dm4k7Lb6hWcuqqmrGvn29
kYg/iydBM+EeHbLqpQrfMjukGN1SToz1L8reISFgQH4ZXRCGTKavRyzYm5Gl+C4v
9CZeDRzgbHIJ3e9FW3RylU/vXASRc/j8jqw3RKAW2tNSK+EIAEj1fo8I6bxl47QY
BEK/gFA/P9qV+Cq1r4e91TYI5L53NrvwXr8PpmAKsLfKmTQZpW/l4Bje5Iwj/DDN
t0hbIcV5N60Kx219zHq6fJtzp+qQ3gIP/gKvgdTK12rlv1zPuQvYQsNUYzJK4qbm
vnpm0NDk98lhOLBJ4T2trUwa3091DnaikMPNvL3DhVUYjuIXKtLRvEJliy1p3BM+
ocz+JhLEp1Nt2C5JKR8ITwXCYaT+oFyGKkEih693B2YbRE9izfE8G1KtzVqoF1Dx
nKn7TnwmRbTbdruIHNEio97Yd1PBFfTGDrGdcDh+K/WPSA9O/NI16PHMOkyD9qMJ
T+YNZ/BZy58EAU1mP9KqzlooqTXpiCxyn+vbToeOicCUonI47WeeqOAHVAVDoES1
b9Tpr5NKAgvE+/Cp9bqY80heMPIsoIP1czWRNYQV1q1DWf3zsars1uczXOd2tbG9
u4SGK2clcTM9E+wJkO05CUOxMUAuHQRKgmK32LrsaCgXCcDud95wyN+iqAWQAmhP
55LYnrvm0sRKeCvaRLm+MMcn89Rp7nP20l4O15Dp4Ec/JsJ3gBqb5YVII9GyIA1E
aZDMdMZzQBGLZHhmjQtrtyf9X+bQaC3b161wpVFxtlBinRwi0Kqy24n1ijdvtUVh
M4X7NxcdCVINlZ/m6QcP6QNP/HHvPTJWZzgTOnLncUB/RMNt2+zFrzom/c06PVxu
2LG/s5q4An3RRxcIDssRpxPOhEPIHMKD/X2aqhtDCnIXChkpgAcsK+vbhQONnn3P
aljvkq0TQHazZRN5W9zuub38kboGTDvs3XsAp3r25u1BAbDxPoGg/wv4s3ulzS/3
qkaZZJEY/Med57szNFpRKLTxU/4Kc+qY5D+6W8MFZNJ0mN8TiKdbPR6zOdG8Np+V
YJN5iVrv0V0ADhH6G0tva/Q/UFAB6CK7pycvwwM2Ea4KW4DRA9N54GYiQ97azSXz
4ylQrZiiDP69J1pFPsXx1gcSrVWtIqkLjw/ZHPrrvQ3ZS7IkOWtLFxz8/vFpuXdU
0pxhSqKOA6aTjFSio/Fus1hknYccsVDlBs23rdkFs+9rjW8V2DpW8O0iA+HdTRSb
wKbSi4Gu8TiGZvQinHiJujLXe++/S1A1plkyR5EQJEszx+NlxpRzO9ln0ul1MuNO
1kKCR1e/ZviW6FdAiyYsXzjcdfQ5ZmycBHE1x19lL9JNeDtmk1J9B4bG0rQuEug3
jRSA9lEKAP3OXYZnARNDKIck2PtM3iMz3kt0Bu4oUDDhCsMaaRBVXyVJ/pqQRNH8
WOjIOT9+qB07lQOrrSNuqsHsENXHT9k45RpHGkWzHQ5d6Countho17yiedAA/2QR
csfng/MNqemP3i8EvAop4s94iMOH8goMyWfo70Ub0IZBZM/4jj6vgiXw4XsdV3tH
ezxzU/+Y2i7ZSMX4etK3LicHGhmjfT2lsobSrsZFoF5M1Dbj7Ot0O8c7Rwwp/CtS
fMIx/jM/IMKuaqEO6P/RksV5nVuIaUihUYFbqyzL/Cw7KwzAvg6N62Hd6fsm+bbN
Dqi6WwbpKKps6Upd3TQFMf5kPxVI7NAeHecqfpHATH74TM/iQ31ZMjJ1i4YsgeAG
WIJajZzqyOOmXjeImfT+/h8MCnNmX1KUj8RX5aFKVY+DSS/Gt93E0zd+QnM/oDQF
30iAhcmIgSgUf2Cuv6HR2v4juzmmiU8uvqpSenNN5EUu732bZ6QAaSrhM7aBm6Qs
U/gJI3GWtL/CnqnowN6myfzNp+7qOyphQ9RTRKpRsq0bxjDMOZm5Seh4VCxv3z5A
5YrvogvKjtEEc52cNe3QU2M9BLRtMeIOIGdlYFjFgzbXfnyssf0aFcyEKBibl79+
JSxEOut5jG0rcm+DpziPS7ZLb81UyU5yc1oXCCWJ9MKbagEqKmD6wVAhMg6lUZ84
PhtbWGsAoOexUE4m92VKpDagLjnr6HiVlxAxznDXa4JP0HIHFXIBr6V6czYKZKhs
4W6BNjX1jKvc8+q9zk7tHo/1YYWr1PP7m8WIN2DwfVkoEFFk17VkKOk1h2yCjjtd
GHFuGxxe/HJUaBcW5HOXJ5aM9/NnsewpW4f+QSgwILqurKlgqr+4epxKiN1TWScD
efxOjew1JqBVNlU37OeK+avO/lfroRr8mx372+i+q0By7PnGPrjX4Mg4CgZlvoJ+
RLXTiYtMF40+zS6Td7rz3dtUf4MSMM1HWh5ge785JAl0nvK7ZQtQcmQAosNTqgFB
LIaWtlVspOP0CjtxdVDK3SkYBFkhhb0L7dTdQB3DDfDfSGXebvkrGgYzirw4C0XB
CkZjgQZkGcUj+ZGWOkVX8/xfEQpZnWSq+hg3eYJe2mIEuCie++tD+TNndjcoKz7G
YwHAhvhlBKTuJzW7Cu3zA32EtgwBINoKp7G3rlr4UeUkCATllo1uOW5kf7lpH29S
qPW1v0CgJzLh6JrAIJ24QmurfFjHPxnJhRf+iLYq7V9DUhq06RCtst92t+Ilc+Mu
aTTqFvT2idHgKW9aTxnlif95SdhU/xDXaCiEL5siRR5bpKtdGQgo7WeWoIHVWfkA
8vsBvKhliGAiODt7iv9uyyF/N0UZSqg1GKvHc588nOhjWTMuS8pfw5Dgx+V7BNDC
jqkG0wCf1E5YrXcQnp146FQ438hRIpmep50CseDwFxq//EUE12I8CvFD3poY59el
7qX8xygmfSRmcyTdtnxXaUfBOcDItTegXX+DBfC9YeGWsH2X/gsu7VU0VQs6zLo/
6mZi9DC4Uu55BwqWvOke9zu8kwHWhWFEFIUIlGgR7z/gk/q17gLeIHkXODxEnpnr
lJWTWaR6NvR5FFbVdFOgyz3UDII0akU2M8/K+toq5Dl9RVy5pryvkOVfLOsPuVqF
SraUQ5OmoUV0iUJKp8AAgB9w1UoyRoijdoUfHMHbMCUPyxzSIHdwj8GEDL1jAOnp
d8eu5OAGrsEZzu496S+dCTx8oyoAdxrQePH+xaCteGQAfZjX/xA5DswdgkR0EJ/6
fbLUIePuBUr1opnq9LLSKcbLbhacNJI6X4Vqb4N1FPBL2yXg72VgzgUIhrJgCn1x
OI8OfCtyfB8dzsy8WPeTb4vsef2pKGnGhJ/3mGHnszM1Ii8fLwTpBYBvwIUyoi08
zCTXCgb2o3ZLAgNOP0NqALb3TbIGxIUNEghDxOuD+LDdrueDpxH6zmVsjKsG+OBJ
8t89Q7ff6+bDnWyI+yCcIZFsWnc1BX8Gkdh6KdWYcgXL4pmlMWHsIemZ5YJoP+/T
yzzW3+qnyp0WW7GetlrATgP+hLQms9Gjq/ssiNGe4s0x6U1ueKcrFGU6jwRvTPyR
eZUGov8Ft4d1nLoGHexpwz6YyQFPtSuKqk8URO8bm1MTzkyB6rp8m2/svU12BA+/
rS0mMR8DAmNlHSSLjLpku8LfvTDS6X4AfhHD6SFEW49S+B1QLxKKviWO8Mrq6sNH
YmCIwAQdrohBXcDuCJ+dhDgVDx+ZROKTKgi7G3rCrm8YXIVlrCvso6R+lA5BhBij
oyBj+IsW6GCaN/jak0JxKl4q96f9QrwrDqAI0phXzMGYxPyBq6+VLI7wtNc6KGIt
0+MBnZnMoMPNeWIrEREqEnTWE30lE01FLQsVPVYhWM+WW1qUXrUMKvFQyLS4DevH
dG+lor6p/8UjPtSvkiQEDsQ9B7qtMyHzR8cwFEc3bdoxva9OWlTDbee6XZ0OU8oi
esQPkziJvBVWyoM7Nk0RpUO2LnBjSndb/z+zZEyEK3wK/mgZKiPaOtQXKWP+1ae4
rEV9UrdDRSsVxqcH8uGYpma89eAIkgIBt4N829OIebRc8V6TkcVwbKjKmF/LrQS7
Dfk1pZ5YEmCp0l9Jj53mnW/Q7QvyozQ061ESE8lXs3NCkSwbOA/Q4rES3+9r7LVQ
jdFqFn1yDKLMVAf9Ol+qhopmFYS8zZ/TlUWunhIsAy3Bs33WfAkN/HfVSI3V6NID
MEBzPJ3rK28PKK4orIlbNku0pb7ncsBQqa3xXdEBN4ajMc0rZvHtDD7LkX6iLTra
nlFfDpb9EQ+6AtERnAtNuFcupY75tEKZvGNy3YvBpTFApZQq0wiKQ8ixZTVV1/Ue
UhDI0uxnOYbxGywiC4KwUen7V/vPlu4UP6J8EIvafkuwO/2US+N/QUwszakwo/1O
XlVaQwgHnwFJL3vWl1RvLZBQ9Ge8tfh5Cp/mcXXG9jG+W/ydPIHN4FjmplNxMZAU
jpliAiwOGtNJQ8kjRJqw4Ruy+mMLWEIUNj7swNey8ZZCALfdp175/Wk/hCaXU1Q8
WM/2fDXFbxPbOZMMoykliwDGldlZ6nttuK3JgWTpFWmWngvapCStGD8BocYMfyu7
3PjKox1MfVT66Xx6dbSZr9Aru0VxL1exjOYEaKlU3XrXoKYJlfSoVvEBmB2eEuzJ
aeum2u8Ay4nFeXEmuD+D2CRkhpl0v3dfNa1H28XQAr0wGr2AGjZcA2iF3j7HElsE
AcYX0o2MZZfLyJUk/kOyCZlyJLOD9Rkz4wfLPU4Hvn0k6KNQ8wpQKoxUtokQQBcM
J3Gb6Cp0Y2g1Ad2O2LNjxsaWhi5k8mSA4LuP9B4PBVr1Q7WbX1cvhIMc5Idp6gIN
wyrBH4F0j74XXpMy9akXmwZ9BiQ5f3LKWJ6vhSBv7hHh4jmZu1yOuldj3lhFSdir
HGolqyZEXt3YYydYXu6jDQ6D/l+Qv2VGM7tKlmreuBzbU7zrcP98F4VULRJWc3Wf
KjsStvSYFCS/cqBZHy2Q+pFuV52+QxfIq+9y3hRZ+f7fWF8zKwGjKmHOxHtnMYQY
SL0KndgPa+3fHVfvwKEFONVh1me9IYS4uH9IyG5raUSkpFPRg32dvmPKuGHyN81p
kiI/NbjWJI6794LR0M9mx3T6SVzZ8yeDP6fQI/DH3yj1d8YMFExvtDyexAweRXmD
k6fI9q3nwHLz3rI/L4HlGioRyJbAf5MWFx1rPPaRgSR9CEUUBrmGcgHa7D11/j2C
pl7hv2eUL68V2xdSe07KzLWxsrf9f+dG6LpRg+TcwP/GZVdBt8Rd7eSpJpibYpyz
tgIwZ6vZWulF3bANiizF2T/31xkl9vRFxsxZJ1mT5ZUy6ZVWPwGWSYcUx4uxyfBL
HW9lDXawWCzJ4iqdL/28SN4I7GD0Qe4IVtNKlJz6DSKEhJ6kZCgY4tfIjZk2JgNb
tD0rAyAPxxFELQx8jrOpjwNsoAH8958pbNA0AoIYaOp+UBUbW0/aA9V/8Rtp/+2b
DxtuGyMnzx/FlF9Tbryy6C55Y8LSdjtqZ2ziCTKs1Rl4BGVBulvTva9U3UlDMSgh
YGMrV1GcfGJpD5igRqZWZs7QKLAoFZ/4pKCwpUV9CPl0DiOuwgnwBPqiX11/Bm6o
rqPNbn5motrGYNsr+oxEbNr7bY6KpdDxH99t7lut76bcfnWObdpaMviJjwmiYKNq
IGY2RNRzow1wHbh9aHSk8R5UYxAdrF5gOpk6CWk7IP+8vbd2qGBfFdkhwLDOShtZ
C0WlnMDLKFbjBz4Ux38aCZz3nw+ZG8noNvcxeByW+SVqavqpQoh2QC0l7vfWte0V
qxPcav4i1toNstXuLohh7d51EV2fNp/TFyHZCQ4KLPYgBzfvQ0M7/JtrF8DR7vFN
epWlXNjRSNEcCysVrA8AEaeWmME9kX4hIUvGZC4SjD80OzjxYFFNlxq+kal/b+SV
NpuFabMgkynuQr8PqcEZC4BH3Y3DjUCUbIo1hCPCcO6YXyjiyXAZdC4WTWjXAnpF
AvAiB27EoX2Vn2ivZamDizCfxRoW2KJpDq0CePps/PjbiatRz3ev/Yn0lJgQ0I1/
Wc094/2Dj4OZxx/S836xZkYouG/4HxSypb+LwAErn/yi3ZmnfU811CMeSmEvcK0+
oQ512K77ckK/HISO08sMv45QEMZNsX8K8MqxqXvE36OCDi19fFybZuLcyZGi3Oom
3IDc/OFkWFi5+OyMJcO0ARoBkKgklFyNqPkK/dKjNYp9xs/qu0F3HSFnHkGPUO7c
VFI92vUwcqAIC9dLZtRktjIOlABz74bb2shq0JRuFe9+xtA2rnIXmpSMCzBB2wAS
XPFy4ljkG8TK0aFu2rBIcHgtGIszXBnwqryR7eIphQD26X7rTgayDeUPEGOi+y1I
hjXJmmLPL3RdSK5jiHfctMY6PEfOgN4ubZooF2xObO8ZsYaHk+Hrvf3dPtnQYKkq
UF8DQU1MKHyaF/a9pbmfBMzjjBbj59uWY1xMZwwe9RM5W8KVm0CxDKZpxFtRB9Vw
JMtkaJmsFI3KPD6fhSPxJuX9vt99uN2UgGexb1VVzEpIFnuxq1kk44YVNGRX0rZu
NOPy4tS5hqqaAcWoXT10dX0692HUeqsMG8igdI6tNg8hpEPUSeg1wtdPUAOVD/yc
HxavtMxRN0v9laIXQD179JF/J3Rvd5MDZzbPKS829CBiNyePzkZUKJnN2LfYMCJI
rk/k+4S83MPCBYAdQkUHUsw7L4dSirX3MXLbL53g0VhOExef5h9M6ti6gmuyhHcM
A3Uc+R1EPaaTLnICxkfpwoTAsBDbMU9E1i24BmtuJBx8xtB5zRmVzX9G4pIY9cIQ
ZuQdqTSbYEVL5bF+S+JgHrj/MrXiFsty/1o8NCoZ7rU+fsWJdPPPKqOncR899KDo
q2LGdBAYaQf+4lOFV3+7IIzSWZqxAWNquOMXAiW3C8N6e4IU/LqGJMT+TcDRJI2g
uWr6ibzDQnuxEwtS8jOMTjFLBpC0XKNVWd/7M93UlSFCi+HP+X3pHzXmJ/f8RFq/
JNs1xaVaDbMuQuZnLcUUGhNLkQgpvmzgILFjxSI8IQulkQO+d7O+WDSooAZHJte0
8Z/k6E+ih2aLjqc02ymwySEhjoeM1DbARJHXUy06WKJAP735aRiEdLc2eK9Num/n
c+X7c2Ci+j3PY26tUBC/7++nfmkxHyTHawiWoplY5Fk7saGIqkZ3Z30ghEMgXaZ8
LWIQsENp88ZaR+3m4uE3o6eTJqxqFHDqYN3eXIBmm7NhcRuKU/ddLAW7bKvV6FEW
q3M3D1yMfZp1SF/QB1lla+omYqXjNQ55+fKwXBkf7VDhwGhP42Bmf31Vww2V3wbg
57N6oDqeoBpfjDxu9w+RB3MPbDf/yw+W0EZaCCDkewlgtciqKh28Y1I+EOoiURiB
ws+eYTKfbmAWdDobHW6VLuxu4LJM1iZCmsrBV77GWVdh8hLJhZmrCIIgiSQv52qP
xpGn5m6KgSLcdvDR4Cg1qOxTbR7tbgipc3hIN3v1hNNkbjK5klbyV1pJf9+OO5pQ
FFIbCsdf27YaiGCboY9N4YiJeSrOdyn4oh4bGzYrcXrxc03NlI7lvMse6C7g0A6w
LuSI9F/DPPCKYLrmVqnPGIaxpJJo1mhsV9fC0z2T0mCc4x2EJFTAi+hnhqP19oi+
z2LuXbvWut+z5TCiQynB8G84D9UibSoYFmYtv4+aCyGs1i1+ScmZSjm0froNwoaZ
ehkrCNkIAXc01gsuDRdLQUlq3lPEPm7mPfGBfchJ8CJXQ5YfEhRLq+4aYL2TJD95
EEiiW2g2Ix+CMbjPTB7xNNBE9Q9hLgxH9CvGzEKnjjVzfqZzfl7f+MC4z8OTxOsU
12LgTUzXbgN/pInEIQMdEJtKaB5N/5X4fvus6NhhmnWeOTUwhbm9+9Dyv8WtOdQf
IfbDP8Dlt5YodzshBug5A73NYRIa6M2UEas3TlcwaiW0h1ZEiNyv6QgTjqOx61V8
e/6ADVKtdNTQ0oID85FAA9aaaPOMGfUUTzDbmhFp2dk9vihIha/YOFnnygaep1Lb
Enb5nFm8CzEOzvZ+wLNLY8qVQlnIsURCfH0U6r0gL6y2tpcxgoYKoOT/fHlIJwTu
1YC9gmXxhg5qVFLm79PkWKb24LwXJjl3h2lqJRXlYJgeBUBy0RyXoiimTSPVynoi
mLQ7/N2TEHNRozrz/ZCYYmmK1O5SH6MDFc+Hot+PjNK6WCMhC3SGwEZRCbcG2jKe
xt6X/GdATPKJ2V16NMKFe2zHMeyBl3pqj2+3JMHcut0gdueEbguXrIkF9Z4J5O9Y
e6Kk8nf3w6LnNc1oquRcfOeQTd0lCMVAMVf1+UuYRcPM+GOfzX/aj6WokteFBWa6
ftv2LYll0b1kOMZU0KoDcE06cK5r75MRy3GtmynZyPqWYZaJhzdi5EoJDv/7Xbj8
cRIMkLz1FotZ+D2/fePTrt5hzsFPaKKMXlleBFK5tPaQa7lBkhE6PyMgeLd5PwL9
sjgIwC6IavE48/fATfA8rNQPPOSiw+cM/h3jydzOvTOR1bvDDl/js0wIkXfHIqMw
Dpc18azdymUwvQBtL7X9jPwOJmM0P3kANAOigd0On10BzU0RQ9+4O3JB+WvoCrR2
/6pOJjt4u8Wy0+A1jDVW64ob4D676A/AADn4d4ngk5IdD8VSQg0mVQ5Yoe6OpHkS
cBOhXuIOuFJDR7k6tkI7G4tT8rFF9H6OCyqLubXgL6wFFR6wvjUIfHyY4l4XN0bz
awzSmgHN6kGwwDr1PLe4t3S/zkM/4TSVHOe5w4kdE1w1ufl/A2m/yK2sBqTws39d
cyzfkw3oRNaSi7YIH+Z6C1aRQDlMz5geTZJEce4Ci0/cYpvUl66bqlfiAWKioIY0
EjQyoPnWbht7n1UZuA8m9b6BzVJy0jxTfV1BptrKBhnsKrYTX64B35slhmkRWS4p
e/RKKTzcvCalW5dcU2Fs379cpUSLuJONSpmnfP/q72UIP3RMmrDJMyPtiPxIVvOj
ZIvZP1BgoI45QBeb1Vip+q+bLeI3X88u0np+ooP1PWG67zJ6HkkiTXfs0SwxSy9d
v6KSVfiqovgdGQ4ESMRHcZcztw8OZopCrkC+OAIWhH7098SgFcrrENioeCusQWGF
72BqjJbUU362a3rNI2kQeHXfdzkuEmXyoBBuJZF9dmnElmqyrR4MmTweuvljMJbC
OM02uBHh2Veoxdl8F1Lme4rgjqB0cvXS4VAHApVPw3e6IxLB7rHJxjiDPmNymYvf
efWy483N/kxUxNqEDMi0P/KfBTfTnEkFQogLj+36HmraApT9DRwF4BKqkCoqh9c/
nVFNvYzhtlqoKSrHSbKqqcxcHm4SwS8mIfQj5z7zXa+OJFZTZfFBJ+PWBn0Bc9MI
ThrTmjCrI1fmTKgr/ZHo4v6mIrAq2GkWBCkyMz6dBkrgO15QqdzR2aNEcuDbVnUS
R5wFsTJJqj0ABRPwmTIUANVWzto090EUP4+TMA+FD0CBMsV5dwCtE/3BS6TBU9xz
XSreLyQA+4SHLfACFj0QUHD9BVBQlps0aCTDw3gYX07B+aJMkVapb8KekR2PctWI
d5cfQ9gEGdcW2KQK30XYLHDycr6Lox5m5qdb8KDNWPe/aUL1DuwMhqiZvtz1b59Z
8azuJeaM1iyLLTQ/R8lbZxKO+BM8dgv/2JCxePJdWqpPspkXu1B9Gx/b69WJKHHe
ZQWRgqjj94AbgS60DkyVvRvCUrWJf2a0uMl/6QG43+l7DRuth2X4zkuUYssQzG78
sIuqL7K/KEUS6A8MgI0F4OiDBBxrW10yxHAfLFJrc0jQyHZH5HofLDHJNQgVuHq2
42JsRPMBq5kJO9nPWTj03rNiHYp4HF5IMdS0glTOnIxkuupk6JKy6NiteagcO4oH
LVklRymsR6CZcndBmdaXXuLdJiA21Wp+zmLCXgGaBRhQ1TRrNxJ0H1GeNwZScXw7
fV+DVZjyhCPXteduhvgXkkgchpw/qls3pHwFpgQ2hIRbmzgNBeRLnCZROvA4TYao
e3LvWnZFow6vQVxoaMpBeINZ21VxHSsmuXV8KS1B+4HA7q9WvOd9uLY0b/1ygdxH
kbXaiovyc8zfzLpGa2+zFIFqu1dohOHcIkwv1CRq+Y8RseV8khrbMjhFdskBC+h6
V/t18P1hIAoGOJUCec4N1ebmRD6WazIrk5vT8kHT//ysvBM0Nl/X0y9Kp9oCaK36
ys2ggZN6IccCAxpDDyHaF8oirFoX3oVwZNR3mGV+v4vJzb7PmqAPLDh6tJhDG4OM
T8mceCHSqV8rTVJE3UwX7EESpGofeKiDPuuxYc9+LnaqM2bZozkZraX6VC9BVP8Q
q+wsKn3sDpqO/QdEaT8YovX5MK6+Teg0JDIZpKWCVv7g1b3rz3IdONO5V6tjS4Bx
Tc/eIMyboLozvwO2Bo7YAtqxlfILX3OrsFoecGtH1b1640610gFccdcAmFPvMKY0
y3Vi2FJniNHTllKR2bmuzJ3NcfghEU8uCLJXrHsXgFE3mhhlLt8hZ0Kp+E1/LCt4
W3lqIEHCpMyPcsVySSOOhUPlust/bIl1EjRI7uwKLPRzggpWspMQz8xnNUT1Qd7d
kpbvHx4avLIb8cbb0hvN8hO2RuSUQ4GtkqOU1uLWfjt5mpcIROy7iDRLnmX5ehji
GpGuZx1OM8a2OG2Yp2Bf5rt/GWPQUKpCJ3bne36Fs6Qbjge1y+Q76YN+fv2xTgRE
sBZZjKwGDoT8Kr8a5IM2KKk0gpvLQdd5TaSehibkv03bzmsaPMoRw7cuynAUYjFN
oG0eamELFm4UnLhGyRFhUxAysAasSqtm0i7RC2y3Mbwxmjq+jGTGqVO0C3CUqYid
bogZw1IvjSFWcvacyA4axHa3MUtr9Okk6k3HBa56ydvkDDgsWvGHwi60/0oe0z3Y
ikvpn2UVPJX1cxXVLHRGkWYAqar6QN4h2Vik0rry8lZOp1PCJDRuF32RD4WCnYCl
9rQW+5nKe+wfo+d9PLUB292mN54TsDwAJjgt5JzjMo5viBHjFytTcp1cZ6CiBeLt
k6zp6YL6HRzRiGQGgNg7QUzV0NofjMTReSOsSnJaXLkdhwZH2KsFchp0h6KGNpXG
SqWxLp4NVz5QAl7mbQhYPV8UezRbHGA20qutJFt6wa85y9pTqeN8AAhUDRIozqwW
RBjaf1d6MWrB8iJlLszi1JkQjs2HUGLaYjeQlIoAbDnvqlXB9GGl8n2j8n6ZvL/r
bx2y6LeiR3SHOncHs6bGBSHqANbDlUtUspevwNtYx0xUHQ/pzaqZxHf1oNkHDwKd
R2illhcco90HBiMrvvx16MWvX1wozkkzNcn/ACXqkiIhitk0wWlqStW2RTToyhCD
2/l3CQAc0Cc/nSFLEcBEMiQyABtdwdZU/RnCk4Xgnf8YumUjmawID/7RWoJH9dya
Khk+v6vL42RejPel50nUqh4huNpHmDvnkQInI1dMyVhJsFL3qYqPgzAhSbfZKalP
eLvDqDkWqsISOuW8PPUvhlyovOf8cPZIoQm9JCFNlK3ov6MrBzwl47sGsI1ui+us
kPPKWQ7hosZJiZJzRBNfJIzI6vwR192PgvuHiIIjhGFVWpkF2deUMFb4R11MJyJd
HXGK+4kctRg9nSxh+TTL5FwZwc9PTdQeimgnjB/hydebzz97+poWq7rcevHodHVI
IxgT3RH2vNfSETWU3FkpV4BHfQLnliMz2xZPMEeiB95DmS/C5PXwC3MMtNhGM0Fp
w7UsnJhsDzfd6TJ02o2j2DrksHmndA3LxsGw9Sssnxa5r5ZqY0agzWLtEdbAIm6p
G6yKRsKFgryNsbqtyHBVjokhEUooKR1tw0n8CRIVkolGSAm24J7m1VWyUBlpNn9f
TdHfV10T16thEkQ4b0LfhdtuVAih1nyeUvGuglUJpXCSfyOcmntzUKCfnV5uxW3B
YT6DexrnV6SGIkUsFHdxrqtykHihC0t0KPK6FyoGTekat0ex3SI0atjOli3x+Xjd
V/Rt5NU8inPGz7vBEmG18lYJKcKGgKH6UcIJRBsGnqvBT+75Mn1g6FVcAPj4nGas
EQ9ueDv5FgBcxSXGRwG1phEgUpXmgsjQcIHerB4nTePvYOUjgPuzU/NUe+u2tKou
xKQk4oRZ3xLATRFlN30Dgp7V8M4IH17bp9kBBmTA+NPaqpc4qZf1bCJe6AncuKij
heasyf8D8nckhN28iyJfQS4+3yC1VPErLq0isjfJQr05pA83u+Vb73e7SkXWIjvm
ariaVYUmVvWP8NIU9bMv+yedqAUPk/BrFKHwCOgij5QkHTDlE0URveTblPS+y9Tm
RRLCclCkUGr72y9Eat+tJbiBOGCeXsv0zyLRIW3+2H2gnMj/OkXswxpW2hk7tgyJ
NMFqMgFEi6qky/+MPxjM8X4rP5kNvEUeGJmWL3wFrPWSd7vCh6TJSCFw8UTN5/f1
3WR7/IqVtbeOQswdYDowaVlfwnPu23jDuLimGW8hANoOadO8H4+nmCY3kEYYUEB9
TqEwODCppKu3kcAXuo9MhP+ce1buVbyaci7TUcbhkU4iv1lJvwiQ7+w5tS6uOthh
ECDk/m3jIItawhN7z90YdEQjnX5+6PWlW+5NVSKxNFFCSC+1VUrg8Bt3njzBsg+0
0wvQxfu2Qv2zfuB/drR+684ScVP93H0BpuSeTp3ZQaLc8jR2OPmReWPst5iEpUEl
0nBzbKXaO5FF3/tIPD7TG1EQ6/EXevyrDNtrYRpDXFkk/+Fe2WnwU3yOuwgS6z66
x2jNUKTLye3bhV+bnWc7M+QZ6vhADgCBFjCJaO/HqN1NRM+42fjXYQTeJod4xbdl
uKvtXevsoEaPOF9aS7rz0LNFBJi37cBiIYIO+RVG05mLOoAs7Iq8iA9i6w3H/4fc
sNrQ0arsHeN76sLUISb0Mr/9Kjwjqjb750XLTvxyAyXivgpwI0urHDvcgHsS2CQ9
SP3hF1PBDw9VCol4zeVxo03j82Tamcvl6K67AzzWRWKfoixoHN7oJHEs6yVZnfCL
dA0cHjzwPsbD/eZJADRoPCFaeO3dvmmm3L/7C9o/XaisjtC03fmKYpYeqlY+d9Px
6ptPt1a5HnAO/0FBbFRvUN1bpI9KCdIQv0dor/M4xfmDkpggGjmxKWT7aBXrvsfX
k05LxiHj+NxVaiNKE/XhBU9otff58934jvkUWPL43iRV8jGDhj/YS654ztR5i06W
Bz80lUrcDzGb5aJ97SHHd3E1StuaDwGcn8Vhjt8STmzxC+rTZKSxv0u0ea5kEgYk
gpZksoLmut+h6B3BY++Jhg0RTHF0w64qoRLw71jTZ1P8Cu1lciv4K9mOlOw/5Wzf
GzRJ1KNXdVtjbfEubhslba2SoohK7QtfrMqeqMFVGp3jE0qYyRgBOUrsoPL4l0st
Qf2+aa+hEmFjS79r72px7Xfrt6Aj64xxQg6ZAQHJpj6lA4IF+z5qaKoD2sW0UgeH
Fa6QcAOUm/gFOyxsx5UQv6pfyeVF5Ktjr8BKdjajNAhn+rEjkv5ImO0e/N5GCIOW
vyFrghhA9T5nsb7u8PvC/oZJWOcQjVQP5s1RGonKLKXisbEOY2PNM4ELvxPTrhrG
lxl0EixYGmebO3Rj713LraIFhx3h2wrvhgmp7rlaJesT577ZgYhe4/JXSzpOE0FB
PEm3QoQ8YbOZOUESR5hckG135YrSRtlewPd+2H//ORYlNPU1JFCOE1/0Jc/j+39S
tEgX4PdUW/512WeVGZ/aSuFSrmwfvqYpTGRxPRQBcQhA+rl5a1Brb+KR0IkTCLG7
crv8+kVd+zlg2gV46RyoKxHFH3fjQsWCmQ8uAiuyR1S+ViCXFzG0rbo0AnNM1OVn
OiW5h8mwsFpAVzCZGRfe+aqVehPSFvOyncBrOW+Y+ulKAkepDx4xDDvmGTiPvuSq
H/8fYNm6ap1CP8gwcwO6BeZGTx0EY73DUgP8h/lN6ZS4t5g0+gattDjtdhyQ2A9E
qLxZVYy+K1d1ZEuntPs7pnBHg0pR4gK01ISvxzeO0fGBN5rcWZPBqc92R7Khkr8h
6d2yY23mQUZSB0oFZRJFOmS+HoMJ5ufN7ezv7UZnz1ZW97oc+jGo7CUPTqTV+b5E
xSOH1yvfS8+shSoY3uEiwgxHADuaEnm9DJubiXe5FG2P1yb6xqjIxNgq4Ynym4pd
5C6bOu7YNstS5EoQLIOpg1yahQ8gNErvr0GPehuc3v3MdynHfnq6s5ztqYVJMFh5
0Cywx9L0uC11/EZX/MrcfgSNhM452/YzyZJY6FltO4fr9d8nLfcsRxTyStajCjth
SMFWYidBsO6ME65L3P8hXKpY/2GfDahAyrbKBNvrxc0gFmD46fgpnUkMP0DclMdm
pq0vv1ESburwvFMuk1v3YSEmJPJQp37L6DpAZejdLyQR3CZ9lfaw4bIH0hBK9KWG
xo6KchxAWLjOpcW3B7GxCdiwTRmwoETkkBOdPApyojh7LjsZTIiUM7ygoDppuyfO
RlI02XwZvH0NkiTF2Sxa1Kxlvw/1PdPa1kduEKvLmSOlSPe5AKr0lhkGnQ6+nb28
ZVB2/VP9AyLgQWE6Ugp//QHllbLufmE/+ndCaQo40t0tc9IigTnsmqK0q1XpmGdW
s2g3i3x5Zc3HF2eSINOMi1ioelnylXoMLC6ZPnu+K2wS4tJPYbMBG7hYwOsvDjN6
vkuN7wU9myAndDWyOccJJU87tH4ipZZhtfVvBDA+HPDd8MMthKwpWw+qkzsb/FbU
aoAAvSoOiqhXzXunr7o/QNI0L9DFZzMSXedrXT1D9KZIWSVsEUgb7NSDfzOWQ9bk
tIW/4XQNW390ZYOhU9CNMaTssEO5FgtwP5pV4Y7sUqaQYNlNnd76yVoY31gNd9MB
ey6cVEJSJdqd6o/VEynhmqtwlOrokto8RF0Z6H2IHIhZfuQg1oS2bqgTb5SjT5hd
S7s6tWRRe1STEO5D9Y95LcUfKcydqzOgUqfmg4bermSeA0DTHBzeDu18qoMCJAaZ
SD/QYZ5ntUjyQPduTw75OpnUYTHT1ZL7GumhO+gPW3LL3HG+OoFiPveLaq+npCQX
Ln7xLLFM15hD+NLNS6jT5yY3FvVomavzVQCfzB7MPxiNRuIljp+QZMp3YRhsVRiq
6GrKDqcsz84WIIHV5Y1R0BI3yq9MfDI+Fv8Qy7MYwWUCiXPHX/TDe1sBkUXNvQ2R
kveU9IOstR98tMdozgb8Kuvbz2QclaLjbJBEKxw0lgSls+/2VkB1MaZBDrPQYlgy
LSA+OuHqu090gapCr3jXPCk7alqkR5RMc0Zmn21FSZTb++dMnN5lvcGATuXisDFP
T2Rze9QU7SHno8ZHrblxhepBbyhS5ZXmikaCMnM3pIGR1d8VuG2u2NpPRnR0D9Dm
eEh7bAdmdoohhSXiy5OWaOfP1GiM/13XLimybjrJ21Zh6GYFucF4jhQRw6Dn2BVe
gKAUHQDKKv7hg47VPMw4ftdg7ZQAJn/BDTAw0qoFFjHwHMJTTqfnFs5FoIh+9wgm
ADvh4gamF3js4dmy9VNjXXe1oiE9h4Hv7m7xilPUbNEdgNfU2byZWb92Md//LRaC
09d5iZoz34AAeuz1l2LrmQBIMlOKBXksmTfJKmIslXNCxwnOzVgejOX45In6Ry94
zLXEamRIr3iviZfmPkzuxnYKbphI3s8lxtxiEu2pGXDMTTMtHXTkKJZ3+Sz2I/QY
9xMDhxvXK4ZiUC06m12J1lzGyN6KwwVtly1GDvz1Pc0bSd18qWIcTEFiNN2GiYG1
q39JgyKfYmceZ6YNoCRx9vSsEMTUi93sjsakQNtsJ2jdef3QRJnKFSigneLtq5t2
3GnGS+pxAAwap7fhLd4IUhoHNfgmMjC4SHgBoR2JYRMfulwXQd376GdTdOSzJDH8
l0hKWZeasamvpjQm5U7U1Df2X2vf+ZWvzoWXC9Wb/8P7t+gXd6U+0lhpsX0FTC+f
Wam9ywDERFROJ64Bof+8YhHWgsYyHrUeetHMa+Zw9ZriORoTudCCnDN5ThHF6HLb
HBkTvzGKDeYGb5CFLW/L9n6r149dA7rIjJ3oqZMWb3gHVSiha4aMj5hglGaY0Mx6
Y1R9Ii2pBcLgZjDZu6LweZEHzaFafi3XoM5JI33/ZK6WVkqC9TjJib+IQDnVBTQu
oOZ4q54r8udNyNYuhEOI5EqI8LMvE+CUgg8G3GwcMmVfVzNMBSp0mVY16N0fU1ri
xtkP/Mg6F+zu+8lYDY+1YxA7KxAE/kv9siua/tvEttM3/Ak80/CCtj89U9BdQzwu
OYrTzzzAuWo6fhl4R5DWW6D0bWJGjnKorWXJrWvagkxcxroLGgebw9Y6FSLlNcNZ
TWDo8sFD2xHBAvDobHxeFCuP/rcjcWktuH/GAOaC30MprTzOfU+BkBr42xaodpla
WgSRn9edFtVkTDpaaLzg/xY/e9GhCRcHZsE+u/zUVxig9hVevRFcVhZA1Q4T2TX/
xsvo46Psc8E2F2j52WyBsRVxPtmsY7hFU1aK3O0CyMFsR7G7FZNvRxgCSIT3srqO
0RdQ9tw4qT9GuhBp4iSmmlp1U75bpdQvLHth2SdMUL+U0au/LhNO2QKRo0NPJ2eN
8fa3vy9ecgzRbgwhyC+HOVvdtpjBrhUHi37QG6jIYIinGSzeDkYsMSBlEuVrZHFl
0CTZUNEpfaNVqUTd3vC/vmNbdyOCkEkQqcIqvvWSHf/BbG3aB5fCvSLoWf85Rn99
hra0RNAFXXSE/CfCrXCNEUJtKDdzTuQXOUiNONIcJG7IAaWiw9MBQVoLsT0kot4e
gUyPORKf8lFbciEeyOZQT91dzD48JDyUZ1ac6iYp+xANOqfq3Ri2wF++vO0AxKeP
9uYTxz7c31XBEQgzTeX2T0L6Lfr4AnSwZWtcFCYqSGKC8UiBXcoIXBvKhlebIaEP
/anjFfCzeGZDLXuqS57l/DqSQQNT9X6+eUTkzz7fTv4ovzzYcQZRUSHt2Q5zX9Ec
lyA8hA76O4KauL+Oz6t42SGUvPWmrDdqIU8kxLgOa0p+GXyAHAGnxbe5zeamRmZm
Tn10H+hdtvzcUhpEEACnRTELWN7mIH+9TNmK+yGRQozmwUmCrB1MPxOYLG654q0B
AzLb+/PUcSFr1Z7GrRpOWmfL52jqxZ5oJSQn9nrr06JAQUQdDkf5/5ALDP+2eE/+
GZsTnAjZ6S0qeoApkEECemOq/lef4mM23ffgNJphI7jBruYZcpbj5M8NkKwhEWZA
xmYSdGD5qJusUuy0BKv4+nfh1MhLXTAVTcuL6/zkgWpIbRxXHnOmLUSKP9wyvMZ5
am+Pv73FEe1k6Y3lLg6PUzhuoCKae1d2P/c5AdNN5DM+hnPZvb0tetreObOKSXah
5Zs9GoOhxcGS4EkZCgf+allYtnwbtESIykdzwwKWA1fcxyEK/C0mMgkHcUQfRTk9
26zuFxvDNJnkzr9ysWdqMsZVu9cbVRfjaYktGiVQ6LkgW+Gm6iDnqxVy7oZSMSn0
HWSKoHK7/UVZvb2SQ91mPpYpJYS6fOkA8gGu6g7F3ap1nfHVH0civxfgN9WWBPNb
ZDp+ubxTHY7kIJaf4mKEh172HOWGS9B/mN/Ff+7SshDiLrFOnu2yg602C2yUkRZP
krzBz77BR6PR1hLfCZ2GrWhN/sWChozgy868d+bkEOTn/YLRUAAeA/yziFN1BlE9
sew5UpkPfQljBlGJQMH7ISr5LXNqOZ2k2Ysu2RMD8gat93ug/ORMeFCgra2tznuk
6bD2G3QvKAXzTJX2TfoIz/pH6a7So/QfT9DSarNtx0iHvpyWGEHcQhIH+ZsAukED
rJAS/0+LHwUnAZ3sli9CNkydNLjIIsZ6h6FweYaGUsaRlRxXmlLNZjRm7rwb/615
TVBSN6xpEjzTPkCW8qFEhs6Yu8JctJ226fPFbTl4IBEqCyXwbeUaqamNGwYd2fBh
Iyd786CXqzSqlQfyYBruqM0tnr6reWXfZP+F6SuiL5Ao7CaZXkbQovVx7afMtOqB
lkzULhdusYBx57XEvS6yoTF3NlWTC741l7F9xZSgY0SsBS/9qCd/5zpL82XP94Lo
qZoHj8n3eAQ6ky0DB0QDW9p+DYzmpU4E5jmRjTna+AUjslTwZhX3t38GYXxEWbvY
MeG/++9fwReLWGVAhdn11NHV8pRYpqxRv2GpaPFiYpd4zW4lS4Y4M0FDKjO53aW1
SvABiehnyJ05zyZFbMiQnSUeB9YYpavXQYZKUrs2L9IVt7mEuEW0JM7g7cwtSwgD
s1nyDjzh6X6RyEo5FoSntAcjO9rYZAFxsTCea7/kgxXsmlBvV91tB/SktGvg6+Uq
xLkOtR/YC+Q9I9VYfL42v/Ch09NcTIPc5tRM2an31f6K1ein9W0JOvg+NyQakZOp
x2cG2CRGq/GG31F0Hua4x2ILFIZz0fh2JOIW7n9iSU15XciUHw5GGlsJCRAMvApD
3p4Yu3pDNU8DOtx0v7pll9Vw3itLN2H7KcQxpsEAOj82TGFFHL/v5sCh0e5Z58vv
GpL5w+JyDCYGLmvUVB2wJIAK9Oe23+teBf22UxFWipL+YD8pdVQPobOPLqtXcTHp
aT3kXoJJQbLnYwdiXU7JVOrFz8h9cjh7rP6KBHf+HP5QpEYae4Ee2jz4nfEaagb8
mpHWb9+CKl9QF5p/VrG043jvVgtjjFwukXhywL3lCggL//wz3UCP2ZCR4fXH+FmW
CA9i06Rjk4/bk/a8xca3aeyV/v7ZDAQuCLrZk6/og4BFM+YUt/uRqk44aMTDsRD7
ON0QSLtOUdrEdCFl3SEg7BHLGaZD/dErWFQqkpQH6pPeCjGkvVbNi7cmsr9ba3Iy
B/JRN/kMw6E7Sxzm8fMsZ8SGJPeVBDUXOfxChaqat3wM6yXIFYRxu5P6kygPwzgn
3d1vCIjCRJT/z9hdM09NHKhADJHVr7Rje/Dsv9ukbcCYXILVAvf41/v9xV6yHL5a
aE2PUKG3kumjJOH2kr4IyV0bTBXlmgigPkN4Wi4P8cw1W/nZNqdfw7OqE0tHlwuW
JNdRXs7OyIKPBbSBgIf8OoZSqqMMWBN2kUeYjhXnjJDH8jaYL4BYxJoKN1+KXXYl
9gj3hcSA92xmN2vuqajUvjbStEks61LvS5klZ3vLGoZkn9iZ82jNON7RfB/o0oA4
A6UCgWsnNbVjf+/JWMIHlxbUxhBkK2mxeZbHk+d1yRAZz1UPFBshgR2Ps3kA9ldp
KXe8if34lBVtCs0DjD7yVpn3RVVddYcugpeI1sZjdC6XeIwXv+mLlHOkLunKMusW
v0Dr6WBq3GuYUaBJwU0n8rYoZvIOXh1/RH5dJEc/2l5r1DLSMO9uRpi8r6pF40SS
jxX08Wg+yQXfjgH+VcVG2kgQ5N4JYMxF5f+rtX+2v+FWvw8dby9qtNpDU/a94w6H
vpW6ejCZe1qI6tMnDqjFaNdFzkbyCGPAOjAZcHUvH8MK8sOPOYoZaj+iCJYLJS1c
Uf8Ry/SHbtJSSvwV9pGZPd0fid8YiD+1EqW4SOUrbMkm8b4p8LIw7mf0qfea6Jj+
KepMYAsyA8+nMkDrnOqui6HBQNiJntIJoLW2KAm7JRKP3TFVvy2G9QwATfb/tv1O
TIB0vJYSu6GIY/8H1av0Vtgeo7jHu1sHEjy56yAU93GIlxlmQvL/oUishUcJUG8p
DjWrT/PynjWO4WJSnazZDvVl21xtvtUusb6BJH8Dw/wEVcdLL9yHtMS0fHQap2dN
BufwClMTWiOBF34Dg02IgcyBZnxTqEFNsSFqIUhlq39CetBWfohMhslXk6QDxPtb
9HbKgDNh5V9kE6xISy9HOxdrYi0R7/qbWioYSi7xWCEtJ1xLIvuplM2BDr7z2DiR
ysOTug566KLa2b3w/gBGInOhTybsYQ+unpxzwBFnsJw8AfZu9G/NZv3lQ4RiYsiK
h4Bz5wJWKILJzj4WaXOac3GccA8M2cqwY9gXirH+ZJL5EmnuLWcWWC+EweU0Jae4
XZ3TD7pyNLLgljS74Ny8jtBieNukBlVczF44TJ+r5YLbYidi9uuGEUN2IyXNAv2l
GJAgxJ3UlZKY5TgCac7t021LvQA685Znhnh8vksGYQELQRU6u83XGo+1kIBGnio/
5QOyRk8otBg5ylJ0t2ydq1Df68SucQfFEPSDbt5xCU9bdBVxc50Yh/V6sKUcUnpv
LsNfRaCS5owFs2gQmLj+CPixlKxR7Qq+FDoypCFiiB/zzWjg1lnSC7W0GmGWhiSI
Vc1K9Iup5seCAfqCUTj31jLWdCJkWcCLYgOtJT09QP+MJyEk+yGr4IrE8Pf/u4QQ
2dM8Z4z7jJKca0uHpgh8kCtFxs0J6m+fu8YW9qOpaavI7mGcBnlQW3JFFdjKCSQw
6infh3vm+edoTBZRErfLSCgDCVl6msDswT296hHpS+smpNYz8IY89nBGcpL2D+Zq
Se/LevDLmil7Hqif5cbluAbvgdITIMOuJpfLZNW/n4f6I4hInvs/cFBLiPZXgOF8
dq9gvtfcKm1jBaNOi+DwLuIlOioDd5npIpE+kvrUR3B/ltwNFXJn7xuoQQg4DJ7v
1R9LojXLGZjaScA3ukcCu/3WavOrqOu2WTeYzu5T+V0AeiEFYyA+Z8hDetnnPgHt
vLssaCqVDfoPmX7nzusTYyUqs7WiaqgHcXpfMyPSUlWWUlbSt6WdPryfHDNPdUR0
kDowy5T82o3M8g3K24kWBihdFCsgRIYdkk9rJnDtXGW4EUUARcA0soI9ayUOOCih
2faiKVmc/CfJPn8OHLMhHxSlaMJ/oeyzBvJpREKqXBcnDUxRJU2zdRRXbAjI+lo6
Wn5yNsURk5ARJkoreRGSqMZ02spt0my/QymSnvgzgzaM7XABa2PMOOY5aO3Uvxu+
qhYW8+Q3EFUKzF4b3qh3c/AKoR3YXRQqgOMRfWZe9NapBbVwsgsYdSqJyNPeUU6E
odPUnvz/yi7lqwFKzo3IKJ5wzdeDJYDw2FyAsZ7XhTRJ/Ttb7EcRs+I8svVnN9+U
vJ0tP79xMtQx0cu+5aubYqss8rtuNVthYMw1x7L8Y63KzrXh3HG1s5I5x5zH4Zln
IZyZfFzQJe73D8+eH1ddvURJznnxyIUd+9EPr4AW+QrNutGVCkYXoxi1KOTaQHQt
Lj8rgnMMSN7zANH/kC3yHvsicVd3uZMo6pEeu9juFdOQr/gLQ57ZFab0ZcZfU5jX
N9gw3BXz9XIZfvPHs8o54vyr1k202lsrSti3tky9XX3vmsPgctzmsh6hvBpdY6Bl
vhbx+p36kEc3xbe6dAyO6EnKBYfGoLlCPcYCEZIZdZAT5fBNVmfseWw02muU+quS
eo1tW/jMdjEv0ybG/I7hnJlQDNNJSSDlOXDn+dwsML7wEs7Uyge5BiB7knco3ICJ
kvNWel/UqCWE0rxlK3fiG8FMrf9wt+IPQ2XpDLvTTjBN+Ur942nzih4YcDxdHlui
X9civqogzi60M5TJNQ20RpwUlFX7u3ULxHvLMKJTim8ohvOVDL2dhHhe5BU8nYsp
2pz5vNMkwdhVPH3FWr+KykheBejOM3V1RKjxp7dKzZrkN69u9Q5xk4vPhgC6VbQj
ISaud61Eu4+L1bjTJZ5wtRaJrWMuG6fF2oaFEzl8l1wFbK3aazFTA6CkLLPXJMLG
xOaXVMQxtMYi08y1Pfqfh+3nxcScf+uwMQCW68O79H+kZvh0lPERnYn3AcCEANZ2
2pLBxMPhhUFdIuYnsQxw4mObHpzyikO8iu9Ebr8h/IiaDIZKfq0ty4G30wQ+XLq6
dHSowiV56tC4IKDGH5Z0LatUeC9swLTqbNbc+O0Ji/hhHWZ06pwyAse0jiCcyHaT
2/r+tB1SUglUiD92hsFCwJiz/oNSzJG7ccSHtDLJZwJwWgRns5lp7Djkm7s8JOC9
njvDvTJ7dkP1SgXU3ySTx4g27vc63Sfvq/FlqL7cC+RZzx9Zc3z+UdXqhARnaLqK
tcMxt5X4c6/qDk5icgobWXdrNdEDfGbHQZjw6KzxmfHn0Tt5QssYASvU4y7lIxOm
5Nsxbd5yYwUJ1rNGorduB0dJ01bqrYENrZnkGABQT4kkWYTW3Tk70xD2FMV49k4m
VHHALCy4wxM8QNKvuuOFuLR9ebFxtFy7MaYcIROAU+xPTMbBMDMaMYevACCv8oVO
F6Mlq9IWxLwTe/0IkdJ2JiYPZ9GlZN/pFq08SV5CRC/TerzLkEPgHshsFgvlQBUW
rxhxr4l5BZOyePdH+St0NDeNdksV92jVsUsJF5+dysYh05gURBCxU7jM8DinrLD4
gX7pZ7SD3FAtIDYuFF4+tJ/nyE+anGqWL4FoWbDui2qWQWXZKG65Sh7+mdf4MVcc
HkmEXLYJiS7ZkVtO1pXsAO01VOKjQKmqukMSgPXtAlRXpjerNe06PHwOzEsoGFz0
dMMUcL6v/e7Am1omSBzFayUm1ronBL/jFE4LnnRdx+sUk3Bdt+spy/XhzKUBfUov
TVSRHb0HisXCISVMvFNVp8aSoLinAbESwCXWMq51yP+E/DeD2u08bDuq1qlmQLvX
swLghYXUkuHbcBFws1woi+bHSAFHewXY+03Ewk8DwVRtLHJW3tZR9N4X80aXgvnX
VSS0ys8Qy24do7u+NTrIWTCNEt6oDzR5msMZ5nAc5ETLNj1WOmjCd9kt+lTLJZz8
zbACbUFTLfkAU0I3AYtsDy3BCak5l0rMYbfSPu5ndLd+12EhDEo7Aw6BT8MGz5vj
TvOVAL+4lCHtNz4BJPbncYYEsYntEswN15EEQXPiiLuNdKqSyttGi25l1A3Yz3Gf
g0L/T7fpWJN0P7iRiQ2Jcc5jTBjlUbwg+6QApCGnnRMw4FATWCSN9l822B5+Ejp8
2B3O6nuej8x8B6CAZBhVDLTKHmCnkgS0+wjdzQzqs6W1pvgEMowovi1ysOGtsWWf
OyLnmjaBrrGuWdVHvfm0JAcUxQ88l8INpTfGiEZNoe7s0HgQM4d0doCKpqN52uek
0g5TpYrrCUgHMVUJ24pcghIifAFfwbJwDSUVtACntYw4VZ1EnaQp5DDV5k5f/5mQ
mm1ZGllugG9iXEnE28RWOZYRrKLy5qhbcK0iOc0coRtv092Wd4pehEeubi7fvYE0
zcTUsrfnDOxcVIsONlxyz51WvTUlSVFCSDXIX6/5RrWpZZXPrThRlqc6nVARHbx0
nnu1+rG1Ow58rG0dbfmybJD++wre5s0U2RDGIGSCIHF18LWI/CW3uvRYgsWEWUzz
nWUhJtmzpn3sCae4fVyTY5TDExGjuuXABZJTlVuk+BsMZiaXzzWKJks37zIa+xZR
6q8T2+YTYkQetcBFWT/2WHcN9TXTXb9Yy4oN7xa1GjYgDEK+E11Nvji4/djbfsFc
NrRYUB7aP66qIcaT4G7fTlTQovwpHhcb0hXnLV9Jdm2120XxVApn/WWNCfslS7cd
nNUEtUVYN/2KT97qz+UdrWpXjhjc6updL6U1GbXYMWTzTzTo+zlE4akRgz+dUMsU
pEbnZarhcAhpbKYWMwPuS1ayhmN+xe8m9kY7ykICLVzsVtzGysGykWPcp57+gexO
cV06QCAefwx4WTQL/QjSLlWbmAUmBO8qAxS/N3RVPvwdmXLGx0ThtiLpN51K4MIR
/hymHnBAu7VLBwrDfkARiwlLyKbT7cQzHTGRGfrNWKLw/DM6qg5wMB37Yt6Ztn8H
n8xCEXYA7xIa1Ukd60p/MELdMrWV0Ubr15gHrX94W6T9pGehwi3SNvc1Zk8xMJ8t
SxDBZLmtFrvH38ryXhg5SHLt1mJ1xJ/aAV8IzNiqU/mmPjqjmAjKPlX2LkBnbSri
WlQayQsmX0Rh4BNYIni5zScz8mjeGZEQii0p5tW0ibBX4Gabei064mvnQZbfH3yw
y2YbScYXQ+aOqPVDXTE+EBNW935SKMkLP7TefooaPryKxM5QmAqB5Evtw9S1p8fJ
fKaapy63ILRlG2dyaHlS5+I6pvIj8BeF5aVCGUxD18Jdp+E8WmUk3SNFpyE44ET+
fxAh3QNT7Sc3ZlWAY6uQfTIJb0uekneZU+ssL7O5cYYhh97bqXoY/p2yy/GnMmt3
0e7kd0qWnUBvef2waHe6XbluFF2YbWX9dUSjaK4oSq1eW4/FgAYZTcZghLpiw1pL
UEicXBfYLVzLMPgCYsbsWyHTiSSXfybHKlC4sdhxGJjRuXVZRa3RNSYknXpVwwkw
acAmZGN6AP8o/0nCC/0hAfFyZKYarLS/9RaAWOE9kGdg+I4Kpm7pGUIAOpzjPh7Q
/sR7NX1umsayzxBQCVU20ZUHP9kBKAh5+/N6IkNDi1iWxpHx4E1rTS67Emks9AvE
7qOjPvtGsPJW2qzEmZLUsz8IkjokMg9TZ8RHGBU9kmKyEOELc0qoI4w1SQ2e3qWF
IFDluVU4zDqn1XPv4BzNIEW9AeBaRwY9Ng4Oi4jYNb5AYkQSMF2X5jYJsYpjWkNP
aEIksb2mUkhao3zeiDzVMlDr44Tt/ym5/iXcKbqlWUJpS17Y6WD5tx2c2Ip0mZgX
TNYHKIzQXCtwGGd/Gk0hxfFzueBRpWQBjCVxfz7DuRcaIZ7bshDSqkxPJfpEgttl
r+iHp0eQ8nEDljvVtBP79fIfcHoEtTNgIoy6oBF90nvwOY6xambDjrnrnKgw/u8z
15eLu8QWXTkPT8fjha14TPsa42vUNfTZK3SJR5bVy+IBtpbj813lQyDoeF2TRqOH
3SQgNzk9aQFe6ZgB0ErJa3lt1MIYl5InepW+bGBPDiN39srQbEgfnYetBuqlQsdu
tJvLcJjzBm5B8kM0ljfdL/aCVlu7i8ATCDcHH+IUs9vflVKFLQJ2E5AAtURWYeFS
TXMtnwVKEZninfQUDtVMSuXkFzGsR7wmezo+/y4QVtVp3LT+sHg20NUWHYYI1qb+
N53JNcpOr23Cdkn0zvblz+YWd6VhD+2bE5RVM/Q7I/tf4uJtZ7wVCY6YRKPy8du5
alFPMLxRbzv21mK5xIX98nkoTTT4Tb7mshQ6n+QX5PXqJEjSvwXzfc9LCM7UEffZ
YsXqsq9zboY71HTfejI7HRt58eikO1e65ylom254ZcAfE+zZkcUugdjpOBxaa+Tj
MgFJ5cWAVBY8SCQBQKjTrj2MyQlsx+OFwege5qHCmS1SLi8hEt+/6eJOUuDT/TB/
qRqmzkl7557qV/6hDOfSlQ+UYZMaJSc7Qb0FY6jPR2zN5qDrfODBLlCy5JJ7jNYK
8B4NYPTkykeDbgBGRKUncqIf6f/kluEmMvTEJWyDIR7qZOsks/6N3+sNDPg8olTP
NoHyxQwMG4zykqJ4KsC/d3j9nnOLc3S8ORuMrQSLrbvlW14Ovn6LjBAh3SwutqQ4
ialTmZPDH9R050FvvSemt2gaGqIx13RAnsTvX65NwiuvZXyu1sTGA8jmdp6xA5z8
QBiSqMtokRShdkbsXwV6BQc+AnmEVYrDwt4OOxyKUBgQE1WksKippvIK54cpvybd
mInKaXTA4dmpITe65tlnShJKiUEaTwSr1Ch1EYqOQxs5hEgAUiX5i0aAlZgV0yCv
RHQbOfNh2ABhgVej5/QuluwuxOATpfVsencMRKWgIRzY+dZypp5jYok1kNroV8zW
FBogKuC/4zEg+t0VdGbVjhYY+pasZLP0pIagl0y6s1fsC7v6Ue8lSmENvL8Nx7W/
tofTX+Rf56OBw83qtxbglDwk/32tiU6vgJjEdXg8QbWevlQF1Gg59aoVVMLudDDi
OcF/C0cYjnVi1xcPp2tFNesqDR5gdGKGs3viLfJvMvqUPPY8zawqpPFtCr4QyKyg
GvdzobhzNagO/Wci3bWsFjEO/LW2Mw2JAaTfjJgBWjnkoZe4XF+PeY1rvBLrwzc4
XMewrUH70qreE0xuVMWQCLW5gq2iZVEHAyXMLRZqLJOocq9iKmGXmBZ5LteSbCoa
9wdg1LpoW/TuoUeivkiUgYJSj6bfROwVC7EpMEgRy/NOXWj7n8ETgGn5RPCHIbY/
Oi5U0X27jbikohB+KYavWJ+S5O2OVuFSncjGwIG8PF3JXA8KkrmPuTntoAZ6DyEk
H6ZXgZ8MIuZrTrmC3dXPiBlp39H2MN5nOt6sEk9GSE6qWrgHL/N4PX8P9pnDZ67m
kdJindopo+VWISxvc9gSeDrU7WrPlXpQ5t/nDzrEQYtoFXEdN6YCTChjqh45rlmb
aHkykHLw9CMoF7ZzDCr7036gaAlEwPzcJ6qYsW7FtN/IQtqnd0b+J1QDMfpSxmli
3FVJCjDjpF0iw4KK//u6R+q8gBKO6lkjBj9GYO0GcKhwptYjp5asNrRlqyYdlZVn
7UAEamSa8AtS3gl/yEZRfnYB81GH92+OSQ+79wcBkf/QPJ2aRMsO+DPu4sawQHTJ
KofvB8bo4crfgCAaZl4FnGc/XELwMajh9b06OzrIw+imSeRz8e6rAsRt6hRtRznN
0sh9E4nduNhp0V7vsSuV3X6cibO2XroY2LcEfrvQ0BM+mFedWfvRwLdDIzxSeINw
07iXg/d2a0AetNBs7DKcA1VzXAdquGWZwFTPqC6HHeNfpzecoVlgXTYCD/XWdSx1
YuLlCiHyLeOp2B6HbOi0mKkpqhysQD3DqRYbMcCBKB+I7rFljQ+NhbUEwIrKwXBT
Dmb5yr/IJCFJkO9M0QCl1yDNGwgow5r0BNTXDO0ZHUlQfLT81HyEiXVT43mkEafr
CnG9RVFGtD80CJbbyib6JiO159YfvAA+cTZAQaM5mj6n+tuSn+jjVETOyebQnpFe
FHBUB28YzO5HOMT9c4HcLwLcZJvK1lApob7+K0PweSYOC+N4veNhEmR+QKNKBuXU
FdgbU/eRT6upG27RyoAKZ9fRH2lkg2XztSBTpfx+qctfE0mg4ZcQJWK4Mzwxtdkb
AMcW/2EztXonK4UzlCnGDNNHysYKCzKpA1mIQgS+neUw586t1twRImTwOzA7vmKu
WuRZlisVkB0RRiC/rrb/wfm/XsNN3XqTWoC6jiUPLxi/HPfwYCQeFjghHzBm0yEw
M1v0SaQzDS87MjAEJb0ljUKPvY8Vi1MqvDOtFqaFsPOZY+lgcFYNmDiJCEOCkfZ5
jn7QcswWd02KMYqRAJx7GAm3aEY8IpGJrMH/VYVzZ32erQjkGPekbBYMVH9z972X
nU/N0JZNQ1PXD9VME5fWGG3rWXGqf6LMRkL2pKaht4QXGZLCWHT/kkwTWwXM4Isv
wXB40fxdMomVyosFIJN0Yelw+YSkMxtWm3+Zbm6IWDtJAFzUy2ReUMXjBgsjboNI
dpHCUBp25s6RWmDBKFqUOafeqrBB3B2ybaaKyMs5b8nV6koK7M71wXh4bNVu+AUW
6mcVXss0dHknYVALrdVN4bGyi635TgHrKyxLggXE+7Szw1n8+eNm1jkkbnjgAI3s
nPGbLA3UHrkUQJ263XU40Mxrll/PoRAZ9HwZnVfqpoO1RN9I4o2PhBB1a7lHaBEQ
FX0eIbuE+U9jYqyGveXkPLu16A2dzd86gMG8aRfPHBmhOERb69xG4aayB3X74D+L
iC2RYBNMMj75smZpuKrVa1TSzBjULndkCE4+mHdbSk1wszjBcp+Ae8VW2f9IhQE4
fCVBB3n6gupmEGNGPahbf1bQEwzbXygEtCImS0BrS64R3Oj9NOssL4zUXKicJYfI
IzELh7qKG8tR64Xoe7BjVsM9PHnu8KdGbfMkKD8ZtulwiPySUkAnne67GfRKxaMu
zNM/hWvA91q1hueKELOuMD2O5XwFnTDmhD2f8mp7WPLgPlzEZVInYKbB7H52s4gl
PXdaML6IQXQqmWfL8B60Af33/ZdicMAGN8YPuzVFhGQJiKU4VzSupEttUOhJB0ik
65LM39qKFq+YbFsdXuYNhIqRFppEFVvdb8Ch746I4dPF8Yyf3Cmdi4TrNfQ5BXgS
jv8DxhlzvnkKp6AwCIRTq/tOkXaDsPRY2wOQb9sY+fXR7NTSqAl5t1zmd10MwseN
tkafuSqdfI2FALagaah9Kuh+wEIJ4R7Ri6LQdjuVuwE+m6C4UebhwcE5rufilzeh
lpiWZ2LPa+0GCMQB4gTHoTzFivBACDd1ukfpjad2MAyJMG8tKmURoj6Zhh8GwK9+
CwhyuPx9bsQTmMVXmcs1i64ISwmGChPOuQfr6UpprbqkHr6ZOBUJR0Cp9cZxtJrB
1X6dDkDIiM92lroLPZWr2OLBmJBwlL7wy045qYYLec26hkKuk12b+c453gdUy2Jl
Ztv6p5r+9Pt6Uu2LokdtwvKOxOn7xOV2VESBB7SE2XfOXDdSwRac0b87G69mj3Qf
3AR5wj5M+dzeEfhhtxNStIsEToToU/3DKC9MLXRMCchI2b3cWU0isen79wuzO0vt
N5T3FucJdxKLcyz5n6srVehKpT0TTvgTRDkQ5+C36RXhNcoYHHKHTs3hk1yTF3R/
/Kqxh/aWLN6ZEwDHLb+FWILDt3GodHRbgta3oNBRdpjzg/sbkk+nKN/aFjvbFS8B
J2rAJCtOzZiCTa9S8un5VIyx2hk5qCRO7QyNO+HQ05ARwi11M4j4xp0dauOW/FLv
301JeNXIsR8kYSHvCRtZLSt2qXv+5EDolcH4taSHge1V9KPztUxglbh4gKvqLcB3
yLjboXPhybT4uzcfs9P7OZtT1NgM83htevmcCXrj6jsiNNfz3KcKVcRawooE8Cfa
vVgPLWqZI0US8uZ/muX3MV0HNa9sI7aYSdLSTKwsY8HdMSF/xK6JuYJAsr0lMkkC
Og1WlG5HHvhftylKyiNFYJ0RrW6Al5PCnj5P5lWm2toJxF7hFXIvBtnHgymJN5Sr
aEY7hrKi7sGvb0gMAcAObrqBbITlibFe8Fr9sJQ6cz06LcIV0UNN7uTMnAh0WYRA
SkO/EtOrjtGyVYmdgGTG1WutieCQhmc7/BhLfcEZJo534J986Yp6xUxefPJiuBS2
9lOfEnMWRHBkm88rq+sNjJjRBtlgk/DpI725Gz2/FWTfsNf9tL2sllv448653+s4
K1kMJmnhEFABqLkdy9ewDFXFr0a04ISJ8LxpY2+1C4rM146RmWxoYWIMYpBtxquk
EZkqr7wV5JWtPbX9BPIrglPzjzbQvstIqiJ1IAKTLoK17/q9ACRVTchJGHxPUykp
f4pmfTLoZ9uLe84bCO2+OOW8dCc1ApJ6Vbeat9svSr8hnoqe3dCpSnkAbYujxPfe
ho0RFrc3tOr0nJpVFwPy/5pGaSmQpVcVtg8zliID2n7Q2fIpBTe7GeZW26H6SF5V
mkUu3/M4IZBmq9xDp7whUfoEPAwfOjU2qHZP4QE1wBKzG5ltfm+BVRcdd7E+BOEP
p38cUx0PlKLn2IQwuTzXMkxeflIxpH2RXDmTO8tE3EMYuDyZOIxuKi2/3QUPeoHi
YFHcgQtfsObAsuIZHJWLwB1G4YS1Ius8S9+0Zyrnz8433JKfUqPnL8vzQquZYtBG
AbGzzCEr2uApVL6n601qtIfpLixYoKakS4XyAoWyGtOMJBsNIRQTbEsDxP9rwfSM
mXK2cjqStVHlxZuB8BgjWDIJEtgFuiQU+my3i4WIVFQczTgqpnkjYf5qvO+1Vpkw
yr7GVrWN6m24YPhZl6nrOZxEBfJNbL3s6QKfH4hlmLbQPjFsdlHtripiOwdCngyf
n85/LkWeW/8BIx6BdK5ypb48XM0XRao/qx4mHABt0POu0/KL0p3SMD2iE2iwC5WJ
TQ2sFVrRIdQjQvq1Ege8VB63CvX2SBzRmSeLS3/YZ27qGjmZ83wzvsx1J+tqp6SQ
tEVi9VwyfOOGJZAASN1c+pDdBbELHZDa101cKpjFIEPFH0TSL5XqCEX0GQfu0wzb
khgJ3sTV44Mg8Yd/I7QC/rzsmMN/VcSfYJWu+KZ2D9vNO2WByPjMomvJytbPDaNA
aCp1vv6df/gvmPzZ9mTg8pWijmm/nmEnrwm2XoqWYt3iUAPQuCZqGvWHI/X3ICfn
6+jtQ8Zy3xTcOoFIv53wprZ10f8KZF8cJaYqxZrHfCKrYkolGR22sAkR1rxciDVe
jKtORlUZZVW0V4PXjYMHKz7ggHzPlHrYTNrViNNXmfgUHnjhUsxsO8gEl04dfch/
yLP+XLZs5HrqQlYljlImIibxwCYZeEDXNbmwzDSwpbGb+sR+QB+DYjyAN2czuIqE
yOLhUxLzzjDMrDVaD/TiXyEaIi1lZ+RwkWcMg//l80Imu4dyd6glcE1kKmUvDQru
ysManqBAknDmTPpImclkuPzkeApVUrzJlgZUX1l1z66WFUfPMRp/cnVuQCq2/5Lo
bNFoelvtHWgexy1l0bNKHs26JeRalw6uGZbl8hUVzwR0VoQRP8V+Pbe/Hbm9/Xpb
IVcu7+n14c6ofwK4jcHvZqFLIa6f35Sj9yRa6lfsdKRVafCJG9cCnKqaFwOIdQEi
QDqqd5iCx+Mkf7gA6UUgF4QfKRhcAuyppsZqx46ckuogkS8h3Dzc0zI5RvrCzM/x
5AKow+JoBD+o42qpUhtnmt79JkTNig52BcjB34sDcxpjC+z604+LLOGWRQdG5NEf
YXjh0o2Ll8ETYc9xN/Dia8zE8I0fp6IL4v7D7tDSls45meaRuzfF3txjjsb3cAzj
ttbAEnmm8Hk6PKmzjeAtyVOQRIMWUpgFgLxRvLwdMyLTKInpwVAQ6JmLbtCih87O
AaMlah/YlTSVgK8NwLU5xQIe66glWD6zDH8lqVHB4H0nOqNMTIGV/soL725BAayx
NhnyoJgF0nvuVVyQI7wE/hsowBHVF353Y9UfslRtCuBY94TSqIPXA/ZP3Ah1jX0d
3oObl+izPLA5G51JQztIr+hvtWUYleu1OCn37q12WyoRSxdJd22y9ArZp19t13RF
v+qPpwJ3k8Ul4gst9c0GXJlkf0OTC80Uu20YkGlhz5a5qeKixM3OD6CAI1G5Ruf9
eQg0FqteRjPryuFEtgeT55xjpuAMmtkPtOicNBXN8Fcis+Izu6TUFLPss6bjJCU5
nj2dFHlMVpUVE5iOMaDkX8NnY3VYDpfWudLQ4j4RmWGZuwbuGg4UUerunjgBAfhA
roHixPApU1SnFRkuTwqTWz4QYbhU0HaVUaGnIf1USiVc8SWU0UxDhpddJ9KsaR/c
x4tL9sv8+cN1OSKF7HBEzyR9j0cHo6iyvbB70h36QgYNYb7qiVYCrqdYRxSw4EY5
c6L1i7cdCm9LY9Pt3/RktER5juO5kAN79V5TaiWW8LqdXN4WRNXuUIEA/OGMhdfG
agrXX5pCf8G8XetERJKypAHOR0JVp+c7vMqIqUCCp6gGRVUQKPmpL9rerQu9fW7v
mx4Ej+0+WfEItAFehdAQIM+OZk21UttQlgeKTFExUrYe+ErQ/dtN4ufTJLY283fr
vbZMvTgjGngLkDF0il6FHq/A7xDtBpuPvzU3DqiPkdtKgj5jKo5B3d0u2ml5XA6D
qRP58rtoKLWzg6AQOa4UTXukVHCibixWcreJU+oq2qUgx/igblcZOLarpAWll9Ws
AdtfHJIwsCcGyhFnCTeahhogRktYLYyKsGZiKhBZQxMOiveBiXZkJYexxJf3QUjf
yCqyrN7Rp29JBZFU0/FwoaVBHa0bdD1E3T91ha82OND3P8yLSACctqesDR4Itt8K
q108wu8c0h/2Slzirwn4OA4c5xwWI7J+1hw7npLvpSgTeduSs6l5fCXvGSqzdlPQ
CltGgVuSh434HNsJLmf/BkoxsbR8eX2b627vQk9hz8rrU3LicfoluwlaYTefnBFx
Hnncb613S1aQa4/ThcT84pelEH9ZZJeS5uBdz8N0KgzZ0gkDhwwhqVgKiNcbXy/r
2stNraKAbz6jcte02GcM7FI16QtBt6HYKnECu/jVHyeWK/syoGR/De84oI96Beu4
ZJa5p+7ZGoPdup4r4FtsSrFzV/n68T/9yM5wmQvFuoLI+QJxcn+SBy+ma42kPTWf
NybhBo+/yEyLofT+nKMm9wcZ9RiyIssxVAvEARLW2ZTaLjMQuIPGyNU8pEhjzvq0
xpkymk3HumOMRuZB0z/Jci4FiIaM/12HphjQqBTvYJFzNrXwzmR1V4OHpxATVhGF
qNKhaUeaMI03YrbrEUtqKyciI9q6HdPXbOxVTuUVBrbFFn0CzwxYovMMgffYLgM2
54Ys37J9V+J0phDSuowS1TKpbj3sGFLZnZgGHdbtfRbC4DSLhv17LIbAgcpIJjSN
3bPapy5fNhELe2xsW5w/XVUz86f2VOJqF+FYS3z8aZTj4wL08Kbed3VXOAttp4qq
Xp4ogAuQQdVH6l4x5zr9a/aQnHS35DUgs1kHcb5vx+5ipsHWujv6+z4CJa1MChPg
JXxTrwizH7xwTJR8PRybIR5Rm927grhlu+LkOUqvDAwM8QbpokakYvE6zrVAOZ6p
cvWdvlWMzrVPmgXLe4jzn4rKxKqgOhUBr5Xb/a5uL7cfch9OxqWLrWnDMGpuqsTq
jju+v87zaL7yjK3N1Fv2e4QFe/c8vw8bs8RbRm7Vds92cqh14r8Efm7buul6kPAE
rDCdTbUK4CUZWRpAoEmz4MGHRTOHjXOloioTY/0Cg5qkL5Gnpp4qz6Z3nXV8oYy4
KbybeX1wyaaDAt0FrgrmdyUSqff+sOR96wZj5GlUlI0tHrGkCBc/flwhNx1LQ1Bn
Q/TitOPUc6vQTQqOpf4zsDOHgSCao7EtkBrxBF/UVpegrtAzQQoxVYn5fxKLfLpb
DweQNJVU/ctzLqimnpCRzZqGKJbmAkKkJelKLTfw3yZaqooEvi8pR2MvLO06wuFr
qm98aRKK3MK9j+YLKZgZNXgX4oLivDAhvVv0+f9f7L69AQi6chRU92/+xg6w5OeU
IO/iCKg3rYvkVt4mWqhzq/+c8B7Yr2Mb2YrpoHbpwDLWbaHmNXXleadfWUfRLCF+
pxH8YYwClLmyInD6th+E5+mVr1rT+OMI0Zx4ItpHoOseSToiPUL7nD1eDD5f5DPH
z5M/Di+y4FYdlXhptv/o1krMxnQG00D1nvkuEKFGkc+MH3/DS5zOivD2GZGL4qGB
1FV1nC2/hKUAUeXe3TgdheJ1Odu9K/PwPdu+mCmRlbe9Bh7AbTkrOg+Y62IruBex
gFmsWOoO1hYJYzclvaznaun7+5anhvhWpC0mkqxWm/5W8oQp2QXTlMS3ivA1ILjo
XQHnodg9IF9cG2tVqu2oAxHZoI3N5fI9rXz0J0Uf5x6llibL3CeOBQBxQc9cvl6B
0uPG/OQiOejud9iwVf0Y7HdRYt93yQ7Q9zU4UPJxSF/DTJetiOCBnosO9EX2So2V
zh9iFZUJfNfuFkDL8mJMawu9wustT1bLP8sbDNPRYJD5HKdWnPVsBZdR5e5dW5nu
0TbVJlZVQq73+3SZAZMYjPc+LTB+v0bvHUQOPF5bCWPg3TlnOMjWWM/je9QX41if
fNd7Nk6NYEGlKnYQHs+ItOfLfIevs7XSZtCdV7JV3C5BdCQEGCIFkA3LlRrAA3Z6
dzAHzO0TG4qoC3VJzvoyB4ruYIfhEve4AArFgbb57dH7aF4i1Ms0D6AYkJyMfL35
CwJ+MASZr7qbwsR8YPYxpXyPDaoevO5ae09G9FRggSRZRoxMGo7+il9s3KSPFgdf
VfxevNb5JyXjn6koE++v19EiwffPwA4/uznKmPNYKsokqXUrObLSl9hD9V7Hj6Ym
AS+e1RzqUjYrrYK2bFSNcoEvFFLJAQIJb/nCJ6T/LMzJ1AyJzRtU6Zq8Mev0aa6s
M+GyGtyo73Wf8oL4v0K3413xCJQH9PwmbVugPzC315RzutQhc5KdqOwkN1j6rXDD
CAnTmUpbI45kPS7JbdZRTWAcIlM9huSpZeIuKvVutvHcNCT6Sw0UGRnuUluugVuq
gTinftC2zmW/BC6k9mVKZIu3h+sKhooKJ2a8hZhkZctbt17NxiIEBO4SNRda1les
6LRSH3O+LmgDs0XYyEl3J2N+BHuKKm9gsq02TMFkpeTuBEpMbgJyY3JGz6pyXlZh
+2Lb0GDzwWapdaXcKwpXwt43GVE4ZUTJUni1TGYblsdWzCNxrjDjvHriFZHccdrC
oaLBEs6sPlSsahFdgkhrLVx35hI4Sd8+OgrDEx1l+ZmSX7+9JpLRwK/FAQq+uIaM
I6IPAqVM7KyBAhc3hpHEoWqywV7MV9VdPH5gtrAePylwV/GwchWzxuQcLiasdees
l5wxQR89mJCoRRIkpxY62VFyqhq4crnmSx8VnbSGqzhO44OuUOtMEMa9ja6969HV
jiHQJGW1xdOqBXyvelSHW0f/GEqdk/IisMOaBEdndi6FCVukycGyFNBkW7YUojVw
gchQ+uuxZepD2GPs6yqIRkmGXjrJdTbxmlPCb7FQN44rmv0Vi/IJro6wrbylbr/w
cC5aGdWZt0ry/Aron0dYv+s2LPBKYRQaASJoRuLbhfnYtaaBrWtLz2yGzHXMv1lA
E+a0qLjSpo6A1LDmE9eycTcPLBJ9pMQeH4AYQm7oskUFRwODiD0W8cJhosSr9iIp
B8odImEZzoVUq928BYgImrljhlRhpYsE0jafJs55kIDT9UdO7wtkIxHhjiYFnwzT
z5Gf8Gin6yJKP8snUVLmUH2NLV6Qy+67+LNLrK7J9UmiwsxKO//MOOVCsRJBvOT7
/C3uPIus8LiRtbJy2GbLwEQ46mopcqGCXQEq7dolmUb3a0HVExXxFYgszmIpYWe3
t/HQZS+9R0lZcIGy8apon3x13Q9RBUFwoZ5AJ26RuWXNSjykVEVWrL2Q/rofw5UA
5TkHXPGfx6jnTu1o/jlbMR162spm83mQ4n05rBVciQQDkX2tilqHaqqtr6wtfi5r
72TtdjQdxrrFX+El1Hls3uOdHChiUlVK5SjJ77y7vzql5riBJR3OnsofLSJ358Zh
Dev8C5w9liSxBkMhdB+yPCrW1oz+OpBdHoR2nHpg29R8RKK8IEX7EBt0PHVrFSD4
U+oA+TxIM53UU/XB0m3NrC3Yu/MOPBs1qZj+64LWF4us1/LjJmguuVEGj9Rc8NLf
ToyLoZ1aDAIk7X2PYehQ4cH/+ac7dZ+dEQogdy0ov5Tuzhy0EWYzWOqhhNO8Qwo1
i5TUe7GT4NMPQycgGww9GrwinnkK/xc9caOAvGOuIcp3RFj6UFZSryHNEHN7K64+
IncFuO+jxGCz3+o1Bt6TpKClJj3UW5jjMdjLZnRXeH6dC9vgoNGhSvk/d0/C3tCo
h4eIre+7yGjXsEDKmZM36Yzjn6v3jaSOKs24DyIaH00nxa2d2ZzHhqchT3ATRiT4
w9SywyFM5eZrHo4p3hWB8GJn/CTlJcMHzPDmRE02OcYeKcTp6bQUGS16QzavkU9/
Utioa7sBkP5wkQfhmF7E8wmzORTGbJU99lPAdRz4eV1d17OfGpXDIpK8HpKUwc4y
dyeldzh/douHDc4bQXcDbk7Lr1ehOCcGsmKMPR04FKFliiyh/7W6hXSjRRLa1O75
IOU2lz8V6G4XiIRcdvxhQr0E8V6bt9FoSkpy/eupzW8Vd/yDyPsXfw9RxijtA7hX
dZEtop4r4HzlJ/KZ9IR8a/voR/eZzJN6CUnDkuNEo6FzKEXKyFpYvN/82G0j7keR
vytkmIdpMcL5UW0Ki9UgDhRbVlON0N5g+4Jj/RUdsbPMhOrKVPWnIi0kU3Tuf+i1
BR2gq2JXrDvmN+bBPjN4/EoYWc0a1jR4OHNRZXMVcFgKAZJeduICwLQVVsKNhOUu
K+30ODagwk+5HJrNYZ4Q8+rJxHF+oS2BKMTfTrnsziR8x9kehVEWnZF4XDOQEoh6
fheFmlR4SjUCALSrGT5WDD37hotAoz8qjqn/y0Kk/iKaKMQukC00arLDz0gMs06W
rw4mWUnWeg9v3Zibh0xcpOcGq4CgYJQEMVccdu+NIwu5W860q7pDpDcowqOT+Aud
ST3uCEjjwdjt0mUUumyIpdC2z3Hj2BZa1s7FOXs+l83Sw53WfvsKZW9zoM2YgCMS
Fv7zzUpGUV6VwxN8t/Uyj0Y271ip080ouUGu5XH/aPlJuLGlzlYhXz2mndcaPG1Y
JfnIFsPWTSiZi+Myq8LxN9+LD7eefhwNMnNa2zwAG0/sTDpd0VRBsFGTTBQzmbaL
bxbwLPMNiGmVRwXRzwxRrPlXeJFe4v+zhVyJmd1sLoouzVzOijt9UtyMy1vbG1TV
/wTQKsy5Iw9PaJLPjA3Y/TdINb7+plOtUABlC1Uw5WEFY5E43URyDuLaw2YGd7wb
hfrcKoqY8n3u0nYrnhoR/zmwI2CQm93xwoHtTqsTvzzMN5M3hFX9j+4ke7bEee3G
QUg77XFL24TqdXuDLZW5E/nrjwJUGfx2yeHnlnizsNhkTz5eSuek0E4zV+7xd59B
uKOSzr1VKTMTXohRXNq444rUyXa3RvKIrJKRG+o4uzbHSsw1wH6gI090/HDGdtR3
BU7BwpMHnUX5tTMTDAvj12ApOTg/haGoR8DmE8ja/bDhQWpObjo3T+nF2vMKalAT
ptfLiyoUGat40OUw2MBD+7Bcr8WLrec5kRuzqJVBWEZX6zHp7uDOb8YjwcNLydym
5s6Gyhtlp1X4oDcpdmT76Y0cz2BNudi0R7FDSppQhUKgyAQw4iSjiOCJaQp1IRRj
db8Uo74m2hVp9Ig4pi7rUeSolvHDyHOyzM+6Ub0eFjwEecEBuGMiEI8NAtD/WQ7c
8Ecrh5mGJTv2I8X1eD4gTAng0jtI8OHcbDQLAms4hbECj1WTCfDDiIbVIFpkcE+7
XUCFKuO2LutoG47VRu6ftZMek/3ER1q7IdhjNLhEdcilLPswtS66DbLXe/AOyZrO
7inWUTESBjKZeQbJkhun363EYukJ0K2xQIhlXs8cPtI504k38UZqdB4dqk3G9pcu
Hp8b1YAAInCTMZnUtbHLNqNVBbWrzCJGbPZZ2igg6Hhb70K6m8/Nx0QB0Ba5U+xj
AaZvvjOykxKYLN9Be2UWuqeXSG3p/roD1c7cWpgz+57uUVWwYXG3piMKQ4CZ8ozO
TQuYIshHHyHyrwYAI/E5O3Lr/cD4ncOZbCbipq9JHCf5FaR57R1UiB1C8Kqc1gIt
UJcFGd+L6Z4yJkaNGviQpIzhIw+/1d3vsELXePBvIGB4g0oTGg6whb3TLrak5UgN
hFvq5jk9Ub2bRg6g9gFhYfhdMIpYH7YSLjGkWfPWocfiegaEmUjclzhfnsFNSp/+
X1ysvSZEE6EqDJysYGmF628BB5TaMOND06qfcYOMM2P0nOyBH3itgC6GOsVWhJFM
POPsz7uOEpp6sfdS0g9TEzabuogtC/VnNGEr+Mw64P0P0d1zG8tjhyHUB+V2lhwV
vXcLO3M1qoyrPTf4xxrKS15Rxw5Y67R2Ulo4dTmla4rhBhQ8K+QO/EEC6t9SCYL3
Y/eAcldsv2R9/IyAuScMdZ7CcDE9dQ+S9PlIsQS/2rJSIfBFsdcpXDlPmTJcym0l
9m6l3zDd60FhPTciG7iKfoBiGVC0cMQHbs3SI5fFsjmfCN4Yn9mxb6SvNk5pPwNE
E3QoZivQwyCH+VHPou/zLz3Qahr8gKY1RylykeTybuejHecm+7eb+235azm/3FXs
i2q/u68xdOHn7HU+mdHothpWgzDnrwGnfmLrs0+FYd7kl0bmyCcRbo/AUE4IkN9I
JcuW/LAZ0CinxCbS4UVoeqrdCAw/TAjvwhGW2ld7DRm0kFYv+mi1OPHuJV/cGpA+
nuDj8fYnFdyjzy504KGbayIfRYDEYfV/cGN9JX8EQx5bvIOZHej/edw4wjS3JnxO
khXNLAqvx43/K26/qFE6Jv4A48E0/wWjHGPGbZKWPGnQHX++jqolXoyZvzgb6Piv
cIoGVW1K6TOtngZYeeA7PLhPo+YOOUqqZKBX2wbyHZOhYqLBunguYBBQ/8zqI7DV
+hQveB9YogW639O+DLqNnGLrsr9/mZO4xKQdTm93JOvoMS7ZC4MVqz4CXNTYtxa6
RgE6xq6/lVlB0V73hohRsImPdkqZM9V7Ba72UCpi0c/cicSJuBkTN8tEy4q6E/Fc
8R/GTnh6nTfSqia3kL3zrIqrKamuVJwaQUHdOzMbAoTZLQWHp/ivyofr3EOil/mJ
lm0aLJTRRLnoZGa7jrfNPcclft/OjyDE9Ce10dsZ3CVszlfCWm3t4xnJVbLsfv7S
sR8DssOHxCPvsmKUz5/NqsQ3bEtFUIi/HY1wUCsLDpzGIiIClgMUvkUQFneW2p8J
ZbUY4KScFa3bvQjazLBjfgdw6P9Rpcrncc7fxiBC/4Swf85dhanFgmcjqSVYOy5h
etueGoz9YiMEeKjhUCG+T9IvZ1N9tSzsB6UaRBIAlz2wvFqxR3SBHQo6T3k5HmLG
aXSIv3fxfrt4GyQLTK1qEIk7VYI//YCidyDkxx1U3vE5YZt2xYSVsobeaSFz6KXo
T0HcgZvZfCDcQnWjjkrHTKPu8QYqw72oyf4uoBV4V3Atp1O0n5qOcsZJM/TmHd84
zzMv1XsSfqfGShrO6ZuUy5z2SZg9y5xVl0YdDCdCsnFMhte3tX0Fz9R+7FkNby6t
1G/FXtUtTlQQH0txVCkzjrkBo85OhHmJ1EVbw2QNq527prsQhSyE1TlfTBHkJWIj
w4oufbVqnvngpoOIbjM8pxGViLHdfGUtjjbrbvWehzBZSvZ0XBGBnx+F39THkWFD
hFjpWrn2FZIGGUhFMKlFl2NlXtJYerb3VO/UiYrvmgdy0fakvRPMeqAC0wQbqkMI
oDzFKz5Utaq89Jp/r4qk13XHnh/uyyqBfW5dlbvTOvJNE7WcEGf1FZ90hAd4/G8+
Ebm6k9fBGkXLKCiHK04mpsmP8kxjD93fzg/ONlQZQ0peGPMXpWgEIYg4XJTVXMn+
XNb0hh397nbhlm1MQDPL05OWA6zS0iVTZVvqu3/HTR2ZDHs2zC8E43ZSaE3Qb4q8
U950Gc6jAkSiBzUuDFdT/L/4FCvfrGK4cbJVzsboT4ZvWBwaYekqZPb83GpdhAoD
bjAalSJ4w0ggy/6B4msbecqbfYOeIPULaK/c88KdMkAiIl1qcvGenF9jTUOZb6Yh
NoIzgkQWvU+ZAbxVc9HYxZh8nG2Iuv2PEFWOrDse/gYOHM86J5kgNNHfMpWskalB
CvtO8/9EygpSgGkmLxDS0j6HCXwk3VEhhKtnTSc4Y6Omy0oca0jm0jQw4OgJNgyG
xnoKWDJUehmP/5VazLMGS5FcN4TbTx+BLsRgmt3H3SmqCZYn7saDlc9cyq7oD75O
AKhvq5gdaERo4Sd0HBnMcWYTkUmZMATdvknNE4VLUEYlx0LBjoSAphso6xTqCtSL
O5E60hSjldhhh8V2jMl5xMXmFZk53lcJeztxoilY6WLxoTKthiPfQELCFLMZyOxr
2ZhUWxSbr8/TXCoIW2mtlpOqCZ6esE8Bex19FdLozOOsP/Ed5nR6jsrXTVkQ4rs3
NDlvghtOvo7ubVHU0VsNFOWyyOiIi0bHAEFa7cbipXGXmuhLk0UMEghQsFzvKnPx
BJQ7jSsaxXgLQFWAtQ2BQ78SYhUdavJiNc7PzvGDjyvWIqbEXsOehtTH6BxT1r+x
RRQQgDVDQT30deoE8Z7W/w6SocuNIxb9LRLE377v4SciRVWi0s7XWbK4auqYxv/c
xJZn/73giuNX8mS0el6I2+VzZPIaHHJW0ElE+liV/jpZEZRt+g1+QiezQUc9iY7e
z2uW478/byku7eNbUsRUp0Q/Jfk86IoFelA+KbbO7hPBVXpnLoWEC9Mpk0t+Vec3
TFqtEynxKvjBOgN6CKxdxswiGWvKmHqKeLbmWduciT5o0rapPecvWe3MWO9sbBZx
eiJVkdTJ60HwmZfEphNrzTVR1317vZwgE4BofnKFX3nQk4SjR5MC8wtIOV4p1bOk
gqB/Aj9B4TparaFNlN7AyvaGu5gypjEgqlglHtX3LLMpWnJHIYMCFeyqPh6yexSj
W3Y9vcFYqteVfSmg0VUx+iqkZwVGANsfgcmoEePFNP30dB2mW4NNghsUfpsGFUIq
pq/GlY3jTwVWElDeWaESZa5ML3xeEkNTGwgRnbOcGAtulrV7wsu0bP4Rn86lnOIU
N7X3vXVLCi/wL07bG+KGtO+0ZGZPrpWc343WjqO97s2cja0y6sf6OT2uhHlzG4UG
2BBbC1OYMqr0oltM4kww0kzaMgWGvhPeI2Bd5GIiztC4pBrggREs+LEWh61gyavy
6/mxRVeh/9KASU7Jp499blJOuFYSQCstD6oD40/Gdj3pGXkZBLxH8ENGyeBlJOd7
PhSLnywJJt7DtxRTxw6KRXY6h6X+yPjcv3sk7gO9oH7q9n3DYD9AYrL+kg2aBf9Z
kyFJe+AHeSGT3GrmVarZx3qb6g4AAvowSLPf7IvR5deTXDG/44xlvVYRzZUY3lRp
+bFyFBEJbk6MRdQg0EdGV6sUTBpNVvzuZu4w452XdyGVs9/7frMgF6KF5q/iUpZX
WewSTFvcMtDtyk84bDd0dUiC3dJwHykM2fUqKzpfrA+pd7e7tcJeQHEq5p6myx33
6lmVHeL7VRqp4o3TZ3Yp5shJUbAzikz2ZDty2u09U2tkai1wOwikszGhAbJwCrrT
hOdyg6gBguTK55t5ymk8OioKFAEQTYkmMijT3gDaOsBoFA/l9Qkhe73TOTLrQWad
4shylI41eu+N7U/sy7DBDapYOj+k2BPBnXl/FEhR7mQ6ZodTP9zpu0rb3MqiBsf/
gy+NkFzFl3xuWHlB9CWdo88jty8cVyBmNPOajabczDP9vs1a/jvy7TMb0K5CMD1M
9+tye8yefJB/9EJLbtZmVUIctHe0g+VGOdHuS7qRZ0etkjF6HdFp/cY/AjClZ3Ar
FOv9Q5zX6IJtBHFeb+IvYQeOVVOKtwd4VbvkVTCPUTnsqQKZNH9sEO6Tjzc1dbJS
VHC5YgxCoFtCL3xZhXbsVT+jQq5kxeh06lI7O1CL7zDgR5RycWia6dZjlifoBXAH
4nsXrWp6bVH0O7fT6jv1Q73LE3rYMuacL5QumDDxqPq2v8PPUFAj0I1ys1XEFZL0
goTUk7rNNszWpoYvfnJmwoKVoTbHeFcXpL31HARX5LK2yLjD9At/FfQRxwS5pV+n
eOIjzs+1WmZaetMsykq/Bx3LpytlHuI3T8knICTfyGcIBSz4Ljjtbt4FMVPOTKIy
AaWef09+28Si84ELMQRXIAjHSDOx4JHMajkD4EAJnLRDobJ1wq6Ad+zgHVr6J0Lv
/USciPACqCPEyu4qEP9vceBv2s+iZvJt6eryhJdobP2G19aZ74KXqKAHmBqEG2bO
G9M6c3w4YwQz8C4RvifKpzr8am+wbYEZEr5/CZ4aiYgzt+nM8H23asBIhUjlcm8b
diKgGzb8YOZlzTe6IfsMdBjxUXSogBBiqBFYJWjEDf1pfv/xKmujB4UTXmo3hWSY
WAcGtTl6dR4GlvdgxUkIe6S7iCXjj6EEvILg1trWxZl29bJw3qf23LwC60EqejFY
Nb4b7hWk838p2g6ClNOYHVGG3nSt0kH2+ry6MiBSx3txS+2mpPbtE3OAU6FqlUfk
MxlrkXHpRmzrsScYQFQnRNxq0AzSexhU+PAX0SDL7IB0qXcisqdkyrO66mq+mOlZ
4DRmcPmzNnueaWEhS4pjV4jUGj80rESA6GO2rrYR5p7Ugs7zxOXN0cnPRyYlJbM4
xd+z6ryK93/EP+AHebaAO9Jd4CPDu/uYHBuOSIJjLsRnf6N0UQv4s1hFxx+JDqAy
NWEXGJrBY7TxzpVJB4W1th6NDKjGZzp9NZ/jFjalBQ6VBi8k25N4cYXQ1WXquGsQ
zewk+ya9BrhO+5V0IX0F2JbazrW8HMsOzYrc00eNA8IuepgzOhkpA1MKCVDYtuAf
qDBn4+v+YxQcCh7EyeVRrORDOwuSeSGFYDOAXAzbEhD9CuIzRfnc5QoQVuMuMHgZ
rbwzrMcAfOng9nBmAJtEt+BmGiiQ51N/UGZxlhULm1OXv//1xDIs9QA9LjLaWV1H
Vf1LLUpfu10CSZFGbogS/sUezPIL4TMwf6v6fHBPZcOZREbJ4rP+ZV6N2oJFUz+/
DckyLRrVmHITnRqKwoK0G65f/XxjLb9yge+rqgA74A8qsa1uBZfTbjH/qqnhC50t
2+sbr/eU+82+5cF9QYd4Qj4F9IJ7Znc6kYgFCcMvnf0W5l6W00eiKC6PO/tLIFMc
wuHpmgGI0VB/GiehDPgGA8o2AsyV5HnkH00gn8fVXdWUSxMwbZBZqf6sN9QlzLYp
PE9SYIyyQA+z4XvDZ4OTYBBLq5LuBNWFuF0byO33lnYx4MJi0xY9HM/2HgNEH9nX
QmidJ2HwpZfp4epB/SgYTyesChkAmNPhEOv8tXLRDeiMhoKPuZVbMHlxy1+Dvimp
yqigKkPrftFQXAVOsv50QWqKutxktCmkpwEdi1NYAyKVOwgc7e/Ceiub++oVxGFp
Jl7JaEqhzg8hfQ+xdwR7nUXGBh2rvOUywBtVYnFtViYHs995UHVmdYNEAYOjWY3q
T/nzkH4Yfo3hd2WNKSWIt8pPUvc6/QyztsZ8o7UHBGT7Z8SAAUo3Ts6xVKWi8V/V
me19lcLRW35E+T4kJ2fWLNasceQIX8ZBlj4XGDaGe++Fk1OZWf7toRWIHdRfMg+b
GLyeDRyBgGJfgeYaMdgnevxmfZ5pBvabAZwO3/9waY2wna7cA7gV0ZMp4toKpJq4
5Q5B2BYqQBZ+lwh65v0g0GwFzETIrniooXxZzOXNJ+Gv57wvl4HNeWZe42ZN5HhN
FeOwe8GW3e+r+YGx23z69dFIRA7WREI9tf4c8FODVoeoZgiZc9nalYJu6DonN8yb
mOj0a5gj9PJRGF/kEKZjZUCWUiRTetIr2nMVntojIboZW2lGY94Bl8PxDoa5q1YB
h5D8w+kW2bD4DBg4casgS/Z7bYg+cvCVks3aQgFwBkzfz6Sat3rjo5hgF/c9ASvv
elwwhdSNIgkpYqvxovCw3wUUgvvkp8tuCHS3p3zcaUkG2g5mCthcIG0R02tElcme
FSJoHGVCUaVDEdb+EHeaQs0vcVjvVSBxirJa24ctg65nCdl8LGvWeEF+g6CR70wY
unSgBgPiHct0wVZL/DdtgKcobj94tEL8aZXRSAN7svdB/sXl540fV4Qlgvv4yQu6
LBtXkybpB1alaIKsVr4/faLBPXLU08t2W8KR9XPH69hbrFvCZvJKF2mfds6leIo6
QfRwszwZIuKqsE2TYMDG2ZNrvhUJc9yAyQHYbV3CwQu5C8XUoAOAejOlvr6sT0i6
0Kj/pYvLu5Yl/TaBKjvbAJtMWNJd3cKB6XMPcYfnxEoYPkjyhWKj1WSHnLe/LxVd
OtO5KFgKqOs4E+XVrjrkEhzv67bUnxmXwwMbDe9qrR8T6br4iisjZ8Oq1jvTOvOI
ZIDFftzYV5fhEsMWwVunOvcwzZgajfjF9IE2vlppsHwd8Oubs8YRlcqbFsMfwuNb
1jISbC2rYCupu1ZgBrCbawv3KWbb2M1sDh0x7jbjFZMGLccRcMLYviptU0IBko5U
PV/Rlp5sOfXNuCzuKWP7m+uXmKYMtu1mjTGacrEOunbCplLj+kOQXma5eDEjTPNa
+3b+rUl6ov3fZ9SSHqeECTbJO9a5vNTQH3pXTI4YTyMYUhAcZ2B0mJV3NWEgY7cl
2LGHPGR7b+LLK6uIdgalaKdMqU3u7W/oAqy02b+wP938UGTrp8SN8E9EwfDPiHcP
Qr9HkuY7W+jajFlwjsWm38o/k0BcXSy/X4Br8f6slxf2Ts1QimlffTyYfTTAhqer
0nTkmjXEkD2t/VRsYhUPg07UKyrz716V/U4gn9C0iPFIr1PlhEzPlLvUX/zi0jxW
nCFXFea3QrlxyGY2/qk+dxQ8qnfJc0xdku5fAbnWfttIWpmVFOCfct1NWlJIhCHQ
y4vy5fUXXPbGpKTfiyB+X84AepZbK/s+l8E6OXAOVvBlcodzatH2fKAbnBu6wTP5
h1paZjg0eDeNdXdG2BKP8hWSoVZ1mHbZdGemDgyPaeE/FezYbm+zhabUWgVska/r
8rR5ZDg8VNSgfjve2f5Z4HpSnUNXFoEB0gFSPS0jLS795cYNOS1j/pt7TstQ7C7+
CF8LImhGewBAyOEQzY/daJP7O4XXFBA0doITS5iHzbxvUJCmuK1ckBsnbUxTE96o
i9fVH+jYgTTIBqRYW7Z2qgr5UpD4nlwySVHy+cfvfBopLBgu/Xx3rY7z4Dw85Sjv
cjFBU7DIWWM8iikE1TXI3i3xN6kYtRTw8ny6AoQtoLBYakSMB+V0znNSlEUNfpnE
lOSNMHITCkPi9hPx+bc4+A+orjJfiW1kZzL8VHFUzwW3b3KyjweldBktLegl7/np
EVBkFvuuxz8dPD5UiE2IsdaXXtLPkMk98/fP7/UtEMlvFozhMh30myd9tZfpZLJI
hkiU8LnM3Pe2d2ZS45r6At381zUOezfhXWx/4GGEVm1HhIp5ioe5zghXYazJICfJ
Jw8tIOa78XkYYcUuHx+x9MTfSqlhG+M2RPfBMyHmHCS9ou1ILu1yu0DQ9Ey/+HkO
H9s+tMmOZ82u4d06S21pZvA8pmSq+G4heyuq09N/7ND08QU/Mbg8jWwncGzkrZIs
EhuzK1l/hX2xGICEiGUDMxXHOrhr91QUWFa/MPJVtKeybl4NKLj5Zigxu7OrF6jw
RkEbXytEtDyOe+aAf84LMS1RUQeGBiRP9Fsr8pOKud8qsHGcqOfNx1UU+Rb0BJBB
ClmGU+PQ5Wavp/P3kFEHdECyXYlNO2Yl+P124qPdGVmQEG+TBPtSQ6qBjnALOlzH
/etKSBOusNW1uRaWnf5zKp19T1capiU6J79YigiQmKDIZUBLhV5Q6iEUV2lYz4AT
NYYmfk2ogQhdSZFQ5vwVm5bIjE1PCINd3dixQjiBmuDA68kj1F1WUKRXXE5zHbtQ
fbjE1LLstGL7eijSz7hbE44+boAr9UdrOUbad2C08kFxqe98w+qnYpg4D7Nxicdf
RW7P8KfLuc6g3TRER3n+weYT/SBzD6jjt6MsaAHJqE4/89f9d8nfblQUeCuHsGjl
o7CJCFQe6jd23f0siIXwNY8vS1Z3k83EYcYdJ6PKA1mmBzIHBWLnFvdj0bmrEOsb
J+DKWcZ61/enYN/ptaJkainlUFEpjM8j4MjmWAolpjsqgJ6Dhg/rS6yWAoV3oiaU
hAzJG9ss9WxNDEK6PIA/Ibrjyj+5ErMKsf3z/vNKtYhEoCvHwRtBOi2NIni25Aoy
9hPKrAl9RBIynUu7qVOkD2GXWUjuM9ea2UG9E6WYV2a3rfjrNNqx98x1x7gqNB8A
MMlFEOH1ksxcPYo3G5Kl3BdeOBZux4FF9UpSlk3J6GpwMGQZwezml1HRBna1c+wn
86aMcmNQiOPtd6z0tPOcEf8YCbF6Eje+/YqAOqalLIz6Yhi7tVB7VEdbgnv75jSu
5oQGsQ1l3j6pAlSA7tWL3MK/LBweAAkCZLAj8loelNoIcitt4424qePLQ/GXs91v
A7XuEpmHtgARfdqsvvOY4/JU35u1+y3yuwIEhCb5rUOqV2jyKaKxTh0mTWhuPGas
kayo1dBZ5J+Xk9W1mTFl6inZeCZ6VP21gjyjHrCtI7/k/0CF+h5rtOHTu0p2srex
68wINO1U36R6VbRKdb1/dgGCsucooc8BQ7EkTMOTnjfn7v9nOXDBpjET4gueyMhS
+P/2bpVff6q6P5YCz1v6xzqH2vQVWPhlAuDuzUYrQtivXX3+VP7/+hsZptm6cR4b
QJjxug7t1KkQh2RNpWvy0z3Zzj5SjrqEBPx78a3IhhA3NW1dBdHB8SY4GeC1svL9
zxpZFIpys8/QFNpcAWEkvtgXT8W15g0Dl5ZhD5TCLnAusXhEK+nz/5P6I98C7i32
YwyupxD0kUMruEYFB1sBTxzvprqzda1iCXB1SWcyJCmrAjWciXEHSfrsPDs0s63M
zHP5yz5AiOg5Qw/tlxuPiRiwrPohBXpT61lvA3A1/3SnVuPl/qo6K3NbnsL4V6kV
DwL8RbMAkocM22YW73bW8qEQB50RzPm9niq/c5kIXm16lR6FYEl8w3e5MXHOe/Cu
jHHSXFHL3FCwJ9cy01p8J2ePcFeKl4Z8DBOyVGE+tlA+3KDk4G9mv7qfz7/iWcxM
FmZ85mxR+LbqsFfCwnBuORVVuQK8nkbAzJXTN6m03PQ1t4DHZzAGhYUDm9W4J20N
B30J6v1Q7x4O0PRaGF7hDegIucr4ETkOw/lsWB8TQAwQDZLVgKNWfxElLyECi+JF
iyKO5CAwo6SjSDiXHXGD/Y4N52Up9wXKLTDfwZFwofyZdNxxT0HO7lJiAQPN8X4Q
DLCNLpXJLI+DbeajiZBa+wm5NbcvCb1CGKSayNsTp9WxVWRQzIctladYDqw3EfdI
GpzRdrDjBHuy70XEhd9qOFXJaPH0QfAQrale5tadd8ulkskaR8UIaw6LEFWCZ+mJ
vOTn/PYycsFgJSTWZxzPRBvwK7sXxQ4C3QSwP5IEJi9LJL7POMhMLYSzfXPoYjm+
JH13MDGwSSsgC6SfHdEVS1e8m0WEsrpWg29C9AyGj5wnNZwm3/PnmS9PyptWd/E1
iU52GIAPbwr6/KcuSAN4Yj/Qp1ywfMP03GXQJedYqLNTm131dnCUsRKkTulruu54
MTNi4JFIqCQOsgAtrHmkzmM6L8uVhJM0jMr0Xz+29aNFTSz8OQ9UCK3Mxd5U4chK
/laUdSPy/nT43wf5TuKyFtCFWuv2K1ptWmvN56/pd9vaEuMVIzVbXvNZIFoHJRmQ
m/sFBu7slTS6yHI1+sQTVJ4fa4VWZvSS5+ZxLYhHriV4vnH+fl2tZlbUNPHWiFIv
WKchP0D+J5K9RFNsRtMZhaYri9lUALjFzQN6iKnkXxfb6MEPBfYwfkslvYSoMREl
mNY7EshQsUQSmQMYBaQ4P0bIkp9aAJXVg9zFI0yvvtcXJmx5l13gtdj2g+bjWo5/
mglbQPEUgIYH3x6CvlHmxqEYDwxeeQWV0h+0NOIcvoDv7nymLy3n94mmwVOPTGcN
8phd/ZTOYGlXuVdrdNCS3ALu7iMkor5pcopXf4ZTDYrU9IWDDWmEPGw5NZZkZfBL
TOkSAjc127N9DbAd7a9CRm2U7qQTjgHDr8xLM5Gv+mGvHA5kdi75SwKyruO/NJ84
bW9zbnZ7wgl9c5jU4QnlG9jO80lKllpKfqi7qR5avfChjCUeVCYSKbZnQ0r60QBx
eX5d6mpCq9jadWhW+oGEcvmrsNtMokj4QJKdw9DoavS7HhMYw+o8h4PWPuXRhlgC
BjZr9/WeNt0mC2gcQz3doBpnMAO66C8S9sJqPJ38/WSTYCOuzrBQu97mgUkCP3TY
Y8fPHYWwOhlz6qUaE7r8DqLhyA5Xu42ZejKFG5sMmjiyzohGUPvARnwXt36DaAJ2
9P9nD/W/JotdjzFQBIRYDlCQBWnWa68PkXB7phMzR58XMaoO8P6W04THqRtFxL9L
Ct0WICse/XBMfFr/FGSElhodgpjIw8p/rVaIhlY/CQIKDPuWppOrAy66DpPxt2pe
mbgmxfh97A/y2w3G3j5NIYyLVgbm1wVhDsyGeUlEyBQgTSN44zyXJvvyjhOBYgn2
abN1JXv9Pa3Ek5ojbNEQUbJRTFygPYsVANj8x2harQGy77+IuLZYzY8n59FyqQGI
olDbfewHou4swaYn3B1FCZn8UVmsDnLjkMGraLHqiDrWxjRn6pV1xgOzzJBdVmDT
kuEQWaZ8XsKdVEPpPbhu8spPcS0FOL9d63Nrh0Ud0X076zmzedm6HdeOKvPpa4hL
QyQkM3HFH46GpRMBCoxNE/8eGqcjxdJTyrfjdhq+Hc4K+qmL/YYWFY1tws7kLFOV
jXwaMU8CDDkp2kCkdOI9QnWfb6UVWKEot6bXd1/UBX4jcQuDMtBg5hXh560RlmD+
XZeZuxjfX0EJuuTNrfb47aNdCnF3ssODRffFRKOUGSj2lbB604x8BmgcRGeJVOK0
HLObg+L3iwcf2vHntIG9KH+CJSCn6EMwjtAP+Ff7qM2+vRMat60oOKgSemmqRJd5
59UoV8xIRr5SpZ3Gz4OuVY1Wk5k8Ozy71KLgI8VSkjrITooEgJfBbnJFiYYeRBMr
fx6Gkkl+RAaHtH9nC/yqT2iuTMbqRCCYiDkDXY4VsJQFnjYeQogBH3L17Axa7Y0y
QrfZBl4NyGOUlG2jeh2XTkKNDCu/e4TTqQCHmMv7eT/9QoO2XG4Wi9yzyzYa6Qea
nh4/5VW+rUNCl13wY0fdu5R1oi9o2mf23PsNFr/i3lfFhYaseXUVByS8B4Kj81iK
YuBMAG5YFz/oaYMnGGzmMg/YEzeIwL9oQj+sxNfIjeGsAd8RJhb9srF7msWqkrz/
SOI4y8h+B+F4lwLXuJxs1LyeFSMQasxe5l+x6OaRgXi1X9r5VvufD3c/mOqVIexW
guy8duuI9p2c7Lv63DvDJ5yLqzcNSfFYCULfPGEFmfk7VwCg0aIIg7CvTdsy3yYy
0kWBSF88WjQRxzmne5sYUy0O+fWhocr0KDvPHBfhbs+IDNxogR8iNfHkWRpuyDSr
T1O3/mHNaNQLI/SGTv6hqAS5WFW0Z36OoNVPFfwjkw5ewDAlwnvhpgToQHiIEdA6
E23LoIavUJNOztr1+gyntI4/OG5DXLc8syecAqd+qqQyzqLuVXlyGkI0iR7rZ+fq
vUMScNjblhHwpSO4d4jMSN7KJ4j9FN3x8ZpoEdaozRURlbjO8wT1WnsRjLLwQoky
xRa0mRYWuvO+oR++vvf74DRX/IDvTzlSv2ZY8n1W/zQ7z37a55sK4nRdqJzg9jPq
9RWi8CUQ/C3/dxuyrRlyg1Nd9QywBDjMIUeJ46AzySeXsl3GI+uzS4ECdexwZ0mw
aH/SDhWov+9Hg1a3yYSxNgtc2K8HTsZavR237XeCGwCKAJWTwZvXBbuQLcLYLQWX
vH/0xd6yY75gjKIA8yskIZVQhlOMitAUCuuUgVSAjYP8IqbSaCt8MZ6rEY/WLRZv
A4q8ILhGkr7cCLid6QtwRxf2kfNM7bW04Vcv4YaUizZKhMn6+5uWf0SjDpc/1ZAS
FtfGhTG6SfCY8+GhEaJ4WtxI/cEFrasdyIUgvZRpYWP9Ksrzs1A6UgTGKzSTLTgx
mhSoKHNhVdCbyw8qD+eAEkNFBu+U8qSNY11Boz79lpF990YIb2Bxr4M55aEeNA61
oBXO6mGGOo0iqk+/zu5RCK7uWknqf6MGuQUPqmn6leKcNf4TC4H1NsN3Q2oVpgTk
cIYS3/qEM8tqdyL7cQDrrRHQshWDJd4crXD0wkkf8/VbPLSewXGFtmcTByXAn/Sp
px+Gn6HwBPPDN1c99RTines6VleNvooAXeTHS8v/Mdx21QY+Y23yZWUi//rLxMeE
zPy4oNeWFXzto15RUrpZN/N3M1v8E+HV8TCKX1uozVtPTXgIsJaV3YbOkUUC9ozL
Xo0HJtpZoX4sXNc348LUpp55Jp2/k8VmIxpW5jnRCN00ffDAgWCAQv1JnxqI/VgK
VRKUnqRqQ88aJMQ94+d0dU/mgdrxpnB9OXMTDqh8IIjlxG1sgnvXp3GZFppzy38Y
ubGtA3nIB2cPgeKxG9p2F9aOa1gBBd+tl5mBsdFXYFyoiiMsOWhEjiFXA3lG5G9H
jRpQMl2mDErZdPUaEay2Spp9AHPSbg6qnkiAves8qfuUASCXPuMmkE41S89XV53E
hIWE9qaZeKdIJfvD/+3gDVYVc8ZLO0v8HOnXZnmu3MsUlSP8lvds21gpCSwjWvWj
+ITdjMeMrgcuCMXoLFlA9qh+soopga5HKz2ieIAsdW9i9sYjyT3qvGblpDbbzkJD
IJI+e3uY8LZVi3yZ1S0ibIvwcKO1VoMiMp7manfxLjKTEgU0kpwhVB7e8Bgt2aYe
AqKugV1QRvXHu+Ee8mCttv9qchza1xUha/c0q+dhcU8rrJR0gT2ZX1iQ2oKzODnN
rGuTUCsvBte+Q8iFDOttREvAG2QzcCHLMSMgMtYLESM53cfkufC+hKU+k1nZH8S6
pNljsDEepV88mURJ1R1DyGngc4SSIGK5SN8mHLedbdfdCpI6eQQvSGuJuCLBuo0g
Gv2+0z5QPhpDoEkdtNWLaqmBNKNBAzjlqx02xXun5Awq6iyio6b9QBzZ6XGekVMo
CMGMZXmDdyH5vmvBlgkOQ3dBY57jG1sgsmEeHKOQNLx6btwT/LNH/EcBrY8RXV+R
en24KGm23XBmXrIE1erZWWaKV89EDQLyhCkx32g8DyZ64lzRwc0hJHgbg5InmFPO
JZOYvAkVDUCULH60/+DggFCciwOs4wO54bf5N9+WqPOYuPC1JOKUkFAJ+NZHVYpk
KRxkMmMAIEy7528QpMJBwQjgrMKW3iJNCjlc1H+/SCWFL0nlaHhxKP/8jDVFDLEn
c+xbJTWRBZcmcjF0IYzm9UJT9B31YaoadLMOAJ4F3dbH+HGoPKZ0ipj9rS3vfpgQ
ifrTxZloWN/oL3V4B+VeS4vIusmaAFbb383k8PXXYXFpJYV0/ZE/3X2bzMN6WceK
Bs0UUsJMrICn1ymA33IBgkbRth2xdgt7XDvc4e0Rvqu9v7uv1BT/jcsdOW4Z3m3S
m144HHmUBB3WnyWuObvpd7aHgDjSiPx0hSgzb0LFUH7sJnrhkQgdgOiLnH9jGwDs
H4Moc6dYjlXdWx2bP7id1w2CS5ofB1fA/LfUwP8qylmWILBzL4WGCNt+Qq/4zwnJ
vUuIfhUSNOEjsL+blA85XZNnWJr9RCVKrEom9ZFfgbwUKZvTalthVRXZbDaXUo6c
+Sk8oxXW6BOv/bDWaG9ro8jQucSr+LayRojpJD8a0jZTnyHGUDsBkdM/tLsWx9Mi
jlEsDV5osFJluxJvd0PkNJqdOq/yA6P+mFgtjQYeaMRizHf9raQGxdSpWxw4oNUu
4LB9Xq7/Oj9xYmgktgAxZdb80gdXvnhmDcJEM17o3JO/r977D7AhnyIEVj576mST
/YCADMNuIouvbtOJNYeyw54+Ov5bTQVlwVFpL1OnOZzVOA2CUrGMVy1vWLVUlxpH
n1FYzw7aHE/Yqxmnwj115yrXmvT80cdFw8wgtjUpZqtgUSAhU2AFgfjCB+Gkr24c
R98IO+EHkwFrb0kNBB5/O1ALYIUyAhRAwV6DdwZrKVzJhHad4fG53xhk7u8EkO9a
tw053wfjJDIDWySkgA3d88qwjBKSmpS/jpEjdL9GbW6X03iL7JwYpLgPKDEHJvJA
o4oVEo/s0GzKk+k9ToKInhvaxJ4SyMEnPldbm2jt7n8+3AzipUqpC3yEeD1eLSa3
yZ88UUJT8P0dWP1rckRaKdo2CxqqjpDx2fYtY/aZfknUKbCw4lmJOedtVeJWSZFj
EN3nZ8tI5Qf0d1glsHQK5zmoxl+ReziwGf+d8GMzH7v5IUx+EHTKnXVY8SkxVumJ
IiOiepK+BzDpv1lQVE6Q89ueEY4/krBjOjeTRQ1cNErAg83yuj5JssJN29QZ4ANJ
znf36kNQiDPePBt9ourdqVRWLgueOxgOYPDL/N/2kLQxMUITWmRkexy09zyWi2Zq
p9xuk0cDJWgEcm9aD0P2cXT97D8bfPDXpklSkTOXJ6STJQTLD/t7Zk/G1SdNcNaH
t6T7SgOTqhEgw0DSERLAJjSHV1ro/54c75Tbr//T2gD1i949v1qcg3EvOPywVVx+
EqRyqGoy6gQ4w4KtW6aGmjIFlyTTNLle5zpugEC+M7GlarM1iqWDw46xw2qhLwJp
bqZt4hkej/+oce64liZAqVKi9utlbl0blFNaSlOwIg9IKAU+QsAV+nQP05Fz6R6o
1kOdhVKRrb7ujeR0Pv6Tj4281IlL9gPQnAglL5Cv91tU2rg/sHVA/iqFYAvFcOFX
RNhpvcWbGyuwmAYGM3axsIjKhpue2XWGdev1nfGFr56BXr6KU7Xy0llTGZkym53M
+p8vl8zeV0YjsaQXvdXZ5s4KC+fLBt9eJdh+e3lC8podCvz4t3YnivaqjQT9HZBR
6bHGGkIVzfvOcILuyDgqdMqU4rilGF2Uvekp1N7h+jHXQngoYK2rTYdiyv78kS+/
9Aa+6XdnCS90JAzV8ORbRrjErUm2Gw4GGE1ORlvpPDTwg7kjx/MZsI+9HdYFlm0y
cXaucFaIP6tePBVKK3atnUCqQkkXER1AqC8rY/k/KkyH+VmWNdfAfxSb4PuXwSnn
EWWBhiehPICN4bljP3u1IuMv8KaUAQ1PFWGiXXaGVgQ50u5bt3v0qxjmUNDQVcHJ
VS7P964wcYdcActSAnLq7oHRuu0dTlTwBiIO9zw1670Z0YwNdtCBRwA92y5CGm/z
WR7dNZDCNQCJ0UUPkmH+m+9g4WNuYo1quZBGW6M9DSZnFduD++IDdUsbkqg0ez26
2925aiaVUNorpvFZLa9ZRW7qTdjJ8wC2npjkGwFNvMyKjlP8PyF3XpA1FXJkV8Af
hXIGGrQauE6jHp9h0A1pQ0EzvKbOEw31b9jQG9S9dPcXZVu/Yc7x1Fh0G1/LxvD+
/O0hC8HtGOTeQohqIEfgmJ0lffTBEdR5eeLEeLfjEt1TUEKqxGzJzACfc5fPSP0e
ZakTlbBDodp+hZy8Gq5aO1oyV+bS4t7Wew3E6lZe+Vth7OrITVfYlynFrV/GiT6P
YA5MSh0a6klbGGzMIq0w23ZNQphfrPqU7RzH22Xd1ApHB8AH1ViTFBESR4d4VuYR
lUbDPOz/OQNoViukhLa/ryyS92KOdJXsmBgDmy4m9Z1aXwPz9Mc86S3rtvXSQazc
m3eZtmJHBdHbclLzSOomUDsjflmUnv6j3yZSDNKg+Sj25564X6GLqS4FuLr9KM81
dovzWMnnioVGI1L8spsG4oh9sMk428aFGe+F86qwQwRKlKn22T9js5o36tszo37n
JJeje8AowjySs8LNg2yV9oFZJC2EZyoZwOlCOai4YKZEqn2XsrENNefaKcyKAw2r
EbbteTRysg6YGulUMo8DzpcgZrFRUh4wXDyN8HqR06F89ckQToYUNMZWT6Ia9o08
qUM7mpdCgC/kd6sKuyBRQxaDT9yqQ2pWoVM3I3qGd+NSHvUcP2TvSoRJFrey17Sa
yQaex7iaxk1S+D9mlTKg2fPWJx073t8GEPzA2bCLSdq5FC6k2QNmoKCnv7QSz957
Je/kGZlmqEbTlmKTBHc1ARBjxvWHiJDXh3rNtA9lMCkc/DmDISCCTex7cRNVglbP
ItZSYMpYKacQBrXnuH4BtSvruxEx0qtfgh3gMdUZ8D3UYFuvxWX42ErtHbAP8vRJ
rKyoZp5jepRuGATJx47005cGHl/+0ojA1PrOiO9cMbmbN+Y8S3M46piDvKQUsjc2
fUGil7v6k232tNHgPoaF1mLU/HhfbkH0+3HvRvMzInsZCXKoFUSG85jV1aCGp8aT
dRBTCbVHZwgY9TA+lVPcwarGKd8UoXJhgnQ2i1wSO/c3hK2Fuu1RnvGbtsGwU3Os
HhQZPYNnq12GCTyJW8xd0pHWjSAxl6AfBKsJZ5HDuqmKzYWCsXTELLzBq6wflv4Q
tq7D5r6Ouz/Pd2soF6C+WRhebt+FMGfX/awItoInm42edhfrs2AcVwMjVu+VAsJW
XNpDvdxICroKeAOlKu1Z/hUrbnTSRUbMiHJ5vMZDdx2Md+PfiBByR6CaxqJspKMr
WaRrquIB0Le6o4G1XCoAI+D/A5kcqvKhyrBG8ERcxz22CBrLgSyk0JoX9Z+75Qe8
YURjn/IZjo1h4Wdk4BqdJ4ZO0uA5QBLxpdmBeURZcG5Mu9ukQNTEaAnI7uF6W2Zu
IzOmnXP7JXLeyUFj6WRE4HRav6UECLUcd6gkgpgDwOsvwqi8gh59iUa8WX5ovh8I
HvLrdCJJZVDah/1BwX+9nlo+8lN5fmUb4yA3+1iRatAr5GMAZBAskbEtr4Ydbu9q
5yNImOA+6kLa9KrYRYH+HI1MqkRSPtTLG4dstAvNqT4vtILDfpT7G0grQ8K/2zeA
WdkU6sj3Gvt4X9G41xCmToqoBNYmt3IUNz5Vam4doDbxN4xTGTFYjXoNDU7U72X/
cUJ9JNcL4LB7jMAMyhY79FHvvhn9/1EVVsixOguHjJX3fevBkR5ju0d632uKjw5A
/dNRaP6Et9/1MHPZOt3P3ozGrMgVCaoWnmo3vDmm82PbJGLAXcOTYIYK7wGeEjj0
wCWpqfdJPdRwFbH3R+rNGImfEn8lWCuRDablElGB/7DuCoPEe9l2rQGBQeVMSkH0
zvkvz35OR5p34lvaYuZ/OJk202HmBDROUjiXAbDDdorNe+x3a6yG6xsRmjVCuO/F
eGmlLyaxVR6eZrkeF1TXpi2yF9UfNeo2kJ1JkkMDRxFbskoL7+OD8csHSEQWWjAR
MwakuMes8E//VcputrIMbU9Xb2yXFPoCUZQZi4Wsqgyn07Gm4z9h3y/YPWcS3Sd7
7DSFMcvQcR+glfwQ8k4rrl4Z3s6Tlrwd76ZAW0rDzY8CHb4JIptLj62SqKtuf73P
Zr/X2cSBKlIk41TAwZSwsyTnZnB+rCgUSOlN0gQUKTrkbTxNpIbZRXC3DgcGrMiv
rlbt3kDI64mIUCNyINTGaS6oZlqd3Tk+TmjYJydA3Sdd0eg1ZCR4ZKpEr+GHGlTy
YORgz/wNDcYk9eXYVVo31InbkXqG7F6o25pl0oMFCsdoMb9rDZ3Tmjta2ujLA7CU
qpxzyRoHxwMxMJHvfxeHzdmPIA0F6tVIGQ8BekIr4d405aoz4NR3ZWl81EQXWhW/
H9ouvs3N7j6449hU/V+tBncUN7jNdXKoEnoelASEW263Ou7vBoMdq85mP7ea3sCm
zyV3aTs4/wZbiGIL3g0yjvmrRIg9jQJKL3Wf2ux/X9Eo7BHX5gO6pHbJHHL7IA78
P/ht1zqAoenUZEZ8VHfduJizscJNLSVjwvjmKGvYAsBkeOhWAPH5DvF14+cxFrsc
/XTW+KdWCmj4fHAVDod0GD018qW06lxmNFiynnMPoS4Aan3md5YC4e5H+YxBGGer
/yBo9G5hg9kYZKKsw1bDFIbg9fVhf5QvqsGdRhx8nQ/pkEOlGLIyRi4td4o9y7ZM
y2y7UcBtxGoAM4v6xsIVvdyvFrSNSe2QnfgqNqBCao6kqwlxqfshINACxwXbpOBZ
e1ctlCA8fSJdL/wOQHlGppTERZBaej4eqBWFSTWZXcMMxKZk4ysE+i/nLeG+JUBU
hPzNGrb6AW3/QNSWClsXJA+HVoZwR2kEmqVB05DPp6+nRKjLt+WsfTl+ee+QpRIx
AvO1k3IK+MhAtD+U7DHkNPk8EaYBEotqOF5wq8txsiXLSOEusdhs97PkgPBX9fIi
jTMzavZpQa2ZmMzL1fxjR5QKYmdcEU/rrTkoo+uj3iaU+X+Hb9AvrZQhRqM747/E
cmmAbOYdCV4NwGT5ll5rPO4f6Rxwxpb28fpytfRzWNtrir36k1Q/uRzuryicxNq3
AepKOI32VHqiQmJ4HVXRrP9cDVXt5Y5F4A0Q4j1z2dRdlfAYCmrdog1Xwa9i+cHi
aZHmLx7U7H5sPAhnjacGOWAiY2Zrw/ee/ABZdnQFvdyoyegcx2yj9Q2a6R//dxlN
9gRUk4SeAlYzwGLbqw/f37wmb3VGTxoYScI88DOoNh6FTxvoHlOg/rJDOufl4G/m
lmx/sFfU4xWJl/NcwjH9SWy0u3tNdPsqyD/BWRUknHFpaU0vRpaAjPusFpag4OQA
tnAcwOA9NRieergpvCABDlpv8GUga7ix4kbGysjyZpkot+HBVxZVN1Vfkk3P7k04
wrFRupnNrTAM8UXp7lkCGxyUVSwziBCKfiwFayh0LdkKxUWZh47zxyt3VQoLf2fN
nkPA3Ubaylm44NnldBARWZRIa0APIA3w1vH5kQXB7TZUAad1tMVDMz89Nr2Pck5I
24Txn2jf96RfcPfmIaozecA+CEeFmhzUyE6hOZSHk1UeHt+XZpT+LbyHWKm6YGml
/8ACSGZbImE1NQ6Aa01wjQwK2QbEbRnWBwJxVk/NTbgNuFej7IBpj7dR2sF2GRiL
mBIq3HUKboEM1/XXxOj2uLKfaCYqWWAVtbpdJvhcIcMuI+7LUT7q/IQVFdW1kdDE
w48LTe0Gzbdl3Na+AgbTn738r7TGv6DEBFApKUC1z13HHVxtywPhk+aHvJmBcdf8
0LZRwS5G4GMGM1akdCpVSgMISZFn30rFe3w0EjzyEFFOi8wN4mqjCaM+1WV5eK19
zCPAqdG0orSM2WvWffafJGqxsn+B3Q1czQV+y31IWiVyPeMenJf9vtZHtYW1fB1Y
Ip9n7b2HPWbmwkhwzsjcLovDSsG+kg41pUWXiO/pdH2L7fBg1zabGnezDAWEsCMS
IhAQQKq9Edx7SnCnMsFCt0BUFSZiuh4qQH0M1PZMo/I3HeWHxlIthTQlPPPXcDDa
e9iTPRTnPdpG1bG+MTEvh+tgTJ0KLCQK7KUXmGmJNq1qZxZeL7gKKlOzL9gaicGe
pUq39zDQNeJH9Yr83fD+qXm1kje4oPrOokblePV0CxJe15eEfjJGmLxQXhByc82f
+5wAXpIhVPR/J/b1m+PkUfVDgdrXI6Br23tsXIrFC4Wx7k+C8wyXMM/NQBOhhWnU
DVPd183pyVCxbDHtbCt4sl14BtR/ZhfBuu+g7fHwOxNcM2CD8NnuPGoKUvM7njmR
+ZlrjznyHyRFj36xepzmUI6A7cuUcb7UUdBLYKsZdZ/jfCg5KunaHESZn1okgOWm
99ZZjihtnUZeS74lwd67WjSP8WQys/AgUHiyi26fRHRigpFeR+9y60raFuytp/pH
CiP0WMF+AkXTgyz/YwWUG0f2hPx+niA+mgy41dKjT4j3fwxkEevytM91DyMjo9UQ
L2iQvYT/PkXIg0a0zV2FjxsiBZvhthmwt0lkEGHgIsg2EcDHJnHpYPLzHnPT42mx
Af1ykRcp4IA8JdTNOna0lOECOHfmy6DVLga1ukSeJU8o1PmGXJCVfnoD7LDTBQef
nQXKQEws6Vqw2CzWQLdhNqs0MFAiLE4H1FqCq3VvD4lZVputokdr7NehQonztpFz
3NEpX9nruW6AYkrs1hXLm8X6arVBc+hy3u28s24EvbOe0pemJ71WWkxXKJZI7mDC
Z//1eOCcP1SWH19C5c7QW+qXb2vJH+zF/5ZtR2Tvdcy14qestTdi1QLDBKt4+1GE
JLpd06+X8jkhF6NYHtwvynGA+DNy9Jm0uNU4DSlv1rpxMevCXhu0y9YQdBhz60n1
bz8+mwEukfFvHGolFV+B23B3+ZFdC0KNrl93naPzNJzMQt2v0TmlWlY3RFFjttFq
yYOaQWMrH79T4Lk1OVedHwnax85dENaNk0IvahUqrNhqC8Fh41EToQPs1AZVd/sw
eq4WjR0zzcyd+2QrVCf/Or1Ef0kh2KBnRMgmprfpxl6QbL/NYeO+pz3huANTQ9kU
i9a4nXQUQUH5fVIVUWdsKfzqKlkFREMmtgueQZuQkRMuw+E692q840mGTgu8ZmBR
9+4MpkpeUv3pOFBvgLz8ghm+YmPGmaaCID7SE2VJmCfJRHsI0noY0mC2KO0nimuC
qm//CPTM4ppAD+cv5fb1Zey+pDIsDUPKcEsapSqzkArOD+SmPcpCpQSTNrqDZlus
CzMusAFETd6vm50qidqpDLhlBdeteoauNRg8YTZqPB7nvQYjrWHkDsjhNT7he12R
t23yeOlnGeYwLgdVHQbgZ80Sb+uVzqgnuUEW+rZS0odCxMyJLZLdvmzbGCZJgjMc
hb+/9L/mwQxdbGrmRFHzLEnsiJ1FtFKoei+b+Ux2XELFXLRETuGoLFIUgRESfwEG
6Dm1RkxaYNCQoILlEFCKWazjFaCYf4/oyfvwiamXaTgxiBZrs/yPpUWjuUdf9RTD
wgWP68L3SUOdWdcWOluWiCvSUoE+FRXWBqSy7BXGxyUz0j9CY/u1yP3YYtj4iMnI
JqJa3qqCIFvaHp3bsWSP6Nn07BVFTy8YlPBhifSLMwYNVQF+xv/3KlPSHBhKl6Tg
IlC05hQplkLp3vcOxFebNTHfj9fDLXFf6EZPnwI3sRDuVlmp3IGpW4/J7ebHwBYI
GDHqW0VwSo8/et8/k5aehuZHtAp7mrkpNmDjf3nhNrSWCS0MBqFYLB2iGv+ZpXgT
sT/ZKo2a6NaLYc/k62V4yomQg+1pWWRU2Us43PITXrGioR9loWU/5vBGPQU2jdX8
x+MUqkLX8eqj/nYfd0VN+F54BnmcL/Y6gPV7CjqoxmlJvJaVd184ekJJrSmU7F+Y
81f5dX6Q6OuAtpF3kTGbk2t6ua1rrYfZlGUOhmZ02Vsz71qHrGlLKZ0zRJaDaOxz
dCvu7Ia45oKVLHrB3+0ExjMPwjSZQBZlYpH0iJ7n1AyHrtmWpASuRVsthKlku7eb
UrTcXpZI01mQ/RoGANthXUyFCIsJjZu2Vq5kLMDnQnKDQIZtd7acl9avtOR6s7G7
vVuawWQVArPm2uAoi9pOIyRpul6n/iYzn7SS8HT5IjKD1GnRIeWcS1HB1iAtnCMn
tgUZXosieQ8RlohPlpZh6MdIPR32lyDTAiwYcALkGNYbS5kEfcEU8u6kcvTVntze
c147GrVu0vnfalH+EHk1n95JvLPpEv34he3Dw+NjIB8+FEYiEGcKltuKauFS7K5t
+pOXarlH4SMZELQzbBMxqMgqDLn0kCbVs7CcPy4/SO6V77qLvOW1IN1xcF8WcdnW
MdHuE21HEk/aNmWsd01LPQQKJPUBYPw6dmggUvRAqTRph7eMC4Jao5T+G3qnRLjS
tOBORpkbCnbFGfvixvSr6g3ArunP2VFFd6cIaEY9GzMYmJ1YBeqgXQSRnr75wL3E
iGhL43hS4dVBt3YgMH0YJ9DWikiXCjhGN/DpwkGpHeeeENDQHrjsgv1zi3fr/2/B
kiX9DPJeiuWU3w88gx2tJgWr4BvIeMDw+enMtxh0T/6w/yHBmdFd0mu+8iJUIfYN
i388JjCNO8eGDXsaTBxIU2TmJ4iHIyVDWwANVmO7EJg3ksn67uC7+Pn8i/BaJ8J8
uC+WEQ3ltyF1RZsbTY5nIrCFgd2q2aeIG/2DVOq229bS1CzDlDTHQlhhryTScMVq
iJ0UjPjB3IIEdAIMVpiJ1k+D44Y15o4lQwItBlyguteFY8D+PGoZxhhrNcGAtDR6
RCYq8TTjtmEc66aojjucq/L6NJgTzmwbR71eHoqq9A6hme0PBgx6BDZCsQx5Y88B
qrmrPXsKllD9XMkscPIVoUu8sOcD7Indoal+6RzswK+xHqOXYQTzNO2aos/Urt9n
LcGAWb8fD3l8hmJBXkev00sZKiAryBJ6i/GTu6av/cWGsnHCBBspGBD0UVZbUc3L
2k942JS+rIs0KflBF8vfk7W/56nd59MA46/Tb8Gt+id2AV23EUYUsXBIK7Y/x/Ay
ZpdUP8fT9inpzkJwh9oexQFVVpRPcxErxDnhnaw3BxCHTvPNP6Pi+dW/vo3bIKtu
rB9gKGEBQVBzgsGMagyGqYAUyMR8zFcr2FiI3XCtETxTsIECHoeX9QTWZDu9uFAV
W1d8FV146GHORV9Tdn6nePxHYz34HHmKTtOFZEWWaydQ4qwRFF5byqExJGowXMmb
2u5X1jx8jtc4H6PLT5GvdGQblK/eEVmvOPLn1wjahbIA9xSsb6RXae0oWsUwNEXg
AA8VP5snRy5mRSc/DKt9gK36plfWbkiMo42W+6G97HCPtsrQ3J1X929KBG2xwkyL
Waogh5a3OhCNebuebifPic95lWVPoPggFHGFdgBv4nk4WnZ58KdA1leUk/IH/B8p
W1GiEF2qbQSCAPXkvrrmGREptsPCismA4cqUqpphqkn6yWbcDD3keFy0dhnYmkqd
19hKNpW6gqKRCzopzFq+FaN1iw+g1zMkSUE5Vp7i7gKB6G3a0gQohwlSN3u54VDt
ZrDmTafAZbiMjHsU0CDrHmVLkxWP4beywjb2wJxr/7TgA4detdo9g9RXg1OfUUlS
fIUJ3xJuOYHnmlhyPgdx2jNH4fBbHm2WK4aPfTwRdbchnjgF2+dq8Z9XBNlBatm5
043VPztEWsE3NBsNSP6tAllm8n/weYy8WkW+xCeVPJetXrry268UGYTgYYEZRWPv
JW6xnPQAo2q9PkirywZ1l4CIeO8OZNFPsM4dOZZQpLjLdz46lWfvuRYezZEtEMg/
IHfi+xLw8tZRmo8ZDNoqeD1E5LpygyKeObNGI7WP601T5xn16cpOO5mFhR2o39lS
FIWnivDG5bQmlDDo4NlBJvLKe452XlMujCcmeWhU36ITZwFwC2C7wnIb8X+KmQtY
Vgq1PMs3/h2DkgOzFftEy1O0bXDL7M+PLBYdvPl5FZubJAuoqG9WJu59bf+2ZpP3
juZSDu82u9fIVfMCu0ueKxXdSC3Fm8P50VJFqUMHFmktq8lSpnwxd6ft2s/VIz+9
Ow8sg0jtyWjct7UKL5PXP0H6ieHT90J3uv1F1d87y0kB+xjr/QPn3qDgwfwpajFA
7P75YXBBD6bUkU9DQ1kD4E/lovbR8Op5NWt81MDtliTOtHP+VKDyVjD73I8+1YWH
mNm2LSdbAsAIiPr13td9vcTRorpUOjdGqdZeBwy3KPgSkXIEdIpcvNuy5ZCjrBss
N1mGk/Ann0II8LtFRrNim4/hZBZcQaLrsJJMnf5RrGOFNVSLBMNl2hIeicFbR0G9
di4mr/OnYYDqG5M+Tu+RWyphM7QVHEroXyWrruhPbXAP4gAS9LgV2eoA+3ZLMiX+
AufhU4WnV6m5puw1Q4qZ+glgX7e4CarsIjbAutznO1jTbt9x0HO535HVFnUIqZOQ
oWwVH1zzJQEGUf8rACeQy+/9y537Z+l2X/ROdRuvhmY1/HGuIuZExcDTTM5TTVny
YM2vu5JouikmwfOqlXCrQknQaXbWWxAYlpKWmanY+iFZ0bRWpeKHTciiHZk6Ye9R
n02oYpqxynJqBEGG0aPOn+00UetWbtTmlNZwEijXaY5wJz4AFTIfX+NIvIxnVNKd
J0KH+HXps37EdWXNNyfCy2UBs8GejWMSRm+xzfiOyim6eGGaYN3M4ReiW4okrsr7
qJh0QEnDbl8s+3hEPbTc5hDD8sOHDCQKYOM5hFV1cyRtIdoHMGBkXN8yybJTDoUI
3QmG5ajy87rOpC/0Z0oj0svQGPKJ6jF3WnrUL2oy8JqJTyFqv7T5ZPkpwxmyNeSj
/KVSToJbZ1faO7Jxm/oDkgPLLuTWKEAkEXXLZaJZ9HrTGlDSZmC3+bjFmpEt2Su1
mXMUiYM8jMRigH8oqx5VeqZz7XdIeov9375+EeB4IJpdaAK8ZIP+CGDO6PnInwge
c3EbBkb6bv7r7e1u0K/JMCBv6S3WbDmEOytRIG+wMibBxPoDEVzZahhSX7sqC2x1
5LRe1jiodW11X2ru68R7fE5MjiHBSDAnjqgmj2ITb+N9Ufw2cisUSPnEPJyfFexl
Cm6Oq4ChpUrnCK3Eml/VC0Cnqnsh6F06siWXnZG1vbsfMmeq7PGGayNxduEdStvx
UBusXUDHsh9Sn9ekOMdYc/fcpDDjmPDRPhHuOOHra6ykP5QLyaQleQvtlyPA3re3
OASKEYSEa9lUZ1/9VkXnfEIxDqk1GBJVMrzUt52gYeuNhGneHaSkWQaEZWiQk1Rg
UnwxflkZY8b4ReXE3gK4If7Q95/4G4itfaygoCooDbAi3wSK8DiWox4B6afSnVLS
7DsUQ6H0mgEN0/F//m/Mbu6I8G3Teueb6IBRZ1EOP4wDbHtq80l3o8k7hCANEyLZ
2iYgvCMYPf+waI8ME/t7coeDWPt53ItIFTcK3Hg97v7oYVGUl90ruWW5agPTQA2k
9nxJ9mesD/lP4C6QJR2OingcmbpM50eJrm5JRBkOOMHi+nNqcdMdFjWyPAFZGhq9
d48E/DxzhdKxmpuXW7fK/Ci09VDFDWMIX6ukJ6Dxu1ksgEdurtRWAWmyicHmFBGg
1b8/whoULrE/28MY0fb6p5/ED1t5t4iojX5aCxS+dBzDwNLfn/zIH/9owTfqH5qG
plnUMQEhQWSbBXuWaFHFuv/g6EfIhdnwYQFiRktK60bVqdobV7pefooQNsfJxqoy
XOWWOnXxkbOfjjSODPKBrbf/hJ7RTtszILOP/J+5yk0sVTlDQwJQuX0zEJ1WKWu7
hlaACFZ40174qCXLtNQ9HDV4tehltJ3nnVk4vrayUdenoB2btRA+AlMAc8FpBfdh
mESbMXuxpM4ngm9CBs/17BZbWjgjsZZIu2esEtWYukHjv73GAh0IopAmgb45sXRB
Dob2g0PgH/eXE0rVvk9fLrB1wAkhT1t1TexpCEWsRNvMkGgTLyk9+r8i7M+r2APs
puPjr/FJGN6RcrFHAwF/C+csqLhWtYXJqQkoqS6pA1x6AweuMSuBUn9RwRyS0Uyt
yyYy+cHBrxwjRx3xE5B12egQT1GXnb8TGmCJecN5ClNCHkHp9EpvRKKZIIF/pEoS
tX8INzygIUVbGV1p7g4BnssqoEM6vXZyMRqrTwAbEExbiTmUSLmHayRRGWZj/KYV
L81DC8JkbJfv9o36c7VGVHlpizIVuNtNO9UeElpESaGm2dKh0eFjC/UyB9L17eMW
5OExtOWOEjrIVrkvKxrdgVSL4Z1/ISlZ6FQhpiXm7nNsn7LczIi34DcD0ulgSEyk
LFU4Ce5lSYvVB9Yx7Jshogtr1xD+oIJWaRcS7nRW+93lot8a+goNKxq5PRN+2Dcx
Du/QGliK3UNpyDSHhuF4EoQ3V+JVNfIVFHijPkXUcPVGPnX/ul5CvDpxXB90x3Kr
QphTxbfDGRiQZ/A0qBNICbEZV1NSSIRc7C2eVs+3YqBbkp/9qKl25uNjTpNXzbIg
9yc0wQ1Pk1WmPVISkvLRGu8a1GCAw1Wdp30VAwOTcV03N8DoiY8M8oRyYT5fSjt6
5MLpGmg+M1XqAQlo2JFuShuilIuHKRfipsHKMSsp4W6crXh+6kBo9ANQ8XQ9G05v
ZFqMgMvbBVwY68+Y52dqPM5uwH4DBhlCtlvTIjJlNHCVzQCFVKZb5f2ZFa88KSa0
bZjEhQL2NAyGipIwL5C2S2U3jdMEN9X8j+2VPpyvhuGnCYb3n4khcel1pbAlRPGp
xZSodYS7snzmF3DBs8TGVhygswhALbKwU6Tiwls54XgS4BJsMVq3Sbc3rrKNrttH
mMg2J6/xWztPuw3twpzWXAiCYE1IDYC2ZoKwRH3+oAh+wEcdSlX5NUyM0wK6H4Fa
hEvQUzQSgh7rDfqw5KfRCCiVymoF6eJSQNfL82QsJuZ9HhxKoo90AL3kdQ5u2Esw
YfdNmcp+HwCmHifnWPv6tyRwDudNiYG601EcT7r4M16hWIBsRa5YNZ+/klsCy5DB
9galEcgBhy48qkTFdMGajZruDzfEYs8RTkU5QCImQqVq3MTvkWAHrqZRHI5gtCNh
+yudb1zz9CfbdT7ohfjZZkAoJQQQXUwQsqWYaBDGRdHEbgVgpHoG3+g7BMeGLXJe
t3AMPpZ9am2W88VF0IYY3qze+wf496HMiudGyKYZrRSPaV7HcfqPVNpJ49XH2Nzd
52ciPtoJcbGy+WL3A0SztFlXxe6ggfiqrkybz+MfHv1qMMX5gY4ICaNA46OnUAjT
V5X6WULH6IoQMZQR6LkxR0rOng3pAVXMAHF1OTmzLzbCids9yv3bzfTbbwWs+i6S
5+3kyH/CvbX4KctAH1WhZrrpVidvxnrZDJ9KIT6GsI0xKgp4zEjgC+1qMll1UjZp
PSLg3ypg7Ic/f7I/g0Dm7VClTpS6AmabOF52YY0F6nSniorHjCWhlLFLRnSu13b6
dR5mcpogzxsDjckN19SUuRFvaIcdSCOE1KO8dyNFuwQ4C6FbDZ/TpyOSGOURuwzL
2EbZF0XzR0fYsUCNmk6fhdJeLzL/mVrj4qZe/u+ODS6NmNHgDP7Bc7MNqxUyWVAA
jXnN2CwvdkTNhhbbm40w6X19N+uKElwr2lF/7Q6bf4kKRF8Er1f0DpsSLPpgUp+G
Vm8NrS82BYg623ysSkNG+9ZTyLdAAjDK28B6f1MIN2pXNXfelEBaIAKupxsJ24wx
7X0Ov1Gyum2wVGLqvTH8rlHxx758/L0aNyQFhYv7DPRMrdmoG+lK7m3Slwn/vJOI
T8WZCyzBOVecLzgNkJmjEj6YoCRrxygCEvq6QVQu5y581YehOBIZnaj5uJjEbHYh
VmpRBInqjPftb+v2ZkO05OTsoloyUSiY/PBRoJOyIA/BHkmqQl6a8OIjPD4s6CFK
Bff+J8NYzqrWRq1ULqbOwz7+27oaCVi1hfSXIf32zHRTYHH0HFD+ElkFCd/QvOXM
Pq9sl5vN1JWtYQ5W2nZHjSNyeIpVQw729U05WdzUcx8KfwmbFcIAR8ri1s0p/ZMt
U/N5Pq4QPD7o5dbXMXgz7xXzw5vkZKfA2UXdWGXRSe4ebv2CTmyA5BQPdJMQCO3g
u9R+QWBw1NAu6AhJrC3ZjZOO/OFYzErraKVxHFdBzjwOfePFPjpRt0PZbmggmmgH
xbo7v9eMOId3rBx3d/xoREIK+14DZNsjFN7hfbV2Uq/UwPo8hSIUZkM/CJJUnpS3
fzjpB+fsI/339WB1NzPANacKH0LmSIGwqg6HeuEY57Ew6j8iJfaS5mLWbLA79qgC
lqMao49doXpkiodNRKUFGVPacLwl0x6AsoynTuEqQFpHYMQABxJHq09JKd/Wlm0h
x68vyxEsjCNZB+YMtVZ1PZItzSx3Jk1NAptfN3ZZlwq+93zibH3s6PrH75rzW+PZ
ddA73oIPtMlAogvoq9dTcvgcl1ArOdFLE1Fy4jPFdJlYl6Q7Uy8qIjlnLf+o1Qdg
/gWKnmFcJIbrnedilXzIK0P4Nn3yUpxlTEQQDfJJHukoQpjEB2AIyAX/uOODX5Fv
iSEIDn+pWVfIDqsWQzJ19OvKoZNC7TTxyraNa2OCjjeqvT4TfFNG/vYqd3WTo1Ag
FMBIRxJI4XG4Zo3Vk1ljjCh4fDAe/meZDfcgvU2O+a4d/9P5oPpE9jdIGLW1HCXs
fVYxwEE/p7rugmMfHv1So3F9YH73cFzPNC5sjvWij1HgMRevMB//uTjAxzmZfgGS
RKLvvHvdMNWl2W51D+x4S7Y1Rq/bX0S/M2wPyey0UqpjeVu6Gg5660/IW1QePgbc
H3GGeIQvLG0ZuNdyJtQmjWr/3QGCxv827Dt2zWLyOvIN0xcEhvdYL9UfCZfLpOvM
iBb5NBEUAYjVi3qtV5ubKxRyGoKpI69tqaqev6x7sH4YoZ/nZJo1sFLHBkce9i1g
gvMs8r/6cy/5a9iFQLal2ZIErJjfgAe1XmxXK7sCI9Dz5qQKpBmXEEI+oAKPCkd9
Il7iJycDzRIR3I3+/6SV2WW5NOoPTUd140KOJZcRpgF9Xq4tLC2wDZE6lHp8SvE9
jmIu5ss+VAXujNzG2qSmaLtWhSl23QUMYa2bEN6t6p9hUB4MIOMlKe6uZ5R7wBTb
uYDLw7s7MR62LAHi5jUfenOOr8Pwaq4yQcW+Wk/q6qIoUvomR20V9IgHjh6C8qO4
e6/1hRYelmXDhVBACxi3t7ooBl7yIJqEqs535f6UnSvRNcrg/96Qc//WzXx0jP4V
nUq5lw1qMlhE8DHk17FiEQ2p8KkrxJ8553ZkJb0treovVqc6lHKNqx6Av2N/mIis
iYeAcNa52Es6NbEcLfmAtEgAMxvtJ9eaJBqRlhLL5zWcZxL8Ko96agv0Qw540r9c
SVchKoRGAY7SsML5EYrWDOylU1o/IY+Mty/K5Jgh0V3HJR+GU3ftufi2k/1g/0Qp
/20KBNy+DlNsRu97jUysQWab3dj88MMs5t+GuzElU9lcwdqw2xNf/seBxCXHsavU
NMynEPkJ682vvEKejYGc7rRs3Fzcb4Gf0QN2lwQ/Y5gDlpwuIjb0jOfYwsgebFC0
v0cPGivxUwzervc6OL19WKkJZlvfBEg9Ape72EC07rvfWSogCWEM8BpbGwveUvdS
a3RLoGpfyAKx5qTi2j/OvF7HsZK1CgZOF5Ho7IYqhA2QKNHoQiO6fuYZrgfSt55a
7XI/XPYypNB07P55RghowwCu1WlweF8E5CYxN/5uGUlJgiOVBkfCxT9/Rzco0CQ6
Nj+t9+WNGPP4ttPQENwN/0GhZQj0/fTDenT6e8LaCzfDBi1gLh83yJO02ylrhpt/
fip4wbvfgJntEiqTSzgMaS9LPpxhf8iKbLmRDX7w9/5OhyYXEyXPOi+la098rUju
dxl28+MMweKN86yZy2dIqFjGZYcndHJ5d/fyu7zeCFbT/k+DtSSTd1iu9EhHBuuG
p9WcRT2CaG7UT+ke8ssRQxdksrswOrvCuV7TEvdB91mvsqQx9SVXKzuVFA3z2IV/
qyxGO5WVIw7E4FztYyukbrDRuYbRzvlimswE7VzoejZlMUWMHQ7T9aMRd9OuiGQL
/hYosMJEwt0Nf7mUNZ/hpq5HWCG0olvePpg7VMJO3VoLb84CUYgcvqg7AYwD0oo9
O7MCqikhQy/2ZYhshSKQwQhHR9pKS14G65u/n6KuUIDq/1574WP4//U2WFWaH6iE
aTGjc42hC9e3lAagzeTQ85UCEQbLh7LE5fBEF9tLJ/JwyPbOE0gqvqAQa2YZ1rAy
KaArtLGGuDmlyYRudWzzbB0Nc+QJrFqOMSUvWzHq8xxhnoNgrEXJHgJb3yNyPZiD
L7PbnwUVaC6M1Zp6K5dB1rIOlQfl5/5aX2Zv4S7qWqXy3j1io3LT73ORxYGytVOt
rT5u0XcNrMOXrkChzfnS2IAJ3+2ATxMQ6DbTqym5+HB55t2a/DfHN38LKr9eWog8
hfgRL26lEzuVnVdpqv4Cbvdl0U4j4GUEzaejNTPtOqhvqm5ZlVGcJb3LH3c0AFA6
neILnDgYBzqUXGsYtfQNX3HTkZO9rHlrFrZ7Ctwk008XSx2dBBy1v4ox2YbdOSl1
j5Z/i0B70u0jCcn7XOit2t9Uirjnu6QV8xCyzLfmCrHkbpLbm33dC0cZ9KktVoE+
YL+GCFjhRUghcJqX/r89lDantFgHIU1s/YmVkWvgFePDv3pBNhxSrPTYEwGxu2yY
t43WJ7Kc5FuEh91VQUg+fVc6+CaiRJ9RDf/Czb8N5Tc4deya44e+e8FaX/lnqulH
uUTePYWywi336t5Xv+0rjy+LvFsOjgEgNQ/ajfxqpWu2kywEdR+mzm0QWJKwYNv1
vG1ihidxsf3Bet3GRcy1yxGzTDs03dVncvMmjZDIh73ZNXAOk+5PcWFG26r4jm3y
dgjbP8jWhmgSFhFfJabRjhV1Jq4a9H+4lzKIE95aoszI+0RH4BO00MjF3oZf6Tqw
uB6UV8Pxz0/A2+TU7UskGG3PG+t8LCfg+1GSkamJg2kz5xQgvpPcyi6nx3IbFiW3
WMUO+KrGzdh8KpqDv/koEN3oztXT7T6IofArmvFkW/Y0hm3XUsqw9RZhqiBsUYuh
jI2bgT2nk7mVU3p4qBrFRiP/Gysp5qWMJQfsV/TEzedTa1OaGMH071ef3b0GRwJA
9v8bBt1pOYQ8ZTwhkhfDSi3E7bM2wdJKI0RvczsiqwlzXp+t1O/2NF19WerF1nUd
2BAu8evhO/6QvrVv2E+ZbUjL2LeKjbTxF5YMVnyq/m4g4QPM5LwFMkICzsdq96Zx
EXFUYoTh88/tJj01BAjqFGB/WYjmBQVTc/3/kATGIKspFLYPcKUsC1qMxeDzEsON
1sj/QsgZvqt30ZUYhvnpWsC74zxuhYpq5S+nwJGYThCY1UdKDQH6lDW0veB9wmsd
3BZT/2vBZS0aQv7qIjMbJCKJwUK4xPhSAc8sZQ2q9exxgz03zL0RjchMnvLVPqp2
qTydjYsZVIxtRyJdjnVQBbOvnO6eAREjX0os9pB3Prh8RVVp8CN4jprmfL5mxpj9
PTtBj3VUgUO7kN5zlKW7d1egOmJ4HbHGVDB/iGdN4qg1UyH5SrFq0QGFhK6TuK2+
o5PhiUZrsiBn0XjvWHE+jQPueQ89QzuSxydfOg6MxKjZjv5Sv5hqBC7OmIsRbGCr
KSn+9d7toAiAKMuTCLktLIiZZjhHeml/mhohKTHOWetBnoKIjfiwf6cAhXdnZ4c4
4/iq8tHiP5nzI9v0VbSivPKveS9v2GCTRw+xc1pzRej7g+MX+qj+C18tlRmcy1nD
0zQJQzkeqRpejH89XAMUSb5YpjLunhAPYOv1XupjeBXI2n4/hUqjU3+imjJpfWvd
9kay5PNRaHL2QnaiFKZovea1iXUH0Qjz8By2ZJbilUDp9EksgDEPUd1jjsIepSIn
PKtjtr+N1XmKxQP8OKqj2GOX6Z8eT0y/BsWuKJIeT/+v0bwtycZ8M7d4dyMswAC3
97GFYSmxu4cVOsfYCgdC4d7IMacRtaWNu5jRRUUdVkAgQi/3EaZeznXwRR9pxTD8
293ejFcvO7lpohopUlzKLM4P+c+vnz8Z77VD1T7P3D99mk4UkSdT32cJjETsyz7a
rhFPg4Vi4o7aGNDeHz1jBahkUhVTQZtuMaSer6viPoyFD2LYlyx58XailX6ubpYI
rIpCjv2OsR+W5pxhJBEg4qoE0dmYeXGpeEYkty1EkcIfwNGKgjO2KbzYctuW/Fxb
7NBVBqIUBU5KlzoTtzWBbwiGVgxt2V6Wu0XIH5ptEQrzN/8jhdWh+YHhkQ+DT5eA
AfUm/bTNYk7K5tTwHH7xcLx+VMHOEynwgEJYPi5znN898wi1DRkORAD2PHjlu+6I
yc41QZygY+ePlw7wzzHusJIaXJNh1o0JS8m2YFNmQdVHwBV4SnNlrDozw8qLBgFw
5p0cg2RfkeQ218J0eXGiwqoFSpS8ZoJ3FKhKRqVZymoT+D3fMAJwu+n8XbPv6lUP
vsweBANUkuYGUll/JRlTZfpru+1S6Fdu9HFV+m3XhAfgQlV2YXaBkd1J7ne5JvGN
9CBjslt0yTb12Iz6uTvNKHa0J6YMVvkHQaPbg3eS/wDcw5ew7SttKZRs9bYysYo/
oPZ71aPteM81LRW3iHzuQeZOY8CtEvLoGXEbxZ86qYmxTRezt6eHnQ3pXBDHdDZe
B+PQrL5mNsj+Yu/ryVBfJv8jSgT6ertw2jtHUB2M8K6frJ5HBaAL9uZN/+lqHqym
etz4nvE9ll+ZFl+em+K5KaWuBWwL2QsXP6VoUvwmUk8G7m1bx+sU1xZYVTt4TzC1
hCRZ3yyB/Z8xSBY8H1YNPROKeO8arVIp23ZN30ilQJCac/nG0Q8ODqocZCak+ck6
uVIxlCVhj9Sy57O/ub3qtrXZAAYmfa1ltl76dPPyZHLrxOh/8WMfNhfiFg5sLl4E
LIiLeCNb8erw82ySxA+784kPvCkU1IavWUbiD10zYRdw2W4clzTfryJi3+9pzQx2
PtoLsGn9qcENbRr7z6Oozdhui6cO/unvt4xpAWB5sQhW+BsM0wxBnN+SX2zjGrh/
LDsfIBdJwgNEO9mQSDindRjdTjYRAthOpKU6Q5SwXKd5wv9dH9xEdS008xSDf4WT
lM7kbfIz+JU7O+rdOcmxvPZeispcMwR1f7DjLpcUWgv6qcdMWN9Bxw3nhDzsj3MS
mmDOv6SIfATYyx5c28eCqWPyfLNBGBp2Wh8DlZmLjciqttR0MWRuwbL+PQLsbX72
6LeMoy1vqR/7kkU4MdO4dQRgB7HmEkRwCiOyJqiqT6kftTTiWDvDvz2MkZTxMEMe
a4X4KpCkIHTvpcqVGdqb9RRZkCZ4d757T3eXZQw+T7KLmKIVCcHPXyhZU+KFfzKh
Zbmcb6uarA6dZYJsdofwZSY5A5JaWGAUESFfYa+/CZHKtJmcBxh7SVJx1/oPZNKW
BZUQWbDGhFVJiojALzUKzlX4hYhce1GGYABmiR8GS3bLrtGaO1flyoNd4U2j1SAE
Io4nvlNNhS1V64lfqlD7lon6RV9hTGQACfJkN42Oi5YtpvQiO4LkzlcewsBHZetE
m1/tTLBCJ8m911k6UgVRZO0foVUVtYe1TF9cZpU7m9TyKfhQJWbH+q328AnnUNBS
bTRVFrhe+0I5fkUJdQk1K7zrHqfVnagerTiPWYclQ+xP0ihbTgsJ+llb0rUUpt51
hDNYy26aKiA/ZeRacmYdNZ1+Ra2Nbncf+KEzfkZtdUHziFIxEMTGI7p7d6lIjS2W
m7U9rCKEjkj036GNYmO9HPr66acy4mTCyskbaxFfPs6rSvY9Dhno8HqXNrpRxEUE
T5GCY9OImWnnCA++FrXWxnk/crS9Xv2CgDhdzVq+0xC1EeeCWqzrNp2olJzsVnAm
nWhkRUrwPpd9gQ4TTHYpGUklnYrnxIo0QPxLIw1cCZmkU8rB0/TnqIqp4iV29OL3
42/2OqjHDOIDSYNkGBiBAcuKDBe1GCzT6zbThnHzCI8cOSGwO3LcMxSwe7Oc9acT
5H5mEelL9je8X6+rJ5CwPA3aJT0bMtcY8zZSl545KT4YuBTXYrnnCIwM4iw7cXLI
HGYXjPLoLU66hL0bppUZoIdTdWfsUPd61Kaye4O29j7KIL5671d0YLVjxbmu4fHu
VFpnP+oJfJPLOJsvTyrBHHSl3BfTTE93BOEI0IlBMolpbfszf4OQx9FL17GWMqNY
FljmsYWWC16f2x8tYJmjginLM4u4lSX2/8XZSERgPkO53xKH5L5r2/VyaooCTm2F
Mv+aRfGPsMD3KdOJs4peC5jKMFZ5UfBgec+y2xEmCw/gH9mRZVsG2av2Xjs72AYX
F0GTVJ915x1QadGNvZsH1CfPpz6VWXlbrXyLFy+0q0EdH6nxzSKnWwWscKfhHmsB
xb6EyeTeqGKLKOwuLFMo+ecBWdVTIDUgx5+gTGvOKdbOLLmdGoGuNb9stcv7/Ok/
urfRbV1v6GrTD2OYZe4p1T9Uw6zZ+kWlMEIIlnym+j35LMsp63vGWyREQ2/dd+EK
nlQWfJHrTMedZnY2z1wUdvlci7oK5r9vPFEIv3jM9bJ/DRdp4FJ88pOQEWyYrgGx
Hh6qeuXorIgdyGr/LRTZXEVtQp7s6yDCenNVzOXMR4hNG300jniBVDD6OhCQJRAU
fwiFtKTu5PfzajCpL+OjkKdeDmqYWWXNb7VS7ffo6n0bu/I3ryBYr4MchPAq/l5N
pZYV1MxFvGHZrW+HVNEop7Gm21J/yaXp5PKTt/F98flKhjpnYTNnBSvtHW+Lb0v7
+1Y2BrSgv1DEl70D9c4iO7COGLHIjQZ36qc4zWJMJGEHJMjG45nsOPG9MS0XBv+f
eQBmoHq3YaHYe5e/Idi1xavUWuI+pBjOArVmLCGOjElIQvnQWyYAHaG2Lwle2Hzb
vt94V1rqM2hSzfR3/SDHEBMjlA/UdKZhxdINisuDmW6yQzjA7whnD4EjgG14X3dT
fJBv1a/B9Vc/uhnfHB5FWcAzSs5Ecvxjgpwrx46K5Q6hPdeeF9qKWzEcmek1Hpy4
iSeNGDJH/cw9tLjQ5sUGUS1szyuvvMxhTgGRplr3eW60Lq56Kp+434SjQMTVLlCL
2F29oC+aMpwA56p1vSL7iMCtpi/KOAusvTOAftRy8Rv9WASBDJASo2T17amPwa6G
6GrUHgFK9uepLIrihcd+sZci4HB8/YS8FjbWFc1PkQNmonkz22Zndd634LROU+Yd
CDg35GYf9/huxQNbU73UuYjn8uDAtNTcHc+LPRB/Zo6Wah+VZG4J0K0eK0U9gTeT
6i+Gpab1r3FB7rshPEtP1Kg9CvjnReMr/mY7oV7syL3BbMJ55XlZrijZlB2ONj9+
nlUwkE7iJKHrHndO+DdP2z8DluuaFOCKuUQQsfJJvtj0jRFvCGuuwVdj9SW7mfEF
zZ7esWvHQzA6Mt4sXDSqg+LJ5DlairA1lVgQnLA0hsnf/N3hqNH7CE4NzTTEYAul
pBKF8nn2cTj/KtS24Hrp2Ci79R2GNoNwwWyuopANqeVXlQPo8jczGvZKiq8h8oMo
C7m4Nc91YDeU4gz7J8trCkYVN/KidFlbcowZ6vPl/UwygOFwQtIPFn6pWsOddcb8
VdOfp+7C6jGodDfemZitM1XeZB701IqcNetuZ44kPH/p1zn/MK/lZsxq8qrEQk8J
jzQKpiK6aCwI4/td4Gay43GihJOoYfO5MRYJWqP4wo07pPmwJs0rbyktG/Mh0X+o
mR9Z7yRrQ8J1bxeGRa3mq+wJSbXtymLNDoBVyI/Nx6us+y1gdECGIqw4OkP4FZyc
l/Ls9sCtQZ6uXd1y9+WKSbRm6ujDm3Y4u+xBCIOIGDvgToseUYc8DwRuFaHUVpP/
jwOGWE98a5Zp0Xi2Ivl5EPUOEgzcySTYOGNFR/cmA6+bbFQLk07tOb+WQ57WfICG
v1d5ty5yldJNqLXTd8CgjRzMnPoO2w1MMhwmLr8CvaYDe2o0vJO1p5TQM8IUzPVb
yfyL95Jxl4sq9JhkjPCjoYTvfsZC/SVi4JJOBdntkVuOfsxy/iV0n0nsWiqusEI0
FlfWXJD/b0Y0TOIYsdTUiPVpdcDLOG7gwp/KTZpmlkbtLnx/SCN9RebKeYDi84YG
M0dw1C2a+oDygHWiKyVEyTy5gQGlk9fTDIyWGulylPHocMDU6/GhI9e+4SFm9IM/
cWdWO07KoMmIWHlV6NMvtUNWs2aYG3tVtkDNMS6Mk4gOQsV3Dxf7AdcqElAoVuj3
qLPp+u4k4AmZqwgHuDdG92miCehZGXTbVDr0wZjs7D3s5z3+KkdK4gtK+uhh2Suy
y6qZmVpSmUbGHjio+/ywNMP9taguVQdH50BZ5u5lyC2gNkZM9aqwmU4zEIRic08T
zfkdXscyI6HpUbwXdYPQTGQo5FgHYYziNgcxvSAusSsEGIOi0+mWlT583eAqaSBq
mswxd8gWCsjr9YJ6gElF/gS6Kc5W3SMY8OQO/bzGP7jKkRgAlI3RejnJlKSZgnL5
EVVqAZdZC43VVOROUAb3e4R7yh6I+NaUYawX8BcEWqdeQc+tA3Imu6WIKLbHMXVt
MhLs88GCmgB7zAk1b7wU3c/x8hS+FpNW0HsRHy7wYAIqvz99LcdU2D8x6JOWP+HH
xno8QEDAhiYnRpkJOBjEftiVCpJ/Oy/WnKWGP4iyZaexlCj4fA4RUTQpmf8JKCCC
dq8iz9ilq7qfctzCwcxyZ9dZA4wafv9dBec1K0aVfovoJbl814h8kIU0y4nJ2epi
qt3nveQP4AK+tLO/BZoyZ/Qjp/KChAu2kJydBxMhk7SrU8QgHu5M1VZD+tHCz+h1
gkvvaOBx2qjziWejxFovTxDBCca1Be9sVk0sYXN6I/yaJtcA3cZCZHH8t6pK5aRw
VNlCVyoCKbz9ei37R2Nj0N/CUQZEBcVgNWGEzbV8OJmpVgvSYSCL96pzXynvzfkV
1UWwXq7Ln2DTvRlPBDC5aOPkVotaWVvB4iEV4KyLFRlGaQVc679oAR64GZg/O5VK
+/tDypEiR2yC1IosIHmF3hkRubKNHOvgAi6uoyavtjbhgq8Gj+ZZ3CpZsWMN52NL
xvUubecpJyoOCDh7kkaGo9qqs8VVq08VN5vEQ0F8kxM9rVJ1p1IuWwSyl15nnaMj
V/RDxw5Ud/ppnzOq5i4pA1gktBwT++h0iL6KpRrrHAykJIWOApENLFTqCaMila1m
yHXExJHtZVUPyonDxRFDCc+UvAKjPV025Drb5lLOGzbb935mfEuXtM3A5WOFJDwk
hukWez8RPr7L6t65f/lMfIUpvqEKim15go1UpfzsPieE2KC2/jd/yy9bLiZz2FVi
/xbeCXB+ciySP5JgYSjs8y4LsYO6Fjsm0dFbsGKs8DTkq8myMsG45eQarBmVWDUB
QHSVVur4jInWEmyYlcRS8CYoJjrRPZefT1vyOiuvKC0h3t9SJm5AJZrmXDgGwuyQ
qQ91YwCY0dxOb3d6k+XEuimceF33SInP1i0xFAmyeyIbCeI76VqctYEQuI8dqEUD
Nl9lIfln0LnH7H5/C7b0Rq5mCwwRuXyQysG92W7SeQYOzFyfnNOWYgIcF3bYeEZf
8qcUU5PdWjLajNuzOcBfG5r8jod2xAt/Uzxt9qP/SGAFS294PVT0U8QkDZL1vP6R
h3w3pQbSZ7hRkVHkTidrps8eglUB7lcUru7fllCGIVGCYVQay1C1Rh6UMLCx9CKm
z/dZG85Oxbu18JWtkzsOmGmpEbpit0uLbppP2EoR9J9hcwvzJvtvv9bNDThd6GpS
y2j6AwwXV6/r1vtj71LRRXwS6Sm7TrTBVw8az3sVPPR9q0RMpj5iXVesh8u4hL4l
KSqrl7ap64M//l1OnWNQT1J6F70/t7yPbBu4DvJTUa7AETp9cgfOkFbTCUgsfrXE
wBMCCSpeCWqnw4q3ojGmtStxHdYDKU2wPYhwm8DA0dOCzY0LssZdj8m/f7qWXKKw
jD5oyrwyOzA4ScTOGnagLhpG5Hzi1LoXUerxlzLUCKQfSViQtRwUvfkyg8OVB8gD
vVE17mZ+TBc88vsxMyALBUWeVa8XWlbRn/E2bBH1pl8CkEWjZe2nZjz3+/vtR1Id
0DnrJ3fbq8YeDp0yhJzp2Xq3SLKbZqNhz+Mg/Xcd4a7t6wPitd5k58gdyLapTBDD
i10U5GwDxtimjaOtjVujHmFKN2uAT1lLkJyrm6Q2X+ZwogiGI9n7+z0EOl2S+FQ1
3CQGn3TrKouoGNoyNWZ2jwE477nVRqEdNOiG3nCyc46O6mNOurVrE1f/oWSg82I0
1uGyGD4ssIjQuYqWjXpOrIxNRuB/t6BtwDQB9URIUFWhDPTBax3Z9WcFEdlgb1jz
z4WGBAF06dgZn873d4NfjG08m3UaMP9fESQMRWanKcUUnGrxxrbz6ebEfKcanZS8
F3WQHfUXrc8e/qtrh3S9N8DGdi/RODLfvEUH4/KowPoGSuPA4PuOchorLpxBaTw7
jwAYt0tjqcYESh+d03/kf9P1Y1MCqNHHBC2N0zy6O07Q0CYrBAs/9N3yEnyU4bqx
tUcVghWWaw87IigeDwZ9T6t+f0mSw0ECM3mwS6yqdbtdsIC/CW3dxwZ8ZYK3Gfj3
fJcM12E90Qbsxk9pgHTof9OHikyNc09mB7BrcaWWGJ3GGiJC+EAw4RBoYPlxCQt5
/NTkdsefnVsEtG3c0+x2batFZHIl2mU9r7MqeOH8oJjOeRSAFJyMb6QXt/55sB+J
Nw9/00/UOk1Md/v64ioxx6zxSEI+m2wu708hJ5TJQw5C2IKd6TlWgIN+IXOULmbs
snYhWiCm2givdacM88XyO44PFHgHwq0fYoHsOMVWIwyscKKZp4fU3hg3mAVwlKi+
7JHLqwQ3vqz8605slP1H2OBPSb/2d2nJkUF2eJmJ7E9cxxIWO7CVtsa7lpTtLk7D
F7M+3KNQBr0iqllyMxJimvgK8bJqKEp+exVg2mItzxDivOL7cG8J5KwAOH+9/wpA
94PUCLg/lUu7MKLd/W4mET8Yb0PxkCPhHsC5jeLJh0U2gthD1zWYDHBb7NZ8Jlzq
LoKv86fo192lMDltWh3qNWKXgOCoLf9aVClwfL6EIqYHTUs3t2CL1IKqhyNfPwnr
pLFza4o/808tukEEagLl98H3dyb+2JsnDVB/OyHNQtr5mmy/6DZthQOWFNNMJZ5r
hCFmpTANDOZbkTW4I5f3FBxXdPGqth3WP6zIH4Jn1thwcuzRRZScBOfw/yk2sYBc
3sNgfVvn2KMacrvN+/HDgbi4Xcay1pTSuwxuhqAXpGqfEwsZh9QLf7uPzCqbAUcK
HClwbemy8QSTmhZijRorFBiMm/9DNtVlC+hNs/gSW/B+BYRSJwO4bfLRjlFaDrvr
nvxDq/2TnqHzMj3rGCpNjrh1/69DA/tbDHCTu8hlO2P65qwec5UeSDWaIIVa6DvP
zsH43C+b602jqd9dVK2t27LKZM3kw9oy8Ckm4dAkE4JfcEL+GY8dVlE+KNx9tEFI
pdGSFnfSz1vPgdytbdqnFAdFXLKYFYX6VIgnkEjE+ZpoX4z9FTwk23BdlAqw6buT
5TGVURfJkMJJPTkgMN22zAf7X5TJEfNWkYwGXfWwoCM7UBebYN1pNtlgCbbqJUQb
A7D5DGRjEemUSvBTm9b5MD/DU7E5fF/A1Lqs82PS9hgxuo2Mp0MoiFDW+4Ml1bkF
i/HTC1xOn91Vr4XXtbm4MQETuLSZNcO/a2S9pjW8wy143fFNw2UNLulX8lylVSve
mkNv2MmYqZ+u1T/zQEoj41iyu+MDP6KNClSaxS6Fynx5djpqSq8a9EgxgoEu49ra
EKZyH+DQQ58Gg1JrOMF8ga0lIzqW0A4x4bAVfwW8hYox1s4rcEyl7EIh4Y8cr+bu
bDc/wdcrWFhsJ9VVYZ/xjclFmvRQksEsej2AEssonTUGI1AWgR1Lum3JTUdovShX
Kh4+G4OLXYtHLaW0lMbgn7jRJhD7fTV+dv3Yxurz9PLjM1M7GoJOt8oQnNuFxUkk
GdrnK8pffl7FGsbHO5LKXV1dOTKSrd3kFIihks/OZ2zAuNaHd55mmAJapzkU+2+9
ZNBInmD66VRnREp+O6H/JSbykyUZ0k5WoOaFRpJx1Rmw0R+7TIPfuSpKIPLZi3c4
/eDo75HrIN4OQbJKs3lIRypIEBxfHAmnAikt7/jfz5ikFzaKm4iREvgEAYcI44Dj
ygJIVp1S2+Aq7dPcuwiaBt//nJm0V0qAR6SXcUVHiHV3/K0BuDxUfShyvU6tESsB
HTS7HExXspspeKDMRQTDTiONj84iTcwSYew5b5jn86NwRKH2OC0Ag+aZl4VnC8pn
FU2vNmXmMivX0EYXWvvBEc0p12nA9z5WUYVND9RdnoCOYACePadh95s176XVUpBX
5kD5RmK00CCr4s4uKKnm61VRMGGl/HRQkieicWi9Tr+XSzFUt26pzsbo1ye3cPuO
a2O0pDi3ntpc6pHCRx0VgHraTKoeM20I4EuSnwJFsCsBz54/LOV+p8xFM/4QKKQw
r7UZnAJ9DyvZoVgQgKlWHqT+6YEGajW7vZWNEN/LOVC4bURZByiDADp8qtmXAXt0
EBfYWIaLkmnW5uhe95bDieR17tWjz8fInIXhY/wKxTeQYfHlnmVXCl3Q6UZaDpup
NLF73srqv09R1c1iSaQJzHERs+uaKibSbkQ5+iKMy7OILaqHPYq7Wmw9WOYSH8Ft
hqOT9h2+qkx5ligbam6UbxOZGoLB3zOOz/kYntYsgaQBnUCNMqbBSCeOWKszm5xZ
IbENYs0K6YDf3ut+R+ppAqxawUytT4JIp3taoi8hz79Kwge+mUU+ynPANDO6J+nr
I8bT5FCNEChSR+xMWdnWm9opofLfTbGAFLFq1PhaMUxfl1RqmGZErxTAQ+MoFnIw
HdpnZJkT7e04iA1SUNIw0TnoLHDEfG68VUWMtzsPU0By16HBuwjlstu8GUOWLC9H
6EqaQRE/sAFOYH5rq7q5UuLaABkvqROtLncWoKH+nX+4ZxAw6Wgo5290IRkNiAx+
ntDC0AYHu+VzWM3aw5tDt1mjyjME4XHYtv7WSUiKUT7YkS6fODhQgr4gRY1eYRGn
gPSegl68Yc77oKFIT0xiQ7xTYvOQiCsdcwSgk9lxkkMDbHa+x67Hm6GoBOg0jpcP
CW0O2fdV/BglukvygydDeeXS4CtSM0he9YgNst5SOLD56UJIOP++8emADhDyK1Vm
HsLfS9wLc+13dUpZQgaEbXYV/84fUcITQFbdNhb5655Cljtoj+A3TrkqU9lLXRAH
tFy5D5RHKrOEg4tIoCHslXdR9GUtMmWXh8CjwydlAcEgBFdYp16x3aN8ZEvK0lYL
TOVLnUBsBJ6m/wYF7mFSz2bOaKO1r/pjdrcJ1k9fWRdwZNemhalTBmn+lr19/qxy
3IL39HiwcTUzSRfVYVKwTmseXKXlHWi3KvpcWDfLazG1VR5uv9FXkhpiIM8HCS3r
wXV85w+1VrxwP7b+cOApNgFs1P5kZBLTiDcSK9m98DDKkkaL8AOit/iMUqlWDOWv
QsoIVh9n8LcqqR+KcTqIeeYX0ndFqAOnxLXigQa6rNSX/Rb/eW5oZypNSru4U0I+
qCyJ9KDD6lQHtOM1u0sWknxlJVUDAX4rJ3PCqP5hVZ8SskUJWCa3+CU3VX/E82xE
LUC+KNee0r+gLkAek/9MB5Uzap5G0qMrqgceEO2UJSdyY5o6hhNoJdsavIOF5x12
//Z5uO0wko0OoAB1XhSikRuS/5564R1ioHLRsKfUr99vCxeCrAP9pm/RJhDCJfb4
xl/pG2Lm01TBji2y5WhBWBDqzD+9nbZKx6xGexxdsNcrIysrjxLXbq7xH5NTWlHP
DDmmIlTWmjkAamIG5/ZNG2QNYaDWwPlZ3OyQZ1o9ifmi6b4aHclUgJOE58pxRGtM
WOyRRRND9NBMoYpedM3jf5UAsrNfD7CQv4gtiW5SY6wgd2W7tGWhUAszd0I/ZKKd
c4YlpYodWE6Xd8ILnNwUQNDZpbjiqHmU6sCGibTAziq8N3CTMmsD5c3wswbu13wI
7t4cgFcoQGyXp/xeP3QQk34j8MUv0wunY09D6a5FzS9fi02cHCsguB/r/fGoHzux
HuG87xDcG6uQzl0rMNWRjnuY8lCobvB/kGLu8yd9FP8iiOjrxNA4SKH7JM47ZYwI
18ZUv7qdngft4GevAw7C3+F/NB7jFsY2Aqd9D+KVsmNYzoFty46DrHzzGNUxUarb
l7giAjvgBaYEO+kizQRLKHQN4aIiDwUIkeKGUnaJNqJHArgbWjsXKpWvEOliYmBS
ue9lNuJoQGaEZPy/pGctGymioTVXfpMsyOn+qeK66EJMtaTUhKJz/MJrvn90s59q
roYnWI72bt70gfjUYnrn3XBOJd2plaa5gBvz/ZTl+/dDziJcqCnJp155DyjeFP7T
/6dAxaBVWGNwJUrNxpwwjEhoayn1S66AFyggCPDtkx7PwURR/ym62tbj3+Z6Q+Q4
PFFhAvqFPKChBNUZ6SpqotK7MPeMKYROxw8XMIOBPWwifFi6i3s3RZ4taOrqiU6E
OqLuTlUEFfcN3xm6kDriCcHnpyO1VdKYuLL/53EZuklEn9qtZdsjR5cE7j4hnfYu
i5qYX3ccPb4GHkCCwFqfnQSJRYZg+zEoKPXuTiXiTx2p9nS6d73wTOn+9D9Q74K7
yv5P5QBaHThfPoiljlTpMVm/ETQOjxK6GWmyu/nlJXajinIFulCbfmPPyabHUFHo
dXhxdw6g3f7/UulV2qcGWlKnIvP1JlKUo047e3SycdS+YPzbuAgf0QRCGbWj2Mtn
uUGmbGxeZOry53RubGxA7+8X0Y4dQf70dooFqA3sZ+NaiClXBHN1pkZapcZkgSfM
mFgqomaqW2ZizAwoCrb6ZUNUPttNHVY9crfw1uliHyeGkXZUtzzwBCZrxnYHlZyY
pi4CBR1J+pXqLfq/GOjDPpjSYfK+RCm7VqRHirzSQnU2edMH10BUxVnU2t2hbjqN
GrDRJGY1BZOrdKddkUIG6xrSkdhaIYYl0RJUuMyJ/W74tKh+3rV3gZLu5lNXOpcf
G69ntwvjjgSO8OCDD1GPe0dhqXWQw8TEbzbJ738jSq1jZmTawgkJXoifj2u8M+dg
qWxCIefbcVaeeJQGb0L4iz4wyLzPwUU1njAJ0x/KjeDBYSDqj9Ka6VG6TXVOu1sd
hsncn9eEdEB/jK9brViufyjapeJIwvgbiZt7noOzxOM9JDeJed8lopm45k8jADhp
HTNnRRIHBKJILqyXG/M20xpE3sepZfZ/SoC5R56j0rvpqNRYWsxnydSQ8lUNm0vb
camixi0XtR5orA24il+29p0yrMp3mRz11+H0hyGOhUiKIXjCQDq+xs4IsZiDGODV
nHNlVkzBvU2E/iMXCFXj30ba/BlFPHMm3sUpeOWIMeKnngZ00H10su4Jg2SnGZ5I
7O0eiDk7EVY2lBBwFws/0Pc5I+mrGmiI0AeoVsdx3Bp2iEAzSxDTuWQvIg9Mqu31
YQCJ9/t7E61u03f0L7cvLNjZasYogfVmusiU23/cd5IIHhoLdBHqZkpSuN+YtEDM
McNgO7qlU3AszCanD4O+lccSrlMbZ+7jQxMQrGw8ToYryRrHKqoWUeQzmE07Esb0
Q7WGHCd93htCcBfZ/10GCm7c8f13sZzib2cZQkBmeW/8YbjvEXCurG8LF357qQJr
+e4J9EdHMpmJQjt5RNjuH4k8UmmKu+ym4YNeFUD74DI+WKu1vJaMD+rjgrVZH5Dr
At2k0ZOwPXWmtH3KRkooGuW10o95UjU5Ip1KpLtcGmRtlCrVBb2cOyoxRgmdUmVO
6IXWlJS6FZ/aBR+Ggu13P5Mb7gUvIyW3YOOmmVJ2SNbEdU5bYfwN21yAIAKIts2s
uj8WBpaFhHDqL3V3CiBUYQd225/y8FE58H26nmIJUjTbmlumz58jjQBTi3lB4DnE
17iUBgG0mYr9r2vPIGxmDy319UzzyB57gNrTXooKUNpWMROq8HD//JyMVMfAX6W8
5qMCFM95jGwNN/KFMOaiwz8rXAbITkJYb/LK0TFISwdLk5278dC/gAb241KRpEDY
Ymj3duHGBd6zqZaEBST+QcCqjJqH8oMPYdwSZD3JG9PFTvfUJXVYjXFhlpMywOHo
fpNtsfA2ccB3tF9mOXzDLOuE0k2PjYHrHgD0CpU+0WXlmsR1u0pGoOmwouIg3eXq
VAMuEaWYLNdzw8oKPxvYYqjt1UkajDdtJ7bEpwXRqQKL8fSpcBQpErrsWAd5AW8c
CLHNybqm92l2MB6wce62Z6BmVOHUcHrgqWwR+b+doVIK0xvkaeAcwWpsak6FijNw
wisbq7/xb3mgtNpz8AHOKpEoHLFRjHnatWZqIHACjCvMKuFtgeB+rjA0Q1LIsnKN
khvLespOJkmRxZPgmsgUViXMOtKbSXI1h+D5xmjZsklXgwZHQiF0qHt52K0paMPg
rdCswdvGqnEigzFpcffGAilLZepaJHoe3c83hZfFaRjwgI93olMcI3MivlBwx10C
khU7vJTQZbx39G6bTZlXd0POGjmrMaOZKpX01MapWaypgmukur5nWwIxQC6atVrq
/f88uPmFMEU95kVjK5IvinOuypbnLV39SosP+kuux/p4QUM9e4mcy0yWlpZwuosE
XeYGxwcGs0TAiH4WERLasf0ft78f9vkLaOm/Ab5YYzOq91lkLHWKNfWELJ47V7w4
9SJEYKvtU5lTfpVcNhbKA1rDQ+kBqVAbuft5mGal6Ca4OYs1asj+JA3nLbsNvCGK
z/CGl8pVDMpPOS5pwwRhWT6a8mVTTTjEj7E21qeJTHBEQ3CUCrvd0b4WALLvLnET
tOgaI9vooygHZfafm8Lvmh6ir6kCJu6U+7tP4kHeRv6nwEuz3nrWH2FuwcHVXsB6
sQURjNBkWq6/ORod6zYstjSKtA5xkTL0+UKEMAxsA9jDt6AYYGEwXoKUG05bz6Wk
JAS/dvG8mMcawNWILOVzlIZ7/3e8bhHkMOwv/IN10qlY3xDE+qqYFx6m07UmCkr7
lwIH1lwc0tVY6NkgMVqWm3Py0OtIk7EQ89GDzGNC2iEyg4VEYx5cM301DdpFfv3y
lrf0Y+C+dpMDaEcrdAAiy+kEdr0x/e3IZ6UVJvBPUGSekO89Q/ufq48+9Ds43Xj4
cwOEOb7iZo8n9/70y0ihMKrqo56xG36ZZ/0dhfrO7AzRQBjk7AG+kDN2HRf2BOgu
nMcsH15l884dTRQp8qzfwX5qIeJN5Ip2bBqRp8FghnmRt9WwIkpGIazdMfuaLCDb
4VwssVQp+3G7elYyiy8RQiejgiS6Ynu1LiuIxzuK4wvw0OMCZRRsu4qv20cFFht2
ihhpKfWKDlcOdkdGzn4/C4zHQmzVVfqEkePJDvDPdd6UMR+Q5ylRJa/XMbbMDUvD
2Zl780JsIvHtVc0ArMpFteLMXTYnbsrw/0xm4TD0eUKwWxT4kVvkugYTfJLmDeKL
WVXk4f9mHshYIabYOK42f2cAr3qVPwvBIezvlaRf9oSkT+sG9+GDqOkpodi/XPmq
2dkKBGUsYggjU4rPzIO6EJe4tBJSPgr4zPVbHrVKMFasxKNhwyjQsXgVVh6UMrSc
ceWNwgsOc5Q2oRcFrfmMAt8M/07AwTmRtK+v0d/+p0so3SRxL7y91lmgiFr6Ahpu
WQIiUmlW6q9eUgxzw91W3p2Dp4PByB92IisEZFHIXI+/k15Zomvt22dh32Hg5hty
W4UuT6fIe0H+J8oFLezEJDkTC+NypkR0wL01yL/Qw7ZNrI42ghn9Pc/AXKQ8JWXo
iqI7tsjkmXSD9lPMYnd0whZrjxfRglThdlQRuExo+aLReeuFPjzCK/ylL4T86Id1
iIB5ygcBA/z3CNYDSBXZ8oLR/SHF0IpnNm5JfeW9zAPMKZTk+v8lEKVJS/mOrW+a
pOOP5kBACHr87FwRJBctp8sYZCwLAsFagG8vVi0rgsSV0OnPebM4IgUiiN/bXsAM
umNdbyxlmRS6vModt5OjHDrfD8U0BdEsUol51ToJBJzQjYbGteszyR1umGYS2lD7
6J+JoxIeveTQEG1qB4D6GzH23OlfBX7baMRJxT/z7qCf942f7r3qRMzR7b/bk7c3
MeP8dPN4alC+FweIgP+bHDFLuinj/nFjcNh6XnaIpoB9OSEnMhetR3vAWx4Fn8vl
CuIs/5OxRI5CAisK434FzbQuvHlfRE9Uze0UzYb57XfAxjXRF42+cWAUpIMAlRwY
mSOZjkDrD23vJ+03wXLbRTKdTGBptqKfNu9cXdZPxWsuO88ryJRFFE26DXbW9yNM
vDbliCU6uixxwTCI1zHvSM2sUrvD5CYYf5UyKS3bDPsOl4uIZdQsPw2TgLXhw7HA
pFoGRmUt4AWFQV2O5mFDwvvwyuJBC4xkKfhwnvtnReyWSH4Xfx1O3eil7bzgmqyh
d8a0EkuHyv2kR5G5XcjxU/juyKHdIbeZrtCr/WsgsB9xoHQ3N5cy97SaBRRyPoqU
HsNyzJSmN/+B7Z3m0e0qFPeK/kI9C6z3byWPHBUoZehoSno8JeLCfVCY2NOM8MYl
4LZqDeoWSHT0OyOmx7Kww+rN9j9n2G9dWfCHT9dqWPDeeczVU+qFILr9D+3S2OYI
OMrTDnIzb4HWLcrqy20pDUmTnV+RDWNe6qe8S6JJiSdU5wJy8hJvg183uxnmZwn2
vtoIQu61DLfvgk1rwjjjHsXpqxN6yiSoXgf+iux+/kzb8lCWwd0teUxHEgGx97m8
QGUeQ8ytALKyVnOTsKzyh1peGjLqjlXV070RvZ3aT6SeGK6CqaWbDRtMvL9FSzKf
y7EnXsrb/mBX/SkbNxqYCMAW6GVG7o+FC9lb4FXXGBKBM0hPlTFuuHfTkZ4iyLCJ
GLBIwevlhGXoVV70SR1t7TzGV+HJ8X2WCxasGB1zPKi+9dZSINH2bFKd1tH5GWzw
1Ver0PsEOpF6FKeCD0XE3zpeCoQe7iCx0Rj8d236EyIphM6I0p+lTc7b60SiwwZ1
6oDLO712H5KbDHmCQgnOl7oIvoex8fp29ZLOf1KexlkNckGlBGFc3t8q+qRgMu5t
SKd7AxomXREDp8gArkvZpFgHvMoAhJcmohbWVzkoTDVB/Sy24NF4JkNN9nqowJY8
NyGTDOS4/sa1oKI09259UA77Snd88JsdnuukgySHMXKaBBpnQAxKmNjDzK23rFZ1
g3FBKLqGCkKfiQa4LcESmCoAKDvm3W7NrpkpHjdW8UKa3U6kBadN7ZJFjdBtxDXv
CPI6S8liQthe9MBK/TIcOVJyPMPxUM4p8roKoUYs/rhKqRA8MSllkcP1fynjwaQs
ppO4KOJvlTspSHV/M1LiYEVlemnLR+z22EktZQdC+GYxu9JL7a6StFJnwYd5m3+q
FUlK+dS6cDIROdPrc4eH2NybQmbxCdLJTtan99A4wudyCLgIDTC12uXQymAHa3CG
F2aGEKGy62/ze03QQSGhSgWPCq4T0o52BmPFQrWRd2DdBKqqgDX8O5ijiH87CJry
/+5Bdyg+RK3AMoai81l52CII3FzzN5DQ30uJ/0xmo9oDtAN4SOGpeyL6XdmBD4Sv
/90bzawn5lm3mRn0qeV8vBm8F/+orZD0f6O3Kq8rfFLkot9ZRoLST/SigIg3XwIL
RciceIGK9rPlEKOBLApKwwQ5OxEyiRwj6K+xh4gTPmbWeIv5pDYbXRI9jbfanIYZ
AtRyT6cuMHC5c2Bc5JfeMSgSitAS/mLjECeAbxL+RJgyl+Qq0QCe7n2EiCiWGAAx
BnH2/QhbItdS2fYxqXop7sRmHPtoJ54fwZHIRXVaHm9SWl2N2xTVM4f3umc3x4sg
5NL3t1qr//et7aZsi0nU2TQ7NqDrH1BttbB4TD1fO9vK9nZjEkdV7h0vqTOO/geN
aibWHy0wzFr7KHYZX32EPz7z3Ld4LR3zPJHjdveePGK/Cb4KFmRjloaRyBf5IAd7
nCPZAQHDjkvAaTk55USaeH2nKOmGQlABD0+usE+dhtF+1g+XFds7OiR1yzeJIm+H
jfepY+9i3YuVbLyR5FD8qCjVTKjS190VHYyc7eSdnFrGn8vxWWnTYewZDhIE1ep0
vicYhxWEbA+ZY9R9w/MdJFnOuqxGHtHU/ALhiMfrOtb/enJVxhyK5Ry7NCCycrKf
tF2LKPnaU5/3hAM0dwbRT6B7BOzAgv1BNkpxOdqQbKimFD6vrJfvYVRXCUhTZNjL
QVmooqQFLMqgy4l2slkm2w253TL959O3Brz53Vkj0zf/dxKWFr5roSe1c4M/pn3W
+fxTKMHhc7YZNIBcyMcO98R43ZgFHQN6JLeriP0sAnBn4B5mUlR7NxTEdg8zQWfT
TqWLxtx6gx6OxVAcASVOje3k5yLtyd8FY3xxgfu4VohhyB77r+KveM3ff6r/kwOl
LA2VgJSjdA2mmvbYD8oBfDpmLGN33+VyO2feuNTmSGmE7Jl4cuzByAwzgXfzHrEn
e9PAZlLKJU6R9OE8F9Mzrd1QQxhyU4w3iytYjZ6v/SesFpEYFPLaj2Y5VWaaE/0C
fREVku3CQJI+5sO1F/4Q7qm0yl9PRmwWkdcp4c6bcGIYev2IrGVlI1/xWh2x3Izw
NApBTkvOYHJKK2auqMlUoYtzLHNqK96n6MB/7kJXJDnp2p7AmokW6V7cGIJ5ZKPr
JVfz4EbDagZXsIkrKAGePycj3eCGqK1GkJeiH2vi4kQGTn5Qqx6mxF8i1IpHcs7s
4V0X3ufihnoD7zYiYYRWwDXSS55AZY6bdYvcmVk6Jc/SOtnWU+2F2lUTZOvyfpse
RgtpgaJgANTkyFvsV3lohJ5bdY6DbzmMyrNi2Baj4DDUefL63NkDiRkBps729s7Z
HQTzqnLzijfWimGM5oGUnjBvCQ1LNNZR233jP/tjKkNLgvDcmD9HSscKo3YGaf2W
r6j/7rCSguzM93u3Qb5h4ZkpKhYd5PFkcThijoIzSV3dbM+lnwOlZY36C1FfxXjf
DP25EAuX5ItaqnU+w3ZtnzgoQ6sTmPn5FbXAEA8AIzVlffp1KE/s6v+uFQEgMR6i
HjIO+DMToqg3sRFZthFik+wIL7wg1dasb6Ipa4b/EVMsU/Tz9nGwJehNd48Lh6St
jk4olPIljEYrs8AdZadN/hZIskKnBtJmfGGhezDOmGCJ2Hyaa6jy/Tn+zN4lP+NU
A0k1+R3rnPWQZrshF+u5Y8pkZaRu9BLoMxbG/6hUC0UhuK4B3qs4wcLkl2j96OSw
OhTMnrjCFwUjD6jqyhiuPJ5xuE3xW7TFrRkDpSSiOSmfyUHOeSWULEjnK4dik2Cj
fcJ7PrHimYrml/NojD3WDcBp65Oy9Y7k8sOCZwZmB6jmnU/VHD2seAIr/7umha1C
kGQ5cNogTFck1NQwS5/i9/iXZapc6KIj3mdoRBWPa7UVJOpDePTqoBhDEh6kT6Oz
hJgC2i3f31xogFsiZpQClfB2xfBwYQvvySCbbczDvHN1fzc5Sj74QmHYJA1haviT
p1EPhJUh3/I/OguIsPrQkDVLQPJ3PHK6SFzFsE8hk0OJ+Av4GSzbqxjsFGfEpjYV
dbC+lIjBljfMClIjhcnCzoCVrKBCZgI0jy9JCOkH3u7UWeRNrTd/V0PvBNMlo+ga
EhH9uD4QugLdZI9JnXzu8xqwwQfMhPgxcN6BfGmzjW+C2Pcf4DaT8/uSIZOarm7x
f4WHKd2pngNwYp4kd3jJKblI3C/bmxsIMoBDmNUD3pMVoyncNbSvgOG6Yc4Wrefv
wo6f3xVdVIkwx2bOH5/dtQFcH4F4nOB+OmAFecjAtDUPUS3/jdPZkLemeJjMGnW4
E0HHPsoQ1WCX/zE80A+CBqdD08g2R424/bgGzEl4WqyKJnNbIJndQ4okZ6+ESfxg
G/V0P60YJFNbLv7boNE5akz+BQybd3EVC89vZVzdZ+y+2qZA29AZ9d7I8aQ3G7Gp
617pRmUZmHO31Yn40Ew6O8HGkX4aU4imYWpNXU3w2Ej3C7/POL4KMWY58/CCwozr
7usI/WSh+8heEg8djOpns9HvxYyLxX+u2WtUhj9OM/s833nRP9UIDhQwS6oo8rn9
Ok0xWFCBDof1gi2xpUpuOwoJHiWua0wf2Rk0RevL8EJRaWWUhWK56gMdcejxG1hp
N9L5x2qClWVZlxc7+1bLLKkk/R5P+A/SvA17GcZUuu8eXKdScgpsetiWqjzcrGMZ
mWGgoJu9UDxyhWPlxOsWZ/yXyQEtucqI9l5neiGgAxymjidSLfe6UPaKWAwtfdr/
pWRkQgq3aqyoVG9NvP03/WYgxGIC6Rp6Drf2qYJqhY1OjDmuvXRUiN7oD9Mtfi8Y
ygJyAFnX2uHkn142l2k/t8q2Yh1bXRLYooWb7hlq/09hKEjvbNdOVCVEjR2UEsDE
GMROcowiSLHCTA7KO0FAUFwct9CEwlP1ku3zk/YZO6ho967oVcdOTwMpQ20vZMZT
dLaYQ9NJ3DN5X7lNNgI538Mbqk2qdEsiohPpjdv0V/+B0LTkYxJCqQCt9VcToOzz
o3oOjG6UcIBBf7lKY0D1ucOWM49G7asdnm2n9c6aZfzz1Enz1HoCBpgW2FRepnSW
L72Jd8qGCmc/B/koEvx503IhNn5lhXL/aZUhqGfHTe9heiTwi4oagi6AwmXWb4pv
CRb7Tgyhf2K9fOTDdFzvWAcne5H8Q58TT0t+BNygmqxcrbqFcwRB+D9+CkHfxq9P
u5RdrBQSsJdyB63UDbjnfZm7/Th9sV54phESF60qvt1FcgWYk/xN5/rIR0wSDb58
44YgESjpmowNvuAJQU6t3S2SHvNdOPOWLBhiB+1paHgsLaEm4DjBRpKfUCO/mEZN
+Kzqmv0xd91fIWzpVYC7WbL2WmX0x2Fmr9RumdjM/PYIGzo38DiyuJiTERq2yriB
bOBfMcO/qLPALk1j5RDQ1ECtyK2ttuTSvUfCXVQrnDhF0n83O+4mgWOba9JxI1n8
QN+ef53maBOqEHYVF8LLEVuc9uQBieimK7Lme0F1fqZfl2Q4Gz47iWpNudRS3yeW
vQvUf8SLtSHE7pzp1n45SmG2B9pJ3T3AzMeJAPb1KHGqEgrC3S2+zzhLwa5wXGPq
LQiX4JbhJUQgWAlyuisS2MCu3XULOJjMDIJuRzGQMzfSV5ZbP7FRvD7IXwedmf9S
vZY8FiX39pl+Etb0w0kKCPqQjGeCvKSdPJCnA6Vv4eldWRavBCVZ7l9adLQa9pRD
SscO6cGc8mD/dkjMOuHFcd8u5XR/bc7wmbDBdDrqbrF4nqxWgeAzl0UsjQEWa5na
mHoORbzcp1huWMkKYG/yTYzq8armmNwi6BhHk1VxU4ble1DuxigvGFPVPFKfez43
BCxPAuz/u1DZTZjpYY/BlhwbVkqUsmgJ4rv+s0+mfNAtmenS1VjYVcX5/S6Kysk/
VdKEDQVo3VA00C2LQ7EfY/RdXcQiePmilGM3q9zD9Qjq2c+EJavvL8Ry4rK5PetM
RPX/83LXSWiPaNvcQMy0zNKx0ke2/OamVYroYraL1qLdEN9fh8txdgyxgkKgqEuv
Mj0367k7NcEOBbwkloG2rpwM9lTuikbA5KAywYN0OIAVcV9AAphwzMMjPXozgLjE
vQxa97QgQHFwAFNIcIY/j64epShl8skh72974Y0H0GyIlCWpBycqOvCsAkRGlASB
SQt5cI8zqnlQoYXlCuQdr8gRiUyzCoEr8ESBc7ZiQNpu+dnlEbZcfL2QEGSCZFlJ
YNwlMiqVj+GBiNl+aBj7Ea2mHBo6yQv8SoCPE0c5wDRK1YIXBUtE6Nr6NU7Nh/GZ
TrRLefNZ+70Pfe1rLK6d6CrFzj088AEY9B9EMs3RfSOdRUezz0GIW9bYjIszAPwR
kkRLTk++Nf7fQD2BiQcnucJqNrvjgDpTXX4NgQKfSR8VwE1UI1zWyaqXtITXcAT5
kgkdPXwCKZxZ8+oq0qmwQM2RfPl/NIzPPm7ahG7p8NSYGLUCqf75rnTQ1YXXuHyC
ZjMZ0Jc/nTwhM0uorxUIDi2ZwKHYxuWNw3iP87LaCP6zfnSGg+PNjFpGHF+T1oow
jO1xUdw8l613Myt8ssN2o2d/DeLtEXkaOV9lQChN3nWWLDtE+AkerQCWf+5/Ex7k
mwRrSrM0lsOnwFvVvlyNQYfesM1DqCMRO5lY61qCd1CpM59Kq0vymU/+o4X8jhaP
gsKZR8dSxWCGW48t11EBM+Vmadg4cTcmrhrA1oqbEgny4Xagbl5MI8KX/xXDguIo
DHug0TPc64PEWwkO6xA/oIZMjC3FcmpriP8NPzbFNl+UIJZsdw6yu5dKIz8OGl8t
SSWeUlpB1K8YPbW6XUoQBQPgQTma2LgTZH/PsKS7P9b/XhJzQrQ0Kvwkt1mtlQle
Pnyfv4KkA/dvGEOBxYdRxSnNpKS3Fwf1csoVvjM2KeRKOWPbMva7MzcovEscNJi9
HqPzENNf0Tew15aAz75Tzwz01098fXv/O4pG0EPEyoYUcMJdsnGnWsZzICRbq/Ns
jhAusYPurrvAAqFQbf6cqpJdYdGODVaSxWRH2vbJcDc2Gb2sB1F6Qrbl7hWTYnyH
40gdf9rhUFHixQClFOXCK59jpSx3Z0QcnGnOlMrZbKDJKfL4WEXOf7Z8eMZK9SUd
XyrGQayl4XylnmU6zmKtxNT/HzN9y3xFee9ZXhhfhgYFfeLLG7cPEoKOBqmTra1A
0hgs1tw8/4peR+8/CIOcnSsmhqE8pBPyXs207GXg28X0ilfeJb2K6SGwOOwIRBt4
8UtHPxNW/btC/2lVcnPhQuXPGMpifYFwrhyp5j0mwBPMGjhkoJQTYCEJ4NhxsEBq
QxG++0fi8QWHZrlhn3iQyhrPtjZVuyKbGqaSuNx+bTYs1AM0YqcsqEiAnfNTBhFu
teISSsVugtvPBdA/riywAuCznY6vhqg59uVGJMEzAcBnbLOvfWqjSeL1IkTt/hqB
XX67zmAByJjigCwelbLfk3cqxSe53nKHGwwMy7FFKGRQIS3xu7tJuHRVs3haaLQC
Jf100fsoTzC/frMaDgtZdKoggR6Ap3dZOPMbxVpR8XHjj5aHUnAlirYopGiSh5Vt
SGCoEVfK0B3GwnFr6iWHfSWhkDmXn9/iw/OyYGF5x0yH/Oe6fx0+KAjnKCndch85
852+S59tYmriGfKBQYg0E2+cG8AKSL6cvS9A7aIiK4HYiD4HwRMS9M2h0wo4U5Dv
mIpMaMvTGXeCyKKJxhEyLSF7IgtoFXZ2odpMpxQnI3vGRyQa/zcuEAAOIsm1TAuH
FbCu3l/8/ffZF/efowJhN6W741JWTeEbVHZ4DTw0rzRZXyU/oCZoGLGjiVQKBNh/
J9Y6eASfm8MQAI6dNyyZhbmmq0SnHEr57kfMuaUFkX6r5mRuTxb/fGdW6Q9xPCuL
4+851G+QFlYWyyg8z/Up+oFIkzwTsp91IZuEDtC0QTuBMDR+5no1bpxUG8joZP24
qVQ19V98FnnkKBEvhBvJ7klrHUBOXVOVZxkIIH1vWIJTAXYyKbBz68t0en27Ahmb
JfCmTolCsMqRjfMUN+efRY1TD1bZUj0ZFHbiUkxaGoBDwGqd+XlWGaTgVypishIx
lrCevCHK3DkHr3XHmMwRA/X4Yh0uXg1hb6t2g9zOYZYM19kVgK2C4Y5E7HshNR56
lWcJXCnOz82D1VtjlkNSWPRKJhZwrEswg9zHgNE3ORJgpYOHg5sGfEF/wH5Fz+L2
8i9hTTWJCg/Zde+bUE7bPh+0cxseVnbTRK5B9zpnhtKp2hSrwyVlj0ZM4doe61a0
MQ4JQvkKD1TQ7LcIEDXyo5K+g+Xom9EzBSrDMv+HjL1JWAHFaPTPjgpzuskHy1rK
OW+VnYR2WoO/4oQqBN4KOqnmgbw6F2uFlHSG737Tyr4KjcKRzWiIdsdR5plOiZCs
y8C0HktSjZ7DUvhxlPIKh8jgHTtjiXJF8iNs530LDjWXAaVtf4IgatVEhXnNqOoq
pCAp5JjjUuyROlDfsi+ySlleYoBKYO/3ytItgYlnSG2+s+GC2MUg/jw4i6LHQACV
G15W0nRzDUvwa8hBjWiYViSvfIDJ/dTFr/8RIgcD+vpnfOo6NjMIkDkfERJm7oXo
JzLlHS6nNvhKdHn+41elM7uYOR5LZgOqqgqgLwqIoeTS8z8bVh+dpBGhrFm7gmiY
NpwzgCgl2IpbtjrkKatFg4R5Wrhl3kV5ee40Z+7PRfsse7RKzXBeNkkcO4CZbHXr
+7yFke2b3Z6DvisU1nLsaWnLS/FDu4VulIQYLZv/Mvkya6hX+5Q1GRKpjEdXpylx
BsCpzwkXAyl3OmOj+XpCALBec5Qf94JJPQ3rvahVVzlUWBmFDCPWx2jQ6tnr+wTY
I3/DEK2+mwJ6UA65A2MbmdddxylUGIOPk/YlM9Ucxd12DozSRcfzUShBOKaxK0dH
GPRPJPExH7qgU2BvXBgbUHuGgq1UyA+nwxJtPn4shrgf1lOSeoq6F5JryRj6LAdu
IXjsTiTK3V4cEPdWcpL3QKXbaRA2sx8cP8WzT4MSLvTyil3Jz/FijoB/AevCqJXN
UHiZVCDVWxi3zck45TIk27HG4qd2YvjwDxnyaJfQ+gDp6X65TDB0LJfrUAOd8lwT
JUyjAoJ0/K0kG9GeL4HoFP5tKZrhK8RLUGhvl02DO9kNwBaSio4ijKcxnFnQuUR2
sViL8OYRdC0Q/XkCRZpdJOkEl0PjZbSt87xjQdXda4Y6/BwKOV0kDn0rJ9BeAE6S
9qFXW4mnU+vu1NgBh0wovU3aTS9OxOEcAShOLrPleDQrqqNzbQlLx2ZF+5QkXD/t
BngRD/Fd7avYPLSP36knJ4KX8wK8sPVHhk+SBUrfLwUP9nWoxafJFQPuDmZ4F0p1
aCx6lPhNjOi2kDnAgfAbCPi0slFf16M0QOsGbLsHIBksikWfIPZ4nxmhtkLLIf6C
0amt3fg0IBOFi6c0xiPz5Z6HHh8IFIdr810MQWRat/EqMsysLZPHxR+E+JS3U63p
y1GBXZSWECtyUuoD5JQvRmXQZNP/qkHvK+MNmA04BLt+oSntHhBYJG/FAkCp6JBO
+JJy3aP0yMAMGu8rYwFLOwdCd4URD89evHXIKiiwQm3CkfTQ2okImxhojF4YR0hN
Z9xuVX32YO9dOTxRDwR/4ycg/j8II9j8V4rTbUICTs1wZRn5Gml5yST/BPBa5EpK
rs3LP0XZmgpympuo7pz4k0IuMxnXC5G7+v84tmo+fVHaKkOSwVM+Njw7AgNau5hk
eoMsZuQ2VhmGj3F9JULSLse1/Mp1xYBg74WWscfl8+ziflCfhHDFpkGoOdaJOz3N
kccp9c2urSQnxUdhPFDi5yOzSBvO0al5oxLxYKJzogrD/N48Y8P3BijYTlGPPro3
FVSienT0y0It252S7Or8rv5s+4MgZFX2FstYp31Nzn4Il1m7ZZat8G3IonmrbDvd
HmldLgyJn6hi45D1fiTaXZt0UGKQ2GQr+J0a5LO82yIi/xYPxdGSwcsfeTji2yYU
voT4Wr2NIOH2ffoy+TToblTSFra7/ontaJ4IQnayW+j7PGt5fOJB4Rt60z2EC2s4
0U7LQQFSgsg243iOJSFjqhsInSLW91WeGJSEfXcUin46tE7P7hxWr7JQYx5ood05
dk3x8tQg1wxC2y6gCz6mPouxnzHzgXwEhEmNCCX2z31vtTALPGmI7HT9UT3I4DVe
MzoW5SGo8xc1zFey1/L7pyISgGA6erckg/if3Oj2epDw/wRqojmkHNRVZijKj2hQ
WW5s6gLU50E4L2LM3aSo1kq0td+MnMGxdGd0eHRMz6inFU78eB0R9oxVVCanWSkO
Q7mOIdIkh3CTagkB8GsZZV2nBHOcDVqpL5Kv59WVtjDx7QIIxFlyFslbumbsiYiu
JSNZ8racFf3T6c2XmTkzo2yXByBaY+UsitIcv+t+NEHdAT71+OccRPHbymPVnxKG
IuyDKS3zvQXLQwnw93mSRqaSFDJmljP92EJb3rqDktkXOcQmJ52aH1+u+iwoDnoU
H6K2rXBy9Q0zgCrWlcATQ+QyQd8DTrWVN1LRotRtSlu7MqhqCbL1Kd8gKzJJ0TOs
GFTTppPyApXyCyoeXGB/amkKgk4UPpmrBvuvh8JI4+VGrt8RQkL4Lh01k1XLQF8J
NZUSChDehsUvOy+t3jwEKC28wyYj1pVniqx10CWGwz8GDr9EM1rsLbOPAzHbfbck
NBvGjmqWBjKkKWCGWy1AXVk73DNLnKP9keK1f0MkwSh9NVVHUKIVMvbTT/Rq5KPn
CMR+Z3/RigAkp8IXac74EkJYisEeP14+MuNaucgrbsRw1SVWB7xKCOCCcyGx6LV8
+VgMcHKFCNzoIVU8FXOfjIgRuNxBzR9Umuth1gX0JYaVDIl76mq1JmfdqHVgjfX5
ycpcCidloZTxe3aYDZEGYDKzLauqhRXYNuZCphByIjV0989AMMqx3EHZ0cLt58K+
1ehGOwx67TsNvTqxbXas3/Kbr1iT3gHBLhI2zbkWVHQ=
`protect END_PROTECTED
