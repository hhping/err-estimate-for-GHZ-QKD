`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+pKnlvb4ls6AMvfwrXPaN2UdsVWqg8JXwDLtTM62H2LcQ6H2qcD7xfNuHaM/2t+s
jX6IZT8N/Dp6OvTelBvOvWCdM2gXMmxfkCbHDgmW5RH6F0PYfsm28ZFTRRhvz3oM
qakLzRbirpSkIGw+VR6KFaOkY0NrJ+yF1uNtvscpM5STW29EGS4jDhgn4353BmbV
/CZA5B6mk8+kx05K6NXxn2ZsExX4U0uzvRL88Z4svH3FQ7dHpY8okdF+wPUx+a2h
q7k6uCVhcRnBgzlB9l1CJtSzyKh35qSadhdFipKzSN+IYR7yRDd2sPrD9HVVSWNx
Lt2ALHLEqwc84dTCWSM3WzT+ddChZ4DpI6AokXNBaP8WQAxBw+R5KG3Zkfyxv77T
3x5RvpwqTsG1rhQw6fLyzCgtDFAgvR0u7nCjK4B1A/XNQ7XkMdfVivee3q6KjgGE
UlJMBpIvOlZ2qto3yHixjp+BrMhLFVj6WevyODIASFyoIfNEJLxirRoYtJjyrcWx
mRm0MUmxa7CUhB729pSVr5EiSi7xsS7uxC4WNJMpqDZQtGVapIP4eJJr6fhSYI69
`protect END_PROTECTED
