`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
os3qtZBbnL1JrqVQIaUv2Kwd/p2Zm6gvpbvvgoWW70nIvcALPfQc1xiNLiKgIkum
UFcQuD48jCCVdBdA7e3WpgFXeORKtnEVICPBrLBEO0mjpedN4TD5gld0qVBRY7Ru
/jfGu82XcksE1MjEGfXUT7NatUYKMFFUUvJOoxWVMgZvY0Q5YXvvye8xLwKJM2yq
ZyKEvINvwagIDqARAYyOjdbxplNhLtizL/lY2xp9df6UCud5isob8UBouLE293Xg
x1WFqNDXuHKwoQxuhJ+nu6Axh7KpzPFP8nTayXPmxU5tsAyJTfdzXVDyy/y3ygAO
Sl2VBXc+y6InchqadniPgb4f1/MQYIpskGFFXgBxZsNQD92o0KZzzFog3C7/luLE
wUcEtDdaPRd0+PMeoX19U5Js+U1t0rh0/pbJC5XqQ/22aw19b+SVUBVLEV5cvo/C
+oUbs6ZvE3jNf1jqR7ERNSdKTe2GViCITweDW+Lf78VwA6AsO1i4T1ZceRm1pjY8
0eTtS+wzFujXGFE2J+ZxgZ2bf23d4FRLq0BENuBDIPdSbLHocLRDnDJjjTteMPd9
Tl89SfNVhunw1K9hQzAAIvrtqcKZKIkfLypzfwbutcAOauPySFahrR8BTKAULnQh
AZ1NoV9cp4trfdhhKLxNyg==
`protect END_PROTECTED
