`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P+0uwy/pZTGkswlUpQ36men8fVGyR91WKfKP7xvGdDj6xuxX7/A1/LL4/b9rYtwu
YMP9YHEddSC7YuDT/N8bnoLe1qd+WTxr1WkQMV9IypxYsg8ds8cYSP+9Ulys6gCJ
CaoSYVdNDGtxACLcHFJ8POHF9wjaCP80CjPU/DV+gJlrzy3oUJ+nPoKIZhzIzpKw
OtfP1+IIm9p3gn6MYlaETSzhcGXLcn4JwySb1OkBngg1psTns+GYlQfeBnjsUAm4
p+B4G2dulK4IpOZAgasNstGN2LGjdFjhtQOMQywLwz4SeJPfDUIJev8pVxuXRZ2k
EO3ZHYUWHy2y0SqEf4PeCc9GWv+EaLOPbIUJ2psOE6J1i8wFabOa0NdSVDifvnDt
0xYpXDv8GA2h2SQ9tanaQcY26Bdx9RRj7Oo1ac4OvOGSLqMsO7Qv7eaJdkeokdpJ
3uLU9ELxpfmdBf6/T3nGPUvMrzNsrBtyN3v/DpwQ+cqhGawntrgyw9hSFCrUQgUl
OyfxjkfvXVwzP8i5PPjwBr8q3iv/w2fa6m5zeD1fp7CeJZMQR4kYcDVeOGJXLng0
z2c+W96T8I4nDlCeCWr2sETy+aoUe8V+Alp/VEF4z+IKnzPzjab1kiThfHaDbGR7
q3Vi5KLh0D5MvkvUSmnZJL/537zk1rNKKznLng2c8z/Q/30pD8l8T+bnYISrSb3a
J/7PzGOve5K0v7bJdU8R1TsgQ3/yFgFP3QE1rVMG6xGAsoGotR26ERIjNO3B6048
pgxXq16p5E2uaCNbh3I890s5dOr8MVZPG1zRx9ztfot3AJzLf1se0efGRMAYKeQF
cnsv2rlXoeYRZo9EujibqHxilX9CXw2lXPAvDseelRSJArnIw4hIbb6xGr5yle+4
Wme3NhlmPPUyDprgdMQd+VlDPyBXbgF+4ICRdiwGO0sXGy3LAifZpZFxdeOptHHO
bml0ptBUOWFnNOYuPLuCv5IpKMlCvUWxukZfbQQTXOevIR40eR06LezPEZP+ia3P
k4mutbNn+1Z5qPvUDk8f7tBG+Pw8tSZ7CEbQ0fbGLXY=
`protect END_PROTECTED
