`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RNLSCYURcF1SDvhXAiHYsroGKuBup59SX5uKA43AqlzF1iC8UXKUo3ETwjEx4Vue
aMvOODjGfEYHq2eQt/BT0jgfrmgFAdcO4BZrpx06EiW4Ny9+AXl7zkreOt1jbeoO
q5XsbNYE3QjP5AxOf0N2tQ3Ryj7pgd+BJv7CAgk2GQwVDZ0a0RR7sV0n/byUqQmR
Nt4c3i20zfvaPLQc9Q13aBKnkw3OH2AsjQpSPoJ6JPrf4BjgVzVjRuJXzaWHA+bR
oMQvqqX2lGTCTZLyLw9A3ci4BGvgBSebxGZ54PwxrSIxUoRLkCLIkh2VWsTANHv+
3fDsA+xpI+CPCye4kWfzkLqRXcj3MYWaF+tMU37jnAtAMMx6GqGqBA91jeVvA4Dn
z1MuBxXlq/LRc7HZ5CGRs+5wpAYwTmVuCKu4LHP0u4g9DvLul+/JruEaMP4h8xMp
RmVILBjZs0wfW+OR2YJVn2bM5V/+q56ePT+w5N3nkiO7cwy0+PuQZ9ehmah9ZmDZ
FuvVo4mbZcEBhlS0RS8M24tmCXspBQJ61Ifr2jZYed2kgq2P5aU4Amf/HSOTgqVO
rjeL5B4Yk0TIY7AXxrxxtGMqkgfPzyLCXAW7mCiClBbwHgNGg9z7pQKAE+b2exoR
B1Xgsdn3rElfeU9CpTqfRDxgOOVnkH8FQychdy0hQG0sJd7sm5wKft4dsyAs3Z/+
t9hpf7/TXgyuXCVVVG/gZI1Sqwou7Dri/SunbuBLCiewhi7co1EBfRvM0n3slf3D
/tREyqk9J3mJqeRmTvYpXzCowOuz/n+4HT2vs+r7VleQrG9pI5u7UG6XgxeTgymg
i/+hHw37ZALCcNjOD52JPA3Oew5kaj8LVtXGPxpG+Pw7U5xOR+By+7rsc1fPUkUy
t3vH09BEtR85eKoEFEJH4uqEiX5gNNZLV+hMg6LwgqCK/V5Zjh+FCnwJY4Ss9lC+
VPg7js4zF09q1DBm1dMfH4ie8FlvT+CuXFlrQkQ2W3Rc8MNbyBpUCI/uV3h8FhE4
Etz1v/ANtNwdUTk3hjFihoPQnpD85NH7iBbJ9IY6KdFGkrzrLeO9eQ47GBT+6yPk
pz+dprXhQHem37R33yAbpo1AkVz8+Rwy1tEIDVZq+9IW8KVCtGkoQCjM0p3nyZ/n
atJ+38soUzz9UnZIDWcIipVkI0ONV5079TYF81eXrCeilPf4em2A5nhM8mxAtWEh
UbP+MHdxed2uXI+oWYaFoCr42UO5CIxckGNxOjSwDBf+TPFqsSBM4WsIMybg2vd2
PsEKh358Onag7KgMLlD+oyjnACT4URugRi1aNR6hlXenC3+bHiwLRrg66deLOicT
zkmEgl6uofwAj+qn0zDZgGs0dAOICO6fLGyRfw6yEFWrhsGQ+UQuMzi9HbkooaXY
P/vutTGeSdzX5MIkNo/14qYB+0IbR2EJ0O9i7aK6NTQmMRBpiLRg+QQ8QgT+iqjT
jKX35eZYofBmojhuyzJiFJnZcujx2U5KljN+cW0b4w9hedQCY9nVs8vhLK0rZ3eV
V5DSRaIaaF++CAaCm77jWqiSKWXoYfnBMGkH960ZZb/BxHSgDkff2gY23uz2QKAz
OMbYO5dxJPFpsJuK89Ld8O5/9D/1HjnKl389kEqK4+XbRsDfvFunyIUcZaFFr1ud
p4rtdpPwkihWUv3fgDCQc4EaAQWXSHrN5EklmMo30YBOx2gr7OUjzuHl8vniUdcI
n1/PGbqpYo7otX0LadvxVIu45NxBiQcHfC39RENU3E9IE/3jiCecx0arIiaKhTHb
1mSgNLnlNaQ9KYXiMaLRtO8fN66egxuCgSoXxL8Fj4VdvOUidvRAZQmMhMREbyND
kaiypfzqtPTrlbZmVkVnjcoJ/oQcnGd8mCM15yWh4Lboi4u2hKaDpS6Z8cwFPQ7j
1ZW6H69S50IRCZu5ee1DUk6exA3LQd6uuA/O+AxcEXNuLjWO7/xzWMx5Sx0/aWAR
Lsj6kMvqzjyTRMtbiekwRU2DF6vIHqVs7MvescBASw4f+guRfvjKUOZUtsQdNpHI
8PIgUy5hY4X8CFFMb41K49kFLt4GStNkMKZJO1+q3r9qkIDVxo1aLB8vxpwxRgKD
7aEkZjQC07Ke8Rl44SucgqJNBNc188jNTm/ecXtAOfSDJAzJUCNiFnjCqdCu3Pa9
zGvASVmXPTJwtIWnuwKYJ0qMRDDcPlNA2IgWF0iwJUJQcQeCdD71c/rYx7vCoaik
jxVE1nPxEToTZFgCvYIiSq8alyh/1AIE7TEJDUb7on/l3YIwa8p0FrRTpYchjFkb
/6j+NrcsrnQA6DJqAPFAnqE8RNaHexJPnbSODBH0I5ML6hDEN/5Jt3SQvpfhTJar
W5lW7YsZ+lIwDXUE54xga0x+UUTSJ7Qo1nMH9Hvj5xtcEAElBvru8dj1d1/88ci1
tjegH09W2offtd3NsZszSDXdx7aFM/f+hf4IGZC3I3dFyuVyWErx6etJVLSSj9qD
zYcGzTZooLh5tw0MTMjH/gJuSzQe86wIGTlED5mrzD/jB1Cbz4mJhDEL4jL2Di4R
y3cdiiFR+9avAG6GSeQHGq5+V5o9RH6+/wCMApK6ngforQSTq3U7uUTl2mqDZ8vi
`protect END_PROTECTED
