`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fwG38UXyNR67Smh5qgV7zGNIG7sBJbJfa1e94oyHL5b1fKejy37l5Gtj5uat1NcA
rPvyB/uIWt01DmvoAUawkqghmPyfpjuSnorSHOcp4H/ChCFiIDu+gHIpRrfhYrG2
TnTuq8pP+JJyFGxF5ZmvyAmC3WuIB8sZvrAAiJi0ST9Fd7Ry2s0a8YS/Psq0H4CS
VdSShP7aaimLTECTHWkjcS8OtrAw7SN006DzLg4pNY0iLn63/nPTNUfc6Meqe7oy
RDOrlwUar+Gcd8h0/GacPr3FxWuvCXNsNJ8pBJ0OmgSQAKGZvpGLZLm56Q7q5vFy
mIaDNNJcukYgnHD2wU1Fb17Eq5u+pyDZJkbRLO2qvI22+BGkWRldHNFQtXU4eul1
aRmcNoeu+eqUKCIav7uqewTmFivNlO8ONn/kC0NJWXSlAsSq+q9jy/n4+BKx/0Zd
qgwAW1qoohCWd5IGk8GyD+y1NP2hBKYhuMkpxfujyyc7qcZhMyazaa2Jc7e+rDii
/35RNV8IRV+4HeZ38h66LvzJg/We7B8nArjT0VVclFr+cKgKMWp7hYTJb9f8dcJM
YH8k7SACyglsvXgXyj8NTYD33qffzlp5HLvnuUr2GpzE18FkIZ/gu5r0WT59WRk/
CrM74MvqY36yFNH4OsToi1RkZ71LxX1ekkOUkRcZculj0K1g1QgmTyCTCJ32wd/F
yUBEzwy1WRm1PQ7z9OjertkOutW/rKOPUBaDyk1B+G1lFSJIf7rLsPISg3wORovg
6dVM71xcqohOVWSDMDeb2g==
`protect END_PROTECTED
