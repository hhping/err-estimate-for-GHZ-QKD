`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p99b0mtlnDM49TwOmImRcX8MX8z9bHqlUh9P7Peh4bp8lGxZpoxOkemoGWlfVB+z
J9ozc5Af/NmfRXDoNiaP8yeJZpNHScPNnGu70ovMir3jiWGYr++PxClTK458+Uy0
QVr2JRPyuasIq7KRUa+ZJ9ceNNp3343u1lCsJxSVN3BGdApwPpOnUnQcDApojkoi
yQTDIGmRdAHZbIMRT9vDq+yLnX0B37e1Qsc70VerQFXP5foDUTH9qKOgNvc2cEeW
3q7e4omonO4Hp7zMdGHIT1nOyNLnAfjQUSC7E6x9JF1HwF5d/Fd0qtz/eH2cvRNn
`protect END_PROTECTED
