`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6J+H719N2eRlYnfCJL2E2Fkq8CCyk5/xkf1jHI2nqeyAvvIYc2RvhUauwMZEh6ty
940rNF0SJYZil2Lrh/nf9u5URAUsWVFAVN8JLmGMFKRoyI7a+an8QvdKprCr2sPr
JRxz/0PXhJw45P88NcJzPH8Bas/ISoMB7vU6IDOj3nl5Ku95vtpD0HSzK8oiWW/C
XtaC97cBItOHl5tpPH8iuUap4ABYQtWReVAOoIJ/3okWBuQ7La29FUCWs9bApGKO
RNzY95sa4XBAMVCzgZMnvBzmRnL3V71tOjzgelBi2LmB3BdZ1XW7C/nWZm10/PE1
wZiGpPgMU7+nyY5XVh/9deyWm6jmSsMJTglWJL1CWCZkri3bqDgEKWlXgjTBSNik
kTHnlbimRSmjlKxOWD9ykm+Y76lsfdwyMlzodqpJ/FfEiiruWu/vlkNWSvE23vfG
lSFglSwp/WE0yfGkMD3yOF3l8fgXaN50Jtnx8RFV0O5PrAa6GpHqnRwsJdoabDxE
MT+77Rswsi1C3WHL3oTJpjCIZK6dZ7WlDFYUWot7b8ehtaFm7ramfl0yFZkUQTCs
TbDt6tWkKxswCX5ZQ/ypFk10yd7PzjdmIXCxre/dJknnIrS3voswJZ/cLBAfpmh8
Pjdfld0AvLHP4L2cQuMeXPXvW2g4+0b6IzgV4I/EtK0AxIVDPrj2bUqjFhJSZZIJ
daiG4kCIBlyQ5l6QWAEtZuEhCGNoyVwndXVUD0tdRTXqnWTH7ilTQ0TQUE8nUEH0
0WJCHLd6gopEsOOay+zG2zeJWbFI8USYDfBWSaYPG6DCWuhw1zhpPr+09Bu6Peva
xxfZJ2hofxqoI8bJOM5ZopHUTD1wm7Fl9+3k86HqP+5V/aMDpzhqLv6xEI9Rh6s1
E/bt+7v1kscSsiZCrO4vAfUWb9WHbEW90YaIohlavlrNXIe6PBSKegmOAdSbOv56
zHNNFzWzafK3bc4dzkPlAAbtZm9I8QRbWLxknL9qtQtPYF6LNMwYA7Iz5pnrnROk
g0J0pHKvQA0XFIg3zRxPE/Zv0uoQbLJmmXAjB87/ECFaERxvt1OPn4D1AVy8/oam
uJwVfmO3zJ0nafQpILVN2QD49LFe6V9C6GjTfuyHDxUfvsaekNTkwzo4Fmr0vxLI
r0CXRh/aeDRd0lmgJ686qMXttAsyyPj9El95pCn0myPzMd5ZKrmNa2IxzQ/FOyzz
aEcASRgWToKpqWzbFEI2qyhtAvjfOtfqyoPVGPKrPgRhzxTKpFjzM3rROQVRUSwQ
cjESo7BALeuAln77HOSKo5db5Hp9tK0POtofv5Q9QToy6nKBWP+exin2c0maJCsm
/amQweAwN7DBja14EhF7zDsb45tfzKBg2ni6taQumHI=
`protect END_PROTECTED
