`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kCDE2pcrijCiHAQbfmQunPoNAHsuW+lbNNxZ5ozDOw4OqRIqa4sco/FK8xpnrud+
aX5WO4TGkh0O3cZudkQ5C+sV+YED+XxUeks+r33dJFQtJgnrLSG6QdaAt575v1w8
GuekilSJ4JrAPuF2oioRxHRUqhwgjKjbLglIoSRyAO6BzF9Ft3hrSUU7+jrlY4ud
sO18Z3IOgc2oViubc+uGr9JJpR0JaZ4HL6hrQ20Sj7fjOzGFUmQ4bY/zVQ+MWoXK
KKhi45DWWfVg7s0UrHwtxo50r9AT9Ut2spBHXfDMXlOK1tfdckSGxl8HHkoW4+9R
iz/IjwpTjmaQnNNT77lCX8Bjt8FJdW8+DP3i8dNYD77F9cHp+XlDO7oBLkLFTioE
bMMQofJfXoy/sDYzd/04gKxHJpjM3NYwxeQYJl9T6cIvxKV02jeYmu6+KXDTBruK
KE8bk5TAhJQJhgVpiU930tpeINkX031nXj00qEF0lBj3rI6LGD+XMu1K/OBy4iBc
QWD1abU0GWHWpPJLYD2Ki3YfkZwhRA3JbogZYVR3XUI/r3qFmCNgiFfdFbqTMFsn
gHY2OIs3YtswN+cDRbWWm7qV/oqXhBFZDI+GtfIPNBol1tk6Hq5ashHA4bPRavPh
cLfZBwHxLkkED7AucOnXSfX+LGRMzCkZZKf0vbarjKFx+SDpiDWPsThxUahOLnsg
Vgv2PFNUIRMzT01AeZomUXd8G2Zdzt7qjrArU3LQor8Tph+LgVUcWzKv+nogEanD
hYSlCFDamz+AydD7ii734ESUt5CF13/dV4b6mYY9R40VGP6m19bpPXvqbdUz1ybT
T+2872QBDS5IsEHfSLEZmLq59JgcUzspjNraHTIKAGWdz4MooIZMsct0UAmSndpY
`protect END_PROTECTED
