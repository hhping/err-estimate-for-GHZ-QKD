`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ufm6rgPCd4EoI4ns7XdTnG2477j9ktPOfQKn0az+4hHeGoW050XTwLpulx4Ec+d9
QM1KKstQ9ZNKQDmyEeImpWE5dlFsmEK6wGOhqiyq7CEDnR/YOL82bJMX1eJ2WVh5
KN8ngm/IqNYdayqLJlpAwHD9TMWQ8RjxOHijxI8spLuRdpMI4XerbBTZ6Cyeu6fy
WJjIcCgBz44fx0PXv87DdbqurRiRp5zaI4MsorjoR3GoFRUJ9b0WhP9/J/2jy7sl
+cxwAPxSslU5I6IObCSFTJGHOPVbNADZHsKzttOFQ7JWaM88edOAtzUPindJoh08
z88pTTM8azdfdy4T45K5v7DWXANe5sReIzO3XB3gZ1WqRR5rNZVTNc5Cro09J9nL
fXhQim2fwbtE8+kkOh5fZnopuGX3Qq30S+ocpnEjd3rIxVyQzn3H7awNywzr5ErD
tskvLsaVRP6+WIVFOKgjdVqOLLYHAS3YE/XjCZOTl02NLWgj1zcmuBseBFPqPRCs
KocvTywq1Gp/sG+dGvmGFP5G2sQfA25cnNve5priBoiIoe6tX8gKiip7JykWSRtn
D7Si4HDTNaruNfX7rbf2fl0SoozX6sLr04QyEa20E2PTTx5BUDjN/KMqzpUOqOdY
JsisknWx2DZiqzvY0OLVyE0UWi8zPxnvphD4kpSSXmppTVYYUjMaV+DpLiFC7HjP
gmiyjU7+8CZ6hAYHiplmx72ewP0dcOs7GU3mEbLjZXxxbhQgeEjTeXnZaCBWZcDv
GMgZQt6IKkLLB1Kbe7cthBLn2SirSOsawoTP1aMc9fMFhdCRLI1akhZWnf6q59uc
HZOd1o+mGH5NiLSbtv5WVpL5rkcz50dE8n/3yWrLubZY0e37Ft49Ng0TVqUtVp4o
UClmCaqWS97DyD1MHa7g++rksqswMya582AdA77x5gkotaE6eUVIojbISX8bzDyg
/5HLH4isuAVJCql03wbCLDavzXHTSkjy1qLAnZIaXeCsmw+DgzVoZHJQeZrOmCut
kY8Ja7sEdh5FDC1wY0V+M6UMokNdU6Qg/QF5+zlU1tkHgQD3xdBLSMQUXRy6EM6J
x+zzlJ8wcqGpgnU4SEjCSm36FlkdONjRpIvHKnpPmHy7sJt6xBsXwpHVkIiHw8ty
iVo0pwAaevMGpkaG6/qELHAnTvXr07V/z4sQRagoDMobv8D12ocwNl+58vQIEITV
1PN7nt22ZMR7QrnSgJ7rLDw+53j+m5k2M/o681/EJg3dJZ4hNZK9QUm/ne2YxFRI
wJSe17BC/cztaejWlnVbBRDw6YkYxaVV7C5DrjqCWszVF/PJlczad4IQvE8xD65n
JfsX0T9UTAoDXOzT5N2ctT0SypIWIGR3anvJluoRkpN57KebAEDm22jNjHv7xscl
RXy6vGPkdKAsgZv+Ox3qUZMXMVxY4hrtDv9rje/VeWnSJV1K94KhvP498+nAVtZr
4LpHKFewhn0Y80lQpPQ4sxCD4XecsdGreVwcfETGL0WDHdd+CzTYsUkmbmR3OZ18
+nVLCBK60AONtWSgZEPRi26DMVlWD5qJaUQiaw092fZPikD2P7jgc+YqvMCxuPpn
6/rvEgSpum20Cyy6qRt0NDQv7mQ/BaQnLmxmXEEMp/QWmG8JfD5Y03VGlxNwgei3
998RHOnK16t+y5JxvusHAbQGAmEW4SA/HNyisCJayVZRjgQI8xTvtCyrsz47Y0FY
eXydpbKu3P94zWSfBztfj5IbQJ+ngFOAoHolzEZzQH95WLbyIxD4EDp5c+kq+Gcq
Yei/E+a2zQMMhoK6YpZzb2H1LcNo/Toa0aOo0qa2lFLWzIABIUndERkn+mijLo+F
FLHLO1gReNSMo5K+Ee1AWTbEj/3/zNylQ4autDwZ5HohZd7SV/nOYpn+gQaBK3op
zeTH6SNTY1LIAm7RWKciv8vaDdy6tv8qbH75gspYcseSbO127s8NflrSO+3kWITz
/AyDq+eUmKFiGF1wbHYM+XQgTugQTNMRI1AGphtyNKxuUXHdfyLGHUPelke8fdEY
0IyCame1I6aIAgS4QRD4E6r/Nhkpp6S5ax5kd+qJhM6LYFL/l3glFeTLxa9V+3C/
pbBD7nS6iRr6uxA5h3wFX0dWH19bChm8MLsMLbSZHj+AAoT8D7m3wTGDXnv0Yh3T
7li78hIIxxghfSPWfJGjaCKQfD4/45Uz7bpcCGe5ehUOsmKEYmOZ3XOB/jIf1F1R
Bca5D0Weth21PlFI5ReraC+FthcZi5SUMchFd0VSGdwi0k/TD2OB/xl4fAH2GHlj
v/R6n6PmMhOFXd8VfR9cbQ8xf0f/2cbFhCiK1YBipDcSs9m+NNhvQa1AV0gvS4BJ
3Aet11yJmmVqMUXLbYAVQvvuBhejsdYXonj/giopLX5xjOn80wJ/RhalHYtJEyrI
we6Tst8uwJNcZ1v12QHKapqreY2s5VE8TFXBXuuVa4eZeF5bKPrwo9WJU/2nWJsb
HB8EaQAgUHTvgaIaLa6WRliCXif12Q8HEB0OVPAhfoKnfZVSYnDdc2wpVBII56ze
5l8pZg/KHniN5RsSe8v4169qW6Y/ezMfIAV1b7TjMv/OYJYHtaxkODerjFG98CNd
UGDNsNtcwrbf/N5n7oVXig7vF+YjbAAy+y3ckypmj7wNdKT8iyP97n+Agvf3Qa2c
bB6WL2OKftma6cXDjRBefXBthx15S5ypQdWkS9hLkpqAvXGjsNagKofUvwsrkTBn
ZsUyZN6B5x/Nc0YcKsNt1vZzVGcXhrAd1+1veBCumoPSE5XJKYorOzeKhyfJFu/E
TAjHfesNL9xkVNlCPsqRlwIdbN/gOKFOEamjNP3Bx0e7G0HTVpLqiYhp/+Pcah2K
zTWGJTwdbbTbykHXVaB2E1aj2BawkYoFhZvUPHJ9Errj1KX+dZJ7D4eSGWP1osKR
VES6KpXMlozIOj9R31X5eJukGCB8e3ux+zd9GnVveXodyBkilaP94j+quEbQmE5U
JIGSz78MhwpXKsMNm0iv6+7jYDBQhDVDhkWjPCjcADYEf2qpvel0ujQnCANCkTlc
pu2B2pkSv/e4IRMbcMNqnVDP8oZVkCf/FTV6qhApN6czfqDlL8S3F3DcV6yaWihV
8lkX8iIzpLdNvtF7IDou8W9pBne1yMqkJxUPQHqm8th1fVEnpFpedDUpXgZmBxmC
ggFRgHshoagM+qk9pMBdX7Zd/qQtTJ7gtBZziBqE8ybtecNziv6XAaDdLYSp2LdT
FFxCBNW7h4gx5QtOW+QLs1ZVvCU4F/1geuIUVDDYZ/513JxPrE1jDeiKKnk15kWs
x5WbMRqCDgPrL7V2WNO5NkpPDh0bQebtoeTX/aAseiUZUnSCl3AGUryzimQy/V0m
UZJru0/5o01wK+xONdHzhfIgNmqi+ogx0S7Kj9QL1eWvrGYso91rcxVlQBuSzcDt
YCtbo60T9y8kwoGoGsRcKFwbKfjMeE4NaPBDelkbFyiqBAlpXc1SUbhxgRQ0sW8b
u4FTq7FIC5sNjeE48QKzvzMDGWv7OyqRFaLbbbQCMD/GyE7Jn7M/blUEe5Wim6Wn
m5GzMrf+lj94FnSo+OLq5RNJqDFM5qsW2lM1JkCUW4lpRNgHqvmbQIXHaPOsxadn
EWtiOj1a/6eNEqdkiQ96sqGRuKqNxmapxpA/T4fC5JT0beOiAZKPAzzsobJFAyX1
4jPQBQ90rLNQZyKEbVywtOW+fEw2fAt4E0wTGRnaSFGhohioHK6/zrxh3QNZwnRr
YtMu9FsU65UqvrSPbUHov7iVvDwxb03iZR2gf/qqtjIshhLakxRTWV+DDqgftQE2
YBx1Qh72WP+EBbtDA98CtMdSxd7EiHxAp/B6CET8H0Bbh74mYEuasHO818chgluJ
9HwD0xULk8jQfEHP1QzL3i6wsrMEIS4grO9K/NFD8Yq/ENfW9k6LGTldEd3eVlRD
qpU4+oq6O/bJfTFENPezK85RHiB+vAhU6078kDYH7O5HSCRWrx8j3Xp44OwBvBEL
r5LmuSDzN0aNgwppjy3LYskfE8hJ4gwQfOHzR5rz2dGVn1S7+l1GOOtSqx8VkpET
mIegBofbd+MkWXQFIM87655wr5dHVQL4lhjlk2GuaOOaAzANgc7r1+fdklbhStiB
ZxkLjx0nREQw5mScJCI62Y/sL6iVdocqxBy66rf72EQfKAaClujTdsAERSTmGb+4
YuGcVXqY8Np51clCX4U+x2247Lk1vQd0uRf+zKNwW2tlcmNv0G8hWhvmB95ekh1D
WqAQ4P1Q8tITHkZelWmUPWBqjucDn2PFPiL404jFskbaD5Sh4S+eq1o4NW/3GKgl
8/NT7DzhRKgFyOdz7hj+wPqL7eHd3yR9fNaki0nnCPyrwQdVQEOxAwjkZi3ph7y1
0zDjgc5S7A+PodHGsv5h3bposMTHREZCNrWuW5wXdINfV/rvSxQ0nwkwaXfhbhie
rBhwJC/VJzQVbQfTy0w8d528bp7s5DishS8e3AzRW0R5G+Id+ZoNh/cdOM0klhqo
L9BrJmqYvFD6T1PEqetdZck/vSFkWI7Fcm85bz8jFSn4hLvh754PGMnVaNuwxglq
tDPzz7QHd/8fwyYhfiUSCcMn+1uesO/PPNru+f2Cdi1X8wlK35bRzMvthVLwcegM
toQ22u05b5N2rNFP19nhZRemN5emmN8dOoDsMS2/qGSiH3wAo5WCYYaDIiPdlGgJ
l7kdWFopTvRC3Y/KfqWM/emHDmoDSbe7NzFD7EWXrRGgWRbx39nFwOKwaeUYGTZR
fLcqsXgIubhoKsnrVQXXL66ayirth3bzfFXpHtu1tPgnh645oZLmpBWB9DYFx9di
bBpf4sDNgP7oZ7O5YfTYzftKbBxNr+8XBbcg3nI/+7DxzzEaAw54/ZoUkZTIp6st
HBuYW6XEhs2Tx60xjLHD7Y2eCsaxkoXTxZ/uhfIYBBirE7K7XE8G7XC5k7W04XN4
ab1fExw4ew+hXFOceAo6bh6Y0CnwaUsAG6k9uzAAusIfkWz2YxL+CFDATOnRI6Pq
Xhv92+jQjlHgjYtmh68vsptqrY8/lLZ/YAfyt4NN6aMko0qtqhF7Io/74OKlpurR
r7BJYv/QhYe9zdQVQmVPAGk02DIhjjP5Ino9zOnhUetAqPMpgj1OrUxZoBqy6Af9
2RBGlH/YlOm4c1XFPY1LDzs8QDf2zAoMPZ4acRoBfSxov9LHKiXvQJmtAGfGzaGq
y6lonF3tqVVIKSH9Yr/X9xGV8bE634fWpd+JSSF4hmv7H2vEymT6J2ycJS9n67+y
6rEFfb6nrt8NUa2uz63+3YuUj5VZkMovNJI4OJ6lGROkJ/DW4bZdZxKlpZXfEZo3
sUEj/wbnlAMbpBHQQtcrnz0Oci3jheZXTFZ9yJIN4C7NejSYfxPcDByvJaOIbaG+
8E6fzUSp9O7mxhjyByLGCZphfDLYUKojNqs0P92l5fo/jpTQ3szWn0bL/qZi3SuB
AXHMP4/Q78m0+8N63dF4LFaioNbwYC1PJp5Tdv3MUlE9aeqBcyG/NHH0eKJ6ugc3
40Wkcd6Ek1DZWCVKCtWRSalQxUHbDeZ+VcjSIdU/DmgV2E9XXkUHimgByiN7juaO
AcrW4ebhiuqOpqVDJndVn9fPf2D8CCwk5LsM9My3NdSoOG+x7jEOCoBK5E27nQGb
A3Iq2bkaNc5mPmFwlPNgmhOpNtP1VJ1egKa4GmKmmtw4+u0mCmU4ptim+BteLfoi
xlIUo2yH2ysXX9h0fcv9fAe4o/BlgfC6mOExlxOMdShoMHdH+kDHakJZz4EIMGIP
i+iXzptp7ai0ErSXFH9asc3FfPJ49QXXKbDo10+i+xbd92WWAndRa0MLTBBb3o4C
gSeZkYWY9cqXzxk5EVJF+372F/IOqmMK92K6oPO7MQNGVeZkAYec/CjBs3vaJfrx
VtxVvrVVBLmvZJBBguWuV8yPQs7YcKOWi3dpI4cTNvAaVIr7SVooL+uVinn7FyPr
l8YLuHY/Zhq0zZbyYNEvRjsJd8w84ocv8NmePlEg6pqLuyCkk4gkTjFUYMLFEKZZ
IIIZ1O8OXN3UDogKkqEeTZSYusWOsw1IOc1qH50DnyLa2v87leixuXqnSq28PeQs
Mw867nVyzfA2YbYHCv5Vpkb40+1Y8iqit5HQAwsmKnmEqrBvCuGvnHa5ejtHrBfq
t5BbRtHc92KyUBcEs26uY+YtpyF2NfLWQysLoNaTWGtOTWx8Mu1aQLRvdFAvOr+e
LF1XDtHolrVlwQrEw3DBp6FSV9tKGU1dgOQ1mswszJYygvLb0szKNX4VjSeg+j4r
0psvHtXda/1w5MjDXxxwZiMziKqXeooNdSfOoboeXPphXkX7Se1NAIlSw71InI93
eLcLuhsnt6BFehWXNlb3UVdFGyUw5S90SzxwJr/X/be+SlgwmATA85O+aY3aiZx1
JP8pTqvhywoDn50yzFmw+QperIwlWiwhifbRFDqjTuDnMACbhe+dSbMuExet4shk
/sx0h/6pS3WTsWLO0kTBhz6NEBjtPH3XHH2Pwv5NpfeT7GomGuELbAVwTCyJvwvv
JyeXREVDhAp6f7Z6x7NFtw35C5okp8lm/VMKkSNUafJclagaYf28h5YEOUzcPqxG
jmkO/xdYAC0JVxHQHC7h9QH29o2AZyXjYSSlTPfbfCw/i2cLJ7hIFVfrfHuX1iY+
D1kaT3bfo/a0Gn1FaAdrw/4+vBJlAnkjqfapmkyC773jg2LdtiFjOriAt2tTIspR
+DXVUnW1LKD8hnPpTTl/jWADaW9JYsXP386HqsVr9W6XJG3LJgaj5iOQMgkyfqkm
rqtnU57WREZJpbLVUn2CmcseiZou3y+903USUCvRlljCDuNs62XyEl+l73vjjj/H
2RMobpztE7z5nQOiZIA/HoktwnRd0YjfX3ItuhIjEeEPb1PMXBf4iUSqOpTUJ0an
eNSGOEZYDidG5S29KETmG7dLHbufEVnoyxa9qU4uD9fe4grNS72ZWgdXfkgFfbbT
f2fLciKjWgSEkqFxHQccEfzVeMzBSDTbg8vD796NFt5Xntpmhi3wxegy1EIBBhM8
shsCxHV6c9IcKlx7mQCifG2EWN8K3Jpya4qtviAy3/lsbXYVE09iODjL89QaKm0j
RpYmybDSyOwUdtH/AJihG4qz5p7tYFBFnFMwFPhZSYGSthjWPWncCFebt1WZVpMV
sm9V0v/Dtjiwuh4g3OzDffX1gJ57H90ep9BInrZDqF+EY8itov7+ft7ezYMI+R2F
nizUD9Yz9E+ChhKFqgj2V3M7gNg3awRjGJ0V0TzBeODYsYJwVsda8HP6fz6UXrlg
Fb/ZJobdpKySO3btLkqIfa/VPep17hE1ouhAeZbnftHBA9P5tu4Vke5xe8r1AvI1
TmI0si6dh+YmgB1tExt4XTjFcZ+YxVy7Pa77l8GL/hD49W3ID57MNYdlBggImGhj
QEeWNj8yYq5uiFLr9FFaeN3cvKqgWggC/sGz028YYSfIgBhpwB04vjduIgdYL2JY
TxOaDiWKenazMk/qC0COHk+UC4ETo4+sTlgxgERWkCQ91UwQc9MxmPJZqL+ZGg5K
n+VziZyJmn6eeONp2tK8mlRNtaPKn7WcvS8/tXLHv+bHxevjFdKy1v0ZYdy1Cawa
THUZMMYrwKLYCWXSRRuWdaevJWCacwXHsd7uW+Z9d4a74D2od0DrYb+FiEJHFe9R
ohmNzqMpz3N8moTZBB1UmvWV8SzLKnwNNNJL6inlwnoN1iR8M747IluxS5sJe0pq
JmThNU5KxNj2dxJihnYvNfTtmgAr9iXiV6cqz8CoI4mOnfkRJKPabmHSlE9Xs4yt
kQbufydHsOZ7ZjDeujmdzoVqu3CBtxYpYYCGg43L9yqzf1WqE/VgwSzgL3Q/bviL
oC3syC0i4uCpdVEc218P4H8ZgJrWufjre6lK/OQCH/lzuzBEhbx2LidEPGiUBpL9
qsgebQh+5DtwiomdZDvr9l2nYO1AX9lp6WyKQA1NTlHzCFS4We3TXl50p5i4zhQE
KtxzBRLn3YTFWXHcOGricDhTFDltcuSmS43Z/z+W4F6ugv3l0j95NGPp5p0n0xKF
prLfq71IRrqHOGC6U/7OZW5dWbyXIoe1/EIg923cBUQVtBPWEb9zw742LS1I7DaP
fTQS+muEZ5UXjzODlNuXmZu3tSo1UVLcNPxZlrnx3RGvsTS2LL9iqJMXbIjskWos
CW5ku7XwZ86yiEL3lMpiR/dIn1aiaVThRHihSq57/G/Z6rhAorIFYz5K9vJ4YmbK
0NNhdFbcGIY6qJBZKrajs/Av51z9bwVza2G6cXCOAqMSej8NmAR6j+vmIyKqdkk5
ab2On1Yfhwobaqlzjkca7BAlzFOOUXxK4GjkUk23eZTu3bXs+Pf8FGDpUSkLWD/s
LlZzMYZmvc+maoi5rlYFFc0syNBgu+oc846/Y4q80nQryeftt/HY0dKs2YRQ86il
d/R3mBNi0JNdrFNXk8k78x7Rfh1FeyqhhO4+coTJomLy06CPs6VO/C3u7R+VXa9x
WXKNIAU9jEUADunO1x0LNrpZpyuH2ARf0Hiw8M0hEU4GW7MQK/8mLAj3qllTjeDD
UvzHxOT1Nj46SJOQcIujFuKfvGh5SimNRqZXJ0UnR4DAZNKOqTIx85cm25y3h8Ax
Rykf3QbOCWvp/LENgGDb4iAaMxs/DN2X2DQEuQhUol2WE7qJ9EmrOgNdadTFjjG/
NX16TOrqb8fJ3DG6InFnt5/fN4hlmppNHskGgDweELNBtyei8Dpa2beeNZAmKu0Y
88ncYKKtdrZ13DwYtlEWCu1GmKI7SCNZO2oIdfsWyaowp+php/cz8mqvLzoZO8la
1w47of2sOffgHwmpfkbG+kUZI9XR28tj5vxmN3BYS4pP1+3YDGwx6oEZiNUcK5TT
lpgAlA6PCk1Uzy0DPFP0hlNxG27opzqmnejMkooa+WjCmsXJklIw+z9+8R4tTy6m
4yq2GMOOcZgqadrL7ndiOOaU3cUw49ZvAR9dDuN6vL3F1aUnCL62e/NmQ+ejNxRZ
oCCuRrNmz9XWnrV0Z4/oAdgBETKv+PpI0wCnVoTjNMJAETmGE5w5p+l0zJ0/3go0
TQYLXZuiOMs7buPXJ3s9gXW2d8gdF6jI7evW215CnXaTjJNQIECTI+lVPEkHEqXg
MRQHuZmeNJ20lHmLjibib0QwHfG76BMqlbThteZ9s0NnZ5XI3WMMWASWAsjfrCjG
Pb9fzeuP2P0qz4JUnA8NrNoEVslkXvMpFg3iR33LvMKFjd4hHkVR0Bd2qdhR2gwZ
MVwqn9oGXwmw02jQkJphBMCHY+XAbFbaPuBCKxshDOCRvNdH2D16XfEzXUCp2wEG
A0sjAN/9tisvKvhnttwtZrGdS0/CgJaJ+EJX2SNtRKObcIAK4jkTYSeT5hn0ncsT
9K0khXG7XiWhUkl58NW3MBWU+50PDgRGf6Dgz9tbWUMKiGS/xsnIrcSOFgZ7ehk/
x8wNYtqD3lcLpr+kd4U7C9pWk3Oc2TG1uwoAKTKJOJenc9Xv60Vgiza9YTOAOP3P
mmNaSzQEJOoyLHJyqwhksAgra6GWkU1Ju+USymCd4cWCGXL74SLgYbEJYxWNQB4Q
/NLGiQb7oIA/RSEVf98aOwz69n2uIdYLbdq6YWOarn7EtHWGlYBjL9qrHt7/fk6Z
CQZQhemuN+HuYWPRR34H7Ud7AYM4mT6tYNTFrkT8/CkNih7NttC0eD3a7GFKZeDR
UTyfQxEutG/oUuG3bYiFzJQYBtO0RgvluRxiR6j+dWx4IryPgdG866NqMXIF58Fq
Itkf2AICjlimWmIT8Tyrb0WePEgJK7TY0uG8VRpFzOsEmZpEZ4q3gMxgOHK91Odp
vV7HdSuxRWbbmDkqnDfj02xUyprvRuCyD4pP/alrUAntPeFqU6E+NcOp/ZIFObfW
EtTDntwOOyab6kcAbLjzVFdS016dIoTpe/JZ4nOr/ieRNUJwxm4g1W/GstqwUQxw
xpbWFa+Ho2EtlEWfBIlJu4mPHOSK5PkjqYzuXyH33N3eigkEea+LNgJ2iTxCwOWE
MwoI4fLixdmrRMqfhQHHGN7tLBDQ0BOaXhq3Ond4fWn8fLBbDWSajrIm6KoNQkxC
J1EtOaLZLLAoI+qcH39nRif3B/svjKshJa2h5dCFE8dI+doaFsXdLUog6IVJpF5/
THbS9Sx/7BlJ+Xsw9+tRaN5V/G8o6Ov8MiUpnsn0zb9HGT6Eq6owz9+lrilzz7pL
6Vg2jeX1U1kHYnMcn6Qj6ikC+jVtmqexu/DZDasFnxhOO4S5pondt+Y5lrgcQJbp
C5gWn8EIZNQzX6M0IQrEbRjlbJN02SDe4Uxd+M6CI6ozmEC4V5RXcPO4ZgOMoXk6
9dCpNJq4lXZJQ77Pcl1hWQ7x1zU9va2UVvZsnCUYPYUfjMDBVf6jOtjSQwfyVKlv
rL547qr6C25a9nvKm6sNTEEtgcyymjG8COR0sxi6DlZkqvIszVQg1H1hEOdl94+0
3NL9J2xzZcxKmDIbvueUxyP1rr0+uWH2Sz3Bwyf2z95jQhuTM0Op7MAQnDyZWLSF
3xfpqzfmukTPbFHnRZ8d0LC/hINMueepKToHaRE0zB2dOwcylBBq7m71+ZPp0p03
1pc6YPTF+KJ9NaLU0mBFkAZPUbkDbMkgwnY1NLOi0LlF/iVXx4KgHW0gcWMG/3VT
S+BKEHobN4WCab6eQfP/3ANIr9mIeydHDNhiNLZZY1lauzQnzu4ja5Jei8lNC7ZT
ZtupFL7sT7imwskHCxzlqOUHEZCTP4zCg+hFiEY4LuR/xdNM//Tl6yq9TocSjYlB
gjK/gN/qXx3M8kSBWoMzlxnO9BdJ+FoSNKWVK8sTRCV/cG+f4SiGmSFwwF+wXsAL
OJhrF3d9NBGqAkIG5MIShuqJBerS900ZsagTRcShZKwDIJp5cNti/zhtb0uw/wTZ
7JYuRq+yFhL2hvh+D3WcxanzGRFyUMNSwNoR0hjLDptoZru6LZWbeq+c/UWhpwh6
2uQ4PR54EPMJW/bWB88x7MqulnnWcQrDaeVH2mICAThqymwPjx12cjfNxWhJ5KSj
EmXSk2yvOqpDyS8nporqQWz8/BdY9TLhFnaBCFA74AMLh2DeG0mXV41NiWeR1iO9
Yk/4xs/yLWocj95pFw2jzsL1fOCOwrh5DSD5GGv2Y5oHV6dDBKfNWmlI4fx7vh2t
WYA7WuTE6fDfHnPoQXkra7nUs6dVcQr/I0C2Z14YwVf0ly5keZ9xnUwT/HgUeT1T
0r36rph+gNC2x0gAA73h8yXNXfOEyjYikWXJjieGa/BMMVRReBkW/9JhUmMgSzFi
c25Mg6S0XO5xbE/7UTZeEbLbo6FycKwwzgMurcJfaVXNHtLge/Mu7T3fvkpDF312
ylhV8PlpflWvvV0uHQQrzVmH7U3IIHZ61I+kl+biuPOXso2X8zO1ei0POsoxIMt7
NX6wMcu1SfYAEVEwUUlrSqz/ygd6mHG6/qLpq4/fOKpW5rCtJuEQ+1/fgV5meQ/z
G6eAc8S98RvUbtl0BYLHAgxOuyGq9g5tQBGstm/uME9yTOwtUtX0+r1otj7ayGj+
Uymbb4Jh2Sd/VsRh/Lcyh17GbhRpoZK2dl0tmxC0bfLFrZwscqzIf6PqaDWrTkI3
4m5bRIZJDvOQNJ391/C7m3tT8wEed4qMapG+Ivm6dKVy73GPT352P+l/H7vH6Qt5
sh/kOIAEn0u7x0k9tU6SvEc8VekVmp2N4jCFQXTNERdtDVib1NIZFDuMLBQiRm9x
xySTGCuXxMJUwBJsJJU3tNgOjLHOkKEh/dqiQA8MluFe6rmqWF9+RZQhPc5rL7CH
hAc2iCpEPJ52XzwYZR2zATomkywd8ALhalMBAljy5aQBR0r8DS7VGDB4acWiT/jb
i5D0glPwfMJV/xhzttfoJMvRoMwox7WyPtMc+VCYDfLbwIL9BIPsZtSC8fQY0Nwd
RZhPLmKvZJPlmvAs/k+UZnUTVC9x82v0yOz2G+pTuNQpAZkVXuydFExE/g7DXShd
h1yVRzGhaFOLpQ2TpSNiNtO8DJFTCpfG8ijhcXLlQm4nqyRHUhg/NIsV/ljSYJOt
C38/ZcY3xUei3IQFPidWUtU8TdqRZmZYsAI4XoV70UPvh3vQ8INEc4AI6tqW1LVS
GurYoV/ANjJVUEhha8Ypms/XK+CXB/WZq5NQHxMKPP41ByqLdVGTniQomSEZnTg/
IGVTA8GCTHfpFFqc6UN5Fe3GUg8nv3MjI+/8lOiY1I7lAGad23n6YgdpBtyLyqHS
1lkn90pIWwDWCc66xkngAh11wfPhtDdn0JVLQ/7lUrWIaSIvAMCtfrZ/jnq58N89
39ECdJCyPgqNpvjuTj9jiuqq3baTBVfcDdHjiAhRV4xEvoUa/VmTtGDMf2jBAb/C
UFqMKPRtXmYAF2ZLjTVeiWRh3nx1a77RAe/NAMVyQ6O4R/JKB4+XgPTalLINLrM2
dOB3Ew6zy5Dl3z+2FDHkttolyTQ2GbQwkaQFkKfAxEbHDBbo5SpYqzyhZnHaRqw2
WHFf96q00rWyjPdm/vLWeyyTkIT00b6+rAuJRxqswkqlUPsU+6uGGzMP1CRxtSv0
PE27YzepeLJIPD4lcRmw90ne96eZvbJj7PO1D1O/CCqnlg20L8g9VarC5xUCL5uF
0NVuvnMb3FDbMAl+jYALG68mZKzJ0JR++bTGwekYr/AwztxeJ1cZkK2g0j+5yLfh
WOSHWz+2hlzArit2KIH3BeNx6PmwCfDS47okbnHKKeYCcpYnetXfpk65iTvnr5SK
l2hrGe6GnSFwEWajhj+kRDVeTpPbU2sdJ45RMzaybQI0z2hm55iqP6/3OxRn/cJy
sxdIX9zMX1NkTRUC8H7oMhjSOg6Mslluw76mzphPk7J0AEdD+mzycAb6HA/KuJuA
D4Q7pnMzAf2JNH3vrp5ZUTAsoLSzLSl4onquHEly/1yKO6IKtARYRzwSoexLn/bV
+y9ANZOcuKWyYJERZO/sOR1p/T4I79ipHK0jGCDyMhtiZhT69XVhQw3vT8oF9i7o
cIeaYmFwWDoj3i3IIuhUbBIWDFQlFEhiKvLXFnksAAsntSysC9wUZYomBCBJBeQo
1SpNzDllOSPeqGzT7a+Pzxc0JM/hjMYFXxbxtDc5duXc7LINzRNoZzTbmTZ+yZL6
ZbpnWUKEJBSolyG3TuFVuNh9VIwaHisFNX+enWmqdYLbTct+BIqB6OBzXBbOlX++
3+5u92xL0WbMO95jEGbovHBhQNP2TgxZ6SRkGd4uSOj6mOsgDFS7mPcYIBBS4jx3
o14s/esNkA7BU/n6W+d6sq3ZCyn5tPMaUJd1cPexBOeIjPmIEpLGjQZYT1E+a/IG
`protect END_PROTECTED
