`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mvSH3ZFNuGEhoXyvjNRFt43XBCcauio7H6FyFjDDasC768NaQC+R0ozChKBlwxsa
YD9pfsGtstbB0qwmNHGJNv90V9jWAgDLE1R+D/e9suOTNWgziAAqpXBdjse1q0UX
aytAuaPxTDDy7O0LGHVDIChJ5FaZ3nOjBueWRRMalLHv0/LJocApWBvKOtlSvyag
xp71i70IB6zZSXqTFCqX8wT6zJVKt/K7wKNj3vjOEa9ohYs1MAq62kOLMJVcbx2v
yChwoTvQv+isGz/nRQm2eFdcIz3NNM7ZhwkyJIw4mW/Uj/oIrTY8h6d+dJZiz9Sa
gebAwqrStQNNcVXr6cacKPQFyG/d9B0mq4pzZGysF4Juvjs/SevG0kXSte2jq9gl
GsgJPYCx42z/NqRRekCYb/B84uDGbr5QJ2VbgyDL9FQray7guUQ/i0c4aiZcs8ef
xLxA0EziJImxp0m0UHmeSVtPTdwiggRbMC5zk1Xz/SMOf3sbIvV06Y9hJb/ik9zK
SyHsnWTMBA1B4I/jJKMxsf5VQVuUjFumh85/n3VUXJe3FB1IQUBh4AejGdtLEGQ2
jd2gXML/kzEmLHKc6+sxmezlheFiXjlaH98Cov0dXtqVEcE28jKdnMg6jSjBtqFT
L8EKsYpBp9G98+xr4SAou/ifDulN2PZ8hhkneYyRupMHhoi1Bl4qsNYndFv/IvqD
DKrO70AOA55NlDSqog4Bahfk+Q1mAkqDLmFJo1/cIkd4rMYwE5o7xKp8qF9ItvPo
LnwpvM+oSch8UJpO3+viuXGvXC4s0YBPnwWMecGDF70zHI4PiOD3VHi2iw2N9chC
fFniXWcQ6chHyDh8pMl5OrXHASjcEizjROosDxALg4hUr9f0x/8PXdikgKiEKIeu
IrymvC/1LcsjHTp03wXTKw==
`protect END_PROTECTED
