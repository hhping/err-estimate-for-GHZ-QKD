`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J83nPU8ITNIyAsGhhf1JSzLrk3GrRvgSF07cSlc1myMT56FySLDuRU3WPoDnWjAT
/aJLx7QuYKfJl79ZdKagGJ2Q+VUVuevyCTPil/qrq0nw9FNA4eyvrLhRcNefrWL8
6PCl3yMRUbu7PFJEgC1vGlBfLlqufuNpVA3NRzBYhJnYQ8HisBZ8XZle1cb2Rn1F
tV3vRBvjrkQg2uFwx7MYOMtkJ8iJ56wMnHs7HCMNBqEYIXIpmmK/pcVHsCgJuj9Z
jonE2ch6jhl5j6fdPJWptXSetjLzHn3AWxC19kHVt4MgJJ9fB+erFzF1BPVgpUYG
airzRvOJMnRhe2QQZN70OEKl6WikQjQcGESOXOCrVU7ajG2tbQGEujIQYGAmU3ys
W9M83NjAEp+AvnCcNzHFrbipr+QC2tPGrvLW6TF/QmILgBJ7Tr0ryoii2hJUE2xA
UiJwBDoZ7VXgXfMP7yzz3xccAX/hRkeyqC5SmAO1ZtzTirE/2RJki4ALsjNz7xxx
k1JB/DxO29rreuOL3Rkrg0ezzspUKDVI1tzuIVG8GpAo+NrTiXG8gxXLDnoDOroz
v0/AzgcBI+ij3rnpkcpmfEHsnSOoHoDkLPfxaQMhHEn6wYZqIOwTg5xJBkJ7Vkx4
4yICP+E8INdKBZa53fJsKA==
`protect END_PROTECTED
