`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4U9/iLJ3aDDyz+4D0ESqGRvnlZrWueSD21RNxx3rcH3gxWJdYdE6ln3XxJXvVjrY
quzpzg4vAeHDnrH/wpkRY7Yai8I3Z1wBkXem+ao9d9SAuQRo1m4yKPHE4Jy9hPyO
g5Q3x19Tc71UDs17AkU4vWZOf7rwlukBIssSFy0ypLPjkJfjpQhrRnW4pRD9iGqL
xD0VVgcmvVl/Yo9FMxWisJmgdXHVjw7wKMJ1n43pUutiwE+ZhdureAekyy075+tp
Bp63oFMfLH2F1J64j+T7jbomifzxgQ3xo7epsjMWUhbsPvCDYvlK4pfl4L5RQF6K
CFSGcqXDgkZPRuOzOjmEsUVAHEzfcOLwz8gV5YVOYW/FXkL5KCEqWBfqc8XGPBDX
qHOJHmPuZQQFzGFbNcv4+HlfnU9cSxQO42VPvSwlzls=
`protect END_PROTECTED
