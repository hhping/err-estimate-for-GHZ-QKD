`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dyIbgVV8avVTa1sNI70Ki4VPeWL36Ers7YL9cq2ete8n2iOGN3e3o4bd+VZ6WsKZ
q7QSt2I0+6mgq7lu50l/bVL/dxQ1SkX/XUqxTgK/EMZzH0AbUe2mGHxvt6x6+b5D
+rpP/gT/XHMs3tg2J4E7fJntJrOVaZVbdnmiyqmZbpDXhUNtrcWAxIi7raVv7CUw
jV9tObkuMnXRO41LUEs/XPob5EdNDzuI5sqOM2qFlP5yhfqRGKvC3S1sBLw3b7c7
Yb2tCzQF/+cFfECGdcO5086xpnU9dsAtqiWahJl3DG5zHl5uO7F0RCWM/ktAY535
fJCX0rIeAFfrm1Asn24tlK6nlM/ctkAGRy+zsTyfHlmCmEDkzPEaBFd2UE4VzrFi
051uOaFZhNWwmB705awYo8BanGOrXofmw4/0WrEJlphzIWjjr+bnuH6b8SfX3UZN
O0dc2qpCExFh4RpAXICV0p+4kfZ0aqsYAR8q9eOWImgdNCdHEorYp0SB/EeiZ3Xf
xGxNjnFSoSXed1QMP6EY8hB56pReJTTsJMPYnwf3uvE=
`protect END_PROTECTED
