`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hUo+yKprQBPBPslI6+C8uslnGlI+NXQPI5W83ANeuU0apSQ60xyifAzi/myP10jl
VTrnXBe+g5mtkD+97MWsd40j05fW0NUuHAFZNSnDMIqLKBD75TPWGUWpW2oax6Sa
YRR+CfN4Tq5NyPeCrbiBNy+bcssUtCPWXb9wWONT6CR8NciI0/4tgYTSSfLJNv9l
KiJMOrUaXASGtlkYgl1TA3je+lLQFd2udmrnvOfe3/v8UYXhhD8ttQP6qQGS/rEk
qV7sZbTrdwNL8s7nAUy31TWv+mW7WPlBMlEh2oyW5qUBC7oyb25Jj45jv/naF94I
mU8Or7F1Yq6ZoLp/YPdpWPsZ2zR3ES1V1xjiTKx1DFpOjyoiYoTWrripLSk2HyHN
xgPYXXyQMhELvW8JXG75iSwOOw4oCZAUxCOj43K0coKrISskfc0nvEkL+WaDgG1k
RuIQgdblyAjE5EYRRDAhs0FNfV3Hl3SLNO3Ta+2CbY8Cyn9FxKOtPMB0YMuE4n6M
MLH022RbhOejK6M+OcjW3DJc/D1XKqS9ZpvMvm7EC4+blSJ4nN2hUJ7sAHPNs5TC
W3s+te/PsCXKap5/FPfYF2hW7JonewHs/Yykis+wwYOmAgY+dls3Xy/e/wQtlhhE
S1SbSe7EQ3BKfU9w2Hzi5hhkuyDhjBrg7AnVqlTH7VfVKeBhIWD6fafl9SB4F1ny
Preu0/ss8QQNPA83xvLv2aotv4qH6nWn0p8FvUuUdNfjmyv4MuXysXETalyZsR2B
GVu5HK8zIYrTdeWOHuPAPa+h8sBA7DDC8H8QzaRODB32nQAZRaiINcng2QPeLQMs
EoK1X+MXtTTBKLrP9epLSr48/3awNutZwL+LMxKW2tGOuc0yofDvzrfBZF9B8yaa
SBMkX7T4RKz0BNAgQGfbX2LZGX60+m6I12d5ipBJgBPVHEoiZuE49tNx/uSVXAda
`protect END_PROTECTED
