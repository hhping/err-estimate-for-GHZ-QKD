`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WKHoyCd47bFYOn8VE198ZCUAL33+ohzrHxxf/GIfWq2Wz1RxTnWc98F/6Pk/X4aQ
ctnZmp7LkGp7GiLKI4gPs5SexUitm+NaJEhYtC3mqLAs5l4DY+3O2Rwd2mpJ8Dkk
VWcuodHRyxINLbCid1hXTYr8V1suXCvBTHU+tzzYRLI3hm3gLaYNNYE8FXAOoIjA
euvYRBRUXq7TQEKOn1YbdShOmo+LpUx48MSbBaV+t8v3vhLzInp8CQeRtyhw7IJI
0psX6IfKw5H0iXrCSo1WDQHqrCVfwvueJlPuiApI81lrRItqk+Bsq0VwnCJtyMaz
Uw7sCcbOTx0u6NkbDAF9reMI+lg+JfFbI1/tapCcuRti9M1gVHKsIM89DiqyG1Su
I7oj7sYIybJRFbW50SgbQAsaCFvFdUgQ8q1mD27rGtR0bU0iO4yDEhztubwORXip
kfAZfY4x+ds/lfc8c2v3GkPkPg1+foaNjOJxgrMII1c1ujC8oZP6x8Cm0MZrXcag
yda48hPf2h9vMRSlWBWHo20R1Ce/KYI7k0ZH7JNQNs96XLxsIJJ9POOC4s7Suxi4
B2Q00Pwq4jLXSYuz7h8rKtPZbGKaCNo4Xy4G3uqiwS71R5iQFmBEcUuTOmbC9m0e
2q0kj+nN6TTaakuFrs+6RFup7IC5fwNF8OymNQTgJTeygbIaiZZiDqz6ls3NsZYU
NAnLmihn2yIezAX2oa1rwH3DUJXnqgnGZQB+/ZInhQMK5DyhnVIv2l0owyRIT766
FrZ+W2nY8JqX0q+Z8vavO05bR5/HPWRfFB9cLpP93jlgB8ILIaR7FV0mFmiVQl71
9hlDgYMbAooPw8j9ZMxxO7K53FMc9neG60zXkY5NgWrZpK8aGZv5yywTzI4EVNq5
KCecZFr+myXmhO4Qrly6Pf3A0sFFBpYuCk9CcIaK3DLymfV81KLgwVCuwblQMLjr
nP1QcclmY4C9c2fWgRUn/luMRHutTaqmqN92yyH/REGNn4uMK33Jhb5HKLHsJK1w
hx/RA5Vz3M1vxdS4vXfZ+JhiWSGODmcgO3kdybCgec0l63ooEGBmBWtRxD/O+Fgc
nVS/O9DKCp2kMMRPukIwgeaR3h7xKoPfZByThkMEphZl7ZbYv1Xyz0HVtEbkHAbn
9rgqmVIQQX2fmHL9LC9acO3/k+SEPS2pOPt1FbXRmbGOIbbdckMu2IW/nDWB0ry5
hfO9Iag84SEAny2b+4KKbTRXuOwSRR1BGknlKMxTTBh17vaW2PWrWASzvGzM4b6o
T4ogDLKrngvQ1K7OxnW+rxxibmsQWCeZR/tT7q4oU9WRw+NTu3MpzwjCoNl5r4xm
QaJvwMFR/+radhonYXXIKP08Trdaz7DKiYtRGDNHVW9pKI9jhkwrFDC8LcgVHD2Z
6y9AxEXgm7NtnFHf2AcYbY7nhu6XYNYSrtPUW9e2T2JMcDuBCeaRun1mbOcyjXO1
RFX2TalWadRNA3hpIurJvYeGlmk0/lhqNvYSX5UouwZ155YQFEUv6bpkh+Ov1YxC
N5XqXsgJFgDNA3uApCibSU2wqN/39p7/Tl4WljM/mSIvvF/0daev4vdDEzJcnUNt
qRCMVCK96t6KrrE8I5TK9rdpFJZCjZC7GbKb3YWrX2jbjr0/zb9VGKVpMWH5Y8ae
bx/bp7HhRPuUWCQMcaixS49u8EQ88vIcJjzFxS2Raho8LDSegaa/GLy9XGYROutX
9PHNj0p5cwsKwJFz4yqtktd2TLH4iUqPPvP5M452GMffF40apAKvkuMz47aKkk37
NuzyaioK5xw3ITvbEKVSq1dhJyFiziS+Y+QH/QUbbvP4gQgsSB5wduo4q+SU02QK
fVQWfFqI3V7uUx6/5Q5d5A6UduLyrk0ZLZgsjhfaTeEZXipwB3xVyM7L3659E5xa
0NvxJlsz1nRWev+oq4MqBJtzVuVvzHmRNgsKYcbpgZb7KE0B77L/P24Kl4I062TR
zujTVKKtmMxJ0hQgPKciOAgdxhHi3C+h0eraPdXKuBR8hnHlwDoEXkl/h/0jrbR2
WWZlZCFpKPontMlR2jEddlKiXxnOdcQl8XkS3B9iQAu+GTUoyLcnO0VwSenE5Paz
NazQ3C2a0owltJE1BiaCT3WcFb1+XgW9kJOSgDLqC1EQGNNJrDai7yjCBrAC9OI/
ZXNniUO2+X/9cTfoEU6tl8jpjIDvDUtqgXHg5VoPTNARR3/vJcggZxuqrlxUJdIp
mt8wSjVNmQ4l2mtvhCi8Eb9guYCyLWyH+VXzpr/aZ5LKUaKYeWQxPq+WRQttiqoQ
baOwpHSMlRKKOxcn7fW19at2QkfUopgMt/jNPu6+wUAfIRKHIcZYLPVhYKQoukxZ
UDX3zvyYUu4oa+Zt3nR5WFBpEf7oxWe/QY0WvDaYg4wkOnR4hNVrAg15Vw0F0FJm
d46vmt5ed1cHXpqDLeoKs50g3Cg0o/Hk/FaRYVy7FhgvjsTWwnNBkxBiYJUxQ+YV
H9ZbTYf82Tth+UqOP0URp1r0pBsiqgLz/+dk44cPTX8EAzQtNLBurwJ6CaSSAokK
wMBpEImVKEaA9WIfMq1urzF7qzmz0jRuQ79Ld6TQDjRdtDuoEolsy+aU6acESN4Q
IJ/jZ9D9FQvrNrob364RjZsF5ei8y8OGLhkWjz3j74GkFEyimwC+WuBLKt5opLiD
NW8iN7hcOeKRPvTdbo2xE5vPrBhhnFeqwUEm3j1INdUcBN6UlmAzBCVg1DHZwdIF
x0FvpuyXR+mFNjrvoNOoJfe+oBxTuwB1srrltyPCOd/NS6XhvYK3SzsYcOnTRhF1
NuI2Ijxnm8AnOj2/+nugNzvUnAUoeMUUOT6VMnygm1m3gXPn7I1cK+wCakgHpUuQ
eoClOSR2N8ecRNG/qlxXDmJNnAFfd6+l0oWU54gVRqPl0YrknOubx1dwEYYdge/n
wbp/XvRLe+nLQ6GA+v82B3gtkfvkhkiUXf8fYQ28gIeqXriHMSnjtWPgjlJXn63j
`protect END_PROTECTED
