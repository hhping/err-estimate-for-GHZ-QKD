`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gJaxTQ0QfG1Rjnyum/hYFkp9mX1VTksfm3YQZJd882nKBu0XgTa00nssyBQv8l1a
mlvejvIsl7ByqfmtKkBzrUzC+xy6P6UEl0LQkZqCQ8dJPx5Swc8+UtJRv4In5yfY
ynLUQeKfJHuh+Ksr2TsYpE9/GLrpP8o6UDb/dO/fMtNmQ0N/t52QtCwVDK5eruB/
BwAYKR8sxDVC6DwYNAQrjNenXpZh3vIz/U1ahEKaHkq70Psa17UOmtbRxT+yszEm
gFgRhM3F0Gx8zrbLAFFeGG4b+TT9r9bQT77mUulkROskp45jmemCfnV3W+yweh5d
YvuHgm12vqYawH0sCWkMmIjLRTzYu33I+OWLBD08iljA8YMXyxSM9hw6Ui6feMcL
DrM8ADIWwg2zsger3CxNqXcJ2rNG3Nf45y01cBcYjTYHMPZ9nLU6eTSNRILNr03I
SUqHQ7kVQBVhOBo/lWJErivsZGMLIf8k7IAwmaVzESnRyCMkqiTMv1INPf1WUxwd
vC+JYdgMttxj/mrKy2P19Kt2rliwCr069kalhboQJD7aItmZRoWqVEalQiiOiT8F
C1mlilpxTVO2+uTZ04AY3hIx0RKdNeSWgvgxuR4+Q4ULalbjCO4MkAV3B81AHIDT
LJ7xjtgcjZLR2BuWQ61D8hN4mMxSqPXn2ex3N/3Msncjznj0znTrQfYoLVLRbeHk
8LNFMkXAmGANzwaA4OwKoOw+mzCvovnZyl1fzBlx1pRLfq4KswPqySUKrOiBMVtl
Wv4paB+KRG+zOsHC5P/L/vSRR6aNAZc7xiz9u52q7SS8jbiJenwTaXRnTHhcooYK
GANH/RgyRwBB5Ag7Uu0gPSkykxUoW81c/fKWI9ruFhJPrMewCbxf0+ePGc3yi/uI
l5k8H2uWJTe3IXWeM3RozapDhFTiq3ME/CI2AQW5NW6SieSUaUgUDe2krYFRA2Iw
kfIzB4QraPeL67cL/yv/E/g0A4UPVh/uocdCDJ8S9j0ofnVuV4CGHCukOn2XLAND
ui63j8pq1/zI2fH7r3+OFE+104LnSoiqweqWM6rVred2Z4cGwfz5pwSEkWArb2Gv
QHXcAKywXknCFvBwypNu0nwgiKIkCOrQ9b2lNxamyY/icLdhVe+uQoLsazAD64k/
sWDxYFO9cawlGe9SOUYUdzlgDFuO4kzDEVNe5tdl8Og49d9EYDc2rJnflVDbYmuB
`protect END_PROTECTED
