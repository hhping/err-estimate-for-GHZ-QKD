`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dA8QVeBcBAJ9St6jEpXCQ6Dd/8Z+sTHbDrk/Arq2XPvySloWpMRxtjIfGsxhodVT
/jOD8A3q9nexHKCna3p4aMfEAlJQDtlp2t5CpkrMVqyuTlRC5cEHpovVmvT5XuUN
IhXq14tH1Hwk1qRJpTMRVPAKWY1Uy8W82dKnciEV+0/fIyY77uD8hhHh0gGgajl5
TsNDk4YbJKwbChk+Z/g3nRmAehxnyv6nhAL9WYCRu1bvl4KjlU67/h2Eu2dtOJ/d
jkuqVcucZEzNGRgwWyPJfRnIwlcLOPoYnAOO2i2dJe1iLLbL7ZpPTcT5ieRJkGxg
vdbTqsFAQRilL9ePtMahWNBjTez4K56Qw6cJ0S3a2efNOCIvJNKoiBq5S3dQVoPu
He/0gxJnHrgIUHDVzMTDTQeKkiyeq209VS8vVEphpj5XPVKKLE6nFt8wAhnWJ4H+
lOVOyOH6BaIbV8OPVViA+u/Na+8NxsAXzKsA/5jezzENfohGFvj+6N9vG5eq5G7a
YlvmI2UPmKXzCUlCTYeMA+Yqm2zDBJv5NY6vR2BrX0M7CEd3F46Dvkx3cR3E5yg8
Ga2fosY/zSAPiU7w7vLB3orse4vdv486OjyMCW9yzUCcfNi9h60QH3md/hH4mhz1
VlhMLmL2jKdrCiraLqUKGEBzGNTFKPyVwWVI7n8ks9Rao9D7DmDFkQpeRHgkmVq1
nog6huL6jXC2n0GUo/8rjHUZJMTENkHclJZIgmBKcyMCgG8DWh+O7BZjwI435/dO
wovtaKi6Ep5OubxLyu1Lck+C1h088e5oOH9LIPUX2EZsnpJrgjE81Up+idyRURna
3HhKjQcl3nBq64gjHFGpHrlD7HGeTx0xX8wfjPaDtcfu3tE7bvEx8BhuYPS4DNhN
cLu1RtLDhNlTMtmw5Tk+uTUBmyfwEYDcs/FIAPV4ZsC+cDstX2Bv66TjOOkhhwW+
fguFPvt3Rfqy93Za3eVHE85m47eWOGybh9h8j/OVWVzqfNn31zv0/vS2kuB2nMEE
0vbgQiUesmPHnDm0esV/sW9AyhWbQswEA6u9lBRKqLo=
`protect END_PROTECTED
