`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nFCucpseBJ23GUGCo0Ja2fnL4sWqCzyVcePNkL/Yc6tpErElI0ylnpe1mzgtvIKq
VsLc7JKFUYqNG34LNXPXfXxSDlQs9ISZ2KnilIr6nMFUqNJuYS+DMPcDJuIaKe/k
EhLMq5hLj4U+8SGKe/nDCET9X2vTAEW2642Q6BCd/18qZJ7Wtp1/RpTIoioj2L03
1VlDov3bFBvgTcplOVRMa4ekJ7129/WPmWWVl2BTmqb7VkKiAj35yBn2ZwIEmXSy
WiggDhjoHat136MQ6wC3Pcr6e2g40zbFhCh1Bnb3mSCWKoEy45A57PWB++r+HfgJ
ZsshxcvYsq7xo9ctFnB1SJ3eFkWs1F7CDWJd5WPrC9csUbTsBv4EuCOQZRBMyyly
LOQL0pkLMQl1Uf0VMd/MYFNz4vblyZWFz9Oa3HuM9n8Ev2BjnfvdhEYlNnaXmVvI
dzYVv7daHzDNzY29XsRRV+K9nTj6a5+LGAhK1wQwDGzSU8UFOA6VX1XqMlVWM4nT
5zgQWS93Kk9pzszSB6wM4ZfoOli0uh/o7oU/kGp+4FSt/pYcKfIIJUmqIaznKmS8
rNtiXP4bogkSe5ayaJmAlH1pwIMWnOCXoKYGlq+U65RKM6tU5u0SREvfabnZ6WVb
ht4fxHhTpC7nxQnyTaOqJjMUyP/mIwOi7cDnFx1fw6W7xtdCCrVNtRiTPei9Hblh
OS0/lLMTzydBIDzTNHSXgSoZnhrbcvroo7YvyUYk9Hnxw8cFYprU72tnW5gFh7OM
0x7doMizgX/27yf75n7O7b669riuEqwKG8YjIDvpUzitQEALhAnKA2tMD62Sbqh2
UUp9QoyPbpn2eJo/VAu/9Xy2D94Ji5w0uA6ExRZWrU3lZMvAT4Uuo0sCqGr/fCZw
UkUmEQNAcfAWhpcNxCuz0b87mg3GichcmW0ABI5Wb3SvmgSttoZnIlQMvDlXa1hr
O0tgqbnBSOPfjq5hOR70FFKtEZJfzaQsOkXYQkF7exsx/8penSQHTcqGhTrrKT45
cbrUaNNSLaEdyBh0WrXHCXccmzRiia4SrF0mS3IDBCbrArlsD9IAP66xN1vnvt7P
sDhA5m3+NETjI7CJhb12MEN3J6rCaA1mB35/1WeXninBcv9JY+Fu1YlPgogbDXDK
wvQuWcS8fsATxR94+cl0jpynk0cGcsD5/d2eTtPtI8mvgNJqoy9ARBnl5JZIkHrv
TKV4qzLw4QlmXDmaFTFC6lLlXdJ272jNIWdsMDZ4ujgRWC6cvzKnC/G7HOEFOLxS
ix4QMmr78lg7ZZMMsfYmbsRrXUS1KpJuyn4qHsKLKdej87Rztzwt/tlc8oIl89di
t3qFZ8kenKTl/7qRO92aWCPgTdKVSfhVFrtQYskYe/FZb/ic48sg+OIUkbUZIm97
tCwuO1wlQCK0lAfx1JC2m4oWpK/1oy5JqWYm62BVoDYXsz0QoW936RFgyJsL3aNA
4UwvJ33d9/c+ZpgIiwhwlKzzvZWDrjZZp7+sAzvfP+t4AMykvVYrSDpSif7LIp+r
pW0gbfQrIiCPxtPcu7fazrN67A4nIzO3tOjXWSWvl9XuR+xUqSeBQaJAhCjiyg5C
Fi/rQvnCH7EJh+P4GBIglPZnuuEemmrM1Ujyr7umOejbdtMGnspR++t6h4DqBE2Y
YdB4v8eIhCkce77g69saCvaBnQG7psEGyv31ki9rd7U3f+eh6fJfnTAiS8P9DkMz
VNQJ0ggUC83lZkmVCH89FRenkaZkSUfPeXwPqIcKtval3hd1swS97vCi1JL+Nszh
dOQFwuT+Ho+rLDHoY3bMRQIGdo+zcyyD5utLlj3LNza2/i9XHTC6Rv1c9k4wvBPX
/X7EC8hwuBJdEbqMGM+x8aZvBnWQfI/BZ3TRYQOJd5YNYa3us9OftKDRgGrobQvX
B1DquGZUlZEXBUyr513J5D6RnoFy/xLnUQ02UkpM+eBhsH5+dZgiETJXsU+rzb31
lFajHitqFk0bHM06r6gK/2wUalL/uQ3VbcrqDv99wHg2cM7UJLOk7s5/Wbo8QVSp
8dp4A/D2ZmpwzyLbWfWPNvYafqLjuLlL17fsJxFNJ+SX5sMMmj14LOCrespOUFWW
V7YEEwOqDAvIHlr6tWXdhk9niozdtKrvhKBYJ7RhIlQAk+/nHpjOa+OWVrM7QJ88
B3P3Iwg9ADjiJH28k2s1ZP8lxBwpI8eNRKPpQqGpd/C+i17juMQDOjuDJsUdhupj
JjbJkRddO7biDC+qpgo804CI98ufky1EmegjZJpG4QkWhj0OYA1eW/ku1advKFsM
ttP/y4336my6BzznQTJFz1CFpJ1lUKbllhM73XMrkhy7SNUJbBTDMc3X19Lrid/g
VGMZHvKOD9QBRA7em+Q875X90FayGJJX8hdKNxQ2kgo4igyozG3nhrRu57555E5e
7JsxcY7Pj3fALAHwOuSmVmGq2LM5wBa33bKYrKRZEQMbmZI2OJoK3VC2ppkATVjM
ahmuCtppBuaPSVPBn2CqR9RSNEaaVWXjUGbCcVOyiwsnG3ySC6TBq3fnmsu1KB9J
kN1NhfQRSWn+nyoTqYoLinRgvtHzBFHeMF+yXgG3QwGsbAp2cSJIj42c4Z9ryhZd
wR0T1vIoWeUgTvynpxuLOHQk94fppBaaYQwVa4qKbBDYyoK9/MhZ46gEC8ojQbhs
/zcM4yKZhMI6w3vd2ZL8YTiQePvBA6v5yG9ANRCkkarkr+YOgLwdhMDIYtzfRjb3
Z91+A4AWKI1sJCszmKJ3YX0lMWGyKC/d0a/wCj194Ot4nFkNvpx/E5NkCyQc9YHn
4ypIQH57vsTL4P3HJXeFL+1vnBIyVdNuqSkQgV3o59wVXoC3F7VvzkH3lZPvFJNW
7zwa30aSrrrTqT3IUnFnl4E6ac22yjd2iyLKn3JlEEY44ZnCi5i4CBvcgSiD+pkH
IsapiQn+7YDA87XhyKaLFXOeJ9PQtv0+k9OrUPwWyNdCUV/r9lmknGf90fGT9xbe
b0bz/K4p8NO37qiVKDc5REV4rjMYoFo/tzHFxfAEd/OTa5+om+cD3LLLf70n//xd
bT+zY4zmADQhsm0f4jZkrkRKJeN/5Wnsv9bt38wk2lD3/+VZLi/WgISwl2riCUwD
L+6M3iJB3KlYISsDMMFwq+X84mUoAoahsmgeI4B2p5O7j47Iwki/XdFBf4r+08QF
vHDUm1Rz08KcLJjMG8AL7uS0VF4Ms6ZV4rV8ekhFneR4lX+/U3VN21g+diu8lTDl
SyaO9U1DoqoemMX/o4qCmx1a8reYLpR4KNcrKeRVFglCQDehzyV4YKLR2KEa+v53
mWuI4V0S9JWHhl/RkjSX/yL6JPmvEhQORm7F9xMeCbVYOXyu2NpdUGAY0FjDmaGR
FzQEV79QeiNWGYg7TpnFkXM+iBOGfr4yJn2mnqSbp8dfugb9EtJJEejli5jxegfg
msORbLYIDqH89/FeDSk63ReKw4+gtxjBtj8bGlMA1oZeIgIJzv/ydx0GjZ0EusGB
rQVIT5+XPO4d4+KLe8Fo8OXooUzRTp6e3oUO7CSe0Lbaz8GmtMb0vFWYe0U9IzC5
Avn8up9HU958CiWovyZrL+/2l4r4gE1ciIq/09dnrvKHCVg7Aivfl9Yy0Nh7wIC8
X7UfKZbsYEwCmCwDzk0h6qC0wWDC0zyETKzTW6TRoLDs+ADG2DSpa1s1WjjglfUg
ESDSDDzCL584pvt6/jXm22gLkg1bB0JFiSzkNaELYbKRmhbYCbBcnw9jcOE9Ml8F
CVEpXPtOD6Ku2XuFlJ3lQSMzvpS59VplPSCMyVg38v+T/kgfHoHV4Jli7t32JZh6
sbtSFc3msisD4vYgjMYWtJMu+yK+e/knEXDybU/HN56/y3beUMCfo9hbWtLNDPnz
UU1TgZQa588FzY8EY5kFczPEN9LJYUBdW1qx0XsUvZV3oJvKDBh8JvsvL1dXfo7N
b1vWsNna2WSrUkeEMxYX6AsaatEi3RBnB5E8Spq5A8L7c/LgD1+aX52N4fj54H7q
`protect END_PROTECTED
