`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yj/a5opB/IcMgdMqSIiLJ+tIeBZ3wY6okYXbv4diMMXHm8pKb96/ZeLXQwGfrR90
ZJTMhomTPhTq9RPwBnqijPxdjcY69ebLJCaBB5m/6hvj8pWlPU2inrHdqmEnPWqE
AZAqBUYmududFcIwob+Ifv+dKdZjreRaXOSyokppOMk2FaUUAIyfkgRnAnQGAABz
RTAdnvCZ3MtOMJzIfht6AEdW0ii56y+OV86JFVQ2maOErE8NBww1Zcj36fVWNmv7
qUKMxo84mXBkKf9BZXlQN1A2VIYU1xkvgOw5gvn0hr0x0D5qHeHnpUZ8paYqCmNL
5UoJooEAgFXD9zshgArbDyS0ww+Dity2JT7rB+IKcQozgfZ4ybRlavp/CG4sighl
ykBF+GzCXFqhilm2JU+BpcAx2UTV0Q0k2vNjoJ99GZDPFDBdYrTLBZpSZl3rStK+
F1TH6AlKsI7GvrGHTVRvkja9m84iovVOkVa0JnoyNne0lg/1ZtAxdL+S+X5IfsMG
`protect END_PROTECTED
