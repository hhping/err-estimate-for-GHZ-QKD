`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p069wCV0VJ+ONAQVgE8Ir12ShUK7nVJ9irWjsKsB0xKiW2FlAvVDK1HheeX5Pyub
D/5Op0q028PShLTr+uGMNOwtlM2QlNAlAt+F9V4+0IPITL4gWquczhyixtbPZv8V
3royBN0XfclIy7zqNrZUiSFNv5xf4CINSKhOzhSCyjKxaRUIxA4vPgS6ndlS10o2
tllNZwBU7LVavcCZW96bJ2g2/nbkthVjupSuc4CZD4xe07zgPeTg8MXvjJSUwSJQ
VqBLXNqBfI8J6y1sF3qF9cGnOV5t7pBpgaanAeLzP+unNPHPzNm1zF5e8ZqayTGb
SFWrKkyk9W/RHo5ANRAnIOdlJRuB0iqE4emwR0NBqYCfS/y0Aw86rUTzB22JTqkM
C7HN5qXXndR0jRXus5cT56gtpthfDI6EHflYtclnrAvZNGYD35FQ7wBiGlwOytin
tYiI+ZbZ1ehY2l+fBAPNsg==
`protect END_PROTECTED
