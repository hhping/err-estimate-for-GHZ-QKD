`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zB6WH9LdGBPcwdbiGR6z/pR7O5BVfNimAPwkFIMswyWvqVmN+Ptymx44VKMF3gwv
hxxz1iZBnruGHwh0whPxPnEtew4cLdFKGjmo4rsK2L/3qikkaYDRqX2LlA0uwuj5
Yu0vIwEAa3m5GN/qylm5fHBbVFMcNv1e01wNXYP6gfFcOwHTGWBMrQp42QPkxvDt
F297YpirBMilBgqzIfEVxdDKQca/rgshTRJrvLDM9/mtFYRRMEvStlg4RAd2a5uJ
jEA+9IcAk5+w5asIVQk60LaErKz5/XufU9/jKkYZIpYeOUhjVFXfzaSQZvTZzPWt
XIj+UZVl0fV9vCEcvsJ58b2mChCcnlb9Fh3tii0Js6kI9+UpCfC4zCi/i0NxLOWC
VETx8OLidFGC6phxJK97b4goLdK5dK0NLZpWkCOZ1dPDWjQnNs9vZrdarILZ2cW/
ntg1dJX9czNfgHYNMh0vLQ7pCiBixhrY0RSIBtRWSL87xAnhEusexowfh/unrOWW
DrX3go33DW42o9pJf6LiQOeBTP0dkAZ496eJHVNKYfzjKbFhWMY2YOM1tF5aP10d
xG7z//uawS6ZRmo041u4kmdQqihJJ+A8LMthHe+A8lLi/jQZr72ZgydT5DsCGnS8
CNQRw7AlvcbvAV/bXYSd/LpGPynxqwo/eOMDBraMQu8DqRZCjFiLbGC7b+ZwSzWZ
nKsEDw5+baNWoOu9UsB8CjurC7+sgf+3pY4QkvuCgi1+GHYo7jIX5sCfhMF3FA+p
Kl6u1OX9u01w7Q9W3RKFkU8biXFTPx8AA4VdiBwuRP70Xc4VaM6du4qEuG3juwg6
XgiyoCz87sBjxFKDc0GSgg4d4D7jy1EMXNv9TFxEvXTEFL6oy0YB76iuy0WqwQjR
PONmCh1tOjCkeNUp22agaQI3zKOqrg9+4Vd8CL7CdAw9Gr5QrVIDzNjjBubNouVf
O+xn6YiksLB4KOZWDSl4vhQKUDLSjiGgjiCdWHoG1C8=
`protect END_PROTECTED
