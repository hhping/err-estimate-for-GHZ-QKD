`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OBLUyRynZSV0WHacFvc8uih0MdoyzrrhqU/qaO2YZSbb/C/G5HWjcS8P/Pw06Ic/
1OkRTI+slwDalpE4ypKxtuNsU/GIc0NadvCXppGfzYjTqKXTHN1+rK+eG2V+GYk4
zcl9USg15MUp0/eXM2d5GcQZvx3oR0+jVzLqiarW741l8w3ojj7dThqjRMzMjIHN
fCJOzMzalsLRLV8Z1wTejGjDYiGInC+xW30ubwgqHNachLQg/ZzIX/0i2NEq3Ei8
yt+K9XrdCFz71TgcjxGtr7u/B6hyIVK6FLdV3r4bdzmL7M9pQagX6nO7gGKNjbK+
FUgdaYcSV9QFSLmguYm3wy9Pf5vJbx8nVaFJ6SSneH6Kl1NOav2l6zWCHnkIYuND
ZEJEbe/yIEH+Y41KLt5AfA==
`protect END_PROTECTED
