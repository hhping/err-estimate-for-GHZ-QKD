`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V3kcfG4fsoWxuNgeQe2bxrwvQkNIsN+zOW0BJdvISMo4lCj/nfkJdsgtWxbbPlZU
2MYkfku5VPcqrrGSuYcLV6fkqERan348M7lEYvgt9g6RDtfSyKIFoKXTukZf2ZMW
EvjGilqfKu5Zg0/ItNsGm0ANqKEc3gtIyZicpxL0ZBOKx7xlraYC/8L0lz9Jg949
3xWEb2xCij3xfg1DC2ffIuyWUX32caRf7hTiKoWaVGBujiZ38srYCqE53Jhtu+N0
0JtCpTxgPMd31DcQL51ii4QoKjfjlA1YgmOCjQOJRR9gmDWJ8Jck1Fa1FYH7OO3W
uqxh6KuHxKUFObwIlXEWjTYnv6q0K1w/avEMoZsD0yuEvCSH+MSSbqF9bPaRmA/M
FL5Cw5ddViXRqQWJZUs70ybse3wYDLFQMBgyQGgXWmEfeeIq7BdPrm9GFCg3zaiI
Gn1tsIHzEqDqCD5TPR29kiXigVBcrTj2gEky+X8oyRpBxNUAim92GfjDHI7bFtim
2N2ESM4RPnlR1n+6c4V0XcR+wK0U19heMt2AjMIsZtFUgGErWtHVg7V20NiUE2XP
NAHOfr9dXNszDw9E96mEaEB6qcPfSIqgBMoYR5E9Kb/bp1f5rVNBCjX9kU2I3Ce0
T8vGdKzkxCZ4lsdkhTeiHdFEfYuOdaTvjPExUJlgGAtXuZqzQ6y7R5kO1nLG7poR
h3/7T8k5Dau9gG9P6LzrSHCySn9KAjpdGphBRa1XTnhpCdsAcusEkxROI9AWQH9V
Ehulapkos2qSwMXkUUpxK3PtR+muc9KE5WtBadLZ/NsUYNywbt+sv3UpDalTG9z3
jrCugoZUbStRTpfoG8/JzH90AYfvJ87tRzEOuXe4mQc0lO5Kprv8MP2KIS1ZdyPl
7fFU+CBZF59A4Cq1DMchN+3Gp6a+adwzswwaV/8O8tVRtpYsudFKKP1zeJ8o4Pmo
FLLDtNrz0KKlIQHCvWzF3Eiis01Q+K1AN67hgQm7MbzQaIap9UUCKifSTXxNfnvR
WglZxmjnsexv+xOgbDli/hDStG/EJJghTBYfRvM9j6Oxal/ak/hC1WYIIIh4AdcW
uDALHiKL7o9Pz+SOtTf2kYEu4jb+IUdGHOjM1mT01XmiKeE5rQes+vLc/e+URAE9
9yNAIonSJamWtaNYjG6KbD9TgtHDmrCJEg7edtwFRkyl5gKbchKR6Hz19SL0rls0
npAc8/TzUD32x/+8xiOavoiGLc2F/SD9wmZEWkNag4M+0KIiHGQD1A7E0B+YzGv+
df3fYjE3FAXkD5JduoyzhCOPQ1NgHYiJ3r+E7XWwk56YtoabKCoCnY8T+2bDAIIk
KZImZNdP9w+eGFO5KT3Kb3luJnuh0pCdQg30Y58zQ7UWhZwGKGzau8xOGTKUP0qB
GhPs6jPN/mzhuJuvTqCDw0Xocy1hU8Gnn/kbPWZJmj5XdD1nUD/Mxzr9nleobD1n
rfQct7dQp4xM0FsiQXDSyWYYaA0YKBw4aZoMbCPXAnE7ikjDTyOaivFYy3o0kLdi
`protect END_PROTECTED
