`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8Sbz9thpS2sl62ck8HW3AJzfXUR+L3Ax04THsC5kV00XD74qceSsYtbHk3OOoqnU
bxUCOxnt3yffTOmda5JAZvfO24frkYXgZ9UGPHdSsfW25VTEuAjU+1WKkeRx2yI/
yFGLb3RMRPyzcNy0YCVtROYrRubWE16U0cr1zxO7zuHBsL40YvRPyUeTkInWC3VH
h6eK1TNEgxaP0qkB6pk6HhfbituP1NvxTRQm/phBGNUiSaakdHtCCdPC4pKd2/vQ
UDJpE0TRM0c3P4R15OuFu+Da9d1udcZ20uqCkEtNAW9Db0XzQEfI4W857f8WmII0
Dpdz5Lj1AwjA6se9403jdVyAUdO4lbyJWPfQn4dqnRs8YVp4FBkB8lNYnrujS/P+
X09r4Jwf8nNutFXaEo67oczEV+erkpaiQd4kKsj4yTLdfqVdXeklrPwteJkkTfRd
7MhX7aSbQYiDdABR0AKUg9ggbLh6vaPOhh5awVe6/CF+PBP7pN3ftI/H8KIj+jyx
19pbgX58Ew3vkeE40OcPtVEXoWIBsEAHjSGuBIekjcJAIyvWPEGkLAJ0qz0dwxRC
Q9yUjhN4gzyk3oiSYhvIzf2AxAtObU0cXRX24z71uzO9oGFyGLX6k8GpRT7N/NUJ
u2GvJ76iy5pgIKrwiw7TKal9r4dhSP5WElrtOS3UtBJkq2tOhwxB0SPUJZfD3Ao0
RfL6OhomhNgy8XiHaUC8Og+U35Yu2X8X8FBz6mDiRmQ4X18oFfzUZu/h03RiOnta
O+NoxCgSpuy5ofq6jlYbxnIL5cZvTEcYmfnTBZukh+xrxmiiSpM5HZHz4oKfWuq4
hJwJC8In+hVFFs8yVu2PucQ5gQPlFYUp7KR1MZYwMvxUoGMimf6BOYxtBFMNvV8X
jsghDymth6UkDQpDTg2AAIlEbGyG774m5w3/ckeovyg+hi5I/ANDj+/duibqLU84
CfvdSyFQH4WXlB4OMokKbQKC0bU/E2L1sJpUvfOo293e8lQQpLGXGIWSCsWLPjR+
cQr4VMEmOUGJ9XX1dNV8qzVZ+yM+CwgBaSHrb2i0H918CGTXH+tqmMg8TrlsasoA
2YQn3m3p//U11Tf/RQbU8sFN9cftPROsSuNSyhhw+QH37fbFjkcqTv6PuR4fVmNz
vuseNnaYSzF8XY279nnI4Z4hMLxVDbsimI+pMIhTA+A=
`protect END_PROTECTED
