`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xz+O2+6VhHtFHuzh1Ioz2cC0GY3kGqGk3uRxmQIg+FIubHiCwbCD+nSVbNu+SFbJ
EMwRyQb4/Rejw0W6iO2IlQ5KVKANfL0dK6J5THXjuBlvdGGJzCalEVrRV5X7x/wT
mrOCisSDu/At1i/l9dXjPwjHwj/aTz4Ff4nDz34qTeGMiTF/sjyEtvMnSziKhLcC
9KxYzoNt4jHHyclQWuH2ECO+PyYwkW/MZ/Hb7M1PRNwFfo155buYi8n+1JmUJD7p
4GxfzUdGv/qxfk8qXcmBqv5okBp0xneyg2uhjKhoxolifQppqRw+bVuk2Ogap8PF
9tcCne8PpcDvvlC1wxps6d8aCVU8Rj5tJ38y3RhcLDXP++G/+r4pEU/wnMC2gBHW
lhTTh/Ki7a8vuqvShBsDOc9+0HAM2roQNOiJapQs0PQZ5tOAG2Awa2m/Vaqo1dNG
PHAqReUP9Q27/bZbbwCATIRRxyvIgYdg5sNoFY0HIYAg1DvOjxW04ATPwr8Uy1FF
/wMeSepXbh+PUwrGud7yFAtVaCEl2j0VO3fdwP+1BKRMX3KdTLik1jzm11DYLuLl
G3TZeZapxRlY5l2UrySnfAZo16KeIPr1Al28YgwAuW6oKolxRYa/ueIW1Y4HgR4y
v4ufpVLdTS89jpMMMkMHDBsV5WUoTem9IhtzvLfjWkicB45aoXSwypdqse9fyiv1
VZvaJsnUGua4TH4dcdtFmb80fmMM57PEOfMFargOVt/EuePWzIVBmBsn9QP57Qd4
3aFWLFNWmSBrUYPwUgr7/HBt9oV7QXvYgo2dul/sLw7rz+WmlVDJSwBTzbbMIFgV
ZtYTLLDwzIdpYhk5E42IKVB+hU1Qi7EAiBhYcE8UCQlzgWAXJ6Z2EcpXAhAEy10l
vo7LsOO0I1wgGBTxYmGJMnRtB49X4qYXWPTScTZu+ROy0m5lN0DWvn7sRymc9mfu
8eOHGFbzXVNOW9KcKvAclvUdH0SsqVNpB+KDrto8OMlqEZZH2UZWRPDfoM5YUrIc
br1ck97A4xUeMLRG99UC+MCef6rbveiOCbpl+uNWg5ha6gZZPF3X/CT5JWJR5BDm
GofWKtmeSuYny4VsmzaxUTMXQQx+p8hAFmIVqQcZy1oQTOYL4PnknMvpKdcR1p6o
WhR5FBkb3WJ6al6HErxSXQjMxrZCmjNVQUm/AXEsP8SY9BnZhp9SRXFK9ZSWJkO8
NLWEMfdh4pilS9B/ByCrTLMR+kPr3FbmoMsH3mDUPMfVCDd6HmU7vz8J0Dep9eTe
RVlQ+VSDeMg1M4ulBL54FkdTGdWiIWA2gCR+OPuKj5qEFRhRXKSGQfdCj6pFYosd
wJu3oiMTb0pg280flWTza6dzPJLBWwrVEwUUKVH2XWTnFhsmCaVbbNG9sp1JvZ3b
6Zaxvg0fETD+sVO21eyvDC+Vw2fY6nh50iDB34DTICb6QmedvcU5ahTPPk5Lxzx3
T3dIYYM0f3psfd5Xs5jfblDJOgKndKY/J19uY2apQCrLTxiJPnQoLh8HCytgbDao
H1nsO4fNhcM4eMu1bfx7Bk0bikWvSDtwIF02SOby3Ht67D4Nk0PK+GHcsFTWQNBU
hPtdJy8XFg3PRZQGqVh+mZAN02LLJF3fw4NsKNME6h8IGZQ7TywS60HyKHLisHNl
4a2YUeCQ8LWWpKJuFTyPEYSHsITh0i4dv6wDF43y60HuYQQmEJTbprMcahsz+sQv
TcFaHtgRPWfmftGK1Ro5qvCLm2RuUwqRiciVMgisvFGLpTxHl1+B+m0N3ezs2w6A
c9b+J78E4b5rOYtJ/odI7v0pSnJHPkyndz/5xw9AIpbh3gcaGAMA1hHCo0SVFDsI
w6BFlptWw2jNW4AZLROXDdTyGWkFkCysioadbn1erXtSkOdyNtloLd9UFKhh1TDK
JDZUqMnMSZV1gwJCgQiDlzNa4Wd6K8CsDhsdaHNk0BmSdjhn8lqVuNL1opJCccf/
2KKvDkVIXFFhuY27LBG7OCFoK3bYZDYxpHuhDyglNYB8W6NwCKet81SQIvg0hydh
oJb/8eoVk+0c0mnMRCWHdARtvZnE5HbX5sOSjq97cAb0h+GsyLFglZNcsAxEIpMj
0wAZEBMTd1XcnATbpgiqqkViF5/dPGF8dPdc+CdMJ3jbZqCysBNne2hFlEgNX0X7
HyMcnOF4xngdJL7zVE5Q3Bk7KZ+jR7hEO5gEUdowZY0rGFkM7NmzbHpbj3UD/0Rl
zPlvucGAtJpywo+/nZiGItaBJk5hNfOdenN7UBKgVXx4+jnemWMKqn0femHCa1Vd
b4BzNDYM0yAROg9RYQPX+R71ubrh+5uWQjARvDBcyYewag7fvrIQZIhNN21Q6oKR
3ul3Ec9Drbm9DC66PmdArZc0qBDH6cD0qzYJ3uZmb0xWcx0Ho07gkb0SQ9xRgKvK
Woy+ix2IiquDzuvoBc68C7Im3YR7XJN2qkWaOr9qvR8M9K+A4U/HXnagFafkoryc
7+/tbEcw6BHFZAa1ZHP9cRdkblY1Z6GL+9NuEdIdu9+TSpDCBErVVvDIQv0/XO7u
qu8q8BEazjrwVFT4nBEgtapfYENPZl6gHmeF5ux3eZBTvP25qghgX26A4sKXzNlC
5p8Ug6XF1mIgqYtL/tHkU5ePIeftYkipGg725uF6jV3jcfBSIBfxybSbfFfRgwY0
atbmdbdEGmqo8UFrKvUS9Axr/ZiHHTLXqTPJI0EgRxRxdnLZBM2xdzARTI79A2JH
SbZ5m8un4wCAnvXHnYkdXdB1T5dBlDcKkDbrgMfBpGvzkNbiLRlMvCm+S+1G1KW8
n+7heNeUlJLQYZK6FXJLrdRsvuegXcvxMuHTrOqdfw2h1TmmSTdf5OqS3r0Sc9du
EraJMj/NZ3WFEcEyfQBAWCgAgh14rlNxYXnUKRYGbE5px01MPf2Wa6dCf6z+kHwm
apvfDxpJDyOGUSiM3XVSeC018cfAWQpvwr3wvbJFRP+JWP9ok0RKhcv7kent5o5y
4o6f56xrVa9uA/j0g8pQh18452jMA+5me3IkWCjp+xdLDm1pDcSMIQ7s4w9eHkOD
qXWTBBEnYsG8vMk7puXnkEFpGz4KWy5IEP/vgVJIjldUxOuIM+v7fGZvHIPToyEf
M+wQ/AyUTAWOy6wnnHeE7OBWaTVIwF3jyvsMUkQsbtsn+13enkpqrWdC+sH31Dt4
Q7CpqRYmRB8DtCU8oezR2MRQUdD4orGeoHhx36dFy2xkHc5URqUpyDQBrMX8tbD6
x5EvIhDQ76DF7ZgzWZqJOhImpsS6xUIQOsarp+q/C9gcfUNeojPhmsQKIfcbyHZO
S+cKyPa5aetCFfQCviTS46MJVSnWc4mc50SIoYYv2rwoGFeJVYKon2Lid7/WfzaW
PTsUaLo+G+xNuFO5Dff8EEDlFBMdTldQS+a6Eg7aaNkL57+xzHF7tmkKzPmoXL11
uLB2wFujkQhyzRcGbaWE2CgG8dds99C8x1T8Tgn5jkYWQyLOZs5ig5O+YSScMMFo
SRBgSBn9C97cYCtdf0riE4kLZeO/s7duFjvjtQXtha9w5Iuqz2uMxGS5fQwkTnYQ
R5FgWndXBk8x6NJhndGJFaSLRhZ3BkmWQ/uiDPGUw5Dc0fDz5ZkwylFwJjvzEpp1
rYubXAixg+vKd5notYJsj/fZhrgbFDxUpVYR+krUWKSH8CS+osBTBs0kbuDih3HT
BAuvZEIj8YJd5Cmm79yQvEi1drCTG3zyvHo2rieeRLjS4/oXjO9olBy0D+7h+Zxw
lVl4HmXh16KInp2DEVDsQ9G8q/tmGqaqGpCY/jNGHaQboS7IOx9fq9J0MhiXcKCx
Bfpb8yrM/tomOCmoHP4FjhyJslIm7PPZblx5jurTmCYtoUTrZelky/5m39q9R6Bn
SXV5jYY6I99K6zNG5zX4YnQ+WxixoDRm9RPDnVGMux9NoLwYhyNDsG0fIJWN0R7l
N8V5N8585+51f4tavuuTn2odZI08uEz6y0EGLVXiCnUJN/Bh5x3x4ojyLis8/XkA
cOB2WA+uINlW6WhLsWu/r1xTlAvOy9KfOmplyR6WvLbTabIXGgN1BWDBNlh/9N2U
1WLN8bMtVBbRfU2o4xwVIgCSgKz3VzHFjvVScb8RRe61pxGPWLdsNmq2zulNxE+y
Mb1MhXPHWSe3aYhTknRy6nfelPLJmcqDGn0ywxVmB9Po4BU9ZwAU9qze1/29CjLU
fMq1VtD0T/XyOb2n7FtugHPQGT8HVSDlHzJPLgXuv0KQFumLqYEptVl8SdIyyQ1y
QkXi/vIel3sRUsQc1Lxrr76IRfS/rlcuP+5sRfrYleRixcewPr5Ev0chrw+nYa7O
35Z6hCamZRiZ1xXyGvT8WNKs2H2fFhFAoN007MoUwy8Vml5LSON+1W6kOS//JOai
fMwSSmx48w4PGOzYvUkcGPYRTFnvhQRRTiWCrwOJfF7Piqt0yeBN0QlGCDLRBVkY
JQ5a2VH809GrrXm/2SGycz7HZCwqtq5jw9bmX1+nX5S1sEh1Xyx6nuu78vh5pmoH
aRbGzf9hqCWi4gX9hkJYwyxik/OqM1iMooy/ZXBtyc3e7mD8Zwj3vSEy3OJw9n/q
Pg2yjZiiIpzebrvCMX1sAXlxJ0flF9Pus0W6GSbXv2fR69FE9vjy7tk47pk2zadr
mnA7EolHJM2rOBZh2kCtML1HG7v4FClvB1QecMrInhrJa4gpnSPUDj0oBsuu/ikE
cX3YFul5v1ANq8QpRcyGp8PUfKLeJaKhkgm9r3/KZA8tP2j9UZ2h7zLK4MNXfauR
Y8ho8tbcCK5wqLmDzn0YWcnU8IW/zGvvW/v15RUCVOpWj/QWPvJbD5M44dBhznOC
gZoePMXNELHSuoP+3IFPI8IJdBlF85WSYTe6FTJIUA9zjxWe3xn6Uk7M6Wb7s+MS
TPfHpUijEFpOfytHaZ4ZRtcRMyoRsl/JskTNDRNU6TFO1aUtG3Kqx1eZOIFgu3ua
R9HRVl6JJIAqFrffS063Yxu+mF1rlbmp7dqB7Ge9yfhhAq2J1n291q7OiE1QgUKx
P0+4axpd2izeiWM9bVNnZXuevSa3s0pSBYywN3YmZpnEVF0ItoeCG37rWfHjEZu/
mzvAiqYplX8gJWjRdVC5bOjey31oQjTeFhAraiqM3QFNBo/YKjlJDE8wWKVLQzgI
7znaQVXyBF1YC40dJvw/JdoGTronrR41zkTqjzVz+8s3bL52SwcA0rMbubTgjlvA
oxuPxMJvfikuKSYdpLoevrAisgd3dJwAJ6VhZsz4olYYX3Cet2T/2WPuvMbGUm+n
jt3qC1Srp9WEHRhjCmCenaYxdnHn0+ikTPd4jzlOI68YLuCPk8nnh0k/IpC733jv
KrHyDUQkLTj2vd9uuU4X98hb79WB4WbfpT1qBqNJug7Y5ZBB87+c0a5tWD8vQW6e
aDmYC8Fxz53zRWn9cyLHhOskhn/KHoGWwJlX+uV+Qj9i62zQ2DQxivFMFMQruSzr
v1hU5ZmLO8gd6qFA0auBjxzvHiwBAshcK6WRHvRnWAkHntl9OyN3Z9/UYrU0YbmX
sSUw+6Q+ZISU6zvqEeyKt4Yb4M2ETsCfB2EfW0pXZ4PEWpX2tcyXS49GV2n/V0YT
6kKo8uoy5KN6Uf8J9CQPJ8v0C0K/6tVKAvkVHX9GB1tEOSr2pigS2lWpjh9TmwD3
8hYEb5kr7lUMg7BbQRkRoOepGIJmoPmbK5LfA4DOmj9M8XcT3pfVCVoTDVxBciDs
167rmt0V7ltAUTccj+6Qe24aqHS08rRmveGSNIHuVuTzHd+MxHFrTYT+4Hzv/0+J
HmJs9vJEfgi9CUY4g82D3u+mir/oYPBGXMYHlkOTx4BCDtTziGNDgbzqvlJy5pIi
X/a3rMY5nG/EuPgERYu6AbNhYW5/pNCBkSK3md1HuVA=
`protect END_PROTECTED
