`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wrsZQot1GcRyujpMBZUhyOjBBMx1kpq5cbwtWwpO9/o5E07h1+yJ9gFvVz0pO1gT
C58cmKVfIjDsa2CBnPEF9I0nnW3rM1AgViEhDsBbYoVT1nMYBWJNjKKEy8IMkwKD
Airh10Cj77Ta+f2qcfgf9bZuIuuK31E4cG9FYBhn/tjYxOI8Fohx0RAOPqx8w2Ka
EATQt96zwYCq0aRqdx/g3eHkn0MjqV3wgniG31VBr680CVir2SFFJ7eNK2t5xQdD
N/Td6aRxMLbuCLdFnm8jaJgNTQ9Mj3GMJB0GGjGDOluX377eaI/jpPCZ8B3hnB1n
Uaj3yx5bVcPoZf/aHc60Q4N9caMRkDHQtj9pPdAEUo3zH/UtxXojTW9rLS4OkQ7B
KYsfIUgJglFJPUUiuN7HZGIt/kE2cwwKAicXa4HteXrj2TeNxti3p9SJZMiLZFV8
IUL9OgdyiMkJ/a63wd8fyWbBVJQ+11I99KGMEUqQq0EuGOobxE93BqZV7gaymrVU
+oW1Li9DzkLM4cfRS/rN3wU0ziztZSYHagpcz396UUkc7pWJ36AMAtD7Q7SMMcw7
MyCnMY9Kzn8kthi2ksOZ4TQ2fJt1jHlWPxYhxAC+n3cruEmtKmgfqNcCmTSSRRng
IS4jA2aI3OBsy665x3Dj7UgXv7e9uP9iDfPruEODds6RjeFVLe0zBTSMpUC4irty
quPCqhQ2nikda+67edK8dJlAibMKn7O2b5Mw/LtFAW7LvbnvVpPGS2450JvbJwHN
6O2JkSbLJht1wmUMMb84/Zcx+XAwfx/Ie7gR4qajyLYc7FqDuU0WPZqkr+sIc0/0
OX6pts2/c9HpfL+5VVh7xbOEMOlhQ0WEEInpy1wss5IuSMAfayrNq8vLX9dmoYf0
6XkxNZsZUyCyAz0zDEs0Kew//IHzTsVQDStzwG922vMjRwAL/PUr9Zm+UX4ceXQp
+178jIh+a6KQDgRgqI7ZSR3ECU1OdyFCIcb7V1G+UPwj+U8XtbX/EvQrmc/pQj7a
p4ZDQFx+sDkMaqIVAt4TvUPDoKFe8kTaay1shzannG2IVWQprZX7ZcK5veFonHlo
f/tBJXffd3zt0RldKRzq5RDHJ07tuxLY4sO+77BPTwhA/9K6OQmlLNAEZtlGxJHl
5J7jjX3wLiaryfq02mLDwhkUhVp8Ntw/kWbax0kvxCCC9PzwH536AKAS0NfP36p6
otUL5fsgYrIMLtfxvw3rrR8eQCIOp6qnu4RWxVNnohunbPV91E+ZT9vDyR1L/Im1
4oxqiUjlUW9ETxTjg3bux+D53tAf6zloHXhMaCqJE6upYVnwCJwNpO+B/CNM1DAm
2RyRBg6oU6A2e0UtjshGzEJAXkpC5raLJog5haj9VDOyBA1QsqFH+PlpF2WeluLn
guGQTNqnCURQh4q5DPPKRL/kGIppCQ7llhR0nPIKSzVrVgOjYjBKpwZu3t/Kqa6i
w63YZyqB3WQJjCNCrWCXbk5KNmGZm2OHA+8k47x3NmvRieX/qW8PwbIGONzhm0ZP
OSD0jWqFkeVAr6/OMgKq59kcLyd4o/ADkx6quMSqDdDh9a6R7eLctikBTn/9F9kY
DxzxNvseLdU8LcLw/MSwxUoTdZBmx8FpRnzLKQjq2Egig3msoIcmCeDJebORkEgN
nWLo3r3ChQe3gaVsthwmwB9Xey3FOtXVilep1nvTLYu6wfJ10yYCn7wXCxVuGUHN
0sUDrT0YAouKXClZ/4aK7rwSyeq8s2u3p5g0QkDMlPMQLQiAsfUg7kk0UL8lULFe
7SV/y7YZnodFAS2Hue5D8Ll6mrhpSfhUn+3Q6ojmsU/h44flkNzzYDJHUVnGEGpS
yIoi+wyLC/SE8aRWqt1Y7U/0kW3USfnVCEx2tRtvGchabyFfR7oGrSpGm9AYDo0l
45eaKuwL/z4U3RfK8VyIaraUOGJuNJL4H7xR510LNLIQrHytcX/p1hDo0cdQXGst
vc7CaGiZuMwJuAtCQj84ODKoBR8BFuRHaDeiMiBfSpTz7iajTHwlLnhbpKoaOwSL
T2CAf3q3yW0Tq9fc7yntOIa+aGg8I/aDtdzvlN1qnzRq/cnD3VSFMmhw7iiDupxt
AAz8V2RlB0qhzAf2Og5d1+RFYKpIuZ9pkBx7DfbaICmlItoxIZKJRAWTimgJ93hq
GNBhUQUbCmGg/q68g/r688kpOvy94SlI+HxMgJAkL6E4gFmsMTeZPQLi6Bd75Vh4
MFoFg4NqXpl1tVEoOyh90dxTGhkADJsMCqnanQZpOtJqfMQupU26oW9w1m5C5Jd1
iUZrGpKgyZ1ylz+5z+i3miyQfrKHE3AX2XYt0vBLh92SV8+jAoYG0L0BcPf0JIYN
HPI8YwaSPyqH9A10sV17H9Oqun5GEhzWXGWG1vGrNUtfdA0xPIRCiLdUqfZx2Bsl
uLxrn3FksNOOeqZ17Z3LbdvZaMATGcyMgRuG4NrFND7MdYLomoltIEpCbbazVV8A
1b82mgCndUtH8xz6myEuQBmTJtIPlCYe7rX32H/Nu+aRjRzBuyAv8FZyMQb4WTTy
mMkNob6wnkJ7UcaGaa6IRS/G3ey5d1TRa/1LdhCmUmfYn1cl6XVCWJ+3hmEERHNM
ykKB/WMrT5+YvFXzD72FeQnqySMIYaDUOIrS8LHKQx4EIMY7iE9fBHP25SRRi0/J
scPzP8gLfdXWA9jfZnEK8km16CKHSQcEB5buzGAU7W4R2OAsadRioZO0W+aNS6Fb
0ta5VzeeCe6leONM3kJer5q7sj1X+6dMNonOPVydAhNiv1eHHFfRRbeJs2YWjENC
PzB50FDA6auRzBoCCUtckkyd4psOw6gMQzgj5svsSAEa/fuZEKKT+98YGbjoncNU
XnKvK0VBEMQ796xbAGXDCoSf9n2/OjpxgiiSWNm59W6fcor1LcvoyfkzBKLF1Umc
AxMFEYOuLwVjfO+oQpEXkDzwYmkNeY/IUqiE0XGKdGlTY9lDt0VNkIuQoHZCc4xP
0avvpNnLoTzYYzkS2PkrF9D49wINL0zTyvvm9XOTs/25A7k4fBwD0OvPFFU7VrQB
WobIaf27qTfXWbFzwanf0m44UuSUQaG4/U0IbmDMS5GyGD2kglrynR8l2YhNBF/5
4i/1Pp3W6uBL4b3h+o6/1I9tZI3QfeVnF1OmckoAvsb7Gx6S939PbltLgRRGOQiI
40IwKYPivZAuncni9WXh6sqSneA6/BE7n7lh+oxvF1tD6Gi+6Y922JEVjOHWSBSA
74iwMb/yIVAMRbh3M2GWfNWixQDJKvXXAFopGyegBqcdks9rS7LQ2sXBN4OgQWKU
VK7yc3aSzvL42ZXf3QTg2mqC889mDtpMUTCrG01UzOr/iBetYLb1zCkUHwbl63sI
qNHXNr45SpmHVRtsn89i61uZfJfWZoZXkgFVIhxJJfXsOHzO8mL4w4Nv+MDkOJUc
02yc9YR4Bz1faUc7oFmZ8aIG7cWG6gbhNjUQUw6wYO0ZtFyOGBk9sHbbxjci4/oy
0FHe6zVW3noFZKUpNoYNNwo6GGr/SMtEZMKd8w0Y4dDiKdsa6bu94b1uFD9r9toO
+n2Mj42HyUgU0qWWT9BoJN1hqgT0iFj4ns3QDcojko+cPwTLQ2w1oXNKjjzw4y2I
5AFL0vE+vRZkq/byzSJAOI/3fvic0OpjJ1VZm5L8TobnqxXjbYPGIRUU542DezDE
fvqccDS/5qxr1A7yI1TJf2U3z5VDVL3SZqHsC3cYymzBAURKt+czdegHHnHDaonJ
qP1hv3jqwb4+GKHpLtlsCg==
`protect END_PROTECTED
