`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r6NAoN/xJtVzRQcoYNv5QLI+CZRV6LxS7QGmU2DLeQmKRKNc25hR7jcNSzjgKBWn
Ed3onfOyHF34Ru6h/pSdoZjx8dL8ql/gJgYSt7xHYnnpFWYdnI5J7Uy/M+J2Hp0+
rx2ojP0FDrneW4h6z2I/+79QvwoHX3YtA+fMVyFJz5mFwvFZfI6m88ebqCA+D87g
iOGMICp+brR9WzQ79l13uIXfj1jZkEZY3lFHwDRPIAN/UrJ8/jvLam36tAXGTtHR
f1yTSa6hGxVUUhC90OMKyyXWv6+7o5F8EYeGxXNJtQEJeQhFjKrwJtKFS+OAwBVk
KxNJfBHzkCBODn2ZBcNqrAwKYEtvJKBjk5+cmz662km7I1Ffgm95lqGuTtgDVFH7
vp3DWDXHY0lUHZQ6XGGRq3wHIuLpKWR+g0bIQX44534asfphNehpf6IVyGjm7GDY
dJXCOiEW+G3oXHmg8XbqCPREbh4eFflziBvXLCgvP4RdErhJbqm9crgJFPlkg9hV
l/RTdxdxV5bItLQmVsIeu/z1TAovtz2dAy29ank1R64qBpFjHxiMJmHaUbUhWr82
xGEmbMVTE0D9Bw58Fa4ss/fKY6E+d6rRMqrIth1JnogKbLEoxBp5jCb6ujJOIBo1
vgH7VhjbE/2iHCRp92O32wZxsoAI9iDnTFHWsQJf4ya4cg7lEZBUq0H2mU1GAa1J
RThSKlcSjlI0J7XgJraBBwHLIGYIAlK80F2PmyVVVxnY4O/Tj+spO5zHzXW2ztyk
yNjj5UP2BIPFHDNSafpvDsRg831vtyLqqTcA9vGaH6T/qRyg209wACDcSp1m6ELn
LlEZk/lQyBnMjwFp4nWEPr6NLsGoCFl0Efa4zb/EorRduCL1u2IZeYG1GdMD1yDd
Ceck2GfhjwBICvMzTIQQPQWsWUxFwEnIrH8lnl2/lMg1m4HubKKW+dT+4EJSXbBj
HfB0clEFZF2vgnQULp1Hqmu4SYPwBhvocEtK/gAsOjto9lHIq25WbUtqeiDXRyFZ
7H+1gMBf2PIBkJzVW3DPUWF/Z47CgDAPWDvdaGaaXd8=
`protect END_PROTECTED
