`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wpmZEPC0GNYiA7E0mzKNNo9XY/ZjSgR9OvTuDHcrSSQAlvaSi7wIUQ0xD0c12TgL
hGnPpQp5OIeyGSjd1A44Ey2wxgGTDHce9dqeejkBAt+CZDFEjPd1188bVSo9IVJa
6UbkTYkxU7YakwiSrKzteLBe0JwQTowCnmV6Z3mIBHnWkYgxyWZRv/SRSA2IpCxi
WnrAaiwwHPPJXHHb9lOXcneimfgt9k3UgqhKt0O3rYSFbZEi2xrhs0X4A9Hregqv
jdnWqzGKL7b8QgL5OGyJw836VQrmEa2fQACPTuTDRmB2991X2cGpCF980r8bApMH
NySZiMjJCSw2aOW0b2QqOFHqqkafy0Hzu5UpknN1S7LZb9qBtMbBgTxgGtl4FEDF
rSG9C99IcXcheJayaS2+Vaox5AhUnoce79A25QImhFgXiIzsmn09mB/oR+cK/mB6
OZU4Ty2xRHPQxma7eSRCJdCXq25A/y95ITjnE5AeTH85WrK29J841+0APHQINbN2
deKoEH0F2p5K+TMTcXDqA/wllhBql4b32GGp5hgf+DTNInOKPXN5c+Ijc8+VA5dT
E6JktNmtVjRxMlPUIc3GN0YYW827xrOBGOG/JtEgyp5xkmdk+Rh+/vKT89+kpBoE
cuM56ExDhzf/ACL/SzYOhfLpyjwuNnHL3xkAOpYa0BY=
`protect END_PROTECTED
