`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nsRxYRuLHCD7uaGyKPDDnyjRTm6/3jc9oxd9U5Mo7MDYPEq4A4zq/eSFe3RUGXAN
QEYUrUh2VrVSH8wItZAU+ggKEVwQGjDn8KOb/H1xGfG3b97WdSlLY1ps1jb8+Us/
6jPL4a/Zw5NsKsbkUfXPwSKc7+kJZP3VCze1o4l6/bbq4zjJUs7VqPRGO2xpehDU
ZXF9cREtuy9bIRWqDEMJALqONNKrG0z8EkeBc8HnYZOV8jynXou7syw3g6XFgekx
bUaWfKqvjI0YTeUoClmpeyCkAf2qUGD05g6KDjmYJeWZr9jOM+02NSJgIPodbfcE
m1lhntHtpn53oo0IdofNkGbiApAWMWoXUWE7yzPhSx/JJZoUlR77NH487pwn11OU
ACjPH9Hlg9bzZdhBywe9zQnPJeSTjIku1H1uo4AtN4Ji3S2JqKEV14Y4m0AZyYMc
T1jngnuftcjy/kGyRjVYYz54NW1Xn9OvEXZvxjlU/pJ43NNgd57S4qgHB3hnECXW
Q9/p9s1ej75rSGz47DevZCzbhqPqXO+YX0MSpFiIFn1gAJ/XBV/gxp5r5AtV71Nf
GjZDMaFM1tt2KUC1GSOseEcFWdzH0P7avj2vi7oWVxOmfb0MOk8KELK9TkRIueUE
LuLJlCpc329Qo6duaB008KaVjHtMF7mervrUlrveeCQwzg6DjbMF90xih8u9+x+Q
AiQ+bspXKawAj9C8hfSbVPQ57ffN3lbeLuhUheGd93MiO4xIQx2oB3DNMFZ42l6f
ZaujN7+8r8hm3VGdZx8CSs4BS84XbawmqMvHEkSNhC4xY8aBUUodIVbY2mnh6iH8
3rqj6CUXMcb5yZ1SoEVG7qMMRwimYAuLQOQkRuCIB4r107QxsVct2NEQd9jgv8XL
g56wdR3S2zI348YHJD9U6ReTYzfwy7BLTJVdhgrKPC4ZZX8AGtM/UBsMRj5auCMw
4/u65nXrwCu+bAjt08RrJ1aE67OrMVzWr0kDXmm6yLZhiyUHTdwFL0B9t36mLRb/
6M0ud9u+X9t1U0yN2QbvF2bJbyKvC09VRpPkNruMJ9oeh4weMxzozHtl20QCOdIw
3wMjqU13TmOC6xLmj68CpttSDvveSGn8w/xyHkOPqB4S15qVeIfTFjzUc5jVURIv
wb/AaXgKtrkeNnexXXFmZey40db6IoGkKiurD1UbCQcrpIqKQL9XnCfg/gdrxbbf
eryv4/OVzb4vvGGB+S0mULV0xP2CKBOOWtklp0DPojbJqI+RDCstcEhq06Urc+eH
2xMM9ZKYyNteFbGCHttmp63Be7aDu8L94cnAPan3hlLZ7vVZPA8kMZAR0AAjfwt1
lYGxu5OcWvMxP2Q3lZ9GEmIfQgdyLlziccO068TKMrSmCFULQHSNYvtq9pX952+2
pOOLE06t/v3CaXpj48bteIaU+Kv7eEVetnsmLCmgrWhhqosIHu3PKKeNLUbmVHuC
PU6rRmzzSb9l2xiKlly1PdYaq5E8MrM1gPBMZilMG1qdB4kjN6oVtVq8QZWgWwvA
ktyyOuGqHquDbgX3NpcgmYJKe7c/AvF700NpXYVw6kbv6BSbNXzbW5cwiX8Tf+8Z
Jn2Jlio/KgdxHffBBBSD1txIL7DSQhb15gqE41mUCysxnYm+w4HD2DIVZiXzmUsJ
45GbhhzXVG4gujOLtN4GGkT07McUBNiCCQGp5202rNleBjYJ3Q5Y8QABjcYlGSDz
cFbL5kVGGPD0t0KOk7/DRj4YwKLq6dfrnmjU1A4GsHbfYYSJ2yFRLmTgaoNdKIwR
mCzJ2FzMNJJcJl0mPloKG93w0HtTkU9ZKlhrOGnkj6DDX1y26S/DU5wq255DpkrY
PdEg2sehBliIx7KaR9RfQLrKJgOL+xrYYhbJsIwatc1Duu2AKrU37r34tqccL+fA
ftbRo4KeXnOx6Beefi7hNdR+Q8YwcVL4S6QSBB2eka6ZcGKRNVFFEj3bu04cobhS
nhH3xxNJQowN7zBE5JA80w==
`protect END_PROTECTED
