`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gUReQzM1OZsTClSs7/rt1NrcuijFZ0cyRSfYrh8X+bCUSEFtcv5Kn/h0SZvf0XWW
d70bF1teW2nNFT7KmIA7Hq22sVhtBzB4Wus0KdceWFIgGK88ZvVIfW0UhRX2QCON
gBTh2KmP7X7+CrlmTbSLl3x19D2EarCYnfE/LKGBzAOwathXF7x6gpX1l7+TmLnk
MfYl36aPPCnTNtCsMDN2maYvqEangr9JHBghDFr2YpUdpeq9vJDJCGnv1weHIx9j
6vOPCqb3iVSLcfHgMvFUTZECTlqHjFc1LKG0ZhsJb6sXA0kK+K2KD0ExRQSS4/lM
`protect END_PROTECTED
