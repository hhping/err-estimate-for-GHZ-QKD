`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8G1HeO1a1EDdHnOrcBbf18zyEIX9Jt5xRfZeSRaLbnl6A5s31BP+pnz2HvRcaJKC
HfO3OiisXIPfA7JKWQOVv1KWBswSmz9TzagaseO10Nrpo47PCMcC3Zxw3yMFswKY
HwLnRkE0oWsZnuDGfxLlhV6unvE5CRFf88kKBjn4t0H1hgMTm5yhEiyiF66YPjqM
9iLDlQ0C47759IMub1mdMetVEsuHgsSCipghnpU+TnVIWmb6JVaMnFwF37Iihdol
c6PTuqtbN5xb1JIkrKzQUaNuSv88EG5TWmC6Ygu53ucYXSX0uoPe2eiXn/YwDgc3
rsvGprEyYpk/yOO90vKdFfmvNK8+sSlX9WKhBj4qDuG4jfeqrymwzhqbX3HnhW2L
wEpC7m0MHSe86GyInNqrCfNVoWqe9WnL4yWTeil0ERY+F3qaD+40hG1Y6HeYkcDO
fbQlHykZ3QqgbfdZJbB+8/AhumjbOD8aoC/34Dj1eulKvzXlt6NWgJve32dXB4m9
AtfVsdh0BG5AbGEWQOG9oH07cIXJMwkfOAok3H1INt6uIRruPvMN0VdlUYLhoGQf
Hl4Pv0T7xk5sMemt4jiN8RbXOVYLSlBMOb+1kNCzZ7Rx4ceu3oItA6woZjsSfDmX
jcja4wL0AzSLhl6xSc5PfGIcSwzVIqnKreVs+78gb7kHHakG7NmN3fFFkbVOaGhT
bHMOZ9nMcu2tyO47O1ypkpQweDbBfj15qIbd1P55uS3iLv7A4RhC+Vt2JrVHCP/J
xZF2PAktY7MPdfU9eFMFx/uSUWYPwtFGi1p1dHY/r66cLmD44oHwWHMX+bAXC7l/
UKF6Kj0Uz7UHilvu7Tponw==
`protect END_PROTECTED
