`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BGZn2a8tbNa19LPzHdq8ssNOF2rWuiEXNgruMd8ArAXUOfE25wZBefjvoNyyjOKi
ht5gwOXxo7ETrrO4ilhuRkP7NJWYXpQJfFItope+KDYEfACs8KcqwXwfSydfwZtG
/77f8EnYUM7HeoJHQrgI7Y8EadAQ/XtSwFVKWCGwnk9XdQN62wjd76MQYF6i9SlM
83+4o5YIg61uq5akLEG9ws4OJ4hdPJZh9vtmqReN4W76U0YhY1i7PfnT59bcL6m2
ytzLJ/Fbc8HsrjCydkuT8tQYsTaCYGeFaoON12IuWxZSPaE7pDeCkoY8Dtkdu1+d
gRq8iaGZ1Sbiibg0RJ8fpw==
`protect END_PROTECTED
