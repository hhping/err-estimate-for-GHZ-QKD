`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TYnDL04ozfF6qHS8oF4GKAGOnGcWkTGAnC/BK6MHdf3J39z4IZ/W86mdj00bylF8
OEZVrbOVjnHaizfZ+DJT9rzKrAw8XOwkGJ4xwISTbAnBpvrM8UfJ/Gi/dd6alr98
xkcDYWSgpbI7FbCJPfkEodxPWf4KkipZ+rsaIsyQsphj0dpLkiKBcZZTPZ3xI7bB
E9WiLWd2RTunjAYKISBjahon0MUNRRhTa6DuIH8NQa4dHmLTz/sdPN6Gn0gw7o4A
zay40YoZdM/oM1uoV8Z0l4H6M1jICu2qF9R3QONtDFMBtbdOBzC0ZjH+fS4PZwdO
e9SEjYq6IU2cCS9mkqDqFB38a2M49bMWPVf+YjAWScdwJns5Zp6mTo8/CpKd6MmC
Mja8sY37IYo+3LCpXO1XBIdoAqUK8Jxsaj2t118xoPDlfeF+dxfjX+pBBA6vnFRH
AZAKbGi4HRboBiUsMNfjheEdEVLpezBhtxiwi7L8BZpVpQtkVCAZhUWaZOHqiJOS
1zT9iJaeNbg2zIG0hvIwHA==
`protect END_PROTECTED
