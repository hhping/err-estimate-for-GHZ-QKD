`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IRVsw1W+oZKcXa99Qt4DJMKRW55yYl2s8bUceH7tePIFsJOz9+usZTwnv6e1kE/U
tClvPgKy5LB/KiiTorQ/JR9egxDHQgVEtjzS0FCvomA3ZnAxvwrQ1yggjPr1W7vE
2WHxF2EYsdlLZB++IoEu43sNNNwT1qrJ/+LD7HoNPPxy8iTtPUn2z6ciPFGLdlib
GqFMgTkewC414gZTIYthmjKsF+WFEtrqq8bR/4NC1JY2qZvmSi6Vb8m7VFvIqIUf
41sarmc9wxn4n4DjvdoCpDt6Qm6LHU05yGCGDnxWYLvVMbbmS2XfDw9bYJ4qVQM1
N54EISxpRjPv7v5Kx3x/7l5yxQyzcyBGwJ1i4oXZyznmkaiDIH7+eSZYCxsP7qZx
ryRfW39oEAuOnvgGsT0hEH+H7C7eQDer9addEKj10hp7cY+KggDynkIGB+2rNNBc
NZ5csK8XoLWthCzzKkuXmRbbD08gGwhV1pqbCNa1LV4ulZXo7VwoqkCDBbIOE58n
daDaVBcSXYJDaR5zWc6NFGMe59RnZN+tpFm83LhYi3S/1QYGJ4w7JLanttKsjlzu
RHb9zEl2YMORV9TDEtDbBzcE3SNnQd4sESQV71grnwZcBjfubw4z7Qy1BC5j83ld
Xn09Q7+X2hc4hihi35CYL378Vb0gqBtwMAMOQppZy2ePrsMWPVX0lt+8sF3dJFnR
VSQZf049t6KHpvluk1gCvTMC2lJbWNVGKYlsF82FPYBqNeKvoN5STKN8BHwTRizh
rPGqqZ71o0zLB+5/HkYo9w==
`protect END_PROTECTED
