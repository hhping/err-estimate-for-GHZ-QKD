`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bi/NsD6ohYSq2Sf3U/wW6iYzpV4R7j8hwZNDA54EXStD8VTKWTkZtf6CTn4vl/h3
0gEurCjAWxMCd3YwU6GDNI/QaMoJaTMWLedTTWdWgV2cR4yXkjtp2BN7hVPRAB6f
aSTDaRZLYDoySrNgCEm5rn2Mwr/NTX3QjVIK64/29IDlbYbgLYEtQJo33N0Vfj1k
rrl4jUvzf33hAgs2pw99aP9dppKVHp7BwXl1qaVLj4i/TIHcCEGIXe/LnrTPSSUc
JgWDeia8Sss411D664OVpNF5LXq6Sm7LFXuervDqAAgmZLMNCeT/+qVJu/S/9PQq
1UFt1x9tNRjYwjzMNabPmf1DDg9ly2LPPsvOdqkje43yw4Bc49ADOfGYL6tXS9up
K3t1ZilFvaECgnfdQt8zDa455Tg6iDMbxGpVAal0dRJOoaGPgLNvsxuzfGF4kwTF
Xlpll3KDP/T5PnOIJ9rUGHUox1CVEhBIIH/XEkL7ECrlMFMh6Z6nlne6Oqw+c5Fo
8ONlqHn9G7AIi6Gi5koJ0QTgbrDZv4y5k+rN+nIC3r615q0ow/dev97o7cVe7sr2
3O4HcXxeMBoUbeh3qVeKahrUKj0JXI56pGOqXZ6Sy8heWg+FEKYY/gh7dqutaUKD
ssYF15PtmdY317WxRahSHJkE+1m2yXRH6lyGQxy2S+p5v0L0uSSEc/OIJE5kzwIT
mDgb2H4ghPNP8xF76jlRwHS4DLkpv7/2yocG7yJDeCyAEj+B8zYBhaNLBU1AvDaW
`protect END_PROTECTED
