`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l6api38BxEwAWqVBMoseRU9MKpSDA9QZCQUCZljOg2RGw3QgBo7wDwVbdA8cyIlB
KEGBMpnzPnug6dCA7ayfnkzyp2qRoRj8ToNLGuH8ouAJnrU9KLCux+z56cDEidy0
V9koQVODFb6cKZHkLmBJO82hwZNvVBv0q9ki7RFqWMBCCOt/jCy0WO0fcOlTQzM9
u6KJcUJeLwlO4PMcKQsKH8K1fqbEQ8Khb9xfVF5JBrT6IIVSnxSpIMT9c1EdiOox
NAtdDvNwwXsoZKKL2yW+rCD02OqE3ucuTBz+uXMCdqMXW1bM7psmb3IeaphB78AQ
6N0+r0P/wSamyvGacp1rHa1oRZtgi5h94E4hqukkwVmWQCbaxG5GVLZlt9+s3Txy
QcecFkwqxqc5R3uXk8hFn0ISE9zMlbSL7TCntcABZhOfkKpgfADOW46oY4gqBkCu
0YggzBfmwtbPYOxlvQlfrQ/7AxkbFTlIB+acgNsDKq/VQtvgWolRaJgEnGLJFeip
ojv54SzEARk4cV0snHqOzaWD7Z1zx0/KrmVMV/VYldwj+6D5pvvphJ5Zq5I7RTbV
yeQYBBRTwL6/FFM7XFqii3yJ+9A+1XDDngoFGlWPx6zaqX/UF0csCBlSwadC8zh/
N+f0r16/rtQSwB+jBGqyZy/Dr+ZKsgmrvLXIh0+YkZc3oHXomzu4or+PU4znSDQc
qTDpUQxkw5W0d1UwQpfgOUiRm4ZfVyhddFXjHSQqlMTCLXBuf3phbqxD2BWFcQ9/
`protect END_PROTECTED
