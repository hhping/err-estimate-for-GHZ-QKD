`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6x7qET8P9pWGvHUlivgnXVVLGEWb+29SDNWT4aX7+utvhgvVs9OQOCvbT3HalxBT
dEdmumLX1hvH7aC2EewCFNC6kA2nTTh52JOb03J4k+dPz1Yuvut9AOB5IVL/zVgq
dSKMYo5NhYZ9ei/aedkHLXJfbgaQVxXq9g4Omd0I/gnzdbDPoJ9wwDtxut7s+bxH
OpeW/x7wipBaredks3HYZqt8z7weUvyL+Cb/aeaHHMgNioOmcTPngXNzAfiN+Rmu
i7rP7U9QEahtuXWPmrrfCNW8YMmxW9Dic9xC4GfF26I2E9zKC5QDaVAk1CAyLGkM
GrORgICnpLslXRO1idbGmrLPkrk6/yN9GrEM6VNXAA+yGVRDaEUc8lnbGyNWi90k
oSJtH7bDeiQu3Y1rLuamb5URt+EZzTSITuC00nuecg+7cHuHD7w5ng9OoA/QZiTl
RuWOqk3mfqfRpjMiuGdBuDmlMdR2m4zKHK0OOa04ZdzgOFGl/vrzqJm9YqOoiAhO
/jI/n5pHWhE8wd023jtokHLVaRGBxJRR2gTcDYArTTck6BTbIJjh5UX3noPeNfQ9
FWT+MQnvObNSmE9p8W67QeiRO4qS5AQPbAJPn02NOfL50a8UtieA27VQGYLPGSag
53Pk09TJO9+8p8gZGtLQS7EiLOn4Ci8+1kht7GeyanLabc1aypKUGI7bchTx1+Xu
poX6Chh8yN7aFIExejLw6Qn3ah3bV6DzMjpOe74sCNdsIvt0Q0oz76cMhpk47Ar1
/rcg5vOjjNBTRc1IGQ3rKEQTcn0wo5jzaYn+1sm+KLg=
`protect END_PROTECTED
