`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PR0cknTk/qbzLMUm83DW4fK9fxDMAbPKwwoguZjEoqRIQQDdor0CuOAdF7F1Tvtl
OfbqTnuLj7Qzg1IDPLpwB0qFvB1N4ijh5Z3HerEVMR5EXojuxy69FFib+m7U8Rkm
uSN4bEgnqa2ZER4tuOOCo3NXizZkkibUWqFNz4kT6o5INIodfQqO7YHtwSTQte/+
zzcugActuEZPZ1GHy9ONRs8zzINuo7ou7gOYxdNwoGQnqDWl/2sqd2D19gSmfoyA
qFuMpK+DJdD1u5cE8zhNdhL5XHPu2QB4noo+uzIl2U24aZzst7ST4LHrBdB2BnRP
nf8jDnLdEUez8UtaJhfqsNYCftrnFufS6oJ+KagEA5HYCMKJ7dYXjoyX9J1GS+0t
JJPpjIxm4RMb7jN/Z8rBX9oQOqhL1YWmXYlQsjXYNTvrBIMyp1ngFGOOI3JlMbMI
eYa46Czuu3/aDk66ak6+5cCm3/+HsRbC6k2Y5VVqrc0y23SNDnnlgdv9AHfqdzSF
riULpYI/VqQgsO9pYK7q7UfOTxNL9e/zQcj6kt3Nh3aVsAtouzbXevkikjf8D/r/
MbF7w44fny1K43Fk6qrL9jfRh5KEuuoihY7gYbIPb7+HLt3EQ5PZT3zQvrTLrsHk
6o2RdoM+9+Y6qo1UCHXAcRxNVIW9GwpoIuQqObYPcoDXnR9Apx2LMXXsM4lnkGOT
GTy2J9PL2REz9Q0WsLbXCPaUtqF2d3v9YkhKijw5/2HKY3VoRVYMuIn8Rns0pVdm
ncthDrPeMuzLXfEclEH02EMN4k3dBoeJwdQYQuxebmfrVAUuGmTa7Tkc7sx2BxcT
qpAB0CdF2hoiVuw6M04pHmzHHBHRlwJ2rl5FhUQp6Uf2CbdUEyhGBUxUlVcRbkM9
qlAfu704J0WSgDBKW0OPcrxj8o+8PKnSZq0E4+W53p7SABJ2M3+UdT5jA1mL1v2M
OoTqMknWqyZUsaBIOskHRkcSv4d2bR1+fk/EET6GfNydisN0vJCuid72So8qbJRI
y+UF6ncgNsrLCzdicQsYWPKWWzxdNBekENeywKSAVacZcIeyWhF+DvoMmWCpG64S
eTsOl2u98jhSfWL9OwsS7xFvPkF7dd4IRmbfwFSBez1GM8d2SnFt+kkwT1h9HKPg
yzxMdDhlcTsLNwTDo/bjY19S5xvNDWXjYTqNj9IYSSAriZ0R1rz71JmXHfi5Zh+p
ycLrpiy6N+pH330YjC3jsAEg16Wwrg88Chl/eZjMG/PIeLN6HWMjGC/d41zTBcdW
TMXVJiV0KR2zP46t4h7FLg/1+90GpJWGWouVdGmw9Hc=
`protect END_PROTECTED
