`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N61I9sjwqaWsc+opWjHSC2gLL6bEbanK/JhewiEMIsyG6wpq0UUAjU3XsaiIH73H
zNkT0PXh2n0zYCkHj3Okv9da9oX4Q51o3xuhMujOlNxb9XK1rEQ/VmxWJmZfp/1k
8+Dy1A7ArTTUVVnur1rxJBk9R8my5FhUdk6yhJhpXPIe4UoPwffM+Ml/VgeuuWbT
hDo0nwguYCF8IkD5KchQ7KgBJ3yKTocP1A9CTeQX+v3hSRFK4+QM1MUZ6aeQ/kte
IO8BOSSxhT7pnrPW6LMJkYVn13CREMRd2iLFoahXzbJgXF/7h/VRf49QtBEvDHjo
Qb53HsFdgzSi65nLBFWub8S2K3bGdbNSqkS8Sgp2udqqXjSRVlIviKF5soQtHuyX
BuBGbygUp2OJ5Mpi7oB+pl+JH859QZwzPhNvdu+fEADxmOb1w10NWgE0KSQ54/Ga
tp1i+KFuzOx8yvTAJccJxJoAIKZ7OfK4OvNy0/Ov0FzM72EhS+PyvfCdJfhJkXiU
VAgcysO8oSoioubcndJ/1Q==
`protect END_PROTECTED
