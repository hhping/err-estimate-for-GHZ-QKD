`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ER0jBb4bfCof0+NE/OnzBQZw4TTzgMdeoJLu1iXcqhR7zp/3WhPMV9Ap8GOuzQ1n
fgT+xtUY8xlg1V8kOrb6PP6NIVb+arPm6HpKgIC727wApub+h8N8zckjVmeBGOTq
DHKT6hzex8D9GHy0bC8+EsrTcerKpQRJVaVVPb0E9xh9T47X4y/AtCIgL5XLoEsP
KVNjOvfmwDn/6RjXlv63s/7ZRzRkDKtWV1jHrtpgCYlmYKTj0wIwMu+hangz9bo7
ta+qVLQkQrJP5nmtanW88M1l+C2JeI/zWeprwc0gZI0vPGdShpfp2l8H1ch+DmAB
FDvANyuvzqEoaTTQ5XLZdgrRfLF2IcX6EtN5wkD3TElWYrxONM5syr971fwoTeDY
JcLm0mxzyB/rHvgFvHTMIwa8dPuVfQLUGC6GwSNxzpm6lfk7dV03B3NJaemGY0T/
Yp8P6twoGFUqkh+PGKPi2mnyrRM0j1qJL82rU5vFowgzVnRC7+dBqfL5pYQvacA0
Ls+CtILJEDBWIDffVt0aM2dYBPOYP7tPo+tPlJq5lyQVJzBKRsMo8irza1ipfZ+P
ipxKLchXeYns6Wdr0oQmFg==
`protect END_PROTECTED
