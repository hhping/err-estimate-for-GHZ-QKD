`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+Df0Hqibd/RqZouQJfwPyl2hw/JtP02qbje46uGoyogCB7Bwo+efePw7FTpJTLNh
hEGEjDUQ1nMdmCRjCHGi0c6Zuiu999lBbuK4ovTMECPSsRs1K2IkPI3///2sZp9y
G5P04/GYATs+fEtr7AkBKwOLj5yHJqqYzAui/pBO51cBHA7F6eBWLSlovhCGAJkK
oE8E6lnaPWcq0LfEuZvFYax4ypWjgRVoiwP/gPjDpz4q/ZNA38j3mL6B26Gd/uVM
NrnVGaaesIfqg9RJlh6sTB70OsQCS/K6TapQnjHK1Y33QPhCx5fW1gq5WjALKznJ
vXiHbzRWx0F6MQkVFJSG3mNkiibdVb4crIJ7degdAHxn+4B+1//ekeFxmFuBDFR3
1WYqIgtep5+tCcBssNnDvtRWM9EhCDN1RArtkKSW411gYNmG68IhR3sVwv4q0lpz
NscRMrkpnscXaFxzajpBqqM2obJ9N54X6HOvh+cOOsx6snqC3VGRfrXxl6ymZmcU
599s19S8JpzPUwP0oqMXtpo5Z/qXqqKN8unliO5JT6T/Lskn7KYNkhZknEMiwdXq
mSofzKB66sid05rhcXFlM8/TfC4mUaBEK2vZddwVVnvEknLklm5fYNu5jqdBPgrz
DZajZVL11LB29jUjLVVb76pmsiAhZ1+B2+7daO1wIskaThqW9MVrXPoP1kBH+ZW/
TWl7anJqYnLG3bsHKaft/z3G7XC1dE9znCHKliRe7d/W7F9EVJIeHdoq2OsqnAJj
opE8MlieD21CuAjrp5aN9MXyMOqSEhD63X9PUQ6Yoq+ptsnqX+qGlVmAxloMPfJd
yNeYlb659N4LjahtXJ+YjyCP4PwZy+VuYPNt/sx1TfojwPbYWbnyBVBO7Fh5bwHo
KHGARnV68U324Bw9yUqolOuo3suIrMebPYDANCnEp+XIUDQeOh2nBlE+y/whVDu7
FIVI9tlgISPkIu8sS+fzHKpuOTaTBp049GSxBj6JGO6GArUEC4Lq383sLmGZPpN9
ymQITSWFS9T1wbJ3EBqCro8SAUSkUt7+5Ez/L2DvfKfPQpjsGlhoI4e8mekDesEp
UVr7GxDhxmUWubuM+S8rPo4J1mpYY2Tgjfe0qtaZ+KK6J4CashaULqn4Jbyi7oep
ApdF6sMRDaNFRl+HQf/Q8CREyBni79MBJ/gFMdl6fDUKtr4VF2XU+yC+8TarnKeg
yk4TvyOI8Nedgc9FBg6MIzyZjzZSDcpcedghvv54x5l9mrSOHMLXtAveqql6gpI4
FUveD+MJhxykMinzzxUv1qeUMKSRjaTRJ0sOzq92a99OTO6dCnBt0rX2/clvNdgV
D7kJrV7emxUdqldEDQQxgIvbtP3eyzmkVzfII2OHUzbzKY2GbCaF2BvhGV9aeSy9
xoJ8cnLxFtJooSQYoWKTEbi/8awTUhDqVwmxPkzmnL9aE7L1JsBeqXz1hc0p5qir
x9RHTrpjJXupv9o+zR51hjjw+Hd+QKGBee8G0K1AdROYYke0BQcaFQU66gSD48ja
FyFq5vevGXaB19e/3e/6aAxQrpkgjmaA/MqQ/hEAnf4upG18RaATjCRNB6Ng1prm
U7u9ovqwI00IEQ+7GUwPvTLjr4Q35IYkMxYN5/iwCj5Gusi89w4f3bvX5qyz4dd+
8lHldXxg8nq0ZUa/Op4asataVJbpSUOL2TRCpqxPF5kiQ74vy5/hLsKLQbJdLkaY
gv0Qqq3EdoaAkQpWEDcZfFGqdw4co3y68Sk+nY2KMdVVrvIr0k5xGWVe5FDF5Owe
VtGv7SWiJc8v/nqYQa17tmGMYbyHRQ9902lxfrQBuEBAaZjwq6ssPX1PPwq3USgA
uvJXMNSPptT4C8LsXJgZWd8goE8/1Th0ykn9Lunb14qZ0r3GzFcHBNHr5rJ8JOKO
yfe/JGuYGl2wrkFOxyOJ/Lklv05OD+eVxer4t1INCuBkolil9kJASKvWKGpYwCS6
HCQzydf2B8pNZZ//1bXJ/A==
`protect END_PROTECTED
