`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8pcaTSZ/5nF6KgWwE9YCPHBbeXaw/sikrX3kQwyMZZuxtBAx7br/6HWNGYpqopui
4cE+38H2+dkOHedwzlJccyYowA/ANZ7sm0RPo/DCcTUvSXPfq8QSgc6LfuIBhBCf
Mu4ItVUwaQup8CREkCOsSnZuZPcvprw4GMfUG2iq0SGZp78hLsJCPK79yVHP3ZK2
2jI7quWLjwOs8xAkY+hnptNQuGgeHxoq4zmF+WcQDjK5t6LCMbaJ7cUGLkBuWW4r
FyEgK7J4rpBs13A2jDzUQGNf6YaTjMhcoVpZlNcRocd48+YwMdYG8X04CU9leavJ
1xjmhphxj48dx0WbPKjjur/ZfONUz6WsFLQfSEo3nv81jA7stNZzUwPKnb7xCOC9
4pPrkIPutk1lDXU/h3X8w7P/wS/4fCQjhwq99V0Jvfa61wktH7H0+KBhpqOabhJj
71wgfgCsm6BChmUzL+fImdo9tu1KI0mWqMO8TCUrMwPX/RSFY5CYUiMedG2/2KLH
WZZcr6NU+ppmjPJ9FIweKUR5brDzQukB6DIvCd5HKZbRIbUI10gJcl1jiZJbJt+O
RiPLFQsEde4CeifM2Io3oUXsZ2nsiy8DwERxCMGgol4lmqWFqf5C5yKnxIu/6llU
IazDFgFb/HlqQHn8pqMLZ6KHNlDpzMt9bDhuszcLVIBsqbLv7l/wX9JO15Aoy1bm
bcGO2SZj2yyvJS+NGG9ipXkMpY3Fo6PncduRWgn4zgsJfXsX4H22jgNSuLmQHZq+
PwJh+qt/oFDDlcCy5uU3tMw4HBkeQmxvFgs8cs5Y5qth8hJgzVQZNSuniGmtmxkX
Xujb1+bWLsQ8N27yDr6sDul5wF5CdXSZlalcXmbnPeDv0L/PGGuULRGuTjp6SOtX
PjxCkSZGaMWqWKMNvjINFPR1nvuZnzgKU5ec3HRGyrC60ZrjL4VkcUO+LUEtkHsN
JTSW2xRp9v71mBCX2rVXgwGa2K+iJrxA935vl9awp8OLNz12I6oaSrnF3f2KP0M+
+BMaojI3ZgiGl463gWu24aPhix0ZDMbAIpJXcNBUAOLSGl8BjsBja3oAC1mXVheI
mrVXcaNWcHSTN897NN4CKb0GkATj/CFCM6H6uykaCd+6NqW/bX4xbJIM4BcGYhNO
2JrQHPqTkm9V68haELbph6i2wnV0JQt4/iO0rY/BPj8GZYhDaMf5OygytAODFNgF
MZb3W6Qb62UGroyPRAgu898LzWwBMp93rdyieEmJ60W6oagjsT99xKjda1+EaUO3
Kr3F6SpAYSSvecOVrr/viU1q3xyv+UU7yBKp1NGSIE4naOFCx1VSPrPvmVmPIi3y
70s8I9RQtAjm13jMYJH2pI67NNarsy9Euc3nd2jAdEvpoZoi57F3nOcAAWVIPcMi
xzOeOIztXooIM8Rj92gzmBII8f4sVEBw8OAcUsPJEZ1bfyEloNBi4IFa+lylq6d7
VakT9xCM+n2IUmrzNIzaOJYS1vZJhn7PmoufPRMJwCTJarP9Vd+5Qy383komp/am
1TVJ4iwVpIVSyfU0ENe5ksF9uTZ5UnVWa+gc6STJEIrLHaujvX3cTKrDIcnOuzvr
mbfrIBi4tM0KiuhlEfx1SFP/DTEocwvnjG8Dj9hKQRggjWA98hj2Kpj+0E2KIvLf
+mcsQr+2V2Q/4eFAow2VlQMFlAVE9u/Av/yOeVtVKJuFuALOHUvFZz3+ltnTi92X
Flw7PJlUzohR7YQlGtZnT+iPbz73caRtjFcELxt/7a4dR0427TcMlItreNrax25y
38pG+yczgoXz0ddPTMk/cbm9L2Awu7CTQ4YTpagTQQoxQBttQ+PkB4Mh1eyg9jqX
Q2qYSdFlzQC4kEiMXzJ1DryDQOmqyH77R/2Jo/Qbut7CLULdGLbgeip5kyLwWD9E
zcOX6gi6I6r1lizIV7Y3diaD2tk+0WPaFecOFAsUXCGHKwdH8eLzgTy0Ptkl2a9R
1UvWRZMIyM1yP3J1PxmWrwYd9I59kvUoFBrORn7jJsPHsH5YpRtGu/K9cLqUqVCV
Sv5RApLf4CSjejxlekiGprYLA0eu/uZ1zpouzprPIBtl6ehD5RSLzP/MioO46HBs
JAExULIdoizzfMY3KxI9aQBN+cJJ4hHHevnBnAVEOZ27AQvGrVDSs5KynBR28dwA
A0fdeIdGJFU1saq5WFYUFW+gWvU/lnxs2GSpspiAkLJmA6FVoKhI9nQrScOIaV3a
OBO698tWOXBxLNw5o5z5JNXEb17GOb4enfgIWOJLDAP7UbnCv0/xr+kkY+Msd4pe
Farqx0Wwjak+rM7c/1euG/5I4Ou0XK8xuM24p6d4bEInQC8kAPIKv07ge3b/0VOW
yW+KMPllgcQ1LWE+ZYtsaMJTl09IH2g/vcO3zYrO0XDsi5b2SJG+1BX4XzRPu4Hy
iBAtk/putsVVW/JX0NCiu2Dkh0T9TTRXaIewLF8C8J5kv8Y2RrSPa/u2VK4sfdGW
+2zAzeGZ+CsaXsljKoZAkB7QVls+pWIH+xfCBPPCLk0aITvjJ3zmZlEnqWUswcnS
Y0S7B2ElONyC6HAg9sBHtOHG6Lnh6NEWsAlkLwwTY3QTLPJQXSqJadK69MykyqkF
EDEQRG54e1Fx66g1O2Ub0mLgYmETjHQPEBQAHjyxi47YhWlL6/WfG5+MoYPRIbMK
8uGsUSPkWfVjX36rJBw2FCQr46247wapnBFIQ1Kl9AHEdAgmsTLzTRsfUcJ7d84U
UlQgsjJrRVlaB0oqWp54uaUhg0k9BfjHhl0YTm7khXBFlpXkeGV56M9k+OK10AgP
nWOf1nplDe8q2hU8fMo6TmUVoj9FfqBXC8Gxa8ADpWs0QSZKBB52kp/wrALgtU7X
/4kM3La/psqYNlED0ywMHi6xNd4PRZsr5I7rXV7urjkpeR6RZoGYrKQVaxW2IJpU
LVUuoRvq0b/u4RFLFBKWhZ1Q6QFbBUF0M3WKM4Og6JxlpEltF0RbRoDzieqo0gFe
3ekqqIeDcOOyo7mUG0nTZNU8TrV5sndf2vBIWaHexqQjnlDUXutlug2gSr02cqRi
D/fVX8O7USgQ1dq/0tX1P1FCMkLJKfqS/WvepCyfS2GX/qmeIrOrKPakgPxT56ss
TEP7nadCA/yGO6KYAVsUnBOLScMq5NmKBFJ/hGYNsqOgCXawSebofRXD61hpPVYE
+CRHq84nAcyX+HorAIT+/Qi43kx5CRUiLuTiGL0jBa0yWkQ03WGwFlp3ssi69JCs
4/OtGBjjwV0If+M1ngmajR1Fs4RMilqw6BsmWhlcQ29/ppNsxTDQn5JjnrYvZ9ND
goVAxpKcmglvUFCG2w7x7sjLEehK45neNo5R7psCVzu1RXu45Asqy7Pb3O2JYUFg
iP3bFiQPVUumUR9AU8N4TyltHCpIzbFjwP7WF+jeQmz6ENiU+JHKKJ9RWcOMjmh4
OwtR6msGZJbpSLuYCVju3EZWZJSnAvRotVfcEglER1ZI8jvw5SgQc8MhbKwuZGkz
caCtMxmCby/inLt6wnznN0wL619CsZzp+50SMGkOam0jfjESBW5r241dwV8e0eO4
jiz/oEAEbmPwvx7HZwGfZL+IOWKnZMSsM4gB+Hdg3GHZ0rbJjveJCkL359021zVE
v3vTTlwfDpQ6RZFeNnX5+3CQ01DGJ0CZIFvD8dNV4Abgr1/tp5M2IDfg92uELEFz
fv7ZX0W/QbC3yI4KPJC2MITcK3GB7MBQAcMM5YAGEjgjUGLlM5yDuQi1ORor2RzB
1V81l6b+re3lefPO+tQuJA4vmtQ2ZTCGRo5bjowcBtRk8ekPlNFiljk4FXP0LxRg
hbW6ESXa51riKgjvlsc+F9iqrQ3fFRm2f6vvnu+nFKG+8yR7+M1+ftdfwTC8lNsi
SiCcXi/a8LPEICc0RXhnPmpwbP5ysguCMIZ+ODSqVaUcQtMVl2z3sZh9lQSkPBzU
MbpYHErnVwSWMBryXpi5GUXO2nLjbjo46mESgY/3dLKg+Eu2HqjsHInF62zu9vGl
T0kbIViNCskOCQgCGoSPp6MNr6qHYCUJha/S69b9y4edQT7iNNiCuhYj8YHPt4vu
uID+C5fUqvTow0r6ohASBfJRxhD971B9HpCBENqzE2jYnKsBqNoyuaDbyz7aKpyI
rchHOO8CKrmRgWCu+WVB3WPSpWxUtF8igM7Gc26W6AK7MkPoYNJ0yL+gfW6VoFwa
hWnq/e+DIfXcS2loLbj4koGrqxw8p6Z28WzgDQDgfXyqjVHr8jgPc8XJmVIFxIqK
pCR+M+nJyUux6K4T7n4R9OlocvnQ7facW9OdrpR9evzBfyJkOttUmQdrp0TXnazV
Z3i6dVcxshdgfEJO80gm1r3HIQXez+cGjrtK1EwsstGJqs5DVdXcJ06sBD649eyq
o5r0rjt2Il3HETiU8vSsCl5iHROz0jgRNMquca26saO41jc3d7xVBbwGBMNFgQgE
uLjbmYDpHZYjTzSPWwZfAPYiywKLAOPFVFcI6dmLr5BB66BiD+FdF4g0brRHQYix
XCGbbVSuu75jujF6ijtU9gz1baZWe9sP6dW4+N+Nw1vlW0iT7MH6foqEELErO9i9
IByC+ePTGP0h4+3372LDmxf7pHLbKt5US1ANrxkdMyjm+WlEXOrpfs52Fw05zNLM
Uo3BV9/00FyH5GBLZe2gtwbag2jb/KRjQJD4xP+deRSYhuv2WHdkgq1dKnyHg6Za
X73v7kqF9REXDf6hAuTT2IS3zjO/dM/nPnkQLIbFiSt5o2HNJI5dtXO/DihVIhpd
rwXZIYS8+CwpUiJxg0J1WjXmqdNG3AoFUubNF53efyTp3RNhYXQaN8RdoYlljwZo
n7T9piow8ZyKtujS1f4114cmo7tPA6l6el5Y7w1RjJpIxL/Wggc16CeDw3OACTlp
CqZEV6HAmL+DAQp5d67mHA3pMO706ClbT3yn0NYMGPVkffQclM7X9EyCO5TXR0VW
o0j2WSD1MHCX9025GPxSA6acMUlRVsLKOs/FmoR3gFgZQj9iWJP2wl7r/vMxRWKQ
6HM05Oq6NtApERvd1WZLcbrBiSyc2in2YY4V6kFIOzx/2DMu1yen/IQBxOjTiQFC
Ky0CmZ5akVU4GoF7U9YW58hvYFCqzHlT8LX3+fbB1C+nV+4uIf995uQfpg9JvZ8k
jEALLIDlEZLNeeq66fFaLRvy7EyGPptLsb9U//xaxvLjto7NiGm7FgdufB1NR2oS
9spGdlW4ETjaerO+nXd7dZ/4AwjXg3ZdzRudYZQzvYON9cAewvNPNl9FIoSRJlPp
EIChxVD04jUy6ekUC1hftKGhI7mp1+GQHt7Qa0nOo0qcFXhTa7jTnS8MCrtfPecW
FgvkNbh7e2mCewR34p9WdFtOEshL1BMNdxrOIVk/07Yv2wV8ju5p+Pb8imuQ5fSh
wM7yAAs4+9iO/4oKO9H6bLu/8r1LqxiP/DckPDTXow5Ki+T7swgQ1B4aop9q4UDp
cThji6LBbm/PRG0isuOPAcBN6fTwEUzN/c+3Dqs5czlq4VwdnLw5Q/L76FA30ZAg
UmkN0MEScPdb5EhysOGuRf6uwwOLb2vOT+nIAZFot3UVqOCxcmHFyeuNUwacgYvW
6cRRacJomhTGVktbjyRZ/O6anIdmn0AdvtZHaT3HPexL1QeDy1UCWi+GWcTRu4ka
X+CrXM4e7gLDZf4qTYmH0LrUcyyjLZeCyEXYel78K28opPHZoDNm1d5mDpupclKC
f+nuFnMGiO4sSq6d12T57cPN1uTJjEiSqrda36U2+vN9mgNRGj5LZ74LI1EenTPn
P3mBUXwlHAzEyJz+vGUWLPWl8xwHceLqHUoJNIE8v3J+i4mWuzt4qYlyvohQcF5b
gOf3l2Yqno33ms9byVnepPf3aaIv33tMgqeZY/8COjZpUZTvbpjEifnrcifxj7Ro
RQoFeGwgA5C+o185J5bwazJhaQxr4Vv7Rn0oI2gO7gGkjXvkeBXbTudEkxBLYkUN
dMdLc2BE8x0yo/Z8IiXUnRCRz7yBEi25Hq5EA6yslOyEU7s688Wsh3dhANNymoao
C3f0TbPXWBE8OyXeipKyv7Hpvq/hEZ5WMCrdWoivASFqIhgTj1L9t/iZtmvlQ+1E
/17zAKSkLlWGVpbD20Cp3KECEimatMv5v4YqxN0bi0jBtFyOIqhYvflfnoK9JcvW
4DjqZCq2PLUv83VqIyPGOicueIsErFRNHyoRNiHfURXNhDZWbtzzPp/hcln14Mou
31wS4FbizQIvd5s9jzSV7ujdpo4KC0jN94Xp95zYE8vD+iKD6eE6E7bk146dkXkB
zVEKE1N1hs152sGSzq9KPG/sDRPJlD3xSvxe1hcMW1XOMHRAeOksIW2TtuBV8MxC
EAwYKW64FF66En8U2elZy1LlKWxn/+Xqmg4cKVcIy+ZkTcYZY9CSlcdiL8XyRZPG
LVqTxGMwX7/WkjJ/ORXnxwiyDS1O4XftWYEjoDeqEyZwXjimEvpOK1LykFOrwuIf
k0F48b/D3V2L7BZUTwCn9SqmR06ZtafNJWuvilTtSSXGqUZb7jdgMU4iN1ckvEE+
1DUCWCO4Beu1kP5XHZtb0ilE10AhlY/iRnO1Ahka1XhQWu0P6ow71vEpUyKt6Bs4
S7gvxUsdRHOzG90pmEDt9m4wbgXndgzaS7qwveo5ycj8zBQgkd6N8S/BexGtcHO+
rJdX8S29rieuM/8RRkqyWi7Y3OBhgSny7l3Z7Fvw8qiGhS7zjiu5idAsXSX3IAKf
gl0/f2RXSxqiqcqotAAY/UCf7w1YVvofrrnPNUo0K9Q4WjjqPwQTueXIoypBlMhj
Fy1vDPXf0OAq6FpozfQzf1uXxBkk8XoN4NS51+eTwF0nYPFND0WHriwOl3f2KQrB
QJqtC5kx8RVHdqnF8lQ8E+xYJEac0w6QgK+2QPlozd/kUBJp8HHc5NAW8eYQ+HOi
ycwm5HI4cOsrGotFg0Yb0Z5djnNpN4+sdXl1gRcu+N4XBvp6DXb4PLTTQDbD0k3E
F0bGCFtwK/aeYX6Xc57tX+iFOgXxSBgNZXJBZDq0AKmE5wg90sm9CpIP93bK4pfK
yjXG/V2nmemYU6xMyzbRzfuHEoN91qLVC4wBrlt3Wb7RGTGkPFF05JVMZ42l5bBL
naH0GbCZ4qbRCce9IFXbr23yNeAufIR0zBiImwp94v5PUNyHi3BwkdeVKHk/w2df
ejp9B1e2altw8faOMvgH/FO3f9+zs9EpGQYFMSmg7UTfTjoRKTG4xBZ96svVm7CN
UPf/dtynQEAtYMV6rwupBak6kp+PlTW46iynjg5fCnOe5SRzXiWFS9sCp3r3U5mG
2nxR7l3OOTKkghBCG2fyXsDP6hW6/kexOUPP/cJzUMg++RAQy1XYywbY+Idgc5oi
me3WuxrI4ba7J39RuzDDI4LNwEHEGXcGpTBSa9oBkIFe8XaXAO43GUXYvvgLcWdl
IXl+LNQY7C6akJkxHXDkHl7A8pmFuzlTHiXPlFsj/fo7onDXopZtrunXDR0td0Q4
L3bnpwNz7LODD1FXiGl72/54DpJILdbcnbLgwn+Pg5dQT3QkC9Rmb2Ax2lzqtw3G
mt6y/mtE7xSJrAF2L4d/yAbL2SLa3AOqEshxGidJOrY+ffH+f+Ws8XI2PqUULbBj
qRMp2B72GVRS1r+RNlRgeAdUb34RYv7V/ACQurermMhQ76niPoumR8VwYsV2UtuZ
O2rwR7LlVgbqv96i7+a1ZQEhVIMv1swS5dyFZfftqoisxfO3qD/GEdQZkdsXJqP/
0QyJJ5ogQKPlo2vvf/oQzvn20nIXglib8BATvSaII8dBMpLmqF1sAqSpaNChJsvN
mtD3WO1RJtmt8/U09G19YV2UJh3YUmEIM6hGPxP37OBd5jrJdQxjYH0KijwdLgg+
yC44JtA4bLhDRA+I7MtJY6TmVRZwGnwaykfyNuIIm4c4JhpajyMqtCPyfiVLvcUT
4kD9hlD5pCJdepJ9uR0IxbHQ9jy26ATOfmuP+kC2WpqXv5BLEB5Zb5EHnEeHoFtr
pw442RT+f4p22vZRoDGjPclGUGT+p8CpyEh4eg7WzQC+QYJW33Mr1+LAalxy9odH
X/1yTauMJqA8hMnk7KMZsZLyfFB4oDUcSN7CapLyl2cOjcRclFB/xp+tKJDBzilR
8aAW62I+4H6T9PPtPoghUtuaF01DVaSsr7sGkn/cdxT/k+Zgm79g+5LPibS1B2W3
2h27L8LES4qTZMXA8a2aG0Spu/sZlKeRZSnZz2bx95NofMfB3+tyMdb/y2fst9He
AJ3SSFN8lNdxivD/bEyq9zdXpwQKg2tWMefL8hEIe4DFU//mOLSpa7g9a5MneB7h
6yySVSrYGo9K99lqsadbvlY1JxjJg8Zk+D9gHbaWg4MYQuCKPu/m7DFWT0vPrjtF
ZAncIAAIfpD7gL/0ZLrhV0kS4DHbUwkuAf67BmFqaAA6p9i+Yw+uNGPMZOT/BkPg
nvqG5UaA/IgYA+ooFppFNz1+B07+ZyQUt8XC59pMCTD2DjuSTODxA/FfTRhKXZbm
M79hy+W4jZjo1hJGHzwt2NIanjnY8nnQkXyovh49qyjhk6vBBmOcrt8DCUj9dhgF
mgiz1k//nNtV5pIX//g9sxferVoBPRAMCh5EbQDj0Knx9HTYcwAPQ/EE9Y7KcsVz
zQBf9QT/sMbCo9uKUuKvqtJPrnau0St2HYy89edzb4SMUMJ4BvayCnJwMEnWeupf
N2UQCBWJyVZzfGPJrb/2Ce5AP62Fqg8Ere02Dk+uRPL7YgCN3EEjTaWItDlEvHGQ
S6lzfvwlmGyTZOcmbPoWRqt9AxOAjyOGLJm/R3OZcp9zOD8UJahb5MWmqC5a5OQh
W3dnTn0m15MiCehwHW9a1nYq7Ef3krmV32y9A1PScrzsgrvYXLQdzasAHRnbviIj
KwXIMyHlxdtOjbrkC4/5S+mrjvqgl+DSJoV6tnUB7Rxk+LxP4yC8Up9GVIEI1RTk
12REhvnu8cziyWuCwCjWvqPPk7C/B4Rnhhu4FfdQOmenWJvQw+O4qqDTKF2RG3xh
jcKbI1akTIkX+azxgqIng+FkdpFVHDa19vm6pd3GYG0eG0Yg3VRyCT7L5FIbYIi8
hPNs3Z0mJR77+T2m3uwgsW4v7yb2SBZFj8eYt4RIuAdrEBRG1KmehlTxsnr6egd6
esYu8mNPQWjTixuZ8GpkR1VFuflV378rRRKPkBzFuQnI3LlcZ4Vr9sJXv+AlehtF
xdhHuhLe9irJTIBg5HVsiPNAqHf5NRpY6zknHiRzcI8zqhGB4unfTwLf7G7u41T9
HmfVRzWiBM14aRYYpxJQryWsKcCYTV/XDTJO+3Rt0C48xMcOvw7GoB/n4xd2CaFP
EJ6MPUJOjGmImLxnfkb7E6WjToSkZoXEz39gpYrfpegQCXVTjfWNUmokI5dW7H2U
SnO7fXKNhmKjCJdu/PzVu4AT2vMbRRKnWTG4uINMptsLteTFz0/CeDEfDLiqUSf1
79FUf1wkxMsPbaMSB45N841pK+SaUFOPAz/uWZ9pv4WlQxzxP8tolzXvOklEQYtY
KALa0bJFdRnZSB3T6ff/MEe1ZPGqOF6AvjmuZfh8hXaov9Qfgjn+/vJ2xi6zmOH9
LDCCK1ZDzo5kDcN4/shXhgVHffisOfp6U+BdMFp39n7jerqw3ALtXTUCuEHsP4de
wRjXklAF2c0aYocsRlJPM0I6JC8FBETXH32nOn6utTgr7R370ZQWL8Mq/tKOiCet
9T5mv3kcqZN642C/jA7SH3GSjfKLzPfAPPKSfqQmtp7j/Y2gk/NNtgalylOEd1Jg
uF92Cc3XBAzIqM12oUDd/Jak+mZv2kh429UKnkpJPkva5hCt+H/eMFvotHbyioZW
3VrQyYkVVu8PxhZipgTRMTLQ/CqMDnXunuAZFcHvBBDyGKCxHYf0zq2j3R8YVnyE
ttUhcsfuCe6NKZKdwabr8vysk31yJ9MH1CIPkhhOUIm6pvte7P/QI9EnAsR4ipO/
TvnT++Eel5jufOiWOvIZYWAfmA28MW0zlYcTSlh6sIswgwKbjaiIsRJh8sQEUXv1
IVmS3LXM0yFIs+FDpPdyRI3GGKXybv88KILF1DmeZjk5bcSeeBa/zocQ3tBDXxlu
ZxEbTA4rcv+K5x6XpnQN/Aq/sTMRM1T3ZnzR+uiy/H31oHxnfzDO0mfhJkbPLXT6
XafGFOEys6RxHSM+7N6lCJ5ThTJwMLOOqh1QZ4yB6hO9VqtJP3QJr8Ipusa4jWrO
gR6fJLq7jSNhpaL6rk1SkJSVoZaKtBk5D8AqOoZo/w8WTzEqFoDcjB5BbhlIzf5i
431onPsDq+HDFWkAEqEXTeGEmCtpU/5ilQcNxg++MeX9cCLAx2BE/E2GB93RBa56
dKouLF/UV8MwIkDlX6OyslJr3EyuIBLEReE/+3YLkC9lVZTyqZz7iMODQvPgtgto
jKRH44DZmZk6HlG6qfcalYTYLGCzyq2H56+6M9DSRtBTiRin8rlTjrsWtuamkgaF
S6A7wMPSFCQQy3jfW67Dhd7PmsAWuAZtr6az4utC2YV6OM2NcP1rmFEkcZw5/L4u
/auF9wTd96pbO2fnpseT6MVwayLI64Tv3lUhk1rzyQlrhD4v2kYc+qvzI2enJIbu
uikbhcCRiaRjZ8mYT0fridEViD+8JSMj6m1wN9DAbea/HAwhms2nUzeHV1DOP2tx
2Gn3ogEkFzDvf3qveTkxvO1jTP3rRWzB0LzcC/9vUbbvnlqM59eBxzPrbrsjnkKd
ji2dmsRtnSKyb0cVWouBZwEomTh1y/TlrI/9GVDKM+92H5fDSHnFFgzyjOn/qIYN
icFQu7gQRMWl/ycEMNesFQuDcP0Vad1Y0Me0zLl5f50eBtrDXL/DHooXkGkErEdJ
ocLwt0STM4ThaAb9dDTDvVy4drQx4VfNeZvhR5KYV23G22oLlpuBE9SjWI0Gq6/t
MH4doObX2BgF6/ZaBn26Pp87qFOly53o694zEFi3wBcNRjlbCFsQ1et/BVeUp4fp
EpZB3L5AEDMYM25uzDjV94rwIGBn2cpZXwWPmhg8K5NFWI0VVKxDn/ffHp3mLcDP
qKq9WrBG4ra+aMZu41hSkXo+27YYNdtj0PdaqdTS5w67TR81GfdsCty2T5GQtdc4
MYVd0ovMSDxU+Ke1wiB60qbOdwLHApyqmPP06bgHZQjuetfg6NaJ0OwYlBvWSHve
R0Z3LJEgbiSxmNh2cu71BkrEJTrq3N0imayWpFaObqpf60smQ6hRDz5VCyOl69a3
kq8IiD/z+DTU9taJVaocBPLfVSmfl6uxq5RkHVeet70yNt6pnIJVEEZt+QOcG7VQ
+e+U3oRr0RqnOKDZFGU80IIWQtNyxa+0OmRafQgV0xwitKpaLczaI/R9fYrTUtdE
WreMK2kPjjzTxWJyerMjxAVOleQfJf6H0QsvlGVyfTZknNhFgIe801YycwX6cDOI
T7VXTSkdtfJUx2mfY0UmAhUx3MgauuNUe3/odOtUWpH1GWog4cLoWGS/kWbTC3Ss
zhXImezUccMb1uV1p9jo39EDFvc6nxRPo977lYekNARnCBCz/AHxKd/lIPeutmhP
cdU40DcQ+SZPUufC74uU7o8CgadFO2E+wY7Od4yoFe3mlAJEuLmBIhQvMVp7LZkF
a02kmj0QGrcQChMf2cWroVJ/H5jhUJRoEqGBAvs1ha4NDE7n0ChsVbCOTfKrQsrD
I1KL3f3h+20sGJUMB9h7zQQ/DXlOXemZmHDLlmMNEprPjCfhe7pYF0f4xoJnJqHy
tSVwLs4cC4c+Fgc/kOx8gb2QIrlQnWtLwUP2vu4kSBd291Xu2hP+W4hSJHrZfkWg
b3XVDfNXNeud0o3rJQDWVLaosr2+vdE1ZJhH89aaUWMWEKYb7F8yp99CtSAz0tOG
oCRmdeHRqumDNJAO5l1aRucQpq0apcbpx/TzIqcPf4SCFzBhq7ObOV+KwlXpuJs9
XPDFxnp1CinNhjdDvglE8rVGZzuXkxtIGK11KDn2BKxd0C+h1JV2DtPGC4z5lkF5
RYLLqUhGvE7pm+/TTQhtTSYgxP7PlQ63MxgmNFqjfmPG2TXkwEKGsC5rY1d1uFwm
PbiPZ2jTgfWaxodgvJ4tfPEJBse7xFUyL4Inw4S60y5Dc59LXg/ZzLEr15ywsHjv
LIZ/1QRr5rXED93wOkVzaPzAvGm9+QkpI4qbHlfM891SN8actvCr9BRQP6w6mxPd
vxdPhdW6rkRmgtfnD8NxpboHnAoyXGY9s7tBBu14hr/YgpNtS67T/GxaoSdbOc9K
TLxUl3sx9LaArW18l8wLHzlCKbf3hs4wFtHVdBJbtqc+jTpBfHiTidI2FDqzBV16
3/qNAXi0mRUbcyPVUDhKUA54UQ6UfIRbjvGUXXljDABaeK8fjk5wtP9m18vfPMKj
+o2ox+sPTuqw0lC2jkmylGDanuai0zTEBNwHMh3YBAvwj54yab6TLxiQ1rKOqutH
YfU6ou27WhhV0ukIUO1Ue9VgTkW4uM/JTOarkzNs6+EUZdRHziexFdOeWdc3eRzJ
x8a41MJhoQwLXtiD4lVja/TNpffrz97LbCuXehodkwnRSvEs4wp5XZj8cNQq934/
Bx13amkgaLfL0J5CRwvDMkpO1pZ9JqhWK6w5U8passrEn+/9RoCg8Cw1Fd1d7wDp
FnEiUVEX6Y3fH1z8/VQivMaO22/RSiaFFVLfYMYbvxjhC92YKFW8Q6ctNSg3U+O6
9CY+bbrihgclV/cE5jo0jPVk4nlKK0v7BzJE5dJTDUfk0y2k/z/9rTrmTrvM0Y5w
FABohfoK35gd/ppfANfTR+ILcvg4NHtNc0PqyMI1BcM23zzcjSWCUR94uspDI8H1
vEKgaO382AUaHKnMVIeH7kmTvoDkt2gIcdw/Bf5sACVqNMUPg221Ft911I+wrKni
IAYM7Det+H13B/dGjZ8hM7bnHPEhYdpviTCtWzN6nQHb6DDqqr6bY+ZtoyXmQQLp
QWKHxcJfjMMFPue2U19bUqKUFXMAvfFFw7Rn6R9jZorqQIErY8Rn3/xJvK3Pr5on
aGCD2eNX7lTiCwZ/7eTX8w60ufLROKj/G0dZpZnJAQqa/EGwT/fkGsIIbByEpzTf
2wTqAqfxZxoMeUEOCsLoggG0SFfVRWQc6ELNAfMbnWLsUCCcLDQMkVEe/Tl2KpUa
cUts/cGhIgrheUVWtHMZuJTjXDdMLkD6gZYwPrPFFssDDtX84w8o/aMJqvrGoLhr
+BGGBAduKbP98qjx3dR4X0wH7tpIpxCwdMNonWcDxgn7CMXAtDb/ajHu1JLj+Ssl
PpXkoGDe0z5I85XPquFkc3Aj53mesvdEiTrg7phun8shlrvVSe5wIG1mUFBntOhN
jxyKNBXvC0oouweASN5yuqUGpbuXresIZbLkfTRiuSmgRaoBFmvbDEHm84qZqayT
7E/kDggo8dJqc2oij84l0zptaihRrCpkfgPmNscNoAMrVhNrgY1vPjOIdEqmKHcX
OlaJX8wY+cUpeMMF6d4wk8FgWXQg6V6eTyddsrjmM5k9cTGfTuQoyvi2FbqmRKTL
zcJWPrgtefX2bKDCTMJFJ3ete/4XEMTosK5AEkOV8eF1lTdGRwaWJnVnezZh3iOV
/vWVVFdi6c4sPeAP+9NvP13jshDh2r1DtiKJb79VgjCzMk7c3hWNf2pCVhMfWkf+
x0z4iiFJbveQeMVfExkGmOvD88Q5oQASSYRGtF0NJfQhIogCdiU8NJNCcDIJkxsN
AYtuEEb+Av8C2cCzKBAKs9F/NUZTfslTxtwDkflRneDhxsInCdAQ3oQC4SKv2sUX
UPtH9O34J/AoUA0iLEv45zTTM+6rMubFSkEmg5z3dCBnX6hl2/czHmwki1zTxkgB
e3CxHCNDp2OvUFKBmWCEyLgErBxQZgqGzdC16TuVyjCzM/YgUganKRcWhty/4PuG
yGMhNreWHz558SeuHewZma0x15bYuL4dPgcBUuXTBZVbRptbem/wdWhsDyjz07vt
em8IQvQcb5PNALRqYBZ+bafdexm3ouX4qO+WZTIML3u6m6y2Yaz9NdOMU/Yoxsez
1YKlOsLhJh01XtaNciygU6ZUoSWQZL20FdxUYTJOkuATw4A0Yo+WiEt3uMDHEo/Q
FBKWOyzNEyGEmcBDYMqd+ih+L0cDxhnUVlxr1mYe/Qvdsig/ymMqa4w9Kx3BMdjv
zFglEpDv3h1EpwQgIA0IQToxU74126trGKkB4Apkyq5GfBNJvy/Ne2zRwMd+Sxql
U4RC3kvu/HQMMOPMqQVZQS3ht4lcdgEV63FDuVY5sVgvGtAQ/Fzh0ARwdJKZj42E
0tmQGqSsH/y7IisjitGbmAqrKVuf7pn2fIlj2M/Gx9KG2/h6g0MWzUW5Zav8mdbv
70n3WLZR8le0J13Iu/jfsjTP8mqveE7tMwmi8ERYcfv1gbkzDGP/nY81XWi8t7um
mEevLqa8HklNUUFOC/BSiiKaKC4k8NbaFHoNGTlGgHFYBgJB5n8ZuqP04DH8aY6r
ypaRnyleXMCP1xzoAw1R1TPe3PZI3sNCWXnaZfuT01bi+uW0WEKarJD0WGdwk17M
wb3EQWzGMjasiHwU9ftIP0k3ugAr3bXQHqBBQBcDTrOFbHR/VvLWCxU1onmdyWu3
uOwEHKbb4uWd9NZeMQYNpbF9zaCFaLXXJBPWDDJ6JTlPYR4G1TTc7lwRs2QQPS/+
TawNbnLcWt6LwUDS/aVyCZxULXobIxbPBzLhCBR5mv1ftLJCNXdVoUFkzgnIoT6E
NDaoecmlY0O5HJFM3v/nxKNJSMuypw6rwtyer8Jy5O4uLW2sIAp9Fgn9VSqbmHtp
e1/f9mIZ8Gp4YbnsOTBNdKEPfPdjYc6wdhRU199GSM6ht0sFeJj+sf6KDEb84076
mlR4bY8TaRKbpVlPg5OlxWwM/jLbf5zu7cNfrwi6ahwx1KADV9g6iC7Hionn0VVv
6uIznfJhGnK7yXAO6vG2Erl3945tQbOCT6fLJI1udBCVGt+ysSLOnJwWcSWqLSPH
G0eJqEso0te0/404f4hHGjVm/7hhKboU1PqpL+qWI9crgDafeLhJ1m5ohLcyjmNH
oXlGojuQ0dTgKeMj4tNJlD6cqoICCCHK+24Ex/6eYTF1a5Z2EKJ4r0R8mEQ17cKs
EpsoPlG/2SyQRqKPS1w62omRYzlB0dfdCgoIFIc/CgnEwzZVvfTEnVmEESKaBwmR
CGgxa9aRMii66Mvo24I+PH2k6yPIlrTu7afXzxoi0kzjSDXgXN9cZE++cR7dsSal
iJYf5n7wQNP2gkIVb88dF6h+czU8xqQGH+pd0uPTVJywytbtkXB8fhlb6+k+zn6p
p2JIWR9etwz1VasXLtCUYrPVdyXEih2P2Lha3b58qGujt9MjIphhM6zSosW6Nkip
iMOnEP3P/h2ZRFqT5DE7osbtYBg0A7DRo0hTwL+9W9bQBS2ziUbciB2GAO1G760q
VpM9V9KPv5zKBlfw+UfjcbblQZ1OeqQfW8n8E69AfDu5u5lyhZzL/fQUfwg/Rjh0
Cvp8/iqbEjox3rqCd7fB9EdyVEPrbuZE6vOOWnAEBFBnDF/N3FZFSpK42TL4WBBN
+u/yxcunY4xaIkbK+CL77RGfFbIDBO70zIbfjy/098aB2giqMPju6YLooZlVlIhI
hkvg2UhgvShe9qyvlvTQAYqvU2V2qrbKn9simsYNp0r/CNHE8w85nDGGeT+Fg4uD
c1f02xY6UB5E7i685Rh9ov6Vl25BF/I3kenl141v3Ysuok9G+348D5hSqP4fCQEl
FZENVT7lHnHxyjTvOUIKTvFbfYK6dG0N7+xXcvRjzEsMCyxOYxHyLsgp9Ys56ilk
NJnEu2WQQUfl3S/BW13NL1nf9BPZaVw9RwNIWi98ZQBfhDWQwFvr7UUbdeifqQS/
VHz5E8n+zb+Cvu393f38zjK9l+0lRcvAIwY9y2Dcca6jAHJCEvfFJUiqXLMox9d9
Ws++fDJRwSY6ZZTEI1s5S1Bg70NC/b08qt9S2JFUC4D4AKQ0JXiap6WABgRhCOyM
WPK7oiK+sg8Cir+R7JGJNwfcUNCQavaNYh1xfPnxYNq+dlSLEBhnmWgcUJDuGS7K
8m+R4AL56LpMg0O0ww1sw8jeRqCu7bnnYtHtnjS4oiwvt3uOXBED8AqBX52E0Vnd
/jVmq++F9tfS9VfgX1Q1cmxL0Iw/SBt3xdlYsbPegV8r1IFY3YTLJkIKAnNGLDK/
UxZXRREpdhN0H5okNdholJI9LGbvzLxXoLlLXOH/JODP3asQkipMDupNJQ3TWJBa
MdXXs4bA+B6A6n2LZ7CnJ0XubvLKvMr8EPWowDVmN0p5uhBMwgzYLX/Y0gMpHSCt
qAZPPIgOshNo6vANrQjCQnaGa1YmCaOsR76FtbYqVmFCuRVeWy3InOcjlTV1LP/g
e3rz8AbdXahANaBMTuIx3YbiYXqVSrB4I5vVcLNn4ZEX0MRCLzFRRa9tqntZNMOQ
lVibFki5dLfjrXfY861xw/UJAJa+wmAVrHbWcIdl+aIK7sXQAGXPjS4FveINdqEm
DJU1j7I+8xIDlUJFQy97va8su3YJsx09/zDO/qLivOiJkejQ1Pt1TE2MgHuIwtke
+lpC7zm5oBapN8UKLsN1OutEawr8tNLW1URNuZCPO61PwNAHZ2XrTVzcJ+A3O0LJ
Im0qDzz0icTfa8RtAkTn+MYQnNVoSTzzO6Z+78L1U50hbh6gRLweaqN4be/gLRcv
75mJzkH3bAV0+zfEQ+S6wMBnGUbxBTO7nLmDX8sqmqvAqtF0pTuyUejI9RPgmX9t
K3UNEFtd8rcunN/5kne2tI6eRaZRh5KisNZfSXmr3nGCj3G3LXmAeNR6ixux+4ys
ukr+gqZyXF2MLrF67r1bfWptlg7MO0iPpxQDsX8NrGj+jaszpc1Y9T50xwJPyppp
NrMbjampg90KYY8K4MVQpaKaWAT0oI6UBw7RqH+XVFlhhSQA920qollBf/p91M9s
va5GhOBFlv7+io/SX/tazKyRDbJqve3Hf8q8Z/Hgx9csGD8zcp68a4ELLsjJIsS6
8tQMZhX9iFqOgcGKfIDfo7sxUy+fmJaDuZi8nzzD5YMBcYIp3njTQunLms3o1CRX
uPvec70mP5D4JfLsJMn2JaYpmJU4Ac0mXccQVxC+4Oj15byfEkbM64tNjkspfzTi
4kqLzvzuLIShH2F/W8K8fdvyLI5kfxv6Hi3jRldeJiqT6X0pirVPjQ6SSs34rsCg
Zlg31sNTnuh8H/JtbYqo4BP6Wd8Kbyb5UZ6hiPvDAFXSrvco8+C+JB2284X0yqky
Fyn2N/48E9KU0Su6+PqEFdYU1LeL5gDceg7AemlRqZczwVkh/WFxipYkSRYohA5o
toYDh3DoW7ewIz8Avehb53uXT7IFcysScB1oyfmsIfFstfleOkYXLZhJ66tz+oQR
9RpDnD9lIWin61O1rh3n4AHvcC+TnTw4dzb/yl3G9/WY3q/rrorO0JGGAWkjhdWF
FkIOd6htP/MlUV14cl5R2D9tbZiYndvBpYnEliHn4la8GtC+EdI9PLo1LmhvT7hH
ZaD0m3JyflTb/QG577ZeQxUJhpLneus7vegADmV853nCrnRL0iSLPgwI/1L38tJ9
NTzhypW6x+AoHc0D5gKUuB+j9r45v/WTsiH7jwq4ONd3wyPrvJoujGqtr4Lov2Df
DoxgWNggLi6E3Qfomj3KeV5apc+b+hlY/BHNV8fT2DGxNuvecd5ZP80lhoeCFA3M
AiKy+nh7rOE27h0lTJciprf5K1yURUYklAaGToVgF+UWtsFzlTV+Gl8sc3eRqp4A
wLsXzIQrUpgSlm4ABSMgC0YR06lkwK2etbkeq8WXVxmm++dae71HthXrIZ3THF8E
HsH7YyIpRuzzNY4B4UGDAz5CbArqFoAS/7XlJyCj/28inIQ+OZBn+Fssvr0ofYHU
eMkAyYi69mW8Q+t2OyXLQs3IeEf6DKuggf25ji4ClCC2l6EPZQKHrsyD7nv7aP0D
ZQNkBzL6m4TSkLXRc95u1R6Bpuuer7TIWpHYdmFAuOJm6HsljrsH1FX30Jjc2bMB
2qGHtAAnNcDX6Ya5RH7hyNOArCknWnBqNCsqxzYYN/IzFo+5rmh6LaS0xJUqs2e1
oIbsbMoAtpyYD/Nd6w9ryyofTHMxhhlXsPHQWNWVfhNjT+c3bmU0az03q5VTdrWL
cdLuOoan2h45S+x57px+mpbghunHfdHAwpT3LF8IZ6TbcXCcSrcbzCX8MPvqaN3J
tDvhAA95QsmtYos/tPQvfCzpK9stP+MfDq4K2gEl+r3FOveS8cT6yWNErfhIlShi
ShvPC/dILPCV6MXs1IxcER8iR5Aizz46GSXTyUg1BbH5+ymOhPnn9aMt5nH+b5gO
rWXTdQrzpnfssEojsqaYWwjrTXFzt8qhNGlQxdrY32QHndmUHHxrOe3Bpu9Dm0uy
bUB2fXZdOpkAmrPw9KLxLCs8tJh8hd9FCdP9EnK9OVYROeJ93vcgj3iKC1jgsPkS
U+ioXeEA+bk/gaz9KdESmP63tuex2/J1N3TLiKbfo95j+ODbNYqXhxHAv+KuKShm
0rc0hYGoqWlu3s4GiHQm8L0ZzlMXqByPKn9VoJtbkeL4tdj2i9k4es9i563xgbyZ
zoPkQR0Ov70X64TgOo8JG1RFc8ER/bA9nw2GCyTu6+pMofGWw141vqj6k15ZvFLO
dvbLYL+rHSBEAXwwC1nVTQZAGbI1NlTahK6HJiKCPf2Op5jk0VGIo9CMLvCBHHiX
vzulJDfuhdCXxvwG7wZ/Ih95heg0vkryGKrTxHK8kQTjfNHCzvHi+vtow12ilTHM
P0idoGeboSk8BRnGMdhMcNImBgsXEKU8wzbtLcPdmae9FmTtw32zh3sNCCoUqgvh
Yuhy8LqyM7IVvKFLY8erPx3MV7riAR7MTegJ0JwKhv43fnCLqsctdvcqV8tWCk/B
QnOPj+0cpYWlqyhaINSkUghOyfbvffm5YfOzknEGzaUe63vqGEfgYEJsKo2vsKkl
7iRnNtceqHANZWba9UtN7vFjZH52SpieI3GyvAM+EGVkNYTRa26bPpQfuREmrtGo
1qtt2FcDSNsrRkFw7SMyzFWWikuK0Ce0ziC0UdItAmdECeZ1jKXRjqHWqrZyB4V+
qUjnJr3P+PHjCYvP+xU3/uEYasAnoqPgXjgCt9lZQ5c7XUyNs1lblybKapLIarem
gZ9WYZObFFxlXgH8nppo2UmBkTVC8b3trRhLuSZ/uzQsewxHhsyqdumhdO2Mqw1e
AR/dBbnan3TUZff1mKiu3ye2STvZaCKjpQc8Ze9jQrel8+llbft4ppiFPQ4Feoyd
MXMohmgOpRta5djfp65jo458gC5ZxiyDUHYrNnLmpJy7D8Qkdb1IxjgPvb+QMEwX
7yCncpvfivz4Z+PMthgGXJDdM0k9XY9XqAd7JGI5wUsivTCx7ydEALWyKExsO89D
i1tkOh4K/+RC8MWXPWhA1mZ+wJWGNz2gdafBQ3XEqqSL9gwiBAWzJ4engbH9Ye9C
iDvFYQPLgs9bMhkmOr/fbapdyxGe/NGc3lNRXgS+Q14xXhPcTO2+dULx7S9X3Sau
CaamlRepsSJlrq3muHs70v5t867kxiEVQFryAgNakAzfqR7NabQjIk1YTPM80QxZ
uwQt1t3TDweIxXEfKyocb777gqAmI8nRSUkv3b+5vE+ggA3zgK8TR5/U80nuMfFZ
48RwLJBOlDqgbGPVsK6EIGrclyw4vhG6sMHk0r4dKPQROKfeOeRagBprkG3N0tPS
KmS2MidwbaFRP4qCG0nZCrT+sfzupmDcnBD3mnSaLYOdeSb/9toQyydM5E7T8T66
bGV3+hDZu1ztbX03X2+XIO00f+gtnNhZCmSmtIoCvtKJL0pAk9aS3GAxD2H7D7bn
FfdyduIbxTQBcxlCF7JIx8Cy/RYHjfEBanApA+2tnPXMNwb+oYcMqvDT07K0fenI
Vb1DHOwROUIn3M+OQ7JpbJFJzjf4TNl3+6ijl7SLE5+VFSxljlD3e87SeC2ACK1a
avB2p2hhchvfCyDiXAzSzqjvHb2g7jQhp7iu3+xeFPgDdUAJfOfywmsixGxoR1sG
PV/Y8CBduFn4tdIpRReKwgDI/4dmg2MUT7jA2+I+AYIJx6NBVuRycsPn59GpKLe0
9S/IBWDc7nyl4F7qX3OCkvuP/WJ0OWt6HxFdvM/Xw4SMkfcQtIO8GH5fr+v6VxT2
3GEPNNWyxYWPcRE2oNFFAVtyvgZR/q/l+QRisZB0LlJhE0TSxJHIhFGEBVijBr99
+8AAZwA6M1Uhug90DEKzosNO+/VtpbtzCyaS2sdqKUHGnLc4u6Pts+p7VrENQcrh
fB28+m4yabP963ADhJOOW4I9Fz3XnvXp295EW/mi6+AFcOnIWLRCDs7PsK1iybfT
zbsgfm5P33Le49dpn5P3926QYC1x5gJ4Ylj5CArWZr8hZM6tEfFrUFBNuhz4V6Ru
xRbm+a0A4kKGJXgCJh4LGylIb6BW7P+WY6JuvptbfhnRVBGSYBOI8KQTM4IZbEdx
MBCA1gsjs+N3hbibd7IDKz1NNzMHuelAd+kWrN0mi9HTJmP62NGsEkCCxdVDXc0P
/tNcGaGtIC2IkvnwZ8UntjffDVmLUBunfY17yLLSaG+Yp1JtUlwNbnK5gFlHEzjb
f8FB4FMjzyDIw7WH7uGE669IzXY8NBIdd2aQ+RPkKbrgbKryV/kFQr7KdKzwcesD
moeeE0CaGTRygT87k9c0EtYpyoddmgGFhoYEQPLqrRO73c/nvkjf//yUHbeufu17
siKv33ab6R4e/D7nR+NAMCoY9umswt7EM+8e/7OqP/VL9Ls4eNMjY2oSx1zpXQ+/
A4/js6At2ZqEUdCoTKpgVWpPRNeuJxZ3lHD9B8AEcLZqSWD3xdlW9SF7yJh1ufO1
JwD+9Sz4VqRLtr6uruCaox7XDmO0SftaEIn9Alcae64EKwbFLyyPScY4R4ND58ZM
//y/0iDQL9UIZd/cxktkDXuC96yyNbSbp18vdKrYpuQv92LF6Y3rJQ+cxZG0H/mN
tP4M97yOTst+DL0WF6x/rAnyaQ5hVwVQ2cDLH57JkSzQsIh4b2TWfTZ4tJ8ZQhU3
RxL85IG+KeNHQ+EKvr7z2JvvNU4e2viCPGkQkLeLyYI5kzMoORKguF8/kIJAQeov
ip5ekRtJqcaar5iBvpUb3GfDl0+rGahyn7A0/l8wU0NUDNN0+GzrwfbK3QUDGXAv
4EyfntcAifACistAts0lbRDYxuHk1qU5R6AIj4spJ4IyvqMKkUcna/rvDGGyvuby
NcCIoYSDzea34OKA2lEepNJcHjnXk8VeAGtysVgBlS8cAQOgLaMxNYQxWBqcPSRj
x3DGpQm1zZuwEuEUT3jAJR9KUOOJCtUJHVrrTctw4kQuCJ4pCOQ2JpQ/RxHE5T8T
N+007QM0MLg0HD0I65GyX7W/ZhxEVqn8j0ioL70voM7zkzXkO8gf5/J1p5xpUhVd
y6qGBumHXQRVgiuleH6JOmRQz85vX8QUkszZwOV+7VaL4LeFK6WTX+dynt7qr2BS
/NeW6982dh114XIyVrjvGPBbmkcJ3u63Xdh+AP57TqXrIqRkzd36C1dJlDbdQcbJ
UeWgRPVMss3a9erZU4KJ0jhOXxnXmu9j+9AOCbc3Qu7mVh5J8qJAztUO3bKo6t8O
uq+H1PG1EsNLiog7somsH4hYz2vavdIwiPjLPPQE0ecEZEmqMNE5aWSfAiYJnC0E
CgltMGlKo9CJjT4u5JQy+WJ4BFPmeTeFHGT3YULq+LiZKOOq9mr/I+WFqDYHgCmR
PhvHIhynrkeSbLbY7UAdYIncB5H5JzNiSHMCld5ltOk3cQbsE7MrzeDXkB0b3L3K
uXPJjhiTMBOSa9e9tBWBwK9fbfBRUDy32PGKYlHaY/cfiE02FSFMcxJFEjHrD2+9
LVuXM7LFFcKNwkKRHzpZvghQwm6/jsjgT1dPpJhTINMxmEuGruhHFGG8Z2Ho4F9U
QCqwSV/Vr+TLyzFYC4HKBA1qBU4V8V2byAKjV1ZSOy9LkkTLbX3oB2xO2EluSe+F
oy/9Ue8BcNE448ZHSxc36/C7EBulhw3J7mJqJ1Sa+jioEsEF3JGqjyiKD6mRWcGm
4yC2wEJpYrP+fS+B96BPzZmNSux8xKJEjHPDtUT5RdDwkZyzINxKPkvPy7Jrbg3G
ftpos/LGZ6v23+Nnr9vogmbOSQvuq3hOnAWiHe1RZJowHSclbmIrjhNDsxQVFWyi
Lv/45XjLHCP+w7lF5wSlXbOH6Do6ZGMlNLdcBfA7y8HePQHaLHLtK9mxO4eFZWzY
cxn9p9/tc5lREsT5pxECckf0EIAN1Z/MCgkG6/+dHGMwC+JL+H8YQxh9qMC/7gsZ
IZ0UePaFn0X10lXYqSLPIvcs5RKryoROIGZJPGkKl25TEkozhwmAd7QZ45SLRqI3
3R3oTBCsopXj0eCHpKatW7Keo3Zz9pd/Tkh5ES37QTOwVepqzP/+RmAA/9FU4YyD
KmCzm+dStl4grhO7Nuglv3J4H/95NlD8WM1MHqvUBJWpAwLVUxX5vUIi5STx7cm2
fHzRUbAS6wiIFAa3s4CSMOsifjQ6HudPLWfbo9t8Mb1zJWForBlVzzsY2X31vpUz
yIeEI+CUykIMyhx7XWHauZO3BTRfyLqBlKZ3VceQIH1pf3unogsZ3s/XfkmAnKWD
6JQLSTN3kkDTgPAk9Eir4VLVsFfbdK3HCj8DtBAL3iMynW9kv7G9jmneUlh5eXQX
YPT8OAj9f/7pb3OK1PbkAR2DFMXxhkRSmFpnYh1lI9627dG3nAa7I0vqJ673X8eE
QVNjHiy8QMuX8adNOb3lxNagcSDVPO6sBwNcKsmmfu3k34PbnHs9VWMqqbmq1R9z
4CuLqUZAVcTwi0LOuodHhOrAgynUdfwVzjvmYhCuY7kMETc0t0ca2FCogqjYD3So
wHuKuC3zgXprZg9fYuvTdGLoPXolNmrO2tlVhOyRpw0bwSTWec6ee0g4yW6Mq26w
umiiEzbQDA173ZOOakHcDdAiliqU8Jgynz5th+RCOFL98SoN+8wwjCJ7BBcI3Ut4
mdGZn7kI8vOaAHbPFsEmCF0GP7ABCJ3KNw5EoWCCI6NwOGBj/ZwFFYch0RtJybS/
F8rk74Ss2TXBkH1F6SOnZOB8SH5iBjXDyDAE2duvp3x3rcCJ3pjLF2dT+nvYEvW0
iQb/UAPBBzcT+sl/6qiyloP4IUjnTadJLBS7RbGqSLahCakaaTCwhGC3UW95CC/V
MbNFab9Lh/ybRsGYRpkWByKifPU0MzBtQr2htR8E2UJcRzCipdkpvO179gDqigFr
QJ/QuZ/q49sP6ZKqFadj0/twCNgsDoqc4Pzb9ZTu2IjqVcf8hUF4eSzI2qmiKceo
fIzaudTW5zg4DNY4Fa0kdWCirSfED42FIdEeyAB9HVI9PpUQFFEUndkcGSArBCU1
M/VgP+ieorjIcSzunO5rw+KZQKHolPWr2v3bA9BDDtly/+bTMKXwwkzXXjUCIAov
XHReXgkv3i4s4qFq7KyRvcRw5waxDqVphSudElxg4eYJcSI/8NR6l7E1VPZbYAbB
qarl/TuA750nm3Z8l8g8+NecfYGlS4bsknYIig7VtJgJVI/nAsj5URAzRQgcm94x
iljl8lfC1HEh/nzPFEPEJ9i1j/FpjhYr/y1KXR8eCKyiqP/K3QjJaoo7MEGT4STO
/Y9RhcQEk0ppimz3BljcWQsblqIBXm+yAV8p9hKjOp7d7ao+KRz6fktInI8KmNp7
nJmOIJxHVqwCgkkEwdBlH23eO56pQtvhp+pusyf0oYxIClKk0I2hWEI9RWHgcxih
cXSQ7ECwqQpiTVCAa00uo7+vkg4tdY+Fe8zkBhyJORoXS/9TLH6wa9cK0tk5fIu+
Nw0p32p9bGMBu9cpQfXFy3RCpj3R3+Xw8oDxJtL+7SNoy6HeR5EzkbMQLorVx6fw
blh+X5EKjr5+2u1pfNxIjRjcePoKv7AErFnKzQk3ZZ5dRY13FWpj3c7qBeRb3mfU
avmNpK4DwZjP9yu984Q3t3fp1vFCg+aa/ZFVFR2pn2jDsuPWDEzyfQe7KPj0szsz
cDAZL+Qzg48kTtZVCMnOrXY1k1lh/uQVtagF/WU5G9U8b2JdG26uRmYlzuCm6RWl
xNM3SgkLleVDMhq/GxbGnHXLi8P3d+AEbhKDbXF82YEbEG9k8DgXyuZZzvk93fX/
1FrX/wU3zK1O0Qus/+oDpAYynVrR4ZTR1AKHe2FxXL7rsJbjckrQtyMSRW6H0MHe
kfbsYIg7Q87/Vz7RwMbAQWWmTrs/JxFQdYqkvaj5Lq2jBmUz3nilOO/Ga+6E+6io
f/9JDnuq3NlDIZSRy3+wYS7fy80fzAZceEAvYbkEUrB7cx0qcEKxP7Vh6buU66Mf
o4LrumTd2VeXuGBD3oPJLBiFtdEl9foT8NRg4bJLqw3yZ2w5HfIy4WVEW3lFYZpl
0J5cIW5WeAHwkEPpqIpKL+8tdIE4p+PeYK5SXMLXIAd/MbaNyp8+ofKCKNEPQc6o
I15GlPRMSScfMEUH1gvRHDFpW4ZPsn7100zK5Eg5DErmpTa32Cy6iuhoJdtdAcbJ
E6Zz8U229nUOi2nNsCyr/DG9Er0SM+tmjBCfdZwwZp1f8sf/vW/KksuZcmCpOvf5
rMCfVVCCQFn4vhwpbBpkBgpxhpCU34lmlhkOxLZgZ0in1Wyg6sWNldKmlWvVyi6J
yEQssFWyYzsbwGImj3E6T7Dyx30aMleCjsYANAl1gtcspn7wuXp6HXRAqXtB/7qR
axPdFZqtgxl+X/x6eqzCe3geU4oLrJ8Jk65C3tMtU/70CH/byDeLqMm6GqOm3WBS
OXMAQigUk+xPILJ7T1eBzRlEC6S0JPN8dNimvYSjkaYH/Voaf0BCD4hOeqTxWvsE
dQReyqDpsFpLp2J3soVMFdWhFgPOgIaY/YsLN6OjvuOqlS1mVv8PwXCvubZyQxwp
VcSOdaUIexRAOPZajIocgAAkzsY08gIhpobl9y0qx1nDKTjVk/lBPayADy9M+HV1
DjgDSZDcwOytg7yCSl9BRpLT1vY0Cmn5/GzpEf5pLXu+l7ZH5aBfwvfL6MdhMS6Z
eAEWqaDqgh4j0G6Ip87WWTfVi/eJLL58FnKk7wgjiNymXicLN+QxBvwkAjgI+zxg
zzGmCyJWK9z0fMnDVf+6tpyFpKgx2/9nJUEFwsDSaEWCt4sDA9HL/cMkWyffy3/C
qn8KexsQMwpq+N17G70TV67bXm97CayviVr8CHg5Lh8sbhQ670BgpaKIQNlmo3Hb
lEvua3ptudznGMD78XDEPajk3tbrFuXCR6UeLD8owLrhCWzGl2tJSr2lA3VPG/P4
2GIoD9ByZWsdVnTDTLEI7PxNd3kMQjRIHO5ZC2hwzebKuEC8cvRMj7+/QZ00iL99
fYzA+FR09RhwOcsRMKqIlnP710Hi33QmuI7YGSIVA9gTAnqbYqIoepoWvdL0fFjE
SlKgy5VTHxI1xnovF73/0NB9sXdxYmUEItmqY5yqh4rvcB4MYOnvHK4iio1DLbgb
Y7Qg74fv5WlD2mlrlnmZO8Ev+7zecmBAjlPfkJmUbCmCpxnZGFrfZ/fKmIBrImpx
7wgMA7ZqGU69N/eFTvF789ZmR3f1dqu663BTIpK1T5xpQq5p8FYREJW91vPUN87p
dMvMTDaxCYZT6bUIQIekPLIUuGz38S8Zsfe09mFdl6BWHDemF0+2J1FDuKavU27x
CRjTcepa7qJf839GE4YK/98F69N1BiGxf8T00RYLYqjCErjtbcXGx+quH3gmCUbU
KEOgQJ3+dsQ9vdhOb861RRFaQQf0ij5UA0qlxsxs26WVI+VBWioIf42/HLVLI4Cz
uwo3ODa+8s3Y7r9Vgg2S/Scrw2VBnk4WQb5vMO49ze3dWTt6yhrFRXQzqcY27Z/L
iAFHvXzQeF9oLHFdqOapaCHUCAhXzOwk8FT1vi9SK4biykxMbYGSYBfIL4505MHL
xvCyLLTUcRUZInP9cp7ficYpD5174vdVECULMj+8T8biQEGt19scdySpKy9dXd8y
+ANnIElXYH+eyxQ95AG8o8Vy0CazL/lSJVtO9x/dWo+nzG3Gvz8LVXDTeHt8XWRj
cw33Ns25kD52MZdBkGpjHh5Y2yzMNW5seAiSCxMlwQDE2dHnzBQ7LrB/S8P4nqTS
fZaWEOmTfETxlQlDgzkuOgl0ZAeAxYfX7OcZnn5d7DBF7uJDIRQmXQikiPhjirau
LhRSupx9g95RPktCi2aLLidrcY5cx24K8eH/eJKSShSq7YKLNb1jSEC4RmR/wII9
mO8jpQg5tceDVuNpWUroxPvbf7/L4aHV5s3cB2e61LQHIihE1aR8wd+x0SwHlRt+
J3kn9K32Aj4TFZJaS3Zxb9MMIBcN2G7PGu58sG6yZXcPi0K604EsiHjRtMzoHBq7
Fb73nlSrDNVrLnFFdWxUIvSE4nP0hZWXbFayuJml+Shi7BoxOHgMPwWFNBRnQrpX
/lm3+5KHEBp0LzA4ALYKBOWFewCAYndLU+zFh8JdT1rBY6atjTQKuWubaNYk85zE
IpidjWOg84AxqbxvlPQMcHXPxevttRFTRuTbOyvXjtWLfJ6Y6Hm9JgWUTpYZPADK
97s4cfq5thAxJ6UFvagJki78nHtTS7gbUNXR21b2c5s+Aq/n9IO8f/OLta48QWeu
mKWaNGsb++6UT/U0w4Cu1fkBhTEdxBCWVL8EZrkozcNbtqMubOrGthXHy+xqrfIV
Py07phjm/B6ff/UuCZGlB+mnRyxnoq4HixRA69bZpf1TXXyceqU+OpJDXzgGVSRR
DGVmMQPS1biKFRcOaBzTX4xvm02CIjF27GhS6wSeggSPPPEMUkujyrkRTnwVAEvA
CC+uQiuRJCl2Ljuuob5E1BFIbQaJHxQ84YtHPQEU6TsTAoLeBzP84OBIjIK5+df8
XqOwdLr0jeZZYvUnyqxdBDV/uXCu3tZszswB1XQaP+PRkA4HAlSEXVeNanLttFjn
nQ/NrGXpOlVT45LLxNotYp/nV2a4r0/WGc1OpC68bUZ4bMAgCWtpHRrW0mPM358i
4D79//EYBpeH242pxdePNFjxm7J+POc7GyH8t+HEqRC1vWQET77XoDTJCfzisy3K
qj8z72CdTRsizIDQj5upc4Rl+o3ck6nB7+ubRUyreeqVuoZNpn9njW1DY+qTXdSN
Gsleh+ROloMCzxf2MtqeuAKkHdHBMa+IWhnyw18ykNgstM3xgpr3J2/wfboNRkpf
ewoHIig9LsbfWln2mSdwc7stKp3/c+6c1oonfVPKjEA+a/08KJcilztZHibSRf7U
dHfgdVTwPtCnlsZ1vw2xl6s3EtZ9SaDVkfNAGbslWDcX4udOFPqyO92foakadh9E
nnoJ8b2FuyBJ2QOJpTXuiJ1A3lMQcFu7CFCvMwFGCqBPkSMEAM+DgPjOIuFfslrL
u8M+h5cE3y83jZbgMUVO6ftjniGxx5MqE4BGwzNXr5bgr78JSqFx3TTtRHfDiJgg
h3o/MlB6AdZ0jsOHK0D9g18wqVfMPssEJAjCjyNFUo8AXbnXnXTWPIvCggMVtADo
hjPGl+rtai8L8EdUAE45ahVUquOPqqCGnPxKyMluVK3R6dGD7V59WamQlPFyPeFm
oIUdOSusXDcWC7t9BbA2rIR4jssOy0YTVh68HsTHeqh4I7+1JtSDlWITneaaMqxY
F98VVsn8I6fzdQPhhtD4NletW99W28tASkd6b0pvHchEpDWSpPusloZNd3pLgwkG
GcrgjGB3fXt+19m8Uqk/6XnZwDkyuKvaliNEmVPycq9g2OUgmZw8nIb4s6hEA2C2
sQ7ZlE6ivJhniv670XpKt3Wg0k3GHuHQTuj1rnNxyLHuZUfiFtN02ZdYyAZmgGXI
myt1YXOuiqALBiWVOUUNuRbm5kFHhoUlMvLxNEY8Pskmost7/p7/22s8LPo3GQfl
IGMKLcjOONMEtXN4erbi+Z4KphBLGUGqPtegdPdKxuk4p3jYEb7muyxpwxvi3fk0
I4FXwXHvyGNUm49VLcp3Hl0qK66rwqKSWokchHIP4Xf+bE7n+a1EK0onT6KQkug3
q8u9plRFee4t+l/5nL9CeP5TfSVtfNngflmkI/XDztya1eLjqEMIbOvpwhtGYUXI
Fez7+8X2Nmio2h5ltJXFmcznX9ejX9GWK3/bxXodufZsNj+jiCxn7QcRc9+Ua28D
TY/MHTkBTu8ima1GKIGGP+3Sx9nQyaq5WjC8Q31dYRExLMTrckVCcfdsbNPKzLBW
UdKhfzvV7Xd7bB5uvkrrN5J7SjpveiVuqfcyJP65OTGoYzrXBknpvFjsOgpazOiq
6hAUESoqCEfR+0VN8eyKDqX030poeF7oyj5tz8oZM53QL+1sM4H7FaIleL+7Ddbk
zxUEFu5t8jrXk64oXV8mnibZXCBJo4Xr1JXkkvMuRyN4E51WxuJm4d30/ff/Wuwg
P8vcxl1m+pjL8lsNK2AYJqGX71mV90IyJQ3wi4Aou1K3OJHhbqTmMFEAZmBYp84q
cSgF96a3kbdDloDlpgcFgtVRrT1Qp90OtJdZr549wMgBO7RlfM44992hbx9FT9hp
RamolC+w7gsgOwrChSZrd66a8CQ3I+lPSwKC5L0DkTwhx/dl4qalDoS9KSBPWfBH
X7bw6j7zsTghm0D/440MT8bT9KkHAMWS4am8V+ghrARkK/3bIY/4qE0r4nYRkxJk
zF4UGnHnxHLPmzVyBELaUWUF19YHNSH/DXY1VB/kU2+YAw+1QtGwHTaxyaYucZpV
Qw4riji+zXwdG41IuchTpf5cNBmtV1OwNXS6CBD2/k4xyA4ZvvzKvcMf41FJsVQp
d2O23djGvFATbhIjodaUlPsYwXZM/3WFgOXEWtog3grEB67H/XUJj0MhQJcHLKYC
5lxxNWGsXODOuHUZJGF2Sp9pjWjRMTkIwLtatIYkDmpGvZYY7ujrxErQV7D03N5P
vrUEUhFuPMB6hK7rcphSZ6iOYGSxXsgPG79NHvRon9U/QDn3yQSHKWLbFJQPwQ77
DJ9Q7PIGjpmNDzGHL8QZM7KAPDN2dtHAVlJ8x6QI9shr7x6N/vgFu8gCM8EGdLtb
d4aAmVgCpB3N4AWk+uEgfS+DCBz6hp/8p1EuR5WV3OGm2TJMvsCLHbPJ3493QiTV
eZzvtUhOnyx+5aMPRhZsWtplj5NS9YNOtmcrNso1i3YTBuw3nb/SicfsEXtlCm6i
3eOCin8tmP+sjF5ymSReyXKA35YZQs9gCrp06RZr+zv2VbRoYVgHvBZZr8tge0gb
k2ejmKXEJO2qpx1dhB8uPcYFX8muOWLwhB0KXWpvxs3mT3h4wmzgaXIvPWGXsRh+
yM3l00EShhZBkfQfc8M53SyzSGjGZRDketLqFfhF+T7D2TspnSV1qs01rWF1oAo5
Wv5JZRH6elBCdqV9XoQVfuNlMC/N4a4skbIc4KWyX2sZMaKT9FC1LxzgJUDBGbMI
t4i2vhMwCBzPApN1vHFdHTr0rz8k0GpFxomZvSWud3m/DdENrSHiWEfOrpVd4jqG
aGGqKkJ28oPfj0qpHfpcA7+kvTXn4z/eS9FWdRv6vof3I/+VtCeMHB2wuIY1NA+a
IXGhHc+1k2JLTSBkJ0Zr7YcYqCq8L1c/GtLyNxH9ypv7D2fvTbj6NPpUJifPU6B+
dOsa36paUd9aC1mCCroKcORdQ5zh7JePkC7kbG6PNAMLfyKQfrEPPb/GAzfL4yf1
5+iTifDoIcoy/TzEZ5N65GXZ1tc7IKMyRCxMdxPSOA89baShgC/2UEm1jQwy8+jk
Ps2ylncsdWPyEGK9VHBr4bpsx5bFHnhIPONMH4rwDSEJTrRaOuHt+yHSf8A94rPM
twIij/DaJob8OFW1PyRMGuZZZSR58naL9HxjzoAa5lCVlJY4NlMKZe5FhI4OTxNV
IxvjRaGfy+ergBzmWZ08YKyr0z8vTUCMKSoxUbZTMWi6c0PsDLZj5At6OhQWyWwz
msMhsKuIAWPjrb3KI50YHK9Cy8Aaz91JpjQgljgMffHkamdCcTnC3Q6q/A7Qaw2n
21ijgveZ2j8kThG35ydiyjsVfI7QfyGTwx9VhmSpPJy1cTX2bemLcQ2KrJn4RI11
IqtSbcvG0Yes18tN///Tn+mk86x+BOl/1XkgRQxvT9+s0klQgD0nutpoRkJvFFv4
W9bngBFmtEq2r+31yMqAX3zic02SfNlasCSW8JlAEq93CsIedbvTZ0n1JSEHsZ0v
jy+WulPJhPB/z8xNzHtmY6UhXnDdr7rg80DbqwsHHGTmIYxy6W0v1f4ieAmMjMFq
fGLGXQfZRjxEFV+AEmgiDGgbMoaVqzKw6QGtpV2gg5ZRq+3g0+OmaBl3zuCU6QOh
scLtUhCYF3ku/R2XOTF9HBLOWe2D4fhMZAt0Q3HLpzqxXPmDp3EX206mGDt4uC3y
evMsUQqFdQ9FBGAnsjdXlTX6DjOqpTf+epIq+vcBxHksuFwn0Gm2ZiGiR1cxzSOc
dk6xaFltFh9bYDKQlml7h7Qr4hFUptZ8LW7WseigSaD44zEFyjY+IZom9j1keUOY
7AXn15AAJVCISq/u2lgUzdWnCW4+qXfMwQLli44IUrcWbEIBqS9vWje6PZxH8odi
IG0iUOuzNJ39Mi/yCiGvmjxgKSPYzN+Z31aZ/cPD9u+AI4llObUwAM8/L9DH4Hde
MJmhc3X2bC130eLD9WDLD8d8/nXJgkFY9FZBhP/f9GnYdyXXCe6hOH5F5jt0+ZUO
xa/mw5iyX2XzOyeu5HSWNfQXL4aPicJIMbniLUJ24wZzFQHjVmPMqY+y+jpHZQxx
UswuiiQHS6PhyvQR0/buj/2X8PI2SV6UKSuzqElHAQ8kTDXQAxxjweQjwvqan2BB
R25eeBIDv4D+Y5KI8RdYxjuIrk6GTqPRAO1UuP+98Xrh/Bp4HKPvMnzCVtrNrIj+
VrSeerHy+cSD9i16ZCQTZwFf8he1XV8TTEFH/HSMWFdgR2Kccn5dpD40D0MoxhOu
DRK3+HKddTYnC//ZmC3ePOLPtpeKVvhLUyZfLhEOTzGKgHYbZvJlY5vMDk85KADe
clgJ1TxqBbJmI3r10HRk+se+ws8CHnJqoob3Ml8Y2ghNxQ8GoKc+OIEXA20evine
paA23Eo0G7W4xCfso3aRwLpBJgfTBgx9UyA1mNjzWKBWmgt/ubFFUpsrkb9ACCuk
PA+2kLlzuiWBZFMoIV864kEdzgfJX8C3pnSkgcIRcqHCWhvIsawwwVkX/5jhAi5G
KJC8rp9rsh0cCzvbt/RrpCTxuCmxfLCZWB8kCRVJ8SjtrwDmfpzRUWUH6vM4ZPo+
TfTs/4l0bcPqZMKsn3Cw8AP9kNmktTZWYoiSbR2FacfUp21CKMLqtTbSjHdQloai
NuhCxFng6DWNe+lRvI2VKEjtbJUEduUjtRBSEnuDrEvyu717/AVr9nLqDUx3bOj2
796ryOdP61+RW9rCK/WEHQSPdEvdV1E6yULe7QPaixArPohOKACbQP5nX70A+Ior
XkCycR5ylso5j3osN35hd8pdE3/e5zS5ahdMu9goZgat7VoZv2VSIJOYJnM5woyP
te0LJ+ROyQ43b0WtkeENmeWDtN9ZVp3VSZK/FE+O3QpcvI4dBfvN3qq7E7N9WngP
Wxsb6//lXnqou4D3ccFvWcmhc/BZziUWGBOx708PXDR4dG5Bm0VVxODdn5cJ5Krd
5KBTEAyvGfxC9B3dqRXO2QiXqAeBzJMV+QmBjAx6Vw22XncfMSRq2wyGwOU21ooK
zexJHuEKoFT0icVlPJOWgFmtWI+g+DJ0TapQyxgX6cIBYD3rNT2W492BbBVF6B6d
oljb15KXfQEe+gRf8NZvDuTHqPj4rog5zxoE0da2mKWfNCMjrXAK7o7GtWgTzleL
a1z2wojG0TSVpet9nI58Bl7ilYABk70tq4C1BrqZuTWllg3PJvLVKzx2lf168WUS
1ujuLVapGy4pdVdJurH5vKDYl6adW6iP4SZEE6HEJ6bbnvrLzuEIYDxMEmH0fNcJ
+9QkNJFCs7ddBzIfoFasLpj2o2YPviwYFFICwT2v92/KTypJQIki3Z+h12LtsJAU
oCz7kxCGYwbpPKAH4Ieu/L54bU6iQYUz5U78+NtW+HvDGlWfqBnB0ec1kMvVZH09
UtdVYUMKv+eayXLCvSY86zgML+gpffrh+NbT5wzzgO3P5cnAhqqbF9EtBv0egiJy
XDauvUs+hbPuuYQctJaG/kYsBW8VMAaNQQ12mdH2SR9o3ud3uBOF0aOQxPMHDDyu
dhZjyaLfLyWl+fJ6hwLJ6uRjCN5wMJIJM0JQ1roXfq3Tm7mL+8CSi+4B76otLbAy
o+26AIM6ewWIwoH28ZxNHD4l2Qa/L61LnaGvXQH5T0ADvk8fqQhB0y7u1qCO2k/r
FCScbrybNgiaLP8k+dkHD5W77yBlo7XRFH1tqfjERvyswvFsicpN8mKhVbIdNoMe
s91H+2ExuWOG28bw2bfDmWZ1Z7OouIaBMQGdwCQ9b/5xtOZhEBb2LnNNr/E575re
CbfmcfccCIpdnzYb/UL3ko2v8+4auyhVPN6XAUrxfdxQ3HdW4Q1aNtPjFQhG6gxQ
k/B21Cb4WxLDzNz4S/vblHqewFocFu9/GIziOeyDyZuhnIgOfROyTCnV3JVMeI1+
RkWkazNnrJ6c9gnUdjqwP9kgZkvUyePTQ5ecCJSYUrPORDh6GMxnC78UX+LpCq2A
3U/n/BrU75s17aeo4s0N6ijCuvJ108sgWI/IpnW+G9pZ/9FxwMdwoeqvwuGy9n11
AZGYLcZEPw34oEKLb/zTFmAk0f+2aH46pqY+rnXZ54CLhmEyI2Bl1VAOcY4KIRUy
nKs+Ln4EAbohl7Sjmtl5Jst0OeLuW+GODbMgqYyDhUbOGuAbnO+NLJbvWwDSbDPt
yNgwl4C6imeHi1wiI26gns9Qovy4hHS7TrPG9qcZ//4g7Y1ynlyLAsQMQQga00l7
u6JqjdntPQD7gfoOd5Cwh+TaI2Rge+tFwYvZvIin3BZPdk73c0oRJmO+SCCQaavU
Ui6/OfZN4XXvwh3sPY3bKhVar8wgmhQujlS6RWSYcWdMvdXT4Pzle78GXhzmTZrm
/4CKzB4CHn+jVVCzalFfyGIftCOr5DxPnz4lN340EO64uQWu9wf84E7JCcFau73p
fdLaQJBU2CwdPMJbL57bdfC1c/h49LJJdsoina9JXuM5xXgUSZ/nRLLDIfKhsif3
fsQdpML/fB85JYrlCGUZAUXgHN7WVMlZ3tpL/tXVrk9RJlneFYRFpkk36g7NxGPh
HmiFxB8fDxmxlwwvn2S1UWkSMJZLaakSAyundDnfbBB4/TBCvYlxsNPKbD4KWtik
XPySi+wRxero5M5oFEXU72a97d0HAdjktoyNiMmustKx81NBFep7iJvUIXQyhIB1
RnCh5C+tBBV5C1VjFzEQQ5PV20EF1EidrKth6oBMEYKcmFt4sNbCrh3OY5qbbdaP
K3TRjJZiWwjNiiI5clq6p9MT6djK0ryir9O2swKkgBAfIA/pbG9QvsShpJOe7w60
ixgUvf3VnmLOaS8Q8AueDORqDPrvIGTEuYpO3BkLNT5fS1x0Ln0obkt+qwFcUJn2
jfAGQ+kNtsqY1LADml2U4iqY6Qmus+AoQBFaT8TyJ9tlv1pjFmythkeb+dTSsopC
3sdvTsYNC6RnHsvS+efs0osn44m2MIwfn4caJ31srtn0vKksHVUuFXSklP6I4Qqr
y/ZUchs3YD+odeFvmLHaMW6hFdShKKZBKSfcacXUepJdi0C/oJPS0/LJCFZUIihX
E2Nn3QLpek0oqxL+WqCEB+MROkwwAMEWaCJEbOP/zSwPsvcb06mUQWbhKKpJDplJ
4uhKndTQ4skg3mlDPWGSqww/SMr3F2ItflJbsIo+mfBdsFCRgHJ30o3xiyflqvaB
DBEd6IWGAoPaVtKduxp6e4Twwxik8BXTrtbepQlVUU6nImlL8H4zcpBxcKj2mo3p
mfVMZRiV3Qz6AcntIvvM23dfaggJTUr/iEqjYg1wA98Y7LtqmJxgFkAk/JwvMTOK
2Aa2dUKEXY9fSsbswUDyWSnxnyVHjlW9pNai4dwdbLJ8wWSRqGJDL19R+yfCvbPc
Sp6oybb/O0K/9hFoDzyqZ6gXoRhmFcezBP8gzVbwFWUEq6ha6D8ueYVG0CYrntBo
1kbKWbsX/9fAIeKx0lIQL2X7AREuw8rAq+bapjYNxC/RQUWT33Ey82sUS2IUQ+AE
HlV2jH11M3C1um9mQyYDilMmC7Ib5H7X9gekdkd3zI7IedgnWYUpuEKd79UJiN2b
HPIHgo85VqXcCiB/g+6bgvgAvm2P7MqihTJuqt3nAvWZUiFi2ILnV/jRKUC9Kiio
Uw2KGBdGEVNoWxhzUUxl7r+Go3Wj6BoMHGmXjVKmCtPSFfO7EvVQjgbrYezZ1G56
azGA6OoPd3QabD+wSE5BuKC3XDmVBi+4oAlWeB0s4j0NlwGauxjq2W6SwOf0s0zb
y+WL9okfYIZelkegyQg+sRNS3RjzMXc2zmqmQHpf8R9FHyYy6ekEACiqkSTai1JR
vpO6rkIUhDeHZp/72uuBW0jFLs/xQOLFhmFaf38eXPRjiILZccprb8lNHkpxwPk+
4PCxVcw8vjpB13o13TnrtRtNoyBoMGXtHmcOjmb+zDcZ3m3bq9HYrYv11TcyrcXj
mW66JdRS3IfJAHb7js6TLVV9gO7Es6ZVTZx7cyhA3hCJLS8vu49nq+pYU3aRacMn
1PP2Jg435qPo9Syh4Of2yoCwOb0BmpF4HnKogZJFOPTZMN5U7bZcKdHFroTPMRjO
BOCEYbfXLoeLLeaaSBsPEQXwIQp5uSzIqz81GLaYNvMBR29Kd3wcGYRhZ+Xz/JKY
hHVSHrnSISq3CmW2tLqHV4nPj5szww405Hq3FFBaH16JofOtHrn00WmqKnbVA2l/
R1PdIHUb2Dtd9JwaJAVgtwtLhz8/6ij3zybFr8TLKmH58vnRyYyYZY7hqXb94WOU
o854rqkb/53dxOibpDcGHzkR9fSAvROLH4Xhtmuo8VH8XByUD2q3RKzjtagk1AuB
gdAGEZZWTJ3i1vqqcSrVECOrVOxf5IDruxtiWvL3DQngltrXyIzOUxO1diHuLqS6
6mDXLDXjici7uQnuRqmkyJspBYLsaEN7LgHaCgNI6uPaHNzEgVy/Vs9Ur2sN/jik
KIf1+M/YD3u1tQBq5zpu/6x9oaGMOylzYgIufG7D5ibm4Wyy/G2CISgHVcyOfGtU
EtvhaYefLCKzQLfJzyja411KXPbfBDp+gqpPLZ1FV1RXaQS7HIWlxY3xAJtNPvCH
L/beFHXFGnBPZdgio1KbUSdijJIeznrCgGL56JwWfZVTxEXJPM40m7+9MAmSgoRJ
LRz3xH3jsnH+SyAo9m/VlIQZZNPF/WTA3W/8kVMGOoG4GnmjI1Sa7A3foiXWyfHI
hcwLlFl8g5U7O13LUEl21t6y92rlAFzI9byc/g2GBd6Jh2O8gxf21F1NJXvzcOPh
DlmM0IMac62BKQD/NKcg493/BHy5OdTi6r7IF2DAVsDhMuC8QzWWdObfq42uVKX+
CsIYJa2rjgh+25fuCfyVWW6qv16TfN3/OHonhfIzU06PRP15szU+oYpkdRY0zGyp
HM+AO6Px1qDwS6UV0OJDmv/HAXcOGqz130JGY9ZvxDoVy4ILPHM8QXkdnnvzYRg2
df8x+v/rVLlHzpnRzx5JFToawQxG4GRYIQQVi6dGZniyHCk/h9cX1cDMkQo5bu5n
AZmVVoDUkQTp94bWFtugLNHtKG21OnquY5V141O4kYRXvzT0gfz8ZtWoEug3OBoG
6mr4wINlMabJ5tFLgvcLTclq6XySBQWBcTMmJusJyPyQYCrPPLEU+Awxl2Lb8rYP
IR/Jhfw997uhsuDVrTHE0Ri3AaYeCPMjDkwebmb2q+iG2F8yTYVPzP1SkbWsDqpL
9oBBl5IuG5TnZNmRwDMhNNWMjbpaGh6kmcPwqnmH4ooOud83WUjgM3IKfRvmmC6i
a2UyEPCess/C3S8lKqVtWfRA0uLq882qDtmdDK05gAuaLag9aUbK/8bEbXjBtqPq
mcJWcPfy9/yKVXt/j+LL50Xu7I1C4IZm5FUW95cSF+8miuJ4ATbg2Z4pswTJzC3V
qqdCnmFlHMRQP3NKKK0W7TCU1+Evy6g0iDUr1DHy5B3r/JvR35fVgB+w/T2ScmE7
NObOy/VXWg0rTSvQOrevm3hM4e7YqCoGtZJlWzyUAWhHk748/OPylXq3ffLz3K3U
V384novPDjP/oXCTNWkZ2Y3OGGhW9kVe0F0o5wWOoBTVKHJBO6HkOb11QHeCGudv
TmpYO+uka+Tdhg8rkXur7LNX5j5Kz15075l2DiHGb0flRVP/gOjpLdearSs+1iYi
fM10mxuaqYfBL6UAU0YlWIE76OW4a9UNEmS2X2N9t79GzedIvKi0iPWH/DiDOJou
wjn6/nYlA0je2TGWVJ5A3LAkUqPxTj1RgO5QnuGtNek+QGSTZOs0lo5gnGLjKmhK
DJNu67JCBhLhEoMUe/nq2GZz/EhPlOgevh5Di8G7jdNC1GmgUxEvaZXdDhV26wL7
SjxoBLaKcab+BUOI1zcNTceTDDaoR0H1nOQ6rCGsHsG9WXu7SCVb2YqTH2SliYJk
Q6JHvhp9Z/E++MSt0tHVLd63NatkCt3szAmjbiAithPYFTJ7ab5cdLf6PjnCOfeh
E5CA2YOEvYfyMGOxFGJhRb8krLB3GSVq5euE/+YWHSo27dWnOoRKGBma6cCJzcyB
V9/h1a0Lkus+S2cRv9ppORHovaxIsQ7uI+xCdvp4kGVyoBGtyJq/qXPwOcaGKcEI
sMXFUG3nnJJqVz1L+ZcilJqnZ8TAd6oTfmJXWH9bUuK4AzlBciahHMq8lOF7bRM+
asxwcVukTs7ptiWtTmGNYjYznaoTLKKxvuXgQ0CYN7VCAEwbQdbku2ZNO78IUQWw
Uw5G0cIOGa15VcTU+I5O33E7qK5u3I+YpmcOWn4yaskIw7KLyzGwfpE2Hd9m69hR
hJGM1T59oLBqvaMCCN9CA0b6R36K/v/X6XQaorjTuNmq40qkBFD1u6lJLcNjnBJa
/xTAvguXuuDGOaNlk5gXSiOevCgQ8ugoCjBtTfRoPaZvKzPNXYv85SkZkSRbEOSR
5dxD+bcltCxfmoZB4GWlkJaZ6UZ+RekQplh+pBd6EIbNDw9ugoR0IjBa9VviSXKr
MQ+75nR4kuQOCBPePMqiBGREtaSlZP++B4X5+vRy6GCroK6KMYtPPskeeK2qGQb2
UGA8yBGYPzkpz1y3gXo9HHyzdY0Zv++prnq2irVCkLjrt+JPHht5WfPri2Le4pAy
KHpn5FR9Pfpr26p9pzgFXvjv1//ZzxZPyKH/YvKyEJNX3wyNmRctYtX+Fl6AfWzO
Cg9fibQ8tvICpqfYifA/PCUgWZWLdnjia1l24cz6wL35Ge3pbik+4Oevvq12u7k7
Ing/kvTltKWk+Do6AqcbNSVn1BlrB0i0f0kXR7+LtNBa0mqUkmDCqiIQXcRO2HVX
dUdqHVfMJ56+B9WyjFJKeMxHUh3X8v7cRYv13H30r1GEZYWI+6wQoVUO4LxXA21p
Rjg3j3CGII5/55JpwqBDRK7gtIJ14iqxoRkUtZvwhdz1fUsg3AkoaK+8VD5Sk5CZ
4bITeiaNkUjJMktOtaJCwQCxdZ56f433LQ36yiFOA12KAS0GhR1lCEh9gCQbKx+D
v8k9g/LiFpWrbDMobOi6kVNTF8nXu8PUPscyfHptbR2n5awTzqUw6XA2pyUhTKLE
uygnNqYW0ozHSHndH51omNGOrabb+Vu+l49cT6U+rzsHE61Yee62pfwQgwysc7cp
G5elLwiy1+dXTxZMygsj2Vofy5n9GmV32QAuJ/+EkFl+Lv0efXi4ZFoWelkABxhw
aAwmi6c/gIJsf111eRIdedyxog5ohNPkhsi1SsJZVGev1Q1y9IoX2NC78KaQzMoQ
1n/Zirn5fX6q7gyvwulmUqqhYbQoI8JpRN79vBmkaWnPC8cNobtP+N/Hp82+qunD
v0kCPd4hUFbOuaWB3hUx8GWXoEJ5XilqvjLlWkOsFaD5vuN8inyBKtUMzBHFZKkY
yOE8RgMNfyDPkqVk10OKWwwmGX4beDxLow5Tkzv1KBsUPizbPIj+oNCkulOjADP9
Rpy/9XSR9N5q2andERI8k2iLuuvoDDHkdB1kErao7xIivJ6dGxP2U5y5jB7PDwGg
OHSuoLP5LkzC1JV/2EdICYjmmmwuk7E+i4ocslz5C9BbAUo4yorJ0uKHKE4eRjEU
FZiO1m8y5xOnHQr04kjq+B4dAuY4iZFM7DTmKYXz9N+yD40AyVI/tS4RZqIalG6A
tVAVu+eq+GSLhyYF5s7NPWOBQ1Qwqgw3BelZxKCchCc4ssq5LU84iXqX9qP1tGhe
rgbez0118ATOrNjigAj+pUbIYkxt1gdm3gK5YgkQ5f2AFlrdNfveNHsdfIUtc4qg
pof1YDmi4mQoj6Fo9pmr2evyQSBF7uZs5Wt6EabGyaDYDlvEr5/rHUUx09Kc66gZ
wiQllk8N1eX3EkNjJKc6gaSiZubYu1BJV1LehqG5ihfmkfog3yN5hTaUAkQhyzgt
13O1x1rapBAJpWAyARQQ9gVBjU4rIOsMgnTmVVQAB9LdriOdIYR8XbswbHqTMCs5
lXrFxIK2v2wHZr5ovDvfPMmPhuX8iC0fJeOAF7OHEoanzaNoA6ppJwWmesiwRXSv
7IZAy49Imz/wgMw7MZNZPd6+If0jVozCjL/hTnChHRSxAPwtkJjeT1FRpaykFjvV
c5vPNE+g9l0B3kLeLPtjjj1YkuleE2Ig5Sn3SkZ8oefvWFlPQKgTi51P8nyslPWH
SHqpF4xfvzn9VsF4YjFlermlO4Vm/d6KP49GTLHC8bfu2jExZWkpwMujDrbrLHV0
0xsJxmzaWgnDCPlX7GuzfkCmb1RAWtjjfs//KZyqjVvyZ1QHGTM3xFlyuWeMKQux
mbyKeNku2dVImmxw5dCySntMsLfrRsWS5J8EEfWw6sRmC997OJ5j4TMDkiyIjUwo
iYsikM/4DEqJ/l4fGgx/SLc5d5fU31Hr/Ds2r8BOuP8LdwyybpEem36z5uyVjXBS
/fdWehT7nXLitMaZKNTtrGPbaw2GJTQydZ+VGRkiQzTzAm78Erc+jLzIvl5BAHdF
EXQFeIwG7VCNbll8ITaSZT+U80vsSoepodPs+80ItxhtKSWdD4mJo+ucbZHFDw/J
RbBTQM3T8QYVnqPfuGx4VyAD++CyEAgdVcz1lkY4wKfJKmNaURx1R7S2nyz1d/Rp
IukblGPTQJ1Rsoa6Bbyqn9lzSNpJ0aXuwL3kCQtyFF8WHGUfsOfrj0yoGR/KIFxl
zZWAQXcQ7x5ebrLnM4P/MYA7PvvIKQaKCHSZvAPmUFaFgpZWiMkjbjkXC2hQS4VH
vbirORUQH6lviAjHzDKAw58TLQtAghmx2Qt9tbASxB/Do/60hDv4l6XRucO+eZ7H
aMtxKnnmgu45cM4NphdNxNdCJPjCuFwOdo9iUXGvKjhotGY+Fsv/JPfYcMrOBKl8
YvbkiYsg4DyBDgNH+n54HgJEeNm6n/PXUEIyD6EnmXLObfGZPAXb10dLhEw3K0nd
5hOhJR4PdjI3FOBrMGOUv89PK86nvJsXxImqWzE/tWXgVewgHDJXrSMFWyOSmBPb
Sqh1ixhc2e8aUY6Po8D/c+1AkV5x4xZ4kTdhM2KIdjn8FDknJyqwnpH9Q0j5kE/4
3PnLlaievPf6tApilYmnP+pfiXUvYgVKK31gL4fObnDVa+yxVX5KqMkHXItZnWfL
tbVev43o6DpWJoDs37MZWaj8Gb1lfQW5QGn/NyMt4SBRpT3Mo0hT8n4/FXzxn9uB
ZCGPO2UHVHJgVHpVtiyG1CTz0PloUgZPlE/ToRzw/Q6+7gUlNg+9nixvHdcrn16N
Fo/DRWV+wt0bI5PvyrELO3TA9OkGnB8CGFTAKyoDzTamR+iLgxMn3lO/eB35x9BA
zo1RNaDhNwJNxLOIFLexr2YvRmhZlzesDzXDpGLwq6CWMySgctY83A1AhbAbOU0P
y9AryJe0JxUdBJcIR5C26FhsPb4gJceY7BoRJ+mkwLaJY1eyP6o+NyssuJ7eCLzx
EfNrxcoTKA9ltYdK0f2xtpLVvOw/HJLA7t8KNFV07AMZhbItlwuKGfOTgJWEe6BV
BbvX8F4ehlHZWEETYjhognv9a270psbXsNqw2fppSSTPwL/fPpYEtgH8phwGAO9E
Tl5dawn1mBvEO2IgF6V9P1nJtivwnwPlZerConeqAUx+vIHBdRv4BTRSxT8YtDtH
EotytpPX2F0bfXemOAyIle655YyqxTHlkxYPkjZ6vnTCfjiNVqncSNn0HoLIsfcJ
y7BGCoE1J9aa5uvwRu1IBy9vozgxlEFqwPXZSkZhqjWJG4Jj8pUrjfF4y5mAI14s
VWN2xxwiJm6/dfYVSKYNPbi7HN5/O9CckkbTidJRdX5EIUPaWlbnLr/sZfdetWWA
TFNJcs44JlFFVYAhure9mfU/ELGbNHlni++SvwMkIWOwRDEm7KhuCP/U0V16ZSlV
lZW/VgumZy97OTDhBxirANyAPpRIwCYpH136P1gjhsMk+rQoxfuxWj/lTl0qXN+u
CBx2Rx0RbFIlAuwu8KfOjgsQGkluRn8d+8gho+9BjJf3R36XiNk+MrxprMO8n6/w
b3Znc+Yalm+sW+Ie+mqPK54A53pttqZJ01CzH49mxFQpRe8qBO/eMjbIMHleZXCb
fW4qPlGoGnlLDPUHxjmkO3oSq07Gxo1HSHqZWF2ognMnqDhwGNfkdRnmNnkN2GMN
LIdjl7b4DeQO7CawuT/DJpgRc+orJBS2vYrMKse0+0bPpcqsc3+p6Rd691Q1Bxv3
fw+OQKy3JxJtHB04cVAvgAmho7qBqP+U5zkGutDO1c1itVcL/ar6TDUmGqF03D2I
SIYnloie/ZSXf5fPy5IjM9CGvYZ+mEazMViyB8Y84mEzi2MquFTlf1dJObjeSXlt
Sh+nXDOgEFgh3//MuR3GGKGgaHJSCUOTAR2gfPtfoGYsMcFdTQT3pZpXOhbzBMlU
XyU7ZEUC7p7SLwuOhucCh/3O1FeCazKiV12/utwcmwp1wEKXZE03z+vZ9H1ba+x8
E0MXY9dW/+PP8BlwCipeN5K4WAUG7ASncre/JXB33jH3T/W3c8pcBQM4CTp+oCvV
tqhcNdNE/Ftf/vxhHgSu07ipkxY8TJqDNJ2lZIBuWGWxt/Q/lCzYdFxbgow9p15V
nXIOCZUfWwvPzarNTSBHzUBXj2ijIGGAzJKuebS6GA51/2mlfi33kprRfS2vnAcN
YedL56Ir1DS92J05wBSAia+SfeA6KsEcr7+yWQCHopMZg41JyCjhPhV4ttPo9zBl
mw5JKPEf3ptGOLn/W5nQEUnNEigcWyBDj7hb8HiKLJsnKM+ZAgedcrbzvGTJe5qc
Yyc6SGtrYp/e8cCigtWstvaS8YtZQSF4NuNzwqJ+KUC3Ljkbk5I+bt3f67bsm9nT
rOhtPnpFB9sRZRCECETr2+oHTrl+qsR8iB/A5HJOTqDSLcXYp9ErAc/aqwi28ulK
CjlTTTFImS/DssC3SwldzlNSh0mfQPuMsiJvUFHjuASV+YjjIzafO4MBNXW8Cz9G
hFbT/d/7R7cZmK8wbmYhLX7NsAz+42/V8WlLA7ikeG84CIfKNlf9ktMx51ey3f62
gzx6+UO4zOhWXdEdJIoTwhGFYjyKSBQEeoKaCbA3xCAHxYl+x9LZ9erDHBvOUaC7
nhyZohmWJjVxXZKCckmpvCxO9lxExOoHkK7ng1t8rS0SB+OdTXMzcsT5PbUD06RQ
+ew420vxDuFH7n8voUB9jWm5MTgzHdn/xzaf1B0+FVZFzYC3TLwRbRUMuIvryWyD
8/U/rKDI/15uBWbVeKjxgxOW7/szugRgq/NhZxo5TqpqXLXMpCdnAJxcnXNRBmT4
fFhhym4NFGBXwxGhtilkDKKPGJk3ChXPBQnntoQihtjGbqzRSuuDsfgwrYsf8mZs
lUMhcrF/b8aTHuXaNRlQDQJ06m24KTYZCkjPSZR3kILnHGWo3QSaBlY3DsbgH7Vb
d+02Cbn2/NdHwJ2zGGANyG/aR/bhnyxRPYMsCGpa4Z4swn3BDQ5FL1naykCo0mFZ
0i8tFj/Caue900t7AvdDFH+fwiRBAYbv1ol7m0twoJSR52lv9MFDzDAi6ptH8LKz
oNVNAxZgxuRrqoXAtKG8ZvZCYLdXRP+T/sC5ZwBFfAyRdvPmVqrbNTtC3/Bi4KEm
E2dLKjH4CnaYceq/wBmfS491QdHZJeknWaoBgbaC6Aj3qY98g7LUsexvnrsXGMTI
729VIenLRKPqdsT1m5d3z9+rf4zC6IEHQGN77/jozQpzr3gugmyMEuqsuIKgyN4q
Qd48Ta/wk3nx/oSVW8dxPzcG98n0ouNqkLMtwmcJSUNcO575Mp8s+kEhKExfWRu2
4L3fR/MR+q0fBv900Fh85E7x2WKvsSEBJ6UG0280RuOk0y7LsiPB5trIlw/+Vp+W
7sYh6wS8DxEfOOyWrd3bHlWsNHRywyVQKptaqjZKbfpco4eOrF78xQAaEAuEkFmj
HTufyuJkIZul3mVcmI6JFalTkM3q2/lq0Cu3CAzHXD7MJu8VRMdmDs2fgbeGhaY3
kuIlSTNzeXKFnYGEx0eOWORnvH0G2ASHsw7m5sg0s+bIn93JNmRuViXyRCSON9Zq
uSTrVqHwFR2U4wvru+77E9/ByxXuh2hTY2AdDhLCRb2CLRh2KS2QCTiRoSM4e4f0
ULtIPDKaH15ZIBLv/8treHzdp6aIIWOkARR+a0cGSQaZYttFedIk8BnHmMkpQUxj
/zXYKt4s00DNzvpqTM2tFJUWN7NMHqSDXkBtPKC108lX+TEb41typiDbGO4BeaVB
0aSON503/WyfR1+ZESzvP+YpLmjb41a/n2ogTZsNMUuTKQAVgjbahVX8P/voTdYN
1UJXsxsT+WnU083Vga+3sQ9cdoD80UnD/bASMqbIKHLzWi6+dfjgVugrKhVC2Quz
tODPF1N0slLVmREP/p9qOd7DWDQGKE/Z/7Ik6ah5GMz//pJocZ1GxJtsM217WGu3
j6yh+bKQ3VXmyS8QE+aErkWPYRaaP0WhaEUMHdQrHzSC+IG1viNh8P7HCpbnjjEW
LUb1cUSn6yp1WVHkbc+aMxfqyuYcq1uJcfONJKKx1+R4k//bkhYol9pyRFAl6Vcl
3RcROunPAG8rWA22YncsrZKvnIL4odqEcCE1DuHNMf9wqKSbJQTV2nPqMSQcai6A
/6SeqIjG9JA+cvHvrFYhXAYP2zuZCglEauLHNsyKDWb3sLbB/lK8PUc4J3hKs1bO
Q3l+r4a+s32WHwJTWSpL3f8Vg/k91nlCnu+Zm2bXDwHhx3RFmTpzCjlrj1ff0cuK
dHymP8FjJcqzRQ2AZoOZdbSrfhtAnmMBsN4S19t9ddCMiEUXrFYhyFL0eX9k9ogl
B5qtzKLKelbtcgCpxO8h01srNNtPJux7SgpMn0swIA5mBz929TQFf01yLJF4WMDO
bVsRecIAwQYTI4IQTySzACuJsT3V1GJlMu1MH9dmOE8dW5/CXSZ8UGnOarNTX6Db
CQLMU3mjOIs7jXsAFUyR/qHVPtbI3acLID5CcNsYD++ngJm2MrrJ7jE6QylGkA0G
MxcZzeTXCQ18oLF4VPXKJ2cbWDNIer0/3wV2fr/EOfsqM01ojdiLaobW5wSCtnY4
T5eoHbGIYuDuM++j9v5bfaV+Pd2bdxQgTLSk8HUiSgtIHQbc2MEzmYIgeqb8XJ8g
McbXynvE2M8Zn3P27QYYRUXaX0xzn1t9LKAcjER4rpZs/Hp4d0oIriBwS5Wo8xNf
zruG5RPbjgZ+AsQI4lqv0nShZlN6eykuG7oNvkIVfsR4h2+wAAt7A9rH97slhvfi
3Rt753kM8wtQFX+pfUYPufkAS6lAJatTiKw7dGJA6wRWKdOSgrwj5kzP7/UaYOwN
Nxcuh8zsB6RwLVaXLrNzMM7koimBUd0KnDUSn11Zu8kQXjaUNxuDzLeSPCF6XNVc
iJimJqLUW9tV3Mc8ZGwC7HrfLe1pWVHDgQGfdOPZIg3EWu9ZBRa8Cne/Bf7PK0JW
r1DBdOyY2uooTspxuOmUy+88Vem32L01QGpgTtiQRmDkIEJvCzGr67rnaWo5CHUJ
026zl0gFb/ZjMD50Rl4ladWrnZu7OqKQblIgbw8bXlZMZ+Drum0qXAFphI6z9KMJ
PvkSboZYNIU4rQ1KuMu2ecm9LOs1uDWQaReIf28t2Vq4fAGKtLWg6745G3iSX5+z
oFqQcafUMJpvRFGyB3FrxhpF9EAHl3XbkbjLvc7xIPEMMUgwrXadzE331XjzEtLm
VYx3RKZVy8kWr7qZoX250vRURnHU8zAsPprJFBDjQGhqmvgS+pQ070W0m8KjA97k
KKenQV4+LyJ3PpNejqsoXFgrv+Rhpdt0O/jhVmYGJbNsiHDX3JpTAcfiAjXwjIPO
3b2d2SqbbJ/al0wg54ReqgtGR7ylGKvVLLm7+Li7hX9Z2sBL3HwHqldGxA2sI1Xk
pDqVOq+l6KYGk4/juinhG/c6OgyTOqj3tvy2PlFCDWFnI8yj3IlwD2KNzz+TSR0W
MNIPicrmfv6FCvOc6hMYoYVKhKs1tLwHOrXpPYA6UmsdcE5A0Vfky4Sr/ScAzgU9
AYHAemEA8Nw5RKHkxDetxo5/ZtjCWNmUX+Z9SxgaZCJpB+ewgFnBdV57RDJ7PrXt
lB8aNmv/fGAbIzFWHdo/5Hb3scu01/nZM3LJq0TVrXZ3UgQewk62ZfvWJC34mLkn
DoaZZwnstV5bjmH3puXiGCGGxXwhx1OWAjSqcOcC2vxeks7RV25JsvrLN0EKMNL+
iweeFCkuNwNGF0pWn52erRYChtRg+WErz3V5O6nOyRBC90v8L54gkd0UflC8lhUn
9tqWOiTzuHTysmJ2/ysI3vakNrDAxAxI7nvK5GeHfkoR/xXnLF62u3yvs4ITwTcw
D4GmFv3Ze6d6K1TuTEc3T0hy3qXqKmh+zvG5x5SbjVF/Rft4UYbAMJmKseWi0VN3
7yHA8dPGKGmjmXql+qxYQUN/PlLlh5krvYAj21ui6KPBcm5xmYpfhin+GbYCmG3m
STnDXQYpITGHf9Hy/I5bQI5URM7MYT2Fxh3X74BoC1CaxdUYQxeJxa6RTZhIIDiA
qcGvDpLfa+ZGaAaQOPPr3plG6nk8kJJPj2baiQlGc1u3hl3nNk3T+mtXVZwcjhwX
6NTO+EG0zfvbqwNheFSHHczqUDOBKD+Cbl3/mChJ9l/PiGz9/uP8LvnabDDUV7ia
QZFWc97oGVzQwcoJLj+PBlT5npH38TduqmKsuM+azUSTYaDWan/9AVGHlKXx87Kb
G70+pYsQ4kwb+/4Zq1gNJ0e2M2OVPZnzGv3uNXVpr8bgVgkA1T1sEW1MCOSoymXD
TFGKlBH4XFVX3NeEVE2GQx7Hv97kxF/uJ0cXhc8kn0QA1rpvUCD9fpRt+K6VqfRg
g189mUhVHB4zgjnT93+v77obGIELhKs+jdgZq96aRtu+7XVbwb0q4U5opZlbcH70
sSP7VNtRaiEHrK3OS17FH+i+qWDi3SWAhDRfaI5DUC5ab7UU5qnYzIv0vsMSIQLn
rYX2iAzMvmcCu+xBwD9gq382RozuxOSQZoi2AUrd/ejC+7geb42kQCmVG5izQfn6
YmgOZQFY6ksKhq/ZeBJ1nK6eJFQmKROzECkGHGUNbAkBpEZYscbHl+FVXVm/Rhv/
VArZAlHladodC9ovmgP0Pa3Y5cZYwel7yCeqOjOILqdH9ImaFEuYMNPJ9AadlwL9
0ir7415zUZbt+DTUlAkNO684fDSYL1bc5v4agz/TSlEbO8vqGD9ybdWwpw1irXrB
83sbTqh050hlijbJ9PIZgvFNv0EXz0vDzMh6+DWrvkj3MxI4MbM/87X2sskyeXxS
NKgAEyXJC+iNl0eOA2MoLMB8ZzE8sBW675vPJIRwqkdedJ1YSYzh6T+blne+6qKu
lnyzvEnw8hj5dbVvqu3mAG48kMCNDN3Vwug+RP9HFd3m/c7/LAw7/u2EoAze6F05
03DirauPggTw86NwtQ76NHXj1ibG/ymRhcaARDoZlR3VemE0Tq9HhLNidUpXIhJQ
kXfBZ/iRzLZOMZJWmHDjtTNOO+FLaLEUoy3bL891JldGEZiFyFNot+Pq/6o6/ixx
qvtlegWhgZxxwAjomnJl6d11ob7/l237Eo55xvXqeuWXdh6bdBXOjievinZUcYGA
AIqhSd8A+lqjsbJnXe1Nfg82YzDQgsuHcNzwuE3d4ZPwIW6TXR5mvwTzKaXe/+af
paE/KdDMF1lLkQgBKAe2DAtC8evMOtazYqJRhB2Oqt9EedYAUXJJs8Omw4YScWuT
rOMNxPLkW5cB/+juWmL0WuYaRqt3gDqQtRoGIhaxfrXFh4qZogLXoXhnUKRxN2MJ
fQVOJoo0Eb3fnKhXQPudxGvwmDMD6oI/kiv/C764eALrsbCTTUEZyimzeJvzancl
wbe+4RYdVqG1mIEPxtWtSvlBMTD+eoKxjOLPtbFsOu9AgMPYlkWf7SUXaANHM/DA
kcaQfUxzPysXVVDFaqPWDf3O1VPGB+4XtdVZ4qZZiYe/vDiQbuonK3bpe15THupP
XzY2liG7gG+Ta3fQddohtFfxZPUgYbPYQ+GJjm+LmIXW+hSR+2WuIP4Nh3H0NJuv
xTw9Pr8VwT705RXtxF05pyETGUI29O4P2HKb2NIKbF7c6otY3/gEPRJaCmVpRt1M
f8N1yes0pJlLE8ohInuhKr6UofW+RZtO7LYMIQ8QgbfMdj18fhIF8k8Wb0xhtd/R
Ft+6dtCe8274IPPv05AbIJP4kgy2nPuc56tvuOiSwg9yfLwO3mihSoFHBDTqGcZf
xJA1d2kfG8NW72jtPrCUPn9NUTpQz8YyFhuXSg8l2G48QzUmtSP0suk4542vwi1p
9zkA3m5ISt9D7EuFxBHneynxF5o3uhB4u+aJ9RRmb34UoEyL9Jzgvr9UJt14eP6q
xmk/d4/PJ3Iq6OyDlO5pRw5MvmtAHBIiffIjpJJLVosyc2KLc8WeHXipEGQT5N7V
8TkNjkHHg4mIs97jcGCNsgFDYIZkrYI7aUtKkouskQQ0emKVyZKQ6OpfwRSVLQYa
aM9mEB9uTnVAh9c9l10wGMwsQBYNUSyysFLEDLvqcB8ThCK69lRPQmMniGAcd72L
lM6bdAu7Iaj70m4EDAsNJ3/egFlAnestJ8r90iELwqGHsiApNKYsLw5KKugSzt9F
u9FJsJxwKnKfgI6DJ4sc9dOiZDv2A73nWoEv89UxDoHCWyexfS76faZyGaXFApJn
8BC6mLldVFaiMmwo+rH4JTa89yDrz/f10Xy0fdwi3c0ETDcsb7oiXFweYzH8izK8
ArstndWHmBRfPN2188GcN7rcBsr4l7GFhfyNeuhgR1h+5YVatmxEELCNWfaeOG+B
eEUbafpp1U6AZ78dW67fMrOfizACfWJTvTPaoRF6NEE7zj7OgvXxzF8QtcrR+Bv8
1Zqce3POcrUeoAP2EckQkazgxp67yAKhvvhBrzpl5KzOVtGz0gV4+gKIVsNNoRQ9
jPMMSvIIZQMNwtPsSoA45h6p6nYpQ7bDIJEqUjFS3kuvnBgvBeuaY4dPW9N1w+VZ
CrQa/sQkovgvLRSy29+dpjCAWWs5r31R+vCzHBOqjFjlri8Gkjbwv3L/7VBblJOv
qABmuwOj4h//wLYLf2/+JiQT0OLyqBMWGhzr8jLR2DjbJKZQKAMurZcB3KEtsKrv
0JqLET9V0ReyR/yFypZDtS728y/+vEOJewdlQ5niCyqIvsPGPLLkuWO/2oywDmCe
NchlpspXiNv+pTu6wGGx0864lRArnF1zhlP/Agb+hH1VxQ7L6SkoJexMpO8w6Iz5
ealx5wOTA1SWVOcbexvumA35CXa7CURcQ2vhdofbe6MDzWF6Y/dwHFMIR1q+u+zk
OIJzKdAg3cxEJhQT295y+vw0muiE4GlKzQlLsr/yz48/kbJ+Fq3dDzRCDD1ZqsjR
9W76YNu5eDf/Wr1ErBP8bywsS11DWamY/RzSkI5YPKHOPm4AlKwSw4kJlDjPkYLZ
8GsgUIoagVOKdmYtfuVigOTGjLUevzVZlu13qh5OfZuqP+JmHm+3LTguZPJkDDol
ugg6abylGGzOPuIZmieHO95IKeDyJ9XzitgBvskmydiT4AaDfUzX47opjuI7/OG3
2rEQ3i7cWcXW7/ixFshAWbV5M0gVuwpgumhVRqRAJWNO8+MH1oJTl0qQNC4rNAZV
HeglXsB6EZSP3ucHGGFG/eMcI2L0W9wXfwv6kP/umVfB10v9yDmU7hvP1MsC0j4x
HFh6e/+Efn2NEvZFRLZUC5FfaQKzrG6eZw1Tua97bOyYy+rJG9m6HCHk45MnuRmB
CvUa2k0/DP3TEtrl5C7fHLPoGnPxMKKcwWphigLRDZsqMngQwaHXi5+CuZfJ4JJ0
yg4zrKfCrDb7OhGuoPKEpfGnwM9WGl+Stc7uHwgl0im3B5S/C8g31buDWlJrZ1ge
YVHPoKUbvPrxrAOX1VfhfaS9pM6vGR/NHDSKNr50bZHhklG6CzVi4ZV4hogeVjSG
M9xB53mnK8q5whcwisIOclHzZtZ+oSaW6wAdSyVTEbdICmUcwXOEEV5sPj65ELft
FFeHTrKmxULNkVkNEKQuHu20avwW02c/2ZuQcLaucrOuLT4ymwFc7rjJcWyy205S
lFsdzb/iZP0gmPy1C01E8onCAY98PgjupkcplrBxYrwuJRt002J4CpG0ainvCFfe
5YFRcgd8jEw2rA21dvk3iAzfNmiwhkzLQkE/cVjBSw+BqdjQTlhX7NTtPSPoVkIL
Epi1FiP9+vXm21svk+oL0qTVXXx94cAuHUZ+l+/eOWG2MWTsqONUxBUPjg8yWSAh
G9ooXbodQ4XeP/UY93CSsG00Jw2yiMbu5lQCvlyDcfZ1340+UStINaF5+94/Ifqv
0WfLi2TgNEXQuraeUti8teasuZaM5WQPTgKqrPSPaFl6RW7qOZDX6fRTHxVALFOp
MvRW/Q+ehf0MtXlv5hNin/b9vNt9Tu1LBR7elNQMr7X4qEG2sEpcgtUbFPG06iKL
tcbABm9pxdcZo4S7iiilVz4F7mb3qqomZpIjgp+lWJN3mQ6TYAP88KoTbFyd2vPQ
w5H9khocVtDZqnSMtTURA+omDkfXoxWMrPwBqDJtBH5JUz6GHSn1a7o55tUA4ZFM
U7fSs2hl+9Qo1Q7d3b4ECuIFJqBIIQx1evCQkHBzS5G90B/+cRe0euOSJthiWOoU
8u2d3JjYsNE3lKuUk7Jmr9QgY3XnlkSPAYyN7NGX/Q9PWIY6J4XBJNTQ8zB0H8BK
d8+TOSLW6ridnqqTkQd5UIku+Kouk6PqV8ZGBIxNy/Wm9EjIEIXHS9KTNqE6TNTG
4PjVMIHzCuuWTx9y2ckkLNGpA8rpTjoR1XacSfmzwdH0XS2F7LnGm8f2o3GlLCq+
TVn/sfyIKBzcQVBsIlplPiv5JmgLnPu5RbsnDR/wEGEve8o4E4dMzfFOPEX1GY34
KnpOUUUVJXSA2bSPJrAboqzN7/k2GHbSkLjtkCZtMt7fmR8XtxIXuOq39q4vcj3p
bPVtMlSTb35e89fmGyijl5MA+W2qNMAV6O0c1JdId73pkIuas86mBygk32uiRJHh
0TAbenBcDvEiYxMRk6cG1xdN1yDCaoJSmyJHm/Op/STVsqYXNnA+v3PobmGSRmSM
G9Yiw2UOtom0GS5ti8Cpjw+eZD5QdECm86NY0cCYsbAjmbZvJGrmKG3oK7UBRCIw
s/fHzhsanjb7qAZ0Oymj2hbfXzXcnTa3k/2nmhV6pv/An+ASSPrSfDnuXmhAOUg7
YjyfyFMD8AAzNOzV/IBXBh4tdXylFssakcjjofF6KaVwMezCYsZ6VyMPyXiyT3GI
cU6NW0ASsGPOMy5xIDQgcDEo05GRMNc7Yq0vM52cwh8dYtm3jylcK8sADp8kj/GK
+b03tSCADOntNr+AJH3GWDB2gKKAApMKHvY6t0rxOLe3GnCnCNvalHRXTeK6NyAg
b0/RoN+K6qk6XxV1vodwVeg6NFHL8Vc/aI5UKtB9hJHNem6OXvgG8WoUyU4pmbTH
nzj6uelOggJZR1bV1PzERzxEfnIqnyDjkNTjJWaePVWXV0fv/xz6ZyDDE5M2NRyx
IOWVqCtWBRkCtRnvPPmQ1pAVScAWYoou9m0k+MmVFDyarskyti3V6a1Fh2W6lmku
iWaJwT9/K4YDXsHCzD7qripkFPX9C9ch+AV6CYp6R3BbJV8sJkT5iCuqJcDQ3++v
HZYrod4NSAp5DizHXu2afVepotuGV23+PyDgjHwZLqxF/Pkq1+dttKQ4XfX7wEll
tMYHFWS51SUN0tfMwC3SUGCC/TmxXAM8phypS9sHMdgE+AKZ9JradgUIHsqjjB2Y
bF5GG1ZoPMDNCrSpwL5js6EXig6kwv2KNJGl7tHO+BTaiLgayqmT5EOOhb8XvKIw
i9SPZdToW5vNqQAirgGaaw979Dk09a7ErYdjxCywKPvf/0b1NqSqwQPtz8v6wbmI
+M8sKJ5WssAbmx3VUSvwn8K+pc/i4PIw8IwmWOVtMX3t1PkPY3xhzankyWAI/lFU
TsaRasXNf+BZZf2HvGOlR5wNFUUqziF8PskFAjqGdAaMkTOLn2abjQu1bm0xuKav
erhk7jt1WIN4xTp7EH/nNxYE+tDTRnq4fEEQenTEzTu2hOwwYce/9+0wnd/ELTvT
fG9n/8cE8SXtlo9Dz9bNh/jgHZX8xZYaTopiSwllzBmm3fF2CaW2avzHiU4DpPFx
XHanDBg3sfrUYBl2mdSMfImrIIrcue7C5fmOih5Wnvv0Y6CoBS2Mizxx/7zeME9C
jggsfrClOvQy4mcI6OMWV2KdF2UqnqzqJGfKmfyKQovMb3pCexEwCRe9mFFcKSKo
iS72uuNh7OtmCEKgoSkk0scPmmBmVHO3E5Gkz+ADtcNbdWlas3CeyGdNHEaMq3Ua
LKnbtV5DyG1RVrlJDnBJNc2jcrOxc91aP7PL3/uij9TpDZJox5B3baIMiTLd6n35
2sbU+edR8vcnuf6qHytk24+MjarCviFcj1Hpb/TSoCIVjYAH8SUP5aeyxE8Y5GPE
kO34OH2lOo1c4Xy/2CtZN3yyssiCNYkJPldJDtSqODk7Ff2MR+lVXqP9sW5Tsy44
jzIfs1yIObzB/nl5hyG+jrIizzuYqy4u9q0g26TlqsoR3jvtzM2DSrQDMhg4Y5qF
Hpz33QZsppIUS0LW6ZsRM3LyiHAvz+Ey0yezPPKXB/iTqxm9pcCyu4DnuXsnmb5h
K4mhEoSsCNKEWLVxwFAMGgb82uCX+T8iMKfxvOOCc/EQ7jVRWlpvSKMEFzEJyz4B
VAXPJH9187sm22m+PR/uJFuYQMa1oEytbtTCGFRWLpTOYr555D8DP0FOmYLX8k3h
HPOc0tjscW3VXrTEi3b/5f04hcb7zPqpyPN8F5ggQxM2S4/AlnOuzfn/xNHEUG2q
QFR7Tc9HE0de7bzrLPlMg3owHhyvQnLZ3lE0inGXNxjf12fRsA0RKx/rr2XUvtpY
hkad7aFIScNnxlGCSMbDuEwMAglgCr7dS4i9UHwqVf6NsICs9EuIoJoNtuAm/NtQ
f1qhbkDutSXSPEE2ATufehbs0LYeT12gZ+20rY1XtDmgluqWzIEhyAKRQrXA0TSz
dE8faSncvkH1nFmJ+N+9qW28/2nAlSh0jLnH9kjFGtWKsBFlFwSyR7gOVuujsbzI
enBRxAlh+DSy38/DnLx9E35MCBobD+1lmDE8vhgnkE2DC7e2C75NZDRaWfUZXStZ
fE3CuBzKVNC2OD104aMqXingfSLw6jnz6749mNRCClrdle1WbARJvEt2RhvsCEAA
/m1WvE9h/fxoc/V/mXtIWn3TUmmgZDZrbn4RGLZLzaeXhCh+y40YX4mR2uA81a0s
GZLWkC6zGtw54XJU9q7qet7inrJ2AlF4q7DEDXd1LFH2o1axXdj3Wd9uTNErsT0y
5c7Lsf6n+qo4+ubV+mmaOOwgu4YPDNq+U54sq782/xtEvzo8UNP2rmwedBRyyM6I
+qfj1RCb0hvfp8c4K/edM5nUyBIaQNPHel8tG+VgLKezqx8m7ybUWad7JbFA24py
d69CmtVGV4B5pcYfoOjgsT96OrqjGUaoKpQlVb33SkWGXzyKa+HyuumKyTHKoBRn
fAEHOuGpoD3cWXMQm/h2dti46N5bIrNuf5OPbuLwY+0BjBvGyRMsRghigOqCRtJ/
bHD7MfPa2iwHUjHb29Hci/LTVBtnc++g0MGE6RtGeBq0Ci4/NOXkgvlFPxTfRCom
IqXUb8uun4llZ6ZRgcLBIOD0S1tEV8SUax8k6XZOZivJEqFPTWKGZQvWKt4jPI9d
BXipHlVNsfnbhM4bbFUeRJOaN/YEk6tWXziAlzzMD0xnRL8l8zTuTe1OsmlGsEgS
flXR3+bTivtQSmUvItvQMtxC/Zcjj+WR0PBIMesb8sDHvbvb+fhrYPN30/e5MuSV
Lnt2eZmZzFZCVAGedngs8PtCfwF9xwRrOqg8OFh25LUxa+SVUATbC3rNYuz3b25w
JBRremSB2jMR1OOH/AibCeR9Jrbpgv0YVIdG1LQWrfbT1FMWxa2FIIqgvLzGfBYY
FdxvQByt0qX6gUVIb/He006HmyCD7mpthGRM0aFZYR7TxJuRwmehwkZytUHthQ60
tLWPTpUYxAU1y1wZ3YPRUlb0eE8ua68ZG5A/EqD+5Z5HSvsq3b2mvzs2LqUncLqI
2MkuGKUQTds2+33gu3r+f+nFAaOOtSJ4oZO0POGoxPtijSZc6mH7F+iFaGCJk1Yu
WYykw0pRiJg8OBTnuZXTEA7fXS5/w8hGGi241TriLKrhIP9RE7aa3O1VeJN2e88m
rfgh3XXmJFsnRMRTTodfMLepLDMWsKJROGoAB4ObETw+wANLj+egXpbCq5QZ36c0
9G8/Kn5QARfyx9Fy4MCcgI9XUNCiwZAJF2AU/BIABEB8wCFR/X9R7VPck9bKvapQ
VqB7lEouK1N9mjjCZ8eB2B8ycKHolrL7yCoRhKKcpxP91VzjVDVuomVklg4QL7FG
+0TZ69aGdrCI9oqGapJ5gIcNyhz0uvaAsXKXKzPxRz9i3WfXVHPrasgRHgKJmCLI
pbII0TwVuOVy4AlcuPSRvJTJf5hH9sRyF3lXrrHvY3aiO05AvM9jWXDSfOXfAN5u
ThU9iKC2AEyXpsyqeH3KSHvY5xJ2Z8Z4q6wB8huE6b0IzroDU5TYMR53/AiIu45g
LsKq9nhxXwMw0OH8iIkUf+RqTqiixVSl+07x83xaNEq2ODP17z6Z1QsGse+xQ/ju
ohM0mz6MMjkfBZL7XaqUK2WZL3vkWQIBvQEhIZ6e5uwRHXsKd62Dk0SykjTm4zMJ
PZRR6lmmNM7qyNVO+sVhM6cutWdBoy86XvToHxYH8UpI47PGnybAP5LQaXuLR/ed
TcDYEFaopl0EGZ4Go5wpf+2TFgbNF7rV+MEWz9+pX5ZmhDU6zya0TlZigAa0jfey
2zn0sxAGB4IOdy/V86am6sJij7zwatjUL3THPLPB6HhPCRNmy3ncS0+wOm21j9XZ
eUWOz/fmP/x3a8uYG6WYoBlF4aW/KHGKe6Y0L4yPNFOBkEtbAfJvtWnU4tTSzctR
sWi2Y474OX7uiyokB8epB8JxgT1BSvIYDu9Q2vFfxMyr/SgYGlTBjr74ISw9uiAS
1iuuOmR63yvyuyAQGPPsSyar7fW4U1SbqMsqniJiv+4IwCSewaznq4iqdu3mnjD3
kW7aNh7MhNxchTprv10R3s9H84rEW8TYxE+VbgoXwMc8FK/TKP4Ws4H+Ye9bQAYt
l9ZhMqt6ssrWIQ9J3Z3QNm1L1wd3QLBqy1BRwC+oK0YomV1BPGI73FknLRLag5nb
od9Ri/XOvnK71fMIvrl781D2iEnT5SZQlgSQ8kdw+AxJ4rol0NBxC/tBcFxjhgw/
arbTLiq+WNvUg3pwX9a5Z5Rb5WP/Z89lbzXjgs6UOIfVN25LDqMUu0gKQW8dGa+g
rUiz3UCgKL4/aoaTbKGpVvL3bVaR3slgYWjJnoXUKB7r4mB5JLpHfRvL3Md8awYh
hDsvXJsY067taVC8N4I3SS4dsRIIgdfmv6jHD4xljcQi3aYPMGogKal8p8QtL9ER
FcA4Ospzt+I7bE/VZ95C4j1FQKw0qrLEJYt9V/1qKdsBRrI8+bkotc7l1XTYBOfD
jPHp9C60PNpMGANCJ54BNxfUCQng325DoclvasCbmbjapKsu4527f+wlea6jJQvF
8rLwA15u8BL+6T8/xWNJNX1KqKmRffQkBy0TrFqeNx++o5MU9i6b+iIR2eP2FSq7
MzVaQT6oaPiXrTKuxEWNdeofrNM8u3TZa5iDL4OXSXoG1YakjOYQtr2Byr4QBKYC
EBThSn7Z5u+xshYw9yoHlZ+/zcwnKcrDTSqPwn+nBMK3xWA8pmwaqDfoPbyimX7c
aedtpo8uSgiqjF9pttOQk++35lWZAt7PaBRT2WCdmKCwCfyb4m3p9kBy6dQszXUy
rCrLERD2dQ7r3yEVCUwEeKij4f7PaCic2/Ogb7KTB0mmZeOMFcwpGzUTKUhHZqyv
jI2VcvK2iSpG5cVCCzsIgDXls4JGety6q1DHpKouXJsWd2RNNvvtl+q13ZAXEUmw
bIHJntHr93WaVV46yQ/8t6w/4p2rBcvkRVkwBJqB8LuWAbfsCo9qXxH40xJxq8wV
4n7ngY+1fnKmExqZwFf9GMEpxv6c+TLb/aI+Vls6k970z5nZ7UTnM7JUQq0wgGUy
tZt8qoCFAKj66uSYBadz3DMShWfVMGt40vzb9rTDF+x9hmVtcXzXaQbmN33YGw+p
SRrYuxI7espN7QBVkRb28yMRE05ChoamwHlukpoEM1oFbyu9Bkj4l1p1kfRcRQhz
FLSZ/oONJ92T5Uaga+T5VusIZVIJhVDTch8B20PqnL7WiwI2PHtVEKZDXIwvx7Np
x2HVAKN61bLPxospOQHx7h7QggOoJzHZWOguAswOTIotFe9nBoUf0ve3zaQm4wRm
8qtZlGkLR201egHoJj96hUrFKMvIc+ChgnT6CdKhVkcu529a/g7DmMT0c1avQAHB
9gVTSj3nMm3Xq+vXq9X+mh56i1NA/EOyEQ+jWloX3ndm7/K+x6+802YQEAz6uhC1
yKGdMN87AFydnxCkfFqLBYRcsAHOun89PTr0Yno25AQn9uvKlyUpxx2DNzuzPNFT
0Qy4/EkUYbuoITPFYiaXyggQJ7vptFwCNmkuPLmkw1aLN6hd1jWEdBCRY/izbFLH
YGbWS3x0+goz2yqvnH/cNaXoJ5gDhSDbX5xoIVAhP/7cqlKYoIFT+5qvbRipGihg
/OLThGU5Jgx3E3zU3MgShsCxtOnBw3faUAeVdKP5ab+mi1obvoWAOjhMEpr+wi3X
aC+Ro9b/Qagkcux6yfX98f85GhPYF3NSnnsQZkXOGldi2oDLMLXPc1SsQm7slmN2
RDV+Y0LLWiWyQP43y1s5uui8naWKGXAf8lzoPyIubfYOR6sXGrv/I99Qn2PjrMf6
Ub+iYm04/nwtVt6aD55VsEwND1c34PP+SICcGZjHSLv7cQhVlAjDsvSP0Q11ARo5
z8UYJFViTjRYy78QG/57OkLwcNKM6/buAW6cNgj8LikNJswT14csWEn20qFiJ6K1
BVQNgM9xDXw92e5Smzo5awy4QVVsb0Xr8tho7RrTxi9RqPRo3PuTSjPFOPaHadiU
beKb7jBVkPRRdUnqNQpEffZRrOlhqa7qfphVBFAxdMBu7MVOzAbPGRziYFGy7M05
t47zgBeuu0WW3rz52/ojiTDnxce1EjjrRabQ03CNADsI9UJXWYgHu0h9ajt/O6RG
1Bzb//kjnUUaxyFvGEjWOdOWRdk/XPdxZP6g2fzap/ixlzN6sIua4YkLMbK66tP9
f3HOF0y/nAEND6gAxhC1iNWlKDnnY+dpK9weSbvphkvqFk3M0oF0AM4fVUe15oAX
kiJpaXCSbuS7wqgk3xZ00EWgVN9yS0Pe976jD9uZqNrpK6HzMEejBvKyZuaOJzZa
ORfrgFvrByGkp+Yuls/sbNAWBvWevdYNt/KoQ/jC/HefwPME/LA4g/54rj3BAbXV
FpYrcaiTJyeT4EllaaL56c1SVECLGKWa4CR7QvhyRycACR+441Xxiwvqw4Ndj0si
UDe3cpMt295nhRHpqcvTLuc1nj/xnTYecwD3gokcYiyAgTWr0XYpZoeW57EtTMs9
+K+ehpSTO68bhuI5fmYCOG9SpGbnlVF09Z9wMPPnB2oj/bjbq3jGjAqzZAbuYMER
KigRO9mjCqN2n/KlYyN6Ya8vmt6bDOYIv0Qwuih1s9ASS1NM6o2CNW0LF5T58aGG
UR6lC5rlDk/254oWWM4CrQPWsCUmut2v25ta3J+6MXa5S7QXuMhCMClapVvBt/AD
tRkPJ2Nqk0NdQmZlI8IAofR98jnRlvgWA+nANByw+Aok+xhGX5VHbKk0trJ4PUCI
i+vOiMQwaIUBa2b5P0ZOVB4iBbkPPSyBFciHrA8M1lwN2TbUrawAd2GLT/vJQYRv
KBTm1vnhNiS6iJBS16xf0o5Pb47DqxwFzLtn3pg5bsRDI2Hhe/b3Urd/kKwrGlfW
LaDs3hTGasKYS+mm7O1kWQo/KphPmKYRIxHYzrPWlgAJlA8hYoNvd6xG4t8SiycB
kqYXOOQPNLd92fIRYPug9wp+13Z375ebGn08URbrlgelA69nbcvDP3jfwAWQQC15
yyrCtPVVUwIbdlnzr5MSwiXb0oBhvC9v+5JMEVmHWK3dMZV7WKNml2dDL+F8pGaK
aH5H9n2YdrF+g0FXby//hoSA3IDT8t8f/EEf38dVrKrQb+2na0skmaSdAcbOUqG3
AlEVDVwNgytlteJp1HoVl2nVpNrfDyhoHGOKd8sXvk0/jfifVcQ9zicW3WsADpoK
mMOLlh5i3Wvy4MAy2PZS21qVkWOL+azc78lf5gwBx8oQdKrsIhAwBOuTZNsF1cWm
N1vTewhbso5HQ8kJMOfd16Ml0FXyxV73ndUz2zziFVwxLLiZs1lOhJIEClUUguMP
kq3nvgsalYQ535NX64MpP4zbMLAn3uPGEnSPo9CsQTyymEQcoLK4vi7LUNw5UHnF
8gjnShWu9Mw4QT8UCzkLwojCLNITwgOAm0h0fVf91YeGczCq8gDgF18hjycXcSjs
892gY84utL7gCRZWYfWht/c/KtzXCl9n/ZDve4UhD9JkbDjgrdUs1RP2BqRfQc5B
nnamaT8tq32KfFggnWJpgx2rFGybpaqYZfbM+sK7nb7jXwYApMuyMvuAzNQwIZEf
fiCyR6FfpYdDge5ecgXU50vMcZl7giPQ6haz8ymMpFq3qEBNcZc4bYbWBiZnedIL
VM3UGuikeR4eEe2b/2eNJqtJZffjR+GL8wl1xIVDsUWTMgYnEjpT0CaHNH0rNwXy
noxdwF/UFUUGKiLn1PEH2hhR0CVzqvExVYhQJdfgfv33yJ79h6/PiqGJ3EuytIpv
jI4h82PtLHRPhTIAhFpwvv1Nkbq828eaWWwLZQiBRxzqCG2MUtrZ+0nTnDkJO9qP
p8jHHYRHl+/UWHw+pJChmouaaB42sFiin5f0WOSg27hWyrv7ZLLILm5CjFESAXJd
H6jpW6yoB3EGqcd8H8QO8Z9L48XGtH6f45+6X1TPqXCq0cog6rO6PbCpHyQ65+C3
awkLYeL1M/U3C5RRpzGBKUDgBZfh+rUxYP6Wtcujzn0dIsx0Oid4B+JZrTXjMRhk
KhWq1uDd0+Ho13PhvSgEzDP05JUVUnI74NUWvIDQisKarb5bcEYs65SwRIrozu3s
ddP9nXmYMTfwsFbfd0MEUWqy7/EEHAO0ELFhHHGfu3RD3jf6da43wk405GvePYFa
KnFAflrYHUPdSnADqH027szWaGhDmAYhuZDZD3L7fT8mPs4ATipptaqRa3JJA0jI
UfolZnDy+JePRmJOFJrYKFgGB3MvMtAocZhROtkGcIsQSvPsUMivZ0qTs1cQHQUJ
l3Yb9kQD3jB5CP+aIJq9iqR2CEO0YCgfs+In+o5zTxWKSiQi2WP3hYWR8wuvsFGs
BPikVETSEtUPJ8gijWc5zixjnCvtQXrb6NrTg+OrOWF9O3CYgYu8aggk4Y+XSgBC
N2yPcgbyscpTrY/gGCVFJmJZFlb26+VOkmahxZ9e7tkhoyaIZwVNmI2MFxHsCfU9
4/Ffmwn4a4pfjEUoK55VVtJKCqSdd35SstfWsgLwYiEaEn2VpGw1Sg+EwhX8yfDw
ON9znBzfLISbbAF3uFOYZAurYHV1mXTbo3W1X9rkDixAabe8TeC8EnFk0RvjF6DU
YIqJmSG1VJq72qww3Fsf9u4MkxXeJ0nwBCXucCmdznsJCYfiiuEgeMk1r/rVizZw
KAvxwJTdGgcVglsUfoQ9/X3Akxl/hbJkQp4eBzJL7pH9PtXqzyLJABghmi3Coca3
XLnfYUqXy+5bCCNvjuUj8xLdIFA/EsEwN7YKLgAVv1meowNzWYaz6rlIdfNfgnlc
DSYWgh9BNg7qTVSnS+rnFSrN2DmJqjb3jCpL/60hUYBiLiDLt71Irkm6XN5b+lvo
TDJAG4huZbza8UGzz657QceXvT63ENiptDNUSTtmPqYJVWtlYBDxT9bQtut0+f33
939kIzv7+hJMPmUQaSvw7ASKF5WeKFn6QKx7r2IxUXFPc2SOtaqcbM9YhkyDfVyQ
FD4QUi8jm6X2Eq8AjKush1wXwwYuxJQ1W9NNnnrdUaaFeZGcdH1SHbimduGJ1Qu5
vydZVpTydSgVoLHhlw2zL3zY7BG4mGktT8NSx/VW8LNHRwsogDbPjalvvh5AX6X4
GA6qUVwC+CWPYTBRDjaU3CKB3MSbkb2ZwoUylp5+YVFiMCgtNQl2iNRcJHBq+jya
3Uy2q4sDZqppW8fTDBeRWDluEL6IOAYgTU92vn66X2vCHx1ZGC7lGJnXBYUy9mBL
oa8rMxjl3KXmHH9IThjn9hZ/5VCvlS2bEEmqfhbkkjOVxgIsv9REJrvGbhebkvgt
lXKiqQbCB9Hh/+OpgCklTkAUDj167PwrHkG0P03B7fozA01mS+NxMy8HYTLsqICj
lLSuLyBQ31pdITLUQ8WsuW4fH0rIM409gV7V5/wof/pCriS550xk/QpyGhLyyLsC
dnYigIFjfKuRehlR9M7/6VLmuxXtAeGck85BINeZL05nEvbnadewAb824rY5hrCH
WqE6XY4kWXffGgzXX43qTnb32KNOjPAaxP2OF/ggHbr8SIYkJRT9rw+wTd9LyG0y
AUYLgBPkSKmutPZl4FcpOpNwsYQBBca8hh9mkhF2eg1wAWlhzpYJ7/Q0HYya+f9N
WYMljN07BcStg74I6FrDEX2Xuw5UaH9nUw8aP8RtmFV4W6RpPoEh5j3PKTuN8G2s
Amt9IEUy37vG9Pctz6kKf5EJUgD8zyYkVJt/Y9lHYBcmgS+pPDmww6jkDafEGOOL
PPv4XeN0FBGSBfwfSQD5NEHRYSqbqSJ3x7XngFYJebQlmy7eUZIcBnvM0Q1pPXDm
Ong/f4+Knu7MVh27h4qBLSVzUun9CaQLqz3EGhY2EyM=
`protect END_PROTECTED
