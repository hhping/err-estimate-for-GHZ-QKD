`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O6z4vdhwMb/sjrzcaydH9E6jMCynY8WnXj6tKf0V2WTKmemIN/NXKowKIUGM+mv8
Z2q2Tgpydd7AFRiaXuWGPXn+fFcgjs/BgHvEZ8+x0bHEnDt6E45n0T9OfTcWD8sS
p01WTgCAb3clfKmYpVjGYl0tGfuGP0lsr3YoVe178lBi7VVU4t3Hi/mlIf4Je90e
aoNQykrBIBLErDmW3hAKQjOPakxMbJMyfnYwU0KDKKJVjgmtdj1EpuJMh46w0auw
SPCuVGhH67qbRdnUDxTq/t7ySMzH0Y6vey89wuwM0oYkta9JcrbRHyJlCJVYcrLH
mmGjWgAqtKfVmJ+IjJJbxrx1TheJUi6uj0NXtbRmdmA=
`protect END_PROTECTED
