`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NMgQgu9JE+O8rEwaNlYm5TfMgE9VYGNmGiQAk7+z9cqxzSOK/2Lo2LO0mL7gv9DI
s2zQkISBQESyPozw2wL+OP8AU9ZYiqfulCLwiRbQwjR8E4jPHRzBMDpPeFe+Rao2
MyLfi6HMptAQ5deT8WtjPsAlwsXTRshhYPmGDJy6egLtEqhr4FdyPBqQ0JQI9ekw
QWnMvk5LiwkeWWOQIbxRyzRqQYCDJ5mVv4BYAlvCuEDXbCHN4NkGbZMTy5ygzpLb
ci5822c2ls/cvEgKQUa1NkUK4ox2SQ7LmveDBLnroFwkfVe07ymOcKN3f0tX9sZP
uN9vQlx90ui2ewckhsIjWqknw7hZeYRrGX/h4w1Em+9AdTn/Y3Vl16z2R383cChm
fazrPHbVZ3IZE08cA+0zyodyoyqtmGw2ImvLACHQldsJjL+gwfxs6iYgYgtQag5P
mybsCh67t10mU1icIKmZah0XF4tqK9SiXSxtAO6WgSRt5uoaDVE4/ZvV+HclVMo2
`protect END_PROTECTED
