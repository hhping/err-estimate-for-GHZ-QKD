`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1yLnfjHfO3kUx+61AP2wJxua30/6U0nHUUHtGwGy7zGWxyWDjT/v5zVq3p5+UIRl
u5hFIISeb7S7lv4gIuiuCy5qPWCMV5I4zmSOMIkpk7QhVN2F2RAAhs5biA7OBzwc
HykZLSfBgQ5nSBy/EMLye6MSS7GJhs95E6wy7YpAPc/YeJs8d5gkIJ1OHOEEjzjN
xaV5WhKgLsRmetGG4jCoyYi2XRHvWP36SE4xCCClaKXcctKCd2Np1Zt3frmOb0XW
gOyH0EbMMLGd8PDG21xwFfslpfb63LP77N06gO2buEnwm3YTGDkhHYPe+29FJLGc
ZGheKTLB/eSTfywq9Z8J6W6Otx7+Ar1/8QPoCSDMZdx253TGwg3tufhR/6KCBHkn
exISAxcXj7OjrI1pJ6B2MggTBlDeakFl1q56Wcbbixh4k6IQadaRZg4Wz+nYjfzg
lMlvIwU0U7pj52Wisgqrb2yy5wNKcspuSUXrC9BCrXYm3vSPCW+lB3kx3pOgEroU
zEHcOoLFSkRQ3pWbEBuLL5y3itp9pV+qWGdVTpsEbO3nEniCpHXDk55uLrUxu9wb
BAuyKO7hf0tIgNyA98h1ME5aW2gIoobtr2WuoIDDm+MWhothHuqWjw7J1QiD40Fp
ZhJ8WrIOnkWpEDtdVN3VFEITQNSikL9jVMxcY63ZebccPgGBSy6trIaK9+5DKNaP
ic4fYVbx9Pp4r7mmbpJajSNSTLBJihdJ8xNJyYvhuSCP4qPJpSDv7qvzVbu3Ipxq
rKr8h4MANiwq/SHieXvY99LVe08g2Up3eY4PymIOMlS2+i7p1esbX8/YbvFUS3oO
jh7X7Ts07UvmM214/cpviHeapWgeSqIXCMgYkBSPDPISBGyVDVM2dbJrQQnvBjL2
cNa7JlanSeQdMXlSQnScRduKfOqNpS1sk4nmzDP/a6T6/4OI+ayHrqOxXmN5zDDU
LT2woZOO40nalGPernODsYaX+AHjBG9wIfN57mGbSn4jV/zq4psMoOn4oM0BytFE
wv2rJVHK5FIazpTXAa3D6WW1szWg3OFFI3ocxwiVa8tS6yGeVxRsHoRoeZ+G5T83
ciu9lwR0mjSBebmpU81aTMrhOIeaoYa5scI4PsEeYGwn671LDYy3YP6gQYIN76YE
8dnS4lUjcGQE4ySjZOcCHg==
`protect END_PROTECTED
