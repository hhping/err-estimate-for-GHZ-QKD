`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h5WYPAphcfqs9srw21KLAfe05YGnFfbHUOeCrWpJC1V54OrG6E55+8KILRnF3sJE
TuWAr8Nx2m9jfGa8bQOvt7zAkyWQ3ApQSvp596oh9UFi0NWD16AfeQEbb1UfpiP4
De2/Ui2TI3GNjwLXrU9VKIRc/nCpvj/bqNNQuki239eKboiVZkQgN4c/Pg9LmURe
MI5BFd9fuSX6ykiqMXXxK5vD1g8qzqM1slwvaort9Q8so+s4dSaAh5H/suP6gEbp
EGZqrcWKJFhQTyZrNCdL6Fsz3xbwpkZSGGhy3dzCooOKAPKJY2h4bPON1UaJbJ7V
LWUN0V7ccq6qZ7X+b11sUdf3z4kk25ybOSKfVymXgC3pjPysA8UJKt38R02pVK2y
FEIC9bJtYcZdxJgnrvM7lF5SogmWHFPBLLqrqqejmLXosq3NVMd0bLN7REWrfDYq
bJld+y+IdH3NrYVENg+XKxJFlGLfnY4nOZV1Q04suT96EoGE0ySmwFr5Ap0J+mNq
31dZonO4ut2EkSJU51XgI4dbyag+TDsv3vcTf/Mmx0Pv82S+iBY4hl1vrMZg1HVn
4g7hjcj4VKkepEfNXnrRTztGmRzWTmAc8tFP6pydhf0lE64vP7yxYcHjR3KEFj91
tHHdeUIRfQB3WxG+eJzMqXOr4hU40RNoH/hkE3qDW6wxU11w0VdM83A1pAZVak3G
c5X2AnrZ6XczMTOqfBiT5q8FP2Cu6x0Hz5/OzgNm6hH2w9nDCqsEmcT+Hv5Ldn7Q
qNmS4kxPepYQXdtXB6JyIYf1qzHZy1UwOre6H/9BuXiy2EcJdjCeJ7bPH1nX4Cyc
yl4f5LvOEWuo8JSv1jT6cGrfNFPSrxPAi6bBwL5dc610kNJtNrhBNWDapp7H7nc+
PbW9aFA69oDDF21f1DPCaqhx3md106evY+AvO+KlRkrAPts8ymhwvKStySBbPtNx
3TgeeFot711rq7aAwLwI0B6Ku/Jns+5sL4VF0srkNeFQKaqwUZqgURl+LviOhCWg
94ilwhwbiACvgdNsJSMu9IxNU02GS0by0XWCY6ABXzRSnogPBVha/4C5Cm1EH1Ae
2vytX/ZYcgY2RmJZRE/xCI+mDSZVAk7JOr2Wqfut5ySOkdDXQYN53a2YwUh44iV3
cO5HqWpSccYduAM/mHljNIed/dTaxmi684rbT8XtR8FYTdQfPz3vUNeX8tljHTy9
dTVbjHmtPnSPNtsf8SMFQ81hQwjoLY/nJ4HSXKvwMvnrPU+wpals5XDzjrKUB4zQ
uu4lKY7GR0OI8K0TSCznPGSy6HsM449fTZABmgMFYvaWfs0k4RsEht4k899iI/dd
tpbbT1px/LF6Xgcd2LvP8kieMpPVb6z/D0UXpeA4cSr71nQUjIjwKQGlQ0TSAjb3
ERfWf3cIOzzgXlugXC3GO12ebFqXhox5056qpFMQuXZpfL9frtWECn7d8z6L5t6D
jGRRSQc0NmgUOXLGqgfjyma2tC421Ds/6t2DJ8RM95fKc0D5TP/SI97mMBr1ej0K
sr0cxvdQPL3bwAtrKXPMpiL8bQt0rGnMaZzQx92azZh6X1tZAZAJqYdrL59VDSfd
m3W8GaX7fnpUxue/5f38ZSo+SxIXTBAtfATpPXCLamAcYp7UzM0YD0U+J/3TEapw
NpOkV/mz5kmvD3oAPK16esapMgu5+p0vZR7zn8XV2Gc9mZzS9aRMboM0Xhyung3m
P7syQnwlvtUaaUP2TZ4ItD4oOHqHnzPRj/6po0mfE/TIkTyBoTGqs1Q3gfaMYoO5
xGxBKCxoib3pPS1bbaerTTzgJgusADVKzCEuu4kW9XSW0IsW6QrIDVEmf56S5/DU
kiDQYSqTshoQo9A2zmZ38IvI4upRWak1zUvSjUwSf30rHNr2YiqQx1J0InqEXbJI
pjM8qE7UUo8UVSUA81x3ZvbYIYVzM2nC1rBQjW19cLRBb1/MsII7PbGeApNkt4R4
isWaCnupFqKAg65L3GTPKekN5KL0i8GWUugNBs1JxOiaxrBrLwpg3ARvgVYAJSpC
cZUfWG2Wt4GLOL6SrQ9SgoJsaa2v9BCVrIlDogrAjTRzwVmey73TuwcpVC8LIvO0
a17B6//eqqShcyfVeAkELqeZmvNFG9vanp6dc97Hfj9XXMVAcHwzLqMqDqfzHONi
LT8dSCf+RFSxML8cbBxx8RpjJQ8QPtt+V5EziOCXu/t34uT03psAiD76IzNijHZG
ZpgHNH2g5gOejYasQ76J5PyxQkw3xdS4HR0yv0/pOYjRvme5hhDWZi7sMXTpaOjD
+86fbaa+gFHNteUBIVJPJrJ3aczMKpKnPWMhhrTD3KPV8Mxt3jNU1hoNXg8JzT83
++7dClh5gEIhKwWwBgvl/+2c/b6yWestTQKw5rcna/AqSVQcrm9KD2tO5kNvgGKK
woYwvT1lYNRdU5XMx0z8Z+QI0gCOGNfbx1JYRox61MypgLnjltS4FAm5l0SVLRrl
EI9goK3Ug7tbOcPrUNbozRWQAR/tpdAaYmbiMdwW9ZQzELR3FLDwG6ftpjjEAiCT
LXUjpCKqa1MY1ZSetJvCsutwH8O8YEYFSPCX2H4EK5y7y8DzysrvZNV7FSnXjfyk
CYPyd9F0yMatzfFTOJwU7Bz2x8uSEK91hkDsGE30/qTxdWj4dcEnXsiOe0GkbWN+
js942uwRfUoRhXTzUtMVL5AzulXmgbAgCaEuB2NdH13qBS66TTpdu4tp15Qi+13n
E50kxbwwWTy3jRf4U6UeRWwVyR+wouFLtEgDwBkgetCyvNflPH19W/xPhQMVbQlI
BZaIokqWXeKN9Rspmnb8cWgnH0XeG4Ln15pTFBzkQ6FeE3rgYEqOKy+G4fQDmEfv
VCmyXJUQPvwbJSGJqpxqxGGDtCmaXVAsivEnxtUwNwA0yxfWi8Iei0ekcXPlQer2
g3mmuySpMCK/IfFrzW4ymxD6X60oeRRHDYsZU9SmG0NzqpoZzlDqAtOcjCfiJfCv
ORtrwDWszIwIOSfeVRNDO568lKF4jRhRYME4faSQW5LRMu70ZyD7lMMGgwUx3WG3
ayI06sro9wyF9BEKnavAw2BGOJuUYO0v9v3P0er0cZRcOiB49baWRB1AXLLohLft
29W0tJ5fTYmH8evxLwjlw1wGm10dIw1U1drya024t0uvYCwUaZt7xAz9/zj78UgM
BnklVye3k6jhyYIZG+qTmuJyHKoUzwYP7IkOmBI8tjRVB2tztoZGhNApYdcgS72d
6POAoeGvTMMu3XnNYMOC2g+ogiRZwxDobQiKd1ehPunFGFNhI4QSNVMwMTQNKuZj
VX2Q2EfaP0dZYpnZkD6SIIuMRb3QHMPOiDPBMaLl9RvTuERngnoutC4rodJzHRjE
/hqO3bjItSEkjGRPeFVkajAQOYmglHxX7/xY/Wl9JMzrU1UsQUB9p7/WujMwY1QH
TBBATj+7weVHab5K0K27zLoc42I0fzYA0BC7+dFr1nsebjhkRqMqxJSgJ5CCI7H8
ooJGhJsDEZYNE8klmpRg6e+V9AqhTEkrbibCqnauVnU5bblNyqrSlW1KPL7vFjbL
BXjjPUygoetcs1hELeCeL/g16oCNKPxTM0r87kkyWC/fT/qcNZ+JiH8rPWJJPSQI
Ua4MvqeVLovqWTJEVyc7mpaVdnFJ/sbr0uJZJt2TK4ag6k7gfVbZ0gDzoGpXd0+8
Oq0Ns2kuMb79cyOolZqkCVFYl60d9tcWgveh16yWNn9k5I9Abt2x+WzwXW5FDXaX
Q17j8MG1C5nI3MqUQNRcIly86SAG3gYtXg6czCBIle0ZqqJe+4B/EF6L17A/bbW+
0NQaoLqqUj2rVhz4oClBUMuzwPCUi3SOmYfuIQbka1UbipM6VepCz7wWnXMGdlQ+
U7G7R+2i52ne8kamNKiJook0PT+Bb3bfVxoh2IGRbF165WPM9OKn8ANgmTBJ8453
OO7O3mFyFDVW84++Y74i+VGanE7w1SlMLIJKpeEU+Ng8+uLtcZieOE7nz2nhbT2z
rpBTWxUQLs1bSdAHUvzDIDyZvt2Y7OHY1+HNpRr/tn6Ww+fnkHtmgKo8gky2723q
WSnyhWyCAb9i7IJSee+CJSsIJDu7IwQYMPqPEVIOQ0ayE1UqA/pWQKjWCTZseUXs
R/AYbZOXG0uHW0oCjaSrzGuE087hRJOHtjKC8q5vDNONZojOtTpYsIIZQfR8PTf7
eKpjWQF4sCd5RQ7nL2mapXGcoP/PugpTh8FZ7wn6YZCsXcSZsCot20eb+cQtvZE5
WbZfQuihnHENecAtwK5xEK+KXV8vQgJCdiGy1oRuhAUTW0bwnXqZkyXSYFwZCb7m
OgHjv2B0gdu9XOGG6kNsuEVJNfFimqGPAe+q84fUWPvt4Yu/SLQU4cJnePc6swJ+
eXB9sf8Z/FYDaVrinpGnKG1j7xPafuvkOOIAD7iR2C0=
`protect END_PROTECTED
