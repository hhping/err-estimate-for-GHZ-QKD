`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M0Gbqlu6LIidGHthL4hbX3clLl5x+mdTbxUoN1/9sRp0Ewd2ABwIMoqkjE9eDx3C
XxWoiDTC8GUuCMAIQJ45XwIN5YJg9v+R5GYJ421AM/WwE6FEkg2VREvOISA+eZbm
bJmHB3hXc3UxnbCp/bhYvL+Kui64gerKC27W01P/aY17hm9TGITD8UoAdqHdRoFZ
iCNcsZP9hj9M2utMjAnRjHySM5lMcIYzi0lgtesZAXXSMV+SUFCfPtSa+QVcaecX
vLfWlI6oOPLvFdktV/fDo5WSmpgRbO/cEu8cZzTQRWju+s3UCdLyo0N9An0ngoSQ
4YNHXZWQyGg7mSFEqYqtYaYPihGE7j/VHKM85MPqFFE8KVxVKtYaCgpyrZlUQGR8
jRwKstP08K4Pvhz0Az1uO8HxHedz3ZW8+cBYeHQ13CWSdu639IqgxQfvIoBE1g74
bZEh04rC+zH5xrGW9gh7+/DxSMkF/IIX5EVsFK15A5cjlD6boNgP9wHgRlmr9yNf
aVFu3j7csmpfWchLK2LYc1BE51BPWhH9Pvekpb9ClsWqjSCltnSnFjte15VTqQfk
vujJD0YJpuFnqc8bsNygYOvJKLHTNrUWJ8IFDadZcNH1NXFfHnm5o6ZGPOEYLx//
w+Ddelgaq3wZ4zcVcWXrRW45mQXg+dEaNsKJzVqSfut+P5vq5mRLIijM/QsxeY66
nIiflOqAeRsTdS6D1Mmfcmul4d6CkCHd8IdH92PD/jzG7Wfs+1WRNR33vVw0jJd7
9UA2AhNZlHzuMpgDmOEoZV4rInXRCAy2edAdwFzXMe5qP7/rl7DpPUXiCdcxctbB
psK/p45ACCOpfmwXKv/OE+HYrsNIvRRpIC16M/J5bgj+cbhOrFj4jh2G2AZlbBub
BqdmufNLt3bOFo/rrLiuhcN4yDehtd/q8gv57JGuhUymymz1xGjusIQEDORAVu5k
zW7dWP/0CxjBs+d14Ik9eJ+cAjEGQZloPa8LFgoQkPisE9k1jdNjUXExdGum8RCE
GdBpmkBL8/TJWOnmdheOUkSRnGeJv35qg3ak0w96ZrZJltkOcSnSfuE79rz5G8dK
vNmXdj5Z9fPV5mHzmtD6malCXnZ991MnmCVDQ4W3u0zIOeZkQ0gsy8POo92aGcI4
wB1lo8aFvy74aCVfWJ8DyxPDvWQDcBLjcyVmiLSnYY9ctYYnCqmBtjeMPz2RLn7G
MjRCWy2o6NToXsroKP5HMmVsPYI8gWTJUZ6M4NBKTUenDdIQDoUR3xcxYtsXKMca
qYFA1G52uVnHHpbLZ5Tu9VXQf1EqT9sUCr+wCd8g6y9z5gqLsqKA6bmyJ++nQo6J
j3i5mm1zJP2+8aUD/zF1Cg6EqYF8uS2AN4o8s0RIskyylWsfB5cxfQQIKdgVNCKw
PmF+jmTgwmPqAF2FrxMjiNtLFxjQwG5R/HWriRc3vY19+tvxo9Iv8gHvkhkKyzw4
7WKXrzQtgOD9Cw4+aCjSYUwBonOEFCJmSvE8GQtzE+yG2nQij+U//48hWvYljq6X
SAHl5uO9ZoYzmSz1GMCNKTMzYUvoPgkb5mLUNNsMOiaYy/VFBq9BHnMfyQSQEFZu
LEganL115qq6tXE0oOn8PaGzHDtIpmwW6H5CK6wXyHDM6id4v/94E/Y3hwf+nKMA
k5hzfjvk/mnjC0NNZ5k132Oz6bofSZrKvYsYGIbbonGAQ/GOxmVKjnMkQHBHk2lA
l2dee+NFx6BSPleq2J9MMef8RXpZRJSrXHJR5+niikaFQHRXVuu+B2jc4GFIOxTQ
sP65W/mr8dWUHcF9liFFKpNHNLK9hRqk3J33J2ir38BkCRGfmXtcpB1wwx4AMj6D
tnV0uA83pr4GQoKfbT1sg8I8+HJILv7k9n311C6toj8F0eBWN1yo1v2ElHgPneyA
Zi0mAljZ46lr8wozvaeBxESxUrYaEWjZS8hoGyAt6QwUaKm+FxpXkFYflo6aiNkB
t6NSzwApjrADr0Dq5wIzlGpQh0a4fjjfQR/QhP7Puq4LMReyWK+ZXnZDkqY2RqkG
G7qTA9J/kBDo0Jf98MB3uGbEpFqpknWgHWOsOkKXFWEIZlDFjtp9VX73nmsec7EZ
q56n8Bi1WuCGZpYYPdeZGUGTq9aHbh6fFxmI6INgJYPNKhlt7Zcfd1MjyqI5fGRI
da+BeGXoQ9zFLz4ASMSvV4H0ltX1SRIuQ7evle2d3R4At+hwaA72hmKCwskGVOua
H244SW84mSny9NayQ2F1rdIShis0WbOHkI7/dn/FG53s+vn+asSJO2CbemWtoQbE
zkLpzDuz6wKEI/mUQcBVfqgXLFuwFwv3UhwKOf/Oj4eBpbPuuwPidxmLyseiBmBM
MR/v62iRH47bT9mj5vXl3d4DWArbeesWIkwJBU8vWgjLyHMA6iz6pulki8252i/U
x2+Xr4vpqyL9qBICVjHrVQbetYATq3IiaIohaElc7o2g6V51XKozy7CUHlkVeff2
rZBfgQT0sAM7NiTR25Yd3qBk9fNAFloWSbF/jOk3GP335ZP3YuG3gt2piWQ/uQUK
gSFLCJdhMaRebd05vAaWBFyX8+Ou7ZnLZ0B7AXLOSYuGJohvPmrax/uKKJIh7yLs
PFOCNjMBGhb37NUhhwSlq2KAo9ibulPbhJsOBqF+eZOLwvbvml32h7HS76SC2MCX
iDg2parz5Y7Yt/gkAHinNoLgrDOW69w+Wz32DcSmmdZDb3YkEQUGMQ0t15iJ9Tbd
nYzHeApNZgTKDETVOlkV0EfMVV8JHER5KwNhGW3vzd6tJ5Y1dgVsagRaZBan2qRN
BYl8BDbqnwPQNamyaWaC49jrEUkGw8FeAPhrO1ogwwA=
`protect END_PROTECTED
