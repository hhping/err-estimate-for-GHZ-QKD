`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RCGulUPb0P1s56PinlosUpP4Flf9BEdQ9LkH/9xYWNKQ1Sz90lotGYVh+9yr5ey6
t5aQOre+rPOCbSKKVk3rzIyBeK5q26V8pUNEzFS6q+kl19vldTdIXpLPGRaueMh3
P7V83xQ11tSHEM1rSPBehL+Ry00I2ELseNmgtONVSLZbwG8+ET9ZHp2r2RWJLOar
VO5LW9JDztn0wHBJ1KdMq4LfwiyDNUAaYvpblg//nwOAzc3OxqGYL3lxvhQhSQeK
hk/O/MaMYOcBlC9qjpil80lazaqAEudCcYcud4E97Pz7Y5Jmbg0reA7tsR7A4yZr
2GBYMZqCR71fewKrY/5OTfT3uWhUSyRhkvpuiBGBx/ougi7//EW2RuVjkxSvO7CK
n7kZ0XQqBvQ1bnKkos4qleZAp1X+ogHvt0BZbhs7wY1dUYYeFP6Pmg+mSl7zxah+
PyFzB4IqRHpqpKOo+xrfXr/JhbXYHL0CKeM2maTAvpziT3VxAAsnMuC7pa6wz+p9
4V5hfoR8RnQbq+Cf1psvkiGOeK3hJ/Hk0l9b6YctpxelPxQKHI+vImLbqxxIg4Sy
aeKh+gkue4l3XbcI8JK8C3ucGYh22ANBIy9DHMcj+tkblrjn69TzQK3uHyrs8Gz0
VcoCZx1f3DQdv+HmuCLfCg0/s9v7l9eWa9DffQOHEprbtjuLvMF8AM6F2/u3rokx
x1mQ91gw7ezgC7LbdrKD3YlHjOMXWuj1VVjPXEjW0SZP1yl4ESe/AZm9oipHGAxL
cv+c+NnTtuz58YjfbE7ojUvbcGJ/0oct9S8146g8mlPUobxK93PbRPmJvOjmQvDw
QgBkrCm8sE3qeoxhwavx0RGZnP/caveIgjVM0ihbZc7y76Idii0EuwEPQElI9GDB
xoLeSkiXOpT0QqyxASF7Hq5XvQzYQOkZsySfTMiQIY/maFfts9s24C1t3xjg/NFN
4D1TAKAMyZWNbo55MEH7obEAcrr15ndos3EXywb2V1/PHGjMa/di/zC13eDGLxnm
t2UswK4bIArSDjfqT9R/qnu78jDPHcgS55W6lzvy52PMayd0ZZi0zoTmdZ/RR4Rs
POXEzCZ0J8vcey7IxxsTlTIbTFbxDN8aV2xUpkrEIRVY3/O7Ccp424nw60J/Qx87
U23hnCOHHm3tsIwPxh1dAH/dkHOb5BpWGSwD19lcCZur4VU8MJO7vXCEACqABLbG
BgPY41XdHWau7WKB/MwQSWcqBQMHXTX3HBnQGcBIj5cpbz7ONvfUS+RRJ14vBLw/
w5ezJ+MAYNgtBRLeJC2NSkUcLmvDU883i5A2Q2t8Thl3WG/xynVLXTsUc6mKrHKS
Z6AbL1Yehx18hlCzUDde2+d8t4dEcCsXw+usdrBtqnpud6+om/ad5DtTFCHILRzw
pQsXpM2N3B0DOKbnwIWiy4lMm2v5JToiVlWDY2GEBpn2Gc6jf5uZzpnByXuEQAPE
Xr6b3HWZQW8l6D83mxk2zPAKh+3sXFOJJxWtgF5URTdaZXSgAvzehyqJhlrSXlv1
WuC6RVzxahLeUprF/XZ8rW4Rr9GtiTIyGpFIizSWLanJfKw2kL/UrWz8786j6eoB
N3JQAB456bMMKpiWZqJAszVROWqMrBzlzyJnKys1Or27WYug1Cx8pgEq1X8X7eYk
2iFDHyDRI/c/cf0dY7CGun193kaTa8MzpLf1T4rnptYl0RdDcTZESyou7vdHsYrD
auFQQnP6xS9DlPLReT6q5qUTUB6fOyJNaXHITnIYlKe20BB4h7FjtCgklOqh+0uh
TRCXHL/GEWlTOp+XH1z0MrY4hj4+h20ibOlA7YcdZfzxbrzXbcdTX9gt5NJ4CUyh
BVhFabzvq7ba//3MJRd3rjf39JgBPypWDfcikmpU5nnNZ88VfZ2avELQ18IV370Z
qC5E1UHNVohEYnV8aQRL3T3aGCZyp2di6bUJE+k3ilDHuiud/+0TqdSh67tmM7gU
xRPfOsD4c1PatJpXciFydibNAC8BgOkCY+qHgX0SlWm6A4mxCcEuuSjz4u39nxYN
EIfov3rzp7WvJN368cR00NUdkYVQKaQU1pH/pSaQ8f6ChI/UnEnfg79u5j6TPPaP
+cu8In3/8PjHYbZs0qNkqD46kJhrqtWNLROOO4pb9r5nX9hyARxjZy53tlcriWBk
gh/lQb/BJq3zzfnl8K9/1UzRA2jRDNP/uaDfBHstJ87OgpM748kgPSV0FIe22P3C
vors+wBz0ZoMg5ZlHtn44jM85MQn0YFRsE/OhKIJaYwXulnCiPPCVseouv6evRNm
YJaiVLBWdrBT6y6hqyNqpTYsZvTKhwC+7MXJ9C6C7CoWgYO1pMKFkr2WtOEjjiCc
xNEuERYWq9oIYtTHrCHhl0rRF5KdrlVXdKHrJpZCZUtg463xUVF7UnKxN5ZSHQm7
wDGgsTLwB3x6lG3ChS0GHWQIgrQMsmuABHe/YlWvcM2EYs/MNG7E/ftlgyOcgfdt
4wfjNWUsy9RhReoPa0OlGE6BXN2IO7ca+LBMp4Lj1KvlSFX3q4iQmsnath7Y90YA
/b5NeeEOh1ELdLJvu3API7XhtdKXTj3AdgZKlNDLFaoDHppUv2JZJmAbX7fv9r+m
jyci8VyKPq4e+wvGqDR3wNeGbfOoL4hlZXEjM56K1pFkB3dwgtcKZBiyzQuoo7ra
T5+VY3mZ3zmuTa4X+TY9RnBJoABaNT/50080Cm6FzKlgiqQ570RUOuQ5gIZOYgv1
DqW2YIGfaTHyKF09yn0+Q3ZUXO1aPOorZFqPdsIZWwy5WYDga35cw8uGpjlBScT3
/tVy5FjXhqsvO3jbhI33dhHdcBG/bU72bLd8IJqJ3NsOXAalDd+7HJJyGSEIjVda
HR5T85NtLmGi0hO2z1Bpg09HuHS5egPHr6p/DrS9ow2mVIEjh93GHzW5xSrHL2Td
+wQKmYtDXFCU+muHRawKj/m80GtG1F+olV8kgqXHeztp7nar/w5LtRwfkG3CPS07
ydhA9t4SPkpLzxl7uLmwaKmGbyiu8v+ymgAKG6yUBIv5ejP9ysXRz0bME+fbM9o7
lNS/Cq9FxKZNvo98WxWuhmYw7RTDNmZr68qzqRynKzLnv/aiEHWNUhnUH6uHsquy
d5iYxLRFRN/3wRpNQ+DdnnpHNotoxPjnSXGjg7a01pTceicHSRrbzl88wns2Ag3c
jIEw2Q7ZP7HhJTDuW5E7EAvQIBMIEXr8ZEsKW5GrhWegQt8Sv6li/Py4BiVCLTNQ
Ec6aeluC/09V5vhvp/qNq0EiTAn/tLKT7+xRc08mczCNMNlb4rcJQ936VtlmPP/8
x8zeHso9tIU+bi/iOxQARAQi3S8uB9wcZ5n9/ROKOoy9e/243TzN3dUXY64ruPcX
FqCtrn1U0/YAwYi74X8RbdSdYzJm1vVMqFibW/nmoKcIfxsKnAQ0kUdqRG7KZwD2
6m5FkOwhIzjto1bVT3cf1OluG3d03OlrLkE5n9DNQPnmuhUfjFXdJsyPBpKzwHiQ
Pe5XywBRaNW3pOQ6aqIV7dTyFITJrjwVZ9UFuSXu+5CSmOM4udtc/mS+HyU2GLlG
SkKM9yLuF4NXsqusmZaPQnpbjuQVEVVMOped9lbzrn8i0tmmgz6KPjKCJl9jhaE2
FD3f5veqKKqHLFbTBtWQbFFsCNtyh6k979ljlRg9/QMP5xjlk/+aEwrjAw5FUPZN
HCwP7mY8spQJMfDkOxjnECaNnu4UpLbWGvfzF8w5HSA301jfivoZyHhCHnEoaMeE
xJbMQo8UttiuB9fQlhXVbjpjbm76BGpt/35js76Uia5JNwb95Q7iqnexTe+TNmOm
/MemlElx1A+2PwkVDtau2wRsVHGCWz9SwUlqmCEfUTcN6PL2oWWJzrjGk3cx2+e1
fJMtdA9rLHlkE9AA2xg+0LJvO2ckxFCFQ5ZA1YM3LwG3OlKoHT1zsVUlZ/DeWj7e
ebwPZpI4rmx87bNZD1pf9x6oGi0YkFEjm+V7MzzPDwBoi6DLSzl/gfd38n2fS/ph
Ea9TyASkSkSNun/fB5b/trUSbbvIAM0K2JisysviEcrnfwrf9kx0IT8/KxT+dYpZ
h1B9nyEB/N7q+BdQi7e0gTz+BkPfHzKZrxgs79Qi4Mo=
`protect END_PROTECTED
