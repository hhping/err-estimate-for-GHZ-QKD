`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oczjjb+WqgpObf5l1X0YPKmFwfp8GgldWzK+GNm8M5O4J3c0vnctadVWrlti4Sbm
javafIgtscuPIGwWtdhubXn7QhStO3kEyTcHWmgVZ1v5sKfty6AFtSofS2mMtBRi
fZ3o9rZF5RbfatMfVj3ocvcQpag0O4/1IQG/7eyO7ZjPAmCdWzirE4RWQC3BMwFW
4J+58jpf0cbXnXcXoQB5e2nVkeBovgPZYE+RpP3t1OLTOQeS2GNMelQW7rTE0nog
AgqF07X/kvkhigmwg5sRBlKWDuMKxo5oDkUIMKUSBdyolseck84608vbXHwDIe8o
venaoMZpQbH5eDWDS2gXyWygIHtOgCNyDHoF9H6xLgNdgGPG1ChzQhAufvoutZ5B
xr/q+DOSUdJaJ6ZxV1SBgT07VdoPkEZjlItrzjPRQUmbFhpWjuNsuCrVdqMMJYbS
CT4IGfX8P4GyWPxClhRW63QlGPBi5UumzFi6zPpcnXAvaFE1j1Ct7EOWZOF3tFAh
SZNCJqv9V04+tvdfH/or1u3lPQcS4OcFnfMaZt5vSrB5u7exp036pTTur+fmIPRg
P7yA3f6EZlVk4BwdRRDNuXvLhUBE6jwnrkgidCDY2miuOu5Esht+1H7wEkAFd6+A
cQYY1MDmVzEyckb1PWCbMMPM6tAc9aNG9XTZdPXgY05lwNJBgQy1s3tTkzK3JJiC
0g2A3TMxOXLTxuoMbNOZBr0mFZNQIAjcLlQP1mperKtcFu6mDLfGVcp73+eWYbHG
pqPYOfGvNrP3uBxUTEIoQ4Pq3FlJEt5ChG92+nGH4AYjyiOhLyQ3do0ZoAz3J3Mp
lz53zpZZJ7s19KdH/tMkeBdP72SRIHw3SxsQSuytOuEcSD2DWX8YRs5AAHiOhmwC
bwtS+eT/MT8ardSx9be3E1vW4ySTtSqMJ6Ex0AnrowjZfGHp2w7JA2blfKYGov1m
El8ta40o9RSJ/UwZ2xeGcpQBaFTkIYFqvzchOFU4hNbVxKjf4yOdajCIC4xuSRAb
pWrg2MsJ3dKs5a9YF19ItXatXLeB/OAjrA4KS/KGIMMBHnKa3hBJII0yuaVAwwZq
`protect END_PROTECTED
