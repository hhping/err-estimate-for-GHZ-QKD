`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8/g2HZymTpu1X3v4fwJP+B/V2XQYTs9WRZz0Jk9jGsTVsl4Mx1Ed6mdKdZt2X8ki
MhnTH61/bBILQBQLSlcmIwUDQYOzQ7NjUR9cJV2CaDNFqjGANtxVkzpbPk9z2yR2
kvTsnR+SwGRKh9N49foDDqqxkLZAya2bHN5GnI0yURtcXFptoir/nIHo7JgXOPE2
QkyWQLOi7grJwbDBw/X9zXp5dQo2BpPfzuGIlTwWarSt3fpwg/lyjooqPMNixIvy
MjqWWD0NlQpf0hUQhKX9fzPQEOaGeP8FLzCrpLuaHG2jXeqpIoZ7ke80a5FiTSAN
alf99q5vB3Tmr3Rzv6kO4bEQBhwV7cYFEvEMp9/QQLtZZlGIuMakaEs68kYFzIhn
sShSBM1LXojtyWOu9MoVvhnjg7lDhY9khSX9bdIe4MfJGFkSjHCIjSX8xvtFUd7s
fGo8dxWb5f3MIpBwYsB3shhepTPYkjuJmuA0CjRrenN4OZBh5oa3y40YaR8CjzJb
2mMwadAalauz1yLfq9Wxv+wyXRvRSOaOboi6Djt45OwHKdzh9Ss6g9kDypru2k6+
GCkj5hAKaYBbuJGyycXKtN0Uq8c+uxrk7Y9LCuXZ49vVVR2OGmTjsZW2GWJg15hP
tNjox5Q2a7eFZP+x75nEgSBQW/+hdo7DESX1nf9xGZI/ucvVlMM6AP4pu+ppukGP
PdPyzvhxTMxCcmXqjLUNU+cJo363lr9zDN3RMvMybV/n9vwtBk/6euSQVinX/lu9
H7BzeZ9XAM3u1Y8zcJTcVqI96Z7oOWsOzpnlj/crRbM6SsP2Rx102PUadpBYMBko
t8rGoKaa+V6gnq7rzEU3uENGhNrkj9IUWMrBDiQvUOGz330byQQnyMZQvX56Xn4l
J+l5TG/x+Ym4v2u26jDCalHXQmZRbTLYs4Cd5TgtKCRdojKI26n8rGmnDjO7KpYq
1phjor8pzGHxS8lWcElvr+nSLM5y6EoKpo5NQiYzYegOGHt2QU/sxeHWcpiFcuYK
3oxlkYsypbY7d2CN2eRfnawPSBkHkv1ukZZfQpEB/oPkAucaHR5DHYZPsx/5nXp9
/G7emX5VrHLLIGcnoZq2Nb497DOSsgGgfYWGdqFnMCkmQ/aQXB/HkkQ6LDoR49uI
Sc+L8rqh7hWYEY6xFZ28RMd6iz2kND8HejfLfjruof1u/4K+OhTv7xm2EUNo4lqS
s1pZvbNtjc90y2EGrvzt9cVvZW487mKwRG/NIWujIkx829pDxSgXy5GOVZcN6HXU
AaO3EXBPnsjRj0mrIBSmOHmrpDaW6RdYEL9vnV5VHOfnG/BCIiHe0bOS9jgB2G9I
tQTRIkcmK36RCfNMXE7yagFQGaT96K49lSmhND5lszRgfsdmk3it9I+gA0T3hd1m
S9TUjbpepWvh5ZBBf6/sqlkLC9dKBqbu4Kk7aZ18oyUtPw4qLAJYPlxmTTAygjrc
hiSP7m2a6l0VCl7c4zjz7TCngbsHqlZs84Ck27tmcuQ9MD4BiV8+VqWfCafghl1F
MprpJ4znm2VuuZGcBJ74uIRWqgEtfLbO9eSyCg7vk40=
`protect END_PROTECTED
