`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w1SJTcq0DZPqA9oLO4NWKOWw1FZNOXTGtSbt3Ez6rdfVugK3hzPoOrXtvRlX+rkt
VVGq0q8X/9gPOSZ9G+hfyrKP7J/olr+EXOfFF4yf8bBHzVRLNBzl8UfWccZjMpBJ
F2zk1cNKT/CeS/wjOB3ZPJFlZQobcBXVBkWEaXT3RTMDF6X2L0NIS4eD+SCDw0YU
Ma93TbTGPWTHKAuhRz4BubM9r9j8TTL5eps2/wCmBn4GwbLil3GegpcRHUUyKVDn
5mAL/2hUFgPOLen5awJRcEoU4g9q1mSOmP8RgYrr72pRvn+/W67zUHfkx2mXQkFK
jAIvOX1PC5jP1C1vgg02R9vfJ9nTQNf6UpaM4DH9/z/6hM84B/LYgogyX5jkWY/s
hOxYZoRSFgbGgtOP+UnYOTW4iBjGihE0rKwCGfm+BVBUTeQEPF/hJ+k4vIM2RlYu
R2dfYEwZGK7h5F3rCpd9FzkrZzFNKKFjZpeI1VAEhf6yceGkEE/ahBcddwEydHRj
odBZVcpFvIhYg0OUXwZQdeHqHGZ8d3n9s7hz3waFkzXZ4NfNfBXj3BipxEQ2R1Fi
+HJBnWvxeOd9V9dBQXpldrB+CkH3t64eMWQQPSVRRtQolMTWBBQSQSpcD0Kn9Eze
ZJ4kOKQz7hI08KZihdWzfAIssQvC9w1m0X9dh6LkPMjHxYK6JM7wwtg0yqhFTony
J1l68gjpexne6LilGW9kf9omlakbIbvDXeP4wG+SiDbH6KpyaYJBWRDf1CPAVBY4
LtAD5HKeSDI71OtKFnvEeaIOx8ztKfWzX0hIavY+3Wd6vKqx3RZX6TOiSTNT7joc
VjxEyW7lM7xVwQcAYD/uPnNtzNDdOOuHcIk8GSGtgev6vtpVkxt0t/m1cu7tOabm
pupiALmDpnRoWX9rGaDtKUEASzS/334r+LLJeWscHLj/v2FcUNyBZ/ksMWnQpdwg
NEWmc+J/w4O4zFMynI4f6ZPbj88Hdq6SSC5ftNIFuUlEpo3VTpauILg3vKftHVbi
zK8+Bihia6/KXS1PnycqbIGNNwy7BwNqubOFmB6Z4zeBeeHuB48raOW12qn4UB8C
26RKtFVmP+dfk1LvtRZK4gR02NKzQH+zMZ1qYxgePyzE4MYUDhlmtuZp38MPSO/6
F+MpIAXMAOljQ6VVflatkC0lub/uABG9d7zPjWAAHFODw9OEToBze1O+TNUKDh7i
bpm0zdoPAPqyKWSQtdMb1u7BaWmuoTVufXl9qJfkkSGtf3RXUMYvN9o1IkjSWj/Y
4jqRxFygzvm/SIOwP/JcKjF1AdftTdxeAVCfMRHKoKsLgaaRm0xJyUH5omCQCGJC
/kvGG6ItViyVPaIAR3QYBM2A+TcELm7echu5gxpCEf5AioDahbe1urbY2/IHSrK3
DTN3vyk46tfP6Drr3hm6INrVHAgrDEIWIobe6QTUWajCbaoRAZfUBZ1tGKlq5Cok
U5OW+GMOEjDE2/Ft0N951f9tEV96N6t4Lz4UFuhTAWxxQl7ntizBtWRqtF7fKZiK
ZC+ACvikoACQL8XYmlFN4XrAQVdg5HBh8pC3D3ZzFGt9ro+6H3rADq74795T8kVY
xofNTmG20gypNjJogQ6Y/et8oaHsr/dRAkmTnu9xYEx3gksxLibYSt+osUIautx6
M4xfHn/NIfrZqJXwigDJB86EQdIHmVzrqDi5j0qr15DkWPBx6BOQpYJ3sGD0l8aD
XUSYS4ECoVM2v0Ewdchfiew/8+DzDmBulaB9MxGhMeXup3IyQARCyKcYZRTwegBB
xLQhdOUJw7BbWY8GKqrLSvFR4dwwc361K10Z8F6NfroKfM5zuLTmFKSUixnBX6Zg
IF9u+HySyRcFixeSfgzGbuR68dTD43OUWxao2syqsgXkKsxtQr8/kkXzXL+qOZpq
6AChy8UL15oBLZ3IvbLSinObzk5YU+0aFovyD/ABCASZIDULyFo37g57zfvrl7zJ
J+dhpQjdyJ9VSeGwZZIewK/Hilfk9tINx1T9PGIySgxyDu41h7FivNhkmNl1IE1G
QIvCSkuD6hlC1J6HWq9kjzXytUqdWYSbsShFMz31Csl8b2DCKCKLc6GGDtEgOQhD
0TxW2SxczN2pBrUku1ll0Lc+V6FqLqEizVdiU0qzhyh7umssoZdUuBImfVb6iuvX
Xl3AOYjRh2iHTwEpTmwKXKHr0QWQCEYK6e/kVROzpgMt9wybyZU5u59qkJKv00mQ
CD1a9IeBLqxmNBcOueA7DfJaFV+O9k8pmBwZTx0t5NauXbAZTvAQbIx6MbsLPdMH
qr38YLm71hysqV94Yv1bHQUMjq/VMywMJeVYUUSa4yXYrjoPBX1Mad6ibG/OnA5d
oZfu7enZ3FsfhInu4Bavn+PsL8KQXFBiHST6w/x7Zii+6OS/3wTAhTcdCW/9EGyc
KDXJI83BrPfshCLYnRgWAMpGXOUItAuEs1ycgo037SvlfWZuSllE4969edvfFiYK
tFidLGTDGdso7XVN0NMGXuKQbWztMNVfDri35nHUAUGwH5N0LoeHIox3HvzdmfZ2
8AQjx62CPFXLCTISzbVfcLhc1Orew+O8+bTFsSdBVs7dz4PoNMvn4tzIn39A4si9
MieJ6Wbk0d3SWlxdD0sV+lvr3Lf60MesVKYZf+wRvFy4XSM07foHTKOh4AAfB5wU
OW3ZouqKuPZlLf0SNNAaLA384acZep2ycgqXXNjKn5DFSmePeTB5KnPqO1hZQTlC
C+DDZBk10ECA2o//+KQX7P00gzDeycdR0CJpV0N5gZLpqMGJjxHpTVBpuVmIxvuA
Jc74G+2HLmPUdej2VT1KummzIz/hCKdr+N5QPqXm6oBBxyqBNug/a1iMSn8dnsQM
E782KSA8hNlIRi6JasYZbXd/9iLhtCydLltIgAIG6+Ihg2O+ttz1g2gb03WmXPa9
mgdUgXf5ZBNw7fesT+4+4Hh8Va/7n2qXCV1KTpK5ZQhGqbt3ou5PVNftsn0zmNTW
UtWNgjKmzKx4GeW8cEpf8euBagLla8FUPisKo0/YSnI0dvW9XIaCW21mlKLNzM+H
3mUiRAwYppric1cWDutyr9SmERtiQYpU/yluAgVdjhjDLJGgdC4LcYiiVNQvfMA/
2Hyx+x5ftnQnI4pOu+Oz6Z26OELV15QayigyQNqel1hbMIn2R029Ig7NrOllx5+K
YTh9PwWOH9SZt4V71VhA+Wh4A19sYlnVjUbY1oKd07e1TBshrcGOXbQEAI3I+0kN
xXaA7WbTkuVXuEJmI8GtSuS/dQRc+IsvRcN5cJ6U8uP9PjfIUq7mN7DACZSQpFdj
MXb9Hu3AoXM68O5OKKhxonsxjHuVs6SW3J539Pc0czsulsSNXe8BoWSqfiHKG3lq
Pu7Z8JaDevtgRvqHCD7D/zXxjDfI3kLQ6pl3PLT937t5ZrFyK/K4kNN3HbP+ueqb
o9Tt2T59tqkelFls/yf6oL782LHe2JtaqUWdDm9afcI7VWXhpBd4xAT+cr6F9cPy
kLUEyo0Sp84BPgmNfhbNrNk2uz1c1LxJ1vZm9fqoHTzVRvDH6oB+/Qm7jyO3lIdq
ncDJ+mCE+VyjS2q05gHcJ8lkGLsl1+2zGFhRZcrGFdEabWo4fvqMSTp7bfV0WrKk
Y9GMom4HXlT/r7FM+OAd5x5ZPhgehEF6llk5Di9YzUmwRojOHuIbycpigNr5m1Ya
qc4iDf9lt1Nwe1tC+ijntQcDqj8xL1jZCMBb2gQ40UpngzV67QdxKOchYz/FOV2g
+pK7PYXzbOf+vzVHkmbS9BPFljiwOhSLNISAVC4Gea6+3fZh8XyHxOv0zNXPqfFy
ANWN7AuA9ZMawkoHH9PEzb3B/aZEt6UGJ/9Mmx/tQ9CMdxW7NQjLf/SmVCXaHjw7
hs2SKu/W/tx7XDKfbH7cEeo/u2yK2znYAkz4g+BlbdE6UqA4XZ5h63OwFvIPvuFw
LPzyDehbLA6N93HPOPbLAScmfUqYx5PROkXZ4nVnoVvtR4F4dONMAIhI/2QmLMxe
jkEMbM3lGY5DmUKVjKC5XAltQScmIwn2rZD3LAJcvmT9kqPCBQpgSd4yiFv8dN2+
L1r0dkXGRn6bhTzF+mIYMih8mZEZsFYeFBNd8TJXKnMLApfSbkFNUOdJUvIJfeci
Fe2tFd3iSQYLD2B68zYv6/PWwDlkiOsOB0+fz6eFRCIU4SqzcxoWq0crvYLjlyZS
YhXjyPasqzPjNAcAqA2pSiWUoxhwTOvbRFU4/hjg4k0KoStXUyTGX+QWlVw0rSGt
4zMugVTwK5qjsv9s4fEz53yOCWBwRdBQTjLEo5mxhxJLQJT7cjDGYmh3RCppkTXM
nL5LuRi4Gmks1KfJkDiFlaXFh5kYhro59svk36oJWaO+ZhExTVewt66fvYWuTyPW
WNjH8PBcwDp6eUlqOwZr1mt7Z3cTveihZHwxWTwNRyEP+0bD8YN1FZixbsecgY2M
9o0q8Vlv1nLZ7M19gPCE72px7+ILJPqRhEUrDLDoq30NQfyguzxxezB0RwqVDk/Y
mDTUaF3BdZfRRHcVAK1y2et9sBaySQIX8l62HfpQNj3XZTmpHs98C+v2/2tW/IRt
GRVL82Z81vMGixeGGBjMfKbtEQAynlk4D8JHk+CVkW1vbk0gECVdTYaSTRGZRELb
wQ33x2vawyDvlhmV2l/Jg9Mg0/nJlKsBEVOOCnO+2klsFHzmh927iAEp7dTq+5bK
ZXKJAONj0cVOOcZxP+EsWDFRmJDWIZQxMA9xWc8yqDPtXyeRE6iReKeLnFcshrw+
Z5QgsPrgLg4DJ5r+XDr8wdrn45boCDjofU7akHdVxgCFixB2xmeckLWQieAzmvBm
+CWDqQwnYem4eJF+kInBiUCz9j4Bqpq62mv5V8T/d8f0Bi/I4RC1wZbGfeNjpk5W
+/GS1Dxy51WsKEwAbkQSmxNq1loGIkrUiXrE38CAQylW8bdyR+wVZaKa9fm/iUoI
7io8zpNIc4napsP/9QDLev0/jP5eru4KMfD8mL4yGxWo9das3Pc/dR9W9moXaLkw
tnIOFatErTXIcySfjUlVNN/iUxJgXjiFBDYvJvKsvae94wVXSDFCdbpWPqR4OfET
RI+e50DQb5JK4S3FgD3KFtcI1/qp40Escbm0ib9WPGFg8x8bNsN8UnLZXJM4q7aG
ciL94qTV7S3ht81BZvG8CJZ++auoGDWQ0kLD5a65HqUCW1xM9KB6PsT9Vkda2U1c
87fI0dzdjI5XRzsHYNjQcQkZ13y4SHLO858zgOytT7gzZbwnrWXVj3FANrAHa70C
C5YxuxXmB7n4L8jTWgDhpNa7DX155tzRywQfqCFJXOUvmafkoo7oNmplgRrc7Y13
43WgyUNb/aNqUXLqdVwF3DMHCquGso1iGE3hzBwSWGW+saa/8WuD1pj/n2TxAIeR
3V3zk4Dca0Mb6pw+sKtP3f2u+l7Y4eFGb3L+q1DqK1DPW1kEO/Uy+pqGw4D18Vsd
CsBO9E/CW2/iG9dp29abom489je2lgRPnFFptXaSdtdMg4/rkvA73Pq1FvHjL7ww
VwyZKHUOOjlyTXx5ssC6nuZXI7zQnQ5HSjF5X1U+hB50ReTrpLag9oDz4dwRE2CR
vxIj9kPFGFn1+o+ZVS8OkLHadsFhqVo9jGM5ALtimfQYTxrqXjRlUsR3kAGfzZhs
U2/xMo2qhrQvipkb++CKN7JB2MErjtadnklPDX/Dq+AUmSAdZhfddA9QRxAwb0/R
mUFmD2DS9X8VuvpJ6laS6qQi+BNHlDKOhZRRYYWJbmjCYmqUI1pURrUtFeXYB7Mf
PVYgfDyemDyJV73uhNlaeFgJAgm7Jo3pRgJ+kHwBuU4B0naIMcIa5aO0Z0/mnetU
7+nZq3RDF7z9iZz/ERNG+rMBHCYOcyB4xt3MK4AmzW7rfWLwI3GtLWAV9HCDJM37
9Oan2yjSD7NP/f4VlVb7HFkYcTkv7uf9evGRvZ83Z3hVXliPmhLNzl7A3/z+DurG
6JYF5y0yfeCKqpeL7kT1jTHZp8YOEcWvz8oe7VnTXU2X2SgknD9k1DPXCfU8zTgv
dw8/XwUq32XiaQF/ZnhSOMRyj1tzQ+AMEnwdM6pfRqIFAVoliE3t1D4z/gFraFzp
F72rXm31qHj+7uBeQ/bnBB+0luVYYIHfEGfSFMtySML7srUGG6b7iTFtkdsIWDcw
qprtm4OkdGr+nI64KGMs1m+seXjYuoJEN25FtRXcg4uCUgxEmUxIzuqQlC8aXF5T
EMDnQPjfbI/ECR8XkegI5gLP6wfiRF4UrOzbAcvoZfPs2G/pCS3nVL49LZOCaEIk
jcuHPYiFXGVBhg47Z1AjaQrkQGyGYH68JjSGAWPves2t0KExgMX6srybOqBIIY/F
SwsIRscm7rwPFLtaHBBnKVxd+DM1Dws7AcqkhdRzJQSeBrHH0hFDdZE3OnZQ5y7P
oan97lcxwWsS7mVIFwzBZIHBI8VIYt+N2IrWivPeAXqjqK6vvyv/ZP9lFJ0Aht7i
7XZ4mnHHuujO8xv2/SjWYZHcXX6ENA7vh3FRu51SeIL98PZeQT4hMP93qemC8R1e
pF9lHb+Lr1xoMTWXiVOR/qwB/aOg0peC9Fwu31cbfRxUcOyIZo7umiRTECe2Nal5
b+tzMMJE+iNjqOIgOtfIl9dG0OpA9is4SgPCe2j0O1alkziD9k3Z6wTJkhk+Jx4S
CjJ60NyTeVPaQ0Pt7qczurNIFRJjjE548Dza9IJcXivbKib5Z4wA8XN98w3LjG/t
qzUxxP62yLtepsWeJgHZr9U74DUHwbug+BaBsA1OyktoknRbQORbf/QsBrh1Fliy
/Oo0kguubgs+W6OLOtTRnWpohp0tGFQ9gXiHxrAZFNKh2acvIik0m41Y1Bfo4ufk
XvZfE1ZVMt3UOr08GkKPe3avqwW1kLgJUBYAwD6ip05IHCeKXxMn09VTwuw6y6Kv
zSwFysqetn5VX1iOttap3WEud38ouYhw5EI6V8n82ysUq1EHyrTQWIV1ZtOkBRwB
9kpZ241IyMUBaGTLe60VUGXFHwiJ/EzIH8m+ph+vt0gPZyZQXGLPqqtk1JOIBk69
W9e8Uz0H/GKzyWUkVes8XfzOlHBHpovNXUPYlqdig8t9a0cVXUMRhxx6rn6LWoNj
yQOUymIAxPbqeOxIEXZf56Cgg+XnqiyBudiwoaNi/I2MJlJYAhylzEHx48UpKiKs
2txNNhY06oXD7nUtTQZTe1PDhEqZoaqDfLt9QBlDE7sETJQp9VTEmuM0XAzl6tY7
vSkWfXvFvzAwX2HsQx2oKAFp7/InOveJ3FgL6ZreCcdORufk3O4x9cIpNhkWncKA
V6DcTWZZWzQp2eSX+58e/2YV/2/ODhv/e9hxZNcfBAog8YVoDX1a+qwAH8Eg7g9k
yu7CBN+mRK2+y3fhr8ACCV4UwdIP7+FjcMFkGNwDE6GPKqM7d3EBqRjd3uV4YNFj
H/KlRY5ZxE+pmFtt5JApEIjcj2zJwM3v/T9WfnsOW27XMfgr/szTB5LwCtpR3rP5
lcnm4swK39QtGIy0RHZ8PFYA4EkRX47CbBtmtCF0vH7uLGvHE+PPWZaHHHKCDjbh
SMj/Bw4bGVzR1DKGni98s4RF1pVMlqvqsxW9C8VHdjUVII0S3aANYR8B6KIjCE8K
3V0+lQQcwJrGFK8kAWpN4LQA/MTNUFRvnFV71RL1ihgyE8P5ailqnhXw/p23GJKs
vu3wiyvMzuO7vVnnTu1bF4848i5K8wZ4yiunBjIVG+sB4MDthhsFWqf9S8eEdEkz
EptURObcHHI3GA4HGCIxCnmjIaiwzwU2bUdou+5aNxUa0QiNK9izyKCvCdVwTphM
5+uip8BkrjfSC2yEl6hNs/BEpZfl73zw3kobtt7bwzhnEFusKMwAcfRFfXYx0JC9
64HSU9ZpTi0jf0I+roAdHQBdbKyGBgmBisJ0SBIxTTlBMvhKs8c6RI4Xz03LnDRH
vLPW7QJlD2fJf8CR8/Zt4lusR2P/PnTmswur5pcdtTggKI4K9bkDbwu2Yyn5z39t
jbC/DSFIu9oNRNVqe1IiSzyxmKg2QbhWnBZNVOdNihQNb42KtszOu1w0OWY/p1ZW
7QtTLm/82tl+DWvA6eG+j7kBSDLPseZ8WrVtD0JJOSYVRkEdMVHH5EvOREi83xAI
xgsmOwG35s2K8u70541WQszIfCHdLu/NhlbDMkaK2IeUurf+D83u/01dyvt//Fcu
P3i2H65Nxv8qN7/9s3k6xUcrD2Z8qjnfYTMAqPdywX7rfDZq/ZQl1CXECmSBqY4F
YyZUMRPTpumYfq/Brp68p8zZwMxZ/cEaLFkPdXJwVBNGzLO4nUWf38LEpegGSNXM
Z95RqFghgPCtS3YHA1CGpZMcLuVTltPA4sLbzAbcfITj7TDpZEUmZlU/Ms2FdtPg
2p0i/NfbQiePEx+LOKlNlbBw8rTyiGNzLAbxSrATVX+othzwmjW58xMJSKzvPfrH
zJ2yukfMDJaNiKzOFEMWJhTLQhzSrzSER7WCC/5sL66FQiV4+3NDJ8eqwFIAm9o0
/FVW4WUnp+Z5qt+7rFpcBKTkPImx0XUnIXbytaUnRjoGKQhbv90O9cOaL2ZPOW1n
wDuA4UnP7FNBj5FS/5+2eGnXtBzuBLgFPe8wKpY8eYKGvvoFhyHXXtOU9fBDZCOI
GxreSi27Set4wjuKTozGy8ZhKBWpQbbaPlugcEyq9p6Mq7ons+k+WT4tBNr66QAy
Yo6jW/zfHU6Ekw70fhtwJuY1LOyDSctaARDHNcSZIl5NZtJH0Dymwlc6ZNuvLlH7
wMxBEr919wZk3RQhc90AmdFHJThJ3/4Uq+W6z7KwqeltWLDtrSAD3ORTn/Nocms5
sXTWEeoOKh08UqyyHrySBa4SeFKdSgborfh2/1kTAhoGrJjU5gqqwM3mbebju4bb
bKmHqwv9FM0VGCrVF/bmzMt9WcIkWtUE6Pd0Izv72kOrPBiVUVIMZQ0uB3jORmyi
KdLUcxjJBAoz5Z8Ps2bPS1ID/1o8RoU0wy9rqPCHoOmgqRhBGKkLlAKuxCAFnQGy
t3qTZzjL8KkTXnTgpMpcAc/hBfL+GoMGMmFl+YCzMUdpv6IiwkmQ6p42rkSsBZEZ
MVYicObReq11IoEPYE1bK8gCpG1ThE9zipuxpnBVmXae12yRZbbWzAjd6NZ62/cY
xoiRZJ1pQvkGZZGADdVcZ4A4Co0z82zSemsSui3U+zXah2TGY09HmaK0e8K9FYfS
ltXno0RxvjyY3cL9KCVxB1VjGLvBrpKgLp/tSht5/h0MQT5VEPjpg9uIwYxQL65x
gaLytczcq1JLto1C8WMXJH7h39eb7gJfNbfXuy0ZN8FSYk33jUb5ryNkqLG850o7
6xTHUuVb4fLD0iFu9eRqGMw23DhdvBSzKbqd2uxkEkaWwu2ez8UYSqsmw+rd7nIk
IwEMDKD0Q98uxHGWkAMk7pGxHz85YuP8zdRwfK9ApD8bM+G8cPtUtOgM++uFvE8b
YvxZ7geFIsxhC4S4WI8AQ1AtsRFjHPCdSECmmJRjebo6dWJk7IgEF82OmVT7s/4N
kQa2yvIzsyp3M/yAfyHltXbYcqD0FBonGAdzNmuYm+hhVHt3X6z10SE+wOJFBu0v
Jd6Ww55U5FmbR+gslO6+FK9ynKtsMHXzGHQdRCqPrf2jRZIkXZSt8LkcE2k7ZRZl
zwQMqT5pXGEYVdpx5UfAI6Tuv58Sbzq0qP05BnHBPh/kqeOenmA6jVUU+2XQS4xH
EDyMu2917pas0rtgiUiWkxEh64vo+S2F9pPMiluz5acg9jhZD1d6sNXLe/8dv9wR
6w0//zW1iPH7+ZAAisOau0Vm+li0TKVs3+35Ho1uj1TGRFVOACesQMyDzgxJJNEz
IKbA3oKSuS3WzIlslaGF4OFjw2iq64z7B9SbxKsJKK6qX889Tz7fS7+STHfAej7a
sy4L4MkFGBXsmdK/pFSbE4pDXB/T4A/VfcEbkRIuPcy5JrwRV1XAmIsremNgSSS5
2Nj77LHwEmFfQhw3EOT/YLM92mtFZmG2ilnGZmon5Eb0agl26hB4jBSlMsLZBrsI
z782JYJBmIGmaRfuRiCkXvbMkL03VBQM6WSw4T+SGdWvboAEH3MCwqxdfl7EFh25
rM/ropROivaDPV2zwPEe6k1nal/pF09HEA8gkbMmcd7ICR5mjc6Z34mEv8yQbIGm
Q/WHPctPNEWa4WiMEO/D8SonWd5T0qBRVhvI0LeprHWy3VryQWMijh7STnk3HY1x
C14HrkVnZgfnpFBAMaQGCz9jOfsGMMMRjXTC54eb9T/qUvjizGGcjkTM4TAkJJx6
+YYotk3V2pERygxUZdQTAYeA/neCMHtQpkJZecvOBFvCEOdN/UB1ZW2bNaVl2KJP
0s5rsUF95zah+DhorkRYx5jnHtc/fcu09ZsN/6oBXO/cQ+s3p0HlDUuyzd4w6mFa
HPm/pIpvOcok+qqsbV9dyiA1My37eza+VSw/yQjEbnnLCPlA86jECnqfzeyJN9PB
CfuuVK4IvFkvAkDduzD3hsijVKzRoZyIUf1vAxKeC5iOmBhoS2rdBmynyTwojr/J
N2POHXwzr9d+UAC9b8gsDmrwBQAu2Su7eLSa/Yh/yH1pyZBa9dQ/MQRTIt0cqPxd
PvvSmkuEu66/wXbtcTIWOS1bU6wQotcNpW9qOk1T2enmVgZ4LlnuA5PeILc1d93y
qG0b9OrIjNU1qAQsdXXMzvk8KEa041PNUTfqUO/N8ny5b7zSBLwNbhIyn10APoSQ
4z9+wADmSDgY+GLgiOCIbnCE3McGaxotq8YOUxwIpWldBHT3O+h3wdzaH/uXWp9f
ZkzSUxNvKovCP3/Thur+cPBqONCZs1xioOw4NejEXVq6pCYm9gaYlQgvfRaG5GOw
ZIMcIZHQOuB47j9blDIFkf4z0jWxcOGcXFwJ28Dv9o0mCP9XJ7byRf6bIQRhahdo
+zJ+8u0J6ZLRKNMOhYimLXl3Ro6n5lxYuDTrlwEHdOTRICcPoTdMalXSBjbc6dUX
Th4RKEuu+cjLXR/FPsGepf10E2lSzZKZfRwdtl7JwNZXNH5a80jeL1qT66Nb/1ev
3s0bFahInQaJ/0pcN04FTeOCr/Yk3vIX2GI4KaQ4rMCCdd6OrfYPJOp2nvbMPvYY
LsL0MwEDs9b0jloSPrxWpZSsmImmu4Fg+NKDurBYk9BjRDvJQSpr2EQL7tGVoOYC
2FYhtmn3IyXjGg5YL8IYE0EfLhvPlTCvazDCZef9KVyVZTqEDAPuQWAi8R9IEZFI
RebcLVskCXOfyvxUI7pWv7vBvNMK5mjpyWrL4kncqNtcwR/dR8maVcV+i4bfHpXA
+3Wufs5Sh9MHQue91POZG4cVP584zKW/pTrP9oQXdmTOjAlUtrs58ZsdwGiem8f8
Dm3G88V4X7RtumHW8amC9ZeVXzRqN2uFhGsYZhEH2OCYyRQ4Myj7HtQd9ynt0Gt7
kDQ2HqFaZ+0LrHJC8S8CTmqoAxW0IgIalFCclxyqUOESNGd+OqhKUFTR69YzPHvH
nwObH8L3IPqVtS3YM5vXeqGuv1s+Kc6V5LmqBLzXlpIW0SkVq2kezdL4IxMKRA4+
xMah4eiuRIQ3u8j2utTnZH/MvBy0Ev2m8eaOMEVUO1CjpjbPPmGabQ5VkPEdjicq
y4dRyjFfmMfqnCr1hQsvK0q2tU3Oo+oqRLOHHfpQAAHnv8lG66/5oy/lHgMwV5gy
YD3RQErgSWoQHIiEDDif0LiaJGosSf2ORaxJ46Vps7XtpUCOygk5xdgLmdFSLdQm
qBBlX8L2A4cvG+DpoxFWUZCvmGKK0mKkzZGbp2D74gkVnZrTMqvmDSvFmdnEfOkP
VCRcx9IhzVh2/SeUZ3GAIfSE/GSwRHGDLvi8hZYeF77RMiiyZ7Kv82nCV9We/xjR
r2NztY2vhFqbMjbGiPlRKD9O9HkvCp8mq2y5SACy/S3YsAIGNlqO6wi+C8F7SbUo
JLtEg0Udgz6G/8VUF6k20QabgDPsYhjL+/JoSgxfGhQXxQ8v39Ys499W5tzuO/Mn
fHuCjTFKa7zT+clej5p1/kVQNifI5dvASrA0hHooTzRfsV/BT5xY1nvIWZL+s613
7wvAbOw8ruvayPbM7zUUGH39z3itvhQa3ZD9coayzmi9tLmMUN5krsCVt0sUmc7X
DM8TyIuthzrp1DnW7LdB29cp+OIYpxIbVqfdsHHuqSfyv8mwio7uUfqvrT3OoMR7
sIHBCFlk48PP8mWmqUtNu8a+BmAKmFJfC4ESjcw4D1MXUc4JrDkAKaE+2l9/jRMr
YTj5Qfw6IIgcJStaKOp4bfAWEkCDcFVH47/gPOBHYfShm6cpEr/gmL00e+dTXw7G
HU+A+qucsK88Hge3AsPfJsA5ME7v1d0kUms1gqvQuuccGaos8DR/tqw+ajyDa6DL
xRO0OeQQZ8/L3XLMG23TTjpfjzBBJpct+5PPY8jeUsrY7mn8t4lp8wzKx4Numz4A
TbhnwGrJxkUriq19JcrI7kNa7wEbVKjsWhf9Id+cm7LaIsBwgd36wYh4OmvGXIrX
ZmcQ2Ge53tklVqAGcOq+3sBI/iBeSmn5Kn1YQfg4AwPpZAr2ExEMsMAOj9ZC+Yx/
itlKdhqcMiul6/E76kIduOpTGPSh11K8RX7tl7j2MwC6bKvXYPmodg2A4EBRrsJj
2igMJdi83GQDx1fMzsqtgLBRTEjKjcHZ3vSd2rHDV29BhLLCsiG9ceqGAgA0zylG
TtWnygr75AMyRfdZx316pMzSfBz2+TzJLQPUKpA7cdCObKROEiNKRPG/39qaiKrN
IEnWCDAMxFtRpox8PH1QwYTJxflnWVH7xA3cGq0qOaNERGneIOw+ZR2vOC8TX3n+
yTzSSF6U0DRE0fwPlUpDsKRwGZ+Odi7+3PEeFPX6buSfs/oLbhxk9q18q6Gs+7pO
jZkvHBbwFvzVdCsqSXk3uNAu0bx1ynSBOhPZf0UOk1hOvi9ooCbwl6D+/i3ZxwDu
R3PHT22xFUnCS905fOb5YfSySEUN588MKMR2SpblYqNUhUt2W3cNXD7FNQR+zaHQ
ZPFhygXYx4MWWYn3YUopDM2mf5x80yujrhUws9Zi4/avLGPMIUbJJY4IS8Z9oNvY
ItPd8NJcOQp2AfalEwt/O6feIL4NHjNKJp8eqQ7zDVlJAeP5niniCvhMmlP6ykS/
JZH7BD1oj27sgZ+c90TJPvCMuzvNOw0C93UbSKc4CMwaVu8EtpMeZaE7Ut1PR/wR
jFJPHjRfcELtiLUDSpciNCSSCGXuaTF4ch2sZ6jiftI3bTKa95yNbhv0c2KdP3Ga
61aJYSaRMIRmUc3HJYuZaW6Qx2/bQ/BsM/+VRGOM0eIy6gJb4hL/xYa8710DTF24
1ne2HiqrJhlG0gmAUK7vc+BdypauRd4LI97dbTWjea8mphLPBvRQzn12u//L/HAp
GUkOFXjPO08ib0+sOXXXlVRp1AcgdvSqJVMTsVgKVpQUmqldn+lmaZwtqjfBlUlQ
+0G1knYaTXQK4PXTQEQDYeAxIiesyGVDTwmnSsvKlaanMQzBH/slvb/lmGY3fPQo
QZzUvx7YnLNob6kkhsqRV+nLlbiYZqlz8w4oohN2w6KmsvQp3yycA9d0djAot/Sb
dI9WtMzgUcrhPYNzY8Vqgm2LuKvp1IrqbUzYw4gaE9wVNk/Pb989Y4d5R9MA79O9
qt1NPPr7Ef8dp8OBZkeA3Psf6uWnKmL9XJAG1ORCaIka1VUGegPMneEWr/Ih5BGP
RMw5wjXhwyEwYLwZ7M0KYMF6UU8nHN+TO8dCHUKH6eXBUURAHAWbRLdIyjFchhgJ
vEbVtkD7goKCrq0RDmnZcFnLhMq6389rRnu7F14UJP5VNBb2LeE6PTHAs5OdBczY
znOn/blZV9wM8odEhuGYMz+9fLP/3/RZihwV5BEXaQy8RwFeV6vIhp6EKcmS/JMo
sVLqYbocRiLNrINy4IhXm5GqctIOzL3wx8sRB7B2yaKgyzRGTAtoXrJXVGuzpFav
rnHR26djDG8HII1RNlmbEQHfMGUMHQYGNpMo3G2scXIDuHQzOwK3d/iRJYyBqCps
u0nJcbFDUnvzfJ2XtQXUJhm3t4u6Nzra42MaPV5BGKOYytIHqpBIsF3Jxa6ePHGN
ToOAoAj7fgpoqOVI59Ug+YuQUPSyNov1/P2JMtMgBeG5I4vEs2Iz9pZ7vInHexKm
7SOgB1OjhInd4y9sJBupnMiCiuTenjZF5JLakNnc6uJFqwrgqGpIfpCM+iRV7qW5
HgtCtqaw2gRvNPwAeaLvh0p7F1mjV7XjlIRn5jw56D1xbL7kSbDm6Wd3oH8Cy6xH
fp0xYkQyl2lZfrkf9qhYTMyN3WcprF2B898IWysgSeU6xHAV+UfWecVhI7BIi+s4
4oCpgGz020MicsVA2/zQk7ZaOMPWStM43H776iCM32ELKc+RK8esnsbVJ1orNs7m
JwBpRtvFnWi6XLPQXSsKufWwXabIlbPOEmj2EKyNXzknqt0pOU9t1m6UjS6obwU2
NLdTRyYK5qKxx5PJHQYFUi8yf8vk6jK3Tb6XGEAi5tfrQvAOvQdyCO1dILA8ujgb
fhS+nsUkpSvLPZoRHtZmkX8nVDAvMWKoVlS4BUP1bpmWSn1UWHfR++R/16XjVMmL
KDJY+1Jf4sJYBj5y3F4s5xvghQhnEioSTPUnVpURISVFOO5jg+dnVvWcsuCcdgia
aF6wHWa1zyFH7XjgHlDESJhTCnd8k+fONi6XdRfZQi8u15sP7bJZ2bpcQHrD8E1I
fxlK6/KOPB8xofntd35VnQxVkIIgq1i7VakDnDNmYPl7+O4INi/yqhqpEsihWOOC
v9mk/n8lKdPBUkyRhQbrJnHTZeFWpsBwFhA/C/pPgXMv0u3p4DsQwJp0Mm1A5vUc
NmC/V+OrUsGbImLuTsfGQDd7R7r6qWdlxX9Yms952Kb49uLGjz/eRvS2zeiGsVXZ
l59LeU7Ogx344Bb1iSmA8rtZuspIlPaliZmkeHOG587MnpU7c8aYLlV3W959nttP
KESQTA2gpe9NPHhjtIeFEISE2V6lZd5zbJAbI9A5i67rGOca3wbifC4UJOUAMhK+
We6z3GfGwcC9JXB6423CHiZg4ZWWz+425i8QimJC4eMV34DA/4/9K0MIUe8pIK1D
Fu3bwwlAMo9JJ/02cm2XjLDfxYPEsNA0Sxdv5IwOFJgw+dhN4y9ELfjgUMrMAPd0
OPrlpQUr8wZu8V6rRFRhjveVHB8zMG3BsgcKKX7MQMrRhmIWZbStdyPpQMlDAo3H
x21kl0bmF0HJVymU5PhsMdIr/298aP7duBR0oAg2aDTl8iUU8MhYyyc0u0EQawaF
RRaomNqgYItrLMwM8wn6spSpbk9OpuVsw20EZ/ABx6uFdEtNs4WD33guj8QKy+yA
4W9XRg4SldDKn4QFffCmTAqM/8sQaJryxCp0F6ev4CwRUZh8uG4+SOtA+TYs4236
qQiQHNX/VH7TFN1WKCNeTgoRB5x1tXBEhOQmxc80UZRm6A9vZ+Aqdap+2S1iVNfM
Ma8OUrHmuvNUSH2vwwcn3siuq+TO0pT2SqhiONnEB9z+FPG4jL+9QQH7QepFDyUd
DPVGNTgI3UC3nZKAy5XeUiROSmHNkNdZmJ2eB7yU8/nmuN4TiGsfqwQxQS/HkKe/
5V6MO/iOcdNRkmyQqM5sbfgEIVdFBBsTtpoJWeTueFA57aKCXr+8nGmGzu8gDFl4
ig6RJTu0pr/AbG1uNZtio8vYNfALjP0Dt713JdPyPTExJvOStZQhtgcf0rVMYxyZ
i/3FAPT4XwYxJQPRoBspBKurI2oHjhlVyr2xAzF9s53WxQg5jr/suALQZmQwUBH5
XS4AWQk9ZzgAvz6ASbBc+GduOJdYJlfQB81qkzqmLrsLRLmyh71YbQnvVls1zdKX
RFMAwE9dv7oX7Hv6LFpMOwn26XdHQmVJVw/zXlBzLhlhXZVqvktSdWlw6wSvhZgO
A3JV3BNe6l8gSyZeX8RE/7vdQ3PZLTLCiXZ2dxeNsToAS1DaawmpxG+5dL6FHTGr
Xe6jVcr/JoVFg7dB2MtW1fAe5Z827bKuci50Z05vYfML5dTqW7ccEqYba3xJY8D4
qxoNW7N4BpUw8z/vAwneveYzi9ZbIB/I222YC61kVl0tRtf7InYx2hPTICm81+y2
lBoHf7c52y0FqeBu5vPAVtSRWnqAGcVikbiwWgTXnq9dR5kLyFTApnbXTV7eL4Gi
ecGmQTH+7jePCQ/SQ9dFq5OqmVEGvR7Au+vjJbC/aBGQo2Mu7+IKRckj+moE9xRP
OqE6o4daePesMgC6/pZlqSfdfiHUwL9xN8B/ZU7oCM94WjUFacvnJlodZMf/5wub
a0TW+fvlDdLPy0Apfdo/Ge2iaBpSVzXRk0ZGq/SAzJonTt+XVblFb7WDQmPVVNZZ
wY+MO5k6tsIMjEVUG1ee13ADHx/SBJTphYNOEtq5YiJOv4zaTRh37l6GXAnI8gsL
UKWSIB3BpBg2R1WNpP6FHT2cUijO3wUx0POss5dTfp+2m+UpaOsqJ2S9zbMHRhXi
1OLiYPPt/Tospws4qwb0CrvFZIGFninJqJDtN0DZzHbIhAramUcT41u9Vo/rKwun
JknzDT9h6i5p5eVVMQ83xfaNc+NbBCIxLbU1ITmO81T0SxXpRej5ylR3e3drjwFF
0K/VuSu2/Fs/5jTlCCRDOiEy5qq4ZbR3OLBjJICiL8+cEVMrxCBJxtf5EZwVoWsC
aB45nzXEy71YImue3fb7BUde6GzPPjn/YEbiUxrsDkp9DATirASr9QTtKk5UOW13
lTpd2fPczM/Hbx3fiHysujwDSKm0UiWAbpbPNYr1D6Etgl1/8PFB3V1Qbe+la0Nl
SASxBqVlEliQTKeU1lQjtTOLoEajZLrOPl8BARif24AAVOvh9vRSTV0KQx+go9Oz
u9vRf4glHslDZ/71Z+ezJWKig6IOgHDG7z/sijywZDPCYuJfdmU6lo2c9sJJpGrN
tbA/IxCHHJu6CmLIt/Usa0NsxUzPH6dZiKtdNM/hi8Yx0/u+v6hjC3mYo5+YMn+z
dlrR/l60DPRJEMlN8Wcy4njkeDKCUmrjP9vTNGbGJKQFq2G+428Lxslx7B+ZbE9s
z0JW0KV1XvKnP/A0ty3RQBnnFLZ3YFrVXonNWtSpZMJfBW2rXRfdwDw8sgiWDw/b
7H3Ck6XvVGYdJ7EfpS0HARPuQEEGqjJ1nl1G8DsG5+naw67eek19ITEROU0D4uUg
Z+ZNKSFE6Bk5Xizw+afycWCESbwolsASEdF01oN7/lmLHaU6CLxncass0qNLoqIK
lPPaJFiUnc41cXleHkdQYpzIISJZVnCPvJ0Hlas0wcadX3IuRGPVvRvCtjl4BSSW
sZOJ67qsJHormhganunXKfP8dSVQ2PH8qwLG1q0cYx0PchUzUCBQVTyIAwZTNNyZ
DyOWpMsTMhReqNwW1sPK0IWmmOO5PqVzr+47+k+EJPlgOIWK9dUUkn905Iet3q98
gVvVNW0GUOpkuR/ydyADYRgtXRpRe0vnPm7YEyNKtxmoh+yOiUbOWlr9as1PXgar
zSwO+gt8mwXlDW2HApZ6GLgG9zXkytblZ2iy0qOu9DHcvs8TaPNPgzQep9Jk4VGU
yiaYQXv/Z0Dm7rWjqJ9hTT5R74zEmoaMahPnpR4yEZNIIgIhs9HwCvw4uZ45we/6
D9qDpSkYgi2pGTAN74OEx//uj6fsRIXdLn9/juVynMf/KbEUHf3SDTOLoqlJ6DJB
zvcuhAZqoo6xgdf1o29NSsjcwaC15GcntApKoGnM4aHO9EoGvaSuJyIUiKgupJEy
ONYXY+IfbduZ7vRYFmZ4qmQwcyh8Z+TRAnHRHRQdQc8fJFLO1cKrnTb6Qe25QgLe
kAMJtWdVPuUkOVElDAOIiJ2sSlHqI5puNAVc8hPTjPZXN9BOaRmjFLIOoj/kYh/I
+TLjNhvqhPOSksK/TMf7SVHXvkf1EveQ0BvnINx8w8JZJC1uRSKWPC/RLcJjcG2m
+NVN4UnpUHoC25cqzB6xfzD9eHazAtWYGYohlylVYrjLqZNyk4S930qiS//LNuCx
0q1W6uoNgYlciSmJINfQn+rb9WwL6YxvJIXydjnCClnvLfg3BXb9isUYmBIZxlwo
2jzyPHjmOefo95yBZyZj7BHiEMWOrKHJmrqdH8hBxPbq2ll1IGG8yZ7D9pELPFbi
eJpwqwvJ+msOgurxcMibOclyNL0vyaypq5SI8L8GwuYIDvx2dSBqWmGGlfqXpud5
1OF8Cp/aI/KwIfQ98rdt5FIZYMGq5zlO4x5eBEQgxBoatC6cZef74m3zpu+DLyQ5
Khvk8PkELMsmWL146p/jkdlUi473928vBtlFK7ZElDfs17+JDS61zMES+RPpJk8i
NCPiPhz/dV1rtrF+cFgLAa2ud/wdinEpOS3z9BOdLziy+7212R7n3MwKd8SSe1D/
ySZHmDr32d8RbNdSFYNYjg7Mjr3GM/Dy+TXIaIxqtEe74hCZ1Np5MVkH9snXEo0i
Eti1alWn8MZ/O0VBHJcy+O6BFSUPIKdJ11XCgKxAzmRa8qyDPhllIfyVpg1w0LXk
+20htCwJgLSRFJJrJFrZJeCbuUrhRPLGstR89gd4hLRs1s1Or0K2Exd5JHJUlHrd
K9SeLfITuKRAG2yEX6CbXX7vxfEZfyK8XBIvPlOtwQBfwd2q8PlQ88nsC3+5gpi+
F0kMwwuinlQhriIkVOGdwquErqgVhrfc+rIA5BEgp4w1MZO5TJx+ww81StRmXjhz
ST/izEwkHfbeBrL3AdUsrM054ga9pc4IN2vyOu2IFfG7OM/9nZ7May9SkHJM0Bac
8NWmqIajtDs2qHKI6SWalQAyzbS6GtawXmwaENWpnhfJ3lDveCqvi3Pq3TZvV3AB
LX4dYrsOrTFnXSYaR7srFyIpaSgOqujEeZUNV+tZ9ilFYDYpBHQIej3hh3tgezqp
+2hLR/2imk244+eb1YbVHh4a5ZpsVQ7BLFX3QdeeSqimOZsVDyJaBs11Gu86CGu3
GB9Ca7XN+DCiok1ZG5Um82ZRkALhg1K6014CnEnhFM9cXaMURQ0griDBZhKoGMtY
2Cj7DqSfiLDBJKm6FdgN7NH+4HjCy4Ff2+3WMPAL9pJpt/scafvdthTZoS/azIyr
7fAGVzpz7OTwWBARdcLCki/mTDg6TN3052smuO+/77GbZExdh8pLdN4cA4YOss6f
OT9qouKI6BDByDCryrk+7na9qYgdkvrBP2Jwsr+1OIqDv8Py3DmdhPab/waTB6O7
JAvXetEK4FbiiG5EviNX0Emf0r6KReQ0C/cmspp2MeyO0vBxN9QmQm68f9/e9tCL
0tT4IJWMaoSad50ok6Dqq4+GQ2HcqnTqTjFbV7pKz9nwskAZ0bLYP1o9OKMouchJ
ByjXn1lvOfV/ub9BPQO/AFXyb/1E/CDIml2KJA+6rDacdzQj0lzNM8Qo8CRDYpJm
aomcbjqFL0sDsXdfvDoAO5+rIn+ZA76V1e4EpWHr0s6JeK1NbLC0C4U8p2pBhLKK
yj1kXl6KYY/VplLg5rZEYtJAyzjqgumFiaIfyKbNdxivu6DqjZxGvHGDRXQq1sqP
JsgqAD2DOqesqoUlzBIhPHD02V9Ikyy0NqM/l0+rYvw6IEQx9Gp+ZB+dgPeBbC0x
Q1p3bPrhZg7hXEUcLR+v306LGWinK2c46J+XhAkvah+52bKlZ2HixZ5FP2b/KgYs
sh9T5ys1Cem+JkU/eVtuCWc1wEJraQ11fSSHdXOm9p5ERm1AZU1x6bhF0Dx1W9tK
ontet7bCjlRNusahuIpnSxqfkxxtTwHiPgzHFuFREbNkjS3wR+IqyTZkYfRG6J1C
ocb8580e546cV5Ps1VYXrOreh6xgHI49B0wz84GoP+3Os5HrTaupF9L5Ug56auP2
i3oNUvVLab/XpgPwiOygOBbCJ3mtlQSI8daZEj1a1eX+Y5UQ1eWZffBesTIxs08F
+bnr2gohwEX46fqC5KKqSmjtiPdtIaupe5Zn8LUxBDRi+D3E8X/IpDSHrfz39Qik
Gf/UPHb6c9OzoJGi4sm2erzA/UGFn0LvobR8DjX9ThinNe1HWm0xwaOBowOa+S5x
LM3gPag+p5vrkxxic985vGiDNp9+gde7JJj9kVYrcq+p7kcFUh0GsyrZWHtPOzy3
DjswMoregiXmdPxs6rMHqh8oqg5Jid0t3WHQ9q2ESQZ0udKkubVYZb2Ovkrydoay
KSAUwi5j89o1rLYz/NXKwvYvzq3mLe+qhTa0lophwQlGAEafye2Qp6C2/XKI9SM1
QscN027NoBN1HvopPOVrlDqDOfU7nCr1+PKGApQOpCqTW4fQldmk5kmpxZDqdMlb
OspKknxiyJ6x6ruww7miQ6b+hm8SW6bFGrWO0GeL9dydmwKvqG3eeHKnxIUMnWUY
4EkLAlis5I4mv3uxovwIlrNuLBQkG+VcxYQ0BC73A4Fm25hRMIKav5kcY+minapb
3ZTBK5mGW07vR0s0e62piAzTzhqBUStBgCM+dp2EkAcK1HsDU5QFPId08eYs5E05
VMdLh/jGca8sjsgoh8CT2c2eBSvqzNY69IcSCottaMkQiye5ahplqDrXjmt0snyV
XuT3bXp4sA5H1ub0thFIZoiZ4BnqDiZ0eIXbu5TR0M9mpTIOHzddjvKdtaRJBZjk
Iu4+OUWYCXL29b0k3oRl8IH9K1DunOcdvnjQOuyp4Ao8frr3HJpjR1Bfm6pq/FOq
Psc7RXikoPEJWOxq2e4d9Mw9pOJj371M8GshIQSFJA+rZBj8S58PQUjZug0VJcZx
4MEnIczlgeCzu5SqzO6nLcouIHtD38zrck3R12vpAUS4zWGnwbSeRF16Cw0ZDYPS
rCVqsnxiaT7PaW0Lntxissh6NFStpmx6FDIYQCSEmZmAHkmJsM6ePSVyWJ0EQPLR
qqbSEWbokpJWtZx1iLM/C9pC6VmyzE8FlsvukZ+l20tDP9CcP53SPSk0tXITI9TD
v2948iWlBhTRaOetA+ZXco0rORG5P/T3S0bpQd4cIs1xX98a4CDogmAMET0l1tS2
J69VJKJznVqczF1cM50m+WT9soqdPhkR1fiiM7mOy7hFU7epzm+JwyPfRx9d0tjF
L1e7rFh8rZiJvcRkDyel/vYkMPWYY1PoNeXEuo4+BflVNMDkFoIx4FRFKrv8zKev
E3Ua3HtIkcWIeJgsh02+MJ+uaWOSzNIKcBuuntprzdNOmADw+u3CkIBiLn3l7AV5
AXetV7KE61yB7R0lh6OyebAetGc73uxgsh3EVH88kSgcdnm0PfHmTXKv53OEq3Vm
2dF3VvoLv3PiVFQRiFObPi+AGHP+8tqcGdq6lrOkCms8RP3zVe1dw4PkmP+tognk
26qgm830t7ChWe2gneJQCPTrSmdgGnrsvfH3yZbjPx0btIDeusDdiRaovsqitfZU
2XXvax3y/fynOxKo+SN5tLSwpJuzovEJK+LY/BbLAPC7F8RaZR+DwjLlf+0/99wr
SYIwg376ASl5cgx+T6ZGNeyCmxZu7cRhGx7C/TzzvqsNUc+WhEFTm0NRJ48bOGcz
rK2eaq4xPC+lOXf0SeYJFKbI3ppy8G/pKmesYzoOUxkTFFvcxTWt3UFxfbS7GC82
uDFsDq0wuYgdsyXa6PvD7+rB9GzeEEj1jpFyYZlHyGm0wszOXJmLp7odem5APl83
Gh8Ilh4abVkPTsMX0MwWwSUieM6AxiItwH5xA6SFByc6tMgRUUdVfEsOoIgFLkKX
OtLz3U4NturQaT+3Npl6Vpz6SjJHfY24P/7HT1ATNsA9/C2erQeU+wviQQ9+Lcwq
L8xRR1+csh7RXUKYFx5uzDAgkGpdjMf2+hd7Wqr3CfzkupiSLI2AZ6I2jznLjh21
JCTDSAPR5JySSjRleJj81ULBLX+WCUSTgPVDd0ON38j01ZFR+8dnJX21/rPsBNDl
3JEiFzVMDuNR/wlaI1WqGNBKOgSgS88kDaVcp56LcrvPgZDFPPNCQOYpvMhI7t8t
RipgOJm6oLUqAXaK3iJtuCIhPw2RZk4z/4svMq5zJoQ5OqtB+NXY6oI+ZvAQzyaE
tKH5WmLZOU5KH+MLe/WAIVRXzfNtS0x8enUxI64NLIsFMcXxOs+VkH0Pxm3zPJhE
SoU2SgA2nWZdQsq4dvISKjZbjtmDcgua9I5pvEBsZucaiFbc0v2/8YUwL6ih2YW9
Bcn7bzidCn6LdGDtGtsDL2F7jv0bEk0KxeAM7th/MCIy7ONkyG0lis67tIIQ/d6X
gdN3BLMUUelymA9YduJ6fOZzqnAnZ5fD/w7YmnLeIc3vDGeAd3+aAqARdDNLeEK0
5358AWg2e2wUhrBTOTVjdXbeZAhpgdCRXn9WzrDgWwxx9ywq84gkPdvP/waWqcGB
0mNdTJI3uDjP8yripVe7yh5Nz0wK/h0tjuVxLcu6OD8fuVvnFq43lcMwH81dBa35
zWSUZi+pCHH3Wdc3hT7X6pnNGlmBlIsKdqLtSGszGZkIEiKYS0PF1SqgVL5aVwC1
D99rG37sMmcA+KhsHXxsppiFg1tGrtCVVXapX7Q3fhBIPmhF0hawcF0Qj1tGysFN
S2igxkgu9F9CX63Z5vjI4axSYHc0Qx5Zff/IrMtwfcskgXfjshV4nMGZmdgnTcXS
ROyxpG4y1BwMbOLwWZELNBGJbVH2+kBOv1uqsB5dx1cbppZNdagvpfE11ZDAXcU9
C0WJeuiavYkXLld4MFn7o74R3E8Gl/wo07vzMSVg+vDGnvUw1x4TPQ2VwbH+UfGN
Rdi8NoFfclRqB0OrxxDQU6OTns9u7wb8o+jgmn29CgyOCLhZmq12tUfeQnPJIYO2
QloTj4XEPESHh3mwEe9+TygOlU9psMGZFo8Ukp/NiMcqexiAqUHU57KISRTHQeUE
h7ofJE0n8/XwYwqEKmpF01IfRHhGSotPeZ8JjzCxqz5sjISgKSsgvu87ES8a2Ivr
i6sBMQqCyL4DgH7wlDJN1HFzP7Yu6F/FczvNt3Jgmb0EhvpTCvR3883uxue0ywKh
I+e3qgYnuWWt/zgtALsuMh0krhF2DrFKU3an9nFfuPUJGVvAoXRg9l617+Su+Z1R
Jd3j9adCioMjZpHzzqRw5kkji7dwAHp+jiCjtUHBYb94WRZzEfy5VJtEoVn458hH
zuRKG0SrSWvlVjXtvemE4pRv0yIvn3DGTNz1mnqtOi+ohDJ0dn2aZ+0oHKnMcjYC
cQwK8W601Mh3jlKs4Ygt/MWTrW8Lqgf6rTFpOXPkZkNsIHmZ+D7Kgl+Vr7qO+S9k
IPo8halhUgma+YFvQYRXGai2ur2W07P1/4zSyK05NpTshiqYI7BA5iqULyj9TkRU
3GUEwbEEpPpOFXIlt4ldbCvIdoaAVuL+4+aJ0bfbLXzow/CfNRFbuB0zxstmpd9w
4N/wnaANLS1oMiaezRqnaUM4X2zECRb1y0AeOvVXBJK550B4lW+hcoMHc6Doie3E
4vvlMKZ6GRSjiQavzRaRlT7tscVLVx88sCYDfE2RPMGmKgbuaR2jZqVVLdgwbMen
V1qcRgPspTww/VSOmZodN+ToJykGe6ormqvSiKR/R0jKM9saYaETiQPWkq5E5k1O
fkx4lZOSU1rUV0WoEkI3Ot5CCyTyutCNUsT3dFMjK5DfNuh4NkCgjpDyromN0091
30wFr6yVdAN0gGabJRv8+TVWedSoDHZ+rYhl8dSOgtS0444rBEtO+rHOhrtOHwHz
QF4aq4sUkxyd+wN6uStJFeg6kZsWm46p/NQl2yuRraN78xH/Nh4tkuYczi1YGCxE
ZUI5GgrwGXnUA3JBNpRFJeFGWUIGab4nRBvrSvAmVpYquEJAOT/2wY5PiyFh5RsU
JdYw0iV7wQ7x8kBCivA2Hj+ll0eZIg5C8Bid2O1D1M1tw/Goem55wbc8Q4NKDFuc
o7BJRV1t7QdZRw5ea1evUnZKC5kk4JGQONIPMc4/rniaSt4H2MhZWNfyeZWz3Baq
sbAkDhmyvVI+IT6AWKEiYFpUjTrSdC2hqBCZ+a/anaDej2vDEmKcbLg2qE+47If5
JFCaRbfMH7inMkXmmUAFGzm/eZ0A/8e6cKN8LOTUx2ZRLxFkFj7nTJI30zIby9Gh
t2Wxve2sdK6vCU13fVPMqi05VNI8NiPgO1vFSGsuTUBSdAwbuaEnkkg0QUgY+5Zu
EQ0fyWk2XONzRKSlXItbWB9t7fL8sWuzkMshZJssXdXMS76/fvdAZnxEBPrI9bxL
nbdH+R5aUyND/w5DKy5BJCfvUi9jSf5PYdXws/r3rBnTVzliUQgTsXc3uRjZbv24
ytzf4lXjI42uCVpHpA/f4idReLCA3TiIw/Yw6tDn3WiQae7pk3AxlWP8+YqK5VEn
g2sZMnOp6TO6ig6L6cb8Pvr10Ouev4AubyLJ3US0pPPeziBP8bGnOm9365WX2uYk
wJLl2GLrYEgxdCNFTxiXhSzRsMXhaWHlLGcVEEUBHt6dXhvAOUAO161lEl2r0KK9
jJ6eybYSXsl5nYtgmSs4Q+yMbw2LR7Z8XbkAOIgT8W+ZuWM/o/juA2utyx77/eT5
owgjxx7Bl3YpMv/m2VkSpc6GnCAGeGn/hFUnvM47xIAR3Rr7GjTIopHWyyhDTrKo
30xXDYZ0mcPxmB80qK7IqD+/H5jgzTuF2mU18QvWgEFHWRw/7oNk/zzcGutcqmYm
FDG2tzUa8aOvq1EGF80knDaZVFuU9QUnEbs3J9o72zS/Qh/iDHRIA4pMiAFkP7Vm
oCHdPXIwkC77t7Vlwc38hQasER5dDDkYme39W2uXXNGtV3z1HvjX2RtM1NxmFehA
5Kb7uCgTGx4jF+xrq9Tc0TY6maM1ZXQEg0QanjNmWfgQPVx+lSQqGbYqoeb2ENXP
B50UTgCcrzBGeyeLXwFdx4Is+72+V4dZxkcTbtYEamI7QYd4upVzicvd281refk6
+L9aYp7ifmQk9kVPnTg5OAvmJ4Kdrjy8hT9dy3q2IghNFINdzLHKX+htO6fbsnXd
kELI0Y8ZjYfiUZT+zQ2f4CAvz2KNoVrEidrJwcMk/EIrbfwVnJLY7TrwaZ+Geb4o
ZyDQmiAkAkXKwjy93/DVqz0MOll34j6gxR2uJBa3/+l/rt71QuYlWT2i0SGnvbza
XljytiodHDMnnG/24mRSjdw36VoHDFNb9oBMaYVM22ow43cldbPsJjYYgTXaKzVP
RVGBalikRYWUGs9Z8vH54Jt3n0ihG52Mu9B/K1K4mUXOcDRKWaFdRbd6GtsueqWJ
5vjm2ze52/CAdwxmnGN6LhWsdUJcbrhU+yLpCIC6et/dW7Hw/WyA31OEV1c964em
yA+Yn1FQyY9Uld2UlawgDsJ4E/T+o/BCtEQDFci48fkKunn6xcfWJrNfdY5PYEeK
iVk0aLNvc5MHlPN4MJ1MiFLK8rZshx7j5hpSovG8TF2/zq7mVrElZKRDTgeMG7ml
w8wzK+HWSpbylFCtaCKzpc2bQUc3kn0aZhfB/N9oTnFQrVNbbQySMfRGOBAg0pAp
uwv/2sdgIVRg5r1E6cCA1jfgdoQ1Wu13LSql40O8UnS+2HZLFvVELc6BC5YT0UGI
17okXziGjc7Zb57uEMi7VeWeCTwIPKyAsr1BinZiqwMlzJZQyuq7UHtg49rm4p4q
JlGT/yFNyq3G0QPV1cC9k73Z+rVgaN038dXjAzhN1hQkoy7/jaOWZzU405LSY+wF
t1jzitEVcdEHDef3MIZ/HefQjPzPaOyotjhooZI7LTyWQjJXskSotyFktKBPTvGm
kIJMPwLBYrwDspatHkmiqwO+MpWnz2OUNQcRcbC4LV6quJWerhsCpaUCYwUDNusL
OR6/dmPD5GJnFnEvIGgoUqoFx8LXnAA7FxGWtsKJbUaQoQStopE1d+bmjM/jjFNH
615DvD2tXPTiQe/6/XQ+s9gUXXd3QVCwFanmTvLMrdquBqfkWElTK4mk94mCyY7T
k+D1QEUst7nDKh3HCiVUN5o0zgV6dbRthmgIFWBIHqA2pf2pLfJraQcickazeNT6
kgvljR6j1sMXOVKH/YIsjP//wxLJ6jn4SSd8j+FbfuuzOGng7qxX4yQjABk6S31q
8rZ6DfONg6KUmmOB/SqXFE4X8WXiN1HgOgXT0AKoCxAX565ie46+0pEAxUtDoZ3S
NqVL3456oemKTCjgvZRkaW3hvgb48naQmIX8OH8tMTOYcwUoAHL+obTzkfidYfM4
Tl3QDx4tnRASN+jdXEsVAoixOlFEx0sqm2pdU/l0ivNxstafqSxYx5M6b7e0/k0C
KOPLdNP6nUPFA2qKXZdIxtoDjjk1wrry1xw4pu8cMzS6m0wiVI8boa0HlfbWIKtr
7/qm9ke+lO/McYK5dtUp5g0AdhrpY6+zRk6++kpMV82GqBOeMJ3c9hiWnWJeL+JA
WHkszmKaDbhW+ZNhL40xEnoAQisG34Tj1nE2QJxrOyjHQvPozu3aKrh+E2lhuhAo
Cz+JRgmC5806454TfZAz6WUGXPCJQ6kJQkUvEhjnKuegIKECnpaErpG3iWKP+0CG
poV8tQ7BhrLejpAhY4IfeP5u1zWDC2diJhGbWNh+dZ17C57XXXV5cNNQ3V5i9Bcu
pwemBWdxVaKVyfHVA3FzcxD6X2pL6+Qgsp+1Ksg1hZGehgBPlTI7ZU5ohJopZUsp
n3Yl8F9CGaTYdrGbPEpIUgrp1LPR6t4BAfofqfK9EVrJLuZ0AtcokpCFGCAvHSOC
6J70E5rXn6qNaFOCHfSZLm67xEvjqra3Y16vlcQjzYu3NH8KnOLCfCq7rXCjSfqW
IUzJhTi+yHHna/aYQDaCsT9ms1FekWcCAZ0Z1Hgr7MehIW6q/XOO3o9b+JfRteSO
GqotuGvVDH56Q2rULM/sBj4Ai7vFMJtThj25raKH3uPUJpwNYD+Kfeuo152deZ33
kCE7sJoQvIiyimfaaKl41KQGU1Wf9rapIOmm824f+bRP0rRJNetjnRBqWgkshlQ4
hswhNU4vCLXR6vYtX3U1g/Ww2EIDmrLYA3rvv24+JhEh4vgR3FLusYnY1o4fGApP
/bBkGGYGWEYjY1BlkAEVEKHWnfiqQGSt88navO3BmbLtqjlBWVOova7KrV3hHOuS
5R9GJ3coaa/KVpr9IAHPIsRYnFQCtr8ZhZcEsEDwIc5aYBrSx+HTcsEw16Lkz2Lo
2cEeRK1apiQ+NhiunCHBuhD5Euiv5cIUZvlE74D4GNN7t3puoAXjJB4TZXsadnFB
yKFtUIeyccg6AkJogMROhIBXcLeLTXoS40HSDMmuqzkQRi57bbuRtq2a2x8sVZxg
2NvbeD1tbr3bF6w457NNLJVBrtC+MAyDhSYO1RL+CyI+AM2vxxDVGng6TNff7KMF
Qsl/JL/o5AFKA6ATc+KE67PeSholzbQeHuM4gzHgab/RlzAAvFSK1w+ge80lrIYs
5A4lorPRI/nvVfZ392gpPJxOH7b0hAAIDuWqDCAElctC1widNTLC37ubPACjYA7M
uIFUyE6Gw+yGbRg4L0p28zTrF+2Nex/txIR0WtlkaS9G0AiCQs57z+aH8Qt97MDG
3J3Egv37GIOxG+RLWNBppsNg5j/L+I562YGo533D2xtN0jQ9L7MS8upgjzVkpe2a
ug56TwIRPQMLunHp11CoM/vLG/3bqXR4he8/hsdMbGpW1gn4xVi9R8MERikhHqxe
5Ja5hNDY+qsZRSv3QemeSYxLsd+dMG9CghmfyNEelTod7up9rU4pjPP8t6PKW4j7
AK2dvxpxr2p/v9uDWBPzepsejD2ND3JVLC1nZ4e+H4/pv0b9v8oJuFGloKrOOP9p
+8FNIgtrFiMeCA+kH5A2TGiwjwTmYwd9uYdNU4zpHGC2+2+9SgkxzTjr09U3dPkF
hNnnLDdu7zozDYRnzYJWafGBT3NGTWJugd5IM0a9F/XJG++ADdPRVthFCM5QMaER
1ObqaSWyWq1U43G93e/7XEI3FA9ZmX97SvQd4MphaL0xW+YAjf7jSTg+9oeq4Xg7
vwMhbDZXNMK/x3wN+WvsHSXK6qUA04xCHhbgBiLe8Jjpn74uosI2mvtNPOFjU2ep
gtbVLhq4+ABGw1xP2GFEkUhzCP60bdztv7JvTClQu6ZPPYvZdqqC9dmwJQ5zC3/3
CgjHjVr5N5qm9vVNg0pwWgUShDYhVkg+KdLuqVcgwvM6D3FtkvDZhXIv7dc49nSW
tox9vOOwCwokRdyoo4tMuDVHtzGzgFIp7BdjD70zFJNewZACDE9ep0Zm/IKWYwub
BtCxdCJmh078v8bFG2Pxb1tarIR2GkUp6kyRtUlF75pWXZUDm7jIqvfWxIHsKwPd
gPNq0rjRPPr53kfgjJ2cndhAZVzM+8taQRhLYFJSln5KgvGCE4qVBWCdHYAaF7qs
+1ZpPkCbFP47NndrkNpAOT8N3ZgCXbFuwqiHPEvVUEJUXIdlz/P89qXZi7ob63XA
pxzdyOMz+bhOGdu+A3/FxpCx2gwlB09DBTZnvExFtXRLYpfUDA8teB/De2ugalxp
hBrqoCHUId9Q0yGNMWy7Zyk6PT4pKjMww2t5Ru6EpPLe0+6KdSDvqfJYtjYCXB74
kfhhy9ebrhBAn6JMngOFSUQsw1+xOL/x+EzIspOnjtl4AJxXLeqGy/dcblbzqYZY
XnPP4em+Nx/4MMun9VQssLdeclAjDlsYS40lZB++hJ4HweyIeHd0pthJYmoEJr6F
2ebJe9qoZq9HklD7M8PhwcPPqyGjN31jb8UWdMuUPUsnxbjnvUjMUJl3JXrkTxjs
ARqdcT93/JUOEankwHbOVPLKkDwYKeXS9KE0gJMoXSLzzEplXcuTyykXDruEyReh
7doT7k043Eb6sIzX8vvbmkKetl5W016R1Oz7DWi87F1JTK37X6xQtXZwpE0iJkWt
sPgPoKmls47IovZlNp78zIIFJiuopeS6YgnzZQzaGpZ1OWhzv4CSxMofhhKHZ/Cd
rKPWanYPeG98Hut9TVUFSxyoeWBNQCw8OI5IJOM4WRHXIMxKegUQyoJHjspwX5nq
Tq16SsnGda2Xi5HYekG4I0lYeG3pzt38m0cMru+zeQ1j44MgE3ecEWD5Ar1liZPe
GdcSxIWxQEuh1AN2KDIw1Zyokiz9bs7SJyJrN4LpK9g2k4jpVd7W4+Tc/A+7pbsd
FDIVima/rXxX/Fp82/DcGGfGF/kAJzFYE8lBAU9QQcrcoYnTebzfiBZF0XzjDdkj
KpGKgh9nfNDKnKCzk8UP/WlDva1TXw4tMIUXhWPL2l3jx6a62LFeskwU6jB3+S92
Y62JCPYBUWTR8h4NSBUarbXCc6iIBrZQdKXsnQGzsbHp3/nzqoYy4iLIXKhQEaHn
1o4PfK6j9M5me/9Chwq0niR7qnss2W2OsrQerYKkrrkk5VzdRw/pffrXk4QGEtAj
EMWpABu83nWRMGzjqo2+LPN91vo8ug726OMJKJQBfs/ddzzAI4dxgMWhj8S4BvbM
rNWVbE8a8Z29FRBJ9x3bWpFuuGk5H3/DvOUJcrsE0rO97SeVHJtkBcsXOSpFhjP7
0bzzpFMeq73a4/RLtS4ff3L1QlZvuVGfhktGchCC73QGPJvhjBuA4hm0OAZfvpsV
FMJT8jDJpM5NyRXS+Z4i9MpEDPKTw6zUL2g2oqFOOi9WocE0uf9eQl6XX3GK42dx
4Vmt74JY4ygwxAZxovYuXxsOWGqCCvtkh4UpTxDRarirN0VswkdK8xVq/mMAc5j4
mfso3Z0sDzpvdrhb+ES2pwuXhkBj9zzRRwk099j6FteIy38ms9cQHj98+9XyMSJG
zyM6HWP/q1sBdS2lOTnxbelxgStf/ECDPHWvDcEmyzyJNONy6/Jqi+66XhDu5hrd
qgd/7GU/zWyDXlSGGnsGjp6/z4uqbinnpgTRcMpkD6TDkJKrUm3bkPhbJH8hK5u/
R2FXTE/CTaJJdaBlDQOoh6ws4ZLzqB+lxhbueWm29NV4OOD3buyIKb9EoVlKnVs0
t4/HV7HYhhM6rCKFhlj9HGnCrRjK2MKUMJW4NRARieB4x7So/0G7SQoxkLUTAkQ8
N4QRjij2oe2WbUhLkURkRY2pH2HMYXLFeBjf00pyobhb/bu8iZn4ndYxgSt8Qg+J
Qt/E/H3RB7g5tp7wu+ux9ExWf66N3JK+GDgFkJVWsqL7JQopPe4HXHExbv80XdKf
AM3s6dMmXF3E0oHqHAKVryACF/xqkDShMzu9B0ttdfohqfk9jdhBIBUZD3AlcCRq
66u9kcBUIWf8twj2w0yNpRuae4K18ZDpptJNExLJ+IsYsM+Mv20aB0vpVzdegamV
2u1Yw8AQfLx7F97iryI/+jJU3B1b8gOZM1OiMJXCr2CWlfXWS/3dPTVVxEGLq+c1
cbYK9n7fDZhyoj2QLBvC181+iB262YVy6RsKOpHkgHbzXpI+asBPCf2KdE6cOud+
Ya2LDov+4OJXlxbiJaj5jUmJoBaye6xQQgyaeCFSojO32haFNv5NxOqHjE0xGyZ9
tZpOwgWbwXw3dBjqZBdRheYBUjs3kJai03n0diPTAgDhX3a1VxmyxhhY53oVbffm
/HX2KAehDbkmrpPCp+5OUgwKmU1Iz/lSNLtr2HwHNAbbHELv6n5RU9yvsXN6iVgb
tXhpY6oJffStlGR3E9PWKI4H3T9d9Hmh7f3gRy1YOMrqWjMIpR0WvMnFxl5UYRXn
Xzcvv9RN7DVEdRYEdS+JxSLUgJEmyEukTv5xAsmvzUmKUCh4lHvn4bqk207RuEAU
LQ07Q1wrWYAmWPf2RTi0ec6hvF3SNd8KSe85Sfg+ELC97nucHoNiMDIBewsiviYY
7x/i7G+gDo8mzgmGVqAj4WDIzec0Lw3HvEx0fINRzdjxwpvM6qWFOIe+U/YHkrd6
MewjAGWFidbVS5KPcThrS4AXfN2fdsk8kGla6QMEJ0FdmSmVOYzsOzs8bJaiYaz8
LCXXSr6wsfU+kJDvMN/2IcPFpkTSQ/8h7LrLp5VNgqqwppZBX2W5PSB1bvc9YTiq
Mi0GwkVWDe1K8tognvT1JyZBm+a0XqSfCbjMFww2fsxIpOFW1/uM84LFqpq89fzQ
D/XdOT3kIJvx0xkGKwSacA6qVvGk6z6TgnJOnvRPKW54eFEdbOxKsV3Dkufk4VYn
qtCwzAtt7ud9JUC7sVyn/N8H7OLRLwSMOJMSiTUc5yZ9bTSByxIZCMYjc7IsZ9uB
Pplc0duyym6No498A1G2sVR5NC3mEB6xOtBwCJNHGjP5W39CkO1y60tRWjvsTppV
hvCii9iZr580bjn31Jhko7qAXUQ35hZESJJ/idU26rIA7ODYOqCm6y+F++ALcqja
zbcGZkMnjQpC0DRRPJe14mu7F2RkO1Ysb4AH52Cbfq1uzdGms6hNgoWA/j5R/fTj
GtTUEDDMXE9/S0TwXzwUSVWPIQ91/GLyPODr5qV4agNyDdIqcE0xAPKr8wuhDaDD
c1AWGX3iAiywk58X9xNdhwKk95v0NRE5sk0ANCscufyNXvN6LxpwhhDTs+hKb8ht
gdVAA5BGEza9/7SV6y5HtPcjgZxwhcsL+/oaqPyy9VqwzV3sU3YH1ZlrSJy4QsCO
3TyBHJZDisP167YrYQtcPcdGF8dvQu0SVw4Sh5Z8ouSqTWcNe5UU6UD0q7pqfudE
Cr5qmtmz25HPSpTpC424QeFjBRvJjs4pEfybZGgL6QMdxkDv5lcR9rxln6GdK4Wd
fxbOSIqOH+Wcrang75IPduH6+qQEcGzioyc58qbevxaMJxwyoDH6ymmdgtyTzitS
5SDZy+uBbGysZVvS2LRDrlnnudSPPSXjhC4JJGPd0BWSNpqsIb9ofrorZyIuXYYD
4Jfz6N7CbYgJWZeLgCrFdOR3Vva76qqSp/pGsdT5wSIL1NRwAcE7LhFAfki3VOxg
eRmhwbfiQB3oQBxoJzYfXYIaTci7r5RA14koUDgpXTp6CwraDxOAdZbUQQIT4mML
zUe/QuJx1A1GOpwcQTFKRYzURgr3qISs0ktg50uyhuu8lZ7qlY4j4lJs08SkL43g
lcqjfdNWApSdpCJLGyg3xRah6lfkqP3YEfOAnzFaSJ5q1fGrZpOKVmEkbQg5f9ZK
pEa1eDvz7UIJb1dVy9MyuZcQJNTHmo2KPsQBoJ9iNji6KtHiHySSGz8Dynjl5fdR
IjdvLj3z6px26CpRF56QidZ1aErX8+gyGiTnlxVbY5trblJvMkzOvaMIPrDHeHP5
qm4yZRUD3oLe4NkVUgHn3XRaf1OjTjvnXItrIqlJ/3WhpaBvLTD29qFN02RtJZHL
kk52VQulIesdvFaz8cI20ibpxx5oKpZM4fFdyI6lp/m/Xj4Ag74A+uaBl1QJoZwd
QlTAGWNVFSj5zSCFww4E8h4sjpCQh5B/4QY2ytHSrKB7B7HURcvhCqXsQD1t5gKU
AOBtQg6jNzJoEeaeuRilUMabLUEuC1qwXF9Uy/9ytsknUMH/jXA48w4y5uIaYt1v
iuVyBhW7fYtW9O2RXOYD0+rN/YTwaqVPOohD1QUWS4/bysBb2qzaZdOxSpdSpqsd
RFvlUyFtDCoRbnJq2ke8lp72tHBqs72bN+TuNDMWspWA0LBODLaFU1a/XbIvWuIR
ZOouVJE18R1nw7Mlp3Dg8EUs5KZCn6kSdODWWO1HGS5MShibh4pG7IKnhi1kCwc5
KCIPOMKgcnLaQKxOvJBBYF9wQkELrbR86IO/R7eJBts2AQjTj6Y0RFyQJw8FXyDB
uRvOPCl43ncyoRlPUXz7ZFQz0vd06bmomrsldZkqTDU7T435TNsXxUbCFvOT61YQ
o31jW7MQizwKU9Ne8+hHbmigFRYLDEVS8okLtddTypSkADt/VulTfYlmcVRtYBUX
ho1JuZ4AEE/a95m4BITEbT9g74snikRT6LDHok4Tc97CzBu7r9yAN6Loaw/VbTY3
eg/OJtS+Y6tJgY7FrJOBMCvfVLr0aVcp6LtCoICvjW75J3Z6hVrxaevXbjuUDFz5
awuSP2rf1Yhfxy3TpKqlFAfyuBJJRvWWFtHTbSqvLtzwwObnLI4Hi+p2wteZ13wZ
Jp9SfVn4+5f4m5zyWSPNjVzdeT390o3/hn4lYq5Y5Fqv9V3Dvfk2bszTmIXAhmW2
/CgR4R4cWXvWAAeM1xTtZCCvRjOaF8PHL0wRkXekAtHz68MrqknvH8Bce9xBUf9L
SI3IrJ/y/5UHeFxjpuO3JH4kaBj7w1kQNI+W1uXCIl+nYXqbfOJaucxjvPM86C6T
HypazG4FfcVM25UzjGQXNy4ic+Q8q0iKvk7bU3u28/wNfEnnK5Ufq26Pd2yMLB7c
okJ64rhcvcJYc6v+uuY5cr5kUyFswuDalo87eaqt8/0z0BXXnPggsd8lTeoX4LYg
aVke+6ultcV662WfLw1IbrEch2QHVNWKxCRbFUHpvIPYwTUipCakgcqn0K4A3lX7
UX/IaSxOFmuGG4QRgWOO3ocTJfgBt5FA69Xysn/2yLa0eQ7VzFyoBvuuzj22XbkH
pQWX0M13rGtLlyn1pfQnJJcrTdlTHK58TYFZ/JXz06BnwUolfWSHUqeFdNOm6weK
NwkvVaGovOpyyea2wFJFrUoKD4hqxtlD/se+E0c6DtogDY0GdLbMNyxCCtZ9yLER
XVtzbNjkLTR+9jD12C0XOPzAlw4sK0C4glonbndpRSfDGFQRgKJcbZTxSWEVz7gv
Ep+G9kzfMcUXHsB3i0U5Z8uyL7mRVpF0IhuLSyUeMkYNrI2gaDml/3d2G2BWwwUg
8JjYzKW9GJsznEGf42QaCztyqREiWZ1Qoutomer5I1NePd/SbLDNppl5psVLjlKo
7Qc+VWTmi5Dvp9SLCHueusgYlJTTAzjmzWD+fw3GsQ6MElhzN7j2qspNeTcqk5ss
ph2cbFD9sLiKYUXibNQQ05WBE52nTnqMP3nsEvegCVirbueN5gxRSwm2zNLM7q6y
U5yuJnyIZJo6dkFL4TgrjPx0PUuzqHuDRbq97K2Dc8VVsyj09892YQTeveIA5MEy
lGbFdVkjHZk+WM2EW4bW3SobPCmc3HCbYDVy0zR4IhioGgHWsyt5SexFrobLY/rG
bFfQlol93e0OZfP/pu3/4ZM9GWlcO4evUVQhCOCQi+BOCSv+CyJnJl3MJ8/be8k9
QCbFxtZWTwHgSdDCXPdraO7+69fSC1mvpE8/lUCQn9kdxSdklCje1FqUdjthddn5
8hwNTomCl7q9p1lKSowgCjxQDka6KVngFQP45bEgPkot8F63gkwbbWPQmGsPSAhe
rQKJB51oswni1YY3sPO3pc5xDQdl4kl+Kq5TEbwak7XeH2s6OSrsH2dlE+qpmyj6
JcAAmpZH20VxcI/jcHK3ooxQB66bgwPoQo5dbxr/QKosIGB0hSRI+wHMKtwx6V60
4qER2zuFcdtXbCIlkzxUzPOYQ08hw5V/lFhifMF/Y/NoOAjcL3BN4AWSHjKNFpb9
/pJxV7YgaHrItf3rGRcztwsWCM0zTSA9V/L3VeJiCmy8Dcz4LYQh+uG5nOy/M3S+
hupLwyHFPCLSRs4ikmk10NXy59pnXnXYqL/76GIvgHyUoFhCD0YfwQ3Irg+7uhMZ
tSUTvubE7yd5uu0weDvPnkZ63pILmvoOjyTh/gokWkL+YHi2laks8MNjdi+bkPcq
J+PDoN/MLAO7fWzbj6vpfon9hSHQjM6qHM63+u8f2ur6OfbQJeRrM4kQNFvzXaok
DPLrd2L4Z2G3O27Am1p2HtmoIzSEPxI1v8jp/bGdmvfXVHB6gUW5BEdfu+iMOCHB
yZaxw2VHC6bNX4lLY56JZENoMGIo2mlqoyyCtP40xnObILH3fh0++poAg6+e9RZQ
GbCd1IRaZnzHjuoqPs91zCqvaopkjfsUMgap92EuKDeQCEUN6j5wMdx5kBNA+Y9Z
MnVsF5l55CopjAvnithY4QE9rridLQe37srXxaWTIsMVWijDT5lelH/IlKjH/LUq
8qFQ0WbXac1yCObNMXQPNwuxrxFFOHqVkmAQ3yXfTone86MuMURPZm0sVzSDc5ZQ
3hzSc/O3WzBZMUo7YDIsGtzMv8ai7K676NHaIkbMpajmLUIIdROQRMSyVtLOdknw
NBJPrfzGnrLSZWYmCMsjUgqGgthOD+MH37b0lvqMABrkn29lh9BXH2qO2uLE45ME
rM9XeISMJPNPluJA9sy1l5nN4q/+Nw1zo3zphICDugg4BQP3H2o3ToNP+lTmYdzK
Lk5QtFI2MdfZ1GMkZYkaK4nySxX6BNyRuqVmlHj40WMqYXrxrSBgAxrPEqMMCYJx
lykSafenL8n8LZgSS3WWVgrxnS5RJFQDOVblp7KWHwl6PDW3BEHyk2jblJGQ78RH
/qIpWNYLQvKdEJQ9RnnhTOgEHvGzUcQwf6D2qcaWhnAem4utXf3hXZUUNHFor6sF
RaekAtHmwogHX8ArB2Kfzbwyr+y0emKTEdSpagR5pFnyV/bHfTTRv3ZBUCu+0QCq
UZqKQ+f1FVNxoCjZfX6yc5KFLrqpIWBwP1+B4hpTccBuoAuKCUNdGOJ+MVTfp4SL
Eox/ty3Z/4ltrq8+WUIMcwy4Ms13M2+tHXC6NyNtp7SssS24PHLuceDfA3nz62UM
1K44VfaU+11LhxKCCt0qWpUfyfosYb9Rff6aa2PoxKXcmCrY7ziCwqodYYX9rU/A
n3BRCwq0Xu7b/IXTaDinJ2x0szKzr7pWfo+Skcf7A7xgEpP4P/6gDiITH1y2M5gk
xusr23FtTB+leoR5vNppiu8Go1eYm5H+nd/F15IRMVCJo/xhMAeP7EkGxQqNUd/m
c2uLBq7p2s9BHnegADpgvR6G8LdCHJ0H/T0XWnjCMxMfuJqRBZddUmQXTlALq6Km
DZkhrJYXA9L/XgpJX7DNggQ4jh1m6jvZiZWb+upi+QNVDzrZn+jrrs03M1do/o+a
Rnp8VE4lh2ZVsDBCFMMd9tRvu/P6Gj6GTGFKM8/72DEdXO43xxquYjjZtRPbydIw
h01FhQ1EmSE6DicQT8E1wAPYtDxp9K+snAGden/5+wME0+xb4O5+eO+8EjDpKgR8
hnwxD3L9G5yEVnMpvHx1q4scyMPbZjKOXePDhbcKlsNqNbdb7DnRSUAPbvG84W/u
lthWWTkanXkUhqumg7xhWSySIIDc9nhPQUkxx9PrqezoeFfO7Ok5yOX9ntb0OiT2
LEItEyjLpOJwV5G0izCvPkv7AtUdlOUo43YONRZZRN0ZtxQaSVVn/F2e7Edwflo3
gilU1DPscto+ACGbRKmJ2Pkq79Vycj/bK2fqkZbmmWmelIKla1mentow3E1B6V5l
l95oPYPz41o8i3RY3pQwWv72HRNVxsO2LxaiIHqwnz+PqUVlESz62OO9upXUzjZu
mAEK04d9cQ/4AjlvFy9lLwfhGJZxi3UDO8+oME4f4LK6U5RH3TUawL+x9pcFd9H8
YxSuDnhYVv5i9SkMtEOvxDo2Xo1845wwi6Mya9kucP8tq++mPXVyf7Q8lES1be/3
iaSeULuGc105HvXFUzmfI1l2vAK1mCCJWQ1bewKEYkvmvg7IO6ZKSiYlmt/xPSdP
McBkCVGJhRq1ZXfm2lUnltt/JaJjy9wvTdjcd7UKVG1eVjOYQ4eEaDMDbMvVNSmo
GClgSai6Kb0uPKrz+fi38lIzHf49w+3oWP4gxGmYVF9ucZx66NxIi5pATcQ1/IO1
Cp/Quw7zfBSJEVaWbSRuraqfdaC5WxgOKhpiJGV+is0hG6rdREfhaP2Zai7p0uzr
FwuNTKKj7Rkq+ykLu4wCIV1IelEZNLHTEGKPp61XKGTABsrZTyL7JpitGaB06lPO
k1rHm0WkX9/vbQHdnIToj4HmgymHsZYQTxODVjwkE1fRlDKeRGVhVtiLOEvRPuei
khkmtiB9d9/nYjA2QMLjxozBAJTC4pwiBnAOKpE8mhAmQxUtHDm2SXT9oV19VOv7
7LWu9dthMi+XnXMZccoCaWZIGLypcQFblHqi+oFbNgrYEdTjbsQQBaDF3BXZqyay
LWfIZcwLDSIhCdEmZLfzfNu27Lz2riy34ueh8JraF1elEYz52pVUKDCcCY8KxTZq
Gh9CRuVlgz5keMK8CCvjeEy9OgHjnfbrQE782pe/OBMitvbaRNdDZVWjXhr7bCQ4
Z3eIx5Tr1EMR9/C9CtUjRAb3t1lxXt/C6u0UxM2kqhaeVulZfU2yawQ33/BilshI
rZdRe3FlxmG3Tax4ptwVVIvOTtriCnaO88YyrH4mOS6TXbUqMJStusNM7sCxCmRj
gfLqrGt/bx+CO04KyOBoDBRKJHqKPMZR60fC9Dc3QFhGdV1Jug6CeeCkyp75j/xN
iwCMRW6jBt09O09ITETH0MWpn3CiBmJBEDcwe9aQzGje8E3xc2+PsIWGxN6Ead5h
vrPSbpRtD/N5/MIUHTZwnTFR3Pc7jaBJiaxM+6uVF3r91E8JEixkr8zHyD6X8wMO
Vg0o/ce43Ps4ydhrvmD0ILZQLdK76KsUHb4Una8QLRwemwMBpGbWIy+U53cc3yIx
8Ot8YUyjLgNEkyfbPA2q6etsAH2LGJlbFJWmKnNbozsi2qK0bEBJos6tYiQwftWI
V2jApJcMpnW0jjaPuxLgiF/+LkUDJYaOMatGAx8u9dt5CP80JBuh5jdtl0Fpisyv
Mmfrv7VnxgpzZiQq8u4/tLLxXrSvMwiymm9i6Dmy+t3pi+GgK/51BS6KolERTbRo
jFFs5S3H70k/4y5Qb1ap+voNTE6UP/lm+RTBi/j7iMRpl+75KeWwSDm1Nrq1hFjG
v0fozLnum6yyOTkOjIfuVdXzIEI2hcgsZj5uECj57TaX0sSyxr0dMn4KCeRgiOX0
SY4mM34w2tPTI7BOxrZ360zdqzCMpohe4NzHSBNxH03Bkp9d3VN5XFbbUhRXzTIc
xZjaeoz6mo5jiieU7kpVVFDZvOy/PV1pXoREhQT2fmW5VOxn2KgqV+vQNo3LAGTY
BvXTzoIp2t0uUeu6btb8O5cD4Ig5/nBdVIZlJe3NCN6ZcsA3ELWTijh+B1FIfa+3
KeFlgKVrbZj+IdrRtmWakTbK5kHpG9nmVoBgAyoZXwdo/YZoUNblAQkGWoI7QenZ
AOzJR8zOvVTz8nCpViV7CefpII3o+YYL7GKNlm3OlL7cktCX3YIIW5/iyUrkKELV
l5kkKpfsc+WXOMcbsAehmmm1NZ8YWGMrRjv4bAwPmM8PyGYTa5eirLv+3pQRzTbY
N0cSkRpqyWLZUutAI7BTLV7h/tRSvoJQ2q/h68oEVASNPXNZ8UxDDBv8ZxGPal3X
/iRPYyxKqKidiTv2cdPhvPjnF0sVOpiFv9JjlV0ZIkntQ4SgGFpvgZy72ss2MaIM
w4Pxdjf1ggGGnFh09Nr9N04H96xrHEuw5Q/vWk/XuGNNZ07njlGIzwRVAhZhP7Op
x3bAbYxBtWGJa72SjKQvec0wZw2slcPh/SsBDGx7qiz5a8M+eCi8k2Sksn07qcZf
d1HNNV4rymKW3VgM0/t+KWN4/R3f5foNIivE91Xjtnd6+9ULCR0kjCekkaZlUvnE
qSGq8YpBA9R6EIwr5favk5wlxC/vY+x778OdVq4isclWh8yi/eqwlHm5jo/9SNQy
HHFesm/nfr0BWxg0zIdlsY3a2P8Q9RI1LjiQHoARuxAF5nZ1GisDyWyhYcq+eRHv
hG/amtPoc+3cXQVZ7TSPYr+ysReAJh8PWM+JD0PQq97vvdMXrJpI6/yuk5EfZj9K
BmNLnhhqLHUDY0V0/lYK6GyhrYJGSPwGMfD5nu8Ayfn6rHALOcda3JQ6cl68Ne4O
8HNPSknJDBoeh9OG+gidT2EIX9YDVIS5b/mgXR0RZfK/pDqAcxYEwKTBc1pTEUYf
dTYqw0vmazz/zVO716INRKSyg1XOLWSqQzLAAREbnrpQB0PcwhfXuxsfP4tLlgQg
01VT3+tndsGvWtBcScI88i8542BazlJE1rjCjVUQMMisoqUPN/ndSdosHWYY/wfy
CjJ/9I+Sguq2ME2ffK48MQX1aZXfSKNezk+g5Qmfju9jCcZ41e/wvw+olJCBX2gw
WsqLywDup9baRAwrgP3oNX2HSCEyLt26qDGzpkn1q4bXNSHcXVit45EWKwT5iJnt
JI2FJuYvNycTKGoqdhuCq1Zwyli3iQireS13TZPoqgZ6uWL21smxRAYks5WYGdyt
PAEUD6euhIvj0ZtNmq5QqpkJLYswr1xJ7vn8OBo0Rd6OKY3o0QEu9ghAAsea4I/O
TtX/a+QH7bYNa8GflUSeGGY5uZOUGI8ztsQaqbJViArJEAa3cp+qWuE7oJcXlCvH
vlXBLeKIKpbqmBv1yQMeVkVas1BcEwji0X4N1SakleLComoMtBPBWPsOGOmgeWaK
hQSpiJgOvvjKZrrYM6FqScorm6zwDYl1ypJyXr5kwY+8bHcw5DdPqaFOiignc3xf
dR4YUMw6AE0/e8lv9WibuZ/iDN5CO517NhXZVRu2iwJMSx8q5hD1VudwDqUj19cS
Jty78j9H2xTZZPEdNbV0kuKV5w79U8hofcrWrZfISs6w7g7FCKYen+LT3xwN9SYk
+CQ30yhzefDmheCd4WfsrLzq3Z5IufB8US8Dhw311uRI6BOKroq4Am4V7Ap5IGII
aP6WSMSXeC7cU+bhoDxum6M9Y5OHi0geFKRB3ENuCsnNxSspLJIz5wsKwX1Ou8gW
N/S4DgMNaKO12MjBuTT8HZN4zes/qNhEGURDZYhtG2pIQY2v9xxhXPTr+g7vLjjD
BAAPlPfcm6quX5Gu5vZXxY2CsiO3Db6ZzpdAEk+FQxcq354SvAPcAOhS2SZFmP7x
z9PSU7O0q4APtxhDa29tF2Ev8qUIWFaaD8Q+9f82w6jzOQt+5KW4jSXrEkyPuBsA
znWRfmqzmbmPpplY7hsZxJeCWVcW3Th9qWoVSJvuKvPFi95TQgHtZHPwT8h8V6Pg
KJqeBx8jI7ao1o7A38pCLJ8uA/ShtOv7PNI8IM4JK8BOdenxRRs/7acG+Q1kWzgt
5+nS0AyWV3l5X4NXTaDfQ2CVFv0As8m5Ovu4wWEEYF2vhjjdmP7fCYwXmD6CCF54
qo2Y1ZdJ9QLIFsdXYEb3UN3vj6K057o2hlA2VO9kv5burTHudzXm1SWNQ/ES/jOn
7kzveeaxzPI8tpoaVv9bzX/ekr48A+mC/xfBFBq+ny68TuoxJgMzERCyPu1PQCme
OBu/rRjSTcLTV7wMg41kMLmd/oczF2MXQqf0/7Gi9sj2bnAcjHZKu8SmrAOYuDG1
Z4jN+WZVHv11CpYcNyT2/iw8aPcPt0sz01UBxqYSi+4y+7SkTsNHLok39WfnkdAa
KWu32/R8ku+t24gHkixZJTQZx7+OOwr6lBwnKEBjupasKYM/+8fr4cb0zw3yTWoV
lHsCcW5jgFYLF+2jfSHr3qO+O9zfdks+NDIbhmg2RHcUTZ0BJgcCvT8uE69wJayf
mVYxyTq1naYHfIFcr/aod3JunUXy5TmLYzw4qOmxOgjmZV6BDzLWPAkepp5mDJgs
XFtYxRdmhpdZtQ0xZ/S9jJrpOpm6YVuXGkxliFF3JnzDjUegOMd3E6D4W/VlwWsZ
DQfCz0kixYgFxN4uyS+Ur201Xcpn5QKyEYSDUVvDKbfFRt2XW2sfTpTKcHkqllYz
LVw8PZdoF2llTqTk2Ke90ptDwB0lM2dhkAAKe6QzjGByLJioE+Oss7ZQc4mQBfPa
5QDPPIyZHvsLPN8+cpTAI2CpI1FlQKVTTfLqmMHzCd2YYo3vfm/QFBAqssohuKUs
fxh4OSRPEmn13a42HJg1PZeS1BaR6UShlCPRaG/QWjjaQrXoV1DqHChp9u+kmsj4
zyMpOYjo2tGFSMbXYQJUSka/4VA8dCQklHOvg00FfIAMLrUpk5Znb2bfluvzHdua
29Vb8/FndW3p37Mkh2iswzHensK+GJbT1akcs6hhrlk2B8vcJb7NPdYw8Bk1tEgb
GodUHeZM+PTK+w3xQMDvAkc/PvJpqh1ZAHCg1L4BqDkgcYcgN34nfk6JtzOWqdZy
bjXwq/xEzkY0MZKeiDFX8tjppYKxx/DJBupq8XDA9PuhfUCun9WlfRNdd1mUoSYD
c6tZQENIeEf9a5scWDuyXQIJ4fFwY7DTRO5oCNSTr27kM/4jvEFn1IbIkEEmdFtW
+QXVO0P5IulpBZn8BWISqvtj4SIdEc9BoAqw7b8o1hsPrB23U+3sFDpUx04Nibp0
B5D0Q/IIjzY9YB09E2cvLSm+wrwc0XzYJzgebAbE15OLL+EXeFZleJzeG0FYJbrG
yzLLVLnIos/iWhWQhd2CWaOMuUUQhz1OW/dXiJHPXBz6MaFlkgVrNkS8v9f19UQt
oPxOO99ab4aZgyRvmi0+a7f0P9x9OJOPpiqCcyfJUtUvAkGI4/OlyShYzek8z5to
fsswt5UhnXur8tU2PN1mAoYWkNi2z3z/JY2hZcYpqY2jX6LuZ4ak70CAo1BFa/PC
D+KZfuElfih6ema8gpFtIOefcDIX6ffOznG5iTB1CkMwJr9DRy5EVXSAZ7PdXCen
GQxEg3Dg30DYTV2E5jjQqUkE/0hzEQCx+eHXEG8DDIBBqKrR+Az0c0cKhKKuwchl
7f03y5RAJtada2kto2Zk0nIugHTE35bsAskImsVX6hisjRA/oR7QoTS0GOq1/eDb
rz4pDJINsbITRjoAcwp6I7G2UkBCLsE2eNqIBZ1bSUjA7nUaf11sLHn+IPJhrke8
2qqex8hJ3Sk0zC46RfrjG/EMiHCbAQyWqX3A77SX5lmTXvArMSWtjFc2x8CyHgVt
/ewQDuNqEsGMntuXTV0gf29a6oMeZjAJlxBBvB+H71IC0kfKZ3EDjZDp/ZAQHnEW
eKOSwXN+Zrgg08DhyVb6YJq1l/cvGol0mrrFPDxmMU7nEeV/IXPXhtTqGYjytaH6
x47vQ8nBafVuEyas6oIl6pNib7zG8rlhgYPgzGkYxJchEG1LuMdhRwrqFq21qwRI
O0xS7CKLb2mtAUpNkgQu8v58D1cR0Nrasr7OB8ADJ17NQ18tgVnVYZtbSiKpTYZ/
w8H5W5c51TJ2AeRkrBFzqBYzLIP/8SJ8UHemEL9HICmOdnFseiJgCb/11XEggyjR
jUYUEH1WZRZXyXazpGir5K1jlSHyce3XcvTdMDahhrs01jMTUWxmQfXvtMQ6ncIn
qGJrtBQou2vDihJbfdB+EDISz9ysdyd27A36/FU+C+kPenJBK33qsDKK8U1LpBX5
INWv5/ytpTAvrbWlg7TMQMDzrF1RxlokHEbDMnAmEqNWpf3hMEaiDBflpFdhxKlP
UxRauO70jR+bpM5BSK2bX7CiifooQvmY8QGN7wk37AFjlCr5yJkqTke6QwiFkCUt
0Hi855vX+ZHQ0yzoS3DrAlzndT+eCm/RQQZrppRn7MFkI5B9+/pymjZRnAQPEaoS
REBQcU0ejXznWyk60Bn/WjhJbCMWNxgaySA+cRBS6pTtmfmDI+s4c8ImgvQuUMPS
Ci+Sa+lD+rnBkAFvoCNEa6QH0UpZ3milkHDv6YCEA68FGfmSdBqdVbraqvTWRZuj
Qu8LbwVHGJ+F0pxAcyWTnhd4LXwIgJJ/a1E+aUo6Uw7h/aICMLhMGF59FmRlKRqY
nv4yxkzV16liL7wPb66Pp2/Lps/SiDVumkcZ/Z37hG/VAxAUfQqVcRc1LGI3rVs7
gYYcDeWGLnkjPo5VfeZUleCAPctcUZbkKqwNxgux0H3RjVr12gs7Mefc02GBGjm8
yAqJVAvLPbkm9R7ljYzes+EspUYyhDwT3dSkCFDcLc89D2i7/vMecN9C2hoSAY2Z
4h6ifVK2T1Oo/d9iegMx+7juYauydxMMQnj5HxpguVwBN0ComfBjMQU4q98AI+CL
MmztUUxr6PBtZ5aAYyiF8G/bxobaLcP2MF0wrf00pBRQs1FwrHCr0i6/ImV5kNtJ
VePdBDEdjClyD/45R7Rq2hYWHaqPnZ4GGWViDpI7+4Z/L/s8Oqm4Egj3O+LfKTU3
JquNroX82q6BZr0hpGQXjp8e95RABSJewcm+GiPBjYtq4BNpsir0d6VfdXHsiFGL
31SuSA8auY+8RNc1eCKxpak5e0xtLhnBcGzswnVYPXmcwtzdhLvc/D/HTTKFLQGF
tqSqFOptXY9LMXhrcMoBitY+OIw3fydBl5uc3xqvL/bqwNVrHEb8R9K0W8stAa9b
T5eMfwX0pEJP0/G/MCBBJU5/WxcAkW2C58CPssi+pb83y0+X35V0XvMluruJbCw0
Fk6Ma7nJD17Gk/WjHg4l1nW5Z+4BGiYa1CyQ48h76M+etlEXY9FSkQhmTu/knbwg
U+wHuDri/uPEo8EAmRYDuD5u2SjqfzC0bxYR+hSEPSW71z+SQXXZ0Afnu5cuagu+
eDUyw2npZ09TWZCGWjJyfYGwjtE8jRhBri3T00zSP8IsFkxXHbSjGZwkPlN2yXFa
mO9fl0w52Lj1zofZxY+4yNlYHP1Io7w6swNxVNqJQqHgg3WyXiO26Lf2csP+BUOU
mlrziW5uWdzB5VvA6J/TEein1MkrC8fTijNwn51dRnMOs8azO6tkBiVjE+bPi5zu
rRxSDBvRpFamTBFXLOxpa9S54OtnbCDZMQxG26CYqkT7dwBMtOk4coRgC7mfcGkA
G8jqq4GF5teCuDvwHeT8YAVua7HSEtr/meYXWoJqkZf6fSYI7NWQ4nrtxIJcj9fI
XepyPUCb9NoK334DG4t3VakVlsHvA0xiPoepIGaxqo3rCvfnRbUYKRPor3/WTuai
clEL9Yybv27iTzC332sAj8QioLWm8v/NkqjltIm3u4VcrO0KaFh1/zHLqvlneFvm
l9sDlLnYo3Oslf6IeCppWggDMs/eTor5uRsBYubPC/RvEiFneGyYOXXtdD/HCH+b
1v28hbajMKejzjGVX6HMEJmL6IWdqASlm1mFg8ndxXm9Ygu+Lqk74Tkl7s/nERhn
K3u3AQ+7b0gh+HasYHwqqkQy3d2WLbIuyA4meaTivO4a4p62pDcRPM7is5L77rj9
4cb3pE9mGXtFQIfBwMepgY1Avvyh++lHntmMNZBVtlZszbtWytIkxAsNOky5LJDM
OKzS5ZHVALGMn984igL3jxB0fV/G0BQYgA4QFU0kwMWVL9EDKIxAK6Ur/MdV+jOd
rIFbzFGjveHDy0tRUdTLKSn9MxYdzxlPDoFx/GyVsyZ5BuQoTsndOePu+gvrAyfE
yRrC4gquIJtNSUpmyM09GDpj7dSF9dR7SBJfg/+q5D5p6QaaCUrMT1lR87jhGgkO
sAeSvsyUxta284cpF7t7/aHhZy8jkEWIsfOtSaUtCmpudIWJi5Ma+hCs79MzZOdv
SuoEYEpySuyAFeJpl4OKlBCqmiJb56rmBG8TpR3WmE0LYV9vK1HpN+S3WH+l/G9e
HGw2jJtvUsz71LH019k4h+oWoYv0TGXxSRBpMEHe0c2sxiW09bY2KjEWAi4aSf6m
hpqEwgwXhKO+1VK40KPwbEFYvt6ENHZm+HWb66BxzSi6Q10Sx1b4N7o7DUh3vmHu
WIjUfxHION1Pk8vSrbCeu7lDyLdbg3/kgkCljqmj0uDnMbuAv/716mekX+Aa2Q7V
SZFPxg29PvLfyuqODwXGDoI2iY/7CtBhZJJgmqq0SSH7NBISVdz90r8DGsLFa4yE
BIyJ3D5sSeMmwRVc1h30lQA+2xzyyf9Ski938G4y49V/wmN2wn2RoW2sj4rEmCqb
OsWPKAIcarg/mgvvAAQUK6p7U15CxHIjifz1JcJyKc6X5+FM+nT0XO0kfNClX4Eu
bfIxF7pm4wrPSbzjdF3T26HrNMetxfQ4AYqoq0LlcrD/PqTh0L3LEKruMczj34GB
DpNCEXu8aC8BA7UYZavsKxaVnRM+S/xLT3taRE5l0UpjxDIgaiWPDYINOLDgd3BR
6PCisvcZvEws8Eco4cDMA3B8f1BAQSc49oXlq+cSxu4/gnT2iAdNcsSQ8Vhw0vJE
JKHdIv1lFwvjCsBw7wN9xnuB4cX0nUyDafvtZtB2LHWVqCRSDwLbgzOvy9I0Lm2w
U3DSTuLWw5ww8aa3XY0bx17ILxu9blcrtyaCl0tJAGvXrqsGeW6YLi+tm3WYkb5F
mo1Gb/jDOoz590Rsl5CcdGdwD4WqMgxsFPEuf0LkBY5A/k94F/ODUkuP/CsytT7B
EWuyD4U3PW//XuDptPoshLkhn2esc8vEplQpCgJ5fxA/hCbJywQbhveNW7LSi99D
wJbaJqNA7+ZhUqKeKT+Ghyo2A4ysCgvsUTEx147LnlSbmLkqYNJoHpSs5gxFsJfW
FRV0/MxUsGuD00WZF05jjQhJO2k6Fs/8zmpv0lMTogfj2Ydjlgqw4sxssMmIsnfd
FFSMlxbbpJjIyjV7zUYHF2RH8/ywO0VcQcKLxkAxhIA2sOp+2k6WzwgS1znODOtM
5ZFb9pn5prbigWGukBGtj1pmK6tIdZi3tUQ1AcekFO6CVXVA++LQKwGQ0oQwCeEc
MuJYrEySoUGmnAhPXi9AW9hIzbR+oB6UWPwQ4l/hnfpgKS7I18wTyq7oTEnmseqx
Pusij5UxnVyXtWrWTg/DPh7zsZkoOFAzVoytNmn4bYAk3KTh7AWWq6ZKi4tZFJG3
gko/8AhE569QEG4EAsZ0UzFr7InDfF8FTKlKZ1Ak4EdCFnKKAra/F7QAR3mDEYj+
dJjoI6WqsKr11iUCSRA3ovE9MlSzQytc+DEm2kEiFy8SThtor1xGlRn3MzUztD48
jSgs9zjlZ/OG8U0mr+iAU8VltGmzYqoTF95F5rcBGTkIOvGduAc/yl1mAsEDdUQC
tRZr4Zt8bXxdk2zRVbwvdqLW77gM1UX1M4EXmVbyQ8vftUUyEt/rruz40LxAC7GE
gnzlDcxCOwIYz4Zf4yN0rpPg9n2MbuRp0+GTiY3glrZiXTyK8pyVMCezHGz2LtEA
HJnIK4pjVtC/P+XkX1YQOr8rCxSannx+ZZD3ohuau3Oj6wO87Cgb2Cl9TFw88/0G
/eiLCUGC+NcTcJxRh/dphuwhMBhSR5rVnZqQYcYnxoFLjsITKwGM1orzCjYbETZR
68QkAuhDl1EcfMQWRzhmaaEDkPWYatgQRdDhwPYfeJoM4z8Lzy66v/KqarftI6KU
GyuKUTUJxkyjbNw6bCbFlWwDoK9bwXELaAfTHuA0BiOjITqyyn6HVOyQ/i7Lb7cw
ajfQ8phkGu0WRnGhSfKaH5VDfRX7uxsgptiiUmFmo2+d6BmYJGDaWk7mefr463a6
/otzoe1mttcRvRwYUj9tXK+NXpLpXtn6qiMnAG4eTqxqKhXQmqs6zRGUrP15CGb2
VsppbRtSAJ0nokZ6FQdD0IQpueOcpTBrgLEjpXUe87fJqUMB25otMbyAUSp+mSqw
Gaa+b/jtr9UBGBpV9bi6aIcNnUi56t8aJlYRrPkZg0zQz4wIIBKj2FNdDMWIuE2E
Wk4zFlZdHU+z0wPdZO3Jol2R2uqQN1dLFO+cETlyVbCn5nwqFviyP+V5VszULdYB
VPyhxALKamrjpK4tU0V6bIgHYBYSy/eQZnzROMse1IN+sVNFr8IiCqaDZl9ugjiu
/jtrg9BCpl+dLkc2SuL6ZLEJo/vk42ubN2LsyhvG0Zu3Zs48+yJg2oh7I8YTVpxu
5BeJNjydwurOYTCLpOt/AgktAja6Zs7OvI4dUBZFxz/iRDTS0nBMfRHXRC69lLmg
lbsrcQXeKzgZKjGQEY8Qwr35FeK2o0JfN3RfMjB9WHhAQqAd68iKn2M8R+xpzk+g
+M8BYh05cgDCYcc4kYABjwoOXkttZN/jAkuRdFa8OiHohzYOWLjNmyQPlwcnTy8A
jYUjLeVOBF69woFdaDT5BC/n8oSJKdQcjusFnFCOtJ7LMxEvzbOcRTrtqoBuQpLz
5SQSvBvheVfzJiBGTjNCwwU554rMwAvqH6y5NPpQ+JxOTX7QqqbAomwRAEG1+NXy
vqKD4eLtkelUbkg0f+Db+bXqRTtNIm/LCwfpTdyxDpNMgF1NuAOQf9tpDjSIe1E0
z/eVWLaM4UOHplvPUMSmZFlPRm6GGCCqk5tCyEgM9mRB/NbxSrlVdiNYMbLuHtsx
OVqrIjdMe8RwH7gsYW/KiArIFrBeRmH35PpNzFGt9hHX9weU+pfnP+xHvt89iHc3
gh98wdBOlxTUxLwzopXUwv814rbPyYu9NOaCAL1Q4IEOaBtQVTwrtlXY09O40HMG
UmgjqY/Y9jZ+qIhAR85WEsUDQV+dDAPmA3Eqhj6KgvYwrZ1Xjl4VHi6NodmR0bIM
yFCaYLVXZCpeJA0TNt8wUQBcIKAcIsqWecUUMwtE5qUJUzCkjYbAreRpZraI8rss
TNXMhzqxlu+LzbDSRHQurxclogomE56/Cf2QDUO3y75fNVNpthiiJIk5bC62jWNb
zeCQMHWQ0DEuJo0uW5C1jjiyedxjW0r9Qt9bU0DJTOKHDiZqe7LEkO0W+wrsKiGg
6ORlGRqwyE7gmCelEs3tvg1+bbW8Mi7zDvngp3Gue5+VkrLPPGkcLR/pGWFb+PM0
PEaClnwAXC8btkKKYDFhv9O8AvR5RWcXFgdplf8ipBd2gKtY+nl9K0lYZl7sDo+6
+Yau5f9qmhl72SkMqpwb5KN4kXMnS181Ic9EzEdLMFKxHI5lT1K9PBG/YPzXOGhY
tRpA1QMBjF5R2BdjuInzqABYCR+c3kzdWClKHI5EeWb/X0YL1lqfKhQgHEoxjdmW
MCFpmy/LcIFfGRnPzTkY6nSu/2oeu20K4tAdd7O2hUeSkoPQ/+OYcDsfSaRWgdfr
dVc7U1CjfLUV3asxoLuDjGoHgOtvrHI1chu9sqGt3q/u5xFb4+lGLqH+EMHHdCak
xZRm/FlDYx0wRPuyqUYaFten0vzXliAnEdmdat9pG/XZHtusqzEzrXRV1qMshyBC
y+v92Fg3S1SatvJ3lMGCHi0OmnCO3UbIPpsDkJxca0G41v19KpgfYh5nwiRZKszQ
gVXxg+JfgckcX7rvEY34N9FsaCCDv/anmuBPlo3QhEimWswgAviKUwFq13jb90Gv
5x34OIDi2Bj78Df4I4TQOWKBaBd1eohxJk7bBN29O9ID9TbeqfkXWqg5dMQgFGke
t3T2yvO8sJIU7SyF4ysMguqInbwVxomYV60ZrFcMeVQG0sZCnde7cE1B5ZKPEN8/
0zjQHDs6XLLPDDSwv2uVI2zK8uIJwGfyKSLOYdru+Aw8ZoH3UIU7FdSQjrFpSFVJ
11Iezi2gcQirrZSVO2e6AV6eoi9w8PLpjI7IqHc9hFCc+Kq8CD/gohJsoOT+uKNL
En3vSpMv4knVQyDUdzON4NdyBFUTUCNCCRH4Tzt3sqFggcs8b1P8yco8wcCrpDNT
oy/002zPyNgiYngaCQqb4NCSAuW36QROJD1OlI2g/KMUdJkh1ACAksJzGpEUVEbs
FpIAAOxjetFkAKGLuCC86WIPmJiTuz6TJ6VNTeSAFgFKblHwOVlh9v02TeKOSn1f
qeFHA/XJCBov4ZunGiquV61TG3KG9SHkY0UGwUoznT3VagdNH6Xex/Zow/GMB2v2
uFMHEOvqWD9YOxPBSUylkAONHo/UxIEXzAHNDplAIJEyIFzwmQ+gDaiSLcdZ22S/
LWinByZmTQxrT+gPT9TMTlOu1tudrKpK4R9d3XbCNb2qTinbVO9mGsGJViE9V29Z
52cCXx4fsnRg+b1Z0r0a86HTM35C2/BdlajJZfP3VlBLLjdrb3eDHBL10+dX+CPj
ZNF5PlcZgeNzc/jhAxACjZSUFUvfREbWczNGDmcFIm+pu/j2RqQcOJmSb3Cak8JE
KMxzjyosWd2Z/gGR9iPOj0KjHdZdCkka3Pi4zHvXgERT2nkOwg5m4WgE7/lyZCFI
pQKKsXCN++J1n/RtFM41D2tV+A38+ItrXbWAFlbsAwH8aDfZNVhDW8rSKSP7n509
K/0xUqe9sNPLefbcRJYRvZNzAHL+t6YjOnJjh4PZ2vcrFnHcbuhydVpz1Qtqa5fi
cqWpOmqTAC1ga6WlkpQoWbLuLSgUdBETLBt5L8m3q5T/mH00C2oMrhGmg5RZ8Vvz
pk6ijay4UV2+H/JTMjdaIczYLQm2UeLxCASlYH4htOi9sTr8fSw9/kkorv0dlhRG
VkDmMuNF1rfPZ3r4VeUoobb3jvNdjzYsYqoi2LSubDQGgtRmD2ek1fmeubp1aQsq
tZ6KskkgWJhXntgafpsa9EeytGUCSVkhcz9+v30L8shj+KXsPjE6vHmMunho9B6d
YnKcYaEHJYMxCGfT8zGNGKj+V/0BM8n4PbeMDm5+zJlYPzaz1lldc492woFazbSK
wreFyHIiUEidPjeHFNCOPwqUsdmYQ4xoZBvDMN/Y3tJ3SZY/uJFGSyfWQv1RMCK6
sJ5JcsYhPP1cZD2t13NaMccWoUayaNiTRK3UbaiJWzwKS3EUoPKRkD2tvvsVW099
6CoDUQ88Wwn1BGMCqitsC/eOySNOLjKsrgATUxMj0W0yJ89MbEYnJEG+a9uF7sF6
RcIE+z8QYOzJt5IYK3jbLaOwwK69kniSBR7RfuDIuVt3jJbtjZVKduFTqtMdhiII
oDRreeC8xsINqdTgT2kLOe2VdvVRvMTf2b2NuGPoPMUMzos4EHdGRCjicCOLfvK0
5M+DEgSZLt6tRkZXmHswHOcILV2aK3Q+HyskNIKyvlClDzXZh0eyA3PDvXAOxyqa
G/GxFDwGGR8KghaHAXXtw1n7dv8XWDjJt73oQfrEwg0TymrH3p/lrIUqrntBhk7o
9vGmFNwliIgmi3GvOoyUXazIy/xNttlpp/PLQTCpY7TO+XKBTIcY9sT3k6NG2596
abjhyUfOniOuZE7Z1DvmKKh6warwBQB8SJP5REhuORov/1OBmufqYxRE2kbvFtVG
vLqyzhmt5Yt363F239Qol82FFfhhCY2YkzninkGvHqNRxZp7QgM3SR3saqOBxL7d
oxpDx2qj0GSqWDJin6sulZBqGziS5RZi0gSzoEhzuGxX+Lfms5+C3PW0md6LZeZg
2uvNM1uZInpEdsH++fPZz981pNPKAKTaaQfIReHIj9ok3XLj2hk5pJmXpczymlmU
RWyg1BgYyrqEKp2Ds5rXETngrOk2cR8e1pxhL+8BJpOEUdzUhzzFl1ug2nGCIbuf
tEoppGzuWs9VqwmblcBUeIKjL2mVnX7Y3NBbHJlWFCMkK6FaR+N9iyJV/iVcwu3h
2SP6OH7FADnht2D8IEfmsbnoar+30oQcI2UQGcscHEXbnlOvjlyGY+xwgKAEyD4Y
yx9T9ngbloLpyPKnIbv8OTAk/fYc3/u2kcxtbrkABLdBtynmvmzKreFiW7IzxLNW
QQtQ/y21IKtG6m4sBPyuN2/i8vLgtltxATxzBvqwzwDqskovJLA5dCwTkSMgY2Rq
2CfGtC8pH5HVd6nP7S12p7Am9erXYGr965ngJE9/6F1vs6oSLslI6E1uXWNSPJ/O
qMcZDuxFSBRWXCmdkyko3ijbud7HvLE7+aaAitBma/2jy4kIR3Vs/cAun/3Oeeip
RguXZqIn8u60E0G1AbZM5AAJhY+8Y86o/sghUJnoDAjIgxpI6s+A3uShSqdkkdR2
yg1vcprwb+30vl8tZpLnXMrsdJgFkLrRCLgKkVoAaeBUwUU6C4Qz5+J6eeG0GINS
Z873qXRp6jSVZySbaaiD6kOSa9Qs5ixE1YT+YBvb7EtPj7dP8O6FAWhzTkMHhy4r
kmE60qt0XSm+FtQ+G/ki1u0QsfE9mPhCNaFfMhM1ysObAuz8Ginn2XPI8e6RrKOw
Ecx2E+PeH26E7tcNgPiJm3utEhtEBzigaSAadubWckfPX+ZxUwUPNG4l1FiJgtlL
QXOO8xW0CcntDmQ+A2tekCUOmS1mDWV8B/lj9om30BlNdU+vkOi53mKhpsEt4XY2
S0MBLWwqTcuUn1oO3rkCD8poq7aPrdfUQLWSDY17eDJUXxWdp9fLtL48zs/7lKS7
hAkuMdvNFU8etzW/Z3KdeoytXrW/Amt42HIcnG7QOtzFBdMnNfAumvkOECkdnz3E
z7Gf90yEOjW2Syo7WLUtJ2/8z5UHPDaReX2JbX2e8p84JV1u3K+r/eWdDURhQ0ED
ly9Aoyx2c2MDhKpAU0exFE7On6zelbZbmHvMlTHQWCA6uCHvm5peXkgLeRXSua2D
zaUwD50YwMyKUqF84+gxCzOClN7h4f/R1uWKmW3cj0IbSursFmwPCK/8U60wUkei
1tsH/gv6mchMC2fyzwU9qQ4+lXvx4QUkgQyChf84knjTAEO++aVbx55V122Ql1cC
FJTRjPjQlg+JML/NqnZ892vr3HT5Kwgy3ahMvcfazjKnuhmPyoraQygRW6wUbV9g
PycZUuq62XzQXoqKDzNatZcCfKL3qIdGCFKjC60B0V0GJoh1HAepepuf9dE0kLpH
Xua2z3VHKGEqVITK0Pv+GpeZ2Gsnx3dKSoNKXBz5f8whhPiMT9ytb9OB2C1svIUf
tsC2Nq+hR0Eb/hED7dVbDbkiZqwerjZkgQUcpr1sRHoVafepj5H2fHO+H/ZYro1i
XgAjApSG8ycT8xaegoyA5Kx8dm1jL0H1cuxiP63CrtmyAPesTXcNui4O12KUNPl2
R9em8/pkDSHt7CfAMtS168Ji8aNygPczEC94R/mvFHmX5YG8c6u7cUirRtF69Set
bNYO1XjQdsmn5PErnagBL7h020h4Xl7ap03pY7ZKMKpSV/JTCBWpsSpl7IDLIjSD
IFrWSPD+yGljD7OBjchnBbS803cT+v7HOwGcJmTqiJ/hCq/9ttKBL5xXJzMIisrV
zJdeud+ozv7qbVrHE2Pm7PRioOlHxsQwDP1KIsqDa+txbFU/kLOx3pXtVBz7CO6e
h815ZfOkHZBlTswdKK25ARRzYNTypKthJ9/xuik2YXZnq+zepMu3aAlArmyRKN/J
iJZjapcYJj0NcZ4sStx/XLLUVo8IVXDTfXYWdzsstF97SOC/4t+vLpsqF80cR8Ft
wYWxFFHdqdjJRq3LH2UjfHgK7gBaSsSeirin8Hya9HZPtJGenqFqM1sChxxw9twG
lksJpg62dZB42B+JGBU+YyVlyIqXbmTM29wbu3/OfX1tk8s0wzWA5Gq+bEOvu1RC
/EfmREbdLBR5e5BtEd1un+a28DdJO5DX4mHrXF5aIg8pHL7vDmnkojTpwLvxWBXS
SkMghjXuHPwqhRQNKzkli56fw6qHIgIzT5ef+IltQ/xcqJSo/yv4xJmAWajEPhhO
rErzF/hgLNut35+SJstkLRnlOEqUivcWyeQiuqFQ5O42jnaVnsMrBFq5RSx3FagH
fj3JwRgYYck71GLhF+B53BBsJqYhDDFJMuq0qGfFzQINdrZn7LzRK9boxhtOTnYe
SPiALjkyidrnOKicFrraNSTZ9BMw735A+bMSYS/XY2S+a8k4C1wqhXPFu7OCFcZW
6Z32ahO/laXsSL6JszLSt3Sgnf4DXMBru8zgdj4zYXIuDMrcdmxtTqNCmsCunUoF
0qdwDGhaNzsA6o0gk6KlCcwcepZcgE1bFG+IIWbOeGsuuhgTFVlPPqe7CK2bAi7K
sqz+/0vLLIVbwCzsmHFc68NwaNGDU1YcbyozWgvPsgylVneO36rQUTVaLmSXqGTy
vsmAINHf2Pjj6lonv2qsYZXgyV7LO9wdh67tIRUHAgwRjpeTLabMcj3ALpA7apBi
j03Vbl4FTtde3MzX0JA+59kkKzZ7RjHaiDgB05dcaC8HkngwHLv8I70xHkkXsLN3
nXKhZ/mnkAVMTcDGXnYhvnWc5Ehf7YWsdomIiuioPP6nC2EydD7P38fKV/aHou6n
RVq3/5FbHIQTKsU0kXo7dMfInmXf/fEBEs9E7ZWov0LcjwaJSVwXlumX+7ERYtyz
mANrcHtXeyr/Lmh9m1LZ84VFvcTzQhHb3DA4/qn7smxZ8MlH0J3P4pusS1PvGlMn
lkvVxpytkgirVgPc2W7PwFq7y0ISnW5F4xpFx/sjn3WkABVOvHKZVjlhkY0Doi7T
lr7nzLR76BxPbW4G/U7mSTFeFXFR3QjapZUjRHlqDIrdxx7i29KIOpoaLyyAqV1F
pt7BWJALDcdWF/aPK0kVSaCkX4U9KMeQOsXjOaiLPKlXL3ddUfpyvxI6Qp6G6V8+
DHGA/WNxQWzeaS1ULEOpchH+K+9tR2HOi1tbj6sSlyyLtWnmfDSPtY7hPG6G9w7D
/tbRZUS+j5Fmf3AVNj1TyQH6o6RU2Qce/5iYFniCLGYBl1jl8FFgW9sY42WfEfSD
buRBu6oxz9RukbW/ptMDno8uUxYGFanmuxEScsjQaCMmsaK6ZQDsMaKfxvpXdGgx
ntOgwY/q7Wl8aAgGDnpXmtO6LXfqH7+l/djm/apgPs8Izx97KdIsA4FeHMTZg93b
FK/zKwv6+SNDnpHErHo4HSVVmC94tQCnQFhaBYgp26riH3x3ViLgBBR+sEfIntmu
/MCQMXrt7eXObv1FXbFbm0BfielrGbam+kpaVKrp0VDjHDs8Zrxv3K2qUlk5vy+Y
G1ZPmT6dtHDP52tALWPwbC/EtY5N+vfppJqMq0zSovSlzR42MQgnER62oLUSDWts
0VNBooGV7G48jWPmOD2ffw6/W3DVAbBrShtPFg5q8sEmdRlU51MemGaTIGP8ab36
rsO79pQ3949d0IZjccDJgzFJuhXOrpsLHqtvkbufrTD/IFGXYnDSGbd4wBXjpRld
OwXKyMxWDSjMR+UpbuTn1i4re7IlPBW3aKuekxLWuBFO/5/lXtQIuC1jK/EVo02U
vrRHCGIO77hKeW2z0pkKpoPgPDrifnlO7ZUQDDXVVrWmSXSvPflwO3BAVS8/Nx5o
qhOE6rQHADT1x2DBiLKjkRl+X0iFKjUwXQ3aH4uEkqdh5WzP/Cx5pmZuBdU9W2TM
rYwqRj2eihJ78YcepUqLjbpNP7PK3mj7cfGY6LY+bb2U9Md3jo8Bgg9iVQV2GuVg
WW9g9dt/h4bmlmfTCi2pMmsricdrk38O8GB0nDjcKfO8v/o7kQVtBHfrT5ViJJBF
1qQpWR6syGsVe0Q16DHQqD/7t+Kts7eHvvUhdxUOzxMXtBMKSXGyxb423DnKTXjJ
XIKblHeJLnsHhgrDR5f4VJ+1pv2JWmvt5MgoqBrnv7RnDZV1FYh3UeWz1AMv+62+
GkKxu7tJo/hETQHjEwdLN86hgQyuKIUpPkw6jm8OG6Hut39Hq5QkhQgwg7dqjo8V
YPL+iGpGWaJXXhw9Ry4lckts4dw9teJjF72n2lLleEqLVpeWpIgKnyeh+towqCXm
Z3hnZtloEcbSpQ26jhyohUyAEzPTm3rtPXrD31f8YIV1LWJJwrmRKQmPsnKlSaLW
/W2SLASkPOoBPOP2K3uUz7ilks43u0u+0ENRwMbEjbwyldkznlbrVmM1l96VvAA6
+Kdnl03g/fHZORh07nvQ5XvyMkcCQq/tGp/qtKvPdi8K4U5De8JJ+BK+MKZ3zt5a
FfIYO8QlbXWTHXlEZuFgrtX/wQC0DpIkhSDRMpdibzuDivsXEtCCF90jHriT0S5k
mQMrFpkD7zwLgeGwEt0iZ6Qb7ZVch6z9By6TA0GY9c4fzF6ulCzBR1lNs93MAhHa
U1d4DD/zec+mJByBi/XRhZ/UvUKBbvW9xp6VIJOfQJQbMPT2rK1edSSYlS0X5o5l
b5mX3or01sanfpugQehzl2zYObC9+sovGYm/VvFtPiDLkAVrSpHU3YXgn2rZ2hDd
t2Sa4SXEJOI63lt4P+bsyrY2PuYXFMso7Kz6BxSVCwRG6EG21bsMPHbsvnSoRvtj
l5JlZsxVMJ6rpkubK2EARe7asvAFqTPRe9TlLBLLkUKFZETb2v7fTAlTdgMR3M1B
zpPt3D3sN+HBJFhYfW5rn0Rpfgp5BLyCqCihrmNCkUlLBxhOKnQodeDC/Prm5N9/
tXBymdNUCozB/7dKJmF49qjLWxRVhjIAwJSNOKj0KSUrA0RfkZ+1KejPZHzgKTte
B5yCXZWNGnKC0OxUhvawShLkez824+NGQK6CDdrSZNQ6eEOuulNjw6k8qZ329XdT
GwCvoGILP1VFKeCJgv2o/qZVS7tl+HPa/VMriNz6YWVYxi7vGPmAaTBo9niYFXmH
pO6+4oCL8MLCgCjNdrk4CIYGeI2Ht0Iy/S6048gvrbkpOvbmUimPoqCML+Sx94by
tONxYDR+PzU01sReEn78kx3ptHn2Uncykt7645ff7u5uJ6C+ihG1vD3CRDWz2BsK
8LrvjCKLhc1tSymsjSsssp5j2OEBou4oLMNeG8LQcfEU/9WSBf0XiJBZgXgPMn3i
7v7yglv0oNLuMtMsiIZlEGvncQFaDzVIKnMPxEJztTT7Z/4WdZ+4v+C1VPujj7OC
HIuxuhv7UGdnJYDHl66TBqBR1lOBMMVtoKZZ1hptNhWDr+CPns8PiUh0/Y4Bee/M
wgmtcTgz7B+BPrFcn9FWSA0dYHxKk1rQ2g8RD3yiKenBs22JTDsdnl1pzR7s3SjQ
5X+Qwa+yZBD5e8XMVmqmtBup5ONjf82LPgP/OHVO8tEK0xySA5KUYTWdCx86Ru9+
BI/CkLKfDbnXkpjksyOnrGy78Tjsg1A0VxKvogFvEhpRkcIf33tafE885z+4+Nu8
M2eGcPDQ9GWcNArtZHRoZZhQFicA/pM71uUkos+MByeY3R7WxwZMtRMhU+LC8D97
temHqi3VvxN+UuMoCS4TQBtiYSmrFnnDJH7EvVP132SprjtZrUl3Da139atxm9vj
BfKnO21UeALzEYatJXVQfxFsdFBrttB8GxR6iqV0qWTTLWBCUR5KPpGtkz8Sa9kb
k0ELTvsz7lUFh/aNOKWvmr1ECHaq5et0G90IiClq59e3Zd+UH91vakEQbS9YhZd1
7saWv/TDstaITT4mHrpTa9uvAwa6Uze70lHreEh/7a6YzgryYiCt1HWaOWZkR8xL
q8YUgjahiKu6/GR0nnpiejqW+onlkEJc/pZ04WJPp2fMN/w6TJHCzcuKzFPsyDmS
G5isLe2iuom4XGImTQy23NbNMjMaDF1gbcLt5cS6KLFEhZzDJYzvBrFSzZFfu9Yx
U49SxUDV13FiDx8oHI3v8H9tUHWmTafSO+QVKe8oRf0UgORRrV1u1vEN384J9KmG
p3iXN3FZ9B1yXhTRCzrCE1YU77WJWP/9i1/qqf4DAY/OD8wcoofCvLLcaWQqVazv
3ikF5th3wIsEc680+7OuLM7xNVfI7jgFn+glRwlt3aznqUmoav/gdOqQ/xrY3L0g
BghD8N+EWXm9W6yhbzizf0WBD8hs4ZtzrmTSGaFLoUKNmeAdMLwZRlpTk4DPbo1a
rV3br/ina3II35p0ch6OD6NBHA2hRrQ5n7bpg86uPVEfnX48bviKn1dB/Ehr99sD
hX7fRrvgyP5STB4dm9z3I0xoKO8TqCbJn27s/V8aHuzPOVNxh8m4AaXAGdCpKEGd
DOw7GqRsD7SD4BzmaNNyC8cPtFfcooJc06Yh9qixAXvMNPc/jIgxVTHqcbD+araU
2hCiSAjpqdxKa5gmBQLvjpH3LTO64cMfoVPYx5Hi0HnXTq6OWFO+6QNc8nE0JCOY
k8/mk9zcakgN9/0B/0mdb5r99QqQanWvOVVug1peV+sQTGWahuH+u+TsEa9Wk4n+
p6DqN/vic0xubk7QvrAwI02E5eysvo1lhhtBHStvPoo=
`protect END_PROTECTED
