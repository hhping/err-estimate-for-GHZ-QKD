`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vQ9t4TiSZs93rDnLzdSpEBX+ysLIm0iLbtNHM3KX48yUz4/V54b9GrQwa8dcyeIf
fYwyte4WMyPdIC04XxNznk/8n/0Q5LVbFnIa9IaMgrR57WvC3Q7eI9bM2ZDmApyV
AweETxfGFtUpzbO0Rt/X5OmqTn3ZGm+aKnnM6fxwyXZHwQiX92t/M7zI2pKYBaJ4
a9bWtpETdQCvpHtaMwmjDlP2kGJ7QWNc2Q7Z8xQsJ8v8WEu6Wh8dLoqyfD247Nd8
RvZr/MVWl8XjV0CHPciBir12pou4SekO/xp7e671sTQwxuDXbse1x4iVH75mmFBC
6LuRCE3RYfKNXF3NH6lcNpX18qaDc69ecMQ3Q9Lv+W2ooycjAN2W2dvBJgN2YinD
5k0mOh1yBWVPx9sHxmrEOfJxIzDrGjgRr0YgglqXhp44TegN3o9VAwPR7Nh9JjWp
jZuOIv0F6+EKNeVDR/s9aXvT45KPIZxobTn9QkXX9onu2GkFVRdW+PccfPq0wlIX
w2P8qLZEMXr1K9cEQn+yo9QNmzWB6+J5jzAOzfl1EVlR31e/3oPdxzHhXsc0/ccR
z2ru+y4z4j4hrkgOoCSHWUB9RQ/PLkin0U9/b8Uvx8h4rQod5GURHl6hIEX8NPcS
5YOGhE8cNBBaFmCmtz4UlX2aK89eLjB8FnP3Ml+kq4wN0AKUZcQG3ebZsxFC5+Yy
A41Xlcoej2slwUtJ7lHOGYD6Jr3VfhMjPlm1zALktOhDxBCRFl0HUVR8HYArRTEg
5ndKID6e1HPk7S/DYYK0+64nM1p+jWjTW+kVQOdGdzbAf1LDLRx2RDelrK+cPbWv
yvWk3lWqlpYHudZzPTi1OLQZes4t4yU2oC5XIGULgowqqGagKT/y3Y8kkEZklONd
i3wX4ket+jOvz5QCXJFvZh6hUlNVKge6CxLLPVQBs7g58lanrptpdCy/43ih2xgC
c+vmyVnd9uRZz33yYCyc5nS4u59GXPWEHR0SS3/o3ymSycZovTEjDm0XdohS2wkz
YLEFcQ1aWFhyDs5ghfdS5M2R0LE7CUrp/duy5qkwN12e9Qw70FFGmCAPBSLahW8H
+xADn+36+cZDAiCyaPHjTLxwUiKnq/tZB1BvoVMsWmnpdPSoKktllt2NIWOwhX4Z
QTFNxDRbhb2i8okLxjGPZ1T5IIB1xPoD7oKG0B1a3hiGgGm9fbDUdGN49jsDS40T
srUcQ/qgcHK9H5D5b/8omeIxsGAy0HHxIbC4Hk8++x0FE/7UzDVTuCN/H6cl2W7/
qJRBOdl9QjG4dcPYanoFcsXXdHvOP2HHf9kMbmZ/HvHRjsL3xtm2EoixQWqRvECO
QecgNmXLOs/6+DMugikr+EbRiUT+ywJIVLUuBZE1QoZnIeiu8VQbl1YzIv2CPHRS
PE/vwWfuPeJsgpfkY9w10B+RpLIJzZFt3MYmiZAreLAS5MQO7z71GBlxkpPpO6FN
1g5M7jhVXgSPybQ2JKCNWPzVUmuDHCY5YirZ+XQnu5SBIsi7wnf5S/zEiw2lIZXB
Lmnxg57QEa1v6m2InEuzIvH4aHarSWOYryjKW/tMAoo=
`protect END_PROTECTED
