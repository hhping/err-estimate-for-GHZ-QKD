`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w84wUTh2Gf7tKPt+prIu4TqaqdacN+GEmPkN7uyH+3LVsKNQGrjcdbz6BVzlJL4z
OQRfoCJHEFYXrT2j7cuVtR8Nw8CNXd+TdBvEBZAWAb00w2h/xHZwHD9978egz5Kn
is9uwwX95BIgyH5Rs5lEYcQeqX7R7fIfNWAu87frbJS2ahKs5jdX4ii3rEkEI8HZ
txX3haD3WJ6HiozxtetOqlw81OHvj/SuUjNkQjxTN7iyfOErbm1EclXAOVicrDoO
BFSGgxDlXtrpXgd8M/ASXLivlD0EVGkJ7vYarKwzh7+f9eAzHYDGbx62j+IQqU3o
dI1EIYXDe6VPCoCdR80x9RuAB6Hz3t3gQ4j24MkLUyTexW/iR40tAiyHqHKQ5XV8
AWU+cMEoGTWM5ymR54fgP1lgCQg9pe0UGQHWYbX92d/E3UyyApwN5DPtUjwuoN2o
5b06ukyM3bgkAIgELb7Sag+iTJsVGj8fmewOkjMdT1Jq96ageg+Chn9UV4TzoHv1
2J1QiT3/Dc125lZlNBSzzN9sTxNf/67TPNy79MUZJO2sKJ+MgWauWvQqj8KT3tGn
U28YnCtEmuP6Me7jKUcuW2uib13bn9D6XsoUdYE9FB+uaz2X6bK/AXAAtRb5+5BP
J1tyPj+ZPxhiMqwqfhelkFiuyOQT/FSEGDTXV3FUTQdqty18MB0fnPkR5qxf+92/
bYKxOxJDmlrEjAv6eO1KP8vWf3JN5zaXmz93DtM43zc=
`protect END_PROTECTED
