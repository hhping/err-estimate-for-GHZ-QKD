`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VqDKpzzrG9R95IZXEtodlacgDna2SQLal74WTWKBpNVjp21fpeCHZBlISribLBkP
FlFweHEla2x0RnsoIAyRkZud1PEtxMuDM9Ozt5JcfFwpZQFXfCym35406JqV0iWs
IvjuX31vAh1UtCF/JYzw5NdTCYh+ndvfkJ2Hg5vr2dRq4/F4/dmci7HvLynQt6i1
zezFyJVA+T4ojD4X6oNlUVfaJMF+ZMX3aE+jhwmowN0fCWi6vZBLsr4L9bA4wJ59
o5MfSpcp1YS3Bf5gCCzMaRyNYqaC93B8ERYzUhNXwSfVaeejS9OnsPwRCEdmudVL
L1FcXUY9QC+q8tzJguX1eYIJ2LhR8d5q7q7tv8BW8TLP8YX1GWvboZi5uyUy1/mW
eyEquSPckQr7nG/v/+gMwqDR9cqyMS5zTZHZaP81ONzCoE0Jj+KDKencGW0HJ6je
Wmf/b8Wwd3aNcp2pgdFydsZKbfWxy7wnndTT1wbfg84W4fXE2t5P3MV+3tFodHc8
XNLCcDXI3MgrXcNPat7q0/5lKHnYma6GOUQdrkaeHnCn80+2LL9yYezNfTW8PVnI
Fwh04PIjhn1RMmfiR0tw0bmrrLFHUmORbbtdBONToGVbB9A7HZDkB6+guRnd1REw
tBJU8H6Ha0UkIhM1b8KWSmjz1/s2gwKL8WKh/p0TS8sQUm9c+jUDOk/8h5hpBsdm
bBm8IiSpdMorTitZYO9d+yexKQwOR92uunF35y9b69saWnUwbYhjlatiQxpg7Fxi
kmI8O3wKdlcjESuSLEoAXIl/Gf4R+Cjr39d8FTaoHkWDVjH+GcR+7A+CVKPhxD0+
c39+cR0RBM0dXwiDv+QTWHVYhJLQYjsMzzrMtGK3CfXcqDSBK4tiRyPvu9TFdrhx
D0uoQwhBTzofjC+pxYIXwOcA45ou7yX0FtX0qSsnikoBRD2iIXN6uiGLp45WWvr5
5yIaL/e+SUyLHS4W3Lp9qdYmE7SzmkaI8VSlx0JTUaipzMtnzfUW8U8p82jD9FJ4
BxPdSyPmCPrdpQ5EahefgN4PTA/xf1WLaRqpMBE2db2F2pE8Q6i1k98qRZtsiu41
cR+1V8xUC08CnLdHSReHHvv4WXOJk3r+VQYVRJHlMjG/EABkONn45xw00LMGcdwB
tlnv7u/u5svY3CobmFrzFXDhKUSTT7MwJiWKaaSYbSPRAzP9lxlorH6aRBwf4cxx
cVqUSxbZ1l5cMWb0knt7g0Hn/2O/e1+roDbrjSepU54LB13MhJV+fmxLIWVPuDHJ
yQea2wGFj5jcHpE4RzgmRkA7Md5oXe8tTN+hLujW/6ZV2sf8hhRAXvAl0y5ihXQz
eLFDj6IbLZsrP9EdoJresUszgaMboX/R4X7z+sjNtDLm1n1fXAtS1DvRGxnC9IMm
qb2Hr9iYRvaB33LvlYP/IzaK7VJAbwAAQeae2FTnIqIdcg8yjrMv1yCw3DduvylG
F3RWFXPg5scSCPqbFU8QW0Vp3c8Nv4mEOvzZhBZFi2xmJLQjLXGBAXzyV/IlTqrV
b/x29Q549E70O9/G9sxzjW2bMAlTsoi0puWYtm+aeVuEEqye/C/9jxOO3QUy+CtE
Mr4BOc6W6rusizcQxuigmd2nEjGrWJZM36+HoiEkK/m87IUaKJUND5EQz5UHUsSm
IRacRNIn+tUjv7YmFHNURKJFiZFoAFdT8dVZDs8UYwbDhu3l96zUXaJBUaXGdE1s
hmxVKnJWKh4xhQVT/WCwHr3gEFD0o6h8S7C/0i9j1QuADWPqTxKdrEIwK8bnDuUn
`protect END_PROTECTED
