`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jBUoYFEglsamsi7FzYxgtSPqMDr/seKAKDihHrbvODTZ+cQkIa7YRdASnhc+SuUO
VrfuojTFakZq03ZL6MP0rFRzvwfJqIuj78YxB2smxWKKUmTjOqPFO+iYasA3o4PQ
BHSWrcEkUYN3fOZ71qH0H3xTDxRlaLh+MzwzkNtAs3P3qH2kPkQUvUNlRqYSfJ58
CzmQzjivPyMRIGy6m5SPQrW5EyU5vo/P3bwZvceJ8F1ZdQpCew8e1PU33YkfkQvk
7BTp83prgmp84azj4S8ueB1HUEnOGEdGG24ELZyjnh4wAm0pTwLqHH6gwUp5jiXc
nD8vc5nIYh2We7weGXxRBem8vr7VzlYeCCX0gZBBwZzFP1Vv2k913QG8oo+liXib
Mp7d0qQB5sxwSwSVzIt/QuaWp6+L7lQ117Fc2lG1SDwKlDQyESe2LPUgrpH0KosF
CSYpdEydVj/txIxUKCLHvYZSHt53y+87b+WxAScDIGT6+fA9aTx6ip9tCe1PfUpw
BNEGrjzBv0ovwsMvPaQMUd2mr6bVon2S1/2pNQYUeCw74kMVM10FoDGIGk57rxFE
42lmurpsrOy6MXHZ2RvtTSA/xUIonQrESXFYiQ66388mtpSm/v/0jmutWoNGfPPV
T7h0frUZqpFqX758Io6f7bVb1fL5LqG7bhdYZoc8d0qU5bbTD7iIKG/OIeSvE/QJ
k1SIUPU309ouWvO4J26IAE4ZV/0Jl5AozOVb4BF6zDeOgE5aU1AzeS9HfPJ4jF5j
RxOihJe2V7Ci9HBL1RjEhN4DRqL0d/KXic0fYkwpm7byN+Ie524vNgL5jxQzF1M2
`protect END_PROTECTED
