`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TK8szzuBQdRAocwH+4VO0CkUNlQIHT3GDeFDLlHfpEXELJDYMpFRs90cWoAJmGCT
o+CnHSmpMb8WMjx1hZPNncYalVvRx1l2/LoIWSR0UyD6tTD/Srs4w/G71/8UX50B
vG6VdYxc0mYZn12mFy+EvmvvONRlGXof4DusTs+f9UFcfjsFBZGLfmMhMdkKOKN/
9zBp03BEK1b74FmIDHJvBbpyHmPe3eVMBmXxDq1m1sLY5UMo8k2583ZOsSlQ9QO9
hdjxduYcTvF4oQhbXDeBPk5Fff3MgpBJF1U9E0l3f7AHcQJq5yFHKRgfxef7wQQE
`protect END_PROTECTED
