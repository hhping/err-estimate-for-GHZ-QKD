`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RCCEfSU4E0e1GMAorMiUSE8X7KaJp5sFFvProVcKLhzHHF3GpEzQxm1rS6DOeaBX
CuxiYphyCkzSJLNMgr03xdRlcKpeGdspaaZ6blu9Wrqh8zelM6jocOX2GSLNIi5X
9l2/lzPA8sNSA0nEkVCQVK/33sM04iTHG18DIo6bf7R95VynRjxfXwWS72n2Q6hX
SxpltSX3MzTDWGPfHqOdAthlbnssjISJCXGacBUdCa0JBPgaIl3X9thcIsFx13rt
H3xBOYcbZV07Xk4mCXFwQz90l3eXNUt2RZMnlef9YjHfyQJmP6BXp/apBFQZDwY8
nuOj/SSJrIedUb8JTiGi6llFiTPLZ2HCXugH1c7QLeKPH73jZ0qVocESR3xanSA2
8fH5K7fXf7ssyzdgjhOtrJmQbzTCAOU84sczR8xICVcQeUW/vr87FIHHwAMriXMQ
jiSVTQbzC3OJeiu8yrtRc8fCZRd9ct+73RmVSNpjP9Vfq5SIX/j6JSXIN6iKUVka
oKhu/vhhT1kUk7xfLptc2NQzzICOnhH5L7ZHPtk8FIKTal0oJaiPJ/hl57aEHDRj
pPPvmk2SJBP//N7URatlripHJD3ZPPo6vld4cOwC3hE03DYo/fwRQZ78HAmA6LOQ
ILjJ5+2/cVuVBWUGgaYjf6Rb91c17an8NB06KddLx2rsP3KpMPcg4X2SJcJvRPt0
fQQK/RVmiKme5RL2a0ol7K42XLVi8dMo1UVPthGapn2klP0LpsIH+6ytq3a/FYl8
5FGNn176atY6Bg456T38y5pElN8UaL7ScdUWIYglwgnZ/Iuda9MqP+0fPvrbDXqq
RUC1djra1TESRqtSJ3IBmKW+VieySaKVELlTthvj9RINHS5WleD669coTfBavcLo
rGIco9qUnBj3di/s340dp6y2PL4IvYmPy7EXLDq2rqEBGz2FgioOhxUv4/2L0inp
USEeDywwscn3tHd7ZNVf+G3Hlag1a651VUUnZbnjbd4etws2wxYiTFpLa5F2qDJ5
Ax/DcvTmOE7Ec5ehm90tbN3HyqEcxzFAXO0BYVCqjtJKG9rlnPSYJMrj6Oi895tu
uMTG26bLYCdlGm7XIzUTL2yMWqEUzvX2yXBwfAO/T7BUkxO/XMN9zwE3pHKQO2f7
jM60TLcTBKXuJwKkxnFHn2R8EmJGpslFbLxs6xRZaY0u9nHeMNATp/5roOsHBMPr
QftTUt1jbdb9cm33updD2QhA02aAhB/8+56WflRnV7Kj33l+zUDmmOAKzAbM8d3b
4MoOZyDcIUAemYYFNzD/8KeZLGQgM/mt04m7LWLU11Hrl/tRVmInUi8msOZTqwNw
m+QjTbhcwQY2ZV0zY+Nm8h2Fw2wZ8hgxn7mLyQL1qjzS/XQWgDDrfVk6/+o/ulnG
cE7PV1BSUW17Vtv3+ABY2h5e0fcc3V6hLX+KZoi/Zq7sNDuzda8/XXAE08I/rvfr
fNVZV+A1iTealBpv3amjdQkAnW53iveRaHXk9z53M14G4nchoi1g726XAp/HbRDi
yBiDLH2LGhO3Z3SIDELgkpe82mmTnimUYeq0l+92J9Ds6/LK/WUeaLj/Rr9x97sb
xb66MOfcgsAL/GznZfWygNEU31ylUeOMkm1TQI3yMc0NyqOJY0oSf/vSNmv639lO
Gff3CAClZ659eL7A/NbxtCNiUgdL22pK+lb/SFhiduO1Y9x8EEWUH2qlXseKJrQB
Ua382uaykC/PptUGcB0BGM3x2AkB1MSeuE+hdku8JG9IhS7tO2ZsCMMYIxDgfQ7j
fadr6QkNVZ1YSZptbI8/b2w0EiW1JCYzVNGJWTrnEqeGrvA9H/w6DI1h48FxwM5H
S/d3escdv8VTHgfkiH7LZnEs1hUkJycZxtfsGsPdX+YbmgyA2iUMfcoSEuRpgfcR
qT5JiFxX8bg8w9VbC1B6yAulBocnuUsIvH8Cdcc9u4k/Bej9Y17n3HAf/BlPxorD
rpDfoAoLySYJ0lHN5XrSY1JsG7AF1oTBkPUAVd9QQP98B9q7KmeIfFi1BrpFa57v
uJd+gSkjz7blKCUA2mnobSsffvZktCk7ebneG4xpBDnIeKAg4UOSKKb/ePpgWcQg
KIxx+mvzGZS7BmLkFBhwFUvzmBmgIFpfZ07ZmoszRDcqvsF+TbNRh6YJj9wwqGpd
OsFQxCY6L1VVOoD/7DRp7qtXSg8O8+QHUxdvdinISs090V9ECwKepibEpYcrlGDt
CsCrXyB2gTE2nTPEKHwrk4T+D4Wh5VWXCBPe/roYC2SkaLG1bkpQLXOoYLbf4xBo
PSO7HkHMnUpI1/md8znzpH95gBCBK9E4BYEHf9mQOp8PuRcY2ZtftJ4j0/XwVw5k
AT+7qyrvNEhFaqmvWq62B2+p6SmkooynILJgEQAxGRb3+aqTRrgUHu5iTDhY4BmM
YwpgCVAxuiLnTFSVgjt7m08oRh65/scTqe+VFZvdxsiBcriHTXXmH6rBS62cd9Sn
tc0aN6mkYiTbjtKKzE7JmqIJWUQQ4X4WdjeTNN6n06sDilGL3d4WQIe3cBA+fWgn
UAC0JoydJ+rPTSr4hLltR6Jeo6VXPRyByH33waB9B+pM05alLvAp6gS7zwu98IVd
CG1F0nPi5iK7Eatbhy/ilnym5za3Ut1y1eYbNlBiMgSGN0BI8J2GU673z1X326jM
3affU4SlCWuTX3kQbQsiA36+0liU/UQbInzahRTEjobUuuBw8yIZhqZsgmQPWks5
dCu06VN5ArfiDU95wtIebJUhV4FqNN9AJPAfP+ZHQo2HBMVNzlsJh064Lb3gwX0g
x8xL/H1gZPTjP9g3tJk2cxai4VgySakuha6JzF6pibU08ab2L/xl2GJjPsVvOVYJ
8XgujbaxnAO7GI2dc9+LeT50cVnB2FT/zPHs8ces+vnJjGvydnZwuvrZLpeWvQAt
tMyMeyD3hN2tSHpObirowKQq5280qhmDinKCE3rjtcQ3aUoxB6dXc38g2mb9RVAp
xeRC2sCHqty+J6IzHc1OMeuQMHxLzalxIGrULBT70c7PIQig+dGSlFvq8atNgTBl
0/XVPCVLKBHjXEJljVrH/GUoMj1ew9UE/bndnqVEPKxxyIqclM/GPwKFJviVDNd5
30gG5NT9UN8+Zu7ZjEPV5FSfaD1MflycwLd/EjqmpKQhkaidH8aJdqCJgd4BA0u1
GT7U0S/+y/rmHueUYa1m5nQRdLK53TrO4Qeu+FkxiBcn6nbQ6dyn/4pea2KmDkss
HNd7U3vz7GXc4z462rNHHiWLrm3lZYGnnmEmtTQ1EC4eAGcI/D9uQGWpLLC9Mx6u
Cy7ahsNxXA/lmUVttExZW7mABEgqBMxwXAuVeuI1Gtz/m2N9Zer9QqrL6IFAyO2y
NSQfVngSGds0eO+oZs3Vwlm+0i1ykaH3UmjFIjvc32wJQEc/RdievfkTfy3rOCa5
aCrlRRXib+7en0BTtgDeFo0vRIU7Nt4dOjoUaLpOagS7DEnYFjkrUIPAS14Nbwz6
+iDvciq0s/ZHTs7e6WI78XtXBTtROU7WQmtRB/T6+ivjBCt+wzGels5mA88Dff4z
9/3P4L/hfF07QAWocPdHeu53lfXioCXjI5ebmFBYABzoaXvxXnKPBsImGd/VW69v
XNmneTTckvcvOL7s2X4HsiWpHWX+hBTpgNKSmbSxu6RjLMMz4ni9XUgoHUyONN7Z
VgMLbF04AlbH98SFYspnQ2Qg7TQfDwOMut1fyAStl4yWErjkhW/vmBvGP9zH+hrz
UODp1zpYGpcJKDB3jJdNvkRT8IcTMgxipZh/TmAf5RD6UatFtBsy8NLtZoTgOaCi
ApD2HImRkgS2Upk/frnh6Ugy+Ka1rUb7aH6c3sGrgUsyCUzisT0/9oeb0eIZo5QK
ByQcZaSxE+UrqKnvjMLIHffb4yTycL3rInIO+pub6Z80qnqfKBbt3/oZ6r6A8SmH
9l6Cz8A0NGFj0mYrnCjX8hEDDeUUTjVbXa2ZJwUQeRY3PqRJMXUfFY1RpOBS4iHU
iK+AUA6XI9DGieaRn8VNviEaVVSRJgGJLwM57MSVUczBQxwbALBZ98ljh5KpHEvt
rhl6mZJ7+gKHKb6T0rok/IjTBmfLOgZ71TIYzQoN0Z85w7+pkkYglGdTplFRsBtz
bB035SfWEkxn0JV26nS35xsja1WbzJ1pIoknEQ6rC4vJ/RfppeTXSWGFd0H3J514
0qFFq9cpUqhemsDbHw11cQq8WhuvTWH8zDZ4eEtoe5fDcZl8ExbZJcX/Q2Kz0zmP
QKFf4ojhpulz/iQs3doareE5XhilG+DxzzA3twjWlmC7AoedEptCScL2+iZlya9U
y/oCYDX67Fh+ubJgJ1vIEq2GDg7x5/bvX7kjWhaQ2/p15Gp3x97msFR0gf63HsVU
j3zXNlxAQ/dSexrRF/+wLYQCyrtVF+zOh4raYAqRhzA4fNpu4gAUSXhMcq64qwCf
iSTVjKKyvxJXjlOlx5NfPcgc7pthPVmNFIQsRVvzRxjYyvedKm7BMgihMOg1GmkO
ENF7NggXmhYrMwMxIo2Bcg==
`protect END_PROTECTED
