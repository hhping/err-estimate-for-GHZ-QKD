`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wS1gK2bW8OxG7J6ts2btw18fuewTUBmdRkEcVuie2odK/XVoDPL0S1upqYK0MsYz
ED44jmslThO4FRdxL0ySYPBTxoAm/htpcIapFvNbXAZQLltWnGli53/rQf2GCflE
ud6M7QMxh+S4dOqYw/fb7lMvpVHxu3oxv11UaXEjULT43LzeqLC8QPxlMF93xQey
etxJQIsgQb7j71bhzA2Qy5d6Fzo0qJTYpKiXhe0j3pPPOoW0MWflvZX67m2os4ff
V4gRNIyW9/SaWFY4HrF542PlSx6Vixyj3msapxwDEqq+4NSgxqT14qholzwv3jIU
ZfQJj4oatLiRPk49xmS5dlGt+tvdgY/Ki+xHmOzBp5HEdFGAgFmg4gzlrwiLAwed
NrT9+Sotqex9js07od1r1UyyMZsvAd0b9wj+P7ng9d0JBWDYpKfWuOSO/SF6YZBI
RdetOT34NeiMV2w69dhfie94p72K6kZZlaDLPTs0vELQKnGfbD11sKPAjJvGExZd
h3IMtl+60KpfWvE/29BaGMP38HVw05ZnET77FTFikgFpHEHYFY95zzdlSDeDrX4u
iuR7gyjLKrCGc+U+NnjZ5znGHNwbe6yKAiR1Al+1c8txacV4is5/fyP/blu0RUZD
oOVgy3rFpgjoM5llcYV3UaQrganqjWID1Ubn1qen+i5AqRRgzlaLA1aLxrj0QpNO
QfNAaCOKEFoNC4Q9H/X+g3z0akljCAJoCJkn8jsrwY1HxAamX5b6NtEwZOwpFPrI
DAQ2zuBZOlk+Fszo9aEW1ymknx2MqoS3OHu3zC1xqrnwj/vKPErv4MKKxkKzBHMf
XpBojHGjii0fgMWIs02X3pE5UXCvUP7arZgyo+fzJp6mqWDo5xvbjffjhTnJB+ff
rPsqBHKz/ah5pdOUxZJMs0LU/8uI+3EycsgKZvzEw1zujNaCqjWh6t6KqYOKAhEQ
M+fSUqXg+5nHniH9otntoTVPhaN3XQU7Y0NxTClhxtbs4zoolJ7CxEegOIfpS9MC
D0JMMRBWT37nvIpSuUsHHETPlwwGtlDPYBHUJHL8dYxY35GJgozbZdq8OHx+vHaJ
U1n/xTQHbiuHl4yFrE2u0G8IF4h1ph/tseB77k9tGBY9gO1VTxTu7JSbZ7C9495s
t6wi18dFUNC+AVkCym/+BX69QRwbZMxFNPUDqbU9vYfaWB5vqEgHtpekBRArBdGu
pFe91Mt69yGSxY7ShhdAsZiDAC1kwjjx32qxvrAbdwYwjDJTyC++olu1QYaq7aDB
t/sd4X6Y62+xofwF+d/5SLK0YBGS0He58nq0VCv9/uv5GKYAImATJ6/Pjhcs+Nt8
pt1U3QEYdcNV7GSACcgL/R2vu+ztAG1xrMoh9ZdBFzW4O1x8NWIpLbRBgClc+Itr
trA0OxQ6nq/zdQYybtH0WLhFPQiND85QhZGIKGW17igqrnTra35NVr2DQQ863fE8
7Wvrou+nLEJkd2cZV1bE4uZ38FkVDk/aUrWvk5CYfqsmOF0b3Ki0NyOGDirt6pSY
4nRCBqqFOBvWbnEI5h+2/jeGjo5b41xMN6Xa/Y+NI7+JseOfgtahhwVW6/vZ3pvW
OE4+gdDMwg1NDyR81XF7GnZkI+HnQrYG+COQFDCdHesWDJcmg3DuxSdBMU2L0Fgc
Lh1QUwu/57h7v2OOrwv7vXwKa9hj3zD6Gp63yDyN4z5KRWLZA299y4mg+qG/5fuL
XbwOEICwIQacsXspoTr7fNjRF7jOn5xbqNCWrvx1LsRJVSEzkgHwfvfhraURMXsk
dmChDZMmBde3Q9Md7uO4Lt1H08tji+irJwQ286j1ZMxcBNWxEnJbd7cKxwy8dVGg
t9l7i800Tg7+DgOoYBEZnEfTZIdWCa1dBi9dZM+KGxOH66VKwov4I6K65l7/cSro
HI6+IVu+uEJvzWdeJisf+c64wXaZR2Yucsr3Pi5mzFOqdpmi7c3hYzFshKIhswkY
YW0eLcfyCe+biNGfW102uw==
`protect END_PROTECTED
