`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/pyoM5dhr47/ct67kIOxcFHspVj5nOfD/0WDqKasCNoc+IhWoN9fHisEGGyKrif7
eaWvr0eq1gwJJ0Nfj7dYF7fB8MypG1KSmVRzzkxCqmHYNFWM2ayvktx6/mOx7bvP
oNpQa/mP9bjqklGdQeniUO3RTm/hC3i50TQV1PDFB819ylTJk6yR2fE2yYWaNvB/
yo7cuKTzAXHHeFX/VTCd/HEiVgj3ptI5wo6S6y2zOQvVLUMRUzY1avvTIovX/TXv
s7D9hnr+gFbdOX7RyEa1+vpInkfbhDbDOb0Mnp7Zag8vSvHgUwnn31ngdC0RLDAI
AZ4g9T9YrrI8i5RwXE9lt1YrnhJrauaMnRhMIGoP62R9xiD6G80KXP85mJjfbtG5
pbyCwN1Y8gnRke6AAMEqdNZ4Dlios/aJWjGKhbkqwl5Hg56DVzeem1U2JrLorGgp
D2CBRLJxAKboKZ2JEutcSW365k61i8YFaqOry2sdLoQijmb1iw8b7nikYbdcvITJ
`protect END_PROTECTED
