`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aDXmsfNrSb58bLmgewAk3z4Oyi4fs16JAmzacGqtuWPZh0+yF6WFhAV8uunHxtNw
uxYQ0+V2yPL1dabaiVxBCgJyDSvhKjor0XY3J8PnbsPUhtrBXk2BoGb43oBc6vOo
+B4Nr2Ud2c3eUXd3Z/ZZQI2BwXZPg6QBiCM/VmW5bCDTQL+xfkfzvpBLA8PNqJno
xUYw6tUU7jcIxo1ocvK521SGQeYIWnR0eR8oTJUI8V2kUOZT8K1FHS1k/BVKYhtk
t+Sftpg01NKu5hI6Fys+my0HzA3rNWeUxHRIghLdUdBN9A8wdDswd2Em6NOhYjXG
Q2HeAE5qaI/fOvRhI/3H6haGmE7vTj3nmIwz5oAdK9tUOgnZ/RP6cfNmyRrtyHXF
Xa87ilFnd2eOKv8yZl6U5O1EVSTYvO5bhmNJiWcTD9abHJfdiDDZlt5spw1Lx9bU
OJ/5WfeKexpxFrwc2k73TLJdHmLjCCNRa0g2zc2isLbJi/1AAvzyTrPJVpETMIlr
zveryDNvUs3bqQCT9QpW27f7zKG8Hadn5x49+KSLvtsvVhzufdYmmlvJZeTHgQwt
/2pVhhy7HYa28nFjENLmHZrw7x173fSP6FkC5agdlfQfs24tCfGRiAPDa5Jncg3+
OeHc2hAyXDkWD3yZtXsM90iB4emA5iiGuXOAsntj2JzVrGa53pHXs0ZWao0opPwW
vu9qfKzDrrbsM+89htWt7kVIxZelO8ObT1JzuF4+Gpc3iYyWg7j2KX0KstB5nk25
vC66s3W/W4bHwIsU6d54ETjTv8N/Wk9G9he+pvTPLYvOPRG5wZLjp0VAXpj4GyoI
/jMgBJpcGIOR4VMhJSD+D4fNrNSw3e9ljDVMkEOqNQRHcVOOsIseMLKJ/Nl82Vvx
Zyuyf8Mxg/GjN6jc0Vre48z1j+/bKlAo1MRP/BVU+/uvKP9qaSeH7paOlLxbqo4o
1Ms09OhVVxkxGc55YwTbLKm2SbQi0yROJyeOQO9jYBGvwuMdh5eIRCucdeLCsCKa
u53Mhc5d9W4mN3DoWszfLYSWeTyftuYhmegGH1650MdPpLUBO4zX/4SvXAWb3Hs/
V2nSvNAxzaOQ+w4K7QUBxccQbklvoOZACSQHiZ478RNh9HRsMbmK771IMmUE3V3L
hiAiUwT4f4rv1RoZoaNrI3jHXd1Uqb8w7+nkn0c4G2dk4n35T5XU8GznjPwsUsUD
cKTKhOXu+L3pS1d+/iBoglctnIXQardGI21Uj13ftGO3XHofl+3W04fXlItY7hOe
+EsVvU8dFo/BlMsZ7a8o9/SsFIDRCBNYGhzVi5IFcNF7BbgEhp3GzciC5g+mU4Ih
`protect END_PROTECTED
