`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6jRVlrveC8g+7ehMvn3ScDiPsYe3otU1XRXq9xalIKFd5EmtKsrTq7ukJxycRigp
l2viJVXUqkm+XpRwYkoR1v0Y4SraFMVPYnAX01dEONRKSfkVXIBn/L65c+42LNQ0
0p47w5s+qFIYAU/sh3FQHWTbKz+oHz7lq/AodkNcVmOf384f1pnA2s6e32DCnJdz
RZ7WmPKZpAq/Wacgn6aAqalEanBFKgVjkYdSjyHyX5BR5NrDUL/N0LvtWbenwx0l
oFhQ4lOOWyAl/usiW5PLIe+wOri4miNlVfd6tO286XHYGBC5y+xqvXHuGOvkjhAb
qeH+VgQV/CAs+X5wjVi3XmX+VOZZYAcsiECbrFEM5Q/1LZC36onZ4H2y7ai439HO
Ez8+Q+PgJzZn3Zq82mklAmL0U1O8LhZZ2ml+cYgKEkRwpOmOIHnkgnCL4AM5T1/e
F/948N+vIw1WdqaIYfohuYGYUkupP2RSSu7LWpI5Q44DvgbsBtyB3PKt+KPBYAlc
HgfFG6kTzPEOYer3s9PdaTYzW8h2nWl8/G9rcmLLrKO1uVzKLstTgTu8vQqS8lTr
PDf3vlvYY2fzeU2s5mB1iBQacDBmEahlCWB+Zgkt71wZc6Pzu+5SYrIKYeKljtsJ
v4ZB575h0ZDU4Lzd3UetHkuNdk3Wl7u+xyQACzNRMhjquYFdw2IbMfg5Jnxz8Xo3
IMFUEX8qIjeCH70047Wl9NPSvOrVRw6Hkz+ewf1r8k4S/kR4yTknz7NmHxB2t6wN
GTriyAaguVkJbWX6u5Pj4ONmpDHJGVF6dVSo+6Y4KhDE5mDyvIHEWnCvRl2SOdlg
Xhd3ur6xBD3fN3mNUiCk4z8aw+LHkVIbUt++BuFCkixbfJDwRjCOT5+qfsBDjvjm
eRp2PU4e7A95F8hsvlvlgEKoX5bhyPGg/jdBHmrTy5cxAdzsz4W6Rxegz6OAKbHo
2ooXy2YNYXaqXRhNoVOU/PMTDc/6rPORCeZQf/Zf2/BF+d/vMjzkHEksEUGq8iXT
6vfsaRoSRcfxjKXUjqoa0DO5bGb61rkQubLetTphOOleg8S2vI7rjg37q938Bh/U
lN1f7ppW1p2lOMtMsuuBliypCXh1L+NTkqlKJ/K2rTSKe9VQLES3ExeT9yRxI7ZG
Gwyzd8qJmfpBk2F1TSvv/sb4onQohl5IfE2CRR2zBUt6eDlr80RUW8W0ZJC/xWMH
oY6lTLXGd1c+5ZhS0bXTIJoQ1jFn8Qb5KtFkRZcI+nFIO1ty5sU/FfLA8RquWQGy
imzMkhcXvCG577RCJFfYK4jeDUB/7kXbra5+KXQotK6Okm62DFH1vzBhEHtCoPiS
B4MUhxiJ0kshQrY6AKAlJJAtUG1LDwvAyQeqbAf1dLlg8uJP2yjdvLn4Q0O/F3fQ
+RkBUkI4uwdke2g4WPqoLjGCflYvesAjCmhTnksLpJIL0crpxq7bxpjgb3c002W7
BYdqADdLBdlXogtI73yv8xX9z1rn4/z26V0PO89l/oc=
`protect END_PROTECTED
