`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
molsJhTucNgJW7IvpKdSdQaLab2fE/As9iT9v+tgaVYyJEjwknWlwDZTKyd20sj4
aUxddI5R3UbrK3gQs3Lvz4RmE52dM/lXE7SRitfdpSfLkUMWI6HAr3kV1Yb7x7YS
V8ohkDmuqccQQ/6XJf563UnmsS6QHIC6DoVlz3J8ZsO5DC0evlA1AhtRrwXUZ/Hy
ZesM4b7KiBXKtS4DMc5zR34YwRz2Ycm7Kcb2GLMklAWpRA4x1cWfb+uMBdtqUFWd
ZAduzi0N2DAvmXPiky12o0JN+/kP1WQDiB46vEKNbR1EpERQSBXu15GApxh8xpm8
Jwjeq+1ruyc5smAUpZjaJQipZ1NnJNcHTjJOWUqe0m7dUZkRtmtnZXAziURlXUSu
ZK8lo4RpS9KFF3Cpd8e2RVvwsnSgpvKFVfcHt9HbNdwd/Kvm0oPiAc2efWEpj+Xj
GwgEcbBsmhO26kx35+3ObF1sZAQrKjxH+WguzNMMZ/JRjmQ7IPutoG+9uXG9Fqcu
guqXDV41Tju4MvDoyR6gp22MivcyVd0pMERIw6/uEwoodejZXpRVTas019GdPXWd
5jbmq3mH8CCSKyj57OF1qQMuPn0iww2R9AsHPeJ/hYpCsNAHwDneuTtT6nkLSB0U
cT+wWBFbH9F84yYXunpu9b3u5T+Bf72ezRTGE/0ZxMgzLEAI0dshZmo0h2krGIxk
4if/Om6e1GFcXqOPpqj8D9edHqg9I/hZDHzUmw75W/CJLtY75zDJzvIWXMzACb+S
`protect END_PROTECTED
