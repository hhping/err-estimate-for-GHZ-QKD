`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7wIAQ6wcLjh6CmibvH6kBvFhg2h+5/1Hfw0GEOmLobC/ToC8q3ofVr034EH8WwpQ
lmRUULUEfJZH+Z8EG2GeJ+acCO/geXp0WN0uixbv9E19mgv5Sl8Wn5or9T7D9BeI
TYEu03p+0DU3ARwK/86KUKAZsA3Tw96pZlPC1WUgeqHLcLS6ALqsuOz9dhlW0chX
k3pO2r1OvbOWbP1TCD15ftad0fSK/F+Qb+UmplGoG2iPyfPtCYTTVXxpNykKIqa7
uYVBR389owgHaUAhqaw0atfkhNrX0V16UpwjMNMJqjZten4OQg9c/ejrYyVsrjYe
2DaMJdJOwp1ystxuv6U+o3yoRYSvuRnICCh5qO1YraVfipKmu3F76EUyEwponoUx
wBcudSviXmZr+072PMieM+DO8e2HMcZ4sCLGJaqdwoxopiwOisK4DL/jwYXi12Tk
LxJETTtMTMls1FGyDu2frnP22gvgxv6L5SPL1yrbuaZ3hH1B07/CDG2ChVYygWSK
oyJaQSGk/mWzRHMdv124kDPkZZtIi1bo67OnULqJRElLoiTaEOOyOHR3zaKzvxBc
26QeaNGdwqottyXHfFY4rgkwzLavDgrWWohAomQ7agsjFWeFb0l18hawpQKqS1g8
bCL87n0UO/OHbvnBZXvLSd/ihtVMsHaBI7fGlDJLHOWON9r3I+58vdeKW+KfbU53
ZlPu0XcUEX+z1v3dsry0c1ilEtb5cqlZNFvLkkis8hFds1FZLlyGWXgucej4WEgi
tD44MHVlKfqfz4mFVdahuemnD9NVadMAcJmeX5awXhiE0Y1R9GydmYl5P/uhes4G
S9A5A+uU7QWFAuCJdnsqqflQYRoiWec1DGmCkpXnEL02pNID6JsnJTGke+Vh2snW
TCCwkBX2vMxcRYzyBNjwIKY9XNvImiR0nx8F1BWbziB0KUWmNT9eqdR4i2OLEzeA
5S+99S5Yh7cA6ZAv62MWemyA+TNnZPGEUVfLE1G7JQ/JPkooNLZf/XgWCwFIlxc4
aHdC4G/A8P6J77QPHz1cB2clPtp3b97WJuUhCA28Cy1NAG8mLkITOOTrBRJtv49O
qT6nZ86ZWIts8+rbdjzZYQE2z/LCEFe9/VFn3cF8GyXt/E9ZvBWN+m+yl+zVht9O
cgkLTUFQAgs+XLdCh6MPjg7NRorie5MpAV4Ykdys2FUWA4O3YHv5oDZuwyf7miAG
xvtToDq0Wkvg3RrWqUCYRsLSEIDvNkRTnyUCfYnbvtph45KilnPUg+p7zJ9AXgx2
Z3b2s4NJ24LX+B0rNXrqOcF4tX8nLB3o0hP2WuQnTfPqUDlb4kRxCOmyZY2BKzHx
Ci6Eb2KDgCAJkBpmMVVJdo2txI7U+DIDam5Mhap0qjCmHY8AEmXSuQvgYh76jpEl
aax0yeT0jIKxrm0HQVR4QBhYeaSljCqFw632JD3/eXhiyosEL/Y/PChOZ4muAHQ3
6ZBX9xUMMBEkBi1ZvTzj3xdE6jq6VRVFD+VtxKXr6OcHTpRIS7nDSGEJPvzzE25E
jQdcpBmy66Iv4wpAH/8BS13RMhozo+pCOHKkb9Sq9WHaMhENeKayv3aSF56FSuBO
2CJOgiPYObN1gcH3Jp+OSrec6dFh52zbTYOOiMGQmdwhaXmMUz784by8GL+AqvoJ
JOrVo95rhAYHC0NVMAsV6OEYZ8kJH+AnnsaOcWfYDr+v7Q67ZsOCl8tTP3tRvul/
HWRK+IhOMFaEG2yK2uUHHrgNkAn9BFMLHcCiYUvo8NGvmrr8R7E/7fu5fiv9EUyN
P2l7xfRpOqgBOlGuEHe2STTxRTFZ7+Hc/rzzX8IWgAABF2wmCAe6YdaTeT43s1XS
BB+igolvnFbVS7pV1l6yHh9Iern9y70r+I+ELUOLy9bAvjv6RQVdqu/t3MIKrPW7
TowtJO+Qupj/O9hqLdbeaCNYepjs/Y35HP+0IpXL7/HSxWvklimtu2/a/v5XSMZP
2DLTdIwx/9VSTk2IZQhlnWNvF1AyrKY9nwGEpB2m3KLbbLwjcWSQVTmFJUx/KUFr
5DzXzEKo+sKeci8OrwNEncpjuOqh8hVtCe/U7azxPLVLTN8fvQYJ4njmdyZLt2+j
w0EArVekTDGdp+/cnxxTeTOJ/bWnRKBz4JBQNIKjwUOgUuIxDMQ3Leb+JplmkOQy
Sgi/UHQC2FT6gYztqFW6pV0ec7OuG7tzhqFGlQGL6UGazIfYS2PC/l5n2WEB5/px
6mN6q8eyBq+fs7I87CLHSMjrHfLucY54vX7p4/RCXrCI9UbO/RHRkPzpMv1Jn8BN
0NmIUk5+mk3VVAmTrsGZqDLmqLUCmoKYXc0egwsBOI1uVTXUO6aTt0CLATz6MKxc
cCUQFNREtHs9yrqiuc2zcVmn5HwBVNFMEPpATPmtONWDZq+vel2k/wFw4p3TOLpc
sIAMipj7/Nj/1nXDUx9BiftaQaoha+lmFI5WUvmYdFzzQOAeB40uXBrkFfZ3WIcI
Foy74viZWR2R8ztHxg60AR7k7hrehbjuU78Ag1woHJ55M/f30eyQQA1rpq5lJKwq
4cnmlVXMYkAicMvwRizkyGyLVzKP0tnWeggVDz6MZF96htqu9fW3uuqRSByHrjDk
W8ddylKQI2+VRGObHtUUpfqscD6y5WLDSNbNy6sjvNXbYuIFTkDRB7aTJ3daB6Sv
3AOTfqe3s+yPkKOc+DdQmwKKo7zAtor94kDUfj7fpMq+SeJF/FuK61SHY9vtn/AZ
9NB8S5Lon8Dcvx6wEYev+3OUSYj9mXiph6hBoQ0rMH9SJyxr/J8ZHLBgKG5Ud//3
CQh0u/QeolFT8PSIAfNCFBpvOZ53R8KAtKJMh2YDoOPpW/sUgUHssRmPPxJ5FIE+
ZKujXlZg8f81zHcC9erqG/Lf1e6EJAIY6UfOg0M8a3HEEJ8HFJqNSr+obsu7pWRu
2fjLpBfhTkK1oV/1x4yWzBhEylikgFKgcQjh41gdkPYS5LazvCHy0y/SPXHZWnBm
5S8FuAJuyRKdYuVCu7Y9JuVRpwjwYCIlUrcqTUatuUdIgHdxp/MQfMeon67qJ4Nh
I9eSVZ504BuWfE0E+jr8idHSusVb15RTkwjEkBlPEWXj6DeRzO2i7Dw+5dTezFl4
t7Wu4oDGSrb2YWVQhktrko/U7anUyVHGv1XLu4AQaDUDXBFmj4O+jUrlv+Iru4ol
W2ZxwOpKssaUF6IaCb2M9RiccrGiNAZmgOWtD+c1Bfzszbf0yGuR98uY4UFptLC7
skxEvxFdtcvgJhoR6rPD/h0HFHqGAeV53BUX8mBOa6WvPQpqhRA/fWQPlzqA1S9Q
ll9r54O6O4sfgRyGYkkPmUDFNj9yy87bIgj96zKnnF4JA4iLl5GFIZ2I1AQuVmAM
QmspZ0PR1MECj0uFFx1b/bhYdgMa1TAm75KI01VdZj5aZ2+Lnq8JZ15cuwirb8CR
/NNqwWC3OJxKUNTObtHhK6Rd2YrHasKh2FqZkktDI1lI1DzFr2FJz7c9Wur/shAW
Rvgntovf48+C6SNDjjGxL+lXImFvN37LMjsvdz8TswqnjkCfeBpU4q4r7QnOuNEo
QOOBiNIiESUoadY9hVd149LA/JrBqsfBF4WQsqj+RX4yeADNWfMHa8NJvbf++6ec
PUWkycO4WnNk1HVfa+seYM7oCTN6BX9RDFwy+rvX5pD7c6VocQaxsycm7/GdAiZW
bnci9D2dARmj4O1hR44sZ7HT0T6eqJpxt+7z/Fqxw5dQqHMWC1ew1/oeoOPI+41u
CCarMOEcWK5VRX74PXbO1iPBklPyFtBmZtFv5mhBHktdL1ceGwtIl6xnNJQhNnTL
HFmFrgkGdqD/8fFZ7jqsT8RGXyKF76xQ6+Z2rYxtpYhTZDo3mD01Rpa366FNtLS5
VI2WMy2vOHgwSgJF/BLbhcXPRzOBrztLDGH4hfrTb0Nb9g0QZXpNbl7L6WQuVlZO
Cc13LatLBSnNOBVdKWbKo6cYFF39sXrzW3SKDgW2LhHqEsrVsQmPuAhoFzhrKnZd
Z8R5g79TWpD/rS88AZOEGRLZI/eAdScCQW9ChQmGL5v5CzQfa93+t2+OL9B9vcvv
Cttekq4gY0uLsVYoSIRtu2a/RWoxQztxckgIyZCrY6otDCBFiWNJQP7GDDa41uqO
JPg/9edbisNz1QTXobvIUlyePzfRVxt6fNE5eZN/UDpR+3pYlXUo7DZFKN9hs+Hc
0Ss+cHnikoL8O1F0VR8MR2dxuWN9ce0EpthAJ1GxxcVUHiGQC19BG3y/yltR1PKA
f+SfORWmXtsjyffyV5tl7CUAgD6AZ40ZJVKzrDwqqPCHD7pw9IAExDaHukVSAQwp
45nvJuRset3HV2rAP7jVuKgHuMyN0HAidhOOCzSAzmjs130eKdpNIJGZFzEP0EI3
+KFnOVUZkejPq84evOL+t6a8mKLzKQlftL7q6+IWoFomBL4fxo+//JoniTroH7sf
jAudYjBI2/mguzw/D2pK2VgioD1G075ZM3/tFSfOixAV4pm5LCsfv9rKubEMXdd7
6ciPY78aYiMG4WHIiPBUYP4sEixDEVznP/owGOKtz2/EeQT2RXCh56sKh7SCR9bV
4VRSlJk9g2fzJz35x85BMic3KbqeAwj2anmDcc8Lg1OhZvtYBSaHfLjcZow82xNo
FvxrAt//+KwLT6tbFdZBkXqoXVpJ+VGaWXYmOwQkQopyHLt2uAkCbvsCFAoDD4/Y
/yktGbtmuq3ygKbZpIyOHi6h0IFu/Fpo2YH33VR+cUjoIwX5K+y9Wed6gk6UUjDz
QULywpf5YT0IwJLloSx+nmES9ONo/frXuPzn9E9nbsTcMqq8fx9hWWbeLV99lc7W
dY4qP5Y8kW2EgQNxGhjGgiuyGDLpZpV2QlkbTL6xpUXY/C+w/nW6NFpTZDoCpMGd
D/5MbNdues1WSVvMuIcXib/bWrTtyMduJMKW4EpF0q4mggdSIcl5L4qZrvy9Sxyj
V0fdJZar8rF0ICZgHdarQmvTA8HAYNsh4IMCUJXzz3Iza7fLU3eIWHegVwfCVMnV
XTsDfxb/i5/S5Bdgg6wl69/rOs9oxTZqhMbqp+DWdXl5k3xh9Xj7Od5F6S5Mf5hr
6KVsLuRWn7GkuWPE3wMEhegpKwhml8kPmEBm4/iyqbbrLIN/Spx/mM+6ZvNWmkoq
rqeIJ8ViW8QoYYUxa4POrHT7DNshoHdqvR0+dWIrxfIwPfePS4TcxO537JggJmKe
sDI25f1BRmi936Gj+xxmhhnuMFDpwW3MEqUr+bkEqVctUpf9WRFqyj8c3nEyCuvt
SZ3ST+t6cXncqDgTsymAS7W4FqFLzF0uUV2es5Pww9lF7NflTzAZZGUB1EAhH9IN
Z1sESe4EbTEp8hdcw0d8u7YHw9Yjd10RBRywcgmMWIKL/uDQtDf7qqXj8dxfBiSm
PhINmSSTejpRxyTKwrLkmARqzQqM/61/BwaBqu5kAd3tNHgaTv0766Lw9p2e5VSv
IgCShwA/VJyYAxfYUH2tpdwpyxEDR0W/LQd4bFHz6znRU8nhtvHxdL22/uQN9Yxq
NoHRZ2IgUwRIACdJXWc1ubVQHFExgB1R4YDI34sYyHLy2IpbjLg8vn9r4BhYP1nI
XyAhx7QrxqVHDB7KRR0lUe3hFqHiO9ntDPf9lsA0w2a0BihvsdtFv9hPctRvwVLW
uyz4dKwc8/Q7P6T+/C7TN3HeVoq9JNTTbZPdryV1J3iv5kpCNRlBVu0nLE8AXtZX
GQctHPS3uuw05OP4mL69XIPIYw1UXs7sv0tZfH9ZBuBorbnDusco7k93RtSE2R0H
VqIHepXxPYhw8GE3A4p9B/B3jWT0znVlVoG9ZFpuFfsoRwlRPgj4gl8QX7FRm9ul
r2iZmBSuwb7IkPzcpdUSTfXyKheAHPIP+Z9IUzdOSZOUa7xmN8o7DGwEv++2DuLG
UtuE2s9efstTK+A8PTJ17LbwHgRXyqyK1STQ5aGZ4i4R6izBPLCXaphD2ysk0Tml
FX2FbgqCAPEjzyj/oSIHPAg5oRMPcVLN7GxUaxj639HHnNvcyEZwhvWub11Fjfzq
WxuenkZQMMPmJWrJESaYLm1uAS65F3d9wND2/UId91KA8DsBhyByNGN1GZqB5tC5
Ual4WL9p+1CMfRTv8H0a2AIiw9TQmsr2u78OXOM4DfhYJqXweXtR5ywifMMSHl14
l9Vdz+f1Nn9tvvuxiJaa4cb1ywEUuk3L65lWd+Usqi1OTrxuVsMz2j9hYTIzswSd
IZWhSFQPsOBAVZSk65bf9n+JJ4GwBLKXJSZ7S36Vrid8ZZeyy+9bPsRCb44t99DI
lm6NVEChGDv4V4iKJUcq0iDGy537PDhC0Hz5Ghjo4IcjynE83QQLQNzQtLom3l4l
3519lusLXoAPMnZvRhxf/nHI1F7q0kVEFX/WJ2d0hdDmA4cKG7XP/zelUu4TnxLh
hM7sYc+I0/iHiQ7aJCZCvadXeJ3ar4H66C06i5Vdt4AMFfB/aMZWPRnOuWdturnn
MwGizhF/Vyzfw+CSJGZBNy69irzoxu5aLg7ac3L1bWLongzYyIPfl/H1QuAMor9c
D52KTfPtjl+V+89BkuMKxAqnZvRYZ+eCPO56HnEH1flxYTMZLCaZKWH0kuT8FHt3
KyW398PpinFOvM9QOrSOG+FXLhOKVHtSWbXt6NgaJqo8F7nFqJHbdQJXCLV5bzpI
NXeWzxzLf1auXdgIwnzVYJKMVWX6glPjAWU82/efH5ePArzwlGhwXf81c7Iin7m2
fpp+egiUb9gaaqcKY0X0j6DDzjy9UHtcFIGEHTWLOISDa5pLsdhhi0+CRDu0Aqea
aD0AfJGfIxx3qqXulUOoaHCJuztERQAv+SrugdUnYKqMaz5eDOYirUrvqfZISrjr
Tncj4WrsPBV0Tp3UE4VrS8xOwMTukOZXR6sMs7SRM9VvGZX8jPJp0EubSVAyUF/h
Sd8M9kAhAC1Jidog/SvaVhl7iApAxxTvGKn5nLLas+T1FqaEhx+uf+Iczv8H7jTz
81eOMkcEmCyy+t1zFP4G2A4Gxt8ZVOSMsTkFWb1+2lsK5s6e0FhU7fbnX77vXTG2
bbwabwO1NzGCkDFq+h/TZwZXidguavAsL1V3Ls5suT4ObtLgxVWdcHhMhd8SKsaD
4dh27NdmttYTSXXTyS4DfJ09IwdXQ3Q5koyJpiYljpTT6/RXDrKhu5nEo1VzDcVO
HX8JCOytBcrymk8e6R9Llm2ivJY8QxWaXz4x4OkQl74KehUlW64BSdfozcJR7e8l
HKz8m7osK0sUdlzMGjSeTVFmj9FQB+qYEHieB6kI9thwStWSulVZbi0tWB0yhuHW
cLyZxCDUF84mVTPl8kf9WLpeUtG6rUFDxCQjfDKJO94EbGUdAxar6u9LiH0zGVQz
Uqlym8drXF7BUc0kR8LyYVh7J3nmOyk1eoS1GENkrGVMkra21/9GZtNlmZYx9aFa
CHHO5WLpjvYaJCM7cqgAfRQeRTSo0SJuqUUn1Ek2634Wo8Pbf7q13CnXG+Z2RoCE
fM6LVR3Utsd6C7yHuRAd1iYZcsA+A93qYUVlE0pFquuBImXjkMJOoIzMDaqBBtf9
PW2P+BfXprmtlVmjiAHSUETOmUFXBoAhiTE6At+NTXxKqboYCNBGfvHa4Sq7ezA5
UnoYI1sEFafEmr4Yyll91vP/wRzwbcHd8hOb8cmEEvTg/1TvuhTdAZCiSrw9ztI0
oYSS70Onga2XFWAfJchCAUxTZg3uxbXLgUgB08nzuyPSI5m8DNMr+dHoVqp4w+Sd
ZRBAHX+mVqWLE7CrrdVfmBqxJEbtIDiivDwPBtGKq8nOuNWSabSDXYDH178HmEOs
cbH4ACA0beYxL5zvq+UU6nGDEH8eJNN9CuMEnBo2T10RSatLhfUtZVMEkjzNOPaE
1DWE/wzixkXgKzjR4YEByIc2ZHAb3ZxGQgmU57xS1JQA1to4TwrjZ7dGUkIcYylO
OcxKxOKNC4tuSeriqgtfkrBfa5zDcGL7NLaR9ANKonGCQe7o2AHjTYh3VvdUfWgC
K/LOWCz/M+B6OK7UBwzVRjtfk2z/C9YVpP2527u1l5MHLFWY7NTiTfrxnU/ljINd
sbpqGk6MyUru2Pz5BAsZGHtNfR/EdYDiVXmiWuspaPL6qsB9lw24Pb7PbVg41gNj
65x7MOXJHEjuwY4PZHl3vRtCax+mlJINMM7hcpQO2piBQ4unGp2BNMd/OnvHLt4T
+IDi0DJ6V/tKszRIk6NByVaTaR5Y7wP/4egQTV23HHXPkD4hJadFYsg/2FAgWX0U
B/0RPjhhRajXOGj+V0FLGCjoCY5+MjwuGCnIiUUVf4ZO/fvF908u5W54UowFT1KJ
dMdl8iIQcXb+z8LGaX/Aia3j2wegxybUUUoRW40kfQD5fC/iQEZRqJ9ZYFaZsKYo
gJEz2aUyOzyKeUpsRyFMsrOBfFG7J3XnMGt26AWwqYQ3CXfZs4baaa/XCfmCn3lZ
xDyBnzp2oQVCGzcjS5ouvYHFte7cJJhDLnnrP/nZlcH4mwg/mmB9SclMmOHyFIxy
mUqzrsZFeQ3crLdIkFosLjvg6iECm9xJGSUoK8Umiu1bLI1Wj0RaB2T3KOJBe+NT
58FSGIvB5L1Lb10+TS98dlkK428vJAB0sIxqJJhBteXcMzHo4GWAS0i03m1r5LiV
fAIycaODXrs2AMk6djD6cXHmTzYmISScO+hv2DOVgey2igkxOloPM+kQtfO6Io2D
384Gmk1qa6KRR8tPtJgKOBcrfEnTMiUivwa/7tkfb1qHAJML+hU2YyZIFwkhmNgd
LPXsv5pnIXlW/ICJ96naAHkC8zX3Zr/0FRE/OhhA3S/w8quAntVNUvbasf+bVoPK
fdTCRVPrLPsOMVtmXJ5q+mxrm4yTQTXOSPs0B/6roXpZyZcGVPFv0SWJ90qfSNgQ
doywpAAw+6qZzJfpJ7eJFlWLQG6pmOrca58i/Sk/XlrpFHNgwDrF10OiAXQqJv2/
jZT5wvmqVcMXCnLgMIAb44m71m/NRf/B5KWUpgcXOH88UIDKl8DMsLK4WRifwSjX
rrr2IsjnTJPqV5TV1TrTePpJjPO3YZIoi0ncp28s0jv9/kDks6qOLdMaSutnjz/k
zcqcGYhjYrvsUIgU7SDyWzU3P2tGXLA4beZ/uGfjUocrAuF9LBB2eVTucBXboVg/
1nr7+8qVIKR1yyn0O7u7etG7WqHN/Y0EEQx0g3p1HTPy4f/MoDECL2dl0wzOo014
OOjiugbm8jZcxrzGUaur4Pzl3lbxjebbVnBlKkkVb0xLGXatqB6XZcGzyHHiB+Gm
PISLl9r8jhuSKEXeMyX6/ybvkvTCHkxABC0FluV29984ZnALHeACoHO30wC06KlL
BqwTdMENwg3WvKLESQDdIaNJEVP7ihbzbjkAWKT1d2ZagYlirJn63HTpBDXYykGJ
ZELgPXyTE7bIzytrpSnP//oL10D36PiNZzSHdtsIebfdMwXjt+tSAUBIoXx3RbA0
ikzi7f2kxzolluWEZvEhf//1O/Lo/SVW7HhBnWy67ufNBjeZ3aiXKTZZ6chxiKZG
OzURaMu3BjWJW1DnpIMsSnBk6iS6QcVzZz5Bm4PUvgsnEWxH/+3/M+BTYt3LRpeX
94kngekqUnoGt/6NR3JDJfaRwaKOCYbkmfRN9mnpOTC+oHno2dIkgsKOlrQFxDrs
ApP+02N9Uie11fIUbpLrFPzCkpzz+XKgRzDpa5Ey2dkbCiQ9HJT8Bdu3mfJwtc5t
sptFxBw6Dr6NjtJ5R2/xGe7L6PUqx6E19WMApBsm/G+shkUu87x4mpTvclonoUjq
aNJS+Fn8mm+xhURGru6hhR0mzGOChbpnn2bt8DBWXD92+MEVy5JvrVdXZz/o5T1b
trIG1lSbcT7VrHfJlA449k3JNfQUyeb/qJnOFc75VpX8iR0Xirw0Fc1iGWaIVm2K
oSUZvR4SVMdVxEy84SP7fFy4w7C4r9fElJjrA7XROOFcAzYaQAwgJ9cQuC3jIYGV
JoEPGtRWTS94oF59OV6onieFSz9klvHIDpImMUsAhuLAx1vdnz36e5lhDoNuFE6u
vgbRg3310FadydLU6m77Rsm1AfJYVANP3YsbGIqlzjpVCvj9mHWT7nBO4fnlWlAp
pbmtfCRWrgx7YMGkvJwH77ez651dH8pZ96ulHxrzBM3L9ulxcOOGbY8jwE8CNCMS
EWKTHWCa9cIiEN2/hbM8Lkz6Z1oni8gOAmkrMDvCjVd7ZTJO4Ea7CGSrEAHTge1M
AH8JCagpiSPT6LFsufCeFqEXA8qpUp/EvbeUQl+yoevDzG53eHpULug9Rn4AWvlY
K5sWTiMCrbtnsprXfAIXkr6wsbVqC2J52+hE0K5NDCmn51xeHOvATFzuB2oA8+2y
+LW+2y/UfxqowsxtKs7Ibe2AgrS8uLaGHPM1540SRl4ik8HX4SLUVQB+L6pERWyu
YanUkUN9rhmiZJgitB2ORYtY1j96Rc8w2D0PI74Ww4WAZ7Dbx5PPvhtGqkUMdL//
3nBcUqTgiQog+jAZ+mNdlQm8HtKPj6r4uB4MDIpYsxCJ6KwFRLgQfbO2wBBZ8JG/
vKOtkzMPm53xU2x18+fXsUW3ImsSX4jkHvAjrJGwFNGhrwl7gDgmIia+Pbyw7Aus
MBpCbjW1AHy3pu31J80RT/cKfImePdiBiYrTvrbyPXpqBvm6oGRBgoRYWT170AS1
EzljxZneAmbSJw0M+CJMd3E8xflcztCWbrtV9p4KPUCtdTj7VM8FFtBnGEVnfUo4
9i+alE/WSokTC540rKnZf7iHH+sMqjBxCctbS5YX26RPdxYgISJ5d3KDuumeuTtn
7rlNngrtEHakfLIYjREs/cy4MzkpnpuRGOxrr4czrl5ycMNZntOr48rbATfwDTuK
OjYNhF5SYtHbuaK79Me2VBA3rGbR9M5espKYMchYsCCU6+uvwb2OrbdagyZqtCWF
lwoKXxNiyOXxhc2Ov/M/qy3UNYKvCFWYfYWO4GdHJuUwowmUqJrLeI3L1UcF5Fih
K0/UbeEzWJMOdMxI6+8wps1Bgm7xSY8D8F04Vw6swtWEvMTHt8Vlg4yQCqZZdaeP
DVTJO084BIIabWF9xJbiP+1vYIAPPwvKsyRHUPni/5HGEDbJK4lzOomKT9KLd6JE
TzNh2/wwvi3QmjSRBkgz1dBDDNySUkIiSWHso329vT39g6bmPLd98V3AOLtuDvuK
yP+M8r7i21rKZD229gqlvZKzXcSxcYPPlXwWx69uw9XGFohLQWNfMAPxPculiiiL
nTNGwSaRvatye6jDpaBvxjVlfHg70Cm7r079xpeg7poPd+eMWyfMDOo4OECy1l4v
g4I1oz6wXLGxXooJncflrTw2y6xzle26KpNTel7+t+W+tqaAqP8blbPbqkH76DnS
fyhrDQIehWGFayRvQ0IgYasWFkOgUGoGT08kjLOcWV3nov6531A+R0553kFih0uN
pI9MyB00vi/QICUBydGZBsJa4bRWifD+w5Ef9P/RGb/GxPO7Iq4Nxu+asVrCKREf
mYXUB8OEnCTnh89xD9pvfmVt032B26r2m9WGh1YfvzRrlipAj3am/lnzHzXLjqNX
J+zu29gf9oorLonaSZi7Mk7BlVIrERy+zRN8W/moJkzzPaNl1HJDZwntvBFZHzIt
duozAbfwmRbvbwKKg40suARlHetbCaUThZvhLFffrSgaNahTLgHZXIfjhl3z4L7b
iLDNYsYCd3YvEb7byzCtPfenh340lkZHi8GgB+EGsQ5gvkDEtgH92vF2U+ozOa0K
5jjyxNcGWyOgzAt6guOQawbG8g9mFqShp5u1+rfYQiG/hsPZq4q4qAeXxLQRS7Mr
U7zDob1yldRM4jba0/1VQ+sSJD0kIuAMljQ4Bay6mB5ilI+64c0On9tchpEx2Ssw
jWpxwsLjHtvP0ZSZe8+4lo2XsSuK8SxNmiDtl4lgiJR/8+MgZyKu63Ng53okfX7N
pUlU5bh+MJOTueTUcPxpihrYo0d13eGB3woQuh6NFBiK4+63l5HGCbuBu8cUlnde
kvQgilxTfzThc0HS5YE1RGCE6uIosvAWTD+4i7hdDB7GxbUGVe0u8L/iyi7wO8dw
npPZB3xdnIca+nZClWsnVolAdTAoDmkhCxMNVSgo2Sl1N32/wDh+HKXK9TiJa47P
p53gWPA4cLBdQJyoY6LHsp+BaQLfJbjUD/aEg/VXGHH9abtKtHChPQVVunnxfPAg
+dRkD3i7pJIpizMBzupTUKMRdlHj0jfAgg5k/z7WDIZOGyCncEpEvs6BvAzGSP+T
/4Xu1eUzdtT223abzaWfqGK36x1a4hM8MOVu8SJFZdeJEDmNUO8u752XhvUYhmqf
J1lkqFWyhCiYjj/JYgzk8vY6ZRtLt4Spr1EPXzt5/7bNpwY70ivLqEmYhXd+8rAS
NcgIv7l+shkaUrRmuMCaHbxdekLW0/GaOKW/3y3lGTCp2KltI6dmNECEYbrjL97i
h2Y6f/MiLhGDuxtlzoWZXnRKBmBSHMiptn/dbQ12k4ol4vFiY6v8Rcm8vZDryIdu
sAVOqW4bulR7yW4+uUsx2HJOJk4WZPesRVoVHvKGOPv2ko/RpXZT+rCIpUsuUY4C
jqaj8TyvLHgi5FTDvPTTwdGkgr+Pl2lPgwiKFO2FFI1gKGkJBkI5A9mE+rDu7dv8
AgPV3mqE5zpjZbSDrd+Yf/0qXAChxQalPyUt1iLwBls38y4rCXKu5XrzQyGpqxJ3
on5NfUXQncHSnWqe7svnxDgdQ1EfKsjGbw5kFmSGbGHJuLW3ZkXMeRbvKZEx3vZW
lZqz9qkriODBjxVIRZdrPd2u1Tsb3Zs7rL+irBzgYgXwRDYlJ9D3hWFaaJRtUvmH
tE9LP+uuDJjuBidR1jIXyF89NUuCNXY84vwFXYYRJVDshWJiZQwgBxl9RV2fuvqH
GoQGMnRoOdZ1oTbzVBzdj80ylPg/UDJd3c0Lfl6YCFNLdiUqH42rXsjKws5RzA32
6yAEV6B7TkgOSRejQdH7nFhFUOhl9nBEwb56PFIfXsnl975oavw9Q43zudZME+1q
IArzTmq69ZG1xRFtL03VVt9RJFP84wvdDIizhM90PFQa7UI5hDRBob2yssrh8ebF
IDI4lHx6kEBPfrmYZYHDpZEzB6skR1t6/mk+V3Jcq2pPMxuER6Wj17lLNrtI1B1g
C1Flrv9bScAwhDL3qoHjGpqyc10Mkh5AprbTHoG2A+G8Hqv9qGXGIBZQAxR0FdU0
4stiLrg3hZXvOZpwJcMnplyiUXGj9WcRHv12XZtLvL3q8EGHkoQPmWtJr2GoUN4y
k8/iXAvCI8UGbEHCt+DUTuHGzyH6u7XONcWEPVGkx4nZERGHWdYibnbDDrW8vcK2
kJvjZ8n9tOveA+4SsIOZmuot/8wDi7jqNnCrTfMDCmwkQphToh7pN97sZnyahBmu
jchhcl8GpxKMd1yb3+iIlOJ/6RS9BmPYBNbdjZjrmHWBmoUpcUT1zL82B+8yYkjW
zgiU7VHgmoyHsdSyCDOn99qHwao1yWZLOH9vt2TFbRKy31msllIzTkBN2f5kCFFs
1M9i68oWnXwiQZHAazDKoLnxHi8r9K0gPwmTEkFvcw4hXy0fMRmApdBGiVpDnUvi
QrtdT7WM7SjcK0u+XH4ixknAvxkek6OSHahMoXKV76IpYqNPkBPcPeaJFQSc79Lg
uwKljWl6qtaDPvgoKozAe6wsnjFaCXa1Jh1XPj8d8rTJnn2m85oLI/VRDRqzkOm7
/WUOBGdS2RfRi0YqqlEQbYf8bLZgX+ioF5G4xKcNBBQxmKj40XT02Lfvk2+A5s2v
TvvM88OBR4bJPhxYdv83rj8GoW7GG4j+HwQLY8PwoxK+WEvhz9WwFfeQhOvHdK9X
vaU/40pfQyd80WJ1NL4zEnZNGIhNQh6nM5AYQPMZRM+8zcY/xvpyk/VVw32D1iTe
f4seJDU1X8dEX766JwoZZ/5qnAusZKCy66XCW5PPKbsa7neYXWpjiWIzZm5MihLB
mCGhLB50QdtGGrhJBzswESRF7ZGs8DJcAvrffMzd13pDfYn+dlnF5+3Yr2tMXmkV
TX4/0zsbcQ52CAA4+SbBM+NUQC0h1dojv7YXK3IJ982Cnz9meyRj04CDSmYdIDoh
xVY9KwXjNuXjpFWjBFWdIzC7Kg3wQY+JrrPOxm3/c6gTCRlKxyKvPBU67gDKQly/
nb9HAgTti4UwOP3CCOSKWN3GbTrXIfrXj3q6IQM/v45lUaFZ2kFaeHO899DiliZM
p7NVYc4BTH34qucUSHU03npT+vtYQ8EemtiO6ZAfAqs8sXegi6WOsI5lWTnWmvZC
JXx+nOffI9U/LWQ/t6glOif+BBnqVzyFWkWhsMQgRnJLIitMaVwI9e7Y2gB0wv+Z
ojCr6DUUTomlhzMH6wR3J+ODPqBYKc6MNvky/GCb1RytZaMgTonVCiDoPOYBAxVt
UDNuuDNKjydigxo7IGJ67eyLk1i4FtA9teFEPEcSNiz+ZwuWZyN6KQk7jHdYKAH/
gVeV5XIIbeyc6aNzkbJ4zxWYviQ1GfkV2s0Ec1btiYgwBIN77xtnAZtO+k5rjfwn
jK+sf7MUJMQkaRtJ22cIkurFW9DUtu+m0uvs1Dqpr7kt0PqmNAFBnxAFiEZ3YNGq
bGpPMUdRb/rTSye8Cb6wTcdpGFb8CFPKIO6wmXOhSeObLTmAUcvYTwOpHsWv3DqG
6pfCJ0sggS5tb6/IUws+ZhZI/pJ8txqcESNnbmffOuYwqQNiRQm8GtNXAaiQI7C7
GfLiRsDXeQNjMcbs74QS5Y5pZ+QeE1jHOfy7Lp0iBOPjJ6iS8oj0pUzRd7ZPShuY
GKBKahhywPeFIvVW1c6bGHqNsHjYzaz9qHzPEzAsT5QjfZQYnK7zYA8yN+/XCJPs
4Bd8syPwIx5MGy4ylU5oMzvL6CXly4o2IMsNKHh8q18kgTfxdH1mClviISnmG+W/
StdiiXMPknArvisi/kJao/KLZZLS/iwzZTAVeCwfcpimKAmDJQqpJlckSNWT3LOL
2oU1UlUjJXj3gYaj/Onop2xsJMLnbkGzI6vAPKZUigGdCJT5fRS3eZIGwl8VADl+
cLxBZj+6JZochPIy3dBtzV5TBc0DIJhwFoRpI3y7EKjBJi8xuxPRFNQ/NHcP9JWl
dOQqeRAnnZ6n/lujZXTYsNdsUABxFeeLxIO89aWKN4angsKhHuyHkC4ydiZvgpQX
aCRUuPRwHPtSx9bmL8wLixSvbiG54cYw5yESoNGuNn5PoeSECTgpyBbNnmtTxObw
ZqIKxoZaieYWfCBxx2Rlx7VvVygt9075Lo6o6Xm4MxcFlkv5cbmS4A/pR+jjul84
AoFeH8LcvJH2E8bxwk2AI7oxgtaZ+/HRMwLU4DIKdoHRjuzCzSmG1FsUOWiSiuv3
1IdB2jQzu7brtW8s1lZVMqTqg+Tv296QKiEFeB+zBmDXMACw9ktNfHTHZYgjA+Bk
vg6lGAbDZiA26jdT6LNqpeYkx8sBtfvA2xPRSXm+DcpD8JH/FbJpiRcYVt4KhMuS
mt3cqig0zITgz4WWXlH/cS6B9n3EdVI3DbkLDTzejZVjT97/fthkAuXp+gntRVgn
kqdKr6NPENRoaIubp/LK87DVCmm2mG0HSNAep15rU3Rz6BbmSp4YbEMc0YQg81zJ
zc5AynRJRCMSqcmbBesyWlY4LMNPKwBJ8feGZIYBcuY72lqrMaobPOLyDxHSYWI3
ADpU5LRR5xRah+N8I++ghWBmMQoyB9fAQDHKo5SD3olqbKj6PlT3MADn5MrmxWfv
W80sd8cG17dYnMrwEXW0d2v/Aln1ZO7fpCERQCFph+nwRAghotv/Jqa7HTYbg78k
hCUrc+JhBrttLxBOV/zPbOqkuKs3bW8Iq0XSSzv1zrGx1rrdiAxGZb1DBcNDSfOl
9s7ip6Jhp0ntJHYXaswXFjh0abGFZ03RL6AHM87hZwXaW6lbAF+E08vlrVE8TbVM
Z8yeAVOcVFY8O84+s893Mv0FNAKq34i2W10/pof/3v2CPU+P8x7VEgYlqzEbLBty
owDMnX+5u931qLplEYM53zopCYw0L/jUoYui6HLsyrNVI3IQCU7gkzVlPBjLab0J
s6fTiHqvFNwcSdQqLeolO73/Ak1PNZ1cE+YXeIvb880ETKMsFl0hR+S4IvYj6vxa
z4ONL7tkBiOwlFoQw6jogWnAURJCKOpi9XhZ1g6Ajw+li3lCVt9F4dldDrIhs0hQ
nHHRl0schTnZruJz//j7R0gAaGzHJIT6M/vbNPofWT/Ki93F8W1gCM76YOJXQiVk
ghv1EkYD05VS5WP5mcOvNzI2F9+Q5nrgvIPAKGer8YPVhHvOGs9kZ/nR/GjwOlBR
YzetIpjA4Tv/po0q0iZrWYz/wao71UXhVwiqF+OBIUu2W78y+9zUT8sWdB8LmE1w
0NiEzCosbCZklOGOhwv1OlY0DpvadIkWxenGa8fIAp3NmSUuVAQo802vnyj9GKHz
/cp4FrqnaB4StAIgApHYbOeaxzGdszqdkB6HCxy8X6UB4ftbg2skNKH7DTYEuYSk
7EAa5M5geLRXWrc8sLkwz7HsMlD9ql3IqIVFSEBsKMy2kPDwLC+b/GD47R4n/0wX
g2zXdqtsrmlyPslsQlAz3f5Pz6JKqmVvJ6fe5v5J3TqKVJV3wUxBs2q33NLJ8Mkn
ay9NxeCs9T4kldIQAtU4DP7wZOZKqOLNpf0WfKqZj1Nd/XJT1uFEKg7v3ruMsl6Y
hWcDCd2XtVBEnIgxXhyBOAbRPHfvb2gfDnWE2gfRevm6txNnxbbR/1HON3XN5yMn
Q2+ANuXl724wW4tet1TeDuq7fOAbW5mwRgPmUWjuGOV052SFceSpQbpx4gmd5oIb
Ad/tPxadJG3E6kppKOPi7NRRQUidLGELex/t4Yqkv+Lq92IccTlyMCY8Pa4nvqBW
nrzxuQuitLpybDXncChvVd1lr1FWoWQBC1KlDDMEtRVKc7weWhccjB7/fcSIY1L4
3+hc0KMTq19SQ81nIEBW6GAXSdzrFmMsllWbi7odfKCjSB6YvEboYrfhf6P9ySri
KlSIuGIl18EJWNNkupooo5dAsZsLrgQoiFJprmohUkwb60mi7IfgtgOxA3WJQjIi
OktQEwFcujRnHstGQTYvQ7ERDcQT3yDRLPfczRQ9F0FOT8I2v7tmfpWCFuY0fhcC
ajThv9oju0ijLfpqJOsz/d0GzAFKiOIP3uEBheDBtCsJsMtm11nCE/pOe/r1FnDN
SPc8jaz5INYegITbnWOQ2uXDfFkSYREMFDtj+YskQrUHJWFgOnTFvQuUrsCLy4bJ
sqUPmbs4bOwijgynoW8B8at4cwFUMCdNiYDJLINDuhol/IAa9Hj4MhcLmFaUVesM
8peOab6BZCy7uJ3JLbQQDPnEg84XhCyTk/E7MVH7qPNZP2OLQRMzTK8HvsR6Vp0F
oJZKRwjDTVbXCmXV/fs0Cd/hArQ7QoHQKw2QuxhuONY8O4UFaKd6MAJpQE5iq1+Q
jYFd6/56cNKCcCPkj7VGlWfytmlK8UYiPN0uMoKm5v+mV+6tDRSI0iywOxOuxm4k
/xyWW2kLCQ1XEWfQlWQs/nI7+3VQCRzoGbEvRrx4PhI5VQXd7RWRsyOhhewzgscX
/i1rYn0OAku6RrTbeB3+nUQ6Wynmr23uAI8BpKffszB852Q0xYbxDnI4mooXm+vK
D/D6zBtrXikf/xKRCmv+naxj1xWHTCCe4JsvpRWPyKUgdNAP+Wsx62AvQeptoGyN
u9FEjlC3O33ft2qICUUWSpo+20DOogArSLaz9vl0zNd+jVBG3YAqNuoRQMm/4GtS
NpwZ0BQwnmVRTjSvu8Pi27RxIRUnIvhhicW7l08UJH0lQNkqFLLMpQWI4mMo+KkW
gTbL2LpS0MW5+UXXzNOFW9w+F+m2bPzoTzejNjP5EuI9lmnObmpaY6CdposS3lpF
qgpMBqt0wAi7chZ2sQVFpsJK2YL3ajJmdIbpxDF09J1tbM4O4aYvfb2p1kXc3xsm
EDdlfpKtaMy5FCIKTCvPUXqcUYWW65wShWGnkyDd0xAvvfCYSeLtl4FrGMDz7gf6
6Lo6mcax4lxRVRDamR/WNfl3bgbJUuXFu5AK35Jaa4idSyWk7pgQT7RH1aYaLBIj
MZ7NHghnpaUqi6qqKsaXZHOH71v/g1vBzpP5JLPTFCgCBPzDmTHUPgv27fCJRpHy
F/YxFRjNgcFGwWqTlvmEts8o0irNeOA6i7ffWpLbM5UxiVgUWpZzsh35eEdoHhhX
yFsrO2Te1KjrM3za7qxO5SOq6loAcrFLoJeOwDNoE219xVVI1d5t1V9c5cNFldF4
8BvDtwq04VYdgL14E+aY3CZwZgJ1zYP1grlvBfJ4/qJDqJzzlKbu7mgOMh6ASO7x
geMQo3o1gR/9tSANofUO433YAXc9XXPUopNQEq/HubLhKi/tiN+1Z/kF0R4dMP3B
fPaiig8cnCjhdXRJm3GVwptj4JOtx806uN2X6xs7RUTkCMAVUmsux2yqYXJ9fHCr
9ctOVu/Ua/oUzyx06696ZyJvVyWegZGnb0YzHk4ntBE4N6Y/1/MDdCUuYCb811VX
2QqBQ5C4wuL/kswVP0JzUP87gZZPXv7VXYydV5RaUkaKKOF4hywMXfeFkz4WtFQJ
eWVWOD3630LaS3RGq8yaDNYs9eUO1bVqSFgh7KT2A4J09jWXBYsdFn4IT8Uerwrg
4eR7pxEZ8Qt4IJswTPerTEeomS1TPMTSYGoCE5OMurG8a48ubpDeKkZXRWAL8q9A
9Wd8sWf7PXhUvpOWmdbSSRXYt3llri38mMbOef9zFJKehRAi43BDiylLV4vTmYEh
8bUWP6ktjArUh44+9LoHvEALnbE+5e//ai8qPGVcpbe5KhJQGfs59NZ2qjaH+L99
cjW16SPV6kpgjlg882xfhpi0P/r0uA/OHDo5wm7lc0mWlAmS+OwGzLleBBeO84sU
lmHy/GD8E7usOE/VGx3GRUmaJeFxDyZHJNIL5gGGAwfErab1XnvnFMxSF78TrZZJ
KibZ5VvLchJKGE4tFiO3KeMB19AHbeQMnLYJQ3r159GklV3vlj5z52823Q8XZNkh
G61ainbFEANjNHaHUYOl2N4mzbx+Kd3Pu84L5THIyBF0dg0dj53jpQAcpl2wKBp+
nZ8wJY4g7adYtCAIsm6N0oa6ZR+juTq/1ZIRzbhXkVit4UvSqMcmqP6qcQodDjLC
HTRcf1HM4u+USxulcGgL/aftb6QPVlf2h+c8e16CGVNwIY0NRTnhzuIuVVH4GNyv
7N1kNa+WcHloeLpOO2taM86w1Cd/dFdfwjLiJ6VhHs7MEtZgtD7TQnrAEfgi12mz
YcszXyMtyuzAplW3OlF+qgQ0TKpbNUp5r1KJkrIlJ+WRtlcAjvCLqclok7JXxjhc
LJJCBXRvd6890pBcfhCwu6I8WWZRYneRpMvzOHWkx+6GbLSzvlBpnVN6R66kCKSf
JUSr2Rh1YbSXBax6AC3/OQHQuqwd5zV6KmXixW0zZOq5m5Db48S9W4xl1tPG4128
FvYgBXKmPcMxUWH35R1FjamnL8S4vl8qqNWAdYVOyrSjLJn+MAwiOnMr93x4m62u
qaaj33R+3Md8gsKTI1JnqY6I+TUnuf9nTFssomckxpVcPJZXBynPgt7RHyp/Cp25
tEV74iOc4i4yzRwHg67AdZbwwlgO9KS2laLipfvs1+VNMCTRkC3hVZ2ZuK/FgOAt
mzu3omvnYOokP8sTiQ4JawLRC1RWL9lk5CiyBADUTGIj5/cb6erdOuzqi6LzZHbc
gEtx0DptLzC3GuvqdYeam96vtT6ehImsUG8OoYu66nPFf9GyjQo6gCzALhXS5s7x
NXetvguWuH7SwGiq4hmXsvA8dSr6h5IUdjV0JbgpgWjtAScbCuOTLMVCoUELmG/4
ysx2jgyrz8XMrqHKsoyltA2S58R4PR2JttbMZh/rwO+wJ9jxtTWduHGSqAqT8tGf
/NQo1Vch1rfkXzvn7iZPJ3n98UaVoA2dwuQ6RcpVBAA/L9u44p3WgXkNUXxZelIZ
XZmnzWSSteYe9fMv28ofI1YAAnsql7DCttnTbFJlmYte91PiqCjSLbdSO74SQK8s
h/wLMJEk+kNBubLIGKbIhnMssIkS1J73fX92AuXIVJrOv/1vGpghnwgM0Fa1uqoZ
rYXTucch9S/KjYGssbCZwCjqbe/R7mtJoMFSMAnSwswVSTmhjk5YpyRMgZuygNkN
r8245SPsUXKf3dmfDn4AQK1wn/TUjhTW9Q2VKqVHdwv8SFdtR9/K6JHCGEe6xukE
FV3H5T0I9VvIZ86HASwQr1G2g7H2uDPE/tYHp486mwXi3sUiCWfvhioMVRm3PMZT
1PSG9WePoQ6ru6mv2KYLu5ORC2Ode1yC5gW2JHutCkqKR400zETgroN/mHyhz9xE
d2mMGiwMbUixtHTiNoqdd5A+VCfQ/mSpvf1tdsFX9Ri4Xy1WS2NWE4p6DipLIoWx
tWzGmUzAju7RatcwZ5d44iCI34hlNAw15A8r13EVRuJPXBBrnwezQn6VSfvtf1hL
wi/Ar8yUS8ZIVpviY9fLRv3rLac4OdwC78f6ihCY2qbyw+quawDj8z8XFwXxl+GR
8q9wAuJSDQ4ycIwAoMBE64LXuuDzoUH9hREuIuzh+yO4sUzIH810uaLF4un4o5fY
4pM6OXjS61q0S4reBT/XQ/3qxSvmmXkuTSmIkcDWSa9Zuk8XP0rd1pvGCWJLuwBK
LBtWG6tf3L/kgpYdOHj7U20OCmvLTM/bB08oVHutmzZdIRrXQbBILEvlMv2NQI+U
OB9e1YArhkbUNtAMXKwyeoUoXh1BWJqZDCq+cPqegfJG9+p+nyVdv3rJNlxtY148
F3DKCK+4tDikUxoSfIOIyCfrtc3TIVynmdHAKMg4HQhXeyLzyM9QbBy0OIRJLO2F
vC0Bz7TixddReqEvYYPmtd5qfTXaB3H7LgMMZukfMVuMZscDl9G2SdjIHSdroEh4
6MOMmZdzQ8L6O5grnDCZFLfO4Zv+40SIzHKtQ7zu2u/V6CoI5FiiqBnTDplVZ5bZ
ij47jD1UORJa8ANYRnblb4saAuJOuP6SmOvqKl/bCE2sABPf+D2eN8Vpb64Yaydq
l+VhD5NLt+T5DOwmqE4qafC6eGQAu0YGXw9LpK7y+CUJqSPv91mcb2l0/si76Po7
ABpD1rCQN+ppoPvDGCwqZpEqLCdQM3r2SJwkTNFMhMoGrluGLsKlhusHBhgTNZ+q
FNBnzudS7qG4w05Uf0qdyJxA9vyscXiXojxgu/LeDKyT8ump1Rj6JdCi5s6Jwi39
S0N4eJxJODRNYz0DyojLxWATCyFNxF9xDvR/LXIjZIpSxb78s4IDpvM0Bh6F9jdD
pywEkPrGyig92lHQCj4xUSJ+AWIWnZO1GXsZ1F6/wPpZZXAVapm33bxJdR55XqTO
vdZITcrWvBJQvl9cCCBlhqdkNEd0cKNm155uzS3L4CM7cCXgtkEQS+VFpz0bCE3P
wGt+V60IAoSuwBL3/40uSC/ONdTkYsfoorsC0waiFAWXR4Yvg2ztkW0iQ9s/XNPk
6TvemgvoCaTb4mbrOg7o+OpHnfFtjHLOWXUiDhqeezB+yaXzULMxShG8ADcO3WOf
7QHmg6NsSZUVHB3p4YS5WIXIA3WFWMayjD9WBmqNhTIRgZ0sIZTd/F+r5Fe9Ylxg
d4upiHPQBn71ZvIyRwR63q5OXlWdCTA9MTmwi24+fQ0njIlNVLjvgW5p83wVx/YC
owrlUT+x5JG+68sRhQXj4M6x540mPgGGxFiIOILpH5cishz+X2bz1rGxDCMm+Utx
gBtlO0SbiuOIKOqBdpIj6G0ScMlCc24fRZp+KwYVB/LikThTeJuH9Lfj3XK0y5oT
XQqyS+pHTcbnyCPgCfhAXhywoSIxVfUGxQOHOIOrS6btj+9CWE8tV+bWQ9e9ypi+
Uk10iJZbvzTn1CqPPb/ysmmD1ib7Ml3iUyCBW1sE8dpw3xAHoWQKfoLvPYfnMFF6
ihHsQfh2TIaM5nII/tU3r5qiVogMVAReqh7f6N9oEAgReB6dKt6Y6BUAducJiwR1
dA9l5SZvpoJ0BbaUF/KSTS2xSaw532aNsLWGZdmTnwgagXiI7C23XHia2Pn+4Tsk
OfHlB1XM5mYoQVYFwAMmWvDEwru2cJtxSycVHtSg9qKHysXvwoUqov8qKS9Fhm05
DvrpwQJ3sFV0ftMdyOPn0lUzRgQKzcCX3f/W1uxeRDKmnFdsvrdJ5AFUuXkjjp99
Uc2Y0ZQIxHZovVU8CHmJDe/OJUbbQ2Dfzw67/e4NyhzMryjseOgyW8t2jGRJ4ox7
7wpnYMfsygheitTTATimB+EI0gZ9dT2bU/Y5BDn4DF/RfviKT+KYW8Ov8dUHxD79
uN+4x/XHszFUP347fKwDkc4seSCJYvgSzOmaLklwVieCbfYqsHzsnkiopyqr+MvF
8Yr2jgfw7wxZxmSVF+nnymg1Zis8rWubbeFpRl9bPnoiFzTsZ2y0rrq7Vfs/ie2y
I0+V7ZA0lNk2WvtjMJh9pgKJzb14zxqGD1jdF/M6iN5bfkkCfhEY+IzFh75rECZE
U5MSBa1a5KfrfsZPiHrFVLvQ0jpagMJ5Ir5sRLF7hj8nINZIpc3QXm/+wcou1/zD
FR3zsXGniNOIyK4JAZmTHiSzZE0uTY4EUQQQkzIbeJ3pMoMxh1e37R7bv9AQ3f4l
wMGAEQopdYNUjVQqlCw6hdjQ9KiFavOEqbHiLq9ESxyaYeFDH+QxuvFXoM2yPk6B
pQcghbrQUeGbbpdQWgUwLazzdrplIebQJdlqUx4rznjqykXLj690NMr0vT1ytxlP
7Ok2bUTtW85C09EOJwyDR4welDkIdqXIOLTkCEj8hnYIFs65eaJzm1oYLQmNK2Dg
rBCZPFYVEYQT6pdF6ao29r9O4nRMgYildFWM3DHzg1Ca3Cwq/CHgPJR9E0vCAnLk
FDxUcgI3PWzDuW+cxNTpjbC/dMVoPHtwTuljCP7Ky+RFI4/GbakXOepTM8aCQpxB
YLTAICdhghjitCzbZuam8nAeLXaSUYRMxWupE/2cvjb3nLG4db8eXh2mUqxD1pJw
Z7eVofqa9zkdzzZxhqOQSDq8iY3gJKMdhGXfasgXsKWhtiXTbDWKo74Pmku3Lf3d
PS9ZKYC+45auyiIBAg6s8ZjFGnfkM2/1mwpOQTs4RgYWCdEeBvBh87IiomhWKIIa
O3hkViau/ON6sX7Z67DzJTtyDgvbnXtTUK+yeSXweEcm4nNj8dLw6LztG+yYsklE
RIwUMv4sr1VZ3AxPkJcv+cJ99G+qkyXyKHg0e+U4iV3AiBfhHxLzIqnRIFiE1wQk
34g9nhudr4KNVCCM8h5HL9iiTaZoklID3638dDm294/BbrXXBOZ6RjJNhj3dYogW
hxxfzTlvcEicJTTn7aPbFMLSxOa3EtGyv4vxPN+vQoJ7fpfr1QROBwbZbbB0TO/M
e0VXwvpTm00/J/sEaJlXNHcsLzAYbw14SQPgMtHXdF2urf8SisdNR2ccTTVmfPgB
WuUw9haMYv6ckyvQelYub3/FA0vqwd16G9MB2tCcEPfLfQc0TAcoriFLmEyskBB1
yW0T2ImjjJ6n/LuuWvzVCILcOq8OBcFL7RyGmhZoFPSxilp2pmG+jb60IgIV8LrG
y+2AdZrMaKbk0isrIMpwHiGPWF36VUqvIxnMJ3M6O4GxM2VQ4w+DKg4ppFgbyUzh
aCVHAKvWDD7v6jByscfhm1p4Yz+Y6CZA/ZiBTwrFEZbP7ueNUO4mvq+w7bG8nyK4
O50HeuSKp0Ppib3Q3q7JDoMLEd0R+nKYIC2C3rQOUEDkCtE4+vl+DRHyt1iHdOzo
sw4TA0szh+Km7y1l8ER0FmtbGn1DcYE4fCSKe55NsoY6Sju4l7jLfQQKWJnr2Leg
8J9P9xxPBM2wGLv3YM09TLSIkm+HGUOUvu54RM3oVUsD0ZMgIkakbA1iH1g9BRhr
FOMVl2ddZg+n+3KPN4WUQAvlXDTAeJLsad0Nn0jkTWHtj+sCe7fd+ergincnGYTr
KZbSIfwJhuyBixs6v61tIKHfhkF5hzKYagtTGaVsXegZzVVCNitemdOr3rNMlc1d
rUqkNn6KQgyb3zNVzF1xawTzynlbXy+1XQTPmojcYu3pTR6psV2WkfRB5A6vj27s
LeiP8UAf5M3Yt5UVrD7KsKbRuDiyxlhrY0usrP/cBHvpdJRCEkSR+YqTyhvffdlZ
EtimxlTtrI7ITfmdBMdZ8yLK2e1ip517IdU7Pkmeg7E/7UX65mj8lIiCHDc9D+kS
rYpAJCD3eQWXgdd3hQEUybDdcdtUJxC1sXbAf81EMkI6PRWvj/g6WuJswzfEvEn7
i+4jSbnGsF1GELGArdt7DPSBeWXSfv8aNow2YCgvf/IEaGkxztQ0jfnlzvMmLhed
rFZSWy5wzJHw/I8r3X+wpKkjbdvJ1U1LTZ1PpAIxe8AS63nZMp3OY9wMOXBaxkat
EUEMCHSQw4eHj80VAFqsy2VZoqqjNJKr3FV79kO2SFf0MUXFS4pceGuMw+vHJcx/
J+KbC8rmmCKy4AKk83VL8mMCzA6zWuZ6fBOzlXGC9Lt7eRa4zC3oibjdVipiBN2Z
yLZq4Q/vU88eMZknAC2xDS1tLVLxqSctSLHwI9FFgasRkA10yfwrfFGa7YRpml2Y
t+sYWH74v0ssk+e3Dip3CnFpXpfPG+HDIUW3Xg/z/XBpZHRTryJEGeOj7UXPg0QD
CLdTYcFQvmMO4dSyyl3S7jOwvg1frddhv0ifcxNfF+wV2dL66nmTLIVuEq9Fy2xN
7i1AAGeHWxA1OLvFPKAYYw9iXD+UjjaW0P3hdI/O4X9cEGStrwfJBgYPiFS5NQqm
q64zw2a07xXR8tRos16cqa9nyDYRsWCebKN1AFhmVcd6WtlCGjcEmxA5ZM+PLMmP
uUsL1r6UsFXbpSOvQ0+d9+h6bWIe1cPkZ7cCVXqJBZR5cw07GPudCXKDkPFk9D+u
q9gNZ3cOJg06u4g4UBLt3NDETy/3rWZ7L4sQPMbmP9CCQDBf63IN0J3wrvRacQrp
XOavkTpeCLykgLrrI9GaqshifaBIONAcZYBAl5buXuNb/kdt+U3uvJ9+/vMKGT4M
rj6TjCB09VTw1rrlwabJ+r7S9s1G63ReK+orfOvA39JNJTzvFFB5yYkO3YeAZiO4
TJD/Hd5QB04cq3tSqbx1zLSILf1boUzLC4W/lu9bAO7WSCow6JuuApLyHUbFJ0Hp
ZHAgkU1n3VWdtGEkEDEMguLbt2QUC/984FasP/8kWsE/NwlLaLpRRcdAqx5wlQ2+
MGCkKfX9E4ADkA4WpsYSMa7gAELAPQcQmbVzWxsutrDPIZKPVkPflsF8Z85cmSll
KLZzlY8mpozxhihkEOKUOSa6GsPYYu4SQk9qgfQuakB2fbg9dvOcfosS0K1nH+0V
X0S/Dzr4EtcG+socC6IfNml9k79y+lGgNb999cuxrJFoagvhHH6OznTxWVlsjfPu
Fj7+z1nzaJuZBKlGURmpB/RbSL9pOiIXzz2YsQ9wH0LQezIKHHkRJjNaimEaC3vC
ZC5zvdYNhRIiB9MiyPCgyLdvHLpxJW79+jStBxl7Rw54rK9VIY924j1yKANcUEOG
8KQb4ES7/fOSQZHWYhvRI6tXLDMEGPFLeMsCtTAfSEBQiII21XV8DdL3mkWUSRMG
MlvUpmT1MTG7BhQioazc134p6ZEyN/1Cb9NP3BaJ3Ilt5OFvrhjGBpscDll6JNC5
OKNo89qmeSGOhexeLfMpUC5a1HcuUTJqdG0tK1fon8pjg/nsYvQkfYDa/OGIwBf0
G66KL9uRuYznsoYbTHgnqfVUNKOW0oSEc6VR6vm2Aaz+pDpwBtQ4lGthUf9AoZS5
ebJO7F39sXqMyy1l3vtXybQpz2DQV2FpectCL5BGJx0hPLwiAC9cAnXbbYzJhvA0
3WL32oNPw3GUmWjPR9Vyhl8HPo7esDqVSGTolQcVso+jTeiB0vdF4Vp2PITszkLH
ZagdMH0NI1XV4lOdV3WVeJixIBK1LxNiDjt7Q7Dg3/JslTAT0Ej5NHU943QjevL7
fUQPYYRWrRqXw8LH7fS0EC4EI7XzYzA1KeTWpunpXcFvazL89CwnwTbRzEqTAJi0
kPAk2qM+yE577JY3SMX4N2JJMEoj16zKQxt48VPdQzK66sgnDe99ijLGGRd1NZAy
BU50vaeCp3kPJGTWDYTx2Hwtht5FswHzXgxOaAazi2/xPWRme7lJBJhlbSm0vFQe
BxOc60a0KBSHI8ipRn/9eR6RvIMXruV0wgKZp9+2jKsJDeMiNgiDKQ3zhmP1UAWF
PMnYK0emFYNA5jvd1NxZPeR9gxIlcxCg5petKElNgDTxrJpYLCTyABiOI0Ited64
/0OHMrYg8CNh3Hvyfd1NKSNPuM0xuuVq5o48RjgTHIObeJV3nu63f5PJUyDJyijO
DsMqkX/H2/0ZBGlEapXENj9Ia63n+lhZfQrW6OchmrzYifguPZn33FH48rt2V3LO
8DooE306LvUmX3AsoAQX/87/SH3BEem5lIpun7tes4bClL7vmD8tj2I4OE4k7UL9
nKI/Pct8SHBQjfZdibhmxLbfDRt2OdEw04v1kqc3yd1j4cuiaQ3yHnEYHNxMwHpC
BhkNo0XgytKOsm2UNc4rsvFhrUYLT/YSfV0Gv2HBxtBwWNj1EolYupCuAO7EbdL4
3Lrm5/QAPH95HigJxnf1/LjflgkmzfL5+mWtaK/BjPl4kz1aUThRgZ3t9DRszDKP
+CrPcSBDq68T5Et79k5oicItEMsh6YHKrIXSz/94iYBHUuGbw+8SbkyGhAA+joO4
CX1d0W+TCQjRy0f7tomIx6afi2QOfsVJMkQYfe1XbTs0tQYnKyg+sepGpmbGgbVI
kutg4nXEok0qWFTb0WHiPd/XE7RAPBS+xyBYt+JdYZBEh9RQVHjg4ypV5S4ipbCu
LyLW1WZW/8g+03MstLEQg8sfL+vb9RSJuNV2qMoK3pO+KIXY1UOH5B8IFqdkSuTQ
oIM0H1vVjf1NhJyopIfzMUUJUT0gnZw1xEbXGa9XcbI40w4OMq65Qvap5IzjvEiC
1KGAFwPEuWGjDaXZT2H4STm8tndweLP+k44g/op2l5uOqII8tSO+q6IXAZYw5BJV
aygX5LHzTymRveMyS0/5S3CCaz/T4dPyoU+9cADh2kfoWr5W3Xqfpilz75xnc7v6
oIywNF23lLyIZobgl27H+cgyp9yZLEgPHTd2Y0TEXHSCUTuEPyed4yjqH8Wif33S
s/AVwtntn5LbjbM+7oTH2/pA0LriKBJNUAa/7W7Te2EQr2xqVu7CK+BptmwQx4d1
uyWV2ozA7jO9nrkG+W5eJNFTX9EnOaZfmkVXggqxgvcA5CwOJ2bSDxfvJ7WQZr4X
YU8klqdWdK1bGQcGEB3+2/IkOcleA4bDwmJRc51wvALhmXjSRIQCfwmFGD0v5EK/
w2wnBW054TEsS8Z15YQUFN6IVS3JKHKzD3IZFXMEcVinhiDR/JyGdD+9nTlwtkRk
DNf+c8CzlgJJ6tfnKXz0r4tqF05UJj6pMCI+qxSYTOUl+K4nH6pmd9yWhc8UuSH2
boFpdAEKacpYTEMMWF/pv4WPs2cfvI2ahdUQ/BFMC9tFBErUoGA6tnCUZJL3dfwL
7KpeWCCh7LYcehizP3WiL52ENjD4YUGwU3ZhOpkBVuWexlNVIhP2T61NhgIrH5oU
Zr3WA75HhQpL9QEaB9Yp1kLrSTPICaongjhvgDUnXLg4FB5iqxS8eSfeDQM+W0CM
Q1NPGFYx2++TxFd4dKeA6KZctKqwVXrQ40iNcSWJ0RACALFLLCXLBPZeT5FyDjzu
FLc0sBtIg/B3qteyJjsve/qbu00SbP7Uxl6+Sc8tNQCD6Tnd/06bQRun232jzUj2
7VlBHv8Kq7RG5Vx2nhcEMPwnY8WHTaz+ZNXvnyBq4YYTir1UNyRERjWXQOTVn2E0
lC/Dow5/+7coYs2Wfn2Xp+kojGyusfGaozaLrv2j5JtObbF2tGLcgsIWxyA6pJIy
LE/bwXGWftQ/fxtjKVY7ULf8dnVNgiHg20m750xS2UNWn/XK/zy0S30p5nINO045
H/B+FHvtJmR4gDHnG0UMG2hZ3dbHk2UUFlSWM6Y05dNEHz+YKVwrU1L5xOC7p5LT
KxzsDtF+ZTrpklQbl7zLVfgwuphgXShFCMoS2NeoH4A8TedoYv6RfGQU3t9ua33U
vrxGe/6A5tU2HE5DHVrwNRdb8fx9GCRuiJJYQZbAqOdCyX4slN9rYoSvRjB9rDKU
PPGOkWWLVVhLcPhkA6LhAmcNabl6JueJUb1ltYBWbZwua3W4OsejKguXUjXmwKGS
gH/HEFI2rPda7oVNhIO/btO5Q+tRwNKqwY1cuHHXNsrJreBEjpAB3gMZIMO3DP5y
Beq5g/VaHaywYrghK8NtML1RxjAuCXI3O1UZZpSKung/XimK8znwaBSR5JbxL6qn
c6HG7OcSPp8frUDgoUwMp6P+EY4ERgn79Y9r+M3Gacma8YTadpdeqDGS0Evxcj48
YyJ1s/I8VzfuKaMYcU9xc07txtnSZ6ShjkfuzUH05+p2bLTx+fRaWTqSc/RZvIZw
HRHJfsqjOk9FeTmj0xQhJf2l0G5xtVQBjf8YR/iMx7L2MfxZLHRMjjOlk+tFwPOL
O64A2RsxYII3slN0IAU54A9haljNuHUwMLCazWmHIrraAeqjY7nuaij55nXQhr8T
msJECXcHFjJKZySymvGbp/82j888Ql6MGHMpcPaW0YhKZbzr4/A/GyPILo3l2yfk
3XhLPbu+jA/3Dcd8ea5h+7Dko0n+cBl9uQQS6BbOY++Xsl3Cqk1TM7g32T4XsS7w
Gs6O1SjRWCVX84Sm0iFFlwlBGlXiWKQkx6cXR/v51Pr2VnLLZMWJSYOzx4zTXG9h
P1JgQtki3vu0N6WGYoi9PmegnQhcVBJhRVwerQcYUc1bJ9O7Tvv2cjUWL1IGnkf3
y3Pw9kFYfwj8eRBvqj4DV9xDLaX0YtP7VuA7TLTmFry8akcrKvNXBxwxtMmBw0Hb
HisBltVA+s9uEJ2zbfWlz5bTghIxVGE85+IicUqqASfLAqwnyCIbNGjm5WhTgY2L
A7C+9bTkiVQhaJxGfYD0vlYL1/VlayQwjq0Dvy6136SYWCI7CDp99HehyzQG+dwE
jCOKEI3wXCxLsB2KKQC/GBVnELaqDRUH6wZenOAJajuPHTjAoMuL2LvEfXnYfZHb
dG3XOmazkfPyK5rZNUIXuY/QfUuLa0yu75nKaV5Yqzm46gUwCuiDOwk9R2eP8k9Z
I8yQwNS3or9mSmuROaJquuJ6/YUQejX3nCOTHhlpt7V9f3rz3TwHK1pyRWzAgrqZ
lBeqm4fCAT5eZ4NpknSJ8V8aUTCxHaaa5q3Jsv0g5QE2/NgZwZQXftxIPppJdpM8
WV7gHF1sHt8DgGmt6BUoVvRDBWN2r0dc/p4hBNz+SdnBeHlCUf6OHlDkuyd5oiIt
Ylkvkt6/rsWaRk21bilRB0lXRoVaRVHNyXDywx547LrOpXzAE7qT8xMluz8ESZsh
ikl5a1U949Wh7QzqWqyTImRvX5xDiC9/FZgUAvUDfS9cnivfabFeTZpwdleiBU2m
oyj4nSWFq0crtKHKQRgTU2qX9DZXa89N1aRmXpJeGy8/Sn4h9P9SRpo/kAOt/042
VTeEFtfbGBMPfEc4guyoIKqniPFn+XS57asWFXRZidKADrQQ1pQWBZ3VTm+s4atm
2cnMWPIKeXPr+rN2IRro/6ic5N6AuUduhOu8Ftyz6hWQjfdIr9DXwh7pDY7gE9HR
Iq0zRLzVjHTappfQRmzUqKPizW1ggB8Ng9WyuX7rKIVjKCOD35vRNfmph4B82uGe
hMwv3sRgDOtdgKe+M1l9/w9zNFF6LrqzDup8M6azuJINAe1D31s8z78ngqOP+kOG
BMy8zlMik+lCE38F5pATb5Hdo6CttUp+grZnqqYmcYC5DMYtqS0h0qmbtvcZ3SHd
LRQa7py7+MxK7T8Ygm3b79v1p8bQMN3Ac0t+yBWxWk8k/yOlFI/voPuPt0goozfh
8t/E8CaHUK2P8uKfghLzqLEISxV5NQgrjU8TBZFN0IX3yACCwk8aKS1hpkqHVyzA
oA3cdWnwc/krObLxPpTWhLtpHDa77HoSLE689/qU4b2olXuxLFiLpyBaQNy9P8ie
GbKVAxiXxuuqX44FnDGMYgvdBO8DEf5VYjvqA6uMhmg+u0sMJR6W0U/CmMU3XMUM
rUWQTx7POMbQEUUV95SbIBNO01thqrqMs7/p1eGj6qWe0rDgMExLi1zcaH1qNUBy
MBRB06R38f7f5U/FBPyd/9Dl1Li4Py7GPfvRZs9vM9ubz7YSm5frxGq2bAN+7IBg
mx2G0cBbqgu8cJpkb6Qeomxwe+xi8LCv9Kd5rO+BrAl8QRkDNLovuGzPHjduazLk
3z1NxZtRsf0G3AcbFxwN4l6EDeLGit5RiITjnoDE9CHulF05LOt+h74QeE16kgIo
IZhe9NHie1yL6/yvZAuISQwWzsyOvwHoJ9LjGrYHHQZrkN8ksR1KlyT1u6dz1P0i
bmEu87ynp5z1lDjumuY56pjYKKcnwRq3hiJvAkNlnoLgk9iPUOjD0AkKOxk4Fxp8
IBiUwV9hAaQgDlAklGwhIk6wI+CvNlVVavdpzu3CwjVaLpRYAjJ6OrcQRcgErvRm
V85WnGL9DWCQaBw5qAS/uspVhHdEU80PRma6piPmNpLLeQaL67mIaGFC4HOey7BI
wtR/+a8/CcPZl9TEPFBBeeLLnn066jtucQ8fVsgHqrb7s0KbkRp/7k2lVbW+MqrV
uLPVxhp+zJ4IbxWAApQU172gUYx7p0miWP+irsde/3p7fAL7+ab97uKDkETRYODd
lOTkzJAEV4YdGoym0ZTI78bnBYoBEhK1+Tk3hvXweW/Q2NEVk3gyrGupxQhU2Cn6
7wIuLnJ3gNGL9Qh3IS1x/a2MM+gbUvZpC9Qd17uZSK7GNagjE+/piWDjkLZZIQj4
oS88DM2OVOt5DTRjBjelp9kSWWcyge1mu7A+pbsbVbiH48Rw/VMHjg//kUfYjMhf
JpzSqjvudC4NY9az9Si2SlSGBQzywVchedwRpRaPFWPKa72/Dxqw1q8Hyx/4L2Cj
05Twh+zeELsTfhpXrgq+fZvYEB7gycoGOBM46dxdov1sYxypRYug0/0aB5Uk8EAK
nSJl+5dUu8NZlAqt/4zFEuCk7KScWrVnF5KLprentj/kpkbNn633NDf8iqmd+w0A
oAV2KrlKWGC4HAcZJ5veC0+Qq0KjfE5GWtMRkAZrd6qEBl9Onp3DHFNYVpNGpyrr
mbX/pD1kv9tiO3ONkXjV/hlR6EmsD6BtF0ypxH/UTxj83mwkLPEtV93OjFxpWTwp
8kn8zlLMxVqY4gsQshYSXW/LOfCaU0WRFj/D73/dONlHXA97cXw6azUiOX76x0RS
cW+Q0zverRyhe3Ue5os1on7lDw/wIAuXY8l4R/RV8PWoUMrEV+Ch/gZQ0/l9LjUJ
2i6WO6EDrLIX/Hg9bzS95Vz6p6OO9SO8Jkq0NBZd7Ei6ylQOLZhMuq8f7G22NbO+
P5rTKoZxtAmDslB2aYEiroWx3hfzTD+4vcgvDJ8Z/Cta/NtOiaXJc06EdH1KP8PF
DivKCvtNEIRncjmTnzYBeO8rzZLXLFKCJZzn1W4pK/GEhelXnlw9aQ9n9rJxcmIN
jR42ThP30bJ2pRTDBR7NzKNTMhTsqIew5+h3qHxbsAUol2Lxl124dy5XkY5JyaWN
SSj5MdKhH1rZOfEXb8MyFquUENiGx/yhkKowPmwF7SZ4DmSAs+RpDBU6R9cXofJE
Rvz6Hd7pQEj2bclWTX8+N4TCX/4v1c6LMX6jGzys8AfccjrQ/yycttT3HU6e5Yxh
fC9vn7EC3QC18pK4FUJMvy2v0vpOukXNzTYBl5nGesJ/x9k+IoxLYq3YDImw5zlS
jYnVDnkxDdB+DZnoIrBQ/ILpv5Sx5swRr3CEYtZPXaqQd0kepGDLJukS7PAY4m5V
iM3TZD/LhPt+MvHEbbztOLiyJ9OD+7yuuOlA0B/0u5U+mtjFo71vuKgYbHEegUlX
oxF97T/mwsfMaHrJxe4WF+3BRnMmZ3cO0Hi3VKZMj/doj42tXLXIos6xNuXPlv1j
KCAvAa2E29527kHU76W0lAz/JHlR1qoVCAoqXqbf8PE4QgNLbJNgnprLh249qLvC
RngUS65Kj5FojjmlMWS0ZKC6tp2/M8BhGAZnIbQfjKoS1kSRc7SJqlknfkXCBXIj
qP+EnWpoQZXuibzofuPrIesgdVrhUI4BohRaT2guj1fzjYARpNK6ljlcfhbfH1sW
TAKwYQCxbRDQfhZn2VAJrl25KBQqQ7tqolijWsDySz/lnU98HLz0XknHnVzrcX4Z
zIi/HEYO9bnfLX7+MpebTfywuPx7hlc1Gb8klxB/KhM/HiqjLQWkU+0sT2PzJ7DB
iGeEzrbwD3M024jQD+wFFIFjSl6MyYcGFRZPtP8dWZaGyIj+vvnWacJpNjynzRXV
MlTagGr4afSdra2X6dWbnaIr3QctiGYU4jB3i1b+al1k+g3ak9HT+UNKZ+0B1Dck
rBrWXVDH1c36Le8meEVsClZUGTKEqmUjtjzBcn/z/94y6OGF+V2ou9m/OVsk0F7G
HZ0cuQq7lSJ1i6PgXntw+82x+glevsvXTz0ApsrFdTuQjbtDUUT0A3X+esfd3t1J
9cdLftmhYiaTOxVRB9rX0dT+I+bUa/vPg52NHCzU0VZ4qWNHQxniAspAe28/37ai
fYMj/5MiP5pqHYTF55g/M6s2hUCVit44BPhObTdlQMW+xIRF2eV16Hm36KyiwDnA
97fasStzTEeW9w/gQ3uq6yIvzm7zGnGErRDGBjvHzj5YTXdvXi1JZE1j/2bqLQun
zDMl04iJymUUTLMpv9LlktAaG+m/IheHa+wHctompLbQ1apOFesjZmHe+jBPGUNH
baskJBiFAmpKpRyTEhW7I4y4vXImv+gsW6d+h0Fi6JQukazXxVbpDDEbjAKYuV4r
w/wNdbeUxOQHBm7EZ8rumLCBbBZYsY0RgDJI5v8PaGjODZqa1AiPrUO3YkRn3qVJ
00XxoTszoZ/Vor6+ZknikcjGJgo8gsq9dO6Uu6D1R9hnUjToonyvm/zyEc4Mo/QT
vnDw7Y40Zf1cxoa1FsUuHkCc428mGeb6npHwqpRPwTKtcE+yYL0n0WNvzOMiBUW0
zToFFBqOm8gvM3Moe9jb0saT0F9nEzx/R3BxvjG8zZaQYfGJ2RTmwHnSxobat1YF
/a+No4clR+t+sEcvLr/YYGzU4dcq1ZpfHk6IlYPXqusHyohFQknAOl8NTBAC+iHg
zJykh+LaxkF/Urbye6Xl31e5S2xUmnikc8kc1x7qloLm0fpDnuwUJxGrD+r5cNTy
0/JtP8Ah8+v5q7Uy7D0XdK6VenaRP3yQKz09crnzXaAO7Q/lMwUzmdk2kRGuvzTS
xwaTnTn6/N+KjUWD6nZDiYprzdqmKDJh3C8A8SlCA5uEzfmt5huAO01PYSFyr3Od
I2R6V+6SxG6j5XrD7HhdXLLyxbP7g4qaSAFifhUcv8bssG5kf3/F9LkLhJ7upyfG
vjW1f3AlClo8XOhhX3RiflybsJMcHQKkABGyAOF2Wmr9CdXi/JkZC93XoBRCX0/S
44sfs9djxEwxCxvIkEokFm/4tiSslKSk6bWAV+MqthbDkMwpHIH1OKYFz7Fszxtf
AAA1q3MUa7rKeFdoR3h6ZkpwqVvmgyg5rJMhVO0Oh6HC/bGTufCbmRUzTkG0SkjI
Afe6LdCByzy15ktDDS0jD5yrgj5XtpgT9O5MYJjicO2HtoWny68CmcBY4xIqdrm+
PlGHeDXBVTZ0P/Tm764IuvK4R/ozDI9VommhnDqSkSFclgr7Ln5pvtNaTAwjdX9D
0WHPokTdJQ5qeCnvQtbrNgPnLkh7JgGSZ+BzunBCWyolw+W5WEoMDruqMqQQHHDy
hBqlK3V97rm10OA1r7NfOhMgkRIU465qPehY0K9X4np/ACngy4x/ucK8A7mYcrk7
qNGh78A5n29XGrakWoe08EETt13Q6bJlr8fKnmi4fNsfk0CZ35RU7JhtsiWDw8ZP
caVJP3rzrYnsfXEy0PAELsVwb90hoqqIZ0NB44O80KtSMUST1G9NAXScbKP727ma
THBrZu65T3gSVKVluBKagDUCdyYGpee/9K3WyJkzQoEvEKVPa6XF9MDh0ScGWs3L
LMF2O5mwIbYVurbSlzt1S/GBcMu0f2+af68JFWW4ypNbhq990k4DY3NOVnxZBrm0
IbLIMpb9yKs2g0s5ZtWfISjrSn3PdKN448/xoR0XAD5+zg0BqiQLUSwfEvsPQHqj
Wt4OgDfRmVPLRu7AavYZTYdYlvjv4QFaQ83DKvpZur2D6TMfxjiKaHxzymFCNgjC
DEwRI46jVJNEywNt4Qfm6jrwNsuqhVpectnkX4h7tJdnzo99y8p6c2ziKeBM2O2Q
pberZUyx/rYQqBlxcYrEfxSAvdQHQB4XoanwsR7rN16/snm1PmFgGRzkwOx/0Iax
3c9Belc4VlBahSru4wZdz9WtHcEaZvA1VE1JX4e8g5KSTl6Wxh77fTCctlu/1I22
9+g8qDmaa4iM+EFgbBPsc0S0rLgvyPJNTaCgL2vZRKC4aTAM7+7RDtyysh6qWc5v
C/OtjAlZtoTQ7fLV79+lhkBFBBm57X1c/I/EJmgHAK+PpUi2LmAVsrJb5k5TyoBa
5oHBljbWQjiSbSpZeWGcNvAuNcmXazH7dPbwpPfS4JANh4dj23l4zowV2jXACu2g
VBA948WhiAbhBalYZmkkjYcb/UBxOLPd6oOX5AK886Rzof97R4dXLY5LtCFaoBYI
9IFYBI1lyt+JKI6S/lNzV1jw5fJq6wBrKjSz7353L9qSkFyQHTyQEOGeU+q0K18f
Y/4qHTOW54HFhZ2TNjvkCyjb0WftqNfnWull96TfQCEtuZcGktHs2F3r41eI4mmC
zl7TdpzwGNUWXyuldupLgGkdh5dAD/pVa9x8yPe80ftezfewR6fkSV864AV+tz5j
hQGMka8L8WuT9ebUgafDrJgn/007ytdDPJ8AFJ6UZqRNYWw9mfaEn89yC7H/bFAX
rzlkIGuMGlgp/NkXXloi5jquX+r23w+XGGgsdKz8ir7Qai8DOZFbtm3Fa/Ezl5yZ
J2jHDl1VN9T/geEDQx3B6gQHh8VYdgkfeYjffP6A4zkeyUuAhk/hxRjnqcY5S7Ve
E552Fv8sC0v3SJvGzCjhoj111XQRZeGzZm9+MvZatvAmDV/2b0vB46gcnCLBmIKy
XcnMnwTKhAgExvqAuvOAzPTHmhayAjyU9KC44mNwkuQ34BLGE2+OsoTjUkhOp+Lv
G6R4W5Za4XsnacG+309GMue2fPbHwx47WPCvtTWJeTPtQBshSi4myysh1Iv+Oa4l
cuPZHTP2Ouc5J46ZvOWx8plF0QZcEnEeJqEXQj2sJYRSjQ2VbZGJl10mqngu7XBG
l2Snd0lc00fpSOptfTAQo+IO0O0XljhAXrJa60UF5zycjG3Aov1JwMRv559voHEO
YZNCTzJYw29ZUiF+yOcfzkxIy3njYWICSj6v5OCudVvzbynsU65irIGXk+LEiRT3
TFhoqA6LZxwskJubMDu9uvo3P2BTP1jYg/rLTXfL0OqHnuypTV0iMZc1hJLiBUnD
ZUHNeMLd3VuF6DIkMQpnnSvABNFEypQhDf7071fyn/4Aeth+Gw1AzPofiRZZcrg+
8Pew4YmEEzeglyGi/3DgqiTVBVemaJH4SqoBuZwayHaunomKAhsbp/LjEcyapvYe
8mkj6+Ya0b1ae040KMCVabDlSmkgKf5DHLriBeCFOd/Ckw6xwl3qfpyN8v8cl1Y0
kEb1A92hTOUMOgbTqd7G9dZAkPrVsIbiWqH/+JUXmtd6YIxxkQIxernozfbsMSbR
YVY3xzcI5pcCexAnsCOeWyFJDhHM+3k20cKxCfy/YILHEH+kybtZKAklUSa14X5a
FGY1/L8SQZrpCwORbtnuI2WIrZzcoUcy7EoM6Z7V/IoDvoPnxin1W4bJLmPRSwqe
I/Ljo8FMsWWTrMpAOwzuzpmG4LdNMro6AYmWM6pf190NhwOjQCmoG8hTAoiCwWxa
c40KP0zwOLYfQhEcViAUsC10+8B2W7fMw9Sz09Er1OveMvYhqcAmkl1uSUFS8u8H
rAoWd8AF4E2gYXGzVen95GZn06Oo/gs5cmf/dsjL6k8QXVkU3dYjMo5oaV3jhNyI
rm350Yoizd36ElkOkxND17a3fjzzmhkLN1e/lOoiMKHkEBZthq2Iz8iu4hAe3JWi
Xp2L59yRJfeNGfrSi126XbcA7qnG7wCScihUU7rPJc1hX/p93j8KaTVpt4wjS9Io
BqSJc4znyaZxg/5XjMOXm1HOLmlzjwTVkFjBZEDwpw2OfL4mf3LIHyPK14zIl9XW
Dgj5PTinX6m7e4K7yro6mpv0SuZMo5a1ubzyXhS1eXgDHcevaKAJeBhz3KkJmC0q
i7d+Wbmrzy1GMTN374ch9qeKbq3VJQgi99X6Oct1nfKK+G1r67WVi+JasaAOCt5r
BvRGy2u7s4G8368WHvnOyjBLBkoTGUvmIbb4b3cYJi++Rkga1KP565KK+zfh9qL5
M+Ujh42z0tol0ZEGFOPlzrolRMGDZNhWQxghWPfPhc8DIgn8g5aPhWow59ki8y8L
LSBcIrwNm9jbxwLmKHCbnDs0bUXJIlNOOxAosQ9ZEnUewgRXsNeAbq5jZa1EVpbL
qGJ2nTKb7MLm/o9pmcc1ykOWjZtjgt4332LSUbYYb7HcicrGal8lup028D2nZyua
7/C7uhFdbFWg4b+DPDyvrarMHeEnRaiaEkTZ6Of9E3uW6412o6UXZ3T7k5AykZ7s
3z0H1snqet7jCdt5IZAMtBOBhb0sodbi1soruG2+VaUSquH+Cpr7Pmng9Ws85HZg
bgaUeWHBez0r75G0NtfRtet0Lv3IW6AKkv9GrOYHbg5HYTfdumQSe2eyj8p2vKJs
BgPbRA0ABsGkC9/SMlvkBTrHht0VzDoN7vA4uk7o6R6jf/n2zEceRoGOhNbzugnD
llnLB+mm4g7pvCTJVedd9A5ZYaqEUj1nTKRWYmHlQiNYmYgzY8Yz/Ab1YFSO7Hic
KxnBRPKQU32e+yuHfN6I0oyPAk04RStGu4h3XDhT/MoCEPmRfj45uVOw9+TkkUnd
KQh/VlSRXuH1HRMgkmPhYoaIUxsvy+Vxy7PTQpyl+p2AGfcytggxlrlXnC6LNkD9
j5M5BTfgH1KUvyVAQdD1bmXsbOvPiyqik/kbEiNXWZCzoFxfTPmSJEdkCZrNyE9+
NlJUfBdBB/ofB67BNWhWChQqzZEIohsWDcaXFF3KEzwIWxGqOlaI6DVzi431hlsc
LetFPO8tP+4gwSEP40KCl4gtTcAsRBks+PB6LSil2OPlmHGD8DKLI07eazNzCqpg
i84iXMWwPSrWwyUWcRhlteaSKgJy+YF995MX/mNyTku+At9YPh+yO4Yg+KsYJmv+
NGt8/bdW2vGpxP71km40z5tCXzAvbnfknwrnyVhg1p7ZVaVSpTwbtOyEG+uBL3OM
MtJKXk6NFOyYUzXDNzSbrgnjpW9UohxGsfP8LDAXcBWLMgFleUvRT5QkUrKKAiDx
kcrfrfX1GI/EsIiKsgt0Kx+64rEeBAa+R/WhuNpLdLFFRHs/26VcJqzE9Il/sLMz
vkDOt1fTSp5SsIhgencnKelxU8/7SCmSIuhEIxn8/8C8CcJMZJeP5STlW4ZNQEMQ
JuO0aw/Y8K7XLWG1aaAoPUxtKf1j2I/cnfLesrreePFXKPEKKqoOs6VTfQhsd1+V
vtUD9V55sJCByvpwmByMIrtWf8Dbn3Y93x0gpPuGJT8Hn/O40rBQVaWhd92W/XbC
EO5V+M/AdeycZIVT2vkon1ZGKnZEuzdcHytunoa6rrrMbxRMC2Q/gG//LHKMl1cf
pgZ+G9XfHuJXRiZFiFNc6cuoznwwS9jyPi30DsIVuMn5CBFeOqMKhymRbKj5Zy6o
jj9UFimgiPlQL80+zh2vZTd40W7SeDF4Iy9/LlbybiUAjxf1HJq/mL3l46CqKBbm
zo7fulpFazo9up+DZlE10JKOmrpvfh7/0XbxdLUu4XER2cPQGmYItAEqwghacoi6
A98rBVW6vXJGKffm3h9KHp9sWcZeHCueP9Ons66jJq2WuWeMASuAKxkJzZYGeAR1
wk3zUR2zZBEjBGMXRxMJX9EavF30irPtQ9W2K+liqkppigOOIsz+4c+ON2giNS6S
9F4FGx3Er5fl2MLM2FfaXxaZJJdnFH+WE+T1PuVbUYAUKfLTNPcFSdR9ZMJG/SrX
mp4JssrFDkVZdAAFNUYL18N2EyjkuZOl5NftdlPqXGDbOxklQZJI2Y6RPGh0vW7Y
6qmI9H9+TEwOM4U2Fa+89Yt4HmOLQaOFonRs4w43Eky6YA1DmGOYgKz6zX0+xbu7
EgH+86a2L0+HRgcBcsLVxNG3RiDhlXv3yNQE8ANnEc9FUWEmRJeo6wSzYcztupjF
kRyliQy/cAx6faHNOEJyR8VTODk0sceg1Z3qHq1Yvsfkaqc16HsTStnoP1P8Nj71
miYvm7kFV4CmTyKl3vCdvmU+BAJIGW52uvaV7VdEXqDXu9ngyoDr2Jct+fJBz91b
wNzn3cCaBxn/a4rbxDn6W62c8cAKozSlbXjdglM5Sfnu7MngTMqGXlICATkBLz06
ce+gPzsAeRJ1EE6YYhIxXCTJwX+fRyexqGJX3Pa8U6ib6BSpMdqOms+caj/VJYMW
sjiMUYIBOFl9PUZXpMd9lw1InW45tTM/WSRbQxEC4xlheBZTwLfzQXwd6lOWBmhf
FnkcM9w4CA0P7Pp83q/pYl1fLBKpW2aEZScy3PuQfzxt9nxZoEH5ipv9vyTdvqnI
DJdmacHQsDMP4uWNFGfvD2N9fSgaR6mdxjrB+tt/ZeSjPfGJ4lEaH5yCmVLlCQn6
sMKT3Rfeq7ZAZE/HxY5DdDNQN5sIyZmlQT/DSHF9MwH2VHFQ96Fd1n/Bb0r1dM4s
a2D5BHi0W8pgwx3ZIciTfOuvSs12Mi87vlRSG5Qr37mZB5iOPioURXeTbK3kSv1a
z38iUAjHnTPfg0CLIhvNI258O2lNMQ3zdW/+OitpGGkUZRYJGkJIzTK3U0Yk8leP
M1aleQddZMb/GDtFGRPGurOvyUxajH1p3J/czV/ptLWtmo2VsErFFnFoPvgeLy52
pLXEm/wzWqZCbeMsKHCD/rdVc0idlWtt9LukcarzPNb0qT5oP+a4T4kWm84f8sjw
nu2RYVa+2YoN4ffF9OI8KX8JKKf6zjFhLEd1J2awJ6zqyynLv3Fwl2TocDh6Ziqj
2mAi3lW4+/LcgbXESEVhXk0T4za4Y0U6oh348WeHfzA6BjrhA2cDumr5Ki2PzQFF
tzflmyvzuU6KRdK+0mC7DqxbOVVlzMw+2M1vc8U8clciSpQSM25rVcGnCy+B+keJ
JG9ZAJc/86s2DRn/icOHIKi0Xl6fQ2ICNeEQKPTVTWQqGcMqiz6ti9VCyFFewB/4
QouLabC/FEE7wxKhppjbKe+ttqSNLRCT/BD2nGBLdi5TeTxXh/C0O5Fg/fDlAyh9
YKKNqsYSektBV8tCfOWcq9w4W0cQ1o+9ASGyTsb4ij0OhczWwiPIha0UMIIGYqL9
/Nm7Hqr0f9hrhIugi70VvGABYgWzkDTaFY2pRaTtLLz7u1BR628s6+l1LQ63WCwH
tJM93u8VckciThleOcB3GoJdLCac0glpP7lDcF++ylCS3eXb1F8tRqwtxmpG9aPL
sHWYo3k/ZuJ7ev3Q0LItEkruOKsF+/rIHKXkIMUAkTpC5j2WXZYSkafo9Hr1iPR3
Dge57zu5ves/o+mYTXDx8QVk1ZloCB6lS0LS283XgmbUzO82UTTrtmWD5253GsaB
68ECCpjceyL3lNB9pWSmsZbNo3kjrIkm97dCNZM85Ntg8X64forV3EHlqwimLdaD
5AMyBa/K5COqAtHJfrp1ONDqDCLUNlFqfcyK/wANTANEojxf2mWNiuSVlGWxKiJ/
S46Thi8VTpICL2BYFbisYArGmuvZkSSxnhHgAtb5CBgBwuWnmRd5l/EJjQT1eAy+
6wFdEoa1aW3NFM+8ohv2laXL6A9eU5Ivz2sZt9GAu+GY+fIL4B1mBhWws8GV2Oa9
hDTV0imvdH7xPlW+FU/Y6zPsW1QpXPuu8UfDmordtHEqwwCiECn2+pcVr4RiJvD5
0PmvATxhjXqrr9Oiv3uPH4dvCBrf/ESKj+mqqcoOl5jFkHe4IwIcUk92EKkFrmyU
ceTRY1M9TIGKIz7Qedht7G4XkKjwm/G7e1ajHPiAYTxKxez7Alr+7ZURJnXJ3ozo
J6KTl9SWt34sxfKoLlFb4a7F4+RQ2uxTv5+bE7YxjhpoHe9C1oQFiTvQL6U/cOfr
3SGVH6Twi+Tto0yoVeqXXLRX5h3CrSLUexUkpRQVssX4ZZhlldhgE3zg8lrKeH9P
+J4WQ4OMrOVmFEysN/ZCSJajM0uK300v3Z4QzoHxdni9o+JrizTi+OASByXvIPK3
YTHnpPoC7BrYAtLCXiGj7lwXWDdOzEoDkkjW+dzyFW9q33oBbBBsd3xwV4flKDdg
FRVAwztgUNqQC5qv38cUmOR7SJu3aeoiVVtUQjwoMH7YAyqhbq+5FO3WafoFXE32
Sb/2zUg0KjsAMoD/SBoh551KFqWT+sNc4KbCowhzz9d5W9VeIbxqkGLRhGAeBNfC
Xv3voJVUFFl31o/gfB3gAfoSBz6JJ9GM3FHyyywA9Kucx4prLZ6xKoa3votqjqvn
ZsiFn7AHd9cWQYQ/eUg8W6aECi7VCzc7A9sL7jr12CaE4rA6zQClBqvXWspQkaKd
QG4oC6j08Yn8203wVt0PUhxV2RUalaF4t014LCe13I1Q+sTuj04/AxfbYCtWatUh
nmIlufds5KhHQpIakQaTaU3zp9HhjA5/SIl7W3JEviMv/Q6MPp8mprjfRPvNeEO4
7fdMGoqdqGe59NObF1Is6D5dFohfZUYNiwIdl28C9nDvX1hiIMngkD4A/R76s4Ia
D2nRiys8ichslX5U/kH9CQ0nhSbBNTtjoi8rmMJS7kQcBEmWg8MwmMwzrbIhsaf3
JIdU9GH82ESEoR9igObtPbdeNvcv+WAZxvPxVxyhiBkJeAJsJ95k860gIxJFpnQF
lkjLL8UeuA52hJgT3Pa46L9iwCB2JtEOdrNParzHSrAwYxImztLE5k7e3TLFJZXM
9Uun9fw4MyDgA5TILgPQM4EKUE4Quo9AFi966sSbPDp402qgizR7sOu4eAaqqLbq
d4fmrj/HI/I7b5c6h8R+oY4tP48bTOcr1sJa4OMXBEQhJ5fpfrTIdnLIWkQMYBgc
zGOmP2bBCacbZBqO1MSCQFXgdIMX7bcrq+3FLKCRUe9V3sSRm+tokI46UQCqvY2w
zvn9mJBAGfi4b7z19XqfQ7I0mi1M+58VniY1oKllUP4+Kdiv7O5ObGcADz16h0Cp
xh0x61sb/YH7DmReOd+sxBGoO97GsYyz+LSAzQSU6CxApu7dDXK/SSNG0n6nwFR8
8nms7HUtytNhIath+N9ZMHBVHJGRFgVrZBQZ/RLTvCPjbCvxLuXKCC2rHCbUn0X6
6HO+UWU6b4zfYEAeuz40Huxi3fnXIxyaJXutNRHVV6W1uGiztAhvoxwTivhFoJTk
FXdRtiz5zMuso0NxCqrzKDg2d2apbggMjNHoKU/vzA+LJzukRWOOBCBQ/CYZi1yF
Ipmxob7zTiOb7n7SgAQgLlHkPL8ZpRWMZQ0oYJ7C5AcKZu2LK2Nex6fCXn3w6Ef0
Jm2kSkUp+RUPcHrLCX2QNJd0dYRtVzscCTkQes+2IofywhEkei6pN8lRbb42dtEr
I23uYgmnHSxfEXauRM1I2eIuqfdvI0F4POLoi+nbRmXDeZXi5H/7Lq03+yrKOJN2
gpshNVR05sq+g7CElQ1TTIuaTW4Yqk4UwbMMZ/UkU8pElqSCu+5idAxsPS5EoT4j
fr12+b4hWDxy/K2fnq/pUt4yC8g5O5m+XabfVeZ3da/1u2A3GctsLPvEDMBKO+nH
BVbDi9Eg+iWvtrSKbLLzVwqWp1OPE7gxpjifjsVu7E6shg7QNZTL19NBHrKn3Dbt
B1O4vO9+BxiwFnzuUOqrxwySgwxY7reWVc6zrONBb19fsqvHuCOTF7n6fckgls/C
avomIyqDfwdDw213m35Nq8AuBF5EPAgH6DsI9GdV+ndIgn3JmG7weyL16i2nJdcT
kW4oM5BUZc/vKqZgRz4lRTgnBMano3IxiG76o4ScDRDdXf1m+qFGtzV9SoE2/g6+
gKSPhQk/FBAv7AWb7povzzHDQO4NfOO6UQeNqGqFllnTKAni+Kpx5n+ypICSt0BO
ZfI3qM0LG7rdS6IF0RtjK3dKb1azgnuhakhyx6p43xsRFrPIMiIfsV/SlSaMJSYf
EHbeOJ5M+aCXJ2AYx7wUYJXmiv9VvD7uB8n+tLJ7iJUGBGjM1G97XYVz8knWxhxl
5sgzdg8Uj0rwPzgtnPQNGtsH6kkvCxnVEDdUOnjDNuq0gtr599dH3M0R+O8sXrSM
CaX111ryVkMGNmMDvFxYE1eFlIqiB8j9UVj/CPq/mkVIOmhX1TEbVa4tNB/MhISX
r3wjhWB4RbCdYPsQ1cA2hhZMZ9oC/8CnTDR7m6Nojfksg5G5MLcmotfGMGe4jyQE
DOxvdSGQQc9WS7AU/3xkYi9quRIVZ2EiJLnBbx5YbYW77E+RrtS83J9ZmhK1V2PS
cO9LaulSINWnh2JCiyHOZyCe0GFLr5/WzgRtBpwA+OLY0G1V/vLOlimxvtGLTSy6
dszS418DgkFleYYipNkVJpX+LqIi9srDd8KhxqKu0EM3MtnXY8XCAJ6Aa7ZvV1Vr
TPgj8YrK3P6G4xCY0y1iixfmz/isf/NSw0g0AKDZ3jtiQgE1pqM58W3gmfKWiTn8
h1R6QNfzqC0GMyySz27fm/guyUqpRZzsNk0aLjAHwTpe9jeJ7cZXzqCc2eI/qIBA
kF+uNQmLcuCIegtp9T1cxMY7ektKb1onqHDRL3Aw1Yxac+ymvSSpam3tDQL29dVT
PbhxznmA6/voE2ziKY2WNNGItjjsrBGyb+1E4I0PZ7Zk4d8tQvxe4fdlfAnRWePu
WSDyyEXOR42MyqXAUHxjq1iOs+kZhTgvg3ZVuDEXtEiHaIyUJtbdxeMXURgjEhpA
jSN9hKyhWy2debiIazPGqoiEAsRmdMXSnE+3z0Xz5gPK06YPouTaG85lLeU99Chl
7Y9G6hODT0pau6wZ+3EykCiIyG2iXqXgv7hfs+N3bR43mp2HkZXZMz5naX65vo7g
v/nJaVFs+fFwhcjTD/Q91q62MSzwSeoF8FDcntOREz+2S9VRY31eY3rkxRsjLQoM
J+9m8Ft5Dx2vZ4KFOAAriCKNpk/t3sSXm6gAsgb7z7jFHCsVK/TTppnyOoCNe3MA
LGDFVoWgyZe/N51Q+xg7B6hJ3o6c19zGKTjMRLB1WvTCYG8/+plh9rHX0DSsV8Yx
OExtziCd+ZiAf30q+/+oe6rqWar1Ujsz7U0Ib3Wc4kTL7Y1rOCG59RyqQVsj+I6P
lJtUIXFHElbPyO43BkbQn0EyhzEJ+m5a5qLVnib+8MAnZSltd2Smo2DGWtMjZDiR
iGwir+3zUgJOlEtKeba4rkIokCkLbt4kqtgBx71Cl2D2i6XpHzTJpOvPlcEXbxcK
lkKyyNQ7KWN0oH3lLc8xTWoeqDsmPMFpkRIgGhFd95JBsFAW7bV6CNqxHTwIqJzu
r+Tb6FGYSPsqPyAgSeDCu+47vbl9xD+3dbY/NMZ1OIyobM40sqfXwRK3xnO83u84
En3wEUju/zN0z5xisfUeIsDxGcxYwiKfzPdctsA7ryksLNwH+rgaKWyGcdq7KZQK
TTL0CyGGFKoIP3eBAYn+DBzxknIjlVWnglzw2eXKUIOQAvC6lFhBAn+2/f93tj0e
JDz6aiBCgAfn8vw5HzPRi1b2WwyO3qjjLMwLSiFL89o4iCjVafJLspsScAMNMvKZ
jjdteS/a7EfF7AaDDad4G3xp4h0O/oCrOVYKlDvek/R3+mvpbu+7CNmUZofPxMG4
KqcD/eTD6w5ZRspPIngg72FCa/kWWZXlKjyQlFi8toaSKWw2/d9xCS/9tWCfv2dS
2G3NDFmcigpRsxMpUwsgF0vX8U3c/jql5IGqPWK2AWAp5GxSYCqKLXiNFLBRVlMI
+v0rlfcWi5atGX0ymH6eCripBXlqgxh9wY6ubxZ5BnXRF+TBjJVVg4gR5bIeB4Jr
JXj3SfjV5L6XoSB4v2V4ykQFozI1ls5QCN2Q82oZEjci+n5wO/nOaiXg9qxOwmpG
JPMEd/sT52agf6tlrlG1pk96OXEYHQFS383DogC4TZWETki23Nn73CrOVeGQrXms
EcKkEdz0zIwXXMA8zPvj/gpJokckeAJH30JZQHtZj/0E8F7jNR/zt0QBDZ3eMIPE
gzdVxOvoiBZOwEPOVW6lPS3CyCGKxpXeI/TdMDa6L03QnnLj0CSvF67Js6p0mkw4
jfaSEEOagReyBDARCLQ1foLa1FGXLgfB29bowZnkTG4Xn/Uxk6Jzg9Zso1AOcoDG
Q4y4lHBhsb6l7ZAfhQA1NOOzSQtHkj+AAy36RhBnJ8Zdm2cXLcsKj6vUlRQDLyQZ
0AjUfruvmzGQtbJpiNUaEbt3PPyKsVa5U8u9UQyTA+0sfKb2QD9G5zFNtTz6ldDP
oiKv1pn/6dxIXMCf4WbCe9EXlX3p/Pgn2eemixxl7EIF7C8aZXxeIBFyiA8FIta0
FEYSGKxAue45/93RzsjaatwrJQ1Bh8f50/4FRGsADpGOn+zZY8y+nTlOKcHgFQ14
Gb5zRWzytX8qEuMffyZjrgFMfZnLdf+mHOkxega1oHt/jCNffOuuhMdklCfMDy5j
7mjxhqoj0n4b0+4SgiaZK09wYldN8WXVEOs9CqFom6y3sL+etdW43Q70a99BrHPU
yXal8gQxOxV9qGas0NvrXp20yozNokFjfMve7SRwxXQaR8YVR9nLG8QQ9LOJw0ta
OfPgiUB1HiBuxnckwyezLOZ8s2d2pN099oKhx4ZHlPKGUXvYdzxyqhmee6PcvRNu
T+GWw4rEno67M/Z+QYDxHwAUHqP3tCNRIMJn4UiUAglYy4dgD9n8JUta2UMYfdnJ
EZMhPqQt9MGkVywcz4+S2hRSb11BZdVNDsLyUuFMHbPrOPWDKIzApst//MV4gBVB
AiHhxxXgatuaYxL1q32uztd7Hvex2XcSE1EirwMT86vkHfhYUcGF47mCIrZmjTJt
nuyTFFnqoKSIj8WjFBf7G/jIiBHttqIF/UkR2WjQX5Mh8Nf1T0kM/faway6grn2y
hx4x/KeXMO+iO0HfCMWoIfoRiVu4d8yzKZEAmg/T6qttiUUUln3csurB2FdZrWaq
bybENKHSvmiUlTRRPwDk8NhHsVU2MizHYv81hP2D2yw0hkrjdN/1+D2pUv/x8W9+
KAhPrb1NWEbGkpSB461u7UPmO9d1Gw+3rCzZ1NsK5D97PKQekczyPODe17GQk+Bs
0hcFIQzwohVRwn3jfegyeo3JH7uUdC5zYGosYRC76ybFT06wDEePCPfyXOR0QFmm
xWBrxceCvv92ufvMYMeDBWv2xiaKagsMSfKssx0WmMGGtT+zb/0WwvR2DFwiZQ+w
OFwkp+VsyXeUdTuyHgQtQQgfc0S1STPICnlYcQcaxyH7K2plt+OeONLy7jmhwxgD
P+iURqYNS2UVNL4q0Qr+PN+/+IDWI965qRLQ16qE9w9sTM+e8YvmHCOQGgb8Hn9g
roSEX5b/oqptUOjimM3Pz125MgJ+Pq47LSLwd2bM8ZJYVhO+5IbHrIyacAtOJtP4
UiSu9t4HS4pCwUXvepISE35R95L0vluQTNMmaEYDE+WK1EvoEw6gH1dy7MhO/mBQ
VvhUtfYjlmDQshW5twR9Ha7YsywfMlX7Uj8M9w80BwKqTYS8zraBeXlXpJzKoehX
vOrcN30o8gsqaSgYrkOpwZ70xv9JrqH9W6DXTPeTEi2qo94Jgjx3pcBSf5axA9rA
nNOgRsSd+/y5RmWUSPWgXPjCOrYI6uy6YS+oO6C4RkashJ6gtjkeunH9h0s0q+c4
fNi5P7wNSj9BTHHsHeZc/vgNqYRu0BjmNPA2f40wDaL/eRZ2flv3Fru1qO6Wxc/d
Av9t2fvzuaGbnBraOxNrsygT4aETEEJ8gp+RUngApjoV8J8HbStWX9ri7ekqnRkC
x/iIblRjkBqgmwHZpmoDxdu33vrC/gXoX5FtjXi7hlgHMTYo6H/hXKyADJr6oKWm
Zm112o92HqWN8TcijzyRZTsrcYSPzH6z3bLsskz70YfpzhWEOUF1sZBrx30qSfJH
jEnom5hREurZ2dTmcdmJPCQdr3zD0YsoyhwnuuGKmlr0Dnd4TboF8sVQXN/xmvKS
9MJtNlPsCYE7EQErZ7UTyrCQDoe0wDP/WI7QPUDtFkz+vii7uOtsaOoe1QQb6lup
6yF65f1VIzBHH/PXO7jcAXeLOPOhaHrhDNmwjNu2RVe060D8An0RwzrHYFUDhTcp
2P39P++omrJOma1wExXsjdBoFSv0TnnL/r/WcNjc0HprQSAYWf5lhmsaPPWYMZ1G
q5DU/BbYHOj4Wi2D4OAwoSFUkztqipp3Y4u4Nxjhgy7InUKKAKzgK96dQk2BlIrJ
v6/XKWMt5Zq6cevOJD4r6iVBDa6EUN5kIC8si16P7xtHp+shcDyRFEYmTEP46D5L
DX8iYyqo6lVNXyYbZr76Z0DWXV7own3Vw9b3dB04KacUhZ67cbcj/sm5vPFcNRie
4rDTiE6LvsBPHAVYjISTm4JIdqmhOryF/i8/+UFl0KniiEWbjaX89bFILTP9rVPC
rYNhhbfUlQO7tdLqvkrCol5yfl4a/Ep9h48xp8/a9sMprQduwsJsqc81zOtHajpI
mnrycysJQ/QKWek8cjvz7zX+ADdJz5N3Pb9Lh8zAZfcfWO46Ylyo8AFBsWTbXHCL
W4JzjC4Mq0xRjFMIk8EGEfev97dyau19YMpWFuFrhUNBI96T7TT/59iCN9D5eZTx
MjemtJ4q5yu/2j86JCNiD7q5EceRHY9ZZhgimq34PbKBNMGkl3GX1uFBGK3ook+6
L2t/uLm8tzkPZA46MsJH/tu43dyrRAmFlnPEfwwLlIRH+FGTWxDHBYUiu1m4Tgg4
AzH61GjsCTpbiPeK9DTwx+NNtxzP92hTxXs5FcKq6BhSskUrTtm58e916BJDkkih
Xil49e9fKDv+IU577LL9hio4+3c5Njf5WVkHBgUAZ/SeXyXaERrC5CwNwo/2c9nk
EJ9ei/GNZQzaDt5hRRWGnX9ZkoflgvFVpDF9HAZ+eQ4AakY+tPDa0KA85qH/+TEe
EjWfqC8ikCrz64Ag+fUlXO3LvSga9Y3Dk7/EqHKkZTD7QLvXWrW03AWTaSE7JITN
IjK5joTRqB+Ny+H3yIKV3S1d8/5/dMIfoBfwFsmFICbsnxGh6iIs95mOpYhsLuw7
ZgO3N9vrR6krnKS4ovShHXJTISHoqfFA6ED8GDXylhzWiiMpgMjlQh0ELWdkoKae
qVxwleBcZadtFOKcxdX8vm+4rcFakqBCAqtTLphZkZjt0zp9mdsWoBOj7e9shT/c
U4RFEhe559tTMXNdD3LueE7DOWc7kkzrIKYcjqLO0wkNHbnnjTnH2KlLKYJYGYuz
MPqZdJbtoVVrk0lwQs5tGOyTLnrF0rd5iFefhRgD4xz9Wtl27LuSDJzlVWQkZHai
XiO/R9oG+C0d3jGNG3k32gf7NJlW7uyezqREq5AT/yc82/Z0YGLE68YND7+xFF9D
+rpgHcUTk98NLhwMYyZRk00PkC7rzhd+1n8aYFcRjA4B2mZ12DSJFo1hRiAPxTyP
qIi9/AcR5f8pcNOjXNsRLh7o43dWA25zTx+QDFXroLN8xNkVVhrNUhujeY0BoENF
06nTXy4XiQe5lqx1xeJMAYDYmyZ7H2wg11z5+8SVTeGtewxinWf5Y57fGBRWLdo4
Kovc0MkNJ3wteDengLZ7VgY9z1MFgcf1Vc3JSPctWuElRUPTRdsx46gBSXrZGNlQ
OiJu1f2YCJAHT1NNTg3eq2r5qUa5x34XLpJkgVV2NSO5Gxco1zcuYF4EWRG1hbHv
izfENavGp+vHZ8NdVBNDADfEy2mtEJqQfvinLqmuYJfsEPvCEWkKb9bseCEzfx49
UaaLF8yQHi3muUfTpxXNacmH2YDcWam3uqw2kvkxpRKcmASKaJdHfzyMlrL/nlk1
PS7b0UepDy3NWGZgcuGE2ESj87qaYkVnJ2u9nadW9DMHwpycwdC2Zc+MRpfUYBtN
1Rm/QJ0mqwDo7W+xftSmToRuHWT90gr030XG0bg0p4boOWIWFTQ9XkkyWuXgUrEG
lFeUxkeoUbF20GyxwSM8rVNVaRIEwUxdWa4TzBq63EogMT/rmz3N0mqR4234jB+H
p08oZKQq647kYeN8rG+BO57FoXrHvOKZlP023y+qLgQ8Myuz+DzAf0SwtaTVvVua
UvX9aHXbLhoyzKKTJK/GeHHKgljvqQ6Wjfoq3YS/aXe9ABN+2mhM3NgqeVlkXXFH
/Y3zaWjSgBbzHwH119tV+mZUTmMtcuEaGJjpUOoey4EKWY5H6HJWezP0m+tMBBq2
ZsiU52QgPmDtVKxezQDVAPa+hPotqpwmIxUQrSpaDhC5rGQFYhG6SFJY5X6qS2XM
xn5+NnPqXknrEPRyWjs0B9g6uK5HADl7RAK+G4qIr7PHyIF4FjUxze9OylMng7eT
WPyMV4XRE/TSKFW48ShcnqKulPeJlDCcCEEhwBr9BwDGydZ686UjLKop3Pnb3xM3
bFZdxyVaMBZFIQoulY89dD0d8tfL2FZbJTu2Hwbow5SnhMuKwRqNbUEQlKjJGcmh
8lhtaCK187MFeWcL71wLWuOZH8J58SNQXo5gd2vU4dvvorACyxGG+iAmUhgN2yXy
PbP+LjSTIYiP/c836Q1+EWPSK1CxQa3NsCbX62346VOIY8aLqAbUqK9e2OzmlKuv
acrlvjmt4W7aBXIxnBCmbLAaFjsQosvy8zokjmtvmrBzMpiyLTBmGk/7m8wb6wqm
z9TD8ZiRkh9aTgdLEM4bH9xte1IzNuoem2c5X1DBNg61n0N3CgN4/yKpFFSsNsWh
VED3d7P71FyUSjVb9MAxfJtw+wQP/Oxw7qlh2k9G/flbFDP4uslnMBmlRoCYsWtT
i6QmMzyckMU+HAvI3uypfzgcKLWbTFCjn3D1gVqSjBsWUZkTvBqLVx77Um9JCerf
jQ9WL5WGDaFxUVHX9ZlGf//n9sHX71NKgOd/+NVp3Kk0MM89+DM/B1rAAg8Af6i8
GvCEdwKh6G6+SlfFtpAxfZSjcsNAX/f9xIxP4FMVLh7ylC8mcIQNMppE5ikguNqy
RWw/v4ulNgGSUYCR40PoveK4cwpTbzLcQjcXe+38VBayfTdphZDk5+X1lHioZXip
qfnQ9NPsAiZhlPAJ9/sz+nP8hrhHLJs4jjSczs5tEpfe3VEaNBntB4bGPwOa7jKD
wp5ETBBEJkPbFtuEy4q+rhtxQ7j1YfUJSmZNeniMmlJkLqVpQWt+uA6glr2d7Rvm
E7dFgmHawDLVZhvG9m2+RqYjekJ00mpL4bkB8lVRArvsWBZk9iqmAf7mnSCM+/T3
DZxkCrAKgHlRwQy/1mPDpY8Cut9vQa5yIveI2CQ6G+Xh5gVQrH+78eCiM9KbQ7E3
ruNDJKSsDHEP9ueBigYLOJpmRIMcl55p5VP9OWgjphSbifFIdctS539fuOnqRBBO
ZFU+JWiYJH9rDeJLVHHUrfyE/lohjH0xwH2aOGe6tjD8RedtHpxR60auQtKV495V
GZJ4pHep1z85B+z1OwSPJlC0tAYK1Ug4yHt1JoeOZhlj3fTQsLPawaZW7NWAqW0I
fh16Yxi6s1kO1ZeVveCbjccGSq0TNO+U7OgvEOhj0xgU10C5mpdhKi2Yd8Kpea/x
AgdD78d54XqE/kGQ8wKxzPFMktB57aUUAltdvHJI3Cp89HgPHZqOoXZXDojINtpx
OGTgQxKalfQyaL9k+Uorfjz4BovE9N5Dbqq1ktTQkUXYWWmYjsxZ0PSJgFaL4eN/
KfQm87NmhNIVXA7LRCXEKlj3nNGmkx6aJI6D8hWfmEotU9AcwD1vHUaXsJbnvLcq
txSG/31Q4i+OWO58knlo1gtTfjEpp9lhFYzIkN749jBKJOgUP2WZ9KRHlGyaZlVT
cIZpEV6MSv3tnycG8+Lc8DfWUIoKbosNfKVjb20RUQKDys2b4NyfCVvV8Jf8kq2s
hZ1gFHHq8HEOqd38m4/YpX8B+Tw7ueckmwKjHT/DvnL293Us/4dCyddTgWPhZwF1
W7Cf+LVuQDTLiz3Wkuqhc1xRywn/ZyJn0CDqHR2KT9dmEYe5VDx9Ic+nd4NQrIoV
o/eThDYsc1Vtfio6AMJsTi//DYBhGoC+buuLVqsnnsnNU65OJRIUiXLaSpRV9dcP
OoJ7nTCeWTTE6GqfKxLtGB6d6VU9rFt/b8VMu0cc5RuzFvIi5q7ra4VTF86y1/sS
gtMnwG5Lqnq2yyZrVxKex5I8dd03r9rEccbm1LLw49ycZA6R5uZjFNeTwfORCLXg
Rs90xbFqvxYw/oUGDN/pRg1ecMJiGjhP/RFavudCwkappLoCCrHfBT9wfFtKlVyt
7ahT/pAJeYBFmJIZLn4bU6cBO4SPTt92sFIo3+HZvaGKO8zniswR2aVpsLicJTvr
bejutcSO+FAEIKdAArLlL92DdxbQxfG5ezA6tPJhPZmucdUClBiverKivtONyF9Y
yWc7ZHamNBzmYxZyRgw+g15Ch92Ozz38A/z+0YqLscQLt+4ylmjjFat+AqWJVIQZ
O9tAf0Babt0PKVrMPuzZmtZEW8QAIevM+jCDsl9frelHv4drgHVoNgqJeeiR08C+
1/mtBCPphz1BKrliBj/023UsRwXTUkN/MaFE0zqefO84B290FxgvMamnoOxfHjuy
5M0e5lOsGEJeLKJHQDjktMJmvuObVwZDoVUJWYkQq6lgVxlY95J7hpblEqq+KNyy
ZIzoSfYxs5quP0/KKY4JCNkX8Zp3jhwG4euvvgXabEAhK7+g0axy7haXw/uPXRJZ
Xgo3O1iFyVdB6D02GGNSqHZNY+D2E8jBJAtqqbDGO7z9HbSb90fZCv5JZ8HCE1zv
ZIt2UpE4nnFbeB05R/AFfovDwxCOXb20Sd4ALhNC0d5u7J89ZMs936Qfj4F1zH4V
7QrzceRpYZYBPXwFUqIV/0KOM804dpf3GulfxjeUjMDr92lSLNQSUAwajwpmWNEs
ZdmnNbk+V8SzFFGDQD19b9GTra/OYP+AQ/8GJfpzizGxelvDzXoeAnNh4STd8AMN
HM0GobmQNycGnaOnOI5sr95ymtpNeJ7m9cfYGCC0lwIegSfAHjEjlEWFATQCjT+C
4JeWnntZ6IKrRoS4+U7VrYruOLGWrw/MfA+8NM2LbZ3P6+EpXpSYr1gtpbanp/XB
X1PHNHrSOUpzuJbk9l/8ZxCBdFNIJ/bN18xVs3zegufoUphuIdxyjDfUxlNMdL6W
EqfFHA+4QFuc7gLK9JnHXPosG06JFITINrpwPtgWYLdGDGMv/9LQkBtJ4JLzLePk
puPHWfM9raF/5kYAPcZRM7J3Im/fGcfLjnpmAIdcJ6eOINR6CrsGuBZ456h6V9Jq
joPdaTBeASJTvgrT0YHmpo4dsk7hf4APAPR1UvrJzt3y8uTEuJHqGl+65gracNY2
XpkF7eR5B7cPgi5rfDnEuNQ4G5sceRZNW2sn8t9BcxvE/5aiXZ/dPOwNeRp4iEL8
ZAi4e8h1zp3FH6FhmgsdqNuMmf0jMldBjfC0co45a5Le8m/6XZno1P5p+r1yr12B
yCcSWv9hoRRbkRdcedhyOS8IdDbo2bXB7N36pmbSIsL57DpyeKxRdVEucCLELHI6
AwfrIcpXYR6CS/d4LuN24E4F9I0y+JLsDpsu49l4Vi7wpoGjZqdsChJqt+mHkw1x
ljhXd/sv7H5EY3iATHlh+/z4hK3HDlxRzVrCnvLWi2HAsdxBKt8bDXvvx08yifbU
DryJ5TFTg87mPPjMQXzmIxkzq1zNonNfFy4F8Cktyn3ya6nOrbqRPzGfSs9NVeMZ
Qx1HGzYAyupbFPrTUrnmuFpHneA5JTXlLNeFDvyf+izcDi5vJpVbiqVbIcZ+sEOy
8jHrhs4jHLzz8OyNnG/KuvMABIi8O/xXe+ckW7ZEQ+VXIVVCxRiQqHXdlnzedSrv
RhHMX/7NsO7b8f0N1/CgbbuUcDYUXX9OSLG/Txud1uxsc284VWXM2KH+XjMmyMqG
lFU9VKnYALuZJgg4o5hrIx71ARDI3Sx5pNz41te8XQZDoS0qexsJqjJIiMd/vo/E
/4+pHjAkYvgnl2RUYmdRvTwlou1MICV+I3l41FIQxox0jPuuWHaERMKJ8vOK9Dcl
36AgzlOCnw3w3c/doMtRxnsTwVmY6lIErBIc0Ik/21FB8rnYKa9DYcoo93iu/45U
YZWFj2lrqO/RP4kiORvftmpycVbg48GD6rRU37E6JX8ELIdLf4+K9Jx/JCJ1SFYn
/+JF6BTPuKyb1iotXBpz4gf6LfnvGxaw9PMPUq9GyuHpO+w3YWDh+PSvlLYfALmb
rE5cOaVMqmpe8E1Pm+DfTg1/FhZcidNEtNCuOlXRSVnkVvq7uttHYeaxWdkjkKo5
dq/nCuGmQ+Oa78IBgKz7kmU/MaytAal+udPLhQM1+iGd09LM8k5Iu5QLKghw9tUW
fotlxrFCMOiS4EvvoCVg5OeX4/igGP0MMgSY9sDPGVDpmCFK6nxXYGAlDTn9flp+
Cse5OiwbRJDcTKxSts5FTd9zoG4nYLoBvYdmKSGPIeqW/EdHakix25mkaBjZYl+Z
TitT91CQFbv87eFuCVuARG/6t6PwwgjC/XX0KnyaVx7iInuOHEvoBHQaInAmCx8d
qgj+1nOdvNPuEze0USKjCA94qoE1E1HZcCq5IGbzGleRGDOMQkxLP/35jkh8+y2E
LZOW0MusP0NFtx6MEo9pdG7vBx0O6xsG0n75ULomk3xr6JiqbGe8Ck+cWIMB602J
zzoetvFI2tQKkT14LhYx7LkCh+AN/GvzTlqOxiSyGKAVt4wBs9HUiZrF71j7xy1s
o1u0NgXsbpSR9iyP9cH+PpQIewvMkGaZ63QYpAu2h+BlQZRecyhXcOEV6VxYPe3X
dM4LTQd0ez/UUWhVfk0omG2thqgK4qIFGkggIyOlBr6rLjCSggTsAzwqBe0g3HJV
TVMlUy8MJJuxXl8LrU+fXiG3hvm9SR5iATGHsL7sDBRvOXQd5Ga3qFCXS+7pnJQG
fIWLLhUuWF3FAiRh0yfYeCqESMI6DXrygDSAFOQxD9txn/3vY2OFtN/b9mID+Yno
YFoo3GH5Qoa6k1UfVcunQnptHofiNLfAaCzp3Ehx7oTYnjbZNukGG+36rFY+qpLc
XUpL4wU0hbTBc5elnRp2E0pU92/QHIuS6IuqC5jsACweFxfKm0Fte2xTtvvyANID
mrEXCYcvlbF8B5vbMWeOeOTihDUoQAUi12W75T1ELStlLZHhihtomvhYRknJ0FPg
d9qUvyt/T0JXge2uK1AK+67mEm662jSAm9VU7a6kXrxzFSRg8fr8rUIQwbv1JFBM
zn9eZQy8hmM3zkjp1c8foCWpX8Cdqtz3KMh5Z2mimSEvXuqa/TtqwjJZxq/NDcpA
dvv1VeI9KL2r+6UiE6lnU3/seCXjKBFADKJylAiQq1uIlePoKnQfxQM+xbTVefH/
EHJGuGLhFv2NfwExWjxhEBuQh11Tl9GbcIBvhLYoM2sn2MGowsvAN225rq5UslDI
p8GZMRtDwVS+afdN+DHoigChVtRnMir4X0AbgyOrqolbOKfbkNkA3weHkYYXnMzy
7wdjQz0Y9m2PblPPRoai9oHD0cSHfn+FwFQEoTDrBH21kO5ReufUpQrEZ7EiULIC
OAw6CEGaJQpMQMv4ek+8RleDc1OWM6JsvcmzSN4WnJIH31zzeqkUqQOeXRu7qtxA
tzwBvjN97goccIid8z9B6OJ0dA0HleMbUXZWiGCHQRj3QSn8sBsYy2dyAVkv1A/r
b6Blz8tCxYJTz+of8TjsNC2X7P6rrsgBiISlZ0xJzLcmY/YeL7X+I9gXBQZd1Oso
pPe2THDt7TwpDMD0uth6D9CGgi5Ug3Wg5ULiZ7Vc1EGPusldLV0R2CAH3tCXgatS
bcO5ZxqjRnnWaE7qTWmHHFLogLlfvonzBGe0Ln2Vt2aOAjsy8Dvau8i1312a4Ppi
aO0doj/KIRUIiHSLqtPiWb5s+D84wZ71+lOqf44GZm1+09Ph8aD6E8b1trvjZY3a
7OoGahcKpx1BiHi7/tVXyBWmQj2H+2ZQCCKhTMQ8vGzEdhUe8Hy7s0F9Y6fVhvcD
FeJzzCWuKD9254rNTteV6Hj/XbTpvXhxtT81Jki71uAErwxxDvgWT/qlqYL5UI0c
MyCAPL7S/EN2uhyur8gfkVG9KrStdEQTGforC5ElcgZ/Dl4IbBGiGtSC5EOFqC4B
oFxT/En07TWrOiauC+h2y8OaTY5m/pAkINpz+qVAaMqDKJXPtoqbWU9XNBQBI1Mi
Mt7ihamUbCb8IlirXtwAkMfEbV3eRABox8gxq6dVvTYDw3m2RvSxO67NBeUiU4wp
e6BZ9h/i8cFNfYulGGg+6VkkpbYw74DMuiJ5+sdrS8vJt4QhHY2F8V3poyYT2rZc
C1iOmTwmHgjSkoG3cvgIaJjho+c9vxL8SHlJcdiQReexge2xhDhNCmE+5PD+e+Si
qVqg7Uzte+KD92ropL0rj2q3/DwkT7in6Ftcckdm1BBxzLPAUB68Oh9/3r52awkf
+O8iwF+vpWeATgiSmfHb3pyBwyGTjEQBVlTePNiorAlg1ZL5jJrgUNJuSyqSg7VZ
790D1Slp8sfnJN2Zk+IlLffm0bgPiieNGKPqYxIERrbn5B5s8wzZ35sgIM7GsCKS
rZDoKAi56IoIYSKsQZnQDOmIosdd4Btwrb/Nkzz0rmpIQnpKuiv9KLz+CsoZxwCl
HlVspVl8yNMWy4R8J59xLBhavAbDfBqfKuTaGpd5xnPeXHN9/AvWJYV+eHWOYlil
ZUX+LQJsU0u4rHTG6oomq62xp6sdIAHEyEFHE0WsSGeLOhmk3Db34CJW2mGfNJNi
qeOsB0fn+MJkXUHFGS7H6wo2OZcCANuaS7iY+/zvEC9BvqVjENgS/MVjG9iNFbkh
biQSOjANv1aZJ7jKQ53dHLa+Yi0nSsBMwY0+/5oNteUN2Z6Pzi22uBXxf9rrhjwi
+1yRHBWkHSecveRFaH0lLC83cw68+481sE3+l9vvPUHH48YUsvHPKuas1IG10AT/
fRibfWdhoIbMf91SPYRqT6jt4TK1XJoCZ2A+QvrAFjNtbzSbkXW+97aFJEiaiMcp
Wk+yP0h0lf5WLQfBmAho0Zu6KqD51xMMIj4qbTJVsheSws/Oy1YNy8Le/pXWe0KC
t2+JaA+nJRm/n3ytW+UNKsu5pb5Oo/FuUhYLG4siWIVz/qjwVEeOWfsgfHrhH59F
sFO6W+pMBgcqJJ79VUpiWyLwgDFvPIzS2SrBvkMJ0UbUKGPF9/IM2SGyOdhTvQQo
vC8k0JGsWmKUyjGI0VuWbUd9c8AqTu0ptXI5YS6ZJr+oLdguD5J/YZ5opMzjWOtD
u7NDTJ3LFnCec0LwQbmwTCQKKhOxeAyRf3Sv38/t0vKuhXNKIvoLgOcT+Y66rD88
fu0LcSRnoOPIMvdkAQjbfQHwkUn4VfhEcVQtIcTEJFpj2p4x6oI57d2rPs2HoFVN
G7W5/M1sPzaQWtUeepeSTb79jV3m3EiXuXH8RBuuWwWnazfw6gcEt6MHSlhwvFeB
aFiwMWKxjkxPtHCI9Ah795TVQ3WGHhWk/p4GFwhgQWhJVLhSRthAKCE6bft5fN4u
jWsvq463rPZ9IaNXFy72fTRIyRMaDfiVLON1SASfXRIxtN9evZBQlu4zcKeH8KCh
CzaQcDn8F3IvAmXyTFXxhZTgF/LwTXlv1nNV8Cjtjo+y5kJYcolpw/7wuoQOKTiN
ldl5+4VZvCC79BmuWuWRhoeOcHg0g0SEZvN5EuaTsOaQctJweDWU5FblnP41RyYO
zFikH8mJHNVAfm6g19ZZwVUO4Z0zkH8VpZaWoXxTT2dX8WdfrKOqdMGDq7DROfhd
au3emivMWxSlnBm/aKryopL6sJDUfL+NfRvfJzh9TBxxM9mdLErQ2WkaEDqH6y1V
gS3SrirzGSLlLNpIZg1cIcrR4bEVh0V6r76cvWcRIv1Kk/qJixqXgjg0L62mJiq0
B/8+IbZMwsYf7muRAAQN4SVFd9PG1Ramjl8BBnlLcsTJDAux7uGiRQNyoWrgWHop
PFWYBjv9AyTxdpAxOq91i5xSszfbzL4g3ug2RbevRuHTtbzllab6fmOxPkG5KVvm
q/+B8NJRWMUy6Rn39Pe2/ax9XpT+1U60o2JynBBLpSjJkLmVZ69EZEmSru0WEU2b
ks5SKQB2LuaKTGsi5Lmxre+MTCt2FbBKPashVPfi4TBqRSwmsLvU0ObFKj3gDhdR
gaPZGjKIfWdCMTlNn4hrZ/qBxh5fBDWuWvWub4WoH7gV1huCl7ofSqeWs0VXXny+
gFAuKmN0kdWGnsa3l6PBntUE1sjPvwe9Kic/4Vi7a12DMDkc7kPDT5cRbGdJHoVZ
/2m8wz7awKKDZY/YbxVh9nYJkrlHCIH/ElnK5fSg3ZidYU47zSJajnt03zF3vJWn
QgoQ4Fv3IME92CVdOwgssh7RQ204Jgp7z3sPgycbK+FoIESEhc+kQ2mqPuK9+MSS
VkgVMT3E1hYzaMforpeU1aJ6rnTIIe0OQQCA3FJPSQ6TzuBuQpmFkXctADcFYdKf
/G05WgcwX0kDd2Wq8iLzhpgW/rc1KQ2PyUe8UKHq7FY9l4eozXQ6eyosMRwXsNGN
CNC3qGSLF+++KbOTnLb01wd20qCOds1ULp37KIBVjFe/Exd+epkHo9y5jT6t9Om1
IHeSMZScwfOg0a0H+27KTVl424WxkBPsofO9QKnT60SlYOqD2V93g0BPUi+Xwtf3
JEZguEQOon8VpJHWXT65jkWaa+H17pBtErcBC6xGfXAXqQtu1sDpKQtvNsAzMdPK
OifUhOSzeUn4KB0+EZbDBrT1OAlfBF7BLrCuSyMrtOk7+m9s2YkDGRU4cGYZki23
QJlYm8RUJH3IEsgX+AXin48diCokrHDaEbV5uREEqPylQQxAhTfO62igN4bnLCOt
JxdWEn6htj9e+JF6cWUvMY2zbu7q85gAkE62RKTxu/5ezYpmj3ocbopzKKVQoecz
4bUaximoZzupGrRp/lRuSYoUFu56twXzKkiyP6QP2XLPgD46QB3kOHAhMGbRmRN6
JC0pOprpGKL58M10SJ3QvneCbBlDY0dvRvntICSUd81UN0Tj8vxVtJONV5Ppo1pW
rFmRx1g05Z8yc2j8QGEsv+2wCbB8DEIrPW3ueDQY4CRd1HQMQ8Bw/FShA7kOeOZV
yyWkluBxbj5iyp+MuJqrRlRL3HG1aSukrn7+1tbnfDHz3nvm4/bq/4H6qBPvE7a5
i+NVimRy4tPik5mmtpNd6KEgQuca9ORCwk2934oxSRTzYZex/2UVYX2/38Tn6aO6
vioMxofuQa+KKFlt8+MgE/6IJSArjGV4ceFGtZVl4DViE974PI31X4k4I2Mlwhyn
FsWkWLExctueea+AsK43hw==
`protect END_PROTECTED
