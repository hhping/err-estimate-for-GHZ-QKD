`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K73ZoILhEZHlqbKFMMnKoGpDwrGD/D4jJdO08yA5D/HXGEb6td3U7Bq1WhPX/shH
c5ccas9+baxyJWd1uZeoawBMRN2N3z4+j2mTNQ737pLet47Ckudh90w9IXMzaCuq
1RGaUI4Pb7AVEPDsXni0Ck9KC5P4c/5Bf6qw0ugYsAMJzCa1F/zPvPtAwgVdP9Kz
9TpWsmKixFG9QisMb5cSLnyHRRRpLhutIkSxHIGYz9CnuHUYm5H6qBk2Y7Qu5Wn3
8+zNTed175SAcR+hSKHDucEqSdzTGU4UqGbN3J64XDdhRzpxARJwCWnkQgn5SGia
EzyE8sN+z99y7adwKEuBKT8MnohqV1oMY7KACX3Q8cnS/gMHjAfeM1lfaprXzG0p
bs2BQ/3n7/ZffLApQfekyK/6xSUxLXlzP8sswssvKPT+yc0wXQthrEfplQ3PMLrm
kDPIvO8FxWg7/vq699Wl/orbpbOvoixPPFOxqlgEq4xlLcqJu4UVCrnfxBnbQZHD
gvO1Zif1LF04OSc5ppDeu53gfre2OzhNxbUtT5B6vYSMM8miXUZ8Z1fEya6wL4ph
aCjtLUKxYBSAQ28JCYyJ6IhUC73hkiBgjtfC8qslVK22+CX3IvrldflTt+6CMrQL
ONJDVkDSP+Tr0RoY2sQVE2e63ePugttpMJ0HsUJRAB7boT5E3TEHJwZqwMyjy8mU
PrEu2weMlPzd35IWJeM5gj6HW2ZXrwXaE936Rx7Aly0HUkAtrnCsLmTXmaWml8HU
Bj98K29R1WRDyMq/fGna9dXOJiIoUh2xlbcjcYQHx7X2h7VbJFEeGP8EU9OSm/uo
44WEYBN8Es8v46QpJTtaB3d2u4jD54akdnwrh+TLz+byIN1ifhZd/x7eL+/Fn9Kn
96AIMVTmkrxTZwtfproOhwbj9JRirnyUFB8Njw1iuAXwUzYjdCRkf7tXQw9XhJ+z
1WmrMKdKVuePX/BD3va2ln0WHbfRGTJsyM9jxc159cBb9XYNqHJemzPW+j13bvaS
iXNqe/nGeVISXWS4v7EwU7nHPSuWlnpRW0jtzGtBBCsn2vt9mQ0YoDx0ox1CucYh
J0mcCZx5/kQwyRoc2LuQId2/kIu9He5QlffNHIxiUY4n7+GjYRyl7ZUnpN8fh0ZN
hNkGV6yQNvurQ5ZPdm+UKkbYFulemnO9L3kokW+i8hTNFQjkPPW3NBkFa9I2TIS6
vXMDt6cTvJQI6JyE4tEkGs9pjZi6V7YBBWP5x3klrmVQYfMZwDhfyehNtqz2/crV
tQuJvZdKLQ8YIxXCzBsXUNjzWBRUlJCQlj+Wfb0dz6j9V09t0ChnwCU4RDcQ5uHS
WGbAGvBTNgmm71nM7ad/F/qEN8AewBDgJ7NZ5suoXAEtmJR86VHbt9dhvmr9S6OT
ZBhZZ5T1oIjqvm0IxFy6dG4moS2r+6ScSlxtmCwwI5emG5Bo/U0GEjgBb8mJEXYw
ShJ/z2lfyUmU6PhQgHoYAi0l1BCoYMR97YO+RZaLw7BCT8o3c6FeaNDyLSqQiPC5
5uAd9tjedHkC9Bo9JE4Ybj020A2ajO0nZL8k1pQCxb+XoDdH051lYqfKq3r1n7CH
L7FpNP1wMSdLNN8BsXQqgpc/UZgqdVXxNc1GbpYjmHV99gM+3QADIORn8mEJpGDm
4R5VzguO19FOoe9S6FSlHMwjoVO0Qj3R6U8N+VHmTltUQSYcyYrplnZyEOETneDq
OBMSAqehjwqO7KbD9UrZ4842nj1BINfREb5yMgGlc4THiC/1p8nuhE/Rpvn7apoL
y0vi+4QGPKbCdtcAxk4IpfRi1lHMDRcTZ9XZ5gE6tzSmulpB8DUwHXhmxt3S8LDS
YdpQdB3Q3AbKiTv9+tYYyNoqrGieHSrRc8cAtZ6F1nOSsXdg7orqcpioAOi7vI7W
+8ECwo16mRRPdIxmDzXhCNHW04L2oNuC95/aJJk4nCUtbDB6+BuRGyt5x2mpxO3E
TWCdhSksNWcngHokT4aeou0axF0Rv8lzZmPKrq3LH/4z8++ADmZhwlG67DB+j5IX
aixy65kx3qY6ZFVCms9l4OaeB/xOHGXLrLIsBdSFH4PDVb/f0AxBI4eK3cVxU8qf
M0pRDAK3hA1vGuRhcjXPcDIw/O5m3OFRcKj8edjYFC1Jgw5gx+icsRW4jCywdM6D
Pavf3kbT9PvmE/JdOqZy8HEL+bDVqUaHWByREH4/AmLB/MA3qvYNu7s+3MSyyLg/
3GORzCpCP6oWlxKaeB2nIjVsBs82LzKHFR5pEjMK9gLWuYvwouVlZ4RAsUC0So7g
l2vicD6VWxoMtkFHTcWiE1hkkBmEBa1mKcuSD5YnrNJhHOaYzAeFEKwS1qDAUVfY
0ZP6vzw6y2nDTnLf9IYbJ5mnRY5YLDzh8qvjwWpedlwCRxSUZp4Xv3k11RX8X6dz
TnQh2qz3KavUDqBD4bl989n3E/cdZB3ooh05UvZQNMSpE60t+ASdPhXnx0pxk88C
ctRbkKgVM8XbN3agcpxg6pFjZanKGiuHt6S/lJqfbJ30I0DtQhSM/8WwDMNhEq5u
q+cWTT3TIPYENEtrD5u16Yy7cZbPnX/d7Lyg4OZyTAQyhtqMGgUHoj0xNa+OaiNc
kt6MJzJOEHDOAIbnnBPcV/hEFdbWv7s0oIJstF+UrADb3FRTItM1D6W1aSfhNWYe
/Ok5SL6mAHiVXnT64anOavjIpWe2M9TGoPw4rzcyJLtL9SmnqzOrXllKrHtlG6tJ
eG5sXBFIr7LjuvSgzl7RLGHH3yVCJnHcb9eVwiVEwOPGI59Qrd30evg3y3IZyPlI
HN/FEt0FmQ/EuHxX43Ik6nBMzzh+RBWJmhSwCvdvb9MPzZv65RjYHEsq+bBvxHpd
KUQQ285IieJn7V9kXS6AyDAkuF9v9O571WLYdcTBdH4O7xd8DI/6Vn04t/RA9wb6
SIa+44dclN+mNydcWQ06E2tlr29x4h/mY0WwLmwlPnHaNBFj2C8oUg8jPidtuGUP
AdyYarYKIrFUWLOO+6gIp5K5A+K/PMWTCYA1eRdL0Bg0e6HikLwHnaEyhTT6lRiQ
8UyvsqKQFlykhMVnEUwesLpYd9TYyQharXoZ5kScWOh/v8cGvUpV7UhwqcfyKOz7
PjXM+rv9kpz+LXxqIMdG2G5GsBrmLdfOK9muSFp8VUc1/7lfmQ/IMO/SSSE8hl/K
Qj98zpyYslMALpMjS3g9dzArfrBe8ZFBLHmrabr24ALpgGSCSjD5GiDVNI3/3ABT
+MDMOXJpybBHZP3oiA3I94x0o+AwpLYbwiDKVfObQG7103fMYBzZLKAxuNIbDSDO
Ztk0g2BesR46Rgpkk2II6zFj5Vi12zUuUhVHlqitSy+Bib9oI436zjAnRxFU81Yh
EIch4FIG6Kcy2y6w/llwhU2L9cpG4gjmXqmc8j2TqN8+WKYoHM9dQvdX8zJ/8qs7
xdKTZ90hB5vgcBX+7XNxsTzeejx5JENmVk+Wfwz2PbUvqfIGF3I0pRIll/CLo+rq
y56mFTlhOejaQB3KZQuZlan7791+XAbO5S29saTxzvTmZNVtIYdM9o65w1pp4YbM
Vz2uwB4gnXqc/LRZK26BpaKYv+uiqQkTAXaNvgpHiC+V2BJk0PGLyrMLRBk+FwiG
Jq34uo0+kcStH5+OHckGMSvV0Uxvj2Ar2H4rVxSy3v9iuX0Sy6mJIXQFpWfWdBKE
JWosttfoR9IM43Q/TgblyoehwcjPqr4GPKubtKRBtcKzFsid59UVV3XI87CQdpEw
PFGDLQbHXZp78hmanudxjVYloT0J4Hk5wv8mM+8k/dzNbD7xPhyZs8/RxQ878xKq
H8jvA7tBzkYlA66shYAF1fFzznwwzuAELr9Np8zkCq3J1X37aJ5Kcc+s7y9Txpjj
gKQyrJH/o8bEcJ0zK9ZKXglfzdpkM80hsqMRFfKpDJbdytG1JPV/+hzNNuFpCihE
q3Mq7dcAErP9KdEDPvtaj3r20c2Lhbi4lH+OwyGAwfKIo4VxvSgZmzgbfgSPNebA
Kkv6Jzq51KP0HK1aQSeelpmCcnvyeaOHhazJEFsMf2smkLIG6ofcjXpXI2T4YYL6
CdPxDijaIvb4JGWFatmNOSQKEIEsY9COu6z/+VDOuoStvJpVAFDXiP70C3Yg2Lw5
rCQ7Iq1IvnZg5OznXWzvDtMli+nQpZQWNcdy40lCbML2mH0W186X6sWvj2jJY8VA
rXqeGaL1ovx40hQTtKLATUdLba/s6QXCrWDQXp4f11KKeuB1EUONiucVYYHVtNo+
9VyoX9sR+886qPxw7FR0t8wOJ+aeUVWPCGodCDxZpzNqPGuSWXS8fP7ecmTaBKfz
VIkzO7bjqXCoVFZRH6HkPoJKJoIDvj44rSqAXvlsKFLg0lZT2Z2vKGonKpCkgB6Y
BSjEOOOZIIe0kcpGIpknreVYSOyRaKMrZCTa0N5HuXb3JN2Gp2ptVshswHGKod0v
HBxq4hcx6MunQxd+bsAG04RXMtTIIh/XR+/e8di8BY0A6VAECiNyiffo5dQeaGnq
PW3nl+IlJUgs52YKnKJqO8WSfiM1O948ykoIExy7ZvY9PbgDe64DdcM73gZiFnnj
2EjC20nzQpq8mL/48pBcJeN5Z1ArPwQglqEl+qLhP1+PQ1lLyZv8qMJv6OzSeKrO
NngxXKZHmHBu5YlA9WXohTo5ALdTjo0EZUn8bBZPgDTwOLhTfW9FdKw+vne/Yx72
RGFziqz8WJnbZYFTplufnqonoPYBy/xGGMbhS4HMVvMHH8iYJU6aUlAVXDpRa5w2
0tJLcKsPfMfMJsAx7ka3S404PPmSy/qJjYAJe1UElYoC69vVBb6JGOs6rc5slChO
tADuYzWr3A6hwk7XwGE3lvSzvqj2QfpDt9dnNow1IPuP+EezWvyl4X72alo8T6x/
f8hq6tonGdbRuOXZHUW+qphDz5SmiAATfY7bU+Eyv3pY2eQHTl+GL19qXBJ6RhNZ
wwTC0AKFZV2d6YJ49fOzTXNG7BjQ2Ra0+4BNnyuRi0K7C3pGSFqdzUMwwT/OWewa
oItT9PEnKg1dTrxNz3QCykxpZk4dt2OTngC5zTPYuZ60R8/pvsvtvlSCr2+IfzUM
rllq02bLs+KEyKWrE/zuBMSfM7rn8g8jGcBQwfOxvZ+2CTyQuXYAlJzArRq0Z8TM
eQlHvsorVnMwImHZytST7Fghpq1uI7OBclKztXN2EykZJNY7XkeV5XzaMVuJN4Q3
UJ6PbOE87br3Kpf/MBF2OcbK/+ACdKTwNnwZh4AN40cCwWqjivbG4/hfqgSfvRFt
8Tr0LM37nL3laMKjuZY5m7pggBHnHnNPZ8E5JOBkQW1hP/oAt+IO/kyLmiXU5isa
Z5s/TAehTB7dFE1/sUmFcQf13RHCFHtA5z/gFfw/BvnrVEDjrxzDE2zNK2dld+3x
GV7FVUTTQBI/1hI5a1N8XOXMwf3sNuFwxg8HNfUMLtrZkGVgJA4Z3bAhXMrAsO4j
KKYZjhieMrFyMyVD6zjptmx1DjF2IfOe0b8tHJ2ZaFxw1Ay2KwJVbqluhOkqqq+e
p/lWS5xR5NaieoQAx2giZc8fOBcVmFz99+UdezLr2xsJdjwCBfczrDm4BVYA/x1/
XwSdS4OoZkslIwm/XCSu4u0+FWHSuUP6tfLFu5kCuaAZoXjMQySs01Pz4FzNv8CL
PbLHAAmjoL1JI+ljJeuGDIQ3rxSdDt4aAQy4GhuWeIhbozoEFWSclc+/EdiGJQv6
MVOS58uPKgegFGxDo0o/8G7g9l5omHUWpF7JifHit2IaIjpELRjJsg4VEX8W7BN/
Swo6capA8hG1FnNxrWTU2CP/mQlfGTYmSCEwHHStcDQqJ2GhsZ07gmJaf9bVsYa2
NHU52hIIx6n8RLm55Hre3LT7jXBqI1jim+TE4yG1RSMgdifzteTzfxAdCYL14zGN
eX+40qCLGa6lYZMuoZill4CTOnlMUYkJAzxL3p8wDacGXX3iVjVUKBdXz791MiJ5
KbzTIzdAnEsHfRvaHepudvFnzXjqglC2UMwz7rLbunX3Xicd2gi+7wLSsUv3+Rpk
QRSvlJ3aVPC4qVy/txGbcy16IlvgC4iX+yd168Pz6wTsr058C/dv7HoEvlQEu543
pUHnN/MTJkD1wcW073pFBDYbrZrcYfyg7/jVVvoq/fEIiZz/gyCZU5HcgHwor4pg
eKdD52crR7ZjWBp3eUZKKhQwG8a5EPqQVzHeYz0Q6djCd1XIzHpbBos7Cpx+rKSM
YyZmoKbt8tYRYlQRt52JbA9yY+Cl+naIRRA5H0Dd0eTn19E0f1LXlkDRsjQtO5q7
F278XJGj0sFVv70rwUH6PWdvVABhA5Bdpim6OrOQCFIaTTrRjbTyHIJjvNhqXcV+
1HhklwvOr+4vSLlE8KXKTMxNxhczjwpKTJ7LOhtNDzCOP5rkLOr/J/KyT2OAoaMI
EFXZBTrHwpIUkf9VGWys3YSnnJi/ee2AW2zNCsTkmn2nEQvrz9U+LL4FQYAh9Ghw
MV4j4HbIlYxjyxr6Y+HRvap3E6jdPnDF1QmkYf2CGs7G8x7Zey79hfqoQ1GmFXbZ
39etpuEJ8xVko+Xc79T+5K2moD4WzU5woOKM2AF9w7VXmCReRRMHK22IpJA15Coy
r5kdizWTaY7CYmy1HnBiYQxIpUN4a/ypsdVwmk2/04wrRQFqipsxCIu7brcAFMyf
yLmzKEsSh00r1AaYtDjdTjCnj71bv4FiqDmQQWxqnWgsbx9iDMxjpKtwAEp6NNd0
Eh0yzs/DF15NwFNlDjdrOlt2CQagCUsI6SvPwSkU0F/qV/fUwxd67Kran7rQ6F1z
RWUWq5/l/G9x9jhPfLNzsvlCgGry98MCWQ2Oe2rAxM/sn7lXFlhPpWTKjAxFxggD
9bKyHqq45DNnRlSjUTrE5rQfoyUsVzXD9EtPgRwZoYPIE43Jhc41T1MbzQj1mGRW
IXZqEIGKVFXDrQNcRV6FAziZrSlg1ASbvXIQnXbQcGWQR4G16pBpZRto32icTpCl
mIRiKs9YxICj2M2qjh0oyz8vt6RC8Z34I+gyCdHxSrLpo+lsyxeCprdeIgGIl4SI
ynKVHMyBzgxjLHPXMrzVDZaJIBWnx6Bos+SVsEyMevnUKyV2M4CQqbeV72WYYOBf
8vL2O1hUzAg+WoeA8IGYARmAXJECFX+oSZ6n9h/WXGPGmetd9wIPChQqLhXmaNM5
TCiHGOZrZM9PP7KZVFHGNwHnfgBfyQxPvINYOgmP/RplFYOax0F6ftiJRTn8jzzA
PGnQbWTOpY0SYkEfMzeJV4NnqbpmPUjhNVj8NcfsLUO6/3CFW00BHGnkAVHTUr0L
AcfLuz2oLRRH5sNccRNntyip1CgyEAB7VVH1Kedv86KLXHebPYK3CqYpA8yMJoDx
SRPJsneY3b4qqCiJ5a2fvuAOxEhvwjUlc2Cj0VBJsTIuY2Vp091D51BanHnayUQg
zcR9hfCtjFtxRNZgXajlGRsvRTyWYixbTUPxwjccOct67expfFqOx2SNRlbFn+xs
cDdeGCJp8CX0x6bfvi3mOuyBxR1FWZqVB944amp4oJg3EpTVjt2ZQy2VrQUVyMhO
V0hxsYpUlwUW9twqIq9zJu2h2l075J/owdhp1I585XZQScoQyh9ZFaDI8gOmxVQ5
GHfza+f+9puJ3vqFXS1mNl/m4Dia1nEqPTmap5AAojh177MccY2zPz1n6vqdgN7w
ClF/OllpXK01+TiZPNi02RWOsn9VE9FnWgBlXNKX0kOLJGok3lwuvGNqqySHocRy
djeeRK7htZx9Vkc47MSiDQLJenekMOIrUUtUoVW3BaTHBCl0dh8YRO41s9IWK/kn
ltWOox8bn6Ho4cCVPM513QfQn6JMIPZ3xha3xoCNE0C9m+8ch2HLMI/h3GjftNKa
MVvixcaZeF0+2TB3r3QuropIeffh57TIieeNC7PDJXhdxGXM8VnZOp/GNx2xN7kI
ghu+hPbnRIeSPbzii8+6s5YDiatbZyaaBY3/sOuttjGVFuFE8abJcBesjS/u5yCa
ELaA6BQmeToKQ/4m8qnSaQ8bikDOUDvZqP2SLFeoBEaolPmH60EnuUjo+4asrGWL
iWCNPKSnbgXokpK2UrZMhNp9SBYKLwtYs3xMV7gZ4AeTFui41bgHkTnGqNuyGn79
9ev2ar03Ph9LEQyRpO0oVyJqvYdLNjiqg6FNtSyuotQP05IV4/BnNlV/tjXDMC5Z
HYxmncjNBvm6mJDGyLALzQQWnFP4sMVV07aFB/Uek2QdkBhip4p4T7JUcVUGuAD+
O0JtJ3VxCCPcDog0DXXcKE/7B+sYEmPM8h2oILsZB7Au5JcFoiboUG2MkxAJbdXW
SWccQyrMpR34J0lHQxG+x0KMaAUXZWW0sfDWhbm2vY6uoZcGS4qET55orhF4CIKP
+UvzSWCWX8JOCpVP83RwMyAsiQ7lJa0CI21Bz0sV4HOYgbtFrTeJC061pmXmn1rq
liXOvV9bbLRIrCX/W98c3fGZHYzubS0joVbTOKJPI/oqYC1qUK7C5n6BduXwt7wV
YKr6YTUENA/cNtynpz9tqYItML+ugxbRkBAJBx0mHc6f1aKxtXDrgs5b2/AkZX6r
6CCJ5SvZjZuQF+I339c/+7zZ0YUCPfQFKljblfFsni+WjP8/YjgeAB1i6/iGKYrX
zYEf4Gm63O8y616TffYqBEQ7SJ1EYvb1MtQJ+bEpRZzZtSEhSI48OnGoOXQ8yGkO
1/94BLyiMYGLx3ZNqVeQI6EYA7CsvsdMCDwZAmRD+JcpYRPqQj8RiXADXTG6cx3P
MG+lZMsnwKXNgBh7qtCmJpCwiTCun33Kkt5ixGqCqp9PHOq/GP7GBNe4CNYEIfE+
/vqbUoyKJB1JoL/PUlshyGmIkNyzsD0wsoxNkwXEJGCuA97vbnpfyvFv5S3jPyG7
ZZ3HPxtGiJm/5t829yq6HpUQr4TOTVkz24U1rBaCfF2Niq6uHT8pJhEUf/TFygmd
/c0y/JWNbL+NmacGGV9a0Mqgrud00jyBrrfmNjCb/JIQ9agd6OxGKiVU9iskjrZr
BbetGXi+uDRxvDM38r//mmZahrc00O3wu9fBujgGcRJEjZxX6u/gJ64vYYKi3SxC
wc6/oAzMYuh87EEqhN7z0/FEsCj0E5P28N6bdJbT+VmRjQZcq0Yk6FeLOP3+fzt7
Jfo/rzDYVawohGwVII3ytIkhzZYZOf/HXAp/PoGYTjZeuwioiVdsFrWZCocTXd+O
Kg+nZOu0A76zZXKvydsY8ROQ+vuSdlUX205QqCSYQSWQCMLGTij4Hb1BsII7k08w
gPE7Tg0e0R1Nl4EuqcxZkOiYRdBR3cub3fE0fFZjM5QLYYNwrG7qAhF2QyPyNgQg
USRo0sx9lno3Lmc83i8opGdPEh3SZd5GMWUb/rOT1QTo/R0xK++aj9+flDkVoYgX
cRMyCKfuVuFpBmkKc0PO1tHbb2MGuU57WAXgUhoBsIsXzt9g4x/kbx/YjlubKgUN
EwYQV+Hy5c611cw5fPpdkaQP03Sywt3j7NXSGmKGerfoc6w63auZvIOPDJZk4p1P
CYfsSN5tiqj99z73YWRqmX4pVLBo5BjvN+6rnnp52kTtyGaBqiC6Z8kqBlRY1S5L
itobRoxpAd5uyc1In5/Eax90WtZ2B5rujexaaZAqAvsHozesvOxoi2ieLYTZa02g
wwxogpYkQjGOM5maB52MSTTfR0rJmpcVVpCL9NhI/S1kcyVFw49ohqc/iLlnzRTI
N9GE9iF+j8BYUoSdpwDuGTXaFNJ4B7g2OE1Bf9P4IkFWrioZENqSPtfC0htwJ7HJ
ZQYWxYGe0CScrrXNK/ZiiLGyOg/l1XNcLpcvAUmZs2NNga5ThOP967IJugZyJaEB
2UyEYgz229FBHiOHPBlRDWu05jTNfWpOPxXquuOywTDl4GuWnsMs2RsMrKDkLNNy
jCyShQ2yNxJvaYXyHl9GRTMRpOGIEdYB42DvQlUYj1SACsTSC3MM1kB1JsAK5wWE
nIRH+q8UnY49LSqfOUrRXI7oSIRSSFOsxfxFzldSaqmYEP3mbdFzl6CA6urjCJ8R
MzAwI3GYzBrmlHxKx0AkAyXB12MO95DE4Otzq1nIN7mqWMdYNf3whe23RRMr+smQ
yEj6Gzm/vP6TnUDy2jMS63q2Zn7HP/Qy/M04dyGgbEGwm/OUfa08h1UN1CdyISsk
c4eSSv0oU8smje6b3K0Zp/VCkhHkGXP/8Drk6vH5OUjipkxzsD/FBlTkZk+aRmA9
+vH4VSkJVKUu4EIb7akcoJmRQ39zdbfFFNQ/TX7Hj1aejMqsVPVXztNLFMfKqXRQ
zneXrze46j4Ib10pgitqrUyo4RjDQ+gOG1tdBmmZVGw8CttnfrcEAKdOAQrODEwa
xqVhUwskUMFGCFB1LxIlR8phs4uwC4DyqXqdjslApRvnodm3tRdPasUeduaSQpWr
wvagtdVTzZLr3WQMEeiiWc0N7X+mA0A/lnkecmjhaNyIAdDWR4zduXKhrP2JGbRX
XmBpQKsBbGZZnNHj7rj2OWDCt8UaJAdq+32XauKiDi07lmcuXsDPyP+kxrind7eh
VTGyq0Mpbm+z1goFH0eZXdsnkTbyiTPCyLZV6hmnASFrHGt6wlIbC4crUxMX6sxu
SFvggums1VRpDEJFsKpm4RRItAns15OdFx/W5+kTYPtbtTBXDRHUKj+nLn6tnJ9V
26aV/373p0w41DbNGwSecGQVT0OfuVdExpy6ejnteL5g6J5tj72ztNQaCMymbi9q
RqRwMjoyxCYIPRK8zaXwEIQwVdpANkHSeo6ulvkxHDG+dfwLI04fc/Rmu67i8TuR
KV1UF10KvuDKAZ+LIFwTXIL/UYN9m4h1oSg09Cnwp9pVUac3+h2YEWVmG83TiUCk
lRkyLXQtscyn7f9AQAqhQCISs/s1eEb9Wtod6v0pPY/dUvFjcOe9eMTgE9uJPiN8
0cxhSJJXqIkoAze+Kt/31009YRmGJ4OOnI+soB0aj5G342tLOuj4yqpZutrplF5F
WzzP7nwLEvMTKUbfjEgsRkOM4glCvXid1b2yz0CvBWMTXcBqSuXI62ARWu2KJZiO
hC2V1ds1QR61UfMAXxjx3aYkLiVMIGVJZOUNSNv4OsJ3pouyjOd0p+8BOLdXtHg8
Y77xz39Yzh6pVrRoZVj53L7hWym7F+X22Ody7f1ZUv97U4yk02riK7fJ1kXjD/DV
zw6/kWVxBCHFV6lAmLecUyQ4DkNxpfZUn/73mOzP8SbfSizgDhGjEsRMq3Dq3q+n
/zUQqK73UZFaOazk65xhqUF1fV2iA/jO9Z67fM6/U7TrxRqbEkhIWmRKARceMrlT
OGVpNR2dK4Ypu49jsbDddxBCMX0au0jAhQWyfPXjUWy6RDleIOAyficxeiBKwF9N
E7PLrh6/+GgYPY39VaFRS2uUiJmsCcex/k7pvV7FpApPhjL5zXdJN9C/h9FG0U2x
3NHomopp07nK97zv4og/fKoQHtoHVuIKncEQ9t2DprU0BMZpzoFgjU8oortwKj4I
9oAN9XgnThGD7AS7IkoJrEAnUPGsgKJbGop9VnrUoDKHvXqh9vdiZ5maq1QBGNYt
wKyCox2DKOHHUPFZsRpkp99C92ag9pqJu6YA+GCzGjf5O6114bmXC8UZM5K+cwV5
J9vbQuAG24lBULoC7qpDWi4jJ8kRGqybkjBHYFVZofJHThuABlTlK9oWtlAZqh19
8S0X6wxHgzguRziYHZs98JtdUbYWjl1ygAHy3XJA+eaaHFm0VmdFUyPIJzDk95/1
6SU+kFnCkSU+F0uIyhlRXQx3+6wVMn5Ze6mw3m276XFj3YKlsgvkwQM1/XjEekjK
K9/mZ1fmheojYP3SGfCIHCXROiCrr6ztwJbz6in67efEpjdbtFcbflpABMKhz+x3
qnPRex0CucsbPDCPwqA+EU+tD9auxoPc4+DPrNRuWbdRCw+n1aL1ItH4BWvldjTZ
Wwa97dLuGfggdU4ld40Gqj1Aj/PzCWeBqDcQKE4XOuBG18XTWBJGkksQnQpH4Lef
Pk4opm6jO3+RBXHWtck5ZfqlemSDQoa7j2dKresin1gSuRoS2Rr/B6gjL0lKFpkc
x2z4k2RMRhDnM6p0wxoW7Yp7v3luUlCfkMAJJUnGdzrF4o+BYrC3eIt2ItJN32i8
tyPTchZFsyrHS0EThvgvBYhaTSs+qu2LjcIRxHYBe1JoQGlXy45xRAbZqH+KDXEv
Z91Jky2FiBghSF15eE9v6z3jiQNjepWmH7saxn+gETrJ/x6yWDGdQGYf9VToiFLK
ytC4JqVt11oB9vSoxLXFs2rq3Cidinu66Rr7Ej/I0BLTqoJGm/E7BIdz1wWZY5J1
SIvRownenQyAtgpYT6laIWY76XcnVUb8ATabAyu/MfITuZLm+9rA7dVyreXgCIKY
LBBXJnjcKE84wMw0mEx9ZCtP8vhnFXF8pnGQXAndEMngmevFohiOUM+9Rk/EteFx
nPxc0EjZE20aVuzs/32LAHfpnZ05dGInembMc2ZN8j/Ic3jz4W6JRy5s/lYcFK7P
xncSwWyMMRf3goJ79LkCpJqJnySGKi6hbFGS4LOsdIuWKQ+iMhvzHRAfzJu7SAaq
e7y8yzYO0QIZpC2fV94KpwPFtBjK6/qOtaij4zN8BRHYDKrS0f5mVlmly2c6wxfL
DIfJrZiXAgvYK7gujjVfYO5prGuCfTT9DC21MvvJDbmqDcdbG9Ai1b246DiuMYD0
5ifLS4p4ngGO6lsHvmlN2a9P+dTQTX/0JpQM4xLiOr88exRIZbL0lKtdHlLjWHn0
yGf7BJJtBstVcJcHdmwYc7L0eD+G7x0xxhQS6+4zzJQk2sMnDVtSJLAxRuSOa8FS
3HB6yIWusA5ZYGjCVLEM4dtA0I/rIE7HxXvx+DkkjRGPXL1XBWeeoLkvlYovElNU
g+CsNqeZb75j7lETicpWLn4iKRrAvPjWbP4GdBPQwcoEZM5/Or+llwNSGeRBMXmC
U4JoSgIOeFlskPDHsA0XHqxcXmpNqCupCYiyWBLLLJdhpa9p6jg9jbkR2LgUjh+7
/pVQsJN0m3TfxeO/bTRqQ71wzp+HqB8kPyNYlsOqaMB1gZjCK0ynFMtMtPXcKWRZ
j3zxx+AESw8K2Xx55aXs0IJRKOExFm9N4Et41EtI449T2/7zX5xUa210o5yG92Mt
mYJpqSxg9oaHu8V7zz26KGhQLiWfBPQos4xQi3yoW52ZU1gYdhLbCTRveIXbsi0S
pD+/f3F5OAinM3FK80tAdBpaU+9uSPNKOtHVIUohejVvgub17NSLDhs9wZ3a0stT
0Ywq3+Had/ZZq59mwHBEKtJO2iygLElV99SuDiv2EzuZTwSk/qHsxbF/9xrfLq+7
5LgiEdvf0YKFhFH1siz4wEK3L1MT0IVKdWoyQATnnid6ZAgq1TW8ksYXZyiFSrgx
zezJvoBYiaXZ4JUGOmuNT5WsV9lQggo3PFotjJGtWzUl/0zcRP/Xy7uDbXR8YhLJ
NKjOUCt3JtQCUSM5DUWpfZ1BhWPeOf/6dwNLb8PsY3q/h0Jgz5ElgG3lfEviXbJ7
lIYRC8ECQMS/3z8vZHywqEKOI0MKEw2VClgqO6oE/RbnVXkjGX2ZjQCTZZsCPR4x
Uv52XVuNq/GH9T+mJdSH8bqjSMM1QBjc5n5Yu/9P4uC63orxHX08TXSe4RAPqutt
zVfpysuBsFTXhiYFDsmJppd0UGof9LlY6xn6DhniZnYh6c0n89D8KlEB9wAbrcqU
DlyrU2yrUmMzYRcogz5TUA+fBPukUe+EJ3guHmUC+uLi+JTzq/HjEpevg/7/TpeG
JzMyqGE46UUhIcyW9QX19yG2kogLn7bW13hS70KTAITS4zK7qOPaVkMw4EVhZY+d
ttX0PImb58oMc6twFQxu4yvoBJK3GycYYjFnUWmRCGoG6ViPbDWTtEcXxxhHv04i
nJIte869Wbk9urgAKuYPCUeWlSeRKErlYMPHIxG7v6i2R9MJa/F2tUlFq8FjYBrI
dRkcZ33/+CYOhs8TgJriKl7m6VhFoAyYETPPpB6XLgEHw9G1AUGGS3XLlzpXh2iA
K9Ed/Dnh5dBcK83kdLUqpe9b3i/rVl4QinuU5DBqYwNYXF9IGkc01sdo2YqqfDre
ilotrIRvQkxJFjgcN52ROfs2/hW5JqKq3vNtyZt1jWGyuTBDJVFqdGWJY/niQxdt
LWeo+WH1mCW4txmad1mtzugmjZFALcAFf2cwlLo+w5aiG4cJtnmPM3wc9sOWbO0a
uYD7JayP1vvoJYk8By9If2mpYEPdiAAfsu5/PFV4/nDYpbOdfUAom12ryijz4brh
EWewusE96Gdjs8f6wb0CR4JmAnk6VCD3xvJRWMtm/iZLI58HRVrZu2BfwUmZLt4q
5F6cdqR4K4O/bkRkcohWYGHiSFNXLty+hs+X5CgZlUp61jrq7/zjkCNm9bQdRIj+
a60Bg75kR2DK0+DCyrxNuBbmFf7zL8p724Eb0P8XlQww5pzgSzONjwnvwGE5cVwg
dzQ5AZzKoFEFmzA++iivWnhZftZG36H+n6gn2xRBQqGPilLwJAAkoQcP3CCyljUP
ZyZLIhD5t6B62zGPncLLr8lKpBpYvdMD3AE5jHjBI63aI0VlZG5dtD0O9Ma8i64J
M6gnRUCjGEx2RK0r5jclYWR4BniYYXwsovZX4iIRQyQBckZeNw99X6vgLSRn5op3
5n7gK7Gni+cHgViglZodEz/cL5R3zW5uC37iYd248fAUiYJUs3ysByH3S/GPnyS0
8O3sA+b/t+mCWDH9e7JqxhuykCmZNMkrHj1olI2emswhFasNqWt0BF4AGhZGbFR8
UQx8/3VK+G0wSbdjiCvhO9/B4uVRPFO+312tGz8qdPXaeMiz7qHChNALsOHYmLnn
U2aHHW06f+zxb0kemcq4SgK1EqzAvYMtCcR22VCGedDXRgf6POlaU0ENowOnEvvA
iXoTxvX4YNd7TAOnYH0jucnu3YlaeV3gFvtjZN9XvH9vpw/WxYYsfql7pDvNZtA6
I9lzX+ZDqx6ZnnV5i3MjiCnzn8J5Z9PdLgzrxvzGmfDN+aJp7zrxFV7X715mS6qg
grVLUOZMMBCGJzV7xREBLmg4x6YqM5E+n71zfJItDdWprmYQfSIxXULp5gLgzP2s
yB0+jfpfZ9YqQPODkSiBGaY5U1Yu0Ho4gArq+sLos6noflPrfLfpXfxeAKhJjULK
ZiCd+PjTdY7ccszpCTvbNOMfbLqGzgWXyd/J+10oE1oCdFFEF7inG4l2X6SI8Ehr
qpBuQQgU7xk79XVxtGnlpllWn/WCDUkn3enC9yBNI2pabTjBhD6t1qN6q8vOCcyx
6R6X0CUQpTmDfFZZUg3BqUtV1QnkbNA0lZdzAD8Rsba9w6Md/GmSjh5X7bDR5cRT
BytWIl+Qzed8bK2kEStdq+Fx5YXA3K0uSj+jmwlONDgML2aUCXFYtnPEtQF9DOqi
P7j9IfxHHOokJK9IpoetsPU7s4mjE2BUKzDA86TP+i6k6gFpnzfBwgne58Ef6Xd/
E77HaUYJYlBw4ghlnt+LEhu5uz3KQt832MkfvW+sOkhPB3RVbD2HsIW7Wlg9agsQ
Z7VQhCSpU/wF3F+qCLFbpyG7RDb56TbhDcHxmAg+MQs57pCR4T8BEtLOJ2lsyqdz
w9vaSZV4Lv5XaZ9fgBLljmWo+FVi6Niv593y8pLHZNOX1vRr8JB84uzyWxigBhCR
6whpOz3F8dx8NTwFc7SA6gSQJ00aWzn9GjxMKqc7eUKmIOtA0UvW4frNWwzHfJ7V
faweDRu9ov54JB1+YL1uyUkj16/sXTeMFC6jzvIac8ECaDP77PAgoMw/ndIRdCrb
4nvgiR1R3UuFC+0qeey3VJCNFN7Z5JyLy/iUBRYX11nr4fdThHCbO2zPWeK5uf4E
ZTqpoRTYImfT+aNJ2MvjTSsfteyMSQK+HFUgJDwtu8alsrFXDBaVs6e+0eiHRppK
qkWdyAyZVjKTeY7xeFm1mRia0RYY9krQ+CGQnFqyTw3tViSO5HxGjn1UaR/UcXiY
M8ffmgrdr0f3IPnLOSK+E1Gu/DVlCZpmX0Uih5G26z5Nx6ne4iM4fOcrBH6A2+qe
AT+43QQA3Clm0it7FgltDpW+H+V21RLYoD9DugCo19mTj8OlBmAk+ju9QrY91guO
OACsVSK7o+9wZRcCzui2WKVlYPq1bG08J5HhTI9/YF4xWNyzmvIsx8yDSPaHCy3B
vTDNGRKcGvxGEBljNl4lJTRH5/3InYaS8Jzj2mRhpMmX3nsJJTYSEM5YsAH0yFvg
2drGR2d0/f5oqn96pFuUkcaChAhxJiDeL7JYhvKDWQx0IIZ3yzxa8/Rtkrc1UDCo
rI7WR9h/GWiTdLrvwTjfU3e3Yo2fSrPRbzXbM2aqgeSiAoyXbpDbTnw1s/TXKDzx
aGowhfUmqWXJS5NyqWJ03OhgNRCoEcz/5nrwolx8eNNka9nNmk3yFPGf/PPd2wfO
I0tPu0gmwkYjjX66y6ePiiKnnViDpi7yGdDWq7QpambphqbYP4NjgqXRodduBF+z
wvShSzybRSghU8R5lLpeIFvK+Bsso347mZ7ggPdchydcyPDqTGalGqI4pdbrOOgR
/0v/8TeqCIXyxb17XUTmvr5+D4m7ulADFMVGdKyAwQlCfivGvgofzE2s8pT+NcjQ
x6MRjWPirUBkKEKekXbPFSaJLf5UZVFGxVZ56mjbHZJcSEOklVmx84KXebLv5lWc
v3vnx18OoohtFGkyx05Fq3lmg4jtd4TpzI6zd8KxypDJcdt8370nRu+dyXrW2q4o
aTlCI43spE2DPx/aRMsddSSdy/UVbEahrHuzI9L71+2RhxSbFJNAjgEEhrvFQCRX
D6WvAgg7SS5o+8qUoBvKJ/euQr3fUt6YhOyQN/g4RbnjEkG+9pcB9EUCiZQS264s
pU8sD50hqD4IoK1C4yGTvUgxiB6TCN9D+zAAc68pKdK//djki48z5nhCfWs+dElV
WFXZfvU47P0o3bCeURIjwYqGHTkHvzUXQHZzEdmVeldw6Cql10qhUJnUuMuldr5e
Bb56AOuvyhEBz0+lZJZb5ruExQU+X4Lh9sx3ksrU5ChBGkVSlN7NEKDvrQg/dc1P
Rsa4D/WJgCoz4WM48QmLgctzNVo0bVxDnzTHrowPpzQ3ltBW/4PVOPfRdtwu4tl1
YPGk3PM9BvJlYyM+JVTva5BHnxVp4x/MAd5NQCw+tciDI7Z9PUXbHH2bmfw5fH9F
/7Dzy1IaPom3d0V0SeXR6AwmS8rSjzLv5saPrNOOn0XTZEYSVhF3C2IPZtlP6RIz
256CnWLEscO0ru/t/AX0cdCgZrexOPMZBqym2POPn1sU/FdDtnBQGZ6YudMotlpc
mYQ2y8bDy3YFTQ7HkwwPeQtcs1pazXyt2iwOmkqNd9JUa3qhqvsV3vVecL9O9Xw+
GdlFS8eqA6iuK6+GAMsJZ4LkRcaRrpLNbR70QV/tJ1jrhANiMDDQsWQJQWkI8X1W
ij8aMmD47AeA4xM0Nma50+sPi58npZ5clQ1xrcSlzPVRcIjq4vHtAli9w6oP6MZu
0U3FGohWpm7ICf9fLX44oJtdsjuTZR9wiWkoUY1R0loVsI7WM2iMztxTneSQFKwP
Y8N0wplWyk/wA2XzewLW4DWgSxkwncnW9fTEufHxnT538QasjCNUVsMs2XsWnmoW
U7Lp149/WVdCJ8o4lBOOL4XEE+Lg/NKNBhkuAlv1iWl83B57P/SWBx4+mVJWWB0P
4brx29JvV9JFhMs9dEwj0bi6PlrsVBicdWALqx+SyOc6FVh19kXs7yuqNJ6PdmYu
l2rFZmWbkYGUw0btjHb55BMcN+RfEO5UJlQGeqJ93BvDFJX4Yz41awkBr+pgpc3B
qLBBK/NhBMPBv1JsqmKe1ChlPgbm0bMz/pGC61UHkTsIlUVjGNGdQxX4S/sqkXQX
2hEW3BVEuyJ6V/ZP9W0GUk8D6Gp4efuQwXLcZ5cMvercSe8BJpAtBvZb3B7ZoC7W
XLTT7pqDinZ0KNOcksb+5oKhWCmPn6W/oxW2divRKDg1KQTtnWC7vIXwQZ1K65Lg
KKInt0uzU00ZVFCxGkyewWad0U4JAElFBk9R1dXM6ee93PiD1QLjWXcThVFRnHjT
FURkYOd7lvvQcPBrWuw4DZMfsrnUYvsakWevGg7+EtRlFmU9HGJRlOs/TOR1Q/ef
irJ6VSGM6tjEZo9iayiAuzyigDio82NXk+NkuOaQ71TmkI1S6goSo1dHTYwyqf5l
zZW7bZy39nLXkeKEoX7g8shHsrJEeYmI7Ts5dUT9pJ/2HbPmCMjXb0RGPFeydRRO
PGOzE2TAB88OfXWJSVfVFhYvZ7Dfitxo3KbiEjURnmmbhc2Be7mMVpSYVSubqycS
Da64LAx83OAx5J0M/MczId0lS/wxNfiuwEh0PThMINonM9r5g4nv8omZlvKB9wro
TJdFB97pJx6i5B5Y7c0vWdVok1xFNOFLGw/reyIXRevH+o2LMIOD5YVh6FEDPWqi
JMCG8D3JZiTWWEucS3K5xD+lIhdLSjUnOp16twvlTdeCFegMNzwL0fuv9KUTOpkp
YXfKbaB2WpxK3s8FiYUb5hVwQSUDcSnVXg7v4tDjvqD3JcTLXTwwEsl2MHbKT46R
+VzZ0TSLmu1nSFXDMtNd1AyCFd0XhNvzik98rAb2H3FaHNgrjbTDSYPl/bgojaEI
NKlCKZ/rP0qXanuNCF0Kvs5VrYm6IQn/ULqe+E4XHonOYdfWx6Hl2Y//KtzCAL05
F75Ujb05EpdUoNzss6TEl3hPfDocIs/CJ017AVqQJxUtO3Oh6VImzK2fHFmeM7lI
e56jbOHj2XoANWal2uLeX+sDdCCI8zv36r10YTDlIcdsDgQ2ilkFtSRkZHy5/Nuq
NMaYpkm9/v9fCQQa5ohaH8aMs0OmutdsXwQnJSq8o8OnKpy3lYA2n7NajlDJng2U
c4GwKiQd4PmfdGNP0Y+sTu/PiVUicyMA6QR6ENhGwA4h6XZs1VOtdmZLIdlhEnVj
mZSolf590kSJ9SjBQVYDw5yRhlMN8Tw+Cr3Jh5da68AwjkM7zExXhjqjYPTNipcf
i+N6XbkCjIaqClc2r0/91XPy2JLS+JP7ZxQzc+LunCxKNFUdsOmLpUVkNoyb25Vc
T65i936jB797xkPfs/361k358E4dNvJ72KTvQucyVXocwMxsdQOWaaFOl4aqIyX8
Nmboz9qHGBQU8sCr9xbMpz9oqy1vuj63U8q/87/b0op00Pqqqs9vw4UoXfWXJcDz
w+vXTquAENeXBQOhWGZd4WenFoemE3GmZqBC5rXjV+2y4vFDrq2HX/sKITXbhzMv
Z0i4WR6ADpxfCx8gxnU6Xwuy9dmz/7W+gVy6lqv4KI96iRkjowgmdxVO6NYYzXQc
hDCnGiSZLDLUjULDNj0H3sxi6Tlk261/x/lMCN594VdhVi2380+eBqRI+/zIfYQf
R9kK81AFJgQzI26RRmjc1qgjX5pxthcIeKDRFReUqGsNar4YZl0JlEJoKedrMrty
yfQLnltEf0oRLoWR9Fn02LGue3dno0m0hF4uKPxBkWGTcNRKw6ELCPwhVAmUE1ZH
QEJXVhPw4QtZMCUdTmNehTxddZRExkbYT2qJbanz8GZ4DuIuOfIYZbK6tjeaI07/
NE1xBUYbAzJZE95LLN4AWJiYFURw/b3CYVsb0G9R7oQptGSZgbEHuINdJnTYgBrv
vkoLRqc1btVLf/ilLgmZjVnwgOaojLznFAs6bABKR5Tr08A3Db/pQn5C7JRwl8WR
XfDLYMyqlRUGwzx23GoCufV1FSqbF0lvJnYYLTuROg78yih0cpqVLX07Emh1/jUf
dZZRqZdxwWGmb0/Kk+cB6KLkv5b74Vg3MbN+xpfZo9fzmfuWsJCny3PuJ6wHU+TQ
2P1+Ysm0t4TgrY3eBIP2X+P2sK3/hUjcfGSKXTTho+JHdyp7ZJR5+iIpEmZ4nMKj
tA+0x4M/jHdKHtAIbICd2X7ZhLF99dAPUAJ235iPh3+xntBidFojJc/IzKsSQ7Dw
5HDEpay469gz5eu/W3lwu7JTChprXDDPY5tU1OK82v9wTnpMQnyzkWfwPU7skEh6
uG372PdR7djnWZMMiYazCvOHN7BklPiqUp2Qpr3Ox6F1VqOb+Ub1ze3FziW4ILG6
JiWAPdpwxO//pl6TeMFu5LzF7C1UybFT5meEXO231LRk4zc6TaG8j7w2j+tTPOBv
B4GqvxJdwBWag6erjdEf+SWGvDXrWSyJVHe1zQHuUnbGD2fJEtEvZ9YVVhor3zpb
RqU9R5+g7M1NQ4t666vddiY19+MvqHqtrwBr/OFpaiooDEZQfe+hUtkDtFJlbOH1
8hSbcQoFP98aAE2+I+RvqwMr53yJTGbxZQhS5x0Zs52PPJHDhMXE7p6WNKPlxLy5
AdNrMa+JdFlPiRCNZfmRht8OrG5UhFV53NYwUTVd/SigL0HXUDHyHGvY2XFpf9ku
Vwhw8z93LO3jbf8ub523fWITpFu3eOAdihTHjBaj5M+6yAYrklNgiAAoP6bryaNW
QRh79RdHrMUKV2sSv/q2B3prYeWZQedJMaJj2JL+9AYxJ6hF0yjzjvQG2N2mMY2U
sLkq3vZBOttWHG9SoeeppNfBcDGNmGjh8nPA2ZOcVMMVnylWw4QwERNIb8EKsUPE
9kp4/yIYJxfnemCFo8zPfUZmB989e+2CJ3qn7xwbPeHFz4dcwj56+QhUE8a4l0Mc
r1uJ/3MZCOVTnpTqXDBvF5LX9Dwn8jDIqtH6dwZ4uYVvaBWbPoMg1ltBLXn+BwcT
0LNLguFc7L8FUK1g8OcYQS/eG1539TRYSMowbxZm31aaS8VyqZ7TSFFkp0x5ZOYJ
WPf+aT+t1NDzfI7iv5SavqT4w8DdZ0ukmEXh8AkdhdVtE/nHektxe/zsVKf5jQ+e
PFSHuslQw+7IE3m2nWi7M+NUPg0JVQyiHdhoZkuwtqTdSGZBeNR/Mqa+vOW0A582
/GBInMaywJMywuyv6iFLBY3ZNaJz+7usRfWeJ5XRrPQHWutSYEG3h/Vpwx6fq6h+
LYBPYOzcXdFpyvnZ5b1sR0Amo2fauRYMwjlO50M8xsj8ZUANHWyEcmK+sXdW0pko
44xREifywAtiATAFxBtqhd+qEJvCoToD3ssZfrnHVn/lIXQ7TP0xYVUuRqfpLgC/
VNOPK7d87MNZM8IpUVS+TcuQK/v51Y1D0f/hrlbtK1wxEmRVyvNHOIUFX/uLPpzH
TJRH2bvdUB7JKu5px4c1fEiTiKNgwA8bVZH10jlRQT0Jt9DFbnFbnVS9b0gMhgn2
I8s7qpR8KdqjikNFbOUhhXcgngO3qhIrcrXhwCZrlnWasiRNA2FYWJlWqJqOzLV9
5Neoa3YsYnoqQWBYA7Lf6QZtHdYkAuVQULNRxDbTfst0FkNgkqzFhHtZN2HtbcBm
k7peN/UkP6o8ed2Brr7sTTaywOyvBNLb5N2lOSExPMb+JPIO0KorbEP5SLpF6VNd
LNTYlUQQ+/z+WgFQLFir7uKmrHX5/GuVD4XUqDZaS/js1tueAKFstnb0HvGIEZrx
81NnYu0aJ8pWyUtaLOzsfmqW+rjLKCFZ8jXcJgELdaDiPnHCheE27qmV519samtJ
fL7P4duYZeYMmQzQ1t9LqQtlAvZ0yK3+XHK9BspbBwKKys/RhpDPr9yKNKHBxMmN
qsSGpOr5e2ngVWWo8xA7c06B4NOtDY6VNflg4mvb1zGqqSFIexwdWKl31QJP6FAm
CDbdLOUUEwa1uspEZuCe3DtmtvIz95S/kgtUPuT9xdxIAOzxmR4syJL2k9/sRcfk
6PTco88vFYHH5zfUtNeO6DGZ8dxsygj9L5JpjFmRXMSX3Au93ivdec+A4wFwytHd
t3SbF94k3rG66U9cPgNdjS9Dm+lXoXz9PRqULKfPeTa6TEaQvnbeafRNCPCv8lF+
c1G+VhabVhiNiA/YW7w5+2L7+JUkNajaw92N40PTra3/Gz4tbdpEQCmkfEeIvImW
b2/MriJxkWF2B4MVmcJnhd6hedBMFUyShY+T3lGlcDlIroCiiFyQ8Q3THn0h/3ZW
lYSp5+IHInDwQ8oncnXA3XI+j1SCxIt+eiZRg+KAIlgH6VhHPtMH/3OIvYVvklNi
i26Peep+BzJFP3IeZWbtsmkjIyvbN3dnWJAaqusDQiuX8xwIH++fIov4ZwDwqL94
Tv5OmUu/65+dGct86qr8punT+nFi1BycGa8flUEIMTj/hYVWJgypBP8+wg/3PVHf
yHUlku19NdTAKCl/iRcbXrwBipJ5a668qlgmCOoUbJ0m+B7GjBCpOKRXnBVz+1gu
i/s3D1RlKdYlIZa97JhcDmfZU0VoQXwsL7CwaBLJSdwH5fJLviBwgZPLT+FfFFne
lQJAUwOj/nW4dpkB5jTLNop0ZEfwJl6n0qN8S3Plgo8KkutMvojy1ELyJaRSPds2
PB7HdES9VT5iwKnD+dQTojsueEzot/TkUacse8h0uYlW+D59AkuiKQchUxJxQRRe
2y3C0mnsWQGMQjGIjETosOhFWH0EfeLA9EgxduqPqpsunoE84DJsFXgM3RKcqYGr
kkU0nITt4F+UGkrHlpP79G5EEUXF/pU0t9ivUBf7jgrxuYTRyjRXY6H1S/oqVCzq
qjPuQ1RMY+poiJ/pJFVGVeSEr8eWPpZoUoKFKxbH2r26Zluor90L1Myuk5xy/ofW
9FZziuebplCGT0sQJyZK7f5izkBJX5G/bV1KgUTWACWz5thv9H4rwBRoQ7UapUAQ
0MkGIgE7Ova8cQzGeWoAK7LTuszttbC/qOhcqDn9NuS+/ZIFmflZKD219ygqHdrl
fCtHOz+VpQYrONl+7H01fhL+gX7/H9XiICW+3EPngBjwgJTkmH4Hrx51ISTucx1P
xp1Kp5FcujCl2pYJBlOjMPyubPmQmalAJK8dTPpYRfeSTKjwVY9nUG6ztDAyS7FU
emAtfpWx5ek4O2N5qHg4w5H5bFoQogVIbRIM5EKntM0PYozIXN1KZw3SQ+5H+u95
yuKefbIqilhvCmcEMsvpASB3DEFLkJidtpvRfVAHOgUoBVbRmLEa7aKOSVXcfgvJ
qvqf/caCV/lYGNQmv/rTSb9cSxP3MLUo2f36OpMyrOBn7/TNcyXIO585TZSmEiNl
JTNYwkEL0xjpGQx/ASOm+zb5Uiac7b2C7G/RLmoZo9ZHFi99GKPLtqd8BBleRrge
E6H3OutY+iuzTnKTijAuE1sV4eVhAgPjcuMG9VvhAUynN3+9N2oh2D/uYN5FnaH5
fRc28lCqBfHMRWeA/bCRyd+ozwrjiaul3bxedacQCgCO2ekRFbwRrppLfL/VurRJ
PS1h9rP9jzjMFrm1Ry5BERkhr+8Qj51Iz0XC0RMQxfRdKkquNbhRSjQJQEKHtYxC
XGmftKsrhngXA5AuqhxOp5Xgl1QwuFLQDkkS9m2y9RwZkG//JMm3r2kGszDt4tm7
TS3it5kDgekGugZwrjp1gp1SVzZTbPUKtYxFcuDJwE590/85N5TtZm6Nrypiep3f
fJWMoVzpstJGbQUaieJ6I4MKTkLDUkOZEHbIh95iWIQ7arJJyo21u7x5tUF/xwMZ
k0K5k6DlrP6/CUshB0tYdwOCfENnLWyaH7Gkxt9WSWYASvy8g2gbJ1oODhcze6fQ
Te2Pw4AeYd3WjeB5l+FKQlY49vJoYAP8oZYJBc6bYxlhUJnsAk9f4MUpy8CtZYpx
lxBra8ooWLeJiVuk+TaQ7VdvbhxcX9V1cvyzwlAFCiXcDhnvJ8bLg2RVVvF6k7rd
itw3l7dK/C2GlZNw+p8Wd2MJF5QfiWTuFIhCEVqZfKSHNazCtuyBnPCxbXRIYiyh
LyMR2uSipY+oGIVHGYO6eL1rwNME7+ba5zDatCd5JSODOnSmShV2Iq9J+VnhuiqZ
CmvhRIsPyzjuNM6ErzshH2n3UWv/HpQYedbHGqi8zXgZ/oaoSdFYMRuN54b2StNS
KkuGEG2zHykw0+SyqqHSJRzJlnu+6sSrrv559OrqMmrnPz9EZYPfSdKMxo/sc1ei
PQRuGDMCTFL1+HGQTNr29aTo3pfGUvL5T1dzksdUdBTgDOXrAcO6j/P42/OKi+XY
YQ0sC9Ey37ISWfto3wmDTGykAtjldnCKPMbnC44xXCE1fAgiJlZ4anzyr54xvbjQ
304i92zSVOb7d+LPcfCrcJzDPuSO8Zw+DbM5QXanVvJFa5DMn56SOD/X2eJsAcKf
Pek4KdmcA2NTk6hxUgsqTKgEmu9gv+8r6gFsoA6JZWG55gU9dYso+ErSnKF4JzvK
WfACpZhRhFzoBnDFTSX1/Va40JyDrAjNwMZ0b6yKm8gtYmP8/AWfx0tRSgbK4MCM
JOIZ+BTza2vmHdui8xYpIAu6xU8zEUsVPBflSi0TKt4FmmeCb6/NsbLz+qTBRKPr
twOjsojtBTeVtwvlDJCrzxirBxmhPUBSAGG62JKlloZdUI68fzQYvshd7SRwyM4D
mNZ73lW/aBePl1QjSB8of/H81v7zrj62Yrjcr9obK6SWM6W5MOiovPGf73nf/Pt5
9K1+N71+xlRt+NxuhpoLlrjdVrXG0hla35iedJGXpvuqVSJtd8jFhPQr8w1rQ2ae
tTAJYG3j46Grk8fu3dkYx/xHvvQkl5PEfIo/2l35iULyuzDwDkLrL3FVIU00uLpj
wVSEwds5WQ8BEqwTHLUKgnnUdJiMCY0H/ZaecDHZ4AprVlWf6wMmYdHQzkydtWyv
R5YXODDF0tNW1Ioh6CgzwqEG3Xdao6VP+RdVAUVNeOOUY2KUw4Bh6f5Akz3X/iNK
HLKguRrgvf5nLImwQ49jHkSo6uW4LceDb6FXpvQXMjDy74m1OR81AqmCtK+WbcBW
YqWwsNh/Bku+7wdYIvvcDzq3NpUkBCIoNyRHb4aXrVGBMnK8it82S0zWXNHZrA59
ieNHrC2LtgZGZrRAZ0C+fbpL2cXbEAbmbUrBsHmy2aQefavqCM5nlUGNxW8m2UwJ
oUc00JcY6+zjP8uJH7YxMp41bQAXZs1ODjqOd5OTxLQ2RmlKCSahMY3ifCZ/irND
NeVR1kKDiIMwDfVuwdlDt5TM+4cwL/qojuGXJgh2n6vsAQanZQcpbMXjfiF58Ztg
mjOSMeSqvpLsRy1nW+XHRP8gq+JcMKpx1IFIvMBHOMCt8wL5xRn+PEn6/xOYpzkB
1KVgIc1IHdsGNHxq9FolProRy4bWY8TAn7QTTPgdpFd8LCiHlIy88HFOtRU1oqbB
U9UV/Ztbh27kkE3lqv0fp4LCV57PxH+kT2vEzWG/VKMAk+FRmmtI+5FRmtAGuqYm
kIr7ZmQfPvSUry3ElK5Rr9j/cRtKwMKqw7mqjxl2vNgjX+DAlKub6BOBs3vhry0e
OSNKWWZKYi7F0I4NTmFMbtjzYptxjTjzBW9Nc4+jlcO70lD8nPPlbEfhlum0s1Eb
EJEBPqb33tcXLOz0gjUEIVVR5XCHmbfQ7J7UxjxGA4NrAXaIA5oqvZ7Cr3chCvsG
wwTZ0EwfcbLq8Ggvmmm1g98QO/0cpXtBL3XmS+ywyr0rVGjilZspco+rcJZXhNb8
+pfG8oqNTFDMzWcnY/vM84Z/S2tZICI4gKtrbYOfHX67Vlm4DY90EEts5PJ84ZoT
saxFnmGdeo5vGQTRq1K2B70vSw+YXODg6ax5FX4BQtKvkKrzIsX37Hy4DkSzJLyw
IZKBXTGV/dj5pJ8J9eHr8l508BCkE+a02Kddhp3UAjjU8fZR3XAxD5GnTLVgYUJc
ggGegaRHkkhKUEDntie7qi/gX3sLx5/F60nFJOyNixVszHNIA8tYQTheAZShYfit
TGxGoRl4Gke2pfIa2H1UtoIOXf0fmWKErj9iOsU7+XElFaw+CnL3sKwzgwVI24kW
vw9+v/V5LUt5HnnjnBj5H1d1dtW1nBKi6gG3S1IVQ+mX6VWts9TZvy+0HCnTamDp
1hF3jTkHhTPxG85FuGug3SrTekOsZhvxPWKTp6jRCgbWkgWD3Apf3ryVsX+TsGdk
zqZrY9GVi3sh5K76hAB0Gyk/dvT1mPlG0/brx2nukkXjPCDmB3s+sGIl4w6sp/Ht
NqusOrgvdcGQsxF301+4P9yzPMd35u/YEzSihIjxb80OPRVrAGSQ+M+MYubP6TN8
QzcqG99mIiTccp4frzfWVyR8FWq5aNa3l8OWXFfYQvQFHG7RrLX9Quu24dYndvi0
2eFcE/uT45ovCAG/gdfJsUaIGJwLIIQBclEBLM5YsCqOGWx9AE7uaOUosJBNNp7u
vyQWFGVFllrVvIl72B7tYo2o8w9B4CsV1Ty4p89wFqe+qoRS6D0OhkApBWYGY9Zw
YkTSZUDS1m/+l1v8WCFwPbpaQFN5+0mSGjb6Tc64OvCE8YOPqHPuqDdC5gFg64yv
0q/AaMQ5zBJzgAZjmr6Xm8TAL2DDYC9qyXPpKhVidf2VZjbWyZ+DjV0TVnVoRu9C
qgkikryPsPRS7/9qDl+XpCuJun2iW2JST0OOXwPIF3mU7Dc8K6raBlhSYbU0xDM9
mmlsO0pedNEmdN3MGQSu0pOh/vwDd7PX/a2dJV28s6HlCI9Cd+qdXkyjYnVTbcwd
pNTSpNlLFT6/A9PFBjguq3ezjcoVd5Gqax4/D1NLzzkHUOOhxOvp7bWCFqUv3GlM
r3FC7AMgk6ZTaMQ5g1sgq+fE4x5EJME1pzbTO7dI/sXAic8qbToZyiLVoB83lZoE
KuWU0hm5HLKGxy0RJB/vHv+JTHgYHCwCWnStiG0GqlHaPjxRH6S/QHYZlAK7Mlgm
kWQ4Wr8cfhyartwav7DcSKnqvgC0XXNfjPaJ94jOfR6UI9quZf4dKIKqhMDWJwCu
5RlgztcTATOG7PqPmpPgelsP9z2tfSKIA7VsKi4O/7EAkRwQZs6LiGXEkBsh6iRn
gSQwLXy8vczrQXOXH1qiT5B9Y9x1e1AWOIWsDWGg6EJ3HL+M0yk8AM/kesrZygQh
T0UOm9/Zdn7ZivVEjv7QaPakKP1Y2PaUk2ffj3PDUTkrfnyYCDIQvY2yUfEQuTZG
K8wk32faJhorLjixtaF9bLDf6DLBQdgPfH9/DMz93/dVYq8O3mDNebp/WOgZXfM7
m0HvYAfIgGbu1+srer7jAbAZNsJ6ZMEpKKS2glusJrQm8TK7V+VyArpUYtlo0p+b
6mCtydbgeA2/BaIRLipb9G+nxoUvW95NpgzmLooLl626Ox+f53uz0ZdgOV4ruZyi
ZWFCuOtSv6KmzPIhdN/PT9TndwkoiyTx/dfsYPAx+PXuLjAJJ+puEOvnSBwjb/s4
RecYGDqSwq446duQmJKaDlQeY/z0zRPGiv0irxibXs3d/4h2trlZGGTFm6N0+BvV
QwNImCyZOVdo6y1xjG3QFCNWKUW9kTJ81Ob7nbfEdBmiNJ3E6//B+VE3XaibH7DJ
Z4jJlz3G0LjPFBkr7A5Pp2rvYkggWh9f8qDxolDjLIARpS3wRVitnTLGHl9Gpre3
C4VM85v7XEjg5ujUOfm2MAOVuVWS9HmUeu1peE6EGb+lLr6gIWxEzzTd8My47nNd
/2NnHdyVktTbUNCrXP2bTM303Ma2hUi6pjon4LSJHmvSaVVS8/MJI16x5FNIXg9F
UFlneL4C7E+5lXXOoYyVUhHAWXDWyrzpc2bR2y0k5hZQ2F4ISND1QHWG8sVCOkzu
Kgx3zIwHMv42qWXt+sAJW5M2OMCCDIOfipNihX7qyzGlnfPl3qOVpUS40YcJTj6w
AJBuT1zYH/BX10lTqemTTxl/uaXkOmqZbpLuzbPqnnE/0jVneH/DJK1zVYpFxa5W
3i0v196FPx5AVqEE2JQwk421NrfjWqC0mPXm59tcdtV7FDd5uv8oqG29CGhA3ys4
1HRINcm5EdZTuTq9DKiqUOGZsqUJLjgJJtB6ZEvFCsNFtSNNwOibb3d9i1EKsIHq
V5xMIlIi4JL8o/Hte5wYz6nTPzN6rMY3c3fFPEYa3cTIE87SJM3sCt3ufrVmL+/w
NSzXF8dnq7scyNKtXoMHJAQWteBpcckQS4OMvmE+4sok6ZHVV1pP9X6oeo/JE8YF
VkUSBbSGsnLlxcM9WS88xmjx9GFyfFr7X3jr6yetUoI9NuqCojMdSl3p6obkzWzi
kXzzw2TgNsSUzp0F5HmhDKVq6yKGEJdFeMuRRcBvvylTIO9TzxBnSQRpGnbz2fdv
LwcTNixh+NqjfC4Hl6PFOxzQv8uTT7B/LebA3SXK2GMGikbNZD479w92dSY1rvZB
tSJravz1n0EBj6n1ar7PTmsP2Idxg7ahHEPPgcn3c4wCiGzUXbmW0zLudWMF50uU
XMhPAdLq6FZ1Ja0ShTF3R0fvQrnp2S9jTM7J03YE+14UhSnf0oPMOdvN67FQQe/j
X5bZKExkzJbZYoDLXL7s5ewCrI3JCn0AMiNUyuAHWa12gLz1Q2Cc76e920pxmjqb
Qs3PELQn5l8nm9YV3/49EQL8OQML9FdmRZZZj2LrYEGmmFCkWleVioM7N5G7OYB0
cERy/Hd4tA9YL+4WzQuqzihWnQ6xq3qzF+Y0n4/926H6Q22bZrlbD7lP3267W+98
cs8Bkq2HfVHQrTOSSq/xlsdk4fOmSiSvljpLkx8u9A2NJ9oZg3m5gO3c2sDrZkiI
7w3H4rg5DcUUJHgsFcmyu4QgBraFost387tGYXBmlXpyO1Kc73Qam1yrU5W05bBA
Ec8vgozfBwgwNyD4rhZBL1TOn0XEzdulTPGy1X1DXCeuUGOjgmiIZXHpBh/TDNGN
1yxdo3IgBxCQLGvqZYsX0PAe3oBr3yHPMZ3vbFpxapk2vMGYCHJ8Qgbeud/9TxOG
FXFImDIwdga1kV0ioKYg7HYyDSJ8z0U00ffXnn88m6zgsZnu5OVTaBzyySgvqxIL
BlYvEG+hkECxHuS3Y2KnHyX4gYacTEf3lEQanRR0TcHJevQRo5BFrtZoGnYdcdPZ
uDDzsN3Els6WM9bBM4hwPJ1kYyWBXPWSpkv+gJm7xo6LViFZUQHgp3JGSFVYCO91
uUL7qnfJSyEIKn4X47WxCImxKrysRejF93j7IVM1BSPuZhoiZvLhSSu5zrY753Gv
FtHnRqRrW4upGvPho5P9H4TbVoU3OPTu1uPblExD9EuN/A+zGH3rQkUf3hkTiyhk
M8XEsafXhgt2NTQGhfLwPHzunkasiKHi3VYuJa3i/joFzd0Gl4/aPMjDS4CIs9/a
TFqC6/O9cOR6sm79gWl8RQSVGlQ7N4LWO1hSkYyxAhhRCbwGRjfTCt9PtPTsESQE
A2e42wmq+smCCBuaITneG8GUQmyPzKiX09I4JNiSbgiLtXlqHe/g9/JmHlex+Mok
HpoDP6Ye8WlZv1IIq5EHhiPbJ0ghxMkBsq2MhbEsMoYkEsBEzIqVF7hHfn0ln3n5
MrfsbilQn603U7QGS7xK44Zm4XWafbtdZmV2m7a9d1ffRmlwRMHeCmBV3LBfbar5
Oc4qwpW/GK8VJSxS9To6VDxzVxhP7Z3clT8nCr0E/A6uf864MlqfZhXaQM7zpgWt
nLVV3+s0awoIVD3b8cKJKSx1W60fn8bFW8xlsdrKLu0hbWFGTxvUzgK9oCam6l4W
Vql4Yyv+0AO0iyouGBi1+3D43v6WMflq394nDfvIiJClKIUbnpMOm0wrcKN2Wtk9
PF5jA4QxScdyFtDuYdEd+hL8unU54V+I0kMdgenWlASAYkApXQia4LTswQXZ1+ks
RtPZLKrgDulosN2hbjEXuksT4lvUvOe9rL6bJqVUJAb/ZDU5NGfutlM0tnV6mEra
vQAw1GLcHvHLYujwIKhyrRuBX29iT4C6f+jfhKrFkJA6GeIalmMhkFLQqs1bpejn
Rb1ZgAGSLxLFMKocx3yZO45z+bTkvHHJ9hP5TlNYQ8uS32XK5BEgMjgoI8o49lKf
PgJCGVRPEfpgnQO8G59GB7kFQWTGGjSWxiCwUUVrhF9tBCBlxnziqXRhDyC22m6+
ORVU8ex5MnoZON+R3DXMthK8PrjtJiXiTrQBxar6cHi5QMTmun3cPn+dwzsmOPgZ
N13i3ehFKPa6S7uIr33tt1xm8jYMHXVOeOx+Va7yjEQnUmZehxIX8wszNdwFmtm1
fglMMp74hq6gn4qyc624okrtoL3Fp9icIQELIhnPyOnMOkNOk7KSaQqAn6f3bPwp
1j/VqzuckGx9CHhs1JzHGe2l3QsiD4ZYVRRsngHNha6iA/z0kC1u0P/vQjmfh+ar
9R5wf4QX7lZ/wn0hNDJeZ0OfQuPXGLitRGWC1Ozwjt1KJZ2Y2bWjnpMKeVEHShPc
kNpoz52a2Mqvg6s8MpeGf3MGvGpdTv6R/ydmWj5jq8lI4HMHfWAOgfRF6TQLfoBb
AcFJWKewPYvvW5fV0q+XLAcMMsq4P0UnUB/ab7rVFsuSA7kgTDO+7i5p23erf5Rg
tXVQuSd7VXpOnkKFtGtq8zVdn8FxIp+y51UOL6xQf1cfuXGtMMtPNPVErt13DDeE
WMleGi3m3DGGoK2j0YGy+Cr+rlWUlKiLnEN5W0xQdWDxYDubLILcev/rHF0csep7
QIXjmysnx4LWkvHptyvuINFCFMGVbtBVvPQw7vmzN98BIXNb857EDvOfoJs/0yDA
wsY0Str38v4zkPBBVqwPrYn5F0K90plvEkZfOwuvs2mL80+qITBWZNtz+KvQwfga
TodoqwBtfDc1t50ElZ0nGZO5CwK6Qs6iVQezLNeejq7e7GMyhoExMEnVWFO6ml8W
GLIKohmpFPJPm5IM/PBqDmXZ3lSIuq4VjRatk4WH/B8NC2foxJJepY3tMf9lG9Vc
Gsjq0oH7PIEMVivwQgiykuUTiFp9tL5iMjmW/ST6rwNe9h6t5CG2XR8JILYQuhQp
uZVy0a2IXhG2LqWw8KGPKpw6XYzIjcDzHwWmVZpPBgJfDdD995uSaHjm3cj9Uujm
9KM/D4kCQ0bHGNynUOZ/rQAxGtZ2ezzA6WcPVOvYITrRowXW239WBSUqcjHnQkRu
y1a904EL4CrgHTn3TcVRVcU8Kz6GdpSwiw/zsxAFFWBPwLsolhnU4w0wmjY1kUd2
UWRgizuOzMAeNrwVYtPOaj4Co7K6TUFkmi7B0GpSRj214Y6G6Su+LNzTvou8tVo1
hJJBLipCVTNUHky3Lv7x2BJtOtQpslbVBHEa2EfISrocvCose2Og/1DaerULjCMG
ObqXJtm2AJCeYI/H3ZZA6foVKAwXkpDIltu5U2ttLf6vCBb+BqW9rz8ZYjcm49Rk
Pl+90vhVWFRFXktTu6Fz0YPh8gWP/CXkHVHX+/SIrMhtx28ZYdz3X2emsQrv03Ee
iCi1mYlrEUU1HnDhIxYRnIq9nEuQ/7C7Ab3OD5FE2E9ZTk3yxgbj8clNpyI6DjZy
PUL38UyDCgMYHXHSvCEzqdvNxkGB1cwi6ki3aKkwT9ayxSfXTK7R2P6kwFxK1MQ2
NXCQz/R+Z2bW1fE7d2unXWrtGFeMF+/sjtj2VjMxjYMli+fHO7gPA554Xq4JGWiA
bZ5kllr1jpiWwQzvSK6+M/u+oCiY4r0yEGaTw38jLunue1b7pgm6jl+G9faoN4IP
Mh2+0VBUuwy9f0HHREh5mZHv/GDOn9hp2rHIGo4PEwQGPflN9yxwMi6nlKAB1W+o
eS9fFIG6e0calj07l8xbbM/lzq0qoKYL4TL7P+HVCMMiGDEgGyN08mBAFg40gX4e
gMxtlbXITHuwOnyY/ui8eLOrMoIwTmm6OA69iz1OVYph+RJ6pl1sJqf43qAZx70m
YoB7lLQYSHOVXBoetdCBKbvRJ9unMxICLdnlNJRffh8cAKFKyx5VzRCIz9KA2eoX
ZS9JAGzLPazCs8qPJ3oqvj72LxilhBruSCEOS3/UXQj+ioF0MEaQHGWQ06VLIv0k
NbOCeSizkkQ285TRk0O3Tx7pG4H9HER1UDwHyJIDL44r4wQlQJP703aW/c2MzFaJ
8fbi4OEkQgDyVD2FFtATa14R8g5ir4frt0KKvoHSeWV6fJR90X89mC6lRB/rXPfw
wDAES4KZSqkhRH1KNbGyIEtfk4jmzaabECMsadx6ZfQdg9D0kps5+BeVPF9Wagjb
zlzsZFPSBAOVp27Xl0bPwU+HgKk3hYC8CJRLrOSiu0IBUSaE/Mpu1BYx/5ZBAzTw
uLvWkEjDyDUb9jAfLmbVzdpoA9X7+nOxat4dZRouVfRUOyO1mKgCa6Z6Lgboobs2
Qg8t1d4me4kyX90P421uDIBt/nZuixExJGceQc6xBROo5nDX3Z5/m4QD7sLlAw3w
zIn7G3lWXI1z6c4CWNoKXOKhGb4UnDWmNFurTeP8YNpPiUUecEX4OS+e2MDgZ9UP
BYZsZ56i9PFSVlB+UXK5acPXECOwVoFv5jeMzeG6RDCjOng9NTq4tu0V+UJ4z1H/
3blN8dnThSC0cERG5/KZBYQLniUUC3GSJRFLknb/5gPBOp/+sUYo6PPZTz/nw8mA
pkuv9cJUWrCOZ3TaasbY1mqetaB0dlMzA7BK0t2teQ/bltaP3yFoJ6Z/QxOy4bJL
YfS6LG0zlWCsOSX0UT8Ag6r46P4SAe72XcVSr+iZaXbbn49+KdZP2KU7oYl12Rre
qitAnIkrRRNYYKgY/E9JkZ14eXZItMcItrCNK0PV2mX1GZCZ/HnuXJns41eh9YxJ
xo2Z4hXCrovU/AUoxvGRRTfqDblUiCLtIIJIkFKSOAn3eqXZ02+MYaNjIv02mK7M
cT171K5EkgeOsLa/wIDpOaroIUR0aXS0ZjiRb+2v+u9/xHGK9kh1l16gwKlvNoIF
EkaVyWYBswNyZv47hyZMz8cVLBooBQKcNPGektoPl9Yzj/IqBNbHlW870D1hu9jE
aIU8mHuQioShOW8I9xTQyIWUvCQahhG+3U0f/55ILyLOF2qbCtfKyA04UYsmX3JO
5USvCucSDUjm8jF+5QHyaqH7StqbWdQSYE7wH/bm5SiE1bE5G6vm03gQ1heIdIXo
ePDhc5Vd5dbNzM54m4Cku2CKNHqYKJvp0Pbj5X3elsZDPpen9ojzVoQ0sC4Cc0Gu
ON//AdCbFDZUN6BrTwcxHr4rJnMKL3Hfgf5jyEEM710q5OHJMv42PMOi77fvoGgd
f+FbSroLhwDPxYGuVSedJlLEu6JibAG2FYgeKavyBuTx+bJsT22s80FaWQeHac3C
21Epl54SNIZpnJM5EezXk4VKtyjtW8utGVYlLzMegNFXi0MmoEwT/7tiufMOSUr9
IlVtbj9Rc2koaR7VJnFW5aMXKLdHV++7SwRk70vxduG+1C7qIND+7wU5cTKf3jFV
F32sRB7ThYns86fL3SGUDBL0s4JSrqDtT+33d7cC+S/+9znSKJHpoNIKWvkRiqeT
1aoAmCude+0HxhpWTgk+LQYvOdFJPRbVIoclQtLLMUgbq0tOW0LoBxE225/8PXgQ
76Jjyw/qlJVsBu7j0dIIMEee7FtBK4l1wd+utVBXSuJp+VwQ3NqznaWikNJ7JeGr
/XPTpz0yQnqE6XPMVWQe5yR1MuUqszlG+nqyHJAsGav4XGXbjOJ5TDg3ZOC5aC3p
wn2VdZGLONrBRtbfOaXUlazmGkBXXqNnJj6jrZ+ApDlamfB0Vn1OXNfjYYN/6/sU
z/G6KrQlSWpwaMlri8RwhhGgsWNvV9htOzYPFFgcoNTTtIqk70EBxyTXsOxcdnvU
n+0EsyM8eKmf95nA/fge7jHGIP6uBw6Yim1HBpKfLozw54hpLnBYW2FwCt/6NGSq
eBplejX+RuS4mPGIPaYdzMy4GyorP1vUlQ6TQ/vcc+S8MOkWKuxX4cOJynY2hBOW
YMmSpeMXOs8/RrTh8R0wNP6GczgxMNjLYx/1rcmi8WMrpDYxtfnA4UGaPgQBT2BH
YlHSSaFvXEsDWS/1HzXtaey80UIbUmrcF2MfqfHS6TkP7bfS5G7sU0Sph3UfOOym
aCtDMYmZpubKk3FmaZnIWFBVoXDBTjm1kcMfdENsafFSYkve3yXG2LC4Ak49u/do
rook4pDtpiMV5LgkAxnJ4k6CTQqFXIDJtKJNY0eD/Ttnzc1mi6++ZPE7w82HJBe7
zHXXWi8ZEAk3HvKeXmR8NMXW4FALQVtw4SlxRh/6RrXIFs6tvS7PPolVPLq5i3uK
c+Ukrlg5JjT+ReBkWc0IhMPRXqXKDcg3BRBkBWfyDiv3L9nVK/Pn86iy/Wnrv59O
euXPle6gVv+dumqt07Q3esLQcquk69s86w6cjWm1I6ThdpjpzERSDBkn0Q6hiDpu
Fi0WptGivujVAVPugY2gHJ4aQHgbNXoIGyYSQi0m7iSd9N/2pRh/J+EPVanv6F8G
m+U7gxRcXtG0nBgAIGWtAYP+JG3jmMoss4Ie3qf7aq67v/objwuuUT5oF/sIsT3y
jogRWxDHTIHHQOMjeGQvpvW9etnHdhQeGMfrZw3jHvCFHBAO+n5nUJElAJGBIICh
mTJsDGj2HiLRjmN3OINlGMJqgyrCBBdLdjkBVZfihk4KTVTkpUxJXwyrwbyyuwaP
i7nTAivaBthOpFIbSqNfyVpr7wDA8mGpHaH/zR06Nzz70aofQpscl8CgBwYG2Sbv
p+/9zdvIT4Z11tFrsJpXS1wbvyqypVf9nVDAlZ0QAR+NrHlq/Uf9K+ZWBddjcFK2
TK13rTA8OaP5jDGCaC+gICvezK1BY6mGhiuFWDqKOxaZt4fcdhzjrefXw5U8yhDn
NKxEOselnbF3807fnS7UbI/o0nIVF31UfM2QsILVhrPQyk28Oo0BfTsn/09F/DTn
yxCr8TuH09aKWwwZE92bjlVpHmIbIRj8V900u9IGUsIg1ThEa0Vr33+tMiWhXQZQ
wQFTxgn+12c6KEl+r/GufxaTw92gzHHmI4lJTG64CRoKzYTCng04C2JqamvXTKvh
cJxLcmqeA9d0M4KecxSVR+aLG/kU2T21KiqIluKblb2/Hq72qo6kEiaybfvjJDGl
y+oHCY+NR8jpj0ZpcQEuesSGLAkdyfVQ4MAUg3kv43iVrCJPFdUZwkYLFWcfsnp5
YBUR+ic2mIcIGya7OsdhkLF1wbQXpJ8ckjNhxr7HpSQtRj10B4aMhPa+Bg/CgY12
+6L1QqNK2WrZmOhnhjOD1qzQlbWFO/wSwACCMtjC6aHCdMfGIeocdXsVALBPMfXV
3oh7yHnDqAFVp+jR+n+PmGMwu+k77fueAA+fBAQ/7+/JEbGEAOG9Qp2jEAHTx9oz
TUHaHmQ1jUekWaNw82B0xPuzVnKeDZIQNujTJ7yM3PzHTpLQgBP4t7Nbb6IXe0O8
QbyWQdyPNfxmG5uQNWZJ+Dii6d1YGwfEQhw4x33SNdFGE0nPV4bgYyaftqoLNn02
oxhMOEEuFdSg+HaZZkRnJZWw4eVrtkvlXAzzH23e951QsR+OW2FHPM4VTQ9KEZxq
AUH/zf7SiqT6jNpB9rZv3BX5SoIIHVUHgSUNUXiR6dIEtE0hSlogO1/b2KTrMnbm
nAmov/bn96DHiVwVtXfxQALjfiownulsxvN90UjqhqgKw7rh/2cHe6S+Izn7/KBk
x4HglYBr8Isu7DTC3Vj0TO1W2CPpptH24agnOtCUeX3/rQGGJIzDKHA+czqxElqI
IGswt+slfSFAusnL3t1FOVXN2VpfPVxmIJs0W4AtddkMgpOuLTj+HvD9njWlxLJ6
8HYpUz3zJrMZ3PcoFXvyD/EKX5xPu9gfSLIXlr7bf6CNs8qZSsE/5yCh0OIrH0AV
0IIJvqc7s6t/q68g8TlZtHAO3h1GJP6VnaqJb7ER2LrDV5ozdYJqJ+gM7No8Ha27
TmVNRHDXLufWuIihi/zwP02307IQCdtY/EbdAuthe/Z+ElYatBBSWkrXWOokhgF6
XoYiYO3Yjaq0wLIn8BAZGtK2eHfnmVpj8sB7gpgTEryBoiE+XTljDDkZvIcEI2e1
Zgi43o47DIXOX7aHL5DFjn0iuSyB7Tm9vO/diX82ws/56/KBcBkhqEom6WbVnF0w
Wdc3YYGUzb4v2uCo2yYLIp6YMo5X6v5v9Ny/+o+/PInkzYLNe19sHFNL/3QaQend
I/shr5q7dpGZy5PhKyR147B6hD8c5z+EuzirBzeH/E0YQ1yKqP7wkhlPfGTdXBa4
BnYsiLlb1ZNk3UyqviFO9VkRn3wSOverkllDR/dlPIyKXSN/oTIDnqTj9sj0JZ0N
FV+3G4fYv5nv3agCKHzW9ARQfSFn1S4CTlTYU+MqhXX3jhPWiM0JIKy428Cwmhjq
oAytOebKidPuc1XFiz7rsy/8sXNezXD4pyH4l1gwCtD7B45te+fOCgcpBwdcvrKm
u/73wKixcXiXK4SHbGHGKZ/88jONBgo3CsACHIb0fQuKUPabV37bTEZGZHb23YQe
xk7mpa49FDeEY1lYjqsZPKLMxtT8hjxSGxAIzML1apke5PCYIyMlvemXhdr95W1w
CZ/1b5JEqdz0IA4bWnfM3B2IrkoPwLQTK7PH0nZzLfYzHw0KuiVLMoZ81hpLGln5
Zk1Hjt+F4peDg0BcmfywEJU2qke7Xt3dpWNFGlW8Cnqf3BCKvIjQfw0MHYVuBNdh
9I2OIuNnqv9PMjP0UrGvc67zzdjCmk/i5zKkBsKFF+hO2JMa3ceWD0ShCJSsW3CQ
buRdouB0AGNVcl4VQBFS1XN/GsrhNb5dSNHj8wvkDYbp1Hj3Vv67S8jQmebiMjFM
bVCYspkBUrC4mnFbA6wo/RvbohHS9p75Adn5Q3+BX88Bm4eV7Fhkd9hPXv0x+Uwf
w6qlQi1GUpHbskzZhXsMBnhN02OcXIgnudxWS2j4Lu3Et0dDcCV9t/z27DrsMtdW
PxuTJq61zDT5brztxg8dy39OHfeTHkhdNdGLM4XtMtikVB3BcFbpaMtwbzlHWnhE
bEYyRFUIrg6R3AgPU9gMdmSBbbMRng0gSIZ19+gZ/zVO0949ofxL5FYwfLuBKOcY
zw7gdwhl3UnD37pjdnx7JuwSfYBVLN9x99WAEAxf77EowoKGbIDPUOJrbizJM0NZ
MKZQnKiRGhuI0p3m3huPHA2/1QQY/fCj2NnBJjyBgSeU6c/TsLiy2xFdaE4thzJW
CY4WS/ebu3E8l09Drr03nxvyG33DaP/j1CRa9+JKWjyZ18EPkNmyzOthEE8FjjjR
g1syoG9vaZN/UINhL6Xa+KCRKh+CBfwoYrIkr+4hJEeWgqkSGLP+WHj5jJsP3Ona
fk967A49g6Uhaq7ZFaNfnurNTIk+optfmhimumSuz9GeFteNUFrXsbaNxQIKeLSD
uJnDpOAKeWr+3tbWZddGN0lmmYa121QEFy0yYOSfgapz64+MBCYqU+Z/ifw9Ibhi
lUHyyf3TIrN9VfjHk7c5eyAMw00n/PXMP6+UKl0PdzIrkK7YPizUIpm/zM17TXZI
RonUPQlRprQUEfpzf2crDOsrhxM7ZRkZhcHc1NUsfnhSw7rFh12Fif+rWiq7CTk8
qFWVxPBMvz/sqea2hRvxyb86pJ/jpjR4k9ap5yE7SqC947At2AU+gTreDNKO4bcD
TifxJlLUNh6cHKit0KMcBQflZrTInoB1QHYCrXLC7KPUt6mnIDailZhZ/Xt4w6uq
kd1BFujfMRvcf0HAnscfVEcPjWFpe00ao6n2i6fsk7/kg+opTVXhQT1bZeR6hgrk
pw9r9E/qQtUdjinSQZ7iNTOj+RnQwW5XKEOea4hjb3cf/KlaN6d01gVO3xvJI9Kb
iaPsb392Dp6DCRy8k0wqaNioeL2roBuyfek3ybfCDzxOZpWOwewmkK13YdAwq7Mn
bHtyQMwp4XHdvPInet23kmcf/f1jRTkKLZL0q0fh9mz9+IH/H5e4uqoYE3BciR8C
trwNAgeOQ/9/ju055v7zAVDbYIXUCzdt2EPGN2XdfVY2jaoDgLnpF0zT5peo08I1
pnhAlpHm1mqbFRVSr2+m673eKrNoBgVXOGjPlW4PlGr0CR8zBQOiaNaQTbg38tUs
FwATqUZKytBmKVSMFEU5dA108sX+FO/RarzWmZi5XVc4x9GUrcGqGomnXcTgwc0d
YdEO+Iy+4f0dXrGRIsTCzetmvcbCSk8EAgYFkQZiBMOu/wAr7Yvfw1ShiWMH62xS
nIFID7bAPyjercUeWoaYkrMREBaTCKv9aOvG1A56sra6JPDUKOpS0AJmOvFfgVGR
ZI4dxR524VPLQRFTVr3pLQhx871LAq0tA05UbueZkD1pIRjC4fkqUZZ0Myz4+V7d
/ET764IhxVQ/HzYSVwJGFChZJVwpC1qXYr0ZqN6cxwkLCXUjQ6Nhbq21xJrWKB2G
mvKi6R4gBnus3FILjxPJ7Kxm9HowAGF3HWwKgOUrqxa3XOT/9FxSPGwVc/owH11v
7NtX0u3O5l73KYRmQIra61fH7htreB1cwuN0jQNMyqwJziJNJEii1sFYmxcS6hkx
7YBVsYzjB0NvnNr/iNt8q9FUYfr/93o1gjGUWU/gWlBj+gJeW8CzmBiynoOAOy0F
E22TFDdkJVf2E/G9N574lqzphqb7B2LiZwoiqHq6Dz/DJ7JV0mKSw0Ip29vlwm/w
Udob5EmwiXhr7tlD1Pn9tiE7b/PulbdF579ZnCeaKhRsdUYdZ/GI94OQ5CR7W6lk
fPg7+1fy4P8hBxOFQ/F7wkmJmGHm6g7I7SFMCTvfWWMBAa5MYm9y1LYI6usUREoF
2RYeAyRLT+xD7e23dZbAUDyzU7Zm5Mji1pDWF7+JMdKnKHJbNcwSTdCFxBs74uCu
coqr0zkJQ/9lvm156HHIGPDpejn78YTAb1bI3XPUGCZ87iPxgHslLH+NLZEFO3s3
zHaOgMeBgnsRi9AiiC+poQ+3rqogaIPSXyUUqhhpvijoTpWTsjbtT3i/gKxbn9Nt
V1EymD2Wm6ZwnVvOgbP8TMHteZJOYQExaAKo9mypQAn6YGg7f8fv7DlNlfAUPAOS
BrPzofpBHA7+nTm7bPoTEBOdYqZXe2a27UZNW/Fs5vglPa1Zr9iyrMGUyoXuOPdZ
12M05NMCgCR1544fO3DygHZqHEbklIehQRtL60H0ehtcexllRbIARbE0p5IaetYp
0JCq81THJglmSWI3LZIqTDcNmco2j+s7BzLERt4QV3QH7+bYFLxpsdEqwvyv1aLj
VE0sgPOCMNiWASQO5fvSaE7DYVbib8sr0KYucgKfGuN7HlsBTF3ox5KMeNRSw8eC
YcH20tPXZ8bE2CYNoY44j7efQUkGAG1ONPDkBksESBUEJHpCSF1EXB3jClkLeYWQ
RoRpgoV/ZibRSc970KHoIGMsIhYJZUjpXtKSnu0JBfkMw2FVUwLVn9Pr4AMhBxfC
EIgiQYdWFctY3IsBTvKytdRHrZnsqkMGj1m64e250uo06VYR+mLTLuI1NrACiJff
jkESBh4pmqth15a9xx7G++YWOCvfnrcYjgmCxCyMokZAvSiBP4uxa5ZIcA6KaxvY
1Sys1S4KVEc4GqWK7mXY+Efp8I7OWXjssfOSI3RMJEag42+XGiVVvL+KVjvNAt3X
e+Fa1hykRaI3qKpb9j3N3b8IcBwCf/isTFTUse3U7nQmuM5MRMGHQeAXkit/7/MJ
QsCHdHGM8/wdmD3D1c8iSp1YTyAc5v/lGSxEIlu+n2CMoHQxIEpCwDrmkzF/v+tI
zOVhpcX/uLaeXPRuQVkXtnrQerwhfp2s0wZeQusIgXJSzG23aAf46C/LRjoeUAiM
Ds5zZRdId1FD9tVFi2yZmrw9ZbSr1x9WJp4voXZZA4EBim2tG30WPAQmUDrGg3Dd
qzYo2Bvo2/mC8eZNVuKg748ifnrQ0oh0qxoasRY5NsF7fl/2mJFFFNB07yKzIo5g
CRP7tNOwocmDefTP9YescPMZ7bLHgvVnycKAducfcaMes0F7Bzw7VJPpQd4nbh3f
wtX0EfKCM7XTuR0tJU3ily8R0J8crRuaYoQ3ncC7sLLJhc3R6bYeFZO9Ys8p4Sk6
suk9LXPkVUaa1NC5UqprZ8Gs1ZxU1q9pDATwEIAZWX6LoUy57eQRpHPE9fuRgICX
Ohi5w73fbJqmUJyOqYFuWbUg/Vdrzd/BlSSpyxQQneBjbp7E8ocqdIfkmdQg1O2r
bowxZNcHCAuMZ+adeOdUdS3bXTPWkr5L/n1EN1QDpOz5CcmzZNCbGo5WFfmS7fj5
tXJEJ1v2zH9UBC6sHK3cCaCAGA5LV/XMhWo7ewkMtaJRyP/kWUtj+rbNb4ebP9U0
8u+/2BBsrYbOw+WHegErZkXzizXqV67DEY38ENeXq8bSpJPzZirqLk/5WkaiNQEG
/F030Zknh/6z0KieI9R43qFyVvxlxSyb5eGGfm9qM4YInPSKLSOQm1illbumXx3x
YmS/lNYEbkT7WmT/ejbafELEtR4s3T49S32A8IkkWyQadUK22kuT9TJJwSSkMBHZ
uBoUOi1Ni06zOczO4dpFwAmXpoTAFdIerxY2w9Krx7ALG8XB0b6AA+8ugPtswxM0
XghOOcTgPFHbJOUqAk1jbeYHcVsbw0eF7nnQxBMunrhJm8eY7k8ACIETuQAwLpTj
0CcvEaZun5Zgac/5Ze1H6p5GkFg/MAwYxOAz7Zfhj04x7rEbQjLzZgbDhN+QIQec
peb6vqoOC4xea8qDNvVoj5J2tv5/90M5X2jo3DT7uWiLGTPXbI89a0TJQUwRdMMh
BnjMb3TZWKnWAi7jOiCS3Gz4sNcickbHvrB+4Upazt/YpfgGIkfIOU7GZWY3kluY
YY8vVrNAlB4k4wUfe7sFpEWk6D6sK02iKDtNQKWInP1OmP3cbTS5m0U1xbtktglE
n8QTTfAz3O2CtZC8TUImMhBndtrpggj9B/yoPtVt/18T+h1k74mxxJHXayq3pGpK
xQLLMZl/+2qzsYMnLCEF64FQa9g4kHdXQIwWlHxNIxm929LcqgfOeEqdOf1OKyGn
jlJADf4snqqrDeSn40uLMdcIHcM4xIVDnG1A8YPipMT5lCdnSdKECh8hwMz88lvu
EHiDNSO/naqMZgoyUOh6jDiMwTzitoBVX6SUVOokLEm8Wu7cuJdmAB4mTqTKFADz
CDElCwIwDXcOxsbrAQwOvpFCSwDp3Az9asAL5X0khGkMXuQ/7QuPjrS0ljarkfFg
xtfvFxc4OyuYRERJBlPOwc4ddqsY0wpuZPbfmCxuU1VQNYvL1+3196ssnxzpHlm3
tnOJV/zMrITyjzj4NNGU3jX67j2uVVWqb8O5w7kzn3ULEDgBXfH0zDUYBt4R4tyD
dxm6bwJpolzETCtQoGcZn8mIS0ibmOBtZ529YnyLdGOW219qCp7QF/6gXiM+V8WA
VCXKY5GRoCzNjVQTCfgENcsQ77qePMeWWwbXwNfp38PpKPjDNu4nNjr7o+9rwc83
vwtF59WL+0yiWZo5tABxYpGEWaHhO6z2ZlbpbqTbOHDe3M4xZEY7S6+gzsMwYFEN
QPVou8NhLlv1TD+oCbOy7PZzgH7+LZtwDv47olgALCimk4CtxG6c2avnVsL6kLvy
PhR9Vd8fvNrVi6Rt4pjw2iaiB0JU3na4stBO8USN3LK5eGOD4yKnJoLO88zgoBV1
mcvGi8mBDfdEJt/Qw7DYl7cZLsDXNwQh+gJiWe+teq3AUP+DVOlytgbYECPopzN3
NBJ9ALi6GZSoxVDeE/Zn8QR7otmBfrKe1ZIxY1OuS4bcc/tZSszYjylR8grD5u9K
8/qTatu7sjuTf4yxa+/u4+yopDOhiXAwt6aeVhm4yBuT31IUa6MC/xhfrIUq65nJ
XO4zrmJ7GntUCCWwO5oSWchWhvwIJiAKZQp/GXpq07YYKY99KMx1Do0fZNu40MrM
Ton0+gxqz6hhD/Bp2tvLDQRQ955snRY2t0ijFif/02+KyZ5VOnAjvt3LIRroOBqS
zeSyx3Yyhtyq5/bLBJoX2vJGMiaoHyrAPRpSbPMs6gtc2HytIMQ2NB+29g/8oIse
UrR2L6/dwWiIU1riZFainh/Zy9ETbYYvloTibXGAKRtFfoGm8S2OwklcjJol92A/
WwJvhj051+30f6D85V8sZil32kLpkZYbfsuapyKvFyEW1Iz7ODgk7rlhCZLnGaPN
2xrVP7XP0x4l0Ouxp3nnjSBaNtNA3EwzgR8MrLynDEX3xC8Qd/OoDcpsJfO0orS9
3QaZ+SlrCyweoP637UR5aw/LaCv0sBmcqnN6CqeHwLp6Bzh5byFAtsSi38OxMEM2
BNwt13UcX3Xoau7NoguimQPrfvHbY5RtMcIioImYTgnbkFWo54RWeVCpv++lvIHd
Gi7VqnSycaLB64EYfijVgY6W8Ec0xn0qif0PJnhKRekZCcvnkkKa/5M9f31siwn6
XwnXJSNwtT390BxsUhRnr7eUFL1h4RE67LRQciFPKp3lUwWDGAK9bhjVXNPLEwd8
oQFQ+Bz82kPIrBBdLmJ7W56AMqr3sPnewb5+btqSYaKrzSgPAGjzq54fv6uVfa5C
v75gt0/fihHWnbMnwOKo5rtXcEhKTUVdmLig9lwjruNtglkdOenhqpcES5kSmzBp
TlfnxqsD7NY4g/rROIeHe8LuAglyVkcEpBIqJJ03wLZT3ZaKm3ZrqeploXjlhMnJ
G5h2Xaadra/MYJFnxjm5q27XhQwMw72LfGLSDjqpqwpsgRqbULBeI0kFMT7XgWEh
+YJVAlSLvI7LmmexyUulDQ36/FdEZa3ZuFTLQvBFlO2EtPYZs1uW7Gv+lMBWyKPb
OEmz8/S9Jd3dBbipjlcE383qH5X7HWWIXAoUY5HG+IFdfmKHJWpfuyHjZVuct1Qo
T0DIj/X22Len89R8tpaobcr/OFdOSmg+7zsEdDRkVDz/wloin1zyQTcFpgK57Q5w
3vfXL46jXKNnOEobyPB+M1HEBEwVgv/b9PWiIplRRGzcgiEwjMu1CiTYeNuPnmN/
lex9cNAM4jS3wf7UgNzQTvlNU1vAdOyRuVg6RITfVxOwzSEAS8ThabUHRLrREQRx
odaWl6zfkE12p9JQ+xlEGWvRrI8xGKSiW90H0V/s9gjML2P+rK1gdfUVGC0MipHS
XTEBjzSWKkxdSIs2Bw6jznSseBAJbYdgUumYL0ZG5LRQu+VmehR0JipiySXVb6Ks
x1ms2EKw4aXPX7m9gFrFpQRXnWgOAc+6pXBg91prA6ulVDPSTYEJnA1aVgMqWcN7
ynaiN8p9Ug9XApmMH2h21OIEGeoCWIxl1qd2ZYEaYf5rSBz/6e2f2vDUCmR7WWOK
80OaHE8pa5jKje9ZZzSnqmkgK7MUViJZ3Jx4SDTb09dnxAFcRr2KiReew2l2kGRW
DmtVtEqjExiYIjJOW3P1IrN2Qa4v7HQjY+AknEJjzz9bsXlKo12cYhLjaBETjCHp
k1/WQQ9GEi73z8FqYwGxPu5Sed5HT0K+6jYgD4F5pXCjVYRt07iLo58DDKTCvz2V
weaJ6QN06aQcDl0a19S3isnVpm/j3DyGAEima5TbRVwcFIJDgNjdLi1K1GDYr+MI
knXnqBVACMsfaLj3kevxS0s+4QrPbcsmrcMC43UB1o7ALt0LfU7u5f6nBUvdvT+H
1VKtgLwei1faAdzG840RCks2plH1zQh7FFWhT52G1N4oZuQRNMLwKowmg+/ZCD6g
hVooWRe43aV4vQGiOw7iskxRNQtgPzj5IK/IulfQBT44W2cBMugj5AH6fEKazG47
i2iQnSjK1UjoajJZ8GrqOD2tssrVmHZPQEeHF6BVQApABBtHVATGA5SZGDPeu3Hd
+ptVu7rwhSLeDCPxugT7+51otiTEQ9oz+Oj+ejby1xiaSo66DG/9JZ3vyWDe+hf4
u0kpj43yN3W1GltIpra+weDIe5D4OTjGlEWyjCrMAbIkrFgYcziYmUtzD6BGM5v+
KRCuGDbT4H1uhYBJ5mA/WH39zxr5PrU6W1jX2tFtOvsQJbP/Zx5PTAlAEpZm5ZfV
cBNjoKdsRxz0kYADfKazly7M8aEtwPZfLZCEcNldxK3IcgZyd+csppX8PQ/DmwOb
OYUFQNzx29yWg6bkdO1qJrtbd/lmqB8tv7Emai+bhdaec40xfX6ImisA7HjvYNbL
ZZyFyCSk1UA5Q+OpiC182acRFBYLrDA9b504K2sQlPL0DEvz+hKD2BMGCVAJ08zx
L5X8NBVk/7xcH8BKM7pApt/wSa5wN3wmmH380vLlmEmxFN+6suKpQ3/p2NxHLrod
S3rd79I+bFtJVLiKG4+1gsNpFLgFnDnxzGfWgOSq+pcYyMQ4yUTHg3vvf6rsP/yq
eszJMfyZCKZJMnhqr533lf51wx94Wk9q4pxhdmin4577FAeiZaIjuQZsq0R/N8Kn
KIowteFu6YVY6pg1YVKGkpDsOlz6+wWgtysRylLw3JnPpAjl2fqGSpv2V9+Sa/Ka
ntwt6IgFoff6tZmDEjv+BXK+vjp2BMOvYhRxgcJsbGJIFvdRv/G6qBEImdJMh91u
p7gz5/rZz1huep6/ImaF+5V1xHob4TrVyOeKEWtQ9HjDAvUocL7chLO+ZOZveJaN
S0MB6eVmK//+JwbW8JKbVHrkOQInuaSBpUYMkaEzAiZwNtCCFoKyOv6ovS+k/fen
j65w5MNsR5PJprzmPfvQ9vUL8ekRaZMK2RW5Y1wnwHgPy7J7omuQ/95QeBbGSbYG
Nj8z2bCfCk4InA91ZlEpZOcSOcQwnaww48a+kTL5PxCxtuxwVNL1Wj8BbjszAw36
1Q5DC6nsm5hOOq3d2O46jz18j2456f1lr0nbNdVdcacBSInSpAvkC2oFB93HNY2W
ZGEuQ6t1e7sX7rFNdhLRoiv79pM6BWnk6nh8srQVhMcz6hKVDVhENHBZJR1dyHID
+XS8NYQM0BVqz1KcRl0Kl0N763ynMGrQV2102US8ZJXmp6ZD7MkF4KEBHpVVy2az
r0Ejz49JAH4huglq1/MDz5wGUReNi0nCcCOuFxo8eS+0mA/JbhgcfweApWoLHIxa
96idzvgUsyQGh20SXxBsDA1cWKCGDTpkVzIcUPEAtR07sbEhMPDoWlHad8jqu5Ca
xvdJVtOijsmbggCVS2tJH2Te/wGCFg1rRWwItmCG7O7J6qp7oPehGnLsvcfH/rGu
kliT2tpNGLkMf4LAJxIGj2kHiwTNQsYsuwJUp/SZuzcyLsdji72oqI2dalr/xxVv
O6lxwUSphLTvbPj+v6l0H7j/kWU8Auqy9s1/vTq09mL0SxwHAizMVsv++vmCNM3g
pg3G8Y7Qkw6snH5ceoTxLBP4yLgflTvD3GHmbaBhSoMM60csLGx5rHMmeO0rGiBi
44NWIMBsl9ys8LAUy+iGIwegBeJGZaWLJJSU4xNDP6aKuPOnYpbEaKdUKoF/fPdb
/CdAYGg7X6MuhArPqx8z1pXG4gAXeHYEJIBj01PxXSqssLepDBinBwCpkWFS55BV
WhZMOOOmtWzpQMSeSCsmmeDFMye1G8YCAl9BoCBU+jxHnxFECRJZ7mEC7CN1txPH
yyCrrleOqS1pgFAiZHXoHUQPLXc6+yGBwSwRqKLZavp1rPYtymbeTG1sjlt0nEIw
eVRHh0VZgWFYcduAdmZoq9uMr8W3zG7Oqy9r39ZPGsf0QALIb/yLlxosvFmOPPe3
Pjpm9wgTedsSgFg2vUQJuJe4dtVR4PIYp0jxj+QU0K3zHgV6wdaJ/AdgPmW0Hm4C
GGlExUdylzasRUhGkpkaNpzKDVVBc2/SeQwps8qdYr128sZSPOExlqwH4Z+lBp88
gZAKGwuqRmPAJ8oLqmpxOe8VCaGeo8l85gghg+HG+EP6ijJi1FtbEE7ZmADHJWpM
SF+ytgKuTMycF/SMTkTeunPJGDCk/FxdaFsreywzxq5JXlCMJZDPoNp4QH2aidvO
OkcK1dxg1vOX703ITilz08yx1hQz4YLkiR/cAr2+bhA38OJdSfyQZHczA++g/hGw
n/EIyk8vOgG7h2cehWYj2d9UbixuG5Kw2GSwijmNbgyTAfzChNUgYIUSz94+HOaS
8R7OKBZ3aP3+A7L3pjYuObDAns6VLN4VglFxKHtJ7JsoTsCSmkJFDDkTf8EuN0AR
2NxnyeXuKk5cW3tI4xgjV/XX3awauocsiaIrrhuH73vW9FvXEFOnyCHcGZfnoKfB
uT28ecc42/y9sryV0AaLrKkjQkZ0Q4PsKLenOMVpxWznLc+kU3VAVqhkQIoIBjEH
Fv5OXQgb7G13z+irWQFLs9ks9ZxvsPGwS6DgxIus10vnA4QuQo3TbzbeLEZmjKsH
5bLbvCwtZFTUG1W791FrvSXxcNGmVPurDgnTunwvzPeZaWi2efvTQHt5XQTJsg8U
VOvoTJRnOOXLf6WwQAeP5VPnE/ce37r4mnPRa6HM8SIKxkWDFEgnAfU6C4RMFKXa
vxpdMPKDREvkt/yN3B/4gqYuJDtXw8a2dlxyOM+2Nrwk9trI3zc5n5BkzNqg4Ls1
Jmx9e44ovY8XmFuiWiVFQmccJyb6XEKVNqv2q4Jo1K1sHMLWeakVA0raU18fXabm
o2eHDGNvNIYxZs6gIJ8ygCJAxXeQ3eb3oFXPrRpgYCqelaXOYPf01/2aNiWrEOIM
AuZk+MhS8IrwF6RHXoPrT2x1LqpRg4bm6re6mU8o8q8YN0aNg82ij5f5yN1WCQuP
y/K8bgsKEjup06HffIGkW7PqN8RIKeOgL3xJXNgWnwGhUSYWgZ9bUhDNctnjQarE
j547U8Q3LYyK2AIWXOHi+C+zaXWx+V6mcvsWreixHsimAY+xQLr6If/zGUOT4Wyr
mcGeSjMSS7OIR4BaPflegFr92p/7079OTBl2qQBhsNDMi76LTRiI0kiaVoaBbkRj
kmWXry9OpAU4eIhut6pd1R/UkotD8u65tH1+ITVgZOCcupDmjO0KJROw+xW+ynI6
x57o5/IcgJ2tIMm9QVJSSm7tOhhyMMcg1ZQVPDIVlLGBbSkQMG+z3PxdnT+B/Asa
SU5Bwrk5T3vkRKI6f/2BILY02+ACkALrfldaARXjSIbvoV2d+GNiiT/Ru2IH6vWl
G0e6f8zLWBXN7TFKj/ZmZx1KH3vIA0yevTCnYRML1r1lm2Wdp70o7jH5qv8D+lyr
ou9/nGxr4boeoSo+2mr+WdYz3ihucZNfuV47etPh5M+bRuNDy+kZkd50XbRBYPNV
7LIj/mkc/EYEXatUQa/U+zZXOYWwFAtnpY3BMcgkqH5UkshL5rQfoQ4yY3FIVFux
ch0NiVaWwN8H7pjiG8p1to4cn8eqi1ZuFNywaBIIoa71ALVHn8aAkCyeHYKcqXME
cf8iKWaFMNWGEA9WuSkSLbKzo/q6jdykIldX2sARamUzwiXPw0kcq49KFqQ3jjdm
tTWTXyvenphQ06+G89ij3S9/h3hTci6kkOKREGXGv3uCNC2Qp/zLPDfrFpus89TA
qWyAh2jE3Xe7ff6fI4dFGNDNBkkGTz4957Kymd8GbjGS056js8z7MjlIoj5QaORf
k3WKP3IEAHgZP/Z+l6Y+cPZfP08qW0sJWI6AAUjjiv/u71X6FfNn7ZFCTNRHiTuY
uMmAmchQIWD8qAeJcW7bRvO0B0jm+RP1Lamksyr3aPyLhAPbOp7eCXJKzOPUtxgX
7agbWTmCM3nd+McUKasmCqxEjKr/pEVpPq5OmH3f/3cdvxb8yyX9mtRIK4B8kdAy
9MCvl+zTYjHNfiHpeBzz2Hu9JBC/7mwUr5K96Y7aOmSrqYsMOttNbEN2pDr/p7Ai
yFny5wzLNLPcMbU73sB5paQ2EnnQyNwgamfdF4o8REEL2oxjIQX3I4xGBdM5pRXP
kmIpIm7emKsiDNJdAlXXBKeBERbRLcwKSTAWvZAoOSMOp54XAgP3wmzvRSmTJ263
esNigR44vXTpQVaCOdGSFAf9TMxMiGka/8Ey5jFuEMYj2b23MhWpwQdzcCHnTJNz
yR8u6O6fymw8Bdv7EP3tdsvv/CZmw6XOQQX+dD7WMyHW8sv/b/kI7FIiuW4ERMkk
euhCGMmg57ei2rp171n+uIaxbc7n6jLLh+nv8q3I8l6pX+sCE2SAhcBT5wI7cZiV
/UuPkIsV6iuVQeyWNiMIRrxcuSLpdFwl1kcnfvOgSnA+Zc4KmV/AeFO148FyUo0z
0IdlZAGfFV2JZ78danppW4J0fS3eup55ZwSmOXAzrjn7eNBuhEI9aZPso5FZ3z1m
rh6pYwQPyM6Jfo2ugmdr7uJklL6RtF8cvszLQPQgRW1B2Nx2y21B6AcFxPsrWYBW
nKvfP0WBLqduWhBaZ4bpgiLIr4TCReKaZ/dumaqvP0pqah/umWIjUQ8nPQqiHJ9k
xY8w4FH5ralvWbqgDuUYp8UAQYvwBVpQu3a5tfbM/8LP070diaHuIjfyoUbsLrbV
nbRqTLCVw20djkzj4fH69CYTDeZD5HMKmop9lWt9DKcrNYw3WYvr7cI0m9Uhmo5T
AZFoPbzZuZnXeiiV4nCKiAFl4W2COCRInaYXSylIBBGmCF0CPrJyVZfUu7I7Dabt
uopRFRfRf68/b3egcsR9pYVghnNe3eo/lE48UcHEPV0MsU+8TZmmf8+/aXQ4Lxsm
IZQe05twPPTK5A5pcTJ97NdXAvzZtcSAy0dSFWqUGGjTZwkU3Giq+al6BeTrc6c7
HLimcUKdnlQ69t2qkj0VB3QrLZ1tRQP4L0oArPGLagdSRfVLtLYiAlPcH98KMu+k
TA3nSlFXkP9QFdwu5Qfu0ce994Ov7dxfcZLzaOuCc2sIluzC2V/s90aZJRM8LeWC
aV7b+cXO+bGj32FWoPwB6UFmzVqbLomJeNgWtw+jBMKIxUj53DKJvggJqxtCIooJ
LuJwgAdl8ZXKHpr6e9rjkjEKNmYAcL7IwUHt21iwFnrfqOSuimnqB0MQnw0rhjGB
gNgWZF5drEiSejlt24mtTe58cW3XK0eN8dhHSUUfaq4YOFh5DLkKHC5rU/EsY5BN
bSjbszShp3CJkmtucJSy6SCLjlkK/taVIaSMxoASHWKUR/oHdfOD6PuWP0qpjlJi
oTHfkccKxFVVlU4Nm94758rZKoguCrJmpliDBbb8e4zhRwzQNonnXUI2voe6kvbe
krV3r3vCvRYxfm0ucF2vIixXa5Urr1WebBNc9TY/X+mygp4HJW06kRs3OkE6KLVe
PNXTvVG5DKxMxBaxn4FvAVmWbP04DPB1URQ389hdv3ixxGIgStkoO6yG2thnSbhq
iHdhq72+bwTJdVjt4eT1m3La7BwdZegkqOVjgAyS/wcqVxskHpeKDq1QfT+STsHG
HN2O8dGwRoGX3x+yaiv0xCfgVz7cNvyOaRoT19VhXRVc05Ga14YWmaJMiP8ZYrN5
2jbOVJYIflLqcl5kn8oE9QO0ionG3VE83Ce6cUiM+eI5V2OiwfLOFcYQ2DxDCdzX
+OlJzR3ZL3gGzuvDj3/HTtL2NW2HQ/QsGUZs0Wrcehj3VP7EXDMNxxd4TDbYoyiF
zxLymqkjJjRNpQLzc8HxTQp+q3ZIwed2i2giEVA1+z96reZQeBnIaVgmg2VXmCx+
xBKFGqmD298ad4/4k40vPtk5IWEVkFBZTw6Kfznv4lvCmOoeKS96j7K7Khc1k5T6
pVp0b01FUNyU9Wwc/ZvM54lH6601bJ4px6LvTxQpnVTgYfsqz1SXCyzKU8xUf1+O
ETWI1ODQxP1PsSJAUjuPyu8UH2zSHl4wL7Fij8YHF41DQQTFXaoBusJj2Q+zMfAb
AcWoeR6DusbXMLNyj3c8WWQ5EdiNN0x7l74dYToExH85MMicm8gFn7bk9Dt4KMwy
MydD6GtE7zsxB+LwG7k3cUd42nj4fdAMb6s/CHeH9PVStELnMsSWPyLrtrJIBeKX
nC47juHbVjUonF1zhHZRroac5NLSupEs/nWKRiu6NPXsU7+XWIsU1DQ/zSK2nMmj
mxURdScAagQMO8hMdusNMgIFN46dd6U1UvwarcaGbKfrm9GBDO+u3bG8ZpUCwWDB
vOUvvaWZKSoyKfjbJw+2zZwO77A7K3j4jVvneqBsvxd3ZjLDZYNbgEjAfVWlSJP2
CXRBI4VvbGgMBwriXrV4sYJtA5U6glhj+N+XXGDI2CtK0MIvyuiV8bjkKlAQ//BC
VQEi0koSOdPXRYogZf034/pUEQbQNBe9g8b+cnkGrKyJs5GVEpHIW4XfEZVH2Y6/
o0QShKwUPlw6pj+GG1+BFh4JNi0NdF5s//8fPbA13n9sVp4pCf0OCdPak2wE3M8G
ZBxRTkO/7uIeFlmmVGMXA3MsGBkkm4OR1N9sZWEQNYkcRY9Sblw93/BF9NFdr/zI
SuOt+OlG2346+jJl0LTOMgWIVOFLs0vyBrly5T03c2yXtf9RAZh7xAdgG4CW3LgL
ECw1j3PcGW1MGXsc20D9N7v94NXtYUSEd5mSza1JFA/OUA7b3aEDydc+aYZYo08T
K+o5KDcIdQCw/z//ZDUnuCYIWO43Jl/kAvm3mi/ENysZhg4utQAvBKX52Mwmo4KB
XRCkTLX/G+IXKVZF5szXcI5dbWJy2xhVB0wr8GhGfObgu4kq8D7brsNs4LmOf65x
ildcB0jGenW/qJAH/mYctG9esLgQODe4ufNwrbeTbV/pDk1Jch7M/COMhLO+TdpF
udlIXOT47jW9qGByGRNsN0s3MQj2wVkmkvzS7PYJCB1Ot7XxLOVDgtTVNnfgIEhr
gPtQD5kQjDB07367h3uC/4Gb2OQl2yLZFYwdyrij7pyDgJnH2mbTK9ZgC85zm8Vk
SMZ0ZMAgEb9nAhtIhBJEnGr7qtgXLruPIJJF9gtoTXjYroJvdZ+QH7fCTmt7gNOS
04nRWJdhKLNso1aubpP8GrXhb5Mw09FeFTg6DL/ZSUDhWVTRmg/mk9kEa/vlYUNK
BL+RFVQhG+qVQnqOjf8SzHrTrodPAYVMjS6UJsRx8kHZxUfnT3ZX1kD/8VG/KEni
kCqk6rLC00uAt7QP/TPouZGSGghxulEvLFPvd2YsxvCEYvrBXJWMJ/dC8eNh+Djz
BoCNcFNERV/9zwszvoAEnf0+Hok6QL6hVBk/FcKhCsHC/T2MuyiXEMmoenbvup6C
kXLGX1LMKnPqnebAEyAm7WFhoBEKCulrrt74q0yiEuQcBRlbqvIQ7USbowqJXaYz
iQze+CslIFD6C5ahlJBIi2ml52ZXS2PbWgG7zz0jHIU3mP4gtotjCpQgVmMvtIoD
ynmnZxekxwGvTq58AvAqyHirygy8xWBtbe9lrZm3UHkjMZWgkY4LAL+m2Yf1qc6s
3eH7vc6Q/Cy1GBwHlmGTtcLF14iBhZu8jfxS0o30GN4+0RU2fCWXIhLA8bCXUIwk
+yio/DTXkoh3Awt5Qd+OJsZlnxvUt4Gldf73L1/8ADF0T6vuUX1zH9xtTcZrIQdS
0biGnd+vpTQTCAY7gpip/gHNYj8sdvIZ8lSVE7XUA7dE6oHs29LCztV/6TLx5nj7
yiV1FAatic6kQrULm9MaI7xr2iGPzXhWvijvSLl5VUPWyPqNmxcVpy3WHr5SLaij
3/arixEhwNWm6wd6oPqq3nHIGkcicTiK0iu+FZSw8A+fqiHi6d+GKNA3pOsnpmHo
q0+uhx90L2PlvtpZwaht/gpkwFhQt+CKynpZ1DbqLJye76fcQFJHqyIofdMSjYnz
xlNVshrCYgZeun2tQ6Znd14Hjph8t3qAB7ZIcg/YWDmFQKhb5W5WW25sRsy5b92U
5QXVlq52tHUCOsqOLIEpwJJmDH10a7QGUNPTxXX/Qcqwp2rvo7hwqRK3iChLqo4F
luMLfG3uU4vhdSd7W4rxGrVJsdsyLF6jxa32oYtRC+ZwniXdMre4ZDbGFAd1kfpC
oXNGIYji3YNdxcuLIapS+qgU9QZuYw4J7CYRV9Nw/tcjdhC0DieMklYWkbb7oaE6
V7Ctijfjwh1BkRDkaZvL3OdxYuwS2PsKGXATQhv0nc+4ZfxRU/t17GVbU/Cnmq/t
ZoDhs5mWiaAEvU5hTM6XwaPd6DohOYxyI216TyA012siOJ0cVq9alCztSAQ81WLq
47BPsqRVcX8LnD0967Y5TNu5W1dzGF3bALV7gEVjD7sVqLUwbmZci1lbuyw7GnjR
Lq84gGA2fe7Rkm22g1tyPwAkifuIsOhkO6hqwBAeZY5FqYtjhuAW2eHNVRy8RAX3
ouNth8s11NIpdU2z9jz4zpNye1TJyP7b5J+xRTuGnDQ6xVvdxVf7Y9S2vDIMSP0X
SGdf1+TGovw5JAMDk0fRbYwSZ/9osuqZzsREs/IbrbPLmeqIaoFjIQJoVyq6rqNL
qPHy3WItdhy4KHHkWZTPdBppYDITC5QfUQ3PzNVvCDmZgJwqKSkzVz24QXIkqRQV
77Hl+mnDO7CdnOSQ0Zpkqp+9oRDONnVnpUELifxYqo4saewgvBjQywU2cy/hxIJp
cCayt5Mw+iZ6v8/AymBstVWGCAg9Bz71zRS0VMZoZ+md6LlsYYJjXAAzjDGaRjXe
y3LCOaHFMJI1tW1C32ilpdotndjvEOxVnlLwNqSbzxF4EWgp3AtWLM+CsF3gPeiQ
UVnl5nrVUN1M+VBX1aAJLrBzA1k0dEW4U+oZtti961bhAjid7MbRgj0+pqj7U+AI
vFYOyr+qtc/8n5UmHvlfZJ1KgvJiQwAKz18mnJE8eADxz7KGtZxjBzaHiS1OXtb7
4kb+5SC/cUAyp39KmJT5zMvF8YeBGmEGlSoVlybDCp6JJtVEFwpX+eYrisoRaOUj
SXLQWdtofOEYOUwA7QW3cYvlmJZfsdCQ3CQU/I68P22iikrc3Ojx8Una0MIRGOIl
zLIszLXf6fvsVUgcTKGEtz6+c10xcsBEGq/ghV8/UwhetX06UaJX02pmxCfYY6Yz
6l3EKMQlzJSlQSn9NWqn0qpuMjfzO/JdJFhK4vaT0/7cidwXl5YnU9Dmi5xDo1eB
j0Qw7SCDj8sDU1bSdWMM4idNz6FIjxkdt+pkJdqdnpQZ534ufvhp6PaIDkNmHSfJ
lSEgK9fPn0P2atM/pzvcejt/Yj/AUS/030mz3xiy1RyXRUtqiJ24oWf1Vck8uPeG
Y7lKIRYDPxdEGWOlfUpQ+fqXs7K8QgOe1XuY8Db8SnzArglifiZvh4HC0RQignJx
xL8Em0KeJ2ZCvx8o8FxC+hnln4IvWp964HAVZmy/IA3TFrU44fFSDGXPwJWSoYZx
mLOwnB5cZEtk1ApawKQL56v+w7vgn8emAyA2UFVXU7rDRYw7QmvLk5McSawxFSnK
IZbfN92CHAOG5ydjV8/dOrdlcKUcEw24o/gsb0ILx71jBYX0j6hwB2aNFN5yKR6K
KEyB+f5luGyCsgakJJ9YxcEHDFMSrLy116FBBGO5ncPPyi3FXt2pgHcFezMoovxr
74nDcpbdqn/L5eEM9GZPQoBMC+0CmLbnxYaBXPKNH61V2eB3/uwtRKWSFiEE12sr
YE4IktvOBClth3+NfXMFDPDtOZUm/VNF+jOc6DD2dx+DweNCuTI1x8pczIEKkU1W
5lgE/ADgLo+n3P5pzCMIxf/1mmNW77RJ+2zDyMcuYgaMtJYAV74nI0HbjOT06ao0
nfXzYaaT07lLtHWa7eLgUr+DmiVzu7eJ2n1U4NpgAHrVHNhHOt5y4v6c5STea0IQ
qhd9WfDUlBkSdV7lvwrP/Ck604hSD5qD85Imiyqbuk4KQiW9nOcJkVKkWsFW6ArG
l3vSr5MjXZnYPaeUsIYNjjrCQ94QKWZEddMgJypxHrur0n+nfWUnm4Tl+GEh71Da
jNiWiVKmnGWe6DUXtrBq00uc/AcaFEnDVW51e3R5KVe8A2PBk+4RWL45d4HKkpzV
W4c76bfIvNcdofJpffOQ6luDNFDC0qhEKrjDAnF5X8D8uiyRf1NHJzt98JhygHu9
U9aWmMxraX8bB4USVm+9sf5UAM3Hxy9hgT8mOxBOIAGbeegdOje7QVcuRV83bDiK
CIk5bw0ahoVQypdTEsSuzgrMW65mKdWOYroaFultn9Rw3pHb62hs87zVGwbI6NpH
JS3eDKPk1YSyIERdGT1HkYMjNQw8fIyvLNHtne9mhD6/4q4bm9Uxffdo+kYw/3TD
dcu0k1/3YuQoGCPUHonBMCnQTIH3K1jJkhyB8Px0YFZBXqxP2ZVpXDlzhXEdugu5
C2Z6zFj3zccLF8eFlWsOjie8Ime5h0PCvJLM5saA2+CiI1h7ihc1hHdOxIYS4IUI
zIW1xII4jlgJbFpayGeQUV5JjYmz8si/f80tRegfgrUgenJb0E6h569mwXkmmHNO
4b/71P3t9qsfuJLtGtLKNMdAof5M4xQfmBbJ7yORHzp7uq1ZtxOlW5GJCmyCSaey
nvF/m+t8KyQRfhBHTr+5MdwkFbNp/3TKLvX+3yX5uW+s5iBMGpPcOgn9hb5nVos6
vbxM+fpN0nkiFB5shYsbwV4JLtJNo4RAEfZ1d/iYKetTl7SifI0ysPCp94nHc37q
/hfkJps9c39ewx9Pdc9UdlKkU795Sl+H5msBYTrCoVmdMe8o84GRtoQ1zbihdzeo
AvP0UzJ+M0MhhjPJKPOpI4pGAXGPB4u1EV+GSRYRALCXv+/FXqShTNo3pDLSggHY
+21abA+bgIQZXKx9iMLu4n+sQx+avqGi2D19nk8uCSp+UmWtjeNcn8BS+wOIn78P
ldIZR5/Lrm2g7fMIiAr0wQlXIsistX8dIXXSa4UkIeoIMKAi3RR6TujMgJOxaGHC
7Vl48vSKyBRDZjhjtFC6mvqEen+NP+3LOVByMwMwTPMV88ATEbc/BjfvohFlybxo
sSJljeuOi9gmdn61FiC+7ICi0s5xPH+zeLnNvk5Rd69lHXWRjhN38XJx2N97ADGh
fMthnR+tvYwWGa3rzV6T+q2yGmdA9Nl5Oiwdy295PbCcn4QUycIxNu2cK1RfY9RP
paryqnZk9+hg6YirlQeRChEuNUWItikgo8L4T+rGEvYZTwqCVdCN+6KyzSh2ymPh
ZTe7MTj6LiJZ5lVVO/5nU4nfwE4wmWOE74/mYVLRduHjALSeCIOuqVP/M/u5XooO
2keEVJ6FwUrbZAA5wgTgDp9HIu6GpGK726dMq0Wb8Vc7RkjTSjf8KNaigX7Ihss6
l8+ysikj1sYl9khY4qWcEPWwkvYtAHYW2UAO0dL4kXtWhnCe7rIcxRb+2DqP7jaq
7ClbhG91SePhPTckAVFn9s0xG4ZASdj6kwkGTNYGtPqrKZXP6V0ToTy4317TRZkN
p62MKvlvdc/bKg1EEIb9sd6IbxW++tuOrtSMriHRQv+MzfAvpeXvdSoZ99bnTgve
Yd6EYWZJ52O2gtPb9//O+m62Xpjau3urs2qr16537/KiB7NqiuOkUpw3nL/p5sXt
mnAoVhQfGYdqYjaiEmYy8zWzOUNyq5jLeVKPiADqM/PJ8ALJF1rcEEQ51wQ3OZpf
Jv6bPtbqre/TgLB5xqkiHB1URDheF2ZFBJ3dmrwTWEUaH4WGtdhAZoICD93oUgx7
uxM2d1HQzQGkgVsPLmorWDVRDnw5tgOKdyUeDX24NIlintuYaU8J9JWu7izr2dYl
PiMjz/Z60Mr8waxlmKjISE5Bsle2YFYVem8wxzGgN77/d5fNkbB9inLGGFyM7qIq
I14FW6piYQGyOOxxtBD2pS+C9RGOmeK5/ctSl18kY+O8Ns5affjEfNwi3eLNVm9J
9NjwWoWeQRRpbbXKMXoQg2hDAtGL1qDbxcVE39X0i3SRIK8g4QSrvQCkk+0W6OZm
7wxLd35Bs0hASnzqK3HZtLsbCHXZ2A9ZpVXt9Z9ZSJRzOX9nPkB2PtPj3JcRcKZp
UMHR2q6/duc8bbNuN6GHT3oSgGe4ugXmH4x9f7aDoyYS/kNVaHOa+3t5JRduWDR4
eu/fR2WS7WqqwQCGjG7H3SpLn1pevX68LDNoOtwaRbXaKY7aCCf/5Ex7Z57BsaoY
BxSFSzMkNkwrWsWC1F9DZgJ/94YjkU80JNR69qAgVuruNEbnWODf3kibiH8MVv58
Glaxsx/+VZd1pALwiuJwB5Cwo5M6AmgCWKtrSL1ASokaHrQOAd9nU2/gCU/eUw4q
F2AaNTmlsjlP4CREhnxrg6rfQ30BFCyqPWhFLrcFDmGVvvE/XbQdckNjifLtJpsE
dIVp8NO0p3qPyDiUUPaK/LxF43berQM7xkluuftGdiUC449MUB/nb/kpKcvUra6B
wkOAFgex2jr6PS7V1N2of7CNvikZeDB3wVlGeCXDonhdWOk4TJ+g3PmHX3Czb2JZ
f+SoW4GYMilSsU8YlVb85tJfNL2XsYP7kG1ZnYUVy8+4t76JLrxN4Cc2rRdD3mgz
WiO0Tif+3LvP8FEIdNl+9N7Xt4k2Agh9f6nFAHLRZrF6Of5ndgaShyFPsdnIbAIV
mOCL37Kb92XDKoLa202tKn+JUILWpR1TJ0npVyfucfah9L7WPKCkSC+biI93yDL+
BxyGi6IsaqhMB37gzvtD5SocaLnk/cxcxojDTTB94fu6La0wxXpV3kKd8M75Ibvo
ZiONXht4JEqqojn3HxjpK0O39549ZpujXKT5tc/HK0yHeS9g9LigErAsaPZiyOxp
UezfsAJfepPekGIxo9Uk5hvwhZSEJWx/t9V2Oq9JfMh7Gtjx+YgoBJTZKpLNS8pK
qgTgrMLkK/svGjhaagIckqrAJ1CtUfeQFXVSGvHcJ2SKRC4O9EpeZcJoYa+xtJjf
LOexCn/m54HuvqjZixl+BWObJaIY0DyX1+AEqbB76ar5Vo5vb3vn8oBvrU0XYb+W
Jjv+WhooZ5k1YcdwBsKQAH7RBV6RNvhs6smyHjgOz1jCWbzZlUuXhM8foz1di+UD
PHo0DkUQMgji4wsz15FPr/a4F3KO2Wu22thsZ4nYZCiToPYbdEIR0VIKfVUyST06
CU4/PPbnSFtrx6OaXHo6F6OLhleOkjJOwbHJ/ZrIUN9DFXjmoiY1VhA/21UAAy+h
VBma7YPPlMTvuh/hFihc+G1NrLRY8Ab31EJw9ZNoV7Waun4J1AIMgUDK0DbH+EGK
xi6m7V5N3zG4KXa7xL8d+KJikPJvLfPOOYYG8eZ1khq1D6ld/zIocTG5evt4derP
RsHNThvQGr8Xmoz6Vbmny2PrLi190TvebuOoiUOAhBTy3dd+DUJQqLZ/Du1osuTJ
vwHXCf/NqYAL8DxSIvStUjty5Cw9ZbHeXWMy5yTQ7GLuzUGtcf4ZH/bFKqyromrj
0/RuFjBTFdcaYH7OdpHWGPPxuaapy3AClZsl/HY1RIgXDdGWPDQexUuzRDfSh09P
XeEsGETicVv3S7JOa+PJsEe1ANW6RIbpfx22XkdO/GU78GYB6MMQb4QFWphTmiEU
L2seU8J5V9OQFfqP9/A8pKnAWaC30ySptgTP/qHwpX5g7EGj3oC9TRsv+BmyqQE9
3eFkxzGBZoGj6/Cv8QAPBhrVgE9piqmzqjNFIdMXqEG4aCbVDJQOHQU/IF8ljLwp
F3Lt1i8uxmmy/lhOnxcvK538gomJZtU3oEIamhNe2hfKHOINIhA4cBIlg7lGYJAv
wS8eEHqBDJvX7ZoqJ9bYtgfsGE1A63V25n8t3HlhRQSHfdwxPpMrYLDEkYPvIJsI
ssfa/90esbwsl1j15/63jf2cWIrzBmDWMX1sPI9A/lnRUL8RMnefgikRfvDkrVit
+CPtdlMjrZdJZnhoXulfYG3JWjJAhZ75hqNqH8FLgH+iAQ/NbP7cp8+nUw4RGRlM
Oy/Ulk23JD7VxlBrnj1Dg1oP8wuFoxhHSzatO2F1mqeCwwr9Aji4lqI/nBZdayga
ID5A45Pz3MNbV7WCYyzCOiZ4SafmkskTTGK+0RdKoD786zyUj28Xrd3DaF+uFci7
sBd6YvqEHNsEr/8EEO9sF5nRU7E2Fe0k+HeM9IwRY6GZPBDRUByOU8x3bVWQIybU
nuRKEZDb9qJV5mYfs96qvqfZ8JWOPvaYBijBDSsBLnj6rCGZm+BoZ7+v6qtIEp+p
cZByf/2cIlbrK2CTwbKogglXMk5ZAyYxtDVK6ruHfZ406xCbn5qOE93pgGagKqe0
A8gShBk6iS8c4tpUDuRYhct0LTlExjr/iZHyfR0TYIZTOVVjmoF31vGfEdf7GwlX
gOn2USfHD8js2NvIRKumkqtIfkiWoROkDvjUBDrQK0Y1L/t/AMSWshbtnhBjvMFe
HDA/jvO53w7LRfajIOeWYgxgNeo7zDRM88EAV8HfmaOZlO154WdhIsmUGkVkGYXg
VH/MHaxVxMGMEh7o9s4vtVArhndi1wMZHbInrNexnn+mNk3CL3XeYH7jmHTDcNiX
kULTrcxGFP904crnFqNyDmZC9r7EBKxO7xWqqxuRQNMT8hw+xS8zs/FFrG4siHl/
8PqjzdCFer3izMX/1KN4eoHeMgjY2u800OBmxPvxGBB6LnJkvzOfrkpRQEWweefv
y52q8o1JsBJWItR8a1+bu7F2XWilvv0pM+6onIIU13W5De0xeco2iZW6c+RZZo+/
OkGeBdQ61g2kUAjSzLlJY/Z7L1wW58I1shu7S3/dpCmzP6CW1NjVaPB/SRx8sfwr
itrnD9SlxcpHhTRMejkU6lr0Bj1HU0gAd98j+OGYpI9jVFuUE7Itwch6PNRTUBBX
Ermu4NVyEJ8BJ9mhpBaOgi+5acdvmUdTGjKAkx25duh75ohiM43hTwhRrDAxkc8+
/jWLrXXOztets0kDP8La/xEEj+w2VtQJD8xfiUE86/mZb/JjXuqAlGANjwz2VGL3
T0sZ8HC93o7pSV/EAFSmNmOTtr1zW5tc+CQsZOnJCzAvPXberinW8S76vWDTluIP
hIBCoobYdlXPxgaA/pmrRzwaC4uzGKouI2gejbHDTferMtezmD+871yy5Uv1v/WH
6wCx3NBMdoaGLM5M1I4MLxtKrIbcBSUGpmIPDywzHD2yK9MMV67a7EqkeSC9a2IK
hkUNopl/RgMS2ukT6+rQlNX9RUYhHv1PE269kh1wYN8b1PpQGIrTk+YMSKygae+f
gvz+9RjBkT1sUrV5dVsw9xag/trdRfC7JyX2VmtwVGvXPEBAGYlKbd5RWdsHbXPs
0qwHPQM0ECmfuIiIhcGUzpoVMaoUPG6xenoFFqgZhmCKVRQatBCavZiZwBgbLbD5
dvwAK2C2yElQ+e8WZqIZuGi6jI7sHYo+nFfhamSgXFmmAWePZ3bkZEWY29a2FRcX
L16ysahTUX8ySxcOWOqPFay2o+z2V7E7jd2LUv1dTyxJgX1Y3IHxageu5YinTjW7
VcQTVsHTRdfhJLxIflJ/RaChPvbsGhnaLCcuVpSDW+m5WtoX4txd7Ptbya2iBcS3
D3QW4LYI1rXqrgbIeh5QT5mT+M24r7LSWundqfnvOU+YXiinaSTOndCbMXeV6Wuq
2Hs8RqDzPVvDdTNe+WOWX9vcIBWvhMnfna3eSeJ61lDFlnLS4jI3yGA9h8KiyeAG
djW/Bqz8BO+JkJ4IGlNInYreo65PRw2SMeegkI/m7adj609z4rU2haY3PBrJ+tam
mEnlK7EdP8OsgIagYTBPod0YazsbUNHMeMlJqbuFI3zTCe+hu0ryxhYIXCXP7i/v
sPmdje3KdwlgQXW284eNb1VRafMEy1kYT7lwLOUe7ke+ufYJOacyE2wXcPIjlMNX
K8xDoRaveK1fxhjFFoh2nzUGWu4S3a6smoyDMaGiIjw1lbPfrugMkQaBvH5vc+9+
Qz8961z+tSeSZhR7OcvMUldxEKKenSRY/cB42xkzzm9H9GAa4tzvIpiWoSa6zkT9
KWzEplvvDO2Re+VYLdbREItJqW2n0SFQcLRAY2Im+v0z9ZU0/EZyTDn9cgnUWS3g
9hlY1y5gg3DKMAFHD3/x7Ag1ba18WvmEug8RSRBLZ8iFFxxVaRw9OVej8hQ+oH9m
LhbBXbxyg3q299QfH8uxAwtttwoYlBGNX/oBq5+7p8Osi0wfJVu+B2WfTeovhAS8
QZsjdaEWLo6JN7jHOdEjQE/bxzPudkursZrGh5+rpj2/ZrxODs4tsTAflOuQlLGC
/118y3b7KFJcbJYOTEOGB7SlHNTyK5oGV3/rHdTug3ZG+QLcOq5YIbQUw4RNTftk
ron5CaavXIMoKTLxWTta9C8K/InXv1KiBM7xzqKbFyL0Xb28mTfd5127X6R83ZE3
O4hkXyAFDMbkHEOXLXV5sQkkZjT3L6i2/qUkvAxUpUXx01F0elu8pbHd3fxCY+4E
1c/wObiO14VX6i9E5ICB34IbkpoCRbrsK2lgwXIZfaT34AJaxiUF941NHTqNRF2E
hLqyXIfjPvPf4fq3l08p2MYUbAdhPjvwvu2CIURd+Ng24muDvwzR/oSfD7mDDEZF
T9c9t6H2wEcc54k0sWjbBy4dGaq9xIdIIF7SFXIU8TCejsQe2JY/lf3+DxzNMqkL
2B8i+b8ZjWxOprOUE59g+VfWj1lp3xL1cI4+UpErkExVPEZD/K5mrqGaPgacUMgR
CUNs+BV+mR2YAge4n38yiJljEitHZA2CrGOzJsrm4doxnslMjFxgZEkzCwQPxvcl
QUDGlowOQltt3q84/9PmB0XpQlaBT6zck4jb11Pei/hcONW7l7i3g//Om+cyYH6F
DydoOIxRTUAVginZ1YDfyo5Z3TYbLMLugvcna2r6OjHyRjYx8l1haJ1wLXCnePqx
OrGvfd3uQZs8ITKKoUFO10gZ94AHwDsRgBAJLRxh9CW9qnfowJV6kmDrdhMvnRYf
l5qb4ftIVXzbZvveLO46RSxnQzSIDqc+Fa4SRbxOxajoDeAZzyqvdhcS8WBIvOfa
OHYDsp8sQQEezs+qOcsM9A+3tCF3n1WAwTwx8OBZ2B/MCg1W8m62a82pZ9yl8Vqh
9I79gx/Hn4Aot1LeTbPMwGc1D5YlQmQ86zV4fhvxnitTtkQUD3fSQkx+PV0+tLpF
M1rKa4qkqfoMx/W89ytdax/GRDTsPQdUfFlM7VTFk1rEgDclHtW/LPny8oIY+EvH
Sb4vkWKjsP7Ys8+qPIC+rY7Lltfq8+zZGMaFG5toJ+3gf1DFmOwkJ0RAEKyxJOWU
7TI8UHf1BSdTbVxj06guld4eSzzx9JWve1z1RqgaJ5s96c0W+tMHMexIRz07zzJw
6Ghz9IkO+aFYOh6NfkQYdB33yMC1MjMOzTVZqfOR3Q7mMf7OLPx3lDtMbrut2LhO
eK2890pFfgeVbKaRXAzfTSqM9O7rykx5BTZFe2wTgxuIqxHxbN7j83iwKQEp/TVx
KYuuK4PL1YMPnJWs+xwCfXl9VFnJ0LGfoegHMBgJFDz1NlpqZaA/Hjd2AsNuAZWA
MCiY6ZX2uMLSI6haPRx10O8FlW4oN9alzZpMbQbbFHY+ba5IesLzm9yz7B9Qo5/Y
uPB+AREaUypqNwNbPzHzRr6dEOFaZqhl0sJI/wNfoXKwX02sMnBvc7v30nI5OV8+
+RGIo+m7DoHeAw39iwG9/WBY6GfmKShqyHglEd6dJdY0FsFlAhQYx9PV/aA+HBKj
JqrNg7ZFhbb6eVV6aw2ydIApU/cQTY3giYx+v27JtIwh6a/YYGtcIqRzUjQ5ngxw
bm1V1QZvomSBeAZyMPIMRlFiqguPf8NZH9Ir1Ba6QmhBTWkfs0sdt3JZtYprn9AH
wYcK5QOa4sc5KzT0Gs8zBYQnRGqSGwV4Rur671LKibpUrnfqGtrEnJJHViBSY3Ui
Tdi902lpx9Jk8IB2RIw4UeDQZUxqMa9UZxL77GuNS+iOyGgZVtaP2zVeSCI960Na
PFij/+hnFJkCCmcRRjbqUfzTtQpFRXPqDyJzJbnA2gEQomlBWmf2p4DCsymotOPu
pCbkfG6CWHE9XIPdUdTqtP4EJd87Momiz16escJJZJ6gjvn6uaeSjzlzNXXBO8oq
Xj5dBsTvpgpCT69Emkzjl5VbWMwsMvK2/Jm4Uy4Vl9qHgVJrK01Kay2GcBinxcQ5
V7pD1oER51yLQnVFWU5/Ml1TYjaaHQ0Dv9QsqM9PQldBEjpR+8lOdq1XLPxCfYb/
jkypf0XiDZD9Ta/9kYtcCV16wWR5E5zX+b3fm1x23SI7njuCj9fJNJGR31wqgt+j
5HcSPq4mFcZZe1lyTVADl7M3R36b3J0LiqaEG+oF8WW6jGPlJqJHdzkkdIa6oE8U
ZaimTZZCLcOysy3oCVZPKzEd37JuLCJOF7DpsTC5ZaErllhDyyCIWAE4tO/SJu4e
VcBCfNq4u+1gMMbwsUMJly0tJbCIIVIZ/EsnCgQobJrsFy1iHELXSQnaiStU1gFM
qdy2tHsW47aRYLRAmsvXKSWeflcgK4rh+Gxs96ILW6si7TKJhb0zIVEbkQvEDAKy
Fmfq80VHsFx4XjbrG5WjdthojQdgRGimY5fu+OjMTGsgMo+EWGcMAF+B4B6hUGPq
tHUzJqXaQyazhrTOUSDUb1D++k6zbzgA3BZObOKQiC+7ZA0T3vqyH8hHD35qH5JP
QU2sB3jQ6chBWPFjsZaJwhBbdc5b7H9vkCh827pGJWBIFBfPEBjghrSt+grFQ8tL
m6HiB0pTvU61DO+LoAM4GBarJOfOTltNq74XWsmFTPPowUEx4QiChaXoRqSGR4xM
H1GX2WLBVV+51J98wNTauHt/z9t240trqnz+XoVvUNk=
`protect END_PROTECTED
