`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FNkb9YNds1PdvJxObKABOmYF1XTJAahrwBrWnITqVn1wqPxCnat4ZK+SGC1NME72
c82M3ovh4HvqPOKjMIQAbXd6XvoRQaNNzeD4PVqEoMC9z5GrcIwHvzNybcPGiVnj
USAae2vzw4fbWzz5Xjp4oN6cKl3uiST0Px1LbUM6qGEvYIl3jVGTR2b00OeZ4Sw5
YLgDP9FNzq4MjlveZl8gnIBFIRANBX0UnIFlj8vwH0R61cWE1yWqlLxVO7qpRgaA
lbx7pA7QfIqeWvCIPVe/SESKISp4BGcaCeQUl4e+i8LakJNWNyj3AWoE1YpUdQ22
fim94bbyT09i2IPN5TMYoiQ6l4R3DXX1UONr6nyOPIHS3RRkrZFre7XiwwEaQsFr
avhpmuq2iTD31Kc4SWiHxTb1DYRLJTrFlVz1mn2LFKObAwXRjzZZH8mIaabkRA9p
Fo3Lh7h1dvVmgAKdawR9cRAmuN8gGvJIs9ORMPY6Q9YXYtD/5Z2LH5kfb1W0bBbq
ei3ChBtggqXumF8aDutulU+8dMOGWaP84lHce+PBEU7cQ1IihQ9rk6spvm8ybK1T
IQgU001upa2oQd7NKXKq+B/1USmBNDoWtKRXjtyOLk43wfBdRhf2tb4y+jtA3vT0
5jrosh39QhDliSHPscHZkTfl7twexCKdEYwH4crZICWC+F7r0Vfb+udzeYANYhw4
BE5LASZiagupckLAoxrtAzLqWP2fDPxOp7eNjVE86k0fLjNdd3ZpTUCWvN9rhHAx
dhPi4FPYYjwIR1Jl3ZcvDU74YCdOGQjGpaH1Dr0Hu/inoD4vGSPgED4jIskQiEU8
TfE3kNqLxIUPjSKLvvtZzmroCmIP5P61zDB2WvbvXxJUJok0ADl/FP3Wf+uOzmne
nHEt9BhMG3C4o8KkDWo2JxQh93RJsRUmJjV84rU/OwVhYeko5hRuMvercG5KhwvF
+0c1SzDCDk0lv0gaBaFyKdzcTwljbAb/xcsk+1svFS82aOURF/FoQ5D3em65N7vN
qd/79yOavGXw+7/pnXtDl4+pOml+jsABQHfNPjzg7BdsZc6PcUnMxW7XWWTMRRwj
EO+Gl63WOzK9EDMjrFBgMO82BbKO/+eVXbKclY+bdkvn1pWWXtMlR2iHLk1X2T0z
Lx5ZH47Ncqa2TmMeEXJuSTbggDsdTiiSNkUfvsi90NUcW5/ek5FtE33alVu40hpa
VhL7khx9g6D5cJQJovD64hzilQzIQCJRtrMwnLmpiow=
`protect END_PROTECTED
