`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jtROYT0ny4CdFUSjeIPV0aHlK105jMEPHHGj1FRsQIwtEZUNF4AZtIhsfTSi6yer
lR6INiaYzB3+GNkGSBbtKbK/PKNDBTvhSEWoWOHIUOiMMv4O5AyXBrZowOcrYp0l
l7QPkP/g8EAxJ/lYrKCqE1HUVZPVxhbu+OUh2fE4L/BQSO2eypvFpUw7gycwHkr9
ogSRrls45w2v7AXbLWoZJ5pLlpYdL0AcUefCYSuMaK1tjG1W2U8Bx4SsnEyFJfjJ
JTuy+ttdb8QaXlDiT9ho3bOZIdiBHMSVchZUeVnClC5bnqPbooJ7E8rxGSvSkJNm
+6TE9BiicR/wL40mfvqypJ0xL0K+NFv2zOEOu794ftYHahUl4cEnmIPR5Qq5cNKO
jSTZAdcpsVcEDXKhc7A8uEq30ETrF/H15XiHE8dmUdezNm3TMWu4wuBn1nGw+fHU
AL7089anGCnoQXMXxUvbM8IL0zANaMfD0fqKyQLgVIX0gtkHo4tw8qcDCmIFbVtr
sItY/7symBnAvh9cOL7PBStWBnEGOxcZNpU0kStEmHA7ZmqodiMiJpC4PhQEMhRG
bR1rwBAhh8dG4sisAr4zQAFJ1E7wSak6zfjrAw9sG+Al8yviA0upDPwOWOte49hy
jBTT1HKjC83/ktxxy5QO9lZJZCULeQIZIGYcLrTRUAV6h95xzyb1Xn54BLax5h7d
hno5Sr2UUx5iFXYzbdmSm3HdeIbiJmCwt9pVg3mWnOqOMmnoHt1Llronji3WIBty
3DlpiF3bsnWZNWHrZo7ramIPJudP/Gsc3r7zNZm9/RqZP+OYWKJyRwyalX+ghEjD
`protect END_PROTECTED
