`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fhsiXzV1t1/HBIQH+Bgapw+/M+qBcCUjbtaIMqL6yofCuBX3X5TeRiiFoBoxlS5V
R6JfI5YCPvOOtIlEkHZ3MpVh5q2SQQWTPhMVlJJ9xhOK+m11i4wPkmxVymlElFxx
9P74gH+CWYxrAiuXBX3ddeat6WKONFftRwPkOcEmqbPAnaQYP+Y1WuaqIUOYcb9+
fQTzPAF+AfoMjUJz7ILRidjH62O/d/izVRXTNY9aoq6615MAAO1il0ePmufSQeyY
EMaJLLhoWzBUetpEZN0UDgTSqklJ0xgIv8eyGjLGLUz1BvJX1pNMC9NaPYUYtglh
tKzKOiak5IjTbDuJxR06tofulH3x7UFD85aee47WzDFeU7rGyn72cqeU3tPPQ2aS
dE3z7E0aKMQEG8nTUZ5zkKq8D6KPo09gFFtbl82sjjIyMi/BMewiDzknrcllhb3V
eKqXmph4UtGf+E7AixqSy1pVmUOUaO2qREo2NLTXbtp/VPdfh27isZ38ZcgJ1GHS
9m6DhIea7XMPdpa0HDFUQgRGCidO/S8nX62ik34alulYhvjnX9R2y3M/j4N3uZqT
I6WZ48+ndf7ayhx/ITtyTYBim5op3ZwCczAgsMXD89W3qvewFibC+y9Xj+xxZ62p
zU7OpV6LER3Azu9f4dZC2GruvJBSwmcerzGz6KlTTqnaaBs0jTgzwplvbAjxvTQV
/dp1YR5/4B1pfWepngruWdGcEK52SOB6lUzTYGQuwoiLdIBEeXCnibYAdgWG1XPv
N/q3aAED1saPjzGb5i7geOw2vjyyDTIhXSOPxqrijLOmoYUto8Yjxjb6v4YpvjWw
`protect END_PROTECTED
