`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TxP0DeZzCVbpR7v0J329ZeJi/0lA6XxRnUxAE8feDvdTSrxB1zTVGGXHn6GFDxOX
fa6419EedD1x1V15FqwdnBOGwVcajAHN30GTP+jwxfK1W0oe9FI8WpRXJSurNFR4
yUbFxZn2HzMeS5ATf4j1uBVQygsjiYnaSbpBdqcXWXNZnWcbJvgl5qF3R1xcjNLc
9M01w974+PNEYO1jr0/2MpJS3H1mcEgkfnhPr/4uITHvCMCqffKMiSJscwudDK5G
hBqPfaYjLL7o5LFaOdf9DYUK8D/ONyQnF6TQE3bed9+pVq0tbmQWtVpGqpWk/m/M
hGYgxKY1yB56V3AFhOtGD58dUKqY1lcH/ddkp2GKDY9T/nArQxwfAfeT6piPg1Tb
hwJ1P8KS7Pwxo7/cKCenrq/SNcep6YpigZtkFHJW3HYByM56nxTxFZfNGj/EHxJQ
P7SnwVFyraQZjV/+DBzrnsij47/i+ADRJKdWm1kmcZBM4MUl3vhd1zjn6mjrtsmV
a1BsjBq47FHMHX0iJlieJ/MydwJb/Bl8bv6Cu1kGQqNY3BArUtABplC5sJN9eA0k
dR9IlhoGkTaAOLrtJQLBxAj17vQG+jR6UUHl6YzpGRUFL2o1IqC7q8PrzsKlopWZ
fZAzkcawlX18wcYOe73WViJjku85opIGu4fOeDEerJfsG195hXdEUmnp7+wwlJId
clAAdLrQdytQf6vODAEna8RgfiCkGYs5AF6FTHFrCJ//s2RXFkl19pl+ruCb4g5z
b8yqu5b78BBOTCdrzY5gfpsENMe+fpmlZsWrcRvEekPfZhYtM6Ahn/wcimRPN9Wg
aym2u2EcgvzHxDNNTLBGP8e1mbjtRE5q+nhReU3Yt04=
`protect END_PROTECTED
