`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2ExGN9MgreMDJTyOiyEt63goE3Z77kX6MuQyeaLaWTHXSTtoZ98UxBJFdpQl5eL/
5OCTYF64/XUDmdSkZFXbUb+myFrhrUTjd0pLJj+I0+jup8XbhCpCmDJ1XDmhkG+z
0rXximaz/1FDYraDuaHbY8GkAZbRz0G9u7X4w7764yusreeRqJ39AdAgIxS6nr7Q
VO2sFFh+qvjReNRjx6Bdz+8hpcXSx/qSBjmkZeG8pUW8lfKIos8o1IgpGodQeH2F
b5i/9N9/jSUBxwXiQ1O7OPkTshhB5R7NhQ2KbT2MCqPgcced9lWwyiVKmBV+FeZw
hhVDtVes7YjiIiSo/WxuhTJsRKsu9aF5BM5Ylke5nIcdfmhTj5GJaleGFyjlFTyt
VNO0V7UV6BPssfPE6DGX/Hhea2eFJjNzqNli8MWyMmcjDZi3HKxiRuwZxj+u1ikx
j6CUZbjfeu2IDv5ZJDM4clU5xMd7At4jbGndH4VSQwkZ/BGxk1MHA8hrmvh0Wb/n
8J8kmQ2z27mP5c30jzP1+f3cIKdEIAMMR2VNWQx9cl9vcZsXMfXezEGtXQ+H+dl+
b+QVpZteF2b7FywbAGJPN88S9mzXSHXx0j00A8BNWBhl9qOe51ml86gszpYIcjl9
QALvnxcf1SOEafkOkKf2QbCCrapTaavAB+68g3O2oGSAGDG+eatk6A21DzZCfUUk
+nvfAm1AK0HrKtOXVsuSULfViUyHsuKgehyj7SaXsqFin0IYo+rn2ZnMTBzClmeo
3m749sfSHx7L7OiIiMVkmw==
`protect END_PROTECTED
