`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hIMAikARhfj1c1dX5Ug3YQKViM3HOUPfOXoh0X5cbNerKraArcvQEewX8DtKFBrq
NRB9G/Ekx30Tl2VzdT4X0guemf5Ub9I6BQs1WRxAjkyKtoxQKp941DJan9gR9AYj
ybaHS4yLPRJ42pCoVmb4ae+3deF6T9vy84zwTERXOH4=
`protect END_PROTECTED
