`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j7iCFolf7jvufsjcdi2T5CxiQtiWsUAvDKw7ixi7t2Qu3KaWreiPD5eJJ0OUagZx
hIKsGbTCNLfb0D64AZ0335KGI1nqGSLXh7gakF5aB/BT/nMF3rRc9b1Wpf8XRxZq
89JKskkiGVM9ljw9nRRKonk9ZR6e1DGdqENjFxAfaXGs+jZ3CXHEQLs2K3js0GwJ
EqmgxnEjP3sSOQshY1aQwxQ/GHlK2warIVCbOl0b4/czxl+f4Dvx3KKKW/haRqf6
dQt0CLEudRIvpoB23o2Q1VaspcmpxqVDETR6X9jMs4bIWf3q9vNcvp7rQGfEys5L
oIBW0ni/n8gzJA5YhYIv9e4KqEgqLm+q3NFwOIsrAhQOhwbQS28Pe/8eivUYhjJZ
TMiRCJwk1V+tsVsIqUzylLghuNWKrhxGfV0m6QzkNRP1rvsFw+2E7PF1i076y4Bz
4tOV6u0CHVhUsmqTECiLISwxV7jU/hVfW4kFVpuVCco=
`protect END_PROTECTED
