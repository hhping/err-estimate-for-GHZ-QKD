`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ODCcXbNI7xq2aOD8v0olu/fDQf3No5jYxuwYIFRZ4BFM06rD1DViKwTNcpFdFk8l
L2z+fmX2Okhntl5AIYmZxBg1Ghn5ABxhjAgh9dx6sEcp43jrVUZFl2Z6lLl9g8qX
IzT5BQTCD3Yg9z11C3jd5ZA7FSLsVjI19kCrDVnu2E3iLusZLqjN7obCxoiP0k7j
8qDOWnOthdH15cqDvkkQ7ly5ekEAqwYouAQ2BduuCRgoGehB79WQmeecgzCtcb0x
B+NPXuOT7zz5ZuJUgKx2hgndO5UelYOGT/WzCO/3D0ZRy6Ug+lDHjBWWHc6arvkx
ohlP2TPTMX0OVgiStvR3x1pK/umJhD1+x1rdRBgcif5L/laTok25X4dnOn4rksSa
6ogqlo32xfJR0vnbw83/6vVLgFTYmeQ7v7IpTBkXr+6M0C4DkU9GIk8NlaXIbJiL
R+qtH01dpv6cSaax2QDWi5ljToijrYcKblFNYm7vB3zVChQEhZ9WqffcpjpjGoE3
cBNmJ4KXbJawByCDV8Ik6qRH2oq8dddXc/1wZS9W+RMt0kpFS3tpNJf5ALunDQLF
6MfroWgOEDhkznNaAKL1ZzPYAPN7EgFieGCb2D+VGBmJyL4CVeh2Y3Z7kMOp1gTj
2ldAPwmPeQi4z44M5wH57zM+kaY6zSAhkuFZU8gZKDeogmC7aJzCs7tPEUeThASs
2Fy2iZwi9T/DtLHy4fvlEnmHGS+UOSPjFxyAhL+hH/Js3o4OjeQ6c3huZ+/vLvO0
UMkeIBX1Ma7e/qtfHff0BDBRCyUPnuT6wQG9qFjuhKcA79T+bteZDmKd/0lEsGsS
AbPRRUyeF7VrZt+rnoPiGPRfnYXLPognMUy6Xduy3zvYEn0t9YMHc8Hvf7QR9lGW
W/OeWOInrcJqeQ7839RDzdHierWJWZQQpMVwqonJXsS2ZHbsAw4zXDn6TEkKy74A
E2UZudWgp63fumyrdrs9vg==
`protect END_PROTECTED
