`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QgZABtEz66vznRqb79OzktcS0BnrXJmkvdxsZYldgOBeGTMBn2zNaEi4ufLo6w9I
L+ECDiL55TFGzhcygnINIDzduJBdkg9iQF//kxqJqnPr4M01bYlHAuKjwOc2TbH5
ixTtW4cXp4gDfOPSomAvKPBVsqs5xiPrCMFrKf8zR2T78oH06cvxzHQHJC+4u2nF
nKwPaWv9DDgmN22uCSrnp6F2AjFBWSvOATD4p23D06l6IlxuCZOF1t1UU7AAEyhu
zezsEdaH8tkofP0bBfaTpyIXYQxtMrKmjhnY/TOHy+o7Zam9B5NSbudhreG69mIq
WXknnZNk19b+N21daa90rW1cVQvLa64iXcryN7mcPOQuUuDn9phG58j/sWaawsEN
ogU10BwAzKbteG5iUJLuzfkpbwUjN3LzgJBK2fJMO62Y9yEVsHYQcYMwdVfguK6+
Ez4s7rBW0pn3d8Kn+qdo/Bv6befBNb7KzTaMR024HGWlsRqyVyfR8iItnF4JXb2d
OlO79YBXlE4lBF17zWOoKTpIMplzWnc3d3kWqOP+OHo5NZ864FZ1Zh5VFfv7LrjP
AZWZWTUpXwEBnzEO/Z4Vk/xZWPXVQhOpgGEPFzlzO9tt6RwwpLO3FpjiYOWFwZeF
Bjpna2fPt29ZKliDFCRi6y1tT/UIUfn00ynAj+Bs26xfttNNj3HvCOlXMIILr8A3
+tqbwBy6CFqV8ssJloqhye7Cpx8VSB0l+wseShzsbQoaDmQ8+r2QlaRku+3Adlub
4Re9z/182cfdLMRqFEjRHioq1rGx/IH0L28vwYh3MQyyIsG87EPn4gKI1VQbkYks
wqHl7R9DqRdsjkwCMwCgypeK9oThnngOMUfggzK1bbKdV/Z/jC6V/gk6kYIuHXst
e/e8xslRMT3aIhGyuu3spRvAMEbAWggQfwIjNNyj1tgXclj8AdP23K97hjm4kvMQ
tabop7C1++fPK8QA6amqx0dysb5CJ0SqrsbVmGCWrv5MV0ZmIY3G7/eaGBf6GjN9
iGlFwlMU08PwIu3c4GimjKYsPKDOAuX9wv58XqsnMv/gJ1etECJUiWSvCSIN7XB5
Pjy6kIoZcP8t2KgHOvG58pQ26Yx/AVo7WteJ8GdDOuixCanFjHzLhXejSDpwtomV
`protect END_PROTECTED
