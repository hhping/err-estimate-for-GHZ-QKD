`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ngC5/oJ9xco+Yp+20cbqyDcvZIYkdZqC7lHKlYnAMPXdMWSAyrngVF+1nUTn4438
YKP06NyUF5NvKZl59xXT/TciwGEmSMKBR8fyTW2cN1vOnqaejwWj9fcI1vKVsX3x
1h4oxJtEi0Yw6OBdCXixjH0d53Jlj4u1BvTtGRRSjTiDl0qOUj1PqdCplEKSwLAp
PFKDyBUZlBkd+OyXzL1wlGgAwpRZBEattjw8gqqviCgOuNNhxUZ5dR06yG3bpwBQ
zyo5wTOirJqT8d75Wv1imCEQp/2qH5BbOwTkE4EMNZH1nbehd0p03vR7JAxQQy0H
jaUzNZUQLo+mfrgKaq5qJd070tP5SwsriUrC/210YcQla5PK2pfYrzc3Ahq5S5KV
kdmSjFglaBR9IogEXHSXlfxwWX9D1k6bqWrE0P4KRnhIo02eRKTQvaUD2Br1oiJo
O+TRs3oCH6Pdo5wxDj+HPd0PXSfb64t5jQKTCT6lmQfEcu7eGQSu5CQvzdJJvIZY
ZY62ZhD9scNc/6OOXi+8ef2C+UrPjzh7U9rUW/YeUd2N3bzlsV2/S8AMSORyxixd
cgHlAY/Ly/CLF9OYaVc4HWtGMSvOhcit00/l2SHJaOCiU+oBpEHCxQ0digrnc+BF
o5AYEg9Wp1aNDjsItkCDhnvTI2eO5mi4XVzWoecMqKTMEBUbaAb6vZkkkvsAyBDU
iOPaK7+QWQm4EvUNKfprviLm2cJv1nGPVLoAXEeqT8nF9EK3U0bbZUgXqQ6I2/ce
NrYJnKXGhbrg6ARm6wuYcyIR9+f03bDfY8CezbZFRzTajI6M0nL681ZvpBAnpMak
`protect END_PROTECTED
