`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pRU5BvxJsAk/ObSou+FOzWQ9hBoE/hx+eFAXGBTYk/tNMLt4h6yI9YHvS8VTl4NF
BveqUJEdS71NgeMLSQQBiD9ivtE5kbxpFZlKX96u+ztBYpyKs0Ehgr6SuB9eHtUF
BsH5Tej/9lnyiRw+AbT8I+wiePZFxi2J+P67h9jO3lhA2/Rh15nnj/4WNf2JYG6L
2TAsPSwlIDr9A4gSamYbWEpvZIv/pedb0Dx2DaYQjG0GYK7Gy8jGy0YU7hHvSqcc
+YnY/YkWCZguxAogR5Rm+HXUsaZJ7dTahDdK83YOsGxJRqm6FwocWKKSGm38TNPm
BIklQqIwwHvdIZF1+tCH9Ng9bPxdHbuwo0cRWfaXsmHCjLd7zN65WokfTYRxRwE/
P6FGuMXuh4TXYU4eh7D8YMAl5/WChzxWFLsPNmfFG87suY6bWd+LE4ElSBzaP82t
M8HZRaZxO/jP4kgitQs1+bbwK31W6gF+2fTWZ0BczcFw3AjctU4rRufqcG4UOP5a
w9wyHr7rdKoGC6JFfDfJGHq82iUJHVPn02Rmq9CoNN2l48Tn6mhonKnwj6dQ65GO
Ki0T2LqFJQVAlHqqp0Jz2kYrKd0CQEMO4U8uiz/J3Tk6IqWCSKBfbCk04ZFvs4r6
kcJ04e+XqO3EYb6eCdDbsU/K3Z5Y4YCGX1Mkldwq5jc5PNp9BbSTr94GSk1MR9jH
AWztJGVnfCtKYMHR3lRM/GJMwrmB1HiQn1tNEF4wadjgPmkROMexQRTgYqkv+RXb
JdLNC7vDqxKOB2Ud5WwGPQ==
`protect END_PROTECTED
