`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z/sC9NGtNYDXTeWPvmb1uPec8BGHRy4r3UJ/JBRgjPQLbUKtcHZ8EcT1NzQShW6s
rYgkygiyF71M6+eDccNf2y+BH9lrqO/in46h4rjXbcy0sVZQi+Nw7WSeSKhd9myE
qumhGzh119zynzSyoEZPfi/TTVG0rnwrvdO2XyPUzhRHm7OYYee+m5IWTPrQ5ivG
3M7RpiCmZ6PyyUca29chaqPLn3D4c/CqkpCIS0EvGr/wgWWBpY5RLMkZZ0jmTwWR
eF9PqyLQ4oXud8ZAy26X8Rsw0V9js3CZOG2koiuxjWiWEgv2nO6KvXjhUXNcl3AJ
FrQbXI8jj1h+VYqlnLAs93onJctSIsJ1w/mRBorTwsFtfW9+7wThVLAzTzCUpbjs
s5HXmkn5JqilyOoC8vKs9vUwzedeK/PT/+6M5avz9pBMu1AO32R/7ZAT1PPIQyKE
3Eu2EdmFtt5/7FouHeoeHGoyGcMpOx42Rt34cqf/Ml7QPGFsjVE2DVefjUunLP3n
ZGltUJdIPMlkkuhU0stsOj/Zp6MO3y8q+bKiD75nAL2EtpxeCe7DAQ0dGvnbxvVs
TIXr5CjfWQM9LKHtKOXE8gni60KowhKKGSySgGR/6FtW0NKN69gjJB65XEzjYofw
PZ4ycIvcOI6ybnuC2smzHg==
`protect END_PROTECTED
