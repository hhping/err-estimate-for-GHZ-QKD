`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OrCHKLUK5bPm0EQfjI2bubwqJaryysqOvH2JICUfChtSjtQ9kYn8SI+S5+lkxOct
rX3CndUMmAJduABregJ9aMJR0KPjFk8IqcDGZG5aO16+VZK8kaYluH+QXTsV6/Ml
MT38NmDzoJ4HLIBIRTngn1amGScpavtCVT+UTs/m+EUMPTpGoTwr4ZQnKk/KF/bg
vID6tUooY+xDYre8/3czPAJpw9/EPUyfoDCZAaTYwkdRKX0qJMjDo5po8HfbrOPi
6EqxrFtm75gRPJhFHSSuFikN8P+0584RLoaNpd3YxFqIeMGoOEWFphg8p4FnGYce
9JmTEpbftgFH3C8rd2wrnRREKi99LRRGT7EdWks82usPCpOndrNB1UhIPIfgMKbx
2gY8c5JvhXkOdikn9J2ByVW0LzRXEdvaxt2i7B315hkv0casb6q1OhPta2Gk0bMF
MCgY5v9MIoCWuJqjqcC0ydgHLQkVrNUrJN0ACTgy0Lu3fNWUukG+GqW01wEmnO+k
P5j9JxuraKVHzdxf2cuFYBVNWcEV3LbkBbS+2ec+EAmFFAARUA0ck8rcLGCniQKb
j/oAUPwwMure6EjeyW26AUlPBQMslkfF8q1JlDKuBwAZjYIoY3/+Bxloc7oYueC0
5NqGKkSAiSPCo3RwPGxbK8qE4Jd+Spxn+gQmC+4fU7plbVDBGC+eICaYzsIrVYTz
V185eqw/sS4x7OdhPtudDByQREGl8GLQKSr99PwZ6/lKlzWkyjoJUcL+H8oXxG0Z
EcfQ4mqa81oIxvKERIX/VU0Asv7oxmMdsFgp2GT8U8nfbZvI5wNnueblQDtXOhKd
/nRaCBooMmMIVVhGJmUXW+Ww3nnGxAzDjIKNY9hIFWhfhv4hNUVGxMNMGBt4WkFv
dBQz/eWVtEp7gc7ylxyEMUY+ZWAZjEzALOokEnbfwpTmHPHZG2IV1N5CHbwzN3Xb
DKOahdKXU4B1Sqt4cQG+CK3q2s7rNZLnO24NwSr+kmzqtlGaxkGs6LVd6eqZaVLU
wLfHvm3IdwOjcWniN9uh9XfFO9aXENjaN7e8hZb+tO6jCg4lyr7n9oPYe4NAe5pC
pEcRpQJFF668aU1lTNE7mLF7XGM38cmRgSgNaJN0tmYcf2f7ceN7cRw035TCThSs
iraFeZmmTWz3BKcX7szJWOQrL1PArIUJGurO2MmZmpgufd1STvhQkfFVfHAInI+R
rXp/xosBJEzLGyBK/+Q9nfAVPJZpwM08CHCQb2SzrQGlVIfyWAmKjq6bsdmdo9lb
1lPrAnjDg9+cyuXACr2fJo4B9qJWWs+s97Pe477KRO1HfEjIHW3jJ8dte/8P1mA8
vmgzhLEkEIYYnDCzO+UWZ52U/VKI7oOQ1pcU76NusLHlyYgXjol2NVQ4P4XPTl9I
mGjO0ftiu+zWI/pHRv9CCei2hvvrGpAe7MwIVbL0QuvC7a8ga4493kTGFrWTvE3n
YyoY/GwB/kd8dAmC5Dticqsbu6bqpTqY1XDdIpRsdNfnvCy84Oxc5Ak+Zs2h01ff
ulooS8cxX4r8jhcOEEHf1CyYGpy0nv+CZe4vZmjYUM8=
`protect END_PROTECTED
