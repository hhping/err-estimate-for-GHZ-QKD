`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oSgwhCzs63y/8dbcvgWONMP5nLWRSs4fSgtjC3N8s+dxxS9yFcabaQ/W41R0NXo0
JfvwGI5MLjFeKcdY9+X6/fkVqEZHTG0mAhMMnN+3lZbN2mSzGZr3zYU6HuVClVAu
JaAJGUyjG8JYf5wF4WbLivYAE9Bya7fhJBu9Kttqg9KgjFDBOU/9c/A4C/Ilb0id
3kXZrIMaq/E2f+bf5z8qTzx+KNQXadfwB9vQcpmgZoOOIwEBBnyvJvgxOY0j5yUW
+oA3Czuh9pncHu1hmDSjWhYfNAdjgoIyad8GkPL0QDW/90c/hX2Wm3BEYStUgsZC
Lqx/ckrgWjddkuHYyREvz6bPGPGOsPZ8ecQxQ1vfySEMK+g7eWYYDUm1h8tmpnwi
FvpZKSGkfmk/mAllwG+0szVIWd962MqcYtBWOWNOb1VA8Q17PdOG7tZ5AWhF+2u0
G/P4MlbylddaM39NFb5xXPoAF6zg0jESH87LEa9nIexpWnrVez8nDi4DmDa+9Nqk
4hSZlnFkkJzDGcOquzDkuSBKQN+qBzgwJZyvKhZqX8puUsQZJkh7f+7jgmKXYPBc
v/xH1cryxa7NMIM6NngI8UXL0RI9o2iBExy8mvwCp5HIui6DwAByu7xb88PswZu/
rbhtCCjRZcZclO8tCn0CknFWD6oh6KXqj3mmHhIGFFcm7CcdSjd7LM1b+i/QiJ30
PY5bXLm60e15ULZhA5HEzY1qwem2VafqvhdUFsDNTLA5oTr2aEIbU2IwrOazlRZy
zXG6fhVRFdZuXiVKVrc0dMAci6kxKMHQ5jMr84s8jMlZ0AUJ3d0Txmyg9c6GLMwZ
CkhZRa/j73jPOSZaShkcUUQYjTCp0yT0DCM6X0UJjeWYu3fvgN8bqt625rtVWEOG
Rs452CNUEat07ptR0+ydjbMCQSmqzJi6fYaKJ+R5Sq5cW105MDs+L3GHFLE5Kdq7
eFhRKZwT4tKP5NSdsxzPCJwdy8xKL9kIA+wMi5EhkfOiABcCp7eNKN8JeRPlimo9
v2Pwxbp0iV9ywMSGOXq29tQJR8u5hY5IIBKCD+TKQ0ZtJ+SUdOseYNPdqugC+w2A
8qnN4k6Ha0fqbMnRIKwalm8lnEeHhxdldvZej92LH1Po0QqGEO7lYTQbGotrpE9l
tThyYoSgBWLFIfmaDvYao/ZrcpChKMM0azHe3j6fSyz1CZYID0lIQNv9UfnTYkIl
NUIeqX20vRMc47/sOtYyauMju3F9JfZMkbCpmkkrevD03bkTJ340UVMABu3sCD9r
+Qs89MUKIk09c3DSdHjXbxoQp8CMg0uymlNH/kt+Ieh8i36elgJjBSHsL09RCIX2
Mi2jMyqlnVKFlRxY9U3y/GQunXLzBQ6fvp+E5t1V0bE2wVjtoyiGoSrT/c8+gGs3
809Jm2sia81Ff/trdFblSYtDeqC1boPrIxDAZrTAxcmArcBUHyeNeIBbc9mu4jyE
P4gAl5wdP4/WaXQoFQMxIdZfAntzl4kbUtW4Xhp/b3O6edJGjdDMEzKXthrmXg73
lZ4yp0jTtIX32jzeP7tJyVOq3/XWem665YYCPulZSmSDr5boTBD1ZaFZ8/0qvH6w
NohZn3V3htBwY2IDL3MMEEluZtK5LCZ67ZvqrhQAxiXh3bVk6NTm9eSxYTERe+SD
kRLU8y+h5yzUoJ0EIq86/9rzI8TUbLsWVeabZlwvXg2msjKXSjHnbO5W48/9cfNE
stoDECo1zJNtkHXQ1Lz8HtPrvsa3reIlnGU1gsFwI35wXQkg5M1q9tA0YJY6XY+R
S3Jsb90P9CWnPaYN0xkJz/J9DPQk1vWrrl7yTj6FPihmFCjAX5uJbtqyrG35Kyin
0wml4TpBKwROGf4pKAw+x5MqOODCD+iF7jaaDfnlMjKDkcRJO6BKymT2HHbcGqHV
ac0grVCq1FSsb5cRcl9PloO41o0nssCI3DA8iKEjZtIrRytW0QB/xfi5KoH+8AzA
iURWiGxtoipBZ5gFHSkbPBTNZxan/6bHGhdCFV7AnIIWqQT/QOFH/EiKdxGfaxXs
acvIK90AW7ukiBEVxL+HWlqGhPnYmJZASVg7TbNGb792PmsoVBg+Qgm8SnVLh6ua
022su1R/fzzyc5lU06MFRcXnKRR+VSEg1U2Nh4192sTMLAwbdbZUk1zcdSk6DvN9
ydnHKxN8JYePuuZ8RXUUJN6f8wbEv9psC3nbByejGJZB3qh5sDEApmEv4ZaqpMDU
R5bluaTqMh0C89dZgahRSHBPW004q1ZgtnUuktBTeoUDV/EKUn0iHzqffmbuCq2E
M3RH4X7pBY1zTzOuNn7gl/9j/CX1/WfdCGEVS5tn+MY1QOSalKy52navTH+crLpL
x0PBV0jMHUWMvxqf+jogLds03ZgXjnseodgyVimwkeL+6gvAewzE3s84FIqI5e1X
bx9RtSYYotYRK4A1pcbMKY2aI9qG+ELA3r7PYAuFiXqU0WuFM/GF2ozsJAaZ8ofd
+WXz1LBIUQBRFtO6z+UJYfD7DTP7sT1qJvz+Wd3QFamMksyeuu+KzBkqEgOM43IG
A24DPf1N+c8vbunJGsTWelhD3764ixvtNB+L6i2z4h07HQFwbnaB0WT+nlXCA+V3
d/XtP0jDeHay8QK5IqbNa6HMQIw1E4HXQGD6oMZd3/uDbaMaNHOAQiHI7lb8Ijmd
tZpK+W/s7i8jFibstFHIrG+zo1CKRuxb0f7Vq+59X9u4FjXHG+EIJId6wxfyH3jr
Ei8LVLfQXTUoJZMv56cCKD7/A9l+T4pzSIUFFcDKulUy+Lma6p3PQLtDeyd5XMDy
ARfUctl6AAju/VwBooBU+Ko0JwB7W6AGbMfqGbHLjeYAHvT1cWi9B3x953PTJulM
YgK/EKwJQr+5njYhAzihS/7G3u6fIH+GhZ4Zf9kjHLR2xWq4OP7PhqN5f+44/HkY
tFzkU6FrucULYKEVT09PI4Ngf7kR5Nu7vZhrOW6nwgE/6JbaQphfNzYbVtNhcZzT
zaXPkid7agmx51GuDXIFF0abRIjM8u0/7hLQy26CBBfHsDkQ6ohaI2FD8xdrBUOf
8CKulyQ+1ioza1hxG2IOSXTTAu3JsKR4CEO96gkuqw1OqoE3GBlxiHb1TTrJFDnA
dN5FYvPcJbenoJLQr5oexgCHnXGoqkOb5HozlL//rvZGBLJEAt26Z0Y+czj/QJIc
v3sUGTvOggjKSChfhOyo3/EBcedH4Brz7SeawydoVdq6LWBG/Y/tki98lTKLzBbi
w4Xi5eXolCBc/yItbWzneU+Lah0z0Kvli7Xzr/rXh1kBdwXApBHCek8Klt3AzC9M
hIpAtgk1bkhWLz58FB5XUlPe3FqbHWJTtJyFqnDRhthThs6FsYAGeTWXu5OIWvJt
A/h6h+aSjIwkHCh0KPsrnvMV46sWV626dp/+M8/sA6evjqalqUaOR8JZW+sWsjOX
DyaivLyfNaS3XdM1Ief7SBBe4rwL0qCSWR3r8dUMPTu6csiL7DHnF20ARpZvpFy7
KIX5rDXwoJeZft3gb9fcGr20l5SZfudnyhHONYC+FUSQCmnwX/N0UIcDYN1h6gsW
vo++96tFbe3nd54+cr2WWRHTGU7ISEDwaKfOMWEYa0yzBvLhY/Jiq6gKX8AAb4yJ
wt37bwhQWkcjkQ2+nvmYT5AWc1D7UzIVzKTPEP6D62SK9PTSqzduLf7a2CT+omd1
YNbLaLorQVD/KBoRJCt47nsfzAb6WHTq79ecv7FGQH/Ycp5tWyzEB3VocEGaj/M7
0gxTtafZX/ErkqAOzDh1FFOgT1pP0Wmeums6p+kYlFHkMUgemFlSCqoXdG8QfNDG
4TYDNzjO2nk4d+bLRTtTZn5RTalFJjyvYH0QmQzDc4dXAf9voPmcBTGOhhZg6aea
LXl1A5JY0hmfszEJJScaVaVSJmVQ99B36pldRpG2ckwWK1d80sHYiJlSJLGARslE
AvpDyeH0a1/RnQRWPmi3PI7/eEChdY/t7wGOTnu1rEJvT56qQ9yjgtHqkywMoxwJ
2nLj+S80C7qnYP96UsyCWIUR3VzkoaS+ZLCTEqurTlCXiE9vrpWWRY2uCuNIkmTx
pyEvNFOiDEuaeUJrY4EBZAY1wb6lvui0+TOoe22U3iUgCLJIUxq9kJqRFlJmXKaW
GwjXHp5ixkn4lwOnPoWkmL/jH+mIdVQUCCwg4LnxtzXy2zxKdUrnrSPJvWctoAxe
YaVdsp5+3XcunPkuoYlvtCBsJwkYSiRM1GV9t/L6oss0LlTf92woRmsjugDGYUEj
nhh3OTqmP31FxdsZh+hUJQWIjusot3h8G+yXSzqV+9qQ2OdlZqu1k7mwFO7R9L2n
rJ+hyrJekxs9wa0r5rhA58angjfmMyZiANoejNbPMaYmcA9oUs3fNhB826jTlRBM
/7nSDNUqv2/BNN2bbbZImGvWKJMdKtgWnjKR+9jx4YGKdDW7rzHskEeckQJQJhjR
oQVnFKCfmxTCj/jr3BucTrGMTypIo0iVYL0F5WVAHIeBqIjfPfBT5mMOfU1s+w8a
7KAZzIJfgOl1pWtN4BGuJ47ewqGWomFcCIb+Ga5pDBVleWckCakWGEyiIXYZUpS3
+wlKDvwRyOCDfCBLL+9NLA7/PqlB+Pa9hU5nKQSk5nMOSSyxaxhLWjIJCt8b3fsV
SImIT1mMQzJZEZ/zlkqUXv6cNtty1C+Jg62mbl7O7BR1eCIonojixpkR6cn3K7xn
jCCEIOi7M4ca6aFVpqyUb1HoyHR7sbiuhGBPesXQDMiRlukFfDDU49UiEg8wdNM/
5TkxKaWTLL5BG08T++rr4GQEH5A7S2n77VG1agyA5xumx3L4FRze6cYbLomaO9yZ
K6LuF8oPo4X1y2PqEW2GQK+3YpCpQy/HcNFAhFyXPC2CfMMb/YLmUeHcB3U4bZCa
qxlr5IK6M9YnyREBoLbJFSRAQGOn8LAFxvbYnXshgBs2n1OSNryD1G2PH2ZBNOvZ
EzXBA4pyf8/k8KWi9njm8KupJdPChEA6Up8SoF1SWu1BU60rmigTRxBa/8DOKmnv
Cn/vnvDDtJidunn9G4K0KxvVI9rgkmnthl3QNNhD6kY67S5Biqx6B2kSYI/5jDkO
OzVdr6a1WgBn5y6f91nCvXb30kctHEqHU3YuimW6xWIj+z91fXOOLRHX0HefRveG
yNYi1mY8k6EGN7JNyCTGjQARicO4CjyVAwu2kPlAqIFJGtwNoVB01ItPDBt6rxfY
kR4bPNzhnmgOY+HlICZLBcdVcxz5vSA0fLeZ2u/X1HY5I7uAf3jM9DgIWBppU7qN
cLt9xAl78mK3xdajTR18VHWjjEeDXxGlP2/zrF1nLqCH810pzlKNnt0g5m46w1Y4
xcISgQdpq61+y4ViAlcodJtv7jDbjl0eKWSBIKHhDOiTbhpzM1W+s2RiWeS+D5EK
h2rOMbC+QZkyW9phiJb/+b2KcslQ3+Q1z3m9pzbX7i5XN4+N0ysgo1bIYwDF9f+7
jeFQ9YPNwkRCMno6pdip9zaEBn00JkLaLYhB87YzNicOzgy9W1g9dlakCbEaxX04
hIFdbzFA/SlYFW2PN3BaebmP6Jioz0znj7fg7BHsIGzWtPTSeLwnkUBCOKeiTDf2
gQ7dJ1Tt27ORAshuDO01VrBWjO22jYonGhVcRH3XgIpTBWnYGSmawt/oGcrHNk4I
90QTJQoAi3+f5/UsBBYQ71Icz+nCs35DwDrOJPs7CEa4PIGHau8S5FJGiEZpWG12
WdVFv871ouoRRWkMhi7DJDM/YQHpOIJGMra6rKQ1VnmEoY/jC+g0KcTpgC7gIg2x
D6W3wyrf7KODGHys6fcvkE2C0369BpeohpyWn+Ptpjj4VIRmh0UqqMAYpBDJodBw
QRBWjcy2fHKV+lVHXj5dFIVEX5Dj5PvyYzV8UUgboqXW+uIg+q3d9hq6T+uzPZkm
grw+v9r8gjfyXVn3UVRV3rLCYSo3y5zUmLKxfuuiDNoQZHFQYjsPRQQg4Gs6Tq6d
WwLjw7bDXCDeMpPbZML1rogIsi/uVMcnTXeZFjO2mcRqz5affgJ8BzNC1Rq14PID
g4dzCXAYRZaIW/g7t+W5dBdYTEH6+0FDCLXaFt1TbEvL/+780z19J2ZV61zILRdP
h1QYyvGJZh6M+wy9b/ifkl8aIErlFLQz/bH48Syodihj8hVD2pvXhh65JxJnnNJw
L3q/yinpCRjkD88KBIPoTe4xRUJSuf3wO2cVMsoEmPKwbUUpQ3Ji8Ov25Pa19pm3
ZHNENPwQyhJwld+FKgxjhwfUvVf62CrOVK03AHM3KwmJ22SWYFHE5af3FlYoiA49
PpL+RBkveqOfuk/qNRTXQcf0mdAb9N89lkjxOzj3xE953E5Vi4v0nLRUBq3DlTEj
1yo02X2PPYrld0W1ZuhifQpNISkolYraJcuQslYutVdjyVVWCTU3NI5ZZDJUy01/
vjyUkeRs7a8jYdDu5/+mOx8Jp8l7MhjyUIf5f7mk3ct0vFi2xaDS2vX+wnJ6Wk3N
YHMc8pSOaGXLon6B4UwZNWa1GBee2tNifZ0/S9hA9nWa3vNAHVZdBTRkwgCLWOER
/NbshQcFgWMF/sK2RcCttaQzfSrllb60lkQ+XRvQ/LzVn1ORN0XqFNWqesY5xO5J
v5hzjSBXB9OMKmBBMue1IT3kA+cvdem8kHJFUmIU63qpw27FlXDNVQS8YsNS4JE1
jBe/y3xvIj0kjmvcRdDPid5tHvYidqeKBFUPehwHFHypBnEge5hRckjT8A3eVZNv
eyjQYXH6Xkv9S8IW7VDGqI/pyb/u50sQ3lKE4Wg+h4+gq7F/sf7aR0Cvlnb3Grq8
YDH12ePFYu2XSBtqFbCTha32CJ+FTKUME73CmNrjD5O8AZfemPIvdFZmK6gmCdWt
2eNta/SkwsuXcCDJrqiLunbMosIU4n8zg2tEVFydW3PbOzAzpMEqZP6kuaTm1d58
vtlHfOTsUyWXNQR3GHfKcaZ6wDHZowYXTJTYBWrhimtz21sohbIGS5TeZF8zdMdV
Lt6uvBViRSNf6qjDstq8G/WHTP9OYYn/YJyc/jFaBjCTltry0fSXwz5aSE2OIoYk
vzm/KJv8AJcmC9Uv3XPPzODyjtFhH7CQIJInsyg20jmNI1tIbQ1YRKOsxUaXC4eP
VLinDwXlRZTgchHccHZuXZhMZUwWP0LtQ0dki5UZFX5gSV73J7inkrFC6XY19LzA
B4IPK2v5ENAYI3rksJl3Gn1a89cG3P59mOwuEKeYVdf8OkGl44Ll1i8KBuauqkLn
1gVY55QwIuHmdAexIBxNMc+Tzbnbh8+IrMmXKk3pWFUzaUoQvQsYSgRGQ7IesJ8B
IOav7qltJsLW689S8bCfefZIYg/kW7EgvqGkkpoRz8r5jfwh3YIS52VUdnYP29FT
1kBkgBvxTNYfa9IF38nAm9zgnarlTA/xaH8Fh8yL/b/ttPPgRKQZjxFhPi3bWG8C
buNaU9EbU0tSQW5HMKQzQe0jJ1nfBlKCvCsHgqZtSPfjfmS9Vg111AHr8a2MHcjm
AnF3HR5AZK10u9zuxqf0/iMA3mUPS/kurAyyj6odNautGu7jr2hWEoxGv4L9rA/+
/e1cBNXRnOGokL3oa/PQXYBiGBV6tXR9ILY4w1UVuOPs5TXbY+gK4d77uIc6vXzi
xzCjvuhgGhNxJEhCNDmdcSWPWKA3pgi7ec3OgJOboWn52Zss9ohQYh1WsO5RbyWf
EJ8abW915Zrk46p6oE8S+TVzZSv3R/8v1IDG9urbUTPjymM1+h716zi7qx5dQ9+1
rDhNvf31g1mXWfUopazC1JMWysc1Fbh/rnXOK8BQu0pytAF5VKMg0HCVQgQ6gHpm
QairZ1a2Q+h24CqjLjj2hRn49VxpEDRit13hsogxubowLoaucagXEM3wM3cFUm7J
fQLJxgn2alx80fyHYLvdX9KTzNiTcGe+Ci9OT9cobyZF38pB4IAXytwfEf/eiPj4
otG9PU7j0M3ufu4KozdQqCX5v8C8WtAuV7PCtAvURNtUftntD6p4U6GzkBrzF0L7
Ht4x9e/4XjHz4rORhyqvqBHT0SDm0yjHgVxhLeg3bZKaSqBA5dksy2mrlDlate8p
KOyxKnr+slYVHIOYxT5bHsYYdgHgqVJQYd+17WED4tfrGUmgGad0FayOMLEtgrvs
MFFIbQgZGSodk36QnPQIGqmO1iUa3oHj03vh7Jg1WpJaJdxmzYB9EhXQIlFn4ZG3
jVIZT1HIBE6GXkZwOIqTP9gm07rFIXM0KEcUmCcUUS/ABCHw+YMqVHrgWJbjKKLw
0cS+KNW6hpERF8RzZ5pmNg+qQ+qaZeDHRnuLYl3aIHpIziXXBkaeGkSgsbLZiQce
G79FDoMEXUDZCwun6GvFgmE9TvEawnECPU238sZ3oDQI7AiOT+e/zYjJIXAhQDah
4YEavTsFALXwdb2bC1WCWI5206FE7plv0+IKkHmBuAC9b+8lckn/n9NDH2kblBEu
76+VxR6LaOhI3522mbPQ2R0KV5ESpCGmjU8yjzrHsz4aT42iGim6vJplyIx22/pO
Mfgu636niPL/jHFHVeFAI/xFIv77MYC3ObtpBn4c5ETUkeDgBBTDb6SjVN/W9dzj
nfd4P4alFzJqeQypYIysdMMh1g480QJP9LnXBf1SXjuzvzURCMH5WYXxuCc8629Q
N8JeToKCrabbzFyeUZKQ5dmTEXu7fMPef/ZJ5psIz3SW+tQeTdTMC7aQMOcyklQk
eUF/qxN4BOEEA9RhOdKZ33QHdkiVCCV3H1KMuOfd2SabfBALI5QOIpfRxHUtM+pG
LMkdE78tVxfKdSNFPG3Ae5rZTCE3GtQYppAKWFNmxmwxFXnX/LL1/k/rmidvcxmA
Ll1IPkVlIjthpJuIUL3GYOIKHXRDN29gUtr2GuGt+rdNWG1/EBPYyKgXYGMdrhSi
hbhvD0uT08E41LGDdMlxxynssJC5GiDwAPs5Ayag3v9XdBhigU3GRWXRon2Uu8H1
ZaqokIvcfrhZKu79OElGmF+uTCSGpV+f1UiN1Gly5XmfofHqqHtTUi+Mqzps5twB
BRfxCVVc5zwCn3tqC806FbiNfu/EJu8JEcnMJbxTR75b2F+nywWr6QpGe+4AtyIp
/byqMWA5vEKwSgt+PAbnw4CN5EqvvcfKAP80mjSI++4TfRGfxQCsqRKPeFI+aY/3
Kkxs9RPZ2O5NnI6H9mYxTuynL0+EJBwKr1lh9yeYxpoaRE/RZ8gkT0e5/gNpSK2T
ySlcHf2SGH/kLGnNfx2vmDD0XmPk5ON3JpPBQAfLtTj8qo6ZUkoNiRn+y5/k8paX
zMpgVwFyKba8sOSnHiTGefW4dQxx6OH0HJlf318G5k0LHLI/7pSnitG+GDoSiYtC
nPcq7OI2lz1EwnT/P8E5VUT6cGhSCbthqocHp/ky2/1r+l6PKWp2RFLV7HA+8ItT
UGxVUFwJZ3o3Nhc23+hH9eXS2MCiw4guy2BSCdHk5Ctk/8aRdnbGDn7qy7DmhmcU
hkHN4jXkbUNTFBBwPN+yurNsXJ11lZHxksdHhq+Ju2Ep+WcQ5x0bcO3kNEMiDjZb
5y2Cko8IRngwe15VIP4x3zECcPCsJ8cQZPw0i2PLadJphxILKiylLoq/PzprHvea
kZVM9z/9lWsWYf/CJpcRKRTfpOHZtpmWhIrjETDgjkdAFj/tzNwD+a9yK6YKd0NR
/5DCRlF6M0jU4Gn33MeFkqdwAYA+3kmHJFlOeMBO6XDQw4uPqak8/LUz3uj99wjl
YLBAA48rdvNwHOtGLN47IYhpGYX0psMbotUcK82hViubr4BwDNzUo3D3FlxwZ6KP
H7aEZBJ4KcQJ9xAs3fERiA5uvyy6QmtJhGY6rj+t3FOdsIdFqhOAeu7weAefOWzy
V/3dRKL9hXdTXJIlcW24+YedIHiNMo09YhjauQyecmR5hXdEwM6E5KteY1alWzHC
+61Fp0eQlgOCQEure/DTXCOD++EckMTnMRjiSsxi2LD2pXX2Zm2p/6XCo1aWwsIu
8Fp8QlTNubm21AC1G2CA0rwfc0ijnTw8rm1KvaOcY7ZEKWzVsBlh6K/oB07XY4pH
jRcgRlwco69dldc6gdktayu9I3yN4zi+N+mdm7ciSxr/MnAl8JZFalQdaCYgT7+R
ZtCBFeILgQDtrEs3UYg482Cvx32THbsB2l3K3xJDa5nQssWpcARDxaz4XfNlFwL7
p0ge42d2wDGXhspD5BkouKqv+5z3IUm/PxVAfJAj6ba7CH+Az6jegHPpnIOayBPl
ocal6qPtjhxa6oWsT+ewrcnBZ1Hn/VLiT0RarOlOWjwDFcTyVosPe3tmMixPU2dK
weFffOJ+2rkYDvEpVdsCyOGNb8J7arGhUqAuI4cZJ1m1/RluQccxbQvH9qKXMIDd
dSrYFa0ln0R0fmg0OgnyifOy+zaF9YiHecCRHw5AIaJ8epXyRWtYeA7sXnnSg03q
+dCVC7ITo5Rs2R37cPYq71lmt0jVN1m1S5jUlLQ67Pxc9xvlc/TunVh6TvuxJxIB
01LHDNEAIdG5qlPt3s1NbqZ/6yKyvKFK1NPITFu91I2HxY/CaZ8wgam818yZ7t+v
PiqYsFuoX3wxdxrcItHG6pTFk7eTasVfjpFrL/6rMJ/yl6jN1ZpmngDA2ocUsP6e
/WahQaLdk4/EFDKb9KJdfJ7HveX8xilG6tiHoNMB46MzEqROq5frqmwCB6QUQ/Ak
353eGr7ku4XbqPZE7BKuFBgWL+aiB46xKs+prKxCqwoUTBcE56aJZujNsi2X9M0v
hnyFFMphwRk3x6bpAff2G1MgsJFahM26ESvPA5M4DCYQ5CtszhPWHe0Mkftjk8yL
LMF/AHAR9Md/vfp2Cy4GQ672K/Lx0Vny7kMv+5dgiJcr3BSIk3uLbw+rR3k4jc/Q
pVDyoUipTXTOq0ra22oVkpsqtrnKJ25+QwZnsgl35OLVxHt6S6LaahysA31wDMr6
wMS2jhAJL2AM4q6ysfYkBItSkOuEKI/MtJUzDGUoFyGtfOXM8lEJGUGtHpHvfign
HeNTTEwEW5+U7ni0q4xqFe4oh0vB1Qu5gXYfmkXJSzCm1iIuH3H1OGyr+Q7w8I+s
Y4s8u2XSrtVp1sV6cJ9wKu4VGLXmEeUQOPT36nKaf9ynSgQGCjsSyNeRP3/Dl3Hd
nvk6gJF4aw6yx/SqqilGxFP9VgfgwzRKzLUlyzhMJOP0EoxbGqrZpFHMr+p087YF
Y9YEFkF8/tXl+iZNy6TvqRrg4B6e0Kkrl/gbNEn76SEXb3cX8Co7SDvoogC1uPez
SBD9yMFGHmXO6KWlWDbJ6ZihF2OEYT9c/LSHr7WRfrpLr6iJ67qvx7bg4kWy1R/O
x0rz3JGRK6sYNS93QzNt96BuKFUtxommMLFVupr3XfCsDodnxgWtZaIwcD38btDt
smen9K6eH7GfRFLkVo689GO17CrGyH6Z3NMj8Yn+ceTaZCTJlArdKtIJMa1eHkrk
YsL0OYljOhWwCEVlG0QXf5O/narOHXi0+rw59DU9eFxIJs0Gn59n5cUe7i237Yaa
bi38ZqjKbLXU7qUr4W+Hr3ruMQFRmCWGcgYVV/HBP+Nw057pnYQGR/wfNtdCxScl
zBnJ8Y6gEm+d7fHADVkDpRonuHCOjBgOWLGSBeZwBdmkQQWacBbWTWlwI5XA/FNQ
bD6KAxtOc9jzwJ81CVR4cyKc/9Urvt4Tfm3DajuPRZSae2ss5o8CgXs05ZjE1zOX
irlrhSnbiLdx6lzKuwJIzasMo2qQueYOqDuI6UBEBv/eFdbn0JiluphFrglfLYG+
UeyDbdxWx4tMY6ONGh2hCLuf2/WUmvJAofMk8c1hsduurUepGnk6sjwOFUT0L8Wm
94sdeYDZc1wkcduwdwPnuIGs6G437YDXvBcLC4ehNeTYqS/fSQIZAM+CddZJ/hzf
NKBg+W54ZjGwcDtOtM8oG3v0J0bjYC1Y+N9Og9z4SCTfV7BhN/V10Alh56HHehHH
731J6KWUFrREkrGGGlP/QY69toYrwnw/HB7Pvwhxc7J05vu8gYjctsplTFgHg/Ou
LqvGyPWAAOTvUSN2DIKBJdtRbdBX+ZZ6jfrofS5MjlTHDc97ZoGOHgiqmU367lAZ
rSu+9g6Jr9RjOgxm5NIW/1VAlaL9aBRASy/QR+XIHxWULg1KzD64DiOiWueBjgMP
PfFzmycYUf2ua2Kz5w9yzJQNnm6EqkDrC3mR2e117vcMPVbTZErrM8/iJo/PXKVY
6UgwCMGC4nPVqHUk8gY7Ec+p/ugPlYs1HdyQuR7Ldu2nfCIiuD9Yw/eqogNy2olr
yA5ZkmeqDVc064cYgjET1SKgJlvlRGJE7Mh7UMjE7UCXm9zX1T2yDHUcvKiyBf8X
MaZZUH+RaFCBRmQRpVNINiiLC//Ht8Dx2yHbUP5S9Ke1Rwd5plxrZwp31SIERcZr
DoDJcOZiY7FmVC9fyJ5KDqZZp76YoeO7PEimHoAuyR9KC+3/NRnhq0xQ9ye2RFVr
2mkGobOrwCF1aLoPNNXkAY+lpJUI3hCGDCmZTUx7AxGtVeWO5jsNCeLmZNHZOpgu
nYXlLJeVyL03eprYHlKgvQQMy2u1oZ4bqKi3iq/fUM27fY3ZE+OTiNDu+XkLf2q8
z+ysXWzHp7EI4nxNWh0yGuPuyJN+NNEU4HnVP0FbsAE/vCR6e9HT/xBJM76ZRhB1
OPM/IGk8qIG6grPoNoSjmOMg75nasxazzNSHEdQEoPLEVN/fWDbPsMVhO2rP06Cd
5n4prNXEpmmVD+rieffDPc1GBCII6z4nh2wuQmbClFrx4qVQcN/vhffbsSevv84+
pJlUric82vBO3rYiwb3MELmFFI6ZKnRUsVjxsY7NhPJHRbWyWiNhxtDGutj0PeS5
IuO3lYcfReCYPA7AVc1NZEzvLDJkPi/BxZv4FjbYnA5+0cY3he/RdaTlT5iwtykm
jkqcfLatVFq4FwWsRNkgVoV62qhbV+4UXyeMzNQ+37wKFW25VSjOB3SgZ2tKKqUv
f1FHHcpHvp8VjORcnT7RrBfTVyvvGn0WVBU5a4UXBWGJVZwwojJTib64hUJyyVxt
KFW91BlxRntUjlh0NsnL+0BC78CO59p1uOvzXsmrxpcAJQvecfb9t4d7NkX54tUS
s0KV1gAFLAUN0x6fb6pY0KwKeK+6UP3YYI2I8mpf+oT3Ifi0Y3qvKx6L/xEkEX0f
ORNXXeZEmt+qx00hWU+fF+qVu5+3aNASJ/94JUWbyLh5IifPVvZaPk8aX08ok7oy
i+38uO6aXwgFBTGhZmSwJoNDAkQbE0hcVejqV474w+h4zY5r2HZ+cXcmk1S/XhJX
khY4W/afehWWov99spzqccY3NgMvhHlP5F/D5BUqPMRKwo/M7hStXi+cBsdnkkp3
ESCniLwJhT3hpe+tRyTypPOUrzamEydIuwOwrsdkQICxqrVvYqDjGgCv52qBcQS3
w5wEz83HoVHASP8oeOBiibGLPEOMF3Pzp+qMnfk9cyGGGQ02CIEl39TuGOY8Lk53
OME4Mcvas61GUIvpcrB2MBkGPWJvuXcV/InYWYXsQKMyrCMkhFI/fShNwvy1UcEJ
qBvXCwclcNjTqZ5sBhZpI2pArzb8iYiW8AiLqq3uultNsMZcK7VM/qTvfRJCPpjm
s5OxMqH9KHh/suLIUFToTnrzuaSVpsOv0DPrsD3lRX1/2twqzZU107Oz/nJJoKuR
xh5Kc6W1UkowlkMhhGT9jkBPZ8puTeUdYYpd97jD3LIybCtZ8yShHWPAvIZ7DLsv
P4lT0LIMse/jKae4EneYYm/1VfnyJF8vKpAwHwHBfNH9N/ClAyhJb+hKaB/DB3h2
EfYV5cxSgB3K3rV5QrOBsVwVOxoxbw3XkMJohLN4po/zoRtRmllgYJIOumJjY37a
8VjQmhHBIp0pBk0d73FjgqrgS1uaDuUEorgJ2gfy0H5xLITgPJBDP2mfn7uNqLHv
1oC84nGE/XMC4HTPTj5ub8wH22SHjDDF3w6l6miblH08PZYcp+b3uSTuWk6crtJo
sNNbFqj5pZiGgacVlMw5mAUQgbSZBonyOp+x8uXFaoH8DDYX7EFRbMSc92uodDbg
/PVGX82aPaQJmmApB24+jB8YIdCb3u/wwfLchqhSOC7TZn+dTusBOcg2PIcXz3Xx
hv1r2gXhJepfJDPMaKjcE4Zt7OW9ESHZEzpaG3I1CMzj8Gxzl2Tvp1UXQ7oJiXyb
DWmQPPHjPHou/oIjhZcCZTVIUJ9KSuy5ESXtPc/ljyaRHGVf76NhA0Zqn99xfzvm
I/DAkNvatZ3PAXYdy7HhHsrpeHsHlq7TAFRgUKo9YKhZJZvq+xX/mi3YKxgBViOa
axXBTNbs+EM1QYVCfHrHN2eS+gHN1JJATwJDAslbJh8b4QzPOEj3ZAGG9fOWwBCw
i30mbIA4OUTszKBDcwZZ67trKARCm+HCAb1V/3STG1E27MDQuBPcoBHg9NbltjOQ
5ujASJpOta8HiTSgCrFiVofmfETQh8JFfF5QjIdYCivnnsYR7Lj4cY0AYY+vWH29
+IF1J/Q32rD/vIeCfIXAJ7ED7Fg1eN+Fyi1PuwWY6ocl8SWrVw3LbyZVD1/waE4q
ZvUn7wyVvmasX6Uoz+9zatVvhxuqq8W+uW+s8srgfJl6zKPRCSAT/Cduzugh2Qwc
jFs01cdc6feUPwt+M/eBh2SjwpRmEUTRkhJl2rLAioU4Ek2PdV31anhNzhtR2LNM
1s+iRASCC3iEM43wZUFH1rk464od1Gsw8E80bNuZT4iK6gJY7FobdKSmRWagtKTD
dlpiyksnlj4l17dF62RlYndktrnr5HWmplEd2e9IYiJyuQy/0quCuPxAFV3g6Wmj
h7Jd8dhGbNdlHwGv4uBKnmTuOKp1kIxfXnY+kLO9SmdjgqZxKVR4p9s7pf3uSPDe
N5dfWfsrs8YoAlm7EbiKCeH0dKJsRqZKWUzP5a/7zGwGoEMnaKaKDyX/NG7f1TVK
pX7R26t0MN2bWcayE9VzkEkGpOFunRi5vaR9FoiV9SHFOR7nXKCzpQcs2d1By/xQ
2HMiBhnevL3LBk8vb7JY84FvJVsGIkln9gT2y3azyKmFHYjKkBppvfQ+lnSIggvb
C9G4xitdei83WlGoVnhizSDYY2InnvD5XhcWyvQSjiHazeayrNwpfekJdg0GQASL
7vkGcR4mSGJOjoN48du/LQShs+lr932b3TwJdt5LHZHL90m+zLEuK9MxQYV/j1tp
CxlcGMsDQw+0BxQcqLtAJOvRlVbX57EiQ4rqOcifyMk+fPcEN97fJXlTZwGcCFKz
MiV2VvMOOFneqrt5h0ORPsMMGFgsqnFvXGQZK6IitkYcw+biuW/eZ6r8v3ClSAT+
ZOOKkxZPl0tkohGAmzDcvWiV4URqd980lwJ3Uif/FMF84MFGO4BH9xhW8mTE8DSR
XAPl/p4q4TVCRO0ptphucVDr8PpDbefs8GXwv9S1b71aTb8WY1kWVBNe9qrwgnpp
NM+HOf3Vc8b2daa/07lCcg7YjyH9sJBzD4eCqi0gmLqDX6N1OJ3DTec0lirbbeVM
hJB8+QNFH5sMqG+3YK1+dYgTCy9nzyxlZxyKc3N3aK84X7krsjwWRY2vpV/aiW9I
7myXSeXzEg2zW+Odo2dOKWJSGSD4IgKaq7n8pVK5eVIkV7JrZBUS/g6J6l07S1Fs
9GjqNekasAhBU5rpDH++Gk3NqkNfUgTnY8wPZ8NvNqM4UaVEvGLkiis3um8yLV5x
6toxOeGQcqY6jXU8GokFzkMHHhiDwDmHRqM/cpgLe54I1sQqK97+G1EokdV9YAEz
4di179h0rjlHJmYJRIiCWdgnxJKKpSPoq/mA1cv766knw128EJcUz1pZ/rufyKOX
cWUFp554mswcrHthZD+fDjXeyUbv4uYFecLkToj0SgcwZ51VqAG9M+1j6FPpuVDn
m2UXtZAbaSg09/tzsjQBuii16NevdeSSD+PjXIfLixOwIkAjrrVALLL94s+JMOhW
bi17f9sKVHRIsvVapHp3IJYg7bkUmBqaqx9mKWDTuCy7M/75HnAt6EuDCBfJBOkk
mVlzVC4zxxjTcASkEu2VHgQJUm6hyTnOqPvM8hdRgeOi+xJH6kbI7Kr6WJU0+6UY
fJUXw5ybA99vtct0r8IBUdHtXDB/Kq8xyo3+jUxKo67vH6Py4T7n5UXmdMM2BnKk
DxMxkiVeVrKdbDyNRQBYakItRjTGBrnUmJqdl9lqV2/2Wf+DQpFuuruvyjMOSPHw
ddp/KODb9Fes/NXTwcv3LZtwq03wKKltH8MHrCxxEfN18NGbFFQ6o5JkYW7hV8qv
bJXSXD/LNry9w9XwcwQQK6wLhvWs+fw0jAu6oaoJdOaxkeW4j9wJ8ESs5BJxloza
onzVxQ44dABKLlor+CYJZ/exrnC/XCoxwpofWt1nSjXR6eCf51lnQ1GQA1LFj5jy
B18rlKRbPq2GInjFpCplVnjP0f18CZvVgdMUH+kWkGu6j33kYJYkNVr+3yxPJaZ8
AnY2rZ9vCE+8mIzpkhbl1foIFu4zyZb4nZ339ScEHiJLtDArnede3Mn2RQFxF06J
YTozEYdQn3gaLU9JU5SzBtn6T0/Fj2ey4gpSw34tcFwp58oxcBKQYE5SSyBDEOXh
8YiDXZB6Eru9Rs1qaW09pPefZczbn0JRvDibST4Bps00j+JHgMWgeB99stiwjYZK
3QIuUFSVeHWGis39VUqu8pU3xileOwmz111MXmMAVetRh9LYABe/C1DvqW/3HAmb
wKZJKO81OE5tqXzkK4ZhCitmnIYxXLVBhJIIg+9TfHw61l82baa4zpoYjAg6S1tn
Yai6Kn/WdZQNE0BpoG0FjVZ8qSpZOgueHHES0VZz/l4Y7KlbuoN6RImwS/WFoERI
FoR1XYkZwO+5D2B+1uqMEHyYztrhN3hjVXHVCTkFOqJ78R6/n1eD5GkXe/RcPcY4
jVtC6vcmPkH0k99CnrKk89jmseEodTF2BKt4vjKhZBw8uukqSpWUSLoZg0iZGEYx
sTiLdmkNOVVaJdkvOYUIacYgvFzkxzD8YsRNr0KmHy5vG0Hv7e0SdKAWmqNXxLGD
kfV1FBlUwEDK54tjbWOKwTDWOWgi4ZUYD//UgVN1XH0WN5ONcS7zhfWksSWs5RGf
ttyZENOVR2i+FAgW6LeA2dcrKX9/bggKa0QB74qP2x9Nx67ybQXKpPX5VmQ5IgjD
Gyk+sK9NGWLmJAErf1cLW5ZzoiyOMKQjBhqcErngjPZp/A1uHyUsHDDO9sbHb/uf
CXjLpTxcMONgP0yHrG+3lrSx8XN9iBXL4LEAvJ3rv9P2h4G4V3aiZ32htlSyVxWJ
5c9qKNZvJQYU8izLvNlNlr6gnV+Tq0thlZ6Ck8IzGXcoEzjQAB74s+eHvqnkCTuY
gCsgxvqNDi8D9rbTsALnmkpJj9mc58FwTYurL+35hI8Tyzqdm0XMI1VBbdMeQTNY
dDPZJdHwztg7SCuTw6SKRW6HPAdoj2jj9nDwSKpo8Yd6eH/LDoukKuDTOC0U8tdo
x0yekKDKyK84ZTPMVmPMCSqEpzzRqy/LOBq0f0+CYrtMw/nDTHXKhUKsnIBDOTBO
wFDI8n3HV70nGfGMJG+vu25EyPUe+zL6vsF+3DqjQ8KV1CMfwDg48XCkmCjh8o69
XRsU6eHv8B26meu2hi4rMLGX7ZIUhplrLeiolp74NxkHhONeGbjJIe9/uZvvPMpm
fhSTaD9qrguGIdjwuRmQlMDxaPNn2OxpH9+ErJ8kyRpdJPvB8BCqmnaDzgdTG/3I
jEGyglLUEWsC2EvlK6OF7qMkEvtRk9SjM91oFlK9BGhGR5lCSsaOFhWMmQLnWKEK
Dqui9rWoaVE6Jul+cCF+JNTruXTWekSEm830yAmi1T0jznJ1lZBvvLI1044B63m+
ojgC7cGzI9mUh4+/oDONESMrk59/COmU7sTXEE+ueuEZFoK9jg7eWH6NcjGEEnlf
bMmZiRNrD7bi3+jhh6jRjEHHT5cmHt53byNb60hefIHmJF6VXNq6PoijQ/EmVWi+
SifgS1NPUSfwCeC/vcjdVNCOToK/V06ywXeT6WBUQ2lfk3Rv5en4M0s3NXDfTg7A
c+DJcuYMnkvXau2yoboc/UfHs99Zq7A35NmB0yt9e0smalp4jFGQs7xLs/MQ0Z/K
fc8mW9vT63eyLTh+/x2y/fUT0iUkTOCPK5Eksw6XdocJ4aOnc+ga7JRNbcYblCq1
n/1fkoxE76iDxorGeTEuKINxqDhL9Sg9ANP2jfoblnCTZcZGZxZ9F/pcZwwc/CxZ
c8bsEEthVq6AAfPR2AU8XCeYk9FM1kpV9TTzdgbLMZf397tmBITke5R2FS9g8m14
XNzC7lvQw85hYp3ZNbH9kgj/0B6910INIcxZ6toRnUESJ17N4QXZ8aKsrHXLx+bR
43J+T/IVdc+dvYL8tc6ralDmf9Q6wjWhh+ac7vzDkxQLCUxOAlHEQ1OHNdYnVNIg
jtv12nnEpCEPFItdNQP80kH0fmOr3vLMue7p8w8/XTow6/NI3HLq2B/bgNFUFvyH
VVWrTdeaRAwJQGCDGgT8y45jljywxUSTSTGsydUh3RoMG8xmdvIjLT/1Gq11JEUv
UrrvAF09rKhoCpMbwChHeKgejJuELegycNXObdkL5fzkHr7Fh7on07GSgkBoweL6
cay4yKL4X2j21p+Zc3SgQNEQCOKpZY3y0s6LMzcw6fV3TnIybnY3PGwCanl8ZaCP
Rfkl72HbbxUTr2yE0lEQlcu24u9IKbdHoYpRA/lcKCa/7MEnmCx318fn7bibw0Me
6m/iwq9B0cUPtzyb+rfDs7zY5LkWzDFPOUIl3LqqxkAiabEDCTb8uBhPrOiXvyJT
CfuENRRpasLuIqmG7YvUT46U+Hu4tw69sL36fQOq0QXINWPoQxrwC0cX9XXUyzQw
ojgCprrwqWL9erIlDD5LOmCkpHIzVLpaSX4XdX66vWj1FOavgtBrBix74m/Pxdth
pAe4lLw9CwONgFpqy1X3QmuBjQAgRlBqFYr+yBJE1hn4OU4+d9pqVhlcKXW0gzlC
FayosFtPJqxFKbsJ8iMoD3cbi3j14SOExDydfoovDm9/ghA2JX/hvQRgtscIptpL
AFP9uNOrXX/F0eh6Jy2iioNU/JcXO6GnAI/oXRsI4xU2hopM9eSGO4Zht1pl8phb
q68KycAgUWFIiEMj6JbggSYmIoysFU8Dhuyiu7GnTNdVMCBuLwVQPwkrnL8ieF7k
HO5dchF/m5zwkyvgR7P00eF1aouwxJOPB/WA4NF/4KjXDSmb96MREtvtAXMbXY06
iMlPY3tnJgrW1rV2NK5NlD+QZTXQLV0i6n8bZB7AGT9DqKGwQCq6RIl9bdDMUF+I
Zvx6UxxYP2TYTqFAXRr2JjhOqZd68LTkrhYmNSyGhlRqLEriYx5m/IxKog4o8D77
+9bFvfLRMd0TGrclKmZQCW1q2v5JrYa+LU+oKDdRfAUS9KEx4NLcR6WB51kUMoH2
7GbTDuympzIyKyc8rs017VUqvvK1VWfDZA76vQ67KH2LvhWGpXBbZgBfzPd4uKCG
wuUBbKQIZvtqUdOaKt8mu2XUPmh2fCQ60ZHelf1MFlTPsW8cTxflYPfkMgGyvFwl
dMb68+aqlX4Wkn80yOckDCXyouLJ8vGksITFk7DuBW/8fy9CTYaSKJx6u+ItCri0
S55pjGDd1aoltcUSwKKrCyErmAMoujcaVQ33qmSIbZg7d+ZCdBJ3wLs3orsnRDrh
1G1qxQGfxnaQrHuSITsAnqp0PwDwSjLtb61NBAv7frPyNwsF4hmfgsOYDINhMQzz
U0MD/NebxQQ5DhJPitYK/lTUBSK9hbMUhBIjrIgOEZklRdLVT9Rk0Qj87Z9UckkD
Y28NF5l/NQ1YfTx2UavquY/BfGJko7bBci+o+haHs22p9xULOqkXzc1sefXIVROt
zRx3Ac3bWoKB6lLwJ6MuAgNbux8n/ToEQVPrCe2hYkwHjNbEGwgiYaTyiPnw62Z4
kbj5rYOy/mPWCDNv2rYHHnTF6/hLRaMQNLzzvHUu6uLSATig/tsgJO0UkRoAcM9o
MDWoyCQSpWL/Bft1yxLOwHZ6dDb1/4b7x2IeS2Y69g+/lD2ySVSR2QcOeqsPFh52
JFMWcXj5EPIUPh1QI+EE40M+4b25/zize0MDO2Sp/dN9gGUZxQJbsIVSJ2icxB/f
ZMOZLD/hRJEIx6e0oq5+kCS2ZVP0QAxwgqMnzIDlcMC6+5cumvwbqa66fXxlTYoL
pwcCEq15wOeyYX5IesxrABiLdCiW34cFxPZsnK/E0XM/+nOu2mlGdf3GbMOihGm5
bLupP2hoRNsguWV3yRm9j+Y/2QHUQiDCkqVJBQD2ncT7XfDPXA6MCWXvJ+BzfSWz
d6XE9nTttR5izjBX59VDux/ARijY7linHS0aI19puoCuUXMvVyaqz5KhhyQhBof0
HIU/b6zBjqpP4MSU5A0WgwyrU0X6EBv2KKHc9+f7dQJWXFeGNYA/u1UpJl8Fy6PG
bkg4wmwV8inXQ58R0lVB8Szd2ndua/Y4wq4LMjqW7eiPjObj5rO/RAWIX6ceriSL
P/lq7oTQ0Pem97suaRPmsMKMxSNTLS264x8S5V56L3DMeRU4VDfA6UxZvLIP/8NE
agK3wy/FDae/qyB89CF59m1yFyCwxt4jAsLaS+MdxXoGe41YYP33YmBQSW9B2mvb
EFHZggb9KeSFzoTM04ywh4hV59BrO3yTCjlZ7ifNZEJhNkhKzPiLGqNMxnmNYFMo
iXJ2K3iZOJDp2fsWqWB3mhl3E2UIAM9KcYJyGjlPJcf5rV2025ab/+BkRK+fp+0e
szPK4Be78OYhR2Nog3O8S/hGBNGkG50clNDODOpTs5+glRE/DK89JQOVobZjzPaH
bK1EKi6H+OpUcUORG6OwQeYzO+9D34lVzkD7EF1TKl3FJg83Jye3u3L4B73n6moU
W5D+nPpitHvb+Sz3WC0lNEDL1nRXRXAc8cwcDVRqO++M/OU/LlnUAzOFhiO2nWRN
8C5lVwPlCoBaCB/DqM5q9pyNSVvZY3cihdnWSiVwMbYHzdHgqPUdEk9f6EMz6VOT
0BPNXzBdwixxFAdMuchOIX9oPbDuFGnBNQnii9VRrTFlLZ/D304JwMzpvoIjVeUX
ZKAfZut535y4Vrtx5T62ChGyEcND1QOexKgdbVoNIZ6aBmPWBZ0F1HZ5kyxBhsON
HPs3qdMxk0xM14kkTEgfPUERvcrTSlN21Z87k4e5vx3gT1VfJxykN2/TnBW0vonB
YPcB62QXtwkPniGnO3+AyrN/XZt+Db06DDOQANGkJk6Uwkc7X1H54IVJnycveeBa
ZylMVXXQoH4dHenfYTbfpCXF5p2HZMhmNmX/nQ+06y91XwX0PbAE0mV03AZvyWCu
pjIZqq2jXolkj4FtR/cVw9k2a4wpf6G8Z8+zLrypyxSOVv40RE4Wv/vM9Db+Vu9/
qoA3FE+qsCO7zRzJhX619Q130L4scEp4Mee4mGMBSFxj7alM4JuUm3Lyh4buY8hm
sbIRh5uh0fvADcnr0NitP3MRPnr2gOnJ31mKJjNKMzv6ZreHKhKy6Ooqx0E+/Ngh
Tslp6nvqToyBWuASY0LcIdLxfXyF5FubKkRn5KCEmroQ5PzbnfaF6/y9NEZkHmYD
Ba7Fq85d192nStwhlIFu8zIfgmvd3NXv7QuUB3MNnvLkxAdP5QLWhSdUXlpvM2xC
yApv1GBGlyWWhKxUjwa2Ja5nK+e/xq9Q1ME1c1/h/hQCBjrRaU+CORY8kkT+2LF2
mymbEC8HrQslep5WNh2QAeOOXllz+WtXvYjBYifx29nberSbIo8vlTEF2eQD5jPg
pjgSG/O1+Ab5VNVG6wfvHrYjKCaj3Sy0GVinWBCwl644qh/j4wffraDRjzXsvhre
108VYVWrEwYzBGgWC3Vl+RHLPSEE5zX8+yZT78dQOuG79wqYGT+4z/AcllyLe+l+
Zru2WGnPV+ywea+JkKzyucoC3sku84kemB1UGVbVUfN7s997VbgjNFILELu0dK7I
66m9KsfX7oWsYTNo8Bkca2Hb4LPr5Ac37elqh75akwfyJNLLcRadwTx4LuUbx9ek
MG3FTZXTTnwup5fMCpzEEXlicCv2blSQAklfzLB0Lr6PQcFb4qWsvPNdBjs2GOjo
E1Z7zZOXo1Qm3O5nv89eqN61AQI58j1JShZfLb6UWRalQOdoVnQbvZaQ+8/LXq5O
eSpTtogKT/b3/uluOEhTD6rnmG80UCtpNqY0krGzW36OxHZKFRinHmb8DmXbwm2P
oSHl+u/wRtMbDHqKJy1V0X7z045HbDbiUHzIjhRUWCLIpO59Kkx7UvDo0C0xsgpN
9Kgxxml3o+YtDaURok53MG/IthRBDJ9/aMD8C74C+ll4pTLamL3PQrx8bCGME1Tb
5iTLdZXC/NLFIqwF74rO1sHDP55dxyjnW+RKcSRPlqHrpnqzjIe8Ts5vDToRMm5x
b/XK/+xIyhDBR0lyWWmIPPq5qdM4HKeevFucy68n9+enhinT4+w0qSEFPnyzdTb2
RYs1sdhroWzPZKMzX1IIEa6tVqak3ySTPPrDy1OcGPG3pqF5SYh9b/zybYbZsRmY
J0hBhDtrL2cPz6Ufhj2Oowmr47mZmP8OEPJVeiyU1h8SEi7NRP0LdIc9OxgMOm52
G5JSPi1sXLROSDs0JgoQ1Vef/RhKpq6wyw2AUxM5Vfp26dyxmAxYJ0jjMkBxAexM
fy5jbIhuuviXt22AwFgHDSp5ynfKvv4n5XPUrD0op21rhlkK9X0q88jFfjXZNECY
V/j9ZUYy+Q1tKAdBmW7cMI/8usSBpEVLAlBVpuDqcyVnghdsiLPAofA9Vlc7fjwE
wkMhS5FmoQE6IqsZnDZM8JgpT4LEihhGeUTmH01mTztyusq1UhAjmHAANY4G+F18
LRlQ0nx+mdN8xVTs88QBpECvkktDWbvP2gmQH1bFam7nzSzXdKXvsg86e5hEs5fw
ZvnSHNlq1jOi6fb8gXhhbFcBDrkHg4k2eO5EIjxpsm8vEU2P6jHvvHw9wg2rPadG
dac40qtRDME9bk8/FURDV4lffUzwvNbJRFFEdhanf0w46fKJkXQSnNd5dHFQZgy5
c/8szkXWsJY9dWMOCtbpDI4B7quVDS+KHgrWXHJi89Y0JizmWLDIoWMdi1CA7L/o
jtPg9JnDRQz9mQbnm5w/Qt1XqOlU6gYVZ459vVi+s0nYP5LFXOPMtHawSC9DULqY
k+x1fH5UX4VtVlA3WDU5Lm29YIJPmUbgcEWhcU2ori/z93qkVTdVTHpiDOFKxaGI
h9jqQD0o5rcxcW4Yp1roAQE80L36TeiO075ptDnXBXUaMh4s8N/1eiG9VtsdcjBo
ry2fmfxaOiENY6OW2bRXWF++bMrA+mWY4MWC/MNw0PhqAuH2PiEnCEcNNVUThZCw
zF1zWWA1UjiVb04fGZURuE4/PV1/V7EKSlM9Uh9f6fVfwE16QDgDkrQyisOZGlfy
sGCYEVcAwnT7fFQoyRn6V170IeHsqnOqc9+PnMtRa9AyqHcVvzw7W7jDEmie2nKN
ai1cFUCjJC8Gfup+XXEfD90CKx0NVGOsmCWCIkIKZSyCMV8QHA/A6W3JZMYTG9ID
lCnpOTxe6s0AWb3bsDyUYoL/WM8b2krsBmciKIYldhiF9I891ZxukI44PqjsgvOM
PNyzvRrnME697aT+msJU2ZQfI8XRDEDmkP7R8PNIoZdpFlSajwTusKjemJuVILdC
JKrT3PdzxUOGGje01ecYVJWIJcDFg1ZANgac+KOz18hCUHIz9cPeLrkOc0ocQ9Ti
YU075/ysjlHtSrXmsXbM1qY8g/F+Wxdo3ilfQmTqOgRWPGVSqhbQGYEqco+ntZC5
S8NbQShVLSHtpMD7baZUzVYhUVhPXZa1X3Ggcb/2A/S6VXj5zEN/pJ5/HYxzBzSu
DyTpsA4kdH4Cf2thYwOtY1DcetwqHQaJFxHlsfKDXqV7gCBSyi+BZJFUB3AFykg3
1XYDByGulTFkDLGk5pni6dAaR83l5ycgavJCU0YutA9B2VYwgWgOIfrjl0+FXJo+
FaOqZ8vCTX8Mxj+/LOO6qZP4z41H8DuZQE4Kr0EmkVD7+vTI71kWQNJkq/LcwvTS
GioevnU+80ztrplRkFYmkabSKpyDT60afi2udewuZjcbbHSTBHvfgSV2u7AiMhXm
gTpBXmqvJQ/vEfW5yG0kJzFZWnLclFiBNpISovAAg60tg/NGMkkbQfM9XMpKsCK+
sUh8uqE/Ur2q68RLOH4REGGKJw7ZGpPO38cf7vMRYxZ426PmF5i7MzVFlhQnXiL3
rkX5vnZdS8MQiNQU49TYx8asGW+XalBeZp563D7VAIAThoUdUpTtlaoPsHIyvSC7
SSYFc7vVKwD0Sut1xsJ7U9DMj5jtcvugo1s4dvE8TM8SkNBXH125r1FQVQuI2V1f
fbDFj6nBfTz4CqI7HH4BYPmFwmp2iswMIgHwxMRgndES68Fim9s7txXzyCb5Q1Iz
pPCRGw2nDUEHXsiBCzOBYn0IFoNIxCDsuijNaTJ9kvtPgIGXMGEAenrV2AU9YqWf
/E6lOl4UrtLTVgO1XCnhDWKFDx8dULHRWCV6lVwhTdYf/ErrYrvkhnCAXx4pT95U
9ClGoIoaVQDSiMPW7Kn15HM10AuRE9uZGVq5zskBOKH+7/Dqn71MOVP83Xs2i+w3
P0G8r/vNT0jqYCAuq79G+dibMTjo5YZPDRwLk+1tyPwDSMHT7IS22B2tijtn84zV
a3vv/Z1WiagrjbCRYBcrLktYLdsaiTjKRWo3RZz1z0Z0Q1AVi5s0HSuq9aWAXOA5
9WA1c+2T6UDVbT3BugNIxRlPZZOnEgEvcvjjSC5pUQ+vsy1Ng2k3h5bc7AV0ZAqG
o36Y4x7T7YcqFD910LunfOi2WQ1lewEHexzEi3JAfQLZrFaQZasbP8GftrlyqnrO
cHWYUP9rE3ktSY6gDnCkPf3/T5IBUjLvglnX8rLz+ntH14SJ17wNpbIY5iMVs0OP
HUlU/LsPm8EJz0zFKOztMSRtpU4ZQkOcjjwFd/h0VU/Xb8itE0bcpkMwJixZhXHN
9u8OgWFTTQim313W/nXqf+QIExDF2B/3t1pTQFYoVEtbGt2i8k/o9fOW8+AyWcNX
qx50u7ST3dusVtN/cdOKhOUgTDcrUp0J4LQC3pqdtcUc7aEBjkd6BYCRrSLB1dst
ssQb3aHe4Ei2+p1rT+5CkMNdQYRcjd4orQ9YbOwyAQNd8HuWcSgt5toqzt7ZeIYt
3oaAfJ1klydPAlMJAgVaE/DdKVWandYZk5ZtNiAhqwyiVv+lRMEXTx5V9TZCl8hN
m2chRciScF3lXAQDnDWDC3WfXq3qETPD73H01UbJLW9s8EXBF+roCoRTglhiwIY3
zqUqAjC+tkTdW/vXjdmpLjVzbjnRBIpkDGN5D8DUwRYow2hNrAZe+NliptD8S4Cr
R1K2803bSID26B1XG9Db2wzuVaivSCcpe2QqXULHMzj6mOXou630bV0tbXVYHIEk
N8U3juhs+pM4jKuJ/qOcNBWp2KXUwq5BjNHNKxzK7JurKAWF4USqUS0xqRFiSQKS
MY5t0dMFRIQBFZjDs6VKkfThhUQ6eyLt+xiMeX6vaedeTIpE8X9UhgVqC8srUYTV
XfKyd2gsuRMAJ5XX0Us1oB6cOXpCodU+rzeTkdWpNVnNMiR5+0WvceIo9235cMoh
/OMlzD6GdZD7XXxo/sUE3jjBiQ04RXAJA07u7QVA4mJ2QhQLF5oQDJJsvbv2+V4K
+gIP5Ua9BXowEwmVu14jc5MxsGFoRX4iYgM3RDXI3VyrAh2oy8P1IaTounQAB8XW
2l82f0TAiMaCEDvbeDdVxD/Ag4Wo22mq7H1EPjAyunRvchE0OJsnRWCVCsux484N
DtWJkFI7cqDmJ5prLj6CZUcnRBky5QuwXkkWQSQmRzIV6Ios+CmCodvJi/Gh8/U9
ObCYvK8Rmy7LPNzzxUZDg+WHO9EPRZrWzO03kFFA3DX6KU0GiPVMUac8AhGfDE2E
PCan6TvwFl3Wryh0TTKdKrNSa13C/5aRw70PDqXdnWLIH4hPKwZ9lr73NHkjcint
33e5AioG1x3LukZhHYbZMNBvaSlOIb/5GEKX0pLXTpO3ZhSGq4PFi0NcxsYGr2oK
kZF6yV0FkrrB5HhMq9OtXiDisAp1eVPZFTBL1SI100WnUGoqTItRLtMRPcGlyPpj
rdevspGoIVIPh+dlUpYjBkpXRe5ItmG2ItKn9Sl56D81o9wLhNGUpwjnpuXP4uZS
SZ+hLqK7nODHXFLVNizRB9woYO3/1OetcdFPrFSBFmVB/nMylOpLUx6GJ3iMGet+
X8rd4+cweQgkzRrQkbu1FIVcZf6jIn7nb8K4zKuUpsTJM5OIAT0b3vURWUsRfOXt
ssU6tFE3r5hGAI2eb/04uAHsTkN0pKWvDl1UuAZfLvOsvFKmSykoDjOuy60f+XJa
ColHu2JmEyOvnMyh8/MYNr1MngoMC1rep1fonZEI3mb720Swpp3v9BVYRnG/JH4z
aNkm6nBuU+iGB/LfTMNn364fHWjlRFW3IfTmtiC1erW4i4taHYZx2Bssjum/w0DD
Rwmtv+1gJUZrLCMSLMPCfsc5U6GthCCBrmKY8bMGNfizjkXYhtVhJsvuQpd1keEg
eENxiTsEKh0TAI9axjyEsRmwkLpnHORazK0IwsrgRVa5nJQgtkM1/ec95rnpPlFW
jMAnhGpbItSnemozvpd+bElfmGbzZayBfr5dS52QF77+OEe/urVIpOEqyyEPbt0e
53Z7OcYSm3Wm3cKjMmBaKvpqZTLZfWLvnL498v7iitSF7JrRBSNud8iKOBFBEceC
ydI+vykaKMylFfkFwFUvG9q4natnyQL9Ro/3q+W4JJCGKGiUV8e6BIE3N3V8kB5R
5oIwgN8iVhMm7Sm7YGNJtulTFXNpII4jdq9dYoYtMF2rD6Nf40WPSI1UOO7AvVwp
/YVxhL7NaazYysq4g5/hTfIy1XsjCQ0XjHSN2e54SvBxPqc2+V13gpbYQDF1PvsP
c/diK9temlzvgfLhnaNsp7f67FtOI9HGYVjbTVatb8SO5GXXypxjcouM9wjYovj8
e4xmT+Jw2aArCZ3+vry6JG/yUx3cMXpx0QdlpP1x/7sqagWQhJAJkD5p1RPqE2y+
SPw1WyQEHvBexrI2AtvFrzumm6mIJSS2Yqyi5TQeZOY96aTYPz2TQWNj/LVppkFo
ITCaFS2eoojW3CbzSaFFIfsbkvqc7Qbm496cucT7Bv3PD9pAVUfyZrDNeNYBl1Pg
0g8x8sT8CiERdGtbCRmMvx0KasbxbG+RXvM/uowagQDpXOoNDsGglf/3wGE3AjOk
K0I1dMC2++xJxyotdRnHrYEQ+JsUCSjQepKKZirkT+QEKr+H7XekKIRY5sxkDFfe
qyC5MlkLLrQ0BPmqjZzbBnVOwGNaNV3JVCq1hrdqukBhnVGspRAXscKy1quFkzh3
o2YFtgubynCzagrZMKHbdCMUTS50l+RXoCmGUw7P/7URyyNM7geAuek3UB4MlMg+
l3pa5hAIQlN8T+vO/i/WmAGlbqbR+SyNaxOnOa1yT5lTepT+dxAlq+W80fPhNJkU
jViIRPAmKr87Ek02UYCR0UkkpPTYhmAyOMHY2TwE2kJ+uRUc2TN24dn2C9wQICfr
VZgbAa+9YX8VlsmckYTm7effDTEXIQ1jp+oDHYtd+yIc2CMg3DTWQ2mAHwKzE8iy
mHwFU3yf+BMIVJcBsCYlewGtxOJYsRsPvvSglSA3xJH01KJ4gUN2pdQw+KgJJXBy
lT3orWuo49An4v32Dx+EK3Ccq8zbfM3ZnDxG30fLNaXdUNhiLnA5N+OT0CHVahEv
waItIHfut3dDtPYcUBXX21O/nxi8yfrXPKJiDBLPRLrHJaDjm/fRUJe46+w8PkVq
C6wJJXJB3nP+hdjyQ56gOoyBbkba55a02CEvVf6/ctj8oFKHa9bQ9Pzm8FBo1PNR
SCNXOKt7M5v3c/c7Jwg3gy2MZwsA/MqrAcSBdPFNezIN0d8GgHEHZlyae2EB1EWx
RntGsFq9L7TxKBvIPUhtTt8FZUqGdbRh5GJUOni9lzA/v9f6B7xjlHL4BWe/izgj
Qs4p0DDYFVzCfNAfQ/Gt3U4fPNnJ5z8OQE4qZsSAvswnnAkTDN3z54nFsGTA2+cp
aGb1rjh5zKaxsJ4qgddguvzehL34E+gQF184yG7nWbqDlobEVWP1/kyX5CgKJR58
tm1xTx0vyBSa/Thy/iZx8pjKmuNMY46dM3MScbt+DNosqB3Z81tBMk1OW39bobAy
P/fdiPSutUn0VWY72pcmUE+JFQ2CyPVsBS0ruPxXcMH4LLynTyz2zxstTLd4HAwt
1xx2nw00WctaGtlYQwkzU0iPUkcXOwum/NTsqA8A4rtxpeHUREPuPAbl5KfaSNVN
wXd67Q6h868R0EJfOhUNEwXOQuVLaDk71hu7/DhjCGCXS0VBh1nSdjPAMjgoBY5k
CXOukeX+ZqKUSYFm9fT2nx1JUKqpa9m1hEw5LI+rg4te07Dg9O6GA1d6XlITHzT2
PqR7Jm1oAGXBB8xBVW5ZHC87fCF93RmIuVCi59h92aX+YMqVIyNBmsE05yr8BgAj
o+hVyuADsH6Z7lXAbJqCujN+E9M6lLJckaXR+FlEA0CcFn0AAnoPX7eqkbZTrZnK
TLIRUljKTA/h59refYcap5IB6Xdh/5FO3m+8XTIeZss3fUyFxa49RnqrxSkoCP9M
EDjD5a/rJFuEATEimrunzFobo0d5KM8ozx9AQbnYMezXuR5Muq92l75DoTGZqWOX
NWdxtjvZp+W5Jg2trKwTTLzSOv2pgqZdHtX+TKGECMtYOjplpSkB/prfMWoa8Yrp
V8VmvfYB7YNscyDtAwChqgdqSjOscbsWppvRDjfUARbIejeUce2BN09hy9Wk092N
GylgwiOaWFe9W0eN3p83zeiznxN2pV841bzgZdNW4e1IsEyUnV5cf6zFQDaqEegu
37YyzrOwKAOQuTpa+O3oMUD5LfH6UQIELzRahe4wTQE5PD20zbj/XvSfV2LP/+WK
9HRfYBpp3baj1lfQyY4H6KBnYBqxXUQnUqqhC0io5utz7xD+/jsA6RX8y2jYUKMe
O5MERHC2TqYwNwRJXI87O5zVn9l4M5Nh/TRc3GoPO+FnOOJbyAE320AKSCEF18ci
cQ3ZUQuZ5AxfER7nATPNo1dZQdICpnG4t0NS5xI/nvIKBI9X2CywtnxZiwxjiTCV
+4/KGFy/QkPCIMsLcxXbFna+yY8Kc6CoNVj6nlgIRy36ooFu9IL5hrnvUaLVkvzr
OVkytdxel5WZocYW2QIoKPd8r8NpjV1vjc7yfdxKf2QZ5N1tVFgM8InqHDV8U1cY
xfF40irUalb+8+uxumssJVq9PL1B5TCmqvuR6fjQgdfYEOVp8/Zn2p42RQSn57LP
Ec29k8KZtICHRvX6IX/brDeNTYg7JQdBUaMhXIEfK3CW0YQ4eTuKmuEx6PyA0Yef
HlwmZj64lZ63GI/76ZFhtmDLbZAEt3Y0pzAKLMBVjrTiLrqZUsLWqrqB7Stcye31
BHLsPh8EcDRowj4GXD4cZT4k+1RIxJsTx1rI7nnscTBdXw7YDnSh6a++3fxAs9gj
vYV6jnGdvV6w86DBiqypA665Ivv6FBZZkPmaOknOwKNvNwoGoSpesM4FhU7kC8Mr
IXn4oy5EPb+v2usCIoxGyVKpyV/eCbcVhJ60xepSrSjH5r2RSWQC5l/MCJAqIpbK
Am+rehsGvpdzIr+CiUAG0i4bO4iXOJQZIudNIsnlFozLdlFRj+ZNTsBHJ0zDni1J
VuFbfaMdPFIohODXbUW+Ve5P1unUo90Z5A+DVYbmqXyE2JioJkKEa5l0qTr6jV9w
wG6geO2bUMPy+va5WCfXal4r5YR+xE73dWxqbf1KUjCNHkHU8PbHKMjtuSX9Q5nD
nxJle7FJEov+S1a/6sK9QrHfltefTehF3IMa5p6oU9fFMIQRyWdOXYevGNXedO1o
qAdNoxXq/G6GN17TuR3O+dcsJXwSLJRVD0q2gFxRqDoDQytSydSpzTY0Z0VYMHfX
K6IrHkCbwexaV5TPBm1z+5dPlk5vrrckyQbj+GdKQNRR6iuPUBio8uz9iL28oYzH
USNU23cI2lYHuIZyKLVR8ozc26idz8LqoVkZ/4MIK0bcxs1yUyPZhCHhennMcMzy
nOQcUxr9b0ujROz+Li654PAw8jUWYAH9e5e6k+FPVr36aJnZvhm7Xn4wS2L+B/3p
pVEtTu2GuN7rC1LOJa0r4YD7ZlQMEHViJzcPOEJP+n8D8bwqJJZ97ti7TQBBbwrE
qPP6CLsRWrcfRMRiLuvzLkvxsEVcxEKxRGPrQcid6E3mHTQurUcsB/BLfvsGTXAe
LMFMOKkLNPraNX58rI5vAA6211esD+s2TPvvVwbEiYx6BF4xnopuDFntkOLJSeiZ
qJo4hAJDDearitSXS7j2qbmgcxOWF9X06fJPCzSJWHpff4q62jMzx8+jHkVAW2Bb
ceLNmvpIB21cmkd6lSSjwBTTHKFypCmLxlxgrlcqcv4onzSdqB+5+gHdJ0gCecwa
L9zwtxvcFZ82S9iX/YoJvqYqKWw/TicavgfY38rf2yEZ+fF+nMCHzBgi7rr3m0zs
9mgZ1tXT5Px9YD7PHCvSIBnmkIT2Ki4Q8+JiwQ7g/QKC9TAfzwdv+7UMEj7opMX2
BVUfZ8TLW9DjpkgaPH8Du/yViLFHFF1EW2vMM4G8hKvhUEhiDRI/bFp10RZevfGF
wSy+lukLno0p0lguKgUxwkoynpNLvEhugk5dPZdxYH+Xq2qwtu0YRb9dkPDUkbPw
FVipm/m/+XB2bh5n/mE8EC7zjH3T+kiJkVQ3pW/Nm/bCgnMcZt+TM5hpINiNVeOv
Hh0QrPmrxcaRHMGqxGUi7eOHoDx09qyzuPNOOCOjGzvL2g4hj9FjxxoNDj1oNZYz
NlfTTVepv6IVeNqt9w/ZcmYdb4sL+QGoTZKCYSuV8/jX/whbozF/hPUcWnWmR5fD
c+u2IYn5aIWwmMhBRBVY5s7x/RbjJ0FL8ivMppFwOACG/83vTlpIlLbewBEfwxWN
EbFYRCpqlsDXwh3YVLKwd1yvpDbX5g/7Y0xu9P10s9AD9N57vrz7mLK7juTR0lBJ
rpfIjldZReUag4U9s0EeefuOTojpXqm6uYykyeYhDdB3yGGYZVcHBW+SRehjR9DA
Q/oBh0yre/+We/HIRhwI1ZEZk2zOgtDVFi/fkjM0zwTdZywzLqEGxsfa4J+peUBV
d9PCmPDJOZdYFNkcWGnT9wgw68bCqDkQRbYPhL3mdInHKNz8Ze4bXcZn7PyZ9I0u
93bKbpjJtGQERKN/+1BpnyOTbj8gev84OsWa2mfj5LL9cEpBBnK7wVBskCylB4r5
udvgpXQ5GfebDE0R/n6DrBOxzCLerJV/szBISmP6IXjAJnmNQin9dGX7PM7kt0fe
eFDvFepDsxnE+gy7lmoIV6L3LGKpfBAP4Kmn1GrCP8YoHDvdoAaL6ylCxAPIk7bu
3YQNjUWLYEt0e5Xyfy19+WlPkWqyqQtyGimENnNIvbbjXISi6oGabuZBtVFEsTZs
MfjHEzQKt0hqS1ZfrhcJttcJPJ92qEei0kkeRK/mHCE5BzCAiB4Y9NgvaldE2mjC
lowm5mMN/oAQCC2L+idGKglKgr7J3mcDAoqzYA9pRTPeAeIoNriPQwr05zhsTrFP
uqSjAT48DIdbPKXoy5TC5xhm/7GJBCFJDG5UeZW7/76NLhptFjBnmKFFP7hQ34I+
A0P0n9VxKm3WCUILlkLfcnFcBoV34vTstPiMD82n6FDZ5+ijq9ho02v9vZCeWrY3
tzd6QyePfkeI1VdB4mzAn+QbMg6sQ5kGsa4/JqCDvInvpf78NTmTY2xUhwwIM9Nm
0ic89Hk8bSVoMNEjP6lhxKTT3LuLzqBjhjnbQNQR4rZ1bKE0YYtgN7YjNJuWYF6s
vyqKG/vcVmqipDzhd/jRUpyGFLnP4OIeWe1dJuejWZFjAeyHmnbdzBVQLrHEXl6l
ZxQNITW5PV7tW54BQW1nhqmX462oeZLd0KOqhgIv5uheyH419jY84fThGivHJ+K2
obAe/MJoCFomL6YK7MpyUlQZOTkHhBVwRLZx/1gFbiqBsmaB6aeHnqOV0I74J33d
noAblAiIUnYGvmOeWLYdMtnWhNRO8/OJ44xRfzd2obXSed/dLMxE4KEHccu3WO4E
ytQpjOg8U3QkNPNFyLgcEJx6LtN9fxR+Hjv0fe1OrOeI0sPvBf35iAw49wv4aLY3
09MLnkZoS9JBqTIsEn08UQFHmRxV0awczDcJ/trX23bq3S2w6wxSiFGNOiihZgG5
xpkEY9tMga3Cyn0T9ID4gkzLlMZmvt5yoyN+OZhewOIKOrlSbtEHQtt7EcCjrZ5n
lQR1TFLBFAyL42uWUEIGMatyaKIUuskFRjpidb54eWoXIuCJSJ18yHHaSjKGet3J
B0tCYpzZ3wOvRaqXhus2xGHcoBaW4TTEOO7ggTGdrHp7E+0mtGzx6rsf3mTudiuo
U5ueLILFf5KVdi5YSBT9smY3DWZ+8QQerX9p7bzVdQ3HkGZJRfofHSmGWq2kOmIT
CboWoB7sI1PBT3ZdKkZjbPsS8b/9a7rohd0v6iQW5Wuo9NThOIyB+oWUV9xAJAai
H16Vm0lyhn8Dm/KHJZq+WNzeiE0jdew8HXuVqG84BSOQUfgy+I+KnNJak9+m2LmU
aCeq6Ys9oGrl6swE1LeiN9pe1ZMjV8LlLm21qwPAEQnhUefFkhvlP/7rGeBL6yeT
keKzpap1lkTDurhi18keKrjqQxKNMB6ZtKUakTfgCKrq1xVr876t6B1rB21JJB4L
NKhsF1JHbXRW3FYnwFlOo5slW3YyadZBD0aXJEjEcZda0LodICCpKWHdLbzKrwHU
pZVqwXpcXh5yhapzBmAettqMO6JhpmyQVIrCkbC8iihba5H6qmYeHg3oiW0fuD/j
ay6z8RFxW5wZkIIoEU+yg4bJHQHq7eqQ9yjROLaTaLu9WEAOy524sMjctFRoJw/A
3k9dmUnQVUd5Xq+x0+J6U+94THReQOCerQGXE6usWchyqz+q+chPoCB8slbOC7B/
D9BNpgeoJkYMhWuaUZlo7ACpb7an58AwDWoW1Fq5VIYrhOclQIa+pgQe0ZGXoeYd
XnqVDe9l8AVYSPxcAhCVfmbztz6fjY5dhkTuheCvi641u7ulo4uMNUZ2vGd00cic
+7nO+N/0FqeFWGBeI3Kqdx7Woo3pBzR00eo+8mmkOMjdpGRMs035UmjUcKNpOed7
pmRb3zzwidrHLeKawrfhj+EfKCbJB4nlZnmHfbAvMHJaJJuK8stdhUM1Lyr07j2d
pjMFQ1zgzHUAkZZVQ3w1b0gVM2NZAiPgNY0bMbMShJS7VDmwFoJbADlewSfonN2B
uQyJ+INVLh0CgXDHw+lGz7L+Jlk3kJVB73V9GOimD3SOpeY5+kQqBJOZ7h+ydRau
P3M1Q0vxWHLM5IYwP0Sc5hn4lAvHCZ8dp9W85GYBooqAznqXkxDPTI/xYozPcJCP
2rZ/cCAp85uzKajdtg9xeUQ/dcwIu+3wdnQGkzThjIWW9a3SL2TLchAQ2s8rkBGB
AehVFcBwbhY7jTT/dL9aOqxMLsdmpGbHckoNqfbJVPOrEVXTwIw/AHlICRcAAAJB
lRPvYYUC7qu35i8Vx6PPJulBqbdwWvYWxChEvVPChT/nTMImZ8jSK2WOIqEFGDBm
SPfqJ1Ff4MVNXnDSwmgFBdaxH/Jx7tngmShOFhwyegTquSSHDoWkfHDI1HIQl5pC
fgo+S05lnG/Ru3Z+CkdLUziPAFGSdcdsK667iCZTgweXOOHPPiyGJwnjicPhOz/Q
bI+jhb/dtPSK0c4eIlFXDfjWI1vHyGwuGaVTxgVS9J38aix5nbwCYeZMNiVtbahO
P+AEm5giCNEZpgwMZkDtk+gxSUPyf+pZHLkZ/kO5Ep2toag1MgctXy9ZAB6MBgAq
CMbNZen4Y7vxUAA6HQ6DT7h/SIjM7G9eh39gEjsGisU78Ouahg1XiFZgt6PARMvc
D1dxoWL2x9zAlTi6WkPY6J8N70hqBHUA/sOy1/gMfDtDtJ1fZ09XDJz1ctCj2J4B
yvQyVpZSCbHAEU3fdbw/7sVrorleuDW0OLSnlZ3YRp383WitDiiGnpcZav6SWZ/0
XlnsupcOwF8OV/EUTSMm6NE6b6I24r0dTzoDeo4/mXehalXq1A8sJpVkaMEYRfl4
DZGzq88awqVZkK9RoCQeKQ4qossabZli3NclAeOL/XIYoE31ZhkiSD/bhW37gAqw
4dLVkHleLp6da2HRsW/4XtsVzvhx7lIWn4gA7UwkhiFCEWnxytRRlcurDFzmyCXh
VpslCTJvPqBijqKsg37IbpGAE0Qv2eAqJ1iEbpeHZz/dWW+nDHpsrsA11rGoW10G
/e6QHPqEygyF8OeiOQQnQ08XjZ1yQsW8yqkzgL+UuJt55PoPAYExfNDKoL0zzR6F
OIYiPsACtneg/i2YC9+qW+SVjZgtzW8z4VZv6ikrH2EMqT/H6r39I9DwVdkJEqkn
ffQR7MxBq0xXLN4fnT3LnJO74tGapxxeAqKRiLD/DqMtzVov55HMBgltvGMi+61y
/OWk3jO/yjgvhGmZo3WrYU6Z4+T+nTfg/DHK71sj7lHbfr17zdDI9kPcYfyM/0RY
spwPpHBmcdL2n78PWD4SVeqom7Sfl1utuRBFFtjGg+rB0A9wwE05OfzW7ZJ4eB/1
QE9+iW31xiHo85+CsOPLhqZZ1laPddN15HLuKK0XUNVNKGEMAFVYXvqDODNjvuBK
SwzLiqXLuG04dr5ST/OgIBHGGQhg6oakSZ+b4Gr7VUCw9QdgltAGzdRpSjIpml0r
suxUZ4N2Ap1bRzfpuEVpmW0TNgtX00u2Ku20mwIvo4Griv3pRA/Y9mGVGiOqDthv
p4yOF5CScvm9uGFXE9hGAhQ4MqabsAD48NH4ozMvyty8RooO2qI1nBY7Ow7Og5Wi
FnAuTQTffR/SVuJrTcIdAdDY9JsCGKNKEWlR+wjbJY5rPSybXPP5P37nhzQU1LY9
Op4S4dTD0ITdxZmuYyNhJ06ttUXUe5FIH8oVaIlC1Y3AlN86GEMQxqb9eeQ/ouIr
4QetHW51OccU49DUbWRLGNqNJbSeh25sQCPLyJVwDHHp0lnrWdj98Z4XABTggAr6
ac5t2rRUSilzcRUUYvnT8O5OWYtSFCOFNdgqnyS7Nnj6YMoMF8rlUYFUevpnhMno
ZExHKsQ+zOWjlkHzJrk+9Tks7p5KcMFvymNJXcYajo530BKNSlDCk8g6ApQOx/8x
WZwNS5QEwTGNIForHQO8l6ZoBeqIVd/0yqCTvgtcO43GRmTT4hXI8RtlSCBb/6eF
O4zjtPLMW+MwN/4JZlzoQNfZQvzzFtGUcos82GaumMGLz5WBX4zSSsYNpVyu2ZRJ
G/pziENDtexGQWUe9XujtcPXSfWqQ2KhTp2VP1yC7PUoo6y5BG/UfLfzUBQ0q56n
+iXR0SY+XS3HytM7we4PKo0Xh4cUc7Xc3ESqCXunBLRRtwj1molKwfagOOhsxvwo
UhtpK9fyq0zX5mUTwkKw5kYbXWQbr4WqgD/ylB6dxUZOTc8yCMAs61KoV2JHhuHW
ViAyj2Vk4eu3UCNnj6hOqrFO2N6eQ3V3wYbqV5YiAVZ9vvvfH/jTDAstJX7aE6B4
P/n8plozyZafHvzkK/px6oWsQ89k9d9Yeny+TLCx9PCievI54SwLpmSNFl7JJUDR
nXBo6lxPIU4J1IvYfc3zRryOqotUyLSgO4nlhIeikGzBRqVvkDptF2ouuM0Y5vPq
kAV6o2bJX6I90kswRAzgV3ENZJuPCw6Wl4vbnEKZTAAzP1rl37U+YeOpb90ypCzn
8CahaKAYobfJSd+u5nHSSvKC23rEDPkostT8ERgNbL8y/KguqSc5hvL0egmwjKub
lb3dDvYJGKLiznp0/j2w99WuDNFmxdoidA/STkaaf799ndj34JrzVJX3UN1qOuoq
ZQJ+EPCIeFkFKEI+oIXnu2nnvKkC61g/P+9OZ8wT7eeaZEVu7LaeCsnUwPiT3mZO
V48ph0iRtYZEgAR0my1QYawjRJUK3Z6h6GDm1RfgeTvi9PCIttBj/NPZBnoQq2G3
d1+1xeTRfHfRqU+H557XkrL5UStmCxTJD4h9kCKdATi2Fdbg0FvSqoc8AefsRlLN
16kwW9Yq1R9mipCPDG3wMmBzOZOsQoA09OqYjipxgrTKjuC77by+zg7klHTWNOUg
5ODbL/2HWPAkPzO9YDcx3arJ463F6bm7ATgbK7//idOpSPbpAXHCMYWgNlXT64QE
SB3gxbVWic7HgUq/Wia7Uedlc3b/1/gFbH6g6Li/ENY6zt8vvDXFMGwo/DAna5Jt
h2jpl/07Hk9fKGw1LZwpUCxnn9oamqDJQ3L07ylnjHkwnkNuRrpf+FLQ2XyNsWzh
0pK7Y2iq29DR4Cg0RHtLQkT7pkrCGQk9hM94zj9ko6lXos2t7nlOo7VxHXarlSSE
D5obSbQsGquccEwOU8ZAj/zBlxRvz8IdiUT8QVWaIfH5p3cVBZshqaRWWGBmQwXo
8eV/c4doG97+RlkScJykrvq2IIS4atHYlBPUNRinJlQLjezNjK6l01wF6BAVV5r6
w2RmsYWmEAhiF45P9mUkqqZmGa5kuyZcm2Zc7UQdDWvWHzVWTAHqhCVXRoQHiAHe
5d3NIIm+UnZuNp4aKmmWrnPl286sJrgWLh98AaoZHhccN5iPHYyGzO0CVubU0BWg
XmBLfnsHOjVTGP74Kag+g2fNQX3gb0v2nVbW17MB6NmejbVdmL6LdL6bDiMxHMGT
oOC8yljwks792Pc+5UWmOt6qbWIQpd9GbVdYzA/bdf/AHxe6PuiYGviU56WokxvP
QISnelxMOYMxepzuwBZwjbpJn1WvzBuk2TGOpz5AKp/gzWZ3erw38ydLw20Cpy8a
+fjNS7XOCt59IJNaa13FQnJxqfnfkCZFkGEpm96AEKLTG0jup5A4C5QMWoQTbRPu
prYnvm+TC/01gKHFiQCS/2E9V/uXrC5jHnkZbRKKYGemHLOajmyGwp4R9V6Yw778
e+u+zjq2K7iYkPiD1jMtSbgYaCdUVrFXSA+pdsTwRJy+xmSbrChxzC1w6hhEYtMM
jqgStJNjuLEKR3Q0wjBK/IaFSRKTnoJtGNuLVuOXK6GMRfAtNJaUUWkvWoaUBaDB
BlsPfv1jhkm3pbBoszIj8Ta0Pb1GtrjMy8lvMHYNcSpZ07+b6agGHyHbuJQYourD
9h8gqeeKLYUrdfalPJKFy0NYyLRNoR/NUy3tB0R0IK+kvPYIYvKMpSbaZa6/V2/C
NlmruFCGyubLqqy4pUZmQG+v0KQid4AcMqEmnZV9nlUroW4htRqC1jyztFpwMd7H
ICeCU4i7EPc24z9dUH1eyMri8SfWQyrW7iv0i0IH0U3RG6w1MqrZ7RqdPSQxDHU0
oej3i8J96+9iQblQNR3A/ETZl5ujk+IEWCZz3XiaNQnJ0WRyGqtpu+gU7fJwqjeD
3VGcJSnw6NXL+gllpuvoxhZN+EGmpGRWFS8EtawPcAlbTHlJkEe/hmVdICX04NVv
nO69CXfNeW4NvHgttFWO5Bc9oDJGXFmiTip7b7Pqejtp+DBt9bDGGyIJ5th9WlD/
cg8Zo1N+84N1yMKNKEr6lrLkjbbn0GehLbpcoIFUtNvG3xZF1BmhHT8ZQ/TnvJOO
kLB1X6v4JitF8Q+TJwNsjskkbFkmSgxF1rk4uWifVfCRAmtimtcqUoFh5FAN5+pJ
4P04+TaVmMeMzoLtjRng0UXmPQ8YI7++eOUOXqh19+p0TDVUuVmx104Sk1XpRrcU
pHWto910CgLSVxBVXy3Ct68J8hffrfQzT1mC3asntdUuKv9PI4N4+yJURtLDj2Cz
r0eGL5Wr+K9KCXLKQGqCKnseSpebGaeoFa/XFR8a7+XMV/DEXULtVwkaXyNzS8IS
4dKHpGCHUs5DAmd3zGdx0pWzfrjx3kTDUfCD26JJa7A7VTHNrhMkqxlUddD6obLJ
P8Ygiequ3Uge4SSC0NpcbSm/tHLKHH0sJDbmM1KPak0+sqMKsme5iaEVa8KjNjG9
x2ScZIPW7r1q4xxyFwKiyC713RAhuni6uJpfhVhShyYFKQvgAd7HgihQUl4siBB8
pmCdSiwmgegwJ9l5ZyQmcoMUXjjvrdk+kWwzuXt6Va6QFdVOdI8ZXksmGDjo74Wh
G34oJe1AIldN7BqAyY0vy2yotYT3QtWqfRRCqMRPPnVD2Uc8RyTcMw4WGrSf73qV
fs/ur9UB3L7CO5jVpkHRJr69on+ahp8hNQ4WxEHqJI3s91NFWkoRdIxYdnZeS/p5
5dxZB/aUT1FQubxJewmhJZ66ItEuksn0sl9CFbvO4ktsRCI2NQHxKB3VUrnRFTa9
xyxFZEZpIctD5/pgZ2JNKaP/yWhLK3H+FiqLk6vbcmk8lB9Wq3X712w9kMXR68KD
FWXvXWNZZG+0c8IkFl/YLO4QjSnb572UZkXw6xzqGJ1ZUIYTuKeM9pxoykQ3OA+u
ln814pFTMrXn9MM4sr3uDxBH27q9+8w/YjXZLrJPujR8PGVUmW+DkWy6+tUIhsg4
3oqJR6lSvyM+zl8dzk8QtZHuKC0RxDA35HsAlmZBZqd4sr02bRv6wIJ074c9GZlY
g9aEsu6DrWyLyzdNUuoohsmCpCLxkOvM1sgLCRLNrVLymKp4mbW+xSg11wxTwYE/
Lg/NQeHt6moG5fr+ysuusx8/e5x9ydiitAdEK1tycj8FdzbT4hzx2yf7NeXUzQVF
VQB+NI6u/FTLdJKIIgeoyIo34obYjXI0ssJQivObPAsBbQ09U8Dct6SmYtZkCPTS
jHvZT2ooeb/Q2bugzfKVckh9BrgawtU1MNDPNb1q9vrbfTOERrUP0wnbCdMOOzCm
UfdGG0+wCPDY8V8JyAyAt9m6nNnizSHiBD1Fv8yZLuUM+qdLWHAIglKvsvM4L9Y8
+Bvpf1RZtXr7gx8JhM72zqhciD2GillbfJx/jHHKZOgr4juNVZefJB2Lsia5jOan
PMz9Lh5jRv+iUduwUJpzKAUF9XlzwvYc+4IPVw7p8dcsuMgXZupG7+XHIP+GyVol
xs7rFfcMV9A1o1ZSW6ln3vpoYTOnDYymiUxPoHQX2KY8bJGpCS3qqoP0/+fv6/Ya
JSHpIFKvIWWw3BA0Z5ZoCGPohKoLoI3Gr7J/HQVaVsyHu0wZg4mHx+5rRkms4x20
Ooj3sfJ9eyRAJJP/Aa/Rhd2qQtS58uelyV6Q+jx9XNR2EG1Ehs+DP9gZtAVg9luJ
wzW2F73E9fcteIfnYjleJlHhybIOASXjWKYxSZEX0ocuWjHOuDAxfI8XSc6/DQuh
/t+4XfSkzFYn7+bI4Sl0CD/TmNa4F0Zo7xvnPpgMMRySnEizO68jwZKFX5dFVyDs
GCaQbNDFKffXlI6dzCFtqgaPLmV4t3kLddPd0RqFu7SzsLq3opzebQEESQvjMHeY
BXjUshC4o8RBQJQOreik4KeIpS/gD1evmSE5S9gHnSeGHmcQVw9oxPTBJXG5Wuvf
o+Jd4ChVLAP2/ct8RqzR8sl2GbZ6li6TWFJ36y46XJWQ/tfk1YVMKIxIu1AhRkaj
mxAJc6/qCX7bRm38RwQS2beBxcjITYcsUQ/cc2JbFFSzXdcQ6TiD+sWQpAU3K44l
bcc0CMnZL4oGA9tshPpHZkj/zX2OeyuPZdYGaAPRjtpA1VTr/mzCDpEdqDEbEoBZ
IDGJsZhGMUn8JgMdlsKJoX+taweiryGSvyxUs2sQqabvKZrpkzz2RLL7MePt10Yh
waaR+pHbosBhzWuYPbiwdMKW9tQUo9M2dphmj/woXLoTHz2Y5nKwb/l9r3jkMcsY
HTRhpZ/FNoethsq0nLZH+LNeAb8nolZ9joU364/TUhIWiBqaLRolt6VtM8ujqCgd
o0eU7c19eAOc/i2q4Gr0C6dINbItuntxcMEV58NWk/nJGK+YMQmLR1LlXrSwR8ra
eCv/o483DygflUtfeeXMtV1yXhUfSsrq7ooWqE8R7NLj2CPSykwdbuWoD5ASG9Fl
RsCb0TFIVlV1SJKmfjFASpFOGP7pPKXW3eurue3jQtAfOaulLz9dD7mdoZYYzZW2
v5LFllPnIflzuaWeEN76aZi2WsMCBHShT5oCmoyHX9pZy70pfwYW3jk+gLLE86im
abR++Y7xAPya4LD3gJllGbYBbAT5uN7fx6MwXDbhvbD8KhZ8knG5hDJSLWDOpUsF
oXgknwcodq+866yCzdedXJR9kpTsI5iH/KHt+xxHOSb+KjtQ1JakuRWplazx4hbP
RSCusTuWSzgAG0uEkINkU8bPtuHLY/YGRhjZbdYm1fFBPhXK10EPM+o7ZG6u9i9N
CcyisjPoZMd0o/mKOWtshOg3XIBRiwL3CpnH17e3ri0I0LUdCoH8q3q0lzT24nVN
h4m2gWA+uHaT57EiylYLUZ4lFF9xcsdir+AbPlWWyuKnPuJxxl5rZ1DPckgT+R4O
L3aeGBcmBEheOtEua1ycgaqBOpQ8UtOLRBEwKZ/n0h4TVZtro86rlJcEcYAjYhPM
MUcSuW9KT8dZ06kut/O9erCGcQ7hh3xe3DuFm0gNdCFkM1QzO6s3dajNZf3Nv+Zi
wh13Unh2B1xH4yJYtxFtI5qEHbH3YBlLyHRxa8AsEAMVS5j37chYgyDF3cVvweOK
LC5bYrtsD4zeuAXLz3oQiCmJiq41ufvRfRJut7cp1fZjn/w1OEhtmkmUWiKD1CBC
kvf6P/FEa+v5qL4LHPi9dULjS7Z6nKrSLPhuBSBp1H4W+mEpiPjBKUrP6/edPAl2
qJKq5tukieVIjXDDEFtP1Z/djeSykZ8OwAI+y4dLdj3AoIXZu2SfCZW6KSuIP8VF
fdkWz7HoxO+2BpJ1Lz07c32DpXFcYETBwGO4JTK2deE7+NeVxux+EmaKLbbgqTmv
twc0eFbpZSyw79cmXr4p2sAr8lLOgOWTNBItxplNLsUCQch5u0dfAVI9MMnu9q9e
K2Yhk+UZ7byiyuqq3ukvpE+vkk2dtlVj82O4/uFjgUkJG1cDmHluyJBrWdxEqIZn
seewn057O/6a8MkpZwfZ84lcJVMstxbrLdFkVv6AmWqSrIbJWzXYD664Dj9MeqoU
nUeuTz55HPBWZHRQMTbzJNOYUFrSyjWmDZL3RjQ4fPFQ4ccbIXFpy/UDacT6gpV4
JP87q++Rv5eFKypodQF+32CFg1MtZ0EqNpG7wYSTuLQPBkI/7Y0yNXTzodF4oBqo
RGb8CXue7R5b/Udd0dqmxYG2m6xUSZ30xJrJuaF5z2C+DP+RsbknEfYYA1pA4DH7
LRYR5peSXMysAuDGePRVJaXKeVoicpc6jFkXnBuBvU1dEHj9CY51pJoOvCWOr09f
1x2Dr1Thq7Rx2K6/pAVjC4PuC1432/HRQuws6aSLm0wDs8fOyLuhjFGVem0u00cJ
uVMBmGaDJiYYDaRY/ZsX+sldY5obpch8IJJrxjCSOT+wupwaARtZIk4mzilTGlFe
H8rhOTgN4rhTmputMbZ+0wAPV+45THFPaDMcJbUFIMZsLm7jRtme4+v1gFe8MsF+
gfOJbOM8ogJ/xReAWwQ6v2enV7QvNKAcBJChQOVrwPhgUh6FdI1xvco68QvtkXZE
0YWI+Ob/zJP/u/l6bXm97SrdRWsO6FdyQmnmKIdFAwvSwkpEwewIk3kXcdR5wJpx
jmIiD8YCoUsybwluhpJOIhWNAbwwXZuxgRf7mBirX3SAtlvEwOdSUM3sD1z4+Ksu
k9mi6L8agdy34MZTaxSosYA78RnuZaSJNuVT/alJFpjVkdoueTPO8mJOCFXsB3gS
+gDrXTKXgVHCo3Xb8d2rgdu411QmTpNQDKXAzWDCm3T7ezVF1ypZCWMgIw1t6GdQ
SXmu2wsqhijNefXrxO4FgaGF3ROybyeoxv9oMaVeYNo5S406CFSkUdW0myzNFxsG
d1xASv+JGEXGL+EQPDd8YwlEiT+IKmkiWBer9+L+ZiLitwLIdRE6c52HYx2nPGqD
f3nyOKDXpI0rHkBEm047sZO6hFlNHgcFQIKhy9L7tHfH1piUOqs8wqt1IlyLlCPs
D5TUpYna0iLmLl5safdopMRGqv1v4vnyY6Ov1FYLXiizWHrVW1gQy9AIYzG4b+os
KwgMcUtS1pn3LIBdV09v8qX6MU6Zl6tFMPxPdPU7JcqMg50noqU/GfGON+P/45ih
ZgdyBaBGzYNyhPqQS4r7vRemNKd0J04o1dakb5HQDWaNptVBSxlBn9/7/tzIZdWP
8nfJmsvIRexYBav4j8/ASdX7vMuV22K2fr6jowjX2yLN+MG+3nAd8t37Afk6s5C3
GAywNs9ZBSsrkHWB/43MRJMesIVJu7e/Qsvnr5U46kHlkD4ILmozXOGv9WoLhzEN
nny0lnX1Ovl9YydwdoJR5ZDLe7BpD6NynShlWvN+VddSqHEYkAnK9ipDX8Tds15d
uRwN2KtTE2IGaSCHQt2s/Y9xyigxv1DBwOyyf+oS2/upcNbtrDXHdiDSc1aSYLCj
rhfQzb4MQGvZtgZ2AipRBoEqj+7PN3Di331BTTFHG9Qo7bjOK+FAzRlQKc3Y9LPL
BW3K9eF+PJICl+8SqAXQK/1jy7ez8nyYmLy/BQdCoLHaHUP2FKgIa+ba6fa1Ffy/
LLyPNiOb+y40n8sj/orWDTH6iJCUpLIVuIvJNxqSsct5MbQeLVfWPS4afdzOqPOK
186eWJ/6jqSlwef/kYuYSuIERZ5jp9cqaFcerMW5x3qQktIBvwhpzg+EoLqHf9VU
3HCdJJUza9z7oiVP++FNZ080IPlqmdrM382nfcVFlsAjOYoNyJdQpi/HEQyOfA4l
hr/T2I3wNQS71fM8MdB0bYGvws0cwjaB7Okjq5PvA12cDP+3OLE4IcSXOilq/2r6
M3SX35FkShZDi5s9ziBI8V60hsYGC+m19gw4ZQza1Lop/pyb/G4OQzu8gyUxbnV2
GfiLxR4ASDgal9Un8rxPor5rHP693ciZOJ/S+B4gCpj+UdjHY68BHsKjlPofqWMZ
7iVo22XV/Zsuor/KnxjuttPx02xYQo03z0LXNuRws+GWc+MGOVeTaYkFa4I8jMMH
ITl+sOGUfM9xJ2ZUzMGz1n9i319H0wU6lbxbmhC2feusn3ZM5dWD0EWJSPIvNfk1
e3LEWlDDkPFCNYMRHPm7wqDfTPJ4ugy/vnq0wSBhq3P+o4Fi+hy5rwa/Qh25xhrj
gm7hKIqnww/6+G5Ehg9eIDwBrWlIk3x2JbBCY9tANeHmo0XmaHnC8ss9YvDR/AFt
nS/l+8WCkP7iQe2Zzlckz4kccahqXH/PAaX8yFe+a7XUkoTw7NNcb5pHP+k8uBDk
Ik/iVkOXmknafMfSM8jwQ+lJArHIHZMj2ZZHy73AqsTMDzuwlFEc5omwhSq+BSk/
VYBNZs0CuTP0KAA4DX3VNE+ZUJttgCxAqhKoSdP4Nphv1Kg19+KvSKayYm8mBZZQ
2nj23RdGM1Lugb0aNbKm8I+XJQaIT3TjW6/D5cJc9N1zJEtvHgc6aVEQoh06bSi4
3Vn3CXv/+Re5SBwR2Blh/ewENmcLayN8O90yPxjDRO3Ufud7wJboE24gBTvYDTPe
dld6Al0hJwqx/aNdoRZ3ENMUg7QoAdEA0w0RprW7oB9TINyEF02TDfzh69ErKnhL
xlvg+F8OYunW2bVzj3cNoigipYaHnmiA2KfIH92DivpHoftEfV8+2LOGexkTQJYc
Pis4YAH+JJHaAff5Q5AgN8nheerM81d2zKh+vDCV1cfj9s/pb392PkyJSaunqWAZ
IJhdZluWycyNZ3MZ56p0lCRFu0pN/YPOlKN3KCZPysA8ovSqAuXw/+AXwUTYr2Co
bZm2o9hfaPnM52M5UPCexiy9hBHes2jeGbQRYTn5fkMeoIL5qMoyeacnWqOy57wk
UpRubTQpRVPK/C3ulWu1A7dLqo0zVwr8gI+Ww7qni11OgabpmdhCn9p7I+VyXBCK
q4m9UhD4XxA90LhP8Yi0GrWAztxlAoAWAAUq8R4JgVm0szPW27EAm9Q7h9AhgnKW
ABh/QjFch3yb8trC9cp4GoXBSXTCNg24VPQBFvQc+drx3s4Pt8+/R0TolOSNUalj
25MaNqBLv0g8/1QhnjBYcJBS1qBy9eXAervy1zP0Q2Tl12MZ4hiuf26FsPaHJl8x
qcJ+lFLMVQBP7ut2a+en6gc+zlVcv2lunwiA8ywe0emqhOanmCAfvKcn06SpwVRj
/MT0ZLuWJZ7Lj8jNxZVDZLtcl4FKjvX6/ciTRMJmVysVJO1EfiQfjCXNBcBE3+C7
qREJ6BLR5I6jimNgSUW483AUQqC5zJg5pEfp03qmwWQ3uzCPr9wFZrI8v70x5kSy
RXDaOpLYIoCCDVy4PnlBL5TGPNFMnOd7qB9IifYkvo4GKuX2/N17+kVAe8dDBp7H
6BelASEsIbsoMM9gR97pU9Gk1BvReW8Ufbkw0iOkC2MdwPuj2t8uGDayu7HWIMds
xtTw5k+1FBLTEYBcACQ+TCYrmngeUZBYHIu/+YezXmZXtNwKFxe50R0FtjS0QrVg
f2MEm+1wkGVMc4MYkLA2wuDgAJ6gi85/L+0uGD5a3YBpnEcTYfc9DzCZ13AsTul6
iKRYttV0yCAwSpgfod3Gho7R8xCLR/UVuUztY1HosuJYehtbeDFunrn8nykIj7sA
t5UCRszIUlyMxUF7kiJyoxkisuD1jbJrWKUvHqjLx6TfbzDLRb25Pwo1r3AiepSh
LfF2r427ltiILPx6eiB3IOb4b9Dc8FQZeUwte4sx/FKO4bHJhPDNYMXgynISEQ92
Lhxw0g2ZEXo58hq6pejDFEzDB8cKWOe+zfi3geoDLPqJb/QyVth+CAnLdEsfSCoW
Cll8G/HDwF65ctmY8YtFb/26+aPY6cNzHHPX+OjTuCiEeW7BVm9ptUutMxfBEHug
L9AILlD1VPcD9MCzShHZUjlNej5MnNIKhekFtYE73CI1wNJTAxmyjvJzbZqjoQja
1FnhDlwL7SrUTWABwUfzfvbiSORvlxyI8L+lMnDlALBjsuFF3Be1ffCRgydqv6dE
G771YCujP073DSRpaAob/Zbv0nNPE0AQRTB/GVNrqhhSvJwUHPdMceTT7krludWb
6kenmrlkMfpGuamcU/86VuwOx0GqcIKaod+9k4Mp1xvVXB1F+s0NQxYbxD7JlOBC
IRulFR20CaP2Jz6byvkV/Hs81E2ZjsBcoF3mE49rl9blX2v0eivTeYsYsAmqv7Ip
N+2qVNIm3m90qJ0tai+m5rA7ctt2SFTiLL2OAy6fXxlMDHCjIeBbmHeE9fr/FM+l
dWrS6icb4NKl+KRsUj99P72MIzD4E2oqvns9bqwEL62EhtkFfWjK5fx/Eo4LVbtf
rwSvCrP1QLDVtcDn/XCY9EZxriAOZk8bV517J1qQB4METioeG0JNPEdPAi1KtqiX
iMqTiDHnxXIeHuzMUPxGMnufJTON4/GDsOlZvZRUjAGsNHAklpmq/leRcUsq03nQ
AVInLwWZIftr5avW6g0HjQrnmXoqfH79Oz9u8SoVB2/0WNsoqUTl7xZBVYl1GOkP
8jpcyUvkdHccsQOaIUKFw9ZVrYp6dshendxhRX0m6HMlsA3n9PuAs4AijwouoxLU
SF272moRyTtJhVSIDEGd2NlJQs7jSD6qKmfSFu52w53tcyCw9IOhVSEXMu/qw0Rv
QqabkmK/hHaUmEqZ96oHYkV0NjzJvXzTggSWvtzJS4JX+Ta3NP7AoPQBqEq09gSV
Wm4HYumV1wYmNmEl/kXUJjj4kLWDCny6BDxR2Xnm/floMqFyzsRPWFpJIplHbpLQ
eDeYzYzGSasbyDTGxtzgqeE3I75kZoGMNbRbCjX2D+ctzXjbdwH/7cwB32hBNC0r
M2DNKnKrfg2NS/WYW4IMWmTDeIg5KMDPXZyPBe+bP4l17gtRRBMuSpi4tAMJ6eMQ
95E7iWhEUnMrcAGcuNuxagGC8/RtbC0s0TFubh6HU/cdKIRjOU1pnaGmNz15v/Nb
NUD0KeJYIagqIg28bSqMQoHDyU1qd1wrcXJA3BALB6VcstH9PH7qU3doRMDTOTLG
+SbmsFSK9zBKxQQMEoeqnW6kv4fSPJnczBaIGPy5xOKuVY+N/zdTbPuA5cZMGOkI
DXd/JjFNJkaYgh/6vrzxmNNQF8W6ie1mzeEYKW6jP/Hy7lhuZvK9ffhnnbu8nyO2
1dAWjOz06Pu7rCWuOqFSG/y6kKGv64DemDhEKPGpuVVcj+Rk59lDai3Q213MCJ/t
nxQ9I7Xd9PSuniEixtN5hqW8Y8zIGeETpqeAJCvesD+wrJ/8pEuQOWc/f5O5pdfi
KE5cP/OPdmM46MAa8SoFDJMwM8+QjI/P+VAinYtryo7KzwzM7vXWqDoQZon4uuUe
3aQxgXLczrGlXW+m49eA1q2IJVZzaP1S7103W2FsNZjyEt1U7boffqxe5TnSemC+
tc41lrYQqOx+VjDLq9kETkQf/9D8Xrs0m9uaHDWImtyNEYJcxwW2bBexWZgUCV1G
yiKNCUfJ43JnjBRyRVkl1cWsIcR6tGv/l1atB9IaFJaAqrAhDH51p2cxnjFFjIx4
RelBIYEOCFHDqoUZ5dYmfWLAm2J0aCl1iNtqQ5JWfJQICISycvOhtkHhIMBPNG1H
ReJbQ7Hc8cFIdBRmoZfM7gFdqlZ5JLhs71FUvSFHxJeO0FCZOOYZqVZgJymUEiZq
pvwruFh4KKjkD8Y5wBDH0fz85kfZAkQuu5COCkGcoQdW8LSKVU0PS/ChVZeYDVFv
865nrKBOpj/7JKhPcgCDt6pUdvJO4OqJiD1xJMyQzbchhu0zaD763iHHYmidFkje
EKtvmxFzwwd9q1VLvWM2zhs6Me+ZEpA3ZcL0xj3PEAQACrw8Uu+HiXPpWYOyARHa
7dmUFs4xHlAUNxadkdUNI6iFkIyDDzSHq55iAV93pFslkvE3/+qThZo40EHluniW
eSF1/e4i8ztTQ8CoPY9y1PZtFouvdn/bcKdpZhrNOun7+/yAwkhuw3bYS7VnoNIt
17T2IpomAcmwy3jXuncSu9EyvLcWVDaqzx5aNklWysQJj3DP8vCC6zpidf31x1Yy
R6muyrilR0EArkD+OqTGu0umJX3TQhN5WYseb6+5hTXtmQtjILr+FpZfSUkF/0y4
3+jA4TtEymYaMrqb6/3Yr24U4ZEuwJ5MGoHCDiQB1K+GN11wnsL7mKu4UzTVaQWE
nmtY8/++mwPVQ+a53Qw3vI3h9h5lvxwAg9RzQu+8lxkUxKZvFO6sZsfImOSfG/q8
vUv2Bj/42MOV40z6ffMFF9PcdX6o8ytlYHeS6cx3qPEXJR7gOOCIQhfCqEZIO1/I
wVHfRtebkqdzYz36kj7UHSu/z42kqGCswRYoEyAKByN4/zNjqAlMMW8ovlWv9K+u
2bF54w6SB4wjve1sXExyi+1zNSJIyR1UQiGYQXQi0YMYVDElYaRTSNWRbGwLgsh4
qh97QQIkipsMMycLsPfcd0k9H47Elj0r9RkesfFkPLRylKu8fHjtuXFMooz2rFKX
T2U0uw06G9c4R+XCXl5BgEhV+jMofSPNjIGUUJ+3gR8aMq0ltPykLBSWZRe8B207
uVNpIeoHalYIndh8e/mEBAd7lPlUU9Sby01Z2oxUoiEkC7sECwO1u+7OTC/e7+9N
mS+K3zxgjJQ8mRbyaHtC0ChxwXriBu1A8qDAyQziHFS8fi/CWhKA+EKFjyxS87v0
qC7w02eyCRUNW4OJQLk9ySNpFJsEFDhspBOHhDyvJWIAUUqc/YUWLSj62+roRN4L
Gi7J6OAHA0ODUkjwC+jecDyWprp8mh66LuBL5nXfz8sQr7ZlHgc1Isoyqhe8m7WH
0H8AXcFHhGeeHKiPXUf6XAnxqtUc3IWc7ve7UPEKNF9RPzjSAli5biyvqHPnIHPm
XxoG/CzVWrMgrvqJtS8b0ZkyW/Mby4L77mzxLBOYoq9UzY18IOA0MWLPQYGG8DtL
A1LsHWxF1f62H+qofvOh8tBt729k2J5289KDzpEGK/X+2XhsGCzY8IzLpxZ7OlZT
s3Xqzcy0ufpfOStIGDz3QFp47GBWwpnqR5HLUJ5YYOwbesSKOlJm4A3s3rz2Rcct
uBvU8pWkpRsj4DhKkxp68MHVlcD+vNDUB/Zt6te2p/Ft9iZqHR7p0+qS19N1p6pK
wxcaCMSTo57ULGHU0O33D5WdogLu7nFGMRgOKJ/Ukr7RYbZ+cNVi1aIrkk3L3xrC
il9ndcHHTPuAxkAhgz4abhGTv4ZZwq3NmTAYjlAxc2aKgHuk2dzTC44J2Mt1kYL4
n5rtH4++/xBkcBwn23M1a6EF86Dj0NDEBkselH6AytMzkGq1PXC/XVczIAxl0YSl
LWriDkFePHz2oJbDtQs28tW1YuFQ4516UwD1f7P8NrBQsCQ1MKGojkr/XhWu6DLR
HVu8FletotZ/ho5obqfwPh/mb6nPzM0wROZSr9dLExEDjYlIIoh6ZJUPrKr7WYM6
fTSZU4oX9NQffv7DUHSyPf4bjjuP4dTK+Cai82WeyrvPtZdaJNDdbVAHpNUkWYn7
lnqrMtV86IPt402TtLYNdxfvefaXZdoa2ftzCZXnwNn9piiIRrsIzahnTP3zuE3I
Q59yNq5vYInPD/jK3zv7PfAwDRy9WFC93PavP0UJfOjHz4qMLerpbwl5lpRFNoJH
N/sqao27MVwaAPjrNbCWo6L/rxIZDr3G0mrsbO0EFW4GAAHUoWP/SukPTaZ6GEJn
ECcOWotZw/SkL8hBET7gmJuhAx45gZxze/u5C4HeWXE+pX76jiKgoAUJlSZ+90c6
3xpGMxw9+p3EzH0oIBS8vjrPfdTJZmUk5tx5d6kQYUAnYzHhd0g0YKr0f9iZgO1A
bwoHueYXEOy5nDAm1lgqzrtt/UZQs1/71kdXlAxmqrSSuM75H0ltuWM8mmAEs4D0
o4l+Y8r2SKtNRXetDVFYStcFIhbU5dIQyKN5ZDoctxpUfzwOsDXcqzi3FzknawP2
fNcrVDF686VuVxTMgE/GMlAuxDwsaZOyeRIz8Atlu4OQgn2+0Yx9xloHNKtBF9ok
xpmsqzp8YuX1MPVuacXns7FnQV2660g16nGFb9XmUOo1zthwHYnvsWM8ZXNOXfDX
ZrHqoKX8Qb5h5covuwXa2ce0Lk9jXTstKWUZDTKmBH8+nw4jyu10rcKmzyEzDkoy
eylXfm8mr9AMim9Fj2fE159x7G0VobPaFS2FBE/hvZQY0dmZVnPwfQfbx7DsOITm
jqlycX81Zbvgw8yPsl+gMWqIquCtFASffATB/BvYYwslyshE0pCH7LmJSS5FuwQr
GpJFjtGYgy0kj+m9pdT7rFjtgzBlsfpTzaaVV8j4Rag1GsLdZxvWDu1+xWaPfQou
juNV7r44LGSNakjeC1D28UoVO8x6Qu3W2aPnbnSQTaXXVK+2+KPi8+RS9VREVplX
JiRlhjGe5RIPkyt1w7GlMCBGudya/GtsRC08KXS0bHceBmQLpPn8mRIKtx8X+WUN
VIllMsP8708KbgJqdDOThJRGhB9nEHXy73qake9dEG5NHJDkejGQH394WDBFfO7G
ZWhTU103qnrtUIzzBXa1BvPhiilQWNKMH6tRI1FVNN2UOcLmOB5m/BTKcLN2yjoP
w2mGaZb1+4sotjJRayzqusIyaUn3dEKp2W9/9xIChbLY8nciZoyoUNfI7eE0dG3N
7KhIoLjyBNKqV8TnazaYbsmeF9JntpmJ3BxBJyu3M2hwzSfJ2Qr7qZhoIUZQOQna
qY41LyVrQx39TpnnUFQxcYCp4KmoIF/iTcip2cZu4+9A/EA+fSYQBwpGU01j4DVH
XAlQy4IkuDj6fkKjCH+jYhNkTitbH+/5giUg0TaYjoBkcPuO3DCBU3lnrGJsg46h
PwcF+ry1GzJPFiTLsX/AYKZAUFD5c08rqpUnNWeUY2jyjwutA5qYCxe9m6U5rA4S
B8L8DKKNkU8VJpj6RGi3OIiTojt7361CGl5GSB1rS1+P3UE6ovlH518bEFFhmBUG
nlVtSfwmnyUcyoQ4oeNMY0akyL6AbfbyfqMTK7+tE42uoAJ1Zswf/2S5y9QsXZS/
Hdlc/KtOWDLMaNje/jJb9yo+n86jSqQVSrThLxz5hcVqwxrk4O6gMbEHhyyPP5QB
X1d32wv/AKGq5KFQPxArgy4pSjdMrbxlXF6jicwerPMs7S8/corlWH0dpsULlnDT
zUTUSWP96LRcnPmhvXSGrxiH6BNEofkOWFoE5rk+fZMzh4dGxCijsa2e57Ira3Ee
QLS/7ScJFU1f5WpGg6p9q8xxf0dEQkAYIIhYZNcXygagIYlAeKACO5Ih6C3OH2X9
UqTO65u2XgpK8SBf9RUdyyPUEbOqR4+EbOw3Y/MMWVO5GxUnVv0Nt2KhiBxslNNe
H4yMNRwBAtFNHybIkzElYEvwygiJytbdCB0ErM7WCr1h5aIXMO+FQaE1Izjg21Jw
a+8Yyh1ec2rcmxD6HJleY7mYnFoJt+5OBPxJD84IXLiS3QA/jOexCwdFcldHmr6a
pW33yFko5HgxfBPv8UUECK/HAIKAlFUA6J5f6pd4AU8miLgcaY0d4noDdUXywPYR
hiFSvva8l2frHNlowRzCiv7tHDXeyZse9amQe5llEU8VuJy7StJOUTXXiwuj3k0o
XrNSATcJwOTXUVncF/LABHkq/ERxQKUoweWNLbm+An6ocFsA5CSyWkqV4udi3x8y
lEPCU8c+OHFwW9gJjD98DjHGATOVenaiDZOPZUghCo66j5WS6XjbRMCYZ+UZYtE6
NqEgGBc5aGJjv2sqaiqzkUoN4uXOhS3rzXcC/0FVwBnbOkCC1EDugy34mlZjh+jj
r031Oq0oxkKyBbFo9FN9HWjwYhrY5Tg9r3hDkkwmp6dKTQaC2GTKp3fJ3XHj2mJM
XftmLGgZ0kCnM/9YLzyAaajMXw5j4YmHXvg/rTVqxKJDPwssrPRS4KPam8yD7CTK
Saa+F2Rso+A/htZ6RHasd3yUyEjlKukXLsY4U+Sg9ENqFOJ1WY97hZATX+aLYxKX
qJEU7vGfeojKVQmZcCUZ/kg0cSRTpnG6//W3l2iE598GCHFF1tuk/yaGH0Qt8UGY
Bfu2yxBxugDjDAri9uMc7PrPM9iZl/ehsa+cDQ+qTpl9M9xtwo6YsOTmKuB8bgzN
DW6PvnZJTYZroT32dV+HlclI9VthtqBSNSyEvFg7894CcCetYMNY10cvzQGVzruc
nJOgWizxnmgvRELSdecM2NZHCraPdJSj2f/CanNDiHYz5+apYIb+vWKT/qqXy2s3
E5Mi1o0xijatD8Y8B3/c9vlJzFTOD9LlslPXl8jWcnXVAUwf3MJf9XwzCc4m423k
EYCfvNOWT9PXJgqWsIxnTZB+MB0aoU1lU5CgdzdY+sVjSCTtqJ9bsQdF7GD/66kJ
d/M8AOfOr2y/R5wPL55dNEoGZ1uE896m901BIlKI55gTG6SQAVPaKzIJNvsMFizz
/vnrlpGmqRqh88R1BtFnqIHelEyrFWzXR+ZeBk+MceFURhEh08NBnUrOMNWwJ5Y/
+kRDRvWWSxPAdO/XTxa55n3bL+bWqEvddOJE4TofA4Mq0Y6kqmD9VXf0AdfKC6jt
Zb7hT3lCuKx2BPpRvCDv5yx+NimdowbMjKfPabxGCYYTrV7vQG1lzKCsr0g56jBe
gvlzv3j0PDZglSZvNRuRd1jjSYfcHoljMjNAYxgEC9stviGnlJv/gwVOcjsGENnw
J+oBwBh+jEaCYL5t55YA0QmxTSEeA8JruDsi450tWwRRSSiSTVp6Q6e+Y39+Py6N
geJZRqXrVJhdSktFZSRQcMerhxc/vXL694yyL8HzCgkXdjo2nLQhq5p36FQ3tswl
Lv4AYzmL95T1XdkrtkTJLZmYkNotFIodXJO7dMO7OKYR2mSjHOsRManwmOn9AXPC
CvugqpX2GS1POQ1rkyQLNYWf6kJvpW+K9OwX3yNB4UEJKxv52vPPF2+KSdoq343l
pTmmmPz1l19vmRV9wQRWtcpU8hHxvTBAi1x0HKIRYsGJCW/EQ+Z7LjeGoQ14cpkE
mjtAv55lKvOHSbhZXx0e+ci/Sn9ITpSWbhFnMzV0Knx3F9jP1PgFkNtXnm1mItQP
sgTBm3QixVd0nIyBxODtkstzsHz02O2cNqYO4k8ZveE1Y4KyHekVrldK6w/G/WoN
cPUVeZOMz94HtEhdixDfhCZ+CGLGIIG+4QnHPhpPxqd3lGGTr8+xpDC/COOOQ8GH
UJ7NMGG9C7zKYEBwKmFPbGdxtpIacVVbGOHiMRZbOaogFtFxTTncQ1QW3MXaoO7j
dWElvLAuUNZFi1/bGDHULKuVrwr50tkTs/a1HMlU3FLGb1SqIRGWIq676Bq0fSgB
Bd/k+wsy1lmNRSkOVmBu2oyhqbVWYrEA+tt6w4QjwrCypYuXS8Kn16wveokVhk4D
ub8PxeFGlEBXPuxiKJtC0GMBwdPSZHOei43w+9Odb4smBzSYZeeBu0uYo97xm0kz
T1evC5NZV8H6TbYWoIyliXs3NtgVdfl3C2wz2LfFzrmIRu/4+XViOFFrYgc+6TuO
ify9Uh7RhnFNtrLMsxuueQ4krOAUa9yq7gronljgW8AHNwuOBaExcD3vQ/58Bj9J
k/Yq0TwGUVhLFFgO1XoNqbGPBI2egnHZ0SlD2gokN9UZg4LAQFX7xrosf8V1HKEU
Psdb8xWBIi9a2l049fTqTZcAyeAc8SJUUga+A+YsSoz9LwtesCGX8DKYzFe41ap+
7wqcxbwopETrS6DMZHW06k7og9HdkOGydvQj7dxabSjrNYPC/yoPepVcTPbO1uru
34LDFF87olRVSgj/JgeD0FsMeuxmjFEwpEqoVyE6gmwvI2EF8RrKJPsydwEshTuG
izmlz34Ymu6gPOfoEsoTooLOiwOKWAXsBQJ7hhy/o7jc9kw8GR11Ye1RL9/nh9n2
zJprkEe40YycSlIBJvILCcHb5pTGFw9Z0ECI5S9oWcnPe8M5UoEQJ/h/3MJaXBxd
TBeWvDjDJC9s8z0j+hl+hnoPqLZnuA2gKWWQb+vVcqgcwSOPDzhJjPVGAmgWdsbM
eUhQeBImG8cr+QfCB0g7no/X1XLFs+sdLBOqCTzPJpszvKe7cA1tj9E6Zp4BGEzt
+zrUa6+6+pJLKa5ADNsa3Za0dO/CeRPbZ7mOmbNpqhLyk58bNr5mx6GZN0Ljd7H1
Bcfhor1UT3lCbG+FucXNrUbXYR7hOuS+vx9jo4VPJY/wOrzpE/m6+fJY3PCYOqhb
0WwubxjLIilMUY5f2G0tMG3+esbr486+bm1Ly4h2NvxTPTom9cEutQWHWEQ1zMgz
wgUslp3/40IaihpvfXWPtT6gJW6DQ/YB/zFMNa57IqseBJepvyBk3OH+CU6EJlZw
WV9TBeDFwZMg93JQ0qy3fK07kpnSYK00DaKJMQEsFkBoDc4cozW8f22fQVnc6jSg
4GkM+5D7jfKEYVglj2/CaL8FqyWn1F1qTOhTM1lGs1TuENaaFKvpyXfjX5IY1Kln
lIOk+5vazYEA9QCIdxKXrD+t+6VnTonwzFOqYRKAKUIh091QYQ9Wf6mwXlrGzZa1
s2UpiQDb5SjknTMZ9FO4VT95Qp0NvRjVjpoAGhQa2xeuDY5A/jtcw6L09GIcYtdg
nE15X30lzD6N393N+eG9GNtv+bUFC9Fd89NIIrwIy7NJ78etpkm0f967Wa2sUzVX
uZlok4UssNs+z45IjVjzggaRzc20JvBJa4sYkjP3v9KQh3fRTL1se9VIHsRkbDks
fudtScVX1nAJb4mrig0xK55EX5MtAydT2oEpYui1B1bAHi0M8gOmRAkuyLLucoVE
hRcPnrwALpKuiMarxhqn9oZlO/1f6cjf0hJZkFK7Dpc/A269mh+HewJUs54G0JIG
BkR3WJ0YDxafzAlyCQsV76PeYKGjwKnYUw7hYdHi9qhPldHjP12Tx30phTWT3oRW
HXnTXgJt/4wWYktl68+o4OO2XeKZ5gAGU7QNpwjyiy6m+89Z360y4fgMhbXb5enD
mXKxBY97xZR3xbgODm6j0a0+oiJwRWo9gSuIXJBRqANM/oBoZ9wRWu/bxrqnhG3O
SE3nvsEZSubBrQF5IM2SLbi00oqogZYrLlAvXfLBbv57BYVtZqqAgtUXZcQqffU/
EYtPp4/YlV7GQWg1f3U8xTFTFYKyT1NEKm6zMi2QT2WP5DBTtprNOdAjFWg3Gvdv
llydRzZPstCRhDFCTSRgH9xkmywbqRxAobEco9hy+G3Lji9zSqeXL73iREMlNoK9
reihSGJwYFFgLXM0Gy7W+oxL1ly2u6qTav8OtuYOA0uLx5wIm65J/Vb2wZrrkoaE
g0K6lyqZ3WYjGBkbdsjF3jK5qJag8Y4WrcvQEiC27dcQvlj9/eLYDMyzlhlZDEMo
jR8rQuveL35Ddf1g8jpSaHPWMpChbEDrX4KA5rE96u7UJt40K/t+oaJaXoZSWYLm
rj9XoVxXPxuycxeROldgQHAKCxFlD3PjP6CeR3v+U8GDTnFID1fkPDITTnZu/c+y
bpAJtYoSFtwYCwYki22WikLhe09MpIWHIwuWGQp8OW63W+Bv0oTpNg4Ay4lvSe0G
gS86XOHA0iFlA6Vo3ZfuurMy7MKgC3f6xWovhVumFUj6dzYbh9y/+W7RB0tmSHTX
PuqyuAk8WSHMtDuHc+IAC+XqbRH1CQvr+pqQEt//pE4fkn0LwKHQ+LBTPBzOFn/B
yw9BoU7DBQGIsrOQehDK/2iLix85Jv+P58Po1X/DwYuaIhkdn+BKiI/JDsNM87cc
rRoFKT9kINEYRAscj2Xhy73T1oNalaSdAXbDvKqcLTj9TgfsBRZQatQgx8J6esq1
6R4322N7BToyN/YPDTndfQNRGdHpPhAd+5W2YY0zcskD/LAp3NOL/CJMuQ4L0gMD
hHZRjF8OFgntczcYqyN1AHgyJM6VqQsTPhbRagSRhZXy2nbBSiAovUamdo6+lPIj
XU2c0MAncM/mRWgiBZLkErCMFiTNLOl2lgl4tCTtcqJ2pvsooSBk6r51XJG9G/TA
GtA71qTF4yr7r4Yr/SkujOX+1ThZJoonbP/by8ziQq/x+7hzH/FPCxf6CR8+06+M
WCy1wxj19UfAe+nPSe6KrD3ZTP7lNDMGJ0A+McBEBluZSA3Gp68Zp9WCQ4JJLxjD
V3OKKhXh4S+iIHdfxDsTw4PP0XhSGz21EhkT2/1jf3YQgdoV/KmFioPUuVIgfJ4r
tu3UN/Yiyd3p21M/wAjLMU/heMNdxGb5bMMvF6CRQa30STRKCFZ8vcWxWcfHgqJK
fHoZmMKV5WHKdoMzFlgRnbdgOc61R/+uD3xz00MkOeAiXNTYQEEV6ww72NtXJ4Vf
+d4aHn6CLdbpgFyCpYMOkGEguLvrm9V+R8xrPXIhT3NEhEIm8KmqGv4vxYdwkoB6
LrNaA5cf3ApL150V1+m+cEw6pluRmoPYD5j3Mrs0RgkvJh0ofhEgBE+5Nr6/27ZF
VZNGWBfB2UNGtj0k2V7H2oMdqCgIAJ8prBQNQd2Z/xeJ/q30lqE+pwN4ZMVF2BBb
242REw81nE1kfmHdO1f9yw0HvtQZ0pYKmr0FVTi+91MfST9UK3ooCujTj6Alz+xf
7fa+1jQVur3I0kuhIiRQ7XgGs/wBiK1hHACxjYP7RuTsvYKvOGnixZpDpViL+clU
uDIH3XVgccawdSUIiayvu3xmyvBkdLPLGTJvJpabDYRl+8KdsMKnGkzo8tPM8THO
js1Yuqv/saJ46k1KhqLF9KG6VBOvhkAa/LIiKTebuFB63ejbSUFxoHAuj5wLCizm
RPfqEkR/d3uiHuxIBUSNV/pXX+YlCTcwr15iK0TuoeV5f7v/Od7ITyqUYYl4Su4d
+f6SM545h6TB67DHzxDSsjCgKGsY3gJa8T9yQeQg2Q6DCUBYoi2stYbkhbDxsiVR
h9Fn339hoOIhjwQlJY6opIIM0g3lj8n7z7QZqMIiJ9XL3fl2bVAP2rraZrvsYPR9
o1tJkXmm+X3cTYN0zKabHxhjl0zrWWzEB63q8m7/Yu0btDt/ShfFg8POfPEH/rp8
XngnrlbV/GC3fPBQyCcS2z+F2CIaxgShSKfMsh1X/z2ICwPmLym5ZPiCczZR9nsA
DPxxWkSiyrt2jeos168WTRV+LgCoOd7CgNAehjXPmsI1KJo8m0tj/W2NtnNSxtZi
TkeNSRyF0z9EDr0b6zVrxKlROQJKLePKxRaPI+8baZiFVJP5lGRCQmkR0AWHcbBT
9yjBDUBIRu5BdDACT+QBnun7cXTOI58RK8fLpE4w4rYvi1Lg1k+1HHCLAu0E8w5E
SZLDxLMTkAgKSdpgDOsnAHdgbrvrsWi0bb2GMX/eJu5/u47zwQu/gWJPep2OTrBF
0q2GrXJVZ0mZAYqnOitxm2l9/71dtYD5IsYB8tKnQ7Upp1vdeJVueAHpoBop9A7x
NSre9T0QbszMCINoNX5q+9d1WCROs89bnYkbCfQGHeJCdfnwQV9gsch2wDcmER4C
O2oRw9q1SWHQe5CH0uo7Q5vbp0Q9J0Twth3/2pJd5m832ARJhvaD8/FNrYhgyDM2
7WIYrivkxZ8aCkKOeEDDS1diCs7UM9blwJomYwh60oPE8nC1ZcVJnAdt+YCNo/wI
ogdDviTYcUrZU9Sns5qBKdMDE0NPrqFQ7yzrppZJUlzxhW/duYk7HXYLehTe6PV+
24pJhAWJK3z+l7dGIfqOIxlAKGRFhvsmA/uUqrom/MRwaz4SvxuLHsW0EGstubbe
PNOQaLvsZwtbYf1X2IsazllXecib0ayqpUoVL9l3NlnjKy7ZSl/xG6OaGCwBlR4F
0qfsaMO1yawvka2Pog8Pmb+84iSlyjsPa5c1f+LZ39fyBVDfe7nFxJtTyhrULzZw
SV78gCt+DeLVqkgG1LkS3qf9qbxCJDRfRzUBaXRyGWR82LibBxK17zcCEVWck2h7
pwJ3g9FgcFVlp1ZVfPpI+IWUOmlwrzv2XowV/aw5bk3fEul8hmkGvSVSyp3Qa6li
he97H+Z+ghNCJ+l9xgX4ZuUzEif03CH6p0BcMj3dpNCQb7V03rxl3xauRMvNjTSU
TjCF+1HpvsLof9atjxCtxMF4vWT4Po3Gq7mFS0AKzjXMm21rtsrRp9miNunNJCJA
N+/Dbo7Ipbz1kRyKLq5732mZhvqwuH6KFMznKbz/k46RRhKR2PhBBSR0BaAC2Axw
axSaRwXLc35Awc3un3BULpIg7s3C6G/G1xBEcqJ1dBBt0X4nL6z/7CMT7Bq0VQQ2
UV84GCEkv/AFRjRPGzY4VxqLopT/DFK4+OG5QBg7uksbrTDGwaMOBJslKNDlh0Yd
rYXz3AA0HJH2RELP7V2VL8Cf67Rkfw6ej5ySnBER00AiK9+HSyh7dShYZ5o2fmKQ
RGn87GKWJ48vqj17X8ph2a2crOiaHYNzLxfkyZRenVMY1vwc3hZKa75m9gKctmqg
FeMZSZK50j2p4eFZPoeK+cjSNFf8O0Dhs0Nc84SUvBWA10mZj2VTBgje4CEbSBxN
nTjmwT21N5UDlKTdAeDUxRLmG4dHsEcJ63hXqiG42pgiP5O4gDLPqBqBvLUxRk44
Nk6lbw2+4GMC5ep25igfrjHQcCKlI3LfgBsfLXHIyFWC7bgCrBAXhs58P1EQoe2l
YMQAC3Lobdc6fOZ7eZpVFXGO0ZagmQD4PvxUGgTVVLFNLJJSf5H+l7Ad52Hnxesm
Hc/ZLz41GfeRmDSPzcOw0GbLB4PFDOpH84BvnoiJxqnv/i+Sm0WUF1LOkkCygnWE
y7RLr9GSQEWov2dLrS0tzqZZ8w2I1erlKiA8ACUFemTSp4KrtVA6cEGl2miBDg3P
Jj7gsdKYasKnDqrLddf9goAgVzVGrNnJCsYcYlna9Q456rK5oVHT4WJufXGL31i1
YHIpJr85yaI7Eyj9E76uuVidh9TfMRoQZh8Z0+T597qpfIM0zA7JtMcg3tnwPWrE
QCWSpgtuD7VRjVuBF1Kki/Q/z0pNd7g652QamjXMFQMlUm+gTwnnUVkdaOEuowus
EZjo4rkMl3m6x7RZIUZQr4vWDkUFBLqBtPz8vtHTxRjzJIo5wYMPJmGdKbSN/j10
VPFXCs7JJHlnUzoRhrYl1I9corjSnHRdUnirjh07sHj4+2d5g8BUW9Oyl46SgVbu
ZNA3rp9Y41IJ78jaXjzQlUnlHPwLNy6x+AZlEfsaM2i56cPaVoCSj1AEJU83Duxp
4hg7pZIHsDsrXv8zh9Bk2fURNQKoTnvx671+ZInqlUGPBM2DUteA0ySXBPnT3iDS
RhnxcJVJfXP/o0BLkgU4yOjDRZFhzd/7DGakiynZE7oujUgOKabhYb9yut9hxWBS
9UmrPTwn3cS/9CRPBOp81Yrvve/tUhsKEcio26KA+eJrGNGZAZHN7dnZk+Zzb9Oq
rAalPptki6vSSLq0MEos/ZGSC/f147fRt5k36E/RSCDjFuVa1q2On4B1H8qadDiq
VjftJenFPZdmAjd+M3pfS0JEhjFCIa2oH1HmPi4OcgSy8OLIyr0FiGqlXePpeYZA
SttQUNoWTIe+62+6jrCikfJx4uHIk7YqnwdqAkdOQKHXQg8SWlb2hJEWk7fP3SZR
JT23ep6KzSiFAjow1nbsGshADeZyNc83MQwDTp6MlSmypovMawEf5sFbQ4wBBx0/
tciD873cT91W9dz5PRIBT8rWvH5laSfTlpx8vuYKbgeq6S9+hx4NAiL35B565JnJ
fpN5ztSOl9OT28/4WIS2qnLzvzn3vmJE6wzyVpjOS3GEPx7COaoHPSJ/axzNXCCl
eyaFGcTp8Nbe3oaQKgdepg17ECo7uI/lDLtM5llQdRc/0BNeT+7MDH4Bzl9fEkba
9YWhQLM1OGUyf2Wut4c+rWq6DbT+PHbEMRZdXJUAzFtKowu6N6+Dw3aokQFPuJPK
pJ0siP8WzhPd6HycZcIGkHjCpzGa+Wap2EyaxSmvxCjB7it2n2MqRTzTsdRsLR9l
/PVyGlaXPD1vZrGE5j4zqvQb4vRd10ZAXZt9s1RTS5k7Is8ehuAvzkUPuEL22PHh
6IZa7dQyi9rsHQqhYLV8FhX2AW0sSHRMvn3ebSCgUPHz3qJ/bUK76GErDaWvLHAy
Prl5+Bm+Ln2JwhvkuU3ucLJRdFlBQfPJ3vxu0La3t939Nab4Js+qsagZpIKFkKAm
2YIL4udC57WNdnfdevWbIx4ym8XLmJqJ9kyHBs6zx9NBC8ZMroZgtCDSlZbWVK8+
VK6/KgLc8XpCnW0PgB+b/2kkqoe3+3psL2cQ7LEOdk2sCttLvIqPlmeHjHoka91q
MkvSpMtTHeG/TGxpMK9JcwPyGdbg5gXsTJG4gabDDZRrQnxInHvqAL8U8gzwk5Io
kv8FwQrBytnZ9Ebg0uuzHFIVnAYXRVqIYlW/B6GHLv7zxvdwTj8hjCCCEsCeN2z3
tKw5ALZf8xWNJLLRPXyFZgvVQ9geACS3s6sTbsH5h02HM4Ay7DcuXXikBzUmZTmR
3QQCF4dpHfWRC+EsnxXFGLJ8ImCF/aTACOuFUzUIYahAwjwXaNPZRfS+Ln74e8nE
HlBBdF4Savse1hy1ALrgZ8qA+gR7mc5BfNWpfY3u8gsOrG85+ilf7qBqeP4laEVD
Q7uqKFFbacc10MJ3Yi28PDSqbsHECdwQuYWc96kaUoGJup4AiQTRXHtAiExH0REV
9EsJ/46pNq/lTwhjAShZU52/kYoh83VyMHmzPdpzCfFLIlF2zsb3lnFWvICAdXqM
ZkrqjgJQx9iZyjjSh/qWm6YbaFgp9fDbSqy76TMtsnDaHmzrW3aHzS3Z7fM/hEZA
V+qby9UQLOkPWvTYaz5n9gNRE60zj2O3xdwfeMGn0+XuYwTWA3GY6EZUJnQGAWJJ
GBj1UlBWo+JK25J/s4/hstPyd4BAFaMJIC8f9i43gUM5RGsclEEWzjt7zOMcu3cJ
zudGnViV7dKRit8AmEyJwgDE9EiHdG5O+AB2OM2Cp0ntyiezMydpcH4hEgYiK+2b
YNdtaqI+lScGm97GgutusBhlq2WyKjM21LBd2E65XPxSLJQg0AfCo2JrwA0mTPp4
FNG5zQXJiTYkev50mtmIIzh8L8L2/Svi6vH5ABoXj5gJzfWErJfG3/fjXDmzaS6C
18/yc/lz9VdsKAA55Wf62LAJAkrVCj5vChgpgCsYJURPaHxw8370y3CgoGGX1djf
iP36bEeeIH7KBvmAiQP78bncCfgX25pexcZQL4d2OPfLnhqvB9l4pBg7IH15SdFM
z8+AzI2ZslbJdi68oDLkBrpYD64cl8Fj98S39WIJ6pgI/t4VqXznAhjCj25DM3Ty
h2cEb6H0RYRJ1bu7dBidM5gch+ujdVNMN5FA8dkQAIB5DpLog6xAIVxrrr1B72VI
8OT3uOrULrkwgp5rEHZm9XxmCay60RSbxO1iS/R849A=
`protect END_PROTECTED
