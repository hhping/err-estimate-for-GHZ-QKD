`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RjGtTV5RpA704OQ/lcu8QE0sgSDJDW9AH8hCjpDraFOsqHkt3DVgh+n5dnL4fijS
zJegkQm1adfC/nnhKyUs7z1gZypHPWalo8/xOOtH7KbccT2kH5VEbjEaPJp5Yj7P
NSu5Zf4cozLfKErFxIh2deVUyMFnIXqsl9P67C1omEiLA6fZ26z7DtRv01tM09yN
MZtMKU5NmIIf78vnItzjPb8skjn3y7frZoamlHJ/VNp44vD4eGsVDp5T28PvUVS7
4y80Sf/Zd23HsUAzFeZrFK39b8O/+WfAgZWkIXVG+4Hss8iHhb6JDU920kX1NCj6
+wR0u5UgY1wLwMibl1kwSYJ9VgTRGuDnH5oWCertbKUjYCKFUOpfqAQXCK9pTrgm
GjfgkKd26OpxR5Cn0RDfzBRk1Vvu363cznpcFT+c0SGNyx3FdM2eMIiYTBkVrGKN
dzQZaGW4Lc6GTKK6OK148CBOAxmhIa2RHLqQ3z3QJmGAOPrd9BQWp2A4jkGgoJdU
KPRqLk4YQ0xD13Q/6DdKBW5ag+VmuvEJF/DnfcvZ7iDkzOBkFoCKS+LldlE4zukE
R2BFuOkGEFw9aeZCgTbXp475Ofo3rqJi+YWlxdI1fYwa6oEBLNvN0q497lgFPmGg
iVQPVFQ736exW25MhewoYNPRGdNvCWESeQKRHt5GMUtvFf1Zu4y/fKR4DzxSl+CO
qkQUT6RKrHcjhfwDcsrO4apJTrk0i6dHZFxIfdmtYCpkPBAQUPzLSs3+4FKjxs1K
Bqvwk8KUpk0XdRGd/9L2taY/JW2zDXvC/ZZbib48FARHhy+QMaYionfajrgIPwQj
yIIz5ygeQF2+V4a990vgLCjbTaFoXgSOixObqHskuj9/A8bpW/mtJjnIyMsG5x+7
ssg/gTlDQp8m74xal4+d0AMfQPJvsBy9mv/Ab9G1Rc0284HRtLU6PRHujxNDCnXA
3UU/YfDSeivezmqhVoimd3n/WJTqJYNq0cMTktKH2360radY9RI63SgkpCQ2lEMa
LiyoDJ2hUAWnocg9ftimos0sOWUgJ/ccWSrpf9lac1QLcnlGrzhw/CyTEfXqfrOO
X7mJNMkWJNW8uPIF3EnYrpuKFoPOfVCuNiFrrztxRxsu8JlQVl39AzmqucEkV8l6
57I832hryeihhmd58WyPJ4aWmyJW0SsGRAD3TV5vLnPeaY9vg7x8X20RfrC0mJmw
AjzoD87tNjvPwy2ybaUBgn9x8Fsj7tuo5lpqOjpKT5m+ViYnTGLpmmS/wwTzz42M
nC74BGzOD3wNMBzWtdhsL471hh9SZOpYHXqYsUTVM7xgf8OlzOeZRofQuq1SscLU
ZyesHMYST6l0ETAawJux2xWW1DRYups5bWecLj2AZRysI0Y5cll9vUqHZjCuMCIm
a9AopYEPdYItCBR/HDJhuIYcHdLd5z/HEFwtr7LnO3vBQTfrRgezuvUodlWnpKs9
M4IS0hsc9D6Cc8RWHRNF2AmXOMLBVjuT/2KZnblZeiquz8firhr/rXlDOAjUoGS/
upEYhf6OoGFEQV5T5eup3Sx993X4bCx7IX1OAlh0sozb0d918nQuE8j7s16gsfAg
9k5BEib/78jXys/7bCNViyQ4yM5XhKvUfvE9tJgORl/7ZQI98sE9eSxXGft24tIn
7C7FlgnZXGB57rgO3wHksKNIW+bzOZFJG4AR2V0OiqKZ0Fijy/cfHMOy7XWbH4st
Qw0yDdOaGY6KcvyXJP9nuJZ2xZkrHR6DsEq5myTzar2CHMHUjyvj6Z9+8qZkWeXB
gzqHZZhYvB/flPQjAUKKA31ed9S5AXp6lkCWHFKlelM0skVJgB/lHnCZeev+cwPS
FxpPOcI885mXjOVC+Zadee7YByC1z2xyskm3NDk25BgX708j2RO+bt9pEJmN7mcc
nHz1atNynl0ogaZBmGpyd207leEcA67gBJqjFklK9pTwdjGzdtyu2VUQYepTJ6yf
Xo7IGKD4ijUo1Gp2kPxoaqeJ+jeEGjTyqpZ/SPB3yQZPaNslMD6NSz6Mi+/KWIp/
M9kwErZQaoQr78P4fbwJgL+YfUwDFILmsOOqYra0s65MJgwZ/wpr4AXELoVRY5Sa
Azqt+Uni77/thmieHkBi+MVg61lzWUZU488PqdNmIw5Nqa2lppQmiMh1bEijxHTs
W/IXzLRTX5nPMctSUdopWbqr3YfzatEsJcQTE9sDc/DG12wE3zzlQMl3vlU0aiF7
`protect END_PROTECTED
