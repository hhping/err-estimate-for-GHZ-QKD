`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hEVK1uvzE0AMpJ6fHPwaMxiH32FCb+2DnoIx/doAxgBT2zQz6HMIgAYMwmB6EObi
F8rKk6UVLguC++zTaVTEfgnvhfiv6BT+VHWXdXBlCYApgkEPu/1qWJbHfdkPXk2h
3l/gX+f2QcV4cQmDLtLD0SW1jWGmz9+OuSD1FhYUsQl1BLiuMu1YXe/73ZBWacvB
Oechm0qjd4wKga4Tes2oc4UZo7/5tGN9IZtjwrnDihGj8GuYbnCy8JCiIcj2mtyO
/yvPZRA9t43ExULAye+Uut6rHsGB811SQOyVaPzybpZDIrolBxU7UN911ZtxU8DI
m4ejcr9FRFIDwbJ2z83eTZ4k+3otIS91L2be1T8cTqu1jCbKlEfyH7fuyulvxenw
ORIRKlS5k7H16+R5LaEMLAq+hwkSCC6rof4UC5TEpdLkzq8cqtkKC3GoeFvjTZXh
TG4i+W50k8OLqf10YNm12feR9ACBDJ/ijZcwUKCnHAITr0S4ggZUh8QiI17huFOW
I+EuU+q7N14PZ3HA5qSVsXD1JRfn8uUOHbxhJoisEyk8ufrl/zb3xO7xDo6H1J74
CVkSb0mG5DTA7n10ljpMa8lER4T9h0zQsUil6hyzPXJRQH+p7ap5IDqg/y8PUEcn
nFaPyQGDQsOikCrc4Nmf5x2sR4BroTkoIheZr2qlQHi3tyNwUpaTdEmWSp2mClmx
1XJfOj6UU4/Mzi1ivDu2qR6E6RhFHsBW7RkAYYbxDWMB+pQDbmYqOFeBGZFCgSss
XVZbbUhsF/N/jAaB+cy98Q==
`protect END_PROTECTED
