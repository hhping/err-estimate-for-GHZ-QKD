`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+bRTgWfuUnWIVaKk6gsPxzi3+u8ONk51xwhWtwa8NI+OhuoshoAdsBs/WOyTWSnB
p3fqoO7EAPEojJezgF2b5Egv/cIAHpf9BawUDOGhcUyIGtEV0wldzVGhDjGYAxtg
ULwiDUOCbaEHqGFlEvAd07Q+HZnsH4kRqQJtHmBfsPqJn7lbwEJ2Bi+9Cg3OyLKk
zMqH0AlHZW5QyMMfHoIcjyp6rWaZULGY6+i7/XU4fqxH9sQZ7tsavd2OsKyO/Rte
1KmuC71mrBADZqqwnhbOpGiqy3XPHpgDw1fw/Sqve0/0+soV05nZQO138bMzyjPv
4U6xF3dr+Lci6ybFL8GcCQN3wlqKbU02h17gv90zKayRkQ9e4HSOwdqihoIBuRY3
PiZu4MP0aA2XLAQ7MchjQm45ZzxwBH8eLx5J+UKKcEtmRG0meZFimdM0zdiLDmoA
ZhEJLlX3Y9F/Dflx6z5qiFzArdkYZq+4fL7o5n15f5/AEzfBMfUyiaXcy66Gsfrt
Vn/2SwzGrgqlY8YNrz6JYY1TqrKWD6XrFtUIx3eXrfkf8WPd2qa66q3TXItvAulg
WBqlcvQy2OzHWexNrLFJmpn77b76ZgytNhWSm6SsLSn7LF+SIlJ75ugbbaHQQitg
+hEXwTULFRFdgvE5RbUDiXI9UHDidHvm7l6i08cvQWOLBbrSCXB9cDUJJoT0scPT
iuRjf6gYwo6HXqY5jWXpoo71bqt0l9KQp+Wos6rb7euRHMO7dLYxfKlGV06uv61S
M2HupkOqdOcYxgUXJdPqntqMlE4vutGg1U/CSxGMZWz0pEpGWvUq0ax7kSryZmuJ
ZKF+Xo5zRqtppPhhIH6Nh6CPJ5TYtYlYXsSRpvYIypTtPBO2KZccjFoh2Hp8aG6k
+otkHgmTAWJSKutol97IPpJJZtaZS++gabIKccEHn9KE7Pie6K5YbI8x1pp5TXGs
3ftk0BWu1DLziJBAoYiX/JVQqRVICMWMFqOLTwsepl0R446NEafkKuQR1KpmMLYJ
tX3XRp7NuVHO2t/DUVrAZduEllGkqfD7kVvlR8GZAiAwhTLQ85HY8U0qjmXuFr3C
l4vN4LiNMVJELsRlv5bCR4srQhjE+eKOFsfFVMV9OZivIEBUfJ25eskaIrOmB3Q9
1sgWk+vnYKnZckidqbB+dpaCxptZ0iB+R88iD9NOXkqsZtiAdlznCZa+J/InqgXj
bHYmmAXQqucdAibJ39I1wcWhVwrWOdH0mkksZ8PMfm7ojG5oooIGoNLsWDrtHxFK
au4L/32sB1r4DCFGPJKBoIrcmANAmuKTFtq4p08vIpkpVpaEPDw6fnwVCQiO93D9
w9Y0EqYQi+Yaa1spUdrJR3PKFz119uA5JQtWQ79Y90BvLxXW+tB9C4E/93jTTbIq
Yl83vVHP6vhuOkzPdQ13D0ubzpWyjaJHx3iMfsuVi3XRIB7mnYrWYHmPyput+C+f
dWCjnp6+u3kyGDlFp0Q/M2iP0ETc6YDCxmtEH/2GXRM1DsK7nOsbCbjPsEYOlif8
0SfFsKQWGJQWNiqLV9afqzvOVUdF4cclJ150MHhEvtoeZyt+xtxcohTr2DYVDII6
X3wUaN5imRslUBDMX/KtiLktjOFnrZgxq2ntd9ZqmHhRtjQaiRkvVN2l147NW3nZ
tRcQRe7Y5t0Ymv9bYVftOdPcIHXZ8Px9VqUHtEiiA9QKAQFz9JfS9fjQzZC9heAk
GWwIPsCByq9XbhaCrTl6Oq4KmTUnV6t3nNiPJGPZ6aK2CjrQMToLJycBb36K6hAn
/M7vkOueE7NEVKBht2/uCEL7DOzAaPx1SycGwRO/M4iIB6R5AUBlzRzTxNRQAubP
l4VT2/SNkcoUOX9mxopAL7lh0yhCTNX+omKEHjtiCEwWNI1lyDZOhOO7xdZ/F9id
0ROcXWit8mBOzGEWorFM31EUlyprnc4AA7s4agDqkFQ=
`protect END_PROTECTED
