`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h2zFoUCodcNa2Qu6AXdgqYeFDUox56KGsgvOCSJ3AyYu6SEWNV8hkmINcMemusp9
96U3GgWeSrRBopeNTxerSBke0rb9yX71Ws6usK1crK0MFfA+S04uZU8EoMveOQyH
rV5XwwnRDlM8t7LCbQzLePFDWukkvemO/t9xsJVvM99UE2qQe+EIP+g5ULgjvx4D
PnFnx82lIvB8GUVCTrovDUUNG17olQGfBnlsvkcjGQNWD0nJqJOTMkRofST4e8hh
zcBghStPHBvmsO23ODismcfsB/88qNTn3LbYO3FOFEIfmgIY1nMqMnQgKc+5WnMQ
s5ES58mOhVrhtZtrQI8TG9FMJDdWGBVPp4tqTAvg3uunLNLIfX42glb9ZnhAOOT1
TGr0gGF3sZ6koaBJ/qjzF2Fy4IoSoTzAIIBCX7/ihZY8WRio8iFFpag7msPPaH2j
B6/QWZwdIQAJGmbZ/GwHnlYG15wrj8eXWOacWh+DHAg/wqAkwOZZ9EWXpbeToVr9
ybNXksA/xKIFDFBwkoWCsC0KrSP2PgD8ktrFgdzZPzTRXlLuDj3dNMYVDnG43cMp
XTHH8uigUYC1VfGma/heidIRXLzr0i1G2md7rNEYKvs5Ce0HwqKg9KnPccHwWSAa
L/Ki6NlF0tRSmao3iwW0kiiJYD+J5zvGcCtKeQDeUY05R5ZCO38pCE70GvcyVoiR
WaI5XWnPCPlAXwdcQ7LjRQIEzqfQUh9AToD94gqMUOsVWhO5gQzpBeJdM0wu1djE
oZTajgxBvzKwZz5KceDoqb8WhlwV4P0XbSAkhh68T50+vLKqvyy0JAACTLoobARU
RsCRZvc7xRt0KAx40XMBspGSDZyCiX9YQqqEDf2ID4Tu8kQszdoSYVicEtL4NdLj
aJI9lkt1jZZf24KPdraJB4UIoPH1Qy0zJxf/xQdeAnExe9nuu1KuaWMlcmp72wiE
X3f1K/OQrjeBiOWk6PpxmHtUDcMCCYw2ePT0YT6MFf8vPdv4b3zRw/AmQmEtrFnI
xiHa/ouArOM2EneNFx2fSgEZBYcLOi5MHAkJrtTCO7rctiVWpLPTBCSTZyyhVW/3
WZXv/CtDclXVfv8HOfArpdQ5DEr4VJI8MRq3IrjGWunjDldqlKBITCHM9ZjQJrES
kvqSw98ITC6/etXfHaHccaRkwQ2ihN+OZnLzkKSy0FsSkZJOSLQGRzxIquSIy1yE
aBMEtmzQ+91F/YEubfT0gx0YIO3oA0y0qF5x+5ybb4L2V3yFnvbYmUKs2AXqM1SM
Oo9XygNUt2jPVGofdkW31gwLeslNLcQtXVzFxCpPQQou4Bk9urc6ByMBgcGtSx+T
XsC1HdhqaSMgH2p0BatJp+hcSEWKgILRa1x4eZm834Cf1B2qjqBEXvC4tj1t8Sla
9uwhBvwwxN0WAVPX6VlV04uWo3KzaBDXGVpCinoBhN8jYmWEQvqtL/wQrv1j4HlC
ovqi6GsSF1yJv4ZHquaIpc5FfXIMSm1JEv8DLoT+GOph4UZlRJL8+nCRbBuoAXvD
SwuB8XJKEy+JgWAXqixJC5maHwGFPsMwf0xWT+l0Hj9HfDFAwwSRMe+K5lqoGiYF
fAN2nr6ztqYt7jD+rn0nVMx+Y7X3ufpeCHX7kxXhDSS4zL9RHP5Lw1yX9YO4YpYu
qyJJ84i22QEQ1Sq9L+r+hoHpWLmprFp9PALyM3/GPXfnTUtf7CDYrqF0TyWaPTw/
XikETXCCpwx4b8S9eJ5qpxN3V9UE/L9iD5lIXt9WPNPa/7+8zUwfjDHnMN7qLsmx
`protect END_PROTECTED
