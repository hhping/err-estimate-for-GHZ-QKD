`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qmkae9UcxYt8FhxCnhbvQLbNs6ndQ2WkXuPP45mjXVlH6xX3Qwc/GTOspCSBv4X2
dR1Q2xfPuLOCTuoxktJGwOI++3lDHWpFVe8jUAMnwd72jend3F4ojLMx14sCdUFU
492NdaKldbOMWNY5t0brY5x7GhmpVGCdh93CdLMB8dDz+trf5A4QxlvC+W2nM16y
+XoZUCXp7fM8X4o92YFH5Nclao3z6AUqz19c9ySf/D6QmPP8n48fb4f4Q0UmGuni
c54XfgmU/5YIP230TnrpcDL9OCHTqc5j45Fjn7G6O88FhMuzxmpXuPrH3kybheH+
SWCEnZZnMxCfmpgX7UIqj8+5AV8SwFPeUKj/6tt/ZEA=
`protect END_PROTECTED
