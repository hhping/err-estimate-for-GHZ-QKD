`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XDYfpPbZ1njN621CRwxUHp3k7ahT1RXok5y9fl4aEjEJayDsJB1X6YHaFJ7cNBzp
mD84NQY/4qzaTr1B6gxGpJo8pOd1h77vHO05jMW07brngDrwcVcxKCubun+9Sf0T
RwBZ7d/+QSArcj6zA38CZ68EzF2GlorRB+BdXAQd3GaPH00NvZxEh8L1BUzVh7LQ
1fmu8odO+QF7kDjOvS0YOeTTbdOBsIYLAeZ93A21DHkcmnSdlr1MU4zVAC4uSsSk
Qo0Y735Gsgb2Y40o3t7xifD00RcCG66GmNEQswUBSd+R87kjFUhGjPK/E2QFCa62
VRDkUNt7z5ay0RbRI5NhdRzlhWWpnONL80qSX/wtQoSRgsKdYjZ4bibbVgxKyypJ
Ln7ijql4HvXsBNsa64EHAy5k1oFS3luWOczT7LhXNyZmiri06xUtlHfDyFM+MXBx
hYaqQRzfqykzegVsmnXjCA==
`protect END_PROTECTED
