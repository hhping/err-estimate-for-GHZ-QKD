`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2uoWG6K6yG0x0pqd6E+XcebwO0/+Yo8cLdTLQAyY5qKbxo1SkfhbdF09zh+nCs6v
Au2v2sYjP2tCVDMLCkFCO3crzM8CXEC/4eb1uUKHxb/Q5m+OR/OzV3xl0neGkrxF
N+HtmzWO4lPX7PoKonzHtkydj8VU7Sb5zH7dwod+tMErrxUeGddl0/OionzGW4N9
pzNXZlgoJSg8xFhutAhNrlE3aDWCEtD6ysUohlhiNPFMqgKYfN9p3qKsgq2F3LgH
cmSS8e57LEiJx6MsW1VNYZeObtFTDdRXG7IAppXiCVChEAJCszprjMvq8kYAWKq3
xtnuYdI2KXMXNOrjr9G2B7aDTwAvE9qroL+P9oGwgWGdxJ4HIp3UrW2lbCd412Ky
fDvN3QPQ7UQN9rKFNQs4CV+oVx1YR0nPnimNFD1h371QbHal1KKtZh3nQX4whkY9
+KGzueoyj5O4qWWsnLlh/9C2JnCTpyRLT5jsLdQc9arkeyC2C8MX8pzzeD2HsOGs
y3S50MqdP+T6J/5E6ZFYTyOZDZzs0Qt+N/vDbG3gzKqmnQYyLFzvRCaBxcvKLF9x
mzef+pm94FNqo7CtmGedppbMBrr/b/SoWPv7xii3gezMIkg2pCybu6qjIPLc/1BO
Rx3h/mdEFnfHxI0rcDBlJNv2o5JLcbLrXBsqJmLbp4Z32fXvAO7x8nhskvicTlPJ
oc3dfS30ais1Dn6MTb4jq+4+fLRFitXWME2w6BdWooeUrPScX0/KTStjaA1ck8tL
Wco6asp1zWh4pqqznQwmEWZHI4j1vuQeD7OBiawYiZKfPdkDbBzKDBTZ/tDBwKD6
zL8BahqzIpfd05GHPGc/Q/IjKhRiJn2Omd9SPD/AeYDGG+uHQ8agTEus+6hNurkc
GLu/gAfxJTWQZHXhBiEEoCDBXLYlZ2EdQRBj/Un+jMT4Vl5u0GisJa3XvW6X7voj
193kgMtHOu9Ms/kY9eDmWdSFQ8/pADBNnbgEjaMyiw5VzfhtpQHz3Paa3V6r8Let
Oilf4v6FbT6p5/WJ6qbBCC8L5VXhqjyKxjOypmC876S49QBU6cyOmM5QK4PrVKBN
IdmrXPYK1cJF6PLuYGrAY+xFVaLSmAllvKX3vPAJjp3FHObmh77THybDyfW2KoAS
OlcS4lxvGXSZWzHMNAhPSM/7n8itJdHEC5oSS+hP2Q/0BiF7Q0o7jK3+Z8nJWkBT
xAY9Ze7zDo8gzJRbsK8eBxT+E4bJ0nlH8sX7oWKM1NARmMaaDlFgRCn2ffRkq7Ns
bv7uGm6tnIoUTV33SAIyXnguOOMhlxC8p3N0cgjg3s8yA8w61ny5cFcCrzdkWuZJ
7pv+ooD1g9PjtJbCpPTPbgVhzhpsOqa9L4OA5YA6DpS/o1np/h04eJomYScKehow
q2TMrezAVECBkSGZcyuYNuWhDQqH5ib6jL1L3opJC+H56oWfZv9jNZyzFElgBNYT
8BAX7Fq/K69lnQ4Tj4QB8M7R+sBcZBUdMHDq1KCqrieRcJhm4jSB1mUpOzfRKMqq
N74xjAMoLnkR9qlpiwSbMgyWpjJrjmbPQQf6JQ1bkaKEREdqrvyis37gRg8H/9os
basaS2le3edKTU7GOih3SsSXolS12VmfItAJBH+nmqbQvcbyqYubUqGSWKZdsQBW
UFZa9mY3n5FURqv0770XncuhmifunV5wcIsjSXcKHj0Ht9/W4Ky+L2Ij8bJW0sE2
WLoZKb57rIrPH/BhTRaRMjEXo+vjkVRVsFih2xaiOSy3WSiCTpCL1q+YE3k+Z5TO
H7qaLL4n8P4Ag4pZHHahGsSLgiWiz54yY9VLC7ymaKw+lQhiIRVqQKWf6vE3s5XZ
N9Du1uuRU5XZ7kkckaiH21zKZzfjhDDJOvUBCYkAGRzxIVBfDTx0aAV6P1vGemP8
5LSvMulWnOGHqhxjXB8A7YSXy6WCl/82cN7ar4dusJeHnraEwkgRrhZpu/1VTKku
3bb8OTOhVjDCh/UX/H+lHvNDikNNhQrCUiMCdKD4VryDUnlVRjXK6xYFFRA53syp
JgMItYLLQ+lbWP9fMBQwfe3UJBidKNqKiMzCLFu8SYnuxUB2omRptQz5IdmE3EqV
k77pB3VG1FUqEVWX2s8PdMe6Ium3T0hrPqnOV+MTciOzG3w5M7pIfx+bnwDdz+sW
PQ67483g7yQ6tfhJnY+qkUxcUlJKmPUtCWR6uU+P+BCLiH2FLEtkCUK1CHR1UuHj
db+ybMoVd0fzg6SJHlmdecGH6NYChkR9pfQa7mOlBDtRegbj416CmSfGaE3UY0U3
79FlYURsd49CmHAyzSdCeXCjBYxWjGKI1mcfoY0nSHcXcatunE8fw2B0R7Ndr2vL
7b9Hovk9rcfuJsiW/bFFaYT92OtVy8dI0SimHHqIKatenWUiOZ8xbUxISeJ3ixb5
RFHl9x6I2y2VnZUDjQ/v7ofpdPbajyaUiu7MBZCun2ngpKe7Vk+17TxMmZeMHYGt
1vbclqXsA4ByWNmg430nU2epyGL+h8mQcSGoX62OtCEFNWBqXBzILPCbHQBlOoQy
urSqiI0vqQSXejCkc1CZGqBhm4XuOVBvH5+ba6ZozYH/5g6/6e+3ZTO0ndqGaOy1
`protect END_PROTECTED
