`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CMZzRsONfBVRld6oLYNQq2reMGy6zMtX7JaCGdtxD+Tk/NmJkX/rtWmc8wH9hmlL
3HHBKbmkg2ngNPN7AQ/fR00njHgE+7bZQJUYLSBG2Eo+jSPCNAOQZv186/nuxti0
XNnt+IfaraA7op5bSBaZSLC/Jj256VN4xh2quRKn7k+XAxZYg7s036Dr33UjCPqZ
HGPJC3eSPErMbgEQmPWOLHrXT7IywrokKCF4hR2Ido9+JlrveRfjXzyAr1LCcYKy
AltuoFKFF8OLv3MuL5yUefXSogAA0rQLNai1JL8v/QMr5JUA0RNjTze2MAZo7XbC
x1p2KLJrvf+o/NUfkH+E9jjIlV9MFVBrYeCjknUhol+RRb4wzvCvR9vTQGmOMbvW
Ya0zyURrxRLcgrx3pg7FZ0K+rM+W92K1hUuq/yBthbZHWF92Hc1Ts8kcWX0y2+wa
FlnNvurokLSruBB3S7Md+Aos/uz/Nt4kjHZsp/9TjPlwpHuxnlzEw4RgblI93uPg
/5VKlOuPIaIKPzgeu8T60hApKEuuWeKLmRZFIxciGRqjFBkrvGUZ5QbqfFOw8Xgh
wD531qaUt2yt/Uy+3ljKQkCdOiaV0LqMmXNXalanlpA=
`protect END_PROTECTED
