`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
26FZpPjODr14g1S6+Zz8mbxzJgRc6IWl9kIQvK7BwHhTu7rgcTRNdB6mDWrVUbXq
/x3Amkn0gcA0xt3MILQZJQGu6xHyRU7wr/qfzY+eF7hJrZfmwTRVlM094WyxSeJG
dSKnihQQyvJEDfdEIY/0b7gNWMv0TfD82Qh7fA7SFeT+EBs2fdC+hFWxzohvOFgz
oOLeEWWp0sGJnx13NGWwWaIJgbGey87gVRc4uVGBOLk9nUZc0o0dtj5/7HdSyM6/
cddFxg96QRGtRT6rOJwZpMXd9b11nGlhTO5xjfjo3ZVJnQu984buAb1rRx455lHY
PjPMk5VTpZqQPHrsTl/Z0O3Ov/Vajoasj7P7dUYeW3IYd8JV5XIpT7F4uWZ0cFH9
2XvqNUPisfjdlbrdGO+pWyLKT83zUU8lQgQBsbclSvGw6D7ASufU2GqtPBXie2V1
Saknh5oDe3ZcnXNaSHh+GQDItZg9oNBsAaWA9EjJAJOvT5JFIKPw5Vut+pyqaT2A
ZvRQMx5xdiuZqQiV+gzJJs4fdaI0pwMrXaeOaXUm70AufO9i9TXYrLRmQlYqGU9v
PBMEmqwDPCM2tIMC/OY6cQRh3X1ttgxl7ZzHasaxJcNzd7tafYw9cnF8p6xKW/1c
qrOYtCxqCGGzI+/FHpIuEEcZQF4maKbchhrxgU14eJgoW2yHgjsAuHokzcBzMrub
5kcfdoyee1mFJUpAkom+ZMgLdSvEL3F5paodt8Kmh0SVeoEwTeCI2GfCcHFywUFo
+Y2EbI/1vU/is46KpyfgmhIeNvmw47e/YqwGlLCdKeXgjAZJZabOWpvOpHcLE/by
yO8iExomvfK3PS0MP4TVb2oaiXM7Bl6tDaYfuHqu4rdBtIOIeDUS9IZg34OfZEpt
HR2qt573XUmk3zAN5ymkOcEjPtJvLpbAz6qqvwLRJnq/+f/YEuUOEZFcjmGUq/Nu
I1yWEcpKM59XutNnIEJkL9oWlPdjlS2chALYTCklPoVaWtvR0owEBEB1MUJY+v24
1SEznTKVy/6qAIcR/xoKOcvwYtuPOkEpcjyrtPP3orMYrx042kszjEkP8FG9USw7
dgF98UDhiAR2IldNT/yVz1uwKAaMy0EP8hERwlJuB1Os+llaAfEZpTjmhr9MAC+/
WO4iPwhRwTwxUTSFpAYcedlx48K8vKpyjYnLjxwKWLF35py2EGQt72cjd3NbFgBy
JKSKoTjZIpkfCaEp6xLrEU8Djk0nj8d1ekmU/ky837jTvbBaZ2tjr9iRPH7gfQA/
`protect END_PROTECTED
