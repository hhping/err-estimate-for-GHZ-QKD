`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4GaoZSVVfWqGWmKXW3+2R7yUk0YjaHuHRc7O5zvFVWyLdGdwqsUdkGGEcBMa812Y
8HAVzc4pmjT6SNmFPmA+QbnmjmnDtXA8OqeTsJaQ/MuJ8ID9z6ykL9+t3B6oFfRN
rMSqRszqjUGgZI9jf3NQUsToLITemvBu9X2BTnGs3lReuyu8GHc+cbU+g5V8JehH
7OuJJifd8n+DchWc7yVwarhWw0Ems6a+0EJHuBaokrsiTrnnuIC4jegbu/KOw09v
IjgJ0FeR4zqQ3W16yJsAwctAYg4edVbH3xRZLTAZezfcO/X/Fl3i87KyzXFmaW5D
uiBRHcXBOvvSmAqZnd0L8rqVA3JQA6pbI325/YXcHR9F3bmja3HZbpCeyYVCtFU2
bpCdx13pXZ8bbE5IKh91/o2+JBMqfpV1MYMreLU/6kzMC+ASw1oYJHK/dtmG2Wz3
v81ZXMBdX/XOorENi6PTmWcHiB35Cvw5JMB5NnLgnLEpE1AHg3VzoUH+6z3puXQz
0DUa2bL5jhEmYHg2eAnlIDy872uR4wNW5VlXqJownuAZUOj1NtZhXP+fT7081BbX
YwnQJiWk/Hg9lER+6LfwekiExYNkr/c4vrTarWPrUMQcD0QA7Vhj7g0v/HyNPhEs
Pww+BQk7au0MYgju582Oxa+0EPMofzljCTNwqepgvTxEZmq+Smjwnyh5zobrLmit
FGKfSaz0Ewjnbu+9pML/F5hyrgN0XtjiEp0pXswKl2ll72OriHXmsIl2DtBkJLoX
d5t8l0q9UXElp/OBtVnOwk1uNL+iKUHPWnjZsRyNFRu0nhpn06ipwhcJmfFcaR5n
t+Q3MVWUgYZFDXEjAHmZvIq+OHzbnAJRSgnwGRDSaVzeoQDkjW6NLV0VpB5U5WQ/
8Jn94bUyoOc/cdZ3QVi3o58aufGQKWrjbaTAQ0rVMZ2lbaMUYIRaAJSuhcheFWYk
/SUfxcFsRpOChZlgzqzO+rJskOWA/fwOE8/1dXud3cALwktGC5BQNZxXuAqVU7dP
yaJ3KZILG4v45JKq08nf0Bj2UXp/LakavSSaRDSGL5aTcQsDY29c3Zsmo2tIkk06
/twnAPU5ZUMhMWoKDAanCp1wzN6kRa3x6QD4xrxYgLjQXB5rVDXgSFRhjqgCeH11
YTBz/1+Lh7eT16WUb19xiodOs4r2qMCRrIO1csknuh4PJ8AvX4RHS6xXQZ9vNI52
2IWy2l+bSG34wG3Vh0pb1JkSXvqsKdXnFT4gCM2yU3qHClw3+oAkGfPnyNGqIpKv
l7NpBPR12zu1T8mq0Ug9Qw==
`protect END_PROTECTED
