`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ocIuAUayiXHq5Eep8/gYiEMyaWMHWfRrpjimR9E0t3n0OK+vMOCBOxiF/R/7cm5c
7/Ui1hOHBE2GRVxZoPwPWAu+S0WxKAFbyJ9mR4ob0HpaNsyoeFOHg2ln97qGPKWI
3DTm/w891kxTu4a7XmF8va49Jskmyutt6fUwqIfG87y08WgY8A9n9hoKM5r7BGMe
THpFw1p1wcbHyXkYec34xEVBRCvJ9LVEShjms89wZZEK86HgYesHr1rpCoqmbo9R
k2LF8VU5bHk65GNqtO0IF0MO0IpFsZVm5lCYzaeFS3SpU5bdktiBgnn3WMcWcD69
ZLJuzx74NDP9zGj7g7F0GZH/9/Nbo8oH6mIJuC3KAzFhgJIoRl3ZDdZ5cweVuNW7
laHW5Kec31NDO9GkvakDUqMibW0UvPCySmIxdenrQgFd4egiG6SFmgFWpdvyDg5z
zTafRQRa8h8ttTZQmSHj9VymPWfTxqdo3fCkPdZUYFx8lHzps16DNQRF+vandf3L
dzfcljcDYNV9Bizt505z2Iesq/iUOWr+pzbhZuzJSZ8+EjteScdi1M/Lv58i2SZe
`protect END_PROTECTED
