`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NoEL8YAw09STElLhgE74gkByCRde7IR8mr6WDyWNlPERIoZN9Bf5aiMwcUzzon23
sm4RipZzJem2aboM7CvHWm89fv93XOlsYrWEet7T3rb6Motq82DsNPXWc7Auno2N
LeCQBy4hmS0lZpG6mDwrc+xwQMWikHkfS3/EAIoZhuAkWycXihUMkfeHlnTCLa3D
Q/VmfyUr2rm518isUOwtLCKDC0/DwdU7rVz/Z1tLYwUxWxCqL9dAk9WOZONKYkiV
7PYSik9KLCwi3VYwSmq/sJSsOa/IOygX7EQ/wQefxqsYGYqAZFWxea89oG7AkXkS
/UVH9RQ9zzs7yaeHhQpovQvZgHnAk9I0wqijcz8WBc8j6eIlhT/RjXNGbcNKG3oc
MXArGt7ox5eyo4hvsQAOpVBY+gMrFlFv0LFe1OXjabJaRiNfbOXfQ+Lunt7aFbjt
ABSZDhSLRGO2jXgWt7wocibwUPwYUmhCD4/6aekjBioNtVbe24C340vvxAJn8Wul
hJESKfOkZsrltRH1I+Kxk93wdO5Kz7EblxIU20CydGzqx9u9kKCl5DWYFLXqgRnf
7/6zoEjBFycPdot6T4CQFrGzCiGcmddBmxPTXhcV/rs5muhSrEYF7Lmj8qNYjX/O
z+1gt/MKLGey8unxhTnwGmFAGfDt9azVDCkTmT0t+Zvt8smyMt/zev5OgpaxvsP+
4I+DkCuyqpEib+BAwJSAgZiKZpmz/Jgzzr24LImVUMQeSHumuKWn0+5lhBTrERam
N07LkXzAV8y5Y9h1SxM+qI/pqG3V/Lld9z06fJ3olECpqZfI50rXNkx8usR2AfBl
Wbv5IeBSZFeciKLepYH+GqQHHQH+nNkb9VZSZr9Dt4jDk7JwUGyorEXX/Dwitec7
sCEbEkYmLVgZzIkTygNByg6A3ZPHXcvjtXll446LJEGChJc6JItg7o/i0h9TCrvG
LA/VHajEowmoXS4Lo4nK+pYtZPomWP060rNMpXSmXSDi5sfwh/Q9xFRy0BP+eEe4
dw0aYVc11wp+1IcRm2JytGGkp7903bxD/FaaUzR//s6S9sqskwE+oBNh4wD0OF3Z
plA/X4bDZ/eP8begFuV1OcNdJ8Mq2DSDt8bUtIWvgcYIJ9Ud+gZ76xeAUYvLiKDk
UD/5iz7GLIglPI27qjRMrsvS6p++NnAKtc4bgiNnIEtAt8pjvl4VUUdcHDZZITa4
YtAl6k/4sM8Th8Fo+ziEcDnIxxzSF/mA7Q1AF0OQlEsfhx78YhfLoWQMkCn53W7i
tSJRw+pSzENYtrS+gH7hvGUPqLWHSYn7nAQCsVPaUwqHcDGwagTutOiD44PRgG24
df+fk+NSMHlJz4WwFhQU104mSZ0+Alhl1PMzrOmKbcXb3wffAlW2gNYmswyZXz9v
EN64dxQGGo5Eyxqbw61+Mxa7whPbNKrqfXPlDJJuTRwZLv7mkH+dBDnGgxTh3TwA
UAZd2PQCu1BDFwD+DCKiHhhbpjLaJfotDa+1qv6sfZ0BFzphOrFocXgB/iyNUKpF
vdpOFsR6SyiiJv384XtKeV+qcmhxv/hUcG02Ag+DACSQPy3xPY6tagZ+mr2IQE0Y
hqoAxoOhpwsCo4fAlXufc45Xu3oMl4zrfCsqMwRBftS33Tf5GKfBPUrArUHg8jVv
AJS16OHYglJ/oHflLZ2pe00uIDHxalH0KM7AcaI4yghEm19DarsmRh6oJoT3Eiaz
ZBOXWKO2++wO0mrq5wEJffrcMz8M7nfvSWOnOuBYNlieZ8ihRGyi4TaW6P8iRFpK
83Eaf2HzcZ9Y4fzp6b/cnxsfz/1WsqU5FFkr6r4XRRtaC/l5Wz0ojTjfKQ8x8m7H
huaVcHQKXLJRhUaJoxbbRo67QIb/Mn9O4AhzbmOHDw51O3DPf1ezdmPkA4+QbyM0
7ZlNY8cej6M2GhAiObTB+Tan8hEj3qAxWZq9OEJOsLHcGxgtHCOB3Dtjb75aZJwH
RxmPlWGgmhITpkiOBias5H5p0uOjZt/AhOcRKTHrLahHWZN7ucFiSjbndKkHSWca
TJHFPGuU4J9pgaVXwy5hPaNb5Dl6P7jbAqATFhuZYAYvs40njccZJGK1sTeI/M1k
LB4PRYe6LEemr9ZD+Di+GUJ4jnzj7hlWqGLx+6tOHpcl8CHLl16bdSToi4899kI3
7kJr43H9SbuIL083lSJnEs6PorzBb2AmcIx8HMz1DTmI2r9p7ieqYcmNNXWr43mZ
Ovm7Z1t2thBXNWXhwMMOcNfUffTEGoUtzPr+pXebn+eSS+EImXPEss8YR+ZnPb0W
W2pLY9d6iW2qw6g/MnUnrwHomlI9qeBB1/Kel0EJ3eFAnB3fGJ+TGk4EjBMBLOcW
nhDLRuA3u42+RVFTvkM4WI9e743h+1hnmbfkjfRG/KCbPvdCZ1kt2kGy8m8jx9Gn
Wo9u4i1AkNTdeGAc+YycdWDptRCADJ/I/+ZUf6yh9bLDSujGuGUW3YJcm9J2S4g0
ufbyrghibSArA1sKyK+GFnellUonhLoiTa8lH64cilVUGS3dDeeusjrSnT67ISfg
vkyWJBZs2smVmJsfjU1lo3DwYG0rJv+Of8kHo/uljdalTHe2+0uT9M1G30n5Xc9j
3FERBbNAbOz+8pkBLJUUG3YGSH9kvm2ujjFppsfshxDEya7SE/gOLJxRpJJEi9hC
IcK3DWUD8aK1c+xCuOAWd1obCp9pwdR0Ay/cCLnvefQmVlERin7f4MHcgBFhcPSw
vuN+zJzJxxGP0NzXW6ASJIAyvS+i6qw8DwEaUo6LSNCDYwtqU2PlZ5RXiVONHNOT
ejFmtZKkp7/l7q+eW3Cb12ToyBUui5kMxD4/PcxbC1vt4Rp6ouxVMFD84xUgl2ml
CGaErWl7YPvN/1rqbhPBx2smuod5kjLydOfPq6MlTY7ic77fA8BcJPLAwGDCWIhV
LAoMkrBkYxyhPoIByfsbE8yTFb/7LM9fBGhEobEqlJuLw7/LOwrVDwWECEu0T2qv
kp5QhoYMvuEorWEAFAJSRzVP0J5nKLS753me54YFv6XU1EPU0VHbFYXw0Awyj2Wx
1lM5iova8+1U5Yrwmvg8jA59ecP2JdL5yZoJ0EQI4wwsV20s2NHUFZk355y1ldJ9
GiuSOvJMSB67/85/zWFp1NSRA2kuIcJH8BWjEDrjsP3Cl3twhCu/df1QGk8p5rHL
`protect END_PROTECTED
