`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zIw4GWK3R7ccwHv5wt0FAId8R0u7JzD6W++h4ws3scpgD8/vYgUA2ae3eSlSxHlO
9dU8G0h5aD8Zx46mcqmVOP8znVpyVDmRxxdvKy0J1eMdXwKuKNcvHJyNe+ksMupP
osPrgiO5W4Til+Dce33+Knf1aOB2xTrww5TJ2FuE5P3VTK+wBPYoN1HQbJ/zhwqi
maMuGa5/tzaf48bE3FYdOK2B3BxA5MT+5ESdFiesOdJ0UNklU2FdVUFn/Pa5fV5W
Wm4KucY5zZchdcdBc5WNR17ck/y1jjjAc4plCtXsnzJylP8rzUqfgbv7lk+K9b2q
J8qmQBQ+uVVxjL3qz/TBT8pRkqtwedXVH41y64ZmOsaSuVq4roj1Z4c0GQiKhj++
UhoLCTpa+1vwnay2DK9QlpUO92/P+w11KxwQiVHnq0boU+3GPdYurQT/IlMftFX9
AzqllpWdLO9Jq2Wk6k+hxWStQbjbv5dmL7FirDwcbGPb3fcNorD+6GI0r5ImpTzI
w6WN4K6CXUwPoE0XHG4LtTQjnA79oVJYnolU+jdEFUwl08jVr7v2umm/UOnVmKgi
pzJMbrJ4EkO+IStzi7SIaCeQkuC+KG8l1Rb7v+HeIB/qVunyuxXF19rLxUMFeXar
/4pmk+ApRUubYm0lB4xKzJYqW70myjp6/PH6A7f4Off/TYiNa51ajQh77IvdK+Yn
`protect END_PROTECTED
