`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rZaH842yuF3mCXosERxHjMMKz08kt5Xsk3jLak5R1skQy50xx5suUAdW0BDRzioW
ND61Of/j7vdi5AONkxQ9SEP6lcZqFfMYTomwA2quvCVLpvCR1gUtrpBCZZ6hKJvH
hp3vs/SjDRVlsseKEX2XbBQfiaL0pNNBMnTDAJOZGnNTzK3/TPbosVluW2aeP2fH
DX2wrCm+z8Q4+1Y3NuGr/yW0OguPXvOwUGb3XsBhYvll325tVF2Sx3MJ1Dv+1hMq
Wh/ZW3DWCc7O1LuGUhaTDGW5I1/Sm6oQq6hNCvRVuVNP+wQ5MNh9kMt2RXgn9PbY
nVJUlk4sisO1TcavsmJkQrxcwc71MRHe6wWdoPVqXlLrln+3m+azwz5fKPYJbiAf
fhu7XhNGt9VJjFZtW09kLIawCfdonuGAL6M3aXKMTIRlL0hTcolMsm+qw9RJwAHZ
wq6Ph0FfC04V7jNJXALdI4Q5/0VEIm8H5mtcaETobjLu5SeUgYwluXoGIOiaw5fr
IjIBHTIrwb2xuYfjonjxqa3Y4aVMiLajuep/AWvEDbuUn3IorDj7H6/FiUSfXzXQ
2adO87ZWyoN+6x15LHI9XD4SRx1ZVVnJjXw/7wLsdxABDIIpi5rlpXYWMaqV5x0J
Tj74SXiNW6mU7SYS2VFQu5ZUOpAgcpDLHxD3Nntl4FiMw7dn9zUkEwpT471AHkds
0UUisn96jeIBvwreRlcIFLDsPX7ciDLl6mR0TyxiDDaybF6w1AihPx5Q7kpf7tGz
kFbDzXe++P4+Oc30OrUUjnmBJvd+3bCexK9Hf4I8sC1KCuoTWPzTPy2k4iKYDeR2
xIFTD1IU7nbWCL4ePnDti32wCxqyy2Bek/Ptr5ulW+z+oZGQfHQ4KUZhji3Ib6+8
wP2dJ888GHVyn0A09onpCMce78sooSLdyab3KC0UCTk45vT0GZw+7OxigL4eLROe
v6fFM/LIJZoI3XWa8NpKfrD1hsG5s8LV7ihBw3gN2mkcGoV1SOUMk6RSNpZUdXgT
NKZY9+AuptCef3KtR5DVSq2F+p/lc0LykbRvob33Xq1bFwmxjfnlbNLv1lvqFHv8
2qD1kzMyxUFfWNpKi/nkaAd/zkjYY1VMsk/QozLmsLyFY6WhSt5id3HeTPi9E5JG
6oulsmWKhlOuD3BDruDhs0zoiUsIkkEK8zWC0GxyYz9BaFk8OEd6d9xApqCG7D6U
RZN9A7LFMflMNZwrBgMCgC02E2O2c5vHquetCy/TaDR9D4HqQ8FveqrEwkMIJzLK
uShHYpyz+zRPtVvSXTNvzg==
`protect END_PROTECTED
