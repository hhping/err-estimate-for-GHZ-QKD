`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yG3nNUR1w7nOcSnUww0bua/NGJbQ9LTfTMsWPvGlH64FQ5RrhAwU9a0DAWt9+Bpb
Qg7FQh3/wusICSZTRRFYT1BfQZF8459pswrcpdgcBvg8oHnZPL4A/+3Vemlsqatn
SAwOA9flDR5+RfFIqXc4D/Og2o27+onPwHub/SCPs1RqLLbHjQXDURvXBJ5dDPNj
EilT3PaYNSyd39QHg/C+jhnR+1617UVKDSP/NavkFy9NbNkuklWEYmIFTTdkC7wN
MRC+yPR4I38UPz6/ToxnpPXc48b+P7bByKFOqWWeFRhTpxbQN6uj/nvBP5b97lJK
spb65PwX0aJ9A6yP132sY5EjvpdzvI7aR+nOrDIsGQwBEupWe1W3cIaQ3i30dDkb
MGmC9qpcc3uGlQadweywLYPh3iyf960cnaySlr2W/OLCW0CaiS6drZiuwscmcCP6
iDmNzmgsdP8e/VN7mqgkH2JRfmvW5p4F5qkF8idpFwCvQpzB553qtXFvIf0856nP
r23BoEsvFVT8UhiO1juouZqz3jHeft9ZAZtGthnmLih0052gGuU2qyP3LrAedYSC
YlpsSTrrmq0gNQxkv3AQ7gxqrne9uAJjKn8wO1NzPF5uCNIgb5we9O0UtYTtQtZ+
kVChViJ6tW+E6wMe/aixMnM9Q3X7pP2mvAyh5aFFJsMZjhp93yea69cmay3WkmwT
f0Js+2vehXXAn739HVh5Nvij/7Lw0fPHYOu7z35S2/Gqds8hTkKvzrtMPyawGand
ymzeM8Q9cl4HveMEdchqXqd+CBGaxQK3R3+R6dW1TrZsJnijwaH2j5gft3+QqyWH
32gwni44bavPVjrqR0k1NHOjA+e4Ua048V45NSsGpNBeVk0iiNptE8x8eZ0AmdoX
WBox1ZDHC2gnzF6j0b4FUckZtVBAKDOu8km+R/W0ZG4nSvtPCUpvinxFsHt3samW
U6RP6jcCIQ0GvP4J1nWD7mwDbWIrA2tg8rg+i+cqWqhlRx5DTR1D/7lyLC/p3vxl
i2sTiZJnN6H1p2Ex4nIPw2GBrMHnn4tYFqTsIQOznjqWShtyUEtx21xaIsWvKCWh
B5Mo1AV0spOMb34+Q69ja/wyQuo8a7+kDWsA3BTWiYhM9ek5BSK+i8wLV7VOBrbe
WEGwvZynfVlO16Nf+atwanyEkVeY7e/omzd95nadxNc1B407UdrNIWHnGUpDdq94
Xx6cvb/3yGSEfdcIxa4uICTOZTCh2VqQ4wC5v93xz4xeG8Crfzm90rblYL/fj6Yz
cNsrWaclXzpBdSS9blw6dDWQoZiKM5iZneY/S7U1JqEp1oEUzsu1NCNUS7qNk6/C
nvYi/0u0RhKGA+9M+YGZ6UmCLWKzqtXUGnGrD2BMKKAmNmIwys/X2LwOttkAHmt3
TTaXSI9MIM+PAUikyUhPshj8LQ08ih3CWVT6aPzkI7o7+vGV+ytt+ujYt7wERTf9
jwQFfuKu7KR3cBS3HtcFnTxu+dO2bywSg7J0yeYwQSjDQvyFHzHR0y4IJkBMRbRH
X4r54so2Ggm2BLd6Z/55ntpSbC5mQueD9tSnXOlgyyJoe+S/7SjwXdz2WcYu4Mxa
5LByoT0Q5qD+lk6qVhqzr0ywF/i75up2SwZzl5Vc5/GBhtmRA9q25M63CuCE/44u
5drkXW4jI/Rt6/TJWJ/IG70oklKyhxVP7bF6yg4Ucjr+aIyQSHx6R4dPHxypzcH2
CZEhMchI/l6p/TvET+QKXpImAzBLQNJPkY6l8rNTJQo=
`protect END_PROTECTED
