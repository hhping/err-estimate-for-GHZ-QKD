`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5k5iAiQADsjyBob+Jn6BJj18F/kPLL6NVTmw9XjxCJDHX0ddZn8V7UdxMMQ7r1HT
48vnGWR170ykpfPF4yKDFZy0d1kRmsofbAJZQxlbZmXw8npeZxRIV16vz48YcnOv
tkXJwH7f6n+nEv92xpWMrVgl+pN52mIpzFXtok5gY0um4DZKe83o0omxdi+kUh6c
4tjACyiAbHqb82uoSgET4/GfumYuqpyLkuQuULu8Ptw3fMioo+Hlu+ftQGYCp+xr
gklnmJn5SlorNU+DhOQXxfqD8p19HXR4rwMcxn0cb4/R0n4uG7QhU2u5doOZaUAj
+uvjGjYa2MxeFytf3dceGxtvVFVkpSChUkHo0CDrm9hvLQMum5S9HslKgsPYwAnd
qBYskdsSo9TsX0+eOdDle9ltWHmtRqCuYU4BlXGueNaPsz5+cUlPHa/e+xjwGV5K
aq4yd2xdAHn5hxe7qgylAI05aRAbcdJgoPnMXflu7F3ejQmzG4KQ2K1BexWxj1n1
z2mP8HHXY2dmC1V8nxHE9ytE5oyVvw4MZmSoZkfqrCmoj9KI4VgX24nLxn32+eFe
qoWoR1ZXQZ562ET6LqEsqc8+qU3TEjIJP+sAtoB8d6VTMjn8qLBDd/WktPwhfR4g
uqMTk6PYxRFLeMlzJXx5G5Iei7As1VWGkTGPP7OXW38U/vIGSTzyRE81d3nJQyXK
`protect END_PROTECTED
