`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xE02DpCdF95L9aEQu1Xoj2FCpQOn64SM0oU4GZOw2DvizPTT+sT6noNjjwOW5rL3
MX0oIYqTfW5sxBR/N7yjbc6W7GHBW1Zx12bLFGIsP0+pmDgtPLq9dJ5cRdaS7/9X
TWYboAwbm11pbCAxcxz8cFCLk7k4WZwA5DtMpLZYcAX+KjyfWv9TZs/o3j0yQ6xV
1Yz9y/QNiwEle3GfLShoOABp1/bSpi/gq6M64pVp3CKls/VzAS/v6nsjeRpg5IqQ
G02RlHgja+J2onE7cEtndby2RFxxRBqIr9wClxKQq86HXTT3rLVDjgBn4L50wIq/
dgqaDGD8XyVOYCDfkWu/FRB3UqMlmIWdXtqizBDsawqbwaK3FSXS0vuuICgTWpN9
BZwkweKPsZXTLALywfXhvZWC8R/zWSQAatUfzIWNtMo1ZVGHl/eSQCc4uHQsoWmD
j1YzlYCRuqrzYuEXpWBtdnNIdz/l3nPJJyQIPfME4iWbN6LA3VGuxXrsqucNVk7r
BubpnXK2Jim+4sFowS4YEX1HltIsblnwZ8+pafa7uAALfr8lohYQUdGGfzlr4GcK
roPZQXP+bmm7m5+Rg0RxzDVs6dy8h+d+dMsjC9SPv5MSQnxnr4QQaoABChe4wR8q
ADXd2E4G8TgBmKoNIL2OELCF4nBfDdvJnAw5olGBFKT5dEeb+MLjAwTwkQmBvQyo
zaGGApwj3XSJQeWxsod/MiZkJFFjQ7lI/hhjxwfgFDNOO2Kk6BD1VHMGj6fjsrlF
gZeXObq62W/cYXp9wRFKos7yZE4yZi0NCU/6QBXZfW2biMEW35kKq5gXWjSF+FLS
gbgd2SAaqWR1Ho33V0KPcnc9mFdJ3lag9b5ZNWpLSiFBXXLbWVCeML23mHFgz4Fv
YQixpEbWm1IAICEk/ZH7ZNQSrQWageO/dvKkZiIzhvcwPc9RU5VaJmyrIIcE4dBA
qRh3+lpWUa9dzpHdAO7c7NiRykVafkdaCZZxcNTIqkJiXf350MmAh2xFnarMJlRw
URJ07Hy9Nx3yE12PuFDRoxQEz5rlSOGrdB5llXhXyecI5pNns37mv2rWeDAlhvn8
MAF5HwlRlacwx7PZDapuFZzILVv0158e8UlWB5FuFvh8vwgGt8NLFDuEK8DMkzFi
r3ktIZ3NpL0F9unAypjcEzo9EHRMXHBT7xrpte6VljwuXQtY2SFOmON9gSU+qTrD
gTx6Yz+4GLhTUvVaOWwLIHbPunpP0dwKrcyHF7XxPRuCRSO3iaFEdMyYRhVuAOIa
7K4CCv+/DxrkM4pAASqBJXYNHxZvXtdCpx/OAn0XzOyUn8aIWd+o8zc152aeO26Z
E/lTVKOQfgOLj+XyykOVKQGKVUOzS/5p2ODU/7hndLUjFCpPbIf8c8lf9OTunFg/
B3CjT2xo5ciFXWtjUrBJkjk9K+x2YTKliuHVD+QPHaRwk/EFCHMbUHb7VPrbCxCC
9cRzZyags4rZcNnDX9voSuLs5InaDtBQmWMDZFGXHy0Hk7cm4W5foh7dsPlOEFEt
QcFo02Ny3b1suZvqWea4vfLVa6wefG413LCBj/Q7poUgcy77IHuMvKa03PKSNoTD
p+/J0UQtbkwQfCrZWY1cBgMEQc9hnkxCvIb4G7WjB0FUg1ycO4ma4isLUHbVM/h2
FFPpDww2xB5SUypephB674NCvle3zfzis5GJDeo6TlzloZinhuBAlVvfm3m1vgQl
lLjV4EQ6fBbi4G2XlN2tDtIIVMoEHgCziswZ/7xX/5HDd7s2bdMIi6CV/EZwxZj6
tQ7CTJEIGB6W/D4w27PVYkgIFuNbcfTPu/Scg3ZqwLzYS3Nck/S4lVMtPG0rcAgT
bHtfSu/mlaKE9deybG+T6NrLpiGDipzT+U80IhC1toX1dyDfGGhL+g5tlOQz0Mg1
zK9LVEJWG+wcDxRCf76LvAD2wR8ZfgpTc8MHkI+IFwPOmdUNPUynKBcsXFcsZ/q2
Nc8PxyKiugtCM4GaofSndKAK2IrPM7MNTWBFAnVpl/F4GHtkgT/Kj8FfQos3dnXn
YrYEYZCFh6YfeUnuRtyZlt/3Fjg7W0jwfHLKa1jZOrB8u49XCb5PvMCyI7tg5rQG
ZLRXeVhaU/zFLYT43TYeNaR0fqPKb2/Xb9iSWKHaEPTo/0MEjjwcI/6jRYdzwlte
mhdwHadLTmv50zbZZe6O0H55xzSckL4Vb6wyjwnTIuWM+xPxQZLh7hVMJB8cInrj
pRsAjT8tFhgEdzfrsO7tT6IfeGPT5fHyn44LJECeHrZmJ7OzK6eS1JMLxeS/KzeO
VRv9j1xK8egmM2aS6inPDO7HxrQAMneGB9HtdCzZBb6JjCRGjxvFXTEDiwDPOcbu
ZIUN6NpmaLyd0rKOGN9DKaRUCCDPPHdQaIIpfRmQAMzElewbuMuRvpP4nnCk2V4G
4P7c8s2YZODGtrBnvPewm9kjs1hnEPZnl6lyffTAN/xtnqy4T2m5oOfKesDYvN0+
QdEOywZQfOyYNU5Cp9jnL61cFvUcVJ3nWJx+ZJBPii1x2hID/7StGxzB7eK7REs/
JAy2sYfxaom1TimOvP2bbEYXeiRSzgtxD2C+Fuf1jATTXU28+1rpNjLaJvkSdhmi
5yW5bJmII2Qe2hzRAwBjPmdPayAtd4nY5gv4wXz5r2OaoI7yi10O9DXmkjhsmbUK
TgZNE2QQpLv+AgyQEVOB7H9zUor06Ym+Ty5hvGOhukSrtoXtnMHvypVbhxL31wJ+
rGIQNW/RCcHYBiVypV0UXLld2BjxbIDyphMB0pVnr6pVJ/8odGyKlWMmrg29OpUH
pQy4wh1qkFn6gr+R24Iqj+7e42078KuzSh3KsqoMsqIlBu2DCKoLY4jcFW/BERwU
vFQ32RB9VuIDozPtllX3hUBDhZ/vnydVK4UCJM8/6wLrY7mCnKNh4voWMuRwLLk8
iQ3xD15lGXay+wZd2DwZAudCNa1U21GJmeUPHtNkH3OoPVkwiVBgvhbNFF7N1upM
YjM5sUHTGUuIBAW7bw4Ytr334FM0oaMEgE3OXrbr14ijpiMy1VR9EIAVZMXd0mKX
Rq+6LtnL+Cq6zocBGLMLxdnQkU19Sw8NQjffLNamJuOvPUDbaG/ZUbGhgyY1mx80
Mck+hRdfHClpur3WHgeK7AvSc11G8TW/WPvpNEYbbSDQCnQXqrKETN8VxtbCi/lG
ABQiBVwn9GEbT1VWx2+4NI6FUadooHY5KrZvWjuOUgGlrJ5qfoj+v7T25zxDdSFI
xOhzU2y8ma0cchxVyG0kerXUm5bpAJRa3eFzCag2PBgcsTS7w9gRgXxQCYDkcVoU
yIUIm38tqTKkYDhOHr5jqOz5gTIv6wMdTGwA3maIStDd3fZpuCbjMwR6ugWwNyTj
yGpbnZXrusV9EGbXqU0kFjwmQIOY7Ps5wuBdnxLWqD0m5oKAmpm7uex7J3PA9GyN
wJb3dICvCEtJqdVdglHb+Gn31jcU6HJXty+mTN0IUORnT+hNssbbUr/xBAOFMyTL
bKlp7HXR5sVci2Q8ihw9tfWRylobw6UeBZrYHkMoXyxqmrTJrfkC031QiUYZ1kg+
GxK+TX+QhmexN2FJI0Rp8Fmw1a5UVVD7T4jKj0hxd5u0nXJWYZhNOgXNRciSjQBD
B2+h2ZN+DLQkbNj1Eh7ZUNGr8WbeEatcKJK+c1cl3/I30uNx3K/P3+/vhYacoNNp
kKHsiK9oXRk0w6jxeTxack+n+o3s8riHOh9yFLz2MkEu+YlIQo9hly6aB4oWB+K3
cJzMPwloZXVgf6SivbZUM2HEXdPrrVOZiTMb+zg32RUpf2xWqltpZI2MWQC3O09u
s+yB7hKWJUksQyQJOb9528eWz/TqYAuDEy5niX2PxCaSUfvmFfqb/0aUtBDtaT+/
qzjVFRIipcdIOCib+QLYUVvqRpjAs9SOGvL72BKSQcueLXMie+xsjDBclOOx33X3
ILBDbVyBLv8h1ylq8FWg1zMD+b9Yf7qXfgwVTvwW2TY7Ars/XkcBHrLdklphFSZa
xTQFXw47xA/sWvEet+U7Ibmy2FLt337STRo8bo2MRauykZTfFlTX8/KnAw/Z98cX
VlZqzyvNQYEEDe6tPz1vMVxMFzFTUWuFWYX/WAi8WXtzSI0kg3ivo2+S47REbrfI
mn3aKwMmEtsN9eM8+KecPmBv0aUMu33YsXbdGzzlUN+XyZYQ/QNp8dGEJh68Q5lN
Zm4V+MlDevPE/6o9U9h/8qG8bKIe+BbWysa8GY08GTpje6D84f/zV92Bc2sNeVIu
n3usi1m8adDrTFWlzEQDZ0kwPhUywiTyTMh9BikhIeDQFbJpOqK/9xCHRmMK92Ky
YEXUDHP186q9CmpyYAEudHxcLReB9rxOM3Zswn3bFb6XvSeVQxOBA2Oh6zkLKQMY
AauhBhqO7rp0v83GME2sv6aZGPqj2tN0IrkU7+P5LRS80xgxXRNNGbY8R/17q9ly
FJ+HzPUw8TirO4J4stVAqlOfpACe977IFLqvAyLrCLIy2nenAhMa2WnMDHlLB5Tq
9Uz7wfrh+JjVOvbk8yOTdmL6kWLYnAjVn3QHVhlvDhvpMENa0jhQSt44UgEX42ET
d0snSCRM2IVSJM+OwMW38uJ4th1Y4M8UkW4V7zy9lPB/UwE2zelj0TYRCbFZC7Me
qjVIQCXSNGeoKb2utYxNdiOOkNPyeLIj1k3WSH1bZh1x2h3PJbqI6odKn6R502R+
moQPqwjUTAQtGrK+Qptk4LjiSd/5tCbTD31a7215knb1HDqbvZ03npESJb0Xs1wI
0Ae3Ru82Ot/60jrkfQBrvOW5JJRSQvHBAEhRI1DvIQh1KCZeKU68zfhlT0WgEsbd
DTRHNdwM9aPKqJTuAwzx7DZLfDRSVki2PQmQxLCXmKIASB+5owZMY7Z5V/gj7NXt
+Z5uItXcV92dVUCFgCS46kIbA+raPpTBd44bFG4PGA4eHcV23yv0Z9HtGVreCc6i
mXkZnUXB27R6xp+PUnxbbpv5LqBCgo/huVgqsYFI30jLGb3DsX7T6ht4B+CNzlLO
AGiOfB3zGcx769seMWmAmDL+VvLw7WXo4IYN3zp2q7S5211t8Ul/f1VVBbSGygve
DOaCjVnySwPPeebt9tfEhHTegnOaqzF25yRmzgZd+mEsHhioXugK3a4ZYHNoEWPx
6rAH1R2zkVEMmNPkBj2s3hCLFTWgtRJzgklBzXjtnWDyaiRVJjEZAxH0VLwrL6ir
ionsJGxapNMWLOdCinniKzVRRPZ0idfBnFE9gNRIvPODurnueSrPCXwg6zlx7XFA
vdA0ObnsU6VF5Dkjb39PNtfdpR+v/BaZ5DF6PQ4NTwQ8aahv+CM1LfWnyRw3fKp9
/kmExEKnFhAkfbhnNWyU/poEdoJZa4T+JkWeV9oScU/tcJ3eXVqBSr/ndvuJtzyS
qdM0dR2CjdYdwxwWrCK0G0Wr6dsK8oB+wnX5Nzu0dkoABdRj4cX+ny6Iof6jp8dt
7TtQa4V4EzDhrlk4tRHU9vkhi5YkShlBo9kGDsYzzx6fOfqtjmTWGBhawzy5Hftr
ao9hYBFldfyC0Nzct4Y2kf88OgZzy5hJE2UcqKPyWxv74EjAC6jzms0rfmKyW72x
7HeTqVX+C3bGrmZWN/F3eC7q6L7G41Yed8G4YQdSItG0TsUoILZUxNaKQRWCrTci
740v8lNrHAhCxy7gprRXK+Q3/zTiwDlqQZN/l5Rgswgn/94gs0sYFzgs2u9Py6PR
wSboDc5lYbCKWvngQ1WPIl7oUOFnFmm50GucVtRwzLUJn4180EZs7G10eW65m+gE
MawL+fNRUiWIQDGGtMaHC4/l619imSdKoh2AAR+Q7WwCaWpArtlMblsXWI4Sp3bO
plYE4ONA0JgsGL5oZOyfxiAUlqPkxYkC/U8CPTp1Diis8Scln3c0MOR1vDPZs4OZ
mKJ58azdCuQhSKHw/bmR846cOwKD/IyIYdlJAnkb187ZiTtMqmSJxxmo08lBsypg
y1GEsQ/tnudoe1DrEfLRSsfhKlxj7b/YcCQANs99MX/UJgCOvt++rhZ45eleDRcx
DF86ajP0PaQpygLG5t2a85OnNtXImF4HreVAVHhaQe7HVqNggKNB+E/yzb4DsU2N
fx9nBhCkqSTyxEQH2pwEmLAV1A+15NvTZ2ff7DKRy7HBmB410EHXPxkgS8DQn4S8
VMKy3FazUmRUbPl0TQWwziG0CtBgm1D9plsMgovhrCJdc9rtfs+yKW5HQYndTfxY
1TaMkENqtJuD9ssjkIKarwQRqERYn0RM2fqrm9r5kE76G/fJEk7pH3LXWcClg/9y
HAIcTyry6xQSqw56wM9ceik/F7s8sYdKWakAwd+5oLvHOhCRwvIoy7msBP/rrWZ7
MY0qp+ReXbMt49dORNPxr6ptLaYAlcrNmO8+f6lLoLCEX/cly7C53OuXu6BguB3e
sc+Ak0CXdfTm3tdpRCFYV1pROfSzmGNucjjKXEaDdi1mGW6yJKsCQoHiifJhDH08
/bXdcwkUZdBa62jNZq+m1o2aYL/hE9AyvA8X2aRCfd6cBo7qa9cNstda2Ht4FF+7
T8+beGmk6h5JAnKeleB/pSXwo5OeXWj/ZaZGZCLhqddS826467PUi5X7402gWMY+
kkFTolWg/w/NYF5FzNMHds5jCi7pWxYrHft+7VgxCoAPY32F5aJckDZqDCSNqcTn
5S2R81qOn4IjWTLh8JRyN06oVNE5G8fBqjKYvuR8q7tP+Co3Tn5GgotH7THJouAn
jmoxdyIiBmfg4LEAZ56Ffmt6kSL2H/yuwv5kVV2ktlPyO702K75v06fwbO3ic2zi
UF4GCJBpgZmBg6P7EBHN1BFWlGbBAFAP0ma/q8uoF0bHyE8nuZIxxpGGjyJ7gndV
NZWQz21Tm8E6kdz2dW1eI6K42EY+nM6kT8KpATlDCDlJVH2AU8ojHQUOrjy0Yjo4
JREJIMOPCDmy6uQfOqULK0AfqZtTFyxEEueXgW72S8JZ/DgqVAwsL/1nJGxnuwNw
n4H4Van8nLLjAESS6HUTdjY+EzweXAwgQP6zJzeYcl5tpj8L3OrZ4DKCYeV14lZo
04vtfIJZmc+w1Gtn+gYPqnZEqB618XhzYa4LLEIu251C4gtfM04P+RWZbwytihPB
5090jik04qf+xuWJ4lMfqQVZsJhodDxBsE2uHPlL7mo4QGgyJlES+UFEgpolvTsh
SultxpFpeJgDxXq6kR9+DLKna5+Kvub5srogiE3dWWmdmYaAdOKNTE3nvXCCfEW1
EnbNgFwGAqhBEZ+2kDP7ob7OftRYkQLmwGN4CW4TXuHRKsBCq2CNTBDjZGO3f5vZ
XteYA+/IbqZeWOsKdPnuFPB9URIVsIl55O9+Vvj5x7woB7F1Uf2Ek2lNxgQrECnw
G6iztc79/7bAbRwDdT7vBXOQ3fgb0ZYEyRP8NKbJ2s+ap2aMbtcffUNRtW9gBRMh
lqA6jNocCmevZ9FJDpgcQv87lgI43c+d1sW4NmvX3eANMl9FB2aLZLn05zt3/nfP
Ayw18mIB/ipdGszcFl9GcE2yvTpBX4ZhrRX5E5KgGPFdibOgT0xRAyhiU/110R8M
mqYbdf/HnvXMooNEgIKfGxD6tYVCqT0GjICnKUWLj7XOuUlMZUKiFXEU3MhP0OIi
2PFD731ykfXNzixYh0ZMSGaU4ixM1sXkoOWNU9G3gZ/2gn8MYkswHVoW2NC2N1wt
sYNErzsBImwsiWcEg0QVPMZYQQfZMTIWICL4oV12niu+usLN/pYKgdhxwdzNo4QJ
ZDXlUxD7OS38Gy9u2m7YfrWxVMC1SdElfzTR6IQOGF6ElxrnxQwsCNr/anN6PwD/
Fs6goE8ca5HQfDWB15ODzVD4SuS4dkTIhJGb1Tj/aKKoU/Lo66EtTNGYOelvoPpa
UXpWM4Acwh7BdAQ2jKVej3CnO9RFy70w7hAVcwirPfy5c+ZmzyQuTTRbYXXBVVbK
TSTpxNe5MQ7RrANxONWyM3HDS2LOi5in8u5wlnfYHMn4/onvQYTfsg6lST3DgTGq
OsnnNffqsjbXD6AKY67PX6BNF/mfCBSVlHoB/WLkxqbtYKWw2KgxXkrYPsnz8qvf
EGfYNb5qBsnXoi1AN7kndHQJDmyWCoDBaukTc6xeJEtVLZMrj52kne7nKhXccnmT
0Zb8lxZdKLnYf7arqScI558BW7ysjQmzIPmTZ2XAfgbsbcbaXpcRyrfPDziIATWi
ZVAeSoBNnfNAteOgJBh6vFAw0zM2KY2t7yob6cWEkzhNLrYLHutQPKosdefMqtR2
ZuQXl8dCiysLpCUMTT+/rjF4Fk01g0oI3uYvXMzRCCIR33JX5hMxaHKrSAaQcQrn
UdJ537fa5M3kDLd8MZq9R89IsJGx5lVZjbntg0GvGHQNoWrpBZgUJCnb2Bl/Q7Vh
V3gUu9boANB+pmdmNPVu6kInnp+EbF5zAjx5ZlJ4YVA3fAdqvVkj9gN3Ttz1Cv4M
HJTSxDCg3bq+zqbIyKEamRZdcwqN3gIkfu8vqzTeZm5HbfBCsNEG0TbrzeKgI43V
QJQFvzhCTsQWzYkH/z2wUgvlOwhY5Crn1Dfax6MCYYNUjTcJWdcSNLKVX+GUYLO9
A3gBFCL/VbUDFm7PixiEvEj3iJjZlwE/00yciHGkrFTWtawWsO4LW97Zagvh/QTo
qMuYfMyQ10zBFPSNjtTTbs/K4R1XkZFAw8No04nywFbXlpH+kdtMjOPjG94YmK9/
IlZweFUJDmvNTyLxzzyLETWJy1JFysjU8foHUd0iRRF6IIGIiiMz0jVGpoQGLdCH
lHCjasL6LNxqitm4N+F4xJtIDH0gCJz0/qu5tK1rf3cHGuIcT55nseyLxBQh3gdm
CO5MRph8Zs+9/ehuH9qo4W6LdTjWd0ewszkGmQc0tx8DoS5TberuxdiBFcdC2PRw
gwHF1na5b/5ALBnpbvc+N1FrhZK0d+ZvTOiJ5p4VhV9L3ZGkZeM68kdyz6ADup58
TjzyACkW3y7rwK+jArLLJYRFuBth77p/mT36BsnW9UTHd0Mmi6m6YAyLzZRGVH05
FL+DRCXUa3rcwaW9An6Yw4jpoRZkhjGSG+7xr9+2mCzLcQiC7ubuN0QWGw8roaWV
4OcWTy/+bNvNrIZPxO4rRGCiyT2PnzKEj375j9kpZCgQQnYCPJqhRIkk2s+yRwyk
zkncTWnXXBoYVkwbRElMlqDSxbpo/I462JklatHARqNwu4Seyw/MvmF5JEEwE3sR
sV6wz3UgHnRtc+rTFpdIUNZqQ233myzxDBgkR7vnJ0Z3Bdsgf6K3s5p8DEvuPK5d
kNn0pXqHUJ2SBo2kwwfdUOZpWaLBW/hH5Q7BTxVSyC9VWclP8XaoK9Xndgy6ETxN
C+zVfoT/BhtCh3pIpSmcvDcwnVBqYzd4sPqq30ze5olru8GgHv+9MsEfGzhBAAQw
x0lyHg9dLeDM1ElYQ8AH2ERB0cs+tvpw5dnZMz/3hdK6a//+s8hDADEcjrhZDI17
fBfKUTNRsxgOBnCGOO3Z1fsEq1rCQVH/cAgGt0yKviJ64pGpjdhLQjj8awkIUnN3
xGtgDZGjpLG29cAaopLP+Qwjftql+XOHvflGTKebPOm1bfoZ4z4+VLTIHpu97lOl
LBkz9EfSO91TqC009kqhm2Aach1Bcx0nScGdWz7FtrKUJFhnURvCuOcKsuBeTy9y
ZpdIKQbl7Q6DsWIHzuPzA4Q9QI7m1UfpsFv85vk0mfSJhEc8i7+Gx/r52wXdsDVC
fYM+X1ichx8zYhrk0BkahrPE0pndVawRcru0us28TdsSzRnLeegLNWG8y+LK5pHD
2zglPno7b4c7gM2pE0Llhl6YNmtVe2MFZL5IE01+kAPANNyuDMtb2uQ1zKEEkUf1
AdJRisn45yWZHxO3rYS4+7hihCVlenaedRLUyAEbxmfQEbOp4C7mnoy0JK6kT6US
N9n2VlNdcyuAOTbKDlzrqQJmfRiGVU7aGWsmxAXVjD/4HEMdQ6VbRuzfW522MfCE
zzZ83S6vSV2yrD6E5808kOiSu25ea/l/bK2fYa8JeWXuDu/vJzEaopyLeGbqJavd
6x+xlzd61xyJBguLpkQE2TiHnK6sDcnOArbvU+tcaA6xSpemQNSXTpYNagvYjtwR
`protect END_PROTECTED
