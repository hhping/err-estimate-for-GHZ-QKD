`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wx02hnIVrd1LesIJWqk0t+larj92kGJNQ4C2AgIuYUEQYIocPjGMHTxpx+gvork7
hdG86kMjDQb4KFRqihRhCbJjwaar0mpBKjLaS+e3lVaG5AD+KM5mKD1B2IxoxkWC
2dsX1ElWoJ5pKXe+8OiIDbjGeBk4VJH/79mv5QABWr5P0KEqtSr505sjljZpabLK
81zdYVf3+479Xq91SNoQ6M8o22W9ZHN0a77nWrN/a2ng6yzeKAv0gZrk2icbzhLY
AFbja/l1UBbEXOuI3gahLTMO6wHzLTDtjCyC+N9eROC7qmN9uGxkWpYsC/rZUbzv
VJblmCBM7Q+ho1BHDfZvVQ==
`protect END_PROTECTED
