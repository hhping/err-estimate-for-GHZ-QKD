`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5HEZRCRocUB6odUe77wEpzGL233DhPn0BfR16IPNSWNbJorVddvTr0gBKaRO5ols
MoGnTP/31Yf7XPuSkCZXR8Yc0eK7I9wn6aR12FYglbXIjIZ0fPzC+FeCqQhwJ6Hs
J1BLEGcJjn+hwzfihNUCknSWosnE9fGC1EZVomYAtfMpSPXexVMdQIPfQ59ua4SP
COi4FXRtPUwXiGVh2NmwWI4M1QtTsWYI4cploTp2zYKilsfz7Af4PIbVkFC59aR7
G7MaTGR+nibz15QRQ/P/N1TuJjbIvAJl3dHaVYjpPBLBiXiBgo8Au1TuovHZAhc9
TlMGk57dighjkktli7jAUQhZLuQC+DK52X1+g9PdPt/RLX1NjYwLnIZf06Ddu2Mi
Zr3wNzvUkI2qG8B1xc+KswBbrc/OuDe7CpRXHs61Uf/qkZUzX+BKeEod3WAiTPvY
JCiTchMvaHxFd8RHXCrCrhZTSW4IQjMGY6NHLb7977UnRNUq8d0gzWOxqfguOkLj
XVje3SBemsv2a+t0iDzyfULM5IqROGNFt99iDR+HbTaBgdH9eaA1aLlGJH2s8j95
H6hUW4FJI2ZpsaWCuSWssFOVcEfRSA0pNIWbJX1JRsD6W4pprDrcgErWGjcpj1BE
z4An2vm7khjlUykPXEr9RfqCbVCCr8sKVe6TvvF4Hq5vIAQZzOosacnudiMryuvD
XMDAEmZtr14118Bg67U0m5mv+9AZff2ovumMnPM5+XDHbeRxM/yXvA8nvM+WjvUi
8P/Gzt9mytIKpVCpiVvHsyByqwIPkOJ2k6lwoD3wlvbZ4G68tAnbwMMxI6SZV2YA
sXisv5OOnU/+3PSStvtNPZh1QzMERzJc/A61DBg3KRLF3FzNxZ6VLofIWHAmT+Wd
ZMJMDGvjbrDjBNzEf49BWdGsaFJBizKM1xRVQ9Q7/gtswbcq2xLyuM6PJn2bVTAK
FsLh2lSIrA3YNev/pghBKvXWTC88c+Q++3hLTOg+pxon1aOrcUTsJopODPRdBHT5
1ZJXr0Df8Bujjvd66NLyBGou93tl/ffY271BZufc48faUer9QkwNF8Ji/udr9WMX
CEtCQnAGtDTUXqP9TRmq8LHjR9W4h2DOfuH6dQl3+wDbYMG78mKoxgkh4/DUbcgG
xXNSlGMExJDbXMOZipCWy3SxBXtuK/V9eJ2hkT3MORgeGYJacdfhI4UBG7Ho5/J3
kNA8Nmj/dEhF+zS8xCYRtknS4X/ERlvoTgunoBz92mpnxaAMXEyWKZEXOf/k8N6p
fGV1bOvmc6ESUH9S2qubQzZgWQwO9DlAR71FWfFs2p8r0JzPlMxM02AYOmCUbPXy
Al4BWyMNoivNvUE3n6rlYJVb4iFxVM2Wu398TJgOsMmjHXTFl6HS2MtOzxZ1h9BE
q5mgAdj3kW/bgHCg4h4ALDOdszU9VwflqjVtnR9E8AqYgZV79E++tkqfa97V+/b6
nJYNLn9b4vovjev8mV/bmk7bwR/qumzKb9S/1Pfsw9Zh5NRP0CS1oAxtZJlzIG8N
a9GyyzWC+5t5Ef/pRudox2dym9IC+qWcZkNEEqAdTwK6cHNgiCz+OhTxgdMpUwmS
4oHiuK7kzQQNRUP9g4Yrje9/toPbb4kBIZwWnrnFcEpw4IuogQvD7XfYlm7eelLy
`protect END_PROTECTED
