`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r5IxE6OM7h8xxki4qJ6wtGBMahx3uppTm4Lk6pQnIvew2f94ugsZxvTOfW5uAGhn
CF3M74icSqn6JnEf0du1ATxVjHY4FM2xUxLdzfOBSYv/8SAZtAfGHlSSuo20PEdd
SFSweEE5CwGMVP1lyjfn+/dlnEH3NANMgA6WWb/w/oeAE98tJm6FiSMf9HPAvPgq
KhVye6+pj9TVZtRCT0Mvj7/LhkcwK0bV+bsaceAPpL1qX6OUr85QSKNDpghqq1CC
bRnCZIE6O+8KytnvtdG2AxDtEEgyQjHiTgg0GVMv88YiQyHfZfHN7M1TdSj1Q5OL
vFFnoTmcdjZQpU6kWJ5GC5mzh4thYKKd2LMu20MUM6yO694zP6nA9vYUZrBY+5t0
j/u0rpyteAQmwlzfN8uspRUNFfOsQNgAAYGkRtO31qBa6/dPKLPtcTaRVs57d533
0A+t97RTJjATUY2LNUHgOkDqUsJk26jNMCzdFmB7QiZDqDuuXyICTQCzfP6d6rgm
Jjp7Bks3CNGDyqhzlPYh7K4al7wR2q6QEMTGEgsm7OhlmHl2R2yyxMApEFxuvXxP
AsZKwNLEBpCD4xHvWBLMBsbjTKCGVze5ebn2TcnrU9LEffKFi9/MYCVqJscPtiZ2
GqOPzc+Zvj/21UImfmQWK/uaZXYCuMjjTWKBEgJGoGVlfO2ncYmFEByAUJiaM94M
SROZboCpFE8r99KBTh3X5W30Zq/FDhJvY43c+kDDERPhkXAyTdqQQcR1zjE7LPDK
SEBByT2QoqXwvr3P4LZqG4wWKi/Jx9T8GEynE2sxrQ9v85y/Y2WeIkI24zWhZRuQ
9tI+mevX/QKZKoB42EfUYHPnWNLIr8KIu30EY8MrpSgm+Y6+jxMphUxGwSr7tkoG
MoDoiFhlS0QmIOrUVxnzSuBRMW+P+htQHKLHNPqNsE3cBtcjQIrPhSRPI/xMusAU
m77oeLrQUZilgAKylJZ5/YeLSk30HtnDdv342x7ubN0bbQrVvrXZPygYXYo/xMV4
CAlbe2Knc1+hUXnRGlj1WJKB+puxEntz0HV6gkAbOVE=
`protect END_PROTECTED
