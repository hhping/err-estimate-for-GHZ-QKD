`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
riTC5rXg7m3fnMo3NNQNMUBulyIYidaO8HeR+ny9/Z0igoDCUrcExWuQimfbdNXK
uAmX+Bj13RQpyDhhHZYUx9N+uF9v9bF2wSdumOcZduvCc0U527jWi8HH+3M4Fm3O
OUMAJHZ5Reb8i10TIw2e7uUR8CBtlPdWouBkWso7rjxbBKTzBennav1hhBs7FGD1
glrTOPqClw06wG/Vyuzz7++Xpp/2lktxYQW6bQujGRP8/b4AV7AvYGkSjqI87HDq
SXs7Eeq0jAZ2UCIIndg08pMqN4p951HN/lwutguz/BsT2MlFnQIGVvNVM9/LoLTC
t9fbnW7a0fRjJ7Sc5Sx19gEBAGqwf2STlY/FEUW+3wGw/B63qkjRJpZ6etYg33U2
W3h+hF5M37Oo3HaljLvfj8JQEkpHUec5hwuVVcCjQiI8aHUZtSCaccpUNMAm7opt
6xGEtQmSJGMhnPd615+PzBrD+OsKp8ZZUkgQAjorfX+6Urc0JZu9WvUQQ0qtXVSb
5wrFN7+BfbVAPY8hQZfah5kCKezn/1wuoi1jr6J8ZbcyzUagIPTQmf+umKxjb+Py
UDRgpHFy0WGibGDyDBBG4vJOqF3ltcLnb51kJLgAm1e9J6NnQVZKHkeTlMLMCMIJ
kBlj1RpTPAleTcwLHo8AIfExcB673oklrmRGVoTjhJQCWDmbq9aeBshLnL0YhEdo
m2AbyUAIsYmOm0ZaZFeZg1YJYM9saJFEKVUVZZPGBwTnsKevpukUq+IlqlAWPwhj
RvNxhVVeAaJ7AZwTrGNJiw==
`protect END_PROTECTED
