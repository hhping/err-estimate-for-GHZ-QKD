`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
53F2/CpgUzDIFWhW+MLN+D4esHAK67iwxQ6sCOTJejnNhhWjIAeIwKR1JilSh7ev
IrjMMBZtq80y+RdN0kgkaWV7dfCoicg+HmeUdOiONBX7K15IZBy7YVKQOK/PR0TE
T3SbVQ5Fe1O4Qp21JlOPR3yf6TauASRNz1440clRr8nFjHyf+j9Q5mfmcX3rcsPE
itSKES+LvXICb9n/5mZqA0AjcYlqNkcALckwrjGnmkcqA6g795UdwM0I75OgIayT
Rs2pqaS+nwaHQAoLmtUcpCaBcDkdH+VOg4safFAAuJ8jAoXHaJcrnAAu47ZEprsp
FKqc/bvppEmGgVt4DgxAz7Ts5I3gA4qWWks4uY6ui5CkDxYQ+GIObzKoGnM89mpV
HUgH6cIW5nSLQTpJsCJBS1GkpF6LEtvY0PdlThLffF0/i10Vsr/Q1eJ/+/uwlv7Z
ONrlCrvt0aFrBMjUafLVwRh0HItVCyxD1VOD58ljYfCSB12RM7Ce5OcAtzOdVif0
fbkn10FU+srtoWQLBqWOv2ydLyRQOxbado7R5r7duOUyF5PYEpr0w82iECEf1qYE
vuE5g3l32s+3z7DsgC4tcjF+rzx/Connfr0Plz1Oy+L2i4/YNXHJG7xgLMxjNsT/
XvUiQeSCMj3x8w0CrlK0iQ2VSAeUgfFq8t69QyGexUs7CMzhSXT9L2o/rAtG4Ch4
O9ASwlNIClfKKbgSMo1/f38frP3Uq76BXXchJJf4gzlqhXV19Six1kAro2c/AFy1
17A5HlGrftvyjJ3JX4/ZOutWh1T37lmd6EmJxkycyT4qRAmcBOwPqsc5Xu+hP49g
0GrQw+XIc4aIfLW4N9mJ2h0nGfUmEX9uWql20rghIlXKfkQ6YiyFswRiYLm9WYoJ
MNsrWesZcctkV3SAaXTDBFtuucGJ5NLb8EhbA0ux2EA9onuzU9pLCWxSMQbCEX9y
enrkurEnGoPo+ou3cfELqTSya9K0TC4BCBi27BezOGpwmZzErbgGOS6125qGj2gt
cvCc1EVczhoJgrfvy9E0PzqtPEIMgavpVxectfV+5+nkKjKiKsEr1sF1JgyNcKi7
xk5sokKmTfDgRdR7i1dZJZ24reebqnWFWWwq0hJKT4Y3e82kx5PIdPdnaKIvXY5k
2eQThfyDTkaFRR25Xqbkh1PxhUtgnQMgv6HUGhdSEzAtvpEJUWKdqw4mkGj2mKih
wK/O4svX8DBh9aew/xj1uMNYoP4tU6Wmz//QijYhLVN73WNQbx9ySC3sIuCKa7tN
rZ2L/W2fkzl6HmiBkGkB3W2MX6ksIC+3gOiGsOEk5R4Hq6D/gzU1LsMb3yxzNvtT
NVuHK0gTYrg8+vTkbj5zXw==
`protect END_PROTECTED
