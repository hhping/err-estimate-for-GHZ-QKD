`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
811VpAvoosc/CRGTLQuMoa5yeirsJ5o5mgkOdX8O0HQMl1yEwA12YiY1RhtxTnFj
0sl0Pq/y/ovFMDW7MOc5VZhNCUBwClaXJ05tIOh1JS/eeXkQT+D9//8CSaaowvOc
pHCeHuErIgykHKWpCBWl63Nv3lsr/+bQ3CjhIzjy6pIji2C/TBweUpt1rkSI6pBz
ID65vFitQIPX9P2ds/YPJ/FRN0bGtJIi2KwkN3UZ0gwY3cvGhQygQgr0Im22wlse
HftruCtipapE63ValkY4fiXikam4lEyyGS76fJk7MqHSbXJ54zExPSkHK4iBicnh
2Iugq7E68W7SJkAI+JVneeEMx8qoZow34gBE+aqnCtpYhtSeg6dbWbLVaCzSdI56
KUJ4u0AALwunSOpx54QX+iUOOqE3xVhk2hQClaAl+79Mkm09TuF+OB4bv6IpI5pX
DSNab6B40W+il2V4mmLZwifVdhx453+engKl/k3TdP7/k/PR/7qkmyYkDW/W+5/Z
hvk9CQZTKqjrt/8SHmPMF7Dij7MsFBLSuyVrNTC1YYTkPSk+7OfOAVVQa+ceQJ7N
g0/OihQ194kzU3OE/XeK6cSLmnaMGN3z8QfGAQnCj8hjnyC7mlu++8vmrdZR2nxy
/I73RESgccZq1lomHtvKCEe3RaCOPiH0/duXF1d8VeCDDrnGcumVhOgaEgaH75WC
RIoNoAzYiPANuUCFS9ivAfhi6XCM8CXJ5UrS/Gan5njQOdGzZzzuFYZeLOfAnR4R
ZsfSI2PH2FD60X6U4c5TyK85jlltxbAiwATh8FjeJH+BLE7tmLMIWkaINjSZLXPi
sUq1ckM9+bw3YDj1oPtQ6M7J2dl+D/oq6lFmbphshsLiU+ma2pF9scj9cYMeFuv5
4nbs3dUvIyH+0lMkwYfYa9KEFcVWxXT06fr+7iIsHwhNwApx3y27qSfEx+rLifD1
9V+9eUcivxeevc1A9pMJecjf8H9yDJ0ZTDHwk1nfGmSLbY6BMVbUYgTI8JNsaD4I
FGw3jRNanniN4bxqhzHgM5cQGnnDx5VDvbjOVMJ3FpiYi+uR4TExhYa2/trxFEH5
CqGOkusPEOup7ty/0bKralia1lJ49JD/Ubr4HzReQDr54uVEFCOsf53+D7zbBh+I
UNjA3A44rQeG34aO/jlyzA+xFv+GRQNve+lKYQQBSbbqnR03AorQ+dcNPopy+EaK
jdy+Ra07cWzNbz9EYfiP3Gfwzb1XkpU4N6U9BEWKjS0Lm9YePMFxv9py8eWv/46i
58w8eQSxhWG4kS67zZY47GLU/MCCI6qGQJXgksHehqqMir8Je+n+fBl7QzjcZ1WP
OD0/Mg5ivE6sN2TY8jUEIK24ojLxK2Y0AU9ivWssMeIGZA/coqBLOO2mscoV2blW
OSrZexMiNC2LiO9wYoIIkHas2x0w+7cwFxD/7DLEyigzdwbBPN/3Za8+j6pRyOCu
UuPzQV0eWBYqw7neBkp5k0b19K/y8/4gkNZH3ynV7lXuYSZ4ZgQ2ouaNOBa3UexT
AuhreeBpqb3T83BNhQHJDhz+G0bPIsUevCDcpJ6RYsU+s/wbWQhbsLoGqBDCB5G4
pL69J+LXIyw73j7Vok+XYHvDWXFHBpehxgMNTIIYByGQ8UZrSyeq8CtGoqeL03eU
GTMhXgbgMlqEYAqLwd8wBlRXra2oKCiZyOHmTh3XR1wkPsYlvXPvwVnRx9ev6Vsh
Xqx4zDOvv2SLsp8Zcv1z0iVnojSzid6WhBFq0KwwsPfxihJqMIDtNhVShori4ZS7
99y+9HoMZMDwQN9M1XV+aDOFGr5cD5gEpIn14DLWuDK5ADujHjlGYmyYGpT4C/nc
H/p9jVzD7KnIR1n7T9HdDZRL7vSgaEX6U45qIB3taJpPaxByO9kpjr/T7AbUrl/N
TjAPb4Iy7tris58bnJS4yUzgWLxVJLEzG9feZ3vLYQQZwNogU0tEvxcxG0hXnPb2
VNnKh6Ao6EkUkMHk/u2l/bncbZ7L8djR5GQn0Iz5RXRfpHXoaGsbUJwNZfF61Wxm
RR++RwJ2LzqNJ4I44/2kDT8dE5gw2XBJ7w1wsDlQ5Xjre+P825aytXCUxars5jxG
ehVS2dw3eI9SPur27jfLYstM59bqfPJrx5XAzB6IsNKFTNUubHXRXaPtLWvgNA3F
6SHxYVDezSIn2N3vRrJU0wCEoPVLGFpuwfvZW6HbtXd+Rkjl8xTx723wfGWbJ05Y
9Ot7BiQr37FTL3FzPULk6Sotci0p9tcVgAyqnf0BFfiQOCWKuqEpXl8hNRsWCIGH
u54UdimFoz21riE5Y3SYa1INCm4mLWvaAyeDENZ2PM7+UypOIGA1SDmkokL8dInG
p1wd8x0S/LBsULVZBWoMyBPmoKMUKvrqvIiYkILpKWTrhHbJrZ+50rAx8iS+K/zg
xWxaIVtLyjTzXgc6ZZmke3N2yeNDsSV8nsQIPczzThmC0DEsdqeRMqLeH4x3PlU8
iWdCGh07rVPc0QQit1gYfYyCRu5cESPl8Vq6ifQsfUd6ag4WZgEYiuaMbj+PCJ2u
PW4psnOR6939hgmsXqnom/epwyi/fqEtFZKsSUj+mnWQ5ORso/HstliI0TmePo00
Hh33o+G+IZvQBXDPUGVsC8njn5rK+rZyL8gpF4NqUGumhFa6H/TlVI2yL8pHI2TR
O/3irZNT0sBWkLgmRjLy5UHqsKfWTHGQzi3JNkPY2qbw7ZPEXzgoKKWkGyQO8pqv
Y1Hj60pTboV/cRv+vymg9GqQZYODJX+Hv0Dv2pM8DmMiJloRcdw3Iam+jNCef/A2
mipcxrEx0SoM/oh3qshR4LJ10XxmoB/WhZOTSwIvy+4I8AD34LgQXltJ29fZm6zx
HXKAEAQKPc6EtDWyU4OxpgUtrjY179NWZKENH0aLIYG5lTSDBd5nsuZP7cePxdM2
RL/CXp8+OnWIS9M2SO8HuMMMZSE6F0jKqVfqDOl9s3oL2sxLiciLW4sPAMVSOs/R
mMhDMZdYokSHlQI5CWhlabGDeAjR/TDNAngZCS79j/mq0lmeWpXadCzFRAxRZmBG
ITeubeB0oCbIcl8P7IWwDk6FjNpU8HwtIOxbk34nUn+8AfYgGHktW+g44FB8s4xw
iBwYd7Q3qH6p0Eew4muaoRoDT4k8jMKathDOrBclZ0VYeoX17twd0ch4FWlNKEBn
8dmDIXm8+WQnD1n1/spolwaSP2Fbp+31kqaFgDW87rF0tIwCEtdb7iPMnahdPXim
TFZmx7ApeoDiGrzz7Q8NFOgu7XvQOOhPH1r697sIG7DPuf3eZOcmT1OTslGSd3HJ
ZJO/OYtVhCSpSwupSWptxxcWKjkiQL6bK0MoQnI44f9dTi5xpNfkJcptf9vPjUNq
KUGb5V4hQHckWQ/oEfg/+0+cpy78aCn59BpSHv7GNmrqaUMtGje4KGDXDWsEWEFV
`protect END_PROTECTED
