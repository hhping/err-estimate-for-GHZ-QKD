`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p//H5Urlvu1QewSYNb+SnDAIACssVD/WjmP8VkHcgy7qH7+bWJsJfE8cZsPwW7Jr
BaQ/EUxbRYehRdiqbqyCHXZxIDZGAdhOJKOUXjiOKTO2SfVJ9AeiTKeEzuIXMsw1
G2cC9xSPCuhgl9rPvCwwjUcVY5yROxmvlkt5+wSSbIUBoyo3WfJKk9Irre9+sb3S
bKx7Ug7DeTo8Y5fFW82vlk2vc5yPnapeJVKtrjwvp2QjvLIBPYax8VDKjMRlxZIG
1Tm/fyije6DMy2Y4ioEJ8aTCpxqeADY1Hi1aZ9ePsYidNzLrxYY5uq/ENwkjN2OG
Q7accjsSE/h7uDblZydIVSJpPH1QBYorF/esLbZkA6Souf+2KdNVnKxiPeUeDK0m
kRs+SUtv5+HyStjwIO9ajmbsgZfOCIA/QG8QweKI/P5ZRBY4GEUdSeimxv8hNFEN
ZvJXC697nzw/6QTlCUqRAZmfXV4U/MU2zHS+UXTIybqTmQqDGH8/dTooj+8sAjhA
vfgQ1rcolpDekd3321StENaYAXJCNx6b4wHHa7ViZ/eIeKLN+ctoQiGJV7hVEDBC
2qcT6BHw42aPT98kAvdYCGZpcjqYFUmsvn9WHIF+5ep5U9Acq38vaiAFabJmGHLJ
6GDapsnt3NoneFjIEuF8lF+WRoEZ1lJlx2vipnxB0Cjegv8tMqm4FlmlovlIlQig
Smu1MEYGTmFhAK886l6PoWa4mLR0UDifpWGkEDjHnDck0lFbV0QWacNVbJHuBvjR
kIMoaLdTHqaPsugPnAONSoGHHPnQgPAibG0LN66h5IHQue4lrhaxWwPdSaZck3Q/
nC/gjmptkbZ2p1JxYoWxj9cqSQ6ZGIe4p2VlFWzgm0G6G7erORqPCVW1mzf1Ez1p
ufJkYV4b1xvV3PanRATfl7IImhoTYmiuH87s7zlWC/KXhzcajAmAx5hsWbiPTsmw
CQCnxLBHT2G9DlnzwaCMrgU66pCoBQFXMMh7zhNB7mE5NDMl6R3xPwlyuhndHVYf
NLR2mjPS6zonouXY6xdDsvfnSabji6Z9h0IfmZtBPMGs6MRd72pP+RGU/YarqWWq
vzNJd/VGZhIoPGdF3gMyxLiDy+w03L7At/PPt7UA7ejqRfy3h9QVR5X+aFRvq0HQ
gPy9RE+IV2BPIaUh0JWD01he3pCuAzcBb7XpoLAq9f0tnThvfAZ8CEDC3maEVeOk
GBd+ggCX27tSLzXMOMPzNdIQDtsG403fzAWJwM/EDymGAK+zJ5erNZyXOoNRp1ZY
2SG4Yz6lBZjZWvY1nByblBsvAHw2I5IeQqdyq219NGYEd2z5j9gKkhCWXlD5o0bU
wsLBa5K1oxMK7oScl5h29amWVQ4foJZ5IZFDx6BzT5II9s+exCLXj0qsnGMTxlBA
fQKgK7tRkiD45/UVbBsOkpqJ6Tx6QjDugUIFSSTN6rk7IKkqBPHMpp0hQWNtT1AU
F6Lss8POmLo8ywQ6bvgLo39IumV3MIyMk6tihgo2OTu4b8WBsMcfaniepbn2bCEo
Jul/B3dKnRZ5PuHNaeULFO4e7UzuGcISx7r1tG0rmpvXuxAR1XYt+tzjdMsFJci6
w14FzvRyvexUAlxvEJ70Mw6sE3ZLP9jKT31EVThO/fvKMP3svU2WFt6RLoeVwuzK
LW8ggjfM091qWXegraP0CSbalbDb7X/J88sldXtrCw6G9jMfmVx/Sr+NTTp82nHN
hLCVdDSr8uC6KOlvq4/ufB1rMr7csp17g6wDsjw8wV2b+4b51ZfelgqiAl0HrYxK
hZltELAqPCe5iz2Y7eMgFdp33j+w0/bxK7rYyKaE4Ip48ZSAIj1dy9+y4JXFpVXn
ltPNM12L0+Jz8q9XvB6YsrK+J7lbuzNdxfg53wBe/jFWAIZcSwHnTtImWSQnPQLH
JE6dyFb0/P3X2qTGBT6wa3PyBxuLe6U8JMlAOvzH94Y52SR6642BUKyAI0lnMbeV
vH2bp4aSG94KZYGFT0D45g/7Sgr/MxiAI5DLRV5M5VlI2erTwLMdmCbHd9bgCQIY
rXSI65TBDmXhCMV1hiC8lPVc1veYoGTTJUEcLAy3FSEW2iEvOIm0g+k2sw6xs+K8
BeQyfi0G4caOlKwQP7CYZjPvQG5eRZ26BwxtiohTNzDjQDFiLWVkQij389ggJKwY
2mJOBjOrn9d8O42gy4G3eN2dIgRR375+8SxsWTZl834oG8mYi/vccVopKnpMkrjD
gOmp3FldRsdIDsaWAWGwh7M83DTXB0WCxs0JZDfILLYzvXbwvO7NIPZeaNwF/9JC
VSXgk7Z0CYaLFKZVM8LpEGZtlBNF1npcTXsFuqS61ndu+CrSCnqCe/qWJG6Kb3ro
6TDL63PJn4M3JRsf8ZE9bTwiPlzLH5YLQozcGjUxjWhsnOmUHn4AiOXiUX6W/46E
sxBZXb9X8Y3tpX8NQaVMyLA8jRMTrkHBkPFrnDK+oeagIQWyunHAHtdpVbGMqMwP
eXk6LmEjoTXijNbXrPCmNkok9e+Vw8XUU86NERGqMXjIVnX+O+2nYtkLLtT713KM
CYqmai0CEmQZY7BUJHn8VkjwU+XybiOGkwYRWD+9bfBsfo/Lrl9zZ+TKEoKp91Ve
I/ooF9OPCgDcxpxEFK+NH2iX23dTzgk82xty9SeKwCOIuu6sUEb67Qo/EGfTYPvu
5jrBt7VccOG6JQ5UxvM4RVGSMS8gAX7kb9a3UXtoT/mddKTV7Q9dpfPGEGIFzQ3m
qw1uj0ngwptAtApOu816eRHLsOQcZu5U8eG/jwxAWN2zQT4IpcXV9yH5oOhcAG7O
p/USDtDCj1tYUHi8HN8BDGM8KUFOZmKRHehMcavQaeKzlQvTLi6ohnnxQ38npzd7
yI39kYNXA2mOnAzFKFQWhWvHnT5sW5wYAAj/8dl2FcmneBLaIUnsuD92YWUyUKrr
kc2NDKFIRCkD3DO93Qi8WyTdJftSwVYcroW7/prXs5VD7Pc6bpQzlyowZE5C/Df1
UCv47Zz4HTCmifOasIcApN9LugSNtlYZR0Tf6CkWteHkmmlufYkBUXS27szHN1jY
yXYhUwGCxtOr3W3rjeWXHgO+95fJNjplKlI37IHw2lUo9UB48VSjzjVbngkWEvUl
GM49iZIcft2JafEaX48LCSmW/PKHKvt98/s8Hoqrb8MxPr4mvWDkb/xEQ6bZJaxZ
AcLWtb+geqNyR7CDpEuwFOOJ20v7WPt8kdHekXO92CiUQKc3yGYYZygN9z8rh3kf
2e+3Yq8YIiWFK1avY7uRiLtl7YgFlHe+W9OnjGaDAoEQTyNNN1TyINVvCsE1rEBg
tq7HWc8MjL4VIUym+LVSNGsWdeIIB49UOXXzt0DNgN/n1DgZgsVcufTXzv1ARY5t
4TG2kfQAog8oJEEEmxSmTeP3W1zAig7mpN/VUVYRxGHbfHxW6Y8eOGSqdzUpjrTw
IvgmunKtbOYicC0o2cciOc4upr7mV09z5EywJ+ybii8tazWUyKCBG6Y/TZw8WyMw
IyQ4nUsWXevsnwje2ZvdAhujvC5Aqfw0/Ah0l1xbnxawpLL+t5qSnqaTNubVCs2g
UBNaW1Y3cO97QcxQaUH78gIHlmtjtDKdTrotLWY+9UpZNjUmGskeYf5LlecX7efS
TzlndmVJAuQ76UFFawcPklCfoHd+/14FH7NwbgmYvmBIuT7RiZ6txuYKKNkAYPWm
SpmCdBR/RYGOnBPVWK6fmvhhn6Xvi6kIQnwyuNM0h8LpsJAp+MvEpgiFLjVB3EiQ
hgk045/sETXQkEjRk351NKQoR5rT72/SFW9+z2t+0T8n3i0EBGNz3d76sm7lKZDs
2lMQxFdqmEJHd2dmCxpzvN2O+2nP8jWAosR/BuXG83Q8oZXEwIB9RxFDeUdvL+YH
Y9YXTZySew2Vteyl29xRl1cdOwbryebqzcaNpA+dFmgmEoaTOSm22hE+viK4DsgX
s5XI0wDb3dQUsWy3DC5OnxyIluhLFcz0vxXdOKx9/otOliBeWsYOA0hvgEJ8CJfh
7R+UuYW0ciHLBSXqTtgBf/3Dd7evLGzZ52FQ1NqgFyCJsxrGlXyUlZkz6Ol25H9b
KR1ElqJucO+VbMXBAZtaMSIV3Cd1cI8v2H3ngjdmJKcP2/OF/MYI42SCho9pYRBG
4MhjPZo4fahJDLJ2LhwknQSry0L3pc65MdialaUtG5EXUAfCZhbXs1q/FT30NZgR
sCfhN7e2nbB/XZkR2yp7KjQuoh2kr9nTJ1ivSLf54EvjDrvvWBs6braZcb/6dxoO
1xLXeOc3U/UngqFl0JC2vA+801UqWlxp0pAEcJcUpXMQeqwQE1eMxvX2v1XHvk3B
iKrxrcxbFohOT/WijrlJ7pltU/GkkD+MSCjLWfqojOywjbbtLf4K3ICANEuasmcl
92lnueeaiuVikdP26jLZn1yNl0p2V9yBm1UktpKfFMlLb8JvVXbXH25k/4lEU9+W
HKttB+O5ORAlSuEcnPT3QgwJIgcnxqtnvqX9SWa2KsgiBYaZ2dohpCVMYxa5rps7
sz/imn8k9MN9Wxov8+WqYfXGRXIktcnqu69WFXRf3vLHeeOZyC+XGrKTkyveVVD0
Btt/JRuUgGEQNw6KLrqQWCRGflVVsG9MSvk6T2jS6mtGXw6Iyctj972cXCxQXmZZ
HkGtXq9wsGvQWZfxjsOG5OIajs5vEPN5SfMibJ12190Sde0G+pcQSyxnB/OYDR7+
dVrlyQS97EHG/pbulxCu2OUes1R/0lCLAs0/0AmW0TEgflWlxXqmLUPkhjpVKq77
wh4kZ3sJXvqy6321iQe/ikKfK3chixafLDJe5ujm9pIUdjpgQgGifUqkLX8gfgfK
IGz/6gBF9ObhZEmppF+XitsvQjhl3qnuRWJDsoSn0iXIBMSuGx7fcccUwqt6/TnU
xckA2oBhj5s3HG/LKibo8dvYP///8JEvEELZLEBL3seKpCouocS4Kd0Nbx57G3ZB
yTBwexFdPPK7sXj+a9Qg+Xkexm5E3ExEvRug12AGnwhexbElLrYw9WKoMcdwxvpS
SUgVoHkeW1Sh61Eu112t3DKEIC1yq+WXQAZ2NjgOHYuaj2klIr73DmiyVPvu+O0E
gfSQXaawwrtgHsMwAlWgMgb3C/B/y59nFxlTa/7lL3ISe9xd/a27xKws72Td2pbM
0zWhSj2PP6lx1lDUvixAit0eHHOIhS4Bb2N6Z82Wb2g4Nu4PDPmQODn3DY7NJes+
POMwnVxmilffGA/ppGeVOtGPyLd6Qf6xVvb0VAR66hHza+r/SsimVrQglYO1feGD
6rbPfM8c5+xTidZCZhrVuEl0B1eRPDntdm5yQ3w5KFDz94ymDZ9wK4Sj0N0jX2Hb
ZlEnIlMqMqGCcYDainKb3VNkB8afbG/DQPfjDuwjpgQxDDKakDGC196+R8qjw1PJ
JKWIOTKoE1+rece2zeDkb27PywyiDvsQc7clGVAUgFYymhxQ+YpM8tFbdoqLDWQa
wU/W8O8t09QNG0/lvOOpA0C/TkoW3OQAuFejLMUQRBEsrTYT//MpVXlgUdQZ9uwI
fZQkQrMvAFVMAufR96AA12oANXEbQzeFLyCTgIMhCwFFpaOSRPYOt//9KnhoZt1d
opl8v3flKNWhz6Tm+8CFiL89w6FTcZNAXEHt89cBgX0a13uIs0YsxAZ+0g7Wcs73
14ifeLG/mYDZz5Wt5qmUNuxLIXtSuHdcfFzkffxG60cCJrEvkEchrgmH+5H9V2Y9
QNi4lU8i7h/HBOJT7EZGHyFT8vYa0KIRVJtlnuB+WAs6fvKKL7pnzDA+iXFOcNgr
q56nauKP+W586eWH0eRA6/BU+0zIrbmXbGiEHHcy+KI5Y8u75OBUlbKqGlgTLnvq
2fVczlbuuYkxDuAyZ9unYjhq9lN8EAb/xC+58JBX6FEEtkZXs18LFW5//jPeK/8f
y580Y8H47xPUqQFDOqqctCZ/zPEILIpUOF1ThTeVbRcb5n6waJU02/QYcS/JNSsb
HQ7u0mV3xB+g2ZiQjmFKxtYG/pgLzdZB88t7jo1PGIBgDxkV49cfYMEOYTGoj9E1
qJDHaheiQ1KN6Z2fPhDgLmRkYrCPx5rKDT/44/fF0ZXzvPvsIvC1e7gRhke0ysya
0yL5FzY5M00vljff+tf7s04yZF9cJxRhm4yS/i8f9zZsGxfzltObA3HN7nYj7j3l
VNG709ieh0hPEROG2UPrKY6kCf7Pfto5+lHHB/xCziYEZZbIB03Qke9OZjCcdbhJ
puNws3WISWHkI2ReGdhvNICIoxYFrIHsVZZBmk0prDLVDTnFnziagKzu3ngBwAKy
rLA9jmeLnGKLI0JsDZ7pk34NvsioZAOedc+Q8YVw+Eh5wSqdx/uwPtN49lQdw8QP
uVclIHBqdpld5mCokCDk6Du9Ns1wC35S8+S8nmIwUO2AtlZ0yIN5XtUskP5pSFYe
Kf7BZ0dlsedvLyAlFFiyKe32rFg/wt8U1TwfAeoAkuUUIIabGncatajFs+eEWgwX
1dEqrBKG06fu2a1xhBoklUC3MbZcPy6dQ4IVyj+wjq0qBFrywKRNwOg656NOC6Yo
HI67825uQQ0WTb1ktNmZl0Bjc3BnW3KYqYzo/8Mgyv0P+514zDP1vgqmBQjhSw/Z
3UWxejJzCJk3sAfNyrZ6bV1vZUc1GM52urG5cQpn2SHfyjQIjPTkBmZCsIPCI8nb
pQ42CsU9x4zuVhjjm8EREcoT5apQUFkUINoB5EXKVag6luSVEvBuV7lFzxql5Lln
yWeRstY73R09qh/WdEvH1XKXw1Mfh4FzWbcsvleY6igb3Gebtk/gS9FLsIfC6Fit
0CMytTMldrwSCQQei7wJxl6NeBLo76HWPmJCDbbZ1TjGx6o3sD+STeDx6TQ0L2sm
IOJPhEG7KM69xBhEAR/5fvlH0DU6V+VFb9Q4Gy/ZAAOfPtJ7tUm/GXzScGwdjTGZ
35EeaW6dA2aX5SBsSn95jK7ne5ZMb/tVLZlDWYDBSCky1Y+Ju4FYk0DzvT2wEnsj
dSCUNUlmeVmP9woSx4LPr/274SNqlS3B4hjQZCoMNalVKXHOafDceU2UM82QA8lc
oorC9ApVv8hCl2sjyxTm3ydNKffqqXXr2OS2OO21Dikf1TX4u9+DYjPg6Z0BqiQY
us9k3fvKt58iPyH1EhPRqXyrF6P45UYzUdYlLq0g/b5xiCvW2MsIxNvb5b6J8joZ
PgNnXNJ8S4mvia7+S0Fx9J7uYrmBNkBf/rJflHcFQy2IdjElCgK1hR355X9HcfiU
ICp3bS4hrElqkxs+HYqwstGmK/OEnmMqJjp2u3zMZ+3BG06XLSJjnGBIrTnCxWLC
kYhZV2813gdj6v7XS3HCZQxNMw/P9OYUfpipq+OLp3yhV4atA6mk/ZSsdo3RtRGy
KHqexLc88i4My0C/t9j7Dsk0nC06+kn7ncrabOvJnZ3YphaVpNt1erUdW+Jtm+TU
VGbiV1W0D/prjWCGGF67YbVDFGMMLLdWWpM85A0mLmeon999kIBAViqbfdwK9Zc5
TbgOLWUl8yZlihrxN+6icTdhiHm9MIdiCPIBZEOhGZw2Yy5Ry9Gk/fpFujgZZRhp
25GJzq2wFzH9ieqYuL5ZyKr23CO+qfPZ95iBJGlVuW881QMNdiGIZQAcQNF3kGPF
HBcOqguBszB3Scj/pa6hO72SyaRqTVd/DKZOLNCECbga3mfmaq3/ShpIt/iAKT2p
7XhJVqcai4jN/2R+ptaMEMHRpZ4RcqHubausz7qc/CGc63NbZjE0N8gru8qGXyxU
7g8j+fOCPF/IdxIqAZ+b54CnDvmNyU/Mo/IMQyF6REM8HWdCnORjjFaoo9VrN2+7
sHd2OZKKb9i6eZKV8112aKgJ2Kc++PUeah9iL1uCFREPCJDF/um907x9uuDEgp0D
xDr0Mkif5xyGCJA4pdcNCmUYVzXCYUKM1sw0hV4+xIPcKfPSXbhxq/+Ag85FuMOn
LHavfssAMnUtEVos4xydbipAQzr4oeNdSxOODfLaQP41BGLdLrSZnCpnWHaP9H+i
Ffqf29Ztlkp+w+C0+MYPrz4CY28Z5ui38K3LDgu4CJeK3QdqDwWJbrYppaCT4uhZ
uzUL+7sTCNWm8MAcR/Vo2U9wvuKgEfF5hLg7ow6I9lDntAgwpT67Ts3DGJkBIo0D
QjjNJtYhPHJJSkhQ3v5LQYLMCUaSr0WOiRQNnx40ZEXwAAt+sCfscY2hmAuudbM+
mcoYy3ZuLcJjT6p4lJU2Jaul6D36xtxZWj4VBADDVxXkHU9fg/XDbEMxBjB8NZy2
ckZ9qKdW+yrZz4Y0vdgwtaFHC9lokIEUTpWkuYY9eZk0JEgrNE4ZHV5tL1g9HM9L
8Dw2zkCuddbqsEwakHbazjGetNE5lrzw/BZiELj05gRlHt6ff9dxcZi9gS32tf4l
7CHL1nxPoNuNABMS96CAyO4Xlcdp4PQWT0dCMGDmR72vraB049Bg9ao2h3K5fg7k
Gfz/fEKg7YgfIjB0d4uuIz+hNajE1td/4DpNlh4tDV79/xeVW8QSGtuVBXXmVEK1
Xi9Ht5UP974zYjdczmx1oiPvQqn2dbgJSVIsqX3bQWYksFFwX0A/Kt6TdOKg+uAO
jeuIgaDu40OCQts5eV6o7xu5BiIEbE+/NChak2ht9nq1BSFV0FQvSpLlol4y30ba
H7Y8+WJ862GdSpFBaPeXnTuxIt9/Cr0zBzR+zjGE8CpcSxzsg++Kn8U+4kMS2a01
Y93kJSG0wiLWwprfErNWcygNRKg+o9LubCUOjno/sGd+jtRFxwW3XbD2KULc48fn
s2c+j83L0vx2D0ogDbSPFl+b9bvDJspMufUaxhAA6Fgp043py6pMMMy4y0lum2+E
9+5GFXgezqGdi6U/Khszaremrmcjj/XV9QfUj+f5pQZdhZIydLlR8v80k+WJ0KWr
UnrsnxrIoqAL6/WNNRFdD8Ya0VClAtGp2DYN8ih6c56ENvspc9IFS1ohEepHMvLr
mB9pYkqG+pPQrWuTWyd+vcckopGCKXKeBSXm5S7V3RGTGeBBe3mxpaGa3tmqYinL
btYYWXZlNtYNBG5qlrOgJiwIh4AIoaEgFtgBULCoeI6bfRKR7KBCbSpMmgUBx/Pl
isZTIvXR3vpOk8XEepT6XhDH5T16Osa0CCfM7jEimtwwxjQDj7cIB4rjgFs3JW0D
yrTjjOIVlhJRHKj/t4NmAAXymovA3QHg1biuGmMR5QQ=
`protect END_PROTECTED
