`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SqxlmekojBH90XNnqxdtLV8cc8jnLT6ry7y64UI3kNU3fe31L7KYf1DowD5HObDe
8IJC6LmUSVTLrLjJ77lLkkxNK2LpX/N3cM+CvN85VzuCFfr74zjIFgeuDeFTSX/U
2QNa5sKux7PQy3QSu17D+5eF1w+5S3mDSQMfGmBSehgMaNDVnpUmMfrTNF9/cMhw
y/JWoeKE98iAJjEzI5FtRx2j0HeKwRhh1nOs+wr25pZC5ru688yJtQjS8y2Wxq9m
NMSrD6zhk8RJlZ3EjvZusNO7htzhVi3i+n6UNnolwPVpKICTE7MJ7UCk2dlRf97q
wqmv580YCcauREdWHI/ttxvroXTJ/gdj2DWjaEbgxlXpkiCb7cJira7LlVi9ljZ0
ySSonHNkSHCSBCeTAUWAVOuvHyj/TN6dv+EAy2dZS6JjmRqNYhHcodGFW+MbGp0F
sZyFDLVy/dJJbs3DhLTzOYApJXeiwrwYfHapkzcVsoMMRjpcZoMKekpuLYMEnC7a
AkbX2ZibKh40Ifcc3SUNt9ausdYJxch1fkFBO/G1YrD1YOA7pc1RjNyzeIAPtiIM
q8nf8n+4QlfgklmZQNFym4WetdEfHhU4FxsU2xT/wlwhflLpmdAm1N9NuSdOkW8c
HudTWCQvvIg3ruoTCnDnzhwgxoU9IcNxUKQije21XQ73kwbrE0gQVDtXc+5Z61To
kv//irv9agsNK5P7p/sFm6Przv/qMeq5CuT9bRdysgqwjvjB8mHujzrxDtd39B32
hEx6EMPjEnVJXSj6uSP0FgEhE3+C/g3JmwWNulAJadQbBX+uD+pqmmmMJhkkUAZr
oSuLr/CyC/GFfGTPjNdYmd+pvWCzENXl/NZUZ7Qp9pMDLAdVC3XyCExMVszHlOlO
oin1swRcWuSNKQtXlLG02sDOPS3AX3JQnsabMebS8PF1zcZIRqKGAfAuK5rGkcrw
j6YADwz1VQJhP95iqhvYseFK9UAC3PEiesVFC/N4tbqgYAOkVBnJa1AYcTOjMq6S
iuwlIZZF+oPN1HtLRE0nJDkVszazNcCMPr+BanVFWu5kFS+4LkV1RVTphrYeEkJL
PQZuuqK1bOU5jIynIAnrSUYi8/542sZaoJI4lNs5KRRachs+oVSO3ZTok+PEdowB
K6pYxz3lIgY+kYD4kD7iM8HlColgviWdodUFrST0zhMnm4tKtrsC2SldCbG5CUHY
moUanFB74hjVq8uT7evNBFQy9zrDkYt+5rDenFnfgDDAKnUNxbeTTo1TFms2BmBF
9lKgqWqyrsL5+1EWoFF/3LSob8kL+wHRJ58LofdxktU19CT8P6U/B19YreyDraV6
h7jzfmzVQRJEU0sb6Qo9Zeur13zPFN0e+Zuty6Ybqq5xXbS5TKGRREavyX1wex6G
gQgIWLVtea0IhVFBLAo7jhzynBBdstwEeamKAVNG8yFj8yKNd53NuEf+u/dRKlFQ
+EX2CVL2sQ99WRgxkcmrHgiQ4X+pAM4Xu7dNmY+xJWHVaCXkIjgqzC3BPGl/FvMA
SjWJX9J7MB0MO7Tlxt3RauGa2UTR9eFy/rcH+iIz3Y7a5VXhRIayfomw+bbYng9R
r+oBTHJcfFMGWyXFEh8bwQGLG5dxkmsKd/Cpa2q3bcKF7mAIIhORZXoCLHWsFObH
AMQGv/C++xpnNSs11Wpv2QgBw1gSPi94vWSU/Qf1BWxP7gb3YhJs+pVVOmbJN7OL
++38Ya+ULPkT8a75z7OE8DTzyXkT/Q4WSOZbOW/iJYP3kaZgnOffjGSv0wG/veLa
bYzz5gqX17udan2t9WUujPQf2rwlGyj4bDuvdg0vcB3mUKojjngpjcYxHujmt6dI
LNBKFDgdr8FqYLb3Nqa4WOZ8XmV7UvybYkDEU6Vq8MUzfy+CZs9gBVZLUIsBFoES
mVsZEXetvj/RYylqXmFON/hBNnd1zCYe2kIo00+jUZEzhRURPCFN3KsIs2qWwJR6
zd9T/sgWMKLJRQFoABQ0v//7/kesSdWs3yw9X66ry5d2b6G+tLion35VcmAhhNxw
kEQBk3tEb1kYzST+l9PYBPktCJkaEzdtPetRpFRP7Z4pPXrZ6dYbgPrA8DpABeLt
Fuz47aaLxzSEydpl6VXYnVXqltg2WQYwD0LjgYrvoiAXXJcQkWL8FIhw/FwswAuj
JhexJxfImzLC2s4ZRKe6y58tKYfUvF6vLR9lwTCIIGi1bdOzFUF94dfKqSPXd9At
L1XKkAfQTqqNogk8ItwzqRiRcsvlDee09F4I7zDqt1Iw8s/VGWWGfu+jhUgYEZhR
McF4kFX5sYTu8muA8s8titjOklOUBkAPYJAdEi83BYEYURcR/I/aZLJrIlcYPsjD
bC2578OJp7WzDeRFRzQ/dhQhceEN6r/17wJB+sP16dHqhC5ftkJEfki/CIRZof5Y
iaHqFEchINGHmlCJhDq+q72+qGU2V7QKKmNJYgaVFRbtlx75Cj6MuUbs+N3aPs2X
H088NaHQ5G+l9cY2cjiGX8sWImcmiURkUMR0SX4J+VAELoPzb9pyZXllsxhsr8VZ
kAzR5pqhc6M1J/+MY5JygNaYMOHajTyT2oI7l2uu3kRKvTL0UwVsxCGSjqa+S7jt
`protect END_PROTECTED
