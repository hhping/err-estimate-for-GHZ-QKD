`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Et54D8vPAIgHQozEQJ55+6Qm8/4wl7O2TV5fRyctkiQlZF3ZkFLSH6AiGgFz6sBb
lVW6uMM0KE2ybyhfRe2BXAcOul8y+eCJeEt8gue9bx7Rbvmx8a8+JDH244mE4JYJ
c0A+yxPLl8puqeOv0nAwbMlvVJZjYfC/4nkvx5Co2U0x+0F4a5c59jCUzTTI8ghO
I5e5pd/eTOa1e2eUdkvSOmaHgBSu6ZnE3gG82dcsRkur7aOVhg+l/2pJW0YHGa/N
FEJMAGw7Y2zQnWqCv0zY9FNs40eyT/Jy2yPWA1+6rMB26QI9jltUVi1iBiiehOw0
yy79G4BC52UlOwyf58MkD1+D6qWcw8ATy1h9MKL6KDWW9OFqKwFRcrH3aIbMeZC7
3tlBuH20bod98mTwBFiqEA==
`protect END_PROTECTED
