`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZB9AgkHrFxLZgtTUG9Fzy2T7ZUWR9Xz3BqfKyCRpaQE4UHcO7l/9PZwOTESDNtaV
l8SDCpVdf+GS+/1h4zOmWf0k0zMdyX9llm8/yLy6aZUKsPYgxikMkrlfroRF3pzA
PVbYUIxr8ImKUd6bvfChDRSbC9gJ/xzKu0kC9e/n4EB5HemzxmU5OFBttAWS184G
a0Klq5IVMx2c2jKnWN7XQ8uy6DrCZ8lJUw2pAndKN1v+tHmqqBm6BjTAlHzILzR3
FUCFXDmqs3g8Gc8MJVWnxXyzKaz89h+RmA+cS2VeDNEnmeofaEwSI+O8hvhvFEKq
FQSSFRKDnj0JJfQQC0qs36HSUqNXvq9/3EJIm1RkGFPqdCNzkH3TS2r3irluE1LF
qf59uPoQ9UbwfvHQxZSrBbnVDsxJtpCpFiGT4e4SIZsUwTBEpl9A8CzNmZuxxGTW
6lIrIapVNeX2jR54ZerZWkF/xJ7Kx/a/8kzEgkTMAZ+yRDcqLIe3Ethj9l9CAPie
wgjoQZGH9UoTI93E7uh8GLuYgN3z4rNv0KeYsoJKoMUI5JbxCY2uRw/zdkzVR5Al
3Y/NJqD0uk/sy9Z2K8ybD6LTrUx+c+crsi7aA1XJq5ecFMdXDlvMgAU9k1qRKds1
GjM/DEW21N2bfGKO+OHVewAZEIWGtGGMwyOsQOoEsQx6ByT4zZaioH3T95TayDFr
qCCAGiXiBounIutvgD4NIQ65bmBYjFbv1QVKTCNMKLqCoxHjAAOJ7YRONZmwVoHC
k6tntOQW41F4ajRixfCl5ZWlrg3iFiSjVe6uD1W1sdiA8Z2n/Jy+TRF6it1uprbp
95V4l0Dt0ApLbdO4tt9t6HyF0PokmHWqHPA4iIZNMyN8TPy/InAsGjKGi5NpUKiv
XEoXuCYa4usdp1TXCAdguT9c2O4gH1E5/zrCz5WPrvo/dPd95My1YkBptMMpdiFY
OLCZ2Mlgw/BNc/XrTGraGbcW4nMx8JBD+TLBAHSasBwT8dsPWpcsbvj1HhKdhKtB
rG1DcmK1y9HWE3gRvsJJE16CvkRczuSx2tdPWTqTvba2wj6lsb66zGYeP6p3Pkn8
h7epIGewRXy3Grs6YO7ctaRGjAUV//1+ZFsdBg90VvvvOVS9GJC9mb2y9HpWyHxg
FpZSTHWNp3AgNSNWGDGc1/zu8K1FyFg8YL6cgbMwY+Z9I/PL2rewcjDIaW7GzSTP
CCrAxLzJuHC1iYWpFb6zdGslkfb3c8JZ9rJn6Q5egYB4cy/Pcz5FX+nr1/9h8Y7B
o96Q5jKcZuB46I35BX70OIK5GtPE8QoF07y/L+/du4HeFalb+J1nXq3A7HNtpAxx
OCdRTFu/mZCxO+gJCUeQ7/5+nIVBqNybl5e9exjVuXJt69c4QqzwayGozMbgtRrV
8M27h4NZrGNMl9rr3NI3BwM1nKpEt2AdwwuToL09TXGuyJY6x7TjrGdVFRcJJWw3
QE5+v3rjP+9shlkCHuQhRl7uT+nhw1U2dXEN7Gl7u5PeluAi4H6TqeqNLZEHiBAk
2bJtJtwrUIv+r2n6tfCTJ+UX4zmKMlfvAiuc8l/k9PJZofLcqMgwyiYEWaHkzPIl
WVYeQJTUpGuXgpT9dxUcA4Vxgfq6W0StMjqCQSda+4hQJdKzDejon2dK0V8+ZZR7
alMVhoKXgk3P8Fqi02XLw1GXW0XEowLUQcqkHNp9/GjpnnlEwY2OBzuSPSS3hyd7
4NP7LhGdB9SCxHSCuraiDu9fG7zG5OLrmGMhrVb/Nr2WSQp0SJvLyGwDre0oD2Qn
gdfRePTYXWZFkEcCtAAD+UXjkLDUItC8sGgpSwzJ5MLr6j3fE0Gty/rQSNbPmaKc
eo5tLq5k2uC6wnsJnQKc9Jj0eo5zl4KPSwz6F6PqPyIMv2ly6zH8lOxrOIfKRg5D
JbLOzmLMIkjEXYM56AdwXCVo51oHi5QRVXF2WosOdDknrKOj3+4VPrA4h9CcGefn
kHSkneYtNqT2tzOGU86a0vZli6az69geo9olHddvX90egKn+RkNfz6FPrCqorfa9
VkP3F+xfZqLm/c8hwbfYd8WB0Es2mV7hC4uO9XTCle6WsTEROvy6bICiNwB7iqhv
h54PMyn7HWHjcAexsTXK3sjCm2pHHo6EFLnFyooULyzGWaQ0GOf6TGk52FDSO5h+
aPBlud2m8oJ34A5WFqoK7EfrGUEPDlhwN+VNq7p5EAP/G8vzIBtajTSyRtBgwxhr
IJH1hM1Ffq9ItrLkcAAYLA==
`protect END_PROTECTED
