`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s/jXKY0DX4AMqklYAS+rvrw9ZxYswZ5pgUOve1hXBpXsk55qx6JzqQxiE/gy3Pss
vXg8kaFsRGReEd0fGVYxaBWa+dQUyPuYhfgPG4iiXrmBNnW46pL9fZjjOAFguAhU
yj9iQcH2EgQIIINpqApBIWJrgwEVul74Hag/DWCnBQfTkzMAwNrFi3lnCCBXTw5l
KM9SV31z1fy+HC+Vxe3aUNS1YHDXDpDWm9gn9ilQe6b7ZpFbrSP4EPxHlsAFdvCp
OATQiSmp47S2Uc542kQ2LKubRPn+TH5H6CCOtBJn6sUAF0ZCViv7t3m8kSLIiRX3
S5ZSEiWwcK+bPYptrUhL/6DlMOPkHWb43GB1Ee3W8/1GnNsrSD+bHZwL0SandBpc
pzSK6W3jtokRa/gtYmGYIGnxyudL/QVhVcRwk9JVJ1HU/XvIGhUQ6K66N2vrS4do
p934EcT/BZeqrnjMO0dvD+qGFfr8IlkiyzdsEbFYYYeDGB/4Uw9heOXepx9bxFKc
67jRHn0pddm3wU6MA9jGn5X6yXN8/emKEwk8dC0QgbKzsuJ/uU9mxOIUkKl8fp+O
S11ILspDugRcPnigww1KUhbmNkul6rBRD/dvKdc9ZOdyE/rpAD5I2k9WncdNm+IR
dD2Zsz9OayPoBq83DyIomQaYD2zV2ajZAMcRf1vztYyT7ZNw8Rqn8DhnSdGx5tq+
jODMQjbMekclW/kcSO+N8M/9rEAlwKbXnQmFkrNUjv0rT4Fr07GRQ6b+AY5YdYK6
wFs8aXAA8MTTUpdDzebRqvw+goQDqLSjXYFaRuxN9+8Vl30bSjGVNMUq0VU6X3x2
H2rUUckCA60K6OG9Y5Yuo19pZCbgfINVWxUG/oPLKqd58Rd5zjmPK9MQd8iQDarQ
38mp4FYVmrTgjbsTFJxyHOgpivxqte8XtEsrZ09Qu/cp5fy2djBSFMiEKuWO2yE0
lw3FiRPTBtL5qPzayUHuu7dmTdCI7DRRqaN7iDuwkTiNEId5r2dZK6mNPXVNGV9p
ashCyhaKIffpIW7ziGo/M12FqaBBIJU02FqWEMTfs1EZ+aqLfxwERzxUQQFcSEpN
uF17rO+iyniwO+EhIb6dJVmXl4I2u2xvIHXRSOq/TfVATsfQkc+Uo16a0Ac0i5JU
QNRIfNPJ+JVDRo05bPQkvpFF43B2cf05lF5wFA96KKHrUmrcnLFxPP6NgWyf1XlW
i+NYMHzdZ1aID45v3te3duVTL3NxlEFT8Hdj8l0zdU1LB1m6LVyB7q4jm3FcKst4
aPCVsZAaj7WmD3Db/vv94R8t1xmnuPaQw2vylbQn6EYNmx9wwV7REKUFXH2nvOgn
fWUgq7K6McIHRPv2+Z+R55ZzAlw6OlYKdOMrT4h4oRZeVWMl/C7N8aJYZ+yEaJJL
Etj/5POjAWby+ZdF/HYCuUdC8srfhuVjmNrohNtVki7k1hG9Fc9K9VrXmbETcU3z
Bfsu+qonp1nPOCWPbBA73Bw4o65os7BfkR3RYWed7vLNTJJd57hj4dxmGbF7d2VC
eGsVNkzjctBXeR0KY7U7dvNmFeE0noRUDQ7fAccdak5FxoUfZ5HqDIXDsYmMhhdw
Xtrb/9i/mJiD6c3F9+fS9LD/wncXavxHnnCUtbSDVqTMpHNw7UvMSTGLvRa96Zu4
sovypB5St3iZ7RnR8VCZ8xraCR5gvpBnPw4Vz4u1V5hv4+sdgZ6OAtLXYS2UFJbr
8vcafPOoH6jElBfkvQZu0wXivZd9fb0UiArGhw1bNAircBdk/Zeut2qgWZiPTIyT
lkAlMcE53UJfHu99AKPjfNFHi4Mldh/0ZtjD52uP6FJIhyDGIcUIQQERDYuRIznm
1+wAbJJjgTzu2dfqYhqe5veeqHpEZFFcrInJVl3XWT4jKfHDvj85A1LtWH5JlH32
ZSyL3gbSMJ2tbtxoVYaiGScWSw1L3ukIs3ROf2jvGHPv2uMdzzTwQ/lg/mgaZ24r
NbGTB1zNf8VGUIoHoSR7eKETFofX0zM6b86Wjz1gLxrLnPFdgRzPXMoh14WNCjJV
SH4bwq7SPf7i9vDf3bOYeN3Vb2lYBzAZNYqHptOzB5EQ0l8fT25AP9IB89CzmnpB
6CsuCS2bf9Z+3vQOa56I8ywH8MeKnA18WpbCFHAXx3DGn5lQ0hmN2Pc+TxGlkJls
uMBU3U/8OnJYNpapxID+8J3y5qdCIOt2AyfKl3wEa/tSdJO5m5ttUzSxMMbXsrOD
jo5jbZJ3eKvsjnO36jrZu2IT59j3ukYovUCUClIb3+puodsxLTdQz0ycdfBKFEnO
jvoDZD7gECeK/W6xFxJ98aIS2IIv73p+ogSU8HfC5v6BgEEbzhXKq5IXqsS+z065
dY14cjcuXln1tAph5wUNGMBSJOBMp83NaYLwr+2LteC5BLiPdd5UzRO+gk8AidgM
wkScw7pooi2zBO+hZ2ZMXhr4YHft2ia4wyTM+05Q8zjiXdm38UhuweCVFZFEfPpJ
eoe/vUSSOZlQMG1yGuL9Zr/SAk9laoEmhoK48s3hEa+Lm8IjbHEthRtMeEtEXoYA
rKTXvc2hDfV6tM/eYjnu+5Z4U7YAviLcQ7N/fyoTmiPYmsUxMOXm6fEAl5OXGBNj
/dTjmmuTULjBwEKOJNFnxHrxcHGl/8dkcV+RcVm2igX0heHz01jh0qMhMt3ZcY3u
lgbb4fGCuUWKFrorZfDt8ahN7emTYDvetA9aNA+Fp5clCRvplLlgjnvkeoBVkAy5
L11Es4hy/9skxaW7TKlAOSF4JmvJ7bAiM38JVibC5XcAzP0apbbhJ/XF+OOibHUz
pMJRuyxYbdZpiu7EQzWfRXCM4KemUYQGDcgQp2ZL/Em+77YwIymSjkwW3n/qs0kW
BOpKJLshvB4RHGXGHHw2vw/lK+wnrwSILnBRUpiLeimXIA3Ol6JhH1Jk2KCXCTNI
x/SDDyKMXngMoiCa1VWG8H/WmTK8Nkcc4dapLaZuPcgwsacHvhg2xgTzTYKKEoNQ
ozFikhIuAWSXC6CHhQoVuXfEEdH00ATNBwjc7fG867XdP9s+zA/3eScONZ2XUn+R
WWBQ1l8mNIIw/EVr3GL3IqmUyKKpmfOqemJGixC+eXB4QZ1fQ4RotiCvabW5Oq7F
9c7u02bNhupXd5AjXlMJYqdDj4fjppsk126X2lTfJeo=
`protect END_PROTECTED
