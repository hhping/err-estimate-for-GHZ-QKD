`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NpuK6dcF2KVZD6jXAmtaeYzPS/4IUWbJHSvK3LWMpU3ZccCW7Zh+oq+wvnIJRlZ+
DPox2x9+j41kWeCAYC1MRWPYNQWVDtcnmsK1bQnqd0uEVubdwfhCZmzqIL0+rDL5
CP3s8uG0781YIUURTfxAgAjfrSUHMuso/c5PkZ4Nh31Ur2x9AyF2QrR/buy6X6Xu
n4TafHQppdyjgXYY8a1nfGnLY42z4AZR62hhkFAif/i8r1Nio0AkEgdpMRZ8vI5n
4BmddDcDXr2KtASJdNQTsKBlXItpCjj5Q4C/QxxmTKRTqNruXEVhxNYk2FBd0bbt
TpYaIui01ngvdedbZGFPTk0vOP1F8Geg2gwOMV/Bu18328LwFq1pT6uHi/PP4qJw
i8Ecp1gdD8VCiygyYimBVKzvH5y4x49PZ2nsGyM0WYIT7MYVRhL5ah3huBe1ap6n
FusA5K9cYcfWcSfZE+fYUmeqNOaotWa6s1Et1NwPLRzLQL4iZPB1c7nv4O6w00ZM
Vl5Svx2CZAzBW+fLQ3jz4cgB+s4vdmBSUrqni6kR5QqCJzOeRMSvjEX7hxIRomep
anpY/icr6Tj6dSdp2j61GexDAH2/uWWN887l9C7ZhlNo02DoDHqplxIIjE7+DWfw
RRLq1U2W8dUkVIrz8ij1JkpbMNl0yoQieMNnd/ADu0LfAuhcUlr35Emk9N/U4uiY
L5dO0JwZ7UF+8ooX1AAe745GpCemByZ72+YmKkDYClvnskOWxs7UTGnOVv39vQx0
b37ofwTwZo7DaNWW96xb4KXztP82GzqSCeYwUaMg3jytCEWkxhoBbX6rne4mHrHi
QCxYv5n0VCuIurv+tpGBqWV+LYLRa0aw33iVUQZ1KcONJyaqC3U67LuxedfVmwUP
BE5rCxlUajVp1gjhfoCeex49Aw4sXIRGV/w5CGVD9FlyvVKJIbuA2gAYUhpDMcah
VbMvkW/4SV/0MN0PyvQ08aFytzWh+t7dLFh3jwMdwuga23KtKTpUFlma9+B2YNh2
iE7x2REDSWZTORK2dQfereNTYq2U8j4xHvIC2+P52MomAZbzvhBC+cDAbCms6WdI
ONal8j6NledV5GLJ7gnUO3vKjYfz/RJsgWOyKzWCnZ0orgdaCQ4xfTwETPHLmO7H
cWvl2bTYrGAbmmgtFtwC85dQCl8gxFZ5XJItdWy1B+5pA9q2SE0Tga89h0cQMujo
kwRw0JHQBb6OITUJoaNnC5qYL7ftWT1D2vAz/l9WKXNoEgVNT7y0zeNJmQDT8Lcx
zKbj79pxp99D2XIBhrJl6GWSg9C+BJ5chsNoUCzFyXqxwYaZ2oFCrLzGF/z8lg9h
CuvXm41ABlFBUYvPYle0FrgXFZcsWnYPEr03T6lVz7vPlm63UZVCsBvoYSMSCjC7
Qikl3nEh5dZbkuqd6Iyn5kD/d2PTqDbkAhsOhyloBDP5jO8NZLRs2Y0UkCzF2N30
QXyppK2X/EsFs8VgfxOEqd+2b+PmYfg1Tpk34JPItlAdmqP7Jl8tfyU7UAYTvhQ3
eOk1rv7V22YdACQW0vzkXY0NsjCejP18aKXgKcvwD+Ogz70yInC/T0PFVxNpg/UT
77JMUxcOEwoH0lE37KKCA+QXiacZIjslYXedBWvX7BX6/rhOcCF+Eib/v0FzuRpc
WH1ZyYPUjgc1forSK+xXd0gIqz2wm3ydF9t1d82jExwMoxsrgacTNa7yoJxbfTmN
+dDTOcCNDxNlGHlrI+GbJ1ehiACGV5L3e/8c8gTSD2H12/qgZc8/uH2VOujPBgLN
rncWpQWfxVYYM77Sd6ft+ZXXpKkZW6EhZFIyKviJ/sprDmbEQLxb0WySXMFJtJix
KmePApqE8Aws/UdPB1o3V/z75khjvvaxI/M99J3uqW9yi5c41V2Ux3H7OA9KNGwb
Swe8HWCISsHQTLCVIlfiBjOVIb+rF1fkS83Hgn5l+uJveIzpp5sSSszC1rKi2nwr
R3VogssoPlkxOC9AcgYXKJRONez1mZgAyYh2vwO+UobZO7ddpDYIXktG0wNmQgoc
8SXwp63vtLf3vpMgcvOoxMLan04YFKzVHESJXPn3n3yz5MQRujuvPtNKWEj7oBZq
cZpe9qEVfS5hhb89EsC9tLB3dzMfc0Z5/NV5Cql2d0Fu12QRMDqlUWFxvhYemf72
8u1M/GRpqZTAwSsq1h5jmvWs6qWGKd4Y71xV0wSXkssiIBDHKa0roILrRqm1IFiV
3nTjywLmKVirkUVeAhpqEbMkUlrPWq1/Yif9mPuSwi1r4mehXcJcvQUNelrmpK6G
9r8zdTOzxR2H8sYPuQCG0gKTSy/o8Tiw9VJpQqwrSjkm1nX4WxTe3kwyiuXCUkog
8jcYxYwZE+LHSi9LB7Ts3A1YplE4Jxeewe7rZHyefiypxbbGO64X/ekpo+YLGZnQ
LmU2uToUvvL2Jx3AH4CkcDnAdeVeIx8kHcy2UyrpV5cXGW3TOj+gEPptLjRo+3yd
/FeoAwIaIeNdXMTxqBQworAIPmHkaZz6Y21phEuRF/N82V3QrrwNxSWopgALDnqc
AZZ+v0PZZ9f/f4sHC9vtx4ITMGvobXWgVMFY7YPwTfSIWiVU27BhNYIHOjcFs31/
2+M3qTyRBs2aIF99kqIW/YWMOzSO2g6UzkI/VdsT8QzP+RpErijjhKcqcQp+6rPU
IRV02Sx/nreeHCrEp6zLAU5SH2XwkCjj/tiJIdfMB+OI8FD9WGj7jaePN0UXPwwe
XknRcNedayleTxlDPgdmku0hozBbnu8qHW25Dck/ClZWYMr/TOgYW2s2Niqe3cCa
TjLttnGZEcyI+o2RRlZIhrA19szHwonE0NW+nEtNd+PoLmgIiHBe+LvJzRHbpi3+
Y5IfUT3tEpWMVmCijTwglKj6loQKa/u/kcMN1mSREUknUeZ9SFf3Ny6AT+hOaSvI
/zQ5frL1mmM4aP3nFXtyH63yiSYFkPoNmMsxRslOX0wkaiCYwhFFBpmGih0dswei
H8ZMYlO0UN242o1zQY00rt5Joi0zeQVX9PCXnt7WdMeN+NVCLIluITbw3SOb8iDg
9TIyA0CMq1nHatNDgKJhvA==
`protect END_PROTECTED
