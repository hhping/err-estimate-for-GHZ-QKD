`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nnawszUNd4hE7wiagauEGfDomjcdxVH2CgEUSDoDLut6clceIiEtX5bIAEUQAi3E
FSMEoAnq10ifqb1yoS4Zin8lnAKbKOXVnr51mBYwsoiJiTC7G6wFRXSWDvBUlYM/
xAhza2ZS3IQvk+DpIhjxQhD1W2dY2CpGfFnbu3554vPN2PRUSGyAgLuw6GmqGz0P
WMo51MtZ75ns3+3fn6JYlssvqNoo76dXN3VL+la1/m2PtDvC5N3d+d5JTPutmB8X
LiYGCdwTvbaomI5l4zr+XBRM2rtnaPcSfA1M15PryCxOUhYqrDCEK/f+IPTMql56
35oI0OAhrik4eKwg1FXyUQgWnEUWVBWiX/75PZ1M5eV21kRtxCibxBLYPqgWUXff
/WQlEMdS0bXsKUlUvXz2/0HjSMpT14XJJZuFJ2XN47Gw3vPp+HAwoekQVJ+eM68V
09JSD4QzAb/Ny5biHGt4VDKTDDdMkPx9d8K6ObZ2QOPwe3M13ejwzi3t8/ZXuT//
KzySS0qwrfJ26HcCi6BhNPyjNu/7FokH0Ks9ymt0LYqzKFA0jLn8WsNzdDNTpEk1
jy2ZiBM070WhmJ0lUx1nBlfNlDHCQjb/WqpHd+TEYl4e4xjtMrKIeb83uioLqNyp
Xqep0lqqv7/irNendCRph/AjK49yYvr45x814+qjn0C6TgfZ9KQ9QC1dHHQW5ZWf
3iuUOeNYUyhYSPmKwtiBbhuen4MQL7rCnG+MP8Gsq90nh3ZVwiwP64yPt/VLMTBt
92mM3E5kVC9xWS0oi45PStwvxo2BhhaQkt8CH31/10WmWPd7fxy4krAjPz1acJG7
XmBgAdtamXyd2paLMz5HPrOFF4MxlHshV0vxxnqoQif9zKb2JCYsG2opP50YYlbO
il3KDgPkTzbGmJWSkSWLg8gqiKYh4kZxhzetf8ZWTiFE8W9ofQduNvWHJIVcqV5d
qcG+eX1pKUVZpDfvdp4YkFKHXAZq5SQyvsL8C3f+Jco1CV2k+pq/kbMhvvJivWS5
kpT4DxcYryECMJKuDC+pP2ZlBmAKeGZzLVDN/pwWM1mpq3P6zCkOqbMNrmEZy0hg
P1IXT0WkD538YOzGcw4yTnclSITBIu9AzH+EZbKU3rB/Vr2pdx19WvH+JITRjOLo
0FYJbnrrNxiaNgKQaL4djXCQ5TKxDccrNUqovFGjyJgzSyaM6Rd/bMdcKJAaGlJW
aDwhIfYGCifKVNKS/fV6jylbkXPf7b1njRAr5EKYcogSYOwOn5n8Sef1ngUD9+ke
`protect END_PROTECTED
