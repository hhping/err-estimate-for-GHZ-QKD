`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eK2DGu5/DFg9iIWVBWPoKda0H/eLmp06c5d8NNwKLCz95EIJXb5j8Z55RZGatt7Q
viYaVo3+8gO3xcRwiRgIJ/aTYybWmkK33t8+6oftxeWGA9/pWhhW8VTJjJ04L+wi
357rVX5094i4l7VFfpgmtKOR98zV5z1T6Ij3dNKmQWP0S5YhsZWBJJjktdC+kpIT
gRbby8FYJX5vfJmNtF7qIb+86K1/t/EAcsgAEOGSZUTwUVYcYNIUEANmBZ1xMDPt
ImOCy/CPEFDpj+lcyyJiXjav+Ha4NezNdaPaIzOH2dTjsC/3inBTCGyfjW1jN1Zy
+ktmF+nRZWnbQ7HSeJKHP3cDl/zQXqXgBsDJsE8dWd9u2Tg13Fb9PIGIn7qvSFVa
PuwB5E3k9svlprONJ+ZyytMbJvxiNmR5C67ivnH8L2ArLtoGTSvRaf6Ay1+Eg+PB
FeYCKTj0QeXDGw92TaBaLtGQ47GPV4OyQomMRwJduAMTXQmwDlWFO8v2mQASjQXF
LDEbam8hyvU+u/Zw9XG+czXHbo6DHDV+SC9xCsq+zXvdPn3j2s2MJVmBvRi2Xd2L
KyOq1j42MhoT/yeeEGbYo4+WOJthg1V6Nvqa6P7U1BLkkafzimYPBS7NxBo1TEXL
quK/SvJ+5kR8NyfIZW7I0GwLwHN/Hk9QyesfJhHnuEHpE7OSO4Ax0S2JU1DaTlcC
yTRttDojeyTz0Lw0xgBM5sIVeP3LtjSHO7EuQfWgGaZfE22ebOYBVgOHJuctOB8h
MVEZZ132DEgvU6S4cZSuBw==
`protect END_PROTECTED
