`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i9CN2JnmEXEaLfKSlJrGfwwidEqNpPTg60fsHa3E45AwzlJYgSKre41mhy256qtj
Lkqku9SRlC4YyFQI8cTWPiBte92tmXEpQx7GieQ50w9/CDR13Eg60PDqumPuVbwH
72LyqFkhY+Df3ya6ZJwgPlMnDOmrSCefA/WVwvCGxGGy6AV5HIROeBaBw8WznusJ
YkgviA0n+WkwRd1J80qPemg1115FX0uSlSG7GNqLgfIUNOF4wWgex2rx06Xrc7Xv
zbTmfusX7Aa2eXFaBwpjnU0ih6KOiHPrepohCk70YphxY2MnF8SeB5/hD217KUHH
vZ+mSna6FsjTeJ44IepleFkrEOepf16wZ9jZ1IWVycyyVwZzM1L7XpdGjO7Rks/x
qC1x5YZnls2mtDtDHy610/fV6ekbYprb7zAEYjTfif7JPklDBIexGIRqeMD9iyf2
YhqF6DWYCuPJVN8oFU8c3WmElRO9cT/FcWV9p81HyuMiGgQkSdbeXJwrJn6yGhVf
3vDiVaSWC2WhLtlJlRnHFYfxOkG2ZLjxafu4Fm89x7E+wwMOLojlPLwBS1IrWU4z
3FLoSqChp4NZFEowv5KhywuDYZUNALILO1wjRZeOs5xeVSQPKP3gj101/t9qItT/
PNFrpNk9QbOuPWZEDlrmpdoEnSWpSXXyyOUDYApdspKJUyKHp5LwLA6x6PWHu/T1
rbrIQx+OmMmvPFJVl+boIZUPBAnU+ZJZpYJOW3sFl2oXoMJsEeKDsL2RuCv5J/2R
xTTCbpREjDstcYbi40YjSRATVYUCzudrQHKPKZ7fXP3tWBDeurxYV5+gLwVN5wZB
57TTyl9ozMhZQb7eszi+axfBQmn/1EIVJBjjmm7nv3bJkbhLPGEEKxSWpxys/S1R
Z2eGZe3j+5zPcEpCSULdWt1EqPCqBN02/9T1DA1f7VTgl7tlJfCyfKi4d13TO8Uh
gJFYY2miuMgDBD+rHQSJFiZ+OFA2/ASwd+3INoGdmTBkr/j5Gi2lJ243IK3Sa1sy
SLQb0hURU4LqZhkjKrqH/kcBqjQ6K5ptJgdR+h+hNRgN5VRz4un9paznarJRqSXI
2LksZA9tKhOaa+47dxOWmVgiCFKHZn0khP/9Y1XaIUU69759S23x7EM7XZdhAsee
bzo9QfONiM1mj15aAXIa1lfVWHj16G+Gh86fpJtf8vIe+SWjKFM1kOVRxi7kjBa2
sz/xm/ts74Qeu5m3l/Wfpt661a1lPcoE2OByE27kAL+2s+iZbw5ASR5Ve/EzIWmv
AYy8wrjjoy1+NWckwgL5RtWzoYbIEnHnTM64D8FFyZkWmsIb+HBHoVD8K/bKGxWB
BkTscsxHukVzwLA3yJIA0fIDm1jRWQS/TBl7yseE+Yw9h9mfnUVb+aGBgRy1fmLP
D9QkExI7b9lwoMuK5LQmx39xtPyUibztNCf/QeJ9CO2JKBoeklzfpCMzcOXh6xj+
qa5GSm5wvuPg6A5eXKLg9ZSplU85wmK29AaYOrzzrjKJfK0n5+ICo8u2nWqxsmoi
1f4e0Z8S45vnkIc+/9Qha9obX4Pg4xvODArnBb+LAQbJ6I56lX4pWrA2s4OfWJOv
N2jpzNsFQHtaata+RP3n6J+ns8p/gLfGjEKaqcWEnDIMamKLHlPd69joMDB+RmUe
wC4y+SoTiy2UA3SMHEb4GNi65O7RCUb2a5d1R74dZbVPWr0J+lOfU0Lk7zex4YX1
xwFI5UAXYh1nDcZBy2cgXJxE1wIFBlUJRqlz2YJpwy8H4EgWNcNzsD74C1UO/V8O
rII7mSyPfYiffN00coplJB7JEQvlIjnrbLOV4qyBmijpKd+ESyT1exbtej7Grk3j
CrFTfmOTLoK1t9uSpbhTQ6KiOBP7d5HNO7nn/bNoTuHTCYHo/MxVKs3fqpBz7vNo
7LF2fEA9/wkEoTU9bPUedkY1BnVALt6sEVOGVSqbsfsIVGYBZq7EJLmxg8RgkNrk
VWbN1jkNcXLn+Xp2nvR1MezQfDVn3qS33TVXRwsBrCXTeNEFyRGkw6F5ook3KBzM
esHURiIthBuORLbC5asxZCVP/Wh1veggMNS4PncnEyHLdaBKZsKMBa+KoHo8OTIo
m/615OVNuMdCkEs9nAKz0k3qoMQMWZT0Ud6ZfeiRRW6z9uSutUas4IJopi5IEXCb
uV0TgPcX6RxDRg36mlgDs+WBM8TQl75zNdfEUZCWJd0P5x56kizNYTTVbYncK3+v
uvdJcBdS5c+E/f5m60Z4+VFZOQcbh3cCHcq/PzaiX2EsvsU3iZdx40fjO4GAKZ1R
BG/qAJJUVPGswT/DYZTJOOhPfgDl11elDQHLWq7tbuqVuLEK4C1fKHEhi6uNsdKS
8XOFdHpivcmueRM4d0tQ4naFAsKJxiiuASj+M2NSFBjrqRIj3Gux6iYZQAqVfzM5
eu0plGSci42j472WtjuqmNSy9t1vC8rR1wTnz0xhbmocx3HPAuwvZiQPKZAQp99c
zFVzekpqJvVbIkxrPwH+9Ws1Rk4xTbzCKfzps1mhiAbJEBtKy9kRKYk/SiV8HIz8
zY69X0avCg2JAl8hfSY9XzqSqbudtiy4o2ZI1oZ8K2+aTX4Pe8B1Pb2NgXkEYqMG
3dj1nCvXRzIaRTOURJsjOSip5yE8qdUOU68YZ4GhTWWYUgQ+zaKcViodnCbPH4eB
npyERYSl3w8E5mzR+WNR5S+zrFCSA6uKAm9M0Jd2Scb67BkSCIzAObGYvazD6rAw
oL4MpPeIvzJookuFHt2gidZ7ioBK7twQIVr5VcPSVsjeMeKnySsjZHK61vINr9kf
aH3s9qPUBVVHN5BWREdY98cNj+6ygeHsJNQLfq2HqiAUP1vhEuMfCms9euqQV4SQ
VSD9+lVYWrU6xUDMBBFgRFQRivACXGQClbfl1Z4mjB78e/be4cZPS3OuhidaM+Pd
inbBI3fBv11mFohyd0m1USv95jHi3m1ORCr6vzZXWBnUy95BfZh8V3O6FeT9phba
9SVwxAGw6LkJpSwJdt6GuyyatZ5FE0jk8TM1PWwm6v2/SSM51v3Mtt8BppUjzC8a
nIW+9a8UDpWzMFnZzQYf6VEszfER6alfeBJG889pLfAb6otlcuG0y/GR0BLp8P0+
f2Up9BbzHiCBEI0yl4iqpRBBGPTbi6LRF4cdg+kQ4WTSXIcoSpO/dMo+MkJlpUdI
9zGG4naMpAwn8b/dJ0Ha4TvYVrD8PpCHr8dUl/hw444HkerV/iisOgZUXkiCb0dg
jb9xycjzxWJ+4vqMuYKhMOMax8d8N/x8EvCikzBOqmQKe90s7tjqaHGhHN7p2VPl
s3rIEtiOpO8bJXgWTRndmGZdKu/EheH0dXJFifGAEnnpchTTDVq+MB6DYeOEYRie
G+3ugqOvVm676hSc6PMVShG+nUDyWHn9exThOuyQNQ0BJW+f4sJX32LLpQXUhXvv
6vunXmRO0+CbjntfwF9taw4/eivZ0RZ2MwI+RO0pMoIhJw3+WVXyhC6rVriiQTgg
/ndhjN0ZEpGo3GlHQIV3sq6cfRJqVjTy7BBQUqCO3cwATzq59jeb9I7i/0zUF+6t
qBl+UYByaX+RgkVpHOhp4JoY/5Fmo6qiw4zGi9Xcqc/6VYl5BmHu+tdkJGqC3v2j
v5pBRVM3lgAv3L6vEeIP444vf/tfxUF+r0MG4IBDmHN5n7SbCUYztGMvyP+RTs/q
DjHKe+0R+U+HhXMeiFAU7XAIqaiRrkpRgSmw7T6F+05eY0POEf10iXKa+Ao754W4
L6JawcqDfC99dwTZT+zkdQ9DR1b/vyl01DDJSRlkBBjhRnOsL6g/upd1TCuPdV8e
u/JTasvLB4o2lLD8vErk5roKs6+18B76Y1Tgkq9fJBLzUNcArNJtagOkyQln3ehB
SWGofwsLVNR/qMNTTUC4aRuVgEYFojDxRherGMCeo3QiG7b7a5ZztnMUo7/c5vrA
DMECq+d/uGhYuCi6RORtHYWFFG3jyuBaMbyt8356iiclgLxMbZGF1XQJHkqn7Zug
5Fy7Z+HHNb60F9c7ujaCdFs/VAXrREOmytg3JqXJlNRDFBp6+vmG9cyiDXKxgWwp
O4TyVehmxLr98Ug6PayxSFdW9foAVv/onWyASJwHP+X+wgED9qfMvxHuhl19VtS8
6nyz+GTfN7xTCovuiP5dgjM8Hl1+FukA9e20QYWAt02E+Mtc11/B0Lkjp4E7oRg8
LnsQ/f14LibSqn5IGEQDCN25cVtwphtU1V/3UIvBfFyrTzppgVmZ5CRW8DZnYs2x
j5ng87hS/1vLJTVrcqhtlYV/I6Oubr+lxsZm/BHpMibBEdvZ9RsH6FV71H/T3eZ+
O1ZG+7lFYLNYr6ofyEiVb52A8AKOOR0zyBr311t44RLQSRPX7BCXc2wHWXsMeeqh
lrMYHCcm3TM2VsXHiaPIRTwBfy5L1v/8RufzcqkFDbvKh9YZfNqBIEQal10gP7Z5
dXLJJpCGjar2q4CdsLf5cSRO1GVyYZsj0vB2zVmprdwLMOjKbuEr+UJ/piw3H3YF
xycXPZ9OvrKxBHq8ESmSrCjlOUDZzbLGajHX8x5cObKf5vXiQKm/21D9CDkk2AqP
sWELSbqA4zUoqZS+mHZxV8OiH4TTT7AvkEPXmnQ2Yh5hbFKIAAo2e/EZnXkTfO0f
ImOA355cHmsOnPOQUOLJN2znSrlmfeE4yLAlHBQRPy3pY4OzudNoLDblp202gXlZ
V7MIbI8a+Y2feMKsN5CkM8q/lnSV5Ven5FM533fHliilEkAc6HCL+RPLHXbHDF2O
l6i6OYCPClCJqLgYxUXVCek8vky+htjZDc7TCXRdwBiIsrRmAPF0deH4GYlDnvDA
ajajXsfOpikFaDhTlvzDN2ojBT0tIblH5HqMlqb3LC9shiWaGZIch4p/KdmPGFQ6
uQ3Wfc8UqW9xceKSN1MGSCt5nYUAfArXvruUwHXDYXMdB9ogt3iRaGAkX3NII0qX
O1n1/S0rmRGT9bhMTkx4FX5BgiW0d1FfCavRjyj8vINC0YqLfjbX0XLvVAbqwzld
vi4ri823ToDDvuFgZASzF0P1K90sy6jFT0S3flC2eLZdtEU+zYlewTvLTUnV/ifq
Vr3kH7fFoj0azy5yPZplqgHBC4FbOayrCORTkzb+yA8ZmBM4pr7Lu20k8EN1xuqb
y0SNMreBQLjWiQ+RklSxcJG67hU2q3rzVAwF3UJHIH++Xeg8r0ce5POhsS2YRgvb
K2N7EadgnbyS0wTZkxo06qgvQy+37uDkEWLAOoCZBik6ZHi8BljtcrmCnIreY988
udFOa7Or684YnKIBNEoXWBzAaRW1aCD76JuflaCZC34JE0GbpWHdYWxF7Jy2xwWt
YSG8nZjo5w68n1JmfkAjBnkzGfAmLENXjmnDKY9GCAxWFn8B6QonB9UyoEsyGshc
xP9In8M9mWzVv4+l9OCx0xGwNL8A27s6ueq9UMCVBGLUpyhld8IInOVcgqP//2ru
FlK10iwaPqTINOYXQqvAouKTMh0H9+hoGIDUgmvL1uYrtAgE2Bgm4G7R0GAu0Hek
G3k8QJeIGqYSnzHOQpDIEnPGcuOJfU4hS0WMRraij4b2VK2k4VIEfuwyQzXr/kZy
Zt0+yKBOuLDb/Q3raAhWDD4mxBh9ji9m4seaOchb74y1VGdkHOv4e1GCdMGrtwjZ
uNvboLCCU35lUcbzlQb5vJssSI6JjEBAg0eRDNznXZO3twOWqsRZFsg9CmtSw+6D
NWu20HIyXFHjdPnE6KvNIN+0dtxnm7m/3OkhWlYniHvpTkg1Xmbeymb0/HQwwFPI
++5ke/FaLysXAa5dh2zz4oxrg76Plg9CY/5viA9z4cBPvUIl5mkIv864cz90SnO7
ioSs6q/6YWy4MP39dXbBduc67jkaewE9iEVAtvQ9lxQSE/zOTpqiE6i8xBLr5Pg8
D6yMMyVfupRThIUsOhq018oujf0w8V40lBvrbxUXWBIqTleyp38CTQtiTw3AzIQq
AXUaQrE0K+dXSuFP7XlbGyAAunUrkwMIHPnjWw1xmrvbu5aRjWm6XVDUdkGZJ4gl
Mq7sb6mNe0PzS6WalmiFWbAyO1REefgUEKj2kVjCC9AI4+UvBP39R7o97VRimqbt
z3PYX5mOIlQ/7+NkUjjjadhM1g6HLb3RAhzXV0+z5qgWQAM1EWbv6pcz5te92hIb
eml98ULgKxEp39MFJfacL3ZDBrdnmQLXYCZURC1oOiu9uP8jHb0s8E6zxr+iY0yY
cYW87vwYC6eEdQPGve9O9V/M5YbY0Gu6TgwesOzzPgEVmuuNQ0xwp8Nx11cx5j2B
BK176/shFrSwL+eDtsTniIz/ZF9lvftzVtEvPNRzeip+RUbvri7WW+HqW2WyJNck
LX82n6LATXJbmXBSewCmOLOiqh3+oG+a1wMm5wZzXYUEmTyE5tJ2wg537YEVFFxt
wAeseag3Vh4ARPrFS9x7D4F3MKdjH2opfxN7hVbBLYRu54cYyyJRbnvHfn43FC9a
Bbca9AjweafQBbJcHHhQiNVK3aI3UpUdZTO7pupaWkGWWk2MGzx1G2Miu2IOpbZJ
DQEpnwczzXePPSTjbNNYrL0K48o/qVRolx6nylrxG4eS515yZUEzdFFUwhNdXKql
1+FZbwR9xu5wZc3IWLb7QBn0I6IJHB4QXfD6Mf6tPiNwYT+0frJg6EHWfwGvWQL0
a4iznssUIM93uOvSe+RVAP6xsnGOPuqcp7EpXuHCxrTMMEyAimhqXzaBS7vA4WHw
JgNiU+p1qQxoKMtz8NftB1jGmY/DGrlIp/dXtZC1q23WxFkP+E+L7wgMbj79HG7E
LQGWav7h+4FSsyxzhKvTvuNCPGNPPfcXt1hWai8KARIukAnU2GTwwRAU2GFCuG36
L6LUBuERAM2GrIhvMTdrNPDt/z6jWNEIrHZZ7f+BZMAYConoZbnLtUpK3vgY7pkl
0SkVNCT+wEa+YFVIHMTz3ZA5MEGKB8DJeOM+kIXZELJQnjuRgxlxC8LFzHkOER1i
DClZuZ/Cubjpgwc4KPo5Pv5T5kvkgSc/v/Isi/DiDt8R2jk7iY4wdTmK4z+LoRyY
7hX4J+RRktHHp+hpbrNRpzLn1pcE8FzoUy8QD3UKasBzWd/rF7/Btv4STU5RZYPz
ZnZ0+KKwAaOLHHGx402Cv7iJ+1fF6sA1nDQDd60qGnTVjdEeprnToWItbxEQXPtj
53/g3QwzNW6Tj5bSJmKrK34J3c/hXcCP4+INQQlw8P9pL8VAm6301xmrWOqGlQ/R
EpyWiT1wSMSt4jlcnnILk+j2/nWZXPiH1pNSIVoGzglR1mfowUmpckhEt1Be1ZQO
Rk2KD4Z9OIrSdhamLaJnfljmJ4GSXKKYXd75b8r3cGDk9rx8EfxPZzPycjzLhyc3
ZOe88M1CWmSmzazdvomSXrhEHGOqXhzM7njf/EHGEDGodJl2CrFnXWGBTjJi7xGp
nsCcTr7X3j0W8uX6OYj0JnNbLUyjaYYL5Qf1Hv9g77zexijuszPTVt+mvQSlF1A1
qrFJj9ztspF82yQT00ysOdqgAtra6+6P4jfRnR9XrY6iMez5JcAhTOHRpokRFwri
cOvL+6GlmWifnYb7e0vv1zFCqEnxQu8QKgw+u/Bt7R1KQXqWlnNSckuHLvWS0wkv
ZhPdw0k5EwnvrjpY/CHnTWFEiBS2NiqZA4ztZcSiQSWOYZf40WOqhFGygLPmRmuP
J4FZQg1yWooN9FN/HN159ZXIDQhI02mCzIJMZjEgl8EjPZEXegTDAETUDKWlbHTd
YAZZcYo+SPzXid2tFMjxraRVrhj3+sINXf5ASObkAxLdTzMJzJoBWSHiRyT5igA9
5Zzbg40ZVoJx8Ke40eQaUA1js2MWzEDjZm/s1DpgwWWNCEhyMYoKWGScRZQmI9u+
2/e5QHunTW9ofYNXztp7BPF3eKf3hRMe+MV4ZyhIIbHawzafRjY+JyMoCP4FO4QV
NzFZp6CCwsaG5R0IwT5I6RIpZT4LOcfdiYadZCit3LarotSrO7eSfvhKOmHZ527r
5s5l6YL95Q999GEQaM2k5ADBK3aXQ7mUMubTK3zyiH2Y/Du/C2IJGXLw5QSodJep
JAX0WQBzM09a/T6c+cJwIDi8h+fz0iOKcSmpz05Y1OWKIUm1O4+Mpkowfa2YuknH
GklQKHw1yWbYtv1dhbaIC4Rl7wfyD8diR6E4qhhI62ZaK7oPFkQIJZeLxiQQS0bN
0A/HKJaJa2V8NceTKxvqhMChHrliwbXjGPfBJ9hRPazB8DItaue+hBzOhKP0Idam
oc55ixp4WDtaTrybfrdVrlLArX69H3fn1day7ATOi391MeANJnPOGT0eN9fXXIXP
7QCFcP4ykEPCX+xT4KrgL3Dm5v1qeb9rWCj3TM6zTH9DiHyUkjXXczPEU5iuan+h
lCbM039pRWh7Uug8SuyQRJdT/j/lGF5ktvL4WMpr73e3Wn16zJckGVoVtBEOFoqD
jtQSDHqMNFiln2qSPac6HXHH/pIPfXzJPPZDmU/LcrkB0KRYioU1fkUijB9Fk3Am
GisIk79FpXte3cf9oRf/zYQnmU3aSFJImAXj79ko9VQRaVSVNllyEBBdJ3KXfhpj
u0oecUbnQu6lSTt0ZMf0bgt7CzXT/6Ds6oMRQgt1EFNx4XQlK4CRNFg0xktG2zXI
mCCYJpb132DHulzSfFNALh+Wuy0Wu7rjS9pXgfVKBBaDPl65UmkOE6YN3FjgIXrI
DIlXWc357iliEh/t2P4VfFKnnGWem3BIpdkc4szt5X7lQT/b0Z6P70PB09LH8gbc
FiXWhvaO2u0v+aBwocRzLDR/BorV9ft0VoIVe2qaj+uVzfP6BmIA7vFYsKZbu7nE
TlodkWCiy6A9uu/du2zU8KUVPnyNekjY/4gh+YoV6u3v5+xfVl3az7W77nr+Nw5d
UE2HXD8I5iJ5l7wakRusD3V5GKwTspxe2bKYKFhl5zj8+drZaTSzk4+Jj4ZYN16i
syJc0GCDyxZfQl5hXSq+kTCB9oK8RyHR15dCEPR9n4yEWdjoqoKM6QkYkxjU3EmK
1+GIeGBAnFY9iXq/9he3yCj4A3diwsm6/4Vl8QRC1vFtMOuAydgr04FvIQf0zxvg
5yabdURslrjpXy28d89Q4mjHUvy76xaZHkWffdRHMHS2c4T+DvJPiIMg/F9J3ucm
bQawAOvg5VhYEsCiO42qx9AzJJ10C1Iol+vXLWPch/C4ZUCSaHQ0I/OuFtSHv5mT
mBH57kBhYojy6M+foZxLN2qldN1C6PE5Ynv5XmBOI+FWvwChzHc/Eber/t9CLrBv
cW3iN/DlvJeg29MUln2o8WqSecvB4jrrMaPTeS/FvtXd4a0EDNQ3QHM7CKhRPOFM
9shOTogDkK34YEHPPO2evUBEtCA4Li7QFG+q99BfTd7QrSGg0kl5avgfedJ91ovJ
zZPR+IlkE6ASaYhEXEKLgPi6TwCUvniwgk9FtKwkIVGQFwDlJ3B87PcFOL05qznJ
sCUAsqwU19VLyE3LFuc7y3Op0EEyUnWIGgcsKu/zkqzYwZS4S9IgA35wMWBV+FQp
+WZ0OWZRJ1rX1Qsu0VhsSVEebgB/YbdNtOH/hX1knoQq9uy982Oxi3D2ArXMZ80L
xWlEU3Vmyg/A3SUAIlCr3XHXe1NxgEsaSZf14gYDwjeQ/QTfuGVCisRZTRf4Jz1f
t6Yghr6No4W3ddCyJzF0/lGjxIonk7UXV+mBYIxO8IjIdO4bdtdpF8FwJp8woc8P
pG2V82KvdTYCuzltakdAt383AxtrTAWCc2kNgde639/bMdZkoAuTrdygUcEU36Xz
0TMxuPupRmjb9M3sqK4pOP5hWd3iXq1XaP7UaKEvifJKADWlWu3xlY2zjPoN/s7z
8sakfqSQtXYDIfaVs+VnmDrWGYgky/WmJV1+cU2HAvIZ2EgAH/B61KM2D3x67zOJ
RZqkL2ezFAFD1Ko+1gj4J12eYsY7D+XVTDN5xDzfMEdsSSaxBsDIlMmAQ1sW3C8x
1UTWA64of8EvdzUppxv8kWowYZh/wA3KBZpe6Hi+zZKyIjzn4Sj8quBGzst5ll5p
RlRdOBsYwnJNRn2NoMITP+6/yBVJaNdz5UpkhtOxqxcHJVn97SfAA9z4o8hL/H25
eb2voJndTrY9UGpaemyOTFQeeH6rVXw3sw3GxnuTlc1QW68QbZv2UCDkLqBCiGTt
W0hzT2Z6dwgxJ13FCnepzdXRS65pneMPrZK1sTZbOBOqcMvyF6YDqUYTJfeVlRrN
5kH+0zek2mYA9v9XJXzvlX3PmqrIMxP6WRml+3G2CaeI3S5Rm8Gzv4m06VfRz5T+
Ku9l22vJ79jFd9bbQ7s8gkalW7ETkiAxMgCCznzlTGmux7jwtpfSYR7nNLYQ2iSR
STEt2vQXpJbpXO/TIPNOMJkgJLacw0VT1i1sQDzAEvprSyzl05TtOCAVJjWlX5Ie
luxMjiJAKIv57Cz+IicIRaKpw4LHGLbN+9/z3p2+PhZm9sR5CbkafY4ltx45B3zR
TOAV8eH0NFUxXB6ON10YAuTbyq6m761aZSTaZD9S2Cf6C0QQENLgqL+wy05bPOJ3
dnZVwPJoTJ12Dtb0HUk3W1iXpIyIryvu9PViGXF1E/nh3FdELpYeo1uJorPMSMnw
/rCr4b7haVCX3pzcKjNegKaQiNalIG7egOWbvrP5KDsPutQxpIAj6SVmELsolMWp
6hbZOrI9EBdDKZVjC2m1JTGJI08/dqFNig9FNxW1ydev8Pnio2wtkZ2B1+FTjNq1
Wh6hIb4R5vKBMravaop4l+Szd/eLcdhQm7e5OcomnyGs9yDNJSvlTAj2CNby2JDT
CJvwjQZBu3UiKvwFktyHSP2UBQroDfJANf26FljYRf1iydHzqpD2rF44PD68whsn
7KDZGrs7rNNy1ih7EALERbE1y5P5nQy6LqeKRoiT5uuTckmE157xEyMvQNPRkbae
717edAK3TmkGf5/dsJgddNQB61YIkespY+YCyUGgF5dofhCNxaMTM9nSMfVYUKE4
fwDSGFbKya5ye/WNfKjVGKPPID4vNkS6nMMJyjU9P9wsNHVC6zT+Rvd0HGXEsIv+
0v9zxjDFrHJRVaS6rSCzdBeifqFeGw9F9BZRy+G+iUhdwIBSq8ejJv8rk6x2G7H3
dcyr/BL9XaRgN0ErIRwl398TP5IenO8PjjNoew4Ir5i25zInS+cbiBGA+F4dqL79
OWHAR5BB61FcIpGbeOA43Y9GyjJlRKRw8AoWxcwfCB0fC886hxm0chixPVDtn5aF
cJZkLPFXsskvE9tYwUXa4NYChL7HEy+DiQvO/n0wvPTD/PQtWNgBZthVQBEKE5Wk
H+aCo7B3IQQiP8KET9gT3JJBOY69RUpB/Qbe5eXrauxvPC9fBepYwwlQKQFBW7wE
YL3UyIWDP4Nd1ugJpa4R7rpBWfDWGmJWxm0XGsMuBjjRPO3q4gghapVtjM5JyP17
7LxaWk0Yw/M/anP1pXpLjvDjOzhJ/o7X4+apMUVAWOsbwyhLwRlR2NXE/FHve7vM
7xHcGALKidzXrrVZg+g17Ok0tqt7NnYs2NQtA/t20zJI7MWGsXq9fra12Iff/n5e
7yt/znMzq8cWFxB4oE2nc8kNNGWMAmJLHG5K4BJWrehnMsj/vXw/X3OB4veLCFaS
FHHMGfnDCnwyZeFswihnPUkO8cT4VMtchItJ6Hmxelv01CxibQfYUPPH4w4fPTvf
xj+TFu9OQNQzvjxAf9gsxh7nPcg15nev203qcHnpXM6pqLQdmVnx9Nae23dfjR0t
Dg9k6I97ydDZ00UOPO/O4x+trrdrFBoDLQwsg3pRWPrvdBHgUgGi+hG36gpH/KIU
AYxS+QGLzVgVeGNt/UtdmwBdzm+pDOqsLq9faq9HzvrEENtTmA3CmwCVxDy7QsHB
jYquKsNhNm2nwtNe6ISPj8T7kVsVXTlaK46BhSbdP2zhgI1wlAWFrWjeOoE87SeO
qpbXQO0TGQfXkD1+e8fhAPsrLInHI/6Zagof3hdaCUEDgJDkaT7jT4HknIFGnChI
a3ZV1TjRZRJpyGusaelNLY8jK65hzBhyuBwPikR9Y+Z1p/jI9zdtCQlYG+CE3tmA
KQOyq1VbI6eLYPOsULUkoKpR4yxsvXJVd2rlUUlWljoP1GN0WXwoE9K9/rKeodFd
o22kvA5NEAqHZ9lY7wfIzChsw35Km/HftCtNFK+hXKJ6rBP/7fZoVzPIyxcFPVw5
xBaKmWkbAW2UVVwWxz1VgLtcenFDQpHU6SnxKw9Taz02zs7QfpiEnh9fGzsZXYxW
ghaGA+xpcmPGeyUcTD1fDMyaAN61PzMys9sVZRjQjR5dBepIp/jZuqbb9lUOVRYC
RVt1D32HqUrQgrgPRENovOxDD8CwQ1SOt8elh3SZ9Z/zDPwSH8AEocS6nzELuCT1
zPLGHh6QgabtOELzkBRoqsZ6Du1PrT6JNIfk28hvpK2YOwcrt4UamT1XC9TEZ1f1
xWs20W3vF8+f01Qj/7lwbt9dXV8zZmrEx6uXTfNkQu3Mc2R32Kz/hr9wlnjvJLp1
HMflqt/rz+ASuFZQLNlI+psvRO0t0pw5biafGZsIGkyBf5WYakrsry52m2M/RIjq
2p40mpaFFuUgvqswqqbQR4qhjraQeKV7lPnjVAD2EScEq8v/FzVbc63uM2+VAN9S
ZoGJJ0Dacb8mkjVW8negFeJUnnVnB2nWMXfTFeT9sLrFTWv74zw+TGVUutQ2i6SU
WgP/c2GhUTRHRBXU39CMwqz2CY54X6rdfjEMUZQ95beuCsa3quaeUaFG/87/KD0K
OhRbPcHOYmDu6NfC8MVqMI8fQjwx6Xv7rw9cg//6if6uVkv4fkgo4fD5Mh/9nuy1
hczdhjR90NJaQXqYtdVJ+taAZMFl070bhj0Vi8nin2Ao4UbWTrxtYP1TARDfELjW
0XfdiFRI52aWgBdj2958ccLUzJRzYJnDdkMyhQpMQPOFnvALMdYIaE+m8SqQYWtX
+kq5rE1CSh2z81HThTT8O1OJ44DUA5AV2ED7RRYCQow9hrECaZY9Q8ozYXcGvRui
2ErW3rb1LXbKQeI/2YV4nTLEKMXPP+SurW13SKQ5GT2WVWMJH98uGcJGZV6faoWu
cNqg5pY8g71FdSVVk9AyiaDkwvra5YHUpUiy2pT9UuXQwTNf7P9ca+vBbYEzMikh
Fw9yZf+0LQD1ukzY9hBigen3pSGpa+hD8+Yh+iFINDWvN9TyWs43CoMiCeBvwEVM
QU4tTKsoNwgf1ZutjASD2KcVh8kxOud7F9jZEpjd8qtjxbzUNx+ILoJtYtG9jd54
/QEWrHdII9Pe7BPfk7wr0Qf53lYcKj0BIYcrBg0TTA8gGX0dhHegZrx3a9Tph+pE
jhCwV05UPGk6ErAnU9j0LjYsgX4ilpEOL+Rz5KZmrfsneuhR1kEaKsqiwiZpmHst
V+YUoBxWJsIj5gl505b5ckn6FP0JYtLcpnhrnISgln+dAR9R5B2IoB/l8A9kWS30
fmDC4OffQbF8d+saCD8twO7DpZmssGWn5yiijF32p8M2lX9tl/1kbJhcudokaRBC
HUJ8ZZkjM62mHLObjqb/cAaI6DckO1NVLfHSzMsiZ/M7J3WaK7BxKRlSWHexKDHs
llJekmUAgaOGbz/ACbdTRhgfB/7AnfDaSt44VXYkGgUx6LfzI+cCwJcrcKnAqIH2
6VLr4JZrdAX1/8seSM1fv0QPIq4SU+377e2R6OUb9UPM6ZJ74vnSNv+rgsJQIvqQ
FRkfuVkwwK52TsEuljaWqrLwsU/25TIGoOK4eoFNDDwQpO6+ALH8mXHQrUmP8CcD
xQGApHn3f5+q07GKjwdb6SXxgoGvGYnBI/wJaqNBUWYzP44ky3KV21Xzqf+VlkEy
D9qTWFh4ksjJPJhbeoIELnbqfhlr4otzy528nB4eV4VHLNJOYK0dIbKdg3uFbxAb
0jzugaz1IaFUQxoqiaOtVd5w0tKetBqAUxmX6c23qD/aP0OedC8tetNO4iUxsfWw
MzUuy/Yf23zzEWpMiMJ2oZhYUGZo1JmilyLV0msq/KohpHm/fhdyEYRFxZ7XTCpC
Vhnlg9Lj4QYdR5S9khFPX68LIXxnxJrne3kPy1dkWKYFCdertEfhWRNhTAgL2UfZ
sGCUAL3LJcZWzC6pMoR7Osyaxx4tQjJhKqQ5BjDEQsiXtpucBQXo4petAYVi9Pj2
0/u39iUiUBrqGmIeSG2K3xxZBKUXnq7FPyOk+bgFaZgxv2Mz11DUVgRaH6Kpsbpw
B4FguFhIiY7vrILtVrJpcSL1Go/hxh+sRLGVT0sy8hChhIRbtrNhP6NHscqxOonk
eVFDfocX7ZcI0Cf56ELzDSgHO7/28mCUr21PYKXli9l68HH3plIGQkKuj9bJwwf9
6rzD/+tVd4+4mVGPnJoq/ZfjnqKfujSPR/lxdsAI785VABPkNuUD7mRrjFcGnus+
PPqSHQZiLtYa9yFrV3WlTVJ4ZdMOZjeDpK0kzofr93zMy6sNKyOvxk9dbW4EP3ws
iEdCjEe+05Kcyir2kuchrsZuOMCrXtg+hTNzZ3mD/sjDpVHo7yOCYteUdBvXPzUH
OvtK4sl0St3Gx5w/sDMFAuvRI/6AwkT+5edMfmdw+jzWkGJ3S0vujyF2x3Egtvb3
B1jcDbSFYQoH50hJZPvih8PL7tfJIBOGMD5JTyylgzEljlamEMsn+Rqxee/O/fb/
9uPGT5E2aGc/mvmI2He97sTgt3fHCp4rjkucQh00hT3XqZy/A8lyzJ8lSjfXyaPh
BagseXEHg5sNY/ke9F4FXkgHR6J8H/VqWIkMYA8GnUWzyzLrTrdQNjSkE6OWFpE5
KGkGiz1GSiqi2b1gFB/Or7py+BJBRUeEt1XdEVOCYxAHxBVBSWdlocczuRfwPn4m
bcgOK8lidFaXqAd/AJ+U0OZt26Y5lbpzSqKbICSD9QnsnOd+hWnVe++1PrHpxm83
SKVJB52OxKPefPNZ/OC7utNwS1vwxM5d/fsI+7lkwDhbrylnNLozGgsOMF8MkBjw
+c4XkcugesXmjRlJc5G1RjlfFAYx1kzArJ8oP3R2pCBgQVhT6KDrjeAcACXVrrVr
Ah12VGiXS+UqDHtRQf2ffzUDNJ/9SUBZVZVjlwzxxg1tj/DVJZoF5vizCX7iSbA0
wboaK9UXbA/tH51mLiAn9gwZGWyN/isoi+uHzHmwz33lT1FgqLsDHYmdBcNjzw10
lR6CL8mSRmaEXTQO3G5fQqFQMzPabz6sB2yCCZwgBqsc56CuA6/82AyVh8QIKr5n
J1/y1HesSRJi6c2xuxp924yxxiC93d5IkysipKOFR3Xt/l0lAZ5lRjpnXYUXg6NO
isjUPQVRA+g38PID1uNOAr6ZUQBlGStjI4kojLYgj/Dqy54L2rvqVrl0WWnFGecm
r1D3ba4RlQ/sNL+JNkGONXzo06fQk2GhusloB1x730dRbVwgoha6+Zrl7AWnHQrM
HK15qnzVZqL9p1CXABF3Efykzc7skVgL0/MBbWT5OpN5Sxk0goDyhXs5fp7wSW9z
EUp1tpuNidqXImrEV2mY8cdtVfeUU+Rw5a4asColFjIi1b5KUwFCAdwL8cKwMOre
rOhKIrd2ExlLzHfUdUCzkwszNOBoSoVb6Ldm6FAkFgNiIyAscQcdRt4h7tJ2/HtR
rn8L2NbdNxTiBKoav3pu3hyANsRVXYrUZNux8lzCjMhm4ldHi6kJbvkBSYH9jca2
uut5YL1dT9uXxB4r7I7ddc0nnCSCOchDzhngMJi9/qjPn+9b6/TEQAUz52Kf8mGr
mY+nvc7r+j8/n4c3uwzDEhFmj4KpPtFwIPaqMUd5KeQDAY0Y8p86a/NIrDtekOSW
26eISA2A7UOH0kxi5KWvDFscCty7K4W3SopQMPQqG8FlVzjaS63DKm1tHuzGDOQR
m2wJd0QzcpNg7HMD0fIqFBQd0IsnhuagO8jKYIqBEPdRijkdA8FvG+LXRZPQMOCW
Ub/EPB7pnqSTIJ91VivojOOHCfaiIs4pW+CYlOZLW0a9JHwAdJJ6G//IErKKLzqa
0CkhiBmPuozMNmLQa5cSizMxXCRfMPPhhHq1Ieys4caSOMjrHTXyG8xWtZvBQFlD
0D0zEbWtzz3Gb/4WuelPXJxqsUCRTeUtGmg8QdLYjsTmPT0apH8lxKhLoNswz0UN
b1QlfIbNgvU8qu39dP5W3pfjgq8yy/GCYmVxBA/oD2nBUd3z06P9/+vd6sleHOtq
YdDW8HqmyaY+tsDISB2ar8IrC5RQaXG9QBTIlHNj6bT+h3o5yBVg8LKMv/vjocfR
dXf/5WwkkR+T875uhu0lf08hdmr8tjazSSZoEetKxKRW0LghYt5N2NKs6AoDM676
FXMfQF8C9MLxpfBRpOF6IFXDdXvXBOJ7l+nCLwDOLCbH2heR1GCxHuYBIc/HvHje
A6BMtsee7QnAXX0jt7rd0qbN8E8Cq02ta9jUEpKumrmWEjY0tTkBm6ZsC0EhZSuo
s9w2iL6USISIytzO1yBQFSFfjFgkmEP41heMdE2FRfNUqfTdUk/VdGX8GwKsrzhB
4bvkZ4ZwtfZhqvO2pzOcMMYIpgHRwfjLUDFoHYQFosMgbGq8G679vETbFeOq5pj/
TolyZ+QYe2HUeuf6SS3KF/Q1Hs8/St4pX7Wt6XqarmLeI6VJNprsuxJ+Joc2gnIs
zSmI+zwJ5spyFJbpSTUuX048ZeBgtu7Xezhq6M+LjYSfu01Uy3KpY8rz9Qtzkd/0
cub2oHi6TFCrsOj9usoyxu6ILwHU6kbVqRCg2N7VgbI4TjGefgDR6qwRIw0Sj0fU
CUiu6tD50RPmU6h79m1AlyaxJ3C1nAVSINZPZQ84Bm+0Xd+PcFktHfw3YUFGg7Qo
eA4AfO8xaCeR9Op+2QAngt5fzW0Mpc+hN8I3tX/rOWjCctvpb3vXVpUpKcsMq53a
U0kKr6/4xt/z55jJWFOmq26K+gIWp5IEzjhE7kAERbjq7mM/2Ki+def2c06dwXyJ
0Z6YmFQtBX9u1kVBOQUEyRhjSyadEdrkepw/TtuuBfSV7EVCoFqh5pWvcaHkWQZs
5QR0o7yHJW2vQkWr9hX5HQuFhFDLqnVfIfMSDjsoPszNZ26CoJrfRM1ER4e0e10k
w8mhMg410zw2U2Yo5xks+KQkVw5/e1OKF6cmcQq2/E7RlOO0NOQgZeRhv5zKj2qW
8YQuthpUCd0cjy7JKfUph8PGIe7/mD0VG5jsvHqR1M2t1QpN081y7CsXhx8oDGqc
lwWtmaciiqsnPuFQf30rlHTEAbV83SIGKQCX+Kk2WvXPfwoJSO/yGnsarPolpQCp
jfUEUnU9h7ItbHiON5RN6KiwFsmV4zjUnA2IEO7DIiZFu+hhy8vNyAx4ZhnubJdI
uAVbN/hR09zvHsvQh8c5Ig1uk5xXi8yrQt6/vGZP8E4GPGQz9rnrgdnqEh3E28Kh
nHbk8xd+3MGyInNRDsrknRFML7YTiOCG5q1tJUKWchGkXZJ44M64y7z+ScTUKZVc
wBTOLhhE7KMvojatoQUyf9RSeYMxpmgfs0wdUxmJ37k0/xa4uJecArxn0m4kalMe
GMZEQaiqJ45pGOteA5CB0nGyQ5one8IJeP7ybPKDVB3iAVmD08v7gimjXfMeVQQ1
kHTM7PtqCa5NqOHqQkJk46GARzUBpXxhdxF/DMQGseAy7ebJO6k59BIcwshLXs17
wh0aq17rbhh+1KvbeU7dspby6BUnxr7StEy9Bi5q3nxHWGKo1upHuXI2gdyWTTLx
grlXFL3qG7TWjuStVVY706pMYEsBtjM6UjrpCPchZmozZy5Snn5p4qOQMylNdIWM
e5eVFhI0ZzMClo4Z6Au7rnzF7R7LOTO4Mj0wRHWwO0VR3ZvM/CJjHF3I0Y5S/X+Y
o802BdBLtp0xpSa/ylocpBwHb5svvV5JjaKgjTVcg7semiW1bteo1UjoTQkmkV+G
fBZJsQB53p0i5d1YiaaxAQcq0JoyEl135+1qRJr8JfjlhpkJrXEq6RhiGDXnPMBG
bPzAO7WU5Jxm/8U/ca174x0ZL94UBQ7jxGgZMVVp9EmQTcYzxqqOIfCfnEkCph/p
OuvomUj77kVL4GPQCUoGKPOgdO1tvVXHbZC71TLJwUx8eXtJ+N2syg33u6eoFq8V
yl/OpJiI0msZwTyx5F2YCONk0bzLP0H2J3uqJXELeEFZkCYxYpmStMQs1jj+N9KX
dpWt0yj3LMMQrLeBeNC4iwu5jtlt6NrPi/l9XHzpNCMWPY/xzWqJLeWPxkgRHhHH
695s1LWO1EtZBAueoMZZ0FoZHh6jiZuT0hLbtkT9rH4YP3nEX4dRzomOU2wrsK5J
LAob8wB/oPNN3L636hJLEZNxsmnK0FT0J/9davQB2YAYgGfaa0npCWsBTQK/qg4W
2EqrOfN3qA4+5i2VBQ5Wzl79UcLief3ZYbIXKRnhpsHvuOsv/lIIAGw7Eih2WTKi
NVh+3AqyOcuNpLPrx28uvl14VmBSp1hh+3RLDnqT3lxW/JTEa6NZqPTd8nZX/gFZ
pfq2kYgWJM1+FjE+WD2lmnnyuAWfuSRDrtYaDp9LXqzpI1KWsY+jdFG7pBElIwON
1xvFy1jKR/Psr6W9cZxVdhxMp1hJuGn2wcsaApflswVXH4q6BdiEizO0G7Qpc1YD
Bx44l87URpz7fSBq8UWWIID7ov2yCiaA1LLtxKhJQftstdkquA9FABYweGqVIW6J
noqEAFODtv7dT9ne/ykMPtUFnLk1YXWhVSpmlrD7AKXKqURBOD/ET4HEW2kUzGyx
4IKJ99NPGtNOj6p0OI4qhY0A9onrR4pJOQx/ZcxDBBGLi9Hk5iEpw1/Sw5PjknjZ
seBEbAY276PvG3Or/rcQYboUVSzJ+ojbZdelgLzpJTI=
`protect END_PROTECTED
