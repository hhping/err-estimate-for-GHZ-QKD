`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sxvh8twhT9IDIc7m8RQ+0W1hltPiwq0AyZOIST27S2vYAIihKnQwGHH93zmDBZCB
c36byCzR2m3tHWB47i2/AzulZdswV81I1Z03mvzSYZng93Y41qx51SfoFAIUg3De
KVCOfy2ngWQHXKkfwQmnz/JX6BgzIGNe6sodE5DCVf4tNLpn8CrfXffKOCc571yg
LdtIj3WelRdGmxdPxxxF3hich4dGNhetIC3VXrVJU30Nn6Ip11RwvwLtzVvQJW66
tj9EOKV8lZUtKHiU9V68rBznGGprxRhIAiKQi5wjakCRZnIWeCQaQcGFcRcfNjO4
wfyR4RSTJACpcAzvp801YQ85KK04ATRF3sJVVBOsut+zhCC+KeUKGavgWCOHbpL9
3rlHjEBNaoELwEs3Lt1bFjWvBN/4qnDdQz2SXjPGR7Y=
`protect END_PROTECTED
