`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y7dKPUEP9/vSrC3LdavjcOdLQRonasJKD39EmZJIpUHR9lRiifeXYsgO3A5OYqzA
N21lbZksnRqWnVzZxzTxOUEm5ORBYr2I3OeyCp1QKPa/LR3LaP2sFywWKnZuUqWK
Uwf3MtWuTUa5IZ1I7zi3nOvOfmmLqjCf9/Tj0oozoBCeanI6HpzP+9GWuaXQcgP3
Su16qTpZWQiXa8GcImWx1H6Lg8UASSMBriiLkS60Y3VQolkJ88byGoRWzoCu5qJR
nomBzyK7D40+Q61wHtfgKZ1fB7COD1/18z7FRdLlYC4oAILsw4wyF5Ge85Gq6Ygf
nDTSEnInqjki57miqjMmgOP7yZ7FCktt6yPbDeL4etqni1rpqsfovAaKnWxbTixL
LhKoKCj2YXPI7TcbNyb1EPVI10Wn6tA2JM6C1sMLczo07Oy5ZHTii5qecO6gN1M5
hz+rF7iYssZ5z7JS75ReIfkfzpVl5BaCRIA5DN2RAzXagUfGb8I8wcKoQyWufSt3
PQy/KQqE8Od19r2IxN+vqLLHxLFRC/KurIZXYeSvHmjC0DERXfQ5vZCwoEU+WVq/
MSh6KSkDx6Ytlca1jVNyOsY0q4Phs8+Rv09L22InM8RfhSI6zAlt7Hkhjc0oeNbF
vMwH/XziKBIB2w5E8u0NJqdahYMDP0e7MYZF1E7Jnk66/XiLbl6XVcp7AqfH6ILg
qjlwaENoiXVKT/Ryhr6oYUKvNK1UClcbc3UqS73gieNDZb/e/5zHHLwr+ozWpTkr
h8Kwm/Li/cvzLBRaulpaByKiWnPNQVb6uMxFEzCmXc2Ej/fRyJq7Mr9e6JgM7+jL
xpoNRkTXPEQfIC3z07Izbh1aC8DjTdZfz2EB4Gkf9qlDJFqo3drZesn2owQSZCCh
khkiW3iSfQAbR5XLwHULxACIMpoZRT8LRnx5zOhketoUOA7HZ3smoXFIVpqmyfxn
JH3/QhIuzcrU7HYQX8tNv7Bpye4QnJeLLqHvVCt2R6fRtcNge8ttehoDlSKgQzwI
Xlxiu8Syo+03gw8wfj0Di6B9aNd2JGtaSFG/BPe5lSI+z6V8QUW9VU7HBUoaZwZn
OlGZ9EHr87Brpu58O6GDcwiO5t0DExCuUbdJ68lmseVZZPN1gJIHDwARJfLqNBHj
hjNL87KmJUmPsmQvABkJuwB+IN9wK4bbNy+gMWdHi3dfo+pRFriUnIwWM1cRsrwt
l6FmdJAe4vM5Ox/WwJtyQepWYnNJ1ReQ5JVmyTzqmPTtQ+A9+83UebYZXr9fIQTy
S8YfR8C7/dT22hO1+HoSxMMsR1m7WA157U0bR11PCGU0Rp6iuxwGrJkkXZxU3etN
odI+1rJH6SmfS25RJk82UzpZdf43aWkKeJRurhKG++DQo3hZpnsqycBjN15yrCbZ
zkpCtksJ7oqgCB1EDQ06Xo+d4jUbfkwT9gcZyPQEuv7IMz73o/dyyUy4DAu+Syef
EQakidu89NATAmC7bP0mIYy5tcN9dot6mVMm6D7Virw=
`protect END_PROTECTED
