`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1NvsWVzDz1nWRxrP7Bk1i416ok7RoBleMjHqENeecIbBRGiMESYz8pr3hzMYpW7j
LjxhvQ7vwSdHRkFj3WgX2bdJ73Aw7KCH4crghI/sPdW04+g1/nBVf88dpBQCjpK6
4SZM6x7gM0dx5KpoK5OnMwF+UTAmsTQCDCvNALdGRJv/gH48WgKVKUQwsj6u2ksY
W0lZLdfxYl+utoXi3bAO8oSlGZ9imJJWqm3i08HKz6q2I/e+msZo+7SkYpzZ31Q/
nVz/ZEBCqrFYkTDh4HqVcsOKvhMFjY5HNJBDJNOEdyzXHxD0Du34ryMDr/9c0UWl
yjy3EyxAw3a8joK19Z1CDdy/UlMl29Uj6UZQ4wgO30Z/Cq+TE+mw1oFXhO9wyCzR
SfqvLhc3ED0MiGxF48mi/zImIYIAQ1INSefI2GB2/VH8RRW38VhlGoSWrPCIknAd
RUr7F8P6avnsh2I5SER+TizYawlJtQxySR+ORP6c8eVu13bt1kj0h//Glf1lBsCR
Lay4NUcBSibVW4SW3ThiQguHFjg699fUl5Ia3wWZMaGOtLQACnByGjgsUKTE3lpy
pDucmItfdv/MADGC6pIglSp/wa82xav7LVLD0QiOhDFp231Y04Iw/8O/+cKFJo37
gQPRSwMi8zKpcOahIVbcLOUY0xMbq7Xq1Bptyk0uSvl6nDFDknUgCdHpP0TDJUpx
xrVpOY9qT/SmNF/bC6IuxBV4duHNt5lxvLw3Jzww95jUAm116qAWTKALD2m5/QEr
SRtnGMAlGxw6liT3GNY/TT5NT54JH3Ue/TBHZgKH7K/wHdXADhU6rxQ9H5V+FRcD
/UNPUClQY0Q8BzDpzl67lpxJqPkLEY0HZAdxGS5G5lYPjp1TByn42LrFML2YZ3vP
CbnTABXXTZFU3HaLlXUjVkCtwEKBU3a/3RtD8A6GdqxsuSgHrYrTQ57tUODphF6Y
7+DfW5VMJRjxQkHiDnz9UuMOoHpDaUQeLVtTKcL376zhRcaTmn9+g/C04zHoNeMf
+dFcMzIxK/Qpw/2IXMt5Tk+DalxXkjWctjrAHQDFC9TyzDgRR5y099dMuH3gF67g
/bvN6R3UfWSFSqjpy+v/Ifs4SlyMaqbpo+BKfdeSeHB2GHzX6SH69GeYleyqSiwE
GFmk8mW5HfjKbCKn/OTasgEDjW9Rr8EUogxxk7HUAWCax+i33nACcG+PGRBXFA2R
BIMldPjAD8B1TL1+r8ti4u+TuOTIRr59z5HAQ0TO0oCXtmqYT1cVpDAwjQtCjGWw
i7ZXcK85ErDXK0ABjALxJg==
`protect END_PROTECTED
