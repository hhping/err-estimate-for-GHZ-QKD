`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vYorbKYbr2ssJ1TBaaRukLF8Q04XGVZziV+YJ8hP/mxtkJC25IYFf5FJWsanz4O/
zOfTtB7HB9Bfmv6BMB2mwyINmAElpVKtZKnehz54/hy2qXlAWN/xNrWjBb/Tr65j
lkdIjSm9OkoOXYn73ZdHlPjona1Jq1caCEcNVaPMhxk4pKUVPiw6tg0caOzyNo/O
sbPmi1Ei0Nqao64GI5owbtRslKUSpWwR0O/E6eYovDinbpIiTS2yTr3ouNBcXdz0
mhoYdte2L2qUyl4+/NtJoqR39aWCC+xiSVk4zi4y2wOPC+epJHtZu/j2Nydmi/fQ
6lLbqVbyHYNKFb8ZVMZiOnmFn7o0o6LPYCvhmYcyuRe94oSU4goPyKtf5/MGWx0s
zh0seiaUSWCg1ZfNNhBgAuPpEgpNRXqFk3uCCFxqA5crPnTmOGJ8A7F24qDgdZEa
8Z1+BdBGcJs9ixag4WzySTGJEBgT0g88ImhRjqTsk8kmitLnFHjPSzqt0W3iYJHV
RF09tNdlAUfHa97/2jy1hMAbOvTNv02fi17c5SamSC3aaOrr8ww6Y0c9Eip+FwWS
Xw6kDL2nKEw1gngUyFU+cEuf/YsLpMQzc0mduvDoiLW4k0QXAWQVL7yiTt78zaG6
AC8DTgZTArP7sqw8UE/m8QGnV4FWKHYgxVr0XnMTmH8yIbpsScwXPj5IlIZ/L8CQ
u5KysdiLx5qQpJHl7cRzvUYh+9aEMz/Uan1QqpN+gJebchSjUSiyxSU3j8pCnIF3
oeEOW3of3appABEDQGdbmJV51YLUuPL8hItx/7JLuIO5w6xnIZ8FpBzuQV9fvBf1
MIe6u7GqStcJB+R8VOLq+AnJiqF97hhpw/7KoVFnrNNbEZOuymt//gd6bQLiw2rI
vWXEnIaifwyJIbrk/bGhvPfDkth7jUNDt2U8Vqw7jMfDFapZT6B49XtWWVP6TDp1
6kYZ+Fdo1YPXApN9n1zL/5MOqTB7iKnBTTpWSKcvfpAEcTJFVFUQwN0RvqCW/GnL
gscdKyi+OXQGC2GWZDuTjJcwp8/tL+L7pxXDAfVmn1sJU9SgMbnfDixrLjA7sxef
w56ih5zpxi0rRb6/SZ9PDHArvNh9Fs78DKtf5gcx0A/xrknFbfirZV0ab+VjIf8S
1pna6n292sZhl5aQnjVht5yLwkriiimejRBmiRQibIsE0p7HHIMqw4dH/tSsal4b
kR+RXK+zVeAN9bGmDej1wpRIsPGQYdbNP8S0Vbbaq0xMST+gBhWDOQcNJ2fFdpfu
TkJ2YtKohxgBz1pMtz6HmqoIBNkFNLZWQkwTMmOfbwV73m0lnfI4x04Kn6v+Cfmv
qbmi2gNzsa9hKQVFZPTmRLsXSGqXjTk5PbzI02rYNIVJoHX8nUBBPbPP3RDW9rcP
2PK0oCjSktm5Phj9MHaWpieehODi4nXMPaiIYhw/tpsWA0dGQZy9t+/3lVCVjiMc
IJ2rpUgOb+2LPN7TDXefG3eFT+XXYBG7N2h/QCbFDBI=
`protect END_PROTECTED
