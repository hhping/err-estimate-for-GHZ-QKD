`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o2jEV8J2Sru8w7Psn/eIQSgcFeFrKYPtjNhazifAF8KA2U0oZ1epZxHprYm94i1g
+YgO52+4lP/3mXnx9Rv2Bu40lFrl8Glv3+SifXJjju5xIETC5GX8+9cGO5Ltf4Nr
1NcXqfmZS01srocp7uT2XbsowFQM6/Y2bpQp4FD9fwE+zJuP+zz/zSDcr90XRPTZ
T5eExfo1Y2auiJ3H//VhBnF+YFrZEr/hoWoFrbBcQIo3LcLxoRXQ0CcQLPZTqWxD
8UE4i7QgYyKWpNvuFGaiGf8TDOEkeesacWLV1G7y7bEzcGR0jnvlP5VvdpTIK8L6
MVtCC7hlk+JqC5TOIGuQADIyOtPWSc99CPIRW/c/WtPD848kTCVoJ/MMlnwGVWue
3hEQaeoyWppJryAbrO0u4HKzWPm2N1XQk/jRcldsH7u8/rzlRvdBDsF6OaL1VSdr
bdhicXtO4NvRiNEe1EsWPvzvpPGeU2nVJ+Zb4B5/5DeC5MrAZoRD0IanaNmlTFo6
COCRYy+DcNYLjFheDG5NE5N8NC9SyuAIyNaoUPOkogxqsCSrvFjikwJrKHBIHBFX
laY1I7MVWPNZuzsjabtc8Zlb1jaWgiy9FrAhZnC66ujuWP97EcEpGp4xMk0eT+Ex
st3CBs9UTUaE8PwKRMjIgnEtnpGsSbZZV8En9e1rfo73Knxgm++WPY8dA4wvbVO7
W2eBPQ8e0/ZVGu0w7EK89WmLsa6Qs/LqmhHzThJ/hrRnBgCxXXTeTpfyMbTobRmu
GnA2I2pIhnWAZazX+BvhN+PmlZuwV8ni4aqShyKpuNIrzncpfWrjJm491WL4zm1c
qA/Vb2Xr4kqSheX7C3MqKRDar0jl9nZV9UrxY58ZxQR1cswlLGbnHfcj7Q2idA6S
sO3GOQ/tY+Bs0qv95C0HQQdSbQevjCwz+/N1yrw+YRydFZBXBJswN1DsL+tn3hbX
`protect END_PROTECTED
