`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zUyDpGwBK25UfbvJkqN7JbM1l3DB3/+A95sZZVC2ZyDZjxOVHChjugHo5Jh2WAAz
opOx0+PW3tpJbYLj5VOYd8etoHRwwrtRtJBcMO+fJDEVwB/DftbVn5/LGxzM6Mwt
7xSFhtowwpMK6l+q5atr10fk3p6eVCWInFnI1L3QjOwn1kOk3DYiLD2SdNSluxxc
bteCPvsGSbh4fNPU+HIdqrwvKgoWn2m+Kq3bmUCmuGxnogjzCLl5EKCLih1wPc5x
nbluhrneeJi9YZLg4ffOJCKQqb8AZP/pSi7kpe1lqaGNphNGMQpzk4/bqthHuLv4
UHXGrxE9Ibf6KVsRJuLJE+R9eCbXl3fechnC7mEignOQb+trTEwgtzfxBTlZuf2y
hy5dfqUC6bTnkZIHgod+RrrMzICR/EX54fVv0lJvlQ59jbg0q+jdsFi8dOVIkubf
otktjOz7ErQdXcOaMDQrQPli5LCWsEW3xLzIEtEy0iOE3Lfupjt9VahYURqNLk62
2MaRzyeFJV2+KZhLTbbTETE12i+cN8itIV+PFqzFdjIqK0iVHFh0DJ64qNXeaXGa
A49FrjoqK6djFeQ7z4hYDqEFEwUC1yT00/b3gopO3G5V0nRSnDu7JA/uYkUft2xL
mzenPywgExOYYpG2yZ75oxwn6rCqTWeIZH+71C6gFY8XE2LGH1SE/C3Jx3ne3Oe/
RIkd12KV86jlBuYtO0GsY56mX2spRolY7unMbEFHG3CkOLeyH3G1MhyM8SqtpEy9
qxzTuwUiXo1PRG5a8ocvndXomiVSWMAi7gZp/G5nB8bBUwgD+dYbiA235y2ZJJxN
HuCbjCmaSEH8+KE3P2KrJ3OVkHCkILICwuSTEoe4E66GFPjDJDRyFKdyXQfiz3XG
ZoQJ8iwVWDWbCCssC1xwOCJPpbh6b1H+D28yj7SYgW+KYZrVBZLSfA4Oy1bPyzzo
7dudYsf8pwwRxvTYvi1EhVeMVyrIVqHVzeu8aHllAZg7U9aI8MmP318xI62u8kK1
yVcdrLWs0cmGKy+FGVPyb1Yx0kJrgJnGSBcB6g90FZk=
`protect END_PROTECTED
