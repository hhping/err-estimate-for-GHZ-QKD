`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ChTw4OzRietkpwBT/SR6Z/eofvLiOenLGSA8BtiYbNax8hj03KmLhq8qcjjaCFcZ
PqMzudSjPDOSkN4OYbLA+W1rPBDYMzbdkknwfPV3pSQ4pA4DvwJ3B10eaD/GATdW
gklfy6KP/BB9+JHlTRizR/JWGytCXqIyD5yVbs7V2wFef7+uyHPI0vkF9YYR5B24
uKlUig2IAK63aQhDmYg1z4jXd47hW4iD62zlI2+VcLo/Cw6d4XMYSmI1pdVCQKHA
HOiPPqTFkpItb6aTYgbXVrLxljagUZ+GFktj1yTmkEsOtuvl32Dm0FA7oguNWwyu
OpAP0+fAte8JsBQVphxW2/YTT8E1l0tTTA8gD3KHc7+K5NFxsUL2QkEhXVwmTrvz
YA4iQWyfKFe1VcAtQgiTOwzv/31LtDeGorWhkPwrVL8do6HWXTz74L0KwacJ8uI7
MC1fX16PUTsezOIOWaotK0dE5Jp9ic4Sv9AQh7G1tSl9WYjYL2CE1qQDssIIyDb1
cq+exq7RKI2MezXZWhxzWx2s3YLRf7N+nrbDALhNlhunGnB4FplgfgxCDh7BriwA
fdXalNYhM15TRumJwlpJ8f2MNcCI/Wn4HPT5+lAs7aw0zTHj/baFeZTKVHwwfgEs
w/TH3EW8QysX+SeTdO/Plx4wUWJkdDso8tD4RjITe1WoVSARPASrA2ssaKXDPqof
SXZPPhpnZFewSS5p6StxcjRfQU6mXb6Is4Coygp6brwQ7ki+Zl324byGxR/RdPy3
8EdDrY4OD2d2eLd5AoQVL+u5+iqWD22HT+GdbZ8TwxjcVXFXdI4KgYdSWNoex+Gi
wcyK4uZSi9ts35W++YNQlgKjWtpTAWOBxxhT7SqLTVigOKEEL21k21P4+E4/oIl7
NgVfS/uLFomNN4TSxZovd3cCDdQyc5bmj0NPUtPX2Rt8QXZPRtPdKHHMvH4xmhsx
kiZ+qAMXPjEAGURGm4/SKWudfXHRDQGZP6En0Wc9uew5gR1EogAMSwxQKBHyXNRE
H7bzauPzzdIQKM2v58IRulaBkufcl5Q2tpsAFylRfRWUkbjHjMGDqP/YfYYM5CuC
/XycNPeU/34gqpPsdtrvmuE1RuP6mBm/SzZjcmLNy1Y+0+igb3lniRfRbS9k2C7W
RkX4gM+imG4W9VMKjTOo2WghrpNf0Ib16ExrczGNQd4mmsI8b1PoRA4j+A1DGxlR
4zgdQv2eC7blcYbb8V7hSZQguTnhprzd1GVDIwqrz0iUnXJRWk9MzopIBnPlSFFS
4nmNA6VXos7A5OyfoJS4C5JWlHY6BJsGzFevjJpPVSq/ruHMblAD4SqTkODfnbiC
BkJ1zsOjMo2o7yXZi10p55smqsMSeKhRHGNaJl7PGNiW3E3Cu8HV7Sz48/BuIktk
JvDy44KxTSw00o7G3Plb6g9CfvyEYbeB3Srlzkpsji+YVHXxT/UPhNSOkDOTDfJR
IZZeCkvLOms3zWWTFt8c8xZgcT+8SWPl4GOROgiVCBBwGoID004R5i6aYCNodKcE
bC8bHF8/L/y5eNa/WcCC3BmUyIz/lU0qVilUqgJbJ07VAzn9HmnhC1nZiwVP2PtI
XOA+Fkd+ZbTQm912+bGEhdEo7sQUnU1B8MafR6eAxvfkEBZF//hfBaV92zN4r5aT
ipKhT4dYuuZOtUDjQ61ZLh85E0qajh5XMtlrroDPtYcEaAp9+uisi8cf1M6gjlAN
pjU86FvWZhM3MThwLTGksevoSfjfG1v6HtuxmwWdIFjJaejV9tfyhHNLkAoCC9CJ
kBBdcHoPqIjWPEkiOaGCWlIVAK/LNI6z4p9olgAJAH1r+q4jX389pmWQByee+Vqk
EBtDT9LymnfL+pbk7EXQjI6g9TIEdQLVrjc4mFCX38M5kLNQnm+Hafjbov+NTvyc
6TNQcsplyShm9Vw/pNl4IU006z023vSqiZ0in9yYorA5wUjCKntLeeVQeZ4v4Nn4
7uLqFIxlnIeVJ0uqBMmRCmAIm74zsCOZ6l8RuWUkVzZYtYQS4c3FAaLVc8oDOs0E
XtQdhtH4TGXgamDAiA7zI9BenlKkGurJ/KerdZRNHe4LxGIGcJjEqIk7clripIh1
5uy6GFs49Dlr6IE8SW+Y9aUgszFM0MIPuyrrjDohQuZZOXqOnFIsKM88Rx9wQRdU
nlE4eQ/xE0O2qUB903PQeW7/jNzKSc1+MrF9DsewPrmxt6xqDI7mnX0WISiW2r0p
etpgn0dpAOXMWj2tgZsuOBXC167T4YxLejbNYI5Tyj5Gmug0GTwn3akSBdnIiUZ7
g3tPzdFiaFeJnc3JyQRsQ7p8nS4AHuMRfcDxMyDmkqgeyouaL3fFWKAKdYeTlhZD
AiLGb85FqmI9DINfeAjTH4Ui7bXkuU+Ls2EO/TiohnKr5IKo61NqyXbNW/LoBc68
LWq8U79zKBiPfN+dCerkMIMb+6xzTPCQ7qOmnYChcCaHDqJmbLDk2ouPGWVZYK/U
salyDwEo31yLO3oEAtWs2VnNHU/DtW+iTn8ttdwBMTDIViEvKH7AlkllN/GVtgqv
elcNapBZ1g2MopjVOD/ZGfPICTHg4BkqiY6vHj2AerCqoEeAJ+skeOLxlxZgZECu
xPQ+L6LN+5pYL34iQw5HpK1AT/JY5/w69OmIiu/b5MNCE2OVAroI7zlNjwiqrl1c
IgNC8uvYjKZstws7yZIxhLX9tinMOurz4ITowZEfRx6KX+yPBztXA/w5rEb+wADW
4FqUbX7ABdzCVDvo0W4L3LVm0UZS1zmxmaoemRG20T4xlqh8P9Vx9DqvvI10FBPo
nNccc7Nr18APnij4VolQcI8vH8vHU1giH28CSwDL1n14ybnns3x5rFrQUwssJuYZ
oJts1xWwKBG8yNoujwau4vZWBIpS5fcT3peh5ZGpgnQ5KjF+phN6JHFLJckKBRj2
oZCWf3ly22RMKyyAFZno6aoVQPUqpzc4Ar+ynzb9PIZ/ixPxnaGZeqiJQSVfDocj
eqKlH4h3H9iwcPYfFn/aZyEwBF4TGbNHzpwIgXqH2mKDYqEi01UVA+qSzCpPcnW2
7fH6S2gLn0ijo1NQ/VZw8w9GA9ZvGEQcwzJZsIr7YbfyGbZWLQXP4WFx9wrD96hi
d0w/v/e92R3VLkd/Yt+09AIcmNSw9LNHbw/4rx+U1T6HpKJ8A2aPZkuSOdtV0+68
8mrLWDc9dOkBiQkiyypWgffrO07M8uQ+a5g2rUyAOqTu2IOO+OIk+z6tb7Eh2Dbe
xLrS7fW+GWHlrCD6+8VJpuIXXjMBuXZIrh+w5ubRhk/gE3UVciVALCgsD4/L2XW+
V3T2K8usMF3MeYgFlM7efCNJ25ao6/TDwguZ2WJMbojzMM8DlxOsERUbQZlbMv+R
aIvRxJOhNdDXW7AVz0rn84cWhPn3LXRkCXnX1wqJmqcJz0RwYLP4AAzQ/j1m1oAs
u1Im1mdvjBSJNepC2scj8LOkbDHF58sEeW+aeTjZNxhZb17G9tzgwqLv49AHy1U4
pugBto6PEj/fKkSXWYupMqQFleOnwEeSCQQaIcvNM5zT1sjyuBr0khJdfLGNNt+c
AVJqy6fiRcRuxL131871Uqvzqp63JY0aCdmpvM/5gG6tpXuKCUeXfnWaJjr1fLoA
mSY6cLLOgMC4TU24IftjX7jdAjSLe7et0AjcaE/Zgdxz5qNXXqLedSLtGPSGKZB7
2qYPzYgjjQscnPGkl/CdfdMySUU8i4MtGfGYqPH5qGJC27n/W0Z+/OQD4JUc5bIA
8H9oq1g6qhIhWmkkP3GCVTJAGH4rzahQ84qqnj/h7OFq0N4IT/PLP2SpIeIm20M/
7Ijbpfk68nss0TPRyacxE0EubxIEJQkhaZmx7neYrG8/BtC8AXqFf+mXuKG1sALQ
XEHqH7B6vIMJ4wPMZLZuUvJTwm+y2idPeDx0YDWoBP8VuN3r6ahmzk47yErt/ADO
K8LhY2DqVCfzpXuI+FJ9AbqgBq1rowOYIbleEzXkvL+HyTjsS47fvNc5c9cQ+SbQ
kcfn0ne6MQBAwBl0lFVJ+ZvpMtn/+xcEUNlpU1zkm9d1els6VzcJ/ODYmjyc6IZi
dOUNpT0584kkwY//zE3hN6iwmxqlguf1NyELP0zeixhWa6b60kzLauG2yUV7XG3s
Vcg3YAlRmQvyelETc8GZ/qg+W2oI0VKdWk60rFGBvk+oVMtQ6WSRlhpMNdINDV59
yYEsdKl2UVYTTBWWcJ92VnOeLYjurX9JSRGfxaR0M+ZcrWV2viP1yFezTZLBnMmT
ULeKmd+6MlvHf+9c6Gp0taV5Zd8WLtNKS6LltK4pUl1OW8zpHmNleAcPbD8IWN1C
0rN615NwuhNgPiJCc7SZP913ctbotzObBKlWOlx7GCHWFsh3s1q/BDE0r0f/0bZA
HqkpPtKBKPExPSXIChZW8xWuJkLYB2bJLxsDEpTOCvjGhTbhEvMDYAknVZaPrICm
YfB4PdDn61Oht81Ka+QvsVnWGw2IHk1AiYjgIg1s54s0JZNtDILdcLfrt3HO4RLR
u8g0MYkf98I0SqKOK7hstFQrIT+YFLjl2uMqwEQs+Dt0mQg9WMXbRDDT0HZmE29J
+IRrcp1wAASynwmSLzqVdDicfFJ+foYl44xfXBKqUZAOrLJpl7NxWOhJzgCW81g0
TrihfE/azpK4g7jRHCd/0KI0CotDWS+31ddakAZPnwFI3BmGnojvXqwoJZpUIXhL
7ulCn3EeIkYrQE9c99npLBaCMmCijVWGffMxA3JD87Hr43cO7QXXPG+GmA5L9obS
T9i3R5mf/aiXRIjfAUsqVsy/Uldz6EBw3IEuHHri5/QL0rjxwHtSIRWIhost43+x
KpqRAVYRFxw/r+XvhKHR7UuBK9hgc73ZrcTzTBE4lTvXarUPwx7xf4SFUf7a543J
vJ+1laTrCVIob0Fn5AGvWe4ICLxvFhQ1VVjCT7s7t80RLMjVDgIufbOOJxsVKQbg
/eIE2zxEcGJHqVx4BXe71L8IVG/POU+JIUEUUWK4oRKq4hOlHwksQr4N0eHdTC9o
fwTHeSFGkwlrmMfVYu4LLYT7olmblL+LRfVASL9gi8a8HKl2yjNiplhBFwuekfpB
21kNQsiGhyQc71QADJSIRmRMBxvX/lZpHasOCKxql7M94gRLE6CoZizrSu7JCrf9
KDtZPFm8g1ky3M4+WkUTyzTGvIMQFYv3Wk70Hp34vFgTnuc8xNnAKwyWAPuNd4/z
mPNzbjdzM+uZ0kSq+ipxkolK67ijGVvcZmr09vBVtbM6TNypD/3DEjBEHkXD5pfK
oYglDazbf/mRtsVu4x/htTa7lusSpodJPVmeGUJ3hSU5wRvlLZaErKkik3nL7VKd
WVnFNDwB+Gj7MCIhVG+FrT+bprE5GnV+d+vKt7qgkverAh9kB0k3+3hWymMyLtfb
TwCY2bWZSznazzcZkeep5pTFaVe57Ytsilm3hy0BnhG2RyHlf83We3DhVKp3hNBy
HuLwL+n0oTeiKf55CghYuQKVMNzOwI+vnfFrr55hR7Ci/bdHFuWC178QBsMeFOn5
eB7Hi/g29rUzZv1dEs8svk84DzUXPnl2bSeUGx+uJDMDDoPfPVGAYx2VFlIe/UTR
GqgFLxfdb4o4GNWxdJsU/fIkioPLG3aYQcsbEoqTbV6mhfE++p8gxC7gKTsi0g1l
YSc1rcVKLnjiaid5X8ku1xeHsh5Unv81VWOwKyUNA163R3AVz4urxZrHTDdmxtAz
/ZXF2ih6vgAtYJR3T8Mas4KxWBkqBHEj07JoVHcQy/EA5EwLIHQ4rabl+5OtAa41
g4g02VzXD8yDb+CVq6fqyKQ4np4iuyvj4Z1PhJ+7t/46U5GLDGTlBfVug+anxNo3
wqLYa+7LWNSoGpkBF/faH85RpIbCD8XTPNy9MzwWiIpEc29O5gonAG1bNcKb5xo2
BgLvqk8WkyndOajN0lXJlGJglVjsgx7KChUsiO54TyrVXLwMFevquRM5FWH9vnTn
5a6Y6HEcD1mbOeoKyTXiFLCsC5nBDD/tlo46e8OeO+jUl6LLitQ8pqFmRArsy6Vs
QRbMJ6b8kqnSm68iaNr0htYm+Q5A2S7Df2l/9AfB6vd+tKGMUkD3KGuD1xZelH/9
kXTCqp/MvFzZHsmSzzSRMmrA69PMCdj1q9DtaotrvIflCigu/d1cSCbEpfrB0fe1
Hd0ZGZ0IsFI2kzZQH6ffDCpGONLqLo58pBDr9fTgiYxQ5zHObMj2Uh4s8vMzykS+
yAstDCYZuROumQqSgzs+qpnWYVqAAyBoOm8hpxmH5Y5DwPidIljZskoQ5MS7VF/3
t9+EAJfCN6WQ5uFQRiPBIAzXoWILxeAXnzmVPlhM5yx4I20iLHFVwzMzOYqfkzyD
7vKY+jgLLiKXxLIKg5OZPIbKaWBh3ihqYLiM2CldC7BPVvn3Hqaa04dHQwIIgwKJ
huCyrbBuX1i6IhA9gF645wg1WpwfOekQfL9FeJLlnslmd7EWeHzCsP8iOt4wTNxR
1+zlHuwGn8nN/3kO+Zw1cR31Htelc6MB2uvmAb8C+l83Qptl6iUgpJbvI6g2tbVl
Iu6e3Aarq/jkrLsmrNY2jVdQikU1GxLv3bCP1rosjuVXayi5NOjfbdm1u1oFywCM
IaaQU2WBX0PzFJfjmhiFFWR+5LnrV9jGCevbtZyXZUr1XME2IkdRN5EIEA/yGUr0
4eOHX/OHII2VlKETZHTi4XRHFT9hQItrSvnaGAeuVSn0t8UkspeQT/eZkeiqBhZ2
qM9SfzcAMUlo80o+184ZAIKi+Lv8EZUUo2gSNUD/rqOVqqN2O4kHRqRJ2trCjy5X
Se4FjSZ08GwGT3i4zcrDdcsyz1i8Ed8lYdElBM7K7FhL4j7vSxIX11t+giylEY9M
6ORVmiH6YxFQIBU9MDcbICgwU8eewXnhwVTjzKbJYGU1cs2AFm8J2B+vrkvRFjZ/
4zeIH2YADU2GvEBamlIYOWHcWFznao/i2iCLhZZpjyP1jddi996vcJnzAEduRinZ
W4H+bBF6vdKowxX5T5QDG2hoyD6FsjrIJadeX3KldFMYkdoXow85gI2fe0qaUFL2
iIzRGoviNaGn9g6Gase7tnwkJXdZYjfvcYv0Ga3BbDv3ASfCMZ/0/tYBswNNSe5t
PVz5FS6ELtMaSsMSpsR8tm/oi3cAa8g8C2yRsSJM7OaSvUhaaLGi0dyaj9nmqMVE
M+7lNy9wTwMrJ9LcKJMJorrjQ+YV+Xuj36eoTCXVNfG1TCDWJ+GQ2QqbylOaitn0
lUqJsEPBElMActxy5UrKPUl1XQKBfVy29NY6Uj8EWFV7g6ulkvnPrr90k1B8rx0t
K7dgPSHlPdvqI4B6pAVVJ2OefBitGzWqsPA7QQy3G5ky5d5OZk8LM7VYHzd+86eA
cxb40QO2Ik8xxl2V5DPsok/mohIlU+6JlNM6wHqD18ldFHmb38i+yeokbzf16Mbi
p2u72+JSx7ShsAEilrwaauHzISSeE53K2WebRzBsnK1sLH9D33niKnTRIoHaAomA
5G/35tk3VQJxj5cO9ZrzP+xJxSyE6ECALZvV1JGJp4C+6geLM0JbVyEbJwtAjiO8
MEMhSXD05JF9fi8pavHBKckcpeEa/WPWiAlPxh61TVpecHu7y1o09A2aGnGcl7OY
cvSyjcDQS5SZgRJIItYr+WL2psQ57/sKK0QCSB0pJpq1takNT6ZgmEX1YED+feJP
U9SYaZm28mW73b3IaJKK/P2HlnascshukfYAWZ6UAl0zUdmTzpMuRXyb2C1MQWbi
XqI/PDdoVstsejXEGXND7moOpq8RP3a7F0S7bsESvFSYZik60quZDUiX/iIhQqty
ik+YugqgWRwTyaSBsoyE3/hVYWtqDmoDRSD4A8eHojfuBzU9HN6XASPabXlfi7HQ
eqV6WcYIZrr/qEiOLs/IZgnC43QSphDRJpuaEagg7MI/lzqqjuVWvnM1zqrSAf15
qOOooVxBHF1F65ten0zG/sbwTiIMQUWaF04ir0tStR3QsTh2OFcAmzp6BybN9m2G
gNdPgqZubbdi9BCzVnC+1FxsT73eR2x3mRAg2zhcdZ3aIjr/AKeyyCHYrvWeyNCx
EnvsofbM+Q8rg6v4ORiBNMemtyUQm58vNFzWLb/Np/02hkIzVYLWS2mg+U5T3392
BeJ4xhsaRU6x5hCSIkL3zKAyi6KrFChv60Jbu3oZVoLGhwBAOk8y3z4M8RRZ9a+D
msfhbtSCEbkvsglPDMBGeHV2qnhTmxwwOiSdL6TIdchBqgG0PDc3cMmf+ZQyv3BX
j7NbH2k+yFjvhmUgHEiAJIeKRrk7c/RU18q/hRz34HaBLmW8XR3eg8FHlqoRPZNZ
ZRkMYzkO3Kp+NoaUPIt06/xdQ6McQohxjP730fJVRzfLFAfNeuYKGFBSZEOf446p
2kEhdTLY/fSgwLmUstMSsY1yL9cDn+eKLJ5q8GNtGqRv1bjxOGdjCD6yO2bzwRjE
ntYtoFzLYswjlQr2heF8sKIiYD98Nh7Lry5s8dqrMe9BoyvxIC3vfAKsMaOem7yw
pPlDxDSnq9AKj6J/YbBe0bombH/nBPI/P6jS/YqQyWp4BkRSf+7jpZbXioM0GoQY
m3jlZfK6+i9dGYi1mh0VghxNfojHGrczMPp26Ev0J+V5vUqQC1Dv3vX0FG60sA+U
vImwT1DfoTyJ9GTo4KMpehjstGfgHJvN8gnDZSTsp51Vunqmp6grQOOK6gv2klli
jnLwU8crjb2a1PdQcEoYaAd/cjkMDrLgo+YdLvjsE6QVjLEeS49sjAKesHs43kPU
L5Jt0OOH0XBzsOc6kxBQ4DD0bUbnDMlkNT+amdimgLSMJM1O0r1WitbOhUgKXoiS
HhkG4KxClNxus+4cB7ixquw0VMRWqpvYwwRyY1j3ry5q5mDaq3qKplELDT99xb9I
l17e582u7QrfNixb6GjevSb9J7JOBXMD3dmdliyWL+12aE4BpM3GpivYYq9WzyGg
LIxBPS08OGV4wTxCxC/s1FKDp1uaCsheN6C02NWk/3AQLU5gE4ZRbsW89pzQFVVq
RCi8K7Ey68VvQPrNAnqECAgvO2GUuLV5GT9mSENBs0Xc+EDqaq7wkr7KuxzChGko
aoOoOw9IVrLj47bbnTQjz1nFA6Uvl7EEcmY8uWBq4GXYp3ZhSfJ+WZjYzr9IKBiA
ielvkyHZzeRrzHFL7F3OzKoTF+4KI6GkILkGouueJtDB3Z89TlfD03zqRG7JboPW
VZrrPMq+hJS0HAbNhLHvs01S2gXjYJTXy9bNvFpn2SKJMhiY5NO3VEmDVKcHqyyj
dcq3NKSLB49zQ2VONKHKYq9xW3UyZXq2JXokJTjmxv1DsSQpn6Qu6849mKUJO3Jp
khnPLHp1HE93A3aWxNGjrlUouppLRJj503SRKutLxM8k3cB3h8gnEGqLb9p+LJST
BETADMSySk7rAsEXBjRz1c6KCvxrogriY2n/Pny2pVf4GrkLri7ioK+raARYPEuH
qsCGON97t4nqF6ULQ88XMyPtAqQCkbyhVUGk2HHKnRIJMCA+4LJnuKWunE7HH4YO
TCeGXwu0sUkXK4qYvc+eTcj8WKXZ73ck1eKDtWSLr/dChMRW7D6CqeKn66RTf+bd
NI2tDJSyfmX1QM0ae78/8/C+OND0sFmPJlflQtApuvSamG2MLtY8PfBrhbJC/IJW
GBFC3COs/J8pw7sOYUpGhy5LzUlV8c5KujxMidyqjDzKwDPrnj0T/zpX7yXLZnnT
RvuArksCIevY2PIe3UM+CRm3/Qx0+j8ImR7ci6ZNJ24hY0W0lVPZXl8EQzH+HnzU
l1sWpoEIGUGfw9J66qxxtyS8Zy+9kHIDcHLAq++fXe4Jzlynv16mqieIHckoOWLe
a23QddugvP7TB/uOtbOMFxueyQFWZuHFc+Q8xj0dXRapzDnSxK00WJBpZhg4pESA
dzUa1B/kr10vVZi/nkOh9QV4S1ejZUGrjB91d8s+0A1jlNaG/TzR7jr5iVGbIff+
aqaTIuEnuVOso+buC/F9Mvu+/TKDPt6sS3tjyCNnuhAl58xX7pW4ZBl7dGSeHdu0
D/FXiIMwiaAiQBPDJAzfiLltZEwUg+pL3aYL2Wb0Ciz0TaCV9fBogQbcufpbD6da
8nuhBeWGIwgpAgbxEfEQMJ6AmYjF2s8qKBd7ZrQQOH6SDu5l4I2z/O2QpwCM/tSA
4H3xOC8D9o2rohaFTpQocVLTr9rSs3wZEK7sSQ2A+H1a5j526cQlPWrOQq+RcdIa
CJD+NUTq4eTzHalz6DAxQY5j4YWLlTkOGSQLiZC7YkFssvLhcZc2qrZDf5qM0JAi
bmJyjmUqW1ENLBDjbirCXijlx1UbnNZ58kgWAsjtsJKPxxlxtwAvxmjVd5cE3YPm
LpmuxGcLynlQAOjiIXkHc2OSi4/a6pb+sDHRRY9ngm7iqhkWsqjiNwP2LzlzVAis
sXGAgoAGBehlhRUS+4kCXXott5VAUOtrJqDrYkbfjnBlnmXk4IdTI3ompe/sQL8G
i/kChSNezbHaYvWcS3PaCfNHkSgqtEvVTy7g8tlKfaWTcY470q5eb5XALcTgEb4e
FSxeBpUFuxjoirzR32zFs/2gtcrBx66C5M/6b0eOhXI97PJ+hHa93+JX32nhQDNv
OH0GeJ6IyTqfVrM/zFW5tZd9evF0W/w9ZTsjTGNu03J2ATkEiKxLaP+1C8gNKiXO
K3WPYkIG/2K3WH/vWdKYC0allP9n22O5ZpggQkRM3xHIUUjt7U6qL34bdOgWMOhF
fWJi9n/PUtj5PnSsb2lafaasXLK4xSyJKa1NZn1cTdn3IQYDROuUt56XrwlNAPqS
dnc6bgz/bXQ762TwsUujQKCLakJp/atuQBNzPDKu4g4PulsicbVmjzR7X67BTspW
aPCW4s7ke+ucI4N6mODVIPcooF4lHHUAliL+/GLIuC/Sj5lTr0l1Guhp6ER5oDb0
GEYKzwS38QbBqs8kxMJiPHUhJcHG4eZuKIX21BL//p1gXb1x/MtOMmNIKFZ7G40m
JMpXCYcy2gk+MUkZqOHN7fea/lrQs7DYBUCwuNP6sHH3n67MYdkiERqyWjZ5k8q0
LEZUexJxD2gdJPmsacDsGgi0y7H3JoWlv5munMg2e3HCzyzNAhcvfl30NInk6ZNM
D2bRne2LzgFi0cnQGkbqjIDSxFbvZagrJlWfFhwVxyvorqyjtEKaw3cAqNAQNiVD
r2vc9yk5TZOjQp0RKh1NYrr9CNEeKhioMKclUwZzM2vvNglI5HCfIhQAvBHBVRtE
IlgXdqbBEyl/PCyjv2S/NJlIyfypnaolEAGWA9zaglfYiVrUIVTNPxC4tJDlrfc0
woZ0NDL+jx7yR0SMiSo5hp2tUeJNwLD7aWfsriUiriRBE6/w/N0EKkZfRRPscrnn
0xHrNedBgzXwlsl/TsWVlyDRaFOC3xAe9qDzp5k4waLWDqPW+dxBKr6KVIM+DFqq
N8RiOzPk8DJFSwQUnRDaAcehQcBRpg7P/Ohg4nQTjiOCygSy8qoKmmRItHz4udDS
pDV099jUucAY/nPtibj8iB0B4GNntGBveQDip7a3kFTGa/3LB080sAZpgoHytq6K
P+cwJVyf8xkRzsSmsJT4S7IHI/YpE8GN/7F5VZ8yAh9I5/krH97NM53R7PdrM8VO
FYvv4NbVh9kKMo6LE+H0NK7AKA3PVcKxhyWg/dx5sga3+2vMCgVjAaRbb3ez3d60
SSeLMvrC3kVKSFgvb3qfMmP1kf3sKhdfu0wdzi1IYWw04Bi83oon0+TUG3yBslFv
3gUk8+GAWjsNnSOKsKWErCOrFBgbGku5tiifI1EeR/9vK1mtrlySRlIwnwZ36MVG
7ohH/SDatMGQkHh59hCzAD6rFmQPNhQZ2Spz3M6dOO7X1Yu6DTAwoP4/+GmTZTMa
BJG91YRE7IT7iV+Jq964mWjCCCxzFw3HV3GRIh2HP8jaDW7KspiEbRzwMtw3+zmv
a6k1OncsheEm+LsE7PwW9Urt1l2CeMhOI/UAQ/fwFHT7ehdNvJJmZ528u7qIsXOV
9qVdBuIrTNEfqJ0H8QgLr9aSOkr5OjWGKq7UEvj4G0H+E07e9ASzfrYaT4D1eYST
O2/2lhGTxYHSz1k79C78KSCAzkSgGcpUGATtIRO9LlzNod1+iH/Yj3eUn6cF9fnV
gjdNZeic4dSce1aOhuwwDk4DYyhaEJd9SQG3oHbORG2l0gRZ6+oXOvgMGP4tzzBP
qwA1cIhKq2Rbn2l/YpvOnhkdaiQWugRclSc3QpbENFPAEU7kPDA2EgqcmJrTgpJF
2OFrdo+U0s1K23az6OvXBqb3rRF+6aB6GHEbCm5mBgazrgMSxs7OI1lBhFiCQwJr
T3HDX2UGEOL2qi+ek7g68xYPZnY4Mw9H22DgkyLZT8aJYk43kYMDoD9vvC10ZZid
fCX8YNNfdj4OV7JxJgVkNnlZqmOovqp4GBPJ8O/ipee7iPESt1VsvSbZImdtv3QC
joOvKYb8Wq8RlncuizQlu2s7J4hhiRPAokx3EFiijBANTivs+bPwnSxRq3NxySHG
FXE6KsPM14Y3/0XQJMVLJze1PTiazKq8Wrpk0bDFakZJ97dkPc81Yp2GAKaHDQuo
5cK/kDPNDZMGF5i5VW1mliWiO4hZ5BrZDUGh500KGDqSWhDdQSBcmQc7MkOFuRas
v2tanIXgJnAIk54LhOxwWzsJanTZMnkwpE/xqHS12krp8f6wl821PkUcrC0MfqcX
RS/kdJuKMKIkmt+XGUtAR65D3yCipXyUvONVwaiCnacYHbkNfwMaRdKakOz4RVVp
9ix6TRCg8xE9Es+Qz3x+TS3DqrZWPjdH1pPGildKPJQ0ZB8mwNUt993ypMVgSKGh
S35VWnZm63Z0sWf3K5UV+bpEzp3A15S/pu+8O01IGdkP3e83pxX5/kmRYT5bNEu7
lTa+t6Qtk+booghLovg85RnSGeroGmREQko1mes7SyisOIxQ/zZ5YaMjzqyeyDZB
txT+FRLZHnIwxgcLLW+v1ZdGmNQ//o8GtoS0lLxP69qM58lE/40KyMsb8z5BOk7o
zQgMlRm2OfzGlzqQKJ2PL98WQpExdhcSFGVvwfZigJgiY8ZF2FvdqUVrXm3jfchh
QP/gQlCXxTeVLJxpdyegL26WjXZgQoeXJ006FaYlLksEICQHpw8lDQgPCfAQWBGX
a+pI+RC47T6m6SZaB2bLiIcSNTkRJhX8eGGmQ1bIPVomGD1N2mdqJFfD6ZYX63Wu
A9Tf+n/df4+gPI4Yzyc9i2eLi7VmpDFopBOM8ri/3G8EbCyOT5z+TaZ0dCO5LsHx
7G9K9yDgYhqwfDvN3oSSKW4B0rXmTO6EU0mL80yce0sIHwGLRdkZ2hssUQ59yV28
5AdWYQRgU73XyM629T8aLPLJUx1K9Bbdib3ztQZV4JDjl7/ZNVKr369JdpCzS++Z
8u7iwZfE1p9geO2AU+RrCDDSJJf8SJ/VNBgsuzEwJAUkeaxZ3ur/zLA8T9MJpliw
JTtow/NI1O3Zjip0sTlCCbNSL9U6Jqjg+gWV5ygtAsw7reR2hj/N2BWs7re3GRe5
BmGxUGRSRxVPp/CS72NV4vKsZeHiUa+oRrzV4LKXVHWMBrSUt2fijLTWuqFfMPaq
aGa4OTCWDAtbbI6W+RnMAKr5glmixVYEzzaRwUbm/MMjXN+aKgY19BzzHk4oYxBd
gvsA3Dkw+s1k2DDjgwA2Ck8dhUcN10IZlILbaM1hEUQsVgdwUd4Dp7TvcLunFEC3
cNlhi07rxYl7Ho/TsLuYo+6a67FHeibFY7+EsHcmeys5zDTyFzP0Il+GOwgMZD/P
BqozBms7tl1Ylwfq6eZv7Go1FcyFuinpzE95POc2Dz7y7Pv5LWqaVZC/BMxP6pH2
yMbRVRoCT6wT/OW132C73MJFq4L1y3cHltTC0YSRgOwgfBHRO36FgGw/97LeHNBQ
qeZbiserDJ1Be8serZkjuZUVKoaiNkdSA0PNA1F/eNTYHfUeLmB3RO26z5IiM4k+
22txHcI6IzN4gl9cfQ0wiCr9xlPx4gc74DpOOj/LvKvP5Op/fqi5XdpjiYH/tbpL
Djf0tRoAjLFMrizw1zst5Bua9xC8OWioF9jULuqMee7Ury45eoW9kYPnXKcv8RjS
pukoKNWoJ24J2vGKQaMsWRg8HaJWxnf92UiW29zhZd6uGs95eARMtS1liO7cCwnR
5DRVhNK/p9H3OH3+vnEM8ulWL7ik7J33Gqv5jeftB1gofXM5G3UV16DHYOw634G5
Qk7dRysvpFlIAXGVsndiQdGmffst8wyyoZRluCT+K2sqYFY1WzGTUK0XS6h//xDc
G/YBFQ4A4pz8uG9MQUwmnKmsfdp0kbiILv9Zw+Y2aFxe7Qka7EG/pLuhOPqDBRqi
xCMvAAetVQqPzuGua02RT/Hd/bHekGK0OIJ2DJJzck1p+fGohk0oSCzRgRNaTCWB
DaEjbTddGWySuvCCTVFe2mwC3bk3f63bDDb5eNZYdI/i6gCaUhJsFxcqmJn4bNtb
huzJct3xlkVTtD4ykbMk5bjLajjXmzURMtix2vx8bZtogS1zQ5G8U2DWs63boM+N
KlYHphpxg57I5P9CccgztM6EBsTkvu6n/cIoQQcbcr6okyfb+tGIqjR8DtZsF3WV
ZYVC8FRWj183BZYJC6YGO1jAzuVbejNM4S+Z8+iM7CtwypxYY7HrZ/VhmndjGgJ5
YtxsXq9xkzc0QqO1SyoLXNA4g/6JHoEv9PMAubE3pYZnbGkmE7OeLv6NcgcAVtaQ
5ea9HlCnQ//YXYpBUs573zvlrYD5Yxuo8kLaXX/p0Sd3wnFDSP4IFd62ANSBuBRh
QyEdxp14uS1Oh+/hg27v7aN1fek6LgfoB64mY3MVsLL9pHD2iUGWMKdDBSP/kKNN
XaU0g5aSVHDuAgoO+tnczJK4GZzSw5Z091a9+Vzf5ztbmFdsekBgMouMcG/nMKbY
ldJHKUQXVQflyB5zOwR9Y3SwfuTH51n2y3Xykd/4tKDISHJvhNFnYD5tAiIdboIf
koxe4FZM5gR9cwUMKDnoQjk8HvHAyhQCh1XUhh4KUIDGBjuxQEWBoT1eALy+fDp+
wBbJQcLjyAQ6SQmJt5OTV8KMLj71vP1PHjZpHlFHnKVpXJERa2DtvfBGPl59Edvo
ta4mwXQcjByM7AZ6BXnhADGVKnwVfMmMVLEKd/UATF2AiLD1LsM/xAYeyN33wl8e
pCYgouiflwwwKatdjNYPztzQ6viNcwRNjW2xw15NH8fW4w4FkdiiqzNWumhNp6xX
yVIReIFBAnGmlf1kyKITsjSLd/vi3xHRG5UZ1k8y1AuQpYKX4zeSx0LcTuuJMLmP
YkXuyZCFU5bcxhhgPxN0dps8Bq9BQtSCGa3/DRugegp2YfZHlgELmXnjBa/NTHdj
QYa2Hb2a+BAtORZP/OkWQTabYDWHwbhjttyz3868wB6QUNehE2jp3gCThLetx8Na
DfEvW8IVrV5J4OR6K8MoSHlJ1zZ8PEMCwWb8e2G5JrHpaz3sfl1GmHq/l5oeC9ib
9O0Xl81MXjEmB4JMt/Q85HKWV1LE7rveKMZBmsgMyxOGkZF3e7V6I6vJtNXgwJUl
3YMW1qJM8caichbRoAGdhTHN87hckBccs5C3rTsvx+qqYvyeZsdf/nZssqWoAno/
Olin+n0lYKw6ZVXB+ryIds0DDkhVaBzGwo+rYwihcmvCilBLn8T9vQHXvHSdiVdB
uGiQKRtN+NvJV4/bXo/x5tpn0aluFWesl64WUXJpstsagDlQ5FXVPw3NmRRMrTBA
9Nv+FkG7zar+T4FaQq+wBlZ5SKCUdrCZT86X7kmKZ6rNku4MTF/uovGGpBDtH1LP
mINSFvahskEI0t/r2cJ8IYuB5SO6t2ldliAAUdXukNoFHTMe6TcAdxaVoqQ+Ymq3
mXHN91wT2o0TC/VM4j7MJMmxBxyX84vnbrZ8inELGLWdwsHgmJSTIryczjSBCQZ3
zy2xcS5E4XmR0Ff319QMWetkT13JRo0lILk1PpdmPHnB1ofsAAalGKImBHH33NSQ
l/x2OcgchHCOLYyQPOv8lyr4+HwrYVt0S5X99+e6YaqwOzXkqJE0n/jkzztpJaUO
Oz1kCzInNtHDy2KCKy/fZThv0ZNudthHRagybVjicCgBsqTTqm5bfHGZ3ssO2ghM
+c0WHVjoY6Q3Wbk50+FLpTMlHxAh7Low3dHPOH/J6nX0TbtYD8uQm0d4Gciry8PQ
cDKCrxEJlkrIM5Z01AmKgc7JvqR9tLk6i3f8c5hpzLnmWkGoYhDzhWypWzpp7+QH
3S9xhn5unA3YxF9LBchBtAf15f0c/4NdmT+D45M7K1IgzBIX4H4jGTMC8+dqLWZi
XxQTadkygCUmk3j8fWTZUoKW50K3Lat+7kQYa+L46DGoBqXi+AW1giPZDzqbbOd+
sVD648qUTQH/kRp5nmpJH/CSm5yL53ENFBJyVgMBEgFRjIgJCylYW56oXxSDh81W
MvKs9JCxyTN1mxQiJb97EJMUluePqNQ852Ar8PF6f8x/l5NDkuPFIwiLl8UDyzZA
bss7CbKHmyvJT8LvYQxNfx5kBjA62IixwWEusQ/LwExRSXNG2I/Ibeyq7VSMIrhv
tQyvwzAbU1y9B6vk19xHBLL3Nh49oQ4G1mvhZr4uLEELHKX/QX8I0+2P5OpT1e/9
b9KNfbHsZR3ek2YzBmIv3ZtZ74EbzzAFqn/vVHZh0g7sG3Zk78w935TYJl5foIES
SeozwUEJwwUr1K6hKHsO/pfBkPfyTe5fAnlXZK0VttFvPEAEArk5KB5/B+t57GKt
ZxvND/rqhqdbsUeIn5RHvrlqUFQAFcFAgsNHG/g3amCXrEAM7DCVxXO/ehfSTbnD
7j6980mT7yj1PSacdfLf1gEjbqAw0Q2QTW2+Sn5Zvggbdwr0Aer5scpjoasvscPL
XUHtyfL88z0FGuC/Dyl35RJ44f5Qm6MLj7y/CkibryPizzKeE7o52r1akVXLEkcu
2/3zd7LXI+aFqEqs0f6tXwl/qCX6y7Sm+yZW1Fd2liyHGdlP4hsVBP6Bym5Ge8+M
Pj/dU2sYGA6dFFqTCNihgI/vvXcqLjeZA3YGTvVm+L9IRtAb53tMFB6cNRKYb4hT
pvEOpxbzosziaTJkzPOey7kM8epUIHbVB/td4F8Z3Sx+eqwKQGxCAg9PFqi3psfr
AYhU7zH0m6q2eut4klW/UsOmoFPRMaoIhxGH2N1AIU7w1Un0RgxBFPRMY6aTLbbx
IkZdScjK+IuMgI/ZCP9RWi1OuqhDo0FQB4tUYMjap1xC17aeVKg7povXPN6gRC+7
4/EYeRoJEar7ZsfVk9QBDYPTKPUrCtZx1MbuPnX4gLjgKN7J2EwYSKRiTULbNkyx
ENs5FbmaKYL8YNYbvfO9a/OqPyA3hdSI9NVXHGosw7rILlbYXrEjP/vdlzAaoqeQ
PLYd+pYhFiNEGR4N7OpdPrn1KKGHQaYRdygRrK1Phg1u4p9njWA2UdLNO3vkzzXN
Sp8vPXFYG5b26ywB8/q4sEsEb4P9SyDl5YXpSYXJqvOKkVEeR+ObRqkjsUD2Jr1G
RZ2IChBIncIxWYG0jrSL3fe1CQ9EA9QWr9PNX0dqmY9wHs+5kQZ6IPu/7NquCD0l
HYD3a9kq3Gv8eKSiZ31YP25xm3IAMDNDrpi/TWTE1gfpVOlWbgYEWl5eCK3+4tJw
ntgu/S0ugHxO7DOIflW3SpEWwpVoaUfCQwxER+hdM9YSBYpvRL8HzBWcNLUsV6yS
p/HE84AUE+wRYpu6zIxqYdMHq+tHiWtigPV7mFQ+SZ+4HkVEeKRvMf2JBUfWl5dk
592+DQ9P3gYltmC856plXrXWdRJxyMJfpqNHU6RYm8ZDUpRgE1wiV5/0HyMAR7DP
i+T+AJGJ98JisOpgSwe0P58HMWgzesl/gu6brH1tTzdBBsAsdM34o252sQ5UEtDU
UO/tiBXukrFqZoZJrP47p5QRAc2fYhgvH2kGqQzX9EPWWYtkAHqA/SpMLc7QisUv
b2+P450oULTrDWW9290+KpK+Rx4zgBgeq6/Bgl5HEa3pMqNQgNW9rv6SJ9beTqFR
8tPupLzlfvUgU1BZxVuncGpcXdoqWSAZFB1keQsV9yfTPebHeJQeQMTLkEntydLQ
lLOF3A5elo7hGtjU5+GjBG6IkW/QDgLkxKitzdwm7/ZH6lK9GhRk0A7zLNnfwcVs
Yg7EyFoPDnQnHVirBFzqaNaeIE2jgO4HGTpbY3EHd1waPD0EvVvdtlqlI5ntQETM
Zi8mT5HZGmrlH3g4Os0CXUttf8GMg6yfICXnk5i0OhqE14xunAoYgKxZIcqAJGRl
h2jJHJFkF6OeJsaxXtqLNqRgb3PL30ZMizcAqvObvS90FpOv+U0je1K08V82gKS0
zeREUSjGNlOgWR9W4VPbjJ4nK6TeN6Qro+VJkm8FHuQy7zb8ZrOKDIIno442sI4P
ZJGbA2OmWfxZz324nKnpNbO2o43uJYrPjYi12BIxCBWfoTgON+FsWSe/1Cy3ZNH9
xNBC/gUVCK17xeeHHIUUIln48KUnP9sTt1n34NxtfIW5xYL+PyEv34JVmaFK5w+q
KZXwFfB+Njmkt63VxR0YiAC0rSJjHdtd3KR8lC0DdrtiSOei4IR0FglZ9GNmYGHt
Q6PvZaXgHSSosfRpW7wKw6O4mz6bkZ/JWxiLvRpYtZ7SoiN0015fs5mjVZ1d3YgI
7hEHESaX/FL9H1xwUK5v1GWe+ulqp0fkRQD+JUMz7KXSkRqLhtL+ed+ZxMAFWgHk
sEddNYFPIshBTrVDwpWtgiI6hs9orJZlwlDzgeVzqFrpr/e4zHNc7169bIR8WOpG
ixoAYMxK4XG9xpIb8Sjp65xs8D8HR1MLhAmhxI0SeXw=
`protect END_PROTECTED
