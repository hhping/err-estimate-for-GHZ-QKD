`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n3/zDsvPLdN31Pdr6gbtwFTdn5x4sm9JA8bIMraEdnXmzyI3AXCgmYyXHqk9NCIF
0pGIzs84sk3hlVjYXZx2RZVIxQ7Pjnwr9ic/tiliYS9JhsjD5zgTuMXuRh9Ieg/u
1xa244qidfyWShMI+qhNDuT7w1/1b7BPZN/iXE4DB4YQvyTFguAItRPXLgyoCDu5
vniuUiOcQuHsV6VgRJzixnQaArC5sT++DTgNPGzPYV1deu3RPL0adnjzYYrmTwZK
0yAJ7XIPzDSAVUsDV6JkY4bp/eVOuNdKxztneEFkXEC69p9f1GrnHPVfmw/VNXOM
qESq1RrOvkpuSr2kETkVWUKUvQJrQAOhNODAr8/p1NPqpjuJXe6pJotV08JwrERj
ObE1KFD4IcE1k2HwpE02P0giCtvcxYRADA+/ObxQTT7qdRbJvgWRlMlGlmURMy8I
ht47qeTWRLgBLjiV805XHglDO2zAtDLl6JW/C7ERh+pi7qc6h2qBsMGSPtj1Lo7O
86yn5bTVqjAQ/pwfDtwsT3MwI4e1Xw+X06Mi0YCxmkCCzKQFZ/ilPRdsnlTlFy4s
a1mLb4YtVwZ18/6VVghQva4sglZ6485DdtL0vwAPZ18YfWngicjJk4Gc0dwN4cD/
tD1RsfjrLDDP9oMyfMTCa/BpAdTdfMbiNRJBsivKumwl8spWXGB2fCtVCSL+Qb4U
UDPxxoYcF1W8cN4lddwA1f8zdiHdCW3RYd6Ru0BBdrwkj6ltufu7t+rg3iAaRAtJ
R+uz6cABlPqfuoOgFcAtYgMnzPvqFX1BD6U+J9pLJQ0=
`protect END_PROTECTED
