`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aBMi7yRiqbdS6qdxc6gMphhqzrP8EqV2xccxSvHsKbP0yZRB1tFHLmIWQBGfIV3s
liFtxZ1Hp1qSkr3SUW7cpU4ZKe5X46MwB/VTJuGVyMlwQXiZ/KHEw1mibyu8VING
DI40r0H+Vm5qeHCluoOIhLoEd9WDiszNTyIN5pzfpUtIsz26hY9ZVc6OwuaumjUt
YgNK3w5MezxlAKIhvUWB/l2QEa7r4Wb3Oya+YGuPn5yPyoGRLGr+XRDmlqEbXKFn
OjSE8B5EYXXeLVVIk/bqBNxFaaMdPiTngjUR3ebIoyaZiVdp6uB4MlCMTu8rR7FC
4IcfDehkOjnDXU/H24dcO8Qu2jJKbQ1jtK6vRXR1dtE8CJd82zJztWStH99PKwr0
nWmX816kArl7Glb/QMy9KcTU6Nin2GsZ6KTD5OAyEnD/aGaS8WtUdIT/I5ZvkxKu
srrohPKnZ9NrgY9IEnqiLMuCR+9tPV3PIW6m0tEruXge37jZDGMCEBIJjYpzURSg
p2iK5C2+2kWz/x1RtbOP4ZJgClVKk+XLudDpaKMZQD/SR8xTU9SejiEUNSjOoIl+
Nx0Be+9SM9rKD3S/ONcIb3fLAAmZR8nJyABgjq2SgxkyOCaXY3+XoRXy603tTKca
NeHZK/0RS6LIklloSVqrFqIX2a5eBZTx9yySlwP4z847wKETD4mkMZ3ySj1Ebnhl
b/3SJyxojg/MDVRfJZydBwyuJSpJ6og3xNnMDBhDBFzMgJeLF4mA7r7Fu5lnD3iZ
Bfr16CyVbzczfnUnOqssc8b6LWGgVPbX82hZKYMykCw20L+/tzb8z6gCFHewPVrf
ANl+pLB+4JNZc1CH4MHWgx9AlEVwIxK1R0ZFddPy/D/97mP9F5ouMX3twf83CIKT
ExntvSx4Rnfav7x6iSC61+nz3F7adqNMxh3vxPsVtxgCRHD1J6TEAlNy1KNhIyhy
n2KIXUETw8A/YnWgT9WjTn8hpretUayLDkldlZjOrGDgKNniOCYdWuvex+jyfMy5
690qU8ASmryU/9NWMDB95MNTB6hDk3IPD+lD3Jq1IxUQa5bnGt9c9fgu09R2CkN9
dtulY0N89w5tmW76JzmIZ5PHLbHOhmtG1IXmsu6s30IaK04SmGxd5YVUiH+Apddh
A3Q/6wqOmQPFS8S0TwkAa3zO/T215RT9dRpDxcK/8ZABi0BwImhaPxt+IG0fDIta
Au1fVJTqRKLlJf7wsa2WCuaOfLj+qwRru/P5/sU0OwpHI2BN5q4P9MnX+Z3U7WEx
VrpNfZPLFFNx2UCUp9QZ767m/fCluuMWJV44RgDwquiMHMGRluUygpl+oddQkHSU
02JwZYYeP8DhwM7NQrs6rbPNFey9l8RDEiZFtEZT200ouNse4t/hDNZzFfM7DFDG
S/Vfpv8sX3B1ros7aXs8A9/FJZaOltdTuDwvcEkI/cEyqjutLynzEMI2xVD+n5h3
`protect END_PROTECTED
