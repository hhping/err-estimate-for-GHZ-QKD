`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hUv9MduUGYUSKs0ZQosgqUtUEAXdlNw5nRtJM6WQwwPXLqY9+m8qaKnXnyyKZIS8
fDs0hLKvKav0f7MwQLyELydiLTruIKkhtuG4PLj8pi7yAAZ5UCWJ3eKl3iAvoBLu
XDirAN1oTpbaEmhYieb8YUHC548+OXY1Myp+nRMx5U8AkqA3w8TSyaboahm7hndw
LYStGxMvVFyP0zP9xIaqYFMzEMER4EHlfsInzGblhhnBdlURZIrehGNo+wzfzVit
Au9CYEk3rpENrKotJq4jCLseu0GP0f6tCeIGA80+/85CEkTgybmoedHMtLOZmIGc
JkU3fd1hLlDDLQ2XOqimxUjfld225OdNB0M7oeV+1z55WH8aqf2RSz+qoxrvoyI7
1jvJLoMcx/FgAtrV2vdXueMgpIvjI95EXZIKyBo3sWRuSajUeSVCFGRWxQurg8x7
t7NAIOvV+dliVIJ0KecssP9Y5mwIuf+PI8tvza9B4Js9GgTaURYiIv2hEuz6IghI
N2s7KYUR1LkkmJ08EEkDeNGvic6PpqAHGZeC6GWO2pH3N+iTvb52+Ou2RczVERQK
r3hyhhR/l1VaxJ87z7GilIcHAWa7RfH5vn9gqy6ihxOgY+3lmCb1Hpt3bFk9MYSv
oN88abEt+A0CpaJO1JM+zd0RuhHcq3zr2HcXx2SKVhDjo5Nns2j3mBJAuUsqh0BW
TAVGnaMxpqVl/0ABKlu4nr/klU3HB2Au6hGo1/inVSf566G8G0b9j0FqiWy3yc6+
xlwLW/1a2MbD7QKr7+nua0yfeih9keUSagsVQDOupKDqVxSprYDJPxvJzt1juN7l
qhO1vhfWTzOuwSzfUdeQ/vxIpXLr3XwbrCFFkqQvbjK36AXtP4m7DjDqjN+TFuvZ
lJLTqmwLX0ZX0H5G2L52cKDqKW8JGcno83gR7K3aHj7n5f2YoU9JNue4zQSepnqP
2Ef/5/rEVro/THP7/DKOMFcE0hhyOjWE9toQ4xEL1xwnWIR2dkvrNxyu9EKXAM/x
rEkPZzD/3xagOx/lTi7LRyACQCOo6XVw5xNZXwnTzZjPZ/vUu0RdEmh7VtQuT8ck
fwFpBS2kVPM+U8QPUTAvCS8XBkuHVnyoZVfWtpiUPJxdbA4h1rTGzNe5J9MMjS+K
LEQAJL9bOGEjlJCPQdc2HLUf5XYjt5H9exnTtIbmSQjeu5WlbzFTWoG3S1+9gVjC
CM0VHbAUzJ51fBoXKfOv9G3qjoy18+cIFN/snWfTG521x5faV/IgK58Rkt67yyLV
fVKfpJMuNDORUls8+HJ8Fesds+KQCle33dQzb2Dj99wGiG9JiugwABM7s0B2koGo
2ZWqUSmr2FjQFT1oB9hdprldotIs8UTjxKggb6+7NOQo4SyeHmifo3Ct84ZKDi5R
bpkv/28iFuCMsq6/XFhz7+X3BTw4gPHx9tqdg2ESul6/n0ZW46Hi4Fz4swVIKpRT
Zq8xJ0WXUJqdeyc4GiOzzJgDCBtpYNHbSCH0f/qwMd9lUc7qZ4dNW3+7/f8CVzbj
AWTzIxOr38m7+mnY8hci8LzCFC2FDjhRO6CrpSvrYr5WZetGXQ1QxNtXwEHZYWV9
eEYEcLxDDQEILuF3F3h1DoycL3wZxyFuZGxBMqM2GClM4F3AboO3IWqy7WDvu3WF
hu5QS4nML5TpHqxVnPwqU1+Imw4RIcQZ0yXkRjo9qk/iZ6cz84XnilbM61Y44YQG
LodHlfleIBSyYPB1Q+qD07Ke+dKz2F6HBf7W92YJznORMdv+snHgVJZnc7NFlmnF
upgBggiuJqvJvLdcExzsEaK5hZFVwwJH2/JjHePqZVgv9WZpRRA70OUBkVXxdexy
VvLjzxJ0u48HS7svXtvZIwI7vlJHM+Fsaeu6ETKlb1qq53SHRuKLLWs4o/M1sM7k
wWQFTrCUhjKtiMJ+MA4dMuBGIyI4jfxnN5PxOH6h/zlgSbWK6Qy5kY2REKeKJGpU
N4kO+icbE2svvNmjhNh44qc0CCd293xCzebv9N0FPTZ7e5Na+D9ByxxPN6EMEEEN
dTnR0dXDmVhrepo3SrnZpDlZez9zonSeRXdEK9QdMrye6iXB8vbBLiwo/GF8jvwo
sk9wo7sBgLTexhf9LPMPDu/zPggX1VmF5aaaNt7AoL0JhmXCWbiYaXbYPcboNNFT
NhszbXpY0Rs9JvGz/1eVg+aW5Cs9UT6N+NwtIKg89O4iojo+x/WcaQA3D7SqEj3r
OJXolUfgkP9T/UAKByDGGrQA1g5tEbSqmpkQZ87k+5BFoOqWS24z2/P6EGA+Y2AD
I+T+bGuVKIgxnz0/DUPpA9GEUVh0h/k8CpfLlSTl79zs0O7M9F2GwycJrUfvua5g
+xTjx+zWRW88f3deZCGtiEHWlJWiru2CAGdPFw2OeE6+zOSw37YEIx1cQC9ewoeV
mmLTtbf9TDeIlP0g4WYK7MjH5CldmhO276DZodCaqazQ7w4o1VUjd+/sQV72bh/C
84/xK/eFPqFNeIaDOMYsCyXLuTOQ5Yod57TU9Zha2RmTGftSQYA4E/piJcH08m2I
R8eipFLuwsM+XE5XUqVdHY/8GUHZpw+CijC7Mq98ydTRsROiYAM8nXkqRhMcLZAG
s+GkvBY1sDEnV3KMwX/MQLc2hrTWCQoY2C6wCG2tlDnO+pOfsIwal6ymbFSrCmPN
aAQiDx5TxkeMKdTgJCGene/sbbioK65V6h7iHO7m55jVhvDcIoKCkdY2pzSXqA22
dbXZBJO2LohWIXgBs1LozxxHyRHnbvevNvovQf9LTgEm4rbOpIa+WP/9621FflMb
a73qyRgB2MwGHbb1y+5oDqxQDH8boqQC72OaPX3ysvNXxPFnz20jUpxv5nADWVD3
YcVMLvSVRRguEHYP029ulDYgtAjGADvnnDUkC3emnpbTImod7LngwC32YbvhzZ0t
DHQ51KqdUo35WdhASV0EzXCjAZELXh5GEdx88h8GNCGvII00xRm6og6LQ4g7vEkd
QMrafjKr/2riZLfC9Zzu2Xn6aTkqAI2RY/5FMXm2ICYc2TD3BAVKV+KyHCS9GEn+
VvWWp6P3Vu6bwVALng5QsBpjq+ML6y84dpYtwb7i3SqYq6MXez3EGdQDkTrDR1bo
XXjLjtJdZVIod0kCJ0mft7dqX7YRjKOtfSxTKE6+Qyzj5E2e40Lydbk13lGTAfQl
pTRTOA8ICUkmOlWFOVmUtGjqel7sW9UZLpBYU9LUcSsWmTuV0c4boHsDsS/+PvMK
CjuRWSo/ODvB6HA1NLxu/20eub9f9Ufz/n8v2tFj2vTLlaDaHmxPL4e5Ektoyc3+
VLrQRHSaHezo1YI8BdZOMLnI/ClrtU+oORrDDhp/2dLBnVzmad07xGeF2571itmV
gopN25oe1OaktTR+yQZWECPcHNzJ7FDFzpDkl8p4czzR43oxGLnddqAO5TVv+Kl6
l2pxwnp7k3dAdWcX5cjNtl4b0lg7IlJHFloYEiGPyXNlFZS5WwJ+rkfxofx/i7O/
IC8A68IwzEUiq/Jpsb4dJRTXx6xAtqzThz/+Mr7+ZD5JsPKkGNMhlVQWkmKaPsAw
avSwItiKq9iFzbm0uvCOZu8AYBX5tkzo0db11AP7GLdILDHBGyO3D+Zxvx91RSOA
jFI2Na7jj0BhjjB9+fA5eSKIfstQOmEpzP9GPi2f7JON8QOJC/HT9NXFwVDGiedV
NAbcB22Giv9yUJEdB/S07dBchP6VtGI+ssnmS7hI04mr5nZbI6C2O/iKNQYIqawH
TDiR7WwUM3tT6qm6h7aTOndtmXn7LXb1Oy+b98Z0SWdQDeq6dYjfPAN1nETfpBYk
9R0IWBB6tiCCCi9HsRmwH1+CgKxHzibTZxaNBmZK3FqY/LIzP/Z9wW+EewwnQf3w
brXZbauVpsZcSEgRAQzfvTfNYmIQagQwbPn5+0Kp2velAVgKCMVSUZA8AzM0Jn2B
4h9w51CL4kzigL0SIlLCyL953S7C2xjjuTfYDOkjNjJhHRt0SIT2y8jS8zKtrp+H
OB5w2J8h9SsNhopcLwV25djYq10TG57fy6fkhDiLYKKI90cwQY6GR6YUhRaIXa9q
vC3qBAF/ytcLo2zKpbbEan4fO5x8YpnE0n/JndU49G0Ew7w5ZB8TpdmRcfliRVsa
R6i/GpgKq8JtcWDcfbuTeJwYMGuRHhzxim2dTM/y1roZ/+fkjup/2iDFLOlJFDnl
T+xpEs2NVsRCeMIRzty4k6CZI4OjfaHUW9CyWDk20CsTu3K77uCEFQLlLhb/syfB
tryfRDgWMG+vJmj+rpFhudm5TKz5Sz740Ihpl1NYtlHCijIPHTvUPSbg7tpjzyRu
GqATY2a0H8T2YswJISbrIYdG8Yl+bEEX9ZBEaFf7JtF0KTvzuMge8GzDC93VqICR
TNqArufSkLH+0/XFZAviHbp5EzORlpV14T9jBpZuFTX8WQTM+fVG8pdUgkO6RUrS
gP3prXJlKUMRub8d9bjf70f0EFNorQrTsQZ7RVQfTWXnfMN6ZKQRlyCxO3+4d3qg
VUcTzILT+vzcHjxyAoq3mc7ekvPDdGGp8McnXCF45qerHugK4L9YbNf7gVrQcmmX
jENzLCiRyiyYMZXAHMHlUSDvibNPP9vuEd6GzwtLbRnAuw+QRZqY7BHsBOWcWaEC
aBPAk4IG9OKAof2jlnWAeHy55ySgeCAT7NsJqqq8KgjxG6XjCUfAz3ExI0d10SXu
QyLSqKC6Y5/kYXiSy0nBFZpIr6LItZvXRgy5+Tux2YIPKrxrsULoNrfeY1CXeVdc
wBIBjb4jiKZHHWgNQXoD9ZvHlQ8NMa0g+qzEuC4G9ogF1/10wmWFuTT3P3wxXlLP
7LS4rQY4zgBrx5rOejOe+t9q3sj+Dy18dPdwoPrw30f2dFizqrJw3e/AXt2xw3+D
87/cjRb+YDbMmy5fZno4b3LWmafFvPPr8HnyIV5PfpC+oPHbCLEKIAy5ZJsoxqIn
W6XKdcJyFJDA4EW76qRHODEZEVjucpfe36UQ16KBlvb8dYmAXJEaDmEG3bS17yFc
EDoQ3muvp4mdMTmLmA74zawRVCkMbB+3EQ2rh5uFpknjtlTrKAK+8flRGAzzDoX0
anG04xsT6BobWy7HGRT414OcCVEKLxPPcojhql1PpxZCigNdfKGiXtFchMhziGlh
lmouQrxKZH0P09MX/XtCJafFa0OUxTw5GizXTuMX9SsMy1VUsCYJtHceurKX/bme
eCxhZQMfASUQtG8qjtSHfScl9m8beGjRDovI+S71+D6QHjm6kAF4QrxIqwZKntgb
WGAttHVkkduI12NwynmPUyLvCfcax43B2KNrHKXVoQZwnZnSPJxFYknBYLRuGAoN
Ru8fSEPl+G/sLK0OUaQ+tjlh2IJuxIhji8rKTOvQAmUaZ0F+d0h8kd4KXVmW/tDf
qFoeQfZ7iTXvqnrrkkhGlqEOoB3uLBlFSeD8sx+b03b02oaMLACyqcHfcTiK+u0j
FEVx2nYyH9eia8YQHvrIMBWXiT6SsBcsRLTVn/cZx3Lpj2cGKBBc52Q6Oxj2/ysz
iqoZ3vX3XatOMkI/zsvk7XiKCx4kibfuawk6hD0fpunoQF2XJO7/JteUN2eHlA3s
9rxWVkPM6cNLNFpA+VaBAavSKQ+KjW/Qejmu715Yo3Vuw2EPZuPnrLrzfVPs098z
SXEkVSuZpL+btGX0979qjQsdGPS8Ms/e3HLY4QU+zzGXvJwPk8BbmsJKMsqXE4w8
VmIBAbcQ3MGylZCcF/dZLXI+i1vyoTNVzYrUImWpjNJ1tuVn34cNtbOetRMrui8+
xLbfm9aXj/O3wCbJ1hrck/8m12T18l48s2FR+ZP1Say/uW1xymEsP4btDZjyzYhy
8f6O9q+36Wk4/Y3JcP5kLF6bTrXM78VnySosdmCSXuke68KcYvMMAopu3tchc2AE
L2KYSzbU24GelqCHlnUB1qJzGUqo2Zq1xHptUm6KDP6si5EZgJsripnzLfT1WQyt
rzPVzGmWO/xAuMoSASyKYjItN0mNP0HFkDbT50+CMkebvox5Bp7HCBYNIjRY80cd
Jbivm94CjNA/rfweySSMWKzLPSKZSM7sbEs/hwk+vpNzbLkv51K+/GNkdLLh/Xu6
Kki8UJGu4Obn2bdNeCXBhlFYOFjLNXghPkcMtutbJVgcEjDy7ycqc0uwJOwpWpev
T+uarnONFdkwL9OM/cQI8IRupSLwHCnKVAK8uDkrskGd4Yshs/rRyRvkyHWPbh4h
H05kgB3ur9bF/p2A5Ir2xjz/cVDDIst+3rT2tF6jn+Vub+0D8GBO16Oo4hhS//XG
noGvCwZ5LGgAqnxuPnTxD2I9gC/RNNARmWJoOzGgSLRLq1SiPT7ud5p0xofbybcm
2nFuGeK9maYICd3UzAO0JZlP41m33uh8lAx3URi9w2gvwIrQ51bHoKf4WHacOxtP
s6HgopK2JP6Ck3lydXqQ4zZwCsZHy2wcR26+FnwcbV0P9ym5szfA/xLitv29cCx2
lCICoYXB4hBVwHu6GRi1niZ3iBWmriHRZzMl3V1dXEEcwxTMuOKQL4lTWVBgeubM
P7MNawvB8r4d+mTXdTFmnwBp+Qt79qKNOsGChToBPp5Wcuc9wthGbNkgbUQqOmwi
lWexEk30Kd4rEwUCFnPigho68O9mfEHMgwNCKwDKslgZaOAAqFaI0Oui2ufC/ARW
n+nu17joygdZ4+7ucOh3CSauNGtE4LnLUoM8ewonScb9GqEOZVv2ZMtyXyBdV173
e9g3KCixqI/5f+RzHS7a6BTQyXs8T0WbgwzPx88qC6zeWGeXNyuNDwAyF8nMUe2/
vbmwPnbfd6JZdZsakWaY0ce8yYyMa7e9JJmIkTxdZfjJgElQIPNrOZHFOlTcrf3H
s8zOWc1XGW8e5YvYyx2zTpPLTArssu0hdT2qoQzuMxS3iBqYu1wUtf3jgDkABCtD
HMLkLzBiJvnmCSD4cEm3fPXt9Y3kG13ZanxQZXD6eBwi45uike1MXVi6rX2mFoB3
Ptnh8+tLlvYy2VEqIxt7V+NjbBgUbJzxja8FyYF8xs6HsOVpHtkwAy6VAA5wmb3c
/8VOeOMqup3l1wWE51u23dGS/LCWHe8NosTzZFrruGcadT7pzTHirUeNXD6NJ3cL
S52e1T9Uul2LISkICOrclsDw2LhDRr90RIVFJ2/mUWNlSztnSGn64KfohVxTT428
jcUM5JShztK3PRwnRxPn2yrOlg8cCL/HQ8S8f5VDuNHO9viPgbq8sDbpguG0YlaE
r0uRHtAHxerckuYVDaQj4RvtbIVVDuPC/UdhA/XdmKsrXHKGeFl//86LNcrtO+9v
4DseLhZ84TCOwKwavw/R/kAUksiWMkVg7QxCgFURj57BmXgMmGq0lNXNw5eLIyjE
TZ8yo7xauzCybK1XNx7rNSx0kd6sCpmK4lo6+wja79hwGyXVDIljO32a4+yLBWpw
IyUrD6Ampu955RnAEnPekcfoP/pgErE+vUH+0aN4DMtsev9H3BtGSkoEtgDJhV0W
ZsTCMb9LfsZI9Rfg3p26uuOuGPo7xufxQQoy7KHzZ9yRhStBM4/ncPGPI4bANaSn
sZByNYC6vnT9VEXL4x6uPcZM16Rq46P6kXfv1XlANVrRf5y99HF/vYJR9dHVa22d
GzKkRzsTCUqEv3YaNJT+Fedw/AwsuVf5appwRe5TJSaDMVY2LeYzn6TJbsCq2onU
aNNB1FNIeX6lGU9itRCVXtU5Apa91Mv4uCjXpp/AOFm82chr4fuWsM4YA+gIHutb
H5iOBib2cUmMggzxvEK0IVyRjQbTxmQvwEsyRvN2LnKeqEOCodtEZrfm9uYHl51h
s4R4N8XsWrv0SDiM27z6jSiZ/rZTdxtTyC72S9C7eFtNG6YENmy/MFVjTKup2TPB
DiYDZDv0+ocQtrGrvak71zcBAFxRksADgGmL2jMgyTNdrGSoEN3NNHPjnvwpuw/u
ncAotgHKfp3Avszv2hrn+ZvZIvntwKnxiWIMj/XFn7amM/q1o+eIMtTb/FX5HpV/
ZOLGuyulzmrNFP1Z4F1OsDvscD0qCthCtlZ2ob1lF/uHHtUNN92jhDX7UEPOvpiR
htIMXKSLVdjbnoev2OvJO7yKk4br+8oguxJ0L6Bt598xBIQO7s7wXSgxjH0/72B+
r7J6BbriksjtH5XPDgYYApA0TOfj69CtYdRxcNak2OCiiuqiFqCRQpScKBbkY46J
Q1w1PSCMaS0q+uwzx/HKCFGp0VDghNoajQtqlCIM4LSQBTyEOMrIMUCALvh/iXsq
ocPkIJhILeJZpIHTGK3YS7hHwaJDbxztSX74UlMfoqu/BwjOihFF/hEAr+BhIMP2
n6Bwxeg/SoGcGrizQl5eU5nZcQinpuPCpvwuAVgHi9ilVQzDWo/c+ZEIabnxrBSt
jDYmzetRXK5SpAc3KhvLRsPyhJMyoem4ZEtqOuObyf+4Vyci2KUJ1J9EjTNduN6b
HAWaPaftY4JRIUuq9O4lGoB6Q1VhnDB5C3Q5ExuvkAMkoURd+a9bbn/OEd7EZLe5
z6gFKJ59Hi8MXz7U4jtY8CBvRsatIvnzGN3K5KB05hxD4FvF1nNX6QcomCEaurqf
agHp3Bn9OYKwS4euDVpCllWag7N1X3h/h7FcV20mYr3Y6v0sxjt+CBjomOWwVTg4
SbzMpupf6wwG3dogfpjmGYgUDZFLgN85t0dVSa0iMqzOmGBURdqzDOQeaniBECKM
pm78a6e46jfpui1a7pUkxRZAGwkZwxo6Das7ScLCBHygKQhiMPffrwk6AsGlDNWD
Sp3kizS1OOf3BAbIYytP0/DKAIo2IrEOsi1puAIMgsWkYIcOGw8YfUuLcIJr+q6U
p8IjdNmzu2dbyV5H4YRWJLotnXBV9BJ1Jek74BF56slcPaEp6UHp27LroGryDIoV
q5g+SX5qtxFGdXj3ineu1RknMeEgakqTgagcSOdP5hVK2YuVjfULMN1ZXJPftTkj
r4Kl6WnQ4RU9fiJuOGaLoa4kmiQy5Igmj7U9jIsJIR7fJTiY42UhUAcmAHjd1qa1
AX4tpKvA4INcpEEXGJrHFWTayKo6kVvcPi1+hiEg1zeG0tilGGqW8lyreSCtmaNl
9/GjGf5SP3ZAZrdFcNxyHtX4iBh7oC4kbFLVlayqjNGwLtGUTZOCPdCV2mfL/v3d
YV9wWI1/CZVG3kXLLKr9etJPuuLrUsv/bB02vscWMxNengqDAf/mP002sPtcU2kE
Ppv8kGT4qLTMbcvaz4xCBIK4OAJync3mGDksfWkDbcypLLm7wBAdMDHdRc7r9cV7
45yYAxKUPnQ//HhykjXdhWBuDc027HTYYwmcTqSt+g3KWrzcjxAM/z+mNhcnqWZM
DUeiSDuIxNFlyHyzjnnq2d8eBKlddveJ+UTTj4oixSH+NWkGWzAaO5hVmBQNGTx8
Jhpb+LdBNjkw6qoMqLBjwCqNxPggF5LMeAYhYc0TnN3geGEuKUTM4zZEqjbfBkN8
HwDUVW3O1ZyCj2KXTv7cf90DN5P97n6nBwuwYKFFXkxDjBew2g0m05GZpsmEU/JX
WrJz4OeesMk5ehovJMM4hzTGJGU14L1QU/I2vMc8PYi0iNNqEEXBh2prawA5hNTl
DMytm00MPV5GP0KGol+PxNoSLdZXIw7OWU7t/QhtTWeGKxrUqEazy0KIHk6psqvl
5vkcuDn6QCKIShDos4wkTIl9zP5XlwzrJtevkG9/l3Bm2vj+RAngfoDftM7GSymG
bkjld8lFR2CVhAcpEZLTwOM5bcFnWVTRPKuGokwjH+PDa3+FS1kvjFNPb2wQDdRV
r+dajedsPuIBvGtceAcLeGa+SN4SxdAv/I5W2pD7G7ZhUCULb+ZeH+sZfPfY7TtO
nefsvD43wOkDoQGGGa8Jdrw0DxN23HeFmH9zo4/dd8EcT2g20Us3guJ7hl4KmiJB
V18a4rKGKICosFsDzU9TG8tTNhToLgqBAPNrzqCfICQmOqEv7D9xI/xZYc+MQQbj
f81hD2NqqZLUOxjHwT7M3TJ6WRUnsUlKQGClIhYgemb0B7sh1bRbOITC5yGTkE6h
aOCVJ8OaWhABQzWT7A+XRQQP8nDTNGBY70xFxB1x4OZZhux+KdkyvPy1Xgw9hsGT
zDOj51MykrouQmsxY174PITzbA6ETL7fA0vYe5lti0zlYYhDZgEyrCjCDf6L/zxF
6z7wS6Cd4lwY67iKSiKTHqWrkpyMdTHNNbtKVgE9bwve+Bj+Nf5qaz2bqAfOJddu
j+GHOQM6/wrSu5szuErceU2ZyfKBV7ALZB0QBIzJaJKoS27bmUf5h1PU5wt6vFc6
HEhRhr477wGTDYcyegDTTfCYKUpaionK/GzYvYMn/HXJ5VKmsqJZjV6BR+ReUutb
XAozh8duj3EHzFOSxhvL8ez7mH+3rcyMfOvUTwyBNJa/VtDQ0TP00XWxyFAG+eWU
4KgqAZKRSv+G6We7YDnO+0wZwZr6zgA3q6nccypEwMd0DAfAp3X4udBg5q0Ma+i8
52SAGK9SSN2lsKuhB8AWvpdFaMgc8ETWGwij1I5gpBCLhLbHoNlA8Du1sb//y/Rn
X80KB4sP3CermcWq2e0JkkOkGQH6jWam0DQeDQaTmrdHeUJU0E1FwyhDPj/i4lQt
g/vJYnhZCKt3VUqwEqdqa7XwSxsYa6QRhkUcxmd51GgWWuWQ2i8T9LTIEEr9YAhF
HLHEExCMuEDEEggcgZnnj93w6u09FRcHLPMPjsymYTrhPFls8EbRrnCfJHey1DEX
kOtzU7CuJiHwHcPG+GsfLz4tGx29REv4wm4V4RQLXYw4HnI/t0vdGmZlvQJNwz2q
pcdEfjuWEbOpiAb0ZI/s8cwKHBrM/2MvaxdgBv6McuDUyU8gr66Lt5g7HZhprfSa
c7UnxNdsNLSylxlzMTW+cpFI1rnOJIKqyrLjiMNlgaqf9vK4272SsA8054D6yNUN
+nSUYwdlgnYQ+LxKH1bu8Ntm/MDMFYBZ1ru8YTJTzVjk+TmDG1hdiPlk+AV6ZJO3
1fnJ7Shin1fbapLkUXSh3CSkNVcMj8isp1cU9JVJjoQiZrqs6tghn4QdyZDtRvLe
wdd4ter83GGesta3xKJKuuBDFymmjtKyz1YHRDhInxg7qQdSiG3QT9DMCIiw4Kzm
EUeXspWJlTlXZrSd1rWuMlBg1wmLcrsudczlU6GfQab/QeNX6hPQigNfpUp4Emq2
xFz6cK6s7YK9w4tHnfhn2n8urWmAOL+0+hzRQJTWOvf/rly/bx9cejSfqFIXMUfT
heRtYlJP10FbsnuUUVBZJW2MJ484KJast2lOSIwFu7VBtAyz43/AtZ4cUFFZC7Rs
JUCSsrQREqqtE3Kj3AdpJk4JajTsGvfCtPSRXx/BhOmxbci9vQjEgoL4AQe+nOEB
vSh3Ouc/mAMKpj00s5yrfRVR5TO1rLQ2Ke7jUJxMUZDluQHSLOFTriNhxt+slieS
8m8wvU0rx1Ch/WTvJIylRi+lOuQhDvjWT/xOhxaqrPS/hSBjfrALtLzdHbXT/O64
yS3VDGy5wrecb7uwPxb90h1H3rwNTlcf7xUOyMlWgdXcG0IMJxROkOBXxgTeQ3tZ
iLywH1nz6q86Sr4ArE3inR8vRRFGIeLxQXkTauEbTjbJ9OMCFd+ADq//jVJb7Mtx
/FD4I7g5uh2iUyGTiFvimCnI3U0bFb+RZwi5VBRTJ8ceOYrCfK35Bq2Oe4BwGYSH
5e+Xbvbp3s0DQNN/DjvN+3e3Qcoqi8eaKzGNSh1gIHHYcjLJShsOp8ifYinjGLiF
xjCh4WxbTAPa90bND3PKzK33DDUHA3GHoqytxtFOu+fmrAynOXElYgOOXWfse0LG
UHkx7edM5TTDEV8wIPXGQ0kTcl1jfF1gROZ1gF9MRCvg22cL9bakgG2voWyf2k1z
TMy0pNAKun6nDCIpaPFH2q61BeykACuuglBqp7KScVPSslgbvqtAyBOwZhiiDNf8
A4Jh2xWppTg2iBCuXvNddgiDZxV8INctoV2pm5v4fTY0qvtaGlokHg2Ge0SCsLWs
1+qH5mqqpXh/zUdkCF6YM06aODRN/bUa/ptu0G7JD2TqEkKLhm7iVmE2ea56maIW
7l+f6NtGFUc0pF9ALrKtscMYekctWlGNjvGGOanK5pQBL4d59iszTQdqnbCbjwXy
TUn+La2ZHj4iDc5n4nKEQqf8xNooWvuwDyICQbaHPaa8YcFZm5yn24kzm8OfR9gO
IrXSb7yzXKeWMnaNJcpv6Du4N7aKLgx1OSIKjwTe8Oqq1n2VW+hKPNsBMJLXK1wE
pJeYP6BgCRWaiTtQH1mSU+Le9YmTOyfXkoeky50vXN/CJCSO6NmjXGDJ8/8bFqpA
OzFsTmvrmuwrwNR8kgDoJ65HkGYwJjh6I7h4Mo1nODkEPKRC//47k6DoK6zeYJeD
le7ePKN+0OhHJ9T2QyP2VR1pdYuu1CKzeCmZdDiGKf1HsmG73VS9wk2zPXxFp+Pd
xmFbj5Q5pAADgtS4U4klxzW5bzrEs6+MO5vLD+EPu713hiKYY/idglpwdEGhjDDf
L4L66KoCB6l5CRngzZ/QaFm4elf1j/F1joNlZxzMHZ8zf7iYHxCe/t+VkiWpRDmH
4zUWG1T/PUGgEewuCRkmS9aFkqM9ZW+WQ/gVlliqhZobVbu3GXA+jSA3iQd91YWh
8IE9uYRCmTa4JnLTurjQpTwcPWedWZJ3sKe/mj4kQSxN1IPsQj6VTisfFtOa8O+I
esHxSVOooGfaLE3IIoGdklLf2AoYSFyZcdwczQUN8Un/qb4B0p2P0DWJmD7QP7M8
Wkn49l8OyuLHSMbCbwf2BixM12EhRe2P9HbyyxvGYl9GtvLAX/2CuwVj3dpctMk/
mNJkviKABd8EVxDzCpd9nBfhEq0hzbKWTWX0e/g6CGslFxOGhxF6VoG9VUTubNaS
f5f2HX5cXKbb5zonPCgsC865AxdL7BvdKs+HPSLk13NBgwrlaw0dm9Ck7K1KKNGT
qOW0ik+37Amha2YkQ3XibLhle7yJSQJ6mTY4ih4AM7zdrP4blNtRjdI9cYBrQOSq
TCgwf8++9x7Qo3Rq9Ub5Yc696/1XL0ZSZqt07vw1sc/b+7y16h8ugN4RXWRqNlDy
QBqZYsF6lslrQuXtIkTxJWSfD/a1LZyLEonWHQREmtFeYM9pPtqVzIE0/TZVQheK
crtJQIVrhAjSVxa1OuPKdQCtPSS8teG5eU7/Y+ba7jaoJC0nCG7kqYQfqGX2RYfz
tgt86BTWBln0Ddv2qFuUc7eGy24BoHVMWTFsKXHcGCnMP6de1E8e/9RmJlRUqe9Q
yETCrF0a7xouxiBuesjx6Xzz9K6a78LnErUffAILX6nLWqlhqetlY2RWUk8s/cV9
kU5jfnn+8D5K5+ag9Vp6D1Il8wT1KuenI87355/pu4aFyXWX4zcIsXxytPgUAXu5
vL+j5G/LEplSdm3AVepvCMLk9UwfnGf1gAImPB0p8UyI8zwCqy4ac0UIRISLVDmb
4eRLHVthRsrYjhgJTnxppjCws/rZd4gucB/d6xXccKI9UY8vUBTbH7iYYCEV+2NI
gUc+84/lODYOiuRioW81ad8ykBI5l9WM0CV6AgzGjNZHZVCIskV/14jw+yx1ljSx
bajT5IkqIYEIPcn1ft9JytEptbClwHgP8+Tv0kl3Nl8Rlk7bl5YCQlW+T1rXmxhw
J7y+WcH0x0ClF+m7jhU9p5NY61dDczFruU+jddLHzCXK08JaXdpbapbQU4128fFS
iMcvP7hR/RZ7SnvSn67jvOhOvZTqKJsEe3RtnwrY6CSy+1fxnfF/+9J2o5FaWJPt
WdOuntL9xdbo8Ra0lcQnX0LWVxPZaofG03DIyoyNog2ZWjpNcwHmBBZxRTkJBqUI
FqVBmoO3152UFeDgYCgV/WESM0ngj+UyG8xu5GqWlKkRDqWd89pSztSKxMYCUD7G
dumnkozcxFCmQmGRP8AcG4neBgYNENj/+aab8vMfUKqUfpdZerxo4ycFf4pfgol6
DGAOpYKBnNzBQcdLID7pDlRfpr36jjWQw/LPuaP6jscDqJPu8Kg/dveEsH1anV7c
vv2lyHP0Qdhqptn2x8yqTvr5PRBlvrPSSlDL3vJ5Ptb7mMDRBMyuM6PcWEh/IcJz
XRR4KAwbCKplRipx2mu58B+ynDPiPcKvm2UR4cnK/1rQkpGx2GNFmrD1LZDfP7SB
h7s9wlQLUvFrxg3LBftSYeSdOiLmzWYZBS6ftC7N3ZsEEVkfmimSXVEBdcNVueRR
Os3rnD7rLD7Pn/TyTWjtEVISa4UppllfoGU09vcx+NWqZp0sM00+6jxYCgzvuYNr
p19pxGnwXBBUp/yCFExb5akFhsvs8HU5NG4Di406g1X07j6g3Pi3umm7XT07DUL5
U3hKkTUU+yu7sg5iUIvl5w9YVOeSz8PjJorIbJWklUEmIk48XDKa0HLBMJvLGn9g
CROX0fdJQ+8klPe1oanmOlx4L/bzTzdG1TQMgyrEZh9sP7HWS47x3+loYmrZVcx8
S7tFXWNFL724OpaZxl0TLqTNKMiH5wgg73uyORmvQwVsBfEXcKFyNrRjCq1X+dCI
XwXB/xClRZeAn7f3GcthNvbV1vdAzm1js3tlLdzRb0H9AkAtwMdsWvAHT6llHbrH
0JENET/vfMVtsLwKHnc65V55j7ykQlW9SfiJMWcvsBRpO/1bGR1l0iITa7S5b/tX
+tx8F57tb33JEEclSxKhFwIyzfUyhs7ipbMZx4PvrmgBABkd9bnWkhzkZFy3gpiE
G2WtI2lsZ42UYBX84w97rjTOT5BggovfJ6NfUgksjhBGWMePQWSwtj20P79Zgpas
ACpyCrvuD3P+n/jgDU+aek+A+qGs/MKZYkxax+iJHz6PHFzB2QFqeaertZs9dZI8
bajyqq1RIJBla/ScNSO5G/cLXxOJoHbD+cdxIW8HUqK+RUA7W+QQma8jvjUqdh08
JKXSlWhn+Ynjj0Rx5L8Ctm/h/7Og/wQ7ZaMLCnkclGsx9uDs+AvvHdYLA/uqz0Px
FSipdKe+yL07oxT1fFmOB1oQtyiURPjHr3jWyTQcbXUdFna6KpN6MR72pk3HFgF+
5G3mlcSGh8lInu4hT6dnnfOkIfs0HChtqvOX6eeIXoc3uyBiil7YHHYkrgP1Lgp+
e9J8xEhbE4yc9gfQhM4D++I0emackK2r+qRB/OqUC7qurCtw34KJOupSBpx0igRc
hEerwq9L+sJM+7FTfc1GVxVumbM10eIr6bR42n3FUJC6rV++44UKVUwW6fICdoBN
Fa6BFN1X1D/5WZSWO+URHr9ZkqtSX0KaAxg1b0WJ6GsqW5TbnXvKR4LHlqDKsfkE
L5PG4CKIq38wdS6L4DN2Xpok06Gm80fGKhsMuW6Uls6rsULJY1aH8bCwDUJNZWy0
TbdmV+5+0ytsCdwd0dDYatBKMBau3BE4oGfv8y/jJ9oObLi7bmlpsQsckpg1i57+
gF3p6JD+vgcV3lBiMMGbd/Q+dgwStmN5r1m6qkOdsFZPHeTV+djQetoAoQCdgoJ3
i7X4EifjUzaZhY4GeR8XLT3ibOgvd3bfGP1YzhiyaQ8hH84vil/TnYNjiwRSA1F9
wVCSoRUXTVtHSGZWtRJRPXGqHaGwvxF2r2z6WG/661zJ+hoPTzF+dYmk4JVnvzsG
vRdnVXkWIagvnMGr9Mm0kaRscnMZ7h72xXDTVXi4yjJt5+FEWJsSL0DPYMriXAr/
OYCNcbNIx5U1+ttiy+Q8vBbeTdDK8jnAsdwyi4MdMJkg1Qdb61bEQsPVcG34/1tk
e6UkF6eFU04EFURHR3/bwKxX44QETgWmj4Im5IBR7IQx+x/V/7QxxqaFOxTMhPcD
BJ4CwV5JYbvzC1dt9c2VP9//LhDQ9PHHz+GjIXIxnZ1BmrqDRZUzT72blPpQ6pJ3
2K6ne9ZvuwpMjXeMAzcSIzq23USJi0Q+C2hXfvQ88+NLlV4sganYm39W5oYi2rtp
nCIwjLKyZt07s0aD1yD8oMjaVzZOOiHEQbE2qfKioEceTnNdQgD/VRurFJwWS5tg
HCwM4eoPAJj6NNHWNr3O/NOxfQc/rhYoG7hNOs2dHDTdpZhFjm9Oa0JgVTFbrguN
sJcO1i+2wFmNiV8jYTvGvMziXLCUdvzBQqNzND9RRdwf+hsfNLjrxijlk0LAUyi4
s32RYPv+NVZ8zFV3Ctu4OgdmYDAgnzvbIZJqEpGo3ZEzjh8ZMfUeqCF7haetajKS
cPg4q6snKD16iOtuHg0+GL6zVgzBzOnhLRwbtIQQw0SLNw9T9PYemGuRTnUKowoL
s6/IPCbNzzAB3KjgU0oZ+a8d3lP+DvBy77DO90n04SER3BIcnYD7I/4WuJLYbJ30
dGFEWip7EJBuJoHAhHz+7QHP7OCa6/Yzxdjax8MFxfdMlJqo8hJ2tLCNS6coOelX
DDEy60s4LtY/ueuIlzWI5iXACvxxh+o6gNRi0Fr5IT2vgk56UDuynUkWoV2DvKGA
Gnt5WYOp4yOWpFatnGCCjEhzrMdB1DQ3wiYCUTabaOAyLqjXSC4Fk2/ko/mPvSGa
s3sSW33S8/he5goiwUfgGRyDFAlEtySNBTEYJgjXO2Z9lXAjAnhiJvA7KRt8xdIa
/5vB46E8+jUm5TgsyG+L/lzLJEVTbK2alWhbfXFHs6tuLHkNhxgeB/tAV+M9mMsI
vCifyjalC9w2Ejz+xbj7I8IVGmiJx57LQUk3x8fSx5MUjw3qljOrLAAJB6bX5mKc
wwDFQOGQPZSvoumAdNGkyFj/6abPijSeW3tB5xEBxIIMfOIMf+9H2RaHJ+kD2asV
DL1zUSfj5ojVZYMPLtMlt/RMtK1YeuzzbznbdWDlE+7YH8fJLJ1mpscmtTPGO+wK
IiCntJ+qkmG4TqE0YqJxGpsPZDGowYKo/OncnplxrVFVKqhju9qwJv3qUp8tUh8V
8xyhJo6RsSmbmKHtY3NUHtGVZJvTHHArbre4INCGaR8bfKfQhqEQbggNos1QP7Gb
oDV3JWsfq2lP9VhWhhLQhRCJ+Joj3FxNmPs3ifT0dF/Ppwi2sR1aVHB3mtPkLkq3
PTeDPQgxw/0yoALGxw3KGG8Ru12vYBKtWokHEzLkhR7PmIQaCpieFkpXXjejqxsT
s1Tm86i1SBFflg/2SAm4O6wLfdBz7jpAQMdZZGz/hGIiBey2FQixg+JVyeSZkuh8
+vltUVytfphkN4V337IVsvxKJHc7qayksz2UYoqZbYylRaKAT9OoRXJ9cnUoLnQy
Q00j7NzBDB7FEGVjlq2acyoKBaNkUZe0hgiy7c/3ZmH4CTZQmzLYM0j6qUb4+iql
EdY7jAiPISojfcaP0NbnNJFKgE8iRLju7sfdfboAs27b0fS02kpDL314aAjv4TtF
xpCxv04blpkbqAk5Bl5uK4f+N70s9+E3zZgq4VLHt52H76vLJ+8joycwhGUFks4C
JfsJ+N9GW8oCoMwpoAJh4vYW4Ue6qHMGWiKav48zWwDX+FuWBjGGRAIUwucdq3am
ymr2bQMTYSZgsqz4OJKVEpf5ithK5y3XkwcmqsOSiWIU7JVCyIB9zFV6myFzEpCT
StR/3jpNA+75uv0vuhi84PF5Rq4CLCTgh1aewm3KO/FHYz6mQfOecLfJwgQdV16H
WHUoICeDu8rhSYfKXd4NxVAubuEt0x59HUqEpsjBrs9rCvEidyw5/ho+VoITTfQR
/Yn4ivkffcfsJ2BAvmN6ZpgkgsLRwYn0YOplevdikFLIiziSuawsk7lTQIejFvH7
vjaeALM9hAH5ueyL0cqDqPsNLv3XAUtxNh9sZFtDAVgg3LMfk6HszTW7YwI50gHH
JMf8KrJeQj4WZc3NJN8c40r/xCxg3m1liF09MvHSJ7yfLMlGgyAOjI9tJhHWx2sG
wZ0hzR1YAEawPxsGypwIZU8Uq9jn8AWY30ufYVV4XaOUerXQxNtAX5lq0c5OkPwM
i4VMUbaZ0mYInVu0HfLw6ocukQ4JkadpjAfSsyf9Fd06NYkrMn0L+mJQozLwRtdR
Rf53iK9GzhyKb56sVmGDRO9yD5kggLetSCcqPpbn1iygN/HTLJDXDWQItH2jhYYm
pOkXrIQqw2Qv7XQdZh2fz67BoK6bF9nZ9LesmQ3e2x9fdTJN/x5yELqiuV4zDoht
nX4gjUVFBu/WqvuwsuT0RkcgrVFHev3zTw21Ra5tT1uQLOn4f9FYc0u4GFwtDsaL
wrE9vQGIOyjjgnQ/BFFK+owQ3gE+yFewSSrZ9mc1UvR1ALRytRj5A78ao0FYlrKh
/NKxnNhjNUdktT8hmRq+yvIc0YpDTiaP2TTjmkBV5BKwtbdP6RVzP4tdBOhU9uk7
lWt1HdEznBaVfcub8US3f6gDaGpKnRykgzESl4tERViEd3PU+yxknt6aLndEvgFv
wgp2H+5CSXz4WKeNjNquS82K0uB4P/aR60yiWqIJXKs9bZ12cxe5xKARAfaAPU1W
1F6VgrV5E/rlJmLEv7B4fq9abvLSy8C+ZuEyKAExpMC8zcw/cMi/S28lxltZfbT2
EozPDK1W9b9bfN6mdNrmHW1U4/faK7xlBYvRaQVGokR2bTaV1Sz3w8yEExvYRFQd
QHdYvhKSSvrSbj4ga91CgKK8dfM7CN6tPpnd1o9ndzotDo6q0HjG8w5CG5+qisQs
VcdVu0MI+z7Ipe8SVQkXdQZqdkvWwFkosJjvhgj4/9JBcitklgkZJJCvQ45SAYTZ
EgyhJ/xTOTHRYH5/uxepQp8wVqAgrPr26SsKugX5fcm0os4PH+lsa4NB0zgmP8Bu
N8sbpyac0BJh3j4/ktZLaUSkXA7ZnVZPXRcdtJ4dD1vD90Rm9PMzqfLWIReCboGl
y12bj50+E36JjgIPbF7mGBPv/GAxVhkLeu6epxEouOZgZ5PseBXCIPtHmJhpVikH
b41lqQX95lMCzGUZpmHTUrCzxFNWgm1E6ECFNpL6XPDw/uNM7cPrggJBnMPHEG88
mD0ToFvRbuh11v1cQNI0GgtS+qZBb316zflGT+9Q272DT2LELnPdQSO3InghOniD
X06Z3QiyY6tqTBltodsgZgmSeRS+x6nt1mvdqVJNNstfM7r+XYNdVJmjJ5GE5PKA
6WYKF8vHfWvEQrG7xJJvha0X/Rdw0ncbaEPO+aSQSP2o0Y0hkZ7cL1XEn3PMme1D
w0+I4lUTeqRGjRPIeXXUSY1YuuQShDr+bSVQmvBYRyaOGpVsXkoqTzfdAwTGy+ZT
c60R4+V0thyeIo47jCqkr8ASbk5h/ZOh6gifiJOcC1RsOHwguHpyLUcFbq+vkH/D
R2u/dCyTlQBIgYf7xffCbvjxB6EKlbVL3pANXipFTGrqOiRYP2rH51dqCa8L+/rP
9zGYF+YlC0yyNrAwV4ubFz89sk+UaoxND2yqZB++n8tBzuuegG9aA01asr90406S
Xcg0SxVx39qNemLDpdX+6FKQXO0shqql7sRkLDZcGBwC4Z8YNpNU81gHmF8MRtIe
+q+X0nFjCv/t/MjeT3MY1zGv839Hl37w+QxOX2KpFzcm5SA7w0URqgUkADloch+9
9CdoHjn2Ex6Yb7qx/FTxx1nYLVAS9S5H2AmlGt+znO2gWdXWRxnAfvWYKZWiQ2t0
AtgQbWDuHypXWjKTPU88RtVJRoE6kGtQgySCj6mgl+e/cTVuBrsmTqBsHrYK0VsB
97z8xT98QqewVEXc/mOwg/69TLBRLPkcRxL6Fk1vb56OXSnITSiGxdsol7rNdX63
m6tuno3NUuAhB0id1LV8l+ImLJ8Fo1ypylV6J7fUFNExr4myL5sZ+kKSs5Yg9TAK
YYFinsE+4bK665PBEibZsgc+agl8GBJJShCHNfN3hwwiwQJbZdCRxQKo+dU/Qaek
s6MXGhTSIaLDir0cBHFHJi1kafjzBcPldOM0pSImxr3oqKKFn3TKb/xT4SY52+k0
63oNSdqblLjiuVVRHcTA6feuv+laMA2SidM9oS/IxID9If72oh/AKGCiBPslXnfz
bwDNOYjoQyxEc3wJdB+MAM8mETAxTaGHJa65ykRzb6oAQyqTFKHcX9GxD+LfuyBY
qEPt6CcW59APfjyeDsgHG5W5GjwZ8hfn9d/Gdq1GQ8v+HWc1oOfnNzAWkyZj7IX0
RHhbL27x9ntGjC843bwLUjoX/xbZG6lousRFpbGLbsk0dxcH6Qtnin9LXyFg5mV3
RURKHYgi9uF5wBmPbnCPqUV21Eihwb6SWjotLhiADT4fLR1N1Futxj6I82DEFcFk
6vbEPb2ndWntbKPbd+KOT7XK11tyOSC2aBbbYrmpAw6bXRCRSvYx0Wf+ne6F+iKv
MG7I+f2psfblyaFK8kL+XOr6ax6LunexuVw4CWJWcAfKvOMjNBn2poc2P6KLOAvs
v6rnWt31BmupY7sl04O/zjerZVmJ/p8TBsoB8/El1VlQsKNEUt4dIqtt5DMLJjyh
YAN7TsGvSlQFaixN/SQAnH3A1UGHvjsgMNvZKdWgNsXjk0vw8++e0+FcUsxgU97i
FQuvS+hA2P20edYuoA4EEOreNGIi/TD6aBuxUk8sRuekaJa1Ya9ss5nnHRJ5dnn8
mMmnjnZLcGnT/UdoCV9wY33zX/jGB6XC+E3t2b+x10pTeCbz/UbKhy8GPv4nJP7w
77/HB1GIdQeISifje21eW2ilQUqg8QIUAL972GohIuIoM3Azl4uu0TEhCBhGjsk3
ZH8C2jbrLFuIFsU2Dd6ymIIps2NZqEv7wdPcoIRJC/M377ZU8/sIoRycUnuR6PXX
Pt/1mrzYxxSLBhT5gVgfj+IHOMRSzzvMPWXD27wyE43p/qyxl/XePCbSeIkbl2tw
/lbL4yTnLf3JqhWYq/TYOXpc91SiTGs9eiu/eTNN14RBfvcMJ5n5xM/63iBicoWD
pb9AwI8YiVtzvH/p4xY2GFRgEpjCBVyRmHVMdow5KH1R/S95Ibz+0BKY+VWRD2bn
bmrf2eA/ru5TMrDrRGO/ful2hBoC4Dz59zIlJP23KXnpLWyWBtK30ngaYP/B6G0O
Ez+Fm9Rq7+PXsR8NlVG6U5fg3SYFVkH2V7nftHWEU/sRsj/1h0sr64TzkJF6IurK
Fmm3ARSIiJQIY9bMPnZerQLFcLovJ692YGUsIh3IplWqgGVYT+AQNoNH+wEygtfb
6v5VinGs4rMdFkgEu6AgxQE5+rZsydPyAtF14meGLDI4fHRWJlSMAO3iAkadIvHA
ypFM4DHIcxAKl63/PI3QmCPV5z1YOEa9xwsTjz2v5vHTTvzc+NPzH/+hWNv45Qw1
3/MZltkAeADcz87yyg4wWL+ctEIed89FGg+bzbO8hGMJhHYpnacdz2wSOm6aDI3o
V+Jpd10Vc2hulVUzQLDofwEhpDYA+Mv6hFwjAt7Z/UmYoAkyVwppiQJKI5HpV0Da
aAqR2ybY9FV2PkOrhMmGbtYq/2tnY7ua3F0eZSyi2r5eMTgX7taDmomGKGbPiHWS
5ej0KKWnVPierClMTnj9BNybWw0GNw5pe8TS/TV1kaxYXe+lJE94y03jU0VjSME5
gxnNUfjjTWiVsntUSbewMVuZjiegp0KKWagBiAPTwRqh2Cg9ptvRQEF5S8xBrlkF
PfYsyHKUk4khUIUaHSocKzD99nFIf1fHciqZmbR9FTT0jyqBhnj2iqphZ8Dr2pzW
FMWVlRgQjA8R6s51Y6KFGgS6gTbI/eOZiXAdjvGXSk7R2aIdVr7N4X++R/+LrNYW
jUykY1Na65Fc1rc9u7XVy2lj6xIp90UL9jdPWWsJHhTTe01zkNnJwoWymWa4vdkW
2r7qTdQCfCuL8iZ7q3pNWXAbK5ZoaAS8d0WV2JNZV9aYXuQH9fXj8zBko6f5PNGg
A4HLaBd/e5H8Vs9aMLpQaRKUsPC2d6uyGDvK5oNbZWq+fQhwvJFtRhtqCErt5jz1
WMwPWwtRVYjuZIaZdV2eCHX4Hx1aWPn14kY+qrLK1Gny5mKcbyaMOaCsCoO48xAV
RW5y5Ug25a9BnKp5LiwH+84hqUFMEmKwBAd/xdULTHK39moOSwIfVWqDkNB5p3kw
P5VrlyAxWFcvDj/nzfX4JK3QdliWFWKdKSpFv1/tW5N7ihwp7pZ7Mywc1KQ33Cpa
HOp3uVHuXTBytgENG723N6HWhhdCocD08CewIwnzzM9aIGST06MXv5MJZLLwd1X2
PkH2BvC9YBnZq39fCEp0dGzu6NP6QFB3Zpebx02qxWqeD7Br7tLtYsufKec9ZU3f
VMqisIxIvHTYhGFBXqqtSEVMEOUB4dbJvvX4WpPsTa26LDx1RC0sfHevkOPa9q7S
IOoWgmjeXYQwapUa5sRVghq6AQLvKQXfULQfJt/nk1MP07JzqlCzILr24BKXL+cd
Z8ctmNIGOTdKQ61kv9oOAQR/64rf4ca7iI9eVeljKFfFsIugUQ/2TJuAIf8aR6nC
nPa3X9vZ82mD+e19q6Nej98kXH5HMPHKC8vVO9O4Q/RKWQAn8gCs0sPueVDaGO8h
UQqlQvaTwiFSs6gExxjTnRoxpxW47D8rZLfwBbRYwtl+91y2aBCVFjOGRz3r68OC
uka7BeWM9Eak5w44ANUT1kxT1g4QQpgJpry4CeUtfBoBTLXh1O+WqjCX2cm1NPjF
MusPcoIniZEej4qCMUKADfxldDnVny+hCDlUBtkNmWIXAewGp8r/AlHoM6zdILbP
acFVdrf8/2GTS1YYIULzEDKtRP/yxxtt0n05d6a0uOuvXKy1ObfMK8JvV7M0kAjt
yIyDxBoAI1qnebB+BO8jdmLIayMrwbFA1ijuXAfVOj6hnXGtRVtUJNGcOJjfyPBj
boV45RrP5kWXtiQqyUpElfHwtNtQ/XK9eL7J4OC3gUdA5dfcPluNtUrKMK+o2Vyl
wQlX6cev9/3PtAUI8pcQEsqTwFbGwf4l68QOtUD6qEOlC74dNUlZZ3j09fvPfTNJ
yllv3JCgx8JYNEN59dool+wRcvDtH0uFzSnQKVJ9y6ya8S+2NI+Uf9hBZ9rd/KlU
Me3KW8aoWVLOwKyQowNpH8Vf2dw2NiYcw6B3VVg0StZSaqhpwh5wUYNE4xu0Xxc0
eIDLolPiOOcwymHOuqNsFacYhjgaDnFTO7QK4+5ABcDTsa9OC3Q9ikgeHOhr6XRh
Ca9Qu70m2SU8sLdszVGESAQ6iVoNubHl6ni6WlaSRBtIru3NkJZxiNKJ+yCQ7Lif
mNCOkmOF/fMTukiGAVmmq9vn4Q87RwzhZDNIh5iXEPiA+IHVs8Zqx3rhsmW71BAK
QRCUldOJTSdttxihIy7KI1G0lZPmx8Jc9pq+3sijpTSQPx+NpNmpV8ursKtbuJjF
848Zn1OCMkCF2604m46Z5yvuyh/Do0ZpuEPtrAVqjq/ZCZ0UWE6IQe0IXBstHS8c
fQbqKQ1fbOmjs9mriSTku/4BmvV/Evtt9TFggKcf996FEXjUWKmY8OPdN4ShMmKO
PtOaaH2vOZGAJKP7QekDz2AZbt7gFAuxCykqNp1+jiWPOuif8RUkFTANRTYJ5eZL
vEZeH2c8vY97v7pJiRheJFzpT/68+ZKBXJk1Xx8HDszY/jMnwmjWdcTD5IGf4vwK
VszHIYQM/iq7HMYY8IikUBEWfcrQOpNbZYVxeZWGrQRe/h8a1bBwzIid9X35rWFD
UJkRsTg68Cr99ws8l3EyE8P2P4Y68sYCceVNxMiaERsRcR+E9yM9KYyv+1A95ozq
yhKc3dxD60EF1fa7A8ORQf2r4bG1S0WNppVT1Pk8BsZ4lRKlvafpCiA/WYDIdtCe
/XczLETjErQjenxEdmC4x6S1vzgW2PM/2AcZr8fn9WgZuVYB9Hc+/ENUIcIFjcVc
pzD6Z0DHDIGrILrmPrQPAnnL8dCCmk+t8k5FWFOcZa2iCrLen1uV6lV/f8tvz3tC
DM0soKMebxo6B/GZcxyLhaoWcff/37nGx5mjdLSohe935ZiVplnGR3akF1lvZpkm
hh5mEIiEov8em5V9SNfLi/n1WiJ8wXwxQeK2G80bZhb6mVDpJoEq2YSbkfWGv6Ow
xnJERAMrU7e7Km8PdFTjO8qNP8TO4Il6kOJUAZta7QM51MuBvhF7uTSqnAI3KiBt
j7U3Jjzed09J5QgbFSwbAwa72afT53tiKvpnSHjx9uy507GeDWshP0uOxl/LAT6P
Hc//7dEb2rDzV17/73d//5T3PlbcTlt4Drz19w7ahDrevXOYydVqBSswSsF5zW8o
xifMAtqMUuQPgzuj7iLrPihh/cr1eOXItupt6c5+Le9Rp9DLSKwA58AHfVNTj9fd
8NhZpztuh//nOi1LKuct4fRMqhTdWUA2PNlIP6fOSuqf2Dgj9AtkD0T3O6Gfs33n
6k4K60KDOxRkUDqQBDETgUAaalvfGuDA5eeU4gsF6og3ECFjbIaAUz0O6BDEsy8l
v+1pb3Yhblnx1mmxALsFODDcC3CTxtgTXJ16j2wU3gilHifsP3J/J+4WAIF5pz4w
FMwiwWrKCpoijOKZonG5Dfrd995JT2L45MKcSRWJwaR0+1ANZYoHtgv5tQKUI3zt
+VLhrc5U4wQKvCWts5BKr4HZs3UWAEKORAvcK6C7JVERJDCmgBQgJQMPemIG44rX
q1VrvwiTDZ1XSrntKar60X5NKAUwV0y6WMT3dpy0SFpr7afEyTVdptoUR3cm9K6J
B8MszwFsXcxY6Zx2s/M6RZrNjfeE0BTNVbVvsLEfG+FYnj7BsakiAh/GCVGjV0Ke
LqqPItoZTiVl860H6our/8zXjkCG6C3tQ752eOgHt0RHiABU2KRP0ynPdmyRiB8X
bB2mfAzvnuf2zMxLMwT0piddGnTDEkdxgOqubrB/dwpaBMMc7zsHyWx8oNnZOvwS
URhIzsVWR27o7uwqYhEoFq5x/WWbvtROemqS61AVzCauuts4mAPq8l1xAZNk30KD
en/+btS6YLMO3EI1ITD/h+sBjTafSDI2Pp+eRwezZ8coCLlE9OfNQ4rh1oxrY9wK
gkqATYFvVb+2jzahuYTjVYZVNW3SXdXfI0h2cjexxuJH1S3ZrBaiUtn4mPbTLX04
acCw8h4a1/bHerdWHfrSq3cyJhHPKc+GGBT8C+fhQW2/NR1UtNL0ZePjqee1moKq
qxzhxEgxdrUg0oU574EgrkK3Mj72+g3un7QBsf58IqnafG/DTAkJk4TYVcxBykLw
Ml0+bK545WbZpGxgNtAAidyUaG8JISiYo7pZI04AmUrVS5phUnbPMMkqBGGKEwiP
ua5WX0nSqWTCbi4TUNpwkLe/EuuSwO4XSukh6/yza3pEWlAN88GABiIVimNzjdbt
bPTzQ4Ict00ElEo2brjvCgzIHLOItH4E3lEwR+XDtnx/1hP1E0K/8KasQuy5aXx3
0bfyXvgtKy+sRIG3t8/aPSXh/zDcL+Pz2ldwkayuFcU518HJJkrKDH25q0R/Zu9Q
vlO2GYcAiVrxow2EcxhYv7nAn+uLuJ5fnsbOia8aMfRlmlzAUdN4d2hvf+X9Zrc5
ofnkbNPXcpRWv1hMDYsOhDXS0YL94qYw5TlX0kv73wN9mdx35W0oPtMM8MpecHQR
C0AKBxwhP7SKqwJAdfX/Y1QzPxlwYNJfPyzVeKHS/i0MjtgphQAD7M9VrO2ZNVdj
UTu5pHguz1odrfH5711L/CHv6ILfU/fkRLOrkgFj4ROgdOkELi04OhDVUVna7bwF
uNrmYhMYSMAw9ZHov5lHXuNWhuxBGowe7Xd9HHDc2wq4xmFiw9FMBpN5HWuDSv9m
yC/HK6PqJqck5Wi2mfyHDwLgePWKqqOBrKO/IoYkcKjiIg4YB9EWO3BIwzg0JACl
MCQrBYleooJLCUCx/vjNxLwW6RnEuFvWnuJEVmdKRDE5ilDOpApK2zTvBiY0erx7
fV+kRpPU3txPAtX7NhTWgNfYkAqN51XM7dXc55xZGJYtAsa9HB7UaTw3FkwbbS5N
S/aYVuXAZT7sIIGqWvKZ4hNwKtJlXkAXpOm2/fcBBEGaTDYFHFuMrl61nBnn5Fo0
aBhwbweY+A2UO1ZcI/pjwc+K7QQzfZLgyFMCnnWaGLCSzonW5cwldIOQmf/uM8oI
1MXNdgyD/nMBcmOz1XESmdvzOCZ+griGYj84pierBMH9Hoh/uKGsyy4ThUtQoMkO
4/NJfpBhaBNXUkZ4MZQIUQqJkbjBWQxP9hxDa8QPyznNDpITyRfOOfcjdHh417Tj
9YyAo0InpROmcDZu3YYYL0rLToPKzt1vrRIAGfGLLBtxuwVKRDGSq19lvKbDHwK4
1q8wvYKJwc3O08JnNIEuT5JVjgzQqQdGLsc95soMT8JKGwn6yO720idpeZpCSkyS
tm2bIpQFYgHPWGEGYnPqQTaB+/Pitj5GUSFYDrlyKwwqEPHfksqVebb+RklWNm18
oqEBiiTpkvSLGrqTUx+IRoSLIVLxOlvwpPwnmqkL+lU64O8NlNgkLO34My7zV+VZ
sHTXyREd88vjKhQKiWtEHe6gqC5D5tuZdA91DDW2kSCWPN1yQlI4gPCggNQNPenx
WABEK3OlpG9kuG0RoA47lq4q8N1nuB+U5KSP/GrUQah2owJAIAMVBcQlsHtl+FZ1
8dut4I1wbkuyMRlmbnm0wu3zmKg25dqewos1XB5t4drvjdA1Uo5uSGvxeDExeY5q
BZeODSBETrllKMf5Ru6iPfLKJDIpeaf8tyD4ypGRJiJbidcBIFoR/mvvz2GLi7wl
fdkANj2kewPE8a0LwWyWa1kUiIZDhbn8goCcz4CMA+kmXNZlfXZ4gvAoPKKCfBRE
/ZroZ8/i5nWgsLZ6wL42fquNNVZDBxPHexnUFeu9C0zvlfIJkOu3RSJDViU9TD9K
2zInx9HRMFHf+2tVOfUjydDsRdJFq/ESt3ur6lGt+8MDWaX9VOC3gf0tBNZzUV2S
RYY2TGs3NM/+3mzlMVREomrILGzjZ/H5CiZBTmgKx3mRAdz2ZbgWX8ZxcMGJyr9D
EfnJJTGiBoN3Sjwt3aGs7BVbTqNR68KgknZcsjrjFlIS0PXeBiU+sKJT/EMnxz0/
AW2BP6kBVV0FmWjPUsI2Pm/T11RxFmkktmRcCiX9WAhGuq4hT+uNpbkT79jdA5v4
sIRsF5WT4yF9VViQ9YzmRMEFIXTsBMyY9CobqF+WSlx5lI4dfkYNmF4iSnn9KQGu
MuYxtgoZXJL69BHe1oWlS6E0Avi1JpTXi+VuvendLla2xP46HGvupGZddJyn26yI
B4bAanrPLTkMcfmNK0l7SJl/tXYW7kgre+/ClY9eLYPhp4H9myVXt5RaLozvV03+
3PYEATwV/DWCNfJ3rBnXzEAfq++288OeIIq9ksDQkVjAUlrCDWAUjH+7+mGUjUGy
7GdrDUC9+KXTom6noK0jLw4VOTmGepZJQimk0IT9DITGRJ6PBCbjJViRWd8yo9t/
AK2EVJqHkaM+y9Kx4/U5hvfj0jbXUbILS33d4DpKiWYrmLe5R/AX7v8z4WbV+dhB
rt2mHvgW8sbatwQm54udPwntNn6eZXNCM/nBd/3whB/kVnxM4KTke43yodIGV92B
qvddkx7V+XBqgz3LS7FqK0vXY+Yx9MnsqnFcAJbgjRoXry8h+JskQmgo8kGapx23
SBdT0qwg8kcCHXSHgUnfJ5JSeThvdNybROcAEHCwAZGc/3yjn/kc8s7fsJlcyhVl
zLYLOcjKpaPH6Z4eeNjsnn+Ck0DAFNe6guOd4emh3lQTXlBG9BffyiM1odkk2gtT
U6nM3RqozXUYCPUS0ZnU9NzD/ewQVUcwo3zUiH07vgGOhh8VoBmLn8afSzmqdfDR
VLZ9w7G6AIazK3MWR0HQRYXHw8RkcBQhaA6otrPjBIvx2iqPl9n+VX5IMeDHH9A5
gtDJGzXdJmtL7NbFeF8pPvn7VYVxWvnnaDjVc+U1DcX7ROulQPnMUR0EOEcQ6K2h
iKa76IzUA/3IR7Y3KR7Kq4+fKaSUbwsQTnYKqduJfBlISPfyHykuL9vZKuhF9R4E
YsObJXerykq79IHF1zHRu3OL1TXq0BO2VeGdQQknhnPaYyiZWQYnkY9BOIj6gvHS
lS4QZRoVeeYWJJrEaGEn+QzZa2nMUQCkVk3vnpVU3ZY9PXWdIX4BnjnSTIDt4f6k
qOtnoLLFzNKKU43WPW+kXQOdgJ/b0cYP1abYO+bFC/Tp/0HdoYL040gmOnsZjk2h
9Z/cc+/Rh+M8kTAmdAzWP7vBhX8w07Xc0AgcXt0vuhJm9mylgPLMCKH6U6Tl5qAL
VuuDGTEMY0/kmLSPVVfXs7KzFBJzcLdZTZ8mRoWXcmKVfZROJfaCOfQxMOM5o6tA
0BMfixzxmgQOZJB/XjbrDll2N3Fy8Dyqg9dwPGYcDHLEWmyUYcHAyXt8uvsBG/+S
jLq37XY+rSBd5MjZa4frc/TFW4iU+j3kOyqYEmSJq8j1xCrwxWXjfPWC5/j90zpK
JkeGke2C7uLgXiK9DGA5ImjelqS7RJS2xLfywsASc4Va/Y6BaD9KboUGAweBvun9
yx5C5fJz1XDBFSUXN2Jjz6ymDw02hcJyFjP5xaDRwl/fz4o7hCgFylPD+fzzBe0C
uvm5rOFwzFuTW6AlyM2Uml69hMlHWLYbmRbz9CBOub9IX7UWCEkjcYKRNxDfMajU
n2dZ0DFukYK+/17fMZbWpwj4O3/N2XxjG6HlkAe9DNGk/bbQB63XWJS5Gi8wfamN
gZmPNTgirTQ0KkVNLO8jfZbAb/vzEhSJkprZ8SQaARVgWRwIydN27ipoMWQKDW3r
5h6M7QXGjHkYcXZ/Vld1dJTeKS/NtLYMGYjAWiB+yVe2VA79Vzdv2zARwsDFL5tP
rFpaoHN9ObGsuAv5YD4arEh/YB7HVGUAif0MVPrCPOeHMs5JL0/7H3Rq9MmBD1+B
qydnpb2kTD0ZZQMDV+7hJJtdZkY0Wo8i4rtsuAKKMPxQX6TeqgiTkQjxq752VQbp
20i9a5IgKw6tzaVqTWZBqjvNSK6JtuiTQuiwsPTM4CZEz24mLrhK3/64dJ4wlkyT
Vh2c2BENK+SudCErdu4o7CqJEnJ/l6sAyfvDUlkN/TFM8nnvkRode75SPXFztlGs
vinqv3s2RhyB+6AR/boCDVwzu7t2JwRlUB0VuhiyoyEP7Q2Rrvhks21HnH9LqTd2
mg5DOqgcZN5s7xgGcg9fey1apiqcbp22NEUUmR7Q+sXjpo8xMMeQ5B9II1WIUX5k
QI/mRXdzx2EwEK21dIzESOTB7dzy4f4+Pl2/ea8csY/bumOz0cVaYfqt0OOLoUMg
c+qPhgMIX/bTRau8DejBtPhw41vp11z1OtW1btDT58UVWcX832Unt/OZvCP86Mlk
amKjnwrBpFx2cpO8cO9jCOlblKT9ZbPsCaynvsGPCbepcZQ+hlQgtCmrdCjLeIxG
MAgFcYIQgwg8EYzN16ojbcrganJjpWrjRvZ3OSSS20O0pQbdY8hw1nHyeFvq/6YL
lwpT7/njLUL87KfSFQgX9JWn80DJQeOR4NxSC9PDMkF/GOABon/cadGBgRas3PUg
EtphGyLyyP8ae3pqAoGLdOndLcJAyVMOyGXneYZ89zR38LhlkxFQjuMwFOMGJgTF
Qt478nBLo7R7sL68jwPUTK57Yhe4js/+5TwzJXb5CzQ9svkVnrOmF8ZyyIXNHmJ7
Nes/VDPOdmscSQSxy7tyibcGBZryr+HiXgCqOTPePUDB6tzHL3Xc4s0Yhr3JKZv9
Uj+Hf++tqY52T9wUwOYRoFN3wONbJLInjrzFMy9A3DupWfmuLp1xG0eQUPV8PCBY
qh6f0io9rPF3+q6ui4Tylja40yzzMnm0S1Uhz9wJMpViV8h/knkg6keDjt/LnNs/
RpQRAVCGUrzFvV0uNVfIxoITn4sYVeFN/lxBIATzcxncIAqksWAgCdLmykEclqM4
R+EGRX8ZCZjnd+q0bRgvqIL24PwgJlfTM305zZqSxNuG7XvvcmFDkaSS1kU9lfYb
rHV6GATZU4RSKhSXRGLmlOTnoU8X2o5rXU4vg+QE/RYGVO9JygEaTTBx17MOmb87
rinqerR6y+8bD4S0uRDkA4z40x10TWEQpeEPDH0H9OPVLrUcSFTKEKyO4vUr8Ha0
HHgodZa4M2cCkJv9MCb0TPO8FC8P5mu/8mGyhZi/rL1jybSIMv1bks7xZud7te/G
Kmbz3yLpFiaqGuNPdoEtEn4kw5JdvNaIi6bYRP79lMG/n2xoSzvJC0ZeJ5BkwwCW
X2QWw2isOzRQad8UqOLznjtmqHrs0u3131tAFOOd0qdIJeEQcqPQKVsm1LoNb5sg
BaVZtA3tgG2FKNrWy/kX0I9N92TSxd1RGhjIOgyH0qqMYQbv0brylMy7O43iIe2c
N7Nhj/+ycHV2J2qNPwszucNH94/PYbfFFgH1tZVGZLnuAJJYt9iIekWXXD6CHyGg
hlaJbWb6mrXtbkRhD2fKJTadWZ/7fh6FkIJjH3eC5dPf1lFiZiER8WszTF+jwpQ6
dVlNIL+9SgRP/aVkbwwHH/4m5XBufV0A3dUtiI2SaukN64tQX/vF2RMmrdIQrLr4
6/2gxKTvLpf9cH2zDfRnPkjjVc/m5Uwasyvi9t4xffj3b2m8yFkoqUIluc4hJvmS
WhBRKLZvLmuOKPOzHQRYkCKuwuTm81VpVmAj9SlbsCPTvaHtVnMnOzO4DeymIKRT
Cg7qx/SjSUqRpbit+60GRDpHKBr+SmsIqP351xrm4kU55dVB7D2WVIufSXKEhrUo
nSaIERr77ynWWsd7O3JqzljFTL6WfB7TlzhbQ+bRiimu9dZv5toWwA+sgLeGCNin
Cb/5ER2fopl+0s/t3nxSFjB+YJFm4JO7Ptts/sC/ToC/E2+UrEzU13a6j+XCX5ha
h5CmYixkTCNSeZNzRdxvyivbZWMREar8i3BpMmxXuLX+CG5o8+k9N0QtP9ZS0aR8
gQWpn4UjrjmUR/qpi46IHYTTXCw4Fji4+QNgT2L4QRrbUgYyiP5Dpe0ZjDRC00lK
3+nfe7u5RvM2Mi8hRF9aiLN1QlXj0WxqwyzqKxXHbkKPZG9Xesc31JlLlcVRXK6a
YpvmQSkX6mMcD3JJGVMBpMPp3OU+C4LDH6Owv0Emy2US3RlPtf24C2Q5t06MDrZo
2toJoxn0KN7mQiWrrJOVOAoI7svjvaIik0L7ao5Ppx4IrgikKOQ2fDq4YX28yR8P
DL+5MT1IZK28+UKw6Tt2qj96yl1Kl3oR6VSe92M4any5reWTdIv8yD7g5ZbtbPip
lFsrJHmzs2xTFGEam1ktpwbRxuQYbuzljJ76+uPP9jjP0N+a6EeKlt78mkoGHajs
UV1bMSetdoEeXAtRE3C9yyRRogcVKyOjwirtJbCYFUP2J0OC+8bnNuJriHan7z0X
53bWc7Z1crG+9/3W9oPL3N4nikwIivMk4jLUWN/yN7timT9BPEA90DN6kH6Q3KBY
VIkZRNm7QfLzpmJIV6Zg4lzBjcekGfYuB0nl963mhYvwrXCtGhNmNlZMoGoKvwj1
4ucoY82fjtUhDkdoz7482+D+RsKVQFIdn+wbzhgZxF/tYrMxC/emLYutbQ3Uzt4z
w96qidBP9adT6jgq/RmfH5CFIKuZcNng//ZmqHRuC4J88C4C5CrgTBGE889T1pE/
FyzRYrohVJKfk+lGfEm9e7crp/rGMrQU/R983pKHaYNoTZKh9G1cZyr4LX3wG7AQ
k3222WzrM8aenN70+r8mzvV/dqSEd4gU1IrcSiaRyq+DRWtBr03Pbptruhqmgvdd
YS2B5v5uCehj8uwRK6LC8YJmJqcO0IAFX332U0u3cLiVrD1CiX739c7S5/z5MEn2
DBhCuTfBrQORLeUk58ul6SKioZxhWqIcD1wOgbD/8FyPbQtTtEHLeo1KR6p9Zui5
IU19vOGAwAx1U9rg/Z2PMImBYvMOqlDvd/fWhaAHgO0D/o+0TWFPrD6FWl16Gqq0
ngG0m6XVV6lPAabMns52wQd71MTeuIgGqUECy/EICy86CFLHnd9At/uxd628J9lv
jxvtfTYIuqVPhBgeAb5rp0At8QvznvHTQfb0ONIOae4kql3bfR7UB1W3WsWfRhaK
LNndus4/vv0WvTawu/0+YjVHUnhxHkx89kL1lV29jP7qk8O2BuP4vUrY47l6lO3L
gXmmOO8S5QNuXwdaGipJ9PMOvIvERa4FztHQ3G2eHRyYumA4alGd3YC3/wL7j2iw
5aGGug3Az9Xoo71duBMtLYcsHxq019QMieDEXQ4qXvg5hYHMxyrYloeM1DjEcvWT
UB4aZRjchBYXER5A6/IPzZxCZmAqDGnV/9dRlJywRaG+a13b//O9cw9+ZNEVVDxD
MP27gy1heRDIVnjzEwzfQEkyvApVlWb911DLdjseLBw+gvq8Vi3TSonj7M9yfmak
61Hj4I/VxpBY8on+0BTNWIIYe+bUi9CVajv7Refx6LXg4MjwHNcPzTUL0jZD0wu+
bNEU8iScY0HcekK2esOlv32/dk1Ey/93U7i59A1a6zWtqSHWeupLOVnMptxEN7/S
duD0jSjLhgjd0ko9i6UTFPPQj5UjTzOEHCe383MfBU7R10zcHLiE96cHNeY7T0hx
DiVnNCwcX0+4iBcvQloX+BygdxbD4HhI0pSvbxKLzvbh+i047KyiWaZzpjB2/e9H
w/zDzHQ2Jf6rFYSJ8tQnlhSmqxkqrniPJBudmQ5ssQ6vumViC3WiLm8lManjnUkr
rh1TcJlLdTfRYtXCCTeDeltuhMTKzG0kkdr1Ug7f+IdgJCtKvEvmP0YcsDuaGC17
OxXl56DltVd1XBlnrdedSRPMdG4KjCWyHXoQEusPNjypMcfRDqcbVHxAx2PXOZhi
UaltMFL5XWkoPjfJnaRt6KFnTlC7+vmaX4Q8dbKLmd86sUf2KIdLBJcneusNGTgI
+/njaXejhzu0yZF7ETPcP6gXiH0vidDGuzqN1ussJS2dx8PhGnwZegIqmUZoQK+L
M+2wkOUJqbqyNmFOQL9hseZHFdTW5ODE9/TaiOogi4nT/oTzhRtYplHhVWPUvMzA
vmB/Nt+U8Zg3eVzhKpwUig04HorxhHvljPfWJzhLZgbSlVPBUMwqMQIO0HAjTqRb
rAEi+uffyf2kGpfhkZlcWo7stREti6ePv2RxX3EPxEnFS7DUk1pM21vZloEehy/A
VUajC03iHm1ejbGJcB7AyU7BtQFyDHRrXjJYxiZRnuj+T08kHaQkZENn6KlQRxgC
hpAxmYvspIojPnDs2nAe7sFO2xAZDYsclJC3DLqnkk1PQQFsnkx4+y4XlJbfQsKh
pQzbBPGuDqVy7IBLcMZm4oRyAz+gY1CLPDlVXdx8Xbfj0DIZ8HldXDZ2GMzWC1Un
zkiIBwJsyD8sHJ4C8m8CS4snXNNGmxn2rKkKWaTSt9Daymdq1uzqVmk0xLlWIIjc
8wEq/QOg7W8Zmn/thj6dF4Vf5lzD3N4cO7x3kNqceQ9jDiE0BiHWseXENiA+NCpF
KQBbnO0FX3Qy0XBlBjgw8Hmgggys8YpY3enfJZtpkIJDfyZTyWsRnOemoCsEfGtr
X3IOtYOhwLAPU/RsyNsgqsr40VhBZS35176WrIIyL9HTMLzFDs8lejzS1D/wvUF0
6tRAudsuXcHh1X6TTSV0NbaW0XUPXg8dSBKgoW7FELvkN2jfqNreH9kNZ/Y+ugPe
LaYx2kZNdC7gzHDakwKxS4FA01gXZYRYx+gkBYA10mGmcBj3eMFd58FZZ1/2z+jN
ESqqVNK91FAJInZGgyLqujBE37y8NuH0r1sO8rCMUWFY7ygYD3MXLRXB87JZoV1j
GKBKvUf3yedAPFl28QvrsyD9AjYxpDBAN6JZNUoEs/n+OSaS3weQz/PGV50hXbl+
Wbnz+ERmCj9OilklHlGjoSyLYro1U14KFKB/CpSRm34KAHxa9GHAjqm9LowwT7+B
5ji0el2chBlJyDHicVFFZLWQQUE56L6sxc7jN0C9mPAcl5r58LVcBWNsqmWBEl1P
7ta2Ytgxuu7BYVG/G581he3QnLKnoaTCKCiE0bqWQdN1Roigc8vNUO0iqE6UWKkZ
Hxc/nCa56vCMK4lLcmiM9aLSJ3hX8LVqZIGVrh+sGzNgl0dBvoXuUGuHfwuFuxs1
+/UV8R0S/ZIa77Ut1g3XtPUJ5aGuM6BuPWOcoG5Jcp0K+AI7ugoLLLnmkuIWL20b
4SOY72fRzRDUYkXNOwDIqhwDjuOE9kpSrbxqWe9LZ55g2EOxkloGapCHIMyC85vl
HObkLRonKh4K/1x5UHV6Fa/1HCJ0yHf6K7J4i4qPA9vDhLXz7CbzZ05l8fS2jHaS
hVYqXDdiyax1Yr2xbnvhqnjw11Bvq2gl6vJryE8+1kI7liEVcOQkhwvAzgB2qQnc
LBPJynAmD3tQ/n7Z7saS2qTj+UMxVapjltD0yjKl4CKpAr98AELUnvT8bmJ5xv88
vX4fbpjL5OGLsTNk5SfaQB6XAfffQv0u0bE+lKtyL8JSM+mAvrECqUP+0Klu5acO
ioEvh49N9SqXk7Ltxegg9jxLSDDCUvZg4FxZtfB1yHto4QZ5AwfqT4EMujN2YcWM
WO/Uxv+ApmVI3QKu/vdvaVWZFLdXB8FiTh8nUsyxPPreS4UmOkIArgBpJ9bjqaJs
G4t9hriLMd13SZt3fsRRsB0H4RGIM11ehnWEYEYz8HkuMqtPq0bPcQRi/LxaOwOM
yABDgAwYJjTTPHSSTHPZYp9gQcR8pvBf42W8nCmOk5+6B8zXaBQQ3pTAUii38qYk
vHgTnmFcT3XirZsn9QgHnQHDYeZQ/DzaT9Tzzb+pwZzwuCMuJSaE2gASQR65U2Mu
+OocPviL1VChS/z4bZ/rXKFr/ok6ZHrqXkybNO4T6sHqBUT/qOicg+hzxm1AQapb
mUP7VVXgMNgvPv+jxXbo0WZtsR8AMknQEaBCq2KQ5bKLNhECLN1Tnm8/H+xz1xoN
FBIBJzeco0ILnmdUrqf5Yu/j0t96Hq+NvDijpS6PDnTyes6DC2C4piVdaemMUzWl
4XZPchWkkhkcajINY8GYA/SXxw7AAt5QsYPxBcWDksnzMt1/54vzyiWQdypIj4rE
gDE3/ceCIKpZwNlxoXLyDMlJGpTUUdsOmYhtr/uuL608uP2Y/H9pl350EpZMYd04
KR6lIGRLcecCImpfKq38jBOyC7Xyo5SSEZuBcmF6b3oYfhC+8PP6ovdBkLJAhgAn
qf5TY6GP8geLKXiX+c63/kFldDNdvgqAWHWJCy9xcpi1pmNukZIqvQqE49naVP4U
4SM9pQHAh6OWtjWQ4d7f4Wg1mBAbgTdROlbu4S6n1oVzLsfC8hs1M7lL2IZYRNX/
f5Gbw7yhAnkVPq4DOvMV7nzagLxsajmGMdmiBYoCTkCIfCaOd5ooa8oJ15XjPxmM
P/32o7sHxbadPYx6e7gLZTvCNFJUTBhYCbyRhzDlHRPJAX1fdItb8PDAGtI7rzST
a8PspIucRSCvVIRPPkl+/VmPBXNiRte5J7ZcgEVUzyMRdR6SJL3uzWzStoXXUnmo
aHjA85jkv/KPn3icU9NuQxpZ4peg60o4cHEmr/DSe2bf8d3pBkyy/QwO7x2/muMO
dq+7Ct0qh1R5oC8mAcsd5iKKSN5WndYjcqEEl14+uDJewmGGYO/0SkA0b/Si8QcU
JEHX2sOTN2HZ0mYUWAFtOr0zcu1phVt72wNj+/lVcjiSffXoY8SuGT7brw1pNaXq
tXqnq0h9DG6UnJB//F5Na9Is5zjZ3yNhQTpC6IZoAQU4w9WwQnKgl7tuAWfv1ntt
nB5UlHqJHdygKgMQ42SGuLVNWsmn1Zz2mmHZpjTY8VP9yRpEV2PPXerpECHDEtKZ
ZLyPjJy0g5dSSrRyJgeVfg+Zmu0ibIE0GsWr/P/v42xZhrsD6FkArO3IqH1Yfv64
LGCjvK+wqVkUI4Dcp90TEKE4erRkErj2OtnNITrHFrL/pmKwPNWo3YM/7BbJ2Q5E
enExU3yqdhTu4DwjYzmmJ1EMTDXoTXQCYWfWtnjk93SF52b23mEdnYeGMJkeKulU
3Bh/ePtm83AL0EErDHnwsdTz9UWvXp08/T08u9jcKprpup/nqB0dcBMjLHRje909
QeWIYQM6s2R5Gppyt449R2dZymaRlo+cf2mUgA0hXh9xNtquQGvZaCrG4EXU6BGL
a5Tw4/pi3WWhcqby3KpwxfnMy7sKZUmzLwtH+qZHa9CcpfRCjOUK+MtgkJBcf5P1
n3yAMYgONj19CrN5bFaIRXei2o3BwxKIyNQbDAHfUJg8zjBAMTCCUqDd2d7p1oQS
zot32fRSywp/9ZcT2wWHb/2t8ox1YvoKkWptddBdtF9zdjBCrhTdsWNhdV36ec4A
f20MwlQLSpYoYFUPROc3XqEr0yv9LKG0qH2farf7Gam92Qo13UrXHHZjPP5Jm2GN
yPBl+yvbdigTubXU88XZYDjwQYkTWgafgNSVFEf6yyzXEDvuuknNIpzFtjuqpEq2
xqssu1ggpUvbfyB6PV1Hnbu9sIXOyaCa3IK6D0t8HfAft111UvdJWlH9jj9ow+vj
F80G3eiQGZ7niYknqF63cERaHTKkYEWFuHgJ36R0tKi69kkHumPhX9HS9YoJO7n3
xXP2VeVtG1f6RMaF2cmBPS/EWBAIBUyzpvgQXOOMfFOxGeRRZKA/5zNkNmg1jxIk
05HgVlNKU4gVQEjbrB69vz7ftZoioN5Ut55VCodqEBY1fgqsFWQQSphrw1zsEhFY
AWMaGC5d88oseOhCWCUEYrG/j8JVMRMqkV8NzsLRIwg5qZ/VomRwPkubn1BEv0b1
vfw7jYs8mqj1tTEmmjT03qvetwHxFPAqlD7m/8NnC75uFyRlgn9AB19v8wVn5oj3
ZV4MRvft/zgyffzY+I96xQaP3GIq5IxE3H/Uvs1j4lWIhCVDEgUdMVpW6eFFy9x9
SkP/1q5TAuyHEdVmLaU4XNZSirt1LKCnX6YdNGZzDXQuf/cyBJT+0ZOldWWdyjb1
X8GnIiwB+G98K2/sCNfgjZCC91YR3d1n4YKzG0wvFcB8c8nWOc4jBkdE032iJn7o
0qetADIyFWVJtojAoa2TaHQja/2K/GhxmheK0QI+X30sW+YF81FPtLVlf4j73l+u
oSKHovfKRB7gusXHFAcR1duWN4uMnyQTAcdtrOGiPNoiiXJJOjwVZ1zLwhT0tPXK
8IWj82OHctSIEuWfa/soue6FrmKKF3yMSKcOsQ8ezaO9/ef+OmR9/rASGW9G2N3H
DSJ0lGbLd2PzG4afw99t33lxP+eAQdhJ0qapI7rcwbzu0TGGOKGdIMMc4r1gVbdp
WEU7FJpdC26O9gjBDzuaxzZf0vFJM/2gshgROu+qvyrX5PZLxfScTvxU/xqmk5OL
VQAyKJ7y4fn/f565uCtztyZ2EgYBmTCXT85XdOzvAUtP5bptvBaQ7wIjIhXpnkah
ike+CyJ5zEx7EUag+U5i03eNn6sxt3wmntntP6otLFpRP7GmICVhFQDGB3smKXOS
9ayjHzbvNI5Ju+1vRQBokbe1kCEH217p87maGrnnNE31WkUuCElRe13485u+A6oL
NrUTIdHbQOkkJ8JAcgRfkryKeZscCCDx/GsNYcshs7cSTJs026sYr/2mvNOQFJbh
pqoMBvcp5Q4uEPr0IT7k+o/osG2IyVz9vfbVkSApWUL2HEnDWxfdDnjZRDh+nEMa
EwssE5v36PNmkJ6plauiKxiLawlCndGh91864o3Je5sDx1vyaY1YGeRtpPWnk5CC
OHOt4Iz7/8j1B4K0TzjsjC5QM3cmSl5Rkw7iPJ2jnG4YmqxPW5bpS8eVm3n8Uno1
VKW5t2/s1dr7/LcRUHS9cm1AoSqWv0TMOvbnJvPY96c2FUyJyuYukFqLA2U/WJap
tSwNgLUmtrS4NiOAL65SDFF4BbsemvHHaWMMplUPHF1fzbqhLQehlJ5wvy3wEGbT
94eappYDVzgfDzC+EQ5/evEWRGIcsu9WSJwtEWkj7BIKCb9djSPpTbBy2cwHzygU
Rct9JbkvD22s1/YrgiPDCwrzPLmQ+PasX2M7nU7brUeFJfJKxBxLlN+gxo31+p0f
JOBUMHl4iDxTpuOkIHVU7GYtxur8zhJqZSh4+zNCB0O+Gdh2/DNCvMvY8zsvJ4yX
672W8LuS6z9usRDil7MkEh1vktS9SYlY8zz/Sa5cNtt3JLMhLheV49qzCLtAqfUK
xGW3M7BfFV2Kur3gjg7EdWnUW4n5EyswbvLY0QIqu+VayHqeAbnDD+EqjvN3hikS
M69HNDDBcVpSwHM2HVQ7/z8IdYnetpkvoVM5KB8hiR2D2DVmX8u41WjNgugjNuzO
Q+VDWljU5xi7fJcBVKVxeR/dsz1nwqL3VSgiSHMN0hK9d4jMUZ74PtuVt73TGCrq
NorMTvtPjqamUBO1UUqoj3sPP2Iyr7DOtmV0rkjmSATFdw3sp8WLNfzWKEybmugY
bEpAiKBtOozh0/kOZkPVYBrgkiRv8dSZ8ObUIR6G4AwCbOM/xHxe0n9pvxDnO9hv
TS9C0WUg3xDLexR70VW3NBjs8fju9ojrmqxPa2TcGA6A/EMVDQmfZ9cUs+TizssZ
41rxDzQ0vcrGRUMrUzievIXyDCZHEGD2LYhqoKrvCzD569jskU+z1ZvG0Q46wiGc
iJMydkQNOSmZBsvJG7snTME8DdSPVRJl58HYXm+ZmkUG/7CK7Pom8s7SaCL+sNZc
FJexzOy6fp5JgWP0xJcRSDDm3b6nrCXk+gOwmjaHaw22zeDoD9wXmeWCooDg+cXr
QMv2nLe4l3Kp920oB4RU2inx6BZJuUlG0iS8rweRFVt1LUf4uupqbckfkLe3irlf
dQTuLlE2NxsIfAdqVt23ESx3YYlARo32EZxqqh4nNwdexc878+8AmC/fCVyGoFjh
MLVULLEKlmx+unV31coW0Ge9g0sYMJpeyr8kx+haYo+9bKUIUhht25BrC9GXIIKG
aN8jEdYV5PIVUJXYkfGXwnIGmMs54HW5cwT5q61pmiqmPVNknDHj0YlXUMeYz3ca
OFEqPDJXq9t0QBM7cETdlW5E7mVsNKlHjWgp5Eub/al813EBtkLz2n8UtUPEGJFE
wRnBDQ2L7BkDF0Ak5NKlDZRlaqyPDsypdFhsXzV1QPtGMWMvZ5pKU7rHrdS0VLfW
1O9Mj46jwlcoClZ4RAPEUhCf/wCzQwjDBoOG+nZg9+Epfls6CJcN6M1hWp1sGflY
V7vzEQ5XSJl4aK0jt6dfCETa7gaNauuc+9JTkjrwktcjRXfIz+kZwPBh9J8+VqeE
vBPsEXiDZ0ILeeplQD7SBEqm8V2IjczQOng7JRTLeNoyYbf16xJyd9kq/mTBajgq
/XIYGXzuHQnG2e2SIQUsZPIhKOqqTFucbcd373LE/AapTaJleoRruaFcwIjXeNGb
ttgQU3bYknoIB2cjp3XRQzrRi9JcBPQsawlvEpR3NwbMym/t0USpNPPwL99aDcTy
gyU+250FfCuUv++3KvZ6b0u6Zdh4CNidrZ112bqUkqkIFbWxGzc3VvYmz/9yeySQ
ocERQfR2olQ3bWGko0XZWbbR8gI6JCtIDPJ7TwN/u05J4EaLenNDwZusl4Chub9C
9g6hqor2XQ1E96Q3Y/+RCzQW9W5H/cArx4G9FcSNLhNGnX8WJWqjmQbNjZ8RnpYF
QXVBgrE81WKQ4NWOlvmlNU2GgNPidbqC+nNLtcxlJBcys5wbacIFYmjl1briTjXL
6Rp2aP8pqCfpmGlNeyyzl3xOTQmSV0HS4+3SwBxfXYUBXIDXxY5dgIKxs/lvd4xI
DjfOFM+R/jGC6wi+HxoASMZBE5f7/74KCXIznJ0a+xMOl7+Z/waprynH4TIdWsW2
dpRfer7VpLXbAfFtY3Hd7E+higd8+zPo5AhQFtmNXEeWBjur1ggWxbf9FTEIxoES
crbHHjb4dEFnvymUKNjVzvg5odfKmJpYtD8Yhw37wLB6yOraiE9/8jLbG15U4TI0
4cnXk+NFNEW16TjEvOS6gkHcgXZWApxKk9rMzw+aiErFGVAadSjNTabRsCP64vrJ
s7cbvLsfUQiwOXgMxCvJIpMVZ4W1MA2uAK3ZeGZEZuzNcm/dAdP6OpWR4NxYqnCs
gDMf/iblRnIYM9u93XFZw22kYRWQrdA547Qbi9S1xWesDlokCEVqk2egj9XXpB3E
wiDOD2/uP8m4xCwS7Wc+eNN43ccQMDj2vS0HilDFBw/L5/NMw1zbhHi2UQrXcS7M
AXHk5jURy9VUkNWq3+HvzM07CcAZ7Wp2EZ/dorecSaOoNxuhh4cwmn+uIpHE3VqV
mZ8oYt30S53sOKNzRhaHhqedI3kMPULCDEZKe3GA2N826MAXBRLwWso1nqGDcVLa
tbaX0bR2Su3dYgugDhis/NrG9oucU8wLIRNMECs/s4qGnDNatXPwoJzXW1VryWLd
+i85LgxJ6DNpyBWnVI+JkyNB/UEFxZRDQL3A1EE8mRJbrrFm/gl937h+gCpS2OjF
S40Blgq/fpJDXktdX9pCjQYotMpwegAx6UXNhilnD59vzHUiDX2by47v/kO8/c47
VZzGFBRuiK6ZppUw4M1Nt9/9WEI1acZdJJxY4TKosvbKxtk4PSymnaqjPZYTeU+V
lrl+iuV1j4v6NENtnSDW9ARG9Ygke8VOZn+MS4026PkuPPdOKFoXQM1DfDeg2C6R
kFQ8KYsmHYM0yDcl7YR1jMvlYfEkUuXKJoFS73Y/x99ZBTCgKquvZDBFypp2IIQ3
JmVeOXsRYuJba+DeMiRhvvHyulvmHiz0+i5D9c24o412E+2+J8VAJ5B4jVEwyRM+
u3oKAWVYx2pfaFFPwKQIrYUJ2ZaEWc42gz3aaWZ+waplFDcIXk6p5IxCyAd4iKZy
fFMdrJdevE7ktzUsHXkpAqJ1FnsQ8ZRsQY1s3fubhu0A6J/w1HVYrLS8/U0j7k2x
BfYKCIF8qPZVfRSWTwN4JjSbVfUqnaxNsMXdRYZjk+80ijP/AADoFf2dg4S30Lcf
4qM8pyLThPmva3dpna9rxtjWmkqZNV+BP6+xE7zDrhF/YT2pYLi6RGBRwvgjo8Bn
MPO+dRiHbI2oR5YEYdba51zWHmMd0J923612OREk84k8Gmuj5bPC3Ddm1YSvKyv5
oj6yjoWXmrO/B+wMfYI+hzWGMvNCUSPVAlKGiN/jHXX008CwUDM+GozuB1PYgT0x
YBsqthvgbuDScMxqrY1sq2aRCMtsY2gYUdh51y08GJPsYeXB+/PhUolUzjRu8Xx7
Vz9T4XhWJK6XyGCAWG1Q/BA7/eUI2UvI7hUUGAISoTEXMWmhsGhDwTyeO8vMOarJ
YlY1liZp8pj46TU2DNdG0RWsWW5wFPUpaDpOEOLH+zwEVVbqJf/+fJKgm66WNd8H
J43gYl/AeBh7T0tkvuPm+W6gXaI30hII29+iLrXvjIlljyuhS8klrV8P5v7zj4oO
MuJ/GAJ7//57mkEY4tPCcirrq40SYNgVdu7DDPQNTv0ouVBVv9JlxWpZxGWkVXUF
9U8DwIH2vE8IjOZ24/3LxWCtSRFmUuiILkTdwdgcJXIXqv//cJqk5YFS4FaJBmzJ
tgmg3SrX2boQ1kfJCzwM7zG+p8NfycYdmqiRZFBPdKwsATldB1afvMLKN+R/9O9w
pdhX6xwbOyytqjzXTGHxdjcsP8WpqiXWp+BVDpjRYxO2a/4QqWo7qoE6KptauhLZ
4PU/qvmVWC3zCBd+DN9KtaAixnLlHKuunYIjtKZjqh0+ilIoh23Yf2w7b72ybrdv
SPOX6l/ZF1ktkc+60CVeMMLoYuMz5/b0zjewP0tEoMB1Qa/GnIhsngWoD2h/SDah
62JebI/GOn6hX/UmIDOcseM+0rM0z8HZyx+cafSTXvbxYgJouw45uYFItwROviFw
vCUuotIyBMHYZ+NR4P9KphHmPuvJQ9kU+8H5A+vc3o/k77lV8qC8Vl6voLtFTJuw
KrtVIiAKRI1ta9cZtxhef2EYe4/7GGKAI2gST9TfrGkBERlZaUqdShZ7qUIoEXli
vyPMkHpDAALiEGr3ZvJN0ojK4MTiNK/IF+Ihgv4fIvVxFxsIAbqe7Hb/gq3mw7Nq
AFiEO/BEMMWMmGZk+TH0H17z/H9ZfBCf/bZvoPtWQ6vAOouoB96TXeBOtXd5Yra2
hDnV5DGaf5tKdXb25JxdQtYb1jw0g6bEbVrKXiEDAF8+mO3z1hXVoB9u531vYS2G
mB7JYBh7iBKbbOQj4EvoWxEq2ryKi/rVJ+5FsjaD9Eode4RkaR3fNaSW6Js2m0Tm
6jYP/v+f0pT8ehzav3Gj/gMxeBnWMnlZ6SUPaDJumiSRw0NGL534E+TiL7IuddU1
21UoETz2KmRmGyrZfuxI3wZmF183NKlOFswuEqV+SDyGNqcCisoc+CSjDA/DggdF
Nsa1CBK++ZvR+xrr1HRMVAz8ZeiRf5ZLSwfVbwUdzdM5m8hPIgaIO7E/UUyoxEGK
8zUayBluUr6AcuBC2s5B+/FSy3yObd4ole0Ia4XbaYfppkKX2DTw2jPsM9G7JcXX
5d79wuDbU9nPFtVijffB/Yg849gQHFI5bBHXvxjeLYbA1yoMNFyUYSGlEH5tiWMX
a0pd7JVQMuF1a7zIJVp+tniTWOEJalpch9w9cPV6NZ0FhprtAQxtq3dw3gsSkX4H
mP3Ak4z0kx4ithj3XQO+1nt9rAT2/2WLCdY3UJwmZBpNSBOjsv42JPIsztahO4x7
gWtL1b1anAgsKwVnXr4deKXu3nMteoOqjP3Rkt9L9UTNYprkwYSWoqtdHQFrgZIH
ZvE6nKX62jygJUnxxG7hvHLDpwznAWsCqW5u8/4k/arOhJF4NUpGCgBOfU3nkIF0
gVzR3fHFDWOFM/YEjANo+tGDPkuZpJxoknaQ+ghCmite2hEWVLz5RUO7pUFMnwnb
t/3a7tA/mNK5YtR0dJq6DjN3vlJHlQYfdUNj4toBOLxkPM0JdJHWKHNfBD6oQxtt
CC09S3nnOr+s6jePgr6p6mB88hdVlV/gGIv5RcUNXY4ahcfOYnfQcu8+YRxosVPP
996nRpyh7UkysbesKxGIlboTnu9+KaGKpb+Kc8EnUKHmW2FWJFXhQTxCnIUfzATr
8ONRLpmE/2I3GwlJxm30RqaycwHpKP1jIzQf424qzNqv5Op7WStjrL/m4bsJSEaV
7fD7auC5tK1Q0rrqkJoe67CGkT2NVKHNbamfBlTRbmtfaqsFXJszbuYKnMJpNDtj
hObz6pQSvcqAtY6Sdx9AJK+mIjnYeQ/7i9bCsZxHoGm6uz/TbnyD5i+oTftJf0v2
tT2w+zOQSI8/gLi46rq9UNgwobdp5GWfuCMUqg8mgeax7TZVhbGtg5Oawhuddynm
i6EsOMn7ZVvpR3yFxJ6oWSWzKaw4b1KOHO6oJ0+zeSEWEgGaDNZ7jWH48/f1joXY
VtQtm+Y++TpScNZpkkRS+88jvKROJ6GtgOonUuLx6ht6cMLLzLLQim4eDuprgYUC
coFAiuUOV4Fvd2Pii2zZVhIgFMfyfkBtAFo1mqOqe+GUJPTJO0PsP+FXXMZXLB0M
HKz41l1J84SNNPeH5B8p5upllvPzGrynFlKgZQbgcx4Hi5AxGdWl7H3C2DHmOzLW
1RHhse/fqpFuTMJ0fqgRbVfcJz2MbYg072jQq1ijweQLZ6klj/bMeDYRoR4LHF8v
rtN7Kcdc9QdLUgSeh+1YXWZOHGg7E7z/JHDLgauhxxBNBAidls4Mie5og+odrQva
QzNdMhSxZ+6gGxFvTeqGKsnhxckDNpBBYfv119tDvZg1n88Xr5EqVzTG6FIZS466
zRKFlE3FyOG2Kkn6moCf10cWJ+7CLvbRGGO/SQjgAiaWeZ4XZ7oQQmBocf1zZpnb
0RITGNx3CWBd1IlMGUrjODjz6LtzhHIrUVW91S1+8YL/5k60Sn9171dj9cprRcED
TCPHvIlP8nnft4VAX9lFiDL+43XQitqNXWYHJgh8MBC3iHehiiFg8TPCYvmz+1h/
PXo2QGIjrrQpPNeo2rFCkSxDSURSOhXlMxqWKlQIss1rAvS68YqApQeqm6jc/phF
bjPkq0/jICFzmy2EaBHZ36TjT+tpCT5EZz/KHN1SdyKQujjjTzOPqwdEEor8h5aX
ylA7BtByTY/zCc+DEYSM96cQWUi5JQqhR2FYuukSYWizUwWDBAuh6lPG9f1Zbsq5
tNyE9DVcJs+22xoTR/a2F4RWda3sMATJokwprrIEPURZ0TyQoAgPCRCHT6RHsRLe
RuDKxqFbZpv2IHBIblGBJ3c38NxJOGiTCN5d3vnwCjxn/xnzaPilMDA8q7NrP8LH
brMQ9XdZOTvs45Zj/eqzIwEykL0P9pwYfvaOcwaym+CY5b5bMOJoeP/8I+Jm5WbI
7gZvXwB7fAkXno4VfLWvbsiPKTIi/IHSW5K30HlQl/T7nLfanel/lNgfiS3Zgk7y
h+aYRvkIosbZ0epSXDSz/kl1A0baA/QhXhTekXwqOXnfS0t/dWuU0xuWpgFtO9cs
fycv0WW97gL1N9BlcVTXxL23jr2ltUXUhn7jweWosiS294zPGRKF7EsTt2plrVME
KAqOpTGOqAk0ThdMu8aLLSTaC5UOdhzPJrJs2VCoNA6jxRRsLNoWIAXk0gyyRCW4
4nY7UF8TJP5tT2yHm68tDk2WUpsc6WhQsS1QOGmxthvnBAKhsaCDcTO9QWwdToku
+TUnS/QGSWLWEXz/bkSZkuXmVWgMT6UZzLo+GAflyG+4vFvwiKXuNbP8WF3NYdCE
zVrJs/6HLP8dG14m9uidf1cxazYhivwRt5U9vart1AVZiWIGqZGtEfo/q7m1wtMQ
V+2whEV5y+ulQobWshM52R14t70Wyqu+woKRK7t5vQRsn0lYmnJEbFzYXy/yGi/G
2PxXiT3jqHpA5ChmLaZfFfuvfr2/Eew+EAFjLey20fRE987+q9Dwz+bNl75pe1/H
vRhU7EN/0lyudPwJVgmC05l8ZzzKJYZVlFMc8kczevBEmuGsNOnR6bzOzn/A4+yu
BtRr2Lm2eSXE9jNkTb2SKOMBLqJQuXUxVLeZRvxbg7BurYSgkPGxchU1ENXFKpVb
/Fm9mxPtL61AYfJLy3KmuCOZ+6qNSw8N9PZp1QrdvzHPgvt3PNzpqmHOJhHHUXCY
X/oM7Xln05bnUlY735dX5qLp10NHnmLVb3jOXYzUXyczPF1Q9LWEme5ELMUeD8vC
WhiLeFRdAIlCk2RD1z5c1swJvxeBfHQGI7KuRTcxYoLwuDpM5rux3Ib7M1xS01fD
Y2pE2Bz2xd7W8vAnkcNQUn8rI9tjLNT7j6KQ6FA/XiEy4st4M+Tso2jc0bQgxWrx
FF9PckcJbTloKg4Ndni5vkbywGyG2bLjZF4Mu8/k9whXLFUXLeV/Zi79beh6JNO6
OgSFuFUYGeFefgQbegwWNzAsumkL74IZCA4tny73sh/dnkru6vTb+SanaqF+RR+C
zABtxZOkiXO7hCl++evaLkwAwZYgucjZ/+6Qmzzs+pjs8Hi4PzE5w1RAzmT9O9n6
33pa/m6NgOxSN8ElkUC2BQWKNQOzff3bqgD5T4nVd7QR/bvmRQ9D9bH7yb3tRiuw
I/sxgc60NNGh67pZMy0CfN44SXbFp/xHUu6MoHQRKDyD8wBOrDqc3L/SsUhTayAW
7DLKnOBpCMfTFFd27lP/ZyWLRIMpAplcX9e/euzBsDqsW/+BrEXxjAHNVeVb/PIU
W0O3wo0SAErMSJWGvJ3dqsrqURpfuzYjLo3/gwXo5XMmfl/8sFapKYlPu9aFoAHM
eZ0laFcpBLynX1eGpb0H/ZLRDR2Hgp1/5ihsM3HiQr0D2XbHeczOrYopOX+C/kbD
BtCbdFHNPtZp9hMO3MDLvBhhukC2/UuxWgz0iNbxTt7PJbRwqBA+D7ZUfFVlbSmY
CPskxOKXOL0easMB5KMqrVneLFEvgWIXvI/aBgx+ApOcKSq1vK40erE1ZQ2l8IGO
ls7qW82eFiD7oDR7TkAPUzvsvwkLk1ZudVs9O4pbglSSf0Nmsj0MauItPAUZauI2
+T9xZT5SvqNcCQhDxNyYb5InHq0GdDzEKS17zuYcX1LzOehAlJ+6U2/B0UhDFyym
olgptPdA1RyefO2Roqf66MEtbRGBdsAqjSUgGm/bZNA+mWnAZ+OYaTSpkNH3XyTC
VSm6Q0vtOSi7/4F/ht0/7ZxwpgHSZb32FukrqWz8bcRahD5o5DjdKAFszgIc9sXf
fhv4vBt5eNXRFsw1XZkxXTS+v/2yX2iXV2sXv4/Qkv1p56S164F+R4hK7WDtevtS
MNVeONKh6HnfvEl4Di6soDvS5BUezLlCiBfp8se9mSYC/zX59XfhxgkPVM7ZlFO+
xaYcm8mH7JMVH5TUSFyrDbAHnG1ELE0pi9Kju8woDc+u44jYtRjAjKxPj201+Wzc
Q2VihyvbZkpRS0Z9UQcqmaVLVJ3EHPZWQNOdPj228YAhgb+bq5x3w239yIeq3Pob
vmxIJPb8iff82vM3pjbblNbOng7iCjw0es7PbJQu+J+8LVVBuk84TKHrkYnkaES3
YfpUHoecghUsA1AbtMAO6feccxBdmM0aDdX0Ly7Snfm2ZRZAU1Sz3MDG5eKxuhYb
LPtHwtE/qnD3QjhukH+xMejz3Tzwda7Nsa/rW/3UD+Up04cfsG7gnik5V/UKWCul
GrhDm1WGig0qT4TjLihKVUjNFtwVdYbO/IUcgD+H4mr0701KsoCCrajtI8nnWhWi
TLF82usZu1QDnegbeSHljTcGovqjUr9JLuaryROrq8RGbjmGHqokTcvWvTJO1a1r
nB2yUtu3rTGFho2cSLH91j9IMevZeibboCZ4ouB0ad4uSs4ZnaXTYqJg+5eq06th
NSmanOPOCDnhn/PUyTphezWJoOT+5hk6X6/kiBZGEd2kwXiQEL2uNRji9LhXOXt/
4r3Q0SzhhbgfLvymhMiHVn0j1yt7obptVYfy4knpNpydYejc4Ttb19qRSomd5M1/
mnAdnHpUNuPltw2UiWYhX8QnqkwWB7E+sNd6Sh0AbiK6oCLcJ4MW/WGNZbhq1n4y
NYqvG49WrCMIfIMl3dEkf4ewUHQemZ79wq1jYn6nGBiNna1MQn/6gfDRXgtZeImC
z9ePmYFqv5/tukYD0NdbfTuTM70a+5zKY1X2iWk1zQeSvTIcgq+KE3a8WRx10POx
KIskxUkJmEOncikJF35FVj4eR+EbRcklVkq/dqawAKonupZo+5WIkFBq5c+Z50jd
AuUqyOgOwJbt/wV99YgK1mjeN6KV5l3WUvVEqX7s1TtnonSJEkbqpdW4A2Sgdu7r
HK+se4RQT17/NO/EqfbyzOBdTSI9wAxOOiPSRhb/v/HsGMqcBjGwcqbfhTSfa4Id
69Gqn98R80cZ6oKGASj/GaMdC/usdpv+9h75bnDE940ziFTaab/OYwJXy2ZQ5/7L
VUQNz1fUAAO9/VEIVwOpFXmd5Zk9QKKPHgiIMH0UvkjS4WypWl1rQLjx1dNZ9X0G
SsVRVpnJxyz0xDQTvh8apkayCotTfOuGeaaX6vR19kVJqUplk3Dly5wQIQZ5CdRp
ori+84MniNhvurXXQVlSURHemepMaHeZg5hmVQ0w5L/acr7FmLM/KlKY1b9577rc
Xmnv+E2oqSwIhnPCYXuI++onMtwxJMlWTUxvw2w3fgM3AgjYjy1M+UQeVV0930yn
vo2VJfIWY0kalWY8i7/97REWy9g92bbBMjJYxk1g+HXhyMyTln0OuMpnkuRqIr0a
YpvG+6sV5dhBmwEijT6EY9Dvahge21rERVkfAQpxBStPyqReFN1lUEVFXqA35edf
biPkWD/Eh0b1Op8SUt0pnliS0trLHAporFMAvRJvhoKyonDuTx66sgaKVcLxUIeZ
MGGLorN4SPPjvwZn8sOm4j5Ofq/9IK/Nl5/sZ3ePsHIrFus9OGlXtPnj+ba/9O15
9U7geo5/c2V5GvdXqm9A3l63BhnUlTRdtcv8TgmGDAgj56Kq/pKF4Afxuv0wt6zB
IxhJje5MpOQPEgII9g/BpoznAfZj/sLOUmfFDNNEE9j+GPndNy6LBvkJR74kjwoi
NEDydUIDZDDDcI2QP6g3DUCBg9lprNHL8v2WArowIxqkV036KRAeC9sjZ9/SCcCD
WgNQECKdZF3Lvs3Z7f0u7HpO/aGu9l8u4SQansEjgLjgeTi6vZYQZfY7+ZgC44cz
ZBgbgkUIicllw322rzPTareuplaIigpjhJCFDbCZR3o4aIQNgV+O4+IwD3CVbdSo
5FPTfRaNUYFEdEXUu4DD3ff10cqQciIvN7nRURuBkcsXJ711OZtzYlLeZ9zzcVph
06HXddmHp6RuoCTEHr56DzGhVcEB8vMXrG+8Rp3MU6rQPuFFPiQLmYdONr+506Bz
PO3xuwzRSJ6lpgx5TufK1xD8g9g9jGNxMFCf1z/Ssctii9tqPEq1qGH4ic9WFcey
guQJJufkAZOBbXm1nu0TGd/0uRHtS+mYQMs3NOf2ie8seF8/rkq+cOJnxhbZBsEb
zC1/H+IZOHSGJKkYRpdL6vNyR6nmX3YaE6vCLXAq6GPV5LO0gV/XjT3z3Gw/Dx2b
jkFyZll6ypWJ5t8nwCFRzh7ahheuFNivABpIpzPxykZpTu2I0Cskp3zwNBxYSGO0
MiSGKr+j8pb1yuZI5DOC47Y3BsRW/pZQsD4ninGM8OdORvtsF4ZyTLuStoDuAcyS
KSSCL9KzvFFEPoYPUvZHmnm2va1zAy4mbpuOu06/8iuiz/OxjJU+ph7FT7ZQ+BXo
615AnAa8rCliY1HG/5UvDIBvQ0cI/7IVvOpZQl0eITZr2CA2B0Or90vU+Hm3lZQp
6ooumz9fjvuM8H/3TIonlfnPSsfjKkKIWNnvMl32CDbRSLWqh3PWhv4fSVHpg7gx
4gBr+L6JLlV9m3/SeGxLXqXgCYKFc/eOl77E50YWIxfq0wkxWkTjM8WFvHR4yvVg
pmZOPM1GTKDjJl7B7WM3Hydxb4Q0Pt64GTwINVl+2CSyO14ZNuuDPyTKhhzZ+GEY
QF4RmSiBYoovX0KtmcqVJQLTJEbj+RtkIdGksoJ57GFNOfJ/H9LNvVIZOOmL528y
ehsgk3EZO30IQXmGW0bfSl/QoL97IoZNOWO4Mu4T3XQvdRbY2h0kcMImHsVWLolC
h4xPe9d3F9BmaRE7pOekLIJA0DiUM4znJzagvbwMQ5BYI9XZSM2UDAHh7W1F4tGO
QTKs4ebgN3GVFORwwj2DeOPxarQSv+MZHjaWm5HajZAZnqF+gOKfnfoDyCc6vG69
UscH/YJ9H3v898TBOrK6PDAH+EGQ4r/dadrCg7YjN90x1ry071p5UiDpY+u4MJjY
pyUCsQCRxfzzfxvzD5F2IdnEK0RhGdi4bPQhg/ernzqJfHt69v1XMg42oC+caz8Z
y39PEQYpkxdrggQiyDxcmp95nII8jOM4UK6plxZyVPVQ0snjNKGi/aWb7ZPNvA15
7gUDyz5m5HB1hpMxhowTT9bjo82IwLty/nFmfD7FaLjq6P1Y9/r2o91+HkSdSyBe
9ZDEDROEy9vDyXX7cnA6OU6zKmxwCbcMtcv+SbBhwOlwQRNAZv0aBerZVcye6z+3
bT/YK85JySRTdKd+Yo0exIbuzCQmzPlQ5rGj3vhicBvF/HGge24ptvYculLbwgq9
8LHywkPqJ4vxMMb4MmHeJ1ptgCCP5pDB09bOZ4L7kH3lRhhAuJl9FvBIkCd8bTTV
qQbI8QCtBigVGbzLCIYpao5vfjcClxghlBoLzoZtbXrOggnz2ztaCuJh8DHcxzdg
DqYuxnhB6F1tYRpkFSe2fGFYeAHD6dQl9IXltmzL6V0TF6oXVAR1SkfL1w/SMKwA
5hUINDT7RtTE2NAC9Gex8rpitmtEi/ZE3a5DxvU1wm4RhRACudxkrhFxg1y8xQok
55fOmpGoMUv7wTXyrFYk5g+gPtZLdOyVYleWq4aP4UjqIwrydXVjm/Xf4wcz9FJy
gWA++gfFnGODpFEUZDdtX7Sw5s+PC7Z4QLwn7W0X8uui+Zd0W9gKPNdECQScSapZ
9FsfG2UTFObXjT3DBUAPnfSUMnvKnc7e7QZ6gXX32CP36ONxmZr0p66c/WIVnVTS
VhTxCIPieS5aX5oH9tVjxmYwSEgGRtKUYjAYkRYD9JqnCBIL/NlKb8/l6XTKk2/V
7TcKhbzd3u67iig4TYXMcETmQmQVOWqmCZXyRLFl3xWWee6nmDzCJtlc5pP+JIds
QKKcbIrxZ1+19k8s6LSaWiCu0BaNPGgWrDiE9URLx+bXyLuJFEwxVK1B4/c1MwJG
xvA0hH24zqIFYWWrDXYJ0LlPYyu7dQOeLmzr4rvWHARro9Vgw+IxzxaV0YTz1FLm
HoE5hXUtrbM4iUWwQCc+8Lic/juZTAoWsI+QzpFpjV61aDM4OTNDscg1pp62hsZ4
RmJ/60Wqpb8YJtkSPmdKhnGTF1Surinq6UmMN/hvfuhncm8heJ/8oMCyzGilWDl+
yEC8Ebi5epltvhzqaj9zdtJaBMnkg8BsnX/ItXgxEJB9n9Dnv5rFrpK44QLUgBHi
cMqGmg7IxYbEfBowT24aKq1LsoPVXZyum+JxX7/Frm6bct7yV1WGjcaR4fXtXXpJ
2AGcroh80+AXQ7BrVCHqcTGqk7Q+aYNmv+QN+gYD8uuiSTaen2OVQuBeeB2Tx2Fo
5TXHOZJwRteicqxbgwIm996XEdve2vzuupWsiLUeQgIibOi8eAV6Od8JpxMVU6Nd
yNrk+jqIpAudWCgo9gHCmjyan/a+lODDp4+QjB0qRNb0s3X/NB7gPCt2RfUatFmB
5xW5o/0Q8cQwlBcNGj4pXhOzZ8LbT7l+4U5Wc7CWF0EVyHkyXFOAYIBVc9/wVRdk
XiERddOodxgRpcbdOiKGdAtl/sRINGVg9oNXbRaTSoSkKmXeAusulZugGkEirEPk
F/v5pWLNWk7iCToKx2Jvs53HZ+7nEHGQeGc6Zz7AEI7MG/ipMj8F4CsDXmtpDGbI
nkZDsInt9Qm08ZCM0UCZ7AKz4nDQNR0PsLFZJNSmUw80k09yv/4NQ4J5KKALif47
/d+FTtM9fYw5LMUynSSigOU//Z9YYHvTIXVgeHxbbXHn8ee3LevOS4koR4V9Ihyr
BvvwEUkg1pJVjHJuWJudYXKBRHyHfFXWvuMOiyT1FT3yDIKwD5c3OqDhRKGPZC0W
cEQn7hlfJ4zA3LQztdcTtOvZjXEO5GE8BanV9VfEjq2OGPTz+sd3ROZWXv2DRFED
HpuVdEUV7bROCbURKz1+Lrr+ucyeTC1/Ru1dnykTZiEAvV4cN4Usw+awiyuffKwh
9iURhl3u7QzmbLI8HSemtV+/Fbp7gsh8DBfqAF/C5A/xKLtEBITSVauc1iD0dCHZ
UBhMqBjWztMNfyUokkSbQ0KGx75SH8NsY07aOHosVxhI3J7SNCmNICShfulAFp3F
yDbhoyhsZZVdnZ5oByPJ5jXksRHNBtnax/l+m9UZmWO2QEwRnMFxI6sdGntpeLBH
SRysJcPlrW88p+VeabboZ6pnEwnJCvAZ1hZU1pTiaBPELvnmarxFYt+JoJrFulg7
i78UnPr1nTq1vwbOPVtjUB/c5nuJWHkT7COOZnoYBaFAfpAokhYMVFUxolFntc0W
xkHV3oLO3+znq9xSoUP28Drw5DHqz1n483OqV7Qe33hQGtv0ZpwKxPR5KFnSayIh
b/D3ZIzZPTM0wtwjVPpwBTEnQYPO8E2k9/6dk7TJMVLOZWrXSYdKNdprrEtaxB09
+9llkdTTBdLOtTiP37wMf+6uBIi07ucsQPkTrQ/6t2LEXK1JjsXqhtexSvXtW271
/mFFwPTGeJblr0RYIkdSs4EIM3xu1puhC2vfSs6rm+hEyEKvwWelZv/IIxXot7s/
0sdQyanJbQvyeXS7AykKbquWwYz7Gcse7n2P1d0jKWlNjc53MHg5PL9ZyoXlJGrF
JHop3hsFLEwyhQEzFCpFqjHOvQ8CSa2/PI5jwmFATjbWx1vO4uaocvn3fyscXWy9
VVs/oOQi27OXWnc4Coc+qd1luFRFwMJHuH8wwCby8Bji2NsRAiQFhRdniVO45Mi/
VRPoTNRdatAY9UT5tUhqXpQ06v9izW0KG6dvp+hfJ1mKiVjSLYK2pa1f16WeBQRT
1MGSsKPJfHlr3hH2s3DLkx0YWJ2ZcTfH2LxEw6Vq9dFgPoaRUR97iDYPmbIBtSMH
DJOLtwAffBcellAepuF3skMXc2luaHPc7ZxqL1ipFsJXaGr6BQIlks2JFV9NaPks
+lAsNyhaQQHZzFwJUHt9AidYxdy2GQGMKTJXuIAYiW9DQV5XGTIYToVQ+LU/4bfw
d5t85gdKr7DHyAKeG3BYrDb7N7V67T1fMdIMiJjYcOvJgkgVgnz7z/yCZKQ4oNEC
JD1sd1ncaXq7xtHMmW4XWxatisyyGAevluqpJBIpsoa5tn+pw5B+Eh168fPKAeTi
Hx6Wnw7j2nEpWAJrN1C8AABggg1KkRsEPbjtkWRK+eP9Z0Dc0qDZ9MFvPov/PyH1
L3HdiVpMGPnmCHot7DiWgZ4Ahx7mNzlMtSN/ceF5uYL3c7t8qGg5IVz9V6TC76zb
gbv9xNbqGLOCnTAa8rQCOe7V1FZTw4jPrCwoiOouKwxtIHx9QpZuyI5UVJfdMew9
mBEnlz4esHTlt88C3dpAPsbasKdgz0uYf5MMQByPuupxTcG7oNlqxRjSWhEic6WS
uGLFBcZouerD11S9qBzQhsRmT7GVQQ+MxrHLUtpJJ6t16+E09EC+4VhqoWgk9CiC
xWzbN5nDj5RwYguz94o50hy60+0yoMuR5Fo9navBwrJAPKve12aGem0+BEx4/0DD
a7rFhG0t05hqFREApJbmK9OEnyjy9clWDEVK4WJsCm8pDi3llY8wUEEnmbUj2kqG
Makl3JUuzERWKFR6qhOJJWszNOFLumgllGqGUzc8U8GRA9bZpI/I7NhceYm36YjR
yQoV/XBTyykJlmYyfirkxpuUPsC7SELpa1h9vNLWELSDvHEtK+3/N07X/OQ2MYAD
jfMU6ThXLKQXNlJp72sCPQXoVfd01D6nAQTZ41nDNXmT+SVGqYZOdK+NhZy/t9nX
q28CmL1gq41lb8m+HLAHyqdD1ziKAvnJc5VuKU0Qw7IaHwXKlXRvS6QAQ/HpVxUE
3Qpos0OkJS6f5X4mEor0kQhQQJoe38ZJd6DLLW7sitl+3cTxkUOWJJYGOX/ll5kv
N1FMU+V9SA9uA0ErV1a8Fm+KTiWdQ55dEqRVOpnnA/Mh+yjfJ6baZIFj3Xy9u2Eq
2T4+MsZYBsq2PQnQoQTCRPTXGmxR0WTvXxBcOhp4YASZ8EWhfhvoTpkhI1smCt94
yEN3NQIVMG4bIe8/Lsvs+HsRynZJZ2scwbVMoMYY6AKcOzYCdyj+wVgrKpcagnRv
qfE4QYaHVCh450eV0QuO/5RCAhnS9fS4G+7YFmF7/DYVy4uBhweppySgrI00nQIL
c09d25tIbRF2aPBnvlsmnI8wOvcPcKRZwM3ZnLTq/KnWywxEQR4+UZbwFobAiEGR
a7qpVh1PINnFxOsADecQ9p8KYbBbPMiQIqtIcWjEcTzbuK/xrY5lWsPPNYsvxmex
+NaTs1ikfM9QpY2flJSv7lydSQacZODQ69v2+HT1ktscO3aK5PtJyLaulJpM44O/
6mjL18Ll3WT5tV/b37x+TW83ptkVbTBi1Hx8DmDj2hKmC0J7t8mJ3LCI/u/fuWlP
ZwFdt/i9EEqDasCb/OeGfjDJcfXTyXbnMk0KqZPYzEasCjlLZmmRaDEf7V5J2zBn
EyCPHmJcJlJX4SajusofpjRpGucP8kzAI5g9pxwErgjp2oD7qc8eamEZwQEALKeZ
BE/qDAxF2z2VWJ42nYKWl1lbvaQHsYQm5ccMbOPN7jVmv1L3Ffb6ITBOxzbUpSM5
wCoZ7XqVuX51fRoroDtOKv4/1TXmAy6MbRnyllo4WIOOy1H7IuW5EwgqRs5EqAnx
jDTH+Ivij1tELiv7bXQjwQRn7TX0NkFqjKEScsxRQ1bfrYBkpaQvasyUNCbeZw7a
+ciU479LkiiUeRT1OTn2htdDupWzAV69vW1nmjw0D1IR6SZNdFK2q9sdpWuQLD/1
uzbpnTf6ZENluS7xopCo38w13F3uf71lr+RQsJbqr78yq52dRzdYDpSlT4//pgi/
MDxeVPE7lMZVZtiWKw4vR+u0Z1hWlzV4lrKAYlfVu0P5EvakSuPeq661x5/15kVO
Tqproa2akm4hN10NQn8ce4AwEaN02jx2VP6vz9OlLxAWFgH1pjqBQ9E4lgdIw/yw
Sc7YDOgqgUAaM+2NuqqLQjO7pCPwxtl7stc7UxlFpQ4sP6PljyaERU6GAVC1/crO
PQ2cXNHfZA6wf5phnA0Vww4S02zx2ofpuXP1Waoah/XLvYYA/ilgW14FfeNFps/y
k+U8OS2Ui+t9QGSTd9o3pblT31+2U6GGJj6YVMoNsNfETm2Hj67AZIrFzBQwyhm2
yP+6tRPIXpk5Z9bRfio/RBXxGjH+YAe/OgjognyA2E00aA28MRmQjiXoFmRIn1gA
5V7BO4c/zMFtmj1RY9IN8CMGHlS3NVUN7h/7vUK6jxkKt03KftW+SCfzRcE2Hg2Q
B0Dk+wQaVhPpu+uamebBQVxqg/MRRaHfALuDLXGJWxzK7nCAYFn3ixSnVFFY1pbJ
MMRdnLTpTrsj5P2Gr+JIe7oPO3MSTJwH3t6KRbU3OHEjQjC426bWhOtEqJYFy7aH
ETFiKA7LBqyhHJhjZctNV5PlR4pD/+GiC7vvWV3/uoD/rbqfiYryRqC1FFrtZGC/
kpaTGHmZt2o0lehfh4hx9LgSL59SUmKzDrM/BjHmsE1XlGCxgVp/fNWUZwfBWkwv
ZPEs7eTRmBkDk8J3gVmGTQoz9fpaWuPQsvb5HGQqMQPlusHpLV7mr07VrIj5vqQ1
tBcxuK9C/KfcpqfUBNnBlbICnencPeME+NU8+Th39my0o0tI9oH3WeX+lGZW0g1G
52xmDBkLgMT65cw5cv+KKEgIoL3k8LUDkvHb1y7n89URcNgkSjngBX5CvMjOoi27
L6qpGwTYSXd4bdrrP4KlcSMpzi6OmN1zRlglDwUHYbQrijhBrcrCro6zj7RW67N1
XCuESrFHYnyo2o8mxtYvpPXQgwo9HnHyeVlf3LMi4ZzjNrWj+s8ruT5fi2HQx5R3
5mdPYW39vdB04Lahn02o07Govme9vU1Xfptpcdq/lpqZ7cNdpExCVsVNmEOWlb3/
U//wTXxbpAfz3VIM2IdAbBg99FFtqfy17qW+2rpl9+FO1iFRigp5coC4D9JkqkZ5
3o1Vstyd4LUTo9kPTpcHcqWTBEZ3/4SuO64IaDQ/NCEoCAZtucftMrU+9EX/4tf9
10lqZMUx+no6sjtKxXkBbOekttenocFGgy5D+Gptxoy0I66cU/zP0lxOIERR/KCg
Vte4OXFxRdrtW1JDuKIHnNlYv0pdz41cm7pWkjrBgIQO8/pYwd3zBtYIp4cLnYgm
1lPz88Po/Z1MjiCSU4CFrTIIcwSWfn+jCO8fn6W+W+SC86upY4b6CQmEiat3hkXn
wgh2zmqTsdutFAIlFo+hOAzlHvYSiLuEnpdLzFMgizwbTJ2Yfr0R/QnFh5tXJQX3
qEFNfKxOTRo0sssmVu6Z/KnpXTrzN5FclXl+J3RiuSFT5/MiMUHt29epn91XFqn5
rJ1diSOHikVks4mORC3w3w4pseTHZTeSWsiprpGzMp7KqDjsZx2mYQivq5uIafY8
YvF2ryFJUDovQ9/jKUwLe1/HzNaXp9BO2pgLRLaaqPQqh2KVwTN1W1Ce65JnRqUN
ckDf31UQ66SV/AHIH9NDfuuIO5Se233odgbww3Q5gMn8PJmxX8a20LeniqKnZ/of
QS/8+hX+VVNUYyAemNqgWmreGafCm6Z9df1uYvS/F6CdK0Sw/z/y3eIj/siRiJJf
HeJ1wXjWe7D1+HsiXgB/ziHl2uH4tJMibB0vuf/N1Qby7okt2/WslamybsivHPpr
IsxhNenkri9DXmX/f7mstg9VrwP9DmpU9uabjxoXlEwYzskI6+PqCnUPmMLxz3wU
WUD7WLY87CRxvB8YTNEi+fXp7oOOP3fq8XkkWvHT35tbIbRW6zF5i9BVubD5Nhq+
jwl4NlsQYa7rPBYGRiYMeTJzllv71UFdfebMqWaFIEh9pRVg8R+zofnUrqy0ntUF
KOHy+kYM3/EHC2zzQyBihndN0XzRrmxu/ILvHhrchqsvtp/cLNb2lSefQ0i7Q4Y7
+ixaQYFBjGEdgqsj32C3k2UNmkFtf/X1IIrvtfdY2FcWc05wRqlNxZD1Z8wGZn+7
7hxIsGeWQ0zavKdt6KGq5Aj9xNxvTC+u3v4MAPyac/jWlvbHZHiHFLq92tgaeIUR
P/h9HjTkMOUMYM76AsqfS8HtJ1Jc8Uc1R8gMP7k0UmV0NBjr/aQUebo0AXfpWWNn
kL6fBKyvhNE1h2A53t/Gd7vTLfBcORn0H+KG0MWmako4i2hPq6lvoM4OgMfCnQA7
kBD3oqTbxdTnT+zaxEmOGyomwPCXPy42z3FnAVnUP/iEE4OiWtiPcEHzHASU+FjR
oKF88M/V7z07+EPrja9pH9jtucF9YcbecdYqjlerLvH6ICtdgb2DE8VeJuSR01bo
9k68lPiYtF3SvY+BfojHmV/tlIZZE0HnjOZo7qq05t0Xtj/WaHALyKp1pvjnv2V7
gG/O28ttzyDpekrUwwwXx3F0d7b1XbFlP5jLvJBUflULYdd4A0vxY5hUiLFxBmal
YzWQyZNe5Kxc5FBqWxMK2DJ5J6Na9QazsHZZ+s/HNSPTESmVUZgU3Qt/aIZGzl0I
8hBP3ZwGxMRF8RhqDAXTgNgBz7sk0/fLK6eASw1wbvliiYmljXSPNqo3yTCcTRqH
SAQJPnA53M6/BzIMZoi9/0+W2Wpnks4lg1ExR5j1EVQqBm3EA/JxmwtfyXvxgWoc
vtn+yTu48p2T+JRJAjD51ThfPFhmpaLZ7QQTjTuG1Gbsy/AZc8x8Dbj9esMV3Ar+
DNKzCT9Es+6qQAWY7NtKKDSUHhTeKCIx0dKJ0Im7IH3/wu6DwutTgFNjrJiCUwlE
EJVrcuFSQsrvL8gTy92wtiVS4jds69yqKlVNcyh33WWSTL6kTpgg0pwshZC4ZTVc
0U67ix8bHJdb/wLCrqp3gBQoQie9GBaE5Fnx8KPXGjR7ZB7wVU4E/2SPwcNpmerr
QY4+8a09WsTWT08tFYgJzmdk7EEUiPYuKyq19qpkGorG9b1CgiyhUmDcEmHO+Kr6
QFz82JVJynK7jV7BOwYyO+xGVpZU0I9LpLnGi270vcka3nWJmtJtb8P+7kD+i7bh
3zj+GiWdHPahnWNR2Voh0A78uSkib6IzV0en5VLJqyxYV7HKtKAU+8bC5qV1bJat
b7iqmweJSxtLHWUh5riQ72smLbVgAb/RQ2IF5yp/bjxsCyY2i2ozg5yI5d5Oy+s0
C0fMviAQK/DDJJ3k5AEHvAxU35BYYMLHWm2FfWcscZce9LvUvlnY7MSatjTQTxhN
ygnhw/oM4CtEzLHsNDj4hdXB4Fo1qoQ4Vg7hrEuYqRmUyGHq+pLHBNZJSJ9cWZgW
ErJ6aWJrVoi9pP1/9WvlzQouzoRXyHKvbWXWXnU5RKIrNyVGR5W/3roZyj083o/i
THagMnivsV3DLiwQ7L1Dtjt1CdMvfTgpg+YcZBHWUEB+0MLsSlGNuQq/Rr738LSA
thWGjz+uNFtnSIYjW4uglcF9wZJzF+Vi4S/i169W8TUrqXI9EtMtW/E62+S3lDAm
a3qqK/yNErewYh4AAQGSxrqL+3ynsGuI6T9RM31b+aLn5Oz0oWEryDz0wjVztlPK
MRCtJ446Pm5/FPgyR9wFBpmO71hw81VM2UfarXIf+lI2rwrhJLfESj//73Q0ZjH8
zyIbfnJhAekGVoB+jxkBlKit1kBtEEJ3S7al9qjdtsZHJneqXy2Iy18poilh5gqK
WMniMft04VJ54xdGrvOND6uTBdT/6WyZD7KygYvANnZOyyKjqvhBljZp33Q9aylb
VTZlPSXxmwkYBIm0423+clpXcqWiIj+fhVA7YuZ7ekURrirgqm2E+vBZ64H1oDEX
Fp3ea0uAnfyB9o9dw2yrD00z2765WMGIchBBn2jWjY9uJAiUearaeqPeGgUsgY6e
cuKgXgS08snG+I5eNrG8vo5qXyR8SmERvq012AJ3R9Misdr1dvEvYRBVrcfgaCof
pmh17h/57yNUHt4nv+aZiGYdYEH4oIKJjhCTK1PTm5QKHOauyrpsAkeRPMeoyOGG
RhungKCZTUk9M6D9SWauVeM7gNe+rrJNTq76g7QqJXm4pQmdPUO7tFy9/SXomcVA
kkAg0eSOat/ipcgIkUqfN3smbTZyC9uH4uHkk/NczLvzhfpAVn7EdQH4tUYm1RcD
HRRT1y8LQCUpbojBl6lHY94/oD8LnVFJ+UKxxCNr0l1GqZc+s7IHZRVlwLKA+JbG
NGn60w3HhvwCPRPNtpTi02OI7aO6e19hPh+L8bGzD0d7VZcDL842I/7TdwuwFugC
BuHyfaVYO+8noazspunvD9HYghtAF/+eetRVZpNZxbpfrWYh0Gp1/dq/FvyKUBOD
tiEJtMv+H6xt7f5/LIZGWAxhZDRQIOJpuKVOxeCu08HOmz88c6ppWnvW30oWUvsG
XHt7vliVMP1JrdFVIwKBD9jHcT2CaLhhMXN5bdNKymWunIjNknLtoKA3qM0VQAt2
c7D+lvHwprv6eJY6aaoT6GX2oy/yPubAdueow6UKYml8DQvlFFXdbYbnMDf8XH+A
7Krfv21lxkdjpPDS3KYORU9tcjNc0TO215+s0wjag5KV8WtZM+s0+UkXTBH3FLaL
93U/qUzFdLPj0pZKPMuNgBGmVKknu+B2tEeR69Mb60ylZ+oH38jifvmIVfNkB10h
hFdyPSt+4LjYym07RQUoC/coXPUnLM0C07mv7NDyliU6BLeSZHspOx7T6uhlJHG5
1w4j6aW9eDlkkHamvSWAsEP0e93q8CvDgS1fJPGqvY9mhaaLFLVZHuyu9yi40LPs
4X2h0fSaJB+jlf7qqqDRcD2X47KgLAkMAtB/ZmWg2AgRpHN5AbduYWRaRWV20LwL
REFIDbeU+MjYgzo+q/eiVUg2SXxUu+FRJCFM7ubK9cCkSMr3U4wjhAPa27cJ88Q1
OSdBXqMPLAtk8+Fcj9mb7A8vypZt9HKEHkWasrJ8VL2+NDnWCYcH11+dqfR9lXh9
nHcf7XV0r8o8l0FchhObNjmQX2PFtwGyvn5BehoI5uiQNfl+lLq9c3bGVDME0JsW
vm18gTE4yCTti4mgSk5pn12KEiGurL42Y/AK5q91hnserXtZMKROiaMtSJAzghvO
yjdH1ci8gvCwnFeiStQS/yeSZBWHC0i3A+gb3Vz91NTzddTgpd0nt/qumZwGEbXb
u051RKlNJU9PmCotzAUziW4S40+jpBI2ot4CrIAwxBFNHEX0IirUCPLiaHMsjGVn
o+YBe+Vm6uLuYPj3/pxwmvrI+9wNbffg6bWvwvzxwEa9uuvujng/jDoO+oxtKmVS
o79zIURdi9Wz98rLv/xXhlKt5AeFYHX+cdNe+BnAs7MvW04wXBrFnjQ3srjSdtI+
dUAZNFsb8WNj2nDma9oMarrKv7BbxcV0X1vUQwJy6kGLwd66zA1iOs3zzuvYN+eG
zH1XUo5fCGZbaKtUTqOcFKuGfy5/jAVsy5TzZ1TXVP5ouajzPjVqQhGrMT2ft7fO
XHOjJ1w93POqkhQBd8HFUQBwWDO5wlOs3XxWQlc2uJNAV+lJZ/CuMNs8rGe/VpK6
FU6RlX1TYkGHlp8O3CzX9kjialEcvp4EYIyILZ1GBY04emJWvKTTvG0J7yId5YxO
`protect END_PROTECTED
