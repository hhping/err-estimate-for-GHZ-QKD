`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z6y8eMCSjklWaGiBN7i6DxB0baOt0SLZ5bW2AjW3Uvc4vgBBVFdnphaRMG5MX8fA
WW2RVpzxxJ0s7UdINmXD++CKOErvwpyq7NcJyln+9saDJKnPcmkE7GTjxZTNVJ5E
PkytkIwHQLCGgPvGUBWtszfyD27qAQWC7GF4FAeAXvaxMF1FGX5318ERhePgH9m/
42cSgFvz4HnO2E/fjLaYAvSBsInRiqWuYRbWrA7yvT3alcUZ1zm8ea/CgzZWdeqK
r0df08NC0CUNSVAhQVexCQ8g2A9b6GF/e80Hu7BBqIRxBPJQwc4t1wos0WnhX/Yc
nGmEotlCvbwDE7uTVYcHSMuruBxLqO7otS0McrjUENvvEjGpMWglJAwmVjHaMIzS
dhFA4H/i5Lar43Sps/n7vbBqyeCHZ6+AGci3lBIfmPjEeLeuXOhNRudS61goB3In
UjGvHfOYSSO7lSYCR7m13rapNUAHI2Iry4zM1zVbxYkcvXbfnhs6RMk5Ka/Cyv4x
OYHnJyvBjGwpJQNW/h3JRRJx+Hp5iCESe9KWdpZX9nRWO8FxTXF/x/h9rtx4MD1I
FP7Eng9zYhf8nkLsyfU3sRmXB40GubXJ9RxBbwAu0v09D9gTdphW48GiYWnc2MVp
BgRrbp3eumdXgUAIt9wZctUXjpCs04GbvdPUuiWXtdAJj/sD5+aeFz9/HF3BapyY
XkgxrMIkx7DoUYf+H2xLjRToq5+/CzWxJbKGmxwXLNSvNoNZ/F0GWnvfLoD+1Xss
dNO0FdP9pdT887jSoOnPkBSLzvvTQ011DZ/XPaTgBY5P9uoaejwgteC2Zu5HSHZK
+IarcurJtSSjqI6ZnogNTwzlpTvNjFKsmVRF54cUU8fCgDVrkB24MfHMKm+mCCS0
`protect END_PROTECTED
