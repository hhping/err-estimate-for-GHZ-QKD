`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O0FK8WkGzLiS/iKKjbfNg1o3iKEPvjCUL2StCJKRApxporcC4axz2sPf2Ct7wDWb
CLmz441PNQn7fDZK6/DefL7BK+bRpirr3Z6FpG1LUMwu27TpDc2gXnCEMY9phKwH
2IinyGphO/EvU7rNpolEw3DVSnFWCZIfSAOxHni/bUDHI0XWxopd8amrUFewximG
BQaBNmJvB/18L1eAiiO/9dkkxxqKNGF7lRMZHw0/tmaWPPWCYG1K+f75nnxKFn4m
Tf0EuPiHhFZwGNdncpGaEp/MmgE7YCL5Oatcb7nvnIKFHX5s7kWB6PXYR3TQ8MOS
CbJqSOjOlSnnp3m0q3Mva+/q4DpAkU5EUADzqfVppKE5TkJovlsibNjE54jLJC/H
ug3i+0SVX0uAJdwvUvRVoPsai4do36S1gXVWF6g4VgO8nyiDlTddzUzn/xmAUcAe
r+S9nQ+a4wgWNGQPpl/5kP6Ca+OmLXpQntBxVESKH2YX/oKkQv1o7ahQPvCkkcoK
ahXGwkgNPsw7tv4y3txpzyD10L2E0R9RvJ7HBf4WqQJk6fVQnFvJ60skTibHKQFf
luq7UN4BPZv/7VGHLsoKovmy5o2WGk6IY/rzhXDdi4mHqzW0JxnMF+n6HFFSBnLH
Bezg/4xD94uM4ofel7LLB+299cYy4T/r7UjCq/nLaa4ujwhDG6K/GOR9Xep9l0ti
Zwa/hpKD5eN7+Fl4aZvAdx8ryjrzGwzw2xGZmsls484K2e6PUEMc7a+jSZoKsXAP
0u1KfvTIMd92iQo+qMOWxKIgl3bGizBVCTwTS0IVh38HwzvI724HGYFLidsCuOym
hdiq2xtuNxoGpzZICa2LQt5Z8hMgS2dazPwER8Fz9MEMikkH1HLiKjeLE4pffmSK
LVCwJ+75sFFgLIoW6EXxrq4P0xGed6E5PlUnGXwwdAP68ZJyrEKKf/ygJj9YRcAr
zunKfnTwpKujxjKcygonN1SzBCuxvw4GwHJaZrxHTbZNLu/fH7h6etG+dmQDaE3D
32WugklDldiRL62Pfx8Y+ub+f5i8L/1m6iiZ/vODHnASvpIvbigHsPL71DbA4iKE
604xgW0bbx6EROaqHj4Dj6YjVFBhKN3w4mxmHgcj1AyuP6skVJKH8qPCJSKd5j0o
tJMmtLrA5A4HJf2iOsZ8u5GmU2okWq9lpKWfozZrh44ri3CIy/qWZYPXs1IZwJQu
VdCyF8j7uEZ+TljM0ucFvTq+VcxoKQ725a+EuLXBmeHzMUqWSgpVycaECJI8UCFj
cB8f2iwIvAOLulZYu7kkhHXc/+YxyZWHS3wnxZXv8hu1L4K33pVB9U+/o7rTcSIT
+R8PqFqlS3UzRoso14JGGzO/9NobkVvW/YOK6vDqeaFJpN1UTAKMW9fbCmCrYo++
`protect END_PROTECTED
