`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xUlgXf+iJOfB0wvpRZO/qmDa3GQNqHi1IkGgqfBzjj0UN/uDU2/omJXWbfF9cF0n
Ok3iVjW69qbPhHH/iGJ6dbgwN+BpW1nbLgDniqPqL98uWQ8KKHrv/ApSNOwSyV3J
tMgtAY0qSRbr3gEoJwBfobWeFCHoCbeTIngdMGEls07CN4k/UiGYLRWnNcjZkL0c
hc95BMOPU2WmJNiwQBgERibSqZOXBXq40+OPPNJO3Rx6wRJiXnaMiwAQtYg2DC5U
lyuBEHKGB2Ij87bvr7WRNiiCNdufEMQCwFwclTZ+Zz1dTP6hOlAZW3xu3OXmxCQ5
SkCrcoQ5dX9fCvsIp2GGZpKVBV0HkdrWkkfx0SiS6JhyOxFOCcpImCe0uBiUAzHA
KM96MCGrtDKqoVaGRuFDX4M8I7u/QuShFtIdz++2MLZqX1oc0ZPgmH/A7kWtLC4n
3MVG0h8QAaeiwDkWp/a1RBg2GQsazhuXAwpA9ueDmLmI6/FG8pc2cqiDT2pS+BYX
Geyo0bBvcZi508cmpcv+xKHpvIFlXYpHYlTFKjlCbiCzGmJZ3TFEwJPAxITwOmmW
MG2Pq1fLCjoq4jjvoaTnrTvoXW3erjvU6EjWGaywiOuTprqcFcsFzf4uGp9UveTB
FvQx7ZzGdouPlHLGdWWjLAoMVfAcYjU8rOOnDvorUhvlTG6Lqwk7jGXjXGtGsDCv
C0/ZxKzI2NLxxoEb89VF+FZCnCxdwffNVimJtyJFBYqwgYhdLCyPqSsQZz2uCZGK
XsL1jNExFImtOYsR21XUr/DrAgRvO4ndoODyUvgSglYywlIjr1fzSizwBJC6bexC
6btHlwNMdqU9i708OXhXr/m7g6WLaIP1vYsuR8/3vGG+Jwnn1J5L3I24ok/f529u
VVpm9dw1ISLdZN9XmocQIQ==
`protect END_PROTECTED
