`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pKMoauk/fI9eZi4EKEkibBtLk2gRMjjlF6itURWUBXQdEQoqsMrK/myrm0Vtc0v6
xDmaNaTTm+J45wCNtPNQh8F2ATBMi4unDa3leWfhnsVaMKKVmGsJYC/TARgcp1Tu
C4a0IEBJao4ZbhNNGAxCNretxmb8dEDI5HylrfykEpNgTrD+M5qv1ytyojXKHQjh
xS8UMQr5WaS7cV8nmOQigE7imD3ezN0RyRRAWTkq+/j1Kn37Z9nFRlSOUcwXMyeZ
95rgNg3JjpKld4rTXOQEL8HflmwV/vTvYdSlxNh40ntG22eHdZ4snOz+/588x+jG
50rEmoFVj+9PtA7/O2dFaIGRzi4XdmDUHOVD0TOx7Vvix8h8ybkV8ImutNBgiTjF
eM6f+lb8x/clLDyiWR+UfixWho48BspXLmgvZnGzHe67N56ArEwJIG4w4OGuirU9
icQ8dnk9mgKC7kzI5aNiFH1y4m4jd8MjUyx4+HNk/FrNotMYVXczqQEs/9JmnPCa
0W6XiMWXEg/5gOgeY+ADoNV//VRaOSaD3XV2GJIp1PehXyi5jXQ6If5VBw/wUwRK
hhFdUKrizoi8Ar5eraU6cA+Mq0PqG99wXYG8poeaAd24mBvtynJZRWckverWiFuE
K3akWkf4PDiiKpxdDeEEoldh3ysX4Hi6nQF75TVH4aR8+mTcrbbVNW/MkS2vRxBq
06W9g0xKZAnkQNvlLEcH5+y3//lQPt7lPaAErnp9bTThRO/F0nZIYIqOEx4HF42i
Vtzz3PbpDrzN59ix1mUaLsKPkLPxaYvpTc89LRTbbZ0AlGc+DRzh46a3Jx6iaE+q
N/ky8rHm0bJt7v5MEQgHwUlROboLnepgyDzweLPklPvRgboBfO4LZI72G6S+8f7l
x1RxWkJvGWormNDjRsE6P3otqCRoEfoX/bJP1XCcdvD/dFtPvbSkB9XHKMXDr0gs
Hjoj8R30B2IgnaYx4JMKkJ81riP8ckiTjX9FaE0EQK6QkrZ+dLZ/goC2KpfwtZZN
aMdOrRUZg/wfclf8eWi+q42MokUrwGieua+j4EHYyHXSor6QrpGujSrZyJD/kCk8
hS4+sHpNGuo7EOuCIZJOn/e6/6G1KdYfunlV63slRzaEfYXCKw2eljJi5kStp31F
aOi8PTkdwLDkPWa/7BFWCpZLsg/VNCZxSYng9Bj+M8dgK4TcJIBTfR1MFy81KIyr
zPh80dREEubsVYgDs1IIQHysMJwBzjpGlePggukyv+aXOBAYmtD3G/X+axRMs87l
C2gmRAMVK9YGNMmBCaUoK8EYHN457TMs7pu/BcrDqk7MF3YbdyQg/3jnWS1MfwU+
0WEcrFmw6jOH4HItvugsxPc0h52sEv2eWE97BBfBKhnAwRt6Ssi2CXdkoG/35uxp
kVzHdX0gUVENp3S//MjB1msU7/jBHR9Tkjt0EVNI7bgWG5Tsumt3+2i343khkMDP
Da/oLrLeV4kZ46Gc13zYJuDmbrifS/9A5IllmOnT7A/bHpkD2aDOq+P4z21Xwxy4
xxRFhuNGnlhM2HTIappn/707NYwaQwORMjuux+tG8fLo/fb9p6aNOcDIEO3EdXL9
PtdjgxGDE/GntflXMtngQlzLhxsCUtAcf1urbkTsBsv0YzxTh8PHcEZBrmDbJjbW
Ywp+wQKBzvSbCnMLNnR6Z7SiRDusd21bkx7NyQqm/cjMc5qCMoFztKHiaBK9q3Hg
X6JDnWHoAbEzmvk7n9igQcmAmf0RJ5HyoIFDgRcMnekp5v4C5pvSHAJrYMM9kTEV
i/BpShMt7F/KXZL1oWH617tdTSUu591NAQDytVw74A2EgYrvPR23nmV3v7zjQKt6
kD/b/TwNelDjEq0kPUxAhFzrSMV661NANaqk9MLeiOG4nzsaq1mZzkUOEHVw1zS1
vLLrR6m4n6Dkjjw3ZI3/uut1vvdLbarzBdZy7YNJizIRFUEwjE/BbE6wZ2982sLi
GCG/bdO2UT4TGgh9pBK5Sr71LbjiopC6oAkh2ssuPYA=
`protect END_PROTECTED
