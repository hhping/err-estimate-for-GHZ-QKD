`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+Qr+rER8Cw+g4sp72w5EliKaQkwRPZjBlUCGWc8U6FTV58jXWKgrHpTvN1QRYfaB
F6RMExz7jd4vJUgO7UtHP7jfHw+fsK+/iYZMTnTvB9NAq+f3a1pU0MheVKZHzE97
sJsMxv5Zx8jkkHmIm3/lEFbeubA2LBH9ZxEsVrrpTAyrdT9Q20bNcWJrFcea6cM3
PFo7zUztDmAqFJjeF8yYIipTM8AUJ4Bwt1HsdL4Tg4wrAzbzLW2MNaVlqaois/Zc
wlPP/cHxU6gzxXpg0NfnpJJWWojhSWJqQpsUgIfBNG+Ns1+mr1QARxpvXROxv6yZ
zByZTfWFGS9SBr9iNqMJn1wATrSmv3GMvYBX1o35tIG6jqTUsbxH20GF0o4jfWRp
J0sgfRkiKP/8vmBFor7w8vObiXrLtSV9PyRjUi1CqoI48iwkN39e2nXVaHHgsHsw
5jkc699cxRITt3zceDLo7r3COJ9MhrdrUkDJujwYmxjNMmydmBBin/+Y9HRh6eOE
uKEIX+4AEvsm++VgL9oPhoqScSgCkVg52lP74s40OnhGhc2SFIov0AuphYZ7rhfW
IMchC7AjlAuVHhLYgCWJkQ5w6fbEI8BiLDaDP4OJdG3GH4X0RtNH+qHxd0KgqbWW
f7opQbEjT7f9eXeasPXh6EBtxTrbQMpbyFx8mVzvd/SWQo3S/UZ0bYXQXDg62QWJ
795kPMtVW0i70fYF6J7KbpeYLfUw6v/PylZQgs4K0IUvDrtfeofzln7yu/15QEL7
rTvp/u4uqFuEzX4S/bgt/hgyAW5Lec8y5zPgpNGHSSRiT7d/88WVznwWeJXo//kQ
+Ns1jjnlqrdpCPGNbl6414/nyzp3qsL9lhm/2TqionJEbj4sb4OqGYtYg6L2EXM6
BUoY0YZhb+C/u7h0cv1DusdInWOxdxx++8kXNfHkTYxDo9YMrqy/6MLKbEljN+Hd
HwlNnTksvxkb4wAk0/ThJrEZK9A6HJzBGwhXCfZVdhRw6zOOjrlvOjC674zalYcz
mTwNUmI8T/8Soq7o7jsiiPveCzhjOlmiP6myhlT2/EGoQFnDiJoBoaLqbclEWmp5
aFL3HtR+zwrmxFkOOxpKn7y5bZISCKbZWBCb0CFro4Uyk/i6IeiMWrJgz8WTp39e
bhCH9XLAHdId0W9RI44AFqy/6qgMeb+uYCMcoxwC8pBO6MT2UfjN6ujMu89cBFzT
kP0/PtzlmNlV7NCaFz/otgX7eBNrUSDaSWfnfpGNV6mh9dOA7UZv4ad8bYUlMx5Y
klzMiPZQqcuj6L4a5QQVTRuBaSU8g+ZfOIOUm0h6IYNWib2FKzi68KXwF0JAzCrU
OabaEE6IZc+u9bSba3WNbnX18d21Yqx75b/nODt5iYxfDtMyw4Pw4Ofk+NTfrj+Y
etzLGh7DHkXBtWytkZUfFXK1Wgziag6jkQiwCROHfkv3cfiBtzOifhgZONRKlg1g
OMRCiIAopq4C4HPZ20tvYd51QcddYtOIaJGLeQfp4iLX3X6M80UAfzM9VDaQjqKR
AjlBFc3dl0i0Tvu4gOczxEkgUg02LYDTvZ8/D6shGf9GeeGkvYjZ8k+PIDptSsF3
WatZQvMaryi13rgvu6lmhsxOFj5UkTmTqQ9CNfL89AsEMA1ucgO1gJFowP7dRQiT
fJr0gghYZIhi2RKfcf5dlMJVxs4NP3lBEN8927OzBWiWjWL5bq4L8mZHc+jEmlvJ
XDqXDWS0I/NJcgoH6Dsk9gt/cl+8Kx9S/R70VO6Pl3dKO8mY3+dax4cftcLHFcux
oYGHaGbH6Kl/tLU++MtiOq6ldYRZLEwA/0cCB9Emn99W7p5xuYHcFhpt+Pyu0U/M
YBLdevL3hCGJ73k7lbqn+TK78iZtPCJR7Z1+1idZBC9qwHDQeJlHLzG5rLxd3hBj
DgZamy06tBHJHJABLLhRpHduWPYZH+lVMq8E6Z14PDrIhPJf+RgW7WbIPh0aJjdg
w7F0GuW0athLarfS9lQGOzk3NMHEFp7W8dvdb76h/yjePwaD+iWpeNLl5iAs2M2r
1ENgcMYUPIOU9g1/GN5WowahP9pPUcnXEGqOWRB6kIbUInizaKHwFgGZTeWkVl+l
`protect END_PROTECTED
