`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TaUzOQzLnoDJjlu4RYqc/BN/g4mRjQwk3UsvP4PP3bhKmfZr0jSD+lFUQtH9Pf+N
DtVtAm2zaIRqPUh9mbodUhAG6lbVYo4Vv1aQ8fC0JiZSgUU7ZLfFp0t2qlGGIrLR
nnyrxu317C3clcjkEYBSwSCoJDFPSBizErmaTyrVurb7YdTUEpmRYT3lySImPxKn
/5bHQunl6BFb/RLVblUbdLbqsGiAAx2GSLiNL/WwclKcjNNNnbPvRi9aLprW8mzC
ZxHYsxpM8rObpbcq6+BnLK0GI56iWvVcQfktJThR7qNKP0k2qVmnLroRueOll+Yq
1dVuBdihvSZsb5vuBdg4HXBScKdSye06VtPDoU2LnwlxL7kc4qhFu4eHusU2F6Yo
xVGn1e7KGCEtkKjaZ5BGEEXrmRHu/Ajj/Bf1bb1lc8akmvIHpheW8Z6/WW4b642M
zkQM/cOILGb4EkYkpTp8O7UlkPI36NyydJaNi6myDyru4rnzztthC56PvwrVGag2
6ej5JQgf/7rANQY7WUUZ93iRRxvLfKWUpCQyQV4z/6QTgJHOvSmOUXRBRsTqo9WJ
GcGDLuacUasv8RMWmi0i+6wIwa5mhepMGB1Lkg5/JDqG+0oUmv/2pIwRm4JrK/m2
hYYxE8GaSlsh7XVbMYQ6JjNDbokkMo2nbZeJzVIMtPudkoXS8+vo5IFA2OOWGbet
QncUXkI2c3Svu1A+B14ujEt0uQxGUqtcjsNW7qoJCx2At9zTlLNJOaClITw4RiZi
0wacsjqECtwqHcuUUe/SdkhVnVRh6ohD/IaGUh7wnqZV37gdPn9JpgqPIbCA2O8y
qAdl0i5gMW6PTK73UOT/Bb4cDiIWv4wCDYBBXsuBzuJ+ZiGqP7Ks87gHExTTMBSl
reYXAVHWy0ESrXRFUJ6GJ/W5eoTdhAkY/uEvGMSYo7I=
`protect END_PROTECTED
