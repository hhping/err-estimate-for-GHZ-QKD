`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D/YCfq3++PDnqvMsvHfnGxmFhQRj6+i+nGPpKP186UQcc5EGQi0tHU9lly19zgsD
YRLgl4PPXX7cwISkdOZOcOaABwoUQbaaV5rJ795xO0rsHLNQH4ZNzi1ao3cZpxpr
HArqOOfYbfV0qPd/9RhyhUM/6Bl8pk2VTe2YsmaPMFefw9XaD6riGZiZ/oPht/y3
5YCqpY2Ibehzwf2qG34P61kr0h5JIfxHyV6NPF7kyOsAvhN3tPu9E0/53FzAkiyn
WgzmPaHerLGl9ATmeEhm6/XMZjXYiwj3DgH/+qxOafEw3FkA70UJ+qGyOQAis5UH
TgMYGHD0b0udRjN5Sr4O804QP72H01hGqDkFE+fxnGaZyDhBCdY9DgzjCYA9ceYU
5FvziFrFDAPwB/SFlh+a3P3q0YNtniVWrWKfI/qqPcmWGxNLmgjSJ0BtvnMn/Zw0
M8P5aP6USlgRBE90I0ItsOiSbESybe5h+OpkN38cEMjG9xKsZskBlVfGT5pLzH0L
ZB7WWUqG0nezUwbw1iiG4Q5uR+yWCrEWqI4C2x/705yxfG5zmWkBwa3S9vj7h4CQ
IXVd/ialEe0gIN73w7Iujeiob4IQC4lutMw0xhykcW0C65bY3qcjgujLayjupHdF
jtJgKufiJaOd0gxn1IS5012Y44KLp7NnJwhZfLbMN1awFcC3VhYKUdf/NrHewkKw
U0p0J4U9Lj9h97zqxz4Y6ifeg+oHfBE7yWqa7LV57drl4Frg3easPC99JO2sZnj/
Il6qSqkEa2rY+y/FYoMXmUH7KyE/3WtXMDH6VAwQAuBPi3k1GMxyDKXjqusge/2q
JVMYJ7xpuH+4RBCFDYb3VMq+TaGnudYrWbFz/TCO8Y6P/vcFKZUd90L8X9flqr06
sNAmhmnlq9sW0RZzUITDgB9vVOUFn79aDbbyFPa9r9KmrPnEW4OjDl1UTmclRFKV
54SFyFLnS63+5bLwA8PYm9SyKXkKea2f02xTjZyJLsSmViZo7aUwADpeUJTBxWJG
5R5ROv1CEyNWaP1C5R3aPlsExucnCUSfCFhUJc2tFcJPJcHyyvo9v2rjfAfL0i80
1/yJ1f7BmRsafern7czbVs6TaqTBtTdZLd5fKuFbQt3ZsBzw118bAs/jvMoiLuJL
xtZy9V/5ElYeo/hFnqeFXMJ6zJquUn7Ob36UDgzqhoIghK1Sd2ZP19WdOg/BpIIX
m5eXcWL7Ku4y2zV5a4LMe1kwmFoClad7K8j1sc7/GqyeBnyCQTb3+QBs+lpgyQQg
UVJoBpEQUkt16lm21S87xOIoWCD/W/pbk461GBIQhB0ZoCvA64n3oUTKd+fEn0uQ
zQehDMVsxed3fpyEmmYJCHU1BfR9IaX2DAz7TuGvEWeO98XwRPm7rIFEfBL57VgP
p7U6lKomJHTutylljVH4XonviBj6a93AcMZRxVt7A6dCtl/E6HWg18gH5E1t3VW1
nPsEscQ3VtR3Ix8gkOMcYZeJ7+tBwPVcvS689IdSvYMo7cy0d8IrRKJXwnOaRFbn
2Qabc3A3xkZlI02JZjdU0QmpelLX9LCOZvJPXsVuKBVRU/MjZVBuOxOoJY3+LQ5K
TITC5fFMJLcTdw4AdGtQhv44lPqAV/H5YxLJ9AQMTZs4LWXiArwSQ/RsVGW2X4Fa
XVS4g1r0FPsIJiJLp0po0H2dYVUrLFbABznsRtLbYbHDL/4D6aKRsRGnArLLOZHG
sexOjjQ1rPkgElxr/WQTnKMxIada/gPfhYjDOHE5h/HmTKBTnjst9bSpx38jo4KM
xbb6wRFzwW3XdlsrbKhyH1/ohVnWlmZzDUna32iIfybe8IWwJNO/Tt1S9i8Ei4i8
rRrM8BKEXLv3jEHSnfti23JIqNCFT1pQIRavZpo0JKlCT5erv5TDddnz9sxB8BCz
Y3tsv8c6VuBMgekkMqI5mH5b4Z/uWQfE0qfpDlX+pDACI6otKRa2NsRTkBiSb1GB
ouDdGqhz5pmqRoSMOgNGllaaHamSinegwrOHlfGA3Fh2C5K3tnRdEUIQgiv89jX1
w56GM0sov+w42MDXNcScSl1IykHPJwd3ALWOXt4+mPWV9TllJqnJv7rOrdg2uHiJ
`protect END_PROTECTED
