`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nAc90nU4nZL/ZGBzcjgi3zFPZPbMAD8Rk8yXbwxtT5Cle6FIUe6g7QxULfm4Um8U
vCHoy/QzExUTlWGjH1gImDM5Y/sxH6BBqjqqRUqzX6jQ8zo98ds/fPdcQK8RKv0S
jTM7LXDISQDPcGnb2XJyhHlaN0rOCd8BNGS6H4YbCh8D7Ns3d8jfgBIxYhxKYfyi
JNmuPqg7E9eYCDQaWNCeQJTIJxZP1M4x/3dZX36myckjClIZaLJKfjMDoQJeaSKN
TpJYYyeeEJC2A1QHgQhPiCaWQ8+tG7blHRVXrPyzAElVSSUjR1dTIKzdZKiZ4Uul
mx7PTx0Bn5PDz9hph8vLbC0jdF2MeHNZCYrZEz1ee0oYdNbgPdhCnXh6Rdc8M6oS
dwQUMkOIV3eGW+Qqwd47l6vaZglU2N6vVbWW2XmaztHyVvR5IFhEMT6kETKhsaMz
r+J3fvsTRyt1UZBnRGzECqWuvtYy6qUO7xC37ZVCofvhhlzbf0tcUEzaHy70d+V5
boGTf27eSVcanIJGIDEvvclyO4npPofHQ/vwIrIibbTafCE+WRolTl7d3liPz3r4
hvP2UuEK69jzYHEkcsLnQKToAO6RkXYdUdsxUAA4uwLEEuWCyht3ASdT/UqHNC3U
75iotlABEesaPhl5Kji5bE1IFSK0UpUf72s1LihEmMClRKcrgwj23JSEDL9Gx79D
`protect END_PROTECTED
