`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
takxsXYYYP+Uv23MupQ9u4Rd0+apDLy6PJ7eplwlZdMBm/08VDkh51f0bpXyxvdD
Un6oihPSHpqpJMx7SnEuve/Su70IQDMSyTovim+z2Ll/98CDEdKuAXyudeEhqD1v
teltYGEZ5rQGFrZzVaOGXADR239f4GjSByN3cRnnp6OL1qjCI+AfQkeSoJ5hZwzE
NjWc+SG2J1KONTvDP29gBUbbNNPK7hmKPtzCU34QWM4IPRMoUVeqL/LS8Om+FMxU
/7oa+VyNEuZKEeDQE1tEX7ur4Kol7goKUtcVaZ7gOxdH7mRdETglSNMxpvnalHvk
rZdeKC/m6bqJM1KbNpvDzxHABfErhHPHKzc6FILNYO1xOOz6yRFfXJZkYq38+Be0
mmEirQ+4/kMCZuFBn/ZHhWEtSCEuXAgCBl+qZAwEliAdqlMwVtN/JptaREvJFI4a
UZdf6CX58kmZRMqOCVGf8WgAnwKo9Z/LLeDcjJCpU101cqNOQJPh9BGtDUt+m4nW
5k7/LamGNKoOTzcFgtr+8k6DDb0KIOzHuKKyiCYLEXpMKY8f9djQm2iFBlvgf7mO
AzcVdqn1nIRxBe50xtyNp+7ge3UwkCgWe/HzNG3Ws09eV/n+pZFwbn99pvSIuKvg
g8HRZZoz6I54ba1poWJlW/G7oQO7g+fOsj8ZZBUCi7KYWqGqeW8QLvvgan/zvLS9
Mf7NdzSSdVsm6jRmw9JRpPv6j/aVJCVGiA13VQFm9jiwYzb92BUh0WGFs7VTBHOE
9Hx1pfJELPOHeYK5JMp5uFWjwnZ3Z3/9Qqvf9MD8OkP9LmLHuw6cwzNEpJB8RdPG
0IBWO5JH18/tylS5fzwttuJFHlsXQOn6oFJ8Gm8/dy0QZqXdvAiUDuPA14JOYeNs
L34hKk4X29RHbtu6kvOHZXfablkmbOISUhg1XMb190yLvJUxiDLP7vR4YzACpF1Y
wiOEV1vk+VZArs/j9/eoSk/43z4wBJhFaMVTZoRRWH+8l/EjJjJgN8z8E+TxC82l
7qOJREny/25b+AmyeqBFURhLk7aRleLvEEzugvENijrxtyN/pp3zZNIWheD6mfXC
ZIyZgARgXMVq4pOSdkihgVAJuu37WYQ1kY6lKZCMuLdNPbew5rhDDH5Tht5iU5TG
jpmLkc1idbGgwR/HFlb4dxdE6tKcZANOyy6/ZEAavr6xlsY1uDXMLbHmu5OFWk6v
IJMizbu3F72FHnZUP/WUnpE9GKRKzBPSYbqeie8iCUXA4HrpiVQvNQrR7p9kS6xR
xgpR3voZziA4LyOOr2OW59K4WIbrNFFhXsfo5/jeMNgpF9ZV+mCvEkLDAwhNTwwl
YqjYP6tRu+GLrj747RG46lmO2XAHBToyeqlH6VKg6GHQEq6yernrZP4SeiYcE6Rf
1SeanpFiCWJ8AD1kMQKMD3UIkWHDEWwXBnEvmbJe/y9RnHPOOrdwkAda9PK+xWWX
jG5lLWLRPvphfzMketFslaQXy9TG9TzfeB0h1Id6DcyF+xCbt4HyUtIyZ09lLT00
O0da3j93RCTyTgqSB2EgfrjmAlOva4VtpG3gnFNHoR02PL56g1tzg9aNirGm0rc4
BapftDc2b+NIWxI0G7mzdBXfwVbnm72sINU4d6INmJByZ2YOMzz8fjhuxqDJz0fG
5/0qdK22FHSwR5BUFdXAT69fjxbepjNxP6eUwXWH9pdiP1zP2rvfYBlRx/a7x96e
bl7l0PI1Q+XpezwY/u43PgJQgZSrl2sLaFSoop68eDZSRZcXfPqf2kzFuOr7q1/1
j2+XydYS34rV3R3tHfmcMtPTyGVxAHenY5V1k2Qecvc3Rw1+Pr8cYFmXLo6sUxRy
4seuqILNwHAWjsKJGnz1Vxuq7BngePBoqm59vl9UCRa3efETmiqug70W0igcvwgC
o0W8i52IV2UxQvpSpdCKkIHnPBJ4JjrjLbMm0PDZ+4/yshEBXe4J1veofmKA0GfM
ZY2aaiLzuyceaqPtCs3+tjltzRn/pex+Vqzxo2cB2h6Uhm/4CDE0pj0a8Gxihde8
eQVHaQ4/+WqZG9uY/lSKxqemIsII5ZuKGjjbwtR/I5t3CFpJRsml9YmaXkMPTILO
tdxL+Z6hUDGAGT1cvAlX09BZXahBw4vQl++u/SyMVMxZjFd6E1Oqw1tZiCBj7SIR
K83qELCyTH1C+Ag/e/W7wX38X5R5GXqn84J2G0U63Uy//a7u/qcgvgbzZVJORP8x
6C05cNZ2WeDiOxOn4ZDg4g8BczacEFtbcWrlpEXtzIlMlpGupU7mi2SB6PRTSwwV
iHysp5pHi+Fhm+16Kb9b1LTC1kLkr6JhdXBjL0pdPLPy4AmBailDUxkRVg/QBfgl
XQhcglwIj6YaTb4yib2IJR4YEZ9G+JAxSTvb6z3BdcOR/i9YHgISZmqwiRvwk5qS
PoKR7/TGYQ+DgaPMLw32ap09xPVig8ficZ//Gvr1Q7Eg9T8DQzIYR0b9dmpQBUY9
ZT8ydIf9ZzkmwcbRxOD5H5uuZEdGu95e0CTBQc6DudI=
`protect END_PROTECTED
