`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H6CHQuChUE0LczfyYXMQuzHT+h4RJYuB/pIf8vNx/NfVX9Q9cs+BgMZU+YlTNYmK
YU3LnX27Uz+L4op5HsgjGTzfijUURkGiXlDaC5GJPv4mMzchevDieIb8rdxwJb6/
yvTV6fjRg2XucDVbgkPcEnRBnYacuxOl5QXMvh9BD+DpawIb2cckUoCNpQwHv2eJ
a4p9cq8v8hO5+UEbr+waB8fFn2fvVvou4+R8sgEv+BhF0DJ/qKw8pX8E52C/cFEk
m02byJpdxLWR1wqLIrNDuKgKQcA3i+CTwZwCwyXYtgqJ3yWb1Sks1afGOyqzoACo
35Q69tsFtQ94zUZpKna0yIdfvc0PDBJAzg5fPiw17FAu5F2Iz8/x27xC5M1pJv+u
snJlUKVNp527aAgdI5gcbZ+mLixq6Zi2zgWFpImmAKA2sswim/riY3+mR+Lv98zv
EcqeR0naOIt6hEayb0u3M3EWmYUQbzy0q+8Lx+dvYEAhF1O/zmwK5FbUH0cML4y8
SiGrlgmwrvuVZ9cJrlRitvAZFlLha7Xnoh752EbBGCjMTKkS+iZV3XezTwIL3VzA
zMIlg4CuIoRL5XGRysoHMlkOe5CmyRaoNdPwMRNA84b8no2dVVExwmjn9oLNid2C
v7wVKQYAg56L49dLx29ikkQOpGaQa4HQ5q+v+0KI10y+o6dhDexeVk6mh0vgswMa
TMoNKbaO5JtLMxDzBBG09wst17u7R2dY3gbxa4+EsYM00EDCSznz2J8gA/w9gueI
zc9ZvPHYOJ96SmTuKG4KzmKogPB/WkNt7EehGkpC3Xj831ws7FVcxCmpMYdcaJsq
Uuu7B+FUuhqJTDSBju9O2nCeJC223fRssEcLymuaB/BwXoODyX/nLLy95BUwsmf8
kMroZzudLaQ/NeIZwsigRY3F/xVqbPOLyQ8trCUp1iRO3HE4OPd4WNhqoi3tW9kQ
t7JzzqX43SWQEdznWYDHmV7zD7W6EaxrXEGeVDLX2GHRWgnQtJqoMuNIfhIYRfnq
GCFquQa6RTSnlGVv0nVu5H+u3oSirbJBfv47vZlJZ+xc8GLNsd1irfoyseGhwa4Z
qCiT3ouVHG98BFJW47i38XU5R5ISoRzJwyN4MoWDHC6dBqYYeQMVMRRsrw6iWLN6
9E5seb3dbV/vj/NafwMmx7RL5eQbSpLtotWrD5tKnUbZPTgzGyMKNUgA02+FTTOx
1iy8kWTo/98zVL9BCy620gEN+JeQEf4cFZZgUBT2+24MV+9CVwrwn8PLR4Kcyl5C
9VZr4z9Na4d6/EU3kRowEFshwEH9k6dKzFIgAMWKY7t+9RB6rD1EJzSzHdbxl9zn
AOOljz3TXSMSVAK4UOYDtsFazJCiHUUX6Gbe9qO1OX66TnHKNgRuPNPJ79hI7f4a
SyP7Awy3H9F46lR0mBidTFVfhN1cuJLczY3XBf2ZaikUwAMrFhww0te6x1FHjXLF
KRK21EL0/rqMnFVMbUxX2qtXSpvL9SmSa/lS5HzrhDpZ+eUXozNsS5wTeTc70OOA
HRlV2Q6T8lzkE5Ru9Sqxt42QJj7UTsl2LmuaqxsTvfJa8I/YwZMC7ltHPd089zzb
wX+BqSS5RHk4nzU3AlxiUAQoMDpmhDMKj10sJqBAA0JIdV2eb4Qp+03MDyMLKL8b
/eyJGBrvDUAN0xObMpVActthZVN8Tq9Z5e5IzoJRs2ZS2KycA9e3lyfHLfLalpGY
P40P+hwJMSyAXrr+EEC5lsancEjFwS3HG1JdGpCGB/oCPPvEJxEp/E7nGY3nPUAX
4bzoNlodz7HD4JJ/Mal5JV1211V5I3gzEXp4LS1LHhijHGQmJCBSfwK7uWsx5tVD
/xk/HT6OBXT7T2K5jGAJGTz3v2K3eSNgR9iQwW0aKWQZnw1CRQ3ancPN07RXuNgg
Fe7uEZgdpsj3ira0LQpgriaB/IVRJwgVGvcarJIPieA57EEr3deVZMDZiSuP5FuN
Z788tmf31dNtWmNuyGrTZxhZWuCF3lTEj8UeuhBy5uTCW5ylB2W2xixkiYFlbdzr
LEs4Ev2RJhnPYQdsuHQaRLEckoN+xFbQscfSH3TpXtihki3JDtA9+kJ+XrBbhE7c
zJOQkGEXclJra94BCKfht8Gv8qsZqf5JOniqI3LOd42iPeIgwiL27fOwsmqhXX5x
QickA4JFklelEe23i7XunK5do6eso1o3r47anJuUucYI0Cpfbtq/xlLQ3GF7jgTv
tELkNVhHjwChNILyhDVHOcEKgB0sDaWXUtWOJnXla+Hx1qafua+tBwGUXQpbaFjE
RtauY0VhblZq6SiRbhTFz8YpH6EE15PhYI+9xfyRVcixGQsXBZnFZTLLb/rsM5JJ
9MKorsxDGsYdJFNXc3E3gGPkJ4/OcBrhczKak8vaI8AAbyJoSSgACDzb6Yw2ThbR
E63POK3e/bPIIpWxL47ElRMuaWyUnHvYCSQ6gVbeuXv4A4TfyPOB8kmUVpe5Evq9
tl0KVF9VX99Nm4a3D7OQzfylTFULlbKAXYwoIaHBQNABhCYBR6nfflBCN6CI1ZRS
5kacGyTeziR79HJBJ2trjfK2f7kpNZoKCxEA7YXbuIS+pQX1hRg5k4Sbu0MpZ5Hy
4ovwGTte0/QbmUgiYeEbWxiU2wIunFpRcwPgyFCs/3+C25AyHOSgplAVU04++T1R
M2Bb85plpvyQUAhm2jheYdwRvryQMty0QeS1Ud/X80D1PVUHhXC9AxZ5o+0KREvH
2oqTfbLGGEDZ0z6Q25WDz60e/ekxLRTTSwttOFhL5Vwgta1CLz+QeBaEKiw55YgR
+D7LSGXpXO7EPj3NEHxfSAEmzdcA3SLquHvzRqdC0rmQKjkiqfWRAYcJLvJg90LH
vpyeNCxTIJrA+UM8GyXoQAK8W9/RbUhCXpA0z8uDa8dYguLTF1pjS86D16ZZeqqt
PvR1jlgKv6zcIGxAf1MVFB3Oc+XqhrZALqw3ddwucWmHsK2jlbbJsoquy1lwujEC
KLn4A1Zic4woPNFSbvgO4PI+o5qA7wdUGygX3mHzh68qpg7PGs0MfFX7CwBhrImh
5OpgFA7NZ/1tOOM9nxAEohCrY9bEotMdFsxksIIKdar6bL7lYxPaP4S5U+y2ewCj
299eYUhm9Awmpbx3enWlYpuZ8RPPgiyaDfkhQ1oTjrHTSN4TGvQaMmqBFmiffTwm
yaZ+4PPW8YK9AKKsTzQFN9e8RaVS4MK7wkVguSd33+kr5Vfo+cAI+77CRNYramxH
1Yk5Ov8JyAuvrKkGLJtAcB13VaQkb/JB1n/ln4sv10qGIr5XMPVVRUCaVevhWsqq
c9lGhr6LmWnzMBPuY4k0hlQPkeOYGBUhzO42TDPgxyIPiLCaR3t1Ct0SiB2ADEgA
oSdiKoE9Phf5/+kweDvRyws5ElYuVXkWKQIL/rCOCBRE9wii+Wmg+L4CFIoGf3rX
+Ls4RBd3ohYLmBF0jqgSfEU37YpfyYhb27mdij7l8ZknZg5VHzeLECY/20nXwRvc
XrpO+DU3JVBm6gNY7FQ09aocwRyFC2vxbAZDdmRoYGZjJF4UxEj6KSRAQHqq5ejs
jx/xnpiXDqqVKElcnzLMsQPwUd4N1cT3XVo9j4p4L2ZEDmKul/t3XLyChgP+X1qS
PW8aMRfuq01qlSuAEPoljaUvA7pJsp+cFboy2wj5x8lsDs+uWF0IkHaO3IkwKgrL
EEQZjjLISEWqTwpxTBUrVzIfh8MFBrLsnOzK+Vkd1HvaglQ9ZkZshwX/c0xhUh5T
Eg2cOP19VJZcH+bVTJ1WALUd3kZFHNepxI/PCf9/vZYh5ePgLsyUFovmJYmmjaoF
e8hGuWD3zU6epznv92MR2nbpAORR9lmaO5rr3NjlxZB1vt5G6/C2S/YeCtBteMNC
wIC6/OrJeX6mrKJcNg+wrB+Va3+R9p0camzJ5l/3WIwCXrBVHBgcJUTtj27r8oy/
AJl4aQ4hWwvjkK1XSlsGjPIiMEHHCQjG2x0/Q/O3U3QZp9m1+PzXBqhREw7aZceQ
gffNe0WmYCzT3p5aq+BTGJvp/A49N6scVDDE+rbT8j5a/TI/eqJhfZQWYx1NzPan
4w9b0ajlTeIqdEIjloy5kBdMTvSmuXzMD5IPPU3AyLznj5IuQi/OEx1AbII7gg0a
TUEBS25m6FNsrUuo+bekYBfZBlm8KfzU69U6ZFI+TWDdN5rIMyS5OP+ZUvoOdc3K
f6rss5/iWo2Kvk7/gPFrhtj2Bf0g/LAD6PoFJsFzjkx1ODVuY5OsGQsJ2m2DFDDW
PwN7KdYkVDQnCzcIuWzZwATso7PDxTlTMmVvXnyJFuqzlGYk6aCl9Iisojc3IQQi
JXaeXjKL1bU4ZkqXr10fMHZYn/VUeaAmZMeHSJklYNhDl3RGEwSLEq7+XfOZLIMf
tzgXn3Nn3zSQxdrgKCBrj0X+e9160DEe0tKVEB/7mHn8kQhIMuHrZ07uUPw8vgmN
kdmyVnemWx6qYt2UV6wdI12GTEY0TvcSMmofXNqeFGtwNXdQAeItNyxXsQH/H4q9
2JSI+XhgwP2+5Di/8ZmV+DzOZ4VAssx9SpdK/qZd6MVaNc8WjYjJaKBXcGyviEPd
9xMatO19NxzuYFoGz5PzcAGKwTPD0Rqm5l9EFpaE0OYRebv7NO2LNpR3PQY6iRM8
zCDyD13h+8gMqHvkoxSHDI39vFIwvHxUI3yYqJANdM5rQ/11qZFgCW8IW1M7e0kB
TNYcnjStvWUWgWGNsDTf1xv1FK+TkU87HFQXXgR6KXRYZX0uZzA6u9rpAEwNoDiR
DiTYW4F8zjdJ+cOK9WloyYZVdsIq40rEF76ZN7tRu9G3hI14jZv0c7RvMav4XJib
hF4XdG1DP0Lfg1Cj5MGD12znCNpHKgzxHyJsAaO05BJ4UMkX6a+3IxSTQIGspX1L
PRsF09K8I/3errTHyHd7fX0B5+cL7wzi/QDIl/cUZ2JvPoBtyDFfkiS6bSMjxMH/
r54ZravUNFtFtt3UySiaa4OVY+BVYF1S5DgWPT1q0TdwSrIS2d82ru3tnoS4e6Rj
zCswDopNEXzGqlQWpLo/Lpg3Uv2C39twK92MPCvKtbBVjwHQt8KrqqELob2mfiIo
I5e7MipNPH53dbav/16WbJvuhs+ckGTSFocrXd95FrbOnx8Tp2x8a5fXYIllVTHe
3yhu5dn6AC2kLZkGpFA5KAVgWoEzJI4cWIZ6BgUsm/E3vBMrnQiRPkaJ0j+YFMkE
HIdsurr7ytZV0cB8j0qv76AdNCX7ClRre+g3dWjtMLi8/ciC3Z3JthhM3HwhZlXJ
/iMk5DZKaJUmShynMizAtnSzFHX/cRWhvl3zrRgiQPN+/02y/V4ONDAMLDY3gwu3
GxuKWDfKw08o+6b66eb/M/mHOnSwTNrPg1wCQrcm8kDwfHRIoNz0mwn6BGTURmbM
2PJah/Xt1pepn1+NmBuo9fwaa12I3VwXaTw4qhhn04SOJwzH5ys6k20FXyLYQNnI
eibdv6ia59L+gFdX906gzYv1aP6skFnJjo954oPW/vYE51vvIhPPTG+eLFd0cvc2
FAOWGcM2kepTnuCQJe5OzWE6V63Xt5it3xvOEGIaWdLH7vxMKdPpX3mkmNSS8wyr
pcR7JVzO8MD37+TRZkVgLSBDNc6mL/KgY9DBQ+0yfuem4xBxOcW7rLulHFbJjVk6
MSg2JIQe+5lZZggwVY8jOjp0DLZn17pbmk9zdMO5+GE4woN0Okjo+nCOq+fzjjt0
GeWGu5R+V6T74/SLekYDRjaGhvc7Rw1jbYRf5XMzTsoed6pIrFWK3BntB/DW3ypF
9FTqjeocVfHLIb2LKSlnOHwTRT+qS6SzGvm/VHvceBcNJsG5x0kyjEye27TsUylY
Jwsj+7HxmfefJfSp5StetlyKcqFzeSwZxJjj5WTJbNL+yzvCLGVFTfqYzu2Q5afS
CTpcJsrghvlT9PFBMX9R/WwECATYdL8ZvmJjBWU1ZksOGGCeeUWUy5dhBQJj09xK
AmYvpTHpa59yYvnyFYjD7BnK4c31KD4UzE0q4cTvrVFt6jheoJ/m4yVuxUVwvjTL
2bcpEKovLIed0BiE274TAWZi58E8pAMgspTjUfT3Q/QQYm/MDihHSlNeByOkcN3z
HJPlteQCYW6EI+R9dXsay/DKEAYD8/2ZnnMMJFRDkamhOskHga9KceLG8/T6CBFo
NOeOXD9NrQ2+/kalaBaGzUsBqU2Sk4rmJzQUqnBSD6Ydawhkz+bwvNoRBwdkY7Q6
JLqu0w3Xhr4Z7l/ycDOsJJ3zN3EnVv7yYWipKlWXpnqfRW9iysgpyV89qht136vW
WyHy3uBgXoRz873z32w0uY9G4e9ayCkZRYJbbz0FV+uE4nmL3mrqJBSwl75R9pyn
G7vc6Mw7d0gMksim/FrQbnp1RHRY0RmkGopMxM/0zBnNPKesR4Cq7R8cLMgRze0Z
Tav8l8B7kU3nl6covPO/LmW7zUrynC2Fkh/s1k+8CzneSLh8rh/u8z5nAaODeLBI
PQxrMR9AZZekL5TtmsSOq//gAMjdD0spQ8+X6ILVzxrQ7yt5sazh3kZhGZ4xn6Yl
L7Dlc4pwuqB+ukXZfTu83TfPanklx/EOkkwTFYddnlTVedLetueEgbQMCOKBOPHM
SSWWuHj9HM6utx7uYtvP+N7epBgjwe1NN8qDIM8o8uy/mvH+iJZ9wov0nZxbz0uZ
0R30nPXiPH6wT/8F8qDXzjkNri5fHkXKkxgjMsxFrOk8UfiZPhQON4J5nlia/8Js
qvvGlNCm+5Xmx6trciOsBwuAEdkomb21bMF1xBDjWkVJ1gdUvdjGupTMb47VfgK+
fNkU8p/qn9BwNPBrcfnCInPXhaxxbhLIN6XukicQJ80cWSdS5XUrgNWD3U0Q5ALD
dP1ZGrfI5HdPKRhAEZ3S+3bz0aYQFehD/5+FIi5DO6p8xpmlqfxRpqgxgiu9zZRF
u+cWJbfYdu8Pay7zwV5WzmovxJuBacg1CGgOykgE+KG/EcQzNJbilTETYQpFpr1E
+SXZ79jTdT9DptpIMjfc8cZVt398oTYYWa2NueWjqFJGR3gce7zHIHMJ1/V6CVsz
9XaXr3BylnAVCWHiBkDvpgdgLi/fakgNUG+T/KLXXm/HI/W+gsSuXkZoLzElNwYq
miWOL2fOq6/FWsrI+C8ttpFc5G9TGqmG5WDk8AuUsp1/V+wK2B5wWDYGAJODt3Zl
L4qS1VeWkk5wy8mQUcd5xtLCsGPCnoPi5qzI9U8YcdeK0n6j8O5869eneP/PyHj4
nJeYOVGq4AEeCiRuR634NHZa8ppgYZJPBg8sx5re95ba7QQ6mPNf2SiLeRX/Sotu
HI7oJc3xdsbZeMKhbM0hXA==
`protect END_PROTECTED
