`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fNhPdffsv405tdYUoeF1wXG8MLEhAtw14IDG1nYwVLu+5V3rUgMBYPsV29hyBIEi
7I1fR6kAApCtDB2kk5PfsMz+A4OkfZzU30+y95L6dA+uYO93lVN+bMyepSLZ75aV
WPuZox3PLv1+toqTlJqjeZP3WcSsZPfdwaA7GDe0VDnUaFrw+NLWmpCYADnL23L6
u8UzkbGDRp2LjbFR5aRGq7wPICgwx4JsdVPazX6zU9HVSmz/jfK3y5dvZV1L4mPy
ABhzgfvxzB3ZT8OgrVTcU0nxNN+pw4ZJKF0RRMlTUFzBVqwSIOf1eGI08Ekdxzy+
AUNx7hUmPn7C5oWPFTC0XS/UeBY2fXvgRZCCdqINx0P34mPKMbeBSPkWLQt2wUU/
cEVwmF9r6R1cw4dqk8HlVCVongKy7ObbHvs30s9skFwlHF5aI/K5naGQYY3GJGI8
kckHSFOIijoJXyiJZCOjbggj6WJWd8loIZGCojiuT3Ehgo8otSFEh/f+ByRTVr81
ugE3d7Fr5Y1//S8Oj6HcEGMUGZsq4bpe2RlmifY8ygY=
`protect END_PROTECTED
