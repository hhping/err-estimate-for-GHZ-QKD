`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v6X+IMuVEyr6G6sbxUeiO/N0Kqls9Gd8NXiljh36Uz0CyI8/EBz2UToWEbW8v6vu
T+T2FD19zM3tXas3Bt3dg2a9o3NSwTrOVozacec35xq//xPjAm1BeBzcQjC2sw27
4tGpyrNgImAUNGL5EhvO1LD5VXRP5Z2Ciaia/THBfcm8zwHIQwiB9vYdrf9zb+1W
961BNyktSkK7p41wfnFuvulC5ty+rAxgezYVPbKKGDIpMP5hBte7QgMROKrY0enb
buc8TAJx7QaXMIEsayeeXV12hvFwCJSSrkfVapg4dlIX/BXkkyfacxHZjKD/FOs7
WXT7H4Qani8ulwf62D0qHHxjyHJZEc/TYF1lqaNWO5EMlJ1FFRQEImuVpZ/Pu44w
hYIuOLbsf8t1gJ6tcnKBWez6hMbRpmPSMTPg7OfY+xLDoS4N+qfYRO/MDKwJRVRA
daTRN1PaQKozFHMZ6AQ2T76l0pgstiJTnPfCCfp1xhAnozqxb054gmRcWL5hVIjd
zPZSsur2rvNNKMl9XcjzHm+lawcw6qtPylMpyteiYo/5iLKCCO7URPtzoxlcZnKg
ontar3yokfmt9X8E4NHgkgr0FtuQgGfH3mNcdDpsFw0e/EHFpeGXL/fjsOrj/1Re
CGAfnVOF136FOqRNeCFxURv4rVahPuUS4a8jDDchL8aUGa3ftsBLe71t8rfNJ2rI
74L3dUfMwHSi2r1S1UmO2MCzRyRxje2zaS+5Ae4oV2IuNwXKE/3INKaZFNfOV+AZ
`protect END_PROTECTED
