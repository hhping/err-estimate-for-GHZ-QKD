`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6zuR/z1Ic1G39S723bwJvlTnnPAV1BuYP+S70CIoR7M/upo3bTnBr9KW3KfIa8+U
sjSzyj2MQYS92RerM6RFfn0R0Pan8J2aMPlwLOQlv8T2etjrRXTjqvk66U/96u0s
aXVDbAyREEz/z/K0i5Vc9ZMDgeIjJyjJWzG9ywOspBb0YC44+4jd9x2mPZh1IJXq
tg8SSSnESXzbCa7rvRkAzDhSovaWhqUNSU9AJ+m6w4B779T0tWDd6zJYWuYwDxY7
A2kflBGSyca6nVbV/LE/u30g+aO9VAiTH6+DsyhgAIwyJD6QKZqrroGqRYsORooR
vG8hMmcGvz1uBDTfT2kI1Sz1ahtGVFw8xMekFlNH3QB1DR6DJlgZBMh4VTc460QS
lTiQX8JhYBQvX4lZF9STrivEAYoXwSix8LpVzaUT5vhOpNyxFgKGBz5RUtRzpsl3
xsmEWUy7an7MuEnRT9yYvtZk72ulUMq4eoMpRDWVqbvEAtziD7livbJvgFy49k9J
kjI+eAVwrNSnkePGpUW1DugPQSRXGKY9FrCA1lW6GTiL2baZHE7qdEKIBARjZL75
ScWClMHWWP7vuC810sGVH9rZXAgETuGu/lIehOcsxxyDsOfPdhdFeboo3l71jqYv
7lzS7kp6jw3rEoRa6B8gPUurt1YMEs/hNvlllSUSf6x8Wr6yz67VDunluh43cukR
HiaBIkCcQOID1DS3E0q3TvMowPM17kQZlq32duj7GcOl8nuJA53DliGxc90Grqte
HRpeBJIEGDZOMrCIYt9Q/j3e6jgI6Q6E9i306+crfTP1PhZtOpiODr0FpUA/sxzl
Y7qtvPdsDEgizcpwk42wfmQ6lLEJSK+QabpRaJ7ZPXbUWL4nbNa29cmpGGsDwKnm
cLU4OeAO/KaRZS6keFJ70XIVqAz6++GR0S7QVvIP6CjFukbRz11sWB1eiEoU6He7
E2aYuoGwJ6A01uknHEi/0AZzFESXG9lUutv2CfCT7IM3BL5LMMP3JoJY3iYdBtaX
D24V+C2NDsvzQuDShEgQ9RRky3ldu0UN5NPNkThLKtJeHwBieNMK0AhRToWJ+jEi
hBP2WyRqDhbfKjW/QNJmHBjWBVTgngLDbkmJBzwgyiXN+sdQ+BOPMEj1/81G9Fdq
SwAJormhINcl04KLI79nsrmxNnuSbGGDTWqzJMKX7fcZyZXS6+umpyolQtJpWWxU
H4Y86KSA0xOEuvYplArROq2jixspzG+YIxyBwD9Pj3v+TeCTpe9ntcc7WG2BdxF6
`protect END_PROTECTED
