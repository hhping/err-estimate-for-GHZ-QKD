`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tGB3sUsS8T/ABrgxvCbkdILISIIn19qKT87ccCYkPBBy8rzNiiqy45ZgMn6UMxxX
jHILeLteAUrkCMzvhaK+38XW5ycXV0wRPC0qJll0SfIwxhbh5BiWUVSUqdUn8WDi
w5Pw8r/7UplRNKqKvbPa7dX5xmbtWfZEY/PdLLKX5gfaxaEkHnLkklCCs/CfRmZD
F4KVRLY7TpQY3hxWukPm7E1408WPNvpWBsth+MM7ut6iw9MXBU4QIVnBD+Beuhm4
QnN+t6D6EBCPbq4RTriAya43DT3sK8a0g5lYBgip2goilNBrliq6/qAK2ZrAbXVn
eWY+sqkJj6Ugp7yhIm/UkaVfCG3+W93/SW7SCkCZVBUrJJz20O2NCiKVKdUZ9Lvy
hk6oHGF/ja8YYwiZ3T2b7UEHEdJangZpqz6GWAIFYvmhmOIPrwpK15P2WFtXOdHb
5Hd8AK/yUCD9mV/iaBHASagSGfnmXPOMOmbswHpVysa1wY6HCnSNsy4m5pY83wCy
FAjmPLqVQniVQ2pnAmC2ReEjZdL4Qj23rsrQ1jUus0cOPPDK7GxwapRmdJZOYKAU
MI735TCszi9xBb1/gDSYLj2kqJw6eVSvip3JCZ69gEERVh6MDZ8lrJE2dJnBvYgG
LCe/q7IZnbeic/F06Vfr2eNqMunJ9D6xz+EHfM1BYLe4EDP4AZxw1178+yXZSZDJ
DStH5T4omXeKaUgSnrpKuaVRsceA+/E6mzlP5J+4c7hE0o2TTUGPogs640pxGYG0
vf4OD2tWRMl5pK4L3JnU9VEsBaaJ35KtSG9l8PPY+ZW3kw2IfEqrMvy+i6tRjaTU
9VmlmUbkF5sAPH9vPg39bpcYL2fApN7vc8IpDMNXmgCBFsS3whOSbnmPRDzSSm0f
Ac5pUOVpd8Yoq20o7aYolKTdL7cBRXc5nz3ZvIxaoSqRfTt6/CRdu7orY5H4d86N
A3dARXOMnuyxNvEVm5lux08K2B77YIZz3S53r0KTCYij/nbXzRoaRTiFQ12/Xx/A
EpzH8y8jOjN4KNWWW3TzeA==
`protect END_PROTECTED
