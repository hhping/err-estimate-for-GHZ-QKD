`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/8Ld5WTJki3KyLBTjwlzNNv+lxktWB07eq97GdhMAk/xCrKrY2LelcgF793jqTsL
6Te6k+Y/oT+9PNBh/Am1r9T2gyGMWYg4VQ9zZ/ZjP/MaGYM9PBx4Tn3UGUQ2DoM9
jUbX8/mWDMylsz5zi0hSQRu3Vx16D3W87rAsHT/bPQuutMhQ9r3kXUjFJ0KBztrC
nhswvp7qMCTYibTPTZX95YaEwjBaLZrLbrKsQBoAVb59ub37YbytRPYS2PLPSDfq
Cgf0yqklz7SS1ueNkFDodcE01kSTZx30ulYVTTcYZO1GJwULTTxyyOlCAAJ7POd0
TnRIN0kciVBqxsqqmLBOGtn5wO4Y7dtUhweufcU/70spSTQxDMiXPVfm7wiJjpQb
b1LO8WJwuf7n7ZT+Q/XFNgteVGdn0guLNn56oPwHdtR0T7r9+AHfvGkx6ujUGv9C
iwC7vR2ncO4i8A0u+N/KDSVpGcok77UaKN09Ly4169dkoytTpQTy2gXM6i/PW+QD
21ZeQfolojG2ZvDRiNE5hu2wtrxxNz4SNth4nPUviXVdyqdqcu7qkCUp4o57MXlX
MyUKmfhXli40soq9zcjgErBROfblPOwJ0cWxWSFBx/fMxiqmCE1sUu5PLgAQMIG3
4FkcMav7nUV9JtBTC6N+Rx6u1cCjr3KwXbAU4/jM6CKiZn4j3Q8nQnYzIKIfp+Ws
Ct4MNYuAitkTHhx+/nLXAfgq+yKmN2I1hyg3kEN9n7Kxzxq/THwanouVJR/pmNJ8
g9Twh0qQ3W4g77OTrSB7Z32XIBLBBAvRuAL0/qp8KlDqKbaTNSojiCP0sJJOGvBT
ZzeC75lCvu5GeB/Ki4AB0j5jI3XaNEy6HFmBY7Ss5c2EH2PFPTywVXqo5yRaBk6B
fDbFsuO+OPAareeMKXPCFyWLuWOcmwe5ZyhXYS5qxAPeCKVNtdZGE0zKNIypyknM
T9RNPx5oP/eraaHTcWI0HVxzdz1KffUpNoM1IRh0NNqVQDNmEzCGafebJITwJh+S
BEBUhpWSIDNHkAhy4BIa3Bm02HZ2pe+QY2a+8AjQ3IR0y5IAjmbZHPqldIUZ1xQz
ZPQSc8jK3QFnuYuUSkJk9rW/PiJPmoeIGb9z2fn7pxs1QsmUv3RAsgnkUxVATWo0
24kiCx10XcBVskVlVvAWqsAk3+yKsZ/RQtsgm7iOnEIuBFVPYnOKQPDOdIp/zeyk
b87FbqemePiA59dgp4CuZ6qq4eWVHm8ltzjKGfZVaOt4CyDxklzwiJWpVsVDb0H7
jREsWx94dPK0AnY3+/q8EUwNEb8FMfMV/GsOZ4goSJHHbhX4bPkTDVWg3y7CrfeB
x2VYfYlDVzuwDAaPXnSzXpzwTrAijuGlIb8BZccptihBDqrnY/JxK9R3592x7KOM
eOMC2gXFvD/Gs54XsTrG3WdpmY/s/zNCS0ZLu3DjBDunBCWNlySWPgVd/g/9zy2i
gB3+TVdHahSPDunutHZoDGGG0+gXTLl1z5Ojum7PdVmliIEQUJG5Ccu/Fn5E4sJX
kOkwevQ50xf3BJmJSyOo9eD/slEUta9uzHagdS0TRvLaFhmCzXKlgmqJefPxOQp1
DN3S+wODbzMERWjCuJS85cseMn4BUI8L97JRjChcvAnLvHY4SoxRNII7kmTU8HJc
sTVcQmk3m8iVL5oXf1bpSAkxIUr2lroiBPhItOeIJuSwJ4HNs8G5sWSf48VMLm/W
9V5+Si7JXR8SGl5P3XEQ/Wz6OvgQjaWyoASgNcvl82+7f6+uqvfeRU0J9BUq2fXt
9ksOarCzncGfrG9dr61cHiml2Xn0nEvrg50DjtZeONaFgmmg+yGhGeNbh3vuje5+
nm8tB9euUFBwKGqyjbANjfg728knbsPxtl7qaGI1mM3Sy6YV08MZqvyAxw7pHAPJ
N1skaq7KwwFh/2Kwgp+AMM4WhaaOXgnVmdIjk8zc4nT1/BnMZfAV8nwb20fRAQvW
HXjG8k5qu7fyjm7AirkwLjtNAgG5dI59mX4WtGUPkj23UUkuTl5IsAPXZhuiDYp/
bE8lFcnz4vZQ/P61+2bVHIfjis4fDI8RScU7zJ99tPkXLb9aasT8HLUbY4oCZbFG
YzGZC9QrZMvWbLubx4SkVfB9CDE0vOtjmVI1P19TtLMfV7fTcIVuszfPfawKsEWq
/A2notxz+kW6vfLISyzDfiUsvzkrSi1WrCVAi2sw8X0boE7VNA4TuaVZXqu5yA+l
U620FrQ/3d2jWCrO48Q7Wi119EbwHrBYMcoyfq4ZuyEYz3LU/G/Hp6JQaCeRqqfv
8bSMl9zv0r7YVrWApmUfdEsOYVTbKuAkXKlDUZlisvqoHiU1kYc9u5yB8icVQqcu
ymdomL9zfnR1rshVm9bEuxMqFQDkSmBQSHMFksBXypwaamf6RGtw7sSuhIpX66Op
ewmkp044bB6emX7L0LB0+8YnnPD7cYYvpvKxJVuZYd76U3dIPXaugbxQvqHJXrxG
XbdmKKpsLvG1z3KuuHDNvBQuoftJOKYSoUzi2xvI5DCWbdyD7jH1+ol/Y+dvfFs+
8K+acGAhOhPoAYEXOJtTrW56/bB6zsKKfgu5Nepp1JZA++YLo7X2cY6VWg4IYDLa
YYMKhSLSiQ53DlhKkGGquEgWpam/69VmoUL0xa98NOSjPhSPGTj42XDJW1d0cOsN
fgtluKgndp0bpGx2M/RTvTZH91WZ57AsHoGL2PwoXE+SMod/ky+ml5DvsfnQTmDn
GDj0aqRIRtZ34DDp8U6be0VpGxn5WP5O/cAWhiQw6yFRK2CkCKSW7lx/8ianuqfk
kxu/y8oMmoZ/R+JiPE847HcUB2ZsO0yVsAPSUQYioRv65AjrrzCx2qk7saBUE/zG
wmp/mllsUaDfv3APh3y7gdrPI/OqMesHzSgpKEm4rnvTroHojvv3rlwfVKFnpd6E
LovfAhUKbM1LumnWWtsz3HXt7L+knb5T6z7sH4iOKYEndPFIb2dJe58Dx30MRiPz
lh2yKX45b7da0ujYxVCH9O9bxXUzYba6yKTHaZ3K0d4pyvi/abtBLFgA2h58yhk/
Kp/+ztjAOSooUVjWJb6UBF6K+VfyVxnrIOZD9xM0Hc3DSIj1t97vCVFvuh8zt/3W
`protect END_PROTECTED
