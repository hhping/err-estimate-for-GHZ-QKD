`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tP9pjDWW9edsIeifY9sMSfctwoL3NOUtyoDyzN3VKbzlHvVcBGFYoQ5oJo/GXJev
q0o9wRgFFrdx/myT70POO56f9ZPb9scvQs/WVdIx4uQKGE00Kr9MrBjxgOK2MORu
xvCqcUPGEOEeizhG0PI//AGoV3tmlwklAwpJXWENFGrhNWLAt/D9+10m/gRHahb2
ZkC3lNUsbYLastGXy65Jo8+isAdbVvdRUBrBfu3XN6oFhIwAfxO9tBqP+ZrHWUCj
pjxIaQ62MgXpUFGuezZTb0v/+UyazMzrmiOHMPfn/KbTlYIQKTMv4hxNW84dpPaz
NcnV/ts+YTuMN4S6XJQfNnr9QGijNY4Kwh+OyaiqYVU6B1s8xne1t7XPfbiarDMm
YUndfkAXsKi79g0fVzTWb7TW2Mgjv7phZWnl66ELEdIrYOPQVvIhtj0qwTE8L2Oi
f1sa5VMV2537u13JbpKUSaZENRwIlOKUp0TJP1MleBiaxnDdgpfVVqG0ZCfrfsrz
gl+xDo/ehHXHqGH99LmZcUk0XYjPCSzLeYsuIbkmeNx082VP0JvMRmkMy04+iIP/
dgarOkFoGZO7s3dwELoprBrg5tYinB/MKLCoEQRTdu7T5aFpoeGsAWQPOl3IFKZD
Q41KStq5ejueXgGG7+IGY24LEIqnzO0ok9f18rMPe8d4L9mg6dkWwkJYAO9XjcOi
aAYUAmQgvRNYiniy46W05dhP8xPnIlTExs9EEQ3I9dBYaj6yx/HwGAYSdUnv3PQx
8CnbIwdobWT2dNI/YcqYFwRqU1yK/IVlRdUob5b6VsBCOj5Ph6DyeBTs+WgL6tTf
QqLWSGkT7Fm1g6IvwyQN80f7rPa28qpMXIaJQvYn0UISNco0tJTHT/zS4EP5WSYo
SFPtY3Gzcm0yZuu9FSd0VWNi3ouWq0Yxioqxt+JlMd3Pqm2NmwnIcHHukb96ygG2
KXtMwzk1fv4tjH46Bk49OtJJqesGBqeAfSaQGROYiObzvrkjGRKClrGSp45l5G29
il0YwXpJN9G9gpLoRL5XI2ppxwzhu/vQdFEpr0SbDd/P/IMVZ3VOc0wATHPXTFt4
7LpZUwQmKIIuZRelK5l1ZM/5CHQUCaBJeItgKhz5O8Oaf+8/6OAy6sGDE0aG1W40
unqYUXx5pr8YZmRpFT3Tvvb+2px6DCWRDYbtulU73YwbnNGEzvsOE21pNsIZHSeJ
uMtlw0505irR584RJpYkdT39tQpJ5P/6qqDPJCKpgM5pVBDf92N5Iv/JsH+rMgd8
UwTccROuGoJYBnIDmoKCxFd+FFhrb2RG5mlhyklyq/ISadBAZIxTgmWm8NZMMSRV
KvEaprcpFgAhk26Q9vXFwzs07OIFnMMxeeMSqj/RpR92RDb7k/dSW7k/kw7ndZSi
Jxnq38lYjiHH5G5TBLa4cJ6IsXLZMj/HGdhGdDQ86Fp7q9nb6nf+SpOSkhX5EKQR
afJhmBIWmaXiIiQpVrD8R59t2ZnyRjhvhXdkksLXRl4jroM9S1h5dsDQ1SmtOaU9
3MZlALAbYDP9JM8g6Wr0Dx95flAYfG3KpslVLKdVCxCIA8vdv4U366hpVSuNP+Mk
9q0esziPFZRw6QTA3hn9639AJ/gUi4iKUA+GgR7V4OjTr0U/Ybm4JTcKFG7slQeJ
IfdqDmUNSjkliWeG6f4d7UKHCkvgS0BHAVYhJxNd2SQkk7yhA5jSQ+xEAAKbTlmN
LCczUe/jKqCviPW+b4LhYItqGuCQd0di58/xBSdH+9wFUltAf37veqKCTUqHOYZq
ponSjTuBxHbpXGsQKC9W1o7D9EItlQ5BwS2hGkvkQt6O8bPoGfvI7DIUGPxoegV0
35CXOANd+54ZoUYQDyGcMcBTiVFTG/WEpAV0g/bs5o8sq9JhTh5o9n5qN7q8MXsZ
AcBrIGBAptgnkAcwU70XgAaYm4t4EeOmHGM0TzDYto8v87C3wsOA2NIstQ/3chWs
dF4iBz8zW4t+fjRZztMOziXsZ+9xJZNaeYmbmb0PxIHZZER/e25Mv2e8g1My9Rbn
FUxnAaaCkcvR6t57gOOPdDw6szEeX0ouD9wHMdBXX7W2d0hjZBhhMpjwbWRgomtl
rkl+O9KIK2c5nZ36AWLEeNVmz6gro3Msrhz4N/kdOm5wAqp6s7aaJC/YpiQHEEN1
73L6/T/fYbmuNbn3BJ+GpXPPnSxkewpU3ibvklIpnAfYDlma7blN52m1edDK1mX/
VGnvEYexm8hf6d3qmpE1S2go0fPuniQqkzovmmajdkWn4cTykeE3ny3nVUjPUWfh
1smanN+8BdGalVHyvcJo8xlil1J4Tc6s7UqZGoUYMkn1EKmt41n/RArOKG7+dZ1T
ShS5QZ3AlwcUtujAdBm5t3yaflT0/k50HrBIwBrdEelnFtjpTfw6WHXLRkCFWSpX
VtnUg0Y/qEY82gfa/+SAobFB3TR43QkCKNrtWh1iEBIydbq6r7LcZNpKa3WfuJtX
hn3JsdtLs39/rdYeRSY6tnqbxXojCi1BttGEvMItcZp0BPSSUIiFQJJ3meVwnBYy
GGOG/yKRzSz3X9lBfgo4CuJigdPQ4VITWWtQtoObpe7DeYp3PAq4JTq5pCiKw8Jo
p8pfgDG93FXHW5+ntZnZK3GdFX0eamSalSuP+SIjQiBNFJLwCP6maTTzQh49cONL
DY86WwwArb0QtdFxDNJ8eHWkKvA1huF86R5YG4sa1jhOs/tyUBkzQB/7VCG6fmCl
4EBlcKuBs4mVytTLq0ubfhmpRXwo9VFBWxTEWoySX+yoOTa9n0sZV5AdLIdo5gcD
KUIKDYrTvxW7qCEPwsVl/vHzp4X8luX0BBZMJQMdBcenrJ1Z9Y9Afd895XNk+F/D
W/qjLRZ6MhhCT/stq9pR0dJkOR/bdIu40v/pibDkRTQLk+iqDAf39yNDNmPN/cR6
gI49K56yTetnQI7EkEVj5iLHheEO9ZGk+PHbLwiUCsRgT0lXnrYnUdkfPUbdk5qv
h/+nT5QwprQ8AMESw02Fz4h5+71dWp83JCDsAFZrmpMPQNd1ddJA2leHlFpgeKAA
AjfpKKfx18N3jBDmVCXIJG7lQzlDT951GVliYblhNzehDbU8fydf6suvb/hIlgnz
Fupkkfd9Yv1WnSqHCqRw186HZXaZkJGYRYij3DcsWK6fu3TuOCQpgh6IRUD0FBUl
PqgSnknYvbUBcOQO5gu9t6vbI04dgIgLU0++GynkuSLjbBx9FzpuzfNjg7oaDpbP
uFwKLOUgYqB7fqm0Ehw4hWfB/9Gf4/3BAyW14vvaqpBZh7czM9Dtc8VEb/K0QgXu
QMz6FYdUoxZtvTd0jrQtfQJAvjoWyT4Fkz0qo1dClOmejjdLTu+wd+LPpSwwE0Dd
GOW1uS7ULq4MXZ1L9nLV+/qEglJGrVx9d0Qm5O0KKW8nOo6GUKuH3JSaH9vyKlg0
wFvz+Svgvp9XxpcoYJg4mWF4CvBywfD6255xUk+SlZ13wuebjJBvGP0U9Nlz4WnD
cGCjei+QU9fXqoIVXYSboHkS8Adsp8ouql3KmH6NJu3q1AIhpL3rVRvqYebyN9Rj
Wkqk+lBPxtZ4IPHYiNrU/fD1CFLHXSQJ9+Fvdr2Re3+QjvlxhN7MZFbrCdFeMoRY
SxSSdiIQHVDycB7M11mzWGLfkTxJkrm689+lbRNIEDmGTlpZVN33mpQA4eslBJ3Z
+RskyigI61VRw3NUarkhmBY0Z959ZMhzmUee1/Qiy2KlNCNobAByCrJRzJtrn2h1
cxEAFHOIxNcNrqw0uuw78A==
`protect END_PROTECTED
