`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xibvDNSpLe8cFKvJMAXUBmWijkfLdoz/GiFOTk7Y1nM19uy1mqS6VmdmhqTUm44W
N9zp6hN48RkRHEeVgndtrvr2YCKToF8TvJm5EkCaAgibA6qggqsXb57omROIUeLd
pJEZrb74HtXznWnOuxtMMA7FmKxytZI9pm9GRBLwUijDNhY6ieVMQcFfs0NVPqlD
gopJMej1KdP39G8TFbDH77Pq6Md+sAdEGJhLFvL+CixTF8j2BAStlqUmzatk337B
GzXNI0JNUGI4R8GfHP+zI3TJXRUstWs9JGZR64MegInLh4qbPeSTOxbpuZrwGpWK
qpWe8wqvPSBIcC9/yHEXh4wGTNL5yx6V1jMERJaQem0ID3cLk4YQAIDa5OmnJYzs
MMMRQWDtU4JvIstnO2NR83OLkBmUh/zM2dfvO/cqyvxYUBHsNPVtOgu/5JZKqXGO
Ji/kJXl6rGTaxNY5jr3NWxh/ns340IJPU1Hyk+vHxFY/kFEiZPKp4kljoHKc/VaY
HBjv57k7VI0ZTUO/TUpFOS6Y4Qm+HrNbB6AoorAxbJjHNGPCdDgYTcajFDefKh0n
HM9qv/X3jxrvvLnrOV4hASKpEn9m1aUTDI/YaQo493KuDD/Syg4ozMwSEyMMQ+CQ
ZfBWZatXd7U2q4o0IgU3K3wz4wmawrJdP1TNJnsrjoy3tsliyd0Y0glNruJdQypH
IfwTfn9bPCzR8f/5DiK2bLiTw3ctpPPXoVLDcMIs5FyMON+ue4GpsBwZoxLbVDs/
QElOWRAxtKEx9uqYQLDQigHwL5dyBLFhyZIXPYn+Dm++0CVHyQoC369b31wqGdJX
Is1WW+ZQkZOOflDqk0G99FXYbj0t0ClnPE5ExTtnXjGalcaNrCNuMTybO3z7tHgM
IamiScwiXJl3nCrXWnR8d/lbWABpyt9gcCwKEgl7mpwvXzbpDVROJKmd0Onmcqmu
aTB0NTE7naRtGt//EYwKkcmznOWGDZpel61ZJoFJeuJAIkj2AcfsMYUfuJASgoWS
VubS7STYOGo298XnTrN9XSbAy/s2Edut4EMt9k/Vult3LoWXFH+A2Y/EjfvFJZHq
jN1GBaVwvIjQ7O2J9c2HtebA0YiiZfuuJGNA7tDjBNb/6DGntj31vmCFlix2eSKR
9pnXcSpWdaaU735or0aQuArlvkowQ+Pi20Psgy1eJp032rVKOdr19pv/+ZweGUvx
HfoywbGzwJ1zxP6N223DvxmwipfGDcRtkPp5fpu1HFw/CRDL6OD2Kq1g+VJ7qGs7
Xj7MpACKuVZVk+UZJLyMyj9bnML6w95K6x9rF78G7zmg38J+jzfs7EQzSffWwd8D
mlBsxmD4vWff0uCyXjBe9uAaGEOZOvR2uXRtsMK5P5NkGqgFtfnxbodrIyAX6OuW
tyQT18ssMAkbT4JswSXoCbRuiYsjczU+ytLscqiSznblbVf7x8ojsI86NhRmck9g
gkhYMVtcBW9EHHyAeY1mdRUhB2eQaYDHhV1D/pRj7+AFhU9xstJAtkU3ez6JunDv
7nhlaicgmaqqu6+pN5nfkFtUNrgXEMqLEfUhqwtN0+0T846wBwT3jj64oXJkUeXq
Pt16jceNBSBNgL4OGSb/L1B/EDx1OnpVFEvsetNJBEOTIHzKJDnle4INxFTawsPf
EE0YwjiWjBkk/8Are4lFKA==
`protect END_PROTECTED
