`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h8dcJBVHb9p5a5a5oP38sBnEGejPw8U69PA40ej+88HDZySK8F+Qzq8sWYV0ikKF
6s7Kk0MRD9tVlIENJMd260ziCNpn+CSoyqJ0PNabPqcK5uq6caYSe652Wv/Dnno3
9Y/rvhwFYyGDxWB2ccMxyXnf/NnyEPHse9hOFrluYaXGhxoqJavDhwtO+ZFLqacx
uznp7zng1Mn/4pwkdSzirV3exkPtalHhF5wMmyGbPQH91OC99EpEIWXAoW2IWt3j
joZ2kuWz3OFM9SsgK3ONPoVspfkaM+7BMLBB0cqH7gSylvkbn9cUDiSbnKAPbVLd
KQtzgkVCw1VTjT0zpFhRmzJekkeSoKSwpM/Y24kxmlwzYIrGl3IGv+NksmdYFFnp
rOGZHDJhheV4mQWjUgtQHE93/tyPt5NMG9f69cuX4zdzHD5uhnC4SjcrkeIh2XbB
dAQBBJ9NdkmqpbBaw+yNoCL4vSbSrOQR9unATYGTQtEjNzZlrGu8nyw3Yai2Ufa9
ufBy5UM4O/rO/Ayocd0MR1JF+C4HjNZ3kqK4nc9x3t96s0ZS3yCtR1UVdf4nybov
6g4NB5UiRYexNwcS3v1BPFygfDr/3vxxa1yUW4DtYGa0vbrwkhWOHNA/Bw+Er5Dg
kS4tNrEp7fgviNAXr5ybCcyFyp94UcG45gwAtzfogY9iq42jTWXcIHkirqy6uBD8
6iLljGHJX6O2DoADbMmVNHkGNq6B2QSfVybZ7lD7DM9QCyfEIzpPCs+InM+Dan3n
oStvzIBPgKCiTyOxNpdAVJ7v1RlItHaR8Slnaz4OTxk=
`protect END_PROTECTED
