`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PxNHmPcXvTdAdRQLUlTAItcEcvL1xpwygS6/PoHRA6OmKfABafkStgut0LXxrGga
kAJdAXebg0QjjOd3Beb6L3YUXawyiiLAoYuRfNEaoUXyO3zJZpFmOO34xhe2CCUd
LvWzk/wS7YI+GczkQ/QJ1Hwb+V7Z85WsTJqrC69aE7OjiTTg4m+l/xVVQycrciPI
IKcgfRlYfDf7c6TcniBGJxwjGVaoESQkiBFqEZkmltdELAwIfC6sV25ABaegrI34
ikrzAzkADVIjISrS/+KEQAEz28V91YhTzhb3c/+i/aE3x5nURY5T8so1ZX4EdVz0
mLKasKaAOxuShhpO+vbUtpA6wV9hoIRZNd0F4OR1g6NJCmahGUelfJoOqI25iu7j
BdXpK+M2lIB80Glff/PZ+w1gUu8Bpg7znuEFBFcRL91X9ZqxxbFlvjgsWMtNgveS
oPLwHvgdF5Z/89ZTstLM87e3GWH38qhzVic4V7MwzFilXnZMF8oGPn6jgUPT1SW0
8nJeLs7r6qHTis2WYlugCS/vI4GGYMx+9jRvthz08vKFYR9WXpdYrvgyNnKpcqtP
mbQHH5/DWzOb1XvHtSa8XbI8LVbWhHNUMMo9Ex2DgIOXr+2ZdLjEMMRNPcz5iqEm
UvEYwfyu5yP3xNz2mRf835sgrJ5h+UgHa2noDn0gDwsS7Usm/MjcB9spACkWZJrj
wSTJRn3mRarB1Gonu8qkiMPcwazjHfw46tzZ6UMaqioRY0k4tVyu1OVVVVuK7Ida
cQydbJRIFFUWLM+Vw4NWudvklRSHty5Azh+9eOC8cmjyWKdwQNcRuCwcsQ7QCkFa
17xycTGQWOsRrFghIREFXJWxKjwbGc0K9/A9Y1z90vhhuOOTRMYKQFxXWgtUXzoy
`protect END_PROTECTED
