`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9KfGSazWi6C/P3MtYo2OaFRDHHXTZFIU+qrsy+FdCNtPrjokVtu8LMr6HEBI4u8W
wfDqiw+asqCryHeysd2/6LVh81R+w0CG2OKRFRUxFxW+SfFt60VP+wOu5NWZQYTB
MGre+jbo9s+GgZwkQe1C5L7CibzhWWf3L6Bg2p42ev+R2Dv43Mhzw7weJ4GnB7WK
UMmiUY2hcDLWQn6zEXYkO+tJon16g5JJmFMK31uAG9LveuEi/5kc40oUtwxgDYqQ
Hm7o65KmPJS7dDh8NyutBNDlzMl7PvX0RYX/ZPYiX10f0C0dsyKqMAoAmy47MQl1
sFqk6VBQss3fx+9dHa1jhV9J9AhUoBoCshkToLpHCTv3qhSjWHpRjpkuQJ6SeCbv
NOOIqdsoNpYWw54rBKgygTiX8x5uxs0e64D0i2gxuG3BO+E+l5YbuWeE5atGq9Xa
tvJHZ2I0eRPZ80UMd6SVBtugMJ+p8Gmw84io06tqfsSYiUKfVcjAQ2vSGqRufvv0
V5mcKcfJE8cJS0NIInYZ7gbblRKuz0081ZqcAXOs5StnUiRQl2jiq+FXIwphJFut
OepFZ24t1maX47d/t6SagA==
`protect END_PROTECTED
