`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X3y8O5108uHmoYPFshbDu+tKF3SxY/DXgWxF3I5a9OHVqsMGlcPTCS3kaN4oBvqc
Wf4cIrX8N6JAIJw9dqRLcAFeBn93DyHEIRXEqbrktZx9EM34jk2va79JrgMVHl6Q
y1L9KwQO/OC+LneMaxIt15PSjKVmsypFn67sl3HiF0hChb8niyShOw3TbJFuXjsE
n4q+qxaGXpeWweWE+4xamaIW5I0rwb7rM93fOjrULxCnIP36opT4wSvVY6a6WjIz
Ao9vLTq93p/YraLG021BqpbFnrCaxDacsAs6xAS2z3OqQZZxGldIcZ9VEFr/BLtX
h8bUdmm9IQrk6AMBSMe/ioiFVR6tI8uyMqBlzjU26oJLhLKMrCUOWLQi9ZPI4PKl
iA+DnUovaLJY+18F5LCHuEOcjUE3za9vRAaM9mmTIn/LrTc3yiaYXDkJOUDbjUBE
HMzJgw87scStDZ1qnQFzh7jAUFDtpHkpPpigy+vvM0etI0SmCsMvRT0BSY0rBL1r
Vz60+gJ9R/MMKp91he/nJCiqmwqnQoZTccraId2Lv4Vij+TTiJuWWW31HCTWB2Jh
qzUcvZt2ADWAuWsbQ/R7XUQFqdvAx/U3LhcJQgP3nofnkBgD2va6v27HqIc4v3X6
CJGF7kU978smRGM8D1pPe20SiA3ix7FiojS5J0oyEH1buDucSeA1U7zSsF54RNFM
9gjnGgeao0mvr4GvLj57n0QNidxHVQbpOK990tsce9uLcP6U7AoUHqWYB1jga/qa
39bgCakLfE/8+0dfSLUtLreEpAhHaFHT1Mll42/uFvU=
`protect END_PROTECTED
