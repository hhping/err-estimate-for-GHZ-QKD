`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4PYeULnfZpq01t8AdKzltirHV3bdELHOv2cP6UIqL9t/Soq+Y43bNkH1k68Wf+Wt
VBlCxOwHkij2F4gdqXV9lTi6BPipmhNkK85oOC5o79haR872PbY4roDMUcrNpkpN
1y98p2MYTj8e1rP8Q/cskt8Jl9fGprF4yb04RAkLsvGuFval6Tr+Ro4WB7UBHcG7
qJCfEzfra4SOxtVK/7sds1zp4yO/IdM40y8KfszqWTJf0BfYSa9ZzGCoV22dsqNa
Kh9k5TbVU36s/pDmLYfIXs7TipuwDRsAzC6u0EdIVXWtDvfJdzXbXydueRWQyOmd
jGP503I1037MtZPU/H7CwPsaXpaEOohYGwvowyAo0A70aXgmaQI/D0IeCvJTgaHc
9Ppd5xFEAAehRS/H0zLUygX7ZyyjKBTolb94FV4b0oRJWQYPUM6kw3xY3uc20u/z
eLlVm5dOQbBWfJrfzu4NC5tkFSOdXebTQV/ZA6gdGJ/utlZKhY3wBqpIE5YBlyvg
yIB+sukSM1/GOih4cbYGB7CgDEftAP+6TPtkrbNdY1e6zFFOjAo42bHrsdZnXgwq
nA10tJTIS/MHP+d9CWHJeBWg/GX9Ibs4KweB/lGmsjhZsxro5HAOcsZpEMrZHRuk
Fp6dUD/+epo8mcFr5uawmpEo/XAsJv4eckmp5Wu6seFy/4516TCX14j5a+xUlwme
sa0Abc1wYUHBxHoqsbrvpudNnYmPd80+IQQ1U8PP+Xev1BWS6QeWRyZbN9pvOx3y
KWruFlDesIlUnXfU755ASyn+llR7n0Uh9fltrJFv8p15bZZuTRNiHcSicZNH6JOe
t5LxNmbk2lzLQuPwMX921mxem+Erq3rq1oOpphTyp8cN6KtPFXll62gKwqRm/8EA
rttnXHVI2nyBOskulK9Pf0SXcZphrro+ot6JcBTsUss/iH70hJLxGmamJNLt1r+D
WviL4G+iVLuq81+5v8dzEH5NX1coBBRZnBDFb9b7lRw0gtNcLHOAIBz0DJ/qnniE
8vrINKJ2UKBiPPLKKjgAwe1gFoI++5cPqlcjFw413L8=
`protect END_PROTECTED
