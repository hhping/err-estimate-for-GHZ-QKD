`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IvoyJ92BIPiQtq45tIhhY7VzWWp3WGVBBHTrQRSjn+Hi7g0FxoPrYj7NXCEq6aB3
9dCelI9BOAf3mQMuO/zHJFmmCDuCf49VE8j+x6+Lj2ldxsV+YEikpHmwbM0uPXs5
afPo4ePEbSu6s1bxVCAmCT/S/PyjGHfhxmeD539et3IHay9u67v7l3RDER7PKi5S
qgOTCYNhaBzvMOqTqexGuho+c2zqcYB5n8AjqwLI2CctlMOTtjfOrJmULTuTB6A4
TT8xlfJlJRmRsgcHNdIQPx2ptGGhH0JSzE7iASx8Kadkfi6s+blOlCEWKEnpaB7M
wkQ4yP66qDTEkZrGMyN9I0IdZXZ/vOcUpRChs7Y/LIxnSFsyWhLPpfhyARcwObXI
KfGb8UVHF1cn6QeuVJTHBAgdZ4xooTlR5cUcBQuoHx6H82I71pDjga8S/OFJtZKg
ZsBO7Kw/VrUyeZ2AdTh8c81HeC2FHtK+k3sBQptcyOg7niIYvXmaWz6sqhBNx+Rl
ArC+ATXmzD/qSTMpkSFYbzZCt61H0JFCSmHmuUlmFinqc9ZGVO9mXK8CzfDyLR2X
jNrx4d1Np6PRTyT5Tldhhi+wmtlDxHZvZwNxyiz9YKew/2lfyNUqxSnN3j4MfKXs
Qyr62FtutLfYvD6V3lvrnz5OxKAABXztoeIpwFzwbilsUktKRyzGhXpDXsqXWAso
xbivYSe6wtkDk66u0MMfk5rJLkTuS5xP5q8VdLDiMyu98szLyrAGuRYdxDjcuJub
kF5MhxBZ76CqNILsgLjC74N94yrK7qTHzga2L5vA/hiBgei33u6pq6BZV/SpUxP0
R0qvBD287xCUtJAKb6jdJw4VkRAvScSCEFA8yDH2LlX/lhyL+hNngGdZrExz9eKJ
Ia+f2BTYGrTX9zESiIcrnOwodIVCBum/v10pGYXAxLzcC2/gA6c68q/+m3Nxwjs6
83Mv60daAF/HFhU0AJ6DQ2Z//FyIYIhbq0LadAqoypnueBzOmxxbP0sL8wS7Zrn+
BwhPcWiictS6TUjhd7H7iTBlGrr6UDYg47rMLAlwxfn7wUy9oeoVi+CfN9xBoIwG
y24R4kDW65xbSB2zvQQVMd1BWFyRJ5PqJWr2mrN2WHGQKT5c9MWn3jlIt/aYRPJQ
/g2xjabKdoaPhEBR34PH8yy7OMDPsBKzlubdxIsLWICEufGycO6QDwMg2iXy15oK
nFn51MsHQ9hVwhmKP171lqiYhVR6yMm10F2QnDmYmLDPMsawJMGH6i37b4mGa+Ln
Lv0IFAmestWWlHsK0QJ2UTnUDp+YBro3ihKXxbJddq4=
`protect END_PROTECTED
