`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z6uQgxW0rUUyWQI6SrlWXF6ts3Ho/ZPU93RW24IguX8K/ji19vluE/8ouvJoYN+p
OPUkSFzXAaZ5LJ9p5VZ95T1S2TV44t0ZvgoXvh4CtLqrQ8pw5fzVHMNW73fjK27r
PuGsXbb7cuovSz0HBpGQIkBBLzt109gyeOUGea88xlrkjvR7lJ41NbuCQQdyBNmB
XLAUGuZ9FwIr8N3ZowoxLnPD2ek1SR+zSL+3QYdH4IRUYLKhI8zojnpLiOn5rP1Q
xvkGP79C81SPWFuVOgZCGAUCq/Bz2obCkaQxv8GGiSehH7qfGib9/mB+dJqSNL8/
vv5TNF3eIbpG/Kbu8zHlYgMsurXMfdMPxibcO/iDI3U=
`protect END_PROTECTED
