`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6jQOS0QU7hV0uyDLke/eHlvIuebVGnuAYWmD3cN5MoIRpxiLtlAsIe8aB7y62Qsm
kaVbn1hNHxb22pUSAxUvLylWzBLJRM9Bqzkcfg/NKohhPkoi3+r8yPq26T2Rb3j1
0SWPy2fGTo+R6QhRxoNZ0/B3entNNOainOhxafuc1NaSRo+jqVluG3xRgph7LoUh
xQBTJiI6si214Km690qtM/ULWYhj9BBSWyFHIyyKUKApj3d2RrodaNO3uLp2AkzL
KF4aH6RiAx131tK6xGx/uvojZ86hOC9eIDF897HkNuFeAkjJ7b7dJ5EufnJzVz/Z
BquqxmQp2XQFSlE6n91YmIWwyHNrohClN29Aucy2/1VD0HBdHQCxmfz+q0ZxehKe
0kB6GwG0X+Ae+4pVR3UsHuxbFjV6f1bmSahgBA2mTtNTVS8ySm4qjpQtYkBSXnax
SGeQCi0bOLOC7GI0aelZy5UQ+qVdR4zR5HkReZUuoFaf6awTpMcNYO8/W/DAY0KG
FHmB3QsjRWhGJusMTJk5GPVVrzGznp01RqE7dX8MPqyfnAQKHr07Y8RU5CaupFYH
5+vCo//d+83uCeCjhbOd1uufcNlQlmmtS/XR/03l9ROqtWkPpLBoLVmmYyIeRK+G
gjViIV7ztKDrLA7qh+RB/i8YomS36LiJVo1efE7GDrAYCiWZALdS8+v/keaxq52i
2T8CBfAXXZurT0+eaVzZ7K55lbDYccQuYEcAtUemmUIDfpXDlIiHKsZB+E8j/MmU
SLCo6YmLEYFvL0FXd734e9ychvuzQBe/fiTYtY7riUxEvi75dF2f+Ian8VxXYunw
4S/bG78VkYDgqKRdoD44tw3njpOr/mZNtWPl3oT6taoXym6FzVCkGGCxhN/nN8ng
eqEeL81eQQ/qvTx6xVgxewbwM32JcupCy6z3UtFzuR7nvTjUt7tZTDBNoGeIOxlZ
LZ2LeFbdet5htSMc0m41DvPMDQkhjXDJZ5Y+xY0Ned1FWvZCwqbaRx3RRyNGIvDw
NzlI0d5lixxVoek9zdWY+mGNzZSFL3iDhAvG1Iwqdtq1SkQEEt3xepTcf+hIhrrz
Uc8dIEPhOvnSy7PfpzH8STuiWBVE7vVH4gMBXc/PkrexVPsEfZBNdORxqqtcsauB
zSUfGB9Qc16tMDMYuqJWZwh/gnW2DSeNavjhu7xZFY5IH7hexgXBEz6UxdNbM85c
GGB6zWN6Y+tAMm2tna28VCwt33RNx+NZHSBOeyr0ZcKBwdqSLqhGb9CNprXumUm9
87I+Id4KVu3WR9n+gIYXC88nNhNezVcFnY8pgRsEYaJj/YSLaus12ityKpGx8fJP
5+WJPuauxBk4URZqrNXBrAuBZMdKF2Rtxte6gW/cRKM1dlOyb7jRQMZO7udU9Xu9
Oc9i2DCKcDZBCeVnSexPltevQnqD+JIex5TnULW0XjQ8bSrk8WFSJXHsPrILFMv/
L7AvDjyUka2c3u52kXytLYZIl7+nKlHlBE8MxUssXzhhemTQh8jp4O2CYDiHOz6V
Tox1FK/Rfsf2VOlNUjJJjpoFxzcy0DWDNGRcMzi69FAUvYTPdFIdcaiK3Zb8tcMs
3xI3puvh4L/3cGUYtJqNnu61gvWTpHtTir3yWi6YB1V63l/etRtM3FDbnaN8CEAk
+1AqPZwJrWFiSAjOUcapLn297ez6CXXkPl7HIbEiNF/6N0C0J81NmEw1UUbo0A17
Pt6rIh7TCKKiBKA5+4SftYCEd+f0Ba0YHa9V+bpvJMN6oi+BKnBfLcahunMy/N/x
+Byqaf9lpD12v1lCkEWySXn5hd+jJJSGzy0d6HOMxiSpIZnKOfvANJdyhinVn84B
9QesoEOXIjAI8N+cVCDNdz+Cfm+PZWGpkrw5ERBL5YTzJFhY5zamfoeVs+lAzmHz
hA65X7Q/tmHc5Uz0oDj4jFJVCXgx8qMftA7CTR+9+CE=
`protect END_PROTECTED
