`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ei8kVtTx0D51dfbvncr41oSxVnCjIDryUbND/Q61J4NKK8V5C5enzmEIaC1PYtlI
WkY0mBoiVijOYuaTOrJkNjwKURTejpfHTJUBceBjmcc10DkRbm6YNlT7n58X5Duw
2JySZOcUB3yYHmnZhptzrzvzTLU9vbUdE6xok3j7WrTUjQNY8/8OhEKitcd/V2xZ
rXRSRV80EDka66HjK9Lz8gWDyBS83ka7TjscXKRXaDisBWfx7WJHbiyqh24ZhFgG
inBIq0PoatjfHGI20nff4gBLAgWsF0g6uQHacGSBXvKMaYNgsQydXNNVgT0Ce0t5
ntJJH7G93frMGBJySqEVHxxH1vRxk0LN50tY1njJ226uYNyI8OM9JBwHx+tZhxA8
E2slaWa2h806Fk7A84FVluO+S9oV9f4LlLW1NWiMAMfT1lpXH01IhyJZXeILR72H
XE0doaVKAj+5J8AvzpYyiPzvGg+BaIvYhZxkGCrCtxJReupQgJa3dvyEDKaV+1Dh
7jjLn6KKg+au+1aSunmwqxPSrK8a6l70TEVSluLhDdkJKsFR2MSQYmqTxFZRUL6b
OXCny1Yrq3tVv5QJuQ9kQ+gp0SXjPpak8mJTznlhE+Gf4GS03LNtigCtivYwRhLt
+xcEqUryqoUhGZYMZ9xyTQTc8LjoWR9cvWZ2O9QSObbubsHktoR+HdpLXCc+Tqoz
4aWo1p5JxqPhLHlUmDZgaO51JJCrVostBf+lDHneUT7IB6AyDcUIfpbSKJ7+6HlN
wFY+CcEpJFKXDwqY3QXF2PYgzOXU0+Tm+aVhq4nwIcLGnANAFV25mdwVgWtq2A/3
`protect END_PROTECTED
