`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GW3NXPbslR+vnM3xgLSsnYZWzLfoUiYFIkFveuM0kUIaiDUFdfGP2H4ZcIIzNVwM
sRniZlSmgIoYmt3zqg13Wn4Y7FTJIEI5J/LnnJRVTkKND9EnECwobL3KWtjDpMjL
tryAYPtcpz8tFk4thecZr3H0zAtbfNjdDGaZOYN8stCEY3n/sFX4AstMHXWESkZf
1znOMQ/hRXe5TC3pY4oCyYGT7HjGfck3+3+zL8rdGq38oKQXjDZJ+ugBZHN2zZnP
puTf71eTxlCnT30cqNUP+QswJfvoIavozqkc/YdX1NFocORxjgONo0utcsJE4Qb0
dgCWoPVc9eNGGqTv2EILZnXz2PYVObTt9SUyYtKNG/k8QMjgNZhs+CNeqz+bQLN9
QkFm6T/jtJsANJsmp6vih1eYyD8pLymdLoIJOirTfH6gq+CcDEBifWISFpsIMVTs
kdY3kme9M6qlQ+fGIEgJrPqDdB1hKUo/PE1wtrtYmY6dldYeKtzwmoOVd6rIuXyV
1URqm7wW62owlQw+ifYt8XOWX8l6DzIuPVp0DCUD3agi3p8wrYbYcyp9zIArHDhw
UH1mlplG9Mrdh/O06uRz0Jukv0SZA+EQpwj+RHiB9Ehd8C7psnXxgXF384vGtqxd
315Ii2j9qgieH55NViNGt5Z317NclMjrsr38YSzBs4TrkfAL5Zh4DShfLxxPt2RH
1c9AkqlPAumuUkyHpKxUrGJYXX+7Ps+yy0ZAGE11wZVevMJhk6XWpV/gdIY2j8gL
e9xkN6V9NuDlVwC0Mwkuy/HypSEE2P5TXD/mtbCWTGIfDhc7drcoq74+XJVJ3sV2
CFSVOpmi/IEEb25bJKL3kSF33Cx9XvtWr4MusWfkR/CS9++dM5k/qW+FjC4R3R0v
CYpSHurBh8miVOAH1bTgJ7ot/vcfEiDNra/nPBHtFtSnAlyeyUJfP6wRFPUMbmKL
AM0CGJc5rGoos+qpJJdhaOu57pBkgNlSTS8Qe8eFbcZgn4faydnzC1+JxL+iBJ44
UlxjPDyIS3lT/iXHwYROuPjiWGNE13aicxxRT3leoiZj4/Bhen1ZCv2UPtExkznb
bRmv4aqmnQpu2U/CNoo1qtC2idjySIIA/4XqlKkyTdQ2CowvBl1R2chW9mm8/85C
E85ZI7dpGR2dSe7/+2VVdSOK1n/s7tfeugzKO+wofKE=
`protect END_PROTECTED
