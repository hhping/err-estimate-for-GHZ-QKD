`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PJtsTUfcXv6mj8qTnrXjbIoLDZy5vK5Fs3v0KoujmGBAdYGhKARn0jkDAYWEiZBp
3xFrARy4V19UCJJzwqrsu/Z2M7kV1m3CkcPHTAgE+azxvA7iNc7O+5LGLifP2KjP
CfXZmRqzFFbF1shfe4mcdnHNaG78cz3NPngveJ0qeoJ6NQJDmfx+Rc1hK/Be2E+h
c5CknxOqbdiueBxzCFl/4HSC1tLcdpk8SDqZdi7x2+A+HR+jK5kZiP7M8nNo5Og8
DAZ9REJrkS7+Yrxuk/lpuZY/HQDqr4L3isJGTK164UEFwoBf6EXqek0xka4VKzvC
Z6f5h5fzM0BE5/GrtJ/WdKKmbPmMo012WhZxBBvTTdg/dVBAZiqYSQdqhZNIk63G
7GTComn+PQNmYiPHJMOIR4mVjozXeL0RO5qhT792HeLZ7u8ErAXOwqD2gx+Pxjer
njjQj6BfXoK603YVw0obZyABtq3/L/3CjO0tdprC9NeEf0zX/3ciOvhNvGmcAJAR
Fhyev9dHLIRDBgfZT/ScAEqmavqOdPihPOaydPJpx5cyfOU/QVR3NPGiQ/qzzLlE
Fk3ZsH0IJouAM6JCqlnWGZWMN1Pn8GeGQyfMdxT8BEnw5tYA21U3MNS52a0vE1rm
IJ9bo3GQHg2HFPXIuLZQMgtyI+iY7Vw1Yl4jR/lffq9qga/JBtKePQA7nGxBkig1
IWJ8vdnWGor3r803ZVsJ6ZdxMkek0s7yeBti8lauwwAe/GNhDFskUsYaBXVQWdYj
eGzwPftc0iLEKlu+sKIOQ9jsTmt2v9xu/Ftztlg5lRrg7BdJ8CRZHqNBVRz1q8tg
boZ7nqZmia7sYfTbWbJMEgG58WNWGxoN+fKhpYkjLAFgZf76w8np+aWT1G0l7Z0w
TaJE9gzd13HAGg1C1snh4twcAQptLNAMyUIqzWJU1NGle3wXnj2mzljHUq+eowlp
Q2eZm2wWFce5xg2dV62LlxRtCbKg6ZZM/0SkK8X49XZWII6g5hNHAoGbOel2Fd1S
tRO9fTsuUVfT/C++FR6njOKwcliBd95fR44yDYdaccW0mWqR7QgwH1Sk5X6X6tqi
Zl7/nTtcK9IJ8EPwyRYnNSnuKjXbCjKvTFhh+CKpRjoJ3ZmnAZS2O+37L9+mMxUm
Ijl3pccKTFuQfDD5QRVHusgMMevtwcmD3ExJ8qKek+UHgANiDvatGR6oFVLyrKIE
frPDYOkDirqNJAjl/jEJYfl3wpd6D1rQBNacfpPyOPRg1jhUW+dM6963FxlzIyEM
Lq5xzbRbyRaQIDeT5nkcjWg6CTK0WlHw7k431jFkGQFXnehnqLhfbjGcaIeSp80m
PRa2Gy57LCTiVnFhV8Q7xlPHmXO4iL4h9speq3DEh9lFEv88XtBBwQuJGm4taXKP
QMQ7YycNtbK51WsLqUlOP8+KZiXf4jByAAiCPI5h+kijrHoVFWvWemVPj10de41R
gtKDfdCBcWUcL+rSaWmivXkKmQZjNOzegETlFp4Gih91pFhfhbllep5LhgloekvF
uWm4JgmNKWYY9nTIpqMS1+d35FLLs5somNM1T6Y8100tDvu0k+xmsNejBVd1FMwB
W6b7uRVYQ2HBklrd3uBs9b2mxCJQGrIDbhXrieUFH9rcQOvuFatHfMRYO0KrvMrh
trGcOvJO/D+dBnOFuLJL+DK2DM1e8ezGXio/9YwgJvxPwY7yvqg6czmU5AMDXpBB
0nFvIL183HHgW5ojh3WVDyIO5zfxNg0LoN4ZzeSpi/Y=
`protect END_PROTECTED
