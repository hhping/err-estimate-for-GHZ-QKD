`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C5K83PF+ESiF9tDdceuLLuuYWeIhvjKdpn2v7FAotdD7vA2xtgQj/uCohQI62BeL
4XXLcbHHMy6UY4HQxMvlWsgvQIq1WsYSHf7kUaGvd/Sg5WyvK7lCDs9BlYaXoLLU
wrxPLan/u8s/FhgTUkogNzHHyyaanTfGmAtV1Htt0VthLyYl/FNgdOX20D3ghbO4
YGOeZrduei0+tfiPNKN/IxfurCmBzDyxDG7Qxf8cFwl+uMogNUz3ty61bp5wvhDc
QqmDqKpVP3r2kobh1PWTPFSKhz4qJrool5cwmm7cCbG7sq7DC0tZL/zp8GKWgV9P
dAP+a4BaT3QcMsLwEb2I141aUxy7e367end7vWL3l5jmmgvzI/vLg+85hLdc0fee
kSBfK1Uefnjs3GdYTwzhDCL+xB3Ad7CFfUrohCgpKYVy3lvg00AiKOR1L2lobyl8
9lgaJQkW2HjI5duZgrgNOPuWXwLwdJLb44nU3YW8Ic8znrsetY7Pgyac/EhkBy2K
oTTiENEvD+RQIhScvxCDSWjBLjBHTb0B3PXCuUOQU8975SzTHFzquwxN3rbkKC+7
5kfRInAW2T765ofJwWZsE8LX7FLwSSCcTkzaC7fj+k7posAdYzE82ESsREi0GEye
m5+DRjYC2Ti1HkBRCHwnfISPc5vmJMMwewMoD6rTRXcK/74KZsoqdPOgetA1EHtY
e5dYaGFxkCbCsvwLwPoyyV4bXRuR0P4iZtAY0YZvj/JKwnG9xTA4uMyluKkJ6FSw
+KDI7ZFVJXStHJikUFAlVE4yu1oFfWzFadKzYRryENSQbCwGjA4vlXtWwvzdCSkx
mBNLpozHZwfguzjce52R3oLLLWTINM7/JQ5d/9wHenbVpWHYeZBplcGZEhR/NGXR
xl2MlOxRyGf8cN3nKwGygw==
`protect END_PROTECTED
