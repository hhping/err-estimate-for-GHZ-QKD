`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mKqJd2N5hYqbhBhWfF9xBjB8SzFF5PanQjvqAiei2Zn4PK9kz5K7p/4Rc2MGrgz8
mqQSON/vEvv6BnkiFBwFBvM5S/tTEEp01N9tzHHm0r4dFXejzXI0kBxaVyyOY7C3
/YzZrrRo4XpiINuQZPQT/vQ6EdZRuE7ch8h/2qR9xj9gv3juW+jsBDiPeheTe/9Z
eg1IEyfm3L89MtW4lrC50iHAdqA+Ey7/KZzM83EegotmwcZVjwHvQXsWRmLDswfH
ufmPjMVZpoaoIsystXzQaQif74GorNJmGL+359b3INuPt8TW40sTMNLXECPy9zLv
Y6vNPQ160mhtvsqUMutYpjWjWEEZHBxnqneo1Mp8XKNryGcTrU3fWvHysbZcMMUU
mfy6agr7HiShrgpOWIFjSG8Sxk4xE5bzJHX8qG2U1zA2RN6zcdouBaUshY/Wv2kf
iaCUIMu8adLqbPBeLlSijIvhfbC10mcwo4z0iSyz7RQT1m+nyYtQ4DoegQ2sijMH
nfQgsTCW8OmDU5kXdApJwnNXMACKgbbDzpWvE7GUlwKKUVP2tERvHTjUvV6I81Nd
3J1EFmIgx0GDSm0trz7Bho2r22bWnW5XnjoyYrPkiyqoMCKLQJ2U2a9y2D/3vhCF
gtNy8U9c5D9vB4Fwbadi25ujglk7nE45QgsxLoHkh2WeGr1Dm93SyIUL8b545r/6
A/j3388VOcdnNv4fuoE+HZ/xtlYSHAEu+6eoyFSSNbTyB6ZncoIWpip2SScEVr4M
MYmFVeWDQr5B9sljZT1H0OhjJfA8cjun4ux9i38BsjWJwfn7zcGzdNxb15kLXsEd
OrsLnvpozBT9Y55VKUGcJSfCeS8xWPmfvRTsnp6sz4rn3I/O17WHiI7uIWXRq3Wj
nAB4cp1Ss8UluC5JID4Ms15BfBeNXQ1i6eONh9Q4YuFiMUIX5ReWvfUzdxnVsgOY
m3KL1afjJu+VawyimDKEpP2LWVfFaQ9h5EEX5Z4PvBOquXZb3oWZqqFYSlTB8zv6
9jAhqIdKIP80FaPvj76RriSCNk2koE3+AHuyYOYOHQiRTmsCMU/b71HLXjaNBm3C
LXKhPlfmDYVhpIId7SH38PN8ElIWAzqqAXFJAjXZ+8ipIiyD3JJJSrIafWtAxndx
2kvuB7ZdB6BHCWlHvcKMYF/7v6vereZmNtRjWxwi33/MYiOxM+X9P9FJK4VYnXWJ
M1Lt8LQvaWO42sPRRbMFfJDLBuM1OOh8XlX4CWneLJFroq1irTHLQFNqdVdIzwZs
a6zf3y1Y+xXt3q4fHuGcDtCznAp6SiF+hWwfQthn+1F7aYA6AbEiexPXKsyDYhPw
YM1IWSCzOWxc/gfPzF0TeRDKRLQz8xq0B8kvn/QR+I6QSOGvy/iSoS0L37Zr+0S1
q0Dpj274bHhc8gvb7UUreFJ+iLuDE0ODTfZw6LhFvfhNoXEJIY9xlG+IHYihpDPe
Kwlp+lxfxqdn7Z0w3do7QRjKK6W7/tBZSNlKZ26qdfsQ8fYeFSJOzGsQLJ3yuB/q
HH1WNL8VwIDEd/Jdx6viPlMRVoP5PxRqWTRj8zmdqnTCYAcBm3BGp62x9nlgAUOf
FONdYp09oR6WYNhwozl2N2vdep7/WaiGoVpP9HbaMYgHZShCRNFDiuKTy4JHxxek
89NuApt8BR3ek7SjM4iQoVtURFpzfCbBXzP8k003cPtDvM0oWvcjcsapLMiWbEVQ
KHiWQ8JrNCvFxSj4jAwWYDa9LDf+VX8Y7SZKS5uFOf47XfukjsVxMbFh7Ud9fzFT
MGf63bjfQ7dliY6EXRNH34eA1J2QVj+NFvtzA+76uk5pogpUj8mL3wEB6Fi80rMC
j4aXZwt2vKnA2Z3XUIUZGfs9tRNCzZSdzn3pEpl7ZzhbZPGozsRmDzIXL/kiK1pi
cpLUFy4cZvBHZvbf+8D0/f0io1EEOyah4fbPL/zoO+Ia2wjx/G1W2IWDjZNJMlmf
MsttajmE0XtGHxWESNScOT6ygk0281FnT3mAbTQmXUXo/tCw/5SZUWuZmkEy4+Eh
GCY6hA/UBqFNddO2yK4TUnOdVRxYZX5JobutDCTroojQF2MMr21xN10I3z855csx
KHxIeSyifQLRC0dampr8odmpWRXj8bEyC8zU7+SHyNdfgdzv6ZeTd5e/+isGYq+T
QL3iMZzc5NgZZSPkOlMIEG+uP0yY6FxfK2QubV8NoKLEikPns47hRY8WuKY5RyG4
SySDMwSpL/i+TX/2nCFP6a6bIuf5ATtkbwo8dX/3HV9sC+gl/FrvMfKn7QspeVHh
NngBiS+My6rVWvuRRTeoM64LT1jflB+UZbvb56QdW/LW6a8ZCryc5bFCwWszqvo+
CqOyI7Ir1RN2gWuTmavfvEDJboNF2KHMyt4KmwkuHWg+xSgabQ3e+3KRnyVVFTGV
UpDNQ6TcG6urpDWCFCGj4xAcoMh2v/bGNpZAeR7nVpjhWmgWeSUyOx2DH9zQ+XD9
5UrP3hk84+lghP8Z0SfYDe//ljKm5bwsNIPoZJx3+yXxWdNcbw2pGwbEWNhRpcA4
OT3aUeS8YucmmSzuoRHk49ADL4vsfcFuvvqX+g+/0pxVA6dTxHA+3YQiiahiBcGG
+rQR36vjbI1wvX8mE/kxvSwfF7C9CLC86B+pqpCRzGB9l+lBsPT0FccIA8RRWCJ1
fnY2HVYLfzP9fB73s8nPRw7MdKsu0+pww0wPLVuJ1MzN9MKA70IFsX99IChVLxTa
FSRXkbuyYiqeSwSOKduOrR8xFaD1dCfaTZ4EcbRBVEVjm94FFyzzAeDrj1OCpovZ
ddrPZrNVz2CDeq/MDJygpDdTKqtvHZm4h6v0iaUQpStxCsMVNPHGBozbl6VDpf2x
4GX1sIxiT2TI5U/BQOh2MUFEzkUbTiyTg59acCActkX6moMM+gKNXV97dfr4HPza
WKIOUqFzbJP2ffS682Vq9qHtKZcJ3cSfobRVwsSEv8XyqZQS99IXOc0xaS4Iw08P
t19ckRATwBWjIzXj/OW6nS+WSYYfEVIRFtpL/Z1dVGwdaAhtj9vQ8VPhiAUiDkX9
20OIhwtXdPDlvfKg+WFqRYdDcREv9WJ3fTzFy22r/xdfvyFndCvamjBpVXKPFjNR
H5S01pakQ80QLAO+yREjT98OSoaejy3A3JXGjloAG/DzDbbuTJiX3gLgP/iDuQ1q
11RmbTmXt/gg4EPjPwnkTK9L1Hiom5IJvnSQu5tk+O00iu8xKAwd7gjI0uz6YO6l
GCfYa2W0F8e7tUAjWnzDFSdq40c/pwE3EJ15OoSSarW/JSvteuByYnWbSyxbckPh
Fk3tDcjSqHxOsTb+taJx4Nj8PhqH8vMrMyUEF5viNAn0S3sTLzrv14egwSSUrHq8
zV4Sh5PWm2Ra5mxZez4W5nEKEpeo9qugkVtk+B7KsBGcSwBoNlB/NL265RLv5r+3
PyCnrG02me6qAM5XSmXY9WiLt3VB3suSOcLuyzbS0P/EW3iflqpEJk0ODRsUI7QQ
dC/t8d0fPOP4+9rKU68lq5wN62iyZDlRKJNW1MCIILrXJ+QxZjCjQZVXBgoweIHJ
9+lqATbMr56DWDThFVjdOhUIOm59f1G3bzWlwh9xAQB9GezLVT27QIagAXmNiXHN
JX2K0b/DMimuY5yrYpw4WZDQMd+ymFph935qQ8OSiIIc15LncOMhObMXE/x0s6xP
dmnGX6G7cibejeMfJwPpT7cFBQr3qTbgeV+vV3dTr8xmQQAE/QBnoBcc9MxcKzsF
RK5qlNJTYmkO1t/eqBjiN6KTS4jshLPjA0gE2Yv2N1kjP7EdZgJbfADHGKj8ntGQ
Z2rhOty1Jd/Zqge1uEoLzzONUas0I535vvh/cs1AdEu0//fBLwxfCi/6J6jiP+Ju
sown/YbQkJ3Hf3tlxoRVR9BWnDyuGSjgpAz0fOWi8Nb4ow6D4yf3QYVIJnvnG/lt
1oelRKutNpSqlNz+GAI5bCXW4DqiN37PLFytcDmn5xkfy73wefT60sZgo97IvXig
8AdiicjHK7uZvi4x29k+umnbAKwDstovpBDAXjeFUHipeMEWORqqnOpzJ+0pDDHQ
Y34aH1lQjoHIs4lcCK8/d2ubbevuQv6twXwzk8TIwGJ/M5oHm6ll+VG7dbvBcWVX
9NFy8xCrVybDSqBdbwyClNFzxtTR0PmtHD67OhDMMv0BAaVmXguupdhFLa357cn/
0ZKPtKu2A6G7XtmPZlonk/lXl6jP6UAudWo+vBNLpljE1xER8ZpKn4JjRCHXyVfF
tWHzpItwmzYULReAMA4oOU2xhOY64SGiJLxt7TDT+zsg9bPAVoOOoSLy8+8tt0So
HusUKpRxVIJqJaNA83GuSe4FCk9jZfWIYGBQn6xUnJ9xaIz2W7jIJdm7XXakMSO9
ccfMT5Md+A+BMouWL3/ZqAnwHKT9bJtvuPNAxojnO0/USt94xgIYmA/fCSsPl4mU
ie1W7cIGQqw3H9KecbYfIxZULieQD4Zzem92QWyWcEmQiETmEAKATqNeKI1RUk2r
OqSVpTTfi/K/ZG9SbNlZ8nbhR73tWAJdW5dJy7vIKoexm2SjgRhflpRP4z+igOWY
mzNv74cDDMYXbno7vpLBi/ZoU+InuHnbx6LxdKwpGvqGMJo2W8sHJIy0m01aPpYl
tIGRJxAGBYnoyYmquCXaHBrWi6o3uyWRCAbv0ShJpR8502yY4uhBMxpRU7x9D68L
x6Jfuc4Wh1DUNIKqdfXt/BSxnnSsyXsZxEPCQj/XHRvcsfcNpDUlhrDrhhyqaS+p
sQyVfikEFObmHShglDHfaooo9TDBHHgBrkFh5UdZkKi1SZnHlvk1K3yKFd7zCRHI
eOuSOK2kbXGiQ6ewHE4xMCSTn4v5ihTVk/6lQrTZz4CP5JQ8QHn0OKn02SYegQRE
mQXA0ZB2CBBF5ZUTZb+flzgGToLWnXuecZKYKgx2SttYXO+hsVM6Su2szNFyCzRy
fnfYRYq6ry7dq2qQNGJfq8fkniynNrpsQFvMVU648BEBjjnInb9fwAGJeVY/qAaC
CAJ3yhO3vRAHCDrvFGA2l7stWhuEsUJHvElbrCEsFgPI+gkEZfX96X1T8sEZQ99A
1SJPSG7Ph33Xvl5XVEP/YFrY6jTpGX8Jm6RYBuTQ9e2KS6e4/gDlgUmiUugpRZee
0ti3OutjW/1+wDCVWSzlqWCVInC4qGRYo8kYyZlLfX2e/XjS4pZajGQEaLd6Ummt
vPM2nmsCKXud+0J1Ceq6c6EUq4Go/S9tDx1EeTKluoijWhxHCi7olkqf99SjJ4RR
OOQtdrDjOllJ2UhGAd8nY9tcGkHMxKQd37YIpSqphGepn+PlVLJcAVf0Er41cTXj
Jj0sJpCwNsQZ/nzOCQuRZiADNQce/9DwD2snIJ/SvcjDcuK9oYJqwjolJvO0tCmU
DnVbZWJ7xBpdvL3cuiQVLOhmv2CsgJ8S7V2GDoLeC22YJG757/9LJQtk8v01BpTd
QccXLvrrsQsFyJjGlkq82Q575/O9a05OUU2iPvyCzuIcl//Dw8oRSQ7AYs8r6mP3
/FTC5bf95t4FAVFnh8ZzFxpgqE4TXEUccasq7uqseswTcWkAJWrocB+aW9hn36o5
12wmwgULT1V3x08HwrWYYV5+fLctQRlc5AgoZY/KOiM+i0VbA6YXz1K+r3Epr5No
Pl4idzmYXadCUQ89F2929a7BCRZZOISjE7YryOZrKqQ39p6smV4koqIaalioaIe4
sElS6gjVuRDmRMNk0ONvnRx6gdrkHUpBq5DgJ/VPDH3AAj39StCAhd/Y8+ZWa2nT
MWb1S8S+kkZE66Tcw4J6tJZO+K3/070hT6GBe2INmQLXqVH2idYCdHxpPNxRjTCo
tZyoZVX8oxjtwNuKbNMMuQl5kH08sCvjQ+XaU3u4wI69vBsuk4TJLRubk8yKijpn
yvyce7z0OghQVaT+Q5Fxl6kNOv1fwp0a0BkXXoKrKGmNs/45B7fB3jXBUX9YNFEX
MptlJUVaTFGgEOoL4Ki1qIpWiUfYX4Tvt0IiFQuTeyT0EZWcl5fxasVCKljEGefI
6pa+9EGszV0Xthat/JNWlqg1QcA0kIkc8G9e+TC8BwnVmjR7mfHnnB5ilEz2Wjlu
EHOXzNO1g888EZMkygCokFz0EA5dL9EkXTWy3p3vI+Goyg+piSr5TEqBcuNUeQEn
zTnkAlwC41V+GW83WkhLBd+IAsuO1FZwqoUeSTReWMV+7P4kD3+3E/zxC7VGdgVI
iBrV6QXCRbpxNpzCse7wEgcKFWS+TwMLdfpRb5wunytSNRefasI0QfvY/9eR5l02
x5sOBa3OmqCg58lDASq1sHUvELLEYGx6Pk+agSySAAzy8kVAk4nzGz/ljzzkFEVD
026yPKK7cC18G6WCmLNu4vEetDvQk7T75x0HrUj2N8s9DIai2WRawhkM1b/yRz1L
kqMseHdqIrFWqPL7x/hKhyQYju/xPgmQekWAX2nf1xv8zYZcX42N23JuTOYE6kuo
Bg+M+brcrjJ1jsmfSaIglAVDz5H5u+LiBpTA5eZ8+HnGC3lXmLlGSPQUv94jgYcE
HbP9LOqUSK/gRlAD+m9Viyr+9i3dRwAeW+74EtdewDSQaNs1KHX5HB3j87rMY6WZ
2cC8YJVWoUHILh0p6vjiGq1F79yHZ2M7CUbIEwoG7amRQatoyk5MMarQ5HfgeKrB
N0XDl9uqbUeHmFy/prEv5nTAPM1kLhow4BtMzGQQAt2r0J+j2yxsb7Xl2UimlgRO
Jbqu2NLA+STpuEZVv+iYYdi+ZI6o1NU6SZoTIbVlRfXIZfs1vvYRWBogP1mvc0Bp
5+G/37KXQFAxaasxKz0kXoT9dBDcwCOCLimgWYgiXmzkPvqcSX/BG1WGHnBs5gek
gjaXZDLLzk3/llhzEBqjkJ/Yh6cdtF5KV5lJh2u6+iKtadEHzZs2lEMr40vnYTlN
wrzmhrmZo/zNZVDRrN149ZnI3mEG52cnhljmJ2Xz51ofn+UCy7meYF5GsRVzgXiI
rjCwSVmcRtRWlKUAMGckbGGB78pYpfmQpqgOgEqMXznhgSEWeGUKjY9lnfZm+IjY
KmMV2e3SlWaxuO13dsL9Tjbdc//hg2U0teGOmUOm2wovmvE/WaYP9Ar76nBwXRWl
aP9Wnnd98NPDEBWIIMO6J04spaFlPitiiQcxd7VJWqNKptB5Cckg5ukA8SIPKgsY
GCWg2NmImR5YGI01oZbSNIifoBbmkvPfjYVS8Z7Yaspl7AHnTbhLMM8+6XeiXwrq
/Y9o1jzQCJRQb0nsuEmq4vvHymnXzkjPV/iHJl4dHIHfi/mKQHUo7Av/9UItwrm5
ZegMX4+U2YU1JXqhei+RXEk0wm2mSZ4IxChKjHYmZEUVV78oNpCqE7o6CH0Kij3m
5obNP6GwVblPp32uKj/C4hq6CcgCLCoQouCkBbaSi9JrNCjkXMf+T03da2zTzQs0
W7YEVp8qurE1z+Z4T16KBYtBaOIEttAD97/cXMQSfrZ/meiIGh+OG8HxtBsNO2Q5
QBksDIRdxbXBUon3ppJgX97fKx8Y0O56n55UxPIbtP2P6t1H9C11maTWOxpLB4am
3gpbJHQRyYYW8jlI8CeWglLLD6aqSdNqx1nNn+bgot+gZJTJ3e7MsxEvuvF5aXCp
x7ByD6CmXr0sN5G8s15dyqmifBpqN49U9ItyiseDOLS0vSy6vq6qHpTBbCgNGJym
GyN5m9STtw55F8DXnrauYY+vcmJb9cHoy416Vgc8uzv5w0sfXO/z/BfcGQXliDdE
VC3apiYa6cl5tIJW2OPLRy/Zj/gdDjfw3RoetKEfpopoPFRkLCXJKulihKEq0+Fd
7Xcb6GiJaMYECFt/jipHT/arhE4IYmQI9in2+Wdb8kZL+8DJ47DBh2BV4Y5ZIbxR
uDJpiI+KWtedPtytk9frLzRLr7KiK3CyMrQcrWUv2/TApIq9QmvD4CW1csiH4CLQ
GpH7C3VIlk7b/Pv+gGgQEHZeFHdWg9oGP4Vi/FPxGo0xQz+aJvDKND6DZIHjPePi
n6RvUhWgzx1LaPikva8FEoMbfRpqdTjkUwzlHpVdSHKTZZoWpp2HxLGiRoWbCWv9
U762jiKGqo5agRNcNX5K7bh/4Nt/yshx8ypWgnN5BHrIS302OLjXs8h3sILJjfqU
/2V+W/KJUBJKwxiU/6ASANDOiVrcok1Z9iLnwVomDophhcO1hwBmvePhgKPaF+H1
w3VGzkK9TzU5NMU4Uz7sYKwxzVGgdOY7tCRTvxUmlKpbXvlrpiKWW4xHidkyyvfe
QJh15MhGvaqCcF2fOV+ofoQJMwsLX++IZdq+GCJpUYJNOomjm32+j1q+bT9mEKRP
dNBPMad0UhH2mTSMFnOz0NpCBRdez293F8ZcmRRMcegejEMuDcIASY2RslBCKdPh
A4yb6+RVGp6y5vFC1nrBKFeoo60rhKG46uSLYLVV3/90D/deqc46QFOceF9DR+IN
w6B8lT0YA057/mFO3md5yPU2yOn8lPq9mQ4Bk0Dhzne7qWTxfeAktUXvVYmZuxdk
/mWI2okw3UkzYLjyWlsFRazUSqLuT2QC8nXVeY5MflEXHL5r9MHcn66OhphDYSNx
SfMtfkHKbDgjybhJdPmzy0V6YqIg8Pog77GeS2JqkMqKyUVsi2ajSmpFBeoU9/ZL
Ep2hUldS96LODi+njWaCHyd7CND2y3cNy+4rsakIyFBy2M70mnJvOD/POj5XyvHD
9Clj71J5KKmjTTjZvuOhPqdVY9o31RLpMDzzQ5woabGU5OkNLb0NHQoxU/Z0D95/
+3IOBjv2Vu43tT7Wkgfb0oFcSQqGUzEBuGncRF0wSVyr8ayy4Dl2IVYo8jg4cJH0
MA/zbt+x8GHa0rf2rwmTjHGEJd6GojpM5L+lrnBFmN95AE2F3/ORReDCGjj9E9/0
4UJTU8c70DsM6Wu/zXHzL1zypIk2CoetqWYpG5wyxDhpi7zmj5Xi5WBMXdTbEldf
hOd0FxBJ8L9qCwupICfaXNhB2wOFL2y/nQUv80ge6sBGu7RxyNwzZuqx6dwzG4f4
EYC2KTPMJL71/4An+we0QpoEydoGM6e8FGCfvFmKRjjCE5IESegPtBvjXRMxFG3C
bQqWSWGTxljNYmXS9AmSV1YvPsJgXGhkjfVeGMlP/oaBI6DTeoP0SOTC74461kUb
xB7lswHH1SRnD2DyJ1n1BMo+gule9pviluOq65U5nK9pFCngEnoFVWLehzyWxODr
5Bmm+7O5qn0PEZWcv0lItLK466MlskeVCIDhsvAHngml80l3/r4sLbAWrcElqgK2
99b0me5TMNDaqTgSUFShRC7BqdiTYCWUbfUBANfpEcbJT6CeL1xwVDqHPJZkRj+C
ZiMuvr6IAsgQB86IRCC0meU7dagS0EThRxH6VbjyE+yTNhGUt6gz1Yvl1xobC+cd
7uQPa5Tf1C0ngXR1MYv24DTxNeN0SkiIxted0dzjqIfHklrX0Oocqzl1ejlsh4Wl
wBPEnevn/CTxBZshNNmoOuZrWCo7FLmAJ5fCB1RO+M2RA+YMaS7v6HlZwonyVXW0
/3KMmaDh1U/7t90vCuW0JrYhV2lEA2SDAv8Ik522yyWOi+cYyWc0Yk3jnsC8oZkA
UZ/4UE1gGeNOE1sRiEE1u2cUDuSNucAy61YONMwsJbO77tOFykGAR6gCCJhFeEXC
Rd1XC7aTNElYTgNF71tlMjpeK8EiETrpS0E7aDbe00vxglCzDC8ZytsZfbG5bZxX
52AfZDGTBzWVaeVN10SzHhE5SJYXIDjPDKqxvmErPgSBkFuyVhxMC3nDEgtcGUo0
gEcMu6TL06We+y/JWBK9bHIe+sBx4/Rlel8dkI9Hm445eKp9bAoFcCg4YRmBJcsT
/0P6nfFNo05MNz8sJFmsyoT/x2x+ylY2sKmTNLXxSTnNELtpQXa4C3IaP4io80bb
pruMK5pTl0jQRYuX8rgGbvpwQq6a7Zr+KFtNgy5pR8sJEtPgt1i2S/jdxzGvPCJU
LOAxKVhIorZTgwrnEaxCxo1B/HfiF6bA0QvwL+WGiabKFL+bE91NuSxEQUHJVfwX
k8oaCVydep/CLBeudR89kPbWuA7kDhd8Snrnxd/rPQkTjzg2tYFMdSsaDGrrHXjp
ZNXCa/OHuBnqnRMZXWt2mz89FpYSNwwVdQz8RSCS1kNyLOHDKekdBqb72IcSXWVQ
gj17p8y7XGLnsX8B96ZUzyZ5DUVLe5MbhRUn/3ECI+dyJ8paNXK6tFbhhU9808Te
0Vq4qMJ2fVdldGt6rI7Yf7HbzVm2jhllwyg7aujOCPsYIWbf1yvyBvxLfhcj7OoG
Od08SRevXiYvegPstuKGnQngy+bMBQwUcnv/MYKVxKZINR+SofO0/GGxk9yeAYex
/G94RQXOQoUT8jGGuXK4IEKOOWudTnq5btbQFSsxR2kkKTcZfT90T9+RZSeU8iub
ouR2LJAbSRV4Raw/WeUy13rRa1uc7FmbZck0LzPRQ+JmBnt6ROzs4pzwiRGS6OXR
V5rJtrAXTw5BWmMiIfHM4KHD6D03OxXHRqfZWQQD/ZUyyTcwRf7S+aot2UhEEGjD
1bgpmYlLmXNwwtTiL1YjE/z7+YMe4oraydoVU+5raPVdyw39qsKntAvIfwWhyz2V
LnaI+mEcMoB/Yn4rnmndbhgxmf/9Dh0SWgtB7spRXemvNCHpGty+tkE2Dez/mKzx
T/tjlTQBUICbExS7xKjWDIcjcwnvQ56zlsmrY5hghMmCEeaUfCtfy3KWA1nz+GZd
lYcVWl8zq456/oComgZg20w9OnLB+yhfEaqU0Qh/WT4rxzbsYU65ZBvAz3iv/nEv
IaI0+Af4SRFNKoGWcOgPQVFgpBIb0EZeq0j1nczi/5AQdDHccVWRPoLIFUSGQrpd
xhVAICJTsiGNzP3Otat58cj9hIIVSKKn/L7vj6wvVUfBs5iRU43t9TykKBLCuc31
N9wFp7FslHftkndH39nAQsVIWHd7sgvElvynCyHfVfCagNWlkjFbYpOJQc+pHjTX
+lOv6NL1ElOsR1BQEC5OywTBq4KGybPPnqONcU0fa1LjonRX5SmGwzPwGF1YLdGd
ugGr6HLfNv8KA2gzzXfAmFlwsx5vrgCPRSKjQnkNqwYopo6/8vrq+mHvI4oenplw
fMwSvBO5wwurmC/uSbXWjn+HzxZxVhRaTGNn6lv2auUBcz+pYd1r7nqNh1AqSbVQ
C3M0h6NstM5iXA0rF68O9XuotQ9Mdjmjw0m8v9eBQilU20JZYfUJ/C/qCdlt+N0A
koQYj6inzH/UL5G/t5yUeDTYEilQsBZw5s5tPnUnp+TLkrd4xrEBX+a3WPt4p06X
cRMp5I6SIiL+n6TDm5j7QeHEudP3xdbQ1CJH4pHPR8PB2PVatDd9F5K71ckuuSE4
zyTtt+KW4FUzjlrPDHz8W3BxvXm6MjGaR2ObETZXAWxdhtbxpwCko42z0vSSItkK
e+BQqi4buKdkwujwFm3qEIDprd8uhl/1diYOmn7mOqeAClF+kZ1GOy5fUlJeIOnE
mz6Jm6u4WBsamqHl1p+MmuukuxSH5O3P9MIJq+td9sT6JMTNDGiuFodDOXG3daUt
FfCsd89RzkWEakLybcDmEa4Q9CFSKuR+0pmGixBlpY4SVzJtQXdot8XdLKYTNQ5I
74IEco8E2aBC/dFUuPSddXJtO+jzxg5I5BSUUoietzAB/FKJIDIaBSn8EVahj0qD
2BWmgr/Y2gfHviOhvT6RluWndvuAcu49Q1HuJBg2NknIaGBxI7cULoXXh02guB9H
t+xrT3Lms/8bMftWEzgfEimV3YiPTVobdOZEo1ZzUmKYR0NYGlLVJ6N7p00SNtwX
My4IH8iY8Ie5/8k8cN5fiSOO6uNp1GiEUXLoWg4i+Q+urQU86ZHDB4wpZyqfZ0OR
RSZEA8fy5jDMTxRVMJwh0lnUe9NymB9TgNCRs7Id4OSxQc4HjCtpRd0T20LHY87W
Avr/4/RI9VIgJ/WviMGFCVXHpMq4H6Q45yxa+bAL21m91KhjCss97gqjqDqDLgPC
9nsqcTauOu7lJ7J0mJ3CXOv0iHU7Gbn4+lwH06NjV751hli6OAb0trII1v+C6HcU
NOq4Yo/5xsU6Q2Z+Fnvacrv5qBpejtAiysEws1ZQgjIp1Xoft0Tk2DxATDt9A9Id
YsvgCLSWrnsdXK5VzNBmrvNWrsRcCuCr486hVj3ki81YQ7EkutfEwsmjBLJH9cxB
LqJHJ5fRT59MEJbrNx7nlEZBlP7REXZI3TrfWqA40soaPd/WX1XgFKopTClO9kh4
KfbzL6ZC0hHbc51fJI0IQkmxrpYYS7z02eznVWVwr5hseCXJl3DmpdWnhuvnCduK
WVXyZ2H08abtfRk5RoTomQshs0lpBnH7B8KDTI0dxd45Vp74nptRHn+P/U+oacmY
9NXlbLy4oZ8xQfCDAsG1jF/l63L9lTMAr4CWQSRJlVWGQjEqdFLPbRyrM+SCy/c7
5IgHqV2IhFmxJ7kjgYl1SNcL7GS07x+oLeoED7iIZhGj+lQ3wTa85SYYucptqCY+
Ig/oC4VDyEh/Aec6uirQTiLOeRef3F4qa1fdMI6JcKpa7JfjxZiZLlbyJ/omV1ry
yfTHURpSMU5fMgEi6UEFqrvqz/B0jJkMqXZkNnvfD8rPQDaUFSiidscJZDLvsRYy
Qars3WQvYX3bvMR7k4bbEbRlZ0vA9GWEZEtSmu4N7UD3T/u3uE4o7JlpZUZlyWQp
550m0rU0j8t4K+mpz/+WHYJvOFkvV2xp0Xltq4IXXml82pwIcbVkEwMbUiqKzUzl
K7BZjwx65sCc8cZuqNlVKmdikVOgILQMQgWFLg/T6vvUbkgzvGwwc6hxr4OHpIgP
NbqsgWvYQyTdkx6j3WRCtNz4ZBEGRUQLZl4hKdjDiWflZsYSiPKhGmMDfD9kRbsm
dlN36Yqe7mR5cjNEAHNsI5C5G9Y3GnSuquoG40mZ7uq4ZC2C1OdrkqoFwQqRo3p7
WfxZpP+jWO16P7Zs92lG/GIIuCTiKQGkAuKbf++soLriJWdBt9e5JJCOYTuXiIKV
JQ/HeIiO4Ad8iQvK9W0s4fqL6oPVCrS0Rul4WXGyqYblCEQqNjVNmTpClTMl9l+O
O33S6QEqjhfQcx2lfNhyZTd46VC0OsA0rJp74iVLBmqOtn4lvWQtt52H5vh8Loi2
iKJqIW1z/C0W/pXadAmj9A6xLOPzRYoTe+Eu9EgPjEsTnncYm1hqu95NnxXDqP5Y
vPlTRbhtZAO3hLK2SR4sHI06/wIcLNDDAVAkdgVmEqg5UZ4aaM6oQBolhu4G+B+4
uGjnO7kWLACbhmxiRrYzphZbPe1NWmFp6BspJzSvDsSvuoA43f9gAC0s/GJRtIKY
62reSKz17dRxaRMSrwgroekoe/yfD0rGR3nhEp34dXqXup09WZo7sOXU5tNfSv7C
kj7ThOcLNki5qZNDjpI8jUMOtjurLHfg3oMRIIwcgjTEb8wYsbOKudRS9Mjwa8/Y
gD9AvhLmSaXv3S+fp/3nngjm5XmECjRxYDnOiBtvjHvZFTuMw7ljki05c8geWkhD
c0oaO/msqU1+zjXl1cqITG3+AX8StgjQV5mqdPP1V84XQWk1jcrvqkuJ0gTiaH1J
LtmRg6ejTRuHVvT608H8kOk9TFVy50PxtYokDH7JsfQtyGPv7xj7FMvrQ8KHC9N5
6sa/4xzHUH/pR4XUMSPdiH2xin7OWgkM+UY1a2LismUcZgtkHVVlSDGDr+0ANooW
rQA6andOkZa/PKQ2TrZ1SkLqTCimw8r2+6LyWsH96VhNFIGx9ZbDNj9glTIrmeM0
Ef3SSqZb7tKBWS+OUEGMpza0gRMcv1nVkHCX+KrkMTf2fIHflhWrLrhB+DOCWYSe
KxKkS0UKIt+EFXUhjEriGENrK3pkyqu+vMCNk/KYclpbSLdDTwQCUV82Ii7qEnBM
gJyWIa3r7sfms45+COcwTE99lv3JAhKPhPLsvAouttc1zgI+B9AHZWZ2ke6KQ6/1
m6h/jtrot3EhK6M2H3bBKwzrvaIr8IW9SSjmDwdO6LzObctdDg/AA6ZYMQtRaq3d
KrvsEwc2uFESJw/8inwCqqR5FHMzKfahWLI8Luch6zLRmRriY7LVyiksMY9HJ61Z
5PiUjaLwP/X1lg38dA5iH44InN58bZOFWxFEf7WBGvxvWk4LOEm0NcAHSEDAt06g
C7HbI9II0fKXPuRQRLuMLNQvwaWhgdRKsJyTLwQdyAcn3oAqT/tF7jGl075eFkA2
X5evKlaLjKsIq12tqpI5pIKCHhKukKo/C6O1RWrNrhU4AufyjhM+Abgwyj9v68CF
kvB/VGoSoJboEybTTBTSh3Ac8/uZjGW6s3ya37zjMRqqSDpEHVfnL1CIoBCDbf9J
pM4+xoBx3jJvUJ4fDmjPBeImXMMmxictVLIsxYO6vQv6JfNJHASEjbZYgrcn8jQS
c32Z3sVZMarZVGbP9TuRxNQ9adYFzojS7OVYHNkLiFBFgApyGrmPNscuqo0QaF/d
8wZ5x2PqZ3L7mX1yFihZw4ofKV+QQClVZ4V3KE9FCNPQ5b5dmLptLBP5YAPtn1wp
SGYYGH2TU1ffiAJ56B+KdFI9EYjE1JN2jjvjOKbHG9Enp05+tldYE+fbJ+N1W7AN
qiY6LxgyY5ohJsOObmTkAUwil/PCyl1JcA0o4WACn5lwZrsjBe7z4Uy92um6dIqy
AhcOJmNM8JhWacGJ1RU657+OigyIFbVqPuKU/W3NN2i6IyyQtvjzrR/KeCxWUMpG
Lo0ZhiVQhicDrFu7Aohsd4biCoZltt2M26Xs//EwmfDh7Zn7Za/KxTXeJbsyjUPl
0dXgobqmTcI6H0kH1Fpc1ex/ctOridSHQzY2T6uExiOTZVWvuaLue9z0sdBIWF7i
/kuaQ1IaerRJx7/kN9dOwtU3MApF68ULkFUkJsoqacy+AsUPUpS81QEI2vUEjNxB
XAD+I75gy9zptRCH313blDJ2pdwDdvzcgfAl+qmLbsRhzzseJjlIczbqcjXezWtQ
bQfD4G8DbLQIT8N5uN4SNYI/10wsSNSikLSh756IV80Xjo2grvbMTrEMY+2tWAr1
OCK6LWoDoEuGJGQL6XNHVDK/Pa1/7gfIwwPv8wS1wt3cpHe7qk7rDR7x3sASwI19
R7yZAiYO9xWhkWdeuIyU0932/K4C2lDHwqQOQ+OpG9EdvnMcmZhNS+a3wgR+Zc1/
2jlRyg/AsSdMjMlY5GI0VRKyPudB/VLXLPbrB6H36u/QsJtIZbSqfoeaQYlrRKJC
IBtIWBj0fK39trvb5BfpOlVbbi+dfQXtqAYUcOUJjihAgwAwQwKeTQ/JDQHu1IXo
DjgCjldDPYSyyo4FlebFcWYS9Hpz1w8pgEUcMTe5cNVGFhIiQ6tsLKNB2ZL8RqWG
2w+ccNeuwVapGl93rRvWivrgOuY70VVuyO07IihnrmMutqOrvS7RfOhFHwaKegq9
SXNWvKkAnhmmW1MnyBoXqPuD5KqTGLy4eUaVxeqA5rmFIJ4mhZaLadt8ZQI5gteW
qX9g9+Ef0HovKrFyUOQhpGqNjkFG4eetY1OTcNAAEsZK0Yn9UnRaK2VwfdsB21xp
pk2LCtRewQZmW5n68Ty/4TWhl5KMI5nPRCcyazyci9rBIT6CsNUX7J2Rqm4eOhnn
GNtO9tl5LjOKIBzqJ2Pb12ckuAB55S+HbAnqUSgGo+xzGmu7ejP3ZcKBvrLTcl/s
63H27mMAVDxsi9530UH1qqQSoYC8zs/Zh47KONI+y9ekrcckyZXH3pJnGXqR8nFo
K3cX8yOEOrLrCj4uZ/YB3MLe/aEzc6NtdAuXb3G1OPQwd6ej2A+A/bnrBkjq8w0Z
hCc0D7zWoWR2BEgHsNaRgR9j30E9L5zNKAWjnjPMh5DXr+nDtt7veAYpMYil9A0H
2+3SodOA7AgTgNGoKFYCrozFpE4CgEF1Uga6UPwLi7z/fhg8Ns4x11bme7nWId1O
qtG1NHfin6r0Majp8mzDq9gLpipB313l/5Kd6BIEyOWXXUVST+NtAJHYb4BcdYya
wkQHC8CoAMTRC6aE7VoWSNcBHFh8spMLcUVuz8pGMfLtDn+sg3P2rIHa3LY0jG3U
PoIXAzJIebNqZsNZdQBLXhUBFutQkMQZqd08mvbQK478ncgyDgXouJojx41iwDby
Is4pyV6eCfeqGvhgblBH4MFZKrGIiejWhbdfz2mPtk6gyoui8d6unQjp0d5uzAp9
6vnhxVzrr9HAc8WB4wnt5NOgSZ4ZE4O99+RAfilp/XoQDmPeyZTooo0kbdv4zs6z
2GtrWoH1tK0OqoSifaVPawhOFq2VaVY7VjiaY5DeVKtEbSJJLSi3DXfiQFwkISjd
NJRldjSYct78+kL0FCF+g1Ws9r3E3xE/PF5aExF2jtsmMy7AsGhJKB4xg+dClSK/
ruBHJcJq7jmd79R+Ig+1cp33B11RdHrYyf6TXTqzkz2GcTuqSmCayrZWubKdo2VO
+ny2ok7ejRnbo6kPov9W/z4SyCSxIZfpUZ64Gt8gLMucjHFH/wTP9Nq4yjJjpR/v
0sH1Ba3puakk9YMmFBrNqedneIbau/4OOviOn0pObm7nSXMCEkox3kP1NqL7ZiTy
IFJ5PqouiP0E8bLFnajOiMpVNmCBmmadwH7Qx99DPgGb+3IZS4ivUd5M+d45v7p0
4yaymV+wa65Asns2rwYMBBKWUJyF35HfZjs4mm4NGeELD5vItZbxgv+Httbyf6ej
HXPF8eB8kEyMBjzCVaMl0IDGozcAyafj0H9xXOAViows6JrHbmQYe8w7D8/+Yw+2
4qlooiGrbtbcreqV33naIlVT6dklOpNQDmavFRfPHXyjEfmVTuWTa61kO6FmqABB
IEc5PRt9zUwSeo37GDqzwuC7MCWy+Gc53YTWt6znzfekFFw/iIYr0/AqwnbDlDJJ
EXpRsGIANWn9pkZ2P/Xdc/CnLKVKsGerg4TqpixXYbQsNnvrSLa+cerKmkS5krW6
oCjT/efelecxMT6qbFE7rm8Tji1gFExqBIB2kIk7+rB3nCWNG/tlweMV3zfc3PWa
oFLYzjQwlHAa0gj2CiLUozYSyQuQ05xlXFy7+m/8ZW1ye7ehqTlHgkXbp5hiNQNL
vdVylBleXPmJeivLPINYaOFoC6cugO8gh+84mgo0tVwHPciCmXxOKVr8hVUDKhlE
JlVv3e3m6rGudd07kRm9PgkIaX5Td03eEO/uH/eYhAwFfqIUbxegbwnqBlrG5ygj
d8FT1S2/jr0/1blUsv7FKJahXyXkq/9nF9MYNQmJpz/sVlp7vkYaf8MLuVaYbjA5
2AVWVYVLT+mBu8hnQoLqjh+7DSiXEut52mej+6uaLWN7RAcxBWNbwBfvexmvPWsM
oDz/SyfhOds/MBk45rTlamBg0IUvZSNL/dYQceMjD6QPvF10mwDB/q0Atrafut/9
wD7eeK6AmLN66z+AXlQOo2mDL1UHvdBXREu5n5iUMY5l9aXhv7g/Acvz6cOxe3eR
9zVRvvVxQujeh6FhlKHcU0zpjeeN2NAvqY9jp7eDn1wzbdF5yvmWwLAe/3c+9bAI
QCEgLN04zrEaN/yHiR5zyg/lVu/pKG29ghIk6/Q3443BF8fahygD1Jbx4IbKEKbN
G888ts2SYAULoe2Nl5hjgfcLzsjsexYXrx0r/lyy5PVOQlbSSJLw+AHMY0KN+aAs
morLJVJzy9GYkCPJ8lKLzVw1LfMxxmadBIajRjyzI+DvoIJPg/FbC34db4l/tahV
qaf8tDDH8Dx/fAxppMTo1yNXREzYBKDC+MG75P/23XoNcUX9IN9sVXRgw3U2AO7k
H4/0dYARN6riSdsx14HTaukUu2ejUwIYyEBsbpUhaOIMxqGJerQ6FFa9ikXgznu1
Vccuuwgiwx/oM6ZeyrE32rZjcnwKB7rFdyAXg+2hu2wh9XIud9DK2neoqlnTdi81
b6QlbAhCnx8aJPZCSKGNk2xiG/+Nj2mXD0HBedGJsjQhAeytDMjRcDx4EEawJqMT
7ctrZeEk8S6VQz7PnlVtzlmp7b1/XY371DOwskZyEENa22M3k0CedKK2U/Q+r3sx
pBb7UWzX4gWWQudbr8Ni88pAe/0tjvpWRJoFpeZF40Uq1jb72jbA7DV3yiQOyYId
OAb25qjkNWRei3NzTzGzf86pCXrPDFMDEslypEvCSmvFv5Vw7Pef7IumEGJz2bZe
xe5lRXWRR5lk+4X+zktLMEza2mSd3LHlU4/ngez57l6ewVCHVxdcxl2PAAq5HkGx
3AAHi8o9lNaPiTJl38Dh/dMdcOsp2X7SPM3HSom+Gb3boDSpllnztr8PwEFOXHYf
f6PWcR8BOyh6vhv94ls0AfBlZtp6onv3G6rQeKjC9wTbIQiT7N6KdfFAPgDM0k0B
3yYDkxE8188bRz0JczgpkP5ZCncqnpm8BJZBrEGO9bu5gnT56Hrm6GQO3yk4CvuU
jt+aF58pIkj0paqO9h2R9lHK/9f0AcTn5iEiAYEvZmupdpGY+pKejpfR8hhcR8tU
ZtWQGmZwO8ZN53WcyG4czFVnGo06WXlYWQwhkiLvdWz1kAJIxIA6HuCvYNaoTq1T
7HUUV23elo3PXr6Ojh/wvmDJuRvvcIGdGkefpTHAnkiAumzB2qsqZuOBefw8Jfny
nqvLArm9sqkw8bVDxqtDAIvQGu+lFbzLBcfvrc67HZpyCzOIylFXbBTYlm+j44UG
vp+fGomsLoqMivvfYz3x5DHv8CyzXBToJaiRAnGtZ1tjbRQBHLBX4Cx+0mqauaPC
PwTm8+oAa9gxiPDueHyUX+/ke+Pd3VOBPZ17kTCQO/Gku+uLdym4cbdGRJyzo7yy
E1sMRmjXuHYopy3RhWED/X3p+hz/1Pgo2fJvqVbm7nCFzGAgC0bv69nkHUQEPFd3
yihENCNYAYQ0Rx01cXgtDd4tu4Kw6n/a+LWSiK1UVpBFOv/ViXdKFzfpDxlMjuMB
Drg0ksKCdO67rZNf9MkqNUo4Bqgsv5N+9tEzRNweF+NAE7LjaCF8VTde4xz8x/b/
2i4rlchdHoLE1EhrVgdPovP1cfbmMNuXwZvw+OgyJxyP8hvRth0bRHipY7SpFJdV
U5mXtlR+koBS8PJpytJdi9V9CFN4pMKqXQ9AuvNaW7+5fLNBIR0L2AitUqvqehq0
rwUhSZHAaiT57uMJJl3nuN2tEof5jnGnK6gV6XZDZNOultWnmazs2afI0y7JN7Oj
8TfKxKmaP/9s3+igclQnL1N/6PHSDQnXvQItDy0CPj6T5r8jAhhrGsoJh2S/tDQJ
RYgSF6IFC9ORdQEeli3BFgM+Yf1DiykFXaKZbsbHAaIppVYhte2d4Y8f6NkCS3os
cGYXBD41aTpfXTsvr50vrFJgJQaUqbN7FEgK/t0V8YFGzFerUpTNGExNS+XZ/u2/
VH9+2hY6N8n03oUCSCjXRgntEjkAO/T8s0zqO9gHNyHgFtIUyId5rAbVTdZBbwoM
IwjOGklMMoFwz4L3jI6ogwIOovvhAEgvpTakCoIGnH00GF7m9yJLCFp7hMKZo1Wd
uHp184wON+bmHChmxvf/OtH7qwrAhjRcOK7S1aV9wu9dyWXFEQasyuXraC+MdFo8
yUOtmiGj9ae/k70yLhw0cyBUvQlDrCl4E+gB2MjXn0AcANpGQPh2Db8w3BNCy6RH
xru1tfpbwk2/Sz4oubwnoWzd3wNxUvn9VBo5yjriDqUgUuJ6h8MlAjRDJ6lEkS4Z
N3WKWk3h9TpnpMxKEwSNGyP5ErEIk0YCZptNQUZUkKz9TZcZTAhsBlT0Xj0e5+U0
IJGTuvVbMfrgZlHkdvX+GUQPDPvRPCmwpDvmnQVvWQ9OPZE7/za0wJTjkF6NSUqI
rQaN7xr/mZHebOb5hyNS8d9Cc8D2MtPgijbteJvh9qtzlHNLOmnkxbI+qBqFPVfA
7O5wZ6Zf/DDzTaFMrA1bp+YALQejYB4tIb7nY32lAVvBrCxJx742xdL7aj2wNaA0
ywlFUBlwgTHfSLclvGXLPuyH4YwFQ9cD6sbMLcwePzuJmz4xcRwBN0GrRm1DVCKz
pJ+PzGRNLDMdF63y0CWnCGzk9E9wWDPLFaBltSZbWrUVTVPcV6JEQtXTlzEbDGEC
8Lc0I3i/MfLYGb7XyG8HttEh6upli9Ujx2Zf2+rOVxn0qmZQ9DFFPcDrfAmuRuVx
JdlhJOy/YC7nyQ4cq/H6ANpICtn2L2DT0p4ia0IYvM3yQkrks0LHSXebkDlSZZR1
982kUlAdiC0KkaGG5X2mu/KyMBfk9AlOAMPLrJ6pyQ3hb9IFqee4gMa44zHwxm+j
j8J3NmwFhbbVHkbqbBFPjQThPVEUlEkUB3sUDaDvnhXbpBcGGWmv8gDxyyqDOAZI
NelspPOMjphlMEJCenKxcrORRYOqtRqSTFWELK2WbkbnF0ZQjJM3ImI6yJxCBHUp
J7CTe5CwL32P+GzL0PW80ZU7eAQItd0nb6qhla/78dYBKGFB0hh3Pj9THCXSxV+p
PRYpas1/Oy6RNFwyEa4KvQ0k70rI7XSowXjcGQzT1S2F86KT07EH0E5F1YZcC650
YqXUT7xMkNfpbHciN8Acg3SIgNWJIVgYyjsH7aEMaiKIjYEqz86i85slod1YW9bV
xSA6AUZeCvM8zw9FWxAHVqpDFQgwS1YRIckSwAsGTPWDlMv1n27JycfJU/L7PyLa
mT+6xye/yg6wsMuD/HzRpJ1m3P5zPzyWr8RVwMsU1wFNQTOs90ALzo4GMFf8xN3V
O1VwtVOIfozcK0wc2jES07sM5g/GvpEqdIr+LudoUglrFMFk+5FEjpRHhII2/bBu
KcXIy3FoIOXYpnyQZok4tRqYjq/LIIZ8dJhMLrJ94I4CjrgObN+jhgdpGMiR4NdZ
nunO+gWvwgJJW/EoherlADR3L/YVxMfLyytHaQxuRH2nGfBB4yA7kOyXuqaq21Rp
FcqKZGR9h4uuZ/Ipth/aedq1UBTATMFcyLFQcEV4X4rAbi4XbLUbR6LHRn3Er58N
zCkq1SEt2RqadWlksZeJDe85cJaN3BKbadaM/Yaqt7WmIEdD66MjfxHeeqhOCykA
W30jc/c1J0IthwZFqu1jDHaFU1LMohFTqtu2jynHcSxRBPOfscYHmuoNL9ubQH9e
ezxlOsjrdEBlrqCbCn0SM1CiSnmS8qWzdtLujjF0b0+KMoF9IlW7dpJozKdgWiV8
40PzYE37DqKet3XymgbCtJGKRHd+FOR6DlI/HbSmwxhauI1LyuxcesF5g9jh2QH7
Y00l5Pt5kRlkLG9ccr69FQtkiq17daFhje5Q3G0nmLGI4hZAhO9hzESqYFmHKFLs
ItMwyJLnYKKOCPTTR2epEbZ/d2as7RkhbdzU+qI1glo0EArIRNlRP8VMIx9Fwhk0
X1rngOil+hTj474Hws/XxyzAA+sIh0Z/zPxwdgH/MF7Ju9ZxoRHAjdqaxu3YJacJ
Je9vzTiCp4VnN88LP3a/pHi01a/88zRMGtXllKDukcNAUtmf5McklH0WkO51gFr7
UzLXNNhhfkKZwxN9kpLes8ElFPs0CC7BCgnyicQ/CNEMKmHU/w18sfd7UuUXZour
yn+Rd0WVCxsVN5N6kAqxmhE3nWMIfGoBznifHOiicn14Ue59lhSOwqOYcw72qboo
zXCFnxw/y+vKfsm9E2YhqZQdbIFvFQfChqqpyzo2RuN4CuMoqMhQL8gHgOs1UOq3
cP2hVwiGyQx3OmOZK3lFWuRmP9+qtFSmHbs/YbwjRm+FL8FPRtDTFVazW6FrA+P4
y2XbjFtFMbEeG4QNLjxK40suji31eqKxggTy+8oPEav3/+nlNeMEzQ5yY1BKvkDI
m1AaNgjxtfSJCGgf2sgHy92tw5iIqpY6RH3pNJq/KZbg1AtVjxfn4lUCeczHT25A
TKvGUdRRcK07hm+RqWl0HQblBLmHAFULXL3pT/fTZ+8mFw908UwgkjkQ3R9Gs+k3
PYq0oDYAahCoPLituUfUBli7UDU932LZIQ4djTLEibOP09yKyN+7AX2HMK2uA1vG
uZwxn0VvGMAAdtBY5q/t7Zx5hh7Ut2ludtaqgdSmzSLRagGYprE6Y9FSLVKZBdg+
VtV7Ukr58tMjbWO6ulomHuP0BMnQ+y0lM/oQznqExz9G2zj6ppK6ioJHfyVna4uJ
/wqDHAt3wIhky2U3a7qCyVHXv5sdxYV6TP37r7e+9d6AaXHo+PYx9Zcwsm0kFaY7
yJw+ToepbvUZYtnspHvjdOtsOjfxNLaoZVGNCmyE4NpxYMIHPCqiw0Dqimp5gv6+
CUknqOL+4ywCtHwNWYqTDsvYghVsXd/enP7pIfX0jtk2uZfV7hov2uaU/dcYH1Nf
CG3jZ5h6y/Txj4zR/UPlLv+y4cX86h5mCY5NhVNee/I2xdIq6p5LJzK9IVk2HDmn
uJX/Z1MyYZzf4gmK2MbpZF2uxjiA50o2qC+mnzFSe4LKihx3hpWtyXFjhB/f7FeT
x0d8iA8SAF+HFxPC2Hae06qJEdDlH3R0SwvTh6Sci1DK3KSCdLiQj7rqhixz1xiO
rBejhtTANPIqnB9ahI/EkksWj3FbOgBwIYKUi0YkHt1QMWY/e6WAD01q8DQ13LQD
F+LWRYPjw6hNZr6AxAJzVjmMvgI6pfUIR+qKGegornEKQXpXvdW+HBVAI1zL6cWa
T6SzzHtABto7vE9max7B9hQhVICzovpL3nHmaWIwB2Vqp2h4aA91Is+llPf5krWs
BRi3HtUwntc/FXlnwGmBUjpFp7AxGx67l2jVY5eBbSqiOJwIzmSkNpxMPkEGrdM0
caujNff83hqLFFXZXovZvRlY+ZUtRapw4DXQITMqqlSF063028AXu05Vto+ZhG9s
QZm5bvU6mgaqwy/zcyoyqruFrFWGihY9JPyPRJxK6/25y/tzBiPxKmw8S+e8xp92
316AQ69AVhYX3tT2cMUXuc4q3iz8/jJEopTtu8UNnRjIjflzhaHX+ZX3rr24OQuB
ubVJCsyCkS2jEme9aoWNq2sEiEieif5mcYmCDyQE0gKBiISduZflwqWau+5BqWuD
LA7OJLk+UPtMIehMyJn5kplapVre+qgAtuaev8Pu4fhybfKJfr7j48RzC8pfKAN4
41R4JGJnyAPNhOIRyZWJlXcLjXc+++ogkk2kaxfiXav6nbXneD4zhZSbJon12wev
Gj5a6vqjC9A/CJEXigs81A+9tE0jqcySGnmSmR0H4p2sNouOtyLp001FpewBIvc/
ZfrgFp+hZFogac3xwZj8usiGw9nRKZ3fGRzB2FSaZgoW7QABKFO8LFJJRKjS8JAG
ZOeKRAubModrwrIH7NuqneZadtkaPMjzHo0g9RGhOjYbue958vS3ySG+LXy2/8hG
gLs32zJnXokpGWYPs/aC+VGC/E+1O9IiI9QgNexK7f9OD87vxfI8BP8c3HpJffzl
0ZMgpYHi2G3MdletW8maeQOWFoFk/64Pca8N+6p/hCtbYkFbM51DGHxlXJGKKh9a
WVldoOD4gOfEbvrPAGFv2714VpKC5YLJoe/8i1dofN80D6mUKApFrkftZDMWVyn2
T09+fSqhzerIJtvvW3oHutu/fCeYsvKVQXD6L3yfLe5Df0QwnFzEfw3Km3PDnq8o
ETdRQQzBW4kAatosnb/grqfPpg2RDn6pVq1rrJZVERsvhRm+74AAkjZ35M5Q/FiZ
wgAx4koUjYGPQy7/Gka4CX1j1+tFB3YKi7Jurg6+CAjI3qb/U77RNh5QstwC7cnP
sM31MlPu9+ZnIIyeLcrkeW3ZKd23r+h1VcbzUDoVwrgtfFhAPJ/+6sQh4eWxtzNE
4C4N+ZEGJsslOfL2a/MA+tlY9giKS4UabfA0lYF9NdFzqXY9n33xeQE7xDB/R3SV
jaKSgQaFGqFB6N2b8KDQhxE9YFemxDNtEswMNUK9oZjmd9nSKxjdR/LIbmmoMN0d
OGQv1SYPtOyMhJ6tOYeuWGxn4u3UklPtkbwH6Iwv7K27vkUPHS5MA6zpG/4inIKf
9/5zcXlGnN+DZYPAaxBWSUvZRpugBXGGBDlphY/SPVb5c5FWUHQIFGe8QK/4M10g
+fc19vAGExtCLvUAW26X0w42rpy74RVDxW+Hm1+iCcX/k5NF3x4UG8NDzrV7Qgny
N1uHLRSu1Zu+WDH8epj23EEen0DZ9HAuwIHeNayPjo7Je+zXe0C5smWyV/GQHuAh
t7WNqcb9fu8f9i1OOtyDssVSKOeMhhSd7E23EJZf8tEWMXJJTnUCFp1GZ4jn7zIc
/lhVv42Rljb27u67Mswlpz3oEc6ynlstLQe15xpaWyghjyFd4WJYraRgnzSyqpPl
tIWX5/Dp0tK4fzhE7axCp4fTCAJUwRxpXEJ0ogLHKFz9u2gnJdo23OWSHbyrYHZP
3ksXSEWbFjukB2obpfaukRPcncKRPHSVxMTgVOFyPxIUZyqj8ujH0QCADAWNV8Pd
WK4LautGTbRPIkCdIsP35IfEEvN4wHB0NC4OWAUrlDIn5P3HTIkwqxpLxsU4Moqr
B6UbT2H4QWhlswFteDU17NrhUOvBSz8cUVE+hXX2poGzRQDbELz0xyBX3gWBf4T9
Fu+EE+mpZBMy/iOwleIzDTLS72vaqOfgUXBKtfbp2quwmsplCJrUsmxHk74eOg5x
UVTyPe2isNiN7O2Kdiw6rUr74CXkPZBojj+jVZLzUClR/x7sXtAl+OX69e2R5C5z
SvFHByQu6hfHhQ09r66nagcXBSs/Y9AA+MrKX3322vO04+kHd9DTw1hzUVwUOUfG
fOtUq0DR1zNGsMbi6/vketQPNE5KDLEUpiw8lfcZzG4rdDzmfGODO1ucatinwMVy
wZBFLwy1xvawjPbcamVJFW8lZCgnvt2hiqn2tAWF2oqUYpVDSHXsq9MGIOe+Rgec
/ZY/tghUZvsI0gj+HvmbVHwjR7EvOzRm6BIHbP5+PTUlhetzayK0JjS8m5Ihq6xc
fD6cACK8zGki0GcLn60v3Sxvtf3uOSElTYILW9VaM/3NnC1OZDpwkxUFroJIIDkt
QlcIXKJx8twwItgW+7XQ+jhKlhqrERiG87NjN4kvRd7jQw03hYklaGXB6poI40hk
JV/+zso4RFVIJbtLfed7t9mtn8NQ87xSndQUMXW/F4rnRZAzmb7caTBz+FejX6II
YGltlftO+yCeNEe5xDUqFZ6HOXZVL7edzE4WRrB2AIn3tEBxeIIMbPAYr1tEODP/
6sAfF3b9d2QYmhVe49uqA3rl9KEzLwPB4tCVvJpsG4DnWIq4fMaAEEB6ketzWEj9
FyqIYf7SelfrpB/3y7Rvz4M0zkNP8BX/BBYdnCWaYrTvap4zZFwMFHogNfvlXpcu
8kunoxXlyM1+HSTG3S9sv1khVYdqMu12bkifJ0JWotBzMucT3Nik1tNd2JdMrYRS
/+7olaudCiII1dYukNSI3Beu0Hzon2Vr5/yRtg5U5W65oS7DsCmSWqwMRdHlvXIV
lma0sL5xS0SUT7uxTZPtoSS9QwnKQEEBlCxoVrol9BlXYjKaoPK2tCzxUbhFKnZb
Qenv7UPzLiZlz9iVSgwRddDz0223gX4UOYVPf9iAU+ndvVSOlhCuDFNAUjwLT3nN
78YqEFRBPA/cA3WOnCq1eSBlXsfQybc67XHBDyMublT6zzh7lbMHUlf3p30u0lor
dds6SI9YHHwZyMnjzwC5LvzeujlSgkkNnWw3Nly4QieH3i4zegQGeGit0h5SNbTb
vw6rPS/VXZz/k7EGCBRLXroF0ortaOoQFz8IPFh2u1wlfZx65DHwBXVvfpprMz0B
YHV3IjR6ETckQl2EX90mB08poaWTztf3sV5zP7hD5olD5QjZfn8ZXnW3c9/kQd9q
GUMTUy4NIBxR1CNOwBoEuve97aXRkTF4ZvSSusqwyKcqdKW7sw8qi98weLFUI1VT
THzYXEnoWO+iIOnqU044H2Yo7/51l9H2rISLjpcllxdaxeTCKvRcHx/j7ew6kWH8
bIZ+vtuVLkvJvwyeCNuPt6b0TIJ8DPtYWk8HBc2BTTabQ3GoC3kjoY2RFxXlOpMG
6/+hvEq1SI5qGFHwYoQgs58gwnzsRmZdZX/o06wtRtGbMFWKAAkqsIwzzSOD6iMJ
YoSjSb/46R+d1zW9amllw6GkcLY+wHQ++1wGNgAHjKilctuWWs2t5L6/sAPrWY9h
EgR+obw2VZsKtZJtuGuf87fcyKtx4WOojKNSIxvxC5TVuEqYZV6v4NtG2p4BD4wx
4xfKO/U6dlDuZ+yJ5rFH0P3C0l758CVL84yg2pX6s/xPrpewp35SeI00shWPceLj
rtxamVMn/z7HIzV1DquaF0sogiMpROut6ugqERtAjEyno8EtZNut44+msiIDFWN7
2tt4GcSfdJworbQMD1tEYL9HJiT24NNn3L080IUhh9xW/YFUSApkEbA/g4UEnPJX
QnhJCMAcfQlRPh7HcgLHAjjAGgVebfE0oBmmuSfTu7WtOd5Td6c5R1Hl5TKDC8Sd
hcRbovrX/Z6SP8u/tTBxXysR66l5Xu2vRxAX+UF7k5EsYj5at9CfzJaSr30lKo9C
OE9xbBEfhOubRzG2Ya6ckBxzn1hh8428jXLlKO42qAAbKnH/lhJCUSoIPFtt1Dcc
WHNXmn7il/6l4KmDiynCIAfRfhmhvbiVWJ2PLBqQTYA6Cywz0fO0qwwx/s2Cwbv/
gg4JGrcb/BgjtTsgn8VdQSeJgdwhXT6cL0X2FY4Cd6S+Jz+jS7nE1NHugOOJscPl
/LNNlVTJlVBj7rwUgmok0UJjxn5xcDgTNEz7viDCu0RMzG4p5dFpGRzp/0oQFLKJ
TH2jOFcszbtsEpH1G545hV8J6qcVWWoy/vtQXg/6YPZC0uavvNBQTLTVtdgRfOJ9
nV5XRcF2onFXxrSl295ieQprENI3+myMUw8ydlyM9JIT+Z2louzrRtF1UxIKiFWJ
iFmSwWg9x3TDh/Rs+b4eea1PJNyOdMQqnn4h2FU7zxLW1KmOa6dTGDwFbpbn/8hD
j/kMz1bKCOrn+oavo4F6PWR0RXsWzXCLKzUXQvl99Stc9hWaNNUcuZyZhf2uqhHM
fk6OiWILu+NI4IY567MruOUMa8q5zHaeGM3u/IkFHGz20pEWMzwME0iOIkXHBxFJ
/g5CX7BdDCvf38paTRok2EJBnHHgTUqQdkGu6ricbWMlEszFWYKbVIPvQ8UX3vRb
Gha5J8YPAiQ81nHpn4wZNQO6+heWqFkINQ5hiN+oKVENS8vEjTp5+vbmtgoaEt+V
lYy+Kkfwhxu0JghbldIgzlzUcAZYGF5GEvF3hwiK+a3YhezDXr1PYpLTT0ch+fXY
rzvQObvIKdftYS1Y4d7JM7J5tV5CAs9rYsYKroHaJNzQ3n4ULXxOuRuqatFVxAUK
zkiPPKR0yX6Uophji0v1aJfaPAhrL94sLi3jBqKofSX4uMTiRYs2L25Jpvxn2JVw
cBOSUAkAt6F+V5ZaiVtQezolfPjtwDfbgKLbd9g/5S0JO0gg+ka+2IkuAZz77AS+
gWMjwVqERfhnGPmPGuLuuTjet/AHn7JYX6E51H6hlolAiU8ntZrvnjeLl6lrzyGy
JKDhab/7pzOUQ5nk8A4SydqBPlZebeWjSoLp4RRrpUDL2NPn+bfxqzglyp4mtr4z
AHSE3+IVgvyVjgNJnIYWVmgqvpmHGIBsFlAxktTpvB2YBlhxjz141YNqW7IpI9+E
SVlAMgJJzAWjL2n8/8FFbamqDrh7L7Tq7hLAJQQH+wJBTBswuDGZMXWtYF1GKCzN
y51F0JHFiCexiKR7W68IJqcmFRZshQD0p1cenJnbQtkaZwMcEfdTnEn5mgjxwqcV
5qXnWEvmi0Fs7sdcGXdVNDT3WJoS7sAwOjhsrnwVVpV6Rcr/Qn2k1RLDiPEHoZET
b9CxknMzTZDKAoFPP+XB3gJqSwAV+Kr6vLQSqoRTgumPnDS35+2N6ZcRJjNaC7D7
/HC3aK98JXt5UQEu4/RfQqOaF+Al4mWSqIhqpexyS112FLJdi4a1IZx3bNYAmkGI
lH55DpIyBfPVMiP8gqPstn/NUCTm/hJuzTW/YroY29UJJ6rXyBg322ENEDDQpZMi
1Zk895zPhzERDR6VklBF3BnyFfSfh95QWaa0JoYhidAThxFEE78NsKJwr6XL31tz
mqof4/9Tp1lggI1WlUxd7v1ybnjI1iSBcDYYLVQ8wgemH+esEVlOyCml5lScvopY
LB4KfBh2K8mXsSrEGm1/9f4Fxvlx7w5/P57HeD2Zz6CmvS6aL+lgM/FHccdBq9Xk
Gk+caXJx9mqyvCbLqBIOfjEq8Z5xhaF7+h5fsdbrR0Z40nbHEZmLw7FfhT0r+0RQ
3DdMB0Kc/vmWPB2gjt/19K45mOfreGr9WXy1xXPjFBB2a+FRZXsn+V5If8HMxVEz
/JN14TBzLf6l9ZAa88crm39kb9G1m0KIx3bUK1UVW8tOnZXZQXIFUhXAazlSw57i
uhI1VtpUB11FuHHFyGzkm65OoEOVzN3h5BJTh11nZfilJyJY5Us0nDei70zyhr3R
6UQ8qlJyv3u7Cip1KjBgtGFN69WAetfu9sPUnPvxAxPJjiS1I0cf0lTMCQb+LYwn
+zdeeSMmVd5j7eXTvfy16Xwbq0MqQ5oO6WxXgNww+8Vutv3yVzAnSzh8UTiUZuMS
WrjEXYHgtHd7xmnqhZV+dQJ+M4/H1ckpR2w2Pg30ee9jCyagcksjXCjxiqaaUWZQ
U6OWmyIW6tXo8EVNxweRaFREJbdvzIy7PtJjbxyXxATIvteuGYyOANLzvkrYYCEF
DpydEJzNQ4PYBqIuDgUyYUgrOAn9XI3cFT5D1tQwyM2zfbVhquMegihmJs6vH815
PuyKKGSdvlGapwCzIDmq3Bj9NEzW8riO4bi5bA74ktPKciD7cqbywfBxpBJW7qZy
0wUDPu8KMx4sGgBSITBcImbnJwBPD1BmcO06H9zy4yDvHlXVdiY3Wcf+3E7ZY4rx
7u3h3mKPXyj9lKmLAW+3SsViwUeQz+ZLwxvsObXw8f+sEZwpTYXUN0TIovYtM31+
qiGByOsTYmIXj760Ia7QrE8Dz94YDcmitmSbGM4LEGIHp9/ib6iX7FE9ahE5XKPR
6BpPnuNneLmYTZRVWaXfrGDkGUo2rQS7zn/TyKJHWmYD9n2RCROVSSSwzqo0h2Yy
5DEzgymt1y2azS0uBburkzE2vx/TcGMfJGnOw5Ov/T0O4W8V3AQvuU0s7mZTvCg0
9a2y37weoQpAXZjPh5NweVir4Vy43prFqaXdi+ihFMsTSXtt+Ir+4Y1GfVXyj6UF
Lr1ISa1y7byLkiwN47K9Tho2+4J+eobBY51BU7hLUiILk0I/1iKY3yp7Ra2ZDcMX
iEQSg3fvzZ7KU1WusZsEOEAs0is+a2g512rVLEvTjDAjykt2rhpp5K4HNZS+o0pV
zdF+wRL62pcXIe4qFxZeWlbniSS22JBXsJRDejcTPtebTeHkFcf8WTdT2BHD+F5x
1C52IJYUpzZII3q83axEU2JuxCrug4bYOQ24eJ3nNlcdpunEJTjHkKdpvRuCwvv5
Cyu4lXpF8lR1HRLU5bFHZ8a6KvkInDBBZSANR+NgePDsGDYL45bcxMBSCA2tgwde
TXlZtW26Fzkp1isciXxVUvyMoYfEXRHYCQyFDH8RhnsnYCL6q+kKPea33r+W/LWB
Y7zvXDU6qZntvbsk2ThLsf/Y/WngiAw6FnetUHmqGmXN1ZxmWrvf7BYMy+918Set
V69e6dHps72stsLsK/PrpTakj6z2apIZWui6k8jqqqnqzi79gPaJSRTUW9C+uIHp
mTHGfatZzNsKLzKeDJBJJb3jBmB51sgK1e96/EakOeCQl0UWrxbyt3u1QxtiUAJ8
iwYk6LT4Vt8FhzFj+P3opmdX/ceozqXI/eMvdwSZ3Mjm1yUeGbR8jMCAx9vlAkgn
DFBXGtnH6QJzwjM6O7RN61FIJhfHcSJ/QXkP7rGrcyZLMrUo7ExvLrDIdhpfO7oU
2dX4r30Aik+YraioAk/apHckBdYkLs+DbcjgrxL2hP0Z3zPY32HRhAj3F6KiCbbd
3iTAT9jO5HanrdFAowPwdD7U1lkq20hL4hS4lCNWXVKrcApEUEEZIt/4apQoDjl/
okOrOAtgGf/GfiSK6fx/R6yXGxE6ZREB7WZpVt/RuX91EQA8Zj0Ff/bZ59X+xwSj
hdsYAEmHqnNIBRhD4WqTQXxaNruBCrivWx8bTj3x4TC/2B6ARtrw8VEf+PLOVFZX
NcnTlbg3udJwVDqC1qpz7ekOxQnlIxbRbbtq21eSYllE7Gr0qAtujSQLFsew3mgS
Jl6mwncegzmNRKSQypXWdsyAvA0MmQtVwl070XUMiTCGsOpOhjP4JNhduiHlu7vi
Qao9Z6OmUlyGNISO0yRsSTVjHRK0oETXsxVDTXGmvnlWd9ZZT1/WZga+7jOvzhvm
Wvb45wbbOBOBkdWdsTe3PsxRWFOEbIzICLKGI0nqdYR/jB/l8Hev/o99+DOzF6kQ
UTF0WgZqGe3S6iWfknrizbrAqNx5hQlWPS9a2/keh4hqIAmt9IfNEZLCnI199Td2
h99iZ04lmU2do6Gn2DnKKWSoJXV4TXwlCEr6yuaI3MSqtitTNMN+whTOdWHCBiVQ
f1Z2UuEAv9WjrQpw4ESNFY0k4lNL/6N8T8yb+LACH/PL/Ly2SENJ4BbW19/3epr3
CeeTNy1DAR52Zm++tS2B2ob1EXSaK/bpnPemf2iZ7CTKoxj2Ixoyi2u4vjOl114D
7x6j16TWIS/MP+WYDlE19eUorYDhAxbh8ZTh5VvWJ8UJN5faLRPLPkwWcOmu9Rcd
lfLTUtZ+z7ocGDryLqZtOg+GSkgSq0Qq6yDZFxM2+c4kv9LLLmRtwzMsquNu0RcK
B7ltJlqju4ySZpiNm39UYGrQBogsZP5uNXIMcvlZkgx2IlL8qQh0vQxQplQ+F0wU
f4lS4lVlWTE2kZwSciotQj+Y/CmwqqjupsgJZisjM9EL3MnCT05wm8+S7akY/nMr
dtKTu29Y/pkFf4i5jO5QiG8YWAsXjoSrKWp43UkDjB8Lr2KYqJjo5MDNwT1tpzZJ
u302oWkvsH51cXjIpSCT5LspdASnT6i+NRY/Sn2hHsar3RpeteaTqusub0/Fym6A
0acKji1WoPQarWcbOo29D74ZA0rxqsuRDv9de1j3OTqKM9IyTwQ+1BUZZJROv8D/
QBJL+0fyXs3cAN5LyEAngn6n5YwejFWC+am9CkfDejx4ZMBYDoRAtQ8aC60o5VAI
pPjoSuu3sHaoEGx2y/Iso4YGSdPD76TrfOShzZQMnNziVPlvvF9NOcsWeSNK3lOw
TA8/w5xBPUnpCELnkGX6gg9FZvCTlVMgstrDmy9qC16FJNty0T9UjESoJxr8/Rkd
m3AFARltJJhwTtF7PQUqK01WsQsD48FbXA2WWcIVR7dHchW/0vytFGqShLGB/qhL
MAlVRKPr7v/Q7F+S3fJWP7VCjTTpSNGAO1qACSlVdDrlrjozsS0p0+LInYsVcZfH
cOksk3o4Q9YUmlEf+wMiG8BTMjiy8cIUb6bUNIQKuY0BmWg90O0Z/K5T5lAReTbx
ZnbJb93sYtiJg3A1WPdK/itrb3yaA1ujrZn/ca8dpPQuf/w5RxVvb1Qd/7nu5QZu
lDjBQO8BcDltwxF7QMT6ZWrJ6inHKy4XwTWZrV6hPF6Evj4Ph8Qlo2SKkRNIUk/a
X6u7jX8+SkjVkSlL2b3x02H3PaYod2a8382+3/9Po8/ULVFkgWQGHk6+v+8/3pcj
tbxo5ooG9RUIyDfZjWFwYlfMw7nX13Q1k9C7nLdAol/qy7LXJyMc8C7WJvh5uG0Z
SZQx5HggVbRs+EtuTG1RPPEp7EsPQ/0l3gKnrV6Ltlzdyqrwg1uPz8BY4D45s/XI
eiGpnmJ1Iwh+bYxvLQ4smcsvAYoiFhuxuCblTAPldT3QROPhzxf06YAV/eyT2Ewg
tcgtQRJMpIKUNsO1juX1flpE93fknGZIM450e2eQnO3z8hoPyU/lLLvjJcHnvDSl
O8lg5q9kdXYrwfUelsHj6qwwELDKGPnlsFSfGt0FNbtarmfQsC/284NBYKJzWiTX
wVna1W8EKDe8XJ0MwmWVnvGJQ3kg3BuDTUo5dAozcr9pgslv8iNlbpebaGuizw/Y
li05JcGi69GmR7VTvK6MUpha7kNLD1yQanJymy0//VVgHHrjpp9CjYpodjFeubwq
yOjmLkdacDvhlQZxdLLjokhoEqfdnL7JggjA+goA81ejaT7IYpptkkrwGzT1NEQs
g3PPCovl30ZwrKshBuyLc0kSJLtgdYanaaitktmytGLTImXEkwlp7peLsn3mFfLK
j5NZoaF3OzKEg/kzJhdfxsYzSm/Y3PIERXVVA3dQQe6f7q28V9uUzLePn/Y3uStr
8sJXRtkCMb6XMIQX2d1/1gEzV70/+ytC+iUDdWJHo7LR8u47qNifOpFBcNFaQaWx
goqOeulKpOJO+h2Y8tb9B0gmNSo3Uf8PZ4DfxBSacHVBRQXb3qC6aScW7/RbK02J
+TCroo4kSP4sox1tl4g1J/D/Bz+pVSA+6r+6nABPkqaI9ZIqz1tCxaZdf9ByQJVe
U0M8FqywZljnuw7LpqzzYNWRthiWyyjCwtbMElocLMoli0DeXIW3mHccWeU+p33f
RmFj2LP0PgNrM18//6KPbS0Xc49xNr3QYVtzBrPXauUK/ooT4KdfZ01SbTHiqPvr
C5BNsLuZuIDyyH92nChwL5CD1Fk6Wc0cS64D+0+6JxziY+CnJ4to4SVas57DSsGC
D8AjetrOv8Z8f4u378gcV+QFJTez9/VkiAnj1UCfU1T4O72O2HSU8KTFb9d3c2ve
TwAPmRRVQQkI55lLCeySgeFy9DozrllAgWDEBcHUVUT2gVDOE0tr6seCQkU0c1zU
5uVDyHE05wF6g/sP2kx1/y3sOBZdUGX2KRDZTftGxh9d6qKvEZErtGwsm2zjYBR4
yftAay1abH6rih0/JUbUM1l8SVwBoYoGnfbx/OSNwYazoiZ2uPVQhKYmg9S2oEMU
rxQ5duYBkUTwy0cNus1W5k526A6tAjN2KvHKyY2UyjJtwHKrp7uygJF1cEgVFN3K
W/EbqSHF46YP0Hoh7iW83N9tfoGXgOEmI+yWKGaMulzJflei6Wl4IFIAubl9JzrL
t+2MEXVS3a4mQjl+TYZ/szQCkjv//Pdd9jC+xQ5xECSkaywBvUy1jfEAcU77bh5h
VC1qVmzn343W0lkKRjNZ4SAXDczGwzef154J+iqNJjH58979sII7SohsbU10FTg6
R8g9S/VtomVfkQ35XpS8pEktvVv7uXAljz7p5gH8+ahTlwPyuQYLuqYBmn5DA8yY
a+8oLFQQGJCtEWFDyz2UumSJ0OdDm0daTTB8OyKlyqzDcPZneeWUdY8uKKEU0fVU
RPkAD7g3ailEHuVGgCdYamlriPWJSUJ94HFzRArapDA0Mip3bsc3xvozB+jFl0JF
7hz4nK5KPiIENh8qWffNuC1ZNNPvRAya1r9z22zDidsV2QpZ7pXb6XNvaSWTurLS
pk2aeOSYMWiyZXBiIRPh4jGxTVadL+e2dwQaLZ4lEBB2I4QXxdJVroeT0qQEvEwq
Wn+zLj1rkLWfcjuAWcivRCDCyaYidyRFuYsUqvnUjPx9GG4jqDTQSf6VsJ+aQxwd
pIftFu84QceoghSeUEoYBv85wWFq7MQzwGhz0c69QW6gsFrFjKz2kFrkLXpvllgC
+kB/ogiBSFjTw8Uiu3mtxnaXdIhlGVbFJQ4erYE63xeO9W46FEP1X4qfD9C7rIlP
ho3JH01NDVeZZLHw8YCLhK4YPmAO4UCcRVhC9YyYOud/miMMkTGljucB3d9Khs5R
IPY7df9i1oKWOa9nW2wskVXydAg9uDkhyXEuR9pRLDvklP2YUYIfsI3T46pN7C1J
+qa7s65OXi8+0V64ELB2qi8IRLXzXYAn8HfayyVH3Kvard3UMQ4IxAQ+TjsvqWaH
Bd0S2t6IyN7h0eBDHY5hJ/N2MH+3KXp5qFaE5rqGakdTUxWvtYdjGVKpeUMDRInQ
ct79jK2YVmIM2HTofLcIcxD+8D3mbKoaDZomNwF2BzK3DKLg9VVkFiNHzG6xkH6i
ZA4JFHb7fVCWBwAoWT/wQzkltVst+EFumYV/rArbEfOFz3ygqJo38a6KuY0FcnMu
+9UiTDJU210wb0lZRFB9gw6KTh3EP82NaA8yWCJkt7Lr34axHQIq3BlkwCMSmxt6
N+OrBIshiIIsAgvyPGmqpOh6eBUzoMJKNR5krOcO06/lbXboc42qlBsqivF51IVi
FJB7b/OttOoBon570+PNIXkDDIISH9BfYaAIttRYYEYZBREEH8lkxtafdVs362Ad
5jCOiqtQYSixaexPKnX+38N1xnhygk9aivqpmTwBL8dk+U8M8AQnh2zsBW5lIbhX
xz5q3yjG2oD5IvmtIjlfz6+2xC4afbKfQOElN6VLX1FbtaK++/lGwqz21mG4k3H9
qRU2aQ5wfEqnsSLashPbXK9Ma0qLkg6DtcukwijfiOMadT/yTUrtp4+SxjPNT3cd
iOiB4y5gOjgO8GwjMqANGAf2RPEwBrYaMZIYm84EJl4H8FhYYIEAvpK0UBbfqEfl
lBjsQM+Q59LYGpsv/JLBpEa4fiQoOZuKVyVbAKN8IwZAmShTsqEB51UhjYgqgH8s
y0rtxkUUK5+2nKWNnoeG9KMm5X3HbtTZ1ThXkTddSl5emHlXC2E36ypMJDQKg46B
v5OTaIS5X2joF6lESHl5PGm6iEQUlcbp8aPO4MivoGDOtzYBPL83DCCVOiP7dLTJ
0+akq82VxEBxtQQPkgcUmrSM9/cht89j6W6qJNhaNzjA7RjvsgsaauKXSWSlSh3D
6j4yZgRpEBq7xqMkrYIhNujFt+FM2MRCjKERfMaKwmox/kkYAZRHmHHlJblQe/8X
zZ2RNMA7dWMWo/HNjL7hbjb5EGuL+/eme2LzLJeFf3tSD1wUpxcSbiAce43Wlsv6
eX6422FH2TPRknN+9XRRtdCjR/lcS35bLN15MT5AzNnVmE1TOWmKYwJw++k4lUie
HtTLAiElaH4alTIGv3sNoKRIpdu2+yAqozfIWCX+/y/TYKa/S5RCIS6J2uaMUv24
wW2EfpmA891/9Rxn2lPhKDzCFJeee14rc+M3KhIKYo96Dw5XWJG9oJObJLF/DrGG
7f63ZewFzySIND4HXIsSVe+b0U+MeCsXdqMlGSwyC54p/wCwRF62ApBUePyBU90m
+S45SdVHvkXs3JArA7/QzGCInxuS66eu7Fl42TTaqXcUJ9+rKBW+foF/w3jBiO+X
ZOdb34ktbIGdycIRbuAZKIMQ1nbEHFcD3CO7ve1Cg3kpOEUWv6lpzLzSgYni66Ir
VFXQ1+ICOcw4vEvw7Q2zwCxCJo6TggSzcSfG87Porv8TBq0DV5G6SCMKn1fu2PLg
PALOOd6jvJDvQP0zVnb856t8i8mQYibs52TWoRSG+Uzx02tHtGVXcMKQ5Y50a8hr
+TmgcNMOqpTbR4nGd0bssU2ovldJKFGcJIsovviMhFRrqmSkchLHxfjsVxVtuzo5
GmdlI6G83iqX54ptTC/5tCtf19HqOOa+E5pOCEAEJKB4hKSO22rFPmmoo5JWaUPn
IDbGtGqEuDtYuY6VuHpqGjUFhfGEFE8xtiYLBt7yCaDbeO7j/iBjY2phSk9xD1UA
rp5Wu1XAbOUoCHmdgZb3ZRL4Y+XBSKDvR750xk7NPwgs+1ycScsLHVsI16svoZX+
pSlRIiEgm84HoC0Wkhn1ZStjJb25xjL6gHCgWIy9pO9fgQR5ye+Xra+QSrLHcDHa
mYE5oOvZKYvZIGa8yORACH/NRDfjduXZ6XRS5xdRVhocF/HeDCGop1JIiDiaKef5
PYYFByAkQtx8BA8OtrxYZPPw39WYS46jS79FkxeB5jeGmgC+AenfUk7958vhK4Lz
WSgY3789gXpGPr236NTFGusXoWrIc87LKIK0b4v9Hcg5giBOmtJuhRPRQLkyya4i
AxTSSBEmowaxWjFL11qrL6Yw6QwaM+GT6tjBfAEoEkCzR3b9t8WF11+2de4ZkxPd
l0rnG4LObA4PMxFM0ToaV17AidJCah9pGixFNqml8a3iZQtjPCNiPbxBrfAgxS0l
8UdACGenddJyCLDvMzpj+NWGpB88S++KmqVpwSFc+FC/6KS57D/EACE7VMvOQj9Y
VhOAWYkZIDslJHIQOrNuDDXnwu/94UbITcfIiG8DMwBMyByHmgS34U6LbCKmZEUC
dsOlz8MkzTqvIgmr6gAaIEj+aIW0Wh7GmCYknERGfChqXA2tJrdLFnX5LAYPd9yZ
fBgEdgrwvSk0Vk1zD162mis8kyzkNgxCehqDEf2aZTJKTUw0oZpsGb6/4UvyEEXy
R2SCyG8RYqN5wM0lMyJUxyB7Z7DbjwcGc7yvuUkO910Jlf1uNhaDwNuvkhse6jev
ejWkXib21K9vBH13auTtrYCYI6pe5zSBJlU0akRv/e+QAZThqxV/bqVZkUCS6207
uGcIsVbFzsNyh8+BffULHtBfPe3nl6FLo2XYbbhg2TGxKYF2pBIFy/FklveJy91Q
ROaCg49bzNXLIs4CYePnq696Nqs2NqLBz1frYxFSkyeGIhAX53OwKPL7ccnuPNdE
2vXXdooFCT24KQGTrmqjddfL9r+XrVKAbLtuCYQTY2OIQRGxEsrvdziGw6RKK+sz
NfwX9mTHqaA/SZQ4EWcp6cmdD6/U5Wa3KS5MtqEZL3yWk5PkURcETOzg1QpfrnVL
KQrlDiJBa+mxPpPsRrECM/Bmi6bPOCBIiWbEKCnICqaguVKqRtPI6z4sP/NhH0Qk
GW25iZdS5AP/F3Z5O3N1AwyB/cnF9u+HQ24xqePUylGrR1tnyf1JzHlCqN+kbI5q
5Ull8vcX2FYh4WeTvcqLD0sq+2wKeC+E0PCl4ThLHtAHfzw/exJRQQo+qf08gmFz
7H3/lWBpXc1AWnsC9VSYyePngKaCgjQiG7HiJVQXw5XAfegu2Jqe6VDjQYtOo9OW
sfZfaXMD0t11qkI4CRLlCpI15PQB03huP28868bCU5motYDUntXw2IV8T7JvYsgd
TgFTkHvyHqXB3oePMI9V8pUA+aAwjWslePAmVKDBmMtF9ZonY4SXgP0UKCHVCCOj
Xi2GC7KGhik1BZnCzdSxFeIWNdkx6Hg/i8j33EnmBUjyo5HHeKkN/mfRNhPAOcGf
b1E7MC0KreJ9EnRZnOMymSYhBA9hNu5kAPqR0Wl1/3xIiopoe5sghTj6YDBzXJmI
6Uw57OJQViyVnAoyJ2j9vwha0UAzgNbBH1JWe20hqTYf0FcQuik+oln+zSCs8EvF
il7HVXtbB7Uw43JmLg2Qi+/RVONPAq6De0VYxEqm6SvYsZU+NEQzBVAsAXE4zEsn
1jk+Ih6WoiVSq6dsYQ1pF/UAuzidWq8H7mizV5f8WhokAC39sWnoVI1jsnfbjbRt
4HD0zjG0pgu+iQ84hX736MdpwERO4N+rDteWsQu2/4evN75C+WCBJz5fkTbveea6
gSmkZxzQ/Rj+dDebTjWed8wUoLfnQ5Ljt+XboH/3Hr+VR91xyt/Hk2Srl104KrrK
zqmFetz+OaCaZaNpAE0bdVoCO0ToQ5p/Isiv4KEpCFOJi1Iwb75Jj4ZFDv7kCJv7
KG8xbR6jYxI2y7AtNFnhB0DdV0eSgasDxn5BdFCWCr5B7dHfJo/dT7qCmdLLTv9J
aMmG9cEdZwMKtFJFpzA/1VE390MENP/59Si+Y3vhWGfKYodkoyQ3NJ0lb8IZJTTC
TNH3dGUWHkxUzAB953DTK9PgLfbKC/Ar1rCGW0LdVmcyfBQz6k4RPOu0ujizH2a9
kmcUUyxgHHAfSj+i3mTCVbu0YfeSUMwX/2QLLX8U43xH7HQ+d8HQidZ+H44KApN3
iwQTdTcILCWuEiFS4aCkvZpo8J9D6rn/q8EchlVpGIVaDO+WG6C1mnPOsNPq/1VK
3lvTg9ZruieO1rU8ISS7VAZQcPUsKYhNky387EBUMycSdzTYRQGo3pK8n0/uPfGt
VzrzCAmH3zuGXoVxUohmmqyQfe6PTfoc2a7JFdpp2+17XH9tejskk7T7ALdXjMJp
MJlEoyIISva4UDdPga9m1wTHK/UAS+8C+/0c0AKh3ynYkfelnHi1DwPqBe3f/OpL
mrGWJfKsXzLTgZfLOcYc/7FZOHBnyItXh807c8Y2O0bkE+VQCxtLmRs47OrH0gsQ
T6R94Qdn/Sg6Tie6LBvfGYzvjdTnsP8SOfJ9U+/3JXihKpe5pfb5d4b12XgAwIdX
rxBTpQA7PzIIziZivfy8d81csrQwhU6E5gvcC51qkxV3JPkTnC3ajzm0GJ5leCrD
pKAbni1PKTE+B8BBuNAydj55L0EzjGj/HkgBiCKOuiC6L556DICZeoOt824N4Z74
3gRHjz111fAck1+rBCqXsEA2hX3XrSVIN4CpkUks4qgqUtc58WmyGcmoZobyDG3b
4WEjGl3nxlAft7ItZld9xLfhURRqNVVZeugj+aVI9C1QpwA9v4h6DDdE5epgvk99
Yak8cSy1NDG1bwC4qOi2gJeDqsv7HZAFA/Rc2iCbOlZFE350IqHEa2XlAiCbXT31
ANV2kTqxev/EkQgmoKM0Z3T/80zSLBCNLfxksvVZHNdtiy9kmNiWlroH3+B4QaDE
/TuXva/1CUB7RLSLc3teDHb9TIxwpiMlv2xfzksiAJ+Y1NDoudh9h5NNof7EE2Ry
vNuv/xL9FBCqilwqItcsBVRicT6aft3eW5W00TRYe10yw5TnhS3TTIsiYVvNpXYq
77ePVArJ9wsLMDDCYANByCfht9bSdo2urp8ZqDcV9vmtAux0j4D9lOZczNi+/TRI
decsFSXhWQ8JnRQMBDvs4YthpLasxpgGyDVgTRn9duiy0mUftq8xGx5rceH19A7B
i3y6natMkiJGFbgBv9CoJ568G4t5raEsR4bphlwJ6sVhoxYZwBIV/eTsnn5B7SHF
okO0SkxwdvBSI011Cm917YMIXjqOP5baI+Mh6HxJa2DGa2deQcq6X1O5nCkIVxgw
elwJ1uJ5cOJYmBxJMLZA6IMsRYv4m45YEiThhKIoJVm7IvNCAD5IbpV9W+UOBos5
MAzl56sT11D8HJ+oryTj43ygDdQumdQRiqh0VrgpoEKYUzIIXspcu1yIWMNiUEI5
WOQJj86tHpEnfL0sxeK2JInhWdo4BkQ4dwfiYWLO2TCTiGnS2qjjXQ/CW+8WNoNK
jykqeq7DQXZ5iZYpW7o5lxUPx6VCPsFteZVwAFD9p5nOlfIeRJ4LlL40gaTyJQs8
MbHNFemXq/NCgOcc62gi+KvKKiI8E/v1d5g4XZkehxTjUXNzuZbXwL8Cz2b+wW6K
iguZ6/s2k+x9SOmlEvpny48IPA6qWEQOpVJdqAGRO320oM5RNJphe3PJuu/nMOuJ
Vt3Y8/zl5fVvMoaIQnRMGm8I3XyLOvoUl+KGms31yukD9V0Ea0JzvRqF4eGAWZ3E
OwLS/tpKiqvbQpb58nB+uTUZ6TRKCf3muKn7L0+4gr5NhWrAjfz4dJXYw4HlgGA8
AsErdyKToipSpdr+nH4+Q8nb0x3blV/E9WPD9d5CnNyFUHUfD9WEkBNy23xkUy+0
ogT6mGyohcuwlEiSRexgZtb9Uwo9oLJrmnOqM6/7/djVSk9kHgwyNFW/W/w3p1hV
GSL6JKum546R/o9fsRNJxTlPcGTBugt5MOQJDR3q23d/k5R9NGhGEgTOfnVO/kKB
41+T3YeI3FymQVVSic9LUfpcqt36WunfwCsN+ZLjDFFp6jn9ciVFtAqNChGjtDbi
2PSGEQYnLFygJIzVnZXlBF4EIPWHoegdyS2ltHBPeqmagonI1IO58nmVnlpJgCZf
QRe2p2IMu9sNYsVdjEZ579Sxg0kpF8G0TkqsNE+D9Dlab/TzUomd43DvxsI9U9h1
6rFN/S4XsPQcViVmbDvUG7YxJBLqjNkWkL6HPWLXqkrvBJyrPTA6+dqQ5MCsyZO/
pVB4Y15W/AYaI0Vy0ISCKMQIa54jG0SuSnckT87EITqftcT/wUbjsJ0bE7SH2/Gc
cXFwXE9Oiyww1nuFdkjHfb6i1TNLc7+wtNnv4vuwgIDMHwQofN2hC/6eVUGUwIuu
6niX/tUYK6Q7yb9IEd2RoQOVwl2OcZhtvQV6bGx97wN0DtY0mFA5L6BB4WqszG/7
zk2nc/tBEiQjLSs0JGMUjCvUlh/XUizXpa2EAqnwugBakyZ7x8PAJeqxGPZcXzyK
3/nFyTqJC7fiPOkHdpVUpw+IoBZYZ5KcrC3ms4qTkNgMWJl/lADJWQuDKKpKyqt6
X/smQ8O5qLaq2I+d9H9owk6ZZk5aUlaoBzUOcV+ODLgjnz4rUpHhupJ7F/akoz3I
VqMEyAG61gKko69weWb2KOETJnRM8otgqHwHpda2qxjHYsinOdW102LR5RWr2r9r
DRj9X/j39kLn12mu2wl1F5OuCv8mrCHOVffTG0mkxZ1LD8qJ0pKyOKUiJMo21BaC
AhPq+d7vQziJOmj3CJY3CKO0dVLTV53rMRiuscUlJoWTdliDjFYuiSPD3G89ewhM
qP9hPkmqP/P/SUvGupWgz2zrE/d/OPmVfYgOegKtzA/uyJZafO9Th3h2e92OShQw
fO6w0njXUkqQQTwiRcn9WDT4heJNLV58/DPcW/bt9+Ig/Mcfikow2VGOmJHKIvNx
ShDZFzvrP9ET+Pn1xPsa4cumpvPMRyCB+u/ZwepiCXcWo6O1ZQWnJKbQhXDl8dtU
mqALXpVCyYPNKgBojwmOFK7boRXmJpM2/TajOxNca51UMfmRkOZ7y5FUbbuWk0hQ
rH8MN2NRc3kE/CSBqwrp07y3zLkGJSsxXTD+l1JEgoxSQzDQ4hwvYwDGzObpvzRS
NRL63+kNlm1GjKLGUXL+C3w9b+Zx3pY5RZN4hbtbh3qsoJXRgxrrunnU0X5zRTAF
Z7y5bzEOxqFESwu3uyDfTSxWJWJWOVBFkpnbmnWpldivRSgfWNRzKWl28TqlDO2U
zrR8siBu5AufH5WJ0aBSOQeYkzeD3yvlyN3HC9UfVRDkPwfc5W3gSnJP3z6bxzAz
xrR5HuVfZotNRwsAz9VQnSfN6uF2E0WAJgJnqA3SgftMIin2GCMzgHPDk9Ue3TS8
wS+dSjNtFGZywnte+Oa+IIBtFkT2sscFvTr3T7P+lK3Ro0nGpikgzmyhR5nrngJs
gvGxKARELyEYfuBd+0Xf2RZMlqrxMRltX16wY+30snZf3coyFzTPxU6avXWv0HYi
Nli05t9Ls3tKSunW26JeWQaByZkG8i8vSpml72JaiSbd1i98M5QPPTxwgo5Zr91C
Cci6EwdJSe07gcMZyg4OPg/Dy/MAjVQyfvTARx4vG+tn4XcOSYGlp+BRzsxtKqCL
1CkYQcZeLKhXLkGYfX1s8/kLMTaq2/iev8vYoyN+n5qKugnRj09ac+4Ah+L1fihT
B1cCqjVQBrdiqnqBsJ7kaV1K+/fUq2/0DV7A0G+qKSg9FpybowzGRpf1LDKEFA+P
1A/m/5kLAs3MxxvFm/eXJbyBWPl3c9ZKOhvfilbNlfQqIafG+Qw5jAM1eGJQ6RsW
wEcQ4jfKmQQRotj5Kj8eHdvObkdcAdA+FQwh4jwCbzgQ6MK83aj95bUZ1yUyJX+m
ziYVDwuxF+l8vP304UNqc4trk/EkcyAvQhX2rNT14MlAUUG65Pm5KbhjHpoPisRV
vTqlXMo5v+6f7hbqnzv6jbDgnnzxkzDUqKM3q0EJjXObQs1JOBL0whll+/nUQvTb
Azt9gfXaoDOQ5IMDlnuaXgVUY7Hluq+4tXVobhV2JWVVUsn07LqhWT4qS4OOP8o8
V1FREfRzqMyI8VnVyvrdC594prWhsp2+P2MD2zF1karkKzYs7ez9yruCmaGCLL3k
J9JgpJEuW5TuljSXZs1Sbs/3uknNyFVWBcHVBw8JEXq2YRehjtYvEw8rRyNuRE2X
i/upQblRI9v6NkK9hfkEtJPXuUnedE75+DTzwl/oye//q786/IXmi8q9zgCGtWlF
n1e/bkfiPekfWDugtbYif3UeUTyfWrq1sHued2GGaptlNpHY41MFc+jWdCrYNU/Q
4k5rSX7De8H+XYAiYvejBediSvx5uOxRBPZi3Bx1hjjyZjkMu0DFf7ZqaTgnpfoB
zgvabusKJtRzPWjU94oZHkFHRn3hO7pM6gL/C62qn56px0+kUe11zKUtcT9dHvmn
CQZxLLxBGwfyJxo89FpJXU7KpqysuaHO4xau5QuW0gFv0C3zm7s417OM+LZb1SOl
6yOEsU9QS7KGyfvABSl3uyilINKQA3N/oVe6M8LIxZ5K5G80fDOq2i1hXDl8cQWu
Qb72JfA+iqpNa3JAoHZ60ZytFS/XB/yDl4lMj2gEPFp6PBeRHu/PIDMT5Rr2vLCD
5I3nFAI2z7TlUWULPDmY3J/4cug6G66aUCwgJyfUNi0s5nglxkMhbVt2MbuxDwG5
aFF0hkm68VFmRqSvIIKno92jRG+kAZ+v9sgLebzo4fBW8r+a7V6O9c8ZNP6Ahm3R
cap+4xk8sroG8Cg4KuGqf7tTN4QKx4eFAtudlWSY5sIXFBkRbzhj/okwL4Oz5M/9
LB5rmOCA03Vj/e191hX8Fb7q4PtFDYEtuN9NKkJ2C1wPf8h+W5V/RsqsIPlj2afD
+Q4vK5qY34xNeQaKMC0kdqoZOuojCttTchd/s1TWxWsiLepmUK7fWKHwSnG/s8TX
5IfX7vTWoIoHDvZitMVIB9OhN7LQ0XpWaZsXqXZ2wQqcok6B77DpNhQGmsH0m2MO
+cMllocqthEQMVofq2W/F5tG0oIMRhsmU8arZQ5hsILBHbZNoyYSUQ0Kx3wewT2I
pqcc3p1ZvdWQpCqzjXzY1SsNOXiEnnY43RPfeU2JGdSCD9ocOWm8kCZ4qEdag32u
/8VaPpghnjRkuWT+Zsrk30crewO+LqeRlEpsjNhu5bWlFMmAY8N2vj90Ux8gAu2j
00G8CmF/gIzvOIr4sqa8uAyGoyB7yNtOe/fU/YHgDbaqLiapj8O4GugxSQOJj3ee
DVs10/mQmYFf/9gMzjpc/uiSiXvAGdjNZ6MQINxhf7IBITDjuL2OXA5i+jPMBru+
hZyjxMDeAnkvxikhd/wm9K/qbQJuja9INVvzcxfCDCu04/1SyRtLfTq2udirZ1U5
lyDNplbp6hXCLi0mO8ZPRLcmKLbn4xLDhZzSNO+s/vUDgLmUb8qon1Q2JBrbsm1Q
yqbTTwkuLI1y6ZSP01M2VbKvg14H3OiyPQm/zemr7XFBFFQCLQ8GvaCyz3qY5CbB
v+N4j69zSMXeRzdbmhBcHJztinqZqml7IK7vK2uV3JaHW5mpr0Sjkc3lrNqI1/9Y
Viw7IMEjgGM+4xA6OZ0hEoj443U/hVuONUb4dfEF6vODv7V3P8ErWnMhKAT4+aVy
7q0ZeSsKdJnkwzG3yEXo7yvOStjgWtVFuuHR6iCqHagK3WyAXv5ryna7IkDf+mpl
qQSGCIVlB0lHuummpQ1RXHnaWBZ+l5/S1j6+MIC6GNtqM+Y3bodIRENliq3/FJG3
K4XswkK1P1Frl0YmQJJrBuCLppRz0BhZ/Duj9DfnhBjiGZfB74jsVx5j5LTrTuBv
WvyODPGgMyYmBYOYomrqQvPZGtO/v5f9pZSarNmE3vXXBk7n6ZUy6XOPxcFpTSAp
NKzqeSE8dnWNh0Ikk+1KQ2TWG8D9uBV94sIo0QwKW3/XDzZOQvChs1dGJZUweh2b
zdP6tZ26wsEOI3WYrn2UmcJnkXUtEytllHOj43uf5a0VHWXkJf32sARRHSHqNRwa
tSyZmlqccXMdOnmvdt7ziv3nwMg+CoyaPs9Y/nDhmWjGg8NMjOvq/we5Osrcum+q
UkXyME2IoIwxuOaQsAfPYHGqPgfFwrBlSWgwGZEsEdsdZ4jWjS7fD0VThEip0nLF
IEnT5nsN0PMvyFei8fJEo9GRpJMP4WkezOTmw9wM7NC5Dbq8L+dXunsXDRDdzo1E
ya9JmK6KV8rfddKZKjWVYDt4WfOYx5NoilFRQLsio8egnanMMEOBQBerKA0hXqv4
EjrNzbYLbDGwtRAJBlzYLqgb6XCpBLvyThsXrb0uVD/C3Uz7JcvYI+3lWctUXVTd
o65pTyIYc76LUeFEAjn7UlT2/7yOgUP48PSwvXGpuumGHyQyS4K/drDsKPEaEb6C
jgzg9zqyvcBMf7lsVaLsy1C5wcRaCyHK7PwTz7OjjoELDyaS4RXBh8kzT123c/r2
2VGcJsh93Kcu2HfeH3ei8CHxcrW3Z9VmZKv55cjl73EQnRbryI0MPCnpm2UYRxQj
j2SOfGnZ9njhvChNENwYAW39olcJs8+SLPHZ00oJ7F27IMzSIkhvKI/b+esfkK/x
Mjjsxa89vBmyhHIKxtR8GSODibMt3gI6jw63Nn1hyDXQGrtJsmoO5KQYURQvdM19
/TyqnfCTvKwSnBxVcciENpyLBLGsJupqLCjhM140A9NjLMuer5ZGw5xV14/g90R2
4siD9QgyVqpr3jur8rIrPI9TcBaylMUaygDS7THoT0CO4F2IV7fQf5yaPdJaInvj
LiMfd6tV3NE05ricnZlMrHnNM+NYMHZrt81qvhNArNGykMVmRtKwAz4AvznDwyYV
Bwmuu2tdiC5Vdv2y0LlHsNzcb52N26mEP9631vbu8DS1y9mMxS5hUCADZPxRl+cc
1fK1vbJSJI0sw23j6IjhKXf2JyHsp1qoImiPR/Rsa0K9X4dSTkp7x6zumYZqpROT
gdT+Lgy1bqYl/Zwgu7Ec68LtgXd5XtOvDeqZTx7jqrirNWn2JZKaZEzcc7OhYHgg
oLb6ZdTBGTXJG2EnRNwQjjibF1Di3ywsJUeItpr4otgdXA8L+qM9PFd1Wa+RdUya
r3r8YHgDnBVQyWA4ZhOCHMeKhdjYL/UP+jH3lCSXHOU/Qn2xuvwo090daTApzhLO
Q4wQAeSEKLjUGXuLR4EL5xaBWFKh1eZ8t+M2lQZdK1dwlFOfl/ztOdNvjl9kwT16
xAtmKW+u5F1E37qVC9quSv6FiMNKAcRyrC0GGhI7vJS6v7HfVxhVI19v3/0YyYhk
fiOjTfBkh5pIM4WVq5QYL9258xAO+j+DTjhsZUnfQA+xUtiwox9nKF2GYZsVwaRB
7r38mq/GsZf5u4osJ4jt1XsLMZDJX+Oq935ws0pE/zI1Y8HUe/2Wd8cFfPIvuF33
wTSRWHH9ge7T6yKzJYC6/bfjJvNgUKNW56j/ao+IPXlKkMeAGHYAVUGNeuGhBh2m
eHYny7gvQvzVa+GHnkf2nN22bBNQWmxv3vJuy4BrtETZmHWgdhOJxym7BK6/LjXk
1Ag0xpGqjywSi0MZ14ua6bmeznHrjrCpnym9e5jR5m4lY1V3wpNTyFpxehIf4PWF
2R5ug1GHvLfmikPzl9cR+/OPGhrO+jH0poaNXSgc0B6RS2uOMzPEWzcPoBxuuD9G
KrA8NdRpy80sWmSgDIuTkIXphxJYDKQWd+bWVL1pSEQJQVMSYno/tH+4GoU39WNZ
WmYU5FFprwk1sp5ySqNc4fBtmiKgCL/g0B1s4qDQkAlrbh/9PtL1QWO9JSZN524+
fekmz0mr5AHP1LD8E1uRF/pHScYzfIAHLRuly7keXLjOu//aSbdor37i4OfmeyJI
KIfvaf47cRUkhxuVjtejHIjLfARbZikLreQJ8LUhiwqxhd3ivdqfuA98kP9QoN6I
sDXImMK1rNMXoJywSqOreYfIHcpAL2Wx0v184m4GDQ32S0cYV7BBXjV8BazXPQLL
jAuvj+WzdNt+iXXEoa48ihvhqCCCO2B10ESiDscIrkguszkcedmYzsOzlJdsulsX
u9DP9zV+4d1xPVVIJiySBaYG5JRoiiPXC7LZiMnNCKO3qzpKhqEnxlGuAUVkqgms
ZN52i8WEtoYz0YRd1Ri88tXCYxlj7PBpVNcu3eFgQCjRp1uIVjR9wnR7MmYuePCF
kI2sQV88G4FhBkZWALTYWZ6nLBDNRmVoCvi13G2GSCc507nLf/6HhHGQ7iKXnK7s
WF4FKGalxLyKogl20Js739mcj9cKe5ISi+twwpT/dcgSjRFvZDBzOrQ+KWPXlTmM
9jMhod33I71WpdnBnpeTHfgcA7GBY3QnjiDXZPnLR0xX7KGUSOr8VpTsqKe2YLUO
tBLjYYL6dOaO1p83gOuQOpfxwbchNyiVLty1Mm3dftF684PpRsz7i8PBUY9yCsXx
1R78Dot+TzrUSURV7LPOflhJ4BHxL4kXU0AdHOvNVydWnzAZnHo8PTB39g8pqrz8
SCNhybFxpV/Yt4wFzOd+tMYyIPsFx9BgVGxnAu7ylFqTWgaAW1hwjuFI+WS18Sd9
dtZ8jO2Ky47kDrnEQwqHYl/p2Slj9JxkHvjI/3TBk/wsw8uSADMYYgtId4N/nKxl
qK4nfB1jpmEvnoUqOoPNxY5Er6jBeSLgqGMEbX+W8NQgtTboQi43JHu8u5tv/QSi
BR0NNCgEYIjPwBbiZPnhPv11DNMy5yPfNlYi4O7oc+8EDrYkVEZWU0BzxOJrR3BR
0Q5AYe2iOMzn57e7TnP+ISUtCBCLlx2gHkkFgZx23ycXMxnV/vzphs7CUBfF40SC
4VwB0kabt3PjaFdFCeegPkOlXg9y9DusnLv1LF5jfEdc70YQwKuYONt34J7BTdbu
wvfuP9Cm85exzkRsTfJim6kMtHI+H3CWdIOwv2q5SeX+P4WroE77ga7YGB6VqGKi
EoiY0Vn+8p7xAFw8o8tOsaMa7qJo8pGmsa7zUNmU4jYZQF32/1xALh7+eWS+1CVJ
jtcoW5+JZ7ZjToA4Cqj5dbsbZbBTYkxJQjxd7zYg3zDpGqTyiktLmeWZP0F3B7Lc
EA6v5+DUlgbgCCuVKetbhSmk93dPGQVt+zZdFzJI9riOSGFHxKoojqZpkSX9+b2B
hlze+RM5jQOJe2ZYrBXrDm5jEVAzFi64iGDpwGTCmFSGsWm5+jqrrEMfbDt2aQ/u
9+C2KvvyugYHudcqzp9Tc6s72a6RIDeJZTTw92H2Q+icfB0VzG3Z1+zKB4XpPphK
cQ6/+148a8eYLSwpo3QTqzg06SpQEA0oudmtYw7+kco49J7rsPnuNnzUJkIqzLu0
QDPdrMxOpThCdK/3GfzwjnkKTXgq+ABMZRfvaohWukpkMPh2ylpGJES9gv4RuBPu
gkQGb/V4nX+PpvmlKX6TZ18cazIXM0A0WpAoNusQI9fZGS7/E8FyrbrEbDvbSENK
4RVRThW8aa3ei4uihbPRUaSvA7zpQgbHMH/6Up/817aJLlGrSMpGouggANiSMHNr
sWyyEdr2syLoOUl0Lq/M8NcYVpn428eSs6nsCDR6W+wnwEStFA5oH4X//FJ3aXzd
TKmFCFMshfYk3QmxJYXX0BJApKEtisV1qbHlsWeAoKuvIG642V/DwsruGjmhUo73
9JmSPx3pd9BSG3UhgIcMlNku0LnkqRaLh9/1pJUJnGjFkik1cLzVcqp68VsiJXy3
pFiSzEgxftGtfNFgN3/qgpJM2NJdC0QIchH6cjww83PLI+NxZyAIBVwEtdLXr7VH
HukbaLk5+Jo3YE8qRcRtkqByNzVZzrGwtZVpy1+2jDfLdgamw1t+zImNLbKT6wTD
AsS8MS3v1b1fqKBXhM2EbQef7t0ILr2DS4XkOuZzbZzq9uwkhZoRBhhsfq/HZRbd
RxY2eTdZz2uGtxQwkcC13yadYQ945X+wsUKbbq++1xBmLcwevbNQTAoYifmO0O0V
lcwIjP8GIKKRr6cIVRXrtp/SYZ4CquKYVULFK2O3mv8q0nuWRaSAGoCt7HhwhH1o
Eld7/Zv8u79kpCmASDoUOP5De1GSyWwqN2KlpMktP006bGYkXnKAB9k0WIkHsduf
Fb5CL34bzwxNquWOBVQKrKSccQGofRAzZzV00ezvIL9WT6IMejYKFAxnr4DvFLTr
xSMK2iOq4ijKHIlS4NQdh/S7GuSPa2GYsJxzWJPzGvPKttXCD0oZFXdqFo0bEor0
Zfea0Y95+ViJRFGR+84R1RarYmZ7KXPQ0uI9+5z83QQpulpX1LX2W0rL8wshCCZE
9PP0rockOw1vjia1dfkS4Prqfk6nKkptokMVIj+nXhcXbTEzh6C8KPKUz+2ABU2J
fTFY8fi039nJjI3UZudB1IiHzaGq+KTDGHAgStGiGBRhNlZ8q/YgvyIc+MRMIXFg
m38XW3QSMXctXa69KTdef1eDtsExYEzylxHrzJvDr1rRoYznqUJ34gw2Ni0W7jfP
OiT9J1GfopXgXegmxm+oIzni25xcOiBhTd7vtnorzx5E8pEVSN2sm/CImLW/s5P6
csLvGGF/LUXsy4ObKj1mTflPp9MgUX7unLRMNFQM2+f/ajtHgc7usgnYPkt26reB
t2KL0mnBtJj48USDr/82DC3qshuds/04i8YXrw9P/9oPg46GiKqmmq7NGftTg5qg
jgd8UNQjDE4EcmkO1k7rOdBDYAVzTFzpklTGIbvoQ5KlI7v3HLOq2zUvq4sqBngW
7twPXFf0WPqFOOuMkg7QiCTqedZiF+51sw2T9tVtOmxuzKgr1n4wp+2wioRx1OiD
MfvT2BMgU3xWlA3Fo/XqlDVx+FsHB7kjYX5KyRSgV3kRJFq+9qu27MkaY2iKy4Wk
YynGLR77C0HRUJEnaxnHOSRHeyEbaRlQzK9WP0GSzAtI5rrWWmar3ej+Rtiz4AFu
SXOBCodz0yNnpDfqo6bwBYMPunJ+d4FhZxfSOBOjxRNVAzyvJuEuzZ+yJHsB+g4H
duliNGoot5wITm6HPkhlSmMt5VKA3IBod0eLmc0rFXMxjB8zz58CLK8cTwpNcPA7
OYZtD+K0TJIFQ3YRcI2FAKiE4SjMPSZSeKBU3wTh7e0+4qPJk3NkydRXlfYQ3JBB
RdwJe8MVf6ZoOk9816W//uumxmpOBqB2sR4LMC6GEEHg91So8CkhtUqxtdihJCCW
6hFwuIQHw4nzBSGdvNX/Y8Bd3r6sq0Ve9hAcGY4OrSMrMbR3J2cP0Zw8MKP8VINW
SHVEfBJ+FAKII/uYixPrHksegmWJ+aNzZ5+KD+UJ48ueaTLofo9f2t4dAn+S3lVt
sbMxxDRUst70lTbDwEHi5uvZVWTbbG5j4KBD+5JU8YOv1JuzTjM+ccHiNODP6cR9
hqI+WXkmf/r8d5VvJaRLX+mDQ2FgXsE0IJ9RYfJDJUpOqok738gl68xCuqOsKtCj
bCQLGS0u3YrwvWNKAVyR74wr1ZTkDpq1kDLy5VWvctqAPxKLW5930PeSDyDluG+b
GJcT5gpV3N56tnvMChS5nHx3ER7YRUNPo4DOxtPh7XwV+MrFBQ2xrKxGG0MXASGF
4EN5UxrF3ggHKONVvE1dRPygmP6w6neBTru44Dr5yQFCacwvIyKw7T0CR4X7WLfL
CizY87X3W5iyU6VyX8YjvOLRs01MsvPDOzeOF2QSOOABqKewieVxQTgcyJ9KNtkb
4yB82fg+E5hGs2ohcNCjY9OF5sfXLdi0qHzzZIdyyXUHMK/OngTnDSRoCDr/lDRq
7LYXJ0FQ8MzDxplUQbxb2ZEkRbMlbE7OmFsxwjifPeFFhoaBjEQOvIlb8Ji+yn5s
z1vVjM/MOhlf21CBoVZ72h/s482bqOEavvBqReGv5yA/Bkp/O3rCghee5cf7zPMK
qIZ4HOOxmugyiGJDx5RHqwOBBZrRzxuhOADd47FaCoSFjkaBtoxIowMYKksIHCCL
5jBW/kEGbS1yg1Q5lYrdLTYY3UxOBxtiWVr26m0/tbfNUWAv4RBkWBzev6nMMOpm
J/4HsyMlMseXSdCKYn58eQKAHksnNi1s0+jzB9DBo34A8dQ4bHVlN5FHu15ZhLf/
HjYA57D+xntPpEX5W3hBtKu7v6iryFcYeU0T7/fawHC17tABx78/LP2h7P2YMy6+
VzJqcaK+vs8f0zrwBNYiGjrMpIop+n488UfIbKdQ4i1h9ZiU81dyO9j3JHIinnBn
uquJltFVzFcl6SWcnJMbeU2R2x3tBrsJdRWvuljF6755aw/SQZka28NYu8HkoqLp
r8oVoPI1OZR6eSUhi/uqolHYEb6VppiD265apc4dZKKMVs1pitV8X32NiBlVQ97X
CQu0Pc+dYazZWoK+G8LjSm6l3S9iVI5twQanozckQW7pqA3KNSiXFnFY6MoHNfGP
HYoqKKIbBFoBfEjuHB0zeml061EkSH1nYsv4U+cIIdMizD3ljJXBAwOQzBTCr4mn
YxeQPjq9XAonMr6wy7SwWhtdpolk7+14CcASQvsMhUR/AsD2JWeasf4oDgMZrnCB
WcC71l/i1tPVuyfPwk8dAAGDhfGZt6SX1p/Wcf8Bb3NSkxWLI+Yxhx/INn9Iy3Sg
6VYpgqGI9g8Q4wWaO3lMoOSeCb7XqMN1gw4sLIlse6w4dV8hzLQeTVy/SNcCYMyB
9HNushO7a828L8AdKxn6L5OlkzLKTygbsH/NLzb4bwmCelcrJINVI0dgHjhro7SV
GadA/z+aKe6iQxCdR7W1tX0991R25qKYZoCHSxJGUIWdbUMeo49gxpPysxBfT0Ir
WMW1NXqL0qEPEWLEkRVqZ6F9REYTKKzWsMqNLMtulpoCFLISzFWCJJ0sRc6V/5kE
pn1jJGfaYcD249OBEvbl4V3wd39Jg26y5nEFN5RkwBqBMjqC+ae24FDtpUBGyqTO
OhEretAzb5XdxuxOl7BaO9m7HXdbX8gOfifPO/00AwM9P/xnrruX5dJmj6M95xOP
/qbDlO52YYbVaNnj9rHRADcniwLrhcRlvQvwmIEr44Ov7dxfIYW3/4JRtt6kL8pc
SOavdmOVRzWEwFcsmQfoMw79TbEPUd8lSgFkLTwJyf7llrrmffSlJ65KrY7nKcx3
QH6HP1wyxdqDGkOw37r9W68yLmB9/Wuubu8z7H98UeEmrIJpz4Cg+WhqgY3GL7xm
ze0Y7aLXL1YPM6Ng0yelCgLcW8CP5hA0tmsrB2QA5uxzgNYUycwNQg2pZLnAS385
vewff7zENS+n+GHOMy59WMBDUluFclst3LOcvNqe/Uty/nf/44JtPqQaq5nQKTYw
wQz4pwgfNUB5hXvxxRMYGq0qljCsmC2r1Oue8D+C46aZgxO28g+vGs8uUrgn1T8h
E3O3ZM1MaD0rGvKXwnmwHLJKCLpylL/ZsxDZTK8wHlW9ByuBt6dPrvjYazHsBXiy
HrxRRg46fcX5I7XWZyAnuc2lfh1uS7yohrB1PxQWc0k/19fH39icU7WhwSdFDrgh
f5WuTQmU4djMjDfzuPP1ihrYz4J6WIwqr/bBZ1vhzFyXAPKIw1+XpZlo/E1EvNBZ
wyb+IQFxIL/AwPRJ0Aag013KsBI0zXSfitM1xhoa63yGbEVyinrbDYGMFq66FKAG
G5FkpQED/ehdh3tzWIPUykGKZ9MKv62ekv/KCDW1XklG4VUmmzbJELESd+arcd0B
7f8xzR2APKB/UnR3DLwrahF2mfo9CzMDYR9SR0XsmfQxMEMNxQBKTCZggqZvN7Ei
OUptuW5yD9391NHu2KJuu2QnbwDwmWP08XTPjkg7yvDF3YSaIcelgZYKaEOtbPj4
masGDRTRSbTTm5vCUN9+11/oxTpRRm+A7d8I5inyO8Zb7yljmhfI40uUcS8KWeaQ
eATunHKtsfrgSjaj3dOIftsVzbjJ8/fPbQcO2n4orpVoeL7TtFCXgY14cr9Y5Cff
jJQlTwhyod25b/mrG7nV1k3m5DY/qLMjggm9noiCkdBfmOZKzd2yIOUWeI5zLlR2
Zlp6svYK2gI88TqMDPeGwmJOraW79hEVV3FLib2L2Qyrz5VgP+Rb/66QR1VjJEYS
93roVI1vhwLm0I7ZOiL6uBKr2iMupHH/SanGglze3FFbdAevtU2DdQhKsLEaRY+t
U2arHKmfihaI22MYpKRaoX6mH+6ssDnBcrpVtOSYeHI39NKlxy1GetanZuVy0ogd
p8ou5GAqRjJUIu0WrBnvu7YsWHZaHrpDOljzlxeDN6OpFUtK267tEjRmfvZe8CU8
3If5tgQ3nJvnZhjKpH0xE+FiKQUrWYOAEO5X3zdS7oUR49mtympOa8s+fRDhsR+f
lAlQB7w7V+YvNSHZ0sAws4kVt20UsHHiozUuccu+5IkJSYm1FPS/tLyFOd4yI/s5
OvbikwQuK/FONgBNWZSjC+gsTrH/CalY3rLWFCZJS66l0L8UfStYUW0JoBS2F51l
d+XFEdLsdc30bgNZln/5hUFZYP453d3O4dv9ydCtPc6DNz1jrA8t9o8z6oxzeYVU
OFHo0IKo5l2zLQO1CjCQaJsQmaxDhN0I6MFMQ+mrvLg2Ab3EvuazIXOx0NQyO35t
DA1Cy69qC2vFTqeZTWGOGldXGQStnaUvrUtknbwNsHPCScFpkSQSFhP8VqufTin3
LCO/8VChwhdUY5wN3sZZslyRpZaOXRAUjoy+1Qm1d2tGSyleIPsRJgsd9LV8uzE8
B66c+cfaIblUoEtCAcaZrzeOArh0nWn4ZhoTOUa07kFVrE0cI7y6eYmTY1ZLGE/e
TTywUjRcKGkMDohsQqzNk2Ycjf8QVwyzuC1EWTlHuhJTTHBhznqDWw/uIZl5TkOb
hE/SfL99jeRb6WoxVBDYScdJEq9L5mkoYyfAD8N2TnvwbJWktKfyD5iWHYKc1O4+
ik/4Thns3sNYmAbnb0pDHxstGSKIhJ+dHEKQLnhMHaVIKGuyZ214I/kSsrziOVG2
3qoUU1Bv3IbMIdKrPF43Y9NPfAlWGKtX9t0vcfEyZLQxZZLA3D7lbiKV2UOjtaC4
twncSw/LV2R3fjikzr5z+B2R/S5oJDErrUaRCJvtsE1KgxrcqcwuuYr3sCWV280x
jZa5letuDIUB2TFbKru60ZVTe8pW41ymBokpUMAqSnxZ5r3EihcPqwTSOG1qYbUk
FmWkDlprRjGl0/EZhyw6YYCfd30VcgDFZaVmvFnT9+JxW0i48hVo+YYLsn7ZKJVI
BdtOi8vwOuzu8g14YFTrF1ws9iAeBiNsurIbWoeCoHQBiGTPEmAhRUGzcRqRUX0F
L/WLtT+fuj78RYDBzdwQYiWb21dR6DXratLBi+iTBilZNJlVSTYAj5pK62ZcbWkq
019cplvL0AwOOXuL8BiEiwffzylC8IQNFdEMV0mhK/YDnftIYorhBRPKhHgYqFmX
BC+OiMLw2Hrtgei9X8w7LWlPhQnQ64ZyU8BKqh5m/AnVt3//CUoah+4gTjkkdghg
rAuUAWqASobhULVyzVrd18ICGpCSwzbTz60+b/hKHxI1LGaoXsTnGIlbRA5Jd/bO
0c2quSgeXoyjprIiVc0nr/DAHwrKSNZsX9R6AGml3W73w8Jmif91VXmYu4D3Bbhi
GNbc2xLScOY+wEz/0NPd71LzqytC2UP+mESYdmYmw8UUNKWWIwX+Ep8eXL9N5Dev
K/hUi/Rrv3HHa9pGgHBWS5F6HnnVUdfrHLPGSpF09Z2N/EO2QMZcmId3xiK2rYKb
OMUE7Fofp5HU4I1AqvpJwhctXKgzg6ljcEe4ZjU3YgsWboANLTI2FfhvRNZtKG3Y
t4EB4l6UkxDii4Aod+vmTz+4dCrDljeObdHkWg1Ffn0jto/zpm9R/dICQ19IIJHO
ljr02IZOm5PdK1xT/dbur06oR7ma5M4CA81zuhAKYxF5EFz77bVj2zA9YVFgE/+z
iaCVT7wzwuG7HYkOh1ylzWEi1eqVlBZZBQ+aAY0eu2iYlgUbPVIlZz4m+iZMX10o
Ia+L/RvUMaKlhMgXa6xGLxcOYisek8D/OlDc2oe0iJrRmuAmpUHRYSqSBUD+MOSG
X6r2JMJqtR0pqt1WttmiZuBJzAo47ZM1Slgr0IdJlDFxTvmYxhGOz4YuRo6ZjP69
YWbJ5n1porqyy5pAOddCa8p1g1KJyicGa0qhtC4hJu/PWMOfH16mDRqV6hDwJvyh
zvZpX4M+G2W1MDunqESYe23ABXFJBtP18hWIVhE8jewPuDMBuJEQmwn87yNoNka/
uSIv9YFE71sMoOIsyG64f4EQYXxFfFFYy3LXjhbeHcWyEUcB4KrqqFAx1rMx+iEo
UmgQJEcDNMT/AfFVjnrZdqtipCuhKLlA/VvyzqCK8rZ5LNzbJP443fGrl/29q4Wf
2ezfH5qLVdiJTFF4jW3PY8RQpv8lHpCN2EOwjZ32kLJtXKbaOjl1YLViIJuNQBFX
uamBHI0dYgtfLaZmxvitukrRHKD00C4zIZ3IHeKwiVqFDmPWpXIrIRmHnx6t4xlh
rknn9B/7aeaVCDlRW3QZeKFbDv+GbCXvnHtvH+z/79sRdzqnGvUfl5WfazCUNlne
T3Ujd8A989mZuU4eDYhunXz8lEpAIVtgAL17BHc7Yq+mTHBjrFEzQGRiT24pOfu9
h4keMC3IpQ/MPX59PYfwoDmrNAVlKJr52sLRPshpQGUvpyD820DkWwdmIhCp5hPd
nFSUziFb2KPj+BSjs8WkjqUVTrZrq/HxnIqY+JDSO2zscdlMAcFKCjGvoFyl4w7r
sakAeed4PD0aS88HJyh8O5LU6fP4Nm2v/v5BaJideVvvy16K4Y8yc7Wt0FK4HulR
nJSWyfj4/lYr/xzsIUnYCX2Vs7Z4M2NbZHL+NX4717BKlZXSisyufx+2z/i10Dxa
CNfnANoRxlGLDANv5XKd/+Dr1qPgCC2xXldSbP9agaZ9qovA9Tpvo5y4gLrQDINV
Oa6jSYILt7pQPpktcvbwrLM9+Xzxncj62Z2ZGIdi5cC6MBPnH5oBJQADVefpqpvM
B0Mq/pT+zpKwFdzO8ytZwwilsaXDEVm7wRotKJ94zMivug0yZBRizdC+ZEPgRmHT
LZ39s5jPADXDoAq6AH/GqdWR5XYTgfuilI4rdmY/LrKcpkaYTRi5tDVj/sic25K8
9/N4jm6gwUPa81YqykAGKfUEb85abMFdBAMCwqdSxnZiejEFeBEZgCT8BnfEcFMh
cZalppRbI7i/v2iZ5hU/pMt6NR84D1Hqufb8v0D//FLnZaOIIvxla9VgZoSJ+UPb
AloOBU8aUlBTBXcEAjAUS3wCSi3lvcBOE0tzWYxrc89G1xUGFgyb2EtpsBWZmy1l
AgzIszHzVabLkpo3d4uJIbYLM0/gJJIsVads+l7aE/xJgb0vB6/hCuPobvUBf6HF
rrA2+ATZu68kwFjVsDUO4oRD/bwgtnkJPHgr0izoK3Pc4d3kiRh5CoipfJqMP5SN
hSFM2NpvloKgRvQstyC8I6TGDZb7ERLhdMLNcceOY0KvMz5G/QwzpizyGf5Ghg7U
+dV1DXmCuTE8jYAgbmENI62ZeRwjv0uywUeIOatlpyVhekJmdi6/px9oyS8FP9pH
CDkReyWrYrddcPcaoSAYVtKzUz7KXAXCiB8Ye5eFq/T7qVRzhzSJQxU9x0ukBMuI
s812w+cAFwGMK4g5pIVf2zWieWj6PcIShtdbwxL/VA3ITy31TxgWMw/XpcvOPYhG
XK3OR4dIU2QwaQdUqx7yNIMRBWzKIvS1lZofJzgCk9PIN+anu/+jdrvL8yp9cqwY
KNgb29RXUQ0ibHgp2NHU9IYiJrh4konQs+K91yn7xzYEm+MBLpYDpzFXyVQAxd7L
ux7ck0eQMraTkXeXzJ4V+axmj4vammGbzTpY/BxRe5q42oyzXGfWHBN00scw6a7K
Wp9oFgRiwHuK6z3mszagSgWo7EQl01LFteHcxKoBBjNsUt8IYZfu5FDkpLRajs9T
aaP7B9KRcp60cD4MBTqCZcDsOhLqqUF/5iFAJ/36/1YE+ub5utHZpgW6YdmqGBHn
8PAtUsQKeMCqPoYSBut9k0WS6PulZQDdL3rWz50fCgCCFV9KGwBbOgk45UCBZsDQ
wP6t2VdfNC1hC29SdBFX4/iShhGiRQ2+QZ7C1tHWEu8+ffPF8r+e9aNdB083N7qc
TtJuzvRA1ZPtmcgIjWfG4Afd33nJorKpJIPZuwUXwgIE+toLHYj5cZ58mRxGVO/2
p+NeSMqxRZXBYXqL6FuGoCIv5h26aafK0euZejZwTiyyOT7orYt+vF5ea0waHHQ3
9TTIVZJ1EqSKCe36M4+yTpLbvY4bUCZ5s8j7Vxc2f6bzqSClkME9ncSLnpKJwV8N
B2KG+lb1flXGZy4qiRqaCevaIYYmifaU8UxuvkDbbo10gAQuk1Pb5iVzVgV1EFsX
g8Ggdxt5clhecpZA2mqdhdZXe4K+Wk2tgTcIbmvB/ZO+UjxDKtULn8sPZuqfTUel
Lv2YCYXSlWpcZAVM9topD1463S95fyGiS7p149LXVcxcaF0qSQH/AJTNMWsLP3lh
GYmothUWqFye9zyyYMtIepyaA+pqWCVgBRRl7bH4aAi+B+6bTN6C33oW3P/XTnQ7
LllVuUEjLr1vaLFOFSx3elsIi8SbglnrawZKsm4sS1OgNcG2kluh4D2/ZAsJIRtM
uSTVphvjWopuxssr6eNix19BYqalMY7y2MtIA+810Oedm/0hwjjgKnJBx4vUw44M
hAyAijkOQ1CgFvlJUEmbxjyZyTwKlgrEFrI6zqB3nCUbdgQfYYcJHuqhMNGx1f5E
M6xs5jAPobNDtHZG9TfHKHnWiAZUdMs7voYuaxvLCl+DS55bCzDePYn2A0YHS31m
E23kG9y6i18ZJm0hF43Jvs+L6LMjEiThr9+IeZPCAlyevU894o400vkVfnAAY3w+
t/mjkhQ+n9YSR3cK9RB10wPwZQcczv4pQAJAgRb/xmwTK91hy38U3+aXeR8lnl76
ufWdCuZN18PxlmuZ1K7h7Mqjb9m6OerpsyokxMawoLp1envj7ouNkBH89BpVJiBB
6/HsJGIwZc9VzaiIQ7eDZU7qO2fxQ2aOg8yielt1QOwpJqE1/29k5jpMsHpplIZ9
OWLXGOo6OM0L0uRQCqhBOBfNPvT0/sSa0KorkFXwlvIL9x8hvXMnIZcAS1D9Cs0R
2MhBY8F/Lj80Td8RMt+KO+SDUY9I7adwQhT6o/mvlS3H4+HeZhDqib5y6+iXr7X8
vd5UPBjjxl0Q4IcqIx5IchF2UjHc41Qonxn2rU2I7Tg/JKVmgbndyCHarllWrN70
ckdtnnflaGBL9I6thB32v8+Mr+uZdPsu+kyRaRCAK3n22Cj1QaVIZiyd6YVniBOH
sN5VtQCFrgRxD1kl7lr8JmJwROUk9xjOqcq+E41bWNjMXViHPxNrxt5IH94ERFO6
WrMqPWxOEztOLEjYTW2LoBQDspItQ8dC9dFMqr8SVIHNKYx7v28SBaU7lYQC5QSC
u0Px4V9uzWxUBj0ePaNuKuqLc8KmJ2PvNAHyRVFTqw1Gz7zZ4iqvuF2Q368oxbR/
OKCFe9/wqpSedBmFdVp1VDz1i21H6wyk2rv25/aSF+91owb+Ka6IMv35+yqL5vhK
5G/i5MWV7qU/et/p2tl+FBUmk3MUnc9+fueYXu6eP5zEFbAb+I0vbgpPU+PhqnxH
vJwj6hC860oQNNdP30l9O4w3AdoQPezwjSD/bap0D7UeCePf8nLJUqZ/Vzb66F3D
j+23gczLv4yIcaT8RZDdFiuEMFhufxRuZNksMGtcVYXJR0Fv9lAfxG1IfPCwdo41
ggheW0KXwas5TZYrJnj8HUHe34hFJLm15XOTMy9XGCY5DxhXtTIxNPMOs5E/pvXt
WHrOVIvvBhaRUU6LG5DTNBIt8ocmGc0MAxfFmsAwVSIwbsrNQXjk1ec1DHt1kcJJ
J+qKUtZZE6LKbS87UiDd8MGX0LbPZTSKX/FKbMTFUMCPxUqDEjVG2vrQEkbaGisf
068QMmYrrK5fBgAGs6RYMD0B7DTCQQxUo3yKKws/zuMwwS9IuVJL/vBfbkh23Djz
i6O9BYrRTOmVT+6nS7CvV5NdzXb2aOXbt68sBN4DtsHxkEOlU7RqOPkjihXCo8rG
LJjJK9BEIj0UqawTQZykmUBRgwEuIsqZZ++Eyj+sM+s+79tNT84il45qevtwERIv
2kMC2C+926oZMfgiXLSCUnbF4GF3plP8ZG1V/hu1VhBydNQmtLeoteqi4FNBdu6/
CRNveXaUMMH+PxCNv4a33D66hJh/yTdBkEilpgtrltxtDziReivykyrcSYJlgf9j
ehDBx/e88D6Bnk/W+Wbgay0ccI4XMvr+0SVg4a80Ol3uFIP5mmNDiK69wTucdhcC
j/HZ/zsJeMDo3L8DtHF46P0WevH73XkaEZGSTtONlp4mm6rsCTlzR3/fF8uuEd2U
qyZz9xhuR2dYpbS9E3PdKHzwaiGFzqaoGd5RiF/OcvCgQG3BGoUdFr1UoRe5Ko3K
rUm7XZ7v+OFzCSfinPKiVT48VjWqXxTD+h/v7X+CL1I+0iopalKggjmBHQ78IUaG
8r7hYV7CmoYmGF70H0INzPO+pt+oDVgcMGKffHN8fBxewBsfB4oFIarMFAS/RChS
/24EgTjKaFEjbVFtj4etIHXxC0rzTNAB14U37gcOXr4dk/oHTLWyPikYZRQREUOK
vIkcXAaInSsazdodCaEU6aYT1rVSCQE4cie/GPxmmInz5i2dF5Q/sKrYBKznFUL5
s8hM8swAaGjyBALI+QfOua1DJ+3V6++++ntZGbkXxuEy4Au0XmYLdsY6SNJMCjwS
1WuHlUOcHJvEtlPunjP9TeRBh4VygYZnIjmqz+oK8y8CGtMmOEcW0LyzyG4mq3dP
xnxZeZ4QntDos5b4bbHMAQOUVZPUbcteBEt05w8EarVM31xuVv+RnC20QzNFY1Zg
gzwKJOPsDzFb5o/+eYIFM/FyGkCmCVQGf6rw/6FvKfE9Emi1DdwjAFHrgGxaI/zD
T1NOmCrJwG/C+FpQMcB3veyVqV5cLmgUJ7HL9LPr58+x2PX/nVFf219d/EJi6vYF
DIlmejnry3wtLqmBEBfyo5Nv6ZEn/d73IEWuUMnajwKP7H8l0edSADTqKSXLox6O
8cYt3SNJWN3Yv+zSope5cY4D5dlbgeuXUDqXyX7nR+dyGvKNZi3Qe/2/HY0LXjig
HbLN8wB2MX+p8qIu7RwCjI/x93ucy5XPyaAxXxZSdWWp702rbruO7uJPz6eSOMWq
XAkDDSJXnaI6fqR9orb6WACLkVco4KsiaZYKBMIkT/mTBSWo4jBZ2Jg6TjB5hDj7
Xy9Z3EwmiMJIRV8+8mSDizqnjbkJ4cZuVUbC9HdKNr76b3CsR76sWAKB7NhBkcf6
qK00q18c2eSuo01E3+L0FzIz00fJLWf1l9uibzFGRKUmDe23BHVyaRMkzhsD3kuc
oHuTAYNUY7NvfAMs5kAHIgyktuf5hKgstTHesAmqDv+5SqW9RdoFHEskWYg0ipuW
s5qH0FqGU7neih7tyaug2bF1WXYuj6O9EzXEz+1++bcEk01BqW1ExwdXZ/ZAEmRJ
s3xMOfo23xwES3qvvHiTQImqmoFaZQvXRDSeT2enY2zjblCyi1d9oczMf9PqiSGl
xNrwfwWamRwvKlBZI3qxjAmnShdC/MxiDtMqXHvSH2Q1QR0oZ8ny7Lsj8aXs1mMM
7jkqFcXdJQ/wfqRE2eQc4m0Jo3JMyuLZ8jl9/lO1wat1wXb8oT3EffVPGPvxVmKN
hsy9o/YLS2ptwn4XkJ3io0/p7nd9yf+E3hLekY+qYliRyZELt2ag/ANwNhFesHNc
tHTOPdI8U9ht3w9VS2WQPTWgeK1/lM8bST5WaX8WuBnZnG8Twk3mvi9aLmMMdgli
4LIwwyYGQh28fJr4wWuc71NOhh69wltloPLDPjk5fB04w8CA8JDF3YGsEVFS9l/y
9HRakCEQi+Az3upNyp0/K7KXhm4LSYyKc0sZD+xYwMQGfZuTIaDNtMKtKsWXrzIN
NVjgBMdxBSD77Tf2BOFQwge29Z4Erj0DQr5TKLmjOrP0bFML+x0w74GcTn/agID/
y9/wyd6yr963OM8CaU3zmXMgAKPJCrK+C38qRX1sCp4pICvUnhwXkiYWFv8EnwqZ
jHIBwBcRIP+vI5XWyD65SktbNLRYu1PbDpWE89T21VXKILWYsJPnFc9WMwG1W75q
zgIb2E0epzNLYvgLlJMn44Pl3b/FjUmp9oJ9yC4t1YiC8MzTu2WKz4NKTXp9BTxl
Tw/YFq51aB6dYjhC2wkFZ1skCRKpvMQesIfl0mQD1jMv2H0M5FSysJOJmA9P1idp
fu2Jmfa7EiVat41XCTESg5LKCLRcjThZuKtKA8dufMmZyEXZGj7echvhbY9tG1U2
+2V4L5qV6WDSz8R7QfLUeK8OsrwLNUuLflvJjxp351vuy9ClBd8ZkkuDZdjEClE1
AySrCVLCm+ziSlhiWc1FL6QjGJ1S6ZpsjJh02ii/6defOEFVNN3nblfKD3S1phRV
c07TVtU6EXZmY5XEMCHdoMpn/vFqruSLFGdimXeZSo/VxHqi8eaf279cjyfVpwn4
a+pfovU+WGCzfGWDY4FNmj7ybehNGG1sgfveNN0lQhaZMjOAs8kZC0EFbIeN9bYk
l3jhAQZlWK5bSz37FIZUijlCeNNF595x09OK4IPdXENyYBjT0rYnBhhLhbfD8N2D
NbdWK8uOk7e9X970m6vO9Way7jfcw/9JJXc9JzkSm3ECgCZzLmecUehrkdbFpU6R
TdjQFCcyL0nQawgwh0VTWtlBdczsD2J64TQ+aAYQlbU72VOlwCjJZzJsCULeI+0y
Uq3V3Du+5nJlJVU25H6Cn0knYu4ODsSmseZZZPy4iJzdZbd/F6hVdw+pOsM8z2rG
70HHVfJ0/qf+S35cdfBmDnkFiv/QodJTcY6WholEIAQvbJZms2GQvHB4VjCq93dj
JrVYRqTclq6zKg+v9NJo0aiPeqJtiZvt9U4lF3aKaYOokfaXuZNzt/JnCxdP4gvS
8eRmuqm8XjfS4jCvBrIYqE3jGB/kQ+Yim6+r4OkzkpLlQDkPqrgoseE9MLD5mdLU
nc+TNm94LkMUuAOwuChiRglAhgsybmN/f6RTXrYwYf9E+gzUKt2TiLPwUt8e836Q
zpx0/i2tUKFr/9vFnvlcII8Eh2QPOMgnu9LA+0XfZ2zaV0Df9/qEHENGdsPiNoWB
MoLzqboXRKhjoWQwSxtTUFbkTDWZZ5dLoyC6ZJUFuPoOJgRqNheIofD/GFzdwsTR
jxjhr3+apgGNQd3PRiWaJqlvC9n67paXvNKPjhZoc/V0yB0pHKW6w4QI6bwCbuWL
lqtFk/N3cQCBgCwCfDJClGPo9C62nKbJIhccrzXfEETynviOHJMpRsrbFEKVViSM
56LqDAm428dQI4Kh9cZwcdUQuq8Tn0hena9XiBsS/XcEy5lIu+R4oZuk1w0C0MZb
fV72BUhkHeSK3aQJ6WksJlSrX3ohSkweyI8vXHelSlQRzWm/ul56BAux1aiSuArm
sG2f9lsw69NdUivd+UaIDQFvnW1gGU4NNSuNm8tD5/1+Lp5VwtFItjHycYwOhKN3
L0Nq4h+AyYt8nn5Xdo9Kw1n2dXop0EP8VQyLECzDS0JR8NNwGKtujVW4+uNEzSxU
QnAwzUp7xeYTZCzzg0HnKiR/jZoa5BuWOJQODR/WBSBHOKuNZhyC66nTeUljLTJr
qxpFTTeSwdcLJbfCJQPjTsyFf3CE/Yj7vW3H1amv70hpTy/kK4+ZY8j8qmGhZON7
q3Xg+t0HwBsT4kDGO6qMnKqrqwFbD9zD3FVGPZEp+0GDtD0nry9fT4rgJiwWBK20
IYU2GpQcfclIYqAmO/kyHh2Fi+IrqEj5o20d/FC+r6NSH899UQ/bT3XnT9SVIIyn
9y2DkKZ9YYWyZCkOL6vE2Khx2+jg8g7Z8V9KG3hddZzked3in4teZfEw3sUb6ryE
7WHgrXZr5zXgVQXh+XG3t99/iEPMtXt5xMBzTFQLxFd/63QMwKrArEFVaqnA8rUn
IRVXLuIA8PLVdKoTQcqR2HxolnQR9l2vSQOvt/+IBddp6kQ4GF8p3tysArwBMkzo
c8cx8Zzxg4fq+J6/ifxHv9e09Ki7vHxHKdAlgKY4auI=
`protect END_PROTECTED
