`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nz0LjSq4EdrT5ADQyIu2vsM1IEiKTcfDT7NkoTvgSCIC5hPmMm7tMywEdykKsMen
1aJTkL8BpPvya35d2+16VvjSg8RWH1xJ6FtJ+hIIR5KmypzQHUK4/K2VZvLBJKDm
7wVBUw/i+36KnXcDwdDR79GeIbC5LrFIMeCP5RU1QHe0zR7BEay+SRqxUtQl2s4K
xjoLkv6FE5oVUsBcxIqwvTi0AwggSgKSKSxem24iqVkyphDlqsfSWb+IHxvPU/ne
P7t5UnNPkKRO3DSeA0AE6PKJ9rEbcJd9bAgT2hgpWYM=
`protect END_PROTECTED
