`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x/xzE3tuSrlpgz0rbGcD4VG85qWGmadi3mhFYuf/dh9P7a6kWdGJeGibPxl9bGZy
R1HUkcw3ArpdfodqiTTb4Exu8LXdnMbxuEUkQgc859W3YpFtlHb0U917aV2jV6xW
rjk//DREoP++x9s/zKgsT+AWCccw9xHPcroAoJkhfp0UIIBJM/6fjTGGU7hhZCjW
sxQlqkGdr41dOfpPd9xYl9mJ0APWzg6u2UBK3lnnjw9uUHQbBqfoGnn1Qxd6U9Dt
jLM8FhsjjP0RD20mATAFygqu8thLHljOfuKbX4AqwpBZKmtOS2q96UNrxeEpSNEC
Ec90F0uHH6EiBG3sW5BZm5eMOVGYRa9V/uU4QgUzUnYfpPzO2FFu//nv1nWruWqW
Aq2tYtbkKAkuUHiuwnwCP61Dyxeo5oRqGNWyRdCJO8n+51HsYbkh2K+ZLKmmAaIS
6J/7ttgOIPmxOW6WHGVO9MjmWOhAo3Uq9vFBwOHGDbjjH8Jqlc1+o7OV5HrEGA23
yfVe0ag9B2/Odr+9oNMoyGPBzUuJLbP48YsjIczPLt7/7ijeEcAMZOVQUDhDAUpz
m56053DE4Jh99vdNjU7pTVgM8Y73nzFcY5xfZm5yzfDSgdvBYFeB84ikv4FT4W+z
VMyLgY7FKTKSzjJYfWtENbicFp9xieHdLedGpTE5mb08UhcwlW618sg5ediCvTFQ
GIx510T7dHQiwub0Xe/EyG7odd4qc1EGYCJAhLqgWS5d3pl6mvc01xg8dPhaqog6
KUbyxE5ND1VpqfmUnREem2fL0iAb93MaZuv4LFPZSd4nPVKtl6XFRqLq7ocxWFyP
b8ScCJxGZAMRQ0vHX3ZXO9e6+w7+iYViAIqAY4dRImMldwVa1SMh7qsWK8vDJrxj
txW8GW862dsLIJzJ2UADcjBt3NTvePkokWPY36E8yBqvR0HmC8W2OLAqvJ6n1GgT
Jkr3IyQFtJHHDAuD89IfngdUlHHg84KMr+K2FX+iKIT5AJUK+sSBFJUlM2yTjZbl
1pvcwR42UA1EJmeWodVWO3ZpZajT9I1pg2cnPOydxLVmBeWPA3SVjDbcCCrVYm/Q
0Fi6IHZ1HoR4ikG//NoI/Heb7vP0nErF9hWRnv4rJoF3d+Mxg4odY3hNoQ6GqiQm
/df0qKU0Q7zQ+ioyDY9IKS01H9k60iCZUmRb5c8lP4PqiTqxoohp4O5OHTSR6XcU
KN1uzPfRA56DxoPhxyF4BR0hvNA+Jd+CiFj4plxsJBqHMYCX/iYVeRJ4NTGqwynq
rUcw1vlqQiWIrM79WFFU1mhTEPlx9lY0v+q8QCm84Xg9ziRCLYm1SlvMNdkDL2yL
ZudWcCm64e/gujmXKKg9zG5S1boZBJL+vr+dt8PpbpcG8Aw6uZvCeSaVkwQd1aVV
OkyjpYlOJ8NCP58ht4BKd96Bx6+XE4sZGRuAULbH0M/i3jMLGTl8BT7jMV6V8fB7
oS4NBQRd3yhRedjfH9MmmjU285C11asKMvVXB3EgReOkQ+GWLqP0ED/U1CYxW403
3TJ06H7Pe+sP2kexeNlPMgTaYcBUdwk/b8rQH/dyrrWWj90kZc9FRUvAIXfA/7HK
yfI/zt8r0N5Xl8sfWzcfPgrPTA11OoSURpZdLnQScMUK5pktPw1xg8i199Yw40qo
dVKtUcNsV8GrjNHINET8Br8BgDcHnl9w2SYQaiV8FIM/w7PaV7iB0/wTHLQfcMe3
gYuudyZSQOGSprPVhNb+Ypr8o6MtheE5/2Rz38eS4x8KUrRQmXKfJ5el0ymn+SUQ
TG+T5UodiLK+PlztoZdLE8SfpoLKIIjYifbs7xU5Rv9klvLpiGpO06SY241KC02G
KQ5OXtgGEALamOzunfRjgtCoitUdk6kAHYFv7ZOJivdj1o8sC76AjPYpzSQ3aMAr
AHhsXT6cwg4+5JTTliCaGl7MSJsO8D7nGm20KbvFGvNFC0iL10ohcWl75nedvFjz
9XdKGyGxUI1OmzLC5Dty3zYvf1csCuFdWLnjxBBpqh6fcsIrwhIvtxnoxTcQxMxN
aDcUeV25H/Qa6hyZnpxRZp18pXML4if0XNos3de9fYujUsTS5gby/Yqe0KnTkJKN
pcPIAbGqZD8DcTR8jMk8lK79/y26X2OVs2vq+aQhQSgRzI/7H7/fNcqRnGEO3Dy/
dTktkFP0QOloJ4cFyUn9/jiSOVa0cIHqDfZ6UhNCUwcUSeJkPuCkBiMqEgqhK4nU
nwNcckDYcs3IueP1NzZ5RK9FBMLrdpp9569Io5xCv5fG/8XEOgtpatIyugfFmQ/+
pag/uhSGmosURht2wLciW2clGvgW4bRg0LobpBXxY57ujeoM+yEjYIOua0QgmSD+
4t/7Y4z3GQYGYZ/d1vrRoIQR/EoudDqC6QLGngGbSSf0yaFK4F0MXCCJwLEJEF9y
QxShHKJWa6KgriEGS6P6sdu84FMkYAbUNIf1PGx6PJVKo8MsiLCfJppQEKcpoyOx
JfTxXgB9yhFVn5LPGLxqhvEBG9xJHo0zeqt0wXdHrNq0iWdEk8RQcztiqdUyYmMC
apmUvmq2Tp2oiyrg6AaMIfwmsov0+t5ypI6llCU2ijL9DeU2eta/mFCyzBphToVq
lPeDLkdyVTIUDllNGzjAG3tngqZEsmzxVIoa9YmkQssCdQs/5fsZN560/Iy1eew5
yY26qa1pH2uBsdR9P7kLyNjuN32myo0UW4DAysCNkbvMeETefjjOEkKosRoQFddI
vmsjuYeFtnoGiaN9iur/ZH5hGx4ALi5JA1eQH38AxlCxuo/kCYhWjJJR8LOvwmNE
SIrAqXFTLOBTJeSncDGDRr9BqtLl/BD8qNm1DquLTAN/PUBG3AbgDuBNs+QN59LF
dkMYd/PDqgVZQavCRfQJhuXwwu33bxwOADNjmBwYPDl+UQR/EZuYHDk3L8PyfgBK
GdJyODqopACGqnxTZh5i/ft632XtBk66mOIzNbXOLQBfd5j7tyEvu3WmwZ4oESVd
EZ3Usk1K9EJRaDfJ4kwgZUA8xGISglOw84sO3lTSsNGrqX/i88WeU4h1+OVlYZiE
vCinycoAPngMYKVsiV8DiXaR6yaFaNLQdmZLpv/WKkxJpg/ekUQa8hju4R3CoGPN
frN/oIhR6MW9f1SFhAKY4gVeeli/8HtmCIk9VcMmW4xsrBpSSur8ssbNY87iMoqq
nptffKBUTuFKpWpdiLubf8ALFByXhvizWA34HHMFNz/GV0bCJChyHjojbNlk9zcu
cXuhA72sPK0C3Yt+GRxGhQRQvybQtpb2LfygX9QJjEZielAuv3n7n+bxZzKNgmLv
DTA7lGzuHJF55qeUC5j0FXzfdPwT5laFrDHD8IAHRKkgnX1l/jDbQ6XUbiDoXgpt
e0u5stbcpFsxzZ0swC37DK7HNpfpcZoIGnE7ssOoaIE2Ks2f0Db4xd+9kd1DCa2y
KgRM+p+H4L8Umi73DSrIEUAUeJcO0IM4CegMzIUeDMPWmloTI8UEXRqWHQkzq1yR
qqqWEkl6ShjNw1jh3lTCT5mm3D9X1lgG9Im3wvm0OD/KCtk+djhrvRvVlSi6VF9Q
p75PfE/uPfMWd6s3L85mBTyKaTbSZQut7KP4hJiMYwK7Jfznkjn7xw9+tGInuJDX
9jRPthOJPiBvAkdoxCYUiTR222ehDP7st6ZzarCYCUyH41FGZdR0yUJCt8y/vwWO
K/QXOqgiG+AKhIgEGVfTeaLP6acYVq9QEK/CJ4Xj6R/kzbfTH1Hcn7WwAAadRGBg
mEANgBDayeMz+BUhWS6PPLRlfm477XL1qGX1XvX0keliYN+gyaNYX2z2yhnEEZc+
M16XMi9Fxx6PalFO1kxUtH7ssJC3jxARg4g3QSfJfzvnBeWqt588B+hL3F1KpV9j
J5CY+9q01051KBpPEMVOHh29ry/NKFxd/tUpygJEy+PlSFmf/CCdzuolp7ittLuT
8N83KgSL9fcRT+VVTPaaXkrA6El1CBP4AMfTmECDTxZtGe+ILP7H60sm3iLsIRmW
OrduoGHdTn863GHPkHy2MKyBgyYfsFxIVu7tEQsRsBJ6pfOJQS7kChFNlnN+XfYt
twLaFICy4C38z6tqJmrn3KdSiFyJwRi4HItip2L5I7vXgRd7jw5nm1wBM9yGIqRK
5BHufjSoPaWupVZNyZEFhzGCSvfPyNvUqSI2zISomwoa3mNc4x+FqSRv5ydUfZAT
7IOC5FQz7A6BX2HBTM50wRyW7hbP9mJG85lWcX5O6SwY/xoW9EZjHZ8cRp77snlJ
zb8BfblcYBXlOjpj43ExYEzjl+pYJWoYWnuHJfetbKkZ6z5a2GKNNMFPCUdOG69X
0fvYmHuDzypMNUWX6LrPiYwxOl5AtF9KZqn9lhkyexw4IA/ENjUOx04gFlY2BICZ
HqYUmNAq8LYGhgVP1z4SZeSCDB2NpqVvhA3RZ+aLXfJQ0Ur8lhwop5EmgAWgoFhL
Vs5VEmj+7o7O8QuyGwBm/UAVFqQNqYA65gYnn3XbqMvGnjSAK3ACWaoLm7NaSn/P
ssIbRznc1luh3xV0YNFjANhS1HWeSNm1YPqoH0+bEi8HT8WmhEkVFItlVMHNBKAs
J+GE07Y1+EyOQAcrfnCIkbKGndZujuEjOfVgAV9cVwJQSqj9nbb+nuyvYjlNPNYJ
wkaX64cwlnKS0+fTZl64VCzM2ZHlqatOjEDlgS5uzaL/7Vhc3D2mfH261AEdfxLk
/8hD6kmJAhBecpuZy6atRNwZkyFj+VlH9wIkdYmyDZdbAbuNouTn+/sr+pwGURoD
K+BV6FpNcbJTfKDYDmyrFrhON5wnB/SEKV2g7VF/leRO2jFgm4MSGye+iKKwnwiw
/VTSfRcLJITUSJOOO9H9H8xwsDirwyNahOjFud8bMIKCjtRYZIB4LkHvBzgT/IGj
wpoiHTv+aoFzxlae6BvHB+uQoCicaBAbyYs3oknPq/E/H0vGRTOnkhZuj0x2CQYZ
qzRVgYXhY95nuPkz/Vrb1Avbst+dvGkOZMB5/mejZPFxZKkBslO+y6fTJsefj35m
DONqiBY9PWSw3w1wWwK8oSiHmsmswam6hmlCE8lv1kKCTXIaxhmmdNYp4XFp1m46
xkSw4cQpH8WyUwnDdqnN1ZaQZXOK02ye95nSXZsuU1Sfpd/ZjQMilmo+BENZu7pH
vx6T39wi03h7jkaixZJ6k1G/CjWAs0e7N/BC5lh1Xv0YyFDK+btTiXqAXhCxaAbm
SbwM0Esuo9SVh6GkKv3fEw3JJouqJq6jufTqjeL+ES3wEksWfgUfF+Q1KPGMu0Dn
bPdBPYovnUxlhlXg5EWcdumAdp4TN6X15dFkBFs6TDJmydv+uxcAoZoRPouZqE62
fKPDrU7fbZLztezzyrXQV2dCjTABf78WfhV1YQqZjdk2esXMBdvADtp9aBDofEki
ofX4FMSSh96IAk/j2KJPRh9sDXsBBo8XEpQInNi3zNibXYstlq1KqoAK5izTpnkR
d7wsEyq9UN2WIFw99qv/FW4QbBHHSCgSM5gLvg4ADc5V22C5VlF6NrVaVrc83lpf
5NEzEVkUDOL6e9gOa8kT7Tn9MqKQsY9X0+CcRxp4EbzBxij56oyZ611RYlFyA6eR
Dn9kFbAzsoyWh0I98vCdv1r4Fp1TMIWgMuRpo4zfRI7zjB9gr6yJ3epitf/ZxHfk
d1ioLE9tHEynkifkycvxVw/rZ1ovJ3VkWF/rKVx6RKfaa32CXGuZH/6ESZYpWrG9
98Ub+I4StGDh0kwIjo693svJWyiZ3s31UgAOYmgI6Qf1RPH/a9XeBPNZ1QCTYoWX
uof+CvnOtslA28veIAUb5yCcgxqUuCmInljTcqjgpDAta6fSL2V3id6CHMPkE0Vb
EITpvqS+/zKERZQdqj/JsZf55USxfDW+HZsbVZK6p3g7k9o9cmuOjdvsq4yqmQnI
B/X9ISTpfTncMYxUJZJUrl8oklPBKpte+dxyZ9fhUEf86YOalyygpC9g3NLxnNFo
mMScp5bJMiK9XYyHmu8QYBIp6nSewQaTLvfH6gyu7X49K2QK/3FDHD99tTfNjkT7
s8RdauT+ialf+jaeQtQkSakyF8BZpxkYN3GuDMGgOn4kTSiqPJdzRskMyfcb4bI2
i2WTZFrdtMPqdqv21a3zV68VT+/UBvklBx8105Ti4/yOkSYrdOl0KoK9CvXx/Cim
BxaowIoV77XBs1R9W9CBJKZomaalQhDBHZW2/8t21uu/eId9+zyQpMEe8xv4NwMk
W7kawKqVq+gOQfKpMxuXYTcUp0KJZ8/xuznV4wCWLoYTldQ9sV+nYhD9hB99OR/B
YsBqskWxl10mHaw/MCT9TBv0GFNzUR0SFmDmhtaY0fWPWZi4aACS0RqkAzsBnb77
NTsfvizqg1YkQZnuhSQA9WgsR+JZ7CebGDMupqCPhs4meF53dY+ejwSDvDhpWFxN
c0KJV4IcUlR3P+DWFE1NcqBRHc7Qr0NenbbTK8wOgPgHcK13j4asSHm3BSEzOL+H
gUaeoYnnYjxeuKJgoQpa4aVllIOjdFr57bpRXowzlgR3CEY3P+jhA30WogXjdYll
dSh4ma/JuOgkobJLA3yaP0WIGzYgCMSAS5GE80ctiU3kHY2M2qIcqzpG0KYRStAG
PePBSsZqpXHCGrxaRIjhsHitKxCdxMNHUXv0NEHCaLLcb+EhRwmkTPhZEQGOfITq
q8yfn0kxmAzLetzwRBvi/C66pQz2jEikMbo+9YvOUz89Xk7IYP/yKiZVbFI0llqq
W1TEAUfLEgD3ex/SSC8fm8tcslNDGI1HA9CAX4VxXv7/0ckVIpREBnhQExdBER/W
gJZZNUInVRxoLBR5GHTQaQWmrwL+KIr/4gqvzacG0Wm2p3IhmsDsR6JAXWTSexkx
xjkdugalrGez1d2GSH551kwc4gPbQ8H1RyIqWbX/eiZtSIeeY0SCZTCVEzw6ND5+
QEjvxiz9JFOfRr6goV2FNBOuhPb40Yx9cklkytJTlZ+ffYJZvW+0OZmTbc7XZ2uW
zqjAXBxPdL2e033+CkStIs+NCIHdt1oF/JD2fo+IVGkyBBlXLegRZnDpdoG2RWxR
mOp2lp1Kabaz9hqroIdm13TwufikeKypj8F37HDf8MNmf/7PXBGcXdfTfSTC0oUb
CPmHKK2Wnz43578pLV8lAq66BjPjFDQ6Do/s2tQN0rXe02igXaFh+zeBVqRPAivS
3HPfx+sJ+xD0W5gptWpB74RQvhmZdp8BADozxL6psZ9QVt8gSclrPB8ETGTQp/Ih
UkBfIBW+dTslY3ixDlxdT4iO9oaameO6vQxTSXBSGO0eZ9EJhgVlIwTr3dxGU80W
llLrSEUXAxfj1hJbQFOCBhJDHod4PzZEEsbYMzM83FwNCsOVcD0f0KhF3cMF3W2F
u93+WJjXnONhJywwDsMG9WEIdeVI9uQqsjYPeya4MqYLloOcacTD1MVGirOpPWVg
EAsbzfDaXtpb+q/RcvVBPPxXN6Iz7hWylPFWolAEFhPLfpHF8aiDkcwoCG+7lrVQ
0+ke25t2VAsyPQ15MCcrOgqvLNXzOxX8l4VCKLDTpdBiZXgJgcy47Ey6c2lY31ze
C5lPksfJ8woCP46KPRuQUQ0/IgxbNXIsjpvwyiWJRbogSMCeRxYlRKn589MPgykd
3JxRPFag3VOy4q6OFDdyA8WwHvxYifrSQewsRKloJbyk1zFC6ykXI4OSwFOj5/Ye
GHYoAANp7zcLpx7yTmzdk88CXDRVAv5eQS+RN3K4Mutk0Cm5PwlTmP4s0U+8tcyR
Iu71Qlo+Z7urTvfLyX3pY1stReOPUZWUONreGDotW3KuLYyFAxck+jgUnFpBJwyQ
eDEOXIS8kGx2uB86Grk3ViGHpMJlmLoQt8UT20/iUIbTwY0omy5A87j86Wp+G6as
3cPdx7LMS8J8h8rlSL6Mk3e9ZduCg3chFN/cx3C5IOQPWd0Z5eEKljFIAInflE+C
Vw7Wt1CyRxxGxc6y2hhB3Isj/q3xjHfgPxa3FzJBfzenC+Ud2+U3QnPXXv3Qvqhe
khsoV/dNiJ/b1xJV0Py+MWeXET3L6sTJhb8jmTDVDyfE41zkvi4JQ7QFwSk5mhxa
E0dTnK4JtBYdlg4Kw+xwBSPm8regxpvgicJUsG7x36s7dQCX6a25+02ozF/7iJ/U
cWC4FDfdCrg0J1to4xlH4xj8ryyvV/5JgMXLN3bnJg2UKiIcJayEvTqBxLXvxcqG
GMDCXCgFZEkpIbRe0KP70Mgy4RXPy4FOyfcm0Pb156l/JJx5X8lLx1xVEkgMPcaY
HLBujlrmWiSucqt7xccTtZoEjA4rh9z7nGJOl0+ayz47xqqINy0qPESsOGINqWu9
EtD7R8+huV5p5qaVBkKV/RjmPqmTwZvK0gMCCCECKl8UjnyvipR73L6PUHQoBSq3
ZaSf+y7lHdN31YQRzU/PSLVsLD8hlTSp4TvpmFPVlEPBm27aP/UjntkZ0Vz4hhtK
jGED7Tj2643iXebAJoMvJeR23XYRGuF4P7eH7LHUT0V9u7Lnn/1S4lWva7J2XI3l
SwraF5tg9qMmVD27crxy8EisIj43CC+itAoArzQN5GBRgrtNPKHzWjRuNrTo7Sy3
cLejJp15Kz9WhRpRHmtrCDKEXWFfgUXntvENjzvyOvge4UblNZS7hMxzyvNRqvfM
EMS81G2rM83I27I6WbvWXVBnlXYOV6W2AMQbKnmYjK/BPn7xrq7cGjxYMUVmztm4
OQCEo0MOC6O8EkyTaxvAZp9ewzQzgoCFP5iJZrf/V6X+fj6uoZnLcerEC3GVcG7m
AGWrDHi5VqYIqXPYwEoixo/iDDT5oLNKlf9WY2OdyB6Qp7dwJsuvmxf41lA6kkj0
kxibS6I6B2KWjioALu9shhviIE2qCMs3jEOSwJYzWH9biXIsQN4/E75bLTammxm9
q8oHIqj5qqO3bgjUSPWCBGgTjMP4OlSyzV3E5XZK4sNl7vK+kH9isUlWnExbTm0J
YyHHWeFFHy21R9k+Kw9MuLZRVUdaOJbDIYO/6gnDYk0gf2t81ZFBRiPVQnQVWeKj
0p/C1mQxiZ3JR0U9wCzVsagSI64RCtGILd1hgliuiNeaQU/snxcbC3oK2/EtLVrC
+jwtM/A8lrUtz7X4nnOVh00984Yja+HKgQ9q74bQIh28OkPEQombg2hlCSObCrmd
1OMezfdJEWXbY/95wZnI96MqQ8gzye8/iIZYD76tUJQU5tEoC8lFxW7UknA88WL5
4xziF01GtEObq0cJVt+i76jWIBcpdK9+3FUjPV4Nvh8llUcBKwc6zQ97uG2OydVz
H/yEkrzdqx3EA9kukWzfGoZinCNaP3Edms7wGai5W+ncskxXMIhmSjcMzuMtfAaI
TX6KRbqSBDP8bBRd7TXqL0c8xEw6HolARUmCsly9iO6NbXL46EmLG13B3OncCr0Q
zRrXASQGWr2LhQDecF1BrXvhnD70KDMmgkC7OjNmFF70jewrzJtWGYbD+5lRBqil
6YvnVTyouezAUvTZRuCxuwgYKjoBUfZ0EzK2BMZS3vIOmm/Bp6B4PO5Yns/TQrtk
wUNUEP6MJFysja66tWY0HQ1dr+lEuKPkLyfSNlf5MToIj4F2DAoysS5lEVeVEbdr
TPuARBPgurFxbn2Gv4q/Q/7BA8CudnxY11ZqqB7iuo2fFcCZqJOmB0hrNhVYbLJf
nW0wWRvHyWVH+HlMhr3Ni2coQ99zWDJP/3VogsENP9jYRXNwvubs/7nTMVaUfsmZ
qas95UTUUfoPdH4XO+cPsVhs72DWp+3Ar1hLCjGF+lo5wNI/PUto4WGfUPtarTfW
woFzQnJCl16VYjKW0FPYl4kSSca0rd0YLCqa5oyxOhltnprIBW98zuw0jNXSdcFN
IyJeKSUtfLAJbS2g8SvzNJReu7loVYwdyqKuETR4+6LGtkYya6NPMUIlJcAaHSBu
bu/aSWIYvONWz5Oc3DPci3pY9bQeiV0lJ6uP1hl7+P02Y6JVm/Sk9XTlkHIXxAUB
PLrOegxcLZIicrf8sPCpvCDOhmg2EWHAfvKLHOGDJyXJtgRD4RREw3XaEPckF2aH
l1eVC2NDwrc46bERl3tRb7sTDukuFLDynNTKO7GCc4QIf/ErwZbxpBNuK+qr/31G
+HQz/lnSgfUun8QZPVJgvu/PPa/7cCU4LyXKZIgtuBF/KgMJj42imz3BV11twLdS
Of4HuPKYEOdIcJiz0oZweshFMjUWfs23qBpTZM8eDvv3UuCedthkxDIyuF6rxT3a
G6KFia4Dh9wG9/6D9C2UkqgQXdJHk7m1uUHvDk4A6PZDhCX5fWvHQMl4cSItZ3Sw
3vO3WrAS/ZMNeKzrtulSUWWOzjplgk6sUk2mCXy9iprC+d56G2xP739HCnCSL2KB
fpKrwEDFHiaXo/s9DfxXye29mFZcHlCIZd7tiCz2qVVwN/aTBs3aFR16/gqCDb+v
rKrIstpgtIhhSB4MulEEGr/GtEgHD3p5tZ74dPeqgZAgrDYQNQDVJCnABhaZ2WPB
uWAPSK6kDPmA8LA9Wyg6Mw==
`protect END_PROTECTED
