`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IQb99SmiCcuSAcudiKCQgkwn+NVTiskTrY14Y+l4AETTW0R/N30JzkhCb+TshB+b
hWuVN8B5IJRh8s9xGTkK9san1Bmdr2NOM2rvxZNalNpySNJIzzPagp6nbDNO0h+e
R9KRzmH07lkLlnARSccrvUFEhrP19Zxgq7fKuSKMiAis9HpL7++NLhuhcnn08+PH
bSd6CGjlyhaLxC44eeTF2KbEszRFcnogdBH7vNn3d6FLN40ZK/6ZN7bXwEpTmPVw
+Yb4mcOvr52ja7khxgmKET/QbAiusLvZPePdX764/lPz15CL4o4TLoOQ5Yj+rckV
71TPI8A+R6MtsJ/YQ4zgrdGZEyNILH9uMIpk9idnWhCtCHXo9KZAIIJ5Le2m0/5T
LyjqThX7awtQVj0wrXxEPeX/sq0ZTICOr4JG6S3Gzm5xXGfYCjDJm/7j6fNA0vGP
yC1Jq0YCWc2XgUHHODihbYXDdvKTiENDexbvQ29nklChTcFQ+VH23h0iAuo9Y8k5
gxkhxScxXkiyZpTyvNBpiPoCLvZLTjX9g4+8q6cYUdIrRpB1wgP1hSSp1RO5jkLu
`protect END_PROTECTED
