`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+QgQGuK2VxMe2nnzTiepbTe16JL+REL9hgW2DGbrEXNyDsVXa1p7LDrUqxfdz3tE
9fYCIFhfUMZQJlZIbKN68SCF3XnTNAftqc/olAWW9og766XAstlFQHsAzG8FaU2n
s/VJIESq9r+SYapY2k4D5hCJDF7QnY3aS5JeeU7tbjDCC8xEw3K0Pxx1GWq5Le7J
96k6nB+E0FPaOQK/6sfP/8/i6MaWdiJKbirZbveG8sj9z2UYLXmAgE4W/+EPKVCE
Eh7D6FRi2g8H30m5ObZhy8oQGwP/D37F22A35x1W9F4CGaNBp0A901LvMspXy0ue
kpVt1YpBmzYZT34p9ndlu/spcnVZQxuWGRslw/IOPSZ+UzNmqKuHBmT10QjOf+JR
PJezUnJHEpjLbpu+Z9K8ml/8Mzib5VzjrdDZZ0COMvgdr1CmIS8XjWSvJt2EK2Xn
2e9+9dJ5Quulg8mqikdxOrOw+LQNrBjuv9aATlZ3qBmD9s4ojHrLJec7jRwvCC0n
04ZIIMzrJi4JP7tiFkbkglJSSCunjHbaUzTBqeBIjr/M7T7sKNYFRQzX7J/+l5R4
G2meLsYUtvY/+2QtQSIUNd0FrkmwF7gmORaux8dyonU98Cv6SWxAf0Y1JlnabPo2
v3v975J4fFqTUiXQxkr6wNHIFVRQNW6I9lMgr0xNR7VUFbSrelmI3CPQA0AcJcWE
EQ/DwQuoEfL/T+VytNvt/8kVY1PJ4N3luR9/q5B6oYAZyj3rBNz8bVZQ8LRizNl4
77eTrl7KjxVQFdrFaDAq2crrcwJPfRwxgPgo07R6G54xZIKxkwZR2rLZSj9KcZTB
uCLBOx0hLt6fDni0ZCwsrJkXHjjzaXW88hPIJqtCMgo=
`protect END_PROTECTED
