`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ms/ury+U+Iwko9u9KC9jF8SIXTF6sCKPWBiVvnxriyfu16aGthZgjQjcOCw3c+au
DRnChTfu5Ptf1EkZg/BJYd2VT39kCjX7xcP0dBmv3KkWTb1zetAmXuDfb5N8C3vb
/GmlQ8nTe+M2Cm6/hVuKxo14c6Uo8AeBpmx2U3+rd90c6inrTvPjDnciRDsKuHzW
s/dIP7aTBzd+vlCLVn4vNVNZQUYRbcJWNYw04R/60wWcIKjYWjumZFn327zx5p3e
Iu1/TQcF/xOSF9uZqVZrhkr6e7yIbcQHa8HoH2HrPM6Qyt58PGfxxJ3g021M2FGm
acSKMyGPX85mqahPlr6+Q0gEXVtUDQ2CtkvSJG/fQsgYhqfD2e9Yn39jS1cstm8e
lEsbAioMoGX5Em20JTamytL6CZdqxNiln/i/2f/dWu8FHMoQEAfasJDk9oyjWx4k
9Dyo8NWP5fxwbZ/obgb1a8tJGeCW2e+BhEl0HRk8ouHA0WWrV4D3xhJrl7mqPhA+
2OkIl9/cpASOh5mG+JbEoheuyZsnuJ/aUydF3T8RgrsuY5FW/eoN+jqnYWdiPZ7K
m5cLM9LAIrkXbzOtUP0VyZtX+wJ1kqtGWrs5ccKu6GJFNGl1ZJ+MYcP97R8YKwUK
h4PhE7fNDFAos8QFQdeto0HqHFztsXFXEBNDoAC+aS7YUDs0sNUek756uquA7E0a
pIrfNbWb/LW8Cl4f3Ih2CVOeb2P04znB2E4eD7J1zyEUW9w1zE1neyIQZ7/CN9mJ
Syp7RK0fcbVxXjVP/v7/bOyq5MJvkzW1Vme+wpXfkMjm8TYg6DIX89RKyvbCZkb9
uzSHMKqzxkesgFZf1s7qw8F+kFKwcz33UWqh/Rk+DeMHk/jyt2PRYVqpSc0u0kin
6YFnmF6wRjUt//9HxMaP02lb3yGwIzpc+p3oQJ+9L8CkL0rFtXTBqPv0B+YA1GPv
7kRJn3hCIlDqAH9VxJWLPVysBNbFFpTwjOTrixxRbJbfs1BEP/kJliGOfIqAcwo8
W78pYzXzjEn3qqDUy8UlQPP6MWhsQBVksl2GJ4FbYrlPDOKAeTmY9a7YUPwQDvdB
i9BSQBkK9CjRovUMkv/KfVoyvkV9unCPgfOyR2sIpCjLeh2TH6UPAwSQH7oMrMo4
x8Ua4Zu+nRjoN7HBalCkaXRqWxDo4sC1CGGaJzA7UEo2SdyNrctqagEkKIsOpGeE
nhux870/Q2Vw21r5KWKbABObQJRMRZS6w5lkO9ioeaY9MwFyTdI3ZdEs1lrj4kdk
zpDVdmBBDep9dTp2pYi8Bg1Y3nrwcVHjYBcILLiJz+ptPdP7VoQoSjdC7ePo7EPr
rFYuAwoQjur6SdGYgKUQxpTA4WXmT1p451Lud3xTbnkISXj/PqmsoedP5Ka3FJLY
pXdjVDAJLO15LfAxLNBbn9bGvsrB1HPQBBG/qP2vQSSLnVJs2W8vBG8x1QcKEiQR
T8TLogSz1WNe98RzLpH0MC7ctBRF+1ntxjGzGfgzjExqn2oZlYKYVorzBLnLLtj2
4l7Lj53gVjhh3kOW0vvv6/R/ihPZVA/VbcYHIMkcCgahay7v3lMy2HRWVTbCB4rH
m+QI0+S38Gfu54nEhEk5o7C/KAsQ5L7m9Yjj7BSPQLDLNZBa5PRiKNHM1NsmMFUV
ui0EoMpgvwBHFqWKjXRstk/mONTJ3T9SEm3HkJxP5t6qIv6JrZPFHug6KYx45evA
qWEnonaEvSlCxlJQlU5+EERtAqDVjXDbDirg9FEyeVJr32olg8w8HnScRanBHCDN
u7hHKktPnp09ElMSd7+RQ0oIbpNrVUxvYUrToER+mh9OXfSVXIkmw7ZP/T0yiiFS
1pRb9Xt6V2u4Is4QEXfd1NsSSfjTNg53ly4cDxoIJD7GULfwaK2uLe+M3lpQw8Dc
wqh8kadQEkBZgTvlciBt47kIsRLdBgGD2y+/IN8QhHU90SpUk9EYZiCY/ptEHjBl
7uTrd2aclFQ7GLqhpv4IBwio7xnBmFq1vFb/BSIb6EjpYSG1IcbtGYIvmNjSN0I1
pYnK2FGe7rAz0eo5XDFotIeZ02zEjDmSbMKD5eF04jJ7SFOJaCfq+PtRj9XvSX/v
NhwMpNhev8WHCXZ09eko78ttgREEc/AkeoC34PlBI81/ABfsomnXpK/F6SKEo6n6
q89OOmHR3zr8yIo8hBsmBda+iJ0LzXBu7LzpfpsAinVTWsris+EJjBXcfBckXjcJ
AD9VkaV/mnUpdyOdOPmjn4Op9n+NH78njqfvPHsySGekAlk262ZC/zgo4FMSxAwf
/L8XYxwjMlhxnhny/lCfOlMTyiaPZsliyaMruiSytiDiK/MLxRp1gmfw3LPlUpZ5
fV017NuoSwMAViYlfThlxPrIhcjU4C++94MLao8YyQT0ox7ODmJ59MxO+zW1YM+q
p6sjhrYmIYhtAiDix4ZxVJe1vg6y6MgPZItg2Ui79o+TOSWjayD/AmEW0ddRWF4U
5Ca5Zk2g5/9zV7QHkxgkqZoMMaX2+snJ/92Ewcmos1bCmUpjbmQL3eW+khCBpt5j
jXeNWaCKHTqu4ZRdsfb+133KCmcwwu8zx/j9Uu9l9ECWjBjTcjEP4mTJdmElDKD7
8/29SiM/fYnbTtoB3lYe5sKHWd/w3/f3P89Yp+x9hbWOO48wIftBCzxDaBD21fSC
BP5+sNlUQeJ0SUb7fy2pFJns5ZDXEjXrR11GDRboNCQ2uHDv45CjiMOBJrxEV4vJ
7aYxNauKvydDV8xSb0i+IRTqxmqcU1A6yLg9Ys5aza2+NgVV9ii5pGxhjWJPkvbO
F2AOKfFiqnl23OeRC2aZu7oCRShcaWNQXOaFka1oLr7ypeixUEOKgSGZudRcPKny
LoV6L99yN2wpzBNb8pX86rDjnK4ijAWya6jM4yHBtNrVohIgxycBEZgQlDo/k9rv
AQsgN/uKCxQI7VZodPIMmNvHJGtPP90PkQktvA7qOlOiQiXG+svHzTl4uK0TdBfK
3E59zFnm7SVbpulogQoEXTQ3nlPeS3z0JVg4Li+gotFcsLm9s1PIK1tVKXuV+334
zoXlK4d9H1POW8aG123nD6O8QnhuxecIKUOvCIbhMZ96xMuM+Mtv38E1reyfo6oi
UJ+1lXOJoay5Rf/EqgXJdetuT2taaYYXNv3cRpUIMZzsNtFnruz5WihsQp1E3fmp
FPJh6FttDhMSnI/ZKUx7IWIE6k3w6tiAwM8h+y/q4Ay/lczkAtQNDX+TeXvx4VjZ
S8Yd4lUbCC5hyL7aGt9dlRJEOXW8dRjGKcNRKkmaaktoW7ZS0yQFZDSh7jreuFo8
Z5M/1Cnt17ZppeFyzhtb9bzUDVygLMWEAAlJRM90cIdQnMQqLCEEOqfIxDPXnhF9
KThNI8KcQFXrafKPdkpDgWadR0XWPbHh3WjM0OuAQ3tcC2miuQtKlmw+dhNBCyoo
BlDeJVhHlOPoN0DCtPWi0F2p3Uu4AQPWK08APEirkk6OCpyPUCTM4B2yYISbxFEQ
NW7VUl7GLExytFT7dd5sRBiYEdDGUHTN+fDIXB+ZSA/oGAjs7gcM+RVcF5l9lQSY
NlxozeBa0p1wQs1sDim/IGNs4846QCEeY+ETZfGBte1dNwd0ZEJNyW135/cioOiw
mIuve6uaOeuVQ2g8XY5m+Rxr5gd6fYhWWU8/QtE+NB1yf8QuoGzixW370+lHNVEv
vfGKlVaBHJdswbd3HFZMCBfHgClfpVbN7GBZerCCqUu8dUm/TG4NVb3337Ubrde2
qNehGIyYJmsyEDfmvSsusn6RnpUyW4EFtVur7Wniu1n8LDlBlExID4kx7fSjzYzZ
qK04S9DCbM/0DTeXdk5rvphNLfY3b8O6uBzFu8V4PV+l33Sg9kuvqerIlJ59Re4V
rMaviTsJb/uKEQwXb3kMA+Hs9RUZPvJOP6y8ZcpYK5ChwznVACZ/mMgCTbxLNtT4
zP41Gy4bJs859wYfXJBnZYK6Tay6TP9fmV5jp3l2zvze3xPNiC8E6/zb5rQN2w7G
ZHRnVK4PTa8sUX59OiK8RLrUQDCTSHBpwviH8bFzFzzKYSBUSLw2wgjuSBk4ZvF6
cV6UlikKKiVN0dqsbCm8TF7oLAcxu+57MC6NnLWQd5PYBJ+QtikRovc2DQ8qCkB9
mejHNwMxktfbv2aUb2SL7+2qQ9KuwmWIIGACkM4vNcgWEYaiWi1Si6K6oWK3Z580
j5zTJXkzAiavXk/jL8wW8QqzXbVR6bt8zopPmMUZ5doIS3v1xQwRccR2/OxlW6b7
W01Xc/SZOca7j5KwlGTtEe5Dc6p7WamQs8jR4Tmr0np+26RNg8WV2sxXbBDwVGhg
5uhZ8M8GCTih2RzgHG8DuHMzyPzLxubgAKm/eUv5irSKTVPQjDiIQ72YY3wWNYOG
VpETnBuYA8o12/XFBspKl2qnESLiDivurHrC7qfYS39MpnuVqEJBRtrO3TDny8Pc
sCKHm0L0KgKd0cjB48WryVDqqBqIJjlkawklXF6JI0qPmbpyd+P15+T57aa+WZHZ
GbSOX47MCOBFFx5EkS/Eg3DF8q1xZCOMWTVm0ghciHOMKoSCPK5l7e82DjAfEG5H
s6XifcxF9IWhmw6N3PQIwPUlXWMNMbVIzOXS0J5DJ6BxCBw3zL+ffAX+ZaO3bFbq
SYzuN2jMovmMRkgFHDy7LMmWpaBDHwZFdPu0J49SP4EZdlsuqtU2PHvv04VnYgA0
wERa61B/JPovHlQS0xEhrfFcCy47QWrw+Djmh6gNsfFDQhSPGoI6yP2XUew5xzwP
9EjIPXF4V0Nid+VrjvHLsTq2BJnhaNBjlYmo1b6utjHjoulThCNgNgNcggnBwsPy
JjeQFnaVKXwxsWy2P5aOjxAmvKmkNvEK8DePHFmSIJXlmmCtV+OzQ9SOuGOLI9SW
iqy0B/KpugBkm6lVSYVoXwcfQRSB6Js/xrkkPaEmbrZK4AG5FmAWYDNhP8x4H4Bd
9LHU4qkXIXy0YLv/gEnMhOHTlL6hykypwJUzcfNR0jzFRPE4lR27vJIMTe+8BjMX
Trm7pyiBOL+oXZIcUvdZWesYzq6wOQXO8zYUD0VAKRGa2dk9ai1Hi2Nvr6r9QlsK
rls941DTZBuXL27dKWqJNbMS+5G2n4eqNo2A6OQDBHp/hNvqDIwFt+Wk0V+sX4Ec
noI0Nqqfli8r/lYBdbwPG+Msvor508baztHckiHeYc4TO0c4iDbh+5q6FLyILspL
wFsZGQLoRc43D8TFoFTlyUQJ5X0LmBhu7ZhVB5bv+t0HxedefX+B7COqjm1qysh9
9v+uhdzUM9ez/c2crto6mFTJQAQUYFcUU23E7zd0EUPfa+cDjpXhMO6ave4XTQu8
3Jc4SO/3NXc6m5Q56/iEtC8e18CDotNGxtdXNcW60PkJJ+9Vz3sbTfwIdkw1wu5Q
gXTBdDbXoulJROGAkbWv592TaGF8DnLV3oAyLrcMcmt04fvZk3qwApD/8tlya8jN
Q236TrVuYDONZmS/i/Vz8a4ocWcxmV7LTLpb43HeI4pRk/IZ4f1nh5Fn7cR3mJcz
8tlWH2Pbj70gY8oBw/m3fI/Mzjf82ksXgI3J7KTD38hJM8PnaZmZDjm3UPGrTXMh
ZdVHGbaope19/H1GuUoTx3kJKaMkplxHdh3BdEhyl6f7e8iAsiIWSXqBXdAuDAUJ
qRTuIqVyQ8Nr9JV9dg4/IHKzcJRJLvLE+BpHCyxu5FPUhCqXXL304MdPsWO8UdIR
6GaNErBjK2ZTfsCn1yrFuo3NE7gExNpHkWHFtS4RVOgxiJlueh3JqN94RHuyeFFW
dsL6qzez0eyX4dM9id2+sJxFSW6rgafv7RnwqQBwH7MrW8oWDTOJ9+GrWSeBBZxZ
mdIGt5BnRFdn1fL0Wi/OQfUFTqKDGtHx5DcOyC1Fr7CkrzHcSE47Oydl8cfwk+Nd
7fowHFWNEvkrvFqpICXQR5y+Z7luXDmjqiXkjx4XqNaOolKD8KXxcY4DYvKPJQUI
O4QEecNcOBAfl1q+9lHyIzWlNkZT8vFJxq3ZG08xpaa283bRMqGZJ4oFfLfq+6Ch
Upji334MARXeLTo74AV3zUkdXIZutLFvmucFZollbiOxrx0AEbX5Qt4SjyeA86U1
O0EDy1iTJK4erTeXaRleuMAW0CnpDpubovyK2c7W4Wd7CiPctPkSqen/9acFyGHb
BHVKl9F3W7Kr/HS4kb4vklXBD2Xf+a0JHcayUDThVDjIP9Hrhb73SN8MRLbtzBEE
pBs+fwo2GTgDsEyNFGYNkuq6G+SOhQiDUwQP0f3clJHJnxDynwnq+WQdBHs5NdaJ
T41fnNUtV2jCuYa83GuFYOi31vX5JamO2WJcH/31t1mlNNZNK7rN8hLWRUS5cyMf
7KDtXDH0lgqLYCwFaFtfdgkw4JnNgzoXrecqOP3x4Xm8PiXQEvX5xkWrCB6FXS5e
4vNeipIt+oEO0meoG+vNOzMZhIgLKRhF8ZLBflPlIGyxiTbmO7JnqTgNNIkcQ39Z
4bLt21ufyIKjqzKA4AuD+xPfn5RYr7Knk0CsOM74Q9CY1CiVV71H4FCREAzOT3mI
5vchwgvM25ssuA7HIkfbhUrGD/565BtqIfkdFuaUtEDjDoa73ncvQJlH3hEJMrMn
fpYgTwQVusoRAdsqzK8m8Q/774i3ISLyMqO+aWuFTWM3ldK+CQH1J6VUzf3zL75d
Aj5p0jWqO8Yjuwsg1udOkApOVgSacrPxZZCxn4bLNx8TqS2PMpiU+B5TjKFEc6nS
Bfr3pUYui9Ceav2pGG8//790Bh0CgfqV/dAOW+ftYhR3lfNMm26JL7J0HfDs9aYz
IxgvqfHiXDCqqg1OXB3SxvJJkERS/6Pzjz0huMeOfWAvq8k6fZqMusvI0AOz1KWT
Rbh+Rn82iSWUAcsN5Olp/lZAG0edULtEyV2deOsEdB1GzsADDcMlN7y0zriyF96v
lVYYb8z2CzuhEW5F4ZGE9Go1yKKadi7HG/mKsLLY5uvwmqF4thoKCIBVX2OIOSpO
EPu95zVQjj/eKgJpfRU1Dg/rPRpmrztk27m2E8F+sowYyFkclysvn4LMB4wfdmPL
x/szI0dSaivY+b3M8DzP53VTSzJ8IQWuYxpkuLmrdBtHafbohFZREi2i4IDrZIbU
K1K8sIwXLemkSpraOEbqRScjZebMoBfZvLYzdbzt71GVXqiKHNhlA7h/wL+f134R
OqzZXi6diKsKWZOvLbY3bcIx0tfHNi5byFvHlZ+Zr5i4+ANPJVRSa3V/Ku6fyvOw
E7eFfchgNp8Q7gDkCMM+gHg5f01OGbDQag/jJ5GjVvQbYLIO543SnEZGwGlXW/O5
ivQJYHKvgJ21aG+G8rsT1DsGNKtjoEqGSBuZZRdq508X+zplQXhCpZNk0M3Q0fy1
9Grn1vF6Ap8EVQ8tCUU0+S4fdKgCEH7viB2fpWidIlGmXBBrN6pgpJu3ul+CyaI4
QZyVFC+FR70dL1BTKWnZ4JcFVGFV8HiOZ12rpEV6L3g0zfn+xjehypvoZ+eWSu/N
0qQlEKinO57YQHLyn39AoEbWmuNuHfICsezXidhjG2ogvA/bSJtVZF+DqmI/Vtt9
ZWUxmZPPfT87OeaIeL5+LTH5G/IgIZFdzW3UvFW87Yy+MmPmUQhBwZHhFRO4beKM
lcQmH/oNYgO711Ija/TVhs7GNAtbKEZOoJwZkCsnvk8+2KiwKzmZBxwwg8I128yi
eZTB88EHRmSU4LQvl0Tsn2Yk1sQzMbsUjlnjUJ+0OqyHydZQQZb1BNwXJtkP5dBl
ltPjlLb8r8c5pcg5VeXC7o3fSyxi7sQ9r0mlVEwklv0B+8NNsj8uybEJqvWe4im1
Rmdvp4g6vc2oeTB8iNFQpoBA0HBo0p3AomqLVuFiaMkzIChsMan7tJ+48XMLHiGR
7W7jvi1vHRYrnfNjd+ttck9F4ZTBfBe0k+rg5WM+dsZfmwJRDWGLTNhqrJrZ/x19
iz/yeVlm+nP9HtRoIL8Bd04XJb3TA7uCCeOyoTio4UT5KiMQ0XDKbWi2UOo2ynH+
QorG3STLzf9rqxr64KpGtlowiWJWrwlC3lZdAqNcRADV0p7AMHUmSEuBjSAm5ej+
7FJSLD1r2T3GGJtN3Rzr0Td/UunVXdqM1ODBNMBHJ5J7UpAyT/2gzwlqJdVS0wk9
53TXJeTfM0UQCvqfYo6y1ieMFEao857RdyT/mzVIb+8MoMH7tNeoqWcbupp42ksN
vXEq0wMjhfjwpWMs7fTvjK1kkrXthd+q/0vFtY+liZgBNvNuEhH5ujZfOSYWoTKQ
4Z+UYashuTpU4ZdPxSkYfOQ6Uf0hmgS+66AV1a48Vd4JChclDtKrcGfrxsZSMwdb
EwNzyycU+2GmCHRAa/hNFrhWRvV3dW36GoRiXe1Qu9hy5uy9DRqTqf9yRCozSkUF
iNbffg+IkiDr+blNGnV30h9Rjva1FZGrK/PxRDoJWKlDTAgzNgXIYIK95pNwtegf
2igoVUPLUKcC8teiBV9x/JeNA/U7+oOSs+FHKec7LEPTttVTzDiwhy9iBJsjRY+s
049f3acDTBvy/MmN5qm7b0+lcvyVz8c57ez8l/R+2vDP9Z4nYdGVf7tKLv5uL4sg
y1W47Q/XsagEES0p34oXoQUPpXy3AdmF+ZP/Ps4eu5ZRVB/xUhi8IaHfKzIfYU+X
TIdjCQnVwPuqhUnLHy5aARBaLfE+9BmlXBh6KlfeuHvIEvynQoEE8izUcEEmv8AJ
J3buKjbrO867Cfwtq9j3WqVcv12TOxeCH8HufvjBTvavevWCEGYTeRtIng9sWu2V
gELzMTfTm2nGsdh/utEuqlxhETelwRY0qRwYV7B9U3uH1IfPzPEdrKH2mNEs8Nd4
PcpaDh+Dh1e8KTVh6Wljkp5yAgYYILI3IkY/XnV/sF7zOQkThMCrfybfb9l5VqhS
x3o1N9+tSQjXYXeBTjdxBCqgplrJPdRWJ9qv/+moM0oQ1DxQN9nljJHMjTq/qlf+
vv3bMYQfHGFv0wYJQddIfZa+6Edmw93ii57fUMApLx1XrL9mQEwWEoyHPlaU2fXP
ZF3MvBe9Q1D8XyPRIjLUaP3XQcHTO25HOLjcfpfKMUdSfFs3xI0uoXhZNEh8GQDP
9dPvAU/1HBj6yJ85QHyy0I6SHvsEUQPe73UoVZoJSCr2vX3oZLUspfXRDZ0FKI2a
HVtmrixa21W9ynjEjyxFzOynk9wO1OJLQI6MQxDd2RowZUGpabG3X79E3cL1zpuP
PfF8xzywwxe2zsG0R7cqka/pFy9A36Lg42bli4Y48xaH1ZEXpgDuaz1wgt4DJEBs
Ri1l2wzTk/9LGfCFmMGitWHE9j9d0xa6Up6mVEwVQKDpNArT8wAsC5dD6hkUHVQa
ZBJ5eVGxu7Y98BO1LWen89NxFNPcp5BOkbX5JqPyoBSo5t6UWRYEIOeR/8+p3LqN
qCb8kxoDpkC/Y+2t3/tt90d7o8SvEUmRlOOBH8GYxdofNDyTpT6Qr+1mFU5RYGYc
GgNGrn8M8h0FSSn8uJAuhJZ00B3aA6aDxMUnL0tJ0SwXRx7s1XHev6V+PfgeUmYW
wkUm+fQkS6D+YGQ+tjBFUBlouxOexo/n1O/cjYAg0pMDV+DUtVaN5eL2SpfUgZMG
a+NOHorTuLo1i/pFjKGhKqKpjrurmgiFeZ359vyq8+mBiYMqsg7TIZ7f2WSZuaVE
XVfS84/R8ToYZOFM3BmZ8Kc+YPVPxbP28pz0MTxtRaGYPh/W5IS3zOF8Y3GL/M7b
kS8kN1w+e9V9b5uWOa93p08R64V5ypJoSmoZTVpnqoez8H0kt6fCAbO6anaPtHr3
NElWoWPvhdfvDiNqUFLKlR+2zGTNt+42DobpI1O18ygw1WEPEut1dWJ6uXkPj4ta
CuC9j8u9qJkLtccYGqAkrIenDx6rvQjGz82X5gIqeCewFqrfu2dlxHmMW80/N/tO
yy0mHrtDJrm3HwtafU6bpTn1dBNEQL+HBzz1n9/boIvNrtG1k98TigtSWS39cMIA
fYa4ok5qzTWqV1CKmPyPsWU4Itk2qnSMoI70mMt8tn9Tw+XBOyoHXmH1LuUXx1kL
NIFtTMOXHdAEcJt6pUi9DDQ8QLRsxUYnOU8KU7ZcS9AiyG6QFrbTk4IeoaaBOlex
vR2oJoo2gTfkADfbXp9pQsVwXMYPHtYsRHqn7Rw5jiY4tkmJXxJCEj5T7NayLm3n
NphRVX4AA/k/0o55CsxPp9Si3uOnCrAYTQJY1SPWqXsaRFC7x7T42kBSQ1jta58o
tcIkqWvp6Ng5qOZ2WFwAsxNNPUOwzOzdswsDPOP9O/flYg4ghdA+orRz3HZlgqBB
f7HciQZ8PdD60+VJrT5CGnCa3qNkPzbwX8sIpxg3zDnMjY1mDIWVsEWFPoKrrxOo
8A/sIGEZVn8+kG+Pwb10cjzKDLjZJGDmCgzRhkrehSEwnkotCg2aUxnc+OwleHqV
rEVv3xSrzJLjpJ6rw+2N0jxQ9Z6dinm+RTzLClV2q3YL9zsvRznO8tsxvbBe6uPM
+4YFXd/RVPZc26rJ7I9P0hbUaiGsc9PSxvAkDfh3IO9An6jS/qsC5R7cloZJdejy
AXjYm6EWnb0h/7QvDnxPflmtjeqIic9pPBG8owCckOpdoEsvKdbsdi2F1ILhWyLe
uNC6CNwmawodQOhtKkhCmr2nBb/rs7Z+JJbMCHqTdc1kq7AmmpBaHljEYcUqXpl6
eqrDwpvqPwHa3qafH/6+CwBhqrHZjZtA31ZhtyEgS4aKAwPJ1eFVbQo+HsAB7zA0
WdW6xCr4YjihGpnpNwzVrde1tJvIIqRQQQ6farOlUB9XiYx687DpT+HJTMALKRoZ
7vuOMsQ2DQym5T5sEablMrU9h5Iebsc2fDsLZngDQt5pzkXD/TweRBi44tWbxUqd
KHqdgWz+OVfgaU5Z9q5YzN/OwXfMH94b+pu66r5Dk1PqRI56YpTydLM0ZmooPwJy
Me8cpRGsrfTY0dXKlrF45w+rEqQGRB67NNHxJPusjEQH08v+TbrA6Jm3Z+H5LEhI
KH/sTMgLabY+IOne87TwVkf6RCuBz3WnSymBl9hw7jXIj2qvcG/f5WH3T7h+nczR
+H2iMkVpW63AW1BOLNmYZn2q2qKIZ9p9K5AOUWq4JUu0+S5c2yVxY6ebSTi0MBx+
59bC1UI+mAUGS6bUdDIu5m6hJbFvbiqLTPlPXUWPWsgi4fyNmcwqt0TVQ8HDQAWi
f83MNoQK6pbsCV0vl4lyj+4TCyONYFSThCueymR0jCMRPzm0cuAW61spHeJLfn6u
2eU/hpelPnmjW0j7TAiiPJ/e060Hy/2SogWE2FiTM26j/aUqOMLZtkPUAszyNTk7
CI7QA3Gt76fv6eY8qb6d+2ozbTn3QcrSs/P0Peql8Zc07BrdtcxL6STWheUGmfaJ
RFOigeinE0iA1YawysoYPqDNntG+JS/ZZ9Hp34tAkZuXZkFV5lfHN10yQsh6CGq2
LXqT5sIWp3dytMsliMwC3qBDmsE/QhIO+Y5nO3brnHyv22WKCw6FL7i84HEpuvgK
YJJhFb0ztuaRjGDLeZsKn4doLfpYX+F/jp6Z5h+2Pg3KQuLD5DWeIqZ3NazEuoXA
LtvHUvtO1FkM5RLLSKKnXShLUnVOzrYSe/H8upusdCOm6A88rcw4Q8QpiEENIPu+
+PJeV8+zrrqrn054R6SzOfQhAEGzhdf3JIfz8rVs7r89KkTVH0eAgAfx/1uUmhg5
iod0g73Fasl1YSxEL3PJ1obhkm+aZ4pQ0Twswwxk3hxZc9W7di4mTCtJrBLHA5lF
KXLt6NW+EJOdKlWaA8k3V5BCHhvU2BxAF2r3X4okkYPyLWOZvkr1SZ1kGMKgzpa3
L/JmjFSs62rL9LAaYxbiAlULaHYSUg8emG19KGAm2N+3TaNSo4v6FcBIxeICBRmR
OpmbAya+QTZwWrAb2kXIkhQxPjStX8NnriO5jdH96wTNcaAHo+YkH+HkAkwTvV8/
o7UHcPFq71QyD10/IetfY3eipXkw1su4KlSd++fHTWRLaZ5s7beqNa3mst2G7is5
G/IJif9N0xjLD4BsnJAlWMlTcL1Cqe4SaZNdymienG0ba3HWqZyNqo+kI6qZoOIX
H1boWsO3ozNKbiUkQkeVfIBq5VWOr6M9emJ7RfPpqa18PE/yJh4eLhlG1iewRSkR
+O614nB07lCtk/nOX7CUj0nsf54w3gRCETdX5OihMqTZVSIgdVx+mUwWPlXuay0U
SqxSLKhc/j7SUIBSjzFyo/M4iHGGvMmtfzrvAKkl4ICwUSHX41cUeNh1Q0eFxzTi
0nK/NhMKJr73AmwHj6fQoh9Th43j6vKYrgDA/IN00f6PXGDfQh2EqePBN9Jatl3e
KSVpQlYVCs0w4RU6k7AAbOyuBBRWr03gM6iOhWZmN23RXGIX9IrvnsnHMiJh8Xh1
bQ7B1KSacsYn3a6jZOKsPlzD/hZlZYk0pFXwLB1TQzPp5Vf5oSAsF9GGhmNiko9x
hDKwLQB0a482lv/22QwttvDR6xi7CamiJSv7N3s7QDttp26LyjtYhzrP30ajPYnC
R6R8td09cih2s9fsBZTODIY7HTf6GvVHMRo3hCWxTVTOKfnnEel1mDj0T4A13LGA
Y2Bp4z/YHs5vsZzofUiXoVucsWLVfi2+Aia7NcTkVMPTY7U27D2nz/UkdthoXdii
m5JfCtyhehU+vSIf18cXmre07b2JloASboyCJ9bNnF4PHypoOp4OAbnZkEWy1X42
BEzsGiWuwTQAs7bGhrVicuE9cWiYO+OcedWiGrczAU6oFxDLD/9lQJL1/V4nEPaN
FheyMsL+LdCztak7cLDZppXcSPpifiFu/ahhXvbo6EU5qJred5VlR9JCL0g8K3fv
CigT5zT4zWhjBn9Ifcidu8amqUjxgE+WOPvZmKMjFuzogDG9H+byU+Tco33g476w
Kb2/9hKR68/A86qw73gxWvEfYfOHkHI9Oz3yfb+fxvZws/OJ3stP8bMPN1PFAckL
PjPi4UMP0gRaKGZfYiao+wCR+tLw6w03/swWLec7HOY6prNJQw1WlsczJnGjZ2vU
QZM9A3x4vSO/XweOYp+QhEILTbcopZwJNJgI1CMXMlWyuHAfC8qTiXXXEx2JDgtF
SSCvD+iPOAU75IrkOBOqmIq0yMGzjwn/HzlH53U98W7I5rdBjz8EeBIqKJOXuUWl
y5GyosVhV0vstiqVhgYINIe6skJuBMK1733iL6Qsy8PxGS1s4/8F2133MIvHp+l1
XaNlMN/RUbjZqJzAAdLf9jPPJQ1GACkeGSFCCjJ+aTbMjY1VIh1/n+sSCGi6GRhZ
NBLjLmUbDreSvtRiDrMgaN+dr1UnknyZ/4dmoLyFXCwZPKWCqx3vZXLYOUDkgS4A
SzI33jy4iJblwQg3hpQ0M3aNO5tsUBxolXbj+5LuSBQ8ekn6T0rI2jzJPV5hDrnt
Rwgi90z7miaTatJ7tU1FLvPQG4asE82kYtkQcuJRuRHLWS5ny4SEV6Bky8LL1zsn
Xte7EvogEec1NbPYAzD7FHdHTiA4VyzxLFJ+B6Rs0AqbcWYJbEHP/do4Ve3SbvRh
c0uy69N3XBsF/GOy0afRtKYAgJhdfKwLkIv/XM2ey9I6POTn5jbTpti+IWKlZ4qn
6AlWOMcvIJDiTy8lhjRbTAofvdG7ekCs5jL6BVEshR9KKhoXo9vdIohGZY1LcxFa
Z8LjUn2H9bEm/RPusp3p2r3Bg6Tx36eSurHCEacq+Qm6rajOFj4C+yI/elhRZ7WF
kMhxeyPCktuyMqyz3bBELWtg8+6dhV5M6PYGzBpyoLjihLB53Cuq4W+ttm9z9x0T
7rkmpnUmq91dwi6x2XXSvoeT81tERFHJlv5dFBRRT2ZQL8+4Otk9bSOanyJCMpy0
HS1aP9/G8sqS69ymstalccxyL0zE6Hbwutvox+Gx/02PP8wDR2aAA/lretAne0pI
Jkn1g69vQqUCi+S/khIUUCtQFyPkoRE9Fg2qr9jVM5NPVZBvk/JUABpZN8854M4s
No+nsHiAfQdkFabuvE7D+w==
`protect END_PROTECTED
