`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d50IVe66zopB0mO+84+c/sSivESQA6rwOwrWLTx55JKPu+B3m578or5PT5sv+r5E
W1L99XwkPoxIVmux1BM+xOKIDp8U3+dPtVzxKfWszIOQ78IBx3rsgWTBxNyAGq9K
5qK+6SxLKkwHIz59Kmdtl4+Bg/eF3FhZbjD3gictcSdeS47ZQc4TPlsAmJ9eCbnx
Zynyv/YpKMhZ/6fJVJswxLHjG2K0JGGb5fhBV8GTkShgZJr/8mnkm6aTZeMsrMxF
EsAV3ZNzyJLZFWR7YmFDDv9Z0+QcNovR2fx38Bjy3sVxpZ5reIf1+kfQWP/UoPvv
JUtgW4ixAFa3vjH0J5rSnEZlaKrDoqp/EYnX1fqQWOJk7EA9CArGfKoaHsr/14tq
AHldBilg/rq/YjXNh6/qJolxYrkEtcpJ3Mj6PJIrufcDInhjRGNV2SPJTN0+FC4y
oFr+6D9GoQLVTAWJkTRuzkdJKlSs98QP+8KGaJ3/Ty6ObGHnqGauxQxkgEnQ+iG0
CzH8mEkoFORSdVK2CCSTVC+oQ6mNfbwHYYI6NWvAExrNNn2SYLSaheGECfVEXkwQ
WG5vFLHzL7LmStnilHunTkBcDN7vpEAA+Z28pVTaeMXUhuCV5Jh78myAD1M0jofg
cOuDo3Txc/IVUNaJKhaaeLeWvhujZFY7B7qMQYlf4cxVPKl1Lf828aQkCR2ohoju
ZR26/9L95V0IoilII2xVB6fzF2JdnnPqvS+a25Tg9koHE+84m2rQvhhHd+8psTpz
bZ1EOl+aHC7tiOrJ1Ni++zJ9NAj/ff5Eo5WT2VqPObSHu5+yUP7KyscGTC5M3TGU
HsC/Y3gyh2ZCMKvPYCG7I8IfbIwGMA87MZKxGkr15WIJXp/bA4HvyakjR4QC+0cZ
jNC1wQBvIF1aj3K9CpwdNxmUtlYkJ7S4qa5pqRBudNJq/3YFhou8T+GngJlfQDJt
Af1Z5JlEki3jdgsbbRB3QjQ4wpjt7azcKWw/HIxJ6nQ7U6vzKhLl6coIjUNXO+Z6
iYTX6hAP6me6cz6ldxvzr5jueW+NxYPaeKPbF4RuMm600TULM6lGh2uXL8W/bzB/
QAqZ0ENPY+gvUyPDltabGm604ZecDKfLwFqtQm1ZcR6b+kNbS18wYDekkLp0DHLP
XSqdKPiZFHH31qFOXImEUJiTFLYl/Zl9aeuXreV96VKi7MsA7AHgpqUPxQPU/cQT
emrAQt4ztntr79TnMpnBxp2efRIgJhgRJ/xLlVgcNPuFtyR0vKXqjsxObZQWQX+J
mm2y+3s31EFGbe3L8txk1KXUicJlm7i4xdxGCw7sj1iKkcJPlp6ybinn2YTSw15z
k1Mj5xIQhDZfeoO5nRqoqMAgWied8ZKiP0PK0TtezrLBehyoNPEYjbe3og8Y41C2
uhM94rvCfkYOpxjBQ+VPoKO7f35CFomvK0BKrBSfDAX3lDgrWY3SpgTrPkmkdDH+
UlDuvxKTUVQA/g/9EyaKUywBepoQ6VvRTKKiyNRtLpXy9GeViXRen7/BHVZ/QDWW
9iJOnZCPf0hrKtCSMknNzv48vgYFF40GZ13iczkslxE/8LfK11uzbSN5m3nUH7at
RY+NJju9v+f0pTniXXWWtO6rah3ASsolQtJT70VJsAznTjXRmLs0xA9ZMbmRA+yM
N/yeeRuj+/tnC5027EFh0Q==
`protect END_PROTECTED
