`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6a4YsobSZfuzakTjG5BBUAS+mObvWa8+lkMqm56vHDEEkD3Om9SriJaoW33crpH6
ByXIXBZfVrBKag4vsi4QYiUP9JMl8FreohKPVvAoRYDUkbJiq1PixQznRRta7Nzr
oDXfImcqNO0Ww8B3HxFnaLShBzUwx6b/LA7XbuaRr/p3u0sAMcOArqv5XrubZ1aC
ksZgIJbBZsA8JP5ET6MnOmRRHTo1kT0B+nuAlPq9WCiRRaoyfSMkFBaUMdVYRdEV
5pFIL+RBtOoS2sIQ/n5zRKwXruhVSng5Fnwr7WkzaCRHHKAyfHTCj8SqiLmZQxAX
6DynRHDz91gCZ1dbhvdLq9ergZ1Zsn0EhkILre+Bg8UMEwzZRyMMYsAA7PXYTRaM
KypSD/SoAHusoQvRPmmGx4tGihxmznmNGcySrgmpUGWnOOST1YAj09T+9Hp9GVc1
70jnILFrZcIt9LgBd6eq7v4z86/zaYW3PygDIWLdl+17TYep4h9f0zSliZrVcO8D
k2gc8CpkDZ8Z2Mk+bJOqk96Dz2xTHMvJCPRXmFQ1v/nScFlrBXy3zk3RCCPIQhZ9
h5DamdF9Ot0AddsCzMsNE1DjToRVxereN3wxsXx6Prk=
`protect END_PROTECTED
