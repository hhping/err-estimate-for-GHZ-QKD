`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1B0XVGqChKWQUPpKk6//rncRCehkYRub5BDlDzi1GRSY6RDG4lU8OUuhxIYKd4wJ
uM8ifQ/mMTVkYtXVn/X0KdL1wS4cYal0B5x3p2cYtmHZCkoQygxtdcXyedbII4Ad
lsD4iKim/BdkGg0OaejzojeVwG8x5qWBMeKHJ7jHxWnv7D+SsO9+QMExjiQQcxo7
HS9YzMlfTiXJB5OL+4cS/3qys2xffVlHw2/mCIeHl9EBj/5kTTOUy0g3P0fE29jp
bwuG3Vki3QPos051pXJcVRRCueptU1pO7DArTFOmY3UYO2C59e2chVRYuLaAoW2w
0YQccmHvL4tnnyomznHNb20sDh7bG8kAWB56kcRM7xX+4uqGv/zsrjAIwI4DOqjV
mFY1U7dFnArhBPllRloQ6GFEiLEdBTPvIv1xpIB3/aGqBjXrs7Rlvy2j0VHuXqwC
ki4GKi2q/skD3siI/pI1iVzJ7vrLiHlRoNQp+NE9KO8rm35mfW/HL5flXnXLoYBh
uwl+TRmmavhy1xnh3WN7S7e1t10TDzlYrcpq0vvyuz8VG1sg3cZCpRsjdIFK3/Je
RbSB71l2UFJl8FyFIbG386Bv3jrrHAqT6SqiLog5MQGlD5aJriV47+7gssd4Jrni
5fPBhGgYoDyG5fw4RZQEXi28BPtPg+mIaOUe2Q8lQJSKtPBaRCa7e4KptQWqadId
2rMuucFu9Fl1eZSuMgOW7w==
`protect END_PROTECTED
