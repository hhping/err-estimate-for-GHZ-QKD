`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
etGThbLtUDmOW/lpmjXaTN+pdfXxunv9bdgSWqChvSOLMOgjWj1BleB+9hOo5UuE
zrs90dPTGICYVwPU4N2lzUaz+W0l1knScMI+vtOkZLo/m9vGSWxz4rqvJpLFHaPI
1v7fcggPvUobAuCpBDFQPfK1Co1BMNU1phZfggho+x+3+oGvY0FYYn4f9n9KjTIF
uT3iLfUEdqxtfPZYioobatNoJU+bjVDeozvttueYG1Mveo2gG/ux+fpPO1ilj2z9
YIVNCcwJAX3SphpSoM23qAo+54db61ubtQhEyzjXxpbYwYQqYZVA4dHJ66pZet8j
r1OarMyqDS0Ew6EQ5Ly3VyjqjlXbi1ajQ5jtiOB7liVygNSgpExAttP7ljPEQvF6
O9tsyb8CQhrtwkH2Ps9cEDftPEnm1nxIaLaN0tzd6oyUXCJsH8ELwJwqs1oYX/Fl
agV1il9xJ7a5F2IoAQ/nOHsAJRVtoAmnFh6bcjg/dCXrKkSGGY0soVXccoihNWZu
3gq/umiuQ9eBlCbYqPvLpjAw/2nUi45JtcNTuhyjfcdQ8XrTq2feLi/XqRX/VaCA
cR17E1Z2OVB1Cr6x6zMmS2b1iMdTHVScomx/3wqoC/szw/yIU9vvrHlJbu1m0/if
hjaytH0rwCvGbxmi/A52rBUb9GLpRTb/a7KVMFQtjPFERc2lkBBzDW3VmKpzlET4
DEBA737WqNEBUVgjb/AfgvucexHkR+1jbkc2XiaLhMOSRw5vT/K/GNQKy2ixY+Om
jnO4qCj6if1SNb77iwxghS7bQLotURgpBM4ha8pefjnOFrrjMrZD2V/ZYn15sIut
gitbYJKGJRx/VqgpAe+6RqapPAuWajV4xzGVkDbhakHDn8F0K7R57wjrM1Z5q5E4
zXWcLKwhY3GAfUX0JDg6nWKdKJwgQUKMrsDalg5s/pXYn8lYsiQuNVRNIwWpjmaj
otHMEmIR7j4JSzZVB3OLPxcB85FG0NfLeA8oEOtbDROgkV1mrQ0n6njA1cxMBYmV
IbsRCSwawKtGYxsXe1p/pBXEMwXCCvDGG93KT8AYKgkOuQKVT7aghF1xJ+/qOwph
LI5re/1q2c2zuTcrK2rqO/gdnZOKM4qqZ3LeHz6yeK4CxCRyHhw4pTP+J7Vdw/Zx
VrCmPevPinoq5I5CfclVPOD8OGTav3KoQB6Loxo2BP7aOshhT7Mpmv+rrRKfucZR
d+VQgEqm1Bh6uP5rkKGYHNizygy7Zpo2//N3gh6wOyuNM8wkt9h0B+2NFpnWodbq
xYtQKqlEom7pH7Bi8Cjl4OZbpGdG6SHSWMYSm9gHzs/rtjPxa9Fm0V6eZ6jzR2Ro
slznYM7HnlnigPNahqO4+1qhANmy9dauxVl0/aBieFOjOBTsdc0GE/zHRD+X1ewz
mE3LCgaWQKCVfz0fodnJwgS6TDqRWw/4uAOWA+Nubm4d8/jJpkgiXHpNf/EerXqR
4vF1NsvZBkgUIEeos0LQ5Qt1g9jhtxoDZkJJ3xwm6bNEK1X6dIdchIT1OX5Dg4ii
RBNf2LNb2I2aLmPt8hJJtgVl6FbwU6bgvrXdoJO4GIXNs2FmzuLILhvZBNXTGvTj
ooAeFArjeeqrY8c4/EVUSafWhtDA0zHVaWFlg+8ZlQc=
`protect END_PROTECTED
