`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SVHBBsf1+1yu2EdL8HjwBsP2FdnQne7keC+tZxDPof444sDckxb/DnCp56fYpoMq
NXdU6rGQT43lEJN/nroiev0+ufr5OGsUmjHq32sHDXhetzKcM/lyVwmpxqYYkeUZ
8pbP+shjraOl7o7PcsipWxZH3gOrb0EDimNwTbtJCTjrQuOhV/J+PscNwjsv0P1v
Y0Wglw59Y8cZa7DGAq6O45D11GF2G2QHEMP+m741KaaW1KDroCEEHI2FioYfUJLU
IiSWj5SwHsc2v1DXAE9iyb1XWjg4OSKFOdzCAZDKGYBE28Ce/Uy2cOPh6P8f7sOU
tu+0OffF9zTxcO6wg+Cavv96bfJ/feitkRczGPVlcAhrwQyiMPC0NTO8HOYCzVGf
8f67AnYTGwoMOoJ+annhDOKimtDJvJoAPeFAckltm6dIeqWX7oS8CJ8onQZPTeN1
DI8hdCHLyiGOIYKGkmwsPg==
`protect END_PROTECTED
