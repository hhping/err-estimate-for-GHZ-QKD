`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TOmgLD2nRpbDgkS0mqnTAvClFleOqLo276mSaa5GMCmwqPIeVk4nu8TRgDAqmdpn
8QZxYT92hXkCjK2A3qx6yzCYPyidIrMqy7qrEz6aJdvL9/qcKS3nNK4tQp+AyNOV
fjpZO/dY9CAtUwJNBZmvnYUJAp53mEhVWs9QGY2dnprNaTt7ihi2zA8yjBCde4d8
HDRapDd5ikfkj/QyRhbZA1f/Rxi+/ammZYzVYv/ilUMsshRcHwKDscgvV6KeYhm/
fcEUTCB+m+uu7E3w097DwhPuwvQrdTksURXJx8NKcY6izERjyLRiiy0PzTmm6V3J
GG2g3+I3LUK2Pq25uttlQWbXAtVwMnGmZ8kt3xZuT/jAoVnOWMHeq6V2HaJniRmz
zzLv7uR/98ZwGtbQZRQVdckKsYdDTfWRi76wWSwBQarTOFs0OPZNvSLnTqOCLF5I
YP2tf5fCQrmRxyGwqllIZ0W/SZcvcKz0RUY/IBLTf50hqN0VvWQ4pT5C7nCyJbYi
/Tq5iSGnuQvPhrqEBscwaFe+skV6dDFgK5kEMw9LU3sSKGzGikr/MYD06kV/Xpcl
RdXEjo7cN+K/oNSlqAeh7yh5zevsqmwhIWHlwA5DyQaafjoAkUWfOos+4bFAu8gD
Kmx7NbXLRZ6ju0tQsojkt5qrdEeQGN9wXOgeCrH85+KsqsScsPi2jOrjURQdr0et
C9FxnF2uGRU6DHsVoKUSFPM28ZngOkeDNy9nfRzX+e8D4SCG2tyJ24RRaYWVS97w
20XZFm5+R19EZ5+RIHX6ziUBNxfO2VKo9sses6Id3tkrAJ/jD3BtH1V/XlUe3mPE
`protect END_PROTECTED
