`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WXiSr1AxrKA5ahzBtvnaiHextygsI8NZFXlefdujcvTmkCQ/nPJZMOtrkKb28LEC
FGinstTWsGzsG9Ne3c3G+J/USckNHNGWn9lYuHt9HWd5zvdIPM/x6G9efaqaR+6z
IojcMiZGhpcGUfgQ/HSyrlY2UmQxyQZMsN1hsl3VXJNcD3O8A4AiQO5LOJEr2VJ6
XwM698O8Orueh8DSHU1+ezarP7NpjO6AHIELEi3+LAzj/6pnXMIq7OHXAODgvtvs
qykBh6Pg1aIus+mfgBnF+ojlIJ2Jf1rrWId5/WP99akKy67U7Gc/Du7Y8hMJoJ2N
eHjxx3zi2tASz6HkuFBTIVm/dYUDWotgv/+R4QQbEAWmvCW1p5J4yc0Av0pzf/ub
QM4x2yr9/7RCw5NVb/nw2x9j2SaimvIhft2ttktvmInE63X+BpwoMzIIZJpxnzk7
mrjobVZ5weGGM1CMpYejA3svF7zz1HmMgWwrV1WVZuCncXnByEm/ad+OtR86SQZ6
1Pj2sgYJo8RVfBPdbFGFVRffgNezFngS8hE3K4ECBucD+IJWL2HYXi6c/fHFkIwj
4rGUoKljZpfbF8lQu/3Pzpt+LnjYkvTMcsxcGsHFamv4MAu5U1H+2dU5lXObOEr+
vG58RzB7fNj92KKZQpFOWzDEPCHVcJmUmD7aaIIHt7xAlqFT4C3dB+6OKX9IeVjp
MwUV10ov5+awRdaF6zG7Prx9zwj54ZzkJROdS+loevxU//tMwmPp6gW17MGMatnr
SVnfmVzGJfKJ7v61BzH2lFxmHs16kW4ub7S+Uu6JxSdMDiK5Hh+DDiGEjQtRSNB9
oep8+U3FJ1Tkx+1G1F21gzJJK7wNVukBGZBEI1pO7/7vAQirLVSbd/jPtDKMHgcG
IZoaJxqO204eN6c8A7o7F1qpsAj4PKSKq270X6OsrO4pQ0LqpxxTYTEibyEPd98M
ddYZfYajka5QX9Ch4cFbKJjWxxFmBLH74w7YNs7zKvvEG/MpBEbAlUhUY/UQA9XB
NM9eFGxwxDJr8PaiX3xIBNcDlyYbrlV3DroT8XlV+aIifCRbyCuSIWkLR63Au7co
UOVU7wp8168WcJomqq8KYgPcZ0XscTqPoutJ4/LbMA0gFm/X+yH5ErJfHJWThm4n
Ndaeyb6AKltq4B3X8KdMExbLucA00RazrFOeai0bSvWgcx/fgmfE5VKjykORtILU
453fkmhy55jFtFTy4jMfsYH7tMCFmD/vdkxyaeF2GJWWdcYIBt6dNOlPqUIrlrcL
ueW0XwgtcO+z+JdSPQnzZGyDxED/ziEaocHVYkm/LMsPu0aMVwwXz8biaDbm400o
MgChruAGbu1UfvsHGfLwok0Js/cEVZIC0khfdgd/PotD9Qt7+EA3XGRjL3kh7tlY
SrdXgMahBVnq393EEl2WYqJ2BJwQrTeNgsM91nPNYhscXjjdgDrRpHAZVHG4VhJn
SHJeTscvIVAI3GhuFUthQ4+NrVIFZfE0aStZu6L/Q1b0LHjWB4cgkr3FSQ6gEtmU
FyH0VvLArGedpV8j6fLCBStF0agWunGCrVy1GwZt7DIWg53CBhNGWv5z1Es1hbGZ
qPX3n/FZEsDSpU991v9T3r35xYVZZEHBieoS0IVRAhQHN2zM2EMceQvPNLxTMns5
udDzOIXibCTfIxLfQ/QE9K58mozBTIpg5KjHsrIdJT4E50JGbF9E99euwRa+6P5y
2b12cjIAezYQgVrid8hhGnPIk//PSV9fWjM7geMSesaqBj2mCeZqiRxSRBTUpIgg
Cr/99+JgJAL7C30OIs84MiFvqxckR84RwSrrAg9cO+HXFyR2iVhOYtoYS16K+6rV
FZqN9v9qhs37z/UgHs/7/9/WiFOzT1EqcaGSOlinhJP8E9JnPgObwa6kv/1J4oDx
6645uhdJVGE6nf1GQfhQAO/7rdhx8YR5hoFbdVI3RdZYcwmhNtrv2oE4OdIgB1as
K9UcIhWbZnnsqLfHV9aTTwfGAamBAo+a6MoSlp+jlASrJkZxtCC20dCOLHDm4Ez1
jAjLTjAunYRKW5zcO44ZeKzK57TV2KFWCHES+nxpwOty82mmjcfFxwYD5p1h3o65
Q/PKfJvyW5f9BGw7dn7SCvXOOMJsTomtkhdlCyY8UCg96tPIbU2II1JIYSDMx5if
u2KxuFJQrvxnU1pnZL2ZG7zCRo6lwwzUEOGfgxwxyEogn0TOETz3N7AEtyeH4xfj
WgeUwaOyRw0sr1nzJO71ExVa0zsc18Sm6IWUgHWmRWtQ/6cjpA/lzVD30aVeb6i8
t/uzv0/s3C86lFynIon8DHnLPpOJvPEkYf0IWf5srH4pp05fk6xZXPyg9oI3lRHp
q6MwjZss9bTm7vJlgiBVsTY7p3EdNQ6vMTxZuVwahuOxJcfWrwV8A0QuJueD1Ys+
cuyLVb6GTFhp14fBz1iwajciQiiUNouD4YOilxgQ55nzB50GVjzO0MrYkqEa8HZA
rI4q42kG1h9OOXaNNUFGbUpY7cTBxNDMLvZi7pgdnweCY6ht++Cc2JMp4iGGbPXZ
Inj53mSf91UfQfa3xkhalbBTGPr0KFMqKbJIQeZI6aUqo5spJlPJg2XvW4yEQwty
mbANPAgwNX6h5HQjhxlHbeZciHKPNrYQMLTSXXS21hFrq8hoIGSHdw+dqFJZpLH3
Z4o7bX65vMRFMW+EPpElKhCDiZayNWwM+40GU8v8fQlf2pwk9inqyMNQ0jmkXRtQ
dBOcPo/VVgHbLvDG793/kHmeLc6F2W46dZ/hKLeZiiEfA4aJ1xvUILgj+io1qXka
pI1IMCo1wmX6mfvu5/owQmdwLGrc7M23BrjxDQ4kTjkLyuH1tuFMiT1W40+sNHmP
DwtS7KniRP93lFGNDBAzyWszpNMzRsE0F1d4T2tAZXnLmOJGd6X5IqE+WzUTiAIM
Cf+Wl5nxK9LhcaDqcosHzjnrSsF1niyw3LGBFw96+TZkka4pa5RKSCfsO2dMRIie
RExTHumzv7fsQDB+vUnFa/dCvNkMIW1n/tRcmQznbh0Vtzz2Y36huybyJeQNuhHh
bBTFRl0StvHdP43uTTpETlnB7iGvWTcKUEpAxg7r76xt2X5nTzUjrA52ENitrf2V
uh6kTsWP6q/GqQMn0n6Yr4cwj8sjolMLbpGlqsx4KPv1l8t1So+3oxcRnLqTic83
nCIYPdtlbnOZ3n9WcpMvXyZ4OdMPipCpL4oHSV/Tu7YCe9Yt7Ws58t21da/d2dnZ
hcJyinLm/lsy2qe34X5Sih9EP3oBj5U8XENgLAkSNn4DtFJO9HuSUZbXOZ3B2c+A
CpschqxCSrfgQfVOLp0XzFppltxqlOMxPdFjYt7TcSHvzQLIKtew/Rz46g6d6UH6
3RbtqTjJXqygwWZ6uRBV3hI/51QM5AdZgpNSiU6r41Q5+RRLveawK8SCrmmBlVFm
CCAZB+lQSatcGRQGa1avvb1oG9mkGq+ctWoJj3mLPmQzUhSM3hcDiSXwVMi8FGx9
M1kH+xIZxMlkU4T095xEBk63XHWJxKwr5Hec3OfiKYmQCG5CYkcbstfr2cm1rxrD
0mzsMChOIUKF3FJhmN0aQDV7pfdTY+khurtDbQxlEU6MzCn5TGwaTdlmhdBGcKQ4
ZlRgDSnKvHACwfoDsKQFxDdFTksSkT9dw68DjbzxDXrC1FUgt53z2RrfR1qjS3wA
5v09yk0tyxMViDVt2AZG5DaNWJ0AhRdhWLRauarE9dP2ihJ8rBVxlgtPD6p8bpRc
fWKTWcDqZnQGzyc4UNN3bIdDVDQJMBZz1DFtV+Kz1yKWTiie2hGDW6q1kUHcbmAJ
uE/DsrGNNqE8iz23U8t2suo7jEzm6vLRnGr/urGhu1U1eAyKnrUyEWl78T+7jM/F
TlTWmpiiZajkdS1SIbhYb7VPgNdpTHZQgvAXZWSD8rAfwUeOynwsTyBHX+8aSQSr
zkA5lj+76i2ss4xxVqDsyNwucyYsRq0vkTUH6pkrNtDgdfs3pySRDOx9OVgwUtqO
RZaCAmV4Ev5rPdxtjzapV4D46ehY3TZ71fEBZLzgOxAAgE5NhDptlYg4GvL03Rs+
ACj3p41SdhkvSmPQr6SPR3cStUlm2cFwbW//iWcAMT9safUur81TYFu5U8Z19sP6
NwObUEY4j4precR4fmRvOwhcNmPn6gsymgRsZcp6LnLOmpBimoUjBFbvTdcD0Em1
joTuOlL6hENKtTGEWVdcxhCBXxg8QV1f4rw1SlxfzCkoRYVW/nlIUWydkwI9l1YO
w+I5fkBi3Qh3I3X3ypWsTHE/Zs5+wi5WMGWRB+nIW/P/nAF+mgVJfG1SyUQPMcuZ
vvZLHtdVD2al9ynsEuJgPq1lJSrsyPq/IDSLy5O1WxEP3+ry30mexxxVnNAzMrrI
LEreswRA8E8aSFxzZV4ccTvt6cEI2Q2K4I6SLQPnPFQUIeh2IG0IsOZtHsQi8Hk3
4ovvHqJY2b1qlYsRk0jAe/ZI1Mc1wpAiyUMNNth9sZfKXQaY/T2bnDXC1Lg9/mzJ
WMC0mjbyPG9m139wpLfPW5EHyZH0lY0UumSJefAGz/a1dmiOKaonDRWTzdtu1x7g
4dUbsnpQIBni68vPUjhrZwVFyZ1jKfmo9xMzyioqHHJDhwqc6Mj/cm7QaCtbbQA4
mItQUbzuzbess+FTHwbq/2EwYiGqfl9vvyUDORPqc8X6siB/+QxyR8KlnieDXcig
CEjH6S4m0V9fJETekz6rXTbjTXCzz5/Ermy1fWFJzz/S6/xeQWXbiXdG4DedjGcI
Xh2Z9or1iqgZnNK4H8jKEltuQPzXUjk8sdijPfcSdr3xI9wMOO4NtdKdwiyd5rpS
3zstd6PsuJqXdeuJTyYufOHcYqzfys8kxr2eU+YuUhklqwE8Mc4CpHmOX2KcYGPR
cR7nVTXGn/wnshh27v0gBhz7IVrs9SDSVPDW1afLLRntPPObWLBttngwPOUkVpNK
dL3ZeOPanar49dHUwoeLAej1+s5Bg50JUpsMTNAaq85BjT05GsmJnxE419AfsQ74
MZBnAfULxJ//x6FkycxAeaDK2AKlaICs5L+aMG1J+GDZ0MjwBKxm0Awu4ovdU5+r
nzVajTPyzWCaJuUC6G32IOJGn6Jiuhl20Q5+GtF33/oyMInEZRwVEOMXVpAN/MNT
xej3X3uRy0qnBJCKbkAXDHl6NOqt2x1p36sOFrnpZWu4HPccOoGPa01qJU7SnXE1
leaDdxGBeNj2QYNDIBgpe/yJjpMORKNQrBWEmaMIzANldi9oRxHDky+yQYYa+2EJ
y+s6qaR0MVxrTGajJs5MSMAb8b+8J4H5ev/q9EvPQk/LfxHomErjKEyUL0bwNzhJ
2DmaQ8WOXli8fMrNhInXjYw0qj3vVWlJvF1FDf/79YFnZD5DeckSziJxf1nGIZB5
MyM7s80gDNcbdvuUWiwS5WMp3YiD6pvPLPZ95Loiphy8V1fHun4oBu+JHcQcG25N
lzU2yvf+3mQvS6BhJqhUC22MdYF/gqXUaYuFii61NVqJhod2DL9XKfnh0BHAJSa7
+dqkWXD3fjD1SdqZI1mNx3p6x3t5qka3OZpQPIQEnE2SZ3hs5IkfKldApwN4WE3T
7Z0RgXcVSuLz6jivD69StqmqHps+36Os4VqV6TwfrwZfueMOV8CamyS3tDwxfGio
AS/xuTCQDxDrBQYvSlpNjmo8FZ1MmzIrypdLL5WCKA/4ebOkqLSu9W23z4H4mXnT
0s7YSsS4I2rSSlUlBfWCk3UtfxjWR+Ml6bYNIMS2AqWw+WJfLClv5fgkSPHIOoOt
SQgZcbfTYA/OIJ61smV0A+YEfMb5n1xfEjbryu3hT39qlrORtV55Cxp+Y4dyVeDg
hCJ9rQWFL5vIh0BRa6vXX/znQeUPVZNM3vUEsUWmdXi9DKOiY081/2oJj7nl0fdw
uplKos6ZEe/kTz80rbtZiXrqdcOS1zzXWZe/Kv4wqgfUWAHyhWzEgoEXO7pHxtoC
xumCEMXwR3I3OANPMYIuiFtEivzQQ1YQAB2mlF5QqhDs9dufds7MNbygWzKPH4Gn
ISVUjBKKDR3RuyszXntnhQlmQyptVDdEgYFRFqb6Vc1/ezsnO+Sgmta0gPhQ5OPr
P7jilRRuefzto7fh9hxNE6qRxHN7M0OZQZLmu3+01WMhhjHh0PiU6quNLvdypGuk
Iyz/GJX/Mx43uxaEicaQtpZTf/SnGaa6sPnfeu56KE5d7hUcPeVK0rFp2i3Y1jst
PneaXhEEBaaQ81udYhOL3tvABGWstaJsQEfzIXKJeK9MkQ9c/9FowaW2Jo5o9kxp
hEV7Wo31EELc3H+VQnNRlBioeJ2+wA7iPj667KCoUTWobBcVHqNpqYjcUnkj+RuN
7f8RgoAZM7UM+FzvztJY6d30iMsWW3AbswbFlkgVM6Sb+iuF5gtgRN427Lf39+rG
3pJLqU6iHswMc4Rk9vtXyjd3CuGakQ+V/bqVN6a2Sq9M0WS3Scc923JhT4/hWAR4
q9sz8RrQpU4JPAYQXGI5s4aLeD/+MXTaBwtG5UtWi+s2gHSqTG1Ib13HfJFO97zJ
lypfCJAxGDCrLj6dEJEGLXdIVwU1P36wyjdqvnv9NEE4m8+rD096ZnMGK8F4WBWz
Vfra/TwF3X7v5HG3FE3zdU48p0NaFKzhGlC6zfEvIVFkZHXcraDmw6iPIF8MJBwY
vidHEOnRsm49n2n0Xruh5PXcadex9gYPxX8hTavlBGwq+ViixSMEEaclataGR4Pu
kvgXsyiR3k6HKHIT7Og7PgRc2tvcWPRVGH7jFZXHAOwLvGBsUn+6AFRpbQTV+jbC
Wi0FmrhfcCcltSkcd2sVPbVvQu52AVVFTvSNe+bKsaijmWTOh6L6yv1Oqq1OPf6w
LUpZlenpUY42bPr1myXeCCKhfhaNNJbHoQiVA8X27z3rC8CV51+M5ptufWtgw4gV
fjVg2oaLFnlWRAwKMhLnhkiEFdhayLFUHOepba4DWj7juIy59kU6Ow8jL+//A3yt
Zps2Cedug3aXgxNBj2uReuZcIim6Na2LfJWOGGvoBC19w/6Vl8BYxVsyGZkqpN0e
g6vjf6Vy6QLVfFeuSKMYq/qOsUL6Kmbx4dtUSOyh9j4VDqqlWEvYUktD4O1Vcq5M
sXe28qnmWejsNRN4uxMtqKnGGPuvrMnAvukL+qEgMLWERbx/oDJa5uLr5Bm2j/ID
l8qDUNhIdLD2OLqaQ/5jVys2G+QG88Btzrn1lXYRNTusavSKxr213Jg9+xS4D+vN
AryZxy/o7FWql80Uf+AEwMhOMzxDsnBPOw9GtvlfK9iR/DO+lIlaNZU1FRpBl3Xm
ckRldTVxJRsNrAXzyfQNNLQoWBb3HcGwTfqkt2LZO7QpwVeWfezMQko6zHg80GuI
vngde3ER+6TX/lSWzNgYFJZSDjXijY5nt90Ma6msDTEPY0rwtd3hCuxJkcvIfKjN
YOtyu18CH4NLbPNbG1eyYl4ekj1H+74RBTxVZqaEiV1tTXw+UtVjdGL0HWs61Jm5
/XaiD3p8qx0fhki9BUnHehNmDpEImZZtZ8IbGwPoTuwc0L0gVhwHIx2G6F2+W4db
v7AvxUZDybcAO65Eocv93IDQ6SKZB0lsm/S9Sml5pm3+OUlIR4m+OivsnS5avyeI
Cy9rLjqR9v4taCN7EW+m5530eQPn0QO6BNtw3YGjd8QZ3JetvR8Jz6weNzERYnxy
KHMEL1GaS3dJEU6UJ6o6i0HWRLHz1udITO0Q6VGHsBwqFJa39nQ/wZ7+8DzxWeQJ
wIRzXNOuXxhzTHE3kpJhh5FouplmpCngNhkVpqPeu4O8ohdplkVW6whbYJWJPLHH
cG9N+ImbEkrXWu4OGQoFh/Ld5WqFmXEwKW0HORmRA7l5QOer0gGBK20Q3Z8j5AXE
OA9CE8elAxY8gxhbzzUrMDAiyZSmtSvRC7TT4jfeZo5cl5Ew5gTfmjmux3Tl8g8Y
v62+NBEMIxM+4jIHZB88k4KxVkiy3PN9Jo6FHX2IdEA3hSmrOGMErmfDZi1ZsffP
Ube0ugMNJ0zvy75uohxQ3siox2sdNaryOgOcnutAq2vhtQzXaIafdfpIlGsD32J0
WC6gejrQcW26BNmHjoYIwGHut29CurG9MFaOeMDuvb+Cigb6cjqJ7hMyVMLWRK0h
7Aj/eo1eCnfEeyNa+qxfCZWhQ6ZeC0qKxEgYz67N5XlXJwX4SEyg5WzuqajCl2JN
c9T7CFx/+tidK1K2JeNty8+jB6sZhW4wI/yP4nzXGYvg/EFXh/77kLHyggiXwTWx
huBKcgfWCLRuitz0TfncyM0A0wvQ5SMtZrJHQJI2F0GD3adt5SM+GUIIC7bxKsS3
Dj2K6aG4cjrd1WYpvrt8zX3iKDu1e3pr+G52vp1Ui5IZXvt6s/I0Z9LUyqDjNlB5
VZ1uR4Jf/rXcuvYmsIfMOnSe9IlppgxlUBoRlwzZCsSCQGYdVgpurox38oKBJCa3
Zy+rAFfPYXTg25vuNfZZmoJMqyKKLArtv2Td2q2azTnt2MH7f5Zevp/S0OdGuQZo
X6T4OCRVGpdNtJdsbO3zWippmGqt2sk+d5wTfenGjaav6pzYQYhi8MyOaoWfP7gh
XpSNlzwDe1qieeTm33n01QdWDyXSzAUSPSLM8HA2cjoeNdujns5KpPoWDiFgS3Hb
LlPODVsXkswx6AfddUvqqHs0sA6o6Ilzf55iNom3H0mn57Mg+5iedwvGCdhAzF96
eTj96h9RpNUb9ExisdthfjUUsUNWiRTwKtbLLSksER/TvrSqeS4SU1pzfD5Cb8W3
8fvuQQZTnOlClb9McDZyVbYZ3szvG4sL6LCbCsRoZexOfLNohzvHD8Ax5F+BvFOD
A+qhG/YLr1Rq3zc5eQt3fwpqkrLdz75qjxsqTQM1lWH+korvW8exTkO5Rh1gkP7p
MviMJ0QLEGDr8mv+iCJFrZQ/ktnXl95h8outa1I1AYbx16FcTaOq5tExGKBEoz9+
Zw+8DXfAhSvQWSTEi9zVCd8L4YyqJbJnQ4EGDXr8rzv8rHjXg7kxryP9N2c8FClf
04yUvyBxaiNUAACxfV6K69r2lR3eMhB1xiFD6MtTWUlw1dTewoluW8f5uxxs5dBO
qbTSNmABr7O8XeF8exrR5xpml4/sRChK3+MPoxiuJAwUqOFJv7WihE+h1l3mnUwa
cQgNMS52DTBFDkGtXzVzpAWhep8A5ZiYvUZUXjyKEd1g457BaCAkfwx9R7/jJs8p
aikV54CIyYPKnRa+FkoTbl3t7AVOlgTWJdjg2W3qrHrwPnYeq0/FJ1R6fOvhYnFG
IkfAyQG52ZEzdfYPrcIFxmUwEEqUAbQdaLEqP3v0Hgm9QUjrNupHHrsJATgdQaZd
PVveUJiIebohrmz5LumuobOLtcyMByiaphNuuyy0nrnP7FjeD0oe2tio/uhAUubi
CD3g1JYYBkED+RHY3tguzgnIBMXACoWJG1n7SGF208gJi86oRUzxxKA7oHJMOqsZ
ltYn6T1j9cU4wkpbu+HO1sWOQvLciJEOXtZE0fN/lMA7V/gl+8y4X6NK2Quraz0D
o682DPKJ1ookAarWC+c8YQ+LNvIPZkzluHGZVvtdtmrHgAvT0VVFUTWyjKabtjiQ
H7v8hP7R5TSm3DmkWqtzwLFX7NNvTR4UHgYWcnmxxivPUTCVL0vpdQ+Uq5L5WbDF
TWxTbSO3q/rFxOmNSUTIcQ8YauacsynIySHmouAL9OnFtsyQqqQa1yG8ADsquzB4
Wmke8Nk4N1k86neVUB/C8XZLxBDs/qZ4BMfnu54+oTRcW4D76f7lgxSfDtZqW4xP
azxYpilmOTojAolCd7PKXWFSzy6Kus258vf1xTFxCsegsaW29CwC7nPwscgsgNSt
vd5nOS9iU2ffG0uDux/nGprKwTlHaNR6Imu8lGbIvjoHJfEStaJPoa7612SMeEje
8kFe4xjH4hQ9H6x6BUiiEbx/rhMNAZ7NvQ4Pa3hX0ipAQXVpH7msv63yoiclO7eB
FfC4aeRMX+8N1zdkRxCCpL62vGS2UzaAmfBIVwWJkaAek2a425wMNyCaFe8YxhUv
gkbMOV+AY9XRKRR4vyWOUTbHnK4+5DFFTSjdfvAkGDmDd7BZZTu/Ix0SeobUFcbz
qUAm2QgdFbqOGLZNJ+5DN9W2clo8x45DUe/BCV33lkeS44r6XrEGwXoUAxaSOd6F
a8EKVLL8+hv/yD7OMsivVBML4mB3uDgGQ8LdM0QrDI6wg2vNqKEu8KFovsj4vJ60
CQ+nlS7GrHgIdmL0d1oxa4qo+k5UAg4WNtO/BhznXs/Cp9gnG9j6LqMyPGrJ3BAd
7tAXknCrqHkVZ8zxMxP3c6ua7Puq849p7e45kDg7Q9CCmLdQ1FsyghSMKAn7Nz6y
3jKbji/k7PtW9bkQDwLDcIWOievNxTBzeVbO2rxg+STslfbCpcxhxr4ItOChwGf2
oBkYLsqOvHloK+O2bEklfRKBPBdbWClVbmCDgwo7898yWbcrhMzJFGT9gbUthvpH
xYzwoCLNUO3nigCaAb3sXVaymbhGzYGiygV3HrD8yU5I+/Hw4RQLBNz802SkskEk
jhBmTlQBOYIy42F29p71sgpb5jj4lmIFjB2syMjhoh1XICaIfXceNKgZexrbm33D
GrWpCXY22mCkXWVqGa0sH+UrLyoxmnvescAWwQ/xYMxWmDbd6bQuYlKA1xAQU8ns
yW6ByoRxcMvuSgpw5pEulJVvSpf6DvOjM50XtfpHusxRY4Hswpu0kDb+c1/HK7jJ
OIlAPpyzA3OA2OhSV5b0SBlGvdtdWCh2rNhD+4AFpvboM3YIJWHGpluM0wfIaUbI
vIM6VCX9Zwy1UflqkYiNryN6oZxrr3N8DakzmJwdnOfl8W34ig5Kda1lh3WwQetH
dhxnIv5zS3oeZqxO+z0tnbyUZcnnX+TqGcjZ+VGLrmPK68NTocXyfzuJ9mpvP3fy
GKiJPqFhXTDUnpfbpm/it/I+qFPrDMi6MQkkmtd0+DkCrlvj2YCH85xCi8PCwE8O
WO/ipWFs17yqyQjclYKrFGhyI7JllbZnmaFvwLOZAVSr963NxtmuDuNFl9qfIcXG
Qu9ze09KWlRj/306CUXTKcHzy9rC2wOgF1TXId0BFmyT4Nnv0GAyCrPg0ckhMe2r
6ZiUMgMPFltoEV+WEJsGVFRBU8IJHU0duekN5QISwpZput4nazlPBtfRoRusN/hk
LWNjTz9pshJLpcwQMIMxleWGivz+wZ3CQ2ex3ozW8JdX5KTP2Gin00+v/dPHnm1T
KPidHYruoZjJiYfJWP+2JGiCLgga75Eh42A1f+V2TViIdZkp5qE111w0hp0cqfDv
oOxKiUBOC7G9AYOd5hq1rLbWwWAW5Ip0gmzgreFtGvoN5IWMUwYmvEhKqNarV7YU
g0tQyNjgP9L4FLBm4YknI2i95kfEvYc32VuKjJXFEYeWCWG3UxySufh2GZx7SCGY
xv5u3Wp5j/vcf9cf4BGmh+95nAVHrtSD+hvl8B7yKI1GHL/KyCAYUWwE0zYwLEs1
YTMRYdGxm+sQGl+YqrgIw2qJI20ZnqKFGCUo5d23O8L5NXESgUufm21PVyBMXIlT
4i51ugzJf8j5CHz37nJMuF1HAYpT+F7zWaZS9X7UEKHD32GwfnlSJabH+ERk/d/3
xti8WUzHTsy9IyLjTy00ZzOxIx2Zta8s2Y/c43v2gYxjl32ePvHpbvWAa2ebFEDA
p2UzTsw5ByGS3/6guOE4HMCrg/YxkE1ZcOc43vrLviMrVx2tiImrA/jj51uq8LLO
b4e+f8nvTfr2ToBfPEKCm97AH3sSMawsp6E75BJ1aKdBx21T+jimH6PXdDdQJzMd
09L7fsx5XcSdYf8kqxK1YhDUG4KPNk34c2uVpK5YUScUn/VKtI+rQoKM4onyEXYr
86/akDUz/dq9RCEyL26BJwcTGn/b+Wl/DrlLWfyzwzS48HQbsHs3awuwTBiK4RYw
B00j1I0R4jHhQaYwAXyR8yKsETNTTYCuqC+W16oJo8SaLHv/m42DK6morYUhRjBT
/F0oSA8e21qBJ5pmuV3MsTSuWHGoZPXP7TTk02bjHuVEoLboA8QIkkfxa5mrIZsK
fUaxCv+5/+vqq8fNdHMuM9Jz1gtkcjDowX5wBIhLPljpun7ddbNi68G3HvvoJOnY
iSmkQzaaXf6ZwHEVr4mb8ysyVZA9IhxUecsel/RUVoZ9uyP9H6RB9KysfOei39SE
DiZvB6tlehy2D52lA1bNEmhrQbeanu1dTLzHhC/3PjwSrAKEKOdxeti+3/SjXMDh
9IkSAScFA1w2lXeQiN32zyRNAMK2PE9MAFAaGmMGNOroqkxsRd6SyOB57B8z+KX3
fIDHyuN5E8eySiueW2Gbs1xgrRXSp94BfYZff5DUBa10g17uvWfg849ckmwUXuP3
AyrkmHymXCVbovvv22qXLY8UoEcGY7Th6SGyY/jfpza/dKQgDEJhJ0cgmU9GVMge
stydt0PZJyk2BzJebDtYkGX8WUClXeLSfo21lNTWACvDyxzmHfVThz7p934LmB7M
MPrZUspWtvaYRMASj+mZz6vsJFFoByCI3DXUtqkICpk2kUfW0uY8PmdtNc0JL1L+
gvREcmv5gJuICB6gUQKGQOmwtHhf78kPd5l1XyxME2g6/kcmnhtk3QbikpCevJgJ
yXJ0Oj6pw3X3uMALB2ihAhicACwJdHbib9eakLAPLDVwsiBYlcbLjALBfd4Lloxm
CK0USqUiM4MFsE4y4PGQzSFI/Cv6wLSr9e2NjJ88wivoyuI+6TDk/LYgPT51AY4G
RhEQWXPw7EOAUiCiLABMIZt/d+EmnrT3ElIfu6SVqMgz7gU4SaRtecTPMDqhWZV8
r//ZAVJDev4RMOUrTRHdiGF7up0eTKXcEOUykUeOJGgqpySakVr5NiiBNsRb32WX
wsOCJ93vnI2Fa4r44nT6OvZw1wZNNeHO442SY5goFym1pLUti6zX62ei+wIQDfsD
+AU0kLwDb6+b9G4tCn96oJYoOEF8Q6lkoiysKbKr5+LyWSL3edcZKhV0lbzPf+KJ
WbpUw+Vgjw+U+lOhXfctHa0wqDU7AphJk0TwFcPiJA5K2E+7WzsIrMcTxDUFPzGR
m78mK8m+ucgkzReTY4D+ZDtkNnZXngi9r4GV+EHwGE0Ij0WxT7qoX+btNQZFX1aD
4JKNgNblisjeLItYWYo/4yMP4e3yyhMABvrpCnXwqwsza+ibgevr4OG34kg+Wwx7
O5YvwS4hlPKwKBHHnKlqzvXNrYLLLaPV7epBNgM/57e629f6ggSYps8dVg1P62vU
l+pxdBApIEmtuC0JkHVVjRyql4pN6xHhX6p1WwlfHO7rOQhpynF+Y8/CFtgmCzhc
/pXHlVLpnBg15vuUrb9epG4q/A+anv6/YctuBP8h8MteVUxlS5+jV6uRRgzm7sGe
Lg9/liBOhGYavxGmEnC3nFzdY2Jb9midicdVepcX0FWQjqfZ24GOeQjp5xZFmvnN
NHxVuM7eTlBPdMJEj6kC+ZW+yHpcYIfBKNz7WfczNktgzdCChAU/hI1wYQM1FWO+
5XpAB8z7hlLi3gzItfJyTz8RtNsxQ4jYonkunkYMUsCzQRiN+6sPWgxPanY9/LKa
l+cDpYeKZOV9wgxy7IhYGD5j37TrCCFu15aluFkfqUu9+AKgSEBNF5EV0ZuI4hGC
769KWUPxGBLn7z1k9KKA9/ZyBvbaSjbZB/4gDRSSTHalq+26M9++v0LAlypMvNJ9
kaB/pde1veeOBoM+WP0zawfzzYWdd/KiIGyYckOB8HIzFVR38iUUMkSlFDifyZOv
pNkCpKdHKSXBN4Rk5aoUfORK/WWFmre/093J656vm+sAR0u9NsE4gibJ+7t24cUo
t64v/kvzQAw0eKaAdhLa5g5eqJ7xlvq+d765vkNAgmqMtxsUgk24qCWTR0R4Ev1d
IVrc42H06XV5HcI5HLbCIF0IlFJkkTY8xZBrmsRF7G/FraVyTv0Ykh5nXYbAHFOL
uAk3mEjHxlNaRdXsd7fkPIU4fVBvNAtl8yuPf7Qtx5WuDwovHatqH9vRpHR66+Ju
5JiSgEQmVfLbrM0H+aRUMts2MVLtGvo9JLR6fvbHSxZekQhv80Ute7zdl5HR7tXM
XR17E/W83iCy0fbxgSA3lRysIR0uNquYZbgHov18B6ma0RbGbgU+v1/W+UYeL4Ht
HoeXLfa/xTcyFTcTVNc5rzAmWVyMmvkAR828MNUCZ5imFqZ7exP5PZYI1YO5HNcp
UmTSP8L3nuY73Y083ElnLRDigzeRVI37Covx2rTbvidukzleLYcmBPWId/W2FOGq
gWLxinLvJ5F887WVihja950i/5qTmHhutG5D52TCQ72xjD0lE0CJOf62kL0PBBMt
dKRRbFU2GJH8DZtnzNUUZZ7ZUs4wJ4reYgMBMkO4pfbJP+D80mFqy+QwHXA+qy2l
fbfkWNlOVGz5xmg6Ls5S/gWhktbtsp5kfdEQZyB1r5TW9nwIYUT1JgGdsf7lnpAM
et5HflMsNVeoKJWIJ/uZY5Q32VRuYvh8x4iGodLBp4o6sk7T6JBnSnWdUKLFD2Z2
fPl+kic0V95ZeEiRq08SNi5xUKu/YcsIrmvRPGmSRV7PFbfBHpBNMeF8l+4eJmXv
/9nnWKYQd7qMNWuuCEgxMyfE7mm42uYtNWu4SeZahDEzF2fE7dCb5x21G0F/lF7J
dohdcB91FpocQ9YBJwd7BVjaOLUQXF++BFhDHK9IzEx+bgRYAKwjQnI3vxdgHt5/
vnSD+8Ge7GYNnANCuEw4TCqAAyEddMh3YDas7sSFgB/EGkg2bedDwbUjD9J0y+Ey
GqlGokZqKtlHELIyD3SPR5nY5Oa4YJk1P7t+6rfs4y0ZjcGnXAFE6WS6Yz0z2tgG
FdyK7RY6bnQJHEaPCd6jwCmsGgie6HxrbDghgenhZr8PPRreVneNKyLE9xRL3BSv
23NMx95p4h7vYCcyII7TP5V2leDpqDrtGHpyl635clCTWmgVLObIBp3lcGmjqBdM
a7FiSNiA2y/CubRiIaXWXNh4cQRgNIjjz8nTD/IeQkh1xTSvwGdrIn/vQKQeddjN
eX7aru+28BJEn4ayQ6bnMH6JauqVnGGc2BjiBxWuq3hB08UKQX2UpOpjyVtZUabE
WGpOsdZjAQLdWHobeG/FydYDVH6R4gawIxErhJIzGzdNA7xcd1UfrI3fHcSySL70
Mc1xiJpZPTfWstXYoS5nM+jLu9WbrlEWalgS5hVANIwJNgIHkutob6E0lrVojcoK
xSwIWOYjNJX4/85eyYFLHPz7PNsShjiKOR71HOIHkxS4DBY7g8Kvvbb3TuRCWqcb
LELPVf/j/c4DfEH+sXA3bZrBqdcfiT2KFiA6M8z6sapPCrNSEvjpY3iCep/OIQOH
IfzrtCXu1+7743ggm+RW08PKsCTfjcAELKWaSgmvvisO+2UZH/tlnRhuasNISjhP
XZ/8RypxkwCx6DLDwwUHETKAHWdTWoZ/Agho74l2tbpYQH+1X3O45S6qp8YYllwo
t/56u6LwsmcCEjTtRB8Ui0S7TYU8ccikdD1p50fxBziKTLbPy08Uj1Dms4zije0c
oO/Qvf8EdzJh291S+/Hevpamhq01J2D9gCTqMpmKTCuAeEM1qSRfpX8Zot6ZPGzZ
MliRORHrAFDFORHORvoBbpLVP0bTDYfLCNpM5rQrRyWrcRCF9IpWGORL8kBZJaqY
ObLUrEFuzAqrz2NiuvNryqU26YbaTmyoOzL6D/TS59RUxqSBzwA292KhLKFycsYd
+socDzU3nC3n/KIrEvAlj6vBo9RyH+5Io9VUPiJmd5dRW0Bn2o7t3YD4Gk5lwNjT
2p75PUvVI1qbxbJ1iw2ccSoohctyNZNZk1VZH8+SO0gFIqrxHOV2jysQWksFklhf
FAbgXYuwg9pf82SOFuehuETKwDAkTUo8N6wAEJ6vAsej6qwQo7qskS0NlrATUdJt
KE9voM7wvStnZXiwSKMqeMs0op2RADnu734Q9rzvVb39FcUf9yCnIpckAjG/iCm0
ZBJThZ4PrztG6DNKxShVqTD63cPucK7kVuBeXa3yDdLgkFuu1xchLwH9sFaHgQDE
5BO/yXLcELBRfFtMrdBouDstYh1U8d1eVPL2ch4TUUFNBrQDhG91m+Den/UOkqyd
hqB2la8UzzOELx46j+CRYW63UKNio3rxu9ywsxPY7YfVW3Ehr8zaL9MO6pdnxCF3
JBa4T6A6czjLJ+Npeky6xkYfYeKP5E9oLhBNnS0/n24FDxAfuyEIt+dox/aGivwR
iAt/Anfq6bfPRRGvzJARjhj0v9N1Mf9rJWJZBNQ22dCibYrJOrpuCkIqxk/rCFr2
Mp22fsWNGqvmJWP07hOcLmLzV1cQWtYKbBGD3p9B/NBDuQRcWWmBTz2BHdGBA84m
+MdcUBwBvI+tyxbgVW24olWqyVlOxSa33aWYBnMgVbVog5wdqcN2q9Ea2ibtLtCm
I2IemaGuSMe9Q05Rs6yzqYvvTcgdHHcfuGanDMP7B8fZdMRhJBSNOeZs17d2u/Z6
yiEjel8/ag7/AWcf3fcpKJFq1t+NCxZI9OQ23565/xb1daST0Wy0cgtllANItwqx
7GqsnyBzi5qMXyFEPvbbsmBBNgRXTrDQIQOmvNNdecCz+38oGVnWovCyvRKgJnd6
upl2A0P6R0YjBDMh+l+TzdqN1EBTDuMxxLbyQ7obLc8HYViMYQQiiGta/8CszJ7i
Obby7capGjLdPnNQJ01fRMeIxwrL8sAu87dW5A/mC00mD1XZoGDwijO16mdTurAM
I0iZI6JGRF0MvzA3nfZrm8NnPxoWgd2kd6Z6jk31X0oMBy+kkoRxBzvxwZFIBeZz
rQ93Qyuc/yRby68DkXZMZvEwAefC651Aw8QdtUBPiSedpbCdH9UZiyXXxnRSfF5g
12RH4MDJGHa265gG6gpoG4UNFg1t43jes9qwO3wYq8yEDjCczAQMDw1u9VXdcBFN
/5e6qolGXX1riPcPcXDjPrYU4LYh4fUSKwUEE1+7ZaMDTuoTrmTw0h1TsoWTBT3S
RIR03Xiii2ildxKlI0tIckOmGXI4UG9QSn50JBy0XMxjPofiA1Q220B053jjvvfT
lgarL8LJant6rj1/KjW+Zyrs4W9U+vacZSZOPzSp23mn/K5SUUBOzLQwslzCzegZ
gcAchWY8Fy+iNQkkILpq2uZP26oGfqGP4rEXyqIB937X7IQ6r7xC556AeJW1GVgt
Pd/dAOEVjyTRqK7NccIEcRYTy+ir5wF3BYsrybTUEDH2NJ3UnhlIPmvCXa61LH2q
5lhqlDdL+MoIJopsF2NcCSpxy6wm6ZwFMVkQ8yFGw9gwDx39EAkgHTI1YQ75aAst
cIfXmM/wPwEI28MexuH0mdi4ZtG9qHKf0CyYcZOGT/SEqHc38J/NjdQSKl3Nq9I6
U1pLxKRydPIi6V6WcWBC9qbNh4wma1gyYAwMCCnipdUgutwNZT5zmoFneH6PRHiv
NHxA2KFItvQ46HCEpmAy4zFQZ3TJKAlgkzKWnDrwpPqdO3LwAnRwPOPDaVc2wHWK
2gZhX6p1EQCqpkm7X1Vub3WbZx1vK6r3WkXfBp7ykHsa+42pH+d1A3BDQtNG0Rkq
nEX6oagVpv3ThHs2gmFWYxK1Zv3Ll7/+igKD3c8C4rnD3rJ4/VE9BncXgab8ssGe
Axju/dR5yZONWWsjunk+khKIzvQN98ARCCeyPGEbavFrVUtTeVbofkWUdrdSRtR4
Z+e5H1hTYIESETldibT+gxBp+FpT09jwy6UByPvoIRWaCru+K963eVomjL5TxN0P
yBjDluNpkajd3DV8MWrVf3KTE8Al1aLcQ01Eeqzkimu9DXOLrthYTfCe4j3GZTWl
Wx7nYAa77me3UvayJUQEJF7FU+8KK59lybTz+woK2c2ztJtrIdGGZfeLq+we+0sb
VEagQ2lIt6m6ZUuwEFYFgsMQmP7ytDCA+PMnwzs3Q8jkcyHA8jHflcyKTLWRPE4G
B3iRd+J9ALrEyceeq0iubbVuN9IZdT+bvqDqLbZR6H97bcSYFWEU5JsLhYZErmsd
txb+Lz6uKmltQb+n0m5Fqvdm8BhzEjvVGpKCsv98asnfxYmIumKOaJHeKcNut3Fj
budoJ/XcdeQbz5yr4QdY6QZ9BY+0ssbsDKVgM0J+mo13RSN0B3e8ypNbV/Zqn2gJ
ODfLrVWmbxlldjHNYZJvwAHZFKngaAHhGsgtkSW4g6rRytAfcu7ZHzlB8mWsW3Ap
jut/wDxTOocp7jQO+WA0baWb3gn7PgxaQ+79ws47zkGDSMI4yrBl983AKVF97iI/
4uanjuRNEYCCtMAf62IUu/MqDUC9DuwA3LFns9BKCyRCguY6nROG7kEBpd3d+wnf
HTBeU8VS2Nz9YdghCErTuSjfcmnFdFTayBI+j/qzjIykoO0ypwKuzBmqAJaMKuPB
pO1sHKwec6W98CJJibCqWwhNClaAOfqXY/Uxtf9vLpfpc/HIyUPd5v09cZsY/X//
eE+PUA/DUgcgtRi0AUECxb8zqnBxUwt60FWATj6zXaSiXnCgfhkm14ZOKpDklJqX
hjR+/0FwAqxoLYlWia0DyF494edtMztvdYtdJjNek0TtYSaRmzPzzydi2rN3dELu
SZtUow9JGiOwXc42DSkylTVk9Wl9BviOpo3gpqpU305Hld7OeVEMkE5vabPdMZ9E
WZVU+FUatcic7xQuTxtjbcVAiZCCA8VTJl/oIWPKDw89wLul/fBQjeWqrxvgCL9F
PBE6IFlv/4J0vvORiPcvR5esWDx7rhEPLrAvGhrSjDacKUi523dqh+fAUjmLQfKM
WOVtoXGlRDIo4ksIEclf1mG4feHo973sCSOYwKi1GwBfEqlvE1dggha4+6jJoXCg
TdNdfNbpM1wmP1H1QbX8JtHqQX6rAyJvTqNlkJsG/yRYFOFA7YnqnSNsjaG6r0vY
rtTPPuyAkwUFKwhqFaZnPNj65zI2L4LwbgMMFitW56OpnxYv+YxllodDLJuhm0yu
bRhIqxZMK9mTER/sOwjIWE22/JXUPqlWoKM1g/TjXv3XQ8FxcOnSjRHaQyyHwJht
zYp6QEcplS620H4PMkfT2ru1L3kbMv1tc20VdJraoZISVj2YZa79oHXYA/qVHhJT
i7vGxv8X5PPHdE2/9Ie0C61UvKWuAJaorIJCbeMF2GHx9RSQKSobt+bw4644/XeN
uABEYRUS58XQpq8WT5fsHoQtfGsl+4bsY7g8pq6XxtQbXtvszyBTnhaZEixCdXzX
ZkpdN4e95t7yXV5fv6Wtdu0i08gPVo1uLrJzVvFRsiRSq8qOxFoUFZKbwxfB3/iw
Np9rJajsndu0l3hviGUbVEx31dWSHZ1HZA8U3e4EnpPtfLOhJ7JCyk9NJzcn7/R+
E5IASl8XtrKGgcujd17dsQ2A5r9xJdbGUoXDlp5DkGyilwptdtQOKxH8YEh9ZdmB
bePLm2rvEKSwr39yJEI17+SPKat7V3Jf6HMdo3jNWQZ3UyOEw2PPZerizxPFTs36
EnUxLTROMR6L+F0qVwdWXTm4q0JBtI+QnSXRCyRKsQQuFK+g5IK4jfIX2cfJs8vg
dcqCcSf6gKB/ZWB3f97X/JtFVxWLICt92y6Dea76W6EbLWsr5aAC5VhcfuUUIs55
71Pfjmvcx5xbsVMOeR9LSS6TRzuVr94AVV0MLG5nfIbXrEQJ8Lwn7UdQg3/pVJXf
QXp9kIaRRedBiKbeVbvwZdCihwhrDbjk8qAFQgILJOmurjrhcENoFI0tryjX5osn
I5Y9qiSvj0yqSyVegbkM93Xjx0GDFt/EQ4oLfGBMYh7O5nfnMn0fn67z0sGCgo0I
66Fnl4hi5Gx4nMBnAIhdjSlH19gJ790tqq/cMr50ahefQM1SNtlGHa2BZuZx4KZ3
oZjz+NJb50F8py5ax/XSoSlJcf7MSjXGzRFecMZIStzzp9+Xr5oPsMDK6ccP0GoD
9E2vNt+du0XnPh5rOnYmhGSezcd8HVgtrT8Yb0qd/ZOTkRjDIWUQaZiRNWm0Q3Fs
xs/lqJjQHb+HdRROP7+S+zn39aa2lL2TwHqrwCT0ATqDjvWBDQWEVzT6d46GgVoD
CrmnvXcge/Hf7Sn4FNUtDniiNCdY2+KeedoZQlwj0bmve+mocynwMI/83zfM+pWU
EJDG73BVJaS/3RMf1YvIz0cru6wtD2nLdesz0mC8xZ/h2W0gEdmQrrgJbxqdvUVM
XahkIRpDSgOLADQe/K+m/2hh7H87V7LyQ8JGZef2/9vo6eK/jHD0LpLyT3GWyXwb
3Qp5PHV5nkRtClRItvfxsDeer/ToJ+Njx/onGOIaE8E9rdcjvaRqc4eVOvGAHSrr
3vA6VcCxTpgh0q1b3CMtBWwcHWOWjhK30z2uyCLRz5St3nC8Xqs6iILa0ikyjFaR
sqtyLyufEWIhnMCMJK01CySPEFpjO9yuT/S/8myYFtAl0Bt8ebw3Y1LEfQdML2IB
LmYKE+wqVpUsqt+O2A4xILL/yfx/3tYRZ7MllC8NRXHlYtogPpJWeaBsO4TWoQ4r
zCIsygM/A9ei1MLzAgq/aLpdbGLXzdw8/d6skmMRO2GngKbgVSrCx5w71ab6pjf7
CsOAPRX42N2A4C6s3v2gEgzXpIaksL1vfpeWyVOhEZ3bAT73XzuSCPezbfAs62jR
y6flIB/g3qdngvc9TosQgJUtKm3bMidbU3k9ZvI+SWeA6z7f5JKhEH6El5VTRnVF
um2wRCjH1QAqtUvM4j2tEcTKPmvZs/zcsNnbhFOEELOliJQpDicUmx/a992zD6g9
Z56DqhIpceRS6dPXz88sjewrYHa9esVh/UvpFrhm0xm4WGRB3oQ9AxAbTepWljZZ
Cgc0LzpLTez4Y1X//x09AMuiWMOzumaMn/OpisUXnoek322nhBkleNUEeLNEYaG4
zwcnAg1rTumBdui1hHf6d/WASEZz1+q+jDP+yAJbr3PEier6nH0ZPjJ2KtMvKNwW
90kaTPeNkJOkHSwiEQgW1Xg8OZEPygy79gBx4KWgk6E1Rr2s9VFMTSdYGGP2Y4Xm
apRH0q4YfZjCMEzltZOdseYAhloLorYWCFneFJ+c/Zt8ULfAUhywKH/EQ0HRw3Mc
Pl55bwSmgKLpML8Oe1UD7FLwkhCGloXB7U1UqDWov45aJKS8e2OahUNhLlo/vBp3
Qs+cAkYQkYp1/X7w4QTTE6qvwXBfrbEHkHTt/VLBPipNAlwA7Cp0WOwY+p2wF5dn
NTOsFQF69wqM4+TT4Hp5ax9YJ/y6OgjcI6hMP56W6v4XVvhpvgex/5P9xWB/mbv1
+8PTD3bwZGmPt+q6wiaVrVq7p1FBMPhTtcrmdnOJ5h+d3rYNJp/uXHzpZVtMJNDx
1mXn7WrObzimWh1SL7BGU849uQaZ+GpoDymLcJOPKzbQniM6sichCFyoYdmKpmek
2CbuVQZg2UpsteE+/FkuAPM/nhNsssXN6jZYUn1oeevoKew+pB5xnFmxMEeI4O6+
vUfcs/zcFo4Ftfhb/Ax6/vdzR3SLQNqg2aDYiHleh56n7TwLiGEJaWg6UFUDWlxK
J1S30vzzfLnu4M3ZhBf+szhynkoQZH79yxZbjAA612XVFbsADYN1Kd4T8QKfbEMX
2BtOEuUoa2p48KldzJsu0D773MfrIETL2nFxqFJJAOzixLlAaKsv32iihIky8Psb
+yO5plMlUxu1vsu6+8hLJJ0rZqxQcR/6dCQKaOE4+Xp9shj9a+SfmXEY18772SQ2
kvpmyD1qycCow8py3cv73pZ3Ue8mLiZU9USpQOyBjRyfkWhWaOmYCKrOAevdzhSt
DzclNgLgaZ+CQgrsuL5kWhyLVYgrPBXSXgsGnMtYq74SguslKGvtg6S8EdlKno6v
/zhaRaRLvZebCyqz5BZMdpF3FLNRINhUEIWtjk3yluN8faMEJpWEtBl/gqbtrjgS
/j8UqFjpIkX0XlMi9f7UmXk6Ollrh/C5UTII/I+V3eBqFlKogNguomPWZgwoNRV5
jEpfhbvG4H6v+5X3vLO2PYkfbzgN9l2XDhfBpDeVNwavw9o70Th5YEg9SM5MUzBG
8/aXyYF8WdkAQ2ajvKQkkdUcUUEDdrny9ZsimayrFTwKJ3g8US+CQRThji0eLQYE
QeBLorr7cmLihsmv0XybofR4XI8efN9exv3O8Uq6W+ii8wSIc3ur/m6E0NFeidjE
8qnbbkqbARIF/Bwt/jSFu4naQoGHmXDX7gMWv/Uzi6Fg8V70L5qeHY16IiEpY0Hf
QX8Y9rpgR0P/7am+fXJIl1nTg7lrlC76lEyDeeKcFRJvMyJmZIKAYoQ0zcSDI/7y
2uMRNVK+1aS2YOCAzHeHFyaK1YE0PDZyYoXX3Fq0fWqcA01hqZi7jjKq7vQmGXRR
1tfAHmkk9og8bqJARC2ok5pUPfzP9NPfH/+FZsMUvhaY2lfL47kDXq2l39q94tDk
J74DogSdLi3wooJADbW4soolJ5ARFTKayMEsKn16Gi+Q4DwAUte4IbZn8WgGAFF/
ugvt9VYuC//UgLNuh8f9ZceafWZVCI0QCUgVB3mRvnhqwq1atPOHn2XLXV+5N/Z4
Fa0HMlx0mPodOfy82opWoU3Wak15xQPodBPpC+Rfgmrj4V2yrnCdDT4Wcp+JKPdq
BKiuxaE6RrrsllbpKJe7HS8jAe+CsaaghI4YZ3dNkz9hlLxrjARrOidaZC4L6l/K
xGRngXYClgq5lA6tg0NytVIYEZ17ZX/lNMWdiic1nGcVt/RtYLICiAytiTDdO67d
4xKcLnZDZI4eyGMG3antpE+RBcxPVIuWv1zZASTukKUrEsqr0rk6xwelhT4gNgdv
4DWVnWr11G+xwbWEJiZi/+MvY2F3oCkYIJiVvkWCYC/RQeM1sH/PlKd2hNvpv9/+
dHxCPe49sDLD5cyjhU0Ccm3DXOaDMUdYns0vAf/La/uxrGdqrUHQSbFaZnD2+vGb
sS23Bv4MBS69ImnWaDTRS7wIZMqk/slqeQo5hOljV2TJjkMH5oh3PoUbrYgJ1Udu
RYiaDKoQxM/Bn8IFBTW/0blsP54yvdkzoctgFi6J/d0KGD3lXoDkMWXynmM0vS7U
yO+BN7RADFPaTXppz8/ijM5c7GpHK1kuzKcAyMH3ofglvbWMpjBZFskqZkCMrd83
7m+CgYfhpetDv+m7W8VOjPk9H24Uxs6UzdB8xj1465Ev1iC89eFhju701Wr9s8VN
5Xi5AgFz/jdnsp+yHTaxdU4sAa5gWBB56ZIMp08KPPOmOT9RoY3q69Q0fEnb5Zlq
I4venjapo6ZAXFewwvSAPx04xrNc2oOrq/e+7WuetAmm8Jb8FbUFt99UUSNZ93vU
IUSGNP3MNLKZd9HxsBj6+lsmEhEb3STdY1P1h6F2ewe3ia/WIrbTMAJcaEdnyCug
b+7nBXQtbWk4JknxteIFXwh1VGryo+gVCl7jfonglrIxnFMLXjNMvOjL7aQjE7KL
NbcSSyJn2kLmwZ75zz9uR+ixOQmKMUp+gHJT2W2jK/fWs6Koztg9MOaMfXrQiPlA
4wyaei1zNU6hT6Ynti3MHx3uaG76KWaDjbQwO0KrPjMW0ymIJR52iYi7EHjvppI8
EtSowYqwTUDZW1ajkuLHys/m82QZFxutmquGx0oFJcpC/I9iWIMxQb9UKy6uIhL7
Fu3uw49nQsQLEF31GA7v8QQ5xu0obKimaFvYzGz6mr3U35XquBIIHL8ArviAvo8u
KL4TAAFJuYhTjM57DT/hZ2Qqc+v+9E1vkVxvs+0mGqvE4kv0cpZ5bkfwVC0k2OGI
WX81DqqEDHmN49IDLNqgvOiD3iNQvxDUpOGblAAK97QFzk+TzYCnmk1WZ2tUy18B
HkoPdTNzEKqSnBBtsc2vktkNdnd90g9u56c9mUFYfmRIRI128q4d3vdAACte/ly5
RbU6blrHVOVgXM61pVAp9Seo2gAjabR92+v6Q5C3SF9a6Df9m2JCmADBX/5OquI7
nkm2OapveyEVYbPgCpw9azMAMNqOD2sEamyftkFkd2U2NK+hV2FoMx5VBx/uIogE
HT8JVNIGyTaJoit9Q4Vh6tEUyhcDYlm/JLGIAD3yxZweb0Kg0YvYUNLxBBycQoEp
+OhrcdXuKDnT7Y1zBWkCmNXWnvFeXDjeomnvoTL2GN3zdmQkQ/1//Ve7mI6+S8Dw
oddla2LgeXVi8CFkVCXGJwf7cB/kH/K3ccq/pE0Wb7v44OpI+qqm+y1+WrmdaFlh
yCLGlXHj2InLvZFRwV9jds+DkvGv/x6a9IYFH0v41bn0JT83MC5LshEgUn4+qdJr
nWQ2km6/vcE2BJCBjS8SskOK79U6vg4E8Gd52+DgRe5DZF9voSUc09e3eiZZQQBg
cBSr3HOfkfp4LGnMmQYWKhkf69Hn30V/zLxw73rwjsehmNcq6t1sF2COio8dngOd
baao1FHRloyS25Xx96m9eeKfMPkV3dOrL1a+AbN0xCfUWRZs8o2gBIcva23wviL/
CWUDk8vXfhQ4ZI7SVPKZVfypROEiayd8tWUpcUwhvTiKnYUMj1iqUk7TTZJvCTZ7
Lyum/F73VEGz6uqgHMhABMue8rPQvMGzc2hHUnZNtGj5943rZFpCv0Fad0rhz/ei
iFWiVYwwu5lzlQ6q/tRH1jXY1BVlBRJRuG8RhutJAxjCFqnt1eEbpdgqrQKmGaIT
v2lh9QucaOe6mG97kkxNZUxrGtRhZzh2N9AKPukmI4XqB9rQkyhRYC9lfjPlLzU+
zj979pCVMa6NvcAlN4MzNd5IScMA9GLr4guRNSjeLU0SnS3Nj+vF/YLvpaMHrmpa
kdc2V8YadBDeqkFuioV2WroLBgI9pAHGRQjTkxQHmCdiZ1qvuMf13/cVraHYc4aP
bM0k+TagjPmndgaqOWlHVaKQRlBDe2doYamy0lJJjN7kOFG0Lfa1sGISWaQ2/TIJ
SN090AMeLCEjcXZP1FYmgp85ETx7mGLVkET2Ru3++3IQVZIp7D8+0MwHH05iUjvC
9NV79h1EH5GJvUWYWVX0zEhpITWZvsgxLsRW7ZJ7l6soRD1YexK8BzKhXEF/ejtA
LsNAAfawQKE+LoRonJjUotlDE9cykom6t2ufdrb2zMEXpKJ3cpUXC6Lx5lO8cJxZ
jL6HE53dsNoElz+PiZqdWAWrf/zRaXYq37DPsOyf275MbYWIQ+W2Wv63mIeP+ng7
CcCSA5XBTsbtmL5jNQH5nY5a0lYSLNVkL3aCANZkU1aiRGwxqzfPugQs/Ax9jM6u
MfOkN71rJXjU8b15AdEi6bxg5zDDP2YUN4YxVZ3cth/xMtuoEB+eOvBBtH9pq5yg
bGtQOdfWFaVSpkJA5qgVuH+fYbEOBqF/x+bMAtOqfKbZbvb448jyCwVsmpZzEMGL
QuImV4c6I3RmFgA80n64EE72qlpsO0AAnoHxiHtRmi07xBFM+ZfUSSY2Q3n2/yt3
ejGx53xE6AE7dHzf+5CIuD1B9Cxu7fn6NAUn5sP4IlTp7t73agIVQ/wArO4aKAjY
aENKCKaCtH3f+QNbFZgkNWS05OV/xZ1ca03M/EgEnT/dSM0NjG5jEggn98TjMxc4
b+PGgn0ivOIiRIEHNf7wPuFWb8VXKInkY4OPmrwz6avqhFChiBiKW5tUFughR5s3
dSinhrzuqu0SUiqrgQ6aaTEDfJG6G2VJ3e9sQ4nMDo36OJNElaNuSUlXUX41E6Ym
DC7yAyTuo6C0O1RfTOKLq7Pd1dV9ZXfOY38otycgcU07OJ4MZeI4RA+8JrGuprRT
hZMOTKOWSbhSYzwOcyMzcLBZWVyFqyDPqd3AC+uMfvHwQRcvlL2OJXtXd+Z42IfS
UefJxIOu83Af19ziqbtW3Rhiaidg0F7UG4Gdrk8GD4o1wyTTBFzjxWBlXpKyS27x
IkDwQi/Q2PVvHlybvvICK59ekEdKY2zlMa61eIuTZl6/qsufJZh5cOsN9x/E66Ze
6TfuW3IzqoGH8hVNwQUf6JctJxdo+5tY3tcR+LN/BISBYCebrQPe73LUe+suCk9g
685lr9DWIRyGXFgVrv4+0XXKurYGr/lbUXCHoeQX4CZ+tJjPXy/zw/oRcY54tllP
k1ZkS0t2XNdQfI3LrqZ/TaElgUf0Ht7DQnuVhE+a/yKeY3yQ0A5Vue6M3D88wswx
O99JgE25IVl4CjsE1ATe1AWfOKSlhxfzKus00pszgMuJ6+skEGXdiSLHrmax2w2I
lJuII0yc/pU0VCQFHcDTGGArlBWyM6MNppv9rQmnequRalOKLOuCJ0ssF8hht05U
zKfM/4y+qnAOua1uWWllx6UIDR5p44v+JiFlJApGqbBNAdfb05Rr/4rEj9sts8O8
/qMm/yT39JAELfaYLrawsCjJO9sXejhUGGLzJr/3CYCyme+3AD5c00dBVHKreK81
iKMYZA0hYFiAKsRMxAgNlc/nX+boiQbc6/2pDtNW51Zk92c7P1p/L/crRBZEauXL
ePXk6fKB7eteyjCmV3zDx/qGxeBJuhnBfnV2ls1BysNvS3kzafti7Gfh7u4ge9+L
o4A1ac8JU527uZ8mO8ocWU80W9GmnKXIS8uFA3cQ4hPqmOxhk+l6HKwMW96VHksJ
4AzG0VIaunoFe54Gu3QDRTK8za+uHH8H78VD3oBdwyZP50kQ3NmRqzCim4rlxu3h
+ghO+kvDej5vaR/H2n5ckHgO4EIaHG0jWcsHAM/XJlUhDTV+psIy3eqKctkE2nTo
ZRiQ7vpC+aYUN6PiWjUIaYuKiwPnhnJhpR+KirJxv//GmRIAjadh4xCxygFtrgPj
M3N9mFJ3BP2NxxY+eQ3Y5SjAWiJFdbTwFVBYz6BnfA+5Zsw+HTGqQSpzXfp3TsM1
/sdf+woFVZJehDha1tGN7r2gCeA9Al7+ICUzTm8qF9wi8Nc7Q1qTQQ8t+Z9Bu/ns
nAcOwTiiv/UWnk293vYnM/QWMAMX5dEZcimJSwD4lb6k7TSPd5WsUfSp1gctCcQF
FsYGOlBSfg5B3UZatJyRPeK1L4r0s9XqcO+vNIz9Dt+qPt721c177lujQk+51g+3
H4N40i9A2qM6xTwGghf9vq83Zf2Pr1IUEPKmYk559VpNBi2aCMXwlZqH9AEPfuGc
DltUM8eUTC4RDcBwHWAm845Is/Rs6YiKGErD/0ExDIbUIcNVBOr6/ZoJ0AGNY30i
lDwdTsA1nyZLJa9qSTSw4xgWuzganvxp39OE/7MgNE3rR6LCxn7CzTVfP7wS5beh
pr/BD+J63nu42f6/ereZxU36kg1my48qsjcMLXJvKV76HZ+qyyATWZw9asuG8w5s
MYd2Hi6+FRQdoF8CY3QyREkeWZF/rjfGHTGykW0UWiEy6XMxybG0f0nAsHX+ux/5
paZL6LltBIauVUpgzBBrwxdNkOhgLPFAgtQ/TWPBgDQjSNscP3NW9wMdClh103Mj
Upa/Et1mNxEN6WtbQh14XqndvXq+fdYOZ2OcujcTy2Phq0S5fp/avvn360dWfzB+
J/bc2TbTHsKhiWtAhVvWNB0TQN5AOFryMSQ2iDkSMi8WU1js2DAL2ko+zRjH0zCr
v6hR9U/BVMsjlHpdyA1pVsuw7YW2hLr5NpUduu6ml4OODK0UePBEkKg7CU1gZEN/
CY9h/pROJvVNHRe2e7wcQDAOF6RNTd+9HKydHKtYNMeOlN5pqhtuVd7oRFPxNKug
KfvqtRWV7F2mz12lDrLLJ/6Vl7KOgv65GYmLuWjQwor0I6TMxRlV24CjVo0WAiQ1
N7E/GhtcEOl4nZ+5P5lpi5He4hxrVNSNVxeP0y0ur5oQ7F+ZdbxAy1xonanNBHa/
LCdpqaW1BZgVJO3IBZfxrjfZe188z7Rt9SCDRO9H1QM04Uc31H4/AoOYS4D+a/is
tSUTK/vJrSPAhBxFojFFaymYC9luluhHTLvX+VVZZUmSa+6u49VyDa8sCxJKI7ml
Xa6nsJaD1DUb+4nFIQdSESIsoGar9oBhzDloJqIShtOOAxBive/os4hjTX0KHqN3
CiTMbjeKQAOg5JjQepwvQex4SFFqQUQQ7S9KfAS1NysroOMtx95DQUGq1/Xlx9ZZ
5S29IPtCCG7tJzw60Vfac8Lsa7BUT8tIlIvxjoyeuwt6hzNWp/XQ3RKWg/Oa26Np
VOPWLKxJQx78VaxPTiUuogGtyee3uDLN3HLVUb5AGAFSwZXUzY5fI1MdjZSAIgxm
NnvFwxfWH9RrSZEVifv83Xr+0Vpn/tGpYKbFLqgbuA1rQu9H4L7kQxjJN4i3n/X/
khH/WFuMMXeq0QQ11dUgda5QXxU/cqRXLhMDJ+QMaxoI4wxSWxNpxiV43Kc0Odxl
os8bj4xNlvFkghD0yKniBcbBk/9ux6hY6K0mZRlS5saP7SR5OuZqHdDKuhHiDv6U
mbX7jcVaWGYMEbHMZKeV5S87wvDCDABk53K2LgBe4/puC+rMvCidgo9QxQMdrsvS
UKhSBy2jJII6owoQ2LWGuSWMxQFIatUJHye5eJAeZw/ur8RTWi02kQw5yWGAiWjU
3EpljbiAQkq1gy8e0VdOVS2uQmN5sswEQ743Es8CU9Mc6wiiKVlwiULAiMBK2Ff3
CY7LYzK9Ttoe4a19Y2/ipP/CLflPm2AvCdFtt/STKTarU1p9mpclfYpIF1FhZ/Cf
wQsRG0HLU1YcO5W00EWWEYpkTSuXnoAjPQhxSUcauUopoHe/ddbOzXamizW69Sx8
QEnankUyKurjDFu3VGmYYBfcqcZ94f7evuvBNgdGCLiPAEO/bknKLXsN16XNaihY
2xBJ4o5qAXO3XIsJ0L4lvlUVn1G3ySEGWtfeP0CM7y9ad5C3w2w6zBvqwfTUJ9Iq
c4qTsJXIxQIk7qlE79NmPs1sMqCC351AsGDPyZ+3uP6UoPVXuvU6Mr+Uh69yhDXv
fnDXkV09mxULiq1jJH1oS397ZKG+OVsINNuSj1actQtz/JzcOoeOx9DaTR2VkJ7x
k71MmiqhmwvEo3GSvE5E1LHkJPvRAKYVx1y6gK/Dmt+Q6U8hdnutkuwczXz7daCu
Z6KXffwk5Ey41wpJ0u8cLI6718bf03WCywvtRi+1WSXdySKc6dp4uyyOypz8fFGr
zeRgseSrKC2fGh7X1HM+wKgk/+uACGIIfwdNXmCKNIaB6LcK6r8vTaC0cKA8ywZX
UbZkXNBwWz3YKw7pyyjMEth9ov9IUtis70ncVfEitGzb9KKcqOvLnCc6sittiKgB
owuQjWXZg8L92FKxUs1uVHjD69xf0vohDhpktQ8L5Q4ZFIZz1RUV4BEq1zhTC4xK
O1r9MT/8GeUfUtVObGk/+TBNgDS/AressvAT8kXPZwSQze5KdC9nDmPST/7ijsGB
O8VSmh88fgVCVKcyYanrdFzKBBpuXo6ZGxqXW96/pjIVvFZ7K4MYILxSPu5ds6X7
EeFb0dor0TzfkvazFawyBKr7VVORykER/7KUh8KwbAme2ZEZNZIuYzq+F/fTq44d
Iwjr7LKQwgde5yQL+lgNWZGRgFuZaTIk/PDcz1lUr+NRyJ0Me0MJSJQmgpKhCSTM
Af5cvAB+Z55OvhEHysAw6WJ7Ac5M9vilV/LB/5SikSACmB2wlo+xXstMwIRMRTaB
JcgA0gdpNf4DNlDT1agGcBAbPin7F+PQvi6dLeYOGJfJiLfyZ3tpwlAB+96Hrtba
cYumXQUpBDUpNalyu6+j3XqG0rwl//0HAiQVuMkxnZDNPQKMXGxt18Kh+gFHz75P
5HDHSo2ZmzSeE2MfZhASbS/CyIn7lBrpJTUMFIyHQu8EZhmebcic3m8cOpOR5gFg
R/1cmBHK/nXIOmYDr5GPYW3/k5nETEsQ8A51zaY2j4T2hjcuJK29719eNcGOdJwy
S5I1hzRBL2P2SDHvVeP1I05rPiimsTA1vyPG7HmDoFyrBHLvsTNKRrvlL5ocsKTP
BkPunBZCf11GZqqJoXmcAsNEQWe4KuviSf0HKYMFoI4gZviXf4h7cuxWDC5lLBNp
oOR37ofl8E/QWUkWFKPSCSbFIxbldN8798zEmIYgCV3caniY9hjo1qxeheUqaZs9
xZZj4GvbtXuayRAbiDXdBx6wesI1t5tgEtnHf9SRwrxkfuYl7HyBI3FbIYuSpuKW
efRPKIc38xHfnigMS6nMYiNrcYaJZ3MQC2VVO736XN6DFTK2r+Gfi55bxYpq1hpW
leIx0vhVD/mXFlhV3DIvaF4wd7Cfh3xt8LVzVKAmv2hGglnsc9Tn5daIBFqF3209
KjEkWoYMm5LhNW6NFvqy0WNcFMilJJE5sxyjdtEd696aWHXacmacediGIRgTtWhx
KseB32CPhNP8Cl2Gap4T4gehqk854xW9rnQlyu0j7hwlYoLJtVhqPuWHZrNDXtKp
EFa93NSkgz2vcNvyV6PqvURvMrdQDTKcXm2cfW2Zo77gvFZpVDR3iR6Xd1od9/CB
R+3x4vtttO2se6svE6oabMjtdcquvUFXQP2HP5I3F1GYHG90EOMzi5OwNrLmkBcd
Nc2U9SfdvtczRRuiZM9BgAFgdwS8MbdyzNeVbU1jIaqHfu8R3/5QwZt4DhxVLKUs
XOFPqXorzPYMIxBGn83mIfKKxXZJk2WDecnCXlSt1WbGtVhqAvxtnFd3p76BidhS
LKtkcYcFGvdBNmLmkomXmdg5RL2Cny9rPP/kkFaNVOyknAjaR6sVBCRYeQ6cbesa
RPaK8IsIRX9uos3Dll/25tg5qRziuUOunEF6MWv5V3P2veYWQMKOUNuZxsMJYmtc
jgiyn883hjloiYlCLLES1GCRfC0Sfk1DxsMyCz9l2Y6+mUtO43s55ymM3yTIyjzm
pDAWVqORNDTxetIcbU7l7UtsAK+2iwvHKiFpwkt/HNzSu+U4u+XafKADztW4N/bq
s4UYEg+eclVHYyDacaDvUvMFlSB2WeyD+BQVotBLGiydJSzAzIm9rsCQ9EjdOpWu
Vs0PdAmZNDKVBlB2cG7BXVMlJvb7wRTwTkEUAk2XaV8FsLBxuDu3AXZH2/l4drf6
31N6cLt6CqiyeuVpzQWdgdh5lfI7BQRHLRMJ4I9iQHlQca7TPJf4/Db9Vcs+JOEo
BfAvtgMavllndlwlOq637XTeQKT87FYDa1MNeNyEVUQ4h5CRIZp7ST0K4FV9V5Z+
AH2ol9CrNAHWmaqj9K+EsDxfgA20SoADlbXwZPdqWO6ULHVLF7mxqZaCYFNwbFLt
OlClIKBbbRMUvrhiZtn5ynYXP6w6/q0rFbIf/v4tRn/wkJDJvpHoKLYVN83/M3JW
3BVwz/NX5SEYBZYR6/4An0ry1x7bR/xnhVOT0sv1/r/DP1iyDx794fBvYbAunxlN
a1x5HPrSf5+h2iNT8m4a94C6Z9nkELTnJX4UdNVSrbjr8anldSuIKWOJIp4MAGPq
C+LRE1Wbzpl879PiFavw1o8kV6uzwPQXGPOlNygAn7NCe/HzeNeb1JxL0mgJA7ib
R1KoCP1rzua97Jm5qzqj7kHXh0EUUQrAvrFnxfDnok/iL0sK3JlA3IHn01d9vcBj
TqWQLje7MRyyl7jqw+9Kc2AsUWVfCuUw80m1+GgEcsCBQyFNjFLcyUamHxnJTDBd
OcgEwRE4ZcLEcbG6fg4HEfGrFxz8T705xvMsMdTWgYwZSheZ4vq1S27Ov14ofl5E
S3301rGhWnyJB2fCbrgRdmJO506v0Y/BHX3jM8DzfEJ32j63hYWiChPdmuv0Opfb
FCpsmm+1Z3y6lQ2Pce41/qOphH6lmmeJVE0a89FeGQ54cC1XFnx8tZosIdCQLpkO
PaqK/hXR+Tzgc60Vd2iykCrebeysqnowoUTOzaa3DhRBZY5G70A9na2BWmjAdVwK
RBBOZho+tXeMiPdyjiR6TiLgixvad63+k86wiWAXgHOOlFuIvrfh/BQJAZnsnGbu
OSniyk/xmrNE9jfI1VwnJz94MM8Gahhce1rKQmjg9jrcXf3btcH4nA1+RQbZYNz5
f0wpMb4xrXwCCbO9LeVEklka3qlYj5+QWVG8fi0PiNh8tDd8J79bzjcluxYdpaaB
VMP/f8q6g74YmF4NPYF+uBYQ88rhSR8ObYsfBSYA69cy7EbWs8mJnuF2P3d5/pIS
4hP85xRhZ1lrfdZYzdRP1PjRrbpJstZcUclmR97jfyMrK4GpH/FKUWsoYZY6elzP
C52k6SQYNNlI8UOHbzNY15gpNNY0a2lfzhck3+K0Zw5QFbvxgyst7WW+MtpD64DM
dXN0AUhwvOZmMrBlhQzY0otwpBEK9Y3SpeKmpBIlV4TuA1bhKBMm0CK49ehQU3+h
ZPibeNtB0ix2kevcv/TUdaKsAEuhOxRLuwkwE0rLhrcise8tz2rvjI7JdUh+7VZ/
wKLL823TQzZ4o/96/2wGr8MN8AmSdOMWNjhoS0fVnhj5QxIn0mgAZ4x9EwDcp2G7
40oSPoca56zOGEd1XgHQ/iwxLejoomjlAsVd8tU5dMUlMEv7zq1izmmvHEFbaReo
xshvS2qGoujdc34Z7A4okAMSQfHIZWwOMuCONKupNsQgN8iwFYgk2sS1XROB6w/5
k2ONEnAc5bZNUKueySlr64zm6W8lMIwJcH/USQ2UZ4xVDMuDdcD4ofT+5xDzy7p1
w6/Bo8Ep4AwDPAadnu6cisnZHF9Dh9gYtIlxvadYC6VIH3ixFLEXjfS4Vq4ixIyB
yBIXQYRCWp093fgWpgtwcDmgxYPqdiwzNbhd5uadstKPPB5RdXkZgILkk0yTxuYo
8n1B67BmL2L+gtNwduKVV2HEmFueaULh1J1WVMJNSix6XH/ezlACP5MbNlRndJiY
RffW69fKUoLTmQNITSTunC21ogmexvmDpSCOrJDbHCkaZGwb8HzU7Q5VsTV0KJoz
Zfs4t37l6BIaru915rBqCu1nKTqc1Ph5ATMp+oHjQEPoP0qcX5qtv3iyO+ymzFlC
ai52XhjyJWquB12CRSuewSTEBrI9FDSjwE83U2Wgr2fsNLQSTopYod4n6TLbowUo
libnx9Xki9EOAqXMJVhXOXjvXCe3RkZmhpdxjulUnLUf2gD2/DyTBUp8LAKkABrQ
ypvilhurIfk9wwvKA7lctpKW5kGnjK3HmgOSIPFLtqXseUbvqj3KDS7oVVPEmKff
AaFzwX0VSK0Jyr1v4TW1R1rg7NDSdM8u0YcEHAZE530x2My+Ccg4tupv0Vhn7psb
M79bzsuTZ5DSkhAYsRBLTf6Xlc9rUyIgJH6e/WoPSUVGyHXurPANXEI5TYr828SE
xI6SatCqf43yhfqBSuuFF28C2e1XVW62AdzyaGhsYYteNJbU2p6chxqxNWsJvERT
8CZipE7H6+YgQIWHFO14cWQGM0uh0LqRE3OWN5xig+hmLF5H5pInlDroQe3TTZ/g
9Qh9p6LQM1msEL7oMaSg6r9X84MqHZqbdx5pK4niedVQFtV8OuG/cIKoYSQLJYr9
MDYK+FzLSwLe5Do7AodOSzn22GJKo17t0W3D/HGiTjFRBfQw0Y0D5NeziIt4oqdY
C+E8tasDmDua5hpQMSpIC9NU1FXy5CuJWBPj+Viv1n9nZrzhYKmNEo6B7GiymOO7
TME3it36phiktZ+LheHOrKWTy6/IOByMHnULPb4JwQ9fTOsvJ7jnq98wv7cCoNb1
Rqa4vs77/IPN+FD4/XmhL5TFOsbA7Q0ExCEBLc0mGxmWVibVBmVLh9UoTho9i/72
DY/vHtnWe0NUtj79Pf+BrGKqs5pLTxyoY4v0Cm6yt/iGk/0dll6mnBkV6zcdSoXn
Jnu+p2dKQ4nuczsSmBOpjWt9N4YzSVAOVtJEKojgp0jw8bscqqYgwCpNQtCxcPhr
b8iZ8HRMB6eI0Kg0IecZVvMPiZUXm9ZRu9sI1tTvVE4Ym//KZBqu+sFV0iv1fArM
R10l5Px/9OTGYRJpK/Bfrv1OjY418sizkk/OyIMt4h958AgC4N6xQjwC1CrcISxU
nB87R/IeUERhgX/pSykBgnMYPEvtJa0rbimET3vrLQ7x1tn3lJbY/KLOkOElNshQ
GBW8hSI8CWAQzx379SlqNPBHuQs7RAnVZw6wmVnRo/wLpE/G293pE7RmbW3U6ve6
pU7es3Lnbyj/45wnWbtU70gGxR7db2psCbGUPIJwr0blj+0WtrcJp7hUtSbulUj1
3CsyeaQceivOjReu6z8tqkPGODg+/4veLs1Q/8n+RGHMcxwkrfQwkh3pfEgVtRzn
ubShfU3FKvsGUxlIfj3QKEJpNIRvG8GY6Gw292waN93BzW3Z566D4ebnuHGCQYTV
dreRS0qlYsaWDT+JFYja7REQVLCIQQ7H51H7SeCTB9dIpcAc884IjAY1rngrMAoq
kzCjsTJ4JXzD/yrsTWgoG+l8iP7LzYYVuxkKHPQhtiDHSf035fqoSZP7tOVWaAVh
gb+ZUh6kGI8arag/FODDvg4RbYjImYJj5XQKrrB0sE4onJzBuKbjNIJMvQeuKlZL
gawrZzCQu18w3bAjFOdRF/LeQcZlpb4pwt4AHyGevQw5fhSwzXmAHXyLm+l3aJBf
xvxbHZgD7CgcZlz1xfgBoxvtn68npAi6W51295x1uvscJkcURCF7qy+RsbonwWqP
Cq9zdJfTXqBjNXS4dfR747+5ej1nkXqhDT5vXGtYrE5XXdPK+Hq/dN05si0iIZlt
7YPeWpxYKtekTUkzTlBgmqxnbh0qV68SCGJr83DrvntoGBaPfycodS3CHgA+udkh
kwUsLwX6aPY9ayapM4H1Grxj1k9b8kan4OpIH9P1hDMg5s83f/NClembLNfY/net
ZdG0I+gs5B5qTxKMAmTeEebXZo3BAQWI7DVpTJoy1oANhqNkfUKkTUq8uTA2ybBK
XmyEw6MTeyxoVaIt16NuVzrweyWAMX38dMxKumMsfH9vl9VjqZskVkHFkrAKyepI
bJPk0gSQrTquoumVFa50/Psmf0eBL0gWcK3YbX7XMFpuEjlEAONtS8/Z1YdZYmmr
b3ysBppmScb+ooxzSObTqnI3NaKZL1bmL5ioc8nZBcDo+zpbEwXCpESCEVpgN8P2
z8MOFlyuGNKuD9K4Qg7MUIaTXQPlC5c9fchBECgze5psaOjUzHpPZzFO5wbjJUZ+
LzxlqPE3lumKAW+M5L8Qvuc+GTgxt5AlWvKGyIdn+G0cl8UZSUcVvjbilCwbGc2A
J4k7EinQY0ZeFcBW0Wj4v8t54xEvGZiFVSl6K5n+2lJt3yhEEYeD+MWbqo7NLVBS
otCRJaDPmEK3DfIZ1afglgGoS2eoGxm7IyyRJbPov3p23H+jzpp1FExanSVMVQ00
2ZjcGBcsanI2klkpGplmLuSJOceCFUncdyIALZ+SAz1F/CP8VkUBTjbgwDYSX1/3
8PAMwqrVvU0vZU9YaAACRyRPb/l6LFP5p+091bPUQ760GnGFptlcmdTaeDV/dBTA
xCWCBq1LYIM/QDb0HkklVl4/wgyqcx+rMMU0UeyXbNr8ALsGLcB4j/dcKPgdEirk
hDSu6u619THtIGxXPlnVl+Ems/Oae1I2uOPPP0X0woouan/le+N0ZQNUB0pb0gHW
FCLKaUa0vpLx2CmD/utXBug4fuhHcBVTsqp6/ZGTgevA7CTsGo1cmllE9+lpeFFT
9i9dLAp8dgAYa0MnGw3Y1gRyBOfigXCNQsmydFsn7ZBfKtQLj0fV0n8Us48PENJh
ISOxClYk2y1/zufgsZSM7u6pybMWCRZ2A75zyc3SG6gaMOdOoYGf68iDlwsAOOlf
xSjfpg0xeRb+WXeSp1J1EvGeA8el4x1dMalzXjfziARd7aB1t83vNNmyTAt3S6Kw
ExY9I0j+CWv945QAwMD81v/9dHQClCiPNr6ZLuqiMfQpp2Le1xTBLjuQiJM6vEVa
gcgYEihUWFfHQcHgBdCnHjh/nYEZkgxyvtTifYYfbfK+RCpZ4dewdtuR3j44+llE
iGwwlWE2GUUmZfHUKNApiLlK9PLpIUAwAto8sE3EXqklAXNUBYE7tSdtzl6i4cCl
YYOY6r1V5MMz7qppO+fRTJLiFqqIznsZ/UgusUsOEg94K6yDCLTwYyqNfPuDTlhp
ONwmrBrqaoPZ1mznl+hS8GL1l1hnpkccWtWHUs0RfpKBea7UQ6RzW4qJLHxDtOWH
P8QUvSXCH3sap/sRk6KWhqQhHwj1Chp3U+bID1QOjOvegDoBG3WIhdCnicUXM78V
VljVaq0jfWrMpC3VC+24ihHMWyNPuRKqEpCelzItGkv3eQJxWVZ4EZWQBSAmuhRz
TR6pXUKeq7PnRHHgy6+HOyipTdoEKQldAlZeFyRFKiUIuN+mJk+vcFzCXYHhls+C
eMTl0c9kHCTNpiwzREPEKMJqKy9nmIuGEoeJrWjnfdbi4mH5JSyWXW6HtBFVc/hO
tyMU45zxGJoMbo9x+rFYhVxLvSEr6a4TAr8pK9NnGzh1d9UP2BTCaTU5/fbLGoOa
bXaAJ22iUa7Y7pwnHh+ycKsQSDFtJ5sd0m2D+G5WdNiN7LQOdSCb8CE59nB7BMEC
oTdYfO/mrYfxXMwCkup9Zha+oRp5KzN78SSbHiqSP9ypD3wKEdhSM5/a5nHYSeGM
aUcTDFeDkd1DtNLb2J9mx3CiKy0SuZu+7zr4H/E97znOJYJgrQabaOcj9MdTnCit
6W47WGLs5+4T9heQ0pCHk7a5US0z4LVxI7BDmJiQrYMEWq8NuS3lqUtrMeYqXgnG
gyHvvkbxHzTo3uy52q/XlpMOR7AsvAXt8uiaHZBcfm3Jz2oyPKJTxrOoEdI825RA
CP0CzTknPBPdgpWtgEqV9W89AblXB0MbD8tOEqAttagGqPOLXd5rb8YG8AIJuMnA
g9VHjzoskWYF7ayENZr/W5S9Dxy83EFbxFR97Oki6hB9u7vhaHorduy289lK/Epk
P4dR8Ol92PiUICcDMTiv7QpRHZ90rEGFwTFwuBgzesJLd3VVGqUBivYGOUccljTN
4ZK5GkzfU4lnkYkFFdl9Y5PkSU9tBQMTtznZO3K2HOl6qfPBODzA340lFLIhOQW0
XK2/zUUrn2KddNvSRAL5Rkj2nK3N0dW7pSDYYgM1mVOoGYrI5GL77Z7zNEmUhM+4
gbUH/B2RBG8ExIj3Y0gbLhl3XfY1kz/SpIWr6q1jxOLa1kV0GgDowU9UfpkaRLcI
c01X1kPlyEOFsgsUk0OWAne51T1jIOmkEdGVyw8QESBMo20My1ZNpMlMe4Za1ngp
UyJ4ABSdMXySdgQeoUkUeKGfB2rwHEJWpwAbhAnGvLTqiwmKmNyHl9BaXPBa1nAU
Lu98+l5911au1qRnbKSIoC0xgp7QEfntqT4XF6Zueu3DuNSXp7MG5A4zngjvBR6M
S4hb5Be9+4BQkaZclmyagIhvT9uv8L2XufSXgpg8W6Z9syN/cMmeKFOsgw2tlA3a
P8GdQOZsn/plpHNT4WmSVyBq6ZcJqkd3W4Qf6zMG13GFvVoPiHUktP2FlQNjONoA
NEjqK1Zzr8rPxIjVlaextn/xil5FhYkX5+Mic9zJLotFomj1xxhCfccHingmUFQs
dIe3+LG38gS71FvQNK1UYhuHJqaSZyDBtzmX0wdnjTldpc1kwBM7ioXbawkFeep0
Vf1YEpaRfaLrUWGCk2Gj0mmQ0QMwgh0NQaOJyui6SSkZYGZ1IiUg+H28JWUSJzSJ
o9VBqJ7cyNeEUcHRz67codCNrkOvriDxu5kI1xtF1FImKYpFqP18Eig2C8dnQAeA
XAFzsqn8zisEvixnh/5K1Qnsf8bIX64tl7VcI2/kTm4AqTKbpJ30w791f6wGhqaU
zYj4WM2wpBeWp1RqutlHMg9tnkysk04F86geGZcxixIBVMEmgiAtKLalNTW80wvy
ESRXJ0WH96vdwHk+sLuyuKXAGDWM9hwFs4rQpjZh1SBYqtgPJxVXwfEMk6Es5+K0
iLH2OZJa1NLkbP7Wv8hwtCH50elPl2D1ZikHSAwGkYuA636WtM4uRpW84AUUdRB5
O+g4WrzMJO9ZlmIb4VXfdg+BRrlLmUCm21PFq6SiHR0mo+L6ZigpITgPGd4Su1rM
5KD5OzcIVDNoM/KQzP8Nn1Pu2/lJ5cHDso44rmJZNjHibSFdQNSAK1v8/+CpWFnY
nPzx86MDwOE97cMYMoEmfFwzqFH2ThztM1ZSCF/v4nY1mixYpiKzPuBixO8ymEGK
B6ULow0SjMXr51ujYK8Z46xzo9nXdGeKTu2lrlzZrYmrsFtxL5Cm5h+U86V6Wa19
UE8dJXrsJzVKix75PO/xe93kflAKgyvLKNl3uQWionHD3zkMnzgubPdlXo7S4csT
v+50aZ/perhns9SdQ2ZF7Xos9X+0wRMCRQ4vYAhjZlJ51+0QFLaIp7idnn7KOKHS
be5uxllG+MGydvg2ORodzxxlVrjO10kKDkO/XJaV03aeGKYynvyVfTIWZaG6XGY3
tKEIofGqWvPCrNe/BMQrtVVSzW1Lv6cOAEgAvLUO6p/1kq7KsI6y5iK+MUqt8K6c
f817MfVKyDsptWK4sv5CAy/Xnp2T+xUGtPgvhUZj5+7kQsbFZAUqvG30/N/s621d
0FTIJ4FEYmR5uoWR5sjsNn7W8VOfMuhO1yk4ocKgvyDvPJSGrathrJyxll1xSL57
soiR7son2VAHwjJ6KXyzLaX/pLvlhFOwiSYl85LZPRj5k79wASqZ/ESMqwpRIRLy
ve7ZN2lma3l29YRWSuIIyNJQL5yZ3PGw7ppb9bRDDsX8XjPQ/5CbG1qo3M41SolU
J5m6TuY0LCVoBiJnOcabYJN+nyvJROxfrTpGuH5G4yQ6/jJ7a0F4z7ADzT6Q2E8Y
61PrRQ+aLZqP7EKZz+Y1qHjoY3oB/nUtMVWTmoqfJUY6cc8OqU+9NVyH3fyTqUkW
mCAghY9UCgwbP4on2WovX1y4FN70q4iK0KStwql1pdMibb8y14hox1fOxfSJxAoB
vkQt2RrniBQorlx4sO4d4xUHdzT3KlMO39o8XnORgi64dj8J201Qb15HdeTxHD3C
z1e8eEIWkdJJ1vdvL9y3O5hPu/ienPAt+zoYf5Ew44AjlhX70tvBeN4TbiIiTbvD
zFGgUltiDyPYrLW4vBIlgY7Y8WgaNRdJURxoeW/YHqn5MtCB6M+rgJcgZSUFTxMw
ziOvNhLfMqijUrIMbgXqTgA8Oza7DvFmOhXWww9JewGVbZ+4ELQyuNco8q8HetD/
IWo2bh9FTGzKCxAncOKxA1ADlAnoraFqcDXK2307bOwk1k7Hk4HowSjK8nXNyNhq
O5geyBSOSNgazRD0WMiIe1DdsMcC6zKKhPTQs3M0XJ1cnfvMjDmzFxELjfCXNf8V
R8DVgii5Skd6h4ev/ynO236Jkyk4fN5JNiEKZIDa+lVPvgG9+VzVTccresHqmpeC
fhd4/6HLsA/hyxatMdfpXzaWnbteffg7fWDb3t3fl/LeCSrLn1GUe7g+r2XTo2FZ
yrH5OUNR+/8EeAPEEg4HEv0khmj2m1mYKBOjbW0iwVk1kFEC7X62UnUieVPh8hvF
t/uNt9osuB75+SWa8oRgYhPm6FFdI7P9gR6XlVWU+a4ReHbvGtEG5pGZU1GRi1ou
1Y7YdRUKzk2f/aakJElYSnPh00+PsWwrY/NiH4SIKMwRfqFjLEQWMGqoYms3l/jf
izvd7/xALVIrPUuxrILG92+UnYS8wGMflJ5A9VBlsAOo6BiJxVVNXk8IZQbqTs0j
XqcCwUxgO6U5XIXd2gTPgsTuEX+UX7TWOQRFze4qL0wy8sUC28N6sUWX6m060u1O
FIK99sh0wsQHjfNv6IWhjXT6PiIsi/kStCwyHTYzlMhlPIFH3EbPgu/29vedK6CT
l+50Qa6jwQeVIma4xCOaNPEiG/iJ36nOG+pRE9oi1MoxA4eFDjhIuTHrak2SnT0Z
cfLjuRubxPe0X3RvLho4xURYUAhCemz4ADRoz5tt6GI8uuC9RGOuqgRFwfw1SfGM
WSHdwhWd8xGVCC1mvWoN3JrIXKQc7EmRXGM7H+zke1fZCsb/635LN/UsaWWtmOpp
QUMdAXM+RIHIfP4uO1acLTvihH5dLceiu017uqHquSLAppH9TmAW1S73ow42gp8O
w0aiHXG9lJZXyVV6j4LclrwCyggrpslgCrwnycv9u7N+nzfazsYFuqNPVXI4p9+t
9Lu5fKbDJMVhsmGTnXZnUIg9NdITwv8M5Wuj1BdsCTw4hwqzzbHtTJvjO8VqI9xN
M6DoevNLydYwGwkHg9UnSBoaOZ9lFV61h6JSZFiWxuJ2nt9jy+sjGBykJ8Nvx6oq
OT6DFEFf4oY9QTaBR7WoncGnMLWmsqhDjMSp6Hv2LFMxcV+FwqTUPqmvzywqFw5Z
QVn2x5976EBOwkiSMZuPOWn1E5HBybZ7DD4GjjXZ55g97Bi9X7xOeHxnmCsDzlc1
FrM8MuGD5NkvTT7MwYaanVOu+2eblawyTzU9W50C8qvwbJocndDGOiFZUvarWEO4
Rhxd0QH4D2dn4tDEHkWK9e7A8iTpxRUHuy4pca8FRO6qNtTngxErsVupYrjuXAu6
XKulYpLaVC7M0h717lA2Hm0uE2oUcykhZdQO5rimhkIeH/ILXR11PKjpirZM5FYk
TRY6iQGIWX1Dxn+vVXkqrpLPAQLoip+lIXIidWssroVh+tOkCky5iOlPg1LzNgSJ
EyK1o8NlZ4SxpE0OEOMnb9Ng7MVsTFmXPaLvei0TfnuqEG+axo0Cd1UAjpwwvn12
xrkguvPxlGOcx06qKxp6cq16O9PByd4wVtRWPFcxyQF36r5k0pE241rnwxo6MzoY
Nm4oxk0ujfA2/ya/iExGMMSuaYARGkFAccYn48XPexOvaTDpRqg0Hdf/4R9ereI1
H1pwdSTpyAeQCJ5sc/48BP5mUjM7p7qnaKoO2gp6EwfeEFsNBg6hK7lov+48l087
Lv4S8domet2dXwoEqiM/joOhK2et/+lvirTyhCw/EY+EoVwlkVPvN70alkbXcOYp
MMyl6Q6GOQqJTDYlMnjLeVXlpF4tbnXw8RxQWiK6X8Om9r3/bM7XxUbgoCuF6Buz
uF6OVC9VZoM9T0hW5xg5pCnTxn+mDEvCa7xDqRZndt4iHVBfZrWSvDe3G624L4cB
5uxFwnmg5bFYybWIbwpxKKIJy4MgekFirMcsNUJQkdz9RFRmCIyAa7pAS8kk9EGd
MjmY6Gz4e2+Dp6WtBbl4KJ25QwqUN+JWnKC1d0E+xpLJMh3sVOEZupNS81skuIUR
8OBpbjKdISgyP+6pAIkRl4/bdFUtkv0cQDDNNBg5adHX8lFovIwZguDq8HNFpPUX
kYVuglkz++eNiMSGRpub0OeerLgpx6Xp1CfnDEXffvPLJ2TQVKaIWnfYk7fWFmVZ
/mZYCHJ5OD74mAC7xw+IDahZldO9S5MkFUqoDIgjUXVOWQZpvtWikHEU+XEzbanh
RlGLzItr4SityLKLvV1nt+DIogkG8hbK+IRXw7kYlfztH07l1WUOIiFHG+7X3kqh
bnoZ9CzRrjWhDsjbj49H0FPqzDV+ibiHspdIUlsOBCYRrtFOmQ06ZF+H55Dq4hev
udyxo6blyTpuQ4rx5hef7KDDYIUPuWfcF6IMfCM+kmKNaklgkZzaUuAFNp2hrIvj
B3GpgDXpO7mWSt+tlGeO+7lXvwu/3gongFmOj4QXdToyjfjfBFh7KaA9Bm/8kGeI
eqENKd31ir79awWC4VjWWfH/jJ3vTWa7Iibn9q+4kHfw6+azh3MWHpcKFYmH6lYf
cwZTm/6EYFgN4KIaYx6+F2JKiJqMtQayinzKN3ViZcxtoKkVhyXlY1lipIr5yyPe
GL690kisWrT1u5GEe5BBgcRr+pl5fN0OuZe/wW5h3QaRSxW3OgIVOmxvYe9tpiXD
Ob0A2n0LUcx4YxZjf+D+Xk/FpJhvLUzbua4GdG3Z9MFtzBTocQPqVphb1RmmaZyl
OeCm21k52ModlRy9L2Sa1feYu1hGc+0BrFoYd6F16pHmrvAGxOneCkMHtyJ89oDu
OsVzDue9h6keYCDf11VqYso9CdHuuMmFpF8kT0JLUHyKtooSeEyP1Vzb+NK6ioz1
iqYzmeSe25fd4I9W6kFbT8JNvRSsn54kUhFh0o8Cti3ixsJkWHIiTaUpBLdVnqiY
+IYk4wbtMd+Q/RuoXlVkf3Ap2yZe8rOsEiBUQCUl/ttPcTYLVMvI9Dmdtw+UcHjJ
ikIQgme7atsiYXjQQTzhKxS++TNrqBYE1fXZSUvIox/WtyKTcsfKz8e+iLe1Cv+N
dNBoZuz/UYCJJxWvYh/CukH/eGm54RvilniGOvEHW8czpnLWFxWYcotC/OCDfk6R
Jv0TZxtsZftUZkXPgu++Jj/ZdQ7vn+y06tghChMBKWHMLYElGpQzp/XJvopYpIAM
E31QWtzvLUouSbFLKgW5FQ7hSYrE41C57Tryv8tNB6G9eNYh/ea32TfAKwBB9Y0u
DsYi25mlS/Pf8g6QbKi0eY9s2bDJoNI98n+QgzCx9MqdGsA4osIjC8znU8zB3oaZ
iiiQoFL6avo2ddgD9NWP7wXzdG3uaxDw5dDJTSGHmbB37UdC13Ir6LLHEFQ2GKmy
1/1a4BroggwKwfevGPfbn9nhruoHnL42pCnFiLZ8hAcahLph3n2ZdjZ3foTcRkl6
Vakh66mAcBynqYBpNp2M3ZRq3UxikGEIaEwkRn9Xp0i5wIz0ESDNKLuqj4AHYDj7
vzySoLkOw6yTrHDW9VWzZ98CIQxeObr4S/39SfuXKjPffo3ZLh1rrmnCjzeFfGPQ
BnzLhfXjUQ8Wzs7UV9zu0RTK5cxZC/f5dhspBfq+hAV/28Wd9nTwAxYWPDkLdbfZ
cJxIEN0lMtUDNC2rs4gMTvZ8fyRYEcT8rh9WO8r5LMllkCPgAjDpmEloS5Rqa0S9
XPKBhpn7xsAsXqbB/lDio8yY6ub6GONkZdIa9yY+Grje1bZZ3vgtRpVO50b/kmZD
LR6C+sZas30GC1guIByRqrFlGEM6UGx3gYP3XiAtvF+NPP2xzK2ik8XImTbxUQaH
F1SeOY4rMO7VC7aBDyfKyjGtuvjOWSrfesfn73OidTU1uFB2eal13zaQHK4TnlAq
xrNo60qotqdWR+gdhiSeZFvAFdxD79wrexgRnIo4Qd2wtghKA1bGkzIEiYqilA+/
jB5u+EqC714hN6q4sqabB0Ub6z5VJSWxSHDdvoz7BVmmEM/hl4F5wPaj+XWrxKkO
y7L+Zq+Dofcr1/edF6q5fL5L3qaqRXy428gJ1iY0yh1buFPnflj9CNgrDq2+A2I/
gWypR6XlBPMNTEnp/rF9ri3+9W6OH9yUHfBnlC5Xfbo1qNk+CSZuDdj+eBDV2Hz2
xByLub0FBFFBy3I6CLSKaIWQJmM3gWQLwwTlK2RswhM48UtC1iuehfpMBxfosaW0
XELhp1ZFK2AA9sBg1/YW53OGiZhZEkFbLVNroauEArtZJ5Sv9PZT6ykxxocIMHNr
MT0ioq+kfysWzsSav0LB6hPHT+HIKMOTULMAxPs0Q8Rg5cHk7lO7GFAmjLKWfiWb
Sjz4hkImYhBuWczx1x0jWrm3PuQ3w3i4kjMTFwGP3m7jx0Z5GmCGsSGu3WQxFiGI
HZt/48igymDdNGk4I74TaXM+ZOrTtoP5VMkUobW24zxES+LMpuWt1+NXby6pwvop
yx00k2JrMJi/9sZRyNwn8LrOzzngyEnAt4W5AHYx+XdzynjX4EuUzGS3tIcDA/cX
to7k4zICLDu6fPyErt1md03Toy/pstOo7JHJ6rmX3D7vzOuyhgP2n5f1FsKhtpiw
VBi2bp6dB3yuAMs6InWHheFMJvD/pio5HNlmoMgSNKha4jHkckmM3inwL/p9erTx
wtz86pwCBuUlfN+RkCZMQulGag1AT9Ol0b+M0uBHBlt8p7/+xJdPS8sxzRvTKAuv
nH2tkbGr7umkl5CdyHs0DiIntj7u7sVuh1MyXjMHub6HGJ+gvjbIvXZ0itxPyFQx
QwzDcM/TS0pNH2g3yLuoo+rOghU41UtdeA/1yUlDccd1xGk5gZzP07tUH3RQ/1Ck
x6Rw4/ATM5uujCnyHJHQ9SbP3hB3VI8lvqk8Lsw/1Yb0Txhj4r1Q+QQJQD96oPTz
Lh5dGfmYNTFsoJIJnrFH2UR76yIwx0eccm/EXhcKJtaeJMuGA41BhpyBLi7GmOdm
a7Ok0HQTNRdCinA68nhZhFy6fGdK/93Q0eMAtNuCSzvQVnk0z+bEZ/Ne6d3mUvsl
o9mAOdM4sWHCdBYvHGWIr3NY5topH2zXT33zi6biq4RpzfRLbFwfmruaOmLk+uiI
v598Ol4t71wSRG4FEWRy201Bdj/ZTfv4hc7NtEe7wNaxETQSV1eiW+ezIc7cH2GQ
LywA5LMiUc/JcprynmRTyev0cPZqBYWTPUxpg9J7mbfriyLKIyZ1y4n34P8fEOBx
98H58HpZ6DGIxWcUx/Ordt9w5FNrbRN7dzpQ5ugEh3TaIoJR/xdjdcH6/sUtHWIo
+0cUm5xDJsyEVKKMHRtGd7IBNyGy3K6+tgTqwvLMWvc4PRLW3tu9dvmJaEbgrAO5
JSXoeZFi3NnlHPk/+5L71AccXyI5nkggAH1sqqQOh8wGZpHBgLSzitFMjvdm68bd
7+98BivspXG5T9My/wjikVE4VkiEX1uRlCJyrl+E0A+T7e2/6TAPRIHGo8nQYnhO
MDUgHuL/ZkLCfSNyz/6DkBIEz2SsVAvHkqEy1atpOYmeUkzgiXVJrF8vQGFRV5mO
ZpHMEFftH6uUP3Pnsho0nsPL3Z5CaR2/8oGOnmCsPYDWSf2oyP0YFYYklTk1o5wg
Gn6qP1LQFjRagaWhxRchR3nu+4Ajb2IuQJ/nAUBEqxDk0gzrArNWP+1GMnsY2D9V
RI8bBu6o5Nh/avA5BdTYrMM+fvnh0s2ZqPsNggOsZg+Ro/uqwBXKcnkBWOcZ1T6Y
z/slmwZtL0zBP+OWdM5h/An5HmLj7XK0gMhiLeVW+uHqRUpi7apVhbqahfg9eliD
RPH7DnVJbgolahkGOR/fzeVrpfVWL8g80VdrLSTwOL1ff+3CSahrtw/v5rPtjGGo
rm+o3uxjpM3NJ/Jyw10AGs0p851gz5VqbLN4Z9dCw9HfifEVMfIxOlIVs94Om7ig
U1NdrLA4t9M/7aQsKOTxSWEJB5rUFj2+9b0t9LtYBgh68woMcgtnbbcxcZl+VrI1
Z85sVJUrWYKe7/UlKgZfXcCaHfJvdmH7zK9BWAK59MeEroNvWfYCcM5O5/GE828K
lGT9TWqC/FjnBJrQa/k+rYWiO2uL7gY/h7fw2YnnZ27bNpbPbpKiGW3u7mkbr//r
59YyPVQFVYZ61tmNRIdhGO80X1QkxQmj52YJt+4SGOeLFkgnQgMMDVxWiFHgvX65
meA4Y9mkQ6flziIisSTRxrPByWNWpvEsJGzFBOedaJZmylI5LMmD6cfyqk1CrSpu
K0SD+2yG1OxRYW+AnWBH15/QYPrk8e2UPIlXIi+s3xnhtJaOdB0j44y5VGuwC5nB
eW3ck8uZpwrStzpqvxs7ID3nsGG9FnjF0b85ZjbmGDqNOsXl3pp99qgs0HKQZZkQ
YWiDmUf69d56843TQkG7/58c3K1gnQ/SPrVOYjhWxfX65d5A2LbGDzZJHcxKNMie
Xh5KDZWBGTqOEEf/KO/gR/PcD5XqybRqtZLyby56MXmpG9X0DOGXSgU/KgRx9inE
3GNEhGF7PvNVvH1cK2cM5pRQqcSSdniCyq77zTbyBIZ/AaErhAVl82jEcBrEvTBt
AvFvA4q2+ImyXCO1HlenV26HW6Eu9S4LpLwq6X4ECABTRL8YLtYUX7ksiPMstp1+
j5nY7v6BSgRA2f2jb1oQBdSIbJqj/2+Op+zW+822nhdoFJWocLAjvmdAWRsrf38m
GWR2b68F7A5+Uw371gInbjWQTYtKIhDaL0TthpBEbcPYeG5E3J7jQFRCqj2MeEts
AbUOVms8RWV2pfYhpmYgd/7S1J6eEmfe5rwAuxG5JpfMZa1vmmraN41H/ipiAcay
8x+FAlDsA2vAtN9hEG1lXVi80nSozcTbLHK++SXI/FOlSaxFq2yRq24DDM1/ePHE
llDAKlppQEJ+ELNBHzEkbpo2Xbb3Cn0DIn6LIxoyuE6/hUnfN2qtCmbYNa/lUhAU
wvCvctah3Xu6WgkSKhcDQn9/wOouVlyrRek1Hdld2OcOCDY3cjG66oJ86aF8/olB
1pzxQW/lJf5xpmWLSZyNHHDo5JncrWFMw3yZDXT90dveceBHe0q2wAJrtPFlIF3s
tX88URVQezWAxad1pFPbuZk5JuIjshQJ9Wz1kaFt1kxCJi09I7IJ99ytZrRIzr0f
UZaVldLyVJAPNYfSbVurx1edSafeRyONqXz4P0aWNIaX5J8xYPdQkNrP0Szd4Bh+
erHvCo9jHaZt3u+cVrNAjx+7ZhFqCFidH5PNTM++KPeKK/4sdY3/qIPVaNt23ulr
hQLLu6LPqr/VooQJ/M0NU/KYmKtZsCsEiX60sWHNUYZ4mZzXA9PLKQYZT1GFOf9+
SK+DhMQG2witpx6jZsC7ofRf8LKM2uwFuJSgHabxE2N2KLlQhZmZ2t+Z2EuzBUM5
KCQSpTI9UpWVDa8lmZFzxdIZbP+/c3Z7ghHWDkcYUNQNd/8iJCQBDf/6vqCUqCNX
kqwJRaBlGOIkpSvzHYqZVwhx/sZcVW30BXgU2MHzd1NCOugvYy1l1jDYf7i7dkIn
AO6RF96G4dyO9bqsHLXqq4YFojWwmA+mvjnSXWSn47QxaCAtSlQfQb0F8T3+rIRI
FTeMfENUz/2KVpT11ouS8TbBNvQVUfJ0zfFUURuGjZ4YHqwr0v/6y2fahg1/i0YF
vLQHiuN7ExPz+Ysd9CtbBKNXUSmiiASvbgBzMiEzWldh+QXZQKXiTbJ2P2ARyuwh
E/e9H7S/AjzdqBNq4thIVIju2d1E5ItgSSVlSZVdzXRZtAuf7qjpsAbmBVrjCAB2
VU4MvdEH9VGg1D+crG0XFH9jsCXRSKXCsJbNWhUx8ERAMyYiP7Yo3Yzy0h0bNl1w
zEjeB/7kwq3LR/wXavulzRoFR0QhhPnMqBdQYL9SvnsCyOJ3OV6TkaB6/Dq53ouF
O0Qa+gAc/hEIvDtalGHozaBsmLMmErdYusO7vfmzBI708iQiHLpShA7ooRe2aa8W
dmuALn/J1osCXq+ymlfZ4pRPfeU1rlvYV5LVmWFbad4+CoEzMVWGMZg04wxaz9qL
aOPgJ921qj3Bl/m71tzDcUKoGrqFdRncXIx2ZQhJPzeJx/8QLWciGraSTZcoAuun
DZLPwWWjE/GzGDXioKbnpSHsy3dIhv3+hNc/a3ITORRfffoHWGFsf4CEt6wbdpB8
Kx5myzEuvrZrNuTbcX+jrC/Qjdc7xZEyAGJc9wdkyvAfAqAStEEc3aTzQFjG052C
zpvvhciulsqyprZKlA7ltzLoitOwUtDtQ77L4fZomNS66MzSiG+jVgKv3dv66Db3
wElb4NUHOtupKdG6Ko8SKap0G9iR0BlgejI4UGYlmJK23qQ8h+DCGOAGdmPKKebx
Cfxxl4wd2CJkLFBrl3aEBEwu8iXW4qYtAmCZmtn52jvKQ84Q4Ti+dS6kYXvl+wBb
q7BM02CsG7UZfj/xhBE/YGVa1l8UOAt2QYM5kHcTinPk1yo36K0KCOK7hJ2ByJPn
K7l5Z1DXaa7ql6iA9xTAunISeWJN7Mvwg8tlA/yItWbxtt9A3SLXO4EOHM8d5aSl
1tkIv+Wf11WWrOGhxXqYVa6wQ3h/jefRART7M30s8u5UKukE33WdKE62+kMcI9C3
MA41YiM3CFb5VBoQpg7HwqYkJrmJVLWfFGGCEyzIUOPIg+h0wQAsH1PlKLSTgshU
gsoMtYy0hWEDhHhzNgf1ver29iF5mKbaT/zuyummxcArHmrRa1aP75GU7jet58gE
iVBgYT7Xgtx83WM9D4x03d/3pY/1EysrK0SIzLblQ4/vkNK/q6EVhiHS+qFkmrTX
m7e8qwVA4uUrb+snMSkyFL6XqtGDryE+hxTPoWDyRT3+AaD3LC9kxhw9AwsKBFK1
0TNEPCM9cbcSKZWIzY2kd9w8WqGRtwvcPuFg4LcNqL0gheFA3no+9dC92/xmXttv
zS/dT2mYUvvsuD/dAJqpn+p4TW2RhK2+5zw2deH/N3HYR6AcZGwMDC0e4dDIxsUq
EyyD6NWUPN7KARQYCIMFcyhCm9rEQypuQdAxKuerILJR0ibfnHDJs0h742paZyU2
eqcx6LGKUAMBin20RLv8eWfb+pFe3A3BHBnak1pL8oFTWH3QP491LHltf5rEVDPY
rVVdA047Hev6gVQXxIRhMsEN6EgXgZcnJyasjYkIHgu8X/We8FKsCZ35S3kUrb5m
jKsj4aosXIwC1ddMVO+U22SJV90sb/ieZU/00TUtvKfFm14tdfXIYVxRPAne6Grh
U2u+2hRixSQx8IdfSHTfJWgWOkpI7S897V4rl2O7iNZ9vwefFV6Hqjs0WY+sHS5l
fQQdi6JrWJZnzDbccQakDvI05eytW8BOVMk/AzkfVVMsXs1ux1+Jd/cR41ggIlo9
RzagLg24TFY1fTnGFtOEs4xb/Lc6KYCLmsE+I8F/Y+nZdQqHx/Uw5KBi04K6Vyj/
yQ79E+6iY3Fsx3f3d0XUBuWF7B07wiVTjLIFnK4OvZMphajHFxUQ73ZCapRI/ssd
r6/erfGfUzaJcdgUwDodOzZQQecuu4c3zodGHHeHaJqZqV0kfrUWvWg6SoMJPEII
WGbmjHqS+RWnNSYUlVkEg2o/rLehwZcpbUhVPMQT82odccmtVGDDxmZIWpFjmhGD
s0WKtZIMe3NPSvyq6Ok8Dx3ZyJs+FGALelpVvwBE7eAiGtrijZeipUYwJcCYbw+Q
HgppTpp8x9aN4FFA+hvJJvXxvNjFuvgjbN1Wz0jKVNwTwbd0j2m3jzCsYbH0cIM1
0h96tZuDZ1pYRIGRjHpxPCx76MZKbaNZ/qmP73ILCHUU9SCsxclvM+2L3Akj+03B
NsJe1JU9iNa84wY9CAhZU06NX15klQ3whnCBiOxV0I5GpKNqIf0oWg3l66LsGju3
3tNQgg1thryknak+BFWq6shHifBnkZ+SBDcqY3pxZXcfGNCo5zJYge/G81ADKaCV
5Rla527qcFGE2h8kjAuCHm7IC7vcrCskVV244seoT/whQg4bIng77u0XRnMgZPNn
FDnawpdEBOMxsrC6QvxF3lok5qMikV0A0WFQkgQzBp+opTTSEX+8kuTKEWv7obpg
bzIwEqjYFhMhNWkdx2lu2g2AA4mNPgDTTr7jXGq5k2zTghg0JSnbbfr83vx2+MgZ
kYfeDZFhDfitKKBlYIvih9Osn9XhfNY1gMtvPtfVWCxggOeKriO+BFUUO4he6W9M
+5O3Tuchxv5lXnFNkqU11jDnMZLE6oDtvhiv+6XxK4r58ME9jkXZqYNs28p8Y705
TrFGw/3v818DEY+E8VfLPipPqDMYi2kJWYidntvLbXSa+VcuZFSE9JMIjiaZiG1q
3mYT2vqlVUtjlm92e77mksEr9cJNfKiSDY4hzLgOa23LlJSvrrSvoLJxotg8ZAln
cUhn9KqlerwKc+tG+WnidRAa+kuOH+8wIjBOVV8LtZrnP7AJna3DUFkPqyRBKYk0
rZ3gJJ4j2Ym+huUXKmyMmXHdVMgJBrKhSFo6EMkG0e4+K/OgLkQIsTGr08JXykRZ
l6kRq0PGn5KeFzYWqObs5MxEJxM1jolAB3v6a8Hf1XkFQgv4i3Vm4X9a7o3N9ZM5
1aYzlzJkl7fFFRETlB1z7eG0nu99vyrhByvyJ7bO5iEdtzwjB56amiO/M1gsbso6
HpSzdqKDSNTXkMJ/8Y24I947H19MPIGkXip3Aaszrz3anCgLxEujAN4XP1nne93n
FiXq2i2uqvD7Hb+x8cMYo+S16fCz03N7jAPEs9S8Gy3q+kA6jIWgV0KDLWfp1UQR
1ibOr4a1dH7WHSsjfhv6VE1N1j5Q+pG54muEqJOb5+oaYeP23a9GsfltHUSfQ6UH
uqOqwOSLjN4j1qmFEUugHGmHyW7LP4v8fKdvI5UI/yNb1YwHhqisPS36VzcxIguD
AOLAIy/v452I/YqfzoJK4Z1+z46AoKJmIXgX58V4eFfpZQe9igAVjLJtM+GwRkX/
ahmSY1oE8u7Ptr4nhpOk6/GD/jnKMyPi5JIcqKsEjyCY81kE89rT02yqaq6SFTMh
ItaXTYHWcj3fsUY3MZoGCD1SSUn67kHSKvxf7uYiQdFXhCPYukTy6xrPQv2tq5Z3
3UsmUqi7epQtoiA0R18GNtlAT9+3kFr1cozZz2yIGohkzQpRfWxjg/76PORTmdTR
NRLJcuvGgKPRL2X5Hn6oPOdIRVIrW5yeI0IPz+vlJ7MiSZYCFSHUBlS44eSb+ZbY
FIW73p7SQtr5te/Xl6spVs3cVqnxsfjNcBQ6skh1NMYFKXx36PHcVXHjwV5NIjxJ
x4oPZHSx835O1UKVI8HtLgGfu/pdEUjRsFb5ZhRLy0fPu9tjNDIYjM4HmCUaQOOC
etbJksV3/fVJ2HOigjzmgLrmgIDVWuFD7dhpabB+lAUbGUadrA3hNwjzytzLB13N
CIGN8rpLa298z/g0ZBgYr4BRQHK26vMsggqH63m6nujX6oQXg8Mo2ePcMWUVVwEh
FT6S7xoV2jPlZ6/1SHpT1RWU+fTszV7P2M/VEwXEzoqNg0c6T9bvoDPf+WqMs5Ns
0Um4eUmGttSZ7fxdzPvjnJJZPF3bfJXdx104H4OmZBUgQa7udDwRTO1UcFQHUYjs
IWKCwe/vjIWCRSmZ4eZlSoLPpsZ/Jf/l4bcNQma8BtbqUj7ZiTuAoQxW8nHE5Y9N
F9PO+eITl1xSCPIpM2b0G29WIn3X5hxWYLy2vufnBae0BhNFxyFJsBppH1ZauQQA
9tM/8dxvRKiRyLO89qDHirsF4frcjdFly7UUWwkJtCf7ejawXr9UXyPi9fT0Kc2d
dQPcNmmzfE/zDa4nF26Dtfy9Sid2RyqVTcJzD+kQ9Y5aDBuL0p0Da0OLdgjICyXc
z6wll+S9G5oMV+HrgsWPGEZcjARKlX+ji/He8eKtfIy5B8PJ9zKeYyMltENkoqE7
8oFFKFtu9fi/45G1sQlrhekcBg23DEx1j7J2+eBFInW1aWL8C6VuSplmu9FR3X2T
SerXNPClC5nSMZ2950krEd1GE4oNi0Bqt9E3yWG4xEiVfs8AK3bSZK2X1tgsGLLa
FLPcoqE0DlqKBZcX3ctuBQ710XFS/ucjmdnEQZtF39vRQfxKBC7Q95eE/tOLru00
EGT484I0/hW94sOLNZ0j0J9CgR++XopHvCK0J2oSMIGVEEMmCWOZrliKMFjcbIxi
gh1+WvVjnA224uHVckpO8m+zHL8LxoRYz3A5yZsWrkhJueyii6mEOAUA0Ey7vd7d
taRCjymmzirEKK49UG4zsAeHA5etFK5sypPaKRzaxfClPo9JJOT+46LWueZ1OPAe
G4qMAwzP6aQxVDkV2eeIfmTbvw9XiyZpTmln5sQL0AkS+pVc0YKPH+menmyoNoaK
E+Mtc3WPW5SMVs4oabV5LdMii+dG5lvNlkqIdHkqhTx8Wx2rlPqgTtgEDqMiPLiR
g157gF4EUn7wVRZVsyBXUzL2lomzAown1bu+wSkT5ezT/kZ9G5WVlNn4naGZJGq3
T0Sn7w4rbJHv24B6S6b6yO49/9qb2L5YkGMcujea5N+DUq4xGXGPJ5evaBLfcui6
126v5PyKg8y3+X2RBSbsC5ujiN2cGGlG/Mcd4U9Cg0vgDL4hz/TUFzqBEvk9vVie
a+PUWPTEtB2luHzGCOpi+AKlt5QfmMTeDCn2GfUCQ/t5QIPmUIpgNu/iQ2zhBX6g
cxYPp+GSI5o0hecg6j5ierh3AEVd3HVezKiM+JtcVE1/Gz6rOhDR0XvR9cEyPTFL
aKZyAJbKyeCaNu4V/604eQ==
`protect END_PROTECTED
