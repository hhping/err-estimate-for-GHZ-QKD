`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HfROnVfUS6lbF/aDXiqLlJgG5TPduwVw7PphSSVGZCoOfVWZFxV/WjHruazIMxNU
lf4ixFem2EKAp2+pyRxmiBSd8GFEFJyLNlJmgoRdfdxWhoakge/hNpa8+pbTzn/r
oTHTrsQ166wjaiM0XBoBW7oagOM2YMlFTIFqQFHlpuPZwvb8lhjA1kRjDJghb/eY
lyNyDVJOMzlyYnd9/QAs+D/CBN/bc7W6DPpTfZbe6aVmyrXb9aUTtknvDzg/x9j1
l4AU/Bz3N+4kqIRJa5p1XZQKw1ADIrz7zNIfoGv5fF4Ctpg5UyU7BgivOuwt8YsI
+PSaNjW7py+osghaRHf4TPDsGCgbZRvfxFH9son8kgERzOsiiWsF3MP0sGW9/Shy
+jy3TrDkoUu7fOTRvvbjRFKrjuqb8RwU6/uJS0wqfgTsmxffLHTJFFsOy+A11Wqu
u3LuGDAvIs5MPlHkxJaZmw4rXHr2NGC8Bvq30slz9aHyJt6GeNElcU3NLcNS0bX5
a6k11ZqiS44ySkV7WYcFjmW7x4N7fyiDf35wwpC6rEBB9TJiRCmgILr06961wno4
6adzeGB4/gq7g8I9hSAuxq5ra4/Yjj/PtXXtlw7jvWSVuYilehHShTpDoAZ/HVge
Vn6HSKHfKXKw5frfqWBUjIuiIDU0Y2BSpwvuiYCvZ1+HEc+m0FxwyTzLx+SvuZay
c2QJgmj7LQO3bxMchBkdNk7Bvl2xXHh9WB6/9MQO9VJ5gJ4gs6IPvGqlI4YTFWT6
b+5i5/CuEVI4z2XS7PsVJyqY4ldkIt+YAVPI+kaaw4FENgIn9K00OlDFAAX+BzTs
IQp9BbBTz1ZGu95fmx3SxvtYVS2LZd7wZMV5RoSv9KQmOnM0YZH4xqwyJFijvQAy
TrSC6ThXMZWymOuNhS+HraF4JdpMwGdGr+hukao7m9U1lQVs4HBp9i6ENbrh24S5
+I9s+B4o/zmJ4kG0nOCI8Fq0HHDGhZCLedWW2uILbBzkApvjn2pL+jVZoODCkeha
vkRT8hA4bNSblX253Z9uny6VFihVB57hJ1tOeir3mJFVNEo53pd842VoE9K9xjUj
kEdk5HOzGeqrds0z7pV+RMOMCU0Is3xil/QLcYYPzaDaExgLFP+tzYtVVvdXmhtU
d1fVjGc9/2/G6Peht6hdWDiIloXIV5LJQr1vvMlNJVLCmTsXU+IASUw+Q6XUMeNi
/noCdV5PjyyRnCKOgfhzFV5BxsImzp87pKYoE1zE6zsjNIx2q3HirmzcgPIefWHT
3/pDYSjVC89fbFIfLh0ZHf+cMv8rKTkt2iw4dC/h63EVhqMFpf2Et5mBEJvM2pyJ
EkTymfx0R8DYsdWjBCL/rFzgUir93boir5cI7WHrUmgFez3/anWf5KVdWyGhfDO5
/XGVt2BwcyqMxgKZiiFcHdOQ219fdz8sVT2Ye/lShl8r4f7duhfjVsS73YdAOHub
C4ltApt8sBW0fz9t6RksVU8hAcQS4bbxqokBWlNPt46KYc4HkloN8WRWWHRoE4r6
SATuwvfQjEd914NWtuotYqnmMstKnztRklxjvYrG/2k9pSBLUyodAkiKLh712oW4
mQmArUVhbzIYzY4INGapcxbXajwO/1jfVYlg8C0670bHVdf/AuEEy9lvEmFTTiAt
qG/9n4LORWkO+urwi5VBfI9JfZarRWMqI18sxf69NKl9UnVaQjSqs9QL5Kzvoobn
ARLMxsk4M+31BQiEW1qbXEiMHyn4zafDD/swunXxLJGX4WdGln9Oq2Y2G7O3Ipnk
FIPNB9yfhJlC1AqTBxpQ3DCuTPZ9pfbB2dDEJEhOvSoMxWBK0YoJEF3iPRnTGFU5
XkhKzDIjreqPROd5+gbPc+aL76/pmbJfphtZXiicHly83qv+2h01BpSMABtfdBFB
wGAxiqos/ZsYPoLc8suUiu5v4h4JTCPtUeLACo637gy0vqJaIgvOjTBz9hSr8MJ+
KuwvZ9pzPM1B3+ivepq6mZ0yFn+0OAaqaaHxUrYXn5tvGeCj0uzIisNLW67XKNQO
h5WAcidK4AFqOF2gZhKOAM7w9BatxJwvVHQFYfvqiods3PCUL3ZfqbRMLkD9l6qG
aklfSnhJDXKjdskYdzA/wJGlLMj4trRvT/qAoWKSxIzM1glzVKYQLvjk8oZTtVZu
dK3qGimLw1wmQB7Rffvmq7hf1F+67bYhe+ZVGExctvG6BtvXlv1Nm877rF6FiF3C
ovzG1lDLpaoUqWG+XHCiSLHcAvq3mk4enMTwDniaBayOzzc8njFlzEzvEkWrrWnR
FSmADH3LYCsjwWcyWUjOWp9wQ7UKzcOLMxchYdi+PFRaZHrq7TY8ow/tE3tqACNl
OWUT/U1X/Ml5+SAYodWucnMTAI5JA7NI2rVj+tNmmVUPrVUWgH0vGlXBWjdOpNv9
OJt/tGmMRz1P8XGfwgS8MmaGjKkKRJfwz3AZ3WpUyL3q7C+FOJCwM4FDnLjt8jkS
hxEABg0TMU+srNBUiQY0+57POREb4n0WQ9HRMN9dZkIAVzXZsu8mM/gosC5KoOij
GrHEHoimAXp6cFo2a3hfyncYwROtPbokJXOqNVC+/0aTusaF917c3diaZ1T0ZJ+J
EazL6nqghesua6EdOoS6+6z+USfAqbbVGVjjY4l/kmurEyvbnUDzxQtoDUoCXHro
CpXt0RbaApAr5hB1KFV1+1N+j+5iwfMgNbncauU2zvxhDw3LvWoCKvXrMSmSNNOY
uSgAyu0X0HPE8pmiAY7YFhodO//vMRMeMwc08nOZxB6ycPz7qxf7k4Cr5DJUCyTy
ucSRQXDCdtfnYN6D9Kp7OdEbpJDLTYwtpZDdlBhYS+v1n6qLY/YQ37YzGDyOlHDz
AsyUbCpcsOSxssj3/2J0GjivKNaQBzAmx6Az7CAc5NgCNx9XQZuSsLfElYdIV1QX
FwmWJg/5QWtAtcffX/4DGyduPw4z3dWVFQFma4vJWAJZnEI+bOP60QlW95s3OsUJ
4y60011krp5CBuC3Ic9dJFlugHgwJ+r1QbNZBzsez9BH7bR1w6v0hbyb9H0f6hDt
hH99B/bmxg5nz6Rgx6XLaTp1CvIQsmJevYgQ1ycg2VkoB0ykFEQUPSjn/M4vY04r
YHEtiZBjDJ/GCB19oejwmI6MxVqxWOzQdiBoubxo9YY/n0P/lRoo2ROkDnt3pf/I
cCtklxFoPGkYqW6OwcaOmYay7us9jEB3hDBGoMi75jSbPuy/aIkiHwUsiF7S43wb
6POl2ARR81rXzmMx/OkHf3EnPcaSL6rxXZ/rMUXRUZNmDdRcNBybKn3DFu51I9Lo
uwJ6pgfW+BG5zz6xoTUYMHxf2V8j8vxKLGOuPEEAapW2BGMfeOoOQddeH8L4YRfo
pAjy/xP56orMI6A+trk6c2yTjOv5Nc1x0f3DLV49ttzAPpsVytdCEyp8YZrsPGZm
3ToDTeccQujHEKEcKYzU44/d8Pal4gmTmtrvLdjyQNNmoO8guKhqZRktpG0n8r6c
12i7e1WQ78YfbzMbrg27ycegk6siSppTlsb9D/MyDzZAkjBCRMglAJioG9TBg3r+
0D9e7rwJ+8RuVXg+cFGccnd/kmcX0O3idiqHn5jhUi4YRiqUYsUh7evQONROqtoo
L6+sN1qHV3StbWTBaHCn5ekh3AA8yacN61JhZt45467VnqZs1iaYmMwghQo+o5vI
TjWxRgNF7UmqpEoy0zIVd5T26978q2gHLcJ66ddF2ttz874irGqq8VYQq1wR2RqQ
Gx6ksMbshO35BDg2kIpwa32pNXFy4bz9om5BZrN4MbG4DYfZlkF6lfqZrcGNvixH
Zs39t+bDVz+Jv5QBxtojOp3dQiIxBkYcjz23wWpcdvAY43hB/YkDhRXWZgtzfnUL
ARW535OTsyTeyN8yhlhcqe164Md8bGTBgtqpiA2iXYs0aAutvyFRdUp9YGOLV0wR
Usg+Zw0PkyrGzWFSAmRCt6z+r0cvb4Z999PuzQ/AspRA4kkzu0ddkpqCHM7XR1q6
kGbfeanPnC5CMcQtPVOpzt58bkpuKr/CgfsQfwlCHOQxspuEKubrpd7Ch1U9eFwk
ErT0zcMKfjTKJWdcfoi6jcGPU/9W3RE5fWgVrC1qIn2/EEyE/M5OdtuKs5aihjcs
dT+wo9mI5RTaQs28vEf8nKPgY/AdCIziFcWQ/B7noM7zDHb2lCDzs22f4sVj9Iyj
CNQiptf1aImKxS7jend1f3bl6eA+g6bq1chd1/qjvp4rpTqot1+M4+BR4Rzur3eu
p+PK1GX4B1o9o2HtZPqQp/o43SwToArA7IojBXle8Zb/qMYZ+/6qE0J0rHSlpsfV
W501pC1yK6mt9Sz+eIi95PAoKpOW9bKolakv/Xq4MY6uDt+pzfEQjKlztBmnmyss
qN0uiybPNy1AIbzowpMPuOfhCIyt+LpiG4Lf4y/3oqzriO2Di9Nu1ABwAMNlwSZu
0od+h+CY76+GY1OrSfzTBn8v6bdH5+DDneqCrsGK10nQR6lsQtEnpUUWKUda+vcP
ixkTIpVyJod4q8xFjosYdZ+VG8lq9MF+WJWLF6Jq7WvXXQyeLuJNEDVA/t17NF0s
d9bsxUZUGUHXBimDdAZS7/QdEDdAljLYci3jp+WsjewJGTQtwaiXi5oUKkn1PVLf
w4ziVfRlJW4QYKftyc93nATXiVh60rgzjf5FoNvnqHKDMccmS+BDEvud0wQJEi3F
r0OemgC2xcreYRs63b/xfbvNElmfsBszF5IkoSfCCzBoNfSiUqaX/S4J5MXxPlyU
AP7T0QkxTcYpSSu42Supz1+qpF3Bk4GWtzC4728I8OCWTveqUU38fg/4+eLOZD27
FHQfGBYmIMDl/KGdOyouo06KGAedgDJqJ1dbWZAEAZ0Ztyeu09bEsNU5GM0rH5lB
DwDldT7InfEN/Hx6/R143PfX7pbys3JL3YHXb+vLVwnTbH3bbx4T0GcCY2pzlzAh
WtfRO/Ure5gitwN+Scj5xEBRQ4y9uprB8qLxXKizSGv9SUBkcd8S8Y486EkRF2Gz
39IlSXKsW8AHlXuJdAJBOpgmcu2J2oWeKCgdUjdZbDKfJc5dQPUoWOH22+pbq/Q7
ai240sF5adlKx6s48ntVTfAxiIhuYLe1G/HchXf2BBMOhxdiY40AMM0w5XMF6dFY
e0XieG6QgR6AaqyDXVS0fhTBH+HhQlVOlwVEp/+1IjmZgRvcG4cUHA91OvAuUnLe
EfiiReCf7wsJRvr8vq8VJ/e0ct7c43ENe+WrDlprmsvNxFAK1t35ZS3hbyKR4a3S
pr5pLVliEEVl9GnWMS/slFnRk+th/4+hecI+WU0/4z5aknbqh876K62NHg+SBcei
2jpj+2Pno813WxCQ41ucIqHzqCdhh2INnGG3e0kQZRKSwW48mz1rzG1rJ6fPYiU1
UtvLgTeET3+XAzBL0N8F2mo2AtT5/7f0YnmX9sT/zrkYRzQbHk2acDNQ6HDfRuc5
G8F3Aj4dVqcGVH0vZK2n8XCHyQcjvgnFHiYme3QWq+FmlDZxiJKNFzTjbVlcPcrT
GZSStgU9SWNr7VPI5VaHGaL0H6EujGUZLeKieznznkhkLD6gSCzIWpsuyXK+Jhfx
zZP8t1RhDKuSXpVQLxBQZu7mldCekENxUZxzgeR+YVHAWU5YCtR5RsuXSA5LhJOu
7TUi1mp50R21TorMXe4hxt6LD2GRMKKZpVro6irSry4gtjgrjtDo0TladnYanVRX
QaQT8wQrFfL3qBG1YhrQbnBpxiKVV27DXsvdRnc+KTKL2aPfdVMFY+DWpuIKKi6w
nqwccIbLfR+PEEI7pv/QGz1hMLb8SbjnNhmiBcU7lJEcoHxZ+Ot0klo9oEMlz5+4
Al91x3bIGio4oFjjHnvkJOaSh887dJc9BqSdtI3UCB9Wz3zWoHIzQVHeZ2WAg9zW
esPIqBoQDb0VNpz/NpVYuwEExAuuwv9ltSpDqU1QMZf+ufPNSANu9ySefGt0iaDe
Br8RKAOE+EY4hvdF+1gUZK9T/khQO6pHuxlHCLe4/ZTwMK7aS8asRRVN3rcvme9m
0UMFVA4RJLzJfhHQdlg6qM9KVonF2hJv7CV9C/hj6/9pfVOX0aHHAa+/6uR2ao4H
oaC67v0GYWKwkcSTCn9NMX66L1Vpsrx1tsPh91F/uQv6ORTczHImvA82Yum/fGjF
r6cbhz+S/7zW0N+zngSD45RpkridK7jSKR1fjlmNIr04WhMv/PZgRgYh0SGn1d06
eqglTkvWKzccD7ISEoOWT6kcIXFJ/hwt7g0rYm6wtuaL9ts/2XXnT1EuymcGTCh6
yITmmdgJYqCP/FqH+60WDiQu9DSaTeKyXcAnjZFyFu7axrRKrJHPKkdWigQS3FIO
OvGt2ORbPd2REVVtheQYiPANO3MxVP3UhMIQTrXdnu+YkTJGMh2mmNeNZBGCCSns
GGkuucHRt1I1KfpruPOD+w==
`protect END_PROTECTED
