`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X/lhQR/ROiXtOJTKPVIWz9P0IU5GCrkKVrWtMJFDX2e3IVYiSh8tdCT7ctJwcFw/
K0YEFMXLZJGCDBAsMGeHn64UlW9ZcNyen+ubjXjoKXfv1dkcq0hn3qZ7+hNBCWhW
jMjLInu9NoPdpOxnOouyZzM7I17R0jvx66FYF4lqrCY4G5gGzRKiQ1/wpzR82JCO
7JktcGpBVnCByC9Zy887MMBET8SqlQchSig8un8pGa7poXy7kZAbve7qD4a8WV15
B9aVHhfggQ9gyebwl3WoECaSLezlK2mMX5vZ+9LtsXlNjDxxcpogBhRhJxdt5q7K
Ml33D0IqBro934z+Cz6d7hPMeZYBSJbnR9F2xKmwNyrKN6gP9zUmhBfqSqKHyDkq
xMmJDUtkEGmr+iLQvDVcuRepDt3O4dQYiiLNkqWExrEre7CUziJ+9YA+rlNSsS6S
hO008cg/cE3OetRCtY9AUD42eBGER9RDwQhX1HgiQZ/pX6ET2LEDePaP+NwEAgRp
Vak94ToQWw4xA3+SbDL3DUPxuuHgbULbxFGokjmZBzO5h8VGsUC0gSWxlVVxUP4a
/DVqD96aAvncm1A8g+wkZ83+wyiO0QgtloPX8WPgz/+IL4CR8/rpUo5XrxI4NwxO
43rdZ+DEdXQVkVJBSKdrQhYGlJ7lgv5KtKa5h0tNRiruNhKAFvt+lmPGSuvhF7tY
msKOg4Piz7DfeMzBCgC0CcEztixuW+iyMJwdEiA9Y1V+RN84+HB2NukjsZB3ioe0
WXypCQp+cjWOBj9r0IEp6+AQqDpgNvHk/nV7IQeELt4BtwPnVfOBRk0/P1Sp6b+A
I20A8B3AyJ9YplASByOeczdH7VdiYLQeVgqnZWCODQdCQyKWKpElX4B1NoIX3r8v
sFImP3aoM9aJ8TqnLesnKlGQluXP+x4T2AIbWOXbOM40pv3+TM+8P95jVvlZf4fS
Diw8/U2DvH4ztqZXDi1aKU3NVCRORO36MCQVuy8Rv1L8Dn0pvF3DmxLWFlLVEWsi
tGBwpxERB+ARtO9E1GIcqEkgC8T+UdC9k5WrOh0ZzwzOACNkiDxGpMB3rj4l9xoZ
aSeZruvkpm2X/jZvCO5imMvYjBF+0TNxJdXrYHvQFJWcJYFwXudqWHkOG470kmO4
6nYkXnWa1NpXmX7eZsO0GpT55E6f1U9C0sYjl4zh5g8zus6EuwPQDTbbxTn5RqJa
V7dgyMU4S0MznE5eLEpwT2k58xHss3RpgeWCGAceuwl07gI+aYu/rkQHWXUgrlqQ
ouypYSKj9uurEvsKPWisBW6wIV3v/Sn1eY2MZZp9SZ9bebmnng9Ps8L7OOENmU1/
2YL/jhTsBW07DqSYJY0tXH9zKYl8O1Ljk/2Yf9J/sg/TRjU/y5g7nxcduZChpGFr
Fnf0rqnIey9iDcxgr8ZRTSAwTVl1CN9s7vMHtjrRSJjZ7vZZsP1lGj23aCXUkzpF
GUPXUNSoBkUP9gJtKrUd14jODAPztqWghv+Acxp+phQBxq1dyd44bEZJ5GYtjLt5
CmW1Y1IRDgiMYci40v2gT0tTh5j8SDJbW0hlosCny22SkWjta3m3MDR+smjVxWU9
kKFiBci0xq/EOg8TcrEI6fXdwZyij2p3QR/KavCl9dm8ZKiV6qo9LdhRpHS2KDU/
tCN3btEWWOWCsmRJfG9dbf2pYDIH3fwKSSHslcgoAnnmQ0U2Ehl0au73799WAO6r
xi/k9GuaV7aOW/6HpC5Mo+BPE0YlxFWCoOQVDr4VYN0kEDhPMQmMUnrmdkGIfXv9
TjEVC2EOx0rCt69/xzN4EmWQpbPRt6N/iWy+wfPfBxj7ZFw210uDs+pa6cNo7Kzv
JLkERjl7vcEPxan5Artsd2Jr2wrEHPoH74lAp5/wT+8AtN/hMBuXC9CLCZIWOF1K
sam6BieDZRSo5DqR3DGBKDzM5/FrOG4JmK16FRhYk3pBiAKUdpq/0ajB9tkkx4GO
Ds9tkcfuzImS83cPj7UdNeN8PmpAe3RRKDJoxjYVOhvo7yKX0Gx8l1dDUDO1DcjO
QqimaO50Qzznto6YjLMsO7ni4qsixaW6+edoM1mDRZFM5X8VekVsiTVan+Rz99AD
e2m64nEJhd38d69HTuoqfPTCAdxo381ZHBTZPspFR6D9orfcTo/GEEDpB7QB7Q3n
b465DBR1pjdabmwrAlH/7L60kXPay8T+xGdsKORtAlTDQjs6qFtNNQYK4oEoGaB1
n3hlctIIv26t1EZvqOudU2w0E/+i86Pq+qpM2t9opYlJ5+MdMckEZy00TigNWB8z
/KOBO+Y5CO0auLXfUpJeaw17FCeJUkXKN7jV0GBQ1hFFrbq/de64CFf3f/s0FPfp
6AmxBN7FCqoKFvNsCL51mD0ZsGCx19s4sATyPvbiY4T+wdJpIAjwv33nBLi8ghzy
3yuo4Th67xnoafMV/ZqNGIskMRseKc5qcT8uJv4N7OIb3bE10JQjKjrsAPTvLWXi
nDPU/PzRZPuD7NpSZ20LbMDPNUjS/EuPKu01yo3SbEJmK11dRf8Xfbwv8vQM/XEz
mKOW7TwkD6Ili2ZximhuhUY+Fkj0fHrZSH/EzsR29cAuB055gxdVAUPhAzc4UlHu
qyuIysayFkRPPInmOZQ4lTh4Oxq1xI/BngW22YQ8itJpWjVID+BtKX8IEAHv+9PY
d6SROautKd8hMpuw85X8V/GMgnkqUN/wnLLp8VUxz2ihHEdhkQ1BwcPhG5H9W/Gi
lm+Guoml7a3UjWW4hiCS+a9au6/N+66WjDxNHx5CPhkEVHgKHV/h8eH4hT3Y1AZj
RM4oJ8+gtde4SU0Dm9sCdbsh4XT4d4hzbuHcl/gQE9vdT+xuJNr0M3+z5kjwMB8C
mANY1naGFC73U4z08gvELjOUZ0IQZEBnkYxCm9q0aOKOygdheB30Z6R8/bhDlNeu
pqM1SmlYTw8hBf5QD27nqHflS4EVAEU0WE0q856ybQRoXcXHVGymJrq1/GI0Bmu2
CG4P+yF2pNgIwWP21R1EFpgDR6wzXWsSvXB0UVMW2UQAea4PzE0nPBb06cjkIwtt
fRq4sFJL0JcS+2MWVs5Rm/JuoGMSoG1h3T4razFozcuwgFRunLHrps5Z33g+SFfx
bJ4HRX8IXMDzMWzef1BGNhZyPZ67m8b8sCObgMPLvbWHCKxQmY9y95bZuOIVy3gv
OYjvbfBdo6snY+hLfdcI+ZXqsYbxMTjoIuX8IsOduUs/RY84zVg65rp91lImnQJy
WUIHsr4AqUkggooRifRhh3I4ln5p2VdihipyVnxIMsy01Qmmy6/SFV5WjgWWT+Gu
MDnw03XbL6IsD6d84bQdD2Nh1Xb21VwtaVL+H2cD1x6M/7OGk/KgPmcSz8LMnKGb
VY97vbM7oRqXaBUfRlDnrvVimZEU8ms6LfvOWaSvZpXzdRXscbUjgdx670AjeLQ1
r7M2hQE8pvXbispTrHnpAH/IjYKc1wF9qhIBe2VlUvAakyJ1lB32T0cxMnMEQOja
wLDfpfdRycLJ0DB4Z5BHrTL5PtUwQtoKQ82omTQNDCwqDO8zyVD81JuPpRkjVYob
ugzDKvp+jjbwcYZAalLupE6TbbXUxjFqnF98UtS9Zx1XCmFv8ALJW26qPby9/Ywb
rPTX/i+aMlg4dQlETtMiCHWCpMqpg2vpSktUWZWwyMjhixnJx1GzMvVJJI1H58/5
cSpeMQvg+31ru/c8wWMKn1SEndc/Z+nz1A7z4+id1yV4NpezxDAQ6oyoPj2sUKg4
ZIOV5VyBFC3CmA8Auxi7p3AvwsIga6cx0PMqM67OKKRbbD4doeAoTQYPc+cCccBo
009AdGqN2gssPDAvvHKB/HHfXiCmBZyqzRnqJovXKvpFOk5+dh6iAGxuww8qIEQb
vIGUbh3Bf2Mi4Zirt+oIYbm5tZ9GO7dfUSn58Y/EXl+tRsjUdXTWHONNZNZZhQp3
ViLRDPt5hbonHYwOhy9Roc9biFlswl+mJoOe/cmkabLRiivg6Bf0KkJAGlkHQAjr
WtAmuPs8/fsLh3d4IaaKBvT3JSzmPJg1c+l6H4HkFg9Ivb0CfBLGW+wKO/YIX31m
suYwUx7yJ5O9zUyE5tUTsGTPhokJFa4283gYakFfZbsa7EFPJpVc54nAsN1MndUw
LFHZG201JtI4nBQqcaXCqCW8p9qsv7G4PS7GwcCFVYMXwHvjliDoDPmgs+s00bd7
+6QTfGv/eIZHpDTapPKt/qHW7y+XcLz56lXDQcJg7Hmt/dQGg3B6Z3o7bnnHSnD6
PzlXwvmdxtD7E8Or4MPVlx5tj7CwNYwexNWp04rsDtaRhLZUyUoygIU2G/6xzhkK
1SnLMMM/pY9OiFW/AODKJ8z0sjPNWksmi2PDpa7dwv6VU3l6g6pS3ohl8lHHXceP
dmTVmkH0/OCSzwSUkdAzPX6k1SIFd1Ui/wI1uZ3c1CsT1o3dogGeQBbX0gVKolVt
W2ou4aa3hsyiRn0xCQx9An7aqna2jQ/T5Ad/oezzIt9DBDrIi3TEltwlqDSKXe62
XDkfwHq5rgfJfWwC3A0cSbNw75QDz8SbFd1F1m7w8FrLUEx9l8XHxMuB0w/a4amh
L1NaPGlVZF8JxYYLiVYoCORM/vcFobuWR0vUM4+OLDW4+UcPmFnsjkEAjDUW7jJs
rIYRwjV/XNWm6YhduV5L+3rhwSJHeNSacpPhkze/+YhF0UhDcQLr6EATsjZhOKuq
ERzIhqBKgedWMIbTkYMNgYWk8LGU1W4Zu/HoO0Eewa2ebpLL1/3U+8g8Nfi89FcA
FXqzn/yNXhubrAc21sLFOVw9yzXeSF+OoHYbrjVPfVmAO1N+KfIYq6q32zVuQLi3
Y1JCr2D00bSIc2ysogsQTEBl+2VuyHJKefx3AaKt7Oc2Tb3k5Doa4VLoB4fKTDM/
AREcQSmMes15E0MNF26f6MLBoApYDRVXXhj6/cm1NH5ST+p+JYfs+XNxqDfkwhHU
RGxYuXg8Pbkxt1HLi4QQjrHad4xQ6IhFCZoe6eIpH7SkunM3C/reZaek4QyeaGtK
HFWo+GQfiS7A0XIbNw3b3+UM9xGqA3XFzAhngCNB4oXtMSmolB5nuBL/0A0Dwrq9
R9mq6+JPPPjxiDLQ3j8UbWSWT8AXozyyzUNSX5WwdGvxb1a2NvPlFuSnz7jtL5o3
Dztft+6Obez4Lmn+OPO2l5Y2Tzl79HX5pKoL/svZIdozWlFKZOhlccYndrTyByRT
Unpa8q74rcVcESH2O6q2popz5KsYNoydEDLPPLobmo6PELp3u2U337mhfA4HMP4M
gEYh1v39/WHMLcSoNQ9EZ4d3Od71xG9ES6NeJm275YoZRFHEGAC1fQMH0yaqb0w3
SyMfcaRfiG3HYsQl3o/4w0ZmKPXleV008KyW17Rd5x23m27SH7iLn2QZuOaI/huB
9alugFdbqgHfAwtT2zbgCjQNmaqkHlOBPEFF9cVUmg73x0jYaixcuuh9qn3Gz6vy
WpAf/DUKw8BXLQKYYcOsGtABsn9d9tHSOygxOqryAosZsXL2UpMhsAiHcpQhQ868
DQQq2DSrCcQt7uEILBcknOL5ybFtEHcKBL2Ui4bcwz77lgWDr5VnDrFNHPebjoq2
eoL6shUWpyXo/92mM19C87hP0pID8fWbNoeG9jJznkUjR1hrfm5XjJGDvFMnPno4
+SN6s7Y0V69zhjk5CQlISz/5lVoSEwY16TvGOO8nVldva9g6Jl96XEBSjTKveZtT
xvxcaAz9LrN4tU46PAm9rKDKa4ROt/K5aRK9urn/mJbx1zLklvVfTYWZWQ36pMFG
TH6ivGkSqFSgAjCZUwYmmpM4j21IAdgZBcxPbkPl6DL6V/h8rYFel541TBk+K+Cu
t2KRGPwT7ZVSnR/1i6Uj/xZOdFpO/4htXQoWsYWQesEXkemjAAttUu2GB/Y8Q+IR
t+V4RIo9OZ/RuNS07/KBCmRaYqFKxmvOv6Iy6awjFGg3azRQgF0kn14LAT08787s
i7fO6mFBA5i5fFCADKxUleDu523epnoShDkARA22F/+rf008h4s9+F52sVbFnONF
0D2Q+/E+yMGsOQgVRU5pdGi+PnGerXum9WfhOdxECqC7rA3BM6bO073GEJPKxeIv
oQbcVcSGwq63blX/by4ovRuvt682f9Y971HBdkWpPJ4SoYr5CYFKy6iRiyFyBhfX
hub+Vj66LS0jVEBVHWmIt32c/Cv/sebpFFSofqbIcNQI3MCRECwSvOpfSfcoSo3s
5jTkEh2bYz7yiw3KIMp8ZSnOEQ+dOUSMBGVPY49zJ0w7QRAR6fEX20VcuQIWrxmK
EyZ6ddwjq9c5qfKiaTel/azYrbLL93TmsevNOb2WB00coBdyWCre/jyABdGYCuOh
GeE5DDDjI3HXApEe806BQV0DLcoZNKr5aAEAyKEtuquQgOkFdMvOUXh5MlD0gDs5
oVIgvVnRqL9XH/2AAhZQWvMV+ejrOdYqYuE/dGfyH/SSx1T6fymaOKBzjiIYNO8l
7Hw2Qm6xwFq2BOunslMhpYyxt4UpjgQIVp4rhuQxgyWsc8MQK4kTpjp/Cq3pQT/g
I+nSAkIsPgeG/JEXbWT2zFvbMCsGIbCLJ6gNoLKwCQf9WB1mJmarsXhREEo1ulqd
c2RC/0beB8oy8aKotpjTvcF5RTEW3igFFvprbCFvWPc1c61nUct0AkCMDJ0+g4Kv
by4NRRCrK916Xv+8to9xc/YIAKaayexQlp3TP/Iv5gOkyFmUsvXiAIVHkVcPYgK6
URy4re2/glbjxSXkuQ2wG4tVxWt/RW5+4lwZhsvPk6sy5QuPyyrmPHDL9d8Jf9tF
ncptIBNLR1ooNZmyA6MhO7S22tRnTOguVUih09v6D8NrF7/8XUF9ewq2AC0N5wkb
urMjmjgkH6pBMA2g+mpjAca+jyEI/uOjbmoerahNvZMupd2uXmo9JW30eZBteAIF
dBkSQon8DrUlGL3SXQWAcdcnekfDShUdDaOcfFZ0DkPF0USwWHYTBISvPKGtk/CG
CGfjE0Ln5vZC6slQ9AqTZttWtqtyhbRTLKBVyYkGwbCH7eoSv4rswGxnHysqllAh
Q8j1qzGYzBXSyjPj1ppoq9Xq7Plnc5llgNFRo3GOFH4oY6PIEAoDK7CVa4wJu8Zp
QdnlIEHafhBY+/V5jTXX/nz+7A/5qLH8otaMFUbhNiAgFt7MMH/f44lbzC5RFSxC
wdADnKgTKIpIKLQH/fsvnMoZYQNNJ9AVSl+PgbLODYfkws2ZSrzUadvlj7ZKrMQe
PhBsUE0sDAH8dgj+3ptCc0Y/6Mfm7lI+ajBx/ItyXdGkD74xJ5WBA5dVA8IBIAq5
FpILBTZYSAxlHlKjxkDlJxtxZRAUYk1Mfw6strhJ7ANOmEyrV+9lOjpg0fhevrtU
lT+tLCF+oezWLI5Pkow5pLaOLgN9SrWKsPupa23nyladkmC96m7Tyri1/BJ703rB
WluHw5C67/gzX+yFW5aRkp+mhk2FowBN6xLD7hrm1u5Mbb4ap0fet76bGN123oNU
p6qpJMLVnEfLrkCKNjLgNUCeMEtz8aCf2Hu4cr0XR/yaxz6G+x8FSR1wbVcL3ZA4
s7ZHuuO/f4w7RHDiYtJoWKNeACzT9eO3upQvOnXPGso8DQg1GYB2oME5ePpbwwSC
iG3xeEhKFrWdSlyudits7O5GGZB2d+8hDUnETIRqN9JYcElzvGEzdLl9mUhA6iwc
VP0upN5nncgkwTspOiH4yUROWu8riJXo/DWKiuCW8JC8SeZ8oKYf4smeO6Rin6Ln
QUq/iGFVii3xBhprwdYgdev7N50ywwwEwjGaFEMxQYfQ8TVb3Wr81wAjApaelakz
QYHb4+qXHVDjW6cIMfNbpE9m1ZY+dJ/v5eQEJIu5ifcJtt7wZbWD2R2t5PdZ0GE+
7kbnkyXDV2VTiDQAWvUdOPqz7JyykKECyllwcbnt7TN0Vi+kLDuS+UcB1/X8JFdL
vXUq6ruHMyvN42gsYd9nrcDZslhKBBwZOaZiH+wEPr5U+Vn8YNtArkWA7/O8cq/K
Vbt16NC61Wdr/kkZmzNN6BqhCZhleUyNH2vqRZrv8d38OqWgGRgjSyTQyaz3oedv
5e0UYy0lwgjoryrFmshn0543PNuayLuT8DrAus8X/UWyYsqCYtu4sjBgTBwYll+G
2bBFAI3vLRlAsvCxShRltn4GfUmN7KfyLXpgtprzPrfzlAn4kwKCYOPj9Qsh0hS9
AGSG9IcyllSvbcRTHI2IeC3Y+knv/HLcSz3Kkx4MS4jaDYDd9IuqqFE817ja+6CU
da1YFPFlvM525v3J9ebHsnSNub7THDNBIGpM9h0zTBHu/jCyOTxWBQwUlJGfP0nA
537WDPFf3nn2ts0pGEwEw6W/d4hHaJwc7Dxmq0mZPmBz1fLHRXvCHgyJu51qfZQF
+0dGnBIubwJljjV1p8rqiSRJORnnMr7ijBRfRBjfmOXu+mTaKTiN9N3Cl/MKuyeH
kAuIWvAnwBTjOKYortCkhDPs8d1BKZw0gr91WTyD74xiBKpHl95jwNiljLd07/EN
f+wcPz1RU393ZXtCPuvSRL+isq3CcbqfZ1d6LtLgNNsf2vsQHMnUblUWy8JjxVdD
fks6Fr3XjH3YxHHrGtPTdWi0RYCqBuiKTsa+KY3Un6QCriVCKxOGknjCyeZ7kTze
WpALgg7liBV4ySiKyKUm0NxZPP2pVaGzyoshfyItaRFY84la2hik4n+hy1twO5GO
xLnREVlAx+aLbVDL8iGxqHvcYU3fvzAHxPOM8XJKbnFP8tUj23dk7x+FZfZdjA8Q
OPn6pfeOFUEWRyVxYuXPsrNGpyGnGq8ixJuttuGPwNj696gvQvv5Y+ceWdHEjyEb
SG92jtdZj/dvydQrOFgfMSCorhuqjXP8vMIRVECej08o2yug8TMagCtKTeRC0w62
y76f8lWAimbRrDXR/7Hci5HHkoACUOrrSRzoFLysDi7m5wJpkvngmpvDlXWp03yR
rjHgNQZOl3NKrNsDjUu++njdna/PLhNJCJ7sFF/hTaX1S/OF8RZcVllZ2m8KTucG
89zeuElMRWOtt0nNS8EhBykFcWNNZfqdPwIZJ4UhUfbCqBrn5par9mUCV3bKzIoF
cvAmopjkVOL79qDktKiHKld9dMI5+qRGorY9z8w72kOyrCh8m89MT85M7of4SzFw
u61jnxbeGj2ydb0py49JbhIMwd4Ta+itYWpikMKr8bmSSsGrrYMfNdwHnXYHhC9q
jUFBB4UC0iUvjzLlG4765zzpPNXm7BSeZxjjxrjyiAq4DC/tbIsGexiaLpbOnrNA
GoDnztANJ0N8uivhH+i3Tzsy+Ht8zpuvTjwKJ+0npxFu+sUWuiByCO0s1CMaV5eY
P08vCooBudy+LIZngNgZO9Tw3vw6ba9SP3D5RwdcV5OWBC9fTxiIFCxc+L5wvDzw
DeSZNKkDTIeRpUktgiscYOlW1+qKfA0La24ilrgUXsx+iNtCtwi/to0rtC5ZSdn5
M4GUm0Q6i9vAX1UJiFOMDivGWQdvZq8aCazPOnZo2+52Mz2NANMooDAqtfbAKUC2
Xix6edzsPbzBj+PLUp8J9tkGPwY+Sslz6+1vD0aDAvIiKeaxrsKH0MQR7MopP2g8
CsarPLjan0EcRHu6y8a1N2hpR36zP9fOQdLCUS/ZEW8u/3pJaUkdl48s3x8iPEAH
u6RHGbHXIor98bldeKqfUaVLU9IRTTaPcyEqdY9RrWo1Mo4QeLSakN8luQiVSi5M
QWj578hIlhEGV6Wtnjc2wKKrY0EuIzV48gZsNdqxFxeqlNd9o6q6Ub++FXb7fdwn
KLoMvDsyk7qDeEn/wh4DfEQ7Na4UN6UaJOlR6wgkaURT1cUgXJfGi3tF7bGV2TK/
0XnmKs3EyHaxxGFGUOHrqk+58w79GsNOU/Xhw1u3okfY9Emkzs2+IORFtQhDI+PA
QNcOCpb47S/1HSTQpmWgH6E2hpAo9j+a24NMcKBlp8mIpgatGknlBDEjB1PypeRX
uc8ZuXpRC89YakicxuS2UCuvIL0NX5fYqBBkHoUKgQzKXgevUy33f0wHF3QF4Z1r
ISL0sq/pXSZtt429NS+P8FCyxmGVBRzhE64dhkNSBcXTj5sFfVgxkp7l/k+4Xjr2
Vsd63y3zM/DciRqRoCwtq4k/wGvW35O1InPJT+eBJTNs1N4CPSpzByVsx/Dhs6yI
qvkmWbIweOhOWJNbbUO88sYTfV3qTUdxWPLICe5hx7M1bFGZoSn9IpalOOQs/elk
DYplzi9MKmp81VdM21JnxcCoGeHFfofqjzONBNbCmizXSEIcR8Szs5Nxg58P7jFv
L6SDhyZ8d+2UDZW/08RjOgI+sjDvpLknUyjx64GPQbU6UiIg12Zw7KsiCjLpm9jl
wfwkGOgLA+xsW4EVCcnB5Em1E39HMEdf+6gzlMo1Olk4kHzCkRMKRlpdZN3zz4yS
gWgsi5Ma//eFLDq8FA6ZNZMg/GFh3YW3CtmLpbLT9sivhX+sfzJH6PXkA8coYupo
kSvHCdKg/vz6G7qjfFMEayrifvN4pkSubcwkb55RfRzJsPEiM57y69dNW5m8BgYg
6jfaIKwK/3qrgatVdCadzfvpaedKBNmBtbhsok+TtLlowwIcSBFWbjvTAjOxDl5p
pozbS5CEgHKwZkIDJCW2wDu2mrirCvyQcwXeyjphLcW6bsTDPhesyZIHeVqZixRz
eOruZWSufG1xU8joce8UjKt9WZ/5QfjxltHgEoUTA9jG7pSSLXhF0Sz9c+z+IkqC
VRGtbzOk8K3cHJjXiSMGXhdtLS7XxJDmR6fqzslJYeuI/0+1ImKCRrpgcAtDJeyf
DzgJBCDHozy4B3zNt/p84Fcn/OLp7Oi5QNu9BBQv3XNGuu7TEk0NTuH4nx9SOoP0
h8Fz1xQS8w3bt0YOTm5MXek9rqE/NFObV2a1ImYKFVVA4MWmHeb8AbMlKrQADXqG
1BkAZt/lq+CfiUGbJcWTpQUVh5mWwDEfLiHZBs3wmwBgui1mYp6sEHmGejXC906j
6bjo4WPSP16t7XetZqqWTpWtG3Q2TnF/lYhUwxUwQzUHLvqkJNhiNVnMHIdCsv0F
rILIU2Uiw5U25VhrCYOobqzSWfYFqI+PQdW3eoFdNXahOJZc1x5BpmpP6dIEOqrd
QF3NEFsSpefRw0uZY1+7JGHjFKkFtPgB0SiwuQM1BBQiC3GVqi4YDZouuyQ2BgUr
iQBc3zgu2bXzDwixx9Lh7dk+pmFjeaKWvgUz5aOD0QVQHZWptF8eY08CyIQC3EI8
O/H/agXAoQ+uuXNeH191/Umj1XR8sCxlN1Q9F+ah9RZ48SNwQFmQfFFZ3Tmze8h5
6s2mH7T1dH7OH6WnpuWmlMrSfgCR1uRe36Bd6UMxhcgm81uFb+cFZs7qXt5RRC6r
fD8rG0I5o9/UOYPvTvEvZFTHgL0XnbhiKHBZc+qdWTAghynJokdD2OrmLwgs/ClC
3OCZpowRA8jEf5EOKsm/octXUIKrpFR4DVGj5STdXTsYVsErLv8GbL4R/BTiJkT2
Vsux6KfO17I3vcubPhxLXpX3HtyY1JSXxSvI4q/armN+eKMCDbYJrDlxOZ11x9Wu
xBc722iajZizMBm/fDj0MXsXFwiBPaEtnpKRy7B5VATRaRm19iwSK/D5gZ9bPlHR
jXVWMJ5p8n3kn2ZcSbLVP2c+1i33MvOm1LmjJ32f0JFuvokxGZeMtCdWpsSlnREv
3NGzckkdS0FFCWAsKzK3OAvU78pemff7ccES2JVKq3q3zpi5dow7Rb3FOXzZYIFK
iHUAr6T1t3HjS+JtVKrk9AUJ8Apqm48Q7P4Vc+QoqBiuEJh4l1DtykMLCzWMy6dI
AGaoE4MTUxXZkIgAEirqCFAOPug952/Mf+SWFXA0dHoydPAljwF0gmH9vXgExjDj
UqDpXAU9GWvwRs76CvXA4uADeagGNmnLPUICpDbZ3Ehy9gooOY0q1kdE7Kl5pM3E
P+zWPnvmWlYUtKREaY6P9dDGR7CyIRb00F5uLiuJqcKjdXEUPX782Pgt6VfW8Lgf
sQBvmbzo/IWduWxv1X5IKzH25TONWpS3IKk9uB3+h0I1YgDvCNlbI8IcJ+KBMd8O
0ijZfxKsY7sUYZMpUQWyftFgx+T12+L3ufatJqwc4LR4NTbybhWksvkGwmEkAZf+
Dhsqrbzo9KxdYpA4IaUB98/Zv5XDY+mU54Mj4p1IQYzXr9G1fesPpax+Up4VTxlX
9VijVxXZCIKqUiRQ4bh09evlQzkmiPPB4kH2fAg3r3rehXVA6xE3c1NucsmBzkTE
oMkkmYpNPWChtnZHOjM3QI4AhuwxOD+QN5vcn+hbZcBEM0GH9m501FXbtjL6eKIS
MZeQvm5NJxBbkDY/vFKXIYuzk0AT+ypTdtSIPIjzxSOTTVez/08JcftA4UNZ8O7T
jOVmsKNLvoUMq6bX4ap4CHEFEbcPvSHTCndoD6AyZwDSfSwr4PLhu0A8DXgPyxPm
Jebh4188Crs0BYjLUz3x4GFCvWUHE0WLoYhnNvuYclm/BDYky9YczJ3OXc0iYDWb
yPs9Yg+zzB/Au9yLj1TBmQE23IvUBJwMLwYUBVGBOmOokMLAoftc8rC5Q4qCDdac
xPuN6PKAriYDSwgH8oJo0G6k7esEmUVNRv7I0YkcSxwMyN7kQbI9nCfVxBQFH/ll
R+Fx3TKnfW6mf602lT8f2m9uURDPQUf7GuRIP0/0/rF8I8U+w6ux8okdyI1yW4ko
zHddWINAqM2IjZdGtF7+Bihu0KDUA4ZY780wH43HRYGL0qC4r+VAor7rXDfVgt2n
xYnFwd7ExkAjgwGS+V9Y7d6FIwcB0elrojdNHO6puMaMfmvUZaj3SxVIKQKX/6Sg
BoynX1js+pLWyLj9AxDGBy215yk6LMAIsEsN/NjMkyhsOvZkYna2l9pdyfWR4pBE
4wDgDbtcsuiviZjJXUcA9zdw+7mMOm0PDd3h9RXd2euI2qs1dVQiEqqYQKnRMR8R
vEiwKS9VLoMy7+PMCgcTQWK1ftsg1VnDGD2K6Zl+w0yPCXntEdgDO/SoK/V97wUp
4McFnaqqZ0nDbO68TukAiA4E0RhzUOn/odH2mVIA+Mh3/k5I2B+wFAbFhfAJB4pW
tpiHd5eHDRTdxbBnrxuaO3v9p0Hb62ypK29QVz3njZhC+K3G928Zl3Nz2S+QHdjk
eLIVHxvPprD6lzcrJRhD9RQ8UJ5bXfjA2FBHFu6EjIiqofgawUCpb10KqLS6Vakf
Wf7AkZo6NLcyk/lh+5eaCklTsnMYJBHYH+0cajS7lftkwTl9ndOX5LhL6oYZRGSo
SD9yGu8gIUB/jmEpNpNQrrOYf0My3eVQ9xF5WSujDl0V1bnsJauQAqmE/qZjkEtZ
VtFQwduLsKTjF7Yaz8yd/KDV1hOZhgE8pH6e28R3Ur4/h8VYfZq3PUy0JFeVAbAT
yWwm/i4d67rXgAXNl71M02Hnif9pOW8TxtngEHnMkqf3H5VOL+cxg5rW9gKNOxh8
LnZnw/8l9mKMg3XhXJq5TLMbtK9iEZeD/iwxCGmzfsYxEl/vBd30OoiAU6RWwk5W
VO4MN9D7gjJushaKpnFAQdrxidQsP2gg9zSjVARuTSZ8WNnqg6Z3GITP7lp3eLu9
/0ogUlah60Fw69oonQ/N4Fc7Bk11BWWIfIMol5kg8zKNQufnrNyMUOUu9gDDPKIW
JfYLhBdCvQiv22WpvBJMoiO91LZyZqige4un2A1RSNK/AU20vXWNFRODyyOm5r8l
cK9WFzJeM1VxhIrVG27ZWEgzr7lRQxpHjNYjzlyObgOmn808BMcNiqSCcfzPe0ty
hJ8YxpRJpJ+qPk9aB5kzALs3G5j3yuWQfei0xr+L91FvaIhz/q6TvPTci55n+KEy
8pUN2onguBFD56q4tkeh2QFZoNep4tjiPeWPAcaju2QjZDTaB9FPj0TsvPO8w9id
ghQsoyLdE3CpvT7U6ht+gbqq6WwNQgFwutYWrtcIiAH1MsQ0jaHvoPlXLM8korfj
TFwbMoOIxg8V/dygNJWauGGwDtDa0JAoXdoRrG1YW873Szv30O558llXBxsDMgFt
MGp/4Ncyt0f/44evIxyb6LiaH+Z+bQzC23cPIcP6fgyAQoPD2RjxlGeTAUTmjVkq
fKFzSMix7h3x/4o3ZINyBFsfXUwCybuVWkRBPsTsE1qH1y241gw6ZcQFPu5C8ktu
jE4mZrz9j44Zrfo6tRnar7SLSCMCug4d9LHeGOm74WYVVC7sYynp3eXS35mVRLXX
xsfdlnakb93uB3xzVlpytmlv9mVmEhE0fdNjM/vMlOV03ThMjKu0KrnYqchS/EdU
WJLSc+ezE4jEnAe2vIjzWujAusPSx5slOblxkpWAZc0pRt11FQKH2wVgmmUKoyCC
8tg3IqVWytBEeEIaQ2CWdw1ev7p9PxzA7ECxhBjeeqeNbD0pg0yFRTXO6OLzgtM1
SZRf24AZLPH3zek4OncWBk9H1mDUnfqi/UsVu/5kzgFKgucPoMeBoIx8FcMb4c0r
c6VRFCjHidfZVbaNtbXaL9gF/TpNnKpzfIphxlEL5IGe6mh26+3wRuBLoVrbM8lr
LF+AhqkV769a/H8NGk8fZY6j5hUY6hE89JXPZtbQEszBKxiPZLexczfPFW2O1hNs
qIkuI6bUhY/t9jP+ITJ4CY4y/m+KSsBfhq43NancDPB8i+3w+r3gncRQ2HldjoMl
OOAIrFur37mjkZnNfS2wSJBdzjZl4fn2VlBrbLElcvKsGozEfL+sQKrzmsppaGnL
YQlsTVNITu5sAqDBqR5R593f5+zrciYpvGO+3FG+Yyf0e06SXOun5MIjcuIXTVB/
WK8fxA2rFHkdZxRR9f6aUNfWB7cdlnOcsxAS2STlqZeSEugMpDFHOrK307vd9EzL
20LwaDQQdm5+j7UTq6pYiab9VEm5RVvHwqUSJbIHUrjbjJzpTQW9N8wkgu+RTXlf
gEP/5QfhCGUhejkx4SS6BGdK3Si1yv8S0dHPXrW1YimrB+Fl1tNja+aVw/+doV3M
+MuT+bo8Is+WrDoHVLM8IltNFLlyKOgDTySiBsfACr5OE76cucRhL0sHM8WrzRVU
be3ptah2yv5mHUSAxaBjSmT4o8d4eM+5LJHjK2w2pzuVgNT3mQFgStnz6FACZ6/Y
HImHPbjuMpjllHfj8uQ+va9pgoAHZWGDExhH0cSowUTmDSJVmmHy7DnsxunYn5yd
i4a6zOKggbG8nEX56QkqF7QWwqfTdHaCP6ibgWB290JSzk9ldXihOyRrcS/paWPK
re+7kv4GdyJOmnAiaiq4cBg/nlDn/bByOa58LdqUaWUm2NwxLoIgMVCBm1+NhI3v
YFKvUaytJj71CgMhP1uK5q5Kg5T5uWNIrHhFFiF5CpN+tEh5r/tW1ogzF5zQVhfG
ybtn+wbDWU1x2eof2DeWREq07es/iwYYKC8dBn+KcTKxAfIpiVxP2hPssHTWH7ao
SGJml6ofgXDwdQ/1ULP5/E1LdNwr+P/IAI8awpgi2K0Kctex8PCO7KW+mtLZJTq4
j6kD0AlaMrx4wNGr+9HMldBTE6MVaL/MIfD6LLRoFjiQcXT7gtV94dVlIG13qOSS
9UeAkUEyNSycNLv3POq7siLLRuJaGiL/tY8wvw8N+gP6nzzoa0xxskwoMaalNp0t
D4sJO9xKBp5kzjqiZoCIXCtVoBIxMore5GjwEjX+IevtGst0gDWFLsli5f4Cv3mP
fUrvCp4aKeI/PMXL4UdS6T9iyYR0Ql8QWBk+DUWNeUScZLxL0LQ44QzXAkZeawv4
pFvYeyx16fskHEQ/3AZFRF8sRcGHIJtiIwocTrKAskpEWDPWey+/1kiq0xPhslQ9
yBuML1bD33ngUpvS+R13BsZUbQUaG8GXJdOuaY3rBcNzZhpZLRJ2ayYwXdEko2rL
zcYOUs48gaHpnGZVGYeHQvirqjUN5Kb9HG74zslq1URtZBlHCa5DOR4pYmKKr5zK
apht3ImcQ57eCTuh4vdck6NN5XxkpG9EgujvbehVUz/t9c5HCWbS5ZlwrWOoaTW+
Ho+yVuJ7sc+FiW76wg66Qg3K5PhqLraQvtxtVmvWf4sR0jbLmGDTu/ktJ2op2GdT
DOCwcx15po+qnnHigvwkIFZP8Tc6hqqAqSZN1QUNpVqZbYnoV5cXL6bcuys/Lpmg
UnfggJhw0FWTGJKeo8zIRW14QgiIASDn+5qSeBdLskIwiHCMGKA2crIJZrp4P5sV
P8gzW6Hqc51+ERM4MHRizseL0IKXbpqxDWKYpwUK7TWKvg6X++Jx1qDqKDpY1adx
+qGvX1K5G19n5MoMmVjOnY8JKv0JFup3xmmaRxR8vNnf+/LZO3pjhrV9vGScxX2C
PBit+sx2svntAxXwL8VWM/1fZkShZdQrWhITbxQyAKO3zkJUrWGrKBlC9Mft589D
moLuK3whq0T/ooLdSfbrpbFaki29/bV6IcKWgMmpGGC9nrQ2LKybNZqJ4W4AiLQ9
wriHuYZePzWYi+TErelhSt/IyAZWaK82EbL37mPozAk8z3ZAyCpgfDbjcpH1C7PC
szto3OZaykoQRZfrZeeFZEbT2h/7UqV0+1uHFmAQXDl1qhrqdZyPKEdKZ5M8NfZ6
ZKiiePrHmfJMnut/C26QxfZnlAqFYHLAUXT8JHGpYYhid9pATwjliU7JLkdnaIrK
0wV9trXBmBlyY5/ouiXZBNG/s1txdJx9r9+IW1P9HY1zWaobxyMxETQmq/wxGzli
esOdXjqxX/Ltk5yzhoZ4VswmuCK4PZwXTYUxtEXtYf7xetmqjHBA/yXmY773GQMy
bbuFUTzEGc9MblDgmkPVGliPJhLnUHZlwVAPvfM8J2lYlo7sT8Oxw1X2UlSEHEXb
cq0eWwM+m2SSd//+dbqMoN7VMjdsuvFP0Dg54brUsDvAC7XN+eb0NJQSZUjipIsB
xpcnk057iX91nFZ5IB7tBgUdZa7iMjC9p6z3Kd7ZCO0I8kUev6X7w/LZSbi9BHBg
v7NFJf9XFqnkVRHkQJm9EzwDFY/TNSglg8cHvkFOAxCPvO3QesyjvwR3Qtqx97wj
M7xvKCvbcdQUdYS7E6ZrUtoZpSjdz2YWuUVRBHPVNl2hkha6NrHIrnMJ1w70+arr
sxrS+LJe1gYlUuwjJsVB1vGEHFCYD/LW19Fz3iplU8apYL3v/hMyWvprhxh2tcKC
a5wppRnzjiwqPVu5OKKZuuVux9UgDR5rqB+hWYk8VJn/Fk3UgzOu1/GA2PiZ3LTt
lXA9WbJCoWrIejO3tjX/tBjq718DikCShKpZcwd36GAMft/nOFISZioGH+jUvmUB
JMjs0efLtUJYyho+dONqeZsVIu/92VoCgciMed6FcalKrpDG5PYJ+gxILj/4RakJ
PgfwN6mlJ09kx4JxAeXOnlxBR3AME0i+NWJOprwg1L0arTcoe8vY34v3SmgDhuhb
ExWpLocs+4UvgoN6Gm971nnp2qfnrnrv93n2pBYX/84N747ZxaElBN+8JIW95VKG
a5bpq2azYI8TIcRYt6OBLkz8mhAqw2MyPxHLYUAJnBXJivBbr2njRQckanAVC3CS
FSObnpursnBU7VuZ8jgmV9Oc5oR1yrPTYRQYZX985cJebbCs3rMpk0PEraO1ssDD
dlYarJSOegdPpWyrvXnHgaMDddJmVVzX2mcpRr4MkXRTAhqzra6ieaIjpskYN7St
jOmmni0XvanAxYSjjp55sLiCSKgPMr7da8pxwnxwRcbV/+mtljwgaMmLNoyNOpRH
hLAXzwUbyfrVZfbzBEHGPniJK8yqtd82/gy7lnvhqEK5zXyAbGUgicOPagpT8fQN
aUVyFhH+5+YCGxk+drOuLn5yfidFzfuvoaAUMIVHl6Dwb/pWuOf3LFLtI4YrxdsJ
IC3BaxUAWTfdEF9rZ9pRSiqfK67AzrKeTDIzKylbBE0NnJk9eikwMYHQ+m+EhQkY
Naf51VE28f9ogx/NJj3a9BKkuf1MomXchyictXzKgPiADACj+BLgQ32KPCZaabFs
Bh77/9hMUt7npvq0du+KlK2qQ3x0rHTntMsO/Md5eLUgykLFEUkUginPQdr+PRlh
uPhoQlQnmxl9mzUamlqWPxq3/yDF7wmMwIgqrbbxAAW8ZIYUrro0HOYxcT3R59Vb
lDiszak3urg/aNzroFKbc5J6XTfq9dk7LnUwHVq0nT7lFJg+Ewny/mhQE3wiw++W
Ao1zaUALq294aLkdEtGJcX7T8KsR2D6N7OGtWDC7aTnAAd8DK26YR7WbJsPnA5bW
30u1EoJbNKaGsnu1G+U2+dRysVObGFN8MRcstjDKx17pBWVwVoB+sSdZ/BLW6z5z
tJ8yOpiBpR7/juEHxYBgfs6m5Vmdcl5X2X+E7XqgMkxX3MVUWOdDL825QoTZ0FKR
mgQh5T4/9ki6jbNezbraHVIaQtRg2r9Q0tz9s/wYB0cq847G9fvAiG+Jdazo/Ad/
W+UQippZK1hr/lPxrz0E6hTi/4S7XxertusE4zwkRfpCXdLTJKSfV/YCd1DnTaVa
ZZY5GH+wTdrStd8sfIU1r5vV3FmrDfvmaN0zpBVxwfKl4r8aBq/UXUEOl+yJcete
VpzNxQXcUGIHQ5lhy2aFcU57VB66ANWO5t1cqXU0G4iyzyj1AosejEuTmltkliAQ
ln8yCzlVHQnOwPfOwSjCtucMxOppd3sSxI/HBBxTAal+fgMP7NjYyd8pl9QmRVcY
SehE6Trzr7q9UooYlM9ZY3aNx3iPXmyNpmrSWLeTFNJXgBXudjOnvUqeC2Zrehdq
Jhdn1qepDwQkkSdV3yn2aBFD27l+EXqY7CXeIiK5AhMOnYMg9OANxwwTPBmSfFLK
JhJzHYro1wEXE5wMysnIBtBF1vhUop2AhE93LuGwFCEJe6rmGFSZlFvROXgQ94Js
IQPpwxtsbUWuWIf9inHh4l0KrpI1DyJmbDUV6SxABJkq184/3Jw2bQlwklRHMVGn
V3XG05vzKHzechop8bU6goT1urNuk1RykNNPiW+tDt8vtUkZps/2A9VA/zLoN7ib
Mco7C7VK/omFN3H7Y3tasxSMJOp2wit1fVRXrGnhcJy2tV+A9BKj/iz9yYCG47GN
aii5vtSfsIezHSBrZJKWEButq8D2t0eq5oaWaXR8wUVeoz1PHuK2pSAVqAsidrKt
YeE/eCmBiA2O3n1SrVwL3NBbr+3GqqGyp4af5CIu81Sr41Zq17upTA4hRfBDkgBl
X5GMvXTYK7EJyMaHSOZhSvfQsti0j00TwItURN5lU73K4H06z+fKKCabF/mWTual
vsnNeLSCb2oeG+oqK8lMRGLELc6jiC6VjMxVW9Tifl6qwgNjaJftv5tiFmmscJCx
rlY8pqwDG9gA00zobHpJ796p9nduQdMU82xrGCRlT8htNKrU5ranEVrblKNDJ2zV
RX1nm8WF6RQOQnNyLOUTUrNZnCfIwvwiu0pEHdUZ7KKybXEEyysWhqcEcRThpCvv
fvXDwacebZ7T8CXQJX8Ctqm8wwugcQtMEMB+2Fgp4Krvo0nRWwHf7MKWVibw9zDu
88SRDprvTcNmRsQZHaHvP+GK8XShViLyPkdFEtHCfGwDL4KXrQX12teP2hxkd1lX
6kwdWNqtBQLijoM3civgqbZeOoFdF8xO/NEMV/jVIOU6MhYCN7HODOHpjdkrTyc8
BcR4BNTrE8jJqw8aHDVUa2uNOc50pktcgonNPqKOdhY3LEzErga8Dm3d1RxlBhio
VD53ZPxSn0hTytUgizMSmTMFiFyGVXIw6A8ahxCZiryUCwpoC5V6eLI+/Z7hOye9
sPiLu1L0fuZyUV3GUFNJSzkreI2osHE5JuB+zpp8FTWF242QdIz710Z47p+5fwzl
8A1d7rQhp6skcPSd6bpenF/IQi99fvXjjBEj4uWIMnAm5KncdckttpR9zDyfLxAY
gr1InZ4/vSNxGKh6EqdoFTwGHXAsJD2zHh7NXCndThL6OJuswhruxeznYzIpAhwo
KvNfgOiz58cQxRiyIAgL6ViXtpB1LwE77l+Y0FqmxkF83t/S5WnBUl48bHGuBXBA
NTsBK1eIhbIn0Aq52q/+ffNuPVK5fefR47SOJanFzSqCXXx2gMSSI5mBb4HL0SPi
bzCW89ZLYgy+zQ47eTZMw1D9X7xJ0UpQkZh5lOedKU2u+E2gj2PukxSZe4+VJZiq
ZYkIUzcoqyaG0NNdC0QhjyuyVC4NmC562m6fjjIy0WbsatmF8fA7vYMAH38Gm8SG
iATrULGAGP88ouos/FsH7N+gIW7dUZXwtsOG5Q8jS/v1tHugcExSfMqefFdoRBrq
PO84I5vT1/Qv95ePRNkli36Rq3pixMdn6GScllMmEzVdJ62JfH5tyC7KQiA/LS2e
zAwebE8uoSmaOD3dA/t44DBhOuq1KTh0FbdmI7bOzVn/mNGTUtW8co42NrPjsutd
T+3peogKn2wjfZWm06MELALBIOEVC2kRwm5EEMHBlyDTZXU2Ym+9rRjkvCQ929M+
kDkOp2dLUuIHjZ9XuzFrRZdyIJGMxDu2mwRiq1ZpM5sF+3WstviOIpipw8dw8emq
uTwKXTlr4vfaHbVJJBAEv5DdDd5bz8AIpBLNjz0+zo5NSzZwk4GxUdOFpWYZpuOq
xEyKWLjP0X4dqbdiOKqBFPv/w4k7c3/wZ3DrKB0yfPlsokRlojet8nrugTO0BNJt
JTPA7CJ0IjDTLiydj/VIGmfU49vY4ydmhySfPAl3dnR/AyLV96eGsnQK+29NdJgE
zVNwCqrvGMDcFyLYlJ0NGt38QqVZ/pfckBT8J7DR/hpGjZbrqeFvYMVopmdzr+QA
WDvdNssqr1B/vk7AVV/yHlhnvQIYCX6HEQSLadhWTEjwny+vBYxZaPKScFxz/agH
IB3rL5DhJjzFYoePrKDfYEhZbEWKqDkvdy0hdZDEURRowBxvoY4CGgR1nhyies+R
ZZhmZYZaC7QAbJsEKkGuSW+LpQsO57oC2uCtjzcB5Kt6a8rZ7oQIETRUNKE3sW8p
Y4orpLvXL2D3CFWQDN1eGEoBDSmgllMrGo8URy3X4/h7RcbY31jOfep/geCF2uMF
1NzUThVaNsH8iFcRJdySYnuKgxmBDwYVuQCfoxUVNrUO3p1Ytsj/yom418zOBLEM
NJDAgTNLzGs1MDirkMoTVmb/ztC48bLXSmZvtAfqfpypW25Ni3yirLXvuOOMQjPw
PMPVQpq/6Q3J74IoWVoJnSunudPk2yTRSmcFNoNNydlbhyR38vA7+Vq2RVPPwRyS
rnMKI7Oi6Y85pWXZCMuPo4yfrGlRnlrebZFqvkFBJQOTKcdmenn0vtdw53oB3/sa
UBHR4y5OWtkKJ0QkY8M64x3q7GUU3dc2d6sg1CHsYN77YdMH32MnRI0qWmt6K/c1
7+kfrhAIubbbVghBb9IdmxUBeFmU+ZVoMGo6iAA1zwxIzwS+UDtZ4TLnzKg7DoDy
KbrqS3hkeM+9r+JYoi+0g/LR90wHSQlpefVwsNAmAS0O3gm5dhbc3ThczQb41con
rHd0mjsZQFzoTrT3fT+9HUoWrULftr+jAFfPrVNjawbrShaP+clIVOCqPuAz5W/E
35pwxBDIiRXsdUnUyWVznzeu14wfMTk5tHJIn6pExF+kzjt9ojudKw9c1y8Jt4sQ
6lKyENvA/KTd0TS8h4hPRIMKJbc0njUiemVqT9u9dcGbBPuWJppCqSI+ivD6FN0L
8cnPkgRjUNiAOZoRSFV5prBWTWi+Yfx2jw1vmroBnA3QNfrQFsLV+7T2BbHsUUp5
Y0XizzGpSU92UK+TOtP8zzOiPMd/E9gLeUOWAnLVptkQT8cJsGNTfM3dV6ngvD52
hRNPpMngL0ivvIIBP3w7aq2zW1pcFeEvHNoIC51g9OMaY+0AIs62UOW1uTfhXfEg
j6Bdl4buitevoX7qeY3BwgZQyLw1caHIEm/WRZw8RW0IPpFDRwzDDgPeYHckD+Qq
O3cjG/lRtUfwfIdBcHCZhbWLKL16Bazzq1j++eGj0dXTm1ZUoYh1tf8RcHmiLf5v
05vgGRuBvBEhp3fmX98T0KqvOaPu1RdVCZOLnYD3wvTFwTnFOEVZ4RlrbfVJ8yd/
dFJV0KrY3B6BcjoBjG34jKc9eXYWveE50iJbFCAgGtsYy7rBjOr0FItGsrB5sNg/
Fy/F6PWTn4NNKEFmhtO5tZdn77RhqQ1Qf+HK5NCcUoOfb9qTHnlTA4s16cKaNArp
ffBPiDlJhQZmo97aWVXeWOlCnI5J378xq7uT2bwHh8a6aCUP9R2Jbeb/n7pPYtHN
LiD18Jp3NBhDXD4mBuNwZFWlhNm+GdA/Uydxb4rYReEFWP4X+Ag441nViUN8TRyF
YU7MwvcQ8fzIxnrG/8lsZAPCGg/7cCaOZGKzAkJjAP01blz/C5kAn2INjoyOPbaB
EZXi/3ja3WOAOTGvIMUCk+biALPFd3E5OVWUwnx1yaN5CogrRDmoJCPBcSTnovqJ
/zj3jMpWZSOM0KV4sSHrwuO0tZ8jST9K6ZkCN9mNo6MiZyPVdTI85Dd/Ec+azZE7
0gtgqzYotXCE/dJHyrN2gGiZFxHtjdHheufwFpyJq0G9GB8JKthmMMiN+JLcQo7q
JHY0jE8MADvg3LantU5AMB/+Q+Sk1eSt1EjoRNNEXpvZFKkyuxfIOxOVqlR/lbwU
WhK44RjCY/Tcsby/pPxW/LkQNtwrBa5YDv4yGuyDYGAd4Awud1Bt9IOlscmPFK/y
4cV7h0081StQuLEf6bdPtxF941zVSzneFAm+UlC+uoATFDBeZeIsT8+NDHQ86ZdW
EtqvWb4CQ/aPr2Z+BqPKvBqVzeH1uwgcqvuMBBVGGjEOK5sk6W8DmQc0MMpw7q37
80dDMxVzCaFkVK5iKKpUjWZ8sDYI3fcJaWeQIACP8yQJdpM6kUGpX1KSLx9eC5E7
54ub5355t4uEmlqJg1uhshMqpHKxRZTX69lSRKgd1QLWJQ2/XhNJGWPRWukGf/um
R7ho/QefxZK6+mRFozwxwype9Z4czdPJTsbeejGOlPgVkk7fY59TyinwWrOo+a+U
kh7vrQlcRto/ZpHe9/7J229doTDacJCaotM1w8f4xDBf+O3dB17uIiYz4lY7U8Pa
jtJ53zHv78kJoxjpCe87BQfG1tTdbeA6NgwS+Ve0dQQYira56p0Z+5oNPIVUy09A
qR14CXVDUOHh1nmpAbMRPHLUZscerBgEPCo1nWv9GN44jRuS54oRrZws9XPqrtFq
wdKlhdNkoBinH8scx3JWnX8uGDDFAdRx7ah+Hcxw5RgrXiJNmXQvKb4pjBXVX7qE
nM3Vlc/T7AliSAAo7SIwL1MGsMmTVxDH+tkQDxIdQ10AQOHbw399BmjW8zJmx5dl
5+H0h6n4zL+/IEcanE/0rHzPmwgw01sQIm63qHU2qBluVtvL4XglOO5Ev/45LY+C
zP5RM6p8iUD8BTez5Adb9g2tv2BRG37huAUGvAC79eiHQblu3Eg9iUupN0aohiEc
zdyr21vM6K2tXBbPEmlmsBHrE6Q5+vBYvnxEBRZHsZpqEVHD3cabzIElD3v+cxcj
CXpLIZk22JEYfwTJf10dcuObNwubLxw31RqKQHFXbxy2FwYEGLxOYGaWj9fysiQx
AcEJFne9p4GBnm/wQf3j5TbijQ/m6rhyyNJK+i8x+C69tE9FwkpdwmN5Du86cutY
57/RZ1LOyCcL+8stDOu8UPPy3ZqhrwEIme9tXJlhiFQRiqtuVAtMkeQM5EFvUffe
sCGVvbAhtS98JxlxZUa+jEkoPcpbk5O9vm4Neap+PFFfDF6OWCqyGbElieQmAd1u
qUWmKgDtfLE43I+pSWdMxbieQHKjA1wko3cntTujmJYrNWbJGe63WrpVTlT73SBd
4S5ySP4c6g+BTWu34/NsZSk0vqrTxXm3tBmIZPle5DrGkU+NzT3VPCGHIo7p/FLI
+HckPRcHQyBjYowdBpMAToWRd8sRZ5drsMMp3gGRgni/zwxD4DWbQWbKnkGdoJ0T
+VP3ywFIMW8rn5BktfLgzMp+5DKgJA3KAVlO8D2uf76my97nDcnnb1M5Wdou1rQJ
wkIiItT/D9r42vjn8p2pODRPAaDSZinjkT0byZdb3DGn5EV8GvmuF4L0q7QWh1QV
QX5/WccfsAs2DiGqCWpGr2irenuOnPcu8XQDWGSxw7boV+GsXB1LZinDB6CrPfET
iVAcEk6Ds7hyT9Z/PAfzdsy2UOCgWfpYcpFm6/mqdw0T9Z8AOdZdKprVTAy1PZLJ
Gnu7/Hz8H5/7c+eyk/Ikzr+uikZPL9UdCZTEEPoEj9YJPpgm+FMI0OXEMpHqY+EP
5i9gkM6zKaqdB30U2AC68xVJ5Q+ZUui4pZpXKCiOmPpQXH0w6vgUYki+wSU+7VFB
WwYT26Pa5NV66iQjrw+3uIJ5uLLihxaRLK1Kg8SFOiKziai3Fs42QxaqMhUJy8XX
g7TmlVrARi742ZjBSRosYOSxr+xeg/mpVIPhH13byHz6bWbAMkq7+fCsZI1IaN7z
v4NAkWce/uxGsA0O0CpbSCHu6JOh3GpCp9scaYE2ykOTzUcwoGZzIrocDyb+kqAw
TN+qV8C/NquuBsHfnF4r9Ao1KIdWgAmz9GgyBC6ypGLBw8MfMrsUQySDBWxoCz5M
PHAPTUDoaEprAqaAoQKvXnGlLadYi/0p3tOsI3k4OxdddmiJf229EMTSxUiSTLAj
T0G3DnyoXMJ8v3jG7kNG5RaHgHAjhddeB9V4kmKUc5Lj+HYwks2szXBt/1Ar4kaC
QLA8dVFoAHzQzYLpiLEzP76zwwwyYFgw/jWuTn/b2U4EPM+xrvQT6CnQgEqS3U4b
8gdmmz4LBobrKTtyPhQzio5VzcDXBWXyOVsAzesHaApHOPWMawCUjDICH8sqQGhs
5gF1sWMSvsjmehkTX/8c/SY4XOjNZbWEWm5z6f5SxufLGYdfj/OJOetW+v0d8Vsw
twXUKllGXIJecJPPnpKdNyYuIxnf1yV3RWN1SG3VndpK7UVjUpelC90T+Y8bp9eE
PD5AmyhpXAnpRoZ+0ppIqOLtgfTG7hWAnfALe6Frm2dcdePm5ajNPPU0qdHCKouv
XGU8pAP/L9lwvhj0+xOi6T+r1G5EoFhwHETmnod65JQui0D9B23vBms+f0YQ8CbA
ecdPMXActeJEEe1Rre8TcZv4iE6/q8KjziVzefUwz/GWr82qJJq3G+bPi/ROpjQR
UnKBrEQttzptFLHojl2m/NvMb/ilN2JHJt4YoYpcGtsKCbAQD+9iHKkcj5OXOPhM
MCoxcbp48h/h0ahcIt5oJsa089//EZ7rL0Z2BPs7CHqTBG+6eS8t+KTfYtZiP3e/
1niircxiM+CJNW0eOUiQnrxLBU6s5DFXTPElNiUrmIfM3qCXoM7dldNCJhyNuWcQ
q6kZ09uzkTU40jsPClM/1ayT6OTorfKOtmNrjmSPMgKLoerIXSaRiaW1ARh/EprB
NWUHt5KAlgHuM5P1SiZD71pN3qr1vODrcl9w66CgoI5kV9f+yQKFOhkTlxv791Kd
2pNVeOdaVO/l3Qidp7kqfuVCi5pszQRWIh+DRaxqOvNERrnwIYxKiKTzyM+q6Fhv
CbzYKU0SqIMVOlY6xBikjvInjC1Yv7lj1Sx4vBQ3zBIXa4R8muL05nyvyBt9rr8Q
HNbibid1pqsLbo8fqFgLmJLEb7nJtRKWIaLKAtIhTXaqA3sjBOz+rfbFEAGdTkG2
DHRrZn2CTL72+BhNG0u5Bu00I+khrhPk9eaP7HaISTMpT64W/m7+0pPm6eVz5N9T
ch6z3jy0RxuzOrI2fcBFk8QXlSzZcNoq1kiCFk2c7AYifH9E8FLYCAOASAy9mCx+
1BsmnMt6CLGEwpAiZY0zLG/YQnlWrqCiKQh4CPaj03e6QgIwuip6oMPOHg2cIBGk
dOllW3Z8KMjIusyZxnKPKk58a/S+FqY2CrQhRT2Ez9uqOSx/xWW0tCBXscE6JiB4
euD7avRdvvywx/q8UaEK1P+AMAtbpHYq7gP8fEn2vdnoRR1HoiYpGBIj5H1Mw0a/
e19VGSEkIanXeFagqGttG+yZa+IMJvqAtm/FB6RPf6urqemFEAX7gZs5N72gm+Wy
fYntjYOaThvRQ5yo3GfPSHMau+lU8enbe7rxEDfZTH+fOKx+lYqplU85X5dwT0Cs
EGJtJPIcJ7oZ7PeYMoMSwrxmSAgcHkrz4iuO+9M2XtUlixK1y2o+bhDebPbh7YfK
T7NnK7IH0n8uahFO55YmeOClAIVcJydlipPrrWK0TS4HPBakrXkTHQz5GohVf7sa
BM1eCgqIZey9HJLaDFxocZqaYD4yydgQPuZObeIaEYN6KrP1zWlHw0n2fxPkZN62
6fFslROBqVB3dt9SoUMSNcjmTwuY2cgsgXTfSQ9vU2Gsv/hucBikPhri37wWOeO7
IhS3wsO8iWsCnFTY0defE9i4d2r7B8zzeAsFLnHqdqMLA/XFJoiIMCixFsQqsH/8
TqwcjDgld3M5QMuerW6ALr7jkc/0HS80W/OSjz4tJWhgaINL2leLiqnOx1QpB7jK
ONVAkc8y8GSvVHkfYyxakYrOeRwIh/fo3OTxotZNjHb7yhhQZByjWE04XVb6pUQa
B48pIBWl7mRG+0iCAOhuSxFtXtV2x4eUbJHe3O4lvP9IvHpHNYiaG29nZneSTI1Q
dbAVHNvtSzmIFZWtNeZckGN4RCCv/JHrBBUQ2/nQn3rL/OCMVt/iJAYiQUcvJyTk
JxEzzz0EctexitEFppltK1bpeBUXU046PypxVxclU0kjrlAkvyzqYYO+HAfoadOd
FyLw8RJ9jVIyPaH5PFUMVg/cuf+auLtxmxB4bdhufv7XZw5eQ1XLt2PdusrTGi5t
yRRQawKb/kKGNE+Qms8cVvxKm3ZsVjsg0hAomom1J8rtcHNVJdDqhynb45fqM/4X
t4aGzwMSfxQ2/cxB0NhlKMRHqizDg5Bwapu/+hJJduY3DlfhyYvRbl0rb8bjDJxU
wffMbTYRhGBdsdxmfWPe1jVNsmYApoaJAhH/dTM9N0Io27kHoQ0z1eI11qqrgj6T
UCUlfkkFpb/hiwiRSVnR9RlOi3fFuyOPRStf3W/tSNxa/gUL9WC9PiyNzxu0Do5N
ePswsY30Nh7aDtmVrK695AhbyOHWw44IrMgPO50eTyyLwNUXQXe1vVouQfY2V+hu
YysUni9ZnKkj48A5tuIDVOOSmo0U/cT0/TvhWDqBF/B3A/+AIr9FtcRyVQPw//3y
+3C5zgz5QhMA0SZFhHg8RElFdoxCIdeDLhP4s47J/8QxfIKdi8N0JPPUpJUMk17q
+pfYXqSZt+2LBFPFwRBy2HOSe1576M9lV7P+XeYEQMbt4X1lFX7a9TdN9jw53Rzs
Cle/nbWIByhfcsb9HXjI/7u3IRaPNnQsmtM5Xpjiib5BLkr18spXApIxSonn84tu
GrcUSBa8/5HyrXe7pTHwFkiKMeChV8jQ3kyFlWo9IThcrHqaS0Yu4i/va5JgN8Ey
vBwUvCOgBjp4AHHSJXq7WdFNmHi1LDtA/RUii8CuGA4NcRMCo7n5irMXW/+4nTE0
utZkxv7B0P/pd1gbNccna4JqcUyL9k928eeT3JAi+gEcR4feHpDb5nC7C9YwrovE
WyJCzyIhxeiZusjO4DKCH27Cr1675EeDLgef+PlH54khINIcMm6moAxQ9CbtNgNK
TapZAKI9Bi82B7hGs4CsKPRQOca/UThmDGp4JGQvkifNOe6iyuYmase9f0K7XMPq
95hbom32v14JQhKS5wZ2T0Osuz7vinzqy5rb6N+w2JSG/ulZJocBJr6wzDLswpdb
jyH0SGqCqDsZmLc9FExBlhu8p3s+f6T8HVQEf5DnhX2GbeUdX3fhg2/9I7RYT5Le
wwFOccxuL3gLXkmjn0h/50UtjksLQs/zXUsDUwobRtQtXySSJ3PEucpOJXcu1Ic1
zRFcvqwLsdSu46snIhlUf8WDJ4vXgYumigoVrGcHvtXTab5ZeOBphgodgp54VZua
36M+t47z5Vbk9McBJch0RNy0c+qOTqJkiD0tljWVLntlSkuztOwTBRX79SyxbOKC
PNq/JFrTlJ3G+KAF3lVGhkgerfPRpdOEvQfHl8MvYCYwsOjExY+1an0u8fBuw38X
rK6JNH4pS6f3EYSZHsombe/yKt6TN7xlAFxt8IKGWuRJ98KtY7sEnI0c5587SjIl
lEqqFfpcYpR2lGcdpymxmcJJ6PxxCOGm1KytCbrNsnh81HH4zttzvw9Sk+TcENVZ
7NVNk7vY5gxrLRrDK4KKJPB+YCXjT1QE1tTrO/w/eeDMwIp02yCe0eMNZ2VZf5zN
EvUvdVsTDfizJOdLBMc0EP46nkoFTzf5rTL4T/I271DeHs/vWmnvFSC9Utb2Gafi
Un18V1/Q2AyErABnrPm60GMZ0/k+lDkacxv5MCTOdinn+iakN0uYmuaM0hIyOT7c
CW2trChqR36Vv+UvM7lqpPqezMoE81QREAC+1nBVSyfVmaUf1IZHD5IvCSIK2Duy
ZB1Ph2MxyGXLev9nqGWV1cCqT08Cg6nH+3v3zwkQ8hhymWeldDE5PZNRERyVNPk9
`protect END_PROTECTED
