`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XbYfv1lQKdxrHBW/y5SmufOO0hcnqTA20JBtDrObEVeoanXHjJ3r1yAH4bxVaRXa
UCyCDP1O0CHX0UCbNFs5LXgXcWsPN44U6F1wk1jdUNyXPdZJwz8Btvh7yXzCF2kX
M5EgmwIGqB3eR0YnMyrdej9e5J1nboSf8TL7kPsGNX3wpnXPWM9noKmMtjxKxwMN
MJPAcA7DLqBfNKpcIQHaXz06/CckBaW98ptXGYd4zY6NvcpJaZX0FDKc56PnlUI4
Tgw3o7ky1HYrFXLiJBpCzzyHCLgTChP6k2L+Eyv3lcZV7sE466cxxuW+Ry49ySPx
GPXPN8O1OKH99koDjHYn2rSOWCFl2M6exbA/TIhp2t7mEVGlZloJJKDkhlsejMeK
wDfj9bonjedtVU4rdaGpOBI71ZjaR9zrJuw0D0HJCwdtZnNkqQi3CLx7j+DcPXI3
IUKPObCYUehuITQRKr1dWD28JWBkvfSz9ddYEWPWICpLLmI7ddAptmLqt923pW1U
89pxlARrb3OQJ1122rKsp3W3VXLWhhk82JRoU9U9o7/yGbj4T3mMXwvJIwng5Cqs
NruKLyzOOFApfC6MShqEwanfOIFz8Rqpd2bGnyOBlIRfH5BSwo9YhXrGZ8DJJ2KY
ZFv0IAoYrqbeq7fxHt2igC/clK0kF3JRpvB4q3YSonk=
`protect END_PROTECTED
