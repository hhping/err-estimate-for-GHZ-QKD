`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1LWJJyhvpoluaEppcDO7bwOg4SNXnrhUkwXBSdbqWlUfwybslZ6m9lu5ZceYClka
Lsf+Y1kEKk0KI/3irv3/XttAQdQ6I1UMIxKI5Pt2QAUntgZ0WgtO1GkamfKIxwgJ
pS1YxUikYUT5HUyxcIeGAcyQe43zMQKhTKOiTa5sd6KE8yHhebVS3wwm0nxwplg2
dErT/GzJM0j9ttA8RqQ1eIdnt71uGBbCv4zOiWgyx8msz182M4T9mcDcpk8dCLLL
o/PIl1xyi71xGIddTvTJA469Zp+ZP3eskhWdiq3cUFTqjEtwRD0RFy0bmS+Qmepb
uum3VMC+YAukTg9deu8c4MJLPnmtGoF7W1lymKglKLvtR0qynbMjkam5w8Au1R7t
tPcQ8DP13bHBVelDmUpaI1jmj64tsBdIJ59mOM5fhc6Ul6XgnbZ8HpqqvueEvpvf
PAMgPhTI6LDuPuildsUaOHrAYaFwrr02+qIyVZgKFy7U2TbI0z5bRXJpGBZ9lgW6
JIAAEXRPeV6x7OVThVjEg3EkeuicL6pUl9MHwy/JgTbO5yTLLs/LBEZRi/OAAbr7
vmNP0+rvm+s7OM1c32ERIx2jjCJ78NtIK5mvQ03/LNQ5MQcMWeZvn+j9xXCnW/eU
8idXBrrZe721QXeITljJFA==
`protect END_PROTECTED
