`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J0eqEybRx1Gw7nCT0xlWRCWPieKWIcJX1wjqYIGMS3dkGaSlpxteHra2vVocXW44
eUAUFesLRTQJf4aYWeeYa4SSFHuAS/4gN4FKhlNXMk0m02aZhUOYrQpGe3NMXeU5
SZpfEFlR11fuYrtWUv/Ooa4XXQYpH4gYcx5boY47G6/A74dRpUM/J3DZJzaFpPLy
zZ8cP7u+D9PYz89NjIZO1BFY+QuaoC3CmB4Li7u+S7tXTlT0r17WqGO1aVdc6R+t
0KT34PXYL5G2caNMyHIWPstfhm62ZJDMGxrp2welCOJfb05VTQ4YYsBr0pDUVuOg
0ETmgHDKI6rF23LU95iZuYX5g8VXh9ITYozAK+rL3W2oqGem4ryrHABAmbhWJSd1
tjTJ+P0apmvStwHknQNgOlvNthex6rGBQiic4AtL+As6lAvCAfF4fFMnbye2loiX
ZbMhjivKU/DC0wO/QUeGGq0fo4I4d3z5Zx+xqQyMFOB0esuQmRy+jgvjC2vLF4jM
rsBuOfQRytf/V7sTvdnddgo/nTHUVIIrepYX4l8+Ra0=
`protect END_PROTECTED
