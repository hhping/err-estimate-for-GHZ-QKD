`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JG/E6gKq0MTPpZKTIW1ucHoWiW1O79M/WOgmVvFmj/P8ermrfVhd5sMgDKi8aMRA
jYi9RGXbGIpttsOS555sWY7TGrv5M4gKjSMjV+f99I6psjaF4t+04FlSGXW3Cjfd
i7KvqHwomAzK/1DFlFmMLwi8Zz0py7HYjJ5s3frCQgZugU4aMBWy7LN3QJJpuowX
Ukjskw8IBqQskJH/rW3I89WWzT9ChAolUjD+Pqy4/5R39X8JrY3UFIDOtedSgB0I
OuVJsyIm5XNT0kQP8LBfuul7Lk8AzU/xbDJZxZwUIPaVvA0XG4tQsuTczrPlHQwI
T3a83mZqWoQsUOfAMLVBiD3IusFnIP1SaoO/HZ7h2GfUaAyTQX0jb2swdusDtUCS
JgxQi2qmjZHl4pK9g0ntM/TnyDZ+Fb8VPvZ6TFnWgZRI1OALtq9fVHAON0Io89Df
cmorMWkbDbuLECgDPRCQxIGsiezopaZTtl9/b1GvF8dxlbw+76qqWL0akDEW7a6t
S9R6a8LsRHsVzA028lusw0d2Kstq8ybyG5uY+s5yP0+nZ4yw1W1do3HeGRYElvSS
rFyaJsAXOsCdQU85hE6sZmJxVf5yY87Rc2UOWVSHhg3HXkwjvZAWRi1b+CPtSu3c
NZA7BZh8K5zfVL/nP5C5LnvB3VNE1pMODLgugdiD817hIZVS53gbKLTb96F8PsyZ
RQuaRUgHsu55oiV6wbBX05xUsqdiKsckagnKxb+chS+Pw84limiOgSkHsyXl6oBv
n2+Nq30Hv831dT9tZjOM3BIRHXvgciJwP35tWSCZLjjrFHJxUe6sINlqTyXDQc34
4NZxbAC1Umzs4X841kkNsoYXSLFnjVlHrzD6dKuwHjGy2JtA6rOALzFR4DYZfoS4
4ZkfRghktZ4aSHsFIaWb9U932ka0lXqeeRaxDh/xjKLz8J2KAEdNvaivHRAXsK4v
iHrklhtdnMZ672f8qNR5HedYURCFKfkrD3XJvRY1F+kC9SbS+X4FpPTAas0LuB8D
cQcvR39NIzyGKugH8TOh4WxFiHlLVVE9EZWcqDWnMcJrO76v+kEGA+Zf1H6icb7G
SGqapgRvt6drEGJYxXzDjECWf2GjnKbtv3iMfFaHKQmRwcFiof+LKYurDBfgI23+
mWxYokVKIH7Wfu08vQibdc2PWQX+vhVIyx4AynXnMG9rVGfR105pK+OshZJMxxwx
hA3SXNPqV0jFreTPOg85U3Lr0xqdeR3zNa2wqQ7djf4aJIFQltkKcCwyTpilKHUZ
DEdTEzjegVGWanHZz/5kYZIkcqLRQcoPnS7JiSSGsd2GrSqOAj3xsPl3vxRAAUdt
xhgJWqf74fqrdQXbV0D+wQkgL75/tyD2gFxrei40OQHLNDJXeV8HIer/ZrNE3lx7
osremJBZFQjhp647WliCoxEKYglmoCFTvnmgm+NnZxO5mg2R8IiKxeTYO9XQUm7R
9jnbLu4sYpEYkTXm/zO31L+CLEKJCPYSxmXqWLAEOWU7GvwwrN2tXkbzTt7kKVZ/
X0PYAqAcCWLLGMklQq2a1tQLaKsjRdaNG5G2x3YYPPMxgSK+2HkhUsw4AhsNB5XB
h097MyZe3vnHrK0tqnaf3WksttDJiKtelmkxfFcopeYeI38CSTvADLHCntNlPN4c
cCrShihK92IoVM/bp4kY7RYrgROk469Osy2DoqQyh/BIJjF1oA4Nv9xoLac2wZxE
3J9pp1n77aD5aWMrgXDwE0TR5cSI4lrqH3BKL6BocQYzJp8nlG+JPABFoC7TaVzi
A81iaABJsr30gBKpvhMZiFegJLomNve4J9EdnMXKfSzcAcPsJPo/v49FcFbZ9h0O
jl8VRQhNjJUqHb/4X69w5nOCDf8cNTmAGJU70ggK3EfBkcCXvIymp5WZpp2KFtc/
KnoosNuKLZRpNOFp5QiuBPCBiC6Nt+SIz0W+BTm7tYrya2Toxw+rMJjQncXAAVOU
HP86q8OJiTHDaxunRdDK86LFAPqZ3I0KfTeWCfPIacdde91+ar9ZeTm/rBrvBD0H
8DkYwRZqfcWWpaGBAQqdsfjVGAjeI2Geqg7G8KtkZrgyGv21/LQWkz/lyEcnQ0cK
8vFQKWVsU7sPfh2F934AnWFbrD/hHJfaaJu/gDWh4UNVXIo0tfQOTH0LFRuk6oIq
TPTk1Egn6Jy9t2oRUZk20uIi1z6h7UfFMb6D7AZm0Ll1b+JY3GzoF6aNrOgiRrW0
O5hSPci5StZCrunIfb2aPZIZqshX9Xff4Ko8qnm/oLWQQLe3y6vN01xihcNS0shU
IvtUbXaEh7Z0ctCHqrrLtksL94Cl/O/x5wpN7SSK+Lyppc7KbAc29zhRRbw5Q5t2
yeFQd+0zO4dUzqnUddigqrlpa+ey72tw/yBtGf9+mYlqJ5a4ggExbQ6m/Dht+Ctf
UqPoREOOVOHVOLSXOIUt5XgMAQ/HCY2IH7MggmVmtkmd9gzvK65T4qa8VvT5G/St
zMNyORQjrha+oGxxBDxi8H6tjAS5682sTfvyOqBEZZQ=
`protect END_PROTECTED
