`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9G/WSWbfHMaCR2W0J+/bWGbKZQ0Qy459M6cXH5325Z3Q4PHzPaubGp20BfUBivVH
UHPnYC2k/WxO+HwUaw3NsGs2jgl50p7Nvi8bIlEcJlC952fvMIdMyeV6lYDrCgo5
q6EECl3zlOXPpaoFKCH8zOSk8bKTh/1WX/HkgHDydiCK5b6eJLovdZQC94Gs96jm
KtiLKEdEzByMzch3bwGwN8E0ZuNWReOTPwYWoJsAnwBT5p7LOW6H+PEz/ef+3Lwg
dbbsalklG2Y5JkG1zSlDVXQ3JZuhiCGw923n1TyeiOf0IC5ngDHATe31ZuRr89RC
HqOFLGyE9O3oj8rqcscO8fkg8VJbo1QvDcjKR+iRfUsZYEml+jPWYJjf6Pj4OHbI
i6f8/vaH2DxT70Bxo4EFDPmMOJNHyrd1KtT8uumzvrfKD+PmKe2YlyzDLq+XE38v
j5Y85IEwjO1jEvyqOhmwuwWZN5PRYJCcIWXhKdpqWCc+jSstcF0fyegMw9qsBtw2
DHoNOHWrC8RD7Z1Z0NeF55ftugkD+AXnyatrfUZ6J7E/34TIM9XoFOzTdO5z5DUf
MSmB0MFAmEtQHiYuz9DzhpeE4vHJ1eky0rGwaWeLyR2Q+ihFWMtQ9Md5xh5up/Kt
feNgtr0JLHUqg7CEgoCIg4sCkArQyGPXMFRnyjFLPfk=
`protect END_PROTECTED
