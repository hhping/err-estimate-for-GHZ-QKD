`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AOwhT49HPUGNBVROGWDdx+M39Y9vDGwjXycRh/HArvVBQvuG/mQ0aP8CjC6ET5Ji
PG7PId3pX4l9f4x0KsTzswzBuosq/pQErlSLncNm1lpV+CaieG71m1XR7VlWIej8
SQL3XhcyAAtMI6a/s1xtEDdVZKHHyACMUyW73t9ZfnplXx6Nl8XCwjoYZTF5/ojw
fFUMoES0yvvIHEaTziuWz+16PdnOn/PEqmHsjf1yBkm+YZxFi73Zi98tRgXmPDo2
fyvu+IbYV0DmOdB1ZptcHU15OzMuMpgKT2b8w0xtFhYm/H4kQg+N2u/rTUQXUzjE
obFsLzhfyUJiP8sh1GLtZGMCfbHYe/xfrvs3sABwzyFSwE+jhh9IVwfTqkaQCakt
v59WR+F8Df2LW4GPrhW4iBbQuLWxOgAqMdhe1MC9JjBQXSx1nCFYaRkfHUo6QZXJ
YJFEks2QgqfuekHwMid4zlkcC2Ih9+12Ky6vc2wOsQgMP/85WNz3/snXajYdHodm
qLtDiFMp8wtlZDA2bND3a2VZqM8zCUGr/GS77/OW4yAxKPiyXtGaFmSV/XkriGDT
3BsbrP9puM7i3OTIqhNqfDbgWrq+iwTWT2HRG1uDGhLCGN0jXz7EnLlKWfwdef/S
GimRzUHaZXzRu0pnWG9LqMZaoQ1WA5Tf0lNFK3qYyVgz6Ny9mx6UGgIBzzdTRN48
2F2ZMAfVS1IkxfBCpXRL+nIBfxmgbtCwofonXRjJgwB4xkFoLZMoSt+WQNYZp7nB
MK19amY6YMvNzqqJvPkVOA2+2jllP9xD4FisZw0esLT5pJnux4pEXcArBjwvUyx5
xxHZ+YgWQgqW+NReeGTFmPgSA2ov6Rx3SJ5XSTt8yAM68hCjUeyjWmAPKCX0ujMO
K/tY3cGaQf8TEATjrgpvFx6BX4MyukijlbgHVhaD3CLu0Y5Zlykq4ZjlPUsolil4
FWT+sWRFJodWJUKyH1KY+u+1ch19hItCTckAtj6pEDAEFN4mtbIGrfaQ0L75TlyW
oCbKJgHPz87VlBojxbn+40bnGTHfTAwa+gdrm2OrBZ4agRLMbvFYv64fyuenXss+
lSOGuBSOzxyyatRm/olfNy4kLicn05gcpDGjMyERCj832ceYLu/Zj+m7mXymBIF9
xB6QI2HRPNl6Dl6lpvoej1UePVOAFymijMBHNwO73wzK4ELqpTeuOVVOwczKrmkT
o9R0poZcnCO32XOmxuMcr/HJhS+Dxv71ZV+5HpIyGmFlscsmxZ1PmaYbMeTmi0Ld
M9R1gfEIY3PM8Rp2K0m64lZX2UutELEaUjpIcWmOi185LtpTQUHywnybdzrWDkmU
4Q4Wgcr+8up3+tsqIotIcLDJxicIiVsib43EqY89wF1AKhhxUgRCZN+rSxixYLYZ
okP3ijFXLaVocImNF7KneAZtVRKJvzrP6Mkkxmg+XZJuKWD0sXsVvsgt21Z+qfYU
WCoMLR/jSTV8j+0o1QvxrxXw2Ku6wmfS15H8GWAKMvA=
`protect END_PROTECTED
