`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sw+seQjdAxMJSbMP3HA/2/IjUFPH75WXtgdfpuCpUG87d2eZu7hCkpawVsJ1AvX1
kVEHoxvicBkkyv5/zciRNXCQOKsswF8QqPw4YXYe7t7gkvsKzGwfCcSh8Nbk35fE
miDqI/Ml3ofkSVHAEZtXSxiieNrJQBUhmcQIRacifGfEo+2E+tDaZDUMgTKfq/sC
H26QqztRaoezYwC+gxmTx3ax/6RLdAVmUEQzerAofDdGhLURfb5YW7dvZsf6hTd+
4Y/VkEjyni/ykC8ekhPi0qedEuFVo//wX+nIeTnrzdV3+SnVqKUZNPcsZIpYL4B+
itY4uSzzCxZhXfQKp+y41kfQB1/TRsgIhuUl/DSh5WkcZTD8+Zui6V8ET2RPD7MX
2fWQS0CmW4Xwq6bGnY/Rr7ypnVyVj2XVSJ8crTwNWnE7xC7S5y8iGknECdSIo14n
oQIPc8xZIbqPEj9mcReYkIh2LJ1KMR5I9u2IuIPNGTA4eOfEFmoceR99bmosov8q
+bIEVdTYpRC0+4mGyzdXY4OUrf7saeWl6MwB1qCVmBKjwHPnP5JSWAJGJZStrb8A
YS+y1g9TjSJ5E7b2TTmNJbDsA907Xm9TLN+ezCUMiWSnUcZa+LSq3z65Jvrp4BFe
RXLtvD1h3Bh/5GltYime3ehhzVtd9Qczkllar3l2b7WAjtIzeAptdMm4VHWzQX0+
MHrjfbj7755EetkocKCOocm0+evG1XMo3JugsEMKN4b+byRnfbmtKGCyLJVNQyb3
8s+uw5DLUF4BIW+P4U62zczsFCgIsiNcSS4zIuUSdU66T0opdse6yB1tWeJEyBCy
GWrXn+hdaCOYqYHE9TOA4B19xFrp5vUm24ITsxc0Pr7QBTLOAyU3HdOxXWoLZPjl
`protect END_PROTECTED
