`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9VX989CUfHcP/ltkmYo/HjTjAZpZW8XFcmOwcofsuHcPWd7QMT002k+ximwU2a/L
aNXWk+igzec2dCXiN4yDQcGxBTxzvPfJWLa8ZXcjJV8LZMyxzDtib2zZG4sImQgs
dUXch1F2jdQDhn0y0GnTfDt2jzojzEeGc6plupIF2LBD281zbfTj42NuSrQ7caSL
7Xg00c0a8d8PZni1P0pfIf3aelKSqXo5BGXBpx7tFR+PtBJ8jm0LIgFrmTDPFk5G
O3JXZJp0ELu05s+xcBmShMWW4KSjOY5An+gYG1Kj0JDrnLAgpZEfWrXfb2fNU2Ox
FqxzfVVaPy82fy2qMfUXIYHvnoDBvginQQ5I9fwfnk/Doq3jbCn8xQedVCpqu9t3
bg9hT2wYSVZ2g73wfh0zsPN4WmCVdSIF9XwpvGiQHo74Nen3RKbAZwpvjYarULi7
jKqHvGq7dtRaoqqgUGeV7JhCb58QkN1UtzA8KYJn6s13uazcqvQ/dBXtAKADluIi
mJY4Kn7VIujPPnNsIfJ8kRfqxWhI9EJFx7uJWxK/cTzbooiLDTEPbuZvROP3HpZq
peBCIrUzuHvsjFeS/7Aqtqw9lQamKMNWmKEf3TqbI3XE+IDlNXWfId/SyQqcDUpx
fKVkF2IR9k0OK0u2UWuzMCKqkxrJbG+gkpf8BRCUqjpbCVS6X6YKm776EJ50L7Ph
kxjmPn/jOlidh4yGuis2vy/BTimKpiPtPyISyUxbrwXFSDilk5Scj3zDCm9tJ/Xs
Da1V+OlQmLk3xoZD76ESQvSJws71+wqzhopacXO+5TeA3p9Csf3CaWcd3rmEhEd3
Ivhgx74VO9fKHSco+oeOgV4e08x8roWliBAn0CHXxiHkObgSn0g2W31a4C1Of5JD
ohTInWDuVA/+5+EkfcQ8yWjUyZ3iyV7pbp1UZePG4Dbz1Qg2FJeNYO7JQLdowhl9
DBssRrg6omig0R5CxeD7eAZh/OHwAiHV0j+37A1mIYy1TyeocOjgWKcWU5cW/Og6
zfiwXnF99YFszI+Am6Qd+Ex3oTP8G551uY+BOVvdwPEzjdDg1pdDm5YPg+J1dPmq
uxYMCta1ol3BzlTylebwDroiHP92DYl1oj/2sRTjqdve3AQfw9V9JvKkAXwBBb29
WA5d2FUtuRXaIdJ3dcXsK0iEbi41D0H+34baoBB6Na0jfQYyY0xw2NCYa6dsojgm
gvqduzcnkHalHj+xFK2klMUSUGai7bBqqUUI690Bue8=
`protect END_PROTECTED
