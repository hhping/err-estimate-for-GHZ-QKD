`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F90imf2u1FGx575TZlOUBCT6sX2x6jOcwgJbJpdKSHi/rI/7mOU1HMrFZWDBuXqu
0WtsS/Rb1eVsh8wjYcuK+Twti+hBftTbw1ORr04F5OjmujP/PVqLcP9SvQj/G/fg
oz5cr0GuQEPJKyF1cF1onxOU1ookfWY3dC+xf5l7OtooWcLyyQHfSyfcmoLmqg9C
yeYGmLTtNU1sqgPVm+My/iOyibEacnRjUDZWIlLC20HrAaFor0pziJUmAEAZzku6
tbfCQXGUiJkVuX11TN6Ll0yRWwyzCMTpmmItGOFr59J3t6i5vizXqEo20rLbzvif
S7Ww0WNArWBTFION03TI0p9pZTHMc93CP6bjfwCFoxuf539ZU8Ket1UK9yR6HqKf
Mc4CcT3ojDcMnfp6d+9117zcZkT19xVGCrKRdHaLf2iDyJvpKhi+7yx9aYczHbHk
t9ZODtdpYhQB6oOzNqF2LD/3fz9AhQwiRKjRGVjgdVJ91m8Y7r2DG0aORH74dW0t
J4PzbTFzaFY9xHahCTiPtx1ZG0ARtqRqxHl1s1g10EwD7rtfrQh4jAuSBjqGuEui
Xz+EMNGW1TH9qa1dEDlIUc3aY+Mjd/w04S9hk2ErmoZg64WhyYwIrKd8NMyVMlqq
naPr0rC1uAn9K9Wu1C7CLjkXRERFSh+tNdBSrNQViV9vBIIrn5One3IPxOinL/ld
hBwahpwCDRq5j02DjnZCiAUyZ1U/NvIhe1mbljAgChalvUc+M16gasbjk709+ALQ
1qNu5WC0eY+vplKuOH2eGvl0U8BehyPI9a+L1/PqtpCpfzzoTwkKKy0IDOJWtNkp
70GE+DkomItGQN1m09uMjWTEoCmwpgbqm7roM541wFZSdsIKABTfQrdnc1xFkJk4
93/TFvCsLvNLB6ggoyrOB+IGjc4S63sfv/fj7dQMrQF6si1H17myx1JvKOvMSR32
uPdgyS942BVjqu5xJYNw0OrmFgyA57mlQgnwY/NvTyVVpwfsFirq0ib3uxZ4U5Qy
xhigztbHuoFvbedlDMelVe2ew8AE59SOtfUNZLG9Hou2qaxk3zElzxwT/Y/AUdrk
yAhEAaCDBii2Bpd/40R1lEPglzmJNaF6EYBdsgD9nMqVGUTrRPkUiyioaHZVsQBC
tT2W75+AUVta0GTOGt6b/fnaXczVT5Rhm5zAugqh/3VtOxp2/PJCLjs0pgGhiCZJ
W40sO9IFx++76ZzoyRkJZ7YxXOrE8vWaQlrgXJxqsJIiqQPXXCjwAqpR3/c83OlO
bdhKixYbedgWDO5WH9zVkK3M+/Itz0308Y7mXUmmbqupa7T0OWyJDwURDdz1i5Pg
AuTji+wfgZWZX6o0eQ/PaCDOyKIOtrARXQv+Gi2jh2Pi9L1Z9XZW/8EWOhj9nrPA
pbexYOXVLPLsmiQ43JqfLVMCKoqyUCTyNifC4wsvfEe8nWDj74lA1kPw/eonejgV
4jcOCOy+Hjmd1YmAaE8wjgitAy/YmpQsGffnoa+ozcpL6QE068KflmaApoJklfsp
HWwl09k3Re2sSZ4XmlZ5XUOz7mCx/tPOQznYZ8Bj+pPjkNszhBgwJmr6350rS7jJ
QXSTWK2es2if1qwt6D2stuOcpW/SN7t8LBxIogYZxt/kkJjzWDwNAn4gy32j/czQ
sQ9oqJoIiLXPwe8hAbtoyvphMDj7GDUaY1xKAw75A52zMred9gAF4G5tZbX5lqiE
ojKoKsHl0M6xs/XdzxuCz5dC4LmajVRYrE9NhOzRXlbuBBmBolFQDJ4QWnlS2BY3
Z2kW8ndEtXjBKcxyVN7Ni7HW/+yJnGwpXW9veszTx6c5NVKUbs2/WtR3Km/Mbm3l
HMHvAbxEuEOVlN2YczpbeZFSgKtKYJWqxGAaoKo50GtVWGhwHvgRPFoT71rp24Y3
vJ+S+R540DJHsd5SlN37foUgTMTJObyL5Eabeh2Shu0lLNzNvJlQhC09t7aZBx8F
6hM9Hn2IuugouLyHlaev2yN4aaKIVFOOOCP4G/2PX5zJw51D0O0lQN4TMr44GXbz
Up+d9Jt83qguxcNiKsIPwws6leNEjwegFzBVlrlfpJHMfGtZIf4ScnHCy4JOqu09
TEuucfHek6HyG9mGAy1qVEloMMa+hoS2Rh+z717345BpnOhuU8CUe/RaAipPQ4Kf
/MPVzI5D54ic/c/KfVqkYH0E79lfEbPHqLbnW77iF3XwfugILqVJeTKHQlHcKHTL
fr/OXClVjaNB7poW9CAPU2zTGpwT8egnSwBBCL891wZ9Z8Ctjyxm7sqphnEh/PqC
hhspUMOwFv+kvKVaAlIyukJ3maLESYCli898Td8HmI47q77Z4Tx0j69fk0DsarQl
56z20mZ3std6UKFVVazwwCMd5Br/JSw3rENYBTmEIhYv4D83g1s3of1YGx8W695T
1QwrYcs53VgglG6oUNbOzXLsRy1xQ9Rwze9hNhoqF67dYgv8MpE9RwbN7V2Aat1I
J5LUMxc+fAaSQAqmmjTBBEoFoiGCd3Q6olECGawkRPpsJzXls1qlOwSxq67M+toX
q73U5/y/WzQIP4N5Gn4riS+BGqBROvSMVk54X80kms7t07Ed0pQ2QIedOeP5ESu8
XfblJc4BbkEeSLqG4571EH6jPfb/C7ZW/XMTi9sazWMffmzvDxwujmSS/Oiu85eV
9gc7bZeVE0k8wvmmucin+gAuxHe1JL7MgbAGGqAyGCr2JWujQ3rBYIUe90OF9G4z
9xiVWKGHKgJmrNfEYsCRtXkaRHUSpPhNQ9v1NBDCcxssIp+ESlSsGPuwZXg77uPV
ach1qpvzLpinAycEgYZpxMxOJ+vOHpFtdB7NE+4RopfiHrgHoRhEDO4K5iqc99Le
4e1iZwCCZ3RxCcTwDLq60/UXt7huu32qa4ZQwj6iN2jNk+PiZ0wna2mTgLkH2jft
q1gb1ezVF29cmCwkDjTqETyEV2pkh9s4zXgEppXuUSKekPTbrDehKTBE8g2MrDaS
UCEfPJ4hVM7lmrAcpV8eZmPg79Z2sUiSL87dxFEeAYa6qgk9ypem0MWN0Wr5si4H
MtjdBqvI0h6+LwUmsryl4110g010+3BmV7d8mZQnEmeZbXlUFAJ/zbl6gE+qecok
FuTPOFHkRFaVHXkzkXJ3MXBD1he3BE5pEXjPQ0cjqFzXZ8IzqSNxe6X7lENSo18F
LtQINjKor/0VAbt452oMfddgYRDNdZR4fBLlliTz/PQavKbZ99tGCgszhd+4bZ2N
VvCVrpCmVlY22WMYGDawF1m4ZCLAAuRpk3mw+f+KMGTtC1hypGszH3XZEgUj3Gu/
cUjqjq8YKrguL3DLjKWzcZXNl2ZhYcoLxYoOr7sR9fqlRMpxgMyMfIfkxo/chJp6
7dShMROcC98Wobff/uwKr7fvK12p+XU3Y/VTH6zzHPorwiAaEeKv45zUuG17nuVT
eTuUxgCXYzmXGIMpI3tRujetX3HAYfahGkfXm08smZdXL4APTXECB73A0CCkg2vY
g8FtZEQwQ1T0UxLXU1GRLnsiSMN/FyGZInPLMDzMwLIzf02BJtGry0dPaLR25XON
60TSSGSLLKnyArEH08SVryP+7l9WMwBW8QmtpAX1DY9e4qbnAFpJ+am8N65G65vD
TVIzv/HtxUpmsJigXYkiEzf3dD4PEaFvbTcsjbh/DpsuVyvt3dDpcbVebDEVhJqs
Kh2IYT0Rn8BVrg814QY7E+DiBJJb0ajVx+/WYY9LTdCnMnMTFrZ42o0oz2mmjSVJ
WmwgVCP/D4KuGORP+A06qNviAjxvcEFZV8HbUT4rZqd2B31B6uGPV+DA/QQn2rxc
y5raRbumyd0E4F0hLpXmwHzUAxXa6seTp3wfsfuGJnRxHmYny/Iz+tYZ5jAqoZY+
oUaXEvj8422dZb36hIOSu/Ls1bJasRtINsSb7EQAxYju8fCUmo1ghuo2494ImrnE
9T8l6+cGLSDejBTWXIdgY4HDWcxsq2P6yLOg1w9a5QiUIUUwBcyCORwgUICbeoqU
/iofqkQ5ov0E+FF7yHePDK8kA81Mttpvok6KjrOkM/rHbz8chkjhQ9tpKNCqsi6z
ADD9mDTNW5leIvbOiH3fNcQaa2Fp8V5tiHIlOwpYaqLQI578ZYPGvW46ymHT2dqd
AASNcQelQYSgl5aq8VISLZAuy5/6J5qXFYhyl22Cfhw3ud9x3YFcy9a88moyzja6
tOHXtNDkiK8qELql2DUZHKm0NrzaPIKaKSljcFzrauY2kZX6MJxvLjD4T7wuG/eS
YLvU67FlfrGKNLT2qTCqO0SUvQTwgd2BiW7x6c7h8Vr3ESzI1zS7fb3yAYDG5ugw
Nav+lXjJbVo8uvkmmkbfxvT+e4b9dwOCRapQKgTHwRqjdJ9WyBeM7ApVPm57nOGf
7fOGiMNJWmAzqxVUR3zhtO6OJEHFSCTO7uFN41T/nWbGxon1fz1bVGBR0Z/Njau9
pLjJXpVpZnBeTRvRQvkxn9SO1+j9lGPjLwJmic0TRsc8r6ag11uEF1tOv8GIpDkl
omqqWNXGlk7g/xXNgfCvyRA/KNZYazMgpRihK+Fs7h1bPAYNIoHscsUtFAS9EpYS
DKwBrWrIsdO8dHJRZA0Lpw/dJVILnr2FL9byMgGcIsGbR1QwQgasEvmoKzDEL+Cd
CGabo2ah1d3mzpG1T26JCafEMndBYxRb9wpuJ3y3TKBEd/BQRXtP9nVMlsXRmrhA
07vnQ0qXhLEEGo8hce6K3d6jk6GStaO0HdoOYKI3NU6/rZ4jxJ33kfI6AwI2+Amw
HbW8V+NFLc86vD6molVb1D5dMsKLOqiWGnx0qSScccoPzhK2g9nhsdYaofmsOuX2
g78GWjdW2ShyCU+4PsOIhUGOTFJihGQS7afxLVyFUdqpixvuORFRReatBigtOo28
ex1oHYtGl/vMUHdJGo0vYibZTfCDvkGCOtsZ5sr9AT8SSJAzwsiIJMip9pEqKpNt
IMBKA0snKmwa1ozeelCiGgKqD9PIfotC90gWMLH4WCj34m7EOyoGWttJWAYKgmd2
F7/bylwfRCqZPnCB2oaGWS1ZIq93BC7gtOYpKq/s+91OhF8BdvLsBhE88yV5Pv+G
xv+AW/jKux89Bw5guYHCybZfXbPq8HjjdIfmOChECNoZIXNY/L5ItO8T89SIkBvK
ZVjJ+LaZC2LkgiCw688YYreRqk0rJ4YzbFOtc25WUqMln+iaBnIU18SQL0VEve92
v5uV/jFblC2aoYvJh+FQDCvpkH8PUUvww5Xv/s5gb1SXPtDKdUEKwju68snQGAoF
9yDVUE66czr1dG4VwVLm2Z6RH8tSrd6ZrMA00k0qjfd7V0vlbgNu6Nb3Ctgf0CAN
gbB/758vDjl6IpqINOlUMqmhChgy/9ZdaSMUoCcvqDtOjgGTFCIQfZdWz//ed78k
3l+TL0QOm7cTqRaqRVeUiUSLoNJ7sgJD2Sx/h0KwZ5sSvYO8cru8kU/mafkaDrLj
fRMiD9h/wmsQElZz/JH/v//QzQphB8FNW60tQ/pYodqe38sCwD9r8p1F0X43P0Zw
8lRIcQ2Bs008eCj1ndUtdaVV+7j8JrXQaIn1V58CvyCvMj06bgIQWGYRJlvzaJsq
2sWKwQ6Y1QOrZwrqpvI5HNxN9wbKDEIDF4rySy5B5b5tWLmyHsALAckLBBJlRgAH
VNLA9gTa2AgBOXd4tzW0KJJxtdesX3i4kbne52f1kL1BwZMZHM8uwDxdY8uSqnGN
9wmDn4F4g2mnSvbAXw4bDqulTH6Gkly4MrOaAvMXRphwT8VFEC++9///HMXQ+OIR
cphQSnwlfNjvukpj0cas7tGkM9L+F/1iAItiUBNdcp7v8jwjXPxwk9gXCLPiLBn5
KF/2OkCNxpZXsGO3VCYo4Mtn93PM8zzpVTaOqB/QbVWmVe0oRytCXJNvLJLBj1kr
XD1bIx/IcKGQKeruU2Pvft7jL9B/T3IKRfmnFLv3hbqZy2g9kgp4BpkKWq+JUKg6
ItbfPfc3Jjeeryzm4l2TkPAAVdgTlX/e2ZM0p/XCPdX/1l8MmTpGveTJrDaqSdcE
dZGq2ZDObndl/uQY6IXWYMoCUNPXf/S//kUCvbCPXudfJ5tqjXU9yeUoA1ccB6yU
WL42hxwcUFrC5xv84eLNaTsQMkSUMQjVFfIKQkY/2GIPrqA8UI0kEvtLjCt27gzo
yxoDMNX4MI/KqzfHYhUzwEsPhT9DvFLKDyNWsVkJ4eu6x+ULlRrsCJRDZ2XsjY9F
VTqY6odh6dKPUYrJCgnboLnHW5zDbE7usm12i1Ysvx1+tAMSm5KTaqgp+IR4FbLR
57VbpMSKpYpze7eK4+50Hu795PI1M7AivOv7w2dHtjVNR3jPIf4mXmu/vpcXK00C
zR5D1ihI5prd6WBEly8Oveh6MP6x73kkwevvpF23EzHqgZb07o53f3UD5O56l1UE
h9JH/p6HoxrxN8kxCiG4k6cxCiTajUdLi3ROxlrLDKFbuGKhjCKrnt6NZp3vc37l
febOf+ZqimJF4eYJw0RhJwCeDs3fRX20EgIoA7TLrWHtGIv2FYw94P3ta9WzzE3S
lMBLVvd88DbR9d67HGlxzHMAs/Z9e3t1JoB01Yg4TVstJ10lK1+CNmI0MiFjo7AE
3rJ+WzUQXpv0kFP7u9pV48KSIX4vyEhZICwzCwlA/vOWtgwpDpfozG26g9ekOCA7
R2MX2Hi9R+QK0cVksLdFOqNoiKWuoPdqGx78mXC18VqjceM+2BFtl0IAFRZ3hIgb
K44e//tQ5SCjqS6qyPRzQpqnGkogChdlKpm546WpAvzAxf24uGdcoiwzcvfaFT7l
SUjzeE8oQ/63mPYuUX8IinNYvTfqKKNrLK8WuPbzpRLu5EWF5ik87XTeb7E/1uUQ
GlCu5tZTNf7A4sIgioqqlmEnuUlgK1F4s3rdJrttRG+jvTgvRIK2W3TzzPMvnkdl
oUhS/uc/J8BR1Gz6O/KRbvewiL42yg6Nc4tWsAXOvt0SPtbZRsBhgv2JiR+CfRGt
gocrPlpOzDrZ/pdBP9IFFyNOAbh+YwKAl+xK6+8XysWGSqdMDTSLBA1vTsNZAvZd
1VewLLon+tBkHumuSGCAM1/PQyKcsx+hK2cJu6kQYYiVedhJSEdM2ozyGl6VdmYa
Wd4MoZDGdpfKJC35NaKIdXzUQ7AMyFDW/mLGmxrNvR/+avXwf0iXUfIz+GUh6e/t
IrxgumTc25MEvDHPAU5lKwQXpcZ3OWOgAho5YHdE6fa8P/rB27x1MXzpyk0JGKLE
eD4anc85tvEOkyfP4jb07GLof4KGo3Qx1hovNVnwu0hbBFkHdTIXdzihbRR37BTe
j4OURGUB4wgR1AtKyaihrMAKlymjxXXOxgS0Se8BLY4VFtpekX/wWpjowz7vMD9f
3ihPp+fyUo8nygPjVXc0YoUvrOs+qFa3lyGo/tbCBwApAKsYLQP20aftDWs64x1O
WqdjMFL+9Ax5mbjnEZNdte6LfFi6cV4eW/aHj8BMZZSSuMxga4cus6UKg3TlIkLB
cyPxtSH5lSRExsyv/bKul4hOZN89MY0Qg3dRdTPrFUrKClPSL3efcC6J2ElYvtNf
IWmz3ZYX2vE+uBj7dBR1XUfRfXMAWInjs1nBmex5xDFgbAlh2+0ZxVKsNCvmq5IU
j5jQjCCHlDZhPhfp9N06JNigiZXK0WHO02RJ4XsNjtwdkWh/ozYN6xk1RYpge0TK
9B2lalVJk+e2siUk5tyUe+0j5h4gpFXHBSnuGDAXRxLQM5XF5v9EAsOxkHkOcCD9
n0alwS7cRm+9CNtclUf+tRPzMjEST0FTsqbgbxQvrofvGlLurDv6Tnf4HxGmGK+t
r+FzFcL8ZYFLudjYvldWqvz8HIHTr4UcuSpQmSNdgPTKG91R1oPZHWDV5JlGKh4V
HEQImLhmKfVHriplvoI6dWQKPn7iOG91riI2uUQoj31jogS3m2vJlWkYAJDdLoW+
6iXEYVCBZXhVR6qZm+1z+KZ46NBm3sAqo6mWWEpIXFpOJm/B00SGcOKy5GYbxV77
o2kEdHKLM3IGdzZY931xk56du9TI4YMQjtDlRXtCLwvhbT1rCgRFxm/7J0B6lzU3
9n93aj9B7KD4j7rAW56MfdvUuPzaUL+H5KFFy8nGSThxHLI4+R5d9a3Pxr5o9N2d
fLr0rxDt1maob7Cz+XUUv97W3Dl4a+xKYUeTdDdA480hqCVpg9jDzrM3QxdgGjSo
bZg4G/EP7JaUvm2LBPJt9OCqrM1ZO4DCJI7DplEPKaBz/eEKIa38iBQPxLNKGa4G
UNg+uZDeuuDaY/lSuBhP1SbQZwDDtHKc+NdkxXnKItus52+4AmCAJbjMTasMrnEs
WoW1TiLrEIUPw55MJPIoR/XQFhUY+Mw/91OOj+oFQPzuGrMlyOCSwTCsariqCukA
yJ3544w8RwECLJM7x3PJbq7969iHbgT8CYiirxH8YmTyCCJ/taOBAB/qpRZWQRnA
KjFz6gAzvTfxHSS7BgceqQB57CV30nmyYKENGBUUw3a+99dsWrisrE3AkSZ/ZsSr
pgZ2dKnX67zCb9Ea/0eywkrV5MssTbT7adOxBhVTPxn1bx5yhPq82MXLmKBWBqZ7
aMvRU/Fb0/d52rO8kZOm6u6eYsCN5+HZubw16d8fu9Z6JA4Mt1xMT4mtzmc2euZE
9GcgKvFN/NjxuCmR8vKL2FbphPZ3TRPFCr6oYD/euthU7GESY0/NwiAgscQ5cG9V
uzB7ejkuTO6FogO+5StQr/3p35bhvSwJSJIUjMLZOoVNP2HgtMyKAV6QS97kOHxN
GQ54fWvnTPkmjU7c+FU+iCmxdQARlpbzModCtDpwWIBNHYIdC3lfU/2aiRp5nXDC
7VrsWieizSvDXD29lGXwKiU6kpCWjS9uzq20xgvftO1IE27qZBpKJH2qtyftDRkT
+Zdlowr9Px9s12wpx/HV4/amdikjxHj2RvjUDA/OODVUDfqPGK3UyGWEgQFj5SgW
i0g49rsQ+oYgnNhixTnq9yBbD2zwtRBey/VpPcRVU8LFb/VW3xT5DVnglrTBb5RU
7tlJttbjk3ssd8AfV17+Ca01VpYrQi4m5ev8HTBEYoM1GZfmUmx4ygllxYtEbGzU
fYrLyZlBJKgZT4ncmYYsz4PMyeMIfbLw8bntyyd7Hll8qbPz0YDFbZXD1xCiispM
YUOxuHq/5oSLD56fvHLhD+KTSauqyKOuZPnHz/KOVwrUUBJgsCOZVuhc4MWJ9hMm
wotxxNVuq3MkpgaxiTUZqoWMDD9tX1vqwzAT51eR50jyoeOiVavk9hZk8dh1GCuo
yU9V/cU1HMp0s+kqLCmFPKL/+UpBYHhh3OZLPjoJ3SOtPyhaJ+9h1u94RdThWYFD
y6q9/HbU/6BnnvwF7Z8/rdErRI6Mhjjmj/6olVrjBWRcE6MWLY3hFYHU6Pet3x1v
Cnuf0uWU1Vwt0Yqj43EO/tlyWC8pOgWU0vETEKOshmWFLjeE+I7zkQS8DeUL+QmQ
nuLBpblTaJppqTNdvgttDeYz+71y8/W02GvE2EksMcNjW2h2bdberTCMFhlCMUiP
TE30UzY39LHixWF+aJ+AmBYRU1v8U2IIap0TLN4B18yAdLJO3z3Mxt9Ksov1wQSx
6HnzCGUgTNH1AR9fU2wnt+OpvhwuKxZj1fEs1l4W81BtobCtCQidxi7RPi8Rayo9
Lm57iZVCQSmEDLOHxWTktaE5RlaP0VyJhL9591JFeuGb2NmBgszUeL9Tgi1LJa29
r+/FnV4Hv7RG/ACdVTTnv2zsQIsKxmG+Ny28a//Z3ZGnTvBTIJHFXubiGWGH8KNp
w1wmgaVJaWndZiR40aHNzvMEag/j/DlbTIYwAwHbsvTqgTsEce6AdvXdlXsdrho0
twsGU8SJdRpMIa3z2lxtqzib1glDN4uG3IfVppZ9Jd46oDntwKBtzlxFEu4ug1Sf
om9Y/bEE9j2iMiw4JnwToJ03SSLi93EwsTmYbNyayUPNYU7Wv4CiY/HYaG2TEzm5
CH6hTK0RsPI0b0Rh4kewTIDGBKyb/mVNRGv2d71+c/QNvp3pWxcGaxNNyCe3XtDE
j8Vj+7k7XYgvBl0aBmIg9xPLBafgyIP4BWNlzfWG1A+8K/EYBLTVXRrqVZkJQm0o
yMeAagBFJR15OZ1r4nQXvJ+A6UJniCKtl6zOyeOlrO0lAwMyQ3eJUQghmfx8yHhU
IXCkDsV+blQ9+Cq/v+DjeLiBBYcOa2h0CtLVWsReSk57FVJ9U2sAFZ0JO8fdjDTe
oqL4eBTynft8cWNxobE958swZUUL6r/BF6x8qdijCrwLISHPiQKrtkcNJFyFb8XV
U36Rei9n+UDV4J3XVhpsX4z/KUBpSbBsne3vZ7tnxLpgxHpxse/Yj3nWWJNiNTLI
/TN1cULy+F+y4vYAC/4xcRynQ6gJBRE/IkRBkDzMIs4xG8FznP/ROB4jAousuh3p
wTDOeNjPjNZ8fCUPT8fT641ixb45lDxpiZikWZHdRLPhC8ma3LNyOMnBnMDW0pKv
slkpD6ZnjgT5jbb5RQii4nkPgGrOFYenLFUII4GWCpdS08nMrP/gv/Z5BWx23Sry
cwXmbm+O7VoaLmy8q/rIbcxCHUNF9kD6QGuzET5RNm5onytnImMRSTHRdVbBiNhC
lgVC+VH/emKQ+Z9sIPrH+wi7cRntxwyl1k0Zq5PlVlieBkVSB2uGpwTxTKCW/M1G
+OalHvDfOjSYc43g+jXSk9hrNq7A4uWsdurq6xAf/LZFw7YPdDzo2HrSwcf/iggg
MgFJ2YvJOFDCyStaOyQtQ2uX+L1Zho5R1cYTML9oQJKBiXPhiUpE91MJr/Hvef72
Cnv2hwlShoZPwXNqEGg2UCPK+g6R5GbaPhyJtR4XDe5cQGItDhPH/xvXfgF3oDms
OaKG6lHh6rTtjItcXpjIjyl9uXKasS6vxpIIXhXOECNMdkfE2Mim+FSClsYUW6tP
ygyn/D1AbO2WKdrjp3dYHxnc0ipagsDfWLYJb+ZSK6EqCrjmwKkYBFNOmfwkMLlp
yDh0Q5mfYMH5KUbN4TKa/nNTr3it4xBK78z0OcQB2q5pqZ6HOwP8ayEuy1YJi5Qr
gN1XkTO9TxH4pzrw3c/Nb3aFFfzlSgW2fgenngJaWJkXI7jGTZE4nwaqj08UEm+7
DwTIWmZ+3JJ5hbodlSbniHmcvV63ab8xxN87mGB4LkWIKQGRH3C510ZV8OtW/vja
I+8QNHPvpn+VmJS0FubLepLGMRHIFhx4ZIq2aQ4Llevg7GjMYtWag7qCpRjv26KH
qG04UYD49YnDdJ8CsjqhFmg/lNndfirRjofPIHImHC4HKQGCOQO1AlPyAe6UftoX
LDQWDlhBitX724DjZ6IGPHgykjZ4BU23u1S9F4sJzKQ+O77/E65ErGfp35LIL4U8
q4XWdG1uTSGFxo655Q3g4uQc08VtdVJ8ZiSkgj8Go+MHxcfdaOw1/rFw2DrcpDKW
uMUNZhC24PbbfUaZmY3YctSTuEQq9vwWXWJCkryum+wEMDUkLBqLqiLutTRL0Y/q
irLd1pRHrKxUy4axIEjcHKR268dpxphs9B99OoRuQsjvd8XL5VqZIbavmL01IieB
+JP50h0jI3+pfbE14Go/ZHMogZm0FrFjX/MU4HuroR+R6nsuciNOHw0rguP5QQri
ij+oWGOSJPkMAy6A11Po7mEiyAvVejhhMgfJbW4P425q6bXLbi7xVeJgrhypTNoM
wVFs/jHkoDDD5hdF3XGgLxmlZJKKCnC70TdvKJ3fKSu82uQTPFmjqKd9/es0VOFf
ivymBzQPUPk2GBYi9MnI2tHYmukCXQMRHgN/U3aX/rTqAFKn6iEhBJAZxOxb3Vam
f/SWGFwODx4b2Paq26a8Znq4zJJ2X8Etef3iKtOJxiEJjiy/VWycsaBJU8Rt3bTa
qTtVet4d0KdO3DdHN2hhTsHK2/rZJ7pCDWwBjFg6xvdEfca0VRC+wgqdRLBqoksZ
zYShP4Q5IcW+67hxEzAbiuFPh7ZAbGOe7GU5wiURo1IuWSGuwlLj4UPv9a3yPl6H
YphTdkZ2iYKDYJ1IjgK3vikG4TU2PD5XrGItcEPnjhEn1Hm8STETBMbu0zIJRnUR
yyn1/kKj2WucbtG+wgptSrS/GkJl0jQY3tfI6N7MSI4yAuMMgEL5beLkx/dMTU8P
FfkuSy0okCPqr6E4wyac49M7YhrJVzXC5U/XbxZ/2+BTbds8GfNGaQPen5XhnW/d
DkBVvsLvsd8PDPAtDT5cJUppX6iYAsZeiCmPCVdgV0gTcC6TtMSIGTMRpzsG/27n
RSb7bEpM+touq0htQzS7K0uZFOyhgKkaGH8IOrk1cQouiTnphO3LuLUPeIyepYUc
JQE3twy5LhgzHp54mvKbUbGogwdvvgbfiiAMBaNVwvFkYgbzPJXFL2wUyYE5lbr8
bz818Js3JIVctdLa6our7CCX8awb5+rlpU61aWhdKZSQgRWqUs9CL7ljMO3st5wr
uumlQzKYs8wjB+r0mShwIPmIPjt88GtgcpT4AcvsYr+0v2eD71rx24414uq2EobD
gZMNvsgibIGN8H7Wh8vXUY7k4kM/+MzUHr0iVkKP6XOKg2OWiRPcfY1n0sXzicLY
oheR7y0SnXiQNytZsCGHJs9M9atHt60K0LeLMBJ1fRVPIcfcmQ9OAQdhefgZ6nSG
jk0YST5w+LU3CDvrfICw/bM7mukYDNypZqT8Z2kgGabO2BtOtLrGqdOGuvuKRkyt
6BQrGHCqQdYAEqJFQa9xTdKe6/bBVizOmqYvZjA9jCQR3zPN6Kld2KeUMliXp8pe
ktsyxspmQY5iRTLMpIw/ATYl55BdbXu0ag8WoEJRGUmh2Z3LXpqaMSut2Z1mcPVf
ju7n5SsJ1NgJtBvzCuGPrm2q2ANYz0HwlruLQpxKQ90SIfk3hUCK3T/gcnmzEXDl
NtNOGJDBSVcnmlq/98ZS23glkfN1x3TwrjnCspUxGwDmlIoXECrZFpwQZbE3et3p
WGgzW2I+6vT2mB+CxiLkR/+83pArb1SrxramC4+LZfg8nBh6b5udS53gAO5DL2JU
d9i8VqvwxPMWY/E3kKjUMNngfJf83wMW3u80Qw2ZCBvNN274aBpc5IZ1sAGXm0Ev
PM7T1IvwV70A8YhbgNZNnbkCyZ85iCm2wvJYHcg8lTp8+b9/V3exgY0mjS4ZMmHx
MieujRApfgMXw3uq4K6xOGKu2fnF6HHYpPZCyI4dNdhjd2R0q2buNOfeGneHakte
zcXMOwmUDjdr0FOzJqfbFpy0g2l0kAqLWtgTwdHj++FvhtnSMy2qRCZv2rCfaL1s
f9/igWoCeIw2GdldI4SrECfOmEbKZYqYYAS9c8baM0SY3GVFwxBQtEx5RPFl4o3z
y2jFStqUOIMajz2NlPWAeODv3VJm919xliOZoXnCgWb05cLR/oa+qgdvYt8pI18p
/lWjhH7gBMXMSihTVzb8LceLdvKd1Et/7CdFeMit/Pu9jQ1ek5X49YSdEjZd1jhG
nilUUtjNbf3n9dSIY0Uh1EKI0FTYLlUQX5fdG8OJXnCjghsLvGG2chCNISoFhcI4
eQdU9T/Fbzp/t5mlYIfQQR1jDP3/2p/VThL1dQ+dsy1mPyCaNO+aU3RrlG8ti8Ea
m21nZ6WJ9sceNn5UuyfarihSePK0C2dHbT/j8Mu4XjfkuAYPXj+spPzrEwcH4zMC
WoWFtIPHylBqKpFdLOUodXbzrj+RUfwINrUbN2X+BA7VdvlT3SpzbB8GG3mqxtEs
S8bTyDUUodCSBVfHEF5bFHzNYjCgJngYI8RaHKVjRqYcYSueyZ6hYC0e6AcC4W6K
v9UTq4TwI4DFxDtm9b+6bvWja+dj/kfV9Hnijsli5v9VVTuojgV/iL+pQI/cB1N7
RMupHJNM8BgNI9FnTjzMTzex/GETP/fXXCShrp6w8hOioEWb6frl+/Zi47KWGaxX
Rkqhq2kwQyxGA2hnxH9QpNAnc6Fy0UsfuXe4kihevgkWNPBahOs48cLy4GR9VnmW
ElaFbod6YmMMsrGUp8k6hAZ+OcyyI2/ylKEg0CiYlSpgKIaRd0ns8s+WH+/eoK+D
xt8RTQh8JV99jhWOYe6pe7wtT5793RYnsjrrNyORMPVHLx4wlPOGZB6ToAD/ZB+U
LmmXlagt5zGOmEPwK7683VPHe2bG7k7Zps5vapQdK2UW+ERa1F31S5yZ/deZNQub
2T4Z2XkBXVoM+9q1EWbPgCLsApVlkwFz9XiZns7c9HxoXwAzBiEfnKJFbi2au38c
b9poD9cnI2J1/zWM4PDU8wMwgcZDq5Ii4fBvhNXiv5q1JQ2Q98kfSQTUSOrIFPJB
Ctm2U7vmrYeRrIJMB6kyOW3PdRhrLo05rwx/rUsQIlIT/c5qoc5cif0JCnNnm5Eu
8VBo2t7gsz5sefPromxAXeLkf9XPYcUJ639kxlcs9nvrx5N86uw20rUIQT/Uic8x
CUf3q01L5oCRbuHtWQSY2jbLR+3BaTp9erkSy0npQLrIAiiwxq0dpkhTo9dP0Vvz
BZhQV6hAQTdoKVpfNqH51n4lxOPCIkMoxc0o18mwzPalCbY9GUt7DrDFvLxEO3/O
hYFaTRpKEX9A3qNXWJBzRUxGmyFOQmnSxNs4G4kJC9eHWRStClGAQgaHO9vGBCL/
PWtVQu72dzV1CG++lqBUmqAGVH/5pRQfhBzUULdKdv4dr0/+f16l1QdSHNxOJ1ka
yl71kVuubyAHhw/8XSWTFSBI9Nz5hoW/MWTXape55x9an2HM5zNXoJ/ZMsjK7JJH
521Wg9VlQOQsVDAggZHKUHx4zbO78ZLtjD3CbJz4kDD7VBFyYpF1bXKLCP/TPtv3
kwMWF2TVPi+S2Am3FVrJ/N6WpPcDBB/GwoL1+mALhtPhgbAPHT5a+E3kFc8T8Qut
hkpt6j8wQ3XaBqbz64EL/enN14e4s4P5Nivg8KxsvqSvIjT6Ayz/2UBaJ4G2oawi
p0xPhdVm0NuRVDKgMvdyyyoHdebWQz6djCcAf8mTFAS/z6xpZhC0TnDFGCJzBmHy
d33Q6h+CLEuQH/POMDkBklWCxz6dlSYnK6JPd41o+VFHcBZc4xQnnBJLtf6yu1Dq
g9ZOkeUrmpksEf3PAj/PhUoZy3vdrIfEoQzCrVNIy0/WO14TuicgIQJboMYgUIYd
0O8ziliOKSG1vclXGXHEB2H7zzwasW+t4WdiHuzTwwqpRDr59OnECKJm8K086r/k
sMStGvmREXpsCxlqjv7BjYAfmQ9uSDgzgyWlZzgiPSYZvALEgk8sT2fdo4GChrmI
4z+eN4iGYdDr1J1gffjb9ZJHIM0veyhv/oxtJQ+zo8LEcIfqzftvEvLPyQ6nrefZ
e3p44/xJ419u/vODX61F10Z/dZw3GIVawtGsRVuVH1kwbBGy/gUYyXaZYEOOi4BO
bwBBFtqwoglTc2oZneSI5X6Kl8Vjl6OGjswzxLHobXytrNM7NVCGhEoAP0TF/Apg
nDY54Oa+3y14G/gSzD/AM3nBLDWhUfbx3fHR+00qzSNlyxpyvHHqPPNXx3s29oPc
nhaqMuhPWxwQd9BoELwM538GDAQ/EkKyujQsEsaPcKuBirvLFdvmWge8c2GyuIYI
rgqEnSvUyy9smGu/OTvvwxasZjQIly2Q6fXh008heM3YAMXS+T67hhRwxYOtTEZm
EW2jmWL+UQeucUBUrDAGEJKXv6L+8l0C0oERsDI8LZLj/fsdOR0O2ZclI6Z8tOrW
DNAimw404eYD9VwSUOERVEjsEl5xx1oUTpjwunw4AK/XLps4FXKnbeoXTC0sJaqn
17dpCi9OBZGS1ybLKvIeSQiAcuDJqMo1bOfPNixzwt+i3HzNqggW+BqPHSO/zukb
yOyFfXKSR4bdfTUmuya+2PBCVmvTp9FFbKTzZveyqDIOAPtccL5InSXSUtXodbgn
9reaxSRKDqJ9H/mq7ki1rGAIqoKXrbQpljVpbR672CW9FGaN0GObXdPZABok/HM7
7yu9L0lUvjwz5rrJOUfiEUe7CPIiiQFlkZroWoHbOTTNrKCedL3DoLn9Z2CHkrIB
+i63ts5bIf1c0LvhqFaOv7ZoPrhQcg4loyAM9PvUy/d3YR0hPAf9SVyte4KlAdNg
GocL4/ITfv7epv6i6IVJfeOABWsMdqQVQI/qUgD3BFpCvU45lnh22x+2pQQ/1vwt
/zZHB5MKhXsn1ot9JZy3kcHXnq/Dp9qDQ3/qFl8KihJ2wey4wKtnedL5HwrQejC0
upjVoyE6ZVgqeHHeheQqquni4gwpxkzUa6/BU/tmMJURnyfjytZcSsjewwOUCxCz
5at6SaClWeUUB7/OQ5OWsVgyyygtWeu3RD2NbysnGhWifTown9ns79HPzw29s/NI
RjVnw4F+C8Aob3i0jjPF/AGfvnTJhFFFiUwF2RgbqByBqcUliwGublGgv71I0Got
pmsu/RrTxg2pmvhnL6bdVddzwJKPWj47uiQ+S8wXEdaEjxypldRlsE6XX6dEbOF/
59Imsrv9anBB5yrL8/vPOTU34NdlemMbHi1ihaZFdYNnXqIx2Um0sGlkWtJkfvdT
eLuQThwEMMkhf7wxO17jfrK+t7H6LfwZg5IAg0HoUVNz/tu25BW/bthI7HFQRKkL
f/H3w8lTLHJBsVYZBy3B2lVerUSAyH/YSE1zeQ8P8x64yMQMPcYzQJBrUIDteD/v
Io5lIFFWWiI5L4qvztP6tFdNs5dIk8VaEpyJEMmNBKx6nF3wOfEoYqEPeeZz3HQS
AyJy2HbUBP1yAjGbl/7GyIRy6PT1ynq+yEWvhXGBgkmWeCdSUpzw/9QYivMDqDs5
AsqYSsVX+/KnI/HtilnJE6L+a1p4NoBoeokodLlq3ZMK/+2wvTrhCXJIEfGK6lxB
kO7CCG84yEww598hGjBUP9NDnx9ZlMnbt1PR7pxZUXuNZw5SRS8C65+hEIJbM42G
ab9hNnq818HcO3LoqTGw4Cw3JGxtfk/uOOKQS+QWd5WnkqtlOehcSJLJk0dvo7D9
vQiCiGLdnbvZwwuz8ypksQFDOqPqaDKiowExuaWVW4YBhcN7iMsqrxm2OJQR5H0g
1iHrgpvzOSza7FkMpsj0R6oVB0g4igCniBWekmdVT4lztVnvGzgRHjp68HHDsaGW
TYT3UVaOkElRNEhf1+nmPMQJXcRHcjaU71msRHZrkOhR0kh9t8mchiO+HbiGJaaG
ZyiGuQPL32wp3nzEzq67C4gxgduv1uRUKS48BE7LYnB3TRbjxzIJLQV2uwofvwMC
ALMQoMDdXrTu6RkiVbX2Cu3wXrSVE22jFAXm97iRQ8hNsckdwJ7kApDal2b8VDWi
pvqpz5+HpMzFDFJiiu4b9T2rFscibFFzlnXOP73hDn7uqUcz1qPzM4kElBKOGz+2
42RICqjhduzunoNyas4dvb6kHRx/CjpSK9MhSiP60Z3EfVIA3XJ+5rUzdhEiDlKa
BH1zh3NZVS0CiMwFNcl54CPkYXx9spzCI6wZmcWUwc2kRSxpy4myZFGvq1WCCQKl
5Ex8pzkvxDYQmORPuhRC7sOExIIi0iO6F4fQHtpD+J5xbfAP9hXF6WQldao30aup
S0fg+cuo6gt2cyb5N2PPp24pfU0IevFNcYacyyOp6fC0zr1hPsqIaSiEgKYTRokl
CDLfrCKi/Qchpf2mxpjxJBUEWprYzCcthCxmWzkDHhag7DC6GdyNLlNWN4lqz6vk
uMcAHSM5UHJw4jUrt5kl5woj+SGjlerOlCKe1kqwTCJtIb9pO63xeGJcjljZRqzj
CKPeQkKR5tMWWuN8fSQVY4LZ7hmvbYvdBhaGuLanCa0lLui/a+K788EZU9ad38rw
HPKFrni4smAg5oVgGNzbHWl5yvEyi/4stKxazOm/XHDHZ8hpffpiFX3SIaGOmY5c
4HUp1Uk7RZGIOwyDbVyaiDD8A5h8t29JWXGpPHshJu68t1GkInq2xhk1/peXUhlC
osIH7OeGJd+uAK27DG4nZ/nYGOfs9GK+6AahaPbc+zL56KdLQxrawaaA+ndaGi7p
soM1W/Gh1ObDn3Fhh7a62p53+maxHbQ95dcfAWxCzLrFRfLxs64nTYicuPEV6g4W
pO46L6INtbnudjzVbXrPm4a6Gx/DCbSWn0uMpfjucES5ZDGMjjFnwHoyKGtmz1CM
Zv2FEUYmbqA0tGLKuOgBREq3hYv4lNXYEM9ibj48+k6Nv5TQxMKg12+sjQM6FZ/8
IscX0UMeUeY/KbaCMf1w+SQi0o+oD6+tQ+4sxVi9Bi8Nd6sHu30EZ76euRlYNrPO
SR2TdHacX3JBr1Cj/lwTuqV+pHdwsMaL02ArCeM5XNmjL8t1CAaSMflfonm8fa1b
YzPxqWOFf2Kr5ReDymFMvPXbz8PIwYIcYbKwSqr6Y+RXmArHsxVvpmVrgksZuBeR
69fS9dJSWaoaWC0PqKaGQkOD3SrNujkK4dS4MZlSJEOZ4PqSdkXGupx1waNyjI+r
StFOMyTkMqa7ZpO70wwd2JlgIwZbAU1WgqdCt2ui2dwWQiFX8bkQgSwEgfKtMXZR
vIE3YlZZRdaJu/J6+Dk/03D6qzAgomxeqFezOEmaIJ3K4a9sG47PuiWgTNSFm8C3
a01JZDD7Wbx5OdGSJ4e2V6yyIPUqT0Rooe+O6+qUhygW2LOcPHqncVmC+oRGtE0T
+HedIn0hYDnj3qzZ9G4zKIhIMLedzHsAFwIRgp48PdydHCHP1HmZ8pc3Se8kvStd
nuEGOD63JGV3aIdEJLAnxs4exOBzwLMndtj6QUeDd/XIQr3pxC3R9DTOA5fsJ5TD
LMWQdaPeV2XjvWS3WyV22AXMwVKnOzCRUwqtxUa4PJMGuMFb98GrePzN3/Yo2X3k
DHJmbPvRQ2cvWE6m4KPYzpcnSjNDXWA+c7QPwwfyA6Tc0V6e77gJ7lLGnhpg294t
g19QLZUiEMUYrzFEwuU85vH5XeWvokZR1fTzCOqP3WniE4TLT5Xz1H+xHWmlgJrb
6AhsRw/EzdiJ10+9+dc1q2EdO/ZKyrzAzr7kYJcYU0FKE0kpqQo9NxCDf02H+E4P
q/VUyi75lO4wuknH0MemOiIWCspN5BB3sy3mN7raQ81Jr4ZRVeKtUgOw023Vlter
oTEIbq8dmkcZWsuQGF5+ZdHmBZkUIE0sIQG1m6tiWZ03Weeq5v6GAjJcMIP/gNQX
RhLB0+Q8JoxEfd2qeRWceF2+bu6owop4YkUWKBDapJySVtJHj76yC0zcyKV64iim
0hLiTtHXbS7Vw3ODbqNxhmcibXhDI6qfJfqeNWm5WqDpa3jGynF+FYMWv5AvS1Nf
7UgOjooqwptzGmGweZz7hX/NMnQDVENTTasLtt6VzX0HVBk+k7pBfNl9OCieKCeF
mVdNua8AMwJB6KPIg/jIyjiUe/BvPo33HcKr3dhPZo7MFIcl4gHn6Bx83AKBszQ9
9F0VaminN5z71xdFQHZWtTtn4TTtAFrbw2JwIvow7cMLdrkGBGp4O6+HR+hFhSKP
iUJKb5jlPgasebYJw7NInU6QFzs+9qOhV4vGOtNMmEObA94QzXqlNJumSY7GVtMn
zuXi8RWKGI+FfXhMZVe3sOWs1VAyBhNrdQaYn23NwIwQYD52hnrBXBhzdx8xLI2A
BZHSvoiIQNr2Gx6bgpD3h7iDL5Oi5Wsn7OCjjr6/iaOSieextMKR/znALLNkV2Ov
dsmWLmD9BV65A9yHfte/X2WFjfA+sU49IvFyyOnGKsCvC7+Q11VpChkScDNkJ6oH
xNwREGFyK4xA6cBae7FbH4FvNxDTbJ03JMCXBBJ10+WKgpcPQ1GdGkpkWJxEuCwP
K8bc2q92lumuVB5beVc086ZVM0zbWFsMTy15lqMyQPbUknHNp+/Xr4S+UdJA9wnl
kQGbzYRcEXzdugg+z6xQsA794Noc98tU6EhtKhFoml0anI9lFYhYI+j8sMoYMoDt
7PmSlY/KaW8rFNqBQVckINybt3qLcRgXQpkqCYjvT61CqpL3xdjXY2RdIu78TFz7
jDslhyK+1Epwrnq2w9z9Wlf283J9XKwYI9fMQN1nXzv1/UNNuTXgFSnM2JmelT3N
Hn2Y0hrxtJvJw54+8W9A+qGrylekwMEroqYRp0YS/MLVO26GvpeODkxin/1GvQul
ix7FTu6Z5523IMrtwFU5Wv3kOt6+MJJ2PBrGjyJ77BSWLD+8t+maPlsG1GSjSK89
FvOqxEWnkrTtN5yPt8/YrVw59TIYhKnS1gikZOLrSbkcp+47YhnsbDoV+Z/Jr4d5
6qhwht+weGxkbqWrNoI4DvbdYCUPC0tAPM+WgxR+9pSBoG2/y6hELL0VI7YLIGM7
hs+knbsE4mY7Hq4OHhpVq9z+YJR2h37SBgDa1ZXHpTeR5nTakeLu0Rzn/AzepYS6
3wKECizFzIJmCcQvNLVy+WPUNKXWGofP0sZn+g6Ld8u0fXgmvseMTglhXgO5WPnL
ujtpzRbWUsINByPky1/RepfIWaG1AM7aXw2qY9Gufu0mGTOZ8sATcIueyy05s52k
cdYzU/DMEdUAR53eHMeaRTcQNgWy/162ob8znzWE3b/MufEf/g4sphJE/tOnTWT+
f1Ztl9coWfv4hOlgDOJAx6jgY1XHGRaEQ438Wlz1sCtgJf5PV5WLK84ZOw/2L2iJ
JwV/Iqpj6jMZRq3O/9SMKFEO2vVlVcNrR1gS39GZDWgIVu51I4Bd2/bCM8SxmP+2
4lHU8RU1ocBxrBVeF9jBf9B6MYl8uZlSm832hgkJxlZf0gk46Q/6X51/4jxIcUSY
8jaIsQjKpi2XE9UhbmELfqjndG1d5zoh3+Zo63icXD4ucuT6LUWAs+E7vEwvLh7W
AW/rDPKPtzPfkvB6ymcKKrCtErVP9QpSx0WC44MZvxWK5svIyR9Rn6WhfWRq2QEs
FZGIrsTm/CLsfJrJCnXoc2MuQIW1+wr8lfSc+N44oyljY/QZbHR9eF6H5sS8vAkZ
csBHFag5EMgw/hbdILxUi9ml7E8vjXrdg/5jKl+0UWJ9ru71BfuG9LvbXB6wJ/Ef
2IRz88Mt6GiIhfvKiaUXHkBDSsclq5NYj1i6NRR1lHHjq/ehFjBuWf/cbeIPLB4y
nXY+UI8e7oOfyhRr7VMS1eM/NdOcA/CxTNaL7BS9k549GlAv/r1Ze+HKF2S/XgtU
2Hzg5Q4mH2biwNQ3aRVqZmWuJ+TMuAMBehkXQWiD7DuAhstHVPAzzQT7KHDYsw4/
ul0GyOm3ryBHY0KIMW6sJp8LWmj/FiAMEDuRMcjOieAIHtfgbLmbB47+DRK6T2dI
FHTi3ob3kgtLpBf5r5myaLAq1YwGusksLguFFFA93igR1Lv8gXlg3X/fs0VZ/LA0
dp4FbX4WdUW+jHYQzYggjBEUQgrdfaPsY1tevH4oiCHYbAGkUZizdOkF7AJytpZr
Ss9v3P7P311UFjBos3SqgB9JG7+fideC1KIheonGEtqwWuj/rYvTQ+Gh1WsNHP2W
Z+1AZ7dit1V7hKJHM2pAdgYSsnPi7fuwFlj9suwlwdhamN6jGhJQ+PFlzKgx36Zb
TfNlaRIeExNQosQGENqThqiXG/gmhFdxTVi0IIaWeV+0AR9jMTw4J8YFIk/n1JM4
RKoN/hhjcb4Zmw9n2p/SLa/rrCyG3iJ9T7D9Woq7bSLVgecppVvAMDSMq6yPJKip
aBjHGPeB3ieDT/wlHP2VcyNS2S2J8iOcxGgVHO9FOZNMyvTVD9xfqWT5bYk8cT9t
C89sVE3cvkflArxSkfnuPc96mVgNM6Ykq4LBIb6kaQmjg9srjzO0ZK8d+zgPbVFo
HfNkKDbkxmickpgzD1kGAj+hXQKQ7HfOzF6id+T+woashDlPk8dq0xoDPfFGJtMH
fcUiXa+dZL14N7msX0qz1vZr2wDJNDUZTOFLNP7v11qBqPLmn41BVQ1BJk01QqLp
o7jKKd2AmR127PUKG1SycI2UHVrNKKw7RoZOGLqOP6WscqrwS9Z9SyTx7AxDjKEd
d31L5Fm6R+VXVH1rU8UXAAWY0X5aa7QE2PImfX1yEy1Ks5JVVfVS53HRvOt8pHAl
zWATZMmEwsqwIJUbbA8j65khs7HpFw5JCaJl+87YIE9PPc3YFl92Lx47B8gjQJJd
S63vxwTBZLNtkcXcmRVd+3lWY1KOt1StnM1o3O0/PnYpRTs2ySLLnEA74rh+hLwk
Fccau0E/WaPt8nAU4TIdPVq2OqxdlRl9uX242X8H4GMnK0FsMihJWlCNte3s5zIA
AmcuZzseQdNWbAO8I0oKvoBggxAOR6FRvIkCkNchCupVnE8gil7mA7x4QEE5ofN+
wZvYS1LA++aC7avTyH4HZj8VRgbVFWPEYYI8DQpM3WFbfVpTizGPHjqx7kCmZ070
oAsTqJ92BR8RjE8QZomHPScYX+wOrXuyGFYEHWwSeYSSUMiI/t2HuHZwLo1ao2Ik
VJEpS0s/AmXPKw9ErQwlxtdP35VfA10nOdUDi4HPPGHnlKPNqcM+vebHF7V/Vahu
phIpI6fCeCvoupAedDyGtwshOa2oj4JyW+k/LOcXm7JJdcoXHNfgxTTJZ4dyp71C
CzVhZEi9FQLKVOV2zv5op97eh/lqSTDOzmTnA3nZwlPY51SaX2gVXOUTWys6FvT+
jzfhcJq/CfbhvN0SeHFaZpI9MDukHvOfq3e3EvdS7dHrmBGK/pxxPXJ9cKtIZC2u
Dfa91vtqabktJq0YY1cfEmMhoDYvYfeEy7OZNh5/LLt0O4n80ypJvhf+J70vyrIQ
LAnBU9yOuYZ4VkR/H/egWt9LwMApjGszPN/4HWFY4ynWctxAIVc/+8yAJZLcv8hS
z3EtdDBJaOsR1MnK3ccfVrqZuocAjsbIFwt6O6znqwFM6+Bh3Pdbmkhwu5fOFA5v
cNfFGTL/4mnU09zvVx5X46NCEmEF2fCEnCPV48I74Udj1FJmxV/DS9rNIzRBWcqx
RBtDBJcvI+A5702Og/oJZBYQsUTm3zYsOkxLCpShTb+T3bcLNRCkmPYnVXvKRtl+
3o8DsJxe9dHg5fWUD8kdIGOUNbRxsL87AaibNvHv8WXjh2vugEhEk/RssZsHJTkx
nWDzHLcNpUmNjDbkWXJMdmXriKaeoBnYkoHFdmlcg8Xp52TtyQlfsdJY8eQAL0/n
gTeS4Aw7dEo9wFXEMAmxuutBN/IRAbArGA3H1mDfONltCCQc3wU87rAkdHhGyopp
GPE0gGCEH935XwzIiF0gvZy0vYFgLPrdMI5CLElv9OHAKLiDo+rMs/Wbmgt0oaIG
xVQFjr/BNy5SmOenmDvWc3t7F8PvuUhlhof00+W565AO3JX0huTsLsL7WPeoXrFK
dgFriYoy1BRJUvOo85jtWf4KZvtJazl+8ioNDX+I6T37C0GdeN1LNXmnfHa9ZEvD
lYzotOuObC5ayBF2vL0HO/bF7LRcMMNR8WHUPjiXiiT2fBgMi6ogs7EJBQoHO83+
7Lceu2BLSQYfR4dnue8HDMrIqpT9Lt5k1yK5G4FzvymsQX2QQyG6XM4CymFpSm3E
kZ/f8M1m+QGQQQRjUHR8YmIzX1kLaT7ZEcegiYQ8OEfOtoaciYmhcEJM0RrMqHF9
ee/M21fQrXoVb5ZoShQROmwBAOZDG6QG2yUX0BXUcV8ATiTQeWsMxyANR/2WLAP9
d5NRd/Rho3c8uYmEiXZ/5b4yHOeG+zEgRAUSoABfmheXretLHEPzEtgueyMVig6+
pM/+JDdKy2qGotL1/+a+qCfjXrKG1L/Wo6SaPJl/nTLNBKK1WwF80pkw1RAq4/L2
oMRWsJX6w62GmPL1Edm4oo1VERdRg0D18FeHRuKzvTDPnzO6fMKN6yhrbaB/5jpp
XXTboWco7XWRxz8Q1zWOAk/bPVJ7WKL49x0R5updxqP4AqZL/FhuutwzVTZ/XBlg
xSH1cWZC4ykkhq2bLQMo4xRuhuoFRkpJqwbIyJdympMKHhS3xO5ZgpqArdBcUJGX
7ikUogu0Krx3Pzbk6PsoAbBuL/0KWwcq/cDRBqOiVVXg36CnUveLcVOEbbrmL812
MrDgLyks8RZisp2y2D/vnrygvyBpdakm5F+nxVLVktqhZu+EXXBG2CdWNZtVxGrK
E6cmSzaB1z7qKF+29G1gx3x4r+695oH9uPgW+1bPvkZ1a7t0//g4qX4M9eRtsyD8
4lxAAW3IbLjM+3tOhX2irYDanAS39ZXI1mwwqwwBsfXMCAlvHIYIB6nW8iR70n3S
fRibfhGUNqWoF/YD4hCLV61o5WXRwYHPJhdoicnxV8Q2ELJNKs5wfDPnPQxxjSNk
1iOEByjRiHWdh0mHoYldYMVObatXGMWHDHiz+SpoHiHnFlomIlKWY9HyX/LfFNDv
s6d3DOheseS/yDeSiS1AWPa6yqL9RvSUajUrmMJ/rth+4qhj3cwqNiDr2w0xLNty
ggc9far3I0GHv+DrlGSddcCSVgCPHv3t2c6cpdY9Ux9vJ2/CKlEWxpW2aeKNpgmF
79F8lKiNqszJK0aypaEJtnAO7tcKvBg1mb306kBiJ45FReYPEknWfeynXy01LLWU
aiuIYLR/yFuUBLf1/Db5Mj7bkDXiMPG+0Bu5lpwOmbsooYgKDrIzSCV5uiMbBJDa
CaKG1p8qodDaup3Fe65NXNve3i+DHdWFsxKA2CDU6X1svDVOK57D3c047Gz3G9fn
XkKszqD8SQd3K6Mzjb3lCT/fx5P6gqdvb45zBw+5TaWXkQveqb0Ie2S4nua7z4s4
gmbwbhtaUarZ+SqEETfJqqpaVTAnlUrnSbgCFmAnWYl4X7OBevj+RJXmJzI8jkZT
reoyAmio5+kyZBm1th1/hVCp7WVKUzZoMGXXMCay3cuceBSK1jtZzu811sIz60BY
OMP9uW4oZNofZWxF0NC/ciWpnggMviiCC1akBPDJ8k8XOhwehbzj79vjjHVZqdqT
jDJugCAy0EMB0Rv1ms12cqnCNbeL7H6ZfsCgfHcjIadmnCxtYnDt6BHPpUAnw+So
yWKKjzlHUAfylF7465Myx69GL97mUHIut5m6qAXuKrf1GShGskwNffxIkkMS/GAw
0hOuuXhh9g6BfcJha1BAD1eox9bFz/3BWubP6pmqCOtW0mS5V09iXJ17wl1m4A1B
pyytlqJVENkqLOWhbIIJRpLQhutmYq73WQz/Rx+Ea4KY1AiNK/HEyOQinQdLdwDW
A5xJYxj1w7FG3s/Bv+ijDYkmPd8ASlxzULh71/V1JTTNqfwPZDSa5eTILHMOeM1L
3YuCLwk0o51WnZq/q/oH5XCAd3NU3leUw1aOZjMC/lk5prSa4JwYbHwSye/Bamlz
fuT1gSHLRKrKNyfIk7eW1OGlrZZWc9a82ZpTKHp/ZMqAnGHGV+YTWDEK8/uSrSoP
QLRP73PGpQojLgayuh+wsXNHtai3+TLBktnkJtjh6lZ+5Anx9M/iVrC8AU+uvERA
oVTiO0/Xsi+naPNUggau35bzRwVig1X2hy19lPrpJnTWsHh3UkDb4xSbaHJQted+
pRkWhIYF2fyvc0qzpnGamTi379sQvygk/bUWC532i8du3QqJaqt3E8trM98Gzgf+
tHWJAN9+lB2BGOhAWUKnJBiONh51iWvBmGho6N1Z/Wc2ZisoFzZpd6G5vCZJjfoP
bBxkdoiAjHuquizHaHduD+LHHPq5EIuUDf2nYNetKsCWtplTgRhyXAxd+bDVEdIY
pOdftyH8CEcgdIqO+lf0WUWRFLUae5b+1igOWk4HzFirN9JfjGslEi3HUNBCQMvf
Oqe8DIbvGXJ+8+OlcVEmxS6BjOdRuUsFFBSw3av1MN7ztmti8k2u1Lctbz0ntly0
5g//DL3KhZGYLtOl8zSNMu9qrDBNiCi5tR2JKUCmsbQNXq8lbB59pPdTkzNP19nf
sWIaNeSqO7av2LdIstPBYe5FT2oN/qgRSydHhZlyt1/V/ESSHf5SxLnMZqIZYKgV
KaflCYPEfYlRRgBwT80dcB28TVOqtJt/LfgMqCDbexXYq+mcbGu7Wr8QdntVTaSZ
YIBh8ZUJMAdIkjPLfeDB6ae+u0cQpX+TtDiP/ZoP9XFAGEKWAW+b71BFmaKvGB2Z
unTjlhVrf2cd9UQFtfR0ZclVk/TtLoK0CWl5vHeHS87t9UqVJ16l1JMmGf/eKxWc
nDzenofbR/aOVJptuo/Je1V3+Oq6CDlxYO3C1Sj7o4qnq3al7GvS/UFt2+2vLC4p
jvLnH7Kv5XaSRL9VvJwYE0D8T84PljEWqVUbxglf3vNmjQCHqgsmLWV2vS+ykKbW
iuX0Cg2GN9PGGQ6zrCYQzxGYOQEETPgF1uGCuHBdhVybKJsvu8pUfz1yz82wK8h/
2kPz+RA/14q21QZBUE0PRR1GTRkFHW8YrG/lrnLbeKz1iei2Sxi45ewmSTjqkamx
AWEdRnLWn6HjJ2eMMWcnoGOqSPGcyVrQCzilSrMkiyl9ByR8JIyuKP9ndlnRufVt
PHsvnTQUNoeqrkklS+FSCiln2qf/bOhS1zK6GKec+ju5rWtoboQM1HJrfEk2rq1+
02xEdJ4K/j0ygLDB46suosLSg/n8ckby4bsjTx/2uJh9/zfKnP8E7HRRHm7uoMmu
i1s8JzmjHVwX/5cnKHPsCyLPD4EKTxQtWGpf4Uyzl9+vduqUx4Zb4K3wcmCMl1iY
gQe4TpbZC229V7XPaqizGkdLryzwHiNmsmBokN/kqObYa9i7VSbzRTISkFSEI+Vm
23yFu6O264Xb6eHNzzcc9GIGkNcCjuVaxypsWCMs7oCBIGd3OICNscTkWr/hVUX8
Ha+RL8ZKEL8gN/NXWPlfemczfwiuBO2VKVJqk9U90DA1GWF2hYC4fkfVdXlonq4p
KzsZJcjed0C7lczSlYbbe+uA5uxtPk+/vOu4A6pxRGV6Wqk7O3XNZd2Q+PRnKZxr
6Ib1Wol1a84/j3OXCgWRPI50G/KNB3crnAfoMJeek0QO0EsyDX4huj4zRojOvnOj
0ylXaozWh9nHDm3ftw7QPai+mWEruZzS2LOJiRl2oi+B2gHgSQkII0rTmeBkBG4c
VKJej0eRny0iIlIJZ9EZB+zb2b2hzmYstMXkxfFWawdWnKwE1HH9g6THqbrcv5ON
upijUHYKYYpFeMWIXknjXquSPWTUL1iydhR4JchGzDnXsHloBnS5llxGfrY8jknK
uit8RXlnFEyA/nxxicANhLiVNA4L/G33BXZJXmFh2stfBOVOQHqqIV1fcm3ww9HR
u2zyTwkK5WIVieomxTIriIZBF34MvnoA3kXj1cD9qKtDvjGESNoJSMfJ/MPlshic
pNm4T/FR1uSC7jANmwKoOANnGfEQ2e58HjQkOdioMfdU+tboiFYDZt6Zs9XLfhPw
Y7mOhyV3FukpAiJePrJhJEusaUHtlcxj5Gfdv/ozhtj4xA04NL447DZ+3172EmRD
7XcH3H67U3/5CvhDaQT9UaLsiYLU8bCMGvBX3ZL0+keNirlJKKkW8uZhXh9/HHHx
32ObkrJvf/OZE72BYIbIJZEJIxN4E+GaDEGZZ/Ykg3iT/GnpNvqdaZPw4C71amdn
8Rn0+ABJD6V3Sxw6o6dP/iY8IONNa8Fj0j/vofQVgsCLczEdXKbakt88j3SIQDrr
Xga/kqXkEaR8/xg5at3rsLTvLhbxnmAGNwGYYsH5qROirgTtmSRrF7rt7n7YJG6t
RbBRltR9N0OU5tEnYVZGCVe1CdX+P0q0twDyP5KAA3N2MyCdxzfhJQb2w76ifvhz
VOxzcvE+0OMPGfynzDcQWi1+q34rymzJlXPyLeOFLb9bRJdWRCYsLVctgI4tN7DX
RVffKuykYI3kxN12GdcD2YSLG+yH0UCciaDSnvNKroNAgB2n851wz7ovPIoJSWzX
xHJNhlTM7ebCa+yY2zbCVDf0Jw1Y70FM4ZaRF0lB6u5yYf8PpsbOT9/RIMSoxRE7
5g8trTdb3HJiGZTijb7EZJPbJpAYcltqibIBCufPrpzjJ6buGsWazh7MKjSmYoR1
l5+TfTeBGRGXzSptGZFYJTe3bZi6lIpaMrhHf8+TfQWU0RyYxUESqSVyhm7+qDmh
g6T3cAoTGwqzl7XOYqiUrjNUTHf14IXo2fmJqaWOXne3rw7XVH8Th3gbdeszhQpx
cJ5m1duppRzPokAcazpw+HltNhxOI1lJ+811C7a8quxRWKmI8YVUcvn+Jp/IOmTs
IzbKo36uV4CeMxSNhqZgrfCkjeCfV50KBNQHsvDJwcnanAFR9dFrSFriIhOoYy7o
33pANYs3gofODt+URWzTm1n5divojVPa3I63thnua/v/thyUB3CfthQ1cpTXRCER
50OkX84FpVqYv9aJSAwkbOJ+QYWxfS8jFfTsDKlGyFXOktoVeD0h4GtmyFfCnLYe
cGZNdTF6Ty5HkN7/1+kxlFZmkOsNGsS4gYNvTk0sWsh4oPqZ8eTMMQeAXb+gnCh1
Kye5xJStvoup97mINtkO7mHKqtZ4ALtCmn4/Ci60waglhGYNlJ8BmfPuKA98LcSK
gP+OZrnrlSj8Z4tL6GCoskdf+l36FM1AiiFJ80AmmI4KSjyhZgrwSCtux3/20MA1
bkDwigYF77ZwUGdxyNI2U/qbSAtDr4vok3bfhKsRy7Z62IKUNVjdydvkyAJr1jvr
WQx5XpADJPbYRDsAbAbFCQ1PMSC8y861sQBoJ//QPN9l7Aa1EtwI8K9WS/mwEW0W
H2ajplAznrTkkxAG3oPj9E7/TFYr77IcEqHjorb1BVCfQSMDwS2b7oHTppB8Ksnq
nvN4nopz6mK/452UHtTSrtWMG4ep0njwPP5lcmBFLYk5fUSh1K72BwpUUA+OXrYA
6cJbdgSKr4eDZL0d5oojqmi2g7J6Odj5kOH1p1jlt7B3mAc3UeD2ftFGTOTzSvms
JdcrzsNuLQtMa9nz8lmR5dzdjmvFrODmOeH80KtHcaiPGwCrPXEH4iP9DDT82y+F
fMivQILl1M6wt2aqHHHwwuQMVwmJ98RYE0lt+uERY8VKa5RnN/0JzR/YoQHVVVFz
ZDz60Sp+3jarhc6BfzVUfIzSA9DfMFu5e892hszFfT7OXHzpyRXbeBQeWNoxw1Zp
9OQYGj/Y2MxaPgdXWBQD1vpVj9TfZkcR3WPaNoy8yEnY4bUrPcs1TPw0gkwJWH5d
YwKjFL5a0qxB0l2IAL6UThtKWaZFFVt8m9AtkbNMQ8DI/cgSjT39L4LgQ4WPtOxA
g+DgcnYG5VP39fCxLpPYnSkOmFkp6jH6RXS6exKmqqx0q5sqWFSYt02I+oucyp1U
I94M2K0Iucjs6l1pFD4i717qUDT955v9FxrKx7FLLn5e9tbAFrtCTL+TM71jNunI
WVgPbZSsMBBS3aDvi/glfHGlgn3VZluxnS/cA47qNMahJ4UC9IYZlhfuLpsoUCH3
dRIbpwtqv9F707ykw5uwV57eDy2zKe/oajdrSPwQGtizbRio6Hx9S/DeSLNohawg
nzV0RN1HWAbFyGPfzyEK21jD/wyRbywyr30B+7afL5qgEzL0xv9QRe+qMvSZjVRZ
moxTGFQC15CHc7v/UPgEH4rS1ZbgvC2YebQhRWrJ6SzsCgImlZCMfdIY9Ioy84YY
hgquBrtnBRuA29YnmWNVTCR4epDSFW1OXstAP2+OKz/GwC40/Hl/KpC3+eWMFqAd
l+aMmwE3o7rX1xS7HOUEvg4gAQLvezSDdFsf6mAxlzPnDzZCsUPVb1r865ehrmtr
oJA/wFvCoEAYvUw5rITWDRd8KyqEnMtpuPrVAatw2xde02XLgiAeiziUDbNkLKe2
G451t9NNJVFpFbKhoCalR5F3uiKC1S36WRo4UVHMfNjEtxg6i8dIcz6RVqBtC4xQ
jNoyO1IIxCjBiB62qap1imw7WLXfgKY//tw6wLhHoCCESb17iIfKUAmT0yvMcdO5
fnX9UlYWBd808v+WGlq05jZBYivEBnXaHyEqqX41bKm6nE1nzZVwM8l5eE3n5P4L
jzmtBU0krT8dwOl6cCq2LS7I3vOMrhqEEwGXcLzr1rqL7QxQJ27jGHnRQbtX2VUX
T6Y/N+YDYiqkgEFtjYvhruSnG32uy3cFWqSDnivVD1IkAoxi+Q9HWLDPIxhbBk6+
Lye0eDnV/ITJExe7Kq9m4jE4AwGOWmPF/8Q4GOg6WsPZwPfkZVY7cCl5Z9oe8wmp
Hj8xn6iGj1MrrF7AKFkujkI3+BeUJCO+iQbEMhFP2ikOTMBFT97P4wts9pozOUcJ
hQa6Da1u0Jke8wVDBFg+Lb/9Q8dgeHCOsbUkSsboz1ha1saf9uFEMZKmn4Y+gMyq
7MMgK+8jnUuQVyj7Rc+yxvnt03vC84bJ4Pv2DlpqB7C5a1m0pHqpxUBcCp/CxEil
hT4x2XsfIQDvi/81vaQ41OCnj32ZS6iR5Q4bCe9riphcxUzqyBDFQl7u/kft2zHx
+L3RT0BeUcz9AMt1pG2WeZrEmgu2iKSjS4SioiQUhQr04dasQYaDwrGAE1FeLIhF
P6jo744HBzw5EDLXW1InPWRGwTXMD704miGVndkQtjzcB3q16UyYqnqQx7PUU8pD
zi2IQSCUtYVeaJo0dlYBfkLSvCuR+kQd7MnjlCA/sqr2mttJiYalqh3sB3utTUrD
PHacubouOb7GgoIFpVqUKEp1Bkf/OlHyRt+ejGI5cuu+FWizcfDLukqyXuwuKZO/
jIfDCOAbUkeYEIOjVrcgj5qUWHlNEb1guEerX9IxW7WI3oXJHxtoMABxK7ovOm1E
13MGTJwpyShWxkzdk+tK5U0TLOQBZe0MduqUN76XtFNcLgpKhf2YmbOiglxSbvL2
F6XGlBuyP7JFPxE0OHjOooXbsGekBHUzKoPux+VGJNU8HmdyVsnCdvBtGY0haUao
V0+stKc6heuJWphDnGXlMFBLE3MstfU/1Wz55WT910pp9nUsH6jVG9nv5rDMzkuM
moKIW++lPKhs4tIZ2MZY83FYdIcoBeaiOccKk4XD4Vb/uQZeLDSTJUmHmjIlpVwr
vukWhlSbBNEM2fBxEfjTYv0I9rp/kTjxF6s+Oo84r/4TBhnQZL0FQIrWQIw30j8M
mwdFk1DjARY90xzdoRPcuNd4xoEb6O90l278z3UUlD/Eyq/cGGUJzRSSk+5mp9UT
pdsyw8y2ctcTqTITMl4mhUWqUNPMFUZ/gW4wWVXloD5lVMeEpPzoNsKbeUvoTxnm
xmadWVqoPRvn3O03mie4AEtRR4QUXyFILBWRlgvimq1y4iIRRjtDV48aZBEzidoK
58RdpGGnWkoGhxa6UCWBdqNAivrMVOr9oKMNtABJ/BQ6uzw1ZPj209uRYhHGgkqK
ivK2XNJAQ5ePk+a1jaNusJIt9q2K3/J79UqO5wFqwowIdakIWXdoGqjhfYMJFfq3
C7R56W6qixfatG/eWiX3k1PwimHqHaqyD95sNNopKwTaAIAcxR9qEC+Cq8Y/516P
mMVlEf0fr+G+7Ryn8Wbcu4bsZaCbXh2jle3szP3fjN4dKoYQuJfVflrJptt/Xm2v
GkTcrTjaex12y02wpGqBcce7xShhWJzY3Bzk/yxgusDP4vhAvP2hw6b2dIhdflpg
354lE1mic78du+ZeCLEzUCdsWnYWMsRd/HYAOVDg6RECFJGXGpZwBBSEuIl4sDCh
3syMI3ZvKSCX+zqWd8WMVVt/SRYqfLMGKWdcpwW/ikB4gmVDTS60+z5EjsIy5p97
fRRGvidAwhTON0xVnbwS+Zfynkvn3qoiTrQh2eRJ6Z3NEEqkagTi7q5q4wCWngmF
0Y5/dpchck/QahtLhVobyXW99xQ/PG1ymlYtqE4YV2o7/9p5y6sfQM0h3lLcKTZr
63iaZ0bZVkcd/7U531NMUYo45M0xwm820qbAXZV0F0X0DmRhDVwiVKo6XUvQKXdW
tT9IZ4FTahoM9E2RDNzt5TVWqPs/gZMUdHgO61ipGpPJhmbC48y4b/zeERUitWnG
9OV3UVjRYmBrdU3nBhwdFvjwDy/yGR8kQis+bl2qFip1QNLiWcJJbULlZ5OUCjGU
KtIzxvLEeCYA5PhreLQ96F2YsumY/UjJCRFelpZZQcjcEvaAAZ3W49N0KFUQxKpy
mcCVeTUo7B63vXvwma+dr/yZIzaSTKRwRpKzAqoZZCKQsK6ezUj0iqqAhmKL+Y7y
ppQ4kEv30/L+1mkaPTQ3FhMpN58OFRoi8uOJ5Fmqj07WpOtHzN6wDC38bjjBmTmX
4K9Ndpt3L7op+pPV3A7b2MVxeBQXmr3zg8ww0Mtv0pB0iNKGfvl6cpRff9v1Lh4U
eNmc2CN0q3TNd/TfnjJUK3LhPU4iDo0yO9FWeYlIEPqyTahcV8di+yckiYR1TNnG
NObaVvpCbmADxKY64xA+aTltdVxFGV0OCjHZhapjQD4bkaY0IWd0nfzTC6PjIzMt
4Z0aJU76A8yuyxU0dIJxjt9rYqqgrqU3Fc8LgZPmR7gq7YUfwfAieOvzKdip8pO4
LtJdn6N5bCTIcpTPj5vArlXL8mOVZMA25nCZc1f8rFbb+ZMrLiZ31pQvDtsLTlwW
2NY6Qy4jHJdyxq4wyAgsEoc+qlZJN/v0oyL+9G+H2d+bQTeJclVM8olyHC7HE9ke
yvimbTOBLN1OPIpb+NnNythcQKPu5UMyZq+A9qdEZMbf0ux1Hnh0c7UGOJOrLU4V
Zh+VnF0yG+PZBDRAY8gf7d6G+eyGsDNxJjDzBQOGcu2Pj225xRQGl7kxQXbpdIJp
aLzgt+U/YbrkS/JfRfH4oPZZf5wGSpr5lR3ozLv2+FrZes60UEUfOGbAyKkEucQ0
tn7hVMWi+HPbbpqej6YRZ2E7B8kv53zaOVCz7qN6t/6BLZ2cwebHpIegi9q76nEE
x/PjKlrbm/ic5g4766Kw53FmTgSh1tYb3l2ZxgumjrcCceNySeCxLIKqfUnQCmm/
cIspzWIlAqPf0M4XVJKzutxqBec/xDv6kHLB0FaTVsAd/O1OxPC3zvgXsqaJjMQc
mndsCiMdsDu0PaON4wPGYgW6yUrNTkw13ymd639TMMyXXyNUMiR53XdpPx1r1+hG
OeA5fOO5gzl9sEbIS2JvOFTfmtTyGnILTwDuk+WR0qMeCUMBRyhISVygByo/rdS6
fSOkHJeHQJHFnlRkOz8hwuI4lILEaPUGZtnqQ8pGO+jYqrVbiJhPS0MDEIalyeKD
qjsrFq/sQV/hcweoeVxd/hU2iYi4IUoNWjFv+2ryc3yp8dUg5NQw30v30/bkqszb
Pid0di6r9Rn8dsW7sll/CS7BJFhWqHptDbPFntGA7UrQu6uBZeYAU4lADr8qeL0W
gEtleEZMqo9Jv6a1ZCWfzdvdZOSOlM0xkfUo6dAVAIenCqfBBAnq3nWi7FjRbGnR
swWIzoXK1xgrXwMwO1YKnPx7rY4nOMgb1wNzEt/z2q7WDoGzxQXHz8c/aFJ68we3
2bNgv2JpKhOgwlpyEWu1clhOu+cxtFeooIN6gB+ZYd9GvGO2yFMTVue0tTZ7n7Cv
Yp2fohaXXKd1TVVz5GHQxeZtDVrPXzOKQ4keyIUKYniVE6RN7H8rD9FKOGcKO4Rw
1/nTUtI4wAYxKdE21wZFP/ZaMZCv4sRRG4zQeeEbayWlEiYj/8NHufx4QRq7FURn
jDZ6Qxc04Zwspnni3TI/MnjyKzFCXx1VfkZECBizGPewXZwtkYA5t/n4ze5wwVou
5II/otq9QSgRhiTewkPwiSKk83Y7Jwzb3Ox4pQB1/ZlHfY2weLmxyM8ZLcCNPtuw
hCTWMKDvxhzlFsz/sqjVmG4picabWtk/jOobRCwjXQAQi2z/DfNAaFknCC+HT0Ao
R8YjEiMDeAzhZY4+2s3AM/m5qQ1yE4KKZ9JJmOpBxVT62JO9lQZg5ru2/PcQWC0h
8T2NKquECoxXeonxMB3TNyZtNgX14kASSaRbR+LN6ck/Cz9AH15aUWHqeNPRDgpU
BOCV4+OJKb4acaGGq1jWh6vN3jCwuDKElibB+ceZhDe/ky6EyJPxq+p8dv1ImWja
B8LRTUofUaMo3sgVS5PEujAweuFV5DW07DP+uEXL0Fb3JzKrEvqzabrbt59HFYKv
JODF1MO7YqQSAca4WQIWtKiQFwAt/IoyQBJRmK2DviYjRQYCMPGfQNqGPdgMZiXB
w3CEhstnMpKp19HQr5B2NqCzuUEG5tqQqo2AOE5zwgf5D9TLnEExSF1bbM13fBVb
7L6wxQsA4OSGpx3JRvOAPvKRvDvGTijTVZpF1HJ5cA/89d6L+GhI+TIJY/SGgzzc
pSP2rEQWxmE1s2oxSKhE8looGRl1KgVi5AZZnsc3fcVjon4aHkIY+1AztsU8k3bP
Z/Jw1MTvriif+D1b5qt0DswVsdAzQ/src6Lk+euzlSvDdFyxcjP8vbiasJHFBZbi
5vnexXvRRulB6MhTsfoYNwisbQK49Q0w6QJ/t92UeRu4dYlI9wPfKHw+sSUYJ6YB
iqU2ZqkkMEAi9W68KfoJFoceSv4CITbhUYCc8B7qBy3xlhCEee7wW2MfDDs3PTJ+
RreDt8Jfds7ciYXrs+dLTV3yiqpNyP8HcNeCjSCkWJ1G2ZjGH8ESlet2nKFnd6rL
mKmWIv3ead4g1jKjQR4MRhWBzYMYPgRVJT07bBss0otTGxTTE40iuAYw7PesMJmQ
iVsTFBuyo+1ul4fRYqzL4DKzEUK1WGK2KJ4iotF7GgWCfdXZ6XzK6oEC+p9u6XUn
tXg4b959/PA/qoVJXlq5Ko3mzy7zjVNNOeoFXTKrA5GQWY+Ckpuy1J1eyMs2D+89
7+SoBfyS+GBK9yWKIl4Ea9pj4FttVwZV09nuYheFA3vMgQz0RyDLcMZS9XPNoo3f
b/95JRFqVIhZES+B59AyogXiAHgZ7xk37brqdKR9JoSJ1HmYqpbO66itKsebua5t
IruKuSIQ+BW5P2cMRL73FPMCPczKBx3F0sbwUorReibL/g/jf7KIUopaLJlXU9jZ
ComnSMhJsnwoCrjcX3+gKUoXgj1bA5wA+yafsiJ1jXmKcPC++SxCoFPNCtLSy3TB
8r8+6mNlkwksf3qvkPbv8wwA9uBIjEIy07E4shDTuCiChaczyxmU+ys1gnSgKjGv
cvoHkIfVv7Dw/bPZfxxT5lN9zcTwUoD5rqoAIkqYH7NPiiOq3pdoVvmMiOJ0z/0q
5MjMBKbigdPsflIn8AiLgENBxE8/FJJLY8DMDc1rGHUydTKnasJhGTOPA4L1u2DD
7rDu9Vrr5pGqzjDLbftvUzd1xa4+KU9lepCphbtw6d/bezpZM0N6jYO1552EOPLN
oln1bE3YXJcaewpEFnQQNKHJ6D9IiQTncHrAvR1vMtex4pmupOzxvGMxMPOSVzuu
vFKAJIh9//zQc2QTevaG0JmP4a1sz9MJnhJS+urjRFR4paZgtoRMINXKtqCli2i6
ohEByYrJpIUNer89j3AFQ7JP1IqbJCNq3kZqrknPjRbuU1RK5g4tN7DPFlI3KlHR
X+QrzApX26Izhb4NjliRdVM8BJMY4lz/0o6A2QwpxtmbmjAcGMJ4EaNhzhQI5uKe
YvL7IP0mI6WREd1U7E/WioKq7lp8zAnGvxB52MuJQ6+2Q1QVSr50ExYxJbHcPfVW
Wi+biHNiIjKmWyLBOI/yvghP0ZloJl2B6tZeiWchHh4sYkN74azyJyS/ojDRNXI2
v69Azkko6ra50K0TakFEbTe3mrG0DZrBZN+ip4Zdjs3mEktuIJAl/uyepaIZsu5a
5KQM2onM3yVtLmdu08Zxq0C4xmoosVIIKYY0zKdO9WnQgKg+VvjLEmw6iQbjstdg
Z7hnY+m9kygFsTbVN+qyd9z33k4dj40b8FkVghg5CgZqqNxEesiyf/cmOSMlUlH4
2GlWr3QC2SwShUt0mSKlZazNZBzwkaEf35jt5LtbjKscLOUU9y4Vl8d6DIsUiPq3
uVNoZUDGBrR+ImV4mTCep8dGuXV/Nqi4fw+we5YtmYqEaTKMFpXTm+gJpXzQgujY
irKoU0SkdNEsSshytlx7F19dXCsqN+AWXJpV9jqZAmV4YFUshUyhD7aTVJ4TxWho
bcOp7LV+hZF5UN7GZ8lTYZ7vPfwgn6+mzG7Qetz2+8bCQBaGUH1DxPY8eubQbFhl
9VapxkMJ7Kwh5LzIxVQFLnnhv9HANsW/hHWANzny8vGzKJJLcL4yT/eYuVJlKlhv
7WTOIK0bQEDKcFrU4UVKOdX85V9494QqF4DvFepAMSUAm006P7/0xqdNYqHRMr1m
fOu7rc4pLYhRgaLulOLrAWmJ8l9G8Q8dNYyO80tgR6BHzsI7i5MP6sqLEzmcfzF3
7vbWFV4ejmzAz4/6X0kCzRQfytTXAoAPyF6LsB1b5hC0ta+rULG56bfOJVkWKK1Y
1H04Ac+DfqUFV1ZzMzRbDl5he8NTWh7WcLX6hpUbuK+oJC+TM5VqnRtcEg7/6Fbs
4dWfBKiwLhGLen+Y2u+fcIlmMrKRhuqSW7ZgBHT3QEb6fNuGVYqIufyT/cvMBbLS
TjqRXNTNxAksiQgKQWhpob7eP7m4e0Hwulp6fKppdZgwnJnpA1sIp1+BlEBNIa9m
P71Jfq9JsKC2iyv8rJpRWCIa0oIFq0VIHz1pm0nX4SXwKKh0ifCvCwgb11/dpFKt
jIUEb4AtFLr13Kcg0sze3KOh0FyCcp7xPXcAifaLYDsP3m9PUxnKGS6GVcH272yv
r2qYdRKHmzOZyFpCkkXOH01YOCnKMSr/NVzRnS/5e7uyeeaUkqgj6ehgVzzk14oE
tKKUaBHkDIFSgrW6HdfDGGa3WgbRIx6n8uDvPoqQpFQvRKclqjrFLrpRPPX13Y9e
B04j/KfJFtDuHSenOhdwh0y/0kXKzRKd0/KvzxHS7hUBtkgNI8oNp9krsgcxwY2L
VHpitghzBDytwyMq9zsAMZta0qRAENDiWRaSHBIxe6AGIkU+/l+cCPys6nOB/krf
rB/lHw3kQgjwN09BqyhqGDiSvg8yhoE4X6oOoBQzRTW8jLsTZiBKRPPb2S0bdaD7
UU8iEX05nKn8seL9P8lA+eIpcjIxf8LLkUWy08ZqhbXJQbXG/r7hrh7s8e75B8WP
YM70GSpz6iajV2o7+1gJ8shHBqNuXj6yRrU2nSHm6OuuD6w3ozsncr/n4SOJUa0i
orubRlkXry38/uQudNISvxzc8+5FlXYhvyKWZAFvxUuBWC1s6SIWd0Y/08vvixPH
2Wht4gkrZgsQPNa+4R70+C+rLg7I1rqx3D6yKLEgDCzz/GIo/6s0Dl360eg30cv2
sx9a211jI/8yqnk3XWK1xqZa9mIJtUsiVK/+rwfGaW0RCRnk4NFsT21kSHaa2kH5
FcGquhc5PAMhaJ6cGQTqLebXflZFOGyFrMhUIBrLACWCkOXlau0E7GKWmvYC548o
bnCxQd7d58BT7YA85MyNxM2h9WiY7einCE2HWp0KMo5hFHP0UvffMoIhyULd8LYx
R+WTRW/bD9TyoJKGb7ssIsJstfBWaONqMhqbmJc5fVhnxLw69iFc21rKQsGVrEgE
fkbxtdWPhM+3HEYIaOp64kkKTSv7G3YB/bIlsCLR1PuYsEIfiMo8yoxkcBNCcG90
PC3VxCUZ7gfnyhVZdXpnesgk6vH0GaEerjHJnhsCvPAXcy7tmjyGH3PyST2IFrQE
roCNpd8uB1WhagNawKIizTGqxhQhaApUYdHo2pnJ5pCd9eXO61rKzypmt9RgugZy
PEL28Wjvgm89yHDflsxJzy9xWehuC38tkFcQWhL35IKkH0vx4iyYMq5Wxh8Bb5Mp
1k6WTNeJGO3MPFKjfGm37vftCEPnR/flkfUlshetJOVU+JFYJh6AQRaRvXZDLZg7
jiXFx0hClNPhTs5Kbb9We6fxKsictd+knDJ9al2Wg92esrV068641Tci78yUqZBi
gHad8Pyuy2n3YbnU7z0pLXxs60PP0IS4fi8QF2uFB17nerY0OY69XVswoiR/Sv0G
tLEP7EA2bYKKCt5xhCQWOR1sOdLi5zeuo2oHOm69E92i/wT3SSkmu/jsAKXVS82K
jjZmWU2DYz/iM8mhdSXoR7bs2xod8yCTCdiHqwenSFbzEy7ioDi90/3ZzZYxDXgX
RKj1joyEfmBmIa+EqhiIHRfKzJwTlmffABGgaLFZQVNikCiae7+AosJgWCr45zPx
FtFZ13LMt/viqN+UrurYoXOtNi4J3TJaA6zxt1sM9ZcgiZ/wTZYzTYCOYULTTS4+
U4Pes8nbLqhQrqFyNmlpq43FCh3bX+r64jktBuo3Tb9ODjuc/l/oiwPDtcc7RmwX
USq/3ACCZSSdBEJN7/c+UGcGabuHHQ/aUIEqKwvflNChS4Mh28hdELJ70W4Pksrh
+RcZGdUqQ7x9zNsxfMbMFfKNBbq/uX56OI098xWDiwZuzj4gPtaJn1BIVlFuuJDd
+9+Ffke+mnTclIM2HBAMyYPkbX1EuCwhHrmxWvlxTkUIb6eSMlF62kHhOpzI/4fZ
EDpHbpQwG6Bk3ZcsM18QYcaK2+pDhOSuzy7h4nsKQy1t/WEfdNoBinhhAY/p14tA
L5fhcjnoKbYpn9xzjpXvaWhy4KYrgfaA6taL0AUJC+ujlsHO338Ndik90mmL9Ecw
A7im0IFMoQkNXhyaUoom/4a6IW3kuWk9ft0Lgzu8/2YBG8CGZLUUg/h+f7QmtQvM
cKZYuTgfgiaAPFlOdxHJ88cbLv95moYRlinnAjDab+3OMBUvkPTGLpW/KwpPmBeV
IKS1ZSfR5CAjUKdS7Ekk90k0p275hGhoRn43lcN5fA1qM//hArGUA+y3jYKG3uPh
ckSHJG02NeK49qz/s/bxnM2zUvZat1BfBZXOEShAPmukATCX3Ky1yurElpIrHMqn
l8SOJ+fheG6zGre+uyN9yDd5ylChf5c3lFxmSnqoRnFe4KbxHc5pjmmCW9Atwbif
CvJr8uFEeoVJcNCOuCuDAkQfsl5mso8H5LzxdyvLefbfnYu9dXZixFq4QniYbbyT
GPTd4f6bJ1ZoojQ/2M+Xc/DiaLSNxICBcnjxxOrnYPVguR3Oe8/zRNwlKtYFNPBm
RaTfoSMjnZlAfdqF4LJJHmhoETATvr0EZKSoY9ZYZsx6zCR1qzZRaa5rgBCafpw6
ZoLDfPzJl9MQWcCL4WHA8LmhYif+NL4WTgAmt3LBTmXcRSqWQ5FCGqhc1QtbpgBg
C8HQNz5iHcwMIHOh6ftkimqR+tlAWzcdK/vBFabKF4NMEyC7q1/cl5Y5ife7ysSH
XguI5+lhqqIZaKQxrIy9rB6VTpoy8TRqVNsJSLs4LSMA3PC+Hqo0V+qwIkt54qwl
hQsuvV9B45zOAaN9Y4CzNmRkBkXl13ZsJKwm/8gTGLG2hwCbTQb6f0UxBI4cI1Zu
lya2zqOXeJxfyoNLGtkXxNT2K0tziTo4oH3H29USe47AlS/TsD7cRw4et15hXniS
9LirVyQEGfLbEp6oGZay+w42COBopaBMNesrVQFEiOldec5evvSlQ9ZnVu7YzEYy
vc3hZNArABXwshGLL2xCZVo9lag1ZJxgSyyjxj8ujtOAbCxtYRyZFUsNXMdxh/4L
O90VLe+UmhFXRDFlouye3eJAQdIzzJX4siBlLvqHRlk9sFDeENMfVXhwjpMIv+CE
bV+3mcxudtoXbksgIu65oekLIwkP+PA4fQHGzXaHT/pN2q4oeFrrASQ542BCY8EU
nwhRztXasPPGJ+eIWIYQe7gTsDCMkZwECuOalnHFegtpm0H99CNu3T3SXM5L/8N3
JXw8csiWCBt8rfap0+zBQOM7Adz+RiNrR2usXu+uXY3cNECiUsadso72FitWy1R1
6HCiNeZOhy9YfM0X5ewF2Us7IpkCwN3j1sXL5icuMFbDTnUYrwQN6Ys97bvdBNqs
CDI20+RoIlUTxHGLeKltF0LNSyahIe8H2cBcDM/P1eskXUklOq1JDco9KKoD+a07
bbeUfvnbRSkywzWNRjgbvzEGyPzbPu0Q3u+ABWTBBj+nVVH7WICUkUiQKnltiRnG
kTUZ6xH6ntYoAb+8JUYniE8nDwpVAapFANQL8Vra/bfujVdsOIrtr+IiGjzvznPz
+fX3ja4BG1QubBm+o/aVG+08VNEM1hEfBFfh8rfbQ/FglBYcyXSDo7ZusnJ9sZUL
wu7DCHXtcs4wBCynYqzdNUMRsqZSgsA6I53CX9UwMkcuikTnsYiv5evPjGSg/rSy
EkeAZEiE6snbQZCTOCx9lollGksV3PdSECWDE5uwJ6GqDdMIlMkp1OC7co0XVFpn
196rUukmQJZ+7GbrDe+Y9IwVQQT/hBs/PaHP1wAmBGNreAbaAhs12aILMJFH3Owb
gAZfZoZ6FLwEUWtR3+JnGgL0Vtk1oFz5zP5IhWVsXENbmXN7XWzZSOpQoRf0Q00V
GjR/+nYADIcFa7SCCE8MSzk8oJd6iZizsSr17Vw66JmuCtEOU8z0P29f7AuJD7SK
auWaxmw62LxKBbz/2myUWmiCQ+rZLtb+Bjo1a0YXG9nvBVN9GCPMhk2fhrdawtVT
fbjGiqd8HbtO1c6/vN9DNt9bJyPX27Vn2jHJ0GUQIuueY+38HeZY75omKfPrDlqU
u4J6dMnxT2l+Wylk4AMIuRz4J3JFFpriEktR6DUC0ROYkUqc1Vu2zAwZWmfZ6lv/
Gku1e2vQ+wywHhvEA31/anmShuP1pbC24SFAVe9ox/k61wOfX4RPw8KVCog4fxpL
jv6jj//jAHYdevUD5S9pm1JRhwbT6ByAinbFkxcViv3NPhj9O99+D5Xz7r03CKFq
eLSHQQMI3vkZIDmdRwPsJDgAX0KOANDCsd6uur1gKY4rOyS70kqqGI8SvDF8O8IX
ilPegsfglYMZqid5oB2JJT1Lxv7g2mxcRoVTebfmPyTbn3Us8nzg441M+PA6gWlc
ySJCQkIyJ+jChIpQUOTyUw+XJET/kY5UW6aFqt+IqUUxwC8w1Xsz4AIlTVMUuk1t
P7VUwMQpjEKzCC5kSK/i5KnPR5TGb0d/eRJQGAE/Bq1N6xzsUnOod6wFWzQ2ti2R
v41LoXbRfqeaqo2U5FhchegY9iIt4xG7GFq8sLAc1Fl0/7yrryKLmqMuk43cwGNZ
jk8pLPFq/ssEn8C4YG8vtfjfqncCJGUpTXYwn2lyZAT9sgpwSYrAT6qkJdIEkISI
PR3FjkloAmv8eLmUqQEh1NDQlb23TCAYQWS4Dr5kDfOO3Rf9cpBYlARvOCYU9ULg
WtFl9P0gULXd2HqGv48kfgOckGM8JY9rCt1qbW+m79wakqCnDcvuhGP3Tw3XcGeD
F2i7vdXjUfLfxwboOoFcL5kKcsSOOun3UYTiqngfccUI9PnE9I1ht6l1JN7OirNf
tMp9gM9W2PhH7o5PGGg+HU6n539ZG0Z/Z+yYsSykMOj0nwJdKv6v34JtBUgWEeb9
FX4sdKjFy6e7/p0fV8uSu83HyDqsHxC4u4d0mp8hnY0lQWxxqeZHbmaMElVl2reX
lqHvjNQjeynKQbDD/HQO3bZ36fxrO8hY6j1E0Vdvu7+lNFaIFBjcJupXbD3O+Glh
UwC+D2jeoj6pTMPjUJZr3aHsFy+ajowwsSrj/Xm+CwXinWtkcmELUepV7ViYXVaV
c5K6pl6lU2nOZ5DsSdJPr6WWCFt4zXm2Y+XRPN7RhmBbFeo4Kkb35N7GVFB3Gd6n
CFRYfH/5p/OjuDd5pWM9YmP3jFycrrJM7NI5632uMYKquOag9/HB3LstS8/Trc1b
s5Zfk8Jj3zjEC5jThCCIz3mcIcfZ/SWodiSN5O6PMZQ7m9qMu98SBTHexYRwf41H
99QTnYDjZd/LgC4pIHAQg0lKEJhFKxT4OEmEt0ZecyIjMsaAX+x8J6qj2e/PY885
1MS3liEU3mczNLrDSBEkHn7qIqj/D/BkL8dUz6bcKsrhusT+XdQoUJyLhkfm9+9n
9eipC9cpJYrtoY3rfNL4m/i58Bdn6QnV4Qg1ljHognOK6cFaEEj9QoRTqudWN04V
851L6oSxncU+Ds14unXiJbuOoAVcYBPT1ndyb0A43eNTfZoBPc/kJP6NrptBS9VE
KbMTj7NbdLpCEP3m8ibpk0i/LtPg4UIlJQsD/FkNBqlA4SKh0Vn+JKR+bo9IHyyk
usdfxAISs0d+JLOMHs4xthn+yS8e1uv/bTbqqGuVdy3J/joWUpx90QqoUUGjvK7M
2ycVDfvlsELE1o0d+uC8Xxk0KLT99WxBXiFRHL6u8UTGtoqBOCsphzPmNz4HBaXN
vaClRrwrpvFPKoo8aWrrRKKGrNIj3edj2lChWwLWesA5K1pEpUVeQsIXXwGJnpta
m6xg7cDpBnHhELDohKFoNZJHPIO0wjLJNo9HWO3vq9I0SvsDB94Cz/GVX/Mnxnpp
fbqHEJ7xhmgjCVm50ezUEvZw0JiypP2y1M5I61xm09QWv8di46FKBStjfQWurjmZ
ZNDTjtwhJz2UcqpM5gYc7vyrDQCs7y0wpxCBzZOKusfUebvmUWM1WirWcVTGjKdL
1+r+Pt2gorz9HrGzK51QCZzKjRwM9nNejL1OxHongxQg3u+d/G1W3a3HW56ujasV
74qR72g0K4V2XbcMjq0eYs1qEnMkw5WccLNfZKu+FGOIyHcP4WhltexGKbBxTUk7
/BfsvetedY1Z5M3kejjW4+Z34zy4SYs7Fmcj68+2pR+9XfY2D73fXKB57LN/ZNsy
+VlavP4R1ijtziSTcIWH9B8K9zEskNejB/6FYaAzmJ7OGh+OV02HQgGIqy8WVXtT
1qhi5y1xopwtliLmdZX1wdN400QsAgCq7xs01e4N7GeaM2qLXn8tH/ShZLP9NxPU
US1N1Wqmo94+gh56DjvzrWLUCPERsGb60Q968Ip/Xn+QNBDkQ27RsJrfc9wto7VJ
IaxId3xjox6Yh3JaJNgeykky8sTVrXQ2H67Ik+T9LeuZoEjiJZZAKIorEvXg8c5B
n7S6yfH/W/p5pLrs0wy3YOn8V5cbR70KcfsZvfcHehD2Ni9RBN/NdvRB7wkvyI61
9i3kTrwxRBkHbNqtUsv8z1CO62yFxagkmkv6V0tHcPCFrrH8BAG7CJcZGLq3av5i
wbajhtzduEgjQjQmwYVzYU6JLzC/WyHmqOgh3NY6PEq52UtpBcmLE/aQrn0Cne2K
3zhv0O3REtvWkoPlUvIO1gYcPE6PL94QqyD+WAyCHSwDlW/dYIFDRfUAaf1gd9Ak
bt3d9gpch/9MbpvqKa2lpbKlguix+u9Hy0YKifNhYYyf0c412prQeYKGZwVEnOTn
asXp6lVJWfj/F3gwWUoOpYH/SY4GTBGQIbZBzIk+7iitZRqGtNIAeDehj7PjDzxl
La6oH+3vAs1idAxQz4ARDfRBKkjRFGDidCykeJxDR2t7ngVXXfospiGPNdLMQqXb
DprgDTRlwHarRWD04wsgWDUa20yE6CgTRJdAkO2V0b5etMAAo5U3AT2V3PUky5oD
8mu4r7iCTWbLt4b4blii74ZYiHsDRTJoTlr2cs7dPnhGemmqCNLFIK/My/KU2oj4
iPM1Yi1xL2gODCn6j8DccVm7OxONTclKTT+MsNt+ZmC8KBNRrlhF7nQSoPFhhxYz
q9WMhPNNuJwSTF9GL8L2km4JoH2m/8MMVe2wIz8U13UXe37gzMhQy5bAdt82AqcK
rJZ8p56havHUxj3lQchD6jXl1EUP59jydBv01DbIl8keyTKL3dJMY96TYim8tcTN
Crc6Olveb/U0W0X3GJ+eRgLo0zfw+EacBSa8aKNs1CaGTCvl8JmznVM1zLvVqFDO
jjAZsh0/DWiH4auPj1j+IFTCElaUl9j8+UIYm4F05JHhg8Yr0M7sG29bDj0vnrFB
zZXvkkN54/VcLCIYiE4/YJTrAqZVqw1c+uGkmxS9SvE9sFUikTdqX3z7JQMs1QGp
gM4rr9Wa3ik6ew2SWPpW//VnV2ihgH+GxVCfWoeBJMnufZpmk5ZwmSqFzbqcUstR
Sqk2clqa2WL2fzdGOrBjffImenDtWN0M5mSmtchKA/bDvrsLQCE8tfEuMSH8a/rZ
ZbBbXu1ZJ3CgRegXk5/mUfTf6GeKcTy6Xn/J0BsuE8AlgU+IQ3Iq70JzCYF7Ak9F
5rU2D7nLDGFheae/YMzpjHaDYZgwWbr3DERrnE2rkSnq1CupZ4HBw/J8ueuz+jRF
w7ijIJativqXHJIUcHisnNfgr8BGb4Nw8Dyeu3bAL0TzRZth3a8RQ1mEXOXQdzeK
yxxootyGdHlARBK70EziLMYYt6pQtAqljbvofAR42frejMBy3L7dlUIJOIp7p9VX
XYUONb/CKchsmDJX5Ko5bvCB7UYPIl9ESpeaZCBQAqF0umvyrNA7zPWWKflKp53s
fCp2/AiUU/z0fBy3yKuG8Y0Q27LOLMXTKDFFmgG7y2Q2yqSr/QaNPXdUm8RCsF3S
z+t3GdzSCCR3zFXMF7duvHdR+f/7xFG7Z7kl+uhdfEZnC9sWWRtroi7yhyC5EyKl
El9672JJ2no2VCjb62D5LkPpNnm3B6fXnXsnITGuzlTgcNIKW05eXZS6MbSQDxm2
wXUNmqU0aTp3e+qM5/0UeEideBTK5ZJgSWovSqs+1aeVio2rTNk2vUebb3TySaGc
1CVhR4Y7MHRSuX5LC4HDIMfZGbVfkx4xZeAEeIDZToNuqt7KsSnv2dHPwxOJ2BDs
6z/oZaHat8DoXCQzQdpZ7trSPKzYuue6QLHWQQVx+eZ+RyBhBkNmIOfFwFXUYae6
/rmVizKjgHBYEjyVOzEKPzA4E7ZGfEczMEMjnqhL5v3ehgWuy9N46keJzECqtr5U
wu1xunE6ZVJBr0KgX0UT7JN/XdTjYOj1Gs6cBWqU9mDr2xlJQsWG+4ghhjLCTOGL
6LV7j8D4RYAEHE/OL1DkAEWBvkR79EdRFexk19lbzQkwyFJ6uulXDhWjeVF8aRp/
AakydlqW61IrfbGwlKUECjLd4sUZJG5h07HlgXrwHYQ5iC3dQzG06xvOzjW88HZi
kt++9uQpGeJqw+ZFSl+xLug83eNKoruPsafdBAL5PVx5ZVYPYP9dOtabWibspyJU
IbmEsgam8sGnwyL+ThaGIvw1e6SivIMFEUBuFTOEIAuLoNQc3fyBu9ULwuIz0Vcl
3KljJOj7uOFfMx3xSca2i39O8LDzMMhMJXeL5VwJYCfu/CO1QnqgoO9gGat2LTig
45qjeB+ky1X97L5LesEtXzSf3PC4EyszDZzTRIn9o3pcbo3ksOFm8ek3UpjXYtlS
5Nk5yjx5fzLLeSo1ZzIy3bQ5ppDoke+dKyRxZCzGuarr6CxcSu/V/6n0BVB4KVEE
FUBl/cJCtZ4iiIjZ4qc8s4w2ppEiXR/ZAZddqWrpKiEx2dvZW8hJEg5H7RZ/Rahf
sZKrRjN45lg7tEs2ZO39b3y+VdF4uFj80PKOGv+aS1Q12j+6XaHGlgFSPRN6U3VZ
I4Iav52m9K+68WMwVHmatsPD1EoHJk/E56NTqC5/+C9jhXWEm09ZqVWQ6TyDx/Kk
xHfT9QgvJhSkGxm2/88591+SqFaUB9WhHgK9hUT7cPasj3yh8EbcbdNy0rk6M0CS
lF9ehBdYz9idv8UI2W+cTlMGa6V+sPnXTy9+okKkLzCBDtmYgNuVAcRtfNHl20/D
DenMaFqFg20MBx/4GYrhxUV3WNtGTdFIinqKBDGd7/Eo2ZnfrxoASPGWrfcZ2IO8
CkNJz2TKAetEiM0YlG9BnUjjB5VGauzsPmgn6QVIbBASiyJuS9jdvTuon0qJfXwD
4PiGlbkUggKfGXoaj51lbnD2aMqhUu54cawicl4eB0KL1uRUK0H4FJf63xDDLXlN
VilgvVMkCeDMotMgLtPWpAxfGMvtnwB5/IKPCgyGmb8KydqRBZ9Tvf9jR72LJqAP
xGOHJZLL5MnPRCqDJD+L1rVZ+za2BUDosEkfeVYEICiqFFUKv6apwvG6kfcusXjB
V6KAp6geVfX5GV8+4ZxK+jJMmO3O1woFeGksb8FvCXPR10bQFNIdsqm57sQljRK+
WMwHL7bGapRcKFbOyy59ZmPHyqKR5Shf+0flA7nkGfejJv21ObJrAwmmoV2wEAER
/Y6JK5REuhvI9N2wkx3te1IatmXAI52RjWyS1tTeGakj/eUg059Py5WKr3nQJy13
WVis/jJOPD278k0WKuaRzcDBQcGu0AtQ2e/hm8VuNNcDds3J6BEbujkJhR5YwQNA
C8RHhAaFYH5htjOC/0O7+yqbEtnuPwNVOz+pEUy9mkQq5X9noQJCb7WPR6I9dRoS
j46TfLph9RwVDulL2ysg2uzlc8eU1Bu9eCBhfn8Z7YuA/pEoCxkRP0U856kibWQU
1RT4Obm3QkUFRPhkPWd3Mm1aAwi8VuTiM4wiRjsR/yUeEQQ5vzVYm2ZHXVrQDNVF
Y0LAgpF+AZNLvzRdI+iDIUcgclDF4WlZac3IMiRlKac8DSnXyZlQ6BilLCmv772v
DVsr3x/Xy7xV5dQGyeQ+Hnnollu7bkYjSqJHcC7VMjs4RGPxVGrIz2/8xvpsGwYl
E3Y3JABaRjXHPv3ro5hopOiHJboYTeqNY2e+7eZ6hLRaH5PfXDCWAQ5wqqflcwr4
QOaUuZ5+3/yQ0TH0aJzcVY2bTpAFjUFfjqWIXZl8d2LYWloCg3AcWkeNygBYrq4y
3tSFuDgeR8ZIvxYiwzGZJxOsM1agts9dTrHVzhtKPIiN8/wpjGlgh53xjIhJFghU
e7CYa7ZXvPyDYo+bYgeLLppeEMjRN8+zKI4STuaSsI2+FTKBs8desB3EEC8rgPhR
i5a0fxaACkPdpUNLJTJr/AIs11XPVLKT5QTOor9OxomaNgS0z8UJvWxE9gLxoE6a
TbdkRYTOW5EGZr78IQwVo/o29Dz+L/lXma1YKrbyOpFk81tzRAnCNoDV7SNjp093
aQtVM2aAGfE9ekhQDaKQtqA4D4vov2Evz7mRt8rBHO1QbiFjT/lmtp2V3Qd1guX/
3hCNKHs5bnvni+404dskK4EMkDx1gQLVnphRmt7RObY4tQCQAw7+Tt+c44JwxDUm
c5K20+N4weXmJnZ5oD0TWh6A859Zt2vc2pY7a/LvDAVNmx6iXTWZ0phRjKJKm0eK
zVN7C7EAb/O+qPZ8UmwZMW13HWjkEblmRkvd4U0s1CkZGxOJxueiLNGR+70fbGcI
tNkUDLd321QTsG8wU/lZXJOiMAKQonu+lFaWyismrv4knkUbC9QQQN2I/1/IIGoL
gCIk0cQzLWarYm7NbDxVkxKTyy39UtDmAEblnCqullwEQPIBJ2kUlMNVX4/hJNN9
sIezqFu0dIUaD36YL86bLAhcjmnBDBhkdurJmWCwa8ZCf/R4dfW5BqkvX5VFSF/6
aPJWNdQyneVnxJxjMaysNz3Da3Qdx8L/dNLgrYsX0Spr3V13iPqEhpDfnWpsOfPL
04HVxds8KeDCh1VMN/jD0B7IuLQ3TPi/PH1RaKJrCJ9wk/D9FzcLpSuf3fi9SF39
VGkQtC2WuTGCf9YrWkLqvTyXMJQ9NJMD4Jz5TCxgu+eXBKxLadbcdH5ttI70jXM6
iVL3qQHrlFU4uAqVlzt1EV4UraFROuaKgFnOnBh39aAkC5qfy8OPeeN22asst/8q
5nOkCMHiJBz2rcz4VwDzYEbBQ+23RisMpM5SGThBiWk1kOMDVnQ2fmadsnWtCPBS
UY+cX9kVXMyfpwBHeVvW5akdgsOEarbAncvPUzysNyR7IQ7rKr6VmCRc2/AovtFN
j/tEY6Jnhbhu5PWVqCfueEtZF6Rqe7eW9HBXq7Z9TPHq7+nA/4lRir4gqp/PRs65
rPmkRjRdQ6nmG99pmINHVDe1IRbcmNTUAxHuavrgXITu9OuzaanmgYXIdRSqZucr
gXC9ojI8r6qp3PEjwuZ5rYlAzzYBYA+3RMz6mKvb0LxLeHWUH3IHvH7tfwJ48Yem
Ij8lDEUw/Vb5O/LSWTz1SdNei2TIe2SQUamIhFIc9+MBR6vONvWUvFxf0FGryBNJ
FRKgoUrcVsVGQJlI4patWXVV4GdijnTYl3/TsOjksXH8/eabGL8IOpZ+/zupSRgz
PKup6h4onc4OTe2JU/47UtMhYfB5lNiAHm557FGFlVx87KS6G/ML4gC7cmm/ZzqE
npDjSmQi5/sbIrFo1yBDLvoEkidYkcMyBs0RUsUI+xdQj24v6bgEnM2GiHLuQmqU
XtzGLUUJhKrTSR1Nyq2qxfzizyg0ULbFeT5WxqtPGQy8CkwmgMsiAFbHx/HlEo7U
CxECUzjcH2WlWCSWU/MLOqod/Tud1cuxDPKaCACbCqEj81hViVnFrMVHZRC0KLdP
4XoGonMTRWC1ZmeytFXhtR+Ay5qcPEfx9D/oZTl8lvO6vf5D+WXfyXEGc0g2YMjk
V3i2hGy/PIwBc7ieGPGEHN6TcKbPAgJvDo+cPN4yyAnVAKoRZpx0n0uAyxkllf/M
hPj+JNM0G66df3zW4+SQgqBW77uoRkY6jr0t30+ZhpsiEnlDwu9p+sGbzI75wPZD
dfsLWwq2bFZv2iHmSknrVexn4IKFFHvyv2FceZWKtHoO9/du2Sfrww6cxlBaMqA8
SeUm6VGULX7LdvMvYSNse/Dmzg4JTxW9gfVH6hc70OPtkTuY8XiVBTuR6JJp42qr
0Oq5C5OwWwJi0EVUNF3ubAM+DB432tAEYwdv7cKaQrPrBc5IIfSVSubWFeQRHcJm
OyX6Ak+9oPnOe06ZtKOor1hRc/njGy07+syRCwl7rLxzLZ6l/ik7NUQqSY0S5JxS
obMFBKCT2ZI912ZSoEDMZTaBeA3VgI/Xvt4ue8igOmpStaUl0wl1euqVuCVRrrnI
qGD722Pfy9RWKgmogFHx7rYIlC6TED3almOftJ+52YZGRqQzp2V35tvbFXmNbUSQ
l/k7ya28EoV7vGFyyGazfD/Ms6+S91lrwQEHPm4QgzLYeq2bOIeO3aUZYQsLom/9
sl/dEY+LFTTzQ5oZRQUW5cu3jaQuV/aHgz8LrS0Voeqzixl+qW/sd4Z0JeVBbn+O
wS+HxycVR79mxH89283VOjVDI25DQdjCvNQH43yPyCOj7KvUfyfSCcpEHQOo2tYi
nBaiBfRXEsie/K+lUvl6i6hy+9GlT7p9QkarEKb1MGYLDCk7RZbmxJtEU6r9WgQs
PfJnYkW1Hj9sIzzfKNddrelUzhkIGsW2ClARyzkjEVsbkR5dIjwbmadPmUDIu0Fx
IwDsOykoxR40o+rAQW+6BqfTauCdaqCnuuLXhvNaV1aQ28UTgJJxYYw3JfG71YRb
5zzOqtn3+A+V83ARFGMKQQgFBN0HxII51IVWLTC9sezkKfpGh+/rPm7/yFulq7yp
Hxc38yKIh2ITL8/7afEnTGfgP15U8mKSzGPxQ0pdMVDnZbxlOYGqCZ+DsNLtExwA
oOx4bYQynFqH5jLGSImS6QqhEVrLP3VfS7Ju/Hb0UsF7tYJyOlfaIbrnKp8kEKAk
FBEvrKZTK701r4hSAVkbuwfmalfBCf652InEtJKLjYueJZy9ZBIXB+U4RqwpUXkm
uz6P4BBOki7T/wNYIY+upqU4FA7bwWY/RcqSzU10B+Q2pDsyWQxvbiugmCswhojw
WbYYT9+P3uyMmAOji1GC6cTcyEp7d+kwQ+UR9dIpsSj+7szrxP0w/cuUNJfCOPJC
IJ/qpPSF+6tv7GU+D11E/tKwefkZEtHhu2W8zx++i9DvEXOYpeBUegFgsve7E7pQ
WOFXYoukcPHSYaXYr5pcF2JQtYuRtmn86dWDaXDK9RGynNX1zMGnPAlZiu/jXpIQ
I7FmDjlBx8WoIdQtul7utxO6dn+uKJiffQ+w4IwZ1j4hg5Lsu0+pcdu3oU/cDvqA
HODbGXTdCfIH/jHMP1DSONa6nku55ZgmuRvCXKcQcXQZRpWy7rsULG/drmYfwiIr
aG902Z4BvDuJKdsXuv+fKocv0kwPR51xS2baaAF8FdTfOnkhUssNz5fCrktTZXO1
Vg9IJXLI4xLunF7EuFhBjMrgmV9dm9wQyzIMgLrynFGkUbIjmNvKOsAaCI90nv+y
Yt0FxuV/iBzEnFWujF7piNfygGHKNBZRZWO6iwx7ZsLvUH8bDcO87/D6JEMjbw7n
oLuypk4F87ahr3cYATI8fvcKnAdx3sDyMWO47iBFYk80G+EKfoY3H6xlYs/got06
hraTfFV1kpITldiaSK3Q4cWe73ab1ctosdCxk+L9/5swJmez+hrvG+EMW83mj9bK
AHQvewfe5z+LsO5NL0LqVhuiKCy/qCKU8zoZvByfFDeikwqAeXS17aew+q+5taRj
+zPgM4uHr0k+Ob9cVm92FdXZA9E09NJ7oSjENHLPy/1pIDPGJ/UzzXXUdIEGPumV
bOEJ7uX7RnNU5u0WwmJz3mRDtToE5+A+cMvjiH+xQQSYqpdFVnOj3ae6WiCqhdxE
snhiDOSIASGdX2ruVy6LfmDkwP4d8jBQj/ip7x4bX87S6srtxt1gx3LtHW6g/rCG
VciXXLWNUQNGV05qJNiM92VU9ScckYU+zRYcF54RnsDgfisN4fR8RkI4JJcH0JbY
bwbQjon6eKgY4RvDQAmwyrY+nL5G0nlpsDx6o+Hb/S/a8lpNgdTu4wZyw0o6s7Ic
Z7tKAZGlHfvhxkAAHP0xLkgNXEDQ2nC0Do8YDkvaGQ6E934smJXJ93ZssDeNhWPY
rnXwEcmof4SXeeCLVQpWknN0lTroTIuvm2UH9UVdRWftMKRTacR249Ie+oN8bZXu
Uz1GyYCUYa/SnFrkapSZTvVbkOwhAt6eee6FaYz9JiEQyAo5E/vnnRqUof6f8jfv
6soppamAOS5tTmYC6K1gwtWqjBUFpnZ96dmpreGkUzUWmCplqT8riaUsRCx+3A23
w0rzHJOw654lxK2lZ8Bb2is+B0TgSIXE8GEHDhCYTTleVrQkCtYKsF6vkzOTDBnN
/o7hPUd3KOL4+VyBq/BAHsAAoQCu1QZI1H1zOOPF3RcesvZ59mCwS4eauuVXRujA
1H9KLo+WjIAdBCc5Z5RdDowCoybl6GpEzScVrzBjvKoFIEL+3IMZquqEM51kVeCo
oO9GiFtcdVOznMHqk4lTeDCtr1s1yumSWYoM7KOO/qEhdX7RJE6wkL5A5eZEspOz
cNY9WmBu94ZIIlbi4YpJVq+RbDX0Bo1KRUFTPOwhkvH7J05D2DtJ0srNgrVOc+6R
Og/sm3viUfxfYbMZcMp5knnGmOIsSkU4Nzg/iKtrBpjBQmQdVBi3aruKNLADTJKB
FbpL2WaxijN1tsxVFD0lroQAEk9OH8R6cQAKOcdcQVsSB4GorehaG7GRlm9FwFFz
5IbP0Qzp2X6TlNY6wcciPyuyp1/vhw+so3PRgQfwB5JoRMtVzn7F6WEi50038Ws5
uSpjXOgCfQb6LNYyiFMNNYuNPiA/NY44/UHYt1/jZmjwPKgSCXsMXTT7BbPPvRdd
SyP5jSK5QeMiBZykhwJH/tNfirdNDtwK4OJuJaQnJtcUrSjKbTr5QNwFuUp4XNpX
7rqO8WI2HIFHNRCoqu66C93yuZYCIu7WlPe7Kvwq7PVhDH0pGp8RUHsCyB+4992U
CSQ22pdETTS03IngAJk+S+xBO1K2/vRK3cCu0oje4ERzsg9goSEKCMbmipuhiCrO
evyjnsrnEPmt4/mI4KEDw5IrOIqBKNBvk+LDMWk3ytdRFOthdD2BoR/TwAMxVl0E
s6YYln2kottcbVAq52M0X9SjT6sjlDuNpelwE18c29kc8lgRsmVyo4uXkgpywNko
H+JMXLU+8ZXZI+X+iWkfWB3OH8bzVsrWg+zu1zk8E3IPni7hjK/dZyPU9BZlwpy1
DGwGaEH4VuXRLlrIuPhbLyG9yKF2ZFAiSjcu4b6O8pgUS/p05hvQsNNlqF4d3rNT
kiuzIsFaKF2/0MDlOHVX67RiTt7m7q5kNLWQpK52H25twUSVmzMb4Rol9jcSU/5Z
9Dj9MsV4IT96bm83qmWI+Tn5wwsgo7QBrUiOBAeypZGeWt+UcbtgCYtEwkUj3Rio
nsKF0+soPp+urvItQd/HddZtjkV5s9GRG1OD+7ja1srpjC+i53K+XJEtLfKDQ8P6
KXPyAlW7PEl8pi+gvO0zbMxWoTqY/l7vO67Zxx+sbQ6FGRRONTyX/wpoM5WsxEeB
dDNBzXTKnck5yAmOxJIdwYNwQYmXvh5s7fv4GnZtug+J+yQ0B0dW2ubA/Hx62YaP
A2kES7ZbzAwWO7iU5S3Hm6zk3oR4wIbWDemP8a5Py3XIIL4o2uCAbMXlMXPNw4x7
oHzBmyaHJHfSIE1kOWi4WmvnAfejkqlHmONEs3i4rAM1kCsDwAlhpEGOXNbaT/az
kZ0MqcysrroN6zdF3fTk+2epwFIfGogBTVI+CwF53ZyIt574A6PWdAKO2gjVX4OZ
Z1ClaNh7vROnit3aqW9PWoq6JCO4/M+Iuq0T8qAWccq+VLxX//PhvzhiphGcKDOa
IyHZ9NfQjuZ0tFJqrXI/+X7oVfwErGHXG5CzSrvfSn+0KKuaBOkIGQq+8OGO/E/A
Oqh9Rim37v+MVcxYY+iifJEeKgZ2EWwl4AkHCF/hLy/5Kk7BoiKgmmgK/i0DS/lh
BUXsiFbeaxWRZCTdWbRqpledHX2oN2l/rr5KhdtO7rKpnuWM8dpx/e0oDcb2+OgW
I+gPoqqjV8jMgR7xfQZ9PX3HyJ88O4QY39U1cyXnFpH66givZjqjjQV2l3w3dbyr
b/pFB1xWrGUBcUvexM1Zpl/BeWbU7D+lP3fYD+/sTgzpjO/L65oFC7MpOCQnXhGe
6y3eIOjSnagPLJlYMgYH24hZfAMVnsfQT+ERbQXAMUYFPCdKb68SlGo261QJ4zV2
LiJLloh09oiB+roZuB5EpfiXLeztb7lXyzVzuh9AHwdIlk3ITSWO/IIezgOx3zpS
VjJfNEbOSX293xoPmzq2/TRFfsis6Ou8AE+co6CCDeCjWu+1+tsD6a3443gco49A
ewokR5AYcmvM7BEEpp5JkcVIu0tgsTHu76nRxQg0QrQRIhAKeb5/gPyMpTb4w1hb
HxVrU+F3lRyWr3foIEEgamKyxuAfNWwCCAhbtgS1z3lNptpIVguMbsGvzfCa8WnJ
Rm3HLWr2qMO0Ko7kugTgG82fSLG+pEeerZMEzu0I2UHbxi/9sj9ok8A3PIjqcn/u
FWdpsliPz+tCVKaRlikPu5kouA24vJ02ThWlOlU57983HKRYwkXc+ploL3xj3Nxq
7eBSWDwE02nVWJp6Ft1KNsqYjwZhrZDGRiPWGvibzqfPwyHDt7VbQRmvQvwXsrKp
wlB3sUXIkxG8kkegFl5mYfWMedTQoi1Agudk/g7Cuy98QokQyPEQDIKp5+48vXzv
9wVxRSYYL0FXmuH2YenKdDeXiEUtP8Sq8uOmpdFomfWo6/XX+KU+cHhb1vov0WKW
/cPPC1yxXbV8VVAFOKpTIf9Yd5y7sHaUDGiq7Cp/kazwhekozy9tSpmhgXAhPuqq
1PNa1WyjUW3mSHX4oGlc2bs2+quh0ZHRPe1stcJmxR0y5qzA8j3tFb/GI6JCry1r
9n49WlgsuO7csjSj/g8oZIg1ZP4tMUO49x6FH5+sW4a6LRhiA2oi0vhBJe8vz3UO
9uSgKr7FjkmUu6NTe6S8wZCk+3e+QJXsjouh8hEdUswa0ebfHqfGn6/4lGQEPzT7
pHJ635gNMKg/JGPh7t30pBPDk2RJmn6Q1pMfIS/spTDKe6wRXN3elxkVmx2oN1OB
SAlYmwEjxv4k6qbuqGr+lmS3g6luF6etFgSqRi1P8qdO7MojR81kUFugs/W0AcxF
rhsAElGcnsvFVGSAqA70f+BISU01DSjTncuEELqe6xi8ImkmuivV7sMIaPKW+NDA
PaPJ0cxa9YPa8pOM2iCTyar57a2ONSeuSq6Xe3zuEuL45R0Iem1VQqUJJRhuCXRC
MlpB19ebBSEsFn5Y9FkXq1zXWE02BgQUWmrPHvlM3cMqfhEeIV1EOOSJfNBoDZA9
vmEc7HQbEMLWNNdpFdwWOomts9InLKIBFrNk1VIMCF42q7fXN18M5O1nJAEkTaMc
nGVvbkzbv6x0/Rej8vJuPyVS3tm4YXqB/6YQhb+PFdDSq14WQvvhGO7DgwCZH6+F
DKYD7QcnNiPUUipkU3NH14BZYxl+OlcxCDldcldKQUogGvlVDcCHeu+o0aU9i3j3
s43MMaZBM2s5dflo8nnylgRCP+SQsL0JS9YHTqOz4j5ovod+TM9f2oAYrOnYcPCX
dXbdaSvuuAqtyoRjCy6I3s9UXQtAc0/cN2Koe5DoKABcidIgNsxFkWARfQ7034Ta
fr7NYIibfQy3uJTC00mAF2sFmFwk+Rnc2vmI6LKy4hMFKASCbDgx6DjUC8ke1g6L
5Rrxge78YFsm9uXicVMHQamjwKzyKN4AIlnuRt8xNxAGthKAyVbswwP4kjUmhW0q
q8TtbtuXHpvupTkDkMNuU+w+x6ymCwUaaCk7JuXC/mbXebZA3l73CIkk7UZ2Wv4J
Jyk5EflyFbGrvyYhhkF10knaNpm0tRBKlCVAoaHS5I1lhGiTtg6lui3x/sZvjbtl
XZmescFVE6hQ+LqWhfUy+LDrYs8Q+6lwD+x6ngqgRSub3E1CF1EmZclQvyBN7thO
vkIs8vUjy93Gmn8zEH2KAuNW+r8vfXzD5nDWzPBnR1BU1hmwcdzLPZK5sN/MFjFK
TBYUyCmIEzezpIVIbztI9u7+vA6y2ZNr57r1zDXEW1uEWrug1VVD0tE95uJtsu2n
lFxGdqYu9LeHiQGbWA5IRYZWgOS27iMHkBNDJ+x0RMrbT4F8u+ipHZk25oVXzCW5
roitDJQc9HNfSb8QUrEX1A1RJZwti9BqwtLqqduuZxUd6qU/jExUbLfI907R72Lk
Hsk2pnsl82VHA9KZd4hhkndj/+mtXSnq2KKHav7ZxmsS5ObmFSaGbSdyPaFHl9/h
Tfv/+Qy+ziQ44dsleVc4uh4w4cXiiynW85SRbMAEk4RT3sFDozEVnOVxbiJ9PwDd
kwtwN+8MqPpKEixt0WGphwP/nOaoLeiqbawiYAURx3IXWKV7nSC+gw+AohIYksHc
hZDhk29dVIp/wPVbFgA2OSElPhVmtFtWtu/JubuzguPf3ZLH98+tUlRgrTlNQSMc
+/r4U8fLzwtAAjFs/D2zdANnmDmssmNcSKW2GsYwkEalzzGa4P4hCQcPQes+Mt+z
enof8DNDFUOOS5ray59SxkJTD2XSucz1KIAYJXFRckM8m67R8ElU5IM4jmv+41L9
dB/RmNfS/bK62ult2BAah9l9AJ6ADYZZ/MANbupWiCQ2cbJ6rjS8Xj8zKd/ZozlR
RD3cyYSMo/Cu37k+tBykhl4g9FrOMGfJigdC+MGC9zNcKAwMA4iO4HNNABmGabAq
JmC8QG/SbIAocc4QYkGAeVAoUNSUeTGLAlqSSjrE0NicTLEpljgfch4yrVO3I2eV
6HKqYjsI3o0KqvVB6xQ7J2+UkggZJGM8LO63lZjlXxJ7fEaNBLBXOfSnovc7Cut5
0Mg/OA1PwqlzFJPOdqRyoA/4PVj5+oA+8AjrlOblHSqBbEsHsXJwGYwOtzlnugC4
CZOTeaVmCUnZ9jwuifxyDos0RBjbj6XZcl5x63noQR2xaFwrn+y3ZsB6OfkVEHBK
CiD0u7IVxLq8t3SbOJJ39UDjkGiGrIecqFgyg4Eec5negirqpuBor+FkxxRIIDxP
JcVFpN2MWRgpbEQFel5DiwZqYcGl8ha6FgpQaQeiufYttpxCaTn+DZtFLbzb+Nq9
10PqDe7TByQqXnrsup6hbv41T7IAFLQUpskyGB9QaK5c89MdDg4cvQhqjaoWttuM
Ee3mxWkHhYG9W1aAUmd5M1MplkO6b0vhpgMuhOJdk53IPXVzZi/CCUclCVnwA1gH
8fbbPwCcpizUEFNe2RSpgHd/83zyGz5xzAURStg4+ZGij56ML3K40x+0pOJlq0NA
9mGHEtLY1mGP0JZhRSx9s5R5eP7RtcMxI6g8evFurY1a73lkEnUdxKzUKycFpIOd
Ry9KVPkDLC+zRRJ4U+UBPDDwmwpTlq0elc2tCjChGtJ3zOzn9vRjuh2JkGLFJuSA
DSWGyGd7K+Ht+Lj387IwF99Yjwbx53nBgR8G3WN9WO4L8WSeYlIOO698dETqqnsR
zpJVp4qNFDIrpq85g3wYRnCD3D7s2ydnROP5EnedueZXChpyK2D9TpIS0NEznUYv
QWVpqBxm2nesVCYjoHUQNPwZ1Ka88hr564TvJaGTi/TejFIuN+4qy3BcwOgUQdiQ
56xJvYk7WU9TC6ME0YI6aNlX4FauJFAzGophfDBDNHaQyEWOWDNwpqJkCHzLQTXK
j+nN6nDrtMfs7mqkszwFZjgJDq4gXgnEj8Lb0DrDX+Kl7RRJ3gunVy3R1teYsheE
sarifnGnfgB9544EP8QoxvafW64eaWVuupXw0uBEw1ovbxm5+5L88ZETPcF9AgkT
WVKx4J/hU/tgk8ED+asggk5fkcb6Akm1uiIw2mbs8c3bbepXBVr44rrzExyjNjrB
d5pHSwFTvenvHgVSEgMUfSkQT8UzqiOjkbHpxyQWveVsBqDlNApJggMdI0IXw0oT
x9iSkvZ6vgwYLIsP1T6JHsKE20vVsuJUy56WXcxtTqjmJh6SHkjnWLUOiiLc7l9i
uvA5JUvwoRK26SaiDwMw9LELgAHSiRn4vg+kcqYOHBgRLYNKzlmo+Xd8fVeJdEyt
rg7g3FO3JqMa/KmZSvA2K0yqTjug724x3SCyUYoo64CGUOg4laN0lAcqH403i+Bj
dVH/w0ZePaa7yvMLlLVCUZVkughjQwRHRA5AzJn9Xj+rh0x/1XKFxJuxn9C68p0A
f9DxBZOFro5nhOd/VEkmsoUqIl6RurZgkP7aItaeX5Vcs00/9bdIR99fW/mEQ3G1
yyLv/lvoverrIQewKRcycPfi56irgRyheqfQNvQNWTxY/r6yJwUCIzGgJ0viflyp
p2kVYg2I/UGPq+l4GLq1IRQFfwNCjaxVCQmbbfWOF2Xi6ziCM6CHx5PGbIO9nwae
itEMmVdAhkk0JBSwsJwwOIqRnpz9AwR9dBnYqOa8ed03XQ5v6lW2OdtcQkvf687k
1LyNa8hMLycNg3plV0tZM3XVEZsFP/J1PBVRZWtlbc1WSbbxkJk2dyPu1WFA8vdM
TA7OzHYir4mr6JSWxHRli28Ru8LsGbTX/zMIXP7D4B5X8PpEjYe4NWVqScIqzcB6
lqXoYKOvn/6+DCzvmG9wGWF1AEQcWfSSBlVSU56fAdB9yeSmeUiH2y4zHxXerDbU
OzWJaTr2xv7RAqMFFIhPOdPM9cw/c7jWdP6He3RpN1Nx+jySAA2+fExNDdWgS6W2
Tf95hY0upb8dz+8f5XAfXGNuGzS5doPA7xqpSjVWxzPwUx/Ee1Vg7GNv3ZHohisn
1mZZDFXoRwXjoHJk/qao8VR1vYXbQQCEiHvgJmclNpWiSYnrYydAqWJwIavHOnGK
dEbm3U9BIDz3HW0hiqz8fkFoA1TDUHNyLxDkwKubPBvpD9upq9wdKp3+qfyyvIOU
kx2ox5dfI+6wrM8D/tJxi/H/O6gRiTq7UBm42Ue3yVtoA1ieWL4OVRBqu02HORHV
vMC5rvVacv4oisnJtRFwVJHEpcl/kk8zIlqMcZw+3InS7HJhwvPFSFuTk/633EnE
lGE643GoTKXZTH55Pcgu8lXQ/o56zdJGEOmcB3zRXz3+J4btequqQLC/PR9Z5jSK
iq0ohL21bw9fwKvErfcJ5UfEvkoZWhpR0PJBPKs6dk7C6U0mGiMO9bYJFDsarZr2
9CYTNKHE6Go+Ftn+GlTh8ve3Pr5OhoFPq6ZuCg9zxQUnGqEJnrV/xgxPtbKOJHAj
7GXYzEsvTPdA0mNvDj4+S2cSWrzKgYevnCRXNaU2lrnnN11PRgce+p0KyXt5ZAyT
waWxQVglU4LWeo+fP3Q7+9jp59iA6dLqOC8/ox5LEUlQ7huKhb9iL4zdckGzofFW
5osJZyvkze6KHzbbTeVsMCY26f5J9qmvpRmlmkm9BQ0OVcFNLGoF3pm9N1qjvBi5
UQGwg5I6Xv/NGUQTJ+jcrqIFxSJIyrpVxDRgumqpNyRmqL4gj1M7uunKA02GZsCu
JvvRRaMQz05BzRZzNNIiZnBbEsV1XS3c8X7XmSYxrZqyqWKy+WALlJSN+O7FU9FU
0PSA1DlD5k2zx6BeVdd54iIKxI33PnMl3AyoKLRMMffAyVfaO27kBWg9Vlw6owlA
1KtNuHdaE1XCzl/SrldC8gvxq27vgfmT2FqV2pd7U+PnX/1c0PqbWJYOJvUYKLfs
4HMGFVCBnmz1eu1puiyRMZxQtG5xsowOeUCoSLOytwsyHE6gQGdVdpYJpUtN5Ldb
swZzoBfVP+SJAVCwpgqNCYcNLnOOI9FJ11qSkINEg3mN35jNvL2sja5dK+hNBFkF
Tn9hNGpZhEgoAzbCgM75yochY7HqkJGEOj9LY8Imu6sfTmHSwpDLQfEWdMKIMIJX
FFfXIpuKbLJZqZ3C+FGbc7ArWn8Pz1ZTlEhZyJ2itM9YZKn7uiVSMhhSGs3wk+eE
pD77d5rl8dlfchN6aZXqCGaf8GNRAo4MgFFq3FfDjgxQD6gyzDoNbedUwlcsKEqy
UTboAnTL05Om5M6TiyYOJpK05WgG8j3Rou0sP5NE1FRmjfV0gnscMmbz7KJFRjl5
kLQOFfPduO/D6GZLBcU7uZGroK6rC1KSGbMXpwPRG6Q1CJvwuY57qemq/nS/MrxB
OBTYSMMOHYZAYYFC+sOyEBiq3mQyfpwpJwSwvwmbhKMQhTdA7n4cdqxJ/8W6z7Qe
4SbplmvmBPKFKZvt+sUHGYQJ5lURt+kQ9vzlQ96M0+LOdh5lYjXVk8qY0AGz21wk
8bAJ51VDvePBuOcEpPyHU607d+Np/M6ZWPNGkmmEvAfFWAZedQF+euS2ZWZMqDXX
66ROk+AOb91HYiJbFnMSlehSjRMtKumx1Zv3IbuhLg/AlXfpjiQkpWwbHpONjvxb
G69BXJv0gZP9R2iZOXENbFBvE/IyeAah+B5mFy0NHQZxuJGMIAFjGEBVLV1p1cYm
hfNN3rZoj2QxOjuSrs1ooYr4suV93QyHQYbJv8T6ilibDVa7h+ZMIfc3h5iw4iWm
gQQ4Q6wJ/Mrs4dPaO0luj+IbETHKMk03HG0Dg+Kw+Qa6FsQMXOScM203dGvvAKjc
VadN96kzQ2OEtbVrPQ7QKC85sRhNx3G2CkW7KOp5T6UeOVJO31x5wMWnYMrhRqy6
VlEBJlm1+Lv3eLgUpEg/LDXWEuvLpsj6oDuw5BYf7QVHEoUNMQm+93KF1ukidBKw
ebwaGvJRShQf3Z5T4+kKGgeLJN4ROEVw+5oMSQtlK6/Fj9cFk1G1PyqyczRRHtdf
VSthAQbQzbJt/PsTMYsEqa//tcePKI98RVQgnogZhCJ6XNogBixpSzNBk1WHexbi
xzdTkC36+vO5RMaia7+cRYbmKlzla/YA8nOjZ5Qd17cehpKA3ZpnPscTuU1bZJJ0
atZd0N3p/EjqOuTKuXRO8STYUHyQS+UYgEw1bnRXEkJX+4fCqssKjHt4Ao66kHIF
GeXT7CAdSINXr5E7bq12g5p0vhInftLJkj0qDjuwEAUl8fwlDPT4+RXfW3RuPVjo
d4glnoIyIRtB5WV2A7c9XhF4loE7U+WovDpNU/wsejxW6TKlfxMmjPV/nU8XlSqa
a0iXKRYGG7a7LWDeGzHIk6eBV/9LXHE0ydEUILRuDWDfFalXx5XQDcOVvVW5bWOR
gye1eYmvOERblE9u4pLsosx598jnQ0F6eortl5cFv4iHL8r/OxvmbOJMyYCaOV1C
zp9o0dTnDFwDwRnrs7bEOc48O4edJBV1rqLD79JfBaDb7uQIRZ0bg6ym0YTog6c5
ZcSd53Zt37gEU+3eKr3StsZYwdxxJpxbexCrywke2ZUJRkj1IPICt/RfRdfiF0xW
EZREbG8hUMYCg/cxsXIcNTJBQh584tKynSRDd2IlfZ/sq5fWFckrscnKvr/b4SsU
GdLex9CTBrpIqAyb2b1JYItBZ+lvQtNYZ/Ly20sJPVwF3ypSdoYpGRRFMlpVi9WC
liXDt4MetTZ3m1Hvqh/VhXF5odVSD2sg1xdAzlvDf32CKmYwluceGzoDh75IpUfC
GsaSCMQ0gua5n0RHXD/bncYUbFI7VtWNjoAsnlVUWosZK3ywHIA9WynmUrfCQsnp
u56Lx78RvjMQ/cDEZfUQQJ/ge7BFUu1OPDBFUxMyoF12RgAvX63mf5D7yUFQVaOf
c+KktWbnw3fOnw4WaUbswSXcrsW2L3Btm+e32KaGg1ekZ3bhiols9DI/P4UQjv6O
84gSddZACih5ln0QiwQv+G1YRtihCpb9gXzdO39c04FKif7+WqJFPTJwEGJ7aEmo
xlPsY2j1J6wpfYT7pK1YzzTztDGl3apM6SZSCnGtGH1y2qNe2pzfHcCCN4ijLN+n
Z4OkNxSHQp4w/131KkmvWPZ5WRH8Ew/d6msf/sQpXaTAVzoyk4BZy/nUDNFUecO2
gRNxNqpn9jf6strDlat4Gt3p4gUZuhR6K8kYlMl6BnSk/L8nMmmPsJA9TllA83BL
9qKk06vMmOHhzmT/fxjRF1mHql35fzxdLXx4RxfVHlE01pjPay15HW0e3SY7sWXo
0Ka8lVuMCkHPvQsax4PQuCd0ZOZO9bFkrAjr5W21QIENTGLKsJpWy/za3fBSnpYe
L+7GE3wCBD2l9ul9RnAz8c7A1/n5WQVnfPRXA3laCg3i3Ka5eiPnGy92e60spwZR
ofDwz6ANuYfnznqt6ZVsuuATXPTsFJAo5CnZ7Cd/9GwMTcaJq3KUpe0OsmDZ5oB5
pIs9jDk3uLV0g89lu/NeCC5da/i3mTT04FGGbVDHb1U0Vs/FwLd8Q3y9nVT2XDdM
aKAjSlQYvniTvrbJIGtoKn4M2IXxF7WebjYli2XqCArKKbj2AtQsmM2GHzsEyFSw
/VuYZSjUiXBqM5a+ZxuDI7Sttr4iGZ68l4WrZG4mox0EZ9MWdx7I/k/8DLVzS3AJ
xeBVksGicD/Uw+pULIsBDURRn5W9/8zZhY9zx6PntWCMr5eeVbntc5PiaGDrROrX
NES5oUqiZ84VSdnkMZi5bnt2fFjT72d4S6Xp7lHckS5PPjYd1GYQ3+O5sOUeohC2
cG4tF0cqnjoOak1wxkiPTDKuY+m13lTcS4KxhKrNyIB1fhRaWKJoYpdTe9ut+o7C
kVFCHvodwdAjquCMgbz75l/+SC9bgjnY3B9njpqNJxEAClGz+9x/EvyCOFYABXHL
dOUKAXSdwavq4+SUj/BNtcs8S1pltPlUY2XxgdF/J0OIjSQTuTq2F5537sqYH8/o
Fpr51hXgJJFb+eLw8Ri63VB/zKrvV0dtyMVtI3873kcNDff30Kmdky6n4ZuP7T/l
GZxrYMbeSEqtpDKx7BP5KZpbvxIJZjS2L9uySIlqa/IjVXaptRim4o27i5Vqw+EZ
/PX4DzikbLtjJgad2dh7IcHmqAZGvJ1EAsjv0oQtJxORPNyfMkCz+Zcxa2jw/VAQ
QLEmjGK2Jj0WOhJ/et7yUR8igPsB3rMJ82tXNhy46df/VSvJcgNEPru/V2vfHnPY
8GAFSnFSPQEBLIeywzTuqANSfU0N8ttwyRtxV3v4hj8ojizyr84Rpwzp2ZkZxuaV
Tv3Mhd9ERLnpVIUwABGrSD+kCY0mZX17T4wBWaAOuYSh8ULB2kGBaU8D4W1mZ8IW
gennOw4MaRSosafbGSsqZnTA4tsGHMGZ8xcTgseXJBJ9eaClTKYtYqzJq3RCWL3d
M2BWGmYaY7egHXancZoH4PSyoPhoylv3vbPye/06E+Fi5LNy3FMZek5agO3SKN2D
NQwKQnWaB7gge2sc7YJZo1hTzs42V2NwRJEOQVoGLfEa1UbTG7aemOSM+4z1e+0C
kPufeuLRpoZCo6jjz2UGRjL1SvGp6nhGmtJe0mjhctB95pb+Z1Xl27+p2F6fC6C3
rysgEOxUjvp/UVb/TDonE1foQriFXeDt7QHkmh/8+dc4JarDjndNjShGjHOxEJ35
R+c8k9frqcHCS4DQaD+Co2xLjK7v6x7tpnhhXJzZ+zD6OcHflTG9/8MTtNFxn16M
AOVe3orofagh+uHePB6HU9EvWsnL4ls6auEaQWN0t7W5/jWjXZoVEqpDEO18JzbE
wF4a/on3F58OkydvePhKeQ==
`protect END_PROTECTED
