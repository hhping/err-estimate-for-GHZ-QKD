`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fSJ2UOlaBILubkvFxAh1dY2BUJZX7jLLOM6spSqnDri9uAisAS+j1YIdA1UpOUEb
gkZdyo94PtOGSIuvmYnTAZoDl5gW80RupeHD0Hm9cDJLdD5TjstwQaA/rdrMoexb
Qm3SC5CJV4dmV+J1gDWukAe1Z8kbh3594L3RTdAwM+vk5je+D0sD8Q3lUGbnBP62
LbdB5YEiQcVS0XDL1cHPDkqVRw7s4OgSb4gekVV200F4EfGngshZabd9ocizMFXk
NPw9+XpfZMnd85/HA+UDOFd8DuPbid4lcxV48bk340t3XhmkOWfIcz7lXqhxzIj4
xwZ6+B11NAUlsgwURl7SENvQBg3CE6J4kTlBG+mE2oTtejMD3nmOB5smWB7KiFCa
4aTskbJaCJGXTLje5hbAiUNeomxOQooMdD2gB3PT4f5fP+wyXJChh2yK4G8bPJXo
BD77iOE2nRGu0zYpK/1SlK7a8/wIfIvsblgn7SoJYjUg/CTiiHqj38o49cLwTnD1
vib6uKzFC4wVUpi9P18Qdvy581gbbFrFMbirRc1+SWy3B8NPgmHclLSvTrLApWtb
vv4zViMR5V41EUa8/nKiJXPo3pf2wL+DUHNfUHS2bszVHlFd2YfOdtAVOIoWkUv9
XMmAMbWnMBksJ2IJj7Gx2gsIGWml3zPc0prbyP2d1HTg80ASJbn2YIiC4XujUEzW
GhyDc2nAuT/LqN8hQEbRut5u7iTXN1jE6ry6FTjOxHg=
`protect END_PROTECTED
