`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dhl+0KAb+jCbnah63cKW+uQGmtmVs4xsxtNMZYYkj2VUZKdHploKC17dOD77SccN
zeefPQemAmPzrz9s226RP5s/UpJD9EpI3rSi0VD4xgRxRNO/kipJUwagJAZR5CYm
uIpepaqvBpSb04ccoCJZDwQGrEBei0NGvLWfdEQmyhgw/EwFlOCrIZhdZshsDxN6
cwExD71sAWzOz9t3Zss0AbEObgNyr0uwGd3Jxy/Om7jJL1zNzXIpRaxqpGDi5j3j
KjQmbR0KHwDWfP3ywfHHp7DHDHBgK6J13P9Ay/MceNqLofz0FohSoA8u0y4mctfC
ZwkQJ50OMAq5dht4zyDg6aI1THK8RK4vdA8/4/GGNyMpKJVDVDVtqvr5Ofa4PQeH
`protect END_PROTECTED
