`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/UeNXoLzotvxHBtVs/RzOS5hhMRQSr0RZLdr8j0rm19AXxHmp1eLTA118GZrZEUX
Np0rVFDKRFwMU5RB8rgPvpkcOPDwLoLi6cAGjC1q/NWL3lvug9U+bLfzcf7IEOvu
1Zd4ZWtmTFSQ0sSikJbqY/mKt+6DHoGFf3XCYoja0Q9Tm8EUFs8O2RMubtlXW8Ld
cAG3fZbetnHr6EM0luvNtp76RVqq6Jy9+kw0/1lnbUrcJXQkFVqvTcOt/thctRpp
sudnAzixHjsyVD8Q/DGzCRnY7WvHzt+/jjjJ4O3cZQF1aJYwtqkr86QoLTHKhHO2
0gzxxbR4ZrnZu+QOluRMRj05pu8q8DxpQ0x2B9zrlHinicV3beXwaFgiEXOLL9Q1
K3B6Wc6MNYT/o6u91aH8K45sNfmSnSE9xGu/qUQ9ztRpkIerGOwvgIhUa8Ed/m5L
NWwE5J9agOzGLwpwEOdQs4isPSDM8PWVW2FHN85P7Wfdv72g3Hwa+zofKIa88J+Y
zIIyXAtJLoQ+qrM3Y4feKQTGVjWJ64Y0BdPfFpOA+/zSfG91GHR9MHLldbk8NwH6
JstEM5u55zB9/UGqjnBX6PzsDcKnUcCsVOrYhDFt3tK9fzk3JUU+E7UlftACIJ3g
Vr5i1FchN5N+YmR1ZlHYTmHoJ2kesHjvn0nji+6+CTXXygw9BXRBmWokb0FsZ7SR
PADi6QRqlrwcSa/Ee94VTD4D1gobm7xHcjtV9P7QT6TImwvXMjj9bwpt3EI+MK+Y
2uEZqCLy7HkMK7wG4rEfLqqpEqz8FnYJD7TlnENvWw0O8VJ86LRvi29tlCKv+Id9
oh/5AGa5ZUG8KeevhuGMZmsybtbFF0cZRiEOLwMc0Iv/1pRWvAIcwAKrcuq1+Cfb
/DWUP1NCxX1ayVdbSWNtD5vhYro1InW9WSU7S4jGyF1fJqN5S1CAIrGRb+2m81vZ
iEEOJ0B0QVdVOkjkDPACHVNDOkx6nMRw9/RWYwUhaqJKQ4e79d1wrQx6Co7oAj+a
D8jyQo+LHV0VIYfOCDaV0RJYbUROncwa1qu0+IGnx01aA82fsESgO4xZP0IWOlgW
VvjBBXQlQK0QrjQIYqVn67gud51M+Abojysf0XyqS3C6HSWQSU00FG3wbwB1QOiW
bn384m/5dgnUsIFLR5KBnFYK1vxdHq9zX0QKtf3wfZmUB8mzLb6QodMugMaapPKp
nGOveyq3ONQZkqWAMi8EdENI8yZ3rS58OoTFhcD4yWrZRTtSfhiPIr8uvXpeMEwN
Hr79gEb0vntnC/+HAEQdS/yn0yj6xoc1OxBIrakm81Omr2pKb3S1gZIr5i5WDO8+
UcNtZQwuX8GU6krJeK6l3Q==
`protect END_PROTECTED
