`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2dG0VFHgepJlaj9kyW5Dgpdzz88zsoUT6AYrh4P4wfxy85gLJkr72aDkplwXfdRB
kpKvKS7yo9f/NXCXRqke0nUsJKuMd8jd+cbIzNUOkpC2jB9RV8+NQw9Ogsd3oxEj
wre6HJFjd24/pfLCwJlIHXvHEuL4uQB07zSFCNNa3ZP3g8ALcpRHa5ZsWx+Y+H7G
yZlu8wEA31YLeuguYFj3D/S2UOTuQow4FDuT1mJYI8/PY9lrr/OZTnFHYufnjWyd
yliUvNnkJPwVljsC7N8+Srzs0jSSoZ4+ZtpSVvzQsL5gDxK3hzcg5EuOcOmVzuYY
IdnTZYGerat9rfOjOcA/zaeXhdJjdR9E1NaNwubjROyJjkZUXQPVMdpVdPbw1G1W
Kb7wvDIb0wI28Ogypc8J3/XX6sQr/xWu65/tIs/oENDv+L1OfW9ePUJHFfyDQySl
TjQ31YGAq+8X4+Wan+PeOoWVJrybDTSJj7r5+D9LH0ECKAxOoFOBwgL+iNP/D7eQ
rQwz46afwEUh+rzF8dSHtvjXTel1BTfqrg6M4aa1hghXiNF0M5P7/F/w5MWx43M+
FVp9mYwK5e2AKs6JF5Sf+Keg1W0JoMR5kJ1M6HVbmAui4VULY9wsvWyN+kn2vASJ
CvI9knl3orHkifIiOZdvqmEH394YuwinyhW4XFoqSj5ZsymvuyLwBhK3REzxgLE1
3ezY+8kG9LnTjYnkFMzNTL6OlauWFgLC4qgHFKP/MNDin+g593lbj9fi/xioNB5v
aQUfCd+sCUFCopcl64UQcPcjMDEx04HNB0D/yQJg5RhuAS7f7+9T9XqPM3C6C1ym
WvEFBD7ujevug9+bVCGAbT1DDmMO5B46kBdZTe92YoMVCgzydrtCzfhq822Chj46
1COl7z0DO0sEeoTIyX1RbJYq77eiUqBt3feTLXJ+5ngbBZuLyg6WzwVVY0ffwhUh
l23H3SbJDQ5YUvjgxYxIDQ==
`protect END_PROTECTED
