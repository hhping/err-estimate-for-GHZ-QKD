`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qOOxbKxMlD9iXiNvc1nSqKEIBb0P7auaZOZ2blzww5iHT89S4DlrzcofCQmy900v
H+ziK7nGWuLF/jUqGJspOO5oPCDUpXA6TB1MGcwULFr1/NxXOj9A+FThP3Sk5o6j
INOyG/H4z3Yd0xA68gdFzFPYxJ6WAWStx/9fuFKp7yS+FuFGdVjKHq2/ZBdkUDU0
Otw8e1+iGBm/k3YgXG94E9djhuVukiM+IZ+X0p+Qmo1ppXhqh/oYDl+ehMDLtSkJ
LQscAoD26xCmsc15lYQP7XPoe8EzPVcwVe10+o7bLjpm89Vw899Rfb8QnX9taxjT
IkxNcYVSzVRlt/mRIluXksT9Cj+FF2Dx327ZbF8NhAeBkljx8auYvPyLqTRO6Nft
5SJlIwniRUq57PMGlMovFfPEXgNLxpTwDB67lVKbTw5rAMLcqZupmnMrMnkgZlVV
g9ERBcPU0lNrB+f7d0eIOEKbaen+0adZDyxpZUAOd+zXLq0SfF5omeTQUgg45/LG
TttpIi2ENs95GkW5xZwBXlnoKcjg6/Q4ahL6dkEyN2zR1h8mh7SbzFksZqxPBZoi
1vCNl16geGO8DqguKCQhrIyivZoapucyYdXrvoKJb0ExUpD7yTyaQxQKEdAm3Vrf
L9Emwp0JTNIPTdnaAYybmLynE2JeAfEy8VJu4GSMNrVmSnbOWZ3hObV1p3irzxL8
8X8VUdCD/mjd7cEiJrVjJlFpnjiVSE2twt60gmM8K30IhMNEgy9T5mc8IBibG6Pz
/UOnK06bwXtFBhLYBdKh7zgqBF0ztFsvd9Lks+vw5YalAEC6K1lw2jdkMOiiRWZy
`protect END_PROTECTED
