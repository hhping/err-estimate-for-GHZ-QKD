`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PokKuRIylvNchFnqN/dCQxl/Qxb02u3UJW7wgKEOPGqgUZsyFFHxh6Z4CAtO5Bxx
mT5x4Q7ZcssrgxdLEY+cjkS926SsgB1WRh4YWAZC+0+KVZvUVGyEMSY9fMMA4zuk
PRGRCeMLl9ZaZjm5MeDWgGTN4tBCwpoyTcm35dvcJe4Xu2rLacXo+hauOaGfeY8m
vIrN6/So/o9Fqtt8dDORiDRrfO7J59ctJET7Paq8L4ZRBam19MPYdjOBrCn5Zm2l
jRyu3D/514vrErUHCfyjIkXaeDHA8M2aUGQ4DNgifjXhuXBdfn1LgWy4begQnr+g
rzMgA3s4qtP4xyARFJZIevNlSdlOkHMZ5xz3qaEP9Jo=
`protect END_PROTECTED
