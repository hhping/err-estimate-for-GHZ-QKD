`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EufOkIUIV+44O5p5wnMAqXwcBPomLmPj99HdzumQt68chvTFOHDwlfQGUvaJDaFY
IsebGYr3w0YbOo2QMTHnM1NLM/gHk8i/VfzUx9Rgq4DosTsWjFdjyyZON4/bAzPm
cu8uFkJ+8LHh0ILYQQqAv1NZwmiMvds+tT3TWhJaw4TXdtwyv88bTF/d/K1ekgxS
epXGVIQiO0Xk0ky8/W7rYOUQo34Y9emQSkP4gQ7543+Ev9wvLy8EI7szuFYoZ5oa
L+1AX15dyHOvEjK8s1Ba+khKbz8nNiMsY8Gvq2jRZxPTkWirb0eXiTMp9xbmgBWH
37ZUSTqbI6l3u9AZIVIx/ZVTeTYjV1NWX3HNPFQe77ZDWcrScU95zOjeJvzpxZ70
4f83cuu8ADOCqF3GkveCtpSpO+2mlln4XZ0E7u4ro0S0vmA9UIIx4QqDuQYcoI5N
QbFCma0vf50M2CUOma1HPYE7h7fRNXdHI3W3JyXxTtoFAVJTYfnRCFaHP9pbuMM8
1u9w07pjE4uABSeobifCf5JVVaVMwle662Sm1vaT7xq5TvVx6a3LGCZm2DOLT4Js
5aFsDpR7O7Midywa28kG3ETXdZASlXQ3h/VdOLEtODY=
`protect END_PROTECTED
