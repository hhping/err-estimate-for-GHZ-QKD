`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t21xlCJUYwrgdDA5kak4Kl/3vJGqYkP3p8pT3WkZXAgCNL6CVQqRUrhnRrVYeGtq
M8xuy1Sdi9grGRWX6sGABYtKPHQy3BPdAHLS0g4sUljXSIUaHMQzbU9iNCYwX3NQ
YJZLoc1uJgLGDNTN8Bp6KEJogEc6rs/x42R+GndTXB3wNobq14NqJQIQftcnlGy7
NHYNPfeNhYwBE9MQm+Nkv3HBp+JwGc+hVVEPLQVUgLi/62pCAweSqhdOjTzGOobx
6DrFQLkd+ts8sJ51PZexsDeigbVtzvS53ijZVsPzHtnD8lrkrH4KBGkzj3lC+RV7
htRqypPdHW9Ibu0QrawinDg9lGlAE7neHn3lo4O8HHrwttIYBgokDzQG5SMV6GCg
`protect END_PROTECTED
