`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xSy6WHhlQyyrEmaAw0kDtduG4vYFTqADcxMfgIBllnpeTuU28KTxGyaJRybjmOsJ
oXGWrVFYM/FtCu+22SPl0v5VqFdUJCWWrt1TLqfQ/POeRBElvWRjhHCHM10DM1Ym
uZaRjIFGw9sODRoDua/l8Zwet+b+cDC3zJxEXBuulucHhF4JCmWmNMtRTR6NoA19
UGT8uB9+TGZQlbOkcgThEnqlomW3Uiq6QNegX8B24uBNkuKBswzxQiLvFJCND9wQ
`protect END_PROTECTED
