`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
omex9rVTXTe+/pOIfUFmPjFawkla0C0sGsEWBgSA31xWBs7PmII+wVyK1w7cXOnQ
V9J6D7BKUmXWKAiYVUPzAkKxR1TZu44kd5sYF2Dfri9D8Zqxuwby3977+KCUQEjt
0DlyybF6Nx6a2BtuYcjpTVengL7y6bcQ2Sot+zT7WXci7P1gdqfxtbSTl3Ek0CnZ
mlHQ76om7MO3kn1cjfwb//qVCPOVM73aS+qjxyRZATLIA/juxys+ayHfzY4l8el5
GcE0ehDF82Fl+whmgcYzgNv4R+Nkda+ucV6lCUEALZvaQGlM8oUG/W4M16WdGQsF
Fj8Y17t784BV4LRHQaEhfN+QGPHU7bmOpAaYQCa6DcI/T80j9Cl2SDZnlypa/bs7
wk2SF/H6zF4u+umuXfLfOJzJS7OgMjYs03XoFxk28cp1QNDAPigmwgwi9w0zOjvU
m4ciFM70p7Da9jCYXJ4CmUgzNepZle60ltdwFprgVg7fehMiJzeeKZRFfGYPc4+9
bdAivZkOEWaugpK34hRofGpDQrqAb2ziN/VKrfh6vMvPuUEwc1s2BCa4diOw90ZH
mHqCsJBCu/sBhkVFtsJlmmfkVOk/IradgJ5V5x/1wZCu630B58+OMvt3eJgD4+jR
IOoOJVca9Uw41IGM+JzAQPrnBZnu8iAgZ3l7Pz7/UXEfIXzMcDawJ/k6mh8E87Hs
L1A2vw1NOcJhPVi2O40X3eMIPOuE8OsU3J9cIlRuAnwSoWF3ouoM6PN/oHgSzQ9W
nh/E85pY7z4Gve8/erbJURswgSZh2AE56bUvn6H0t6i+382Q1AP5/k4w2/cHL5Fd
YiPeaNCVcqAHWCgEMBVJ1yOaCXNoi84SzI5iYMviO4EZ3cSmNNJC9bLGi+6kG8wI
zbpp7KZs16DrD4r9l2zkUqp2mPEBUUY9XEtHxXsGYDzQMIuA3sB1SobOmX3PNg4Q
hDdlTk/bN8zqMp4hpHxu+Y9hRwvu2ZU0FOV5h/cIrLX5rOH2AtJFmZu+OBsh1Ahx
tqZwhJSZXy2n7M02lg5bIcPFb3w2CkJ3C5/ygIAi9VakNQcuONc4hRO0jLhMQY5k
Ii/0eWclWDWr1pSL9/km+J9e1cD1cDaob5QXKeSicZkkB0tEGinNEb/YnzLcdIxV
GnmLbV4h9axg6Q0R7Pehu+EpVwuViuqOJKWSWZYtzLU20N5B70WmcIqonCexq97Q
8jj2+lbinZKB2sxjOx+DZlmpCl9uqR2XOt89pxMq6J/K3ZNSxXODRLYFWAET9cjU
Y7pa0WOBk1WkyCTJl2PYWCuHwrwSA1lh5ZxeFdJFc7IsdLvIwKIkGkd6l4XT+nW+
HQKs+JZlyU/MmcmXjKwaFeOLsZvyCxMrkPLGDZY1YGHu8bbd5GdJOGZwGljeB93u
x2u2flDSJHDX1hj1yg3SW6tEZKaSTc5XNHc/p6R+2sBxIGHGggk1ODBwfwPXDYww
62lpzHr71Xl/GNY0n1TCWR7ajX7S+/KB5/zl+Ze6vdr50QaJ5e3vwWVQ3el3zGIn
sB1qfJSLxFWSxBnFu+BWEmEPdRJID/OJPvD6Kbn5mvLoUDLnu+xRjEXjBQlB8YoU
LQOpfL8mFpMQ+kDfubAn8m56ou/MZPSOQdFl7o8uAyYjy9QXsHoMrXN9H/9ylE4O
NzaOt9/g7NcLvWIg+HDPrgdBRZr6Oj+uVcOWcv7nCyaVlGPlxh5elcXYa+AR/Eug
WpME6RzruH0ReofoKgiZCU3RRIMgr4wW97hthgVzoL4lF1aAaj0UtHonmNmOeRuM
5+QsQuaX4BAjpwxdOSol9VEpbZDyFXvbvuGPEAfjqmJfJNT5lHDA0+pcNOKMzBnH
GWHN4CzhjjkJOJME8zm49co+jP899VKmy1bnWTSyD04JRcwgcdmxCDMyIOtW3E3Q
EsLceyZ8ZzB5g+JZf7RXjzZEOrLJbgvDR1lOV+FRnPtWqyXkHMol6OFy+LI9W79u
58MpPu6gkJI/Rc997C/94xaQfKUs8voBbLpCD/ZgaoddlOoKzRlwIcwjhMapz5gH
lb5eKQk9NkzxTf7GHtR8HIK+LPgeODtGyRR6y1ic9bu9NiTzFJ4e6HVnucDR2D2m
dmv8fNlmAfFm5Xtr3uOqm9he9n2unL8HX7NKJkRg3LgkYiq9rQQh8TzR1cdI67IL
h1MzderbO2wcJyrUrmgeYkCKX++ZdMDyd+i+jj6rvCZGvDzubuMZecIsJr1mNwAX
oYzabyBu0gvEeGKPuhnAyLFct0kUrhgWqiqoG65C/iAuiSf7Gpbtj6QyXiFvnYc1
CE7uyWBJCKTfQO5Mn1d6nE+GehZtDaV15YQ5414qQBQve1yVCF9nFxNPpUz5bWqi
kvEy2Wvna10yPX4VaDr5JMKYwf1cuBy9iu1KXwlWEy2i2ZAIOpGAgS65nae4Jt2M
g3lE7FpwUrvlreurqrBvnDqksfcc88rHJSRlnJ6yhhWPKu3n7DyFmE1B0talabUo
Zuh1z7xGlNXiHlfPSL0sZqa7Dc6EixZb2vTE2gfaXp6aeV7R7qXgOwKNnhrMNKlM
87/X8Yu2AEK5muqxVH7hUZki9xIjEAyLCN9uex33QQD4loSK+3c/4QWw7f9vJ0D8
qhXCFytQbtKaGgLCA7aJPuweO+AkTCXyHwe7kF97tf3ep7iNZhHkx2129ePniZeY
NEBFweKHi65NYsm/nS2q5sPYCNEP6YXnQyjlAIRVOlmNmCHyQUDrs07gjMjddlyh
ga2DC7zBsKBQ9W44i/yD0NrYz+tPIzo+N+FUXtyaTrYVUjyZrXKZdk1vxswr7CDD
vx+DktNq6eum5qXeq+v3mnCoZgQU11jTPER0koE2cIRSNTGCvQJX/4VClNaBUbzi
iXo3T/VSxVaWa7swXQYyNcE30qk7PKbo+ZwTFiv5d3PLnWThIEXULaJjEmaYuRO1
0ej293rPsDnS5opAQJK5ppzh31zWAuEQyWYeRXIQ6+23rCuQ8RMsV5o8U7BiZEIn
e+MZtMvEiWlMMB5IgyiO0uvpbcGkO91n36796ZQCWf0CtQAsfssoVK5U9vnzXTkA
758gTAcvDuoCLBbv17RVgncG2dt3m+dgyB9q2rAsBd0SJMVjoi4stt6tCV8aDidz
UITw2I5UCDzCfrcot6bzVokxOFzNAB5JSEYODmRpIk28cTvuuh4tk024zya0Qk2C
g+pdbB6gXaf+AQ16WBi+05yIBJYAnGf8RW5smZ6YFrd3tHLLPhAQ3VGyMTDDJDOs
5VTNtTXdkebK5nBkPDZBs7M/d4NYHVeukUivs3U2opq9BIpYsPTTVKkmSLpmc3nQ
RJoetIrj0wwxUpci1GqAou2mM4vjzXZVPGDIlSf3aLzXcZ0TMNmSGAkJTGJ2Z3m5
5eXfMYyc9sPyLYDCZmYTm1sZJTQRoknJviJG4ttTjn1f/Wn/wVAlp63lvhG8q95h
W9gKXVS+nPS+Tz/opvrmiMWmQlHcImNrPpgRq3DnHrcHVID4zyqXpOYAHwwju4oQ
VDdAyNZVObliIrYtnP7cxyX7RRDV1WqUQjwpY2vhRgnWuDfJI6XzNBAnqIN3jK60
xf1bbcriD+TW8UUFtVniwAU9Nb0HedHnxQtaCuONCH3upe6R96md/kYW1FNzIWm5
VSSCEtgX/l0WU2ErVSwP4EJGAliYBN0tQNnG8jN+KSPl3R/j7hZmBwhilfkiUNmB
YNKnqPksVCkqpsKMCb6O0RZ6K7L1OyNz4Jk3vbBwhKkdS3hQOzIoKf9ex2yUu/RH
fu0oB4PvxX5RacfsE/64ULisERnZRIrNYkeUHhDsAPzacVYzyMhsbjsvhZEcC5Wf
93CUzVou85ouKr7xq+i92oWTcTd3G2ByXNtAuN6SPqqtT2zERHnqH6DtV5sxw+gQ
QIBate9Jwq/UU9mtHYQv+VgfpsA3H44YVLwECxBpZ1VzDyctAQiuKD+siuws08mx
j27oEPgwMQgdD2lW8FmAsFfPg1QIcZztbSHk9JFL3tlEf4SQ6X9aX6FEc4YfNTfu
PWDAGQNPhs87vqv69sOrla6P7B7gi2+hzmBDi9OEE65nhFyWOPf8bEejBkoqNqlJ
p91iv5pR0noWNj2hoFCZk7tIYJYTyyCdnY+W7+Isdl16smM6GK7clpYq2oi7izHA
i9fuJ2fRreAkE9p6VaV3kGOMsq6bWnV4GR8inVplPraoJ5g/mSnDx3v3+CpSDyLI
800psHw657kZ0JGx8AbL4NotjHkf5SEzfuFi5RSWG/KkeEBymsKr3HqwQQ1NT5PA
xlf1MGH4U0N3iIa8/glXvlY2CKD2ir5rStILQaWfTj5CxdvNIt8v+jFiWXlYltBP
3tv7B/6pE3DOJj3ecuxAprHKAFbllW/i1wQ6ZAW8sB8Q1SN0rbThzyOzHJRD3mQW
fG3E0WjW/DYaBscHAxipoFaqdU0peFRzka9TgRuaKwo5Nwgg5IiSMqe28JWDtwsa
Gr45DsnOl8+1gMfvpOXlTraK0P/JThz6o7mef7UAIsnz0fSShRmLhBWZheaV30vy
XLuqvehBqmqmvGA6i1c0la0K1avXQ5K5K+f5RVMHCRuVRVnsLuPgkJ1fnsDsyla5
t7qGzospPsYVeIbtRktrnUNW6HbyHLlhPEysuY9lxvZynk/Rf5k0RUkQgkTijONi
peQdru3OrYLTsga4XeoCGyobuF1RYWoHozVv43FFwHEpCB+r6iaNVNQ+nrFxR7TM
WqT7KYLu3vL+QcmZAB5i4wNX8yHeJUfTsoYHJDlJ6+xcFPjtGGBQIEEolvvdLRNe
4aNsuyIhqBkWw++alN/u+HF+9hZcwJJWOUNl51XO/s+qRhFc+WgNTzpL1PKHQI9J
0SKROi/OzZWIDhoxgM2OSYYfrMyXSDiOq92dXHdpN14Uj6rsN/Xork68qhlAYGU4
oESAI6y0XlzI6MoXEYHOe7lPqy3tEawjmk6Wn8T9MXFFKqPn1eB8KJ4Of+TgKl73
+DN33JMws9zNoar4sCjLugHCFZyreMspOPCs0i6GPk6hsr+QRed7zWNzPnKebpfZ
PlQspKA8J78MFRvGqtDJwQ995q4m/HLCpiKKraWF3ey0ntlXU9EZ1do/Db673YiJ
O1fdKzwqjaAiOJCBpTjLRK4Mzlc++31ZzImdgu7JXz1zaaBifqKeeZWUC06JAIm6
OFrsNVFdltj4q2j1cJNXSiQ6FG9/JYPgOs2uDm4ja0Lw8bPh8u+WUk1qi+5dufZI
V/5vI3UbH2xevldGKXZQIZESMW5uZbd4r+WSOhSVhjXH0csrM+eY3jNXIjPOti1p
o6tZqijn5lf9APAW/AUWTzOLpN8Hh2jTVShXbe0t+EDxz53PNTfL4rzNTnfgP5Vb
`protect END_PROTECTED
