`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aq8m4F8sGpMvI6Zy+dmlKzdVY5r2XIZtmnDxIby1wVzKQDwTOb9xD3TFeYbVIwDA
iur9/oxc+PoGw+XoTExeVofgpvv9tn/NvTUfjMOFhEaWMp2L5CItBTObD+P75boS
X/uDpBDOCVdwy8dIPXLAGs/PuwPqj/r2Fk6UmzzqSjwiBJwTLyMcDlP2nYQPQZmN
VroIBRwvPcLsmPotauJsw7Lm8vPXDhaTa5Iz/LB2BfzzlKsnjxWQq98ixHzEu2kr
uhIUq1KoIYRZtFiYsndo5sP8wKhzkP4ckdkG6xz/FV0lHQydZkH89ylcRAqTXN1C
mAkonZ/fg73SvFgRXyBhgPZWHcrmTmQPBQ7jGYvzFsFkBU1QeXM0Vwfz16P5Gprk
xJ0hzBDIKyN3aMLV+RVzMEWOuQeCbWzKOfB2CoeFQX45gcsY+WshC+WE90fpRYQP
1LG8b3VZHy6SepCKAZM5qruKpu7RCPVYym/svCTvNXrlkPtcGOhQygUA+lXS8+2Y
y2oiFAUn7bTL6paJJNmN/FshkAmZcSrYf4HwwNp4tNNRHvmyU1N13ZxtLnouXlSN
VwfJOV5hsQC8xy+6+IVAAPbuGJxgP0lOzj773koKf6QwCJCzmsTHGDOdIBSsGZiv
`protect END_PROTECTED
