`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ij9ppKRDQif5l5J5pDvSK4KIUAg+oGWncu93S5SIEtu126jBCSCBHHyXD+jldzOQ
0ZQtoSpUY7LRhU1BVtf9C+YVqubke7dveeWKT61gih2S3URHHGj5/UI7NKQ7bw04
/L2zYMVPzmvaiho4VyxpHN4/1s3gi8NVYZJCNoOV3y4aTxLzPdMUERbAG4dIaEXb
WFziG+TSTwAAzLo2OXYPJ6D3GpGYqJgttSjVeKicHR6/5jhESm+8si2iXEa8jMSK
YMKHOURA7NasmpBa3f5mKFV/Ko1wPZ2+ZT7+hftkN5bBHhGjYDWczsTon5501178
ZsqkZ3DX3iQl1aT3DcfvVTmzKy8mIM15fWUt0AJEXj9rOdEurQGcTQaI8s5wkDMX
YGJuFxGVI/MrTigprTlNRTSC0NWGyHU5qdJJpnM+Tjvpmb4mpvkaJtXYt056wGG3
kcQIxWwarSA+iQSq+ADMA60ryK3g49HlPiZnJpXV3q29nmcbmShsQKGsG5wcp2Vs
vRcpjV/JzrqJn/FDysUaknYnXPW/q+cXtKhY2sGRXVAIbeT1UWlVLgDDMJyej/Ua
6f8RppDMAMIjNpHq2TjRgVl2e+2mTCzxutYdQ2BZxjaNg64ilJ7/0K83rnRLSd4D
LJ+NRCVBgRjGK/VtPQ/HOpuJAne8x8ompdwEV2kVemP1TLRHaePUw5aFQVWMB6el
H3N+qS3wUmSYaQBs9Td5AeplNFoG8q7SqFHsuCT92/kZYbAEXs/hMCsffdO/67FS
U1eTLpSgMSbvIUYzvEJYNsU2IusH7/JU1dmKYILU4sF5FAah2Tc88bm5CrPSR/yb
4JS9Mikq7RVLT9jaWy7uILbOVv95HeL9xJ1rwg+XECPrb0hZqsKkb/AAngZO/8nh
V1DPDnBr3pmfEhMCbHZ3c7Qfnp1rZQ1He44HRSKBrvJ6Nk1K/rlIFX0DcheM4ue7
Hnig/L3p6rqgcdquT3o85VzC0HaZv2wAnKrXKeA6d27wK6V4G0z5ohVUJQjOgksk
CxLCS81VxfUayvFAgQca9yHQA8aJIgKYwrFch3QLPS8=
`protect END_PROTECTED
