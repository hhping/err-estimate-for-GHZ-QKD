`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EX0AGNduaA5IRVd3tTt+VQ09NW+Orbp4m7deUK0xw//a/5yxC8dWwg6ytHLumjAR
U/T1ppsennylPiuJFwEkLicFf/72YzYSVnRVAHtZDWLu+v+UCa6jszdbhWgto8dO
qD5+MPVz6QhAojYsqRT5TxwVnAsxy4tj1++/XnaXiR6heYppTgUAQlZS1I3y1wM/
TaRTOhwfGkFdygbPQ09+TW12ivOh6TK0ISrrxP42wZ6EzOlktzY9igPa59ZlKqhV
vr47Jeg5tTjcBD+6rZrLdIMJvaVl4s0MfejspGcaDpR5+r+FhJC5VCHBIbMC7mjB
97EnuFMPK8qGow1/UWvQb3axX5kriGGD//OxRaeANqypmCy/3zjmPA1pOBxf8Zj4
wA35WDb+x+wfRIRUzjOX5eNdBVqZuK/ygsGQ3OWeiIUzYKUb4pShPQuxF86cjGsD
xEjg8ddRaYRANOMf/OAJqmT9SjNoTSVifkhpzacbdK3dnDC5Tp/3qep4UIRLMSil
RBJTAz7xWKt58Cvkxkxl6sjLukgA7ZRKU5unltBC1VxZ+CNT3uObYIrlv1xSNLx4
0e/TEAxi77/hO6vRQeK+H7NnXMHoglarDwX7R3y4pmvu1NyUD6cMdThESdOJHLeo
43MPXb6TtaAW2VwqmRUc5eDKAOz4AcmlXfl9UJKxAKNgOveQ8g9z9nO+9Jjm12X7
+QzMAhDRskw0WtYnrHdL3XOI1sDqD6Qk55eEoZDPC+2hbptaZdytd8TTrnC0asvc
rxnHJYqhsHKpBEg3zju5DnDCLS5OWz2DlbgjVy4rmk8A270Ikf+LApz76SVRdZOn
wpe7XGtXMsVV3czXbVJ464FmzlfnJ/rgIEszUjKkjyIelopntn9f/ZdGkMfIKRBn
u4zXlmRgz8RjZYh1VNYR4a13ZjogKIFVgRhnkHSVicml3O5p5clcGiM3oEamHLb1
T2tnr8WqJGXsvcDZUlKMFA==
`protect END_PROTECTED
