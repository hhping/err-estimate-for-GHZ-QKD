`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
peTsohmWR+tsKEulYRjPEkVy7GgPt/Mp7p6GQDrcGJUi68Ki17kCQg0AVfK2THVQ
BA9rH89Ly0mkmhDBeMux2BoV6/3Tx0U/6xrd3akjs3Mgvwwf+DNQTFl4yWxUOXWS
dC9sf1bhai0PFur/iSGm+PByMHfuhO6RDR91zmkL5tixn2+GHdWpjRNFMb6Q61Q9
TEMeNs19Y5J0A0vO18nPhSQmH2hXDY8AouRFYEt1Oog3mzPQXefervjPNfeCAcHH
SkiXWyOCubeyEG0Xyiu0cbDoUEhl6IBA+6T6+Tyeu+CzXNG2pZZVmnUapq5gvXoq
NU9uXp6Eanlv6mOoYSMg4THSj7CCgEXi3wZK5b3nAjmPBVrqe+9Rd2+P2SOABBHa
iURHAGhfbcsqVL/94H3efwnQHa0EYYjgfh/j2RpJD/9VXbRq5Gxm7XlS3Kudit4h
Kp0yqb7ixt2joUgKmZTZx6aeUF33WPNofANgI2rFOaKptF7ek3iNhnDx4jYF97OQ
96cmiDfa0ekVwcYHw6UZDhjBg/jIzqEPMFkTtG84OSkHW7aqZqD6INSBIKqvIJAR
ZXzY6FKMk59yDCDpiiyjQyPvrA7BpBW0r7cpsQkhChbKx3YwNcNiqD8Mj9eE3EIR
dFxWq2nQITdKNhTjGb7lVHJ8WWevYlKb2zGfL/8HCyvYibgUpTn+xKVfOrgli7hF
hqphkWHmJfYoUuoxHSIN6fk70eoqABPBT8mSF/5v2OYK/PuH6l904q1YNpDnh9A/
AFIufFvxtsHGd39alSnW2/zkAXO8lAdL7q9/RMjV/ztJpfMWhqkk8ddJzB6Qrrxf
1srJbyBKU6buc52wk885a6N82s1Dh487CbLg22a3W0NmA08Mc7lV9E68lQCSi/BX
iqWtzoleLYtq6vAaLNMMfR4lbVqIDIs25mrmLwn4/Erxgn62viPmNh/r0rCoRkl+
aGiyF96U9FGYU0lSjH+udVz0GZjPM1y8voechc7gMEjdgBY88/TaeA80ulPi1Ipf
3mgpcZVzi0kzNnGZp13rKKwsXVjiKoPeNHm02kp5aasKzkP04AZXgUa6Jql3rxJM
6tGFF1o3ACCz/ykT+9INQrJfRzqjsIyeJg5LchH7v7wP9JeH2LwD1xKD8oj0zp+y
pBgcJnCOgRuaKGFE12o9MFHbqRHcKTRnCL28rc+rPbAW6FD69IXB81KvXWli+fEc
4++6FBual+dlDFaUMNUkVVLEOCaHeLDBUDmBouwVQKS//5Ejjn+2/f0QrueAA7Be
0l6er/q1+aBvu6Xfl8fWRJbernnJ1rCBhc35mqjLZoHCchN59yePf7bofUzMOw0K
bM6r90jc94bBsdqiePutdugdL736aMHJRO0Np+Wzn/wYFkSuCSrk+HuChg4348ZQ
EG+cxEs2VtArbU04ewA9Ms03YCTaeX25ezoCYp3yyByV469syoPXcNEiGDf4l6mv
k/sbU590hSeeY2bvphzCJCZgCcRNSfGSJI19yF2PbDx34esUd9blTw5zBTBkFNCW
/v9AbnmG3iIYrjQg2QPo52DSB2tfoHA/tVluO3lbu4LvqZG2ONg8989feaTXplZZ
+5s0uIZKz9JSkxoTnnsQYUoSK2gm9azJDZHxdTcC1oqLEgGbxBZ23BxzaQP+rGEN
Ytb6ROObR94hGLYXyFK3xti00nB0ZlNlwR+m4aC8y/LU9a7BfZYvyKYN0QDKbtsT
QbzM3vz6AbGyk6uGCTiVOxZXpR8Yw+do4D9op4qfc0xrQ8eMgkiZEexsupjj8jaU
4RPz0yDYE5XBIuGwRbhDyTPpwEirEaPrDGMUAlETHxtkui4rm6OAnkUJE02Aslhd
0qJakbxQ8V6HPsvFLkFfCL9Oz+JYJhxSmlvci6P3FgfdyvcqboObPmyj6U5J6cu6
m6CH33pv1DWAlayEUm0TlQvtxrZmKFe9Df90pPT0kvce+0KBxi5LqsNS97wRcRml
9K8ay031PvaH44vd01WFvNr8WkMx7uxuFZCSKigw+AlEsT2WW3qEpr98uqnfidxn
xRgd1Cj0quDcq8ZBk9qbdn2+KtwUPudOedTkelSzetpyFOuATYInQyiAJItvMUUe
NgtEOD3pM+prgy6392VstzhbCUx7xg9IqG3UPcfK0ihDB+M9sh1sRgjCmoA6pSHc
w4VulMRO7IXECVkKspXrKAUBvAMjODP+XWORcV4yoYPYRYp+qtX+IKWJ/rv3opdm
k2fx9T7baorQ0ColOjfvHXczlQO8XbGJKjdULyGtXZjXnq4dFdiFoIO3SjAa2wth
iOFBkEMc4RkeA4RlNlXYKSb8s0RnWuhHZEslk/uJaXpfovdOnAs7j5HDSWPFhhrk
Rrc4+kgnXkhQaIOK6bOI8KWVw4P1zWF2+bsA9A1V1EAXe8zdizxahaN/4yyhPDZu
/NTM/Z2KGtPR3ZvkmlRQpIkiSK5uVcftVBR0IdjpvCny1DZTmJx9pQux8h70VzTG
o+aM38FphujkjGYcf6+5cPyux78jlGU3ntzPfU2IU99VgxlM4PqPudt4nPqfHTjF
+srr+zTKpmQpoSC4TeGnr99Vwx8+i42Sg8nI1EBFhG93jfefFgHiEROj3NMjKQRs
9s7VgQAcmqseZasZAtkIi85syP+7isL1H8fwxYWa3Le9KuLesLCRxHmYI/xXsjpA
DGOMPI44YDdLv7vVC5Y4WnbLmE1oqXiEBIeEue8+4eqqjLak4eSoT0HSJ3Yu4ghs
I7KGV+ElNm7b4o17YqFAlSz7m6Qq9zkk1G9XMhBz7XUiFbBCJX/TD67GIs1eKxWk
jzVcHmkNadYi1hwcR872wfsoWY8uXyBic+bFor+HFkxE+tAdwpM/orl1walaaIbg
9BQZNfnA29A7CYCzDEUwYSeiyFmSDtPgrLS3XobiKBGU7S47ufuccvmEVL/sEE91
l6HOc8Ech08TMDFWwMU4+TSock0jSmDPElby5BWvqYus/QZr33Y3F+KnrUNYsXv4
rjiA7ar0HP9IHEn4t0s+mC5Sj2ifN/QLMQBJmk1MvU++dhWZzZA+6KO+/IoK/pjj
zSIOL3EzSo1LCZHZm3Scmz0aaPnHBEK/Uqh0Elzrixg9rIiU9WbKgfn0FOb8oz8u
6MHYyMQgRLGgO/vpuZpTcAPH0xJdE374zR11wWEcd83s36EW3/BtUrX7hzqerAUT
o1ohDIOh6Plc1RhPZohnd++5lPCQFAnS4Mx9Te0TN5txo/hgv6VgoyGUQAyIHUh+
Vn+EJrLDJAb0oR2DFxRbynV/PmBMbI56TCuMdimYf64ej3omOsqXKRVzaM9Fvs6a
ux4DPHJPmK6TsRujdPDzvznlXzOFBBJ4WuSA5UxphCHm2uIbwg9u62ugsPH53MlV
2LKvPt96lxoqVkB3fKLwJt9vTDSdj2tWHlc88rsxUqX6a+d9BRQ5SbhrE6Zg8+JI
eNrtmIupnW7CpBPig8GLMzK8gCb9XmBLS+DYb5FQPJfsweZyWeSCQ50Umm01gts4
ae1ynSilZlGlP8FH1wp1lzcfkqqKHp22p/c6wmZ1GG9HDQWRxhOR/HUMJBeXLKJb
4n7ra1vYmmL3/c3g/Q5/ovr/2rO8SN4bMFDgs7Aavc3FkO9yYF5/CZS5HBMxzMnS
X6uVJuZwA1rai9QoW7PzndE5ZC00NUiBT4zQvWNJy/I4E7Ncq2BRciur7+AOGD3V
k6m/kAhhc77ydzJoYnLs32YFmEw2k0I2fwOPifkdMl/QwaZbQsfrKyO7Zi8A3WBm
XNP9GqEFhoXcpMIO3xY3mexTBbG+4P5XoNR82nNROcE1SLhsRtGDwLs5rVrj1t6q
9H2wmOH48+kiy8ZQUM0hUBN50cUuQVJT+cF5LVFUthjjpv9L4LXuF0AzEf0RrneQ
HCIP0nT6WmlcVsNGsoUwokWHfZgkUj8UoodiYBzbXsdtll7NWZwUhk1UVcWNeR3Q
Dl+mj/wGdySE9rOvQHp/hG+8v744X7TfVJ92NFxOCvRAng9nBm7UeDhRC6oMzPaH
CK9it83po95mLNpBjMgqzpZXURHmM4PwHFdOlAo+/8PVlOeu3GnZA2I5vSXCuLdH
FtI9SZ7o9OjQHGCOAQKD4OhFn8LRZJ4MT2BJUOhVMve5xEK/E8Gnsmz9Qf+bNGUm
QvVUC0GcW3if716Ojmzs7jsEPQByEDhbgufgR/lEdpCCUbVPnowlUcfW0kgPjnEA
x8ZAlEMDP6VmF6RpTF4O3cbYpoa4h5J6PuHWysTsgAGRMqBNiR+U9jvpt0XIOiBS
K7kxymn/9P/DvoQyz5QSKNtjuH6bJ3rlrfjIznxM96vNveAknDM+TpjWJsBg1oZ7
kL9/kCK8FMbORsGQyMC2vOM7zleTy8csFZy4dWAIQcWZGNIgTjZ6uqP7PR5Nceqh
FHNU4P3z2wnKGt0XLCsDY9aEJKFjUrI8YxqDLcizzB2o/RsnLOilLqFLRjSC/LaU
Q/9vRMlT1sVU/BlUa6QpX++IG/hrzWjQs9tLO5jMF+TQ3lP6Own24JpGXCtfb+tR
UPXfvaGMhwG4wjn1FnyqjvpKOitcn5oKUHABi7qCKIFfenD275qtdmLhhIQOC6Tb
4aZH+JRKIIHJft/9LiCAeIHQeZDfP2CMEzE/AoZ41m45jml7oeLcPADkryaCYKvu
pvGxGgsoxQOit4VKGgv8qLY36m7RPysz03MSCa0canz3KwSq7NEbUOQYRliNaTio
NhpSro+4+gONvYsSLYs6L44GqA7TRyXfG8+C7shOXHDfMSwaL8YVN+01hEdpPQrF
eJ6BV/Ey1qpZw2PTq4U6vEueCpkWXq/8YyygWZVzD0M96JUNj6cZFHl6Y/9MB/zw
5dZ3E+TvI6qx1EDB0IHRoDp9mzv6Zk99kaZMZS4AJQ6G/kgsgLErMXxHOym5DTTJ
hp5OXqjFrMtmXHQ2Cw11LGpbiOFl9kY/9LL68MtQS/df2ZjrVXoZhpTJYJXQsUmI
9GbTxHvG3BhsmqlDRSG8KHfaXGBYA+ZQMkrj+f0TohCZmsXuJ0LCX0X+XOZIbrvz
ZUB5KWuY21rSDy7ICIo6unfCenoTf++EUvaIvYhWJMQP//pIVNqOxp7ckpn1t7f4
72roTSxB2umSInXp/iXUmZq4Txp0pn2fHkaHLREMJ3KI08qryjBrXtuYf1IA1aFw
gO2dqZcpQ4XGR0Oxgo29v3HZZaFFbNIb3aSnK3a3kAWkB1ZcRt8ea+Se2xbtorDH
my6Jhhk6A/ZXCPicxK8eFDfI/ogbH9hhr+rV966ahHrKl6p4PU//BKHRQQrpH3zF
bd4af7wVBsDESaSAO6bYpoTk94CaRM1/v8th8n2khPWYvTmREl57LcxMGRfOYcq4
kt9xpy7RN5GSEdpOhwk4LxMWADH/VpFNxY2yUqzulGLNY5RXRQhohqeZAfzlF0p8
77org1rM3ga58QkY4PhO6MP5TTq8WB9tFeUZ2LIEWJnhliM6bu66MtOUgPmiTWMB
DMdMR8zopgJs+R+Z4wxU9emB2VroaI0+Hf3zLLAzPIOfE+yDcdW3riGIjEbuF4Dj
K6/0efE8IFKCGY/L5uY06wU/Px7I/pGjEm91OIezr4uSmUqNOeN7JYJwF5CrZxrv
EccLbDtX6/nz4KmsxQqwSQtyJbsdI3qtsXgxAyDiM2lKpaOoxpwHmEpQ0SSBy0Uu
88dFlRxbDWwHFPkliZ7QISyXh8EXHyUCHlEBKBHiG0//YcpgSlvefTXLoYzw8rH2
0odcu4896Fo5KZXRXlDuarx1EyQwGlofzmuH3CoaVrRPyjusmHk9c5POXr7dVsns
dYYRpNpDDWuKG6FgLa88LyHHCccYt/j6fjy0RJDsRNUHrI74ezdA2wSHfrIjPXyO
FlT3Wno+y4SbO5b1pxF8JVKuwmHzSIGQxHjScV+3NxuH1eY6Cw5C6FXTUBi9yEPq
GxYOX83mhtvKQeyv9NwCAPVmu3Ha4onyqwfVPiomC2Vi9b7/fd2JNaPixFOU+MYX
DE0b/x+dhgX2VfDEe2A1ky3Bpu+lqqQqMgGYb0FtA6k1qEln7Kr86LZnCs1epfXx
a0N52MKq1jffJHxd73/kkzo+wMo+LArFf44twjb1IVfxpfJ3bAE0d90nP/DnhE6u
Qr1ckjGMduOzZdkpYPB/E5O1CCH2osbWdtbJYxFHPynlIvRXszyK+78dLEb6d2w0
JxpdgC2SBXviyJyxoaE9CYc21UgXryRWt66P/W01MyDSIKzkZXFhWBZOFp9AHUDP
XhYNABMf0ujDBSNI2ppw6lABkvIJ+g/gHaxuRYGnfLRNHnReo14onynzuLaEPraF
djbRMDDm7f2oC4i1QUfM/5lQqUrQzXXUfx6qTMxSfuSY5mjrGbuUajo70YorvnKv
LZovpRJhu00BkLeXNioCn7KUjfm/lHJj2SvAqjzbBn5ObBV5xd4gVif0x3d9J+Cg
6zBYQWnr6AoKYlH0SMQiPQNDOIRQ1y7TEk81ACXaxfEvd13uHfzBaerdqG5YsZeq
BKXEO4ZwiE4b7Duk/grSb8K0fvKPldHl5dAYvkQte4864BQY8shy38t0gDlf3Vps
h+/6EBO/gIhgq/DdKnB2+TpwbGQYAR7l95kv4JYCZYhsc6wzMLsBnHlRLk2LChCa
cRd/gGnkZOKemVTWUjNELlzdW383ml4nGP3M6KIP1LFpK/3i7Mbb0HvTIX265d0y
1ved5OgKhBDbUwv+H+jkPOa635CYqzPVRc6jkU+QZdbQ0pSMchTVJYYPqqlsucsW
wF0t3+wxe71b7rxE/jS8V+k1JmOqEUJVq+1Tg/FqSCd3WxRs7IYs5dLctC1Zc1d9
3PydOAWxxrE96aTvgsIVUKJxodgI8FtVAcvnR2+re/iZsaewClJ6u8nCSNqgL1eW
LBN/iJeuhiZ6oqvtooSmH023iks3mxCSh5z4pmyrZesuxNH483rCfaUK0iEnfU9g
hZGVud13Zl6PYyZcssIxmE4nCF7LrwJfqo7RobReVAJUV1RdXPaHgisgd1fzrUe5
KfB46Bv1LbRV6YAgKsSEchp3sCYSTrkBnXGJmB+mynAZalfkrY3VP22VTsjb+Ylu
GZUXyaazyJLT6UVxri78h68RZdBc18TkS9dntCyveKpOKdOziGjyflGwmmoyRqil
kLXWfdTN3aN1ZeDVERlIwkAHVmfCXilMTEoEaCIwaw9YlcxZLo6TQkPxvg+YyGBf
oNRl29Prb0eaweKJmft9RgVvl770peMjSraMIGyUTmOcHC6s3/zdIGn+NZsrHx8f
w7wp7aECQT/JHUPvV/PVdJ9YeM1jLOCaEoccGUA0GrlfCEXaC2v3ZSqUYQmSbDhw
VL9+VAoyoU/QyjA3mXBYqba2D46IdGxWCIJVS2HRdD8zSsz1yTGy8294vRpLPhJY
I5mIZtLV7cVr8m0HxMmutOvSX5Ogc/iUTKLiT4DeCZJpiaxLPR7F8r90xef8SHQx
VRDyy+l7H9zIK+vFS6a2f2P5I6SmLN1EblEeHP2uEAseRaFtza7kXAoFkxWp3Mxn
rbGYXxNcBxeGDZhaRMd6M3AGA6HhEvGM1LgnAifu2vcKRjalEAHd5ErDhbblxz0c
/hDCKiIuiw9krN1mkLoWS6ptCE1Oq8wYzJC4jKwp1jsh24quJf8jF8HfHjKEujka
nB2YioDDrkeGEynGtxOY2+U9t+gVhK7oSfjZxggJDYoPKwYmKfZkXXrE/TvrS5HV
ndK9Owdxl756AWYYFjHBVhE9Ol649DLNnwZBBNvIj8+q28WUkeq5r+NlotIO41u9
gUuf1cY7FUNaYBFL6gDKCpQeD3i08OJwgeaAFkkcushHKQ+byJ7zwsPBSmEFpY6M
3vIuZPaaibIcVx6CvchzSGOuy1+VE9Hna3lzq4VvVLk64kwdarFFXdYR82ZENO4B
zzW5NNnFg+33XeGFpQme5XYxOJBXFeMknxpV0VFOO17TYQ76bnkT+3kL9uIF2oVG
ukWTTl3scs240bDlaAIcUhE0n5oYj1E12AO0UvXByxJb+tD2vvU/J0qyZpn1ZQPX
1O4ovCWQ3+9UKOuF7nxiZQictj7VpZcOp75YXPw4rczWOlHEGyxp+dzQWaylGjZO
Mg5VLyQ11o6YMHSNsYdf2z5pH0dVIjZYKzY42HFVzIcHO1HhmPtqRBbzX0t3dK2+
zOFV4LvYVjOidwZj8tNceXpbLMl6EMAXhG/GXSFxDKeMz9DKWychaNHil/6LGdhB
iLgJ7Iaj/uRS+6WYfbaUYntf53xgj4QfRdDnGs1EM7atHv1He4LCDgFRK9R6DxEY
lTiCRipYLJU3owIc0KYGGgyv9/5Fms+vEoudvH9kYDDvJ8pznFIOKuQY8RmUXXUq
laElqJnmRlle8xD1m6jPw65BEACMHqaOCmWmdTV7a5E3Q3pfbbZG1Y9vaqWWTZMJ
yfwtPoXg8P/DgFvP2ELFq+jERH3CsBv+WjLiLmF46l2sutAVrJWuKa5QjqVwn7at
IsULJjCsY9L6DWeSNpoDfG7VBWZEKakONPrTXVyi3vACGa7oTsXfVHODaJz8j03u
DpPxVZdiXtm36GDPR3Ar6kwk8gebUUVR7OJuYrfdvmwcRtlSGzpmetvuOeSVl/8p
/y5XgyMk3gK64bwVPEyvoFwOSokWtjH+xc3XWWnV4cYm0renOMOPIdSQkuBJCA8N
hItftHRr3SsYHkaolIQNhCOlv9JXnpRHhWyL4WGz7kLJlQf951/Q6FxZsmTBId0q
lErtA5wfnRabWI9N3cVWnNFvDEk/HAepI0eI59N57lnoY1cqrSQDdpjl5LYKpz7v
0+6xsFuEaMIgcayizz81VtF48Fx84sWqZUrlslIMtPeQG/SdFB5/2sQICP+ThYui
RI1Jhh5U5lSGNWjcfyAp2bHfgOnvSh+XFbczZFctEIkNqp64/h/qsOzsbgceQVQ7
L/j7jI25YCvagGxaAa7hjfkv+MhgjnO1ITdv5GmaI2EgyG9tO2Fox3dmYVQ7dF2n
UZJn6eySPoJ1G921fc2wfh2ZWB1/AlcxG5AehbY/tPbL1SNN9unC/nVo8k93GFc4
x257bkxqHYYxDlMIRhxKhxJtNahUGITbhaDNA/CbNl7g7+fXJdIldOVhonesD66P
kBBhioyCeKQJ8xJjEZrsC2vKXZJj3ZSzRxZFxIrM64r4DHbRTxea4wDvsvjF9vDN
fwXinbOd8OJ9Rsr8jLpRFGyketcT2HoDXUL1X2CXQVqz3GlWR4p0z9z8+KcfP+q8
rLcxJ9HqiFcOq84ZYPz/jqY9DqDa22J/1s/X1vji4jZ0x5KzStpbRDQ2+vJoUsiv
qjBJLj1BpBmfhpRmz/jYYSYr99E8/BW5tJqPfIUnSSeB+OmDEm7b0XQCXanr0Nua
FKkRYpJrjhloA+apETyx92jzhFJ8DnsFWgt33uIJgEdKmzMCg846K0fe6XnRmSnJ
uTnuH5Z+7UxUd2yAYfOZwAHjMqV4Xem6H5kCURlq6utDcsvopTFDPeCwG1YkMHbD
yt9yKev83L5Xbo13/bq6M/bhV1DJE8BnPsZ2orpO/YvnpYutS8sLV3/Xobjozw7+
3XnUQJM6bM/fIl5kIN43SG5UxWZARitwlMY8CSUYF6NmxZxW6mQxoRuvHrgx5xIk
NesK3TK8YuWrq3d2yUefMIrxSflsk/QduA9zqZnokJYhHMKFvGEZXqEbhiRBEjB2
P1ohtjMLMyMRcTXlPETb4q2nc11wRbvwC3wBqOPfBMN6otX5uhb8p2Na31lxaGsl
GaGvCqBMNElR/9MSayBACRbhLR98PtrM6VsCjoWCA8W4KqeuI9Pgf3l6tz4gJm8J
8kM97tbD1oz/P32kCs6KKJKxWz43uz61NBNrCJ3irPyFKBKcKc/B0tdEVUOeEW0k
dMhXduRPx3UiunKoUEDIPTTlzA18Q1cPEzJSWbgdnlbA8mOMUIRRJXH/1q5A21vU
jbReVVvxYchh1T3tq7Hci/x20xoS6FmEwOh+U3kCDeUbanE6+7rjYNbrsJoQQTFC
M/AuinzzxqMyEKqVWr4N7xMhZiYKQFPlKgpozOIjsBdVD089KrIpu+fMTORgAFR5
MM0Ni8wnc0QeJMc9zTDA+uczQBFERR9XcM8oS4XUlBUrMFQo9UmBQoNeB41piWBK
Mzf09ozxcdN45nofoyL30xmLOLsYAJnl+uvWsl4VA9PHOKHeyxgsJbKXVw0VgGjH
vyYwZKVWBDn60lLXdKyrfzZ6+sLNWYdXjf3ztkXzTB4YszwNtL3Oe+tZUU7d5Nku
3PuVs/9MhEFlJM6ebq0We9fH/HvsC/zh+bLKNtWmr+9YUHZDCJwO39wYx3GLab8s
JNqzjJKl3hUMMnx8Wu82+LxV/50WCXZTYWzpV+DJF/0QBYfQvkgdTZCemyfCoXcE
xi1dn1xa3+D6I4JmJyxN554e+KHAma94MNlWRMm/yUw685w7fpvJExevfkCZ+u4+
ctGURKZi7Rin70jGnoT2hB84ug9lO5xjQohhskLPFmQSyhvHPlPplKZzoIayyo+6
pDdw4eVDDROgSSAnkaG8hL78YFFj6JMqKZeUS4SoGicNbH7mZssvujT7XDpIhO+E
vmFko4J/NTh2FaPDpFvQsmoIdn/Yem+UAUQVFsxoeJ718gHRiW2MF+geMBA5JmYL
Aca8rQebF4ErWIiuA0zmcp9HLhjzdLvRnaQm/APjYHBii2G93836kDGcCJMvFM+v
3YdePkdEB8gy56dFzWKKVWDgtn6BxY5UwNY8tfbohLAWINd6lwrPV9LPd96TnycS
wUQGIfX72x133+zOvI42FlJfNSrDzscpIS8H7NWKYUKg71ezMOHpjyImiRF6meQe
zfp99P/sld0Z7MY8uVHdBTmj0jtUWZh9SVnBowDGQBoVhUCD9GWKuoNHUCHwErMm
kpl5skyrvKxP0OjAwEENFiVqdlRW6svkd3+451nP2QsncI2qE4Hbj0LXoI/Ob5NV
FaTyYLHYJUYwkYdjH1QvE1wue8GsODCVPIXWeHKiOl1b9d0yxqbinOjXm3xMZvvQ
XTUwOUMqwEuv8UoyyEWz9wRP/f/LRzDl30a+akjUUeTQs690uNdN+V0GrbNxAqLM
M/X7fvlHUzxhfURVl5UFUp+WNgrcTdEJuZ5I/h7f+zaDMsBXwMvGPVd9d7DsHCXj
e/PlCuli1FiD4b3OvfilAj3SqcJIZPpujdjGvx8NRFj/T9AnhtZL43pqYA7tWsSW
vybKTPVNNYA85VvecGlCCLOC4sN+FQzUs/+QNMxbZ6U8sRJFWVlQY2X1/HapyU+g
b15U4i3o6wkHYI57lbJyeoV9jkJEaBJuafy50JWMAEO2RZFfD4nrX1qqoPVeXyeu
gWxMeCkfhji6jJ9G+cBzr/fB4I/i6vIlZe9zUhjeK8kAUkOMjqCFV9N/ia8JNJqz
9vdg8TzF+zsGMmxjkFlqjp6e5GL3kDYINIuDCrSOAPS8g7sWgQR3nUFzp9ju/8Fv
Y+XTphT/ZzUxiWc4wbw3t7xvqxIveERn4fFgKgUajLA5Ts0V7cBn9ZrK2rOY9MgH
nYg4ybvWdt1zYB2YenGe2/kLsQ7LVESeXWb2GjwN/6zKp0HHbcNp7Ij3+1xmKsCK
GvJA0MT2M4NK8JaqPMoQp3lrRlsNVitso8I9aG6IT+kyIrJot/y2DZJjt1QBG03i
O2x1Lr42RgSriOUKXDdVFeQFzrlRqJHnCPx732aHATnS3P7zA8P7wQePKve8nibM
zoHNChrLYoKFIRhLG7KpCp8OzSdPKJ/15wqtymbR0VfhGfDw8bjfx/yK0d8FkaQb
qrWzJx+eT51422x5J0xN5iz/qp6EnxeBQ0R2XVxy+YauPsA084wyBEeBEVCGB0Zs
ve4pUIftTtObyYE9/PSK0QgcNB9pPnuIu7GdxUQKY/QvV8WCyHydWDYINr9txtCt
G2C0WON5wQQ8WhR676yQUUAfs0NdczB4LGkXUmnYaUF5Ji3N4uSYoKNRg54RMxQA
vzL5MrG2jyBxPN1O/1+GC4VfGVm+/wyatStkqQnhbpuvCJSZt1LULDa8Q2YLJ/tF
hWl1OndGmfiriPoZMDYY5ppdyAfDcTA2PtsKdbygUydjzzFA1WZkeclbw/VdTPK1
vflJALVpKuPe9bIxCcN+8retwgpSOCNpbAvjv70lZ9H46Lt85ExzkXT/03ZgXbT5
6haHUSPa97WU416LDmcN4qEXeQtWVON4HXpzm5WIuZ7gZ76H3vzB6OPOXIc6gVmk
gecq5QH2RTSTUJm/8s5w3I+B0rrU3Y2koD75MuOjU7O1Z5tc56hsgcT/Or6A+7ah
bxXzeRyI8oirH7A/3spQv+8Rvcu31vvT/p17a4aWkWuLIqPEJqJpHhiJtXdIfodb
WuxRNLqOCr0t9yUwOXFTahMUQtmKvLp7JJgWS2JMe6y7JyG+7dRk8vxoix1JqIAK
6rkVVRNbE+kochatgd3eEiYYX+8Be8kk0zZkeYQiNc7Hg7P9yko+wsZQMWfq0EqC
x8ugo+dwATaO0gsVVG7s1w5tdtIrmBHKaHf6fZeZzzKfOu1u2aCf0bSZdykXgwLu
OeVC5Cl5j6MMVA2evLM8ErWccdZgOjquqQNnhhujcqrcdPPCNqrB7LmXHdOavT60
Ajr++GkRxlw7ytpW5/pYehWc6Kw3dGxtosZBnqPyIS4A2NVmZy4kt71By/dewTow
bXHSA98X4efnrQESWo9VXjtrdCjflxLhsREQXJAj4G06Vik2/DulWyMqG+qWGSIV
n7aW7j2l6Q4jRqgS3tuQ+oXiDgpCycEw3iHXgyBvJPTKreR6bw7kyeXg/ERxEWB+
1by2X6aiCKZCI36U6kvNO41+qWM/EUxcC5Gg3vtzbwSRJulAfmPzs5NHFgs12RwB
yhIypXGoabnUpfpYSyBTw8ce2GXV8uOIUmWqnenvoC77sJjl8KOtgo8eNFQtpwcR
p72GmT1M0JtZoh90X0GeSQXg/zh8BMHS3Qr5WQJ1NbDAz5lBXxzBhWO4V/RDalYK
ix0dJSQs0D5POTnQKmkNm893yK7YmeD/U1liHEDPbRkprAiLY539SQce1HvKcbts
yAl212yRWsdU7lucozp7O7DKaHAwLc3wiB0x3sx2V3Eee6Nn2ZXHjRilJiGgdgd/
rBVnF2bFbQHN4xOYyaEJxeHClLyWfuT0lsJ5r+Oto+z8aPG0Cn4dI9G0HmEqvsEw
82dYOr6jQ6c6sH1iMMS8vgf15UVZgnGZeub51acOsz146/fqKqBt85GXOqgUQqrp
VRzL1M+YkEVlMBO+u8CeX0S13SFV5vC1m/guwDbkGuyeNq/6ocKFqIjukLps6tsT
u/dr2c0TvbOJB0snCR+7hEnJFbiqoaskxk4LZrI+ONOBQOwNm4FkAjqW1/Ed3x+z
4O5YGP/Rr5IP4tqOoGC7wyfE0uqdr8wU9FEd7lgcmwvXcHVx4RJqofJCqXE3+LM7
E+27JBtXNUU9DqoDr5U4RfqCgWLIIceWCjlvnUdesLtr7Wm9nyrjlgZcZZCuGKDW
Yam6jRdhRsgMV7cyCz/mHEGKNkhb2pWt46qMOXPHGleDr6XMdcQKFWilUkaoxCna
ja/QtsLSb1kvRRcwhS4Y8mMV52LGB88uUUO6ee0D/kVtDHmVKF0WXNMn9vpn77TJ
q3u61jSVk7AbmhntDu6q+3TlInPn0uBRHF3mwfD3km9Ak78UUoFBlnhJE7CCTIW+
dWELJVTnGPHm6TKNw/4ZfAIi8liqrJddvEQ+ThurJfotcbn/cYWw07oNDMy/kwn8
PDKQtLgGAAbgvrV0K/r7CPsiTAAPUUKaYgzC3/gZt5sfq7bDYakU0zfryAfIpF0g
bw14yAn/QN/9x/ECYG/uVwZZceSSAgQl6hQT2ph5YOVcsn/zg92fNv03eY1HvzyA
Jo+WohfyWYjdhI8P7/UbCMmOVZhR25GMEF1glTTacQmxqtfg8tyg2sM1rA4mFCf1
XWnz/c2BslewrEk+JUYgS+a4kPRU4o4BODRjo6p1CD3esQAad32SZXdN5JXU40rp
4WG/egU8LGFNfQ9wiyij3VhSOJ9BeGeuJSyMcznvVzoPmgHGFWtYWSfuA3oHU0j8
6CSpA91ZAPNL+x5WTOixwp4a7EpSL1vGGdvIwCDtZTwFQ/AsTKNoQ8N6wmzribN7
2rewTh2Gzukj1mTquPFvl2OAl/rU7ENLQrEZZaSJn8qf0d1ePzDJQscxfvDZgkgC
vYu/cxVkW/54us94iPxNDhncV6gbW8CVWT4pPavEhLK4vwmmB9H0BLQhgf7txGwb
sixSzVNleCc9mDAHEgMH/url7zYcqV+FlKoYn/XNrE/B6Ps21ah5pZNMYK8O1YSY
eUZBIKmiibEJlBsr/Yltfmk6tf3W2A7Kl0X9IGpHZ23EzFqx0y6YHo3iTsxjBZZO
DF/zarz9I1XTTOKU+OZ4gbO77Bzvzs/wLxNMixh7IPH6JY71EgX53wvu2oqdXI/V
VpjFaA6XJIP9L9lqvi4YMQHA8lu6gV8qnjinhDGgGcw9hBg+avljW/axvY4gFJ7O
958VGM5Y2jnAA4/XFdXtfLTmTsyFFjK1ZzFmlgJ1sA1OS4e8obiHRHnZPSLdR61h
i3qRXLkwv0Xi3n3ocSvxax0gJvfpWE2js8jXOBUw5OxOgXT7Npl3szeVKNtSAXwa
J8Xz1CeKCJoXpI4LJLlc/Q3lqobSeFplam3gjkhuYI0FYKhbmNfCGOB5tLvpY5ir
rSEuMHPMHuIQmPziBS8afX0j4bGtAvk+2CBM8ptDcMTum6xN3ExZpi/hVrSPzlwz
X3f1ZmS/yUlx8Wygmxe95R6pSQHHSvK0H0w9n3FRDEiVj99jgarLff1ikPSamFQa
Boo3tyCmoHBhR4392bl9fpyYT60yFRS9++D/OdXRBXr9tsWtsxV6ZMzouSkIIwWD
15li54+L5eRoxAo3l0txDiPxkevsLsjTcv0wbJ+YJONIAPqrGVdZUgL3WIRDDx+F
dX2YMfCJkVAVY5sd3Ip7gBNcjBnNt+AxUpmM/hmDj1xjueI0oVdPThEIWEnJhrZ/
xXm85nFnGJ7LSiYnqbCJpa2fzPumoZf3XHimEJpRKHJgRsmGCuqMwB9qroCzhysv
xnHJcDO16Lt6cThh6bEPG6VrHKyPDZ4/UVlG8S/iEW9y2YHgnJ1G45GwFAsO/Aqp
+td4irGRDSNulDyh8mt3Gf1Jf1QvltQ7rxuaF3cEdubPJW0rn5A+C5Eh/s1lyKH8
W8sE0n9+z6amLeBWnwKPZhifqG4dJcH+ZsMbv8XJf/R9t4yohv5imy8VbNtt34g8
DkmzvckAXJmAhju5Fr7tp02bu4dfC+IcRiA8uLYmUrMIeOocOjDRsHg21yx6fGoZ
7F/c9bAGvaTOHSUe8CeFY1vIkvxReoAt68z2dCOkrvMDhwW5BNHC9X46uzIGWMhj
cqR7dhqeBJDHmAJgcSMFpTMGUclmmSPNi7AyfH8dzNaKwRP1HXqJNb+mQdDK5S9J
n7ommTWFg/q64LzFn20UvQZMSYJYYXtdSpzDCV0bS4UWFEI+AOEn6ZWyA31+mw1P
BwPsZYq6g2TB592/6eXtCnWgQBGtzVXaetEoRe4sb7qe+JHf5UIh3tA5dLLq9SEr
TiRgzH1eQdJtjZocKJHwyB6M6ev/iRRDUa6fbB05+EuwZwUxCpsYsu8/9tSK7r+0
mOIh1yz41UmjFH2wG7WB7TtT55qGq2PAfeq8RJw5SJb2qc7fUU0CzAN7izvBjvGM
kIWjYQDcPOZaIBbERyYAEoiQmX6waAAbSo3HjV3dk8rgxuvlV3Xn0sioA+a9IXof
b6L25f5Qq5qKLshkDD7tjVK/zfUpMY9dguQjqZcpWndg72SxhzWrkrn/j2uG3BqD
eakpyJCvKO7hYs+OFDRLCIuOBUopweVZOiNW3wwL/y3yR59YWc2Wgiv8IK5hqJIX
BrTEFavzyK5wpwLQAVS179DJ4kvNVNCebu2QrAacuG1HGd8UgY1yhMwLXZUHevYh
Q22w02IMRCezt4wYQ0/IBJXIIaJp0wMOB2cOxpQkwcjsaCVroMgYn4IBa2+smMXU
ksT5HpWCsKE/bGxnuygN/1Q2WEGp4C2eiaUTO2M9yCZKpK5rMiGywZMFkdkYYQeD
uMXPtJG/mhZvz/lYg2+QBLDzarTwWvn8Khh9p7+XJa03/1ZaQ0maoHtobM16s/SH
Q0ZeEedVWDpnR0lwvUXpmLtKah3PHcfy44pBJzi3FEi3BZCEjTauG0EVVh1aNMOm
gX4p4xGQv/7KrOxGknuR2X6vFqUverjUbuzI0OnU4f9IHUfCBV1qpWrwAQEVU97g
RiGi0yle94vu0C0jL0y0EtM2EHQst5lv1Fr8HuiNhEW/o024qc0veT/G5fiLLFTy
nNIE39MeE2w4o7J8YfqXV5SS0zoGFevtXwmCJvjRsLjACtznXoZHK2lESp4VA6jA
si04bTxoNFxJbICAGMHo5Ek+wCN8L7Qt9ZzJZbNvNd9+LApy/ga2p7RwJhYBFN9G
0bX/z0bSxbO60+MAgQK4M/15la7wNWvWRtXgIQoHBmqM+NhSWS04nvhVOzGS3zNr
n52kNqsgtKlUyXHuhwHq7WWB1xB8ipjqRQYJCv8IYysBNcpi0HTPtpryES2xrZa2
PEpNLEpqcae3Eeo9nPfdDWtuIZsC8sFbOuAQZXpr42vPLjSKldpQITaikUy/x/Pu
WxInx4UHXq+lgTae6QKmCRtuMJ6h6yKXAfMTO37qdjXMO9ag2zI0nfjaXoB2UPn0
7z2WjvXcIsZexw5SUfOdMexLCAmkDx1ZrJ/N7NBQ13pKQIExccgYlZ+7+WiamZmc
p0+Nwxtx9NnUxy7UgtoKE/aU1lhUV1VD0UhFCb3HZFVwcllPN+aGEf6GvXIV7ajD
aPuoZcL6z9ahifZS7q8RJoHlpDtvawwwVntThgq8MfLf47nfkkbLmom/s3Wvj3lv
bahZ/s37dXSfQmawVLv/m1nM1v73VmNYTOUYc87C0um1yEu1LFmn58Pm03V7rs75
8iWJoua/EhG0kaM7r3G4JEZ4IBpkFojX+Umnl5q7pertxhX3895dO49kk767yy0C
I3OnieHUvp4cM/L1o4HcJuSEMcyHaiwmMIMPLeVSjc/eSFfigobIZuz1/3FbgoyV
m1/xukzCIj+DuWKWPmnh1JJ95KuY0uifwWZgDpMEK0DOJvcYDmW0Kwup0yq1NONF
Kt71XcCOzQWFO9sIPQWA1IoHFZwiZn/8OmkvALibP13X9ZixLyMv3TvXvQGajcNs
8B4vqOLOcnock5jYE25mvR2sdP8xoG58jaL6/2p9d/VMhbeNvfh1BF/5XBdnlEV8
Ky4OWdpDrrc+hzu5tslrRtzhcJQpuDhPhvgzq6+1NlfrKO/Wo3TWNjR6BEHWSqzp
jl+4lD6Q7wh2+uRk6pLSMRQrUvFvWmtMsTF/JfUt3tokWbftH0pEYlEHJflm8ail
XWPVg+xZvT9DYj8pLtDnI3fuSi0Qh26qVxlfxZgCws6ggCHic9hrGsALHYhDr/ag
b0Q0GMHalDBgLgMqiyqcEOSybTkpuvlUzo9reD7Gd2Fhr7vilgxlRd8dr0hb+3Dm
V0lzy3Qwo2n7JF9nt5tGAQCuTxU4IwEDI3EW68gBnIOvUchbqurQvgUlQpvT+cim
wuOLM3UsHDZbq59o678zNdPZDbH1seLz0tqeqMZ0DxV65BfStCjfpDT8xsVKdxKb
Lww5OpYe7QDz9PxDStzcKt7begYqwMjviFcLGyE1Hc1ycPPFA4P98GYWPsoed6JB
ZbD9sx31y1cL7OLbJchbV9+mqpSpFvfl9MhhVy3HIPnrSIqXW00pSTov2zL410Bp
8MFNQihka/z+Keuql2cX2BHU57gXFrarnLoLrOH8Acm9rMa6IPmlYL8XYcqlkmRK
frVZmpeNSbfriI1SfnVBiiQmg7DXDIOxidpXjooYo14KPjCnDDs3jjKi1gR4mbth
R5n9hefBa6OhcqyPZgSRJ9nLftYdszFjjYJ3Ye+oBx9wmusWjcC93fjHdwcR/Pzy
5L3NsTdLzHmTp6jG4xIWHiJrPPUE2nCNPMRl4KhiGXgIU4xDB2HAaf9nYOjU5Znr
Op10i5oLQRBKD2iklZxXKkAHBTUkRMzXFcF0/PbKhTdgLjMtFOsY+W8UHlPX/2Yb
HdtTHX/9+LfpsyPKNJFMriM2jeGcOlYO9Zcax9n8DJSTuEcngcNngLtV+YjYJlFA
hM2IvR0cpkRLVcZO3BgZpH0Bs0CTWdLpJRbp1Mmt0kkSVrZwJN2ae4UpRcSe9qaO
qBmDVxG2CHOAjpbbmOZ0fAN0a3dwAHZhznQWE7K9QAF9aolh53Bpm1Z4BZO6xMmY
VeQfgwcAUHU+wctAZdKXHZi7uhVHjJqhUElkL/ZcsCLUzBu/6IT4TC40A8G3AaB0
fu8n8Ud9obtQAZnVe0VTTn4sdVJE6IUlqjXbWg+QcE8d+d/Ru+4/i4BsEeG/YIQo
h6HYjnBwgCtsoAvNcMR2fjaHUBHu4x4QFyPs5sAqRDn4bmhOKy0Pn1HzQ9ycrRrC
u/iVG38aLicwr0CYV7FwbR385VBKjJz1ORIM6tRJ5S0JRhAIdIH0pv9kbZ2VHgkr
exaK5XFpGabZ33mfG0mhZOPtrETn8xLrVUHfO0v7SQUF8CBt4dp7RBbryJ+/9zL4
YRGPBQl1lF1uu67fbLYd8Lk47Y5l/Q8vv8Tvw3ZNRhgYGYu2qPlZZXu7Wci9rOQ3
IFkEJIsr4KxN6Mpza8I/vUMkklC98SwJw9aDpvvIMruBdtXot6EpCTXHtIyhXXLo
Z1WAkN183UUxpYSU1K6LcZqz/xg+K3Nvhsur4d7HOMK91ZNduXA6mcVv/HhKvfa0
wQb0qckIKHoGx8Ix8lsDkr2oeQ6KCaJ4Q7IoR6dN8BGLbH9X41rGx6nFCTUeZ2Sh
Uhb3vs5w9lWQPBnn/uVNGKNybvE0r3wlx8omenQhXntzKgi+AEB0swQaS9J/8l0W
GNq9KwK0pjb9mMJImMBllJC/UzMjajM6B+rBhnXqwDyoai81R0lETGjRzzAVANvM
A1vDxMCESuKEzemo21dKgU/CESINlj8ZItGUx9LonLqg3pwC9HfNgnEJ7a9Xlp8/
JK+VvLrwfbD7ud3eEQYXc8lTNzLwuVlAXrMTUwtmmIG2kDooAB1nr8z1nNYCQt5+
wolad/6ZlR9/yj53FAPTUaDXG+cmrcTYGhMSdZL765CVHdeGrD26C0tn8DW3uWLG
PeZbEhqewp2j59jfx4UbLAosCvNOL2i99/kH3vocasqHOUCxK+Jwww/xKJfHgBV4
GPvkJAzqpX6trf7sl2Fpdd4ymfXn63VR+RTpC1rrkjj6/8GMEstOGNHcbL2jp7rq
9Pt/zTPA1GCsImKgqlDRxPDPMglFbKx541QHtlPu+s7vbqJGWd6VAP9hFdFm8iz6
JRaBlyPyu+BGj2gVoo8dd4jYvD3ym1wi0zJsHWadqPUJjmvDDaYLkTCZoNYeGLkf
vTFvurCtbsaAXS9Ypey7naZjOExWA32DyP39oRIWcYOqCmk+Lw97bfOJe+Pq+4xD
3qhN2k+VQj7sVudDK6aV5TWvelbWk7MKZ5gcgk50o+FKipMCWTjCj7JyhV5EPEMp
WvAkKiPC9Q2NJXVkgr/LABgx8/VD1+ncS8TXfyzPQENKLGW74jn4kQ+ydYRMkt0T
xZ29MWh4PCBjrFPkwRBDoLDxQexoqOYu5rPVGk3xLUAXhzKTiy4bGvFiFmV101SA
HhJJCo3RTMXmLLv7V72vTrYq8u+sreGKz5JDMIv5+BH0ktS2subLcon4aFJXBXkc
YGrCHINHrQR451j+9OCYEOPrtbh+iHezaPWg8oiMQ3zHp78XBk/xkDCHwCcWPBfg
bMxJn+0gB//AAwsusJ6vArbjHDyOV0YDVN3DolFQby8TEJ0yorMUKAoo4udmz9+o
3LxswlZWcGIUAilYX1rjnOM33hsle98VSgFMJx58lqz/cc4B/cgXgp28jOZKMVg4
XO4pvUYqVjdIcR3X/TL1WgFlz+L60wWraLsEAMaBEDqVGfbYFVtol4RTfC9CHRj2
fmOArRh3+7Q37056r8fZ1bRamGOp/sc1UuV33xhWFgQcOTZ98n30Y040QJyNq7Ou
kpz7R54Ytm0384+4nynNSpaahtn2uPXtdqOra00aBnjE+NajZmXGj32YmlzOg1IW
P+qqtM68G3/G7lCCQj++YP5+ScTU1qdQ3z5VsVPkwf6WNldOJLpJXTbxKi5yHM2p
r9qW9Qs2FpJsei7kJJgdY7UWPqIV0j6i31fLVf3cgOWXWQ7kOi5TwtXElJUVh56F
UoMSM9F99rfaJnMwM9AQbgrEKbVHKLEkLDvICD7dG100xl2sAKFq/vp8oeatFtky
XAeWie1I57eF/ZHRtRMxmVU0mDNJWOZFSBmoW95XG6BN7bXGNCFzLI4WMXjKTEXr
WamBmjaopTypy6NamzyNmdC4rueIByaX9Lvx0851uXjsvJTyeEUd6rtf4VAm34RP
jCXY0/RC3Vz3KWSze1fsRD9b/iO/KteE+wp3JAZy+OAHYaAVQRJzxjgFOCocUpxg
x20qGue/TXgaGTN3zWm64PvSJ6iAbPYEAXFYIOr15Z/WVTCZQSRY2X/M1dsJw8Ko
V5TnCsFXjlIyUCQ0dXXl1wvo3iMticmNcsN1DTCdf3UVgs91d/I2PrXP5UgPjNFI
t2NXI1vBW3U8YBph5X9QLXBnxAtK7WmJyL634AMs+Ty4a6UCyr/Y2iCinatTcitJ
6OV6CZlC1iI15iylTeSULWLtz9EXLefM8geVPmV5Vgd+xNZD1EAfC7vrv86ES6Re
rGD+I/Uo/Et9sMqp4bV9Wze/6IHpbr93wlgvM03ZK+SXcDu3Ad/tiyCcVOkeviAD
j3ZnLDTeloSn3StG0jGLKjAAecebapAft6b92vklAFf/KNXZgNvkrObn9ryMyZeR
1SRpnFsPH5OlJgDml9BQT1TMUrhf2IFgsB+TY9bwAHILDVL3WzbZ+Bh6+uFVhLqC
uHq2tE+QTCYa/lOy/oXzSdhUe1AtACERucerTwrkJqSlG4FjMH6EA7RbMLeHYtBI
SD8DtQellaD7INQAABTr0mybw5QgKUN/VoemqIMmwlssoVuI6Q3cOY0CIPaPKJ5+
kJTdmpmep3j1/abQMFqX9VJAVGDoHtxtYfRNZK4cgr7R0+nWVVm765hzH9s7bpAo
C7Nrg19CcWr9Skf2hefyvMtqjTj3UJDjz9N/IjiGED/YLjbzsZlpnlVd5dN42VEu
fkNpfomk+RaNWr/2olCjmWf3EzxovV+gHj0p5ugO1IffM6ZRXvXp1AHl1o6kOQYX
SZvSQuuDmV/KM6dJ+oMOIMabi2pYX0yROnDXWnh64yUmrndJwJ7uUtD7Ax752aLw
RMR3qM/AYFajeHZniEOW87QJjtRQJwgpdjpJTz4ji/c0jBQna3UZTInqqUDcxX2R
0DYdjCspKhq7PtsOFrxutjCkdHaSDbDcd1KX0Vpev1N/ncG+HMBQ8zR5qWN8Q0DB
7i6ZIHyv/3aQ8FGQWaZ66gHfLn3rEpXYUVzXYx53uHqGXjuFOOw9dDunJnlNWGhM
JoCOZvmZ+vtSBrTm5jzynxJ2mnIsEm1BdiYbLsyH/XmcAuQWngGgn3OGNKtqY/xH
ORRJdayRz5LxyPTQLgCz9mhWwZFbO1ikHqSN5ZQd+29Or4Fnhp6fvo9iWdgOiJt/
RNTpmUOh6A3OrlWpba41gwCP8z9zbeymRdeZkEEIPx3IzBmFnArH4uUQGiYrW3Hj
a7XdpI4pRITe6TcdW6rtc9F/8IWz6P604FI3vCfR7lEaDjiRzWHqmSYNrn1ua4sT
gCZHaFEZgMvu2lHblsESGaA2U5MKJOmnOBaGWBSRSLxZVkw+mZAP7QoXHcdQM7Ks
oIDvmDWj6hAejcNeNbnLKbg8lja1sMC9IPLwoXv2Tv83EHjs95QtetoExcU+bw39
SLAU7mVCUP1iQqA2S0fAGysB/ESX/rqphLkAsG5oB3/xPUVlxwOb9UpFqXrRKr7a
u2s7Porx9pTX2UnbTHcRPGgDEyYBYVHmZyGE245swlrLO5crKx1ZyDN2Gi3x+U8F
VoSSh3VVXprwJY2fYXkA/iuk24+LijL+aEGMDb+8Eejypx3h7zSaU3UzQL6gnBy3
WLu6l0ULlg2vlbGU39NdiPXSKcalK4sDjNJN17tm5We/Qpl1auqU8fEXuzsTj9AR
HwVIOmjgLh7ZM2PFR3i2HUYgIXxo2odBvZOG6T+btejg+o0y4+uZxa/8ysXFwIvc
YSkLallADG186v9SjNs7dvygkiUpo9VQLEXkxq+qL5l0pzB3iTVWRc7kBBugoAkV
+fQryQCOjMbDO3YxC0hJbSpNrlBIkGOR4pVEuhaR6CjHX8VOOERWHdfQlhGWyYqY
vgF+S1Jx3MkCBfM38KE9Uo+GS1kaAKuLIiWJ1WIU8Q0Mq/RZnGoVpBgkvPPrnDiO
LBBr0nvceH9uYF9R53N6NvMF7rQ8wxBx0Q0exUWtaGGsR1kFdHfACdi9qXckF3Qa
SswYWHv5Sf46Jxa+cAjHu111achEon2ICdUkh4Ij8uUrQ4US7JxFqTxX+2va0a0c
7M8cztDR5DOMxHEonFAgL36SlvhcthFvOyNmEKwL5KDTlgnC9FNJ2fWUGZLDDHyQ
UecqKVTpHEWLUccbXBJ8SRG6XTRDrMgL3WUhHycNybKcPJq1z/bgszvLgSlh9q4p
vMyyOoLtC6o0rq1dMFmulQw51P9qxVGLjJ4EuJpDR85pMigjSWauYZQTRQ1ZF2Wn
DSV4Vxz9oguR9PYJVxPy6UNPNs0OHVFKc27KyOgyyitua7wv8JertZHk+gxaoOMY
fSQ22PsYOiYhJnVPWOhAUui1OHzeMxSaSw8KTLLcvv54cXEtG/x9LrXQkPgqcpMu
nBxeQ+ZxQh/BwRmEsLfafvtWMDlKhmDqJpLxuSjHfLNk745xz1KDGzAJMjZchZck
LkR26rRBNWuTj4SMd1vSzObXSQhQuiSHhDhWQ0qDJ3wN7+WdyxLDWr2S2tbkaPA5
ciH409fBlRY2Uh6yBLNYhz5vnoQmGpbp9Jc5hW2Olgr3//z21RUhXGklPRhJVjOa
BAIs91CRQm4O05gBw+s2cdCydfNDSnwlFd2NhCAg/pwOh+NfXPxQgxrAMl7MpDXA
O3VQJX0jo9RrEcY1EaenUwlQs7KtYzgHHf9Au51WtRY616amWyjJgODea1X1sfr9
AcZAas9Wx6hjliQb8+mBfNdG80rhEK1NQ1CnJZc78R6p/6SXX79Oy4xEWrsST9w7
3hkTxUHsAPTIxpoLB0hkW+aFnPi5XcIfk6jh4waWht4UYtnAzkeqdeyr8W1vpbxi
KJ/LYISFQ7kmq/vBpNMzfjcaZeW0QNDzouDqZwmMZ5UOEJ/AM9UqhP+4WFSn1Eo0
38EHtDJ10x8ISneGI0FXNSrr4RxeQNpmjYARaHZk2BdxMgpZMKo12PCUqp41zdwz
ZK0HpnKAknYw11rciDcNak6OelzW7aP2G1N14moYzwAWbXuTsOBDJXoKSt3Z+5dO
iU7hsO6BbJ/V5QX7sNCSUY6erg9HGBmB7FTDQmhwQzIUcrulsq5EwDGnalI98oLW
PDbAxU9v9whc4Uj53c/domsYUZmyh6rSz3movbm+WUE6TlHeyaAxK3algK6FOEe3
79+NrtWgZL8A2CekmfQ3pw3Idx98qRH+nU6Qe/ozcX+u0MGgt3ns7T49ZJb1lXTq
khhZnjl0xzcB9voq9TH3AJTnP3J43yUA/ez1Ca3L0qAsrNY/4Lk1Yu1dpbni3+2Y
mQR3qD4+KMrs7UADn/5j2QQwO31EEVp9OMGiYcDb1EdOdLt1XEvhgvlA8DhTyPz2
sHXN+KPVogNBWsPmfe68nAM4S//9ewiyAl8hscyfCpxHRO+BH0+eWzIFv1/ERDlS
O630qZfezYBX5RkUYX9Y3H3kU9FVzPE5BSY//g0dV/Wez2UYbC/VU8lfwtgLTguN
JRAjdCEJXVQCyUkhR9LwZK+Rn7nYVe+zorQKb+iXIOGoQmV1Tal6UsJmBA3iiHrO
TnNaqMGAQdM8ZXP+5GpX4bPfZwqhKR/1IRoKDyvx+JMq5WqJH65oxVJAhK4vWFNz
+T7uV7GFf3eROonr6flbaDPrpYqSZFnFIe10cibAJ6D0KPCjILc8pFsfQohtsj5t
b5JF5XJc2Br69+iOWV/PdDaFPlpzqPFGew2mLnMBINS33I8f4RMmYzwpkgJ0ue8x
SgU1TBzpMehwKlfXGb76g388hkgZpqgtIocALMKfWl0sNRIWLEUkz7LAnNN70fiK
oUn7RKD7r0HdgYrFRaot3F7Gu66wTECCkcQe94ZHKb6Fkjap4PBSEJ/P1EqEZBS9
QhAFfh9eNMpQ6XV6OboqddFl/EOBp4dv0vP/PQATWRzXiMfaW83vNFo5B6gL133k
qSfI0n+IJrFsdng8dRmqqACL6zt7HTjNrpwpOAuvFY1vgpu9G81NBVu2GxfrWtFB
M4xIFeP084nxINLBoP5Lq113QZKE8axRHRx9p+JCES0RejdjsZkwYeM/X9W1Pitm
LavTPPnrSqiDoTQSD6dLqQRqMOUloPMWexh+P21dIxKVzutpkpcCA64GPNP4DIWh
zmKnQCtZ6hO/TGdfYw3CnEXxjJkUSqtnUJqj2IhWHeGPWUntvo/TjU8HiEsoVIr/
gs3z7JG6Xdb2EWfAf9DGwcHXm/RYzaFttXcqoRUgUA2nKaURWnxyUTyBZQXVggE8
T8OBv2PJju9IbSEDrQ/imasac1YV+yaY3exaBBb3LzOTAEXbxObP73UkeQ3Yh4KR
e9zzntKCzCdXQHOazVyYq+msAD5DjcEXjLJcs+JUp+di8BqaGy1SxehzmMaT5VVp
v+KbpWDZa+DVxBj2z4v6jEuquajb5zClF2K/cJAHQiPOXRYSahorfDqz2tjew0cO
8BOTFR87g7kBfyn4B1ap1ap4oZqVYUq4ceLRY+EkjfSoagyVLdPSqvkkc9+VZ+DB
4kY02AkBuDES9WymC0pOYUFJvNeFp2hRWt47hjlhCNlkaGaczZ6xc5YLu+eHmDdg
zbcxdmqygaFytQ+6jM1Kw7LeWp7zgfZ/hbGrZcudMBbI7ElWwTpW8GMWxHlVv4Xu
CVPV19Jh18NQcaapFiMU9vGd7g2eAVIjgCAsq6gGbW/w6r136H0w49jbHK7anqSm
R92uaJ9zZeCPQzsap1gWCZYyaC0YSaYh2NEepbXz9KR0E/+Ac/ghyeY6lBR+XCyB
FXMIrOowsp2rzjMTlEG6ybHKD8xSzu3PVpEauaBY/78J0PukZTDAquw9uyVRsCRf
RRyQ9QZqxd1RJfg7xlR5VyceYBudcOD9avCoxidZ2M1UlInocriJdHoaHhRbsZvX
M9DuuhgRCN6GLbprj573ozEM24bU/15in1dt3HooqHFIVfjc54VTkfwixoosv9Nb
U7U7oPM1vDLeWCbsK804g43R5FBhpa0uYMAQ688ICwmb1MzUdH4pa0RpxmIgCtSq
Z0OkITErreg+QRJhnPMPn/ezSCqgoxWW4zn7AGFrJdpyOYdWeflHZWn26E/KJAP2
V7Ky9JkoApNnP3WxKc1d4Lf3nIJT3x9z+KQMwPT0C4njVZXJf553saQZNBB/G6Ra
cwCrguYZc6Tslx9oQDUHZ8dQMYRzXDnHP2Krj7+yFiKIR6D+lobUms0xBdLCK8mN
ARcMA504B2rmHwWUTXwxo5CoI1W2UaMilh/cdd20woEnESIXSdCXKXaAS0+eM+p+
Xr6hsbyfUCSKzCumhEUPkjbsE4ANGW7FFiV/2gUyLk0zbXUzEnJUtDLtowssEnGa
qhDmUrckoaVAuvkNkMcXPznOXWMZzUYQBmbB45YQJcCEi24hz7diVYJ91igkma+k
OVxfYZAAApB14I+QWQsQYPtJtkFiObFOzQhXIwyW4hS0ob4k/xxiH1w1udFyMkX0
jIkHvGCH2yLDI3TyEZNtmnFyrkfjDxzdMX8OHDgFZMsrKIx+q2nC2Fp1ax3CCqUM
Y2un6VaWmFkldW0VE+hk93omyKA8cx461MYLGwYvltIJqkEoefN5re6oYm418OfW
BJR6beo/+KHMZ34RkeRAPjBzFon1tEFoN8W86kVYdqaJjhS9vFG5pgNsVhgRo9Cr
MB9RiItyTiG75/YlvwinFqGYWALRFE9Oeb1apt27AYNv05B7s0NoaSYoa91UpFlA
orePIZLIQ+Otn+NevM3yeERijZ3pwK2DopLAm15IysjG/kYs8Fr0O8isGyTk4G/U
Ozx3WSayll1ylEZo3sVeUYjDLDJrWdlG0AhqzhjVhT5c9nOQWEzlSqaj0QcBESXB
Nark6QIQUKLQ/mAtzo3pm2ZT+xIkexgT2VWegKsV0e9sYl2rB3F3XCcoGOPYjRcC
Xzdj5LjYET7fmPxu1dhCECeWSbO8WK7s7H4eM828VxqwqpnB2NIXLpv9FoU1fJzV
7bs7iUA+kZ4gZs4wl5zc/emC8taL8teWQPRWU5a4+zsAeww/Ryx5RgskrEiX0mBz
aPsbae2P8peU6WTXNR1oJgZgn2jgEswqnhroXtEDi1vZWIDhfiSARpkFvZMhroDU
Fl02MlAdL1Z/M2uLEA56L/9TIinlbe8WooB3cEeKKCH6sa5ykozHrRkAmt8KwVdu
oPXKwTDoQM1ITEuYx9UFCiPPAmCKvemgHtzb3nOlphuDQvheYbukqR+0Z1FxH4d9
fPP8NMHuXnevqupI1MyDEdvPqsLprGoNnlIHK0GubNgeonLklclAU1Qdxr3O+FOE
KXBwHXCRSx4U6msmiLbvnuu53mLLt/iPqjXOnQVAZrhQrd8yX1w+nCj0SCTNg08l
whKerZt6z1bsX3e99BBiIjxiGXELwblGWF+VOYjyBN9oI7gAxqfO9pWrgzjyFQY/
ZgZwD4xlCyHd3fByJttemWhJorIs433qtZr/I1kHUC8swI1tCvVsYU+wuC0RJpaz
XTcP3efj3b1JJ9Ni5jvKvWprlrgEbLyH899O43h0kK2sUzIkON5V34SMfeoHBjEJ
rQfdXV1Buf5hX+qy6xS69yMie25HBOh3+CIanTbJZ7JzBBHP347iw5UIL5Uz+3uQ
x7jkbfNUXOL3WnNsQPOlAH+IYuAL97C6hxt1x8/SFQKK+oS+REe2xrI+Xg/POguj
e0x+L+Vpb+ff/rZX4nGo16a7i/akTbcn4ndz6JVzsjJ6b0EL+ZRISwqUz1cXaFVD
oFBXUymI11AZkCAqrlHnvq2cYiKaQbq/hZj3AFgHwJYeaTVN2mxyPq20JNoUDVj/
5WNyE+1LFgvlH7EZvkYc5l2k5JwZ7FCYdGKToo08W103aijkFlTw9Rgdh7NqUTXA
BMPt+1PMeEGK+GoROZuwO0SEVUUBMEk3y2znSNqh5AN45A+iEWHlLlODBxnMdOvt
0wN1Y7Em1bajjF0AGZs0viSWIY0eoVGuK8v9h3C56O0Q6gLHOjZz632XKB3zN0gg
iH5EO+m83he4MLysa5m8ebiK+h3sVYXA4VSHUnC3foevsYVJmwFitz+wmD9zZLxp
g84A8vqILKrnrvshseYe/5zQSrDoOuhmneqGvMVBO8xW3F0zx/Bs+nVvvwC2C4J/
ePVxCncRbGMUD5Edw+N0C59RpSteY2r2WEYuGBFxeuE4UIQ8aLmz8HoPlR8qLxvQ
zJ5bNINc89QbUQuB7LOh1PLn/Ghh/+Oxfat3qaHixTCPS4/6pZ9klueNrpaA95VZ
pd6OUpeigBgs4n9oyFU1yuFrBAK8p2GAtATjOutvEd3RG15EkXhNpToy6cLsnMpm
qVfjF5nE3Vsen1K1e84MWBAAow+B9RptOZgIyshiAnWMsDG/rlSwz5b55fms/5+L
5nRlSBiQMCmo8Gha5XmntSNYsVmeV7WTwPsH2j0Dtu/hjySlguaWcALaydeU8jRg
r9R8MIqiU2f+U0zKCGjKaUJPSwJVrNjjfSFH3+GcdcI2EJwJLQp16pztpkASxWk5
JSXl+dy6Oncmadl47lQ62CmTekOQiWY4v0o4EOWFy9Ox8ljjHK18ZbLyIUeSdM2j
qdfpHnHjmIU/UVsbkrr8XL+aBKng6ShBtWrMNTezMU/FLaf0FpYoBqaRTlXk6ArX
Of2GHqu9U+v38p4maioqD9ta4xg97G+4x0nfzm+wBo7LcdZVKbL4bmInxrx862hw
ya2WVzJT3Enh+WMr90voGY51yqvvSmZyWioBn8Z6lMTht6U3rmmlmEYGP6PqXVOJ
VLp/ltSk/n91OOzAlP/gT3dQq23jXZD4KzPw4ixrdsMRAgTmSkbj906lk+kmmIQZ
6NJonw0LBdwXXZNUDBCBP5jcOr/OxwVnVISBb2FkgHrdSx2gMx2UGjcNgcNpjKyq
pg6uAtx8b18p1MlEInQmoq/VtIGkKh0fnFmEIEOuxB1mfd2lvSxPtFDwyCvedVKq
2tx2R5zwl4vg5PPjir3xNeesS4M59X5wRajTea8AgjPPce0ISo4adouvOwHtaP7x
tcvtSgbktszC6iUSgWES1DN4RZNi2M1d1BM+WpqayS33R49BLxyka9BHO7xQLU+P
eP5fPbtKg42fmkqCCJhHNFcqe4Pakpg2Xim/CU3fNNzq9R+qqmC353x00DuJKwdt
Cb6Tghw1y6eZaH1eO6v2uDoabkQbruECTgkznWVFPRbh4fHM7rGoF9DoCwD3WzGy
dTyJnzpJdjQzVS3jMbH7LS9f1VZE3zzqFX7r22550g38Wayykwqn8FnE7EHfLjkc
deIRLtdpoUkkUBWyECWrbNdBtVejyecro4lY2RnVzLlSKFthBHPHPL3zsEEj6IOv
LkpM58jJQc0dmZmb+j/ehVd97jGlMmovvFFn+vYe9Bm7agzwlgqHn9FRlQpPs/m6
gUB/a41Xj4GrZbAj3niGMNttYb2Vw7lDKxGW+od6gHdy+YB3v3exxebywW+UbIgR
BUiFoLiN98CanOj+681MU5lkJme3ajAu7Nv9uLrRH5VXdtY3ufESA7ZRRVk0YA5+
wpv0yv3t1voVIzhxpaDl9SIEqmqIfilomOLvpFnaCck78iEbeMz4MXEmZO1yVux1
kHz9Jg97tBANaSKrKKIh4FKg1fPwIkRPl2uLne6t9cWnGA/yh47L/2hrcRMQqVBr
akiMc5FhdPB+zULdzg/1w16HuEZe+wa48cy5bSnViFGYPZ3FsexMt7wtLvQGTVpY
1O58fL0R6eavDVDL3HSKIhxCt0QkO1Ds3m6ZTX8imHvM2pJhec6ADDTh416p70El
/rFfwGJ7RbELEUzNdhmIFVBb8JzHkGhjtVsPMxb/HfIr8X1eFckyvOCJZayc+6sz
EuQaS6uRjks3cVoJsozu2gAqmnLal3picrdvpUg2JJTCx/dRYgLJpXK8tbGMhDfs
SWtx4FAy/LQyG5JIkj5GB5DZQNcIVRbctmgz3SH3T8zHcbF+WLxfEHtcBz/+b0OW
o6Wom0UDHbuSQiAJLdQAt/+ZwwHMQr2LLx9vE0ZCoER7itsQdFf6vKgE3jVSU2ad
OU4JdLs855dfMHyANxpX2/rkRYw0bP6lN3GPiekdDx/GkQFaz5qFLdkyDP1/ufAM
YWgESLprZ5DqECZHl0xSSa+Uq5KEc7vAoh/AlwFaWN32ELfFxqDk1ScMN5B5RhQN
gGlBPKoYWHZw92vV/gIWZ5V7UF74J7ntDTRQgYanqhQcWUic7GV8uujrcGg22HE0
162D+1tTHamoSM/PVERtuzC7Z0p/p3LUE9PcD/pIEYDsQN7j4PXGEmxNnBsHWZUJ
KotgWtGheDQ8vuUwz33jvb2weXjaqMiXTJm9qv9mSnuKdEeXMt2xfeRyFaS08pxX
dWtA1RSSsxd5H+xjLoODx2dVOBGmAap3sMbBrgeBejdVnzvgyt+YEWOu2v4XnSYC
svAUodfIIYnkUBjGfMKxc3CABBXmbtOg97X4yGego6a/5RYLFmUE0kkN498HMm/V
aUuaEsAoqaPqBUQV8kkf9K8XDWyF7r0lZ+71pP3eV48mD3sIWVvhljvuNx64DRVh
bVywF5XX2ktgkqu8gvoGjOwcNbZA7GSClCXSwjmikF3PaQUP1rp8FrNmMwVftQRK
zh7+t+5tZfcwwfgXXU3s6/mTrvacoJrZJ0HQIWfXCQ36jwbDgEceZzU0i+q8AyDo
oXmfT05U3rgDcPLI0ZKRh6PqcHX4JXN4KgCNgZ7csNcjKATZTTquiVqWguaJ7UvU
xsDmI6KWvfjaaD5nxXuByRSBmoBbd/s+oUlPL/0GEUpfzzfuUSB3/VKupKe/uNxj
06C24w53MUOX5Xnck50XGpyHOXqi1V+kyhLpJtJsVRWlrRihPLbcN0JW7gs6a52P
UVkBuVTfxnb4IUksKXRpFd/SxYM9Hk1BDqvyvQIful4RDdmAWWbpkSRv3WXSNxRg
VurYxmxLPpJRoNuw3qyGfQAktGqLnCAxX2pqfAqTHpr1OB5vycvGji+q9PC8UHg+
wm9Bo/7DJ0rRSD5Ne1QiRxw2yDy3KdPc5agOpPYia5CKCim/Nk1lfav5IjgE0Kqh
6EuLa6iCR6n78239yj4jKYenFdd9MGBpX3YJ44FeNJittZhcIfqj/wqRLFOeTqWn
sCwqNdca134ihAJnkCOfHeo6TTeF0S7B5/FsOYrEDUInJJ8WuNJDaLyB2O+o36So
huclLNkpTdIhBGjbzlru9dPbHeCu9EjIG15LliVV6TBNXj6B17gWKcNsfhQMKSL3
wqzQn0T5JAJz45CWOGwy15dB7ldGrG+sp0wRCNuKhVKoBtIyFUx/eFZ9bcMEtGD6
Z0+EgeYXmWLd/+Q4XwSTkNgJcIpc9+dEVVFo2tB5ck4rtLM2VZRUOienGBGvH8xW
N7qwdQAbOGPaYRAh1UAuFkltK083HdLynFgxbBaGE0ZxqBOp0B2AZYIcgZmMmbeH
r7f/vZHAh7BiYT/B0IvILIy5dHI92LAQwV7OIFTSqK3160IoTAoLZEZ59QBuxSec
vNCpmHsUrPFMVMucfQZQh2NwMqUvKhSG+nmspQ5QZTAlnLQv8lEyUbI77JNVp+D3
UbOpVvFvAWW+ajF4GB9tEkY0FCo+eZzUfGbZ2WVATMGl/JLjvuyxIkTFRtVrVolB
U8dWfdt18s0j8kgnJf65YRjGyrQuO1FuHg++bx6cgN5Uo80qx+olt8uMNqQYGY49
4PxgMQfqoz4ohGa1s/b4yFkoKDSrWU48Xx17WqiKMGSrQT9SHDb4peP4GMtfRAD4
x03BPOkO7n9tDowYo+s6C9ugCKFiC8dTpxIdeorAF6JjIxgsOH0h+bTy2CtONObM
s0WCT84fC+cmdm4RJi/xa08HC7xIe8Me5e8vFkGCrV+5l9t/8sVTDHeHfiyORs9a
FgjqIuw+ZacJodS44Qj1beCI/+kPApCXf1JJ3MhkdBWktLc0zKBYXJwIdh3cPy76
QQTfQDis9Y076gDJC0mdQcjdqqE2fsTyNpTttCZiNN5mj7lNkdPW913dtsKhTg2B
lFbg7GZ5FbJeqas7yv+jSBl1XPPJkqTMdFKo51P9Os02KpzMMBOsLs+i2fuoXjzc
M3+w4skV39Ct+WypKGhBbW/xWxM3v9wKYefLVY61vLcuxnrLhzQqYByICym5dtFN
W4qF5ywgwe9k4xg6UqWLPGHlJAUuUpg9WfyZkziwRRtS5T6ADhjo7w4QhDnXSivA
X/TMcj8/JdpYyRsm7duV8B+ow3aWrqw0PbqAyrll+c76jiUCwO4jqhXWxw0V2Xr0
VE6SHRvZNyKMA4VbXGPJiwR8Xp5Bfb1xlrmj1tN2jo/H96sQW2O8nHKdPgz5Noy5
rVFhLSDEadTrQtjO1bFNvB9qpru+btGldFc9q8R6BzZXIEayJzMKzyXjtemlRoVy
KFApej0UfCBdZsV9TUXlvEI7YtS+OE1GcmFPnx1MbdCXuQh7cCJ068TAlwGdgpZz
sxEPda1hM0iAeCRAn+YIv4TZ7gPAhGaazvKSR6EGN6q5FDU4kYUk47WfUAMkIQR/
B0m/oG84mnBwndm2cs4WG167kEsXm5WzL3ICWsVpsDnZPTvkDTlEgLm6B9wJqp/1
wapOWfm4rGRX8+kjWrxneXe268MYV4dTxKpO80lfosI7qv4ajYeqoXltWVtOGvAS
PVphjk+D+C7FRzHOdxfcs3rD0kIUWV0vwAlpq2siYxPE7Vjd68ZPjtqWMNKjrq83
DVt2HtF3y2CM9Sg0QHTpQFG6DuSvh29OJ78iSpxT0hAawE4alHclGJ/xEY0WVQVl
+sHYFciq76T0uBn1rH0I/RVvgQnL/DHPa2KR1NEpJpX3WYPDnDYoCHM0QHAagQAc
FHSU8cN/vzeIymauxtSY+MKla3n4l5CDTzRpAHQOEkVIdElB9Ue9svqccN6Mb7DY
RXErWfaiKrvMi4vIOL4f8R/WmrWAwv2b3N1sy+inzfG8jOP6MVm2GoBDjqtWHPQY
l9LPbBUEizrOObv4t8Tqf6dDN38s6gQ/y6mYVm1L5NmTnUsQfOiO1M3JiS/KM1hy
hh37hOjwEKMEwifL7XYfELoRUwYTQR1DRMypjEPa9XE1JqhcgJKM0mJNbHsIm48F
BWrNWi3L4c4BGHZpB7SGYMJs51AWjmjBfzbSOOQB7+gKpixnH6B6pcKRGyIk+ovc
bVPySe7lmutJ9iT1BqvWTt2sUuKgjR0w6qVjROYe2SI77L054gbGA/vRrOrg9bXp
i/KPd4+uK/wi5O2KiHC2/DbXLRzaETFAjSV8x70Q0QgpCU2EVqIH9mH2BgRmEXG+
83WvPUp41DXIacwd51b4i2nNX0i1ZSF6E+XJ39Dpz9GQVl78ERMjToFwgIBS1+FX
4chUQvrQeJxCzE1HzCp7Cb0PAsVXSSdwAJAchz38N2UhcJte6ShVmdr62TgEdW8C
/UQ+lO3T4MkuCzU1GxhcDm90808P0587/GrCPSpfgD0tAuoRxyWtAeC1e2VEN1oL
I0BNVTJMnzh9qZFlVDpQqCw+naNJknua0j1eqdAA7i4Sp/DtpazZhHhQbOjHTlHm
5aRQl3jpLH5M+D7NP1DC/iGvNmiI2gFXjJOxNA7R9XU3NHqMh8+WbomQX6mQgUxr
9n/u/YqjWxz7Ug2u/l6O15wUiufm2T4xZXtSKIg8S0nRsHjDNn3ynx2gBI8wC33w
TAiUOvELOtukuP4wIBWFuoUGZCl9EHpiMW2/fa48d7ilC7h6MjSX+7txAtODDKKo
+cQlY+NqSRDAusETmzAwTi03Sh8jJuS/CmowJbRcvW3aHdx81FN+9g+Jg2l3sL0a
qW1aVBJQyjpTi88G45ScvYdaCeuRoW6+a4ZnIYkmFfcHODtCvWzVPuTXHLCfOmsy
/8PP39/uu650LOW5WPXqTUBSR0XARooFwj5QrK89UY0iAnZ8jxs1d4njJDcO6Oll
1nvgFt0k6gp7nAmIAhnvQrnPMmhfxDn4wtyrS12gSpYsym8o/23psPhN5PORpIeo
8CKTy2KUInXyd5eJS7fcQr80SR1jZbNcAmbmM0iqAPHtcrmASBh61IjVeXvOygWp
2QMocdoiHhyiziU/HgIuMPNtuL4aoFko1q0hi6SeuAzf9kXW0eHK7XxmfpPtBQLk
grJX3gH7jGMxkbXCj1EJzRssSO/pqbA1kvHbH68oN7sE9slRE0CjaKFz636g/VT0
Ecm7fXq5zNGyGwtWh0n/cGhtD2s8xr8US1+EeQM6Q1I4c7ruwXGrwPlPj3U+lV7q
RJff4W8TrmbwMGCOzH4jFFqt3nBM57RBwJPFPSLPnntslmJbVbfzf/XdUKkcAI9c
NO6pxPxyMYqbUaG00yS8Y1AQR/frnYzpQvjUlr7iDMCIYYLxlHv3GIvazXtqoQ0S
YTg2mFOMx9m6iGKYMzei5b0zqYVNdxRp18cWY527je+AGUHBUolozbA5HfCVsglJ
6OcfyZpQ5cWlPtIIIE91f2x4GblkAe1fL+H8DblzGOZulqd7RrCUBUw9Q9HkAlIz
rU0dXCZ+Pagp3ol1HADNIoDF2z5DFHZiryKw/kPdNjJtTj8/Wcp1vSxR2r5c/9iF
w3DOk4wB71c5V4qS5W2cu+hgpCGtO04esPDr2nzspsf9TA9pMu0tWcz9TNCiy/r7
hJzbeUhLSjI2aiTrI8ZjmADaEEuudAQ2v5JhB0iOAp4Hbp2tZpjmRuoKhkPyvFIf
E39YF87UHmby/tnSksqh4Pti1yFzCxI45pxluCRMW0Esc0eBmstuRXvCI/qkNZG3
wsrAyaMftDlCVJOcXpCZxR02qkh9PWQs7aIgTz5wrC6cC/R+lNZIRZiywmJIEbWE
B387oMTWl4z3oyTxTB0ppgp7w5Iq3kBqpiQjTMMyCKyA/viSPKs0ATjbTCPrRtI5
5csnymSa1B9RPKjpzxJ3mBCum38iTfaEBUbfwclXiJ3s7/ZR1smruoA8xcYCN7x/
x7djnVBF9t+0d/qBE4stg73B+AbnSkf2S/2fbZRGceE7Uj9bLAdouG1tOxXyawhY
Qh4/LWLvQQcI1BBvTh5dX7H6MLxh+f3D0AexNt0y+aOGXvGS+BIsGLCP3LgHjwpJ
3eP6kNzVF+ygXvKGktA/ryNI6teyMJaHG6gsp/SZ+sNfzAyW4RCHFUD6LgUf63Cl
zS87slP/xMw2LF3WHQzH3kftD1CGaEmso08n/zV1Wu7pXx5H5+RSfpwlJOxzmwI5
CcpSUlBcqkgJYDcVpY5XwWg8tzBFd764Uh43ECkdywNWVpLBekShfg5mdwclbxiH
m+sD+Ng+j53lIiwzhJCLbFt5FJrtitfS0gIpu8pW9hE2gvOiD3Q+0BnEX+elC+df
8x0MbVBrA4TGKJjVxBUs8YhHSyDf4b2j3POWzp2av8xgDYhdkqCoT8xzXJeYTwGN
J3yDZLAKWBQJD2ca7qQY9lfZyYBScQAUDI2VK50HJrJo/3tgyhOGS8nly6lGVhOE
9ed6XKgDfq3U0RmZz8rU+YCP2U5DaVHp5ptfvRT363L5PVy06xmnKalovmx8VZ5O
qRPceeJrXMZjszKyKAYPEOxpAhGcW2NAjBtYmJNLa7gRuYVof0TxSUzX6pKqscVZ
U1Jp82Ruu2N+oQcc8fjSbJIKCGbaCcctbm3njsJCAjFV33S6Xzvpu+7+vuOpXWv4
Dz4RWf7RLBnknrRBfsfQ6I6+FONrs+PLNTU8LE8v6f8inHmVmTN22/R0btBobQg7
yVo9fGrbkqtWST9C53BaD9Ug103QhxueVD7TiAO3owGszJDF2tRUJarjsjwV9Vku
YcA91/d1n99iE2sypbOp9v9pNfCIKMYpKOCOnOMR/zr9/ylLMDoU7DsPbK0lBkso
R2e8VELm89E5j5BlJvenH7bzJlBbuehnI9hudEIOrRwLd7TszgAU9Yj35QV4RqEF
5DsaKNQFgGCoSQZ3CnRl/7bWIwzQLbULdZHjQbXXpcsLPh8Q+uNOBiUwQBWLWzm/
8RFgVG+HyHDX61ckh45EjVe4+Jj6YNxojDliFZbEU9nwCzolQPUM2n2p09a/LZ38
Tl1IN4FLy4nvHVEC9VfnWTKwTpdocEsWGbLUpM9ZIs4tLV8++bBT3GjHUrQxtjPT
LnRili2LOZI9CoAx7g/vUocU9UxvgEHjEZMgBd6Lu4G23WR+FWH6r3B+zzI/sRSN
NIDVyyXJD4Hh0yQKqQUVHkkJqv7328iHQRMQ7HuQ79O2AFbn2B7hWZVjEcGx2cf6
lav4r372XHDMXijDXCxOXMeQ9+IvN2nP/jGNXQdkv2nVp4PUdgdRquiM2ziYi5kk
O6Q2Ugso5gPVPPxUHFL/KknzA1J08WOCDTG+qDwJdFysjbuQQlMaItdpxmHKifr4
dc3c+N3rcJuJmC7j+zbUNoRNnAacVk0tOTv7cGdmpmz5J8T+GB7gZOjtnPVGfDAg
Qd1HFuClG6KD+R6m/1YyHdEKj3CdJikhqVTRs/EvZSZ/+Zise3Ydflg6ZkgLTu8I
zxoUd7r3FapxkkG+h8wVjmBBf+WQfux3ASklGKtyn0CN9xuqFbZRH1aO+7Thgu2C
2LIYcHYJALnY3oBMr3jgdeBMaMezcjuPOewc3+Gix0L2UuqBXs9XkIauaQhLiwJz
veHgvFAnxt7iGhg6tayhn7/3W+KnQBzxq6wIpJJAIRgTYcnhtgUNufhGqaJeru6/
bQIc7P1gyoA0QfA2pMEOUT5Krz3PxKdao2pTXnJKUIcXhqPUS8UCnHoyzBs6yUrG
ScYM6Msy9S+/+asoiEla7L88aRuY3aGml5AWynpFNlPgtLll2W8lkHyWhOIiEKCw
euCdjpOzRD7GledfD9OzZX1rz4Kcr56D6H+SY2xikjOjQOM0d0dxcGHfm3UryU2Z
yPzSLlLsGeG6r7Eb9U+JJOmoZXHJGe0pX97u+hoREGG4rnMNh4sKrVf3VLvLoBzC
IjxFTXukCUUFjxH0iYeNE49gUV5lNJmzI5mfoKsiX8kTjvlbipB8xGgF32THlqan
lnPz87FUlr6bxnIeZ/c58kz+3xFeLdWCVZJaBoluaMJbvm63q9z178erzAg8PdYI
uPa4x6aAtIvHFe9IVw+Ka1OBS8tBmbF/M0L4ZXnX10qf+Gc41sIO3bjyNLfahoAc
h6k75OIYcxx62Nt3ei9WmFV+HQHK7GIoI787Y/jdTYDvrVB3zv36jn30RZkRkrhb
BHhxtMNR67E4z8obGXW4h0IGhNtC2eLtVPPl5zppg5xNKhgo+PcvGFYLyKSiI4YG
ZTThWxkTI4WgQIAiZLZ1+8izej4ma8OANTKHINQh8EfyX59CFfryyulDXqSVJSXt
JpSyTrbjVp38Dhxzxq5p5ANppdhiam0uh9ArG2fudhnXL818+XMC9kAzFTxxUjkl
eNIZ8s/JtEGFw/PGdFr6c0MZ0+qv2xE5/VoHdregxNsmF7r1d0B0H7PlkHhmxvUk
So2yuaeNDX6kdQWv0X49HxNro6y6nc1xE6QosWVG0szL3R70fylvLSX0zw3Gjh2f
jpcWoogcZfTQC9XnKU6xHPMJ0DAo5feu01nidmZETmgdzt6dDCkIYmJteLFM6U54
wwp9yojT17lGTt7zmErY9LbxyJsujmmDn+C6f1XhielCty7A+SBRkCZNWGrBrsUf
74xhsBFEgL5u3ihxKWShPrlw5XyNfjKhxNZDvzVP1imxj7BFlV58MiPtp6f3HWlV
fGUMpWTXp5wxceI/4z5iRxpy86I3ALJvRDH25+py7RxJzXCwNPnkXMBij/5v5b56
z4fN+tI/jIe3xeFfizxgAJHmZrV5+Y6K7Zx/8N0LI2X+oKWuq+t98SYNPXUr5Drf
RsaGU9DbqXP209W/oH3SM+gkSKId/BO8mIbsWwIs034QXxi8bjXWklK5uyXnzfJU
rWeKlWv0fjM7RH81CSWG3iYv+LCrvHsKE9M/hfKaRhepPopmkIFWMt/66F40n9Qt
SimmprccotZ16bGWAwb6QBwP6kynY/hqxFG/Y+eO/QS+98FKg3lpLGofHDnMzKXt
v8O9iJ422IuTN/ErPyMXTnvR2q1AGX0IYkUTG8tNPnAQ3eChsVrxtF9ldlMmVwu7
ysOwgEO8xviAgojXy+we9zDIIJAeOq4o+5GGEAN56+vaBEnIC6e4TppUlZ6kvWfz
bUWoHktIG/3FSwstDUIJUcXmpdWd8/H9gHBtDAFQ7PEak9eglHy2PuWm/BDM2Jl3
9YpenMrawaI7XDZ3F5PwHjOwnVFRlaL/DdKLGQkb2oQr5hcuiCzd2OyIX7/TDTM2
NDnsYZfNaeZvqQxMtdu7F2HWVOFoqzTL74W6nJ4l9txFeRXuL2yg1nxKfhIkTzM6
5BzAWkx9h/0Rv3C0q7MwCTy/Kzc0Cc2OpdQkh+FCqUiZv2eavJJ94OGnYon6DF5p
ZBeSpw6JF9nDh+9d2qnxH4Gx00EYphlvVuMosIPb1HndVzZZmFdpDe1erH0XeybH
ucBOfWzF0UFB7zKuwWHOO0YiGJWnOryLFZilusW+PdgEl+O1e3yvGFACeNFmcgu0
XIp/wvcg8MKGoRWG14uppsrdJ+jKbHHuxptsXRIc6lsLvKsW8+xu0LnC/oh9nzqu
yacH2KN6UQxF/5bsFFsucqxr6whXMZP6yYirwSpbUS2XE17Khhf6+bWxtKJt7jgF
+LYxBLCiPN1sd4bPbT6BhKWpKvu0zfZTOeHLScnwJB2MbpGZFZ/nzy0wJltD4ggm
ZyCN0ZIWJcIXklHXZkVgJtr5BjC0G2LQBOBNkLcwiZcqjcuoIbZ0XMtk2WnGgcan
3D3J9Ar6BX3172WBnKZ0diQ6ANOnxSePrdpl9WCSSQGkvsvzxcrJO5bH5ChK8P9t
76olbsh6g2HP1s/nuQZRBdg9N4cxRyG+EYGziKCVO3hXYuyMtpF26kHz5HzVPspq
k6yhj9LBmtneVfJxGgKtylN6Af6XjO2m2nv6TO5Lbzu+ZGtaLdsydrzZtltXbHP2
39J930chf0ZuTy3P+WT+1vtkDkNuS2XqikoJ0ZndVL/EHFvJKRLLP/JlRWLMhhVH
NgqHdslgSmJKVBDX4NfwPpwyVJ2Tbu0IdMuMHBTwzFTgd7/B+FVVblmiyaUdjnFO
VuSGKb0lcCi1dkU2IDQOZiMUgmGASwI2ywmuVMdi/Ag8UGqejaDQtauxxcgYxfte
x7NSgdCu1he01xkYLqKMh6oqFvEcauPwbXViZaoC+brxcQ0R9YVbjDKX1Lzj6u0M
yNyLuCYElKjITqUGz5YtHRiCex75Dq4NQpTmT47s2kZwQKXOFTOcu96wg+WiQg+/
NAfoFewQ+Gf1eiT8O2TVXExDMhxOlbVrizy/ZI4laOEzyOYgHEzC61/aGXqGGmSN
baYZc/mhQHuxWYRqotKZCC2RQ0h3vNFAkYZvb7eI7N/Z3DW+Un50QwTiRWg2tPiy
ewBxDGmqapaVMbXnTOX4LjtaSE/Siq0XTybEgojqTAGurNkUqoANwUetQ1aCtlGz
p1yjjz+L66H+cOOleKkgEJMD0NmDT2+V68Ti7TchxO2Aej2XmNlUn0THEmt/3DGD
NVJllzq7c688uj22rpvuobsD6ULyMyZXZN/fpuW30otCH3j8XaLVOyz/qypejQbu
2ySNXWAxKF+o9gjN2UVhAuK7cpU9kO9It0XoOZJJgNV+/q6j38kPx7+1Evyro3NZ
iwsYeU5PDa6FmudntFZrL+B0vHsjZbA0VOlRwA/9O7CGg1q3G8t1/mMIriJ+O+1j
Yw5HZwbargwYgf93H16o1yRUaNEWR3QLldmaBQpdSdG19CgRfo5nobsbms6g2H5H
5PWcExEbyoEThzfAPtwxsnyqQnItYBwI09+X3MX/FMXlue4EifHAJMLYczRjgxI9
yzWK9pWw57hgF+rsSpDibln5LeUvrzqS5TW1D2OAp/z7UEN62cSoeSG1y4+DWJpu
6ElHOCWn83kv8A0uqXuNkDLa+BMVpryPjQgjrAJr1YMUFA3ETp7Q1AiSpjElC+MG
5E10aO9hHDy8m6tTxEsju0W2ZOfdQxlvMsorM2kR9HoeUGYBP7s6GI2r3nav6SNG
k0pahrh7+7pMb0zZcOXLm/kPcOo5tDLB4EFG1ezOLiMn31XeOta1yqJQjePDfWb2
ZK8j6wAg/XuURsnbSbmJV6uFOHY4wVMEhKA46xnDaX751I20Afh7s00+3m8e1hy+
qbTk79R4Yth8R5/UcpRiMonCzD5t9DIIwBmJUsiDYQqqfdvVrGeoAdMBptdIzauZ
Ks6nepaQ6ryJUNK6DXN1/G24i8EYJTX07Xwj6443DSUrzIiTajhcoQ971igENa9K
PCSU2WuVOKERuoq9SiF71Y88gCrmQ+xgzTFsaHOEI6xrLeZqUpKnimjH1dfeDxA+
DvPAlVf6SAHXG1RtOlb2wlgnVWYGMHLRt4Wn4qDgeXSLZc/c3YlSW/GMELyX7wd8
S3tckR/SUsCgCQugDu2SspdAifYRfXgxSG6WQD4IDSjWU43GZHj/6YgVzy4rVq71
0ePwyeRpgDnAF1s0c8RFKWnfvASgYg+bC4A6mzw6kkYRQnEkDRO84xgYsyX6kGdQ
myJyI8mFaYE2XhNzIaS2iKqwnyCaqun4TVOH0X+brnWpbHMDSifniuhhaZVEWDfm
ivyRMTMY8yAgrfxN2oDAO7v24TJnms+8Xf+rSIJ8k8kX1N0C+ZU8Rap6ci20SQ/Y
aGFQO3+av01rjgiTkGZA7dlTz4XfM2PTN/C9tIKE7SZA2odQQCb/mDAQkywSJR5T
sACINKKv+uHqggLnJpAO4ps3Ikabv5pR4DLGriK0wzup8fvJ+GZl84IpFaF20k82
1zG5qqae6UIRcbohUCPnXxs4v65V8k2YJg9Id+hK/vj2elYlHS3DvLtoX70yfGFC
Ub2p5NfJ0TI6QYPaQjEaB1LU5sc0+MymHBdvg2AwUTcwLCvOjnEKx16hokiTu/a7
3SrIAQxEXfiVmXzORx+O+p6ZMaVPsu8J1LPCGUddEvgOVQnxrSYZcGK9TFr8z64x
LfA7fQbRjL9HK6v3azvNmZD6USf1C76FDEMdB+nzyDHMeZThM40CHKD63n/4QJ89
Y5KXsar1Jk+4ftuXvlnmKkQ265VFg7tQkjaNiFDdEw0XP0mS/CdoLG6s2xhzqdDn
ksSRYr5+Qw4306vk5A071S5MpFXaBaLowi12Clq9nDayvchkT8/2n39tK71+AAJ/
20SxOGpombUtnulFETa8q533dSUt6UPzueD526W5vPD0lu94JPHJMLFW6MFkDFQB
SFBtrWWO3tlpgMqqeDjwVoDghCQXuPqR5bQOKGky73d1RRUj6iH2LAzqT7HbXW50
JNH8OtXTrXddbBbDM89sUql/h4p5/Ps+i74n+5nVSIaVYDqugWUM1MOognEUkHE5
st42fhNPvObLZLs4egTzgPACPzFRfKPl/TWaAZSXHN0rEYlS5/OBeNTqOQb/dZMV
BP0RugHK3mV8s8NS3IgspxYkAttPNsuhPYgf/YjwUBx+vfuJ6jX/bx4pJ/MQ5Pd+
eMqXd2DtAoKxTrAjgfnuTRAa1e5YPV+Qh88ChH8hRJv7sN5IyWeRgxrlOI0Pe+nS
a5p1aHi2D/RrvA/OveUnAzZb9Uk//iDsTdJszBy4NIBMOyL84HzHEd3StIVn2CVD
IfNPNRmFs+msWaUIkf0p9LM5SXwxyLr+Dc+4y1tFColou70BvW4k0tfOYDVckx/Y
U6DTnF+2g9NC2qK/miT5ekoVdnVQqbpD1fP+okTsQl+WRrN9ZBbIfD+YCJeLRdCd
sv6w/zG4QqqSqyDYiBdobV5siZVZmBZYl6GwPDiq72zJsnQ+D1zOwCS2qK2p/Ogq
nLwrjEv4BfYVXjDLbcx9sWIVWls3vNxlRjWI4HhKd8ZngNWgC4IQ950PaKX1yKf/
SjJlA4EPv5i1Ap6pvsJgdZZZCCusbatKb70oy8p4+B2Es7oZVtw6CEjNfxmxQ/ZC
0jOcfW5soyz0+1OSrXrc11QoLwc1urspFVgwIxAqkpWJZjC1YxZIg7xhX9wB+D9L
V8hLMqJ4Lqgx7MKY9rZr6+SwqYKx5kQBn8o+Zq3JGSlpEpLk/qnKZKCBA6YJKF23
zRbQ17rFQt9AmTF1fjp97PfquL9XmAgjgByNGr0dUmUZxuusTeZPmsSYhyAeLHpa
duXK75ykFyuQvhUP4Ei8rbCQIPdzOLK/OgL8U+XyYxlsu97Vr82ub9BZnnY712KO
hIbTHLpwmj937DK7ozw/e3N4H83JoHEAp7BlhlXkLy9doSfnanAOiJq3RRRx+u5R
G9AVqyE0bjBXKbzp7xXRFLZMsbaQTYDm30Ailr0/Rjxy/DfSVC/CiFOuVkhRSnqW
oXl3U+grpm72E5I+4lPcUI77E5G5KdXrwAQqaxYUwvjXurjJbfk48oV4iGs2C85M
+0cL19XHfFeBzh9Caur+yBl4Jnsrz9RKZHzmmWwgpdXh/o7yvcjQzcSiZOnSVzP+
HPDuKbT7SbG5H9DmXMnzKIQmtHYVNriEYO0E/v83Wo6pMUkxV3vH9Vxfkzpd0cPl
5tSYT/KA9bCy7Km8fj56ZfJKiReD2wxe1AjwPDb/Jaa6gKsSmZYV68og0nQ5V9wJ
gemg3czDygNqXx0hwvKBEPNXmKGatVDMtG1pbTrP4zjqaRSJUu5T23muivDDVNGW
TPCUjHFoR0VtbcdOihwNzEBGt0NBGUwOO8+ak+svDr4gl+V/tPyRwVT4sEPJ1xcr
xSM1x8eNabrAVttREw+P4YA5NsfQhOXFmKg5aXuYeuUeTKs5HvHubB3EPcBBVomg
YpHry8bAGydI16hpH6pihXBjWvQLSj717CtrqcQncnd8CwgHqtBTYklrrzKHVxKA
V5i4cbXMXt/Txbj6m1Mx+CbA23MB5Vp6mOotLMM26UftmmD/tYdNvWg3B5kZOVUn
pAwwBW+YYK/zl9aFR0RdUSS/AylHgAZN97siL1rar8ezMfXa/3lj0lMvvmQTBxuy
ugL3jggXCUfLAyIVYCDxcznVpwCfOVpoVUXkOPCLERP2x1KCHhFrnkWz66Jtwdsu
Z1cH4bqmCpLcu51o7vERhXDPI7UbB4qK+rR4JeG3S8UwBXijyD6O9F6sq3F28ROq
pL/nmf3DeWKAl7ImU3ff669Czwi1RZFAsAYbNls5x9IIgREQvlVEwxZb2Klq0AQA
JKAkssK5duoNyQiStitIRQ85IEriQQpNESccArh9kNelYVAjTOif3oGTPPXSVvmn
8qCD3qrK5/Qh31GvvZAx4LqXgBTv4ONHoz3UgzLUD6Rrl+rf7t/oE3IzXOI8CUCg
Qx0vboziSDZLTG2LaEzONHUVqX8uloWDyregPWyGcW7Dwz4jRzYlg4UYKPbItue+
9HG240fAHYdk3QB/2knYMhNt61pbTFOOI25SrJLIn34lSz9uWuFQAeAOXVOGBztj
rGhczhtn5cKAkdDdXTPXaChgWVJvTEspS7+x+xthW+jjgN1hhXF56I8wbRVEtziU
Oih0xSe/QUKb97ybrc5r+jWW2UVUmn+8SK0QYP+haDMSo2OzGItz9jQwIxD2mNjz
37QvM6lyuMz9SHZYfS6RCtB6Q1GXz0XXRjcdBPOZTHMaO1ykrTyB4aOyd9OJLOB+
yBBwQnY1Kc/YAVZSxh/Sa5Ug7nS1Xno+4DE9uM/kAscV1QaN8Q4F8hzvmEeRqzz1
ifcye4zoV7W3C2GL7lLmC49RjSvI6DveNBhYtGXJMM2bHiYpIVLW5qpkiBRamr91
/wlaFzqvf7IxHYqyW5fkrU3KrAgpNvYNXJcbSb0q7tY+CeH716wTF3lVz3OHgqTa
GTbNB7SCAXG+1Q/SMSexL53gRPMZypFR0HKjjRF4QWWSKPocWXZZMSBmjQ/Y59U3
PuASxWVG1NzPEmAurm4dCzDIKdyLzCDwop16EYFOEMNlJQbmV0JO+cEz/C5X2BoJ
FrdNVGEMGuSYyp/cDeUt582c1j8KihpK7HEgIqkgYJ775aXMQvRVpY8tiq6kYnLK
p54oOvASsUQNRbunGCSI7LsoQgN4AoFYX/FYpsZRk9S9lawHOIKBw4qTgW8O/sMS
V2RtB8K5+3/WhGmLdjcrvtv93g8nRRdtKNZbtfx/Z6mwylwA1MuavpYlrTEmpyHz
Z4xg1EBrK5yzxcGU0Gg2dpc/UbA5YnzZKBXwl4DdSq1AosMTvJuUL8bLI43xYAPX
E8M0QaX6w22OzIqFyradGCfw1v/ZLBQJiJ9oD3o8JlQH5NYW8UvvoKOAef3NJ4hN
EnAt6rd0z+R7xbwzg3lrds0pHB8bmFOCSaNH1AvqO6pBb1yNvd13oSPufWw8pkoK
mqgkxPnYkjI/kB/Wy09TogsPpRG6nFQ6q+HmY4740tKsWloF0hBbHHCf+z0BhXsj
mHvocvthm+Wk4dEGqTlODF/jMtP1IVWaC0QiRZgunupWBsFC0RNjTUDtx2BQgRFG
qdWes9b5M6IIczAJJrUvW8sVgoEtrkbWy4AlziLz51QRObRjnzbqzOHW+1jijq5C
QvIr5+xNCrlgCw9QVLOLhupBmpy8gSxhg/Azlt48ibXFkmZ2fqPniiT8ob4MYBLT
T1ki50VryIGZW6SD2Hw/7uLKe9o2Y5KsUVL1RLE/3YXL0r6KD/hmm42Jw79+25ce
YVVxBQIcejRDSlwmfuP1gj8aUsai4M7v76w2UI9SAnYr7/zVDgkq9rgNjh8d1qX+
tOh2YTBPNZEAv9UOTCYxcLt3JRi3ndz82lsn4qUF6bfcl8wOwMI3MHzow8M/eO36
EjWfPPbpV/3qsB0tzmPr1rdKjN7SE5RNZHmt89V7CJL/4YdkrtumfH2gukThzzTk
0byV7ssaM/W1sevxE9sd8CQ3aitySujyCfkaLFykxkhwBwaBtmCkqE283S6yPuiZ
hsbT+TqohVeZnCWiTYhqo0fsqHY5VAPqgOcB9JIWYGipAble2PWGcaKdX7DsUv/X
+0JCsr1cBS1zzfPn0gtfljbFfX6TB9Tlx2Q18FYKgL3zYVNLtPSrr/l8j3x6OGz7
3o+BkqUX2/4EFWAspfMvuJq/m7kDjPN2nFeN2lB4a3OcASs3r5oOvJ7o1bTstmkS
leBXYlryhZePECBDb+lDDSzhucPD8ijlcqauBZB0eyi6f7kEDT/7SCYAUCo0slsk
Zu6AP6DE3i2imGlNz47KFWIieBwNbwpWU/xKxRzrOjvCSFXlHRa3uGf1XJeZPzol
xPk+VG5iAX1e0mGuykUhuDvug1Ahi0RPQDM6ag9y6zdGrD2dykExIZOUuc3PTY2r
sTcliL+wzhHP2gAzFSx10Cj7xS+5DXoMu4fEQwO/4lCADZZ9+CUPnlCsx9BMwtjd
W2qiUftbcdXX1DKB/sxEfvKEU1YwVpYNLEMiqbb47WLSYxkX1hmxX24dPDaTbOIV
WGTLTylxR7nFXR7TJxWdIU6n2iLMwW9wnkrayAGmPpgSZlcAYf+BQnA+miJ0WzjA
3hsA1MCdGltlFbP4bfA6Pmhai2Vohxoo9/ZHrkYnujGl60BUzakcyJjjsetn0+fk
P8Sonev52XPxjgLerudM2w2Ckkl/dVzpZ4O+wtQsIIY5buvkzee+xI5+yzVUKYgw
/h6yVPa27bKRHBmhWGagTTHQMvH7TmmGYk41A53LscFisSiabQL5Y4jmUiZcZ6Gj
4bFyINY31HV67Ek9NRt6+UvdsAiy6Bc1ft/zv4vdVAW+wNmvvZowGqhlMhweweLf
dBH+WmZFziMo8BUHV9EIpwiMxEsFPqnb8PdrwiCs9Qw3GKcgxU5WyVkadfeWNT0V
JMD64Hax4lyXYq/npioZS3nq3ewWyxpMj7DO8J8zHEq2wDES4Dca4q2WOWXrSdyr
Mzf+FlaamtOfmuDn2npqg/fckmeO3gF80agvGCuIJlN/OkIDfwtual6OmmIybxkP
59ktrxyyYPAi8UZI7Z69xhHXOgNwGYgC9ILzHjQOtoKE3dK3jwLz/IvB1nXoEy7p
QzBkL7WNcFdBgHZCZsEBNzHSF+HxSAPGEfi/aNfKV6Yihs4B0K0BEfV+ChkTq9y6
N1XFf14B7BKFuq8Viy/6PRxMZy1xi1uNI5G/Y0aihBDoD0ho/SDKfBDjFZMe9G9g
FAmETzpxg6yDqZu+nv3FprZKklScNwAARm6iGinnUfUKnKTecL2ACFiqc3KylpcB
2CTLM5tVxodNAmJu3kqScxybktn1LrifL1uOQlG9kw5iPwXF1HGxXO5NSIlkfsAv
P7dS6bvjp38j0BdudcVXLixEmqTUG5Hflah2G3Ap5yDt82LVTpRVysI2frfX7S/c
2L+WBpaV9+tM9K8R219KQnFcvYK9UM500uw8B/5RGzo+Bzr5Fu+jc93B8PXoE6XX
4LZo0Qok1OML00Ff6c9z99jeXHHGYeYPZy7ROJgPKrPvPOrKPqHpIslJ3o+u5tWl
qi1nIxyHpt8E5a8mzBk+x/74WslDgfB5bi9Z+FRQvFqTxn4Vi2+pLCYg31slH8np
9ufLpnP9kg0T5O8JJWVvQhtYtga2ZBfJJmasE3sF17iWb83AA0TciM/YQmXWthi+
rBd8HXG5my0uYwgjQ0wFDsNtBQdf0qw4DgGdL7+lkhdBd/LIiyJBNwGrZbfY9TSJ
FBNFiltOcGHQH/x8dYhKLxWNZUfdwqJ0MpyXVmqa54+i5TDv0iq+srYscNrRw80W
iwRSvLtehP5NsgEAxjHG8Iltf4opByDFNB4zJtii4mjsHcSpD3c1DV8aq43DeL3r
l0iIYN7iCpWMRAQgOUM6UHob6CL9CkutItz7iSV+wkwi1AyawQCzVUPbg1GqdErJ
P1sE3m+kFRXXPAEmPgf5mGp/KJL8bn8u/C6p0CmfsKhFtb+ZzcawO+tEWA0VJtLG
WcsU5WrWEvHrEgbvhBJilwJlXaoIUh/pBW/JBYFg2d5fgYd4fhk4GnLGq42JYBT0
hLb/atgpK0AJ8ZQ1PpP8ne9M/VD/LjIWuTS4XiDnv4HKQa2ltJFnYI56R4OaCQqU
DdPgV9x5/eSE67kkpUfJSwy4x3Ba5l7826E+jGQyW39aYFlDajDowPUbygCq4wNY
RjTV1SYu/2hoSBFIznmulJa9qlsGRKC33XCyOntDwWRiCX8xg0eAgce3ZYkvq3HE
lwKxfE++yLfnYOVYBk+/M7+ZrxweZirzW9HNLNDUFYlMNKPu8FXKZXqm/PUMuCof
yXXhzfWOtIsE1MThmv9nnfJ46287pzv50z8co1wnS6mQwGJsfJOkpK67ZPg9pknZ
iLK6x5lPCVJBERmi9yoihbgjmwkOVnGuQPXWdZyTkJzTrODAXAnCv5XcPDbvV6dO
5wv2KPC6MFVKOVmK+p84ImHZFF8SaD5ZfTKQO9RhCqs0DoVdAK30vJwa5U6vrnAD
CiMHXTRq0wlRxshpaRRtKepug2bdJDbWxAF8TIapWrpIBHsHVMkGK1pDjfCB8a+a
oS8dSD6W0fsF07gpSAaT6RnjU62TkoF31vl9wOE4aBo4L0S08Sj5z0q+PgzvG2m+
/vB4aK+cXOn77WYAmItvGNG9I1f0yGIKj0CLM3H9IvoMPsothzCLYc+qL+Q0ryQu
9CPe9iuQIvHDEx/w3ctNVyusGHx7RzsEjY55pZORUdDca/LTHp0oFHYBTimOBXlD
N+/GFR701cA6gWfgSGKLPlQsFALAcyZPBHDNc2cAqESJ2dxaYpUi/l/kr/IIcRx1
YCibtXIZXVz0E9sJmhIufVrdtY1CEnLPUCtKFdsqMZjPo4hcPoHq8bylyOQIRtLU
T8dUnlFxQFozqODrPY8yDaBxma2WAEjGx9GmojOp6ujqqwVbTs11cQs9NVzVvFY8
P01464UnR6VTRhc/YQG0SOQQCocHPKnh7xIH0x6chHz+5Mk5vCHL7ETWK0EcbP3M
Ko7pT8j0jYJXe41KMsV7NkQDSPF5NeW6A0OFtiqrTMtAIgxFEWeOJuOQuIh5NEYm
cAaGH5Y7GMa1VpCp824M9fofDQYCRO+rdhfquZvvxC4Hc0V7qdNAK2vljmxO24tM
8Z/fnjyF2x4VVY59bYsbbvBPJewKIZ/CkjBZQB0zAHgBK5FpHVKguFmcohN5Y7JL
wzB1hGQMiVtPHg8yv8JFTP7SXKSnMyqezdlxIkcNbosJlknT2O87XzdIi9hkhmR6
81fNQHE5Ga9kCu52fIIIdNQ/UkNOJ0qVqFgv8l2tL+L5oEb5rnHiVknsUqfep2H0
9iGeEm8EKASXtrO1gsZJ5HluQe+K9chYH+OgrHTI9L74CQUcKYdqp+vpRgkJtbfF
k9xHy4u1VOjulWC6d6GVyujTWAwOMCbsWJ/mLErg1f/Y+2K4l9tqOS6t5E3qsigS
E0DtN/H4AQGo1izI/5yac0/xb5s6RhPIjPwQbNSbxg3rCX0sK/dnZgTHhXQTP0jS
TpI53BkQ7Lxu18t0DKuy4kOQHIq71spP9GGraVRYmMmtXHKtjEMWrLJ+rQP7LEMA
xwzWENQP5EQodKnE0Tb2z3DyCaL3xL/TORD0XhXKDonzAM3A9IQsARh9qcIZcG5J
OZ6DN3CrtX4+vay9Zagi2FT+k/6Lq+i9eKLWaQTmpIjRhNE6wgXJxs95Sh5jaAM0
y+0lJ4gJdvJTUJG55yiaRZCoE0PNfaJyidqQ/QcbPkTHfq/DcV2izSeGa3MadiZH
mYI8q0rtN3EzXBn3NbhcphhmmPzOqDekMGmDMllX9Hn7yPtibGD0I7lJdTIsUl8f
8KbZE4008cEvL7v2UwvDaclVRr7IHkgIRpONdbtLuipcOZi1l7CFK146hXF2wp1q
C8JYScJcfazI7hVwMl3u64FBudzBLkhMGFalQdXWFBb6QlPoqXWVFSCpVIBH3oZ7
qoALyTqrjbVVZ6b409MYGtLTrL5We7PmU/Q8zzY8b6DxzzyDyRuD4vxn2pB6Jr8/
KS9w8f7BrT1mBqyAt5uwfMHasXp2TjaMtynCir/xea14sqXqg4GA0Bbyki/z02Tm
05r/yZnzrTj9pEU+1FESc+dxqaLrhuN3QWbPUiXDpiGXnR+lAaNW6yhCcMBeF8Jw
pWunu+xgW3iqxjzjH9zq/r47cDfhhjSUlXeQUwX6FQ8x2lvZbitRqFBohAR90CLv
OHMyo+WkebJUeWazJ6ZahiAg9JFMxPRavUarpFM+27Y3/4wPtlaHzneNHJhvYmaq
dkwscxdEsKRrSRgondF9SY/DmaW5F+WWdqQ00gN3FEdoStUucgmXbNgZFDiKlgK3
TrH6Gz8VKYTlhPd0KQIgJ4WSwy+k3YS7HzwEgzxWPXXqm1LBehUnOWHmtc9eKkdb
sqqaPw9AEl7jKyOBCrVf4spp+Bfgw8+BVTODQeSe54oifZnLc898/Ah6k5GItsre
v/XaRlMzCB9se5PebfJ2z4lmDbiJtaSG7V/iu09Vjn3AOCoOVfSMoFnq+3FrC5ht
YJSG+buo1xmt00wLf81yh0/NPxQwq2ocVfz+Q6Su2ESTX+YBc2UOZDf4twqOWymn
wX2XxUjEegiEe8VyXQnecfQL5Sy5Z4RMDhPVuqDLH8voD8ZpqIH4jZWv4mfKgqFE
2g6uq49lqVVYSIFA/HkfG7enXoiMKNwtIyQUVtV4iemiKcMWDlZqzmv85FHs4Agb
LJJMa+A2XhQrfMR2TotWYsH/4QggJZlg1EgbCVbMZavjhkq67KsHmGqq9P5+d1BP
3UU0ajTNc1E3S8qGjGZpjItfJOEU4ZPPTvOPS8UGDt1SeicVqnBrqKMfm0+s7UPu
w+965gy6ieckufDvJbQbsD95jFhmpaGVqyPtTt02fTuIEf09+T26uuIHOVNlm8SZ
lzXj0t5NuU0I4/BiCQCWKKQOxE4CFHoT1gGa+07bHW6CNAJhYbO3pS2bx9gaWt00
KAa6JkHcJ6vHJgbeLqWTbhHoPqYwC+DI1SwY9BmdwukNU8+/vtOep9e6Bq222SAM
WQluaJsXNGq+NvjK+h7Fv43I1jYs8Kkqqowr9FUkf8trTxUV7pGcl7zUNcBBzxvr
ZVMsP2I6XGBQ1JW3fj0qkJafBS4RvMFaZABPdeSVFPhIWOMdLiXjCk7mGoC+UYJX
rXL9xfidQgBor6t1o/fDbitVH7sIokOGcZWsj87G4Y8RIybvF+o9S4ZV97pQWCQk
ZnXt0jfXEaluD5TUSyngeIl26hLmT+yDvcimhf1lb/K5SgHDI23aTS5YK3JS4F+D
RsaW8Bxk1TJ+nkJ4/rG8Pcc1eSlTL6iABfUqsU3l8iumFvCxi8wNmcWGlIvEE6WS
5ua0XTTo0HWPFJrf6bnU0p9ltGdKVZpK1GaR80DpOxQ/2GIJ0282sBUDjVD5yyH3
S0lCIeSJ6S26MD0ITQhkIugW16t36KTIj6pBd/OvjSibZo8LMq1oDMxiNTopXlkn
Q8Hy8zyCcSdOZJkHl2wMK0wpKbsuBj8BaJ/Ka1Ca7YT9AxDBPiwG/LnrQMRBA0Lr
ygSKrjqsXuWGmcQL9YKFvEyepIxsXzQbINY55I2aYVH60IqWx6GrKb0rj6WDEdUh
B/FkMce4ky1cFujL8i+xr8JeNJZ2WtaMkU2C1LNVdYaxyew+qUOk0h4sqb0/aX+s
6vacZflr3rjZfaIHF9Sy1a940pxslg3mbnwbkQmQtpudrLNndB2CLUaRXYS5JzC+
0WfymR5rhRooV+ZGt78LbX53qS1xKEsrMPYnE1jzOhdh5YV6BmcvVIqb6D5aPDYw
e6zhfoNF1oZ5WBJegQEFs7Q8BNM0pvYUpgCvGHGN2R3gIxBbnX2lDdnaRPxk6FXj
ThyVggiTDMqLhEjnNEf5ig5YDCEs0Wsf4CVpSXzfo0pmnx54h5Dmrkg/5i7O4n+V
dnSaZCS07q7aOuVLzPOV1iWFfeE3JTo/1EWXWdTaIoU/4FUaBzAbavEzZiJFN3wk
vnWf3Gou3Y1f8MM4rjS90W8UpuYd6lId4dlFEAUIbX3XNurOjb5/h/T+1TRucX8Q
KRRP3zJ2oOakuRVFcDObUF97mVCgvVPB4zRdMGcba86hOcYZthYCwsMecyNPa+iU
ncXEEBv9Sw5biPvLK62SWqtjzbdiNNVzvll1m9ZkKJiGVOLuVWn5SK07EMkPFxNP
G5yqlpxEzI5yVOxzSVHXM8uzXLYhlbkRnfBqOBHZyV75kMUVknPJg9oLRV2XFJpP
7x0DcPbGUA8FhxcUT+FPdIgJxJ5yazJdAL0XvZRD0osAvaoq9J1i/tgb5BWgKCwr
cZ8ZvfmGQJdI4FMZ4TxpwjeId1+8xVcPpCBmajd3nzRAmO07dRhffYs0NifHLWXu
BJEx/fOrM7Y5Vwd3SBvXQ9oqsaoed4g1GCP30dHidI8Ga36R/wUMUe+FtcLcRjSg
3YvpiAR8j2j5N0rmXmZBoj9sXrcJcdrfSw9fMNT8No7EGHm4fqGGVcEb+wNMd04D
b0uL+2DsMPJAYcR0kdY3YEa7AEU7vDqfzi+WJaYaAD0MZzivNHqenp2rqMJv5P78
kY987t8hVc+gnSc3BBcz3BtPngUJhanL++0Yyb/ZiHbRrfOD3qPGjyXL4Nj3cJdC
tWjMbODVMw9pX78gYJuGMKy3gMDY/B19KXpDRyoGhFK2KrXG/CSnkpNqiU95BZTk
ZxIGkguxws2G1OVYHxUNGnQ513CzbOnlyOytfLPRGlqvtTFwfUPIt7F9gUv50Mot
ntU84nWUjyhGjtTrKxD5t1OYWqrnFy1rGvGCyRkXzIe5x9eWB+t4RBg2xYRAiOOW
bB0fyZ051pvZfpaJ1xkbmsf0RNhq3/iXxAwob85P4kwC2zPW5CMHbYW0gfWihrSV
jSAz/8WOteIdPWamJ1L+VPMO96PJCefkkkFLvu2VSbWUPY7SpR/839g2XL3UwXn7
7fKzqpew5Jeh6FnzFzgHSRUsQXSXFNbOqVDrd73AnxNmnA7SLj7uXwWQAeTyPAyV
HXVb8SJOfuK4BTS+z2PQGfHu24ZkUS3rs3XWg616TzWgp2VEVqU2fXAs3p8waxw6
7oSI2f0wI9X8DUVLQtv32xOOxbXAUymDJgP8JPJ3TP0+dHqUVqhoUbe6M8THGNAl
/OLf6oTLUuyp1bGkhIuRVBp6K/fCofJqQJyjdXX/sPdDLSdgVdc74AV34rXQcmgD
5j+7XbeHUw7wY9liRRVfyw46Lkk+ROM3/dDKTbwehQs6f7H3EHUzmE8WTA/29hzT
fSPlcoCMJyMT/OIjJK4OkL9XCn0Tamu+J2CYKRHOaC2HGJueviktOXUPTG6aBgYA
Uqy2K/dKO2T554yURlOBjCqg2hyMXvPe8e9jFxVyIIq8dwSQC3y6x7Ct+uvlAkvH
R3emmccHaFeoK30Vsp8wPr6XH+cwTIKdfSnEIFtlQ9PBLG7z4PWaAxOumU2ydzUA
O/XIjAKllHZfIAlaIXuJXi0pep3aMxIUJG5VPsxc4YaGmC2Tmrt5Zg6Clag1S9OW
KoWWfkwL4PwgG7+yimOKXo9tm9xvg4uJpZrf3j3CusxLzlZd6V4y8zUyh4ASxXN9
kCuyVfPhcd3JqbQ6xXImIhbOomKqpqvWhxWcekX/E2FmoP2ufJzzLrV9vm5tMOmg
p3GVhX67hk9PAf9qA7ierAzZSGlgHRCzUWsM4rXtg1nt3AOXZ35Eukc+6VB2e/Rc
Yhtl1sIXUCgK9tImAN8YBn9C4eHflxEHBK3S+fXtloa+J9C+VeKuLHgsnh7bFr4B
RR1wA8RY+6+GiASMeR8pWCxKgKO/hRxxWLbp+661gLgp3RF6QkP0cz1SZNeAlk2f
i6CnFR2WXwJ/bPndSAOLrVpxh027G0bbcCc5s4mufhjYXCkosnxhgVWfNrraRsW3
WcfaakdYwCHlNPsVgpCGXAq6YHqWLZK/aNIwX36ampvpJ5rCBXCF7+jjHMCOEcvi
kJDKH4wdbb7SOcQcdh3jXA+Sld4eRqKquXcP87CX9qI9upkgtLSVQHRd3p0RIUBp
yaLAUM1JGQw+5V9L/dxgZNoOb0GfrC7xVhp8UlaXBHrfGvJt4SuYxXJQ7I2SUCg4
QehDxfdqXO1ckmCHDdaqJ4blc+Cd9741xFGW4VGkzG8oNx9PEknlrinCdb5oHoRD
CzWNCy6IdZa3YPGLlPJeproQr+2qgXY5WJyBviWCuylUnPNMHOyeyp3J9g9xQKQB
r3PGpFegt8yPWzRVId6V555Vixe6eg3Q2e6Q3JciWaR9sr63vFdS/8PCtPgg5u4U
41YN8PH8UMYsufhhfTAhfD/gOQvUezGyuxaL+Qjooz1g2qCUCuVukp1uWt3/nyC2
oM0hVCLgnl515eBn/1DQpd41iTdJvumlRcJeaVHAE3Dpraq85HGMNCSm9diZ+DJN
R+wIA63TKW5eZJhfDPGiEA0YuTVNhMumlAAVs7w6t1xADeNNxXOveKORA5nvbMma
FUPYkO2u5UyMFmBsm1stfnoS+Lc9zazq/wwLXYVgmeH0CqVAZDBoALBa+ZO62SL0
ScGiVrEes+0cH6bF5bc2ByVcSrkMYbdaGsM453GHYuuVc7Q51epaCKgtKshNFfrK
LxrUDl0aW3PqJcjhVY6CsFbxatbruP7TxjNHLUTUN9g9UTeBxa1cxCcrw2PXY7fD
WO21v+V1KTSjYpOyxfGBbE2niDwLgXnhxYrfZNe717Zo/ybWkP+N2Kw3KJv6qlNk
wrHNYgZIjALBS3iHRgVhbChWv8IxNinThO8x7CrX415AX2+EsxJbccr7hPHvxege
EwshrwXKTkIMaU+fIAwXhhwLaWwdr0x28TAc8GyH94kO/xCyO2lbKMagc9eExS2c
lVp9HFZKJyckIeDCRUJuQptOv/UFBzqEnntN4WcTtrG7nfilKm3iJHJTBUhNdsfN
Rdt4zfRV9mTukAe2/Ks1Wsz5k099A+1VbQcne0wIt4PvJspOmODEXRj27FokgeoR
gAGjd0V4lKi5x1MQkwvEhnv/o1Cxzbc/TOqYlgwgZ8iMh92vU14bnAUOjJx9U6fn
G3r/hdb8tnOqT+zxwGuxb/SCJ4SjqULE92USeJCWIhyhqV8pszPyH0Hp/kszH4uf
9I2dAVjKQuy4hmPUWP0Px0VLqke075LStgJmZg7XUM3hvcw91kOSQ0GWAoTLN51u
T2qpuNROOc5ExbapiY6qBPejS3zKIBoZ4C8Vc+qfsmC996yCn8q77Ev/WejRWkqm
c6yo/msv9P8iXbffje95C+a74mb4WVt3+U7kQzwxKFm9/Z2S/NFLobvsWS8rdQov
6GbvYAtk1zqORA4pcl2pSiQm6i1SqhrckIF5FM/Ci/Zmux9t9jqmg2EawtYlqrFL
wfwtBmwBe+qXqRdIM733W84SBT//BWKgT7LMM4wK6DigRbN3MJtnHoBdbdczCSV7
gRlwYXg4SpkU+VW/CMg9+vTZ1u6gzurHIo5s6VBnnv8ViORNW6xcP0FjRWn7YXJx
Wj79YglhMXZYNk+bMyyxI3gwLZUCfuslGj2GKJ0SxfhnWkwNx4a+UXRhPf/6jNO7
/bd6UovoLxgo9n9zl1/Z3zllU4EaY6u+SHjX7aRiMmRrefGF4GCvHhsE3x6O+1Vt
5rxYzQVT7lNoPPwywE24m2yKqxSsyrrcQQoc3PxPXrQR1iutNOR+JOiCetUCFDW4
PW5OC4ckU82gCHZlDmb6Fbt3JFAos28awCkvCGnA2EgoBCIbB7EJUnUh1UZa9dV5
zNck6JqqwFJIRnyTkkZSao07ooq4a9dA01M+cnrdrjkHbRwtMQKQ/RaRtv9rMkhL
YL1buW/fGk92v3XFOY/dtoAYJBag/6U/LEiWkhoTujlO0Sui9H2KSwVMpcsfHslI
ps2sjQun4co+QoN/JVxs9Yt9lim9vxwjm/ihBiyEcFavfkilSO9PFv+Z/Iqc/nIF
JtQenrOfwegh/NAvQjvdvpGNBqGmVQxy6BUKhKGX4LbSFZAe++wuGQ3uzU2QnzHE
osAIzK6r5DhYjw+hnGF63bnYi/4PdJzXplgJIxxhL0SCscAtbPDsUtaoQfsAGiBv
RHZjiUz4RvoaCS/+B9uA/mEEX41CyU26ixnFpMGYrnN+eQgxmE/kVa6gKcNAF8pl
jqpWw+LKd0DdB6wMJqUIhwZaVlbUE+Nf0VQ3lxcpQExmuAuzfEl7MI81F95KZ5SK
55N4qtDigBKYKAVqjgk/RuXMANpcQk8PkXei+kTKP6F17VMap+GeMtGZZfUHgpti
64G+c5ZWDCsw5+FykaZEcmhcnRniLuJOG6ZC10C7rSFC/f64Vmth5VRd4oFiCxbV
TmQiQTFfDF65Gv0u7lr8m6yUsz1/7tX75qEKb7r0i8WxRKYRqqRAlFxzEDuNCDdO
JC2jeYFiS14HiOjNbAtR78cCvXNisEiwkrI3YtLS2gCEVP+Iz160hYT8u7J+IYr8
cx4Cm9jbjs71dOrSztbWnFmdmhGnu+WnbYF7GcbPWNtezlVRajBHcSrIqSWJeFUw
B8OCaRl14vuUOQ00xzpNS/nshEckg6SKECCCMqdlHbzoFgucwWohQHqQWv34hhdr
GFYcrDS7SSWTlrsVfUf3b1W2d8xyWLVRqOGGh2BZAoYl2LV5ouTfjtmI+5Ydust8
kSzxqIrQglgjpbFPJlUy8odWxlAgR1V4cTkREqtzYAKRhi0sg68j0U7/F8UE9+o8
gqq4BDy6HDKQhI6jNj/ipIDcEBGKd9XNdWCoH+pI45YF2mDzXIVUsaRvp7fvgx1H
Gux5a2NFdnbB+YzT/C4gT1SKVGhy2rsnezmmu2UJeqe6H76aPR2aUyenAYQxuimh
fzd4Xze0THW6lSmXE2jOsGEmBDEITNiM/aHWetBT9Zo647Ybk1f7YhNG3zPu/Pis
k4uBvi4FGFVjOjgHyMFrNq/eng+rG6P+jiioWSB+OWdHrP9qs/JPOb33y+Z1bv3W
fXIJ/FU8CGk5CaBBA8bJzCwVV/nsBWg2Nqp6TeRsdMM/xlJIX2LSSHXXdclyjNPQ
y6sgGXa8/Fh1MTkfvz+OJT0pyH36fqgO2XQfzPzkVh5K9ztuJ7Youu7CJTuRrPxP
pLyE9pd4w+bMHFt+UaiA9WwbOMqukeGhauEhrkTluYRYqSH1qE2zjGYmb3ygRtT1
3DaAil8gP3obhx7rRPb3ppq+djvmmuvRSh38tPvp1Vjz4MMfctLU8GUNhKhYpG3R
Qctup89YcJ2MIOwXPtXQCcjI8CMcYe2debQesiyWmGBWCRzaC3NQ6TdD6S1dp5LC
C5B7+wmhPBLnHhRHubsyONxuc/hcVc7zBbchAdYBu/cfY018yrELbbsNQ3trAz4U
d57qEYWyWgiVipKokNghVZ2rf5JH/RijP/e6DDuzZqaff5w98ioDkqMK6TDK3f0G
9xI5u09BMrrm563oGaaxK/IrlwEv2qyfLkQTInL+uanLXlsrUqNACPQ2ksfJDXyK
ubmcxafYUc9ZgEgn+6LYbnw1kc26nnRuP+8NH74kiwbROWBfOsMzMnVQpGAEZWF5
lB/6IgC5e7MRlRk1jsVYwEybbDNgnXtcEiMTH/YY7nIdKTM40z7VdzoOOYmz537r
NYTqJQxTeK6/FntXLoX/oqrbBewCKdh9cx8a6+DF1aUJh6dGZGKbcG0kA9gWXvV8
niuj8rdik5r6aknKrTp4GL3bM2zkp0VSIUljMCcNder6JE07F2NlvYQIjvjqP+Yw
XwdLpU0nCAAHYGsWKPUIJqqTueskVbRgzSzFQXfOtdSoHmDE++PAyxKULXo3A3uo
cFVpcVetqIRb6ADUd+SePL3TRlMKNEFcyrCIFQMaBrsUVm3MyrgbfKx0g/t23LkL
NYa2S+FChk+Pl1APspV3x3z3wbVJLslebLmmq2WiYmiZIqLjmYQkOqiupgkhcTv6
M+gF7/OBfFxDsTrx+gSNc1jRHrTDpRbFBF/L3Atr2GQ6rVW2/Nrd9w/cBhBmkYSH
AnI4qnWIT3Hh/+xWLFt3haDBRVotKpOmOOIlqoB3pq5Phtb/VBGmOTZ3NPdNQEK9
AVCsvzmUGSRXQCU+2ubg4nXIG0yaBGsW770WLVjlY3L3NKOIHIk4KOjmMi5s76/v
uPJBz2XVR1dlUSyr9I/dLr1D+VsrP86nfi0a/6AQltXspn3bJg2Ry56uzFif6Nnb
uEebxKz1/VTgNwfK41hcQ8YXMbrLZLbAVFISbc2BoY4/DyBj2wje7TB+vqjZc+I4
q2dJxBDXqc/FfkEBmKjtvQLH+NhW4lY4bkXK/JAsN+vBHYDuDJdOv/0Eg/BVb8d/
TWz/fmzsTM3m5sCp37G2+Dj2IdwBIp/V4DxCTTSBiU4/UE8wnfFriiFWMzR20bh/
RoItJlWlypigZlNEQ2tz9Hb9nBZ50fJRAExAZD5KDtg+SOeNnyuYDaH7jGfSnOX2
k65oX0Hs0/yVPtd70ryRErzFB1mCfPONWuS2ILRXBqYeyHONhRnuLowVnOjXM5ZO
ZQtL0wQMMNIAFVgQ0SfSi9OdizeL2AfZo3DoIBeRRuRfBwwhOGjnf+7+xQPMhVMc
RwF+TuYpMXImdlarE7KOcsq6QwuLewF6lSNETn3lcispV65K3xdN0pMdvczE8cTr
EMyjZb5LXwzaxqH4Z4RIvwVyrooKfaPN+MSV5RafEyMojtmpgD2U/bgCEk9HB8KW
JPndnYKL+uhP/3xNwV5znxt3qkC9Q9j5dExvtz+H+Vq2iGAaw8qMyUba2rGdlLdM
b/SHnyELGIu6Ot35q1jqQ5Sp7KsSm4HgN4KkBMAxBjBNlACucSUChGqSGWV0Pkm6
GJkN2Ywch/o8u6AnfGwxT5L/XjvODpWjA7p2uYS9SAZw7JmWSXh+xWbtTxKHu/Kd
TFWDp/g97DPRuZaHPEYb6bIJfcfOI7cfat+mZ6ZtL1g5XqCTzHlDoRz6EVvmEABD
X7Eo/NDgFiSODb4KUQWW1oNJpesDQYqi/zv0RO0jKA412kIvU57OOav+L/EW6K+h
4MAZrfIxMpKBtj/pzk5CqZViDWbZoKz2fmVGwxMbMBoq7KQyUzB5gmmppG3UGIhH
mODGzIvQ90MHmw8+C6F0mKhynrAf3un08HvJOxKj9b4zxEVmyGD/NO73xBhpoj6d
xCl4EpVdVGQDBoKXB1lashq2kCxWr2S1bYOYPzYgqdu7RmVoKXmIs6tYDL74WJnP
8taGiO6qcL0MUwUYo5qUpf6D8d7Rm8ZjKnjEgQXZwWwsnNXOQlgLTc4qERSXM+DM
lBR32hE1IK7bCrw6L6wAgYTYxGN4GGx97AdYzIismmbewfNRx+tZU49KTseVoQSZ
2s4fSVYg593SSynjGcoydRD92NeKG78UONirvgFvXcChYirqgpSxFD2JyP92+Xys
ZXMx2UjxxGEOQzJ1CDeatkJrLc+r67VCrmMKtBiNxp4h4PuMM575m+XBpvB+3ueK
7UGha3Re/MlBogh6m32ttoPLH+7n7CoHzPPuUuWokaGCALVO/IYea6/OH5jYw306
xJoC3v61Qa6TeY4+06S7VJJszH3XJHoTtGXcFUZ5T/JM4T+qOh1LeEJWyQSvpNup
wfaob/6/mJd+CiE2EyIVtZvLnKAosnw2miwOrElHqm7/a6CXBN6yg8xcAVGP5QTa
dBdgET5vawHrcIPntR6bkWqY9kj6/SM8nWljcl/zBKqB4Dnu5cAAwsyCPbeffmhk
pSSVlGoVGncYFr41jRbC9gQTy70YPCINs8ly5+uSv2ZxYXOxR1RmewxHwrDmnp4d
CCVLl3AmKX3KpqgBIWbttgWM5tQmUxCZTM2SuJ0AYr0rAMvovIBQxLWx0G0gelRp
xAs/PRVqpqcBMHZtIndilQLKjSa22SZ2EC6iNKplIACYHV3RtxOy6zxLTnfB1QIT
gXr63WT1iaPixhh0660RcBsKMkQEpjn6FAxe5Yd4xqoCwZeYj60+QdDqTSmRUinu
ExyGlaVtScoysS+ZFbpdIGSQLSAustpue8lh3JsBoIV3jc4PKq2lM6EBu8/h0EiN
xuYZXVse68T1vvOXkfzvb9Y36Li9cI/np9v/er84A3sOqXnf8KIWcD8k7inMp1du
t54JFi53z5TkMkt4zCIVfjNHNfh0M9ytL3jo4Nd8LX4HUUg4iKW7qbnWXqglhjrn
ckiglP+jUzX49GTI3PXen5rXJa/71shHvisvH8DlUctv1tyBBLXNEUcndWkaNtAd
RsDr6ygomOz6nmIpJ4b4DuefUF7cJl7UCzTax2ZugmJ2gTIPZjRZD14ApudbMIJl
ok1G5Ii/FxHXXL5UDItvwb46TuXO+tCKxNh77FSY/V7EHf0nTvsNIgt3zHIy/aQG
3ngcbNtMyJzifez8aQr5ZMPj7AUKwDt+IBJ5T3Zd4RTimUyCbU/AYPCDT58158xW
T663QN2kPMmkD7JM5ZRz9q/8b3G6GGmc6z8wW/CWNI3Wx53LXsgqSt2LBmFYYRGh
d+RY8hiVHPgrV1bOb9vuWjcNpQETf7XJGX858Fxjw19ZGl/vt5motffvFpiR3vXz
7VKfxLYfQm65kEJIBZVXGFK1P/jCtNQ5PioGzN11dbKyFqiztL20EhypauxGa1M4
r3ctWMI5DwixTWWteyKFzDmZVzfAzvb+VIg9pO6RnD4qZjH+Yq53b0xqfQRnWpqo
s36+WRwjGCUDKuidHVmdH48ZG+jedK+26pHGJXsW4rS7xALfwzGhtQlIVUBnUoGF
fDBaHAePa0Cc5wiZUTubvlavtw64Uli4/+UKjOP5YUNO3JfF1b2UrSQsbAUrgRt/
wXQyBJOkR0CqbLuj0nbk9blEcx2WXFD8YoJ2p5E1W7gpHJiP3Ca5NBwXI+xwCdEt
/+WOIF9WvE3VM0DTDDhdgg2vwP6xwGpViU9gYxvA5GU6e/x7J0QmgDV9fws3JTTO
rvBXc5HBNo6t/ls9P8RC9hLp6Ae3uhBKhwveau3ysSzorYyUIq0RLXS6Um2qYiYY
srOXR8pB1Sl51NvSXp+6v9iMMi/Kki3vNgZOMwsZIWcAHVyA4E0swDZKggX4QoIo
+FR2x9UBH8KQc3uxbHJj6YP1XoNjcH9+rSST8ppy+/rY0soxRz/hxR/Lmn1FC49Z
Q072v05i9Ur2bKBbLWMf0qvmaeUjSyTWyhA6Dcb93UB1WiPorsrBuLdVvAS0D/Hy
I2graNUq8yv5mJMdj8u36ZpCNRZIk1kgj4jAc9MyAdS+7grh5z6tBCiCawqRvtwS
7c9VxJH+qCS2DicWQMtrb7d1KYBkSqFjFv3jYDav2Pw5mSnggCoQBSf+q/qfmbf5
iMJu+BkgxWnuPa5d+enNiJI3kCpPZ96lLGuPU1DP/ve3Y1jfMcn8UHyUnKwZkhQ/
h/Q8XVOvdKlVArDbvMbCC54O2W+9tCZ6dbbF0F/WWUnjFuAaRxHeo1I8+MYZ8Gkh
ZE8oD+hv47bM/bGw6kH9T1XPXDv750Gsemc7q+IkqlYmX2g/3ULFxUGhPGpEj5ei
xJe+Jaqoosmqudc5a2rnhNyNybuvNpzUbwzgNa34oAev7eYPylwkxeZysX5drUMx
3k6gFuYDhS/Gp6f04YG0zS60lMXXmGIbDvje3XgExzt5t0eMSmfglsF+dVQ2Q/8F
7PteVFyEXQ2ZKXsO2zeqFd4Wb+ZHiXAxaSVIyUbRwp6Q4rxedLN4c/6ASt/jJko9
jVV1SghCCrIt7RX6lQES+ounewgehfmHt0+ny2CuOthvIXg+A23BSaqxqDJK/rS0
Fp6018MPhGbkUSG66cg2oFsuce+nOL8mJEVA13WvWQMV7cIP2sjvbF5Ygt59ich9
GtW//2mBrn5rQ8CjzHCj6oURwK/AWeIHJOjqe1QbLWKKIy5WytsXpgWDjS3oaAYr
ungcVT0gQD+jzg3ygEgLDlSXW8xG6cZqODeyFMtkroL65I3SLurmOaI3HAb1MZl1
6W4hHPRv1S6x5dxL+FYOqj248yag9D0nt9sieFyTz/afNXhIO5eELmL15BBb7/Dq
U8UvNt/lPLDziXzpNUL/VY1n/b2X+UzGr6dmcRoXos384hJp76nrRC4S2p721RGA
7bcG6KGDX8dAxmghSQPS4L9UMTkAEa1M51jZ2E1tDjcvBqi1lkrDYWCImaNvusaw
H0BdnkzqcPdumPasObwdni9ezOIRk2A8Yv+ewK8LDt/xYV9UdlMkbJ3Aq/j5ddu9
G8oVVrIwwRIkQUypFT+lLTweKugCUC4mVjKIy8eOfDxg4xQ1hbcvY9gg0j7HjDkn
jbxQN2vcD3I8wTbKG1iaiVVjetgJgrIDoddD7zn52oOZ9TPIFp9un55MilF9dTK1
otRhfE3AAlOP9B7R32vttrmROxoy41NdbvdQy2c0yM7ipSGJGp/ubVIz3nnwg2YN
gghqQErgBQdup2RiakWRhhOzOQERJ+caXghKkwV/LZFAlnDnXH1CfnZum7RmJLNO
0hZBq131yKpAeMdSLBLOX8oD2B08JXaUNmzu7HZHqYiAt6+dTYtHJN5y4bQSiz1n
JEEVtHbfC1N2QJs7CnIVKhKZzFI2PsMdrziz27T6dXKOVnxv9z48WfoFSVy9CwH+
QL8xHwW2aPmy/nEgYLJr2n4J06USZZTWkaOLWkzZGkPQVO3bATCwws84JOhEjjgP
lZxDaCkp4LFKn+9/7zAdKZCEFstbkO+OJwRmXdQpRNQCyKDVwff881cIczPBwaYq
Z61FUVEjOUjrjBSAD83lk7G0X/ilttR+JLxjhSJx2BfLC6eGSnD/1q4G9RLr8/cN
2cWOnsYtdHOHNp6F25KN7uuCkq67GCveCDisQij9Jo3wTpshcG7hCYZpqk44olWo
vcCaD7cPnUgePLpn0/nYZ3mbutAYErrYaT4MzSPNSswKjBCUw/3dX31bwEnnWtcl
L0GUl8WvLuJ0h0+W9+AHLdYdUat/VihuLpDboQ3dBvZxbXyCEKzD0Ngq3SJD/ApN
hFCSHXhwlA0maQGIWkTirpSGyq6D+2XMOAkezmMYoV1dZBNeXED8rhL0eYA1g/7T
BWquBWpbCorh/NYujMrNUtnG9gLngH8fqLzkaA6vtErmpey/d0hRkKEBXI1kNKPW
gOjrxQy1r6jmkT0Ci9vvPjU0DK4PStGfp/EX6JzPspYz6ASWsO79ZlME7G7W4aR/
n7+V0NQJ7j38DhXPsNrk679u8vQ1c446BCjA1xjCLqUDV++mSZqwOoDqdRAsoz5F
5l5N6EXP5tN9IHEwHTK4ukXcpnWYLwmb/Zx+omTtDhqAAQzZVvEPbh0KKi1zuHqH
rYuOXJRP9X9OttCF64qkQX6P6cy5Z9CaS86VJP3t2ffTD0/QPui6WNE4eu1j33vz
JDI+WB3KvDqhUZQFdZKIPPol+BJBxPMusFNvKdu20rWvCWzDojF3m3hDJQdxcJ8L
x7Sw/fA1BmmXRXfvs3ytfsO3mtFvLt5HWl3CtI1euvuIj8TksKVKtQM9VUjGscMG
SiS7lJQdBLw7SyqxOpLbG+6DWBRpz/WjtS0REdYSq4QNLhqMdaCHyon/HhNCqeV9
jbmESNDDhtNNZA8us32gGtx7naC/FHT6VJPuBRFmIi3IE/if1dN8vRCm+pfi6ZIF
KutHpThwJfSMt+aRiR/YmZcow2jMcOL9zuQzgSBIzhZePhID7PzWnEOWlRbZm4QI
Z6Pu7xavacoO5YSGcA6owUBn49P2J9RjMh+NTBa/3Y5YHxgadnSoDNlI2mi/P2fk
jxBtWVK8PavrXPrX+CW+IPVhMqhugpbbEp5A+eq4i7/vOPUaOn0wqkR0U6Q5/yjh
jQR9SKovlrottSGwA4OJlO4uD3dv+C/NJafZL5t+aF4di/gBzVxULP+j+h09vXqj
gs1p3ZvsS891Am46Bh+nimgikUxa7b6JpLRTOJ+7SWrQzfOW+828ktnvzcgO9dQW
MA5OIYqLdqbR4iAy4r/dsDoLTsrrX1A9Xw9yX7jq86pTXaaoMmC3zqip4OAHiioj
/+qrfi4ycMqtd7qJJYm54u50ArowRykNDhFDZ8p3I96Jx7qcMiYQH0jee0tYpzPp
yOVjjWW3T2BGsC+uBBuKgauGdOcyRCzihYMd7bsF+yq+dUjDyHhS2EP+bRUkQnta
NvXmKs2fqbnUauHFG2mb7o5tUmIP9Aenq22rVwJadqcIWEXb543LpZqIYbUnz7IT
3d36xyCiOlZlkzytHGChslp40cy/JiP5OnFTdhybHAtjh0oJ6Xu+nOCn9kPu/M+h
Y0M02CZ711GnrB6iMjb3cpYQbVpvGEfVT9iqKz7SP4Cl9meMGW6s66fr7yOFyGF0
smLjNflib6JVmWrXdSnfgvRpH41k8228T6VyEB564YP2lKIO2PdN+0PJwX3Sxzqi
zHgrIzsUHawalHsjGAZSm4Aj1QjHb00La36od00ct6eEAQrNHxmh6XmHe46i97Az
0aXVbLUQCO2N/KGEhzp2mLxXcFVT9420o/T5lv1X+ug2el9kykhbf/6Uc69BLyzh
XJ5m5XtzSWr82LSS1vNQQOjuM4dsONFRjN2hkndgDpULFPy/2P26YWvG8y8cCC/4
Czg54JHKnX7M6lnTynYXBMrvOZGLdNmPjvOJ9jFJp3pbHKDHWuq/tRl0EgigRulS
5+0yB4KsSSabwtM7bteLQCQo/Ka6Ye56x7y5dfubYHjduI/DgqV0AdNOfVx3cvWv
m/XBPaIzFCFcfyAkI20DzHggccEsu1LpE5ZccOq2ootEHC0Ne7MFv6Klu/2v3/f/
DJuSH3eEIW1Dt+4bFIjE9oawnHwGtLI5ysYMmunXFe1iZeH2CqJwwgKXIVtdHmyM
OTs0vUDgfNttSeEwQkxvANCHn3lz2XtGxf6egs1kkQ3fIdLz6cn4dIs0yrMwNGBD
gpTJvP22j24ONAGwjEp/2scz0WPo0WSr1gGf7ty6Wx+Ek9bg7W7bTAfGlxD0w6VU
xgWUXqu29UBImEYYeJRt1lGbxBkZEcfA21uU8Xq5ZAG0MirOSDj/zSs4iGaFCvmm
EIjdxzEMSNK56+rE0KCaaSQGTYRQzGqe4H628wwlWyiIJuzv1Ux4Q3gFRwo4Y6CG
HTJPb+Xjfv/5HSBeGzANarfjngN9JZMrKT4yrO0X/By8R4b6z1NtP0x3oE8Wgm+5
9xvtVw2N3FXG7bmr28ul55YIQLoogD57+4pvygViUI/9jv9IvYVPnU+CngW7BmdH
Vg41qJJXh9VBvqBpJROlM6+65xjuYguVSx4bh9w5zbJJGd8M96GWRv665LpFYB3C
qwSxxOmbBLIJnpA3BzH7vxSTT+pgl/iQ1eppTI/Lk3PWjjOwtHZxQ4MbADNI9H11
NbHHbhwO4BLuEYX7rmVAplYm9YzkuZAy5qPI0YGkQwx3Tm09cyEpmHsdMLA7LO5C
1KlpIYWr/rX2Yb2CYW8/oHNY2MFxb6hjOD5sDVBaDoeVn0PkI2//XHLxYTXFn4h2
wjkLYYZuGyfOngQw0x9WrazJ8HiodWmMnfQTt/ud1kBpup9cI0qPuKOnHtvwuH8G
tL2oVdF1COSQniJcwj5KyYSnWTl1nirRt/UM1FrcYqMK26lvEYPClQUpYaWsHSgl
B8ggx1OLnmWqEbKyWF6R42cN+ABi/cmJ06B9a/Jb0cHCmKsFv5Np0NLMuwF1BoGA
yMfqtm+3L2mydNJ+SsnjgwSUXChHAWYLU7SUhQHQ9lo=
`protect END_PROTECTED
