`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yVr+ISNDBCDvv5DKHWPrQ7RlIOwAEIA84hJZ+0MtLKnmHBDwmcdBOOkJ9bKwXRM6
7PIbBlcK5tv8f0rpzVu83CXj5bERJOvYe2DoxhFIa5hG55W5FppUsHk3uTbukUCG
VkeqizJ5WqhVLJuMALpYYqz/Ch4sBUojES5TpGqUdH1aYIJicRNOckSuV2VkqTLd
ZLwocgWDhNYWtYbXSiiFeshQdWnwhzlY0P1vfi8MyQgo5WxXBpL8KbMzmdJp0G42
47cWs1CcfoVGi1gNSajg0rwn375YiLsWkQHlnjueLL9lohWgUSnGH1ChtFSHgi+Z
ssac1StbkWcK6VNr4LSIgank3tYh1heocAUmoEgSPq3TA7qrplljfnG034awaRwC
dORiL9KH/p09RLdNJ7WVC3ERNTjWvhwi7/UQazg9U6P28WttS/FQmAbk+QdYVk9m
CEMN00HuFaLkSeoWGy9zURjFLCGyg+IJv3adwQHbbnynAvfxInmPVo4M9Gek0XsD
b0bn9YYqKtNo3B6HzZ2JOEnFqbv7EqU4VL+nh0eKpmg+X/dbksbr826zt3k42Bpu
Zg+E6vqAMAT4xh0UIwu2M3TgifiN7YH7/r4XboKVhVXvDZ+/sAOjm6qNNXjadHWd
Ghq9jYO/H0qR8ZrzxbtHLyfnnsovj9+hK8ctYmjRU4pctW/QIzGtKiCQNuw3q751
CTTRbsVNt2mU/wagRDDkAo7F2mssiuD5jF0hAavthes6QTiMuGwL5/xqXjWaWuFA
U+rR6sr2K/YLE/37krDjdvq930qrxbJTUUy1DTwQedrUu2dxTGIO0Kqb7SYdWq0p
lU7JoZ1zD91ouJL2inTIBjxjzCIdQNA4siT/z1ZMdvbe1EVLD8LLtWnCDn0RgQ8c
0xZptwFUbJHvveWbuEhbIqcgZ77yKOZkhfhoqmlQ7HUbSMi3oS9hO5NBHrSQhCtJ
zSoL2Xejg5cyJapWJ2OV5RXeqIJRiub/inXWpqq9duQzfKgPDU4fhTXvC1szkU1n
zJKPzHGa+xo1hL5+Vnbybu4vujKx/7T+IgO0E5UiwTgP25bmPVT4ulqPSe5fRiuu
AYIuNUf5b/Z4ZcCTOdV4p2GjkXfPA+wHM7wJJvS0+mMiOVbAGvt3dlqgaPJHDpbU
xXH/KfarTmIFO5FBC2dhg02bNgJWLVe9wzDr1oAFXE/y5YLjLVQH61D6qf/hyg9Q
jsaSGdxgEh9gPHUvQPWTH7Q50fuY8GXOnkZ3qBl5kaqv16s65fImKs9eFvFSqYBZ
SFCCpIDZ8JndHDYsST0nuJaLP0jiWwZl7KLX2OaDHWniFL/l7/+MGJerzbWyLD/n
51+exr/7pHJPAkFFOACJCLaVIZpJ+xIVhvzuWEv6AU6JOpM48RJzMAd23b0rnPxi
3rGyJHSYWZyohdHChZSA/776INUMf4tr0fDGKdh5/VJtPkAD484ZWyDkJf5pWDlj
xpGnJuYdfnt2xKGNzdFM0ITqEsD30atupTS3rlBYWJCuBeEUKiN5VqEqI4LvOgUj
maMHygvAIrlEc0Eu+zDzRQEyfF0qST41uhKmxaJ6Nmwu1Z9Bu/1/nXUthMDk/COj
hhO6PSR3G4iCb5Hry+T0CmmSgZ+HGhquCJQI3BC8D2MjcBxPHkv/rHP1ZGqXAOt8
JRq3DPuv25XhAPjkjnUVc3u2Kv9kgE4LRohf82RxwAw/JxvJU5sBetHNJ6MHi2P0
975SkcSar6OlD2JElPTSll9G85l0hb+4qOqwzfY39sA3MhmzO49tIrP/smZWVLdh
11yYCBYwbgIax/27gwmA2KUKo3TF9EFM0x7MtwtPDU084oZUS7uEvHXCqMbo4u9s
X5XC9x2GUJDlFQ+SCdj/826YIjNS/zIEeotZzYwXAJMFmQXBwDP1sR/OBGtvE5cR
rBOit47FYEQ5GxuYER22b8fvPWBSZ3JHwe+xLy4mgzpLR4cLs2RiU1WdWzedgzhU
`protect END_PROTECTED
