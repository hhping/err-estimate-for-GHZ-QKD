`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3zvq3cPGvqnHYhwPlf5cUPpcpG2JgL0zZ83zVF31butBJU7+csn2BfiUutzvlqTQ
hC83oMx127ztXeKqKlS2lJE2pBcNQ5iP88SgloDtXeEApyI8fWw+R5wRdF3h5aMQ
ICghmay1dxqU72ATVdrjgT3BC0XWg6RKxtxcgDRBiK9prRiF3uHKhlaYgj5BuD2E
zYneh/eaAzjbB7IQpddvkgT7FfieQZjRIOPruh8qWb+FDE9qWBiyULt6HPly2tOb
ik1eHbdy9DE7rqPrpjAd43+BKxuA3RWd3kWpQg88EiGHYP53O6NgyYXe+z5MLiZD
9wd2SqhJ78nHJuvv1iBNduAeWW1BNWDVqMZoe/bGuGpg1nte90xxLjC09MrkyFxj
SEJLmfP4kl2bmHs2UhIcj1vtNZ+qynhO8yX60OTJyf6mML3d0vexfQAJYYPOEwV6
VADXrRJBeGqb2KUSjgwBBlUh3HSA2y6cBP/qzRaEIZzo7CLYy2RgxypPYUNZffKH
qkYYO6zv68QWzs3oV4UC6O9AgjVAhpoHDj4dG5vpx++5YKCYpiWKrRpvve4a+Ibw
VxvJ4ELyRlCFk8X4bu9HNIw/P8O9cxK85Rx8TDrLKSu77O7ARbJOIvzDABQr1t88
8oG21cygHBlIAQgKG1A002aoQbSpHqr2Kw6YYQaGD78n+ButZtbd9lIdShjxPkqs
9AOi5d0+pL1GqVaWBY/GwUMuUZPEWeTnvCq9X3KtEryJseBbMzlo2npdouIQs/r/
A3W+XGZCXOxThHM0y0VexWs3ETfCH3T58zvp8U6KYCPbYSMKXR3e3KED3l9df/t2
PpAOls2Uw9JiN3Sx8DMXCAJXVVQzo8qCAl+JBC5f71aMXCRixU1hFpzVqiLeqj2c
31t/Mh65gO8mn8rFMCeZx4bDxudn4m6VNcppvjxpE87fYY63U3qCBRlA34ZkLyM1
XN/eaf66XPCjLvWW4jAG3g==
`protect END_PROTECTED
