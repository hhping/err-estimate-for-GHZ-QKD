`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vywoH0o1wvKPhqtCKDgUOIPUPdIB0vXzujHlvLUx9Yh7AxJAGx0ZWU+Ek5m43Z0Z
R69fffUyo8RHMwWvRfwhSgUxlYPavLvY4TR0L6/QqKZhYtpGOU2rHZy7y0U6PFtf
I30Rgxc6kS0e6/iEADEV+7QoMYdFiSWpAjlpKh+sAP/mvjnLdI4pnMXeroYd204b
WrHY16/BO/7/zEMh68O/2nZcsE7n//OG6chO3w9ORz77rfbdKubQHSgFetXb+EaM
VqOPf7V5tyUoLQV77azSpaWiicQvRdTBfPSESebyLXAATmLZ4Hg1o6DPXfD6UZuC
GNZ0VktrdptiwcV7vjsLhQpXY2QmKjogJ725ZtIOaJior05n0wREWYlkkcW2ibTf
sJs8pfx1tI6qufrXMSGa+pHMoB/utiqheoFr7KDQkaUBKJjbzKT4joyJVFp20DzH
H5lwuE5ttwUPBhg6bi0xm+oRGkgYSfBYt1/S3JgxJOEogND1ISkucxubCUauCBr0
lvjBi4FGTVhZMhH0MRE2KKnjyY95QM0LT2hNc4EX2tRFbl1Ju/F+/0UY0YlJ9p+s
iDtN3I6YdnusGnpkIdPrC3PC5NWcFnTCDQuPGUO5ZbJq9OSoma3yUHzB+Vmb8tGX
2qdvhQh0NETKpjLJhH2XVk7EnG0Op/n63flvET+sybsXToyl7IC4kRHOa++gltBd
5t6bHc53k//XcwfQfUy5+g2dBFGtkfRFAO+RRrx0Q8uzL2ujhOVheAlaQs52p4a0
Pu0ssQiFYidnK0dHZM9dr3yf++M8VuuGV3deJ/s9CnfgbU6QBjjxOLXedz70ONA4
7lVD2n05nbegA1RrGnlARsorbIcTZ0SuICkHXmozJgi3XMoz9Od5viDo7jjGn+El
WEv35mxxTyHCW/7Z4KGFh7VOrBpnZ2vWG13t+lQYVfWPx4DIRgLIGmGoH6xscp4N
6tOGRwjCogCoAM0E9hv52lJxqwR6KXark3+TQ8nuQtMguEbsBwskJbh3UcN5P7Y6
gCUAknWuWmsx5t7+TkxO0ecL+f6Zg5lNXVSSGkzbUKNPyR77+imiQFrvMOhcrApl
Hl1HY98YSULjLK9zjqN0o+114PhEj+WK3cs1Y9m4fYx0ugq/FMXvIWUW9jaUppsz
`protect END_PROTECTED
