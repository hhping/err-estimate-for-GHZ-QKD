`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tgG8bLe46Of6OkmpH4eBwqqUYDLuVrBAf+i3jE5P+HCVJD8SMvCjuHgxbxX54F56
1x0XfGjMokW5lqHvWGPQRhXTJIezEsBDEmEH8Ud7gVdHtBlrxcQI0gi8Qv0Ua3ro
aZmj+rN8Uz6zwvqcOWeCAFotACthS16/bLdJ4L2Nt48UGGc7qqCxKuFeCptYaapp
RboJIN65NDohk6pnVFXK1lKF19BaxXl3L7a+9Icn8WPJ2GtAJpBJVjOZ9jUx6uqI
OpkMOdHx7OtnJm2dQfEX+QY2J6/BMqBK5vRVsxv9atJOmlcOp1JIqLZ7c1zNJMWz
WtcJ6oADFiJ0X8uwsbD1E0juot080nuM7DFLpJD2htSc5HI5iTX59AAwhOLxHb4D
mDR2jBQy3Tn5fecRDEy2VotUjBkfHyWeqOdfelR7kWXvfeCjkhPBEgbnr9fAM3PK
PJTn9Rjvy1I94qgTfosdK7nshys+Jy9pn4knwObdWSuLgAB/Auj5O9fTmGBv6HWf
68cjQDGk04kzyDATtP4TeG5PjSI4U4rJMKrpJ4UToMXV5RQqxSZK7UOos29Vznm7
6EZ82FF2QZSM+6ujsrgzCZ9p+g748dfKoYYgZSQrPbcnj7B21XCkGizWLMwcvmzb
+o7yGYxR2Lq0rVfVC4Wh+TbA2g60Ny/6qxYQ/UopgqFjtrCQiQGvIIsobHdghys+
knoHnUcxGYF6jIIBUft0bQPaKgaG2xW5DMRBdbrmlqAQ+vCUwgpARhd+Z9mL38ne
efipWs6GoBJ8OKrfrD8nSv5KsbMyh9F/Ny1RksCWxC0xYUPSJ6mc1tLfD5ldCulF
apuJXrQgxZ36ezLwhe5ofpSxn4FRmyM5hH6BcDzQQXYThFZxgLOCTcnfxlBnpv62
LGxLI63TI86fAzhmm3IDHDkqSazf12yyle9cd75a8rWxgYYkwIPfLK7hNjz8sKOf
Czqq79DJD0OtbQTi0ODMQGK5zYLl/uIoyR+xbTcsi2QRVdtnHHilk0S2PWyV/CU4
eElAFLvvn8BsZp851/04A429v1f4q1/l2ie6meZmJDvRAVOqG0Cxrj8sL6MkTTeE
mmCGZJethRnb/CfHfsQl/py+Jczo5G0GuAEBpsW4hKlhL/uOdOiJCAGw5/MdpH/J
7xohGYqXxiXN6G+UVB2S7d0T9Q0gzlozdOZM6e7t+eRO2YvZZRwBFExInpPWSwEE
UHvLitbLeJrcNK064ngBLwtfALSHTw16Wwjr8uy9/jMg6UWKXZCnddn+fKzT5/oR
93dFewKiDNhlXzkgy92mNxctsSQOvd6c0hsu3rt/dmYmz0Pq3ZxBSVHFcYpULSbh
DjMMm4kimbHHDrDiNm0TlFQPDw5FO4frvT3mFxdmZ20naA/YL3ZFMW2UHA7VZUps
x5QDOW/Wzo9ce5dnIa40d8o3Pk3cBljVUk8ZiF3S0gfF3u8bnzjxdU7MTp7gEqoY
fsaiD8+AevTrKnDJxzxWHjWksTmtQR6SeNI9pgQmasHrCNcwEQHJ5QoNw/QKVGg+
RjHZYfeEhHc5q/QwqvODMbwe2EfABo+LA4Ue0uao927lQE4s0nGFu+shRx/faSiw
vECxYi3MnQf5VnMrUoOmxyBtREgFO/H4C/dwHtMHlMwYQDjEzK1eZjOpl07xuMun
KPAJ/b0EhGshcRElOwvLWJlLSds3mvb/HXoRuE41FNW8vH3D3yItqdQgWHBaQIEn
aKq6+l1xODB7CUBl3110lhqNiuazDJyKICjPm0zXAjaURcbiZDm5zcSKBLFUBssC
xNI2/zN2MMxR7QTG1meiRmtc9slufOo/IG/E3TAAU9vN3zxZm88zXsXJxdbnCDgg
ytBIWLceXeqSD4SfgfXAOnSv4jKiuBzJsT+g8BGYSgGTLzM1HsDqUSdRuPWfXIhu
UFpcYRDAdFy8YHkENEblq+/o/mb67s69DCS1XJdqZlF7X7LCeHARxL9C7Z+wygxt
SC4ycIIy+8uazREpvkDH4XhrldfZUUPqhlprGIoNruvlaRM1vr8t8yXVRMPUq9vc
J1dXRL1BiGGpcf3V6O+lrHVLAkClgRtfHLNPB4Xs1XEj8xJt1uv+9kW0ClFmrVpZ
gkYWiJ5HT2IWebkyqzH1f9y4NEpqXtIqgZ+TaoyxGQwFD91YBPIvL34WPgLlZCAi
KnI/ezXx1bAP1+c2CBD2spdP5kKp6OKLafAvjo79SDCkTvQaC6C6qUwbKvVZJ/+D
q2pEfhqT4PgPiFVa+u8NHIb76Ozn53DlQn7J36K99okEZ3aGC5DuSa2mJQdVQGKG
iBSwA/bjvVGRRx2tkxYGIPFzs4ZoVzzXZv/iNNn9O7e0q3Hd5tDpVHkPu0qv2NoM
0IaarEWyI0EFo5C8tagfOyHG7ZAYRWx7Ps/UstE9iM97xKwifbkwbjwhQhaeRRQY
TKouxV6jKHJgys/6nGNre1phoZY7ilHL6KqF5sHpyuzsNEhFoGgzog10DlRXFZ9p
RFlVk90Epb8NUffZH41MRP3dtMgfwp2BX8+RJZRlwLuIxry0XlThUyt3n9Co02G8
IWKmq5l9mc9ve8G8kchUAKKySbyjZpoTQ7z1OFBD1zVo9XFjMAtOIctm9KWhwmw/
GJ4vvHht/5FxkgIcEqqY9ERi/KD8TdO1g5xwbCWvvUrBjuQYsZz8G9xT4dCMXtjq
6aG1ovmqEXHIL9wrwi4UpiQI7EQxPlg+ZT4cQRZco9wSE3ebS0CSj/z+Uc7X05B/
boyq0cE0+TqEnJkw2BGV0vunNTK1LI5PUuF1mWTUsWLxfH0vt8UfnYWGP6AUE6hF
1/H8XMERZoD8xXOWJTvvjg0Nd80qSAyjh0wEMJyqkL2CUC+n9NBlsoNwaMKoc8de
NSUvHtsOafRA2yAuAty4npyfkHON4o/3UdSNUU/Q2KhZEtZuKLlpbAZQXARLFwTy
xubKAw7L9vY0wdkDonaRHmXh3evt6/Ed8TsOnWhj/gN08DFjTI23UgdAq1LbIAPU
s5M9HYzJ0pxtOWIHBzp5ceLCYYK/4+JRDXwG7HebBsbacrQ2pZZ/KpEKGIyF6U7C
GZrRCZrrdIQJg8i6sr0rsVeloxueUbd1UYIMLfi1q//JYNdHi5Mq1NDxgMxR8Fe3
cqOpw9WyYJ1efe0SlL+IHXxAk+g34LLQb0aNtMT4VtxJbjiCAV/66HytO+AeWcHl
Xz2KyeomGybVoc8YVokRswendTSJ34zxuJ/BXUcA6fGRun0Yqu265otxkwvQ+wPT
gE1D5WnuvyH/O17oO/4MDrjfD91wKiAdQBwNRt6YuYQGQP1DVJdQUTpVla/d3osb
65RTKUSo6sVXYsRTAOX97XR5lEbI5nk1S/Z1GeJ+4YhzyQ/jlIzkbORDxUzPrdeI
0p/8paVggdmmIUYpqOpkIkaT5wYzUq7ZaYBmbvMAPrMh3RpfthOZIsBT2TzkgfCV
VXhHdDNaAnlC1MBreTSrrGelYEO9coANp4MIvOFwC1KKynQclx0X76zIZlFXbfMM
vFoObZgfsKTIWXflE4sYDmMIIpRYE5dDGLVh4HJkhKY=
`protect END_PROTECTED
