`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PlxH/yGM44552ufX3kYpN0gruBTLnVoJFCh//GGXzuUlW3wYNI3ENBLD/1zhh/XN
l5riIceDBeruNxMMK/w1jSwUPELq2R/GgeqCbfKdrZW7jbam8JrytGRHxoTU/wUZ
VJBoleRP/J3GOP3n8ULvjWB9ylWj3RHljjFPnsENNSh+ohBH49g8TdnWqVGxv/Zl
8CcaIlB3Q0oWFfDaohPqiq9Svie7I4lf8FrzsKrxyNaz3dPvwKGJN+ew2vwq1tdH
gElWfuybkGjIzHswuWZ8RicfcVwsMUhl/qh/rat7pX4UPCNnCQBzYDnO8kXlIV+K
Yt5d0KQk156UwRHILabiNDSih7y1EerNGTB28EihGsvxtFSIxbp2zuqM1wNjkc1w
puSBkGp37etF3XKm7zNYoZdCC/IBej0ah5RyZGSv3xlUeFL84QMUwQHkRk87yqbx
T16pDGNoyIJjIK51EsJ3RuzMdfK7FsMbuv9LLcxKWSVQnghQks0NfTcy6E7Vri6y
zUFC6KXn4wF/vwRJkP/Cy+RIV/exjfcSG4d2rJxFXBwqRYow9XP+fsaY5NapG2bJ
LIEfqBNG4BEJJZnGGrlQ+whEza0gLXwP3OOGcvgpy8wiiVeRFh1niVl00Dbeg9fC
OorDxlZBhMveoj0BHHKkog0a3/4D6nltgFWta1ouQc4nv3sUk2cxlhEsIrWDfFYk
hO1fG/q3XiBWFBWXjkOAjWk44JW9UpAfvIfB9HI2363JqDp+s5bn4AN5MbZjmmlx
qYNNEz6vPKrdwxsGqETvPjzLw2+7hNGbBdJUElbrUP/bL60lnxCXovpyblF0z0pZ
le2UdCUgj1fysMovbJt4ScrPSu3Pp8TXLCwAN2HnqoJQuShWiFeSrrPkWaSdKy55
s2Tek3GyM+pUhtAMV2Dgzf670zSyB4k94d5EnF1a3ABtMXg7nQvFUwu1VEtlA7SD
6vuKDbA8w3DcKKvVTzWQXjju0bunY94y57tw1TthdPVbMhN5Hn+UuJ36oYrB8ThX
bVVw0zfTGOJuRlkTBRglTok7JyXGevTCov4w5XpKo2/T3J0SeBYyaWd9VVLGsHE2
vV2Dj8NcV0hKcRwviYN/U4ziUvAYM0M0jYdBdOo2lyrj5boyggKJVFfEHgIHBNrf
rr9I6pcejwMkJ63ztIIRACCbsrIfN7ZCdBqSignHexg=
`protect END_PROTECTED
