`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4OCwhqxKtS8VzMPrKOpr5YdyvyX+C/OXdTitJfTarNujZoWM4WZ99n1GRICwdFu/
VIN6VV8YHv1+5+50cgjO1or0P2J9bceJ0SfjK4/oHYOWW48fps22vW74P7hxypvo
B6zu9x31bbjsUJ8j/sfuCrYRXNpDNM+nOB7H8iekRlc98s1TxpXPhtp+xVxp0x+b
LEllwlHZHxUeLpS4yj1geKlpA5zifP/BNAQWEJmSYnwUSdiw+NkTjE9C2rmrnq6j
OPTGsvhw8kpgzInlYCSEK15athTc/fIl3Yc2jxcwu7ApQBu51yLi1/tZZ2/bHx9m
+IycHauVmsrJIK0AsaWKYUJg7mK4t61Ihzmdo2AaRhZjxf6adV+WHnhS8lXg2s78
XHJAZts+bwHupyHL1aDyXefodDuLN+yEA2JIyt5bmj8=
`protect END_PROTECTED
