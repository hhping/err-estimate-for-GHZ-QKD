`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SJBx2Y5AzXjwfGY4nKqqy/GQ9tKZRv++/pDs5GPPlTYd1zLOfVNM19Dc9QK1vx2c
WDXFAdqzZonfe8aLko9QJ28eRbxZEV6M7xnajZ5sx0EbWQN6jALby3WqBgtFAoac
xGhMdbjOjLffS/GbAKTEvFa2PepK7vRpvgK0ctOBIoS34ED8qDTKb2kw5Is/6RFl
dRMhKvAxE5RZOS8YVyZ2uQ9xfHDaNbhp6aKrS+a0qIEpcN0wjqNarkTVAh/cXqaJ
nKbCEVLDWPeNWNg9QYVlA8sqsFd1zMiNZBca9QPUDFX5+BG4vxccLESPNASo/cWF
DKNLicrm1geEN2KlrLXzO8WoW8C1bsytADnlbITykifiStKcY/CsCxY69HnjEkST
q6G2o92FC8e/828acJ5TaAUUfSgvHjJBv41ctnRqSqYKwnQ+iupztaIh4m8TUagl
Ux23CmstEZLqGoiv6PmJAPromGZ4ofmoFECAQKdBtWegJRLUcCievJuYQ8oWuDi/
RlXyw8mHN/WTjJhvBZJ5UzvilV33v9dQLQ2Prs1hKmk=
`protect END_PROTECTED
