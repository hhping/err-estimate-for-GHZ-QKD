`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gFd+cY33XFMkP9U/K5/P+WFmgsLeG639+6EDHuCryUnhVCVDnPoM9+hmvY5LUX7n
g/k1y1ZbrZoD8bOKaLBUKkO08y4hGZiMgL40H+Luo9QnTqnfptAgLyzlc1p6/bwQ
VOO/TWg5mCigYqUk492W7Q8eUsVvt7XqiL5q4Z4zaSVKmRrL2+VNqEYmJgIzQ/hQ
bv2NWemCFKbV/LfJhzifGlgeX0SpnTSNKuJ1Hq1kqbQqfdcbnNTWRsj7CM2wCl/G
gf9xy57K00felKBaQynNX0Y2/Bh8lclQrGZVbJjtDJuCkWL/zpCZTJ13mgc8SIin
EjmYEFxNFX3yADqfzxmqAmEPrRzYvf+Us3x9aH4vWjlqG1SUh3QWZoRVUB2LRj6j
lvJT6A0/NstqdvHJyrMaAHVt7A2IMak7Tscpaj6l7X8Lm0CcN0kaCPkDxf1XaEwr
HmKi/AqW97+OoEAhONWiWs4yyTUKhPlMvNy3QQsEeQk00rvYDniw6JJhjLfh3XoC
OH8Tj1wNOl834M9ti1ku3ZlA5B25KqV2xXu8lXn5Pzg/GM+krMPsDsWLTwfwHuIO
D3Iczq6PyIBUvPd3cZfQmd7JRHbHa9XDTQaepOMu8OyK/ubbXaweAAnIGfAnbCb0
uVy0G/0BpmAcvk4rmNZmCQ==
`protect END_PROTECTED
