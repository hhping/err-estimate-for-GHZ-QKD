`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0YyrWcusY60/LA6h4fD46iarWcP0rquM3B4nyjvP/YJZy9cBhh040Ou18my3gYTa
oGtNNQYnBfredDu6zkpFjsBXkVetJCxQ6+e55ANeGWXey5irdkM8yhfxq1G9a1g7
muSkaBIzK/sy5wCBNOvgEsKfx1DDmWTdO/1+xxsjjcyMc/KVJDys1BsyKNjM54rW
X9Qg9t5kaB2bIAyUHz6+Ef1bKrF80vuW11Pe9g6ZZAov2tqSbor3y92CyYPSm9xQ
NaTqBNqJFb6IigJX1LXIjLiWqrK6ZI9ynq+U24j7Fr1Y/Kymn2ZUJkHuTCjyWFXh
1sR5QJfaxfTCr+2LcGA4hkmp9zAHIu+bsb742PDebogDb0Q7FXLskckhFaY26131
F3XFk1XkKUAVeOABFEE4OZiVrjBIKxYE0vnDscah1hxjw7DaLei5EkLsOy5Amkso
ZUrjVb7HFoJYV5smxXPlFcpmb5Olep5ugMpvZTKMNTY20gP1rowsRmz73p7ogNOF
76COhgY77HBj41OyXmMdXC28Q9Wb5C3MXb26ft1aAlEdftr+QKXAmbhz46PWZoGE
tCYjbxoxScoebCk05fWDicWCyL5E4j/eGs7CRLy4ZBzpSfaO4M6tlBQxoSPwSaAe
mUignTaqDyk1woAmIj9xH3Qg0bg1V2O1wodj/asUqhbix+WbT2cwySzSvySHTVFE
fPjp95D3FHgDg5Uc2TAda+nQ8Ydi4nYFMXSseCPgjQAo7Xx4iYvHr0uqzZl3iTtq
rRNa+eR9LF/9wgF7xJyESBxebtS4o3wDOzloc+w28971AxL8AiKFeFxxgcD0eZOs
aHFkg8sC2TnQFBA4FFEahTjl0eJ3d5aCIiw98/IjzeYWd3WHLuI8tap8WC4oj4Of
QBHfSOtEXYGjlnKU3ZeYyMtXZ7iXAhhV1MkXIqeY8H62vkQo0P6GhyylDqvgAMT2
PSeby4p4/HEXka01sSRbgs0Z+dbn3zBpPJtuht3IC1cL+ZibvL+tGQ7GXvVVMKQ9
WeresHtsEBmPY2r8DDFPs4y+0bMQRkyzPjiw8KvDGVQ3AXp+hPvnJ6E2sec4Rajg
8iXUskRg76X0U1eVoQ9T9jpYQ+26Ts1hBb0Np6GxYil4UMsUr2UkTAyEiOHZ23Ib
sqXh4Z4S5g+lRtU0hypryqK64s2EJ1c0MRlWx4FqxbeE89r4KpBOTdQ46vNoAAyp
wqq3JysCdirFgL1VrebpAKYbGxV02qRI+5vtwcZL1h1N2KToYbWlN3dXTCXRSrmn
eMHrpq2ZfBkYPBYWJeEj+KIw91G84Z2O7FIMYxzAZW0ldMZmwXnGVawBoehQPTE1
dWJFf2AVv6YKAufVTCowCzedhxR4bQo/8O/k0IAslDN1KyNhwDUDk0/AmK8WIPET
9h5sk+3+xSIVY82rSR6pKGipmqBMZ4WbtA6CDrkKqN4YlZX95/MrMtzzSn1K1iEL
vtAxP2Kv2bZfs9ze1mhr29xmvezqf1RobHvjKI7EOFQ2m9F5OLwIcK2y+lt3vd6Z
130Msc57bN71eLfuAUJWW/pg0IH66vBBLbVvC3HlpQbRAjvOb/d9ch5apO9eFl6Y
eYtNcAaXBT3NTbdfJiKXmN0HQ/f24L48efqKO1tHHVE7p5WnbBIP9qnnyRuXrCd7
O65adkDQIt2kyBnWMp9GreWoM1otzu/ltbRWa7NPOaUbFLqj7jEEBYmUSJU3w6kH
7ygkwBnRVGQTpjJaXqbMHtMgM9bGYfNSAYqAvhsGd4oZom1wTaF+9CopFbe5iUvO
4ZX4i4q4AQptFvLzZTdMn+N6F8J1vjHUMZldD5oXylSbRm7CxPDhURcAWBxmFzEV
yE69hTduiGfLTLVw3+RsyOyOMCIrPTAYaab2g9oYVRBpamNB7T9unaNxBd8bNEdU
7mgCMPVcfmOwki12QMYN8xY0B9hB6IUKVtL/EuXCwJAlV4FIdJ9nBO6QY2xsT1+9
laAL5BpAW3VJI1slymRPJ8Vjtf6pfdbw6noWluLCdW4txJQqKbwnjja4Kki56/4k
`protect END_PROTECTED
