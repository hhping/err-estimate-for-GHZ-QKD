`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xeqjwsVXI3QOqS1GethyaY7/Ilklv21WkWzsLaAzc458KmzgoH3rPlMKii+IYLB1
nB8XfckxIgcWZb6kaTJDuzRnVRprkqfyCQYoUtaJURplFQYXoBrNNo9mLbcOnw/w
i0lesDhklRchcF89HOXZlRbrcf8QvMvw908QaQ46+tWtl+vVwm5YBY/E5ysX8JRA
m7LXlqiN1F7ufTzhN0ALPhMlg41Ym076GKnpRKWZ3VeGBDOUqBt0PvmtjJs7sxp5
Nq6eVmn9A9qjvLO1sRDqLgHA2W8zoR3HSzEzRsZSBht8ESMUoue1k9HKqHlC67Id
67xsDoRejLFmwBEtUQb63jTxQBbaE3k5l4Ns93vdT6LKOlj9jDwgHFaB4/p6252h
8OfX+Pn7vJOj4IxEdxTtEuU6muOgpym39XXmtJB2BruD4outmfOPNGwFyJB7LueW
rh4q4pY5iO+jSkICFLUmeOtgQl7p6rYNPPGTliSU27eqpbYPKv6OO/S2aKPmwTsJ
jGGadGBJTAmTLbSybKQoiWboReMDDI8VzW1R/DqNp29QshNXvRxoUmcI/HgM/FbG
yr/tuX6B4pyi+jckDTUZ3/Olv6VdDYQy4GDQeUSDL6ucd0mh+EMbYCZ3yddO4f4n
l9Xu2jwLCQ9j8brHG4NtQjwv1zzvSEpS22CtaSt4btGKM0twmszNeUGHezf/XMiJ
OswRNXBblmW55nwcQSjF4micRuzByuDZFAumNxVrxtNc6S4HWmJ3ApOae5l6BAhM
U33elxv+oiuV9UN/KKHRbw1ospXIg7jbkee6SUS8Cv9WjSPqQ5qKHxocDtQVLzVA
UURJVabB8S3ChSaHux8ImJUt2eLukKvTFAQlf2kGOLbo6CsMaA+ELbPaB6l/YIDJ
vRuvwcSjHkDQ8RLqyZN00BitDkRB/H/QlXIOdxbaqZpgl6EA6xr9DOn6jdtAcb59
AboXxGgs+b/jj8V2SWsqL+Qe0j5s7yE8geuryibfH+5k93gsgRD4d8CC5urBfGAK
Vs3qIfb8Zx27BwtJOff9vw==
`protect END_PROTECTED
