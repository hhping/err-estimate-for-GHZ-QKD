`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b/TsEl4lTBDFSRffvxxBfx2JkqRjEYsm7Uf2F+hAmOhT65KTLfQFhYkW4/6cFM7H
rcrVxu5LlWP2kk7179b7vdWKgH3wP4CC0UaLghvqC/RyBOI+wnTu+b7cTzEtCAdU
Sn5ZyJimzfRMQp12Fh53XWMmB/qSaUDFUg5mHXgmys6dJzGooO37XNguECOBCxZH
5zt2z1tFyCN0Y0HHWDoInT22LMFLad6mwQX3Px9pI5mHUXtbdh/XhTXCAxkD5cHe
HrpByXEkhH7+FlshsvCO11l6Rlb5788j17U/tgQkOSKzJfSzKlpS2BWEqcCQATuY
xHmwtkCiUbW9C4xcwR1oAVNpQ01g6gSidK9irLQX1Uf+NHsQmnsg5Kbi19wDBKdJ
CTPd2pcSBIAbZmY+2HoXjM3AMu3DutM0OwrqZeJLNgqgkcuYuUnZKyX0aB5LcvP6
sPMarDbVgnu8aikpSsJpHuj7hHfz0nLF3C21NiyP87VJw7rt+73kvAP50v5ESkQf
cOfXCqha4dJmsFuAfWt9QnR8nQkxfv4WzAyfSk9sGCMfJEDc9SvMFnftZd7+aR4l
Ot7pA8N3AOMWmVg7LYl0ByMsnTr2VsMF2oGR8RcpR8uE0qz5kodhsSbX6taadj80
XBx1VeofQp3NPLi9vWKOPvd+CODz09J5we32fpgg/9DNYCzER3GRWeyNFagPxoEn
bwyKCD65Og6SATyTAST+km6bqc9eTgX9TgQrKSzU7bEgXSChjWR/oaO8jXFFxaGF
Hd6PwNPkhdISxlCKVlULinD78PAo4/2vOaUV+aI/Sjnrx3cmaCxqmXga8hCCSKFq
rtgvl5GE0E/GdXPCSZmUpwOCPYtbUKqqz79eGDNsSh9xGeI7E9gS1qQBUgCzz/CX
mMFm6OXJO3mreLVzThVrL1cvOAgnqmR+7z7apaniw98ZDwdrQDSypoCdjcm8GP3M
UNgEccGHF0xVH6RLXz2x16j6Y84BEe96O+hNVSBZ6GaNB1h00y4aFblgsbnGm/2k
vESPcJxEc/YV5HmxXVLcWnxzdKZbckVFtFFlqsf6YeHD4gFY8VYWUrOm6rMiJhjo
46yNGA/iPyTJHIOjE0EYsN0JJbfAhKu5uO3ECjF4WgKNT+Q4GgHsOIocHp/KV/M1
6oLzp//5Y6KUWIW4cIe483LOujLUmlW7AMja3QRj/wQl78btHud9VlCIUnXjRgun
SrwkdDytB6FsAkPgfJ2gUkmZF2NpdBoZj1AqqOb80rpZzZyrbzLrLka4k/A7VbG9
C7ummnDxSFUqp8m7RtF4BHvyN6Ns1fPP8bQgHKmiRWa2u5BGQr48A8hyzUJZ5bLi
2k1meqpWsiaMdWr9Cd7swvFoINFsLAtfaUUqBOrIxlAXkm+5jl78FPJwLLiGFUAc
t9JpbK4XCLYOOQsidkINC4hi4I3LWnkqq1/F+8oBqEZ6M3JqDVYmuKGRkuAzyS8G
Vepg2DgNzdHNNBxOD2ldlTgHszWYEFfxrfb5MLAaClTOpZYB1FhDoszNf+I5MNlS
u2qd88Rm6XV5C0Sp/TJsgPDE8+SAhpc3NHCMzbTx8RkLZD0k90WonOdv4+g6T81n
BG9hY4ptFrrimxiPteljqm+22tl2qNQ+xWlLh90UoocOSCybuCFQMf1KOF9f2lR9
8dsngPZU5sSsOu4FZaPyiVJ8PXN5rgcgLFNzMWmPmJMUczak/uJ556qqTMAdR45G
RKL2Oz5IndpPU7DQ7MgX/d0Ma7VXi72el3qY/1J+rMBsYHc9fcwpiwR2qXpEAFSP
M1l662txByi0M85gupNxC17u8SrUiCv/CIf/Jmg5hwaqJmkDxw4tfUqckxsPQLNb
gLfUmsbdZzzIBvxyfbo+qs0fkw00I3umIYyAsJK1BXR/xmWbjWFJ+EItoIVAE+GJ
oCNvM2v67qvs0lkj7AKSv58ngyhosWYFeQjHwZcKKgH9NK0oA53Rrgeak6NUWm+r
0s7GS6wmFW1IL4HBMsfWOgjI+gZIPXwOq69EzL1s30bkgajI6LIe6p7rZt65ioXa
lIXQNnVMe0OYty4sjqEYEgR0+oRSzpS9g6G5NUtR3vO4TlT4blm0PdH6TWSSkvwq
QKcx89vPISy4NkkzzrlTTWsosnqoxP3IFMrMQy+4ZjdwKJjxCUN03JTF/X9a87a+
fAb5bv8rk7ehm9hm6maPXeWC0jT9qYVqCN2WPLVx2pr5CxJTjRRmF4eBXM+pIx5i
40fuuSFA9QozPg3ryJ+Ht9JzwZHmk7zl1GGP+cMShzZHxe/y/93h8JfihRpV3JoB
MMng24hd5OlQmbeCbs+4BYDASs2wDMWO8VHTXOneiT8ZJlcnVepADQmN3k0J0rDP
EWIjjUaaNmxGvUM1bXy4crHn4dTipAEgEUM0YgelFA+HQrSAqsMGk97OQMdmJfo6
1Cdzhj9J/f9pntk750R5DMGrc+dHhXkSq4QiWxQ6rsgZSCme1iniyJAUFfH5zhvO
MvrGpqffsK0hmaYj96Xoa8RklbPilre1WuSF9d/Dxp2j+Ef10GTzpeuRkdbjRmXo
+PXLoD1qIV/W5xtGi3CtV7igIlMcUcwwmFqgXxrk6lcEd6wWNd4Lb3Of/FKiyJJk
CE5qqcqXYepTRBB3sfwV6u08mYj5SvayGbdSjPwtm77JCHEZvn6Jhc4i8t3fHNBf
L8Or8dRWl8gHAW6cENVAHXBiM8mrdg9vOMyhPYaSvOAEtWRoDHmKjyxmVZYymF8S
MEt9lhnyauNQBrS2SVoSqpLSZwlkRLxAURvyjyVnajnp8DhDyPOfFnYBHpi1NCwV
J1vskhA69rAupUXur/Jd2UHaTDJbSe9n/WdI+X7qVlbtOWxCEHN3WyCtw9C9vJu+
cVKw46RuvBkbAUktfUKoQkM71z/KtSvJjqhsf5U3y2n/5C9rj3Fq9KHiWDdebKZD
qpYGlZ98NEmkfB4GPLQxaaSIyKtxc5UrZ+djwi0fHPOiK5mgPZG5hDxOXgNDP9mo
S5A09hkLAKdvFeC0E8oIZLSwqz28l+c9LlI3V0s/jOlyn2cSQDxzDTKUfPm3ztc8
RRRstyuydJxJ6wKAqujJn6JCcuz9vIi45lK2B/S2r4QAGjYObEpwZcoC6PnJ0s1N
PakWEKhhQ+RAP+Pw5MXJEljisFlrHM+eGPZ/hyz6FzS1QiM/kLrKM4G+xbiNTD7i
66vg93yQWNEXMR1JfDiiy8VHCPxfNX5jLtX+g24Zqb5nT3GEhRPXUZhiLZppNZIj
iKc1M93ZhlCJL5SPUIa+ItHDxgDhB4xTI+xeXO6uBGWwX+UxwrMl+yNiEzekGdZ6
tLJ1uGWbl7iugnMIEYzXSCS9Usq92ekhVgYgrXC8nuDgD149brloxfgD9hbddbXc
uy7MlhOUsdm6Z8snBWlSTJU578Z45i4QhiLZmsZu7M+PsR1nxeX7/w3pFcEVfyl3
63BGfAKqxfATaUA7n2okMcfqEWniNtgsPWxSjds3clmfyYbUf5h8LasLSVZFyt0n
FU/ig80sabw78mu5cxGDVzmnVmo3GDUmDGsZjuW9458WD9u8wPljfS69zIF/VinX
A/VLSAM1asWk+0lIGaCsS8h27xh823UlBPKcxTaObpXLwJg/6mebN+spB0mbq7R7
kreQoGUuQzUGD6a73eQEzdCCUeFgCj3NAhrdzATiJzVjjDdpRQ0iu2YWZSIMvSjT
q/42djwC3amT9wIeMGNJq6Kz/8yz9yeXN/vo4mzRdIcCmOEYrA/lj4xK7BpJGrGq
HjrRnIKYCxLKBGCcf/2VxdCuC73cl865KUjw0X0pxHPona3wFMbHvvJTm5IwgRO1
CzihZyVun58MUnAynQ/fxQ==
`protect END_PROTECTED
