`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7+/vYiGkXYjbghvULk5qaf9mElHHT8CnlXUuuSuRFdsVU39NoZp2HrINcu7qAIE8
WGd0EjItv31w5luPF+meH1vja/kgGwypH8WQMvMvUmiU5wiTmjvWilzJ72sqsV+/
jqX3rzdCFlCpesiMaih5J95E/VRb6mV78K8ID21ZY8hb0s3Y+GimovA58JWkmGh6
EFUpQ7ws5dAwhYS1fIgcgQenmLnODqtFSWl6nV31F1+M2zVM98IgZRE+NFCwxPl2
Lync5DHA63HNTNjTh13Mnm7jj7t4WgIKh/NzfV2NQsk3q2Eu7ey8ZNdO2lsu7EFU
Xf2q/VXkhmz2MZ+XkZt7v+BKBo4GtI3a6xzwfTP8xxBF9qeEHnBGTEzaIqLEqQzG
6P1E2IPOlrKOtuQIhwlz7IulwD4hA0jbPDygM2oCA7Oubb2iCkBCk/fapmDo+/3j
jPL7+Dqngem7HcX8JuEEpnp/BQzxLG7IVViJJYRJq6YFRXJVxamjGFBdmR0wl4Ik
8y46/RA6xVY3myd/7oB2qXT9mNbVRBxLxrslLi7l1OzwbqmTbv6to5oLczdVOBWr
9WyLT5DGgC/0IvOytg9sRkZDKh6V+0q0fLDJXhxEOFEJHqtUKA8EnDWyVhT8dTl0
nA/3XIugZvk7ksv6eetEmODJVsPzokI06ENhJWvV6qa2K5ngt5TrrnWVa0VcSvoY
dZxmdv615k0tkOF2XS3HsetYOFkn4UuouG7lGeS6ET24UpEGPQmNu/RTX/kKkDQG
ZOFp+3adDTxWXwFqZXkq08/gbM8UlXNMPTXoBGaW70u/3VjQubKUmWrPEum1kfkT
9FoKuH1/+IedXfjaA4ykAM0FIyd5lTgL3zuLKl9deYxK9oD17OBKZarjBVesF5Je
Nb9KZNIgx5lDGvl78iySf7CNAhiqeuWeE7E5dM+ZlYkZxryaXFJMCBQpZtHV7bcu
BlhMZN5FjVaZTQ/m3wooamQf9OT+khe28YaPMgVRBKI=
`protect END_PROTECTED
