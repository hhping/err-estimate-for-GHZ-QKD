`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2pwtCYDP4ArX4V8KeM7kd+tyXKNbXzpVHguXAVAu+aNG/At8VQjYmDZzGDOz5CDA
71ZwGCMiRDEWCapH58QJ0P+zSn+mUQDAmu+2r1VnqSvvSqyLiWOcw61pmSwqUgUA
z4gSeHONgrjSVY1uZAAUxheNn5tV8jUSNlSUfsTvHDNbfbUZe76SewU+Q558bdvN
k0L+feHSa1qtzFJrUGWxNpgHHeiKcM6UE9qoDNkWvTNv4QyOl4gHU+lW9a8vFt2y
2zD1EP/WtrExelsxHOo3ywJ2t0Wh7Bjsspqwkd8VC2dLIX6UANJaZOwdhWFSOT72
EuXYUkpb9eI/hl7Pc3gRUl1N5aBedhvuTSgvXgSTbNc1tFvrzO9XXyMmA7q4DNSZ
iyD5cOgRGzwgDSF1BRrnCM00rmC+cvxlMDJE4GXZXBRjau4GY0XGCoVV53LyeSVb
W8e/pTdNHpdi88/xC5vZgK4RgG37xVVeX9OEKTxdvjtIYPWc8+vPvGKnGh9fcXDd
`protect END_PROTECTED
