`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5z8zP92X7aKpuDf8CGbvLM6rWM75Z6h3739Olr1UI9TAGNo9ytrXSPCEN3Y26RXY
8vh6XbOEFJwOkoTiPhOMXESXnO6aW3rrB5OFIwfp5vxcA3/70NjGfiNY9sayOVpY
gNGLCYVky9VvQxBgy3uoyrsBIlLR3t/9FUEjKWPM5Tdpj5R9nmRHEkvv3lHT8bqf
2sP07/Iurn4bC5QnCjDAkUlau37woIFBcPD91ZXESeWeWdY6H7rBq8fyJuyBcqo0
Mj9E69DS0txVgURSmnXwMAuc54b2HW9Qtkwdu8L+bmjvusMZYhAstRxs1fMZvlvx
W5dfH0DWP7S2NG4lI8S9GwsrtUvEyVhG30HxzWr2nhI=
`protect END_PROTECTED
