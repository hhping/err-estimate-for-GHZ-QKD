`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xbwnKVLtbN0Vs2KZa7oYeNhmfvMj9M2PouqnHuY3aQWwg6NkeqN37ZgILdwW9tEr
KAzEL6QXonJjNIwe92Z7eGeS7RBVImXijWzuOf8ACY8n8rdq5+Ri5uLJbsqDMCsv
KwfexijFCQQXBcz1qtFCdhGWR+yoVVUVDcXUKtPGI3eavbqEarq5rppl0kc1fYaH
1kgtGVwkexSc77EQwRY19aWPr4yUlczL1M+7mfbsnggjUox42YZJKd0uYWxGtaG0
xGC3pjvbWLmWkznaUv28cjjrBAyHahv9hx8FFp+hc2UIYQZU+Ja0RswV48l3GS7L
37rf3/mPwqJkRjolKP4IktPtXKd59fkosgb1E8xk31HRAS8zAUZwRXeIT3+15wlM
hUh50106UDLiPTQlA9UhmOOSEs+83AE68PaXhHm1pKl2XL/i9hgDcT0Fz4CPBegi
C9W7Qde0yrW46r08BA9/fxX5h2NhuKVfuNlfnUThcgts45vYhb0tSyEmllTg4hxS
1RF8l9q+jImU5vHAnt9DEJ6YEF22iPt4qwQxaV+5o2FN0KawjvnQRLf5iqc2JNS4
P3K8/wJBfv1WKxVMc5/s16p4DtnAJyzCXi/VxFA4QjI+223EjrXs5II5AGzHfd8F
7/BLwQU9Z7C3dxmecnJ/qKqKHSpCswknyocJIHLBVOBl65KVhaFa7/Xgie6MPHnk
MzBzYyXCfswRpd6fdwCJtmwukkcaJ2nIzDGRVjglv0+VwICtwxZwE7uwDYCeG95E
4jrErJZRywhlfVeuPm+A5ZjkXcPctDz3i6s67gElWmLgb7PQA/jq2R5YURrro1PA
heoRZN9QMmdu4cDrouyX2QmQ2QrfzKM3m7lZVXOomJfBKibRcjiVu3LJ3pWlE8nH
reNZX0C1qhW2+XttcyLSj1CUgYGkvQnZbiV0CrMw21aGJsFd+E3YlSe1AGePcI/9
fr8sC4Nq/L+n6cf4pYgCEatA5aKqLEesH5LfW1zPQNyCBpdrFDbw1yhgQdUZL4gT
9nWOdKuvHv/nsrWKC5Zj3jSlnumbXizljuilsWwva0/2oCaatukPVH9bPRbWBJ3a
kg/Ld1srEUhR4FzAbboGYszfkgNTax1XJhZzRhNu/r02/U7ilksfcsLvbElWBYa9
CtHLkg0OfPhrIIQHd3PdrDK1XLJstpca5UeR2MnC/2i5KPNzxYqoZTXTZphYgcQ7
9V6C1PHeBxGa4yXB+oNgLSg5MtgmdkcTV5YW452vluvXEDnYepLBHvofbYLV9fld
3vr4Q08oFcDrM88Dnkn5ab6t1eciQ2OQSgDWYHLx5V5BQr/bb2bKhDlYwu2MHQQm
Sb2Ve7unPp8I+VkDV4m4hZuixHuk2DU4eY76D+KQcpdV0j3akD77RG1xjJxKJMZ0
+a2qLBoFIEDl/boLOuNv/L16sCjCPNGkp233WBofgVVavfZ4VdUjH1/us9P+eeLT
h+88y4JmcXlhgcqMLTSAiiP7JcSp3K40EtT4Oqz0YrMpcNZLJFAJ+fxj5Nlj0srD
bdJzesPEYA8LAj6TbY9e97aSMWz4n5DFR0KVam9OzHxABxkag3RFCsoC5CTP4XSi
Luboiy51Bae+VLDit5blYVLlfJ3eTjFEohE0NQJpXFMvQbSJ8JdgxOaII8CN7f71
fKxQNMb7nDLgOOuNuR5sArabMFfnykHx90VBdWtoo5TjLAceI5VclZ6MTMy/fFCT
1ghlagaHPxLGuPHLD3JJp3zupZA8vqrEacKxzQnx8YJvyY2OPd5N4PkMV9haGaU5
sW1ybpxDQW9eHukO3lHpAwkxU78k5bMvBtBXlD76PIUUf70mYp1ypQ4piJ79c9iw
kmK2dG7H63sWD2uiFUcGdoELp6PXz5Mw/5KbUGtyO8YwPwPzW8JO15tE49jiZ7BG
nhjo0IdKyg1xj2i5aQ9SPHCFnBfYZn+X1FROfWCHKUtV0Q6y9cL+zRrfEByv3n0w
OfViuLcX8AQUIq5+H0LvACXhag3SQFWQDV9Ulv1KE5HH6h4zesA/tMsys1SMLOyT
ubN7X1z1E0SvLOzt84qLmZU8Ie2Le8ghkqoexNC9o+DmQ/A+5h3BzsktiQ1/NHBO
IDBJTidGQv4bqF1Lcb3IzM6XNGjvNfdNyIjYlhIRzcns2AI+i5eL3QffLlQt0nOY
tZc3AdVWIHp50e7jrz/0Ssu0vk4lHjCFSXCKvi98KEY6Oua8ea02CcS6vvveNhGj
F5q/iLwjo3AZQDNotfzg6wMb3wgaNA1IS9Bfq/3iP7SNxVnntAo15LjTll44LbC8
WC6pQ/fKkc5DYc2e2+avdUqeTwIc9OwrG+8NWNe743JQqCc/C5kBT7WYWwUNXPDc
p9lztUH18YmpWpxC6GKbtjnZjC10hTvmomXJUnHpD4D2rZzoa+sUQlFASSeOvEOQ
4mBnbw7Th7qI4Ap68cAcZH/yv5IIcfRMCRo0kkySdi17ilGLyj/HDZ6CORb6Oywz
XhnGQ61rDvcW4MsBB9hCHeKnkUSMMzE3Kn6Z7Ltgpu6b7KbXIq/TI7MYtBzZ9yOD
HnGkhNrbzdT1V7ISCzat/762MreZKcEixrfrpudeQPLflLOaN0CTCc7ltHgaRYXw
uKG1WW5MNYelJq+NkjwuBCWlW09XLU4PqFUW5E8ci4q/EJq8or2/kXLTF6k2BoX0
JgENb0U6dFpdEUZXf25InDyS92YiSmYa2i4saesRkytq50NC9mBE+5xzTZj8bsYI
GEbbMVyITtMWOlH0KiBkYkEnIVUjc6jSCS8YczjoTJqUQl8ZejBZdN0csijwskl/
H8ufR3siT6fJPVRlFfqFIwkC3yRi2cWFyGMYXJMPKZqKhK0L421UhdMGlL6CyLkg
XHSYmNiSb7pojNEr1WRDcy47w9AepD7Zo4aCGl1nPwIrkuIOQMzXJSmsAFOcOsbl
qpVPMUwDfKr1bCf5knTOT4rRFJICUezW3yrYJjyF2R2zqga1mqqpGsVZzF7MLIef
nBbrp4sQrFanhbW2ZpnqxsFYBxBnNvwTeSj1FQ/eP9UKhentbxMhl1LA9IE7ZKcP
qQl8OLzi8hXd0ZAWRC4i5n7KpPvIOjjXQSOMYRsSwmJILskEGA31B4hkEWwD5ccl
IwZP96fFgPYtDhDEMYlq00H7j0/1Y67Ap4SPeHDGij0NmfObU3bo6/vQOf6M4FFT
At5DvLO1vsAH8B//H/Wos0kqSgaQEIQp6+cLo2Zkue8NpCpsb1RJJBXvKiC5TkOm
uqJHm2/saM5kfdNvEa1YEl/BKmy4KwWDC+Hlnvtt0U2n0YdQ9HEEQqVQZLql/5NI
XtHnuGjipwmgqUA3j9wwc5xYgWLfbhlhSMwZ+87B+DIS0xJ72a/pHYKHc9kmKliu
OtbsPrLbqu87QoHr2EoFnI9PGVGSWb6yf1XW6dhRopCLN6W8PRn3Sew4Qrn/nEFn
Htj6wXZckF+6oOJg15Xw4TCEP1wWjiD6dnS4xLEUb+xlLnZrUYxW4sTXEaJL0/Ar
08vlLXOsF/JEUZw5jnzHR2UWUkmr9lqBDKELbhbQr/UbNW+zv+YuDcPS3JdZwEKu
1PmqguEmfGmwE5f1nvnCiPdnI9Fc9pJNskTuJihaPzGL0WNQq/rbP1K+QNJ5LmlV
R497yROOxPmbuFO7MjHgsxkjkgYEUQ1az5xryZ/jVjF/XayQsabZ2zYO/oG6bFhc
cTbXn5IbJD+1/fbBbPFYc8vcigifgeuFAtFztnkV77M/aAwv0JHHyrv9FEno9x6A
7rJ7ATmu+QTXIXMjT7ssTYzidDp76Wv7lRvTVNNelvNsBzUjBZ+ktHD9EzqAmgWI
t7wYYDXGRQNZx9f/e+3CzzJgwPt7Gvxki/sdQi7pnbIOIVHuBeh7rND/5MJFKLIM
Z8qnhch8jaNSWuiEMOqQRXCqw65lCu2nWqDTMVZhRDQZL5fPeBhkBJkYW7MQ0pD6
IsbYCWpIcMFXVh1fs+LoSjhIPyugK987Mr1e5723mKC/1TmGLRP1O/c5c9Qh7x19
GenBlUSpaeAhUYKKjIlzdv3ANKv3Ilh1vAw2TUcIiPbVmkWUpc2X1xaVWmuu5+Sb
lci1Gy12J/PcQ0meyXdMH/QcnfnrFuCbPbMfg7ofkdE48L3F4pz+OVLos75wVzgR
WfyVRRnHKBWMyEQP4Y0uuCLM/zdrFMvt8KMn+FdFJ7WLxJaidI4k0qfXh/62dF3P
546qegldPC/UodXYCL41RULVNoZII+ziJASGzsOe0/VeDADfQ0wAj+KOr5h8BkNX
/V7kUHWUwXsuGgnZowGDrRtGsW3a6Ljyp7tzJFyPtAgRCWe8tNLBa2h/r8b54fWo
MuWVRHq9KUXiN4OHU86XrXBF6IgMCD4VKNzaDGCUGF0f6vvlcCvvDPh3L23Lo8jB
GKbySJZw4rjWhzcexriqXNjaB80aPkJge4C6AlxiJWrnF1wHtwrlOqi/i1WbWQiw
ee8KA1Qdyk+kikizqPAW6gmSmAxfFJNgMMR1NZYtzwsslfde8lOXaAS27+Cq5Ady
DvzK+Mh2RAL1NuGwkL6YhDk6a7k8kYvEo7JK5xtG5YvCMu5r46UhjOgIIOHGxfTc
Ttcn8WpuYuuFDzICsqI1X+EH5BESncApJIM4rVdg/xGcd/gib9Xc3ITVynGdwzDR
KKuzuoiBDnnLm1M3aGUjtoiw/yhmAHDdMPQjWzjTylpSTsZ56ybnhV0NvZS99Lid
wSxBeY9FUjeCCaCVdxZBnZ9m7f7+II+ULJnu61aOkDIp6xmqo0591kJ5U8aztQC4
lpCUeqbO5Tl/7zgJWYslihh1wMka3OD68gg68N52fmgug4G762rQNvHW68DUULpT
TlzqpRkpOm8ZXPV21HiGvyglBA7wds8oTddXqq+ncd6p5ou2+ADlvQ0htaZ9YQlB
ityJSigYAAexyuYuW1BCkn2rIiqMgbZtVCYTnJK+zVWXZsLjTe3BDXGhU4l8CP38
PXPPk9YnX07cIAGuIwLTvWrCDA9cF7z4mOVjcZ9ozeAIGctBCAgyryjHSncdI/Zx
dkRBN3bvRmYBynK5J9K0fw/hmlS9lMy+VPSrQu3l68flwobNml9UnbpXrw4u1Sn4
CAmOoocCVwezPsCEq2vivnKyimQGGKVMJUKoqA/jCIPhI0osYCUnDiPSvtoLS2R+
x59dlR5iEohPYgxuPvk4cd9GtJvTGj8kBnCYF/LnNfjF1YfWPuC2XfyaQqO0sxap
SbTGrcZC3/cG065PCVB7wKrdxJXy/olicNdTpGPFMP3cMKO5nf1l6lOfRQGvEju1
N45BBAWcscom38I/KPwG1ZG9otk5C8iUyqaNlB2Zxa5zUiE8gZT5cCZyGi6Njbwh
NT+1anlEwZJysdMVGfJFSwbXJLBr1Yz2AQVO3fKjXKr9HYW/yFKOr6JIfyB3EQ6F
+HUj/+BMgqQ4svhDqWWzCeaLv/FrCF9qwAjX5F7V8+idCtWv9yC2d2uWKWZM3fpE
vijEW9GABeBFAYUEZqQVzo91+CAdBpNnXnqoQxZa/3zGzOmxpCgedh5vEG9zzl4v
tps1CYRRUlUgJ6o+nyg1IJSroFvzX+bYLO9vIfinN8PPNcj6Lmf7GInRs0gMsjFg
+YYr8NHZ/YJFB3wmO8K+VXXJFHfE2mKioZoETezVA29AxuZmfwWEb8lrrer9Yt2I
rbjFjZ04J5sFzq3Pj9vjXTLS4nGO+N8mdS4h3za0Ci6XoFUYOwC3ymWhaFZ4W4Zd
xkhVTecv3Fk7AK5qFw9+6nEMbFqmiL89yXFa24zZ8DTBQPLQRZPG1P/dFw1m2+sV
MxUwPw8EdCXAcxDp9vRj7tJUFRIgK6FXENUAYCqwjaL6lz40k/k9sDy1Mmkqbn81
bxY7m1HaSp2an86J/1/zBPlYPEIt7IqRCViO1CWB08Fn39d0xYBDOMr1MxJ19jMh
Um8WY+jlb/QqFxSsvhDZyzg36rOADJAAknf/h0O1lwpnfJIvw2vGsx5Atfb7sbSM
YD2UepeU1psUN4f1dFcXTmtqkHJvzr+TxtxxlQTnBiPC2GPcoW2K6iERk+fHW4bc
YF4JCWRoq2jF8Rsb34hXXi2Qb8cS7QCwPHPM1xydo2ofI7L+HuW+zTR3KCzNAs53
1A4nn53VwbY/bIasf3tqVWLoYb9uvfG/fhS855yGolL6rbdrUvnTlVpbWOkHMN3d
m7nn7g5V7s9TAJuhwOgcB7OMHbVHdEhV+7731vDGENcLDfdpf7Qo4Z7TOJQW2VBf
4hxLOYS2pX4iHNPDgc7yIZgRybhzHWY1rWmrAEWStqFB7a/HzfzV/nLT0u60NPCN
2DQD4Kp0HZR9OeD7LQXoHxep22oRXGVAD7GcbV+ZvXYIxGCDCikDctY3McYMYWCo
YnrSY8Hia25s3g37Ui3C/WPsLxToet+7ErY6sESXexnnn1YSHjjI+uir9kV78/h4
hqHsGKN5HEdKNOwJj91SxjOKZFNdG7tutjmeD6AL81Du0pQJP2+ddYcO9HAYd6FW
TO+RpHkKOLspyTEE+zN596rxyjkmgF8Wa2ARAihMA79MMIhgmOmeas3m/B7Fz/AO
+4kxW/zvxFW17v/B/dceNc/g6QAPVFgdG3w6XmVYJVTlA+fJ0WeTEVt/orDmJLTp
8Gwf6wLDvvAuIY3Wira+nk9bFU2GYiRlHUkO9zGm1t2TdiAn4HJ28XyFWEo87zYs
cRrZ9cpfpv+MaqrkjVHSyUIbSqWmdT6eaPCb9j//+DiMaTTIqUrs5S1y8RH7MBB0
eD+6wze10/8Ied9Br8k6jbqnearnP5oP3z2HgdyEnTUmsF8Bk1AtOI0cuJhdmTuK
vTfoiMTMqmfMIp6dqrR/NCm+/kPIqXON9sSJl9WtHReuAb+SFtBrXZU6Z42Mlvq+
Zwp4oQO0kILPk1MzUtDi+2AKE1MbZeetP+wnNYHPYhoFolZyyWccGz7d1WVqEbz+
iBpRok5yhtS6lNY9fuvlKp2ziYA3RzOfm8HAcOhfShLSt9HvNbn4aWkhtVF5cZ53
VZcWDvj5NoJUfBs6f94pg+Gg61k6IMZf99MvfGujon6fYp+Z+uJnGtuv5D6zj1oq
6ovlwiE6SmxgILRHuRNbsDyyjgTfSX9dQehhVvaqAl5JwTHJuGtiUl6Y+ne2Kjy3
uMJI+7V+HKEPYdEauqCnLg3txOgOxC0zyMpWOT8aXVuKhdvwnr7+5SspI9FFhrlE
tUe3Ks9KP2GGxT/hCWYk366h1kYxUKOnIcWaAcYoN8l3wY9yBRl7EsErR4Igf5T7
9z98EytQKWMzKQY0veVEyZbrzIFK1IsRgVgOfluwFKnaC20egXcsAXORP5kbtuCv
mzFw1Yey5c6rgyd4WqiOKLfpAWtw+p8kqEHw3Cc3ECS0auNZi/+abPmEwgdMkSDl
8q+QyA4/Zrm8QUtuvBI0qGTTclcNisVjwmK7et6driAz8pdFHjAjZgPpFL+OL/0s
yCcyGY9bousy4d0U5wKxNB3RQ8jHeHkYRlQBp3b1XUhce8lsDi4eratsEH71hrdy
1IK6m5huw+BfOEwVG4DNX7Eb4cRq76zQb2TdO6GCz/wGjCy8Q0fjoGXKWdpsAUE0
TDDLVo5PjjJBfTDCBdqSo3PQdWYJE45rzGvpzif/867ZsK8hSjqfr6JdOhkjjmVt
i2ZhXntCU88/syrxika+19kLXxkMzY7oZ+qaSxxh019BhRQuPYCdp19MQ6ANNErE
NCFy3bU2k/jfFRz5tqtMlTEG/xg8IiOxXjYiN04CuXfPfjXC6Svc5iFol2IPV0o1
6pd1jD3Nngq/rfAJtbY4s9HjQegUE4w3EK9YTi1fGPoMYM1HO/zfLAImxE56GMoB
dKQSO4no+E1oK5FoqALNUYYyf/H/vLONiLiEhEnDubzYLzib+6TWxrcfEljrCpaO
uXZeF0uGEQRYNCeI22GKQ1cRcr4yIqaRhGuvLsQbTfXoRstfbSl2FRv+Cpx2n789
DtlAXdWWkx+GL4YpX/1lhf0w9xVyksm/PXa6/0AkejCAP0UHZ6ARdyi6NF3tcfhS
aUxoQZB1CLH3rLc4eu1KcEr0Y3Sj7O4WWjJANEkYuK1qWhxJDIts1LxNIkm4+0W6
BMe+E53LQmjWG6mkncZ+P49N6dVjQV0RMeX7turepDTfYHMDvOBLMRG0QjUWwb84
Um9pvAPhUfhV04FUBMoJFSuscudoBD0PxUX9HLF/NYmFkI1J3i8xtuUZexs90UEg
w/n77Rj/N6J4QB/DG6PTB2mRJmd9QgFFQKyiNf7v2iq9qay7yWhQlO79abfsEE1g
ENY52vzGDY0YAcmcTSIC9k2ev3VdYFpbwN/PsfuHBbDT1t0XSfT9/tuymXe4LMG/
zvDTulCRIDsdKSl5J1b1M2ntlbQqTnj682pgk/XkTqcFTqvqcFE7IgVjtBuASl+/
YFoazmU70asG5vG6MCJRU2euv9sJWUB4AGKFmLBpBEjsHSiMKqRyKn2bWMSwPUaE
iWH0cksEO9mGKjEeCydrMT68/6zrTgZUJwiQ20aWOGJ0a7arm9+oxg4E6P0t/2Lx
BdZ0ny6OsPUv/hLNYzobLXQcG7/klpnW1ag0OQbXT5WWilsvwq9cOxdKsXwBtF4R
u6SU6APtvx87p1oNleLHNxBD5gCLGPs8SEYCjnkx322oDiOyn59JLPuwLEu31Ty4
fdPOABfvHdGXmBejd4rAjCWa1CzZJbEQqizc9YkGShie5D8BHT2PM1oAmQrviOlh
+kRhaktyiJeNWDRUnsmKXl1e0gxmp77z8nvOd0JERtrRuck9Y1VaIabkVqA44wH+
5sNqOS7jrhUo5M2IVlR22XfQi14AVuss1DVTGBiHGoVronhzPd3uVk2bhCx+CUSE
tQYcc1GyK1yjDkIYBS0isedFS1yVDLNWr9u2CuEH4gMmskKzrKZLyXrfyKi5if9V
HVgYZwpOqe8DD87eQYzYLD7LAFxafiebK5xI449bu6FAwhqENgvXXUuM7mEdrLa8
ikS2kd0ukTyWBgmR6NmI2h1JgkVtxlR2LG4jklPTBmo6hF7Lxe3ONXid630aWpQ7
zvJnN/kEn9BkkQIC0C0N+J8F7IXADK8VepZmnBwLZQOJPQQ3p/BTAC4RAcVkSmIz
s0PrNq3i0MjDNkY/+7Ck3jg/cqH412M0EZXFglH/jcMreLffKHNlr64LmYZaVxeO
gowR72ItpDIjb09GukR1WmpbniS4Qb5ikecKjn3sudGCE9hJVaHwXYTB6AjB6SoB
kpobMItoP7UyrxJlY4R+Xs6tENMIQ6/8lijAoghw7E2SciOlvAhHS1Pv+Zr65tM9
F9WAncUq81ZJ5jRS/enMv+A+CQeFLXa+oRmOvpgwaU+BOlRt8RSm8OEas3nZQKv+
N6vjogVdq3TLgxt6A/GaFkzmVBDnDId0k5Eq8RbEu/bP8lF5ji/cbTLjw0E/7QE1
t5k6z34cQsr0lL9Ls0QiNEsNhPPni3Bn8CSBKoJdK9t9X8jt8qBBX9+O0vBRXrpG
szuDtZGuVTsz8byUykEGsri2yAvi9qdC6UTNpzZLFTshh4336z3yutnP4jk0k8Rb
UkY6L9HbF6SUZS0wv6w1U083qywrV5+WpHbSBXfGYML7qR1YL2dQAQ+9TyZiEzZC
e+r3XTJj8b2gw8bjTjpJptUtHUDbu5geGvYyMGU95McSWQAZ6D2WjjkcCFavxReA
Pt6Zu+9VcucdyAvGSKkszJGMg/MFqm4TPmHIyBVV3T+zbm0aoZ7hu1teUNkoNHwG
N8yCA19uZuGcN8VSu02tXJtlmdZpCzgtxKfrchaiU3aTOJJfpCkweQNO+zMBpxny
L6DxH5aiO1Y6KZnC/BU0DBNY9z3u0kIAzlAjfShZJ8pf2TVyHVxtyhowlcdSEmTD
X+NUDCFMR57vSF9Dx4Ta0qC6DFmZ0VbWYWNIUVPJ/USOdGoVYgVvFvGBVkLR6qL+
mQHWs1SMGTW22vSliWqkaszedoJArYp3XI2OjcvFlEiwT0CKtVFQoKvfNTY7n2hL
HbdRFKNmV0B34wbUGbJam0f2qRlXVdlBq/8hYprJ4FhKk1+R0C0JX354Ex/vytv7
okv4BQaukFWDPRpHshgONPwz1dJ5Q2fN2VFTZXaDfmv4O3hWb+kFrTAZQlg0b2jL
cic7OIDIiicdSNN6L3b7bXCQvP3e7n2eP/1xPZfDYFfkh3QGelTU6tSF4Kx1CzUH
t7ewUItfpvTSBYO2YyTeOYHBoPZMlBif+McURRSVUI6YC8Z7n25CNydbTiJqXUdQ
S/LXFTxdzjob3UtjX7DoHBMDWKo+twGgBdG06w2gWV2pCjLmXaIgnZb/qt0dNcea
TYfPWRjzYeCBfYrCWs7+a/p86O7/Kuqt7zzS/3x3KllyDpKRGN87MIRSjUlnEajm
iiZZQA8+Q6q3nRXnYUlbIKbS4NA+sTqVrsm2p5sUSNODHuGci/pCZiSd33XzvK2X
faIyR41ASmJ3tCO8M0elujTdxBkOe+uXJM0VbVF2Znebv9w/Ba5ANfrHjLMsxD7f
tb68/OhKAwaPLA7rmhBeuunlJNY6sC0nLL9x2uZDXIQmD4iwBHKhsguBVD0Z8DgU
bWve0AC3REmOP5xf6c3WRq/yIOK1klAb9r7QDJASIl5Cl8+cx6TNlhJHedrAcgJT
gPP1cTvb1L7aFJi9SAaZBlRbyO0XvD30n6ta+bB+g7stbauqjdAWIYOLNKn5MJh7
Yu42/UM+2yVtGayMDxYSxQhey/IuSLDFIaw7f6T8c9iJyLz+7MYMJHrpdfvzyIkb
LbY+LvRfqfnab1hF29cZYw/zU4xBSlv4fvfHIY+NiMNSWgnroXZC8FgQEz5E0c7L
xKImHwO9kLdOHbX7ZpLpU7TzTb/Ns0MFaEwvSggJanQvjgwjbWdbYD/GlMrhb3Bb
VjyYJxn+ww58CpToPPWe3w39z/dAW3hSj39zA7tApe5SguNUmIA5Z2w2IkjmJUEV
5Y0kqvnlKNK06lV0fZ4dTv5n0a/fspDsofCbH5BVEK82HzrIOkam449lcmyF9u5H
zcMCKh+fJTmzi34CVirFMYKjf7KNdSQB25CrPUe305Qdkhdwoi0rDJwTpVQtZnn+
dsAXtliWZPSILw+n2rKEjkd0rG5M4S5wgYfaECb7R/sIMXffYvQcJefUjWaiw069
z7b9NgUeXR1jMIms0BvZolLRZ5BULCC71fGhmPQU9teRlxVt8CC5KpMZAMgITv+a
K1bo9GaoA9VQv+OX0YHVVUEyCZR0GgkB6uBGGPhds0l2oEWCzy2jj7E4oW9+HTsl
K3nSwYAeSegtP4FOV2kPB/A2xGnVejKCeb80YTxBgGbkeEqi7P8b07+VZLM5Kozq
cHr+vbALuXM9zsd9+9iTRwMhYYiWvCJ6rCEhsi01lcih7vVRfsBDiWSKAos2Eycb
a/ySu/msCnE+2DmI9KHjvnJYAy6cs3rXSgcYgNY72Pi8NjuuJeHHi2EnioeAdF6z
5zrOw/Ol4lPGHXmngP1cOOkF48uOJycRPMPQlzuLFkSUcLe3kaHsEiKoEMdWRfHA
j+A5LrW+YlbkQpTFvfTp9Nb1arYRPttOi71ZghT45bAHkmNCJjlXmtENfHdsbkRZ
bDH9zgszGz/2/qfW/VFvP26mNRWhILnaPz+0VZn5Z+0qPH+piT4YMiVt++nTpnVr
X/qWZl3OtPW8ysMmmL5zyr+fWyYxLsjxGENk+fVa+Vc1bXh6eu/yPZQHq3uVxHYp
4TEGdOpM6FX16mQBJf+SykZiwD14cInNzrTxUFbMnLwYCo6hdUiabppZxfuz2ujA
UNkz5yTpQJRl3HEH2Jaf5oiLDIIyuSUEnZKtcjHziYMrpAjkSbzxqz84M/7IlS4r
Rgj4nWafROzFTPnXD9sFwbWO0PbpZJuGbZz2uiFG5d/UPksz/YpqfLdAs9SCdug1
U0HmMmpRz9BQ2k8ZYE8smrXdlXKiVT0Rp6jKtDhlrHc9U1n8tEkMVdNw+A5UDA00
0GJ4Mjuht7sMCptgDnlErVCjx0vaY6e+FmMwmPnOpVHmvr+sVn4Ddzr+H+iMsMyb
0IcHVX8ZM5xgxQXecLSAqOgUcfOrAhKXdQN/sDBUb4UJYEUcqwaNKkGRZzPZuBtn
52+X5EIb6bRI6yc7Z+WwUVTi7D0rfxlmO6ZNRaOUu9t6q1AS/uG9kxoxjbx41lIZ
I3+SM/WhD2sGzNtmNtBqUlYhIkSKcHH24knyIQ0kWbe/coOjKRYVDYytV/yE8q24
6ggP5O1mwPbEh6QvYdYRydM15tLa4ruKg23PQaZjxKAEPz6ve/4BVCtV1nLFRKOt
v2JQMVMr1FPg+NHezx1zxzoV5hkmq96SYkVLBZpNTupv/xWHBrxZYoiBEIYZPCPO
acYlOrNiQlt416h4CLM1Z/R7N6liVNmDJhw2K3z8z2tXlAapUE2E8h1z9g/CBIWy
lJYV2oNkNEqINKQV4zCRV9ApZpbfbXGx+JC9XDTJG3VCA9TOQrl6wqHUZkukng9v
Q14ATmNp1S3gueHfTBvV1zXM+EvehUNpEDTAwvNSiF0imxUAWX/FQsMGI+5tq0u4
1AUv64qbyiS1XJhpeGdffVniTtzbOe+MIx5Iap0GtkL7yueLWwiONpLPWwCvOWkI
L5qAtcUR5FQhDtAd+WsK87RJGIXMnK1B8z8TVFzjB0PvmHos/d5UpEo13H23/WDo
/Avmgqb9f9ISwYK8+OxnxfRxOfj+w/f0FiXp4Ebs0+Nrf/1ikjbPzX/wklr+J8Bq
JasH9OAPxxlnbUYiTXZUsCKsJypWwDVN4hhoXdZ9VtrrtMExAT60RxuyMAQ+8Cum
+un6bbTORggKhX/k900d0AvsjuBRj+DhdY+4l8DqKo7IyL66YI/MNcwiq5bE8lRi
BvjSeT0e69DT5QkNQx0k6acTGCOmvTSsynTShM4VNixYn8adnoqjjIOg5lpHWRqj
f7eTOHcJAQiEJnXv5JZu1gmWTi+600e47DGHzJCo/1D9umtPtagKnrQiZpW5EWI8
+4LsG+2/WbXGI4VZpRnvmJ9xGMjSEUxRMoZjmw3hqVzhN5yhczJyW2plklZDd2/u
z2nahKK6ju1lwXwABds4dekTazXy9hBripPd6Bqqvry4NikNKzzAMvTyzDeBHTQF
lJOEvjOG9i3h+fWnVBRSeywXVhLsyVBtxADy3GcI0mFMDB039sePxQ/afYR0Pfy1
5lcsWj4lIMTMeWlMgZynH2Ll3vydCHPoEQqvS+UpFwoxEXsfvPBylgu060RfuET9
TL9476vesnkUC6wbT2kpmcthgvKsjCAf57vQ+/nevFnGMn1C/H7tCLLTMHxwnipG
kkNiUvicpaLJgyhNArvafudXkJauiDS4DuRkMgkDvyE7tSzk9JOpR4oMnuRoCOma
lfBac/SuQnb9sbCOf08GSX5WVFoZrS5nR+HtfP1Q6E139OHmTwSbFZp8Rb1WFVls
prZZmxYRMNHQ7GO/L2UBFco5TF0Cd4VrY29nafFU/i2ji+iyYpjaJSA6IGFbNrv/
5X8m1rkRWP4D4YvLTlZ2jtySEBVjOckWv3LqkFX0v0j3FQG8RCbeDzmKdeze8rKO
hnHE3tLZYceYJJXh2fBsYfB0zbk90R+2JRCNr/DHPCXmnu3+Lwa0szP/ySe/EI/Q
ystd1kvMrFWb6zZwqzzdO4vjGvtNzqDRYUCpmTPGDnxQ+i4cGj/IcIb9AELZMfBF
QyFJhoqFJlHQ7eewdQEhIxidb2Y5o5/ZThRXx7RY4+vNsfAbI1UOaB3M4/qZwPRf
xLeY/zdfx+U90hMeLv77atGHhsZnJl051bKK1JgjbjSfO5f/EOjBDl94xFmoprAK
92smNx1JFMA5x/pSUukQ63YjRl6SbQW+Sxda3gdYj9PfmA/3k+ySI1rhFBvUr3oU
D+wTPffCjd2xRR7ACj78Gl8a/dktiy9NA+y4fkB5FdHKRnHreT/E+3n1+32VirTL
UX3Sb2630JJKyi4EcbZPUMbfCd2ONGP/OxA455gQnCQaT0r3vu1S42D7MR89W1R5
vBGqdfB1ukXdYdWRuw6AXQ6OPsxQJefQg6eo9HVkQNFEsaIq6NFyw9lMx7bMQJBP
erdqUeud/CJyXdKy/AvbiQUtDK/RuIjJ9HeJxLdcVS7nXKmwXWCaxb/2MBPIIevW
VygatU2jjiDBjqBNLBcHWPfNMTIEq2PmgSLogUnT5TVIrRdtawETesaZv6hBjKfH
B2xVtX/VEmYg3G1c8T4aHp8JWNwW9K6qOrlA6DriPVxdfYMSAjW1AcnZ3QAijbju
dxy+WHwgM+TNUHcBVcAlM5N07hi0kzKdVi3M8+HKp1ld+wVavMyJCfTBG6Fbe+f+
z4drJHq8EyYYWrQob6dR1lfeccoz6AX+RuxPfSIpeMUtrpUscIc5j3BeuvDbRYNd
2IHDWdPToleRqwcsyU2TBxcUHwD+K5wkDY3SpOCv437hN3EVrKygJ8j+SrxgOcrp
+S/FVpuYEOTDT0h9KwZG5z7k7xG9Kv1xqMwmV6UoefOBOmmZvv7iAT5Uu2+fhcTl
aWsrYboTu0WFAW+tpmJ2C8+2E5iJ5QqambknXFvYPP+voah97/qE9cV2D54Bs1vL
K7VqEY2JqcqD0o0bunuu0CfRB3hhZT4JtBYt29hLISw6t/uOPbI7ylDjx2gsmy+n
R2uHqQ/N8YpN1JG7ibW/TlA1NprsIQyMzZ4S9HQMwwjylYYKrbwPULVrwsb+XzMU
Eg5+JmIVX7Xz9aWyKqCPpRSFL4lkq9EH1lWS3ofQa78F+7rbZrVPTcFDarE4X5PK
1lfba23I9WpSkhGwE5314O32LvxiukkrdxdKReReUnB3sm9+c8hv28szl3tV3NAc
ZtThNp9b+FbrHwTDhA8HABAidj8ttDYtCkGI738bGU5fWUBZVKS80zXy0fVSZNrq
cePvrKLC90zqU7NhXCO3jUV9oXKOjeMPffKeCsOQuphdzFT0CuxDRC+MhSrp+79+
c9MLTrFoXdWZgam7JTsNUNWGVg5vTESQ20yjnRbGp9TMb+twKAhE/LdbZLw0wL1g
Cvp48nl/jmmbNx/BuJ1qeuJrBJEaKfPfmoXTRZujOhWs6ikANvUNE5Eik/GoEgP6
WutqCCe11oSkk4kplRA4ZzDA2b0MW3dcF0wuJgjj8acIhhKz3yHmwnzAZX15m1HN
4WQIBbD/vjjYZnLA2EbeJnQDxjLWHF8LwnuD95uegZF8TCmhQoqcAr74sw+YzUC8
WI1HrMuoc1MPzz5RaW1PYhehG77DFHnEQ4+XNduDl3ehO51SjYXW4OUroDmsR7ty
v6RzICCf0J6VlrmaI8LO1iszkI4f4QhR5qOBgRvICQLYYykipOd5PfLupRYgwutr
7uowpxBlOMJ2lyEqoma0wz+RbHv4Cqfv+G9z6oZyWpZtLoW4HBLS6qlVU+SXBp9Z
8EO+1Mq+cv+MrzaUvgku+8ypZCHgr5BglEMzQtLYOaj61QAlmn+IuaId/H3jVLOt
aSKsqPRBUEiIcUVjLA4gcz4faI7e52X7QV3gger9w6J25pviRMa8bnglUxU3wK5F
+M5R92jfGc5ZBTCOyBy8IxFZGXTazrCM38vh+Grblb0QwhP1vwtn4C51FwJI6ncu
HPyVdaE03zB/A5y6mcWouBy3bol2Y9gtG+2RtmSbuT7JurYrH91mXywb0pBmQPIQ
NqUhTQwI3/mZHAIYoyBl4tPY+EGiEyaBIWoxfGrh+KQYoU7u96DrT5yPZnH3chBH
mkLXpOtqDMVxkC4bNvuzUPi7/Nat+8rqb211RviYvqeW5OaEj3E7iuHKgPE04AFZ
ehM4A3nJPm7R6WUiMVEFPbD/lu0qheR7ujkbA93l4/oLohqUHMiAuKd4NZBAmzRe
l/s/qzpHs0uLL9h+UZPIK6Hg7vwzPaEtbHXTHA3XXC/EVkeL8cg5rNaY/JNNIz7g
qRXfJgnEob9etiydo7ZTt+0/qafE9x0P9DrojlZuzQBOsZqKHglAb1pofRacpmnz
DBHATLObH+UHGZRA0C2fH5jzkENnItSjte7am1FfCHeBzw1NerDRwseSUJUkss7o
Bw6l46Ppn1tTbXBM6ubq28sIzMEOuf7a46+6smVPn7d/5lvtDX3shaewAYJ1Aw2S
z7z1+A+E0ndMi8i+E7g3geOBlypmR8Tn6A/JiO6Yaubp8aQ33+SfytT/7UvJSXnX
ZPPeRFQDu0XxPebUIWyXg6eIpGJ/j4P1cUrdDtUIR20Z+FP51JIGjx2xHqVWMCBY
AHxz9cQRr3HnxVvtU7N4M/kz0xaAeAKOdMB1E3L+/qZX8RwtizdFow33l490kx76
bvodxgtvrgV4OmLicDZ/VO2VqZWdGvKVLPojnUziLf8fNJdRzCG7ZhFo+aqynYNV
l4sznUS3H3vXdLfqLovQChY4e9GMKOeCOGFmns4uEiXUY/WvZxnGQPj3HqzaNcJr
FG5M3hU35WjgoxTEQPP5ik+UKrCZks6NlCUbtFyvPFfHgQoyWddBSNopzw+Anzoi
2pr2Py1aR340eGeikm9qHbiInLm3pXcSlY3mohLnDMuY0mX0o82ZRHfvgbUmOrpe
JfOe1M1XUdvzGK2/qfFViDin6z/FkLgLF5vENysm7ffMaGMTnIduCwEJVz5XfdUi
N9R7DXXygX3KvnUR5mEa+PV/OuLSXValX/MZ1We820tmVAluCF9asmrh4idPU5FZ
OSzS3zmDNr/ikUKUHZAfwWgPSYcIxRiFWhVOKjoUe31igL5BdEgSUlDnTc3oqGJp
HGiP/1jD52fPnacKnrJfUjBu5wirRn+k2LPzUoEUDi2mbUkg0kSbX0KfgfmZy0QU
Xo/9zHfJk5aYxjzuXJ4mn+AtXWOaESkRTFoCudFpoVm3YJNtpN0Qp0IX89GYFtqO
oD8pfLfy54OmVdYHI5hzACTwr2RFvpxADHb2mRSv7nkMLTLJ9GEw7iyTsNlrtyct
AUodYqjkFSCzjFjikmZ9o078ZL5x6zxYIVlE9zb8Ybdhq1iTMeYkhgYXgM06EcgE
FyjdA+HWZB0V011KayGmR1vemHR/ywZFbEwh1RlTm0Bk+rwsKxa0Lu+jKOuH0CbM
gZOaKWkHvchVID0kA/FB551NP5L7UYiYSQwujjiPMuNLVVTYEwIQSV6Z+e1e3EK6
RW1ToOCr3pMFMzbB0FojAqPETkmajgKxjKyS6jHDZYSZrfs4ao6vFbM+nyYT2kHa
g+DxQZ5K3f2WCc5MQNa2atkOO84Fvzp16FQRhvUHQ+Fm8bZ+lhOjq1yngb7aG3rA
a1ESNiS292eqIc1Ml/yxuvdCFOuaR2YmSADt/7oe5p79h/Aur/6YyHBm59VW0jXY
5ke6o9HqU2abnzS1+K6zxTadUWPI5mmqJVVC6DY0FWKH2SAwVBtmyoJ4T297pFH3
6GfPuIywtl0I5Dsj9UFWgDbRZ2+iwItaTgBAPYACXvEZrlJ6a+tVfnwaKwNXYtdZ
Lq/RBp3DOLS3J25ZKlH87WfwfuyMbbsttkZw05HIy/erN7GYkINVdC4c35t5xuhJ
Oxbud0Bq0tEuiVoGkFeS9JQZhTu1yDx2g+0vRJ86Uado7zDWFnLcct5gwt0ch6qy
g+ynE7vVEZhpHmANJ2pSYM1GyiuMj4Obe9FvkxoQ8HWgMWoVQDLyE1vgR6CEBpww
6edtJslHfr4IxeKj7JmejiVs4TCbh5whZzglP3Ir1WyLavoYfI3XnTCwGubnGxxv
LO/BuUEI2Ty0DZ7aINbaUu4m+FfjhekoVheSwog6k9grgM0yCH0D0n8kfD5UlICB
4xELQP2IwGsJFnmGKzwk+7XJKeqmPXdbKidh6zV5v6lRJ0sjd2ZlBnHTUl2Qv3+n
aCOcQqBzrJYWVH94gTKnvQLRy6SwM3SQ19u1aV8iifH3VUx/cCeeFsc32nCciF4d
0zXukwjtmOZO1I1VYaW02hAdQjBvbkzMhUDXd1L3zl5J7JvaDQz5FnjsXjwcQgAk
nyty9t1c9ocrHtkLO9UB28g6nN722KxR+3JwG/uOqrUdirk2ue5wfLntm/pmauIB
jX2g6YxUDV8kvG9xyIyC01zVemAjFJcxbHVFdyXnIm6qXA1uEsF2N3sRevv9iA8z
jP18mEmH2WsG6bh8K/V+brQxR1xugVyfYffOVoPZkZf97NcWJzkS2jbweLMCg0bb
wLYQhVuMWiGA0sT7REvW+f8aphOzSgENMFuQa+K2uX/JWB2T6GG/WnFlbyocsfY5
57F6W37XKmm8noX/TnyuC360q9QZYAHNhGWITtCPT9Y/VrzxjjwqE+QCtkBjxecJ
v4YeyXQ0KHIrWFxLiqkWj/IrK8HOGajcqrbM78syamCE68bkk+CwA99oz7DediTA
9Qio/wPKisYxky94r87C2jWs4TtctDHVGgPeic3vcDjXF4rbhYzdWWF6rEk9SNSu
+v/NjDy62crX7C3Zoz+2ljuGNO8LXeT1aK+x+P4ADyMS8QBhzIBdpoJyHNjD8o2U
GfeczJzHkb1irznfwBGeYES6tr2guLyaRxGpEMvKdsT4JHDw//jbLCKByZIa0UY2
n0d54evH1MrHUI/kaA3bLnVsHVVTCPMxfJMWSiv7i1JafKoJf4wyLLckhTRZ0uLc
SRfz71o2VohYy1KenowBW/IJm0uekzR/XZHYq2H9yseNUfDIChY+0ewiwnsy+HFW
5Y2f531fOyKFCar2lWq7nIY1P5CifKKUtp1aQv9KOIV06O/LH/MQfb7AIlYjFMtD
fg5Qf2jb3juHn6EVyVlwkxd6kj4jtDcbat1E+IxCCKTfUcW2byxKZLm7EXdNanhf
b2PxP8cXJKil3IGOwsfwDHD/00UPam/C7pTAxeWj2nXPTrbeymTjCSdlf44lkaB/
ZG4Zr4MdTdVHKld4YWI03HVd7nl7Dt+B5uI0Ciz6ehcbFL7iaMYMceWOLISgAh1J
SXHjmhDkSgZ9W3hdCAt9ed+xv7FLlkNBP5gN3HQAULt/Cn7RH9VZ83pwZGMhB5Tz
mw5FwwTDHFGsSeqTOMex6U54rFpXXneFVm0Tz7no+ewnZm4KZayHloHQyJQ+KW4T
85pJoOJgk8Q7rrAwVoTfXWbNRnZghS/bxUua3Sr0UV+ba/wUgCY04oAQVukLt/pw
8FjXN2/KN4SOIQieHThCSYEvyRoUJ++MzPGDvnIQUURzJHM/PHC7pqajOKOPQuTM
/OuMg3A6PfwdJeK07eXq9NAiCXVEP3DINeqOAq0e+bBcex/C5T8VAkphfQHzy/Us
wsSlmXMmzgDN6ADWRuP+qoxuM9yEfWKFaxPmhkNu2xLN4T1/tXZE/+z5fpHUFE1l
UIL58ee/fh+n/dQK1GOuSd7oH3JpiuERHMKs45HDT/cinq3YZaw6XrnJ3hRSN9Fm
zteajXGutxDk4sxBD/35zDD3+iV3nImxaelL9PziGJjQ0ejYevQpV+NJUzNRwfW0
XwZQX1oSYhKjsvN/b4OUJb7daEG+HwxgkhQZdWlmAVPX4EPPvJthP7AhiLPHWo4O
yr8cjTZ5qkkUtYSYETxb5krB3L1DnO0kjWGgF0q/jWGptCIQT9sbJ5cYk7MPzFqv
EdE3gjvP9q07o8B0PW3VG146CxchE0J8kn07XZLHVIe7IWt/nf5ZmBykIVWOOKUo
klPud9MIjMSRowPQgfrr4WTFIELj57dxnhz3imhIrdb+/xdATBnFGxQIWd/oiVFi
mcMO8f3nTrTjpHlpv7DYuoZzBpTB0Dw1wrHs7WYZlF3kmAJz+dnfaQJRhEoglbZT
mfpi1102slYjXPJ6mDqFwt/LESIAFACFc3lBBvBJih6JbxUci8yUtVtMoKhuOKhD
hTILju4TPWdoPMiBULarwGcc9YaCxsyC1SIidsHt/QrrZtCNZ9gv7ItdXFyHC2lB
qvHQhS0iUYGbsW8lk3Jr0sYvETfI3F6Aw3SUsKEagQAKDrfdHc49oko8o1IVBhSp
QE/9h5Ixg42ckboYUVIIzs6x5Quc+iJyAEGqZtYFJ0/q83/mo9p0eHb2FM+NQNn2
Qs1DUsdk0bQwoejAugi6VfFmlpQ+L3rnNprNyXL8TfjtjOms2Xzd/JhkD144Xgl3
rpwKiIOadQIFfd0RAy47XjUHdC43gbOG/MgI05nJ9dss/hgZC9CP4SYHyYqKMp7W
CtsxfD9QetrcTLsYOfmHqAukd4gXOovgiyuX7EgwZpVSu1Eug+LHPRfUGYA9cC3J
nbwSJfThxZ9m+SQsimN6CS9NpC/z/4Gw82Px2jAo1++00Dq6iKM7jPRzPMZ87ak8
APQGpU6iAo+A/D2hLVo+l97tBTr1NEE9VZITLh+4Tm0yzB7iCwPfVk1RCbiaLCyj
O1iO+s6TkwDy/+AaDvYN4CDwqvDajW1mjI0nzZD5w5BwfqPneHA+q8E6mQItQf7x
D6eVjSZ+/zl/zgY72518Y5lbD6Lsk8nRHNotDGd4FxUOdp5vW8mL2WSOGKdFcQRP
VWt2B4rVXMjb1YnTetVHWy7rh3m2EyP5g796l74AEpsLLudUt1P+KWtq/R9sEVix
nSPxChpOloXduzjQCXp1WeekZjk9q1RDMyLSQrCWpg9Yx9AY7iVvKxocbo27sDCz
+jt+/XTgWXVJH3y7JmneZq5yu3FWFOQuGcTGwagTbjGVzNE8QnFOmdrVDnVdUyXe
c5A4iAEuO2/Kx6Y7LhdbXuoJY10SLAU6qYT8O1eV27VCILVpxq19wsq3q/VZmBxo
EZLncHmdO26i+i3OPGkIuZn/KsbA8SkTAAJ1zVUT+R4WPnvld7Hjo6zJRy+faup0
6h7fnqtvzCC5rzQA2qabzmc2qvn3Jp8XrYcGY2Y/Gk2unzlYG5MvGbcvnjkE2ruG
QqOsxbAaihzqozVrM/VcT36E1/sZ1BNXzdk2+ZoFBsYljqegESKNt4aTcAZMfLqv
OFYZxrVn5o0Wpmv3Ke7Q8PpeDT+BvwygDZp0EL51xcefM6GNJzvtciGJfVsf5MWs
mmEjcPIh3E3d/chac1LDnv0GRYKh46s+OARy2gt0mddK8KNNMcvC654gsJlM8ECz
VWF49aBf2PbTlHG00w/RS8fQaJWdOzOwEIcKSo7AQPPIE3rNr4uVKgp/wGE1pn7M
WEs5BpIz3Wlec924ZsNKXst+nBGIiT63R1/7EvdSPTwGBdFOnt47QvcnxPl0uu4P
GPpHgyByYCAcLADtfrC7/SrnKDy65hq05jaH6K8hiDovaFLmPyudasxqJn2OTIDb
Oopv1g85Zc+NTabnN7whFSRvdhlRUOFjmvplnND5ZbCybjCDh6OiB28ODPavieIf
XuZxUbPLDZdh8xUwUkaW6lJte7bwLhYQp2JiXA8KwF1M2qrvSP4HZSz6CTvlHDzA
VofZ6ai6dl1cjlm3u3pVQfgFQEiQ4gvX8+LsjN8WZ1oTZlO6zL//WN8Z3SAYNsRN
UcHBkrvyYDPXKRg5KHrsK0WmTRIfs11ArtcM3mOnWREcIzjPi2bx36Fmvfedz+QD
EPJ+5oFqjK922R9RxL5Lhdl/t0U6DbvClsRh9bjbcl6yt+nIZbEyxzFjVqAUOBhf
8nz+FTLcLXLB1Ht2DPYZRxGXmv/60eMD6mJ8/6z3dD56PZDJTgCf9uRw2Wt6TX1v
chVsoOJ4/yEY8cZr79Ypei5sseZetQwii7yb1fhIk4JAKksdhCX992h7RkuASCsx
1r/UO1doqFP+u5vpvsE7lX1/1Ke4HD+0n3ZbZGQiHirTGeLOjhiNmLz8mmA1gsxs
qiyH+aD/SzI00UK71QQwEdLB+nUbihNdOzwp9NMMCgEngqtmB9wggjfxASDHt68+
uyak9dzxj1vIMksrSeW9Suxbv/4OsVnem4K+YFDl6i6K+I92EfF9XJ1yeLJ6UWT2
OqpUjnzPFyxLgtBPYtMtnK9hrIVh0FAYDTQxuOXTWVd7dnAoCO5PT7eY2dYcv9Lc
Pr2n/n2T8P7k8d2lPiHQGshJCxb0Pfd9qCpUcU99yBVeaXuTDq2FiWvaK7EYtoHs
BrFpo4l0MczA3vvUwSBjMQhqmMOcdRJd/HjEzNV49QOIjgarvKJ2vkuWdRi23+I2
eLNkhhUWqUXW/jIvEfGWzkLFn2EfhCU2/9E5kIbcbgCigL+JSjS8X/LsToQLPokX
+4NRuLaAsZKaUF8fZxk7Sm7QXDIcfV1p5Rw2/Dlo+9P4yNAdFHujsn4KyYnSP9J6
wON0rh9YH+pg4VhveKWwE6QMlcdVfpmTjRsrOstsSlydRrrDxTJmbqJmRJ8dc96f
aeig5MTB06KpEwlcwBxBci2QTLzGG3mjYrUrWXz39c2E97YDIYGqpkhvAECCCc2/
DqUhFQBYiUXAd62XJJXt6X6VJ2pZhi7wGvK2Jm7fx/r9gKLc9XBw/nDcyYyemkWM
RnkMgBybc8DsoWtKRnllEm0mKDgtx/531dG3NtRgT3GRWC6v8f6J99Kez/djFr3i
GRI4982kUzbBmaYEOLWohf8mFvQ+X3OkDa3wod24VyjceD+ryaXtvIiFcP02+GnI
qBePiQK2KJJANKxoDprfYKAKAzj6h3xeaAcGUFIKFnJpA6xNNSWra0SQe6OEkN9L
TMYZzHazmVhACnLVED3D8XD/kr9okeGWxw6yhi0PUEk4c8UBGrrpossSXjAC9ov/
9Ob/YVu7mnXXgax5UR0RDoI9rrRegY4YLOExJmHkM4GYrfvuah+vzDv2GS7sZj5z
HTYYYJGhasi5k10C53gCpnX6lReaVhjkp6a0DdN2flyW3bJvCm9rxxdAwe8T179W
hJLDqOygdwhSLccr4usM01KMRikAPaCZ531T9qujIE5TvbFPa9oQPOQQPqdcxj7A
KVwthMlAj/Zluh1m/Gv3PWPyGCNQde+UlautITJA7Vt7jdOyLi8fyZtI2EKH4GNY
VEbodsIn3+1ma/ftvhTydADbmh/qq0GYr238zNHu1kM0Iu+eiq4USjO/VW7sRgvS
CiEc84GvFd5XXrJV7E0LVnSRTeEl5NsbhdwOmFW31bYbxuvkgCN/cbrZsjyalquf
sgB0IEHzATTXI4TyFOcx4Ga6zQCKQCeL3iXJf0HqfQdibseb0/rXwx6IyCudFu/7
G1QIW0o4IZnagWCMu7+bVQWrBk5b9YE2sxNT3DfDAJpEFm8qV90U2PpFYXDx2TLL
pc0rzh58T8A2BI34GXzrecRN2KjoAbfSOU31gHhkvQknwJRX7GxchWnEc9cHH2pI
Nt7nVUgEZkFs1bXj6Qqy+pbNt6Af8Ya/O662eEeakPg5Q+f2NFZbN88ahoK26x6t
D0d4/iFbimDNm0VzV3PuwFCplBhQBa7cgxtdIb5ezuwRhGt3W4ezS455X2Q17yK5
xv+avoZlfVRjo4o9fxIo1lW0DtdpB77fOKf/VN/Xm4muLMOZMLzzQFQI4RZy9UwX
kkh2Zi5PAepl8jG/SCEg2Lj2N0xzr0f17UuaoY5xA+LOz448LhzzjUihsLq3vYry
gdhfkXv8aKXRu/kwQ0cl59b2wEZlZuOm+pQNHe5Lwsu9df0w+kHTUqTNMo+MYnF5
9KYHKks+75vDKps8cZdGjLfU83wrbOMWVgXgvKprHojXyM8nMUrcyVz51GWN5bSb
HyF2PcS34YC5cWqMC8eKuuIUyPkSzudsb52TAkWaH1uBf2rSRoygmB8Xy5I79UeM
Tpb5VcnwV6ZELzLJ36U3Gl5/NKxj+C1mtCucgsYA17mltQAd8OFORhEbvpux6W65
96lIMeGvJN3DTABOBFlKXDtnPuVRcgTbfOm5iSdMx3gkiCYEC5VFs4+3n1hdRAus
3rBvmnm6EaPvHyWNUAt4KUwBLQ5JJq47YYaTh/YHqBBInji9Cw4oomfErcaQMgq+
sMwwY/1z2Oopj9zso2yj/T9pGTD9I1xIj427eqgJ0Ag6iGO6yA9ajyxyq7kRVWxA
kDfmZnB4JQkhXYd4140pYbrnkNporMXhdRmChdYHRo3GXZZ0TICXh4uiYskbw+MZ
JShYc6c40fjGB0ERvglzEeOmuBdP+6cnAj8UswRJ4KyA8yopz//Roflus7gHdiu6
KRFg/nCLpp4thprPuKTUjMPHQPPBKN5tbvgsmYHo1KsoTYtg+HZ4sBnwPOPxjO4L
XDZrLI+d3mUlTfInCl2vyK07TGDdPp4kJiQnRPg4TjHRhf7EAUN5aB6ugfmhN5aH
KnP+Yz7N8vhIUdGWM7ymqMW+WsLWCwxE5ky+pdZdXinV2/MQJFaGqgpBGZD6IwhU
NGhZNAZlYuk/Q/LxHSm0+1uUFhgCGJwR0YOdo5xc+8IAMNUYo2QlKn9TQ8/JN/z/
wHMpU4uKuARTUoGktvEtTCSXOZ3lsElYIvFVw86CRUWH9VCHCBnbJr2Jy3UModb+
6dGE9t4qyZoOGJyZ3kaRQFzNOgF2R9zCxZv9nLHm72t2dMScjMBLUMGgXBnbq1oP
Svo3mjL1sV1DCTSZ2hh22D5ki9v3CUMlHNixrunHYUBbF9VPdmFsxfoVPrBqyqKA
CnbisgWIw2sYwWpowk5vI7yOKTU1oeitIR7T7c2aHKSeARWs1Hhv6zoJPA+WI3Wv
aY6vuMsM1EXS4GJAjO3I9jNvD5CjkkrfZGQuIeqcyGQiEyxNYC/ggShivU/Adn2p
9cOQyJpxkv7CeQgkN3Hl7yCpKxEskVeCP6H7c2/KuSRo3WgaFfgdfjF03Uv2YOyB
ny/F6Qu93g/Xrk4cuRnsElpapnBu6ut//L0JJ4XyejGq72EkXXkFXGuVRK7fIHNA
ZzgW6W3jn3s4JhWkKQUxWeOw31H2wPrBIO32gNhoFT12qCT2aJ9Lg0gfvIUVKnJF
GTDFZJub/kJJpud/PYtcb6/Ovh0thkv7rbhiaYj0e7tsjP9VHkmJJqZ2wLQ2othd
ftKXOlx6ycYLGtgTuS3I/t4quRIYxJaWxrO+Sm8Q9cPJqYUrrIhQFOJubVIYw99X
EXbcL3heV/PIs4o9FXYdzsyDyEEYgKWSmOuWjTlhNA4FpCsJ97SJIcQ+mhFfZ8p2
HPh+Xj8IkCDoduLkImNtx39BlV8AtX0gi0D1KBraA2MPp9KxI/PWd24JcYt7ZsQk
AB52aGzmVL6iuBM0Uh7mxlr5bKiT7szi0pexuuMz53oER7M4HW1mwuwDTcSydtwh
T1leNcwrl9eV41LETkrhH/Kh73m95++pntA8ME2qzgAF0LbcFWfKfxrN1JhvnKUW
KnjXHU2aWHaADNNA59/4LxbDa5icLTxuB43owX2FjuWFKnH6Gt3v7+Z/VPitebYE
U/cpcWpMC4gMQRogD8LqIqlRyGiisLJp5AWyw8R6yxMdXWoQVINDMvWBG1EyiqCF
12Z2JlwBDPX745fXtcP4BZXBSi9oTcL5VseAt55UhJLlHzlcGWfFI4Qs7YkFX0oA
M2uNdTCeu9jddndDDbcdJmPNVKMN7sp/paa7zMuIZofmzJpNAt9kHd0sDkAm2JC9
UVxp9W9faJusrmIjzh3s/5l031/qRvTRHrOG1x0CVZL7yB4BRPGPJjkkAiWdXdWv
0E9CHsTXXISYy0GbFTGn10iGF3ohIOwtdGs7o3xWB+tfutp08nYfqLKlnW8iyKFo
BJig/DudMLrAkuvBdfXHhYM8JlrmIAH90XgKtXd5hphc+luALkZ8xejPJhrBKfwc
Zr46Mk3xqkx8a26BeNI8josEkOF2i/mH9+eQLyDAqSqKyeyHV8ks7AGvbrTPmW1i
w2utpvCN42xI49VZ15iF3VebJtUQb0r/+XygPGea7NqKRraXMPxM/Y/ogvX6gm8I
32C9QYAIPdIMMRYbdh5TUt9h+UWSSHPdcVqosPUcps/jd8zmoetIJ6M4B4xNfSS6
mJJ9Iv4SLD2ML2WQIZapZJuGSFhRJGuWQ1JBpjGYdbQcwzTBkuZiWihdeiMfZDR/
wEPZgz9E+GYaUH168lNfePw+r6rDd/rRoGUtQP7HxyzmB7vjvnws7xEJQkLXBWwQ
ZLzD/isUYkXmH9b4zossDURuRpA+xrinTI3da1a6nFaCCdSHtaj4Ct6n4Q0qD1qT
vdnc2tUq+BVgWOhzXyaxuK0Wq17Doys4xgNi257FWx1ZzDrQ1Ruudgg2tR0ZWdrN
JTfgjJ5TdvgWBaV40/JRn2BmyxgslucyskL+UH01Ltm3dUayt1YMyiKzsLcIyYER
oWPvMQNqedk6tuM5kHeQzNJ6B18T9mgMVGRNozQ8hqpPe10cfGnUkk9oRtIzq/ll
oiKOwdT8iJ12hCKM1/LJe3WzZJTyW/i4gSOWOR/as0jAfbbBg6eosM7iPSGZzrJK
U9Am5fBRdWchgNrlDJL1upjwRBrqD4lDP9elIpVe3IwyRtvojuhSl/WSUZssGKxX
goGKwGzNTqKbq15RhMsu4wRkhpBVAgmjD/85uewVCsLBcPDfYJUzeEszy1Yu10Rf
1F0Zol/E76Hudl+sFg24zQO3UrX46ocKskWuWMN/YK6BmLFEnNkBgc1AyFebnLvL
Xc26Ex/AjUB1UIuVf39nqioqOL6KmZKX7+4bAZaSUzNi2q/rc7+QMDNcH1pTISO4
VcNWOeUCfTS/lTb+62Pgb70ZMCtJVQT7XUvb3ka36SnhNnnDbbv8MJxIvmHsRSx1
EyJDJ8gSOZR0Nnj66NeEMllFcpCADoHmYk5p986Jq2oENVUyuQ5DnSgsO7jWsTxy
Cw27lMEY2cWHJsY48cG25zMnj+kgrAEItBPen6uOoQBQxM60zm+/UzXQYe1UG6bB
BoseibQylgPnMqroomko28a7qDdvVR3Q39EqtCZTyon5GPYwsaQiFjf0QqccJbqL
JxeiefS5pNjB5WaKBGRQioV48eD0EqZWluqThHj6RT79sx3vUR5c0wV3JfCnJN6T
6Wuh9f/TxK+PpkPNLoxjSPDiWJCCCYkOEkPQrMa52GgSXh2TLgDCMFBMuik3pQEc
+vz6+9ZCpcIplnJANsbet6BjuT9T7EkXRrRxORBCbUptDG1VOHJcw32adyGVWV6V
pGoDG3VcxWCq+o5o09ChzJ2wp2nK7BROzrzhMwcObpEFLes8R8qHpBlo+vMm+ZgU
794MlBd4pktl1P97CvwSjMtAIfk0ar2WLutqxVbTo/FJSPJdxs74T4Nwo9bro8e6
C5++MvUbKTlbJ7g6WRHTkzN1Xix7Z+TjutzNmIAK0IFddePqLms1Vabk893aVdUa
cQVwZTQ+vjfmbIjokjQMEkwW5AShEahRZX7I0X7ZQAGo5vOKcrmHCEMoVJFPawR8
qG36MAcganiBZV6QEp6SaEP6mew3+CppPzAxzb9x/ROZZntiDRAuarU7kM4Vq75K
nUEdjINWGRlvxoqfM6S1/Is24kcPHUiUcyWSMaGk9+4ZqDZRMdEdUN75w8+vw1Wg
T4LdnvA0S8sevShcARgRBicLVBawfgm+9Ebh9noGoIGppEzDeWawRqnsSVkbUAPv
lA2RTCsAFPdcscfg+ry2AL3o5mZgsAklV9ZFKKnVdbzl68APGGob62lqWaZQl+Xz
2GomOHCSLCTfoLZUvl+1X/2j5jpOTt7FEJxsDLLBxF4bBaEZ+aaZUAsdvZz8g+lF
VIX3u1nKozKVjBN42YYTERe+r+dM9GOeuTWcGJU1bzWmOSGW+2b7RU2EBFoXqIv1
cSGu3m/nKL4cEErFBrew1U3MA2kMRMm8uwcrVxROxP2EzyvLh8LWUaTCRZny3M84
X7o9lrqHaj8KK5QeBApcyyoYyaxNyuAtMIvOdk8rqkk8t0oJZj8/3Ayw9xLABR9B
Fd6EZf5jpL5sDY5csPC5mpxU7szoku6MUhny5q7hPSg/WqyHv+Yuy9/mMYzPYXAH
NCJhupK/chlexFw2KXp33HYQfmqwiAhKpB6f21sWdZi5773ruggfjwU3solqJtA1
6UikoICZqgVuGokJFWVTcg+7qprcjGM7JAuMgocyrtSjISWPSzjisSHVHGvlRWiI
/5bfALvUo/slq0WqvjE7He/iRpjoKZssQVYQ916h/TExqWJkM3HfcKCEQH5pTJM6
D1P8oCjXfqLt+jL3Vo17ds2eDqVHyFWWFg9sug/TvPWaWVoITNGgtsLQ+9jOevLx
mSu2uIJxh1xVetW/KLi7DMCRba/+rOWLJhYDvEoNcbGPAJ0hKYXrVFnhqNFT24Sx
EkMPG49EQoADbSfGP3iJeyYP0U7uJ/Gl9HTZCDSmCGWJbbAjXgg6KJOdVWhn2bLm
ktGjPA+7ziqKq7HcteqH85M/6fdbwlbeFGdMXJaCfdn2CLCuuiEKsmqLKOYn2G4P
SjAqYBgy/EW0unVyn71m5RC6j0gvhxHfrI/9Hopz1Dh7ctoXrVu+A7WvEbhn3ME5
x4/gZUxkqKS0uXPphZzScTKeMewNUxmCglir8KZbNWeqdmytFRSZ3O6YuOQWsfJ3
EyaRQ51RHnkzZSfvKY1T7ekM2MkP9IbxJPay6Xul1BmSVG6x2voad3WYBeFglQQ9
qJnY9Xh8PjySGfEeUux8QfIgfwkI1iLRDeDbg2483+KgO7RqF4muVYXtxSP4LoL9
yMGEGurjgLlCuJbM5gjka9NCCUFh1hYYuu6uQ54oGDSfgNwAcXUSDU+/NMOvSC2g
Q0RkBf1sKDrv0JViPrOmuOQMWDCLRmC+UaS5rgXC161Sh1VfTkBk6PGXLtYj2u5F
ZgQoNxTG11GX7CQwYHUHLxXUZYR9MCNnxnpZPN2x16GahHX7/xspt2BGkUjT1OK0
VpY+GMSBPgjeOu8fGWwPxH6VaB1Aqign8kXqcwbkpW76YjnoxcjiR9NhHmwH3TX8
p1fhmUrKJpoktu/AcIlM49zdlqyG63Zx/GiA69IsO+KUexTHddy1e5/5jowftwum
rYId93rkops731U85nD3tIwvrXzLBAvZByH752jISh4AfeRP8OZnRBfKP5YDnz1k
IARf/EgHN5FkW80kuRzL1DZYwU8X/WFLDu8fCRLs6afbrfX8GYNOaNRSRdEgpGIo
ZcfZisQTECo+b82IJs69O6VIehya3yu6EwdoLodrahJuie8soK9fDVK+U1POeuge
vu4RG+T0MKA3YX+/fPPARNAUMuaH6p5xO/jUWvp7TMqUdJPHTMPLJEBJxnOLnMP/
u1aJDDmiorzyEUsHDoU363oCtv2uiKRrDjaQQucZaR9jtVaa44vRTzwG3VIVjS7W
NZVEaMQBV2aPDWXrVg03H5d6f/ObaofmQq2aDXd6yqHVEZ3fu3Hv9f3d8lxn0JMd
pHOBrGJfhXeNLGRPhsOY0mXV0KcSMmLZR+285I3KLX7OtMD0GKYE2x4EDrKsHvhg
80lyA8rLxL4+rdEGTFOSxVvIVacr5qRGZFhMugL6sSbCXBT/XUvARCXlUcrjr3uO
5wVLknjPxzjTUrtMsd7BuNNLwO9HK4tY7AgcMi4hEmuRDfJiCyG8bPAcCe60lfMz
KJ5XbYY9dv1kpAHHXEc2eSRj/6qDI3FzVluGCD7HiHG6AskDWNWqDnKfx80wHwZ6
ULr8PDCVWdSTNMlzevx8VtK3lwM/p64oSDlj8HRH28mzGwceXxMMHzIpqon9B8Lq
ktDMTaHhmnwpev4IOtAD4SZCnDUCbLjkv6s3AcepG3XRD6IAVAts4ij7sPsVaqaw
+/l0Ua5dHlXUYjRYuGYDeyRk3z0sWy1SxaVtVQnysUYUavyShU1F41eqq7lh2coL
CmwNqC5OTG92UOQTLJ17R4PAFe9vtr6r8A2xNSyyP3wT7whzppibCz2bEyxR/Keo
EtWFwkT1g/T0rX53jtmHpVXVRMZ+1nMMH/bDaTok/o8JGj0GvZaJT93P+DCZ6vec
aOjeX0rR2JmgV/XoDc3cGLFo4yq//kuLvM5nYgoUIItvqgvj8ZVCDXG+GK6XKToL
T6kDW5DBijs+0Z+84qohcWBv+znViUHZgG/oHDgEo7GFa4yDTFnF6HapYnwQ1uLP
n/vMcvwuQBrnkLh2uCBD79vJgnhivuiLFlqysYMM5eCy62zbX4lb8En/fgx7wU3W
3v4NoqCiDitvXSF7ywe0kcqWWML9jLDNxgOHM43fStAbqZK6AmC09MMrTZ2jfO/n
DzC2zvtDPr4/UXhsV9uEWfxoBiZtgrJXpcEiZ8UvfdV8Ui/Vf9hKoYmkqovGt84u
ERGvvnX3vBGiSZ7hM4hNjEMWtRX8oauvClxWnLpNgQ2Rt5OlG/ZvwTxWfY3K0ukk
oAzv4jMdkvrU9iTzDHCKm/iQ/LPqkV6DdrVbNed7Bma5DqU1fVlcHdt0D/HlOp8G
d3EYjWw/KtTNoZYhY0mwgrKZjwKCUvWo1+4GdtiTN/xYGMqWtsyRmgmvkGhZEObw
epv+qNc8zsQb6Z1XNI8sUEbepwNG0VklR8ntpKFjqf9VvjTPy595cxFUWjqNhcAG
YkDHZc/81oo3eCiB+Q8PKRV2CjGV865sv3M9O5dAd0J/ww7YoRnNt2lgkUz8TH6G
CfuXNWpblsKbM5bKJz6rxVJhck8bCsS87qHtOHP4/uxnDp6LZCdWqamv/+bcqcQN
k9zo25kE5xyaBzae3zKYCBKsTn5KKm9hyBktZ3PZISvhbpVDP+OEN+jcpZPVoNLc
q0WZCsMKLEtQtl5znPEhL1QwI80YB5clfWmsgH88cLzMAt/WZbBhu6LDefF26cZp
+AMAYwPU3ltonGFJyZZJUlCbdJSZKTJ8JG4F0Zw2DgxR48ADrA4Ns92lS7XsHwao
NSd2HvjsWC9ys3JbJUINA8Jgpl4fTOivokagYBRa5DCb7egn/w1HPpWkabTc06iN
6M1mjfXdMu/MJ+ErCulLpigtjLMTCiDTt+v1+8QFVO/vl/59m/H36PgvabqkhX9g
ydSZpIGHzzzew8Ura5KEJKRFlHFs3gL9CV2nksVki/+xbIHywvSGxVz8CmQlZ6ac
jVvZipfeQUqmgpoSDtZM5Wk1zqhTDwZMHvsfAffC+XH2b8RJ+eSWhiue69/K0+eM
aOATaSe5/B7PjdNgQJYrihrCc4UVhmpKWImZYziq9E4r4sQFPbFYubU9ljuQDoj8
NO2nJ3ewbdaMy63741knBMyvKz+S6kltfZmKXsbK+vD+s4a00aafB6ps5DHhZG4Z
DrMOFIlVKzkq3h4ahii1XoorhLDYa6W6wQD37WiXwOerckzz0HUa09cFz2Me9EuR
H0+ijBVhlXAg5tkLW86R2xutI27mls3YB5XnX6eJecGjSMIton/Wajw63SA2kwTx
ZbIxDH7HriR1kAwaqbKtWwYQU618EEyi4uf+f7QT7YOnwfYMI2d38YjKhvxAW5Qm
a9SoGWFx/hgGPUB7e/ASX8AqeshAQGCubUlve2AStkd1QRouUelJAPOznkouqRsX
Kuxbc0FndnglXfjZON8qxgiTKn0JG6S5NwqKSMsuoSzt/RAeO88OWdfWjg57WaaH
upXH3sXskF9RgLCKxCQKb++XZ1p3dKmIUTnxQhWHBH7CC01zC4VB5XK5LvnQX5Vv
/xNCE3TrG+JZos2EwD7TVBRvZzrjy1WsTTM29IEJfBxxjYWRgw7R5D+u134vhoZ4
3cp3mlOP1zTgQ+OMlqUj7qOD44YanSfMkIgoX8GZvPJr457fIISE8iSdxy2WVBk9
RivR9rPeUVid2oVTrbtn2wI0aSCHBKhuNOiWiD2euILYpe5brMx8Gwlqmhj/epcX
khs+sXFXYBgoxeHCP0fEjCCU94SySokL7S/9nN09jSi4Cgpxu6OhHLtlVjyMReF9
bnWP+M2/oUSFpTNttRq6F4fxqp/tLkK/A8lmf6na6UmOYnhDr9UCZqH5JcvqwzCC
k9Ml5j2i9I3PEJbiJjCki0wi1vQN7htoJiUcPuN9esyYaM9nkqPzaZh4X5uFDggN
AMX2X6boNmWrQJBV74HGv6CU9MuTNzY3pJQglPGTLXF3DRGQqCLD6p/WrbLifvCo
S0UUVn4GOtXaDfL3YxnKI9vrPZ74TEsXqfsbudhpMVsX6F4ipa+Z4E+Mh70gAtF/
J8q2cwaEjntqSf1AUEY8Ita5ofVu/E1Cq1fj/I1dt9Zbs2HJ+qABklxcIo23koqo
JUhymTlJLnoludaF8tbr4gK12dgWCTlPkXnsJ1vvaddRapIJ8y2ftAuNWhSsOX/h
pCpxYJLBZCmIFwMBIyHxm8hCo6L+ykeUASnBlDIedLc/1CS6Nsog/7KnZw8tu8vl
QFTtAKc73zMlXDvQgZlAI4YLMtnmDmqsx6hxbSrEQSIIynb8z6c33IaTSeE63qzV
9hU0nV2aWYqYjvM/taaaFo9SUS8E/wsn6C2L8jtTwHspmCtqgSkc7T4KYfNlMDoh
MeWshcHClNrKlVFQbNaaabrT88l+4iYlQ+ULZ/ty4k0/FA1A7+Pw1qq7irZYLV8X
mdlkh3UXHcU2Mwkv5txkoPIUR6R+HDou2HQJMuF3vhfF/5tHxqbYvPmde24QGIt6
i4THvfjy9CDsaDn4/7TxkTCmX6g/+d394fKkkevyf8YbF0qnGxcJnahlwdpxEdys
9J/ktSkK1YaAR+GenvKQh4dgYt8TfGssupf87G3Ogh3tN88Bmq9oTerfAg2kX8rU
UlhElVCePvw8pNCn4g2hBGS6RZWnMV2vxfXbonVWTaYMwFG9WJ03cnXXRPGhDTe6
6O1ikogWoSmWojS/FdzviF8Uq857UguX03qIcIja9mCIgMGA3ArZ0aJebHusd/Au
3xqDI2a0e3Wj4mctTCvNqmyO7lMgjcwrXio/p/D+mClArbxbUb6A0OGDTOuU1fMT
HzeRpcTEJKm1C50LF3Apo0VA/uW0FFKjTRNaWLKIXfnY2SxqYrd/AKgm2Ewjtude
WuJST6XONyjisgp+55cHZ+jT+bv556ztQsG+v5Jkb5yJkP/Bh5zuZWfm9/4mZFdp
2H1lLnOjso/da4g4cbLiVT0UPvOBcDTGpDRAwKq2Iz5vCBvhg/1TLutbOgrrZ6Qx
X8Z+23A+hr7ZtvXZD8jjMy2r1Dub2bVWyuIspwWQOG9LH2tqLlml78EeBzGYq1f5
Rq0+8SoTnMI8a12Tz6EP0YUZYNsDPIyK6oIRUHMl9Nex8ILPKlnY0k5JPClLA6YR
oKlvggdc3VITa/wMma/xqWx+C9q48DEUA2eFeH4ECrGwLvwahrntWGDXzMexS8hv
aTWpMkc2mnuVd8OHPm23Sv6ugG+1FEh0OhoGyPVsNTcRjxqeJHKQoag7A7C7MWkX
oq92s7C4K9gxmG3N354xyj5pAr/Xc/eMLgY4EFM24o4U/jbjWDB2xYNgRQy23lmV
1YJ8Ygd6Py3iTnl5PmVOyV0Y9DHG5LgzUZ6rA6KijOIvKHAYAAOW85/ZySfwNz7t
W8o/5szDyBwks+9cSecXLGYLa2/jcBG81yWk2yB2Ss/I/QInuKpGYqOUJrT2HXqK
qQcev9++6i+Z+Xd2/dJ7X99GfuVscml+/vlENMt+wrasUIRWBbroLt6dRO8fqXkX
wgxUUhwjDMxyg2YhDZeEot0qevCQnVOQVNLy1Tj6P6AosuAvTRlGFIJXDRmfLQPF
nIkXjpKQ5md5cLemSkgwgjNMPozinLbpyOS736P9NpZKesXEdGVuS7mo1rWpuKZq
U8EU8k0nDOnkYFlTMMub7sR011/SHqXE+iSsLeUUtzcvfvjHq//edY/idtTdCMRv
mXyRdIVCua4Geh51aQQN+J1EJPg/up3G/86J9V3RnqbFen347nd+lA6loOJsLLsx
XtzD1GBrrclm763j0qeS0mU+XveSg6mZhFiWsaSVyTp6GaT/ojUaWC4oD1OBSl31
dXQMM4sPo49ANUgdr3pWwLes/OTVuGr3Fh+NZpXz7v56Wcc5C5wPWYW4bPRiXX0m
f8TBk4d7v/UHxfXUsiVKCEo4pxH3gQtD8laxvj+MXxWErSGrd9ov4WqnlLAxR0aW
0t4ZfP7aqU412CXKA/fMCxc6i4if/wDpNVFyndF//Wy73veZiYu1yH+wso3KSGDY
4MGprS8jS6UElr6JS23fAHENY+EnOWKAqzRYf+OUyCEnsj/MBy1w7YntDwVWneT/
q+8nHo3yYL+9RnEMWyr2jNpc2PGTf/xsZjYvVAhwN0lqbLMSE6NHR5p3HDfOZyO0
yHUNwfJgyc14hhF3Lnda4MepDDDMqMcZ0TokbsfjpkEdzPtkiElLFvooW4ZwCUqQ
xiGdmbbjieqqi6hAgmEfV3e8vEx187GGNAM3pvEABo/vj6eThhBYLzg9UGZ0g75K
ICnUE7Px2xrp5IVNT3bQ1OPx9SZRkEwEOluZCT7ki3LcknH90k3umMM3B/6cdUwY
8xjrU9Xna1EJ6hEhZ9s7fr+fr2JDAReVDA6xdiLHT90K4Y72Zsg3A9ekXE+4xn/f
RRAGUj7hUchhg/rNE3UkqDWra3RYMYI4xLkeFJqyc/fYjBYZtkcy+QpOCPG75kAR
gnH8wOcSNX9NoBmS/CBXK0e5AGPFA30KLoJQEXTzLlFmdn1wJ4KMZfivnOp8Sz8J
KRzMuy1/zpwf2qh82xmmxLMZ3NnIF8CDw9mDr+93UkX0OqMiAHkTl0dY+PlrpL/M
gBWy9JL1ZBosp7/ELmtAk8pMl4uXca20I+2R6feFw/DtGYu49lgrfHx0LK5rL7/7
KtJNWTihHdYKVB6G72lId2xyg3o6j50vBXJrvoBb36TY9bPi7Fa2b8V3I3Ax8ryF
7uT1iOumBgAp1whymIBPtJWM6GrBalaJKsApsP/im1PtUlPeYKlUvo+0r7O9feMX
RqA4BG+Juwg3PtsiIZQiPfU0YPgoevIbp/KIhJDN8kuV7Q9YM42xbv5eqCIZhgDz
drVe99gNfvyIvYVMNhUNJ4D+xXNwCKQAYMzV0Mr4czU4/Cxuz1osiDV3NWjcnoH3
8nyvJ5s86wGJQz8D13UJQF8f0QMb25TodlG3+kXxkozQae69lm9LW5WdHYx4/+jn
r5I+df5hGVH7GDyjDOfuEb1qCu08pEmWMD/nU6XX+usN35VjGB01YfeggGoZHsD6
8NHbE8DOJCWc9ecJis5uai58uIMlgtgky8yMljK8vfQilhZFs9C8utoTQKTR6HGh
ckvhYywmS+RkfUJl2HGVPVIta87WauisaZB2z1zX+iiCGMzKzDL9U480na7kh8ON
Jk72kH54JS6xWWRrkY82TOsTVKcH2QlmrSHFphqjhbRWtokBqKa7EAxDxdRShn7C
UX8gIZZ9l5FRtmQIlcqdFnck7bM8CGO/T2GGJOLKyqyGz6rVCl9666WADPKT5dgA
IycpvcK4nNpMlnJoQRFYR+Mk8JD8q5ziXTe4Ditt8ZQWcVYJYSLMWohXEW5Q/LK2
XM6FDoWMRbReVMovQENh2w8HPATueLN1zzwkn7GEyPblNXh7WUipAD3r8z4Xqdss
QdNNVza0Sc/ftVIo4sNb+Q0HqJVlf6Xnyf99kJAwyW6CydaLptrGpByuNwlpRzMA
taprDcGPx2h4XIvS1rBNhlcL0Y0mqgDs2qrlP66NreN9qyUJwT3ZafUVMYLlzC5E
axwpTk3F2uI6rIoS9DdAZ2Hn0bPonM6On2FfZoxIk4SBrFK3DEicqbYb1g1xZSSw
70Y113ArslrcK3gjlZNVAd4S6zFtUFio3n/nQ6k08S3Xr8S5lF0RF+Yw24luOK+h
1S7oA2nSrWHBxKVHv7dnqSdvDLM0qnEpSDXdZUh6z8OsHqVtLZZHhZCrEyXhZ0nU
oAvXAPigLewWTqHZMYciY5IuKW67fT3yR9JPzsAdGt+eg6wOMf7raXaclIjV5lFQ
fIdRFBofIqiMf2JHrIOBo6vOyoFjeUQ9WvmNb+6+BhqAFhwxoR87e/eP2jb0tDe2
O8wCMAd+RvnM0vsPFh/MDdNcMUPLA9XSnzz3r16TJ28lKMNgJsJm640LpXBpXBpV
i9JQbzbAdbSKrifLjOv19i/SijWbceeCceT+NqQt6bb8VBaJk0GC/+c+4sUBKhnB
GkTjJtQ/O2xGdrurCNnXWYwniVgl8UzlFW1l85kHpnZnK7e6q5vWnhI9Q/n51+eX
oZj3SrdhsO1wc6YnmJpJZ4rc4yqHDjny5G9aTesBxuuohN5QOphHHE0ku9ILeFbp
se6yQ7oTYeO2Um0MEIPwob1sMzIRliPfJr+JIn/MwdwgywB+nTbpMYxe7CeozBUT
LT2Lcz7KxGoojXVUeZJR6wdkeuEM3bMTRsHyhNd/qE/m9TKDojCL38DIJ77tsWpD
IuEpKzQTysQYP2cXzgzAF5Wq0WGtJt+coSwq08RVtM5ztIBqdVaNNXpaVD6Arii5
kdLi5S4l1b8ZjdUYWBMdNvG656fMnvnGr3dbQqaCkHIHy3ZMbYsNPEZDpe3unHQC
DwqHQF3kMIZg/HXiTO0VluNmGKfsi6Soh1vG7F3sk47ZCiyq56O7V0jvlOaKSJFu
WoIpFfm9oFl/DFpH84HtVGgMh6kj545/0AjlF0lQ2fpLcd6M2yxOhRjA4W9kCGJb
W6qpiXvl+1MNZ/iESU24ChEKjoq6qZOjFUjnTMwt9Vhlc/00eh1VayXziWzP+0Hs
8gQxq2vaQqY3NsQ012mB/WEh7oG31Z9tTE3ehYf/eIerHcGvLghJuXDxcJ6w03X/
ONba8BOKX6/XQUlmPOlaB64ZhD5jlVe23+tTGrVs97++gFhohdbde+2xMfFKwOE8
NME74rWwCUHBCSpa1P2nGLV5/u+EgOlqKifjNBWii8kDY8yPbStvNAl18XoDagZD
u/pVx5Oiyo0QxfqcuHDB7OEI1pJVf6cgxBOil/U2uTP3S1EUMD42fxwQKZPdHlkx
BUqoZedcz0VedbicYtrbUe7lSuw7AaZN5QNX1W2DoenlwYJDi5fwZgaEbin1kovJ
E9tgBBRyF6tdXsvMjMzJhI/d3kQTPQvnKFquTuEVF0TXwSh+7LmNrYtRkCDdDAbB
r8o0/UpuJlQRSnuGXFy88INx12eoHwX2dXYLB6Xrzjh9heNJnkrEKu+UGdFcJNXt
2jIkWxqBzgDde7li7yr7dq+6AqVnntxeSzgIOjAeJUgabSzDCvQy3CHkkJ8zBkpD
Ch44k9A/URKNs3aW9c+BN4BVNoAxHERX9fsVYFt7oPI36FJ4s9JB5GQaowLtEoU3
u+r8IOnRguV5C/PjvEV6BuAUzk5zBQ+urnvjDJZvzgM+KNlSKR3mnVasLpn35fPd
QEtMopdC+tYqBWuCzz0EeRniI8lfOr41pPKJaA9IbHAVU7XRbpLXrpNYqzIIyVSK
0JHX8RYW+3VAeZPZXG9xC0ObgoEd8VDusYe27Vhh/SnVAxrOVtb562Xil+QYBVO6
o/xPbYvb8y+xrLuDcsZeGByAb+quajPDJ1eXZZ+cvFp2J2ZsGtmHpZyG3ZZL847y
sPuCQRCa8bMQ6oLfXwxZqgOm6x12wu/hCYNS3a9xtsvzYdOn/zWMzkPZKFm5BNXh
3Q4d95Yk3TSxGfohEHAFkaiRbe08DjFWMTrsZWKRmUfkqqkjKpdGf7bNaJgxOjSD
20YhqcFCOW9jmBkXxzqZ3VBDYHoawa2sfLWwji/bV86XMRx/j+bz+L1FyoGVp0yE
QHsaD4v2voGJ94z48MSD1gj/UWcUB9KFMo5HN27Eo3VSVi2fwXjKYgEqNwHC99Lr
OMeyFCEKHkIX2SnZCXI7sYC+GPkNZ3dURbguraYg5YNMVl5MJY0jL7bWr1ewKgUq
EIKQy/bJcZl1sgOB8DkS3ym6Eok7Ete5BH2mMB1dIVeInGEWJrm/AZ9CMmkNPFyo
Hm8wKumUIbqjcr9GXFKYeQcds86VPGBaxjkc+ZycGpbrqWN4yNW7SWl6kMImxqK5
2zaVadzAtaJAJwk05eDwvfAEhMGmMIFPERDyc/Fn1BmYQjWvKtnyPUr5RmUyGFeg
5ADFeAy3f0eCgMqYq4sRw/s/A/wOteewpsyrQFSBMhVk+nVR1/T+ShxFmXoLhGs8
B5mRIJMczsY59yZqDzvAn3yPkYS+2y0I09Cws5YcP4iIRnhemmswjFNlu6DKIzul
B+qwAlABry6Twj5r/KeCIxItyuVDfP2G7jvGpYLuqXVY/K1BFex6YFksrT7ZBbuz
txVQcCtO5MUwZr6bRIZDHiqifieFbIjjiPUIiaCCtGpsdCm440rIljoEJhpCuTso
uB/MaZ55I351AoAz3NUytVXNxjL/SCsTyE0I/Tseyc4cTgWVYeg0GISZQKmR1heh
JMykl2eDGHkYAK16iu5s4U6F8zdQYxjxyI5t3qTtYzK89Zs1XSt2k1YtV9xhfRWr
GhVCYjR2nri/+AwhjHCutvOtVoOl1xM/1piXwr+93ZqicQsPl2VuF3Ud4E8POO/B
OOsME7jnjKaF95zMN67BKm8dRrD51skc+Onv03cFzv/4B0e/mLOrZ/8w+QoifT3v
1lYBSk+ULJfdKwINUsfjT9/60t74Y6zrcRw/Cb8PlB+kfurMhW0lqIU1MWfGifQ1
+vlPC9eVnBizOSKhBKJPW2lNrDBbnoVZGrHqeaNcYz9ODbeTtXDYQlqy4R8evnlu
sboFfksku1/glM5cXGpuejn+kojHRQcAI/sV1NUkdT7PSjRpRHfThY0+AR1ImNTd
Gx6flCrkI0gaRIopJ6RhNOdz6gPMNmIHIgL0QM0OPSjytOZZIsY6ofa7CTHX29nQ
kud4tZySoL0OqBP/2KkW3PoV3nKUjlAxWrbnLl1TVyseYvuq/uZyA0KRjpDg39bT
NtGtM2IkfPO/a6/UxVR9wlmDwG+hjkqtdEkcpBoJtxy4Mfa7k37uPWXF++e6EseY
ijOj8k8MErB9lCbDjqxJoNEQUXK08ceOI4e1r+Hk54sIGTSQj8i6LWSc0ElMBsVS
MO+0tdqJvQbKt44zwXp5BKVbrTngegnJroBJk59JzdCI9/DV7eY4zGjpwrKHAXli
1FRJtebtYVPkvSdQ9IQTzh1d+h8O/7uRwpjbsHaGXdxchp5U+WXoWBUFDao1I+Ax
TAXpS06WkRrPDoLMZUcWi+qmiyqAXtNzv0giqo6DHXDlD9AI5e+ZznPYnZ4TYjzS
6RiGJuHIwVgcvmgUowKs3xEcEbDjtp04VCQ1hwIajjy9VSZ9Y7B5W7itB8f82lmJ
hRCKWztNyFSN+X/z4lugcHCJlDWLRP8HSYT6awOsxqNxLVibdjGLsZgFSnRcg94B
shjmq3bCWnFt1IqvBP0Yx19lA3a6A74RZ6x557JcQ6J0vuXBCXCNely4JzRzg8hE
h4h1zvND2LZZ6UNnv1QgrcCEp7Hmfr8yL9QDnFt+r+3uOXAuydtHdWKYJeA/3NFu
hxyOCxilROHjomCUKDI453oqHSEfje3kwN/J6OgNqpXDPvRdydwt9L4c7kpwYHWW
Zde06wphhbDNU+o2QGwy+ScGmggsvd1bGsijEkxUVjAv/eDMvYRwMKMT68IkRPhA
QjYvy9lzfyi/j5XEogmuM9wKcmW/c8yNiPwLJMs0syRvF5r8PpWw01y/CSDjbeAQ
LhgykyN+b2QTnckncxBkw1gFXPmBWd14j39l7h3sgkth8BNzxFtn6E8FT4CbKh4E
N8sUCKSKPRpN8n4xAue6XOKvRohOjHzq89OjP+eEsMw0NgpCi58aKv1YBWqvfSH0
c/2ZYnPPimX0swPU4ZeY2mOwn66dNYJqnBmxvHZ6sLCGwaQuDqaNozVrMv7/3Yvj
dlVRUMgcUJgxiS43RDLzlDZnlj1wXFu7KR3AIo3SEiNbv9m2SjnfaVaNP4TXEBEr
+HHTbsB/Yh/3YPnQbr09r1IcMLhe0YnUyKJCPDBdge/9nKt5S8tOxagEDkw/znol
Uh32RBEcn2Ofa/IoAacaCR8d12UAmaqSfzvzaMPp/16cPLWJ2AjV82h3LYrYuZ4X
h/xwn9u7BF98PjFaFtSMAcr+n55QzOWD93jDvr4uMVw9a5tBHSpxuywcgXXCqqIH
wMnKBzi1rTGCX19QUToGmcyPFXgW1A9jwdfamF9uAFmzwC9lk+1/Z++jc5jToPee
FGvbsTbKrtxm0O7lVPM0E6oXmkS/s+WCnLbeWayJPeNjppZ6QRY9YGKV3Rnlp+et
xC+2R/PCkLFmrS2PBTmMmNtXq7yWeo3LbOCDZVlzDm/qeQ9JYMSbR7j0YrjXdk8U
JKSiiwCGWYjD9MBur5arMnpwNICC8E4NjFKdSKl5R51Zxxozq/MNBiaoDDt8YDpN
OjCXzt9XgQXZ9dVG3phMgkz1fD+NQpPaJg9LZcEosq2E6zPW31fOf7cHa1V4vuGn
3bGvPOduF87nu9jukTGrirGdSuzMAlBm3u/ijsUUXAA/XJecUxB7p7SpB/nVeEZv
ySr33sJX/fK1IAAXp0gtl28d+m1MctZsmErgQMx0g7417MGsETIKFStcgS7Hxs5L
jM8oWbIoscWIpsfOjX1anD7jpmpHhlGRW0kn7/sNkp9dA6kdKWYIIT4P9vPoEMej
a7CzJ0BQzXxQ+8vnrxmrsEMl+alOilqcUZKSdc64PvGet9Y7zEcdxEHWiWNV4b8F
ybsUXKvkY55M+l5z1wsSUdSkkovqm7diJxCgM51Bd20XaGVHDbLwgFuhnVwsri04
N7BPHUx+kapySTyPnJBy2Ez3nce4y9wgT4H6AGARRVdPoXp30clDofuBaj8bfpvD
6jZ+zVH0KbE9GO8vJP6ZWQYxlPAGj3relSBzdWSmcrG//7mleQv4ryfuR38qFr5e
+5c8xZ2knorBpVHfu+N/6wzmLRJReuKZe55pDd9iZEnOPYgAHn0FvHHtJExeJx09
Q6yprUySQE96TYpP1Lw3iJGdgkyM6e5yaeYyEv5PzdW5t1K+KpTTwayxqzVYhjDP
HpvrCmeZoYMed5p268S+xVukXxR6ARPX5v4/egfJh+ETdJ5Zy3FPkFdyPJj5qCNH
wLErt4/AhenbVqb0YFLPFcnGqc2GR4zbOGMjUi2cQRDluQeP6Kgnyn6ktHJqRmXP
9wAZZpxJ3/wDAUYRh/66vk87w7hA+QAzEMfV3lYDbHzoLKnRJJL1Tzda+yes/8v/
MnOr/NuHrYPjIi6iRIhKfnpwlQC7+/SN9yP/SP43suVV5bEIRxdeb9dkemYyQJlS
DYqiZksNtOlM3tuZwHvLP7BHLzQ+wg09UvrSbgPCmZKjXlyB2B2avBDd7den8WQi
NCzyABZRNpRtbqAnc4RZOUeZK06Zk4PV1I0h/N3RCV06wM4lC9/i9QHrASyBllLW
lK1J4Ymuu/uWfSF5I7MmLhKKez46ofbAvSVeOknmPbZRXcefhpzQWSQahllzP2GY
9CeQRDqatfAw2whm94QM6UK0P1oj/ropesSlTdUdzoE/XvTyDflxz5MJGAPVdnyT
r0UNTDfLG5ivprPdPorHeeVuxCunKyEVkjyVnH7HFJ7+B5tYegKHd88DCBn77rvp
Ej0lqZzX6iZMOXQI2d3Avg3ZnjRYuA0QWhlUg9z7a6V2ncBA8rlO7LBa2a1ibV9A
v2I+rv+0tpicKErlI7unsdzEM8NWxZzlCc7OWTOIywpVFLT9IV4paJpnXEoBimTC
RXaIQC29Zs6+owuz4xQlKzV1ecPWTEHJPNvQYZsAUJE0MSnxIA3AMnZqDj8HFmZd
nT2Wnuuvr5UbRaS+WibvKtXteoDO0hYavGIm8C9a7gm1JKPn2gKXlV+mHCchpez0
q5Z3HAWoeAahmEnOcJd4duj2rt04GJP1m/f43kYmMMjYH5xCc6zrPQgRJx+/Bfok
mtP1zJpP8icLpJBffwKctfDjNLCD3HC5SbGCG9n24JNUBfq6WjX5s4vKctnxDlJP
yGBEYhflpuLv5kpQv68kl5wOHXQTNKIKfeoC4FsGeoRlJuEiwhS+UoEDtyaciqRa
chLUOK6AQTx+hAaEOBXswimrPdgOUj3p7XinR22cme2iO9FeKFkgmjwdpYCqeecv
39uBOAtabSJvp9UmPTHEwBBm/dpVPe71lVXQSbuMS/MSiIW27YteYqmX7yGAtII7
t1TxV13zVEOgCiG6WBIGK5MyuC2fB0oAQ2rxAxDDZDRnXRwcRUlZk3B3Hj5RcskG
TfqXJoDl1MRnQR9hRQwbNw9EMDwSNVrFHipgAYNWYFzrSuiRbqRfzDTvEIk2fG6Y
KF/Ohfqe3xOh9UyvApqrpeYJ2TUseVgcgjK3bsDrGXGsEBlxXcPPspDC+RwUx92e
Td/ulYHmd/jE0/uChKd1SXEQebhNFL2sUJV9FKiZesDyzwx4dW15kDW9KJWDUxta
TKus4k12QA/xvqevljraTFYXVUHajcExx5Xfx4haeL1HUV38ngTU6SRoppjE6DGm
9wTjg+b+RjRp5SDiIMtcTTmhP1ReMYm502Oo+D7L+5nVIQieSLrci+Gz9HwnE5t0
rfCTxg4VH7xbyvjtWpj50HcdpaALO/RBElGzdFp8sb3T7Ku1K8TiZIZqXHPIhfes
1jgLHxnklE3sV2BAYlA+56cs7yWqR3Q4cWO2FGzCrN0ddgVGrGRuuaF7vlizARXr
Je3C00YTpqihE59j+a+TQRfkY9lZSZUR9cnTMpsc/DKmXme8rKicJXZWm0Ipp4xf
+fsZZi3P4r4Y+tWOAZihAwuTHbAIz8IExKvQ//Ac8Sqts8dIgT4BX60doEN0Osj0
lyypQnIHEV3ON0pszHVU9vhEAR8nErO6DK4ShppWL13RV8w1saXSoLVdQzy0tfLu
PlQjuI3y1D4/kIHBwNBTWW59ruXZVpdfPSRNrpJlWx4JLn7O++I84+eHHmpanpbm
DmlbYDN1xO7FvxqIiCEx7nqJk7Ms9QOhI1mDTFbKtcmn2M0ax9JrdkZt8LCeoGoJ
aoPpgh2/nfmRUg+uH+kSK9J9t1dtiBsju/YQuX1em2d62M6YtSuPmHNkC155r7AP
j+NtmFgkdqB8KbXDdMyUrxWulplbDoilLUGm6MsL5Ee5S5UaHxmK+g9CEmrS8EwJ
CJ4qj9hfpyEDfG5J/DwLAumYyWXXnOVycXKS9gHaz2v9Xh9Usxi49E7upPi7bDDb
lVJNLsODTuafyap4Cx+U1SuS7UCcDiSpO3cSIwzIjfphDHW64z8r+NmnZfyNyQOo
6cWK5AeQREY0qVCAn0XlbrvTej8mqsKoR+3eNv9oWJ+SpDkFLf6Z9FTX7l3O6QAk
nolvazlDWLg0+XCfxw3yzq+zk82PlA3E8+sLm5JzNjjAnUhmz51LZlhqUXG5FhNE
ijlUUzqyzTH484lFQKpkfsFQDGQSv453xSV+OlVI42bHLY+/M1j6hYDHvj8qjS/e
32bHqeHSICxxZi+HyNPYswXzjp73ol3CQ9hFfhVgl858kJA4ywE8LNIZAPJtLF+J
6vE3LmPAgMJMVpYJESQ1WxQyvPlySd68hvqOE4gfVaWbeW4vRWqr+jHHKEmEgT/1
HMCNAi6cwOYxNT6SQwjM2m2RCSCjf/BuINsK4V/hXR9fhlvq9Ab4D21cZU8NieQ7
RknwMqEwGadNy0FR+MVlvgkjqQQ7F1u3zosYE32MgbLYAO/rrbEvOn1/DbVZEiXv
2Cqnp03ynfp8PcQBJ3DwJH7CZFYm81hs8JaKNoTHuvv9yNS6Sd8ccjYe0qXA95Tc
dxnzvKYwLvLOJqrf3cDd65yB1/FjCYG3V4DBZFT041yU/NNlXWmiDqBbzKlDiXBQ
liQe9JHQfF8VYU59H/Wxq6W8PlyPPx69Vo6pUusG0eL+aqhZsh3pc4Yh0L3C/Q22
5nvHraZZB1roe7JRFMXMGUYlq8xT4NyRt9JuAiODVY3TzrkN8nKEogfPPHLRYybO
k8AknLepManUSbOGZxQ4R52ZVDnVLsJPfWaVeDpWovOSimEYeFoo7YdkPVC3KU5U
MLGlCNmvEq5uhVrD1ak5YnTXg3sFzAFOryaPek4QAmSAkBwxLDVn9Duw+8/MUQTt
iTC/njR5PozwC7KrEVvlZSQ91EJmq/xo1rcle7LquvfIx1cR1gSicQyV7qDN3g83
P7ZCT5rWIN08aRuo7kexRUQyyXjC1SrmaU/VHEKqAHFxLDriO7/EjcEe/x9vm8de
nHfHGevBoUkusNN6NimYEroppqgVjREXSs6Cb3EhG2Wwq+OPGuymoVdD8hRuznNF
2myge1zam/5itE8KioEHbvGNQnl+QOiHMx+1vBWMfU1zSMpRdoiRXF1ZBTapPxTn
rWhEnrCfPAqrGYsB6OfVNrA1Tt22ZNz/MCfAWkaxWzUFaasTfbJ6sBGjbblFVm9M
TEobnNACFXelTqbgdUd4jgOKsWnQ+pcpyIzqs/7PPHxS7jC7pQ6vNtHrEq5/KihL
bQc+GynAh88UsG9EH04OhlsZuK6WxZ4LVNAkKL73OuSV1PXd91lg9splZVjsvoH9
tPzKejgBbACIEkwB3z7aqExN/TR7FGqhQNaHRjUtVouTMsmZZb82zvRvDfTsTr3f
6BhUA3pPWfjg+cLVL8/YVDTqwUOkPAeTK9a1FCchZW7s1W+qOu0BwSpEbUA70Fi5
EI3iLJMVKK1Z9gJhY94DZRqdi2wZ1P6a1qdNkidENQVB3F6HNeMm4geIuutZMi9k
zKUCbsWNqF33riufqqDzd3YGKXmC4XXtO2+o/BXAKEjEp5HOoZj43l6KQ+TBu62G
9ZAqfQoIMYljCktN0zC/KX2EtAzzSGtd7EEeNiYW1+MaimGEqS+m/qZYGRPvjNX2
bo8f+W8i3Tzfny3982kfRN/XVtVPuLzL/CE/0d2E1BzTLjCb2UdWN+rPi0DxaeEB
I+VYDWZz++NJ7cvF48UyLCnVGInxRGjvGhwlUPqSsJmzmFtq57c7AiTzaAiScms8
arvFc96j6VlDANX8PqSutsSoP/q3t0MET/qt6PRI7KvW1HILas62zJJhUQvDyMdf
Q2HhMTdUpFAuXfeyGRfD3T060l6KIYRTGuMEEuNNfE7DZmYCUC9yjoNUU+mvojC7
7aRkg6szGzIhMX0yRJpERXxfNAW8/w16vht/eP+FFxpaNFKy4CIf4bKToazX04+L
CT3cJ3mFymijWS43Xs5lg6Xrj3SGn6XTSG/vONKP3XpSwo+eEaY40gfNhh9tX3Cd
qcHRCqIfTuFmLswm4dz0PdF7htNRmGHPky7VfE8+VimOkaFd+rewu98vkCvDj34b
n5NpUAJ2i3kquMeueOOKZK1y7Ev44QlCG/RGdcb7Dy1nuyd0HjWkp8H83raXbQQS
BvhaBMTYJzqfZoD97X5to2E9wt0i/qlsxYxVpQ4VzjtA4FCLY2LchNa56NtMrWdc
EXptagyofxhMpObPnoMetP/T1N4kHKjR+RDivClqc83tGFctu2mKw/ZpMUXscmXg
POSY+IvV2BzGjefc7d+Q3N7ZVeRXYc2kaxRrGdvXP7h07ZyQcJPUxlSbYI6vcRXC
3eCBlo4z2L3T/cqfut5IjYrZ2YXkLU4VLPAz/F8ktZCe8ZNQEaFN85bXfD5Wo2Q3
U9gR3zYMK0rkyYl5jv7JZr4ZixOYXku2JSIG/08FWdr8oXbXW/khjKvEu/xn6gQX
VHlAPZo/WeVVG2VU2rV8bV/FukD4zPD2Vivq2pzIN50Ua8C6wvfdWGiEtOcVbCQ9
IJy3WarR8iJ/JtrClbWR4bXeROM3JvXMty+lI/1yvaWzhr7kgaV72gmNWusgkBvl
cKc8Fp0n2j3BPSbQqMbMUcWbAKN0rgd7dYQi6gU2iXDc0Aw0pVBpeauiPGwsIOr1
U66qEKihjCTpcCSR7EPO2htYOY97tyDMC73RDA3Im26FySiDbjfzD8e5UOyniA9S
ySrz02cUCJYNqxvzVo74s0IC2e306xHiFb2v6+z9DQa3qTaCBroYkM6Zmj/ngogb
297CMiv/rbqj32kMXHn84QAA3BdWlBbSHWG/NRhvKCROESB7n5r5ysnnoFDDXJoE
h1NttteEXQDeLtSclEOYawehPaGqJYp/FdXRJ8LEm9QCW3Gr+UArxB46Go8hbiAM
xl6SZn5pgpOE6fd8bVgnBlx0LnzjH2gZOFd8T0BIjsLcOM0ylK3rhLIWSo88S6nY
GfOTRxM4YE5Y+DmVa4WqRirlJu3mlgUUF369pupLESXtjqJX+SMTGSsn6v9PA66m
YU9mb+CH9L4m25+m0/Nhl8/B6K1lJWGCZQno/IG8SrvVFu/HwlyAuai8rk+ZcYZO
HMv2btqMnbArG6fOTJVWQ8PhlghgrQ32Vr9W1BcyqagEyTefnCMNfuL4mAFOIfxj
Ky3ALiFMkqH9v/vlIR/LBJcDe7m+6GFVzYvo5YHvu24bI0O8PlF+YlBXP/0FZ6zj
AbdOH5hpIYXQ705I/npcyfrAOnDY1XFECdB2/e2VW+tUkCHb8je5dU+JeaI1KEob
EOCkVyFq6e/aKAjUW0mCLufFiie9+jd2MMuwnTQ2ZIJuXVVYxMecSNIrZjDEDZ2/
1WIfOWDSGBOyofO7VS6Ai1wxvdaPjvlv3/sKk8z4zFZZaJipD9nrW1BnVQ51Rl1s
3BDfLMfAnHMchGWDdi/7H6voKfl3FYXPqfGumOrGy31732BG/fbtgnldTrs20nEj
liBCONrgJAirqk1MwpBfLSNhfRjICo1ar81sImSYkGlEIewfiy+6fjoVpr1zbzOa
qj0BcMqMiiwR7z1WA+j7kOlRx/hSBc2R6OYPcdqsbOV4q8RiXHYOSN9GdNU1vrLh
bD8gYwuU+mcbRLcGHdc/z689nZgHkUf+f3XW/c3CXbFPScwU7Cl9il3GCck8SzxH
mOWSwT88ZGrK2Z1xJHPvuTav+P+bbfyWNnd41Iwo2LOCaom/J9r2DxU2RD5Q61vC
mqaXatRlShA6jFde0+oCLXf3p+jAo2T/MLXcIdonQvabYlDkxbBEuh+TaC+rqCKO
X9Hls+8c2RUqqhZNNwNt0NbmVCF9RrgCDHYKByh5RIpDk1aPaO/6BTgzROIZl+eo
IpHEbOCgymZo1T6yRAZcCznYl4GHHoOOstt4b066RRnIR5qbhUJYVlzqkVxXBu9o
45DbYNFE4NH2tW7ofBQUgPL5PNXocZhy26xnsb/4FkLzjsKqVLY9/IUAnNDlGTsQ
wUNhgySN1ZN8q8bO8bmm/sHFABgYdSSB4koew3K59/ZW9f+nvFkwxBvR7WIfDy21
IsaPMcrUOTc/Ff8+jUD568AzAr6Stnx88C9NEO5f9/jjbbLrS2n2YoSDT2WKJmca
Yiuy0m+g7xMeI0zefJ10/JIlc2qHwdhHLJ0Nn6zA4AMISEYIVB4dpu9CRETvFogx
8NUkjsaUsiaRa490ybxo2LcOV0CFnn5hYjKCzhZSpW4LpPpZwL7f+IaqBBpBL0Xw
k1rqPNNTRU7JcA9YSr021bKotkDUxKYYV6lkbhBX5XM87LnUKfzO24LDWQduTyf0
v0p35QPu3uFDP9xBc0rYJj7nUkF8G9TZa/2ii2ADGsGsCB5mMitnuQgtmVzN1g6h
q4LL5yuivCDiTV0t2UtfYExUsaVoTkgpF63YXFjtbYuLEEW4sf8sXEWbJSKfEU0g
818t6i0klY3HI828GLkGiHwtc8HpW2cjtuoR1yPgAZ5ERSWvD3Faw0a8qnFTl4lY
TpHiKoM8etWRQ16jEjJ71B7Ff8jDbEgtsScq2wwe07ZUOuv3qQaP7q7DLARpoVnw
SZ3MZR6ZFNf5x7ycHvuLc5Jh0szp+ayX+Q6Pb/4DRay349Wb0cr4bEQxRU5fqLgS
jMRECBQLdcFNsC0xmYLSzAP0wJLrrGLZYbr/cI1ks08RJYVbOGm6XMhC3py94Dyt
Z5s1QAPQ7Gi/M+N4WJf1UZzc17sZ8IW/a5DjQLnDSgK4GKedjp6zNCp0hQjlapWc
bUTu9s37SIL3JBwyhBWpHqz0dIuxP25LzX70BC/RIRpniLOhVuFNaOB0atCOCi5n
c9HrcwmNU9UlYxyxzo69uYMxGJvFNWjuodZ+XPxwMBla4LC8ep8sgRUekvU/ziwe
IWKx2/7fEGhcQkCkEC1lL+v0OOn3bzVaZ/AIefa1PvRYuvzbtxP1QembimVO3SK5
83KsAQ5RfKO/3fhwciDcWxCySOCvLuNNMqxMVy2joASB1Y//4ti/m9CV2SxFL9WY
WEtHGb9zCSH+hk4GOCQ0aiDO+EdpYVXTGWYl9SzvssOT8FoATevAvjmHVrpETSIl
0piMw/Bd6kOJ+gkPA91F9oR/ysHUggDw3SK71IJP0YvVZsf7dMXCpS1yQ2F3VK6V
wURQ7rz2ky/m8fBOe5fZuQhFDGQpW8qBG6LyZNm77gRcWiDxez55GSm/WzDyXMbp
S7AMukB0Rx8+7MVR5lMIsJs5/L1/Ac+UxstihVfcnqSdWJTrlQcet1Fq+TMUmTrf
dwNAtOaa4Bq6tvlbd4xhhJl2e2H0NIZyCDU9msvR9rkkzogrF1qFCJ47QDeMl/wm
2MYq4WQsls9NH8W2FgvtBh/RzLMoxJwPxLRDf6XO6GWXYheynC6YO0L5NXm5zvhy
5He+N33f7klBtdLnZG0FwZB31jCHjVVtK+oXlEKIM6o6w0ivEdXjDLdaq24gqFC5
9UER/eQzWtMaC/pdgga506gefBNsYp2tLVORDB3cM4xIEMI4vg7qXFrwBkjFS1yA
kK2pK18Z5dU7G8YxfwWAuTD/Jma3imqkf0JvPqN6wTK9GrMtEfeTlYe7W3DhzYau
kIR+AU/zgIb+kWZH674b3aS1+cLGZ8Nn1sJAXteY7TS9Ub9cJClQwHHQg0gFSPOL
eSMpPrWbW94FwhrBcvD+irLdCCx+xzYTxGzNIqAQ4P8UP1qdc+5xNHoMDGSJl3Yq
OyK3j/rKw02OzRtGWWH4LjqUHrqoWXuC50CAe0xgqh5WAAHz3/lkon/2LoGQAjES
eE5Aw7vPvOOPcnVbVaC6Ohr9fIhVrTPp3OyQcmGhqkjqhKZyAeMWIalRZy4Loqf3
fMyRBhw812ZetGl7A7BDFub0+H6c3E6kRzCDjDWf+b1k5H82d/RaCf9WjAfxUg1Y
pZmSYn55YB928ZriL6OxHVnSD+i1MnX+Am1E8kCUD+29Go2hB8jtm4s/Bj3WZbcZ
No4sSSP0XfTg/rb35ApvEyql2n3zquZA5NtlXzMi/VnK4NO1BIp/2K5W267YbaED
puVqXmkOvuu501QtPQQMjk7oEMOXqjYG7VHrL2oNrsWjGdQXPrXTRLI1UHLzOZng
nNcl53bOuzzGwalFJatdquuQtVLgNEAVTY4qQ9DXRoV2nnivQQRSSkFBgVYgJW7V
TcLgYC2Q3En70P3cBLAp3u8d2cQKWVloCKQJCT2hKvAkZC4mO/Vy6pDK8JojpfwO
t4i0w7MX7jkdA8j6YlOCC8UCiDpdjAzRqjjvS3q2+sO7keQ/LCqbDNJegqKTZUiD
JlH5eKDZlxnRwqn1yJN2e9OLtRSpJ1iuouUXKMrCaT7cDUvW5WMJHoW8Udtb/KDn
zzZBiEiOijsQeoVqyzJ7UMhFdhT2V095cqwHTKfIIdqS8OFHPBf2V0Tz4zh2wMhw
OjN+Szz4Xg/6vJszdLZ96OoMLPebSgDpzjQuFr5oAytoMowuTIHGbA4YElQfbr1X
DL8KsrxQMmSgQbIZPWXUFDMQju7dmZosp5KgWKym3zrkSpTCDm3xo1PAjQAq0CzS
OEXRkmBP+YOS6PlllLfKNzlWoNdSRnYj6gFjJ1xBkZzIZAJH6TkFeHhnzxwouRhu
LPTeEjvf2DFowp28qR1+8Go7iJpbMGiik9SF/Ce1JjKPmh19nMb7PHqi9m9CICfD
9ddJMRS3KzfEBKICC/u0iBetuwuxDrxnynghC8kjnGtCuN0fLybTd/bja67bL/b8
zJaf/ZzZdRiSU54GhA+oQ4QHGyjM6vsCS2IatgGN8g/i9hr1CD4LDYzgcWmQMqzc
OM6WMzAHrL9tW1ZBkdOXwBkZ/1sbEUx5+qhpn4ovW8fm/tD1CrEXdQqkzQWjjvlD
WgYZaN1O6Z5add5pgXPyD7rUC/HiTBiUBjyLzBet8OLxZAqYzjxlqc/7Gjhzb7TD
USCsKET0Y0oKJRSF+VQxa0/GoxGzo3i/hvExVH5aWhlimkNsgffLY2Kf35ihYkav
Q00v9a1WsZoLv0XZvN2ia4+sfghZBADyf+iXbnmZrg2h+NZiM9juTopzyGU2XubX
Txs1QO748+JxUG5r+07Di1J9F75UN8p414J0n+kXN2VQpSVT7jpHvrQEVvo1EwGA
xBrorZP5RhiyrtdeqAy2JhlZGsQtrkRkCHDiBlpTr3FYzgFEa3MNt9XjXYy+EqTs
gw5Rpsg8qbjVzpvQISZ/+aYuV5CJZbGMCvPB79VqierNg6FuU69rUpAgBuuCvBL3
bX7NA+AGkwpcmgHqZN8hLEhsg5DLvXM9fSym1tUmA34MI2tdPJVX/GAwqxnfFFOk
c3Ny3RMQhpLwwnVuYnOZhvpA1RDUq71Z6jLx3IaadlEwDCgp+lMt7GzDEzn03uhz
7BymqNjvK9/qXOcPS3Wus4V+qpKQ5B+C0JnKHlIzjOFKDagYRl0SSPdshXrdn17o
/uTcn0Op7M4Vgo7Vxxl93pWgJrbupjYJwMGL22asxsZfNFChiThN3ndZmWxrxuha
6SQwwbUNc32m6Xbv2dbQfwI3QahVF4C9HfE5pzwhRzWYlTsQQnBINx22z7Qz9vj6
VzeoMea14l9+RUkHsz9Xq8/i13GaTCmqFBiQ3uENP1GnsEpBUayUDjlon9W3sUNP
LcprqXrJhxBK+AXMAkrEXJDQxkejuW8xp8Rj++Eug/I2Zw++lEa4s23NM2boM7IX
j2GuMqY3tUTUpCMCeH0LbuZziwtFQaUv274iekmBk2pKFf8Ym+u4wYrQIJzuvEQH
3QRnDJs7pdNDUxVRjFAOEntRpaUIBe6T6E50OciIIoryrh4K9BpVGE6yhSI4NtZJ
8kCHJyOu8xVngPo9NicIcfcqmCXT9oNRFsqoH4FJNM2k8iA5gQJrd3NLnTpSeNXg
9D0olBFMSwQvhrhrFhLyaSMI3O/dHMTa2pU4d0drOG9WiMUQ78ZxvidnYKDQXQ/g
ygS7WFIQxyzR0eQZ4TGGfgHaxmEtwZ5g74ixXDj+Sv4Bi413zSm3vpp5hPd28K2r
cFwAu52U1HDVseUmh0jk84r0GUhZSld4f93+iFY0u7CJjrMkwcVuBw3lPGfobdrL
QP6NG9N3SpDXwgl92C3Xxt2nwIo0zJ1c+UWWUzPknYbcCWqJX8b1oveXiJUnuJRr
Tmk5rIDmU50hT6svp2zK0s1d64izLvDC7cJ6zfRHQKpsKZsYXuTR3CKIhHCt7Yi7
i3WweIU89uImCL9kEjpjdw8aIiOOIAuv/U8UE6wgolm6gklrdQILVlaeG9Xwx8of
guPbQB2ds3S3LMsUDWe5De3MyKEgMHgb9uOYNFqqWDgBbTY1jtoaASNRMy5sHsET
84Ca32vDO3Z3MF46UErE0pUd0NbR/3eB4GdcYRwGR9hDIuwYqcUykrpQMV6vQTOo
LkyaGdTEJgY+xazhUzEY6vBMCwpID8zm41Fyn2pvMmTJSIyTdmmFTDFltc9sKwx4
Rohn7qWzha10FCXlPapIBlPXZuUk22T6JpINwlfI0S7PveEhqgcOEyspX8ZVPNvt
JXawNNh8YiNyk2pC7mMVqkdPkcD1T67J+SmWTIRkPFg4aMpuJ46Aplh6KiIBHgDZ
Wjq8tGWoML1YRyjoxgGbmbiyjYoVbYh3Esj9GwdwCDkLIHFhftN5bgNmirTKFmr8
g0EqiLTYmGD4Ky0L3iS1QHp1o9XbyNWC4DsLsY7oKD8EbYhuCnqo7WUbCnyaO/Nw
DdJJ0WxC+c4PwNVh8N+JfqDrNwhl13wXuDMtTA4bJau8FhbM5dExjDUIoNePAQ10
mIcyWiCBQRDiNWylOPdkT56NIPXm/YDYFWd/GlQBNvwFuQRhXE+yo514z7YRgrzP
bwP8OzHAFsbkfiktfV6nZwXxAaGbFKWOtm7pZzM62LYaN6Np2hiKXa25OMySIkae
7j/cg7Fn07+r9E4NAfwapa2xw7t1RBxwzPBuTDGixjTDdm18XPJVOmnR5qywAFnc
xyfITaXcPnEdivF78wFgNx397E6AoVKxsydUxEZQG8MXeWmHAtZgvfZSGqTR7ORE
NdfyyMn+h6VGfIsm6ZpU6+Tgpf26cScmmA3c1s/rPuJV3IeVSldXm/qFc15GiQ0U
yjB0kQS0u/nVGIAE8HmmledoDxH69yI60WN+SiTB7DTajF142P2lsWHa8tTFXkkY
HTReZW7tSxASfTDj2AZ7JlojdpwzuM1Ue517lqMoZeh8eBKB6YVxRDhHLn0jXjSK
SpVHxJA6al7PU/JZM0C67E4wiyO5AvWz1bwnGl3vRM2HAKXlO7X8nbfP27TJzvsV
hJnz7+zAFLe4vI+AtJlVcNjKNshzYnn0olo60CjsrLJ64Qp5A6sX9j3nShbkl2jh
lQSQ1aPc8WBZKjlwZZrODgFblFY8URAFpb5nhlFvPY2aqCAqLQoWk4/j+mb2yb41
jUWBvMDsEMTk7hPP9kjUd359AUbOIPmpCjRQGa2Vnz1t0F9xR9icWI13uSBNoeGe
9LShQI0QUMyYuspKcCCWy0hMe04q5e5Lh4zlffHywbkgD6KnTWcjgDRgHkqMEqpI
i4O6Kfd2O1JcnWZ0QBAZKHUBTOsvnAle0T/lq8SXzC2/yX4HM6gTM/LIe1rQoesP
hQygKbu5dFuVbRfEHeoDKU1kNY9XYEmype5I4YGO9Wvy0zGsTr/+X9V3+keMV9YB
IK97FBSzZI5UztrEgfR+3+HeoBaBvE+1RYXebrOymhwhM0Tu5zo540QU0+gUo/xn
9ak2TpgMHud2qHFXIIkOiz+y9t9eX5oStCY7dF14D8s6ktKhPm49XQt0HtUlsnZK
kq4EiV5ivdsmoiEywsvgiwCxOyqwAE79lVeA3Y2LuOzdVhuU6LrlOJ09rVciGXWx
uEp6966HnYbEr/Ixig5mK5EcrsSeti84DCspfDKtYIb+960yjO9V8GfCrxwhIdrr
DgdMMHgrW5qFThXNalsdD4p0MH+E1LwSTfaAeRebKpImIP1nHbKbRzEt9/pymT7j
MTbrV18mGlfmHjn3VQ6a97+XcKSHmDDR5/gs2HeTt2wsSow9RhrsLjdhWkgtPAsz
BmyinsJtTkQapT3tampiIBtWHgvV2a9QwQ2H1wSU9Dz0Dr+keY8+04o0OWWivLlE
kRq7/bGZHarTKw9KAv57uTJxq9IBqNdImiocLikgWhdqnIYWPcF5nRURsLQtAZ0P
FDt4BWYaYutcCqtRzbUkwhZNHg93W5kEwQPpHixKjmGc4lfNtil2420Gznq8a1nE
bPdP2I/r/tr4RUXVQvsw6orK463LZNKOc2/vt3O0ZQnB7+6ze1MZs3I5PQn5GvZ7
jodMgNk21xekrsKfmmCX/3D12ISvnMNsuYf3V8sZgYeSZxPcA7RF3oLwP9f6mEM/
hRNgl/qiaIGuoS8znFYA8ADXZyzuaJHMmzQlMjC7iuK2OQOGcsv4NtSqB5ShPq5i
gcWMZQa+V7rVtJKlv113TjH41KjimQkwj0TZV6GxL9t6oJtKWzJPfLFf0o4t8KaV
X8ZJoe2nw6C6hnEo7l0DRH16O8fXR781HAmN9HHoOvkDEgvzIvnQvy4B9oVNHodl
UivmQmAfFzspljdbdEHkeHKg3dJ0IoPl+2nSikPV/iye1umUkfudgxdci7R4mjeQ
XAmYVsGOnLb2319aXgPtM73Jq+EgMqN6wJHvYmxS5yUxdUYB0FpfbYYAazZlNS50
h8xMv0ffZnvNq4861iZdy7DO5lSEeQ49LvMVxxNpllVWrRAAEYZSanlXfmoVrhs7
Kne7sXLv7Vx7fwFNvmpE9xBAqWZ4vWxDQmne2e9izz0jGIBUUq/6Wp90r4aTYYoW
rvnt+SoWIn9zu8JZ9HRCchhTVJP36wAbk3FnffMG2vNjsWAzuxU9HKYcfJ739zfo
uxLME85gaDYldg2yrLgOQCMVm1gBLYY5MdZGxAMDmZdvGGtERx8fkEWyMCJ1wlj1
1O6pdgoYVX1PXpxzMh2nTAJU/49NLT6ZBlM19ICozkc1FhvFy3J9a+ClTGzix/i2
H2I3tZLnfU53hIzpccpSuwLPLeoj+mnan+k+aEsNikWvTbnHkyAPTFG8p6YFbzMI
MGX8Zi6bm4ZLwG9/28qR/JKQaUi0XADipg+xzOAVL+3wBmfaJBrgFvAx8DFg1PFL
D4FrR3XQ9NhYjM9ZKPeSbNSw70nnvbWBUNDB5+78E0MmuiAG7LfiCL6jZbAjxP9f
KBINt74593WOB5UFOQwp4cHCL1o+ur14odHDvZdDWeTlb7caaH1r0MqPnYCakTSi
3FQWCVsJ+bCpBQKUWtOpDR5S9JROOE4SQYDwNU3U0z3kQPRNwowTJWIgG0gmIfDo
eQtDFTbIWmIFxKVnN/L9W+u+963cSPfHwkP3Sfi7XbRv/1eSQtSgDezl0qWWvdyk
eBf1SXef5C+AT91edglGZXAjxkslG73++Jxj7ksl9wNvVYzG0fFlbt0Ww7P99+0D
GlBaBraW+xDDFo27q5hqZNzphmc4VN9Bm46aYP1nRzUyMnXLBLPDqX4RphQXyVa4
n+TJQrIZtRkSj7Nn5jkXmv++uQg/iudYjnPS/dkDfdG8bAy33UrgPzcsGCfD0ovC
P68/le478pDWQOeT7da4B+TLvRc61yKILeMmk3FobgwU3fFFsI6qHgTda+wzn7D3
1vQUg81it7SaF3RxcWGZ4E9dnXdCoOu/T0xLtsDBNYHkTCthGgWCiBCIlpz0HBQ3
vJYU3/++CU0yx8HKF3ZATNolQetpBEkvBGclR6jsIJIwBC/Wx5vBgMxudug9me1i
EEMUMrwYcMzI5KmWFrIXHNxBq+J++541WZzT8YLnFdY51rWEzIEavd283B6+8pom
6LlXLqZFYBcCwrLT/ibUzo1K8ZNjekC6fHP5uUWPCVDwqy4bMZPkwNkONxExg5/o
YSwCM5PdVzTDtueXXugb8PD3M0WjWgnlShFLUavr0fN6++cQhzOWB52npD5wODSv
RiDgrgvS7JghNqY5+iApIIJez3tRj+a7ia13z+p4ZHBqgKCU9IyblRjTJG4gezhc
cktBCvSI3xgSz7M0ZOFNrovRzHWsXJ2M4ZKK8Rv1oWTVpB4kDc6HGxHJtz17jC4y
pUFKQF3RhLxO51SVQZYzSwyq03BkCS9uF+zMSBee4Di4EQL8T9E1vW8hIfx0xETN
iysx9YSbuq0ItTMOV78DBPE9z9l0fvwFnVrAsW6hT6XikfGjABWJbSlVYcFKqjXa
zuVENcYvklfHAPQXdgOpM5v+bgQEuSFOJ+wanDaGmG9vaizyhbllcknOj+RZBvKz
Qgb5hw4YShBGD1foJIgVaPskbuZOvO6FsSMjtRKRSGsXmOSR9S6pBGWEDmtmE9Mx
IVLzAX7zhpWf1CJZoDQSCMJvBHyPLYaKDe6W4KKqEocUAetV3i867dLpCKdT8U9B
ppHqztm1DFfpWSc7gkhHaXdxm42051TMja4GtUe48X+wmL56xA6DvdVgvTA6Th1B
jOaUuPhtlFCGQB1qPkNagbg3dpZz3Y3cqVYZEBfMw/sKA8qKWng+fYJKL8FvriE1
E4w3IgezkUmeTdxMvDNp7UZer7HzHo5oZRiSo/hHyjn0Y5Ck25XbUN/TRqcmWbqD
FvmgcMJ5XfOdAVrF+y2zVjk7Xpnf0S9/BhLV83vdV1UEihvxz+KxwRLRAYdYH8pj
+1RhzrgSoOj0dFc86v1F3g4QrkYNuwWTRB6cBFFZktKqvSUpCHzYLBPZKcBw1uQ7
BFs949X8Rig0n/Pddgv5qiKVpmUHr9POjdT4OTfey11+sQO1Yf1RiaGSOfIoJFH8
6kaTTCiUE1fMt5+T1NPbBQRQRC8qEZ4do60RSWNNNK8F3CjOI0jYgZF2Hlk3FHPd
OGRknU7ybkbmY8rUVlb18791VjNWLNXfOVkmA2lbueFT8mEyg4BQQ6a/SgZwC1LC
hdBybB+QWTQogqIjngF4v0utF+gDLW5xMYC8lN/gR4iaLxg7x3HgKCQDXnhxG/SS
Fx5yOSLWT3FREV1cZ607qLQUX+pLPlMcP83ozrAl9wiyHsEG0D+gRNxK94jyf4HA
E+SYU/oje0i6MScCixFAvqjws3Q5MHu5qN/z0l5JFMf+1yWh4zaIuprbpKMGvklH
p5n4+0+au/dlIIEfGKGJNAYoCwrhyv5K/BPwiZ0yhDjlBWKy/cdN2uFWHwkPlAcu
b6wvzQASSP7hrAun/sC7qVlzIh+aYdc2BlpK70Vlkq5HR8wIaxOqbko9lngVmZQH
GbjTdWCU3lP+dlz++MWmLxwqnc+tGk0DnrNxxBI67gE/mXMpq/9QDziK5oMnCn3b
IKC8dpBDvLI37gw/g9fkS5ZErRkKHyiFt8H+WD5INLQXGpvxykGLfXERaY5/PAux
TdGvRG+RLeHpIFusAtygnysmegLBqFs/1F8VRskWn7FqkrpL6uZUiON5J13JKx0w
sR9nQWoCu1uxwIer52cFS6YfP2VOixVR163njjKbgjPToFNOVufcELkFll2Cw4LO
mURitdJz6I/pNjhrJiuimDEAIEf6OmziGnMO8a/E3Abnxx/M7TPcHNReFKZZng76
uUWwAZ7qovB1N+IgQj+V1Rc6BYMv+/nZkpgvHiqDRqlyLYRe5zU89la3XZZNZ9xP
OQah/GYeMqnZmtQJAkjTVmUx8HTBgMPjQf91EGA13LShRWWQzLccnrKQwd72zqz8
hfUkSQWnd6Wuz1FsenIvifMMRBEH6ojsByCcK3qc34IzNXfoZ176nOuZTGk6KUJu
bl9batV5R7xBUcQMVorc1RZbOfv/n/wOV8ehuSds05Wr1bqLnjPBKEpph14SJiKg
NiNDRi4NjM2h1nPckY1hd8LsaYlTqQah8XgKjxddJg3+r5ZbDNewmi7W58iKGpa7
2waNg9gCRIdEs4KHFi/ymDmEd1u/XaWjYZlYM2rC4Yl0nIG1SB9ZyNJGfdbPxdiQ
iE6OX7/06/t96qnsAt/ginFqhONy0c+8BdcXCzF2++4X1Wnn9G5SkDGyZ058uZvB
Xv47O2mtkZzQ6uOY58ZQc1MooH3saN5DBdGvoo1Era5ML8dUg+ph3w3wf+BV1xnI
p5WViR9Q2KMw7MmT61u7OjkHVNPG2XeJcqMyPcr8Rd1vF7+Z7Qqn3FHe7F4j9BXQ
1vExj6aoQoeDzR61WETqSg==
`protect END_PROTECTED
