`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4QMNzrJtBJ3jBwXvoZ3GAqzLq0X7OTWxu42z7stfuPty7GVdmE97CvAbcomX0q12
K8PHlPdV57+gXSOegAo1KvdqW66xzGt+hAgOzeGAe51RwHrarpJvXJ7K6F2MBeVX
El1cXlrAIU+gxPkbjyyX9KfKZZ2tGDytYdZB4nQSPhQkUsf1jGjfhqEJjkjYShHZ
WJZ/pBBshDGWCD8PFKD0jPlZI3NZFQdcJVqiKyzAcapgM4Y0UaSHEVH8KKTX2F+j
DwTNTvi13Nh3Bz0OfTawdGCpsDnv8p2in0wu/yjOuS0V+BMjm855QINp87lrRqtr
VoEyPeGLsN584y+hM1ldHnt7auS0NSJ0OhgNyolwKYNQhvfDja7elQ5+tdrN8w8S
/V5AJURGPN+Cws8ErnIHYwA9sxdUB03BDbh99DkDGagVkRwGhYiXhrr07HMHUlnw
gmD+6JC3X6tbGM/0hAbuRw93/0qTCvH1HYyAzewtUCEn38arF/DL+XwBJYMWiICW
+ZzNsG+aLr+y+vWT9j3z/UKueKLwu5LZRhfZ93x16jhZ3MZcXpQLDWLl3jD1t7MW
wx1752Ud6nCtVYwLI2QUg4n1KzT5puvwhObmsqZTrBwaEnfbllJc3k3hqmEVV2cq
2RrqPi7omryixXpUD446C50m1mNcFjTqIA+gVYFed/t1dMYtXeLc01jIHQL/RbuK
OVnQma+nDo63TAnqORtTX8YTE7EUN+U+NvJFXwVKyJPaAQXPQb/njlNfiTP/FOi+
NCaNTha0BNp+oudV2Amqx6YNrrLvdgZPLuACQW5K0mTzVc4L3aQ/OkXCo7Q7bT+M
vtq+an2/CttlcAQ8uvDzI7nE63TRzsdZc7lEz4nTgifJnTKVuepUqc0Ks6OUOZ8v
uAwviVy1cgYHjw6+wfi+uI0T6F6i1XMQGxL6BfPKftDnpoeIQAHWlpFp9+ydNR74
F+e5RVdxiVdc/NGrJAoEt9h/+I+YFzAtUCfN/xMVOEzw6wbOwHKPkoI1AnuAEdVA
CiUM32eJ+xg4Oju02k6Be/QbusRwHp6aGKu+YBKcRgTmyLrvipRbjK1Vrz0SfRzC
R/Vic8yOouz1guMQigGxjMewHxAjjc9g+FCzuPJfk6ejLbhxd6O8PLjh0geVVqOH
l8xQt2IPPZJmdKmVnnzdxxV9GnzO9R3wByGok1MmD1vfo31tQ0DECIjCSNNRd/5d
Cf2ksLsmaYBHIE0UNIWGGaEmyAl/ct5ONZM/QJQL0G6nQWZ9w3eLQmxiJ8WixmbW
n/FEFsbecfTTIUUcAmPReQSll6BXkPN+F+wIp4xK0vZM9pef2mufWYB95RDDGp9N
8xCxckqpnSq2+HHa5PYc5E3m0YeF+I9rEbFRhapHn8woZXhSH4vlcdKLPLw+8O3s
9BOSZ83ds15UwMocDR91kZXwUy9itvRg0ZpoRhe5kIcr1EsZ9W6qlPBhZ3Czk/Fp
LmWEO5xtQLM7DcYCiuDcYA9zzaYK+IJpHEGrVF9HGddmPkRBa8nZlRGUpE6SGTAN
/RUc7FWcWsXRmAIUAkXb7uEcLI3XsWHNlOBAy4FGtIg+f7gZNU3PsyaCzMpjg23L
OR26dD6gt0YmWRMmFlbAu8sOU3f6U/pnBoBUKEfYWV0D8b6K2s6e3zyTid/enxm8
pMX3a+LCvzzoplAypzq/BFbuk2/7nTtVGJ7iv6ixhoBMmy1lH8/pfu+ZWQ+Wv8ke
YvhoRt+12FKhL9guw1C5oQ==
`protect END_PROTECTED
