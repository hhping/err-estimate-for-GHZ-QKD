`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vaVJrhXh8VSp9zItsX8b9fybONk7MlVIH3qvVV8S113BqpKRxo1F9skxc9xGMw83
+hGGY9HE+Xu7fBmzMJIYb1+ZvECZ5zyFKC+Q4zMtyLFTap7XgGntQdtp5xI2Qjza
dFtJKuvRgiEJb9vhkbUaSgbOHYqb/Rc25JlPyy/i0aXYoHdlvgyQsQqKX8pWdhXP
+h8kNSwEqGn81mk2Ue7hQ9uMv6EQ1/66eYh0/yMoYqRKWmIjX8FxFFnp+DeOdMkZ
0Y6pUuL2Zbem8Oy+67n6/m2U+5KIdlytFrclhFXNDTTCEpgQTJzFPJbRRJ3uGG+i
Dx0w7o+AC9taSItZDHoZhc1xDT/jdE6Dq6Ska8GD+CDbnTXQq1wCRRhL8yVp3z10
I7FnLj24gq1Xnw3DfBNZYEHY+j/UgKulrLOr0S7N3y9AOt0MhoVqcbAmL8GzNgif
92skxwj+O2svc2FRYCqN0aIt4jTta1xmcP67macZ+lEsU9uk6EDN393E8lBftVos
ZDc+Pedwx7HlL9EWrgoLl+0EtzAcHYOb/SPsQIexYyVkgN9IWiLvbpgF5qCw0HYS
sAOxxhNooSjIxQ31PO7D5sMcAKX4S8KJJdP+88+5Ik8ElUZ2IR71nLYwRojE8j04
hiKXedsNTo8lpKdJiEY5eK9O0wPEhPIG2Ufck/PO+QunxLduwJdxbXF4pSIXRAWP
ZrQxlMqTHKOlz0Vdfd4OgsZI5B4rOhYqJqnoY3lyVHtD+agWpVaHPFsa9/R+ugS8
DnjQr7SFso2txOL0XLmwrq32QcFbyRRgV+YMugftdlpWe6yR5yLvoV19MjAdcdIh
AE4aTVgu88qNehVR/eMAu8k6G3K7UiJ871pL0RgCe/nmJDQH0UHbzsuVAfKcWwun
5dxoQpFXsvs1GvoDsL4AEGSi7LMR5d3EfqYc/7qUpzeiyiRIayIuoKgb0qEkgN6H
NR2ebCyf3Despaxn9z2ygOX1UsgcxRVp+r/YSFRa6FAM/1Tbjl0lzaQfdLcx0OU9
yHmjqQP2iaRcDwAcoU8v4pC8pa/wdbggXYDQR6CanD3Pkvze87PSw0SEp7ECtCDZ
mXOnEFAzhHQCb0gpAhsf/DWFTwYOdpKbFX7Td+dBfyvvqnVi/8aQfUtoLefkYpKt
axuxaSqUEGBee7D/Q5Hvr72wuxEY/L3eQIaL0vnLeSFtEcZl0P4y/Qk27YY+VKMO
ecf48UscltfXvpRApV1AHTdQBYHJcSw0K3VrzO+V9ecFpQYXhBWcrMbEfefAcb0E
doEeSZTbdgQyjugvgLVxgiBLsRWHlLfrmmNFrk3WD1VWfDzAO8CsvaYqVetNzzTg
p5cP7pcoWPHMsBnrxAqcDCPCasgIDmIoBaaBhjLIfeYrc0bIYqbTnlovV2Yh2HzZ
LrKQbZtauHv9IuyHkBMtkv+rHJDEL6Aw7eh/cMtHPJgaviy5UmUTm/XDxEd1mX2x
WTvsPeM1RylWZk8Ji/lANpmfE98lja8aNcDRrPrAVaXZQpwDdMCCUb8ALRFyWcZH
tiSV2ZeLtogFCdTZmAje9uN52co8h0mMuVUq32eHJFPm1LniSQJe7qQ1Spi6UgwJ
HFFXSrpRInWymh2hnASw/e93ziUt6U9gJQ2DyH4ZLrqNiuoMiMsKPH+7PEXldM6r
OJroTdGrS+igR7IB0jmkTgoi34NHLKqI/Hkb2Q/sGdREuC+c9F7UPnFurE8V82Cr
LakX9zBVVwlhiEYPGX+gAEvVOXOzpX6o979Ns+dz4VBhofHyZUAZMabQx01io6yq
bWhn3rXlZP3nISi0F34aq6LHSl7U16F37pgOUKY0XzAQuBJfpo5VYFfzm+iU1Htx
bZBImrvph5lxeDVMJK9BQJt9mC2eNX0vnPDcf8TT/CNDz0i1OZU4AgneBmVP/HhQ
LRkOsGVYzg9HYnlpSLTOC0QGgTcaQlXngEbskZr6iiiSKmD/yZJJIncuWlUYXJKE
/dUROXh67I7rJs4zjwHD8S9XoqcURb/xNUc2eNIh4ZaHpXTU7e2S+7Ql3yNE3C/i
dN2+3U4Z+VsRFCu4cpT5+phxPuA+iLTEN18PMEpF7nQpBYkMPSy9LUJR530GfdPE
Qg87L9nyNFSbN97SADFD4VibUG+ZBQFqPbIjAN05VGZMnrSNEu9QU5eMdy/zworf
Eiz2oAjT+y4veTrjkCBeEN64BUXjLxliMbVubOcV8mS2ySpLDdatONmchNLiyt3L
yeFBeBK2Fp8TDxOiAwlhiHawe7/BfBufssHz0Kc+E7PYbU7CRbmPWJwgoetmd66O
NAm8H/cpX6io02f/abgjTJDX66VnADgIJb7oQ2u0cwMVMF5FEbjNJGEwaS1AMZva
5fQML025BAmvKSWBHAiKjkgthw6HbDTZA2I1HgCFAXc21vnnaOzG49lhfJ/P/B1h
9kh5xrUNAX5PkjxJfut0DeEGWjfkYlVjjvK5NoiQRf/M08hk51kNwBZDBgL5Do1i
W8cUs9FhMzRdlUnCH+R8ov/0EzWQSEQYj/uJZkcBf7opGn0QjKqVPiNy4JKi4u0L
0pGisLJF/jTUwKjstVeOTjzU8RqPAgua7W57v0S1CaHc4jY70MKlCL/3CnIkB+H0
sczyDW5d8tM+7pBfgF6eXQ==
`protect END_PROTECTED
