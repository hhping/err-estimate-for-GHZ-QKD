`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
24rOJ/0a2UG3MiVWZCfsZpG9ZR9o2JBnMu0m1YQbJv42xO/xRWepKazGmzHFXnxq
enerH20hZCm0hSklcR3ozNhYUn29qepgPwTm77lDi2KYnGA1iyXTja7QEKA6RJrg
HEhUbLCjbRFiGkwwBnu1TS+QeZ1hvUVSorbfUq8KrxK/Hv1gyLHu0Vib8Tvl6KLO
HJBA7vOUEoOBYV8Vo4W7VA1VfgMg4h+wj8hdQb5G9JNj04EMCwlIgUSMh3eRxs/i
OKrg0o5MXZ+NuLuYTq1lEEzkIzJ5MLms0iaq7aQJ+faPbJ+GMLvVq1AlGd1kM4hw
HbJnFELfslkL19/0Ahscjer0/eNSBdPxVkYYZM28m4DVL1fV6YGeh3UQRSn+AmE+
0wsrNb74pJimQUYT8Wku5lETuVfT0WKZ20LgM26LI+txd+8M4Vul+qOJsITToifA
oexUTPUZd4h6hCo/+WxvllNA31dSPUbhO4iOGvvoOYUDqvNOxfFQMSRmdcmhN6QD
YzWvrqbUMHr+IuyK8QJPXsvXeCiUegrmw/PrytOhhDtMJNUSoZyddg6V0dwqE/P8
Dhgkb5Us5h55cqIfpTito+4zoi+GR3Rjy2NqLr9mY6L0i3jxkLIPYzq6I+ScXRsq
wuYYmXefbwQxOXtAl/t3aKX3XPNG0s2Y9FUQt6i9r3IPavoelOAuCZsNwI8qNUQB
XJaHDdCH+BVcjAldilohGp1dcYXN0C44SYWxLyTAA7wMRoCa6dgwtE2UTXL/lP0m
ARGbexznPTIH3vAK90wCWJGjU4PGUeNGsvAfTuLAkkRH48WOVm/AE8GeNmPCwz+2
g7wAZzq8cfjNKO5zyo9HJUDLxT3H1krfNfre7eZweVfdJ/Th5hK1fwdAF4x9VnLk
oc/WSOfu9rpktic3KU47zreBcBSqC55QigvzUELW7tHqpghXKdzZm+GLZH/imJSK
CZExb3rzP37f+/KkY4BVt72aABYS1+7tR9TB9ogjUmub7Zb9w5GjTPae5+ynfg5Q
mLc3L8cWV9VdstclucElau1xHKwNeTU1zQARFSXSP2nUZ1GgcRaxoA99HESO7kUy
JereLXdZrJ+z/nxwZt+GvkeMem31IeTXDZ/yqkifDtxXdZ47aDJxpQOXcPO1s+kC
cyfV5OxsWvU47GHaGZ7vfYRnO8NJI3qh3lwinhFOGXqQrLwcSau0YU/kKZAKDB9A
0yC5NICbxB6/DqU+TaDj5kunja5ScQ2tyMfIFNgh1H1yQyM1PstRvfoNqBtG0fUN
DuVl+PKOA6/G0ackg5K87t1qhi9e1Y66h22Yx8NjE/comfbxM1lMlHAnJJqoK9eL
tFRwscWh9eldfegx4n2jRZ/kcYAmLtbtj3GjnVH34Y5qvpPlTEepTsnEskrHR9V1
Td7tXXnbtgQIeOZ+CRe9Wt+4LpjBO1TgU0PJXw5H7gM=
`protect END_PROTECTED
