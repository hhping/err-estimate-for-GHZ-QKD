`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wTDe4sHgLXS+LLJgCxp4brG2HI8VmsbWSpba5e+RoOUvDE0PpUsy0DxfcVz5NILd
4xxJwiONr42cBfHQW9cd1NIftXZAgrLgmWaLblMEzDGuVuKoj5x/JjceaqBvruzN
pIjCNRneKIXoM1zFl0mJ6QKOFDk49661rxKHAOtZqI08ZMKpJs6bqnUTNx+CuClD
4tiuRKu0/sq+SfpM5AwLf5L7KISA2AcYD/+rLN511zRVaqiZWT3s8KMwWh5FU9Fg
zlR5IEVNcSsgqSsF9JynDW8cMH1Or0EL6A59kqBUL9bTfAcBGeer/3lBTu6PLIga
b2M3CESPKGjMLuqHB6iRzNuPAzUSqo0qYWJ2rUFzWUwR2oMVkbY4Ly7Q7xDq7mdw
f3Flu7MYlgEjkRn6CSheeSJkMFvQwuCg/oJOuy3TixwTO3X2qpzgHvxnO8iePkrJ
yQzR/N+1+b6jeF6ooetybOP0EBeg2+RFybh0oAJLz8Uiqw7h+9xnOiCLa/FXom42
YvsNn5oQ1FCBaBLTssvMqjUydeszH3KqORC/ntuNuryhYvWjKmx5CvngAnO2jcyu
r14jHH7EEC71iOZ4H2L67opYzPeQCME2oEKcJ+lyefoE2bBwQuK5n2dakzPhduQk
E+IoYOcrHcDZAGv3q4I5C1/OWWKueCgWfhi+Kuv4tG+TjBhNB/B1+qirf1uGLtTP
ZN3P8nx2oLAPenHCOP3HQwxd4hwZej+9dfJ/TEqrJlmrdPuwcGr/qhc0/WGGc1WA
GP7e0eDZVoJTKf5QHHwS8Zrfp5H6PK64ghgvpS8fueKOmoSMxXsDeDcJzYglK4AK
m0dj3xbZvIs39XXfpeAi6o1iLnOwjGHpvTwRpfyg4PbN88r0VPd0rkT4hH3qLrTj
aCQm0FK/JS/5N1IYjFzG/sMxMJSHJeYVlFHvFgrQLJQFrrlBaCFN3we/SPJssmA9
wc5+3mdDWv34m4lbLbpypo/AARtF9IWLMm7I2be3WCD77IkQ1BDnDy0syXgicSnz
Cfih82OaGFwgOkkGPh7khGhFRt+8/pE0bjcUR5R+oBEnAUiixWPvcwOWDO+S9OC3
H5tmLm4uDUWbgO4bjFUIigIXfhToaTW2bJ24b76j3qY1G+bSAkbgarkK4d3sr0RH
3tow71uls1ChqBgReK5HqmUYU/5ONZ7C8HDIRCXmFFOq3Ffoajp/dIBqPSAqeVX4
NhzmhXufAcGedgOkEi1lW/Q+KHdG1xl0ux5mLc060lD8GUrcRO7lao1VPgFvJHZm
g+uMSgSBUn+bf+vssjOSFuUix9gkM9yeiJ0jPBhOdBPEftq7be1biS6daavfnUaZ
kMGudy/qQpgWaFIUGPK4BsR1ztyccvsQPff94lg9WCUv3syG6ovgPMx2BRD7PwKG
KlwjzPLqL4ntdWOpfv524Kd5tb8OtRdus/2w0yAxK3KGOqpu5uLdF9YQpJKY/9N6
O174+RbT5e04OZGjNwkCNtpLk7VPLeUJuRpX4JX9dU45vpU9s66dcKe68R67sDZh
K1Ap8X5z7szr3KokgPA+mE6v4wefLIpF7E9/GVdfWr/DC2oYucDI9wFzwl1br2Er
Z9DVWfdth96tuDf9VfzzWAL8byiH8rMzBFGVEAojydu0FvOJVEGs5TZWmtEs6hGp
J+OutNGEPsMTYWIenVNa90UhDb3mEuXcEV2ASf42a1ZSpU9rwxQxXZRO9IOXmb3e
HAM1kdhWL24zCln3jLMdJjOA6pzBPhJAQbeD7E5FC0YQYBn5AlEQSdt+g8LO3DF/
98XlMJYF97C77Kv8EzKw650iV5UWLu4lmnT1E1FByMcTHkyNuwulWHJoN1+1xOMz
0fYRcImtnHsHMyTnot5CuvfEsRs43/mKRAjeAXAXswMdibUpsGNUOiRKRK3gbP+g
h5TljPNoHmGc4KJinmdsyg==
`protect END_PROTECTED
