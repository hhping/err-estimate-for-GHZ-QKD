`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KV0HKx+qAz7KbGM5OlETEi9Wp4V60xcCCRbG7x1Z0Ycq6ZpgJU+rx7DD4YyoWogJ
+It3F/YXvNEA38goE++7hQWRqUYg63mTysjOEXbwl/p989iDNyyZdR8bnp8P+0Si
dYhtAPBG3aLiW+vDcgleyCzP1uh6BrHaObamdwJRe5mY0HIP5//WsT8N/3vzK9zT
7s/KlCLygnmfn/zaZyVlqIo3s/L1jIEYdUunC8FOxUkojni/5koqdVHiDFzeRyEM
wDpF0H3Dm45iEQc0ESn3ORwbbMgnFrLbqUPE8NFCrT6m1VZh3B6hzxNThDo/np5x
aHYPWYWPFEz3tzXiWuDey6UVYsHQv+Na0Qa4M87bUzImsVMmT0AlSKHiWx+ep3AU
1CwCs0T9GdgXsP6rkYHuMwiwcUX1RIC2g4Ptvf0MaYbWg+l3kUWaekf3gvA9AGHG
f8u7Pr5N41OjRgRVx91p2sFuF9Rw3fWFmyx4CVKPQAiQdflWFwKWGxiBXEbSATpT
sJgFDD7vz3DjZKwpchmDc7wfaZGXqyKqWsj4eSBG1sk45tPXAe2N4lDGPVjm3Jmr
9joJ40PpLfX5ezQd7R+BKCTfvdRrl+PNtn0jSChSsqaKEPqzyWKgZg9qgDSwefk4
Idf8ilMdfb+aacVd8Raypg==
`protect END_PROTECTED
