`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c1xWB/hUBoqLYKlOw90frBk/9rYaqVv+crpCxb0Rb9me7VbyAsa1ishsj4xHjHOW
djIsXrk6CSFWeT9fgc3UFKc/6PQYKM7Sbc9IeXvMC0H11zdM8TZ7RYjRJb0aGZLJ
a/2v4Sbo2jmwQ0bCyyLt7s8iGVrSjTrXjxFQ34McQ/Pl+MT7XcMULmUvMVzdb2Nr
WB1DYHFg8J4o23CIiy+VXCszrcdAfRpANfPNCJuDOaP6WxGdR4pBv0p0ZD5yuo1s
nGpTzSYoFnH01805YgmHHS4Af2bKtZYXeqQl3rIGnuxehFt2CAm4bqKpOMvffzKo
xp/46wi44MPZHsCoB5fwScbs9Z5mqPpWQ3B4Uo/4Kvo9u+yA2rb/SS8TzdLFx2SO
4WhfIJUpHrhTGd8eSliNo0haS2O0oM4sc+CW0uoYY1WqKaSJMTihwHU/YJfppaTs
v/V3p81b/lpS7Z4tJoMqHIBWiXQ5pG4Umx8NaFfcRi0x/CsawFrN4kdbqRlO+Rkh
Bf1VjgesoD8jBSjmB3WR/WTWujg4MEJav+Il3YX+DQNEGIDNW9B6NTvxkbuogc6w
7L8mLZZi4eTR1BDFtXw0ptfG7MRbA1I1vWJBy4TDMJ3lTracBc+T0varDAjJWauK
Z8GxTUAQWm08wcGouQ0W11ewQxo/MLQr/+4D6OqG3kNoC3JCztmFdWGjk78t8isY
3rhMNeeuk0fUS8pRLZYCAUYfIc8CUll2VWNTj/ZkIgow7V38NLWC1aReD2ZbD8oO
gm5NversYheGEDNm792mPnX4TwbKIgtEpjQGPIL5vU0NumUS2Z2nLAXd7AIfndkT
Sk2ELENS1KkEjC0ipdiYw2XvsyuI3SEApDpG8E7oQ2INwUWBuRRKK+HOuuvG2Bmi
j5x8MGFmnN7KsvAnoFFdto167Oml5XA4RDvGCMjkdHfmfwZNQeVMuIgcDV74zgcf
1XcCP21mZXLXa+D44ksxiYztrBPHKzNGDWAQcNC4ZQ1yf4tHTGC/IF2hzCxoVbWt
aad8fO7n3MZWzwXtZVfu3VEXduRcBOEm/9bKX/EY9ohzTCQg7HrTtD5yHtxqjOz1
fjh3vFJb5iToajvh2Zcurn7NL0mL+zPL13uGFtLt3m5ewepWiRkg/Fz27eO+WC6z
N0K6K785a1/462DqlwJDOa1QVI6281B6oik3DV1YnRzKmZrjkGL5f9/ZRs9TtgJP
/wuaINk7B0jHYDtvQUz1N/A2dioCPdTywhLqe3gIiQRHREO3fcGN86ZCPvbDlSg2
Wz9WK7vqFJu+iTJTZEk470B7ybce2RUe00ZWSOu5jucEEYkZj/ZaNHT0Gb/AonN6
eKfQlHVGTr+XxDrNxdwqGQXomGwqYbnZzx7W940syvCNgedFNg1Skg4s6FrkfVWu
5/iAsDmUJMYlJ+koTxYhGYyB4cWCRcaMwsBEtQJtLQ6ODc7LeDk0JGsJQfOswNnN
gfKPzh17ljtiQLsdC/HidCVSludZ1PJYbulB9OijOP2xEDB8NhGJ1pHb1aI/v9kD
GI95jrrVlsMMFJ3pzHw2Qq/mOjIozBxCEg1YaPSlh+VPrHYoHia3pXIDE7mnvmzN
2+1ogJ9pYcVIUCz0OUlMCU5L+HLrd6BuVeoYlrDVCMA=
`protect END_PROTECTED
