`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tua6cCzOlybH7w1stkBfdbCYT/MDRcOQaaVZ+KBfK2hw9Fw3tvf8TYTVhuRFQw1T
1Owz36R6KQzUeVaCxLybOA+QXU7SwzK1dF8hXkDwgXn9I5zYU2N3gQ2KYzND+Ujm
VMp0Jyzsvv24pSRRRqK5/SlzJUnPC8Tx5/CWEbg5Vg3/FP9mE+q9kVxffNix9zyC
MR10DnnlCBnvD+3rZby+YlbzxVseHfJkeqvqMfGIpV+NIkZUr/c2N83PgKAqw2UV
7coIQAtt+vwaR8CoswApGNRzu0pUfPbrkul99IAkVcN7FOBMTkCDh8zqSWFVBKl1
IjLlA3llkb2RZO3LL3L/heqgNBC0AGu24IsoSLhPFtyN3BeDHtRdxwY/e34nws95
UmWeob+61eNf5M8OWwd0sOVpAunalBqE4vtSQCb3Q0sbPLBL7E321BaLbxkn8RXl
tawPspeoPt3OQYsYBrvoFnsnsHM5e/PkpqjC4bU3zLRE6+ZODQvOBq+TRS+mNxCW
XI2cgHFFTTya2m4iI79Dhg==
`protect END_PROTECTED
