`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mUMMkB5/zCKZWz8YCXCCIipjIWJsxV+7qapZdJa7E7NiezP57U6HKso4dFNJWGTW
aRpgGVjrRDKn+YyQ7ihRwgqYllcX0Q1LcJ1IylJuGrrNaFJM13AbEiPxsC+KxMvn
ALpbie9y4CYbgEy2xbdZBLU9UZPTrvtJneNWE4zvZPI+XZymZ/SIaXR297FiDdg8
XlA4JU2pWes5mWlvUHiuYAHFPycv94qT0MxpApz5QQhPWN5j7N4fuZWwh9TwrOPR
z5htwuq5P7w7l4cxrv4j6EWQ6vkzZvQTNqSMhK+R18UYy+sN8ASX9yywAAai5xHZ
xJIbsa1vuVYK3rk30GWFG8bp0T4R3L5gWt2rSrOsbDUQZvvXhxdl9qqBAINaugtp
uNrsRHY2tnv6rOLsEYJ+FWgqComAbzjaI5JCK4l9gZ79mEkafX+MG9MEjn7VDOYR
irTEjkYe7hFU685BQSin2ZYOjO+0RShC6GqH6QK+Vor/KidsZPYSJvyu074oG+jU
8brhJq6fnA8Hfi1w/Sn1QVT9isVeDzXv6SY1zklr7Oh7zASkJ5NrZ5tRs9ZRGySi
AluwLenYmzZ56je41fbnYgq3rjFXzfl7q5Nq+pBWBVgZZIhLhVvL2fPwOY77fEKH
6JidTRfxaKAPOaMjRN1ZkKmH0Ja8N+i2nA220rdKHWKWoyNQgb00R0hxJLochhkb
g0FKjdVuJk8X0yJzNxkpDuo5itxcBgrxgzaI4pIjHcum4Dx/sa60vx3ZWFvMT42J
ZfA3yGCnU+BkhM32WeBtX5A3Mmn/JisQps7dtPZWzjo+aVoX7h4mj2cd9mEzpU1O
1g8s8qTf0R/PVzqsY9LbedtWrxNRETkn5NWafo6kwuQ7zTvtWCtxwOF/dZ3kAtZ3
hiZWWuQRWvGPGkuMp32lh5dtEt+1xdYEdS7Fcsi042Cwny/Pyabyjx+FE9nK7mWN
7baiPqgZpGdFeq5eB/4yyY5Hy8gRu7VHPKZb3RQnjmNO5XRmxgayb3riqMNJxjCl
SLydr4r1Q8t1xnRIrgcESB9/sculMli5FHHWkXzMiABh/LxtFJZG+UNrSsviLTHo
9F3z9qRRLH7i7c1v7HmomKe6qk/w2zIkOTRAgZE/AQ5/uGz3i6ChceB3kJnXPmPQ
9lK7g3LP0zJaQYPN65El579jpPZiJgzUJI3kq61C/FFBrR388ijnUtPafn7dZNzJ
Fe7BVh+yD8WLw5zQNxIqxDC3Cn+d1kke9mZHsZY42XSbpUfVfCr30eBwOVaKJuPl
wfr7gsA51yASlX+yeIAU7k9QtNMgfJEzoqQXVbRdLdYjyJubJrSb39FQY6Dbfabt
e8Sas56y5HswJL/jcIYqO1534evecHa4bX3o8BpUwdfo1BQJSBsuVcFE2GEqy+OL
pmErdENZjsLVeTzKgFoj3GK2EYQl2G5SSD+FLyTXgBdf2oWBCSjhlKajB4wxl8Yh
Mz8foaiHQDO0BmOrvYJ4Tg==
`protect END_PROTECTED
