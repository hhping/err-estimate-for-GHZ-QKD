`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dR8m+A8Zu9/ehPuuTWf3Egt8En1Wpl0GabMOWgLyzD2MzX+E2O75/TPIW0MDwmKA
sSuWuUJMet1h78R41eznr+7NPIzV6Gc2KFLpyKjoDOHeif5hJ4O5YMbFg2pl06l1
2HlDnIYm+WugGr5ljdeTXvhQqrvANvgHm8zLEkDz2MJrfz49GolzafTGV6wrmNAU
Q9kx+GzflrAxta9ErmJQ+gZAf9lizhpb0fjEXrgRCG5pjh9TJLkkGDG0/RJZsafq
qpPJxMf7CEldiyHc7ETOLMCwrKFJ8mpKW18zgxXF2QW2BlafZ8dmzc3ijOPlapMr
G54Z1y7pGVMMRE7Em2YZTZ0syAeeMWrXBiA2qx7cbsXLb4471tZnSxC7ASeGLmCj
2fMYFv1IDkXfk2CFwn5A/J5Zw0s1695+yE7Ukx1U91GuU5GteWBnwCYouJz6fQ+r
3gqf7m+ptOsVaLz6ZA1W/oIINwzx9EfeVMwWmK8eEZY25oA4XCEod3O4s9iFd3az
TedYpUWRmqxublq8w5CTYBdPq2WelSgIUlu23B50JFUzN4lQfkrI/u4UZiVFsFLN
RxaUvqI215JRQkgBYCfg9o+fEYthDmfVF2V11J0S7hsX668DBpxOLJx9AmvLppg7
5QlKXLToMWqUa5acXs4GR15xaQ4j6PYHSfPshDQ+XEqnrcJBwdbnooTH8sqL8ANM
BWP9UIGV8CXUd7KA9trjbYFo8F8wPLKv/aQu+gd+9ORZSWt2XyuDy1EnHGJbHnID
3n6tz07H7ETUxWmVihZfy7G843u1NnfbRYH3wCmUhnB1NC35j1eoLSr9m6z7/EVe
B1ILhQNFUUmzapaVLASlOMKBm4B0ssGR3yN0C+ErUdAYGEszePa2FrVt1OhXWU7H
EPCoyMpTwTgVTQ1MgycVUBXd1M/zkU9whTFCTxn8aQE8+jrMEZ5uFLV6Bk2OlHFj
ah8IH5HGnA8Md5F8dJOtrFgJEp0Tb5ZOIKNvWpCw589f8wXJXSidzNIqOVgYnoud
kgTGl0zSO0BQUev7ZIMk4FbKmyKGQn6yFKESzuhuO8Wlqja8k4DxgVDKGyNoETLv
DeSyhrysfF3+oVjV1VC1EksYNElBrMqBO7iCSosT6U3IXPTH/2HdKRsWjmlmu3Nr
FND18kNg+Y4qwZ+GeJ/SZYBZBnxNlOekrFYtqViY4qwPlpxoZnvuFw83YFcUZHMN
XrLLKar3RgvfZ7II51FfwQ861/d+Dh7doGnuNjuCRMKXczslZr4cN0rQKWov0cJR
UwlwtP6m/a7Usm1vbtBLTdirduHriaa6ZXxmuhiOenezKWkL8AMf1pETTvrrKSqM
uqYyA88jbWhf7Y86ZpvLCOkxi8+a687cyxy7shR0t23pymGqdTZwrpLOC5gxm4oA
gGi0w8FazyIeRFUeykCFGKcMQRIehp3xemFoZVjF+1UPu32xvz6w6LsChJav3Tp7
TKStlE03cFxTshLdy49JIIbL6yB22C+RijJHrVZNPyNEy36oFZ81VSanJDGVbkbk
UA+mG2xBNWreEtEylAyUzdj6AtJe0NtTWLM3b7srwCGpsnC5R5aOWykjfzcDLNnC
jqj8eUEb0ewbczvxi67od/KkyCgBl8FQM7d5gJgSgFfaNF1J56soK9LckbzJHUMG
X2DoJ2NY0IKzoxQpZW57ITrIyHC14l7yK3tkOBb40rYgz2jRpEwwlpKqziSahsOz
rXb4d0nR9Digx6ESewW514a6c3UYjnA6e+5UGsfespR5tFUy3CEdJsNRfZYTvCau
4no+dCeNAM+PSmuOjNrMAz1p5EVr190FvS5D6bD7QlU1owbX80cFDUMedR81sivk
AMSmeAwmBAfbECcScIGDwOSsD/MP65wJiW5iaCp0+kxsyANQ9pRqLlz9KwyFE5eE
T65Pns5s99tnp9fznQRn8/+Dw5wLGHFKkMEETLu85JQGuraKlzn6Ti5ZckWZelDv
ayJNsRL42nz2Vs4YiZMuCskUpWO9Htq9PuFxbIi5576tL40A8hPC4JEDTQJIOI1x
w9pMReOLWpzeJfojXjzWskeaAPfbknipFnpT4/Q6dJ1DjJXamyaxjFPli+ThCA5N
SgMK54yaC2XkaDYLj9BDOp/tO9DyxcdUbtJnXE43X1Oho9FkJsR8PazlO65yfXad
xubZ+iTD85BWHrVM0GPuMyTm+lCJ0HyBJzXNaBBO6y5Vp2Mor+tZ38D7QD3bR0Ze
+PFKSFGUmyYMStP4agXxp7k7NvVe2vQYZo+M/Efi/zJvQpADdJsDPzsgPjcfDXX/
tXSztJWL8nj42BbHVATO8lT5QvtvF2J5hlywute9jTiPHb34gE/hyK6G6wK2lQhz
rN8c5U7b8pkm4NqPsYIz3523gel6sbVkCZTdbTJKfUF4+/38cHV/QrGroy4/m0KC
CxgkSj36Cjr9fvWs2v/9sRaoVJLKKptSCAQNw9ePRJWd7DzG4TexSSf+c47F06El
0DYuPoqvSAGaKxHGb/lLqNPIWjWkFstt3Lml5x1WJJi5c9ne6NDK7TqKu7HKy5Kc
P5Bufknj0gYMQevwRUb5XDzDV4WXl1USnIAsUm4dh8N9a9nY8BVTRneJNElcIvVR
/NM7UbOZgVRDwUKGMHjdsaN7320TIG5K8z9kxD4+HUmSARMqoG8rsbP59Gy+tQzM
UtkZks7oVdi2ubs7+u1/SdCELhRt+8BxsHlrR9g5pUmLg5Oc4Gdb8W+gKJadXWvQ
3cP00QgEA+/whhsbEi4cQtyh4B3nts/kH8mbpSMeuQgG257N7nCDkCBmH4dT3akP
5l71L2r7YO2pTo9cKGpqUqeQvW1NsmlKfiYPo/JQL8EQQ7PaSM91GViDRCaqrARQ
AT60D1ERRtKZT52F7fLmSyBeGY8zFz8TyEBFan2ekRwy1VjWN3YrSWBtqQmI1JHo
fQngPJAJluF2ppalcG9fjx9b5fwgNJ1ZM43ZPSD73DiDCxwUygpg8iE4T+wkBOkP
BNU2z+3YmCXt7OmhQMyVdgAWhkZyUI6FbBFfiOlvgWR46i9DuWRkmi76CiAv4Yxs
LJx7FmpTzCHNRBEcwUdtkfNPpLGCe2jqw+jhGEsLe1aJeGH88HkEfLanlaVdUjHw
2BkEwq2e7S2d++KW1mYEEcNzD4m0EdyPIF7GStZNPnynupEYDGPEako1oBcfjzYt
uxkH4C2GnSGwrDUJpDiEsqMpXNFLMFBeLarisfYnco7TBEXqRiVaNIBB4VmY+jd/
OlSxwMzc7eqXDEysiygpeZKe6eqK0XhWiZoDhLqmHIEsb47JSaayWhqMnJnoCp3L
TC04tbtxofxBHvuPjHMh/4fhdKEfAJW2TkU/Hl2pKADiJmLe9V2xo6QZvNpx35g0
eGw0liBfFBHvQjVJvq5gmOsbFyd4po/NHOzGRNBf5oGtl9gQLTydXeRMoM2vo/AB
l9LO8N5S1vCRgWs4saqkjVKHsiEWd/fhgrW47rfq9YfRUPi8T8AzAT+PgMsYds/7
YawtrcE2LXM161SI7n9gw8gqHYSS1IrEafU2yPt4gWFxATjZAvKZjYBCFnu5MOm0
0CA90aJTjBbeEZb88HKg5442Dw27kyY6CP4Cg6JStAxmKyCe0xnisijWBseqzwQ1
3MbQXkOq6IEKmOWdngkCBmGfKJPwBoyqLxAQMyIjzrwohqRu6tgitgyYP0DLWUxh
pZtUgvDAcI21HbMQ4NHg2veLFnACN+WQ9e91o5Blcmbjq6MtZnbj+8tnpwUtEPlt
TYkEkVvZdIK4szVrcjCg7fmwW8wnTdzoMjxoleqEpG0oGCuAOiS1jvJBVDn5cHRW
45RkX1hk544mAQVsAZiz0DWwQi9MWIlvxoGFFv3qKxf815IK+anA9zVBvfvL4v2y
YNsEWp29C/DbVQW2soSsvTUQ0tv+UjoyLp4fS+esLn/QKUwGcQQzrzWRgzLlREQT
WNLGxo1ChLoftQis9Z4Kgs0vQn7RKibx4FnaPBP0Yd1/gfyS/XJBGrIkoVixZCwn
h0nAE+An0S+37Y4Hl1Kq9onibY51bzkVQh+RIP73H+u+D3rEjIZzQmsTM74OsWC7
tsturGBZPuBZp3mEA9N1iRt9dyeIR1JijX7Bz0M7JDlqd7wU3V1Q399J5FbqRXPm
4ymVJDvsazI2yR+YeqxrDiZVr0QRkmsobTV2HAimsu5M6DJ4W8K8LPVQQ6UNlLRw
OV5cfLFDa3GZwZTt0NfuRM05wqJNspA/OwgvnMeqxrq/kmVCmE2sz/pnp1t+7wZh
Jqc1J1zvpvtDvQfP1uhLk56Iw23UBwjZIg/hNmZTKej3qRH5UyphuBblMLh45ema
qLJp0Bo+UiSgc88Pe7PcTr3e7GCIyB7uCnQX2oFsRLeQnVgBPClV40PVPr65jCJ7
/vW9L24Hs2oU4WwV+/XHH80knrec6TJNLSW7/fjTWO2cVpVfKwmzuuolqTdAtF2x
DhGHmNQN7tswzNu9OVC7hEorghivcMoh0fNFXrzdSR/BtxR0GPR5o/vqRfYonn9h
cfaJ4YFXSi7fWiGOFu5g7qTJL9CPyPM+rjkEUn9J8Sr6hxB7mQr22hyqCPrYKsn7
1gs5s0hWWqcHojGsc0QT3uO+BwSf1liRl6bgnb1YNipml6JOJRvYUbKhSHLdwhvl
Oor1XjCxHrzKe5PZ9p9qK/AI8homgl20bHdt+C7WmTN3CTyLTDeLUzuXQmvwyA4z
DM9g2tSqs5NZ3cyK7Z8F5zVDIIrtC4A82ZXjSuDaLrPxcGXRi7PG13z36UWcis+2
AFd6UAXKIcJHOavbgOFhJkOYMypnr1NLsqQ7NU3GJKRJ9yYo/NsVYp+YcKRkz7Co
GNuj1+KeHUoq/KgpRYRowb2IwP4206gGJs1/6thQ2TkVmOLUTdcYqhX5/mCK3TB3
zVjZVRV9bWbmD4ugBoVvV85QsyhbLO+431lph08bv5NxkvxdWS7ZFE6nAWsgj7hZ
ib/OkIgP+GP8d1AAaNzm1EWe/qvePgyF/jpLpXA8+Rz8J+sZIfwUpunBObvyySW5
jbIpnhtVAadw/CN3JpNKzv2PMgTJMaEdooh0QMKUZAd5xrg4ydulUFg32ri439QV
FZudTEz3VvT7jhJZ916GATKALb1KF3xB0kXdEDlQJjstaghVNBqTUWC/ZwCpDa6T
qkNAQpbE//N4ZicFMxAwx1r9KaAtMFKHjeL8b4QuWhFx49pRws+RRwbYgMOfD+ZR
iccue9slzS3NP5SkQ3f+gzXvX6NNQPHHrgRsKAt090ks5hQ4Jkaw/3RoXsnEWs3s
KIwwlVX3/Zn/FbpCPLqTj2upqwJdg/KVfwbu6QxvrGHv0xzw8FmVkgqJPZIFy8l6
BB+kgITCIemJWPPuF32IRBWJfBEgePQO4t8FbY0NAjc0bJnh3ot8uyl+yXwkVnon
3QgB4LHRWIR9IWpvF4P4237sk1dCJh2/soPMALm6OL1guqdJvd9f9l/BRj88UBhW
zxBGR+rXX6SgzCE9/CTrQ1duXA6PMZ8SoBCyz18ZMpVyTHmDYqyjnu14y5MrpW6/
brQLOKpBg0GSW4NqR6D8ATpc1lnG19X9yQUdns2UilV8B9/Y3cPYYu6baC+8d8R3
scaTuyJ6C1DJNc9kc8yjitoZzRxSeF7X2kRRx9V8WiEDG2ssV2L0xhJGvC7tLj38
hhQpoY6vHbGBxN3YOMvScPhLvUduGWGk2KRzbvH8NAXJGKIYmecgX5KQM4tdrr0d
lhT80N/Z1vFud1PySaf7G+sX+nQoCnTDO/uF7er4kpRb4wO4zdr+q+iL0g+aprII
LWFFbGAO69uEHqQDEfEAfNMq7lbVXmlCqv0Cs0g8buFlyu29SxUNjOnXzRtV2j3U
/cTFcB761VN5sOfhSGJKX73NIqcoCSSOOWp6eweavovqJpB7KurXckYqsM1WJBqg
aovq9AVylTjPIs4voZx07Qu/LpV/FJTWt7WRleVZgPzmQtoiMec3QA+Q/hRrrFfe
nBkHoh9Pqx3ngabVpppmIrkUK8eeHkrZwftNdaLGDlaS8sIHM/gyI2gZckOuQnKn
ICR8chXN5tbzHjdC+4xRsXcOnRet/glHuLlwR+k+YVOHiCgzzX0MhO52rQXz7ZVw
/buj0fqw3R/Wy9K7f6KMV0zj4FBb6PUaZQlWSAHhIWq3dH9YNckRNYbqQVkTU6k5
vVeVZoJTjUeN3Lpt3YDfMBGcRG8/xOoJ1HLfyMggwRUfGfOS//iDql+YY7+GNoxa
p4Kslv0lQSVIHSbK1IFYwWft9hQ5iAKhCTylFJXiiivT1wTu+vYBRJVZFtnLsUsK
Jbi03xuHixx/f5OquFN9aKmImg7NGVJMonxREGOqVP3QUkPiayzJCvCURm3L1Oxv
vBP/zxSFF3t5TSB00BRVFupomugVbFrxHVbboW+gsSGVO8xi4tVKh3GE+VSOMv26
zgkI/WHeq8S/wG1WT3gCzST0KjkZOhXhG4GIAY7Qki7A+d8tcy1H2hW9o674bbth
6xDpJyErRlKvgZdsHKHCneF72RnIA6Oh2gx7FRvWajGkYlh/RDobTIbXz9zxzUdP
tdaLSFYIH4MndtqYZQ7ZCb4uYY0cZ/LWO75njVue0zBBdJ9D39MFAjEdxqupuKCs
dXzo9j/ertaicTca4/nbaivZX5ihfHzsNm9jSfYSNO4T0ZsvOnYCccAJTkZNjpRj
e+jgby521brGGXTdBfRAfVEZB0bFKgG1T1v3C2oOlH1ymX4i6YgyeWaenBwmuFF7
JuBrMRqKY7zu8LNImwt2zWsNkqftC99e63W7B5edvp5787tWn98Zp/eeKkOJX2Tr
8dbodEvhjs5N9ufrcrmfHDOvb9Hoy3FRCLlhTUO+IVdHJa2Iam/e2+XJVd0FyNH9
+RTUIqJ/Z37tflh+jkqDaakAU5rEtlTfeTKHLzkN2BO/OoZ41I6Ys+HFmcmdwQt6
duvp2nbDsp78wXAcPRrgWur2bjXouXpe9PZv8ZTM/1n/mTnBJRyUQxO6QOvueOF1
/XORnV63ThdqRvgTXw6VTtv1Q/L18NXKci5ZSUIFOWj4oMJ7fgrsj27kP18W5xWV
o/x5pjBUd7RDfq8dsjwSbYWUVl34EaKMcL6Pz5/qruhxedZj9bmXDnibxQl0w/BG
8U5gPCV3ZQolN1qpCxlcw9NtC7BxqilH76COp9wVfYGqqof1w6jzTH5UFmLuQk5i
r/mcrG5qeeI/82Mmmz997ZzSD+TByh69Jy3QFpscEfDenVc0G7Ub+zylq+A1oXfG
INZXfoogmf04B0PurmA+U0XPql0C7sMjBzHdFkOIAcnkGtqscIOR+XYWdx7PnqSb
Rrk1Nzsg+00roXFkPNTYpn1OBXvoRCqyJ4rnvAvn/T7OqyYKgndnEL5fGqIqw8FA
U+wcRH1II6/kaUR+6uSZA8aeLIBSmRw2AfmDGiXMCtXMDGf2eJm8slhZAA2riDxL
9dBBpWM6TD675px/fhCvXx/YNjNfAVzUF6/7Fo2fSjS0w2/Am3nDSFUuVMYKfS4B
l02ldq4bM46rajAa0KayQm2P6aOjWf3svTV9rq+S7Gc=
`protect END_PROTECTED
