`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ben/9vH/kXvxzM+PVrtvPzdReVMvjjjXgc8jiPO7zIZT0GJmo1RuRR7BDfID9iLv
fBvrHpuAaLr5QY/QQeW/Uc6ha7NOEn1UXIkZlKfvZ4WR4wpPBtO8Afeb9JaEtsVI
cxIH4n5VcCUyBo/8Vnmk2s8q8SSXp/8Tfd41V/EAJLDhDOZqGFRzWC2GU3iWxI6l
jt8LLGojvnrZpxSLzgFOxZH6LktuKGOAeG0r3RWFeB15Pfwqt7oFObvsPQ5kB6Dh
3FOb8s091cjJNZ/4LKh+lY5+QZVEliWeGqMWcoDsdsv0+hAFjLhcDm5Z4DXiNkgu
/z0wGGK6OsvV6algr7Mn5kvULnK+nRGU3fv8/x87fnkvYsH1BQxB/D07urIhAdzg
nwrQemaSpJPXM9RE4UE7Z4gJDmmzuuWLoa7Lv/iBCl4avLjzZAWGl+M0cqOfHnf1
VhEeO+j6mgqLCI7NBREMRVmStkvg3W/BdbBlz7r8QrIbD0G3Velm+REQaWATcqU5
8S0oOBnCq/NAKe5vWz3g9px56bvMjU/dh8r98HebvpbEbAkxBlUYtrSlmYMxOkxN
Yp9HFTBPuL4NEwIFf245O3NkvJIonQ3zwquq8urG3/IBl9TUEw5L+KFixP9B90/J
ob5x5kB8VKZS4gxpmLi8fQ5Z4zvehr+aM1MPVYPGTw/81pyUdVeua6qNfAPozCej
iPUzPSVTHUgRTaiLTfXphACwFnALfNGxGK8iF6O+yrvyKiuyg0YGhSi1lMcWEhvT
F3A0XpiMfgdfJBZ+AAilZ8YWIBGToOddYmiOijSlu+3E5EU4q95pECj41RoFcJ9q
`protect END_PROTECTED
