`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4IGPU3IVuw3paJsBotuqysPRYqog1YF6MfHu55du4RSJTGRZXk8Abi33N6rM+TZq
y6DsuTKS+5ye6nUkYw/XtGazqO3Qkq/mqcdBzeru16pAj52WpcadwYoNsUtDNF0D
ScNM9uzr3zVQAJ3Sd1q5ZwNxHtqMYCtLlMQHuTrBNb/CeVHCk0Wezabq4J8TyVVK
1Ihm7F6YIEPhJXVJp/Z8c/TpmPjium8ksiM177ouws1OBgM8lxauErv/4xytkiPQ
JBTdna/2pb57PyYVvVVHMTcfrh/DkCpUwolS3bdxBq5TNNf6qKSkrD7C8lfHdA07
8A3XxhRE642WpVfKj6X43U7YTh0oozleHW4F5JOGXUuqbllvRjcQ73VYl3XWvh86
Mz4My6SYSz7ld/akZh6hZqZGVaqBEVcHL9RbjTSF/18Vz8iSosJns6lvlyWYqdYV
gQxLp3v+HpvqfhMKNA9AzFZZnpawCwDJKiyWSjCx2iRKp97GI3pIXvzEngtQ59MN
QrwNfK43vOdLffJcvSQgkCV9rv8M2o95Dkv8NW5GRPXFQFbjcdNCc7YhH6apuCxz
6GWhDsU4GbW4BshvLYY2mb8fvZ/9I0jVuZZ16OsbuapCEFhHOhENtY1JZWRO799X
CzsTZgMnYnsja1ciMpmNXNd5baCfa/IZVqJbDf5J6j+Cl3RsJJ4LMEmcQ55deHWb
dN/925H3zwVJucJG5XYVAetXPgncCasIChMXhm6c71f0ypNARzt+uUHhXHZL3+Lm
mTG8M5xF0rkffGV7P1gzrTLhSbUOGnkNN4RcBmQ9NHk=
`protect END_PROTECTED
