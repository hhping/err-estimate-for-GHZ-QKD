`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SOiDD8NtvDN04EU2yUynQ/72bCRYlhulh3zE/SO4oppnjE5GIajYDrXb5DWa2B7I
OSbUPRJfThKM+VGtLYy122qHi8MB8/hNA/TLclK7TCwO5wIav/+fdVfptMnU6KJx
4KOgNLK2aJTyoUNfO3UP7lzVj2AwGF1TMKR1oXQomU2UZHXufagNNNV7e+edJfJv
0eAvO8jY+FtylG8tSxNRxB+RB/FkuOGG+ev/nxW5vuCpKo1ySnuPC0dNoYE6/cJs
cjmbXU/1YefPFOI6Nz93iGc7i0FwScQONMuGeTQweg/barvILlueRak/JUYQVf9j
D+4bl/Xde5l9ZbxsTLyomZGBW6nGdQfvkRH+2rifFws3/Uh0sTJxalOktw5LVxg5
3Icxv/DOwHKvkbjkJh/A1vOFNecvXecyDjqSJFGREawrULSAdz04NZFvSeXy4Kt4
cayHIihiXhgkkXkeMk3FSUBF1WsxsxYYz+ux3CKqRrkBHk238LYeHkTYOGGM4ru5
f8Ojhm/yhH9OJPHnmOQBB9bzlGkaUkZ6XS8w5REdevcbuC1eM/nFaU9CAH361qF+
hQ3p2LbEHGf+reoYXfd6kxuI0MW9VXsjYr752g5YfwhvQStTaY8KjiAmg4vNpWWm
qO7BwvbEPfv61PZZGFviBa2AkV0bCtdqkiFgMgqpLPViFckz/fNyPCvD8kRKu8No
KQxhyIV+EGBZtTXpRXPZsTTXgEvbDFE6CZEp+77beTJRM8dTiKxPhR3hdMSagj6U
HkKoWpQZWID6E9AE+0Ge4rQnb75nJVePmk747QA+GgWjJ0069OdImYjpKn1AipTL
ZG9ALHgJ3dv2zHKLBypkpO5BXgV4216VRPog6bqqTuxuPe3OcYPM5YXOcYT6kGdL
z4RQX4/po0PvP9a8qIJyavC9IFLQ+d65kEd68g+N5xJJbjGYnU6tAmMbEKKnRuEZ
6HPPH0ZLbpBVqWM83EpeCU1mdNdSymSHoE2UXv2+r1WmojMZaKg41pSiDcr+k2s/
ZtUyQfsCV0VN3rgzOFSgfdDQVeI0IOAQ5xusi7FYqhCQCzVL1hB3lRACyyWJA8NT
6HCzBLH4tpeMQJmCWWCmPl87fopo7j5vkXEj21hAe6hj2qq2JxbbSEv3ZBlTFEbj
SCZTW6On6TY8uiK8sAAPN7oO+ktjvHJxVL6TAXd2j3WTMKEypNSoB9QOAAgxolga
a+nWcHSJUMxon5Js5xyn7cQFeWYyQyXHGQFgnWyVboiXQEydniLSCfTeF5OgNXvt
wIWChOCqbHY9KVXkjtGaj3ScA20S8485APP6tKn6zEOlcg9VtoKNE6Uss3JNFlci
hp9+2x/Wd3dG/2DUWpLmPUch4g7RLKimw07NJ9USZDP86z5fTcnYVMMwJ2I7nPp/
B4znhmSv+depKcTNREUPLCdw29uApWQSK/LOi5uGxvRicQQByXprRdIG4PDL3LV1
7waBOZKOrA8+zVE2mlqNKz1qKiZC1CuaJUstPv+ZwYx1KISvIfECeB099tjnPL+M
lYTncBMTvCB/IDzSZryPXVjQKzkuwcgsnOoyzEwpmBEdpPc+Ll37IU6LBhKOIzbq
jA90ScpXH4Rqn9nzfTXbmAfMbVyA+uHL6upLJhPF4RvWJ5Zm3oYVyECawyxsSOxw
rTwoXdqqH4b3qWvEhYpKs9kKRf0zc+khzoMWuXuWjE6RnXvYjpX5bZjRIOwXJnX9
/9e6FfTIGCJQje/FJxIt3d0jAEOGoX6bGSj/G2zxvBdxhU4BdHk7vvxq09U9znMh
kypseFyNiEG18CLWdnHzjQtRK94uf/RLsQ4OFVC6xjptEJ+yKZ3utcQxZ+F8knuL
djdZLwmkeEzI3minZc4SnH6ly+Rbpmz8HmJIcS9AuKqrTROJw5SQDiUrN9idGxlD
SmjihkxQ/6685rnsy/uF/cEmVHA5hcTTbjGSCqfO+EG3DYKfZbtzmdVUCbBsX7Cm
8UOS30sbwr1o/2gZogOeusgrzPZOoSqEekVQQqjFrgdx9ukp7zWjqo8lVq2mBTn+
u/cEWCXKEpjUJMANPLbujH0ACy9eDfnDSNAlIWmRCXFtA6F3aO2q1JKLBif/cET8
CTFKltasP098wGEueJGcu0UJh+pGtvy5EKR19tFlF11x7zvgM6Ug5TIoU9qUWPd/
VuR8goH6rmBJ5OSw+tR+VJ7OUN9SKlp63H0DYMMR8I0/jKk7Ub4SG7C4qgE1mNZN
VEODVmTSSZYA9VFDsZQ1i5CKwdLHXOri/gnol8K2NxX3oyJ9OxrFxfjO8xItAgp4
GH7xhmJZrYarwMfMr+vE2zLNWtCRhHnHQwYwvx+G5JZOeLFjBUo/j0x5Qdem0pO7
UyKrx2rwDapSeKtgMinRe1MSl+N8nAlwuX3naxJ1aMimMVknFjkRYipp2MWsnzxD
q+KJaFPtHNDNgPPCdE4/niN6VthbcHOiWhsIZ6Erzwg3RCugaUGWWZBkQNk+Oq/v
2Ww9b7pyZ5UhFmcVdZWsJ2DUeOchKZl0xhRw3wmApci1XB2daFs9LxBzmLH5EAUk
xg0p+HJNR6b7MrxGeJFBPgJgyB3TxAlYGzHuhdrA4x43XcEErX0hYO503BZWrGlJ
asSbp3Ni/cpRjxrsd91Ip4K5aNbaE+USYFDZhoTJWo/tn2rhvKNLdBIS1SC+mLeQ
totUAUtl234IsmHNlw8GfQ2bJ+9gyfqYcWmrjSnk04UVsl1QW4L/urS7Jlg25NlQ
vXqc9aMdaLTLgRQ6pJqg2ijUpaPlUEh3nTPA6oc9N9BugLBps40nT0+4+IkMnrWq
kQMHxHBOjqzOPaiwjuOANmCEitvKTeToYNtwPWIZBpnag5HdjHrC9cIyrn8cRi5z
1TQPajBGuTVEBsfHyHe3o0k3OH38bIrnbr6td5jjHXIGiIt3vdm0D8lIzb9kCUPt
p8Vt+l+9iCWm/abJVWVcOmPxSPBxPgj5ltu81EGsGahD3aSM+vWMt+B+ZppP2pS8
CPKWKwbLMfYMGtu00/AJn4u4XS2TgCWlbuXZpunIk2wNLH7GWr4wFNdX9UpkHtTR
OOylwtLaiua7bvmGRSBdMZ7u6c50HemiDCNG016go81CbZ1c5VBgMA19YdDtRkIS
RsU7HxZ362/FjRYflhi6vgRj72d4tRi1KF1SIssHbXJZtWtmc3brMkzj8ilP/9n0
jE0AeI9JmSdGPd3JjrsnfDyrBMydamOfT0WPiAF6Crwoc0F9xFGkr4ootXA9NyOc
cTJebT7M4c81ZEOIyG6WJqRkpGrw03X+TKjZ51SPOMpFT8jB1uzKvT/YXmXwskEP
5Ees6Sy1J7nMR0V6QuxT2wKB4mn6tqGm6nK+ft9RsoBlO+TON+eZuYtKQT9+PLBf
nfEYdnBSGoxf53RR0RGIhhh1gDFEs4bxZh5ZGvrZD3pVJOCYqX/7P0UF1QR7NrgZ
877QsWpYCbRCa7LsNn1fAuuecMXMqg7ZhgTWMr12P4kV8mRg/0kqNnKPTDRpdA4W
paeB0KLMyWngVMKeWua76gWSmKLLuv296jM+DaVpk4CIkW/h5HSrH8BYWKtMp0kg
lPzoL+Ysttn9rJnhCexcqbel4OYnLsiUBm/davTZytEM1bWVYjfG5oisAu0txm4K
whP4vGXsQim2yC/NIJLh2TzdnWr79nom5cMWdetwqs20U/+q4fBH5vT0HUkzJTzf
5ZG79rXIvmjbMfTOPlVxhLnLbLEiTpsaWa64pAQrKwDiQxWNF9ldeLni2f65yknK
mGSY7cqCpVWs/vTXWtIRTy+wdYblDjht+KR0PXzcL0HD0yVXtGkuvF/mCfbyiJPo
0rRPb9rS7nkYETQzLxwlh/edk8puQM0R630KefvpaSLfDfNR/c6DyyPOzTz9j3Ew
jY9ECQYKajQEA/lpDmVARGjOnau1RLdHCtYFysy39rJr+2hz1168VYwzixWauGVa
wpcjhPf7oHQVRp0658Mo89L1zmVvh/AzBQB+sf9NqHwhRuoHHgqbwEvWi35b+y4f
n+z/NSxAe2ddw9d52nR84ZqxaYKJruefUN61Ra/ZkKmQAjqfRnI3IMBd5wfy7kj5
xs6bLTVvobH+wb2VcB8zZQ7XLJA4pjO6YbkPvbilcmGT5VCdTbHiyKx0BpXjMyij
fc5jtX6LPN2m1/j+5NHdIrZRrESIz9faoCZuIw89AMearlymbiERKAq8U93n2Svy
RUVy8lh9DLkQUYWc32GDetKmbMfUBgSz29Og/xcHjjs85s3Sv+AXu2ALL+nLFBli
CJSyVqsLif0kBtBMnKT4XGEtdSyCobiV0ORfJkCt8+wB429jNUkeiOBZkVbzL1GT
9nFOSBswATYQLJiDsYMIbMVttsdQ+VXE+7jZAJ5XeOyKa0vhikMb3yXQY05KpTeN
NmVsleDdEocjpGnjd3tiqIKFx/nNLs8GgkkMeWEeLIkEDfrtXWc5UGYkF/JOPtu2
z7NKEmvUsZzS0reBlIbeQbhcaEbtoAiNnX1BFoJlIOSrFhT3ZJpaIrGdUN1MIPCs
lSyJDLeHpmx1AHlhcVaO67YpN0vdJyk2RBuUaIRAAgnHfLPA2d9ymbKr0Cmsv3gV
vLTxFgYfVaATKwfBhD91tSS40o4PF8Zg/85Rfk8AE427w2mvA2V/ZjIdR1fGqbtL
Bno9pl8pBiCLbLTKXtw8GUo3lx8n8KkEcxQzIpA8HWLfgOUtx2buihIgDpCp3jkm
/LPpFOqbmosMvDZXQGYCgIVS+DxBsn/29AmyvJlEl0Zdt2PcMM2o49jEgioj2dtJ
RUwWD559gnnHPGyKUT0yIRpinjC5q8d+Egt1Dg1RrfzOzwkIJBRy+YRZZISQI9r3
UTxFTDbOurTYJoJMunk0WuwZ/ZkAPi+DhqE1HkFBArEw3RqGewXsteGjYwXUtfT7
1BsJehhmIHxpvpWiED7Qv2nxcZoB2Bd75rZ0niR5lbxIUnLHIXVyNEUleYUwLWDX
SacvsZH11c4Xt7nOvFDUB9BNrOtQC41jQC8ymEcWtZInKffM1kB31msyhDySlVp5
K/GTeMBtOCHrcgNDlo3cvlEBj1ykYzDozHBnGcwjBh+ftdUILEunYNNYg/Pgw3ss
0tIN397lKF7RHcldXTX+JCj2tB2OO8uGWGrGs6pRXrpirgvIIywhjs65XHbhz621
XCI9aX69qmsxq7Y7IpZdAX9IiLaXClU5Gi6SRRU2mR2TtydtSfhvig77vulJsdLj
9MZn345JeLCZx9IFcpmPIuaP0EdAbVz917pNrHYtLeqMf3iBFzUFka/BSUxVfqKi
A9mBwHQbg8O0uO7crq64KvNwVH7nsuqsbzWT9yu3lcIcROuTdZVZoGYfDyTbIFUk
5EZQWKEJUL6iFkDnq1f8PAUnKYL68XE4XIqZtRxeBS9C1cSmKxvVCHnj2z6SjAtp
nqGRM8HrYrmIcKI1rdbLKMlDiqZNgPnSrvSUc6+rrOIAuB7eZngbqws78xbIGjz2
oETWbcp9JzU9FhSrKzYdg4cdRe7NsdR8+/zfGaKG7nhyvliKqNDID9YTtRGR0kZ7
ls0+eytnhaYy4lr2MFUJ+x/Or10qqU+y9gJjcy3iI1Illes6xWbVyict/YhaL0xz
0Ya7tl6llLlOv1YUjRkvyzbx0uNxCm8eqxyeyu5ByHqik66bVtIuDUFBsaR3nJfA
hsjSuT1z4a6LUGI25QvCnVGv+MawC6ybzw0dPbcn2JPAwvjw8unTZvSlciKqqrlC
dihlKnHRiYLkmJN1+eE3SDIv+VK15d2CkHaUDw8Tc7GN5CevvYZAyYysoWCMdjQe
wV3iSSM32DCj8y23Hk8eq0u/zOzdzdEryxWEd6hhQg1vIfGiZjLfC1wTtABD/svY
KLZmC99Gl8X0kJ6MfIXqx38OLpDWQwmO0ScbCQm4olaCKo9ww8jJbpG5xVXpwH8X
e7UJiKgkveT3jyehYe7Psqf3RfsW75XOz1W/shzNWXLFt8ImBe/RSEQalh1nd2EY
RvYiew8WgJ0g7gOFoEXvmmTk0rmlJcOzoGN5PA4l32tvtJaQpCy0cLE8CwB2gxNT
anFmkvThiaKwsZsUGSjDVHuqfjE9mEBBEReyptQa9tA5c0mhhhbR/YaDpjtqeD9s
LVJYRvN6mANIoG/77pUMvo6COyYUwXcvzd/w+YwsLWBfnBwOz4z1YC186aFn1+d4
liu3HV9uUe8I+UeX+HtlzRITYMsttds0dvYfvtOTuVWECNJoYJq21mydAaY55UQx
9xDaAxGthlGWa6XioIbsVfnGBD/5CWDD8BjPalOy/c1nihGHn5xPq6yei5SY0JwY
Srp3/kkj9278QQegIiyTgQrTrUCKc+VLGTQKGuXlNVm0ymSALh3vqsDZcZ3KJ7vn
Ddx0pZBP/Z1qlzZQoR6l/fMMxLRr5RGbUkyAtVtEuxJ5SXSEYSusUD+6Q9GhLY2F
IF4cIf2v5gNrpsb43FFrYimvybuoDyC0Nxud1JbccixKbiRgfLVvHCJRrNMRa5W2
L6M6VSsGP7DzQgWtaGRSMmlS7mWm2cA3dUYwAQatYGMhlAhJFipS4ISCffrW92iA
MM21crUqsDOpMVCHJ1sCKEhj96Zk24+akG5hMYw3bAr2uXsQYUu1t1D5a6VmoXxj
dHoeOqaZoaKOLCvSYql/6M8uuZbcOz2XOBXMydFcYGpnCVGW+xYBb44xG7XZMihX
bhhpS9iPtzeBcqB/szgO9rJdbABn6bbsti/IxeBjFMmli2GXQ2RUbcuc+i61/vSA
uNKhnm/IDGtPO1uYJRhJeg4Z2ZN2xzTZMuSwKYPeBTDNULHDclhrdyCuhoO6lzbn
w2dy4DA6fx9ch0vD0kWurqQQ+I1qPuYzv4ks8k7dN2DYE7Lbo2y8vFBPyjhK3qYy
ba5pa0ue3TP9qOUNmRIAYLhRRk6iw7A8G8m7cL6LYSK9nFBTwI847hFmOVr6FiIH
p3EkdKBo4J/glxhA2eW0qWW2zy12Q+3Q/zBqO9YcNVx/wImgzcEgLkI5/C4oHtA/
/K7fFLQOHqh79nVzj7u+LIg4vrHT2caSnvhkHrNpsCLuPPbWyDle46KVPOLLmXHs
cyap5x5TB8CZ9tWU5R7rFQTz/mSjXSOHMYL5D4gghxMgicdHJE3v8TAdRFZutk2j
vSvO9PF7elwMuJbs8vWQ5pi/IpTxF4CtuHw4/shHwHu8vYqeaceWT7IrmFWeMdE0
zdkYOTJMv4BHzzDJmq1HYZthmKsR6ejHMUyQm3ASWZ7wwmg6f0SJ3yFXn6QZB/UY
U0jnJ2dhxL2IQtKGL5HfJsU7U6L4x47Vc05RxX/L5+7IcOXPVFMrQQfJcDvoZBk/
neqRaW0l6p2PwPNeDnmmglLP+Ag1Efz3sM/lB4fmCt3zGCrdsy881vM8IPeefh+k
2m/RPM3v+RF0LySbsIAo4bcVXC+0hWOZAIgzWp0MMJu/DUAYr7cRB0IJwD4A1ACG
7LXN5MwsFCNfLTr0jZPAj5lvw1AKT5GnpsJQ7euWrXkIEgP/GBhXYPJ4Icz0lNRU
x6NyBdvlkG+Jbw6/cvhtiStZJVwE+oHnsrKnZyPbdJsYMqR1/NYXI+0HID+J8K+Y
5lOCeejAzA2kd8zW0VG5CeIgmFFxH5r1fs7VJGXGLSzw7IlSj2QbHcYuLNbuyBs1
c0TGK1fDZSkB/zR7KzEsRMCqab86BftKCgeOUIhKSeSFD4Z+0cOcBzL8B9WGgzQo
wLLmwOgZA2giOvonKihHtKjqA3m6ZBz5XVzpwAWKAjLufZ72wPqLhlMHw6WZL6hQ
FuCS1cCLygd7s2yPY8IlJGQQfwnvenpCY/PZ3oEdzh3/8MH05rCuR9P35HV+OInS
nsGE45zlVK00SoWduYQzHijpBxmaMYtgv899R2GOm26XTmg0wx7YqDtIC9eD0TrU
0URe5s/AnnrGVsi7mIMcy+FOhw0FcefNQVecVnRlZ0zkQsCRgYhNAz8f6FiVz+eZ
XRnrHX4+WiLf3eQ8Q0ZYuSuJr4u35KMg4M8Zb3WRed6pBgntVM2NsKRWqcxE4VGw
ZG7SJeiGMlwB++jFlxaI1KSJVK2Fc0gquziawdJbZ0LzLDooXn1t/9oCXXa9q9p4
pVqYqolvIdPuTQArbMKW6Ep7g2ojrJ9eAE2FQkQuqRtNwimM2LY7iRrnK0vDQTLC
uVoA/yagN9jMWMY19XtJIL4K8rKFr8x70TmpVc+pQQHY2WYkHT40kB1NaKrJIdzg
A9kfa2ob8hfIan1CwQy6aCFrIiISkDYpmTHflMfuEtaVPANkmmxILJUN2vwspMlW
uwnszYKN6OjigwU/HLKb1bUIsAl5LjI2rgOhKo56gu4pZIZcqhrasjd4rnWKNY7E
M/ms37FxFrF5Pft2m44fO/IUNbDrVbyaD8Bf9wbDK/dM9Fx1AdqX13XQhzWpnxGy
QDiHh703ouUmUGyNLM+fkvtCyFLsj/semG8j3Vtt8O4HFzkt8kwt2ls4iUHoLH6L
Vj+bf1pCfbwK4JwYKOIdjIWGzl6emfo+ldOEdXqeHdWtYmUDnDSdxdtH5ARsayve
FfdmWor7uSvmE25Qck7gcrhwiPeKdjxffIacQV9UvhiMMox+Vh7vduYJbeQd607I
Z+CJMQX3pab9rnPHfYOtQsxQ4bgNyYlaOI/h19mIv+mt8+54iQAdu+JpTwywu8Ok
dvn5vOjqUs+zP4/H+D9ysKE1XzppuOaxfpqOOkTyF2sjslR+/MVIKNWs2f7oGDX5
dmySXP87Vt9Qfa4HLq7iSAmZLKJsADEaJAr/ugJ2hHzqZ+xmS1aveGNnNYB/CgX6
9Q4UXvvc7xJg69bkXy4VRQ==
`protect END_PROTECTED
