`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zBKIpjMRDaNeD0IZm8UhphuIsEBNK8XCwIyKErMc5SsedUQ0Esh/HWdZ1h4uZhpj
ZwQyUvxffZVb9EU33RW6E8biplcQdkON8nSJAiMvoRZyhZFuxkbEieTJKKTqsbKb
ZDdklXm8fZVDQjVHcruuDIztlwBWdhOoK3DkwtButq+YOGNCffVBBziT8+rAkiDN
R4Bn/epKH4fMtZqAmiC0VHbX6A2x773o4ORNhVU7EmjDpnScCJDNCM09k0XiOFpP
Afu7TnFYhOrEWFdr8I/r8Mhy/+dpbULj2aEjw3TrbmvMhdruwpDI3q5QgpnW1Y8g
+RFEcC34bDCFNTjbD2O3c8F743eFd5tX8Z5FXsBwcM0nvoB45exNJps6V8tfl8OJ
IH39IbfQax6Pgt8+9cF5OMczhAb5fSS8EY3NtwpYFrmw0QvDvHWxRIxHqj/CNUZi
yoT8PJMvLPQrS07I66wXoZMgUo2ZZaHccpVR6REnfgNoyfyYSPuyN2UsmkWu3nJN
vnS7GyW32dzZP6ilFarZDZzsQwq4ulj3+hTCFBiwu9tBKEF3XmOcqkpt4VzPqY8R
Ab+cx8YvfCp0Xsy37f9BF0Wt+Hj4tC5R90Y7WE70NsDm8byE9nNDZpwap/HvPX4p
L//nv+e4CZNB/IMm7y55t8y/LFFqA+4G03yieMVkuytY2qs2S5cVf7QYRqGmHVgb
WqaMp2kMPlg6V+WsA5BISuH3T691ihtEtqMJndFFS8EwieEja5/pdJnh7sVTiwIx
VHVNzj7BMF4aC2p5b3NddfjWCnC6qgJawO6RBx78GkL8hXpkrpQohXJKNeptymYe
TB4sBMTWOPiNzFIrRppcWFKAsnSs5lZjzAYL5p8HSrdbJy/UOC6ea7bzYhKmqQol
jkXsy1s3IVuXV+JPKqc4+g05uUEyvILkGg3iwlJZU78hvjTi5O32UyIxyH3vSMzP
5EdhYyR47bnfRWGQGbgmsTcUz+UuMsIqWy0eghjGxnrlRkXLa2XVI2NnykIyKmHH
e4E2GWftq2RJe7mVLdRQywxt4DwpqLEQOvC0ySXef3DhhtYVw7h+LfX7UBCjukZP
Qbg50+okpy8XpkUX6zNknbOxUCFJJ5SLAdWS7KYAbqMzOXLbB4wdz34yFv6cagwi
EDv3y37I90rGiYU+CSpTieStSnJwXAd5UtwLN/gcAzcRvzA1+u26joHztTJBzGnb
RUlYR4CvtzjcHi8T2rISo+vX97uBdDlLIJ4DLsa/XVq0mbyRLX0hY+jleNUEaSv2
iGqlPxs1iyFIBFhCrmj4MC+tonLqUfeBKjyMwCpcBNlMwUYMXGOuHTN8HfgwYGt+
aqoiI1ZmVm9Bt6FYHVmUBh2OZZL4lS0oio+4p0vBw1jabcQYSC3lkhLX3US320+r
gWMPBuwAOM6jWfDw1ezRZSLWbfQSWYgbZBNiFubCNxBQ1rT90J2/ygMshiEGhe0Z
fwq6aMTK1XF1TLrA/wHjQPNj3cYpMWEo1TOiVZAE8QLZ3dc9thsbwBUusZpP5eOI
/iyr0x8ti1L5N0fP3QV25EK3NlPcwJAvICUsWiHfgJrNwlOraBGtHr6dSKutyQOf
mkx/dpJDWbc+BkQzCNf12HrPfHtL7OBAsmdkSiyh3Mx++4lgNeD7PlIKi6nwQsmb
TacHbWYa0aRPQ7CZrZYYxk7/jln3z9JCYuEvJG4kY4+3K48ewGuipcCrlRTlYX4M
1vRebf+Yx9OXrjxRJN+jA9ilvoaoAul9xJhz99ejijGHWMqZqXpawQ0qDhxNKNoU
7mRAggKwYqlqFJjjT0s2pEOhHUg7EPKgyCgh7jO2C7hZTa+Bk//JOLgSndDLeDU9
lagegCrAJYSF9f+BjRHRhUjia7kB69mR7+GxhWL0+kwlzq0DXWgch/XoBwARh7Ic
FiEB9s5BfsnGNuN11RkMVgDaTO6i0chjTqYxI6OydkWP1+3r4DLEmQUlHAtJOrCR
7lCQ4fmzz3D+qJDfADu1gv7cQ+b8ArY2vyiIRkPdHY2/R8dT3QkVbMlcKXOa8AfW
kA1YhJWDYwYZV+7kJxOz2JrPnoIGGdmomQQVeH3RdTFOYwTwMj8ugtrpA/1eb854
`protect END_PROTECTED
