`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fYrkxGP1bhB4wkClPKF0lcBw70msykD1+STViPObZWEl4g17rSQJrzYCx0mKkak4
3+vm8EktsPbZdtAYJq5I3Ll8KtWK3LveQ/VJ0G6bgIOOjDbFbAofYP2yydWhESsI
2b8w93K4BmkXiylvl5s547A5XiTve3dcjmcb7hbY+cknoUR9aqmUMbFA54HPp+9B
Ezbc33TO5GrXz2tit9DbJ+CIuglJwxzoxlTKxEACTMZoa9mvctKRof+ffJ1kEJzq
aea/ooIv3vkA4bcibn71sJpAyxsAJrzhSyfy9wIP2x8=
`protect END_PROTECTED
