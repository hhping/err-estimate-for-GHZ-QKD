`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SMVWzjcNJZqYIeQDpfGAMfwkVkLZz2KLkDqgXuXPjZjyKaEeHQcE2qstjPCE+Zpl
/+qGOAPc/3X3M6N6wB2tEy963cGxKgldQ8ye4c6/5e3eZ2zYjIUB95BIpinAg3UH
6Gchd/zMVqQAEU2WBxDfNyExedTEEUX2zHij7/VF/n88qQix4F4cT6AHzmOxNE+M
XWx3EhcvcB7ISf74N5QAhMZID4ROkDiVvft5ZTUKNCIaVu28LKTZoaHZvOKTm9ZB
YeK/ALyYM6tkz3vCG3FuTuFUC7PgUpbgUNvUGGxMyVQ9LX9qRBIEJaAp2UojaW65
ryeL2EuJ0dBRHuzW5Idqjq4WD7HHcP1ppp/Mik/Vm+24Ptq4oMSlVyDA2zG6Ar4J
IDBbWoqxFcPhqSP+N25X9k9EzT3Nb6BRYNSvHCkpFXj3lPc57zMJQR0y9RiCxLJr
07FsQ32Imhr8dgaJrRD0wY730cUCGJmlgtvUGFMx/43n9xPObfk86doW4sQe+K83
gzd/pnxzKo76B5iIpoKCvqr1Xw4PpPvMTNIz5zG4Soy7dwik1W1LY04+WXf1+BCN
Q5dKXp4em7jwgHlSEpwNT0HXrZI6Pq0YH1aA9w8qb5a6KxCY3USdkMePkeaeplYl
ZmM/npE0mIC6492jbWTROlu6euiXI/hIhSFYOGXyX8uQ9sm+W0S6LFHnKLs5+uPo
FeF5b7QGKF6RVKIiUHyq3BHOk4peRg4h9cQ6YxAC39iiWD54OWaKed4bMyqTfYu/
`protect END_PROTECTED
