`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oc9aFsLETcI9Lhcx6gp3QIHHQvJOCCfKdAe8iZycBcGzgebleDYj0HdSjQ87RkD0
cDNbWNXKlpcmIynHSQubsh2uYCfoLeBfh6IGeKJY+GyevwrSwMBP1ApoRwtdTpZ+
OyyzZ7wgCazzy8HWks5PrLTh5ZnigBAa2cEjMa0ODeKZrskNbwU3UKPLvG1oRUJO
sYOW/X6XF7wUmjeU2xlLVm9TzmLByNf6EnqQBZBehjsRdiP8uaGbAwI9NrndJurT
C/0CZifk174a85yp1yOskg2bupS+rnL7nFvr3U023LN3xcqi39F4kXScik1mZSpP
08kbKoSBS5hJOVaCMND9K9naKSjNBS0E8xxH/iWhKdbukqsN7NHahWU0ChO4zdLU
fVBsCSHt03gRnG50BlOgjj1rI8VHRBsYTIqUL7waiBLnPEhCZkzXNPGy24vHkzrz
DqQL8fvHeyCB00nUqI6b9mikKBKXcPD5GFwT0EHFGZ0=
`protect END_PROTECTED
