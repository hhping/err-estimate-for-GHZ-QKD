`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XFSDV3VYMO+UO/v9yITuZ3431ZPQmt9U0/tcRJUlhT+4YlC20L5A0lLhoapCt4cl
yn/u5oaGM/yAKEMV1dqIn9gADITXQTifmYWf64noEg0WnN1JTuf/kX0Q8F0s8PAI
DnpiZ6/lqOEhpBqSQlBZDX2BkJTFxWasgPaW0IcjQm6s6swZIIXt7qZHPtWCYlsJ
A5Uf/oUmIAWosyuo3bKXCHUFlCO2kUcTgj0N+BAKGhBZYFHuUv1Lg1m2KSVk+caO
6B7qtc+0JJBBe3vSvsq1zET5NDit8aMMp/8F8PfhajCEs7jhhW9X8Ivl/YkSAr7g
9MNR5uMTpCbXqnPmePPjiFAbO9mbxZQPcEopSsGxX5p7PXeMkrxLN5M/hmdQZsEG
U3DWC3JCp2jqgUtRXB5kGhTcmawQ8BaaMjcDYp9NwKuD5qwiygsJAHNT4CqNg7R2
o7JompUKQdRGIxW3eV90HTbySObom8LU9KzgTqYvv6nrf3XgLTHCklvd2kBY5+FB
/jRq9BgIDjv/uZPu85KY4uvCPZvWQrRe8wCj0Fk3rHRdkP21qkxF5Em77tWmWHH2
U6JfuH7JS+ISVGJ380GgAnda7tKbJ15PdT7ZFvd4EIeE8Tnrn48LY4cyJVH7QHgL
5VRptGLcH/IoKY5ODgf/LG32bqbAa8j9TrJTaQCJbJM9C1r1A1cN7hqXXtsYPRB7
DctsnMq6l1JsrMm9iMq79g==
`protect END_PROTECTED
