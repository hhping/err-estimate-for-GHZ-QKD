`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sAt/KWUwVmibLBualptb0jiV22Hu0jbx4z0JoB4eaVVPEMxaQgd1uFstXK9gUTpv
g7y4YTUjQ1y9u41oyY7AbMHRLMDnliaGxZNV766rsntI8Qkvfl9vyuAA4uHI/Qs6
vnpzxuiQNwNEvfNsuByjhLsJd3thY+4V4vS7fYKNxAE=
`protect END_PROTECTED
