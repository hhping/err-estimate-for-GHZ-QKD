`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9nVC5bRi7dl2rcoB1qzYmj8jRH5MQMh0jKUHr/dGThWde7+KcgZf4wyL5DGWLhyO
RyXkFDOGObSVU09wC7c+2gaGkghOcu+zOdWIliqIegSZHfDNBvThceI8MRIwbpKm
x7LpzVVBrYL9G+RPl+viRybUGSZPWT3Htq97A/l1plSyIK4Z7ab1wVOTSWRizY/B
ko1VSDCCcfWmP4DdzFiUe1vd6+HT+onhZ3CBYujXH+Z3dSK/eBPla/0ZvhHoAfpR
P+H1yM7Tx/jCWz6HyU1/NT/GDeOwJwnC/VVZr75z61ORSPsTkZaj7DHthPOdildv
Z2F0JEq0amURvlBlBelOHj24KuxlfPUO33O1+NDVhjJs7WGq16B8vHH6SiYaiQW3
Ju4kvLtZ1kck4sHezNdCXqsoXrRtQ/Kpe0xgQwGwUjNGRtGF3DhX0LVb0iVHHmpn
NBQWhRtb7xhIeiUt4fTqxKzJswBtEqDdEZ3qwnDREDHVlVZpjMDagzg9v9E/wjcV
4qiiSYvYUS/uE6ZPewzTDuft1hnMhFdHWfPnoLp92rMD9aTGimVE+1NP0FfGwkmB
4CyleqUjtZJdm5+pl7W3hp+47sRiwJtSWCfvz9MFRSrmQHovpY0wQAfcJKrjb4Vl
3cRFoIkyzO9E+hz7mzLn7G/RpmTIto67aZHii89K8eNOtsYC+WIjIpZg0JZvD2vb
VJdM0Wmbv+OLqQZ4QdnCOKIEsfAQd3dSU0mqiMjff73wJnb+zzlfo8mpT5m9JqQb
ESafkunGna7Ubve5rEWQUIk9fpjMZnJJAaCh7SC4A6watQXxKsffiZl8u8jwHvJj
TlO+kksEDzPYsDOY8sm1zhtmDYv2lq63gtwEKYLt967xSfLVHiRt9/flr1lWnjD1
32J9T14RGeBQnEyzvDLNHoCO7DdszSUq9ktDKfgjlM6jppM8XHbhgkNtD5pRPqwi
HVyGaqr+wfVjJJXB4sj1t6rSshhMSEyQ7aXY0V07L5/fUiDe4kZVZO61RGVTCdsq
ilMMamyHyGxKfCWUS5uUAky0CnKb0gc3Z6qbHEKaIaQaiJRj9ZBd+9bEdU4Dipi6
mlUybwZP0wguPWU0siQlQ5DmQS1+ub5KnQOeW9g/Oz9NbftGKoBaQ6lpV2ApOln3
7huxGfix86XsgezXQA6x+mTKP6RHrQm9GbLnfbOGvYSesscFKyJDgvBIMJHEOKUW
fkfIDks2lz2EeSgDTC94ERQhSRzS7d2mVZXKFb/JPSZT1yptic03NyybY0Yo57aH
9b5Sxj+ZV5rIx4zFFD93gvUB63z3E6ei+/UDSjJGBpXLbz6peINhNiFMcuVFTIbT
tXDlQUlv+Z6ORAJ7956KH/tnawb4f858n7l2cfCznTUq/g+Zig+ChV3252zy6pWI
RdeD1oyXpHper03uMFwaDXfuLO851Li29WLx/kSzrqSxHuAoTT1fEoZZM4bDAowy
0yrfswLJtxutFYrthd7fe86TtVdvbKl+xaCHwul45iH2rnuZQ0kH43LqtW0UiM3g
jB3SZ/z246mz5pSJKjtMjTMFAFc2rRn/0a/SJxPLtC2TOzpH/bm6NyNCLzp2rk6E
`protect END_PROTECTED
