`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pcmKEdj8Gz+2dqgVtB7ilgD3SXVJDpfCGvvtndbEGq6HwOzl7tUJLx6WYlHDQgJn
tS4MQ18Al+nhX66+3Ze5tZsoziE29AbLNwC/Pr1kYCqLoGPTDrnSRAspZryWFaIf
+gjN4QCIoKrCaXaFavH5eqL1h3JapfYUrQOMbfFnGBYBOpjhvQQx7Cekmb1QtwVA
aAGPt7gjUtAwUFFrsFQ8mcKycLtVN1Z/G6A2iRQWXOR4ZTPkHmKVaUFlb2iZZOR3
Nn3DEPoNephPOv2CABQsalGdZgLrXQfr5/UWZJ97Yfm3zEMKhZ0n6qqtA3nGHFTE
b4ffDpcxUCMKaqWRNuL3ZQ+kOofN+KEY5pJfdOxu31Z9cFjRQoINfHpZB9zWm8OE
aodSTkxZfWcfPtf63krkwTJI+gcPFNmkGzPv183Kue4koATnco2EhhAmEwPdarHS
i6sEHsuHEjlJUWg+ZP3a3u4/t1t6KjwTSt87XsF8jXG4L30vcUfCW/Y5wiYNYatr
9p0t3C9fXycmAzItjwq2E11Io4J5G0+3chjok/9fv1oFbV+x+fjrlZnxsp40RGdG
xCCvUBw5e0Bxfbc/mJ3/kNMvPfCytUmyhS6zzYj9c5M=
`protect END_PROTECTED
