`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H7fG54Gqv9NXNsgt6dTN48vgCDo7AegsZJ8kWTwK0zbN7Nyka/rIeoDCEEVaTAR2
TF0+vB9Y4h1h7U/jeJOInaMZv50dSUBLdydFatwEW4jQ6sbt/km0rgl2yJRwGl9M
WJFcoovdmdfvDUbW6I73LjIYzIuhzgTa40vSpb1Mu0iGFLc9assGvRE4MVY7X1XM
cI1Iau189iRi417InRELw06Do/TanMimmYgc2SeB3ETYn6K8mt4ezy0Uh67S+uqb
rCgIcO7W/wEdB/L1e1sf54EtxosHU7oenKRAPD4a8IJtSUnYOPVq47ydq0uOBfd8
uPCvoU9/4NCEXwRPeesJwgcQHaLU6xNMPZswPrsA5Ins5WTbB29r1ETwXVD+iu09
tJlQabjBbQzpZMHuZBFDRnQwfijI/xRnPbj7qm/0Gm7zGndarNHOf66XDzQ/EX59
iKuLvSOEqCnwM0FJKqLgT92TGJR9RBWYvN1OiRTPiLtINVJcSyjhifR32tyB7Prt
zlmu+klJqEekpLhiQcYCPKAUZAGkpel6am7m+M0z2CN5DD6R8J/YdvhpPcBR0ghW
knrjz8QqBgSrSgvU71xtBDu1NsfwH5ksGNE0ivvYK1+tU12plXItLMJ9A76ss05z
jgB84mR4mJyeQbcNqvwz8gBBk1ifvkwc3DY98O6+nKsctH2kcrXIj4YoOQ4XZKsi
k9Z1zMifSYwpOtEYOj/YRVeMuBW80gkgQqftaTpzDZvR7FO4CaitNZX0XPzR2A2A
lOFzb4i5HlxCTrdG3pEBlw8PlxHS5E/ibsl41eOAyXwszX+ztrRXfeJrkvTDJFu1
WDus7llCuEQkPWixI5Ql80D+i7Jbb2CFuPbATnxx1e/efjzIYfUlTzQIke6iqoQG
/G9o4LrYMHt14+LI542fzo9YFIzlG/DDvvcwDdTL8uuwyMNo6qBf6yENVAPYNo70
UN0xqBkzp3DgR7NljLIhKWJyIuOdpbdKA75bVLKkjfVbKPH7zKxTD/SBYmBPjJfX
6bmztvidfZcoNJoi9meMaowAhKoND+WtAEloz4pBhIJPIIabdxNVzGk6U2Wr3pQc
b8tb6cir27YzzJygZd6WeWnnD2+1JC+Prtx1bxA51rPDYrSbVoqFdbLVW+hhs/Hq
NTCn85JVesheAg55+jnanEh76ro22QZIBpBBUdTpHpGH/JzL4RZLVtYrJvPfTXag
DS4YkFqhc8WPMarVISQIWJP/jOP5IkmqQ4m8hEpUyOGb1AO55rop2Weclkmcfrib
wtHx6/B/Ews8UJh6AWZKTp3MpJPMqwVBU76URZs5RyLOC0d4XzzHO5B4F0+1aH4G
YxqvUJYJUUtZlwGBINA+ROdaDLol3oLJou88A8d7KyrVMu+3zFbEE6c231ao8v8k
o4wqmxSwaHHiieNybkYPthnvwjit13iPaWJqv2h/RqQ=
`protect END_PROTECTED
