`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uUzUu6YcsspvrwLjk4Mt2c69wv0UM7BVr0QWdspTBbxPqLol0DvKxRw7n5M8+Nj7
4TJ+1HVF0trbo1hWy9JRfH0XDyAXUE9tjTPbZU/JA4aZSzW2JV8moGnzj03wiNvs
ID5lBF38oXUDSYDBD7m5IZrIqJBj5oYGC9co/aCljea01eVCcufhcuEmAaj1ITlT
u4t3uDLT0u3mr0waFiEb8pZ0w9wKo4x3/AzPdA19DbTSH8CTo6mLu0i8Af+EdA8J
wRHn7mGSsCkViMB0FI0gl1FybssZF4WqHEh4KMBxCKJc+LwLOA/5znhDylQUEghd
3uhe1iL1J4DZcAZnkwLGxV1vC09fELW5WY9aEpIsklkVtxPSGZqDToCd2+Te3AMc
ZwXfPPxTXxl6yIhrK2Ao11TBO3sCHwq49Ot/4TanpLFSciAZdIJeEoO2OiaoRcSA
KflAo8preVG4IRL7qZN1IR0n4iDYBKWVV65Ze+C9/EGkXLnYRPFrvj01sG/eeRQh
eJfKrD85Gc5Tm5srVLhyX1tqXxSj64k3+6GK7RrcAgE17t92pZlcK0XriQIUQXQq
sHri63SoV0Pan3ZlUSJBDQ==
`protect END_PROTECTED
