`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fYRMio5IH8gbndHkEqdvXdHPkDQJTtL+IJFEGLlPTrjPmDi2zORQ7G1lFWDsNvqF
TCHCjNV31/8H1iMsZ5qMX1kd/aLEt9koszVBfMhDOL43/mFzytK9zZgdi/WMqVEf
cKgmHz6d8FOJOJ0A0M3Rz9q4EHL+bMtIJQ70vVVa9aqLpuwFXfqrTF6Qx2ApJ2h/
qXkAA8aHrpGx4GMDlD/l2k4P5EadfT0tRHU7kQKWtJyjDJ6iPfQKUb8fJudojvj6
yO65VvhNv4L9mzLkjoz2C745cPCu3INIGmSKcjc+NB4c9HI7oT2EbnKmbuUTl5kv
LyuSO9AWVSjvqeMi9dJYMGqcFqWaMEiOllrJJbBYttKE++knRO0pSJ7Or+jp4cs+
nmkQKv8Uu933/poUFL5TnjIYyyiSdcx+Q6boxYXv3eqQNaBow0Vj5u50yIBEkydN
NKOI1qLDA4KZvhxAAF9B1AegA/Dsi/qWTvjmGtYD0Lfn/raV4M8com2QsHjRVWbt
ghZtP2aC7ojGVsebf8XvWbqr3DvQN1ws9PmcoE+tUvzOGF8n1rx50ZfFIZq72GdM
y9x4BY8JwitXUpxYOb5wX8w8KQLTy4TRW/w2H/ICo3W9LMRx89pEoq4RGVadiABS
da7a/iQ26oVsdCE7QWJbPW9r+y/rQvtWUm6QhlDZeqBnlAaYVP9YnY6pimg4PWm4
WOii6B4pLSlFBK8NVvm8osThftPjBuE+YfQpwItj08059jsPNZq9qQiVOAOj1jvs
PTphgufBMrmM1Nn1aYFuzdTQFbEUcRO7q+cndG7z/BtEZE/WOqkwLwWEFjdFpeSa
99QdKDEH6v17pxp5DX/arkWZxOKRFTqcVKgyR2OZE0MawW4hdnqV1UbR7ZL7wszr
rxhfq4uJzvN6sb1KGY0BugFEWEuGXuFPZJw+0bPZqlRpOO53xhjf1M9JbHinzes2
UByld4wngS7v+a3FclF5x3CqxzQRjX6/voaOMP3gUcYzilekYH+VA8iDmk5Ozt5q
CwZEf4FQG9VOumvhHYGYKyP+HfVPLQ4oKQN648508zGnAJK8/itbbiIOmNrVU86L
FBAvmV9PRnSwLuC5dnW8SQnWTpVH+eUi4sg32oVIEHjjsl2N0VRqx5r7D3BXYR5O
DG5JfL9K5ZEaek+4bb1905qas2ulCnvn8DO3PfOdHx7qDedn8UAfUyY2HYnghUUw
d74IcwfrQc3JZd51pZ1Oo2ruaNsgPABV3CwL/DsInHdWt3dbsbXu262zzX9pmCjo
x4EfbU4k6a08tQSmqfH7L5d2QhRUAd0ZjJX6o5DBJ/fZp3bZHWBIWDUOCrhwVbhD
BiyCRafs+z6SBYuO1kTA6cujswoH6Bmi1hG+Tugz4AXxpOSyLBu0X8SzDKoubmgU
hsUke4hotF491KG2c5SI6VnyNkVQrnC034nv/EqWf8TiD6uwLL+Qn0kNGGiliWOb
00CTE8CpWM7w3IZv+Zn+UntHmXYOxDe8tNyrut9DjsZa6Ogw8IRwq+youLMyJYMb
IU0J4zxhDR8P3TveernEcVb14iwIWFjcP1IRky3XKyN+ljlyNs8HYQ8ntBDqIZOG
e2NYrEWHKo5g9iPHz9rJI134kEgCq6iuDPkJMCdB4RP0y925tHde5bwce02FKIlg
gE2g/2yZt500ZucCIIO/D7+wJwlcKdiOtH/yQF8o0jGVK8Ux1sA/9lNfycgzle8+
diAHTZtqOyUqMaw543fzDn1P9r8XJzny3jHAG7HryHjJaHNdfXMf2d9PC6R7jLtC
abnnerO42sqKWvtt06IuGplkKT7Sa7MSpbFboZAIF1IPCwR6EOYX0ofyN/GQpZ7H
+UPQKFQyAKecEfE8ijyLwzrRG0XMaLAgZKgUF/tLP6itDa1SSD3RCespyVi+niex
QsngrJsShBIRS9QwdRsEvSJgkVxfFTBsD8qz+lkYPH+QZi8HIxLY5rDa1SvFuDp5
QMrzOyWsn9gVdMNQvlK/M7OkDvyQqYTzO9C8DMtDs4qUyrlR9ZK2V5jr5c7coSpW
VMj9XGUeFeTQU+BPektE3fkvUZkJ5QjqSUBTSZyYPXNpkGis4EguNJLY7kG2kNZw
2AJablPGRGIWconNYhcdfacob5t0UbhIc0SqorHbtQyNPPo1LVyz79S7zEWL/b9B
5LapDaXp10pBuwEqu7SVQ4rmldVN5k47f5YjAMKcTnoc690jTMf/ijbfLmP3NtR3
rs6p94UYhcbj9j/aJXhDad8BXUEmTfeHBb1gSxsFXQLmmUyQsBPyA7lgQj5Rha38
wngyvy7fJYkSYYRPDKfulsGn/TJB5UCNC4vXZX6mJXpiag2PyUZIOCmigtb4gKHy
CVelcQ3Z0C0Z1hE7QitXYWhgoxJkXQmHrA+lgCmmI2k6NJUVzDTbpQSXMDT6jaAV
VxOloVcpwow0u+SLHCsNUa5vfq6nt4j3xt8jgssX+PbxO3A4OZj1w0+e1pQc3ITv
VPxFimCndqjsZGNrRKyqnLNjhxKMPOkejBdMJ+h3ABBGhmDIabYjNS8oqPAHiOZV
Nxd9JUTL823HfN3DFzO4S8v1SeS8xwjXhSfT0GSfhpD1w27MT/pBzAsJAuhipGNa
xl9Mj23pCOqZWiQJ0nlVPS5iUSp5sFXfWgNo1Bh5xM1g0uWs4VXnPEX9uwzlD0cY
JZr1HA3c74g7OJtRwTzwdmyCqLwja7KFcl8OKm4tWghMTtHJjz0AI0SaFtYaNm7W
NU2xxsZj9t+GhJLije9/xRRmXjuFKxAVh4P1ihicTlUWd+HV+BdMD9wQ+QCptgTG
WzeOBfuwiBlCC9WJu6mTjqCepi2eaRCExSREBg/Fjw1GDLusnPTL/9Ees2xXLEYV
1X3xV8b+IKGrRIDgPLcsbtM5gDl4arj8DxYff+h+ec6m0IA1Y8O0Qh13F9Yy2dQn
1HdIeqe2hxfg22DDVM0yrdFGzjN6XJkDnIoHG73sZVtY/3qqINyznBKVHgFAMMPv
E4R/pCHfhnQYKPUbLFC0Uotbd8PRBeeoXnZB0hq6Sd0i9LTcPu9Tg0+fLH6cMxM6
LaSypN41axmjFFa8fz/h2282M0c0pJ5yZQhCE+ZJJVhe2fURHR0mcB/0EC4rQJsX
jem3pDahkD7oDIzPPqbRNSR3vR2F/dv2MqKq6rWeXsWPWLuXu3yO4JbwTIXR9GBU
/GgxokcFBURbVVxI5jGb2cE0WV3JqBzoDnt1Mgu9iNz1bNzHqSRzIJtODSYyHwV0
kgmkN4HmWxRw0sEpJKJFDUncJ9nMMmYJn/Seal5jQ5e8Bd/AfQ8CZ3i9kgDaT4Fv
UHutfzbu+AhseBvahJsfgN5bGJ/UH6xbC2rIGE+WkJBsMwXC3R5cZvQbHoxI6JAG
Y5BonhVask4+gkNaFFZ2TVB729uItY94A9CCeqByEzq1l2DqMJ5+zGXW3H3JS6SC
EJDTPhiRK5ehT8kmkBGEKYSgmkVM53fjzXLT2+wQkjLdDVjtokDdH1uzM1Dba6ip
LOGMkNQ0hEMo4ICwh+RpAQ6WOfDl/YiRcFiJdqEK+42rU7dWdkTPzUNRcfm2X6gT
Ma9LxLPL1ZslGa8kqnkMUZ11AWVWlEZjhByR95QiynM9ynKbVbimRlvVoiJ0TWPT
mnFEL/zY+pUy6QRWPF2w3uPn+vUVbdv+tH6qGg22zMwQGWA1jxtQgwV1kJ20Cp4d
9mRK/vHmkRqor1vSVrXDYaSOGtZ7Vsk/RxnS/1OewczwaTax4hvdJ4mA1as7MvTb
CGHwDkJNrqw2nhCQB9mP0IuY2QCEr/t76ZQJTbzoHvENHqDFIEhF/svpHKo9fQ9E
jS+F5CGNISAcVQFFamCK4WXWu1mP4dOcfCVlL0Bms7n3RWhGsflvyZ4Jv6xhMAoG
j/fMq22+G88p/Qp5txKMtNsopVJPmpaD9EBqK7vGiIuCHlw26mJjHZkOOIMOGiQk
TpNX3UYnX+SGFTq2ckAsrSPhsgLRdW95BXlBkJc5UuynAlBOvzdMTA2kxCpxLLpu
mA2nJ3DAevI5++A2+6dndzoYYsPGWfO608DLgT1A+sQAq9nkmEUZ1gF+cASUjRWg
Dn/xLVPNGXE/VM8RUhfW2zCoiyaxSSONguqTvsJ2I7a7R2QulaQDZoMQA/aQeikh
XEqSRu4lWtv21hy0uiEXiNhBQsbS6eqjjMYt63smzyddKy8mavxSbxC4LQRJjfxI
GpL74mAI5/Ask4BfgrYba9Xoiz6pPQdjcMoyKNCAHavqCKdflbUTs+9ccfFfCyMI
LJhMx4JSnayUiRw8RIfex21W971XGSpmKF967N193ZUyyAdshNRXR1i8KmnWYAi8
DvTpwJqLyyvoU+iUgoGuPVw5BHwC01n9SQ1E/aQWehOccLW9C/uxTbMe1xv3Nul0
OLFzAdJxH7Hrd3wpA+FuBkRbKs3alHRI7Q5r+OqezcWFiX1KIgPBfPhIMhS9u6aY
2AD7mdKSonAM1107wG3flspdV3ZAQCyEWx/OKIZsqnbdg3Jx6eYItUVaPlhrQjHX
4NZkSbSJERWDXhZTN8Wv8L8sJfWTnN07VIi2GWwziTu1vysP5q2XOivwevKwPbsg
kFTH3Qn+ZdZbAhG1QzLVVacKtFC/OQaQK9fjwlx3JiEaJiLWvLLeZYcnTkKpFqEp
U2URuOKviCO5B+NfpZIqF0DJ73prWCCjneM0OdniP6Fph3y26K7Orgdes/kZUXDj
/m9RtPHwefo6IbhpdA9Zno1rK9VvP2+y5lESLqHGjXz5P6wj1q/c+1bMhAAO/3kl
gkRGIIhIj6FcEEvUV0C1/j28znt+SU5rkjKJ/E9HpdR6duF2v7sV7HwG3wNJ9UDP
C53n+VG9VJ7xaIf71Qnp+OE6m7qqDNDQV9gJa/ZFsZra0qGUjPi9DRwkYBwFUxIK
pX+FgTRbTUlnQmmaa6YXQJjMsLPEqUvLM/IxH5VUVFHE2nurs0CroaeWGFdSwTT6
rtTfK5oz8wUNb0klZt/b9X7z7lniQNtOpppsGV1sWxQK7Ays1zXUjlYX92CC6qDZ
53uDnnLPn749l01YgQ4xzgf4UaNIOQ6hYJXldiAPtNoz5GmXqsCy6CVz6bSW/6ky
8dlnB9DHxBLdWSBtfNh13Bs8Vkt1e8OpWxx0WFGEnVxlj+IPwSVEaKVXU2cs+BFH
o3/B8DX00Xg5n12JppIL3rPxv/21EG5fqw91ESRJxZaJ46azScEtpojEbSv5hs5u
011P3XAbG7WvFfOSL3JcfC9Y4N+CXNpW+wGvruN8Ct4=
`protect END_PROTECTED
