`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2t+/t7ZYKmhRpbgIEviak6Ycu0BCmEYAyjHcadVkZ62PmddsK+P2uBgDbBLk1ejB
NuI1wXAdvO12Q81cDp/OEFHb3re9a/R9T/0jZ7TDrj3vU1c4lgkS8eb4oRNGqC7x
+ko8zYqIiB5R2MXb2f0J3jKr9TCx1olMg41yu66aUbpn08sP4WOUegaaBGbFyPbP
32T+48CBW9zDRQ9c8wwV/Fjig+OjUp4PkbYu2hesikQODM/ifEQv/BkLoYcxPeTY
6XyxynggaEvBLRcJ26DoTwGGy3I1fEAZmsr0tekuPxBuNm3GDuGoymCyZBNvBeCI
gmDf+3gvasmzHJbaQhn++zEMdWn1ZiHYFuSCiajV5+Z5VzYWhi3lEF5G1L1DwKCg
PzK3g8J9GsyoILMAy5aKJS/jjy6IxxFDn/cdFcVI9Up6CXHVI8LqaIsfn+hZlAXZ
At8BJzQnhD557HyxpJoOco/a2LhstadXB7IT2PzA3Nsk5lxcGE7mSlN4VazwgfuT
D/Hd1embYdDP8XTvJ934Us9A/QRN9ZT/JCoDfAZiaT7hWd1lg5352MtuPAcDJlb+
gzTjWw02+3lAKfzJs86qPmeW8Grr7XX9wYEGRPzvh2GPRZCL74ABawtBpt8ANZS0
7xhsjhNUanAmptoKZWqTbvgWGXqTMYUXb8NRjohJIWLK+e/apuUZ3a7USAPc7Mok
uzHgIZx2kGMbQ/X0XrUWGxjuSMV67VthbmRL5QL4cajVG4UUJ0mxSGpQzVtvYSdd
mrLFcm11uUXbIYvWRUrGBlZquSU+bvlhvak6qKbp+BGXWOp97xkoFRwjMlYUpH4z
cW6vtT/XpwG4VYeBE+dOrEOtAdFovcRnTUSnJgpk5fPdlNsH9ga5QGugcKzzJadR
fXMf3tdoli+Ypmoe20XBCeW0lbaJx0vFmgzn7+2j3SaN5bRSYO0jNZEuCQtVbvHu
fhxs8o4SEWGS9UwlkGy82fHuJBl9B9olKZslcSWNDSMPgyjYQsWjIumV5qk17P47
M08UPZND8mcYWQruHNQYpsLLXpCQ/KCkgJn99eadif2z4S/JYnEGJu+QwMP7SRYh
3GHL/5urMAgYux1Tae2t4TmcWS9o9zh0T0TzdLK7kzPKcJbwxsmvLl7dRVz6qLQh
uYTUYXLvJH1pPzSgz98z9NEBb9fjGXO+2rPjrgUT3r4E7ueBidrniHWdVr3BPMib
rOyhozb/iZ1heUohgRq82xcY7DeVGYYI70xwsmPdasrCSz5vHDvaWOqDVCZF0EbH
at8KpoOS6Ehvp0ju2zDJgp8W7XTroQD6G7cxPALSdAARKurDLwfnGyoUTFBXid9L
`protect END_PROTECTED
