`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QjaNYw4qzsqWPZ81pfp2bDzDqOeIg/DF0RpWjA/eyJayBNa4+87kgOB3OfWg5OUV
GQez1MNd8fflyKvzi+T20EwCQCizVoRbMSpOtjLDWV8Y9sr7saR+6ZuEiWkRMjaw
W5DeEU3GxfROSx3vyjy04VVk7kRGLCQE3kKYdZJWmuz7oRuCJQCS9lqF7JkvLWIN
5Plb1T88qrrBLOEaGQaU+uE094RqKO+rBslrOLFVW/+f4B6ITaH7wM+oFtnEA744
jnh4KXesDVzvPOkISC3mYDuq4zFH6R+Awks1SK6touLmmryda5li2H8T9hoeEoIY
cPO4wfhpoG80AKpsBYk4oriHvFV3lD3413NKEn21tLfJyrW8Uj4Pz9AkW5NmdhPA
AZsr88KY+Da7aCe/Y96FikO+OHQB6+qpsGQ0evDoINDEe9u6C6hUBjoVN5GIkik3
7Su1x0ZX7cXGOEWBaeGhSLovCAzTqDB7lwIneI7WxbjAYQHwMXQWuj5X3UqDnIlE
TszGcuiBTBaeEX493/w9uaIS5PoDYzdg84lDx4azrtrLAtZyPb1OxznTFl2Xyn25
0SzF1PzMrnL+G5lBTZAabN7b/oeJpXx5cDSS8T7cP/8ULlZ9agkeQPjmns25YqkJ
Ub3A32/3opUtQSK4I8ashsSSXjsKL5rW2+iCC11Bu0xU/qtzTFEZVVcrcPIQ8K9d
H+UnWWKywWIdeCiw8y0HuHVohno5JhjOOGpt5hMbr9nseVAXnErrefu/NmOq3o1p
wdC9lwGKtWhlwtb0TvWD5wTW9fknBsQHh2lTeempohM=
`protect END_PROTECTED
