`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8VV73eRjc0wKnszIungavez8y4C3CGPADIt96ncn/bJOI1N/fNM/xgYziAs8hJSx
6VdINTv+/yX7DiOemw9BApQ6XcFPvo9a3serqIDTCxNFABVGGhH9hWthWM0wh5CT
hZ2134fiYAkIhNi15feWwC/qxsTy2HXm3sJOPQUsOeC1hSmS+D8KCK7bWcxaTwKO
ahoGrdQ2Tjn/uKzAtgjoykOzx/5jZSJistXnmdeKNShf+pA3CfBIu3fJxR/6+zeb
IB0MdslaRcDS2EhvdBROwTd5A85xtXIeJudmRW/psyd7xcaW48FNUtb0ZbryViEX
6I0c85N0PBNrNw6Hnb7Vs/TYiqSaxpbYECV6mozPH6FO+CAhJJG0pPuwgQNcfolX
+a8St8jqa7oijP+cY8S7AhXP0Rwoj10uf6SxQO9e/kwO01bchHxkC+UNWZiz8tve
LgrXmzzwibDk8Uyo2EEYNCfWSclOepQDHDHPetAmwsl9ns5oyvIbludItLjsPUhI
iA6qp0xBEZ+iqCcat6hpvhbEZi2or2Yye3zUfPzawYY=
`protect END_PROTECTED
