`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NzNdijHVLbJ1W1Ebm8nk9tWAEXsp4J5hdLKqLZbdoybH8yL5AUXbkuGucJ9qHT+J
CgjGAe2xhk3raR4kEvN1V/GPjVtpFjGR63ECs74eLflLlHUuZsPz2YxhHofD1YmU
TKL9h2dALWdY26j43zthUM23d/ZLKM/cjVcxZol/rWhZHZzQtQsQnhU8G2c3m24R
cNDsaBwoaX9QQOeucglvfvZ2kNu6bMLLUA5RZlolt144/Ihja8lOteFwfOEfWbrp
3xuU6Jt/xQDWkhS9vvbwhwtiy/+ljuQd/GeId8egQmRzFfpttmOLEu1WtzJnpdLM
JMOBlqZPWdcqBv1m79xOs4e74fbd1EJpX8XbsxxekEfsvo3VDIBCyEfTfm4pGCWF
I4No5Ffm62BwejgyD1XKiqYQe1NXHpnPUI69BNSTDZlVWTJWzTbBNFSFJeti2LUP
Nzg56AvUdMiDJ2UrtfoVQ/QmCbuIQEHRwVyEXudnPg3XcXAStRmP4ClyK8zfK0mT
bNfoFo1+FfxQaKM81jIZMRCVbM5fAiYkHz7UkKeU23DnyLIpVFzG1H5dxZEQmRrG
OCljUA3onIB/NvlAFMdqIYGB/nM8a2zC0ofC9sJ5Qp5r8k0n2mAzdg1mfHaKtcaL
kR8T9vUTWns7cHmNrYQWez0+nojNyO8JqNFzeoLBXOzCb8enHXJDgv1QDmIVsjb6
glLg7G4Prst+rKCd7Cg+dcgUTXAQ/ffiT0kzn+JpmWZJbssLVJb4vr5KCGRvbQXv
CvEhb+PylXGn9aup4Cndgsb2phAXA/YHb8sdBfD91ULPaaOr60d8YdhHdr0GXwqP
tgx0HzHu1SR1XOrMtCiPeSpB2ixjEy9A+N8ZIYJcRSk45ZgCW4JhMBssqDEP4PGY
h10Fy9rThRJ3j64hfgMO2SpYuoTKsvR9d00PZ96gtDUWa7X1MZpV8MZo2lKE3yeP
ucuYkTozOLI8i64n7H0o6aaXzg/RzDPHpj8RAr39X2bRizyWEJjsX1bP52fv6dXz
6Ia5XxSop7fkxTknyY7ki35Al+XIwRW2j96/OnnSKZ56SnnI8yfCzZlJIlGSarW7
xd8pvWt1oM0EMelu0dZ9+MJLZZqfbw35jsplYlERASoxkz8l72y3Wy+Uta2SPvHP
fhbeFw5vymlEhb21cb8R9Kx0+guwh0IpAaFG2PM6VJDeCS+HW7AXABc1CjltWQpq
82JOnyODiarA/ppPU45+KQxo1Kirg+G2pvZKk4ByfDeT9JDXXoLijxnw12S1eCm6
grXWKHAVJkvQ8fwBOTpSqf9RpSBVj+BWqBj6WXh2wIgdU4MQehZbUIiOt+tmYE2F
gJghsGFdEJ3kQeCWXfEEbC/wYJybuOKOiZualTncT3Wyzdo4gAflIpPl+8/WB7cZ
Gcq+fj23gqJ/4Um6m/nqWTvr3hZK8buWOUsAIBVj7Mlz7AscfYpteJNQ1nvQJUGV
HyQkJJfqrRh3c1TbFzAZ4q/wF7vWgV44kQC4NLrUv5g7FAUDGcXTVDQASJvlNt6Q
qCaAIiAS/Hp6uChaI7ZKcWRpByA6O2EOxd8CCaecGswXzL3iAVJB1AoWaE4Hh+tT
SgTaoH/Ro30oU6xWEP/Ov+lM1uVAvwVYZTptej2FRSRaoVtclqZAecst9aMF5FJN
wrS0yFWX3RTyLGYwA76CvwU8Bfasiojrr1QuxCrYKxz0VKRaogrPK2U6UZLhs4Z8
HJ8TaozzxVCRD6wnI6dQvfzwxspNNW2rSsfYiIqEK8cL9j28wfNQ0iDlSP8E/WZQ
ZHHiclF6TqIXo/1BoqQojPuVcFus/wneswI/FzHQ6V6HhIMZTTZ+0fDe25eRi28W
HLVr1Fxdh8CabMZEj+G2r90icspyci7Fq8um2cFoYe3C8dljDqO9xD/xb6zXZ4g4
45ltKYZoXDKsxbrZOc1TpnYb0slo6xchj9JaPWVjj3h5hPSUXw+436jljo8QbGyo
rndG5L5fWVVTCrnSiWbvszuEMqGPERf9AbP0m2LcAa3jDv7Yq7cDkZ+DOeh4Y0FD
7DfytSq8pnVmqpEQBbxj/9hWa21G2Ojz279Gt/ptpLlBbqU+d7gR1A+qWdMULYQH
I7c+BWfzD6ttwWTgMJhukMGk4s6nK2RMLIg+a4W3rXRPDadTbcIAUK1hS5KkgViH
DQcsCIQgt+A0TZZLa1z6YFEOv6BM1iy/0t+GBFsoQuu5PHgGFZ7qf4uJEZsyAoTt
ssLEKu6e2BT791YCZ0lNJtbtUTbcsmXP4psL+YLfbgp+gM9GBUoIK6xIQQJHZEoo
o/o1of9/SiwNzTODLzsY5Q6do6W4WHpFKdgYxWKcAJen5A+0oVWceCtPhUAx/Ex1
JNiw8pSRcwMVjIj5ePp7mFuo4MA+hgpJSvS3T4QA9fxvE0tAbYAHHo33rDKtoYBG
yWyqpQClEJ8Tz8QSsyl7/+MWCVFeg3IzEzsxiLLtw36rGGupcdYBTzgXX8NQfaVr
RGCUK0Qh08la3e333+Ea7u+XNzIvLNzkvDQ5/UhYCx0OIq5hCR8PIpQXfwLoSx+r
qVxx2Xtyyrz/gKfBcyl8dAX2Tj7/M8/Xwm6dbj9+JWROkqpSSW5bdhqRc3aDdRxb
0FxC4e7PbSXQLBzbBZSVGSULrMGckC3WwIAejuNWxnUqZYVOnSkaDo6pKMvrhPnu
zqSS0RIItjid0igcKdhe5DIIKtqh5z8FaSfLAOBnuVBgvYIqZvZ3/NDdd75o+5+3
uTKx4Xu3qTCEN0lLdOQX96jwJE0WvE0WEX+1rRs8Nl9NWsls6TEgkdG2oGoKqW+Q
FRnCafDZ4Jik53bwnwH4uMEnAmryuB7sBUy6rW1OGBMggEQCDz/qbUaNybegkp9i
lPaMkvIEm8xGVL0vwyKDYfWVPXaFJZ6PAKlTIMdppMxmDAUq3eZmJTch4akqRcNz
+u2wx8zn9VUg0fBIEV79aEEYaeJm0T2YjTT9S+rfKan8ZXVd1qgzPr0BKiCqU02y
blCH2OMFnJAi7EHvN0TkQ0z9SPewu63GTRSiYUeEXsBdwd+UAnpouul70CcJjxIY
gIk5Caeix/W2VqzPp6uUzc+AoDMy6IWLvt5rYDl7d4aAfaKdCSyVqxwcoB/6rl99
P6pv0bM0Bigk9Db/hv5u9H7UjJrpXTidRAOrATV8kcTtreS6MGNsDfDF7lSQ09wk
tKSvRsQpgFAJT/ku3xFgsT+5zw15oLS6I8sDglTzLUdloPaWsZZtWucLUQHbaB37
iGyK12Yz/DJPj6KmOUs2QEFZdMgP9+NfAw/+iecDtQ7REEaGMuNyk0JWw4YCfkky
z0+IqwPdwcJy/p71hnb1lsjSgl2/PrTlGu1hXAF5aOcs7RBIQl89I+I0Dyuy8IP/
BYCRJjdOYWwFaLG+JNFlg3CtdwpQs+8Gl/+KWs9k2wQQUM0IzjgtWONYQqQ5FWEW
Rtyn5vjDP/fZhzbArBR91m86e7dAEnWKLLAxhPQvUk7pAoZ5Q67gS8XJ2IvPSEeF
+/fBQw58cPLJHDfM9XjjuUQFd8zmUH017lBhGfYJeDlBRaoOBWFwojziygrb33xH
qBBEQkw1AHVmfNkgZ6zRnf78YdyZtW0HPXcdeEnSlST/HC5x2wtGzfu1LW6vsx2i
ZveCL5rcMOeG8nolCtfqlaWvatZ6H8HVddqpCVRMBC+T1gaaYmZurxIVNhmyx8vF
Te72CqNZKpuP81WKquIJ/aWsbHmfUGCJmxNZ6GJl48pKYs1vKL5NLIvHlr5i4Mib
L2+7jdZa+GnVJ/2S91frqWnMQ65Ju5JzgrzD+kHiSqrBKQBidWJMbhOpaIb+RUhP
l141QZNXCAw7805x181zZAQ4ybRUkXXFhhnG5yhezicizzf99ylYO73FuUsUBe0a
m/KWzVekMbtTngNvJWhdslapTNj8Ie1zXLp4RV+IRhwpznCqRH4TvnF1xI/7Fuqd
30tnTd+zgRwclk2GikkGUxBJTJh3CA7U2KZbTyQKePowh7I34k+BUiVblHh0ZUfJ
fM/FBkG59mkjet6ppRMD8G1+qJvXDwVkpG50LIIRYdDSKu50msdgSS9eBpv/Hcdj
CXVdre5sdrhOrCIO2t+G/59gSVv/IrEQp1xB2GWX5Ok5Uo8ySClEQHTakhjEk85O
BJNKY1sjsW7MntjRhogqHfcVE/RL2rgsqE/hHA4GHK1KvD+ep1ouA21JS2Q1P8Me
RJ8wJoFzyfm8kl2IkxB8YNhnUlHtDvuBbM9bZjGYuudbkzgR6GxgVIKZacPovowb
JhUB1b29sWEdwVlpCs/TzUkTznO+wiHrTsDWCgk8tR1g04F1lBAdeLjwigwiID34
QX5dAhY/BcV9v+RxG0nqycFWvIvWx3kzGA/8KWliNbgKsdz1RieBbOlQrJFI2r0u
dRv6ypNiTZAvhOFNbMK4WTPFYCj7FAFFpwfWTWkjH+YtQ7zForRIBI6T8Z4AJi1e
7wUEAk3hxQNE2exwWxUzblujGtjsoUA1nxPFRY1JoppnLsgYcM8ZwzYtlbZs4URK
83yS3zzqBuD0e5y51Tfq5Clss20PDvay990g87I5bBZBALHF/Toi3y5GpOhvuXuw
uE5w6SL79rptLbWxMEdsaiiFPzvCD9P2q5qskeii3LotnjfSOt8LG1r5BRNH90lB
D+SvPz+8STW0svjHxmAyup6Da5JcnworL1HhpvWQeO2/nkC5G7vhhhZnJLzLjgDC
ZQB5oczgkePE77QesKxgAlR37spOW4hp5fFoxCaqxr/1rCLIhs/4hhidoZbfF2JI
0h3BLHnbeFPCfOEhSn8n1KCkPoTmnIdai1qXUS0cPKFLIuHbfu2rFuODS47QVxSV
w2zQD4YhjIvi4jruK4YYuhYPymhsGV6ANLQ+dLSMtb/Rq5xC7KK/sxIRiX8KoeOu
BI2beLOfbeMvZpKB0yw0/78Mz9KLxUU5AOUjVy0DvDWHPJp3LCIASfN7H+5CVdgM
T4N1OS1A4qQOVo1NL5MrQD2Z5C0+kMdaG2dxB9V7rTs6NjtG/mlAmuyFDjp4Ebad
VSUdcuApxKeMqWXAHNHE8OBoZMxAfzYFjyPYxoD/vPOpXCd+tQyAPn6tCAVccxKs
9R8UYxCdjcZXKBhF2CwWIMbi6HN68KxiNJzfRyqQvNn0YJJbPqEYzBFC2rnqzRkE
Y58n/Tchuyr9Pi9zlVWsVPiEqz5CJN4WXHNv9hkWwAbYo/ozA+KrcGoaR8kIdTKC
wD3DaGBevvlmE9+G+r/bBGneGVvlz9sJCgrx2tOXxlitrzvTPOgO8vutrNEd+mxp
V89qHt8Ll9HXJRP+8Jt0JQkI+AYPa+8EPOgJ847eL9kQm+uwUqvd1VtazvD2EIl3
m/sMF64DU8GIHFLODtl0+lfqxGQ3aUNeW6hicqO7q3hD6D4JyWkq/F1KBrN+Ejz7
3ULIHMln6MUKPMnTpErs1+IUKqVkd75svdIJcWHRHw1004MmrzV22kNtzZ4azGkb
pw41mrZe7DDUTfCKZTnkKpCFXD8Nku/j6LvdSyx4qgYRtw2MeyRVgvfS8+YrZ13w
LkSSC2EawWJK3g6MZ65m0tPtNXkiYPRsTaYEW6hd0GsT2ZcDzTSed7rCUlpImGst
SQj7e6PBWB4B3MdFfZdvQ97/M5yN2m6QkwoLX8sBI/xfduiT7+Lrf7x33kHwMb1w
qU5PAiFbQLBiYmbA/ejasG5pyxV/eoEHM20PDNvKK+jlrByO+CxMFLIWrsvSdsSR
DScWDBoSZ1nnNp4K0pJem+DT7C+ZcSanTaaLr35WKseYXTD+I8+Ni0o6DF8yJaQr
T8nRdPsEANbs9xKvVfGV/8Xnt9SoWYcFIVExeqM2YtAEhzQI+oCAoaRTZng2rZIt
x0hivUgHZj56Lezz+CJ+NTQFPXCesynIBm0N+XUdQZfUoLG1lrZoQmnPr4nmTAFc
scZYVOvvbWL83H1NJSjL1fgMnui4cSxwdDys/IfjBY0NH4s4cmKbWpbjJI8RIX7M
WWeYaY4yZxl6ZI6PAel3xEOQAN+T9JE+WMc7As4vVzOBqzZMgOT5IR27ZJbQ4iru
+c9OT3DXnRmIqOUYHJIEhNIpnXkgx5taJRfAK1G0H2UZINhv3yhlFU/FBMILubn8
R3O2cdRE3SLnQ5Ld/VC2Sr5kWjmCCf2xgN9nwCsP6zI9679yXXhkX+KU556x52WG
ATxnDw1rrT89oSuH/c7nlFXhJi7Xp6wTD1zn6VW7sArAL03QH85fu1dRxXUubwT1
yBQ8CwLjbv/YRyHl7vfvN7B/gJ6XIeRXUPc/5yJOErZP7GzR3Tc1wNR5I+0ZZ4m/
GHJoGDmjMWr9dywbS2R1EnCysOxTBuVN73fgra7WuASq0mlkl4n1LI3I4UtaSXrb
6tiMWaBDa1n3CGaUY0LlhmtcqLX0PKHRsbekWSUAnBbki9X6TZHmTaUohANUQyLC
zu+5q/XMxJP+if8jK0dz06BeJA2llLWnGcH2fbyZzCAFNFst6WUV84oOfq7i5d47
UBnnyFHDrHb6T4+FJvgnLuHDu1ydbvvE0s+K7WWkZXSA1req7skQQ9hMNmriLDeQ
OljsiWqT2MrZMNqGayvZbG9KqU5clLTEjbJjgB2omBqZkSf2d7vr4rYKLKkK74Z5
VFL9cmgiAwPLesBuOW1n+hEpDe5QfqRxA8zq/ifCj32Ln9YWFz7raoTbHZEbXNgD
zjaHeEfebxzI6uWsPQCYiaKK+TgJ/1iBF9pHu6VT+af9CO99xIcemee5fUUfkOTK
tFerCl7F3EocQH+xPbhLPvTGxk5iQY2uspkF/rxSQnydJ39R5373J99PONB3MwYe
cvr0K7nNpxPoSVcQh3wb2xuJC5Uy7rj4FQnVkNGNxs9fZwI1ViZ5fv/l+tQ8G3cB
PRZsedqWaPudFv7vNn0gVxroOzT5BGoLfOCOmNBotAVyM9nPUS2tbS2ntyIl2umu
wiS/xXxUfwHIXkhhdv2Xpw8m6pq1pQF1IuC/czs0ROK7IABdFN5PiWEebP9KgDdR
gq8XlRBZktTOS2DN8Auz0HZ0bZSqY5gxdaiqo/1JY6M653gP8wiaU0HogtBZ3hwa
flX1B9ufkpGO9d4NSVwf+rAQDgOXGQLx/mUcbZ2g5mKWzqsOLMuZbhHYGR7iaTcD
pqYubbxhriv4PcBSw+BoQimb1ka+0SVw0vxdqmh+xMruyRKjC+eq3wGpiUkgZcAA
l7fgfhoPcrF01CumRz4kjA6cC1HHbeK6uQBi58gfVLBbMBZ2WTWS4Cuu60nxxalw
gm688pIudnPePcsT/pUOwLWyQHl4tnk4AijSUSaxxgMzwZpbyEU/ERG1gu9OAUE6
UY7gOlZCHj7w9lJnXjA+zeR7FnQh8Lt/SdY/n1AQcICQAMRM4q7Hr4+H0b6V62xY
POzeH2OdkwdV7GUf+N4W2WaTErcmXevMdFfCMUta3keGIs94jsRi1lu7j6Ge2cD2
cFBLChKjWT9Ykki0xx8ww0pRYd8MGajnDODYT73wJQyentL5G4S7HEfJALl3OiQN
eKhgz6yGTuuBoSU+V2ITpUXs7J50Kmhq0d3ep/zYebFyKMlXCTgShYwB4/V0SO9q
ypQ2xDPF1dIAgdvbGiBcTqiIMYyci26fD3qx1ob4oDYbpyI3FwMnXByKhaAg/SU9
ts7cjVAGWd7IpDr8NkgalpMaoXyEg3OExwsYbyI9QNRvhLnxy3tzY9AogxrBtZcX
2m7qfaLKeLDB0s+4MevACAiFaVL3cHyQQeTyMSnnO8aDAYreftCyKkdtz3JK5BmK
FIK5klrSDBNQbc0ty8D8B2aXFmjRnQFZMNkTv/ImH9Mtn/hjfQVQ9bQ3leqq77IO
ofwBpZe66SyF9BSS982WpcDxU+gcqUV8FRyQgWP+p/rAnqJwRqmy23dxPh+VDwy4
Uls02PVfsDYepFFsmK91bQ==
`protect END_PROTECTED
