`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iNufpWDICrt+siwiKwWm1MW6EbCAPVOUdbbeJjTPxkpTBTOu4INmw4gOHZyUa2Qa
hYcXQEtX1dnMW+XLKMw1Pf2EdM5Xi9aDc9GMzvpy1jjQ943fOmAwb6CEm0Z6W5Hd
cWY7XmlE/vTuW9A4M3SGaFivRVpclEdFL79FI2A+T5XE0WJ2qjx3KGpPV/GfX2V8
vlcVCoGbZ+utgtkZSPW57crhOiq6yQXSkxNcVg2mbwaIwW3tG0RmErAO0EDOdoon
53aSoi0niXiNyz24kqBOdh6HCNnLRZI/DdFIbKVt6MTSyMcDpsJMmgLHPtvYmEtv
gmDXRxUjBCwKKyw55aY04uwj4JilVlRgOPA3tFPw+Ha1t9+GjB7tEXYBQnZ/jKjA
3I9mgyVKNGxXAq5Ar8NlGTeHbJTpX+vpHQr6AnQAi6J6R78QRAroizLx5uFyC6Et
U6HMF6fSzJKqRrbGdh3SmAg1o4sFpFLqvDzs3P9wARy0ubZCiTy/tLQIfrJhWaFb
KFr3HgTD96zuVFGRlC26k86O5sWgPMKnDYTwRHZfP9X8fy1D6rV9hCHNGWeI7BwA
vsOlGeUgGeEYcthtyFeRPhiwGAXyH+jtTqthCcSl7Jj7RX1iVvCfLajUmCJOFyco
AcfKd1qVSd4Pr6lIrLJ4GHlvI7TUQ+Z33HhdwkW/beOZ+5xM5W0aurM6U3Y41wJS
WIleVxlhpOEyXvRla2+7XFSDuwks2o6v8aUbg6YITb9E1Z9zBZIr8S5nm3TTHv7q
sP8dumoLCT5WRINMCH+Zwqugbr/4BYXuYGW479aHqzfZdNNfmjh7qyGsbzhe//UC
VAnH+dTJYVjwYJyYjjpmJRz5XMUywQW5jiVJM9XVNlFzPpBkwByLzzZcX5MvVEAa
sidt/vIjXN/Fd/M54RQ1f/b0sWVG5sRSqN2cPB2BvfnBH/CVhWpu8jMIGYHvl9C/
uxJJOCqdS7nto+/U+vw6wFtgyaRgOtwHnZErprpcJR/89ZaaC03hCAu4w/5NfGQ8
NEEYM20r68mZIL/hXBl7P6XoGUZIdDYb4TM7CdH+uhGffoQQNXhhtlwQhauP7MwL
zkKLxW+gpFwEyQ/1n+wwAPwNzmwh2t0bNhQOP6O29ymUK3nOIA1vWBn3ej+pHxIu
MhOplbGUuueqc3Zh+5wP+sPww2j5MhqS/cTiB6lktixMauVMvS6qsITs+HhyBN6T
0eJwmIxVXI8bkTofsAwDxG6eZQ9ihL92z1z2QGAr6/qze8qwulcCdccTfQj86QtL
INeAQCFaZIm/1EtsupFjUvGYrD8nlgQG5hFnegIK/uLqbYztcHcbJa4w3NpIKEnh
`protect END_PROTECTED
