`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qqXS/M/OYX72gLzBcGPcbZI4I+pe4JVHR1fYEj/XnGHDSyf8DxjMDDKZLWp/rKJX
IptSq3POxNBIvGAOCHuXRCTflmW3HhOKo8V+ubxBZ8o3216qQuzemywNpgRlY8ZC
eajQlT3JVIFiJn42cDcAVbOF0dMhVngUW2n0Ly0X4TTfGvAc8WWMJe6XsdxGUY/R
uM/8XmrRLz7FfDUMH9UG4h1vkPYqf4r/gNYKBTAtfJBXep5V//GSnrWoKFQaLZjZ
N77sloscIDnry4sbg98GbvXCuyPN319AU6R6s44yLfcWfK6/oW3qQF1hG+re4W/6
UGvuxAPlOLQhRH2WWUvPp6NfHaS1BlndDNG77EdZy76D8DcPgblo8Dofs2Zlr1Gg
TRqVO0BraqIRfSnpmnwymEAY7RWZDZFrEITN8AvZU2EXbEG/yj8OVvwL+l73aU+u
yXhBtJV+6S6IgZUN1ePTT0uMhKLUliS7neKNGaQFNQuV7nlDzKpi6x7F2WdX3+vz
ZDQGyeXuIwDIMiCdJM9maLosd5Dg12n/Enu2wmlFzYj6N6GBbXFXyrW1nPLTD3kJ
iusS8YMWDAzACsAuykfq688LPedYz6RhJUA0Ag0ici1JHyQjFc4m+n4h55JieTC1
76UO6CIvzBbyDbc/l4tv/CYefUh8w+oGNAe9lgnPwzVskIaDttawW/pHSWfhjSJ9
wGP9xiNt9mNEvcdqHlr7P1GC+UTO/c9I2J6+sIZwDSfchwP6gcOTfEvub1rVkCFV
ixFpy069x+IBrMIlTKx1ifhTZX6MsNy52cM3Mf1boIhnIB0xiYnwzA+CeVsWzfhJ
0t++sECRlC3P/XqpaHaL1+rAOiYGrOJNPJ9hCEov4r6e8L+WLdjWZ6DQeXa3cqwY
+4G5RXRz2xvOL5z3ZzEAMnwUEn2kpLg3bjfh6qzSoAjaYoEmKsr2dUaxJCY17qsI
URK7v0Dj3wCfN7maG6qP9l6aZR/Ha21+zuPDeb0NOa0QmctGOPPzTPb0NrYXfAlU
vCzSrnkr22L6EaOoWJpt9VMozf0it7k+3E9GQIJ7m+q4WZh2MBGOex9ruV93L6Am
rkpEIpPydVbTUGR4g8SATCafUkLJzHeYyql8EGReSWzdpg0w57tJGJtaeMEgh75g
UP2AXLLqs1TC7rM/a6cw7ehJNoroHwFupvlsty+QWIgkn+opWGA2+iruaTkRxkUM
bbI1pb7WaijpBzY87gpzs9lcWOM6Mj6+hFQjWdbHpqM=
`protect END_PROTECTED
