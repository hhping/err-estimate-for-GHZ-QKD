`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r3je7zkTq3Keu0LIVahPYzM6iElOwLTnfERlI8R+tHLgxzZVRhHqXKDii4vOJj+I
EQ6rGiyG6lIup/Gk6eyePxWiJ0EgtRRSpE05jw3T4SaadGZf7GJ8XhtjLdxfaKUD
xpC9tpl69cKc5FbMuYMjwZmm+XSINlpetvE+982hUcp59Y3Z7Q56lXHx7RDhNGSo
qC7ABzzIsYONZ9mZ54VtcCGdq1U++GnS14LgPT51BDAZmT/0v/m6U30pRAVJClTt
t1mTgEefaDkpxfSlWa35YtMhvNuik1S6TDGOqC40RH4p/G7VMH2tfulheuq3k2VV
lY1/VIc4aTp6zLHzjOHQPB9c2Tge/0d+Yf5N1gjxjJ3RQEr8eLRl4e9L41KUfcMH
UlqocOUUEn6pjPCWQuBqaxVzJrQMvz1R6P6HwyYwBaiLxqQ/GbRMd/f+zIhGSNzx
ItoZ6DyNJorppMqfKCXcjpypyEAHY082RCHGnGCHvY4XrYd76O+d2ZR4/M1t76pt
JkIZkHAkL+zkLggZ7UjLuFrUBpaAYyjEGqH0aASaOi1HMfCxov1MLfWD7hfyNaqb
bQLYnIsQAHizkX89A18nOW68kDP9t6vkRnUBuXNqOom/K+gtbbNkOVr0QJYwocGC
OCDNo+/jVn12msgJnz/lBwODDBegmD1mgW+hLls0v2GNrYKvkv5aNe4sGp+hXeRk
gF7tDGEpTHx33blJwHqoBvZ+Nqc3WwqGUiuiSHqJoQzbojyjwJ4pjU+I4cyOl+YG
7VH926Lm79tcamq8T4PtXpHVoka5bP7b0zBVBW0x8PgLPdmr+XWgVk+yNGyEU2vJ
CxsLv8kHfRtjJrslKZmSt409DfPj0dzYt7VoMKKlonUGcaSURBkgsjrwLvu0dMtu
b+BHDhRjp6dcKyGGYBhtLTh6iAVfXhXbgjakh//AJUQimXbUePsGngIQZu8obZMr
uafZqKRPrbwqtEB5cZsv1LCxz0z9kcBM/o0ZeMEBHaJ1S312EgG1VzuDIjOME0QM
94IvtcTOSK8mY47I026pwgdkgvyX+DRuOktIvnVsnj8W4MD9b13CviMTjLUbEEdd
oqXbgkMtTIvmJPPzOas+as/ZuR9w+9C7TpSHG62V1xSi0wsI+P7DrMHuYXaq0MQt
I1IAKhdzZXQYRA5sNsrCZ+VmzFR7atQRg1/QQq7vTPJiIvLnShMieV0A2UieIAuH
OPo1BFhNetg5lMooEVV0XuY9NNAaJwbuzKe/Cyz5B7pGUMhrnif+/eqqd5ucKkOR
wZUm+HJ0bB+soMht7Sok+lRgfB9/LnwM6YW3OcihRU98R7PCgzbuUcrUP6M9VwzP
dTVYnUKqEk2+DjIl7AAh8WaYzM6jk93xtVlrz+i/s6EAxlNAuAMsAvh1e0300+w5
Gc/dmhugKQCWB1vVt/Ern1uX4dJaPPVGpij1KokqA0a1mAxmN8vUbXHcfg0oxxsA
GwrhVkw00mTMPQNWDR+uvFSBnWmYHa5b20+JmsVvYYDd0P+7gHJYVrZuxk0XvGRb
MYa+5fWXc0l5FUWK5aTWDt6nrCOLRoPxmrXC0jrCHnia4WHTqww1cyLZX3W8xPbN
K44Uu9pLOgYeJ3zGVLczCGc9V8kU5l0kXyq29w+xAVBVeWjqSTbwrUGjMbq+jPut
i3q0vIR+7tZI5Gxe0HTRd/jo8mQXIWGXCpHwq081wK3+DlGiCgfYyzBOHGVwQ+5j
rYpsDSSNREzURP59iY+jKcEKWlRDcJyF6YGzESve8jfQRKUX8Fde//t871QpEgge
gJ5F9S/INhh2JlU1ytyd2ulazaM5+xDbXty/rpfD2hnH/hbxVlktWULm8W6lKUWk
GVZdb0y+ODY8Nqj/mLPyhCSqsPxRxZvEe23cIBuetm+VT+PCT5tZvnbwThPG98el
dGlMjMJ9xZMfLX+meeGM2UGegYhokap2p8bjTrvFKNG9XBOr6QSq1szwz4Gei4Mz
j5bWd+QcFq9lgGE7ZrwuHLEA+/sgq2ScsazwCvgPs4w08pdqwJ/vYfFHYBCHr/GX
5kFDzJlJ6qy/FDnLp3qcN5nuZ9/J7tRSfvLIWRMkB0B9GJ1YMHwOKg92F8nHCrgT
72opCufaQluql2HlE+DDemnAvTD/MtvBkvm+jCDCdzJc9b0ZSThnKxkW+B9idhKh
GIAwUs+T285zWwt1nnxDeapeIBtWYwQwPl65bDd3SfE7G/EMZzPb3eJQm5DAwuen
DTGqSMZCfT6iPt6iU4hPWQulWo3LqyY9mWFfKDdpFgAYVR7tnam/ICwUU/Se+fwh
4QkcQPvEvIWjTadpJmOUXSM3cmP3W30EZJTdb0R9aPOSg4fdOL42PZYf6PxZ8DNb
H20ye3HfsR9cnvil9MPfIccWlzl3cPvo+/R2oHJDNDmneR8xEteRvgg5u361WZoS
8rKpnixy5quICeftgGYCPGrEg+qzcOZFPNJblkZ3em0157k6gTKOQ2exir+w67/r
iznMz983PkDDyQ6g6TX2KcXr6CHHHxgGhw/vxZVAjq/+bXX1fb9qmwQj9UbtEQqb
CbhJ+UB/LrYd1gNdpUeUW6kLuZlHW2oxLwItRS4DkQzqoJ/DKdRluCHfkcLM0QAF
H8ZcAXonk8F9Opk1oGn5efTN3r5tolvaRMWb8GH3su8dFWaKBBH3Uf9nkE4ff2q3
olUn1Zrw/5+SV+kJ1y7d7LSyWJX8MAX9REgbUkWoXtAVMVYJOVtQZnQLsTgTQ286
ysbE3NTwiJ1//uyO8pu+Z+nY4aOhF8hGpkjmYUTU4UhEV2gWJ4UfUvoBMqe459x+
Rr5BsnBCpyksI5Xgcw/dLre9XxdtoOd4OPExjLDIk9djoz282Ytu521CjD6FfUSX
/Yvi7EwL4NyO4YSmFZPkbqYIclYcn588TVyDDn8FWBHilbJp/KqueY0MJAZRyqot
4+I4cFx8+rE7LoKnURSKAy7CW4cN74392VaZ3qHNWYNjckp0UBurac0s3lWPvxQN
GExLGhAU7PPxOKGrwAd8jJVB0+RLAt756zRtWNzKvk0MxaBxlOiQjPTqtC+JuEZB
gjXFPT/NCGgydKjt8oA8eZGpxOmi09KcMp0Bk2QuUz8LO0+g4EYvjrngFg7+EMxx
yx4EOuRH0J9KbdJU/h/9GtgF6kcP57VPuLEamJxyfB+2K+F0oKa/nQmCX2UIUa/X
ttWiL5MLXdtJmuOr79oCvsnEZpbxrkufrvRWx9I0oLMEiOD4oQxRkvk0qKZMXAE+
bPpu9gqxzD/ePH8srQrnb87WaZlTj2yigLXVoQH5xxUeQNjnXj3HeiLEblpc5PCZ
Bgap0VjAdBOHKewADMNh0sZK28gb9Yt4KgmMJ+McHt4wT4rfeIn/kNTfmUkQ5WMp
kfLOlDfs88mH35cwSGNREPmF0Bv3UNNpBve2w7OIgSTbS7PX4RkWXA9NvIPc77Hk
aM9DuLIwn3e7m5Qwp+VIO4DMACziJxm+GQPGauFs0ji6lL6PgVHMjNXrtV/G6z1K
Ris81Eq1b4KHIQDu3KuAb7QkODDhLKBNIPrNVcH23NtM+PisjtnNTEax+/TXu837
h7yPUHNwEMQRYf6O36Q3mMcHcg8dXZesh3vtv55vxVTRJG1pTJHKUdUgKmicucUN
1JSlufC/lnhm9JZmA0sz5W54YxH9sHEb34BVFbIkodIfv3KdTa7cxKD/ylEEbKsM
RruDOBIfcNC27l+FOG4C/OFM8CCAyQSvkDx5V9MdVsHl1fZAIvSA8KXLA3wpfZAM
+wScouRbXt+dGmMbf8G3APg2euFl4vacRLy7DZG5j4wB29qdkqdznZf4gp9TYZtm
SHzQjOuoSdjkuEHYUlex8owcyTNKTZ2laIMGqE5B7+oWeiksN7L5qwtJ9Xhx/wqa
joWnrJA561r3kpou+u8w3DJKfh4R9oWgvgR0pqb45opUsqTg1UgdExufM+WsA5X0
Jy6l0FUdSHWmthuEUEr3nv88iudWOzZd6fTXngjN/6dS2+lRDKxTHik2Q/EXayrY
Hxirp1YzSgimhSq8s7jRITfurVjJ5KEjW9nk0cgOydggJ0JuUdRWyFLRGhZLTDX8
vDWupdhwbt6KQ1q9po3eAiFXLnx8JQG+FjYestRz8FNoOeDSFWMEe4Qbq/2gJGQo
kPdKtKeY6UTuK1kj6p8svD+00o2L0D+9BhumRNfrY5cHKIJVPR3NdWS9AEPtR3Zz
r5DDSNeqoZr6C0ZyY3QfF9elD0RzzhK/Ji2SgM/W44/CC+58HhtXUW/DuHxIqxHo
GSx+8lSOH/w33laMQ/dW5Vv3ly49K27cncyLjpF9vZf45jRC40LV1eyzIBsciCpR
sgnHZwEu8H2djvqOne5QPcHdX+R5M6cMpvT/BP7x6G4t2L9T0wpe4TMScvCsH77Q
21Cyv4O+FqT3l/i7SU/V8c3PZ4BkgB8Zm5hUNTDvS+FwXv2lOrUD+Yeo1JJlbTyv
5D04bf2UaWI3vFCYuzOqim4Tl/bvmUNToMDzneWNnBKkPUJd5O6clJHvR0ugNclH
w5x4Zh+hfKUdNbSqk2TaBFgSiaAaQIkUFNl0P5UMQ8BrLhh8fEfBblD4OfntASnD
Yl9/PLYf5rfYLV+4CeT0NAwpAeqcLIrARl3QKjHRh7Kje/CTmF3hptadabY6+dhK
N3+dvn0+6m/2ezNxYk8zeKunEcPGqPf03B/tAx2zxS8KdhEgQTHd9xAJGKP06iHA
v2jGFSQJqabIrdX9FN8N9NlxOydmQx1PN7phMP9fyGk0k/ttEsevzO0NACmgiSa8
tmYPyjIx0Wp+Ke4lBr/BIN4fS0ybq2WdFd4UvnJifiL3XFLS7PKIzABHmXzUeyqV
7969M5c3MjZVll/DrrPVjdA5ybA1Y8FZH0mbZu+H3GGRxN+Bn9Gg+80LZfcTI2SJ
I2E/K6vJd9vnJ6OC8FYhZ5zkafiUwf54jY56dxFXoTuom72X7h208WKoWx0xKNT/
JOxPAHC0ElQB3V5rX/W4PBAIuoIPMEaNzkfXddthK+OZoT4iYovh1Z1QPDALfEmC
LJ49t+TYfnNe9XSSWrKI5/W0ivbJhS6sfKkuk34lNd6FhDzH3VS72mbJOVv3C0In
t1sbWbZY46C7TBNHFj/u3INF2dKuL6NofzbPxmalhhkwBoaXFOmnw6dcam57eGge
Dj1Q7UJxE1INfPa9cBGXx+ARlfb7ypL+5My3U8KnwJanBL+2vaeRuqJzRucWji8Q
DI5sX9yluFsab59+dVbhm0azndTBF2ZLLH2j+W+3xp5cVgk8r9KiRxFz+Mwda5g6
Nvtyp8mBBPoNgjMPl/jJ414SyhszGm6q6NP9xuhFQpr9iGmiCW2JYpm+u+XKkqb2
4vLjCZkEFKYBH4x7FPX0XruyMOxNtBAOBDsVJ9O6i8CYwk4tdPbaCMs3jrsaoFU/
wu/Sx9VdHWYWrlXTHJeQFxwC5XiAo5OMuYdipeEoPsIpt+znBo5E1jCsODXvH9jL
AtL9rzMWBMy/aUYtbY+z2/3ZybICXWjqWSCSsCO4aCfAf2GGe7UTzvZGrTTSz7I/
w4G4HDUx4dJE9PUfTY/1OLPSDRCffgY1kCpcUGXi+Nr54tMmuqB0yPfjV5cnu8LK
5BSNy41UfCF58/8RVuiP1L4ok4LWmDl2YmPTZEkWx8mz44gIygQ0qd0SbXn5dKQY
M8ZLMTgGAcjvPUPU/diOoDiYSFYIDbQUi0k2i59h7OFaeeFKLkMSEM/vUdEZ6ljZ
3s2yQygnOJL4yRc1BOHNagqwM6XR7z9H7Uq21VMsvWtu63tHE5ZPlZxOMQ+FjDaY
4izy6QnNZl8Q0jaN+lX7B8q2XhDOgXH5Zntf2i8Yn0sean1O2qxs78+aSY4NgQPZ
UfXg/NH/+8ozLChXRxsdW9bgxsPuUeAz6pKt+C7zZHYsw7lKxHbz3cuSgxI9Bw4G
pzRTQHwj1d2hxzj+6bXRVs2jj/tvo595seN3c2g9J4uNGi7LrqPSwEnT1jLCEKLo
PvuCL2nqJo0f6l5hio1NUvzBbZEyEpG0Vv5BAVEiKqbGyh6pJpsrjdx+2LHuTZDU
lUyslUXBQkiWna8cTaaY0h9cATlT854tfpewZ4fbXvd1+YqGqaS4+oYe37RZXk1Y
tnFYF8rlJGXlCeynRjwTgyLawavact59LSbFq14Lp5AlQD+O4MIyzy92SJNCaX2l
pwddkazdHDqu+xdaCd1IaGJxEKXELeUHj7qv03CWxoGThk6LQaexvrX9pbULS2eh
PRI91aLkO3KzsMSGZKZ9s7yd7JQHrgON2h86sRVe1qZQTS/YE1Iyngyo5dpSo4YJ
eNgiib/9k24Pj/mQcepQXgewVnXWiU1EDT1c8C2zu35wkycqY20l3RvTA9eKpELO
2kRfmX1lA+Z0RCL9dX4yEnkiCu88kOvLq3IqMPQyrz10RGYzWf+6iGr2XSr21Xhe
tMGTR67ZeKRyMorcxwrYhPq05SrBSyQrInv1CQQwXRGhsl7ExGFJ0UQeYV9JkHDf
ht43eJX9fCLv1dK0IW9WOjh0GoP7ebR6CTGyHQ2ohewpxvl8bNQLlsvP3elp+xYM
b3pLgyCl+/7bvEss73wNtGoE9EP5syhY6bqxPrzkQkfHUpOuymlW0JSwJB5SMu22
jjtpPN39/UF+b7LdBYsOSKUNoKzrR+hXVkKeHnE6zsXLkRo3+UsfjPAs2TskAB2g
v06Fi1MjrAJZt4DhFQCeraXcsD325J3KET1oOkbgxEUymeT7xdXkOnvQ+IcaXylg
Np5VnbzlI+gy+PXwSU+ZBgxw3Tt7D2E9EzU3D1/P4itF7WxDhLrX/vVxp/5UanCi
XnBLVE6u9bW5ZVLpfmpZkn760KSqj8Qmq+3Acs9e4x/LinZSXKsPgzNIo6eE+zYo
h9LF8mWjQbYsTT5/L9RV4nTq2z0pC+gvl9V6m/CqCzqs1c6EiEfvLGfnPWGRr66F
tmuE3nLPpA0bzDxfVyRR5lk7KLJHzL+Gl4MRwUBJRTmYBTinTNFQVqrgrj0ARpBv
el0WJOoVAWEm5z2M48ODnsqz4mVLaLaBbBQ+6k450jYO9DfPHbHQCaxokp593vi9
IrA/FM1tDsdDppmWW12cQv9JPwWx+/UxVkUV8IPSoyCRcVuuKARpJT2Rw+ZMEhVG
Ocdh/eT8i1X4Imw2l4PNpIkCDZ8R4wQ9/eqm9YD/sv3XGdkNfbADLhaEqM/UmhVX
4HqD8/RgXG1/ODZWdd+BnrimU1T/yo6K+A38pDtGENjvLh8T/Ph1pfjZAgVvoYIL
rwoM5bVdR2OvpyuIdkBFtXtARfUwpzJOi5/KKMcgejMLkteyX2EMFw1X3LKK4o6x
lnkrJ38oAj2bQIVPbXoTrHsB35fSoithxrIfcwju/ekCKwANg3kESgwvKh/VdN60
7X9zL7E0qMqqc1+oTmutzNYQinufLvDLLjXjuMIn0g87GhiQJL+ayE6TTAJ3hN0q
W5bgJIhzGw2+NlP7jFVzS1KsJaD2uAcmCskIqUmgp/HLTxkbHFOBvy3r8xL3+7lS
Z4oCLynOLMJMUp/YuNmMaVW5FODa0A4sVxsOu7uPY9zkIWyNDJdfykDWUpDf1QoR
DCRsQgTxPahOYW/IvD1G21vgNCOxd1l6GOh6T0WnmOSwFJelCiB56C9POQqWwoco
ICR+db3KHRgqS6RRE87now+hRYSs29izTTgE8rCpI1K5mwafhT34jQ0VnrWD4doE
g7MRFSru1Jay0GU7IwxIJMnnab0MwYVN7UtV7dzUY9mc/dAGzjZEADVOuD4u5ilJ
4rZGQ3DWtDBvUUWWTRmoLcrXful9NTF4u99fffGoeEzGBN5oAobPEokODrWTVE3y
QswRum7gV5jZR3lx7pqPwDMMiCx/dzx4fnJl7PB3E799EdS5OEnA634pxrLAGtDe
VeGHBLxRX5pxwRseyub1uTLzNudOJbJKHcs2wxH46Q5ynkWi7uVtTVTcgmiO8C1k
7Lf7PpDnrBdEwAvjfl4bi9vZHmoov0hsat0itQ93p7tcBXMBCBj55YXRHN/OV+F1
dQpmqQGo7Vf6yx4QZoZG4d5w+TRDxWkMuLxOADMPnKXwJVAEgHcJA0lYZQx3w9oT
gvDF4EPCIpoIX82mUs1hPmq54ksoQhO1srAfWQ1joH6K99WiGnIJpoNRlcSyLNMx
mPU52mTB79ehazamy54G8bPatzTRuARp848PKea96Ux9onhBr5tWhqtfWwPBBvN9
1EzBxBePZzlWgz9XaGU076E3LWtMpcacbq66b+L8g4N+BJqM/a99yhxeotpQLfIN
xEQMtp/aSNDp98S8OsgUkDVvYCwROq0+RPixHRy0cqiWd/CU9GWMN+82k0OwbFvH
8vVaj8RmlOwfWG2i0nSPH/ua3Q1KnqyTw0UadyXkshl7OSCGsS4BG0VyGII6RW8z
vT941yim5NwPs3TUWV7j6di0f+EbHG0wxiQ7ykkFQtiR5jyxQKs8M8fGo/xfOKlR
W1hCS741FO1cbb69uxfib354Zr1mRO6s3JqnaAvA+snqB5PatVm1SNQFSH9FjLN6
lMO0vDI8R6QwoONKEq2mWawt8spN3p6DbjnpQc/u3mTHp5ytnPtv1sSE5ZgeOzs+
TqNGD+27r3hVn2Y/PeQM1qZjbk6bSoCz5NimxfgjVQwnzfrxOAp1clILKbdyFsQA
V4+IQAj8kEzjWIXy7AzO1K6IF9T+U8gsw48yWzMyS0c9u8oVI7usV1ob5pwk5nzb
/4KmUpYZxTh97lFK8fLMe2i5XrqbP5A5l+Azcvv3CngzVVV7vq9cgUxvOt049ovs
/HlBnAJdhUQiKhZLPJqhvI6mWxwW8u2gyXABapnlhBjRBL9HMEva6r//hfMdsjDz
uga5w94PhorRt80PSe2F2iEJTCdSyfcx69fbeCuL/yXeLIot70BX4ZN4rLUlsWKY
Ig6tu2gaFSLeTdiXcG7u7qq++qBEZc6GihLz/pwrZ/y5ziP1G5X1tANo/AQXkBcS
3ENgwHG+V8B4uQzguCtG3kjYgDVhW00eMJfZFm5wSZHg8FipUUxOHJDUIA2Qpufj
eU18xPEvvn2tHgzoH8FGgyIptprGmDDroRQKGrRqpDCLcI9WFW9rtivtHqQIYQzq
B1tqNYUThozUK/+uTEpkRbADl1HANRv7TV5BNdz/sZ7ZhrsIW/PUQZ517tAwhjrh
BQ42qsuGldMq9qmvSXkC4/OXNGDPfx/oBLG9GloZynJWuLFCUc/UL8/dVAjTJYI8
TCkGAdYkjmfGeiog5k0SlNhxqdQMqUvGcFawQMRcf9i25W9MfKVsvGtkPd8Y1Mvp
T78HMQBefTbOX4AYVsyJ3Nx5tUpiAhwVweG7dbSnQDnz2ecxinJ2gijYcJdscjvs
DedwMoDS4zo3C+rzIec5jWrmu9Z+l64nz51b0/1j6JdRkxdY8bSPdYWcszepVg6a
JQrD5moFs+Vga7BpEjDYzZCOni1sWYlNRfWMOgx/joydo3kex/ZwA2r5Mhxjvf20
OsS5hZV0WSgaMYCL9YQLofmGroyhsG1I45/ZTt+ObYPmV7YpOL9qcvKbnExtZm81
aAopqiVz3AEHQsCW5+gNFbV4Jy9DpZypjPPilVF2slU6Q+SorytDq8CPzKJDKRMy
3F3/ps8RuuY6Okghz1N91IqMTmdEbWS9mHx/rynL1qc/Dz95P6OGhqLk1noilneX
C8COmQVWpPk+3B5I2ISorul14P+5DP8oFeQAojzGYYJg52OGcjsXegHJ0HZDOyrW
eoi7rfcZFGYpsPzUSlIiDriGHlb/QVNMZ9kNo/DTzkghx3X5a4BUkTpQN8Ts8ez4
4VERdFXU0mtF20WCNGk0sZJiEbYgJRK0ixEV0q+iLiI+3kwZHLwsZsLOpz+p8t2l
0mM0U5hwd3RiucmfAhZxHZ0362oXgA5na9riORSURAt1UPLl3vghfwGkCO/O/M7r
SZTo/WAo8sWU6dlHM/WfXtfV1a9pBCeskLAinZQbd6ubjSNpgjc7X3w+VaoI6tYg
B4bAbyqjsiSQFbxpJnBYNRTNsszXPUjeDzgQYW/Xoy/Ep5KDvyhhA6Df9NgGhFLY
bySCy9OF4lRrxR1avVMVyPzmL4SNz00H9SQaGzeDmE2bEYRw4qHLUk85WeJ1fqFf
q04gOQWTt9vSLGAG7u68m8QwMqlB7HHVbkc1AW2lug33g6tcbZ75KewOutrYy3q5
zpAJM8WtMjYUwxsy0bppke9Y/8D17jYYWbGLfX3PKuKxdx2wbBikxWdbSKlH+MW6
mClP/cl0Y0NUuRPRAoYc4pGREh15XdIE7heJ4SETznu0uARp7a9RrSUNAdDamxcJ
/WiKt1czJssrYA9VAm+lwbVh7TdT6MUeKKUFFMssJWL051r/EJKEuEVpJ7Uwf6V6
QiGEs8v504bvIsqykdWy4jL4NBx0xoQCRT9hE9zOzElbcnyW9UPojd9uzW90RzxV
aOZ1NKlKvgEd0V/VyBGlSygdD3GUlB0Eqei+T8fBDGKBarekDGTo9wKA+EeYW7+L
QdQXc+aMFpymANoOfQYThEX9rlwBtQnIbqOlvUDj9kdjlpOmwcqkDgCq8r3T0M3d
HZ2RhhISwErYZeJuG5JPrU7s49f4fJQPQ36oysKfhFBYXeNEJAcdkvht/Dg5Wn2S
aIFG/1ZjOnfzQTZl7Z2Zvq+5ny/B8eGzBOA2gQ8aEHTH9bVqYqMjHtfXA7Lcn7fW
f778HGHwRtNPXmQ+4CLgJJbC6rbkygiWUlllUm/kkuoTEAsO/qD3jeaQeLueR1qC
ZGLGzbiCUMuhHgUE5LzZyMsLsI5HSApl3wYn8irq/vJFVXqYFLuWbM37OkeqQSRW
90fZO8HEDuisi6Sdesap2tVagpDWG5R0ThRgvwpe5QtWR4rlEV/cyiPQE8f0LXh1
bPGZelxpyDa/LPBh0qIBz+fyJOYY1xKRSZ6P4xU/cwLBuh7LqkoMNJ73k3dA0lj2
l5bJXsNHvgnGbg8tP0ZWPKqxURPQFrrI/ZC3IZLc2KF2mCRs3ivgXJnAWqHpg39B
qgbbjH1VWEbY6+329txdtDAhiZHGD0fQGqwCl29tLDvVos/4IykG7CPhAISfVS0d
3cTZAtJbdv0ftIavtINgZ7w2bgV6aAXq3SPWLBpRaZGhJ44Kpsv9oBU2d39tkMge
JEtSBlGTlI8flI5RSqit1b4tSe7VrYsuZRWkKSPFSUbek9xihCqyArjjCVK/03f+
767dE6PuIVJIyn2Z3NJa9xN0kPiyvZ3mMUGdOKx8zts37Wo2FwdGnbiKPm2ChL0X
QgqyY/vkkqtZdjph4W6g1UlzRb9PglyazDcig2BxoY+69jBvWnoluvgkrTLgE2PU
WMAB6xYlgJu3XI53DFsJtsQKWDHxU4+m5gpVJKO08yeAY4RhsIwqCCTh9hD2us2X
wUdkkMaSUJntz+ufiLIuMQElCIKOoAtWbUVgMegk0l2wPatAo6B/GC0QlX6DBhKv
7zVNDkq6jKb0KJ75SQEXaM9FxHRjpu3AvXflQve46SIKODMPUWo60fST80YRzqiQ
ZIwpFWXP08zJ4wP/e+dwy1+49eaazDbyRhH7vrjrNflLzcGYWdXOC52s2/k+664d
aeTv916AU+2HSdl5J72pgOlj0EV15FW0zn5ikFQmlvzoW/wM/FKp36/nm45zTpJg
aIrvZKo+4sgHShhFshFSR5yE44dth2t/Z/MWptnZHfPoWk0TeCcylhPuY69qfFly
8vx2cDh+cYukAOxlN0LWbM+DaHXTRZXH4TSk16BGP62fgXrdPtzCwqt9VDpCprXT
2VGMjUoItp475v32Tt9/eLCqYPUu8y87MTP3hwWCnSNultryEOLwrZ+XFkHHFCeJ
hQZxWNA/xgOvYnD5T0ofId9PdFXComAoASwB0hirkaxGFndpZCvd9zZsLvbQa7wp
NByQQCsAeeJVvqipBnd8Zz5soNdqcrEPGPhMgfCF4ZuuW6/ruQ32XFaG7pSgh9gv
hAv+Yp/1IXsEgVNI1OO05ljaxsQiGPB3KMyVP/Dt+kfybtBTUdK8HMpwe3UIzMcF
AOfopkUwc4HViS0S1AvUpS/haP4eZ4J6VebWA8tt3/OBQ74VBoO2Sh44OfBUMN9q
M3tKXsTXCjvuFlnsFi7zteTEcBnn3yoHWZFcl3ehKM0R6OVFyycW468FN628OHgt
Hfc9DlLf88E6Fx+LuKzYkzsDf7y5x6caJ4XfCTP7028aiw4fgOE+WDtsKY30SPGq
1Wba47eE26YyPHwEn+jH8MEybMAwcDfrsmuYuREB7DlRc/q1Sdcg0XV3ivX7DPAB
4RQ/Ik1DQ38XRVaEVFDt+5pCR/AFKubr0ZhkqmDfkHERULLV5928/74mYX55v2Ag
J0d4Nkjixm5Ot6udQm/kBg4hvaGHf+JWbycHMGwUMbmnu93lKYLdggRIeyAggrJL
SHW1/+ZvmJNJm83pz1ZMsgKigx+gdz04CSwvCqPXJWNsT9feRJFOmv54pJw1e0gX
TBIyLjMBEa81pzd1TIk3OwOMLoc+7lnhYKMakA+cs09pfnTj2fbMFA3+uhxsBU+d
`protect END_PROTECTED
