`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hUJavEzAd/HmoFUwyocYnKKAkZ1j7yQDuKxzQXT7TJEddZim7qo2fncTolSol674
PfsLwVr1oQqyP3Uanq5Fc/8RySDt8Z8vxJ4T6f9Vg52NMLTjcOQ6RO/Ynn59bnCU
U0tnkoaOwIs7fCXqI/6LSZ1t/3Ly6VOagDLF8j3BnGC1gbAowORd7gSv8Uw4wTjx
vXmpU6ywQWEh4p27ra+4aNzXhazRbkcFm/M1Ud6COBmdgar/DKJ7Gt4yciEY62H2
8R8gpqwyT0/a1E0Jj91J3spWSCjWWOiIrQNtjMyyXW9dS6TxC/UBtbxTUq56e3wX
WC3cuC+qsQ1TmtGc9lHGRrWH2A1QakE63cvatBSFmd3jmWHdpyeK6rD/wHPl3mCs
dCFvZrssyXEWPFUEdqwh61PkTPhkuxLy+5woFv/fBWCXc+83gSH6cPy6y33oNKAr
kRwOlG87fPdxto8tWUPVlWOHO5c+RrJCkpxSXQTVPK2xQDsnlC39oNUdWZnxhbWJ
BcTgBxgadEfcb8c2LYHO9+FiSJ15Et7T/f0b65fRsV07GP09HiF6drw2ggCvT3Pl
elWCm3VJM+6JVDppPuQUcJWKz6/kUmtVzPWxkv2V+9R3xU+9LQ9btZjR+bF1V/NA
WGKJMfr1Mrtt8JQMC76ciLPjIL70v5WrH2gkqzOEc4acqkQzycthexjdvErFH4yI
rOCqvUjMysKzjamn+ym62whCZov8OkgR/hq1w72XetKkQGuV+3RqPLeJRecLMxAD
jMeRjNg2C7wp2tO7slcHg7kl/ZNTGZERuBjtPF/ns/B8zpiEaNKxzQ4RxJP4xK/B
41zdNbkyxD0mfe4SCmeMgeULgT6Pd/VZjGB3pMvWg6DzpRWRlcHb4bDYmkuh2Q9H
YBheECt481fYcLRRu7L0uWBWndgWRqa/aJkHVYEKhmD4BkycGFVVJIUMrV7g2TZW
PHtf1DvmoLKga/XIgAULrwQneppBu3yze5Iset4cq4OIDvIgSiYDlSA9dVeJeOUH
ilGddy4AyKwaYAYwRwvIgtBGLz6sPJLANgFmLQ2DT6MUMNyVjkNa9LgHZ6YaTxvu
z+XiSV+av/Elf9boYkKruqZsGZs1OpCuhspdFlpfys1TBcGtIfh8NjtKVkqtz1nW
mda3yrgIuWkn76u/2ELEWaP2M3DWCL9bhqezfVWO6X3CYuNNh5Yl+0zibw/bPfw7
9u+I7ptPQnQFs0u/89u1DYE4n/iISu9d/JjG2TtvBVsVlHZfHh1BNRdPjxnIyR46
EV+P2anHTGVt5UQMfq4uMs0KLIzpHgIv8Z5hWlv52X03Bj4/Ma4wqB/6qUo4O4mO
MmH0YZRUwPMNjtI19uzKSPhWAiUXunJBc7Ri2n7jav6R7jDNapVqU9+TgW9RXeG+
uWbDbBBGUC+0UNjifmAvP01p3QE3D4EP9fE6rPacWE1UYqwHKdTWlpIqgUoU6D4k
Glst5R3C8pPeVj1aZ1Rpt279WX/fvpzmUAod0CX/RQpv6rOj4u6ZbrE101IkxUIg
FutOkthKgmJoaV34yego/TSyNDqVP4poQoghZjXKbp3+7X2T2Mt4fd6COJ0XBUxr
pm/LJ+XhbTlCU76qNHCSKsEare7ObqGA9ByFNfWAdWXix8I5FXO3z8/xnlLqq3YN
vm2x1EPIgTNSyPNsvI5cc/EWVoY9lMv9dMKIxZZOq3ykmPpOGLXb1//2g2YpWeUR
8ElLH3RTjHItjsTeuRVmmpX37OwSQm7IPcYoG5Zs9IzrOUx4itvw1dXzEQZ4x5me
1e3g7Dj+4F/JyxsmXa2ZlEnKHxK97PPMcqHxAVsGV/Unpxsu2ZFUAPWiRjVx2Jb5
O1O42ZlT17V8UkWPyBNUiN7HQ9El5KAc9ULN19K1JuYYNWCiyYa+fvKCVzugDcdp
0/qb1NlWGuAgL3sDbdF2zuNvkHqeLKG8+tvc1AilgB7RKo0fQpKNb5GfgLNDIqvj
/BrYra+xHSgSjZjTKf4p+sdPXuYq7vvEXhifIG4UxBn2GYfuq1QaIMtxRX2jxedo
ubKy/vNYDFcHs6m1n2tlvnkFGBG54ukKavRTxCCIDYZ2dFw/Qo6j4QgYhui8cfGw
i8lKmPa2A3gkwKooLn3pQ+xAYoMW16+vTpOrQaqqvNh86YCSnAVocqWH5ubb+GHr
CX2XQWmMJYubBX5ecghdCLA4IT1XenROC/ehZOCZoO9c7Pc2sgvjofN4DwArHt5o
eINQUR00ZfkV7EggWxo4GMigYHLxObQbfRNXlrX8zrZv0dCCHXXsbjzeeGXgbpF8
vLizd2UUWnPFFgo4+caCYdbndLqWlBj3XpVv5FCgsd8s7f8qVud/7KDccaQaYRNN
gjH4sZrcEVn6gCOPDzM8mhMhWrUtTRe+IgRUJmc+BdttpLMNSeaRelV1qT1fAnfj
L/34xGVmDZ2KSyUqt7PFP3xIDSpMrPa5j2A/i+gXhOf8YLVGUBkX0/3c/xBKhFja
vm7BiO6Q/yHQlFIthjb/3oqNNnIvRhy5qa+3bcuFz2rePJM4ndgNEuX1DiUa+u5W
WQjFc2JM920ymujXVKvMBCvoVVlo684sHHe+RRiLwZswkZ59NKlEb/CegLiPV9KO
Oh1lXLC6crLWLh0czfYShmfz0ACY3+xlO8OvDJI+2Wv/xwzPI7FjEct+mxSjCV4a
pR2hu+RJesNuvT5FNhJt4BuxOAiTT9sZl360KMdQ064Wl4JulkOa8828QW5JV0Fp
+lrgCBCOCxqiqLEjjo66RMupKUZArWrPa7+1s1RvQmL8KrQgoviSPAuuSh19G+gb
MtuPNABGAZi4H0w5vjnmdsRToEQRY+kl+iyX6aVXb5DKwsAMZC5f76iXUNWYbnJD
8CVMwjO0hdMof3xb1t4zhCEfVV3sIPBZcPK4YZ5TbKCbhUbc84fLK5E8aTlInHKa
fe+hT4ls/Zajb/UwUe8NCqBoOg+uuyR1ea/quoRw6YzaPqabmiI0KcXc8Xmtnlw6
usPAXZV0134VuTQ7SicdE3R9ZasKlBD+IZI0Z2VR8Xgsh3VsAwmkYbUq+9e+IC+i
xPE50tnKHxBWPYrhbhwbz7AWg9A0QiTU5OL5HyoyIMs44ixgl/M+ZqBNl1dSWhqx
fQfXzaxlzIV53TsbIh918NE5wcqfyfTXlkY5gOElCDT3/9+XU48VlC/c5vVujq6v
OaLgcbLbvw5RsKyOBg5azt2S1X/7aQjEfn0MiKI2Xupfj6sZ6KKgzk3Oa6dVbX3s
c4yK+9kYK/oSz9yzZlb0PvPedIR2/abwwo4w68WD6h8M7hU+EfXc4OkwtTAbgwAh
pCLzRsvHo4RUx7VYX6uyGbbFfsty+kGAJbvFWAM4oo2wTcQomt54mEyrq4J6wJ2t
C/vrsXFckqPW5VlObY9ob/McPj/R7YjWA4ie93hANuQJQFRSHX1SnNYLhx90xMq4
DRmzZBYOv3njp9I2IwQw1Mcu5Mulxfe4GfpSt82DyyqZ4gUjoIPi8YLS3zx//+NM
+Ur+AacZionlK66HWRFMyR07UoMwp4OAU7N/GHFVO1Zqb9p602xah5a/UqXB0U1P
44IlGfn/upO44BAYucJiwTRV2MyZ4v+Qak8G0bPrDXtQDUwYTO6N0pMlq3AogIj8
HytMO9Z5OFjRPqFPpCJSqGZETaMkQsezZHYXP4hJT99+obNJkFihto/t9NxUI/bH
QcrJZfU2wxDDWcwFKTO8VW0bTig7gU2ZvGjbG1lLsaGZ+CgkPKeavAomwaYlZ55B
ViuHw6zHJfxr/SUs9Lw7FXuy1nxGaHeNmM5ZmbN761qoRRZu3JVwlj0bx9MMgaYP
/XutxXtGoOW9oT2eQEVm1l9ijmmXuBAaLpzKM68L1vPdSBy4s1jW28L3X1qQ08+3
/YRbppyXmEnmeH6d0ydCcbRImokNI6/mktLrZw0YBKk=
`protect END_PROTECTED
