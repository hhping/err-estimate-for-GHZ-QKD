`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OJtpoBDBw9WIggOASaTrHBSUzz0xtp6z6qQNAkEgu1XTrj1k58HWzzIjffsMzzHr
a+avfyAvMvzfpBvXAvlaiYvbgF7B90NMET2R1E86vptN12voWpSd+6o7z9Ke20co
QWYGlrOeTGX73OH3JwA1jnHLoxRI1FRjHSLkMxxiTi+JlvvxVRGO4RMNjmiJD/UT
WemAkbXs1ewoehAHOAFcLgR8kRt1ZBJqYWPYnvbbQ29kZvbAfXrlYz8+Bfk2W0lz
EHvhCufQw7S1R35yRq2XnQ7zEykXPLcyUCq/vbze4FE6UJ6Jky0KFJjwvOIhWI3L
4k1k5CuznkzDajDwEFp9R62IsCnA3Bz/+2ieknuJDyTVzhQBIiFYwtQoSLmo3ing
SEKPFwZjJZ1UEkz+S8KRZWabz4lgfgX45vVBM/CPGP8m0NIZh6rqKtQdNvOBgtQQ
eDCNozaJN5PMTQOXiQS1m+EL6+qmI9Nn/OpbyCrb8/uEVH1Okx4FtlqotziWdl/x
tk8MK+1LKmOP2O2FAGMdRLWJ0nZ8A0GXzagOlprsfoek5SGdvnJ+2Bhe8FBPDV/W
eIUcG2photq/L1uAoHVfPl+7loSzU365CFknYlyLTXeS7fBpbcePVq1aLmvNbuof
yVOpagImSyV3k4FFKDtpuIqQJGeIaADBlDdp1bdxKy55pGeCbNNc0Hwu1e++7hDu
S2ILy2p6ePQuOgny8c5SENAkCDiDrM9i4GM49FMzLKYsNqrXZiE5UQ1Sz67CVoN0
tu4QEfZ/dCBRRzxVnOkLTrUTnpN9KAi0TmOm14m0+I96ok/X1KhnJaSIdtPTfcSc
ZYZG6yufISSWtY6ZJ1jEBFgND/RsNS6my64p62k3BrZz00ys1EBbnTqVo2NOtCTn
8VFbFaGgFd7KC7VAVillr1UcaA6NtP3MZMNn5AW07aD9P6HJXDM0NCJJ4w4xZzes
f3R8gxSc+7hJtFohjQq/smuB5XUzvRUt6v1Soq9uWVOLfV5spuX+tIbo/HsEyPLx
RgJmKeJ7LNYprAHwACXeIJLNkUqTbBeq4ULeplTLoXVm5ZOL3R/V5SVFAx7ue+kN
ZXdJH/an60smCStI2/WC7s+m3HfIFHKWRFT/MPH938D5nO0i6vOg/MCXz6kTRDDH
1ZkWtFMaqDfsy6ZD+BThuHyqerxXQRtFa89jncNmkOxrCFvi+9kJjkiwL3xcTVGS
TAmx/dxu7MwQ30j8vIiXSzeWYpmlY04b5AjM3T2DW5hyj7kTymQgSE8IggtOlcNp
voVDXaU4Q8fUrnV7BjMDS0tJ1emIgPKkuoDC5dsdLgaj6ng+5RqTGo80FeCF3jB5
LxvBu6j6sDq9wVakSlydt3JBFTlT62x9yW9NbNc6lGIulCu5dO/WpBNkU18LvvxX
4/7XKK4xC5C+RDFFYOZs5Hb7nsZcBG3hsMpdFEbVeXhE+uPJe/fl/pcj5aNFOOnQ
7UGSVjEs/19n+UJesOD8eplm1vntvy2lrBiaYp9aUHP8CHW9M1qTq9tXtfSGEFvG
hNExlMFUnjW7q9Ds3/LltZv3zVi7+S9ng91JcTCDicBwliurAk2FAR3cC2uZw7/y
7xEGtp31cNkn2GALYbwv6V4L0TnE3yVPdY+bA+vqsUPoqaubVsrcFIw0EhsdGqd7
5EZuIF4EFL95ycLQqRzBURsC/Xjhf+WMAD6j8YapHnTcvzTse0Ly+LOcdds6+Owf
ouLf0q67i8Gb57FMei8FqMEURqGUI3EPbCbsEBqX4pgufk5bOcq1V53louSLuwmQ
DWaWkUIvRfGqMJJDWsiqT3QYoD+quKDPdTQX+9dLvK0s2UCbBIy66mXgS1SsPDbd
Eg+3ympCwc+7xUDTdmy/CMSlIhsPDlJGeQ7401xoTvgX6yT6pJ8WVzg5wcC6+U2e
URqa70sjT+DjF5qmilbpGv9SPrvgXF6c6z3yZ76ajNw+Rk9rNenoXno+36IQYa+4
KXKmFtb2SKK3DTG8TMJZ9ECXrBXFqRHQXbDUZhTUuPTbg40BXona2zN905LFcLUb
4/dxOwvt6647dDYARx2ubFHPYqmkyJni+sXDQcTlhaGHfZCfkvJOdWW+FqXY9rdH
gcRPPBGtQvl5VIlUXrYXyHvzDIQRM/s8CxDzdJ4CNIE1gEdtMh/u+ozq3XjvRwyq
DWci2lsnJt4r/gT403WmE8EkvcgwUN58mpFmWGrwaXfNdUSljOX1hDWL185EHPv/
D1fZw1327A3rZkdhsQOFX9/F27pThpXBXrLB2beGkn8Wu0cpAPYz41EgKcaQVUz/
5uqNP4bSURks0uCyvZvISrrrFVbKOy6Vd77eYktNaks25yOr39DGHSKtf+q34pzI
D285V6c5ND+Q4Cn2xxwGij74gcLEP0I7cHdnKbmsdzg388zUOSERulrwm7kO1p9I
svBbJx/AMTbMz0wR4uZRoZnnJ8IDpqa81X4aXHykhAuIDusZnLXqA6kQ0j0DZSXc
HPmdKCUZBzITu1yrUKnRe1cDPoes4LfJCsLlLNPyXFtJBsZt6axjkA+L8seahHlJ
IOxu5Fvfumar0SYV0snav692Y69KyGmyRDoCqUICeYOmOGBbkiERrMD4MKbEaF87
BJoYFXk2h7touN7HIW2B1KTZfzm36EcN4fe2VWGJDhl60dB1ZJPHyeghdJWmOdg9
1GyGH4XnISqwamJQnlMsANQy+Xuu2VLsPEk61zjUHfxvY6K5SxJIHxSAL3S8FSNm
/lgJrKwsgFBy7ETktGaxjwqU9HOcj8Lr7X7JPPoQ5UVIOMqkmnlm3IFhHoNI9ERT
PqoNYQKpQNU20yjFwTpakpwmlFqF8QxkXmIGGXcxBEGTeNF7f88jCuAmr8HfccdT
743BeGWCVF6t+xqJAFayrbynp2spfFGCg4wasAux1xfSoyQegfLlEszz70czC7ro
JeCUymgdVPWC/hZMCajWXF8Utb73nEG5zbbrxvNozhbd6SXGcV8cMRrVkuBzHEZ7
ox2Y0nSbtWHvbb6AZcegFWSo5fbEbAzho5ArqdOyYa4Bmwvg2LV0nlmrC1QDvgZa
0NpHknwGT8CftnzB/yYDF1JD8BufeWZVs02FA7TAxt85XoejV+S7KwimPnJnlwUQ
jdXUbn7tun1a9e7kjq9pM2twoHaphKamT7iANmwUfJadiPGG1Nb1TGiTpgEThcts
R299vnwI4Imkov9pFGhQDqBZiswI4zEqMSNJp6yv09LW4AqLqSckbij93OUYhHzi
DFVCDmKOJ6DioMOhbowMxJQ6sln9Xm7yLOZVzaLWWD5vneOqNlbZ/usdXJOao0SH
UyQqo80gcXdo+rSVTHPP/by5WRoZ1h6TEHoBNOppiKb4s02e4KKTd8EQLR1CRvb5
RJ46xFpHlcFZrWoT9lsgvVx6CbbFhHvdHtwlfNuVEygA+TFIYF6lFNp/2uwgLdVy
tBK49a+ZlhyV3UBfA0RjDqG2ZSMMX89fWBRzUiWfVxqV65iewNV4ZKAOekpSje61
FmbnZf6wBtlBl2260MMnqEDWJAwg50WVLF3z9qVd+W3aRMHB3GwmFk8yR69j/lxH
+SrPjF1qpDfQ5MkuzqMwWAh2tmppHzgwxHFXFdLb4uJMFzg6n3OwY/ThGxYhteAR
dmd3NnNvpqxp64z43qouom+tzhAf0+wXfbGTu4qKSDTZne/XHsu7yCaWxcA/O0pM
s7q02XLe4XaqESOVZfasZ6XdJMVr3mJbvuXK4Brym1gvN6/bcLVzO5urCglWCqqV
Ao9WccVbYsgSxhJb1KiUn7yFvg5N/TKQL/b0byF4EezJtADvm/qWA8DX1Xor0iJD
2hgPnw5L37kTX7TNmnC4759rtGjpsjwyweAp1FX+nX/WyvIU9IGZ56ZrUJCiA9vB
t5K9HR7zSErpGk8Su/qK1nFsevdtfraz7+w6BA/qqSWXIpxbouTPqxEbTGR4PY9t
cG1+p6bm6+XPHqcAxA8UvRmfwSZEfDaup3DHbQ2jt3p+eCKpTmBTjJirKrecSaTc
9c5XGxnCMctLpCUaFIoVYcF8iWhiXPd6+v85nYYT7/dCN2RQ38SMqqNhzj2E7uEK
4wJa4LlJojGgqXSc2APbrWQpOLk8QzdMZX0m5fpqZCg=
`protect END_PROTECTED
