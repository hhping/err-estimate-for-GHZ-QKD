`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bkeWKs3D1kBVvVLVdzDh9aLrMxzJvl+72/lGf160EVovrTxsOgwzw3O9iOGz1FCp
bYghFIg3gXb3ivrrsQUTVY5xYt8wlgEC3uP+kGQsYUMhA9dgajpeMNpbkgOyBR0h
/xXqgkLpXb1YoUCy6Mo6kCQ95e6QIH5Rc3vM3NaPzH5eq+tsHevRh+TkUtzpikvE
grc1SWF3gFPFZ0nA/xEqSFJPMLOpB0NPOX9sbW1uxNMVQpM1mJ7eA3v16qil3W0Q
39NwbuaXVDJpFqE3IcHpyBTVQ47MAvCcyIosW0CkxTJ59rNtCFezcMHYmktMPdcR
hmeKdkmddhCW0HUWGGUf+GVA9jJzLSVm/BttqB8BqitfLnn2/d2fa9sHrVxFqAUy
fT3ydz4GJQ5W5do2VWTyhAXrmscAl2ZYoLAi5sgFoslTdxs7hj6ZweA8QcGV489F
ANYMe3k5KP6MKzNCA7ucfF3fTsyuyU6wjMVoVccsdoUfut/eKYP8GCLUbE2YwZDu
morsJ2imtSjSDQbRI85uGglSMj/MaRBSYTkyophN3I5Guq7r7Jcpe8yNQqoMoTZ0
9/VdwyqCYzOAiqocgwmW7HH08IinLk4ZxWjUHW+8ieJlHB1PDGicVWaE4dahuXES
jG2mRwvyen+EFu11pjqhVObgejjYPLceBAsnc07NJOg=
`protect END_PROTECTED
