`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3fiwLP0Sj9XIvheA+43PwIw8xdrBn822ib7nIwwmStwvk2D7eCgKZf5NfowT/+J0
WY65fIbuumCs9dkQ/3+CK2svYjNmSMXAS18pnRpSOB4AEsuwSOE0/NuAVp/MLkv2
/uYonJ4JRPhKNdrieUqW+Ovibq5IEMD8uVbYBEcgLQDR66O8AsUc4wJN4u1moRSH
5x+6X1gLhgFqw68pXdMGvXKViY3/dHn7XyYIcNXl67DhmiC5kumDfwiyuwfnqRJO
rcdLjuHtNXpRteVSUhvK9Iof2s742Y2Psobk9AwtH7o9tIFqcysEeiywGY44YQoV
QMR7lwCg99nvxJdkI6M+1pVGMIs6dM29jAdz3OKynIqjjwrBCnhSQ25KZajMIpJd
iUGq7jm+s2FlqD1FLD8/u7ex5LjTmwOyh3EahEStgma38RCtUAFgdCeP5rA95uBA
tFDei2392f/VptdyLhFCw6q/aTxEjy88YsKuASn7wKPq53Iu0JRV0nEYpieKC85o
lOoLum9yu/S6PU6xu4Ke3dUuSaXOWMN+HauNXuSfGL03us1lsvXdxQs2/6qJ34vj
3bzCwcGESq6KYbN8KDI2JlilXKG8ViopKWYV3GOFnaBl0fnk/nXhZDuLoRaeJLMr
QcBDPVF29nITAKz63nNYGO2NQbGLnBfi4Bxl4kHbvc+pVguTLE7XotajOCEE4HbH
V47PE1ETf34qz3y+KmJoy9mPAHfFAkxfkzeDQmC6mfsaQyN5tsQ/CSgP7tqzz6hu
vmmZ40YqDQwEnzG/BFYNB72TfaUeDfwLUcEGiLILwliZFB+b2ux7tqjRRysGZqOM
f6Hax0EJeWgSGUzGy/svw18F96Y745thikx4azII2bIGxsOZE0P64L1Jr0k4ajMw
oUvLRhT7UqpTaz14+6c5wdou+sALOFTZqBUXyiQxr9OdGvrJeRrHjWYw+2jecaNE
Y7fwqp6opLxW/S7ZdCuaGyXTdxyynyKsBaCyYHSmAC/UAijgHzf4ixuV3Pn3xzrG
wnVJNNBF3pNt/W3ERvT5kk088F5O7e7HXTcWZrOr2IY94EYAxQ+lHeoQVxHd11X1
aCfZZB8lQ17EuJYw6hLtoFMMCr9lV8h1maB8LE394yrpd3+bIbEWp0j6YC/8B5qc
fXalCj5yYkx9Uv0nwVcc1UPEWwTSxT/ETXDxaQWydIM3FjhvWT1IDD3wx1sOPEJd
o2Gqp/0XSroUUXUrMTddyVzMkEqkNuQ00+GFVlLJv92KMvR1JG6PpeMcvbm45YEn
NOIvgfUrO7M3/i5PsEPD8YuhDq+imECMKkfEBcara6ElHL3B7vqvINsNa4u5x3li
7sJYpOzAlZUB8tB8xbX1kHbJefVv6oHR1HjrhMX47ARtNKLilCs8N7/gnNqAN2AI
3rLNCCAZ1R1sYOgZZW9WXNhcJ0wFRPqQ4kLMzGziQyFnkhav9V1443QiyLz5lqJb
AZEzCFKdeClWcjjxxG4I3w==
`protect END_PROTECTED
