`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4fQvusXbMsbiHQzcyM+CewirK7yi1Q0E1ogNilScS0qOrgHU7M+BBG8HcYPkUWbG
QgNDLL3SmyFFMwo1MUjQG35itktqjazYf4GOBrRwjCCS5jhqlFto60jxHMP6zYDK
POTC5m2b2/SN+JLGpnn6AwgYS0lXfK0om71KMpsxlAAUpWeSm0yypoGyXpLpKNbi
vzMhKpOgjABDyP7vU9hZg+zdVJIeiPMBI1TX61JEeQPcHjNGZbky3XPinN1wlBbr
MwkAShNLUFqGbsJ64R+g8zaiVQt1N1OW9HxZe4Ryd6SppNiqJFoqZ+d9VxllsO9b
Mib+txNU2xzEiYgDN4EzT/2Z4qeAxne7STKdZhAS6wTWzqbrugwloNb8qpPhRGHM
gIqtN0+VgL6mtp+/dnm2B2rP62ozBsbYABhqOV6XM2lTH0W41OLl+wE6GzsIdG6y
kiYUumRbXSs4e2ggeDCn4hodXBUYdLX6xG0V/l2rhBJNVoKhkrz2VBw0tGiNdym/
hGqyS6WvisMQWj5WDKV1S7tAz9wg8w0ATJ/3f9PEAAtf3kgSyhdH6p+xVK6+I+SV
8vpmCqv/IVOutDvcE52blEmVIf3zE4fKD5r2OEaeKfIBnu5yd87s5a3JmCBNstT+
QCZTswB7avjHufT2098csPboiiuX0F9/tVC5IWI/WZ/iGTZAfpY6p53Px6MURi9q
fohSdzyJ+GDmVTSGNP8z2Jx2VUda7UQTJfxJXEy2TdAJcksJIS3BNyPyMrAM5wB1
kkIvt7obLWlHKpNMGFBAeeRs/KbtDgijzzysu7pNbWOVAKnEhnde9q3IzXdJFc/N
rX/SXbJmgnBnIcM8UQJ7+XUNj9lb8Yg85G1+uKuGFWY=
`protect END_PROTECTED
