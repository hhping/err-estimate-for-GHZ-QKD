`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UaWnv1uhlErqHUhpXJEUxjtQwAOrJJxV6FeMupBkMel97uje7M3xFI/1QiqtxZ+j
mmkdD3+xcKtnlGQwRuXjn2VcE8HICtlDc57Vd283c7j3Rj02Ng0i+I+F4up+j93T
sWsd/CUkirDRpMSItH1zTr/HszIBp291mXz1w91oztWx5KBebXeyexJjMQ3p0bfK
I4mcxF2fb7nYR2GxmLMaHnPIubqmtRDZON5HJQY06HC5Gtm5W0Re8grgGYtP5X9Y
Y/CXJLxGAXkLnysq+p7Hq0ypyvoZtFLXMAgKW4UgVeGdipFX0u/m5o7txmuV9gU9
jtKO+mr9gHbBhqceVSGXh+2OOlVzxcjPmOH+qGffae+w9p0u72RgbsZ/PenjZYy/
DJ8cFWJjYbvnJpK2Yez+m8e8VvVgklBFSqtaILUixfoQAAWlqn/mP9XaCEsKSNO+
`protect END_PROTECTED
