`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Os8iygAITVQbpFbqPySpB6Genwm/BjPWOVM2rPQ+KnFTng9diqWz6Yszol097hSZ
Gdxv1oG0S16usi++SwQnC7YC19OsaT1cQ9wcEaDgVMMLjg/c6ereR5sh2XowZYca
fNS+hP/xJGmeoR6Mu33NVDypubHskFoLYVldwLlmk4wSImyZW/Mq5TZxJ5v7+rDc
17gLmrJe20INBjSIxS08chFUCmWtf1954JH2TrWQY2Mo+eKnBXXXCyedRvJny9tS
PTA0Zv2qtoiQgL+ZHBd4ENex6JeOyEgumCxgyrBJXPoiIUVZ/z+vA0fJdH+NFKlU
u2ifdQRy7MK8g1HPLsjTjlB6bArCDHgfY42+RHttipCRMdTJjJEarANl1xyCiRH6
IjVctOO/o1TVwafo3LVDUMCKNzoMHacirPfA9JRwYZkAHP4ooLX55W92MJTOLXt8
fwLJ5Dng1m1Bympr8of6sNFmzTCBTQQoyBLp/kG4VsDniDILdbA1k/gOD3DbU6GA
8UOTDkCart8owzqoszruCaQe4NMTdSlVXzkFMYfh/MkckX8p5Sa5vNBtHlgNS3VT
81wMnuQ/mMYIcgDb6msUX9sOfu69lg0svSEEKa5WB8AP6wxeuNwEdLfXXW/tPgnh
n9dwnH9HLNWZx1pPmJOaRGZlGCfrcpyeUJ5mulYV3Y2W1gEjgntFIK3OQ+LvyhEX
jjixAdk4xcRKaOrhd52uLHzD8Zw8ed/abruAFeTKIpR5slIZMtZO3R7Z4kgtvxZN
ZYVQ/luHyeU9uD4/vRHsZVFep1qjCwqJ/qba7mvc4jZvJDGiORRupn6O2hkVSAKw
Lp1izM37cOZbEqEjTF2ts+0bDFPjXOxdP4xfSIyelzPfIzoDtwBbD8ZGG132VgQ3
wK6jgcS20ahIYvWJPahz1A0gfclQ3nwS0S6IX9iXEi3vqPT7tfRX4Lk4VI/rlCEt
twl+3XV3zxj70YGMQ5fOZRnr/RwekooMLR4qm2SM50BsUDt9MFTy4q4mPDcGrfmg
JHv+kQhiLvepAnknxCp6Kv95hczizrX7mm70fIi+oabr4e2Z65F+h+UWBqFippiG
XHWMgIZSahOTbAH2wi2BoHji3PabM1awwUpdJIiedVWZBDg3ISxYY4O2deCeaBRq
0hLcF6YZRsgLB9bJShyA50xWtl9IhltVM34x88O4O4++FB/eDe8qHx/aGXFEdJcC
mqjNxFirrXeRaHaroF3QAt3Jti1KdwhXro6YPqyoV5UmxPEriO+X8NCNh6un5C3L
UnqfrU3aj5lvNdfrhfC5e5zOIvd2/fxOY/pCMpp0iHqWyPcx2qBFMebOG0IUJLee
54lAbb1SfxFygsRplgIazgBM4gqPbXvUXTGEXYCWml3ukrqYTtYhYJUSvUcVq5wl
iJDhSh2BSaeHWXoskDa9o+iahuQjD5IvUUpOL8tUjalKpmbN6E8BdYsspz+IhZTZ
860uHA5XKOyNVUyvBACDx1vWxoCd8tpf3aNHnTxXfY1Flo66v+whBK5zimZw1+Lv
HWJtVQGUBZiZaM3DL8tA6FgakHPKIgLWA+7TIDkqhIhrioprWJ+UJLGBFDM1/EzY
qtwqHCfclov9MvQBZMcD5EeJqXECq7jo2/me1xwAQRd/QMREvROIsXndbraQaVCC
u6TOmYm/wQrpcS+Od/CFjPsZsklda32ci2nTyawqrsW64mpXo6+N9gWc1i+J8seg
DKUXeNnygPozuvx6G6+59YtXEIIp+YMRoUlfXPcrpKcGFhl77+nWdISmmqSoEW42
inn/T+d5PwbUzMk1mECd3RJfRQQIgsnDTCT3t5a051kRLpt+7pp/ULKYmyF475KV
cBXu/Is783yQxuHU1gzAteejgJFyBgbDgVKu7vNFcB+4dzAXABAWgxo4rC3TB1u8
9fLOSusAamZwfGf56k/KM4OksWwfpecFKInOx7fxoexaNxavT+8ptCpsLXik+kg0
XVI3LDy4qLr7rRMLS/E1nWKyuU5NMt0nwSD+wNPGOogYrZb88iOIuUewB5LF7WzT
FdBciyCTKX+rZgd6hyEGbZReZeUtptqtL599KXt5j5PxcjpaaSouHPh1I81g3r80
LiRQZXLyZjF7c6bvEd7+faQyrP6zgupMjjQPDHPq7DCa6sbzRKDkPLxY3uy0DBIh
zJbW0MKCfGwl9ZWqkWXrJrQk28k685NuhVT70Sd6dMClfh8FOEYHT//Txqhwcezw
G9oGhulaLUjfSyTpOlpz9tR/euJ54xKidKpzy8ZJ8yOz83szatdTBkLvQ3WTw9xm
s7HFbN4pv6M/+6kF6yt0MLaZAtn6Q1ggKaH+p4mvtyHH8+IQJHsE92mbu53cakr+
knQjRoBqA2sZFMUKfB/FrFXkUck7TfWNvArjrayqPVGLp8hEvqXBYwLP9yf6LlmN
A/T+i+OyTLhA4g9dJCNmtpLK8pI+IKUnM4imr4CZ4hCNd7o6smCTz2reuO8TAlDJ
Cw5PhNbzcAOy8h0Nz0O0Vw0Nsf+lrhMWLqT/rYFly6w7tQtUy2yQ286s1lKE636c
P4TCXPIxg6weOaRpB/SnXTOx0sWbIfXh9qfj/VuEJeFdOApluBINDk+yQ6ki8PaZ
8ea/eEz2bCnCBL8D3WI1D/YfqWMwvr7JWYfebzMW4j34WQFK8CTotK0BDCERkQdG
TJwZZDbG3CvrbQ6STJyozMtKdIqxviSFPRKndVGLMLQqlVOR4dnPmHvUfkOMS37t
kYrWGSuZ1x8aHbDmHM2KOoFqYDOWvgdKBxFv4raimGblAgQGG9u4snZNYbbzvBUb
USyVhD0RN9WVa7qGa0eJmpwQJH50EHt9a2jr9c4dcT9PGRQyppxyDxSfHzrjrC+7
ndP0XG8ZST3AsOs15M7lTE8CuLcCmeqhRWrTqA37KoPXo1L2XYX1AnoVBjNJ1izF
ZRNs84GLAn2AuaAXqjawYVNLMEpNkhMFwEKOxZf8AMA7/SMsXKTiPfBYr6v8M5rb
t5SI3s5BrybbUFGodEFPGREoiT6Gh0BLRG/8abgNbJ4TGIsHRPX1t6qcCzpHaWms
sJ0oK0G57N49twegCFR7QO4fp1YWEyVwbeW6GCGuihS+0qoajyRbMm19pBw0L+LG
rOYVDGliafXwibtjQBpjK+ywUoE4BjeN5dQXaMuZ/Rfy3uZzQukAqeeey6Nj9P9C
m36VthOr4SUFGI/5OTY6ZZG5yGCFR+ADjeGah/uQdpgOT1QtqZI39Aase4tGJd3+
s9hgPqU40lgd5Ez0bmItJc2EHOsOEp8KWj7bQyharJRS8+sbqaUHMJeBLy/Hvo0V
vonhau9hz/Z+j9o5n4wjwaql57QXNrUm881/l8v9PhR9UsvhxPh3gaDdfULwSTlS
wpI7gSyHpq+i1RSjIFb79qs3cx8dyPkut6oxabOofn4um9xXzXBTMIGHHIr32sTJ
Ycno9ifWMRd7NtCpLCpcnkKBRHBp6jYGH9kxmG8sZCbTniw1GY5dNpRuTCvkqIEW
MJfRxAyLYzQX9oIVAizYOFXCJ/2ODY92Em5eutz+7frlrjveQzKHsky3murtuJPg
EuzDIvn1ks9LtJ23CKYMvyr9qgirvQX8WYKRto1CYyqRpZ05HnEKn7LGevGfiUt/
Y/yBfyhNXtqGloequYwtxW/O3k8TT1vBPNjvev9QPrQO3H2XtafpxQZQ6r8PXsFh
zozMfYLpWLMQepaV3EE8OUvF/OClCHaLhUHA6JnczIDEXBHwsrtQGhFL75dSTd0k
brlafVRJcqJgpCVY8RNYyRzPQwRH5uYMQkBcGHy3WyV9yUMktOiYBtgesKLoscj3
VtehJTZD/0RBAkj01k9EG+qxYIZRjtfC4igNOTKgD83naGPLNb3eFcvzUIgBe1vH
QwjVS2UNkCYM/YXChS4zIt8wiNURndkoKB5jFF7K/qUjiSZgOxfrb7WuaUkICE4p
DOn5HiuzbZTfzbwYNv9SuEP3JqgyHuktBOXPilAwf7qqA54XxWw9isgrg4KnE7Kx
vDcgCtL+MK7ga1D7ElZ/0JSQ4a81AxTDzvznTenhQuqnJ/Y3hiKxXUGcKHHElwcJ
tTxw5pmZa9iEEm9JvdhTM0BbEuAGU4mzv8bRwgxMeUYGjmyrTJrBp115L7nK7I1n
HVN1bWZ62uRrO/SEmb1xfk6bPi7CvDKkEsWElI9+nAE9rkZ8RBuMdbcJW0Je2YSb
4+FWGx1MzUKBg5NS9cOlyGv3eVTHD3HVCwVw10l0qahQxdmMQ9DfFqKYD7peZd7G
HNT+HlYAqWCGNy+FF7+HQrdRzyOwhEOEzuN8sX5pxezWBJXkrUHMXDhWn37XYmgg
ml8JwrN43TDO8JZ0f25w1beutDhs7rBC0n0uU9rfyWmyiOF0fGqNEiCqwwgy3CTO
UD9x28heLTBbSFLxt4XvEVa6DkEOQz6LDG1cWwRtyC2h+tG0W99P87R4RSUPb4jo
m5YkGJ0HfQajNsy2y8++G0RMQYC4d1NQSf991t/8ZI7lyb6Ovd/n0hI9Pl84Fe9q
q+QnUmxsGcvk3iybn9wx+XzYaUZXdXWoa525m0FnFxsGm7zRHoGWjsfA6qfu5XoI
c+QuyCs254KeUocFr8iUiC6xefzxYzUe6GG7grp3xI+OiK+JZI0IHsILZPm/hFIj
oJ70SWn6G42YWJrbsVha2kkCOGwxVviG+cvwYIA8YUZY+f/joXoN29ryM9g0mzFg
oKLh1ULRu/iRiwMuxLRL8aZ5fdGPpimc5gcpH3bY/arnNqoA+9+fHpfSGjXKJmZ1
X31ynCDp2kyGyP+tXmx9B0rtlUedOc26C16eGq/yKfeYzgL51++DdG0SP7dQ6Isz
KJkYr12V+fzdYavsjOfWvJ+aeHkw9KV5qE9fjibZMF/znvKSSIwliCJbAwQ0ndB/
krMaRw1643/4JuQJm9OrfCNkNMmowgH39eyFFhL6BsRgdZ/KB5z8ie8lnjEWp4JF
0TRhUc7xlfJxKUYQ2zCiHfFJRuFmASfwC+omK1PAY6PY0b7om1uGD4F5EEQd0pyc
7KtWH5xnspmu+ZIPgwyISYTCRPaSRRph3LOqZs48aQCOhKc8HiHCVQiVKGE8z9Tj
71t+9U6ys+PsztCd/DK0YtqtXoKR+AAT0Wsw6u6eFN0WAKQJoO2DrGu0JQNYS7U0
rJxMxwJs/cXem0JWQRlRAt+BfKHCUQJyO7h7nP5keW/d/yjIII+uZ0bn3NKPaTSL
jijuQ6Fjb3HGxWwcxGn49LyowXcVeCRTH7gbV2oUZyfnvK0x/DPxPK3PcaE/v3iW
nl5/90zkzZANu4Mm62fFue7FAFQsGDS4IADb8fPFAhkC/8m9N90R5MVRtUD063+S
1IVmisx/1o5zBhX5itFappiQ2AgY3RDrh6iSfc1sUxddjYj2KKPI6KKW4bwujuGG
bkO6WlVnSgjeUN6bzxRzGTe1DptRwPc0CvmoHA7iCxL5TMkPd30oKkLuJ3tfAzWL
ht4PbCIeQ1WutysGM3FpIyPpmaUaY0HM2YnuXyTXBHX0DB5oMOe4qsetvBEu4gGY
RK0BfBM9xO44vEooHe0iXHD7pJFBrCKGMh6OecLcan8LDJ4Uv+O7RaqA6mprFhmq
F+uhG1oyIzpdj8VfEjRHFRmlfTiUCGhEpxicp1hWtDocYAv+BYqAL+RxCz1FYvwW
E812YpCUjUKezRgAWwylOjcHPK4bFkzNiMZgpVKzNKRLpROwQZWHjF7Xq04gQDo2
L8vKFpwi9A81Mwc1wb5hwp08pHxTY2U+gLf5XpMF5xY2fSjAW5UHoa4X8FBCLWU4
5LAeczsIFrFDzwQdliiQq0RY8wmnLTriGzzzDxlRNyNRF0wlPhWTaU/4EOmpqqBc
+DZkHMEn9OzPtOjHDoXKS7IsDM6npTjiGJUJFaNJYTnFQ0XNs5/MM7wtTPXJQjQR
vvin0Tubz6WvwhDFhqldpxYRGTiHpvF6MYLSe1ntzey3tFJzjdspI3GNsfjjd0Yv
LeodUwFKZTFGtATiL8KiGT9JM4g4e6K1SE/eXoePk9f9ZLEuIDfucGNlvLEmrXpK
jGgJTitShTc7YTlMIsqt4GlvBm561rL1a3Msb2FLIm6jabgHZ7kCqjgq52noGoxF
c/QCeek6e8HNkdCWVR5wuSeRICqYDJU3rx6f2/F8X7APHfgchsAPUAMTgoXhz9Ly
mAk/jToFyuo/Tr0m45IkZ/vumTYo3s20IbFnA4NAV1QryVuqWsT8r5sRHAjJxJ+1
vTTcvhQCUW4gXrqdUVoMgmmknPAqzWJEIbPUeUF7fUA4ccZS/m29XJV6HHw+oCto
bO92qSxPG+F0emwjZxDSKWThOz5dINKhdZc4lrLSnzCjypUXGvKDzZDT0KfkiIlc
hV9B06eQeeThU617c//PEID+R+bScFCmvjekiLYpQ0e58Fy6jZq+xlaMAAP4USoz
HwbkYaoptvF/9EuiqbNzxHkhFuobVYC9YFGYNRH/APEVodPMg4dO3UdWo/9GmQHM
ajRn5XwkN6ZnNLW3Mx2AsoyVmxyZ7x2x0800nawJorUN8+V5tQMwNkDBzrsZNI9i
42iNSX5tpkBvxPxO2qdzegiuYQAAVIdD8wPFWTBtjzBCPw3+ymzjnFe+OJiE+485
6nM8ts8u4C9JrKY0RiJWp3IOrDZfFN5kjaR+4s2Jfy3tbLz5RcQAQXzePCjOs4GT
OCRACqM4CE5cSN6KOyPqz6FUazzTlAVVG4TqbdxNeQ/iqzooLoGh3R1Ur3LzWQC+
y50bVgc1csyzS7LZhr9K8HuSgmqJ8gt42hITVVdQD0NcAL4gNZ7UfPIjySixY74e
E0nbn+xuRK63+oFrUd/b7QnIUR7jiWN1MM7sjIkWxCf1sJHYVQd6kOktwx6zG7Gv
KOp6nFcjgcU2KxqfjH456ax2yzLL9yvYJrHWQHLT5n91QXWqL40zhtlIjolt8iCi
CztuaGvp1LhmX1pD7ZpJYrqIUlWVP3rZ8Y289HqDh1h+eo51zwjeU7sUGa6v4bu6
ZWFF36I4REscqzq03nZJ04LPFPzGrvIqmibbHGI6/WrGFRFepgpnzj/do2AR7u1N
wEnbaDZNxLnhlsRXAMR1hbOVWST5b8X9oibuemjgmSMBvqxuL0PNj9A2AHn7GBLe
Sywt14yxE3fEwRK04uaKL5p2+IK+nIDIULdwPJT9oJJ0ajTnpRFDJIZiBO6po+OO
scxrKCY8cSYGSN14F8UviWFEDh0AHlj1Gd9bqWW/LWMLPByCqBm+NkEvBiMBo7He
UsmQrlNFP9ePp4FjQAHGUpY7ATnF9wsgkP310/WIhv51LM6HNRFWX/818uzB+oKL
K/HRtE2eBvSY9Yq0M5vIO53Digmzkz9YKkN/swmPPxIRUEsNbJ0IJUwXxYpSdbL2
DkAEke2Kjt8tOp30rXmZ4s4cXgBxXUekVpFwdi9BZrEK+irVDR8sYf2tXMirQdAd
LCa/32A1ohCAjK00mjnuVaK6nrQdJOyRRrj87iZUKCjnQFGdmD1WsH6J/jgxmETG
RkgNxmNPS2QsEuqTwcQ5U6L69xRz1JopMnAz35jB05D9b+3j1rI7IvuK4BB0nfGV
3WmBbQmWq09YcPOu1Ua4ciMzFQc5Eiz8zSDgkSVw+wzgN5FRZHiY8qhVecbxSiqs
LdKqIhUhub/cKcoPaX6o3pibzW9nvIE4V8mVt8dYBrCkHoX/NEltdBjzkiMFomcO
P0zFRLIwFRyq2XYJ58EmWdDRwdWZkOrPs7zLNKXBDlgI+sx+lSJFwCIKqagHxbuq
kudmXEhI0mOgGI/5CiB5sCX50BOOjsydTzpPC2LrZlU1+/SACc3YRyZsYmVSD51c
6gTMUBmbENT5mSpLI0Ve9fabJNvEO4cSpvH5/F2gdn08ZSA6QTjVGBKj/YMNF8UU
IcRgw5egZFiEN3dntRqEZHq7uhujeBjRbmlYTx67klTKRT03avlMBhpmRjaD33rb
ogyxtjChXZI5TpWSdY7rdk0UzEpxSC9btx8jp9+O08GIDSvmQEPYtYORjHhzV6YU
N7OnMFeH7/TJPpeX6/H0KKkHSk8+Ki3ESswWhL/hzaffjzcVR69hxIxwagRpcmXd
3etM6pfwVp3XBpXqR7MoZ1pCP36KDFLDf/jOoDUt/xWrDxFn4Wz31t6mCiQS5sZ0
Wg2XG0Mk50K97FYkQlmpwQ6brbdsQsc2QQ1jy8yrNGt8xljg3M+Pdkjc/FzaivAN
l6/ivDbaWxSE0FZi55Q4TwrVyTe+v6mM4PCgim4MDha8gSBZMftQUhY3MUSYzQZu
Tfu34LKdWMQ2anfYWAprawYguHANjlaPgOYq/LZBdUhvxtGTJMFjpIEVj10S19Fc
fkXQRnpvfjguEWKAN7S76CZIVNU56GEhNR8KxsLDnVRFGCu5EbK/jEejuvybd9Yb
kQdvDsJXA2E4QLLbJCKJSSrdPFwdqTSYml2CuIcrw+dVdq+MOQEU8ekdAlyw+Xs8
FexyOaFI36r3j1RkyJh3sOoEhkLbv2xARKoTCoo818RuZ8iY8tV6x9yA83bTbJoW
4iTfuXPSExMpA8TIVmuXQgTG86LDkJsVA41d98YHhw/J+EKIPkbvGKp0Pnj3NTh7
Wj8hHyVBHg5cowGLzpbzMhgKALTTzrbF0m4df1SFtsh1eC1vjF7RWh83IRLlvVHf
m45pUupePLAaKCVV+MCDGx5u/j7SvHR6vbjcnN061+KuvguCmzynbc7nL0Re5kYw
ep+nJJ5M94LCSMnB4xEg75Sim2IKzV9AyA4QvCDREFYygsuV3b5oWq7U3cUlwA5+
MKD3FekUcks4GCWoI1bubBV2J1ly/FcsrpRNfWTdAJccmIKfR2fA0lNPuwDleaHQ
T0cRhJwbMW6gMQd7tMut21yVvxaTT3+41As80VPLfnkoYvwH0U5gsRzym3ywtEdB
LUTVFcT74ZqCBUnuR47IigIVxpLQiUCYrYR0h5Gtkn1pPm0imSzQs4TBG2CmGvfn
jXHyXxXkx3eQTZetl3Q6K0sDcN2zHmDG4Qo5kQx0t8UdpfrZYW/shgGU276mQu7+
gSEt7Vw1eJp/Owdi5Xono9h6ZqVJeJ2uRtQxnh0LTV3QpsLcboMTEslhr9WEd7mS
ui6d62Zor9oM7O8nHftze6mV9Xlvzvnye/Hbvy/Rq7UhAXPh+e6Ava0CCc6bb27s
U0Uy44/pY4aJIcAT1m9hNDDArB1nU6CnQPnJfjje2veQK/EZKOhe+U+melLz0DWu
Pd+Pcu4p6bOpAI5Rd63sUHH0xMq4V+OKMVafKj9sKR+FUlaqQfdcg+gXW429vNVC
4+TQXSWH/jNSSAMUtHTzA22d7wIZ+LcxhwAJBEmVsORMh0rg7/E/hE5LZ1DI4VyP
xutD5ALm0XpeTNKb+AXIjx4LDCqXuX8CKGTeZqmD7N3eZhxd+8vZduOvMhD7t5BL
YF3lSkQjkQzVFM8Q6mjii9b/1aozPSSBKZRBTc7BcQ0DJXxahBbXnY5XU+JY6uiH
7j8CRSfz7u9aTI3DoP/5wFATtVnvvOUeBIFgZuuQ/19svHAb+sLqDOgp4UHChdLh
kam41j7IsbvcT7OlqW3g9gkoimrvqVyLr/QREisOxtZOlfkIehSAWk4lNQxs8CTP
F9kQV7qU3bdOFtXX0FjEcQ5uBMPC3n51DV5j6zb5pDCeWTTuSBQZxZ0/y2V7YaYc
So6o8qVnMjMIm6pTdiFWjhRNUAcQjp03RQjuYwYrn62xauUidArq8/dJSP++DX/E
/YR3fGzHTwjNu6ghwfAB+qZlAr+dFTFSDZ3mMZQkRWahcrumuWnGPz9oGWAEnABX
RYU+2Ob/7/E7CUB4sYKBj+P1je7ntH1pvUguVJKeB/u2e3EWIFjuF2U5EiOn7yqq
PrVMngZ0AVQ1ySldJPpOBolYQrAAhPmbLSAEf8Dgd12M3u1+WEPMJPi3xXUopTIv
Y4fMVgAv/No4CKHLXYtSeAaW+WDYkMj/1w5TPmcqCo2jz1DvgKAAJ23UCpJL1pHr
CbQtIqONDT0nfHhNd/AF/atXggZT05gNDLskcR0qCoNtkZRDoSOexuRlbh2BXCKM
1mjSTivBoj8jVhIhCch8KTMm0mWu5+6YwlMM2TalM6Ph84oH9gY2wcno9zUJmrZD
ExSmj6v4C6WCiKJu1BROecb7gu8MTR6Ob8ldvMAMx6CiojiJ+G5jd18kRqpTu55F
54Ftp8bNh400zBGIZEdk/ut/SizHel4qAbLJ3JxMosaepA/QrU5ONpOC49aHNMEH
YPzdDeJzZRrDIiWN3L+gXa4E3gEv7g2ziSsrglEsG+Z0Q3qFDXG6o+EqthOMltWK
ums8DuzMS+YIGyrg5mfogBPs/qOjW05/ifL6i8MINHP4nQwmFeSCf9b7+HzMoEE3
JUPBztuK5bDJ5ucfLGw0smTaI1jNI2EgDt4XZ6PblImm09cmxV2O49Tb10k9TwvK
MZFQ+GH/Z0sW29u6uQCOL0nJbLL5fUVwB2oDQ/ne+U6VOLMFDJfz6KD+5F/EkHtC
zz2ofP3gIlb3eB7Dwzar0KVbf3XyMwrldQbc9+WQ/K9TSRKU/bV2awvaVevM4XdC
wYz5uVh2k5tl8SG87H0VW7nVpPpmykNUZtkeLSjnejuMrqf+xro4vyNEfMzhjQ/t
+bihk1C3mYF2eKrkuL1XYti8caMJz2tFNJODd2iMxVNJwyUynPxJ/o0KKE82uW9H
VX1TaX0YfJcMBuYswEsp84QqapoREGkfFsSTzdUuCThHx1G3XXPD6opoeEL0VZpL
0btgzrPvqQo6klBelB/y8OfR0i83DHlkTECF8igmlJDzCkUmPxH8lISnFLaDC6n4
lmMlixgY9GapL4wqTpM6cas1Gd4khO89vGnmdnHaeUfGHev3C46yrK6lOCldfFCs
0dHGVPos3v0Q0Te9BkxeZCz1OoQv1U4jUFDOAYpaJ6PAHJSXAsdlnOnSKPUwzudA
iPT9eUtwv52K4gBMlzbzL34tZe5u1EF+xnxqsG9OSI9eyw7/K61OGWhGMTK31mLN
UXJLRqiWH97ZP2k65xsqYMcrxDykWWsUkb5MMHIP+JTecnsye4gKWgJGm0fPlmyd
helzsUQn1+DhgAIIk7vWiyukOSUBo2wN5+gOUe4FRez+q5AmXERkWwgIeo1GQxc2
umzNVCQ6fNiLXAmL0XKe5E2sAMlZcEQ8qK+u+pJd3qpvlLXIiPoFWZBrgWjXl45Y
edUqmjLBRqIti3Io9N1hFZ9bn6H5bD/pZiAj19Hm6wng9nLWSWhVETwvpuCY9115
wY2T39+m95dWrssugQ7zu8wBysGsQfy515RfZAnlEJ7Jk8Teo75zjjVCipn68Q0y
faLkoYINNzPueo1JQS0G3EykfliA05QqhCOabDOI8sihFqxXPZYCx98LPVojHgyZ
5hinkGE7VZTWvTi/ux8m73WvwARrYuq4nIJHxeKsG/N8JMiPi+yk+KTZFBjwjAuj
g8EbGvj85uueMZwAL/EmiWnlxCeUdHQaFNSo6MpK9DOqkSX2+ZrkNvOqSsOeDI16
uK2H9AAxyOXmMJ2ov/KkNL7rS24mvVd7iu0YKbX5pnGOLucT/GKHgXbVOwkEHMaA
kdEfJ0L2j4ElUVAYfPKWp54A+WRinvD4diu9hgMcmbTaA80coUltOujQr19mBtbG
PDQY0564MlokaCHk6o2lLP0VV/BMkFB3Pfnne/5LqvHDagxoiAClOC6D5JP5nNOj
gaPo4PVP/tjWJFjL9aFTlnqW9YtrxPg8+f1K8xdY6rXCf0LyHEjHVEe7Lr5692Cy
TB9uMWv792fKz8My3z/sUHMwE+UPxLhnVLBNKgRNCCFWcgmWXXv+RAX3gnHOhCkJ
u32ERdFOgU6UBZviPmtVSObXK8r7iy5dxJJWofKQsN2Kh3caly08IK5HXE4PDmtd
ZxXDsN/57vVETSXiZitUFHxXcmHMhqJIjM78V1B2WEvl/Md5GZzgr44uZ5YBdDHY
C4gV7flsI0dtgP3sJGZHX/XiFIasAmllyMwFxgpveuHvNNwLqTbJeZgIAmYGqaqb
6QVuaadFzdgnlxQ3t8XTrIU2ggat84hQfnY56cGvJ8wJWGU84wmi4uaYoIoHVCkI
t903YuXpzGjkKmE9Y6ZaEuGczfwSI0ZX5FVYgm3IJYNJycGGkhVuIoDThOd7Alkh
dJx4sW3jCM2DlSc281A0flK9tLqi6OjlAMYOl0ofGk9g+mot5r13+GbAfBaaNFbV
wPs8dwouPpbr5MOQ/a3mYu3vwEMJO4+kMJpeL1prJv466VjquqtCBegu5i8gpCEG
J5PVQsU2aD1kFgRt2KBaXNkYy8LMQ4Ck/p8PFSQBDeRpvKxQVjUH50LJlYsAcXhz
AEm5Mb9WbCiedij94OTN3wQGb64BxrMrZdR1L8hvInu0YQ8a4PnoFUSnRmkLsjjC
WZqC7flIIhh+koDY0cyhsxGgDPdmXbDhorTTZteu3/WtkuuSvwu3fbpJjEjbCdgz
UAhF3auHcWWh+K8ztShbstFqBKKL/X3euybOT9s+jlY6a9Z73hhwrxxs14a7/FoP
M8T4JhkFCeEPaxyL7lqlZiBJFBvMQ4ylbuz3KFBgCP8vJVRkX8AgLwYejCpGspNR
O+nzEOqBUqo4nvSQK1oTvg==
`protect END_PROTECTED
