`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IuW1tyvnBvy1dmmrxphfvsl56dozYrWBjsrL8hoAWewSuwYUnEmdBn4GQINvCLfe
MsG0VT6Wvle9NdQhrOBz7bOGqvk8mz1g16+5FdEpxoKCMTV47NE3EQq7RZtlvtQQ
HYQ0CW8OVm6KkqTQKZp03wjzGD9RJq+aMdBU+JwjlB0NMXhTBdfdlc04TRdz+TTj
hGVZEx+adZS2ggg5Un0ma0W5Wa3FD+F/SC6O3fln9NfFTlkxsucQh65x5i4rpa65
dT4j1zCE7QJn+tcMAZqUDQ4+orRaBgG1g2/a2jHJudE0Eb1vhckM+CRFDvtidAmq
DUAegUDn6p0D7/X+b/xf9fuvqHr27jNAkBPD0KZoF+hTjz0g+4cth272c+uaFhiJ
H5tYB0piX/+eusoova0ixd1U29WHYPwZSkNgeMEpT0eKSYZ8EkKMHcrX/H5TjVS6
bu6XXQG6Z/C1WnoeZiveyaWSDxWAMkTp/YEXR5MrzisgSDgA/PilKOVl64NGR5GL
J7a1VVyVBqNwgvr2RADLU5f8VH9tpdbBOvWTFvfdSLFb8W3lVuVy5czTMqtpysqR
DpXjUhgPZlaOSafhzLdknSRfJ/ceisijESiCPf40+ZL+MsT3aeUMu30cGSgZUSL5
1Zobcachp/yHNDszdGxFA8Q9+7EPoPCfQRX03Xku9qpDQ7vdixIg2F1CT66A3aOu
rJe66prRefhOHnridcKu6c1ugnzLGB047OHos6oVA7ZPmYs5vgV0Ac39/f6efhYy
0KUCZc1dkenfCERO3v8ecx4IThk1Vj/JCYRgH9RLAMLmBWdIreELxR9pUCtwk800
1mhRX/C5FvYnqSg/STDqXKBL3QJ3toRoSZwwyIOv/cV/uyLSwN25f8j0W7TkVBTN
SkFLOEiorEY57tjT8NzPO+90e2Vr9tDratI2tOKlj/OArg2V+CWi4vfiE3C1ePsZ
QXGxyFJB8ROr21G6BwW/bMRD9jQzxntcro5xiqqTUGI=
`protect END_PROTECTED
