`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I/erek415tXVlnbb3ykH115Jf+tDgYu0+nTNPbQ5O/PHNpsiNHE8eiW9bAQ+jD07
kX+a0zUJ2OhUsBBSNB2Pnsq2vXg7kiXMe6nW8SNR/ok+JejzC8Q3Joc30Tr6MwOE
vpGvr6cKyeqcyt6WFKT89ssMjYsQogvpqJNqCr+Ye+IJ02ecFWNpNBaLDL3ncTw9
ehHAS8cIsBDzSWD2CGVrNuPMbLXi/feodwMHy7DLhIhchkWDAiqJeA/f13lu+tRJ
iJ9SFEUin/KZRB0Ha4H00TRinUhyQKBaDua5/4qpZKfI94y//EBaaM/zeXaZNIMM
PkPld7w3MIdKWgdCxBtw1vR1ngiQHkfewuQs+/6EWw5HfdSu34rwiX6J+EjfCakg
d58DWZaKqh8Y73XlaAQYyMSHCFGMOQX4QafNAfni39FlhdLkCaYdfk5F7udR8Td8
Yh8ja47e1Vd6bbqS/GS8P518wkpmkV/t9KtkLwFb+AUu8I/NUEybcVS0zR50HbIg
Vh9QKo9pCuQwIPVdSLvBnsCIuCeJIHt8sOkfJbSpg5mfTJ7ZkuSJJ0P9Hbd5WsTV
Ak2C5g0DZoupg9qDvbHGTb8ZUSH7/kwtEOxV/m/2cvoA/j+YEvb8MjoKDuvFwzjS
ClGmSBtH3vXT8oKXqLRdVMbJ7fk2mVvRJwiW9d2UVycLUXpx4u8GNh/KmmEyGd/w
HbK8opbFSYwkwmedNYyt4NAHTgB9aa61U+IV8ifxPSp3Uj2No4H8SFvQd1dc7bie
gmmTa4LY0QdBDKhvT8VYJ0D3xznT3f8SJsKX4oKrg+p1uOlTOlshvhaoE/cOABVI
JBF199oGmUYe4OBcVsvqcNOd8+eQgjHaXcTzAOrE2GWt4xKGI91q91Vd7LW/xb/s
WSpuORCD8zrDzYBdXM9xMbLErTMs0HQR6EdW7HbQ80Hu5BYOtQAyGOpg0V9y1Cv4
jo7/O+O/F7favisNR8BaPUa/UJvjBja2hjNrkrUsinPtEtWW897XV/sD7BECAh/V
4NIzv8oTj2W40xAWjEYD6SK/Dw5pngjq42Y9iU2CFMFF+0LbUY9zEOZ0JCyRj6Gd
/C5oRQpWRspc0LsghnNkedTxdqs3FwD+xWBu8yhLnP1Yh9czECKUnD62MWst4XKt
CS6zK8UhcU5ATTvKu8Ivc1n9eO/Kq7M5xZmxnv9iEpxsSx4HzwBQLOldiZpXxjmZ
S3+zu6t0QeBPDLrDvlstZi/twJlypuihL6kVJ2eBIXLkBAPg8E/kRjOgBuGSIccy
AYFw+HZ6cCunEgQpFQAmgqUMNZoDdGVc1grhUv8xwxAnFmOR1DEFNIWpUcaF40hf
JD9YQ/aN5S8g/N+QaJ0MF4HpE1zDsbZI/NXdnCIGgwvfFX9F0ILKpE+gkBhxgRha
UTVBmEQ5uAsj1Psj2BRWw1pd2ot0SpXMQQ3e2WVQPLnYxzYYW9pqTPZsurm477fp
SHQZLFPEPyMF/A4tfff1OeRydLk647R3K9uyyRXs0kVArGLX2ygv2SfZ/iPO5Azj
TNsSfLFLkOowFROLJb3c+HGIWsISKO1jpOx3uk/H5Ucimy4gLds/Ln3DAl3dGA7j
538Qv/m/LSYbNVwucZHaz48RTBuaQjoJGZemL27MC6bmnbG7tS1J4IF+svsko0hO
V4M7gojcxGpxNyWS+T3k3vJekOl6p4mR9HeTLz5xkx/Ztlg4pcLCprLF5G4fgyZ3
bu/85dqLuUiHHN9iGctZRjABiFnPMioUaseQbFoq0MR4+YkckFacYXe7WMWtSChd
UbMhkmXbg/DiUAIc7wQXyqjwAwbS+YTubGP2cTqU+w56IWjouyQXQMOS9sin6j5t
HG49S7D7HJFSuIpUh4MrC8erfj5ERcV61OiRK6UcfVK7IBhTGSWUtbC3pExxEBQJ
LKPNvtnPeA6SO4AWEcnVZEysb2osG21dsE89nMLm/ZtvIzoI6mXkh5O43a44f4A3
wDcO76QDN/eN8P3SZCIrMz6h6xyKfLs4R/28weovdC5JcPNKx81t/ipVd2Uex+Rk
lxYpfixBJoOiEK+Om05koBfiMDPD/Dyz09FlqiW3jo/ENDyD72qgfICQ2aTW/yWT
v55e1TrDqgt9JRRUeQGSegR6ucTmK+drq4CDCKiTa7ADxscNZATdOedFkhNsZyux
ZmYu5ITTZLc+LLiGhALsbFejYO+om1jMMAaU9WV92H5WQwHOCD84HWnZVDvvdEQ+
8jzBXrKcmLlgHp99CaC8Ugr5KcP2SE5B1PqBjtKz9DIoevdcOm/G1hMsyqvtYVL+
p7kWiC7a4ibAXFOULAh10OJDhom0EJu++PWQZdstglhZuvj5llPj9GArcvsFXE1c
/tZVEtLG/njPohGW5wCj+1EJvbqtaLrU5jFq3TFM50halIaAXkpYyxfqK7nCKjkC
bNmwEBxq74OeC+CIrXMNSxgY9s8Y6lwRwhvCKsa0atRYfKN5gsU8bv+GBKshJqtb
Ky0ggSea0yJ0uiTdLTDggjJoM9NP0sktmlpRtjxS+rJoKckf4mAoQ989i5adYG5R
zcXhKZkjQbwoBzzyOySZUUGTYMM1Qauk3sAWZx+TGHKuE5Zy9hiSyHZbnLDEz8GA
M/FIax1vYtr6HJDzIJrCuT7yiXKKrWd1UN0vyCLArnE81J+rGYuvPef9VxetAxbW
5PqChuP590jfaXT2MNO6+4Agt4GmMIJ+b33ad9DQfqBQ2quhpIBCTSRZ8It9UiaK
MIyAVupHiXogxi5XZ8/YN+7dGtAP1lg85l5e47QPPJ6CmYD6RT69ylXv63+cFwt3
9b4dzKxUofqF7YILs2jwCxjSFWfVN+XwkdTwbiN/xPw4yc/InkfTy/CI1glnDAt9
wuoFomssz2kCIP8gWS2iysggC0HfOrRUBG45QQta24CWBnhV4K1oVd4JstIK/jx3
kZGuD45BVH3UVau7tTQFICUsimokZ3FeoF02wrbNZiy7c1kB1v+gtKg2KOD6TAoa
vtAqkjJ9d9gRp7wu5DmX5rb+ezmSYB/rciBrPv0jljzIW6VDUL/x2Btnzjtc4nui
g0nkVgaFiwdVVlRbHWh97ycv/vGxG5Mr9CssM2ABIf5weciVzfSsQPxZETNTdfde
6v/FUTU+6dEF4+Uw2+ADjFfCtX03jr4e5tgSEdiCQCy2cnS2SzQICqfGlPQ+ploI
jkcQpwxCAC9Euhpuvxe+yveYUcp8/jxZ5yhvO77lY6mYLiaQ4AifZfsp5lNi/wFF
nO1+Dr5/hKM+R6q5xJ3Bs5H0iX/ToHH5XMK9ZUGOjyCOYGNzzdhGiMBB30vRhQqZ
MhpUibhHAqGJ+EcIx17iEKIEKJ0Im/pnV181tFH3mjV5W/VUL6HUIJSuMSy4p8T+
GbCilhLaAng+CVCv88h0leCLd1jAX5JrZawX1NFQZqqLC+Lg+mq48SJc8gXic579
9Jt7JHkq/TDvBwyWRK+2ObKPfUkdraggDHyuP/NXxEnDy/j9USWkGVKu5/i+cxAU
PbYpoMXs3QVdCRYLNNnevj3XXj37f8dDqwl7nF0Dnu6wzGUEG1zrW3yoE9e6hMll
AKV1lCExReHRZpePZziKjkspr4QAia2A5cf7zOPNDg75Y9bQ+aueuUc/Hmo5x4GA
sLrIQghtEw9tyQyjzzemu34LJVqjP2w3Ps4ABiUHSMPdGV1G9r5sUWf5ACsaxMVr
7KDf4TJ96WdpjJ9HAX38MiEhFQHZWmqp4If2wd0qzVH6aXaWQz2tsHb6gfEIgKGh
W1WC2XaH07w1zMwldaGD1XgCO7jUjaoj1veOXMPNSPayJTTWF5/B2seR/Q9F02mh
fDeSCLPGg5LgldcLgOqBRy75sc6o8Z0pTH8UryHeWTVphnVoT4rwXAbL0urJVsMm
BIMTgguCxORuGTnqZb95T5+n4ERyw4eozQk88GvE528fGuc1lSwNOpeiHt6risBB
/g/CUZdgLsvZ3J9mcaJXZo6ekVGy7YBPbFLJUIfHS3cYFuNM36m6ZMt8c+GLb5Yj
ESaTQR5iRMH/gi1PuIWebFqX/fJPeCagIPB7b76Re8EJdC8yimo5WerhJiRyl3pV
QwYjzsDEjh0KGJ/nDabvuINhY7rXCMOcquhiuJ3HTK2gFdJ6rIpCwfInK6StajFk
Anv/+5M3fhAhlLygRkcWRXIktj2l+047JsD+7/6Txh+19gsV840w/m7V88lsvL52
iPwr0tFU++xi6qLJDlqftquoGpNMsT4anPXluTwIe8pCSIO1UfU14TvkUzcTYsJM
9Bie8oRreMqeW41MOjJii4YNKRI6XJUvh5NhsnKIT/P7Ph9SipvLuMy6yganEnJN
3XoxwGBJwhcdTL590y6pZXyMGfpTnP8LDfpngl9TazINASUWHShdlO8wOLHkbRr7
/cb291qQkypP/YmvvFpJRsf2pSPguDgeA/nJkLhzKdpTIvL88Kw27ge64+l2gRxS
LfiRV9xRBYUdSCUGCfAyouO9rvYvAOm8Hj1OJK9+sAUgNh47vwnIDMld0ixhfQm3
7JewZl21/KAu414fV5zMxH1KTPDHx8UACPjGYbOPYViKum6CH92tRwond3shDwB7
hVKah6iUWUNuLCbTIAgshKp5d+ds1uYJB1koevdmC860nCcMngWNkxx8yDHeu5sD
s4T5Q8kvRNJnkZey3bxXSNy2qdX8JI4NLutqwNL364uYEgd+FBE2FstmIj088ryo
vEINjCdM97Koy4SrrrfJKkF+GTX19sIOM8hzaNvGejaG8wPDn5EOuqVEO1fVm/dV
iR6bs2DrztelyUAeiDo8jTWs++GJbtJsO9a4lACbqbbTDSkbxaUArzlds0d5787R
J37kXjiLBstGxAHzKcbMtTe48NIlD8RFYYEEjzjXnthnqjUTNFa33lA/Jd4DFVO7
d3Gyuew0417wA7Fc/lly8HLs/1/NRi/9aLE5h9m4dsZ6GUW6hmOg8a1Rzno8vsmi
MZz6aE3WJx4EftJWcx9v2J5rlnOBS9UmS3mq6oUD/OEc6poLeHiDBqhJaDxEaVE6
q47O0jg/ZOXffm7acQn6jb6d2U+I6tUKe7vSGZItGZEo7EtKPQM9TcppNsZ3tk8x
Edy40Auf3pNJWu1CL2zHhRy5SjubT8CY6IcBhwBiUqGsb3lmnb2tklxQup18NAuh
TLVeIsKy8w8Y52nt0l8FgiXPhsBOV3Hx0D8K2qblglgGoUpELsQfvOP+zOuFA6c4
Hmup3s68PCRYwvdAQ11lUJDR9WT1hVcpmpMasEAk0Al5UB2m2Dw58Lzhg8gIcpW4
5bdQWXfgzrtAaa31h+1BxAhG6qI9EmfYG46ShiLDfffoYux1fefn8m84wXdUxGrC
vBvJ+IraQ3FZ4Jk+k/zRUy+15o9+Vt/+xcmYIy8FDE1qpd4TvP6kejKUStMp1wXt
ED5aSUy0/JYc1wZbhXqQ0zuSs9jwecwISIHXqfzaQM/eG24cB2RZOW9ir33wb9WL
e8EAqNeqQHBqooHg4/cHKuy7Jg9VbjV+D5WVgjcyRErklNX9M6XPXI8V2NwRpFBO
foWuSsO2UAOnHqCw7o9eCN5iC+WOCZkhsxnWEmIdlAIDryT1yswMnSWtktxgEc/U
zbTZzRxBOjEu40f564uqhjYKj21ijCIu7TdVNHZJ/75FQVbN78R5qs2o88Sv3daG
Yw7bfQS96D6Z9jATQDi7gQQe9ZQBNdLUUaaDHVHsIlSFgzpcKEgk1NuYY1iF2OwY
K0NYqXSuRVsGex5GbNs19szvQJ1roak/mXvds9R+0NHSB3RHbocq3Yhnu+yBd+fF
S4HD0BVHSG4o0tse+hTFvOTlSYEcZgN9pisFek0RzP50Hc8bv+HzZWIt3aKmk0Lh
KFAh7200GNWJ8S0Wa9muBwUl/TazH2MFYWnsYmb3WGfBGIwyxVF3vuUH77Gp9H9b
gFp6oxYFDcmjHFhDJJQhFN4Zv6T3rq+LMBbFZTWJlg3wH6V5vzRHX7EN5Aw60Q6O
oPTuwbhUr5f5oASU2lUJoco5Q/UtX520H9+F2aKP3zEEkYAu3+Hnrq39x7t+/BGO
2bcSW2TDFzYM/KGZ5MG+586LctAoY7/MKBDsi4moGdoPaI+IemXhuWg7bfq1wODq
tEdgHRx4WN1ZKT5amXp8z+weM2vIHBn9ephjY4CHjxZYjlv1zRWsG677IR8UC5i6
Tf50D7PRIUsFdEByZ1EMZurdXNoPsSCFM068d1tLdw+VsCfTmjUFn+VEGo2Zl8eW
3xImNbSD5GwFCI9dXruMd6Y89nvSrxaJk32e9sR1HtPGAxsl4oBuaD+66QqfjJ1x
N1Zh5dQDxSdoQi+JQOqvHKw02LPEXuBfP9zeJIWQwlw79Y6Hq+xF5OPRS99Jq1lI
Gn13FsbAzK9drdp0HwTyzq/foJX1SwQPu26ZfIK3/k5++7djCobiqKouq5/iswot
CWxc9k3/4pSF1lZvvrG6QwlEinA8KTCdcb2dAOPcUZJy4LrEPeIY2Y5Vmn6Vz1VU
3b7UJIR3gLoWJCrnFw7p9JWKYHfUmMxIBYsj0SZhG+9R5WtQDB66MJALLkIuUfKV
RNWbB3bBpV+ySlX4wdp7CIciIc7Rm596b72qCvSwObNNMBnID1S2cRMq+GjOeRZ+
RAFsRF4nOkNgaNM2iSNVkwYs+9AZByVrxIeBg3CknJuXPlNa9QXbM4JWDGjCWR6w
X4LJxik+tHh5OC9oAB68NI2cPjvkH7VkSCXkoFlCdpHZsZan4EFbX5YZzF98l3ys
CXWhoitEhm5K7T8h76YgEKHTJygSbSghJgc48QtdHLQapONZR6nuq9Ny5zAmPWYd
aqwPfqwaMVE92ldzptWSFvfKAD2IObzttuCZF12leVocfYz/BWU20S4pXAi9YFC3
HOeeyHNiVZzle1pmKUZH2uj83SiyzS00ub0N9iupJENAI89N7LDsnvkMl8pHFViP
YowzwJA36OfE4u2Ay8R1pptfbux5BzW85wXLc1N80iFwJX61HJOq+quNWTL77Y0M
KEMSyQD0BSrwBDdJEdhKxeRGJmhVofpkKeyqi1HOfhTodpav8IY4UcnMAIYrmPAN
AntJumMlEe4ObfS7TgQGozrUBDBTMEvJvOxEwCI9PFu01UIr/5nELRo5ouF58Mk/
PCSDV9yZ4/zZ+7AyDDnK/IzCSp/Zj44KA7PT+PWhRyah/IKguTaak87Ze6asV+9I
C/GHlXa4a38Pwp+bs9y2sG5QhsK9KbVXAdoom/fblJDxRShr6D7/HHHVxEiWql5C
f1T/RftJHA0AjPpio9XPp58IVtGFUCs8aq78wUbgMvWZh1X+Iop8ghspGOAIH8Xs
pH8XDqjLlPZarghfWVDctGxqTDt3EAycJLrqmjm50SnCyoy2wYzUFhSwnjigYemf
HX4qGTl3qIQkwFveVu24w3FMNVr0csDtJa850uEHgG5M/UvFOoajsDRw3AZflb6M
13sWiCz30vPiXBb39fpOZg5lNc0Bjr8wBHPd/aOY2TFntxaT/sEkRS6lDcNrc5oM
T3Qhqn59m58ojKeuYiGCrEQbp0nOQLIlcePNL+Gr1FHgXY3COP39S/NqnGq/Cre0
Mf/Kpo3ZD5L8IXszLhLHtyuA9IHfreKb1XEBByXP3BK7O8FV4zJjpkcx5NRMSqJS
qTj5NR2Dr30GnX3iTgK5ZH9+g1H3kJHCmH1ZE+Qu0bjuRQKlXVu7WoIkm+WKtqe+
tStORDLgchF0CerhJwOeZ2cR0uIjHZBNa2kG5ppVofICt5365Uz0jocIWlykUhDd
GNqrq9nFJ3pwpFU+LFwGtsGXwQjP3lR6SfvELL0nMSAPxScSQKGDpbuc3CYsrx92
lE4vYiq6BIKMOH8QdRUwOPFaSc7aH9LeOoSCI6Abu6+jwL38pn2rgaYLWxSC82i/
odKmLd9j0+Xfav+yFiH/XmJuuNmkkvM6W43asxGOiqTxbbggDoRayzNlo1wdS65E
LZxUav9JWS9XJwIwkOPPetszyoHJh8DraDf/aKJCzMTaH91fPYnByqEZaE5dL9tS
biZOZzkpzvvO1csH4eSpHIOMAxh8j2LW1lC0LOF/Xzz4lpvMpSzUoaZkQyXifHyX
bVSZuT1t+yjqir11WR0iQjytWXd7guQC4Kq8JP3x5+BfLJO41GUkz37lI+lteenS
J7hFjkmdAeOgYJOOQnxj1wm/BpiGR0ohQMq3XULd9b7UAtFU8+9b5h/7N1H4s3YL
oi5N7YMlU/cZXy/JxXLBqWQ4TbPo6m3PEwBR0gB1riiwYVzpfARdehZT3uj9yHc+
06ozqAZjqz9MOuoLlLiSFHb9tpU6dEOSxTIMHo7AYH9vOlt2E1nG5EMw5lbLQfbE
0sNy6FzFsz/h3kqA8L/A+WQ9ZYTMiRGeRAMOHZVVhjLksDHBfmbURk8Lr7AAeuAl
BNUc9eiprbRdHO3t8PToY04JSat4xMBunYcqUlNFE1sUIo6tb/WhokxX4Qh3Jc/7
8TA07dwtprTbGB5a5NVf7VsNlM+EYcfcdjQKJ4MckvMIdUuM/j/WbkqXeRSGM0wG
E782OOJdJudFEdds0pch4Ew+Qy9bFu8xSTEE8kK59ZBwyAe7RmTxyfOWCgmRo4Z9
xAuc9QjwWM8iJbiqEanfCLSft1ytXqAophFOZWbDaOddHnQMAR/JPUE0mnlRr+qH
m9O8q9tEgVucV6+OxpRJqCosXhxoLDgjAEnSJWPb6chiRlItxC0SugZ/vdVfiRa3
twVCsld5JtnVrho41EZ2nLpRcFzdYx44tQ+5pmiagup3VrNDeZn87jHZ65+XxNJJ
zURJkmN7D9ylnBtHJ1QkKdIzPsSam2CIZZq0shK1F3qRtrQ1pKE4DfohIzY4psmx
rjS6vVUL47F4HjFarIN7FIhM6alel3ZwjvRID5DQ+mX3G5FZ4peRGGzzPrIPuFVg
VrEFDUnjduUnDIpt/r8va46q+mKRWRavPDuA9D3I1V1KFEOP445cLv/UFtijBc/B
gtbjgg+B9x5WTNPLW8Ok23AuVuZO0irdoLrxdr/q6OmJgWfcgBrsN9ziavZyE795
Af51iX8kqjnxGtmZuIzjb67EEhFr370vR2I5v7GTRbh82940tjSHvYMAysadCYV0
MVBuf6debDL5iHsn7LzTbtS8EIJ1FiApxz4mf/YJIVM8tcFqf4MOnV24bvdV8ku0
muk0G9QRL53cy/4bSCwriBWx43jY5qfIUIvNdYklBGcyQ38QvB+pVI7zXdUtFLHQ
oij05Jp0u7bISJcUAof1LbSpIWlzL3O+Lk7crChnw3dMvjyYIaNBUehEQfojchQG
TnmC9SIp1gdHTm56rpyBPM9naE3prQrdtgY00eK75NmsCj3p4FxJ4CVuOn1IA+id
mshURyklu7YukiLgWLDw0WBv+uolpw08F0xHnAmLAVPkRLr34NzKSv2QZiK7MIaI
ndmTKHBdFdWNYXXLWN8gnP7Y+SL5E4x8amSjCuI2qDQVbPhsfP1//on0LqaLNhL8
zFj0EXF/SedtcFs6nvglA+ALRZ3qd+fP/1EOzON69miCWqbBwhOYk7M1XY3n0/0k
dZEjiWDGtFrcQrIW+YKF9uupsQjBHlzjDYMVTlHaf0AHARVbOKyn5bwD0cDM0ENP
aQiOxymZ7yAiDNcIaCVWJ2+IGWBUadshRzjgs+Xyw+8r9ffa8tixeKQuy5qhnRrg
WPRfAu+0inBFRKUGo7XDxsA1o85J7aFAfbgyw5g/XlyGI0x/3JEDSqghQ9cO66gs
DyFY4mBPum1XcZo3dq8fB7YR8560oaNAwlOMmFvjyEoLIAShtMHMFF1uJXHUevcn
oDWXQ/GZEqCclWr35X5cEXyYqzS+lrsR7Tv8LJ5oPX4ETSsUxjMcJERcn2zM/4a/
voHUJfZP7IIelVG/f+sqvtpyc6SpnpR/7LKAZMkI/8nwLrr+oZwwVlbBt/Ub5Ekj
WPCfR57ArHDbezaNsoJWYdnrcrsyoBWC7PZCiKXwitfxzgDMb4nfIdMORZz6DCDD
6wDFDigW/+AbTC/LMfOmawQTc3PUuws+DxfJrH6upiMcCIbtNyzxHsWR4xpv5Id+
sp0CjHfpaJ2wq9mDaOCEmS0Z7GaV9s4S2PAgvUKeTvV+ckW9sCCsi9IVAWF8DPmb
MgvJxGzW5a7ZmVveSnopLgUEkfcY9HcNElzs46O8SC8AhmVCZ2G1XIjGZn5+LeIm
iw9iXrFjxgmt8X0e5FF5PYS1rhSJyfkUkL050YPTRDhhEkDm73Sq0PlfYCnIJI0Q
oLpyZmM+NC6j6Nqjm03QO3/KuqY1o0ngFyMZGjY1bighD5a2C3P0LMV9SSf/oJsl
awCcZx+Z0VjZsa+HknpSiq+F72nKWxQUl9aulXjht94lD53B6qbOiujH96OSqct8
HkYFD7EPZqdsPVwk1aFf06pIzWc7N4DhHkR3CkMu+m9Z1ecLQPe859DqGv0M+8lY
AGfiR0BgeyRH4cjwy9uXXz98/Ys4dtFIZUnZqlYSUm5IJbupLA9h1MyNDvullsP3
OEj62InchD3IaPvkPgUVTQ==
`protect END_PROTECTED
