`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rM+3ARJGy1Hh4vvllhWTz6ocAMysJPgDhcK7SguFiIKXeIu0rUcZHxCI481Psujq
dFKtntAOEi5xo1DyX+g8hWscN0uHIlthgybJnp6uLzFCzmiO6r81TOchBmBYl72y
PV9DMgkPRnqhkDx28p3jPtDM1OT1mIVK5LwBe5ZsEL2TisfLHkSiBT6e/psWT435
alErvwtb3yX5aPNAxa1bGxe/YzGQNnA9uj7W/YY1UIX3324dMtsUCmr0UyLookHf
YQTruL3LS3JS5F07gj6KJg8A/GDAcGt0NQ98D2OoTS6g6BmS+49H1W8iUp1RBWvE
4ZFRmjEZ+4aQlCrJByKNLfsIKc6jO/417y+9eEA4RTSOEmcthV6kzOZ0V9gwIKiU
T44h7pZb25MtIZaC/dfwNxORTNAxg0yLDUQYKnbFvptFeKlxooWIzeXCCOXc4aNt
iSWx+y83Ze8Rpie91Muu5/aHONjHfUssYMwIE/cg/KHPqqvQEszoXVg+HRXpbyCA
phvXm/0mwxJJL/fReu73Z/sLnPwbYJ6O4yT3Chg7G/0ZisLP2V9dbBmoVqmMU6Vt
AdwB4jgY1KPweBk1simT7NODlLTEkBK0tJENjmU0eAVAnsqs9o6ct7VyPkihC7CB
konLO+Q9py64NjYQ4hZxI81055rz2UYlzNuz9qhRbaU36h2qTeIvdzGPcEHoE4Gh
8Ci9il5RlH/QWqqG7jYni+G/hIq3eJH1udQhoevHlg/bcOhOrh8xiT0NrRWIOm1m
CgJyE7crVvgnLpCquuAVdihcR5nNV5jk3OQbskHSdqvO5iDgpQ73JzGvDknXhvaV
jd7Dho0cxn9xDyi9zM5ARAStZWpJVxo93NrdqMqndBerXcAeSeNI5MljTO3c4Kbj
`protect END_PROTECTED
