`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8Ia5q9tQMOifEfUxHsaE4qtO+oRaGTK/I5gx9W+wPLAPvotnK5x4B++jr1WD+Uma
HhPeVkBHo0yLXu82WQZT7c5aO60Bi1lsW9LG3K0TCvz900Ijms0U5FhokMO/h8ZC
11WgIlWwHTqFoYQDXP/0FOpnnzesXiggqFCyPzWk0XipLMCMD+1QRuSr4njDvPCQ
2Yj4Mgink7dAeRymNqAzC28f4dkPiBIJXmsqCGYdwLYe59Yk8u0zqxBAcSilfkYB
CM4MloHjIyj9/5mqUT1zeuesJvxyB/F0hML07IwZo/tCz+UNBfmHQQ1d4Jp3ptY1
kr2Qz/1JSOOF9WqDUaPAWqy3+R01iwpex4hY6UoA/w6BI8/0JaoHoEabHzvvUc8N
LWUVvPHIGzWUSqjoSwFS9aWNtPD/KqMZL6ETDisw+h/gnojY2AEFmU85nckt8Nes
sHDxNFxELmt/FA1fKi3A9AXTox/tvwFy0pLjwEytzUMEnJ3MU4sbQhTOLdUS94rW
7AAmcWTY3sN9vOU354Xoxid31E7q8MQXrQGnm7n7XKgZtYufmtZznFjogg9MXI2m
vHP7jEyCgoOD6R1ZHXdIoRBn6vxvb3F6cyi6mLT+Mp9tYJOTZhlvKZVlkXIRkHw2
KgZd00+Z24+IlUn/ZRwIhl9xMAyZlHnhWBO7K45xzWru7hu6GmXJLtoKYWvgIU0t
XKqkH6gcaega4KgkkyzvZ8uel/P/FdXsB/CEatolKy4dll1VDWPZnVDFpKw0YVJ4
ed+kbT8adWHNdb1Y8C+n6385Y7RmfVPnt7nno7O1jiFLlsGZj597ls1hg1HXMux8
k5umu4PRJoukzi/NrVoaLwB2f6wLP5ezcsSmCZWpWhtDAWn7CFFSDCdnSYDJ/9LO
l10A0WUn/LouewJJUbaUwZyjWFEpBo1sEQvlL6lhJntgl0fJEPfK9v8XKWXdu2uV
XX03UxC14bXpZA2LpsHeMGlemIHxnLhgFrYYfSkb1FdW5puo5Ta3Wy5CTdegQuI7
i+WjRmWl/kEXlpqJXGog+g==
`protect END_PROTECTED
