`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TuGfnM+AW0auk13V82Tst6nC0P9KxbQAdf8HUaP1J6dToIvApoEG/4AMlsFwzrCi
IMXgzNxFigcwNot6UfSu3fwBSvkz9Xqp/F2+GJaW1l+wstvVZQs3JrlIGi6r0Mk3
sqmjDiI8qh7UJAEPt7LDRNFOvWMt765m2jSUOxyO4trPiqFjcCuVA/l5Pu4wOJYV
JyQTdR3bjPDwzDps/l7rsSDhLkKv0WVvzCF7GcH+KJJGy/VfFuh2NEyqUNjdNSkt
4HFml8ypgQ5b9nfx04FO08FARcCB8tJU5BpcbW8B9wh62SFKDEMsjmdYdE0ALmAz
OY9hzs9i/NIszw4bEIQsqqBojo8RJeLH0AjwCsdF2AyzCxg7dU1CmqIX1Sh/FByg
B+d4/N/1ClOzarHa+SFBe4HVlCVQQ5pO32MYOtggSrdNn+uRRNmilARJgGjVmxah
5KJdhyPnphp4xm1x34LXP3X7KC1Oo7t5mQJxE1Z5lBFun0ugmnbaU7oIU5kcXwXE
O58tf5x/6HTtyVd1GQwNV2P6Im9Ppk8HeaCzGdgdKN14kXrKffKHf9KWd0Bus+xQ
d+PtzEVkC8IpszchTtjetIMULcqNTPEVQ63GdeTDvqg/S1EGUkb1BMU44h0vZXNn
1w5a2/Nf6+jyYgFVVzXDpKt0L75cmUDUXjijgyNA0ijqtZLwYU7vwY27Cv6r+WLo
jnc9AWrZtX5Lmb7EE5WHlkPUL/AP5bLVgPhVMtucI3ROrB8mliTpQshnUeL6NDLz
tGkTM4iU3sTLlIxaQBzjVECj6u9hlXm4jqEE3YqqTuNPDP/2u6ehuZ1CVKnYttDH
He8tJy/VVdyJh54BXqKYV8T+xEaE749rYdKpQgLJSAbbxtBbVQ19TJoxDD1TQdKa
i8XEaMYD+/6pZKaskAYQIPGwXlDWG9cghlV77GKVo0WaoJDsObTDuDDIsmtO/ckn
ZBzMJmkTbHLNDl8V0nxqk5jRXw+eZmlWpn9BUy1siBubQpd1IZhlLem8emelqKdV
fRmTBSqlNy65KypUYOgbjYG1aqOyGI2uDk+yzUS82CRCM/KJPhIdevNtYquoV7hy
d6j42r9+oWODdcVEuBtQoCUgAKhIeuHu4wcMh8VOAMzZNgzRZWdTtfIRWGZfMr9r
IbTlDqowl3VJ62tHDZ2PhozbEzzKeO2ov1yP8tvCLv+fLuXzqPnzGqrjxSxKurbm
bPb63hDoVQViki1+11u/Jd9rWAxPtpgVU6uSR5YzAHbBQAI8rP+eRS/TrZRPSSQA
fyqyBOlKjyFjSFeyQduv5D0xqeuU/zt98JHEuMnDtRj1+C7qEGLQ5R/XbA3Xt/1N
sDL3AfjMq55vRhgOt+nk5VN1cisVNzvllWTdpDL0qV6wZ72VkoitIbksspLqK8t5
pC2RsU9ijAjxdygtls+jXy6toGLHpOOoUm17lK/NctqEcGhc/ygMUw15ATxmCJy9
l7+rJUWULEUeuYw8I0XzZ0kocwoONUaPrg4Lo84x7oGZFcUUe9UWnG5aLZtQr9t2
zXwdMPfaw4i7NPr4rjWaRHOqrWDyNtvSvhP7bJPQZObMts3tdOuloIO5KfIHitkH
VHRrXvpdCz4OGvEt06z0MDRSsQ4XzIew2P2LaToxSZlnFQcIgc65OBwpUkWF3ken
ZYGE4phfwgGx6igoNe5aUWo/gW6ksBPFenxsd/jTNTjNMumi58HTqs0jXljkD2Sy
nn1CO9IHYn47ZwSl8XhpwTG7pF/3vM/Dewl+5OYum2cXblFdSXCCchy6cDPvV+xK
TtWiATdWvwV+khul96gjgtlOPAr+Nhy6rA5tvpoGnZuElosvjVHzWfDlQPbIRa9W
vv/ovtNcwHggf58SKulIUJjP2sgY/l6Ci78C3psP2rkKCEE+2ocoHFi70yZ8UTu6
NQxv3szcaomdm2m6hI3Xh5A2Q34sh2QQYdUvvWZVkFDbSZQgc0sSo6Qq5AGyVupW
c5A4TX4D+NQBgMiohAk+udrW81xJpEbwp8+UrHv4nC769SwhF1nQUArslg+MeHYq
KHmwTRaW6GsSbFOvVrEEVmmxv7lCK9dMzbD33Rrs2/UnGh4TCryfwavlM0Pl5sl4
hF3VuxnRlsjiQtL8VO2E2f3iQiZHKKzTRdIb2NnIX+pPrgy096g0+t/EQYNF4HgY
H0rGqg/xuj4dRrBwpaQEJVAhgTc/PYoA4rxb++oSYNcqLwzEcXx2ky13I8OArW4z
+Gvzz0adQGFsOqfXDHK20JesjUuSkuiC2vFe09oW/gLzcuWmEf1sF6P/Xjha6pZz
GvcYKXiuURRWFG5kDNkLbyWL34rQP1S7NChxdopT568DSOVfVf15exMnasTAAcbk
RSSZBb/1mg8Ti9ai47g38b8qYACiCvwvLAzHpIIkKunbdSRA/7lmxpMvS7RjCbpo
`protect END_PROTECTED
