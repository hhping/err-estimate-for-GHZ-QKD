`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TjZVBdQEaGaNvlktt8MAYAn3DNhec5Q2wpM7ONhXtl6gjxXWzyQ+RWpwEZaaabVl
4U2w/mA01Z1HP7aNLfr4Ou+hj1gCKnwk1QnXZ3RBLnRcIMXPoUTYfywofa+N4CmJ
2WiLAbJrZaauQKSURDYDTaa0G50aSeOCZYM6TMdyCRvcFTpG0XlmkkoE6u1M0cw5
Vek7P1c71XWPSE+i2tGPGk6d1gciYdPVBOskJju+9ECihPuZYgAL6mAeQW88fw6G
5IdHw8l0hH5n3d4Gz9IdF0sukTSetBggeOuFHAw8MuSiR49ZqIlxGNuFtuHfmy2a
cwnETbutXc4rjWiuiowAh/82J/rAnHlS4LlhpQ76l7KIecfeQlFLj4nfy8pgANUs
aL12r8ZNkfL0Zv4Lthxv8eMrf69+FA6qFneCJTLeuNHDLiwMaXwfSc3zlM8jnSjF
i+JdJTiwGnd20Sjy0+h8ubcZXwR1Xb959TkzRedEn9vWEJV2mWCxAbDzD8k0XkxY
AepdjzbCwdSqaD69Pxmqt6sxNdOy0rOiJD8+eIQZgzIClo2zfJ1rwYmXF/2byM5y
blt8ToK8nmzM96+LCzCMtBA5FjAjabAyjUtldYdXPzsTnK6CsZpIPqt0MhBLeEFs
CggE/U76n5nahj979p4oD/6DCnaQoDdVfgEVe30V8Cg=
`protect END_PROTECTED
