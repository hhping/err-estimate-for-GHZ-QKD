`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9dCslHww1DdGU25s6ae9/TC6/nZxV5d31Ka5boxWkbxX3GPN9LqKZhXSd/I3Rkoh
QP4YBV1z7xeuJivNA/Yt2lKnONPlGGDuftwQ7vAAg9XKBat9p+X5icu087vJDTPD
yIV+wrisHo2ExjFcBXJs8sTiXSdrb9UiMizLrUog6NCz4vlCe8QrEQBLEQx3ypbN
FPgcpfNGV/UnVOD37C7immZ7EDdUzOzFlqwbZ3fOqarioHK78iRMrqCMjvHF+G7g
mJWUJpZ3kv8L4woJGVyVkdFZG6T1e7X6k1bhXtHB2R5ZwYlEAc7STWMX7hYfxaY+
ycW7mRLWDysQGLpSC6Np2Rv8WIVQBqSZfrvTDXYw6qQPnyhB4YH1Ae/LLcKg0Gog
MYS5011Un1wdEe3dtW8rSE2DL4OEnhT3Fax5AeC1N3VuNmYC8TcFDGHG/jhDz1OA
224e6Sxy2FRamw+fvxN82gPH3/VJJ/nvMhE86BEeEAtVitv6/rqufSCe3WDH7Acs
t7dWLHEJCX5dK1AEE2MnZMITFpD1kBDQEe3dvE40cvqlw8Q/4+dRNIypiPswdFtC
iaxBYGKZKKpV3cqPclMBcgjlbimyD6W8Ru3h3CKqZpg/VGpD2Z6tk26na3Y9F3Gi
/sksRPWTiU5rb3fvH4Bg3zrimq/01v7qrJBDTFon7LXBD4j23DnMWLjF0QDjP6Oj
XpjWgB7XA0F0hpOMsQjoIDftm5POCtm/nUuZ8UnVwcyYmu1xydKVXfF8oktzEMJP
QrvPau9hVBR77Q/AcemG+lxIamrKMmS4jsjIfkHnLshQ4m/lEhea9O27esL+gWko
LW/Fo2bgsVGH94mQLv+NdrFsyQCNtv2DlyApXmZLG2mvvtU8/kKHQWYZF1HGOk1w
0AJyba8YVUR9lI5PXy1HW8zr6YxgdOGDh6CEBxvzZZvY+lskQFO4pWVL+nmrzW4r
2diU5tvZ7abRRvxzXY0bhfCcZqmNyynA53JD4tGsMYbVaEhMv+35Fir3eSGRBy3G
a1bfncVgTXz131SqCTC/kSZ5aCUXWj/ZGKHJTitKAzFBdmlrIc+nqurUTNyfpA3A
9/5o8jNI6km+9pbs9JiPTAzKDP6ZIdLbjexN3bxGkxERaw+Mpv/VFIDtx6s2GqeC
efupqeIfnwkqnMOYpyfy9RKjkgLAwfG4Nj7OKgtu69alolkq9qvuIPwUX+ikk+GR
0MQPeg8EFLvZVmlYRPwdTQn1/OSUOksQcdyuUFVz2r6Ic6nU17+DvPTYAv5/vJNO
MNn7PqnNOH1uPE6XKdyWZS0G7gwFBUAatNFNVw8KSSJ30p3bxG7IqW425CBAprL9
qvaHLlGkBF76IOss8dUmo/xEjmbi6i8Irwrye+kqmrslfTj2SntVbPsWJozUIpSQ
xj29m/+2xc24bZVoaOvv7FoOfzAk7LTJcpPEXomxY9OQAO/5jaQc9ViimmUtheWq
tTOEMq5oYYP3cQlzyxom6WvFe56GZzTJtQMyXnw93MNBGhHNF0LA6nzvbEcwrIMN
OpKFMqY6+W29pT7lgcbrqEjH1ymKNHbO1EAd4QgyMzLmaNyJPn38RruFqByiLR+j
TBkqPjHYJAiGqbYGCPdmquRuUmlWUIUtqNeS5r6rprxPXJP0EKh9i+lssdM8qcL9
LodbU0k1SR5RUkxo17fYDx15QiT5hIjcdQPlVPsObjRMKRTH0zD4cFcAoVt0DAn2
7gLwyq0J60DQskK66ysWfOJjr3qJKTJmrOnAYWYWaCjkxJmrkJ/Curt9DJRAPzPj
GmjUEFhr/HIFRAwdqZe2q9M2IlNy1U4A1bQ12XhWtfvMdXtsrpvl8pLaG/E/xLeq
R5eNyVNviwbrF05rhMEKUm2MTIhoDbZj80/8rSmWXtzJgCgCgZnhYyA9f2DR8nS6
fhnuBrryFHyKJaqs2QNhIm2fqMCAgIPQDSlzxw8WMtWU5yubEZlF+GuKjTBU4FTm
urild1EOqg7b8gqYCLUzoNToE1VkUL+e/Zpgru4SXx6yTr0ny3KE+lUO9ktFm+KD
IKa2jSC/popqJdPEFdkxraU8SSPDG2pWIc4pVLJVTYQkHqW5/tiU68rTcTnlF7Pu
2DE5T567lVp7dbB8D+pnr4TlrR++7FOQ4xjYS6V/O1rw250mlNLOMKl7F1E2b5iJ
OuIpNa5EKEYjdtxtR+qYfex0v6KQ4iwgRPx8x66o/zZbjNQuw7+lu+g6lRx6Yrt0
rYgVrmbSKhGxzUMF70p/cH/JLTNAtp7QKB8FyHJchldHH5TlSIgoW+p76ZEE9YTU
dJgJiOfqqzsaooVi/YthrCPMW4cEIbCEuBm25oKQrzqFbxY7A//PxQkgDeM4/vbp
2o2N8kZBCiSphP90rLlsewVBYYmQVscDsP2CxwR9MrPe18w5Pz5xAw7khsR34ck8
W9/W6NUP+MtKpXnWLwZKyZ1jys4XeggqskRPAFE6ShDHprNwVdezAMaiDhYndpZh
bFn6wcCWDpKOsAaxP6YJEqJZcJsaN0m2HnJGM6fS3713NtIRC7GTb2XSbR1HBhYD
S2mIL6VKIdMB2PnOlxkk5wQqINMW0J12XuPwauIgTq9fmCwxWrqJmRMq9U1RN5+8
Ge7GUKu7OU0lk8Nskw3LNfZaM0W0S4IOiOUWRi5bnM1hzUCwPfxP0nQ8LWvs8HMa
xW3VzyTW/MM6nWqMJt0SgBkh31VC6EmZPKjxyiaI+3NXSRZx3h0Edy9VumP25IPt
3i3SgJlgHigV/8As7JSkCUT8QFPnwwOYHON1dmwIPZwNkCmF3QG+37usHeFsBN2J
5j9af+feSgoUshfNuOvf44uMclhn9QK7Qwqv204I3sz0fBLu//qv74wecJC+k8De
T+F36lPTAMD/Gkf+RK4UKL/r0NySk8Qws8tK7Zi7Iyy6C6OuXHVD2OWcbNgpB6TP
8LzXpblv3lSNnfb7qqlb262d8Y9Q81qhjN4u7GuKlwsAJTApQ1qmMswtvL5WaGzJ
RQK+KrJMLjMR7QFWQBBqypImms01alyAHq28Ftbk8qmOFqj65WRAyJFYJZCF/A9h
EwfjoUXXe5a+sV67OhAAjmjGJu+8p1wEBOKCw/EGMxnWCp1rgiVxWGxrGwtGMIw4
M+ObBcdNB2c6am/T94LC5ei757v//5klxMnCpnmtiCe2XHYrjv/HhBAt9Kwetvnp
URiKMcbbdKIKPVNqAzYJIN6jYGYtL4j0AuBN7wED0Qw6NgcVaSFrdmm4uh7EM0II
aircMe42VePi9eD+SUTh18ceL7hdkPzu3+zY80sP8UJJECbzjOJmozRgyJzetXwf
KFf8nJhzjKqHEdLUCF4zNrzvsW97E4DhLPNtn4mgEYK8ec2aJR2V4xRepBuoeAyu
v5S5reYDmvJ1ShjSrgqm+EvO7H67HFqIiH0NDJPI/B0bpU4Qn+teP78wTcS4EQ8Y
WIOFsRpaMxJA9oaxPsFO50+xcArKjYgzc2TlaUeUdhppA9RysFUFWP0ue0V3ZMKf
QuGB9wsychF+HkxyhsQuTeKADHdCMslSuspcA9CJzM+ONtJnKilCpzmMlsmQGFiL
f/H8HslMaaIwtEudj1qFq9q8/Vrp1spIkNmEcwBNJEm9NN4oAAjZPFdqgxnV078v
BYSukNl6bFMDwF0OdcqojmBp8ZjN39NTP+eGND4Hs4xHE6nGkcMoT2dn6a+UqVlB
UeNbTKJy6rncq9efLA/dBTRTJn+MnAdJova3VZVKQa70R1yYz9LY7zlr6+n1vx05
02rJwBDWz2y/PUF9MvnKN3cglTAVOlKg8ksfk8NKKYzY6A71GJNqHSZYlGhj/fs4
g84Ccg0Fa0JnfbVAZ+dMICy+IAUF3KY28FuX7alekj1X28fC1QMWGrlCU5LuVnT9
RvwaGWLt2BVHO2r75EHtV6bjlkKKLSLyFlq1WukhEnks3WR2E3LCKIEGKuxXgaFZ
SxqyDY+f4b377WMxfnghUs0DiHEA6pekRslnJlVngm0eGcnxQBq8gXlfOMpbZdtS
VfXA8I7mFSSBEB+wuPrs9Z2KN/ShFPxXWSp3mQCvdwSnBSzY1t47TEtRNXU2REvy
fPmcQjvGkd5hpBbrzog6rEXxKXMUugex4gqNMedzaJ3qJAh8XSssv4g9BW0cBzKr
xzxrQHOw31L35w6mdFFzCu/VB2tnFhvHxcJHjQpd7cHigP/WlLPwHnahLEnqL1nb
IIRGYMD9FC7/WaDFlM2kgL2n12iezkfoqJ25bt1EFJwudBUS1RwYEpuAQRG6z/IV
apHJA3C5/QVgRpV6aeA0MWv21Jk+MMmpi7jQPSk1I1xm/2S5nU0HvqCHqmgNTNsI
jwAASZD0XT9yXSIv+hWlavMxBJkirULZzfun+Uub8QZGPLuxJOASlXxqeKuVj7Wz
8RYkCYRW/CyDRckUXHNFQtLgYEJjQh+3+MVuhOfQQ3pkaPyb4jZEdzYrtg0DCLee
HSbEHAPaaC5HfsG6hXjruWL1y24Uq0jwlhb2VEjKQ9HQU95hkXLMf/zBXCPMCWhF
ne8edfG5oiH1iYGimtqUPyJHz8yR39IHE7tbXBde8rJuclThwgy8XIUmaP/xeNEy
batKuho5gyXShQz9XSE7V+EvFFLBcyFtyG33MIqtCXs/Kf5GadQl5avwcmN1fLh9
12zLiunDnk8YntGZB1u/UQ/WXY3eD6IpmyaPSZxxgXyIyGX6kMZxBFgBDOxxyB1w
LsNfRx6MdU7amyT8gGtvEhtqV6BunJGwZAU70zty/51kubnMXMKuHxs0CYjMxXYs
PE+ob8ALysBLoWX3VCCH4fZCs1riJ7+5eQDNlhc6PAOBaP3B82HzCRtpsB6WaK8w
AO4pNbMjuiAlyHi7m2Ud0nEVzAGt5SN4Ob6X7sBUgsacGM0RYIanFUMRKpD0UvVQ
iwrs9x92avxVD93uh3+GHCFCBJOfc0a5S7hw2GU6tedje/z4wcPFeEOVlXGNbpBf
/lYtACoo5BFYqNcvVHVEP39xtge3keYxj8xN7L1k5qDe4iEVCh5r+R/LUdC8IGtI
BkVuAqsdpltHoJdJ7q0lnGsV8ptmJ+BtySVeGmU9dhyVDFtIBrWhLeHWqLnz6qcn
khInLzW3VEbYWZD87LS0THm7Y2JJr4pgJblA52yF8Rw3vEVknkJRWEH2eJg8qqxq
8Hk/PhND/2DgQ36XiTtYJYIAV0Fmk2sglwPmx3+RrbgCSQlx3ZuLbHDEvII1WPvd
3WPLorzLI/N5ZqU7E4LpkgEOJT8LLboBOXIE9TRZeF+BxJC0txESLA7cgBWIo0x6
NDFvfuQ2oYzKufqePwhRG2hx1nxTAJASSHJD2tol42uO5telOJdYzoHNepHCAc7k
197Tvx2rWzj87oENnRVLKAPKh5MCFo2OZgD2pZAMPBRLooYfH/ynTpzIO5Ui7nWr
L40gxHcuQ/GNdghdmWJSjjyLjnUQooc8XWWOAipyL2s43zWa9D58h5GNwr44F908
8W3Hn3ewlPGMPsADdSlNu5OdZuNt97UiH3E9EA9ydRa/ylVfqCmzB8QMS69o19J9
xVJz33r3LJFeAGTKRtaAi7aJIh2LM/m5P9CCd01uby+TXLg74smLG0wbSO3gFahT
g89sqzK7YVzS09E51JucOB8IjLdfjzbXQ2VI1cyIlK2PUkscuwU9R5y6X2WsgGBz
zyva6nYAHN4YtPDOwJHfFnEePTXANKLDsgVUJDNstkieS4LCk53YQ5ESe5hlMWcf
HepbiODk0D+BlPcXVFM4gADXOD3LV/Ui+7T/VFT73cAeJa1Cpg+jA3gOEkTI7Gt8
iSjElmi5nqw1JpbeUQ54SQnNYx2dLbStkykJDrXJLVlXV4KpkmDpZ55vwkEGLOSY
ouMu9BHw3+xBPfoR9hhieO4ldCq6Bkqxu8UdfDkBsw7xA5yJbEJGDJSX6oVQMPz4
iOId9UatNHghedHh7LbfPa/zmJbhnpwzlT//W1TQ1uuj7gjl7dwjF/FXK1u0ST5J
U7aWHdfVkJjy/1dU63qqLdwfyF74Y9oUaMtfsP/WOKHK56n2FYAaBmr+Uspqxely
BaveMd5ZiBqsUM6YaItUU796PoysVPF1N+8VclCZAHyKBIF7cm0lfGFEa9FMUpxC
J0824tTBuQvrbzsa6Cs2xYZ/wG8iKEc654t2wXKdXZHQtJZzoBnZC/CF5KqkBHU2
mzlF+AOhalAj1rHxwBMMvAjk3iiumS+bD6Ro6Me/hhzVNzM+wwgry+Im1Q8Fnycu
PXw/vSVuLmf21AoTUW2FJ3HXPhq/8JsHkYq3kD0jGGFTU0Bz75VElAAqoWOOpCOc
crZPJ/5MPFERfyxVIz0vOagmzWu6DO1hqa+awVIxM9dOj06dwnYyGlkrZvujDiVf
TJMdacSjT1V6UtkwAg/Tqv1BtcGemF9o8BMtUsF6TP86FMkxn5Myw8E1YbhhIQ88
/SGviieuB0JxTv8rlBFh2ktrfDwlnOjrZ1upoMnXaOxxqz04FYM/ipOTWh4eRvLt
BHzKH6GSzhsvRBciui1yf9/vx7h7G9pKv21eVl42xpYReJ3HtOzuXAWtoRf0GIyb
PQG6av/9KROTajOXRRWMLFTy1MTtyiFnXzqCqNOXO9mKWbTIP3jzHaucUnhK4B+V
BUJ+7apIdcnt6m5NnI+TiJfIlxDuhVhLbJ07Ts+bCb2Y1PwZxA8K3qOMUxqzZEmk
V9ffTlfi977FVd7cIZUqqoDFnDTW1H+Qe4BdAaFdGUDtTvj9gG72CSH6agBJn7v+
ZfPG7uvdWPOY3EHhV7cGvL/Q1BErMugcFJeAK5eQoUj3c2xvtPVfVvk+2DjKNOti
bEuf6/r9fwF/dnhbMMsPTjugVi9QK8kvmiN72XL2kt6lPgjsqzlulJp4Dlu5AF3U
s3JzDO4RMUor/mwQQJx+w82reNVPsKPjbYBMaHDeOvKLw1QdsViyqTkaqbpcBOmN
hOsZeb2/ZrglryetT5A3+z7SQU2UKoubndjj3m8fO6NKRSNehsErcTALWPSQUq8f
XX7IQJn/KgHhcJlzq7Qy2eGdROhI5Zej3Bzn4/xQwy0BHZLp1rSuWNrB4R4zdin/
PLlNCGknBzNu0bv+aGHqX/tE6nhvDe0LjGzyA0Div5Orv8Wc/yBLGLNUy1tzK46P
OFXRf+dT8pjbhsdOv7xLmF3WQ4LjFmIEGmCp2q2yCRFdQunS4x486ObEIUbVdzGl
vPdtQ2eYTB0SdMaReDDGk0c+DPYmcypdFgfhy6cMxVy8BZGWJ2KjiHFHu9lg8HIN
DfWEeFw00d5ag+JDdHKE7VYFDQhlhYiIFAMWvr4kEq043+4ihxFgjXhbod+53nEQ
gerKEeHyARJRWlKMBIfxvJNBVcsHPnZ8sbJ55LinAqH0zQGagJVPYsnfRGp1Nj8n
LD6FOW64Ndvo9naczVxGb5Jq5HoLeatov0y5zXH5qtFHFTfouRtvvwmCfuC1PFg8
qc5RC6X1KxbOFRYddY2CY60U4H+sePaDRqnVQSkW1P2aN1yXbdQ6rqOPPwrQLiTC
JEfBArCOA0bMb6UWhYwUmrkGG1P0+/8JC2UNKDs1CGQqIX3OSlpwTC9pvLmY1j/7
gsB3DUIwzH3Ibl+7YDUiOybs4NoMDQcUCUTP3XXXx5/0YFjdi1CrNhFbXZlSjXOK
qZr8WxOb3XAhgTtb6gcL0Bo0Ismk40OTDQ6L7UluzuuYcL2zgm9dyvD/mVxepadE
l/z90RMepKocTUZi302rCQrKiIirxj1D54Uz1cVqDPSY8M31mjYjWHPnmKkTuWry
Zmz/SwgcbM3oBABEjBaOPqQjhCQrKA78TNp8s/9fLNntc0tJuR3H2PwO0AohLd7I
NlPVxwlsf7N2byTXmEU+P6GUciU7zuO6U9378DJFk/gvGAcKsbqa5j/qH70EAuPJ
pWlCUjbEO1xbduHESz0YDHpaoyCOblgttNbSPqAuaQ7sC/y5lLB8li1lfUjLc5i3
yYsA/vm8b8sRkmPYEandHoGs+tevIUcKPvMumjTEK/iZmiTxg4Bl3nzKYmlyoEgm
BkRr8n0RzpBr8wfSsHAsCcpZCzNaCm/CatkbyEhO7U+I/kiX53zk4HKLW19z5e4I
rwzdKUlUS04ZWCtLL+kBaGuQSS1K/cvJ7nWsl+fH1TOxyALfDWIKt7gwg8NZGgSW
3y69jY+iHUqLdZxbuJF2sYKZXTsgKzmIWX6MT5QKDWFVhuwcHkRe33J1DljkwUoi
r/8v89Zq5JSGb3a9seuELco5wrizWlQ0Zk1usLt09qzpiR4BA5tUl/+E4AfOKxTn
Of1OUQbF4Kw4YJs97nF+r8tv2N7/GDfvTmO+0uPorNLzgDsWjATmrPLEyNCtrQZz
B+OERAT7pfj62ecq6Obux0DGAXDukeqqP2hT+bTKYN5pG2BYIrKr85M9ndSGGlS4
OUv/bYr7GY8p8fPVs+ZUT3j6RGQR6y4xWI7HtdpfgXzb2bPeuid/yDruY9uCkSKz
AfTZQsvj63ld4DdmTKXPyrfYg4fq14KhpEfTnSbsrDxM6Ng7uIL/W7nBHocj8pQo
0UUc6CoRPbo+0/BfYM/+wMbNwApQOLV8+DrNPMh2i+YF4CDa8BBUH1Jbjjrb/xaR
M179zr1cUN0dYFJis8NbMCCUSOkXZUkCM/Gbghil3UlAf27NkLm0MqmUu09q+tlc
pul0U/nxLdH95WR6LYCBhiNqCNu67sT08mW57d1LzvTZPWbXDcdsvMmjbGu4/5rN
scfF3ciarYCb6acntBv+baWuzKRTH5JDb2m3m7+Eb0utOcfC/vZEBD4tpwU2iSO6
zDTEO4ABC3s5Wc2OwDnor51zSc2ChICqTTkucTewM6S7ZBE7CxWb2887nBho2NYG
jxTaCOO8hrzt0J8jTh9tk8MUTzsw09+jgqhRBBgPFC6P/eXxQNjR7FQUtF2RYjeH
RkIYQF204mrmh8rEvgHH6ihCC2B7vDclK9cx6rVHnsjjWvlzol1TN7flJZBc3cuZ
iRIR0lfHgepU8VDwSwIA6yTqqfRhMHJb420PnjdofUfS29e1GTV3PbBLMDpBPWy0
0UgWUj7w/mUv2V5PH0Pvpqj/ve+ipLetinFzvABBxOUPjFsYOkOSr7iC9niTIkE5
P2Of9SG6sg0rDydIHYSFqH2AFBnUKPbGhmrsInUDngQ16kLcrHPrXU9nBLoVmwAD
E60y2CHEYI0jtrzOQhrAZtPD8bum7k14W8UYSL6K2tBWbCCglnBxZaXwpLi8ncPW
aHgY2sp3HQlUOKpR1GFYxHCnxB0UyE6KtI5h+ehfQtoQ0vFKTrpP97OhZMSoww5R
jg7rDagH253AfTolESmS+Cn4JC7I3VyToNkkmyYTATAX+0gPGS+29RT3TAAnKdGe
zNHYQGuNqnz8fNvKYonQw6pko1mQhT8a1Wi5wbyO6G8QtfaKcq66dx0hvyFH965D
PSocC++00T1wBvacKre85TryVw8iPDcHC2KhHVd5ovl6JqwRQVxB9iuCAuYISYDY
XJShEr+pWxlPSW7Fin6bR31gJXuLDB/l5HXlfN6iVXYF5mMceAHSaWFaKmupjJW1
714VAtklOGQw4P5a8hCFVKWQnpzcuARx3b41l7aowxN/kbhWgfAzfjG63EK8PRAE
q9sV0YCare4+Iu7r3UwCD56TE9xEPpdbBPh+m4pzrtCFVQHPk3g24bix5baA+Q6d
wcUszJC9i+Jbl0LwaGhl9kMZMIKUjBjaV42Yeq4qbT1eSYoBXg4uN5ZTjTdURPUP
+Rk4kYIdzK5rCUgdjQF7vt7xjdQgNiwpUuTFA/xBYtPbFJ7KkSlT+mBSee0JYC3G
uqLLdPCFNM/NBRJMkrTtqpSz7IC6AJbNds/bTX22HkE/JLGrq5hBy7oO6PgPYOCI
yS2I44/+rYt5Uvee/VM9kVoKdqjPKaFhkFb1XcZL8Yci+k2hX5/zE/05CbyRrzhN
WRdCkL2yo0PigUf9PKzKTUhxvRWSoRh50AM2TeIOgrpKSKJmLFZ0JU1Au3m/7pE/
vaijOGVeClz3Hmb87FDJV2zVtWTWTbrrhTSRJVAYKlRHzXvaaKpmEtj+fBoOClU7
27iN1Lhey5DhKdXmPKFfDRBYwvhrZ7Dzho8dN2MmRTfUb7ltsPXvPiNLFUVl0/2C
NQ68tPYTdMweblNmcDYOgTSNTW5wcj5YrjEeUbE2M1UQj16uEq1KegoLykBjdsDk
SUjxB48TkiKopvt4iT9yPoz9FvAvungAYKpjqqauI4yMS92gkDLyjPDBfBgvnptB
+d1p6+1RRh3mmveDH9mHML29JatPAnOQE0O7d1Lx4Rj1VSlqWIwz85pmPO4ifFaH
TNluE6dRI9hDkvXUy2T+6/jiKPL3zq2D0N9oJXLyoapbRH20OWcoelGUzfEk0Wj4
T2nkYAuh5iO9LphGoRp6OkhsqXJnO84/3wj22kM+kePi/SOEU0GaFnVK0ObB3hi2
GJFjzdWh6L3Du9Mc508LC8WTvS0FPqO6AnTA3ut0A72zQNyaUS3W+6yGoiYYQLKU
i4EyGKq9p59x+UCcqShSO2M++TBRX5WiluktlCw9qkIHk6pIgf2QeFPKU/Eb1emV
iNHbmWOr5sTEsjwK+bMM1SpJFLKSdsRJaRjmOuIuzbPMfEh+d6MSYGLqHvRL/87h
IyLrwM/iegAs0n2BOeCi1Qke25Fec971iMilh+CsAh7C2Fu2SHSzP4FAvCQ8Hxpt
+vvFH9YRwQuQPI3V39sKwIL2jFhtEARaZU8C8v32KU4fLeIBT/EeIoI6O5ytlMZc
kV40li91AwgJhxZAvp5QUyslnKlqiCYi0y53LWLCCQoBemavGRtScthTEkOGKUvZ
Pzh4tn2dfIxH6s+hz6B6K7WuSTWUpAeivxBfiJXgxqBp0zC/OtiHw5WcrFKBQI6i
KjSMdAzLhsQg0SoGS6qWjsnaWaGwzhXlAQbfZ2ym0Y5sfRnxjBmXUf6DUCbtgw6j
NmNkylBlJVZz27//KCSXsMVYjnVGZ9mFmGJnekJL90gXRqS7HnCA8uTkH9ogoqtR
H7qHw6ZLifTCV4KwnBkPpcxbfx2SCQylykUQKTCAf1C84ny0RfRKEhe91VQAjSnx
JcVk+SgxyT22zckGQeSJT1TD2e4boWMVMN6v9XeoeC47cwJmRnnUTxkbXuMAEWRe
fxK88h51KVyLUo1ax418kCEu9ZFLQ1+miLD8cNG71irJBkz/0moUIOXBfhPfAIUE
HZssBpLFwYSmqYAHn3XzK6KmlH4ldiKlXH+P3Vj8nxWB2JiVrCbZ2UYpb5hXhHnD
rdUVZWQNCvvLrYpBEfVT8wRrILOUzSDNCU0F6Swh2VChVZy+6fG+uTLb0cCEBYdM
ZGm7dROnBDYurc2mALEDuFmybYnICT0ZFOmF8vovXVsKESGkv0qE5XRhqKVjCvm4
G5tWrpZr03EHcO0AeSwNCDmRepdZy1MOnXqZxBloKClWoOxnbO5XPocIHhTMQpU2
xxZHGde1FDDns6V6BMKN5loe2FRH/FSH4ac+KG8gkq2L8pgH3oZvuir7O036yv1G
Q7elPRNQoOm82rVjvOGjv/p00VigDjEAAKoTJBa1cfpqG2lBDb97wJMA5iB/BFxZ
jB3uNL0+VFBnaZ1AWS8u4v+L/9//LY+SWT+2ftpLT2el++HSwhBYPE3Hu4RocQpg
yQEgItaZZ89hZ0eo4/y/ctbp4SQ0zumG7eIrr8dZMjAZ5cxVOoJ4AceifFZETyO6
fbwR0R1PhAPrrrbRMrfdysk+eRUIw+tAKfL8TcmREiIf/95kayrPqmooZANFB159
8eKMz9V+PDszqphpc1tTf42EV0B5EJDVbMvj/5eHTHkLP/uYOgUhDm0T7m0eYFmW
BI8u0Vlpctc66Jc8K+/EQ+aeotltARWl4zWGFZXaPNRij33GWgh5xLp5FkYVYQ75
+N6FZBccJedw2a3T+OG+ZDrJvIDzCJc9B50HeusuQa5L1XYLAb+9ErxalSNhjcbB
Q2MVGcgXZEAsKkbMfTIA9FCqNsz22Q8NUFA8Wfddcgc3YXY9HpqyFMy8vRpP4WJc
MmbFsFPZH+97vj5THXHWGq/50cyLlfjUndV5HLw3CufT+dGK8GhHrrJzu6lghrPz
oqmz180PD73OSA70x4D+fIacPPoMu8i3iXlHeMdtIsVjIujFierxSmWir8w7ot3L
Vvyy8/IwZ9MuHSo6ceQpnMEFFSbMKFge2BcurXMxSMz4bnoue4k6U9NgzIc4UKml
91s1lP2dchrLnvJBj/vZC9gniXkGVioeEl8mJcWqOt7VDrTkhaBGkXLpyl1aK7Mm
B77kRYrVPXhWOKXfiWgMmZ03om/SS97r34KSIiwMlwwlEaNdqFxHAWjQYbI/IX7H
pksiwNSdjgPjCTc6IJsRAjPW6PVv02GCrHPw6LYphbXHyWb3QolboNKUuyBujbvY
0mpxGDhesc6rCcm+0XDxT4E9Fk8bncnZ9QrquPSk/u8wnw1RTYPNDnbuYMpBu+Fg
khq2+nrI+3fGk7W4fPzurU7MEhyQd8msgwms4mezbLWVQYyfY53/R8aaEx55u4Uo
SHXgS0+CwRXB6Z87KrGPsqUOf4lkcVrM+50jkuiG0TtNAF+515h+rwlo7u6hyGxu
3mL25ooX5P21H/MuM6XQwgYzQgUWduPtGMoe1ewSQp+hv+zdWXnKlcBpzeN/9WTk
CTaeTNN+L+gqGzbb5+v1eg0KzboqL/zkI82c/+yFCtTYgmzzua71duIfuApJQVSj
OVfqnDv7b7smUNNwWL4vntqDqSFXtPzUXJTDczQ8EuO7RC/UTOqM4K8zS9NZuPJQ
fpN4nlF9rvIZfTiqVDdLy9Tc7Maqf8qWIBW+kAS8fOVcggDNMwkUsaOGT1aTlPQp
l5E8nWiwRbLJxF8Rvf/quJBgqF6yns8z2Gcqhbbft4oXkFu1iNjmCW8afhMusWNX
yL95uru6DJJMg40+BR1Ub4c6n4g2Re/ErHiJY5SG7CLNaph8xi+qOSK0ZifHe+Ou
5KCIzTtpePbcV3UgiQwr+KroP+RyQ/0lLbJ79PdCGMqUI+SYASV2w6K7SGHPmrg1
X2yQ9/+H07FfT3FxcgK8RusOeDa1DCE0fh1Zp/vHOsOTeaNMAwq70AsAJtn7kTr0
YbKIkVMPBlqiKNrr+XALU4Z4+YoZL/gN2zvmkNnGApX6G4lRCvH2/dFYALKOO43Z
XAs5MkLKkibHuPJ4uCF7VwUnGZ/M5VOSFeF2WPTKN8zWdQhhqf8CKKBHqX1zVJL1
B3j+Y2UYJXMLT46YDv9xQHwh425G/SDo2DNdT7owpwz4AdwZj/rJwkpdragOwoI8
L/wUey0O4g/t6jWfjX/JVOQDI1oIxsVoF8+71fLOMY0o4bzJ9RCeFRPcqrtpoqGY
ne5WqDGilMtaXp6HoADFCgLDMqu/AyAx4M0AmBccDIorcElCJSTFTjNZpFcekN+1
vAZM76qxLd4IZdav3aZhuZefYLpuAHq6x7ZHKsdUw951SjS5H9rt5vunuTCb6OSR
3qJWdeBXT6ruj4UKemSYqaw1W1625sxd2NfVNiyikctflX0AKeJLGDJc+f6za/Cv
74eRSgCDSRah4l/XF8vFSZ0VFLDl1HcrC2mhJF0ramy4FCoryMqAoNOHEztPu8KB
kfHgbKYhv5BsO6YAFfsddeErwXrfiNcyuuSZXtTxIr8C7EdUDEJ851ccoCQHyNuH
ivCt9/YI+PrKDwLv9wmT1fHGq/l03kVIRNPBc1jRPZg7zosOUgTMbR561I5YvN/Z
dOA/lPeJDEUb6qsAyt3q4yGW2i4vtZjMIjrkYnoSZPWp5oVM9vXXQiTV50ahzjac
+TQGLNL3b/3lGpimPuxYNVdmsVHGVuFybaacmaMy0yz8sh+HSs+bDHhSw5N1cS7D
T7YUiR9gMxkoymqKZZqo8X7MPC4QOyRqREoPf19f0LNC033zIPazvg8gBF2nf6Ne
dt42wDzQgS7agX19us4JRysxEgEuf/wfUCiAFfjvcYBoLCw/Ci6pAPyKD3I0vdrv
oOQA/vLIq3s4uv/q5XZfMUeJ8PiL57lMtzIHNDv7ANSwE2NBqXr3XKiaczWKc8k2
wdU2UPQtXc5cU/Hd1mch8c60USP8lq2fpWL8+qzLy92JUIVqr9WxZB+g6QTDlVgd
fwSvl0mqxXNSq1ki8xv3ZITosJazzRxjOj1YwguqgZ8DxjfFEr173MEsH5tsqKO4
kxmMX7T/eFvAvgFKFJEtZMzjADhFWLmg7FbB1opLJKJQewnmnJpuKAR/l3PPNLRB
RDq+yrrxapZQkPrM9ErFstJluV7EQp3KFSOjV0RHUkZINMJc8STI8CTHbQXsZTL1
MryOiNaEo+cL0+lhRtECJZk2a+IPM8ucqO2gElPya0OiunJuXB9U2TRBJZU6Ixio
TTjK/42H5p7hHjYsd7f5mWsmKf8RfMuE6osvNxbihtk+9/158Z4Ha9x4s+YYGsLJ
3bpbe0j4glw4VjJgzDpkkwVPoybBqrXL+tmcJTzr2tKaMi/LCJ6OUIqDHKFwntaS
wO0Fzc9s8TkSja9S/1v8f6bA8Cu7yoaCeVPaEeWzLzxZaZUQynv5abTxbuv5zuty
z/Ep6JXABkKnP3LVFtM82H2sVS6XkWojzYr7ChDWt3LFuZlQ6b/qiymjm1T9vyXH
2ZM3yOrNYB+8z01sHj2edwgZjS2iaqI6kDQHwty+9OYd8LxChFCISbELSzcIlIUr
4NkZLUSVu+NPBDjT0j6wanxF3s1ajGinsfOnIMGUIfwWmHudCDl+tfNeAUNrrZY8
GlQ7uISB3b9LRYBRD+cwj//J47EfmCgQH1pYg2XoAz+EzO6faEcOyuZ9p22AA5nO
O/lTBaUnnh02Ph0EPT5TmsaiM5AN21rIGCfGHgo4AlSVp4SR5h/1wGpcCG7MRzUd
EVHdiuvCyJtW65WOOBQntf0k6qmRkvzIM8KHuZKfGZL7gFGAV8UskxlRJEzpK2nk
KkeLil9iWHMtPs+nCZm2arTviyrQTHx0+REYIOCMPvPRHkXsQ7tBE5gHvvijs3yY
nyzirU1fmKmtjTudLVKBbPWG4egTxQAtDxUJkx1qj1oEOjLX0YJYg908R7gGmuGs
dXmofH/llgY/JjZgGhRB4ecwUFhz0jwt/vZriAHqKHv7TQ7VtKlLDcM0XwQuYfWh
JtpbxbwK+rK9jr4YqHXhtSUtn1eUzf0mid1cnJyDIaAydg1wnHoj3l2UY8pQNqLc
XgxQzcIYz1o6S6kmHExKWCItUKD3PA/b2Lj2x4YMvcZREfhG0kRc2MuoBA8sGIYo
noNd0qCIg5113B9WwwXJj+mG9ZwJjS0pmkQiUUjvyaQQ9FaKjMU6G4At1qOjdPKI
68PceTYy/l7o3bAxNrxlBUlRe2wMaorrPgNyaUy9bjsdrHcCi/POrrxPanCjkj4i
ZIa5PtbW0OVdtlKXCL/vH99HHaZiYGGCj7H+Gm9ftHL8PHkU2A2Lc2U2qjaXDOz4
wWuwbuljt2Kv/Y0GeMIQ/9bZznCKYZJe0w0MzfOG/Or1kEzZIoebaCD9MkS0S5dX
gHQNedR3BJXI8FiV6CNAawKw1rIcUIEVXCdSxEPdClHBVAv2ri+QVubPBA150H5b
i1gwXiJYGd5hY0y1FmtcjFQlzguz04Urf3SYmHFCtR8s7XcPi7cdGjGpo/vfkMKA
pqq/l5jyCReEhuDxwSlJveghHa9NpI8dF1FQ7jpV5+Su3qxto3ZVNA4bfduzyYsQ
3KsYHFqzt0+WIpzqNYf6DSioPm2F7ODBAzclbWzyp/kf5lqMFp3D1q9BjSmrTxKY
s5IgpDvgIAok0xFbo5hYa8oDMHVX93WH6QxQXsOch8UPvgFQYF7frQUi8g75zV15
IqqOe8rYHnMmpJ73GEGO5DwpGzucFQfcB7+i6GF6uOLf/MoBBDuXZWXeYMEiaOlw
4KniFgXXuliECXRdCc5LNSxGtQVjov5kOIOlU2Sr35U=
`protect END_PROTECTED
