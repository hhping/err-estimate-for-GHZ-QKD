`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kc7sxyv93j8WhSM/mkPrBaS/GQJF4gZ3NNLhGhehCTkRqMJXzC4trR81XNuEAUQJ
EF9/AImlYossG9cND2kp65OXpaNlJfhavCLnKABEELRv7Z1R/XrCIkduh2r5BTyT
HXsDJDpcWBCdsIHqh0JWT0V+1P8DM8Htxn0J/6QdRnHOXYM5/HPqyfiJibPCv9pG
HfeRMjlKMaXkbqBf50MyKgNqO0oJuLePbX8c1PzMU5OcZPn6QENIRR8zu0sYwBrY
pZ9/k2ZM/+7JngdOQExlPxAuo//3XRxU4fHnELYqGPYye1BzLGk198lLcKqgOhWn
im324FJtizIIZ6dQOmemjkXyK1i+5eHpxbMrwDQamPbGQ9p3MaVIanTGv2NXAT2L
0xBjkRZ+HBA/HpSs9la7ANRuy+KPBwH0xt6o0QZmZmjwK1x33LgZH+mfvbgWaewj
YS+vZ9hARuOOL+9oNjLb0tJyV3MKYB5af0gsjMPdOZ1sdGncgWFTtzcC+nEhIFfP
dupWSCs2MFTgUygGQ+aCkqjlZQItgDGwMU3SGdP+i0tfDEqNJiAdsrGhLRxI1TKB
d4y3yAoj4WVw2FcrY479sJMpf1RGas2/fWJQY1ZeOiYJLajuBDSYxX73+hMxi8Jv
y3cmc95zR9/BSVcoAGnmjBohWrYY4tk6UZHy+LJy0mLmA0/HR/t2BwTBUQ1Dq8NX
93ZNyI0ffy5U33o2jct+TNA2BR8IJ0gplzlDAW29WNGXUvzCgwrWAjKD8u0EGNsY
ZbAYi1+QvB4dqvRL3EFjBEMQ/e+Rczo7Cz7cTzOxfbB7nq92OAqLP1UFkkTzCJPS
9pSbBYGIFCvJf90L71bMRJAkEcrUJlfoH424e16JaUZ/otLD5EExKYRmHXpB8z3k
11ID7tFkDgslrm/iVwmql62Am8lYuQUzDxPlFf4DaCjgKlXzZSQ4dISjT22Am5Uw
AzTIhRqq/lFoGVV+x5fT/1CbSdjiQheOfw8XcoMNsOPcPlcgB0VqdQuvp5dQbrDR
25hbhwnue1U7JT+woDv8fYOCbZbm4X/k3W3RgM69EMXfgH6azWfEFvTWtFbGVIy/
3B0bxhjlB8TfYZRI1O8Oy8EBgMBWUaEST3JxEmfYraaGfqdPcfAhWboSmVOZx67G
04QixuM2GcFCfd9B8fkYbG3i25OwwOHNbV5B8JVsaA0BoVufl4CBWc/tIgMwEvaB
qkLstgYdL81QahE5YsXxOZD3m+69uwWMU4F6F35tbQsSbTqnMctSkQblrD/efns1
o/muMWnpr0Wv5Tz0+HeoY1XSdkSHsNmIUcQYJpcz7xI66YWcfe0Y5/pSJBPjLz3E
87Rupo8ODtiBLm54GYPJWADemj79ggX0CnmrBnLPkfrRfd+NleYITYjX9bHp6MgG
uIcrxC2bi0EK3s1XbNQgmmiAGYCETifI8P5sw479HHoPq+urCrW//+6JY/FGQxk+
izM4w2hew9++vNJqWDtwEzBbAaoZBwobt7aUZaQa4A7IiNjvv6bdTjv/IvnqpRGM
vsqJyq18XXdeq6qkzviUM/eUYy1ffolAuGTvNE2e5g7nMt4d5A1PeAf3jyE7wHnk
nZGVHVhDw5Xh0P0FtOeHjWYH5fuq9WlCZSCdhEBGarW1QXHKPv738iv3vacAPlAZ
`protect END_PROTECTED
