`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FzDdCUu88g1e0L9rZSXBK2lR71ktijV8KON+pilqpvRLIgHF1gGql2fbtTJxzio2
jOVQPktWP+LamVA7sOaqzmUARpn/JY3EUJGgydbn+7xsoIh6xEuxhJOYotnlDnAS
tof0QNqYXYUebrRDgKZsYDGOT1MgPrZ2hFt0WgrSayUx9Fkln6pPbzNyp8AwFZh2
tdrH146l8lsAqWRBAleRwywqauekSWSKmkwo/+FGIenUXLPpyvDpIATEMEX6+qbz
8piO0TYpL0yDGe4HtqOBQBYhazhaQ9FErOLQH+1vN7tTYmxfJr2iL7lXo79WeEod
`protect END_PROTECTED
