`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8qZ9+7Lwljx1EvVfMGE44hVDPC2RtW2LPoYrAjS6apvGvuH69AAvhm0nUUtlEQ+g
wHtqgvoqFXYolHvX14DIblqHkwmAF62V7AxUBAEmCiSBDMo4+8vKfzEkkb50bRNH
7FZ9QcBEJz/lkrxZcOf79ToKqICoxrBLhPz+57D/VaGGUzMUC4TfCn2XZ55Cz1yY
vLWlM/TsSQIAunz7zWvOXditT7jXbV6nVeR3U62ZGS5NswQPXVozfSmdeHCLPN/2
slWry/tFpE5WnJkcKPMFQ5d/8RylanF2zCVH473+mRrUsvWrkMx76FgutpzqW+f1
frNid4NhwFVGCJCaxzw9SCDMZNliRa/goB8bdW+RdbMWkgqB8v8QlfM+ldbBqpso
dd4JWQWtx7pd3zlAvve6O8tBOVoq6y1ztldASsCkF6YRguj1JpMAc8yf9EF/5RxD
Cocnqf8UN0otfEpURF3oVePJJYlAH8EbqFn37+bVI+8TbpUXb9saDLWkkcO4fpjC
eif7TgTdpfTTjBbGCn0VIMlETxpUcQ0aIcdeI7dtWbwvY/ENJ/T9oXJdtLZAH8Cb
81PVo1TvJFSZNFP+W3/LwcbI7g+h3XBJr9+WNW6r6+gkF0UsqtUak21bFXvw6uRa
LmA4MuLh9u4jZ19OuN5lH7Tt3UZKzUCPNemNQvfGXBMSCJjF6m/uTGyXqmsT91Wh
ISsceo6UW8s2dRR6Kcv4ssJ8C8+h5eLTrGiDXD8ekfFzijUN/WNHBKdNfgH2qC20
42p8VveeBC1A/pD+ZeAOMLvRHzfr7XnLFYDjBNPgC3ahHPCOfiWKGFE7ru8isiFi
yyNFwUCh1qJ/19w3DCH2tMzkYk7tT9mWoBggKT5x8ME4eKvVESc19u5qVSLi290K
07xTtKgRH6Pf1NK+bfraH0k1TbtIivmpV69f9jdT/xSxFlCDTicxsvfOyfO8Zqtj
dzofYE3PfHbPPtGyAbGkCk3kZGCGq2cp8r1aEUNPcXJ5ixosWv2NZRrmwrAGNR3H
OSUQQ0y95Tg9AgLX1Ndvgksnwu87CIwhYs89c1SQXupGHAJ8P2QlTPaEpCpQVmQa
MOWXeZYzBMzg1ihx7GCyytH1n3goadV65/8pCBGXnAwjt1tAz9EMDcQaRnqcOj5u
7KTwmcFbYV3yIjc4N2Rpw/NIZ/lkLtHYQnOuCQE+mODWTL3lR1DCOJRk+8foxGT1
BV9NAgeC/MW3Tbbe3m09hKjQE14LEXTZnGY+86q8TGvWZdm8/KUt1SpiJycSPQt1
2AJFRJSAyf/BpGEi7iyOA3zyvsZlTfAWVfAb/xpQktCLj0IzUO1uyxjEkk2/hyw2
3IQVRplOXCGRFXJEgiT8BPBW8k5bGeyjtLzDFnC/Q4LwWapN1I6vwmkEMb7yF1pL
xTv62CTTxp9HQW6sg9KUc1WC9d4tr7LB85Z+TXtdYAla5tKcvn9666/Le/Y0nnKO
VlYxUmbw4i45yD7krrGT7H/civ0ehX0R4sCwzShqfFzBDTgqOJvtZYljsZe9KhyQ
D8ODcWgbLWrjtPFzOBLpWOL8QCGCG6Br7ppdZIRK5E/3BjC6Xqc+YynpArPMPDX9
9ydGMobRSmrKv6n/CQjjz5o2yj41Km56F/6PMeVQgjiFeAb6H9nhfe2unGS4uNVM
zKrJ+yg1ZnoBoCSaGS+J5FndtFTdJ94oIPN+sgwrOk1RxXk5DJDzYgGrR3OLiNG4
U6fRc8OcZKuSjJ+QDSUnazGSFa5pjj71vYpz3hUtQFw7lwrAWSZ8MKZ1TBI5bxVg
W0R1dLb9qA58eWkqDObJ0DD7sfYooBrWoXvDDA85aXkXucWPS1Ch4uZOWPWEzW9x
VFWDAZMDLkWkwR77dDrC2n//RSvxQ7QSQCPhS1EXkCfbXirIBVG3q+aPjwuROfPZ
v7/RQV7jtZF4oABSF5KV91F9pqzemtTF59/9olpo5Ntpqmzt0PoxTAwGnMi0G00/
dXF1n+hNrdxNeJozxl+rQKVA4ZewcGoQ9GFkcfeyevml0RGDd/Xgf/NgfeBnEpgJ
O/5X9/swKuUGS+/Hn9KMNGJ/+U+HYw/baTsJaq3aqOQan5lmTvOHH97SINIdVXZA
Z56JjU9nBxsx/eZfaXGlUoayPwk7cigG6lne+FVrCkBIRS1VGCR5dx2AFddXvfpt
eToti8Omtj3lA479luVONUl91I+ReXQLZ9wE9KJyc9vP2V4eDAuDEpZthtrYGxbS
pqKvv1uF5xZ0wUGuiJx96ZLungX6oeWf5qfaiQ8MWBd+7z9SEldK+tT5j/gRcMcS
kAhC18aCIbtsZfLIdON3b5ydFKJqCNx0hBi9pLwHKoxjk8fpCzivECOaZkbxZFUR
bbIRWBt59Z8eLbaVY0dAlsQDO7b3ylMm9sN+Z3EJoXlZn4tTeOkvh9yUOFLjNRO3
PyX77bhhTzOd1vygN2ApNTDb03J2gWF82qBM4v4K//gMBjvY8bC6h6hzAqQyAy2k
AkxV7zljV9Qq6Kyq1LuINPqSqCJGM0zivLyMStscooUwPJVIMGbRpKBPTLZ8wOQ4
TdYvmc+fAeL/gLIswRAMuTUGKRVmsCHGpxgzsZ1v0dTIrg6/bFubNLhIdvKbqZZN
+8+O1vieJTRFulwQlT4VPOhaYKwvA5Gd42JFF+f18zdVgziitAsQ10izQHevnDs2
9x8NW3ThigI/TxtSVv0Fmpn8yVU82OjYJelB7ldTbYEwDy6fwz3w6LGu/FpVvmVy
Q3Q9l2dj2vwbWUxliIheGxcSpNa+XAW/aAc4hbo0WQD9Lw1kPFfDDd1aImrq3vGW
d9VXq5TtCGBuWtA+94WWZ6EXKiLTXqJ9JP2nkYnG6JSddhG1Zxnlpxd8bGTL0lkz
/s+N5FlhvWYDJZkUQP52xPy7hCznpoi2776JgOqHneAJi6+N70NLOUWXLsisH8Dd
aun+Z9eQ/AzU7Vsg7L/R2Pv20jlDshhqlgR6B8B+y6oXhXOF3n7XoFfCvUjhMVQx
cSEslbijRSIF4emoav8q8ZtPtG+dgTOc6YktmPRhb1ncxmt3GIOtz0XWnAlUdp0u
xmDiTmS/pDVTtVZz9Ig29tX+VEuzyjT8sV9feEXM0qEABi43XFMuiAjDRGp+/+ep
MDLAjAojzJeGAqWmbxNVOxOk3oN1Nj+YarfxxL+6529JFOOFPcEwEVApmEZABxx2
wFUeF4MzScnDoDxJIwLlHyDPhpktcrPF/EKkwe23SVoX1sQhmgBRj8IUuLiRXYym
kFHV/QcnBS8uDJnKd4aKd7R1/0FLSP+wZRAcBmETpTC6mjw8mgSJS8WirRb/K8U3
JlnHGi1n/FNYyN2PnJ3GolKWmje7ONsYhddh3bAqVa5SuPV11WhHTjL5XdhmBPBf
4cK7kgNGLS7vaDc9bMgQGYqDsAsdDH7N6tEJtqFUBdhdyDSs6d+AUkvLwFGRj7op
l19dKuPv4vmYclZZ5LlB2Ie9/Pvp/hOPFmarSU3C/vK8AiO71M1O4XsckVqGqQiU
7Hor0xQQFWtxj7VI558widDQfHbSfF++IawHvMHWYFUmdXYMeAGZYvrN7H687tCU
SaJHFb3MU7NhBhM5AAXNQqkXccZNmcuIJImMtUdf79A/AVG+/AyBbI5KP0+xvkwH
Y9y2RwqnIY/bBxSRh/NBXS/32DSsh5+e5bkWLgjAsBils17n5F/Hc6vpgbdNCKB0
dkjaddQcqo84NYQO8+SxicOYQnpVU2mxMq3WuR0KChyGIBC0z64wfpgimTxl+PfZ
f3C2PWLqzcKcfK0fapD1M+fS8dg5KEDEQGR/iCPV5nb/jiQDPDZDDAjuDVZPnFD8
fPyYwx7kzKs+Kop6frRXW0R7nsK6qOQlaehO5FOhFFlDT/IKMiPbBf50JTOxKuTM
KlZUospBWe3ZyIIvyw7mmyQXpYCvBK8c4MrXwzWmO28QSa21eUZuYXnu/hRqMkhi
qRO+fWe9tsuGeaXDVnCJbo/lMgVr62Xeb3/OUXikcS7RYKx1w1MbuP3pq5Wi55HB
UrQqfq4JBq7hw0BzqfQxYGritNFpQyMtkcNS8DO9UBk=
`protect END_PROTECTED
