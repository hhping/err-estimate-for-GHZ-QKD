`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NvC9B7Bh88hXA9rEQ3Cof2Tr1WB/+yv+0Wzl9n+ZOY6yMxpYq/NigtWVxlPHte80
0I5ALgm/x8cYluueST0+aBze99OTla1ymd1PK+uaFiI3rlcM/hAHCs4LGhRWV51/
i2Wk6wAJWMEHIVDwR0e6khpZZ8EFhgjmlgN4yXWkNfLPFxP88B2/6BDICnVn9wZx
KMeYxJPAfAuGLktNNYy+L157SSyZl58Mq2wOHvuOM1ZzraAX5b9Nv8ii1AKPi0/H
SGpvRkbZihy7ZH/oUMYlhBknv/sWuHnJuSeezFDx9dfhU/0+S2+etNzUd/wmvyeK
BKV8AisHrNgyX4x6GpYsrSX/JlXszn6e22J2qT9ksBDgArchFzi2rjNDcP3Qf4Eh
CKZJ/Z++xrULRLIkXyiWtfa6rvf9sjq4jox0L1hMri+kZKJE3vak7Cb98t//Jz2X
AZ6kaRrDURNkqB6Tzp82KSwENzQspv0lJObSnQ5WdGkiPeO1Ndy/sby9xoipDU0D
TuZB/gc38e0y2dyjq6N0ZlwEtibQWsZX6CqwONZmwurwhrdXr4kKcfsQyxmnNN6M
7zThi1k6kHj70iDxg/v8bLdNvYHugSl6S55j7k1H47b+FS+7QbDuPB2CV0tznU3A
Ng2xiBEfUP9G6JlqxD+C1xliyoR7VbhcPgWheDBS9NqbONt1zOLFBYatOMpula9r
fQyufr7L1wrU2gvuNHA283ioykwIS6fkQAi8yT/LegHmejxbdQktocvYwXWGkVsN
kLkW6Q57kUGVqdq8Bpfmwr9HjWN2BFwa1g79487Um1zfu3bq41HRs+fvHSHKIBES
DqHpODa9wpV5HYk5vVr5uvbJYSK07R/DDjvaJgvvLEQ=
`protect END_PROTECTED
