`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x/TbZReHN4AkQZmOi9zEPS7obRNvjFyHnW7PMpSZxiyAwj+z6yMCdin4VCViFPVw
Z9AOx4QErrm7Ay8OIXg+EKzUTs6ZkSK9Bt2fDXc9qqnE372MAEjMQhl0L96w3HBk
PM2v5Lk6zVVHY5jQl7MR5jClKNPfYRes3FkXDqxKzz55kDUdos/Odlgc7nCa3jUn
rmDnQrJbDY22MufiGVhdJz3GlhmvUx1+Utev1uBwBSPwAt+3l9akVDzunKXddbQ1
0GQUVVH8Q7ocGmFQWnK/85qVdikGOnT63NtjMdDfPg2BCM4oyHJHg1ilJb39Xl38
ihka/eOlwifHENp18VLLycwnnK+t+bEo4B3hoZTNbUgcN7kac3byDEW8mI4py2w3
v2jEEX5hugA+a4PlSQx8tvGok5r5xs6imfsddiLGuvw2DttPHdFXGmHLp0WpYacg
Kbtvt/ltdcI811UED8PlNKfBDlVv7wskGi9j9+Fb8hQf/vJ21Ucv3tzz/xyJDNY9
Y3lZ21qjTyK2+OUMRw83OtVUuUXzabuL1ONWG6oQtk7htQtyhaamzbIsZLG/Aeg1
auNDyiOw5tXM/i9mDLivZCXsUeoIkIAbtpooMBSPINA3LGDanZgJ3HcrHmsUfRPs
7QNZ24OBKmWSPMHCQf8fq9sL/v9AahiNwxdCVfNNFX+ADC3wPezZ1Q6RB1JcR8tu
MqK5ijo3dRD3QB13K/1x9S6qOufRorZoBcDJxdje06cHeC0m/2I3XwT5+ibFcFkt
akFV54hfSSrDFNgOYDDyx5GLDhd/FSDoPDijmUG52edqyb8UvHOk5UpKFvzmP5rJ
uucZHggDgnXoPUXvZmELA/x19w6H9NYFyr5qh825Enhz1Suji2ZifT2XphP9WOqK
T+PrMQKV5KmWXE75LkSlYrSutkVFJznyQh/IcPaR6LuuNfGOMb9jCzpQEQIVb76u
HTlFWrtxa8vN0GseohKlLiDRJKd/aIHvCge/KIbjkXltgVNlM8lqFC10oXfcXc1n
UezWpRadU7KGPTmrmaH+NXidRvSrnu2OwRTlaOqTRGzpdFmPsTmQLoO9dppLPX9T
jb5r+c4W9xLA/K943iOyy+cjQbAKY76TBGX+6mlOdmDbE0fEHGPQWTeHT3dFz0gn
4PuXz33H5AS3xrRekNRJ0Bet613OO8EVmmpKFRdpivL6m67s6uoEHYML+q1nCIJk
cg4kORicikpISq0EOdOtxg==
`protect END_PROTECTED
