`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yDeovhec4xL4VKqEOqg7Z4sAjL/INkT4lodnHv5khA9BW0fzWbKuIYfC9HKCK29S
TJbRM1HGk0PIJnwG9ZUh0RpWjcVQa/gTh2BIIyuRlelM8wRMOa1hjO+X3ez66uVc
Ca+AzV3dPHsLCEjsokdsHz0VARgZXDgQPkJOH9AleGemWY38Moo81LsZh4mIr9D0
BCz4RsDUjvJAE0fpvOchPvRGJENv8FHcNZzgZ67WbDNZSBNqF1NV5dk7S+r/A7tu
bvtwnieABsBYhig972n4kOEqhFxCi/KIbOihRL4M8gz9ubVew5OfCK1RpI2gTtlU
+nVHbfx/DxVnQuPf0vJLoI7GrMoRQTte8svK74HPPlBImxkCy7yHBgEN3f1SJLUX
FAOxkhiLOdL2Al71BH250PhM0EpshNqGP7Z1T1FWyA3J8LFW+1oNYK4vACgrMdUo
BqXjC9UqUZrR98Wqp2Ligs+F7SpTUxp35kcljKlIETM1w4oLsxARcaLZ3B7arsH+
CTrr71e7IRx96O72YfKKaG7R5GCOff5CwuV1jV51jDiIJDxixnKkMdYeGzNwEsry
BoTprWxHDhkJnzZ8k9sJyafORL4HGL2g2gx5ZpDbgkRhx1UJ92L33+DQ3Lf8V4Dv
5f5kAXCewctBSO4FLLtHr/jk7XaZj4uq5Zq1B875SF+PULOfSPrhM6/aGX5spidu
Jh2Pi46gYEdpap30LEi5nUU7Cg7MjSyWk0xE1D7sv64uMHuTvo/wQtKYlhYiPU94
IpYgQtoArY6wmUH6XbMNvMfvu2/RtKA64I6zHS8oQRmd7Ike6dAWtXH/RlI7w6z8
8u7qMyFsCXJx14IsbOpaj8AMWrih5KtO4zVpYDHmExmkHUSKl8amZHGt0zUACe86
CiQ84I3hEh7W++jGpCwKkEbk6D81vfXd8j1LlcEZSuwaCmOcsFV/ZrbaWBeZUftJ
3nri+epdLLRgGjzsIEYMQaxvRDb3HVeJTeD+efwJWiYFFCGv/4lehbzttYZO83DM
sCx1UlRQ0bxB3Y0EIs9R7umfPe3lVtzXy41E8Eyoj6nBLXfYYw24ESPiMe0MKgd6
njd1rWXI2mh7l3fDjnzGKM9YPKigEXmmI8gSFzTY3NWEHmDYvNoViDO9up3aJ5Ee
kfCGXF07q+ayJmE/MgBEtQ==
`protect END_PROTECTED
