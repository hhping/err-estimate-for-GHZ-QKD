`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SF5X6kFPGIBIPlYFQQKmY5uciFaTs3C202lzN+YlWCBYhVkdhzCjvx/gD3aoOSvy
EOQakB3cogZAXXeRf8REfV2ktOi5tcXVzJGRCLkTICdJasmHDvYf0/o+x+/D5CWe
yWkYFwUoQ6K/tYPllFM3KqHZRN01PKUI1TKNlRt5l5jlvaOjTO33FNa6bRN5ndyL
VQrZLng4RRkcXZrkFoH8Z3n9PkAmPdC6YtYGeXI3dbMy8BWlHfR+zZlSLgJN7j8v
j+K/ca+9JN5Rd90keGyRF2XOOj1kCz+4jlRxNFOInVYSjFRxIj5p+xFG3nlyOq+J
C/cNfkT9JVwbARfo26DfqVoIFA68znsHttS78/BDOxRDCzN8gDPlZN+vUE+up3H6
hHyejFX90a0YB5Jgbv4GMQ2zxnX9Ex6BwZnTCGLe+9Kz94G+DGCckN6lWQ1qsKAq
HQCahc12oj/efxrV8TyW5Z1pDYLKdEhioTpV2kxS3MBJlJdVUEkzifWa7pMRvES5
Euy1KKJ6iyVsR42FbgwuBFLKhLLQJbIWsgJ15z2CAOsjNusLon9ojEqX+j64MncN
jJOGPydDycSL/lfHveGBIBcd1wHecWjz5tiIHdyAAUlAkYcoB5P8Vq/TKrNSTawR
1BuesK/cfO8fqmZwIoqwrr873H88v7p5t3iCZUuc4M+kkc9s8wOCyKzstaczVJo0
bce/obH3QhXsc19Fa3q86d9TvQxDDopBQvCQ7Z9HqMKsdM9/1dMFJ/vXXkumiD1S
ogllUcnVi4tNPjF63gYm1s/1sqUZ44scJRTf5YhfRMQhylKgucqvbuNXn44vCCtG
TwW4epUAO3UBlzIbrGwB0/MZHaUEJ5h9pVLf8oE7jYCx0d3MSAidiY+2kqDqEVMr
T+htvKAzc079wL1mumf/mq+Ons+0uVjRoFNHGn3zDGSvtNVCTtJpyVMW32G8AqcP
uwBL6Ek9fSd+SQ79COR0xQYtd3VDJFszWEwdr3RQAsZ0lvw+zMj92lD3UfCQCFXd
UxJx1wq2t8GdMK8CBcocAUU2HDDLcSkt/svGVpZhvddWl6oFuY6BGrlTapR5K8fV
Pe3zdrQ90I9iHif194UXDRUbUZ0+I3D/6DsfEWxmAdvlLSrAbKWNt36QMRS68MRe
eiKZO9cb2ndx+km83NMhRuR7IQdyQcK8XPOOkaVtdHRWnzYitikQzp5Ea76Dgmlg
RXb50LUScusmKu17z/F/lA7vXJdCrT0BElobOywcdfCyUKrIePD0XX660rOKG+UQ
ypyhatCsh0ehRh+e4rUEp1hCKmnTA+ji01m1rRHasyDbJFgv6Ml+5hjOWTk75K/V
OZ2IZNZWmGmns7D8BVh2tGHHM4TKVmfjPV5d75uIHpM=
`protect END_PROTECTED
