`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xYeb8mLD6sidxAORRXYDkfYcgfX/VuSRS667CBNmj7fnHwMWc2zkt7UhzB/xnWBw
0+Xxw4CTfVCv3Fh3xaGg0VghCrEnZnu7igVsPFT09nvx9cq+DvmUyQmFghb4aVHA
I0CI3S77Hg/qaiiiKA2urOdfKGW/7h9rO3YxF+yVOY4cL7UH8UR+shRiHPgM0ycX
iS7ox4TU8vYVSjyeU4i0eBJaMPoYKzxokmeOVtejGr1zRG03UkU+Ah7ka+GkXosI
b8ZdeRtQqTVQjYchoPicsxhPDgNjTMafeeVXjpp3Bm5+Hp5Tg+nxCQp6BwGtfyVA
JnZKqezIMt16/8EqT1yrBY6bYewl/WYFAeY7rGJz22RveBti9aUPLed6I/E3ScFj
WSh5foUBJOh8KwY8zi3ozMs3wYIOcloeOygZ7VlHYECNf76/LkkZd729U1ydsfDG
uJ10ECi2GJiS0W5QamPSbcNLOEBrfSD08dzkfV+AvuLSrBve1UTXuGDLyHottkxh
7h8xwFQVfNYVqKq1KlX222g1cfCo3MVIVgQcG14SoBCaPLbkKQ16cRBnORXsN4+f
OEIcJtaOqdCgZVDOG5fY6wIUY3YhfBT9TTORc7DU9KopOP894MokcvLrdNqbOaYP
kZOosygdsNnccOnVMtzBJqxamLO23cBrTLeBF0WAS2wNdLbmwiLyI95ms/0NgwYz
UuRsxDvdVSuPrNKIirnlRQulefpHi5x86dNA1BoW19sPz3/cyWlkMSCMwgLgBEjH
Qr+VoGRNRXAGDURkoS0UlErbuFnTZCIKjkYLIb6y4Oq9/AL1EwfV+u679oIQZFCr
Gj2dCW4IVM7jhCnT7nh8oJpKFwfzA15vsHqYdYb5olKkyzrN3vaPj/pbsOzf9BIW
dcJSHFVmV/ZnvGQRtCOXhoXGq/ZxWolwFmns3edptFGRBC+T3IwG771Kiu7nfKxj
2bTJNxASBpsLq0ySbYOVyvn8ytVke3fTNWy9wHENZOe7LLoTGkOTvz3SeQ2adwX3
CNTh+heC7O6OfgoWTdEBnGwAbjUHRCrvMYJ7GoHnjyfVMWggC9IKPdMLN0W5Vw1F
FAVqmpPXxC+IrTFwvDDZJwd+GUFwYV8lgYMAwB5VbBKvvnhxUZc4IE35qhPGVlCQ
S+a45sgjttEyFREJB7sSPkZ5tfWBQFE3AwfM/J/B0M6T7P4U1v/CI7Cw+JkNaW2+
2WBgVf5LvZ2C/NE78mPRS8RUC+zd3fbXv4cjl/oQfov23ThUaTnftkpFFW5RTILu
VAFfHfsiJnT+CWK7B+/8TgEcLNcO/5Sr+PcIWMVdapYbsJoRYswuTwP8VHDTeQVc
qRUEzUXyj07DhqbLDe2m+kyMPFM8SyRtp0ghZFF8RFk3NIc+wuAcB8z2trX8wCp0
IHOvLOQ+uxnYxUcjiZWAi3IVP+9E/vrhqLZOOj/gQvGti70qZcwt/LR/R6IweUMD
ythtVLeg5HTW6Wl13KnBq1pmUEd/V7rKgTYIQs9HT5TshV80sXEVzFT5Ti5954sz
k7mLhlMBJM3K30sEfjSllkhR8dV26YqLv5djFgaamcmEhd/LDQoPYb91kpKjkUrQ
W4yehHkNsTCosngiRt4u4HmjFFJgZb2P9wwTNF2grYrSnf72Kcq9R7Vcc5QC+asD
WHRFxnJOnbEUUck/9sBNCHkJgv0DpRszncpGIWBl+gzeIdrMKNjPAaFRNbCuFr2p
LQTfxP6kuBwZGC4lNh2kr2SpgbiPFRpKoAxOl1S1He5LCwcgmL8ey68uUUwHNreC
etKRUZ5QfxRDZ+r5fVqrgYRmrNIvQL5PgdHvZ5jrc6uAxa2lxTwQRYP9do1pp+Tt
O8FpLd4PT9g5UcBrAL4q0O4kYNTASQl/FBLbDZFBzOwS08HbMhRaZuezms+rSW02
Y1ecIHIGZ2RCPfwzebJlXaM7G/YsGha1hTkUGTdB1kvmGFxg5h2cnCiqDrAU/Qwn
UJ9DUCgKpAunivNIbuOtTZhfDl/wVzniK9zSxnEMMvo7GPSw4G7Kxd4T6AFcMynv
q7mx5WSH5vzL19sOdKwPFeKpktUNoDLUJDFQ2650BeLPZ3X5Yz3+coxJWvrhRwDM
9viM/SZUJVCjk/b2HH+hWWOwyoxpSzsRNomzj3TNODdbLMPfYQmNj7gvY42DRUFf
h9lkb7BgJXJkFC5d6lzo/VaorkT9yPfiAD1sY/9AKIuC5WDVR3cYkkUisSJjSq8C
nLUP91vxcqBud9TiVExWtOMLl1CJIOlbFQYGP75dVM3MJ5NWAtCkZpGgmUPfqNAI
WIft036/HDoB+e4vQxnUvmRVJr0t0BTFy4htQ4JPQ4PLFDETIioXFNXU5WreASz9
+Iy+WtnjBZ8NMLf3ObKZer9Tar8rjI9RCGGvTl3jHcewIgrgmepr7NDjshhYYj35
jkmfpSgxd+qJ9A+ahcas3iLAaCSKXktPdbqbr96A8W4Mj6BPGHM5MMuj7x/VKzNQ
uHPXbr+tDRW0A5R4u5YqdGZyh555rEPYsPy0hGqSYmzAqPU/WeCg4/Gc+Oi0zqS1
woFR6Zp7GYOMuP89o+wn/HtDpvY+UTRigso/ur4NzCRwPZGshk4rwG10zp1jdO9n
Q/50tPk7w6/vnVLu9oeqc0mFJ+Y7fqaKO03ZiB2+E0VVOG1jky0dhV2jeUILyU8N
W5eS9bKFx4G64wfMUCpW8lYXMIiXxLgAsg5xLAxETGWtaKxhXyOuwb+86KdUrVPK
dKog5YGMExo8zfr/YLltzIvXFrVAa2qAXP7A4BM6cCQWnZY2csioxQD/Qgkkz4x3
hCxt2FjUwT+ochhvM7DqaYu2PptFdGkcd9Y/KUYV+zwO6ULo+qRxmR2BeSk2Kzjz
OiLU8d31gl0QRPwu8U8BYd/bjknLaEm+nx/P9wspHCXGEn5HIvJj9YnR3cBHWL23
8RmnEyCsu9aro2nbTtjbYr6H+/RvQbuNPtKr2a02Bpr+txaNEexOi3BhzSmTBlwh
23idpa16wzSYF9euSrbrH0AI/5nC1im7D7s+KDW5NlXX5IfDp3xIfwJS4zYZvipP
ebdQhFZ0s/bIJkny0YXnu3izVIZTXMVskpF/DJoGYE1Pd67QceoG+gGf/WdzbUM8
oPYRWhpDOkkLNt4sknO2ibWceY1V/o4OkPcGbd6Z74WNwDw7brgtoK/jXqSeFBS/
/T6aoWkUtQ0xHzmcXUZiW7T6Qm9E2Gm7WrEsG18P6F4HWe1/MvTYxM/mtkUlMu3G
5ya/GH1BjY/A3yYn/lfHDEMq0g4Te1NNi2kK9zSN1J0FnOVG7uPXJsFdW4DPq3E0
vXrAOHRF1EWkm/A1BrPp0ziedvoSUAH9wiQ/x+lVKHl7NvgBkSAdgIMYiPT+y6q3
K6xvqVDox1MW0gcnePm+OVLUVKS97h0MefvJhsf4wVyx/R1Vpm4Zl1eNbro53awy
io0tlYkjF0To+a/BmeVotZk2IhQnHU93Bt0lvVkxBrtngVPTcjkBEzrEJRYS1wUw
3t9CshRXuhJ5DlCxjGtV6YMHSnL6Nj9LqviUMvjNK3+wAaSPSZe5IpxneyQw3UDm
dl6tGwaLE+5ee07EIGw5PxGH8uuClrGQ+gYIquEQInuYrexJuKHKniqZ3RG7n9UF
5tTKjQvq30V31xKPCMC2mWagfGszGr9nkJ98CdP3m1GpyFsxsui7s+UAIQblQxwm
dTS4FEE8f9fYnJnb7fqX2IbWtt7drAHZZiXWjM3pKV32HA2eElZxeOH9Cu4B4jgl
c/5LPVF95PSpGW7ffMwDX3NE3/CX/Zg9P2ZjaOr7SF5H+JSnlTyRj7rsqRpXwJOD
APPjLkVKGgxW0Ws5Nc8Vb7vTMh37CwPUfCjchIF5WIxNIY3mJ5qk3/jecoTCMr2F
RM6tEb83DUl7emhJ6+ZS8rC1klGIFzUGPgwYe/0ZCF9TY7TZxmfVDMp1r76bQO32
vPW/RLhDK8b56rTfB69UMef1NKrNF3dYkmcHnIuGmd/fzkP03I2398aLXGmhAnXL
8OEJxL3Kn3JAGoARYCN/qMtzW58yFkzjJh3kfW/tqUBxtLADdGv8V/VMUMlEUZAY
yo6/dHQ98a3sDzfU9jI9dQ61w5O8s4ixtXO3A7sE8VJiIUNUrtrgKJzv2LmOG8HH
RUvy1ZS+P2b0A9KS6HKnpGktMKIZUAwHGTeGsse93oxtDA0FYf34JXvypcduLfj3
vaEf6ZWDvIlU4VqFyMuDRsGkNtaezmcWCPJL8j+qm/LlG+kn3gL0Z+IHDCIwPaVo
jnxdksuJ86bTv2/MjhItQRyFUYz/MwI0Rd5cMVKOWuRYJQEaYBXts2nhmymlpvg6
jRlTGyMSNslX3ebNOBxXYeU2CP87k6xqpvOriI7DPBlBPSr0+XHnWjIkGvYGuTBT
gejWGcGcplyR4gNHMWOhEl1tif706mofvfAoVRq0TLRiteqGzhTgvXmqv+AVjumL
pXkoi7yEzyhVCp6PnIk+medYq/jmKkb41VmaTJPo1+wLml0CWUs4im8rZa2jv3Tg
wE2iXtpx5DbbDvn8JZoA5XTvp6klZGeROLxP29N3hr063SgVqzXV2icdn0KGU0ds
XTk2ra3yrlI6jpKEa+qAu7bgSKjIpAnLqCElAOpPzrZK4QbonvJlsK7Z38S3MvKN
k7e+bS5EWO4LlIbAX4AxHzEI0wqjMhcl19bTZhnh4XfVInBIgAqMH/i1147YTGZS
tjW8/p4ohMajxZe3jJJNRwUIWOBPmhPTiGrXmUntWDcpi3k8fznff/jjZM5NN2tH
5pX3YOao7H+la7Bn4APmhAAnHywlEjptzk/knu9pgbK0pYnRaBUZNSL5WVpen7WI
gB7g4uuqetfwwimIpebX4H/oqxv+RN7+Z/qTXSpxBitc2mZNhTOkE8/utHBPa+sY
vYeoyIaOs6cTONAm+Pl/kPgfH0H9M/a7KxUj73rBOVieTnm7J7SCm+RswIum3Urx
Uaddanrn63v6NWPWu9HERn9DNBQqeFXzye1V4URCbHr3kjLYZtvFaIBF4tTssHse
SPFKjh6HwylAsL82dPH3VTYGfUY4xdkrihFmATggPP38BvaMTP9Qzyb39wTE/TVr
Y7Q3/Wci/CboFDKXl8dlhMpqvpHCsgAlYh8grZ+DBDeokBYCzUEUAyGYRQcvgnl7
+CFIBwbAgJPYCXOlmLqHvKZbFyJmOCvIxQS/SAjYN9m63/J85CqS8HIEpMkeXJFN
4UHeuxt9MwiitGUMTdHbcZiQp983WIxALBIUB0WwVotQqQ/3TEqdm5zyi4imFvwh
b3qrAk8VxvxgEXwh5gTGfep6CErH4M5lIBEe67TR5p4EErwCK8mKf9Pp2vtcU0n5
JkOGMkhuUDTixA1M1bcp4FN8hvvRaPqoVsJ0xj8gu9OyqKzOOO1tY2rfiaV1VRyS
vpdaSo1vDdy64MikuWce3CtLrbReNb11ZZPFNz09DVMyDOMwvHYYLsdzI6RUNcnL
zBWZh6HyP6S2o672BG5qpsujo2KZGVHTBWyow9/Bpp2tvWJxkyjxbLeGvZL1mCtU
45kvY2W/RetKLyCCHtQBGsUeP0nPpu77l72KD9gIetJvvs8+FVeAbdUoDD5OWmcx
rpDjpsUBdrToMhesR8MQyxLX4zePE5Ts29+W4l6uBb7d8PYqmoTqUl7Qvr9yVHCl
Q0oz2r7HEdI0puU3FLmkcJCpzwwz/cNu2t/MN6HYf9nRUisLC7Ib2yDbz4iR8G0m
2L32AjnRgrbKQFl5mbYjkE6dqbfciIcRomMzdzlcWFolW6DHf03WTzMAyIhQb5nB
8lgLUjzmG5X9e5caZTLyXmCYPzLKh4QCC2r8GUvpOxtP5pliRtPnUj6PzBom66kE
hD44uAWYLGURQcfo+J9E1qTNphaCeVqWSm9zk+AJksS9iiutOn+vcrjkx+/pLv0G
TYWrvKMQvDNTJ1TH1JPD1QirZM9IjChstmHOIlkgoEDFjPFUpxL4ZV7O9GFskv01
Qu4FtUmdHoGUEzfFUkdZ0DxVeLcF6dbFVdPgjKIVytWcWEWLC/Z3FzCvuo+1VQ3b
gufdHIn4sgrqSoPcU800GPcsxJB4Ycj9+7ZSmB0iXHmAZT75v/+FFAfD/6GxfjZ3
a8gK0eHQssrRi3Auh7x8O3fc+W29M6Vas0mv3r6iGGzxkkHpMPRV7hX+HvPBWC8I
dqhPkIl4nWupUxXP5ILkeYePtIbFORHkipgQ+zhvMKj5oVXC2fp52MQ+039OT+mm
G5u4qwk6rPQxoUW6OdoHBaClY8b1iDF+T+fNcn2zsLOKU7cQg7BtrpCEjZJEGt1R
cuC1jhXBOkexqw1KzAyawQ0IadFW0DyDkvoewstm6opoYDktfOcc7tpsYnBLlRrJ
eU4tbV+B03nglofEU1cLRN7yU1yzWxC2nvuLogZNRCBF/naurXSD0zCHCdVGVfM9
AWM6WZFdsK0OO51roHOVNBh8A4oWoV1Ro2PJMFEiV3ZtV1dq3pZOBGMF0VEB5TWm
lNxzeaicl8EPuzFxcbgRQG7GQY8C4hqSuYd0R2en0UJbj27NG1hudubcI4nIoza8
G1Q4VeP570J8tcmxMc/NoHoCJP7SI7c18isvOxNnjnQVkHjI/LZ4qjt+i6tzXS78
hT/bg3Tvech4RQejp4ooxpA3F+6krGpfdhSvn/Rq1q2fVuyFOLxZZPK82KWCpKQ8
hPUQF+GsnQk4mD4xMJk2amR9S1L+GA70hoJ3dm/bst1+X27ClK6VpuRjUb6jvF2X
jJzYiMORlqcVuoV0qPBFzhP3RuBvkd2pcdxRn5BxldV1QcysGNkX9PKf9q8ozxHm
b39ZA2LKDZmF7eVOG1sSoaekwMSaXnw2lApOQXAitHPc69tRWBb0+9OFUqHODOLF
xl1rKA9rULtHHOdf1+qZcd4RM0Ygvn8DX8WmTcAk+BApQXQfI4svFeuAlcWJZ6Xe
a3xFszl6rXaZN5Dcjwi3WNgcnjp5LqfDbltiN0C6MkFus2zCOnVptr0tO5tvPLx1
9ZVgitu3m/1+TlnnhPvzn5t+yBxrIbCyZOXRbS78kuBEFlH38aF6h0wK7ygASrz7
3FxDDpNGduhxMujIprlwaOu8TUKynZOwqxUf3ZI89GBJz5dKtLAU+7SZGqH0TySC
UAugYxiQV4ZLVy9KLI0450uBdtdixzl56Isi27O0ZM+Z/vabzXiHmxQpKLfTfx/6
RHdYkIrAylppIaeJnkm+b5TSMbRqyiTzKvcHkLeH55jrzc7ZBe0bINkBnynOOQfJ
i10WRB4P2OvJg8bTJwTDKZABSkN8z9tP/vHh3IBWUdvA6AtBGn/bOHtj11rRSYII
RyQf09itzSyli/Zp+EoXzOOUIzSuXP+v2Re69dPx61ysKdthaheWhJmIAe2zGeWW
ia3/QDbWzOD6SvHKNcm6OAGnHfgKmhWxm5eIgBgU7qif1VRFf9jXKSMrlXTPQYCn
HF7f/AcqPLxKtzw/DPytEaKEmwlzeHQcyQRxksw9BDLqAt347HVH0y5HJYFeLN/q
EALzw9JJiyIANgFs8/52wlUxRVbVGqrF/VNpvSo+GDRSeuKFNHxyG7wclN9FT7nw
KEsEG50DluNtu7CRPziopSPlThdNnua2I27ksX2zJnnh3D6jvHD7sIg6EsgN6tVN
fuOgl/QxpbN2Jkeu36m5s0Kd3kXiYOnznF0yjpxHVmUZviTB6sSNwp+zD/0OwHHs
b9bE+3pwpS5vyf5WH2mm/Y7YHzRWae0ChfVv6FgHpEayIT/5O6Uq1Geas9fok1ab
XLunDaIYhE2KR5FCnORbUiP9l1cNvEeUXUKML4Wm24AYNb8hV87ndGrPjsbv57+t
qZwGem1IK6DpjxKiI8Yv5W9Y2i6EVO3T2n7Mz75Cgrn+4iRKq0HijvgqfsZ4XKIY
INXuxE0O42Ua4nL1LhuRHdiqaV7qa94LZ70GRRXq+2TmwVUOTA1Ch8llMcQFpDhQ
SyDrLJYJ16mLqpjuWcC8cAbTi5/ZlBRTN/wBOya1AapEBDjTQCDzI45OPBri7njQ
sXiBX2iUnk+zgG3Uxy4ZppFi8nQoLtfwDBYFITLL8S5sQDZWRwrZDGwW9e4ERFOB
IVEgyWQsFHDZIYJ/cVB6kbEv967RoU42hZw/yQfO06BlYH+jxpsnY7P99EsM+kVl
Ib/27NMshkdYMUir4Lbjr0amXThbpKc3c3rWx20MdoKWVcn0jl4qNr7L9DVRQm9G
HZEgWwCi3I0mQmRrNb5icxlTHSHfn7vXSkKT8IbL/wXW+un/YP59yNnYIefpzIrC
aMYs1l1K2xnWNidB6tj7FWmwQycfLlfRhE2n5S1EpYXQbvYsF0eAKR5BSV7AWIW+
GbMS8Uh2LBGc71E46LrzakNHHbA8K6QQqnAkEoHIEM1Vvrv5R7+cWPfL2DWOt8hp
RluoexaOPt4K354FBPb0wBWOrpHe4rpIbWWqCADMZJsYSDvSr1MFITpeLrnBIsUF
WOyk1Vg5YcGPccNDDISYbCY124e0nMebYWjkihMPbe+wc/HLS3mLhdP/rOMFQFlb
4r7JINqBMVqvPhxK5PAcC3kxLBXiNWMLS0vOnd54pF+ep63r6SuQCGGOjIfWszoK
gnfheatpF6canbENznbBZAek/3/LmxxcoLkXmMPcit+lw/gNrUyibhPiNu2cAqmt
NF/tcL6HnW3GMpkErOVQ+y8VuWyBifCg8dFVwvP+3Fke9m3LiDEYr8pC+L9YS4xa
Nze7BgI8OUvE+4GQN/xq89E8Rzryhbv8HISQTJTSjf/HQd+3Nw2qru7yXjcBoX9H
CMA69f6HDwuRPFXUtaOJhwaMkDuh2CFUjXW5rwnFHlpOpBC5K2PFd7bNPDCctsmY
94aIqlUNcCBwB4Csgnd99hTJN5fcGrXbRUNdYSPia2Dk/MvuKjpDj68OAk51WWb3
HVm659CW2CSXlbhF2ZzQFKsYEWSbwDLAfOk0X8ldA5zf60Rz3C+WZZVpaAW7sgrL
0vReGzFgo6ofUWe/9OjCH98o2MNRBpKqHHlrplYJHS0mRnrF7nPMUBFkcfXXPygT
KbnCbb6OW0GnJH4sNRRoFX1rhi+jvGYcmg3ZJ9EbjXEkVZ+YXE4yHvdwOKkDho97
RIurZTltbKYKFGXrI9mj/bK/t5nMef33m/fwBGeAZVqmedJphdln3p2/v0tw+S6l
t/4keDf/iDzUPVuPbA6FMmsOVKZMhRM8I0EzbhJyEQunK+46w6t7OW/r5iBG6S3H
ywUODvBqsoHc60UoO5WExcXSqxIvXHC0kQZ/ShuVIH4QrZOmLy7HmiLoerColZiQ
P8LFcnYTB3eyK3v4lrwQ9NvGG42Wf/X6G8OZxhQf7F0wKGkJ82lPJa3kaMRXsbeD
Cfpk7RJpan+vEIyuPQaRBWoY7nHijrm1Wpp9Jxcr4H+/9Tj6oB5kbaWe9ds9+q/x
LhJ5yx2Lr0FaGIqgGZcl2kP41DFQrG/Cla7ppHIyjHu9PhvVkhrCeKP29ENt1LY4
8zc3hWqvr/fWWSiY2TrOt8SNBCYs23ZZ24WcDpd6XVUyoOXe5W7VI9CP3Fe2CRUf
e51uqjrv8Rs2hCzi3BJTJvj/fzw3U8ohBce3M/ei3CpUhdzlq7SH+Y1yWEYyvehn
6+GG0h8vKzWUnr+dZHKZyxqMJK2knTqEKvbq2iFCI0w6UEGfoFB2bivqxFqxLFDM
UCEjuKtRSCalVC9JPtvdE8g8TMnxIfn0KkxIRCZI++FR7Ispyt468hfVld3XqQrZ
T6P6rOjzdS77VitFmJf8gisKvP95T+iluLgSlwsmMni0Vd2vzJirf+whNa+2Y9w8
LHI3QvqVU6jKAfVzlmkLS78xHEyWXka+Jo/kYiVTh2RXXXklbsKjxjX0fF0Q2e+/
OD7cjMQN+4cyCW0cq4A8/9COy66OYVgB3YuxV+SNnZhj7wdABebJb7T6bojOOMDw
5gumVPEeML++QGC+eFWtp8JxvqfMtUDknSpCcRKihEtb39/FnGOlldEOvsVB7C6b
ka7avEH7LM/MZlIBUDxye5+QiG/5ye1MjHEhFpdv6r5STgxukpSrbaWy3V+i4J+3
3UPl8z+S7khwEylzKwogWWM991TcuDXqXRBoLjT3XuzNol4iyavFcePUHphDFkfB
jiFZ7DMGJ19D9Gih0w8NsN87e/TTGgwDMPNhjx+gabWiboYbQ0KwJM8R04iXubFR
Sp+1NS3bMDn12AJ9GpN2NDBEcJTikNFQP6a8vrbbylzAckb6jPo5/lPechx9G4d4
vgRkLD7hdvu+6isaE4TQ8kbiN0qR2oJ6DJ4D3aUWEJWAW6dQrAPK5OQwDWTg6uVm
dQYd9pMTpRr0R1tN9Z1ouEtdbvG8nB25KnkeseNovpjIpS4wZNmS3v9zjCOZ4KUj
iREYohQUMPduTZ+bb0dXWOLQKzDUeLY3qnCvK3AjZKoycBvkEziwIfTTwh8KSf5G
`protect END_PROTECTED
