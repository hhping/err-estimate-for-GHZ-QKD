`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SJMvDbO/oKAYjeM/p2CpfHRQ+AEGDu+GpV1bpO8kCwKUsnyv7sjbsTkhGDwC33fj
rFtVMJT/PwRaVCYJIdVN5PNJT6Qw4Au4mJwsSNt0vMInk08tS5R9Otvvy1xBY6/H
0qdCJ3653aOtkz6EzKssD3oLa/sEQSwaLd/V5gQslXBWbY70iC1ijrZ7Jo3lM9pN
OLJgXl/35OkWCq5Uu1JVVSDBK73Qh5vyt+QhUMeB3HK0vdQ09FIYVRIZzc7WKRUW
aBK3biRY+bs4CHUYeE+WuPVh4gKLiVxW6WbI46DKqyeU+w+fL15qI4VqSHE4YXzo
2qcrGVlHPxqL6Ob9QJ1vA4O56dsac35blY3Gql1b9vCV9IhB4lOtnGG/PDo4Fuw2
xjeiezl237gw+OqXw56qKMSgiaodxxGRctkBUOmMnApnrgMAUqDKAx13zLQ8q5ux
eZNBYUDP12GnAeLujwXdvuHQqpuNG1Vsg0TqSGJsjcR1BmsAwbi5shQ+1zGMac60
9cBNLJ0M/k6rfaeXIPU34u4Kc04Sh/fp4aRjMaRZULHL6/ILPbIi3fpdTb8kKkV3
rJDgyBqrp9SlUEwATtZvP/6jDJIQxoBpcVx+jSL45b4lnnWQx0itTXOQE8jjExGA
NtR6l2Y6sekXPcHPnWILRAPLY8N8mvcnmGPtZvg3VGoYFsMYRptaqUIa+YADxWfP
9N93tBCrzSa2XaTc5R2J5i7f8ntxAr5esd7e58XqIORK/u092IvAaJzfwVcL0ubn
05enZTs3FmIh+dGydeuji+M0CtOF2iAqRSCKwzswz2RCgscOl7h1Qvih801CLUX2
W5sx2LKXg7R9z/8ih5zBVBG5b3SNWEkuv7VlLwplg4tz5mIpvo4pvvPRnVucAEpN
3TCbZJjmmCdYswmb7erPO6NcXTsYwSlaCFmp7S4JyfURAf2jylTxWWIkaIc5aR6Q
5M1H0NrN9Kaygw5M7K5PGuCK9w1ryQtgqSbS2LPniEsg/Fij3bCjqfKJSTnp9cvH
FFhQCQQ8jTtvLixOtnRw+cI1I7fxHpEqyaswvF3cVpT0ED7fwVhIYMNCyCeenXWw
qSb61DbZvZ6i0HSMVicXhbt6lg+2ih0gBAq22zyAvbkeWUKv6GDDZcekAXrzRc5/
mVbJ1mSHoAC66QcJ0k83kqNB/+1Gtl5+4rUgQ3OLWrshDk2MbBexXihxIsiIapEg
BN0SfMafQGAJUTtJVXR930U8UbXisIuM5SheLalisQPmtHeu2FV/SD9cWpsvmEOF
4VDgT2r7s1Fzp+UK7RAoI9GJW+niCbUaPQwsZzVCYCzKyQr1+3rvVOsLfK/Tp/Lg
YjJWpWg+OGbcBKVU5Hu7if/BhryEtIoVC8GsoFAPSp91t6SfAvHwreOyLuyv6+Yb
pAojtCg1nwHtlxryyGctdCrumwPl3HJbn3gmUfIta9zEhmViG7136X+zo1HUP8IL
4dhzoohfkOk6JIACfedbDTqIFCaY1gc//Tn/ri4gtnK185n5TyRWsLr2nSBJc9x4
b6stV+CU3xMvy7Fn1Q5S6+0J9ELNaLDX7G9FyCKSlIudhHtZ2XcC2mG16+iIokUI
7/F4crWV7jZTcgG9kwdmidhalQyfHcMZ1A2/4IGMP8P3Vue+eQPNMMsIUPi66a48
lBX5qlg/3G7DY8lxnGHxCg==
`protect END_PROTECTED
