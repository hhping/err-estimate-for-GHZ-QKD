`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gco+sfwruQVekNa3+rFJLtTAZbAYSGf4HEtkZzy6/Qg88K2Yv+NGhacOwSndynD/
hxzUjoAzCvfZQYKZn1UfYw69VAJpwB7H/c+yd2bLVVpiAswoU6pPs0vaRGGqMaF2
r3//VdBISWdGs8PRXTdijhhnTAUao7x9tavIhjJTiWLQbCxBxEpnd+yKqLXfWOSl
uWq+tVa6fYTzR92a2XAp3DwuuANCcR3PFtFNbdHm13BAlJpft76rbfvKtuh+3ZdE
uZjEg/aBB3OaXYqoS+aN7FAl8nErqsk47b6iNUxA3i0NOwV/Dq/AIzjc18gYMxu8
GGyNcKrRD9mCmQdYU6A4EfYGNV6/t2ZBQ/Kv2NwYieGMD7RDq8Dd7Q5AfWxhfHKE
ahhqMCccJ4qVINH5+I5KUKMjHQFJcOdWiCRpvUWwgCls3VhpTIihLDiSShHGZ1DE
Ni/HDfmWjQPbb+nNbORB4WEVTwURCX7IpPUITdgMEsenTtatFJmVUazh0Rwkpc3x
n56+nbYjDLh1r7BNB480ECgp4mTAnFtnKpfIkMdDel+Tqg6BJR2OIoqnWmTAu02N
d/4ZNjMZkDRgKmallU+YgMvWnVuG43Z4NXp9KngN8QxJGH+niiFO9S6ADifZAozS
BgMvLOXAyL6alI91J+fpezFfR5FcqjPCwxBK4OvvlllqfPenXSQW1+TynnAB1AUl
/a9y6T+aqW3SmErUpvidMEn/dwaCn/uEtAG2ZxwSilfnqBJ59UxPENa8CQCSZUau
mKbGT6C0lqbiQVYWIC8aCnD9xR4WpLerDDR3CnFQkkyXsAxQTNADmWmu5JSfU4Uj
m74jO8TZzXpCuVDNaRYnoSiZllak6RUdsChTihfjYYoMxgxbSNlligjkRy+x3hqv
hkueFAZSfHvRut7ue7jx6HztLXUW7xGlysEqVEdBD988J1V77czcaiB2W5PhZU9S
ym7QckVyNOAUlZwxdSX3ykgcNLoRs7T9AS7P2MZ3QR3I6hb6yPIdWd9bZxRi4Z3G
XLIy/8nQIPOfuDKxshVm1L/YuNvm3BW0JsTmdFLnUzZC0sF5Ai4JflN9BCKVeVry
S3p9szD5bIuVOQwDy07aP8v5ijDT68vXq7zpt6yclEwr81eBKm1yK2LCXtlfou4M
pCd0qNpIgMPjyzs1iI7/aXUqcG5avCrLiO9aqTytBwPJZ1t66PWHDdd5luSe+muK
mITwCZM/v+EBl8/kJxA7DUd7CvsYHhGtciV4rrS2C9o9uu++jpxMNqGtTdh+mR5r
fAPwXiE8F3deJNSbZJrkxhGvx9hx60qGKoH2o+TzGzHs0GoCVGJ5gZrDSoAPUpiv
PoiOWmc8decY9rwcOEJaLcIT8xq6y1OCyzq6ZIXPQavW2s/9Yv/x1V+PrbubwWCO
2A7frUIbiLAhGJJeKIb+Pn/Bphpej3MFfmIDJbnPyoHIiurTmqxm2tsvMbammBtM
RogQFjYLXH6e6UpiuaoFZe8DVeMso6BC8nuTtdxw+Vv0IBtfEI1gGTkkopo2drYu
v+AkXqwXREuEa9GXq/zuu8PjN6LcC8RgMHjZRD10QQKA9Y7Zky71FAFpTJtxNYgJ
f4rqTcrgpZBeje8rTYMkm9Lat767r66xb0YTFzzHCXsiynxOJZgM0XZa/6P4ikHd
nidODLloCaPO6YWSt6qSJ9PfLhTArJNKMybqyxpyzr16/wa4USxMttSZ+z7sZfuF
EippCGN1Jyob00r5gwzbIkmv5pJNkWLd3bzrKMr1Rn7Tz0lmJCYUgXyD5x1b3LTA
o80fqIykoiVLCOJJ3EbHv9234lszVN3jTRKDeaxaI+wwff9AMx5mZSvYVZ3b/LvB
2AjDJfrfWt47SKeat8JQpAYVPb39tQyyrHuOWWOqWgdwafo7ulkfOcH7J0znaCzj
XcdQU5XE3DyPxIrB/RQehz4Pn7JQN480mPjfu9iiC5PlCgae/Ry7E0RZA7LC1Kpd
+Dsqx8C4uUCUmt5SLZs7lcyHlqsv+iz/M72LXlpsoxt8SiD/p6t3X51VJ94lFPd2
MnIwcAQxSu9v8D62A71zkulhYt5+C3RbVUgInsJF8GNXb/DYHNJ8uqPkM1axxhoj
+gMJKJAD+8oyvWsWeOyCnu/6UVFnaTi8onj7kgd5gQnmr/fs5ODVhCUoppAOp9/7
CjO4oyTHqHs380UiverqsmG4vCM2Rd3tgfMTJkUdHztbboXpSTaSasRtbKI6/F04
78qU10QBdrvaz3IJXPbvS6pOgkDSim2lx/7nPmtm2BvLk03zBmZgy6uHu6V5x0f1
7OpsHrIKnkajuUQ6nlzLDq2gRh2ymvtVQqTO/76FZ0SPWjsd28HR/y9Up15WjNWH
s0UXOYvnqvtw+TihDF+zXUvQRbZfY46ginfXNq2V7DFgcISfEZPTYx/u1k3ubLe9
hyKiJcIRO5nAY0KcJraMZfsS1yYbCxhCjvy5yr08TzJsDVtA8qCL7nA6FZhjmtQK
J5dONzaqJ8/mAT6+GU13dXSwEhST33Nh4L0lNHySZWJOuzfl4XqVt1hJg2p+vW5h
x7FhSUmMDIbGQza30PtMddTPSko1gV7GKVkKvbSjrP2KD0D0KKIf1wWWSEa5FLn3
LGhdzxRgX4SFt79VKLA1XijMvAJgRBhySK9NZePEdhGqj9I4j9vH3OkVjTx/qXWZ
Udv9iCP/AQtlN72ZCGIKbT4+SApB6QyOkrzzHAl59dTFv/93hT0YZ9k+CHbvEw+t
C1NSQjDyVldn0FQRXVQYFYxA3K4H7qWibZU36M0MiL7UdZK+5EF5GRrqUYptlcwc
TWKduBF5+qWw8u4vFhz4LaQEdxnYusYXVytUlP4S7wU8YS1i1GwFHnM769z6XDgh
DEmvAZmzWtyPQdZzwCrgh7aqfp0/J/wRqEE2ZTKF6gtccw0xRrENC21VxkCLCgq+
IQ9+xht3d/FJZPXcozuuuUBcd/GytOVJWjkgGEZ4wpUybUteZqItAzRmQE5RGuDG
3W681FHoOWW6b2XYw2nKQvFLlb8Q5uxPjlUasp2lQnRNm1Ji2cVA/jaEg7ceeCLe
BX/KhjZpw5NpzxUS8vCCB03mIxMYo3eAkq1YgnJoQN7R/PtZbhSQZJJpKA/B/qkc
TeldJGXxGmwBwt6TuQ3Yht73KagkjuJ5Tx2CSM8Adu877hsIdtOPTOj6/w/FqobF
8bKTajMifGCMPfsa935MUCftYDeWnXgx4x0sq8+fbhKAYMb9CLnCQK670vJVjhPv
uuISdZaSlA1fk3XYO6XPYsqTw4dQA1f3+UMLe0mDquz4k7rNU5dqTz3Ezew+Hhle
51t5oYIUvtQ9hkpBsF4k9TdqKM+pHc5BBxRTGiCmFtyaqNq9m8X7cwrMimuOczbI
J53cbbHorEX3zTdFBKrHnYXxRz4pZarXQBxJ3Le/fKE=
`protect END_PROTECTED
