`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2LywTpRQUwda5CfeUCYfUdFtxc+HfSW5srjeUsuPAOePYddgZDd9MwPWosSJuMMQ
zADp4Z4+e3wZi2QJ/iS+8md6JCji3k+3hJmq/YrXnOtif6mL0zenn268bdWjCtdD
danYGiIInkN209PEsygrC4N1dRux9tFjvmWXZvZe9DRNGOkJBnZRxOVpKI/dTVTX
4Rxewipnm3I74zl8ON7SM+tcRzvN9CG9giKaDLjHF6Vq3kiMUwoJuhfZQfGfClUC
kGFsv3rsuw/NlqpRxw2LKjs7OCGWrv3/zm+Cg2I/SR7/Ny8wPC3l/mSRJVP/81Nn
9MCL9Ls4K1hgisktDp+nZApvXNXozF4hKy4wKn9wGteJSbzALAz+/wL/q/V33y5I
mjY1cbwqyzWKPSj8PybHsFBJGKJh6YTUVn9ySWoqtJY7+fkK7xcJHQR6t2dmSTZ9
dbDDHO6VyDa1NbISIE9l+jcyxsbhO5vCq5R7slnZ4CCOSW7mxVLT27j/ruZ/XIAO
M8oF/iO9JY7qWKZZAHpazB47l3f+nT3FzyYQ1SZ6l7DAX1YLkxm78haPNOhmymki
5OsvXfiyaKrVId7+gJLOUaXcDSbhaL/NdEeZ5/uCeFfYjoE2V32+4o+U+hTWF1BS
bkaB6bpUauXVoIER8oPCfQUsMesuLwyr4OsPvJabYuiG8lf/IUdqVChWnmzOh8Em
Ct5Rrko77DbH2HnB3I9rtkLas+pN4oOvsBswZmE+eLt3VtioWUjfvmAL+X1KzXCJ
AnLM454g2iQ74WC6rrSXAWKZSblP62lxstB6dAPLFzVLQaiMCh+3zuUUz878WzI/
64SZAmvFPfA8GssM5u//9DC3Jv22purl8Al8ZqdwYx+L2xCKOPX9qBoLEAyiQ3/U
Yj6j2G5UPC9QIYUILvRjoxA2RwWcfPglZOKcdQxJaBG6Iv8sZ+nF7fluH1c8GeUt
suICpYeby8MPLkX+quClKPt3hX2Dny+D6vgc4iEgN0HzVi29wIewv6JzfQ3hkcFn
jJedk0XDwU5/Ztrn2y5tEg==
`protect END_PROTECTED
