`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7JkX9U0qwHFZNZcLXC75fX3glisRgbWivq2CA4msztEHfPRMKakGUii7+qmoZuQP
n+WIreoTGuKDvrBqubFHmeLNAaRl7IN0n4ncDWzeRni6G4hHb1ghK29NqOwsvJAE
9coaN1izPfuXr3HUzXlpgYQrf9a0YEMqTbvQ2tcbLOz68hXYKFuMDc2B4mMdt654
a2JjEdFaiykD1XL0Grfd9/vNH2eLCySh9ExIIDBdRef82CrVj5RbGu5qhR70qihj
VqjdBJc+ZWZ1ut8+korxZCo8/lTIejmtBaKT/M993yGJlDMDxjssYG47xu/DaLM+
xfhK1uz25RQ3OTQoa6uWcMqKGlGTmoLCWXS/ZRUcadL7I/egD53MJb3n0Taxo++s
VM7MoQxvgwGHvCJsxmDi2sAC6TTit6BPDOh21ti9d4/ScD2+SkHBLeEBdqUYDlkQ
yaWpROv4uzxgNOOszeXUKqMVM/pS9LN+cm2fc+Q9Mz3+JtZfsgTFF+M41pFJW/zC
cGm4tTLnAvjAZ0Wa/VTMJA/sWbJYVemKJYxet73LC1ht9TksyY5tIgtD1bVXvti/
mBW+ynuARxfqG1/WpVtzL9y9v6UymrGU7hi2sSk+fNwfNcjZOImKNZ3i6Ep3p76P
Qhv1jVp3EyDsu77/u6yyNMIZawG13bc+7s3L9yNEZZTdD911tcqM04lsp8Vzq/WJ
XxpLa1LXAtF91UUbiqseiDRWE1HnV66wBM9Z1ZgRCYK5BzsheJatPrzZm+md8gVi
Lv0XdglEOIggznJdF9FNRUjZYFONtP0esNiJl7FVH9qTGzk72q6YGSip3qtNCCbm
Ee0GkXAoLImZq70wUlcT9ytureBy252vkldXguA7ZbJaJnvRh1DyPW3oXgEeDH3o
yaGJIfaDZAH9xBvoyftVJ8wSbGNxMEtp3M4nrUKbjcVPmCjghIBU+eHD5NUkTtwZ
0EM0Y2/Te3jOj6KOThrJnd60CIR05FzzQLkOqMBgnSZxcRIZlzVoIXZ44gfulJjU
fFskAKDFCh8tGoDAkrj1VS/1M/bcDLFOveW/iTy2QQALXD2TNplBkfiXKd0XJSXV
VZkohanBc9XXsB62s6hRBupuVRqbBUAkGrqueM5Jjuz6HwTIvCtbR2n8PwxiMzoW
EFi4a+ovp5F5tmjnz954BU1t6Qgj4eKakLGPrv7dVRKGEn7BLtUxJDvYZ5c2lUw1
zGZfh+mpdC5IzyNBQMProymJVDZgZNRYCCZ0ZcbZxFS4a0HiW42lRkwRvwPfrqGv
yC7K5GqIkYbhls5TyNlFmPWZiObK5GxI7csgPp/tK8Pl76pTByzapbo6Cx6QPIWR
ZE3SfIUmSIjzQZOc1/ofn4+5Oj1bSZjE6FVH6QnwQEMbSF1M4a2n7z3DWLit8zLi
MiX9Ktgn+az8tcYZi0VSy7qnND+MIQm9Z/pRF5XLFjs/01ZYrGzDOHNbdetn+Nz4
onWcjIQABZn0HpQajkFQaipzyINu7MdIUfpY9CRiPfwMCvO74nySFYCiVpiTSPS6
dUPE2BqPPCCdAikVL/mvnbNhOjA4nZXTXcXnSptHcl2poImtz2tHyjN2bUXDIVeT
Axxhsopfnt73a0fbSHdFUEMt7ZepkqFHYYiF5VdzcoJgk9T23RKTlcvx1Syv+ZvQ
tIGJCqrYEP98DnSyCEqw56JZsGgbWDWmxoMkJfNeMI06kwSm7quPT/cWaS3l9hEm
pKp03RKPBhZqhd05txbQHGqVb86PW2W9WVoxWv85Rq2/CB6xptE/uIieSFQFX/YN
QjyclV+HUr5wK9wLH+CPVqib0hvuabRr1wltNQlELRgvNnbcOFldukIlcQBGHTyn
EPvSNuKTGSLioIbHN86kQWpfjeZQWYJXIRvxkAhJJ79hluY2WHJ0hbdoZTGG4STX
slXqmx4KNVOw5LYOV18GNISO3gsrpzsekMHZ0IHD17ZWodyuf2Ael2Eh9oe37QAG
Iz66xZAqaABWPw/mbDJGNDyP4OCMQNB7OIVnOhTYvOZmGvQNObjcfiq0+GrnVlT1
DB4QEyD8eipmv2bU/EgKRltykHnA9ppNGP/aOlevqrJGVMK6mCyvDE9dCTzJlMF7
uiVt7ydMEuXUKigsziKMVx3gJtLiw32JYEv4oRFvr9Qb7LdWn+n7aBNwnJ0TfaIO
f0opb9Th24Z3lKgAo3lcEAa3yL/hLX6EyHin/JqtB8XheGS69CU6rFtylTX7H2Ku
SIOzfOvbt4cTPk7aDhsjiA==
`protect END_PROTECTED
