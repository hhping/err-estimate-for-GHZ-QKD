`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
myKcVoHLopsJT7hxqpJSsnfwUI7i6m5qoa6XU3hEveXV8E3FTWYkZ2Sdv5u5c+6i
XtffdOPXDXRXUrli2fOhiQLrfG9KMLDXXZQyGufooe2weNjHvg0TZns4Rzp70ndx
f/wsvuYQ5KEqF+RflAGObLrGwyfwUQkpm1Z8QEPuH5NtPAeCgYHADCSb4xQSqeIE
HGLDKcfcjZXmVc/9WE5pAR7+HkHWDQMip42djS6DOVy1HM2d1VxzJiV/1xC//Qc4
q/Z5inLc9WUwynojfEPN6tdx1GkTK+wwA+l09wAK2VEog8WQnjjIzFUD9TWo1pLw
KJ3nG+jVdgts7Wd25wspOA3iifxbJLYP69X0cKbDzROWvKeGZZkadD8gnMKdgkJL
/PMJM9FnTV+iX2zfi7Xm2Ug6O9jSkAo3UAeMzuNsb8melayi7lVoALqQf9tVFVD4
fV2YmMnMgWoFp+A8Sc3rF3A3uSyME6Wi0+bfttHc9l5vay+vDPXNYWDvEqGh+qZK
EF2dnZrGC3QQvw2TNQosKzDDZdYsnL8ZpR9uU14JhmWTLhYO94P94AR2d2yiyLwi
r0gqWBkAM0cebo7JADZA1XJw45xsMtrn6EzxJel6PWLA6ADjEXt4Y5jHNNdDUnY9
qB1nJV58DxeMhL4PguCpVYakKj7ceAzmFzUDfcG+X7ZyNwGE/Ur74rntj81RyC6D
IXnGOKeX52a7ajSV2UFR5L6aSvxLJwK2O42cUAR778TsSxBNyQ/Wl8XOBCLRpnc3
3L2yafxpuAYEeJBK7cMB+Em+plfthHw5ncjZRUE2ll+FrIxd8uQNjl268pFODTGM
u4giz0T5Mvi+5h9xPyPLmCwO0DmqzC8QSAjMNTy82HQrH0DJV6CZNxHOP2r/Hf09
o8bP2DRY9RtuFbzzs7IgVewhjT5DdkchtlZPVJb6vePDzyfYRZnfOeW59PEYV5Fh
YCeSJ1jFvPynzGOahdbZaN6v/nXAWQK/Zq7K5Cqk9yoJ/gmtaJahveB0dPT+Nlsq
+QiivRYVuX0OTstqSPL095lFns3cwzyeCK26GTS5AaK4hPX7m5UsS2rmUYIdVVln
Tvy9cGuau2hyLkQkEqdUR+fMBE8NME5vq4lwP7/wt4zfPYkAsyG5h876jI0N1+zy
DGGJx+Q8deayeUYxkF5KL3AMP1lfFKKq3F920bnbWWgeOBQbWk6vitCNswwf6oBH
amZ6PvHqcFZa3OG87G5oz1EKzHD3qloBftqqC3oCwGsrUQsmNAEqmHqrlE5fIrJB
PY4kMpG3cxH0OOSd68Hn+phbRmyLkhpC5H2TH8ukvouRFcZnKg27EqT3BsFLegHy
HJ4u8FzgnoIrNnFKYqRIGEdpMk6VzB/E0pXSoMnp61rc8ccz/HOwjMgt7hCbIqKb
BnWk9h15swsvP21d+Qbxw+A7CwJ1cYdEUrFGHvXtZGwB6sdV3dSzGG2OzJN4H4Hz
S5NH+tzBFHJUM2w6dJelsbkMDdsL809DakkI47iv62Es5MWuydkLnMWSWC7ysHX3
N2v3zfBlx14WdEziJPUWCh5py+EAi8avbsWc5vxEdg+4abaOfZLO9CcishuXaAPZ
tlU07H0CN4GDUZ3csXB6z2VNWALfurWG4bddslBMrh9h/YTqqC+/N8sOIMnzuF2x
/9y58njvb+sNRjow8BolZ0P0aRSrGiWd0mDOQ+4Jh9rThU0+fIZ5X39Zge8wDDrJ
clwc8ZMzLvSCW/9G4/8cUXv7bilhkPDLXGHcEbbQX/uE93eRVLYE0PaLI4xZeQig
MzpG6BbaE80RrwF655jrj55GOVrQe0kbEfU4OLu3Ypi1EZ6iEjqyN6582Pz9AbCy
YqsFTUJth4gyR0MDxfCtm7O1rvNwWs6rHy3HBzzeKMNmgxQ3fbV96voQTujd/xku
Paph/Y58oa1nwNNdgwlrold2S9Aggm8hmh8nVA5dt/t4SPRgq6TN9L+rgwiht70I
edn0fVX/8/gmgGBtP6lMB0Wbj7AdeHed2j2Tw/MVZZSGQxHFLayaHz5R97o+juoN
8kmtBKunizLpMcgeA8rwTvnS6EnPIw7gO4h7KYoyWi4PeQUsD3M7siG/0pxw7UyZ
E1f71TIh+Wj8jtcLrJBpfkEkCojIF0x2OMGJBzyP2h0uaYksK3GSrOzpxX43BvvK
rE4He/UPuBcDOJoN+pUP+0FYAO3KSDuCJGw+5+Ank7NsPAXS1h9mxQXS4RM3uXRY
OE2Eu5M1BkPByguCZWXwhnLfLH9CYebe6cPF3Rp6igYKPPRUzZXz9OF5k9UUKNEP
ubEWpdKyulNdIxq/DDdRNmvojdEIDGk62Jhh/sPv7aq8VhSXXwILtxP7pW1AQQOr
q3CUa9GQIVODAtBVW4ZCoq6cNv9HvMPGB6BPCvSQ2xlAxMi1kkKk/g9I3pTMkvkW
rFQ1eocipkjSLqfCIL5YVEYm3aviKW2U6u5RLx6xTKS614gP26CxmB9vQt0QBeIC
wK+O7s1lKjaWFwO9hR38teBlACe8Xe58v2AEZOnFbAiPMHrCe84m/ZJfKcp9GKp5
VWUCLNiOQter8wqxUSs7rdrso7p2+OI5cfEhw9cybHzcIRyfh5e1ceC5MwtFz9pd
nKhd7wBGa3YSMeH7QPPGDttY+eqO67eshcHiebl8njg0MVFzjP3T0s1C60nhBqvG
Rr4mvfiBXxehyWzU5xG0dZK7ll+shE+unRAb3f4ldacI4icX9MTTiNc6/TiuWA/g
v6ZgWyxRPOEDTfEwnsFOv1nhLThirrilqYq5aRD5NtLUGgi3DXTWauBPgCvt19TX
wY96v4TqtUA2GI+HsJc7XZCXpEWYiCQo1BrIRZ752g/6i/1inphuAh5gGh2IUL6h
MmrhaMVOoXv/MQ0LXYXsW9fqANFM1ECO9gMsyB1oZlA=
`protect END_PROTECTED
