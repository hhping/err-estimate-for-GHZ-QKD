`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vTrsnhX4qN00O/fROVz0TWxiaQc1mldEhb5l8ghvcXArYZNt5CYJaxaPLgTJb6Mv
o8wfYlxLDrVGOWDtF+T8nPjgEbk1A6u8S7jdkKa6KMzFLY9W4NYIifJmFdpFqS+H
UfmK6hLaOU4f58bnUd0lRqCcqvyUD4KD5RzXAPTz6ZuhFN71m4xpJAmRwbXsKJB9
twoOMir6FBaD13TdZZHhDRWfCscATzklXAS2M5sq/ardHf8sTa+mdjJxulgkHPFb
ycpAzXt8bT4FZtOwnCZOZKC9RZMGWeIOArXzoIm80/AITruL67RC7b/g2+ym5Zez
PNPRiFmEKb1XPPjFTQgJwkcLP850J3ZK2btiDVcB5k4bk2PRqaVfJ5U+sgXVU9Re
TR4w+/Ua2hP2IfrV5y9RHP5R2fwaJQv1o1x8xF40nNjhlvJABHU7uqy8FBy3KZeW
IQ99n/LulAaIXmIl4UT7ZKM73ZVZp5WeFPIuzjSOBVeY45DYzPZUyvX+Y0b2aANF
frT7hhrjZXGpkOrOIrinNN/5gDc/jc59cUvgrz6rRt9onWPrgat9k99DuOxqTsLu
fOlGo/l7whwIoCAQKm4GH02L5280FTVD7IcMorVeTE6/gQKTfhkrElQPW3Rp/+4K
E18VcbXAqJy1hvhnIyraHOUlMIMiAt0W95NoYS+hLkE0M6fHnxkfSmldQFx4HsFU
U+yk5xeZD9qH6CDLK9e0nJ0Z0FcBEntqwIljLpaMEsGqrBs1T9WUsUmF8emMpoIy
Qzj0cyHqfRUJgu6gVqwy6JG6waAQs4b49AaukhfkUjYxF8qMyReGOGIoGWDun5RW
NsSzpiHwPb2tcEtiVrPkPeIsAWhFX+jUhzc2gv6wc12/bt3k323k4xuKrZOl5EDT
GAYOtCTnV+oHo35JxyPQf9eTNfGU8HcttBzWCGrTdEoi3S7RA/VoUacVDVs/6sqF
`protect END_PROTECTED
