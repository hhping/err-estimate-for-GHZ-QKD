`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fx/0Fw7LeS47NaH00QcBIQ9PVK/Q9FpI2tSb7TLmnnYHXyUWFaQBhUvGn3aKb4HH
4nYlTkl9nSR0oY1fyMNVqH626nYgL+y1yYcjHHc//to/vGmL5WPbCC6V6A3tuF8o
n/kkJUw3oDGX5URcNbPD1kyby1RtcIo4CkR1++xGZSxlnqO7J0t50H/fmqT3mJaD
NGrXCNjH9GF2GRMrUkNQAzXCJl3GLCqQ3n9fSS3Wrw6xOdpuw2HQyKog/Bx4btt1
PtG3a0jpuvdrGgy1/FyqVFFozVXgCqJIGgukH4Zdhix9UWz0Eur09T6d0QZTLYVi
p2Q0mdptzHJM9y5dzq/jmy0z5v2VXHh8sGngksF5VBUx/DckwU+dA21L+MdTISpw
Dy7wsX084TdsI0Sq6g/cy/ABs/MkZR9aL3NsmjPb4Gqd3Tu6SJNy6KU2d4iy2Kj3
axxoDnAV6qQda+ZcL0uIZxPWGAV6IEWbDXKj5VZ06zEA9qhb0Z9sRAoa9m1JEFQB
tyatq4fB9hJcb8IqlznQGQ7vOKqj+JcMGzjaf1EmCbr6KBCTKHayjTLAguandl7f
MakgLJKthD8259DsjL6pDFxub6pdTgCRcvWTi3/hXVMMVc12aAHU2GM9X5Wuo8yR
LpH5CkDYJovSnimIBY5iXSxnYOkw39VnDxcX9c7qVxcZYV/xiPM+wSqOW+tMsA3s
UxEWZ8Aag+bp2NrvV8rggbmZ1SlNVDEZcdRyDV/XIFARWgrJ++Fq9c6HTyZVuf4d
pIu82/g0TDzmMdSg9yzNRppHFT5sxhVeUlQ9ASVHHhUoaqZFTJKIK4xVqjiYgMBb
bHL4hUBfN47kQSwDD0tzo8cwl6YyQmk1wEfIAUbrfs8YD7Y9oXpCECE2x8mXcoG1
uCeVb4Ww+zEcrhZJDLzsJjVOL1E44PwMQ/x2Csq/AZpn+mLNkSzlcBwciK3irc8K
+E6fEpc3D56oWHit6arc1Zm0PwiKjNzWYS6LCL8+N/O6p4ZnO9ahFzZrr8HW1Was
XfTXEOaZ6vPkwCrFC3p4z/UhfUL/IRTM+STLp1HY0MEWm23buHBHCadH43FezzAS
f2xhRyarc6gFFf9qA/YkPk7Hqcdz9d45bG3a0JckuF73E/Flj68qZKsIHyfVm+Lo
OdZsQfEgIX3/0ryYU8wLlrb8SJ6DBOaM7jy+6bkI0tj8WFLWL31hiN72pqS6cdic
p0Ra281cjGTvi7kze/pM1LuDQ5x+xnyS+394RiU/Ig8O34nnDnj3B9Z8DFTw8+LB
AZl0exi5662E2u8Z1EQ8qOW/fK3ELj87sIoqFGqDI0WlSfc/vxLjn+fwkXenya6G
XXRGd9STzI/QWHbF9a5ceAsqM6b4G/L7jlfpCM1hFZn0HdN2gMUs4JEJoI3VJtsV
Zuad1SgEi3pDmroMMF/+tIujIaWx3ksRjF8lrL0sfrmJuj+qHsCOQBk5frL490ga
roKQ5eZFA0KTSjUzULmEFLH7pAxgxNLvqFrXMkjoHCpo1qUBlTgB4Excy6Bfifzn
qdWAwVDCujhkigPjhumPTb9Nb0bMuUAP5+biNGj2kpddoq9ukMUb3FIyrnTiBgLb
Dg6gzUbEgwiNOJ+wJC7e6ZG/ip5lJGuZcSOeQaJzhLtDEf8bQssMWk7w9HVgzi4D
9i06LZsIglIA1nxgyrnugKd6FD2Qa9cZ/4EsYKiDsWjsqQVILCnQjd8OQ9lOnvTf
ynhGcyDuHCj6kUkC678HtNHLtv79KT7X8QIWL7hq7UTcPPZ9dzbvPlw34pBW/h1a
DZfATOMw/tFcClUdpOkC7UPNrjREQA1sO9iGh5QYiNfPGKp3xN9ty/rnDthHIs83
A7WdMC7iAy1aEVc6uDD1PrRnYgjKYwlq38xwxbazASCOQdLcYCaFTX2E/eLY77oO
zLngky7dBXDekBVDMsT6pV4RR6vIa6uMoKc62drMZogruxvl3MofVMbS8+GRUCtN
0nZ0TmiHacYEN7R/0T7AQYuA/dA+0e5aDc2rL+/v33c1JSxB9WpAnVis5j4Anma3
PqKMQpCcs6+kT/JtbgMQQ8ARDveagdXsLwg32lPGF04uJvbQUpPjNCm+G3QyNZij
qr+oScBWtGXSFAUNjBz+4MKG6lIclBy6qBqCzhI7yg4xnT6Mse9ZyZtg0Ub1y5Mb
VweI7m7VlSiorhZa5G1sUhJNTRcET+Q6GV/Ju2i3EgTkLbR36xRCJAwKgkziNfuS
RdbX0lQP9J6iH9GYRt9u+qBdDCxjyxakH2XBYk/+SsP7kYVNYwbSXbv970JQwkr/
d2Ke5tXe3meq91t/HStFePoPsB1cBH/Pj8C5o1zQjQ6phnm5FTERWLINJBMnRLrN
ZD7Pa3yjHuePMAuBzeYvtWT+ftEo4gIa5B8HqNAnZU0f9FuRxzcsD3MbE8LEtFXe
h8mdvughi4wdBosuRwI7JqL35O01UZNkrdyNEaDmXMaCDTZJYbaOFhTmsCEYgGvG
`protect END_PROTECTED
