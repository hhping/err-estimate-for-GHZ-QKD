`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VXuAepm9dyVt6Z7K9OA2uory440EDhgoonosEaGdfGXNc7Gr3oXhdk8abd/Pe+Dy
+6Ng+tgJAgzjRUoQxMHV8ZwxYECMjr679BqC0HtHQiV6XztyebsGRN4YuJlBqtqp
RDupjiKwvsR2Q2bhbVokNDJHydA1dgeW4TAKVC52HeUCGfNbuk7XHc93fbbWGSc9
5dfxp52vJmUziKqYYYDEYXDskajZw+sLIMncq/DeNrNQkP+HwIQU5SbFpYU3qxpD
+xY1JvoJ+wBoYFAfkp+uzCN235D6hmD7CwbOML93ZmpY5Ri36uob+AP/rigoAGGN
NONXaQlSfET4tK3sbohGDF2QfUQeGPUdjS4RlT43F76JDvXSd83Dqe0f0+eil6ZW
o88gETza4BF9C2msSNmXBQiqVXl52p2IF7jcryzOt0nH8aHov5+WbJJq6pyJEE4b
XhQzwydq4fqqY6zZJqUjVtPPiQts3pRKRqM9kwdh7gP0GKDW4TzurkTWIoP5ECKg
DYXrX89Ikqzx0V1oil5SMOQOiAl+dMDHM7BU4TZIwd1IFQRTu5+YEfPYod6DCnT/
hBt7L7++zIjDXhHGQj1HPtwcAKtwAut+cHHbQs5/9CqdhQ6Y6evVNoxOue7rU+fi
udTUklEvq2ivynCitfpHky/z8ezI+FWr7+g4IS9xTyXenpFboTjaAEAif0sJlA/5
`protect END_PROTECTED
