`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Ffnc1cLsz31kgj2qjuDLcovxXfnvBRZyziH/dCFSpdazdRUL1XbSz5b9aib5Xyc
Jt2+bFAO9uRtsZ7kW7dm7XhoTIm0jdHGxa6l0EnahwDGPb2Ak55rWNEMEZN5EUUg
RoK2LKvgMYi+ZErb+eBsV6Hevb5DodCCeBn7ge1/eT9fRwKbX886kGMFGOjoKbuw
dLzHBRHm1+UMVPyYfLInDzXCprHsM2C1+yNrT1NHJC9kff/GDJ9I4l6Pk4I4AFSL
f68deC0ve0zF15/1DMJP1yvPYpqrCGChlY3Yl+UP5kt+xW2JaFbAcQxfn3dr6PhG
m92BdPlztj4ArkK8cQAlHssb1hcv8qbWjKOx12utDPRFyfgWutUBaEU/1VQCIB6u
q5ZDorB7Ptl4aodbbUTvm+DXSehku0rf6Yl0My9MgZvXAt4iYkevrgqUn/8xchaG
wlth6NCYZ0tNSYr6AqebgxZ0bZvih9BteYMOzh1X66B5XeBzp7T5cL0svAyGio6k
5yMLRhDfv7WfSoSFkJOAKQl1yOZBqlh8kuTqp564qBW0xNaW+aqnIAOKYAymbhti
/UkjnrWNgFcRoRpLGRxS3c8eFqqa/coliweK+CvkoILrfrfUkZ4OAXlMP777kqx2
Uw0Zk4oYBukNrG8aS1xZFA34b3Ruh0+lrSsAH6Weuo+f4aF8DeX6CwVGZAY1zEgt
WmgtYSSbT7ZGpPXFPBkuV0CAVRZHIe7iP2ck6lJczMRdSzmvx6Dyqko8vjYAQiBs
5wWQKcVIjAx8hAL4WUrSzvf826bx+TOpJH9I7eRh0hwY25BvgjAHBbm95XP7dOTf
4rVKeKh7FmsuG7i1fh24Jw8yVBFdC3EeSlDb+r4wjqZm5hhnxkwOjVHFHitzGkU/
aRxqc8a1fxf20VzYSHlVgSWPWjMea3agdxhNGa9FNe7P/NQYJDr75MtFsSOBqc5q
dzxEIQxLWx9qAO90REZ63nvBP97BG1NokxdDubK5uCB8cgU1ZtSKueYFanzYyQ/T
D5BCRVrmM37rEJxyMHKNq4DSKC8uYjKO2q+QHqRz0pai+L2DDfBnx/PwyNDISbuV
/8eaKfetSrSjnIijjA9ywxYEAuGtdprfN+KdW+bCkb6xuoGNRF8qLuqDdhqGFFDv
NSH2RIXqaziTf9xb6b1A6rjZkDT6hCK6p1rSPUrq5cT17jZraN/KFxM74NgIDtlY
a8scvYfP8x4PWqntWeJw1gslpUWUFcu2i/CV5b2ggdhCqaQMC6BOAPzPAX0iGbIc
hk2LJI5ulC0pGH0l8vdURV8XTrxMRAsMPbgtFdmRyDHhFIkemkEea+W9Xv3clGqT
QOQ6CpRXLkWE0O6Xl90NsxfVSYlmTqiMjR/YuHKcgCIe2Eu6JPQIJva5iv1LYRIR
GBJ4u4LRmeXfVKLkdms1KTFc3j0PDAeX5P8lzMBSizl5CRzWE0WkBLvkK/w7hwke
8OhpL+HcXaC8latuJN4jFmto8QpZ46ZiPXywxEmAu6cc+sAn9Fp4zWInfUQnx0Zf
12VF7Kxn6SV4sFSLj8+OMeEmJ8gu+rm8iKi2OUPdCQ0Xuy+116SPILXP3mt46qP3
BeGOyuIJ7yuZj1RfXRqeXIUlSIrXQ+HTB5yWrKmMP1iB3ifNgN2ZlxEm2cVsiG0K
E+BPCM3x6imRh9DLkRWu0FywF5bQvFjOnLh4DirrozaT6its/zgdaRZMdO0v7O+R
Q8SCvF4/BEAG+EjhKnzTPFd4/g5oF65koxM/Oa/v0keGDDrZIYC8wGYPuwqIU2fT
DKYVJsh7DLIc5Iu6rabZrgCB96lKrw5+Vk/Zb47tJOPW+MvEdvNrdCe3gdO6L5Wd
PlbIgrMj1CxqtS6edFLn9901AEiD+D4h8rssRcpCL5eemXeji0r0tTghbJRgCYRA
5KWfWJ9ztmOW14ucFBWgABjxvLW4Nf07c5UVREpFtEJpPwyUAg0G94QHkGsK/aw+
g3lkIi2pdnM9GrAPVgnduitg9wcTWpLBTT26NzfRjMMWhtOUiFt9If5cQlygsxaz
pdSV3oaDX0kSXlfxZ/2whzWWg2V1FgFDZm6/Hs6g+E6T6MT/MNw+g/TwqkEpFxb7
3ilUV1u9HF9SM4eUoX06aVpUZ6LVOzI7wqqPtxu299yHXEkG7XLgwd4WOoqFITIc
ObYpAhFgTTP0lLmBnUHSibTciriFSiAFSYOmP4ExqG+Etat4Pi69au9oi2SK2Q10
fCYNhnP++F9TEOKAWHBS/agGS/2+m+sZKjFiKkRhgsQBLtomvKEcOP9ZRknYFWBN
uvkBV2AYCERS4/F4J8fI0/pctZVyL815SL9p3bk5S7Er2uvMub9V++38BqCteGxd
VNEm0sGCSGSVltBVNJfkozqw2qEEqlJqD0mvaVjv5Wa//OdD0wEkIamNplCcfv2j
vCwIixaykcMs04wsLcVFiifMRAoMHJIUph2cwiA9gYvVJ5lKha18aunrTzKmR8Rn
G9LeD+ue4B9yowy22MGsIvt5ZnuqhfuWoPujRTuYPDwdM2HC7zcK80VIazgNd8LK
pcCmELqloOqyJx1w3KSgsSn59hrsePOWnEuO52F3MOxT7NfaGwa6kHKPksYccZZb
FHIjKClldroqlZRSCuFC3k6sN61as863xzeCk1tSbeybWVf448gvVJtnIyP+NHg3
Io6aUQLILyja9BqTKOBWjgfbIKC6Jgy4sBhQHlGuCegDUAN2xFVrZ71cY+/ZfWvU
Beq20gZ0Qm80GeWZRri65m7NyZEryaw5h7z6IKw2YSsbbzJl3gC1IfBIu2/LlqLB
DD4C/vJmLUPsLlc1jHxFqhmNMGf/7b9NK4Nl8QTuRbU6mBAsuxtfevySncJNDxwV
xFewRkBwq8QnZXqyAoKh5dr9rcNQCwn3kN8q0VpPlh3RYQHFB169SRLWOuXzfTd/
hAb3QMCSQN7xZkEJAoQXI1QomdOvncBXiE8Ia8/YWmQaMYDE8SrfLXOMlr4oy4Ka
viRRwF826loHxPou91Fye3iBFT4FWi0llxmkI1B/ngrLzJGtj0yJxFGCp9dRT0vs
BTWQeUH7veikpEJccM0mIPNBbdBQgUixD7cqR3HDpzGx0NPtsp/Psj2r3t2AItCe
Q+mFgOkmOvO2OAMdT+FqmBj/uPkG07dfNuSWVVH8UcZHuJ+FGROAUrnx3ofcmLuX
GuwB0AsVbVlIVTwYP7RWJHLpAf2Sx17wtX2a7N+3Vchddi4wqOLfIaQNOjPabHuQ
51y4Rgwz7TYMV21WFAyZaiKvjC1HiqzWsGIEiBTPTsca65dHx+UY+Qgc6yC0p2IL
v25asmetaRaBVY35/WiUxuhAko2WsGrOEYDPGz0F11Erl1yoYrd/psHrfhPEzKpr
YLJUotWnrNRJLTveRoDvgjlS+r1Ch7aZvMib6nN+p7lulmDBbQU7M+bR1gmG+5+1
PJVSmI7AT4j10WHdDEVK/QjjKsDBv/litVjNcoWr053V64TuMM096akadeXHhXTy
Z8YF+5XNHKMhdlKTql+F9RyouwBTfUFSoaCT5RTrKpwVdTgY5owcXfRz2turm9Pc
16LgCAy9AadI0M4d4xqaYyv34vdzrO+vKLZqn7mSKSe049ztezlSu6O2b0g9crbi
fsfhArlQJjbWL/2SDtuQ0aAwFilW6LT6TTsoqjxa9jizikwNPVWHROxiVemWbcoQ
HUcZF7dD1tfgVKn7wF7GPprCXPiR8mA3IdLhTv+rjmd7+ViCk6a3ZGU0bj3J7tHj
oM86BRWfkAaOkAc3RYkAE4ub82gFvgc/rkVVvpVAYpDOZ7blNE1dn7KJPBiyKLVW
uAMl4XAvEQekD37ohglGZnkLEXOdK2vYZKWLOpsc3JPfwOPWgAs24snL7NmArz8x
9Q+5ufILdRbxwGfWmN/vfuzuEqRhfHr7Q5Xzx9l1MwYyg6PesW/4LRurpWV2NhPM
3a27YpoLCykHuNitkbpclD90o9FMhaXJ0wG4x+IV1MlYkOhNAfHV8cdjlFrzzDg1
tLTZeFMiFr4hVCgtIR/b2bS6pbRf6XPQ+XZpNFFWHSa99Bdi93XcSpBl6bqzM//x
WqD+zKjsaUuqryHg2e+2Cmqshfo9bZRFnNVlkkslObVhkPX3IOn8ujEYzdJVmw3s
IfVaVZOWQuP/+G2TEajkBQujbw72tZJQKHouhxPenbX36W0JaEXWhHzj3WFYcmXA
ScFIGll8S+9znAP+yOXtGJYu5Wuw6GNQaIVyqxc32kGz4qcfY+5fQ3n6qQFmqI48
Fxfjx5s2+vUqYRimEhk9AAnvuKOi6Ks+Hn6C4BVvN6v3UD8QuZ1a1z6EQjNPlZEo
cypE6Vz0RgilKnn5BK05PV1q/DEPGyyKkuMLbpliGv0hWRLjmaNJW15KiW/jtJg1
FvZw5pSROsu7akKM7OeumvbdGCJSI6wGsmpP9F+hXoDoVYlE9Rpq1w6m9ewvhDHA
To7VUuKXNwxLEOP0wUaH40mGVPHR+XfuEUDJU2V9G2Klp0vJOU0LEghnMEUKockf
+ka1lzBFz573WIte8U9YUFCyXcEQh++2LAe9pVO/gjYcGaKeLfa3tPUpzbdvnPsO
EX6Gs3MsPbI6lr0mHjQVz51OPBK7u6DwErwy0HT94ixb0S72cAsssoCFVd+tKaUa
GT0xX4FBAUXGf/V6LV22FqtDUQHcXckgUfL45iSK0j+SnPIyw1zxDav/cWhTpWOz
LZViW9wSBppSfhYSac3fDRHtlCEHoyQVYX/6xIEpFZ3iYSISiOnoRof6nK/Fvx4g
9c2k7W30U6YlMfDolukCDaWy7QNbsLhGIoWm6ZlDhMap/ME66vqzizOI4MGAS4kU
Edvd2XiAfWK3IljprB66EUME0qMlpK5dYp+w9evwptQgqMKcnjBqnUXc5kY1wUOw
IHDkOnoUp0WKJdkF3Oc6z7dR/bVUY3uCDXfGwR6U6XE4T6fszPUdKkzdbHGqFE0t
uLBnOfnVJv65bwUeLaTPdAb2Sh32NKVS9BJgjUecAlTW0n9EDhwSYAa/jaz4oBmD
JCn+sO90w5HEhC6kgIkMjlE+ow3/TH+4Q/Q3JNe08Hawzne6HLGqEgh6dyFBawON
e6MSKyZsKwFuHB7+WcvYYUCEZAiCK+EuF3hglfukxTi1RDDv4N5FVE1MQSCISN1I
q4xatWMSmWTbQT/YmVfhRewYar3sOrsCLM9bYc8mOY1cEDu9N+/tehLuUL7CjEqY
x5cQqQJbklDqQ+PbJ+4m9Ckf2DhvGYwFHJHIFRoon7dTGDPE2ZKv+n7lhmznlC1Y
+lLE9sDd8kL6X75DDdkh3fcK08EPjhVmsJK9tJUUFptN0X6/8oc/HlKuqfPdtn64
dbgC9FLA7URx1EiTFjNeDlmV0rPd3n6l9OY+bXaQSRfgWEL35TTKkMK/c+VO8EJ4
fXfFc80u6j2cjISYwZbTpprxntYWidlLv+CmoZX6jsg3ZR6j6enqS5GmnFiG54bn
r4+5n7IQMnuaxVkV0R9vEI0AUbjX0QPS6ClHx0eQJPtyfJbqrEM3Qcqy/KNN/Ycb
ICAsTikegUJlex/97FvHbu0l/WlsxbPxmlmpxxGMec5+ClPZSPB4gg82H8k1PB3B
5Ds49/R6XDL5R40ZKz3seyEKzpb7exhhlGLPDcCmr+VUbOoF9goxXhfDX9z6XPnz
lj1Nx4T+B78gud5ndNgPCQBh5XiuCHZo50rT69kjAyNjr24ikAxK7/aNIuXbiyfP
Dqi2PcHC2zqPilyJCRgiHjNj5SoB7px8l2IXo1OfGkj6A/Ml4c5134CxCJSaH4p9
D9StxHxWJbeeMP7RLiM1ISlcQHk4ZqLoLtcLpEwqfFkVk2GgGuBZRCioi+1S9s8m
TnLMzkaA5MC22noRL9rkrc+bzY+1+7rp1XxMsAgEDJ1dm0Y3zOnNZV5PJZFeEiDq
5kstMTjxqfVzOlGcD9LLMcyhJe7cy3lBVVpM0MaXWKLOF2OXAzVqrf91/1BjxRLT
8cQ0ia43oAbS5A+1BbQs/f1nWIwuwn502V4D2UpbJNaw/ytCVq3Y+GLIhyArfKCB
PTi5wEd/n/+bolosqg1QVY1msXwfCbZOEx0p0Xt+QdaiROdhEq6R0u97Rjh0Bf41
sqZK7Iu3XPTWk+pmaLMmWelyXNPpG2cZ0whifEpyMxqOr4+c+f7Z+uLmXqjbD49B
CjqtALLK0TSt0mM4NKevk2oceyfhEhUQTW744qzJEbzHpxAmvAk7BLnc08cMhmER
5H0BQrX77q8LsIGUAy/sgPnBr8kUae9evG5oWW2rbemNmKrcWecRfLbqmKPNHqWQ
HODxwuaEa8K404IuXSUWPI7FtMM0o/cRSgkfoZihOUm5VXAx8YdwZTL+qYjZdet0
3nRGvYfLtN33w0kZJ5y6qBaRTz0fM677zvce3eAJersq3klsZIboZ9XitzIdtLcx
HbpdVolhETCFHzK3eN/YEFjYxXtVqHf7QUoGAbbmg1kPjaIKIV/mwrpo2xdVt5JM
HYrbSfNgMSkljv3vE1QJdozq8L7aqNBJeq92F09dwrMkDAVPXVIn1hCM+aESAyi7
8SdoiyoU5mPFhnd0Zb3lTqp/F5f3yP0QHw0IyAo5j53UK9dwYIE5Mh7aZFrKuLKi
OOyx5PnLm4vkXLME25GrSLQAvgPFw3JY+EE0Io0MA+jhlWxCfDwfzRjgZl0dm4G0
OGL+BL04x4LVuwOOuCOC7NFe1ZB5RUeJX6dLDDe5gbwMEdH3ywNQMcZqqzr9/btP
MC2YF+tN5/wg/LEtFKfbXYf5TZbHcvNDIQ5zY4dT/RUCclvvXOSMaY+WPkrF4CXQ
Okm9GqzS8ooUygUFDTmuKyPZ+M6cFvIiwQLIW1L0yPLuS0JfgIFDA1llh35ZnNh+
3qJR2JJj2Xx6lppNljwNZucDnyVGtbEVUWrA4Ix50HolF0HZ/m4Uuvje6Pn2AbpW
Gudq62uyDwhnnHUhBQbpGEKVkhqX9YLnHC1pXcG+0EAz3LjJ8FyoPVRluPRXwbt6
ZGKRq3BnWFDZF8omulhBBINjOoWNMdBByICcyM4e1uYmHttjij7H3GsaMC7rEdXl
tXz6kYQFhuFXs81XU9gyY3c6X0vuS5kDf0Mqt8HeHdcpTqtveYWDcfHwK0gYob2l
3f7cLIK1UQ739EFs1Kt6yhlyzpcW0mNyNergOkM3N6OW8JaQrpcJ5hImduGZZpsr
PigJzxseG+Gdh2wu/p6jjANqgNrMlQ6SB3mTChUrbel8m6FDV93QRcXqEV+0hvKG
AJDWV2KniDClQaISdOdMW1wuyJZ9WPWYyPxEPULItaNpY23F+8LRkEuKK3RuL42e
/n5+TjjiQrTqyLvaqxAql1tAjcrlC50iQQRdIlnSgPGmT08YhygjD+cp7bgk6wDj
aVB0ftn50Tssju72cGCpth25e+RCXAHYpZW9W/X48Mga087h1MdGPOoh56mpNu9b
4tV/VVuu24vrb7d85XP7oZIe5VvA/4BWAbCARgskZCN2aP+VUpaaPsrkAuz99Nwg
78vqhqGYFE2Xdf6RkpmDFePJbJfXw1Ge412gapiv/GtW+u9DJA5OajvDRhm+niVs
wka5vNUs+b5kCHVZ9JzXRnS4JKUCcgIGF8D5oiiWyDiID+QFf+Xoe8Fdl3vf7loA
xNTqvXHn0dATkR3zkWnWhxiLcTNhw9NOO488z59xi+xFWKz9StkXSXtrmWw7xGoK
EM5NSWKf9TzoPX4ng9BwafWl27H3VDkymL84NMzcRKqZk37cKGzBX/MA0HE2A7Ll
Pt4Q0EHz766o7TPKPISD/DRDoDDJ2AS2QMdZjv18rMkY49Av07Y3v1alZJiJBxGu
0gUu9Fs/IyewlwIfug6zy+VaLoGlytrAX3EHxP28/+4mnQt/YyfQHjbGVk+Wzz42
O13sr5V2o2XCtUAJSjDBrvLtlVtwYqYVkYA1VTRGiK39QegCt5RIBONKNEqrQ+Le
LTE+DiZkUsdOP+IKk7yMMq8nQ3lTw0By/o8hUegVHd7OOTVG24odwqBlJXivgWLg
Ei81szz0VQaFFWBW4vCNOTieH3cLTifsjRHZ9kg50F24/Vt1AKqi4lNIxntZ9nkK
XlFJaBXAm5qrw3ohvIFYTTWzWWAE1v3eHiRs5wPLgoJm2h+liJUWpNFS69R3PJG5
jtiUT4t0kxJ8pPULUS6rrciasrGQI+UdWgHeD18ISH7uBEWZZqE3XXRlTKH0oKia
Ozb5+KFJ9EQrvaTS3fjb3sR8GCtZLgZmCp40OziqTWL4OiwrAAK8zhHXfNzjfNEs
X1O+FXkK1KHLsLKywJVu+DNifnD4LIps30Uj3mjSbsYKlJF2v6iBIZeiterRBEQE
Znvfn2OryQaCbtSFb01FhVts3Ox2gmuQGwsjhkY+9BzdG/o8r5rsfjrya3SKb0Mq
AIXg25CRRmVHsO1/owzrv01iWR7n0+T0Rij7v+c7w764oUIPxpBgFjJC5ZZZxkcg
9CHd+pjtF/belzjo2JexZghKKB0Iowf/n27MbWezFiWKOnQ7f+PgmYWSRevm2gYX
tkZFwxTkIpnbHBS9+N979sr1VS8IAZHBousm2pxkCGuYM4KO3dxWOHvIdFGgQ/nl
rlnkS8RFWCSgoBnVMleu72cwRrW8P0Ps7fS7DZGHws4e9NGXS7oELjowwPyqRdbn
Y+7uzxGzgdchwUQuHTgI0aJSwS/Uial9K2cUT8wAKDku5I7K7fvSB3dqCoLxHxF+
AETWnV7l2LXsRiqxHJmLEWbhMYgptyYdtHXZFXzInETWt9E1OEEHNmDoZhEbfDjD
3sYG3FwxnDi8e+2qEs/gzD9awRVqNQK6nKoCEZm8ZPob1ib2qaSwkRLpe/OFVnqh
wjKWOy7EAYS9QT0ZVFIcEl0sTzrX27GqGb+qMYSzLBSfhkfew2/lwCqq6dvczL4P
NuKhnCFUOrtr1NZeCu1jZz6WfedxseI/WrAxI065b/MIQ9/fF97WEV5LF9mzQaDj
J1cDJC9m8yrornSxH9jFZ60Agl8oP2znHYmJ1Ts5ubKA0XfCPwA+m2KqiJXYtzGd
tkWXg/gunYYd2RgqnlIrdYKtasLi5RX3FCNIkALNyOWDTLyE+BRSF6oiAfIsovoF
OgHrCN+oPJdZ+2vdjSiEMg5jf1uKfk205RuqWQK8Zfj7YNrSuBBcmtD+dansVAFH
IOype72mxLDgHq8vQ4LiHRHlf/d+SGcRqceY2GkGV9obRNnTocSZCMxD2M+yrcyO
CrXZFNwPPz2fgCtnTt3XPUlE4Vhw+7V1ofk+8ji8Yv7YHpeXsAXnsw/J0L1+ljj/
iFLgoVgMA0kQEXwD110QBNUNgxQqIMetLwdYajm4dJv/54PElj4D/yz70DfNiw3K
e0+rlFymSZgrgRaLC8PVGbySyG3K9tDDYvgg0bo0gRjlicR9U5cZaA1K0JuNQxMi
snzrZ0K0mMDEgNYy08k8DkxEMwrXYz7K6EGljUKgCSNif33n7fsd7kzWeXkWkzXu
DlFxmZ0XcG8l4XDg26rARnoUoKALEyVVHVmpyvCf4s2iGuNPvE2scLnzOJ5OLrm0
NF0+lvmGc4rgzYpOosJmCM601VyMkLSw9RCw5PK62nLLlaAWfiG+XkIoR7iDpztJ
W69lOezpUmeuH6cQiGaVq4qLzIXNhXHIDcw9fptMAM3QdkhoPyxusnV+x7EigWMO
EA5SKB+QKSeFxXPhN09A361b5F6zbrZ1l1wE2U/r9TkI/TQgu1ECni5nDI3uRdKU
Wg/ZZpP6DMMU5yl3GVc+G3e/+/cguh6ue64BzAQJ8iNXcz7sadowFLMcyWcLuTtU
9r3hdNdW0X8iiWs+CdufWqwuaQlHX9LrYOQcfvjE3btF8Bhhl5pZ3axeEE7z/Rm1
Cf5H6P+oZkjaJKa/jNV0OQI73B6L0IzawIFBbn00xpV6xM3nrGYwgdKqp7YXv733
Z1cpDHbZWYBIBOcpuSU+dOV+zRjVxxy1Le6P5By3AbUWH7l4TPJwUR+kfeoa+tnJ
/fPQmXKVvgpA7iozXeeBmgePEi6XQtxQZ+YqcDCEYEUKr4LwkurbiA20AKD3NBtI
aiKeEWZ/WWtkmNaoBi1TIbPfwaKelGKVJ6jpj2m0XF30I2zVgsxA9CCNS6iD2L8Y
tYQMeKNPdj06he8UWlMMw22EKQdKlZ/HNM9WT3ySuV3RMNljhVKArdpwchSqnxEk
skXKIbm2PAfCyTSs3X8yyd9yY/VKv+ItJ5lwNY7aV8Mmi0D1GvcOcluLk4xjgJJg
aeHhCu5fu7YNSHC8Yvw88/Nje3nsJiMXWz677cl8z2bt/8N2SyyK5dJvv8VxoCSS
I074/ZIXpu6lewvNFVhY+ZRkdjVq7lS3PCGzovHgSSBjlOr0I4J5FfOMkk2aXXdf
vzsbaAxbINvn5b9i8Rw+ocOl6rxEUep9jZleECayVTarEXyQ+xkTr5Vx42NjSwiu
pS7gGoKhl9UySsTqR9EmBRqnnfMAsX3mlf7NsmJsWIsyaYzQ1Ac18HOZxpRb/3qj
LCaC8OV4jt2xYrR5fJr684JyrXYovKEh+sdiKB+3tozLs3wDEY/AsrPc4sHHT8ar
iO6uqnN8gxwQylSm94Bh+BqTaZKOd69wVdFiYIqYxTgHtKIy0p9A8vzWVbf4Mxyy
D43BegPrMaeN/5sj2JC2Hxn+9a2K8zXKjPnYUcyMSoro/JH74uy4fFBNO1nxX1QU
5IK4pIV3YsUcvEavT/hsfVoXn5h/QJ0XAC5Dapk9yfcGCDe4kjeVpgLlMiDchi6q
A8i+m+mlojxRzTELbiSeImYZZc3uorrEvEqP+l7mNdfcxrDVSA0viosbsUfaOTHC
nm//8aGaOX3HV6F0KS9ZKYBQudASQMtS1jzrR0G5NlAqb1i9+VP1sD0ix3NjbeVg
rufH/x86l+JtaP0T3p1ZxqKwvpTc3KE5qIID6l9fAa/UBcr/YSeNB3ynQO5Qf5NO
9uOgTXGzX8P8irZ3yob6Q85z23+O4ngLBw0FgkEgDGdSqJqUMFth/AKE7oSiVht2
EJ5CURMU3pn3d0wvCjUh8FK5biDoJ1+ZEvHq4E/whLSIXaj6PkM2NmXJ9+qfyYd6
mug2kvlRmxnoV+veGS0Z0tjy3ziMG+YXPtoueNzwg4i31Q76PeLGqGb+//2593mf
YZe3t3vyd0YljOiXbWyTAqB9FEzRRX9m4FfIPJLHPn9JQx4JTTI+xr84pQ59oRFw
d5s9bpUOZXbSiZHxLLg9XjZ+iAe5pf5anU7aitwWMvdjM1a4qd/isHHPzYLyCLWw
Q/7Emj726ibLnrBRekUeFGizwdiFiyKzf7YisdMWUgay/NiM+MpbNlbPdfprMlWM
j9SQattyRtIs9XogU+3pDeG8KPhT+SZFxmAxxe1KaS1MQ9PGgI7qqlRtz5rMEGUs
S8AoJUboXT3S+oGXmINQBgXo9ynj5XGsf/ZC1GoFribbYepd77OhqNOrxinWercV
qXMv+q5eYv8rvLRaeh6aAFE+f4U7qGu7YRegaX8VYoQW4mxGRwGRXhk1NUxyCFMx
fWMbvQtlt2zN037t0NuAY2NCJ0JEd06uj1Zt8yE1ttox7Eiew2wh4XwLH3UkpE8O
7PBE1XlW7Ifh907b88pMh4vzCyWBYntiTiMu7nj5xKNYooC5AcGwqCFA7vpwT1gc
foWDH00WkMJbx9e8HgxqhaZuOfhUi96tI92eTGc4WbFElOnw0MAL1gpSaQADGfqj
kNBZ4ssVo3ATC7vNfZ6ai4GI5x6UpGCwXflWK6wJJa3j5BTExZqDF4b0agP/eOq8
CtZgfpOFJE1NI0zEG0hLvnB9oxn/gGCd2T4LxR3qQjLEJgQrdFCr5LSyDBAIfjO1
uZrHq02Ioxy8FopYyA6aiCtif/HywCza5GWPLwyDUd2TGAPjDkxq6zUkxFBY04Fu
6BVWIAQuYJIaf44da5KRaqT24eJFFF+1TARFHalsSYmvKpDyCISj8bUaEq7I4exF
lJKgzB7fggcZ08FnuGa7ndweKWqpXAAS2NHX3a9tqx21MEl4mbZgigX38HX5jMb0
9Uy9vM2N3B8AnxPr73KNT2+DGVXiB/plBlwHvOypGaeJcbOI7r8btbnK8VgsnSkc
aQxI4OQKyK+3cns8RsJ7KagkJqSalivepLyFsF/CGbJBJFOXFL2f3rb4pKq9OPgs
2SQecNAcWELKZqViuNzRa7rx7M4cSteUUb5RoCNB6ZcdUBKJt0P/v0/lKAmdkKXU
QXFv+321GBW0C5ZKL+0PbFsFX5bt8xnh25Zxz7AaFw/4nhtFuOn06MlZqbZxdj77
LkYA3czxpp6EFiFtTtwHUpL3H5ca/oHWjWh14oZhzutmLaLkgSUSj2D8qljTnU+N
ZkefB/WoqkfhqdIX/AbpFEedfEvfvyXB2hPZNljz7KfhBCZ1cLHL4KYRtdFUSShP
ygDZ6VdUWfCcvGWdDbCEpYpBBx3WVyZz9yshJOsANIc2THYoSflUuOL6tAiN8Bm2
JY/r0FDbNIKBupMLNFFiqL8QH13mqlBF4SNqvOFnecbDDheM9UOrHVmT/kPngW+Y
amI5SdF1cgQ/Gk/pvpf+rj6jI24GU7qjvfRUf0t1F5t4BmE68a4Ab52PWlvbSUxI
JNpdYU2pjpy/KbhnKCE7D8ioWwB6N5mIhoJm8tiYDPUex4k9JeEPtRuCZFxtYMgF
MtPuy0UJQ+U5lPvPfi4MIn7u6DF5uU3bRHAyfegmUCTpzpDi8P8jDRzsR1tttRfU
ZN3Nf6Z3DiABcvu2QnSN0IhPL0e/1zYzPstV5IpYvYqKY65+ACBA5xLnS2bXsxM7
Zg4dkp4i2cwclgEM6nYLDBE/ShmaRKYNHqt8+GSTlJ2A4k2ZtKuOA35U2h/rN2sS
FCGOFdnYTqrjtIAX+QA9aBUJdVeN/+JBnXdQR6gp5lkSNBtZnfFr0KM2Al3Oyh9K
63Wllu33NQJYfVNxFlj/gHQ9pGefp2l0wTddUEUAlu3+NcCIsIcPtmfFzvbxynE1
IVzi0ZbhF5/fBAOpJRLM3xaDU3XkGWD9dBoEjVZXBWbVPgx1ycuzbd5C0dBZEAul
cKLMsz7z0nL8wn/jhEKV55OMVNuLgLCLpq9vPZIFAZHsAwBcn4mnzt95svDk3rpo
xw+0I+TZJE/CZvEkx4BPVwHbadKenOzQGoOJMFDtbrJ1h63DNElSeE+B4Fo4AuHY
ISbSGHrG32W1hFWPUYKgL7fWIapuj5nBfH8BbJPeqlmJEoua6Nsgw53AJkcAQ3xc
OjkR6qgZi4VZxMo4nNHpjvPwEOXwDVW3qAJrHX7IoiXgIL8QdjfbUyvzCa0nv1Mc
qNgWXIpW+By9OL6VXqWeSV5uiWvpmBvjgDjHREbhmA610R5Sk7UMCJhvo4PgVl/A
G6Mq3PSqJoDe+JmKBusHXUhwi1AqlCIonLXjqe8ixX5rQXq15f34rFMUZtqQYU5x
W44JyoFTe+PftTPbkqKLxxrh7Vglg1ONPBi35DJMzbhvlRV1QnAg9sNJ9pSFMulr
3j6SjB8/kCeTBRrYxceMJ8waxHOm+0+w0ZzVwJh9VdDTRLYIq4vwsrd9gqy+Vk/r
u4w9AnCvI9JWAAkGrOfgEB5zhKWi9D8jneRjhQcEovll2rNVYw6eE0KhghP3y1vT
/I6NlHC9pEX6hGlK9lwyMjs0iVr9rPwFX1AIYtG9Kt8wHBWIAwNJror3Y26OOhir
oZ3h/IqiofeYz5dzFa3IkrxHTz+l4vBQ/GoMngmUGAjhh8scOhzQ3x6I8TmLpvp/
OghVjHzOKsfwfqe961BIAsvb/b8kxmzDZFohvrIsNNk90+NPGXZ74QxbOtfo5JwX
UIIQ7tw/ipLQEkhc5DOxJpNnsPScIQxBOn9C5f+1nVbkvPoMCFMpSvXvGVW9cTFb
RjqcxrxrLnYuT2MVksiweOmbQ1c2BK429hGd08o7Fd2+/016SGZRWvr73OsOsCTO
6ZTF6Ud8XmRZeVQ0b9TP6hQmg75pdMPzqBe8AjB5FI1YX/IRjD8gaDpC9W8RcBuO
FmBstZ5rGCsJyhNQSWemhFpSgPyV32pT2Yzy7ysokkyru3nbSR76VxBTFgwrKjj2
3shRVStMF1FTBACdNN3B0oftT3X+mjf5kPVu52ibhYAbpj+1cWz8J+xL/x2i6gJa
JnPs/YWyXHsVYlfIWNY8Wd/BDq54MtrzOGPhFInhdd03wKh0KlMl8alW2Inzy6mL
QGADGroee0tmGQ2kB3yMrv5K1f/c3hmRbvyFOzKHfskBkVVNFUDVrH8vGEBDpUz7
dCZQgKD4SkLcMOCRP3u7gd1wyM6AUdJlDEWseRcQX/Eq1VZGk1rDMXI+lftAiq4H
Swm3Oz3zS7t+zZyi73gBZhd8hPDoXqKGk31gdYcRG0l2QgVQVPVT917J0P2tZpwB
0wCtCsfijngBRocaUhagIiJxbchseWfUebKPvc43mJUzu+vBLgIUEo136nWAjGJj
SDcpJqnhADPOZYyC6IpTLzex3FRyC7yLGAcvXC7lbvx6Z9lLKSEQbo9IL5PKbT/0
JDoeJDW8vpOdkUVRCA7noZrZEBVDIA6tfbqbqwZPqqP470SSIliXzNl6IZugGjiO
jy4EzW0p1ACN9I+F5nq/ZkXSU9fs5rJushhH8DxVaE2QlFx9rrcmMBuPptt6a2az
rMaGtIqFQcysf7pA3fwSi+3lAweOndGkMb097bBNtW+wwI+6Uk9w56M3rIFxKiXz
AXp68t08Tes9LHi2UVBkcSZcc9JXQD7YBHFaFAzLgcxS+7avhvbQY+CNXZ8+Z7Ph
Dtx2bm6/mwGlRuC+XY4bY/JP0aDq9DDay2tzOV1lvyNxXl+uSFB99TJab6fO+m8a
u+ZmAdfQl77573hZDT2vh4C6B0EEGF7zoGW9GHkXjyZzmCBwg4753Oz4o+it6YHN
7TJr7SU4tits6KmrYM1kdlR1vnxV7brDcCQPwmypVx0N+5xaK9aIvDmNSnABeAj7
OboVU3oFeoSxJNasB+Jha37yWEwsz89CDGKfSy0D/yCx5hWOHtnYu/HAzCj8Y9xA
llJt5+eXrEIWuqqDdOFmWDJDeJVbWATODhZeJ2pmBfoulDtNAxx/XhoMw6vjpUAS
4kFjut4ukaIq9heQDde+2jfkY+0eXADOCtbLC+ss2Qygk7aaqOLN7l25EB9HEbki
gTkYhl/eix62pjFwTKBV3OkDYqB4b+VUHIsZM0SDZIv3Q0szgTlXoFX9ihDX4SPY
+jVRpTlR4cVxMp8Y9DZ0NR0cLqfG+9s/bcNrBJ1BcCOIboqLVqigM0cGC8TQpi1q
hiILKzWtqxDpDPnQYI9PldvLyQtVi1K7+C9K5I2ze8NaazJyycWGcvsZqQ0n6yT0
0wjo/FlrXs/EuBAYH2il+fBTO1E+t2S1eOUQLBslJPWI132527aiiZH9mhhe9Q4P
FUrrhNrdsPcfCAcE5O8gtmiPSksDWc0Ia7eyEEpfDwTprm0khG1wCU5hgrrCSzu3
cMiqWCNXY4Enud5Ec6l7JGQc20jwXlVbpix90nd6ZPr2A2ddRk5RGqUxcxSBHPGn
4UYgGTATm6F778VtSeSgd/lCPVJJjHelPGcaQ2bmsME50PiQnsy3Zxkb/MRGTWJW
0JLFeO+C6DiDYW5g3v+hAPEAUbuaGxMtwFdhQX+x/UGZEsuX1pjc3sW1YH5lkR0w
P/4E5/XbhLr8h11FFWGySk7+tLIDT+W32HhF8vkUtAK/YLtb2uASFdhrnTWy7wMh
jUmDGqHqqH/QVl9Rj6GZljdkX9J5kPtLzy3r5C1rGmAdMmWhpSfJqfEFWE95aWAL
Yc3DmP8QNssopGI0evyu29l9QsNmw0F7nko1KfICa3Kfb5zfma6pwqeufiDdEK/z
h4gVnXNi5mj8ClPMucL7NTdc6A+HADO047VGH8Wq6SjR51DrBWI96V1n7IwdS1DC
nlqWTMxDg7zeG2wM6+mqcCahXJ7kztkS1JHNx17U70OC6+FR+rwcVtBymjjcuVgP
F/v98Wd6yP4nMpd0bVpbL6YFKqRZrsNG/wK3dlvYMu52Y8aE9Vs4444KOxxJp290
l5gFX8YN08KL1fk/rkdvCJ0KhSAGqEDmcGZk6hioyMi2EIavyYRd8Jb6RMipELJc
v8v6ISLA6gbkZxN3aTeqvWj8W0G/+od+1jH3vZP6oicIPdyxf1DpjUKF04hW51lp
4AgoTJRzkKc/NnVHA1BuQ7ct4mQ7aM2OaqqO3uuPII6koZPz/MxCXCl4nl5QBkA6
Yldh+cfcJ5dHXe+kdOcaEhL9vCQTX5KauTbmX8u96IFFEHGBbX7Gjrk4S1qs6nDW
jfSWTvDWbOzx502+dnlfwrElMqaF4ufn20BFDr/GmB4nichLtb7bm2q8TnxyU1Q3
bEomNhxC04ufwXb7n3DTjead9xe1qTyYPPbMuU1v+340nrPZL//Lt2v0oS58yNMi
SXiZzHaKSpHv3UBy6zbQiiGK0kYRyRTKik4Tpe/lUilOmO3PsqJMsJFxiyNL5zwr
souusyHTbDy+JdeET/6cPv8shCtOCzBB8fP73cY3Wwh5gxziGvImHXIIGQugeYzY
tfQ7581gMFhX33OA9Zm3NytT3ijwl68qU3Jn+gltc+w20Y8ktN1Jw3A3sSCAfJ+P
xg8tRse4hk93FcHK+tf9HB1nJ3TaqHa6Yhy9iDoYtKuiyvgogh2QEi54TF6gpJwB
JCNJBw+sNlqpLgS/MVG6XF2/7KdueuwnjUoO5QEbqIrLBhBzlmzWSASQ6qtxGbQZ
4RyyJusM7GiSFQffrlP5GJ4wR4yLXLT1mRHEBeFL8Uq0XHoA4i4vFQ1eoJtV/I6S
S17U/h7It0UTeQiN7VLOBEtRx9XvzPpHVevg1Fzzi9BfI/dCnnnDWarbBgBjXshF
pZNwEbqIZDldlaARSRenO4ilH7ypOGjunKwqM0ecuuroXifNVKekGLrjUYBytMjI
h0Nyj8ogbiB+0NEHCFv31NlMfVNI8xKQytVyEDpO+5Y3dYB0uJGmm7YbWY7b0lSw
oAkoqNwMTYuQPYKTWlaVpqWwm5yqndIkQ3rzH3hvxgNCnvv2/CDHWYTUwozu1Sii
foWERL78ffqooigBctLMRVgDYzwPGiLXTi/q/4VAV6IBm5kHGIhbNVr+DQaKrhlN
fqigAxmZhUyX3vqBXsjEwpOBZeFkrXoKfuajzuyI3VOlz+8k147FuVY9m3TgrqmH
YTsIVBhUl3lHYxOhULmBQ0KTrtxGxNLYLt4OM39bI3YutLND+vUihwbcgZ6KhFrZ
j4k558ixvP9zfaBSfJwlt0fpfmDuTzfiTnUE9Czt0gb2XhZ1QII+cTy1YBuHWe81
sTtCfJfpozTqT2Qo8jNq0Nn4L1hmFtY+o0OTCvqlLmCxL1EQ5HDQ9ZsnKde9qbMf
Z3RL0Jj+WgaYWRQUUlMXBWn5F5GDsjJcMbKBS5olGVNwSPTLuYtVBjMQf0e7w1wK
6/FmCDn11GeRl+UAP7Pk0RUBbhRTyA6Dk/fQek1qW7uE0lleKphlu0jIpqqI6FHs
Fby4GzJzQh/aDLUZ8IPH5b25Bov1fU/OKDg/T0jeEZDlkoSOsmaXg9L2LuupzLUc
ypC1D7zIDDE3ixo1zaN4sN0vgth8r2yREEhGMS/Um0JWoqa2+XC92f6vA33x1UOu
uaiHeT687oXips4+gCOqjaro8xF7H9ByRSTors0qzgaxfSIcYtDtfopZhcLOxKLh
opS619XdL1mC/kuQLJVvRujdt2NeF2mxPu+L+jFQearVLMkCtOLMctWDZYojLgwB
3BwTUh2jOiN3kJ/M3mHaccS/BAjZ+3Ozzc/7CprqJsPk4lnQU5F4p8rIQd9xnlQ9
4DU5ITfOQ8WuJIHQdQtp6bU7dQyDvsI6O9Yn1oc20XidMlMbGRiBO99wvNLGtNTm
WXe12R4lJcg6B46vXDVup8DTLRS9333OPiONRDVQ6XvZRS4WQB3hhv5phWjJMn1D
bjO5I2Deh2Y9DCEqwsVLOVQh5PLSqfUwwgjBcCWx1FJPuQFW6WmIXODKrig+SDJJ
g1hV03UcBVk7V1F25x49/dLpC6/L59to4rY6q3qzqNxNarARPXrG0kyhLcVIy1jt
dxYHubJ2uk4vNBFdlAMZZOONUbKwxy8bMt6YgP8Dm2xbIq26Mv34UFv0mZRViMGJ
w0zvL9LAdlZIZ4o6VumhoJu0Qbbf+yxaOMRkFY72s4Czob3rSsfefmOHJugSqW1+
ABpOGO3xddieMIpE3slrua4LWfGjz+33c+DfN7GqTF+QvVAQ1jiFRl5vfrYtMLf8
EZMxGUsJJEAePPz04MhLa+0ztOQDw+nvpSTmzlQRqtnbVBGd1vUBIh83d/M9uNIf
yz7hIYgnbriQ3cNI8TJkKCSfPgae2UZhratp8LobZQZH4062sco0+Olu939U9zM8
XHFqSodyLvNjw67HQAn5ZoqtmuNO+RqDUayEg0skrgcndm8BXCB04ZNDOm4T0PbS
b1BgBhonVQz/GSb3PKSD3Z4tbDdIWJDP5ZHPHTfkR9npJ6cSVmZwHcuQMNxKYBRs
lNOZlGA7L8r9tPHC97oK+EkihMZigj4ha+JN9iaQ7zAQOXcF4ni2c/A5LHmbS6yx
tRlhgPd06DwpPzAipodKOL77xTd7wYc0zU/148wdrQy15lBCyARrzLeo1kO6LtGk
lkGOD4x8nW1rRR5XfqHjpByUnuIuRU99aziD0bPbVB9WgC8zVfIFk9s1xsHWGtER
hit/wIcelZ6AJMsDS/i4KGq7x3/YZhn7RfFny8I5Ns9ahtxDM6tOMT0MdRluDG4w
EaSPRlhqqvcYyQ0nCdQl4aE0AHKaOqb/NgkK+GTJ2/aoJhM5vsXMQCY+gw+m2H5X
/fyHlN2qHsjunjBqEMcrJdYjyUM7ql31rA6tDAIJfPo1rLm3Anm+UwbeAUAZg0x6
X9YuayNACKqu1phSihPcGPIri1FZdYrhv4aX8+VmqUwQ9e2chl4rGwPNng1I+k+D
QaCkG3BoI7FLq12UiBnCMhlDkt877baVTr8LJkpofuv2t6n1mu0iOlOBHiuslvcj
rSMW+M/GtWp54YT1VoYzVSLuvqH6iUkq9KqxrDPCIsqWmWHXvd02Q1eMylPnBUEy
5uVFOXLANaznF970bawiUbZPEnUuJDgWRqTSW6fzW13CqzLsjX0RqqUyOVA/QHdf
gJRK+oCDyHZozeV14TaxOnf7oljcH1HUxfzna8NkGEslTiICNPYBiFwg3T2i/1Do
2AFuWOEig71BsEze+MLEbzGWLMVb5/P/4cSwS4BL1FHWEeDBvuyZ7wfJXKuliV6R
3XAlX0of6/EXQRg8Q/wgmglz0Cr2J2D+Un5mJS1Zt3QnbSEvBnz4KK/GD3OYN3hp
QhPixgChbc1q1YK3sAzz9Ew4ypgF3qU3jm/CA/FGQ2+wYhccCLpJytp9gS6AiNTn
27pz2Ee3oUvVHqcvBoovIUtOTeugt/3YwJZna0S8sBimTl4LXseCuh5Acd4xzNBL
FyApxB/5EOCsT7ecBsj3Dgkt9apxvsgJsdhYxGccBLRTJ4HPdWnAFUaLwFmKbQ5H
WsK7VMIfondM47BCkI/ejg3HJ1FN+FubtNhFwYEeXOyX7RXmV8VlhVovUYmc6oWE
RKM524nH8PWeG0lvccvUvn+DU73G8fZVHQmf5VOVH05UVXmkuYM0EAocCPs6w51v
ecG+bCaqc/Iw1GE5AVkgHlIh6IR9c0wC6DxH+wRPpSBmqrUsQyKLR+R6v8BBX1Ud
1OFA06zFZXGlDk6MsNyN55JEUWaVGXA3lKXX0Qf1PJCvQsf9Dr6jyOcTlhMfNKdM
NIYI9m61lmNKV/vlDVGW8REnhONX5lJei8CDZSa0ezTHPas/4aR9H82fEy6D2pxS
4+UFlHPwBI9MO3Bv2ayQDw++qY8b5KXFWrqce6qsq2eOxANRRk+xjmeQD71zZQkB
iuSWn0gjU6w91X4ptDzy/lgpaclobeTiRGBMVcdieRGiNmcE86GpBficl7uWrkny
FxNhPY/OaMdLLQiYw2/jlXDIr3TAhAKynsA6rYq4JY170xePcBHclUMGWIeB+R3V
9QIfn4eCjq5eIoBCfGBNs7B/FsjDPkLE02SQX3KnKVKG+85GNFbs/OO3E1X02sRy
SVQGVTAb+ZrZArJKL1pFpGEFxZD3boT7Bg6+WLbLZ5d2qS6EP5ECA2iOWPo8QJbH
nrFIZpzqUL2Jj8PDE8hbuBxuhdvszbv5tCK67rlvDMAO7CpDaZp161oB4FrwifDR
qdgRvalN1Nxx74j5AHCvIcHdTholIx3in/sJhc5LscsE+Ko0I4TJfWemXzQGTPOj
E10fyfUNOC/3f54PcYir49zO7ydmRtLVyeXLu5NV0mdw9tiEDZg4tSyx7Wqj1NSk
GKBWxnMxD3iOgcUaaU82aHK6Ql0q3up8ApEbQ+peay7XPd669KH2wVce7MwGrs7r
QWYd6FLFyh3/Cu3MGyT6wUhkpKJQOtJ0oePuBZ8EGBIaFs1QcZbxFdu+yvGtkzB2
7DUEhp3oJad5mMKmsRHD6r7E0OQuccjWKMhzwjJSmqTiQFB/9B/Ix9boih0PyCjj
BWAOq4mQ67ELkcd8Cbd0DBGlMq/vvnTMT+1AwjxiN+d3N1/xc+A1OKjeo5GvkgpR
il3l8COhpx5Bzd6pZuDodzZZGGQUSc4zF/x0N3Swd44GLHR0079bYVCmBfljjxU3
ZrJ3ejIGbckfo/XSc4B3bw0icUY+borS1bZxWcwhr7+1JwiOXU4OLThfpFEuwLQs
D2u3E8rExlBHwVAKcew3baxV7yPSNIDa5SWDu59d6pyk51mP2F/6oPSkCqTbWnYT
580+FirCvd9LmByq26xFGzksG3quV0IWJXyeGO0agwfwbrpuVD1xgeyKgvClqDA9
h/OAGmwVGdU2aUaR5ph5MJfLBHQRFT+oqG8kzTH2C7nE7n8Fn8rJ/lHSx/Li60Bw
GyJs97Ua0nlno9LBmE7u3QnA1lVi/rgd9PLRYMvzJG2fuHNhUweMNv5g1F//SbCY
nbcmiKola/wzxSLdFO6khrvLs590GpEd6VFNFN3aEebWWyVqLdV2EE+KmPiPYVls
qquiTmp9EQGFtRc8bf0SfiGg91aA/YUVv+bZTh+LPo21MGgdr5Bwe18H6mr0bCyQ
9V7PZgwvIpoPyNu05YKxHnCJK3l+r3gtgvxhXDJ6MnmSqf1ruHcExn30G0CM2Y1J
IqAT/Jo7GPLH3vgVsdLnlxiT7AmkfpRCb00Jxq3dLrfYYnloTLrIIPdqEQIveTCD
ZHohpGmTby9YjGL93rZ6tAKII4QJvVV5WspGpBiDFQvXsq+tuVIB6vYUBmyPpUwt
gZj7C7qHM6lzkpXYun40+hRPT7wEsO7Ow2j6IikbBGRjdUZMVbfJaN4Y9wFg80kF
wu66M+TLZ5CgS+A1m4JyoC3RUpTO6IxtqdUHqnKRxRf4wx6rH/NCQ3foxqTaxkUK
j0K0Zj+tJ17jBa3PMx7CvyxbSpZjOoZBuNZFMaXAhEA3skG7DKsyqoaYeb97ZT9n
8a2L8xD2f1R42uYvwhlbw2nU4T2MjfBcWIr0/L7frU4ekDUD9fUlbXz51J6v9vv3
WOgxKBUnB5Z9LbJ4LKxADa8YtXi9tL02Z1ZqgXY+NetTce85O+v4xQAjJpKo1mv4
u3pWy9SyjsBkcSenxExz28SfTz9EFsWsPBIMxEGnPoAR7VxkaW2C70FGMtqTSAKQ
G3gM47RTDREuxmdFKvHWTpaI0Ylo4MymjQ7Lf5Vz+m1jBdmS5QVxVoT0lHFmQq9u
zz4N3YIOJH22JIuZoP9ezC9djTVFJst768Z4jmGPlz/nw0xhMiFBgjAzvejmRGkR
9H9pzcA2t16P/iMiwvZ3oAgDb9bn+Smv6DIqKm6l9KM82ug0NfopTE9RjJyYmot2
DrDEmIxi2KNkbwOw5BxmIymWYl2yXH2WtHEDAvBO1DbVnYfs7fI/xhgIOuOHR0EX
0rkHTutcYRyG50biK3eKugDuIuvpNCCpI5U+L0JoN6jny5frtJjXJTmTXYyrCHaG
Htfiod8BuDPD8Z7yK0QCPojip0D/lH3FV0aRDJHDPwTMsYwpB9mkK0BlX+YYW50U
Rj1YNiYhDx/wcFHfvw3h/ZKl9MSpjEuj8sPwn0kuidCR6Gmyxg5nNIMs8CoD+VfG
HLABiFWQPAzp12sRkPrGRvs9sfn4dSA4D2o3DYkA95Fj/FdukCZDgThyhE5PoJAw
wHThP0+9BusYSxYgkBo5sL0zmGxLRNLCmZmQWh5xDtBaUIAyF0WIvJK/kjBOWKFG
qcVNavg0u54LAA20Ob9mm/wt7mrBkwnZU1P/451CW+B5mE0EWzy4GeEDPCzwg8L2
mWAcTdryLmzbqYi4HlBwnCvCttpBl5vxow6k7gEt1a5yIticV5IwUhDluMHbRDxf
NFoUi+x/NJ3ZvTRM0B0Ua+/rhMo8jlwJs4tQvs6SxTDN1YIbDaJGg0rBdyXJprBX
wFMBT2V1Ht7liCz1CICUmSSzhX5sCQXFOb1PNNjrtjhKgNeg8IjlQxnKb0bpXzMj
M07xfyeozLFRGwmK2kq326ftcAMq9Y1HLKdqlYsE/spGLZZKwr2AzwQ2lhVARGkB
om2etlw5m6aQXLQpA5dwGvMTuPSffkWk8ra0Ra/whJqVulVURzxLSV+FLvZZgT65
KBrHcupqzxFVgIR7JCApxrCoWkFQb7D8GtqVVQYPZfD5jADAbMkJLz0oeAOfLwdZ
13q2Vj9ZDRXgLJpBZY83He9MPnGqc89FgyYKj0Sj0C10C4Hl6I33rmkydc1Dy5bF
7wUniFVOCsGAd9FDjsbvrYMUnIGApoSvkfty9JRrM9tmimsuv3uvePrRUdIIFfOa
jbyDHHIh5tAGGzh75gIq2fkBtZWRTlPvonm8T+/vMNK5jGm/eKqfXKX/Vz3AawPr
y2+xCix1Y354DJtfFydZhUBoGEny1xNvS4xf7fH8bKLw2ToOYf7yOP1Ij62YBNrx
vVkYh5CXf2zfM2UTkLhpNQ433FyqIeh+BUoW/ufDl97dc8wxZwlz85V81vQ2Us0M
04ZV3APTpP6ZoifnnrCkAMHMWz/S/nGg6VPRVLEEAHptz1O6OFGiElkOZmNGHxR+
iY/MY67QnjkwqSMBk8D2dfXLQzymOXenojYBnfSFVeG8w3xQ4jCewaYeuAjdr4vj
j+MKgoqqP4C0AbO5eC+aiFel0Hh7Gm7kpBBdQJtoKh2exPUI/HfunutDv6RA+b2R
s6G4IjDkWCopGw/NOrQmu4R2gFBstnvwoTXguVfqlyEsaLqw4jONlauApVhaGaQU
mv05G5B1TO5AmWzEvotDVkGEsQmWbPJduOVx49JBKUcOiybzxy8HK+eM9sUWUFU9
sA1hkhRqAHWl4zMSD+pNrXWxPkANCxqLsVCMBKtfxmt+SwvSHQuWqeTAdBB6Fd6/
ytEi9g6R2zl90J4og8/P6I9FEuuANV8m6bOCYrTuhTnlkR2jY66OQV1qgw9ewQA6
ndgzDqXyGWtLbbPbvgjU/FxsEVZcb9YmFamAtFte3Y3DqBQHGPN8DyDlzUgFwwXb
/SSbbwsKzdvpkiEG6txqKYvaIMMXvZZgt+YM/5maBWcqlpdJLyaJFUeO1yd/GrBw
a/js+drWJF2VIbjifaZEHDnKM20QNMrPwoLRVlk/+Zi7K5G3kjvhVux8sICH9V7A
qFcjUyZ/8y+mL3ovK+cs1aShMbiaUv6uD2EUgJtJKUtSSCS32LsUxk9YVlJYOmtw
klVyAN8VxM0ZX21qUN4p/u4+yCEB1O5E47eX3vCqLQVBwHZG1p81jAiOTGsgbIoo
EEHrELNXXhagFEWGLi7ubPKqmOPd4M3iQJiwjI7AJIiD5hNUVsjUmGOY4eG7P80i
2QcaS5/SZxwzlaw8W1JaSHGrTAwv/o004CDwyON1nmfxFK8wCPXw2map4LlCok2U
N1ymMMPMtn4BnWuws143imaPaC5FcmzLycNVjVuBO4jPI1OGlDN4pMf+ryfo7+MZ
Ua84Pp6huqZ2mndnZ3OqsOzPecjMMfO/y2DwVH0WD4id9S88o2VG/QOo9vV5PK4b
kN7hL/+kL705U7zXQK3uPhBcyYs9zNUlSu0GRm/sbvuAASlQGjhK6Jr6aKDdDhkQ
aiygQDS9JZeqqTk6fGFlpfs0LBECtQp8ReqfcqKco3o7SuDgUK95YF0UVkgfsv8p
4WsKGsoyzmBKtLG1emAxGZkf/YjZzWAmjOTrgheXwRkkbo5C+mkhOWYF0cr0Lm5z
TRHnkzmKEJzsU5qt5MemwuyfFUXRW7QSU/Te5Ef4l3/MJjsVE2I+yZlal6Fnr4Fi
2FpkjXSCVda1mzyB+Y7DbBGViIskC1Z7zXxWD3oLDpfQZtf4TssjinLaQdRU7Xik
MVyLQceWcTry4gtuBuDl2ACeo5TCEVRknpnylk6W9WSl/SN910ik/B58Pm8k56qH
JQpLmON3iSAEYH5huc3QFV/MEAV0XC/mfN0cLaJmvlH8cYD2Ky/ajoYW+2Cf1ltm
WuiSLtI9cKz/3N0SRWqYPkWQiqqeyM6Aj3rdNN5xxCqxf/VWgbXsXgKMlmRTGLqa
4/nCRrdf1jDZXBqjFTV1R48e+v0geboOi8ZLExXdKfwZ8NJG4Px/LLN6p7IKl77J
DoguLvbdVV/ylbSdOp/UMlWkVkV5+aC0CiW9BaDIW+T8JZcDMKPi5/HvcEeZEnL6
yfZ0S7I7Emt3It8iPwMCwPRBmxjd7XAcJXupeaazNF+SEi4LBZJjqzQtV35HvrXa
8ZAV5qGVVekq68dEJEKgsR8p9ZizLBYCk7bxXL8b38wL6NGzQwBkBr9YRwS+17b6
M+EOtZhuUV5HtstvZG8FO3XSG8KasjYMg+fjoOalXQvdtt/Z+OEHRfjOYSSt4r8m
br90kpTHEQa9oqQpSvg8LHiav+5LN2odJB4PLF0RDbC9iEY865bgauFg3+CKCLb8
BXehgZxIFaO+oEfUMN7XMWRt6Va2PeCd6p2CGSJFegC72QVp24B3u3Kp6r01X6Od
m1a33nCaYeaXMmM/SxQFLtXgdtDh+FjkhEVAJpioIcbwObOt0u/JLtMagjuvRsnl
8/fZzuC1zBFkC6uCYrU+WHbw4uitK9AZEvLS4MJM6x/v3CNari9yv76dO1VCClxc
gw/2IYQMNwoL45MnTqLwbUH3g9lERxojxhrkYR4uhKLh5dSZ3nEgqF8erWEb6JtT
yVh4/5vppoUU6hPk6gCAElr9HsAPdLMyeQAKKwNnYTAG62bnYn6uIBLwxX3FLqb4
g1PP8cfDvaXTQRXJlsWPgnHVNj9GtBCKu4RRjKU4QUt/6TNqEfG3Qc72Q0RVMbUF
QtYRqvB6MJwQdTBeMLxRcVHofUXNRdPOv7pgAemxYLEaMem/My7BRSEtvp6Nz68n
7Ky5xM59+bjREkmalHDDM72AoY0ht+YXaz9vFdFyd+3fatO0YRBKPiwrzVsqCpXc
fHmFsaEDU4fHl0SQ+EqFsj5dJjfBtlKUDwZhOH0ovgsbbLlTReCBin2X8ScVzudR
KD6bOzL+X3AiYak7eIZsrq8Mv6bNVynx/JQGgyeLcaWi+qrwpvyUJc588P4k6tc/
hEqtyFdJbiqZeRe3lckztXy76vz/s6nn2/FGUf4eDx9xVsOjuHxn9W+H6nGdptvU
zqZ+cWyTQfbdqJMhTAFG4kT7Feo7AXNPf76WpRW73p9tebCruSc1FQGZ7LjPNlRq
GAMUf8HaTW8XJRsayEiS8UG+NRmNBk6abO7D/Myk+SKvd6TQ2I+ZEzHEMo906Msv
Nti05KZRpDmCdDn7x4s5J8Qh3a0dCkOa1+OhNkkdKOhqMA5nM9EemFGw5RhrGZr/
EJtPWZFFA2pbKEOm2xUFLK73aKhqJW8mr1Diffom0AjY3xDbp6Z24D+q3Tfz1mwx
91pDAVPXB73xD6SRZYvNDT3mpkZxXbZmawqfV3G6GBxGcFhvVlFJWBhNgId6UlW5
4r71LxLCZ+q3QPClAc3H5kPOEWFU273zzjO+jhANBHfIUnUvf/2+2ZtmIlDYH9Cl
LWJRyutjSH6ycFfahVq8nojlzNnMsd6NziYVnP5oopP4ll8LhkEJ2lQrvnSwHiAk
5NTiXdR35Ee9utNBHWZsjFDSVHWVq+69QH559HsicblAsHuuhsxNbhorgSd/bwv3
gdk/WAAe2QcqOzoI6VUu7RhpTd9oJrxSJtiDe1FB8Adg42rRPS9rEmMODmqT5gEb
llIywPuvIhdhwh6WbRisfRULv2fWa2eav2XyMGL5Jxpv5wy/XNICXH68DznppYsh
ApCPD/0Qwe3DWzbepMx3cClGcwEQKfGoz1F+ZASWJMFaksSZVXr4jKXiZwG2eBd2
ioBRyJiUxrXjshWUjGfOwv/TidU8JxWnQmQkXbTQYeHhl9RUyJyfTUggj9zUVXDx
coFQ8LQ0w2TMr53ZnrXGrU9dqaTJoT2GNviN/WVAEPkuYhODqJZ5Jqvnj0vaTOYf
J9IkghbC0oy5SvxQreY6vRumyfK86sRsCDsbHSWGl4Ujiv07KQEURA9+KxK/O4/6
OH/ulpLUEVct8u3AD29MEXCN/8g+B+cy8COp0Hjd5HH4V2iUUrpO8Xil+hCGNRmJ
xd+ljwrruXscr7XZ4nPDQOzXFUlYOfsx3WMiZc7zQu4Y566j4Jnes0u8WW5nXXk9
K/17dGI2P49IEOVvIFMv82tQ7s8TaE+9VFKvjkbumDNDS/AKMRzXU7rWUQ65Aeg4
1GUWDMZgRbPm0HuepfbNJEbtVgNjngQcjr4uxGh+m9eNJfIDoJ0Nie59hmaLP5GE
I3nwq1Rgk3tpeKFnPZEVLbwvAFiH4YvUlb10UiDwIBYvQJHO4ehMWsbAboGLr7H7
xlBmkwFLligqI5Von3CR4DhfiFtCUcnNi2yY+zDK9QnznGDhVEjilFszJbDo3jEx
F7DAl6N+zizHffbNnsnv//wNbKADxoZRAHfFL8i3OgQWJiZs2u1qECacKLR46COz
YHkZZc1RO6UUdOpOwek003s9wqf+T1VLdPPsmuknIcmOpY2uXgnr6zBMeIDNSrG8
5XtT5IUK7YK7KRTwxAH7m+yvslwjfS6pmHbyDREGKv1/lOvgVt90Qpwvd6mMH24/
QcR1GOBvV4XuiOEYU5wgtQD2weE1DtNIEjJoOASwmKwwEY/oURVdMUwkkpyCfqrK
dWttTNJ1UEtLra5z/HRbofz4ciozxo2mEFkH0546hwSk5fZuam4YNpSCCIxX9hpH
5H9uFubo2K6aqTy0gY+q6mOcL5n6JRHnzJyyygmEBlGKH8/DLUiQtlg3e0PEjY+A
JsU48mbpxuLFEaqc4wk8/2fVeO2SAcjG2t1KHtGZnAK148dd9rnF+8E2jKyVYepl
iCX+zXRa0X7iRxOjrQ6nXsKIbXvXswJ0jLB2Iw0iGVQv0Z/w9DwfcBcCbGT6xlK9
H7XApdTmw5llVQgB612moTimwEVsd8ux8NZEutsuE7y3x9ccUD0GJJatBvfthTMl
1Osa5e6AlOzffMBCchhaURV+kYYjt4Kp/9VWHbLXslCTDRp5cTDwQcBeyrt4KEBD
TAuHHHFbpGunhkMGVjIQlhrjSk8FJlzka8NHKUZImuaDcFVnIzPdAohmCFVrpk7I
cFHyrrGXwEu3Ahqu96CQiEf8DTwLl8a0N2CYom7VZ8bEc2/Tn5OOi/x328kW7Ool
EstYx/hz63OhTBs20v9xHebicZmr5bc4RH6mqafpbbfnANymEaEs1bGGizEh1dZP
77OTRqbEJXCRKCEYoIQVVhMTERhYS20AhjL7gfAviRNH+kU+5cLTGfLClIS/+f1A
qvBB4a8czyqnVNVste1CHILUbZP3j7uBk2RXohUMQ+DnPCYvN8xu2QpsRxuzstGN
ergpXP8pohiGioInfbE16ZZP8pRldvQudJdF45RgJdgR1uO8mfMiaIOzCpfIrlxb
t78m2lOLhmpM8KYZgASANwz8eatSstW16G/RRj/8bAfByM9r8A4jS6aUgIGzmMFt
IoMGfSEGKS4q2hdUWPt6d+R2aEC0Krr2EeCkXmsPcUXlsekqnQw3lW/VhMrCE52u
t6RcGBOnFQoeXwVhHQgXB15MumzkPikffakZz49IsrubaLcbNndEtyGFwIOG1SAI
RIc1WiOcunJtF8hYsBSDVD/8N9YyaZ+Lg3haX7BwO0WzIOrcT3rHDag4qEP3zN4H
+p6fcRKvTrJ/UrLHF5eKDMbSCIJDyJY0wcBfwpR4OMd2OqjlahKKOruCz8cmY6eH
FeZVg4nc7skKQQ+8YmMVdHJx6GojOyN+HNwMX9eIBhLo+PGg/53pn482SpbQFe72
uUWQn8cN+KTbL25uXhQ4wXuNz6+9ufzStzC4xth6c+vWWYSYFl/0uBE7dnJ1Uxeo
l7ywhrG+5eKXDuLnI91Em5s+xyChLaOLJaI4YIrSri3xBCBSDRSmYsY8/0TAm9lu
B+LTBeP8Sua/wLJBuYqPN6IFviwJt1lX9pT+TeTywP1edwyuacwiL1RSedBKAK1s
R0HND1+CGQRcC3PnBp9/gLw0Vg1xehaVW03IYT6wtuywy2OF5eye+tVvOBAQOwOU
EN+MZ/dkp0G7p+fe6WL9Tdk5b6ctY5ce8yZa9E0qXg9afU2LxQd66IdH3z/7iS1c
oDTtBAnFsYcvrk0gIy3+qdH9YbtvP9OYSYptKi6F1e52iaWuC9bN+dcCL8cLNRQi
YDzCxqamTX3x5SXzbf7jOmlLP0jXdIfMH/qV3j9B5zGwPNnSmdWAeKXCAzCRf5Js
OpP0IAZ4mBWKwUFsyw2QmU+VD3i7Hh0q+274HFzlz8mGRLAcjKi/tcQBPI5wrUA+
qy//Wc/3iMGDWfq0AyZNYIsDwXJU2avm2hrc6XZJDUYh5ssUAucz0kA7F/4czEJr
E3Uh7++42dRMXcYF78o/19no+I7Acwp0K00ZuTmErblCCZUDOsEmB99J/tqgy6Ue
j/ufddyIcF8GuQra3sI0Gkutnth7veJs5TQs7iYsSP4/h6+hfs/+ln8rHQQsHU03
g4elLG9UWgxvRBjrMk7mccvfn9U3yAKF/TtAgNnA+psrY1p3sEJJdB7OGognt148
s5dzf/X9tOZgOE5m7tm/1Q5VhdrMHSr/8ubUc43T7vCTzfmVp3c3FxzCkP+7E3TH
6Lsu+GrZ2z0VtYvyy+IobA9QkK4ZPt6xyH7fuGvTfttGgmcnz95fjEaSzFr983aL
hEh6B2+mmB9N2qXnaWDuQaoQtoLblftZCZs//klqjkFvRN3SPeHmtsjdI7I+aZ6H
nFitIuJUq2fPiNdsbKmgJ56mcqyYgML0vJLMESLsvn0PHuUDD3m15rcY+k2cd0Ys
+pM00hIVXVucGXMBCi5GYV61aC1LAnssJl39myyWjdnGr4lN9isV1UrFOn/bNA4a
vX1W4ZEwr1luU+dwhp4oeEtSiyTOx9zGEwDFPHTPPUi8w6LhnNgluIxTth+julwu
BWnZo1h8EIDisdCVfffqB3H/2GD9Noq9jA4v0fP6Nvq74mShG9yWn2qI10rjWw5+
D9FRKhHezqo12oitI3m34Gx2EkhDZxg3kR2WV96N+cAzzfJ4KU43xTvHBOMEex/g
CKfY3vBLxv25PspV5lt9N3JC90PWdg9Wz1vc1AIYPLuU9oHX/3LukcEK5p/nQsFi
j8uWzglSY5opFlX7oNDKi+rDLjRtyzuneHp361N+UauDRjNSamcVBt3+B011yHcU
XYeaB9cILNQSt8zRt/aVIgPHud1tFIcY6kVhh2mmhQYOTflfRUs/XSLiN9p8NT4a
OMqfiR5s2amS73avLvVovtPkV038Z2RRP3c9XPydJ7sJ3sJobrdU7zP5vYPlUTnf
pWL8Wsly9Z1k51C6vPUfcilKSD/Um7e21v8bciRzpZ70ohkDXkZZWT3OKFO0Rtot
zSRsr6PZxHbDaWpT334lKKxPXTPP3KINPzc0tDQX5PKoTLAgRk+rHGjOy1TH+pX3
T6a+o7zjiwra1ltQHmSF9Z8gtPklHX+hnNBCgBMi+Y0TVc4CPxc+8vX3189FOUIR
jJywka1TbPMUKt7oYPYD88VLhxRxMoo+016K5Bk+1H0eegJmf8ejxQjNWxPZOdKA
vLzpSAX00uRzRoRrJCQjnCRd/g3BPyDEIlR/t1r5UP4z5f/9nNgYYN8N+GbazTr+
kKUvJ+SU60wHBEqNYz2ikNqDcI73DzLLfyuLsqXgqe+cJC9Ha0qHsoj/yhUplOoD
A0gn6Weyy7oAQqzZZHrLseQNKsGhFug7Kvwfs80zQcylYheq4a7nzleXvTfPLukN
yBWLJo8KXnA1CzQSNLPQ6zL7QPObBU+QmQYOoAUHt5g2IAVCnKhLIZ02zZJkLEMa
VYaHzerYv6bcbB3kf3Yz69ZKr0X9SbLfrXY+fZgf3lKYZvxJahBCilAvXlxgP4Jx
K5anroYbCjfKECAzaxDj96VSrSEDsgWqOHEfG66vAvL5b2fw9y1kE7rbRg573mHE
dA/aL9zcwXW+8BwGFruWCwMGPi0EHTX9+WrJkaQT4ilOa7dXiMLSFrP2ebOTxzlk
BejQeKNGWu5Kr67hGQxD4d2Jbs64M8ZHGgA9JpwrFREmP+eMWgy7XunHvIB4P3GK
wWH92O7hMwdLGkO24xANIwC8odMLNUm0yICfrDF0brfHexqkWzu0vcwhdFKuieXB
rtvjhHPIFyZxlgl/r9T2qsd4zbESwnle+DyrGrkGgKG3YlCiS5E1aLHaG8ftndZh
eCJetVkBPELvPfjrf4vAqNX0MTK32QGW66yOcfA7ETfPFJVJi0cIwUaZTd+My8vp
rl1/sfM2MRbegH/qMmwhijeeyIqjdP6Q7mhk20IvuGcencR74MnLhbqq7DxJj41S
+R62xlh8EA7fIi5djrygOAB+cF6qnJzHfUGBn4rZRPGbsJ0rnAIhHfUmWXNYkZQx
YtktS400rESA0sQ3Xbf8UFhqgSxZCecywsXII4GXg1rQECYlMPSpv3UaIsx7W3jR
RpLCFNHfDh/3fxAGzYmR+KawagocAvnt/GL5OUiAjv7W+DdP88mt0DnPjuLfqtW3
R6BLztL0IySOQO/IhCgeoL03m7ej7bFDR64BTreSXpNWVHUs31tAFyuY02NmygtD
o4qoEb01vzdKAbsVCvm+ngY7zNmTYyj53cf9aqF9mh26r+dxp23KNCQU6WXGU0rx
Rp+0TA3lMgAVGu/5ioNCfP70xf+vJUkqZMewVZlj/uFjCPRAeBhYFo/L+xkSOO7z
eBgjwmFw1VOt+de7RXn6ee1olf6xw/ujW+FBlw8EUFCdaGTH4YWzxu/O7dg+85zN
n/Ywlf/noclSBhUYmyFootaVAFOb7/ZqPxamhu4/Ki4e+FuGxMJi/nNFfbyMo94q
KMAN48rQQxiyiDrBC7sdz3cSMDwl1L+A152kgh+zN7UWPmjkyRG1iROv2em572jb
D+gQXd1MO97mi6/J92aVMvpT29l451SxnyTXuji2nUwTKFjABhluXiPBjAFW5JYU
R2hf2VXY68i75+9ny5vwc13AVQCjzvO9Hpp/O/9u3AbDlNSr/eyeWIX3nHIjU/x4
WriF/fyQaHi/HII1BuRobswYfjnVHDXf+5basTL42ZMrd+y/p+uSiaM0e6gRI2G6
7IDN4TurAU76uDocXYn8eWtxMwl56sPPfy/KpO9kM/ebhyGnyu3YQyqm9eDChZYR
1VpyHilh1ksP8VtZvP8GuyYzoV6y8q1WWnfTY4dH4dhevHBEEv3xvW/xvr/CnGbA
bivdlaKNl/YQ/KmVRaiy/4VtFid5UIHNuzf+xTi319m7dmbL+5mDRVMB0dOz7xy+
QBOJesBCGGqf9fHQJ04EhFzvCQRBb0MW6z/hC+1C8poOqyrdodPLJaDdIw25mbrZ
UpORQofOHhAYHXYqmWCU0gCNEXnWlSIytK+F6MUpNt/DeFK0c6DsSHNK/GbgxZMD
zbD4W3vsI3WXA4cLo/bUDLu9MOkXICzH6ktlET2HtSV26FSXCLzadJNL3kZT9EQE
uX0hpiSLq9VXZv/wOaHd9Af1a3B8AvE6E8XCiKJKuagzCorcY+hZImloUu+MpKBH
pXhdTPEjjnJ3pvVnt23sqFS+PjazJxPwbwV179z9OoU1AdUR1j1v70FcGMUqpZee
dV+/y0RZGAG+dGu2o1gPJumkohJJJxlK/sF1o2MOmkQy5DX5Xd0cQDaXroHxnL4m
V5ZZpTXDkmIB9hfXnRDehjE3V94mXBQBjFUCPdmr9Dzp8+60zYYDaA4dceylkkAO
34ICBiXZN4vXQPlZ7Z8MJ27zjVy+Y19PicfkbOIoJljT7PUBb+mSJjLwo91D3I+h
0csby5+0Vewd5DAJ0JbMzsfajIzen4jiSGDRiIgCum5Mmi+D7rrxC/X1FZeiGqp6
Dk8LAoRI1SKph3hfDIj0Wm0hDl2pwbHyg5NhTX3YAAt+GoYJcmN4e/3SsYiVeS5g
7Z5x1dWoDloRix7DKR/44gyPN2jTykUFxJgvxsUqrV/Fo8VWasLCJmYETrL9xJVJ
FjiBKzF/ci+vcdXF0gOpwdRYiWqo8kFXFs8+1E7wIj7pxW4QrP7QUItHGORdcmtS
wjPFGp6eOwyll7oNxsQ0d6WP/UAVCQ3Ql6e7sDb0MRnxtjdT0lZx0Cf/DDrUQXRK
MR/STdhUahAk3eOCi/Xydvhm+U2IVKRIhmLtPOWl+Egq+aEygaXDpgDlfDCmjbrs
YgZA+kXxI/GOSKPsjJblaPC2piir+cNkyuHo8yv9teRWW4XxZdEPR5y66hTohABJ
6gSBPp0bhdNdbyvcUpvemnEx1zDVF1ugkl66SbrICYPMFhWVu3ramb0+qVCQDYtA
lewIoNqpT3XOZgEb6ZtSrm956XDo0gYtS3qGZ5FU457hn5hb8WFzJG3rx3B9y0Jp
kf3E3vTE5PIQ1Q6jm2grasGxLpI6mT5EDtXkRV1MdNRTBAVQzXMuEn/j5lK9wMwy
vIe9DqMN1VVDx0m9OfHgcxBW0wvwGtnsNYsfnMJv8Ycqtkrsx1MZd100JCnMelKA
tdstGkBhZYG3Aw1hxc5WHdKiyZaJMYiSoAXw7gtRRC3CTR7YbqQn3XlqXHtqBzgU
vgT7uK9xL15CoThcUcEjIPdU2wXaJnBuIrRwsSPTYhWf3IUynj/VmgAO3mgFvBlY
g6VxAz1xgFegWbifxjkRJ/fRVR7ptctK6w3EaHYzCyb8AW+nSfxstbaI/pB9s2wQ
D5L7NPVkcweMS3vlXzcDQw1Hxmr8vmKqGJLdkqWJsUy6RSGYQb1N/xZm9QXJaANO
KNER7k/VtjsonSO9i1iwcPqIwaDq3dCbjDUXvWUrx9dBpgg/NBkhp+AeOyUW+8wh
DEFsvs4zozmOWPmYjMEeSQuNwRhTC73YDJx2PDsLdqhYU6sUjaVQI5HRyS7S7juA
4fvkNPDkfqbwXAFqBXd/9xjPdOj86BGHR+IvDKAgosh8dIn9mtOlGCHQPAaw+MCU
fIg5MVdiPk1kNRkV+HPhrL390zDJ46kmOCdP6DrbPvERR5TpG+HggmO8V3nCCLVd
wEXEWFWu5Fw8Wn0bXerSi3TuErjKCYHmYX4duLOcaeSy5ZjtcqdJC7GSVJkpeyMU
W9ypUMRvyz64ogMuHUGHdG/gfgBoFn3bKERO/CJAznl8Mj0CotgOceN0FYocI92B
xm6xsqXTBpx4o99+VCUtSKT088qJ1HrH0Gp/oFkB7xQVuqHtnp8cVpFyaaTqyesz
6zQI6V8XqBM/OcrpUlJzqoJAMGCBhQebv8UtQOmyqU665+LF6nIc0Rry+/MmaazD
QWalj6d9xkL8sWsgIuxrgv04K8NTqHWwqqRth1MmfcwVcXOlKGwT7cFh9wM4eozZ
Bd8+c4QUxggt8Sjb1oOCKVt51JpNTjlGirXn/cbgGPqE8baNhaIxBkrCLJcbdjOV
DdQMLSNbepPZMZsfbT2P3VvwAnST0wtUbua/MAq7XwFxBLAtku0jzmMQYEXdJGdy
him+HCEK+HcgyEJZ9Sm5PQLdt1SMndx2r8AuCXi4K06r0+n7gMAjqyFHauUpGAO1
59zZ3OhQbT0TBy0rAuwApDSZDCkop08snQyqjOQp5m2ocIXOgRLuWWJV/MhOWcq4
2Vl8ZXu8idotAvZZpWGY1SZgX1NBJGVETnlN7tgQUH3VyOLr1K49mu7Bp8r6w7hN
o5kXKhOutAfm/29TxTOxCT2F3KLryTgByrJVdApZj3J3wQ/lhEnAl4PCKx/Ofj4l
BdgUbtdEynAtBbiRv19jzntLjIb7qJ4WbmD6ahMgDHZ7/5LMooTFJWgPhJAREWj8
z6XaioFVSPxKMW/wBC/EDcDWgmdWsREH3hVrG5++qLkbx5aKw7A1hC8qr8ocEYIE
x2/Ap9ixXthmUb3jFqm5m80eTx6Wpbc20xWzkNM5O0G/AwpNl02mnmEb+sQuaM1B
lpdbK1mcc+rIZ0HEHKiIKM1bEYpPc4kkA2BSv1zvbv8kfeDZ76yWkBzLmqEt9WiZ
q+awL34bBboqTG/xS20cio+wCnXqF/O6nyNkq8zEaHtI29zgSANFwhBh2va6/uw8
xPjVP+v9zkun2iBHrj7k/jcK1Ex/+tMSrKVZhkgTg8xVCozQhgsI5/jcibo2NDAf
wDfOyO2PAtQt2HDtk99Eqn/i2e/6xEFQjEnQZwXCRyRQJUI4QPI0HAhsC8VCHWFC
xHCcM6Tx1ZxV1FMtBFnH27BuxbcgJJ0vhoycZ7K9/Xmm8XRuNjPWDr1v1LjRr6pH
z+nFbdn3cXCyR6druXvzkdLD89XUu6aAdP5+zGvq23iZNu5fEqZSjBoijynNExsA
UU4F/HWRNiFSrnh8U7S1i4IdZFzsMQYfPnEwGaAgnkGyk6Ajzy5qH9qo9T5ynDhS
lVqtZDqqx5VQ7I8O53OYXkvKFQrLlLtRvawMH9fbMEv57rzZ3UxKrKLin06+8sbm
ZG4ZxekAV8dHCgZHgJ3zMzN8CIE4ps+UihU/oY0YpMBBfzPEGyVkC5iemiyyVO3g
cAyMI3cwpJKqLPmu7wsfOr9GLGcd/8z1nrdxFLFUri5qzJLv9kDj49/fA5uiIIaq
1YMJ2LjqHJxb9g9irVFKcxPiCoe8dR0cPZG9NY+ROn5uM/XD++3VC9uMkWOXy0gU
JxiDsuyXu5Fu7Yh4E6x13/CX7yVhpWqLc7rROM+8Rej8iuESyV3J4WyvtC/luVYU
9QBgYANbd0W8doTyN0Y9aW/4qxgAIeeHz8WcA9RzI23j90Y/50ObIBVjjEGPH7sT
Qca2t3DA9aEwoJ5pEfgvdnsfM9rREu3Ijzkzq6B9lh1ExyNAQV0hP6QTG4A1cEAT
IwG2zHvfAoyO8pquWVyFGDqxUdpzhmfF5Xd1eu8YW3TLnSwKIsWUOu4GbHH77uOL
HhyoMONmqcn8x/AxOjeVhwYfPO2OTFr/wFQdyskxsDniqQ+8BmKng9BrBWMaxe32
2vSz9a4aGpzhc1FYkyEXwjyc9ebBphzEbLKWMU0c5Eknz89axfxk/9CJBbz4QSfJ
V7Px5drHdWDaKqruyrFlz8QVGxe2J7K2SVKQXYuyTEQQWeoE5zDpjX9S1N5pZGl0
JCUMUt9rXvOzZKoQCvFyJdh49qZCOM+0jgkDa88ex5x2jej1rkDyIfBCKj2vOoMy
TDPQXao2miyuMpRDp3IPVdEMpMUVlcFJsrExZiNXWDD3/IjRQCByLYa38gRA8hdi
CtDNUl5zTqWbA7pijA0K/mg7diOqheXWy9NTes2RriuNr19Rg4i1Mqhthv5pROQ+
N3NHOryuXKZQO76Ibouw65gTaZI8GQEKptZEOfJkee0GARReYs8mKMKKCZJcKA+L
TVc3iiCZ1sw61KT+YFS3Pi1QD6hyDynYpbLC9PfsUE4hodCBcCjmwZK4muW+X+90
3FvUrXgs+jzedvNCWZLx4NdgPcYQ6lr1HYAykAJ0M5jFJTc/JDKby4RAe8r+LUUe
/+eAi7JAWBtZToQY/4Czn8zCFrlSFAVAnLUoqMT31TZRaiJdR3Nj2YsQ2MoMtinp
NQGF4ScIgi5Jupx5m4QM88jMw7RQnCP12TppO+3gufRsLuEojV/Smp7XCkB0NROH
kFnyLkDWVV8lEmOd9o8zWx66MNPdMOKEcs7hCVVsLcgnZcFSEkJmmzFEReeC2Wh1
Gxh3muYMLMxWdQY93gsF/tWxfxC9injPSp1F0FHbMZWlxwVUhNEAjZHxvIxsNIix
uEAOj+SFQpTRXv7R4a0MLAuh9Pos3ttAVaoc1xcTlY7IEgZVrKf3oy0M1KMhsHX9
7NvtAi+ZLK7AvJHzFzdL14w2z6p4jmo2ika9AoAFtUV8x72//gSx1TJus5VWmB8D
8ZL3n9zk21pj8QUfBoL6+XmOzybWmMj4L5O8FdjH3CiIa1PCfyDLVRywpICqjr1p
/oAx9gUT3ymV8/Ag5LZ+UnjL9cwTLoZGC3cjlG0+4DhNp6IuT7EZfVoys6/BUN3/
u22qRontdC7VvbEfnMvx9BxutkG5YMOviRTrp47zJ56oHuyUu1N1Zx0Gjkar1OoB
FsHwo+6DlAab24N1A11dJKRfeeNY9+cbgdAR3adPUUy4M8yQfGvQ+BItL0nd3yUI
cTv6mTRofh4pHuZiXdQQaSLGvnQ/IwImowcBUwzJJXPgI6goc/96cphtGBVKi9VV
NsppgFNNI+WfrDwZcevf/Qq2HO+55m9t5eBMAWKzVAtfRNdO/Aep3L8MR8YK7yMA
AlTe6JgBhiuWPMlqQUC3AxLHoHtogN+j7UFxPMSQRXu4coVQ/V1E0ERs/JcvxAxb
Q2Vr3MCjHmZ6KTpK0W6FLsenj/0Kj/dgq9iWbs0mn0Jpx+0yXdiSLmcr6Kk3vIyA
yhLBS8vyxXJ9qviJN5+vR8VhoNRaBX6xoecIjtk6lCxZVarHu51QDERv2hUfcBM8
Nt4wFS1re5PoenDPo9/JnWebW4OKpKeIlvRuAGQo16XtSDMo+zGt73ogcBX13ZIR
8rsTA2AS+MGhd6QgtEZ8QIO/GP1eqm6a7z0faU7lyqhO62I0lak9vMfAsCzwt0Do
yghmv0gk5ZKoJ+QxBhx1lKib/FGnujUoR83MGpRK17EWq4mmowxycRA/RStPLIR7
FzYWEhTXuBIai2hHzPSxURnlOPg+Gkj/hV2u1VX+h2G6Hn3JQAytl/KZxfT8hh0g
Pf2NhRpQev1xeeUB9xQD3//UFLvbY/E06QpiSl9b7iEyz2PraNQazJLKa8EPp4Ow
DOHNGbPxhlvr2ebWGOZOfdMVtO91PgBLvJ8eVCiPshLh+6V1eBvP47BVxgpsP9zE
Aem8W/0ii2uK3E7gSo78Nhd2EtxSfQyVS0DVqYouump4LVCIQbcPO4Lo6sPuJOB6
BlUGI8gU5FsOfvWzcZAixqBInoCyjWLnfpUrbvUaryaRZQ88mXn8ikv5FROyxIdx
jmD9J1D/9WhyW2QrsnLV9mlqiMMK5zIVskqYe5ufhrj1toFBL2Mwk4tTZif5CNRO
5F4qL23fSBYaFrRweEbb8wRYqFVv5FrDLxww4BVbYDov7ibCtOuQ8FD4V2s912OE
mt4L9cf87LPUk4jYPh1VPoCNeEI4LhM/3wPjD6y88BednI8bKrs2hZyC3m+BujQ5
0a0IIX6jAzHPKMVvcD6NqyAWZ/osKsRSlS0g5Q2m9MZCYOoM8YrR38pj9yDWpVUj
/skQpjTSzHM4JyJYWH81CsTnVcESpdYTn06D5HYPqJZB/zQ2CTG8++XekuwZL3pB
NcCsOM3Y5VS9+1bkk5e0UBwQOSmVCr72eZ/rtl/sXhWfTUWaHj9jNml+rT2am2Dt
/CHrLru6OjApITGBnAyzYlM/lKCT1QstJqimUgVK3KztZdQ2vfjUSSx85bwkZJA5
Xg4jFaCyHRxWjWyE64H75siczouiQ/5kxIudpDvMja77G+y8R4X/NXer8LfKAu7u
xjtOy7OMXbYGDxBFmWDA3aEZ3Ju1ed9B3zPv7upk5tS5cob0SXxJvkDIOro+NSTe
X4qbNTl8Z9JeNLRtKBbLQt8u4NPCdc54EUuO525Vxuo+lcKh98XA0i+SLFDOlpmw
RSML/bVuUjR9znwNxJ+3pHOuNUAhHPVdqeY93Y3AAFyV2Byixgik/3761txkdxP7
TYM5d55TGTbHQn431mN8UmK0Gnjdx7Twa2W9c8hRlJ2f9MbAUcbkgiwnMUiyZ4zr
HYZxeViqVaXutoJ9YctB3AbtmGyaVfTwcMDo20iKDhGv6PLiiI8nidCqLHxzVfJu
Cdks8Mjb+ZpRsRyValTykwmhW5eSHJWflzyL4NzEWWWYcpJ7aoLahMapNhQzTvS5
2tZimrNt3K8hmh+8dT/as4wwahW/PRT73cK2myf9rq04h3wStqsaGVsnAapi6qMH
tv6wncrxqvp0Rn4UjrmPabORW5KjOq2pPcTHlTdHlfCrxyDesVKlG1p9M7tP6ZAN
Y8BkvrSjsrA7dC9gC1+AA4nx3WvsFclPOOevikYWEHuxz0M15f7ocM+hRrkvjlw3
gglnJz9gYdykd/RYmo3V98ALmaKxCzX2yeAVjrC5L785tFyS+Dwxp5OxMYTUhInF
D2GzHHCnsEZpsCp9jhEp3AAhRYu+CMfQUVDWy7K9nuyZfWNU4PlyznCADiX7WDvx
Ow/I6L0DqJ8gHhcKQC/pzagaR6eX4VobSL3CICELRPwOSYt20K8Gd2xDK2HW90q3
cQmcIgUgp1pL9fNWgBAiM8TOc/LBEPZjHXHXVBbkwqntg6AT7XvQj2DHGJq27cg+
AAovR5Tcp54fgJhRSwmg/RdlQgj4iyGvsIzFe2BmP5bFYN/rdU2KR4/ovJRLiXCu
rXxQea7ANOQb6Zua25grK1frXcDWGyHETzQQSMSQEhEr/3MFfNBW6uwyRVG1EB4B
ucRmKU8xgCqqfm8vaZsAcKqUbVrJ/NE1hWpTITK4ECTRhdTptPDj5E/UguHrXoiR
uxtkwxdeoPvL0YA7Emt9G2dtJUx/EP25DlQurKdn7z3CdgGjOs1zAKV6iFWgFeAW
Q9wKOiI+EUlKuIVf7KEb5AYf0SOEZEB9vX6YSBjJ2YxbYc33aAgjFmnWR1AUw7+j
Yi0ygbb3ZyvAgZZGtKPa5f5K3yayTOj74Xl7oi6a8prPMy970/cjP1aZ0CXNSwlD
NKMWwz5+XJuQbPLBp0sVLat2WtkqsYZAkX6pg8mpBbCSeKzR7KRWNmSF/dEkAfJu
Pilwxl5+DOfEGmRjJNAk1kZsD+hqBVuE/w27ea+HscC3w9MKwVLPH+7MDeEMevga
YqXZKlpALBsVA/1zaK2mpXZ729JQjIy8naFpPa4vWptIuWyBkX926tpo6+0i0lpi
fI6yc/XcSW+de9GjNnrRTsfcnNz8qAaHcVUXgrMleh1o/pt/Dwu6MnaGm3bVSw0i
D+PyLrwkhQ1PMNN59YYtDRW8hvUe2c/BL1OCuZVHQLiASHWML6eedPZk5ST+cvIp
M9DRfujrTMVah7J0md3UkqJwe0kYsedrNbGJuH081ucsM8fguW97OL28hBwW9fml
qxDZNgsRbt9MNCM1FaCETrSJYVo8HxXOKhYusTKFkcy9ASx9EUwjOPtHBTf3IsF0
KQ+1X/zKZvpgZwHbfx2UHlS5tLhEF4RqI/prSHl9Kux4uPncUX2Hh6Ui00UuUt3n
h+voQEypdrJybFwEGuxPoE0lcEq0QDAJRk10yyzhRzoVnhvcOJChENEG4IhETbAS
z1CJod5f6hL/w+ujAX1bSIZlRdZLms4yavfqWnpYKxGWjzQTfO5T1unkBWBUASLf
jsqT0AOqCSk/+mRNPU0SDGmkWmRnu331krmJ08Lfm4jTy/VQxFqKkwiWHdMC4D/t
GBN/UJOsAbTkJvqNH11VUQQzbZ5sE09RbN8kyN+dOkkladi0rU/j9OSg7u5jLOTo
uO6YbnWn1+SYDZp3jegITsbATDIYFhft90RTbGIEGUQObRiui+UtSRXESS+xN1RS
C4GjQj7SstF9CtzEGLNiewGftepj1WNeQc/dZUUALkyN1rrMYEyrMSEC7YPOi3T6
w4Wf45MoQFHfFxK0TMbFAKTTqT1LAXUDBgFyb/59dh3knS0Yo3inw8MJl9/plgTV
lkjJE83nrFlU2Rn2JzWgfLa+i/AAwLVem6wh8IXuRiQZjBil35dWQx8l9s1iHIYQ
sFfYclLbTwOaLjn/K35jDThOzgWgvU+4LLT0u4Ok6czrZuxKMgQDXfzX+HOvgHBr
K7Dhg13VZz+J4jVvERi/fflWDMWWW2xUJcKiIBQARAFi5yNzAoc/iMxpcRyu8Kdv
QR946dDXw4vA641ajo+/9iN7dT9dbd0+w+30fqz3wHExuUuqQd22emNAp+p04CsC
0WwHGbpr4Sq+b7YTrlASHZXtJxoQk7G/0e8GeA9rUQcfuxakH9pGfhFDJemzPgdU
8IgHVsImOM4rIc0tEPdt8ALIfAHKp8lt4l6FpnnPlQVltqDVAfoqPXV3HTcL5DXx
85A/+tnezG0KHi12S9Ca848TyEmd+I20zFekAqX+jYsEH5NbkBy6ywVFV1JPHmZC
yRVrNFtYCod0w8XCvXKox300m1supeyquvBne16MSANSyCigiaXExylaFMQ7Ubm8
lBcl7SvphLBCBMKAa+JHrbslHfsGHt4F8z77HyCX0Qz/l2vM+539S8lpFmWWEDsO
UkEQODlc6c3c91bI0iRF+mS1YPwCc1n1AUM+a3pPmJ9FTFWEi8uThz/RRc70vj/W
wZgEKb+A2rgOyFZloILH91MOrujcD+sl3cDXKp0PZ9bzcNYI5Ld+gU/W80ilVDrT
4IW9EUF66QT2ZakL73FO1GI/61tAY0T8yiioYzZ9RqlEyHliGO8s0fe3NmllhlJW
wXuDV5vkIzN2peVEproQ0VQ3JSbnK4xfWrr0hU1QwhBMARFZq+moR0z/VPK/yxl8
+joz/oGtoTgCKvhpd+tGdwVOTcY6l9gG2Ras+JV49bMe0YCSxZ5h7PQSni6gyD0Z
O88t+Ps31z3dpEOQOyi5r9dzr5W73Rum7GJUKk9CKWdZj+M+yXVroGs++x0NZRyG
y98qHViqP0mFSwtj93Dv6Yh0jJYyJsDZ4K0Z36bvhD29LUKQTWuOX+yz5vmFr5gz
8LEl4M727zXTHrCwQH6H0KyY5fZ6YIuVZfoVAQlSCD++QFIPCzCbfADmbiYqrftW
fEkx/4J4aw8Jn5XvMHo9DJ7ER3P82Zmkd9coBrRMWvECxWScgEvYVHi1fih1hEL9
k/hi314aIPN2YoQMKajg8y4V8YIbLslp+/nUCsJqtC8tn0swBVKgZ1RIlzXBHrqM
fTYZEyeJc65GrpUxF4re7Zen7GBcwlOgw27Fpf2+ERVOPgc+fJAxVycRF+woWchf
uhiZEbGpPFQsyjok/BNQ6S+9H1INXQB4eZJAey7hQB0uWO/QZW69HOCc6VhpRwpN
kYasNkNZJdpNyRWvae38f4BwAxnEJ0xYFA8B5bfZ7jfxK7no6sKu4Nl/EYDaN9d8
vDDi6W00dFUSdByMwzxbaQsEWjQbmaS+LFNSQ4ShHp7cWOJVq59/chFt7Y1cCxb6
2mlli0g1R71C2wrfj5izLtN2kU9g8TctvFuHsXKmPWH/aaunDBocRB39+A+quCEh
BpZ8gtKjy8O+33XoRCMb38fGrfjpcWPsZnbyNpueZe43In5PN+GRomi0MqCrQsVD
TyNnEB1EzaG1gtOjqfMxz1NCz5jWDdBLfqQ/osmoMgb2jPpWL6SqdZK+lisO/J9F
2pHgT/6tG7x6bP+Q8jUneZ0DnNnCetRN5ECv50kJaxBiwYc32c3hFobRn1m3qsZV
JuTVg1k3ZrmgLk8FW/SIR/vlZCIrfKLewiuE9M+uBuPejxRw2GkBhOGMkyLIUNFG
OOoO4WQdX/Tfp3jejIOYS1TOonjT/S+xaXl/jVTArU+7GwD2pJZ73oNACCSQEtkB
pt0WWmrkwbq5j8TpICgKO+Mwpgc60NEZH1+d10bmokTgp4SuZJqemSSrLrZqUhyM
zZvVWLenuf0q4KHlG/hrl1JdQ3Ay16HGI7d9Oj/wCoTPrMZQM9LT/BeS2AhpzcCf
BBuW1vD1xcCuLijVq+sOXreVDddcmdyUinrNxBPnEo6ve44yMs529omPAKGzip85
aJ0JM1KzfS1MoSym0XzXG5U952CmvE4aVf+ykhBrSv6gRb3ckwTrcWzSHO6fZ2JD
ZFPStqz5kp/AnIFKbilKCW79z9RNbwTCrAl220sis07NeuopDcODeKo8Ej5Rs6Hn
RS1qKZOtXCq7ZOXCQGmsg2H3+a9UNJ+Rh7witrUv6R/FokNZ3O3xh934pfqvP7g6
z92eQQHyCDl6d3ogoMWvQf3vMEaBZAn0hVeagoqpOOnhzuzlYEu3zPgKwBDk5j7H
/PCSe6vEZvslzHkxTHwo5HXQmTpgSAO7DMT7s/OnhL3jlC05PFiu120q6YRuYxWE
AAHAK6BYtZYa3zB77dYxbqRbZS91eLaucMAieztAY4JoY0wGZwkaTgpK8wnL8bRx
fmxm/QFt64/qtXugwT2aMWuSECEl+q8xsxjBYuFWPUeOjt0pJKJU/mYgYX5HtVEF
KlAhVpftKIRmGkPUEzCgwO6GaBnTnCQj8qoz5qOlDjl6cOvoVixfQB7iKNGOc2r2
6nSt3zK1UnjM2Skm9wfdNkmQlwXXAUSu9VJ5J8fWm2YFYge0xlg2sw0IG1nYCrtk
Wzh2aIzm2IDGfXqG7CN0O4w0dYragNdM3K4YOAODTPzuJnV+StfDzdwbRgPDqLJZ
HPTiiZObO5RgGSR9afKVBZQS3cAXiEVmM4PJRQyzuJxIMcLkeiBzMx+93ESdmmov
9+aTvpnCEeRiW0VsNamkPB77NRcD9YmJA4sjYysHsX8zmf97b3kk93VJLexVhU9b
tFf/4242hexbKFiPJYQzxnBdwz593sGmA1wdlNxrwNeMngaeV8E4E1Aa/WXKS8uz
BWDO+d7Dscrx/dxCOrnaPgMaQmBaXRpPuuSZPgwWAEv8qiAjyEQmatQrMXnJ6SOt
vzky+2Qj3mZcbS85CK+FNd+saPmXVwto8xf18adr3UyMwVfv+64wActRce6ZF7Gw
Wwvlmq2tnEhsQai4+UA2wX4tGuUvKcylYAVF3rQfwGLVvUg/ELuvIocjzED4RIpq
CZBd/tK/DcZvnMuZgomzwuFtMq7KEmb2k5/zAT0UbjA64aR6SMau8/PD0jLbGR1x
XMyHpEq6Rpa5jwy3Q2rMo1kYA6J/eltiryp5Wn1fYBSxIs/GD1FnlXtmvImzT/rw
xsJXC9T1NNamDgxuBigpUv1F/89fbf+UWLjAYeemhvDk1nKs22sUa+8eT0Ndv9UX
zjQ66WYmCe3Y7DzPDf/Su7rKRonaOf9frfeI12OOPTEr/z0IddyhvdyekzKD/NkO
/D3PRdj50yJ8JG7w0UzW0TaSR7o0pdf1i7ktVgXiGI5Ik8ecNdKDQX5EO7yL1RZ7
cnRHN/7FXwk262koRGs661v1lc1KbjGeW8/j74H3dCpcC1U5977PrpWoDqzIzvV6
+1bqsw7Ji0ouI7I0cfp92JdMslKrVKl11PCWm9erJdVZEN7LaYNmrFmn8ZzSowmi
yUpCSCOl0gGgyxE01mP6MXm9kMbg1xuOe6wzPnTlcFFso9nk8uuxqitvU9Ak39tH
x0WfQdZBYeOMHg4SiCNTV1iNcuikzhL5uwiIQIy58E551qAN7TfZ4UXUpG97tIMI
mWhEhcaaT+7dBp6UNWWU30E/0SjO9q6Lxp3dTogHNgrJ6UX3PJK47/0XDAYTXh6b
52Wxj9pgUOR5kybIumHTcbNNpJo3+LePKTi3FDQkCaxzp/IncFCfStUCqyTROqgX
ft3dalRgROm2Pd1VZcfKhJsRNuwpZNnP+1ERSCaY7cUS8RP3gtR383Muz7wUJjYT
UCUXoY4d7zu6B04IByjEKnvMhhP2RjcWREK6SeQygOALkXvr0Om/j5i9VNmFDLF1
u32a9tdXYqgIBxDI0K54JHokFIcT91bCKXKUewakSMCTI4NJLoNQhQDszxVyxMJn
sYDf2OALzCN1zRCVweHR28WQ0YHBjm+j10zTh4SoR58uf7cJqPRuKmR2kE7dqsSw
UmrQPve04uKlfxJuz963Uhg9Qf0QqqrO7kukLfoquXH7M7grfF68m7t4BA2W3x3k
X8VNxG8He4HG24jyKZRRnxu/QsZYtaFTgSgmyoFJvRxnnPlRmnVOkaeSTj27Q4bq
+yf1SmT+IlvLFjHpzwwLhKJT4OKukD8rHcfSJaXfQQ4oGXM/AkNz1nFXjkpCfaLd
yhoEbyhqMdNC1m9ZMeP5kosFF6AZzhImgYVSQ1OzrjGRSuXk8nz/b6cHWIhK+l5F
MzO7/81KM8rRoU2Vf+BNMd8wrfX1YPLm6hfPl1pmfh3cudT1/StVTKFypP+QxJLK
qeEV+4VMUWQGIy30xhYRxps2FDVu+DMuLTiX2/ovYouq3yvL1pBpr9Ie3Ll3URxx
NuZbawaUzEWCXo3evz37xplheoO0R1uikCgFjObE8p+fkPRKbcTJMg4JyLq6G8Db
FFInQPSMjejilu8eRc6+qfycUvCnEvW5Vmp6EwuRxkelI2lHM+KhAPRduZ/IEZhz
iTkkCJNsrvPNofIfUro23r/i2Olqoocvc9VbOVH/SHGbfP/Rf4f9iiT/V8DTfREv
UfpGSWNHbJ4B9ItPvOmjJv+BkUonGToSoeBqKKgnJHwbCCeAr45OvwSWdMAba5GB
syCS4TfifAQI1cN0aHVy4g1MgxyeCMO8B+SvYeKeo/oIyfgN40pxb6axTIsm04+T
RsbK8j5VWGQlrpqv4tsYLEPn61B2mpyJFQ+5KMIFpAuqOXN3x5+9S8HQ4S3DAWEp
s2Scp+Axkpu2U8Xh4O+uY3BB9Cwf9W7AWwpzdklWwrQhFxxQL9hE2Iz91CFwUA0I
fdWVF4CuZdEATU+2bQhmX7+a2OFG+YP83e6EabLDjxWt5iOx39uQpMpGhcyrbLlC
9570/5Svdf37+HfDYvfKPW1ltd6fESHGfIKDXjcyiVZ5g7efSZskuMg0Jgdn9Dti
DpoHkkaMm9E8ybY8cX5NzaQSErIs/9wSppKgtlrVy0cnY0zHTsb2TE/YThTpmOwP
PFYkU6y59ylbLDOucLGnJlVesFD2L83EBub6Q8k/dpQ0SNqoWeTOpryyXlCF8NYm
eN2fjjjEPoG69/djt6aT/W2jWOsgvzmrDYFWYht0VNv+Ot3NHjPdyggslQDkEAsn
NaVcBvP0elXOa+Lz60XiqzO45J5poGnqg+gSbDHcmw/MumA8wO7VIySwJrP9k/1V
wL6VXVvwrYLadBNQ9r5QtBLCyLs4Vb1+cwJV4NYUcHbxUHnlz96bO8FjR0L/ysfq
lgpmgmeNkZaz93gb/tOurd5fTwoRWfTdZFQm5u8MbQ7rIY9X9ztGujLR3DiKgM5H
jHpXWy2Y5HOzlDjWjfJoTsRMI0702BR1Cqi8Y5C7a7oRS3SHUMKPH9MXn6p+infS
whz7tnrKq3HuTlMqoNAqZDRHJXJyImMZVSvU/1Aba03qItQFqtE1azvindcuAwqX
OpmpPRi4/yUR6NChGnKoD5WGFlV1C0rK5QPovyhoDaansaN/uhIZJR8+VsW0WyTz
x16CSq7BlwwcFbwJBW9iDxoPeAlZkVWs5hGIfO9sI1OEPnfapucdBZa/LGWlMk6C
hNypmjiCsxfs0nxp4LUNyvWzLvNuLLyqdivM1fePB0h+tJWy5WfYIf2eMKcto36T
xWkQQRY1pQ09d1XFj8YdKqknZID3tAYXjbyAI/pVWlMZwbfP3Fx4NG+JrX05W2ai
BWSTyapdC1Ebp+p8C2Z2Ilx49SFedUUKOzokO30uNsBiBmU/ojyuyyY2+/RWypHd
0deYBNL3WI+cdfuziz4DT/+xlW/eO7TRqU4qm7qENaZL9L8jx9poBuouxjeV2KVB
ROPHcpjkU6y3SdFXmYoxQCx+Bl8eYAbPRmdEGUkuUiBbqv3me5BbfKVQnrWx+Gu7
TBr4aWXI0yx+csLiWz9lNi2Q4KpOcG13KgjspLkYhw7xQgXjw/eeRvkvQPV8mPdL
bzH+2syIM/cAtCoyUpn7TSk6L81e7Wx40CxRVCY3YXqhuwyyvvTl4GwEeFYeTVwa
ySit6DcSMiyCiDf0zy/KQqQi1SggV+zxPQrgJ4yJpeGRj99HogJf5+/jJEPU/RrA
xOBfImeAWP313O4lDo8hDF+ErIkokQWIZ+6/NlbQTdc6cKSgeowpWIvxyunhCRpA
hOZmHvPrn9qejnNWvV2exam9ol7DZBkkc3wrzhDptnC1ziIpwB7mafRDplooj2zR
xqGULUM03a74Pxj+RuOm6ykbSGYTeuKdoJ3X7Tn1Lesv0vHkbu81d2rBtHT/VFD9
8OPC8/c79vzkE6Tqi4tDcxrVOvMt7tCmDHMhUC3lEqq4WKIDGjA4d3YQ5jWxmbRS
Yml3uHvmtV8WSBtY7+rCXe5Jk+NBThtSf/ZI2ELAbl4N4G0dsWl45YuVRQRJC8uX
yFJIyfl+ujtX6ggXoDHTHhgoet+EtBtvH0QxsdoWWYF5zsOtGx4uyLkPGEWhW3Zk
Fy/bignk2YAuTDFe1oi6+ew3qoQSEVA33DY4zVSOMTfP0eqhDYfA8Rg3MqoWO/1P
pLaR4EyG0RlIsZdJSi406axvIzdneZlHyqZ+3zIVYST9FDl+11C1XH3HoG6KxBgb
wgas/n87EmSIXBHoQaz5+oCCAq1NVZFlFk3MqNA9wmUVNfH6mtWYXo1gJ7ofO95r
/Jm70rASNQtUQO0uOKKGJn603UR5GcLqjssLl+JLRb7I7rJNyfCNGtPwcprBeFSF
ZFF5MNkGh3wdRo/7bQZQSIsPV6IPdrC852lFpeDJzp7nO6VG9YEIhMTorWruWjSA
9UsjIsz/3I4mEDzlnDReqFioxm7NPhg0tEQiCEOAVrKf3zvdgoAhK90QVOFHzoBf
psREfJ5KXssUY1zvuHEnLd3hLgiGgoc7H70dQU4LFgBz8/L5WzP2dvpgboAwNKv0
t0meejgZtqL9P5fN9ehz9vgtvGIDt6HD+xGbC3BHRIyAvL6J62rgMdjoFg4IgH39
eHYGV0rNymVaVxDwU/ewrgJHTZNxf2FHO3GTJvbeDcP+9heFhXv+HwIU7j3t1dbu
BI9JnUWOK3iZjrKli9gZ0QNG1yaKWAFMzbVFxDznGZKqGxXLqDk5ZM+oQJ6LfBzE
FFJzbkx9U8+AjTkdj9C1vSpb5vjGxOZ2x7MS84EQlMjYdwiQTXn2R555nbh0dK5W
1H1hkIA7ky6DkBZdu9TIhj6fxR/DJuTCQnBjS8nAfNq8n5abEoD8xTli74/FXbcG
L6ti+nyTMyvkhA+pojsi+2sNjEU83e0uFFXXWXQbAD+CqPx72VEJKtm5nZMnx4UA
Nfgl8XUg9XoHo35K5OmVMV5MQIOfhuKJ1vtTx0a3+cJSz4tCB9BBwza8Zm2O1IkZ
CrIcubRlVxfaY/o0yAw6q5oYbNmbe92dfw2ZFS4IPfhkgFF3kal+1fOYoSrOHppE
qp9mGIA2p4II8o+McWTWJnJlLnggSZBvEYagCMRGW6UWjf3wA1/8PGEE+og8GOfl
WP6kZ6oIWO0KMP5VX4Z09iMVH0vwaTntEhxwWiDiYmX822gXF5NlTRmlyXF9itCO
Uc4cFKOMqIKF2Hbce17Wq+8oSZpLSfpafOwTHoHuQM4UZW8PTqVVCS3mDo6Cc9zY
fC2IetzEzavdMg9/L2ook5Kck8g0QkAzZM6N6Spc0+C41WS7fVKc2J6gz3rZK3ul
nVjUmRgNV5Py4xrVa/9qVVm2eMHSogmilDbfPRGx9r/avUAsnZVaCLUM6MUhfkUo
kWy+Pkt1ophQYaqw1Ka3Vea6r94DephV4gdS417hAg6vKAZpjUUHtD79Y10X1gHg
28NUjUnhcFhHjvULyLNSpW9CFMQR2eyGq6oYagScW3xersJw6zX7UIl0AYppM87c
SqUFO95jrTdQSprOvnbA55u3W2ftlk4H/dnLfWPTGBx6KZETGKkMN2tphzYYmy1/
DyJzsgVOgPrfRs5Dum8zsHJ+MtWEjUbqCRJsNIDXLnvUj8zoE8Pxlq3MOucGZAYF
FKsCneGwikNg4flVb0i2NpaUYZI1fpv5R40CYBtxbzjID/5z04Lv1r7HCRqtdNPH
PjJW6S/Qys9srD94supibDFz/X2tD2PSwVLMUG6iXdt7vH20BnzPjrz0a8twdxmt
fDoHT8llsGf1RKGp7QJu/nj6xo2dxoacVDNQlzfepS9Wxz3MKdNDCEX/vWmw2jkZ
E6Y8mMrJw1cTMOpjmyiVBNNtElhXvvq8leSiFTN0IcLpFUudJKRA/sT1I0HM6Jp9
XgLdWOO9IXzg8iGrSEiogTBGlAa20BY99p5+mGdRllsA1Hfk+9P2UieejW7wOaGH
psul5rnhmsBvn+OM7C5p0T60ngCJ3lVofB5L9qJJOQen2yc6VovTueZnfTfDYESn
n9VI0wnkJzbCtmrpaWyKLe6e1QvYIuJI70eyxFChMYtFuQyWaEDKSgn/AkbKdjWs
bUWoyPffO0JXZVbtmaaM1q7cK2Z6b64MW0sltTp8xJEYyaq2SZWW/uaVMlILNJ4F
6UMvXxocSd7kMo2Z6kS/osErA5ii6iqYVl5h9u9COxvgTq8qu+KaAdsDN31HB0Rx
YqH6wM8XL9yBG+b/6rgUnBn6gJ6quK5rGwn9/twbOOHJ/P+Wj6J/kK0oR3u/Bvw+
/Onai14HmkJH09Xu9oEnqqgXs4pOVQ4a7f6Y1Ps4k7csTWFXEywh7/amXJCFdxiw
09FSGfFRN776+hDoKn+ZSeKNaYjrrRAQYtVDy3tB6V4PTXE+Bc7schdTXSe/hyGS
rHwXOWAztTJK5Y7HCqBxlvnbw7fZd6C5QzRIzCSmJ/sv98XeEVb4pz4GElkBbxzz
K4wpXFnUIsa90zq8lj1TO+D/68aIV3+Yf9N2iCKax3l+uRxuxfPVzLUFck+Eab30
q8zbCddtP9kkZTtoIfsK0OwjbYXSddQ4ExNuhNVParAcehj0o9bJDwf4hMdpVzfj
xGbyphE58Fvv3G9tCrcvgKkjKHY+GKXKGG/U8GLNNfwm0wgR3DZx+ek34URcnjzY
/UpBOwstV+1Nz3YnsTZKJMNGKdaEBa6ZJPq+kwUI2ItfriV+rO4pFg5kYa9DZNuF
CXWj5tRkoGNCNC6AdKSWSxL9Q3H9jRlEXLBISr5hpIQ/KzpzlFZEmCVa4jRFw+8/
X2auA2KewHuck2KxmVuGrKBt0pw9AyxTWUdl/cI8cyUx5c9Cwk+XO1uXpntyo4fc
lVbypnJ1mC1+EEPfLApoyGnhIRNuBQXGk/V0ZWlnLkPd+Ad17YYZ4Y7ba950taA8
nuDcb7XsO9dUoWE8XRCayS586kRiqJEATaFE0cX3TW4p+JGttGxD1JepZrlC9oaZ
KHZsV2iNvvs6EtYi+UoUUIA5O/92kcvXhTcgDe5WkGN3leNQ4vjK7VgZR5bM56uT
ehEGuU513Re0C0s1XQZimaA7obGRbMXehKGy47idMSpz9jSApbIHSIijjXeGkvHK
Xh+rYXtLaeTCYTPMZyG0/Df6c1yHOG+736b7xAscDo9Z2X/YIy47K4o0HN6yjatM
jwJf5drNPLjXDxT/AFaEAW+56bJ9ScaehUgfZ6+GYxQ03YYvcxsnCQH3uCP9MLi7
pD6wwe4HzkFig9OJXFI33UKsHLAl7POnAnhWq/wkxlxtybUQuUWqzulCsFn3/KvZ
YbqlqIufE2hPQciMZvndlu6Jf52NytQtghuIe+3j9TQrOUArRDRx/+RWBN+eAcfp
AOcTLN9aLdi4OZjlNsk1tG0NPrO0FJld3Vyqn3QrUG8+d+RprW/KvvT74jtZJWl/
fYrFju/I/PPJNrM4ModGVuwkopvi9RP/f9vT++NBI9udTvnZc/LlOAjklrnGFFDy
qQYGoh28hkGvBtJ7HiasvfBlyhbHSmyz+q0LfPIYlRtkdw5PM2lk/98xjgAO6+LL
MYbfOkSThUqrf3HfIajym8pWTfesUT7KHrLJfH2MZGXeNYeVVDcjxLwNlAsqCluo
44UuTlFCr+G9bVx4e+FPvvUd4jmZKyiNQfR7Jl9qV46cMTVvrciRXBuS3KzMMjAQ
hXacVvn9l0kQLaNWqyIUB55Gy6Hb/ljmUj4UwYJUS/RscO+VSeds38umS28cSy27
4g+lk0IkoeVdGemuRW2apIGsSny/8EJWN+Q0ewKPbNMsVuRaOMj41mElMJngD0Xw
Ocq86rOxq2hv14EXAO32DzEA+3j84BEA2+Jgc6PoRwmmUWwsNAKB1sD/D1GKA7du
RxAVvL339LsR2qNkGkzSu9Ed5uiISgcDWDka1fpVAf4LoUsiZh2yx8Instn7zfWM
YNsbjtPi1rEIwb5QEKCDjSlKxKNUaTTTMb4h99yWQRB/qg/wJjnuAZ/AzJ8pbrzd
kKNf/kAgo+vWvTRnarJrK8day3hzcPMxwf0BuSu9mKgUi8uZohwUyGd3xYUyf/Dy
OBofrjijVH6Hec241+TQVy8u91AsqfVR588vBM1K1lXizTw4RHiGzZjOiUnGR1JP
jdeRNpcHRn7TkK1C1vQfinJ/bJZ1M9+jRcL6sT1l4DhoH7OqSs41z4InZRn8HEK3
EQS1fKgyNJ7nG5kO6fy6pzPAOmyntrF5qw6UT0mkcMstbc/q2EH1xfiVxQUL72/H
Dt6+Ri0uGa4EFPEJ+xE3YlcixIxpnttzzIgQ1gV96wLoj4M11wVBrfXhDpTl5e9Y
r8IXZgnw9LoEF63nE8v/k/kUJ0gxbrGeZXJfE4/LvqXeee/5YzH4dG2TUyvA9nQZ
z/zxLn07xsJFVxx34BitcaTjceIMBhWpUq+u1SoG303sb1jCEeS0/zNj3d+EF2Y8
0lShdFcPtweYlfDMLfYdrZmCYQ3rTrxAIrYFfW15CSXafewqQlpVKOiTsOPPv8JD
BVxcEPFgoz2l0vAJUQaVHJ6bSHwbVsGy3p5hCje/EBSdp/iDRFs5xczztYrzPLCY
WO54lSLc2GP4Q8ks3ryMpH4o/b/ySvN6SQAOz4E0Q4yLXwA+BOv0qiWnMPzE9QXy
PFFcMPHAkUbD94PGw30lA6XZN9+QsJUq8QbSr7LB1l5urgYAT4GMXd3FHwAPqNXV
Ctb4m0IzG8/068GVJw0xXXuUWaAzWEVpK/FO9nnN46TD16N7tjHcrss1xkU76/fL
Nyl8NVqjeH7XKkS+5TNyIAUTBaEZhWvmU+TTFgB75yIb4mQH0x5wE4QM+3NQyHc0
aJ7Q5OgW75wAzzBDWuNm49brRgHhozD0wc9e3Vy51uZjHZq7V1o60G6xQo0L3tDk
4QpXQYNqhsL+9WHfXvZ56zXJDKcHEGG4GRLRCPlVrFOLqD3lL2CjSoRqcaOWOf2Q
wGvLsZCM6R0MXJST7b8OgWAiqA0a8XvBIauca0SUc2c47KDvcQDaRCN7zQhvOMr2
4cJZHxkZnYI95f0JFiMY7MBqbhzPupIUadzUuR8O042prM0FvT37HpmvWmZOv7u0
dvH1ZNdfwz3u87JghITDw1A6lAZgK8uN/lZzIXIiTmOuyWChTXAVDNdByBp2waVA
nN07gv64BNWnaqeEqDMD7njpnc7eRSanSgoRbzNzLniuw6UuFeESCSZrY7SSZZ5C
nhgStUzRKoDZ08A1jFU+MhcQW9TVo6Jdjw+NClUhfrtdWQ93ZsQAdSCZnioZkYKn
10+fjh+odVsTTvpPrjauamuGIpnzLOpdnhV29SB+P4XxZU6SDF297cGxXlUpIg/L
kbsru1n32LXr+zXwIz1Fa5kKKhjEyv4DNgu4I4YEKpUAD00SGoOq1M9JqiviT9a4
CAbVEai95dbbMjbNS7k/rUi1sO09vXzWj3CUfe4O7Vob8Q3+LHz9ebN/Kioq4pnF
p9lVo0UNj0K2yogXuUIm6oPOUiTvpo6fIl0ejIKsiAYePSH1kEkvLDCZPIHLnK+O
O1tJa8osqqvUxriHdQsUCQkyEm2X9/hLDlkC1hXA+hukbThzAjpXcrtsFVOzZRcc
C7GiQCNSyRtSVNobfpY/6dnZYJphy+zZOPQSj0H6ESH7aKx2NDsBIIK0/sSXi9vQ
l2MoyEWdvLXLGKI3ih5tTXB7WRtXfBFaAlhSKmHOdNhxIvAw0oEfarZkDZKZJJlp
9V8wbCMiPxsUCMzCwMarJ8c2RXXZTY5U6EOHocD9rjGzYErrnSLiM7FUVLN1SePV
0KM7HVfRpbjnDzHAfXgDMAsBQKEXXBGe7Hy+XV7mWGIvgWF5jfyvxztqvq0wp2W3
3Z2J8dtpbSVjiTHjr9tkjrOdA6ewv3sJg2RgdjYC4B0gcfzycBhZYieFhVkrwQL1
MP3r4I+k2+5Bk8ji/d4Abh+gvmR1xzC12g8r0F6myORIz5C15HTL+H1IYCeQuJFU
BM8WZsUdu9mhW73i7C98/XtRe11bhznyi0RTaghj3DgGniXAte6OZMs49tbYNZBK
Rjtbl/1W9BApPlxo1CqCr6L2G/k60LVWatrUjYK78uMFr6MKWkXhPXmwgrvhE3iy
NcwIbZ0EV9W/lTt8KYe03hD2ljDOCAsUxdJlmRNkKFwmEqPwlZJ6bYfQY3JmUQUH
L2gdJFqBareRxXtlEJYdOPjdta5VyqnGetsQQXA1muxjHZNuE1a6rqyfuXgZNvEq
RlMjp9LsPL0EPRXy6CxOKGkkH1CywD2andWJJjdHrzQy2d4fhgrv6/xtUjFoDGqR
N00B1jIOI5xyL1RyDJu+/QBML0KxqFM/BziScu1/bRtQX9MCUC6WZJSsW5qXrQAJ
/IdSzDWqh7K6MT/knDD2nJJ0HQ6b8VzodkhprVcIuLz7saSKq9PsAoYZSn98ykHp
JE6OhY4dkYqNx1GXVn/Zenvbc2jC+wH3JPGhn11l1PweVwqqV544HzaohlXHox6T
v4pWuDncwmWhuO4MA4KouqvnUzvtXamzHrcvowxdOpIdKYHWCdGbLqtpDV0K9y74
5XQxDwDeyKOqQ4wNUqZ/kiyumPnIM+DSyOBuu03gQQ/ShaEzDDT6HR0H8GDfkJHb
YoYD81tEIR94w/P8angetn8BZNq+zp61pS3e6FrH3kBLIJJ5Pz5iZTs7qiMiOdeR
/f39KyMe0h86aWjkJYIZqDgyvUpHeQD0nCvDHvMug8TH5EyDgHUsL3zNw/wQ+80M
Nk1RfBC5k1R0b/dyHft39vEfpgDJMsgL1K9zAuihc+BXJ1jCLOJtiVzK5KvYEGlm
25KVEzeTk9dHF7tisd9iEhny5zdKycrkT65GnA+PlDLlI3RO2MaMrUYNbCj+DiIi
Yq/BflKoGZoJjY2MCMNzL3JjY0YvueD38U8V0EqAv1MjhxIhyWL21GaYmosXLB0z
dRbfSXXYW/mRM6SlXejirEEA7DuNOpPWhVk6m3nJBzsH0rEpYTTYo7AgrLnyCmzj
TlgT766giTgtd3+8b6KYufI2FL9TJo7tsdEjwnsobO9y0nEzHqJjJ8Vd6aSN38RH
lAHK8ZVa6vEP5cS+uBC69K2CTVEzoMYsJWje7odD1xpql7mTSuiD8NvEkKdYNCyQ
whU3KA7EHueiiqghfVLVRF0JYYAtJnK3UEOGNe2fhP2w8YJ5X6BFEFSUDjXffT9w
XVCfCg+Z7081j/orllsKzJwxIIgsYH1W/h8CrQnw28lEaILaWdx3qP0xeRQ47J4M
n+x8xLDG7nmMiiUvAI3F8rH2MLzYAOvDBft7ac7+UokiOBr5hIyMP35R6v1aRZ1s
eOHU2bro3kav6ZD2S9U9BYXy5z1icOttMZ/6FvH0bx333mOKssRj+isxprjdxE0i
Pgwlwmr5I8wZf0YQT9NUCkXJZD3m+fCjFhpWDlzp1Qm2eNk2xpSe8gXD/ixpdfh3
70eiyUph0JLWp0+LYpJbE/d0YmzfnF5AQYkWomTY8JsWz2MVXyN4XRE5oNoOVNyU
9J2isT9jMN88kFDx872/7xu5Ebq8QaHe3YjNJIf7xEonX7I30W+FYXVDiqofbNos
C0E7pQIllo48IXRXwx1q9o8G7qMytnVDZEqBwqd1B/ksimLqFP87laEntOEOV11d
JUAk2nP6rm1DQr59VihAPU1oYi03DWGWxKiFsjacYjVvm1cPbhazcNNWK4+QT7hS
Ct2H2PbORNXeiSXsb4T4sMY6zTCQejGvdKVsZOPImBktm5JOHEu8tmkseBJ9D/dL
oURBn4Ud5YppllJAru0UEncF/Yaoy8MiwlAVer/K+OW4COi8vizKaNZi9Rf8qX5A
Mh1617ruIegpgaIfbPRa/NIsBNkB6Bs+WPx66uldXlgLZZuS4FPDSDCibiiAgtMt
rS6snEHSTeH7F8YIe9+98m5nkwqlX2bcjiqAtl0kjn88bqqi0yEIZRJXkk0cqp6i
mf15WpePSxVwpfgmuprC5mj0IKLkrj65fikmCjXWFkgeeUJhMb2PB2RmNFGUuJ9t
SIpXJ1kcAMMl6pmIEGqPbpVhkwVFuCVlRseSeQergEwbobaDVAcmn+QUOc1ObHtO
h+4ChDdv28OfYBjqRa4C2nbRy+uE0I3W2I4Qe5v29RqC+P9l8+Sv+rCB0BJsL1ia
8EmL9xZk28kqIc5LczlY81HquLHevY9VHjdyj7Z5W21d5Lx8VbLeBLznAHFzwt7N
1DaPqjzjIUv+SiK82ZB+wzNE1odsHy2+eqOn4XnAZKnVW5ckRB+7+9bE6ac2CgEj
m6I+mSKPU9gCTQR/tH6AV51jtOyqjO+ut/vnUqBvSklnwYNVW1IAQaqGy+DnItA6
0czBJChICAoa8OXGSJ1pesh9laE/K5Jswr7fFQp0qdtKORVkWe0uy5SpWMYRa4uP
fULae65zQNSbWI0UDcdJLr2wrYoNhwIxOOCoQvm7s8SyAzPXj50XeK1KlPOyagwJ
HLPab0Tddb4vr/ayEgTo2+Qh8jwk8FpXF01xsiCst0GYsBE9oFFb5SrSe0KSbmVo
6Zo0v/Ro6E6/nXm3IabIg5sym3V3NDa6z94W4fXe7WGCmKKCgWma6CY9KASa9wUp
bOx4N0JiZitCmmPmL0JrDVhRGD16YTriwaTV4Y1t/I3NHQJzQjusred6rZ2ScgHq
o8dFyqA0WFrpzpolCHmsIWiPE8gFbX0ymBmOwx8NKEfYfqxCIW+tyUU63Cn6HrlM
nqirJ7kvNxWVt5B6j9O5K5vl5wH7xNgZ8DorGIqNjUEmo0xSXbg4ooriu+Zbkzub
3fPTPBz7ar+Lon2NvYOi6jhu8Dy9c3wqPwIkPKZb+BcI7Wr5ZJeR7JbSsgmx7ME9
TOYLlJQJCohF6HZEOpILoHwmLHbMyDG20DsvRWzBvUwBeH9DKkp9JFqD0Fw0X+YN
rsF6W8j0HQZVDHk1IZ9CUnxtggYI2hdzx7a0RWvw+EjNeVYtMOOJvpYmnLdAgxSU
9YmI9vdwvMX1Q1pYfRvyDPfVqYueWmigCN3wCO9w8kuGvuFU89uny0lXII026eAi
GwCYJh9oEcr/g7OLdR7VIsVFKEktxY/xG2s1tYbvGuAMCoeQmpeUe8GIxdXkwNCC
YdzwLuy0gbZOenUES8yxzr54qj03PziDpvc0GTSZC4VS/JWvMyy+8H2TtGCPbcIB
wCgsjNB2t4rSqOrLzdquuuwtpxTn/LhBeusaYDLmm86sgZTXhYBfupUExFwFbBbj
l5bDqlJX0eZIIvNK5Jx9T15Xu30HeCisx/M2yDTvh/d5JSK+A0aHs6XxIJ4rPmeT
SvEPwhXT+BR3hi0WKZCruTxZa7TJ/khzK5JGnlNp9mSxo8/1T7mOeiiPMwqPlrbP
n/rtRK3P43s7oj+dS+3rOD3WW6uy8qcqjxvSByFed2aNR02bR7MGisKgPMk9BhGe
LFMHauQgu5/NIwn3A6zHia62X+AKWdJx45d1D7rMHpGjEttJaus/Dl0uqbUz03GQ
2PMcRxZnOISKi62CSTcQSarZVI+aMuCU+5wWjdhR/8JzlBqpnzXzKwz73HcGLutA
NpWN9lVsCyadWf44Tfj/Qq2peHcMnmMXQ/CY96MlcH40grp/zyLrHwhcLvN4hAcs
a7rXaycawdBkpUSqXvRmkKT4OCAnkQQ6VWjEW0D5rufDZ60mxqP7SQYRX5iILLja
GApLRqLpygmEk69pJtz9ofxK7rbEdJx4wLxAu/ilYePjJQu9+g5Z4/kvGEB8Bi1U
GY4XhlrAnhrhA4vVWagNIoZU5RHpPjZRs+jTK/0KOAknUsHNL146yEA42bqtx0Ej
Q0iCrB8tvcwYhQslLaHlQxHiKu23u061XCCZvNSbcnUSIldVY9kDgwKMzI8ST64u
znybsUmYxuOPpSthBvKRp/g7HXaBFgAQn64wlDYb+G8PywTZ41iieyODJ7iFisxU
uwwu3Ja38WJvy1Lr+rKXewu4tMX9nPZ2o2DgeVSgvEVyhYePtvqfBQzRe+jWm3+X
hYYeoavVcyKW068GwKp+nAENsEcDe6co6rASRSwQMn64fJ1RiyNr2m1slgqp1duN
AyGP1nIRqnLDnw760jK7i5uJyaKhmI/3KJpVhHP5YH3x9ErDAulQGqzK2PJskqZv
3zkaGT5lQ6+e2AHWOKaR3JM3WtXb5UlvaJ420qbifJctA/xyKHiuh4EFuevTQEID
f6LRtBI2f8UvU6cHoP5AUeKAUQoGGEagolYgXV1c6yJhxY02cesNJXI3uBNyrpl5
rYdImvaweZGQEAPIws1J/hllHvtDQjO5DCc2XZe1q9TQlCvPtXVKWBYSDZ/mL5zW
pS5CUFE1Dk5vczb6bTJW8Ho7eSvKOuRJJia1dVYUM7coArJUuN1mlEcok5WADYt2
SODARgV3ck9g3jEHOribFoctXci54hnBHsGg33HpDgb3xi8dZ6BtVNYZLj3vrWJJ
eiiloGz/LTkVSDW0/vTDcin4uoeIWfD8qQqyCjJYJOpFoJ2ZR3fR+CHWNKUIzcNS
S+BPqj08tz8LDC8gSXpFfzknurbpXfru21ViZ7S+PbotsuW6z2lePsoXCXQ9c8Yq
jxee+IjrMOHdsRD1vTzL+S2qEK8KcEAE3rJAQ3Tj36RsL97c0oM4fVtauS3d6xVn
bm6f37rjNQL4pMUfOzK7mDdOyq5hHFl2ubKFM2LqGSaf9lhyE/hukoBqbEDN6HNS
9DP7uk3Gs8mR2/sXUxM3aTowx8LZak5rO/xoNR/TzZrLRfkjn67ooSMBEYTaRNvl
hbq6AcsQ1GRbOXqaBwhwdk0aXccjoF+lkSMDdEechH7hVgiyogXthxUPECfohgW8
QRq2wMdehEjiFnFqMSWfGKvKzwkQmAHhosDwrc1V/ljDryMjrjiuK4O6MxYiVUTe
OaD8rSluMsCpRgDttGUP5jEMMnD2k/2nKJwrTsO1h2NOkCBYNBu3va/RdRuu3uZ/
exD8r1a+zUo1S2KiVPo/7ktlcF5ZRtSel2pi6jDgUKMsdcScfNzasu55Dphn45Hc
jjaU4TFlLTVC8r4OxqeFDTr/k53KGvVtDRf3k1unXbInkmK9xzYX0QIR+JuChUIn
vGviis//ibgNDzJ5Y+rDVMaHeJ4c/xhAkyOlu7zu+Oh1ME4pFulT23u1UETmFWro
YHqLK2mH+/uDRDN7Cp6GLN/emkxUbc22ydp1d0DegZ7Ggg2YyfyW81Tz3N6w7nsm
HG2dvdJISMrdeKmx1XoOJuEgsSaaj6BqFkyXPlstZFGajxJeJZUutI913axd6+YF
aOJf4lDMaApFUFLVGtHv8J8hOXRKHpjidiDExPR+iXm0Msstfdi3YR6n/Jq9OSkE
UAi77sralG+Z8ucuapbclPQjD1eus8CfhoYaUqrDNDB6fXnjorFDE2g6q+iQV2tN
q1cxO9K4L6Um2a1B9Cj3qqbzmSS5X1Rwk4OqT6g7MlwjdvhluDnN8vEDFLxD0YH8
XwMkia0i9AwWCp12XyS/Ky41P9fu1EMxwDh7dIufNgaLAL9YPOisKdcNwJuicK8s
3lDnmzsv3AQx29X9f03hPMbt/W/fvwgibI1xih7BladXCGpR105BymKWv64AQFVv
ddadw3RMe6Uw7JnUgPVcf3iZCyFJXjeTN3Jwtp9ch3hheYZdT9/onaD9q9Fo+Umc
Qf4HDX+0hqLkg9tTXrZnSRqUSbfFUTek3WvoCkLzs2hoXEO4R9GihUibXsSDhGN+
ZXdMsKfPftwqTlO4inkHi+Vnd8GJIbFYlIHOEqoJp4Sq3HiZ3stTUpK5dhsKSqIC
UzMrpXpFhYxJkwF5SrPaTJAwZPPFBkxZ5qNRVCNLN9uLpjbIFeiimiZrmenNFin1
E3djWuBcXgytxxS1ACnasclcOZbkZaHo2ZBM5eWl6nEW8Y/2eAkfsoQqNiCvpWQo
PHVcYTk0iJ9E7E0GEA6xTgvAXXdLttFOXta+OnR+0CcbYkjsqCqwpWarZpUoFNmr
czvfWLAeafGEa3LiUO+X/66Ob8pSa6NByJSsf8ZcYmZmrtT4drc6juTXe1Fm42eL
ZpJWdCbqENdhACYvfE1kXZ/gHuR/Y5cyeLMVvdMpJc+uDs9r2+a7EXJSI2/ortne
usgMvKUBWTiJIoOoFQRSyOSNIH+7Dk8wDhxf36QfCsUK8Ncy3fBDUO/pXnPsFd9E
2FQvw5IUtYCyrdpw7bW/9f59cmYLotTcWyI101RQYJykSYxW3E4/WOtiaI9Fi7PJ
Dtmt70sx3/m3MmcVoY3fsqjRhorbqmDOaCan9L6qE2c+24ronc9zZ01FqRSIxu5B
hkNbXW1az/5LII0rqwTZrY3ab8oWJ6gMvHJz0JOqvXnpTguMJnQ1X8upokqfQqyT
bui2hmeZeP+d6aEGgGBSAIBZfou17ChLmFbQG5UjDTLnclZBUGmRK44VSrEgEVzT
xMeHhvvVpb+GtbmXw+KgU9tJJ8Leqjwytr64b1GbxJZwdcf6qTj46S9Pd91GR0Zx
FtQhatsYm/vfZiD1VaJM9tb0If/k3zLc+Bd6Gv8w12c/bjmTVsEwvVbi5VrGYStU
PEjGsgmKIZ7KJanjeWAx0zJ8p4aXSP/bBAdNWB/xQhz+l9d+p01qrtYbPydxjLV6
HbALnoFZWMgnaNnLXg7+FPwLdboUdxQBYvUAOcV51DqyNOCyIScwi1agEvdrmmvG
r6Qjifk5mo5A8c5yEMXkI3WF/iDSnH/qX3XHGn8cXbeic0e5SwFRhDrWeqDyFacy
6y1ozxSMOO/hixGGg6ineSNfx3XrWfAR2Yvt9l33GZ80+no3Bdc6b2M3smTc3cSM
dwnibknTyLNoVCaRg1H1loM0YAIJOKeqUefo1HiNVa76YOlw1/dnpbFN/zkX+iZ2
Nwmiet9YhGcD0XYeKZtfFY97Q5w6NWbWuNhQ3i4Bybj1eoAxTZiMDFE7QtV+ct17
cHHJMUWVWAueH5jKYR3KiMKC5GPbBoU4aHThI0sDLTus3kgh5fAwlxFEqGiggI1f
R1IOwAsRNHwV34RyAOBvI7jtnP5tBU3Gmh9e4kHzAMohLtbr/aw4wyvLi5AiEZFt
+NHx7ywYOwLztCG0NzFCys+RbY/oqfNZCwoha63Z6dkR5qZgUF1L9GBPuBKDycPc
X1B+d6ixzDqRpMph5FEK0U/zHZunxVW9LM50uKHrBp54oipGS7mIbTqkeIL8jQqL
krkwlIUnKlsegIYYrsHI5yBB8iv+yXn9XtAGM5AC37dStOxcCDzW5+8vo91ifzjJ
YyOtqsqRjSyuWQThVef+wOY29F3+F/cGvzfIiy0w7MXYp6ZaX0nw6tGv/auDi6sC
WYQrgDNfq78TBjO8QWBqkPWhgk2DKNwWj4TPBhema7kG2Pgj9q/o+Go48GHvSzxZ
StbJ6vY7r2JSQWLD2pkqBr/dO2q7F5475uUTn9SVQrpM3LalwgvKO6RIEBQgycxu
O3/XGUSNrgNMT2eHI6ZDvZF4UkHv+C+f0F2pcUdi6PTIdimB9V99TRmL6HFLfE46
2LB7WkV/MXH5jI5ben8lGP5MNZG0K3xXWVFbmQdSf6+kBnHv2ncqqQyvNf0hE2wS
mf3l3o3+1y2MLQ7DO9kPsFO3lBl+ceoymdvkZnSYRrRv81FHIEHKPZG11NO7xZ8d
NCwpN/cVPsyYQ0oHZDe1ttBSaGE1TNZxOS1wh/eODG2siX/HhNhAe5vQY8YJEn8w
mTxwGpwL/KfWqoLeLESz3f4PsHoFjo7rjE2EheZDoHeGt9q1F8onFrqDzxh5/RVy
4YWKIx+FB5qWRZs8605xxkkJG4ipCuU81ibngDfa0GlNkRUxpeBpsLv1EC4TWPwB
XH00kbeaBZbmPrAC5J5xjs87ELKeT/D4P/qGDPK8ENU1SHrU9BMYNrZQhhoz1jHA
WEZs+taB6kmuN72qKZJLsdusvsufl+tP+msdTyZK8wtUEj0RIxVWH7a6rOf2y5/x
yepC0OsrsZLRwhmIYIPCYaIi7G/NxH56u2LUIYt0vNTgCLldMKyBB0EGo0BKFf0v
hkDN1+h/mmuFPjTvCzSHwBzYX4fRaxivHdHgxLrweU71iAZ7OOHIzECfugzGO6k5
sdCg0EtvGq8s7RWTPeQdYR3PndNQY+4kh1O4R7i1V8Jjei2DnZNuhNfOKgwhfcAA
8yeIt9IMVNQE3/OGtKWH14xRl5BKJ4zKOE9u9WvVE93SYHjcObFZJXoiKgjbLR8p
014ZnZ4yyevnr2WdPDFazDUOeMKl0RVCC8jI1uythLgZFfDpRL9CJMuJsstbQfCH
HPgz6C1lMnNadVLzVyqRVQBzXSwFw7HvOMlkcQmXlTEy19Iu5GLNHevBLrtBKzPP
WAOH7ih+zcZt60PIMjhZOdfBPjQ4xyIdE0EpF1y1gpXH9TLXNBzkA+6Vrz5oaKcq
4P/yjJB6BDEDcGgHq2Bu0Ederwrc/1uLc99drGv8hWcXsmYItbORXMrnzM2azrJd
0GJUzn8qOxWfb0eBHkhYDh4IKKoXQ9xTq7h0+Jb0J8yEcRGQaDDzLCkZKn99uFOJ
JkayD8oE9xWmBkIIIorRXKpjphUUaw8AsIy3mj9dfykplcdCA40EDZdK/yxtJemm
m/5YuhbaJLH/OpuWmKaloCf/zi22nWTNmw25uD91BbZQrBOf0KufA/XLbTzkAVsY
xW8EV0gqGMdVpJUOprzY5IwpyYAzKs2f367oVc8A0UBi344yeSjhbWijW84R7W7c
pU8zZIkiouRy7Xmz9Zyswpb2S8Fd7P4xNCtdt09cN8D2mrrY9BBKtu7MNRTqsmW1
pNiEgTqo9oG/ITQqveU8bdLYNqaY744kCJAXGUTWh2MRATx0BT13JNsUlAEl8/Vo
42H1NJAnG6XpTeX4d1zdAy3ClTe6+5y+ZGhMoZw/aLVw7b3bFRTG8oJ21XNk1w7l
T1d5UZv6z0mjb/MPWVmSRSXP2p1K0VAg82T+b6dToG/e4EOZ5CaOe0Ra+QlM8Ujn
0xsa0jHbjJKVjZboU08tHuKyHP75vYLr18IHTCHDCszGwTUuvew6XvGXh/qcX1yK
47sip6XG30Kc4Bai/tylrMxTE7q3M52TpzTNlvQE3VSVei8HWw37k2dwtCI1vd7T
LUM27MtrGgwcrWshfI1F7e+AesDjjObQb/c52A48IF5MWbeEYAvPjn86Dq1WApRs
nffPmitM4y1d/ZaDfP7u/X6Wuc9qoK5GdP+4phLN+keBqxrL/8AJBc+VBvIxA68j
sz5P+4XngQpDCZYT5vgCDc6exum2mc7jdMAxEOCGroaBkXff5mxptMBx4zwsK3k3
+HNaCYO4eZGCGhEmUnHwQwMmEYuLVwiJckLL/jO5jyZVYeNh2ddOQdzElGQH3IP9
TnT4pCl34IIX+vzR0Rqe/ifSeZgAAITtp4Du4fKt8xtNdFPtTLdA1hH6BHucJjLf
Mxx56xXtN/ew2pH9Ve6fNgQJdVk3VSs7sKC5fZ36+X36qO565WeaLfpfi/NQpEw0
156a9FXrbq/+pe6pLAH3ysKUTddlyqe1PWQPDQHNCIdcjySeicA7yTK8CtyLBTlV
/4LTHchRNT6RCI7po+/auoRyGMOcdtGSsANDuBd2cBlBS5M6fqjlKORLCTaVxnhs
eMorYaYExHXW4u188qFFxjQtxsAWl4jR45/t7h4Nh617z+ngU0xZ3Smmw5MsIC16
PuBHCXLHqQX8TbdSmWpZhaE8IrJs/SHILnZ3u5q8BC91mxVz1rqE6fxZf6p6PHTW
o5yE+F27dfgQ9M46EVHiE5cCKbec4UGmZR44CMIxtMXgXf5UoLtqUzRHIxC9aKgR
Dzg2IE8ftZ9vlA6zD2mef7VkMh5xJnR4hnJeNKF0XcDsN4Z0BQTClRn+sxSTPtKh
UZlGhd17+wtpNDvIfnJMfBpkyZmTbkKs14HpT6ZkAYXLN0AZ4AD6hZ1ms8NCEfXu
iySElEeUSIs4OlPq5vUpKiPfgykTNn4gUUsLXjt1jQrbCZZxpAmcGnfp7pyKpy7x
0rbCQj4g/hUWAt2mFQBr15urTN2R5kfs/+lBEg5B7saluV6y5LPDhVU2YJb7doia
y79RQSpoV92VjfPGd3WLAN5pUQ2dDYtlqcW+hnuE8bNJ56AVu5/pq8mkc7KOKtVM
MR7YNg3t1QZlIlHH5+FlRVn0UOWiD6M8JXwpIw5CW3dq2fwRk8a3ZF7/OlpB8+4t
7lieD+vp+q7+cl0jXmXfZ3LpZn4/irdWGLSys7X0UeFPpt4oi+rbrTHlmWSYpqjh
gwNvJG5MllxPDD7GYE3239inF+6+8qWuSWkrG64L6IFHiB917a1jYbB0oQGMoCHy
zC61+ZyhEWMWVljBwN5y2IU5NcQ977Jb/DQwbULprAeb1xsykHQZJnOTjGQ5PhMO
BzWZA/OHjqnJSZ5WDvMkXa2n6n9/iUnPGr/d3TtkiA1TI53/EmviUOwgZF4W7+mr
8wEg7/lKqlSUhXSWdnv1fVDEcHhXJzZYKwIR6dbmBD4=
`protect END_PROTECTED
