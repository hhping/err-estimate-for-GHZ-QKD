`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z07cJDD9V5uUvpF+E10sX8hwFlO4aAp8dWxCoroC/J9abHoGds8cF443MXkmj997
phrXTyGMiHGZUhUktSpHATKezLXnvcS7AYRUGsPkpQOxTrXjEErfgUN8LPN6QWVW
DorBjV4BpSdbcQS38513Lnijo1R01Iky8gJMeKTykkiCNtcC1XogvcD2YGEO0vln
oExgQHy3WKTnDTp4UKhlNmBtjU+Da26jMY99VqI9ErOqYiC4tL9QUvrobSDc3gNS
JZb0DtXIQ4b1gBbuc+2iyBV/gUfo0K9meL2ZW546kcCfky2flQvescTtRN2EUV3m
T+qth+ZpdLTXYjdwsZRMkYHu0PBmUbLwkUyLqdOfsDPgerUyi9BCgi/JC0RAiDIF
4lzMhvMyzzVmOiB5ycdPHXOI3kKnKUcF8jkoHWL427PS7oWNoyDiPqnfiJ9FnaBs
l54Y5mqU8AJyD+DAbyscHkqxg9onqrSFl1lFqg0RWLHgxhQHqZNvpG4/MGruBe9b
BD/cZ80lGQ2qkkvydbXgQYTlWtYIE85baoRoyuxbGc+gtwYm2la8DJ+78PHNWxA7
+7JRvC17OtQsK+TLIZOGWwy6FTtaSkgNx6t6qpbUvbwacM4YNLyrBf1RI8lJLsP5
LDoHVKrZyMESl8dwISd/ZLcDYH8mdinpMcgcprPEhJ2dtYh0+YTmlgtSvRSn4hIW
gNGn70VW5fSqjPafgzCLmCV68zYcYa7hWrmebmm5xIzTdfXNxJYjZqwGsVfszzRB
`protect END_PROTECTED
