`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ohdAZeHqma2bMvL516pPdvvJ0U6TB7BvkoiZ6CeszUFg+/5pFcpX5WuB1TTVvjDN
zpT3qkG1cwzOhx0/4UYlwSZwxqq/gBukXipgF8UCVe5qxHPEkIcBb/i7kJxgZzt9
6/R54HtffP0bEldXdWtl8WCb9wB2pwKHJL5AN/OuQtHTnLu4kvoOUVTmFmng7VXI
wqzYpH845ckQ+6fLzBbntjS5pNi3sFRDrsXR4biBsvEFBsUf0+1gFvaYC/u7LiB7
SwjoAUXZgqOKSFDrxM1a8t1kl74u1OYfsjH1Q1wonc9flOmIIGimjcr+DmDk0sRA
//XcvXI4/gI89HoZy6Lmq1Ncw0HkyN7q6tQzXz0tVc89QTjdSErik3imXe3XtCrD
VWDehdPBqTiFIumn+ZM2PgioDUgeASRdZpJZTzLwGwwosEpMBCH/iN2FTb9LP1xE
NP5bVo7yr7dQEqMD0YXCpbqDPGEGeE0GEw7Nj/3n7QbkVhw0xGNRUSmpw9EE6NO5
v4jT0jJn9K7UNpYbu32MdM/jhfVjI8qILR2L3N4LiOIgudKbDw6HKQIHjcTXlfhU
VU6FDSoazephXZlhllTmrqGFiu8Gptm56gw9yxvKAZOtUlxw8FpY/4b1kZCC27Wh
reook9RcKCtA49rTC/mx78kFCwMjac6Oi6Yfx+7XUz6gJQsZZpHLI+IJWH7LlWmz
5cAS0fRi4xtKh1eUcncXb2eSexKto0fa8I2+nvoDQkiUeJ3dRppkRpWv8YMYTIOq
yuq5yumjPz1i5eOgkQgQfhpJQ8mn6RcdeflKSs11qadF+V0LNsTl5pMMk4Qq8qws
bhokyCT6w+SFfUbNQ70SEY/KPS2w6pgZ5cqF5pedreK5TWBO/sJno/izdFGy6ezL
6A59vp25wsCOKX4Y2xeBcda7gcwjpJPyhiQXRevm1RWor/dUAIr3QHWlAKHHa5Kb
TBI3HMxh7/tlhteFStoOFiKQSbvNzZNMKcYSXG8cThF2hJqJp13KXWwqQeMKdfHn
5PitsGKbqzaajmZHLr91QJjewHNEaDn+1flfxELYtRHURNUPO/GbKI9+TL+tOCJk
V6muhT72rSuwfGHYkyd8QPk1mZWKEq14t1T1VfBvwcVVZ1Ftui08KE+2Vji9//CH
rq4fq3IwIUQL2S/Lkkd7WtYgGJXctiEqvDvtR43CmHmYkwq0/rS3MDqb5lEMD1QJ
1TWJeeLLDQcM9UYAVHFS9cgBXZTiMlYhpwZNHIrrHsMxMKP81/ul4uw76UMf4b2A
JsPu+HpV2uNkppvH1+ZT843exYj19tCsKKXn4/xCnaq3nnaPy0Wg4RcO0K6m9ZPW
7c/m70JL2LZgjiT2cnK5gCtZdQ4Rggx3fHG081wtsHOLKrt8/y5KIyoQIqlp3cco
XT2g5DTWuuC0l6DyGK8Vuw/H7em7Ky2gv+XVf6TEh4rfxkzqNhCq882G5hQDWQIz
QfEXWXwP8mMKyHL8jfKKu+jMP6qrle1G9QFVQMLwfXfzXBI1a66UA0YV1pySfHPR
C+sJT3wWVGKkx9A3yB25Vpkp1g3C2P4I+/UYxakOUfgd8dBAnjMmmYp+6bEdSbGZ
vcXn/l6qvrIlIiBgKsMeGpiZ4hstrXpc8CmcreE9AgGDboPnVBFSs4Jx3orQ8cdj
chORQWVkLRWPwBXSy1TDJazzhRxBHpBEbgDNjckEXqY7rf8bscPp1MdKNPfKbaOG
RKf9bQLAGKn1Yc00AnEkHmwJiMgggPjQl4WYbxu/4q+nK/RHkH84kRDa0P011tm0
FktS5Wkl47Dsgwt/6gJrTaSvzXXWhtJx+3NC2TsOi+CTOc9c7FqreOPpTZ2BbSFV
VsTpTf5q7jYf/JadEnYfakvl9YhDBOMKyiZyaAxlU9LIfX1SQAAKlhEP53vplnLW
ZHGVheHdSoP/5J7G7YKVLGfCOC0rmyNFyEHhGCV7psEEveP59PU44IwpU3YijAd3
Eu/mb/qSCHZhB7o+ZNqDM1XxI4kdUG6/9Na6a+pD8LX5rqfFuDiqoxCSf7d6Fkj9
rRSJpbx/7GrwwQrEjE7KL+joeOv1olhpI1rHZ/APS0937D4vly6CkMB3Nvrr4MF1
9LIiHZRNFgor3jiG+fFHDtnZxgvSN4ngN4C/BCMUtj98WIECS6tsFJsmtvIq8q/Z
3tZl0K5g5FYGhdDiz1tr8AKV9GE2FwYZRXjk6gOR6XOjf5xUaQoJRTTxoxMeQHGh
yzxNq+3vvwI/0ElTTTvVKQYwrDXXef0p0tD6a97Cac+1Tw61kwiR7oGEjM+9XR63
gcPRZrsHquKWFaenJ5ssz68g3khmFwhwpqhiCsjNR6tNmzGFm3spEg0XCbhOZYoj
PSrVY0nGOcZMEFYV+mWjQrRy4j9GzP+koXgt9wqukIpLmf0+gP3ApaiC6DUGKxsN
m8msmtgjbiYnFKl0s3SzXl0pReFesCR9yEib5fdCem6q4bv4FSIwE/U8sXTCM4Xj
IecixxawkY/f+HD2+yLd6nh1bU73804cQWTXgBMNR/76SWB2nVuboIVk39bVcUzW
pfeXMsWDp6wasGrW2aIts4xAdDhuMoKik0DaqtiCmu2HzQhsJj1OOy+FZ0deqPcK
ow/J652XrTzNR1x0X4jWu2luNE5AdyHtr889i4Jwc1/JVS8ie9wQvenZjWSZvYSM
Jt1//tLkT5SqChI7l9YDkBYYhNKACj8emgGZ8aswgI187vqJk3645yKcXEQyvaCa
Z9NR44Y3r2YcU+iCTndPXkmXf4QjxS8HANApi/C3r/44uWo0B1E6lS0uHJJvG+v1
NjBLbjkUD97igsDJdK4/3WprSTWnBNndPeAS5ufj9RGXync3M792Lq7kqcoe2Mte
gXqPSl0RdlVaCpLk7/PcdZk2uOFDEpZG0O2CBhNVrQ0+sdgoqXG+/d/qXH+vPXlB
IEf+Z4A9DV5KMfNPjGUqIgiMhnZQe7Lu56JxQoxq/L8OkbXO6w4Wei1r1Mz56dGz
`protect END_PROTECTED
