`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i9/wWJAXEJA4NLEqul0WvT/KWeQgU6SMymeocXB2bx4nfx41ODKrE6lo/E+gOixZ
EhJjCZ/U1z8Y9Ugeh6NpqC0WS9bZC4c9lB+2FwSdsaF+lVTNpZHDL88/ufQA0AOl
L0Knh43H0ywbXM3tNfpisvHXRpDTw3BEXTsH41iVlN4afxLZCKhK1PV35JEC2Z20
+z77FSTcDUBIspSXlYbEGDSbt7jgA8FLdY/vSwhk69rHtqLQdwsye66KY+EA/ovV
H9gTykvREsPw9Q3JLRr1KKDTxDZj4Kh2T0sfwiEdEvyy0zt9ofNpIlRUK+iyzgic
g292kqMeSS3nFTHvK7pPBCKPArAWH6AeFHeKobM3B9nnCkD4DL5XT3LMRCyRW0qN
YjwktngsUkGVQORq5QoWuWzngOEHZhk2nUf8aWLkCs+60iCllkrsZAgGTniFcrds
PUpotyYjZqRbwi3krxleuZ4+srEqp1PiaOhiN7rIzjWkRK+vcC5RjyjfWnYgnMJk
0O0FcJr16u2jRCwEKovaxNgA0P+RL67zb3sNxi9PHIaBbv+2cP/iPihKhuCVa74v
qSW5qkfNT6FKXqVkOMLJ6/8J2M4Hbv51Ved8zOEH2Hn9085hcTTtcZHTZLj6Te0N
kzPbkOm0413HCv1lsWWwLA==
`protect END_PROTECTED
