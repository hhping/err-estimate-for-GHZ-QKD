`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U5YcJXP9oDX1Ui6AKmVh26bi8KUussG4o2zoldpC0OOXKFJr0VXeSiBbd59rG+CC
32TYElkpX3grfZTtlCT+0w5lfpYkPFdJIcx6Em/0nX+3nTukrcQnm7c96xe9QTRm
F635AnFGNo1qObqbQrniot5CkdG9pGEB01gcc41kcmkFfVk8knk8yVC0qmf2lzgz
3Y/C3bGU46So5ddqZ2ieozSu8OHYR59G6GUXNoEk60Y6bi52XAHuiuL6t4FXvUjb
6xgLiCYJKn+QDPH3AJ18xxeV3CG8MGIKyJbQ2l+4LL9+qrd+z5SbCbkjUJBfhDnd
Ss6yGrRF2dhf5HX8inBobjnWDugkjyRwGT9S/xLOgCQz4N6auE3mHUC0JyT02AA8
Q5q3D/qvxVC0BKfovb1a3oakifn8XUDYdJA43DJwm4/BtCHjcb6iCt/EREtPVGKZ
OL+KJbNYNfnxR66Uz1nGQ4AnKNRL1iCeSWkUI+22vjGQLT6fO2ciTXmLKxA8R5Td
QtTKDGYoN6L7fOvGJ60Ej0LpY7RW16F/ou8ElwA0T+8KK0o//fl+kd8ANz5m+TMQ
YcCjaNywOatyVaSz7OZ3jh9sxo6ig2WGigg6uDvkZKCKs+EXpKne1krDCtdaGJyX
Ogj+BtEXdulKZCppYDB7sBK32JJCR4NCSs7fEYfcAyajfGNw79G6wr2EPZuRe6Ii
W4HUb7vYcwUXwG/XYwArPaMt7N6SYyuDNnqKkBl29IntgCYVFH1QQR5hrj1OJDD5
I2d9v4pshT+fFoTJnIBPEwFZMaIgt/8ReJh4JgeMyUcEnmMOFY+UlCR1OmlRXjwI
m+Gz/vvq26OYjpl5RSVTf2daOoRYQ7PRo6NnIyTJPmShHR+HGByrQs4OJNP8LSLb
b91BRlJNZauQTu4hPHRpzg==
`protect END_PROTECTED
