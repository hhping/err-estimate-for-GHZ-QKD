`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LohfFdrxI6sNPyz9Shh3uB+pWWy5JodkbU3f/48UJR46WDKeksBxekVix6kjnqo3
3AXrUT0Oqv9Xi5Uy5rCnTWjUXc0x9nP+kDctKsCYsEQdgPaKcp4AopyZoeAkVMkt
0ILHmbmVrrZjiuhhxxF728kgHHDfEJXgK3RDCyezkU45bzf7Rw5CxYmI8c1LG8zs
b14CJ3A3N2hWA7o+Kj0u0s/sTihoauE1taX7j0xJLhBPAppmy6PH7rctG/PK5cSQ
KkyE2fQud4kWWKgFCsl66BurK8rjik7PEpx26Nk0OFeoanp+VgqdHGiwtyH8OfzZ
KNNdlR9e25bQScnbAIoCVDKr5dbEVPx3Q1VbitBx8Od4/VHwzQV2hx6syfzbDZ3F
/1zr3Wy4ZMhvNGMRexWxlKA7/FZUTbPiAdqmiQbAct83+1/PME/4ZXZOHr9PeBeZ
bpPPPRt/HzS4eA8f+ZPqW45jm+lWWnUCmJqToZQZJXe5aboj73RPHX5uE2ZmeGVc
nIH8eTFW3OQ6JXZst68bEJzBnF2SKPVnE54f3+h0ZP/0KN4i0CQexWL2ddEP8JFM
L7diFoIMEB3p1DUjj46hn4DX3bCNOCmneo7OtJNGWdh5U9NpvfJqI0Hnk9Yn5xdo
JEq/pGkMJXqN42ZpbVkRgCLeGyUZQFy2TkOuqLsc36sqAjAdSWcFU0G9N+f4sbf3
/hZb+9ECOhN4fT1/MWFHWJZCJ9FVLSrqiwRe6RMg9bs2LtwmH1oiU7Ow19+DwWW/
RLQv3B9p3UTUkkhvRDEmEO5BS4QoKHTJw6ta2WR1mMjkZeiRuBy4DwVagDIvU2rL
QzYN9ZJWaeJTZqLxnbM0LBW/9xL4H6OyiOTjP38GqkOpzHWZhOSdPGSiJMya4XuH
rA0GswSA0Gm52v1Cq32k4NtKiv/AdOfcHfzJfT/3Lvm0a1IHR7emKge8FURvJ44r
dnEWgFntntINcAKcb+Jf8hTvwzbX1QNrf7j5RhLKFjBnQNfZvenzR+ggMISNYHGl
VZlFNzd8Ie/yeHNKaes0ltJoRn9I0Stjwy/aKqOpodbaudlkZWg9O73c2AifOh7x
vCoclwbE4CUVsQZ4cMdvmefYeD190sL8aeqNq4hd9qiNIc/TnmAMP3LKTb92Y/7H
rBVrY0H95NbUBTw6EbkykRWFQXQuf618+qx1GxZKMA4f0H9tm5f7vZ65+49McwJ8
dKd4Hl04esSZT1+bS7+YUtY0HRRqziIdDaOzHEinOPiXdVJvi6VktolkpHR5Chl6
TvBtKiX9r/i9RET44x2dKhLnBdlmnCvJWkF88WXR3nWx5EsysLd2P9ILgqBmDJ8w
8Gf7a+4b1ahf9kndVxwOOKd37hK1SZ6DZeP5dqnqxRSeIxzib5R6p4RYDQ8Td4ZF
Fl4nmb1eKDRHsVLp7UWJXF2xZAO8p701RqbwjuodSHxIIHVXmyyFeP9qw5xOPDlw
JmBzanIK58zDA8QcMQ9J1DpE2eygNi3hCHC8H0nT97NNr1j9VyFZRYgq4w7/cM42
08M3nN7H2n9ejYZBlp5BCJBeG+rjM64tQ91Ms8nT2lg58qMZTr9ZSJFAumZu21lF
3KG/BbnvT6Xq0Yhmpxh3JrKhwUi/PiCrTC4omkkCDKh06mvzMdA3spvPh2SvTejR
+4es1CmuVTia8911Z1Iqmj5U1Vh/2gMk0RICyWHvqqXR6F4kQVmN3TTTQRuQmRoy
kZHY/IGyhkw0QfVwbcXJ3Qfsqb5uD02b3Mb4DSZK5lNpIDsgOM57t7phbTqBpJJ6
THYRKNfIS8xDD73OsDiAA9NqSYsi0HVe+AQCc0QmqvgLa0+WS/FdVVmIdmQDXe9H
T05Sbb2ztByqdbFIMF/txWCOQxuxqOCgC6B/51HOqQE/qILdaHngITScXLHkDLYM
sLnOEdkjNPHi1z4uuP1F2RdH2dJRRZOXMXWVKSpeiRbK29ZIojakRyztpDCAgO1G
atFm0tHJGgQT1p44S0hts6hIyQWkUL4v11/gMw4r+33cce1Pdwa1igIgBP15nGh9
y8kr6UJ5ZmWmPeUeHHWIk8ul/ndM/O/GO7ZYrdKF7XUT4XjwzYArNZW/u+GbPJoV
wDgPe+qEAJr5FjablEW3D1e3sSGMPxml6YYhqAX28QpYVyZvct5LjA5YUEzhGVRn
KZXhgBzRhI/zHmzQ8G9uRR6r5pBfKJYMSihNrqsmOY5FVKECvhVQo5FGIRxcxRib
gMziagCA3XyobPz/U6Ok+RbesXg06cJo7BMxHqfRS0e5YTQbj2srC6ySRjU6sm/U
Q8cRhlxwv0uaOeAhXhv5FSPvzelNWQy2XawuTiKTXMkl5qX9afoe0BfT7El8F4Mw
TJAMhjnRNRO1unjQknBSS/Ujh4xGlCoOojv/MFtUnkKDnpbYMX8aaefQjXLBJgez
HJD2BK2QbCKgLzk5VRjvvBWlloGbehgrq2YsUhV9wWI=
`protect END_PROTECTED
