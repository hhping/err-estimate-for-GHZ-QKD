`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cSfRo9z0ckSZY97wKXy88dFz4M5fehEVY0U5AzjJjk7I8k4UlAVhmjg7mV/N3Jds
GG8f6fmuh5zEJHumbtdZ3Bz2tJay7ZOFb07PNMonc7NNqt7FnXngByzUY8HTGhcQ
y2xx5vViRuQNaxrK9yFVDbJyamXgRWn5aYUxJTmNepSHK0uHA4wkCsijZt90Z4YQ
LtLOFLt6n86nRJPXMHBNh3jkgaP6R3ym+4ix/p2zWvpcIvsi8aIdZ39n8FV9OiOH
ysHrQH/I0cBi1r9swegCML0+lHpvmtI0LlbL/0cCqj2by18a2YBYvU3iz7qw9xeg
z92DZ/nIIM9dwoS19FBmVKjQhe0FXIqOGdHa5ufiMHhhtLomhJjabog0iiHWdgm5
UgRUF5ZvDYkzjfGZin/OCQfuDI6z/LIbCmS6eT8u8ho/3HL/Tw+7u+iHXuObCieG
BkO3CQEsYmF5Q4ZncdwketiF6bShM3kfVKKnC4nB5q927Rg+ikm92i3QVH4vqfB6
wDUow9TPyaiXZbwzQCYS5ViIMeuDoZ7j0Gxc307vp1Ovid2c1vX+8c9AfLdcDB/V
xK1DYC5DESaT2qOHTfkCEQzr0DgZXTTEnLnkqjAmWU8R4wm6QNWvO1AboyGcHirr
ky9TXsH/+mz5F08gnTbbK/pHAtn4iR3y/goeOFKvhw8euUaf4tJzw6X3L8YmgROe
MYUQRY2tsAbyZa1jfGZNtOQPNr6gh8xIUa/r0bH2e3M/6UH9s/+5oHafvBUT2BK1
Vent0AVRqMZxpo8jR5MFuWtA4LPINLCe+q2qDLQY3G0WC8VMHgJvEObJXKHBhI8E
ztVZFaroCGS+08S1/Ep07dngYW1RVjhGobzr3HPaXOOAa1zBb5S327BHiXJ9OZXm
8WLHZUYOb2iuOLu9oiBYP1CnB4j2AiQhItb6skQifOMoJLNY8kpw77LZd3IK0Tj3
l5uJcnOE+6/iE9/VaPYAKw3BO8kwncSCmYMez8QrmqfbQfZVCluMuswWqgfBX2Kt
P79c/0EPy/ft2QxFfXcEOoKo9or4mQ/oVLNiQAZue8PFyplfp7nd0PZxvlEJHRid
/rdl75hGfrDWkv1s6O3y6A==
`protect END_PROTECTED
