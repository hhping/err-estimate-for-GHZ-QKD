`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bC+z/FTuFnhotothc8RzcopUz6YsyviE0lmO+7UG+nlaEO5eIXWsQnPoL59+Uvpk
3meZdQERHjVn/XzO4t/cHF3mtj1IFFENCGxbAQCNWjbZVeDTJEBw0hDDss8cEYhO
KfKI3oVwyLV2IiT0C0rEqXcEcI/WG8GMxb9/GzwafRM4fvo9EX1EcEHNbHrSMBU0
xJvl6tSodnUa/5S8kSGINGWs4PLO+nNSW2lbVEt0ythySe41MdhP77RtIAaUAOLx
TLa/NMD9XncyKhR/M1DastavSnWqgHHIoZjXijKP5+QvS3eRB68id3YZm2bIvSd8
myHqZ2pvq0wMaL50tOe7GoCWsrYUWkK1gYevB5/qifRcV//CsZmanAYEpkFzA0Ae
KrqH6R7MF+sLf0WShmaOvhDgFQW0I4/3dOaSY0KEIECehc85Y+SvWeDuKWtpDH6t
XmibETUtS2OLXJQwpNcyLqIwuDC7mEdlJdqNiS1Yfg7Wp2c+9i6VctjCmNBbFBL1
vbB5qDSJ/+UGPaHeLBNiNpWFcmUbmCayLnej7bcd5CuLkro8gF8b8G5Qm1kGR/7t
adUC0WCmaXJbL4HtG6N7mBK6RgK6s/JIZsawSlchtu9EXQRFZBBoD7o0u4Han84p
AA9cvSIyhTIupS7nv3HMzdr22dH97SzwnPX00Djs5sJRM8qA4hWsreRDDCKXPOIt
y/hFrfVm56vuctqezqcGSF60lYwEZzYpJx8aFjTj049CEWq+WeBu5yjd0mC6tVLQ
lLzyof/la+h250JHN5dAaXHNRHz3Sz2+d07HXdBq0hjczcfxXAj8o8lTv9sDjClD
716yF21PNxs7koW6pQfbhigl0UhLyGNdJZniGusTulXo8mCsPWRIFrKe58R095xb
bduPZ40FoBOR8QgLrQx1mc5P6WcBziFxIW7Z5geT5AGq033rnemzRBeBASi73kN4
6Pw1LE2xYjoduk/wwUVX5DNQsA+32KoUAGER6Ob/Qq8FdABs6H23CS5QzYqvzP3r
NLi00UHNfu2dNOvMJvh/1kRis+wpQILWzob/bgi+hTReDtEnHdziMC+jtSB/lMY/
S0kekwbGVod4HuLMMhaACLv2eIH8RHQPVGElqki1e52yE4fZ1fsi7p9D/Jz6inLE
84QetpJclXki/0gKPvGIGn3QkomnE5VvD9nIpWYGexltuVI9H5JkHm50Q1eQn3IL
sNjxgrsn+YwVJ0UIwDzSHM8ZTzxzFYh92gNDIf4U/vI=
`protect END_PROTECTED
