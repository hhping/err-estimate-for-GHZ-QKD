`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZHd3JyvtdC3UhENBzlAfxnZk9hN8tzfSpF3TvjROk2QnF9XU5GCHAh9Y0NfE/0Im
6tFbmcs57Vra0WHNcPMBAipGPMd0c38LpV1zXJdSNrMKZDXE7NGvOAVOj4I+vcyS
ut9ynvN9BUarBDk2PYfFm9cUMKUnFK5Bat+bRXJp6PrTL9mrBD+CrUIpeKANtu3L
Z7PFGGTzQrwjE93ItQhgjMVr7Y9z/+VEbDhEK9+qXLIIQqQKHjQIY8zSFj7tBkiQ
/T1y8lcWH5Q+Q4YEfNBgDeYEIO6kQC9AGuaJlRleO/7KF+Obcfg6QLAHn0t2Yc50
BSIl4nYvYPyLqsP1e/CE+6r4Vn/B31OPkd7byZNrBsf6VLUdi23DB5oMssduNdrm
UKvAqvbRS3dHsSSRS9RIF5eCsOK28Gpt7nONPBanMSuSGWhS07sr84zFbRDKTs7E
Nt7UnRjD4b3FxvMhUrHUeFxFHBxAf4HGchwx68xLgO5Ft58lDsnjGRwhuv/z4pWO
evI/1+IgLSVmJDaf7cJbiPEkqf6D21XhzPcQF97qSNZLJGi5ocaeD2xDsV738Jll
HhUHTz8RAtk6vK2xXoawbE3vExusejW1P1QfQaD4YaC/SZ8jryLHEXOAfen6ouh2
`protect END_PROTECTED
