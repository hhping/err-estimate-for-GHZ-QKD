`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
scvDn+UYRrm7ArjPQzcCTYCVJc8Cbu0ZRImro98uGbycNKSfJR6vdiSws2M9t1yZ
rvkEnkLZ/wrMSFNa5Y8ND0YwM071HeBGFHkhaKN7/Nlonhm8B0mqYnUV7SBS3rTJ
aCjVbea6P4RGsI6gBEXRAmJpjyox28h4gvzw2yqTXdMw7scjPAM1iKUx4KMks7WU
DO1Gpu6TR/cAIX7NrHSMQyWzEVQAJJyHTkVlRzqn1bGyUtxc9YRAdBQC875Thiki
/IlCMJsqvx0JIp7eE+bXGlaQ96l61kTg1Dkpm6JIyDxPTjJSuz7qk8gco6jPDCBq
FoMiC0xrPTDsYrkJhI4nDGUtCp28aT7mt3UyvR5r/n1b3+31GZY5VoN7UqeigE23
fwyD5Zf4WGpIUIEpMGWb1291KXA6ZZ/Q3w/gd5Ynre+RqxlwAh2AOUpv7d1z0SR+
xs9jgKijlnN2ectwAKpgBQAM+nvIDoz7X57YS/kumWv+QI95Gdu5n57FPVbFZ8G4
AtsrnDzdq4CbcgW/Q89ptTzKKPHa7dFBQdPsEwzxpNQB4O/0hpTFxSG3YZy0Cfpw
nEEHKrxvsrZ9lrprOFLOYArr4XIsAtJTuLOqOH7n55hSiDN3c5jrSfphVN836D4O
bJ8cvx64rdEZT3OXTlvkPwej3ZD1bMijzCrBHzFGD0aPUPp/Zjqh90JWA2uoOki2
UHmQtB2+RAViH2zK2SfbQwA2Bht5qzGr4iqvRGsTTH/GZB+MHXkGBU4q1od8BuTL
ZYvWoobOVWwIQRXIoOQ3qwsuJFcbEBM/tq72doUMnx/czkLBlkIy6tvMmGk5e2WW
VCzcEqoXMc3//LIOUzQtn9X6GyhOldocuTkcwSx2PfHQEbbncSoOofb++FwVzP7A
wIImvBou0CzD3Egn+KfCub/hTz/8bnyOI0NZQFqfMHcoAxJvdkKqbYJWmWLG98Dx
IuuKOnJWvthkoywL80A8OtTw7/DkMZzZlalLyPf4+lz0aMLD/JwcscoCUFMF7Yqr
3Z1pFztrGsCnOzyce6FGzmwRHzTp29uY08MM5woEwIwWm2bfvN3jkmLT4sd4s6QO
kZl9fRnnRm/pf/HIX8S6OLfB5HTcibOe/tkhbJ7s41bBrYgTjRJF+x8zu7fEapuU
zw1kV0lv/UtoiVlyccMvE5WaxFH3K2fqNkY03Jg6Phf5m54XXATTKRqvvbjwCDK4
tPcKYnT7trWW3xwgLu0cYRDccFOybgEDl11ERwA/OzJLpX0QCknu0RdEo4jolqTQ
MCA0ZunHAD2CswU/XXcTGLCoYGAmMQyTfh6cLMmgTvt1dWuoZ5/WaMpcUOhZCCaN
2OQGGWDcxRgExOu+wOsmbDybwSjRvYSZZiykGfnVvkaYzsAa+Bnwv5g7uDGP1upU
dgF/SZ70VyVeBEhSwK6vtDPnEnMgKYR9nIaLAX5qD83HEJg2J/aK6dmqXx350fwr
O1fR1Lbd1l1OjeRRl/NtkdF108Rgo/8rro0/0VRRgqHV/Mj9e4lgTHdWkKh5ftbl
qdoXBnRufEdbzOxaY/O06KkUpSYyPW2dIKWQ30R4TKA=
`protect END_PROTECTED
