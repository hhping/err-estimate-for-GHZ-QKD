`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fiG0ztRt0HyahYWO6sR4z2RZoxy3afnWvynCsuYoLuts4oZnhFD2pXPDQM3sCAaE
huq1M5HbE289rVy2X1Y+B1QdCBxbfV1isf7W8Q5evEzC/5DctndiRqT5y+zzQHAR
LvW4GMmJCIyYe5D2HqX5hWalX+rvk5hQOyBCX6+aU2TBFcZNmt9zzXQszAoYwL1G
rBgCNNR7om+bjPuBu1u9CpvGv52PeVq7rDWJBM9tH9jySF69T60YV+hDHHd/amW9
R9isMcLapBrfh2csOYAlY4yrIVEboMIOo7Po8ZfQD1q2dXcamsSuyfZ6GA8DinZY
NxDSSn9DR4oNi66QVGQUXMMmq7nOOyf+33fYu/JSaSBLq0cBHT4L6JM1oaVBSSGC
4u2CD8HhVTkI1hwveI5PiAIofs88mN8FI32mZtguvddgbbeBqeHuaVNteo9TgBSv
vyjjTf5AffoBzkS5Xi40t2ITvn/DHo5mRoOPZkuRfGxucUt6mN1nHw53PEk+8Xi2
lRjqPSVwm2O6z3nBmLsIuC759fNrhp+m8eawf/wNsySRmyicxhmDT8faujMOwlT3
/UVbjQ/+Dp7T0lr9N34gYv+KUPtNlCGqOytfZeqSjS/v7jODPfqbf3ih7G5V8kiN
WYRUjkmYkU/xyW6kHfjk3Nt6Z0VlKv8xTx+69aDXywI+kpsgf8E5HJIR1XXekr9A
XKR9hkw6iw9sv3LRIbF95+hStcKsUjiX1u6lmC9htUYTap7Uz3NZQL0nD/rAb0GN
+/2HZdRT6XnxuQXNjLNt1xRau+H6uadgGzlbWtcVsWZUx5/K206FiR3u7yas0Zr/
2zTPRucJPJg7VmI0QWr8WKj7Rk/aA3bZxeAy2iOteqs2DKlEVM/7+1Ko+Obi3GYH
l+ujHeXIlv/nMZmeyNAN8iquo25ar3l4owjLmwY5vVI5rqfBfUnL/nmOZDvwt0Rg
PtfcE3mW4OgxaO2bAgNMcq5QfqVElNa0gTKcFwCggpTq7JgihoXi0zNL+osdvmZ9
scJ2dqoOs43qQ9pAVDiyUoKQ9iWy7Lol0BJDoDQxedwwPhcv0qcV04ekSP82El3Z
eMDMNxXYIupMz4AJ6Ww3fpS9eHH+ChsD/erEo8h4FFivtn0u/JKCxD9c95sdhNl2
5HyoHMTlVvESEdOBkXm00teh4bcrJmO3J+4PYeVVyVYkM/eoKdnPhqpxGi+M0oWP
vtTtr44BigrjSxjmYtOnKsK3cEEz3jYNgoQk3jvnQlDV1GzwSYcxGsEwtCN+yKF9
XnJXfbxYKMlkrkudnT/1TgQWSOtZBC4R3d1uEXrc8+7n30QPyGWTwQyBPKlYTgio
FWG1oGWFBNBfEMyeR/zUin4kYfHEziHtMM9/kXzEK6xxNo3MdOF3Pt6GxtqO2iWT
7ONJSCYRMChY1wZuoJoZoynF9l/ZBDgqeZSmKzhZcKU=
`protect END_PROTECTED
