`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H9VESAvksxcP9DzwcKZD2PpCcKgZKh48ay+s1Q2d3BPui9RfaKffDPakLFCo+KTm
e6wWmcvjAMOrSdmIDC30BFpCzKlVfzllpOiTvgYdSSod8BCKMOPeS21N0x7Nl8Lf
MApuQcI60mzD56XJuoIFowdAA2lyKWzKuqyKTFWzY0LTu3zjfWvvOrHfD6EpCQja
xOY4Loe/WIjxz4oseWgq9K9TG13MA1gWfwk1ts3GTrwIrCpwxhKp9PK+Qkm26M4I
zqeH5+yJDp9vXAYxCXlBucgn5ZXY3bCYyro88PkO6KVz6ve3y6se4W2Y15lYydSl
gkA4EZEtu8vNAZ4ctygGLcQ7NYbQ6TbJ4V9lO4iD/oNsDjIheBNDnzeiPv8sJk7R
LW/PJ8lAuOWToamEgpOaKvhphfaUVI2WZeyMAIaPg0GPMzhv0sK57G+kpqfatkkh
QQUnxMw1/c1xFCo2ZOmZCyY0fvXe+9yWLWS9oXQdi28g+sunQcqBG0no+vKOqXAl
7llaO52qI343bOvv5ScrwYreUHpgH61upQDOSIAGxFFMLap6dR+4EHv2npIPgA1G
FXSmHGDPlZQ/HRoH0xKJqQDqmLaamSc390YrA/LxaorDf3flQ+xiFVMnD5daWtF0
vVigIeVIv3NWierpHRhiVuvWh9Bsx8/LIkRLC13pnINsNCEC6nFR7CH5UpCL8iWf
aJc6LcPxBNjggA5rasYnhVK8Pp/ywcBz/8PtR2HydbynufstsWE+reVvVoH6+HVt
sm2nPWTYjIWk+FB2Gw1K+MbNaVDtBqmNnu9lVMA3nPIkG9hh66x5jwfnpQq7ZdxI
4z24HRRws61jcDsaHOfym5Qw/za27Fskt97HxkdKhJiLwHzBQtempLBEFLC67HdR
ReOGrDLJ3YC0/bJV5hIZ7np8Qvzk6fXlP3LQJCDaOyEoqgDxw9armTStx9Fy9goo
8iU3mGWZddXNa722H+Hk+yJSLjIa+M+eos+dPRLtfa5xZXhpD9zbq5t85Uv36b4a
AcRunKViruCsRoMHBlbEEwrIqtYqurBXa8G4wlg/138ztBtFJuBtpXEB/Jg7jXba
Kid0hQB3wH+3wKJdsybDUKqeepzHnkezFe4TV/gE4A1Yq0H3qLSxeoHs+IeHTNI6
U2QX2oop/apzgd7Uj8hFs+imdHH9ztDqHTEjDIvpBoKPOCRcL2nHX6Q0tuDTYFsT
vE/m0aKjTmxv+L/22f7FP7twVVtySqdGbtJkmsy5BtA=
`protect END_PROTECTED
