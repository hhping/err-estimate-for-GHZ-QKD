`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f/VrFD+Tu+2Q3U48msrJOwKBnGQcNp4GCA9ilklt7btv7OeiilCwc563XT3fvVP5
KZcdg8tOGYWgKhyqKkDA5/nocKNe0rNNzIXPE4k6MjjQjb+QDcKZApdYsUeVGdBm
tZpiAXn/ybYKzPxfgoNvkw2HaFOBd/F/qMpxkZKbvM1+9fykum/pMpFq++z/vhGI
p+9Clzzok1ucgZhxO1672vY7uqHGovttUsZzrKV7I/CYJVNIQQrm7IHJOgIAqmcm
UJzsVqQ4W1Rq3UXYJGWQGduiXRe/PDzA0KiKNU/DdYNRX/eViDR0kslrFXy+Po2n
N46YtkwpWLcun8mfpu3S0S4O+DlH/HdMFmHQzi4Lu/Eif/G6F86LbUSSZBJKh3jZ
YbVjyeGhag2ifb0+PRp44Vp/hYg7aBOPcPedHlr1RKSQOCwmDEx0rn9utkuLHNdP
TqiC2z/qxOlxKSxYiHgKqDkm/xpz78ibQDFhiT8GZkEYMChIgJjUUJQ2Voolxs9h
uXkqdjlLQfPkn1TkhJWozwWk4B8mRZlnZzmFzKXpaKx+KHavJ80Z2ngeE9OPyKQe
hLiEEjZv4bIgg+mGVk/uNa8QcG+8XVAGABHM4120C4Q=
`protect END_PROTECTED
