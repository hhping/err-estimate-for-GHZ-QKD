`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b3J3DGzKajqgrwqNJ44FSZ91hso1F/UvGDrc85qmC+WiaLh1EcVB6homa5IkC7U9
fVJj36J9YK0xdNzJDf/lu/0u+etQYb7pMLJL4GqkVE0x1HToCSzsbcG4qHxgDxUX
K+S5cbQVDBL00BbVlFE5fjOYx/Bre8oDBY4hd/NF1O1gVh0TgWsFGbBqlyZfG8BB
L33LD2oEhI7s8s8XYzYM3vN30jr7HMgoKRob1cdmJxIyb9ws01B+gcpOS3uoHwYl
turo6GCLpZB/dCZKhB0YzdYI9JrAkqlwr8f3GmeMuQ4iXyOOZaBU77pSm2XXFk20
IqBMw8+p6XZrPh0lzTTl0Sc3ftvzhdu6OvswEATngfxbOkFKXu1UnGksx7vHqd02
ojl/e4q0jnALc0Yuexj0iY5f0l9PzfzonOc3oiH87Jt9/GfYVQqrP3k+Fr0zwr3s
Bdb4bA1MTeA9bXlA+d0AfgAFVxktii2bldr1YjQc9H0wngdmAN47kz8jWTgleqg4
Z9zcqdZAb4S9Ll1AaRzhk8pSL5Hln5S4rp877WrR2rDvaSFvgQe7lktjbEn23pow
xJzV5GgtixtnKROTAWLro7k3+lY+nb7o0KB2c7o5YSgCp8FCMUMab7OtmoqKzRbq
rt9kdLDBIey94DvCoRGDiHQLwzdLPZiYgmK3v79mmIyothxEXkDU0D0/PKTK+x3p
eAh3eF3LxY8aKH71qNd7w/65CpaHpQdBwYdG/GeuNmK3jo2S65Qhe2ZyUsnH2N8r
9nLMGzml+516G/f/0pobDMiLHOYWWQ/uhTXXlA6g4tlRy8jEHdVHqkhSUAgsybxa
pitEzEzfGc+faaG4XdjE0COfxIV2gKCIiRh+9P1uhWmeg8lQP4LXxT4cGbVOG01f
gT6kgsjOuvVXnY4AGrDD9kTdGdJSLn0qtP0nNObxTZLw119zxPlJSRV8qATqYqI6
vEvy5t8W1F2AhRFBP7f0WihPniQpN+eQ0/wAL+PKx3LKkvZfI2XWDe+cn6bxDoxK
9/QII7PF4Dw4epNhmfhWQonZIXXVWVx9jKk8FJmKpyeuLejzeY0+BhJw6Ok/WIEa
bSBgf1tEn+Zq1danouSNsSY3KXy/Cz72hAlLOhwvMqxx0Ew2SblwJmPxzLcIg8ZB
Uu3rYHuTtO4FhHt/vnhyxmK0idaYhuxD38www7yjAonjnCIln7pyQgHvm56BgCXp
gdjWicqMQCVL2YWDhR8izXpvPg3lg6SUpvLSr7kZj5zrGZND1TnMxbEyJydOLAfM
vH/PP3rYxRvhPAVCgZBhr8T7V71wJSE1b1n+BtBniw8eijOtbHGOtrhKCd/EeHQj
Ofh6nWnIB3j55Rxdhw8tqO6RX98Ny6JvGQSB3r/aQaB5ZUYJFup0raTGG1MGVts8
CD0jnF3u3Qv+JRUgaj68K/e8E8P0cAwtxpSWVsIFhPGTQxrkQ1MLz5+5Lo2CSYOq
ziF2niX9uLKZRyw5z76YAzBP3EiybET2UbV34fsl5P0MqMMwahho0j73JFAnV+Nn
NXkePmMgFNw9RqCkLMeGLY+PoHlPgNlWYAIyTt9ciOHHiuFTDC5FNoEiGWt7NnN8
AW5hLx0s23sPP6GjbzkaH5fpxmoEDQ53r4QZ7cCXa40fqNCEtdwLe+MKfMjzMscj
RsEmvyfH70OrBSJj+cZk95ePAuOaQbStIjCBidr++UksTddDiHdo/BSDJPOOTDux
3wpUY82QWpvNTm7/jZgb0+lzdmFTCZ3UfFkXB/4dRRyGDUwu61qXBQsE6hc287Y8
EVWbR42izBjAlqM9Ia9VFd3Frvt9vshyjMtZ4IyyDx/+BgBXzLoruARhsOuxVtBb
T7t0n0tJiw87KF4sTadMD+0AGkErJ6FQtZXlATX7KGJGfVoh02b2gZfC8T7LQKgW
1o0m2MmjAKJ0H5jYua4PmuJaPfXBpEeD6Z3dLK2x6YI6QP6UZa0qrFaxSWGrXjKw
j8qB0wXCPVVttfz7ONVyj9X3hKdGLAX9zpcCZa3b8gPW+y/KMSK21XfHxx2IfD8p
x8LH5d+sBiaJ309Z51Y13B59lmxiGyMqLfjwiDhxyWIMYYET90XQThYwJCBL8gNO
nCEWMkI0hxwjXHR68/xLxQQvEVnLhtq9iMyBSlDC3TGTrVKr/MdLnGf/gPEobLdM
0Qa/rVcgySCrpwhj3bjgmsLVnKZxsvZIXvZj2/rWdo72MwF8HKTd/YrTAqLg0hbR
vfdmP/Z+VjGeZ14QnwbWCJ/VLbqeAlZexn1nGC/n5MJ0FwRIo1dCzq9U51O3+5Xd
mpyYZRSVlbhfbxphHqChb6RpvliRBsttcOUejxyRq8ZLIoKVP0Q2naPnws4mpP+z
nz5LUwBaaxtzuzpN4hA0rvYB4VyF/bFLasBpM0TJC4Niw8Gcv/+RyNFEHMbCkCTW
G4XBUdTJQHRH2KOj265QbPqN4GNr4Kw/UaD5lQSCz6EewDKNXfC/EefNaPY1uRz2
EGKxEKM6mpQAIqzzDyawCA==
`protect END_PROTECTED
