`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j//IZbS2XS3CaEz8sF/TkVdQ152XKfsHPb8PnrvClAe3GaW4cqNe9HOpxSyhKRri
TfuzrHl0bN2ulZgtoty4xhOKqXTqBIw2PbsnwhOVZ3JfRCJGfk5XigYQl9l1PvBg
YuwkoS4JAHNTKxKgU9PZimXJwKpBKDWfQly9njA7AIRDH73+AraAU6+Oh2+3insd
iOk7j64g8yhnhL+uteNv0KKGR2yuNQkEE9p9sMnz4j//q/jPNVE2leVLFaoHAIeb
pooUS8l0uageJsIukjAsu1NXKTdmCmumzwRXaAfnvvbroio2SN+rmYyNNpIRIzHr
rXIO+tYcnvWfU/QOmmVUYDZy0b/GM+dRO3zgGoj4D2cBTPQhOkkdGCpSfuCoY67Z
x/HW6xP1FwexSHRqgmltz4divPKFwgOrCi/poeD+rijx4l1gh7jhMIp16TuGAeVl
anMQ12AMWM61e8YPGe5iurB0UbdQp3HQgfo6Ma2PhyMYaSl08HsZ5e3Bzdj0gj2b
itWXYWrxQ9voKHMrurEsR6RTCDlnIFbGzwj1i6mflyeuL3uL8qwrH2I9avyHIqUs
kPLYcu2dLwIE3t5mv+OLGYwB1TP4bJ7BqWlEogc9VZSmpD5ThTeCNptfMXXtTwtf
uY3RyIDmV5fD/VxjCAtSjqOWlB1pZNB4IvN47BbNOavR6VdmHuAaNidCn2tFXX9j
6qMhWRiWomw9F4VQNXDNXuXmVpKssGH8L/ZoSuUqb9yCxfA5t0G0X86/XHkh1Dcx
WFahQq23fRgT958ngZ7vYleZX38ZJBKhr83N7Gmu6RbBUcWeKhSJHE6nw7QIqK03
rRtPmSmiBkXbkDtE0VNkJIC72rNxK5vNgAev5d6TyiL1iEDbGZbLTDLLf3Z4Jn6S
LvV7TtQoUJB7s+hb/OrIIId2RAZ/CKkLq7Tjh1IIRbcALIqQj3a+uxH8p6NFGthj
0PDdcEwKmhtJHOrmTfWkflz+7228kVxLuAKrHxtBZbvsQ6AkdecylWlEpWMEM6do
wsbKXkkPCUh2P7KzIlL5uirnReWSCWyObT+Dl6A0m5oYfJS4b+iOjOjn4VLuKxXF
iiGX812CVAcjF3t/8fvrvbWi4r0BMY0zqrNgbHhwRD8h7VN12JVs1Y0Y4PsuaMBV
FI2I4T7nfJ6bhdFYoosv3DxlHF8K4M8XXyB8ykENXhy74NN++Pr1YUwSjdq4J+7g
jnEoOTE4veBPiGwVobykvkBoLXfPBvMzmtDvGsyFN6tfynF5Nm2gKuHHMEVzbww1
aZ91ZE/LJdJwUgjAMiJhb2LSJGog/33k9gyeq173rRs59xljH7e3B5hVFUlnReE3
pbxRsQIh5J3pOINoAGQMgA3zPBJra8yIRYGq0zYbfu5Ctk5t/zGZWWuPbWl9fQ0B
hBxYApGfjCC9eZ+UxUR3ncqxO/bKMfn5bHbXg4IjCigAVcSc5O/jfXyTQp1MVnt1
5SLlu7Ku8yE3ivugbIRJuWT2+dNLWG4zCfnQgV02NehoNMM7QzIPBR2mqefAxksn
X7imvAVGqFiH/adQmXHSaL+o/zAl3E0GYpX6q7kbH8sXBbpF89wba6gSzsoJQsWm
qgijrHAchcWQtmlmJ7dbA4RfZ6zV3lqN90Ojdh9Z5NLr5tlu+FCqiVuus2AG8G2U
Xkj8Xc5GEx2IojSH8Y/rbyKUiGUSxk5mr9NVCXJ+oxg4LT76j3uayIrEqjIXn0zM
gCHlyrt7OSlrwrP1h+gz8eV3Iu49i+bpfTtn+wG3kfeMmZZqkt3lDuZs6RiDTzbl
AiS1d0nnlaKsk38DVUMcZaqLkbvhDapRzl61FUoCtYxvGPw9FoXZZj8zQiXSQdfr
bEibUYhIG85DdQPA5INKSO8e+Ju+0rTSj6FvBC/ImhPwhdY3ZN9c0+YBEyqcG1u3
vpP5KfKOTZuPd2h9ubsz2+GfcolLiQKHKC7mnqJnlV4paRD2uw+0m1Rk/qNuycYf
`protect END_PROTECTED
