`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jgmhrn9OXnqIkphX6edZ7b73p3wkziHvChR8nTDjyHV5glWAuU1/AwE5sxsPcbhj
KfEFK+lo29UOAo35LTAyuyj9tV7lvCo2cdbt0i0PvmPgCTIKPy8j+rY/Va+LlAow
2xli2uZFOmgebhEyXeWVvxZ6JJgoGDshJkhFCLuAPfgH6n+g16LcXBQzUdHf/Wqy
k7V1BqpiPU14T3ha7SSXy4P4WOU1ni3Mnh7o3zfUa5i+VaihSJBCoUT3CYwIT4ti
d2P6JEBYcMQBdbKIMZvv0ImyK5O3uC4VNSscBzKOepQOUp9aNe8hVH1gHrmjdhgz
OSPN762DaOtsqvve1kK83Lq8oDeVheLypsmvq9GeNuArhuAQ9mlVVrv3/fhHbY6K
lBvOVYBeM8Wpxxf9IrfW27DHZxI/3V9+N2E3rlZ8pPs6KSlz+v4aZC0qEL59X51w
xKoywuHq/ACSpN5mzkXcZZvp1dqSgkvJxZyQ5gradEM5JH46ttJJsoocDC73ztyL
XVMis0IOczCVG7k5cM7ymKqtMrPlKwRcE9+pDvnV2QOmggQJvEdfJTsicJbIcFR0
P7geUaeJG7YgyXfDUXV2prTU4/gJeBs8Pp8ulA0ZnjMjmHIx4908uPTHBSob4VfL
0IZ1t1jKb8ovkbw1WK/vqzYdk+3S602n5pAlBhDiVqNGPEBP/XqzZBwJahgeLRpr
CtSyxpYJXmjMXUtQlMxYPpSZS/2eOZsULAVhzK//+6uR4pjgWPmDyOVomjQaXffG
14uT5AFiTVZGr4crPHA/Q58Tg3Xi79Z+3reMdCs2CfHQ0/mIr/cQJnONCUUwi2K+
ugsgFRvZREmp3qXL+MncSqO0Yon2M9hCmI7G2lUH+/qEsi7eXC+WaeMD18DZMXlr
lO0+CN5sm47Ef2FOhp6613YmU/jza3JmzYS/uH2hNB1zrvPaQ9y6hbAFaQG/QqeE
xDQe1JLfLqEum04lhFZfedPkX8yqmeIYVHr6BCl3NMHdXw6UG72S6y9UBUjRhLt5
Qdwix7hZpY1wD1WJwzmjOOStQIiuzZzyc0uieAhOop8kKZbIWtKAJxslrIHYyNBh
v8xnYzsB41tVS/lKDEMiSdnbrLEnG3FmFxUFx27KCoINwDcDdYW4nO5p/ZDGqfs6
tXrXHG5yzYjaxrXMBoI/JTbm0l/7MHHMqopkO18tW09f4r/SHdcF8w5gCk++YQ0h
BzL7xvcjbw5vp1sD8weEr5OHqNDU4RSRrP1zmuPJ4XNOmxGK6YTB61wOqCzmSBwa
YUh5e2fSWn6MALOG6gOnQhILze7JOCW0lUzQZf88YNX8rxARIt18f87Od0tV/U4e
4knq8teVO4xR23Wyt8TlRALnUS6nf9WT1PAoKuO2kEAe4kxvBKWBkK241tOlUuGt
wonGA9L185vNwGL5UHmF88ny5FJbMdhxPxRyPmwuCAra7C4bDpJ7NqZCijKgDmIu
bfrbt6LOUSUvjDHvujubE333M8eIaxIr51Zu4jdCiTVREvVS1CUpyuAKMZBXX2u6
wWbFYDQZLPNoJ4Tu0Ncn27u6sXrjU+EDW5MPPPuIQgtR5Il3aXks3Pedit1s5OEI
9IkFO+cHRKjZthQ/JHmhZXsUd4weo6rdk5R32wbCCdvjENjmw/y4zVYyrRWGmiYq
ozJiQXKnYJgQhdtcUPnY92rpuY3lquzCJe+AfwfR5aXGEHYjeQkkE7u6H2elFpBF
LM1omOvnKXB3jPCFzc6FhqQ2FFJUPaALHho3wxRh9NhRGvnS/bb7YCwHFsGRxfr5
ZgI45FEYbxNWGxPShmdiFDoOpGYT/3og2QcA6yMbjcPvTuD7OGrpmF2wpYG3Y5ty
zvcyowThilPSXB39WNiZsFqKiN+f2XgpZeztf4G0PIJpbmL0kNdOzf+f/RRjrRTf
Y4ozvJ8yKPbutd3raRy0G0JPNFBp5uqM4vWUQzmH9WWCFFLp9ku4z87HkJu2HCh5
PYcGiVwnxc/zbQDuR8WVGWapL7JMeqjcNJwbw8Awrz2Aue7lfCVGnO927e8ZQH3X
XcMYqeE9Q8wUGycNahFe3MZEYj7+i6D4ROCYAbUueYCEzeAzMzhS9MVo9CUJUOtc
GrdiXdOsebWQjtItbTkBxe3FXpDIJJ8ytGW8+t/n311JhCHpYb7f7fDr4VSlZwKh
zqZb6vyecSWf2/j+KoMtaVHcb3nmo2XZ9t42t8OKOs0vZeCcYrLecb+z+1fzx8HI
9FPrpfpC9J+ybR0oCHTCzZG9X35rFQEwLMOxLpdRriUkTXu8NDMKffR/blBIf5uu
Dobf7fRKMtUv2S1NBoUEcDIuv7pD+37B0cFSEmNAJsMfoMVMFJlmn0cSD9aB9Tx2
Mkw+iFbq8gSP3ir7AEZ01L3i/LFCT92lk1XEOJoHbpFjJ5iV+3Iy4RLk76Ou3Kcy
QjZkznEeCwn0nphBlt03XRvh35583mrdxuORuSk72+nhdUt5lJyGh3EYnWXOXHYq
kcyXOygyt36Fjkfs8SDXzLxQ3AgIAL61EnpqMYHS/76HzPAWwh1PIG13LIsPjoYM
IgH47IUWMrYZ/k6glxHxaGYRjv/EANU1b1jLO5AeoDgf7prGyop+G+IZPmeS++/j
KfVkE65S5pM+k0exr3vTOzUf5ZQCEBGzrVicEnRHdfXk51l48UbYMEo0AmR1wZDd
Dch2Euk40SYWHCAq+al2ioI8vFtey8ed3fKYt5cB2/+ELd/BBe0bVd5ebg8L7z/T
vBYDiOywvqazEnvHdzkyrgHaP0e24Zkgnq4oqqajE/opeK6Y+4vZ+qEPpZyGuh2+
GpEGmhCoCH2GpN7WwcpgIVp7FFm2OddZz80j1D3gb8uj80gt1ztCr4IDJIvhHcbb
Mb3n8YPPkMvSHe1xhoHznn8YeU26gPlEy58kn+OWajEpsyxNO0aenOJ5Ki1L9i3a
qstp68EbZJwJqnXRHsB8zIOn5CzUElp47ae2j7m5I2gdf13VEKEekvXusydXoZ0q
axMcQh/qrxpbXuB652nHoNpVR6KflelgtOo6O0pa8hxV0P81/ujTKq6/F2x5Q+6d
KEHRwsGVXnYy2w+hjXJDZz+Ky5WwxC4vH7p+ENcl4K7KvFMjg/FIzlx+SBnEAgrU
HyzOdk9hEwzKO6vz0YLY2vY3CrvkVNLlPN1Wk3otSuWqJ+RYfoyQxeHTkTCTfk/L
gcDBbmw8Z9NrOBkcImntnh8e0atf7BY4CUH5CuXPzaVr4RxY19Myr1Yg0hxY66Wr
9nCIxu8dIVVRL18WLVfhojt6+k2zRRk94oX6NSY89l1G82S+3rYWj5vvKqA39dn+
IipBTupSNNHHQfaf2KFK2MEVDCQsLseJRSzNkD/cKvirY5EdLKZbxqnPgNVcRkqZ
1Tu+PA2FtE96MGQ7TBj6bUHka/ux8nXQieE1ur0WUawCEIBJVSymKaX2vKUMbTM9
OIdWRTrGXD7HpyBE9Ys/StYwsoX9p7Hh7M4LSjbLMyzXYP6Kz0UiFprigXnGxZol
hdcJ34qLwz7k237GKQbIbUOVr6SkSQNtFaCv9dg1JrMUsz0RVlrJenuw1ZDtWXMn
c9peLghlWpda9n/IWDV+Cm0EbZSklrjwWDx1FOs2GLCdBcbvi4fd3B/53KeKXfpR
kxGt3CTTiw8shcqd+oeKSyNA7QZ3Hc6juwtIxAR/A7NZgST56KwVKStqzuQd+fQT
SbsMjXVHedu45fpbc70VYFKHPCIJOzxFrtnyf+9AjJ6zupzH0V7gJ53svYmc+IPS
pvaQqimIyLehMvTZbuof/CLJFaQ0xvt9k4NADl6xRXuYJxZR8OG9VgdXYbT+0lKg
UjMa+dwlJsKOHoDRS9nL+KNw9aFqCmE7HoddtbK8+3SB/NjUgy2fwclkiFH9enfX
lxxoCcAN7DgeNiUvzVwPw8B9qni8l7OdAAe6UkBj0lhdazXFh0FEiYgs0PyglI6G
XNiFW0cZTLamZ3pezt89cu096hy8ylPjRN6O4MZoLnWuVqhBFsY/+WKih6cyI8dU
MOKV+sJSMOgRh5w0eO3xOrNf5ON+sAc9RJcd5AAa5PeiWDjFq/zJC8J59uM9n1Po
pCKqk2pY04nzN5xSeIW5VqwgParqFFfUtScNS+0C9KKAGJv9YUg67mDdXQou5tSp
ixFF+RlZ41kl4iqdtXwCKHXAY5RLIDVKuUQg/a6nD5zu5UfQl5jAZ82N/NJNP/Md
3iudZIqSSdv3AazF1SiK1YEmxamX+wyE0sCNS5yPwwOqurGiLUejaJhmbrtSUpHV
7O8oYfDRaSfErgyjo0rmyNpAZgDkFPsgJTpRISv5SsF4Cfhx0+ZPdCS5fZHqABKL
6vqZt9J2DDJnGrogzyTA66JqPeFR9y+o67rrEy04EHtN8vdDcRo341j9JZiQj7vD
9VsFrtJkJWaZXVkPKlcWUz9inVREAeCIxpfjn6XcOqO3ndpp0gaAmtXOzo5b/0aN
3/dxpRSCNcy4lbAAm+0XPqX+RDzfF9Ehkf+BCJTqzFEVsaU1YZ5+41ooOqx1uQ7g
92jcXAu49NZ8+VOHlpeY0sdrVzy+E/p0hlbZeOt/IZmEi90hlnEB7W0VudQ5g4X7
/XDRd8X55GaQD18AEbO3/UJpitGJf7oNFzljwmCX14LDhAYbSoEfP2xXmICoTTy0
HiKgNw7aroIpp2aUktHQuFSFExrYJJbtkqqHwri0PkzEM837IdaiIfi1R+itEfWp
NAWhqNEZgmfTdDkamCsoWiVrkI2JY8PDNzGdDEKoBb7WIIGolHzofTpCa6cF8Za9
Hxv8ryI6Nkf1Sq5uLo1QofKMrnpes/sUT73PbVJ2vx45NaoRkOGDz+Z0R06hdvaI
YdmMhM04hxCD+Oo0Up7TSTkW6dNq2bgXnkyGIDwy0JdnidpYvbvP35qGpxaKEjya
qE2Yzi291kQm2E/HdgHlfG7CyzcMzvrxyPM/zvDaJu0ifjN8uNYUHgdYSHP4atRb
50Jljtv/BrPMM8J+SIl8kHXHh087AhW3Z1xzk4Xu3o0XV5qyX0Mpwsu3yIqdVi6Q
wEK8DcfBC1SMaCMn1E4y96FfSNhQ866ClHCAmd44/VmvUb2FNJHZZzPkLwWA6OyT
lDR6IAyFIALSvePRYH83jqdtWC68OJqf6FNkSRk/zaHwPPjS7U93yG4EcdSKJOsf
pjegmKCQTFRtIPGb1sD7f1uuhaLovqCUYoVZXQTEZUoymm2Vsk9ZHNfj99iAyPEg
f0HyWWgD/XvslWIV8kJb5stWd00hd/XoijvWu0t+nMa7v2WdmTvGOK5XYMkD8u5d
V3PhhRIm3FwTXBlabtKbm1jUXC4m3FuWVygDfnVXSHm+5nm0VsMq9w0KEBSjzjz1
JgIZA1NqmH//WEgGQZhonZ6G82h3YS4BUnAAKuuKUSV4rmHVIllAA+lzCgyJ0u9s
ZHsDFSjym4MtxWeblN6TXK35+UQm1yJuPLPIofYN88w/4OigLUgitVUpiiZTz4uH
fpmElfjpiBiLxfq72q0zIrzZufKtIe6sxFEgDwt6WinZ6aTI6rCRkWMehRsasxzf
gv3lAiqnji2ePTcKIjyETBm3Lj24dZWdVEe+SOmPdJtFIhfVH6yJ8KsmKqMNQK4H
z8TKgw2UeWadwZaAWX4PGWT8OEWd4Hanq3Wa1VLS2OA7ybRI6iFNogkMbidyv6kv
yo7oNlw20Udfd6F6EzpV83eUcp/MfaK+wB7/Q+2xQyD5soj+b7jKCKyVkofrYUiM
b20jkeQ/vi6mN6i8sEZ+fmYjBO1AtQ18ZrFzI/eaRlA1UJjntCoF4Kkm/gwcnBGM
ybikAWzb88qF8XeV8JAmkntuqZcbsYNlTgELkX+/vOGORUjTTHnJI5CB5MfE51gQ
X2lpKiz94MzB711pKW/uVIPEIoqFNVnjzOE/EjVKiGpG6W1a0iMGX+tSKeWVdMrO
dQc0p5V7xC01XMIlQHum9Nk5tui2QvqsgSrrcef4kjWG0RlX9z6ZoSzrIv+Fe5sU
68AWBbb0rHnwbtmQMJKfHUh2UBcKPvVtgRT7QE6g3OHxIv6CC1tu0giDXllTus/e
agggGG+1SdIpmf2c3rmaY6kZsdjj2m02tZZHln/SniL2eSwNEs/GzA5s58rv48/p
6nH0VExNeRGu+6R2U4u/aLe52Gxu+59Rvu2F2K9c0IQss0/SkOxSqXvV6OoIoiyd
QZy0JSmiQxZRaWDmfaJJucSosaGTdRduJm9iEZ9rxYRZUqovbCLmCdUDD04Pcahr
mCNrK04aocM4cXZw6tjJ2xMniSrn8RVltnqA1PLtSoj9uaU8FeiFXITLWmcxER7f
KsJqCi+fD5wYKJNgK3j9ZFAvc7OrrfIIuNfIjwRy/S63BqMcZ5wokU8dH4om7wQc
NdFYfnGGNNDib1/DwK8SMpKA4Z0DVHzMnmo+u6hqZRWDPMwFi4j/zHAYSKSGX8aE
/kY/9P1cuisqNsihqmEQI9qdvkPrKgOne74Y8gvVseWEP1DNqsp+FqVYsMR3QWKr
0hNrPrFvP9n3Hoa5aJYI5LwHTmj6WgaM9vm4rfamz/76WhwsFM/V31m5jtICQKkq
WPFXN/gmuzkSNPY/fjUYHqVBK2cpjb0hWZfkKrye3JE8bewK3tMoBWXXAoxEoHCH
P9qYX9PLi9ZMVvXmnCt6rYr8AxkNAq6GXxUASsEJnSQtSDFMHb3Itq44HDVwmjBM
1iRpNyx3EpFEnFUk6Osn2+pZeE2ru+S4mwdvxsEaToIUn9MB0kZNVVYwv4+Ap5vg
WeUrA4b8ZTADC2XWtml05dsJLI7SvjW2Y6cccUzG9wOp6+XJKgqWv/uVeV35sHXD
QoLeuVUp4SG4anQGx25+SeC5mQSYAIG/QKmZztPfT95Bon/DhTXga6oCfUUVl43a
C0+OnrcbEePWg96synprghbTFpxeRgaOQK9/Ln0wm9UNMmxHXP1eA4PtRMVus66i
wbofPVbp9FbK0UMbEvSCtOIv5799qLeWhEYu0VqNpqHWO8TmOAB92lhC8zggVOag
/6UaigWPYhHSKtv1mNz42+/pQI3PdzJaReLkgA4x+R95DgE4GUGUvO+OaZ6dtg0X
GIZ63l7fd2YhTFGgzW121CgL56nOVNvdSCiiNtXnppnTkMxQuHLtfN7fNbpx751W
92Zi4nY+z6K5Ie+TkqPwPmwOoTTPbouOzM1Em9Ns2Rk9EvcE0Qp6HHmsV1V8LFsk
YQcVe1Kb5UBEoid8Kc/cyrUnMAMijtVpUb8KF6lnJt1Bv9J4pQiuvmSpGwVuiqBZ
0GEk3/c3TPZq+Mx267z/6sjZTuDR9VmnLDFbm262EZ3OMWGito+iJPujBsU+GgbK
qPyLwNd2Tic6+JUjJOje41Ws/LpdNfnrHfR1L3obsrSWC/pRPbL4Sa0UVK8YJpvo
hhzpx+6RL4RLrV1OPnOupB/37GAgVLZuspL+aWKEGINklUQdW9vALfFjZVXCBCoR
dctpgwn9883RXf2WNJoWJUwnTYiTq4PQ5CEC+yzHQymGhy9wRj+IdHsT9j3ADQUS
NVBNRt3BbUqmCoTTwNfOJEGPg7YtdmINa69z763QtmYa34mIgnhs24Qql+jXqvKB
6hy6+qLICJR466SFJ7+f850BmffT1uituakcaRHLLE2qxfUmkYosDLD9sC7FHDj8
igd2Epukv6IsY1BnVW9oVRlOYEbOzdQUkvU0mT2XJWpvHIutxAVfrPYOvA4icTSi
860XVUAJE1Ls/Jjk6YqCZw9jrZFoJ16SFVk6yArM5J3h7/j3X9+ZVAkGInR/0neM
3QUQpviN0+ZChkkgLxTBd206x7Im2LzWGIfWkq439HdvJxMX3nn+TILO9I2FVjmA
fOSewWg8Z7oNXWmwXsrc1HSRkzx/GPWEtb+SSOgpCrS95M6fZWLpWDb0eZwIB9JI
Nz8e9qOqW+uuLt/uReKkNnoPCW+3+lsGJW/FyzZx1X/uo3oaqFqDSN42Suzn6xyX
RrDmGR3aTnQANREOrkWE2ijqaM/DL4cAJ2LCBmw9mP2sMdi8ZkzIIZTxmTgrMMQB
r5vC7QpkbgcXyM0q3IHQMToELsAJiOpQGGg5epcMQaOzFxqQYzgOjgF58ceNrxBz
mfdZcrRwtO2Z/I/3bapiti4ATJwQ2SsTYu9t+jSOPglt7rdb5pT/CByXu0hVLJv8
2Du2ifh0MIGflYxN2LnNTcY/Dfsd5a6xx3uyHOnobtI4+nOiGNIAsPrO6X4lxFJL
zKhAouhwVeuYVac9w9US8v4Qx4g8TuILUCU/oMCAOpILDd0VLqKcFq1THxZojQmg
1UkqHTB9rpaYc5c9AF6rl9+LhYehllKKbIsusyucXLrjdKG2LcvP8EQExQ73LJq1
GnmgM0Xm2dMuJbwj9uzAKVT25NUoLJwjGW15v4PTKSLyVvrB6OnjNr9MMYtY1J0w
VA9kwI1VNICSd9nbnBlxdMKVQ1GKcQJslcsMG1VEiXEVVGpUA6NAjVzodATAJ+wq
/C4i273XhWIge+zI4SYXdp6HNT/Hsn3OhZ9E38H5KZ726D5mQbLGMDsuT0d2Ves0
Zp8HL10lg/mKs12mm9AaSj9KoG26x+oZC2+aSifMu4239IDw4vsiGGNNlymB2mO8
Nv/lhnaCqpy68GnKHfHzWye3tCOsHG9ybZqTpBceOzn/aTfZTRVw2wDDIbeV/bIA
e7OBH8d0Ur6rKML4NbMqZp1sOhnbAJ3YvOfj4J00NCxjkH9IEFhvMVPQoPfQh/Pt
MebUq865vOLZ1QBTFaPyHAeMK+FWVOgQljHQKU44r2HZoEoIvSf+XpccFskTgG4h
UVZppaeM5KmZu0P5y+4N7nUrObvB2RlUvOhVELfhpHCnEMWyJULDqn36dzDwHm2P
BhJ1DjRJ3/GxKvgwy9UyDhzsBcVEAO8c/OT5iI3vA3mkgvEAeaPovQV9qAIoNIPJ
dkRyooqDE0BgJl5mwQ0MqZlth9TkWW/jZJT7HQK8Z8eLtzIhuSH0CQ/wgBuiG1/b
HT0k6DeXvgxI/LBO8xiaIXIplIwOxFruY10jT3cngDZT3wriMFgVEu94cQ0sTnAM
ov1yWXkGaPj5sScNq0bgs18qXbwMh+Ap4n2luMJ3/sQNrhgMaEl4pO0YhNLAWrzN
McgRxMc+jmWPsGH9Lb5amj+067bGcLUDruCxE4ZXw0laDatpYscRYcTsJIF3nRQb
mw8uKyxFN9pvP6Cj/cCinifdL6z4S2LxcNHKAqpBQYfmgX0s/jW5UjXuXaYC6bkC
l0URCneVkanSKzmLx4u92dOf35H+J/7dp+BwCAe/1yYL3RFH82XtkYGZm00KBBol
J/u6SP0tcI5ft4euYhiXxKZavolBWMLmoYjY7mkZ2+vXymZ3G8CBEkJrJUz9wLJz
k9Hq/F9Ljx/tzUa4aRXYVpubMxDz+Gn6zX5Xw5IfUCpE+gvd/Wj6trSaDiO1/WA9
Rp5YB4lgfgBlvnS/LT2yhui1o6ObKWxnK/pbZCTuWVBnyGgonFFBoj2RPRi4qLRx
4l5zZdnRxuM3oI0zS/r566l2PQ78+uSbyO4I1L03JX8s6z33XrY6X+z1ZSoPeJRG
XDSlTFMDYaey6IXqt2udACTeAZMw0WQSAhH/q81+6m6HT/fHp+bh5rL8EoPGeA+E
GL9PwuDWtrO95FZX1RFtUAwmz/zjgq3GDQFj2jlVjbLziNyqT/I4Jlz+Oxhj+iSC
ItJSNN7B3QTCHKDzp9MUG+YT3kUxlYwNNXqPqkzTDYgLo+qniXGj403P/WcNc/Fb
1Kqk7h8K81lv4U7KzzyOphIHDJzS8LYl/47ZYAUXBi4VSj/fyTMV+T0ZrWGhgDdQ
MTB0DBS6QgMHWd1UIqriDNaX/udbaRg7j9PyxXCiOCfWPlgkYNqJRKGpydjMR3Fa
mvi3djFD4S6H8682AahOyq8mMUk+t7LFPL9CfN8cgSWOMe0Q6ionDYKk3NRpRpF+
vq9YhSq3O2re+qSWYef9vSBxnkXr707vloZzl+yD1xJxZAs630jgsGF2mdEmKWyC
idKdda02oxj6wugbqhvRIvhVXCEE6gTd3KErfc61cBONp4qzo6VVyJyPLeFPdLuq
yvJp7OddMwzd7cInv6eDHF80Wms+vI8h6MbLeWiVmJk1KQBZLO9+e7k5r6IiUGpT
5ib+YrS6gJKNZw+cpv4rbM3rHG/gQ/8wHWS2i3feFOculwo9eBfg7Cv6TcMDx8On
vigd+M3VKkFXpuL9nEIagw5LBJ4xtYQ1GzlhzKJwvzfO4ydEJcX3gGyrLw03QYvz
oVt86AiznDFX55fSKMpvrB2a98YYN6WCFgOiO1yGnIOTIai4GjU60ytlYcifTzCd
OivXlj3o2blq/iV80U4J1PKmko9g3EFhl9klW1K8HPPN4brEVVFnZsjL4DANjgmq
wfmhD0KBByCq0z1Us0WwRRJL6D3Rtam+mpjXAu8AXxK3C8dr+6Btc902nEXYGzmh
BMQk26FGT0+/+5B+Ik/oO7FTPyFg7/FbXRVl/6qkiZGUAXIIhz7OnZN4R1aDU1jd
kI3L23+TjsnN3pdiU3UEL8SojmSwPW0xszHmThJdY2pcu6NCfF+1oYBz67e50vu1
CBM+X2TMwwD8fMqJaIRUVOmmC6GLIoIPIw4spz7TPKvvMw8dTdgKq9seFFtW10yo
+Tc6Sfq3j2nlbBOF5Ak2jFPqrFJPVe644sfBy9Gdf5Ar+90uDRA1+N55N6c9OGU4
PHwoNpa0RhRWAawqNbHN9n4wo6QH29T6mudG0yje/GwrZCJ1tw6hdSKhtSuj+8b1
gouGZt9z4mjUTjBW3KTGQKGPGcSFx7/AVvX6ELGfgwwua9xDsu8Zw6TaN+T+PXPJ
QcJXY95nUMi1hYRzGbIKp3tFfWZkvRNyhG2C3/+iY3UJL7UT9QB9QbZTdnMBAnLA
mGkgT3NuM+wVETBKUe/bvTj7KNbe6UST2AVrIfwk9qvgRmTD4rAzoMquiRtaPb9F
wq3NbKA1mUzyenaBw4V83ZfNuYmiQxSQJLaz0DB7TJbM5uoBA4XHtdOeUdpuzXuS
+nD+hzP9LSG8fl1DtGSJFl/qC7GiaSbtO87TD2esvXTjcHJ2XIa1bXNwzrXiTPvv
SWR7lUQbnSBDXkwN23pM4u92RDNhEgmJvt79Ho4fhNI4AoMveRyy3VXxdFxIIvwn
YN4wrFonuU+f947by3JymPYAVb1jBychGqIgVC06Ta4et1Vo+JMJvV2z+C2MZYf6
TBY/J1lpdWcRPo8Bni2IJBkM0cc1n+5R1Qi+3nYsJASy/b3xCE7zKvdCtXGGnWIF
Kve5jhnPa/hT2AXa8DAk6IqVwCbkKrmYD0BTH0oXCOE2nAX8KRtjMRvFXZ4GFa6J
Z+BHF/9ZwbL9bb4NTEpYCdyX0MaxN09QIpmHcgt5gIV51XArBUiHdU3jCiGcayuZ
vBmnZrwNf4+TPZM5Qfsxv3wf3LfOr+heDx8l8Rvzx3So49gyF7fRHxDc+MgRSam0
owPdmV/S0fgXYOxozRr9Br4YOma+xcXZaxLyqpvLqLR2FahmMCiLFPNdzUmxdEZo
ddEE45597JSLAWF3bjdHb7D9629ZW6sx/imv86N6CzY=
`protect END_PROTECTED
