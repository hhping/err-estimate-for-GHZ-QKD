`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+G2xtgwFPuUmjgrZY99a4dSrf7cnrjKPXuFi+1M4xX+m8v90662SEfifJp7jGCmw
/+XsPXrB67K2x2Y6Vuw988yBJaWQsxGmipcs+E7VTTic2QIg9GnElAkfiTSbKgZc
95fWJf5JIUB+JZYPn1FG0Gl85uNk0L2GJoJrtXpJ7048ISHb5BuJ6zFtXCix/J3I
U4swIlQHvkG2pEpbhVoiJZFIS4q2mrtG2rn6QnAmlHiPzTEEQWDAMyHLg4kIjDxT
UoXB3FZJuE4zhaOH5/PFy1lAw9abNK2O5btwZ7KYjB99Cl7E+qRuY21RuXWx24xX
x18rQ91+KSPPWQFjQjb5uHEFCJQj/YpOU/IAR8JDljiC/pXTP79JgkzOlqYIjPY7
HerVpAdzVnE3lOnNTCzOxW8xbfAffnNJCeFY7lwRrRNE5XwVwlawIJp46eMz5nRR
TqTHiStJZJS4jNWaa2EK3waWtvn2Pi3cpT54W+uaf7hkWbnBgBep2xAGqxQLzSNM
MUDdEKNm4ozLucafBa+XN8qDRBT49oZIvoj+JjXeqEsUl0gKBk/HtHm3/igI+2Uz
y45ssCMBz/8ZvF7NybA2+Lrj1Vs5Jzcpmj4wdEWSt8woB8FZ8LHwRkMn7DHtDsRS
0Eh70lCArVjuvWMyKuttztATo2QJ0wvUZoW7o7AUF2wuKArvYwyy5EkwcvBUuiBN
YpDFho4Zxc/Wdt3XG4B/oyhnGnVtCit46tjGfkhWWc1l7NRWUgjuF668OprD9qt7
6esnJL1y5qYv101yAHc7RiDFgzbBT6yqDiaICCMJaX3MVF4jgc4c5aMk0FTXzgJn
7leO0d40QyMZRo/OAM5sIqxG3GUJi3MBqLZrp3z0zA0lX4oogWYBWKJKpHdjOWbq
47cSuK24cVN8RPhICkkxsDZFUHe5L0/26VeXiXVlYg5XHFAHw7LqrfaWMHqxjEr2
6NMC//hvJ8g7tsSz08Nn5oFFKcC7GIOfXSoHZYB8KObABpQ8n8cZXB3iEXBnpI0X
SpFs1YbWnghJRJJa8VE/MtCAg/LoESeBVujZrqtQ6hnMECw6nQjMHMad5/O9nUTn
gR/dDylcVzQ42FYjDTiyAYUhEdVlJdcjoVX6v9m+9zkOUPdxdz+7XqPSMADAxyKO
ccAbk9eACD+yI5wCGf0jkOUIKjyzyWWAUwK7kfBH8eEyNaSWJ6oa6R2hU/ypRMjn
xRUadivnQfURxNYwhB0rqjPHOwZSbz6psyjxVEsuXDR09Vu/YyR/irmKhVCISt+a
dD2x6/6AlkXCikqXxj2nmhUpTLW/pozvUS0DEXJjCRSquB8xcMZs17cROyYLJ2In
McWbhuy589rymP1d4vcBeVIPTwmhLQuMd9Obhc+UV7AV8V28S+DeNFLlCKX+oOuR
TCsa5zX4BaTKGmb/yaayy7YQF/OiFEIebatyWtOuqsGA4jl9DRXwNhntO5lzDl0q
cipVtjmQQSVASAxe3ZOrwTIy6VGrc/ZIyHjt+TdJnsTvjt85K5ns8HV3kU80e663
i8n4Y9V40puMIzYCYYxQkYqwMQ3PCcHtCwlnB/xvW+oR2XDbR7CGugAkUsYMjVrX
LHXhH2Y/95IK1a0cjLWkFiOcUZebQPSumlVWGj9YgBaAr9dBWFBf4Zp6i+tJZGq5
NbQ908SQ69Fj3D2V6OloiWGMsrQP5Qa3TUtHrT8iRoCllxjC81WzeQCCS7cxS0CL
bHQc6S0x48hPdNuTFRBcRFEMI+IzTCKcZfvK6yzcD/aKqO+Fw+Q1LTiEen8cuHVO
t/Y4FB3jjY5O5yDCeSOpZfDp4C9b3KhTadi49mnOqPkXlfxwXtI8UH+s3UyU9IY2
59MzHWPnTsQhoafUiKrlC98b5kOSCgTO5/8px2e0ue13g+UbAm3HRgT9CS2kUZuY
/f1DDya+Mu87fNr1LVsoAjnJ6y6e/tIxhnT0OfNXQWM88VlHdn20U6cw19Lw8692
`protect END_PROTECTED
