`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i6900XSaSrSTAG+xcp+Z2nAsRfear03n7A14Km8Ew2L+WRZD0YAlK5WRcZnZpe4z
4klYOfg5n0X50NvHv30rwLYyCFBp9xmXQVfsb3bC9TNPucS5Ibr/+FG8g976A2rj
xFYq4WQLPCO3Yx4hG//bUqLjn1Pst02grtfoKYoL6zfmlpwBtp31oUWg5rnC2hA/
DqiHGAlunsFYejLWdD1Wy5ZRH0D8thhXl+eIfIhgOv3TFnkMw7D28SFbJY9Nrk86
MavE+/WZlfkK0xo+ymxGinh5OAnpZIMnLn8Y5cGIKfQy30N/yfQ/bPIRb3owdL3j
uc7grOFQckQFc3BpdzsLgG9ULIc7ddFquDQv0yptfAMyadsTAeaJ2QZXa2RSVlTQ
fanEGYqGhdEQGBy+ag7IFFJYF8xJDMZj+CxRl82xXFKk7xW6DWCHlUyYSoxsQWom
zFRt17U2uC4RCoLRYgjesQpdC5XelUfwz0yXGzhbyFA8XLkSNGOxfapIY3+nWr0t
CHO82n36s01JBBDWtMDaFSiLkJ1NhpkrQ0icUxZL2FdUjEHvXElWz9tQbdL29PQj
dGEYxJSqqkYdgtbWiM1M4p9UwxNCj3sv5E3V3gikHlYVJRatxdl9JhFQYHOts8uh
FYxEmO/U/hrr/LLUSSiOSgDv4eyCAtQIWGoarAiAd3hH9sXcehpyT/CJ5rGTxto4
kxpoFEzG2ikehVc33JO6Ssxlj6WLTC1+v3ZTyGih62l/ea1xWM+X/ZDsOIQc7qhL
Kgc7BgLNE1l9aurlh8NxBFwJM26CeBVLllIOedl2SDY4TqQ8C9yeLiaeIaxguiPp
4hLGuxriQT/A6/s9b18N8Hzj1ajYGphl+g2+opY6jo4bqoKr//0+HCSiDNneDnc6
C4DaAO5oZhkoXvt0OiT3BoNWwH7sExqERZ2+7SPQ2/zJTsh30noMU8yX1tvCl4BL
UeuYaSzD/9xNj8ZMNDibOc5droPJkbUzvmmjwRNnywQTuJNFgFi5grPfNWToKR8+
tI7OTS6v3He38/t0wpaipwyKCodpVRTlB7mPGfmjwMUyIDl9r/Rnjk2er+2EsneU
+EzfpoS8UpRBguceB1JegzLpUzZXwx4i5Ru4LLfjMNeCz0vYRt9RmQn+lGG1pvwL
Qp3z+R776+4zLDG3NcPHUPUnkgnP43/6C1BpHtGQK69xgUuc7O5rUc4WtyMJEqfZ
HLDRI+lO+lPtwG2SvmEp710U631mmrqfYK1ZjlN0YEVMr2RKp/Em3AaLOe4kw0wm
DGCGtq4xQapdxrxd39mYhDeO/z4Z8FIgWtCLb6DlbUQw576j0UWLPTs/NWjgX2NF
JXmFYuq93MDb2TVxZ7LKQdw3fapd0mia47oe4J0k04XNk5yQ4KAju7jGqvJ9g/v0
Ls0hVD0pxxA47lMROIA41ADndGGull7eiVI8BciulJiuNrpyl7V/I+EPYlJaf2sW
/90MjG59wFFRXS010isqNjG9NTNtMDecz0pP7G3NDyUgF0Fh+NAXDWZO/rsvfUMi
n3CCHUbnU0Lh5CbuCfjlD35H8yzF5Qc/cxmQS/71ZE3CirrYbn88GR3EBezUHQpT
/CtUsnHEai3lLXKgV2sriZ3Iv87JDQjP4Iif95A5EAOJ+FY+/GYVUVLxDfN2SIQq
Je9XSIDy/2m9e3nO8VnPMKL6YGAqQ5XYSULdTQ+Y9hcFUQlZdh920moOxFQRxXOm
9gFfUWsde5CKUaDmyq9q+xwhI6m157rM705cf0/gRh9LOEYByClqBL/yHUT1oIE2
SHOMC8OQhgXjXgBXaGdUiM7LdY1/LprQHRWVIr2pJOmisdM4XfmWcFU8kGxWVUY0
xfEMOQxw1rwJstI3/mW7sXMnOyj2y7CZg3jRmvjjGStYq61Zu7r5w5srxVTBF8XJ
gfaQY6P9g3NubRAJaa4bNVzLAAIytjL0ksyw79pYxA+mA8KEuqmazCvofMhkQ+1e
brhTbmxK6+BlNEwzNhQ4VQmX25zQa5qsVHNlLc7YE/Oz5i2HqSVfKdntq+XWdhWq
+hxs1dNffaZ7PT66BqPns3QB/TeCkdMgFKcyaRwrtVJUVgAueH6Ryjh8UpCHwBlJ
n4tMFzD40qEWobc4eqi7WSXXin93u4n83z69jnCpSJxWFcz6OTDOCVTWCu4PkhJ5
E33TqXGZTMigQmO7y7SjuoVtbqSmvJHBXTvyeJXU8EhGnuQXQ54D+Nu1zWTjKVJ4
zHXU2uzFyiN/LvW2hThwg7CZF84pYPhPg5PUtQiMXso9lPXhZBLlX5YV7cXUBplD
++FvMbH7Licjj8E5xl2YGAOjSuVzQtHBwNrQpESeaLrxXoLiuPn9XW/7QZbwQUDI
OIj+mA5e8/3Rx1mtiGWxqI9q562RFVovJQIYuXQeFj848RnnnWeEY3CZxjCtxB9S
shEhR/C6XCao0n9tAqfwF+zh37unoX1HgSJ/4AKkW0/crAh+iogVWv2P+2ikWP+o
lpK7gp2iHQ/jGJKRY1Wxujftzp6U6SYvPi6pr0sO+vHRh6gGMzRtpH85aolpZvAo
GNxhceECRO6LM9Ds+DHB2bTsEiTv0vBu4siWs+I/502iFTjR41PFIv4SHyVXx8Dv
htfxHglEUTZMC2mNhQ3u6KetNUJ3JocPWH25IsMNcC28ciiacv3c5s5N1zKeI9XU
nMGK7m30xZDSyjfTBs6VM0jAU1Dso/EMN3cTHcpoPkTE5MHbv8Lt0Ozq0lpXDJ7W
QfFsr1kELzrEQlMADQNlkPwdrIX3WP1erlEkvj3+DNVAsi6JQSQp+0fMj3EEn6z9
3QIih9uBfl7+/EtdfGUK44Y3BbsIUf0htv1f0KFmF3NzuoZkkhL9d7pgbJ7lL5eR
514Te1+VotnGRKqIZf/4i0A1+lIdmXd2gQE1aI6DQjtlIAb69w5R2732LjEDuiRW
JwLu8LO8L/w23mCQ/0MDU49Q9MPuxFS4CTzuEU8yGAvsq7djL9ITFRI/Jp7F9B4a
jl02THH3xDbI1krkWSulPEVHrfVWuA/w9uWt9ajwLsObVKXdRSJKHt8OlM2ixwum
aChbpc3QCW9VKeb8A2uyDQkCtm1WmfDubacI7DDfbeQ36PmmhdPZRORRN0EeTn7t
RM4XZmgcreyhrraffhcgNcF/ProuRo4ZAOZceVdoKCIDJzP7yThjy8JKRPeBmicK
mriaed0xVULAC8iXwhECcrro7fQ/KTZPIX2a8h4UsvWZzKcdIAtqB9m3X0n80G4H
9zCak+ekQarfYgD3GEpzTkRpCnwMSBNpqO4kHt7tw4WgzSDkcUZNC8MAjKPdRuCM
O3k92GcXi3tFcZWa1koIF+2UCSbmfP5zdJnIZj78+jnnBiu2JuK7xbVN4yM+YP9l
gRJ+O922QdQZqr5xq2JJI1lw4/u2Qq26J6mluijSNdIOLOYspwJnOYub0DsaoC4B
bU5FVJLKom5X/fdqPjs4vtMjkVAmIAYDA3TOfyP+L10eN6DyBLp9TpWlF9uoeb02
mVcbIDDk7mrqdJkeec/q7i5Nj62eCW6TjeiPpU/795Q+E/PPZjTdBWUfOgaDLseX
NTL/NXo5qIibij412e4JANmuJFVctn0wMGeQFHcFFjzdT70EdfD41W9+s4gNF9xK
LNncbdXdcKFXfD/NpXIq2hpcbytYFQ2OVxl/dDeJ1/Cis7qbsaFcpvlg5wxuADvP
3mvi15HOmasrLGVcQkIA/2bXbpo2BWKFInIzlOwqhlSzyibmsuwKwDExiH+Xtdfz
Y8FpAg/wVX56sEuPtB4Ha6ljDHko3d2MuZ26hpcFIBAPUJuu7DgcRp9QMQnqNXwd
mYjCWgzTcr5fQQgd/tgoUgmuqoDhRmElOB6Jv2K9e7yU4hit91ju+UQUKXWHK9Te
TAdMvKDo0huv9kmdPamrvdWAT2DB+OTZ7aBB6dAZ18B1aO+DtydjQL7rtWvLewHy
Vxh+c2wNrmM/06yMsmnrbXw6PL1ZTVTlDN4/78Asu8lZCDMnwDOjmurar6O3M8IE
w4DzrD7ChAg7onCa00pQ/w0VJxbF/X+w9vIVEdEp7yzSvfcTKt/4UvqXElKul3bt
TYKkvS6Q2Uo8FKXm9O6nlPCTPEOvHYRwdnhveehrf1pnDAd/fwoFcjnGqlQCm/20
ufpaTYie4yIrEX8lnFgewvspLMimn+afOPavIrpBlBRpclBOhXpsmTg1DxWvQeeu
K4BbOWsuviPiA/DFWkHq/3oNZBXdWyJf71pvNpziJ9S00CrLn7U2UH7TQEfUlAoi
L+sXBR9eLZzeVIXPGQjQg6iZEs0kG4f10A5NaDsk7v9AUPTLLuOyssWxvHNTnqSZ
JaG9ddesCh3tOVdbMvX0x5og/8wbJ5vfDqghFQdAMYHtbQ+0zdtkK9q8hrBXK/jp
/2DBFAEi1unA7R4rNLc5eIuoua6l7xzB5BU3M+5k29e1i3uvGGoJIKR6WS1uUkK4
TCso/7HAShUdW2xpBTcetzwjIuvtcrkB4pbxdG1Njh4pw6pj3gN0bziA5kmyyFJd
Yf+bvmztj5gWOkROblp0s/N0vHwWJeW1/SvsSP/rATnEYY5GTfe6LTT9aeYBo7/W
6h8b21HZoqzkdjpcXICgG3nKRaqQR55ImUvLsZAD1vfoRS8m3XMLGUBxXX2FzbVh
tpcbxRCQqVXArev7SXEOybJHYWUHtl3wsr5Hocp8VkF21nA99c4QL1wQQMQXe1Dm
AnHsIAa7MSW1eL74+vI3h+zmATEKyk/BgeQBpcVBoWPoFmUjNe7GiU38GE57x/HP
NuE1m7GBUiaXgRFIUMzGbtnbl7pcogVfVbarVrXC1gjo4mGJaWVN21+sLaY9QXGS
PUB6S72FluHE6QTIXg+yO8RekK24GMpjc+d9fiF4sAlzcKSuWIMBTiauGVmJvQG5
UCsun2fu4uxFBw7LRMT3Y8VkH5EOTyJt2eDaOF0JyvL0Buo/Y0eJTBw2ybYbdOLj
etK6StaIm8b6RMnK7waBDrCcUwDnrELIYLHUAcw+7dCd3RUV7ov9szEyipWAPvVC
N4hREd0QokT+t0ETHgkLbbSG2sj1dR3Lqz8pXQzVVYJ2rm9bKUqkJlaQ7wvmHc6R
2N02Y5Pg9jgZx8He66uoxPdsUUiD1zOJCtoONXIplY9gAvP1Bzj8J3MkxQDjM6mP
WYCKks0pXFE9IsBRbxsJSzarEOFoQDFqQhpXlm5q6MrB2Tl78nEl6geFqihkxpGC
dWQE+IlSUrEDeblCNuqdGV0EUiVcrIY9FD0zFReeEhESQsYVaGvWnHeZKeHSTTrG
YgmgIFXUI/xkBytSodRPtKMMRCShU9nED2JyGg8uJUDbXX/j0QuZPAaQ89WiHZL+
Eun0SzbAEbCua+KKiQ6wmECnbEUAb+QJUOI45aNeE3zsg4snhXqGZGBfFeLkGhHo
x1Hn22FRsVqWHkldjfUVythGXfij/26DpYIYdbip/pKrxExBOiHWrqcxwsm7Hhth
NunM82lyxj08PRjYa+flXPhyirUGTBI8jmUtXsKQ1uxBvc+sCAT2A93dQohHxwh4
Hk6qg0S7nmva4Wt885gTunBPlZKlUDvvy4Q32N3NnteiZQi8f7yjIoWV08A4PlgJ
7Ke0F2oaecu7FonB2lNkPmtWMGNfmVb39cK+tu6+D7W2rAj3xjljWnNkvgMFYK+N
6JmQsAYGf6/j0Z0V8PIoKlobFj0AxrJRyIwxHBhO3jE3HTKQDoTkbLEzIyuRKWbg
er0abR9rNGhcm22Yb3N3RnoHLDggrAxwL8ISVIg+V/bOcq7qSl3wYKmjFLL9k9VR
55U9axHrEomyps9jBibV5vjKHZZC3lsrcbG06AG3lxL0YxGcr6M4XkAHthHonHjS
S7T+aiwDWKdo/+TYcQEFTu2K9giDuv7Nu9vXprEwOrTJpN+Uo0bG7mVTZREO+9F3
O4zkqHJDWZ9+iDP2vZy42kBZwYJZS1I+wqFwL1Kv1CBrCBCYyzFbMepNDFCloNdQ
EOH+DGPonncNiUazYQXaU4X25qA1/Tle/pRgsP+dinQD8txW6YrrGgqFTCbhF4Yp
4k8ufvSTOk6ObJz5WDnopyarmblvH6u7fQWpH4/rV98/E3cuewOFIEu9PDRveCJ0
Losj6ggcGPgfd7CclRRY0DIiSR8skMU9lQa+LijBzlqi9SXq754NRw1zJUyZ1GEb
6Af4w/pTgVavCrXuy9Z6uiwgSdTi3AAuLkH4s5rMdsEWe1eDCQWOF/7HNpgESK29
Np/8Lx/eqidFEtuE+lspwKrPZQUucLzhet7WzULRSeYAQFG0+UDfEY04FrVw70/m
PTMlwu1wKuqrHFgTwulWiV2SA/FA0WL5qQ0F+iytRg45b6Mz5Nwqs4MXEXXRiFcl
ygJsVK51VuEdpOUeq4ROl7MalzX9qFSC3I9zjxyGP7zuESucC4ThCzIQYD1ADaiM
EUGcjwhaNkzSku9XjwVuUH6/A2wbm68nQu6zlPQ3zXVIVsN4Z6GEtPHrM0KtQkpA
eZZbv0xmc3KMjmBx2LizwuYGAnojIvGBLvF+shIN/XtpwcMntITxKJ6vGD+L10Z8
2ZwpH5Ouf0OwsALDZxRCYZJo/9aEBAPML+iAZFyP2Kfun9w6ZcVUpgY1sSY+zeAl
BZ95qK4GsHsi3UN9ZnUIfWrWjf3FlcMOiq5ZptiLpZgezo+GGXa1U2a10Df92a6b
gtRzpK3aXDGCoc+L3kFJSoXzwju7Bhe+IAviadYSsEPef6GdYofBvtVVa5fG49w1
RdpiCnE9OuxX7Q58mINhlHI7tR7H26W/W+ljiCxLu3YDtLkMKx3hZeYI6oU0EW/c
YKkEfgTxD36L0WvZxg4LjLzxky6azrUxsh7gPQQj7c2AfWrEaVEjGMfF7Tj2Paa6
NdAlrSkFu3yDcVmi289sMdcJNJUu/OOAV0txBWELoo6k/UWsSFScJzdN1NSkdnTd
AcPdqjnt6bcpH77k17415/w/Wvyh7Ih1+oNpdMjzfVfTb7VsF2xyINtYbTZrmuGp
o+Jct3SLF5gyQnkhziL9qkuyonm40APdiPOsW8MWDhm678cwnNpZI8YCFEbskw45
QPSbwYs6T+MM74LUdUTW007XNflXRzTL0p/LW/3jzpOoeTUa0nFlN0wiklRluNRU
xgsJaI4RAJkmdKhOdbpaJL7lz268qxOj2cxKFRcT0FPyrtCUT4lAYINxxlwDn3mJ
M8j6vNWu8wMJWtNsM15lPU2uMnC0/Y/CwLexbjfeq8m0XjfCh0Ijg3lnYGZM24vR
tY3Tdflg9YjYPlVRa7anQIST2G2/BW+k4H+QshH3zfWCwatc5golzvIJYld31yfP
pzBCKK560RGPaCl4LYCciXkFH+y3NPlX70FHi/ZJoXqI7iHavo935rSTbk/cHHE6
G2SRmLUxNoR8vfD+eX8DvLgt9Ig797ox3Uv6r6A468V3z9usMGC9N7E9nQfb0Sod
6haxtdBNK+OdPyocHJo2cK/J0VVnU7CEV7xJzZn6pGS+nLSFu8RruX8YaXbnDx6R
88j7ma10/7XFSRMrJI4/yepSUM0nepkpyKAXwbY6ax4jGEjExiZPz2XLZc+zwY5p
otsoyIUIoQuZwRqzFSn2zJHg3fOp/z9h8s2WKu13wnG8vaN7xoD6wf+G67Xp+FWm
/YfffYrU7GifYGJevxPgC16uRAjtz3Q6uNxLwrPR8nJR+KF4BdZ/Qc4O8sP10qpK
0Gf7eHTFb4DV99Gqq3tL97CkRGVZLTNLF7O6W41wEVI3UgKd6qoKA9vvfivn8uMi
pKdL+jbuj0RmFBSOLjaCSioyMLJ1e9NYpZ/R8GvotEjgASLk6mGYCOwCxUVyBIm1
VXXjLuUrvj1ov7s8gDsz33lK1waA8VhpSrrlrvmXgDOtX5CmJYB63QsNzvIQXCPj
WYDNdgBJZQXhONRBJ705fnkQjoDOZP2qCQueb6e7SeDiRIwqiYlLCPFeENlDSjeB
SXnHMJRU3D65W9jZprHm4RFcIX2LdqGV2o5ruby7EoJvXpa55eke8VYybo4Q0fIh
j5c70J2ogXPN4j34qK/uWWSOWekPRh+oo6O57Aao5izWI8CiXtl9z6I5+T4/bXyw
8sxZsvAEwspzIB4Wj8489FyUch6xp8zQXdbcmAy8PyxkEJJVJs03s/FjA2T1+iKY
9bv72r6KYId5LHuN1KL0hsZEtqoaaMN4+T0qUHI7anzO+j+3M8G+peAjm6d/h6yM
ap1WBiB7BTBNxv2wsUY8CCliOucdnOY8KBftV25pygWCAX2ov9TcsBhoc6bOjweN
syEeYxE9XnPGU678TXvAKyr0gGlZcUSugtqDvqj9yXgChjZsN5JWJlfcg/VSbQoL
e/UHDpYUXRXT9qBA4tuAAkb5glxTnsNOQ81QR8AuCFLSq2KX/vdILqCwSg6ZotIf
pmXt1EzxfS/4PtVzepgginL4ctkYNsI/Xjox0uVzYTJRlJ6lcDh11qt0Bh+5b4jY
wvYcNxysgYPpEQxSWbUFwT3jrDEeAXGVNxhMnOgeiBpxnDaXSYGnDL05rbagQIBL
fdZk/kuWfQ9dL0ZktCDZZtjRto7j+Hf1PXVM15sIc22DaXEEINmR079Ld92uQ2xy
6c63Cr71m8BKisDNq5dq/z3G/T4riHp+gu3qhOLWKYASSi3xjcN/I2PjEoyNVQTn
Ojlgje1bJzVCHyBtlDwnffazDViRIEC2hef3T75uqSdQM7Entlj2sGeySGFvNC/S
W157jqhXcaBVOR8DvKcf3wQ69qhX4Dd9cto5txe4BiL2CNiNtd+x4gh+VygVX5/K
6sq5TtkUF9ES8Ay9oyj9HBSrzXCBVVY+D5a0uFH4o6vswN/6s/zy4kTvec4nuSU+
npa7iALWWC4BVpNAAlQQ0SZGR3x55xjSLM4wKMQWsBRLaIP+UhoJ69slUy+n//cV
F+VOeZdC++NjMcvDPZKObjuLadjcTCPsEERXyxOc8okgEBpwYpY8D543vXGWDsta
nL03RZxRb42/V5Ntp23Xe28k4NSfzVmnMkpoaTi9J000YZSAPjrxoBqTPWL0uQcu
9mf1wMsSqt2jHGHcjr4sDaF+Qi35V9bSCJuS0+TJDkAPtMMyHpsAsIbQiIMTEuGo
bDOtXZhRy6tLEjm8xwxbSaYxLuvm9xjIoln+sfOTm0sflvsym97WxdBDTLw2OsNu
QMqmKbX/x9KsFx6mif2bOh2vHzhQf9RhWUINg9Kr4vZXjRersZhLzrrEIxjjNknY
B8NUz2TsLoc8538CcYFlKMM+J9zOFJjS3x2v1HbP8LrMg7a5m6GkV7ltsXVamvaL
7bF4cGhX2OzBqnEF0LtJeCQsV9CGTddSt2HQc9eB0awclUHSz9nSyoPsXDYJhnNa
8pFbZBzkLJnU4hG3E6APB7bGhXGWl3wq342C4KKdfdUJyasbD1U0NSX5MzVfr+vB
joZvwvJHrk2K9eik0SXP7T8AEgWPSUjmkps+5xeNVA0iZO52uvvz2z9yJK79ZuM3
ASln3AKVR34AoAZDEDD2RLoKS9fLfKHw6ifC9McuTP44JQpQ29hv9TV0WaEK/PGM
wZv7NzJOr5q0wht11HWOWsbV7sC2wNzPLOInCaO3e9ZLH3CTakOVjeiJFkS+dORL
5nRrD2u5qLrcrqUb9fHXbXUQ6uFb4siUmhF/1EZmrVppjjsMYbIBybDhmbsoGelv
eDSI/Jg9CcLVkFUAsSWD2DLjJJsiDpJyLxc9jXSTNQrl11ZFzMbSOCxyFnH4AA/x
S9Nk/nPRf+CID8dFoIQ3HX/Ko5b+aQC3x6F26eKxsvbrheNmwCXLxRcYUR8CTci/
uv6hqTUK1tuhNbJvYNcUAFt7fs4Mswx03tTPksie2h8fOL1RQyAs4FzkmavDwp90
FXt4eHSq8+IhGrteoLjSsx9ciDUYChY34ljI3/xuIxRxocznD/tm2rrH6KzM94Nx
qX9iXk4+zB6+95zWiYhAHap8vhva1jsE4JTeLHjCsQc3tALdkcXGq50NpOhGA4W/
qbl3BBMGdjwOGOpGy+3SMTfE0RZsX7F79CJq7iymzcWi6JIbzlxbqr1txYULsf3z
TkWJVRRwKZ5msXFUua9FidU5HgSr4wPTnOFZJwjCdDr+u4SqFmphhDe7KTc/+W2y
IJK4ZPi7uoHNFQ681L8JbfsRTRtulU2FwszuplRUu259f+kokP+I3KiN1ja4lM7P
C0GY4BddMLLVv83Uq1cFp+z8K0XFllVokFwNKr9GIucxBmSnED/BivW6nuNbFSym
c64Sa5TQW6ReYXvXasQOJ1O6vIPx7m/89MBhR4WHLITRazOUD0eLc2isM+ni7e1Q
f5n7o9UQmGMC3KUKb7GRR9EcyGy4TpsN26N6mUonvVmmvGszPiieKDImQSAL0Np8
jwuaxjoosQIkEk8CPDznTB3+KhJyvldj3VxF7J6Q3OdNMKWIRUcyove40/HJ22Pp
GVVc0rcQWqULGasb72Kc2j7P3rU3FBCIV+nGSS3FeAGFHy/c/FSwKO63PRrQIxT5
xS7s65Ly2uZo+JuhY0wQOCPRNnikz5WdSeZFo0RjH0Q=
`protect END_PROTECTED
