`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2jtS+z9wUCKiP+ehlM5Zjvu5aKuUzsGjDT6ldHBDKLFHlf4CnfpQbZIgdJT4lclF
ZzOatZvxGHge2+nB9J4J/FWHfKdRCiCDs/tGzLlaq6+PfvHdCuAfTAvonrY44jtF
5FXstfCZy/zpD3Vb/6VW5kQr1Za4Locjh1xvJAG/5KTKwj/kN+u422Or366iLgt2
aTBpdLTZKzKf2HK/bTlttAEB3slPl6TKjvgeeSCbvxYN6Anayn3R01rhCz1EB6Gb
cD4fuUt1Gz8uka3ojKhUaAld4UTMGlhmagACsdIJirmIelPlt1sraYvx6ghCEgEv
BKCe1OKSI0amea74IhRtiK2be2uZNuur2TPvmSc5Ny6cEERHi7tonvvf81aS8xS3
lm3QrI6nj2y71UwfUgriMjR6ctNCXHcz9L4OLiUgyTzKQyc9o8tPFx3WHsT6UxRq
nzmiF1lu301hZGULE0QM1s/di8I6i2npZohEymOgzpKyYxZtYMOU0JySMCZ0zs+x
55xLnu3dKzORaYs6Y9LnZ9BugGynYRIsLNpk9IIfdO+g5PCtBg5ru+h30IBjJPZ9
C8eo44sg45weOrJU3KTuP4Uhl8uTFF/Ad892yZiEIMj4GtMZojHxdf06z2fFw+2G
KO4em1F9xGYgXr4Ll83ry1EogGfC6xJqnflBMYvfy4IBIt6zxM52l7HvMT+zsqXa
DQbd+SQcdKESdonRKlOyYhihHXa11q3w9OCSmZyeVbHRL1IA6m+04jLwYZN6Odmz
ICMjrJ/zoSF5kZ8QmBF2Y38BuN2v0V2vHsRcrNdv5uEbALJpeLaGx8dAtAVvUiLS
jk8EgGpFnn9/Adh2HVAVn+k6Hus8rgecB4AYdQ2eG2WJ4rILQ5njlGxc/TbWZPkq
b4OKlv3j9Wq+yCJ2RPJt1/NT8Vqw00tCMkS+Dk93dEE7yVNVKWBUDj2GhXl6ri4g
3UO0QxyfVjXbIi0li7wmpZkhqWVDXkHVEw6GVVjps8/vYtpgEpbcNGACsz01lGAg
FlgWMKz1Ig52gkBcMUuEffWuRnv0buq04eSg9n0DD4uOXOhZKUIcT4b5pm0Ha8GG
9Ofllm2HwtrghGlCTW9xw56vMnr8j4GPLPGjaL8cDSIdQnUm5jXgRklui8A4qfio
B9/dyqdhW2ISLd7Iupm6yuBlvfJyiZDmIeBa2wLqELCh+ekepRBsvZ9y/T7mPTUY
8mu/ab+gcqIPBh2hk3xJ9yVrqjwXRfnuPjGDViCqI6/GEsyPPj/CbSs9ARZmLa/h
/CNVKCObzxiRexdWR5fbP06L9MmPbUtrnFqBbwbxjH4yHcwbEHXa9BnxMJqR1/Ze
Gb/5Qzey7tt929PC8SlzyhLw4/RxjAYVb+j5OOaBBZAjkE45Nvy6FSIaPBSeAY/7
6iIJpRMsDnxCDk+kaKYlsDEXXK2R/gb/+/+pK4kH/CBBHPhan3CYhNwCsGL9ppQ4
OYnqYZ5SB1snOhMQ1jYW/nPFl4IxInwHrnCih+C/eFUnyg+VdeTSQvqJFsbD4R+7
EFKrffm/fGii37ElC/Dvglo/eC4foShy8o2tXnaoAs1f3DQ9hpaQsu1EIw06cFsP
cwPzjIhb8dkkljOP9d6CMHu0N31IZAtpco0daq7rKy9QL3RqEAek9R72SczA1s/i
w5+6teswH8KrKfqe0z2Kf3taQYEraEOuVT+X+vO18MEoMN2tOlwRXoeFbhkLTG+r
XCy7KzdmC2tVCLKJqroFIf5dfXQ4/wjQJVBfZ/uwzYkR49EfmR4cwntR6rltPWyF
L+VLuwNsfNkjKa/+NvLe0ubXo/vADCXpJuaP9f7wG/iaWDNt8I8k3axGCehRRQoi
tIV0bcWQ5iMuR2X2k6x3+qGtz3N9RKkC1XvI3JMj6zpKSzgafvX8wP1PScyAtn5P
W8OzjknoYOpMQZQDNX4/pd2HcJomQRPgBm9+zckmQtiBFkEsDvo8CBnxkfAnAXz9
M9f/+MXW/neeU7cX6hy62uGlBC3T3wyFL+nUhi5Bt2cDGNPrN3SvpZbC+wPFND6c
mlcD8ugAPvXxGod89iLMT6FU574VgesbTSYfxYdJkBYeDwbhs8H1yqfrV2zRiZxY
sU0x46Ui+qhWTP8exdkdcinhzMWsFnccObUmsCKBGLJ9Qv+CqSY4+CPZhD5LbYhN
4fvaFMp13m8T83Xe6yj5QLVVX2iwU1BjPP4WSuSp3y4MfnGvXxtWWxR7f446Qkx2
TVwTZ8pq+/p76tpk303F7y16Q/e4scckAw3GVAaIUsG61242BhKqtDUd6YfKvx4B
zIH/MvLW1ABFQW8GyVXemO+ClcBSuPjtJoTpokEQaSZkKvO6Vgt3Wete1q3MYdFz
7Yd075//9nTFOQfHisKgdV6Yz1SV1MS1kWFSHT984UlawNov35E9f0d7n0mQY2gq
LTBkJ21uGua76hz++Z8wOBZMqcIzkv9ZgbVQP5Co7B3mr0rDxNFq9+QGPpLh19OG
X/dpc6YshcASz8gByaw/DoFo3ezzvVmVkD76Pg50XXVNMguwNR/jEnh7wqLGuoTP
e2lOzEGSdrbYgvlIno5cz8ijrybTt/7SlGYQBpLCYi5qCW74W0H/lQtLKHI9SOXy
CG+lCLoAf68sTGc2vUajPBQCifd3Jx78siPoNoBEVpX5jInOFUNEKL5EjjSAYvvN
kN5hBlgqHbHVKJrk5nmH0MPwvM+8hq9Nga0Hq9YOSm5gtkFC0f20ABrB6Nme7TjQ
VHGMBkiey3/Pb8Li3xoJB0FHzdZT9sNIkfcn0pZPXYq3haVK+g0h6MeDq6IXPYMY
t/D4ZoAVffdSo5ti8hu3Ep+6mNcOpRXVbSl5GEeGTg931C0YNGmQtmmRxq8RlatR
hfkFDf/Ggo6v81FtRHV72qchOmqxDUBfA4H3mqXdazTcq1xsfOaCpP7YuQC9nSBI
zvI+LVRInY+zN5u3QRldQfVsU2ona39+6rH9neOp5TJuhu8IS9MvaiIu9NJEAB8C
+rctiJoHopvghhBeZyWoI2U0At5xDQCY0ch0wYuhfpI+hF0vGfeWmtPOIp0pC31N
NSA7kzdy6FdpGMuNLPj8aojqAypL8GuLbLfpSli4SkEfRBfNFKEq9BO69ClGSmZ4
`protect END_PROTECTED
