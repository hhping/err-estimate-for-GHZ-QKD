`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z0wvNpzNF5V7BL+0IZnpBgJINrV0D9oZBc+lDC6UDR5en3CwCAIY+oJ8d40qWcxK
GBc+HmK82J17u/CCytdW5Gp+yTm8Wd//V+u40R82zLbSzxgfzP6AFSbsoe3pW9Mu
MgymszHVZmUcKABmk9IN4X7ry4EsIXV7H0ASMYDsQHWOApILQEq0/rS5RiFjF7Ow
049nkVxfFp3vJzABpZnQHndZ3qw5r8dhrhKRKeKkZPX1Can4c5yHPt4dGzB03Dc0
ZjKgStc9tjpvRWVL9zGQnyysdJgBfXtxsAdqC9CvVZDpaKH6I4c7+6RrQEawVag7
RzdyJpjOZHmD/G/Eb3P62ajUK7ag8DEwzN5XM7VxJkjG+EOpg1S3joYaMAB1Ah6g
ijnOOgkSUy5F7L/MBhpcIBjPgxzCaeN04v5b00ukv7xzD+Qxxim2NpOZJjhKldeS
B7SSgijyAAs89aIzj9VcsC4ocui0C7jhDyAZtJoIpykogGtZds1XI/srw3dwO4qD
+g4VnA+sIApVgQr7vNXHBQEaJZJXnc4Xaf23RFKJtmGnzz+pbwQHQEbDtht8k3k2
UMptypfjado0QUQ8ZDsXww==
`protect END_PROTECTED
