`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CpHn3j2uON/rUVEV1ZA6+HA7XOUxTZFHK07p0KD9LS0CgcDGGEPSYZmvyvCdZThG
WzdQuAChapg4wtaZimIYX3UWAdphKjJaq1QhMJZ0ME3JVx5ODt9suB3/EHURFgjc
ILnazNAWPIdsVf734is2sN1/ARd8rccO0fcH0fueyAVCzbbGBhEpX+dDpiXYSp3q
ASqvGRDW9MIq3sLPdFlfscaIOpKzmVcTuCLBbR5arm971uqNWUBiGHiefEH9U31C
i51OgkVpFtALSQp5yb4i6Ki/+1IWunC7dzvo/tD9FyNQekkczgpeVxuPVFcNWUTY
8bwkVm7rjdAMJKeWj3JoCfqNiTLM8gl1kvhvjrkbxSSdcxg88W+CKJHrmwXpgxPx
/xUlW3cSN5TNcrZvjvuStqR+HVBreC/B/nxpCG4/DQg+hfBdO3sDrWHSWNNUw/Zj
QWGS4QUiTO0wCUhwdA/+2XP3SrFx9nfSr4OuaWbVqriaJNCUJZJNLtr1aQN2XkBH
DJay4vuTqT9fWq8dETfizxR22VMYsulFXskej9n5M8pj2p341xT5e1zYfrth8n5m
XhzoyE0CPsYkBZO6ueNjK/rDXrzkGdY8w4iB2qzQbFMqputYOqbdMEy8DM/8QeIq
zBN4doPTG0M2wo8Mjt9eGAU43vqOGe1rbaYVet1TtRlYsKKLTAVduU4qzCqW+Qlt
3Bsz6tMG0gIBNn4EPxb5hYz94vsm3JuayQPVceIPXSfY91VLwEg4khuK25N1gAp9
GsDJ/gpjCwZN4NKhNwBRePDhFdSXm8s99uqmNqVEaq/t5c/GDtizYIJ1BtGBIefl
xkl8zKqje4gIOAh3oFtoDyChGABOx27xuQz/ATMT2/CZZzCVBjOFyNoF4cF/5pwJ
BW6UZ6qPSWA/ewrBOEY0ZlP3LyzTfEJ6D8CaJiwSL8VpfZGgfHR3KeIlV6xPdStJ
cum4V97cVxnpu0fTqlTtlFgbeS5/hlovi0ekkMeHhsNeH/8O23DdSCqfsKJsJ6U0
bRP80+KLLMj9mPOOYn8dm0IYU4IMc/1mynTaAvKK6bx8/Jy6XrlgDkoKok5dnuo7
CKvHMiIYpJAAyj3WK1p+XeI6ijMHQ+bEU6YwcUsyQVmenCva5ppXGEX+8YtaB9zT
55hp/KgMOfEAKFn2ktSz9ppzK6vdE3QCVHO/F7lxAxWEI50ewu8I52iYKPlRK5T3
oCh+ApIMnzr9Z5jUHPseSg0KVTnVPpI+yPPV17qzEM3DBW+H4w6igGauA9gFhSPN
NWrl0DDeWncIzZSrLdVek35uP1TRiPG++3KvwlAqmH1yJh+UkPK/Qrs1PVx0Gi6N
ZYKYO+IcJjQcJSbd3+/kMHgFkj+I+lKmUqKsLUpBCbPwASRhnPH5Jm/DYVDaI5MP
5CjRwIM1kOkGutiCRlUgYe1OLCJuyw7JPdNIjt4LiqcM4GBFJJV9lJVHfBw873SK
tGKMTHFNm9Fiqjgil+V8ymthUJ7d0FltK14saQYZzTMd1Gv89apcN2STI5AXg3m6
Kh3BIMsQ9SF+8mbOuLJ9S0iPO+R4PJrqtNt3AY/jtYpVqx+aN/ro8GSfG7ydGNNq
sw4/TOdkLnkQyDirVuyui4iRJksJUPXIqIB4KeFAMevn6Si9ZgdbOGdmhaOnpmDA
EijYO2NFxuap4P9/4GTAXIh8JVxBqwoXepM4LTJL7IKUzt8ySoCneCGcYEJQFxcj
puvy8tyrMZaucnovCP25pzrCofjAUMnqq2G46VtL8mprr1rXRFPDUq/qhWG2+emd
BjiRUNqemi09O4+QFlk0s0yMyTe3wCIpdx1zO8sXxWjs/qidMxi2trYvh6e9tO3m
s/QZoI2QFr8oMyh1IrusLMVSBwHq8ZzNcxHUIuT4t1v8j8HvjewSjz3Nvx/VIBlB
yoq5WkNqHJeFw35hh3vD7kxoFdRzA9HF8FLgqCle1AFbG8TnGv1Zf/p5XtiDBWDF
kK1WYPNj/HjX4TgK+CXqSsdzo3G4LrE6/wCn+qVLbvHYP3AxZlcE024qqLISVISF
unEvMeug3u4exmPI28uS/JZN0OFW0Ca1xdf+lPBlfOXg1WGFE6dXNKRYHWal8lhl
XYcLQj2skM7TZfTSMxKP5Gj8WEEPk0RnvPk3KCB7qTix+VE0nk46odr9QlBBB/Uk
s7z4lZMXV2yJHqCSyrD9Gu6VEX+R4niyKIWot4fJLQIdzoAO68EPLdDSo/wHPz13
BNtTCdeMxbBqNI/iSTsexJesTdQw/tKcGKjv9qTW4r4vZBgehXRfpZUIIt1oajns
LZ53Hz37hgs4VEm3t8IA94KHwmudYd5QdWu3cvku2GdGq6nTndLPjjFynX6aPZbW
19Kixlir6Tko9vkg0iJBJ9Wjz7RlF60FIP+z+EPz4dxLVqxwvfqTtd1bI+orzhBe
U9l12hHm/ly7n5TRgckGYHFjZVEx3d1/2HTOXpfwxmT23sHD/74ODEe+InI9zadV
OnfyWjstI+u1RbUsE8Mcfl/qAFP086U5BTVp4nkv2UWb7UqRw8TD4i96Oux/mpoZ
/0SdgC40l7DGedyGfcDDZjj2ytjIbrvmoRceJ8+zs/CNTHK0uKZZa6AsLZAkVm64
Q567jTxy5rKx5GTJhCTjZOxlEa29ndbwx0q91HaOlqQzE28HjvZfBRQopgCSt5RG
sHsZL4xiGiFMNPqDmOprgUUVuhdbwe7igDcVnRc5hUjB3MSUC6X9yKtrx7QoWTqx
KVA56IBylAEaWuDTsBoiSM7cv4gw7NAQBxRs8MXHen9kzwqSSWI3kt+MkAh4w6un
AAfVv3EcxOSzb06l2IS58O3Ga4IETVvhUdrg2h9/nET68yQAqt57+ayKkGE6DfEG
JweXxZkAV0mCd4lPERL38Ya1Xk/sJ29CX2kwQJHpLiOVBTMVyhP+axcP2EEgCO5K
nEMfdj+ikAodvCsrONTmlmizHn0ivonfm4UxMZDUz7DfqIc0KOgFaTDcKAMWDTGq
qCX7FemRDy9AYwuWotyZRBooVWN0mD5t+XXzyt9UTeLR25O0W+ZAG96koaa+ngsR
Y5vQQvFTcGkhCpBOz5WAp5icKuBwiShrj2aEz0aNFte4u8xo3VgVGk4QxGnZ1mXm
TQdyeg/Zbv4xqGfYbLGivAP4mj24guX6Tq5QNwMs3eNrBTz1VPvNHf9vu6YKgGYV
Z1Nx8T9X1N/Kk9GmqjkPRtDwxeJr13sapEeyia3Z39oFJTUNW+pv3Ef9tOwSDm0I
4fVoRmwaneRBaf00d8JHgEoiUF0fhZZ2mHs0mlLMmpwh69ZEQzg+amLfHuMwOSdh
uJlI7AZhJjQdwKNZ+aLouV1Xo+gpBu3TRCfXHaENjdhrEghobILBPx23FxIpciJp
4U491C5qXT4UJL+D/h5gJy05L1mkUzarPWYAQxSgkd1xpNC24gze8FCwm78tGHfU
rtvR8eyX1mVT7WZdc3QoETbYEFjCFMzO5dIm1ExLb7thJmhzUfqYAks1v2ms+52o
Oy0UkJdiZ/tDf7lTNshBxYjBn7WdTU6Kfdj3/E8XfnWPRw5CxZrIsHgNLvpospJq
Mgcp5xfCxgpPu5CZpZ2dVrx/siw9n4//aBKTvAR6p2dHZac5c7O6SgQLTbRTUr1f
h1fNMKl2QtC8VdGF5+kz4N36uBRFCUsB6DswoXLIYfeIVmcHb1dPBR71YxJKHy+a
tUWEIFwakn2U5/9k2oAsK2U7MKs+h1fueMImjYkSwJPQqg3UUe+m7sDBT2jL9MxI
JeyXd/DZAUpQDk/Akh6Ou0Ic0FPMYHGH5GlVO4hAVWLfoxA3y8+YdyipqDBNYfaE
ap7QEn3QAywxTPpRgF6Vxs/eWXwgxmjuBeCcpxqLKmAeX4o+yTjctoDOCwPfVj1W
DdhZu39mmmxtIYT+nkaaz+ypbWT+9J91UgURp2OksznvgCcRXSNY5f5sUM2PBfHZ
kBQZ55LGnLNgLb55CtWxdakk0sI35hUfumM2NeAGyq+wO7A0DrETP2vVLRNDYGJF
9WUCQ5phX2q9jh+rc1iWODYzITeaHaXBSuH73J8r8TUdrkGLakI5Xx+bWt2oue/K
rLvqRVmHLrcD0OtXCOYqdBh9EpEepa+8FEeX24fmpOU=
`protect END_PROTECTED
