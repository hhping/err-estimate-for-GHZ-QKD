`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6UpEBIQ5dSjg1ekPiqcxGDef+kqrjzkWoHjTeFME1787pIE3ezI/xl1qUnRbETSZ
d6tEmpUIPULko7gN/r/ZUhZFUk3Qm8EMzjS+AIzBqXpPmCmX6oj5f8lUhjmfmukx
j06pko0KjZcAO57Z8VU9leAho1lRjvNcfAY6Vhm4HxnrQ3lRgtwA60wPIHfpJm1/
SSkddfQ9U2iOpOxFcyMMr7Mni/llqERwzgT57Jvwe8fV8rRCL0RrLoQaZ92u0vck
XaMKqGTGEAr35SXVz9mEbnRaIOAWGLIyxnKV1K3atZltdZS6HgxSGAlC+ggFfDVn
zc1jUIBN3g5SZkZn3rDSDNJeAYgmZLAafMyCxMCs1Pdi4+zgmwWW/jEecjkiywek
zVxgeALZxnxB0geULNs6XGsGLAQ/7LtdJXzPC72wkzxjWWqLwH8V2jqnBwPJx9t0
sSPyNlYr0pnQoKcZ9Ly7sSmONQO3Zuhj9Cf6i39QsM1GEV4JdqVMiX91WzoYQSVk
HnLfKX8Joxazt8oqTbWGTkckE94XzoMvfJSfl0iZI7UaBPmAq+Rgpqd3S11Qu/yr
sYzqDaT1NmKC1wtOVI5jTlBnlBKK2sPt2C0gaLtjA4wUzndGWgEZYUwOGJBDrDNA
sEZggdpCDDAnF7E0Z6j8fSR5vnuGx5CN4bvReZI8mPRuU1tuFySZ7Q41Ddfh0kSJ
89rE4N5b7AERUFwr9jrkgM3ewECAb9O2iWR/9k7mUXR6sjujNHfRbbesrDdWM4qL
i5wEp/+WSGN+EHtGMSbIwCAraMjujasmPwuQ9ZpMyNUCaDcJDU4cO58IfJ3LN28b
rkkJBGTMvcGaSVZ2utPCF+g1fVlx5WaQZPMKMEoCYzG5A6IyLB/VRljbXu+SCQh2
bizqxDsw346DPU6xzITgfoPplGduTH3N8gitbAOzj/AEj4rt2fh3ciUNapExq6iB
/2YFgbBoxEF90GayJJDEMqpLyPOnjOkx6wixSgMRTiuOZtHJhXLwRKRh0mPdfZnj
wvzIrchzfhK/MvGAEBnqnA==
`protect END_PROTECTED
