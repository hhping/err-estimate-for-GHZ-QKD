`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X3ph/yMLvP5yGi9CWqhG1MKu8imFDA+sPGBFOOkxm5JYyG/D/9WUdhEoxcmri7ku
gwzsqrYiFxuHd8GqxGqH2/zRyRyZ81ccpQ0LVWQixH1JygO8x9n+EWEOg9ILwrx4
+n45Z3Y3Arf+WfFJARfoud0mN588vSVNfxXztKF7gmPMXCL2LaHG0eDXPB9AFKB4
ZSKK+N63yRk52VCUnNEI49WbaW94i57kNh4SuN5Yp//4QvKknXAUiiWAumoKcrT7
59e0C8ZOI1H7lsEnZGoCdkMQ+CFyav3FJeGEfp4oWIkH33f4ddIrt7L9bZFNLwdk
F4N0L69+fl9Y5QdpJFlBLswqx3Lr36T6VNDjsBroM7q9cDa02gS1QJNZf4dPBr31
NruM9ei0A6Wvroqn5Esm6HFiCRGiTsldBV4AIqIgoMtoy+fmxeVKqh7NA1nKYajV
F5MdaaNj5Afu4CiEHeegzO14Hq3CbqP8U3JNw+5Xm7166Ay1dbzIFeh7j1fDuDrB
Z6mh6HvXoIRUvj28pRjdO0JtAn6oEBc/ugmpKGcY5kxMN5Udt6JlNP4LFDivn89h
mcescxyf3f8f70l/8ARBVrgXJQ/u+MOVvHRXJf1ptjrw/FcLR8ygKWB2L6MpEDmb
6ptacwnioDWdP2DkUeUExpVfRHE0D7Zi0MqHEEBONPt6aYDLbyqzqDCeiaOufF9X
jI0UVIisg+j2TSKDhfIrmkosZ6ScaUsxdGeLDESYosuoxB+KFGwJzydkyUQ65tut
IAlJPth9wf48Mw1YoY6WXQBm7Br/Pp2J6igHphlX7YfBDDXSpOXLxJWSRCjd1YsW
xI7p6qgfSrfQV7dnGRdCKxnHJc3ZsJQTyJKlh6lOc/vdQZJjknJqkWfGrQzb7xFy
0PI8Ujyu3K4Lo1mtAZMamuuJbcXKVvlQ6hmxQOBqlY70CUA8d3EsOxDpx0cKiwW9
EMaxNoJFxsRZe586Q0REBJDVfGlJpFbLgP+WARwYlbAANtFxkffzH/2OP+EkWhZR
FiIP0kBwfqOQzEst/hVOlwPSCXTU0r3LymQYR2aqkAjXl2u/ccd9s85vt8gy2ba/
MLDoPFjwVHcx3VUjKGbLJIikk+hy+GsDkhuZOkfMfo3j72Ezd1cJvu6ozg6AnNw6
WCVIEpLl4wpkWJqPV6+T9lCVZAgixfvpb5aOg+QjkLJtOe7A/yp3SX9+8EUkBd8l
a4CbJbET1taPfctUPyNUUw==
`protect END_PROTECTED
