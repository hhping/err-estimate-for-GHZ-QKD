`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N1nqgiCJ3+gzkEh7IlSFRoKfE7TaT9Jk2Qb06eRDv6tcODUKjqm2/toq26UCWzYE
kwyTh2CicgEhDiQTdYf3LQ4yLXIK+a7hiPdkBNBqYNK6PRYH/C4K6czLxyqtXPc+
9qjyP9OBrRCrAWJSYa1hTHGZL0NSgckTBVZ7Z3CFlzLxFxj2GzuCc9n235kNLHgp
C7NC+qXLSe7c/kJuLjPeQ95rRwEEXaW0p5OdgucspCY1LvNJAOVT+hWWOqMbkPtr
5XJiyNkPps8Mi1MNAgDTWy0U4nDWRhNlOTHxFt2BHNnn/FLx4g55AnZxUoCtk7tP
5tEjXAnyLDGrfM7yTTMNN+ftNmgPKnaOTC0bempKCteZaBY0ko6kZyIs0fbpcVa3
FjGzdp5nOZ5QQtUXyymzqHGmMc9NLGI5yovYoDcDbJKCRNCM+ehy1LFpe41sEfmI
dGTfel13d83jT6OwxQiRwMg4pSoXgf3j4SITykkgdwAgL3Lb6TsWU5aj//9K/TOA
/4Esg3kK68gCa6OGDaWfCyoiLHBo3AmkrIDtEf6jwtw7y6OihsJi+6GNfQz35pAS
xOGYUmipyXAn30CCNwI2CNpFbCf4+9ueeXVvqrW5pxQ=
`protect END_PROTECTED
