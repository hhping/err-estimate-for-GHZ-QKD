`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lF/SkMFlpa/ayT3VdhFmDELRVoXdpBFnEhYrSGVIqX7elO315YqVthY8D2e0ad05
s0S6eMuFN2BXcsYLFI/+8ol+fwJsTk3a9b7l+QZXEj6cXmPZ17KK1mU1Fe9PeDFv
CqOeolOtH0pW2uqoXttfL7J2aOo/f8rMXnGRdvYuW8VI8Nb/XfzS/MzFXgYOm0TC
YzazF7URYjIaxJ8OnizVHwGP8L6JUNKIQpcF4tBNGcEEwakDo/zLSgazLctpgkYj
AxGj/5b0Cu1HZZmxu8PcypOtFRKOhtHZGDdSxljFAHNEKm8lkoAJ4eq45UhZ5bIy
CyjdQCvDBjJZ1eReGGTeyIwPjNE8RPlKIT3ttP9rjuA7eUMLuUxexSvtCSQUEu/R
2G/8SQmkTSzfCRo3BKJNrl6HU9Lwl2+KewtX2Yv+1Wo=
`protect END_PROTECTED
