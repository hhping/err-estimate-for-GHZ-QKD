`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oHfP5LhX3D1Ekq2zQfv2BMxgi4JMw2ahDoHWPss6epRAUe4sd9W6V1c3HYdXH3Es
7CkYQ36Tl7kluijxk1WgVmLzg86kqXQrnsmv0w1t3D1HkrR9L+yRBd31uprj45Z+
oUJKJd0/k+txOnIkL9QUlglKm34tKLg/Iv2HtbimC7p/rKFEHAHn3N/qfjS9fL2w
2Xkca4d5tWkAfNPym+SqulAbhWvwGpl6EG4u3RwovkTKdHH0lqiqYnGnUoGpVrXn
ATGI9tJqmbuBFLHpLEeClovVfibnqzUxlI4QpXoEXxBrGEc5IRbPVUSOBD+M732x
ymgo2QyIARFzK4j5+d7k/qnGJ5CDoa5fXWSM2hO23oZEIm1i0cs/hqnWS0m2X6/S
bCkzsg3LQxoAIjEky88aNOklaZkLyVcLaL0p79GQaQ42eYTNHnYad50EOiP3RR1u
1JOIiw3KKa2vUAaPPnSiG7+1KTW1wmaZ1IY3O+/d2Yhrby/2Z20s+e9UjJ4hBqpT
pS8YmSGpZcCColThdhh/aMragotBfW16pBi9qQDnmOuQhIXd5DX+Nm9v5/lwJmku
sIK+ib4PbOCABTcGyZEo9LfvkOhmKSXsqPjZitL53sc85TZIwHsNWub4I0i0aKRW
giMLodTfqN3DtxCURJdWtjyeL45NDWy3Ql/W6DtV4v6aA6tH7HoKEIixmQ/lS2j2
t+PJorxZ9VLhZ5AoqNpKmwbeZimG9XCSlJ+KYpqpyb/fy3jgYt6MpdlUhzf1OsB6
DJGMeOzNNL97nfkhY6ZoNTTqJcxkM+n7ahoVo3gADuNTY36OU9xFiUtZPjS4Ttr2
fWusRLAt7yKMY8RV0kfpoJPxEZISK6MdUR+YKTsQ2WPDVoev3vHEVnup+JficHLE
Qe8KJespcfDRlre5JSQtFLx7jhA/o4g5ZAAuUYv+XkFE7cUXBcEdmk6IseRsrYaJ
F4dLtjmGBXeL+QWF0GPot2XDG65w1hh6OSqlsHrYY06Y9mfw+/SLvxVsSkujSYDa
P+pUDzvvUWTu8/6gsMKJIw81HHsmni8+L1OSWmXLU9ek7rZEKRN7POqwVSoJOPFC
tZGRBvVgQi9UOr3gX+wDwhgHn7jnJhmUbTmnG4nLL+1QGNZ6zNAlL2IAay4SYZ/F
p4S6jfj+WuxqZYZ9oPLTvnGmWFQ0uYCdmLpi6gKdnn7hwRSXEH3j1WKc5b8hH17y
H6yLRXij/QS09Kel+C/z78W6OkyWLe9P7EX73tN55oviYWEc0MfPYch+5O/fuSP3
WKfwkGy2yuA7JNZCWaHOpFKRs7FYzoabpUTdRzBj0fe8x6Fi8UqdXlGWcAtOLqv2
lMQGk5TYwKHGVMpyXKFJxs2VM2K04kDhFlDOdKYVZT1zgDxpkr3Viru9PBmosQ7X
8q4Z3ieThcK724mOE5jbKdUc/CNUUooXvCN08Dz/7wrMBH5uAHTf+X8UpT2IKzcl
XK+OQwe3dP0sKtANAsh2W7QuoWu6+FKNYCDScpoLDzqCTj1elnWSDy06rvFJPNQH
wQcsIz6XrhxrFiVI91ACA6ZgJZwXH4Q7gPvsDHzGIeNxz/WebBKUokvWYKeL7tbA
gtXVGxIVaC08oCOAZTtOTnABXuvH/cMxSDwdPeRViF4Yc2p62r4NdxLUb819YAtV
/pEwJvMzmbpxdLcGYrxa41ZfipKUpBS0NrcUR59nvNZyGIEGORpKBaBpO83k8XcB
4Qw8AYMyYooc8Dh/NsYvsCuDOsxkQvjfgmGhO+k7dgp0HnH0yJouMv6W+sf55WAJ
nRif5CV7v4JWWcFmgCRmOYFEOm4IfukUYlYYIhMSdwlg+gDZ99oVWmEjBEt6hU2h
fv8KIJF5SNsY3muJu4wj/rzY2GtRQYFJXmvpvhzWmWldL1rwlFnq+NkQjFzMflLn
`protect END_PROTECTED
