`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
odDa28tu7X/vUPZCx5l9y6Wq2M8imD5Kpl9YJFypATv+CwKBg7Ounld6qccSAtP9
7gGSVbxX8k+hZMtKIMZsLux0lyaeIUVxuNiflwXB95IJLoPt/8XgP2Q2U0uPHv0S
hXwhWumDh3lVIaZSaRFfWUDlic3H59sRd1pVk1enAFRvEs1Zm6msyCgkn5rnA5TT
znNkorXupCHMQ4VTHcYwlZJ/usmRduXY8PPzyfrFlD3XR4ruTUb1zOCgAeWhNg7m
AHN03q6jB741uc4nQfq95BmRB8lA0kT8+54+pzGO10faTO1gnwCH7fwvjxTvXidk
cTs+ve15CEfwa1WVEABskVZgXrJYkQguw2QTIRdB1HGI6OELB5ccoYt/MGmmOF4M
UW/dqMJ9ltmdqow9NPBFonkg1awOjbDVfhACJb0yDRK27rCyQrwQaDjt8zi4OMVt
5FP87TZxZr6AU6uFjUtnGKYcyaSlX9mh3BPdeAUotQ8slYhCmdz/t1pVzrJqer22
HJbljmsG4iF1VzY75xypFreU7d//0vTq+m1qtzFsfxhKn6UNftTkHWp3qqkPisXT
W6fFkGcPLteofXdBH/7rKGINuqcxdCQ1vVTGi75qFwMLfHaVU9yVgU9vT9kIe+o6
5PK3oxlzHRsogYdcVLnuLUGM08bLtHC9vwrGsdoYSnz0esJrAAAKkJ3NqLQuEYLm
cA1CXHjtven2U5RGdfG/fZ4PtqkAv+/BHdjUUG0UCJ77UtCqigALfWmP099yHSCy
2yarviu/H+TgJGu7MBag86WKWPMnmF4cnCnTz+7yHpeJnIuwKk1OeiSs0117xa/h
OsaK4NgVYbGUz4CJ8QSdZSh3wgGISFMsVJ3sHVS+s2zJkUHX5BpsmdAZZs/6WUkg
OFsCGQwjZm0PyUQa5bbw1Z7ms8iuIxHtBAt/gxKTb05htiPNRaR5sqRhc6BYpXPK
QksTCCGbdbFVpl65upu1uClSIwzak6c6agIk3X964uH8+52fwQijIbVuSIbpN4NH
fEoR8o3Bvcw7p5BG58l4+BJOXmLksCZGSeOkDQZTskgLGNX2xo3wd7XpEZUZb92U
KOQZyTFJ3iMJTUkne4piAg==
`protect END_PROTECTED
