`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3yfbxYfYNGzm2inbDIFejg2reGc1uFxREYxN4362WxUHDzxgVa7m6QcaQPhEG8hs
RUkYsFPG/7pkH67Tx3AwaZ3vthfq5tcH3qa54x0gt+YfJdMDwVe002rvipSQcdOe
r3PX9GSRCekRUTAx1leebm8N5c9tDTZMgC0H4qUXpH7rcqXKHlwco2nf9l5ZAlDY
wwbZO9ZS4acKEVjdBrvnclzzVZW0JO+YwWW3TVDAcEEK0C/oJqlsxFLnGAS59RdN
fxaeagGHQN5ZVQb48qP4aKJarEvMD+Vgy9L3BK90nl4ynIoFa9gxQQhFLP/4EapK
kh5zcTa8O2taaEoZh+G6cTM5x2BT5qatfJiE0Wt9VMfgEGXcPg54ee4MgpSz5P8N
VnoqEnPEzsIKf6FCxN/7xCxLliJtbutsVUbeQmcMl4g+E2HsyySCIo43LboVXu6t
NHsTjXWE0/y70lnctDWJJVyGSTrdDbI9zX3VEj8jHAonIX7hpvnrruHzLIaDb6bs
8FGtUUkB54RXi6JgnkxxSkXzsCe32ahYfQku6OHmmKAtzUX3roowmv8zsPyRva8V
hBoMUPpno7Q5raKek5pK048chj9K/pTwHMFXR9F3q/w1Xa0bbBUB9SeLoJUMGoN4
h/tQTenfwfftghQEKqUXuj7WcAhdzRQ4PEkGlMHXFu+DlhzV/Dt9Ir94eIJ0rqgv
bXwpqnarq4MQ5dPOnfD6qPNkzlL1+giHnqgVb2rRH9sCbmFG4GMJtmJShtMcx6Vt
+IEcDlRpu2WyiOWkHrINr4lhdIuciVcVjKzcan9T0tYWPU0aORV3yQAiYyrsiy/M
bC9fbDk9w0PSMg3yKi/CTRmZ4qRlE4jJ2bN0BIvWVdgff90j2N7FxYAYMeW6mlmc
4m57q8g8PO1o/HmEDWSgGN5oKVGM/AjmnKPGQ7b77ASK/hbrKNHI3fgDHpg/f73R
UTs8UGNFCckC8aMrgGrcQuBfYQZNgU8G71jlgkjZBYXnSlQZQ/lv9+9VnlJc/9al
80+bKSf0+bS3jGcsfoidlORj5fHTTYAUaGZfYJqx9Ro3N5SBzA1SHXB3QKo81g3W
BcKvrHNj9g3Osgmo3Hd8nU/Y/RT9ho7GmVMFIMznjzzyxunxu6d7RFF0nYVDiHMZ
3bulCuD6pnZwbMrlXi39EWfULd05f4MjcfSMAdb1CjHB16Rcq1SqWSDbc3AJXt+M
NeCavvzSmxfMdJev6TSjMlnSSEvMC0/QeMQycFjlkXjLi8bdnNlWyq9nidVcPJgr
EePzveUyw5lrnkfi6ZJ4mAGq/agAiGE8ayZvaGqb5jYVblTROjZ4FY36ggMChkD7
wIPGQqLzIW01yB+SNkv9M8DrUOxenK79T1y7k0bi2LuB5rNTlUl+XFOkH0CStPed
+ymKWj0r+I0QujZ40+4dvenvIFXJ1mkHOGUMAT0JhqzJ8zIT9Ro2S993TrEqYLNW
NJgQbLmXxyJI44MtW6fyWcOPFBlqzjmicOyBOZxoEK+kWEj6LtjlJy6QvZXMQiL2
ejrTBLxoKU2XtJMP6rYj7T8Fza2ioQYpiEDeDtUZLF4Fn7IVe2HsfwUa1fk/CDy2
C7DgCjfZVX6N8Z59pt1YbMwQyuASzcfCT5WlV+ynSGWA4AfmnFNz58G/mmlUt1fl
TpATetf3jepYDMkkZlbbw1ubeL0cU10qbCIpAEK+lPwECfT3UnZSMRjCcE9QcsnL
mOrCbU+aAftzt94nt2vXqm6TcNX6DU7lGzmqNrLhzu/pHOjxBco8VE5D++2FUErQ
CyY7+rjfzko1qvoxLk2hmaF9z6aPPKAi34wpj9Zvik9cX6sWLSaaaXvSuHMPXUpO
qkA67v/dM5bhupcuT+G20qsrOr7sfbF2XbjumsPi15p5IruLNwn6xZ24zGdP6DPR
tG5EQgClJPIii05MH+ZMLZ5gWTvrCH7cYvJZHT4LTzWqJwbeaVJ71xm1pBcBSO+T
L2zoLnbbWVmRWwkQtC7qxwXKpkI7ob3MbQ5/z3NF591UDHizG+p09XCpKrU8qS2/
xpMdhVWGUMno9NsBKebNu7oQFdjDUjJ1nrr4J5bCFjgGSRMIllkvYaIjFGSsBkAx
hWzmYSmpcUHQ6h+C08Dd5TlQ5XlTNK5UCoYw2W68mWyK1I8THhm50dH8sDhuaFTu
a36D1oVMmoPDWnmMy+aAztNcrey2F5onxebtTcg42CaCVMkWge11/kX18lKL+YeT
AII3fOMTSwLJrXDwRyVhKEVBbCea++jlcDevjhzREAZ0Hqys/QvG7Lo2BC7q4TXM
hZ/X0wN/qnVPy3Yv08EEKwnUwD/DHfUctdeEKSR2W1HOjat42GGJARsu9uuYXS8v
qXSWZZ4KiU/FqqPB4YUZB7fcqZiS99KK+Q+mr7P/r7HyztfFbGakFF9O3O4+3NKM
pqu6Yf9EexjsrjEBmjslNepP3IpXGAQ/gCmktsW55IUBhxStxgvh2pK0yD845I7P
cLpmzYhJYdrcRPCGl35sRGg6xbbtVHeG0ObOhsjWvuI1hLrkXuBiIN+ur7jzXsjT
Av+p6lKAoD6vwLzpeaw5d/H5aZV496imVS1o+kY0ZaXqmz0hkgJoyHb3/Hny3duh
jfXAtRQouPmpgqVosIyiH2hGaUAQvq6sW478KMDXVETLyAHD/ES4oQOI0rZ4T9ER
aRx790++hN5esK4KpBTPrzTPRdEDIowGWyqTL0A7ZOzXPmEx1zdXR7bNH1mpfdEK
++LCxGBY0gqS6dAX5oX70WRFDgGHk/gOyLt2Vb/c20kb6xqxQR3Nd5ekdtiGjnUn
RM2z+3ypW7t8lRCnaggQaoVNaaWZoeScR8hszJrhoNIscv7kD4CmaUiXeA0mwxow
eWDfp720EdxMxbVAhWnaulhDvxqRmd9qHSFto0w8oFti645eb8+AcJku1zBTew/l
b6W7b8LEWt/Gy66M09NycJVZBxURL3CL7SJKUSomf7UPlEwyxvZI6qeDn/WFtZ1H
MciG8lkVBV4Phr0JRbYMgXg68xnO5LbaExqtDZgCYfFQXnbITGumeLdeg2mvNQKh
Tiy8fzxFRv3nqP4ZBz2WA9UAet5VIh9JpTbixf9v7YIeBJ8ZvUoPQluASI1sV+aR
6g0n0bxkeAIRBN8CrkBVHsfPKpvVrfEq9rpwKfdQtr1st/iYuF+gRNz9SXOiSwvP
J01VuZ0SUU1Q33cab2Z7c2Wn85q6qxmh0WjoIduOQ6niZSJ0uQCZ0/cUMiUpxn8+
t1JmKK3Epo6NsuAAiElObXJiuE9bzQ9eEFfN1u5nO2iGb0JUQwBkRHGTrQ+AEUwA
TQGREfWWpEjI5ubPjrjSDDi8jsVo7yRmwADJdtVjSquAJgBbmSiD5T6IGXDVNH/m
L/aapn15GrGR546Pe+BsgSKiLpW1xIaWIc7tcqjaYSltES1rCYQb0l9WmSghYCm4
Ujdar22ClIhA8PSN1fr0QJttn+BoIarJ5KAMbLYXFnp0wuvBdXmgXEZ+dwoQkbKL
/rJwBnd4uPp0yWjVguNvfkBYbQAE+kiP5JC+Pui4qgNt/5Li6eRthE8/Id/1QPsD
HmQJwE4naE3eL0+hbq5ohTJHAx3rMpau6WXifMJBdPzk3kHeXuqy9pjHa4WMwXIT
DYvLgdNkblK8xPOAmzwL4YzWQy1nzESefgCrmoN4meSsvf2H5O/wRXfTMLw1Lnul
eUt7UEDbJw5cxxL0sRd+EEVhrSu/YBNkN3rJU6hAtxO49lhXY5V2Ji+8imy1QeDL
ympdQqEKCIxhLd/3kl2tCMecZW3ds8c0DSROYV5DM0vLaSyg/iJ+4aK7UcsKG1s3
g5PS/wlZYCC+uKzHfRh6dooOBUzYHbD2lPui5FHKcilHzXYYoUmlcry5ecSE5KCd
YxuWEUt/ZZHImZh1h3pHRtn0ecmJpWl2Pa9xUM/nLLopdS2yMbgoEBVh6ywYBme3
JZdkOPN1TK+sgLSdCasDqL4qmzBYYxAqv33fOWICqxpuld5GV58rA2gltuSy0+bq
u2ejA112NB42RLuhrjCtWPNUkv27kfx8IJHlO725vykCB1104ENH3ZBIG95hh3f6
TAlMzC0MUyPi5s9xmqRwoKJy6ajmV20qk+rp+YcmZpUhXCdcarlZkpGXWOC7qatz
Ofoy3WBWgPux44oDAsCxASVcS0uee5OyV8gB7OExxE8CxxqWzTjKMYK7K0IR8tjZ
aXnkTX0fiL1JBCzsPkxbwy8t95GLpu0bD2/XLMPxbGX9bK0pdGlp5HYydTxJhV1C
hT2RM6sOyQmWoG/kBzNMk1F4vhyvgPx9gNGhhy6hlq25KHRPludpJ8E4GrCcmk5h
IKREjtjiDuy708NtjH9OX8+ki63DJ/HGobj/7xK7y4bODGmv/bOV2TJ4mYbBeQSK
exg3AwWp/DPuMjuEN5CMoLCn+T0zH+rEz6IJgy/ek0GDqD6b54FH9LfgGfQgIJyU
BFVfFjUyF6lsg0pxj/ZBkVD0tIpcAf/3ugdvSumwg7X69YiDSMEwaGiubVGb9plj
eSJr7CX6aZdZeiG1lGoUjDYqiM+JM3QqjeCC1fMlMK0rk4dZl6Uvy1gvvwecmJ3U
KER9I4ueHRLKGL7uEoVXZRDIJ6AKRYnJZ0NAoRA4SQTS0i2QWskh0sRRm5GJZy/e
2wl77QZ7fgrRpJT4zphVUmqDr9jdw2+kyJoaZuz4iTcJmjG7qnr3763HHuYEjfg8
Js8kXb5HhofqRbC3tbcPQAhSEZru0UDNw3EcY1krf+J51aoCGX8ZiaE7qgIufbLi
T8mMZGI276D9W18esHVsDTC8IhRV30Rt2LOwwvbVMCk4iC5xWHTyohcWrNGkeDkL
2s4OM0yQUyZIOhWNHm3MfnOj9odE+IZKS0Hpqrr9cIq48Dc5JVrYVXPEq60ZrmQ9
lgedXk5/kTVqY0JhLZmEZeNY+0ATk1SltGdz+rfpuJvZTepAYWbLekPu5WTYYWH/
7mqiBWCbdIqbBxzaG95q6R4oXmJaENfmyU+tNLzoWKs9/0O4oCWED30SMz89P2G0
ngKgDYjlxw6xAONLC+3fZyCcPmatzU4OOpwBgNoJLXZvEd/RTnKCYWN7beqnlHTY
eAmkbPcNUIHIcva9oxVjXNbR3D8zxQZwZ9LoNc9XhcCjKJl8v/2fGGOhmHwktZ78
erccw0WHJZFMwEKQgqwSJtfdcI9J6k6L6k/4Y6t7+iyPzrgPPzS5RkE+tTkcP9xH
yEnHLkIQsDeiBwdRuNB2kAQ5P4QEjPP4v5+vyiAuaBhmdWNsXhoAPC59y1E7gl2U
nebcBM4NqtJ4F1+tSoqqjJ88rOeEKCpW5nMMpLAepE1wJXC5WiFcYOOrrpg2xWWe
MH9xVhZyol7zfT0IgmQMWT55i0XZnqDOuy923LildOymgqdAVxVhWEifNAQ9YSfg
PMup0+pmqVrV4ZAiPez2/X10IUyEJtP1GPDLB8/2b6EDtJElDqYEucrJD1T/WNFn
oLYaIPmUk2iyHiK6hlvN9HB3V2BiCbc07xpEVmLhZGf8zBm0JK+CUDfve4/y21wm
M+ssaw5yeEQTTHOauJ+I/rocXCixCa44S64x+tEkCMsYnQWJgamCnvhGYkls+DAa
IJr2Myq6xPV8UAkLUemPPalNrFw0MkV5YNazsERq2FgY+LYIzpVz/Zof8rPbG3XG
qDXDPlznvYk1q4sfOPDySTq92URb4g8a/lurhfzuaHPu5VVjGbzNAAZ6wsGRp82c
/e9p3JFE2YTk8RLRQO1rMycPSQldmMF4eYpeaCvBRwXqG/9njw/fcLOmWc/L4irK
XyqDJt7E3819ixRs/9N5rNqgrbpd7MXa3c2vDZ91iHXKfDTRe+iJQyOAVyUQ+qFn
DB1DkjO1SyFUCrrrZfubidNlegWr6wIrCoDcjN3Qm8d9bUpTtyg5Rf3ID4BisYks
MCHstgBjkBIuu9iqRegcpDOasc6Wcg5aEirJkaECuq7ZCace2JtrhRWZR8GsnIQe
xQqHIII/qY5dghr3m3g3TLVcqM4aRZJOmOj7a7pf0/kElhZIpTQtXOYv60VQQ7GN
c/CriGvGB5R7kPOtSLgiug==
`protect END_PROTECTED
