`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NCmSg8zdGLVpIzkY9/FDINFgyL/B7kbhV5JQcw2FiubA3JRqhr5xeCQ8fc0Fg5Au
rfAA0LQiJnQ+i25uSat39t7uH/aPQPJcbZpSzfXDLIao96C9NoESlYtAB2a0NQqB
D+1EVrghZfFD/T3aRQDcX2KvkC1srl8eccDcFax+IlKmQ7klkElVwMmTZmwvcTH6
a8rgedegIMW0JHYwSzbN72rlXG21hRMEkXbQxmp1CG5v/SzwXX+9HFajieaeth0W
Fy0OtcFXS0qyI60yfB0k0CE4sXrub5gLOhWXpOSVUWeuZjNzvQk5X3Eh3nFYKPK5
Mt53kVmnVx4NYg9kVa0QJas4WR1fxCZEifam7CxKQRMqz0kZOCv8eEE1OQasJvrQ
qVfbmZEfqLSbbxST4Q2iyTG46HKHqhIxEl7EGTqxcrVLfG9T8z6aUzUjBveKCdxL
ZJjwi+R8IXm9ce77gZOViPXpwKL68gXzVcrMtG7hui9RvGwhaNnNve9kPYdBuQPp
pKHFK6OZrNvltZBaKfV9ilW3MtRlQBx3FEp1Ml/1fDlqDXeaimPt+TIW0918NDbC
uvB3gZDKm+B/y1AKPgp39ZqdicWUHk2z/uwXtptYGzKgO2kuKSMsuIlmcIUHC3g4
CA1u7+1XxxTWbvvS80m2gHrMQEMAOntkn0jVF16ARmeZIfOG12Z7FNuSbCvoKjSq
Ixt2RHy64g1dGxF61t8H4fV9ll9pBxSUBIIJC2a2Z7Sb67947deJgxmm9ouOPZHw
l5DL9/Ctcs5kYqIyGctfezH6Lrs/6sMso2WkeknbhA1q74hFlz2ZjKpcqIdP/ahn
2LUqxMtibV4LkcsK7aONNN1LPKw8uNkL54I6Voqi1nb72F7Cnibpais5wzt+dJbz
zFXpXhjykctJ6li5DFZLgcfsljpTHUk1iYXDLuN4NvCRscK0f7aDigOM80HOsNVH
PKbI0Wvqy6yxHnpVUjAmKei7s59HdqySvQWYYjCM3K+htLkSoYLcK6nSkUUSpqGC
zWAFFIqgIxQtOJWeGmeTKebhlu8cVpMxxNabMZDms2C80/SBBzKpH64ViOBuXQ6a
`protect END_PROTECTED
