`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TKt7zveGDXFkcSEfwnloTiJ42o8Ks4c2nMlA7MFA1o2DajDgV77BiNLHvN5GvKna
jbzWgOH2urSKidUS3wRbn7YgVsYP1dfnx31X/puSJr8xrQIKDi+UlyMzma+Ak2MU
+6aXsr9iEowK3fkyH4HIlUdXUVQYbEj9Rp/Iun2UPWaM3clkKfGP+caynRcx2zIk
bNBX18LG5gEG7uMP9N8CJs//RrgN7sJsF1E1qhHRuGofHy6+oJrSvwnvLfKUpgK+
3uWqXikBVZoVqX4D1677fn10RYywPTPHtzJdj4vhDTB5M453wDLPJhyRAf1q7JNt
sVwqf9XA+e0glXbGusrBo8I9R1hVboVncY+5MHa9VDGGC+qd3BZJReB2BQMRzAZK
LAU7YJ898e2zaDAq0Cpaq5eyRm3fxyqpMupiX4M7uY2SEU/CZcz6gD1B6BtxLFrz
1/3qcv5GAsJeWBJtx/rDprjWc1f3CI9RWaJXorMnIOgpt2wwXYcy8yRPaQUQMGhO
Mn9oxNpri6fadD6uRd6kNa3SRqlXlVKiGBBWsZJUm3ve8fizWRDSbZhGQy3UjhPi
HevJcs3/QG1V0K6RGHWUyE0owz1NM+eYrnYkRcJ8VNa3BbaKkHp95ttSIdGVp5Hb
qu2/k5+u8+lyBclx+VymjbV3LQErLgwuReEnEJvKIWYvc2y/PUaFoI42Eaaqh6Sq
9Ep2JuRdJZ8Sr7SB1orQh9ef2y4JSDQ/fHQcxHXp0bcJlvdvLYegFgusKMDOCfzS
meYSkX2RTIg7syzHYw1sHk0C2YUQYjVL6JKJGeYknJFianZpuQZLGmnnrusdmV4B
hszT8UzlrT5f6xfeh5IbPSExwDOkulDxXSiFKc9fPK4bxMtCq1spVSwBiPYhnEsh
xguK7pG1EzOp0kt1KvaJczytmUN+Lw4XjvXFVx/b2U4jZXAO7imgHnkYfMbWlxir
N038LErs18r395X2CiQGHDe4ryhYhgwnVRALROgpuJq6J64xtwgthMKnKA3gsGIF
Opw49wkrXyAjhLAeTWT+TwO+k4S19Kn2XaS9rfkH2MDCZaxqfLdEz7o+iQk4gtzT
NG3t6H0Andn61e9F/LfpbhoBFDTAsw1x8dCigOPuJLZ2nmAQI1VEuZr+IbhkSrGW
siZ8u5NyszQov4n3N6fvN4McSdM+S/r3vIqzrrmtrQxo07beakU65XPK7HPDJsNW
bzXEQpClVJbPqIxy1urw+86A0wiM74gk19vGNun6Ix8ISEIlc7UYmgRQePVnmu5j
jAYtCap7FY2s8J7u95Mp6JGNb7MjqRQthOKv8ftCEF8ble7ywSxS1KGTp74DSNkk
WWeKdE/eSu0d92vLbe5lsNNXzwGbIPt+zOdPnUQ76vh+N4uaY8Mh6NYHWvOMv5ET
XO0ngAiShTnVXKmjjadzg5uZQzFwCFOnp8MUukJh30wUPCl31xtcrmdNruFoLyBA
AmCz0m1ixskZEINC027c2dXBhL8zNep9GMqApAxnBB7i5TmEpzr3BTCCc4NUhl6a
IdDa8Lb36Vx9EO0Mz8q+INRs/rC6C09xW/JBAY77i66Tv1tDzlwjBBhGHPspJmv/
24j2JD5FbwbkvzsBrhzBZo7E096rKGyuwtTQSLxTK6eUztDxnZBngvgfeMVmxsic
7RZXyZT5PvLc/xXKXOz1qaGFT5ZZeP/lziepO1Se2wLiM+bef/pTcB4Y7caUPJGK
md5Js5o5eJlGLTUhXT03/j5mQ81AUens0ZB47Fh3qajL/tEO7mAIjRBHq1zLZnO0
zo/H/8YcaSHpzdhZuS24dCy2mPbn6BDLCQMJqD5rm0olFl+kQjRl9lbnc/KWQ5R8
G/QtN8go6cnclUMMlRqR6sUjqOjBQzpuQPNyZ3r7Z+XTX27OR4wGbplsU+oSgVA9
qCg/GFuBSL7ZELR2PJKbtAy1I6eOnXhVNADgzAoKNUv4hbhwfZdVa+HVPeVe13fn
mdm2h4QvqoaziG1tPQjpnLKPnrNl0J93kWfTmO6rUc7wiT7ZONS32mTvJWt3Z9An
BfyqOKXfZC9Sabfn0OoBqrNjeI36uM3/64K3jbgG9wSHFlVjXpKm0MMfxNjA8XCZ
xznkpkNHuDij7Fx0zT834nHABhY3yKl3PK954SzU8aUfyMKdjh5jm60MyIBI+8On
JJfv2kOfLIo7f4FkjMVxKW3bUuBrWUw5qzCyOUpEisk=
`protect END_PROTECTED
