`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wCojYUYAKKgHj18/+qXYEkkehBtiyN8AH0LpLODdvO/2Tw68nwk+OFGqpJWyx080
qZRyqR+RNHe6/xEKiuKya8vweKsazIg9sffP/oSNvM6byH5sNuPMWrrGWdz0/iaF
8AFRKWUwRL2lEAlt0laWKCrJ+veskrvsFHavPE6SWVWXWNf5PaCZO6vCvHUtgdrl
d1vX7Qf7FhlbiRPtFOys8W+dIMxpvZMR9b5DNK7iNK6U/N1g0SZ0ZJCz5iUqPdUr
m26vX1vxFjbwLyaq0GRj/h0frxR4XiusmXCcksII4dE5Rh19UUee6FirzXLunea2
JNty8IJcEXvVuGu2o+/8XQ8rAQXZol5y1aS/qHDDNPHKj2PLN+6SLCDWpKbrw26i
FirldSOb25FnJovdZzqMQC2b0aB80jxeXMcnJiiNbbar2uKiyxie9sf9eGxUnSjU
rNbW0rGsAs26T2SMGe9dqel7JjRgZh4h01nFxs/3U3sxgGGKGsGL3wuh8zBuNVVZ
R0+1QE3hJlOwxQDgchLJj27/5VDzUBAxKCJwZ8VPbEgNOdfnpui1cHqX+vlEwzfM
TJNiTQPgiXYV1WgV5eAuGAe5PYNSYCxGa18GhAmvbinjB4/LULfp2g8BzFvuCYww
EIE5FJdhcYw9mj/mJgW/APOljSnd2eLd7rbHhBUfCJl78bCEtpr80jwzw4Y+pmfI
`protect END_PROTECTED
