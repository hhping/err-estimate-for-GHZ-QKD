`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B3cFDjUWBXATfK6oiMCzLNAxqsY1baD5dEVTG3jPoDJKbp3C2LQM8FlARCi8pwAv
C1gZaHif0YzNXXxv+kh3enUwFR/6xC110LKzwSIasOn00hmobWgud51NPWUJVjvB
ODVVLK7Ut4JW2Z7bFrvDChYeKjLjpNzPt4GuBCyRn1vtN5SQWCEDPC+LWupSPivS
r3DEO79GTGaWBsfdAyRUaBRcbIhzAxVKNPBLY0CjvHAJOiljbJynWNpblYOIBpIi
eaf0K7IJfgom6fGZEs0r9hwhOLmfUJ9fWm10layX9SnG33iEKXQLj3Rwca5UpxoE
PU371Cbsoi3BTyOCMl0OnrXeQnXo8gWF3NJMFy5C3DcW590hhO6SYGS1ga2JeXC6
IGtSSbOHrFJAcJqvQf9fYK6Kx3M6z2baMyJsFnJoZztQrxLouwKAytTfOmL3RBaq
FJtotZnR/YS4a2nuN67u4qlIXzGGI13QM9cWK8heBzusz2vrggtUibmjd/vZ/+sE
Khfd6GEl8+W34nfMmK0tP7TSEZnIe6ish7IKY2FY5vtOH+MlMtUgWqf3/vC1aFxb
+u7LVdeY6UVewny+MQqbmX6j8mQZSZ7voPWfkCNrtdIQsTjAI96jWCUwBGEz1Zp2
muBm5A5f8M/3DEiNPY/aolGXrQleqaJ0b85+jSk2yAZBdeMvtzLrrpP/Wcqvc1eT
0RNXCLiaqWjVRcrR6dNmp7oixZAaJImljnajbFddwZ6w333kUIgwBX11zmcNUbPH
UMinBIJJW3dec9E0G0rG0ULrCgWM8V3N3YLf7hR1pFbmt0nz+vlhCLytWrnke/ib
KSYjk5TR58sToHgmwKvOqPVnFz51ZErmhEI3ihnApJ2WC6EoaWjQ8SCmmUjxcDYQ
Tdn4eBHkgMi/rSYvH8MG4kECfRICKIMwonEQvvA69plezHo0HmYZAFybactjbJnw
e1vav4n8V5V4wtZCa4s5P8dJzFSn7sTQtINpmj+zNAZ3xPLgbt4z+6as0r/DNceg
/jx8jSp1ITpWxbBQO8i0f5065Vg89LSaILzokHxgD0eN85CdH+f82x3zeuk02DUw
EALKlzCDMDIRLIkOHRZoHG6yG8+8JgBhEqiI1CQAQfWYZTm6HVGbNRwiQGB9xjbw
H3Cro2SDU8xowdac5zWpovnqzhlybT5eMkcVuEe1eQc=
`protect END_PROTECTED
