`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Fn4vmIeM8GNexZcDjO3/EYpopeyuzl9OKwgAQcYRCV6jRbNhsSLIrnX81TGNT9z
nf8eQAzPOnu24xyQiRJcplM+b74yiom4N7VDMqr4SAI4Vz8BbIeGR0jClaiszRJC
C2NW4LKZ/0PTSs2GkyDmwuEsMtPIF6khkfgW9lQDOuIIlI5qpiCsOSqYPS1QWJ+x
O7xo9Gde20g1kz9veKyO5AuyKO4qs7Z1h1rCdXA4ptQwCkMy1QBdKD3SDkF72HFu
oSCZqzY8smsqanjUng62b2bXplHcwP5qZCUXpq+ZXrEWZa9DzXvvknOHQIP0tnwR
AEQWN/hF8HG96cIgrlmNSPmyS8lcjptHUQV8LvRDE0n2SAt0+kLThSFG3R/Cuhbg
VuyXoJB0ZC/sHw9/7OomfsZSdtJ48J5TXFXPcObRGaFcc9d8wmNl0ghMQqf94Pis
WnVzgSnTI+BzlFAO2kG2D2OCFcu7oXESc/ibbI5qVDUci1q+BnbSen9PWW4TeH1S
xOaRb6t7qwm0qV9FbWfZ2lze53KXjBHdtGZQKlEwDx342IwckZ/XPVITGA6Kce/V
GsGMxRCRyXOpl4jj7wKhNHzvq/xbPcXc5NIbECLey3nOGSaYjVoLNrRHqatOZsow
3VVhLVTa6MvdDM+hBWlTzRY+nFkdolulPFd+CK4D9ncN1AmG3ViitJEn0Gsbw3pI
ul809fzlcd90gqoqWLVEVHfgDL5zQ8Y1J5/pV8AJG5I2o1LHZW9uAJOltXHPZOaf
s0vMOcHmXoPWZmuQa6+ehvQREdxKAIbypQt7wyK7xedckAQma16MdUf41Opnof8L
3iSbhJDuqc/nRy/QDIp4946kQNRSnIhW6/2s8qMsF/qfL0N890wicIM5CGqsd3Ha
Op5ukrnw1GKWIZr211CdNO06tf2C58R4KgCumdXTPkUVQrWZG71zPKmO7+WLpaTK
g/Mk5F2hp9I8fljsRou00gtbf3bama3XWjbQBz93i/yXaSXkiDpJGSuFcDxR5jLo
657fkCH1ADRqP9J92n2d67MYGX1h+/OaRihSfErmQrdJ37Eaa96TdKDndsVnnety
lbosTyqlOsndHlDbtmiCltvhgx6yhdn4uY7uGr90lqPMjpLOTPuP5uaTEgLRwKx8
+AvFMPqoUSGx4vROcUCacF1WekpkMPWUNhdkgNM6X2gVhjyL20Ghn001LFraHfXb
3sMRlbYQbp7OQwyBKwjkb/NeRbRcleHaIZH2zecRySGqFvOBwlslu+B6tFvWTNUm
IXIJwSwEznlF4upVjxc23kuxsBRDtHmOmlTErYJ04VjltzjJUrDysTrCIcG/tyC+
xJmleV7z1rjY0lkZ+KE04tqodw/jf/0aZyKmvn0KqkyON1O4W2yEq2x2u9GRdHDh
PPhD8hGiQs+Hvq/5ly/Zz5lIx2MjaLvnzwzwKPQAbvm1Xoq2AtQMvj6g3pp2mM86
SJZO0WF2IJDZqFtI1jWtL5XKqCcTmxZm7b02mjuimxapuIx79SRBfzLys4FtSfxa
x6nislt5Njrmsp79lexWawYKH+UQLwqdpb6kfEQ8vAHgva3LZQ91K9r/Kuor2HSD
mtzKDin7njqXhnflmAN5sW6qtpe/L6IZjYSRIxS0SyD5jeU5UDuIXj4oVpgNYjhR
ARBpy2EycEAG4DdWMPLps1hzot4UfgmK1231+b/YMpRAP60/lgZZtmaUlLzpG43v
mH1flyrlLXper9I9JhxTTcc694kiPxFiDDwtEuwW4XIGa8IslOkLdQA2SEl0TIEV
GDE5+C8EK8gU5HSKzWYF+EAk0V2a7uzNsb5CBf8zxbVjaqShk+juXjfeBCg+SVwY
XK8YtZ+OC3vUz0rOjvAxKW5HyR39lo5FoafUgYwNsG3vEhw54SXsdDxhja07/rsK
x7hBhi9JnOtIHzlBUemf9u/MXUhNHsD9Ejk51kmDU8s0qgif++Jxzlk+tN7KBicy
K7NYWD7dJsEv9EG8OSM17s0oD9+YlDsAXqv5t0r1spG6QEn/mXx5FxTua7Y5+YKn
t6YEYaMSgugOrH+EqWWfiNz67A+uVzDB4N4s4haWVcREeHG79SKLXB2FL23oBhi3
S7WV9Lcmynk+LCIvjgdMt/bSca07QpetPZnH75YalZb/AocfSuMgdNM6Pdeq8FJM
fbpy1vEkajt9JgkqIbrTzN5vODzio93NLecVo/fP1Uhlm8fFcn9HBfUy4fobUbxw
lKCslgEAAHsgVkIh88CJXuPw7s5SLFHdtLIkLBodhan1w3JKSbOUgijoj5i3ZMrF
DPjlV3GxfQc5NBKmO2FJxVlujtti7grQLSdqGrOYi0SNUnGCrIJh2hDhh2QdeHg/
g91J1+7bRSiYv3H15M6DwgYU+2aeZDFup6AbCgAZYvN/uAmKR1ewf+3WJgQge4pn
BdPb5h0v/AgeJt1/vsOWatsei6MFishhAZYxmu9/yagTyqC/E3qFPHwis8VvYbs9
2miqwqJ5FF7BLxbaPH5jhb5QR7lGDYRiX+ka6XQ9vLM8TAXwrkeQdLUmxCdaBm2G
nqSOeG8WlmaXmJABXr7Qyw+x1Ev1ZR4HctdCn95IckWiHRKNUpRlcVK0AKukPl6y
9IKky1BiSh+Zu0nf8VAba7EUtkE4gu10b6oqp/q79SjiQiIMT/rMqRqEKyUk87LG
jebux5tPlI9vSfygZnGKJ/C8Z03mw33EwRYOajyUNCpY5XeP/yGr1xwLaUOEPQBT
JF4NAN6jUMeWxksPTK+nIU7WULXc4P/zIKANqrjteo9R4Bktr1HvWgQquxr7+ZiD
P430C8mzIGgiNWF7tKXWRv+yDfwsDooMMV5AzPATLYRLsELznCABXHXFNpTymi95
FCKpnIoJVwPeMVjpPUZ4tNe9Y/5uWsxzyM1p2PufbocQeXzdhzyGbyi5lIMcJzet
QSiwcDWdlCmzAfDNXX64NPkF3Bct8Yf4oG+uJvOpq9r/GKBNYoaYmJknNw+dM4we
y+7zBswGxLOHAu/eT/ecMhx0Udv8RQ0PIpbcBBXICRPU1ypU0WiDliZob1BDpsee
H82w8/kk+CL0crgtHhU78d8z4gYujMFVqbFvupVzFAGy6N9WU/+L+5lRj0IOSXSM
ONpCacmMupcRS6g8KygeKk2ViP/TDofmAWE6r8g8UAAckK6DiOFEDs26w2zfpUri
JWZQC0bM0yhFRxjA9PpaExmRxhXskVVnfmNZ/uGXbGjeTELZkPw3KoWfxBCpXUEc
4tQoYOiBbIyQRvIRUqYXhGKpvlNrQ+lpkF8IU8JGeeNJ8kpTDVG3ZyclKOpDLKkQ
X1BQp353x/MgNPKjacWcU1qx+/5hQSQsUkJDa2zDdLy/PPG3PoFCPxeFsSk7cHx5
U+OQD4C+JIRMnYdmuWAOfQZfCkX9wssBfV7JsaCtmq1vPlO4l7y9W2ysq7NEcFhf
egwZFpKaTKiFd4vZGqJ3kt+6BvadESJ2OV3xbeLN6JOP14x7PhKdKC2DwhmMri/c
n//ABDJszW7nBgi7xF4AUTmlsyQ2mp4TA09AI1zv1pmNhIHyFjtB8ReMEf1GY8B2
okxW5LGSVFG8htN6ozApFy3BU07fwD8RoJJ4BbqzPUv+ap2oCHM1IAm2iJMkK2wi
kdtV6xZ5P5j3naeAIdIEBOSMyvJXZbenGbBbyz9kxQlaPYOfcI7ZJ++JVIDnosfE
86pChJBQk2ZDaFbNOHq/AVHwmE+OxeMX5eSp1gzsGGDhKUVPdsI4swkfLiZOMnqC
vQzKjJFIQJ56pmwDPoUc9O0An/AXESyq6NaQIJsP+ysFzh96Igo1/fHeB+M1hbtZ
L/lUczxeu9mJxW9QPu2f+p1Eo+tzBpfIHhtXdYZqevl4tBoZiiN4x3tEVbrmPzUV
dMiDVNI7QwpYnriOJSWTLIsBDxMsmczWgYI5hgWI5flGW2iq88p1K3BQ28yTa/FS
XOCXbbzotf6pfyIZOHSjYC3JSS7/+JOfKFLuyU4scO+rVXGXEKAt8iRcCxthaGKj
TXnEPyZvVEUK52pIAocL3F+1DPiemqt32gC1cjUbLLeXhaLZgmv5c6vnNAy8EruA
HkjB9NIz2F9uK1RQy3UpuXmKv/28RWaeDCK1ZiAjjztRTml3w+tzd4ebsucaUvBl
5cVSOHCufwDvVrlZiLkBigGcaf+X+84UedMxNzMP9zLneNFFq5xzugOlWiJCdtS3
rAvIKZQf2/Ji5oRzY+OW9PsC55Ifc9YQZfAKQoxtjCs10Yp/52Rw6Y2MmUc56tX9
iQ33GACanaYW3RiY6zbCE92U6Sps4MZ1i+TvGM+lzJazW1B9wfzV4mAyUnR17J+a
2L2psphuXE9f+CbOWZ0atcgG/66JhgPsO5YmXj1Z19cvlM8QzFBMxLxdrpQeR1YT
M2WcSY0worgJj1egb7n2AQ1dobwTNivMIB4+a2FDcjPquFyRFFj1wuBDkF8yUw/b
ItIGHufv7dahJw1N9FT/f3fdhreU1sihXYAGB8vMW9hFWDIVq7OOtY2tOT1B4OAy
ubbgKiuT4BGJFi95eiuLhBH+OvhhRTq3fhIQgyv5RzvtpjXY56cTg+a8KgasDynJ
bkc20nbI34qTB7ZnvniXSiPZOfHP2Zcla8kYxnfOSWxfUrz0xeJhYRe6I7POcYx4
WhRG4O9uT/HVGPRvc5myApGXQmMdWMihoQJdMN/5Ptr9NMPJjpGAPXnJntjXQ7XJ
macCIddJFqHZ+kyx88MagBVwcoDj4Nd58c8IUFrQYm2pAgZa1rSazNGftj7qBKKa
1alBfwoTV7fqKJahMlMyw1gGpzE97u0J4OD4eTkbMMCGQzQlXuIbYGsmnvbF0E7N
BrJLu3uaCIsXK+Y2n0NYjZSXJ6bdjzFn4FpRtXVlC6npBSGNsIsZ1hOEd2HZ1Tqp
f+hgoJ/mOfZKlvuHCcmv91dVzpCd6jQ0DrvkJX3s27ojf8zWeJPReI2z9kg/uM3f
28LDLC/eyDXTa94RFHBLTQdv/vNz/gBDd1FB+Wmu4LdwotXrBtaYqJCU9SnPtjH2
eHcyDb3sUnQk+nnb27FXDSbmjes2yzSCX4zeN8GmHxxWZo1/0vaovQldHbDlqigF
TTfQctIhEhuOaQJ5JXfIKaz6kCFJKUjIcEqOo8hUMkqcEkmZBwsdxSpZQkK25+Qy
ZNRcpLOIwA383hVxvcm30RxaFOvjWjgaIFW0Ue7Kfx0koRYuvDoiAsSvO/AG1FaJ
lTUOazxjIvv+rnnPh7/+dT6uUBqavnJuHDZCvxWSUHJeb+xDXpWls5f+OrL25Kkf
oOhkNOvx0qWjNCKOL5tPW7bUPQuSS9jp4TaaJIthi2rkCrbvQI66aHkvmvoFgXHr
bwfhVq2eFljqaAY3ovVdqg86e3m9HpYowI2rJ1P16ZlSQPLdRrUwvZLOyFRRdzeI
FBpyIZnFVPzmDIFvIDTbWZPFgDDwhjPtrryXc73S96iSjwxbX2dpgt/SLtucOClL
SVVgri535nw9gUprnJrMgo2/affCO9IgpG1Oav7khm2xafXqtMid3LSwej6Y/pHR
ge7ZAt3tRd6jtl+NhqDZRRbCVwNK0biLbJhRKOW6c0H9VekD73SudYEQbfZRlQif
mDfMfP1gSLX+0ZW6AAcyRh+xOFbqUaRJPkIBQYmXW8uZ19QNQ8uH0EuFeoRH4C+2
PtFlCrrzbXEUVgKV7/FHBR6wmMPfRXLqdzm1Y8DbwkqofVOBp4vc+4Cb0pbU7NZR
itpNHG4Rygbq89Nm/9Ts4ZqyVa0vNEmQ+4/90nFVQo1KmBHhqOHjoakjexfypvKk
na9zI51M0c4BU7hGHB9ugNzuHNGGeoNKrvZQ3XVkUYvuN/uw7XOoO7gDSkxJ3Vcu
3RnzMvhXhImpPCXfNJeMdktdo9zROoK9lF08KPEzcUDgsI+ZKF4OsYbdRW/efQ3g
IVOTSFuXAHKnbMjJxMk+urLsJtfb0BG9VBZbgt+ctJR2dodiy/SDbn0Jwm9EEqvF
DCGTiGgdlcSpnLSCza8Q3nMcl7Ci9RpCIJWWb2IgTn80xChxTMd1v66Cnc5s4Dzh
a5eaysss3PkHzwNp9WH1HcwlukceZm2me0+QEcEUdfrdpeXzdHlWOVlm+EPwdcin
XgLI9W979ICBZ7G7j+trk56hvDmVCbHtN9fga7PbIWnA+4kuoEO/720h1xe8y//4
UumVnTuoC8xKBIARwGOLFKqjweo189i1M0pmoMfxtZ5K7bCbOIk2KJvAdqEPoevB
P3XzaiiwI+eOYsbiRQ8OhbTIeh1/7vZdMFGx0lA0vbp7OncZbHy0OXbr9qM946r4
7aL/Ac3UVM04Ig8eTgT3QcE8hFAMiRx2sCBvRapBOiBi4mI1a88PC4p9WHWW8liu
oc9CjxoSWfcNNQZRWFrkksVrp+lnv/067so09mh6FsfayS1VbcB635pmz1JbH7J2
li7yHaDNX0JaufzeML9/47P3fnKLhyJsXORYDBZseXqLPmqMfFmwgLLnWI8IuHxc
FdWn9lZrm2xTZxCmzbfonslSVfCd3Vj19yGU5HL9RAh9UFQuzjiNXp/Bw1ouC0SV
nbAW3c3yia13F6UJknmFeUS4b74yOEr8gRj8I4iPQ2YrVH+Ck2YpeR9KH14NoCer
/z3wTZhe0dVr2i208gvlRxJY2dHQeyRMFdEJ9+1hQSw6p7g/Z/lW9vxn1brrgVGq
Wul3AFCd1tn/O7dmU/teJzArjzrOtWcZ82lHfmYNqDmc1aDLp7Q8P9K051qNoBaC
doEmshw4Ci5oPY6pWQpDlRgfiG9f9mFt9MFqraGlRsohVkcoldePrDj7NjmbuC3Q
Swa6VzZvLqum+ji9WBXPNTykSrRh9CudzPEezUx40i6ohtdYf22wosdPo20BeR9Q
zEjFDll02YyxQ7g99hHBRXGTcvQV78j3oO20ellewJ2AsN/j3Xi/+7/jts6eW0h9
LVs05SShym5PNlLo5b02pj+QNQT6FEC8z81BpgdaASHQqjshU+3Z9yqy0/i4PPmy
zQYc5h2tAp9pzChWDx5uTqPlw9guq3HsHeYUIcHXnxW/Kcxj51YuzNBbrxQtDDbA
qmEFJavZUQWyUJeY+vjkkui5IL4Mg+refAVbGWIMh6ZP/6HaX1vEkuctnB95ZLME
gP0gx9/Htlktx011JrEvdgDziGsyhkfTZyzoIviAqj3p5+b+TOTP4Dovviavecmk
qsmRrw6k+9AybV8SCbhrgb/TqO0tlxW3jUbIMYf1vGXfFx1UniSMbxxXCBKlH+aK
MWsDo6zcF7IDj6p2eJC6E1FtZY8Too6MmFdtNEfIVGFUlOxrDD6Hl+j/cZ5ZxrTJ
OEyeYCtjJiuZ25juMvv4nL3CCW1yTxcED8N0/n6b3S0YAMjGmYadT3ADIfrjh5Ej
Woxoyxc5A0ADerKTKAp/K3nPAjh9BQjdqWV7uRBdlYrEcnJnJNaQhVMFj2buiiTR
KBK2QRctmqfN1NAGW/GZY2WENY7PmcsFIh/IRtzRT+NgzsS6y7BguvWfI/KK0xDL
cGlXEFD2gkUrfpg6O/BA3mvoFf86qPv3N7QiGfz6p5c+FpXp6fo59f7yVB2rwEa2
INrf2q/1jWk/5fRrIj5C1vdwLytNTJtCVGOsK0MvP70R5KZT1O4ejwD9F4QKSJfn
lpRAhjenFkARq2n64S1E4BNoQ5LseBneTPLCo4SX7A3qHtYzXICI92n3qZAa5/U8
i4zyZXhWU316ELsconYORgaqnDmak87RmcLNgeMlNTDxzm5ehwjUeZ32AOgpxWa2
DEFtoqz8rSPdUn9o9Fw31HbdzMTgZPv8kB+uSwI7uZcauFb4oTsHkDVwrarL+1K5
yjlPQApkWJL+OIEiLq3RBtnvhJBw29aVb0JAWeq1bPNi6IA7MXSnFIH8gwOjx5fN
xb161J96ZQgEbSk7WtTAV0QDkwAZAijrq6mJrC9LlazbfIYiFdc7K5fSUt01kNox
sYZkGTVP9xLLfmD3wazEpRkEd1zPdnrnTKu38WFNVIucHTEJ/pwFu8RPaBX4qhxf
DBhPi31VGzPsAxQ9CtGCJDwW040+eNGXjQ0s9a7W8PHxHO5X+7GIxfnNCf6wY698
bUHrNEDEtqeBOSFzyKT9h9cNRf92Htsy5Ox9TPGUFb3B/brHaEr+mHvDW1akVZ8Z
bt+M4Bfsxfck2xTKeAARV/dsVdu5q5hHnIocJmEl7+kYa0n2POukMB6d7AQTjAo1
6gPAK9LBOpptDE+SyNkY/dD+B/Sc8HkoOnCTARNYBQGOO2zBaSEBMUtI+8Cat5sc
G1whUs386zgFTFwtvCWjY5axcgnl9ZW2c4y+kB8PzsVA8nTyu1USLJkfMlkdOp1z
xiL+zUolAhZQCumptxv7Sz15UTbAmyeonD1TDFTXnz87WkRplaeKrtyBPWSnGkCw
6/deEQ/ah6UyhXSBh4Zf8jwFk87sqUF9UZZAlTtuQG353fLabwyVIx924bfbVCFL
2C0Xy2GmD1dd336YeW9GgLGfu22K0Th+2QlE490xJBholSnvkKZvoveFBpfv1Gdb
pe0XfohMxlSewKeSN20APFv9NAsZILItqBN26eB/z7depWQr9hISFv7RwtGUFdqm
TG82UcfkEYZgMC/NQ6s1Q5K5j5mk3WH1InGyqc7uePQnKHBrAgsli6tLQp0Vha9e
FZIYYrc4CNgQ6GFCTNS8YZsre9vcKefwg+7byncPbErqGoZQ2tydcEfsBG+WKH6y
1n95EldfQCnMJe+2WQHplU4dVTXe18KKwwk6mNcmH/o9y5PbPN4LSOD5JB9LpJ7E
mAKJJmGvkdTHBA5DF+RclZRqrWxvSZO2X/ZuFDIAx9B1oD7uV/7g5ZeOX23OmnnG
PCfO8W8MhptxadaeoT13DyZfBLusnyDyD311pY23PGMlEDkyJ633SHSutuYAp5v5
mOJ2ZQLKHP9LW0lKdbSUdQAzT88L76D97S9fd/sbauKnhDyeDt7RFl1BYJEDxRlq
8tvkAaaoYqSCD3a2JXc7qRO+5wGiP4qsATdysWs1kD8QlMvHPFUBaCXBQhZwJKH3
vX94Azrj69TLxH/RCHJPMI1JspTF+hpTWLuBimRxHzN6mC+S7gE/Y64O5io1bqo6
ZMa8fnsEaVqDDBc3m/xnsXk8yN8Ooxc+GX3lWdyhkx4RapYifYmSlqt8CcbyCjeB
T641gm/S7stKXTWmqfxTr1NpEk2HODZYB/nAZxtIfWiMQSyIYOuDm8OZRKuRPV3t
x3sJH5xY6wGID+CHbNFehNhybMw65/ubinLLlRHElWGMFF0CihNd5zCd6EjRUP+E
FtvBUm0Kji/lzZ2KEIyW//iCQRMlHI8Oqs/O0F1x7g0CkUY3hTLBfa+Klkv/cjI/
wOx7H4VUe+Njxxb3MzXYBRHTywspzScq203j9AYxApYwM/GqqEzVrx/H7kqDvAOn
MK0VI6j+zZntOUN5qmTJTbIb934k8AfmqpzyB9bYvMECa1LhsWWU93v5uM1kg4fu
LpUKfOxsNXuBRu86fhh0GU/QN84wgiwIYjqiT1cXurOQECgLmo7ATx7a6IPI7UeW
G2/vBLF26ZMt89DGyob0fUX1WYrFc/DHv7Z6ANfjkG1L56RgGM9A0MdZQwsObWyo
YnQlS+Ag/tl4ATWkBPNJR6IZqJD76/0DoLP00p7pbEhnCMXymbCCQwFsdaepNH9m
V37FyKUldHPJXWzqFdAhFyX4TSDolO8+QK4rjpH2qUIPgGn5/p1sUUOtVnY3pVvN
Wg/1sCe11y2Yaf2/SYN+ZStswAR473dnCd6I87Psu0PQRpswQ28Gj+jwhN1b4gKj
JHsUm0JdQi3ST0c+N5G/yu+JX3r4no1mub/Rtpy6DQteQGUFpr972Yl9+uVYRemg
fRPMKmr/W8dtCPsTCMWcY6sFM6V8lkgcAdBhAzT6G+lm4uCJF5c37xXN/csg2FZp
HW/9Nrrq+MRO1C8SvQXlmk1cO48j2IZBMyqKudo8aT4ZlPaGxBZ8qVRwabyX6Qsj
6BYSsmf57Zwwrbpfwacp3+GQC0oZ5aVuw7iq03rzTo9XLsgBa/rdhVay9FbRtvlq
2KuzcFnuFcH6WLh0FeAeQ5rRSW9E8kMRP1w0GIPIGA538By/Q/kSPVd+yLkPEzqq
Pfwu241UR0UMpQosSm/xJHhCLxkh1K+c5LRGXM2ZNZfKAod+y/rNwsE0O0M18nsI
JdI12DRA+v+Qegr2GaxHuy7B2N8GJI0ixv2eHrl2dAm6+5hax556iBPvLVfzYOJs
eg8oo5hidKMkRnEqzztbnsg54pIO+UCRNfM2lYeVZQdjsPY+iR0McJy9pZOJOM/S
NRL+XpSmglZueEmffuJ/Ge4kPE66+SKyxkHCIFFOlNmEVzG0w2Q0sOu39Vo+a5to
26YGkxdVjofxiY4OVFiQMZ3PB08fnNIhjv81bZI8sY6kzd4yeyX5uWwQWMeQJRsB
XaD4dOlfe1NMM1/O+wREyD+Yg3dKiAv8THA1/IxVUIV5NuskIXpmMBoCIdth///u
erZXgJpzDCQ4S2D7EVgy0+Q5SSFVruprd1thOUJNvxjg1F3RGOn53g9it2X62vJb
RpvK+GQZOxOQsWv7gcLQfRYZJoh9K+ld8y9n5fJyuqrxwUmoqZ8zb3cdH1tWayvS
Fy8dK+g56ABwJnZIIildtgGESf5ek/sHFPIofOX73akcOZst0dfPF0JOhqoE43Bc
Wbpic9YOBSyghcSyqs4/xqk3GCH8B0XhNlQJbMaM29KbTkaiN6MVvaHyW65lZshm
KhRIUk2e4UjhyIH/fe7A7X5CJG/ZGha9zBt83TEfQ9SuJznzb8znXadaM3Pxnxwl
SnRH0UGBitBEQV6LyFuDFJQFwk7YuHfp6ECvInJMBGq1y87qR0J6yCIqJ0hbDpzB
kTCRtMmLbOJAs5ichFJRwRB1A0LW5iYvQa53kkgjXvtpqRMnCeb3NeiNsE9ClJtb
yt2ivcDNVwiFE1QglCXLbWBsvcYYFjT25nF1b169+W3S5YUIRgzpq2uCQwersO/a
rHGuCuVa59Ibni2DXPFyjUCt020ViDJ3y4KQJ8r0fTjIrjB5+25+/3lFj5QVdkeE
ZvQZ4pL/46HrDu3DoRCtZRZs+QoWrYkPiIU2zdmZAXvwZQYajP4kzWL+4so7z5NN
N/VI7Q4hfTrA6v44ER1LpvMsn+tAj3jd/fYaNxqcCwxhgwFYTIiNxaZuyA0YhKRL
bFszx5n4KmA72cr798aIRmilqhg9BbufDPw3f4s6oMJ2bDUOxtS7X4OUIW0ULayq
WioSr8G5PrrVaIuYfKeI1O35XuIrsMDRU0Bfn544AHPe3MfoUqkh0V2wPvGxAfmX
0pDY8zR6DJU5AaVPEP6zzWC4ZZ98t0NKK/MuU8I9mQgmnfgfFXvX4/1Eq2sy57za
Ebsz36TjV403dl3wUBtXTFfYzGK1LIMn4LOd5O1QRvI+WQvsGAKVxKmdsmLzP00C
UHbHeioScq8y/yFnRhhCsSq28si70B3ubsuLQxowsy20SZRlQOcdnrLNUK3klJ2G
y/zCEeDMwsJmHkfplguW4U5Gofaoh181V+QZhHd7Q+YzDsdik9SxvK4gStd3pIjr
chLsXgIxzzKVUEuxqL3HCLwwwW70sKHRfetMWEU/QwZeIj6T5ECqtbTOJDpOqjXo
+pKtbcZy23JO+D9WmzOA8U6wMTme+QQ1mL4eXNDsp6VsfXRvjpv5IV39Ti9Yd/p/
40Q4MTKogyS+gecg3K3INuZZZGtWQhCWeAWKcojcHnfKsfwXEoDU35QUw6Jk52rL
wDOVjOYkwOyWcBLRvHem3mWGsSxjIfUP3DC+awxYaygLJv/WP4srHkKK3sKsWCpV
XgcdRVwe5m/zOLmSiDwY5byvWfAkehco9jm9TXYdHiqQlhSRUDBhpZdgAhAKUPZF
UtTfFjrxtOhoq2FtRE6Ls5uWaBg2Wz7vrSQ27ue8la1186+FZVWIXbhrhHjEyCo7
FbIR8c9rk7hyrjBIOly6dUfurubChQuYZxOos6cNsIJRauZyTL8cDA8BobXCPqrn
5DdWZYgphT27BEKAmSaqTiIFXlNr7AYTXRW8l1Z3/7A0Wb9udeNV8cgTID+isdxe
5ilZOl1t2ui+xc/1CdpV4qwbn9CbXNXCdqX+LMrzOp1uh2phnYgrWDKVMw9v2YiR
zMirujuFxlDc4anIuYCGVuLZ7e5n5k69P+6pYIxWlpX9xFdrOQh2swtutY5t+gOW
EMKQ77cfgkDUzuLFAtUP+xSa7MikKslhwyhQAh7cqJvRm36Lw2RT87J5yBcf0/hP
B+G9ws7GaPgVszkoJhx8bkHUnzuRiZdB38E7E+9gdliDEUq6ev63y3AFHLf0axHC
t1N4PIgA8rgspCBGUiIxALrX3PcBzCpZ+cPrXfrX1wZKREHKIm10hKcqeDUXEAtY
a0ODRu2FcjRBIkUDAth0WMt8cEi2oFx49KlN7OalNkhuXGx5dk/p5V2DD9cEluMn
J7UvQBtVIqtIkAU5lvUZboXD84VdFiSYxDHjOIKo0l8Uapzm8R3LbSFJvAEBrgJZ
Na2yB0klu0Jd11j3HjXWQwTJisY09N9YFONx0n4ehHR11S9C26XbPhNBgVEjpHz6
X387cGB2UZmL2psRSzjMDWpv84WtfB83jg9tfJ/xUaxhBxD3WFbtJ6pokhMpuIeo
IRmuRearDMBsgp0FnAFGvloaCXsnzdSA8FezcKe87Eupqo3DjLetAh8iAMD1TUmk
H/6wtKU6i8hdOxhEnRvhj4F6e9vLL0XSLdo8FSljuZXvxP7aPu86d+MtpZyu8wA8
hRqp+huXa9YvW+f0rqetBcGvs5Eq78+3vaLNqWvpkoxBwO56ABWL3bXd7RNsZmr5
lVlrL8tBV54BnUyYKRsdv8nrUMVS9JGexN/GJWN6v4jRHZxryca0KyLbvkDsirnm
Ge2PLEKGoCaj8zwBR6xKvV2bErzy+p/YEz1Ol2ypkBJt1T8GNT+um59cVsgARLTe
sEILZOUedU0v884m2ySzgkbbuWLPPltI/l7h7tzolozzuf9At8NcQ9KWPoCDv2Aa
zlUdhvVxFo934gCrEcwyTn1HrZ8K/Ntb271a9e0FNyo13xgOusDoCc0h0Bj87F8+
uAw00DO88yL0xhuBYaZlYFl/yg4KUIdOvm2MHcC1NUTfC5ZT/Jt+nAp+vKcGd5+h
W9iKdNcjRp4/KTcFyPzIWO+nPwHEQYZkbylX/maw2F7lpkf11DzoKAWNE3o/APMp
B5jdh8WphW2Y0HPyekDSJqfNT9dTV2lBVKVzJH61Mws4jziH+5s8sqg9navjpXzI
nQYAgK+eYsZDx6XQLu0SIBm/V6P2HxHNnEADBYn50rQfXbq7/Gc/h9m+m4miy6ED
3AgBLbZy09uqbmGtF2IGtfqP63+EhKUwLdPuwSWiX6abYNgTAinddUZ6ryhvkISj
g2+K0qyQkGAvo4RbGN25+NA9ecHFmo0DybYVpI2gIzjjGqDE2Ki9KF98S3FJNT7R
Qc5vdMF9TOp12aIge5ytSokFBqjsDu014EAFCQ9rNW4XjKZ+5Xp6RRbTaWU7dpQq
EQnQEj/Cj4AVt2ilFgvWRF7DYsbmYez3XmBwOqkKrzdSN2nHxXNuV5RFIfbD/wJK
`protect END_PROTECTED
