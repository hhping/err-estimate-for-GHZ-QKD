`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mxX3GUsUepOMg6S/0oQ9nt1bGTgviqW460WIAoS/G/Ciy9K4cpmf4lxnr8kCpu7W
Mh4Gw61/lLPcyn/O/wXkh3deRWaXQPxZ3fX5ePImzwGeQ/xv4qIVfYrN40ccMAvb
rZ2LxmBmJulDsCCzXMFW6OKyuOaLED8aQQdNO/DAHkSWtmHEN+Q0objtlnp/nrea
/kBhxzas/DSCCJsTQhPE4lQq/C4mTQKj//jI2k4apjT3yhtRyG+3zzH+4O3x5dkT
7vriXtjc6HsXE54LSUN2Uhnt0wXea0+ErW7ZBxppC91hovuZnbTymey0jpzKLoA5
4LjmCHtbLQGSPPOrK8AUKiOOlFis2Y7BqTxMdOKxM3oCDcpLVGMNBMCMmcqVDqbU
kgGPtrAIXhg+miA+Zds+fEgv052JZSD9FDCYDLR/DOBnXMjJ92+98Xrsg41H0f4C
VNkSp/SuBHXvObv5g4SRk2lnecVS6XIImLglWJbENBeI50EUKYz6kULsuFVUh6kA
/KZsnEAGZAIsHcN2wnoU99wuvuhWDzsizOOc2M2XsX1kwfXvV2rTsqsUUSKT4mP7
DWxBbD1G9x90Fn7TRkdKChG/azj0dFm/teXQL/wdTCFli9KXjaBJPDCSfJMy4TmU
l0fmfmURRXAXSmScMUilbeabIjvUSVEvjDrHgvSVMnfkuDxYlS0tZfU3F5HuwLTp
V+vvLlxtYCmfp/ThjEfQwSJ04bcWr7XyGQdlI3Lk+8a/2CP0w0ju9MGFKsqUzo0+
QrzsdmL6h3XlucTqWUy9UwCXMthGrQrmwOFZ+xK2jjjiOzrDuTUAGB/NI6eBUF9R
pozvfkYv0Jt+leYDVFYrpfi3h/k04F6UC+4B2MirA1fQinsINugGIGmcDWlTfZBA
Mgvjc7XjFK0QpkxIe8hZjqhndGn8/jd0GYJUKi+E5QKwqmNe216uehHeaGI4q1RS
oKv6pukv8wD8gTwv/iyLBS60Jh0Un1L7mbblgpwbWmuGkh3zqaCWT3HwgrZ5CNTF
2GaWf/XA3jssXrPR4rSMugqUqDLH6nz/LdYW5ov2ZfrzCoSE/sOMgkMPiQsIiPR4
Zbn/nfl9jP0AoDXgazdxTpR+JNdOaJvyAkfkVoMPGxkmXOmM0lPxMaw2o2Po1fhD
RSANqAQXK9xtE2BBawbf6yXpHbNh6BBIZPY66aLQslPNSaLhJhOiqUGrK3W0WnZ1
/Lge/TusGTdwDmeNFXmMzhRymrEezD1hH1XskJXCUIwxiSIsjwNGmaEwRIP1IxPN
Ubm9v9vpgzW805PdYojy15DBFJSVXFxVmXpUBbQvVfA=
`protect END_PROTECTED
