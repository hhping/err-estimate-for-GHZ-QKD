`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tfO+192O8T+S6m32Gp68GYoJPYQ8HqiFVVAnrti3uvSoy/DghY7/tdzbxikar4Op
IPCQoo7PFl9WOQg9SjTYgRhh1M4TtOHmODQCf+SCD6vu35H/DZwdLpqGooXrXQEo
vEETgfs9IrpS5ryBGkPXmEJ7csNsDunrxi0cPmtRepEf2W/i8DAwdKLJHZEv73xY
nGvcHPCJdFzmTERxuqlzuaK7RTWuiBMrd2DR2OOvYCjrIY++bGcktUY3RCCkGmOF
djpvjtnMs4/fi2xATL8G1P1q3LdFallIfUfh1NjPbFUoIg4athD5BjnbmenVJuXh
vc7Abx/+TTyQ5XJn+4qt5SnCbUU9CkISXbCDEzNPjNT9+OKYtcToklbTwi7HVQQ6
/R0U7KaJb/G4WjphU0W21ccuCXWHIS3G/ju5KBG26ty0IAdRtrvsdfGmKCt2Ify6
RTqfX8yKSZOfjzBEHcP3DuECh0VZKVY0UpvGotQFQTo4h1swB+rVeHhu0dOFdxzr
SKFaM8M2coA4CShH0ew99doxoR8FKhzRHWSORB/c5LKDLdKr7e6mD+ukV+FEnYWg
xuCCewex+NJCfF8fR4Nz+oXO5u7JyGJ8L3NGQyi3ZuaXet1YAArqGChKX7XQoxHT
GHsRaNl0+C3rmcfX28EXRZhZE1UNsnr0cBj1egZ1MlxR0hIoQbPhvAIADKdG8nvL
aD1HjPGDZLcXmdQn6NV55mDlh4A5/I+zL6qafYUTPD/Ei6DfLsnrul6yzLmS2sZb
FVoaiKdU0gM1I/AX7BS+hpUTiXGel+G1+glh1jUGqZjkxzCGmTDXcoTiNzN5a0+e
JL53NgYsXaVw0IJmndOaCIkJgJuq6Vbi0arslwO/Dm/rf59AzY3+SnmtqRaOEHr0
vEquDfx0rJTI6Lo4nVOeawPgnN9ZNQjyRfIUBetxVKnliGy6k6BdGJycvlCWqGHn
nf8x509TTwgTklYF61cMsnBO03lDLEd2pmsscuUhsriBQXowLedNiiVP1t0r9oLe
da7XDG714nYBGSMZorlMnlu6E51mwuZX8saqK3PRViN71N7kpv1lmhpMV575HAWT
lk8pRDnoTW6b/FOqmppXhwTHoLX3g16eGh92BNWIoi6VmDce1ViFGNewOJYw3ht3
iRM0V4JaqPJdNsaVEJDJhTEvydm7o29MiNIh1koswkPVxDefSQKHDFtHCpVuCQ20
zNs1ceyjEwP69uLYc1jtLBWIw4gQhm/9PcBj+diB2yxy4Ce/I+xVML6+bsrLo6jU
8cObVLN/FXnxzDXcNotE6eND/0Iz7oTRgP/qR/iFw9pVDzrnIr0vBhHCHkS/wXVM
ZyEVFan4RplahnoGEf+n38kki4dq2zIR4GOxOKvagIBVi9mpaCaLEb5NY/7SN1vQ
uRM52XGGWLskrkhJ+/LxBg==
`protect END_PROTECTED
