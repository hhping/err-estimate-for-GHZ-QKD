`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M/hMLG33XmCm/n2jSGA0NGsSLHYopnFeHCss9Cbh0OmyRzLgUjwQwF+54jfYjcqi
5FuOOAayVax2OWGkC7pLOZUUJU49eoaMFyuvi6nIT8vGYvoRufz5JKRw/ajokMNv
tsT6Zmd/Qk1TM1IiFA62WulTKvngaZxLSEhe4Al83adI/hVtqyfny/6Ytjswua2/
T3wBycmzPbMbgF5G9esO27Emljhx0+EQuRo31RT5oNfqwtoQMurYRAiQBOUgXjnH
VPyc+mw0gZ2xCa5oOiZEUVwMf3O9d+aNYo49oRNDTVOzRHonZx5VABEu0eUJzQt1
tR9lDDgvmtKsE783WUSQdUTZwsP73uEtRWqycRWTX56tFdgmQysajfS1pCG9ws7n
32uPkkN5CZWUSkwOncz1FJpx3j6QEK7bHIkkzgY7bVzP+tB0MOA26jKO+JkuWVG2
yvKXw+3NIgxYgZ9SewO3qb7oQsRbFwWxcPTt1b1WQkzlCtcP5G05wLDiNo02HHQ0
Ka+F/4vmv1bw1Wc2TRICzDDbq4PNwJzDjfOOBBM63AxfAKNYC3JLXxOWCqulh3hI
dUxQYtUY0iA5LtC2w/VJWvqts8/lQKl3ln642n2X1kKb44u8zMDN1sKIMVbjD79s
c/ak9JQjXPBYFbbuwOWV/4jQI2fHEHb14TD1QESmkOhfOeXsjD4ModEkGEtPjdCA
TFo0GqMwG8r0gKAdarkeko25A3mECGgXM/rXZJA3t1p5yXzPjkh59XFyfQgTQzBM
Tvh4htR8GfMiVAc9MJ26/yIxdKfVmmMb/LJtjedO/qzHjps3dObt/5g9+e6lUTCx
e4dSenbndYlduEFcF2R6BLl7ysXaHn3aFSorcZS0vV1FcD4XzNukZ+1Xhu7aw2GP
HpExsrz0nvlBj+5UVFlQ9dGXUQDdcKlbKxMKhlesazFnQqQ/ZUtEOJiqmTDWqUtv
1eTKmgohX7C3xMzS0kUan8CetX98M3ddA4ucDML6VToVrSM9/qFeCciNnzY9FWZH
BZBvQM2BoG1pyPgxoc0dgXfu3AaLfNck7VRZpNmfti1YHMZyOFfkPpUHOheGg4FR
FR+jp1q2cxB8IPoFWEnZ53DYU7Mkz1Way4YuCW/sj2dnJy29mNLT9kmdB5EIyVnd
tXZgh3rOdtJOR91Z9lsQMLAOeMGjqNcMsts+BT0TK7QR4ixuExqpB4LB5b7apcJY
ONGD+D9mv8y/lOiEkVwCeRfTthVpRE7NHI+MWCgk+v26Cmx2DCPBrrwsdxnLti3U
U124V+BQR5KZVUgAOo8z0gGStVgOAR5Kjbm4cwOWZVf6B7EKa15wGDvaIqi0v2gs
SY++DpLpiOYChA39DY3omQeI6mhZCjtiyg7mei2aNRXYju2BB6j0a1rVrVXtQJnA
d/hMyCTT/BZ6CU3Cd6esVHlKAexrsDNlOqwk1aQlVlTmMg530/MfmOrkd7uM8EpS
kvQBr8vEBJwmpoHgzxgWb9AnB5onw1Go4mJsiN6Jev1eiw99uysuafauzLef0hLH
XShDxMzcCONHLsdATIZ50/GGSrktepCBZMUDZRT4GsMj+9v5C1b71VR4klE6lqIG
YChesZ1kvD8jZGwEMfsJNIyHiT3ny6Jp9IX3LM1IGtOk3SSI7X748ONVUBKzc2ou
KoDZzJkwgqBjUEMeQt+iO7VMiuxMsmMocd5INGGjHNjCDJ/C/TOmcRPCJ3QbduM8
PJwY8Lh7FABQl+TicwhkfsMPcXCUPKLTpo6F5ABPyFxQyQkM6YcCV7mkEF7iAqFb
iTrZo+VKI+LymJcePP7eh1hf1M0bNM2O+wXFdcEfCtkLQCemDLXqE0CAvnDqeyPX
ytUctBaNkHOTbjxDgAJpdeuA2OhlVpZe/v9Xywl74rJXdclQHPC7ETC3lz0uKJfa
`protect END_PROTECTED
