`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZROlqTmjUWBiDuBMwVB1D6ShCyRrwf4/VdnM4iNd7aN5ZYs535FEoLKgGiIAF/Ly
p7tdwXfoU9gQKbgVFQ3non8f8C6f5M6j5Ef2WLxBOIrakVQRHAuqWfQYYkshhfhZ
3qneFeu/qiEgSJcgPmu91Ssb9IhssEYNg808VkKnibyybkR++iRZ1KyQzdAJYaVn
KgpeQZ+s4K9B+xEqAfCFL5DomilHeSVtTa61zfmeK7IgSXC38kYbkIRiDYeo+kwr
1W0l3uXA8xXMA+JT3g1x4XoFAsdH4kBkfGTu2A8N1BVBsVZIvrj+8jsY0DK7855U
uzJ7Yx85cdKrmg8TIOQzz9xMZ399tcRoMgm4aXC4PBMqnQnaRT36BoJcXGimHA9W
`protect END_PROTECTED
