`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jgKSiJTzvs73kQlG3ZsI2n8kEvwrI1A9aOY0uJs/vil5PfwpoHyvp68BkzeEW7ZU
fqTQGU7YyVRIylyXpPhBjNY8ob+GG8mUzKawpVOJ5G+rSrdhelba/i2bziMKeIUa
MfxpedWDMbBmBIoWPN0OiUQF4w6Sk2mqhomQuwY69D5YbAVOTVmg4/rLGIVKFRAC
oLZ3MaTQEwFN7bawCGeVCzwX79VVUoB1aT/HyXk2SNEf6m+H1mNt5DyJ65J+HyPe
QJTCUooo3tpjxHW6PadqeUSgx/dcXig8xGrV15A/4fwUpwBagTgsP3Kc/1ugoh3x
bfXDpDngByJp2TlLboEac8hf40qTtZusts+n7e/q+ueIamPmZv6Xt0LOtPw57pyX
E3wljGRU20Ez2EGTm6J6RxcclgQ1OoHraQshdKoj6o+A58LEeyd0V9EpZ0l8dy5M
Tn+WeZZH4y5RwN6yHc4Y+O+yqobo9CBBj+guft2+3Pf/4W4UjXSPEEPp0dekrG3a
5JQzoapKVkZra422r9jSaA==
`protect END_PROTECTED
