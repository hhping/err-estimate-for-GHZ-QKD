`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Raq7/CT10BmlPbYdJ1iHw03wz8lyBVA8yO7EMj3hic0x+HkkffPsWVzRSPgWV57s
7MM7IdkO5yDE0sYmPZ5KM/9vYsNFGXbYv1R951onZK44jRM1a+5Eh/aUPYRgVtjK
vTsgCJIyz9zWuE9sw5rkbNvK0jEER1zlUHVRh1i1gyGnjzQcpIYm21FMeV+pF6KF
r/ru+64+7Wbc4qwB066E4Q852h0/BaahLvTjJreuUBQ30+n7jXpuuz7l9UvixylC
SDaYR1dS261iF8cI9Tv1ox/arlDxwKDpp+q0GPwlZ7Kg3S6I/Byi+5NTfarHRJbS
1tewmHnqEV5SVI3uX/5j+qm1ZWNcltfMPsyZniqnT2bZCc/2QUYQOWMdTrLyMRdo
3VCP9T8vcp9Af5RJydpOopcdHYuK9MZO0YW1C8Ybu496YL7fMcwOUZ/j+/udrmzd
PNLNz59lNtoILXcD/AnG6vafDYwnbahNMoUoP59sFGpPWGO11juutSpYAL+El8aj
TNOS/QDXQzMP+30+2qaTp5cXo4E656rMDuf2HvvRLDi7m0h1V4V3vz+uPsKhP540
VZlmnvX9YGPCOD6cA0tzzA==
`protect END_PROTECTED
