`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y+z9WkdeiltSF+liHa6j9zaqdYO8XOS0RcmW50sa4I3fVJ6vXT/35CetEBxJuvzb
7tu+H34SR8gR/iCYHMS9ciYrSe3Kn2qSPkXaRVYqrvzXXmazU9/zGbUqTgGpzoth
Qq/afCaszl977MRQugbp13z2uLkRsWv1+6BT0u0WxSn+xRlZ2iPjqhCaWnYxn661
UxIo1AC3mStMYB9CUxHbULqvgf1gLuDQ3zXm2W+bZq9FOclnCwat0pg0C23RxIGk
qE/c+1+Hc2HrqJoAFT26uaT9ibXqOaNBCibd+DfyGLTcm7ykCgxWv0guSUz7nFgW
HZuRA4CRRdmruFMKFAJ2IJC2VLyDzIn6PaBE07AkB5vCgNUCub47v5L1WdXt8cuK
GUmll+vPy2heTgHC/nO+T8mUW7WphwpAnSEf3pRL5uqg91vhXomC+mkTsfo6jP4g
OH3d+/wIcNQ3vRJm5sN/4jfHtiTo4Ih54LRELlweDS1jRCa8I4XAAGkVNqBr1SNB
wLY9jpJRCsQUrgXDidvx8Q+1bEcwu9GSDr2lVxYxqwnTtk+rHHRnxbVyWpXPx7Te
j366ojza852A2GAc4Gj+Y+BFPaCmayCMsrIOW5PnsBn50qKcTf8BO4sPyzal69sc
okgvtoyAigQfcFothiMSpDnm6Tvx1cZi9Zo4q/OYKPru/xRNeIN6OT9FmHFYQONy
VVvgAUhCpCABr0y8aGtCwKZPHXlEPm0upVavwsq7TK6P1jdcHuTCXPXYVsKxoM6I
ohhcSSK9Hlr0F9tfeLkeRm38lWeCuQnXcS3R6AuKblqpnRpAGBzNa5Q3XTbqzI0v
B/Q2yGqn7LGsuoRIX0pL4oCPLjdRmq0e44io1ZthJUwyHmWjOMsX5f5JttmWO6+J
yUQgbmMnc4Y7vvITrexb6HZOdsT0ZbLh0ISg8pGh2HjQmLlLo7WyYaKO5djJ9z/N
k1X0Y5ZKoUEHPfocaKMplQCS/TH+MHE2APqFu+INXyLxSc9CRwi/9IKzsSi8rT/+
yg99aBfz8stzkEzjmYv0tvCEUabrmJnuwvI7oIH20a26gIneP/1dylKhvvIQ/Hj9
QrOIIXBsXgTZW/2mJHkPo5D43j664j90wg4frxb59e3LxAN9iLB5z9BWEWalnDMs
48C94st/aun3EoXOO8cIWAnifjncm07JqFfinv35H5zLoo06UqLGsMs9lQ41T9fo
VJPnnqPJJGqBz+HFYKoMblStC21APMwMEvqRnyLrgSxIQXg+X34y7p3/1kTWBAlc
UA1wL4UdSE+WgDv40zeXY4a3anYGbqkiuTnqlFTwA7mZvJRKNDX/NTkZ0Txt2yVN
BlIr7Cfh8r5Di8gIEgoGf3Ctiz80eaEkmuFYY1h+FiYyapd+M45iDdf+LDIh55jw
kebtDnLFdRSgXjezlztekUZtjSdEHBgAWO46P/kNGJu2oMbv6ERZj0gxPQ+rN9W3
qxS4Vr/JaVIvr4BQl3SYBHkdjiU3DSycXe9CYK5CNw/WBQA/CbIA8SPtfGFClgSU
WEI5fzeOz7PMaWegX9mpGBdmG7bDmazY9VQU9AnFpKFSbNUmM6nMwaOsoB35kGWl
mxogFB9MneqXf7n1g5bPIpqD/nqJ84q8dFRPfvVYuY3jpYM3n6nwQUOxjnh63FOW
EN6mdRdtY6AXbZ493A1KxCGAPdiEYkueRx8U20mSIts4C7e+FNyDLib+gDPQK3u5
JFQIvivRl73FBKi9/MhFNm526NGCyEsd3uktNm2gQSpFsrHMH49uuINqWSmzy1Ph
urzO4Jgp+VzsApiY3K4wfvtD02vr34XouB5qwcpu+oDohpTmIVdyfs/D+vSMAKsa
SzFHLpphRePOaV2mUHe/6tTsDJi+iRYVQnsgu9HQq+CKuKGnABb7T+5QBJbeaHKk
dTQmjbgMIZSiytEW2B69nzVYKSkV7Y/m5gi2TQJNabfmc1hz6Ohidww9e0RzCgo4
Bg7JV3b9iCBA2y1O80khHoerHAXDZ2vWwakEi8Yx8lFSooc4YRl6wOt2VIy+OICl
bhe6+mfKOfoHkAxOCkg5KEJigoQaZA/cg/x7wSpnTkbxhCIqpIAVhCe38jui4PJ4
7gMaI0674+UV6uZGCacIx6lhhzrCKkJmAQu7zX8OieeKeeUBjjj+FCayh4fivaWI
RaPT5sSdyGRX3AcltxTuscx/0kHXbuP54FguZKHi12BazEvCltIesKN5wPxVybzL
2f1UvdMHzShVccvkGCGwLKxZmJ9SAGBHb2eM9zWSx+akiD2C5DUHcGEdu1Go53B5
EGZiJ2wDi0a5f1cq0/5C3Hm6ksQG8RlYxT28QMfy6CO0uQivmjZPMuhhpbCKsIxv
nG/dI6L7U2+bP1uI7U0djIjgZLN3lCAbpPyK3dDR7g/R3YKB6/fGhvB4r6pnxB2n
p7SOpACzlvG7GFPNkYvyvt33NbmV9Clcu/mbLtlpNukKGkobUHbmrR1xz2CSZOt+
y76gttibbdH9fH1YySoPRIN/xEI4Gg1n9CO31osdky8oZaHwhsvC7VgTADDd27fb
F9I2j/yOemzSQBfNKznCGRJ9lgMxzdzf3RtjYwX8ts/Qie95ITFsO9G+tYAAAcJd
JkIzml7nBDCXhnlBQZgUy8v3AOAZUbrOtyw47446lHLcJ9huwnVqA6CbGIOWaZy/
onOvIYvfQtZC8h0lJSa1NIbq0MjRSRu4sx4EbhqBmVn75onwxRqf89fwTAjgbF+t
`protect END_PROTECTED
