`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wekrE79EBbr+hwvolPPMVQAHnpGhnX5hrEU7A3E8ZmNaF2JGV73u5hX/O11FMC2A
W8yk5uq5/Z9f2gcmWzr9CtOXdFJweh98+vsw1jsy+LfdQTCmIJJXaOVk5XurfRQ8
vaZ+sW3anYfxGSoTUuctsj/ByoM3X1fdqMyvvA2ZnrbPHqhl/DxtDjCXxbaqyS8c
bQuWV9SwELKG0r2zhwy76diteL6TBxHAnAg5XX1ay1ZRTOloHmCuwqV5eE6zSiDY
xGzf4B30TaUKrt8ScqaINw+9Opmh20O6NtXX+mFH/Mn6rKdG/t3gZT+uFTWXG9E4
lwplUWDGiTGI4QaVFE08YWJo0vbDahipc4cIZoULxTeZs1MElYkXvRlsgvK2PUaQ
BLkQjHC95cM6x3Fcn2r6CYW5Y+mG6xmFoCGauzwSOs6XJvbqf7XF2m+vwjdfztr4
xGROjX4sja3Xzlfv/NsgWnsBadxcuDb0nU1/91Ow4eM=
`protect END_PROTECTED
