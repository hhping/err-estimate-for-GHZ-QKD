`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3WSFn94f6UFszpDIdSH7Jwpkwk0MaYtKX6AswmMfMF+nr/tcnhMFhAvxg26yxeDj
VivELDN++dROF6uLfJ3yPRjKUOtZaWY+B8jxC+mfS7IMfZncTm2jWLuHuMUBQgNJ
Js7A/y2N2Unm89GFUEtu6LzL6c9gRhfwawAHkIStZw1X5D23/tmMh2zaZ6UBVtr3
MnN5EI7+3eoVU0CZQjX2QuyArk2tbV2KZy0+OckbEFFLg6Dtzyy81lAQ20OGBOtz
boJmOoQcTj2pnP9+s9cSj1gkW/CVaCunoXfMoi9dZ4CeDapeJ9J2MJ8iliHYwIuI
uNbe+r2Uh6JGaXlcbwVE+Um5YjObS0hdZ7Bie97B8fT1jenzdAzQ2Gi1pRvgKYT/
LcXmKGAwk4SMqOpw9W2PMwfHcomG1H/KTfUXRWygQBJmXkszGPzhE8OVSvlYhA/X
2GZm1EWey6iMacBsrxi1CmcbO1ZtKAEY8q1LZ4Sudvh4YCSU6OcXTEfhMrNwkZbi
HsgN2W9t1PjGfaI0zs0UxCesfzahRe3kztPY71CEGy85R01UDOfnNc2s/AW3AR/G
pWDJ8VufIe7ujubuTh3zqR/5qeN+Xsxk4/qgBK7a6OlAm7GQMXro0Sw+zObFi+wa
BNTmgqx/l88gcWcmjnq/IWibEZh68cHuNKDXiSpkwE3ouNqOAQYUuDQ3iloY2FVs
bmRbIEf/ERo6GK1BpkXVXqXmGrlMexrgHggndg/maE5n95z1g1SNN9dwmKSTztxh
c4qmGVHrD0BcUzwe8Sq/vgN63Ra6fs0WBjSEM9aBqg6Fs560dETd6HVCNq9pu/Gr
0vNF97d4nn6zmpwRjyFQbnM8GQQPo0lhZDIU64VsY75N8RtPclV/ehelz7GLjmJu
mzbUgnPdXfQUw07qGslwhXQbybJf69qMOl2eMs3OG8QTEsPk/pxQpEl+KrjrbtNI
9uwQzRk1NaBR7IYWWxRx4jdHmGhnYcfhparZ68P1+Z+o+GYpOak8WuN2tUWxwJKe
Zuo0+ew+HhwChHgBCkaZ5/yrzJzCKa1q104YKN8Y0APQPfF/wH3AbAKXtWMdmQ46
8EB4weSPt7xuPrU1U4qlq//9ixjOvuPK16r049Pe+2dKrJJoYXwRB7Z5u8Xuichd
0es3T9UNM9JN1HxD30d28WV4T2Fj2Vh9hL2YA9TCcJBqGZutnMGsZ/jYsE+udC15
GTlRLaDe+/QbhczH371XLOvOb0MYWk9KgecpdAoOYYpVQeGrmb5Rn21HF+lfAiPm
ha+sYs0nMJCvA32CUvx+cNMRiDDVNCKLMYn7KAjodyBXygxqvMaCHTcuvMMabMmP
kf00mg/pBu8BoEtMLpsCOZhW8KH9xsyiAWhGZ/HdclaGP+o4ofvU4q1yebk+iJ9o
1w/B3W0bvBkEGtv/RSPPL7I4sEbyfDUSrKeCYFPWJ7qZbW0YYFCvA4TjrduHMFsh
aIaj8m3eeN/kOJd4tGeWoRwrxhVjqHnkaYaRKojeLqdyR8N/Wgdp5Qves80S3s+h
T3jntnSGrIurV6jww8fS9ItnIrXRsWOxAJp6gTTUpcEoX9PBL/P+6MlxCVPmLYwZ
B84qEQHD8MUVBOkbdqPplsb8GzM86IkQ+A4fgKreZkZGYexa5lrRPFKMBXi/y8do
KNFtaQiF5JDuJkdpuCgEK/60ba18q2fms0M5zT5jSlVkXx/wO4OnA0NVgu/sVcLm
5431DfyEjKGxaw2rPP9d8ZlZD2LofQZyqneQT54xfnqt7QlqqqXWwkz5/HZvC6ug
0sqw/0LKYL1qaqYXDgD0woWp8DON2f0fKPRr2tAchYA3z9xMzvx9oT4lvEyy+6GX
BhWhvu9229TaNgFhKBdR5hm6TBaG9D0LdlkzE/onaR7zvNYhO6VflkSmIqTB9M89
aFHCheQQNSKCc2KJ2lwpnfHL0lybXUJ6L25KKuM6ZA+L5rWU8RUQaBPfC1gypFjL
5U37nxPpyn/IxushDTKodvI5qUzR06weWpEFTh3YiwEHuJt2bL0/OxrNnE0Rtbv+
KCYPPaIx8dsPH0QbBN21j9qxYPPtCiXJj7w+jMcsysx2P9hjgOb5TtfhCE/2VQTP
b2ecwb2PTOv5qAF0LA4WD78AI3fCbfvfWz1SSQVoDdixoETTAu9MTsStUl+VkJX9
xdWSGmqiYL79iaOYaXgG218TGi+k6A5zEKrqK4a6sG4JLW0SAwVOdGwIU/QycSvV
vmAV+tX9cdURkLiY1aHt8dPc6jxUyYAdLALooVEpUixhpOqEHA22s6JyG5LF0au1
YTzPosJEZ6I6Gm5pPARGZvRNA0L3OBEELIHgx/gTxZXMGQBqKEf9WXLCjrpuPDEi
tlccLZSIa/tqcH8bQHGCsKn31c6dXfOgiXsvdkJI/HzQVn5EwoWU9/JSPRA5Hy9m
7786FY8kqcbN3JtexB9shg40i/SZbcWV9c4FVMhdT3le60L2uC0sgV9KJ7EzmWT5
Xy6WICDEFmdXx5quUUDSsZreOWSQsFjPDKBY6bEiJfRhlxXEXrqjrXo6tpQoBKDA
1bQBtVQtYmjx7Xp5AT6R+sOLQKY5bbKMZtYdBli5zrFQ0pBzB/a0yhXPbIUAD8rm
vBe+Cr1+JeYlfd6EYopHMx8qDKWeA/dPwrQt6wyggHphX2v3qAJlT/dfWO3xhghK
+cI+k7XcX+eYr4BQ3SmzXl90dyPkpKhG9JvvQqLBVc4q+CHCd/5PvehAI7MyhxQC
2FzznoC/FcI6xDkabXY1uizC7R6/jMnmZ1JYwB1ynoJNQ+ZNtnQwOQWbPGMiPk2b
uH07m9aCF4UYypS//rqMaFmmqVHBOCmOWqCltA22Kb7U1ws5U3DZtaAnIwC6/TXH
0wsN8avR0EyoUNqELd49Dlrat/CsyLB9Ql5GpE1yHI3NapsV60bojzrNKEd4VG0A
V0JbacQUZ+X3CSRemX7tNC9bgMOXxGnFuCmZa66KSeKxUYQx2EymAdi3ofrK5WeF
DMnv5zK/FCyJM+w9SkdSHJuAP3SfeL9UG2M89yG4+XmRzA8LgzBQKGBemfQeRt1L
Qm9nwPqPoCO7JADQBQDtWB7pBa8SSKry1PnjtE3cjobb5uPHBixDxSENA0AO1BZo
I38K8qOPk/bG5nj2NQej/LGDo+oCH0/GzDccCcZGlmQEJ2lQCD01AbFwmvBZYwoG
Kdy2+GyzEB3zhK33LUGibOIPDDJ9KBxlhb33ETzv7O/M+vciJFrZJbttApYQsaN4
O10x5N1kaSnvs0O1QI2zxI7C/JmDi/teEUjabEduIU1PM9rZGq1sjFIRbikmcqXR
lwUEmOAWtWymA8qOVct4pUhmWb80GRSZo6WTs4a5VNVRR0oKHTZq5e51f3LV5ykN
NhUMEpeUARAVAP419eP6CJyzRs6OEVSQGtv3Wjy5zx2FiLGa23LhsY/d9oh411ue
H/Lp0JwBBpFzRz9TR67sS4MXfNmfXhAwqShsDlvblZCIjQN6zoJM5LNP0y4mMPah
tHI2+p1fA9pZUIxy11VIYjvMUdqpvw+6E+u4hM+WdTSLAwYYTf3mB2SzZGZML7AV
TMwWAB2CAiR/grsKYvJvGJp3xFYzQ9KIlGYlZYNzFnMtPjMnEDqUs6POxMynOMpj
757Bpeu2hJab6/SPtRquWEkZ7rE3cUauC21rtuqcCbaDMPRS8sTCUmH5Ra+LMFSx
JmRWsrcKG6QBz0FyoOwog7Wc4An5AMDy0CtrBvypB46blbtQRmajz+Lb7e/YAi89
tPH9KU/24D8175rEoPG8IpY/g+9mxTrHAo0eLrufmsHDq/Kj8MrbuG0DNjzVs/EK
AmxDn4TwAZQxBknbaEPiPXHq4q2+25+NkeWGZ1ktzMYNnloFF9kAaXH6JXljShED
AsjNepORxfFRefVLIbGOvf9kVCdUmPmUqEPBpkqHufcXXERGesYZEJOQZDoE48iB
S/9WdnpU1tIr+wmfu344nNwTSfbzWNFges0ZI+Xjo4voUy2bEbsCwl22ANGhAQBs
q0R50KJtRdMb8PH/WPqkD7NPe34xp4ryeuInqjQssuthjmV+Fxyjhd6PVERGSdVR
maCuZTTqHNW8o+gXBF4sYd9odGyf2rSGrJSoVBi71wB4p6lHucA/N2JMsFcuAkKc
Jjw17uD906gi57w4XwC56NvsynqT2H0Y9GxaL/73l9+3Ayik3Bw1yBn9ANLZh9rb
C2p6EzCtDwme/S1++pgETDut2UR624L5KO3TODI2yQ/Ur6BhhdQsJm0CfkomZY5x
IHS+JT8jY4XlxeYJtczeSVzNJca8Ih+ep5Kpuc81zw5Zck4+79K0zbyOwSikz9mm
NuXnHWoouQDkwmPRsbqnHi6IwqGxAwNczai7XnlV9cWyY3K3rVxzNELhCzfUWryx
uqRfRZGdjEpp59DuzXTD/nIMTZz3/MCKYYLvGPcNGZDCuVTqMj0aAPaIyG1DnA0s
QRw7dQrpDl9ReJkHf1OpR/r8ZNbtbKvv/WduO9tkFn/4TItOQ9u4EkHIdnWMec9B
F6deW6ROaM4GqnLYLkVbG2uQeyIam0iUX09kYx9AINusoaFWhGg6/Qd0wGQxcBuL
a/y2a7rn4vDW7TZoEJtkiosulwN6uzW9b1BVt1CUB5fIqnXAnva1sYuMgj/7sfE7
ZR89t/r1Qlsbm7CSzBgbWr0Mi451FZDMzbztwLQzewy/Ts0rREHF/fTnWrvIgIDy
AhorRxa4vO2Hm3yCewM7lhDKm4mM9TtiRKI8T2H1cl4KmhAnvqdCKncod0F4O/7O
uziEv678cq29z9OdieV0KehqxtpmeDshWbyZWZVtbckkQbwNLEnXSZuxgt+bv8R7
u6QDpW5xDIwsF6ZGM1Pr040JddDj31WOVaSpOcmdSbujm211N+m8tx2LDfwOI1AY
uWPHW22tlQiGBVKymxiOIKVh2kWpxxHIuog2rTngEz/0bIuscJpNP6KUOqljiG1C
KQeelxh2CgHwOx2ShqdDE8M5UVGmGEHNSjBrr/XHtZCGb+31GuuUN1CkgiGq5CJo
6pY41gWGoJQQeXnUcgn8DWMInIfbrOq3L9edVG7MjkiG+rhZqI/r/46CsbSQlq4U
t9gPd6hvFxHkr9Yx6Nh0/AMQh/S59Ytxp7vJOiG1CxFS5l1+EAWcSYxmEXhXY7Qi
BoYA8KYiLEvQ7lr5CJlJXz9bUcx07vItlKnAN126wbBdcYmqKzq849gPg4D4rh5z
I1XX4a0r1NVXsahvpBayJEGzBQ1Th4lFtb4LhUEnjhU/OKICBN1X8Z0MkH1EN3Ow
RX21RTbWt+8mP1it5pTM4dE3RhkUkLe9Sj3wdd9+llr60hBsfpYqM9O68AdKY4v/
JKc6sIB5Nf/MqE/6CZkVTu0Nf/CDa41tGoHBUefgFcG32xYjjxE/o3h+JrqOrJZM
EYny29JB0OIEB8szvmcYisWqGa0pDMG8xYxbEkZtUr1/QQOk1dV6IdQm/Pzgaovi
coJt1IQR6slwAaDvWEdf7bOhpEiiBhfo2Mu/E1vyRddY/OlcyoTKgJIkOto6eILW
7ge3EbeuqZtIPTqlTsBcKm004t852DC3glPhlXX29jDL2/GzxN1vqw2qwoipSUyN
GAOT7fyaXvcJbqJcnjtp2UNyMXhCOmquLE98XuH6kSPWkL9ivtdESOR9CTo3/PQU
YvRUTj1I7PuFJaugWtBMmttG9qHHcwgQIfqT7vwKU8JmQnXwvpJcm0cm90sPwevB
HAaInmQuN5cMAyFrYBzn5k2cSdB6ZvQrDseRc+DY6FkJIxUtFNPhSBKJMh07IMXI
DhCe0TpreQL0OGGWneaUc1zjVR7vT8pXqrRBCb2rB5X869sQ4eNkYFsw8WtM1gOn
DYjSFhCGtcG6j7M0Bh71QHx+1zoakcEvFb1xaG9KN40eF2JG3slb+sbs4hlTliKN
FVeejAWNypkksoUNxQAWwDbq9JgPJ993tRKPqb5RRJlgst/80LbQ5kblpbT5Js/G
SAJ7eyfur/GtcWzZt5vsiuJsok/uWoykBeV311S18i35Ne2YzG9Y1M38E4kJcjO5
WsRG6ogejAL0P2OxuwU3lIUaFL5fpfO3cVINJPS5fzoCkshNYsApKstDiCvftZM9
lCQpSBmKqB+qbdTkJwqnJP0cyHo9ee3XwgMlRiDCH6d05wfanlZJTHn65M+G+Zm3
jroO4/+VAJf1T4t5wuHMoleDiVpLKRm0xxK7U0QSW8rPcs0DXQByG4HyBvEShi80
ejVTzkUIsIyD8lbJua/vZOnNxa71EsZ1g/Pwb+TRUHZ87DZjpaykMWQEO+S6MW7T
UkqWCA051tAYMu+SkAKZfu6Rh9vYAVJDYo3guacG7q+tJdm6yd/LJmkQnShdLXy1
e304u4aUtksV+mMbHt+Pzb2xbs6kUsZeNWLGL5LQava/rcF718CEfjd63IdsI8Gd
+fWBaBn1St9Nh7y8+R9QUv3c8uRrd7WUGtWa22yJA6MeLXixJ+Ge7A9W25/ouBNu
wFZ25Rp06RvwGHyeM+tqO8nU1BXvpXSdfn1joasT+G8g2kJ1KzaoIFNYS9WuNfZx
kjTZ41vwO1aoIXBDslAHxQJP3sCstrQdLIdSsAZ25n7eKfIP8m8/dOD4XRmUgMse
yPvjSPL41CKvxE9HgkUFxa1RmIXnQYvrwVW7ens/jhFrJAsNkNU9zyL0YG98AGuO
d+cuFy4gj+m+o81UGGBYnNIZm9K4AqN36LZ/CTUsV3uHWlejV2IpSrSSVjW9ev2L
sXqDgFw5P0YsxAv/s3V2DGGx4GAt/K7xdevrsde7umIeeN8lnYQ1j7Gu4IWKC3lW
9fihEQgFfCBWO5FGBdGn9koiSVnRqfd4PPdd105WnppUoq4ZZRkCRrHyhOlw2Gl/
SmdPHhNGXxybaI2/pnC/nNT7xlnLAnXB2d0aNCoaFqTXJAqT/r9X9nTQicvX5dzS
9sAicG1omd7oWvRMIL0G3zxk/7ioQaDBjrkKqbHp7sSUXs4aTmmtr1HsBLOzsjVQ
op+jKjEH0bBpcz2WEuYIzlOoQHsjZWnMuDMm9KkPEyUHF5zqSnyYZVJUU2MANnht
NSrH5Kxf51JPgaloHfahS+ed7MS/m8eXBSrttG5DfSX/QV9Wl5kB8aFNemT27NUm
93ESHPguwt3Af/lbH7Dol33EZKoMymJAzpKPTYwcqJRvZgJS18ApvtzmhXxBypOo
+mA6O+PRN/v5M9Pr/IA6JKX22DrshOUL3GrfX3Vrx3DXLDm7PClnMuaVn0UHmCL6
wVkD9jf21uPO4Mo6n7ApRST1kAiBwhlusAQ9K3W2id1SRJaiZcljfpcPBlFpv+eZ
WMBWIiyzm/RXsNJylygzXFYW92o7cQj+Kpj3fP+js414DyL62KhxSGkOxZBb6M+C
eFpx8FJHMQ6IM+YRsp6lEl5gR2d1WZ9zKhFOdfZdrgWTrdtnZ7ODJ43nggvBOK1h
ZjOjRmSpim3jHkBQ/rYlgInIEH4T0L0WkE5yTBQBeHtZc3VHaNWHXTLSMFZbawVT
PHzK6H85iaYprUl1RR8SRbuQv3Etm1vIgfObTBjJ4oBPfERhaAkdhMe7wvdKExSv
TItM7g8ma4RfLAZcR2zsNhlP7iyFyqfTi3dFcqYNdyxnJV9L6GG7mKG8dlhsNodG
cWlalmBUQtQs6hj+GkXH4vqIHXyoznH7Z4fqYbNO9m+Ofl4zNeDE/2ko644RpPIL
Oaod7YwC4MnsqEOOWjDWCsjIhzK27tcuAFotXzfjeZCQbYBaVDnMyA6jIpqb2XWI
PJwZgl3JptRY1pRLGV94oAYLVratIAhIvfgbCq2rMQB6pJ0VWvqEpylJDI5ayM+8
ZtJVFGsFK8rgptBmuVospzZ4bUbv0zMZAp7SA++WlLOAs3zzIGObSHfnmpsjAVP3
0mEHHlOBD1hiJffwjnRHlEjsRrEjlg+cvlUmztopLNKVdcJt4Guw+z/ocBmONcPn
E9JbYdpoexd7rZiO3mPGO/Y8+1NIOJMQaYf+Elrrk2atTXqJTBZZmLyidE33yW1h
kst3U7Bv9Bjp/ZVhwLMGgYIMk9mh9znIiZyQZH0ZfA/obU75dO/hBCKrJEkWHOFD
GrOT7JOOl18Bf8O3cMn56jXzefz/EF1pHNMb3NdLfFGXz708IiM6+yildanMFiM2
kl1VesKzRgp7vb/K/A4vgE61pPrMkDklfpf2R4NHa6D8Tz7B4ngGbD7HjYVpuLpq
he+hvJozqCXuzqEsWpYClhCwzdfU8IjPAITHCqOyvjfTzzSywiuhoeQegNX/NPCU
x8XmUOjgunk+wD4sI5TKZNAr7PgJk04KE8xppMRin+DrBsGFsNOj4gUHl+T233Dh
uIfCpxgj45vEIJKYdt9rNEgOwwzuym2qLNLTQFqgxERjDZnYektrkS+bJkoaBUV3
ekG47zru/EqmddzpJgdqrbdVs8RxLd7ggH+IKSNrE1mvMzsTKExOP5Y3HLGjrBeQ
TF34sqXlM7/bQktnIdNAZeQDCJLVGrrMO+fINVBOUCngU7MKGnVsCHa8TY4xAXHt
A8KEBfi678ZwvWgumQtOxs2CMmsH58XWvovZ/KA30zooP4iJI4xDYehuSmwVQ/Q2
WazEpoOiZA5rDpfPw0mAzGdzurmo6sD0NUjmrh00LpDZ/MGn+g2WDyJ7TCpcfvXQ
V0LOQ+kuEB0/gK887M2UaV1FdiikF25UWKvHL6EeSyZd96TEQwilT0/P0M34mm5p
luzYORoh5ZgaxI3oOFcr8mJAww9/aQ6qqg/6kicPslpK39DUvICKEMYxM5JxIv9O
fCoq6pHJ3x+jcDJeprfPQSkjcmYQ+l/B4AC2P09A0EPM1lxybv5eXaJRO2zOFK9r
KHEkfkXa/t9k9HNmJekwmOSPdtHRug/K0CNKEWGaM/BZUIZUuRZFJ4ojDNnA7YEH
4cYk6P5kIDtjxlP+ztXyMHf7+Y+/cNZnbEedmx6J2ay/+QZ2XXVZjXgd1jFM5Ewh
4Whj8E90n/1youlh7jcCBxZffVypEY+GddG15MN3stTmmBlR5/vRcBOkE+fAo73L
KJvvFUI9i7vnxmoxwQBVycBlSVQI25WrgRkZJy71B2ipcPi5359S1723ZT5IYaf2
W5c+UIesHVquV2Xu5qALDFis6ntpM5GqvAvaCTsBzRY32dPeSUlO+wVEqUu2XYsg
dRNLcUU2w0IVWNz/M58+eq4UN0XhCpZ7MZQot7zebYNGZrO71VCxgPcNyGLU3epb
RHGcHWHh942vhmH5jNbJrwvx9z8suW/ki1qY6Ln7mrXF731SESMXchSq0+diqEY1
ch7VPu/ni7tJJkaJhTaMq68U88M+z4e56nh0a4sfArR8slguBsfwm2GaS5FncOYD
yrUKMWpR8nD6uu2yw8dd3BXnRq0vKZ8uq7NN8d6GXSBSnmq6w1D2yk5hjMUsLNSe
BYT8vU3cf3C7FYvay9eQOg52NXFvhg3UVFDaBqI3S4klXsRHNdiqgDO2s4DyuZIJ
WwQRA0vHiF2XR5R9g0YfS86L9neekijJ/gh8IouP7jdtIlD1lYoiqh8QfkhPGx+p
41RGcfIl+hdxR6weP5+Lmw2tiJ0uLpD/psiqY+6KPkX752z8GsUcnjqbyVwKYB8M
oAAOvIsZ3wvXw+t9JDpOkxoOgUHCt6Ym7hya0/tgG1PterPjJg5jW+CM4XDSQXDb
16g5eVzCxhS/Ig0NJvIk8Iw6KoY+FyWBRpJbXz/xhrsKlM5E8Dl120USM1QEQBe1
58iKLeEGluRtSi8dW73QCoHrF8l1+tGbj6OGTTsDfhlumohrgtfc9yzQN2C1o07d
IsqWY5NyqfYLQK6fusS0PKkfytoCn3hy3STDcvoJsRfZriN8fy4lmQSTz3BLO4un
vBQNtgTMxRLryawCgAjnBkMhwfKhtI8adUimU/rV0z+yn9q5fErXz6GjWqAZFnYp
GC1pDWWKoMUpPLSypuo+F7G8tyd1ccs5z7CTp9jrz+PUHzFnqYNb3CxOcGtmPjGA
h9jIodi7OTT1LP/9XbBdsN4hO/01mIThlQZCI2zdarD8L1bISDE/SCuadT0RC5oc
BFDHYXPAmLLtlkuQz+v6Sof6oxtzLa1qCqia5bL1Gsg4gXh3ntoEUYFK4IKJd1nz
5dy52Nr9vvKN1AO3bEHajWCSaKMLMWERzjkQ2yfJkQctf0AJX1utIehnQK0+Xu1p
0DV2Y0O1tC8nxVgsfbTC7i/+av0HZre0rtaGz5TitIeO3E8n7m857YLHaxmRmWxM
GTvK9TW86daAtogzwTrKqVCxyYRY7m1RaITPxP/nQHYCE7IATBThNrTkTlEHwm1K
rWF6Hf4kni+PVFhEBrHnUnjBeNCybNF1x4+ku2NZDl3I6C3K10FmjL78WA4PAffQ
ny1gs5MbBRyXjxP51xwnpvU2l8R8cdMqS0IodyUCzPgixus1Hatbtp0oQl9anWcS
YDCWf+KOwmKjBL9Hh/nRjachAKTFs0u6m6fU4SWz105soIEqFtEmyZ9ni6IygDo/
miU3XEgkaHQx1I2szK7/hoOP0FJSaUajOtVjF/0bECb+e7P6ZTq1mpTIKSXansI2
zcweuKcSWeX1pjZVT9ePJPibvLg153BWflUl+pcosipyYqT01mBaXjW220FSI+1j
SgYuyL/aWixXeRFqEyA++S3+991iSR/F+2pKA41/OitkgJH6+68GggnzMYAQdSj1
4ml62WiATmRXfud0Zoi9qqVEfLhSSQJoDNVteiVmqX4+opcqTqs8DFGM53ZuMsVZ
GTiMpyyAOS/iXocPLLAUciwGF6KknkSIMPGvEldao6z6Sde9qI2UAc4bHxyusYAP
6IEgAyLrIYwG3tDdF3x7QzQKnQ2Z1QS/3KzK+vFJUM11pQjs5Z5pUH7AJ9Gi2Vff
jLAtwYW23PYNC4Mi7U+c5CMZeUpQmGdV43AyUn5BY4i/E3fXxfBL8qmodH8bwSXN
C1AdMXnI6+SkjuL5cSKZyIZxkQt69iP0XiJNpgyEJFKdDBcQy93KIWDwBvBimuV/
I6cjQ6eKEV9iSVCjXDEehyEAIJ6hAbXsFC+URPnJ8f7KN/OSrzxoH4UufGnEIMEp
R4h3q2I6RO7yr2N7un28wqsiQRJHmk4jMs8vTQB2jyqq2bRvq3otoYctvDp5Q3RD
gTKyadXWSFrgfqZ3ZnFsRWXXu3UgygQ5eRAfK4yi1YKp0UDbBnn+PjDnJEwSGn8s
sfJXFH85FSBPpVXiHBnpEHMtn4lqhayPFfWXnUnm1NKpoifsCXJt0tvcKytCJyjV
Tu474nZMSbSXJT1btJucHnavLuHi/MFHzThoFZQdd67jaEYEgPlzjt4UQ4ubvtL4
wyI+bJ1AqlFI8qjmwk/bPICgqCWb+bOdkvp0XYTIsmmMeJa7rW4POprcglldiGu9
bUGpGAwpMcDuXffnc6Yat+djRHBnk+iPExHKnkWtgdowukpbvhIWnlxJ7je5Wn9T
/htpmufYj/Scj5v1ylBYkvj9177FODBtTeu7j+KGjfMjlSk6fK46yv7GncMLdTUs
qCYkSHdBl0tSMl7Qu1GrO35Rgs4HReehCv4W9yZrf16YwacygQoKupZkdVLZPsAy
y2EYXJDdphDaMd8ek0VQVPtmW7ZPrWJisUc6oaQRpdvHdC2zOJdDt6RgcaBFsVN4
7DktxFZm0+aJVKapa+zpTvWMY+cHPqtg19w2nTlfAZEtAv24jHr87AvGAZV5UITX
KoNoTZgxmnyMOp9WgXGuwLN3dxAEIQpZ8GWGL4kNaaBjMO5tKK8VGf+VWNNzjacZ
Zm3FvuUkdMaiTDRRj/qf7qrwBVP37ys+80nXINOI48g5aR56z/saIuff29diUGdi
citVmZYrD4BLch7hYV56QD6QcdFyNm5lDuJm+8ilTy062zQt9EZ1+jHoswIE8EHI
kf1V6KEUBLmXYkhk7OSEeYWAHVabAzhxou1e1IBVXeGF3CQNI/UE6u1qj3xRli9y
obCx218PrCVPJgz1x7yYAA+DzY30yNlYEmw+V39s0sGauDlfBxLZyWzvQBD8z5oS
HN/tj9mYJJh99yPmQ2gztXAsHwDUBFk8+egZDS51RJBzHISjDVqKfKvBhv6hxjgU
1XD1equKJhWOgEvaDSQ1kdXjHvdQ5+IhEJt3ZWAsqKmsVghvXAOBtMwxg4BRhyos
ySqaS5GVIyTAG36LiaSLxup0tut6NxWRM8vVrxGEJc0Iex/qrNinQZafqunlVI4w
guxUO1iICv6HaJKP7OffM67NSPO2DN1X/OIbCPr8XPMk2xeY9UjryqvWwUtJPXH+
m8of8/N6Fh1BPp5eA9sBb7j+tqt6bT8MHZTOCNNj6KUec8ZrhP5xfgrMRwpirOdk
dY6CVUHN4fN1pm7wS67zo+M5W+9vR5PM6JXiczl8+sr3+LHN6r5906UnBUeAWQby
mgF1oL5VAqCRNA8w6AH5+n9e/WFeFLRATHZIayurqrmfgAqmj3IznwHc9+I7EnAH
Nv4RWh7LUVO/Q60AHeVAqTg3tsUYu0oOg6C+CApmA/1Nnf2xm45jG1ITZlKnCqU2
Yab9ec70m8Tj9QbTQOGqbzvyyIxtRhNKC6lLPvOOo3+YGj/qmRiLB2x7TJJj/VvM
MIIvABUO4LFYMjRQohiumbh/87ASPqE7RLcwPk7i0Wu1MGzzdUCxYQF2SKratABT
2xajx3p9qvzv0iYlb6UWB6BFe0tdMFbCQ0uqU0Ftq2PaOvdtwtlSadLU1aoVFaZD
FYZhxvgUaYORdtQjbNIinHC+F5ns96O/39uif/fmS9zmag+0sR+fDl6I0WpdZ4rX
NE6L62rPWNRYpF0T6Sbo/fKvazblAgsaIfiAEPiNI+fyZNW3et82VqgauZLaVXba
TUjJzUb+aoiSNQz+3rNxHv7/sscJTraS+J4dYPF3sSQsDGAZacJsS1mhKzdZhdhD
UKeIo786UlHpMh9Yz/KgqScQUir/1caxKQyKC0wPkG/BV6O52icjIIRKXGr/4yb2
4UKxNTJPK+7NtXTW5UYPYdPu5SHfKvQc91M4sAzgFpOE+MZGoLqG14sEbMADnt64
6+8J08/dLDZgJbdphx9bGtIlzUMDTAUdh2rI8VVYkamO382TjDC5qIhLbSF/Da9E
pJdJr7/kC68Px9DWA5zGb78HRrTwihrz8XtmcakKrTle/91sNvTOju/LOrnb1+fl
vVrk+I92qnDOjLfu9b8yaTK7HjX9k1/920kOl60FDjzl+SUHzPTA2xUAMp/k8DrL
XlOKrJC0jsreYkveAg4SbzBcJWrqFK5a4wyXofn2x9F6yitpeugESFKcueKRSgBN
LjdhTqitahdMMMicYEgndQFqxbcujMvE8zdP5PhrZSaphnyCbQ/Csisg/WuY9zZd
lD8ExJtIX5g0bY+N3TbWf6AavFjwflobyS2mDOeNkif0fwKGVmDu7uP4A4Cz2NS/
uXZUkqDvid+3RDCJy8bRNy78RwbL2ttTPerbHWi+UfZ6ok7J3C6dhFgOZrnY1EUh
ObmBSbyClQ8fhclt3Dth1zCLJXtXSPEGvLX2PBLhImBqHIge6KtFejBlzzjc37hq
aEG/SbVqE8sh39pFVSYlobfqIynHs+f4w0n957h/Q3igjHwH4SSJGLIF3ObtupkB
HwAXT3gFOhdDijSBjda38AVHNMs7TZlWTkVfS8P1HuY2J20y71ZmUZM+ijr58R4O
eBlm/07P8rV8ml7vLC9Brv0agtgYBC/AoyLAKC5sb4eVD//JL8wv/3XjzgUwqkS4
bJGuMI1I59h2qMCHvA9lEP7HJjy5+Gk/+Y2oeoO4+2/lvCaDmcn8Z09wFX+jOXu8
e8YNH9nw5vDKZjE6wS+vDNBr5/aJ2LTuCNqqndz3CexdnIZbnn6DsJioE1OcN6UJ
6xwJzZLWhRZCnbLE7jMjtED7KdQV/KhR0fp7vfmctyLiBXAdF73Wc5S0QR08wwdy
P1IdSXiRj5TMTIM3IWgy2a9HIQyvaCwel5tYqdqQ44Y=
`protect END_PROTECTED
