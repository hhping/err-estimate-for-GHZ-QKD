`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2xs5nYnHLBG+QUP3YyCJE5HGwIPX8MPj5Xw0dcz7F4tVtiwU7kyw/0xlVJUYcPog
8j6kCAV5ozPF4IT4SWM5wIpn0r7I0dGjQk9BeRquh+/6QsEqyhX/fZjQZNO1JyeU
SpWoeym6FvBqd2mgR9o6leaxA6FaI8z2Mo2b4U19eTd45heb7BNpGgW5U4xwPMAZ
kH+nH9n3cF8oDHFD9tGq1efPKTPQ6olEMt9kFyw7xy75UVWXvxGtSNttNdQLE1lR
0oY5sDjBNaLmldNQ4cT4FrA4w5SM9c0Sf4h1S1vq2qZYqxXXJVKkcH+L21yF8V5H
VG37g7x5GjOHSjZMY2b6GyYxmWVJP9ptSPkSJUskSO0iQzUuDYG/wh7To0+MwCil
ZzI71vz5I9zJ+SlGDclJT08mUlyU+PDsnRKoX8hQc+sth+tcE2XpAP3ConWNYhuP
POvTA3hgQvtv//QSmOzBiyvA/ODS1LBF1N9tiVJFktgRSGIFjFRiSWFwYdy9t1LR
kAJBSo4EQzBr5PaLYNTdl420AbgX036fk7LTGum++q44poEtgHZGVhSjRF9OfblA
iZU1FpRrcZ58pnRXy+wbMzCZd8nPzaHzD+oeBfa5Kdxz7J7KsXFZvBhXYsrmUouH
Cdfl9HJdKy43H+hIKIJwrJpsAzq8lJBk+x0tSyH3Wjw21asdTn7V4/dCxgdXQrQy
Tcq/0RGnJKNzUEy12SUBcu4lr1QOW7leCoGdD1yXbYQ1+3X83AZNSKHqCV0u43rE
HuW+uy5bz5x2qKIqyivXEVK84N+Ma5sRHGMZpPEEhXdqHqYB+qd79hQN6IGZDE6U
0+AZFle3RuzgZqcNOXbVVwGRUjAQfO7h4iADA7xSSL6MHiM0Uc+EOHkPw8dKmwn5
zszOy/bQIhgIMEYdDJXQCksYp8czkFK3KVQ3PGcBVcKzPGNrvvZYDLsRdAo9NyBc
cvuWNDlmzbX5+wWUOagQiuDmjrtmFDd8CmHfsEXpZy66w4AMr8rJGB7cgu/JJqD4
jiO9hDyhR9OOXK5LhAp13A==
`protect END_PROTECTED
