`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8F8pCCUhZMjDbhxd8OIWTqJGQcie2aIYGG9PMcJdww2qmSU7IayQBasxvhLH1FHz
Us3siG9ckwf45iuCVuqyT7RcJ+XyUxLK2jX53yC/l/mrZuxj9q4oFASorxYBIvVk
HEEvyLkSEEa9cbQ+8A/IaEXWDlojRpd1xp0l5g+nv0LTqE0xFDyeKcOQys88IQuy
JkHXotXtyjhvX/2U9glAGxNZv8/CxitovEjiwK8KP/T8yjQg9fBODxoM2+q8f6IK
K1Rw8yLM3JoJQWfSp2jzVYZZXYslENdIdPJTmu6ERoXeUINf6TLr7b7VhxTg9/hK
Q8VEl58kviMpl+i5O+RYLsU0G996YkG0m4OomoOqmBeg1FAfEau1TanX8QZktF2o
tpGxfndI4nH7508V6MgJGpa5dcxBHaFExufn34t677G9NCYxyJONU1WRPUjYIvWF
TMyw+YvdwmQOJ67ZjJtIw/pHnzqvqjcB4JCafElTECRQ2jHS3Jqc3lMPQDpIrxce
BLXBT23/725KdMj3R14vXdHIBByL8jZrmQEHLtKfM1Q0bTyJpbOEtNUm3ujjHZIJ
HId++Gjw1HhAhA9DAB9yLbiOMbxuF7RrWGw0a0lDdq8wwD9/Z/xN/66o6bEb1vbV
sYjMcJx5Ja202fkj9+hk2yNeyef8Y4G9TVAqgwPGjCFpZKfUaTAw+X0iMF9icQcK
XHXh2WboOP6k+rCMjlRFpWAS3ESYUWw42dJrJfm9TOOrJcm6yHvlQR48ym7X4W9y
s9I+yTSfv+BDKVs2uDT6l9G7sG7Ql8QvZsP4UUCIF22sAUNLSa4pF6D+FKjapxET
UZezLsPjgsG02htoao8zW6H+a9SEs6FldZQ2YLWM/oywZEmLwnKtDMwto8Elk6sT
ejMvt6tcgglYeYE78GX/8rM4KuBSDiC+EZDfZultZ75SBb9JLhrE8leehy+/3hj9
jyc+N00AioOZl9c+iaMw5PXWD7IRVIfe3/IlwJWrFbI89u3TnLFg3dvVcq4Q7Hwp
3qyxCFw+SpRM9HqBeTMgiBdxot4doM/N1Ig//t15CqLZuVZH5jUB4f3nfP0obaZV
pedQEWcWQUFAxpskPb3bdTCNsquLdlKdHE2gdcsL3CejNAoOf5vr8ONVXwZpJUM/
616krPTDrqZdAci44Ov80RjOspfW2cxdYh1SL30lEf43NpTg1Vi02AR/SAYCq6SV
4PHJ/RZ4kI6alw+NGAECuLU0kNBBaBd44NZvsc2uZquInUymp952eXz52jzpLWxO
u6xpDBJdfKzR86Vu7NiBPfUSkGgoNMUZQeBnQ9RxlOtt90FviaaCM3f0neFWMCb+
bFy1B86lsMHaJIYjJ36h4AsSLWfmplyLTUDxDS3DEp+sgw47PgRN/zDQy1sEttyK
SXBxs3T1ZEyJudn+sWP6hz++3oKf2uBHmO/ziIPms3fDJ+8IXYjBEUwTfUfMRV2p
qgGJNBIrcWUoPN50nfF4FfQ68EYqrgy3RUPrHaok4eIgGRPUo03iuRZ9WSQ76qA4
+lGStUaNIehpX6Or21UIKTHG+b4C7Fsw2FPqMNbDE68P5xrIsZB+o7UoGDVNX46y
8/Fgy7RW+PWLxWUOgiXndCfh/PXSPQL8XPfl86SYpufMqrRBHj5QY1WQLhJ54Y9l
b5JEgmTjK6lLFn/v+Ty7Uoynq1R11vVbhLO6+752S1jzBZfHUDViQbyju5XaRPJ5
rysxZEvyopYJnZ+isyuZTLM1Cjf4iQERv3iTsP/6Z/a/J8mWMuuSW07GPNyIR4N0
SBZGoTyDTxFl+/S5uAB8u7nWfro/B2yBrYqrM5lJo6YSF+SWra2CVsMQQ1XBvhe4
WCpW277tgr8QtxtbBxzJZZRMwx6Mx226onShgGjV+MZtOAOELZHaB0jVJvHsT5iY
E3BvpjXlT4mBlCruWKiEQoNj4QT+uBGw11zfnWrPeMc=
`protect END_PROTECTED
