`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
voZ6o06Jf3kHGI6JGMT9cIQlkIupEZjhe23P4Gua9vbykJjxx2J/jBBsH4KzCU18
i/A9IwOEIO4620NmCMTdr7QBUKon5zcalC97hOeZd6wurgDFMorY7YSkSAz7gUuY
xx50JiWRb7EtcCkGAzO5I3o6C4fs0V2BnGC3JRqv6zG7VNbobM5EqjCf5m2VFpTh
8nVbT0k0avMw9NhwdJ1NiClm8b4xPWqqhCvUq9v6/D25XKpoUg3UNLj3sAB/55cV
bMO0ZzWEj5r5PZsux/IHbS0Qw/V9+6X8wCLuUTmcn0PSwt6zQxXNXmhtcqY7HhKj
Kb1UwOX9mBv6/ajb53fh5BP6d9esb0A+9xz3Nw7xhiAvrLph2Np/1yKGSKAzPpEI
oWS8FvX+wgQomflFwhtvbFt7Q5OOv7vphIBl6YSmEpDGI31K81uLt/y7Il6LPPnz
VXIlMlx4pBgKPzf4nB7P0tg6WqwqyJXsu+V/p30KjjPfUCDykBPi0fnerEYjrPaY
LSjyib1i2HB8lQd7tmmXXX3EVCe96usl/DxsUDPa6COMu/MkmdGSZKu0jgwy72lS
C6baAcvzDYOK6PVS2JIdY7Pank/PAjS+BqByGgjLWYC50mdoI4WGAhQ4EQxPZ6Nh
CiAzBtqavKokLjTTz13sC0ev8Rlt1pP3IVLx9Z7epYZBqCi3S1+0qL9ES3MIESSB
uAFvu2ZF+qLOQtDL8OTixgqHSvsxJAqYkQDiJsLGRVqXNoErMn0+VDZGUw+z7jA2
+OkJrIEpJd5BRRplpEIjSB0g4t+n02bQC9NyiOCHhl/D2d6CiJG96mJtakb8+0BD
Z/N0w9ztuE/ALy9mTgFov7sJgBo+ohcvPK8hKUW21Udzl6HnERLPSOePB+2fn1wU
DwNfAF+/Q/Aqnhx6v30LHHzwO9CTyTisc6sdXqDs5bemHAIMV2FxiuZXHoMMFmLs
u1tXLW+hJ78JT84YkwqTv8rAGNA4+BXgZ2RTK5Zj0+7Oj0z9tqf/NJqoAp/ld6U1
EaajQrq5SgdimeKrESeW9HrYZKRKfMGswc+wf1nFW+YMnm2irZCDyL8+78V9Jk7O
hTmnD4RkODQhEQZZLR2L0aRTMHFB+y6PvVECSlC//H2g9JBrg8JM/nVIDycqLbo6
rNjIwxwOSZTW3JwFJV6qAQoBwlmlBsXbU2NGRu/eAlfSeKPycHYtTxmJF6m0ONmf
MZ7cYhZ88VGVgVJRSIGkWQVTs2YbZxpiedso16uo8kphLcikz/0jlRif8s2d++t0
mBR+Uo3yi7b9fcRW/DwAtpKYz0/DB3nehnmmOKhOi41FTevFElzc8K67G5U6gUcI
4cD0lHaoO3N9YAkblY3mvKdRONnemllrv6xyRy3lv5I6LKSb3is2wECYXXnC68xh
bwHFoxBKZs1IR2jphj+15gPgD06mnVtGj8u05v/G7ANAES8qbUg9TTnKJJ5lnGCx
BnCMKkZyB8UuyvXi9gh5off0LYn6KcO4aYur634yOzayKQe2oOX8wH+PcVqRupCz
L2kfM8yrOIT6n3bcCkkIbOPaITsQNvqvIj8Ee2EPJ0wdeBjQr1DzJggVnJRLCQMY
T76zKSHyHT1dImpgW1tw/qJgbxxiv7rBD547ielwn+H9Urz+v1IPnWX/D3DOee+G
7lbXDepwQ6qml3zlBuzIMJ3SJvPWejtbZp+wEHc1g6er5aM9x9t6XSjdiCqIiqNc
c9sXImdsyJIXba3vT511wFDvAB4ESM28+OFO1h13qXTuhKSZAXkhl6GNb/evwMhO
k9O3hsfNWPI4QQoM9t0XbKnfvEHh252C5Gyw9xeduHOJzkutA8JTi3fL+9qR0zDa
RwfXe10dBb+QDh7MXLvCsJQ2pDy2s/jYLxuOId/9x1YxJuJoot2k0p8qN7EnKLZy
5soeTjSrbVAS5lM5B3AJdyODZl9YiWc+td21JlNIdJD+FtZThvidVLMrq7sdAx47
0GKnQO/hf8wBGKBycXIQf/hgBqrUCSnJLCpW+TpIEsJHvNVocPhreYl9s8+SvDoQ
DGrXVRUyCG0fstcoqObMVKs2D5KjtQHPzagzWbreHoFf1fAvVyaD6q2fykOs5sAb
D0Ssgn4A2RdyrEE5VCo2KUJCJiJYTE5Ll5kJQuQt0iFJFg3toKyxNlqPwgFu9xN9
9SDfW67duEho/q7Rw+4nd6KSLX+oeF8b6VDoNgiQUV4hqvuKvol5hEl7IyGf7BSi
EbKeZnOZycA4W9/JrhZT5uuSlXW+9uGwTlwuGJbxDiVSNwOMKI+zoqeoTolWYKQB
TomjdIWOYESqwbzuYl4hq1PXwyzTYWtiknPNBiZPEtytV2fVSJhOTETUybd6gUBb
KDuenDFJbAvBrg3w+5PkpgQRADgN7BKmyAQKqk25GNgebWpcM+kM+kuGY+jHLh/n
5PGgl/O6PdaaYTaDglBxv3Ykk9BAOhw2he2+uiWZkgkRbA6PGpzwuvOemJKj22PL
WwXj++5PlrHpk0crSLPr7P4B98U7/GvGmzmJCqGNhd4PdN13F/6wYtjLcy89gX9n
tp2HL7KPLc910uZau8XxOaIxHh4n4rpzHeX8rOoqCxEi/39mmNXkFYwv8slT8Qbd
M7mCr3mLtUQH23zOjT3FWthyeF75De2+CqCu04IGVrHm/IH1nDU/fvpC7PDItsaR
DhZF/X/qGmEK1KqaZV/1VjlHLkvKHYwQ40fmhrZGAPMu9M9VjpjdIHZ5Wi9m80VV
S3HJSVDC5IDi22ERaCUI8dBFWQBqAZjiPRzJ7NXTO+0kYBl0D2WVj+b9s/+izxHS
kPLra/KLhJp7C8aYj05mySsXGw5KagOr/2PcNV/d9jarIK3uJv7w/zviQyOj938n
suKFEE8ZjkPFCkByJAjHTuvmthTslD08X7qEXPzEgRHYnNxdSVbmAR1l6buehsXr
Qpe4w6d09IXPr15iR10Ge1yAv+dHGBiyUExkPAWP/U4Hrs6V+SsnrdLO4pZ6VAe0
uddhhEL3IiPp15aOBkcYFYRUjxn6RbVY+THFDPjfQuOGwz4IH1zjzsWs6fRyAvIH
e+FlEAyi37cMpE7CLb8Xyj8I22Xy7prsh7obV+QJ9yrIgpgCpBNOUMYNLbDAe6U8
yXD4UeqpRmey1U5PJZgfreClfdvI4D19wAoiUSc+h6ps/Jkf0MYrMTYi/8eR7AxM
wwMrYBeHu/s6Zb3tYlrhRH7u88v//Wb6+00NoIMbBTUUz0RS/joZNjFm5TKEr8vh
Hccis8cMLqDwtJ8wCJzjqEjC6RzxjFtvUgTLblKZiX2mYyRQd0eLCfYjjdCQbGhe
Wbu2NXMuvRnrNRbzwoslx7+A8BXVSU7/2gMQq7bdbCbqMbHUx0drUn8W3gxZNVUS
f43IndDg/v/e3+v8utkJ+za5B3wyh8vw/BqwQ9xfx3HEyCzanFwKSDBg//5kQdhZ
ZBSBrkdhDboFBcc5kTp85JLBIJY19z2zPCeqrkopMesRAycZGYkeqET4HWQbP3yJ
+PwKzE1nGSERATyLjFCQ7ZSvei3E0GMOwf0yTT4+rdSRFRi3ZyJxDXNNtbcn/LF1
ObeJDYRJQiQkaefvnEPEtlH7u8MBNWYVeqYtUN6xSAUoYWT9T/SoMI8l9UF9UaWw
lE0WagvgcixdW7L9W67e1CX8pn26HqFMJezEk/dRg2IIl98Zdtlqn2SLPQBVua0X
zi0m8hg2QyWhnF9PKW/CoZXUlRd5Zj57veDCQHI1OXk3JatP2uN+U332CidHy0tn
PW7BTpyTLbDRuEElKFbicT/olbHMqE4DxwDvqFoWQE+RHfZNgMJn+c4JAL9OqmCX
bf9fbQ90iqMLUfYIFLcixtxnniRY6+uhYrPIddukgWJC/w6Kg+SzP4YSs5HUxvrl
HRP/FQAoe2FOMpcV0+i7c1WD/hKKKuxKCafMzw9sSdZMWW9R2lYMphMT+hpnnqIp
k3954v6vKbncd9hiazuiEEUwTAwoT6cK2EJv2d/TTYY44b+oRtR11C5PF4Y4UU59
RjUfOOH+Xfn9CRdNC2ERGf9hgwNhAYaT3tS3b7xcuB65ZsUDfcXYwDCFX3LDmGvL
1T5Q213dRkKre70ILY2gdnyp2dj2nZhEUebFoYOp5jWnYDllhBfzMk5ydEXjZ7TO
DAsBCvnc3urPek+hC1UzO1Ou72QR8DoVHakM5lHXepHA9KEmtYnnPbzj9On4thDi
cqKii5VcsQtSSQToFHmbCNPQ3N7JbGs+jOe0UZ0ti0dNxaUWY8DLJKSVIrvEZSUz
yWoaaJgYcF6z/f8ihoRBpxoI//rDC5yj/Zu74Ub023qnAlC3Jm6Z5santuztA5s+
TOH6rmuhjEz4EiLToRAWm2E85pK4JrGqh0DOwTKDldEYfXiO86u/puwQBMXWxV0j
JXCkTPab1gmZMXhqcsNKczbhieWatvh89u+2NusDPaQVcqzGUvQmwZ0tGLHsYjnG
fJjaoMDpg/bmc6WDcCpHpPckDsBD7OaT1Lt9A/j1GZ1DJhsvU5+cmPDXZSEl98tT
57bp0wLifTdtwUcpRQYgncP/C7onJDOVwGToC4rcf8zTWFI6nlzNKBmDo+InuqZV
eJopF5bS+hGC3s3KwGbbT1e+yvsiCtMyUTaYr7H1Bk4LW1naRG+ASVPeyzdu9tff
zrrjtJM9micbtBxvNTRsiO6iRhQJAfW587pZYPTg018qABL0tN/nO93k0jEO6BF8
ctaHsNa5aM8iJWDRGDN8Jxuy4OInLpOeTlgtxnsqhAGaWi2NLEbsSGWOpCQCKj61
aeJ4neXt8QtTzDdgdN+dFQJHAkIeCgX2KTCxFXtQZFyUV3QSaPC0ARcbTuq8ybmR
qsdLgL+f5ykCWYvy6km29J7ya8rIMK+QFJaZblVGUQ2AD17F1zDoY9Ft0AzaOcEw
K1Ev4H9G4ProgQQHy9oNtjpfGrIH7rWAIjsVWToPaMRc4UiAkQz7TN2r4BmrtRmj
5/BIGLaf/FWTeWJaScmwJ9su8dDw3jTkFtQS2gYPod8gbKBFoL47eDligJQR3FFK
IRECxyH/7gUUUAvFA79UGJ2MzNMz0ESy0ormtpjSSnnVQCXfshifPIYlkOzMXSxE
uHkiTqw+z4dUAWUFK0+LbcJYAynEfwluyxIuq3kdkZApZOsPEWg1PoSGeaKZOGtR
0DbTTu7kUkRAcTNEjeTiWE/tedFrJsd7DVFbC9BLMLsoF7qZ2IbibQwBgcRXc+mG
IkTzZeKrqj/vZLps2mW7LcwwSWe3VcXGF2wuHaUUTZjhDI7ufK9MBkAS0pEY4+0g
A3RoHcxyDNVIh+8qnln5Q0N/t/2eef+Jb/f8nJnHgtVCY0FI9kJA+CfFT6YW5y5Q
t1QR+UVTxt42d0jFgDXnrOqm6dLVzcVujtBBrVAmJxQ+GJnVxSo9thV+Y7lw+Iyr
GjhTaEuYmqUR9dmwWfrH3iX6Em2Bc6iwrV6+/tI3rKV2G7/MbVybCl4AOpgX7rpZ
JsXbYVk+gPzJDXjxBz4+RNT+68iyhhM51S9ID6bbTmcXaTNYFAUHFv+izf9gpqWy
RZd7VSmzyPYnhQooc/lRnDwybRYS98JSbpW99IRmmNfA+nLAt/z+usggYH+5b0jF
JlKu7MpQJWSrWO/hDnlbJRI++tGwutC3QMAD8KdlSZaPbli1ORWq/BuDoo791fXy
EP7kvo+DCmebaJpQQuhyeAw1vZHYQNN56kcjfBbYMmJ3OqkaFpLaXtif4xkgXL0L
PxAmQktPHaJe5O6HUjVzqHzgzLxX1zrFFWZ5CpK2pXmKpeiHaIQQsYcyYji6chCz
nq9ji3CuTPHSNeJLzGC4GhOTUiCgwLdO+St69Mwkwoi2zkHqBAeSDBCC5X4wwEI4
NutydDvmhPsPbxcM8zdgS4LL7/LOABLTLYgInKQ72nTweKCIKfuPycxmJ84BXjJ6
ntKQtezDqRSx7tCud/xBefLIjLd0ujCGDG+C5tk27oJuMAI3Tmo90NE+PlPEQJYz
pCZQMuhhcIM+ND75uKLy+VkXxZMpuJ0TGdCfA2kxXcwv1DJzbSaRtTuOEcoVLGv3
MbLv6WEuXyUWZuuOIzpWrIvg5a5cm24LBegJHyZr7Ec4LygsW1B2SrNv16SMx0YA
Bq1QuiL9Dbe2G5yZjULNLLaeOQtWfwshSv9eE9tS850JwvumSHj8gm1zTSga4I9r
qUYkcOKdi39PNKWGADI/x09Da2KJXZpL6wB29/3FGG6oCu6rISTKSa4VnvSvCJ32
/8eNt/S1kZpnFBM8GBZqprohPyZ+ckO4DFVuqvN7bkKrUtWb+LKSE0mA8McrOtqK
ABMMMo5I/ZuPfO0Fk4I30v2Wsk2xJHG1gBHcMI8Iq/F9H6RcidVKRDqeowd1XH+b
poDc+XGuoWDfZWOp5tAPJywAi2Tmoj+//Bhgf9U26oFXJt/yPGdmXq8L93PhPnCA
vTQvwx6Xj6amSYuzzS84ckuR7a6mNQFG25QD1ScYPXRqPIW0dJNq8jACvauivCab
m+QOOeVU8zxso/EH/iaa9lDsWZt6vg3o1nG2JOsTKZt+6hRt5VS2h/NVevno6b9w
TslK4WCtlrPxFgz87H+Ze9q7axqbm/te+c2uTmATb0P4ahkBTDy3ZIQKGVv4odtv
lJDH2MGU4d0/0fhdiEwUbSlu2epeWE07trwwF9SFKdVc7OjwJcgyJas6Y0jWIYT2
KvlabwXknqJeptPa+BpWS+tdwg/eRRxVvPpMvFXfSrGdlwoVCPyIzNKKe8VaMLLk
HdWxBzfMi8EioYr/zEqtwMFR+aXN/oGC/ABkzSSZXRigknSpmFNdvRHbV4UMW4pd
Sx0kre7wPVeYWlCklW8JwOyf3e6TMKoNoc5pnhNJ9X0Q2RRkawxIcB76SVO67e2s
BebPf/CAkFRHg1heMpbD6/Gm4/03VDi9P0SjfPhTfjVdPjaSAWmn13YCY9Oft9/U
kKm11JwQpYWwdaOXfON3Wq29VN7T4LNX9rYoMxZajehT7mW65HsrvGkjJMCjvqkC
1Ka11+7LASnMM3B+ECPWSvBJhBYmHRBiUMweIpbcn7KPKyuR0+0TSNJGriZsdaL4
gZi3aXz2eiaanPX7Uk4IDMo8aSCh+Fi1UzGVOgda6z0FGpk3pdF3BVFI+YKM3Jjd
N+bHrVpbbTDbbLo+2ZmmGdVnSdajc3xCuvzK8ZJq80BPCXqijP3P+YfxF71QxYAn
Wz6aPqGqhi99peB0cuT+iudt+PsQScS+vOEaugv6MGNQbjn1YkmhRAaFeF3PCNar
JYDeJdxqthRPPDmoiOucOAaz7qeJyZZQV1Gt+yefsZSIYgSDgQxByrR57L3J6D2S
Fh4LpxNlklcnl3YcH4/LLTwxw/BtbUXauiRcPgv+LgURg2Xbj7fmAPfo/WiEg0LD
DQCmbFsrOJjmS8ZzKGDR4u7ZTUWD2kaaqbvhqSPGJhr0v+OZUFs5+zRgPwTefvxz
RFVzzmLqPFaMyn+/p0ePFRJzCUq8mt5s6aOqmVVqWLrlbPErsQOVSJFs78+U+VvV
7Off2b0XlOyKwovuU8y6nKwJPis8IO2io4vZG8pWjcYsTqS2gBDSQS1EQlv83Mw8
8euEIfcjrYefEDwy1hGjYhUkJqxvL1RhQX3RJK2WbMSlRlJtLkWJcYai7WVqszp2
Nhkwqkkab0bFodZKVUwM8TSJ+BMrkTg0x7IWc9hGZKzK5OtkyMSMJEKINthkTOcZ
eR/qxUN2oxBqrzkUGHtXquczzApFCO9EupAcLtP2zkUhqzl8omxGXlhErrkC7Vaz
saKz0ffeSe9WuMZKxPrz1OMp2obHza40lgIwJ7XBRrJNT4xgJ9mq+GMOLaiXkuZB
cPAJ/KXyHQJENRzqT4+kLmyFYAKgCkOp3+lZ9bW4sOCV9bDPIXJVWLUUUKLXfZ+K
1JnX+viL+hBSLX3MCzIxVR4oA5MAFJ7m9vrcp2ilFZt3oym3XCVdaJ4AOSqU92So
q+6FmPWvhJOJ36vQK20suo5iiHXTWmLWikDEEcaGHLsaCg3mrn0/B5Rb1ZcFLAs8
H1F8peIJhWRtPsdiEJxDvozrdfnKYPb9p2/LgP91so48cVBb7LW99Q+jEwLHZwBX
fntRrss58XVb4MKlVWjR3T8WQkeMl+3TRKM9c4E4mfuu1bgdsMmt3h0jESQ5ZAfx
4vA5QUyhf7QnK6TMvPsEiuuZlQWgnvmRkIB5cQF1i2Je3tNo+th9n8RHh3cnD4AI
x7wO94RlzdN0QL6ani0kJat9FWMG1fnitp5O1nL3a0cDIzNQj1cJan1S22Q+4Lvb
oljzr8JIfWdWR8vXhb3IXdvTeNrtpFF3Q2srk/6lPRfncsMxoM/+wZ+kRBS0UwZm
CX8ga7pLyIYwWtvYVtuLjzbQul5otqg6tvMbRLFZAgJLpEAp8bSrwT4PZ2UzivnH
BxMA5qza6ICNzOF8owDGDacVSDY+6o8a9YGR+jmebKNYM3q0iiNR1Y1mLJUE89C5
b+MREAK3oDwvG9IYXFt7bxZME9jLkUQYqXoUEC9i71pLdBGFgLn9VQh6P29KiN8G
q44MTj6czKQkRUkjekOHbBeH3rBR8VjfgAa7Bs9N6ghjoaREDpuGSPwLb/6rr4CM
0Ul981b7fXhiWXfWCt1nFF21v8tP8/1manlOU8gM4bwDhJAKpwNjd4npF+89HWON
q/ZFnjfaRyH9ccFEiWoX3ANs9M0eSQd0sIKfYfbo9AYQUO39aRikZXMpToDJXAjK
+j7liPBvbRILf3arTFoVNnLozp7QP7VCEHTspWrT7KxxXAl6J9bA6RINfdxKopPh
otUJanqmh0EuUQE/DHV7z8BAEdrX+ZiMMNp2I9cxistoK/yxLOKEa5/4rzAEivts
k0bSqXCYkbW4G/QHX4JsrUWJOzlKAp13AuqULCg2uBtC3f6eMCDXk1NK8zLqUm+C
DarHDdt1w5eZvm5sbnbkcEN8Jim6zt1doSmvJvggyfXsba8zZc35cTSlIS6f/0Cl
UL1WA8xQZnkmyiwl+BjT/ADoJrhSdiey020QyXg/Z/HQ2AoAMSUxO0S8nfymKExV
FWvScu8wtAVHFeUhLSTPmxtUQT2eiCihNaoppkR/qbW6uXxaeBOVWp9QHDF+bznX
cAipFYcReDyng0CX+YLJFOIkznPdh+FAbkFdUTxCOPJW8DyxFvgMLktcsdjn//d4
+kOITwV6j9RYa7O3jeTJjTr4fH1HIIGkbD0XsIXNvgwsBGWtJE84cQUy7YHdenGC
RlP9QljPWYBUwxFtRKmYDFmuoQ2r0qEEXusSFfsNB+aynqFPhzrXiSe+DMCFoAvZ
hTjq0kVdRJkUGbPN5qKaqUY+DEYV5aZZDbeaspxtiSrVbH/pjF6f/IhSNcKkQoZ1
HZhYdj7yP/H174qS30ERFLuHAIhAibVc/In9J5ir809KZF5FCaETfmLcEQ4TN7xh
sZkHc1M7Uogi7QHJtZuvR/qhMq9bDDVxU8zO50W9U9DDEnjtabs20IcmwUQ1xowm
rksFdokWLXFaqSs4byX3nrNYzLFWnmZiQEo880reyh/xhH8wXnlZYCY2hQ5YeFQ7
ilFoaTHurSSe4Moc+X7ZHm/fWe1u9v9OaeRYxXlKHQZausbqmUx6mn4cb6qy8YKB
rLB+DFWT1OJTEOfOntLoMKDXqzubyNOjJsbTKp/8oZMzH0AwI/sYwYUsLBqI+6hK
S9PC0X/RiX350yDylSOCjmJyYepMZmHnGL4+aS51HpdS6mCy1ZYFuhNlqSFdj/kI
lso+bTmjudW0yKcXp9LYnECdK0yBR3ooNUrRWV+R1D8ccQvqv/8a3sjeZ0auFcpn
+gR3W5cd+6Ustfy0odIrR8JAsW+fU5AmwwloGUdJr+t01S4jXjku1R+uaxWUo1n1
epAYqXyW1VMU27qPVg3ASHbWFHgvv5v4odD4EteIa44KoEiCd8jK1mZZN4eIteZV
iNxVtqAEeLzlaPOLFukGD8gWUjB2fzjH7ljjMWQALHdZ4ZpekthCCuUHVUJXLMje
b06j7RJbYJ6rwS6+rFxgoLng1jgBEeAgTFUeMoWHR169R3BfdVHAsbuN8PrxmPyU
fU0cz0p53rdIF6jRTCiNwkOxMjlFr+fxkGU2jbnVK+n5/4x63Cai+lHI/Nx+TR8r
OMCxF/t71Il3PFsIP4UCK6MtkxAI6EuRmcQFZJymxHPMRuP8mvF9LEjqq9sSyTX8
PSlUY6IOjFgvhitwdiTeZd6hFLeJ6VGkCo+TLjR8kMwsE/BgPEREhIsxgkBMnAAe
kpcJ1O+KRwyijL4yajhVvQQoIC+t6s+jhAbHXLVaUou4SPxg3PTp0mjuSyYeRVN0
JmoEEJ41W203ypHBlOq4+QED7r/AWwuXKs/QCZJ+1sNlcgVtHz1avHBR03iJv/DW
ULp4HTiTH6R/4yykrbmrmgdPaGgMEIPd1gziQ9TLPb40ytAxI75A08zsRzBnsekP
QSwJAZHPIQWNkSEji4vH/SRNth1pp7/vdsuVmWI4kRQk3r7E3dxKG/pZPbrfnSi9
Duvk5+e4Vns3BH6HM/BaFDlhLdPkEuxmHnqcrX5QAiW2ecpdr37oTHKdbHY6RU2I
LM9CzuBNN8hxRuSB951T62IMEJQSuzMYT8ioBlu11iZ+6hLNVv7fJ7oEZZk1+yKU
ByvoyDOF/1qwZkxVfBchS2/ABWAdiwPJ7hnQIxvc/5lLUgm2CgrSOCCo4i7BKuqk
mLX1JomE5bXSQ2uBwc9KpSkj43frtA2Jv/o5YlnYkyMDF8JMTSo31X4aFB+LRrRT
iPdyB21KtDHr9Vx2x3xYRI7QO6bvnqpwHhwyJLAq9D5ipbhtxwE4+IKtpgBIbMTq
7gmzl9P4aAyAb++HcH4VTvd4sJ20ADyc+mrmBDeu8kvt/qDQ2ySkXagznHKHHGcR
UYdmS6pfT3soMMw4WbIjuOpiezM6xsTj/iZzzXJr0l+jhDr1MmH+BnY+g472JFpt
quG8rAjyMyrhDmj7/qjqHoY56I/sDrFk8KseAxE9Rx6kkHMqTTsPCz4b/hRSDEL9
cxxm3gGpS8AyeSzCcZBG/R3HAgVS1LVZr/SodIQJatDxp3UNUqwVKqcy7ZAwg1sb
iy5w9ZmBeZrIZ3V5k6vXBFkUs22OHiQnEFPcG5XlAOKcZmzX5JLf/061zvLhrG0v
YKru8zvZVRAu3enqbdS/lLHq1D+DqM8q4OQ9b9m8NJ0mHUVsqh9kfuQxJ8sBQbzn
RgMpKGSWxC472Y8V1D9QHOjsZVxB9Ko9OnozToRHHita+91AHMcey4JZdgbqocmt
KWVx4PMOQfnTpUA3cFdK6PQ8qw+6OsTUq+7S3ec8ZdKjaqtJjll4fBAZLosM5H9g
E96vlo8QWFjypB5LjVIGaK4dOuosfij1j8GvOSATTDqIb+dbhPfH+4iDOf+C07J6
GbxbzWTn0c4Yizh+U7tTsyC5sAofNVgdHQUv6eipj68lrPB22CK+Nl1OixdQ97sJ
1CQDqlJ+KGFXml0nbeieGfaLS2dd2l8Uzi1ygFRY1aoXBqYodzW4IU1RQckR44Ft
5wTAorfT25mZu0XgUktIbbGfgqIy7ds7//Ni93q5+nNXWKxYqAP+8+IB2k1ajTQw
0CMQQzhMWhoQKXUToaq0oooh+R9vhM798R02Bi8OTG6bfZajmUB+MwsNK2CUwS7i
5FQg7clj509GNvynmbpfwT0cTB5hjafItVrUGh3GaRYlYuB0oU7S7kZMybkLYukd
P2Qadcxo3u2TX1mciWvXFv6VXwJMzTaIXd0KVl1rix20xnq6/Uq8wMzQa529f6bO
vmjKRLW/F3EcugukB5SNbaTS7plQYCqUr/qa7FVWruZZopt9dquSGXJ+w4YjuIOk
zgyyUDovc5IE/T6LObDfjTkQwoK1gFhj2Cgsd+GbcFApClZQ/dK+byji+lxbubd1
wwfz0G++8UzBHx7Q1a0IKwdSbAgCTB0PFc5bs8NO34R1kTNkzGiHSNYMlJBZbBRr
icKmnUxXzW856/CKlPo+1UFfS6Hkc7SY2bbq7Wfx+7KMdEclXzhfUTZCDE5Ru1w/
w0i+bt8bcM2/LVLOp436uZI8upm+7KvuNt8ZIIwA/0RK8b9aFmnYM6iPxT8X8Pga
eFTItWK5AKDtF7BMBwSerTmJdNCvknNgLGhqNeb6q9KmOHaznXRLb0J3Iim7TNRF
+IsZPeLD3AHVtJelJoSS4hoO2kEMagBMnhfamlE1GePXfYn2/UrKSrNUfaASMJGa
Hkp5AWj3If5K69BJ7+ibEDfbK51+755LKpKJ9ILzekhVGhKYAmoT/7WBfToUlR7C
Ouur+vk8E8KMdMcK19s/UARqqkQRc7QhGwcR141hJAiB06QpGyQtGSmauI09yDQm
XUD8R6HmVInLBPYcp1YcB1RGo4z29g8BATOKTfDxYGUbXJh7cQOStfySpo2LAiWa
fO73EZ0QBmJyP/vms5IsbYJRjvYUEmbhBKnEKcCkznBMgZWOpk5gYe0XOwqHUIP5
oEXB4KayzqKTY0a4q29cIwM8TFaoYjlODsjfm2xI0DSN2CISF4OthjSnHH1HfEQN
g97PjRaQ+Wjp30JkVX2hMPwZckyDH6fbk2aT0uO8g1tRVkJTFTcpQMWzQhyHzlX6
I4B8NW+O1Den1XozV176sr2hygSW45EGKox9pVoIsSzekWYKXy4vZtbfF4OOgR/z
8DBjsnlSxNdap6Jif5Ld8htJdvjTiumLXgDe/aSAlJ0/bwXSZio8UhVKP9nF7n9U
tYVgMOnh1QPLSXszHb+i/e/nlbjcgJU0EJe6JzejysvP31kUtD7aVd3itVCiarJz
CF8y+9I5VxXbkRerunhB75Ye11MTJFD1xsiT7gl3lNTP+3df2OgSwXLbMEA1L+tf
hcQuhhhv7JFU04GIkY/J5hNoPEG4zR54NLpQhaAFvmHmuH7c6JW1g75G+HJrMFlr
0T4nEphgMfN/b9edOnWq9ERAstYA7h3cVbnxBsDPFwEAJA1K8ajNYgFrTA9I/T1R
uLienJa8wROR0bMiA1eA5EjAGuR3iscMQNNlsJTaxTgm5jl3L5rPfNqEAzytt3BK
gtKMfTRNkeg8PrMd9tqmR+80JU8oTnIxmTlK07I3eWQO0RsnC8jaKCSI0ez2sWtU
JiqbdmHFKyGdEHJggPG3SZJVNZcY8XFOJD/vyU+epX6HOBIz34L+a3J0mDUMCIPF
mXB8fx2MffBmzmDWSz+dyFrYeezWxJawx7Hauym17pAdYyfbDyaeWQSM2NLPh8rZ
QhcpJd6l8iubBSIZz1dQ9gmMCoyG1N3RBs3ai5jy2WMJwwwuDPkbWl9xIHRBvHO+
+yR+hjl0Hb5OQwKIZ+4o9fl6J9rP94tRjRtY3c44aPyVqFA5B6KcWy66FwXi5JIj
eiTHfy7aaxadPl4B8+/Dd5Ew6EOis6IIkvy6aDliW/90Akkz743FYHvjxo3goUwT
1+0loPjYiZISTLrppl4C3I8HdzmsvNTVA5LnBehO8c9jbj3N+/0CJd/1NwyN+hmr
sAHIv60AO9H7kp2y6DkpyQS02dGq9jXBV0+uYqeFUWu3Ohxk/3n8zjzOO1vfR1Jm
rkLgfmHQe1b39hr3F0lYFNfV17pl0wB4xf9mIdJd7tSGM2y//Hi3v1KY/u2iSTXY
23a0BeSrX5YzSmSXqtY4VgykBA14DkFZZ8ETIPZtDw4vkkE3gNi2LHMdTACAildI
VhChLGGOo4Zr4n10f4vPUXn3/Ml8jdPRJf7pAL70q6Zsg1PfNGdqb2l3WUCjMmwU
55dlaMe9qddazK39P8V3bvcbBj9cryB9M+bfyfWD3DdVFwS294FmY2DU7PKaEeOp
1Tq5PRN7deLYuyaXaTZ2ObS2Cx1imIYXFW9FHQSCn1KgIZaHYpZxB/8fIRGCWUWu
s6Jhaw5jR8aHFaLyxSKDsiApLm+oL5HZOdFZdHTwwb7oEbrxnpMJGwxfkZiDVIUd
0DJyTvdShmIBKHf1eWIJq2Ob8TDffoEjfEQCO+h+jEq3jdsTn6RAAPTG8T62POGv
GsUE8VhZ5Bw5i4jv++dVK48Nd43p1D5MlRyOw3DkO4kpIEB3aaQCIT6e3f2tz2Ks
gHGa3V4ieUIPwRGlGFHBe3/d7UJRPE/3I/lM/CKUzlJyWGs/B6I2mMo2QVhVIOhi
7b5x/XSfi7AYjKV9ST4l2UF76PY1m9cd54AGbmPCEVmiJucfzzPgIIOWoNAFeAko
4i6YDReGKFKcAiWgPrHEs7bpT+sDDLCvjUnrDzv8/NI+qIq7YP9nRHIEJ47uqJmS
iqjwsw03KFs/qnXxWmY3mAmEyppUtq3doIFKYVI0fHwDAyOqym36pD+IFTxOpOBX
z8VUEJ3X450dM4WHLWXlwVvIpX0Tmoi+Lta809UPqgljEhdMKN7PgoeT0/GtXF8B
Qj4fwB/aafh1C3iwUPv+UJDHnh9Yfg5P8NxAPsTW6rwDvhmm9CaiAEDbeyZsv9kV
hlcvKnEKBq1AgHjhNTTBnN+mvRUk2+O0tnztHffqlh/F9Wsf7b6lUettMRAdZInd
pA4dMQMlZj5qXAJWjdCpkBVPmh/UYFqiunXeuBgEILmKJjNwWne3FUodYzHbBF4k
enreB1mhw65v0AC7Xky+n69mUUNrNGu0ARpWuyzVK+TdgWHAQRJAKukC5pP5BJmc
74UTFNJfk9R150j0kx8wkmACgL6fM+JW9BQszssNsQS1ako+xpV7XkNPTD5r2AWM
uc8WLUpYFQ533+F5uLvFel4bbR2tPo4Q2qdk7WklB1AjODKD92wBwtoY7g5nb0/5
419AGk9YtTU+O71/UPD1oV3D7VumnCAkt1lYHL+6siM+Mz26wKXRLRs+klbTc0ov
xBnxKGfepy+E1afsAT9fwJapJNPw8GN0M0TXWYvFkXwZTSqnjROYq8WaGuGLd0XP
ISy/RAAHWIVDuzZmTC+ZmO7V/Rf7k06/D/tuAtzvtP2MBiBmbYs3JHiCc3KEIRCj
SfdOn+gJ2zyIOgjppl16JcJuFp4IvSIxVh0fCT5TgmSLUFJG/Fc9pYGiDGFhyZAE
/mgBxULS69lGmWHcAmQN5WzvRxtnr/Mxy4TWEtEzJrg6HiQuvDov1cnb+iq/+DVb
Nwlteyd56QHa4xQLWwDIoxgnVp5S0xON3+B9oD9zdnelQi4r0dlfnnDHtwPE1P0i
FCVp7HepzVzYuLGDHySesz0wM5f/jVxaEjp6FQHNJdii8axFZBt/MRaUvkVtPHVO
C+gv/dHzid4d3GdvtJAZELWSQZhet8XdzxmlMq8WByigF/oLGsNVyOinBAgr00NT
eqeqrm9wPqxuvnuw5tIlhQ+sMqLj0Rmx1tHhQg1cAHjUJ/GzA6te9o2qlDnZ9UcN
wOVvAETxUs2+l8abpNISWqXCcmHM/Jgz90PB2VkGqz3laMmjRm6WE5yhaHICxhSo
eiEwrWPK1IrRAdwNBfI5Yir+TRVpC1qbbgzr+H3HShfCyxNykmP4DqrBda2bf90J
N3PBlQoslOjGx0ZPKlm3MH/Zm3HWr/mxGgkiiZFIJ8jHrx/K5azbAeCNPCp0epb+
MMmbqmM/g5iF694juGBC8Gy64kumlwkzp1lSQxv+kpPL34qh+4xIosmlG+f6QQBZ
I1/NEPkUYIx4G67Zdi/f2eDDWDGSJAAeUHwHaMYQxC1MS/rfetXxfJbCKtunoyLd
Yir7lp+TK7mSYrliUxvY30UybzD9GXZYVa6zg4bdO/8=
`protect END_PROTECTED
