`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QMvFPyoC/26ZuN+IeI76C94bylFTFlIXxP+2MFUCR8MoxbD2MPN01biyKo3/NJtR
wlaX4prvq5gLDd7OA88PqTNQbwXtE4fdE5nmE1YyGg0zYhPh5ShTsgQb/sUXWcRX
iEmDyqZ2aSQTmSDttpx5jqGbB6jPyMqot9vWRyQo2Gf1EIgoH5Qr3G9dOK5CUbYQ
Pgaz+XyErjmXSVj4hynRt6GDyaQv3JHfXJyxOCsRz9exocJKUt6bDiegTwzXhsKf
c50Xhe/9q2Bw+4j+Osr9IpkgeZllgubj07mK0CfXq3QIOs03t14cOjr8tMR/Z7Ks
RcRQ6hmxR/jf2773azeT4kpZM0lO6pRiCFg5t3/GEO/PIHupY/9jO761j8XDzi2t
`protect END_PROTECTED
