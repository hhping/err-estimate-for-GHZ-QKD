`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XRtYpTp+xFwruO8cBvsBLIQbK5Pp7YVnfajd/7HhnFjOhIwVXzdCyfwcpTZTPIsP
5yRy8GwU+c41m5c6F11CdX0Ilac1pSsnCt4ujQO0IPOC06zUVn6geBOo0SXcDMp7
EpW0KF+q2I51JE9OveAeRweBXNQnS/4iLDLIIzBUowxvN1xcsTFlE+09comRpYHt
Br7MFYI/ZNJjrKXtc3H7a14Raf1cdyLMSN75q/7Q0oXrLE/rHuu6kYEbJZIRRw+c
idPLgm8mgLNxaImzbsLOrgPClaABwiEMNlDFvm8qim/aWyt4dzyBKKFM8QmMA41p
s2YkCUzE/kvb5tc6REM5mpwclMMKuSnq7aWe16H/I9mlF4e9AEZf7u7tDKTJy2Qs
RS43QpM8OnplFzDh/o/dzqSiaRYQWuwo+nj+RjM1wcCpI+eSfIr+vnc0sQMGsoSp
3JelqJGocSF35ip91UggKkFXgZBJ2rb57mZWr4lLHJfUWfaOhujirWHLvqNbo5FR
yt+aq5Vcszo6dTLf1D31Bh/fMxFdf9gSRJSoAk3yvqI9MDS/WHWnrk9V8oMsazcU
4FYslM88a68V+46dY92xaAUQjwic9QbHLR+KU7Ix8w2eA2NYhxcnZsICqtVqAAq6
CEVQIuCUNzRXHQVBZe7avlBxOVoScJLne5Gghelo+xoxXlFh47iWHx6sRecrLm3x
7Fk33PRXezGE/y69oapX2madDzHQ2vZT1In0I6JROmfIWWvwDRm6M1OoIdEnH0Fb
`protect END_PROTECTED
