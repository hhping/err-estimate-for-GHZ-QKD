`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rWMS9BvuAuaG57vqh2d5VF7+HlX+1JYGJWUDknZsSNANtInOeWTBvnRL7cRn34nb
QpdfOOsmWdKGDPZNAnIllPhn6nBC00AdYkOLJj3V6l3onj8Lov3eTja/YfyibKpI
5Fq44mRSmlaSWaVoVL75PiNdf/kBNjSS2qhMP7MCBiWbho4jnyZhBIr84yuOpmSt
UC1fvaKnrDhOEz2BayRB0sCwCXfAroAILaDmo7JUuYVULpdCbIZS2VzsgtKDx1s2
WD6jCx4J1GNIXptHy0X+EQKkZcP9rd23o0z+GkUzSMLRiWE4wami8i+JZo1h8OSk
Y0SQl/6X0sFaEKfkMB9/vksiexwB4TXOv2qTrgG7cZl95FzoL5DTVG884LYex5AT
2jQ6e7RqHa3rNfH1xQ3acQIe1ITLE7gaq5Wztzh/OtIuVzGhzEt0iZexf+Ob1Dja
CZnN9jxH4iryNBqtXhe752aowxWo3WPEpeTX6/EZvTbGYYA8qcNH9ZKhp8drVpNk
NPXrv+dYY9IrBWXeWwFC+zUiRWLrDQahvtvHT/kHKmS2nBcAdV2VYrEbuBLp11xv
wQcW0YmS6G1FGHdyB7tKVIRm52QVIXYNo7NlK3HIsrNswhMF7/iVBWtkwGHTewxd
JomYv02UMfwm+ZKEdNfJ0CZH5cNsqGQ4PaLblXK2ODvJCT6nljI0ujzHC3C2HxsS
T5gA46/iIzWraeP259HuIM9HEgym7nofqFvFTO5voMyneg92sVae2wHwyEQ4xoAx
acEcbWGBHJExvXjhYYo5s+pWCcKMYkX1+YZDg6DwAIdVhgWl3LQI03uLj0R2eU2a
95/pOYyX9bJn6Z1YuZ/irrzwZIdiN4QmetCdKSVbtz/vzGEC37ijvIh19pcv0RtZ
lt8pa4XP+mrB30JJZnXRpqe9ZPy9QFKbqbrARZ21EvLgEVG66FtGVEMG/jv4Fo/I
cJP9Gk8PLt1OtBrbH1hlwbwCsF5V3dKjRe+lAcYfPeAIZIN3TCzjwjRpzvfQLHRZ
GxXB+8hpy9r7oN2e3xm/lFKSg3spadH6aY99DHA7o+bAKGP6yPRRsLQ5xZf0Yyoe
8VrRiB5ftGDNtMz8PO1P+mO0YIy6wkgg0qrKzjHfoJMabw6NajExnF3TtaJO6rWm
Qq8TEcxJgQ4ubmzDv9MLL590jZkLixlSaTV8tcy0AIiCI7f7nPdD0HfVsNMvUsue
7+w3PRBwgLRlOiD2wwMt7AkEdmR4d7QofMqjn/MXe27/t3WLQCaBV/V+Scdr6bUj
+qvGPcV6Za0OigVyEkdpTqQDhpweSE51Q/GJPGS681YzqGz5lE9cFGWb+4vth1VV
833qqK5QYB8aPgkg/FxAm8Sl5x72hdNIHp6wNfr/5k74Rt4u/fGshjv0bIJaqUDA
tDRyE3qvpsjTm/3sxgVVAcogEANHaKebKdo942j959WwtaWaJtFiyQOXD37ZIV4N
GLTgIs2YN21/D3rAo9ekNw2wzO4V0DoekEKDCZGYm9RE88H2d8c6/ZL55rYK8s+e
GuCXJpGJ23mMk+rXewWZMUcD+0t2wVe2NBXXizBdyV8HqvlgszVd++pB8TFQagkz
SvyOSKE4LosSvAyrNRBh3mMDuqLwB7nwmRUQeoSofWrpiEWXFNv9PxRWSIsheUb/
vByGJYpDhV3ilKrp5hJ9Fm6ZfjwmGJbrE9Q2DfC9VbkKNpR0yPJNX/IkFUk2QfOv
PAlZ2l3DOf3jgbssopkijIiLUzjmtyEQmet6d9/2W7vbmrq3c/prBHlwsFAuUNRe
7+8IBcrqDJHIIg9Q+CtM+8wRY/uML4DrJhbtFeUOLEuDT4X3SxNLkiaOA/zitBae
KaH1uVgiwt4KIRGboiYNIrszAIt/aRXwtGAeqqxeo8A/rN4QMUG6hIdd+htK24TE
2rI4Z881r6CWfT96YiE3oCjMHfCNOyaufK3T5iVHjF/T9/vT6NoCzdzKagWMpJWR
3tJfvUsIMIwTp17QO4Un+cgu3OJxgx9fcxKK11DX/ziuz1oeoD9BMaToaj4ZqdF0
IuIJbcKVXeN//SxVDLi/rsBb/uxOCdp8wG2uARHr5SaVHuzywm/M0aZQP/esuigY
RN95g3jnHYY3IG8LzEQwmmkZ+hYOj0A4uu+Asl/fiThUgy2OA0JHNL5Y3uMUfyv+
jM/6wFCpRZ7pmxO3Qf1DZ2uMyMavTOGmw9bGuHL/rAV9k/4VJpC0JMZ1CEE9l88U
LFK425Nq7oIoAbdL58salcDmHVlA4BJImjFCIUTzX54o4y1swRHH4qlUZqGcJqlj
ythgM8djYeVenhmPCG5w8LZALLAurqMEAqgP713jeHgbXUJpei/AvSbWQrT1m65f
RgvOFsqfNheEPqiqriSBDSCU5SUY7STyRXDTdHbO2AMtB2oR4H+5ptBKPbY9w0uE
KxxNxTmr+tSLFpNR5Ho25+X8nTe82b+pWGJk9tiJEYqeSK70WLMEBNTdiaMmUUHM
hWwX12ppgT4gC6mBVWidY+lijdq1WxnLL0z6bclkC1ga4ZUEcW6o6XFkICb/VBEC
wbIyE6ExFRcmT68iwlQJH3hY25AdSUwZBwhyQ/RceTNL0nUxPcvZuDEYEBRuDA4d
AIckf21lSfaRetxFY3MCq+KLlDPxNIroNrCMPOJOWOkuhayKeCrSvXueTUHvosoz
ZSD/LDvMgMrituoAhe14BGK+WI2pxDorI+sciMoS4MgKoi7RNQmRU2A4gNp4jDqb
C7JG8fluzn8u8jRwSvcdjWPYjg795WBcdJbRUMli6DY+qvHEQVdUPwkgP0FupFpF
TIflOEp7oKj4iMZ0kd1+qg1c+eRGLEabFwd4+Bna1P1KbGDWktz6MZ1MqkG1bVie
3Utpq7gd6GxwOttaa4plsCokjX3Sp0Z4AvRmS7i/lBziH3OE6alDt/2Z2FCZ6sQQ
mhVrxD8xUe4hQOm/56jnlY2jEBemA3/YKNZFmA15QjnBrdZI73cb9YMB7n+nEJNh
EhRoiPm//t4yLNKKEDIF2LSr+4Ko87sXjabtMRsatIB9MqrEUjwgMZgAWY4FHbcx
2NUTDUEjVgBlEQXIEmHgltY/B6glHIKEMhNdAAvzVr2kLu5zWoxfXGDVx9flRtBP
YmXG6YPMZtygL8ulqjV0QC90exPJF0U0AZavmpI+Xcdd5ozmIrJuEYaYNqoDHXoE
ev5wx0eNkRgkmqNk1Z1rRgbrvHOG7HcmdwitaPCF7v8vuzWWbVzO4RY7y0thEmmN
8pS05URf5d2NGkDSyX54c8WE3hoAhAk+GSRfS636QFxJ47VQ+YEyqdrjNrlXco3Q
kDkLD3q7u6u2qWFnE70puM11QgJ+AP2BatNcQ50LXK6+iFr2y+pX2HummM176ztM
+W3vbZnRSPpG8kQPQw2FlxYaOOyMaCz9Evbnb89b7VIDbD2bqb6D02IigLXXfYub
ill2UIVEkrRMHAtqoBNHFtJmfqjyBSKLjWYOyQzNCPAiqV12e57o7SCsbkLXKX7T
/y/6rFwcS/nmcHvYutzvTUCXt5wMN20tDiAmBhwMZGPh1U41xd1QuC1Amo9DPVXe
LtAjPkN4MGy6A+3jJQwoWIPms7IqzwK5ezYspOhFglXasc6ceuFwpDf5SzW4JiDA
kuNPJ0uZxpwSi8H65M+Oj8+0zbDLSbUvB9AD9t/NdUwTzchhwlalAtUFB2xKSBJB
irngLro8OFOomm/bVavkmI9LoXiV+dBep7TkRGyyGM7PIJ7TxNxgYWN2nRzJuGTd
wa2/VeRjonBrwzLjaZAi728ViTu5HB3VJ0FeF5IW9bKyap1opENTO1B9NeGebH/9
3sr4vpK/0e/ELzdYhg+DXQGNQsXWFgl4yaap3kISkNSUfPAAHRr4DeQ3jnu3fmUG
h2F+XEOjbdV2opqR/rGy9+Igo32RYGGRN8aGSWD05Ywc6vqUKdyAbo99WuUaLwwM
wO/iL383U6rgPT9dPNyY2JR3lEU5FnkpBCiHMRzJ1TLzRAGGlNjDI+1k/JBgLPij
hm/5TpNyIuQ3r+QUQCHmCn/jm76OBm5TplVeStXkYJzfiDxo634fha4DvjPnTgeW
AUaG79bMxySSCBxqdrw9Nh+4LGczGn99GE2joqij09bqIZYkQ2M5cIqdnC2fX6xC
nz96Hkf2Ls4qJB1bHMoAhLNuhv/o+5UTF5vnLmg9jRb845GZrnhJEs077CwpyqfX
ED6B9ZCnOxVICv1FiycbHhMTnuDxbbDfJnmP0hC43AIq+3xW410Y5REEl38nUVCr
UMo/IEACFcp+BnXwq8atX1hgxgUo4rYckHnEojQdqaHEeF8d6U8rQzvKDg4Sqz1w
bIky/XJU0bnLUpmmH8BmLvbpz2mncaS2U+xvdlcd3JnojypRM/C8S7P4GN+JIeGG
BKTbbiEXL/fFgItjHvTipxIA4qUjgs2KCXbMevmaYPkODTbnr3cSRLp3UCDyC+ZV
fCuG5r0TSuYtvnq/1D2/TKQg+IiHKCn9rUf7pczKooZU7dMLq89swxdwz3VqjopG
hN5nMISsq1LRlUkW8ygj8U04KCYjsOjJcGF5WswqDwk3iBKelCyrvvpEothytfyE
g2xSrtq5gi/FerZzC7Hf6mc5T+eMnmlZX65sSjGI71qIkfrlRwrJazZMU0bTCIL0
eLqIqXrHULt/3G8TGWyOP+iGfGF+KzyNvEGBFviNKD5JAxwo98eDyAEXvXzZV0jy
77vUfmeDSmZlA82DjHXdU2al9KqlZLWHlgyWGaN159ejX3y2B/LwcXQT61iDiS0j
aKq5BJwNlF7RQyKqwVznc0xOnIuqXu6mX71wCregAI8eENuxt1RGCIL+/K5gFolj
8P1E/ghK/XaKShWOiQek1G/bDU5u90ONknZ43pDnNJe2vpDF6V0ED4K2yvCDrdBa
mg9Y+iSNRrLENSAfUvdJQadvgPRXCq9XYnMCgTAvsWIkBDkvs8HImIuu/Js2r7uy
PZjZBqD2Ek8hKXH2CwBoqP5MLrnGiuYJ/IGba2QKch92DZJHXM67TYkvr960PXvE
jHBWurKosCKB3GeCO5JeN2Hlrw8uVGwviiDyV1AXfFViJEzNukYNfAPXZViltfeT
xKg7tB5al9/95mmXka7AQp+adC6DHDvlrZg2104Sx6vH36pBlSfJn91tX5rQLgfz
ri5tnv0aNhhOw7bbPL/vYEyflrgklrS9IhjdJKvy5Fxop8D0xDHYphUNrTL5WxZe
64DqkSUMPpPo7JFqdO79K9gSjFNvUl6P5YhMVHe+yRX9YYWVOYvdUUnrQMyCPR1n
VL80k/0LYsHDWbzZHzyaybG1rkJ0UPONXV9RkefcxKN7XV49Oeni0+uKwTGkLorK
/HH/pDW/u5rIMUL1cXsU9N6x0RF6QoLyOYskHXejILh5GVTM/DaJtED0DmEvLwfH
oI9+GzK3hBDSq/1eaJRzqiMCw4UJu3c1Nfm0j2gNqZ2i9D5an210nHVbZspk2iJN
Y8qQ8wpo+uTq0wT7v+G91WGBEf0ROTg8uktjGYvon00dLPxAT3Xm1bjU0ZmKa6cS
ly/kw6/EKKG15rLLYhDVpu1sG2XeQU32jaPKo5OFph6OF2hJsCy+QfP/Crga63DY
GEAQQBCno0RYzP29pz98vEfcv4GnXRd0dN8yYIwXfXgH8+8R4ax0woJG9nj3zG4b
lvfn3V7T0WUdjHtX12W9AiGe0IAG7NtZtdvpJOHEvpu9NXrDLdjVSc/KqUyOT6PW
d8ClgH0bK80csMNndQlSiy9cy+hihlJUd5uwfDqCc3dIBURgxTL7BmX/GXDIqQ9J
qkd/tmxaZHQK2/2JeyYJpudsiP4WM5gwUJfQLe/qhh8sSVTYRKKQD0fHxKtJSrU9
cnqnAiT+JH4OVLuGhURb4V7StqMU4zqvmPiRcomjjjyUG5Gp/r6xqqth/QpUl1PX
rTQaC9UeWAlI0+8dgbPAZwDC9hW79GK9UGgA1yYX9aYjcVo//TsWuq1NGuMpdr8a
0H6anYdXhqtEFw9raqfQHcDuOkMtCEYZxNrll3MeMrZTAOqCs8t1guhn0Cc5HdES
P6E97/9asWlt8xuqrBk68tVLrh1c1id7QJH+1xFQgv8sw6AXnlaonKGqtgVInBpx
TDqx47dePKhkIuj+sh0JLliqPM9zpEVZYSkUnm127HTWgGhzumlDZB+q/5vTpF/J
xbcjywYgn1tfQooDm++SJL/lbzHyX3pfSK3BI0fozIKjB9xfR5FcaXrVuw1Zr9u2
sZbu+c7+pBskiEs+TNpa5NDADdvo/fhf3CxDkc4Eiyxkh78EFYxpHXKX7AWRfOfJ
PaJz0/jkCJAycXqdGv771mc4zuZd8KO62MhgE+A5khhUXANvdDaHIR25Fk16lAKb
P1SvQaosVXmU1j/C439shiW95wQWk6noOs8YsUzTPtty2NL05c83oV9QHHmiZpnq
dqsqMX5EGfJZ1E56DYYH74VP5dhJPLHNB/4aaPs+L+OwV/6j83CueQb2ikmyIj4O
ubXHL83ONBL4/qwUpkF7tzyR5DfbrJoNAsZY5TvGk0rUqy4g6JyHgQta6/2+7SWT
63P2xOEi/GciyaAQbrEDOV5qjqxkdxf1Gzs6sDfVEXIAQJc6wE0NIArvp5E0Q125
vEpKOGgwNi/PSOzdgiJ+wysu1bFBk+7bogfTvf3WhrX8nRI07xNZQ7/RZDpN6axC
sWo2mzcTp1h6CrFPWdf8GhwUt4DAcoqXEbveNkuj46NmrStdRBUUWOMchUcWKw2w
QjTz64LvLwcKILuHC6GWTfYvFcOL9wwi0zRNiCzTlQK7JfmlxslJgDaSFh3bzonR
ODJnm1Fc0vmb06WxeB/NsHTxZs0blNK3vofSU1NDQ0E9IujDkYKCEeM8WCCrxgtf
nq2/upAPPYEzPotFq122h809CgQrYtPqFQjtjP4bZxuiidS2r54LTZsyEc7OgP5N
kADykfGjACzJ9mPpNRLawvDb5Sfdq3lriWAVawnx8ygWdoontegaIAC5Tbetd2+z
ptxlHzNd5U2WQ9XrILOOjg+xSeSlfJhcugLZlhgTSE7x9xfxDBgMNW59zQB/zUdP
X7IROxDOt5WC2/NgM6K8P6TtOp1HUEgwEJ2McGpuZxhZyE65fDZa4Xbq02g1EPY/
N1YiE+4w0NpC+ePPf3ZkeVFUxX46Gv+Gjll/1c9Ef0c3P7hEILpFc2Lm9vrwjDHu
0v5u1zpRGf0zFqdvwMjH6WN3CJHwNMYX5nazCIAq7kz5trhTduHEjAZ4jhIndPVL
9wl84uxITDBc+lF25WXHAx5PR3EVozcukV5Shqg4TKD58TZleIFuxaxGtOkxM/17
3yh347lddTICrzPHneOckACxIgPU+xo/J4hvIic/qBRQIONNwsmJ8goGz7aHu858
mBG8/PdplLcVs9WAzgsWOz5KREs8Dx75wfmkgTxBrA9FGw2N3CMWdYgF61pXfoSg
hnUUaYqIhlls2qnLs47BfB/xgo2ZcY044uxrVAYD6rAC4XSHALugz1SRLEvr0WIL
5gY8F3f18VVmmCtNvOVxS1HSF7iciXPjopzSQ0pFatViJpb3qh1ENhsVBXsg6gUE
Gnkc6KEY4O/43m1YajL0VDEuGUb5LGZQ7/iZM9Dhdqn7jyD0sK4UQdeP/8mfZXIq
FwgWO19FO0j/DgCqFsHjS4PVpGlz3fm+BqUbR7sooUhtCoQkP33NtM2bcsiJgG/J
AK4tcLik8ifbAQvjP2Mv3wjikDOTP/ipBQJKFT8R/s/Y6EaWJOPafnLI3iNcy6wx
GvGIB6lO8TiTej6JRNCgBZmOQCSq2YTcxTkN6J9o2sKRLGAmqX82gNLa0MibKJwP
yw+V5u7uXIJxhfdLW1kbRgZHoUsNgrN2NWYQFdZIFEeV0/CrNcC9Kh78jO4qTHeI
/ZkeIoI+Tmz/ZqEFYinaN+gUyz646+0isIi96Pu1yShghk8mWoElp+ltbhaRILNj
tqbglQDwtNIoVTzq6o+I3o8sEtzpcMU4bI3ww6vBElQHnT70NrY9d1s8YrawKZZl
AItAO0NRB7E8/3TVD/IQubDR9tbaCA0mhFw86PfhQ7iibr7SdyBX7UytHKHqPaiK
pqnjtVeCRD3t0jNwwC89iQMbnNI+RQTVCBksy6dVnG0K8Kj9t1tgNObRY6UAPHjn
WQlcYdHozVYzTAeHZlwdEKEfu1puATBPZVa0a9aeVt4v6BqF3trslXZmFv42WSvN
tPuwjEzrXfKN7oUquUQWbouk/K0U7W9vdRC61xR7CgLWasSTCp1Ooe3+GvM+bNOG
82dNKpdH9hoOw6aajy4Yslb9Y4bE2AkcxOCYkosEis4KKZGMDqCVJ037wkcqnXcP
EUc5T5pH+zHmASgALbZq6M45J68EgUL7i4JtZ0F/yl+v9KpQrzBu73Hhmd7BA7d8
vwmD4PJfSA+jP5FESxTSTr+9P9wVHA+zTxOHYHyErEHOHtZfrwCMaaYcm3Ei+Iik
F8MSe6y0ZyzCaWrcZSl4f8EHZqNV1PL2Pr5yPKSrjRzkLD8jcVGtjhLHQOLNkQqH
DJMCK3reu+CpO5TuNQpsNv1uNEUndKvaJaCOlSLhqX3O6meA2OYUXUxprPGURcPZ
fPbdzeh5flWc0isjXdmf/h+NTMq/AvvtO/LolfTT/1AzXc6CqL8rOVSRjV3rnmn6
t54bLYsUI6KPxapg1AGROgXofEe4qZVF8YHRmZ5dtfRGZGkJkVXzQYa5YeUSAbeU
bLp9H52xkoEYaTvXor3K5y0MTJDusphJS5SCAuaGjDv8etRaqKtGXqklVorLYE6F
dbRH9C903PCFTx9Mo6rUSK0C03WjT6Ud6SFAp8YOBmeTr1PX1QRpdEPxP7tUj3pk
G5EXymr8l+cn72RUHG+tuyVPdTdIrny6gTOubBK01wVYS3TZ5k/OX70OFd07qrzs
nmWOjgR6833fvQnX4FwVYLmwgt8jJ6+8hCALuLaTyCg9vYtJOnrb2rxaZCUxsQf0
+zjxL3xPL08F9DT6M2GaXaCmGjOx5KQLTMJtTpUEGZAmFwuLb75BQN3VpoguWMJb
a7vsEKbsNY2PTgC8m6bSkFJj0nMUGptjfCrbW2rOl1PxplJZikxW4jxu0TLl/btr
qnIKqMdBoVcJwq3TLWLd+tjU6A5OLVORVRPtrExhXnK3j5Y9fSSqi/qc7bEWq/yv
ISnvA66+WmrHOQnO7JHbWzg+H3kO1PV84WNI0s3/4sr+uqJWVN1jv6WbD3UriTXO
kJ+aZOKdOhrWwGELq8ASbv1oSrCRTeLL4M7juPLgVuaxHQNhwm/Bs8jzfC8YXh4a
wjkgkmmD5pPDtrUI7+JOEZZEMPQGiQU5uSuutg5d0LwbSMuII6qNoHJlsb1cCZso
+lvzhrP2H3H0tSL64KVYo6ebGWYxiHa2RWQr1kDe2YBaTVOkfoItR4+5ETVuQZUB
5bPVN5RaBqbOPCtHp4mBDVYY1X1brsK1ciiyu0sOVF+VLT3a2VeTnaHO40cWTACN
7I81sSNkb7nRbBolLWOW1GJ/36JRBzzFowuFOEwCvckAswAP/salmdcBCn/2UDRn
XPtfgbNvtow6OXCi0zJWquvR5UmtGgrHn75+71BlLYEtW37BnVlolQ5+025AGnxO
ObdMy+cqk+/ZpU2ANqFzZwQ1YmHfvBdlA51LEoc3BxrsIn8tEr2V84J5AS0HILHg
oFoH0mweH8u9aEDMOXreaJab+57xk2STc3ruHJR/BwtPHNA1tiP5SlDCkMjh3K7/
W5SqARTLkkAZk06jpwySCD1YFMT08q4PzNSLNgmAWJxFtohdfZ7cy695EDhRAC0D
W17DIMhmI5ErDIIAxQECJ9yJeoQdvZRdBrf4Fla1aRCCW/NQFSRQdyfi6ierQUHk
n1XS88FcexnwyovIRtpwM5lauoHILgzAUEqd514HsKQYj0u7yS5aBk6pakSPAvV/
L9L6Cinz4WAxuho7dBcfMuCw6a5/kR5ciRv+Oi8qFPlurRuSYiWHrPOFemA3Ein0
lNy2orUMbXf2h4K5XD1jBbxTyjxsSB6+blV044wSJXI7Wp/2n4khTB6fn2fV5s9a
Nj6FPPxdpZjyDfYEX+vJzhCBbRlgDUrTtdfybRQFYoqvuX3I1Pqbp0fQZkQep1W9
7DuLxgxy9+SU1Mqvk9L7Bh4F7ZUHClUb6o6STQo2TxmkranwGboS4cdzQEw6SGpZ
jIawEaQrwp7N59ecwAoFye36Evrm/7GDWF3ioRomOOeLcsbdvYAUIneLjpj49iq6
JRXZ3EZ9dtb51cm54OeedVse8kxvzVMneUbVk5IPR7wO/B8D6psNS0BQILsuUN3B
m4SN2TGPZ9yzjhD2yHKw19ui15uUgWqhWj/ncsrbwrpXaGODVymyYMfkZ9rEAkb+
GWNadWM7pgMR9shs8KvY/ink3MmTm5GIdN7DeHA0BqmxTyMDeEWLXOAKZDpyd+mG
ER5dTtUdb5dXcZ0FKB9/KiyddwjGdJdGE4SC/fzZG1VxQTgm4SOBduCa8lwmPaew
Mzz4IJ2hDaDSp0+ZiGyaVMxgUh6arqsm+fV7yjOvAQ/DxNrWJ1eOfY5D1tWuIL3m
FzKZ63p/oI+gMN9gQRqlTHTCPGshYiNnqtKJoonPWz/7iiYF9czLlvpA1VoK+/fn
2HSOSJz1fSk7Af4/X+UEsAVIg9TfO846/o3MQ8nwad6SSFdlFLzlkXo3rIVKV/oz
WRYb4jz+TILj7vEyfDOxnb6tWJRmXw2CedbXn9xosY4JYHzqQcvBCmgkeSvkZfoj
lHdrGNILYA/3iVRqOuQ20uL4ZxKglb5Ne3Uytd6dJfXxYYdYtDFDtkzKRzSJ3aLi
fFfQRAPYU48VudKBqGJnfibixWTFuOLP/2dLDSQBuCN8dIXrjDOvVNxrBXuPUyyq
dDwcg6IWSuVzjgBGPX4bp2OnSDhB8S1183gFURLT9lFrkY8jRXlIp9pdhTPotIdy
NOVsRswh6mGqE64K+2S0DsZmzHaSLa4IItcCizQYh0Go++YmtH6pJ1LQNgtgLmXj
BkDHqCojroEe4zCqxDzA6AxDpBJPG6Bf+6HH4xgmOQqysExku9Igo0lMJWw9fh58
nWPqyAH0pwrWP/LjlmBUUu7iIE1ZtwzuEbJzwr8XcSirGtRiuGQ3dGR2JGDqiV0W
2NNk8dQnuRcE91YpprIXpA3TuDVOWOiu1Ee3+ckm+kUQovNIqBsDBT5MpAs2ZDW4
QA2IYeMlI5UAIza3rnL1xZBxGs5C6GemPElIIJ9a9y9QD/eX4WM2Nt8muElI2siN
Hvc6mgx2beOxHr/e695tM0DlnAFYOhDpU4Y5/QQifc/3I3VishWUk4eXsTKWsMZh
XAU3weZABvlIAuweWRfE1+Z4Nt1b7SbJHsS1niUmNnnqeShYNdHNryYC+9OzUXmX
46nviepLgmr2OdMfwbYlo5Ilbx0OZEMnB/yZeA1ChCIz10dbbNGiyDvp/IcAPWsH
Y0JOuNfNKeytvVBiIqNL0+wkQxVEF3R6yFvr6uQJyDi/WDz7jNFIkoGBbCPY7XXi
ov1TRW3DF6FL3IQPF6S5jbcvmDKcShI7HCrgXCp/A13Py0/i4jI51txIcd+Syvyq
NiUipmKe6T1vwc1sKMk3nY51FjuW5l38P51px8FYGVooG9VMl8ZWcZ9iJOkrc7X/
6y9F6yi+Zt6nu++wyI8d9pjUZoPvztmclM1CQQVE3/ym75FfOpCafohLzitsOHia
e3XYZK+TBlyu1tQNggGNFFvbXtwflv+GpXl7PHiSCkKkID5B/JDZrrm4EwbDmRjJ
luUgb037anhD0jtWso5MyO4PjK5uERDVdiBiNJzGfzyeyzzYSNBZZ9BKU5EycPa6
FR7G6qMp214+7ujdtlEwO0fOTjK/tLG3SjWbPCUTkz+9PdpbSICowwD6EnfnLiiT
n8DElts/SMv8aFVux3ul2eTuDf+1fY+Lr9Tgp9+WvYLOHKDlL0kSAoOLWqkxzkld
03yE/ErhDLzt7l400kHWrEDk8K5eLLUVeh+evoykd1YWPHEKrJtd2OPu49PhH3wo
nkGB9cAuDR/azl8jn9QfvHD7glU/uvuQQngw4SEb5JKAPzpQZ0v+x4UD4NkSiqxx
7sWniba8vit2Ldn6+VGPKiE01sIQH/mD8n0qiVt9NwFqmouqPaQ0QKDiey4xUbZb
ji+TES0VRWP4KLVmV3m5pegqTVAjEbqZWC1ABkpzKotPkNOEBP+Er7K9j1g7lWtl
iBGD1/fS5c0XhWMCCV1oOlbO2PZ1gwZ83Kvw2RAEOlTRCHfHXAb1EDcU0Q3hwM6n
dYeu2AyFXDxfoDk1G9VpI1jE4N9vIMZAUk629J3qMN6fGWQ4jREsjZZlRnQcChrE
Kloj/TuMXAgIsrxOjSB3bMiyPckXwz6xq9eUG5CiM/dZIw8+qiTNoTogjDfL+KW6
ho38A5I1keglPq+xPElNDlb5TL/QD2S2caONOXD9F29pw4crfQ7ta6DkJUWRX2Ji
oPRCI3WX85D+UV720toTWq4pl5VjmGBht4Eogeyde72X9aK0s4s8CKP7WIIDXLRL
I4jUGuqa7f3CkM8e2NiB1/VcztBpFnVdOl7XOoJiL/aq17qIRVvVQV734n7zdJrj
uciCB1vj+dZ+SUAodSu6grqFgEcoQsRZ3WKH1BU0zvdrdmk8XAZrh9tXqZyHhvRJ
z66Ifi9Ib/+GcaLiPVHe7OCtTnY7L1Akow7vzvfzwzo8SsL60gVEgUSi8m8YNQAn
MUmP/UsHsRnKKokSM/gjyq+amLNsb33o4WQ0m0GiqhkCEQREswzEYnbjib9xeSVP
CTo0ZzcT8pASXV4Bjyp6rMnuzcsBqYUazc9KNWkgCDbJ5wnHpziMh3IkJ2bWt9XT
EfBKhqbduVg39e8k11ozSU90Mj3G6Vajwv8/LY3TIL0v5+Y/nqrGGgZ1WnIUvMnc
0MdnK2PKhCtPuscazdqQ6YOxb3yenhfh3QGTA6K0cZgW76OMOpvJMkXix7sBeBYV
Kcs45kR+UHnMcq6A0brnW78j/LTSskZAZ0KD6myL50GSTZp2tlv5OU93sy3s7iNW
UVpohmMQSxXn9NGX2+Ms9l/44826AJEz4LkGTVV82GlMxBnD6nXGnMmTIcIwHTV2
W4il+zQtPOB/wepjDWlrTMddX2778NHLJMW52WjwODeVyVGhUiGVv2zvoFXkS5yv
+2/1iFeYaxBnTgmjEJ/NWP7d7zECjikHBdgSxg9PpsWR3RQrY7Syc65f62578N/N
Ee5PRc4nFQFK8vips6V2Ld5y51ZfEK+SU1uqo3NGsES6lB4bEqjach4UTbePNIMX
FdfBK4+Jkug+6xWfwo8AxP/V5gigM8Gz1oWOZPedfLTlb4IiPB2hAGJZcGKFcQ5t
rhVAAZ7B3HWdghF32mse+chUq55KXKBCN2svCXktXEX+/8sj06mKpQRobxBm6iUN
mK0uHfaff5JAcNODUX9+FJPk2kN+DPfm4nz8coKmT6ct9NFC25VHYxXHN/nLIm8H
4ZvnM9DGW8NRKxnq8/YHUS+AhL/v+M94S3OYf7ffFB+N59ETOm7qqYC9GisIrUnv
GYi8J1Y8F+E+jLBtrr+XvOvzpaMPkgDzvAszqXkQpn++2CqEkrhQuRTtfuRfEZ2b
U/amM1bs8Javksgyz7smnIC7RkyiP71vQvx6uSP6TIoKBo3kBpO0BZQPcWvpr1re
rQNJ0f2hr1BAMb2ginduVQCeMAwSO58VxvOZgpyt+EGQUbdIGKob8xiWtb2hVkCa
aJVYhQCzDSrWJ+HlS5yPZ3vJ8t2N5pgAJFE+QZf7awFagGcJk5rXcVz3hGXoYe97
JN4ZUcIncGBHqNJXO+/EoACBJRueJYPS9n3DRuRtcwmS4wq72H+1iHAdpIXt/rKx
ZfdShleJxN65rzXFCICuOzBSeMmF8A0aUTId3MvlGSgyoyrpfhAxYVV/Cd0ddvSH
i8EPiSeKi5G03aHWmWCnpz7PEYjord6REksAJ2OPuqz7j5kvZikusV//yH3OA+NP
miXrYHbB+Dy1O32dni/JjpTd1fqWpz4hhdFwBh3gjCyf1jC+iiZU5jNAgBkDtnbk
mcxKbn5sELRjuFfQ8P2qKaDIZB57OaG7Ayrwva8hpgrCS4FWpinS5L4ZNJT9hU5z
IUXLRVEDzpwRA5C7BA46sY6KJNOEggcd4Hu5vsNHDUVkTVUwZWLZcxIBZHczcVTy
wZPEURGHLwu9DZhzNId1xoARV84XX7KtpP+9hvr+wxBemqb2Cam3oFQIv9epZvII
NTTKaz+TH6lr9lYeMP8Gh+QFqt/lQM2Er8ba2+kVeXByHyMnvymCqStPX8/6TxEl
FAmpuLhGKIGAX2kPe4LtiYV3bZA0CvoeQRom7caraBM5VoWBqN/pCYSx6dIZYq55
tRaYA95eqYwg6QCN3ltZh2UhBeA7eqZYX1NJ7aHMboPnDcJYDE1B+Cdhln7Eq1cR
ZPMTnxb0GEuiGz1l/USwynk0O2p9K2RX/Qt3OTWS0vyFOg+e++/PKP+zEKwZeKI7
/98/FDxNICtVfgMzAMFYEsB/leYCp/N9r8NPo18Gv589VStmhHQnIJUr+GLOX3Fq
13hGdAoPkJRb2IzqQujMEgs2Q6ttVYxW2PARcMC92v9HzJef73WTaMAzUZwdsHGh
r40dAYLojwlp/a3LybUx/JkxphhbmLdZDV63mTD4bEIdSOyEYc/xFYxVIw8kYgGS
CCApwFTNRu+sSsMa4wyxgax9qQwnDmlG/ToPeqwR9JBCD8reCxa2gyKPLEtESw9x
`protect END_PROTECTED
