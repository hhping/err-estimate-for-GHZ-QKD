`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QvbOeCYV49vU5DetRCoBT4BIcRsHhWmzpQdqBbpke9yHnv6S+Y+Jf0fKtwsbURNA
jdFE5sgotL2Hbc9Q3dQm3kBbGpezk3YbAorY8c7gq0okH5C9ki+v44ijsAxxGLTk
7SKjtORiQqm9NyCVbHZiTgRuOwHZaXCuVX3a1G4YlXLjosOGCDhRnpboAy9JGETZ
lb/okllT1wYzPs2ymoj/EgdsXNy9W14fKfhAknpIpszP0J7WPJCnt2uZB+yVXak3
JqcDnjZ6lz4RzTEMrqJg9KkGkPyTuHug4gSsjbLJQvxrymdTjL/ZB8AZhSF1hJwb
QK2ZFltIUer79zo0CxPpV/m1L1FVKOHeNo+kk1j4LkUsJoZnzcq3w1jkDEZFzCRV
cgzcX8zjCY3xkScn29DBreIxH5unScBGAgM9J2Nr4bwZGK8JLOD9Qe/7X2JwRfAI
dUKi2huQyzK0jLh8x3vIbDz0882YJLwa++R38jo5agmT0f1uXXQq4AZC6bv324Ul
i4+Q+XknMNG18CTz89v4F7HPMVqjpnPZc6I/PFNIO8SCNB+irDOFu9/qU5UCRHBe
SuDqRgAhpAckzDFk9Lqb5RRl3gTD0QbB7cUQTOeS3bWAagis8ERzZLnto2cjGQej
xVc2KkZj2AacuS0hJos9nzcC+1WVS01CzzX+gQMLIQ+IOTdqW6XXZacsHdEfYBqL
I860DUpcB/dzdbas/hOXXbrHlvQdwWR6yvqwUxRV1sCEP6xzSFQP0+FdFdm8eO7q
02tGZbVlDoaBGwc8z9w4wNdwYVO6Qxjr0Etu7aL3OSUA+vkpj3IKsvmVUFt3YTf2
K/OXhWj+Asb2GCVmcAMMO4VuxguGNLp6M8OGziTFQRg7hHfzXAmvjWB+S5J7Ag1l
9YzDQzqT4vCRRYmneSTkpg/sWd8CqwInEGgD7BCs0tnPu3QTRt4A//PFJiniN3xD
VeMnc0dGxIK16vX4foeSN4vsDtdkLAEpqgVSWV5w2Nngy6oJaFZAqB40yUCBv14b
zLz+SM7mmtQ/e5IWPFrrmeFq71KlaStjdEH6nNW3m1uB2lNqkp/SS7hheG3W+mhX
iagrYSnQUZfbb3hy8b7muyVrkQVow6/qoCCg/y3QP/05ahNK05D8JxdGMeHnAneM
qeCgfDDfsGItbI/52+JhhBmWf4BTG1B+jgKsK9DVWXV5XMRU3swfD0G0ktXGXBSQ
zx1lbDtF1RIPdNZoZ4qX4GFiHu+1qdEaLh9LWwQFj3Xy0tvLUg4BZm8rBtnfubUY
5ROskYxfT9QqDQjJHUVtj1rOQMdaTgN01pX6JMXNP8Li9bwngOkOWzZsmn000ug1
3Non2xoFtYnIxhhjo1x09dzHbfNpJf9yv2Q8lEw4pjBasjm6FWmzuz17Wp7Br83E
61XUfEYjsDC4klJ+haeaLdSodx/ElquOMmQVOONw3m8KhGg9YTWJR7Gw65ndus4/
eh7Ipm/OCn0h+dkmVE+t+TwXd9YA5/Mo/va2GXEAWSrGOXEfwh+76s4vofABYnJX
LHhm4/kBJvE0FMhIQVuzRgilhQVqtt3OFZ51C7sjTG4=
`protect END_PROTECTED
