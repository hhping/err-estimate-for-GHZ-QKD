`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SPSdgVDPFCaItS1E1Ri9XyZ8v+6TEHHvViuW625N9lWAQKQV0B4Q1RV1qu3VROHK
NeNDM37IsUxQJoxmGmRTggMtO3STxOf+RRs0Lp2jUJBwKmYtMbpXr+OGBcwPyJpY
b2X3upuqNs2upmT5C9HCnPzv1iAUZ+QncdIY9xp5AFUxvat5T7qkNpdhuZIhF88o
YnyJIFJaex24ZZYhciuHOAlBtuTibpR0u+RFepqT/r9we9uXj74C7x7qb1qsEucT
6Xts+UGpCuim/UhmxifFPxDA8RE/4TUKmgsBJBkOfTogVNFRPll2+s11ftSyEBRe
W7UnZZarGfZPKP+3nlIlWXRSjxO7NBvgLtKcogGCy9K3Na5Qu+ZR5NULc19L3T1N
pqb83ZrnZqEptAvy46xynjBd2Mu5JtB+qNOWSa6kWsEE6W+jJyojTJoHw9gfGLex
enmcu6H+9PUZcqUtH3/7VnTQv5Wq0PJYi/tDdNWLbF8QEH/rplM+Mibc28tKw8GU
k+E9oKsI/AGodAQfLFBGLL4wMN/LHXms/uojjZijMS7R+JcrSjsBdS8rGP+sYF6d
XmMZkdVXB3zLcmnn5Y88RXQfLjRxD3vn+r9ciITKxpEnZrZ3YM7iPjq36JaYG6kh
Eg2bECvInDEX5TpBMgR4welz580HniisGBSdQ13eXZ5crfaVA9KfxHSak/DWUJoQ
53wtn2lsst5GkAd3n2/k/5v96+64VMatUBgDjlNHxXEDBKQoonNMYF2h6VqVrfTM
UBpjc+WPU2/OFFJ1iJFzxzZ+uT0jGuLQCZctlgc1ATdtJWMRAY/HMXCGa0eGLzjK
53CGdqBr8njNjw5xydSl+Oq66cwON/t7u+hZb8ngS7MTN+HoeT3sL2tzbYDUVUdb
2SPUCCkRDKcQ3WEjEDrO/Q==
`protect END_PROTECTED
