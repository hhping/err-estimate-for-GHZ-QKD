`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aJz63QIuA5PIcxScH01n0b4HR2dSOHdRtTDF+4PUscs/nPv734owyLbz2T9o8wer
QPM5UnTcD44/kgrLBjwoIdTlz6eEbn8JhFOxyBblYkIBWJ01H9UgJLQf4sb1mOTo
3belLLFlYJiDPx2WgKoOMZc2kDJSGakqIt1aEBz+dDn2BuX2Xn1jegMFDLm0oiux
6pJQ4Sscvs2blEQu7m7NxmpXFTZufrbDUoRDBOxObD4bIqrFm5GF3bXbS4UiJBzK
2YdXjk3i4cyHzBMgxn8GsE3gmmfMrytWg+AcsBp7uqzGXUA//FBylvwnbO6QJbyh
2zw/itArFK4Uql1GDbIvdZOyZtt16O8UrTKEzptfQxCT14fXFI+8Ta29QdYS+kon
QFd9IP9TW3SaWJlrrAE40IfmuDpIGPCBthwp8dBtRQXBX8tigWdKYXoWUVk4ICkT
tHKwzoxfIYuinnkUw2H4X7Gt6j6EY0Ost0DW/uYvQCHyi19iiI40efYHbmdTJ32E
bxaw6jfNNn0gBO3oKIJt6KVzd5IakGjT2DEUS1ArqvPdSKnVR1IIBsj+OdpY3Jqe
qrUSn/hXT5ZmCqBMdo8YcTpgC9CiVyS1cTmSV4GhjQxqITioRIjNRqlI6gw9vMmA
KSZnIp3zE1r05KNLXemPf9kfqgJ5YN4ABXoW7UBAobHD8tDReffywHeRDSHCM762
TkRHtYXqbh6cZu1lb3/FPXT4NoYK65YY1FNu6Iq+jsyMjpSpXXavjjNz6vOfDhD8
sZ3Jc68we7Hggv1aw3/oGayYvZMjPQW6rH868ouOR7OfQoLJxk+0nbzbVPlcb+uG
2g0Oj4pYEjXLAAIEDMJdtJhPjJ+w4aK1eLm5iZsqda2NaX+ir+8OaHu+74cn+VVz
72oupwxJbsJwq74TFAEv74fq9jc7kjzd0XCNlpOnpt9TG/JD1lLRCrL4loiX7DzT
2Q2l+GAfTViJvS20zsnJwF1LYnn7z5hs7FqNuN+3DiwZZok6Oc+zqcG5/Lt7+sYS
o4p3o+NXkNJul7cVBz889kBf6/N0n30/w4eK98aoNIKCkIHdhyb8G1yw+R1AfMCn
oZw4JO9P/pIbXZ4sOOqHEsAi+0YsG/Gg3FIyTHU5xI2G4wB9VYekRoABHmVwWK2b
`protect END_PROTECTED
