`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+vO4ogVm8eZ+xveZqDZ/X3Q2LuJh+MsijXE9+TR5+a0mcjamGV8fNP4XS7oqXsDf
aQGFyHlo3Bx1hJRXyEVGaerUuq8r6MsCkLzHiga7HDpuElCOp7zs+jW/YFByuF9z
0oXFV+AZ8ibgDu7JbuiGzHwoAQNNbUnnlyAaFf4XCWSp7o54FGqjArEmPfa3Z3ZP
FmnavQcQ5aU6oZ5NqJXEn5lJDxO2YX9MdNDj3EOaJFydIFzdRSgF/PTzSuIUPBEj
Hfkw43wZrmb2aTEv60iy2ST6UyYMrnBC+GKniEohs+NVEmYYDAI4LW9K3BbeMDTk
QiL9qSyX+q2sebQdohzPgM3Kk+0UMZKZKw+wPQIc4rYUsJx6YQmpemTuw3Wz5t94
4V5W3p4ycLoKfwSsTYvGm4yRd5Gi4a23FvdnlKVGiaJhzAPcE9ct7ILD8OOn5z32
Gnd3yEVD1bXe1HfmbHuFeYleWQJJ3PzePX5n6xJw4c8=
`protect END_PROTECTED
