`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ObBdrmUSgtGam0bpjZhZZX7Qg2FSKKQd3zOVCxIQpvCJCZGE/Jd0qy/RD13tigIa
YzwnUstLbaNUGOWb0e0CKTe0+bMMLbb4QSUdBUBIQ+5fdFy+BLVaB0wGwdmkZQ8L
lIhr86xIXlw9If4W9g7Ip6YX2KmyRTvsLOYOZmjHp+lSwo1dtbfMuJWVtQGLE5v2
UO7YwtDDrq8sQ0kBR7JOKBG8OhDOeGap/CMVeWgbu4R4RSK79NNXteN2sw78unpj
PYJuTN5RW6lh1GISS9LY2f93t0YAqamV7ikYQPSAKLSwc/3UMgc6nTdgtxJpsjk8
5YilVqDoeuFBTbUh4AKpsLo/IiY1IukDwrtLbxa3nN2zZkOzKItK0EGxx1eGexJe
zeNoE2lOkIctXETfYU7a/ifF70W/MSz9XvcBALn7+/+uMtZJLFu/Zqyc+JockRQk
2cGUvcGyN9VwQKxOsLQFrgRWEm6/nAypn9SrdTyobXzMs4E/+KNH9yNK11/9LvzV
OPmQ52PDPlSrb/VUXOTS8CwKdfI/SQfwHbDkZ5sLlwlK2i8QccmPEsKWg97M69v/
T/U5Lm44Kw5eLv/GxSH9bVoonGeW96x1Vewc7UpqR71TExXo92LwUA5BlIMbAMF7
2Uphy/MKPVm7aO7DPWG3Z1j9eGm1FPlm/fY84PFYHw6zC37yl1i+SeBnIl1qj0QZ
8q+2MyoiIk78uKsbJCpT1/D+RHhQ1uH7LvikWm3jRfP36x2Qp4wAEB1RsQNxWoON
ghhyaADrqbTTRYgaAge3APSMYa22Aqafjut84YjasrVEZf21xQlBXAVQYYbdeyAF
3Mv9kUQcGby36SnpUu32eFP2j7qQUKCXMOd+ViBdjE9p2p1hXyicrl+3gtViTa+1
4z2sRKzgYqtIq4JhYQuNBtSTGEXpkdcw0zwuFspEewQilFjQqNs8gVk8703tBj3T
CztTppD9rVIj8RnDpMdzNLPq/T8bFsaHLcg7vq13mxg7RwZjOubZcr/5pCquhKXu
C+AgSdI5OoE1oRbnnBUVYP76KG4hhCYFrX0Zg3UiSw9o4KpPzetM6ZVDc6zDCRxM
hSv2wThQGKFl2pWs6NNMf0Ewv9FfjkEAXQa8Agnjh6H3uibEbrL7tZ3RZVlK7DvK
e+Pprz/WL9+Nyd+oWvrUYWMp/qF3vgN8MzxWr5gqWvGHWuwkf/SZRG9473kyHAO4
4cB88+p1cDUaHqBLlTjT4hklhL3PGKCboZWOSC0+txjuGVbjv0WtW8eUd3TD34qW
7BJ/RjhiPJCF3jBnDbLeboGuri7S2ozy6/u5xTyg4GWj0HB9QsuNNqzYA8NYyyUI
H3iPjgqxzREUq5GNADEaEJdTA8tCvM4TmC3BnIm/n6Lki+r5rUDPQ6hrN4mol7wE
bgtwfTIa2SDaXj+752ExrdtfdlMtQx+0C1lnisc/AMaLJUDySNhs53Yhq5zOiN9+
BwmAaaJdR78omokHH7bk+49LaMFhS6mEaxlvQ+9SxYEb8sETbjqpvFpzmP3BzUVW
WjFVbas/DACGcMRQKG8Q9LM4Pdtu7s7O+5k8wV7DolvBkQS+EjoX7owZ5pMY2M71
C4kFr1REyeEMTfzJrPMZFRTb7aS3mlQw2e80u/sptt6dGlwEOQUUh7ZrQ6eTxCex
WJmyn1kovZ5yMjMyh/l5rPaxfhwSme2V3cfbypODBFie4GSHXoZRVqstcbtoAbt2
plKkt7uwMIocR3Qi9YrqMq622jlaj2Jl6kFxLuAbpvaFyY81dB2CVHc1LQKhy3Tl
dlLRSiq6pGp3k1yUcZKGj39VgQrGAAatt2gD/gJdKARCavpewyKwUCLdkbD6M8qM
0i/j9NW8KtZYFIa59UEliEdYrNzHU5YhXFpziCZlhahS18wS8zGPs2Gcdze+RhEb
/12EebYqBwlNKjpJEp9zNaeThTkg1HbT6J1ohE47JQQmFfdQW7U+l+AbJfWHReD9
kWChAmWFxRSEEtyvkUOcYVDC/x5520AyHqomZ5D8Nu5Q1n2wOwRFagAsK35rd0A5
WvJYrNG23yFdwsFAJr4HnRMRqkDw9UHcioEyB81dPQNcjQFDB7g7ruLW3liUd0XL
ksHMFZm6vNa7N56zX3K48OOEbQqPxEXfslRpxunpAcQGnvKWmwxpW3g3xj1WLUFT
AmE2BDrPA0hp2K5THILFndTAOY2AhrutWvhwy/RlhcAPPH79xkAWieTx/Tpxjq3h
yAojUtH/6M8lpKW59uE4eRiMIEkqZ7lcqZEwCRV7sCfXh3kpZLJpbgq/IDE69m0r
eaE4AGMg0Ba1DvdvVJ2Tq79Lbp10ymvUFqAReM2U3bAUqCr61SUER4DZjl/SE93C
1cSwFHxsbQb+TK15ty2U+El0WJas8BVFF6N2pwLSrTNYrw+WkrwldNyFmPIdlVgR
2A5/Cq52YCgLDeX6vpDzZWqp5oGmJYGJ9zhEMLNf5GEtDpJt0j5LzgicmHCPn0BV
Ezggxvo3WMq59X0qh93rqHX7/RDOWMQ0Vqajh71tJfDzjfG88j8gm5dEAsOupYJa
W6SeOT4NjPz4Z0n3agiYvlUq+ObUzJd0PDzfgCxsAxX+Tu2ogRxMNGp5hxTCauxR
JW81wggzeT/z1vhwJaa8xsb1Xjazwwo8pwgI2HMozoN52wrzIcypnQwiJWMw7bJ+
78dnNPbZYIocC17IkrtdZwYRxpwaB9MKxaysas0BQNhzjf6eQMXcwkBP+0OhU3hw
9VA+h2Gl1iqLDgGJSaoB3s7sHhs3lpaOf0JlwE7PQF4wr5QlFU6OzNd1tA7EPXFB
1IfXXymfTf5pHOd1PFq1b318cXezz2SeoJ75TnC6vmq1Q9DniJ7iYx9dzbvHwdtz
LZeS3hCYWAeBYs4sR+z6pr/cZypNQPPGWFcDPH7D7evWYy1b9+Q5B3wOpjNn1QB5
Z/TbWgv5XGprdSPAoPmDE2C4etLbobSGcSXmqlFCluoWSrk+RElCmUbeeKmtZNFP
WSylHqxUTRBQlKVDG6nq6G88DPsigxwL03UMcc+tc2SKB7MrrRwlAkcOiLiTohFD
kpvyOvM5U44TBFxaPAbOvMGDaar3H0hM94zQrhacKk1/AenCuguuGglolAKFnsYA
tSGnIUWwPdfSayozhV0wAF9TfPs0NHQmKJHQo5HRYe9jKyPTKhO+uEZ+3gNEJfwR
3foZKvWj2hZRrk22DuE9q/uRNBkp48E6G317Nti7cg8pNbGoVqw7vjcwjb2eWQIr
+clYBojTMcs1Zb7rvlrWxSd4kmDT1zk04W59xNWgSELXLepyPmsOoCaCJWlVB0Mh
dRGQ94/OfBusoJoXdqCKzklSw5ZSqObUNMOP2h/91L28gY/nVP3T93Jn1irmyVtB
FuPNWdvWl7b6Z11ZpW8ywUBi2HL9HfpOC+LRh/fc7B8NkT8KiVhprkZkcYA6UKrx
lUPhFmLARyqQ9mod6lcqrRncsz/r8SCH40CStKDtmDysGxl0Kc+L1Aw4w4lRrTSV
u61NW4FN47hDQ86Efy0Ar1gxcTFlasvxVIYBNOhk2rohXoU6ZXV2MPVqaBMvaIFW
dMQf2JdRV/gZnBOKELvzlaYHyo8HaQ33UavP6ZRy5rt0bg0N/Jssvhhz8ngDMbRV
C7w+pZno2pb5uBYNR7pJlMKMw2YdNauGILrwy5F7jMxk70Dg15c9UWScYuxKQpgr
B4gLZozYFER8GVPAaOKgY1yBk0rZT2FtSmp7HC6L2oQg4/G0Mmc1e7xO9Crzj3Ae
qaRJduSV5yF01g7q7ko4BjylR2fipm+vwF3sYSp+oAd2Vxtjo1/jdf/WR65ZaBVa
cBvZdKaY/JKZ6mXG53TMQEwQkTeW0A987D5eAh/mqvWC/Lk/hfgfE6DYoSHJGJn+
Vn1pYOu898b4oAJM3L8gB8vdcSGoVHYzIGbc80m60SD/O4eiekZ8WxNsTJ2aJDwx
BFKn4DOwormjA4/tCRTcOPRCRRibrGySBSYEEnwk3d9SCFIzBADfdsidTkpZgvZY
e99wuacPj9KfmkXeoSRI2MBc0a1ZM8fDc98PFvxvn5p1ILKhu6GXTSHpmayBL0BQ
DPzxBCpO1laITyU+afIT3T/WY9+Mn1E3V1KB35mdXx0GXWx6cqJRcVGcy8U8viK2
dgzicnPMgwCB0pKYwdxfoZ+aZzrDVYOnCbDOgiZDhv09C2jknKSPL2Bho4mAl69N
lgsCtokCat9OY5Ln98R+LA1FMK2BKbmUGhj/Nz16wFc1yxUP3Dhtt2lXGQZOz2mA
OHllC5jtEzKO8PVy6xgMx1IAN37MH8jimn0drRRD4o7t+AIMEw6jlkuJvlPBL6td
J7ELlUeG8/fBMMrgpotZr1Lx95KHivtCHh6BklVTPjXw0cbLkxv9yhzMoBZ31GyP
s0k6S0M6hEQVfwaUXivssnqLYBlvh3cRng2/R6qIswRa3UV+i+r96ihW/j4Xcil2
KiGVcZUmvLexyL0kkCzZls2aN58HKjUBSz84XH9k9CMoh5iuCq2IBKSCV1o1DAes
B3Lv/oUBPUa+TLztsw58PGy3+VrQTGZ62ZkkjPEmGf6pXyEQzr9fi/Mj1ZQQ6Z7W
0iEKQUHSSMOoNpXqJqDS2jORLGfJb3qG0h2a3E3NsLFfAUUjpeo7+ROkOKv9qAhX
sWBm6ZjMbAj0zoH7vPmBwpoBcSAdKLG9Jb911RuWIHR6XdazDRsm3yDjh6LypDO1
p9DxLS3ATThBbdZk1MTXrp8p3rEaWhvgdRfQpvsm/WcKnEXSeGf2HFZgXYtutmdR
R4gEaxi9ZR5uQdadLFiwZ2fSr2KHJpLvfy/4NhYeqvToUnS6jO5xhuk5i96/tVut
O1x7NB6hKTNOrRC40wxUZ1Mxal9yQX2UBLZ1yU4VDz1XnTdkqs+YN6RP+ZpIYw6q
sNXWHYO9oUDBbZ2NobkgmKi/DhKeJIbwiARx7yNkOdO4tW9LSa10SxoemzdsFPGH
f8pfBziv0k/hlJzAfgqafu+E2HgxtvWQdryJeh58hTij3MW23ZmuwLSkbP3Vcgn4
YDH9B40emrl1pQ4w3jwpOjHj6/ZLGQgDrdeu3J9rhKkoPtpbv96L/b7kr1H9sWpl
fKsOZza3giLxoWbfXGDlCy06HBQguKPLkSyYjpYQam8YV/gUAOK12Nm4/XEoKl0p
QrYPopd/BO1qoCv7EnSgH6kjmuj3KziZIc9Nf1MfX0YrcfLGhEIu5/n7Mex02oOy
BFevHIy2Q1LfDawdTvpuNqaDUC0Rt6cn6Ll0+rxbsHWf+/DZrD03ICWD/Or83aPY
j7xNkZjCrnaMOvy8mq2UPmDt5HjbxPGEofWcUHbFX8whqg3Az59N9pr4EvnVqyJR
qE/021oJmB99wFJF++Emx4juSAvDD3+7HEITmOaPW3fcCKxUKR3HomrCDukxfCZu
fKC45iuJ1c7tKpCvb7pXR+kfsRlxmwEk3O329Yn1d2FMvjBD7xlnC2gzgMi4H4Im
FFR4uiJF1+CcGruxYDvAUeG6zI0q/vBI/cLc7jPSEnSXidQCAgwPXa2k9PwFaKLd
tKXlBAisFG4Ta/rQRBbdHlB+vVMWSJFQedInFr6hWWr91ZHI6gIzLDU7hSvMaIqs
3qj3l9jgVp25VbgIb1ZpPf+HfjlhDNsjRaoRtxlsOV6HuPGZbf18TMMwY3lyz4C6
EWLq4C9ZS1BvBHF6o7lJdjFHjPd3LPXwMhwotbJ//I0m+5+rY0Tge8t0gdRnQ+qT
dklsRYWj31of/efaVdMFYDJLH4n4cmeba1sTnH/TAjNUsBzBEnoJT5jzB3aHmtQW
fQEIvePtAiuf6BP0vFpQhHyGEfZkgy6ZG5AAVuvH0yU5iMLZvkGOI47cxlDn+6ov
o5XWamf8QpChzerwpfEMLYUabkgw1xC462xkSnD7jVHSruq0BmYK71iXYRIaHlQ2
mUUcc3lOAPMmBZp/P3d4Q30pNol527lnZVAU3sNEjjoCgfgBwhW/bE2/7RTLrV8N
tHrUrgwLu6NknyckiNWhA0eNvGliIa65Mtga0dbctEw3PlMW4wluA3Ji79j2OIng
PZ5ECBmIsCQ5GtDtgrbLwDiuqlgZVx0vzkS2FqvfWstJw479rutgh8oYEz3BonmH
SWYc4/ygvuIP5kk/0JJHqtnF1nL0/5za91I98CzqiEpg4x46mAp62kYG/nTg5DSk
BMGyEKBP3+Z7gszIYC8Z9qehg0XtoeVjhc6lpgLGH3yA6/wgyPanO7BOhOfsi9o2
wSB323B7Rd+btf9CSH8J5wD017iOBDm4wwstR6C7crBtGv+DfHP+yEKYxm2f6xjJ
awQG/jvE9HJXSuCJpCTUXe5jwphzim7KSpXZXU9DRm7SpB4lGs26GWj1Qk3oTFpm
PeLjVKx7jwYuYn1Fh/LHx4k6hd2XfkMQSbVHB/SB7BgXsLPBnQQfMuu/JQJymR+j
YFXWZuKc1TBRpJHBgkthq3vO5qi/uZuIAPVPHz3JnjXrntH/EK1OYbB0M+qxDRmZ
WvKxgT8S6DHdLvOh1yXKdmGog2agkqNeXr+UVowaXZDklyc9+Rf3/S3KU0Xiw4UJ
697bXAHblgFGKA8FS+Rq1G465FvgkV86EFn1smF+djN47lNWJoUoz/xW68vm+DQg
WHZ25IsLWBUiWLjUD64fHg9KFsN2tsOiz1shgl/J/DBl4KnM7MnFb6qzMJUcBSGS
g8aAoL2+vdEwvCopfkpjYMebfeGuc2/1V9q42cCqqryJr3EgZhTexVTpgmENDK3n
NkgmARQVbeH/sC845jymIt80bXSH5Nem+X50Kj5ePA7BCRWc3BiOSB4GReDbbce8
0A+ADA7Q2mi2nv/Zub7b0cQwSaY1/viztjwfjTbAH6fdiLTZ76ArFtm16TbXPCX+
wCmBl87f7phEXG775IJgmYDMvAoU+5Iw7QfsFJWIGC8hPiXuRKv56gxp+WPqgOlK
Byh+fJCMN5zmpbFNN2YEcQt1L0yLYU2fH7zMaYJLDhBCjtCUXKpc+ImhjkAVdLMz
9aIlVmPQeom7BTbnHJMoSjX6pSGiTeJwt7UYCwqnwhs19SHzsvLNDkYkDKcZyWm+
f8O4tMATTuvAJHIxM/IdsOYgz4DkFUCq4mP2m+WxMjZhDTSFgN1tLgOSaBFptm2n
rhI4eyEYlafzyeu98zZSSrehpj8bDRX/3K2tI6OtF5/nX9/W0fwM1JdNaGgMMvyH
nlby0+jj/gUFAfsf4pcGuvDXiAKzn2OFjTzdUfXdZizNXdA1SEs4qEIFlXbbfHsL
ldYhfo7I5h2NEwEUrh0rszCLAB7mDruEtGrgyrVO0tzcgudzHdGAw/8tgYPcW1UB
AzbQDvKU7CfEDcQnItj7SJL+t/QI4ogtFt3YkxOlPNm/ne/J499y+QXUx8ANkYuC
6l/fsFC+o7omumFY894m2ul2GKdso9+Do8cKjWnMzyYwPatudhSUNQ76wM62Mso5
yEqoPmITTajIEii16o2Muxm/dS4GNbbgfq86KaGUIyxt2zeKOovnyClm4aTiKDvl
uwsNBhHze6UrfDqpTyP5TXhXz06Ho0vs/0ElwZH2qA+llkUsmuCMsyCtp4h64H2f
DpkY2tFfVh2xviI0NmGaWJYuXdQIbqzwgGv2ZIswRM/SyGZHUwCNy09rxAd0++4N
TMF2UMbNLkrc9kCddKTttbRMv4n/8uIoEzKBp3HL87iH06nSkxvlyA2T+RUg/BXL
VnmU7Z5nfk2bG9uw+tRZpnn/2TZWBxGzV0keN4VCJXVuqDrpEZJH6vH0xaslQ8ac
bMHWVXM7IL1XEhNZP/G7GvxXJ6dHu3D3rPm2vjeauS6+diUZnaDrCchldr7NPtoz
t+tC7eCG/D2jy6NVq21tHyqygAoqryzehozDaTcrUzSdPjLxud8vrHJlLB2pouuu
y+DQ8GWciDot8MILaaapLtPdk9nwE4oEHn1CiRpuhN9dcu75lYXBkF0JnNRK7bK5
NrpIHL7J+2QT3U5Iq5cfYTKoSb5dxy9F49tnX+sTEHv2+Ti+Z63z2kMtEnxI3n3H
yuD4+4VZnr42l1Uc1XCPPXrr7OU+S4hohlRpNs7VHUSQKQcrvRqnqGaNelErpJ7v
cRkTlsdt5eeF6mAtRa5eR87N5djc0dNDQMjcMcYFOSnYzq3i3aeeRQF7ZeIqVQZr
l1aCLLseaTRrEw8m+u2v/StnFCxjQh2mS80O672NR5cFWeA+MQSg3Xc1I4gAx0rA
teMEBXn0Z7Sj0Nx7iI8wBYnpyo5ClUMoxzNUutL7/Ehu/cdLTJ/adhHDgk0sQ6V3
S0BYualEN9l/goieK4ozHvdJkbgdtBD9BJmb1JPqMFAqH4Gy+eUwKujwmGd06hAD
FasYw6FxuYXeenVOIvRI8odiJ1zUuD4Q01JgyiqK+DYLFPwssjqjMSWt5tyInlH8
OkgQ1n5oIQCicaRHM4AjmzJavB6/YuVQ+MssdMmVqf+BMN6re13E86mc3LTPfBRw
t9Rycl8e8CShWV3FlF3z8PTL9FfMfUdibH2hSZybbNWiF6X1I7UoA23T/kMh5Thn
udObQmpiGoHEjVq6mYXuj7HcwVwtBdgeIfTwBdqZWZC4Aw7RmcDjo42WFXZ/6GV9
nx/RAH1kzUIQTxu3qwYW4COr7rFdA0iCjlM2EYlVZhUossolSY//7KRx72qr1ufW
X639sV3X7ZLBYAUSECpKN1nZ9mO+gwTME34hEMOCjOrFc9hWcTYOkAVCNakUxIRu
zbbanaKTdXGuYK58itPS3vfT/VH8BfJeuJt4yfeneIRoVwoiigz/qppOKNhm0/uf
VuFcyp4poLgHHYvcynmYDMJiTtlL2rCqHSJ8zXWwsFyDnaVVy0Q8GCfOX6bc0jAB
GudVMGA/YMWR7FJSkcnc5r/y6wrMt7o5WVR0Lo5AU0tRhHJ4XpMa7aXDvodp6yJV
wyyNRTvzJrP/js5QwiBzfjQs2BAQcu7tj8t4p4SS7b/6C1L602qya7kPF9mq3jCv
dqLOOikMfZfEvaVEfGekRRdq3x0GyajxztmR6Jn71kl4aO6XAiWTBpRI9XKeW7K9
ya80pER5YrzsjM2Md3tvSYiC/fh7DscsPswuIvk/JSEXhmPKunHJqm7JCSagQMAo
qhzZjt7oGNxBrtcQ0ZL56ILBIwUg5WUuED9hU6tVSuAE0obNJpvubAWJH4TccCqb
s1CGjrSd8IfAB7IykVhZZaQa6z+q3OlkRVvmmq2Ry7K7sAiTP8dQ5VAgdOQ+rNAe
15zXZy29Y6Eug1qLmPSdVMSZvHqWlXkWFKbQ1BTXD27nn3DTWNDnVb7KwC6t827G
ep/C7wFmeK0zWYPOcs0mjoX15EIatUNdcnQ66fm0mskwJbOrBFC/IURajxMp3rEa
UlTNqxjCaqxtWCspQjpdHmOJMUw6/N1F91N0EtZJHaHl1C+fPpQDPEc3/T/14hyh
9bmcgyrZm6cz331R77FEBE7NI1jVHWKLBQVY6SpSp18Q1N8o3hUA94baSv5BhT4H
lfbJb6jQ2oHhItQlai4gi5PXnwpWUXQmBuKGcCyE1Dsa2NqW91pSkn/7mkiIocWH
Mi78JXUTQYc7XYpVZ3nSFy2/GPekX7rNa3oYtWD2xcPWrREgFnbIY2A5DyeFljfs
Rd6JvQjtee7R/9I7YzYep4dtYj510uHxEoGZwr+/BVGNF1p0NM1aBGpLe77th3O4
t5KCj8SlFnY3Gcl08+WF8zTR1IpjjL2GtZJ+HdS+9MHlARD8pqKE4AFgcLcRkQFr
vgKVR1he9AMyaTmvdgnZzm9IBCDLadL/WttpX4W2Lx0+wJes/qsCNPdTZJ5WAMSP
Gb7i253N7APqbbFJwsvHQ5vDcO5sVS2mXoditnKsfo71gfP1eG9opdBguJwMXNNT
c6ZG4KKQEZUQdhqU1iFgJEdv47FGG1LXFnytl8PWwbviZVdMunULZxcLfGzMAUtT
ktbuGe88Dt8JR5037J2Es96+sPenr9yXutjKTYiaO9RcabyxpsnSP8hCN/UH/+0/
y8h9c4k7WtX3j5578LpmVHK/eG1ORHJ7UH3VfiMaZ6cRJfqTFAjSXx9ZJD83YJLv
T7UyIyhgQu+DLZFrE91q+GELFLexXZUKfkyNw8d36L/vC+dbVQ2lrgvBXalVpU7A
aYuPEioOhh6WXM1PYEediTp0Bc/MLUIBtoPnDtm+rfdG6z1P4oetPiAltpLTwtL6
GYzIQktPK0hVFHrma8gUze4MXwi15mwla91e8EbjQbGDtDyQYPrzMm2WSborXFlc
l2Amn8q0u0HXP6TuRVZGQEQOBcMxU4aDOtzNfAGVFkxJvaQZ+4L2qkmeoqoWZlOP
wzM9fqtW8wbinJKL9Zg2/uSEistS4p6Z1B1B7oXfF/cpmHWdn4SvtJqPSVILmnxZ
EwQ320CtU2rzv4dbTfZrKJlPeas9qkZR65LbHymznyFNq+v+hRFRvFOeMorKP8j+
+u7xeOGQL2JhD8qIhDkyn4rw9UCYiErDH6zcUK8pm1ZGtQ81Lm5HfI8KvVzmOr9s
vKXiNyURoPTxmWI+CDDgbXDw5ZWbQzPRDDq56UWKRwO/FWADWAPujJibD35/GhcW
7L/eosTG42gc8Sq9N9T0eIX5zGOnlEpdgp6LQZL4FmdmWLfDpqj4h4E7GvMUByPZ
alLH9usslmA9iJTV0TiRERJwDAXam1lhrhjcmWpO1SsmTsyNErT0id1A6oQ5TjLc
kXrJBmrxLRXVsAau45uPL9osThtfAvPWSbJyjTXSAeWcaOB1TKfqkwLDCxByKt3w
Ac1FIu7u3SE3O2lSsVoIBPRjbs8HnBbDvWsC1IkuV+K5zfQ2j6ajLtXbP/ENkZ4K
66AS/YOILlerlrKC5q4/dE8SGtBnDl7KpUPrlerTqdv1alubetn7hE2hkVjHnyI3
bARnLOf5iAIVwrj33tV7uxKuzDpxzMxmJ8NKJ+HgLfcGpy3tc15m/sQcYtJoSCjI
kcBFMyEZt4LftgU29Iz6EvOUzzUYJkTqAKjJbzhEUBXX5LxxxQBgaM34tvQtwqEm
eZiePGdsuFAmkQWF6vHaj7DSnzSufCgyHCChRytxzimZiblkbR+dO/joGBAhdgKl
P5zbr2n2j0QjrXPxSaxc2CrD/32eBQFBInS+p+5nC5rHB+SRWGFu2ejcTRY9m3pI
l2AYJ9QqshOW4+eAAYmqdUVraieaHzXXc7h+ahXtb67NBLf7gt3GL5wMICp5+F40
OV+lP+Nb6rwEJgYSzhGZd0+y2zP3lX43JLokTGmHrSVJtNMFgKKw8RTN2bMzqX/2
BD1AP1Z4tgD2/XS+55iwEDcnfSH6K+YaY1eZ+BelCsLgykhHbAdPLBBExoEQj0H6
HnKPJ3flZFHnKg+ITma9i9JBzElmOPB5Bdba4WBPrf9XvUHQ1pro4xdfC/m2YKPP
OwEheaM5KnoaYcTJW4CmhLN8aUdOolGn4tnJ6lVseWNiQjwyx76GnbtG3n78yPxI
mKFC/N0coNLrCTSl81fBNgmksrE4xwO+nreleJBPEO7EliBwQOzUpJAoCvdSvBBS
xAZqcnDMh8ZdBXjMA8K5ErRJIgpSceVumko0U7nfvF+xE6Cc+EycUzM0eKxcW6zy
2eJzmdoQHYoJxQzkjOH83P4B3ZFfKUiE7eStyyqsQFqyPs7cJkS3RwK9fhudtlku
9D0GOEIHZT1SF4AbA3waqDjqTsuYay4GSz9+Yj8yxkV5RKMQwrGonkDqg9Q1MxB7
CSDlY6EtTqyq4i++AcUaMjQj3MzjttMNNw73xE2jgZgQMxc5vtPuv6omRs5tZs4K
99j3bb5p4Oq5EnVNUV4bUANwWnIFPbeweqq/Q3OlI8+sZ/ehKhHNRZh8PE871mwI
8GywM7Sc5MMnfikf1+/HKJRuLksCEnXkIXdZUcI+VMW2cofSWKketC7ZDN5c1DOb
4138ZKAKkkdxo47YSz/qDCvMjPYodW3gFkLVFY4DBlTmLiOpD720SUBWMqWudZnZ
6diCW4h1F8igCDbhK7b2Bp1zNF4Dw/jRnRmNexSoJDinJrwqCrIEJBRh2ysf6k3C
j7/uE+U4v02Qc4PZoVPnPNq3OTQXfS+BEIbmF+fW/6r5WCN+fmNheRxj2RlhVbw4
4Zli17FL0tc5YNOmOzZTNNmmjc6ip9DruDUJm16NAyjcvS9/ng4nooKMbvbDbEO1
pw6u/Wr90Q6pDLsLa4Bm4/1gkkTUYvpJn4ZBtCwjveuPxqOmKQSkM5AXdWwoPprr
3IIyvW8dsfVHpedrxYPhYXU6oxAuNJY7QqIv2LQplwlZH3WLBwobm1kZctgJwYSo
nvEP+M1sMOdHJH56hghLpv+RAZExc582M6GhaGNrV/jXReFTe76RZlr+GtG2SN2P
8tX8c7hrBim+0/d7n3nzSQz3TnZeOyj6tD7nTCCVmVGUvlE3/fTBVaZSQKF4jpgq
6IEMq0uyraN3InuFq9k7w5pYyskVS2EAbbB54ae6Yc7k04JcAKnSHqxbfsyW8YLr
aBXGBntVAvePOcC5FWkMCSAbIf8GpXVFB9VNIKpWal1cE95cRQIjPTefXVEYSdwX
YNXbU+67n5KPNJdMCTPAOvqOSUyP3h7dLICrpGfqYJ7Yl6c8K6feP2HKqCiSSbV5
VVqEdBmqQLUAJVpCtaW59wpL3x2ZbF/HXNyz7PLZioSfxOYRDobVYQFmtOGYtBBH
WwmkxPB5RdWqFhPsE3m3KotjnZl3MR2IpXikEoiOYk52T4VQMOb7H1eODa35gXW6
abPAvYNKM3Xqtwx6rf+We11hiDp+uTYtmtk+gEQGgnxua4efosQZ45+zJs0e27Ta
Cz9CRqoqZXLQwu4cK7H2VBCFz+MLjH5kfaCaV3RV6BaEpkMn3K910vzHmgrwmQrj
y10qbn6ItQ1Utm3uqYxeoK2oPEWvqmO14vagxtaLIHGEEuVT4Agc+FfK0+UCKIzh
f1pfnfXrIbBa8G54SYBSk/qETwdss75TagroCmi+DLcTAAdWMcba3EQ4qsQoDKKh
z580hg9hSEvG3qNOIL4+FcXWkap6eXopjIcnI4f4dNd1E+Z7HSeivpC+tJnHnuKz
IjmZOMQEQ9ouaqD6Fi4R9NlNsnoswB8gjhv857mhzeAIAPoOWuyViWolUeqwaOWc
sb3VHqvkOkIDC8prgNfjJD18/X6yTZ3vOIj4D0b9iywD4kl7oE4Tby0cAJN3fl4a
7Y5DUSiJKyRG5KQKJqxNM48Hkf4qv9x68fYNt8d7SaR3lhZ1zCxixfmOlqGTZOvs
0f4ZyzzSz62gszUrww3SbBdJAHEvrOE+0q9BLxHheuIAZErv/Yd1k5swMsFTE5YI
X5fpIai4gU83ochI4t4f/mOhWjPbJNf4mmasSBunvq6njFxlHjSZ0YE9KjqC+rA2
f6YzjkDt1xSg95LH3VaV5rs+SmmOw/i+ftmB6sZz7s92PZJyNv69kEHFg2YWEf6F
C54WWcB/I8Ie/nMUq9cG2cXhahJq/Uxi5kpHQFiUnCCG/0NNsUUl/xtcfrIeXqvo
vyR7USxYTOxPIoEaGEE4lNV64xRQZyF25ToxdPXRXcq6vYHloWjx70UEjmq81ct1
OuAKOyRM1R+SaHzsbj2CWCUmHQ7EMt8aT0smZqzJlxjv9xksE7OOLuMzeLs1t4fR
ayW0xr8Wrt1hK8Urp/OZk6js4ceehrwJpTdTQJ+JNYukI6QjpZ76g42ZS2R2cO6V
pL8Rx/V2zOmhB9gasJO9MDiULmZGvLMNczAB2BQokpAiK8pSHZcdIKcviPC+pfH/
Bd/8sA/8K+48dcFfeye7lQT6P0D4suVKKnfy99Mm0QX2EtqW/grNQsilolD9SJ25
y39s20eExTIm3WLa1Z3U+pwB5w30soCrbYtwQ4ZpPQcX5v+FkRxKi8WrUf62k+SV
k8SuV/km/T+czkQTzZOyyRmikf+NsEsN+S/bX3SlKsQgBKd/r8E+7pnphVhGFYQl
k/vV1x5UXkya97LQcozbJ5WFE7k29MuuvYMkfnm2/jeSsXlwcPshpe8bvkdBVjJv
1f4Kuy3tRlxVQfK1kbG5epjlDUslRbXe87wlODPNElVEw2A701FE2l5V0Ow08uMa
yWFmZmk3zymEOzay6Z1VJSsS/TRaeWtq1G5XQGPLHAD1zSaXJ+8mKRK6MQIqY1pl
wK8U3b/4yWexk3rr+U098xGf2oVP4lBM/Gd/WwDKhTrk4o24tr0JJSnY2MsQfUi1
RArtptJgYJlXNKgHblKk3MRgUVbMSuitgMIYr/xbdsUUZXQOWtM4StF/S3bwm3Vt
bLA5BQdIGSZa8+Zyl7/0HEHgZv5dbgtM5G0IwRnNrVFqOVDq63SxMk4qNWBvSNE6
Y1wuBojCOLU/hFJdtZDiz1tjhdTHYiTa4ZlPOaNTZ1IkwokZsyZHnoGBbvcnwWHu
aKnJO3nQ5ry9TYR8Pu0kuB0etG61cOIWWHblrr5gG9VXNO25eNbv8OstzjRWaJXA
N3iXdSXROIJurjWG7mbQYOTNGJhWHaAkjOOUqdas0ixSxYlu0uDfWyAe/tWaptA/
fQORaB/r812VmrfOVuFH5e4mGAoBLDoX9UGu5+bgHJvP9FB5rUTAE4Q15Qe5FIWp
ExL+mGWwhGVS48IDthGdNLBGB6M5NJT4oX0wPjC8UGsRzxmqqPqb8ysVS6Dk2aPL
gbs/a/97ky0lTA1+L2J9Xkl5hgH43hHaCZxokPY1pt0YtvEvxmmPRMShFgwWOyOD
9FcqXfT/j1FqUPttu+E9x9cMZACs+LLhEStyh7UbX31PruHorFBomLYz6ptFyK9E
HUjtgeIwTATgQed/aEH5EbLYFUWfLuNd4KCzqxg2rAxTglmeCTLkVRUN1uNFEDSW
WngHdc4q0KC5BphZd8lrlOCGJ/0ctTb9jde4BZMX9uajUFzBtDV3KNiczkryk0nX
TH2iLBqib6MgdQejH3NjMyp/qF3fjbA59CRMua+rtk/OxpXUzBsRcbLtUVUIP2VE
S3WP9I78bzTQCbBDmNTzinGhkn3dpWalk77sftQtFYFdN0n75QNrRqQXAVCrCjWm
GHJTrdGO1iPWTQpY9CY2MZKoW8UEcTjFkfwYskorB+zkbzunnilkvRs9/21TydHf
n/1nAST3g1K5UTMTZIeUugH6gjM/j2QgDF/CJgRRHhtTTAuO9xkd+537pZHTNSMu
c4rAD3TZvTHofOGqSvgoERvr8aJ2oFlS0hYrQz6IhhD0FdITRxSiKakRXQb7R6e5
iqUloV3zvsr1rctJ+pn/5J1JMEBQT2aLMk3dOGxeEa02Yofxebf7ic4l+DMgCqCj
Qvl8USc3/FdohNRtj+/dCJtwgH/LpYQ0ErgtXDGQNotjkYXE8BUuCSnwszbDVUcX
Htog5CB1X3g36cs4UaDmaO2udztZEMs1uN1qGFYWRBwEyEFK7clf/UJxSlJDWLK+
pgtqjepdPjXOzZ6inJUPtmXUzjYcHhr0cT6Ll+SDBRUhFfsPIPOiGW4gZ0ltMQky
2jLv8qND5syta2vkxC1dlIDHR1VYDv5ekhZ3QcWr2dbcjge895ufHDkkG2mmUjGy
`protect END_PROTECTED
