`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HjHU1oP0BmBjmgBurSy9ccQKue6vLl9/Uq+1DXLvplVmw7iWIbkQiGJCT1zcB+Gh
qheKyKgzUnzd+DfwuoU+2R4KHCIHANNp+3OxWp6oRXzOVGEX9VrJvvHuQmPNQ0d1
8Et2QGq0eQv3YkCJ7M/nkd/1iJPHcGv2zBXOG2ZKCtfRuelEOrvSjNH65aAEPRSv
lqmVGZ98caBqU/QFInhlrupNT+LgP2oHWcl9AHvCouQzZdtpAN20PCi5rWjCpu/q
zGVuDmfCId2WXl1xOompxt3EBggeohyNdZykznfDlwm+60F0vySmOlp3qFFiu1v4
MuWJ2QsDhFcjM2Wfgtn4TLjSuh7b6itATw7X6nbbiDIgQ9JUKc89K+oc3Ze4lJP0
rxdcabyNIGa+629C4nPVEdc3Ke77m0nqv4bMmmVfWtbxP0nhHr2hYxo82L20dNqA
`protect END_PROTECTED
