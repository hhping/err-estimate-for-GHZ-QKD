`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YWP9z81d7T/AAqLOAMZy2NCiCAZ3kKQ5usjzaMfcPN0oD58Px9gXui30tbM4pPLP
fp+7cVd7tH39Ho6UlbH/OdFzx2LM9CDPhM2jCjvKnOi6fTBQjNj3cHZMzEapzqxP
dbNxRM/ahljE3L5bYGO95RQ+lKPjkgZnh9hlf/ZG4CvO9Fe2cvkZbqPJfi22/O+X
9V++cO1M7LRqTWdH0UNxYwBi3sWh6ilBb2Vxiog/EYEPcCJ6wr4+hhroqOvOc2f2
ilbjceWBwSgraIYb7GxiYkBE3Zr62bWmGgdbR9uIWFk=
`protect END_PROTECTED
