`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GfnfcRr+zOpJ16QxbFXisSg+c0ZlOxlA4HpfYPiGobRV084e0fxlb2wPF2lUgNkS
K1nAvy2nTS3pvzOj11NAQJ/RTrMReFIVj4v/T1Y69HwuA0sk0793GxFfpq9nChis
S0db+83BG7F9pDk1c5ZJuw7o9swD3uuQLafoHmYNmhWGsU1vfQwr/rwUV3y61fns
igX9sd+sxb6StOq+fjsFEY+n7CliJbcf7NHBKcjmZ4pPxTm6q3C6Aqmgky9Vd42d
CieXrcopyGxWl9ceuq7TyA9QLUm1VjsZic8iHKZ554C9Zbb26DKbiljy1FwwJP9n
CWfG8vesJ5XwEj5DMxTpg4bcAJ/EVZF0XDjbBbzmtpd+9uLaO9SU19sgf46uOf/j
VfEtY4vcY6pCjvCQkbZzGXcHwoBAgOlsTXoBRRbPGKyJJKqgVhlwWOPYhmthPzZ4
uta5Or+fvBFGHUt60GDprB6uCgh0fVlmyahEB55LrooBsCBXIcTcNBWNyedlZkfM
oSMDK9AsABkmVyt0tjknehTatX+Q20FmzEiT2xWafR8x9TaSSaW40il220EryV51
R8rh1g2T67Ia4UBF0rA3BY2NroEGhrMtnml056ylP1bMFv2dAiMiO7z/2pStjcnw
QhbR/ShMyg9CPdQPFkcq92mo6lElJS+MdywAkp1WPwM9YVGuP9vHR6wX/PzdFjsA
ej+GFd8NoNlzgE7DSZVhQDL16YEOKAODTCzGMXGX8ksrivVJX0clZjsm168qOIXr
HLaTvlYjygiRTe3RbeeGpSsl+2sUiYEqGbl2dLRyuyGC9FWg2qAyV8/Iysy8NczP
3esSsx8g/JtGAH1rkjFDEWCQi5mWFuoOq+FcORQv8HLeFCU0L314juBN1SvVWanx
QOg+6YHNVnFrOw8vrtdHD8Wr7Hd+OQXW/kQmR3GYX7xLL0dTwtqEnWk37qlqn+7f
xFNCm5EttFo/MzGliL0PbjLgeFyfunfMlz0VgbajU2nQdF+SRoDo8gyLKPmkzDYN
aeWlKrTGkBK9cHGbVesvSrQ+2fnXpReqa6zqHcllHOEzt6olI4ETPSepCyqbMGs4
UuBcfLXld7XdMPdVsw+Z8COE+I7fqd+5Jw+FQFIRteZLQJ+avj78/ZPS+wvJ01Jn
LHG3NPa4N2oSRxnl/vTGTFhf3q1djaDBuSQ/sxLElOZQzzsG71OSyfaSDBy97od+
uVL1IY049iB6r+opjwBtQh0hjKOoHX2rkBgx+xam5VBMGAJ/go6RCQOwbgX2wpkJ
5g1RVZAew4eqzKn6ZZb04uha0FaXD7Fzdvunxdw+bz2dbvC/N5BuJ84vhUgWf8+n
pG37hlg0cxjeN8kxumjSrwUpf/ryl3d5O9QbM0qGskgICpn0K2HX6aj1BjIkRLr+
MhEURFp2E2d0nJlvrQfokey/cRQQObdTKapnUSLzcj33oNB/yQ1hpOkBvSLjIQxb
dcXoHnDVOr1gJ3ReEJKG9TnbiQJclRvzAJ0n4N9ReBDf5UjFWqLerI9/yA8bbIDj
w3bTu3C4GNsfgD41dB1yEmk4VF10Vbf/6iBSnip+/BJl9jwdx6XQQw0slqvWpjDJ
ilcKv2o48y5GgGzVQjYG731jtZxTgs9+iec5C+MYycbceu4qBlyByG9Nn5Sb31CU
r+OraFBq2nvduN4kFt/PYcdk2GO5BHV+3B0A4Ge6jZ79oyPobOIuDZftZ+53hoYS
7z4TRqTyrWV2tjf6UbOweZRhX96n4hM5mNDGoCg9GMxmlXGvHL8ApJmWqBH3XfAj
sLHznWlKIxv5ESVT7T0fX7vI6FwGoqyFZTZ78L7389Q9kF3NqIcL+Sm3UJsQSdd7
scemjcGr7jm48hvuFjGWSNQP8oeC2cjmCJiFbM0QwnSJ2k5PD4dODBaD8gyIryUb
wTSQ+PY2Sd32LRyayGUGDTXIa2UAlf3fLWfqpNgi7aHf+PUHwZnWTZeCecaxXzby
mlLWL0YoMSQ+EBwxJtvtdZ1mH/ZZkgGDgRbUiH2HsEmvBC4mDhFUUj4QTYrl3YRY
QhWLlAEtF2RSvEbjt8FlwQeBQqUdavTCfhXnmOMc/8MX8HzXpXrnNznT/RhICygf
aSrhu3pisay1oWMHRuHb3F7y2yuL2bkpAA+O/5XSaSaE2do9/gTEUBipRp0jvbU4
hXucuyuPSPRVlZgWkimsW8UOmTPsHIlCfrgWJElJZaL01hSnVHrNpnXdR2YVw5si
6CRa+Rro0J9+XwODOcIzswr+01PWKqlCKl+qSOrmB6xeehCAFEyeM3RSrQf3RF1c
7tiKf2em7Q7z6UZJgcQxZlo3AP9xMyuKgxbkznvgDy2cXN4ZSU9ATMTIUOgf8DUY
eIivdYHuuWxA/w4aEKz9Y2ZWrUXoP+AX1HNbhtM6KCmpt3Arai+4LRUect4tLSLU
8cS2fVdnXrVWOK4K9f3I08b28zVyvEMhdhrGelMgZTACcu6mBJwfZXeyNrMGh6Qs
9nb/dPYaXtFQSamMRYiYWB0oEitNTqS3N0d/f8TBhmhIkvyQCJ2Z0JZVnJXTT8/J
L8lL1+k/lQjTtPiRyfjtpfnE+oiee0MYFpF4MLRgo7MBeO5JPK22Ut9ujbHXJXS7
sPUboqPvhRaq3EcaZRRBl9ZttuPUdZaezRCacIGtBqJGOqPmHqeeLioJD2sQ26XH
VAePCTEclKklaeiRbbSrJerTjVYWA/avpy/tR/0yEQeHGmJbkVB9OnRe8DnApLfJ
z5p+c9l0nS5Ja7KjeSFy9S66BJnPuTf/gvFBpC+zPUxeeD2L5xeqQjS8Pz76ccZQ
GfFJgut1HPf8rVVD77+NXWMr8YfdfyapKcykH296XVV5Fn5lo6dzxASRw+iAFsZD
Gj9RMax7YJit+Xe30n85fa1ZGlctvdotUiZ8LnqSBkCE5B1qBeIwsJrcv7LVIb4r
USjghhCbtpWZedGTIA73Cw9g/AnCg1xuuLL8MunYPG7olXoBXiA/ttrF7jmqbIfT
LyPaXFrs793tpf60+4MAU+UiNPeoSzFQFzWkbCwrRDBJRu8KB0lz+11xQoaM/2kr
Og0XNoUVfKHTL79d3o/qQCxLm7FCsKKP9HkZxvuIuPL46OE1/DWPkWOwsOnO6bo8
hJVsH0EZkGBrcXBTd1XOozY+7SXyDwTzG84iU9/Y+9dbPy225shi6bUv6UENjiF4
wtFGWdTxzEAKWiQAZ1JVgVWgz4JctMa8nlOxGYnMH5ETfbJw3VeUC+Hd86Y9gTh/
jLc2EDozYeGwP0gruLX2v8eZhBnxheRjTzT7jDfwSnVV7VwYbFlFStkc5dsLR1XV
+KmccvQSXuy/ZDaBNDSGu5/WM6qG5MVI0IqYRZDIKJiXPiwfp8ikkNOHQqgGuFK0
uWTxR2Rq2SBMi41IzZHuXCvPWfPKo4v8bZv1YRaLYvf+3bglF+TCrYfDl+Tt3Dbr
Jb+KJ1ggp+m7WnmMKYwn53xYQjKD4zJ+3QM5OArGOzHDxLsjNQtGruIGjqzFfjcc
5ZpEiCwMyXEJ3EDMlFzhYbflVV5IVdc4rW1PfnzzCufvdjcGBY06jBPHtoKCtb4P
IeB2mc0CG6TmDNLr6zg/aY1+1ZGrl/PTYFY/xsLt+zrEpXXPQnTb6OzXEoZZo5f2
AxdCuxZLq99tg4t0v6ikKQ9wa2aseDlQjoQ1nJBV4R7SF3zPqxhXVqf93xvre+om
zTSDOLE+49sAC4aVH9/IsBoupxBUZnfKoRn6zpBVSgx60Z5k+p4CUT0qUTJMWINv
lduVfpWK2mqdeExfjrihAzGREcSUioKEK4RX/pX5dB2PmO38613yI8x+AayqqxHr
9RXYgOhRsGOfqnBB0oG6ZRXow1U156VVwiVLEtEBh7GizpiQ0D+SRHgGN1GNCFri
oApDuUkqIXwFcOFYt1ecZhNgKlVoB7KOBTxi5hgbJ/ZvKHz8D2xHBRTb/bmuRvKd
hgSBn0tfpJleK5OkmTo1NsVpXoGuO0smHnarJhOlR4ZgiIDwR6sa9eePbbIWUqaE
pgmmlp1njprjeT70kWlzCK3EXoXLfWmzZVi03vqHBuRyjF2kFS1kXfhQB0Odhu0O
qJfwU7osfgx6eBgR0/O9hWGi49ymDuHcJEl3LDUv7WMBRRFuo1SJDVIDhHgWdcq4
yky5t0dt+LGonum9zPtsKsQuCR6YAGzShOIVBdFZ5l87oHBl2FgPPqgGNQ3N3sj/
JecngL7KP2twWzQjir021uTH1xh25PrLAOjwp/7kU9xxTW31NZtp+0UQgHsJu6Hd
p8seE7ZdnBtTKmqhA0n8rSGRr3+J5qi4EDgIEVPq7/pH9QypeFuMIlJqHHLevQqO
V5C+5S2iVJFW9UBXKyAQpSByt5Zg/j65aOMkpKGHfo0MF2WoNMDUtxwXLYD8fNYK
s2wAvAU6rMyMbvXf6KxuYbP9D8D1r2BL2Hh1+HLT+S0KtW2xn0RepDwHna98cK3U
ngWVKzZjmh5oB+sjf0fGbHtCzFe6en7vgfJiQTPGOOlweH+qyrzS8XceeaptK1VU
hNWqIAkn28y1ghvSSlLo+80Z4r7QfQQ3Hrg3QdLfkR/P5GFGz5/tDVoPqlgvptYw
W+3CCQxcqSgWMhXqs9CNXZ/6XTL9e+wImZRLisZWUgXZWfZyDMGC/hNpSkRa/XCK
V7QDx88MycdtsB2oTizcVlOpqRYlIFogMKImIBLBuz2/vSo+s2MPZaDZDX2XQQf/
MoSr/o1wV+4t2b1PytTEPkKEGqN3ba0HT4UWoBPtFogQvmc7GDLbSRIO56+Xpc4M
qMWVli5Z1UMbCkWD+82UOKw5kxyjwwBdVsFlEESSduG+Lts7UJ46HQ+gxiidVwt8
ksXNn3shmdUfZTdMsLCFHZyw4Qubx50+Bx83Gv0Ga9tRB/SxafiFMYmK8L/PgIz8
Id+zVhyjbYGquBqODvlRr8p+XLo7FNEIYwPDU7ivR29K2WGLSOSvBIPvO8V0w7ui
AHhxLZhHZ6O4lAUhQ7JKAB6Jc8432/chzNlUWbTQMSkCndYOta+ZFQ984O5nZ6Cx
u7cewB1Rd7gTe0pTb/pqox5vwa0wEZn3NCW/oO7lUbXFVw1m7r7avcbZqAQvZdq8
6W+tUpw+tjj70F04xC7NpwbQbm4YwZ8ZwTq+2unaIxOVOJOrvlNt2/WUwo2jXIQH
fqWLMmpUtiq1bzthNcbGogjzxjVpbXWlimhQyTBCD/nqeLM3iliTwvuplMqZmBLy
uffXsnjpwPBMs1qU51aK7GTsZcl4QS3O5d6hvuBEG9q3DjyPafcGDfqA4+uDVax4
R16nKQzLyGh81XD/jDWiKlGjVZ/8lpVqcYBST17rm47f3FjgPsNuIvDBCzcrRtBT
CR7ERyPRv45rMKhfJF5WTg3Wo8xt6Get/JEGAg1/3F0v4SLtchdscMB4YxaUASOL
f5VEl/B73I3f89ArSTMLwNz71PLRn/QAkLAa23qwaHNO0eF49dhjvbQdX+N2CHyv
HySQFU1K3MygqMH55TXKsyMbxuR8TdVHFfwvQUt0fNR6A9PG0ubOet6dmCxdG1M/
cHvHbZQ15P7bUWpBDonsyDrVazGH6uDCj2N7Ic8t7juFk0XoqSVqZPWf8rKDJKpI
4DA2Agggc3NvMeTb1k0UzM6DD77YtKc2CBR1/MwaXV6LOXEb/EoNORDoql8Ck3ft
Xdht5Ug8AmfsvWEvLFeC6BtURX36x7L6QmsgK3nk3zM7NRZ45ICZaCcB6SO+hYnO
7TgBcfXC8LB6S/4qoa2vaCKUNFMnQBxmTdSK+/q0Qn/Yol0KribosMpDH9pgwvhj
k8JWeUqPMZzC2tJU7K8MOC5naWD6EBPp+oTIImUdOTbdtbXQy+N/OLv6vXmkgJzv
ckElXmQJckDhFJcPwTrc5T6wN5Cq6ButOLoigHbOLdwobEKciE6hJyciBNODnuJ5
2OoejSBkFSizr9vn/tppnCSUrdJFSjklkp0x4B+g5CeIRLRGrdp9m1F3vy7HfblX
72FfQsuJ4L+hr5AWbnb4Kh2cSEpFXBZ6vfPt+ASagzUGHLvlWT+czdGlHS6jmZ69
zK59t6HFGZjvmgRhZuqawmT3gqLcf0Y3NA7HsLuK6+UidubUEwzpjJp57pooRK5t
jQYgsC6BHxeeBFayfRrDNKWk26tdkgScznRynFVbbuYc2XVBi5Rvko1QVqFWdQCi
yAAuJJA2FZTKnq0tp+tN80hhY3ZyLW6E7neW3g6AtHyo2ftRMeVyo9KyY72iYtDD
prlY1tKADrAtfToE+baC3Q5Xuj3qURUe+UVrBzLCOarcLeote2Ncrq+U3qyoOxbV
8VXXlWM+n3nKrEaSRgCwdgyKG+S7FDA4cyaicsWgvmvvD+SqNv1/j2z/kDe+r44V
Jmtf0fPnRJJF4xNbpw1gF8glawVq2QiokZqyF1SWBK0Uk8gL+XwjtmnBujSUg3hb
sZ0rUJ2cUZYsMAaECIN+ryx1RDdGT1hbM9XLrIz89dQOFhk0qBBwBCmeo41v7ORJ
RhebWtLXTBGI2mlz3bn3C9QnGG/Au2WHZerTq3toXiG9xA20Tp/t8vPkcDrjTZyL
WlXhCQ2XMZ6OH2dQoDri75+xq93FiNyk5Epf3pNY/2fH5FTaBDDKHXwmvCEOjRSr
sMcIDQ2WqoruzYHDMM0/tn1S9EZVJOMuIgN4TSPk0e7ZON/1Hso+TqQoSHubsUJy
0uYwDNFI+eUX99aAd374KlPiTtX2SQwqBm4TXVvqguCNiEMsvwjVv7m/XB79ek5n
pBuZp4LkvCtt8qmWg/JqV+HlJeFQE/sMgTeI2ivc40dY9m7clF0Shyx+gHADyMsh
qdQG4JJ7DcKmhkxotShl5P4go7VLF6GJLhuVQfnAHgmYhvRstEjHxeDIrx3e0ljt
TNOciHo6pPseDpqDzSXw7xcJfRwQkUwgh8srQFPKzhXuP3jcTtf8vLlCebya/H7I
BBF2SdkpslBpyLoeX/hpw6kVcOOu36vh/DwkLV0Dhll3N2EKYAxEwWgWybcJFBPd
0gEOUG8Gc6neWYrC9T8UCjy+uBM6IBo5e/VWHrevHiR4X4bksThqJYkXogmWc9qk
V5KOOeeMXt1FKtkA8an12WnBLnOoZYf9eT6B905zn7yodVnkstGpPlvBM7In5Nzq
fZ2U5dIl8n32pc4KneXpIptlmF3Zlq/wVOLrt1oSPXbxwfuz3PoCFC1lJzNWnLPX
AoDWIlgtD9k3KUoD3j4gXyv7zkLkN/5gtSNbLgVW9xomP9ax9o/6ocymS1M+IInt
X+BjWXBbBHBM1P6DkLxCSVfm3dxpgm4KalAFjrRYyQon5iXWcLYnmt1hcHUvyN5U
8jfuGpPd57xSpPNMqn9DAf3TNRKHbo0/gI+q6AVjgXISP9KCbxnqw96gduQSiI06
fChzz+Ac8zpSr7pDhmrSChYMp7zmUOgi291VOeQ8WbzZliDj/+xTcvRVBw1QFtZX
B09sGstwp7QEZwBf3DXja0fC/2OIbFXBdVWd7VJJFvSf55iET5n5ZVHoguI7xiuL
7mtejmg+nitu6kgMohzKutTZ7UEjvvioxr8ra2ANPn42isKgn8oDlNJODDZ3biXk
CrAv/v9pWRXgnkgqycax3XbXNoCj+Ft0qKYy8gdSr+C3qt9vMBR0UTttCxXJUCBA
DHir+1ZAzABlo/qoai/g7/gegMtys2XlVLhOMzHaaYaam1aJ3Dbb1Yp/ZfYHzX/A
U3a2MYvAyUqzjRsI/ytl/V0RV8Pzl7XBX3ZIc7CXRKGHiT1t/Xe9AvVqk6xWonI2
/wjc6vItPe6MZ+dD9Xfl3zHfsH64b7KSWHxrRzeg1cRh7jAxVvhh50vfPbYQMUmD
rNhjsE7BinXKUtHLdE4pf04yRC9KBdh6JPiCg6PUyp/jfORXxaMToEZH316UdP2v
9tIL4aQ3ikdvHScx4I37YiRx7KfSTzRJA2DQD7+7g+SrIZxcWSmxSJsqVBRa/jq5
Z53GZEA0jwSY6Pd8T8DurazRAFGkxWJJD844/efiJjm1nCsQNn69bBVsdkdGywyE
0uYWD300QXSXM3DBVK0mwMOmwOjySxZ0gDbbYuuztQC8R5GGY5T+bDT8UpJ6G3fU
7OY5+YcQ+bAHyqULBoBADbuUsIttr9SSkO9wVPF+LZFOzwCurmtYVZJiZVyRfg3l
qiiotoYONHMHLP8lZ5eB/zri2tizCaMPTwVN4B4eQE1WfFpxxY0Dk0it+6c5PmcQ
7ENDpT5uBDNc+BLuRXP+5LOdw5fGZt+EuZfBxM7PL6wZAw+GEF3DplbwVBr+Gwb/
`protect END_PROTECTED
