`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RyhpaGv0SUWDzAp6lG/Jgw9jtqwwFldC7n3aHbiXyLuXkmA7+b+i3wNYKemY9XiU
I5+QOi+0CcYLvNjAac8DggTAUmRJaWUI8oRt4Kw30dHJir9fIQ7+1S4i144nSdYz
OJeIkoh/sUsxWNTCZgtjiL+SrCUbrhM1xVm8O1jrgPU5wbF7cVpW61SWwtbUBova
miIoUlB/YOupdfafAzOepkVhe8uQmDM1XMYW22tOVTf1UOrHD77ZJ7AFmIWlWye8
DG9nXZhxht3V0Hlot1G7rQe7bo9L1CTHny/2s+XfWUwdyz85ubkLPKDrEXrAZoy3
Qm1A9Q/Fho62qJwTYTlC/8EORPreuzVSBfW72e6PsEIUH/RyebTu/hjb5XerVKb2
JyrC/lf2fVQvIWcQLq9a1mVQyQGcWMBepA+sh56wDGAOTtfJbf9JP20CC8eefy6/
066tmY71ze9A9GK36Bp/32ihE2pyHL3z+3Av0ZGhq+zdEChy6zmEvvB7NsWQ+Ccm
JyZMM4qxVFR/iVrUP/Kn+qCoaOvztGz6gVampHIDKLSqUBbYdjql05EwMa6bFUH3
8wKRP87N0ST8boLqWKi/NmxNZva3byDqxCSb0JNc114sqmVIaFyKvuSHFU8YZYqe
ahU8ZlueJLJ1qKeX3p23pvgM6sEFacD93ZS9xl8+gXss5DWYvKdz4AoWOg3omds3
fxuwknUqc8U6wE7j+lIONjM+TADShqkLJt1MmI3LejRalvGkDZFSNZbVxgbq5kPY
qmU3wB62/9anBUFNPTFQ0gDV3hc5LJNXFsWHfiS/zSmecNm+QEs/lVShK2u6VwDb
02bjqJ0XUAmUnDFoKPfzVnoXDRVSLua/EkLAnFq5+iWVHE/JvEQ3JHmh0z86ZsuN
K31eyaJn9cCEc7hog2pzkNJ3MnlaQTXG58Kng1PDer/NvPMECUKDyzcvQHMx74Lc
zKv9lUxBzxtF7vnZJlmzMoJaRP8bWbj3pOXW+LJH9u6XEjuus5TvaP49z8rXEXTC
g43gnfQaepgqBGhxAVFaiYMAxdP+Cul/sKSNnlTUnr54mzIqG2Fn++cTvv+EBchX
GSLtXDG3WMa2Fzzw6iIQUQnLpdc7NkhNmg9q3WMnlYdYAMB79LgneHIOJX2ujBzE
eEDk+wdrFUrfUs0j6XDaTLfyZguvlbiiEHl46IiJg9sjHBpf9tn+9RYDfH6cUVre
irSwJEfxdjhJX/2ee+TaW9O3Man35gkpv0X2xSn92xpiInLee6h82lTqI45VpUZ7
he0b7nVnCEnEaT90GVOo5tH++n2u1j7u+7edYUqiWe7Cz9RigLMyxk1flSzUyfzn
Fw21bm4zf40oEsghzfT3QvpVrUqkslTTfoSfJMXIcw/nrXdS4SvT8y4ULtcMSfsR
7BOsIwNHiUMyawcxiCEHYgAxGSxr+pcwEmwg5WxA95a4pycM4NEZgzJQJTPvfwXD
tSa+8CLYBaTJ46/LM1IrCIYc3/F6TO2I6BHf3DywAM6tquzvEW7r5SKBGoWF0Qb7
t3ZiSY6m/c0eRsxEJ5NI8SWuMlKBBwveXgiwDnK0eAEn7h5kMIG3wZYd3vCzH+5R
j67CuoVqbwqnxpn3Z1UN8MKyOnvoZzoHGrzlZYPsETDvxgZqJHsp1UYFpsNJYJL6
DzYCi1SiPOyGTyNGR4T034HJeZOiuREmFy8NHbLbwlPQmazX49JS6eXcElnUlf9S
vlwZ2qG+znaC1ImtGb91ysji1T33jpff85+DY27q49sSI06ajjAP5aa9pPDZ1vFY
oFqgrBxxNBzH9DNN/VSncO4Bx3Mu3kvAzNwnF7ACFjpFO7tXDk8srtmITugNYXq9
T3OXYbnIwH54N7ZMU9GDc99G+ewj961BVsVU8NykCKQV4Iy2NAG/ih70C/4wLEri
dmMLVpHR2n5monnpcM/uLJJWGau2r+QKTcKFFVip+vUD4xEnfXbjhoxZm1s93Oqb
Y6zZa/k48fEGIV9yUvvfU3hE3XG9nQHdvwVwz7SBnqEgG4rChtxKAnz5chhMwvLq
4j9fYmTetWCxfjKQ4ctxTdifRXw70xldBhy3ImsjWymab+764d7hmBFScKE5hoDu
A8GGgG/PKC/E8zc9fvWgTOHwHSeIpnHy5cQeH+sP6eW/pIUoTdrZikNSCkDekMUf
zkRsDXFWP+S/+e9NFNOwIybcAtzxMzmhyKaB4YV0TlMhHROXdNICYTZDQiSVRAb1
sfQow6gg7RQbl+j/xOZfl6sY3HmP1h1tzpO6rJc6edGJfFO/EFej/p5zwukXv7Yc
BIomDlZxI0qXFQ+0902s39bkgNb2nmZ0ctzvHo68SYPgI8lGfbTREo0pzvL7SSZ3
8t/UhTDy/yscvf9QFW2kgfnAn2YaIOXcefEivc5zCbfJ0TP5pq4v8yNQ/FY3KnyY
zJtzvIjHtpfHSfJhWTj1DzrO8eiZFY+tEy0T62R+PKVw6YlxRf1oSdjLo/B6dQRl
7kExXWyhoc1hW7ehAQ5/pNUTWc1CQHAYAhu/L38hP5poUT2qT4AjGVeCWRSzMjy0
llgqYgFFr9KBw/nMzmYDSF6kdw2LfHzQRFkfae4yiaxBkzn9dr4iqlloFdRoPbjI
rV4NiiV6AsIfsdo0JYi39K6xW7ANPMPHa17UgLWwwgKw6MA77weH7IwwBw8sjIYz
gYtWV1Ufw+gX0Wgsi2DxCinK0FaN72+euTdmgmNGqr5+btB7Z4scJ6WvOZLdmbcz
nDuuh3L+OBgge+kIgeM4oQYIHohvLJJZBWPfyUMvW/ZVdKQf+9zX3IBIrxxVc4EC
zxszPE07Cz42hC/WHX1QxXuON16iOYCC4OZAS2ypGtVJPoCTh7EjQml2pQFGihwA
FzTxyJRTzllMiM6QtEkcrNpxgR4QczDISWsdRjBcOQNyDPyV0JQcuII1CMAUeKpa
DEK4fc1cIETvOi5+5+9UcK38qovDNhctuQLAQenrYlLiJzq1PUrLBw9Hp9oUarjj
CDzFthJYj/OJWb3T4N8/yObk2uDXRMqKfU3DE/F+bBhzMJk9ZNQL5pzdedgfBOFn
k8pgu2T1d1LhBo1Z7nR3RSvi2M7dJQsacsGjPQty8k6PHlY6ktFWkbpOGODcnr7r
PnIdIsNZqaf36TKq74pRJJHt2kXzTiPZojfTnn105FQituZ+WNF5JFk1CfjUU9CB
cqt2qzrrilm5WUwReK2G3w==
`protect END_PROTECTED
