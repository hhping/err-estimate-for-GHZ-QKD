`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I7cDpGl4LNKG5GblvdNTHK9M0r3q0uROJqmDwJZVK/usMlMse7rtL2XEEdG+Uy2Q
EaLqexhwRF2ZIRIb8leOkL0R4zgNQl9zKQijbnO/YVEGjM/+PSEEEK6Jor3zFXGL
v2XxWYKOt02TCVixtBBCU9E8zaENKE3HRGWqcr0C4NKOyiWkBEsSbReK5CdF+imn
8E0JwuHpcMod4nrVZmuTUaI/g2fha5fEyX/YK4SX9uTiEbbkouQXy+Zm1uS7Ixo8
TtzrNV/5IYwH/heFF0WgHh5O1Gb+116tzszo3qqLP0IITdi7KVx+z1zAfPaRdCjr
4LCLwlSwi33eQbLTFEc6l989j64C4JBysK7YTYmrYMXtzTpQ5theLS0Bm9Y/oarv
hYfrGeeLayVn6L+l1TnKY62vpCGiUTfk+812JXsR/3skwr/aIP7pNRpXagr5PxK1
Aqm/3JVsIuk0Zh64wIgb5s7tAvpEe7TNAkjN6tW6KK/xX8jDCNLPmBclwfVUtgVf
N5gC+ch6Qd7gt6jpzQftSJji6E6lYSAeTUGfa5kwlh7aWAOvyaedv6Y7X4xTbvLo
vVVyblAeh1UHvFsCdGNthTVb8tuSmH0ulubsMNPFncl5p2OoBO8OWERLf3Qj0b3H
vZQBU5kMu6bHhs8tWOMQ3W5cy8sfVHLESicsIY7cnmMVj/yyAkPZuAvUIqoJEeei
F0y2kxHti8ZSMY6P5P9K7fx1ywnR3UibtNUoWgKUgKsVc9Y/myd1BAXYwdN9fNXY
Nl1mp+vt1GtFP9vkPjs3oKc8XSDIFEAQGkZok3eVgAQW5F6Stik3ot3eiYUD3GtT
62EQibFr6x5Bne4KAMMUjAJ2XUJe0NcDuYP7MiOu4dStP0C704uhle2oRVi8EPyE
rpzBuiqlemXXBKMsqn5X6cHOWhn/C+3rn9IRmeEeApbrZMDaXINKqmX9qOdlRz+a
uceKc6boRgP//a3PBql21NbPK7w9DUqs4H/yK+u5+cJzc1g6Gd+cTmAd1T4tViwB
UdtWp5f6k7sVGxyuzhetF/Gyf+bCQjLuTY01SgjvnzFpZKWsT36nueM1oSGR5Pch
Eugr1j2XU4i/x/UsL4HZzbgGecqLSfgSdD1CEZwI5CJN1ogQu4FiftP5d+rQXcwY
CPhYAjtAuCKU/0V0n5K7PO62r2YjguHTWgYvsuBYsdbdgcjfwjlmQcpO8L92JFVR
7N12sP1Lpm6QY4d0/CazlxBQWB2q7LIp2xbFks4GeykQ6S086O/KPp32JkwGDssD
nALeGQzjXjZ068uR2+xs/rW2FM9yFDvFfsv8nxOITYtpUaZ8GwT/kXa4MtMSMxgb
WImxOLQ1wrQh4KqZ4JbKwZ59LeX93WB+aCzcRJcFRgxmY40NGjlonc+h5qHqwgQe
2TKWHo7PBvVTWzfNEpdT8P60YNO32enAxQFFPc6GAeg9M3HaDf2ul/03xzUvYbCn
F3RLthG27fE1LR8285qAtXnqCRavIlnjl3tEER9+MT2VtvmyYseeP0zXI8vBz7In
0TdIgiNK6obghfze0lByl3dzzciilJswtGC78t0nOx1DeAw73798mQFztQCEack0
Y6Iwb4jP8UPzm/r4MV1by86at98HcKqSzzzPAqJd9mDml0vrglqZAyDnoS4OTWdQ
ql7sWe9lYlikncqBMI3JNt1TFse7FJ2SYuTrGMoethQocKJZJu52WpJWumd3emya
1GRm/xjAx5Se8bVPqPer25YRS8iYuAE8jSvs5B0fMbs=
`protect END_PROTECTED
