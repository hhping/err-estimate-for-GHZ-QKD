`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vATQhKLuRwiJkol2N4m8A2ReXsUS0mqbuVR1NViDvdP3OJNLNWh1UHhkLHUH6Xu5
i8vu0OvD8WlpQ6tBf5aqZ9kSGuOsdR7NJKRKXASS5Xy9cQiK+Y0/EqK/fKsXaNNd
t7qxH49E+XGiVTFnuZ9Ynag0Lh5X11dhwkk1liqTiKjW/BAQPUCRlM4KpJ+KhAfR
Jh37HobsLKX/uouer2bZXYB3bmvLmnlaG/uJavVUUHhPvj5IWfm2beY4ssq1iRei
pUQACKqaghhT2G7SKIb8Gvpb9b4/Si6kQf/QshjS0ALKi90h+X7G830m/z0OnVHA
yDevBMIWV5Imsk665G+2CISEjtnxADha3bd7oMlQ1cd1xRNj4TPx0JGgEZz6lLOw
1/lzCN7vqjlYRaXJFS1wo+nvVMxzHWQgMvhmkV1zHN3IugOs6ame/MT9Lhekh/J7
sCak2Qrb2EAP241qfWhuqzLDvxytyTwilP2cVliR0UobA1ZP6XaHkK1sTMBQqn8v
GQgs2qVi1eaC1g8C/Q0ffazKGwTF7NGrKWnR15zyxv+KhenLJg+Cmc+iN7NpJQrI
HD5GhISpTUYatcH3PaKRzPeUNBjZH9KUeFYYInq4khcep3SiMBlJSZ/ku94PpRnj
xuXygYWfXJhdgR2fHTbWC5p/GzunAuBQ1iRG/zzbx1e/TwLQvhDJCx3b2YOlVDgR
Jc/K5Dfq+7q0hv7mM1ppgiTU89eQ1s3AYOlmlMy5XUb3bWsPyzUXLoIm2hSanTmo
zakbAjA7pjTFT9kqa51TAFzbET0jNxTGYAWE1u2xm4SaJq1iMtsRrO/5rgvQWPQS
THHRFxQE7vlPfEegXGoTpjoBTKuNEQ/ZizsSmLjzXbJePui8ans7BXwaMLSwZC6C
4b9dv0C11co2a7nRw01FD8+vPo94057sXjx5ctSMRmReJ2UDYZFGHozM3JIZs+Ob
Jbxz/y4iqelIm/2AvCpSXxsaKCXx4NAq2ZPdvcDKWWlZgIoM/BNQGjtvwEAd9KqT
jehA0wGRbDKMsncAmW75DLFmteEdbqK9W/wWFzYBEpDn2WguoFAWzbYF9lxpvCnc
WxRF33tgK+K+hiWRVyREn+BxpwlgWeXiJbeuHTOOYlMHdXLuj28AA1P4XDNFEYtO
ZwrKf2iT2/aD/I0mK2a8ejjwWNA+xY68XLEU00D49vaVML9c7KR9+DLEtWDFaawd
ZeE0lzHq5Ia7HPh9KzMveICkZStYO2aX4aQsoHl3MkFpVA+RgN1n/i41NNPs5K0H
Vv4kFysSfZhggQbZw6VyVBYRvvPBh24aKund5RJwQs+AdLPW8thbI0NBzo6c6VOO
u+DduJ9beRuMWqbpR7GpPXgPYY0VK6Zq+qxddYnppBWYKgxnWJjm23hMMNzcwdcQ
YK8b74pTkgdpLx4CGn9mCpXPoH9KhlQqemHGWoDz/mXlIMowed8ckyYwy4qu3EMQ
t8j0yWYYOPY5sm1WFsspeptrtm/n6MsLj220fn7cTOl+bEcXK68Cr2wRtu2c9G5x
PEYm6KivAgvdsyAn3HnwdmpvNHQY/YZZ6YDLhVUibCUvyyzyVKzOtuMqPWS5VNbH
qpKTvyNKnDgl79X2OImP4WdI6SkU9Ef//Y7vTm0CJlbWZ58B3UwSmENYBoHFu1se
PCseTj2aKVxO+qxa7EULu3WypJwPjt+aBkUSwSoTcZ80jWArhzGncIxEXSKpok5/
f/U6Uo8iPMJHTi9hb8YGEEjVubS00RUQs1VBJd4K4CbEwKjCy4+0tBrG6rJ3WPz2
oZ/05Zue2I16JIyx/PcfciaozfDm1dRBXdOqlsjJ/oFAATNpe82JaVf7cJGFmU5t
V3aD/u36Py96Vj7LagFuqAErEIpZZQHVDAppJJ2F2SXtrh8f0zuRTP4RNliQJzsz
xOEsnNwpvAEVPAbNM2ohXoqemgI6HkmEHlqwdK27ZdR6u4AgXJAz0TeljhZn3m0k
fvh+A47iioYRJGh8trZuWVcKPjDjFuvx8HMwxFIkIWoLqaq24Gscm0wqOqne9h3Z
9jgSGLREc4M7uKRbrxYF3IMn3PFTA45OdcgKOJYdFUCJ/O3051nY73bZ4YrvP6NS
Z1cJ4ml0R3fypN5Rf6lnvln9KCq7WXo7EGEYg/WKDJ/QK971Hd590q4YRo364PTA
SjCTFINMsHtK6x215ofmT8AeiVfXKcqkVKsR6Pk5blDPoT5qjlOZ3JTuNHUpEeid
O/IJCy6T6iw9lwzxPshaTOJ9/n4yB0sLyjey2y5+7cS6KpR/31VBsgLMAQ8PLT/t
dQdPRNXIXt3ndI1DUrJe1XeKyAXac+nYU25xqv/T3+xx0Rp0kWRUsPhDZtSwCP82
rt5WL52k9alozJxmfJRETGiAb0a4H4CdfesiMgtpZB55JkaS/vjBMimi9WArbxCk
xizzNS+JRxaB14B4Q2LCr9H9PY4+T2aAkZhWAtRESR+eBkBQWJuJey8zZT2Y3/Pk
RnhHJ/xOuDSP0jfULYWj38LApuiyFMQgHvVegn/Bq1aKbBckHwTVEGeqkZvSvQCZ
tsGUGhoWsMHLT0iQl9JAkL/FD/nvEf3HA6dnYKORjtJfZGaxV5AIe3EVMeTM+5sx
2LT71GeF+qJhL1141y2QzN8cWORQgOc1fLRdYQwPwJfW4ZZ+RTS86P7N/GGQvjiP
XcrKgr7XFLsCtn3u/6HX5YvXEM+4J+AQbj9+fghVmg2RA6Z8BKP8uzjtBkkI2Ps8
2vkpOLC5wD3Jpy49266XC/7pW/Rh9ygy0We7H4MnZa8MCCZqLVjikwYQRJ94p1WL
9Pk1YfJKmbEeuTKsje+4MnjkSHRq/4xaTprHy/p/gR01GH+icRNHT+0+xs5xgucl
Q/sCBYZPemEjDDB7mAbhTepN3w28F3Mv3MMKpqT3AdODceKv8MAgzmwF90RDljZO
96KTiyWmGMREdcfyif1qkd9z8XcMpBhzEW8jGvu/IW2HKX8bMMknjUQBWY6pIw8b
PqGHPD8jGrIZ/qP0U2eFXD+NV86WlyC6c81bu28EU8/ZgP7jO4R0ZzpFxvBxCa5B
81f5gbDNaRH3AnVtxmiOyx3j1Ky3V1HkUSxHhpErSHCANE9QkicFqrfL5Matwtu2
mTfCk/7bwsd7koTXI754xfJ28O4xov54c6WQSyG8z/tFz3uYxtIJQLYvj9zQ+PaW
9MMvCU25S8fCrNTfDoZZew==
`protect END_PROTECTED
