`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zACqoTs+Kd/9ygbwArRPmP29Z+I5kkEWoLja6hhqxnsV67X3W+l50yt0lXlvoH4r
W9XVb3SF2AkA631ILydQdCj18H3G3sXh76nlNS/Zz/YxnSwdXKqvqdo0iGNOKIOt
4a78LdRnlj42/nix/qTKykGCX+g9OtZ55ow1nsTG/u9T9TOXaJBiO6tirL5wuTeF
pS36PkOCuvLByKz4wjXq6JWAbeA1mSNro/OQhVUi6ywM74UBjz1WIURaw1Y+s5yV
SNwvDvoK8GUGjYSYF7We5E6F7N+yRxT4i89H7aGgAj2bwjhI3tgfRwEMnLTcjusD
fe4+n3jpZULSUhkgV7tEPzOp8s3Z+fo8m8gqlbxaM3GSg4aZgINV7OVmAr6x7XNW
9LUsIRff/BkJ0H4QCyZ8b+HoTvV+yYcofOhNey8VDz9ncJtKdtZwv8hY3ugDDJ3L
eiN/h4vVkIGKmu5l2QRFktxfkgy2/iR6nuFYVh1ZXCuPoTCfZz0omvOnHd/phs1m
0ZeWyJUsovEc8+MqmWcpVhbSaodSZW/enKuUU51Yre0Equw4ZQ+2K5wzYuaz2VuJ
GGRwiCWJDnJHdcQPi0x5sOO2c9y7Jc7/fyv0O8yHGGR641ZkaDeEIW9lu+b04l16
LkZ2dPn7jBMGREU24mVSZYB+gX8bPKDzha2xzrfMbmiNc8t8OMbOIAb1xN5y7TdH
te/po755RYEYvee5qlhKEZNyUIHs8oT0zy4EJUOmLmIR4Dx+9RVGcooV4SPWPuyG
b60unnDgHwPl2hl+krN5mcXGpfkOX6PylaW3wJ2n1XN2+6CgYHfb57D7DZ1XqKLg
j8T7Idqj0Iu5OhZ+BHCZ/eVY6A2yi7bUhtQ46Rib5WUom+GkeFRxMB5AUyIHmJmP
6eTfKwH4rv6tmR7n0uun7zS2jBbfMsNwPuGHfwihdNXS6FjrsZvzOYWZ9AX4cR9c
GTFi+oswzensZH2zIHYR19jbEBVQoHO+UKmLGwqVzr2QjM2jsubvmprkG/0KM5iw
QcwLxAxLFH5kXKSGu2iI1F0rLaSHPL9tu/KNsLmciBTLjzEPvAoy1GINPBWD8TeG
fVLXcGCMgpThY7ncU323pxn5i+jWC8q/cCfjxURkpw8mir4StkbFKTXmGgRPn5q6
oFTg6MSOO2P/Jqy7xeHvC2Zp4cqyHTbgN5h5fe/REAJaqKeiUTEmD6gm6FZzf7K+
lEQpFsoCz6EkWyP/sLi5yg4gE+rgv4A1ucqkK9i+BdkJzQZlZTJb/2k2zA43waPk
wnStbGzGeis4SpXYV+wNeXwmoBS+TBxhP/CrnO1HUjvWN7a5qV96RTHJro6IfAo6
PtgwRRmySrKFGvzRzRb4KdjZCgJX7fbS2/pa4vn+mIwLzgdBX0efLz829uaXziIx
7LSkmv+rQKNfQDN6w0Oo/A==
`protect END_PROTECTED
