`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sjYLxsNBNnvnP8pFMKdsMRsqgNeHr71THYVGSw3ccnoJ2/BQ/3yWb61s5LLcF2Am
bI7iOpt2iTrzsMONJ5N8otZqN6bdppuXJ1Om+/xHzZnJ0Ns1RadIBYkxA4srEeGI
qQuyGz/Se3XfDw76EK6ElkbpkgArQUosVKcfaBSwt1/tYSnTwbyTtxv0ftb8Ozlx
S4ohWbUpPRhLGeVGjP3dUXNwNHqUVPYoo+B+KkHRPVCt05gQKIBBl3e/dR2GRruX
qpX18DcBvU8+up6c5MS24P00hJeyVNM6KnVX5RBALLsHfnISv0hlkZr5LLy3FU4W
mF1LPntFIX3+sHVpk1uGJ9P9UVEMb0gKcXQFdDRYzLztCT7b2A8+ft3xg5GctVDX
KVkrCRrIfVMKEubu2CSnSRh55oRARBi4tHE69sx5UmasE84brQBPhxP5N3V7xYYI
MTfRMDD9z/pGpBW9bEF+ZZSd2ejOe/cACsHKDbrbHl0r+12paf4VGxKOs+eE0BUz
AoJuQisnWPEQMI2OCUM7f3t2wik7d0Pe/Od5Y34C54Hly1PHcH3ePEaPXSp8rsyH
uCqKKduEAzD6OTwH785bZrMTcJ2Zs6iUf7n8KUGy9sCpT4iYzu4eIxO1G84mgVUX
P1L0HvqgML6TtDKEBVx1AjLdCNsJlV9wdd6QNIzempwYtvNJN8taO++ZnwOCm7z6
x48EEYIZBLdbKxHEgwGpaA==
`protect END_PROTECTED
