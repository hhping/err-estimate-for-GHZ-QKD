`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
49ajni7ZOv5Gf7uKw4BjSfXaah3h9n7BRQlz1ms4WH+tIQi8mOx7DxyaO6+bKLTQ
RRU3IGKU0L2mLuglB6sWyG+vp6YrS4gGVrAB08qTYN1o8UI71FhWVixmy+UCDgVI
wjbMKSLWz4/cR+oOOiErMVTE64xA5VdRsFjhHTsBbDx7OANT8XBW4Hu2gB4fDiMP
Lal85Byr3PkHRXMbgDtsLkjZfinKGrZBDW81XjVCm6uh5uzX8sxgLq0MlcBBxnGW
Tyl4TeOlYH3x79CZP0bfFpmmKULiAvej515QmP0wRad46993H4eAcpWIUafQAntv
emjx2ymmdoMX2oaF2lWmlElQbk1ldJo8k4ebZ0cbJXbTwZQfljRa4RgUh5V39WIK
GODS4yr+PYR8X/qaGsNRj6EuKO/LbGWSX78zk9SSuJo7rqelm/1srp6Jo3LsLQ42
`protect END_PROTECTED
