`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RmsbCCzZ0ZPnrBp7WRY9hrs/2O8Q9K66wLJL+AObBLTAsNws9K+HGc9f+ueAdkKy
NMqVcrC6bCtrSZRbPeowZOBNfgIN0gGMJpFsc1wCzqMczMGlFv7MInfkmZ/Thu6w
ginPXCjytnxhkJaT8EKFRlwilRaUy8lPKapLvxBorCrXem7FiuPEZ7nqvXj4Rp4a
SwXQsgJ1dLM38FPB0gQUhhcSsI4QcE2tXvtAKpPBuIWoZb28Y0RLfB3aUH/q7Lwx
q3f1OlC3ynncxvkKvaHbQxx1ef4szLy/4wL4dwps4p3bf6kYY0u75RUZl01pOiyy
Iz6Rg3zBuUsyw1lsGwyOI92ZJs3Onf99Q5ZG3W3Q9hqR9bIjxF02L1+hun9iZIZQ
53fXPgm7EcNhkwX2X/42EMlINk2pPhgBo1lM2mOVGbx+GtoCxfLRgpokdC65Dct8
XMVCj5K4MthSNlbDgyTocuYIbK2nFokICNDRKFoyQNQk6f5QcYSqlc952t1fuW23
X3NQ4heHN6cxdT824vXgUxzpCxBnCzujpkHqyiMaN2sPLrbyaxYerhDScEReRj1A
meOaoSm4yWHi2FXBYhsAbRyZnK8JbYPbihe7fU3QKai5y+wakTiV/pwiWoGstD6A
6qkBJQwv6tzXPdulwMZHgiFFtLL0b2IM3mEgARfvxsBpKgX+/f/HnppgdYs4Ctzu
WqQgeeb41gpEGzfLeyb8xxd5f1KRsmm6q0tT5dnm8X3UTd/Fwi6AaoBfV64Tr3Hd
YMoGauWqvLWGHQm1X0tHNN9SEeXZFcIJHiT2G5U8tGv1EtIsVxn90PXA3EH3jRNY
Rt2JpFMDLe7Pr1xC9TJq4KEbbqBtFzp8Vsgxt7yxCMOZbuFpR1ySfn3tWAWNH6kN
2+4XSHfsSvPvLrBbxJcf3f9dxBJuCVLwOgoc5y4/TbO8mw4vcbyn2cXRtozIPw3L
D0rghJcoja/DbO3rCYcaZ9SBWwB1NsYqfK7HOV7S0FIkBYzqJXQOXRfEDPNpnSTg
g1TNiYsmueu11oFAJAgqdJwBGaBHjoHRCuPsl4ve4OvCKhRwJRTU20jG5mPgLpmz
kPX4XdLbDZEjLRcQNKRaUDQj3fovhuK9CRyq+IRbHBsO+9CdIYDY+d5+1xA2C0Z5
CiILjzG0p86zfm6Xpnq7WeTPCNd3qrL48MNanLGoGP3F7XvKBIELREl7P5ZMciah
DYGpYZdC0tGdeeSWDueHcLhPYfzn/IIQuwliL5Xp9owfzQj6AsMoEkzv1g0d0pEc
d5BHZE/vR6EJ5z6xOW8jRnsosAKlH3LzE0RGAN7EnncL9DZvH8Kp1fZKWiEsLbzx
OpUXLN7VGlzjVXLmSCd70O5S/9HR/Rq6lgxU87DtkmUtjQ9c8ozUZsi6nOAmw5Tj
skasgw6EvaCirdEUgTNmow2TtuHmrRAtcVAEmKFyQa8P8zfNouDFJhgVgbkCqOsu
hD+js7rAPIC8e3FXQtZ5d7On+4ioqgIDBu3hpamiFfwgOAj8KZkz3D4j/GmEMeRK
p0mB2cWEOTSsQ1AVXFFOqOEA8va6XIVZJwuwIZdEIe7IPYdrSChZLXczogxj7URh
MIIP2KoXXrNRcX57viHgHK7MopPcQeyswbzMgnqZS/R+tXF9TbUmxbF6zr0k4QA1
p8ehXOajMCuSKNPQtZb09bKVsStOBnNqU3q/6lIv5VJ2Pghe5y24jwrDk7ieDFni
AZ/JP5bPylGXOiz3dNVf/zXof8t3L5QBEhSR4mAnh8qf6YlESFSZKy/FBiZNlGJl
DmaLtlNkelNDNXlwNmDrtg==
`protect END_PROTECTED
