`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WCxepyC0Ht359+2OQg2X6Umq3IFhPsjCxpNLU7VsN4+fSqqWquRuCYZLtGyCIFJZ
sBXRulMMbHySURp8RCMd70YjDO4a/pVa7f2nK/HHSWFwhPXVuJpgCRRrd/km71gR
YhZ6j7M+JnN/HewEmXs+hgoamciLDtJAQtABWJCaV5eEUKmA6+SlVJI0/GGFXUD2
wI85DnMKavSkDGDegpB3T0rCogMN+Hcyfdtg9AIEjThVNVG55qvhVj6Ef7PQsRkG
n6BJudOZYOjD2XFr4Es2sB7ltynDUiD9JU74GTMI6RG0cxu5QSfLC40N+Zj1uyYW
3K7/QtUHr8Rxm4d51VBDOGfIl05TfKPSh0P3l1jfewsJefAAAaJibcOCX8PmoZH2
EKuWQKEPyV8VZRh1cHTFcQ+bKUQJzd0Tqp/d6m2KlpaWzU644Ey8V0wBaUXvc4e5
QWf+re396JWF28jXjjMo2p9M2Vomr9HwqQCszSyGalmqSmXDK2zSNk1JhsY11hTw
vZfYYtIs7qe+ptylMlKS4GrXs265EOBN/B07qoZNtDluIpB4CJjmXyYKpPGodHaH
FZFLz3kOgZq3QSk1z88d8wG1qPirhy4BD3NMHbBr2UCt3vavoZNK/IlwPzmv6Lru
f+EIVk8r4vqQu5aDEmaWeVXlm437UJpMxzcZHfa6Nns=
`protect END_PROTECTED
