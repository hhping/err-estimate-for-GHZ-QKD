`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iT51deNCjXxZ2VS9yZz4HpEWFaE9lAyJG1SZylKR7cBzVE6Hfq56NLwhgRCO1xwb
yfVwyIJV5F21fuakXYPKxwiEGYv7VPSvoGl3sNKQFFBqKKtha3AdCjwEm8NsjX62
dqrgIdaUVKoWyUtv/+BMtKlJgf6xzN2V9egkrg5OHTBaSVE1FWMKKZtKJRsmW7m6
LMagPZKlWs0TtmJz67UBlkjl++F4WHaRCExxwdm67OqSkUFuaAuKT+zC3AQbil8d
pAwkOtm87i7Q9EZiYz3lbQOGO2dEFHkcBx9VMK6edJ/XnSKd6rEaqaT7sRcNuhuE
yRIecosQTIe8LfUxCM2klFF56gX7QfPxP7LCJt51rVO4+Rf4WkXWDfexfEkFWzmO
l+6atXVCircr2+MQChYnFtZMRa6QJzdMAsRgcOpYoseNWvRecFX9qd+3ICUqUP6I
YFDnS84Y8THzLghFilAQeBJBeuZb/aEEnP0xNzvoHoYIkZ6KTXJcC9vdimHZn2wP
sRid2C95Y62Zz3TlG6Qv/AjOfVKgaLDIRqBQ+3IIp0JiUBeSCYWsHwLrET15D/Zg
+3sbI+BShIUOXNhl42IIxwndofC3c2r/b7vrUlf4qn8DXDWJK+YD2taIu/4lOwv/
wjX1UM7Ct6AacH9oV5wkDLpL3/DZwkDoCZcr96hmkusFgu9+4ExX0y6u88pTpapK
SN0ILe/p6RkrYATBRWhFlT88NGgsASxlDfY5/tNVp79u+Z6qQ/pC1TpXRpZMXgZK
9bBG00sEaNCd/MLORbbhHoecsSr8mVSeh0HhdvPQHWjNDDORIhuACoqbEovI0/oi
4bHqGerPppzts+q6RaCdyVbA3bLNvIhCAs7lXX+bUJirZPyZ5I7Zp+hs81LKlxu2
Wj80YMtTZ7d7gh6BDXoQ2Wjn4yCfgZI9707ruxOG89NfrZAh1FfJ8sEtMQs9VyoU
UmpNEc9QvOfhQvIoN5iZFJXTzfbRsLIQGSS599eDsws1CmN60GAyNr4GySMmgagN
IgmnSek9EWwgOe8I4qKvdI84mHY/rz+QETbimUWNo1B4I6mQeUDdHbolsr2FE0Kf
k9EPturdkUm3nZqytDE4mjV/JLMRRchGUxsAvlDzwyzIgeqSX7sFxNlP6KB9I1Ew
zsKJHcomRgQUPQLO4BOYvcPuY+lOXYHuOz1qxJawdue4WkCzN66qMbhmNCSyJxvc
dUxGWpDThdChyzLYNpLoDOJYtN9aESvweN5ccaeiglSJlIn9IYUg30vFGbs4A5HO
aY2B/flkfJvATk9v08lsl2gvHOtDgktxA9UIjfYbZYpPJtl650yH0hoNIOt2mn9W
fLGD6h5+7967MNknf/ZgUr9V2uxTIHJfrNF/OGV+J87nMOG4+ovd+ArNmC0qQFmW
iDp3QCJ0Nimhy5UIEroKtryP+zbbfpsqbpy2QKBb87bLAXNcDdYHMIkp6KxwRx4m
TRK9ZrwwOwzq173sWYT6dY6GWWWj+TvDtJ3QlYnbWcJr3QzGKaAbBVP3RqvbqBi9
5yWUe5oxpxF6D12sDR65Bwf9gpV/dTHGtL+xcRFE4BRsnIpFOrVvlYNb1sz41TaK
SHr3VI+wIXw82veYFPywqW1W0KcMnXJZ+G5B8EnOXDSb99BFDx+la6YW8erUFsh1
Px9ZLhtzQW3Qisx3TolUd1291K4oHOEkUbLMBNpeYOypK8bchDdsjOMUDsjQY0fI
r9Ows5tlR84R2kGr+ZfWBKreb5XHHqbE20mDtmrK9gdelJkkTLSyAazyCIApY4uN
fhzTR7ZWouX5ptndTzowpNBtYDfebmN1G9WDx3hpYqhIzguRKF4kVuQDWVexHQYy
ZvQA6dDUGigILcpyjjb5iHAB9Sw1Bi583RZbpURTCZvmfKkk7RyunmNmj0VoJE2l
YLH/+BfUsGdDid5oozZQ1pvNQO+iDShgzuJLe/NeCNFMHaKUEKx0U8nBr7HYqH+U
+91buZE1WIylEFq1Hdm6o0gaxJIzf2L7KOr/XWSvsgQEgItXGWhIp16jz8o0dNgd
PzxJRih4EvaFJYPNbpVMZ0ls0QT3BvMl8NhkIGPAeayA4XrDOUgOD/9MHBm0JMou
1TGt5vDzovccBclxmPBUL9T6b7CpGCTziJfdMm2SsjM18U+xPxATToVXmStf3dHM
38mADtVjB2DUJCFp1bsyWqfYBaTo3drb/kV7JRsGgQodjinh2prI3nMPbHhditTv
qivEeF9b8cYkKOErKWncM8CvwAyZBfw9xZdSP92WnZKMGRsiYz/PwIDSm1rDCTNC
CuYU0+EJcN17uydJ1d7b6/QTuz3cSpGySqI7hJbxLcgBSYTkZ/4GJTtU/tm/VCL6
S74jMnSyM2tPHl0T/VTJ1SKTez5I9roQxJE42TlfD3NVnp5vfYG9DX20JPO+Kivp
NNbLK21JeF2fLWDzwGM5hz1Yeh+hqPYFqt/gkXtw8fE4SeVlrCTd6535mGBHpmIR
J2KXnmcrG9Vyg1BW/lAYHBaDiLKLzX/Pidow14/zeVIPikWlCMNlU+6owRgr42Ff
b6Xt1kNaB7ntBKOt9w+Fr7sOwIS+rIKz0A9jKuoFV28DKqoqdn191noh28XdrTeH
GwRi+ziEYY0fi9fBuhrPAEKXrKvFvfZsnpr0y8mtmglJd2B4VaONlcP9TKY80Sqt
s1/pXWZIUmIiztljwDGmsgTroXIf1fGcVAEVfLqOMtIW62n5SyeJGPM0rQSyQums
EIPj08K5dBdXb3bto3ggwG0HY0XQ42nwcTqiNriWX5W08MNDO9gUiRXUj+ThUpuE
u1U7zSr+lJkBFXkiKwD35U4tDXQORyVAT3SoFYoFMoDvyRYqQg8fClX4FETD9hit
s1I8MpLgTsBCniy3tD1wM3rZONKSWE3jIWxRtvN3DH9N3ICkwLV+KnC18GeUUnMb
jHg5iVFFuIZDs8EvB2O2D4dYqNKUGP7CeCjfQg0TXO4fjVFz5t/6g7zdf7xpBC3s
NHuSxcK2qurOsrdmBqhObunM/BVdT+uu/4navl4ciAziKN/1MEK40EvtN5lCXGdD
KCP8IGKOgGsMXpnIYxGUxXNejv7qrwy7Q5zwh30dV21RJUxVZZvmo5vf+nrPQFts
QnqrEbMi9px4Ns0Cri5LCP2PP1dxlLziM8y7fXlizd+9fZNvxwf+b11FWZ+OuROp
oTIMs8Cp/GMHOuqnfR4v+ntFGellQlOqBibcBqjsCora8XNBuNWE/Ttj9+mD+iMO
tQuEaSziOa0r9011FeJVWzxqqjOdi1/K1nl7Lbs0f6mGXwr2esXCOvH62F8a3ZoF
VjCpX6s2lL+3sgC6CAqhScSxMhjrV+qM9nue7couoJPq8PCzjFgEeo58ajqcd7Ss
7v/IUkR0ChcnTwAIbhR8Y6MpFAifuxeqLUOTD5zzSx1Q33a9Mn0Goro9q3m+rDPl
EBVVyXOV0e0jhLG/LfmVz2yduBBbJreRKwynf+zAifVmIvg3ZXy7gyZzw3V4hpJi
/Ymnqd1vK0AK5FDSQQHA84t1sdnYj6HrrjCd+nnp5A6oPBay4KYTWMQBbK7+d1CT
B+Mhxrqajr1qet805cUMEVNQHorpfCbaw3y0Dgd/S6jw9xEb1lYeVLoqzzd70gIb
rZxzf5fikAqqSJkaG2gPdSjH6SVsCORe0YUbrLt45yJ2QmbE+BNK0X8vikf1YoTh
c78/GEl26jE92uwkTjSd1P4PyoArewflbkbFYpfuOlU=
`protect END_PROTECTED
