`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oqaqa/vaCpIA5JaVG31Pu9VevBUorJXNp075XE/jid55xmo4rhCGht8dsUfU1Km8
+Zob/VqRJNCqh1JhCazwrXs0lQtjBdS01ynCYQU4rclQRCRWvV5dENCKsFoPgIfs
+UrRwMT4Aioj68F0i6LQvpJBTTuj2yySCVkBFp45ta05Cq6zuc/vACmN7gTQYo0s
j9AvQgCkbvwf8hjFHljSBmZX/jXidNYWnBYdUDLvOORM5zjix44X5lD7wiQt22KD
GHc8sWkN09JGmyYKHOvL/m+hMd0o8HZVWG60ivAfQ/XTp5YHtaqiIbSAMXT58+rD
ss4zExPHpkpcwIboyEo8x7isl8a5ffEIsq4hDSCr3KMpNgjvSrpi39o7x1v3VXrd
TvCDi5KxEOqT/5ZBvjmFp1aPHmiKcd0HQgx3MAD6k2F1a+cpsbtNkm1sIfon47PU
Z3atXXRZPYNuCKicyUJlPKi0E0A3Jzhy7eDwIu36kKdVgkmSqSj2rka1w/2OvEe6
cu2v82Wulpe4+X8rXVIdv/VRyN+l4D081OvEbI/UtrA1ivU+sO38Bal3lnHsLzZd
BH3ISUOZne/dHTREvWo7qQ0Dqe6/EvE17BBSh16FrrSKhsX9L+mzABAeXJZP30AF
Ix1ghZ62mf3PU45NeulxTRvphECFKRnD1dCR4Ge/9+Jkr0eWqpEEYdz56c36oEsR
gHFh8qNgBYDtiAlbOSyO+urudsZ2ePq4sW51Bs5IPlwzv1tfzxFL7n1t16zg1xbE
TPU+PfJSJtf6zGwFnmqeMBH0EKRaDz6aypWfcWU8OKIwd1PCPrTJxQtAjyr/ObOd
sGTFrpF/PLIGmcioy1WsrtOh/NY/nxjW8FbOOXorAo018bvmsrUGMMrlUkf+9XGv
19dmkMG/Gc7ID/JteIaNlRF7kqyr0YlWIupU5WEThDqbq7UG5b9cm1HITtvktXq4
Aiw7N2/Ol7OgsyS8jafvi6O49jheBABg1Dhv+dT5vOPlAOF97evoo7Wn0UzWohcz
2nObRBMCgPZDJBZrymZzZqUe4kXH/KC0rohpT22fO3i52RW41auUPLtz+X0L3YeV
/noKfqBY1BEiaVmp1KtTHyRohY5GntKHAOcceAkWndxW+roiPp0gw0SNiGvkEGXU
3kfL4J/IGRM/O1fy63W/cdqUZqPSEl+M21g0eRIrt5QAO+GCcADpdljyrmgPy0G3
o6N0C9YBX/RjKkiX8AqYNR5Z7UO0939Oh8CgL+vZ/65YQKtfhj2dz7Ucgn/umNBD
eouJRUy0jltONdIfmGLn92fpCqZ8frGl9GcNoDcQd7+8wxrTCMHuC3kBrmQ7Xjg8
UdQxbnwPQ2OnrDf1fmqbSpKE6il3MpcNzTJCuR70vqourjztfNONh5UYNdUW8HeB
92Q0S8IMohO2JotIJo6JCHA4hs9B4uL7isMVtBcqFKu5JNWd64rAp9l6SQB477B9
IkiyrhaAwLy5CpZ5IUM6d/Q0mj48VdB+xVTZ3dv2foaK5lqRdGCNQt+DpBKq7PKv
jXsBPnWYjGC/pPrUSlND5VpVDphZebvLPs0kPjijnVup9bcv3GwXU8oreVrbm89i
NNaoioDpkN5m0jBR3N+rd6qGsfAQuKdpLU7jyrmy7eyTjoDz+gk/E5DyIyfLZM/I
knOnttcOTistrtbskBl/sRqJuoo0+GccExsvRGqvxUJ11gjx8LcEew/BKrkGtAg2
t+ud3KBEiZnfY/OQruS8gY6eTZbVc7BDq8907OmLcLxZdEc/vTZTuMAyDJxs1eHj
iop9C9iSmUjY5qyJAT3xE/CM4tp7pL/MrOuQXwmkZako4nhS0b5WgTEouUR7dULb
4ecQ+1HuJ2moLa7X767FjtiPA7FPIFXMPlkylG231GLeDPcX/kop+Wyp+zbfyIRo
VbmYkvkyDoUjcy08mZT38odP+vzl4YXOHq/iDW1xMLfRjvj2OCSUwIPKoTMH7NBr
ptWBB7pqI3q+dsqGDsGFWL80UIef0/np2H9lbnAiGXspf1rY3fpG7QArpv05y0zd
73Xb8vIb2xmvUDRJsriwXA==
`protect END_PROTECTED
