`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kJPUAuqBbd26sg0ot875cEhxglVHjd2RRXQqiu9INKLmlKdL3t+VGN9WaMX3uJLT
5z9+z4Z1mLwGdB+tMXgjFFRM4C0RtPnpFs3zqA1R23BLXhWx3OSZEyS/hGlD4bsm
63jmd+uW9oLqmZLmMseutL9QWlDjfm8VTbOco2JDSxwaIO2Ingv43NOcmqMYEsKm
TziW7TrjMvVbGmxoEQZBNUMmpmWHtm0nioTfUhibyHwTInLj9n+SR3G0KXDgoeYn
Tm6qGzP30SebZ9t2DtZDn30selN3GBXJltBcc8Pw8CBnvHOuH8V+ZWFBNyvrW1Iw
H2FizPneOEh7LbJgi39ct9uuWaUcfgRRxC9OkNGmHoDNE8pYc7rR3gu9cDo8L+wR
Su+ulGet2L7XFByWZ2aqcMOE1/o1QHosdI00AV7NaxqYmfyoTs76qAUqNaezTGFX
rA+WzWF79NRAIdbiv39woIC7C+7XKD4PwDKY4Ek8L8+FOBWQVKdji0SzdjuZevZX
BvOHfbSYB75HNlOyi4+9T9xODf7eYekoApCaoXxpPOa44OABKjDMdl2HQNjn1sZk
l8Gltxd4C8eslml4X4J/TazII0Of+vh5R3wQfS7uINu52PeelBQIibao4S6RB6v8
Bfc2oNHEY+Z2WEu/tRzZbioHOTXnYQponSPnUlsWKIdGbCTvDS27Bq9bxjhnTf6S
NIVTcGBhNkk9HaYxm+vIKoU2A8Z9vLwPRC9j+OAmWs/Y0oNQAjIkgjo+R1nTjV0J
C1RxZgblZPhxVRKNQvy7XijnP1qg6/4JprrjXW0UEfHlvUISabw1ELvyXb9CqOOi
5bP97QpETqPS9Y1HT1NlwPghL6RinenlTg8Izx9Wc7B+pgLV8ZUZ7mEkv2M6EV4s
8Xy0sYot4HOP82hSDtrCTkYtW94mpXbe9AAgzFUE//5mBKOYX8vElesEV4lb2PGN
XOYufIxu6XWRqpaBnq1aVJBD3IFGcpPziexx0ty0dUZOjLwAfRdLw9NeTwJx0Mnw
294P7+Pvf3GIWbChJQi9zcBc7a36ettMKseCSKQiguc=
`protect END_PROTECTED
