`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Jvmvw3otAeFG3E+x+aNUsTXA32LNsi09vXggPR28OazJA7bsIrQv2UzXveBhODv
ld0mDk+oScQAqyGlYtlA9x21Z8IB3nRf0F3qKbwTJg8nmrCqGM8lg3/A8cTJnMVb
/1RADtnswhQVucvjLAGEN72O7jtgOZ3A3dHEP6M47Ue/V57ow6XPWyEMqa2qcV08
WJkxjxoeaXmCPg7u06H9qnyMYBN1ryxmS29HZWyB5sQPdfCKO4/gHbu03OgqTQt0
zekObgjbIbyK8PCB/sX0roSWgdQsYPfQyCYB/VI+M/Tv8wh4zTiu58byACTJO4Ky
WRaCwdxIMIeaMK5HYS18oFJo7kiL4a/z9AdcafYrWt6ysCBb0BNWjMEQE8aEnI4j
CTZ0k80agjGIAVvOzIw4nBAf63G/3VUZqdBzkJcR3ooQkm8q1B/kWbSG0Kkzqr7X
q9OMr++vap1WXJ+ypFEGaWRuoZZxHBzEAY73epLw3crQlyj598SGydBHEIqY4/pq
aww6SLVvvCoP64/AUWyOTDOo6PmYBFgR2VkFzZd26rNXufuE3JqzBkEke/9/oCnj
vNXmvixWFG0WDUSPpsUqwpdmyKFLbgxi+NQgN+1WTeB7nPcmdGYPrzV9432yb10E
61SqkpneW914aAlwRMb6Lj6f14H7QWk/ucYI/4K7E9wamP9onD91Oc1ZNoIjgSM2
`protect END_PROTECTED
