`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KoQ6m9ac96ojvym3QKEbNBcXr+byW1ErdbdnPsT3L0IKFc3p/DIPOOtQTGxyjMv2
L2HJoUnE8M0PBaLfXbPt5QpuSmDK6UFgmYMGDJmRKkFsobWrDqdEozyhLtfcqaKk
Kr2LHXMpjV4ac1boL4aK/Iop98kLfVM3OnZTaTE++GpbGAwAR0jwIZJslV05C04e
hC33mKE/zbtc+naS0PRqukpC8qWJLwuBeG2kRD7qdZfpdd96FdAQFe/BHvK01o7s
oElh3XHyOVujpyz8AQYdzyzU4gBFKN8Z1bbqVW5T1WDzopk7eEg3TbUaWS3ZmjSj
xBUuH9qXY9IHrvIUiqIEDphxS4tYqhwuea4CIV/WrZ4r//ON/2PrWf6LedfACasV
hQEmv81F4DEG+OqXGUY16MmnJ7SM4Ho9r9qssU/GiaZbBDBj5o1MJlVWC8aTpk4h
Q2xPQgf7KJps3Qvn23CUUxDpDskoo/j0v4IMWwfEaExdADAanW4gmO4QSeSBIvO+
mDi7zHwz4d0iOs2+0FYC5hUtr21EMLgUOhhk2cDakX+hT++Vpoc6Sd9ue7dPZVru
0UzSEb5cuyygAO39N8cIhRDF5hEx3GGzn3WYWs67wg1tcpmeZgYmhCfWH2Bxxq6R
WO8JRtIgBESzn7EFBREb1JMkQsb56stWPUzKxkd5rage5+12gwZ4uojKp3TdU8ya
ZloaRr85y1oMv9/jMKjsWh54Xdgu9Mj/g+hBGMJVoYuusH0T0mxIEivcqfJcge12
Et/yg3k237tC6kX+m6SlFZaAbDBQU1rnQdcLxU1eMDeI4lL96M8Pg3vT9+S592I2
XpklxsmGQu/WsLt0m7IqLBa+GHANwZ/9E7U5lVbbET+mkdbl9Z8wKHVwgUjonPxl
n60//b5HoohvGt9J0E5HuIJLXv0fODOYuP4OXPFm5F9rSt9pocy7JYBSTmck54tI
SDU6oNBgXqmLv1EemDz6wMuiUELYyLikGamd9TcHnFrCKQDrItg/0jK6dlP3WhJ6
RbzwRBRx7wmsIK2s+XMLJqlApNhCfvtDRjjotwAZTSX2yXRiSCV1Q/tWUeS+rimR
qWapoDgchpO7kQuHWx75yIL7+gI+J+Crz7Zf0fB6cSmJ8nYNd2iZb2LqsRVEe0KP
kpoSpZVQn1IFfC8bsDII0ybc+pdUaZgjVNYdVxpKHKaIPbRTXEPD8AQEsEwLtlcz
XcSLsKMvoq3EbCB2G1+6aQlBdiXfb5OQSJjvK8SjPV17swk83DSAg08UQvr4mKzV
/6SDo2cpDB4E8lRTNRmevmsWHrkU36aNCwVx4+F5PkFXHbnnWClN9QdZPLybyjkh
pwNf8ZfNsXDB/8CbEaMd9Zmy4pZXopHoSwXomY9Vy9T0umQjai00+1ufNWkSa+/y
m7wgdwQlrY6qxm5bWQOEskfQb743Kf2Z292ficaWM7E3bIZXneozm1w4VZbCRMSf
EzdJxp4wxQWAx2Qjp212Kx1xjJSu9XSt3FV0++IoUSHD5KkhWTL752sL4rR/UONU
JyJ109Kiv7x0+13XKlL+KIPoX6hob9TLoU3IBZcPaE1wbXNr1Ov9veJZWqzCD00a
ZP/b47cTaXafMirHus/f/U5qddRpT/7XTdRzHeR7ZHXO0i87FRRPLCn3fFgPwCR1
/XRXIiGaT5uz2T3oWF2F90MAvrxj7ru+RQdZuqfvSGXAgD8ISmPihcFrF24BFGCt
H/Ixmrb6h5XwimxEyYekhDuhgnWsMGm/O53i+29hdSKVtxHfI+I2Yg5x5DfI/EcU
1tDyRLjp7HFWzB60UNEoPHFnRUYZcZeKsdyUGARF9frGqBV1zAEL1ztkxorAxGya
JQF4qMGiSMYPwrfQan1runt4MF6bE5LNbYeoTNXEurP2rTtLn4Fnztn39c8Y8Rrf
A6VlyHWD9p+7jcTNuN8uQbFu9H69qnh0lMEtcq9abFWrqUkHQnW+rug8/mOUmqwC
3M4MFcZbGfPjQjcN4TOrQk7Wrsf4kCUqPmuv4mfYXqIj7h4ytSV0qZprnGboRsCO
ANBuk2h5tVDh194sYaUzHEjjE/abtasIPunziTmzh+VVNRhKsaz6dT5hZB941nkN
Q5Ic2waVd0myKU4tlQPCdkoOhd2Tk5A9pMbGeZZ7ertTBFsbLHWYlNCJsj/ZN92W
IDnsCvdzjN/hix8eVis9dGEp8/h+cEayeHeXx+vAPxch+lv1vtUOTIZll1bT6ihP
PrlzIiKprEwhRMqfE3mmDGC+R8tlcFAaGn5EZwuuj+35Hz2qR3rzeLk7iGGA6Avi
u+KES4u5jwqhwN6Qw20DlZxpEG3DlxJy6G6jR/uWZOVATn2NufhQN22wM2UOft6t
KemQFA2f4OVJ3KKzHYYLOx8BzNrVs/mtnozMKWuvl1QMWLJBcaUM6eSmIlSpzbUO
HkQZbJ7hYWqgcj3RRJV1BKxrYmcE9Rgpb7qfH0kod4wHsUeDBDVm/BYPxUamP60C
V11IpRryLvHKytsemNePjYYVrCPPumBsIvJqgi+jEp2j5X/YUbqrwSzU/5EmRRKM
E/lGtoNS39rGzs8CuvPahpFlV89kL3nFuKUbS0VE4sgkScjpl4bGbSpoDdddKKOo
8aN8jG7aC8q+Ty/leOyxapwx/aLrrmMAJdkLIpAT2qWKFBEgGAQ9GJt9Y8M3/kPp
v1z5GXRtO9gHzqt88J+75O3ADExJl/HVl4GB2uRI1HLWmNgoQSn5z5vlneFstuhv
NQFbnq+OFk+1mHPypVqMOofTolpTztJS3RGMQGKTQ1qmvIdeZGAue5sQhWzuLtbP
0hAt2KRboNMZUgsbBq49ZS0fdA9cRCKpihmKIwoHLlvhepoM86ourJ83eQOUZgAg
6AMiJv15B7voa9OR8GbIq+fTev9JJeZLSq+lGS2XLIeE+YdfoPYFz5Y75pUCvMJl
XXYGDMivyUSaxl8C/PaY04d2qBEKUavOWiRHBdtaClLFO0cT6XWpQJDJ/jSq/OJ2
4HkMFb2tY+gR6z45unjwbnArv+Cgw9qHQMSvI0vsG9MjEjDxOrpCocDMDwFMSyev
RE6rYW4QbUjTGbINwEOqrmeux6xmYLhLC19as1g0I0deEd7i9GiZeKcgRxNXh8FY
p1Yw0xS5WjPVsbtA0wqbdmLykFXHCiT1XebIRjlPGdq1SX9NvYb5ezFpukEnuYLk
LTXsjIIjpDKhafXnyvcXYBAb0TQogGeAE7PsjfP8/qqqI3JQ3dgqGE+nZ1BcLTMi
tWJrN5QMLBcnc9D9mDWVmH99UYb41g+1+nDkjJ8l5bJ4fdtTo52FRTYSk60rYWpG
nrV/5nVZXDfYt8lSGy/fuE1gJ3lyGyR/O8woUsl3qjvfIeUjAt9STtTIdhEp1oUm
rjFQ+VSCnC6iBxxq7XQyLKS9op6srcG3INPs4hw5fvgKnMsMaCPVMbDP4I6RiTWq
FsG+1mueTcRaribAW+6QcRbdeLUcuQ1wVr5gpNPpGx5kxpzy/SoOzh6j7cAw2xJt
POxC2+lsQdyJAozkXFiPa1E3c3o9X8LDS+LXSBbo4MX7XPoilZpGOiRuFin0fzJl
S7+0rBjJfqpX8NV5PW232gUsCgfYXK3/zoGLvZTmLrBK2UBHYsOGd2k9LBRqmCrE
OzGWcOVs8kUWWbey+lv9mEkoGpzgWCstyGRgdez5xpMu7lAl5GpNlychgItRS3Ih
6/0RvC7Co8C2jquMuZHRC8tLNn4pANDTI+dAIDNakn50IX9T39PCqh9RkRqL55KU
ud1nJGtXBbJyoy8fwsuDMw6fHPoW1tw3Jm/GtEGTygc1x33BtMVdV73ZVfzkg9RY
i+vjeZADln5HjXNRyAM+zlm+qoGiMnnwLnl42nnzR996jgTs/KzM0XlPFi8Tj1KD
PWTPAJ5W9jw5GzaGBaEBN6t6T3u5EU6bGxAtPsb2M4BR6WOenkRYg0KXNbAX0V4r
s7Hzh7ORlIwgMOrO4uzZJrIRy7TdqFvVd7iBmnRGN5M05OSVEXYX8u1jIskKzck/
X/HVhOaf7gp0fik13Q7ia/xacAKPsc7/wo8qBMGCwXqaryXjm5UEDIZMjflJGIi4
DnW4Rfr1jnYxH1zNjDFhvZ2rejQgicEh8DbnqHSbxXSYMaoBJm5ClyG1Zpn6zpj5
bMa+D6ZbxSTzfakA3FqZy+anYVSE3rZbtrZtPgvB/Y0fggTEXD2tx6cPi8pf72Mh
d8WaMrNIkMsNeOIION8SEtY0n1Llgn5+coSXqhtNVg5B2navg4stFyC+vvqWJZ8A
wHBHkTpbpTURo7moLERJamUSiBH9r9xOWRRwZSqgwSQCS2U4GBUjEI5caX5zY2EH
l/RTJpJBmiWHvJrPKlvs3OX+jLfh6xt6r695PCA4WRyecF7Eq5eIoxOmV4ogIrcY
WFUWukOhHqD96ta4AyHSCK0L7QnOE5S/rPQEDCk6o7FeygMD8IW5xHKPEfHTFPsw
6yaJp0zkFEJzYw3vVmWTSGdaT1VsFxZWM4vt4xX9vd1B992DoarwpzEVQ+GUdIo0
mAYtCw8QmoVE6X1o6VhVqPMm6cJm3KCsCAWPAM1AZ2Cmw+gL68nI2J85UZTWB1Bz
h3wP613MkHH0PM1ankwd7DGeZX9a8MGwYcV7ahgJeYOouR+ivtUMyc1KIjmYqh0G
KxSGmDln2cllY7brEb3+JvSGNK+wpXTOfyeSPh0mNKSDU0FyYXI9Oj9velY/cQ1J
OVEb+ZIcqkRhJj3W8H94HLFuQ0HKzIZvduafsOO+hdSFxQfV1f7eteJKANPs2kbD
KqGRbqRjbUXS03hciUNjifa1GskJvhcVLFnS0lp7EP5sBrHnKJKgz3YGY6MIYOAp
WyHHH/QbPmmYRi2KTN6f/0PdlyeNos+hTbj+Ko22460W8gIlXZ8w5gp/uI8OY43a
l2n33e4gpnStg6JP5YxbkgUVHukOrtf2Y26I3q3qycZBTv9YvIj/yxUd5MWUFguT
QLcuP7+qbXqtnAbr4pyyZGWu1hbocANHMTcrNE2C1R1F2TZWvW+CWWbAzEBdCM4+
h4EqQJ8MAkn7DmLoK4kNnVc9R2zStPI1ObHjexHuX01naN7ojIYoiF+6vFWwE4pY
hFVd+4bK8eRZ1KdGO03EFcdEHM4rSuKDLd/8ekaMwkJc6VLb3ZGUrwAWayhAWvWO
NLwWL6/e+bBe6lZhswckyWJ7Ak2KZ++dSHBTsO8KArqTuLB32fTQmZJrKD+dYmOQ
CJPjPqTAKGZHssRcM+HEmBQ9JqfdvFrLwsz/edwFNQSo33p4S43dUaCabgHspe4U
pOmfEF+cfq+cOE22g+/sK6HfkgndXh5LXhkZYk5oZP7MTRHtfsShFuP5tzUTKf6j
90b5MX5BvuIafZqCc1naCt4IRfZqQULhFFHNPK3HRvrZ+4BTaX0ckPBgspPaCdOB
E46AuI95s++CLJXO8uNZICgWEbQmt9wd9fRT7cu7nGKsumCxMgG3r6QdJTL8SnE5
p5yFTCfrIkY6OTwJ7MOPTiXb/lorFdUwdwKlsVaoaUnFu4B75Te9gySA9/Q8gX5d
UECVY1cKZ6J/SBPPZAMbSKBbIqy8vuRC9T/wgEX7NdsKz3DYsQ6qBp5UlCGYa6QY
6s3ZvAHvJ8nd8OHHj8nBqWtC0u1R4UWcaFIdP0zPJ3RwYj9QCWDPmHVJZ24b3eA8
KWzmUlufOdFbQSgCN2+uPF/3f65gDuovNh8h9ozI3TKZhOwZ4EQhFMl8c9HgAwQh
HNfAOR+EJ1M4k41UAlJBouHn0aCATFbHZSsw7lwY5k2uIb+Zq8E/4eWD+038K2Ug
FGstyPGlCZ1t6/x20oQoySTkxoAn6DyaSG4IRMWZBVIGGOfEeFI4gtfGu6j+7QiG
B7pCUGTdgzUI38/giX1qyuqtg1Mg/sG+6gPCEqdQjW+PF5s7JV4UHUgPAEc+kOQw
Ph5399bJljuUMvgSd8epIFgjIr6IW9izp1D+sIqhM7l2W9ToxE8yZKqbZLxcgqv4
lGlEegd0x1Rc3UDDhKZf+CImZxUNoZKN7U3XKeWKI4aWn5b09/OL6VDkLW/tKtJg
0H9HnMZ66kQVK3jnzfvtl9++uQgKQD6AbxUp+gEKoILEv6RjEyuyJikzFBNCLqI+
XXME8c/hMNljCfDPlKyeP8PcHSq2jEdjtAq5Ign/ITFMqAbscAqE/LLjjmptJTkV
wvphLW99UBH8c+TMe7HRGFK2pVTCujExDtsQTY1wyIKYJx2PRbvvr8YIBFJOsN4+
MB/Cqtpk9s6BltG7Aa6xck5ag+RXNCYy0bliLX0io4LNTkRm5GMvm0fz710bIj2E
rBmM7tb8tNzWJJr9JM+F5S8oCq2MjqtI6d/+c0ezWtt5hPZmFHzULlHpEiaWFNGH
GAzAg0FWPuoSTYOl7SzMw6JC1e8+3VF5FCq59PQxvEwjnKSees6Hm2yxARoTInUL
TP1UrdB8ZCvxzruM70M/fO2k9PCT/rCVO3WNqWfkwVN1nUJCSggktsAPoEIz3KAt
JiJcCwpjhURi8pMfxG80j9mdDe3Sr8cHln+gW2OCsoU+l4l3tUfWnY53E8i4tA0c
bXqAz0NdtYq2GBfRLksy+MTZv+0pwwNV5NTd1cB/OEDvR/YjuS2UIS5O9sWI0Xr+
jsl7bFGQQ0YMMqs0bcctG+Pq/wJpiMuRM6kzrstdrcBU2OvFTujChVX/t8qMVTkT
ELamNzg0TZ3Sup4SD+nLYA==
`protect END_PROTECTED
