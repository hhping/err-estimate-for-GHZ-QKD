`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bmm3vCthS+OXmIRwwYKDzMc0x9qEy7kdRuC7b5UfEAdW6mueX5brB7lfEy5AqKTJ
RfypOC0qb5WyXz6DPPK+bUJvPOS+DXk+an5rsSDu61t93i1vCqZtsDbRE1D+3s+2
Ak0lg0LWjg6OSQr37GBi2j/70TSAbZZgq7X7t44qOdAWqAjOEhDxP58hfvT82aIg
aH3KyHPkxhh2bkoBAgRETzZls45QBrih+m1Sj4R+edHSYk/9GJh0SgHgUt4RdpCS
2c5mj2JPcWwod0fd2NchJnrfRx4un1bV4QHZiDSNQrWN4NpJHeCaZnkOhrjsKhB+
ZRVBeNzTe+2KNppdKL+G90fUtqAEULIHksbNmLrJO5E=
`protect END_PROTECTED
