`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a/Raiz3XKCv+KLhIu6yuhxMp9bU3bq3vxEHkPkCGfwRCK74pMWr7MS3MgD4KQZwd
wSzze3XlvFHzHzRpuTRRkXd52X6nzXhMF63cxCdhwY4JtrXBBSRSRaU64ZPMD7s5
I2diGb8pDowJ7f18+k/8mFkqfFIMzO83pMtaJCZgVp6g2k2yOc9VdU5qrqx/Pe23
oU9NqI1sezRhxG0+qVH7vROBhmtficiZUEhlHD2M1VmynTlKjolPruVqnTuiFjVT
hB6u/P2f/AttKzEMLxPIJofgP5UhQd6oEGjQP9tdig7qkCtB99dH4NEPr+wvFwyM
WtTaPZWou0hUt3fJWDYuLbBkimsKKsoI/ixdmjYOwZaPiQSgbV7slvmZiOKrY9Rf
xDLSBco57Fq6W/RhswdEne0tq1fr2iYKUexOk/TbtwgSSME6UXRLArmrlZSQZPii
3Q63vc6BYwxcL5vEn7OqXNqjTtHVHACrkcQvi1MU/kUhs8m7Bo8otJFs3TFNrCqW
6uEJhhm8a+EoT1f5JUSnB77jiNxjIcwaICmp7jBLWB2VVv3dUUYmQo7vBLtvC5/4
3zzOehdgwJn3o1KhjucPxOOoUPHexbKwHM2/SaTpE3JY4msGhzoulsbUKnFzr5SA
8gMx5LVacl1Oc1vhyUQufZEn3atpIcG30XGZf4UZ0R2PCnpY8dHyV42j+uNkKpzC
REyUZy/mYdKs3ZRX6U2kaRPLnT2rE8h6QkMoYu/bBsw=
`protect END_PROTECTED
