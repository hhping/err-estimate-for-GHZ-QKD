`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yAavNrkvolfTfxs1lXlwdagH0N+qQRo2pxNCgw+VbC5hWhgiY0oBGNjYghsTyMPe
BeIswsBelepNE0656EKZaMl+zKvYBkiA1ZKFi8CmrDJbw+7VPMDDv82u3luTs9Tw
QadVL6PEOK7AfDJZzCNnCnna4spr2sdDlGb0bP2jQcb0AfguHEb7/e16RNuLz1s6
v4K6D4P/IBrjFG+jlbdmLnztFncR03YuR6e85OnBPPSvQNBjuhGNeyW5QVrxNiTi
J3T+xPMiIjhULzRe+Tz8Mcxfmeh2jzLTBx0xac4cADf8gBwVts6ZM+Dp5uCJAewk
LiMrl8zBRXlITylexlM9fg9uSBXYMTbEuTUyZwQAaGesKwOVXwZt7Khjql4jmyUd
FP7hs2KJq+Xw0COWMF8HYI00dVy7b5AjH5bKrlhG4zJbjIRmKZs29ooxMq6J9gki
j+X9K4nnvK3rFrphWc1+3QWIBUrrOplc5urU4hP20k4iQlw79Ni1KXDfBCm/Rzsf
S1/1oqyR1kn4blOH/scWyZ1L9i0RhALsJrij7zZSeH6beJL+q8zS1fpb00YplyBZ
wdu5NbINbDQqBZhi/rN8eKjenJr6q0pXAoXJJP8q8SpgSm+vMX9+9CE2s65Cs48L
KGPbK1qhXf7VjJkN6psBRFVAzgJUuNJaB1ulyG/SLusYryzzs+8TyBlUBTM2m+vu
NAMZ1jBP9M0/UZi3TUI3CDXcQzYVdC+LYpUaG4ZmE2MZ6rFQxll50h4suZt/ZBsH
+Yy9st9lLP9wcU9BEsb1Ry/VnHQOM12NbMtU0nfarCtTFw9whtfBaqI7nbQ1eMv0
MdUKzdtrixeEbNs3ADqbAnLJxa4rQ1XT/hymHMZyT1mT7mB8jN9Fsq9lkbSnYd9O
HgAaVZCAx5bEh9jZ4o9wm/JwfvtTOPQpwKvON4Bjai5ErwC6FSyuG1C2FzFClw1U
SLg3pET2/hOwYSNYbd7eG4wRlK+dk/iWAkyVRDhVAG4ksmVIu0yZaluUAEa/MC1v
ONffL4j3OoJpkorUeEeteHgXuMsyHMkCDGpLjDKcXkJrfl2/7kBatMls2/m6mWp4
0ujPEzFhW+JjkJQTkpKPIpJNvFRip+kUc8rR0Zicy2THqsDM7ut5GO2odOuELukh
`protect END_PROTECTED
