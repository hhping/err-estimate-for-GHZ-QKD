`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vteH7Vgf/ebJyFUqUAd4E2GeT+aY/SPSu0A9q2YDsxG2s4hTHled8flSS89kuwiS
hcOZccayGFEyDc3u2tYNTuykR8z1TW+sFBzao6ftmDkM8lG+eHhsrvOfeIQvpvoX
xJgMIe/XDz3/NN/4N10ZPqikhAjwqhBQhduCzeSk9VdLO8Y30jp/Pz+qFQWn63Di
Ntmdrp4TcBT/2kjvVeu2riCS4x6ZbXWcXr+i5kVLOXIUDocIXRfEEf1LPxvFGk8n
QNzSyVlFVJOz25+PboeCBWrmwI/mEhHZagqjbRzCTjfC1qdTTfqg3TFRyHLgxqdm
VsNvmWOeoEtcDZ1cqugoMrp+sZt7vfeteewz050R7X9nEDe5QYHUAoM4nu7oC/R+
LJW04BAGlvuc70UtzWGpgA==
`protect END_PROTECTED
