`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eizWQlO+tLDvLjBiV9IBb3T6D6DU8dJYei6uqwRR3tyB38fETMhkwoSodPMC+yyR
huEnqughQ63VAxQrybVXRbI2SrVvtsCRR1FeCc3XpXtWQPEZQw67PnLkjODSfahz
xrkUEbIBpjjIyjOF39XHHhI84WAc4ti+U+DFiUFEIGqOdEXS8U3TumBYeW7kMyvr
wuB9z5JW2V7lem4EIx3q9YsgNDBjYjy1ZL5VOqlqY4ZGgsJvJz20Q7wVTxnbvCMl
CXwr5I5CzwiCEjuG+FN80tHQ0yCJeF9KzU3tychZge+7uheh53KBSUq+hvF8PHiM
oWK/G8YeZGMxGjTnEiwxuSa7KzvyUMTww/nZs3ME48bIAk5XCOzFWmgaQYJq/rgL
sEHx8pXyhiA6BLKTRMXy7rtcLSxwzDUqhJvS0JQUyNw2h6KAa1kJHwZlJu/rwbfZ
Uy0w2TToCh3DKMK9WcN1GL8y91yfXX0WI9lj1/Zemj/SznRJWU1Tj2irEkyaka5k
6sUY5UI8EsxKSmZqWLbe6vOYktViZdgW17LGY4Fr5heSVRB//aX4ZcJfdlykYv6p
PmUIjBpp7HQRyyN7TySAdt3YB2eU80olgMlW2cKoB0ZQ0SlAq+Wg4pL3YtMfgJGd
yYmxx94y1ISY0nDTc++cujo0W3192pNDoL/iM0fN/MtypfWUMQrjMwck/aAXUIJ+
rJPKVk33n+lwFe4AUDpHyOn2VMRTjd8Rn3MlUZIo518P0YmuDA+v8cDu6JBrCbcF
t/8gGfrBIsAoGa0rnvSwOMlWtZtUmaUmlk5jsLZtw4NN8p7GNOhFvbLU1ajn2tZQ
uUbbLgGoA/ObUtpucxgDOh30KLfOfygQ/Q14dKoJ4ecMnS8SBoIr0+oAoOjw8qur
8dK+NM0yL3wkWfFWWJPgeI4G+WLoRAPp2XK+cwzRTlK9jbVKK73MUVV3Kh1bjKQ1
hTH0qEgsNbVBA5d0eLvHNl9CxmFLiKFkoPH7QgVrH1a/TG/ks15tmgdjI8n2dGb/
HRXTKKRCf5ryDt7ueCZXNmZtx9poT9b1PCbP2tVR2wbVbgbhTvoFKPhgMJks7Ve4
7tJV+FBtvPtiqXYPWrWCbOHGq0rzAk6sQcnqC1ux6rVJ6WbhSYnNq7Ab+3PxdeRR
jwvN2ru73O1yps/2lFqRoYoqwlglb8U4TYRkIvMS/5pCa8LufMKxu5u6phn8nAnE
lm3ZahANtuZF45IdMdxC8uQk5l2VKT/4UnfyjZ8HAo9ZcoK1iurUpcNH/KKKjc0y
W2skgnjeou2vE9+Femc6VEXbN2/ur8LPBXDUNeSpNVJHYUH0+NA++J730MsGoBp8
MF8wNsFF0zLeTL0GvGwkYQs6hH40zZNJ7iWEuPksCphj+brP/AVTSlFGK0r8VmbA
TiI3P8MymwxGZvRFQLsuAK40idvIOrAy+vzN0IyHgH+vZT4cLpS/8xpZ/31eU2/E
JUlvhexoVnATzehxWP0xJ81R6Ty1FBR5rardovw91Tb974eg8qyuLAc7Je1Q/9Yc
2cdbK9Q7wMdEPCq0AHAy3KGz21vVlAyaDcb3FY2tP7SmXwrJeA0FQVd7/NOcI+FH
t70WqGkZCKEwKBZwSWVR1I2hnRWJ0V/wrQorT+e49p6OpW6+OkYK+2krIeJ35VET
36pCf8UvH6eJ3/69jjklzg78gikNabcoIat2QlzCopMjSDNTlJe+YiZRaVyiiQIX
1FFP5PW2y6U710ofH6Dp78AZmM1NqC85C/bRdA/2Kn8whEJpQJf/A7dCO18Y6CHM
yKAYYOFFRCfSyEU6c1CWSoOOWUJAOKFHe2Nsd5AJPeaNGZt5+zw/HndxnvTaRY1B
+S8luldOm2mT90q9UA/TViorqxVnRQu0eiQvWLZ0gQk5AaVqHm5DtiEpKLU4Q7Jn
HgRz6Pn9DCXwlxDtBucyJEEX66KeeSvB5bC8ky3g+YyECCwRCkIpONO8cLFX695S
tsRW2J/RBpnDrYGJx6ZmkDSLci0YNB9ju/yIzWFWMe+L25qivOvE84YI1GSgyga6
VE4KWRJ5NeSyXNQ+MoSwjzRilE0x1XqOijUKorF55blLAVANmrQTjpfEM2uh7foX
RAg1Aa/uebSjnIv69T6hzkS3sToHnnIOCb2RW4qQyE2jUvgkUkEdo31XtllxQEDx
Os3UKtB7FCuTVzuSpR0Xk4N49bPoqqHQCtaQ7LllX44WfgNf7vLv+fRes3WmUwnC
rFTNn0/NUk3ACZ6qI+3qJxORCgvjS0ZZzEdI7SrTAOqY8BrcCpyRG2m5oFVxF9lk
1yHqkBz8o1OzLcOrZukteTgtR4MZYssFiUIKrdfHWwKboo16nHwU+nv61piF/cre
jaRUXmlsKHJ1aZ9RWxSeyoPIeLtrBo/EgYRE74fHcaW1KL2VJiEkso49j9wM/tJB
7I7fyX9lkj0Xn/Ro94eRmhtRvkOxLL/FwnDIPRptv3O3jlXEqkcH04c7YXOGnAdW
ZPIrcbkH3VuiFC2BLtqyJzu3ZGgXihV+uhXUxxOJ0dE5pAAPnGTJhmPObPCgE/Ct
0LVzGluRBjA6CLW0qzio4vpC1gzNMdVWnpkfnL+OZibqEvFNEfCZwr/+fPtHnHav
BshN99GZDUMNf3xC5GNtRTJYTvG53D3X+FSa31qYpK8+4xmZvXLIBoLvqEl5WqVT
Lvv8RYHsCdV3p28260BHgT5yhNEs/bUBb9pHm+7zPvFckLLSn7WTdKI3Bwt/o6NI
yGBMLKPJ5WBydTjcj8TVG2AL30dpRBwsRZt8RvwhxYZB9aKcLxsdYcd20nBuxDvb
JwZff/7dqfqAtkLitLKEM38GU9L18TmTpDzzbdji3E8h0zfT5kzY4xPHqb4C4exr
l8QCYW+HxtY5GmkH08QvmU8wO0/ug5siCzSPDO9o35EFpkPOuTnXVsqhsRY0GpqX
dHpne3u6sQiysZeXYpbo5CxcHRYpNBgsNuqUn0zVDpTuwZ4/UekmYc+yAWTP5tbf
ftJF1WusUIP8oiSupA/NLImeqrl66XJzU0QnTnw/bo9GMM6BILIomhTVQCJXdo6i
qLnUlzk/uUmYW+TDhys5n2YlXZpqYPClbKScSNqHkrz3HXNhSyc6dkZxyEYJ0FL8
tlrEKE5L5uhSquSC9lRLGBW2vYPJrN+RCbfO1kQEgn9jFUE7XWnGtAxLFOpaqICv
`protect END_PROTECTED
