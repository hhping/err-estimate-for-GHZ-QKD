`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oso1zOyuR1SCOtZkztwofilNxHBmpXBO+Gi+tv9Aab1AeltN3bZSCeUCcf11yUNY
VaajuOjr2ggjPHvKtBVKLeRJU932Jv21cUxCWv0G+nzc3r6vqTr+1COLbg/sZkXA
gQkyWnCtT8wJwxeZUXHfKvQGROj8JVAbRYzrZZLNQfTfbs6pmK0TESBwAwmpZx5m
ikqqHtiRpG9+a+ESsrXay+RObja43n9mJtkdhMl4yqKIqfQC8R+THMVZtGKDNHwK
U82588n6P5CwM30wvvZ2Bf91F2w6bbcrbY5KX5LRPDEruZBpv+guWB0+9hZRp9eI
7xSLw4AYuLzHBpkaBo1LwruyHvjaIyKsSJxv9xGf9PAh3sXuAs+xba9Eg+lZ06NJ
bmcTfNolR1v1aJwvJHXz4Jy1syTMQVfBs2R/kv68GoSsun5CBTd2q/sSfV9lRkMp
GpUZyjAfdBksQDSMoYquxaiaXUIClXDKtb4stowjE/Y4BQ1vI4g2Hbi7Fj4ZAqBS
mtjUHrRT1mJIq7ka77cH3A7kzSnB1wMBMjbcQltcTYWve5uHY/OZzD3px2AeNkpm
WmOTWp7kyo/priLF0GNAs42yEA4j4P58ZITmPbhIfliidvnAOpa6B4EergRFr34w
UGKirxT0oScy9IfmW/+bsA==
`protect END_PROTECTED
