`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3XeeX8m15dfdY7N1tjhH2r29NqPeR/nufI1hsV2txlqhsBcaeaw7TOpvpm1BpzxM
mDn7dA950Q7OUzfPc0r4KfSzQuDwL1AjA68cJXOseGFJOfwXsl9qG07Pw07x3LSG
WXtHbxjUmS7lrAygRrrBzFeM8Ag6VwXreF6hG9SdYvCx/fG/VkxsmifgnY+7r7NY
yS3KO9lmAkmFXq0bnHYsE3C2w2PDtJf1nJyPsiUIJODXLNYeW9KLElAWq+hJkzcZ
DU/Ach5pZQSKCe2pGTbTldk6s1JGWi7ecEXdcexg+YDqcBdFsmOyvRktb7pZRpFo
2Xl9AwHO44caNSdsRpsm6mHw94tjjLcm73uzPEZHiuOgx3AprIcPtJyNyVgTih7+
76KxeJ3513/5PKzrICm+IPC0CKRswbZyUhkcIUhSMdK0JU2abI8kkchjYpOaHpb7
bGzJkBpAk1zlLTSeN2an7SQIcKv+Qpg3/Kuools7XSddwWV54wIXujskR1mxg0iM
6xA8EDgid8uenOHmBCaIWcpuibwBRBn9eur8LT+/U7SOEmpJFQ9ggO+jgI+oPbsU
uSVstyg5cziQZXBK8OmVv1ncVmO8Y9kXWsKGkpYMbUc=
`protect END_PROTECTED
