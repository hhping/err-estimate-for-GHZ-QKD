`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5rc3ipIjv7rCyXZX5ifSrOXSDgFndCqs916gyg/z9Dp7TMcMQAajSRH/FTXR4QL9
S0yRHZDsSUVF5Q4/BYML5p9jk3onY50Xv/t9raJDO/s7SdBzeAvKHYvYTcWXVooJ
LBL+IHNg29BLUXyaBFBWATWKsS+Eyz5Bu3J2Vpx6NhzAOrkD5Kv25PR2wSDZUTTb
2EvS6D8iAfHCJ8lchY+7zvy5L4kSwDHUl7W2T6cVJ80NbE1VPHREW5VgUeV2ncx3
Ct/G7WzvdaW3kmxIQffu1z6bwCMghYKZDspONes+XTYJFH1jNixnoFZKrXiZMgDL
IaWCVH5rcX3ilcOT0U+j2sJlc/fNVKcaBZvWAZZ1i1zRpAwfDPdlOtZRv+bk9w5w
3uB0KWFo93EJUoKvj9efqKQ8cTWg+MYz/kk2iu4sNUaDYTc7gMQ9Ymm/bw6DGEKt
yxGaziSP8dfHPHUARfq0tUwk3h9QurbTB03vLwoJljKsI1Zno+8e5x7o4es6bKTc
VqpFk9w5HScO1PfaTVgVh7epba6z57I/YifGtcvr4zamRt+GmuplXVHPhG15iJRl
d/mAZYwh/i9DQdD3AQ047lwjU7PGGSys6+NjxHfZWiqf92XVwL84NAUVQ5VHksi/
tls6Cg2rxm95qZUIg7XEk1CzYySFeWSIwcP6qO9RAK65SQ+cCKQbGJqopIIi7sS2
c/Z5Jhig0NdjxY9iCooHUlymmVezPJQX2MI2AqclE4WExtXUzbaEu78ORQtzL36n
svwhCmFhs+7O3N+bYd7fZAfEhgxiX1FHIPHc8h9qzkGmm9AmY6my6R/D4vQUEJo9
SPmk2kTgMcibi49Dxxu/Kety69WTbR3mhXWt//lIXSMgnzDeHSgKwrzvaiSHXQ7k
fPrbG1wCKxz6gDxrA7e7Mka+LdabqT0jexlzFsf0oj85U6tFkk1BdgWLPiwYKqH4
GbwXkaT0NwhEZnOms4z6BSDx4tUY31nozbCrLXl0TiCYybrutpeXFdy9gohmN+74
SoRSCruFaThXI7kBwdyYh1DmREA8hqw2r5XSY+OZksf5xZS3t5seUWZMnGdNpZz1
KyRUYx36ZgkRU+GsXBtzFUG8JEc1rPn0OhHQ3xG+bZCWO+UMZwueuT3Tsu3YN7iO
e8bVzh09bPHqeEcIOIl1K3cpNRaGMTFlKsF2m6yddivRcCPVghcW2FLOsNW2uM0j
nYMmWrm5jPoWESDmDzxfIHQ67EtZqWkieMJRox6VQF5uwr4nNBdS/5gpH0X1b5UL
ovX1lldCJFFo6pPNvzLDeyfaz5Ulr8Hq+8eGMvkepshN3IZ+45pE3becrgUstD/5
634Pgob/HVqG0ZUq2TBAYb//QhO+Mv11Vq+DM/cn+QEWa+54sTcL4tr5Xl0DccQ9
uPc36TeHwm/Ij8DXO6xFWa6gAWmLGiwkwI2SoaRXSYcNJf6trZiaEYisuSlI67ZB
iU3YTx7riu5oqpC8bvy72LKPS2qL1CYAvZFK5QDXlnUoL3xUl4syXeXBD5HSXSOH
nptH9by9xIrOJxoQCBMMxFDWACJGN8hGbzlgdiQLGe7+D/D9CLsaacUTM088eMT/
Fa0OJNxxbsX+QN58iUf60S+GDONtJguaczoEDXTqXPtlipsRHRXVyBMf7JxsIiak
/flRtYj1xiYsrDoVSkg6OiK7gtoEbbh1rEhXCUMGigrgiap/Qn7SHHBzDo4u6IA/
nOfjPxVTgTjcxaWBEeSG8fh5hH0nG/2vrwhdhecETgUY76X7U2navb5qBG0SUAmH
PY6X52tYYuHgu/lAss+dNJEKJXzO5gxe04K53z0L7+272Yrmnxz/+Mcpxk++RNOr
ZSk8o4qBGOcR2dBA67Rcfh8RSBBFabwSBoaIeUr67InH0mKfvDh8pT7MdpTBJliZ
HXKoKLbUOyWUfBd3imM1ZxiYbAj2fxA3ru17lO80ZRDd68Mwsh3pxit9ju58RwEm
7RUGTHYX8aT+I4lK3CB0b9wH/MpABDlJYMuVkNKHDudRogvcJgPH990RI/d6AP5i
pBF+Zis+DKx87uSQHJX541Be82GY4jzu4bYI0o693gYQQlMUKv4gEzX64+6n+BKl
jvZowtNFfw37EUtU7JTptNeByk1SrV8lO5omVWM/ok35X83kjs2QDTpo+PF/8U7h
6yfEolDDcDJVQPrRi/OJUlKGm3xICvnhDcJBLV53O0UFAdgkxygQ7UGgAUF5i2Lz
`protect END_PROTECTED
