`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T3QdY7xtH6PYwfjyx3cg0PiOKPKaZoj85BunWKbtJvZ/Mmd1KBKu3YZHKtm1YogD
nxIydD7yVhMi6ZeMEwxGC1JlmWcrlMXoXBJiagd4314QB3id+xRmhFlpcIaDw6LO
SDIJJq5UHZGis1+odNTorUs7dOFanDV9EZD82Gx0e0h4dKn9KvyBPFv92BLlNYor
dA23NRZdkkAeZiG5BiaPv5/3ivxgmrjvv1mC/3ENpU3NOzn/1QNk5MuSX2GP6BDE
URM25jh/8WOdcwxScBLAZKAJ3z6a2oLJzH7TgXQ7orcFXjqgqdTorGcc9wdYnBVE
sO79nzlhGiT5t7bB0ZDOsz92tzaEPAn6au0bLLecBIw18g+95cfLL+fggIR/r9si
GfG0HdbW/769bIuAor3yiKk6ttycWDbQntMyQ1y9mkZKeQQx2ecdlLUdNty61MOF
7IKkqlRd78PTDQ0Uo0aoK3C+SUwYCtDsE4EcZLLw9ZQPsLLJl8ntR0tCrVk8IHlu
er+OBbGEPHLEFDHhtVLa14rWE0s6kfFhABU+/Oi0MwJ8KdvP86bckC/1rlZPiJr2
sQD4v4I62256sqY6KQOi74Obl75KU1e+oswxWt/1VEs3F7oi7xYNzjR+YiqSTEZ5
HyL+6wEuULJTPNJv/B8SszfzGai71vkNzPgSl8VLtD5PbIiU4K/qd4t03t+HeZT3
0bkaOQs3AViK29Mqvp/Vi4sTpkk3r+JHmD4A4KK6oDj0cUGAx1odw7XYR6Y/d1BT
LzjHDG8DVlvktmkkfYeHIrehA8lPuaZ6UXt5frtdybHDBxRkaTUO5JFrwQk8+83E
NAHKzbm8j+q7Y6wRnj1V9BWc6Cju8JtnuMWtr7YaXAb6PrdJiSLPoNeRVY1PU88G
/zy08CcYHVBYIRaK9tMVel6C+sehRtgqJohFqS1r94VG1Pwap1x7jA+Hko2CBbi5
CoVBeYvqfP+e82Q32hTjCztqbMMfC658l1d2M2U7vXTIvJafyHDXicMF7L5DXbla
HhhWV5wATHWaDoIZ6XePjcibLrho1AvuGQY81vZr8Bf0aIIlXiRWZqBvXdsG/uSu
z+mW8IITP/3jkzotuzVeNAuToZ9MZ+3ah+dytd9iBaztZ7ykqykB7rytJXI7aqDd
9PVNvlfCM99ytTFtquvRkkcr4vNBttdheL2fXSrhWYvwJiY0m8CJKgll+1nkSIny
oEgNOcITsVEMNCUpsV3qzAGfKFmU9YPY1UGpy9H1zYPbesa68Vp1XkLWovEofOY5
7euOIpRZKHQY5NeBkdVY9MqpqDrhfpZjcXCQ39HJSDtY518hU/0+RLwG4I62WQtb
aTzzPPFbgg2n9BgTgTNDeSGpv7wj2hHOl++z3BZDumjw7UHTRbs0339XO5Yo860L
N1p3NW6wsrHD+WEJI7xixNvBK45/ZI4iRzv/8mrSMwInmw7xJNOGKPz2YU1oLP00
h53uw4FclpwHJ9DOhAxc7qShP8h3LKPZmsz35Kf0Q39SH1vO18LlUkJ33RtRyt+a
11SrfeY09SYyTeEjOwk66gNtSKUruHDW0loOZh4xgG9J/kxFpte/8izXgEi6SK9z
V3Pjrzrqk6YSpH4nADBbEtCrel9yJdlrhHlZPx/MUaJUDJyH6LyghymiZEZICwIV
wyCqGcN/I6Ens9OYTuACkiqSmJfVkj6OtdSixD1zGuTuKMm5r9Gz30qPNLgC4XdN
czzNUP+vmjYC4fmaPMGCoSA6GeWYzmvR+QCrL+qC8IkbXoMG8cbAztNYd58wa1hL
jajk27BsoUGTJIzxgLVeJTdJQLMD7wOWJ3pVseMANifjfnxRzIw6aChnZJRrtepp
rpx+NaMDeU7iC4EoqPaQ13YaRheOJz8qrzrfwqRctc6rf7N/hveH3I1C2i6F/JhP
BRJVPBiTQlZ0v0hMsOYe7ZZ+UtvmUL5EebUI4Yir6UdL/68ND30Qd65cQukQCpXb
4xGtxdyYZi7iu24eExv6q5T26RdFD5OdVAVbPEsCchgN0thFQZq3G9P5iGNIuMMH
xecDDzCNfO46hTIVyvGOHiMhMjyU1Um1NVrFAcGjK411XqE/oAfQdZyxg9JGt3ow
LPJ2t/WYJekpgdCHb99tbGSBJC2VDbhrYI8WeeU7Lcu1xsE2VxoFwF6o15PcIUmP
x/ud35VZFx+l4W/WMoOkPowlRFNxkA9fIXSprU394JV3Fo2UrmUm+jWmwegO0xuz
aR6w9G39b0rt9tHTDWHhZ6K/y5l2p6Y/fHGihvb9W1kK7+p1UU+kZzJimEF7Dae3
v79FiTIuqgpFxgEpoeyEmObaEChDX/aSFAFcyPSisZJRrZQCCKP8T12XvbGzyTwk
m9VqZpC8eoZAQmMYqRQuN4QXM9m19kN5NTL0uzOGNtsmAmmdT9wpOcBg52E4ba55
XqltbaiiYgTB4buZKnuqyZfMV3N0YSlgFP4Mp5CUJiEsMSSb4gIf3YHW4A05u2gl
Igz8MhmKUUovITRwpE5cYCb738zt2/lv9QbdWCUKoYWt+rJDVwdzQ6pEYJvloTa8
5b/WMqcKijTYupRKApLKy+ODyQmE2s5bZ9O0gxaWyla11tN6QBf4ObUi9ql0J/0Q
wByHjE9kHAHDhAdrlNpVPoCid7tJZ3jqrE0rSChZhKO0hSt9wK3JdmRfCQ+JTr6I
fD1IOajHw2M7JSB9gvmaMWZCQoigeh+qSJ7376zeIgclEGaba1QPpo166m5ZcVpV
FJ6UzYxhSMAQgFTSaSLaEllB4ODWu5E+VnR4mHvW54+yZT9aozm1aOBr6Dpj7TMR
/hnl2yZrcXvbAhf/pqcUWNjkutmuacFskCU4eJEM/MZ0lP2ULMS3nKPH2dPAjgWJ
bYfYfOumBecom3hi9V7Oft4RHqjAZVkJILqsFzFkZ9puefHLyUh4Xyw3VQnkaRit
KOmAhw7oyJxhlHK5YlZSFnRJW3f2/XFs7LWxOtNzBz7H2eN7WC75Gws5Ur9y/dc/
pDEZ0CqnBO88sYfD0U4Nlaf5/Nf7k86PqrPS+7Lz/F/gtStaM90yWZ/wWXLI30ew
zwbYOyyjbJOY0yPkxFAAG11FuHDejR0/S8jQqUSQ6onjyCDVVoE5BQ1joOOgr7kH
MrQdlaU6KntaNgTHlTuJvLAc2NVVCvajG3JeEiDAHkWyU6I1WS/0bzrSNd7mEE5R
DseOlJQbOhVrXhrQrsabQKchVJFJw4gIyo2QG399IrhV85Gn8dGRr6+Vbtv9szq6
g57439itLqbZLfYRbtM7XlOsWkA+zyb6Q6JEfQqWoaPyHNn/7G6g9KHFgqp8hml+
lDs/YZs3vAl5tp+W1qRNGl7mb7sBsplebgROF0g1Z27wfppzXJKSC+khJ1G3jABe
q2MB59g1+E/M4457zxkL8725tU346zTzkmC2VSXyTzuniWxl9UcAgfrHc/tf3dO3
Rc9cXQZDGWwh+eZdmxwEAvQA3HVkjHJcUpO0c+Qp8SgvdSUIQH3h1z0h5f5XrfYO
z17T4R2TMHzAenrzfjhjjkb5MVlsQBlw4ZnlWEid+E+3p0sN7PIWe/vPhHgglstz
BgxxvhYJfy+fwnWcBcgTeds/uZq3T1f++YDl6n8SsuGua8wg4k7hv0GfgHXzv3To
0Esk/fJ5RYudVSaU87PYYITJtkX/Bdmcc90lzo++TiRNeHBhJ2vPT4H7SkfRe6t+
akenku4Wt6mwlrsH/wVxMrc7ishtKAkD/U5LtDyMqjUcMw8EfalrjQzel7tDOAfE
0/Wg+wby0Mnm3ZD61waoqKzHzs7NPDsixn717fK84GZ1a8M1ftLAGwH3IlUED3HO
2TWPt5NNj4fIIgf4BgTRUegqH4Tvr6onTFZ/yccWUlEwIlTPCEJAsww8NoMdRzgq
YF91zd+nK2PTj+NZnWVRhO85xKVSASBnW/9oYW5cFHJioqiITBkrcuQNqUlSOgsZ
gm1XRgcYNHSADzQXmccU2oMEZe5v6o5F/aS0tuJ8RurdL2yIOxNvsK4WbgrwUrET
x7TEd9/TnqfjNWi3+lEAFVzTRSEVjPZ4dzk3i5C74xbK8lc5LQbatCbJAgra5zhP
PEsinVApl+zvAG8r2QnB5d8yMKXXmoxuJvmJ0tm9iJ6oAMUIyKhDeB4aEI4LD4g3
M19tkcmPq916cxA7RbP8npomRjeekMSyeH0rft9cJ5Qi8kKfALyabNInfhNWRPML
YyJw8h/Twys1ceGa01kmjhjyHjU3X8X+DwO7TZ57ZpmtgMRt+Dnmm4YIvjZD2ohf
TV213m2siCuXl1+ap0JaUsctCOGQM50i40LUsPGxU/Cn3lEy0UGt3UX3ju69qY8Z
FQRopVxUWQ3uXTlzYQOBfZJ0c2PO+Szi1z73baM7xUvF842K5OOv0QohoRni5ZM/
gNiprVQxhxadUfKirk3SyshpBG2LZK4pMOC5tuIfSlzfLXHs9c8eJw86XP59BMZO
GqwjPk7bTwLKM5CtxBGVrWFYdEvBfg8jTp4o0Aliy3mGrzZBR9a5ugwxcVb3F3Z6
Yqk2AjIbMvx4bcmc873+69kW8FvstLWCwxhI7cpleF9tLq7DmPTNtbSSNNDJf2Qt
TS137qs3/gzai53Vh8/GYeJo8nK3NVAxcdPH1CHug+oi27b2xUYaP9Q+gCHdfwP0
9yeFm7mRU2RHaU+quTfairsWzDKD7tGs64ijeMC2Ff8P4MUmu4miOYnGu/JtUvG5
JF9odrekHQ6lpB41MqLAhZJmHn9NjZRQk7ngxxxvHyJADNTbteppyfjew5c5Tyck
AJl47Zh5MAFGUkBt+0BDeJF6ER/nXmb4PaCS5rglmCE1YfuD2F6PXoOEhU2P6dmN
1gYc4qvkktdZFHJNYqvP2EJILGc8CJQo8QXUgtUCFefTenW0IcTHUJo7PsptCyT5
QWbxhiU/bOHRTW90/+DkTjydAjsHdBQlAywPLyYme9iOQATA3Jjkskl+aqWoEJF1
n/PnZKhq4+hO5RD7YMkhIpsUcLehia2km3rrIg9/Lz4kCA4EO4WcT8jd4reeAeSf
ZYBaCmigYlJ9yUqa0ZAkYET14dxydIbPzWobluMEXf5XdekGNlviTVX1PCI8Ghcl
N2H5eJPWdBxR5GLvn/oAVmCPg54unQ66BrAY3SDQgFaPIvJAEculcKVz1jGctjZ5
8n/ShngtXvI9xCJM7hZHP93oHfNIJUXyIykXeVS0YCVZzHqLWQe70vUwrJ+d+SUp
qrZvMnGci884wrcadL9D/JymzPnDuCwuXXgge+GnDprppSfe/b116f+zMWH6QwzT
DjDggEZZxkVfksnQEbgqUgYaC9qYJfFFbpvMWNhEzGUJq/AVwjpFEgTA70QpVQkT
cqWE26OlZ84l1oAxpItHDEIpRzGg9SUedmnhLOVTD69ITOiRdJ32PuXMfQ/uObwz
XqyNwP4ZGLp2/fKgIlbxf72GY9onJnnXypTFd3JnQiWfDvN1MYsAXPnAUf9gjatk
RB4f9JeKCnce0f4hkc2L297TquJl1eDgOf+Pxz+f9ryfY9lc7mdQvikrf7wjodv2
GQEYvbsximT/G5coYCBqK2ajZcxiHnDOxPg6Pm4vV5Hz6uCQe6oKxgaA4Hf9ZGiI
7Sw/5imzis86dPLKmgPLJFupwwuIX44vO4Uu09uCfXMXyOCnYtWgUUFNiirtu8Oa
V8IgceVOBFN1uxr79O8F92jXy+nXBpuLGC6X969KqjyHagOFMZUW8i4qd110uG+1
RyyLr71kKXWhfenEwTesl6QybyWpn7FGQBdZ9VE7NjOnrOfOfXWss1EK5oINeITj
IOoJYwMngkW2hwEqR9Ck8hzbmsRb6lWw5o4O/hGTzr99NAjaE2SMuFRNPKkAvzBT
q3FtX02CnMH6NbZBf0PKY+wUUGzyC7Bqg9JGVWOunZVx1uWoKOwTX0BscJKICQkT
fNYtKQoGmS/dmvGypNDS0q3v7BN/+PNGY1Ypt7xzOIS4pSwpAdmWDr/nQHtpQDl2
VXi33EhBDqkL16xoEkHTWK/bEBbq319e6oifnLUAGOEc5QuXzvqmuoGno9XmiX3C
pjgPvshOGn7s89yKdgHrtfpZbcRbFTF3a9+56X8FLUVThlI6JvIJiQG4K2gcWDlA
W5wcNpeBdVle6x8+Hu/CPvbQZE/SwLWrSObnpEF79vY+pvsDuMEUDcFCNlnFnmM2
AFvq06MUEyZ11fNNF+34qHoASmvs9VhQ8Pp81l21ZgxOreml/m/0Fotfcbq91H4h
bIWbCU8Is8iE7jTOF/ng66k/RIKWWg+wPhrZuGYRXRHLLvbwC6hDG/hSwUUDMXPE
6nPHZzDCPdWzh+80zL0NG4gqiP4duPu10xBJP22K9W/+3pbDpaJZaODxyHZGfwtH
nELkJN1587j4qX3i6dUWBD+WbTeSRugmsNl4aubVSENuiuALegbHJY+NKpzStnYW
Ov7QpHSry2ikpPCB/aTM1TQC04Iwcn8cANH+qP+7FNd4tT8skZefdiyrVyAjnTaV
J5GXxYDicS/kezgFG0LHgf52qV0OkuKFXy3Bw6z52uXdUF8aIzu0m6/jUYHeN2IB
zJguYZ6HN0eW8XcuCUTYU0QjxknlbQ+k9iZeuXQLLYyLf8+o1Vzqdlaid/2+bJRH
zmboVUILKWV+fOD3K7c7RiH8dDIGTwIb6tNIo9GzeX4dIQv/thgRDW1SEURJ7sDf
IqaswRspI3XIMPub1l6vZ/a8DvXv5iVZApKsykwO51DPEFfca4XbnNObGXwP5jBu
lrcimI9SBkd7HAJKysQQ9KvXFdsDGgQEZ8p6nHF0w9QPx41TxvRfEzhDCvqsanrh
iR7MqvcO+Fo/K7v5V/Gc0HS1SludK8Ws0fxECjilNOdBV4kb3PgrMgbQ3fOKsB5Z
8QGx5nRo1RWZcm7PuTssKW0z0RD46EDhX/m4l+03ivu9W1MeKRMHeOn4KO4lOpVb
WgFUKwmAiTCZxgJCLYHeeyE5PXzM8uVWTdh6a1JQ8gPFnh68DnRVwAl8waTD8yGd
PN/d04DwsBlrliwenVNRhyMzbaYdj/YBqxblfK6IEr+/xwITaprYG0XPKOmPSTpp
6KSlVPLFoK3lSxVC+vhLvc6Hi40PLi9+QAq8Krds/ukn/LI5eDcpj2p4Rm3pRwCN
NLyn29fyVrMh4j5BMSPxMUAHrHntCn1XnLPVlIDyte22McocnHwJukspiZe2t/G3
VWdgY+puWyGLD0WAQ/kQa9HkgfwfaVghVq6oB74mDrWQ5HrJc1MK+9DUvfh7DUdG
CiVvM6UajUreI/C7Ay/EIhBIHLGBMXOvS/Igi0h4TWBxAKaC7RW7CMwVPARM/F02
m2Q+L/ZjH8enqlOeQgrJpGvVMXCaOu2n/G5B4IRuRYWCJfU1sdL/KA23cnXEqe/N
6BM6oaPNQlAExrP9eG/zmjAlTZfvVa+6lO/lt7/M0sJ6yQeEMQ57uCoVgpVre2u0
s/pHyg5HUkqG/xlgq/VILOE/ZIqKqPAPFcLEgsa5zDohgRs8cY9KEveS9Gz0avEw
ZPWYfyVWUzy6p0kUMKdhqmNjsQrY63A+LNGwOSz0rOjdjxGXDaY0cG2y5fuSdYLI
V7K2YfU8ivqfiqE+E+b9kg8B6HtzzZI9dGumcu+WRF1/bqsvgLKJTSyWR8kyplDI
HySDSVn/pMPYL0igOKhYdBchLacyWeg6Q72+xvl0a+xiye5dXUs1HnKPwdbGl8Yx
0Cnud1QiMgRAZrzg92YScOx+2DVNHp6v+/Xyt44rdc7lOaXcbLVi75Gu6crtb5c6
Pz6oqjgHnYDa9nlDTPDYjZoYtxsy3eHyGrSnqaPcy0LuIjkvTUou7c2+RcsW4eAo
S7Hj1mbOC6uvTJdopR/WERelocnVBK07J4ekcA/EiibU15ANPFh6LZE1Jf1H+37g
rPq52FOgPHDsWgnQVdx852hM6zdUW7r3qoqrbSn5RruvPx5xvLfFDzeAcvsuRIj/
0poy8DWF3S4QOecuXqrgyfA4P3IyfZ2p5tR71//+ltz+K/jJ1aA8tCFhOPLY1WB5
3StBtLbOaoyADSQ0jq3BW1qtwb6hE9CbWSZMb6LtpDTCfVeFMqHvVoLHhJvVlasc
HUVhKhqyjAc/RcfrTPbQ6heiDk5BmLij0qiJ2QUDOS6WfskBsIXDrclF2sc3HFQF
dTarBVlOODFY8hx95lnddvuYmO9Q+u6yO14EkfIZyyoEyLtUaFf16xnm7Zo4gF5i
HuYMpdM60UfvPAvb6jP7RNUJScawoLhyp11afq//ibzfr30E5zOfiuc2z+wn5ucC
g8iAohOQNeVFOilk1sYNwJBP/x5lrwWcAgQI4/20WhPLQXkuX/gXlEfGrnHcur/B
bxxhMQa5yoDH06v1RsBrwXMIR5KZRH+FnM/uWhA2/04ts/20Z/wrwUdiCOtGifT6
hdP6NOdnHTr6TlZ2CVaDTJ0dLXQLR9pgYt+zS1K/YllLEcOp4/SNCP1dhklLvUy2
i+a0mZTLIvdk3kFK4DsdZENcbVe7R05CqwHG5gbg4folkKIMb1geOCyRUJIGpZwD
DRerllfZMzjAzocyGkSUaoQ3HaKW/LfBm/PRmGBAuEf9Ja/taamiD+M6rQipHXnr
ORMFTZb1kfy2Pgt0X5h8PToAKu/LmlWTbVmZJ7Egp9LUNiLuL3Aj2k0IRFtBDoHo
IiKFCToi1Vyfk6B85miu8lnlA281a1BwcnFzVTQ0hmIlbKGoBQ0GVVtzl/0WFTzK
zs7jXAEtfhmjlXZj3Xq3k+RSqb3ApJVrBpAiYSb3ZEcm1d1eG+hOp5hWfToyYffR
XGaiJBF2RzL+5oD972wgyJS6pJr1OO1s/2JvmsusdZVG0brY3A4gQPef68sB8egk
2bOEXjaDoWdNQ26ABdQNSbrqJpSFvoRvIx+nm00+6UFq17Zusuo2D469IX5CpDze
pwPekvuKrkuygLq7j9KuFZzWukj5Ff7SYiNx2FF1bCJAmOxvB4MYDOBLyR7Znt0H
ueCWjwImj26Nx5+ApRauGRNCEUtBKygRIOhciNJYPisSqTizxGgp2RUyxSTjgGkq
kEK8rkNDCMgbDr9ZcSUaohw4MeHz70ptTTJfWlmUYIxtUCRpaEhldRljIlycxlmz
C4DYKxdi5qt+McmG2QhWFP2tj/c5jF7F8lGASji7uGIkFEEkEGrQdUfWy1dnn2VY
uE3iMSvdqFNdoqzl9PDAY4iTz7b2HG68MOG3iN3cd7tnyHH/N87qBMEER6RarCgl
RK/YHe/cbkSGjon2H+NWkBbJ2qz6rQ8euZ3oSEHWsrZ3/mLJ2to+cFa0Hk/FoA0F
ennrvdQSbpFVfBk4dshuRm0RndgTWhvcNbetdoKxZxOok0mhH/LZOTQv7PKSSu1y
Xi6Di0gBKL2URPzks6PXbv3fv3sDvXxZrjKG6fG/DSKbjjqsinahEGzK40ovGDTX
0RcAhTrQk5xvcUCX/tUBfxCZbjgwdqgRkov0KnBrRM0RazmvfiJtomnceqfL228d
Ppw+R4W+RFtRllmHH9c1pDsIyshbRUA9DORDnYvrZW17abUUylYlxcnP1y6iPlpo
Cj/gqUeiVmQidjJyvWh6ubGc+fL41rIu7RgipqeHIUcm7KX5r5ZQOVpq2muqiiN9
FRSe5pTU+DwN9ik+5X7Z12/2EM+Yk0zS+H9p2FaIvyngEPdsxMf5ocfQBKm4YOY1
qh0Vnwt8eXnkh4Sd2bSKSz90CrI9yB744MJ41n89kTqs5E1sRwDilwT0YbkWZZD1
yk3NA8Gs4IppIAC/a5C4k/516h6dLpPmrZ+8JDfnIVvRtkX6PmMwAjMMoxjEsNxO
TPh3Av53inf3b1VHGwX2+x6yMuzRyF4hu0tLFZy0qX98ko9WCg8aEi7JiCp1rz3l
URi1OcfVJnKbo8t4Fkd3NqipcksfZGY0xZ7fY4F3RJnwIKqMp6633eeU0Wtwb8zd
T3/98FH8S8mr+EAzROgAPYNFppuojk/2XCyFD/KKMPWiNn4J1fS3slAQAYJbVIsF
igbAF+ScEhsHVuaDupCgC+OspcAq3bOsKG8Ow5CcfFbXb6086T4p4mOn5kpPwz2F
7KI7nATz4jBru3ahJFLOBcDt560gSdUmqLEKX+etUJdILCXmKRtrA1YkKXhWN1tx
NsXa3EbjlUnHFZhdNJb43SPS2Q2sdOTkxD+zt4nkU1O6aFwP5sj+DdfAFeMHfEHx
g9Il3Fi3NWgiUC8+rvWjm4gmnkdKPH0ytLF5o1dheAwMZxSnXo4uGN20DfHsp0A3
BJU4ZwG/oeb/VnVe9LFUsdwZ4HoIpkvSLn8eNQ3SG/1MgvZgSn+svNUpanM79oId
Q5pIDHRMwlQNSzkK9DmeY4sJPmOZqzHxJF3u7Hp1qNcC8oHsbobIe2grFygVQ3a7
qfnYhMVHp341+0R/AajAhWND6PXSU3oO+j++3AiU/+bNl/ASXPR0+XqdLHZwwHfr
rGMNDk43nICVmoKr9Rd4QCpTNcDM8ht4EuGeyEyjah+kYCgAzpqNkp/MhJ4d/qBk
Jsy9T+ZM++6bBldKuCFSxHVegMZExT+yAykruBqvbBmoCnDIUfpc7z3pBpN1nobR
ZoB35badLNwW7db5IQOYcaTP6pggo7F9EYv0xw+zT98QerYHigwVoYLtuD3VtoQO
0TY/huX3LVWGrKLHEO1PH18kfNsur62t8tpABfTHAe3v2YZRIhYiFDMvnmBn5e6X
IBorWyx+KUKPnfmJjcGu7QbVqTe2OJp8vl0kxMdTOP/dy/7R+2xowI9WkYX7FC/m
dMh8VFI5ZL2O9zVG8Bv15M3/9+C8Uk6fiUP84kDg/FTXLF1bf4QkxUQV/4wEYh2p
QBNXW7GJIlKnQ8pIuO8qRaUtjq/DO64rfUtG/R3+bKwkWPYHaaDhNIVERwIR36MP
rRN0Tlwm+qsqyRbZL7hV5UUbmS5mzoZ3AQT/CJkG8BI=
`protect END_PROTECTED
