`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xqizNwJDQbl3nSB1TpXqwy/5NKrLmPE9aICwu9neB8Ur1o4iI3pCsc2VdFYU1g4z
K7KqVC05eD5+QmrEACmcktNF/FcZQzZaLKN5rkPPZOEn3fkC94EMs82z732t6AAu
KhUs0KkP1tF6Ei9gakgpxfm6ZCUdd/2Ru9qEO3yO1Pc/xPL/gmDuAeb1ruM574V8
9/V+TLW7+RZozaMKmZhM6CW+uMZfQ8rBvyaLwd1msNVU/VrTcWT/WWLvESExInry
NavEZXrlngf2dPGAudl03xrIjvt88d1lJ5QBcYkH17VNALPpVfgNbmnybP4+ed8f
2xDEqXBK4tclbGnieZLfNzmHFbqVowC5x+9gJ65CwMc9SxS3n2E4wjd9EUUPIOhN
OyBC2QMM8pAnoYebcZaPgqjktY/IbIe8UMtEKfWrfX2kDImzx0tm6VgHNoq6DL9m
7tW3xL/vfnULyHQHcKA8gSVAWZyi1ojz+fZQ8VTjMKA=
`protect END_PROTECTED
