`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HC/xLC4fk+H2ajXA4i0Q/07+1dzWyHt+hULaeFLUtjCC9aNMOIUg4jhxGbQBLPRI
SPWICRNpTcoSCGo7lgcKN6Lgfiflmi5L7atvadKO78174Xg/KdCZPyRBvEZxJ19J
0Sae2ltdgArf1tf7LeywI4o+KOo+j/oGsadZH18rfTlK3Wk3D5PlGdbVR7gc581Z
hurPXDSbCvl5dPXzRgDk/rudttNxXsSR3S39zmP++CY/xjfzZni1aJPnB0XhNOBP
hgcY1MLRV99K7U337U4eb2sXuqvZUjz+MTMVLmHpS25pUwg4ZjU40lUWFX7Czpc4
D/6cp+zAEpcvW+9/fkfiFHQwctD7ZuCk9r3cTm2U23oLglHEJiLff0qWbuDqcrR1
t/tNiCPHEZhSU1J8vGMJ7laS8ZEqjoQNJSvPOx9dPJXWNpK9Z2dOFh3sTAZWscwi
+oc/j6qIwsgl4jJBze2V/venjP6kcWpBtMbDAWDvRvMbKYiaJAES75dnQGTFoVKK
YWpd3JBQ8ttuvL0+JIrxnqGpG53Yczw5M1bN3L78IR+sjsuDlE/XLAB95RUkVOp4
ExwRhOry31yAptUGUYGud5WbT13AIDCK8tqV2MiR0mhXrKvBkyC9heW/DoPT9zfb
+xC7X/nBziM39U0X15rVJLpEELxxEaVhZvyI1AsaMd6Ll0NHLYlxTBZgEzFeNl6v
iy4LxzDNwWh9Y8VPkbK+bvCOWl2jJfCNh8ZFuFYZxKgy0fkLKVAEM1aMpSh240N5
D+aosjRnnKmHoaqu/xpohLtQMgxdvvrueBDtaAj15XvnzVlThP0MTy8z8FT40gRh
18sD8FyqWs2LCDcWjTd2rAwUXMZ7lmGQ4SMvQlLyL9rUlcW48r8I37EsSzvx2sl9
i5pv1QkJUIeFA0+fjSA/dqp5p+U51sTMwWKoHk/3LlGmowrfopIj5kxgawkqbOZ6
pB3AUrUUQtJ/LibG4gzG+MOUvhM0gGfBKY770gPJArzcNyeRYar3zTeoj8GI0zuP
v5rQiQqbYHHb6wC8kvj5uk1Ngzv8SbxUFKTVpyywHFK4BNCT2vXlTNYceJRTkPRE
sh9bkr3D4eLWrSJtXoaSgBKOY0+HixQ6P1DBoQeCeN7VNTCyxJxSP65uA/e1A3oT
/cOdFuV546ixd6qC0+Hf/BcfGu3ZjjwGw90tfUanKk6GYDKEcRtkslg2d+HGI102
StizDnRlIgicJ5v/yxyjwhvR/PBorbaN1fjXZkYxftMZYKwk73jHyiiKl88mMAsc
Dq12gIyl5qE5vGY7xtWHNnVS6T1Hf++1nfCq5tIcjmfhNbuf7MnB2akWxGPMri7C
oz8iZrqDJroNWGd3gaOOJjCxfxFZ4eJRHRBIF7MgRfzwyHqk1Yg0KBUvJkAeQTYc
1h7FlfjMelMvVQrmLYQ2NAGIuQJ//2c/xLYmiHFL8/0DYam9EhlHw/mm1J5iUG9v
6ZQ65Lt6OFLo3zenVLUa2rQ+B4FJwB8eu8mJHed7R6CUZKunFJ93g6KdECU5ws/R
tZ7xbuEE0V7wU2+Dp88MEvt+2E2knVZ5Xbv1Xbc9h2+LPR2l5CLRJgn72RX2B6jj
aloYRF2V2Zcixq3/70Jo87IeNQ01Mz+UIM0+QSxDB+3mmplnmgC2e5W8vcszS0fx
1BAqPPZ4+ldREvYYufyQoYHEzNBJMGfWLgOdnLbI3ZcqbUFKb2xbE81pclqbRs9e
zWGymGYOUDQtxitKKjyz7Uxhc3kQc5qClqZwUo2m8mLz8TgzFALbYzVx58s89t6i
KhB9EbWNp4S3uwGoZ+JIDQ==
`protect END_PROTECTED
