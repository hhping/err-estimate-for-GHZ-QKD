`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ek+xUT0xSrBY6LDj9w6bUagS3uAqI6jU9fi/EqEDp+IPMroXGisXLhdTxoW7hOkN
hduV5ksyxvt538RcSBjmMtt09jQ1/ktluQYCM/3gewuSfemXcyH2FqU0lNzPz9Ne
50q7h9iR0Nl9+vSHqKarjnst5Q6fkzsqZlb5txo/UU2tTKf9HnH8kBmCvc5grGnl
EThjfPoKSMQr6ldwmi7jTAg6W6TUBh27+37/jzAYwEs6iaE9h616RtcuD+/1JasY
Gf9SpRqVNmUygQS1l4dtT9AjUqSeIygVK55CBDLS9PNal6NSaaPxq9ZvUvYH+IBa
wSvHyGT2DLQHVQ0VJAPg7IjPGF5BqRQSTegyYvwSv1Ev7SZC3c3keSXDi9ZMXHFx
cAqYR5kC9rP51R/CbJnn+M8mQqxNPfmdHA0979+2RRZM50oRehwt6GxGlWf6W+eX
6iSQUJyfEkekkuI4ABYp2W6eGyiJ8Qj0yEUPuagnSp5PMQnaTQmQg8Vjk1UhhZPj
plva5xLy8lUz+apyj4+tlLBBdmYxfWQaRMA8hxWOiAeaj03q8RMOREeFQI0uV4y/
p9PPjTjaLUuCIqhwAUWs6mV9w/5MrMj7ThwurTf70XikH+au8tAflRAr2KgbY5Ph
RU0IYVBgNHtuV3uKvE44eJMBei1nB2J5lsKEz6lPaKqiyXQeUdGbPDSVtYulvGu+
yQ9Gj9q+IA2SkmahBsTuaLeBAHYq/KzJTdtlIaNvHjMarc/u4/N0TVFLtGdnjMf9
tRNZXiYBSHN697khbkvMkGFM0ahswbYXKvUU66GpbY5Atyv48uRJP+8enXaEU7qo
xSR9xzIXPpHxY94gf2iUbgu5QPxouR/LZf5gIqQh3VVkBpcaT4F7pCesEj4eVzTT
3EpKXE57u+LqStF1Nr0+IUQuyRcYE1WDsflJT9APXTHUMlNJP2qsnKae86VFSj8z
woPqJp9tfplPuGCe9QuFYA==
`protect END_PROTECTED
