`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N/PsVBQEepxwp6BF6h1jidPiCcUcwajDSGY3FlNEx3l/EsePAMw3Gi5J1O4UM34p
4Usoft/RGb5FBMh3nE8phnaWJXvppui6MZ7DO23wausOu0Pt1PgsRzCSDQJteW9s
gDZZhAMJGCdDT/PbOX3gR3H1onaDPQq/R4smGrW0sJIP2WlfWnrq59dduf6/zpWu
RcLERbVcIoaAwrYB32L4/AfWf4cRePvGx8AVb0RYCBLlnrAHYqaKHPiv3209tDC7
7GmE1Ot79awhTUgeEYCv5QknQCe694mTqoWE3TQJYqauWM4LWcdMBxrCboFH9kaj
lIFvRkuZ+iubU9rxG7tYRToBXz4iRZRLXtyodfowLFECnM6vvieYzgVox9uARsHu
Ge+NZiraVf0r7JqkkrrDYAXjsEXP186qNkJQDsmrGQ0Ip37dVcT/GJoiTukt8JCO
gPL4fWtkUvTFwINvoiimzZ2d6hGQxVPanXa6ZBizdttl9KKMKfcIQ06cb8EJVeT0
z4+MKUEN/g9PQrZWMFXupjhH2nB/dFa9NYIRhNRDIwHrhh5bWK0e5B5XELl8Y46n
l0pw/6brFsJI/1jQsp8MjGD80jRDIvAOk1zZyrlS/6B1OQSqsoxwVL1n4BNNQRuj
GfoxiFLhaVne/cTjv94ja2y8k8HQQomzQVmyZcdycWTijHYa6mZjwbQjbb+fi2Vp
XiKBvDKMwH8M3wtDTnliZjRtGHxSJYmUNqtad1p//aOo7X+DxP7dzRRNcArPjCu4
0M4fHeGPvy+alaMBkn0u6mvAQOMQ30f67Todg5mDnGZ0K+YfOME//HAtdf9bfG+k
TFseOGtNhSkZ/EbsbmgFn+yzKFnAlG9ZonD3RIZTMsdaXBi0P0TsS5Z3pP6OlIpw
HQTprOjlPWCvWeeycvk/vMZnnql75VSj6QEYwxljuRM=
`protect END_PROTECTED
