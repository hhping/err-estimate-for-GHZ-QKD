`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UCkt6JJBD/p1By9HcuAeZyJp+Ct6Q477Kco4MMaYgikD76RWG1fXViXeDgIs6gjo
ZzeKxw+rPCQgvwG6FFXbUo1RpnHEiyyGBsZZ2L8Ttqk1XyAK06k8m7l7mNAD+/B5
J1CzK0h/Dfi9QSoomupLd7OWt9RwbPMgVANg9gl5Ln8NHRiQV9yStsp20fElLHa2
V6J0pVo4EMrf5CYucR8XX24CtPkHsN83XCrH/g7dzMbliy0D39Uj6OPmWJ5kqfLd
cPIPqvJG7YjIZIYhOkUtR64JnP9rr8tjtKxxlJbScMBN51U0RNWjxNqWokQHM7fx
VK7xC+QAlBMNEEulN4v+J7DCmm3a6H3uIFz/p3RWgxkodmBpWDxY3lKFyiTlRivo
3MM0bZ58nZQ252e+Ge72BtZ2bqFZ5OQ0VmkOVFk+ygH6mSFxPM5OM/aD+5z4vb4V
8bCe26aVkBUKJRM5ijhbjQ==
`protect END_PROTECTED
