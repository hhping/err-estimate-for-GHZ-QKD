`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5N5cImQJh5T0GZglF+anv80VStz0E1EBKrEWVFyGxOELftu+rGGFSC192GPop9dR
Iqa96WFWCHJYj2qY+vHgSVW4vfSJhys9yV0Mmt3qygcyHzX3rLfPL1O7acOjOXbq
8cm3757OSZeKGagxI+wt59ybH/WCda4wiFQkzWE97Cw+TZz2rrmjWtZx2lY88unH
HEj5J/fXsrmD8ZNh/SYEn5n/kfyhW7TlW9rGt4S9fB9cRqHyn1s5XgVbmFD3A8I0
3jD1w595Z8fD0IoLZd8V5ulaivpit4WD/Y1PhHnqRxkeAVHbpGJFUFZaiUzsDvUs
zHTLd+EwMg/kzuxrAPLNPQpnXRjCVOv+6JEeLdL5yxIWZjQL15eMvT7J+BlHwSgX
q92uyjH3bNvLTKVwfDpiDkTJ/EPGSxzb/Zpw79cCzJiBKvIwtXyyVMNFa56bGXR9
ylHBd2AJH9KKgOXW91M6FYjaimbSp+fCRBMxrg7rKEBwj5vCZHW1oddKI1LtdPDR
Rbcs9WyG6hNFE3QvfMk7Xe2QuHKHg0I231yot8cxA4Zj6gp0/lhM1zyrs7/IidVc
xAJkSf7FTIc0aDF+B1br5PJN5HTGV5aABgp6gR99QS9Z9kEPmhLj6Wfuu6s2yDko
OiELsxZg9hFLGLJgIJYxh+GQmYOD+t0RrOgBo+lkshQ7W+POS7LQTGKw4nYl++pn
dVMaUOA31RRww1FuKbh3BsnigKrgxYXBYdFp3jhtzFIU32iAwSbETBDiJT0pXPaT
cuHxM+ovT71ijBn0hjz+zg==
`protect END_PROTECTED
