`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9tPKZywf+HjUBDwQTkMcLxod+/K6WFmCqBtc0xCqc653cEMBO9OfZAIUigcQatqX
y+LNRMEOMw6FXE8Od7HG4OxeD5UBWP9izZO/AuJSAnz0p4xhzW62P5j8YZ93RZAv
VtH6TfoetLg130aR2Y0zzIBeEsngCAW9SXhyQJHUPlyqiqlJPmDfSYpDIea4dmSx
9Gd3tUl5/2enQOevzzRef36r+VvGbULH4tnLWO4J9J3PYS1vfKVBldRhNyq9IH1H
fpXwsZ4xuJVNN/+DfIDq0pufTcW3vusA9jwOxZvHpWoH/WhGJq+KacJq2P28cbHg
0vvvwdmOjDukY0d2FpNaCRRviIhmcMBtCwLL2OX5DetMwvGlEKOQUYmLhmupBqbf
71sryzwbZZ69CxY+MvPRfF52iAOKKeIdh1SDff8x7EluRp82w4MlWMhKEvpNKQ0b
3S7wWAzHqyjqp+TIS8qG/Dew8POTdQ1/Xhz47mVaQb/t+DFpEOBrZlcGg+IVGIgs
20HfZF/5o8y6qrOBJ1ItEUVCbxvQHGm980Ae2DOsLoTn0xC0JIu7zatqMWb/HCI8
Gq/UyrT7tlKPYkNd3g6wiNZSOfB8BTcfLk96UwyzmLs=
`protect END_PROTECTED
