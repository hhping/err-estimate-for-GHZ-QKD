`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BfqZu0sjawcBXJiGvpu7WUUlrzXK23fmDYhEc63zGA643FeM4FSXNil9+6IdmwDp
QnuhfN6g9/botPhCayiGN/0c6Cfohf6H44n9XIZ431gHc4Q65khEnJfxVLJ3EifI
xFyZbqAqH3anl5PN4uxB199vp9uxhgkEk9RJqBJkscY+U+9OTJIlukJP2j9wqmno
yK3MItWUxBClGL0bXcHJp6cJCB8YvDtop/8hnotXBX0NNFxfMz3XXSbsy7jwepFC
RhrapVY0Pf6pMPyHx5qICmmiUTdrRxJoSkYbsvXvtAdLEWG7bH5w76KZ7LcEoJhI
464F/3f+M3RR47p/J48t03UUZ1SI70S0L9mA5KbxTmw8qypEdZ5ZoxmLN08SVMcR
JouZpj21x1UKWac0nGLAtLRAMPweW/1PZ31jJug+Qk7txwi3b3c/oZMKksCUB2kA
O82h5mdFx9IJOeTFCnMrWy6E8I/FwxZIxQiOEBS0yFRRRp91EbN4sGo7nztPPnIo
BRYjbwRrGqtCj+77feRtjCHCPQI0ylg87/6OqEC697egdEBe9xuQbpFBPue3p3jA
4vtA2+03233sDO/BOz1RiD2znqDqLDMMNd2wQ/WMZKn37+lyrsTd957gFNDDwb33
GcBvTQpsQFQCCqb2dfnuMiLInQnWyJWk8+FHD1AXUD8EA7nMRUFJCNsMAS7sYmNR
TbG2s81ajHbG8ZjZmXm8mAkmbcMhEfDSMv34zbo9CG0zcLLffaKofxhDEped7rJ2
M2kLw3p6alqFcOb2sojrXDtWGXa+6Zmge92wVFFIbPtz4A/+8XRqrYbK4/pVU0iU
YqtnGDqSMrtsacbBMvCx0sjYWyK6d3pGaxtbKijaJ2JLJs7HNhg0DNHzlJBFysy/
RrR6tFkZJzqfzkziZFXDcSlBhyrvxlKUI2aRBbb2uXKY3NWrHO0Q2IqLRThnPxAg
/VDdL+UaurimKniJNWtSmGyMKuJKqy8IsDxwyhzLrElVqJSsi79nFCQYWFJT33gg
aOodrxUlo7ZFOP8D8EvdVKhgSQ6pQ2Oiq490sFeukOtuw/hD1XaRzERLmd0v8KqJ
3lQRo4vcPqGBlldvXCE8JwwKPILltpYKIyjzWkp1MG8K79Dx+ZkSipaFsnY0Rrnj
DlkYMtsuyrutsE4B3FhuwC0q9Am9t619Si+pPSCgehNu2W99FlFDCo/nQs/q7A41
gkUtpuMhdI7WP4NvdabLrgDppKys5SS/OIYiob7iZfpiR8rsUqF+eFoN8D9x2jc2
XvfgSeyXlL2wQ9T5QgK0AvkdUmi0wFGhKikPu6VddO43VQl02txNBCiHjMCwBJSz
luWLIaLOc6MpZ3sy8Tf5vgNyACEUPTjjmb2/kChpiROb+eFjUDrDfdBk5V5J5L6z
zG1axzI0tkcjSCysDm4Q/rsbh8YQLN910JaiX/Uzn96z1vyrzqb6fhEgtzvmwrSL
GO1BEcUgfYeHDrjXCG5CIooYGcv7HGsVSAR0Buw3sO5GadZLRziQCUPPkKdo6pNv
3/k87CDUVa2kGORa9EIIehiFBNCYKiKjzj23WgqgapbdvlmlvUD4dw+uPkFEidSw
XTIKwqvCFjh+GNutlq41j0YLNMHq+Z7rBwA6l/1LiYrqsDRmkfBevCDiLnqshdP6
ETDatzrJcB/BJmEwzFoDbLV+Qqv45N0Y4nnaUwopxN2fbp7INR0Y+1vkYLIhMvJN
TG9SuVcTtnOlEaKLw5tceIWnLmU4Qjps0cEUt06lcD/98CWkY3YfPFOQw3c5B0f4
HlFEY91LNrlDpYzrmjcv7gmhUyW61EeQgABXZkGsMGCULLSg1LWJNgP07S270YbQ
2CLIUn0qMrCFE+SDdxTGG8FJlu5J4WgOOZ8Q1PBSD6bljGztzX4wHPkBmGs1vNhf
xWIM+N8l8iEIs81eegkd96Lnh2JgsCyjRZKacyOvcrDZkUejqrlQynv4wkKrLqTG
xKmevRLfBECUWZW9ExPRpZpXiNVVLIQ6EAdqUm/Sw1U1lHKYPIpBddm4zU5a0RLQ
TkzPKGRWP5sOlXWBDtEByLBq2cJwPoBWIWHaOf/5BNCKUgyAP9uMsGyueYwPR/C4
DjgHyUnTbj3qeevgA5Ft0SUiiJt6fTiHG/QXygzqLSOAXqy8rQprBlAuv+lpJJ9I
yL+UMtVcFBH1xxxAAfUXbiiaxVYZgU9m1isWnHjFbDxjxuTmWO7hY9epOzcUFVtL
QMBvLXRMRLUNenztWasf655gkASteBeTewRfFscHxFEatvS8+9SuTVonm7eDiJqm
mDzGfa5BzqVwPjcvFWNiU9PPb4lEu92lScpFyjbx2M5Xzpu3X/Q3AaNZf7ARJlLX
yDc/wrGKdkwZM8M9loGS2n0lEm1A292ZIZymXg/Oi6wmDDzfhQ9zbXFs4asqPrlK
S9V1PQDPgBYLVlKQqcwL71QgMPCIIZhxbvwMs8SsDXf8Zjg2vxnHBtIctMCEQO0G
bHQEeapXy+SML5OV7U8WjKC+RTVd7lTpaHdIVx1T7V5vxxuyZtNJQFco4dijgUzo
qHTqHK6pBystjt8dK5JAReXZ+Bx7e9AecnL46b7DBCUdRwu+PbryIbam3MfXgcX5
oHjDfN7+6Sg7g5NKvADrdPkkTxYMceYCzg+mnzlI0220ZhL9G3/cQ/8LbBb1rQSf
Bvg38sCTesKg/PL+YGwXlaDrwcQ6oCUGfS0ZulChiVp1cpGJfIbUFCijcxJrgxeN
pgf55XYwsuHyTOkeJoa9A+I+YRIZa8X0Yy+m5Y4Pgmaj7UjecpL8HwDJnzH7UJmT
dcXRRv0i0kBQiFBHMc5g9cINGNG9f1IimbjIHZNyfmS7OYqOZTvvXrfHVR9O4GFc
r2Q5XgcaPUom2DhMCpCR7dvn2nWRzF8gCMbDer03rS6+jTbJY5lET0wHcsAr2QQj
7stjpGXtFI2AZkZj7BJAgPWGPV2Sc+zFu1vwS8Gxe404CPv5ijePGA7Wf/6qeSGj
AYmDpTQt9YCKBt4Qw0O/voj8fZARC30rhwMeHiPXEn0xCxfL+uvQi5VTkhGaYPby
kG9+901rTvM+cYIaKuClnWXp47A+phM9oD6e7r7Pm8E7beFcrnn7aqYAbgsmzbdM
F+dA0JU3owlgn5ign8tunbM5E+MqNlrNuxI1zN29LxrClmhTlyWlUK8vmhGqHdNI
kenWP5H5rP99iAhSjdqdGXaxb3agBZYy+V3mzPxlWlMUF2kWSmIXzrKnWYNVyOeo
gmpcjdLrCqkeTlwe7uXWRdGkfk5rlc/Yld8urT3q3ehS1MnzIPoxEOqiJQgbleZw
CP9MP/6QVSWE7tdy8ye6OirOmgg33+9ucXOn7LMkp8jmj5+RsZ797m7F+AOB/F3g
15pjT3gqZDMSD6N6B8OLt1qllN8DLw65+c5kDVTmjOJ3frfi5n8RLkhGQYNkxoSS
IdzHgXzvqihxDh6DJOudpv3jhb43vVITrjKT5Y5UL6K7wgbRW1U4Isl8WO21ube0
0PvWpAwUAI4amW6MUjZEV03QEuAqSABdxCQhZHcJQnyJqgKIZ/65GDg5AP40pbYq
16O1Y28oeJYDvHbt34V75SSs7q6BECQQuyl75F+q29lnblEifc0TkZEB+EPvsztc
9jyA2RGBseTfVH+RVuPxf8+fWbFmO16/UzW83tI2E48UHW1mJoIhoMCph9GmPF66
QRu430qQV319mDF2fauOp1ATXBJU0QARWENJa1ilxMgAy+G8ivfYVrsZFycfi2xK
jUYPBOTbuD7IIotzXxiJcoSCbh0oBl+hOKSIOx82hF1lzlYhb+UGaI6JnZFGKUxe
RSZS40S7LYU1FeedtQ+Azm3WZdVvzsDUUZplHZKd48VvWdEzyqqpdP7/afgpCuXp
9PuwNHdKq7yDAaH8RM8ijV/bxXcd21j5vexBLSJjf6TiNxU8qvIcD8k3LlIROnJy
AnlMe6O+4Fb9xR25ccnRuWvy/0HuIj2G2dZ3rllnayqxWUC6LASW3chrQWHq1Wub
Hz2yw7b6EHuV+B8XpWOeWYg4gireC+4oXgQh3HNlHYDL7rvvKF+BcFRU+AwGTnia
9fsHf7He9N8y58b3QjheTxAUsLdKw2QSvtes8TtOshO0I3KpOJOVk9f4Q2yColLv
uu5BnqDtQdZiqg7GgBv37fkwCYtxv06tNsXSZOGROEbv5JrbcIb6vvsY41lW9WBO
K7KuUMdEFD9xs634CnQqTO9dRdqRnfIKL9z6H0dccXQBIA9KCFV8yUh9LUYDY56S
fFvbJmWPWtb5/pI0os98nH0bl53jmNn8inc+/ifbO/h8JndRtH743yie1cU+ACZk
c6dZe/XN22z/a+I6XtKM/p0LymQYPovHar7FlBrEgrbB26PpXsjApZFz3RXJKSW6
n16eSPfZ46XgS0Ek3uk6p9SV2OlLOlqZcYHI5tKYhSQbfDuHlZsG6JcTYrwYSxt+
GloePj2yPI65h4VtKjOWBD7+E5bwalmRCIv7wFkHKMV7ZW2nUD4xCKSfY3SBmcgO
JxXWO0ktoyCDUTBEbd1YXLGEufXAG2jFdXK/eDj2Xmn6mGPeFPmeDShxqFdritrX
myNUwygnnEe9K0Sw+rsfCcMDsxk/wAHz+NS8ObZzzKoZ15ODYL3ABtaB0aqr58N2
3wMXQyoi9RE2XnDEwkXcbFMZ0vHudckV8HdsbvFQRhqSqVspeLPigIygMPt43k6/
RmER4qPtxyNa/IJaXxsNtiSPSj1G2WgjXWBFjFyvRgnSd4P4ygyFlFiFtW0iwymM
bDRkTZcLYNRhHN8mr2FPa+KpaPh4MExcXBgO1t8moa4eAYNMwuuA2egBaEAV9ClQ
0Dr4Rrnq5kosws+f4gsEgx4vLQLEFWytoCmlkRIAZYiz9fDq/V0wlaHKlQKde6cq
O6gz77H3Rjs/y3Hffl2BTOIgqLTEEqXB+84Q8x3KeXwl5zjUVbd/JEGEq//6+uKn
pKpuip+Mk2lYZ31ruL90nMxupkVC/+Axm38dTFvs5wsGWcJnw84Z7gA49+xJg5/y
t6xV5VdkTZabXDxaeHk8w59bOeb8byw+2sxi+cUmgtjG1DR0xzU4Nm8oMgWxNRPh
vxC+dpb0uAwekQ8hiU8xMWVu3bKaZX9rP3nwsNgSR31AVQGPMe2RNkm/i2G//20D
38fXeEdf2HLC73A/B5vO0GkEB3VfBRR7wrFpUBQEE3cPkC2nCdfpM/6I1ZyLizK+
c5BbaFTyWuR+0utPLP53AU7d3NCQFmoS+hks9eHzl+G0nfmrVPcc2Rm9i6sosxOG
P7YWCE8T4HY5OsJTlO77c0InZiQLoRoccA4uSbf6WeXPD55CQKsV4FUfmrJhtosv
PbOPg+06JW3hx3QYNjFaJpqhLhk1O3QY5OwK1v36H9AY7ILokUK9No5rD4m973DZ
W+ZnUHKjQrouN+OMUq8DuDP3yasOi/BEtx6Yxwpvw3W4pq64S6jiJo65TBFvUbzy
cyuvcsNR6WWVBOnBIdAKp1pRUPU4GNwTEfgcF0dJo79/ek8USBIeILbRDX7d2pCi
oXjPFWczVgKbSjl2xvneM9uWEigg+IcgT4dbMlHf/lK/umOYBQYoS9FFLSeL4ZfZ
c3q8fY+YlDiP1RftpxxKGmhN+BD3qOtWbyNblQyJpGWCL69GZd7vwx5xXpWIW/bb
P9bbYjCiombDYppVWiNJdwa5hXeHznuUG2rpehpmDOk8ZkAv+CzqiPfZGsYeCGzx
gvV3Ht8Hq2k/APmB9mxWimF2EjEJ6mwGtJa0M4HZbUX9kaNwR/OFGAEzNTkSlNFb
ivDtQGgYG8tlXzYQU98fSFndJdyP+1Ha9N9NZKsLkOcmD8orHGJOnAAp5JRXAeFY
fQkReTOp5SqiO57ypEpJEprO8EVB2eyJfFHiOZvGUag5WJ8vsI7kgi/YRWouAVB/
ToR613BBpRCUdEEYl0pap6T/VocuoMaUwAxZPMvGfXmTbSlpcMjhMpxUe0cABrLu
VbgnEFVTNit4n8uNEhy8HGTC8PQrx5gC1CW50HDLk62McdlkwR1Ky22T24cE6vN8
ZLyFGWi/pPVWpMJZOYOUKhmm6F+JHvhNovpkWfFQhU6lDxUcV88zy3X32/242L8S
ZmZP+QQSTlQFoBjrLjgmtEa/ovoq9qFyZ8yu2aKY3A4a5xGlUAojkOIm4LmTAEU2
G115zJMJRGwY+0JazUNRItFlxO1JCxyxB0o8+41BbBaogBywP5n5IA3AxFf5kS+P
oOdSRD2ZrROPFwKQru+np5qGh081VNjopgH93BUO3YFxpRywOfbL0gxEwJV2JLyZ
J+g0d7ssrXlaXnyDWJm6G4Ucw1m/hu6l3nGOOtBJ/ByAxj8OlKeq8TXbyO3idJEC
Rx5Hpf6J58ymfdgGDEWbWposcvYurZcRpccEPggF6IpVD3I3uXZnLLfaS58WXVgf
psLv27k6wQg8kfn2v2GK65Tm6bV6mxoa8d7jwPG+yCF1pVvm3aa3RRc6XF2WJquW
cn2F1mDqhzJpiIvIiTOXFSPlozyqa7+HFx0125ZAxRQSjDj3tN5JXu/cRIa3wYrd
wBs70Jt8HrozroarxBO66CpB3A8AoU2DsDCw/i3deT7LyRs1t5m6EUjB2lIts2KL
C+UpCvdmkA/qAKMpdbfBJcpyF/YHf8rcEWvr0dzsqc8TD7lOPIPJY0Jf2OJzEsC4
wHxzzEQCbJzSEHDRpAnVxRdrODA5mrzTvsgltRwxHrZiqHnMVcw6DtexbGDYfW/p
DtYcFfEYeyARXxYLZdYPiHvtV364DIyBJ4ZoSMuye5quYpXsViczCCRnWEdV2dC9
x+QJKI/iwOsFPLe2dM101HsSUkZYWJe3U8+7kbQLOboyENjBXJcKU6SsTmLvHTNM
wH539UxuaNIOdKq17VkQKFfmrbzA8BBfcJ3UH1xBBFnl43df0YPwexj1P9RqF68w
j7HHDO9xvDFZAq1yWTiKVRr4QUm4qWMF2Rw2Hbp6FPpeU6O+jHUSKdcZRBTyrj5W
EAGQ2gOYBrQd7gh+stvzfOpGaNUPTQ+FlGd48DW9VwspA19pIAqg9lSZ/xtk4p4A
ls8kaPmq60u3IXkNm6A/Fb3cO6N8xaVOfli2q9UxCbSLceFUXMXg4lOjNroFP7DB
byYoqa70ZVmiZMB9GB60HSvlb12glVORuQeppkIN1xNh1TBSH64jMy3/edt9a09l
Xqx8nRNzKaGI9BzTG8B9X+QlK3VmvnHFgRBSv25xgOzF6Mr9GyUqHU/XMIhXGtfe
qH5lqJhslz754RfP1QQ35X9H+jxOnISu77qHxGdFQyxqgAtpdw+WxSksZ0lVtHZ7
Xp2FGkpow+aIQ737JR0yJMzHgZ4ZRNsrIyS1h6TCeKGbRFs4moonf+O6j+bSSchc
x9p9P/YZkIo2hr09n5vLPclVTrxtZG488JlRbKZhgLCl45+YoUJz1kK6RJdqvQnj
jJhWX3Wb8IdFMg84TjCVVgQFGICy+i4tRagsaN35Y/TkDwyCeO0l9vwmcYXtWfAm
5/tu8CYkWpxes6RTVQkwyj/rpFoE6Cq6yazP1duSQSsebFY+tIqtuH1Pyk1B3Nuy
mP+wV7nKAQRAcyzr0QQsofxsD+IDxkGLSJRiIQUtZPZZ1tJhNwc+8uunWlRZvgB5
ncXCeWzqI8E+/TecjoGIv80EVdPOEB2ec0oakny7KTVHWutv/nEWQu36YPAVr9ds
bi1H/Gi4vkXqa47rGbsEC661m65UXPmXbkq5k2EnvVLCdeXrh5wnBMXma9Yj+v7n
xhCF6/V7KobOS+GhLj4X4qWFGhaQV/OpY+V5hJWNb3WFKs5zubMeIcUkfRrOymU5
Z65ppBf6qh8ibmw5Mz3l5XmHRS8Q+Frf5exUZMXLt8S8L074ReN5nvNqIlbukaoM
ZTq27ZrrcihA5/X4Z/a8dMl81ioTOEZ08ksq0F2dC+S5/pjqUVvcDvgZrn/1l+Bc
vMrMfzRDxTyL4rG40CACgpwj4wKtEkItCghezWXUtGB833vg9jPYayrMMEHD+UsJ
rzdbc52Tj0i9vFW3WtDY5t6uCOejOGYhMGP9eIBKMsv2C0UlZvX3T3L/OJhB4QXB
AQoVbynsVjiEh37peWhvWwc5T8hP3CyRf10/g4o3Gfj1taxxIvNsgRaAjfqCHd6a
73QMwF1FOqb2QyfGGkJgX8krRBjOydbJf16mObA9oUPbC13rw+rAdr5ypkO54YGB
99jAUVnvoAqFE8n30PtzxMCet4oTMGUjnaZPVE0jHpf5XqJ01OGQ3577YRfBPvtZ
/bTA9EDKx0/6p7GgONJ1yLUTKUhQd3xqTtr06tY2jj8AVkI3YRU1g1rPWcbTT9Cb
JnOrNjNkrU12RYR87A6KQxFcUtc6dde79wtqXQNmEKL2/x3s4stJFMof3qdLZLza
ZNnFmyy4TWlE2D5jL22HgQ==
`protect END_PROTECTED
