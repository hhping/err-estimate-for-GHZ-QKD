`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uzH7//MPc////o9L8XMc/EZY05v5qf1QJsC5TGvR4NJtJXS753IFZhO4RqcS1bys
2QZQmfI1PGUhmCax+76HTYufBGSgLaEcQSi1Me3sCa8hbf77Cow36c77X6NVvmbd
1q5hgFGeGgjdTX/0T5yp1zJboh9Lwiik22a004Du9jYzZ0R/DVrVfQmXkuXGFM6E
8YgdZJZQjJ8+xUQU6ba8Vzx2eDGj22V/dPl1difZuTmkwQshLbD8Po0TTW9JNeBg
q6KqYJO1eHENnWCKLHuqxcbtJgPBzkSWuxNMoXJg5TX7yxsrWEbhkR+DVEq6dI8F
IamlFpcRFRZ9O9LuggCQJSWkdHnVrmGPImbQdRSPtgMsvov0QSHHqNen/OyWtnkt
7PSsbTgAWL8EayaQoGfzc1pwO/0p94KM2pRtICCKGmRKYm795JkCCMaVBz9oYHjQ
OgEDKpFa4Yl7UI/pARkMXCu7T7GcD4NkSr8xCE+Pox3u9TAV7q7MJHXxfKvycK2S
dKboVoIptM1eKf8tXKQulOyDweMTg179mrHAaIG3YwKZvBBAwXPFnuCPXO1qixPH
JvRMLAHjEzlYjfTSuqDEyLWPtJNax+O1FfwD/sWb+nevtAvebrYH5o6Rxc3WurnZ
0AypiQRDsf0FYGdTGqLhjQ/QNYNf5BU0/HHg/wiPatdRCrr2A8oeF2TVEjnaUOwq
+EhJY5tMZr1qq7gC2M5ZIy85q98cSGCAElp+aWM3CVF1IC3oJUhp3kciyGHWW2cn
QaNVP4O8DUmx40cPVT2a1RUMFITiUEmr+FZiAxp5JfITEbD1VtrkLEDKQOgqxttr
DWi3PQfTaLVzB4HwyJ9WW72F7EBLWrhVxr8kNB05Kh7nRPQECslDcM4nSqP41Wzc
4a0ObYrO8HQ8ZUVluuoOJJFGU/PCd5gW9Ohdc0btwWY=
`protect END_PROTECTED
