`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iOkaXxGwzPeOVsrELN5xsNP6fjmEsZPYsmbU0L9p153wwjQjCzCZsddiqBB+7/k+
u02VcT5XqDeipghVtNKAtt2bPrptRCkeTtlNy4DXR1rAznJ3TjJUUKIQHGFsLJFx
cEl751X7V088eflJdUsat9auP7YEM1bj2UVJC/KuGU0ZDynjb7fbm5Xsua3CxRu7
rMfXX3tM6GB3JSJ8hdYDgtefQ2s69vOaTDZpUspjPWOt8Xp/MCGaU8QDiYEfAEKK
XBme+v5PBFHaIVFKmn4WRtgS+AXszFgJk2iPTQ17LJ2ofgcbV3a/5lsREkz84a0w
B/RhAGYuuYOe/BXJwZL7LGKQGUTvEv0qFeontp4PbGZfBHXVWn2B1pWH4MDAdecI
T71cykmlRcnAU7mDdR1UrbZsGWeNElAAG1M4skzSt61ri2EvSahJh8sfy1N8Msp+
8rfl4WZFY9DkuEPCnZIblBX4spyM2hxWWthrb3Z8dr62TBjwVUUyeujdBbsSKPRB
oANzgMI8AqklBEt6caSep17Z6Xwlqbcev2cUV2AR0uCBFw/R4JheNMqTg0eFQDLf
P098kE+ouUOZMGr8zDMXo7bJ2ThndEY4Mn+mp75byETQ57S/gpNZ9SBf+XAOf0Aq
zJ62bWi5fZQrSgSPU8bcuH6gCVp1RaqX3mA/0v5MIJSjkreC+wqX0PwTvveT/DdY
MZoLHyNW66O5jnKDteyQt50PacjqCBkqp8qE3+S9JGXm2wfc7Ktd61/b7JNR4FML
+nZm8umTXy7+toF1S55dZifO0kL612jGxn2wce4O4uMIOmxQGybt/HIRYvYk6ms1
XLf8qLyypMPNOItpJ6sP8I0enrfF4aEuCTpybn/5SHVtmi2Ou2eSLZHKfzdOGTOI
8t6ZrkS5FVgPjqEON5zJGzaoWJ9sZmtc8X1nYGj3KQQVwAPvoGCQcBUkuwCs7xQA
nXlPJPfViLFA83v9BXdWJxn/DVCAXutxZY37kw1G0P2y4ZK2OzyGdM3MoeJPf29d
0kpY83j8RQCi0AwGQ6gtX72OJnJpm/ztmWd6YHd0fcV9ViQarGCWdKY6itwMWjm1
QMYcNcs6iqQjIBX1BK6eD0xN/mxxuMT6HbMONnz7TCAChJRC2EpEoCWkrqJAZ21i
RXBgzlGlBg16PfpXPtDpTT5xbc6HcLmsne0hSkCDRUOiAvR/QPJoHELPYboqM5IN
bbJ5ZSa/fWyFnVFZcFZTx4iDa5SnDrPkKRX7PSZhLu+h1Xw3C2WAx6Z9O98FoaKY
E3TswMiMa0WfeYq46rrFKFeVaCe3cQ/3z0xtSDxzCfl6+TJE6Ng1sX7wkd76Scye
YLE1bxQrLBgfts8Rg7F+fIarU/qgB+DOeFyfYuSqsq8/DH3Gv3xmN/axkriSYBEo
toHsalp+u3nMbjRa9SBSAD/Src0fQ3VwM/2+vLpTk2gFham8cId2msgEjQgWNoAU
cJJnAX7TLzyu+oaC+vr+PS7dpjELrV3PSBY3OkAchYEswEn2wwLfvNgTVCJq9qvb
SUEEa0mS1vJb9pv38ZG93pAbpCmaH5rgO719wwnU7BZUUhpPvU4H+SjH3PxgMOBN
ekXjGKoB++s0i9kjaDFIC6E5/A3+m7SNwc25izkcPRmBqPtxdCESB2czjKs6Ci/I
SriXwgR37tLwb3V1Oj50lkJRHYGBFEPcfEd9XhshoT0lRnlChnJLm1Vz4VlUphfx
TbVipg1B7xuDQmT6kPtiTSu/Wql/GrNyvo8GfejeIqNoYJ9sh0hCT2yrVE7li68t
j9HBcGmIQWCPXxnWB8NkPSGPazB5j3O22pAns0eejIMX97CNyrd9BcmJwYqNyaZ+
vuhu/ECUKmKkuXNR7utckjb9DYeRhUDghOL35nsWprh9Md4dMpo28rRL6ubm1K4i
VJv0SjLR8r1gbvkLAdqzY5IFpr0YTnj4WRqNtowgV6CQ5KwwUv52rVc2eiM0FmNw
NQbNJ8w0j3TXwytw6kvdqQIw/jajyghEWYlh9ojWvg+JKaLX7zPfROUWkiZ5qzB5
N2/h8gVWRHBwwAjVt2T9enYcrXyFQiAtbMsK+4zCrDVJ4KolPMYoepndqAt3h+F5
5DOkJXjyTPs7dGYisgyq2CCNiW+jUFFKhiwitay2iChsGpWZ18gsH7BA5OyzqXYq
brJWs0SCCxUiO0OH0TWk7hgFVX1tbEzqHAenk6i8zlBz2zutqMhjldgzxbaYttc6
A0SvcDPI5aM2/Qd3jyU88OAsplUKF7zK4Qo/WX35Xcx42y2Olj5+TWgjfuR35fPi
e00CmEkQ3xn0htPmFoVCzYXaorru7p6hxgOz72QmTNVqq/ooA+cWaNbT90iTM4B2
nlLtQNDeErjxC3JDsJUpjajRiZZOzLpBg7fwGD+Zqt+rk1z/4nfRl43VUHrxGtsp
rc0axynMZ1ZIOF2pQcvZpWlwOG8xZnLvIiBo7bmWjXz6jR5IoLQzGHuSgj0XSVrY
ygQxjywPbdYsSkyPjFErMs7xO/EJFO9LouJUgS9ISymNFXWjqKHwuRejFHEDw3ul
Eh7gr62SoGniB9unIma/7E9X8PA0+nX1W5ugCw3wCseS0Ai3fwZTcv0x7m0Rp2Zw
772jiuN09Y4kJZwhkauCNZ7RUT7OeeMx8Xa97yvgkhWym4/R0JnvagJcdyhskKE4
NHpgLCU7Ht6WYdIRY8f9MnKm/XIVx0JY0C3cv7RpliA8EV16pW2ta3MclKVQZI+9
Re0U1g6msnQh2jbxgIjFQvUSN9wkd9bp/zBnftE9Hk3vpf3KQXjKZ7WpBF5bxLDG
NWOtiP5/ltOlysgTplgQz1hgkUKqCAlMZ/bLfVCS31g2Ufy0gUjfLmjj5WoZJD+X
5vamp1fwExXyQo5nLr/ifTzXAiW7+4w+vvY70S4ZYq5Y8ZUcqDK0I/D0+FnpwJcC
WhugBn0XhkWXAUOPebtZVdSDxLVypf0Pw12bwpABrQemnqvripX3AILHMr+x5XIp
romiAzdYJxkC2jZrWNc+5+80T3cdq9LW6+WzYRVU2sYH/0VPop2vxkq9G4Oco4tn
7tj6UKcp5K2KnEgfYplX1N38hVw/ngBEnJm8Wm9n9JURSX1Y3Ugt83+h/xV+Kxll
kdAgEUMV1cU6Yzk24RFuhV6NHhs4EurTniY3cNWZm2IJuiIrEEakdO4fULAp6Rav
aoNKGiyUPQxbQHO+Uq4ojJgjMXr78s+i9w/yY2EljEjoasTTNZBaRiNzN0HQORNU
bQo1citeXeQuDNn/squdJzP6K3RuZFaLX9UwqTmMke3dLdYOlxxR6QklWZMXYVMk
kQD+XZLI1PCQmo6neUd+04Fm8ZpU0TgkTMqPJvTXrWVd6dFXjA9HBhccXIqlEV5q
Kz8ebsoqw6UxpE811didb+yEoIBHbdmgjHKBdIJxSRIkisL4rqRlftJh/pHSiXk8
zRGZ2ZrjwkS5Gyvr5IWQigj5zObUTrL/PkwZrWoDci8EK7tz15OtWCLxE64/PKfw
OIentkV9JmDudCxXN98xAsMjkf2KEd4ld8p5vYlyqcnUr4xXg94Y5uuNZI7x2dbv
tJDoN7oJ/Nz8duz5cCcc2cpqFIjzIGRJWkRCJ4sfoEN8DCKaMW8G712XJE3VH3KO
dR1Kx5IULtgPR0SWj/hfWjtxpDsdgg7ScqMSmScaVtmNsK8q4sGzOTmWzhAFUv5g
0Qi6hJNazsYfG4u4k5phmKEtzrXWAIMwL2cWY0k0ebPPgx8Myfg7VISr4C4qXMik
2yE/aQeh7qOsK7MIZ97ZKZu+MnV+r954fMmJkGwCUqjoFztjIWMYUzeB9pSWeU+H
gA/q0njGfhysnJDuT3TNhEfoZ9HlbeChw7iKvOSwSZYhPrefvtloyN5DyfZtUOin
y+CoQW/VA4tDyLiqNN7ncxpOE2XKmMbBAl+TGX8KpISvplV6xdsYnCiqY3epdGBV
GMWv8FgJnkcXqec+Nu7rpINbC93NnP3/finrHbX9qjSss+MMpgO2pZYQrTEo4Ud4
AheSdUQVYtg4+9Ij0WL/ZE0EFQTW/kgZRqWhV0Qr3FvzRVSfwdGRwi3CMvT8IFd6
O2AVjPmAUUupsu5/lOuIiMEbudisWfZawqRO/97/MV/yFtTg3vX4SKiUe8YMGqDn
VPRGxgtlzLPg0Lpbm8Q19XCHQg2oqcfy9GCih45Us3Sae1r6Epwt6v9ELqtPr+nV
2xemj40DErmxuiDrZqWt3RHbAtMWPJLlFNdPl9RwbsAmkH86wVmHbE/7jLG+NGaL
3G3R94noJKqS9bc8VASyotfXsQf4r46X10vCAyYD74QDrzrmWK7eRkJfyP0gKFeJ
296uMcCc9laM2tBkfRcMEksjFY5KVHB9/fUetUsy2MHYuCsYNBHT3XPjT8p/wg/o
+O80/71t3fCu5oVCO1ve7zYPqJHJFhj9P0IhHkchby2Oi97HmuEDhWAsElBShZrp
xFPt91HNNs7vEvLn/LuO66npthuw4ig0r80ztjBlig06mNzg9x6GojOYUzeLbXlW
7I0G1SkaYPv84QkNmRSWxoVmx/lNH4UONgWKNWK4O92WuiN8EhGv8oXae2HG8Pk9
EZPHsWMhsIqKXbafgA2gXgczcK7x01Qo6ZhjV/3n4YTBL6mLFtPKj1JsB9SCYP2K
D2PHqXu3PKGd9hyU4DYKG5L/KxJ3cJWP8AX8wHlDjudpKy1QYs7KOErq5u1u0ZsA
pGGJOoev2Y0qeNj8U4r0LJWoj84XD/rAAj2zyh2kgpueQfSbRXkmTxriPoMtMGZ0
CFuOdTwguc/uMURksUy24ZGocE71ffBc/EDzthxzG65/PSoBAW6Q3FCGKI1p2Nz6
HNPwXFFLWzVAEpk6Tg1sgj+xYoRnSYh4URKCik4Lge9O4b3mh+ga4jl6hFJOUyCC
qY9Q0vDfxSbx5J+Ce68e941d65njvFBC8GSaxzP1+8NOrMhywg3XqjgSfgq0mDMU
zo0+MbC12x8c/Y3PdbijmTw+A/745oDcFSqIQFICv6oSWc9gjMPLbPTqPG6M5i/i
t46yYCknM8hMKTC54KTy4dSK7ERSkcWs4s1YFd6z2+DciZsX55HMVfJffMEqNXEi
mSyhIUNTnWUebfifvolNjysWXBXGO48VBfUxR50TyuWKHDEdCOU48566wnmawsur
tMvLOL4Z8nOMrRl1c8667BDjYZBbgT/iXngskPo/xabxoFurCzQT5fuzQZWZdXWI
lpVgX4gLKqHv8gFyE/uWUUcnpl1SKUJBI0veWvbo2tSkbBZIUeUXg+1YyAWFXxvo
eG/KiXC5uwDWuRp6RV7YN1anOOOeJ9aK3z82blsHmq5b2Rzy0uf9Lzho3TSE2Wny
eiXfrrjt1ptm6G7y6Fa3K2Axf2gRYQ60izgpVCfwWV5STnPI72rG7u0ZV4sLp07w
pE0kbAgRIDYWsuv3kT4Qseh8TMrSu1xY0ofqRYU8TM60SgcO5+uOrHzLVoYpLeWm
/PKjFqURDGhS9WlOpW1uVF5TqnL1lppTbwWJrXXZG5SRgrGLlmgqi/v0YNwF3vHi
4Ne8e/NLTcJx/kXTbplBtLdhZCGzb9dr3LVWdY/spgb0uH8Uccr6zMQjb8eLH4MZ
kTzBuSIkEnPqnA8+Cub9YzJkjXDDTIXnUVqMQ1wthxgGk4RJNShHeMTK9/jyM8+V
iZJa4mxl/ymCH3Nfw5iKZMcpHUxOgMk/Fiw5xPTbt2PwTXNNHgPj+OXDVBecBjss
6u8PDpbta6aGlnVdnrGpiJBrgC8oa/wXp28P6SnBKRlFNbqfR2GAiVOWm7BD9zUi
X1Q6jdUNeFyY7dxAyNBH41bjPX2lmJNC46E3xQ9srpkk+YOVH47vL+TiST5Hf5cj
MvrAcIMp1E9OnzhDYal6bHjRTi3eVsfipJYdH7TIcYLjFRRQUjrdfIgmtHBgNMXq
k+851tfHlbsNRNG4mIr/+cd4t8uZs1EFrgeJt4rsOhGDJOT1nlndzFk1z7vEZaTW
ptvG7RsQGbDmceR5b2jFjAXeNnSZW+slSWAnCe2N2fKLaittosmtBNcAEk41m5dh
YFtn3FozA5R9p7K89JDY5HGY3VQEg6+gZV5Aj76bXnSVbqRcfSFopRS1BouxKXG0
Zny3dBojXdV7aaIYxF6X6DKZGAiyF2HjnRyr6vS7zirJa1dzFvLivY4pt372XoL4
NOWQ73hosWvp8dBI/obtXdD+vyWhzupminBn5+gHXkCjzj+fOhheAbXcnAy7a81m
BD6CTTCggnHsDmc9/jplclUaDXTM8xZUiPWaftwvWS9/ZAbfZYBPGMj1LMnktdZ4
KmU3igKafYCbRD8RwH12jTRdP2ale34xFFwQLkDOHLdNZ6VbrxTqmFPRMzLFji2/
/9SfZQrCezuTitCa8WUnJipB2+Xr5HwK7fWv6nhlV/LUCFLxRq1cwkNaQ8ay7H3O
9X+XYj3m7XTdBZVpS/ZT+cd35JbYmjDF90AeZadmeUkJBJCuI8i2UDO5b1FVZsKn
NVemyYsm3zxyRecpJVsRe4B7RUBdyOAQlxVl9jzJr/uZi1FurZYZO3AzOrprPehm
VVtKFoUEaNACGKdaxvxTE1PZZa1kXS9hryyngZ5mJSpqCmoAY6VGhctJJ/EtnvF2
s1UdVCYyGyoJCVXuaj9GGXxcf/3cVIyeCgEuCarWHtKpEN4NmrtrOJXhwwihpagZ
8vl3WBGum0FOrbKWpJVe2PnTkVAp0o2/jGSiVdjD/5+Fi6vp57CCD60cgJC4QGmX
+b2TcQyi6H6aGOH2jSzgCo/oITXJokjETg+R11ej8TtH1+4skPJ+PxU5BGT1gdWu
0P7Txcketva5Y/S88tu01AhPJjQd6Rdyyg65YY+XxnyfKP+DJn+74m/w30RNJhO2
gXwXc5HXBDQLTtspLZem1HUOG5mNDkgQqwpVm0E+4UJ23R7BSdcKhcTOJds6wsWI
+5KXRSop18MYBdEnqD0ycIXOEkwbekHirFCqzXWB9U+QMbE2g1oK5N5S8kosAgHQ
TEEiW4FlbmVsPejkF3jknQU2oahdKMJwtpmz8ue8jb6zKterYGXblqhweQJVQ0ZI
M8opXOVjYEar45y/2kGiexczB4uISPT3K13BgzPbwgPtiW9ih5w9+aKyTnLCowzh
ZeYDzrl1i1A+bZjkD3kAEAgfQgjLmtO8rGeEzoKmoBcvkQkb72Q2BexR0RyQsSXw
ZwWXPADqG6WrkBDa6oNUVz+m/uivUy5fzD+yHQdKGQcpDcwpVSgzqJpR6srmfXXN
G6YVLtLQ+w5ot/dkTBR2TeHpYaUBl29Kt61nDhhuYxRIIPd1tcURe4YOjWBMuqE+
44Iohr34bfW1ZXG0klgBBItWcmR8EToLdlZK4UNZzB2towugH68OQoqZiqsk/Gk1
g+mnd9Hnfq1YMCqYeP1swUD2WeCl4kHQS5rr5H+P/eR4LEENXgpFpxBeWk7pdphU
urxtWuUZnWBCD9HJgvIEbrcU0L1/fm6sMCM3jHlWmgI9t+3lHsYnq3wB1Y92oFRZ
APuZ/kNY9BpjwSTZODePk6GYoY4Hd2MBSuk07U89WeKqPqno4wwT0z1351+4hpBl
s7YjYe1yse0i/pA9V+7coQRW94Fh5tenJ+wJu4IQeJJE4uzuoYY6EdywjKO7+7JO
HCbkzlEtO1kr7i07F7JXWqVSBCM1TuOBd5ptRqZxi3XTDQozjuaem10mFJiVwxIn
dkNJUa8wc/wOF1Gd26kiBCAQNgUmp9DpHL+639ptIAwUqB8e3Jy/fP26W8jOiDdY
96OhXQMI6zyeh81TVCCsfv8IjKvqTdDhoMMmn+lbl+/fshUmvxjzqrz3gHsw9j8K
OhXWiIUMxyWRhaD9bGehoBhK1+2ONez+xSnrJB4vQYWJgFjKI+d3pLzgn9ypYL/t
t7YscbH+p0V+7cV6S7QvNdmxfIvQW0nTZJBtzUoBEUZANFfgN+VK6SwAKZmlE8hp
NBwQmz4fGNXl1tcpqYv8W7fXEyDLEBqFMSiXFhzQH6s1sv/J7OUCLhy452oSD5rO
pdq/gkLpdGk9qGI34SGZkwvMNS7PZqYSM4tmxAygwk+IU5H/I3/bz1r7Hhzd72KF
U0KhZocEPdQ+4JtIMUZgS3JHCiBDt2EBoER23l6cdH9pBXA2M1exTQG6MFjfFzfO
G67sEJFP4AxtDWSCyDo9oTJXhJx8uYl5lVJw07QG5Lqwr4ygLcLGlvjI3/hMF2MK
F96c47l0qz7XcAtqogn+wCqKIuV2ggqLd4GoR0UD1SkvXuwNO8n/IKwYLDY4oNH0
rfXCeuocQzeZ7E6CxpOGqDjilBIdeRKoTOcSgACHE1yy5oadWyhP7mVNCknaLA5r
43OFodQHrZHFiHVsCD0FsCek8nN1ZhfLa/e5P37AXi1MStlIlEfbB+Giq/ydAW5U
WH+jFecWpg27q+e+l0KId/H2Q1jX4sDY5yEEGBF2JgzGAVTAVXRdcpo0+/dLyeVK
fV8Iyt2YwAksEKHutyI+4MqkyOHLP7Zvi33JiCCZF4BpBBddnd19PQIShlHpJRDb
gZ18a05POzi0K1lflqfk92DGS9r4LUQitphEFNMwvJqbVlQA2WJA+Og8nDKQnU2M
2Hmz1/K5Wz/WvcYOtmi1wlLhGchpCigheManVS0lxefcdx+z0ltC2w8otfJE8k8B
w7h77D885mkWAFZ8iPtWOCQMxUX2ecLzkUyXdGeqtcU3Z6qNpANcVJWLxTAqfF/1
pRRkuaze5BNuiyCoJKuN5Lg/6nj1/v8F4fwHMM5mJwa9+Uqzs4u02jf0/apR8lpO
gr7Uz8rqpVLoV+O0jZnaq5hSAhNClI/09/XFTPTYnCuHz+3a2a0YdX/54awllgem
3LCP6zurfRzmsegSfTQOswE5IpVWyh1TM8IhWnqowYNc3M+Jjq3c/vKQX3rAFchX
gWJH3KPavFCelPTIIUdb5ayk5VkQdge2LF+DJ9ui3oU2ccPfyRhDFBNNsVt4xQCi
QK6KSIS55OZtcMfDrwrr5XYMvDzUaE76Au7nLW64xn9Byxi/oUhwkk55wD0m62H8
tBi2DFd+d7TcKVE1O+Gp+ZeZC+0yjEAnSMMs6SPsW4mLUx+BvP05K75cNX1AvBGD
oUeT6hzXM1sjGlFVuZRVXq15cnSXQdz81TEHxNI597tMLnEb+YV9USuly6zFiMj5
YVF4QuR8ZvjU3BgqKEo+FZi54/aObU5nfsNpWLsWtutigL8Lbmc7WdyE5Xm4gvNM
QRryXGJ8CEtZs0RWz4JC7Uy5UXra8HeGVNsR8m3TxP6dbKoDNVfQ4YA/7v1D1Npj
hzDbCmPU+tSsgzjAgFzPNrIkQAeAlUKGfLP85BjIWNpu9KxxtUBzqVAv7qeRDGjZ
wnoGJP4hGRNI+tLgzgPA1VKx5nuHbXQbTz2fKfo9zMYIcX3p15xES7+RNPScd44S
2OYjpTi1OYwilqjOMC1CMRLF8WWDhnqBjJTvh+Yvo9VXZsQ7VHc05im1tfghUcep
s8ndh9DmaoeEPBqHGRJM7GimIv2qxMiqQq1/fFhn2jZDYuvvtp2I8Ih6seBRffnc
8e/+xDKhL0FXNzUwVK3I79q+Tr92TDH+KLaTJBi6Or9SeVx5vbRZVkenz5WHQhGK
C1qQ1CObGD/kPMJ6G8un32GzxI6WN6plJJh7CXVWsnrmTacgb8Fr9Hr7WnmXjURC
5DIiLkMrupKd8COEN71ucNT5aKRlJEe69oMxMlTLAdiDrCqMzTCgk9OZBT4VFak4
SeMzaFasaZ7zX/ouGAnss8RPHWvvvXNvnO85YErcQPAQ2x7pkwjMwfRIybwYD0sK
Wrtu5kAfPrztrVn0xS3Cl5LO85jfCLQMWzcQNL1nrcbF3KgNa/olxA+BjcJYqys7
1FSXPoTnTY8IrVjYSyKEKV+Xntf0E0VUwSVQRLLmMbouWsnmspWyzgph7iaGbLmB
ahVF7a3prMrCqXdaLg2hOmhuk7hJgoigC6j5DJ2G4vWE1GdNNqP9Q/RTlaX1tIri
x8n1kb6lMclDpXacCu1Xo4hKuj92/YQpsKAhMrZNxBruQlZwW4/xdQUiWsfvNg2N
HWqSJOSLFbvweWzm13OzAjA4/7fI+UACEB3+M2UCx4zsyoFJnbGx0U9kL8+1YKAr
5r21lB8tHLgGWtFxSddkOKW6X6m3lxpkz9IZLDoa0h7EnGoT/H7LcsjasRPMFeDi
nvWCJA766lmHjfiUTBozKZ+EHV5589azZfR7xDzlbiLdHlKTtj+BzujmQbkj+bPh
Hn0oZNMS1AgR0HJaobZ/lT7hiclChaNAr2JkgQjZ5HsAY4suFBxp5BtpJrEeT+xN
hYJ66XJRGicPSKJsUDVEGe+Gt9EQjAVIVkMCW5CBpAvQj5Xnuz0sBBENKqywTQ6h
RvFqDjvoNM1sSTIbTwOB9mSFmhgN3M+IZPQg0ReoXhbPwSK3Ak+z5s5SgHVKJkYL
DNzl8IWO+JfVblA9anbZbAXVDLOGQh5axH0ua2VrLAybQPWrfG+/PlzXW0k1BDUy
LxjQUv+n5oQEH4GcGXZr1D6YS890To6NUzhRSwVtfIU=
`protect END_PROTECTED
