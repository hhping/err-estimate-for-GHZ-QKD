`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mZ/copzAh7lFPPf8jRGYY1pb2cC0oSxEkJ0JnGYPTTRZxP0Ld9Kjj/g8Vi5w4xMy
iQCSXXrHrs+QUasYM2KtuTC0MCZv8KMqwxtdPviZjf00MpCle+qcXVs39rC0oWBV
OzegKCGLGUPnQEQCKtUF2BvrSY5kySkcIdGlYAEGI42vmCI2tonx/krlHcl1/Oa6
Akz4rEBOT+ckGS7beqehEgMrkpxoPlMc/+0IBoKvJb3ykEBPW3OY2mauE5zwFiQo
SJ/6Bji4TzAhjl5cwaXDH+MQRVTomXQaZ1vBzWHH/ArFfNTgjS5aXoOHI8MzxZBF
TrY5cDgheJ+4yZXbyyKBSpTF6p9tR92+xEd2ERGai6zEGP5oGP0ujydaMGHnGR7/
KT9NLn7tKr9Mu/GwGegihTbSQI+VZYOpHaP0iFY9cClKsvcYal2Gb+W4wFl4tvvd
yln0jWOZk3llfBDZ8iIJXpyCrkKSb9pkkz2n9fnNmbashSjG8R39vpkCI3Ew8LUu
/CHnwaTdvbjhR4LWI18W0N8jF5uJoyEafagOabxKyJqHdkjOz/+qLplwcFuzWVqc
9XGB5XzF3DtY1Ckix4w+xyDQ7ZQIJrlej5NHhJqfer8Cc+aU7XE5fczijeuYiJAw
GlWjwNw0bpgVr5i9u0mN3bLONU5/UediKGK7QUFWHaLj5idF74ab3mo5RHT+bhCh
qi7NwnQV06v39Pfgqa/+GL7jES9rtSPbH/pdegbkmwYs6sOgypRy+PDwlw5K2tPc
lvFJEi3J6VTjLNzB+jyspC7ggipw/TuakYK4JtiD5nwYquMgA6bEvqjrhJ5Z0mIQ
fg3U4rt3XaIpW9kmGWHNfDZSJ+rC0RZVahA7fhJFqwKOlcPYGMFn67NM1tp+smNs
/tXTPBYhzWYRC40yon+bJBUmuW8haFI4NsLBsoaoifJesCceyjHOwH2WWbWBsoOu
wPK61zOuZK1cRkruENSciDnzB9SxdkEBZHNah/On0qHyLjro7mGNDHmuZ8Ytuoj+
iU3RQYJBdk1cYgQ5HMfsRo16lmHxfD/xQKvOXBOslkrwQzWrbvM339Wtls7eZITa
fefI78Zk+7mqQHS5awcfYuDU0g3HyPScadUh6pZqLBJO+lpFb75rBiqdzgqVpOgD
DZLzxXWXhNzu3HB++HK1LxmzY5Kj7RbvWTW22kYhchA0ySE4cc289CoY5s0pfLwq
ipHe9WEUAe4oE4vr/EJmIhDwAJwNs3Q1J1logT503hQ3lzataI8pQxT5/Vx3qYv1
tbWq1pJiyHeJ1MAoImr85cONBjNdPLQB+DsMgN3zAe5rHcJqfiJ6729mjvRUHbAR
wD+G2/YOnYsGebIGpB6EMJmHi3SsHfLgUnN4HhHK/LDCjTqJ6FyI8KWIw0lgtYvE
MoE8ICss5FBxTKC7O9g5zWcFGVxMepbM8TVyaZ+6r5GnLInk9ANpzQSickLStlyE
Y9FvgF+/zIcQ3WfO40uOLZSgfisJliJTXSLZB5fATpcyUDTWboS+OmBCY3gHWSs+
3WknJZfEulbrrjnW1b/qM45yJCNn0MSl0YEYUSqGmSDNN2EWNz2HeusdYaz5AXOo
7lSJ4p8Bs0w22/N7Vfq/ExAYwc3mGl0vBlnIUyiArylFoDV6fwbnyOczUE5odgLq
57mwBmohOkf2ZE++mQ2I1TiX/fBtmj1HKFVWK85TEzuqHmWvyfUF411MVdIgBIeS
YkcxrLSGbh3SwXbBk3gzsQ==
`protect END_PROTECTED
