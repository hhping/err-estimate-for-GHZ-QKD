`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cNJdRLhFJXXopGdshfsDeDyzoFx1WkHbzHq8vZR/f2bwGUHNTuky8TP97GMCZnXx
QXsWp/6/nU88FnnI2TvcsjASZR3pP9SC0Q8LyTpByK77mHEh4QvF0xZRgpCBoVfn
BISQYpiFg3TMRBWYJSTnBUVs9Aqhu+jwwn8bICnKHbVuf9KLBv+CCm8uEvmAK3rE
6CjOSOB3PLKD0iq8ON3T3/7GkkU+Jyhb618GiW9qi5GubyZWVSTaFk0TLbH8ovHh
VoeAQZvRkiky6XUhSgBa+1SykRyQaVFuWPHy5Q7mhcsfemoEXzjvMFNpUOR1+9xa
MWmEjrTuTwNxN/z/lXW1X9EWwYzJz2Wp7u+GcDPmtho9rF8HNuKxF47eBHOAHIfJ
IwetYK3b34/yzeaykRrA06V6I/YHfisfhKszjiLfIb0QSgAwC43lOu+9fs0R1Y4k
Ssmp1BR6unhMzKxl5A9SaXdbFzcwMEm7sbm2weD92qgy9TmgyCREX4bCPdik0OJ0
g0F93SLcBw4TMrR+ItLNeczqqtma0QrwSXwXi0BsVBoDhvm7/Jb41ewRIaiUq0DJ
IXCSsBjx8v2sIfyB8/Wot4fjFP6NGA8JmRZ1vJ3Czw6S62E8bPh0wApBwpAR4fyg
y+3defLWoTqeRRXrMD+it76cgxt56viVonUXYQ1kgSp1eTqLo0N+jM/dncx9hWXQ
`protect END_PROTECTED
