`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vWxTZzxd3qbKUnH0nM4Iv8tiZ69WYXq3/0NcKeJT2iMROOplFlM7qEgR2eHD2uov
WUequ3vaoY+qiam7MC/RuWn9P4GPK3iYKDE5ggrXgQciasitD4FMzjnXg5PmnU8x
J1p4U8gXFYahya3uI0zai1MKf9FY1uS56zzSz8JVlN7QMwRE24QNfO47vY+D+/p0
B8GPdt5kjV/bywE+9so088+atsgswk1cuMU7TjyoTj2lgZP+3Gcqr0j2SmNJ/kBW
7DmgYqdFmibHOi+lCTf0Q11kTE+ETMgLX0y1XKZ4RrpqN+RvDTVScFcbl82esoRQ
5IJ2CJzmg5kY6kpmTd4zQXUC2IKzyBSNyx38gkglp9c+HAXZ9XuPDvUcZdSjihDU
kDBNQG66JjrJNp1XpIpJUU2bpebxgZJYeMjxDNu9lG/gnHAFAnBXNBHkBlc0P6zt
zt848LiTqwBDK47TOQqz1RCB8kqC/4pJX/WXG/0WPFyiGgEj3mH7qr9U37cOTOce
+xBZF8EM8wxfdgXBSTyR1Mgj16F7gqkSRqkjTpX8c7RpJqP6/JVklElSFu0+GAQT
uwnG6Jx40L3sr98Cfsat8NL+O7a7Xz4NBuxYS1f/185loHrnCW413nqWZJauuTov
FOWJwg8HloohasoDL3nfMkuRJ5wOEG8DSMPQC18w+D5aTHsVQ6jq98CIMhL4G7JR
YBojG8KI4EF3ByWJU6a6GDypISmo70l8clCwJZN1Wd8/Gsrm0E2v+OB/k+tRLbtX
9i24XNzlK4bqy0kG+GsMuRAuY1VkH6VPiz2Pa6c13IsamzMNJr0BZsyh5lb957d9
ZprxrhvTTxKKoMGYSdb8DLn4cmssMI+FDiYO4Huhtt2u/4m0WUknURAhyh2W3dfF
11f3s+X7tEFr1ceAlRuX3xcblYNLoj9MTMfqNvbHPGb46aZytS7Yq88ycgopAq4x
hZFGxHUKPyRzMkx53Bq4R0RdXg6CFUyLS8Dt+h6c9kPeUQHOqkuFzSR9U2PMJPBr
scjjroxE31oW/4pSITabJ492v/K1rBP70KeteJ9wVQf+yDWA9hXAj1vkLt4FsyZZ
pbTJpsaFunF3tiUx1Vr0l/g1mc1+NYz4/KVcJhhk9bx0ReWfkkwu+O+8FH2SeRXQ
`protect END_PROTECTED
