`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NakbbGuH7zlrh53082JezKmkJa1//0TNVsIqYm2cPRVDp8GrHtfRBmaJ+sCNPs1I
7l9MJTXZ3cbcSZYEJmQ5x9KergEXK4g6xFuzqzv9F1t4QRLM8XPOOVmLAUptjHie
BsmnEGKlsTXmIBwe50l9W/esUFx1u/K6w/bMCRIQot+HPSA64dkWXAJ+btMIUKQb
G78/Zj4vZMYiFVMysBS04SlyI2JMLXflq/Npv9VVlkIDS1st9DPz8F49cogk9+CL
bhQ/VV1avokJ304OiM2EEwkoiA/ECytbFqsPbW35DnYg7SaAX3MEVXwIvr7cwm2m
ce8RqNhGoI3e3kwm4JT5sb8sTMN5e8CSLtWaK7Jk7yq9cXd6u6X1xxP3emveDSXX
zHGlzh4LExYZnHHkqPLyBGojugf/grqtrrxXTlWsm9a1JFpR/9qXu7+GCebNuthy
l+EZBAqJfjQhb6qfH0AR/w==
`protect END_PROTECTED
