`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yzK1dLijpqQ7lNeh2hOc6Cyv76nkv+OuM41RFcAsLqSN9serVYCGT9NBOFq7DETM
SWyxGf/MfUOEtwhboCe6HncwkFkw/D6dODiAy6UvESobFN2RU9UEmk2e0UzrML6C
RIECy7C+q7KB/UxtahCfjFOF0tzTsAilozuXgKj76i56x1TIaFyzc/ZNSTQ5xZFk
fEONJ2kNwQSEN4yGEnvh0cA6ukOWCTPDegPVwm2Ttao8eqAewYKc5KTz1W3eOSRR
ijmPq1ktrMfw58T7n2AwuGxC2TRTb841j+AX4Id4u9/edkIGjVhN1csOBOgNzSlx
9PAut04hGY2bQrwUB/eEImKu4Ts5HtLfvjB1F3Lflv8RGhXP+gnnPLie33Iz2/wU
FzXF4d9QNprL1La9Jo9MD/5xsQ+GShyb8lXyHxzlwy1SWby/YBbz4IhGMVqcTlB6
9CpiAegKjzqWyc7alXxyE3Df7+fg1rb+okNSvAryZ9eSEUDB+JPubv11YP4kybzj
w8IL8CRj413noO/huYChafG6L5YPjRvBDuW0qT8//NVfq765ILw++FKWiMzx8Skq
IJUvlq0V7haxSUnFK10AJdExONl5F54HX4NpvDE3YY5jucYLHQrcKA6rCApNJAgj
maJJKxs9p30W2J0JQ3IcUIkJOre3EFZsHTBFHM4pyuII3V/4/dDFLTQ8tMNV/rbJ
vGjKV95iiE1MHwtSkmNn5couGzY3BBmAF+9K9B7vZsO+u1YSr63c0SykA9b/T0LR
jzwNFEGQppNNmQCGKUi6/PzUmaTAN+L2qSYcq4V0RmBJOtNlCg3Pq9Xp4JnW84ao
oyO4CWnVm+A2uIJzJIg2Yl4g/rclFyCVsFO26s6fC4+aNek2mIEmRtg/b2TwEjmB
8G3eBNOhROeRcpzMC5JyVxabxMWelhiHCSVyLMPrxlKMl+4b01M+Y9IEX+GD6IaN
/SskmTynBNDv37fbQJ7Z81hMzYWL+UlQGzrWOQ8OReiqM7R48QEqsoeQVIKZnrCw
sJZB5SMkYQGg7oTJ+aAhYVFc96SmYNod5hYajQfQyg5T/qGeY9rLah75wZhe0jrX
knw1RDhxLcbRwEIW1C7mqBKFjgUD+RqNMI29weBqndi3OwHNNYU3vAX2pJIir5up
amxYubiQOT9cWSlPLKPUkmEgIxCZ4nf8G6WQgxUOAO80n+cb1vKOeL4kl+eS/A87
wjyjeg1FhGGdEoEvCpTAC+9LKA02s7IR2SbEPGOgkAqY/uVXDGaex5ZTq96cyclS
jLu97zCV/7MuDgofGrQei4bWzReXB82gu10PslLs/QP1MmHVLPvFOxZFJgodYcb3
giQ/Pw2P2xT5bMeJOzu+4LeFDNj6HffCzWNH1YhfROW3okC+4YwTA2w3dG2R8MVA
oCOgfXyvvEw/AoBk2MPqW+e6RayD9VtgiHHlabiZsV12r1jyS8j+Zt5oQfGy/eSA
WKhO/m+ffOqEwJ9uad+t0af6W+SAuoUR93gAHpbXli1YrSxnpzFix+GkvO50EoO1
dKMFEOlXj+WiyAQDDE7yru0c16aCXTKb/+i/BmDxpPgfYvwN/kO4z3hhq8RsKLok
tG2Te+ZaglXniV8ugXk63DpenMbDfh2MxzUUHBQ84EKPyIPudueSFUwvT4slM7eS
yF58ieXkwruN3LuFUZZ47zbcqhQPRexZi6zahF80T3/637fkFZ/sDtMAvoiVAikA
3HYUQrVe7XrfgBCUpkBjl9RmDk3jWiPkKZgciaHg8vjUTeTSViSIqL2Byx2pc4rx
NsB2q3fE17+BfHVJ18kgQZGxxwTFlXoCOR6pbEXtBcRCzAqU+1IiAhUgRnX0BZzI
7S+kUjNGzbRcV+lHvJUcFlD+NBzH5307ke1hCmMIfKfjbRQexVS1bqUeNKhZLGzc
CfNIqaqD9/QG9IZCqfKpt9YtQ9/sVkxpfvCFKhSW91xPWU7gEFqjmr9bV1nYc47k
EO/vVMEJRm6HP8wzccdq301C/s4iDG89ugHnqJGV0CM3GBBG13WOx/cA138y6Gmz
XZ84XQZOv6vrjMGx3Z7Ihe8p+DJgAGt1JycneIvXZCGEVjVDhgRdBFIorVEvMdSF
9Wa4huPWrDRraMNKqsFiOjByaaBFvo1G2vGTEa1Q1tYeVu+Jc7q+VGC0WIWsP+kj
C8n0k/idarNgNO+F50HVdah2AxNHhAnVvFeHqzgVdG36jDIq+grqhBP2p85d1Fy1
hHusvvzVrW/CuEmn+ABOc3aC4bJvFP5AYTrW9PaymjJkLCxRu48eP+Git1+FcGZy
3eZMR6hJpoHVOvkpziFCIGuUQqCPbDSJQ76OTgknoWfnlPsaLtS2HmL5qJoae7Fe
nIGauxGnHrzJWuK8O/i/spUDVbmICGMe/X75JtpRTG/cW0Wr/2UxOZ+7rCMxO10x
pw1D2miKcag+oMTyjnaFFbMcK6yDUZPOSuAAa98MZwdFnN/jiptjNzdp9tVm5u/H
Kekj5Z2leMgafpsqHnSSWEbl0HQGpZROUP/2hEmSBAA=
`protect END_PROTECTED
