`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bZQW12qkGmRHOOKqdurxjQC3BTaku/NeRGIbUL1kraI62V/oCDna8QUafZPCLi8i
AxkDGQAl/t5hr59iEzDI47b7E0dIFAv1PnYiA42yl3HGggutJL24AjqFBja/e/+X
v92TjawiObLdqoT9mowdRpI8tZy7VCHg4BJAB5t2ZE8nfmcog77UtxBn7OktSNdB
6YUADhV9SN9EX3DfYy3L+/uv5xUdUO+I0ni1ynj/P6puACa+uQ2eoNwj88RwIfSG
PQ7dcjArHr0ZyFDkj8SXGhjKvAe2qM3BwvsS/HmxO7Wmi9PpKXuMcaVn+V8SoN5M
VInroEK5fQ3f2iNz70Q1ho3UQHZbXg4J/zYaNMQdulJ/wk6bmEugo9nKLQm5MjWt
Ljeqkh28F2LrbzuH5zRulAS6C0ZEuYsRBpwWmV4ku3cielB9sxMC+7TBZiSDPwWM
RJhyrb1/4UjHdg4iWzNibh5TbF5o/G9XFmNGN05JMuxtgRPtW84/85Mq59HgDSgm
Tc5nNt25UPsAPnHe797ijNHB7byLMMkUlCBZDzy2EJYESbBw+Ohtiy4LEeGJRL3s
2oStP+eUZ20Ured0GFSE4hpRSG6CBGxf5wjGXNZOGnwSdLVxH10j2c2+oCW0uHZI
QCz+2VyEqhKPrh1k5kPNAlYi9SR3czXBCKDhnTm6onukQlHHHLRokfDEO0+gsZ48
2NeH1ewnyYH7Kep3isV8ZYJbsf9lIu/VRdqGwllHiw/3Bll/HupvXSeDkHN9Rnib
Bb8kdOQokj+NUVjPh4gJFWYtHsdiIBClLZ6KSeg1vAK7hC9YbAgy0Sd/TsLo5Wj4
J2u3+kcRuMZ2ZN5rpgXtpHeP+Dbj6pdpeQaJ+zjf9ySQiyEepm8t/+0wQcSRhfy6
CDOISh8gxPiCLhwZ/IYFzYI2X1yis8NDBJt/yVyNT+u20TbuAKm7wvAcnhVp90YF
4QVwrKhdHC/5uEKNuyq+PGX23jRKL27dg4IGw7U6U9mJ3sWmx/4w+ueQc0qw16dM
WNP+lzk/u4sbOwYG/Vd5t3Xeo4uU9SER6XL71/As6vSFZEqMftNIFTgM3/Ng03dZ
Z+bxjnMZl0Jox4RINZsM6lvF7NFiBQqwHdiTzYfQIdgQCj0kK93+5n+qEkQ7zxDs
jrMJxR+h2QTi4Lcm7rEKlTR+P3N/zH8pLrUGVFdYElMnhM41ffObL7ILaQ0yW0Ow
crW/4fFBnPvGke4nXWanOsgkkSRIh3f9oEfptLPByRQCoawSvfMVbQuOdMt1TrXh
ogqcz0s2wnyZ6BWNgVInDoH+dujpPinkicIbeeFMVqrJVLAYKNZFmzsFgybjuG+i
221Lz7/jZ034GyvJDSggb+vWw+S/YpU2zEO1oE6EAD/KUOYe2lzfpuSaGbGmrj6v
CKS+Pb9JlFfS78+/emktzxBgg5VO4Vmmo6gk5/tN2iztdVETg2rwoWj1Czw7lK3v
F/5ZkOxSiasGFVw7sXGIwsVFCx4mUcG2r7RVECFGMFtDJpyXrB6bPi2/uKzBmJOR
7zKbY5lRXWAr5W3WgjjYYQ+qDWIXOqdDiS0W1Epc+9L4uO7hEQQxbxKvNPbCaM3F
xTdUx+2pqLzX6PRHEe/HkALAFRYL+jjrjDptjaJtBo31V1eFuMtwdLI2p3X3tICQ
FnRIMLa0xrPyhKHweHr90/3gMuLkcSAMTzwOADOCJKmzE3Ym3sO3clmbmgQ4YzPA
XZ+/ZDPZhcBQjDmLkbhEge+CwGBuMCtJKds8j5Reoy1w/syDASrV77Ejd0gt0T7O
P7dxQZ37r/XmxEcGGAb0OBbKEPb64EijXqM79L5nNT1N/Ea+T4Pdkz5OA8alJ6DF
AI8xXcp6Qo97uFEwwb9+JA8PScVg+kbQ7Uz0QYPCkVHupuGAvwk0tKsbH7kHsWuH
dCa6SYP4NRpjJ0b4HCx2IeF22VEbk5qX3a8q4U+qA0DOGLiZd7nF/aiQyRIBvqnu
mZFUIi8dM1x99l19LqoST4r9eBauJiiBmHoAiTpF46k58G8Wcq3zTN9BlOWchLro
m/K9KoxoRLkVzNUZZlrVXHgTzi5aCwaAMmGhnRLE143VcDelKpG0lHaeR9Zotsfu
DlB44SQNcyRLe7l+53aMYBCUU8BB1+LUDnHzWJY65DAKv8HdV6PPe7TmErGBdqQm
Rin3PcCUnyaoBsLXvVIGCaapFqYtWSpIMu8OQEbwzhnNmHIcLBxys14gUmXszFhU
qqYz02FcsQkEJ0VxmeRTf4mu3tKnt5vearl7iQxJBrxxqRBbFT7X3/4jHncqc76O
UM+I2P5FeJkkIJMCFiY4YUFlXmd4+sjQLwuhb1dPGhI/iqUWO8fy6VvBKM704jfZ
4YWFr1HpQbzVVP1ffMWxieLh7HKo17+/7773csnI2ONCoYZAB/eHYaC6UmhUMG08
qf4bIjYUvNHBgFTjK2MmF3SmlH5kIfj2aehm7k7Qms9FaZQHCXKe/FgknbhMPoie
pJvwe2a213BY8ZGAVTT7XHbyGTioLfMXbm5VTTU4p/2ZoIcCEmu3UwUZIgxpUB8C
IvTRF2y2gQr8B1bcav5E77o9SeeD7zw38Kf8OJOHMGa+z+kLt8KPoqR36WdELhok
mR1Niun6AXFDUJLklrx/6yivnp4C3ucp5AoGfLcc6UYWs+Q/MdnS8AFdvnagAfPl
PKNJteFl8mBguUfmdV0cIqpFep9zQZbo3O+za8hHzzZ84ynsHu/hMRMnlnxWXNg4
arFPJp3/CAad643fegWiErpJnblFtYeipo7Hbo62sEwWPc8osFwQ1pfRcWof7PYq
`protect END_PROTECTED
