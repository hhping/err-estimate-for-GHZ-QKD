`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AM9v4+Q7cKzLviV5+OUfVWj9g9WS6XEQ9esX5SmAPxYE2ne7hGal/mzEp6XO1VPi
dkgGVmMsPXgR8wTQATAbF8sd+0Brq5UuFCc3tGA/v8NeAWm/Npj46PTdRyWSP2Ab
uDlkz8c6u3ftHovH2eef+2KYWeItfdNKO0DNt3FrcAiEfWROnRtNmBXjSu4rCu3/
xg2LpKfAmcEURzew36r5T2e+QPAgXsrctCdgRdWJyMb/hm8KoulGxqXJSTwRuZZ6
BFmkWp51zgCb3kdn3jxKjauRp5AoukyIHfa3z6FPre3+VsqFEThtmQDnOZ3Fo4F6
oS6McHuWfhtOi3rjWoaEES6xHI1Fv9MTzMof/pKfOb2ycbx8FNgoeqT4WbatRoX5
Gx8IlquxE6PBt1oe/gctiTz79U2yLxMzyct0HwFGYT4BA0v6JrVEzMzuI9GJN6j5
cgzxTziND+MjvW6Z0xzjOpGPKZLCcNy5oUffuDCWJFI7ZD/NSjwI56welEzlF+tx
n0nsrfjhUEeEygRGAI4MbWTSJPi5dm2Nv/OFBnLyVgTniurZKfyAIXPj+Ub+5MPL
FmfAI5aGSbSGhx6TK3r3aDNovZ8UChLqTw7Wln9KnkjqLj2vgWQuSNJnG9TQhQMI
Gu5nPP4gwxWo/NLfetssxKSf8rBKuQ3tm8hzVO3A+ak=
`protect END_PROTECTED
