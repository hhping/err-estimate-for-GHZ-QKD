`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gyQoU9laQC8SiNShK5HCoBMj/rPNG4H92dvdmMVUlQMmiYyFNsvN8ID0rVrN9t4t
DkI9Kr5PrSdaQbESW55lXRUol4SuOUoDEo9SN2EVJCLmznv7wI818qN8uQzQNo92
QJ12h/ZBJZ1v/ZAgBdHz9Gm9Jaodxvm1RDIoUzZqA6Hj6BEC84yfsjt6V9pwjAQx
YbwaZ/KJrLdP6mjvxncRcie8pzk1Xa5CCEvOvqvPTMpzNV16KROHzHlDvYMau0Ec
oiAQXQE/77bY1gZlEkhdVlonW1aamB09GmOATmj92jsnICHenrl7C3uiZhVdYG/1
iBiNqBPPCJf3tbv2A9W6oHyZrt2jTB3q7CY28fYUaiw/ReVEX65vUZ9RZQPPRqBi
gbRVFOD29UIcutDcmFxB7VW8Ew0jO6uGcaKunfkK8+eCYddXWNChfc3IenbSW5xB
DQSxOE2NKymmr8eObi+rEQ==
`protect END_PROTECTED
