`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bQIut9EALDjbqqB6nQF0Gahe79eVy5jZMlwSkVqvm61ithiqntivuDYmY0OL1W95
c9/OvaGAKWnYbZEeIF8grFMsY7KLv7DCQJNiA1u6b9itLuKt6o/MFhchirgCv2UB
rdaqAFfykc86rJnHNTQHFYafj12DxjkgQlFmp5Q1ct9YCcOnXbg6lyxdzKb0VIB3
KCC4P9KhxJnjBcNRdpYVHXJd3htbfb1+uEVdgGSQXEeLNLVIlqXfqYyAKVM/Xefj
GrJS8Y/hbHd/M2n78I4EehNONovM7quuWTgtAy+VBlhkmIj1c6Wp3OgfwsgSQmdk
E/GuNI5w9oWWJPPyCfYIi4cFhp8UKePSJGSvEdgzBcnElWxRRIQH66kS0FTSiNpy
t1nMAVBwI2Bc4qOI6i+xURskkGrhy5LtmX4gt8Gb/cs859vzq5mCMYaWG3Y3N5/l
GlHsj+odyzUJbMQYEsGIQiwxm0EN1oprUtY8kyiQ3qMFBn7SrsmBar0nV/TNeNUo
hMhSAul0KmNWO8trys+7tUJRc0VQucsKgN0mNKeePrXhPBXEz/gzR6ccL7+KgWw/
n9JNiP+RJhsbdMKQQ/FqdV0snzPr6G6XJpGZYWYVpCP3sCQuSQPCOscu/BoEKTrS
AOvaOhNl/NNw3Yo6BGagVS+792r13OrMzI4GiMDx6lh8Z0dSxJPzU96NbzMIN+sc
vfjgIt6Dh+pIqdoNtNQzCCTxKstDqzjWW0jmHUyxfkuq2Em0dGFsOivNuLMSpPzv
hYz9Fqvqb5WcGWf/3Y6sXKrnsMs0OO9tahbhmUb+N30UQKHQFwJMfHNqsp+wpuq0
gJ6mBU2jSfbRjlzi5zL92eueLgKan0mNOD08qw+bqGZQOtRz9Kz4jOlJvTJRWQsf
xp8ISrWpvYGyVtDu18tf0XFLHHLUP/jvgLOPjg2NdEwHUz+0EOylIr3Jd9+HBWhh
tJWO6JzC9SM6VEL0dN6G9YlVUmjaOdO3VjptGr5NNbbKimde8dplNI4j0MojS+t1
JMY9yufhfdwXpb9mnkOFzySr0NzEpYPJ2CR5m6MbttYPO2HhC2+sVS2iwszwNQjp
cAk+1gbOVxWdYUu+w1Gvix0jeXZBXxsWmIQifEzayKsxnCDikDs7STgn4eni8Sbm
HM/z3+YC9msY/6u5v19yO59fMYfPom9r+MRpZOFYpG6qD7po4QIo58BUiQcgwX1M
f5BFBNlpM7U11bfKvvsUsAALZzaLSBIVxYJe4C4eVUTHdAA7ewy8cgWxoUYppILu
AdTTDJzZ8bQL8zUNzqualcxIe0FkCtd8K8pV4DwSkuW5cWn+mKd5lS8RMQbjRH5z
F88tWYsVnF1fWivpPdfEhRfXHc05QG7qoKNO/kav/vqYZ3V1drYKoT5FSVY4hcIb
wJ5z6wS0BJm5VLHPo9Hth4h4XhXvXJ7jYnNp+kw/OOT583h1nM5GNJz+vrmqaK6V
xMd9SFnY3UXWWWgn1/Mn85CWMIuo5dQox3aP6DDdU6Z8c14g4mA4SwAEtl9qIOsn
d5QqhQRAnMlcrfoB41i5/594kmP3vtVjxnfEw2ykjSqH5DE6V5qxVrYLay6JH9+W
q1PLrKi1E6QfDMVKQkw9iR9DClhsilGScq7xq9KxxJ3kSYCHZ+nUO77SKbyU0O69
wRrcy8/Nd+E7QJaAwUTcKoSJJng2BBNxvsmqPtyr1BHGfEWFBluXAb08IJI45beB
pzQAvLvquR0rFHTsEllWJY9ewSz0dz4PhCuXVSj+RRzZ/WGXBN9DiEbdvcr6FTK9
JqjFZFY1HwsSW7YLY131NR1wnWRR/5dADgBTyKANoDafEYTznErxcmYhgzO/ZAnX
ihH1Ofy0wMluwayHrn4GnrD+nbz6T3Jdfg5IBHC6W6RU1XI0CY2pcP8Xk5fccvZK
TdcQDhdjJbH7YV084t5RKaJCW1ZaY8R0iEcZ9LGI8fV5F92ofpFuu7RURdWQ6AYd
z6E0H5lblR7kLS42QzT1tBuscRkTdeN128W2zh5u+B4tRy8UfPdWW2pGvBmsSDoO
lJrkAhc7EadYtouKJMjfiAkxUeMw7uOi85FJWDfFZ9xTN3c5jWG8vBL2gIVW7Buf
41nqRqkKIj/LSyLTvmMDzQ==
`protect END_PROTECTED
