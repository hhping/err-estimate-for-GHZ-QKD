`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IK43GOH/9R8L6+zQoYyngMji0o38xVEsKo7w7WRQe6shBcVDW2xsPSk/Xw9s7Y0Y
JgkxNb2JfC+iM2vIV7jDzUk/z7PFTOFIXHl1RQ3z20q5VyEjqz0Xb8sHHPWl8KzC
dKxM4duBgX8ie0b7UwXm66lDEr/N8K9843C4Vcd6Tx3g5GjcEKVJeL5J2xi2l251
sftZZADLw2JojeVodwJqaEE+VVnbJ2vRdDT9gtxDNp4HMb55cfvod4lUuxctEiug
dWyJrLfF5W7bxwkixdr0sVy3GiGn+6Ru1ajEw7f6SPulhXefs4tDBFFsAEXz29NO
NO6jsGtQI6hXo8uRPVMZCoxPE8A6zHsN3O0rVt/r6+lQqy+wVda37DJpWBQu4GHK
HWK3kz8xUI5F+PtLsZWVqXz9/vQmsBdyuzYP1vHtxAJZIZp1ImoXI6Afcb3q48un
PXcxg0wHjDkgRHRf2b53uLqeMfCCY8xKZ69VyE86YJg8VoyrrobN+39FS7NKmIUG
jYFejNaj8H4SNOHdpt/ATDVmMzS9+LO5FexjXWuC8qYMj3t3XJsbtF1clCyjgjNf
2/LhqQJgqSisvUYUfbhFpOI1YM1KH6728YtdGXORHMS3qoDX1JE69h7lWfnHcaLW
rNagb7sBwm+OvaqBZk2yPgFWtV2Jfm+B9/znFT/ZvQ6+f7/4BQEo36gyCFJHWo2y
fJBP4rPyixBZuPmE8lNWB03ADG+ljIdoEmkRI/ORMBKZ8J8gaGVZQqn/paZsDhag
/RPlZ/fptn30WEHQyBZTiA/JhiXU4wQhaeDBI7ZzuspJ4ZUPtq5yeqDIWmLSofva
71/VnKZI8gU5rE/uO5MXDqBOfhHKrmWfaAKHLg4e1LxpPkuq9VqiAm2tXLJYUYNI
lzg7n0N4mK9Cg5rF6WXIUzXzOC2A7G7fKpD4o9fsJHAQud2w4k5rUpLA3URSH/f7
66OusIjryigFsmjOCu39IwmoY8c3Pxd66sGOh+PCvI0o/i9G+G4bCUukYG5/Swvn
SzfeKy/QvMGQjrmTIzfRikcSPHvsmyb+XEWJDT2TpwJYo0QKkW/egnNg8AuSz1Sg
pWgxCRtfrkrsopdYMp05iuRPrRVBr/zTwazIf5nF4JJoAP8bpclcB0zIQ7fsKBZd
1pywzJXdNY/Mar/zDsvbjF6qSyu3rFzWlWxgAHOiMHr/NNPn7yGTpLGVXTu5uBbt
onvBxmYAuQf9M1u+BuhQfALAx3qj4nTjuPLTMIn4+o187dw7C8ICZLuyYxRfGlWn
oBBBMrOQMaF1b5Egc4Rprge17JMoxKkxGn0EamqI3XbmqxZD3bfG2Z5BhEXYETH7
57TQ6bYKB674+OcYS2kok3ACMbVslqo9wc9BbgJ2rpYvRh5tgJaFIPwm4w3MGDBz
fTc/tj5UufAr6tpU833vF7g589c//cZUh4SNUgrBGNOFyDEbP8+jdhhEt+fUUfUw
fkvXr0t1UdzKDSqTpkWKA512IqyM0OAwejA4oS55cHY3fOCrnSkQp7Ac3uS9m6EB
djSgwdmpmXXRuLAPmICiJCfO5HvUxQr3ckg+L2Y2/SCIlnW3d9eSU20Rwq2Nl4T/
RZ7NJvRcHmKsKYJ3b9THXvKh6ncvR1PRz0kthmPE9BJl3+IjIctqadQEj6giZleG
LtIAav9SJ7OxNfhzU03D5roQM0QBbvO+LCRl1dPPswlKCM5VEhaYxCPOKXfSpuq7
n3eKtiDg+Hj5UIjk8J6xJqCe/zP/y5NOKHdsbicmjNN75+po92ZY0NE1ErdvniS1
TYCXTJsjBcwODGBGkOp49hqYvEwGm410cjJSM3KLGRs1nQgXynKJjmGN1MFOCwCF
lwrm3KlMRVx0dXyP8/L8n7LNnz/y8tCotFZKWmUHF1PIuVIKd5Qxln4vrcgGl1Tb
O3kM2wPEOPYB875fwZQDgZ2v893684k7eg+vr2u6aOZhmr+wbq4CkDgce9P8m6iM
czGJOxzUbQ7gh2mO9rmDeEvMs9l+9m6BbdVBhO7G7VxcnDmln9FbURZim7iUhoo2
UIDHntz8oDRHhQVMo44FDgLm+uq+cERjwiHatFjef49N0zifESSq8orhhG+MgG15
VEix/bypYPDAbeZWFyEwVXzqj114x8hAjkFsOzdMmw8qR+tJWMQvj4R7upCmDbGl
3jyNot8B04U/QB5nynt0ocTddcCxk4J1blsFeRS0miyZJr7q2DuEwTtpFqyMXi5i
cCxmUaCrREFbIq1zxB7fZbuzV9u+/18oTTeGexX51k4pAqFLUqqskHLWu1aWZXpz
IV4lnDJ3w8K4nwscexCMazcaR51QnNYgSHx9OvC2E7WnGYiJdFvvFVCd7N9wPe9g
ceXZ2xOhHOb78F238hm9DQarLHSwmf3G9T0QniB/uGiyBE+zHmbfnQ/A5Tj2QDQ0
ZBEThtYr8nSvmLDR3xm0I/mlqqL6Zef2wLY/EcNPKHC5oHGg2sSmCwoLeVloiKv/
JWWSeL3AOiLp5pRceWeD8ANz/mFFNouVQFEmpPtm+rIqr0q9gTeZokdQenacyuqy
6fEFpUOAJKU3lIKBZM+2ajeKCRobpuVPPNob3mb/2knq2DajnSb2yi63JFAbJM3U
2dCVNLLYv/yb63zcxVE5BQzrMeQQzWD/iWr7HbF7VlPoXCt+EKixek7E8tK0FasL
Phdpzk2DsVCJaMZIcta53s5MOyoFFmPiOI2iRmx0yNNc3U2DaNS/QHpWL6SUWJMr
c+MJ87apx+GJFra06KlDGDF25XTN6yhEACF9+btQSYhwj/kJsYBnSFD+bN2cWOT/
KE6avL3VNY4zXfTLKWuykQ1spIBR2Ciu+2QXpI/BJntB8H6nvSI+ftEycS7p3/24
wVvML8FwH24phZnGMJIEKe6VGI6tN5WtPSK/Py6m2VXW0zhffQ99VUhNNjsmd9KV
we88rVSdd/vSbC4dKeQj2kg+HcDxdGNvqMXYY1DtWkPG9cjm8agjXRDf+ZrBkODE
M1U4YTjEJSUaaDDlTdr98tpYm0o9PXToD9r8HPhKCTF8tvjeezn38pB733IQOQ8T
cYutSD9ycyX4xrKEb9eSfZsCvjZhdMf2L3I4B2N9EmqLj0He+hl/Y1ibrgnAh/cs
MMMRgLqAmB2vjpsR8o8+qaOe0r87X/OMcwAR8tF4VWhhmd8V4NZGiOBgg+H/oj3R
xRxb4K1qeivDve+7X++HQkaHs5z8BmSx9pY+bu3mOLeJVemUhx24kN8UG1GGGxBt
fBUS1NklEzBSdyDIkFEyE1hKaBLsjInY6xuiesnp1kKqa1RtcH/bvrL4wJHlaz6d
pi2ZfSeEcKf46w0H6jSBctYr/rEf/WT0UjqT8srIj1NcYly0UJVFJdN0H95I9xQ3
oki1D/9CgEEjYf1ptg0kftYg86QKNj1XkB62ErkF7Nw0lrqEMnqt6T7GFoS+/cT2
YggSbeCsXKf7qnnp4l9m2xBpjtcwQ4X/YnVApLykgyiMMXsntg1gY1Svkvdiknng
RbooDef9wpT94Mmhnsa5EugpUEckKEmDqS9li6ySLIKg6vx8CZkdNRu2G3WKUeI4
G2OgHPzO+HHNqY2oXSvg5IDbeJuVOHqSDRpe0oP4qmmKf6sJ+8W1GH9wHYhkfawJ
MyH0OteE1pYlDkxHqIKK+u2qP+BgYPuaHrRJTLa3n4usG5W73z1cEExe9dIMz6GT
k5oy3afz2101svhir3QSrl7mRTl29+nZ1wNDkQfZIPAiCHjBTXR/mpTV23RDnJCA
MQqPyqKQueeLRNPPmsWsrof+LtSiWUtKiHPhQI2LGkuky9lRogoYiZg9LuJZrv3O
A2i3SGFxykT/QAPQUP7rsCGBxugXnj1z4LwiWShVZhuKbmeJaH+pu5hWQ7zbmNwf
D+UV46DHMtFCEXrPh45yqYXyIJoApnuxbeg9CJ0um+eje8VhoU2s+cxc+J5OuICS
NsQLK2O6PFoOBAESGz1ybC/BWv1IrxZeOPqCMSm1hg0jC9nvkt7Wb1AtqhL6VbHy
V1BSYS1WtftWyIqG1XJXEdpmCH/pQPpda3Ttgqykfmp3hMKWUQtoMIFfLm1yAcDl
F6Nr1em/JTHPLs1lM1A2PuHVY+gKvysAP1w6F9fUtQ07rApC40gCDpE6U7jJf9ne
fYY6dFn6pmOMrnsaKMuiBPEjuZSftNdOUWWfHOarMUZZdm4LNknxREvkqUkzfPA6
gYsRYP9kFD0qBXTSKfExrXYRTs35dkLZibh1982IrgU9Mf3OHJ748R94mVOcEgD1
L/ue9WTjFsOoin/FhzJKGaXRYbKP4GuZ+IssuUA90wKe8XvWRrISa87gSsqZQm4y
41RzK3HvNKLlGs15B+3dPIYFwWmVUMkOWSgvcDLPZPA8loV1xF5Bhs/8ggzuiWV+
ILmdZQwgCZD/ivYVt76vWQFnRZnsml+NcgOHVz8Xz/AL7kKtOM+/wFGU6xJp5AMi
yV40QxVDKre5zGrCRPGKDLAKCKsT+QZ7NzeY7o6XbCLQ1L0GnaU1eg3EkH0MTKPj
mhkjfWSHamErNdzXMU+4fK8k1XeyXgv2j8ZBewvCJWMyz3lM2iHO+7IhS9Gw8Uje
kcne1xYINuwA0VWYewH6SGL1tSgeNQbWhvlLyGvkbppNiTqNp8VZj2/4xrN5OE1y
K0Boj2XumY9ZJ2jbtPzeq1z4Kej3l+ppAPMIXBWAZ+dQQ3F4BS/Rw+FkDSeLSVyd
4TmTbb157TndiJNQnH4eECGEUJRYwYSPT+KivwHl6YEteYArte//EPtJOobPsuDD
0uMvA08gvNHmVr9JYBCc+apEUEDwxOsycfVsvy57/+Tg9HvnsWOhJGR8aK0IgDsK
d4X3Ywj4l8pqeFjmZFbNqV7V4+TPhoYAiUe0v2XreZey09BGHVTX1s0iz6ZT0AQf
roxFCnXm1TxtvIs21sUTV8ScTG8SzaPDB7eOjVIOzk2vTXJXVDeOujK96LltojQJ
2eIJRjzcT9PX7PgtQz7LJfwzg6hlEGcljVyKiaW3yToeJI0OlcBFivVWZtbiAbt9
JS/vp1Pc3OWR17wLTNHQXOehqAFzTo1AHiqXuMdLIq3GFgoBbjNnd7hjLxv4BJ16
m1004PxLmneZpjsJJuoRi9BYjjjFJzLDfB1nmV1day2Krgw1Am9mW1uZ6oLOwtAE
HyA17Q2C8iC4jVLqI+Jd/QYOwZKbVJQKG40Bt23R9J9oXZdDSiw0NxJSf12tVk1j
sRmxkjnhfp0Is0hFfpUuROWYdkwVSZbl7sTyupvikF+0MGgl5JPEYZp7SQ7XOitW
cCdW1l0SMnGNrAbjbV7Bolx9nj4dJ7NbF/ez+A86RXU3FdBTarPrfJV9ZKd7I7Lw
/zuzB8fY3pE9ctt7aweh4yQKvUeo0XDFa606bDJoXC0PSauma/oBawq7Gn+bHEFX
9nC40lBn6gRDs/iVhiJutjhmZQxygCinO9PBsCmy6DgNRkH5ZIKeAmVSi3NKVrlE
w/rpVKEgruGuOR1tWKCCbS0geSt36fcj4S71GG7Z7Mm7Gu41gmzmg94+jrObJBTO
cibX+miYVFCaB65M3++506CyyOR/RlsqqZpAV6Rd1rLXiWQBPHDwVA68TRf5g3KP
dlc2Mqd5Q2VkDxuVg/FeCWFoJuLbmdxC6IbwR3EsSylsgPXCmDW2kW6TKLOPtbLm
t1pFHTnBbYBTPo4janTGl9xVIN9y39ctcI7yXUIoi8TEC2xRGxWSMkoXRPSylF3r
mbKcCgTvi8AuyvL2agxLoXqWJc3qCxYFby7YrSzoly0j4vgslK/0It0VkbK4EXcG
k8QBCjL2o5yHW9ia+BYo+O8BZaRzDSzPfw6b0a/A12fNq47UHtGinxUKDTGL7kwx
1zcSIeDZyRHUp87jOWz2inSZ0OLM9/V/4Jl0dfT+weZ69rif5dExJ2CwvTpf4WFr
RyEyng9qpo7pu1nnNIKsPCl3WEUGMTLldYP6+NBXHvjFK10PaVQ8BJxst9CUhRDf
Y6BbT6bWJIYVb+UkSrmx3BNHU2apd39GOHqk3Ev/167I4x0obVc/y/E59rwqIdVn
O5Hc52qR5o7SvjU6408mKBPnsMwgPOYXRv5PZhsUUrSuDNrRSkfxrijA11Qkzrke
56kVAEkrq/umfjihirU65qQ+VSB3E5BsOr2ERxjRL7LcUlg4Cc+jDB9yHbp8tyaG
3JWSCJljmhlmt8s4z9UZISuzh2b2lGzv7174wo/TtWIvj0IueLOP8C6Bso4DNg2J
B/BqKizue0iFitJlXA97FtKS52dMVoHY6iN5Ddb40DHKRBkidnXqatpj9EbpUAS8
tThC0ABjtq3l0+s4zS/FtE6OYxsRhuB50PLGMOLMFw3hAm6f4mGcxU6QxSitgZ57
oHMu4h21KP1r6g84DKwf+e7Z0KRlVyRntaD3XTmS563WEUrnQ8EJDAVdet5ZxPFr
c8jimZFVRmOWdIHW+oBum0QD9eNq/Fk1OeN8I/wBwx4iqOQMRp+zRlZuO2YBapfd
2SFHxRXqkv+pCtO5bmjTvnxOoDeCfPf+0y7do6IJlUeQdCQ7p1k9cji/BWqOOGGk
0vQGj6a3ohgfPP5TDHVyi3YMWieQ3cn2p+j0/Zq11b4ikzaydml9oDtTmBUdEiNQ
A03sgvOlrR6lw3qX/frM2nGSPUBLByFyjhr4tDOc2FnslOZZ4aYgpA4o392r7g2p
69UVWPJNuHKNWVh2qcJiFQMW77tLZIBdIRiXtTDRqnj6Jg/y82CcNAFtxlctuTM9
37fgmTCzNDrs3rzxzLM62E4VIzGcC4XwiNCSP6MRtkKwybrWDQzeOBzs8PuePcKp
YEj2F8pmvJsmCG7ml8jlRKmNWGTFAK9sY2VQlL300MO/9deKJHTe8NrpOubVXscn
74Yb85BWy68dcHIb1HKDDC9m1V/r7lGBvyvWhD9XvcuCj2B9NYAvvg/yQFFBXai4
SMAaycmj3HokUJV1qOnP2cPIZU1+xdv4GCCwbMayyJXmRrjw2KMQaV4j8DZXIiuU
pqSt2YzE/PIQRn2FbsEGFux4KXI3CQMf4We3AjwkUDVwUZ0OxKMebDJodwahQHTo
r/iCecj+RL9dQRCFVUfXIS27ph3tzztCYVpLl/ZcO7C41plLpqrA1a6YHNzq/Y09
Trve0t7iVBu7pDwp51rgkgeHhQrF0HQLSxbijk9Llr7iADh4C/mauLFaEyBAsgsK
nTJQvh+sF+Bzo8ZuJBCcIqwem2+AIta3PhC1BuAyPKgG+AajbmOSHV0sXVw9gbzs
CwaA5sWxZWddetlUpgowG2K6KRGmZ3r/RaBL6rOqz1aRZvNsJ5diWzYvXXPwTHax
7LmRJyNQZtfAqpkuoguY5lBOagiyS6o5G8Nzn9Srb9FlvnnYRiitV7lfrjpLqf4V
IukUmfZfBsxyLA3CUT3mjxinyZu9t4ygxp6C+qF8ipwvqZmhBuXVbiCN9ErCgpNF
OF9HGgY1/F4EreGhRPWRvnSznFpoMBvwON+doxrtDdPZpanr3Ujy6XEYTBnsfRji
eodGnbmMLVFDDBhTHH96Vi/FDHj5y6KkQk8mo50ZPDn4q/B5V86Svdk6Ij8lk6u3
MYq1Ij0P2q6a2fYpN5ybjCJqUBW+EyMm1wj1wOnJuL4MkdWUnfteq15dCWRfuBkS
jY8BiRmyryIjkJmkx0glk7+/Fk+rMCl0nAVvYd0HLYa+SR5IDsGx07+ug6MkTS5v
2lY6tcUfQ3s7CA+AvHqqVfS56chIDpvuxfbuXU6O8N1XDLBieJi7tLyyms4mE8Sk
C2RiejZMknWhDqcyYSdxTsfmlpsgzxx+EHdhzINpc3yKMuxhvtEDTpPB80EP4AUb
yf9rG2EIrevUpbZwk9rhqZEpDS9eOJ4Ux+0O1la9yT9VlGFHheXwL9Akrk5vYURt
V9jEBN6uSKaxnihIoG8H4RvpA3XVUEdd9IjgXOYwAUttdnZsle8/OtswKVopSgeV
tYThnDxr/c07vsAZeaQRjF1lM/alt+RfvdvBCUYs8dmYp3QpRgtHhfc1PTHUH8NX
QX64MYs3zPv93lbitCFsDj5MUdpoEDyOXKcK/H6moZehMPDeuOtaCynIWp0lM/gz
tPJQHHwgzEP7tWr6+61TObNed2h9rkot579+Ro1JKLr/0GR8yfScnBvF5LkBmU4p
Za6JEao5SfAJpPOGyKT50xGq16vOKqNvGq6XWeFIJOqoJj9Sd/cXEx186r+pJlwq
eUo/Uo+GbUEVotdvKXO+xz5Ntx42R7MdIn8b596hyCN+hVauZAc/MUwy5J7nDX0t
3ooRglSlsuN+TLl7AfFYqkXO6tcQabPhzGdeaWo/HtAeR7uRClTqcj/Zr3ISMedI
FVmuUCiv5h65Mv12tifqME0golgU6vATFTPTBHC2ATbjuxBsyS8d0qhPVR9AjYOD
GUxXyakmBpDwp7PaBnKATl1fA3uvnHPtjyjDmbEzr+FlbuI9ogqox+4orE022ZTI
Wxb6Bsd4rHNBu1i32nqafBZSA6jsqxjXIzRS8y/3Omk2+87L6QBcEM+kyx3zUO2m
jV37OEFlm3DN9lKH75kHWlxuAoLnkLo1hUPq+MYTxoCksIHr8BN78Gffe9JW6je/
wOJzQ18qcDcVSVXc1vtgNSkA7xXCJjzrdxuYJzurFjMVCgdm2y0BMG58NrVFDO9S
iSR+6lKTHb75FLBGUVb3xDE0lb6mARVe/dZCSgAMmD8/UWp4PWEB7BASu3Is8L9o
mmTpuz9fo/kz1WzXY9VGm9h9oREFKRZHC4xnIFWe/RQrO0W1IYgoVdodE43BO7jU
QtHtZkqxoAB7SObIgrpmnCty694NsbFexfN3H3KeA0l/uumtDDTQzYEmikD3ZKhp
5rhN3n90UtT4c+yYnAgLmrkMenMdYq73e3n2o3D5+VKwadm2AjwRv0VrarvH5yu9
fhQarR8HJ5ve5IvrCmda913YtutYVduXciEdcba0n6RL7RGsKKQC6L2w06/IMDYi
p2KtjWpYJfCHD7BIaIUjjRjoUmUSgSQPRjW/eJ2ua6X5XQoVNRTbArW2yeQFqycL
MTU3dus66UuwXHc4P3ha9onc9UVj46u1hEdRerj5Pj3FQJxxkGBXZmACMnPp2F2c
KeiTby4LVdivmsGvs0zKzzpPTlu20HcF8cTN8/0y8yfLn91uMOTuYSaqxIB47V7x
Jam4iTCwE339A2dENDXuiIksmQwIyMQ8avsn4njqJLaYLyajqSrTQlqXqo2PibxH
wN9QKiCgSciLjUSC8F9sHjSOiMf4jGylwVV7asR5lWFs4hZbhjGxMmALf4Unvc/A
AzBw2CiGupxxtJ9/0q5abrEnbatLMFOWlXZYNirp11dYahX58UhuVGo5nPOaW8TK
o0G9KGChjXwsUDvGX13v6nU76q+doqLerBR9TMYXAOHvoK1AJle7doPE+dV3Hwr2
ZU5YOpoN0D2hEGKEm/MFLmeu8MUiv4U1n82Gmg2MR5AsScckbQqi4UU+chBSpKGC
4HOU1w8GcBlG1q/lf987bju0AaLClNix1OQrzz0Xe8sjtmFHB1cTL+4cfx9CX6n9
GQZSaHsfxHyUFWBPjWeV+OPgjKZRke1lCMt33OCSgxaMKnzwHPuuU+NEmEGyHKk9
bUalIAOx1gPQ/bCoAbqO8aLZciV5sc71JnmwnJt0Dwl/POmhVyo8klAdg3edZBv9
/lSFjxMlvSZ6I+YLFmuBxVGtTx+PiyC5pwMaxLNog7VwOX+/YC6zUdIHdRFf/8LG
yKfWF4bQTtJN5eidS7rcxMBSav3ykawdgrPcKT9sWBjnA5Nfxpq9CVHlNJmU0yl2
eG8vlzq7iJLSEQLJDJtkYHUMBFYTxPAR/9XRYE56Khg/9fnQHIVre7ITjghPevDH
fcKTMRRLzS+47qeiNYgei43yc/5ju936Lf/Z0K1coNlYMSPCqtIvUSCJLjS2a7Kf
yece64lpIUv0EUMLOVBuSRN+WrMrxr0G4c/StbSPE363IOeakKGGtAt3cIzF8Hh8
RHO4oxQZios2+e2yASCwFzZjmyQRj0aJC2dkTtRe5Rg=
`protect END_PROTECTED
