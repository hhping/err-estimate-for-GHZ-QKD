`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eatuMmk6c+gDaytXY2ekCgV6XxCyWPYyVzTEto4qKuRlRh6iROUuuR1QgYl/RSD3
5Qm9JHx7S35P5/aQq+cPNCsH68/B4qy0OG7VThVC5/lTnBR0vWMrgt9PSAZbZ8ia
YUUfDTFq+k+AWU/qP5lePKhLBGxCM3L4bvgG7s1mk9NSXyS3cafIOBdfCYKT/N5S
fz175LZVz1vffW29P2ap4a74WRkR7+optCUb7S/sdRNT/Md2Ut/KNqGoqQe53hur
KfQNJLbXktflPbVyQ1W30rNQsMdGoNlXZ+9xze4aloVXyHGkapKEsfFabUKJB69F
dVdup+ULdK8/rlkqaSKLsaN1ytgVIyxHgHM9Dz19AvPb9tR7CWqDEiW7SRIlqUnz
smRSIBfdwkesbC/qlT3zk6GcGh5VwOYMGUQI+hyw8ultZ1/LXZbdWzUnTYwbpri1
jC0UgG004YjWgWPNDfakzfqqB7skNXMfgORxbSJBgcRORmfto0RZ1VsV0oNVqlYa
kD13xExe8ruIe0uRRBhs359mXHGjTuC8rnAE7EYs7wfdA8IvQvsGQzv6nnQbre7Z
Pkr3KN+IRwZO9cNi0FlpSYP4EXFJiazRZbfjMc2a3DroKdlDbwbSkgYwxStYUAaQ
durpGcNFEcMigJNcRkYNXY+whwkjMWdwc0kp+LENQLzB8q58WcYPXhIIn3TwRd9O
xjpsy4boL482YIFPYvJwhEXIZXvBLXtuelAGA9+Dgnw08UdSZY8SQ+YYyslKvbAY
JbVYgYHbZ/d2ZEYWw88/YzjsZKTZJ6lBSpPhLJgppBN4KV1qW3I7EN/dhZKWdH/L
L7y2UWEjFzTmCYYmj1jvQ9sN5om5XoPX557C7fvyIOe4IKmjTM8KLmUqPhrDkvc1
HogXYz8xhTojOJOsdVIIjt4xQH9apqenod6PHlJIwCTg1S90oSG3RYIYvuQiq9og
4aZwq40Wd71NldU/44MrEetIL3MO/KN3uT5C2wfs1UklLTEaTxublV10AU7pRZ5A
p+2kSp+RxPWbmxHFXYMi1/kLJtm1E2w1yhD2aRekq+d5uZCmmq+gL+BD7nupOGKy
8ZhE5ztjmPu7Yr+2bcLVhELXqfqzP5vAnZfimYFGnAfrOAG4ROS93gVnpw1EZDPe
7OiGAXNar7ugQq+wMtviOFn/ifc/Ri2kSdhQ2ed8vIVBM80HnXWiqb66wzEBP4Hb
/7QCxnL6OYNP/NidG7UInvYTw+hSj007kFdvCP2UjL0oMY7rfD/OYpTnd7VgjW7q
SXDNwXKmInZ4B8/Utv0KnF5C5rFcGDCIoAAJkhbizoV0AnNSR2dUANGphh/Xwznw
sGY7XcjngGCiBVCdsopYcI/Sf3WpwkPR/Z08qEQEM1JXXvZq3kMirPdjrZ2hdXx5
hj8rg7QcRmlNJ6f/0neephTeYroRrrxMtL5jMR2DpPIJolNu+EnzEvoYwy8HyY0s
JFtTNmhrekcbBFVXPXIySS33fPnClO9bHjO0gMgd77130w6aHDleiCwRW6KmHe5l
4Brya7sur1zBLeJfdQivvhrJ1o8yPkOWbr4z+9vG6WBAAqpJVyGks6kGgyP0YLUW
UEy2F9Kt00zY3OSB7v/gKRevsrgJflyzy8ugiBwZWmT4bZ0ROcj9i+LhxyBmeXaG
wSvjjJg1riQu8mAzp16RMshrMh81JBBGXroV1EV9773sKeTH7amo/jO05d4otp4d
msqZ9Osb9qxmEr3UVp06/wy+qnAo4joJvDJFKKa3O5xew6cy9ukXrlBaD1JK5oWb
K3dUHK186JzOpF8VGXmb62k3R+RhgoChBxuOmW6i6d/9fL652lwPvjrsz+C9h0Yw
CZLksMVbD7axFI4O8TOj6HcKJ6nDWh4q0W+mHXHOUj3j5HzmJ2C3XUlbqTLjCcEg
hc6fVy1g3YIPudJ14XcBsIYCHoWgfyvOQEt0FZbX1HU4ExG7JdJ71CMX9cVRI0aW
FPjsk133h3L5BcUhAX1LNhfVjH3BV7KOweLpK9BP444VacN5q7TTqcRKnL5Opn0G
ofzKcQjwZcHl/8uUJNXNfPfK8cliTXK5H2vcjySPBkr+c/k1Uv59aYow2kQeCY04
ljw3pc8BLOJzmFuawCl6e7qLTWhopyM0Za3krRMtd6bsDRO8YgH2egZrJpmb7dQh
gtiX5vLpKMTdxwkR6cENvflmJVtUqycTADsn9+Z4ir5DdR5dX8vfW8fp6HvWwopD
EwhZK46XWrGKfD2fqH+5EFVvX9cQf5TdCSxClMk6oMLcXTfYzaEpbSGsp3TmHcE6
vhOR/5mO6pcNJE39tDQScmXDgURKrARYHEQSdMuEg05vtFJ6J7AohtyoD/unTNIk
/Co6hPHH3bfKI/78QASn4W11COeHwwm22SHY81GNgkjOhEVRX3YwbKGz8fNF/dyH
gVaIyb1WqbD7zjAF0yXi1/D21iqRUcEO+a0fyIbC5MdwtZv4S1uvQn1FdMOuFmkK
SFOQfS3qESO5+KhiwxDsmCWINSeIDTOMD8Cx2t4+221fn8N0Ojjb1Jj21gyayoC3
jDeY3fH0Jey7keVprxQu7FsF6l23mfTh0X1CJ4GI2Jky9EVMcL2IHChzb0oRyQ/B
YzpEHRJMXeGY+aKekpfsrsR0Newivkmeu94dsCLEVjngPmhb2Lrnv/p6B33pqUAO
uIjcTwPEqgwCMG+MW772vdCJm/IO9i2YhiKYKcb9S9CaZ3JeBYeRUesMMNtqQ3bp
rVwy9TBudA9UkcmxiQtRzfrbSjiRS5USAMIz0Rtxc2hR/lHaZ4Ni/y4n1tu4uTvp
WMc4P7EKx88Pelorj2CPznXjoQjt10jxI7sgfk4sxArumooF9Ym8CrJY1oLtdNAt
NpEowwyeVReNFM93lMnWn597ox1vzuHXA6GGYAov9wz9xy4qKT4vams9HhGIWW0p
T+y+NrmNMPwVW74K8tc5ZA0Y5709ruyyXRjDqQfj6/6NBK+w+BN+SzNuqKXEK1h5
KMG/TDFtWxwMEfxSjb4TwBd8nKgbxG72L1qz7sjSOyp8hegbiI1/aXnQUiPEJLk2
fPmOgmqa2a6kYBDBa4c9dguywVdEUdZMeHYp0nanBxwBUnJ3ZPEXOdTgYR1nrv8b
08CS6VxPFojTggxR9W6Bs/HqSz9r0d/da3VQnRMKe+UxnZZi4g90/G4KBTXkp28N
xx7qNlhsYNyGjt4JkprN2WekT/0d3pNs8wRGkrl7/Eq4IawQiFDMGm+STbnbPmJ3
6/sLlq5WGeqTA0pvASMVpaAowIuHG7JdIAFJuZd4ggj9e5L2+M4VKdxNbIqmxXiB
0c6aCsvTuSHwgC6m4aVUjE74GE8unwNNC5r6j9I9joz74JJMEpP+VCxdvSi2WmcS
4HkwjgHWcLhAOuDrjnZOgEnViss/nNxJZyVFs2zdqLMrBgXrXB/Xn+qoHNXXMWQ3
t3bpaca09rFyEEeeS/dz6CtdiJ0s3DBi8nZk1XsgIP0056Xw8VoOUdvcX1vnA9hq
X0CryDUI7obUmvKcL+Jhj8VkrxAQ/i3DnzOotrnAVQRUjQGD5ttGsPecElCBeTYp
egUzZT8ic+cYTuWJUXQLTbqC6zB3gW/i2Rk1ys0XE+mDnOlIalpEZcGtixqwwPz6
ADSB4sJP4e7r02V6ZteTXbTS/4vTZfUcboyhlWi7fzLH+ScndoHwb63GU2jB5V53
SafDMEPQt/PH7n+uUF+F3KDNYU+75qUsbYumGaSZrWZxRbpgijpTxwifuDtVd/jb
BAuPtxYT8t8GFyhTW9T/XBYihQwCStIRxMiGFLoylTsKyQfzgqtvPprhcpEudqKG
k32bBut3h5NUE+UjLO3MGnp07nsLfsJ6n/hmUAbfEmvrd57Zp+2C1UhVTbDogphQ
scc+Lo7V3Z44TsUBjTzzKRdqdapABo8P8zSUrMuVYBKpy/vIPbUbuj8ry6hI7F5e
fZrJjs1y/K8S/gO37Sm/DKQ5TG/dsKsBlpTr7FUu3Lzlb2eAhrob/UX7lyMRLJ4L
QT21M/UWgFo20/zQinG/dpBBdDsd9q6+wVGAZ/7h3fAEC+x+bOGRrsp+C0A1ONy9
U7at55tIPl1/wIJ88A6eKQQlC02vm33NSQssZYqLCeZ8wCXFcJlHyWw41NIN1BEe
nF72GSruw8RLDdxBWmFXAwe52UVqUHHAs5yz52Gd871oLqZYpo34WCFGRjEHxMPu
XZVyRaLnllM+693cazswESHshBcjtDj54ol18dgf9w/8H3pWa9mjGYw8Q0RjRxxY
X68U8ab5XTSm5K97IcxHXY8L7nv7fzpyAHalPzch4IPvE0HcLvH24X7HbFVRq7Qc
kb0HwjfmDvZwSHbiyFiS6W1lWoxF0hfC/OecWkOMolBC3j7qyNKOlIudz732OAT7
8PzM6v5tr7b88KOJWPMJRiSbQluzP/lnSvsGqmmB0FwAhNNPQw9T/Ulin0TESXFK
a8hPPTFPgP4RKdsPM8fXb8WfemmmWUEElaLK1Z3GajL75znDV5O0BwV4ax/aaUBd
p9HhmG3U7qDWRS3CVVZHFPe+Re3vs9PdPNLDX/jVG90AopSms/N7tZ2owXsgEltM
Di+YSlpepnHQZvYDrqeTr1pMTcYsj09Dt6P+yb07AKwT8EPZz0gJQoHrY/9j/g5S
CZ9EvD6Ou9mx0MHjU0UTDUdE0nwDL35xalSdAzePArwyn+lYbfvIjE1lpW+7nF3u
0trNvuf8DiqEEBjU+aBQJGSP4TFMp1WE+DZ3CB4bntTooP4kxQRWJAkAKr0QTYL1
Uoc/oLQKTmKEu1Y6i6YcAdSv5T9P503Hs7HlZ4UkYDaO1vfwPjzp8GuievLnH7LR
b9Nma94xweYWP2bOragbQbXvLExXG7VAfza0NbFGYdF+ftJNopqjHGRis5TLsg0w
IXM1ImRgbE1m7WRaDeryk3MT+PQ5RhcG5NSoPDNA2tRoNjoU7MsEpCb+JyZf9pKS
25S/wa2U57+vHKE49/PWn8F8r6bxIKk1qouh02mhYHs4IvreU7GwnW5Rsl7sL1D3
BOVfCxxlQ/3n74bDlXwm2Qz98fh+OYerPBInf/X2FjkQ0u7uBZgnjc4tMyvlqW8u
y32R3QTfOoYvApMfHDd7XpKRLqjAH3di99OmzgoFqF/ICIznPBtrQasxINGO27xD
TLZCZFyECwSj1PHMtcnnDkIQu+YYTCR2HrXKmwxvqJxn8JG1l2Ji/QEG7vBmCx/L
oitQMfoE9lwU5i9XfEw4pPGA0PAqafUf0NDCRu6B49CjDlf7Xb11swcedKUYySC/
zYuu8TNItylhXt16ip8rBTAlhaxam1F9iB8YQj7ofbNvUBoCEOWRxNVXZ1+wUAzo
UdZo3zFAWA0MSwLQBUyXD2dlReXn9EwHILeuHTMec0j3JThZf8CoNd/7v0Zy4qDO
F083349+eSLmUJLwW3djd0/M1lmX9cN2OOBVVK8KUdjU0uvmzXaBqwQWJUiKFUnG
a8/Xl4XZ55ARJIc2BnOY6gVe1UWllbSPSN9uJz2ZfhrNhDNlDSft7PXHErXrJM0H
dTW6mfGXdyPm34k3Q6wXVls7VZ+mkNGWl0/SX/FaKI5I8yyRSoIR2KpK6l/XPiBW
CPtGBBF0upaZWZZpe4tpwcBk4cJ0d2rikxEXJGEuPIKeOqOa0MuwLeGB6ZhZ53TO
NY1+5JUzS1NxJ7uCyaboDdBoPeL7s3u0klSpWasE6igbVn5lcnfPtaFQzFRPidM9
uewbzmQ5lBE858rqxHGVFTRBqTQDbArMw3otdKkZFDLB7BzWjzZSgnKYiebFd1C1
+njBQBovArjMLtchydo4bzb8b5fs7vZ4uv0rCSwdbZenJ98DWF/wnIIdeTvuQoIZ
3SjuZ6q/NhyfYw6E1nghdrv7AJCTcWyahEYYkQfIzGNVCcDxAd4xMwP3zZBoWRGG
eIxAfy8l7x0XJyf3tXrcR/x9q27TlORycZ7mH921TpXlr3ZQCDQvmfC+fVqbG6Dq
yRHt0++7U2lwuCpHpZX0qc98UPFjMEp6+orKqwu1pzioR1YkKNGSjzQtxmfcmY9I
GsLBeDUz4PkGcyvK7vXMKli5DZ8/UG9wRjBlcmkmgRwuNBDtBjKu50vlc+3govfT
AKT2YfNii72LDU+a76fCi/ReQoIhbJ8fp8f1DYdfpteZapdXU8TaTbUVp7/pcn+5
NzKC8gcNE1gSiXBCQahPHO8mxjH45eDbrYz6nZWpIT6XKU/TDbennZhUlfHPHv4m
D0dBlB7kv1SKO6+r/4cJ2cNfxWfMcLZ8Wgv6rGscHnXH1jck4/AqfISCDhqjLvD3
1sljJ6fm4ZQ6YAyH40s2zaKgnnuAHix+BAiHRbKympBkd8ENyrfXRedjiKpEDblR
jVBCc79lpWG9fZQOIVzuTjy+Sdx1jY1d6C/m9oXPFrUU42cxqg8pJY9NSrg0jg8+
ZMkN+w0vxHu7ZEDOr7Uz2KqVjw4DsQ8xZ7+z71c8t2fAJIz018azWcIUu99hSzpm
dUmapkG12D9mr4ZXAtKhAoA3PIcA7lqfgbP/gtoKnabhRCCln7USarWn2n4scCBD
V1U5flob91DE+Ll8lVBbcHDoUIrcw5UOyyyjnAV+gprCqAuJWmIPloiBS4V+e3Wq
CAnu9Ng+4g/5/b/ZpcuokdO9kQ3OuCo4k7QxCmy1jCW/hU3Ez9QkhX+Qiy6tyvhU
lOdK1838RaX2fEiPfeYDNlxPUmu+j+fQJpnEZx1ESCsFdBbWyKB74FS3qWdgpISh
r+5vBxm9Jvp2pk+lmBocqrk9kyosvlkTg025c8O5IELXJ6wTa67eW7OyGYoeVo6H
wUQ5rydh6WHoRqBCfE3KHECQtDPKdVgXTSxD4T5WnnhxbVN/aO12c4BnKeCCVgrb
T53fV7ojkLFgebPPiwhEnxn3jFi2OCsFiS++W5CA2Yo4FxcMwQljogh0Y4wwsuPW
j59chjvT/jzXm7/igDB/ihlfUsB6iUFzD+YI/9fOgE7fB/yyCPGgZB3VKV2ftsWb
WjZrYKh5jhQguvV//V24UZXZ5PYRkK3jxpl7oJF6+0EjGfZddR6Mv32WgFWHh4Dj
NK6QEbGtyJrdWejYZy3j/Z+uWNRuZUSAyYmKTjfKqPAlljEFvKvxPRMARg8aX7kz
IX4xZ6w8tw/DyStyAFkzAa87GhNxWCZM9j4uH16Y9W6tPUJzCr6DTEBQKr8s+W1i
s3G9WrwlO78Zod2BQfshSiRQ5YlHESspP7PCcJvqKrJDeTOGFJ7zL0bjHixz94gP
2+qxTMnVh4hhkWeOp+hVZhbYeczqJ2WuQIhfSdjn2plGI+HJCpfdLjX+/Lt/x9OW
TTxPEGWoBYa/XAxPhFKCiqKXvMMd4A2miQM+92Xu9UvS+FAjAzuuSRnxxTa/Wogu
KHLXluS64W50+/0dH4aharCd987inGzrA694D4dsROiP+caTau7uaTmx6l6B86ib
8pSRdHgdsHR6T8+W9VOAoO2DoCa1PA7tS1titaxHav9HDxxknTgG0j4Y/MdCltH0
hIhwUN9qv5L/3M2K+gEbYGSiX9f7XK6J5BnQazrmYlGGf7LQyDnBEKnOgFrS+slZ
c4CGvXNlO5j0Rof0RrBtwQiTgV2ttjZ6WO70rbaGARJapt73cYsbppBr9iOPwkFo
BPTpfPTXYhqwJhe2YrPINThsVGeXFYNWwkemgpxVEXQS+cMNBK84gr9ZOsIGTWor
juTjsPU/rIZz+RJYr4n4kItKL1iedhKruLY5T/zpL2CeXIVAWpbcKB4G33MyRaim
jgZ5izSKdl48G/SqcKWBOHjlhwxcuVsRpTN3oeZUmHOgJjWL+JlrPVWNahEGQhqA
7m+FFGpAU2frLilnRNwRF3GjFntUWQ0TjXo42FzPnO4VOxw0klU9au8bXQ8tSFay
7tv6S4o0/6azTx2w57CU8FrdbEwDXL5n+rlliBYEKtXtikddJDr6Ybuw/PIZaI4b
N2N0RM91nKs+O73fJfgYgecQf2qtv4SUIm3yDuxQcZk4mzxdMYEd5u5iXEJdQDEf
JveUsgj92ecoX4UmUluUc2FpTLH6wf4ehmVsX/4X6zZeT6+mB1oVvyfv0hCih+O/
9Jq9f1JDPTlqPq36pjJnVRrrTOUuEVo2oyeBtxNRmZp4HJtJCif8HZAhFaYkkbQp
CRZfBE21wRVRyOqm4a45/hCnP0L0nLTT27oJcPDNckxds1q4mjXE2xNgAugArfdO
WuJFYCPsIeyeBGs8aROglC+a6zbDo3qtiaEu6GCyxpHm4Yt+LcvyiAhuZ1nZlnT/
YrhpVWUbBZ+zt5ZIBzy7hNhBhXMoFEl30QN8uueM71oSbeFAc0bkrHLe93gYhfOQ
tpVhH1Z/xnPUbap0TKWRQJMntTQsUeOUXK8y+RM1o76d31KyNci7v1c9F7ZItKVC
zM+eLfCRc1SQBfQO6UrbCrPJNJKOfMvw4te7TTvXL1OZtll8W4EzUKfmBMJrLRUT
c859bSI0Z20zZrupifVHN6NoFYavQ3oETkArZqlo5VW4QpL++jgut14NY0hTBjiS
4zpwoSKc31s7yF0vBBDtDh/dgx6gUG+4ARFmeZHr/Mdg99HrV9KoN9T72v4wTr8t
68BQfQ/9c/zidyQTquWHTCupdtTByg2Nia4GWCfcbQy04Q49aHpStSQm9RJyc5Ll
xZ/olLBG+4mrco2Xc6BRrNp2uLHMzoDrfjNdewsGct5wlDaoUyz2SfSt0iKJv5vR
C5QTubZGnYpMa/RpAl0NEK8v7vbRAB1q2v6LsVqE5dhaGK0uDQq5XxX4mJT8BUbu
g6ChMah+1cG+RtMNhMa3ZsQX4lo4044rNt+CnbmEF9lA6zOKnw5797OETFc6t83B
TKeyTRKCKafUysSSY16MQcmCiYEccvEe9rBH3rZBd4eCB3Edrj2WjPmjI8icIgFA
SomISQw6PtqQUhIIcBQJBiUxm3ziDwe2wW8lyMLK1E3RcjBgVVofaA2IsHB1fpfN
RaF0CQkZqehP2QiR3tVSvj5yINUHyhCrQVddgRIpzYeUB1AbK6KwHD9rJ+UYxCQJ
LwxBsXBwShGe7EMkLkjgffqxd7tpTcO6G3W7MHx510BGHQV2/OGU4oqViQAxJEXc
eE+JwoJrv8rknAOarUZwqIzy1F2onivZeLRnzGBDlxpK71/EQKgJWIMamWYyxMHv
RUZ/SjdbAbScBktsrp69QryyDMxaI1TccpaOCWX63FxjXxwMWttPnCA9oHzPYlFG
lOgdeoVBwE58sOhKMva9vXSk1qQTUi37mVk+b7mhlb3kuf/XUykRa1IQDTEwCbe3
9WddY4ZilXqt47kBEQ7n0b2xP0zMQ3hoam9n1DPdHj0wwlZNqq3UiB2XyLCkQz6u
9EsWkLEOYnWWixSkUk1s/69WnUyYRhHfi3ea+PYNrTsw622HplizArRUc3Gmb9Em
aA0zAEr5kSUZvG9ayfzphJBYuRUaS9rPvtXC1oJdb7NdXM0ioL76WJ+np7qidrd1
Gt1cQb8JKV0z+iRL/Zh4YXb4PkZa9sOIQiDm4tBKEafHiCZnYtf6SDoLPVTjzw1Q
TFhKOyp8nGD6lKoZ89jypf0tbPhquqT68rLHxK/9o3Xk/xcH0DAX2dun/9qn0T4J
odBTLn6AYZ0dCPmiCleu3sHVR1ZDNnV+4gAOf+XOJtINErXIZRg2Am7oToq8iFlL
A6p+lIpAxYaj1F0MyODaem75bLPy5WxAGfcjk2pNKEjWHBUwUe+gcYFEIGLXNS4c
6oL0zz9yaJEEHmqbSzaMnO0NINJPG0jd/hDAFSiw6GhAaba81rvEPoi1a9zk/eGV
aPeoMH9DWowh8r+Ikq7w8Fbe83i8pObL7TL/Zj32MQz+HZpL+heeTWgJR/B19mLs
lStg502VVKP+YLb93g9vVOTlPz8wacS+9Ut/R28TQ9yRYPHcSThPY6TXXxxsctCk
xMz2FP2jzciSg1dIfl3BtKsiEe1SVBi4JUFlTKUd7+D/5YkuKkr2HMxI6a7p8OYT
8Mj3mAeS5+UVuIHJpka11hRi1rP7z36rdBZ964FZl1r7AnXa5vMLBvll+mFrKY+l
to2J8eKFKxBe5rRut167tvwIj43k5uK3FJrVzjO3kszWwx//D7JoMYzymBBhYAoc
8TuQhRf+IzkMeB2ntoAt9CqflIYfsZCmK9KDAKMdIBioELwlL9vmPi23wFOpsRGY
yVVEBsIlVonNJFgE0+9eT/tzE7OXLj3OSiyIkHNoOCU42wPYP6zsHRdbCGCjPSWc
LZel74pJgyYYHLXnaSDQj+8kTpJHFevj37gdlUMTIWAEir1p6Hs9tXvN1Ja7uK+r
JefEB67Xk3j6Oa9nOJtMpkfQ9LP9gumUErHudAge2QgZV8P8dKjNVEOil/3yX7Rs
tKC5l3jaHW4abAaC9DnLNNZn5ZnTg8/ARKeEwOPOzVdoZ6E1mnMpV2KawD4nE9e/
wMcLQSHum6lvU6pmkLfCD/EI5KltmcqNJr30nwrgsv2enjZyX7NCYi+pPq1i8pij
vvQvqXZXPikPZLXxwVCNun4Pb4Eq09/olmcgqLOgba9wb5i6/H/Dv38rpkS9tnLl
lx1iJ86cpPUW+aoD+xRRqR8Zrp0pTA0aUOVDviVGzqRFsEpsRQ7NjOj1nmSj8sKM
iPtKeyF8PHZ8SwpTonlWuFBtoOqd/y/e67HR0/kPgAQJDoCKzr7zf9JKzLOmMCoN
83klV28wSrQVc0Zrayfud7A0HFfRCzCDCE8BTz9I9YEyfi9yJc0ty8TEeepyDpCy
2ooAZPlKqgFr821BJuc19E0eJCwKkjeIVNLXd6ObyT0QuIOfTrYc2NyajubWsCVD
m6WDEhL3M0Q6OWZuNaR2eJwbi5KhZESl1tCFbgYa17p+QfW6CbKUgSiJ+Q5q5FSX
WegVofPjXPvhkRMWvGLqjCWqKhceIAvIit0Vt8pS7C5a6yXK+s6SxlH8hH5NbfdM
9k3yB9oVgb5gOAH4F+Zc//Pr9wzXMcDgSXiMPOd69UBOA2BP0rN9uLCnxsP1LZ4+
4t8BTsd46LzO+VKHOysHdKISduU3k+kbCfZ/Y5JvjN1Q6O5EtYb6TRVfXxnl+idp
pOZNHTO5O+TeEjLxCDa8/U/SvHMMZLBpgs2a0isQcuZ6piXrbMErd6A4WrGBnBd3
ZSG320wmxwp3sb/5qtNftWsqXwi7PKH6LGtoC2JO5wD5EaIAyHEls0Q73daH3kus
IqkqyIiE0XdhonYpB81poOYDgWZyXu31C5h7veOxCrwd3tNEasVdwXHDEA96ewIO
`protect END_PROTECTED
