`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WSV+mJ1P0uEZQT7Vq9QmTQpwc0bHKpPDAn/PA9YPlF7EVtdJi8oVYRIowbS+9SN8
e26c5yIPBXGkDL3ANHRQafEKEXZ+oiChLqbyJVFcSwIwLoeqbi1r5ywLDBjL6VxR
VE6+QeK0xtNPpoyv8KQHOYh+337aIQ8AasJi4i3RIG8Ebz5VISr/7DUzkaZeyIBZ
IgucHJj49IlimY/DtmY5QiQvCuamJ67uCQO7b1Sk+lRURrVJ3GrxjJTlDlJy8+LV
IeS4+ooYhGyUy1oyeuGynaRVeV4lNdm2HuRe3xnTVREEqKQ3i05vEKMaUi/WjTzw
RxZl3yw1oFBqJtsvcAVLrWZ6eqG8qJ8HQ8CjVyR7L0GdKmDsflUMkBLwwkuctPRZ
NhTV6cSL/tYic5jG88alR4e4w5MTzD65FndikVTxjm00VqS7J4g1do27aQIjQ5bB
AGor+l8pJFOFuUMKBG2XcJHeHyqjFE9kWUNLVEKWYgyG/GCocRe2rYsNqTXXvRBb
qNpzc2JcDfVZrabRDMeJFbOn4KzeUfNPoLyRUpnyhW/eXXFWmv5Tsho9W8DfUaVA
VvNcCZ9+fpxe1dpkJzvOB/XUD8toW2dvWzcttrWBmX8Ot0e3U6BYWtBeT/uHLcUQ
UxoDVlC55zmoCaHnaiOEGyv4qNNYcgNF+Wo+semhON7zBYCrom/0tMiepd8P+KuW
DEcBve7w3Q9nWQdwkBTrInWrndxdor64TCGClqKkZZuI0DBSHLgpwyibPlyG2Yc3
iRRF0l9j1SKG+Sozg3azxvMA7P1b5ycUnQKPxRkMKCXYExcbVLLf3UgGfaxUbgAB
NUIGURjwYCQeJ2/mnGsN66gUJZQGALD/X85PnwTx8BaSu0KMDZMvnWhvlZIlFAUe
oO7VayBygQcfbnYxvJXVA8tnaC3G346uUwdaMgThFXeJQa1txw7TjGawmmpE2m4T
l+b3W3SGIJm1G30LSgUXkylklbXETCapm+/kBOJyDvoM5QsGqSUF07djlALvhdaB
A+lu/1UMfLMtX2T2MsueGmbMOQHbabnPP0iL2NWrV91X77iMrAPq4EG06gDRyPbJ
`protect END_PROTECTED
