`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1BG8iCmGYk67ru/Nd6ZdGu0nfu5g1ZfWxSp/LICDBTSb0KvHnFz7A2/g2gLLE5rm
+wxGPRFGMW9ESxQclC9Qvcz1519IVFPaFBb62tI5HT6N7YBGPUEGxFBoCHXsulkn
cAoHUNTXACI+nYFRyPkJnA0yB8VTm/7EGhvL+idvbBnHfizHhvXyxYmrnFag4QEN
zZK6ri1//ySvVC+/Q+C/is9K1tdGJCNnJFdvnmCbbooY+gcLoqQA14d28bNHVNb1
aBQhXIA4DqrkLyeZyoFBdZXJpT0uFTMWqB1aYGX4ZG6EQSjIs0PbKJ8kz3qngIjg
fbXokWPJ+y3XMsn0exGk+4b2I2VMUoE4EXxVH5tFpBeUonQWY3ZtLnV0Vg3uRyE/
5gQ2mjkVcBz9HPckWrr9BtMuVIPi4WoRFU0JHgwxRVbp7WmKcYbdxL5JXcEMAwEH
L7wPsM/jaLJg+jx14hl3nRSQU+PvVzdo2sJ42n/uhoBuOCJOn88SH84ID3isHBtK
i8AtIRRV/Xf1PPP9CAW96gJNrLw20faJdNMdlNoWt/lM3e4h7RlO7LkhZuGhrNvR
FUw1lUMobxHhBhh7Cf8VWjt0RuW8GPahtn0r6Uuldmi5BBulOvZl+SZ7ZJLLyObu
yKvmaTcPDGHDG5kzVoDHqiL43Dd383oL1zk1lvBYak8=
`protect END_PROTECTED
