`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2FpMn/ipjBDzYaKVhQGDxwGUI6/x8HQNDfszcnhvxRIZgc8CqTVSfgKPvMRN3iRL
97UOPBbM3ZegUk5Xa8TPmv9TkoVbPoWdHTjOrMF89nTDbDUuG65lcQUjjzYMVJn7
2doaurNyJG+QyPYixpC5VPLy8ELWzQfyv4sNjC+LIQ5Wic+fXn9dHnMUbOmR/w+z
9KcVxLpcleO16l6pa8lFJ8Qf4FbfF4sgkd3eBbMHZ8kUQ6odGe0Ox9zxwn65h2kB
O+OwHk4ZOLcxPQf5rNbbIYuMYIXRKkGA2NCcfHx4bV8+sFJE36TuI/3UftAISWyg
Gj5lrCW02vZrPHPEAQQgt9eg2vlxZrDkN3Dq4CFViI4+b1cFxa2tEyv95bLGWhdb
mcIEktx0DXkvZ9ntD/7pR4sb2cXJs6q/GeExArWKNNJaAjO/juwvdwjcYtmguwBJ
vHh1uWkZPiLjeo3SpwVfAv56ecE660AXlI9/mYy7E/JFYgXXB2EFdF64FFY+ho3B
vW98UpFyeXOeeMKRXel0Wwfu3VPVWNxjUARQU4Z+Hnk=
`protect END_PROTECTED
