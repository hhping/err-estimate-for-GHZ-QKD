`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UxvySgf8+xy6hiDxHYg0HCJ286qTPUkmOjGa02qp72pCtl1tkNzvzzaNFFhT7XFV
NNpgBr9DP4ZdwJeOxdDuWZnB6da3u73uSme4YJQymJP/6/uHPHMlGltEAo9V5C0C
AE26Kro3rem3NFJ8ZE3S+yMji0pISaTevxg6+TFCfwFGYwnXy9kk48h93NDiZ6XP
qKGiBtrXHZslx92FBlOGuzrzpq/V5fiicTYtcIVDtLiXRfXCMzGuvJ/oyXlGHglB
wN1fXcMuJsMlIWzgay7OaIQEQZe+5fmITMoS45zIHZ7Bf7eN49Dwd52I0IYmy8Io
O6EpWITpAIgOjd4dtaevmSORrB7YO9bUXSOsZLS/cfyyz3FIflB/Na14hyv9lHaA
zdrg9WQfUl8eXx3+E6oL9L7HmUa11wq+TA2dmlEci8tu4F3LbdMVEwM8/bO2kGuI
f8UIBdYhBzBMDa7RAAhdQqsKPawHbOO5l6Kcu+EeFOFnfjXpAO12cken76GXSA4/
jxaYaGYsz5yAc21CwyvCrOnRKlL2v+qJcCwmLS0wLvDzbKJzln4EuVeAmyV2CUv+
8A3ta5H8pBYYh/cbhqIhFSyWsrC3rdhmB4KiPdgBlwpfGhNCCUgclUSnRT7BLbwv
RKVgt2ccEMwzNCJ9oSEZOch4TG5llXzmwB/12AgbmK2so3impOYO2BgV5AFmYOw4
41Ekn92fxxU23XImxGHUBY41GEW2aYKULVDukyP9OPyQagO+jjrX1dLJ87dprIo3
X+OWh1BD9Tg/tErL4zclUHk8c4ny4h5L9zxyglHNeupk0Zoojub4eXvM4sPdkZ8P
/wH2BgUtYsGbk+ysKbbLjIGHetx9/GlGUNUANb+4/itnSsC4/QIhjUnp4Y07hEsn
5mux3vH6WRyfmz52SiGmS7O5Ovj8Sb3BdRCZEy18vft02Sk60ss/i0BPM5yLGtvU
rtPjUR1FL7wicvb3z+apevS6yZNgCYeSkpcRpPkfB/oBAaMRVYCoZMwcVQ+0sZjx
SNk7jNNZtnWTJkrjOJLec+tELjXnRoVweFphNTKI8jjnxDjyjePPw+G+4TdGLDVO
TZfjt+K7SU+vspAaVdWk4/PNK73VWw+WO9evej840IRWqQSxwuxGfAkME4gpDZVB
xxJMXlghs4aA5g0TIwKpAZtcPReHSYBPk35kdijNRfkRlgnbt6s7+HFM/2KhxbRE
AcfaBSkfwB2M0+nf+Svecz6irKQe/YylhyJ6ud2S3cv/2hCVOdavL91Qhs2ZQ9Y/
7OY3213cABQ8Nufi2Qm+F+rMpn4d/RAsI5ubd3QWuWncQc8A0sG4EN4qE27xA6A0
OndwRLCPo7cUuPgtjr2OtUSCRY+7O5Fs4WSjqDIy/cxOei3mljDEnoykliwtNQJN
gVOgyEph4t+9tXX8wARQGzXolQ7ipJbV4uqzXvz/KO+YbvKPru6RWQOMI5S+k/f+
Po1xBSoDy9hB040GQuoF3lectsdnrjl2KklPWaYL1gWBjy80mrwIC+Pc85hS9esV
OkQYwT1n/shZaCq0Hg+WiZjvnQLjq+PwGvJAJ0P0R+sbX1NPkmotcaX/1ga9VR4a
ySbNOEBbg/TOkSCMeg//hmkB07B62A190qEe6h3ttx5mx5oaZ2j4o3kasy5cCURf
WCYkUTM/JVHxsli/SKDkVsQQK8z5muZ4aIGq+94g5HfcEhIwzmIum30e+agqARWD
wPOys00Ym9BodjFGzcUB6dlq97/yQZrD1FfAzlcEfHChYg6dAoGo0Q9sY+MIExRM
PWZcA/in9C7JQPQtLxTGwy32G0l8Q71EbxjxTIFkGwFrsvRq7HyFGF8vCt7/LYQ4
XzK53dhz3RerLJEvvbFG+ehVJE5ijXtni/IenXaa0Esu6NppF4X7DiRP7v6icJ5B
gK5wryYqV+QCwZBgFDHF/gYmaNTXfWl5BTlDzhRHAiVxHOV2Wf3RNoW8u3EesWK2
sSksxPKlLAE+ruoDCzYHlhyVIWAwQOo1yOG4I9IA01u5xDHtMd7kXp9ow1Bipozz
0nLaVbIQFLr9fxqKFD4uMplVlAtRbWLpvC59LwMdYAb5QXLIBvB/VUDWcmEHHsKu
K0lNRtGl7FUqEQaTq22FZhTVR0ju/QM0+JLXKTBn8zncUF7FchohQdB1k2Hby5tB
JxlIYgLvKY0Jk8Q0NJ8ZnExq68AURlWFtyHppXGUWKRzCLCKYJBP9YHbdaFfBgZ2
CMa+1lRiBA9OImrAAAy4lV0fV6jB9HwwIiwtKft237UTPOvxRfVdal/55u/cm83j
1BucLw7HQsBMWzITC6yq/h7ICjVBwKvXIOoPaLLMmzRmvkG31rSDGQv+GFn/uFml
MTKpUNNZmgxK//8bQVuaf7/LVkMkuHOEpnPuZEkSfzRUfWELMEAxwKE890pWr0tp
q5wtvRr6hHmhF+j81GCBF78GGhnVN3VuH7ZPb1IShvaWYuxe+kibXTVEUENdii55
JlvCjTtHf49JLD3f82eXBNY1GWbwJpwF6DCS2fpO/u3Ckv4eu5r1egRdsddE+64W
`protect END_PROTECTED
