`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4sezDBI131r4ms7Qstxo1bO8X7KzhPZj3WdOR+9wV3Hc1iUJm0YJU5HDLCVeIy2F
yRDDNqKyrjiFVWJIwCGRgFApyHeXuCqnOqyHUqwMKhlpg58PJaOCZBGPRDz26D3f
IhQKJLXDqoHdKspusBk9BUEoAiN76lSQfnvg3WvUsE71rQ9+4E3DzEUIzy8J8s5H
7asRk/H8vxNYm2g7A2Hen60I10HV2JyUojMJcbQ2n8gHYL3Zok05kWOiAHXzJFIw
fD1MmFuj56DQuDVwLbOmGQ==
`protect END_PROTECTED
