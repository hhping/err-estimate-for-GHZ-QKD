`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pK769CRj28s397swx+nUwuwfte1GLYeRkqNNu2Ex+mF4FeqJ81YxvkX8SZv+AxmQ
R58VUjkPwHTCzsSVc3U5eyIz00y81vX06NMljCUvxWZxK8SuZKBeBFZFe6BZlXzX
2nTAwv38rYCxHePwdXFRIXgVyAIqQFLLp59yvucWtzsgtwbZNzPXVwfg39vpQguE
fdB//XG32mvE6WtaGFMXfvFtjoyZ5ZHv4FZ8y3FdJGC9nRx7ex+PmHhOHlXo/HZT
rrSxfr3W0TFR+dDRQKM3cMkhcXhZJ/aScN7z05vTLWMt5n4B4RisszFPTIN6BPkk
nwygyMXyBMZNPyXbk1lu2Ih+/FoYlHFMIqSf3PLBHrvyjknlKRt3lKjSrc3hTtZw
kN/peJREYP2rtuzg0d2ZTU98GJiyiTCCA1KRTZbJjOoZfFXnZGurBGFe2aL4NqRJ
pTrOppNREzAevEQTH2TSsoj9/efmhwP9bJZ5kodSoQcdn+zGOhWcVutVj+FlMPKg
4yXRZH3d7y5f/O8XrvNh8tCsBDO7ZHMhpwafXrk9CMlkr48w00XXbAHhJ/dePQhj
Ep5a/7IlQooD5kvhAl4pRznBL94pkBjt6HWV7sO+OURiOMKZm1OKAJ2Po2V2N+dX
ftmMG2Uld5rJ3MQ4bkz6hFI1IUYurIFKT68YDxWs8Rhz9eHSOrUI4AWWW/+7h5rr
LP9sxNCvIeeEqSspy8+xz0bR9otLSRjiN6p5apPy8a3ixX2r57Y8kfahMbZGb1Vc
o83lm0uSheOuut9Mf3adDsJImIqxh9fx2ZUcGnVFouEGPW4UwJa1gW9SqghMq4sN
XPP+MmkmrW7Mfol+IED1h6NdM+QmBroorFnyWhIlgpUxmg89QcERDZgKuiTUCqFU
7mUf7PMPlvujOQMXYh6XAdQS8nVuWiHc6UrukwoWlVfKZHoMaQWBap4IQMSrsNnm
7XQtWjpWC+aPzsUAsf3+WxHj3yIA5rv0y0Ty8d0oK1gyRtfC4JERWvdc3KSFMIUC
JXn77zNCaDF6jfFXpjJ40n8raf1EZhi9TZT/kcK7dqXlSSDXkRYxnitMDZO5RDY+
0mV/x1wqptCB/j0Kl2aNCWMUgrw9XzZfjN3Jn57+hNNBw79ZsOJMC3AOugVhg7XR
dzSugiDqYYwPA2+pTO36qvGYcewhfvlFzk9ucR/5N08=
`protect END_PROTECTED
