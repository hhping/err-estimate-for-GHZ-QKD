`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9M/bAmkWeJSgaFuWDYfq/SYudi8/r0RS64w8te6B/oAbDvQ14+S64iky50N2EOuB
va/Z95jCH8qFY2xYWPiTinHuYoebn3724tzoBKWyZ+viAsznlvkRU7sLyD2VxUHp
OywMDUJ2Wy9vK/2y7GuXabitKGRREkO4As5SYh907bJ5iWE9SaFL7r8lJT5wQSHN
3sONt6aOpq01Qo1YJ9w3RWDKm1SLu2NQ70Azyyb+HXq8Hc6WZpyzzoaDClo8v1vF
/e+GjPqRa/lS9uNTRbrobXjQhlnJ+qa6iFsSTe3bfj5dEDPEl2Golka/WAFiZ5cl
ifRCgJ1kmHqe+YKZ/Xr+3hWzgFQ/kMHfsX9ACvjYxM6K5oTLmq6S6T8HdQKItFVu
Dds6ucMGnEuSKrjbJxKhaEeqiTV3qp9IBoyCp6wifZEb0Cl/l8w5RdNMKrJUBgYx
MG5oLX1vg8VPhSvHyhoaJNoeCiV2RuSk6zkn0RoXFVA68dFpZtlZtAnKQSo0eAw6
t43gApqlQ0W5dtQtHeXFnqNapx2ZDXwzzQZ75ItGKPPDa4faUOjMRiuLahumC5p/
10Qkpul5er4JWvZmxewkRU6Rv8BsdtS0JoFeKwUKmOdIKN9nUiwJRBHTeE4lySRu
DoL2yzNEflCLfjp5niVZDsY1xJiBDfU9IO1eKGL54xKk3evaBoYoqu3zBsjVr7w7
Xpl8egMOODGA6bHL1pvXw37I3h6zDArCyKeay6Nog+eAKmx0cy22CytAMJCi16AC
gvhXlaMtdO2y+KVTJ/PRXCf+pDRZC+YGfxtO3dav+O45gOZP4rIKvtcg7+7L9/sw
28/z8nlO0kEs2HMFy1iBnQ/wwBUtn3n015jttAskPtaIOe73GnrwAtix52ZNx46m
+xG77ItKpEggqE196GPyp9/MhJ3z+d4VjdLFmpeUEQ88o66UdMFZXNtX3J3w1kUh
YHONcUT40VUxEevTWFHvL2f8cNuO6YZYhm2eXdoEEvfEjGSxyqptISEz43resx5O
a8SM1XgR5kuLGlqBWsJ5YvKM6Agw+3YZ3fPyhJQ6WvRjr+/c6DM8TQ5eobkqXHE1
eZm5gO639bAOi6aEcrKrM9vxTGCLgAHv8Yb/J1dVXWo58S/5q8JnGSX32J/h2HWQ
iVzQD5qACABfBokukroc9xx8GFvqisz1aXZhd/BDD7NF6pzhKHCu8RAz3QMK5qBx
`protect END_PROTECTED
