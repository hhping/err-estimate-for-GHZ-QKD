`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0PCosO9sc88sTY84n5dLBE4N/u2oOt4YiaEkjDdpmGlN+oNGOQuA+5o3zHsybOZ9
LCRVql42Ln6rVYf+rrY/D+gUKiZ+S/a0ZKwT7YIBQsp4od7XQ4AzBKL1YJi0Dv3c
1iWQovQVv79/kW+WQogW5s83GrMvW97kf42lat1IAfL8BdumSKMN5n39K5IC4sgU
lk6IDf0r+oN9xa10CHaUCY2CvEZLQA5ObpwP2POY9NcLVfQS+m0ECAGap7f96itr
lHLuEYjirons0+3872pURIHaKpMN/ne1ekYHhIfKk1m7J38SMQwsNI9bcLS+SKce
eJjA3EK77hquape8ux1ahwtvYYZlXPANGJMF1NStL8j44LM1ZwiDMMOTuF4w+QHU
SMl/BTRjETxK9X05Okn4P6Wr4LF6kcIN5gRcVJhTZF6LEXlHkdLbP1S+LWQkslcE
H+7aLz8EUCR4H62YrvuIsFK+Q5VrOL607CJdDJj2Vaoh7EtPMQes5TIzf1YJqEcQ
UP5DS3klDwUNmOAU68A0JhNs6yWo3cQAgY1hR1E8bDrhSbI7VgeXLqmFPkwh4yPr
lETrhHrSGGRVq63JzvMFBdxAmGNxwwGzZ37L1M22rPgee8UrHeEksGSVlmbsTG+W
BX/i7tAK15/H8V47i6K71TNmEXb9tKNL2U6BzAklcDecHIRkpndVTjiPibg5Go2d
F46j9fuhn6XRtdtLFBcqMgtjclGkxbg0CXoU5edBi1Fk4Nby7//AuqGS5/g3+8Pj
bofTVdgcMkhz0rh3r97URFwtn232XdX5+Kn6F9D532+IBj07RuYXO9RYr8Zvhqul
3Bo01c8JGDGNZStYeqOmpPavY77HdaZWzkCA5/8hGdCAggSBTY+X7tsX2bHXDgiU
57xIDVU792MLwvaBU30Lv3bTO6+N4ex3Yf0ZFXwGnGZKLIhBuHPpgY/337rt35mi
3N/vlZfbbTer4yASxrtaH6VRlIn/yYYHzrdT5ZvmhXZjESPfzhah2MFrWnn4dq4o
xhKxGGqm8EujEXf8Z8tDf+hdlK6inmot6O57ug3+KZNx8kfdCiGvfgwiAcD22big
zc9QjoSAx4ZahzFfFLnNgHUTBopbfbEe46ju3O1+PxY58onn67JoS3m2KycfR4bV
RRl6hakUoPpzCJE4w9Fm7eV9Yn59aUUCC1y+JU7OL225AZaO9qiJRWpQ3LNNWZUG
5TmnvSCc/+2XHdtTdXPStFYEHfTQgkqvRRbJIfX8rQmXFs6I4nHDpA5Aewp+UGng
2/QlMJrlO2P29jx4W7p3ELa0dW9Q5c0yAzBdxFdaQK3PYgGAjpR9oQ5axiYphjL1
uoCmfuOs3wlIstWxcU+6RI5n9ZNGMNBbWUUZOxC2vYwvGun4I34wGZaGnKR8YciB
WgfTT1eOqTwm/7kchsat0QI2DOc7hDc74XTo+zxDqoHjiYLBXM0Jh5INY+bH8Pkv
6cEmF1CmnRSgE+UMGEbtl1G4pNV40QUVhkpIztFsqbQJBd6BpQHkmTgKhlzoxnvJ
IaMhIvkL0lM8LEXFoBPaXU3MWLF/ZV30f6WrnVQam8wonvuw0g5KVRMqud7LB56D
Szouv/iVs1AH8g4peTw+ApHi3jwCJkZHosKARL1ejp3U7wf3hvDt4TtV/dxGj7ls
MISwE1g4hwg8fezBd4NLMgYKFaWSQQzNiJbXWhZunR3dHWL1S2BjtGhLshxL4hTA
iUbDmll4GU39wF9+b+xsgADPsN8LxAzmQ6+3Llmt1NcFm6Bb/X1hXciJy73hgSHE
Q/5zqd7/8zWAGckcEeAFfTQEmuEognbtBHAZ9nd5msLp/zfDLLFcZH4X/OwOLgQT
VgkHg/9+sFEgw24pJVdd8gXMFUkezYdBPUfPhecLeYQQC/2Jfv9oUrX/jwjkCKVV
Dte3MwoCrnxfAqwqjSP50v9tiMBi3JLdM0NHoF57sviiNaep4wkD22a6H8t3of5O
296GTJreJa1ok5IPukOpxpCVYlh065ZO7Z2hO6uqTqvY2BpRabkyd1BQ2jiHR9yw
Dm9W+KbQqSTWa5cLntIElRbJeznTP37R37RXZS1CbWeHKuE4bkHWoteuTJQK9AHt
KTFY4GYwzmSn8qItPI9VWnXjh+iAuFbzPr5vua/iYe9DEXuF9w5mwmRDKG2IVJ5E
bCUrs+npMWFxutNSvIxjcmA4y3eHqB4iVMN1XkelW/BpZwty3OVPbMHYS1tt9g2n
UZvzJUNN63VtIOR7Dwpheluv6FkmiYtQdxQ+zeOQNdVn1HK0XYU/8SaoZ6Wp6wCj
b6U1tXDN3mGSPax0gpMhaB/UA0Ohtv5ErhsbCKn3DHpenwDffPeaCapAYGhxDqyI
T9qtcAodhSKl1k7fUZk5l8x+yosrYy6qFmf+gQadjhJni9dxWOYqlA9jxIDUI0IF
sYJkLRcKv0Ib36Et/AC4O57RltS6nIZue8A3gHMazcFaBWQcGZqg4LWG+D+ILBOG
5AVjk8OZ88dUqc3eEYziRP5K7YyMnSwor1RL00pTPR1lvKUGLn0cY2g1VI6yTWXi
MvtMmg2TA8pqjmcEkgrRV7Hfd2cETQLRsg7yH7bMT6AdyTVujkrvHBO0et/yJ7+6
XgiRv5bOqk7qOMLc4EwbFNk6Wt1V1ip5K/3+K7r3ZlqSpNb3g1xtv1Dw/FYABF6S
XeuhjxlpKBYQa0QPRFekxHiGsMcsMg79/K7W1foaXIDEVa1v1cqpPHkf/hMCh5+/
JLrS2E5MwBo2J2bnCGmk8NY0oR/n/tiICmuZzMFStSauLHQlfX5uLSSOHwq7t/W9
VCWUgpgwMwUef+Zk5TN28z7+OmWXFLi5OzzCDFva43A+yOSfHFFWBi3FyUhjraxJ
jSFHuWIfv2RITrdIhObXJ7TWOk/eLPKA9942qJDreBDk8cfEA2mCWDHMBdrazsdo
wDPCmW21R2zd+Vs2iuGG2FePppEFZtNfmz3qU/cZSmTaSIBGt/lrmxrmMFMEV0XV
oih1sy0ZrEueZmiDXm17WGzM4TnescGLX7QpicaUlKWUitUJPNAMmh7mt47COVsj
THeSiyhamz6WAZaHYZUF8ZOKxdYAlD3rRaYYwu0S+hAG7p0ZVBp8FneDObpP3v8A
8GqZGuan36YqPHXq6Tr8fUNi2RQrBiNMqb+7mwslT/WxJm/7Vym5TMu+zr95Vz2O
VQdv0e9ileAsF9vyFW0/RyQx5dw7xZTjYhgelMNEY+7F65aFGdr3BhtlkrUka5M2
Z6UyCndiJhCWHLkoyDQX7HHm3c1PZe+4CsVQV75y2DluHlFYH8JrXu+L21+pSF4k
UkqsGKzBngFAl+YDKzczGm+K5PXpc+UILNSt63tmu4P0R+QJbmmmRuYXykOVknnh
+m3TNL0Bq1DMmkFLcuyrgL3+PwXY3tqzEiMcja4qUKN4VPDm7WfCSOoiE0hS+qnM
CQtPEnFtVNcUSEAy0LF+hOjRzlmXUYnU8ayvwY3NZWQCMG8p4Gt5alBoVX+5yUwO
rBy0mK8zg7Spao0+711SxgoTIJxzEPIHuFX6XCf6LL7vNKVwRxZgMWHHIe4K4wEp
M7indL7bPhREseSergpVbmvmxGesBRaxmuOpA1CI8IxGEIWLc28mVYx3/OqEEr9s
wKjG/wCajEv15fwTL6EfNKcTwzdQ/WPl4CGRhuo11o8Bj8yo4hXjWR9enjd7AQWP
k3GeLkGXeufQHMrnmS7lpAnoiFOAQj6d5FmERpLfwPohfzwkVABxixODO07zvdm3
ZbdsI78T9tWlNEPsZ5n7PYOKksVdX1hnjRzGi8caAus+53Wn6eHmbYILv918c08S
jWx3rL6ltudyiQnTKiVRw7Op+HIAUJReGG9TyJohV7L+KD3hKHjIYwFJ2pz9j8LD
ImgQ/PFKe9Krl2Omtt4urXkCiqHFqOxz9JEgYUJA8A0HEAL2Iwu7+/qkqHLlYyMH
33yHDWx43Sj8Rt1t/1mnjIrCjDRzYkAadIzJ1DnKnkzVCo598WrYuugEUbNmpyCX
8wQNxm4I1YCC3VPF1IaKGjmxKuyWQDHCVg1q5nymBxmLAgAC56721THVj8zTSzOI
aH0add6sfDdML9fWY2Fi2I02Me8gLJK6aG3BUnoYIICCZWzMsOdkY+A04eS2reuJ
rDvxuzii4k3PKCTXcBQLQ//yEU13NcHAcMv626wmdfUa7FMzI4wrpgfGs8WNhTD1
bRToWL2n5CRRNw4JE4wUHjHDQQPua6Z3SX94AKkh4NRKEJBPdsCoXC8PZpHcllap
HD0SFXbZ4PQckdcplA6NJxYjso9shw/CfLL5R/rfcnj8ruvUAxPtwc9eNCOx/0Px
7x6WHVbwFHT9rXlYDkqeLZrv62seKU/iKOZavBS42GKzbSl00nhKNDLu2QwYi7AB
Lpc5Bu7WDAxch200oLd39KBJrWwR9yzcp2FaNlVX4MuVlXIEk5HFzG8xdipzyFpn
FcDGhmxHadE0MKHc8uLWl3FGz/ogv/YU0mCQ3YGETveqvcUfB6FEDdGLzCAZFDlR
qddKlaG4Iu0QkECkpAp+X0yGznElLq4mna5yERsO4N6xHNcltL4zMpmQ1+tVMz84
MMfjA+xLhz5Bk/aNUA7UUwwGna7ckW898n8Q2GYC37crNPbSsGbuWFzNfI+sYWrb
1cvqjW9ORDGfYpWGF11ByQPrLCMKEG7Goxik03I/Yhr6TPpW/A5epNWa1hQXyG7w
AZiiCw+QhSxc9Ap2Z8nZ9EqwXGwzVGI2zer3iVW08i5eieK28qS8xC8BVoGHneCf
ksVmnGnwTku+a5dh4TkdEX0rWUaxIBsHjE/vQk6EK4Wj/DZeXBzx3aD5zWg9MKkO
UpGEomP8pt6yFFIeiXwS/ee+00iamEUVX0+nLPfB4Io/Wyhsc5J3ac9jjAn/UsRv
UAGu9WuD54aHHM4pLCYl87Snzy7Q3QffVKpRQLfJM5ibdsC7wTIPjUjziuBjHYq+
2bXhSombpm8y/8zrtfD3vT8/AhQ4jP7T1txZu51VkJFFBW6+L1FViisVDD5s8Gb5
s01Ea7AQO3unj1YBErai9os6KYHPstO3fu5o+RIBGRcFqcXh+P/toI8qtWPY4iER
1XtX4EhC+FpqQTMII73h8Zb7qJ9H7tJTTPoMbH/QVFkt9AUvKwqVXrozz4/GWXDY
Xvuw+SzsApFm45ZsX6e4F1LgQOLBke2PQejWHGMbo7FjtMUrJBf9+3swDO3hGyjC
a78xf/9wosp4cDxmNf9vDt1Poopza5j29zeXiEQuJkA70DabdHu+xRI8Fhh2rTX+
5aLTnlmqWZymavW4/XpIlwfAvsRZGkAbPVpa3Ci1xpR/zSnaGaLmzU96XLdzqXFr
+Rj78dk92asbKfuwYYxBHSDu9Jxbu75dhWcsvdbxGfGS9HFrbzxDnzk//ieMgFL2
Fnb003BHlmwrelaQ6tA0qKiMclvAZoPrXdBHlMfiP6+LmWRnvBHnLzasXG8qT0/S
iO8b16HEnryIOC+uKMoNMYCo2Qc3YfhoSaatxWmnjiiLDHeZ+FAUfYmrOdFiMLGS
IDracFj/yfdKZlYwH5ZtciuoHNnD3uob1mR/uXDhbz7GBHoLenSK2YBeBa+tBOu1
+enO9/DxX7Rp+LWKGhX1bKBkcy3O+Cw5Q9YocoY/bEOnh9d+hYIK9OpYheThZPnC
ZKhyHK1OC7IEzM/Nwp28oYjymxwdbz66UedJSzkF2WLi3daC81MbcDo41jNVdsEg
oSzU3zCNVPIEH49orXkNnLgxKoAg9p6s/03jcRYFeCPTMN8HuRD1M55aItt9SJ9I
uB0BcAEKmQjPI+OJUOALIQ==
`protect END_PROTECTED
