`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0hRYorMAYs3xb0LgJ4P3RDVzSD8Rai0mPOwDuT8W/n1XR6AMOsoj5QpnVD4AURU9
KxldKBLx89odqd9urEiYOAGV5UN/NggVyjIV3zQqV/BZRe/iT6vABgtyX2uB+ROL
+ZHdQCeEGHnn6Yi+EdLG5ib+aGTGLmit616P7cIXHZ6NXQS8pgieAWBgTfi8caNl
vs0HSreUG/ie42plD1wM73RTC//tDT4JSxph/S6dco1gcdzVWb95FdBzyURtgj5X
6b5WnfS8cJBCpJ2tUepjO+FWuGrmjXxvnui5cp7EheSBIvYbYUIj7ePFL8dm1HZl
3yKo9GebuX9XSTImDjE/oZvlJMrdpepQ+1H6opa77odcQXRgKGt9TWERCvnNsniS
1QAbqlaF/fDSms3Oc1kcVccuv9BAXWiNp0kOPFiZZXMdnBnb6QIdgmX1qx4xBFFm
um31AMgic7JHpqD9yfznz5CIYLh7iqyNTFA0veFWvGb7b4Jrpi3XjMJLgl2Zj0Nr
P2VutBdPJSz8j2q+XpFeMqkTu3HrJO7Q2YgBUsJ6S3Al5lkD+MnCFsbntQFLyoy5
mWQl/umzme8wGEZlEZpdjx5ebXCcL+F+bVYaNGNfV7sUJ9z+4AIPEO5uD2/1BGHm
uYR7SL+d7NoYM/3aYooFedxRWR9jhKPCgEpBi+cKfTtNESrQdCcYlVr4wc/Dgnll
8VTr4c2U59G146jfdH219v760jWbPanI6KoKoEdteOFFkwm4I6SxnSqm2LZ0Wdxv
9rNTOSdqbcXsL7zqKw0wDSYvkC29z4D7IR7ULnTh1RpguR7ZiptQcH1HXaILbEys
JGW93FURslyKiVYBY3hqC2LEKbfvRAVO376JTK+ZgBL2SrHu/o00WSZzVI/0b+SQ
4apyhJjo7KhvBd415KqmMI47UCn7AZbJXLZ4JwkD4F0=
`protect END_PROTECTED
