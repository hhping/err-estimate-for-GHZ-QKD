`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5tXW+GrDBkYQ7DZDum9aj8EMHMkyRmc2CRgROW02baN+q+ixu3KLybmvmNVxzndb
dRyBv76PXw0FBiX5Yz1q62wWsTxCT3M/TM8NZYrD3oGmdAYOIESjBAFSKSGNouBT
ciM4HOP0d9TuyOpDsrGcjtn1Bo9OFBvHn93dx6VRJIpSe0pBTDy459d9NMHr+iql
L29phtRwlPnaUZj5m+jmpyi+XHajIu98K0fAwOKR9VCtYkTdc1SQTF9YTPmWOICl
fOq8fV01VzUl78M27vrarxOQeItYZ2N8j4O4HrtkZfOZGVXeKDGRDOyd3/Yhy6Qe
lDhZWwVUtyY0b3UGz+cgPwJGGCYKuZ3f8V8zsn8RwTz2qlPWMSAeX7wJJ6T3XQiN
fngHbMy3Q3ciagtbUlUNDMvkuZn9adJMxXMbpCMyq4Wub6oUukLi/ud72OnXu0sT
VIX0fTlrengauIF7PcXoatxTiLHcUmg2ZWF53L73XzsljcPbJJCFiTQdMo96T+Jl
a06ZgbG0ZYfFYliX5yUWdg+S5PXkZpbhXxvz8cqUPRwkZwdlc6Dz6QmFQ395F0BJ
z+vGhGzi1srsEXXj29hmfnRP93zcQD2A6jaUhx6LH0baOQY7GK26yaeK3BaVE0DV
P59VOEyyOSUEkICtQzWV13ZwrpVNESm1JwlOdEABOHUTY+m7xnsckuQjxScp/nTH
XVxZy/1VTHhl59XuRAg/rUmyK4k2l+62DqnFql6MclGl8dgjATd3FBtFOzpCYuxc
GVkqvWcFwpR2AtY1A+ygnkt9dDIhtNNn6V4q4uytuU0PtMmZ6PEScv6Asv7yR8nj
CMH20Dqn5Z+ltpPPkzvXtGM21MFrV8NomLe9q2L4JiwtNUtvsDNZSKbF8y1fTsIO
TcGAidb+xrZL5kJMeEFMPHmkzqxA+Z4KZSOmig04hcT/cht63nnUxfrcGU1GW6dt
RTbr+aG5VO07gRdnmo4xHm6EVIJOXbXr8LqnFpqVS+ThHn0LAuGpTpHLc/RVbgNo
lVS83cd/Fw3iS1Oq3RSoiEcgDDUk0G5I5YfieKDxwyd8h1ztMUBAKwG8KGRBW5ze
cn9s0pU7HvEa0q4SrtywBNiyNpAK6ZiynaKP3cDRFrvt9W+xDfGOOaMZQZmAwKKO
8ARrQNJG9XXRa8UK0LNbGcurfRihRqVkoKZkeUuaU3QyO+1u5gKDa0GnwqKmUeBz
6u6hT8/efNG/18lv4xk7j91lQDFCNuDv5UQfowsu/50Z4vmaHNoRFXjzsEoOQkNg
FbCPjOYnh4YuXVD3MI61WXEfnGgI9xW69jA5CKNQ8XAZ93ZMvtoQKea88g4HsPHy
x15qI4GJ9kRI2MlVdgmAs47zDOdjg2kJlInKLIyCtYtTxJ6CmDrmZiuP3wksHLGr
rd3sLCjCOKQajzBSffL9hu0DyRefrteuEE75RLTmpV89BLnMXLsYMkcs0fy4j+/p
looFpjHxN9U6F8i335wq/V+kIy40+roNyhOkjaVMcCWvGmgn1ribRrZ9nQrWlhu+
oCvi0J6zapAFCK4ylbBcZMbf3a2d5eGY+2ELNNtuu8/b3o3O3J23OJwP8xtsqkqL
3rLuQ5PgBCrLwKrrGzyiQyeN3a3TFkSli3XxYsHIVc3DSZcygxIotsBTC+Khn0hz
kc1UO0ABqpme3iRDRBmVTdka11adZXg0ppQoi3UuaUXNrUaARZBZK9FgaX/NtgmH
4pS2RB3ti8kHiHy6BAemRgYSaZj2/rnzIXHuX7/lLeeCxknLtij68DWrIjDj1/IN
7IzmtvNLIWjfFXgVVI5Ehw==
`protect END_PROTECTED
