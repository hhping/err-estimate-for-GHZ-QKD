`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CQ9n868MPPvHuFpoCcWK5FTxTroFyHKyLxhHYBZP/3g5LRw1i0dOHSNxcFQz+AtC
kipu+IiOuDICrWp4NLksNogLCTc1cjI2aYU7OoXP2DbQPV7OXeIdDnhTUbc8MaV/
oRTODjQ66fCEMmZAptMcnk/zBYVf1pmQJg84+MvgAZtNj5Go7gp5NX2ydZtohhP6
DRnMj2YoJ+Qd7MPNXdrOyIJL8rYhm9I1yRhfH++T1v0W2Lfb1GbxZVHEZsxx5829
3oDRW7qYJc1yxtlDuFBQmXKeKcO+1AQVw6UUooyBPLP0RQDoeL2cYiR95WUFO4x7
xs3OK8pt2SANaOfUxNsJ1Wf5uf2EIaZt6YTlY2kbxdgCkygRxy6b40XiNkEbQjmQ
5M3HyxK8ya9utC7uhmuso4QI8WjIQzRS/jEl241PCkoPRyTQTrQ5b3iYK78W8ucA
f9mINLSn4N8VWHTlNhd5SpHpw7hI8w3zT4yvn4yD1S3oVXFLLfXJhtSE8pKCkMoM
8fVkdWDPpoyBrqipQICPFTS7iZxB5sWNIXq1mpQ2TCkBB2w/22/oWhgfoqC3umTr
2+/nmNTxDmIgx4x0bkrQJ68hduRDyERhgxmCPgVmdiwPFeqFjZJUMjMqWPOQuUy+
sutOjSBWbW79kYfxL4+crxjyFQ4KItR2WDUxUv3XlqPZkDmuq5kIixobI4V4b2oE
dijr6toWi8/BqVcDvk1NetfOGlHW3DsHHXhngTIDLmglmsCyzyBeRcjN52d5UOZ+
Ukytj0V/vQZytKvSv1BWIB0WU2tNiuFG6ISMMDHLeQMvMKMcZFStK/m6pgTb9p3R
nGzGe5eU4E2LWQMoU9fSC6pe9hXnYjCE27D7y+S78/rXUFc4Lufheja8zY40odWa
uicBIU8bG8ZYhVaEk4ETAyaYMgGjBOoKHhdGDff15I+v9rQ6CQSztnqfCSYlLS1o
yMNLhmXOiYAZog7XVvhlUg+5CGSKHip3G1e7Il+PFwgi/wl+b2DKGYqnM77FIYrS
4T85gGXGUOGWGJhsqVTXy1zXL0FXv6GWhPnrm6RWDz3xSflGQVNET0IkzHnTNde0
G+RPQnj7ghGkwIw53o7Ooq3T7BajU75NcsYsBBgtXvyRDBf7OjDeHxDj4Cfz1cS3
FS7UWQMoNtfUoEj0n/PdhylF1xPpekqPZuhEXn3wG7vj5OTG1U2PMCvpJA507LF/
vjuCBMEZqzxXKMY5nErXNQH/4NOA3iy+rS4jr1IZJgoeB2Xt92hiQeIw3dB549n6
rkw4h84Lh31XXzolxtAU8Sm47t/R2z3/4y//PlSIwo8=
`protect END_PROTECTED
