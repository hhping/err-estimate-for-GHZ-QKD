`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AxyhIhHlWKc0czZVVzU8K0V1dc/tdEbvsF8TA542XLh5eKM9CETpvn/sE2CQ08/3
o+Yp+hrQ1eLVqOV88PB0SLtCZp6/VoSfRrR/aee7M11eonrgac+k/WrWFRgb9GPS
yb+VzeNsjI2p2oQpRaJc74lZDKGgq2dGYGSC7IvXy5zAhlgts5VDhYw0N5KI2k+l
seLs5cZaNKfY+MDpSMZrApvne0jl3loznf93yIIuHiS/iei45JfX84v5V29BAzfk
MQlIcnRDdoQZQJ4cOvhlYA+WaE08/Pi4gIcmWuNSRdQ6GVMSnNncddsOEvRqO7cl
x6FCsI80T+I5j1bcD98C0drYAqdE4lmmNz1jUr6d9EU=
`protect END_PROTECTED
