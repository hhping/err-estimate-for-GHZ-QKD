`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BUrLwWN6MucCslm7yaLfUWBVW80MOwAhgm7TK3sSVZLfvI6LfOsgMosinmR6cQJM
V8r7qVtZ9vWeLqgO+RWvldBRrWF1U0ZJKwUtnbfXBD0g+1wZdkBueDQniW2jsu+i
UH0s35M3eTWYpzp2LZIg8hkH+HxcK2OUafnB+44yj3VyhjzOPBCOzA0NqWP3gWnt
ukkhl/r3LwpKVpc4hKLJ5aFLLTzg4sM8uVlS/yaOizCCW7FkGZiDz7Y/4avpm8zr
dUWE36YxBKY+4wXns4BgI7Mee3fJDOMaagU/BeOtwkViT+6FbISEEixAu77s79Mg
q58wWuY86uqyFRIjRSfiCbV47jt9bGNQHsvzs0c9alAaSXvAidncnUDeEQyK9up5
ajt2fxCwq4UA4MgEy8oEXnmEUDneaLzaLIzyVgHeAaE0ryQwxEd03EdQvtuOPx2b
QGTavNxRHfHjXeg0GycF5G00SvFPA0pByO0wcc2AUZzkzEPJh1Rcq2jIHQax6HUi
LI8D/CTRBKEOniB594jjsZQ8EXtGTevf7GjrxkDtlCdfgAIpJiBm2G/kuqaMMUOL
`protect END_PROTECTED
