`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mor930yKJOEJXeoEuoZWCPPLKL0nQxvjJyc8hCXtF8qw5uWaUx0BTbfTtRjfKEU/
uUqzem+l+W6h35Myee5pgDMXocCBkRYb5KfTEJ+gcLN17epQ/il2bT3SjESuwjo5
zDN7ZiTWWNL4hJzVj3klXNluJsTY3AeeeSi/B5GTPCFKx0h3A9Dd1q7cPzd8sesI
Hps9DYpmCkkOpzEFXICEopXpeimkx5jOxd49YX6o94j6yfA0JrM8maJ6GgNjLWh4
ybS4i5yNC4sW+htSfOlYlLRnIbqAS1jYkGniXAKWSunFh4nhuZXMilpfVcSmV9JM
r4/VkPzaYa7jf94zQWA/DYH+0U/ccC7ulbfdgVM2J+Z3g/QtO8sTyHUcquXujnpN
QY74gm90pY1K4vIMD0enJkEWyvoJCyZlzkY7Jtvx/nWqpk883a14SaKLzirz8u2+
FQZAdSEG1+NgI7xgdNQ4cYMS9S0W0WMTqJcYt4DtFudQrKLZozNiXQtSJ49OOmGH
n439LPwfTXeuw5/ANnpduUysJnnsbTmpPJz+QzasGM0SAgSZc+lMilTFCW84rJ1v
U0mH/TJLb/LL4xSIuoS54IZY2WbWyIWsCOeAPll51H9NkI6F3cXB3h0x5q1luFD7
9nVyuHtvLbP4FRQJEfcg/QxctHaSyPDUb7b5Z60vrB3krA0a8LHumFOmPI5yPmR9
HLwCWGBHBYfPnWjFSfn8fcHKNxDcenWmgF57MhzkdxJ1bWvV6e9pXwTYPS+Joeel
c15cpzuSQdTKfPdWWUqLpn62hkki4gS680mbNMXU4SxeUR40Mr7pNAz4VREqSkkA
lPCepyWBFuXmdw4sowpfT0RX5CTtTZMNbL5SOWhz73yESRq9nSqvstZu/Rtrou3T
Rr/UHVFJH9vv1muxQMWi9G8LQdZezdNL2EkYYPngQrh8+jrGzrD8bWAfjiq2S1tc
EarooQkDnF+3XvKgg26EERBf9ur+CCzVFQlDziJgbL136yxWpTdku7Co6ikNIYfr
U/z1mRFzthsx/rqiSvp/6C/sNFvPLCOVQBT1kYQ50cadYZsnCG5wO2UZPBZTgV2A
SHMXONBPZuTUCGFqvI0QWtFTBgADfOX2f3D/m0MkAaqt/BLrPbbzxXwjG+2KYsS1
1uR1gPmTlrsfEuIFTKDLWmPkPgXQ9JeHQB1WOqyG1mq9AoImL9WHEGUCuZFoEMWi
NxuGiNyVrAF0eKtMrlqtM+0FMBai+nRUruGyXT3sWC9T86Ds9/8fhLJk6npJQKmn
u1+byx6rZk2xPobW//5KT2iiWCYc/VsjSkxfI9fm3AVQYQNtvNUwh4P+lRLyXG86
j9xP+ZyfzE2MU+rwyN2vUE/6xwdcwMUEIQfY2Z+hj2nCZtRNIx3d5sAaBAnqfv+m
b9JV8EpsTAaZAZoFLlO4/qdbCr/Zh+cwbWLfJEWW2F7JTJW3tyU9w9Sr/KPzin2E
Cqd3SRhRQ8mmNDgRUEY8sDSTyFDy3oIBv0vCmFt6M14ZAX8mrHxMmGzca+NiZKQg
mlXH1OP1tOAGtrTA2d8CZbhlnagR0TLhrkR6BXqgrsDX4ctvWLDvES5kNugccpqC
/PaDpLpEing2oMwEAJPHfdttLixzCx9Jd6giKt6HgdR5KfI84nw0LV1lz5DJwGUd
3PTpOlLlpXZx8Xuca8PGiS6Yv1k+fAjjuH51pW9mu3OkrEE3Pm0nVq/HD1Y/+Kex
5WnMvcJf9wmU0BS5BhxmAggLCfkKCbDhgBMMWQZPq948XJvk8IuWVvrwIcKzBCxU
uJdNGY1jQtzty0V6DjK0MOQaYC+Khn1liSeqPKbpbm6zOIBUjdDfu62JwqyR2Wfs
i5QD2MwwhCmMLULNWKdnIcqP/PMEj6hza5FANNk/27rxTgB+p1mlFhuM7N6h/GEu
qmyL+YyixK5lDhzRFfmsDQ28IfW01/1OC0N3Vs7dpwd7oD5PtsPO2XHA5JDpBVJV
WqAy301cp8MYKBEmSo6SOMcHQ44CaC677jOfl3nyYm27hI75BYIkg6ESNA8YcEz7
lIGlwHwxF7+VUDZaqsAR4Hc5DSoWmhh9x8iCSZ7y4u66zp4JqGPbyJPh/ZJdXPuT
gHRDNCzrTseoaqwShu6MmG24Q/AeiMub5oWXPz9VWCR03OtwZT6z5Z8gU3EYU5vk
wdtUmUVPp5ObxmRFqaSrbhHvUOY1YGojOrsk9YT6Op6f4VDENEmmdlJeFytoy7i1
+tFDqRPUMqbErR2w6k76j4R6wqLg101LfBqrbpASJ+/qTp3bAAPOrwFaBKq9w5bE
50nBkkaJkdqk6R13fnM+UbrAezIvp2VjLvLbVV3YBm3wOzf7x/wIy0iTG3Wwo7c3
zZV7VSnXhMtfieTVkD8Il3K/j9R8dYJSVMkWuQaZmm1Y/m61sTGw51PrShUICyJG
oqdPxExRpGr1GtBrz7n/Rny3TUUouZEmuiUmZYTPVREywaGF0nel2q+OFeXZ2eCA
fEuZmNxtkTz7QfKm0rEVAk+MrYiO2HNe2DBNtiRixVGwCpLwBdOb5bVaet7WfUNP
K1ukPol+7iidcBzCX1U+xBl7+6ykU5u5Qt/wJuAiaYUy1uGt3DjNV2N9Zam3ta9q
i5f3CLle/E+Y5PZCxb2fnsNTaTJmJWHQmqecOrkfqM+eSqhw15aig0xEO8RCZnsE
GzkLsKTaC08o+FZV2xO0Wh836CxkmSLn7IvcTI1b4OdSgoca3Jo+eY24g4HRC31j
tGgbO//OXFi1DqVTxdbsrd3X86JgZHa9i6lRL7FAfB/WKMunWYbCfpcGZ59/kNTt
doBwKZ8HMyQ67IpXinuCPYA3ksYsfUEfI4vZqXPUPY1GDPZN31EQqkD0+vPF8IiS
uXClrWsGicucuPMKBwM0rK3cyZ768MRMDHlQY8dOp8/NuALn0oDcZ66xDiMoetq/
AujuDoevMCHH7oF5yWUMY1rgTXVNpMe3VgAl86kPJFU2qo22LWEPJL1Q3qTolf8f
PRQaNCUCFBcCpEvIfVxPhuxibo5C/MlQIPlQHTfOUNSn7uUG7U4HQ1Iv5ASsaigI
LY3fIK5XgK0RG7GNeQ40hAecQGJk+QPlyoDxoqWnb6toF8HV2wrF0zpGJ7ehtjbq
65ykhJ5v2fUJr8z/y/sddPs0mxra3KLPb6SqZ7Qlm8CqW0dC97b/y+li3QWJpKHF
Vsj2nbZTo3h72NG3qrcNXhST/JKZw7BlrISIHD/K/EbiF/HBIPT4I8+ToxylFqk+
N9ZP/jOEjAEFAIFYtxoCxw+WqFOZNfXERc/+xtK290mCWqcYIlN3DcmpnQ+haZUK
qOzqZDmDZktjvC/W2XQbEcbK8C4Zcrd4VVzdWGrJVS/tb7UVm+orVQNQ81G9Qj/p
yx0DGPB8S2ymm8JabP6dDYvRoX3xrWm4gWnwVVNseUfYjl8WxCZTXUozGoyO5ItD
de2eaFwzi0cpsSwOtua0IQQMq7uDsRWQ0aGatVECstLE/SJHnD12k31mWCK7pxTR
4kvpne7guegZKr+ZnId7uaSVEHcwvKWf+PImffWJyIX1Udd32nTWtY82nmU55b6A
jCowOj/D3WOw1T//BV3jv9IAC+eRh5hoABxwo1r1tf74YH5nY2LsYOFfcq27R84/
uVjJAMPiQ2edsHX2n3QVY02NAcDsN8XRVxDNWGypBNMJvMQH05UnGl9Nv6WDP9Gi
i3hj3ws/roEW2IZB70mpcEW2l1GJ/RHILqrgyZFcAF0KNwylpN2iG0stLf6dHYCE
MECHWcYQwkvyccpX8rWf1Rt6cRVo+E6sf6xuYjBkurhAAZfmzs+sBKDv+Jl8J4uH
qx/btFQsQ5FnmoPKne0WLpsFXTRF56ulqg0oePpEc8VAt3IcY0HRLV6J0AFgqD0L
Gre8vcnjHsqrQfaQ8xmeit+I5aDG5D0i0OrDv+lz/XWQk5+DVGFaTK0VtG077b5R
EPrQysgzbCRiYOi+GxyaU3Kd/g7WM8aNHDsVM4JkK7BSQiAlmWdsH/p5kQdkNWjH
KAkfUwQvTaeVox3OYFHXypIBbT+UdPhoH1JETZ6obPS+2RcIabJctSOie+1Uo1jm
zNCE1j6luAnKU1duOdrCj4zhM1gIGqK0e4Ob8MP9iAY6TqTiow4I98US212XpPGr
mU9w8LWIL+lVXwLWInEyxqQbdO/gQXc+5tBnfpXCkNMJkAp1IsUfXc271DDgt8R8
0Hb9xilpHpMSXAkYZnP+KvRcWg969JfUFw6WCfRtn4CPQRbbWrsRc/Zw8Tb/fvHA
f+zr+j/jfM3LAlOGe6TYJ3jNapf6ntCkfRtA1Qxr4eXL4kP//WRKGyAHG7dJE6AG
4LEjSMTxkG/29OVSY0PJt0Y/LuvGV3UVlPEbVKwbjGtJlrpU74UfgV5OINs2Osal
idwJ5H4zD8TMlEZhFy7ctkxI1JcpRKzAR6Cw5ND2nThFYP2805I+blGOuO/MEpgz
B2XNdutQmTfK1NJacc+99/aHvzGSXcL5bHbfRpg1C1dLcamT8SE56KsctZHsyHyk
tZgaMz8zkHZjBQT3hkE30r6zAaeyc2Ths9SmnoYLnk96lv7Wwy9DrZCoCMASmOPq
l5f8gtvo02+Qks7b120QT6MCc55jC7riZjAhjvUVv9jt7Kj7CJeuvKJ1PSpTAzM6
PJ5052BJwykXK2WBRu0GbacB12CD2b5XEhpTg6/v2bxdnaEMwuQKXdAJrMDagMlH
xE1YLsleM5KDspHbzX6a/6D3Exvjs/JpYO4MBaN0a3EoT2jg4mOKzdgkP3JfKTcM
Wnu1O+3KZA2Y9fDqc8YV2f8AAZ/paQ6PdidaGZFF7gliuLhy4mO6uZFkINhRx9Ru
aRokPifbi9k8Y4+hsvtpox9ZDsZzxyI0s+IBTkgJtuTNku5ITBC2/bMUqfdP/Nm/
5JV3ComW4A4OlxGWcIrimfsEH59bGoKIo5Qw48gg9buJw//EgdXbM61sSLkS8GOJ
k6pnLGBs5ufJTB7kyeuU+A==
`protect END_PROTECTED
