`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UN+SOqwQDEvTOdrwm4jXJxMeWSTFlEWeQHpJxqXq+oyOoweV+613nVGqNjeJo2vS
6voyZsCx3GcStfz+tC15T/d5vy785ZPGRoXxIdTj8E9CeDgJmVq9WAvwo6QcsASK
6nWCIA6LTbFyZCQLxASU5DeC4EbNGNw6hif3JYrtjdSCe8e1A1J6ehBKd7gIfB1n
S1VOf4InudCPcs7dkawKy2/wCKCF4huycFQWFFpDIwMBJdWhYAGAH7y9rCUNd2QH
y2hbDb3Qw4+jcoH2s2C9X01VFieo3jR+6j+5BX5q/F8nUFIR0Xv6E9narPghxgzq
7C+m/XqSYqzEn3lKjRD7auUCNuw3n9diMlV9b0M/OSQhB4QtykfT9suVXLkzD1jc
c4PNsGH5yyA7+HRGroAtRwRJQ9hxRWInglNx6oCNsah1SbpFc72J8D32erAYGk9D
WVMi3aFbLg9yz5RodXfw3odaLzPVK8nosgfeB5A8j/wNa1OvAxP0s0NJ2wRTt8DP
bpk0+W0TJb0BA6RxltY12+1VR5hG1+qJY4k7nIS0zDfi/Xo5Kya0w8A25kgqtCnO
h4gY45ffHWALeOV5J8PlTUObiFMHqAkruNkgeHwqDAqimfRdLOWN2WdspGqUZ1QB
BLoyOAez1Ec1mYVI2IzVtKJcrbqMJ21Bwa4Y9kUz0EuGk/yyQ33sBYc4luKP26n7
ih07xiAO7xEWg7tOqQF85Tvp+vs+GqC1Etx3LBRf60e8ejAYrzs1uiDn5UzYJS3l
CfC6lhD+gpMTdELRZEPJKEF1mMX7nstagFjlbtHtPat1Qu2JdngfUBxUe3mUYQn8
geOWiquzt5SslbIAiSjt9rBrMnJcsQsbOZSZZZQgNzGX6Uae/89gRK7RHajFCvQD
OxNG0Jk02Mm3QkcURvawjx9grPgzjRTi4O+aR3aHBIjF0j71T62h/UcfJXPnm5oK
QIAc6zr8FVxgubwp3vB+lKFRK63XxLZLZRsfkYlW73rCoofdnxZywz8H/R5LJfCN
06D5Gjd+ooNJcll+i9CUWDsahG+rk15itzGCUaDNU6H7GOacFf6u2esEjUIdMI0y
e6MRPK5muQ7YfUleQ+DxHVtPU8XV0kzqMeW+zqhpQB/s+uhIeFgrRoR7S/hRZD37
Pr/BNodMMhpVqzGooeJ55SseKEpMc35S13G+4pPuqgllJzQLBWAlKFjpxSLOOZbu
V07TFuw/2Tq7FvGmf0g1nZSfE6e4Hz8wmjhCjFTIZxrlbSrs2f2fLEv1vqI+tT5P
C0grYEUBj0kTnGokiF3AamhyB0DxUjdAk28kofl3GXiwbkoaM9cmHwryAEwr5e60
5h5YCXcTEhjeO4X6R70S2+Byx21I1AtFf/ZZhOZ4uJ2KBiytoGah3yAzKyEqtvNd
+9dlPSVmM1mPOIMGJrq3+StAkCLwYjnG01yOXcrNusoNQSw66idOBf/oPYecJde+
OBjltaJNvVjNv3W/THmjeGjVBMFvXYVXvA4Gb4myCAtYyFXTENgaF131y74wv6nX
H7XHchtCj/2bl/vqojGZe2UHrwiWnLg2GSKpBQ51kT8JRa+K1uDZSm6Mr5InxKoo
OFZ+0EzusWY083FIAg+pbf/L9g2zM0mQHPf+2doDIa7ih5wl+AG+inzY1EyHxNO5
/v+xV3qqUNTXFcv2sgJHg8LPssmLvA+TBBpN5VEK1HaD2Pp+kAYn75HMtiL7Ub1q
xQMulrBFYTgfIHI+vbZ9hgaqZtCz3Xolt/hHBANN4SdEYjVsWetH8+Kkn9lCJMdY
ilVMMQIs+lPuiz0r3WFPxgXt5T4c9H+F1VjT3frQ4zeW9EG2VWiFjos/6CX9Srre
rrJXW3Dbby0oBJQ/JCBt29aH7x+2RhZj5w+xL1bTVvsQTgj57A5fxpHeeuEB3CDt
wopyvlBSNZqwk3Ea1cYB/wHFT50KeF54BELmh7OvrW91CtlMyh2770/pL0zhU8cY
Lf0RKJIuoqzW5IIhASjLK+fccSOgkf9wpn3hnJ+/ycb7wQAjV5yceQXiWm5s1OMz
mknvpqG13dbe7TlLsLMEIglvH17x8Lgcsf7RkSDB5XX9ZuRP7pJqMOmMn605beee
DJwqmVdpxEb/EWFqtUR94L/UeGOCTgm244Yx0WafwCJo0ygjjAtJHnX4Uc/DWQWR
NOqeyC/n0UcvwLazdv8TPxt0/rTXrzZFLxP22uxvLd/IrwJ6iOvxuSUNK+IYQt4K
udMs5vqOYYGiJQuCQ7PcWstbXqFGRta3UGPWYCvbHY+obkWy2myrWSm0Sf/wLM4A
g1Iy9ZaGTT12Z17Y2JogJPzH1OeXNaknRN4bwh3ImuvYgGconrOF8hcgEE9XEu+6
YTaazZjOXHzq3FIvE3ApeFzZl5hICLviEkJbCRwN+SQqfmrnj1dJyWLVAJuRUhuo
F2tHeLUFUJ9N5t6yPDSpqxp89FrXgWrSo8S2gZCPfZG0PRu3cRPdFFiSmWhKR1lB
Jonuq1fNLGIsGvX2B5zAaAC0Pq2vpTS76WWysHvRnBHBS9NV/NBqaKsqbNVFVcW3
E9n/Hm9qKtf4spxcI9ZAvuvkQEcYgC2J9f6xCdsjOFW5/6UjHW1kw1gklbL5m3pM
KD8egy91WYVXHQ8q/IqCyjdda/Myt8Y/EfHd5kJE8VQ5UHNVZVWcFv+9JAu1eLIi
7teILvKnJMj9cr82v5N/ARB2vLtCWLhQ2PUgNCjhGjlUH/gvqx2NURscbsY1Sb8L
`protect END_PROTECTED
