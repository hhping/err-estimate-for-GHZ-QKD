`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
geFMHvkwiFCAjhjRzBANG1hzSovOaqqRJgOTk2iS4nB03IthG6ZIOlikIjtG22+T
ilBV6ZcmWIVnhsmRCeVtqNisHhOrUwgqpj9ccnpnzytSGP/erEOgVh0+LleQyrRD
UrT4sNxy5ZaVkst0QC0zkIDs0HaOEO7Le8krOMB5xIBY6Uvp877RO2O9EzopW2Ev
y3b/Z84Trza1Asfot8CX0k9BWb3vuqe6eQAoYWCn8xLlAsZR86jU/VhyOtQ1Rnic
pjqI7uq4f0SpVKZnnPoGLc+JOC+U/zufFjnZRPFBl83S9tslpA32G5FkJHBsEtnp
lwel2P2e8g14DrN5HWjaFeer2edu5zQHaBidx7U40tXOI7L2iqZV5OYWNIjHxMiE
z+kLHCih7yJeZQ/NtPHKDKug7kPGm4el1IGB5YvruGZw3dx1Z9KfAx20Yt5WtbqB
LoDrB6VEZJE3z3gYLEgQWKiy8TB3Os6TRuVTmDMXMoDK33GqHsX6uKE/CdZlOggK
01xwbubgOiHD9ptZjOeBHfW97iAD7/ToUg4hzoAEv3Eq+fk8DzfHqog6IepG9fhE
hfWW0VcJSKizGQ0OacwZiK0ajlFDPxKrLVa0sJ4D/xXyBytZHnRAX5x53O7zwieH
gK7iS4TSGldm1mv0/Y7HnLKHx/sybeCWrPl4Ek1Dd4OuFJXel4t+WFEeXwxwwBQI
Mm9U3RGHKGcSuBbDLM5hktKpEAwU4Na1qCfEbSsbU+uI6OqNAmUW+zDyul6FzcfF
MFavbzReXylZVOxtDaUnh5E5sRF5muytBeTMQ4IKBEuyQkY94NF0H6QsBSQtjCC2
vC2yiawOh2UavD6LEPuNnaO9wWSzZeJg+v9VAmi2cKKk6phap15xyfHPVSE/S6Mx
CCI7ENyBOjjhTwapDd2aNuBBJnw11QPneiFVyJpuZyc=
`protect END_PROTECTED
