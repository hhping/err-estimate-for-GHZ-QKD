`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
loSDkWTOt/8Xz+RXuG36rBejbP/rZRIFJcHG4eQ79oedS5qzp1UJ+l0z2rE3eqx3
nmN/8lfvwRSvQXSXRHcyb2cqGZVYGtdXrvVSx5j17oQhYA0TKtMBMX/9m3Qhn0+k
ORQEXcO4dnvzoFHYgGSF7/KPhSkRlmwnId4hLngtcn3Q0o+XeFmKXr0I2xni/3gB
RjTJ0cdjoIj3Gs1Rx2fJN2eB6vlXtspG4NMuZvAs6shfRjPrl0GJp5M5GxlOWa8p
YX5uNGsYFdMe7a9qk22iwA==
`protect END_PROTECTED
