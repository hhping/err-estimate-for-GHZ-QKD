`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vk6PdqbTaQT7yCTXuLOqtcwWX7L8+t/pAJvek1fRVMgkRYRkKWIKwJ2YWBUXVcJE
HcLSjwfIy4aMYsVRGHaIstUbeEkFoW9igTDcN4Nw1KJhadhxqoyEZmrBWwcOzwJf
BKiQv42SP0nnlC4krWEFeR1MOA7myC22tAlZDPpp7ouZAr/Km9RG5hXc0aXMUOxr
Cdi+0RAqR3ZEmnhBwLmznQHGdXHLvSgj4GaENEq8K9eqGKBGszzDtvK5+LJ7GaIR
1ubPjniIVG2osgJQLkn93E05ym2We1Bv/V1ES6m3Jrgw7OVx6HnQxfr+yAd0vbPN
TncrhW9O/sniG1jzi/3NogEysVxO8x5syGIQ3KbZlVmbjzDAK0DQcz8vDtlUtUna
mSP6i1uQtYMVUIH2/+jUXqudn4bNzSYEpts2lPaLq5rlUyion3RFnsVCZ4wuJCPH
Hlp8sNvlONNQjwibHPRP36xmAs/TBDDBGJaX5jNFhRtfw757Tjy6zkK3FfFPofgx
d8GSNd49zl/T4QdFxoPOFoVkPqe9yj/Cbe5w/y5DEYPldtDFKKBmcAerrIVRY2xG
ib4AL4CXKpteRA7NcXOCacDip3DnVAUn3KSJi/CBi/uXOkFF40xSPMy2eaFXOBVL
3aEj1hDXniKa9IPRB0RN5/A/yI38oz7ZRECr41YZb2KzIQqLyOQiUNxHXz/RTMZj
Y4Fkiy1aP9YRdunFKvf4xdlZ4Xh05vo/PI3yhkU1lpFBgoMRwf7KOk4Fq3IGeHJ7
JYsytd8pyDMMyuD7v1Kb/5hR+eR0yBEMhFSfjRzQL9shLr0jQPMTgMVYVSAEOgI/
unOUa4U4vUl6AATei2LQDYlexCKouIj0/a9sdlik0rVNhHPt0yabiqYlA0HZ5h1d
DAfJjgJCi2pcyVjFSWrX4t8pJBYuwEe2rOAjcVP5kAO6ywR8zwv5PvJhsLyK6j29
nn1MbTBILf4G8XB4mZc7FKU+VMFTaI2DvXIzLw6KQmw1rRX0LnsHSV1P6Fjapzkj
1AFYGdZQ7HaDwbDlV6fL2hkevntNCdsYStp22S2Bn9u8rsX2m2uv1hnLYaXL38zM
DfJ6GYf+AaEUGw+4qUTmk4U4Q2hSkOvT6WJ9u572bpB3ct5WrhkSwOVpou4Vxn0w
uiSAxzKHpY1e3EhoYUKCd78F5jGU+dbV3kRim8RQtJUvZ2PAFr81Lev8U3A8qlKi
A7VkjefGWPDLfL+892tQX26Z/LQqS/xeFbs90rmo5wqS7JBsykU9g9hREctzghJX
fKOLirC7WVepq648t2VbiaZ9ePhd4kqxqlhbs9N++UuNo60lSfDEMhGbDwmrOD/e
0OG6VpHl943FxDVeBnxqQp1bieApU80/lvhILgMrlyMfr0PqUotxDwfJAhlCsc8A
OqukuFKPg8p8HxJuR69ATC4siwH9Q/EWHRjLB5f1ks8pVVEik1Xt1kcy9Syl/v6b
vzIWhhxWefx9MnLrHeKEEcA+4YEZ0ewS1SMrKHoVPqWTNcg/Ne61LD/3+RYAeBoW
eCVEaa8mzkooTZMuyeYtabnPKa2nlKDvdUPKvR81zjnB0QCBNGDq0T38thm7DmH3
nkK8lLATUi5vSE49sAPMoOfFnrAqZBiuaLAbTc0oAl1j8uGOlkJqbk1xEq9bxBnQ
6+RSmL/rXHFGHznmKFAX1gzrY2frR3jGmF+drmEK/UJ5nmiy5jh+ibIuSmsgy34N
MgWcW4qClj1f4tS4+KXMHthh246fDWzFRSOICAcUKpb2ycXIp9M/DLK7RlGNbNS3
cDJ9sR7htR4Kc5E8t7a9pLzEg/sXzoteEKuFLaYzPjC7s/sQL3uGq2GLbnDVaHXr
smZuHnUjF9uwJQwcp2Ou5310rbA7UyQECYX3GJ5KVEe9G3W3dc8ZkKRY99gT+zHH
`protect END_PROTECTED
