`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X6zZdVM5heKwPQ1yjlsJQzrwk9tyzkfV4pxscOHzFUCMOrnag812/+Ki81sloweW
y7E0pSUVZbrc7WSGaf1TW17NEu0zQ7e9Q93Zvmtc5BDpgqRxvUglgDXfzHeK1do5
gOvj5Nw1uOlu/2tVRXoj2QPc8ks9jebpcVPeHg9mXJLjlTp3dHQbWlGfhAR2eAIa
l4/l0d1UIcuba/llgJf+sfbZolXg9jo0ByAVyks7GshmLRgaUgPaafGNwb1v0Ryv
Kd236Dm163wS1hw6vc+eG8gQDnFcYR2F7KClm+6UtmklRMQ23lR4dqilI9rQalUz
zhpklxYWv+9bQydtoxqUXQzPUvVJuO9CoIKQ1E81W0DOwh9qGpkGPltTDC9Igho6
SJxb/ejyqxHOpjFuP9jTBMX5mR1/UPqotAW2OCnNPDTjhi0gtWlpBxd8dMvgkX5v
IPdUCGu847X+0qgy9Oroj4iOjk0qgq/RXgRgZlL+cNrCM45lp6q61zqFpBmP+b+o
bGCNWs4On9KrtxKBPbUmJKeDZC41lyExchxbLNvWJfVWTytQ9AVRBsQnPh4HBLLT
jQ/EAy/T8MqnsWX6g4ru7u4EGpj9KX1rznadYsmd6thqo+t8Snuu/hVVipggx46a
b8ue6zTmZ9aLtTF1UsqpF/Nq18ZSlsK0oHdpupLJ3p1/loo6mfJi6zqAjINvHjhl
3xLToXzq6B1Vs65kI/j5TXiQ2oJcXZHsJfjvZS6+fh6n6rMGIfT8LCzly95cAPGH
Pu+cRet90pS0A6u7Lmv8CcYbCBS1WqJCaM1u+R1C2rIjoOUiriVdB42BDmPWEkCd
EVmbAdm7WCVuFKLYFhwTo8JdigtxUIsnbgGmGayBnkpo6elFT9DUZ8kRjGU6ie5O
cPj8R91LBj8AuB1+wNWsvvailHVxF+CAut+riEWCy48=
`protect END_PROTECTED
