`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Nm+9sn3xKNIJISOCCq737E5PXelnqSfiDkyJJRu/QRr08rPMTH7YEcmNU61SKtC
KMpedBH1Yo63zFP/RAkX//yLopxkAyaEC0+tGsiy1m2eOFkJpzvxXMATji2k5l6V
TOGXz4yG7VSBdCNy8tYkY5wpve7kPogX8v25KRtcQbFPRY2eHbxOADwpPbtFEGx2
5Xx+2GG1A6wJVwyc+xJpocOUWCos9rvIsCPV/usrxhTlLeGstCaehknVtz1gx0Ii
oXU2ThT3GjH45prblONn+W74Hdfc6gx9P/z1w1upy/q6DsRaaSCcf9cBOUAa0VTU
Lx7V8NiMk1u6n8rXG/pfJjVJ9jeOarWToQ4n631adzTCRfhEbPeREh6gD5PvO+K4
3E2Tv1RnDM9ZhJf66evCMx6x4gbjK/5Td6di/g9aO+5mWq09nwQVGw2/SMCSBxOZ
CHg1lyzXHpMTKDPOyNlhX3GzYPKBqd/Ah6PRP1BNelyyghBg2NfDDRpp9L+mbNF+
9M/+4gabTa/xAdqxrO36Kdy1PHlPqhNQSr+g2XXkgcxVHb8hkTPVtVYMmzvU5aF0
iG4KURM3K+p+J63XqAzufgQrKJ9ntL+aht7klETa8ExqLqq+h3w+jp7BHhMDhanF
xBv0bIIUcwAltuKapQlng7vrD46u5QzX8YTJ/GdK0axpjG/2M50MtCMRfbFOB+Pp
WVFRsYIHMNLNLgPnZ8g7w6Wr/0VqdEIbG0HnNJFhZJA1gtEsYrFMNx5L8TAA4Ev7
GgoKHPqegvVphScv7Wix/tDi4bwszBFZZ2tSyuissLWyd7bXxRbY+bOQlhNLENrY
eipEfmz5Rahd/N86nex2WIhaeq+RDqm92W2rUTD64FuFKR6YWGzRU6ozh/fCdPop
T+jOsZJwRwjlZOIuAFUEmv/Gnm9wzSrStBknUDrSkc8FuyuyQZRqHCSUjijeyVww
L2X+mSnruEDf8MZqv45g21XH8HvnB4OZKVGcrT3cAjciD0MSUlUUQDVyIK1TbWiw
8jxF4g5xSsGYMO19OnjqWZkdya2mc120F26F3KS64QhnpFVUOvMFDDQ9oiDcfnar
NqqX+M2M39rA7eNKi7LFG0+T9F2Rz9QQF115RQuMnYxXmZSKSeEH5sMkRCwgfkso
Ic973OUn6aa8vlvzDfursxvAakFFrELuNYvHNVnD3lgnfWVHz7E4ds08IGIOHv+Q
xUmXBw/otw/o7tcBlJKEPkTGQZ2850ttw+xJxxSHUMzwWbtasLm2nd0BLiPSWxt0
5+l9jpNhD9BRgr2ckW30W6cLoa5Sqy9wbTX20VhiyFcFLhooTfOgg7KU/AeuETAu
vfKsCnLstmCspfQAWJCPuTTt+XZZ594d5n6bhQVPP/fiSwpI4wGZhFx3XR73BVL1
vQiSzmfdAAW+4WRktUSgGHHmNovzD08WAwCs9SV/ujkSNaIyMbjpYm2I0RKEouoK
22nqsSzrFMBxi2ytRUW3extPu7ke8nowc/EmWKF+Tk1SsGMi33ldzfHl6TCk6/vg
omHUT56DyTlq1qef60Gu+1/nrawE5HaUdRU4tn1v8yyfxDIxnIa5Q40qUuaIBKH7
aSGEOj3+FonHSl0VxYz3Sl3RfDmQ9/TIT2QyaMR42WVW8pheWnttcZyPVhrRLgLM
1JudJebBco7zCcpcKSxpTX2mLY0LLUUUGd+FydVlrViLY7SRz+J/paSFNww/Cad0
qiFTy5pMf2nlAr5iNCdY0wrewsBFK+Or3l3gw+8edUz6W0E/vIhjzMbm/EMnasxL
9XtQnwQkPTAcKQCcnVPdLvKhFSy9AUUnQ1DtRKnYvuWhEQUlMXa9n8+RRveq+Mxe
K2whpeaxUlynQ2Ghm9t3zrURuuVc1w0xsNUdzjlacHrRWEcNMJTEM++y3MOSvsLP
7e+iMOM4o8t5VGc1h9lz6Q==
`protect END_PROTECTED
