`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+LYM+MXgU8Sj4MEjU4lXgNkDX+oyteDSIRNiQfpDxwyXhjcYLjerGQDLTSN8hYUV
DemR63UHQ50DpXLNjkWqe2w8Cqk4XaJ+P84xp8TthKPro60Ufglc0wtbj3MS9WCv
pDWq3n7j4nMsOtto3v6JghtPYagA76utR2FPB6TDkZVhEnsTHPDmWTjwxXDD8WyW
bIX9eSUKBp6okoQIXuPiKNQ8JH8Bb8uGsCebEwa1aMhZJWSkR29iGq3iNnDBNcYc
7Qn+GuQgFeir0X9g2XXbFtz97yZAaj3HiMmtXPYq+rcTsNS95oeN7iBFKYoIxecp
NMj97We5M5AhN9yKJp5h9AJujseGHmodvvfUoNngQBFJA91jPrOLBRqefeohgmvl
D8nRc7ulOHeARV/HedpDju9g8E9D9qU/wzUhNy/ajbZGrx4hIHsTfTF0HqFsiqH6
9VkzEGqjrZpI31El+JkJ6bc8n/LRF3iOyMACAGDU3E6XycohXWAb5w46zwyN/F7Q
s8soOAQ2MY4eVlDCUIEb2mooCZyOutexRxrO5hZKbyPJuFPtI+HXHjzGFlngITnw
XIHFO/DrBcAd0HOsydA6WTYEUQ48SrpYrFcTaegXJqCcJTCqEAAV7TggvFLiGjh3
sMbvND96kr/hqCigf2SWQwCN74KCjVw4gZ/goLVD3n5XtvdmOSsm/RtiIvKH7ylR
ET67XalinL4Nce047ahlSsuft8rdVmh0macFK86g0EtPBy4v/iKPwjqWscXr3hjd
xCMG+i/LkUqWrzXA+3OdNBFAbZ/zfTSpyZZQpeVHYVWqPLMSoECUlLtPR5Gt5FFp
TAE1C6n3gpF+glYj8aJwgO8s9NgHR5kCsVqPp7PG9/eeikRZaUynkyh66hkvdVMz
CF4VCgU4A4YwUD24IwN5Q+WOH/ZuNUE2b6CTlWnpH/PBYFGA10qpXwaRj91rPYEO
haIAK2srMQGE6Mlk2/EaLuXvuGbCyHnMaAd4YZRdzwFdjnos5e5+wA9WkdZ9pUI7
I6Z1vprr3ORvpBRngJADjXpuUmiozJPj+plvNfYPE/04dkmVJr4EvU0QWzS9IJ21
UzJ/PLue8ciHC2+h5HKT1eCwf7P1FMW7vUXagxS8lSCfoER5CqI+x2GPaXWaFzRI
F7xfklYdaHD8PXPJeTzTfpayn/NFkTc+eSdXKZTlX2WKlfbLZqkqaAl+OFUDhuz4
23MwNSolchhxasPbq/zs7MQkeT1Qrab0h4HZ7sKxXRE4WQ4ur8eqh6dm5Y2V2qzV
LPVliJQE1UaP0T9IP8GIWiP16G7bKL61EV81JKadLHT3A92w7qFFemfDkJ+HMkHM
gMn/FGlJ6WvawccvwHAvXOFerR4WEH2ryVS+draEsWSsYN4025kmje9UunwRvKzC
2Eh990VkjmFzl5ZvvZ+oyGEO/A74580ClpiInPpavaRx0FSnrclN8H9AZV1KQXAO
eL5lnp3FaFp+0wI3UEhn1EAF5XlJmwDIOmqTDcsygmtGWSLZQXxGFsD//ViP1A3A
pKeu6+j1HIsHaFc37QpW0xH6iOO/A8kzZ6vaG8IfrSsIUZgakPHMWZjEtyQ3y+Lj
+nViEJdkwS9ZdfpC1VI9PD7uDjE2wXxuCfNhcOlwsCCfghGfheOOl2GALp+8ncCp
vZZeIVUsN3Pe7m4ypdcX9NwJxbzfw50kjnjJqVxMbMe5IZvrkacHZfHaTOFFGEl6
Z0BOyY8hOePOD4AnCl5iXEzYPPx73jIGm20XriTCuYP4UG7jkMYPjV1VoEztpeTT
izUkIOPYJjIvv/GuVfjxnqsMO8hQcYVduanlWji+w6GaBy27sxPq/7+U7uFgJv50
ZtlWLOt0MQnbnP0Ik9FtT3ZgOwz6u0KTtpF+2GZFjCFWP3sHuEIgkVPA2BQgSfZ7
m5fWtCRRh9q+7l4Yj/BvCw/MCAUCKebUpl3i8WuSPawisMjNqKTSYqV5GqCdrxHU
Dbz6gVw07vR5ihCUOSUu4xmHjFggafJsBGqeeXyZfJJ97Im/a2pvmH/IvGjnkhNf
/SQjJ0o4FbEHX7hfam6XgP7XFTX9+08gC6X9avYjonRLwneob+ex5zHa2B0f5Jh3
+s1+BvUoXK6c7VlZF/qZTXd9IJ5VserNio11yPzO6IV4Yd+xsXw6jK5b/0BEV97e
y7n2chfknBeaAcwIgKBsY+1vlQcPsH5ehwmGABcVw5+QPQrQB++ug3Q6XxHrRR3O
qwLWr9K5UzUcz6Q+PgP+ORDvD7+IasY2T3OpXoIcnFjhz0A5oboN5Evl09q2EnqN
cuQLaIoGyGlcJuSJpjpUzLHnEJ/XK/aI3DYnbEY1JUoR2g3Fr8a3Dgu1BSuNwfQX
vdNJO8QLRtD9A1EtRMSmMlczvdNIA47XRjI8yvxEq6moSPEgDm05PSnhV8Xkp3uh
sppVPfflk3FU/A2tiZ6GqC7S9Qspw8cxuUD0fIhTgQOX9dNEQ6aJuF/QSv1+Bqpt
9xJayVlbA5isvbkcfEmZbu1Grgx5E9H9JiscQ62Yom4N8IGVcFHNpiWsp22AoCfz
j332ZPhKk2HKQxpA5Pr3vAUBUnH+Chy8VEVIHJqO5zJWGZSEWD8FR3AlddMqlWnl
mFyS2JnPWSUTfMeoJtrf09epyKmTi0e0XreH8IhL53FbKGWXzVsTj1HE/zZ1lX4h
+hCOADZR+4H5L67PfXg3rJKkeE3GF/mYc2+MU2JZV96N/hdv984GZh8K3RvL0IoC
ebCMLzCEgxxEpUOFmRr/Jb7kAXnTz3NsHh5EP7wyamWnVNvesPdm0JVSnqH1wO1W
+MiAN7NQkteZCb8Q6VbpwemwQTL/xnjpHmU+XB3yECLpU0wsA90Kyc/RyATk3kF4
L3t7T8UdIcudqjusDnyK8BWGNaYLklqHLwIct58Gk9+z1lAKNpidEhwiI8xQrrCT
JtIg83+rLD6j964GdXid1Pv5FSEtblYc5orlB6jLrOxpUBt63KlBkxZFRQjkdgYU
/yB7PxkJvddtWL9aeVuPunpSxPmwRLaSX03Q/XdnXEWUicLZKAOnX7oiimYVfFac
fdT1JwLYQNxiHhZ9JysQttUyOATkQk3IYA06Aj7FyCFpeRe7WUp0qGIK77BaYGPD
7HLrA+qD+BFDlsIPz4L+pJXAsvg7tVD93JZ2y0nAqeWM4w0S83vbFNWartocLD8w
zkm6+YGbq8mH69/wfQiJY/1yGn2wMghL9wXOH4khedtLWKOs70OP9KdsblnGVOfH
oFuoTlI2hBqvCk0cPWb7GARjeMg9kwA4vp/YyNbUKoySxQ2jIE7RvJmeOc1KRTSi
hntuLNxxa3760MPM8XqdOUYjAKS7De1RTAfKdcWAfpLhL7E4px/uO3AGIczhusOX
sl3JbCtABqnC7AnvoYMLtLdTSeenAKekbRDmPw9a8l+ndfxuAoc5NKcZ/Sr9fa1z
qyeObBv/Fg37ID0duMwQ5D78uG4UmPdmxZm51/T6nvAOo7h+5haYeadllNJ09f9S
1H+u+tJ9XxN8XQ5F9pykk1r/YYDPGSKXoyHRem2fpP0GBUk7RkuHW6JNmtMFPyri
idLNWdzBGNjD88Eu/U6MbEP/Z8cbAncC/s7x4rpqrE7cSkCX+fk4xfWjQ81/I5rP
Xd8ToPMmcvXsdEyS4a7I76nfI4QIQLVm3jLfElkP7ajTpTpqVwJghnRytVn0+a20
UEc7VY6g6RLYYJVsuCfer0ZhWrqWB6iCPtNTiyjznRjGh8B1Mjt1Qf8f0HbFO5JN
yPJhZ/lmCupo/HIiiUawMfnSV8HE2MspOQi9oX51rVCWjSwqIhLXDxcbsQcvPMw5
884J3pasjIbTTowGVKV2fMbJjhYqgBks08IqyK6fsrzmlMQnYyu13R3LtllAHC9l
5QWrR0s/AE3sL6zwfySFQgYncppZsv3LQ9xlgQFKy1uRcPADN+FbcidNMVw3QJWU
tLSlQQdXk4ipQhkY+JLnFPPpnLo2GpfHUHiFC6QPfaQ3Ib7dDZ/l64tpV8D85En3
2arKx3rEAUme+r15gRYV2FO4BoCQ4mE+D7LTHQPV1dMEFVuisLtgyonfMjPYMruj
diyS0WX8l0ryXcDhQ26b+T3lYYYsbb1qGEl8OsIbe5CqECFoAtzxRwcKbL/mE8/7
UOdtlV+puwlfi/xEk+zWQernbPLIGVMq17G6pUndswnKIhln7nAKq7QenaB1kH/u
H9bx1mASm9BdfW4R3COXzSvI+nHdZrw3G9Zf+9WmopYdybLJaMlt99iGhZzQIg5C
2It+aOuJyuDuqoEXd1f36EkwPUmiA4ocdswiPgxGUFC291l1IohG3H7NzhL1xWBN
bKtswLtfYjcttPFeeluctwRMaV1Qu0VyCzTuWYENVGERpKtIPslQUUVkOqDMWACk
wBhwvjt55Add8fcRSOj7pAfLYqx3IJmKAy0NcLT1ardHvlEugYqaMUgLvMI/1K+t
TBGMYvFfMzD7nj/BSCBzudQqOR2wHadh2LdPEV3t9oO+zOhq/6a+s9vq/QxWtc7h
N9ajPBweG+eJRN3mtf6zA/wGv93KApWQ8hdWE/jaovyDqQlRovbLt52jisGXT4kR
dbLqOKQRpS0atwv+RPnXyw+5tihmQ/bSD+dhS5klvpKsp1ds8tcgU4IaMMahMyht
FymwqkxCec3lCruEN/6ttJvhAzOIb9XFJMSW2b/g5z8bEc85li+XhVRgT9NGFbFU
GG+DRARVKuxKOm9wv+U3halfx2y27osA/iDEnHTX+raNhegDFyk35pBZuCewVekI
K4w/P+BYqPVXANS69rvWTMMqn2dajzhRSGUXMHfVWZ97vgWXopaRSjGr64b+nwL4
X4e3As8FuovE1WW1QK4J93m634azXPYN7RqG5pLMRsc+GxJEoM02Lr3BjP/GyA3A
5ApFFIu2MzIeTZialDbho/WrqBgAZZblJmXwKmCxzISg6Bd7jcT6QMiDndaBvwaM
TrihBP5Dcqagr8iOswFpdZUaPAP8ShBrsnWW3kpBRLp+S397oIaLAbYkgT8T8P+F
krhro9HThKEHiWDw2KJ59t/YC82Vxe4pwDzGoQQxOzO38kB2RQRFij0xHxRwkyhG
5Er8DsvPMtKFqdOjofCi+HcptiS1utOex8RdUDW0AuqlCRLCSMWMyLakMmHIOEEm
FZtMRyKO3reID0h1pytFVQz2hRo2zC5unu50CIUshN+swGkUBCNvKIqd9PVMOi9h
tu73jnytphLvtOiuAup7yhd6YD9HyVWcqPsRYYMvkwK+k7+3JqP0df7V7pCmbRaL
BIatbt2j+fOFCmC2JPYKgkG/ZVYlBGpIPG4R/HUXO3bn49wRq9U2k98MZayThqG6
J4fRfJQNFFWymnYdFEKwqqyoP2i+IYo0Rk8uzSlLycwcdF8FrP5ASZPQpE8Q+GPc
UjiKKj7mSEcTH/Pnbpq7h6Kz4+UIgXUs6Z1nuDwk9MfzXDqHfCPLJ2N4M1wvapxM
diZZ8ulPHszVbcUeunQlgvTiqD+rzoOT+B3WjxdJEsp2fw/zIIjUHN56tHbckdvZ
b0A7NsS66KqCcBjSNjKamoCkPEwbNwfhhMb1roEQQ6zgKq48Iz/EsT30If6azEaT
NZjyRSXEgP9mokl0tpqlfqRtvGYzd9jXj5+IvWeMHrD9RFoCS9WairbMIcXzzKeH
Ye0Lz4rJILsoglQF4uXzeUs8Ua1JJ+F8E1NFV3uof4YwkdyeGlneaWTw2zCPi38X
fLio4sUaFUDKkXmTD5GR/jyNGPOI+j5SlhrBGBUoD86ex8kycmecZWAPQjZZ3Jcr
Aqw8YF8WNwjFXcatVlq3Sijjl3cYKDdRk1RM7AZeEHhOJ/dYnvs4IMPaBW8v46hc
mvUNPQrYwxrYdp+r3gVRfIbzaiH0qlzx8Cppq5t6yHhSLtUZU5txVLg1sJ5Z3jRl
wVjdYQBcTaIKU6VlpkEEkKJFLugV0dnYnYcCKRSsgIXlxrM2fSfMVtwB7ji/nstP
j8rRKBBehARbmKnSaAV1Ex+bl024FFNc8yvrT3r5ov21Ba0i624OsxVGizhWqNRP
omLHKjtoME5If1EH1q2uFDg72vCF+AdnlfT+Twp5p7lbO3L6IY+dZNDRAztaPi1P
C95oF99B1jVVnbYywWO+ADtygMOczPRKK2L495iO6zvXTGjl/RUCwp9tpp9vIUII
o7H0B86CDGQgZx27s97hR6L13Udz4MybisP/h4YQne3gny5vXqgQ3cTwxYnmb944
fXT5ieo1Yp9beklAp7Ukq5pkTywk01gWETwRi615Jy6sHv6fJLtUoMUdLsRi6Yw6
rbIEPIGz5Yc29rPYdUgEUT/fXc8ggRWWD6oB67EeoIRGfMddkr9Dv0FAxnRVSfRH
5XXC0yTTP9RMxigPEP8SMfM7DO+gvsBv1orm7kVTKQ7bvk1bLpz63+RzxIuZW4Ze
uyBnyTtKXj9irTSFN7frqgUB/NbLPl2Rl/tIyLULAIpvgr3HtDGd8k2X5DG8lN07
cSYvdPXhOcmT0DUuffFQRMi5AEyIeI7TX+WtaPI42MIhWVyLgYiI6PMX4eow3LqM
sp3o6aFK9KlNoq/JgyfuBjbs6JG8KWkyzbKpcuR1plasfABu1QzapGjlYRT/CDdh
Y+gN/jT6gljV6NXkp+BMO3374HHh9ZfxbAWZFYSvK5VgM1x/prJ2e+/Zt/22JW6s
WoVqvGhjErUKlqItF9+7KhdYxOlwpzCMDpLA2Usm7fQz/8zciLXVst07GDTWJlmB
3E0nYQckjzHQpmIeUieSgB4A4AYbsE4bX8mzCdXEsrak3F7i1MejnJwqRhbjrewo
hUpCVFcpr062xDCrbr62uEAzmwqD8gR1nsxDTWP0TRRCkd9w24qJEl4UB0xCZTkp
GTg/Tf5BZNjRm60LrXv3RrkMYE1/CBh5GVRbObPN218wR9d7rQdK++GHyP3W306n
QQzqqxl8GnrNmHX/oB4L90Jbe4xP7Bk4h4mMuF4JBe8JwtVmYCxXALvRdLPGGt83
o5jyR8s2KNTnNMV7GpT5+ur8WoBqbkZ8LWqtWBSGb9cw1GNiHrhFzYbL4NC0rWH7
eXvKhH662aFIZ0NrFTqSLGjLkWzxCcQc9hFGGn5pf+Z+iARs7iIP6mOa0UwZ2xKx
NOXujSTrx923uzmKtyQTKmZguabvuvS1ZcBB0wi5JVBXqhhJVS/m8rpTkzkwOKZc
liGo/W+UjA7H9buurJDa6DkXAjqaV4qvtTnV5gHcJJp4yYSeUm9qjY5LYSogko/O
O/VtW+cJj4PYsUNIdKCxclP9rlTgbOCunjdGAgK4xlbEgDJ4aHUyoQqISKIk3bvJ
CHVIDjsJxzrDV8vmvkrQxyL59jKG9yd2Fnwh4xTzsTCRLkeEMgeFixrJJ5+wICR8
GFoChN5LyTAyE7ZyJVVafzotMR7OqDhEwVrjjjEp3j1XbBV81FJaPsX/aXAuPTlg
jLuQ/eVpTe+OWG8Z27qlDBr7c6DZQ4ZGy9AvRVtvz4TjjvQojToxBsROtAe5+TPk
eV/ZCDBqHUA4qvTetOywNqjp9ZzerEr/dUiitmtkB/KXqeUmsYINjXJf0tDMx7/2
C92YbPUm212HJdfk9UfdK8jR4D+YonunyeXTTtaXfGJns0vi38fdr96bL9u3ypB2
brWpekxos6cRce0aCylRMVueYXSviQoLFFQuzUEBudpemdsIg59gy1yFvjlcII7d
KIbdjd704wlrs9qoojC+lpKys4w7hn+vw0YkQb4h8yrZGF/FXVThUgyHbUHsj5lq
PhBlbnJ036c9FmYkVJW7Ktavt2/Lo6bqD+2/Q2qz2fztv01GKMxzyT2w0jXsFRQ7
AR9zdx/4Tb+KjED5PqxpBJMVGPj+TTjk2DpDpkB/I/qk0vFUdMt7SCx5YmQey8A0
2SOlQj8rPbnFhT8WMTGZG6CrgRyDLJVDN2X/+zfwxOj0lJeYsnT4LyzB1ZaLGb7Q
jPjEOsRIS1hDKD1vGra53jA03xJ2Am9UbDTYYFPz1b0tiC3mVyPigkdqjDIE2i67
NCpGdLzL40KpTZ+057FgmvfcXXOLLiv1j29IxPDiKD34oAoizNCyPqyE4G5ZZ2fh
X1tGusgSoA0vbA1wDyVnt2VKg2IXi4C1bmqGOh9JXQVuSQua3kOHS+tTCUIHnFio
MDW71JLIv0e1oX/pbAYFIN4x+R9X8+JyxJvwMOP8LOiA1VfbDA963CKkCc7bVGWi
yiNaQQN5VQst2yNCe3fN2JLX1rx9IPzZZJ1f+UJ9PZAVDsSarN4fxDUCaULaBQGK
+d9Hfn7vz0XwKcmNEC1YiyKC5OFBrQTKPmFtg8XftLS1Vx6F/02foa07PWTCuAKQ
QUIBomaAMRJNbaM5pVnjXqac5Jsk520LJB2QGwO2+Lpk8g0n7UC2Ye9SblR3v3az
5W17BHZZpqQDBEppixmB9UjF5FrbMfSd23lpVgJdIuxFecmD6B7TAarc4/nNdJ14
9toXhhR8pVbbb4ijnWfW78j4A6qXBgVN6yBT4H0wygL3uESupr7D0kycc8xWtg/t
M6oZREDl2iCKvSoy68nFmsP3moKP0J9fquW2972+vSPO6yaReo9k7YJHVdR0BUqJ
QasprN5MyTyeu7j+1g3vodDmD7p6DFvAS+9Eu0AbtNt4VgDSjYkYWbBt7A86uFrd
BNIOM176GvooLkx3+M/9zszr1eAUwKMupanAyCr/AOP9hX3DGxwUuiKTxbmHcQJB
T1iUrgREiDnET5P8YQFirFB2Two8n9a2A+btMNYeR4VuZ/8aa7fPcfMDBEezoi8f
/S3holVCax3+9p+OfT3/O2ChdyfEkWzD01YiY2sGkC3CWXDiDBVemXVITYQnMddc
BwGWQKkB1pqMetkz/HVY2+q2YKkYY5EXxoiVNmffFn9xy1asMMcMiRVEEbcVFhpV
sUKjRJQBYDmQkxekL8ywNGTHUUUXX6bg/HfjAwi6Bgg7arTZdPiw248abMWEooDj
jDll6RQ32SVHUHOhTvyeWXmkpCqB+HwiXk6D8npVzbWJyc1WAKNM81Ti37ANGH3P
P7SAp4Wny/g6w8irwlv72G+pbtpAN6cUGXT6Y4WgCaV4fddX/tMliEGYs5GD+Axe
nyHSILe7XV13y6jSm4yN6XLxIoQLmriw+nD3rUQPeMRD2HpYeR8Q/W4ox9AprDzn
C1PgfX5d6VBDU9CgcECZfgDn4tnOTDGReXjQwb67XNt3/O6/ZL/ZmTPbUMqgb+4W
4CPOk5QRB85mBnIC/quvH4mYdEujV46ZhHe86mtX4fEetNfrcv0cFiqHqdjMRfa5
sJVMVoMHcttPPjoMp58pDmmjFtp+t8562Dyzzykg9r5t8rh9GcoGrOV1vj6Of1fS
9Yw8DWunRQLgbWQG4zlXE/zSeUVPwG8Ac+zMD3qMVxQmBrKzop2jPR+uxC6ljQGb
/bPZ0HH5NVf9kizEdNk99YJjMT2Z9tz/Zbnhhvn4SzvHZrfCL3pYMGHr5qwsDhCP
ZtJVj2V1hgw5Hui2ghuM+fa0h1Zd/wk5XpW8790K0TFE9pOBcoaCtsRLOzBGiy1y
VzzFz2wU0MoEsCs0D1IB3l5E/dzgefFRDISCrrV2z07JVJOgohFB78eP+///jElx
SHhjxABe6WNi2k2EeKBbPCbZSQuv5b8O84r+sCIWYjBzYfuLFf4tQZMTJyeAZhND
wPWngXKgzZ0Wvi1hIqB7UuzcawfPDio//fSko4mXRQWbMSv51BHrOOL6A9vvMJF+
0GsOuviSpJUMRxQ1URZp1IKSoiXTw0sWOf8CRbObF49yd7teq72uJePzf6vAE6dI
gaJ0dmrq2pNpbblUnpQeZCoGj1od85uOxaDqRivVEiBtDOXjvq4rqTD1sL0lv/zM
KLeRyykt2Njkn80pVFDbGR3TOu4Q3oYRJlAClV5cU39W0gfLBrLx6958N3GKCgHi
2X+xOewdq/PsN9gbOdX4Ay84gAxg6EJgDH3PCtmc3jqf2GUhJYyNq3fzJEw6oJJC
j5HqiKEsxtVatAm1783X1/+hkA7+yRzpwwIkuetHgSiJF8XjmTFkz+Ede62AXK9F
7kmANDKAr7tfcrxPWOfgv0EZcUaCJqr0lzJ1Aien9OHuK5Xa9kOAi4rzZyTTlbsG
AwpRigFsxxr3AFH9Rr7RBCJkJG1kPOW/8G/pSvr/qgVDmRzF+s5tINa32WQ4/gVs
y+G5PSnEuvY2ExQr+11R1htXC/WmumaCCM88p7Y/izGOflU65xvrLmmwCLCg66wt
yck9Js8f49V3Zp7m1jbEvBeTejletBXyQMzMk2oO+SoK1OMyk9TiXYM0INIdFb9t
TISEMkYivkQuRVE7kxfvk18tQwr+SxFRU5BjIK7qrdtzH2WE9P9hs/r9kT5LRBUk
UYUWbptWsv1ppnNk16V5qPU4w3SWOa/mh37HYujK6GKohnLaya6L3FTJS38Vnv5y
/cHp3XfErTwVplN8V3E57dqXNBZUWr8kQU7POIA1ELeDtnGYr85oEeN7USjVkbbu
7AkZt2xbsSSdcD/mIkDtsfEG5HmXDwooGDmuiRR+M6z1zTAqm0IxyNULMdfpHo3u
E6iI6eKFntqmxPR9S5WdF4xD15jTrO9IyY/wch0PmkJvIbjFMYclEb3K5aVTiO/Z
GzHMZ0gKAKd2p90HMnOHAiu5W8/iIfyPmG3TOnXNkO8t11wfB8JKGtmJk5lHN1IL
oCHNiLX6zA3YFi9YnuOLVZSiMT2OR8hk5g/SRoUmnEvpfbr+HNq4wF2IjScVqrim
bmy3Xnru6Fyc9Y071z6xM5omqB6dVDy4jSxD7g9VZ6w+UurLrDSMnSFHyirt1ucX
/mWxtwlDlAz0LlWuarUXNgFXJpn4bVbETCB0LTF9Moh+ZrazvJEz4iSQhhZxgKY9
4/qRJ3KeSSskc6gHdxrfDgSefLO24BIvO3zVMTfbCs+BssmTyhOCf4YmtET4+GyF
XYKhL/iYSPB5YeEfv7DOzvCpp+anY5gS8CD8Xc9wtmKbV0458ME959SrpD/lABjs
wlz41fpMJirTmjjJcvv0+jXWgGFJqSUuNY/Aku7aqeiQqmXwxZ8JBcJQ1HnxR/Z7
5TeSADjeVQYCvGvjd8Rs838y5/2AKepuqdWVec0rGGOXs+85Uw/CIuedwcpp9k9w
2PciPFwGtoa4Z2d5NsHodj6HQNBb3ZnCqcnqL+Y2IkCwNSMKTYCDwVAVJshQHbO8
+AvIylOKKVME2pEG/doWpw4/5JDFPWb/QJKIkNUwCX0bhiQlZQ9TLVElTtB2Xi+m
CK7p5o6j63zitLM5EWSDR2CUxH+m2opWLsf+bBAsTng3TRBo24Fo5EZEx1zLveRk
rgUzySdiJvfk4NtN09HSdZ62UJqueL4g8S1Z4zQ7che6p7KAix05m9LXZqRix4oc
ydDQVVPAtzc5ZAdE0a95KWztNrcpYYGlxA7O7gB+7/O4uqfqPhbMBKDEJ6H2x0jL
TZActoW3I9UueKbof9PfXD7a2PQZap7pIXRK/eZ/AGOoFnZS2kN5m83GNaUnwQ5q
fe92L3+WmOmeckhv2eP4ir9vh1Kac5sb9WOr+sltajbzKYMm8WZk8mP3OhbEtt3u
W3ZPARBwHwBPlpz0hPVDuZEtDp7hbHxZw2OyBAe4G15+EDELQhETGrWHmB6oJuOg
XGueGg+MIj4cf2s8TQjvgNdCfMYlE4Uzv4UwOdKUD1zl2nMviWZrOwbu+RIftZc2
73rXzSsZLO0OB89Jr47SI5n+ov0hlmKhPZUm3UKvquQm9lETASrVaoTrqErgpXMy
d9D0GDKXus7s5Z7rF5fg/U7fSMatLpaddXw+AxtGpdMTw4v4LzDJqDUb6KIwGaOn
HjwQIo+U730HxRR1hYaHP5hW5MHVlUIS5X88zsQJHJ8diXnGawLzroj5EoxEZWyF
w54c5L3MysTW9+xDgWW97zq/GtaL9a8vnj93avsVNeTgV6t4skOqdEA60csIoMXM
KkbPsx9ph8EGcGjCcGPxsRy42ssqTP+1afU5f4jFV9yxXx2hkW9QZmKheCf3VIOT
qfFS1tLLq1X1d20EC0h99R2F78WHgAf9XsYNv4bNJWHOIKboNkXvn+9IX0tiLfcz
Ht3T004Ce+dUCH2Ifw7fQBSihBTHPpjy5mn0ir4O3oPQEX9QTy24Nss7JGUUt1Bg
Yupc3S+Kb9HbGKdF4H34kT5WqkvIV8aFSnXCs21WOJ8u4ysPaD1QQ0i+WWchs77B
+O7U/gzCCBdCIakdbUrYlzQqMndxj1HLYHm34Nx8eKR7JhFYf0oylmiiCGrMhRjh
hnHqgsd87gCB/nywFXiQRoXuWpHdvRIj3lVbYiQeTVXybPeNs3ArGSsNkgeRXzEG
nHpZ/rwKNf3AQ88RM68iccOY2cKNeYezx6ni84BJL+zP3jD18qrlm68YIOVVTwa6
NtZfY8bp8Kd0Gr3cJNvX/wWtBO4XtqcxSGJqxR119URQbYP7dnIKj0LuFGFWzrUt
aN+FYEthE2a6IuNr0gRl/mOkAM8rezbJmu3jGsGgYdcLMNEpA0v0BgIt+NiWWJiM
FEwZddje/EfLrGfV8Nt8D7q9GRIDo0qoD/MUl0Q8IFdGqw0d+sYXpq10s80V/ReA
XZJWxKuMnTVzxTL/wJkxL1aai93/HJ4EZzgSrzEdip/CukmnlyMpfIgqCadNIHx2
nYtyDjrrPon4G3p32Gmd37JKMd1FLDwQmsE5R7PD5AnmbHD8LwESlCdJep/ykz/p
Ca8fNQKDEp0aTKCCPzhWnhQio221VotzXBoqFFHE5xZKvWqL57Zgp7yikG2IU/j1
lxoN54tdTrkdV/ruBv+YMGcR5eLSqQz+beNVkXC2PQlj2IQTeV3QuG4aMKPodBZP
nOPOPLGdTBD10/yn/K4JNn7xXxv2wqYue5duHEflBAFvnVCTcJTtTRLZAqc+1ouU
jC/YQV5pWiQzxoIPus0Dmj/+G0JwD8eOGJxXVCn9E1Qw0MDNsmkfeetg0eOUJVJQ
LWKGSCafl2LlTBQRsc1sPGsJhIFRKmfSOy53kZQW8uU7uZsG+WLiCB9nyyiwattn
CUP3fMN0Htt8EZra1hVvDpd5lYR4dcEhfYSBn84q3N+oSqu3AgvTxGAZLBSKk+Nv
v/GUitQ72XmgxLgb94nFAMBo0IsvAxxDf10qaPKJMf3hcFl8sYs0VIIZP2oEpRxU
eiIHFZLPhNZMq1tC7Q0l7SUkwg0JrEhQMWRGst637bdpbLIROwCJXyTM4xvgCjPi
u+tQjrGYhdrZ+m0lGcXlkRqLaHscyeQsVgvy3mPp+oC/udQyjl8qF0SgWCWIKW8l
YsSgUxHXaFalSIVFPCHxs1QhCczwTbwVG/vpg9imClO+YxtSiTUf9pomKS8gL11W
gLL4QUpV1uEe4y+gaK+HPH6/Q5NaeKWU6ij5Gt9BlX5NUwVIOdR2IjJ+Nj6jmNPS
rbBJas6/Rt+2olpnxbHUBoVHWto/BiXeocSrDrfazFdldJilHgJXZDN7ZtHcZ5Jq
24XGqFGgLUu3ftMF6a0x5DSt/dUBW4aqfL5khf0rb+nf0XB8IOHp3R9l3KuVQfDz
ZXZzVjnH45hTCV3JwBh5frpah4FbhaV8CwfvuccoQhQLlWgLNCXpR67PJe6fXkh/
ANyC6koHiNLVy7lzJ+VnOzgV58ds4W6diHmmAM4ZH28We9v4pI2cYM73uM00y/o+
d2wFvJPJSCHdoQq/PZErrisFjeo7eM72qsDp8EIGZF7nEoEnrtCeTbie8a287+ar
ZMShOxPH2CTbzwiNExUe0Z0DhC7+zIddyT5IXUfZIonSrB2X7Nn3K/y9otxEKIBU
GRX4wB+c52G4tYyJtsVfqODOC/njfT5f4HKyJmti7Ks4Ba3onxLPJd99FDpSqMHv
+cGAncBA5U4YmjufYbTeHeVFEbE7Kp9qyM2R8POqguZbtpqLmi51rudSdo8oxwJ+
Omb+xC27Ln2aDuTvIHRG0N3L/L9CsrgEOEpqrotVjRpkIAInk8/SdIzbSAaZ1JKD
vkKmg2mWy6jZ2vf/TEmUV1OZnMY/QemXMRS/s/cPIs2RNL306YksFg01rGtadCg/
QJh4QYcXugZ5zEG4rWtWG7YPp5B0zYACYFRfKXxVvcqrf2VsLSbrkcRAWqVN7G14
5iSPLU0GULTjDm24y/9gWimg7zF7Y8eoNNTM5UibOfchIJye2mNkza1AyTkdrpzx
El6cdBmY7+G7i5swap488fbMdzlrInQIlP9/fng7CQ6Brb7bk9I9+DymztHcFBgd
CnMTb0q5sF7DpRL2WiksuPSLVS0WnNRzL8MlGPMniGbgZyoA5EFCMwxCC5u9kixX
b4j1tsSPUkbVoNVBUH/qCGZ1zL8+G5/qaHVR+nDArvJQ8WRNdOQtoRfmTWEAo2EZ
ZOxxtLX7g6gQrW3hxQOsal3dF3JZ2nM30NssPA98fDF6PQwappQZwt2DjS29+Rqg
TYNSSkryEXhMxjjxL3EaSn66m8MHGnoJOEQFYQdEv9hIlYb7QMeDS7OWN35JMBVV
pcXZbSE0xxIL+8Bo9EuIV8ABWXwFvKvq60BrToRT3J+EveNtVWad3S4PsKFbtLJm
cj3tqDoI5C6JxcghXQ0q0HGFNTGngYv6fL22CSltL62+DIIHXaescmAGwsmlc8Ns
D0bt7K3S1o+7dIaSZcci8/LtC7uCr1X7DPjjPdDikMweVDpJ0coVQXOzvEJx2QVu
fdCzzp76as2Y5CH7EuNfU+49SkBwq2ZZOgLo+x5Qnj9qbumVmMuBLl5Q5YCe9oex
LAgZyYMOJIpmDUhEKuo/qnLYDDao9a5peuFkVFrd/HkZjXoHohy7DzamN6dofyzE
aHm+VojSt1MWpub8ZpXxo5D3HwyfKaTaCz+wCtUQqjhKAooGFhuBpEgFD4k80yXa
dZlumH3aEB3QtuOHgl+TJc1eVLUJkIDDrCRQU+w8li1H5oxVkEomElkVfWHFQAIl
JloKL/XRak2kvRg9L5dRiWX1lMq/RwnJKurn3V08q4ZWfM7oob1+10t5fk3a1TLH
A0r7xqt99VM4kO17uRBbHoj1KnllOgi/GMuVHRmxQNWilGiLhehxg55TDJd9khbr
e9jjK4N7mgqaH8lVWaPuY+rz/FrgYRKbcqY2vyAkKo3EFDe9P7rOtlDp5GoUBi+A
bI2hdxOmIeVto8/AkvuBdCKGHMkCsKHReTpzcuMLreRMODExygqeCX7mdnkEoI80
wCyFuD7wXkOgMzQ66Mnas5yNmywpi5nnQTR26D0LO+qGMn/hEZ+FWvO8wOXDhWkf
3OSwkSAPw2L53VNKiUxhl7VSgROuRSPr3b7gTh+XK3OK+yAs79nQRC6cdqwVvdcI
Q4eN0AC+r/93Ee5bLrZeT8CnVWowLMMOJNC2WKpMONCCVIS0jRnqHJW7ZhfzTLXy
8NBONiSWCV3RPzS6wPFCItmA6iVu3TzfyXVfEslT87iqGk0oa935y52cxYVT6iGn
VLvaSCvwj5AZykNKDfMYhgnPrAJw/kKfR0yB+DZM7RQJRbUdtRFnOEaaUVGaJme/
FqTuWjnpWVRs4EzI8/vB8vPuDm82iA7pIVOdWSmr5ePCDYaCxAMLSDpMol45ovSL
8q/ExT0rnj4JF3YZZrHekWU2BKFpdG8AvNmut/QI9qd+f6G65+lxnBO1yUyiEYZ9
WNdjFBVvF6DQWovDsfdZ0OWu6QOHYZWgyARnUIBMmfGXfQHksdef+pCos4aWfA6x
4WfChmOCmcNaFdJDn8NyzdhCRrQaGjFrMW5wujpyPDgLn2k4nx7ciZAS54nUO/cU
02EFl/4loPVrDI2XljrwKRBSIN9LQKNCFvHym8U9wc+FjLoLQrPiSXPv933ph3Pw
qP1GziA4V6PZleN8Te0AsILLnPjfGHwRcQTJPG4aokD35CUJsBdSl3nwZprhkfU0
eALuJwnOkMEUItSbv4RqiFU50CwcQo0JO3rfNPQkueSEoNmtUfW8TTTNla3mpCH0
BjYzmsfyR+BtvYQrL0CwcEcQnqFSp6C0DjdfavY3N3ckWIgVG/o3HYApsxWnZR07
69ulxhAM6nzMiS/tQdt8hCWDHZ26Y3PPlbYRL+XQDmuDUKA9YPgxqU5ja/AndpTB
Q3NOrKHsFFy2YA5lVhACAzM7XtoDcTmU/s9RQNYx02cxJ+50yLoBjvME45dEORk4
tS2Rnj42/ENs1KoDeqgThejFl+cV3KeODn6oUdwAIdJFJEQu9eBwhTpNPBvQeukO
IHHZ2rlNxMicmxA6ef5LMhCq3Mpnm1GmikyAgzm1QA+BkkpjxI6oEYf1JJ9ev271
glHbLbxLo0EVo0vopNSEy53jTwR1sXuDPNtvWTRroI2ua0EhbcZeHIYOJy3vGogw
a3W1dMaOz/plQU55LywVBzb2ZdnVaBIlZ+6ErQ/9TiK5bgpypffHMjcEKsZ2SBlS
cuGQnyV8m7bNhOmQIaB4QU4QUp6lF+VSGlwh71TEeaZkpf4h1lKuJynbZDR1b54O
BK8mLMCnn9FAJ3eGIKu4TP6kuOr+LV8TpaZ9C6KavZ98yS+MshhY967lQ3qy+mQD
XB/uihTnmMD292useAbHX/Um38dfE4trI+3sXizaOhKIVhwmqQLaqBY1WehZ6WQK
iUSM+l7rI0mRyhZ60D/CGjZvc2Pwl23pEvb9SFhkUT38+CiyCjI4zs1Do5XdNQhZ
b3xqSm0mTAARg0OTZSrx3dAyBJ7Hpvzkw4sJca51PQ0AiC6azOlSNfyoTLDPYdgm
ck6rmx0iNBlUYj2Kiqtlh9qxGUzcy2pI7xmdM1FbC3LPHXY1NxgibW3RnkdKJqD6
dHcXnNn+pokyN4HfrmSu7SMo4IuY65kZtYDYKzPSXAFXdPzWum1wIatycNdIvdSs
pL0dbFUUGo/kKfMflVKi3+WpB0CbOP2jxXv/N11J5GICDQufshRKJAqlmhcljEZO
0G7DSxX+sn0z7DE8RSrR85B2GHN+obZlvZK7QGUqhHCEiriT3PTX2iSDl5EMWu4v
eTPA0WTzrY7Nx1NrCusUrVsO9A4cAMbLeduHZXIqF+WhRln32wlVXxyDKeP/mErf
NO0lVxJhE1E+mYz2c9MA13eXqBywj5V97aonM4KXB7IQt5U+18+9znLgHYIxZ61+
Z3tS4RX8VJWgayNdB5RUA//wLIH6hdpPgJ3ptgHT0EBhV+B77O+HbRFBrDP0WGQ/
f9KhCLfFv+Ka5TeevlHuDF3EPYht8/dGZGyeUeVqT6A5Rd534spf8jZ9WKZaNzTg
kChmaAQmpB7djK4KyvBaX+YLc0fTbs41G34g6709PMUXHzUGYMFn0zCi7nm7/S/j
E8BUqhdrmXrlbAKmNy9doErx1vHmnoXMCVVPDfCwANwPZLbq3Gn+6WKM7Y8gd6pI
OVexDrdKqhx6/NlRh9YMaKErgRSOkZhI95EoiODaQB9/Xe+NbdSf1M/tz9/I9pog
HyAUtwOrzf+drkdW5lj8tobtRdyEGMvlQW13Y70iPzUscqYPJegTft028I907pqk
0QoAncwb0n3V5uBmxtwSO8NOl5aijdBjlQ80WDYjhQKjA1gT8JRMI1kFP28zOgSk
P3eLKrSK1yCN+43jpb7um+J+W8HV5gB94F3p+WvTCf0PCpuHDFfJeY6p1C1f2bTx
VDJfKEZDpgZotKaVTrRgWWmHLXg+MJp0Ef695D/sAotgG+HbKbVbtANASybZHVeY
Jgdy28GdjKTzesUxgGFd8Pd9qVgTcEjSo7Znk1YzwS6LtEHLSuRZK4OmYw3qVsmN
7TV09c1sMYPdnPN5fel5VWNhQqa6dzz9QQkkhx/+9wvoE6EC96HBDuU3YLqHhL7c
MUIpPwS3KroZLGzYIL0dbhzWu4TAVdJDocIwpuJ4u+71+an6yn02cpSkduLFealJ
uGhES1ayoBf+qE4742L/y1zfU+uNyMb/y+cqDIGFHSi5tz4Jw79T6pMIa0/E04oN
uKxSuS0CdfawE4biR2O6jpRq5CjmOw/Yy3ovICuXpUUFLxvnc8Zu+35XX4mRaUXB
5SGOj2vsQSL/7NRLJlXRz5OFjIPJ8LndUg1d6Cm+PTMyXDbWXDjNR+10FK8lc/CZ
LB/qZa5QdXDvzaKQ4AdBklK/KGz1DR7/uekjCC9BPGW0S0iZ7sUTUkhhol3155yO
jlgoGVdlUi9DDChflwXv7aEcs68ljykQMKUuziq2X12pFxK1dsQo5iJ050X+5Aj/
iucz8eisCj0dNkN3pisI/qbZfHOLyv5Q8s+IqbxBg4QcsUAX2DimeKgLKZVBP1fd
76UILlPU7K+yoqrMTesHR3LBeZjJzt94I3HWDzI60itqMwIve3N5OHeLmIunm+1d
wN97oT7er9YmjM1ilgK+aFJ7Oj21TwYVjL/BOzDqt2BjQHuoxaJs44MJyqbEsUc9
158cLkdMlTN22Fjwp4IP+64aJ1Vr2l6+58ynpWPFDXoM7XzqlFONfKTNmQgBwSUM
LNwoEB2hcRJQB9G3yaHEkwLsFOsKJo5VXqrg0W11FPMcfSJLoBZ/EcDLVum5cMaj
inKIF6Lsb4VXdwwrkUenutoUGi/9pAru224MOrZ9TkEH+p1cl9ovTdzfKF+bRZNM
WgpfFKuFt57MgmmoC/cZC4RI6oY9v2eBTueHOMU3ZmmoKkWI0ZxPH2Pk1JQTAEAD
+tUJvhYdk8fgNkPjxCj2ZHwdeGYxEG6t/3n7KhvY6Ch/eLprm9HXmfV7WSo1WVSO
i+azey5KZNYR9LohTbDTWvJCmO/ndxX2Lr69B50hlA/rWHg/rhAMSwKY/Gbf55lP
ZOrJaSR1q8Ia5v4KVinmG835ko1/5pBy8vTnEJP/d8yYWsuTltt7ojy/SdIoZNuw
1Bjqa6yBrsDYeb4kTlAh5zlVmUJ+oyd2ayI1Kh7CU4Wv9jZECyNwc3UGTFLiqLnR
g/hyL3pKmt0UwUxbqqMwvbbMny9bHgWmA0KsBx0rUcbup/q7hs1bEbkEnfyaJVW9
C3P5y8bwp4jte2TOKlwhO5eKW8ibx/2iuDyKzCFq26oZuicG8n++8Hx6O1MNZM8k
DVZ35MeB/FmpGUxTjyj5HkmNU/8k19ScBZ9cZ3MT7GeklrR6h1l58ztzZPSXutqE
gsPWX1Eojc7XlC3uw94wrX3u2WlEU5zNaIgSYnZt9EPFkkWf3ELv7wd9hZYcZ0yh
HD6ztEm8o4qivxFbv9j3/nScZt1UjOR/EAaZsjSXv3T99BZJH7yujDRMz/fxB+sY
EFYR5iVRnmrhvvldsiV8iLUrNR7z1z1eQcMaAbS0AqrR1UFytjw0DjIxWOyKqqQe
mCyE5EdbR8LT1I7ZtcivX0SdRU90JMqjV/S/72vMKldBrNmNw4irIl/OBO2Tv9c3
XvnfjxHa1Xwc2S0psO1aSJBece2s7pf2cOeqrs0AcMELi4gxhL/+KQwrlQ+972QD
HBSUcbcwHhZr3cGaIKT3u6AN4gviOHldV3Nf4wGn3fi3g17IxQ/phO9B4VTzQDSZ
wkQG6VKy0jGMnNZZfxcUDcmkN697uOyoBQwKejxPkaAdUKrAgVeOC0buEz43JB5l
0c/P7doNAX2Ill8wK2dK/yZMM8n1QAG+hww5r0zBx/g9G2EPs+zKmd446tJcnMIS
t3yBtiT9Nw7MEfIrYRjx1zJg61fZf0IiMr17p1nwCS7rWdcLoOxReUR1tzvuPws8
zL6v8w1WjsHyoAkZ2wFvGTM71L4Phl7tBjOt3KZf15dL/vjzzIqe1/uHajC7NLyn
rhNfbQO+QEzfhJwFDdL5Sc0v3tSF4JYxu1y+E0AnYOnrldb3LNrCeVoipfwqViwU
ln4wymh0sY3l81IfD88LdePnKWRURq3xW7JkxfoiWilx0+nHphxDojtU2uExjTx5
xeIrnskF3IG4iK1hGYRKxGRgzCuWrwGdvLA6pTFy+Ul/OyqHgurW6A8NjLRqFhRj
8xSOA5ia1Vr/3vNnazqK8CpCQn394P+FeGv/IYpAv2h++0deyPvmHlcGlgbIhyFQ
KbL2f2kWla2sh+VqfDXup/b+7AQlyBumWoBW6Yz7U6hT0TONric3HQAAckqfAJNP
2g+rfcP9QeeuEvWHEMVh4md4iQv+pNoMRd0sLeBOdNybnwstaNR/Q97FhG689KLc
vuHZIvA94TRnc2IPL+Xk4s7i8iW0ki3y9ItVWNV3JXs47xjj9m+muu2XyG/as3uM
NuFHS0YBEVWYLUGcQBIFfxxdUJkKBm1osC1PeDsDWXHHArKLLbNtZjaES2JrI4P5
5G0fP8X5CG2v3tpoiTcA+91tTxlEDKmbhacidm33vQSFCdOKBDZIFa0HmCUZfgqe
ojNtBkCHMAuP05v5MQW9nMzADtteQw8uRFd+E7pFtqNPD6y3JTBHkpB9cxwe/W9E
6TNsCQL7V0QRiO3uQy/HUbzZdDHLUUu5psa75QerliRE+Pmw0OLO/cqsXuArOJ1o
+kjJ+kOKCkn1o44yC4ySsoKlq50GYB7Cq/+T2gQMiKjeLqGXafLpRXqX0Rp1VJ9Q
fnA/TJnAqoiZyUsgtREg0KXt/7I/SBwqj4/Ea8Kkg5l6JxdKOJUYZhVirs12Km15
0uKWWMCPHim4KnrR3QpvhdTm7IvDBsAXAHLTTwZKfbbtyLpYa+iTk1N8AwpVd8Da
nNrsk6x4hCI2oxVJgmLIrlaGqnCbWBnSTyyG/If9PxlC0aeRJf01C8C3Jvo68xR0
2RJIVADziuKUCn7eaP8yoXupGBiP/zkojlBJc+CowBSAJP5dq5QETumVQxguP8u3
Xqng/E3WlJ6kak/iVWUSWSchSGFOXL41lnxxDOQryoYGn29bzZtMsuB7F1XC/+5m
G4e9TvvIU8rKMLVGRd9fBb3xKNRhhG6tM5oLFUlg4h0H8ssYW4xdqpawayV77ZJ0
TAkJHjN/A8Bij0b+sT2h5gIykBlMomIYGxuJwHrMqZr3o1uEVBRuZ7AINUOP4fbK
hQl2ysZ/WtGzXvrRQ/Uf708OAYoz0tukh2as3JvkQ2lw+GF8wJbElBvgKut0RWSq
RdTX3fxTKfzL0wGxHhvV/Kc2yFvy+Mr5NzKi/Kgf90w1yztUEKm9FS2MWmALYxSw
5WsalFXxLO7JWEHv3b8Fkotm8MgBp2nKB/6YHaR+lnDBybDO69iZwHIN5cTYPugu
0nP6qwFR23F7cy5fgTojMs1c8uvrt/JABvHAa2hAsMqsRrxkRH7R82HVYwNiHspA
N/vcwNgfohayiwoWfzYtvx2Ep6pdgQTWl1cQ6WHCU5F8VqjzzwjsdpOU2bkJKyhA
lVCKP1LXzXdfgEkY5k5AyH6qchHDYf+PDv8wIIkdBA/aAGE9MtyWEFIk5mSiO5TP
gJCh2UKYW1n2KZDnUzmuTH2/SF7GkZAc0Dl07zyOA9xdyyXEhN+b+g1Y905ipK1K
dEd8AkPMWlD84XFcZw3v/h8k9T33pBeQsp8WQ1W6kPvxwKQI2GKdDtBm232qQ6xx
+f9U6u3/ygdS7W7EmzYcWTWMDbZ1g5SEoSwMQ5t9HwhFteJYAtkH9Wvc5YZpIb8k
NyavdIcvkOM7ILYxDZMxfrrrZFnvFor6fsE7cGNsXHcnu2U1Ll6EZ0e8uy7JN0KJ
UVBj8kvyXHO9R/bmIp4PTXqCtm5QeHbyhul/xFyJa8mMI2rJBiWUd4YMrdfBqKgl
mzWEjcNLg0ZX0lHo7elr1SyxqtAjZ1jxOEa0G2erKIMdy9ccZLDRDW4PoxHmttNM
zWJM7OZOSq0ZquvGV6skdQhC3NblDToe5B7XF7jKl022qwQpawpMBub1aDNUgGec
NFgphX8xT4qKM5yBkURPbOqyDWGPQaFp3FJhWMExZyS9GFsQPtFuFV2b6SucH1kp
RM0U/qfl7g0H3wH2mjQx6tB4Bxh5bnlh40HGfPNVIOYFd5qxcsUNzzv8t+kP5+0L
U6AXKSMM5Q9fTVwjLs4KXYQmi/EQXKIltDEKERH6LYgGDWmZdHqRWWwpfmGcFvf+
EN0iWn7QuW6XOrCB4KMq8pEafTjqwwIFANHwPwUSDFZCBVR36rmLsG0TNUtFN9yb
ZQtcUQPAOSk/pEUBoI1GbkJXRJCdgzWuliZiUD4VvRjyDVBLHpt+Dux0Dn7RQMAB
FCGK9xo7mayX6EkfqIqCVyb3uEAObHwOLgSyGCWPA7eFlZDgppAOpesdubYcdGJH
bN9QRH5UmbRpqW26rJtanDTCD83yuZ+y1HeokFes5RinIORcOsJgq6CV6PwfnaUe
coDtrYECohtz251UDchiNQIMOb7K8kt8N30yFEvQlhtmhfuA5SRPqx8k/WQq8KDe
QtBqQWpEfoeUGQZaKMbau96rJ+ipbCnhv+nherVZ7AoawcR8sxzYSUXsXId5cJSd
B4TBB+zOGSGftQ3DbINcCvpSJECom8WZDdAv2RG7d74dXRmrvgbHleDTBjzXk4gK
C3JQ9CapZz38FMEPlS68ch8zq8qGa3SEnadHaUDwa7DbhK1xpHcEeYnwOSxVOyG4
BrFs9MMUlkNmK1Q6Iy+b/kYGHzarNIzRUkrh+2JIx7b9RXHS2/RuaxH5KlYrfqrI
iy7qIny5Ljmn8jgCgHKVAzlLeokQKM3DjcC0PYPx5nRzMy2k7fhFc+7SfW5ztgpD
fx4gbryoTC4qgxr0P4+AZLI6RKkIJHYZyFWY0qeEwYHa4h9wxfpz89LnvNbnZlXZ
pZQfjUJaQ5eFN4zuyQAyQDvusg/mg4ZG1z/TSarK1oQkPnM7qyTJEQhOslzDEexa
5hS922Ykbrg2ARIP3pWoiqTaJmV6buLVXSJH2BZ7Cf8NIEBw5Sd78mlfkXr6W7Lj
v5DAdq7SQ2tPtyqz/nmNoFjRtTQPthaDhY30fVgK0KqPvoCPRHbCL3vN/TEQzcEO
yai30kEvr1POCfL3myvqUaIHT+qPoiHAxd9b+jPQ7haWpgTX++VEadnMMRJB8ee2
UCirBdoORJRWIU6I3CHriWa2QsXZnTEc5UgaqnbR1UMIxV+FhWXSkCkvk6CkImcs
XghKdoAKIyH/u52+WX0Een3UDirL5myiZcJjbBjz5qZrJHDxwt5onBtWbun65IC2
nbMv+Wvzg4saq7Mb7/o7E7rVd1c1+yZUpQ7/4p+ZyJn2UeF9tK9LXjPQaFzhR9hL
S1xB3LDs0123CC75Tf+2NS4/fqA6/VSEaAaGCMlIaOVRyvGv/gzuP/fVHE7JxxIv
rV6qdTuX07orFHcQbmFBhPkFbxo8R/UY3gX9fBOKnOw/N6EG69DcyqwGzRmCNJsD
n1cHWAbNUDPJdJbGm2rQ1QFnL4VQCNFmyE0EiQDa9UpjnjQvsaZHITvoWq/6IyB8
3dL7Qjk0z3sytw9tKa8po+4w9Q2lFiIcWaqf3WB1QB98Nk5d/rwCxZ3J3mJYmk1B
VR32pePBYWIXnONTIsvPqNnda2OUUfRXEULlIZ2hgFWh9FvGk7efHV41FxoabRav
i3ZpnuUe+l2J5PogH4AnOF6xmTYiYNkdu4WiyvQ6lyPzOjs9wgHZmFtp7Jk2Hc4d
pHJCUjKCDjGD6NkiGhob/RJtcK97mxSBx8XKnAiD2F7jsj8Mj7ZodCBun//ZCA1m
4v0XSWjyRMQTgmZmels8y+aXv7iJ0vVzlBBBo5vQg4Fc1lPkd/KiXXhN5/Iwwt38
PPnGFyZTVap3sAW4htl+gNDOrD6uhaFXIoWQkbFTYJbbuJ75H12b7KAE12Q1DhIT
LaqDH5DKVvYKTh1K7k+DriTeT2e7u4EsOzTbmXyYEzPjMzP36UL9MpOYPqW/qtHv
xVERdxgPEmLafMKAZut5jU6GKPHtLKQYo/WPdq0JcbVsnMPr1D8EMWq8zHQOY8Ue
S6evsenrJzXr2+QPPxohGLU2qSNQZ8nZE9inwE2mAN/xAJ4VsIhdds56UKK/GTWw
AIQeVbUBM8aE2/lSrg2EIUT1qN61QLQIlwljxiL8jVuIwXoo5zvfYadqpeVOb7Kl
/rxU/ciVOG2GJBxDm94bKS1+RQb4zKj56MO+GV4sJ6BC+NLpi9FYlXXx1PYkf4dA
V3ncyUMUofzo2ogLJGArsyKnwv7s5CIJDzYeHwBduum/qCaTE+T7IpA0Z3QSjO2z
zAEVf4bAWiaan8UmbIRbzhRhYDhOFb5qJNoVrMQjLaCWRB7cGigkvwCJVt04k3SI
G6AF+0bDby2F7+Jsp07nkE9VUe8sbZuSa7PzDXROp13pThhEdqnpT+svgekvoj0q
CV0p+53PLRN63Oe7mvLCohLAg/h83QumMSZLnLuATbFPN3am0LnyfzLYSkrkfMFD
d53JKIdtBR9wUulf0ZWiff5HKx4iYmDKBCudtbCdjwjswq/Bt1HWe5HOLvXTz3sH
ss1GmsokujqWF5hHxmL6ZEma3ybwRuwTzT5/vrTViAvf/8HNrxFsSUhDvQHl1w1P
zyKpy4GPAyP1lB+S+FRLv9oxBzzul0c9qKtA3G1j8/pD49Mj41j6y3Ckaxr8uGhN
Sm0ia7/hodriQ/cH8XpoZWK9hGVEULWBYJl/3En9jNRRZCahJJ3Zpunc5x1dNf/0
a/eizPIVvd82Dg6ETBb2goKTqXtfrGKZzCs1UpeCfGoRVA3b8/jHDpxBYMgOB8Pz
gKyKLq5On/sxdlFoNhl+sQWI5xTISsQCixt+M8TruEc67NWyU49j45hjhW+4+xrG
41I/aOk6Xe0B63abhVmpwGz4SsISo59rKZPWIumTryl8fXA3klwYezdJTADnFybG
vrdDp41rD9nkndJ7R5THa0wJfzqg9+X29ggFBAhEej6mpV/luCAJuH+baNxsbfx0
0hL4zXF/n7VdReQgcn4ZyJSyQ6DnAp/yNz53j5ZDGGflvCEWDw1G/kLaD06rWy4Q
lVdV+0xPVY9sL77RjKhVVpHDzEst7VEb/Rz+kkiRHYpBgZGGPutI/n5I4jUDQNkw
uDGajv6NNx90k1UKclIqYChj9pwcETWUmQnilfBeM0GZhYs/2wfVSLU/QzOn+wzx
kYQrEPfEGfbi1nmQgGRTrOlOl2avUoZ88Axbe+60H8zeKMVuo9ePbCoitC+wHX//
yRqYg94hH+YJxG6++cI67HcFu29ZbH2cSAv4f5D7PCQAci3FjdK24AcYQP0TAKUl
y5AUplO0wf999GYZYnz2Cq4joLAKX+VT+WW977PgcpdJJ4KnMbKbHr1LiY1rgGNV
7cRB8zEKUiCgu4FmVMrZ1TKlVX1bOjx2zJLB5FDGM6vucvFrllsAkuS/C5bmRCtE
ZlV2b3B4MrEQBuzEIFcgQGNb364Dn37xIzvR5nWETEnOuoCNPdIypwmPPXWY/8fZ
0rRfpExRwwLWkM7qbmTQBhoLcA/7fLczEJs7Bew8WOk7yyCl7/FwEZU3iWW+CKm+
4TtMOOJRMfeMsuprmpfgEvXW/ZzmyuK0zoq/9eR6Yf/0dCQEm2yHVKNVZkY5UY29
Rp+3fE5tRA1yZ/GyAaCSml0hlWmV6Co+X195LZD7bQ16phC6FnvTxzS8RIUleq8d
2se/puFHnxFJpkjM16HluyNyq0CXop68jEyq02z1I95E3EDFj380HnTONVaHVp0/
ew2+vf0z5E3lysHh4YSDl3UEtd5XSfTrWmIngperDkjlwQ4tjQ9CHRi3bVDAe1XT
yGL0JHiGeZGEOUrGOAR1Z/O3iVsrr3JNEV/wFOIpt/5pglnPVNW60b/BSHTEDFta
Dc7p7NeCSDG1KOCKviwULvg4NWB1BiHWQ4pA3ln6BjRPK8TUW6Pk+AU0NP1v9bak
1DZQERlYgGvkfFu19zg/1qdq4v2VrFVNS3j3OyP0kkVrw0HRiFPmO1Da3X1BdvRQ
PAqGFy1SVx++Ro956kLvWoi/XFJvFfbt8CPIB2SowfXjIH0Cq+Xze9Y+D9eWhbMo
RS3tJTvxdjEghfd64fdgy07x3QmTmNIPWUhI52+UG9MPsidtTPrn7Ty5Jlo+3Wmh
d7SMeDWGnIBfnSI14+AavTEmbvxWFGSqQHMcHC5n77jH6oD8Mnra0xnzNXdVBykU
jsNpqridJOHYWs5gkZqd21Uq0yroklZOXiC5MzC3JH8M+qPIp2EpaNPOFFFD1gYY
JM8saMHPObS7ynNF8YEbMHZPa0UqCaI1JtsGJIkkYMwunDXaCqNhO203uUVSSO3+
zVNr3KTEtDJbcUguZ+uB0ichlipTM1MWvGClrpd4gO6c7PyNcNjOn3ObP2GikOIT
68HHepU45DoRPa0BwNCttzkvd5k8CW8gaunKP4iRde8X6BcqQLrrpsE0C88ESacz
WzU+h/OshDmeElEcXmWOcJ958aEQ5IUY8kDVUCmD4hg3K52h5GiUg29ix7FlcDy+
UH4uxvT79q/GlDEOhdqmE2eYvhaqY7Hvgp+1kfxvvdFC0dzbqDWFWCvSyGhaZec0
vxNUCgnpLSyzEJ56HgxgvhcUBmYHjcTW2Qoz4f22Uht2FbssqBAj0arcgTKYOVf0
wMCw6esTA0h9tna51MlEcPmLjzLcTC2i1DeiRqHOF7ajGom3GcKYgDcyPIKM/ta7
rmT6+Wb7ODhLBpCUuOX0TyKLFfO7NZw/oK1VGMaRkmmhYBG5Y1W3NkD+dN6ojCjJ
6iV/vCke/pHCsEz4Ruuoqz7D4KUzh3EnsOr2GK3pB4vhrRrGjiuHDX4gDSoeY4p4
CwzlzbQk7Lp0HK/TMsipi3MAHCkSaEpS9L1KM0M09esoXQ4mojje5zqHEOTdUId1
7VoDZVEO1DrEwasx7k/XqhXup3zedho//R1oFNzq1J+jkAdV8s2it4FfLShZbk8T
9Ja9YdGn3D2bJRftP2pV/wQzbBZU6upbmxdAISA8QAO6I0AcDVvkLZ5tgiFcm3l+
UI1KCqIb+gEXdIGXcrrwR/E0k4H61eCB2hxB2j6VtXIhjYtBtOhaUuTdw6KfewhQ
GB3ieDBWdR65XDdYMkOfiHyBO/aIwK8nLzkPbfE3wz6y3EaE0/si66INk+ErTuWF
BWdhbO5xbV1kyYnyuX2hhqQA0Sr4fPFH99lJ0ThvSiEzjB+JD0N5WKMPgz9Nsr9p
vfOkhbni9IbO7Y8VJvOTvaJw5REEEVOe9P6pbK/A4+3rx5Csxd1WYkJTZqhIWox1
7TCJji5uzrUONIeZS1MXGRWWkywUvxYFgoNLoVJaHi+7l+IsZXChyoe1LUPH2x2Y
YNEEJgYn2HihFQZVA8nUV/BiMbYx2yGRS3oByc6DgpBauoeVYw3x1/2pQbyZ8kjx
xaE8oOlyDg82VjB0gGvxdCZEVe4JaOvJ9nyFyVjBzHuPCRssAH6OUWECY6x7mkX/
WCvPxYZ28btjW/8i/GUbKxlvmndmJW1ARXIwfduslfq75nZ3k3czVTkcOSObSVMN
AiO11MqbtfBeTCgxppLP+0rwCBd1Bs2zl3ADyWnLl3LWjI7lDYGjELuHqQGb5s3h
BQhkln2iz3I2gqovWprmQJBFJ7o9shQ6XhrrzYJoTt1vON51RAiFGRxYlg/u6Iv6
etCdv01OwAA9eZ4TXngGFDK9atkEJjDHKGV2hwqv+A0/qAIVZaiZy1J0eqkBqLcU
7QhkANuIxrColLYiTwVgsorrrOb3hF/FhcuL7TdVOmeo6O8MxoAWYi1+SiqzzDAz
tYI96OF1dX4l7CaSnp1KIFpVFJfmxx4EtyfnzDlHMhmAe2e/sGPnZ+SBv++HmRXc
tyMcImQ18cZlNtVdUFrraBmZCAm39vG3hMLC7OyJHR6rxfZNmqGK6b5wTHS+0L0M
yt44WVAMocT0qJKlFHpqwKm+j7JZoHiiWjZK7fqzEbaYDeRWp6qQ67zHEA49F0m8
XRXwFEk7/84esbMa7+NGCQSe4o0b7uXQfoD6xOFePLPXJp+bDHeJZHVGApn1Xom5
mVM7dWIETncQsfhRX1QrmIpIf2ld0mLVrwA6WtFWwl+XkzB81eoqc6Vjo6bQ4eAb
lUQLHKtaCoAEDKbSrWTQoPoTff/7iY4sc/jBVJOnDxaVM0MLQ/vldfnM3kduEOV4
h9LC+p2yM5V1TCot614ZbU6vX/fNDaEhCqEMdRG59z2LnL9aW8/3Y7SkZfDn3WPz
+tlcr/1zwsXEgioRVhf2ZaE9dW4cJRcDyaX1jgZfiDG3NqShEJuwtzn1q8yu/O2b
Ua8QFe36WsN5hvrDAojHHgXjXCKWDujOsvvDSj8ntnd838aOz9e/QQsfbRIUvkEy
1sujIr9nE91gklZopcnp02WKp2H8u5KY1cfyh+AHF0997n1gAp92KtZgEM5aknhG
wI5/TQqefpebN1qVhmSGv/zLJqbFtGmvlvJWM+HVAWlsMbPzBYEyXvikuGoYbg+H
cochFIz2MAsoIElS7vlWG8j9lrvwMyi3VuognvZ7OLqZPwgOlUkOkS6XqbFQ7m8a
uk2BDUJzRYFE9C3suDFiE9adqk4VIVnJ55EXhGQiIqzWyMnmP/lcRSkOToKCg+wN
dt2y3XqnFRWgJqd09oe9SfWhmUj/15ejK8RnLKpclYDiPbmp9TpWn2vIGAyAUZWp
9jDZtO33XxbpdH/3tqiXGiTQLm1j2WD86vvh45XSTh8UZ5+8JBst3AZd35z7m47Q
sfapYWbAN4JMHvQPaBW0QexBErRjofdA+meS7/CUDaosevN6SNfxt3UYymvAyJhU
/e4xVvvnwZLlIN24ZZnXfmOz0FmbK06BabJV3kbzud3YSaAsWyEXuBGYn2+Wa4Sl
Yd8SB18PPUWzamlYdODLFQwmXnd2fJxohGg2Ubijgb9MuJ2wJYEef6z1fx338MZb
B6yd4boRlRAAGEwm5rE/UkAkKloOCgdC+abKPwy+cAUgHzDq8M8bVNRSt/Rm4R9l
ItrKMGUuz8T83VEJFCWMTqGSmu+8UdCFBtJ+HlCNM8BA8QMxg4OHGdFfr86XEpSe
VxVbxJ9iuubPnk+y2myW6sh0bB5249Np4wmnz14b0Cuy5YuIlaBqRC5YZblD5GaJ
BhicAOS2x12ahnnrp6lN+xpvINsnBOS1glhlTRX6P0Kmwc+m9j+Vi2+9LTOnG97x
KUsXq/MsPp9JT7P4KVGccq7sCNAKpv93Nb1CCf22U76z9Ypa51aGhsgLMz5HjCOa
lCp1qswsEMCfy3SX4Zaysg6EYwkIp8kx7hoMsgIlg58E8jnkcGnQ55MDBQQSSQ4c
NoRTsFTu0moHBRrOYG87o+7970gZf5SJ7vS3PijUyAWDZl2F7VqkulSnvObFgENK
Cqgbg/d2AdlobIWnGwfrrtzlD3bb+c+FRMSgrK6/ofIf+9NOQul1sjyeCQUCVaYo
g/5zQEgfS5K6Uobmu+Gj06loY41hiT+neRIUnNHCa9mCKWDAex1HNZD7J3aZ1zUQ
Xu4SidASIn1sCxppi1DdwRnKmPxQqomDn4i9W8/0thPyIkMzr/lKx+3q4IGLv0bj
TL6iMRDGyrm1i4q/5RJ+r/ULZ2whA/T5hKpvbQaYpyHabPf6jNRd9XbskS2v0Mrz
whFzr/kgDd8nu4OYr7Mh60v3dxMcTH4DvBW+qMlqgnmHdEtCI45gkG2i1aR8P8Df
Rtigk+uomt6rgYvrAmna3qvJwZ5moJZhfZai0l4UGrCBbAnrP7ABu0bgsvL+8bD/
xCGrO0zS1M3BFqJ0PusiVv8yAH7yIbe2ODtaZB8W69xjieGysECpojxtmz/pRT25
ReLg66EU0CeFHjt+4wQsKhxld2eCt91RHtdpPz0ZGDEMeAO+SOUOn7X0wb0otJoI
T/F5hK6cXVBkdeFezK6RCqzP/y+8m1T2eQ8KkqmfWSbq7lq6IHgeEsTiV63Pb6im
GG+Yfg95KfaOsr5BAB1NTRvJJfXnzn70Noq1FvEq92MouvoqgzptNIMk+A11p2FX
+zCBnZL4ysi1NhPsENVy32DkgiolMy3F9AvbgDeL+KTI0/phEuLQslpncppBYYVN
qz1vmJRGFHFP/r9ZJY9RQrk1fxBQzsak62twht7ToXbyPZNrVCy8joCSUkM8196l
9Ufyz/CpuqZGHOEGy/6dxg2fBda7F8/87dIH2Qj+XB/NIpg8qMLxToJQJ+3cK3W5
pdHbejekkvqE1IvUcSuA6R9m1TzECBG23ZyEOBra0tvxspUYAFThS6n+wj0HLIU5
lnB2mRyz488V+7a72Of0AI9h98fNefpRnWRJVZVSwhD++hmXdocDSUlV6GVDMmvX
+81vdjh05U4pMmcc0elkHIaHUcHFw3s0tobo8kDwWmL4rC64eUMBad7Iegvray5G
XI+0cXR3q2ukba3i/3qz4hpf/pCnYgHw4bjKMwUIc9FKMpazb57jTOLCoiq4Zh9x
i5z9W5Bs+HImvP8o0fIapWd9sI9peVhgC/fYsPx9PZ5H6X8vd/v6Fcq0vUtpqYHz
ey+K3MerLSm8KQh5KAbi8m+4/HMJOtvaSgVs4iSqpkxKtjKWLiW/sdVwKLHuMjT/
+UEsXjbpxMikUY0q9hlRoQg+A2h7BVurReu7cvR51fsGvRLryi5Ro5/gQIAfuzOX
49qQ15esCEf6GlJvTRC5qhwjPtovJuvH0r6t2a/vE9wZIqGSdQiQnC3XULdnH/8n
ihZP8Bmevj6N4sLZZ87XtrG503aA+W1mlSCZVBOXcSavCrpwtGF6JHMxcK161YsJ
0D/SZC5kp3aId9yJ+3nb5NDi49W9Wm1hoYzgHmY/Q2B/+VTiAy8hlOogQB8Fylge
yNiKNqd9QhyIaZ/9ysfLZ1LucUGcmr5CiYJAJsS1bTx7yl3A7AnwkBGS7oJRlsKo
/10mLkYfy8JTSd4I7V4IdlBA9rODUH38qjpfCo5f8wQxnBphm30AJve9hAz2cCKM
yWMB02l3Z05PQ/AsXLfpruuJiMgWSzQNVv83Hl6VwobQ0RPEdr12WF5zqwyrxCwj
9c0nIhncv1K/mBAVr26jGjb9dkNwLlv3fgOLgRM2MiDmEX++ufhIIHeD0KJiWWn0
6SRKrPUjXHTucOreLl7BKzBHqJR7BFjsVmXoxAcbWegTXTofYG4peGZEY6hW1Qz0
8aNR/gpfXzItIkNE1BQibP4Wt0d9r/JzQ1oqr9E5PZu8NCtyx+6nHLznzrb2RUcu
mW6fSqmOstbIgWotUE3DUTJ4NX5OmecK+LMf/GExCFYOUHmGxVNXumCgxMxZTpJS
zYC7YNpNV9n6HIRZUd63iCLXnh8nJug8j0n8UTYX2aISA6X/Z9m5IDs4VK9a5yfX
ZDHzmBlne+AUKIRyWL0Q4Ed7nhRC6SNgnpJZIq2AFeS7mcmu8zSxuXFXqXyBLjew
+pyupl3wlAthDc//QNmZw+y7Kgk4ErfcGEVGU21b/YljnZ7Qig9Ra5jswPkrsOb/
vMiUQILW34VM2w5a+ldA68gZqZYqynS7AORxLxtVlz+OjdB/Q882lJRGv/OJ/DFK
BU3v+vnhg0iE6ar5Aoq/e47ysRx2M6nBllK/cXUG9h+XpWVCoN+j9fPLyawdMUPb
ZvoVS7oJeyTU1S5rxpbOXg6enMiLelbdydFs/o/qIpP9U4wsN1bXeXW3O5qxkBY5
gESRie3drnaOGuZogfdwmzxR9TfZtPDmgRk+tbhsC2JfLMGqi24issCwGPnI+f4T
jXOKczF6pDp8ettCTPz4JDt9z6273FQBElayhH20O2YTpIbv6ZmwmIy9vHChTXk9
0vcJzZJyeg2eqZkhNDSCUAcPYpjh8sCqY3zC4a3Z8sFMCFTfRKcDrKuiByM2D9xf
tvosm3XTktDTLcQ7KLzQ0Z9vdxlY1u8gzdZ2cr50HghSo3INSKJOgVLBpchhdmBy
/h3tmK6jcPA24yGWiYtk1j68Vz4J7hrZZnyUvXYDCNTO8ZtXVWbqHF+0LUwHpAXK
vFAHATz29jRQ0in+Zj8A4sYkECLencSe5YJKWdhL9eILpntTjXe1wj3RHin74u7T
G4f+GPbTReiNaYubVlTidCRtz5RrVz+Mib0NaTxMPUFT7GwqJzUKJoSG0r07dPHO
gmmaKm98W7g1zE24toKD/ZP7fTuDc/zfJgj7USxDVof08cyTG8r5XJP+c+P8Z/0O
uresl0VuBFTfoyb6O5/ZxJ8d0mOPE/Ee4BxcDNOuBMStJRNiEbSA8kRNyVjYqhSK
7vElRECVwxjJBTuDCgkF0e0Z6f5wqePmyt0ulvpPKsDPXaMtYSk28lSs41YRbi3X
v5mkTZJcwLxBT1skW2vaXhsF6EzSg0vhSE5hrSA4FIMckn0TgeGHamiyktUnCsRL
2YQqgN4KxLa9R3CNjs3IYKEK1F6d4FYfh/9v14I1aXeQc/b490Tb67Zt2SZZN6Xt
hswc8mPW1rNyemKeb7hHa1m6e1sxc0Nao+VnfUonvZ7Q96a6A6yfaK4RUMMdvEN1
I1Cn8mIpsy1ldRf629m4/MUMb3WO1OvSzYDch4DL6EE956r4CGZD9ATeWOibc0yv
rGidJKeEzaNpog4hUWy+IE00snQd9LXieVT2wF446uSAvlMjjcCNLd1gg1tRR74r
aK9WaD+zpR6CetEz6W17rB48WNKjoBlEry1DiiKLZBq5j2Y9pJzKgwte7mXJbIie
vNhg7MXldCMJyR38Dfz3sDD+22DFyRmE7WtJ4VIlybZTmX0SHNP/F76T5JuGn4iB
1RI4/iIjMk/o7owu6fkdCFN/4NDeSYvT3cDcHIbLMIRV+fFdf3vvM1f2TJQuHnAf
wmyCqvof96xInxEPswCS7Ld5mD8zw9lWDC3FrnnR47XMV/SRnjc4G8UntUGTj0Pa
An6flA7niCRuQ+U1AlGLSreHK37eB4Vm5qdjJibUCbL8Nhe/Qf/Nxekl31wQCuXL
vtsI/0dZlcGQIRdQlCaNWh93u/sNyge+gn98U1LrQOkaXM6Du08KQoSJ6hNrm5Jw
MDNTYow1YRjGDZBCURG4Dz4pEl/S20ah1xCqF4TMZla18M6GB/OisPfC55IQ52fY
Uz42rN5GZyzXbhqwgCR7KcokKAQk1bAPKLLfp+z5MpRPuQ5D1WvOpFN+ZeKSWDEk
wA+41KiHyPDpu8ugOpQ+IRAuLkuVCy8HUBoAyQWarqV6c+S8/MDGKXlA5DC7Jjml
zEEYqV14MLYGMKTQGzbj5J2DZA1Aj7a3zmLlgqZzKOlanWSXNSwuNL2EKbbofkIi
hW+eEsoSkftEsGbdvCxxUZZMXDGrIBq5ncUB74IhMEGuaftCBCxda3CMkodG6C6a
88omVvZamX0CAVy6rYJAdXKI9V/HJXF6DC98B20cirg4TzywjAZnAGI1O2i6QoQ5
1v8jVb6r27Djf7P5L+p9IviVqvrnDcl6K1inmur9vTafIIBzh7CYSReY1ha1PSPt
hXrcRRak7cLwYDieBvVbI98EL1Whobhe1tOAxlZqEwk31BLznp0JDg7xxh1jdlzP
g4EncCtoAM8byEcnOTQERGxmXyvjBrkw3Gd1HdHQQ7FYECN21rV7bnBwbumIDCdq
/wTei2gS+LKNZ3hL3bKUDnzW4pqtLxPYOI3iuCuAonZmn574cY94UFaep4eVVmtM
xHwO74IyHjBMss/1KI9apMGm6AnOBScE1IA8rAfCmHgg31pLZ34Ma2gAS5pPSxnD
QH/jycfS/EvX9btzN4nPt9H+rCtw7ap/yX/yrjmzErfwgDXPVaqoiD5Ek2e3bcEf
QtNdxGjeA4rWZfOicvFhnvfgl0Dbs1ikwQ+iCun4eQoYVHCdhkCOwDyT3ahQhMDl
nYoZiJEjeymbUD6cWgqIJ9IeST1KLLAImtiua6UkfOAsXq0KII4qAwytxfJUApZ0
u1HGBZjcAxUAU7eYKXn998/LJYp3iws38mKxlq48uQgFhkYLXSKM8Y/ggBzOXUaw
bA6r5QdHO2C5NSVY2lxetr8fvugk2ldXjJmDxPjJE1xbq2BWNAKXI766KuGfsZAk
Yv2cFze/hUMRcNZUbGduG6UTRcGkrUcphQfJKG13A0RSvNYhRAwK3PleRj0jP7Yy
4CslDJNz9QQQvY8zeb5uoUOKAzT1Jg9TxVuVK3xYdRI/ni8UTM2YqqL+4d9foJxx
n/FMU2L9KH3DivUnq1eKWMkMO+vhXxzFAxPVGoUnK4q5WFSwDEF6yGun/Qk2W7WK
Efa8qPD7FMM9soQRwIIJhIZ1Nt3nSKY+M3HPqz7ra8mhVB3uFnvXh0MBwBkBM/S8
S6GewIMvROA1SvJy9k8zGo23d8Zjmj97eAXt7vBnl7+iEgMZGaWiXuUYOk+9ieDB
9oDyoGrUmfnshFifpQSkbFvZrxgahlcn6yh3n5XMfBTMs4BaDaeA8VwdAvITx1Da
WJYXuz208QYDMkVmJntjwtKXqwEch2ZwZtLV+qGI6kGIBAU3lhwqKkFd2l2S//z/
pjECh7ZuWkZLyj80+pRVJrkY6k12QoxtMAycTCW0rA0wGsJWKsXE9NH+BGD1PZoY
/my51qxDfrbonB/JrU77NhzI9CrSUthhuhlvRKmgexXuWfmQ7onXGp0uxgFZXlpI
eNgJpmC3PAa/sTh/78ipKEegSwa1zyVQRkArKuI4OM5cBcHLy9OeT5KYJIuOa7Zv
wfZaABzNozLmBf0jbzRwJo+TUnxQ0RZMQdQd7tSVlGCgdKxJp/EOsv5mdiPd2xv5
GY6tZT0ts1jLE7kqBqDzLv+obY7gv+50bUMuxKFvVYt5rL9PlsExSGwleGiWmcpJ
P72M1CeU6GHq6yMxWdmcH6nqV1UZ23wNcXhZSEXWk+/LxaWHdqG3AdMdk2CyVDfh
e/cNE9CV5KoIR4XxhzCEy6EFOL9Stj417w4dVYBAwVXo2DXog/rNbv5CKddyWyJE
eQecs8kYRnAf5HrceoKu3WFxqCPUtVZAprBENL4rfUtdeG1kRhoQz6Dfymk73rms
8TiM4oQ2hL/ljlW2WTDVRE+uZvdA+rz7yM4h+hGIodFA1iZcMbTgOCf8IDi/DF8F
Vld9oxtJl0uuEb6EZcJinWTJfsxEaQcmaKEHl/+cN//do5TJk09jcilrDNvp8qRU
h7l7w4UzexEXG9bzxTN14aRYHpEg7dTj7UJaI4iciUdcD7Hh1+Ip9ohqQ/ms1McO
K5TLDBIlWLJ93pR4gKUKogwSCx+S+gAW63LSJFqmZFHGoZdE1NsMMUqSrnqptGFz
iKbvMtK6fcBUhUEHGqRqYew3id4FFgc+J0PWHXjhH6ZWD4ecSh/FUUT3d/9sLBvB
ZgQrKDe9Lfl2+zcn758zmfgPm4KwvcpMUp9mV8Dqle4gw+Ji2HfGqkhG1Z7DI8rM
SxJ8ZLouTBdtTdlV7vnJ2QDPm8Iwynuuzvx0Li0HQvB+hn7obpboE7B7FwPamHG6
MAbqBK6x2JiUCHAcksKctIWgvhs8Z3l7uRcaklsxk0Vl+JmIk9ema8WHa6kn6uL3
c3wDZ5/bUGqw5JFgM8dwcDkHyfmaH6ji3L5QCLsoOQFEEpIf+ypKnTtOFtn+DmlQ
o3LKbkAUEvZlq9yrlgU8+Uo4VxOnZwO+TgL9TxhvaNkzgJpWJR4/i++8k4Y0TeaE
PAXKVZQXMRjOYxtj93AjworKjDtnfzKPbK7UxosKKmCluxeARjZTHbZDOmBdiQSR
004071Y5ilYXFS17exv8VywWP3mTUvHxnhc0DPjFPNHhrYVu2bybJiVFvKqyg1d9
WZhRIx3dXEqnSzt1B/2uh2LNGUa8Qo0T4ijRTEralNFdpi+YABMBz+2RSCJiK4lj
7tpLu7l5u6XYP0oi+/x0HORGBio5GEOsBzgaIO/HCWB9I5PoBgUrudUkLBAWEExp
gjMNPpVmqeXjtt/9exFNGIZQADSCbdsI5R84Y+MkYY06QGvqboCNCz6CkPLxm1BA
ESs6r/e1isDpU6Ys/reM/txwSn4DUnpuYCNSwqlN9/RZm0hZCDaXoxrjAgRSWkyc
ds0b9ClkKSil4FksMbW/sUqj/JhRlnSZYD8pC4JbPbrvv5mixYBe06EVcJsCKPc4
lvb8K2MICnh8miAv61cjI7egKcAZMO/bfk9XYbvrmueRWsN3rfhbx/VRDD7m0eff
iv9K3mkG1y7RqZd+am9EQbSiKYXrYf959xsdLiNPHoZ9kHFS7NZh5ifjWtvc17j7
0ukfiIdlOC4gdDM3/+ylOtSG2YqZYW+nvrj+YyHsVrmpPYUPZk1sLc6W2zJD5QC0
qhpgpIV/9o+qNjWJ3+KyxDdKmAVQAvBDrNL+lNJmSrCqouCPK7tI/gHErNG9NIL4
ANAiZ9Q7UhnevhEMgApSdANiMAmRAa6ge/Nf0yB/KugJUKX3NHNp6qwzG7Go5Uv7
aUmMpzxAem+peKtJqROz7iOHUdS/KkDZ6z9W9HGcuPlhZo1eexH4v36gUz/TlBad
8mjkxl/I0U771Km6m9JbGupJcurPEDDXaM4pEUASjEY4DLKlztMbdAUUvHuqV/48
A06CXKxrPq223OoOLrC1Pr1jx4/UIW/sLAw1XyjKJ6f2yinWXdzE7nJkt5BC6Zsi
Oon5J4IWG+S0DUdxUj//SNiDuvoHp+pVOhxZsCqIoPUb1EqzG5He8lPxxLGj5/z7
5gvbqvuGwOTcxDRMvBvvqAIGfVLUHw++z1gg4RJe6ie+R871/bvF9KeDa8aDv11r
ikEk2Fk300lV1Xf3OyB5TQ2eoBEGUHBU6p8h9NIV7I8gB96zfWOQm5KOMpRoRJiU
u6sVGc/RYwR+bWLIUL5z7QSHzdP/aNeAoQGVvNtgc1UXHJt9JskxWh31PcDFmkP0
Nr5RUjsEBIkk6TcDbVVvTfKrmEmJXXDDP7Rzu0iKmKKZsU3LqVG4KIE/Ju6jV4Ts
EAcdCi7fleEKQSuKpBP6J18lANQKdRhoJ7xCyiuSSfuFUDjVc4VfFPpoG9FqMXtd
ePs8b9cYO1ItOCpPJifwqszOcs/xW31o6gYJQRelJbruhhV4dGDnlh1feN3QqUjE
V3Ymd7a892hl6LjL2RvZEohL99Nnb7axVCAShAXmeSnj84ZU+OdI4H6SYh6WFgJO
rbCjMX7eImhERCYMA92pXX+PrZF9eNfYOMlpLxk/+goBQTQV6/g/eRJ3N4MFQivA
jZ7evRsKNRjwWnZQtwIxcQXeDHRCRO9MqPh7PuCIJr5RHObaD38DYguyt8f68ymX
fNeAWx1Odj0hVA/VAftyXCr/bwec+rOySwgzGcYlBO1vIJe08TYZfK1pudeaVOq6
4R6z5FMsiTUHAR7Gj/FfAb7Tpjjxje5rSgyA/UfPRnhfZ0Wq77DPI8jWgINTZaBq
U2CBCOIgWV7gpaHiSjZptlx18YzY0k5InCCeSxOyXBNnLoren6F6gQGvMhNv5IxU
NYRkGJYLyBbre3TU4QTsZnUVCPXYDzMnlAIYCrdf1iaJQqqDVVIBhxX9bM5tvqT/
aAqzj6nYJ/0x11crYtLqjzbajouYPOF/LWvYb1s1nB9/9K9JtYMkHGswDoHLmWmj
lq7y0yp/h9Yyn5XaIKwmoepoArXdhs6RWixQ+5I2UzoANh+kZWUAkQa3AHCorkcv
a1GTEmnRjWZLSsHMbl8L/3ah6ZweCUudsP+c2I8MNNJlb8Gv1YgKMAeyXMkJbGOD
0wzKAmAb4GdI3oary2V0rXxvElWmUnC2F1lB8AJFRAT7hwb1YA0nMm0kpRY0QY7u
ROgzuxDVxwQ55UOb1kX5WfKD1qevevym+jhPrp5b6I8rtGCQetCgeZWCFSR3LlWK
sQLhToGIln1xcu6R1IYQ+D7LtlACJjeaERRjHA/2G42+14WcVTOqZQ39ie6bvEao
a458A6onJw59tsxloGf0VzAhQI0T27g0iGBDfs2fP8pvi/Pd9grXqLuE2EaTXrbZ
/zsOxJbxc3t97bj1m5nwDME/pl3AvRn37YwtuogvKyZ6uBDBC/hsoSXllGoQ3L/9
zK28ik22UriOR5y/dyfMOivgnR5QzTfGah2gu/rebzNWFe0eCylFdD74E161y2t2
kukNJQFK5a/D5BgqEqW4dc13RVSooC8lKr70Gkc8VM/zJ16q0Qj3LP8dXoyKawKu
EUskgxS0DjgBriTxNlSOT1PdB8+0d1ygQInB1mOq/B4Tm8/J6/Ff+iz72huJxVU/
93hQcj1Ksk9yIysbgENiOzeUAVhDt93M6exrRtmDZFizeUi5LpFXvsJGrRQbkVxG
iA/fpp/1oE/AlqUyKBPFhCSp05jE5beG7JUQ5myXhrqiehD+9OxRV8FsiBdaUf9u
LA+2YOLq1D27J+eUTNmHuK3aeOfM4FMVl5/GwbIziZbNJzRPrNrNYdqm+Aa8iMtq
zFhsFEv/n5OyA0xlc3Je6tlFqFfjwQs7nM7//2w2ynOL5+avcFoElhbVNKEfEBJM
BYW/uJwWNLVAaLuT6fuN7DV8+uozKG1VQa6mjN/yF3MrISooDJMGES/I1d4ICP3u
/Bcsr6elF81E4lL94t8YISSiJJl9TDeeBOILfUIPCs2hd6lsYO1IUZbQRe3LMutr
1EQ8ZtZ9EwpVSldNdYb0ka2ICgOU49kQlS/DdKYcggiaOo6c7Ty7+PuxkQ8gbf8a
8mLz59X02WH//0uj5/18CdFLrd6oiMYCkZCAs7jalQbhje44qJPMYcArsZAa93tM
fhfovZcjCM/6Ij8udymi0sRPjlf9Wv17bvaScQ6neitCGCCoAhqvnLYFBjgxLplZ
kr+mijRVNptBhA9lT5L9TRHgTkWEPnSYYCI5ElVGyicI2/0Kryuw9O6MVeezL/r5
pt8tYDrbh0DhOkFKitMG7lPR0vRjg+hYFQQs47BYob7Csat41vDFkHj7Kyu0ypc0
7nY7aagimJLNGssHf/e1UIWDXd3vjvvg1x6GaSjio+wothHHKkBmmnEi7r0VmQI+
nksQlrNXmaRs6DflMpjUWXK19kwBO5UCY5J7CzY2Enh3+EaX9gK9X2S1umS7FoVp
jbSA5p6MWqA6lOuopIZdGDjMtNK2yoVZfqovs6pnVc0zsdz/L7/z58AHtka/kyna
2ea0s1JfFhAbCpmgYH4uiiDA+aUNdC5vwqBhRAGsBmIlarIlCtunaXW/Nl6w5lCl
txvLiDyw8Qlqnil/w6U97SJoGNa4swt3/nf3zKgk2qbTGfgA5a2XvNLihEwnBgpo
uDjLWv11LFxA/TgCNsb2nxy4WBkqUwR4fGKHnMk1vC3gg+ASvrxbunml2ohQmrzR
OuBDX5DYCFanqxh9DN+5Mn+1aTvhBsaq6hpZrUAGvDcbNrM6uefA10IpIXe3kc27
iJ6f+NvUo7V5/Hzl5bZTCLRK/mw13V2+bcsgl4Zt7sK8fhBK7MQ7AbRgwog8PykO
sFqCRgPR/x+nS6MnAFVmhAX7tUk4M8YRWRL9K2ab+W31gQVblYQkQaNcQfmmEPMu
rG4KuGVi4/8qsM58UO2y9hJBoCDlZrB1mxd598q8FX+IYhbXTJWN3rKUCF6BmNxN
wkDlHmhx2WMuU/yQJ6jh468arjuwqRdkoL3edVak6bDmqoj+13o+m7pjEbQL/LzW
RXQu79lJTiHloA3vTLIr5oUJf5kihoYmk439fUMGVQJ6iQBra0mrgR7PmoI0F/B0
OhhUO0KRiUi2zaPu8d+SCQhAHmdfiMMOoT2h/zLQc6mMZxLFybzxFnDhv28XqBJO
6RGEUDVYnVzpohhNHZPbThRPeebfBtKAjXxmkOt2OG7O0draUngDND+UCOt3crzS
S/bjFy5E6zC1TZLvv4oEu1Y/RQFSwC8zjrwUDrImvDvEMRzIL6O7+ftE8kDz7e0R
KjlpHbXk68SWsgB1xEG9djWS07hW7EFYBuhMGnegb99WbU+b6/AfaaDB6zKFUlZu
uTuHhETf6kfbF/LYRUjLrkxPS++vj/v1imaXk2z4E3KQ+FvqyvgajTqBDegZ1vcn
4Y4P3j48VrmqTVbCgbo15+hyPt1I5oox/5ysMEQ2qnCBVrmLeJGbSHuafGnMl3R9
zaRiLJgfbhVPD5GsUATfd/3WGYl4h154JNoFtvIAXnxtNSxEB82X5QhEW0k+wgOd
tg6ZikUW1CUD8JlFnF8V9UVi6PGtuOS31c3qhN/Vn3xXBn+41H1sUsGp81pU+Tku
lWryFx1h4JEoRnuyuGa78Gt43wnFjoWHjAbJl3pZlp2zUYClsoU/Ma62HHlkxSZe
j05GGb5DcI2+FvRs+StpOHM1dKQW3lCd6b3IwPfuXQeZ7vozY1e2rrsklYvYLGJ3
434ZjqcuUTl3y63cMxI+F2P8PR77gXUy6B6E1AwPhd6pzSV3ACwtQyhYk+jFoX5i
wX5Dk35U+lJMoFNwcoGV+B+WVHjHpc3wQ6/19utcH1K2p4zmjGhvWfwyQVChONkw
LeKFzLcNH0hu06DumWTTYt8wewLwvquciQE/aMIo3V1QXmgqkLpq6f25FHwJJA9R
Bg5dgivzlaOMvu0mfs+kiBSdBCZz1tApYWoUviJpo+lNoipqq77ZUx/WkKIwSf31
zRynvMsma58J+ifURnnHMxaUR//4d2/96GA0IYcUTa0KIItSjCUvFCXM5G8XpMCj
FrCVdbuCeEgV4NMMpu8Q2NWGxVOgx5B3URv2uHK8z07G7+F2wv0vZFmF64fM8l75
+tY8uFRDrREogzDk4tQSFuwBOq1MN/C6lLjIeUwEPbOEeR++Iwshl/JZ5MLLjpGG
TpIaFiOmsKFPmXPFgeNJ/G/HT/kxzcLU+a7hOxA9IPIgkSIJWdreDXkUspqIQb4L
G1nTD6SWzcElhSsS3ORyZWhYy9B/CGCGafLFymyibs9k9drGQuLFCPzjSOUFvg9B
2Rv5uHVr9kYr3mTwBZ9PnhRoHjR2oUUBUHEP4Rgi29ppXdXr4C0RYbETofUGy6qs
daEgn1Pxl5VgevdFGutkhf+/7NQzIzU2kC0g3ln5WBSwKoVs4GsSEzc/bHZ7NS9r
LvCZhNccGxJ0hP5z2WhxFtxIpk/ulgto7N4rRpugntTBW5GTf0x1ie99CsdwlMaX
P7iQte9DjHyV4DB6axXREbo273WZBtokg6iYMU8fXflIKLqZPYgXlvlekfMroS1t
+UOURjafToQdqQ9dWhRYUhVfXunjaMEJZArNTmJAyJea5p4QXQgJDf7qP6sZGblK
Ue7WegfRNYwUaPcuwPFzV/KiSqdGWjjH/1VRF9VHk1x91FA8ST0T5XPhDw2ArC56
NGQ6NHaMhmYUdhTBuvBufI7llard14P0gDXQziw3zjx5fOIFpxEe06o5K8VI438B
5EsneCScdmeLbh5ryD6PSszT8jMOKcAfhuzCtX1BoVtRaCuODh91S7hATf84xOW7
g/l620huFTCX+4l7JLMz+iFdJxzFiJ3ZA9YKKCwJ6OCAa7HcLxl000zt8JgludiZ
Wll7lFA8DpDE3u6i+ooNI8L5K1D53wWN1dbNjC1uW0NN4QUtVxTD3h2NcbyGdvS5
MxTGJyStk92jnNpNCJGjAkUQgxS04vs9LLjGEwRX5U+6mSWvY9tP3YDV3gbxEGJd
Tye8YeAqNXI3GjxzGBJQ1gbiX+BeOGt8wSxUYw7MOFdAnFkdhzDTmCw+xxxWfjTf
EQkXpUd1UI41voIYdZ6Np0sViIJO85e9jqMHC1QsRzse+WWpwIz6s7lDp70iGGvk
5QKxu/U61UEvbEFC8GGAcOqcCSHYaw10SwwDOkifsaDOO1RwmWqDAOlmvLcQ+y32
kizsVA+2Mj5kXZRdcgaQ35r7j/GaGjLOgaBWrG4b8qwfOguUdbsmmt7GuTwDqB74
J6x8DASbtv9MxjccF9CgZ7ti1aGpm6yeyiyvq7R3yr6iJEkexcqaQcKRmcun/8oc
SpaNyb5qJRmegUFvGg6zQBIVkAS9HAI1Xeul48k2K1lj6VXrDtvoSlAYJ3oO+w8h
Iu6ghWc+nPjgQW4pAHjSOc4WWsqTAscMrwMeCdFbf30DEw48+S9VWr3cuUfsKCaL
1EGJsjcrYdNjK5atAE5gbnbqkRG4Ih9cZui6lSFN3BE5TsFEfMaRj/sjM+fBs6Te
3/jh67u7FfL7JxUWuiT57SfO9yvpnBClGUG7R0b1hPA56pF13W3RY4+c95oCx7DN
eU/14Xfm7oBDcgX+wl+q58g9602BMrWmDvsWgbI4/r6sXjo+gpJCoq5bZBzSr2+B
HuKZo+w0Q21VRyGshM0VQRHX8X3cvlcKIJxJJZxQd/Pge5GXTB5ZYUDFGAi2D/Ek
2J0qeEYH6PF63gQ686pIgzwfG2fx3bJ0RExN5g+iJD/1HGuRWQICsSQl/SNhJ6Mc
yKTIahIhVMK4/Iyk3nHz7+xxrlhR7UViMzuCa2qUQII86EtyTRQ38f/s5r4X1p3v
nCply09izto0Zd+k5lv3EuIa9x70Xd0J7sl9AXBI7NhTD+i8Rd5ZMUJNDNLjV6o0
2KyC9m6pT3gDhDqWt3f+7GfZ7Ko28xBLLFzXCGEOlq0ahsxCdOFVThEp+SHs/cot
Lnxi5upDnAy9oyX8OtLzycZ+mZ1/yvmkdW9zF83wbeP1BmNehqq1B94s4fFoZkXc
0Pyp/FmXg7PsMsYG4VbFjWbBNqCv2ZlqvkVyxlP9qpvw2PCTqjFTZ8RU35K3glma
s95hMaD5rHllon6Rq/JoMrowUBjUeUzFEeiJoxxyhops1qxx3vNiIJwQUC8fcgFd
9skmwU8RHDiWiy/3UROfKiN5x3tkS0nfZv2jC0uEdlLZ4oJyQcmnnMHrbYT9t1PM
QdId/FCIzz/FBNqNDubgaKnLlNxszM130zCNPMYnYIZp4PIBMNoBUwBWEuCUXhW9
SFPpMKkZgIzJTqW+lCaI9kOSsDzblJLrbDkuS2ySB3OM+syyq13JmhSP5ux8hpi1
FG3NSqbrPcNfMSPXQBkj/wzWHQBzz4OO2HhoHs8JUlWBclx3kiorqgYaGzh4bRYA
EiReBwOJ2VOImaVZcj/tlR+xPxUw0qY+uyeDOkaFCk9ZVwYYfHqyZp+hlnTXpxkk
q1trX88NxL68oWxvHkdkRMfbTtmiqVy1KRIMbwzVO6oBe2K26dmONJvc4NEuhS+h
m2rq77r7A/3YZCbj2P1PJVkUVREnpcRzK8sfRkkYVwO4uy48X90OchCeoMZbizTq
QffL/CbPBQN6QU53jOnNnTWLyLVSlUOHV5qSqBpNToM3RfK1ytg2WBRRE6htnQc4
ZpRW5YiD+tuNCiW3mpbtjBZWri/UJ2uVWrTXzwE2lpEmdfxElNYa2e8ulctpmo0G
Bn3dvv4uvh3GHZi55gpKUvs72cTThZXNn0zLrlOLjy5zy2BLZQKZDTky4DP0PFau
SbD5iddYAeHFsyp9zMPOGhKMcF4KzEWlXmubITy5xF0AISB3RieJ3XKrG0KS9ncl
B/UdUHIgj1xe/chkkhlh3544804zR8UqmfEDtfI33BrE+OncuutxS09UjlNmeuS8
yJTuRBmW8o0sjwOW9Gf2Osyj59EsbDNNz+Rg38YG2Mw9bkHwPVNlSlzpU4Djupcb
zm2/cQiMqORkT8+TjLGLIfG/BAfRy8USRa1HnKyGl+aeOz8rl0LwLB/OJ62nV8Cp
r4t0Oy/buue0BxIBJG4VupN37PFZxVZOwKLxo3U/B6/ymc6vkxIW4aBwhb3RUXLx
Zhnj9XCvbHfh176PxiJNCeao+LYzseicnlCMtj1CafOimnVWVPmFfIipJRBAAR7h
EJa+AFgi6mYjqfn368YzOPgVvfkC7rcCPlcODcq53MnXep5y5ZGDYndnLOvJyyNi
OG9U5oh4F8VgPeLqP92aYFpi77noR0yrCKev/AVwYdWydCZ9n8W9hJf4LeBu8WAi
EM6tQxFFcmK4sAXVs2hY6RYQrZNYO1RSs+MtufHV7bK48YMJUoMnWCOj2+K1Oahf
oUIAwuV0y9gGg2QsyfYQcB2HqdN5rkfX751NgUXCVA7Rutuu188ZsOB9BY9HBVps
TqZmnzX2792i7DvTti3K+ht5CQsxZbPBqR3FmoS+AeFqJsovCvTJhGCRauMPJZ2D
SdpLwtBo6N+m7AsHmBLmlhT17VLxub5HZ8vULfbOR7+iTqixB3usgcgfSe2prSr1
Q3YQI4kZIdkSqh39sbLZtr2I6Wvzn4DMx7X40v82hqP43x3VBdjjnlkQ1zqbbGfn
RXaPJPfvMrN8cs5bmcf8m1MONl2HpOQ4whinSNNo/fcnBHTShVnGLU3lhcHwiBTu
wIvWTnCKzOrO+jbYmh4FhiXtr+4SqkLmrOdJZCvdrm6DwwKwzTuSXW7WZ1Q7Bq6C
52YM+YHcJkQus5wGfWseZGt5VxEAhidsooIXxnZ/J6UXH/B/DOLOuNtCBXg7O9Ha
T2fnKHqxaUMx3TLxVnLd6Qrw4teo8kO3bBsaK7LUgXQG06j5jFbRGa4xwVlCKAEM
7na5tm68FaIvb7EsIETnn3yeyXr7VuylhD2JhgED/Tj9qJlnpTQyNjISGcH5h/C8
y06u0ddg9hWZlR+4/STv4wEKcMyz/N8+6Cc8amK/CeLuGZl2YA32DkCLmy+59vHh
9i+QoCWBATc5DJpDVYCi9+uKTj8Ih72k5a6yX/RVEcK+Dz5eJtJjlk7vJNk7mJUl
z8guozvAnU4ZQMjDPHVD13fjzEg4S6VA0TrBozFfHuWno/ZtKk+Cnm55AHXtpX8a
U86IBE10HHAIuf3up0QgrzXi8AbKKjUuGz7lwWAxnEMb67E27ubHx4yVXQwS9mbU
ECdQQeQ18PAMyE+MQEI2H5DtqhUvnfE2y7au8JfL9AF3kjcOw1kZwj88pJg7Qt0J
6I9/Hhe/pe2C5+shBELJ/VhYBqp2hWiz6L15ofnKo+pH2xUT1CE6/5vNipCBqo/F
GuDKzwqN88zGc9hBZk3mE+1lpEubmLbsADs3lFc+y+TKb9XJ6PGgAH5vHbik5owG
G54oqsGWXfQhIXBgwUl8ZPcpA7K/AOadrSlCuRnwyFePQTcdr/kHvkebAOIw2KbL
JEwWzfTGN2Qo888p4RNmwWfp905vSIAU/2Qtp5Vud5V6iobFfZj9DC0R3Mqf4yFf
O+GbFESxGDEA8C6s1aShyXbSnaJ4cbEYV1I4nIPHeKuLUVyKmNqRvELTU4DPeCAU
c0k+5uJK1h1+z2qGULjiY73FzPt19vd4jNmGayj45Tz3GJXDpmAcfnfYtQ/vbwD/
ROCrZurAArTo/gCHDDY/pp1B2ScaQb07QOzaPFYPB+sybXLnbuj87V7yG5cBSTM3
b6fmbUEQlDgyYY3vpUAHwSF+YJk15ohcZ3fvYXbHuAZNijhkuVOG7PaBD2pwERu0
EnRrVPeEsjAh93wqhG/mC1pSWWPzItxHqrlPBn9yBu1SgRAoJjNoAX5c+vhSwre7
QuBxQdN82e5Nohi65VykZjfEBIsxMoDs+OOAsWZE6X2xJII1sa5kd+US6UDcyhXt
ZvO0VLPRTgxygEe5yrn1HfvhUi7r3+nfSD34Wt8uGUrw6gew+eytidM63a20Tmcf
7Kph2VfunBRk+akPDcpu4GG+aYaB0SX/QgVTJWiJEAZ+C+rDqP7yWQja/uQYEQom
EzS+yR9V3dZyEIpoaBRIxfTauyjmBLFdgc/ocpKArj6BaMXOA3EvwzFEWmk/xIOK
J2USo98DLSbTe178xOXHL19cB0gCoy5KhC9aD+DWQ0VbK+oBkZBN4Z4eRJASmXro
H6qM04yeokJuVQAN5SdUhnLpNSjGhBkW8dP1H8LpRVGoKgo1O5RJ6UsYGMhNxlDM
rj1e5dha9L6wUqEDiOCKlCvzJoAM3WUNcjW3Kwi3l5RO61aU8pM7m/jNDYsX8sDc
02CUN63tjr4kqA21FuuAdDVsw4tbBtyhJLwdE1CKRAjCJFy6GFYGi8Ze2xYqu2g9
80q0pXh1kPidl5CYJdk8Wpfqc9c3SywRpH2S++xSpPujPZDop9J4MXynCj1DH68c
TvvtgCWRnKMCPvRomIssH/k89/qvw31oY8oGOIG+GWEeQxFVU2He7vrWYjlIuME1
jjutu4rs1B52bPMJNWJIFM819GmCBRiv2koMX5ba5TBxImLJkKgmcYO7IELFyj+U
60LrhnpPJQh7Humh+iIHSMWAp5h0XkQnKpyw/D5VHXN+HvBHsh0P3ITPbqNdeNkK
JnZfp5E7OlVrlAPbPzTlnnc4jc52+FBNE5JdzxQSCF01xODl8yQhadOBt3Xt14KL
sAHFxKRok3pBxTbhlVd7HS0t7Z9TY98RIXZjCpWpOvwP+xT5JmmpgYzqXN2Cpqmg
2oK3ttI5EdDN4qajiUaxiz/YhW9CKNYOO8xwK1xTcjnML/gieRm9gkI6rRRnsSeG
AVeS8n5DXQopYu7/AEaXs+4+vmI8MDMoLc/8x+ni8pX0BCigOELP/bpO6UEKDMPt
wRUPoVklKmtmFobBlXFu/p7Z1eyDGftsT4lGgnpngzj1gVCWqgqFXRYUVuyhz0/i
0WvtUz4J2P1p+45Lc1MJ5qt9aVD0JMoW74nz3AyPdXLu7ei70vzyNt8fXn5rY2vV
Jl8Qpt5t5LiYgvJOW8jgpyhf34sB2wZ0isTNFXlA/PQBwbPmlD/ctQXdnTtxJMt5
fjJGM7pWwbk0tts5DpY2b0Vmwxt3JQkzX2D2wmvtx16fHpBY44Awvp/XZ5nhLDiX
qzHjAU5QOyQHkhZ8AoTWR+Gg52fVtBByqJVOmmns+k0HB++9ya07/AKRhOeCk/Ez
nr7sAhv+tSnoA2AD1M+6cy+D1UXBHUzKhEAHo0DijNRQMgmiRFMJrYJMazuqDPak
e7BUwa8uIklg0hrWJhYcZ+mUUOh58mnBw1Joa6IyqAmLiCgy3EUjyi0riFgDsNh4
sDAnIuGoClNUDaTPgjyBjdv3qZJ4Fggj0P3Uzoc7wDWBqY2yDjgtcw4r3MSwxL5X
Zlb+4078nY7ChSuR/ZvYvA8cmdqiqAviJsxOk3Zqz1rqs3wCvs5JTBY/V4+2qtkw
Y6ORU9JP2MzYFbQ5rfsNcqwgR1jfSLSV1seKus4i6xvP3Y+JfrsCoBQlTgn7Rf5F
o78yRAmaRJgmnZ49X5Q7zdDpK461U3kgyGk8F1RD3wHatXjta90QwX5sSC8VCCB2
qK68xmH7zGPMdSp18GemD1O1f7WyLqw2RR9Mi/wL6mBw1yqdjV+SWPBbB3mr4SxS
XFjtchxss8oQ/BnybXCWrcuwS4IH2D/F6DbJrwBO3NvtltdZkiYG5zIc1XaETVtu
9OK3AkMSTVD18Gr09BGyCL3VOFdN3U5u3KwaWTO82k2QcHqHIG6KA/ld9cbxL07G
k5Ta6cqPYG7hsT+t+7dykBjwlb5WyD5GrtJnpfyFcUjQsXnHWgv/ggiUb+RFHOeq
0YsCADhVHIAEoNxjhwEbWJI4mOfF1GEZ+BOND3FtDUBfwyaYt7iH/Ju40Hxe+1Ab
99JzjAwjGPpdQkEYS4Fo6CEjHCVgGLeV/ZP0iDRAx2Xh6MC0vwTLqDEx5XW4ZZ6R
7TbQJ3rnEBcWPW3/ncAZWcHn2quuFYrwHQ1wFAd7eRPqAQvCJjayqbAAlfCMXIBc
4ldHiQtZqjGzE9nK7EfP/bPMNmthpBzet86ZudTM+gZajDHj35CpGktdHJzyYEWR
weCwDEuM6flcYfnesJgs1xfaYFFEXl7n8HbQJ9mBPSB4rNfU96N+W42vmYfLQqU5
vWFtQL9Tfv59BSqxi6BaZcdWaFBmvNi+Z4XPDECDpBaxTpxzZcRYPCC/3J4z3XTT
mOaI7tvlJeEUMa+zTDDf7QmDCSPimhbVEAvM6FuDPNG+PajgbOeC4ieIm20rWX78
YpWsO9kuQq4pxV1u3PprnE7UqSn4syGBF/Epz94D9Qdpqv8KO2gdYHagB7C8eu0u
jtMOXGHX7MmMzZ6H7tSQcpgNvWyc3oDv3gWTb7PvnjYO1Mkyvg0a3Gpnw3qJvwmz
32NcY+so0w6acQC6IGt+ewyzzWmfcjOnvapyVX9IQ60cATNThJ734mPZ+d7+PKri
6trFfw8SfuCbQW146y7iXGoJr6lTVhdI9pnMxMj6FRLiMQbekkdfBIvt745/+f6R
CdKVQbU/81nXhLydx+8JZfRz298Q7BWJ1xIJcgxua8JLVCoZK1ofEaHU3w0Th+Wd
mUE8VcqpH3SHzG8oqVtZ4/Mc7cCbs52+Iv6oRXQWw/ckvPsi6mmACD0o2rdVX7rz
BQNXWAoE6/kD/53w6H+DHBpqNfQH110MfDnXaRk9RFB25jQWpGPW8x2rNqZSMTTP
tbtLJf3sS8MQrFBsQ92iYHM+P0xO1U0te5C5MzYGmZZH7a2KgzDrKtzoVggiW8nw
Qk5IdPibBOcyB/xPIdisZdTAHWr1AjCR0ZdwKbIDbRSy7YDqYtAtr0J1RqIZu4/7
rMvZvuqWW7aHwMB4/cRVvvWkw0PKumTj5Eb49XOuvDeBP0F2D1JX/J6aWgPHKNb1
r3JcRIclGsDxfw7krDJvWBvJinpp1xaAzycvy9KxJBW2yFm4+QOY9GQMJ5VL+0kT
uv1KWVuLkIRzgHvTMmwG8NwMdqtto8mM3BhwV8jJOwqaNxmwZYsQ3j/PBX0hKi0d
QEDYx9DyefWBKwL+qi5HOUCYbWgAaFcjSDE5NqWgz7ilNFpie97WBKNmFvXD7D0H
Z3asTeARsjmEtItBu8+y2pofe/xJO8geQAyrLw5CN/WZZhUDBtcMttPeeSQGU8QF
lOm7XNiXlEHuSeamEYQHNG7kWW0w55poqCsdhtx5Sl91zRS1QVyspH4xAZqN0laP
k9tHpADEdNTwtCL4Hf+B1LdcaAUTwQv8ePZcehPJmT3g2iQN7s+QMmKta2f3MHzD
eVLmGJXL5Nx/qf/hJdlDwM4ovMdDsu63+yh7G3XLrux3ijwrJ96DOpYUOvCExTa1
cDkAqJs1PhptyeWgXmvtxn7GaC9MGsoUnq6/j80oGhifjqeu+3kceAOug4PVWb9h
pRmvMfxFdQ4eUyiF4Lon4nE9ltKZwtMOcgkGRQNyAhOx4LbyJFBwYKcAm2H4kCNB
EMbJmNDT9cJHs1HPsmNUVDbqcHwajzuBmAm+t4Q+EfU3uRm5OEFly1PG2l/KH26S
bPgk6h0Z+F7rbIrYv7SrCsj8/cws4uxKMTsyIVkv5X48RwGlAys2pW1HueqqqtaV
/cXVTGDZLOQQI3RTkv+6P3F7I12RHvjKqT0WBFMEyvi22V5Xb54K7/Y0SoEWt183
hio/mlEWbfgWOXaPZCqmkgxPZnGL6IUVRcQCPEiF3QqaTel/ZjnuSYIeQJ4tjC8r
CoMs9YRc1OIbw8qd3IKBaz0dM/5AkckNezXKLsSlZrlAYsrIw+Jloami84LdeOlm
2vrCzGw1D82Xjmn+gOaP1xm2zG41sQEOVfsLHi6Ic3ahCgeyzTfwgW+gwkjvjnpu
jGs1JtnebQXG3FLg2c8h6mHMXSxsqcjs15mvfsBRC8ku41GtMXjtAMDV8xYGwNO5
vC98SPbW9RK7Y4b+8g8knCLC1nZikeEGgerdDV76W8oFYLPeYVwGhqYs5tu7SgXF
EsdeIfnCCNM0/g4w9X24rGxV5R369kJibKCiiEYjEPeanuEwt+udlaMsa/kfs2V5
rk8zTVik8fbcZeBInncXM9jRNNjKXuQeXOvrbFQmzkl5sN8HPFwuQxMzYzFrncnO
7sFnT2Wm7Uv/uq0x1VYCpS898Zfi2YdwMG7vDYOGaxDvxrkulLXN8wT8P8XMoCim
1/EdHknIHCQ+QdXhq3/jscrq+LR0fReuMTZ2fIX2HIHgXXK8DOsll6QpjU8+qiFs
WGBcx4JYyN/JrqR+ziM5oJplhj7Lu+QwqTi80h9+2POoO+tZL16dMxnwhkWXJL4s
Xg8+iYZSFNJ53tznDABe4HA/kFh9Gx7yRJ/ucvLvEsLCMXzjwvBVhFqziyLy8ZtT
B/RXzE+6xl/niohTooaTh6RjAEO0m6uEMHTv88cEwMiuCUI/kSbVdx1Q9HVJorbt
ob+r8Wosu5d3OxZCzSWrwBX5gHw+OMxtcd8WOBheYkpK/ZBTArgip6otZYGg8/Yx
Z/sngifglSusIwWquxGmkj7naNG52+M05DLNYcp3PjD06SMYjfDHiQBL46q7JSDo
02TBp7+skKpxCsrx7JQiRiTfKQhQr0A1srEhpEKGXVIvzmDKKaZRX24rkQHHM3OM
jYu+BXPAyKFi1JOo6Pm6Lhlj85u/4QbPj+jgevUpE8Nh68u3Sga2/4q35to1Jiy3
2lsMzPNd7Ift2WoFLZo4VVyTEFayraVuAvuAvtP1D/QgLLs4fDrmFKun5dfrO4uN
YAl027/xHGHqZtdfa66UMtlPRgiQQcHhQ3QT2fjd+bp39tv4RTdQvrV9BwH1n0J9
fS98VVcDvp1RKVDJ7oEdNFz0qdi6/w+LSnYUZ8QRyh/4NbzApHIvfVX8WZ5Iaq9D
UEA91NOh/8vWVhe/iL7WA0e3GDwYvhr1B3fZiBm7NIULIY0RSGyva+WJpS4XPDpP
PtcwpWMyp9Zi/ArC1yo3J6BqutLzg4PMlpE5r8pZnW9FMAz5ryB2T3Oaq448ZalV
q2vQjYrDkwrXxr2Vllyxc56If4J88XEqT6R4/erLCgEIPFuLsQkcA5JmcWrJlZjb
T099pCVl6Vr7t9sdxfuuw9F7mABtt/BpKA49LqoXY9oJcHDhDcHCkEf8YSUaFzwb
WhHw7sZ51gary8HID5OWpCLvQDLTJdpzbq0/G+nxzmmLfy7xl5YAFYQLqzfQUvPT
2M7fSqVEVkDLfWobbpi3ujoOsIV9MFCg/pa+BT58qDSnDKWdwMeykdv/YVLY9onV
HllEPDwwlo/s2Nk3oJV+/lXmlQhDRz8ExPAHTseUoxq7kyWCS4kQRr21s+uwobuB
lKH42kQKRvIHOUsCAmS7uAmwCY6NVvTogbUrb1DYIhQKzK5K7OsxJTGVF4VJnV/m
4MfZANuirIZvQtmMHnJoVUXBAmeTyxGJMA48Ds3Q1yyEKtnr/2VYZuamqRG71O1P
3vtO3zozymM5JhG3q4Ors3Y4pKufZZ0KmasPIeOJTumHMZV2WxItXIanXzCEEEVI
jR7HV0AUNarr9MJSzWXbuduN3sQB4Ny+7f+01aaSu//uy52/uiY4og2OACaWyxOB
J+dr6lmcF4yincUObzKaIoOSEhZWzWVVlTzP+gVJxeijcXb7dCVZQNzdHch2EdXA
UKlPZGY1vYwqR0oja4zQcL64iQLCXHFN41T3xB4aNfiTMg6JCnYXRYSHUkTztHY6
S7daER0a681lJedSYhITjQBciKlhcAQXcGyVRNCPdnFH8GDg8dMoG5+wPfovlcX4
Ys9u0zubfSM7e5qnC6hhm2izhvfmot6QzBmvh0eTBBVz54cNJXbmwWWnxQGpnDCi
D4ptZB4YW1NIgmJ/uSxc9kknGjZu/vKtDXG+7ViAu4ToVOlbcglLRRxY1RcGKkJz
CYsQ2+fUWazTJrqm7U2u6I2X64HRYaylVGD5v/ArXHR91yryHbGZjojUOXWBnJtt
sYp5i+CLlKmWj642Ufgrf2hA78sBKEc+Qs9bXTraT4tc4dgB7R9fxA0sovWET41X
yfuE1Mhns0pb/5CCIBk2qQgJ4bPODx+h/VvMgiUPHVJajsFR4G76s+Y87wDL184Z
d7saGanV5qNuspsxi+mse4XzzQrdKIvUvNxpE1u0JN1yPvIpbD2ebql4B4tZ6g7r
pCOktZPZBdxfLv9Oesvjpem7Lg4O3zDGNAPrKrd4sUcRNjjLl5Ds1ap6hSFBeTYT
2WsoI58pJwDoB69L/ro2KP4YniFOnsb2LBiKlu3l04pAwGYxG/aJgFA/rfWsQM/X
qHOvYNBZPTO2aOmKTy/D32f++3+NnFea/kae73K8coZqdKwgHkwUoOxSrXazPmDI
tq9c1HgH1G1QiGp9XDOcHKslX9l5fwRSvjgREZGzCmqgRTTAfCGjO8F2bMOp6PFz
j3LM07K/f+iU/4W4I336l1M+ye6ADLSK+6xy417P861q16fuG32150n9LETeFVnP
ygcwvxv0UweIxDcMs7R1aqfYxdq6eIX8I3dU9ildJ9EhUAS8L9DiLrji/ISJM3Xh
GlN1aqEnmGE6CGAfTm5S8oTACJyBzwgCsoODcKLoKjgk5H8/uM3Ag5l3JLbS8hMh
xbE8RTjRKXXboOHg1zKxG0nvEIDbAEyviuGLle5ekg51Xpstn3Iyh5rk4lvTF0n4
kcWB+NxAHvBhOfWtRkxvVb4Wdn3XMUClQex+xaez8y6wrdB+7ZRqnSy1Up9RJRQZ
2zd8heW0j+0lySoVDpqY0JzAccQDGUXQO1gwaq5ckW7DbSSq8P8C5IK0SqmGQDUV
bRirttHOueBtaiygII4WSEJMIvf+zA61NUSlxwa4MYtUs5dZnAuVSaiHkFDuEesV
J5Q4xM40QJmgIeE2PozlAsqE/5j8JLtwtExyCDSyezRqRtrxHSpP/ueha164+t9G
/8C1TdmL5ZkLvXmMkGlE6et4sSs5DIEAgcErxmENcwXAvPfd5Sa9OqhdliJA4lgf
5jfU/8oICSumeJQxEqvIt62K6F5Aabv1s/SfuucW5GZUmuL9+I25ZYQ8ImhdwJKT
ahRDTnCt7t3MkitvtLa0Z9RsG0h7ww+RisNpZCdqCR++69oZyz+xIlo6euuanyqU
+T+9044JHwJzgpo9nDtO5ObG1MpujDjpR5eSAggzSN7sPFCnFG6k9yFAE7n1IEsU
fSOzFfiuFnnadcbDEF16iXmMUFmXG6+JKKsgcCb1vpbiXz6X2i8+IHNI+NnnVHiI
RDizfidc37H3Sb2hSUsfXrEVmmFcqk1JpEl152kYilQi94yTWfv3qqIMIsuTWqlS
SLNW3U0RorqhgOmP+F1KWZ0kp+rP9pKK4+uH2yqrKtNdMq/jQ/pS2Rxyvl9ICHo6
2yewyKewsfctBvL4qlhe5o764YKhRlRO0m06Qy7A3ssmKywIZXaP5Niff+COUA8Y
jUyasH5ISTB9ybEQTpuNHySJL6vv1TYhVblZDjbPul7eACalLcf8IIJVVQI0jlLi
Vu1iK32dDzWc62/wUH6BftY0cRKuZyX1j8Jd/rlNcY+Yu+BzO5fxXn4clmyqLmxe
EJYc1r40vBuPI5NZbpzKoQEsN54PjAVhlNWBpbL+ZNMTCGtIoj50M7cZGJWjTR01
r92lc4anGr91z5iM2+A/HneS9WyWPhFf1Okerx8e7uSNLRp6WSJW+SXTQ/4o508u
jmjwFM/CriP3Jm3H625b5Zw4TdNIZUY9Xu6/xRiTknVLEq1o1tW6VXeoK++KLfFE
iTuca9QT5HBDiGh8gPRUiqX65/oVkhZ7kkR/N0CBelNTKAj4vQmUnz1Cd717dmnn
eCf9bNLozsJjA56L47LAT7bl8WfBRi0BC8kUqnfihpYODhd2TMQ41wqqLvKm5dLi
ruCQ//i4x7cpl5riOYn1fWWJDq8N7w2oRCLFtHpEMc/Kdlq2wOqhddqKkNfIGzJg
ByqHL/Gs2gJmWSJ3PPX6tES4GWM3TFDNZ8BJDcRYfEvRsDoUo9kWj7C6ji56yy+f
7JiJZq9JEWf1eZWUv1pwTAjU15d95EDiNn1PC3f9oedWQWvNQKiaTgwNV09AC71I
CefeLsnSA+Hk6DF7qhI9aBpKfZICkb9YAYidZyhL1pOpnbN6pwRRKyrwt+1/EOVZ
ma++l1LBjSB1Zv0gCVvP7xDq6DpTo0jfKohO0mPmTCXdmr+1FhaNaYoTdNbO3g4R
YH3iOFm+VG4kggLc4ZAv3ZbNj4Rzn7zscbfkoUnFDgSzqNTMViY5K9BpSCDexvmQ
VtqioIUjOoc0MarRDKtG9KZ8GhIJ1bgb9Sc378DZpftGtSnD5s7hRvGMSOosQXAF
oO9U9Ec1cALtW9i8yKSllN/vr73xqmFYiVBuquX4D+jK8DgfXBnrhWVNBzQl7oQj
ASqjU9sYDMwhXFjjQtuGdEIqFKEoydWmvDBgy/BNURGf+vITVdJTv4KE3YJEUQ9i
alj3X8NmR0QDGLIDxE9R/Ml6KYF340UATTUq4c4IbKn/SKCcCQORVQ7oazoijdXc
Jox8/edbPG/iE96z4JDiIG9QfUnoe4UELR2XpnpVUvRqdRG72/oJw0smqJjPPxfP
UqN//gbpV8vqwO5G42TlIHH+MfGX7zdYU99NzHVfIsU/p3w6jWbPw1XHhDryOAlJ
6Jt5m9CpxwKM6JXane+3gRxVCQu+v4rA+wrzqJYEFDhlQI96VZGMXxiBCmqUxXW0
O7UiY13VZP5fyemUUJ8c/9Ft5fCHUZH0xPwn/CX/se3SmyUqLQ6P92051mdgvX6c
hc2be3UYdFzd+eszILLDiK1KyUy4oWNhmr34vTRUrXImNHdBMNL5i2aH0S8L7xaE
htESGuiJZP8Os2PIi6fjLNZegT20UVb86F2WvLDmO6MIkLFCSnV2F49g8JTRlwPD
ndeh0jLIAyJKDeJTf3WHIpND74ZeMBYRrDP6oUgb93ZTrXPDtVXzfRQNeE/9kNK+
9B8nN0n3/SK71ssVp5/GrotspCY14Wfj/7756OZzC+sEcEtpQ6kndN7qSa6pK+5+
ZvG4Zf+7QZDzPIk7bHD2jWTbfJQZGoR36ZdgKyhININSoCt2jEjgF+FWzDcbhr52
e555Dj7kGJkfZjoHDMFgb71A8yt9Ue2/4Cmn0fHhpTmMdsiCm3GCI0c8njZwBW8a
bFEm/d7+/fcsnxMMxOK46NrPG3NHcuZnN4qvuxHQjILMsT5l9OJVnLMwu5hRFNUm
2XfrpggSrCbHz7Wit4cEy9eQAPIgBJbhnbOlgFKZ5adMXGSrfMBp22gFPNTqu1sX
XZUQKUGu4NEO3q+TRh/Bbcj0D6kSTxmJ4d+/T8cb3uXKR9UPNRXDcnohBfL4yynb
Hqpo5DUNusl0kc904q6/F5dC+c179xg6Bb1SMp5JzfSannnQp/idjzWo8yrFR7PJ
mym4FtQPkXOx904NoadNTaQb22jw1EhwS9urVaTwx9qwzJFzIP3JnxfYx7lLuO23
4ZGHGJBmCvljYJ0fg+Yz3BSDhGb/cAIv7BDqlKx5S7QQjkc3kFGEfed9miH+LgpZ
V02V0qGN/FG3D52FhvMIo/Uubt8u4OTI2KX9YfA8j+6262R6EZWS7fnlxqbL0VG6
HtVw5oPbzoWSx/aLK5bWh3g9qhqmuFEZf23Q8gtZzFXe6qX41RsBYgjxAAkQiUkF
OzgwTpuIoDyeX+Rzppsi5OPysndjKZQq0BVv0xtftah25qUELDm7ABKZCzqzfbWZ
tGsDnYpWXJysv9JhIL+43Wp71UbmgKIsZGlzl2WsqgVgCZAkmaygAeE3fCBOGo9l
xW/vcTxnKzDC03cxH1E3SoTGKrijzZM8Kq2gNeme3M+ENzxz+oMcQUSPs8zT9uj1
laqodpvk9fBPBpcQkwQz7a01tuFhhcFsdSfAIVnCfc3A0pZSBaW4tfmg3QxxRpzp
qy+v2rNQ7ajNaKFaDsAeTi9sCdBRYPF7iPk7AYtLBBhIOnG4MgVEbEUSZfGwQWYQ
O+6HP0DJPMfTAkmkyZJYdryXt9pxO6gCsRSyIgtlSTou4qL27bB0xz93du0WR3TY
l3jBn4VAr0zDf7IQFmDIqVJQ/IJzv/fD2rtxhoINNjclkIyIpPN1U4czxGC9v/dH
3HhRwg7BoadTVPqiE9X/7CDPtUxoA8LNqBMHTw0OUKT5k1eCp3/0xjuks4nXRNQR
n76jN5Bbl/PZLtoUJ4lyw7mVKgIYtbVhm4BtA0ktwcrg97qOL3p+8zdFd8FGvXnA
SeX/2rGFJbNJ51faYVpWNSLpYXAW5U1TCGwP6tWZXA+nBQCXXrEn9kodlEILlLKy
NN8OCCZIkwpAbegIwCDWSMkQ+a6cAkasguF4ezFXMhk33jTzrrhNNCNa4UYDo4mE
R7ui9y701ZvV5tj7chGw6UBQLXf29obhON/5R96ecC1VQbMGOvmvmjt5AylPlQUw
z36hMW0fnQ9Oyw0GiohCS6Xoo5kaEK+/jsCH4Iol7Qx3u2XlKvle4wzBXwHNYjJK
j2YIJVWtKiJJrvQmoQwNGLLMfHPMlU2sTQcsiCi88Ux3dAFSP7Ph6XaiWVCbdYen
MSVb1kx+w+9TvWbJKkVF9K29tKjrGrESe5mdU2W3GcXDF1BRzRiVyfjc1+VoUPTc
64G3clY3FxZUZXlZCw/IikVnfN6q5HZTxsEFd0VI5wuWjxkE8vmNQtb5P7BWvHcL
FTJAbXFfWiwvO2laNaOcgjlL3fyXSa1oTW8hTVM9mvfH4v5biTzTGKGqNm8BrPUa
uU9NeGGNGxbDxlkyscDMIEjjFVNZOZyu1TGaoYWd/DlOd1xOYBqrZanBlHY6YW8k
nvhG8w8S+MIBWFxtV1Jo6Ye8pHrmbhgW4O4fsBv5EiBFixi30KDqQgLEgnVs4TgV
RMOAW8uYQXyMBHiygTN7KtoIkFthPtbpZgy308YxaXtxotQJE8Jr71C5/CLs73s1
KYHkqM68RaZys/WaXFcraWOEuHzvi3zZDdd3DHrkeAtpgQQBKqpX0rGwD0nSHIo6
CXdYUBydigGH2ecf2Z0xbdzzkorx2xGRdN7RYjna7porKVvQ7QSQQ2ZixXwuxiBm
xJSCAOihhw9v669GUNagge0mgO3HzzHw3PNmJUCRwSKEgUdt+Ez09BmvOIbC/ZTN
zZlRIDGPUyjtDoAzlWc0RyJysEemzxCHc9ollg4s3etYTOJvnuQq1yI8xLkzmeGk
ThjNgARSnJ2+mtuWC3KQQRKqrJ+lHgxkMgt3haZVMu+10FgJE8VxeTiMR050OeT8
OgaGgmbtxNZgFCdxjY82+GkvVujsY2ykjweRCGiNfdDNTUeEoW+jHr/8A/J1ixAu
P+lJ0gW3DQ/oL7/idAoKW1bo255F6LLfzE8so5vPPaFdvTaUJqvFQWspS5BLHpDD
sm+5dW2NKyw6Q5paQ6nN7/i/c77GosJgieuxu+VEDoaJ7GveEPrtjWNSnhY7urmO
T1Plu41YauOcQplHq9tjqSncMt2Jl0fQCm9e8oyZ4KwTOQ9KsZnweOnIJs52KE42
JmKc/WuZ7X1Eb5vlMClwTF8km7Flw+MQjXOwbo6v8l4dfCCpkO97ZNZE17dgkxWE
1Oej0T4nbmOBUfEnajSKDEf90eK9t5sj4JwN89yzSh6/acyrMmva2RKd1r6YjY7G
wUamKOSCqXc7GSjbZkIDqkwYidvFwQtOiilDnqhEbCGtNhHR1UEt5/77QjKqerjL
kgpfdwdgcQz7TaQ40iR49Ur9giyDg/vRQX4JszoEadCw9s97TWWvcJ/8cHRshOhm
1Q/oDgz651Lysrzc4ZHSF8c1EiboOSmZj5QbVYSVb1yPzCy6IBFWMX3dfseXFwLL
aUfihWiZTwNqqj5g7CRHtnJu15w2W+GtLIX2KOQutAtIh7N1IWp07kl9diwU6tdF
kPkNoOCTQTHvf4y/cEm8dRbyjeA/ZA0xes4LY7+do9x6D3bei4XWjrbrguLye7jp
nDSbAU2F/HN+/OkluBHHr5J3fUSuu2balPXcvcq67zLxFYvwTyzrr7tuYp2FWhkq
FXvXOt1/fToyCwUGlTcemX3zm2lGqWxX4tKmIe3rnBNweCVUNleZxXL2ewQGKSfd
XvvYu4Ivlm995UOrz+UJ1tuJZCwtw3gU+hpU04kxreXuuaIdkLVCXCNHwtTnz5fZ
33QgK4KNDqNWLn/e9fDv8p028wtmoJavdVaxXn4QD97TwqSzUTaoOhcWA0G7Qzt7
lnhrtmSzqKvz2LRxV0euR7WGSHKiXBs0MzrFw5FJyE4Zf8iV0j+zkE9ouVEWOrUs
EAT8eAnx+d02Z3/CvonMPYs9grJWxk4WRLzUaqC5Tx8XBegjHT+jjApXVSO1vcYF
GCnWbHcn5GA87cbeFAcmTXZqtgHUFpT/X5MjpFibn3NFuDvp8TscXJ8UUlSdh8Yv
wopVa0ry1Q9zOCz+v9p46d0NFRN7KFybeocM8Hmn3qAintDCyd3fl8FIHkg8uLfc
4zXA+JzhxRswub4ki6LWA6sESQTucx1mXLPg/uEgIOQI4Y+BO77lTsyFZgYtA0Nu
Fjpue31od/jEhoUsyguWNySwgPatIjDKPYjVt1GyvzMtwAsZW9+oGcNBs3MXPOxG
hj/Bv4D0f/saVCpYDn6PmmkMsVx/T6hjTeukKzMHyozbmiKOIfGmHIzZkmZy+0lX
y9v63j85Gf2FC4BgWYTe7NvGu76jBE0XbzGOlJVsVwfTrQJohY6SWTtjthihl3xL
ez+lbriyI3o/K+33fPOYUNbHgjspK+05zvO4GerxwTyH0V7zZ2blBMpSPAnf1v0j
4RzxZh1SG7XfQnXXs9kU9oavGUU4TuPNSJ9sIwpBRAlsAHJkADSB2qbAUYJ4uoKg
IC641I0RLXjs2D9gqDvhUDhUXnVD/K11usqzkxi7YjKF6JTCVMURm3UTR34Gjozj
/B1GErGmH1cWlRzSlLJgwjtulO1ANYH4uCXxkZZlBhgmNTrfn7aJwzLIenD+vOSN
/6P/5T+yBi0gRSaiu6TNvQ==
`protect END_PROTECTED
