`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aTif0CevwOyB9V6/1Y3RacHP0kLY6LK7FoC6VLgEcQMHzVZzsjgjOjgmtpFkI411
l2ciGdaHvOyWXM4L/8Hw+b/lN4OoBLPiKTIHguK5Xxqkw85iPPV7ujRXfPpUrGOW
rDfxr8Lk5TeUUviOW0PeCQyBYK0Cjoh4IA4MmGWD6ekXbRxf6NzTBYam8lBpO9QU
wnoh3aZuRy+GHPxMSeWPphc3VPaF85g31zIOIuOkc1XL+PRNc/nlWI3pPOVIvZQq
7mAegV6I6OX3SlVbECbDwpEbKI+zJTCQmYl6o3Gp744IgEWNQRYaEc5XfeBD4Hyc
0m2CFW2wrpovpkY0VzN4YQv6J8gKapc5UErg4mTQ4tVKBdlu+ZZCA7bZPgouJYzh
TLHs3GGpyMy2DZbpdHS2LNg1YVKSF88ABcfmcMeSQPJeJfkhgrNK4LNNLI8PBJf6
Lw+CvxEhG1Nc7RjZk+0mJUfL+L2uHMqa+IaCRF0PJ6fYyquH+H2N8WQr3xqnRinB
fzKA9ET5zul8lDQ9/QvX7GwKk9OpsULKfLWMGgsiz0BCmbU69lkM4kubu6NC1MFZ
EWprmSJphkW4ODAIJbxUDcWN+WE470dpLJLQ3UtRIHqyQzWh/1Em3jDzRR+GXpZB
MCFuhZHA7DnRW8TzJIX9zAASx/oG787kWZ+s4JXJabObcdMAE0zzmEDSAML7zv1Y
QnaYBatpnSx8M1UHAebF7GVzuJ8ydBRSN7aotKeHCb5ahObmkJ9aZJLBPr031luR
StFFd/MlnMrJOCWUh8D413+3VlE54fr+aSgI4cPJ2KiVgQBArc9LhxluIFhLTJpc
4qKidzXPY9apn4drn3+hDq64MLt92avzlqV3FOrJ8cRkYHcUiUpWEcAi2KLs1ynY
`protect END_PROTECTED
