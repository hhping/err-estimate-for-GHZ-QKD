`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R6oZmPpbKotfANyHynG194SNZ2Zu+gGgQq86NGqU58yNNC9OYU9iT9xFqFLBKBH3
EewVfrcAMVT+u2T7j70LLGUW/s890tQr3wcAbwpfKv13IIYccMlh5awT/F3Nr0fy
Ope1E1v9lcXQ30HS2iXFDiaZ/gFOMnuvGnwh1iOWIjJ1PdMiF9wy7qJKQ4d0GgsP
NpIvO3SoRMe94Yb/OO8KAjp9dZT4X3vZhwmrl8Jfir9K7RNqSyx4ZQAXV5HBnn8B
nfa+IHxS8xWc85Z9WLFLEjDD/MV3KEc43PlHyDQeTWettCTSF0uyM4AW70U22Vw2
rYPDK/7Hkcr3sIfzneXrETegB4tkCNffa34Notd40roFGN42GOnhE2SclQ/tTAxU
f4h+MRMn1Yku7TkU/us2jreOqaB7XGfVwibw/2fgQ5bNty5dAVN3E94etvJqjjtu
017AmlY11EdHZL/WRzOpartBuXnZDM6lTmJHVmAGMzUtELyFIQRPLRMvpY3oi3xd
oy9uCt1AvfYOJLMdN6kfhjnsLVMIKrRmSk84eZaIWhs=
`protect END_PROTECTED
