`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
owHc8dOsJ8SUnGCUh0n6qv6Xv0/pz/Ay/D0T2XAr3RrXkx2+mCdwLnjQDFdb3cr1
BbxaJyfQjGJlgevK94kQdQ4Pljkwg9eSWFFWDXx2MaRrtNZQ7alLhO+1ILR/E38T
vKYG35kSrjMA8a6risKIkyama5qwjMIY9W8kAaWvk2zqBxphrExAwpdvQXDMTlup
FQj5zFhgQ4d4SjdEzMFnk1MFSjuKs699nmOIb9YMJLdFtA/No1JpFD8qh7LH5tpC
jttdt2LWMrwBwZpE7mRAIGpYhe5lF+ZioOc1gp4uY/Kz5VW08QiyudBkODlYuHvG
rGaQSnQE31zqtgexNktMAqD9+fqaK9TlIhAdpFj7fEPwIFp9RUnsoHTkcIC086Ab
oXzJPcbkVUUizGzKrj9ihjbS4AUsWSyiHJsw8vRJ6f3cw+xqGJqSuj71dVp0SGoa
Fal9TmINsmS2RYonx+2eQQjSRwrMJ36pboo4+JxjTntGnYDtqcr4bAIuYwTGi+wt
rGWybLp13ws6Ir0YPNAG1DqKUl98kp0KMEThukCuWvVdj/Oe3pURsrRBEg2PhRec
EIz76F0N8+egm0qrlteo9ZeH8Fl3IhpGxOszkgENKza1xESFsaFtAwN2jZy0Ouzn
kKxHcoOPDdDQDr8kodGbvBEe4hfDOgcyXZ+9TbY8eIDymVITwW+EEtm45x7TvQaV
A/ZWXtxmTuG/h2HfajHOIRkfTSklCApA+1L1Qap1509oSX3eT1NiDHSwxxGFiUgM
`protect END_PROTECTED
