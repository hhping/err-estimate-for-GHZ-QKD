`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jpITmB64iOietjMH744CRPFfa0GCAeukr/suUuOM/zJE9Bh2x+thMWxLGGx4WSEl
yPjeQlnC5U8iUxksR6Cyqa8R8MGJbgS6X1UXTeN5wzF9IyntoKd8cdM1w5tccbJp
Ac727ku4SgRftOwS6qzJBSf2qbvg6RevgVILNmVF8v7JXOhaLQzGRvyqIQPv1FER
6ZhENwE4cvIJ/UQBcxGy2zIXW8DcqHpQGTmlLJf+2eZLUnKYzmirZu1CBxjCiwFd
OSJLt4RMqhh5raRzblG69HU1/xZL3yRUQwr5PMP8Ocpwp/MgFKaUV/mez8yGSnQj
RLcR/GXuZkJyL19X8RZGk0eEaZtyZZPxf4l8Pp2G2oQHIsGnScWTTw4ko5yxzu3U
RtKVU1Ik933ptHE/ga9ONAHErODAWUWv2FSSUY1atWUl97cHwfijMM80M5QRBCW9
JnF73BxPzUR3/BbmjNFZmRyLe62tpOCw/Rap2DknpR2S5T1IU+L4SYssQYflZ+Gx
eR+BG9Jyf0WKCTzVsDeHy6/U533E92JEU4fZ7zAGoP8fWqbsNa9n9NqQ9QI1bhe3
0MK7p13jgXAgJcm3vcKQeK9AwCQz9d+s2qrvxcwTpmfdkxcAil/xj6MKnTAI4qvb
1/15+IxcgIdpXwDmDAKQdV0SfOITTX7c+O0PU9NHBFfIBx9hpOtenbl+cvP3pf9f
/gsrMSIpqBFIFTWGelYAiSy4C0YXEoyXYVktJVnwnNQDn0exVAp2cpnSjIJ+3RP9
0wniCQWJ6Nbzx5ndFHcwZPAM0pF6sahC2Tt+nj0mqkONY5jcU5gZVstPByvQtiRz
eKQAXdHo14AtmNt0lI65aaaU92xoUsu2z+l4so2pKZcKtjNWMW5jTdBjXFIcft/w
/bdgOup4P8Twn5PbOlQfTcRAGOZbHMOPjYFizbsyX8KLm6NXynng3IuvGIEkGdH9
jvgfoYRfkuUAtzZQxcs+J33DH6n4LuzXXZ825NW1v2zRbv1fGpm1iI2gl9OalUY6
ruPWjj3E9YbNAvq9zjUFb0BxAVqDsb96aG4wv0T7knxv+HWiIdP3lj0m1q5g2bLA
E7yMdnkZ9L10f3pUHD4JJfxDFugHZSS8iUmz4ROsIOpyZ6ui2geF7RFzBz/77U2j
B1et12b6XykGPAXJ10+m/xnnSpKsoUuaXdr6053iuZGSXc9/H9bD0ClTmTX6/g+n
xoxv1r3SXi+hkvx7heRTqplcnhgTv/8pz2GFuulqRv/bGDHEkdHRWt/D+WJAQZuk
mRHeQ3wQ73o+iUZxjz1dgLGyxnM76U9sBIEvufD0TjottPgPOp4sk4QRgpYfoxjT
vntTciGwNf8Gv6XEq+iHF1+isfO3N1BtEVlDzK6IfTntFaaGEEsVMl469Cdsjmn3
ssY3+SABJTbPCeQ6EG2CvOoiKu/dmp7J7ejalWV3HFvSFSG0pKfQTUMxmyVXLYhm
XyaVFtuVUzY3wWVIJIrz4W78lxy953g1bJj+07PzHLIw1nX26XuLPTnlWffGbOD0
qeM8R9+sveXHhdMgsSc303TxiYBkdgNATITwo8H1VPRKrW+lH3oXPl3LIrumbiix
r0A+4dPujTVbHPdXaymHX5+3oaj9a5TNwru0m7mN5g0AxmCsQOHN+jWZfC3Ta9xL
JeIVnRYgF5DxCybk3M4UMtdP1X+LTSnr+fs+IvQMXxlitW4/LqVEsfZWk/I7pXzk
JhbQt95LOttEbiGZKn9ePHAem/sRkThB34TrP3FSu2D/fB1TCIs9aRsOdjVfRjs1
D6c8R8n0BpYaXCHrvTLTf5IGjz2Qu6fOctTZRQ1pAGrcKMS9DYqU+CsnORrzNX5q
RVHHoTYM8NTVy4CqkH/qaOa2NwP9gwanHjkrtcf3LJk8WjN++XoPLpUGnfbLBa4S
gDC3fq2KaImgG6ApJ4m+vVZlH4ESUt7D2yffIIzBk9nBk0/90PKZCcN9DXQavy48
2Z7S57VZ35hE5aFhn+CUdKxjz/0a+7doYnWbjffI1wT3VVAMdZIKfiJB2iNHdqIn
pwgQWiSxgJgTGFnn0SYV06KWDC8WKjLEJSno3IMLZwToEEA4VI8DqRg9ug3vrr6E
yquraHH9KCMUiQxf50WqrMowNXSIkcWVWM/aMIleEEL6ffm3S5YrgKBqPMX+XWUP
OmgJPhYxC1SOBRmM3CJu3RfdaTziL275EMwqyZpt53vZwmrsJ/g19Fwiqp8ls9Fp
gdjKpZEdBWWQ43szd/fB9osSBA3zjEdJw6uTq/8kTGSMr843ZQDXR4YFjjov28yX
NvDC6o00FQvgXgGWp08RvStorf9whiXjKBtYNVAw0yyaw6m7n8oy/OfeMQub9kkd
A1mohHElq/aGWmPI3RV3o8oszKY2SEdiXalKS1ROq4BTHCNAcI8gHjB7n0VJdnbO
rMOjOLDIWbR5xK6AfWB12yAT4GSUSX8eAizWBQHFoTle73fP3rHQe4lxZkXbxxk5
mvJDuzkAgeRyp30qVTMYNvf5teFXV6HNLhpEwA1aeE2e3HcUtIHX8u6agh7kAgzt
M8MASI8niW4p6OMEMAbBArBGsMFWzyP6X4KG3Inq2sFvefUlMiM7f/WwrJ2P6JJm
NEn5nGxFo3UFaW5BSTqjQNLnoZkEiQMy079rbg1T0I+feVJyWcrqwqGJbJa3h5ox
aM0eaQzpqLb9gJVi3xhgpv6/IjVmdoqP6qpveBCicI4r75p+Tnkqw8OIlKs5iC2X
AKL1qRXjMw+JiSgQlwajCWQqmDH0nLIjMt/Fx+PE6qx7ap7qpW15B9pQdsdYGLg0
6D9xeoxJrU9aC7J/CXsTbv4EnvsMLtyqkQEm9HpMpj8n8wgE2Hf4sFPZ7jjQAhrj
`protect END_PROTECTED
