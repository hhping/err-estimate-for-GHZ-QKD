`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pvTc1GQut12xlgzi6wK8Xz+B9vn70zD80n5fhbVXzCvLQ/5jsD+hRAgo0fVxHSko
5LRl0U2oWI1ZJKPhhnZ053z/mw4P+7AdXyXBKk+ZRad1WTkWs1BpLJbkXhJ4ux0/
jywtfNAf71VK8Pph0Z90npJ3HEv6eg2IhO1d0BxnI8YiG5BOjWY+1yCqVvsuE8oG
yvsDmH9MB1G94oF7hJW5YETFyQLePqNtcZEgBRJ3+dBgdLRDFpgF0kerWHp9Ct57
68kLRpsqy/l9iX0Vi3pwCOuG49S8pAIsCAnZC1xGSnLuLolQ8maulVMs5+QPygOl
lF3X7Pp0QZTKNDxUvw7qC0tGLY4azfaQ99dBlmB48XNxsGfdaQaGBTMYA28OeelW
PjvzMvfCNXFY03n6Hpbm9b8rrGIZ1Oesv79RLGiH/a+MDwQ/oovCGGbINSapIirn
/amGEyuGCP4H16at+Zl53mFhMrpnHGjYziO+HJlScn7qbhXJoIjt9od1twjkjx2h
qSZ1Ix3Istl1DNr+6R514Yj4gcrZ8KioSeP81BijZsta7HcPIS/cklP2f5utI1+I
x8Bl1VUdqE7wojaB0SmVRMsKPElqaaeM6iirjTrwE7Z4LF5MSJ5DNuQo9RDIqg0B
Ikzqql2++6l/eFW1CWIRsNVhjdJ51dFAdc1Zy85qopfdW6s1R+D+7aGkct7tmDQZ
YJG5yfla/LZZ6PquLWCyAMM/1dm2M78En0V0PqbUoCjDFrm9MHCCSxX9mCys685/
myad0pGmdE1DxZ2swmE5rs+YwEeFQ4LgiMw2RqV8cuy0HjFO9RkSWMYadA5sPgfk
oTR5dIKpsUYqgiAMi+X+aNzjhxNDzVsNxIL1zcmS2liEP16YYXVs3AzTNDLwQzVe
R2eT/Ogl/AEctGSDGfQdJcPWppGFemrNYZz/2ASf5BQ9Rj/QXPa+avwkhIxniF4j
AySd8vkMiSKxEfhqp9v3+yJRKcFcCujv1KpYrXuHvYd0cHkLh8Ab4b6zvPYAetfk
jcBUwH5PzVXa0Bzi0nqMlsTPxEW5LqLq3KCrgk+3e4jgldg2TcH1RrlzwxMeKf6j
ZQGgbMO9Q/9SO86bkZcoQaqiNojrwsh/VBU1Tbx9uZUd66iuCkZKZ3LazTZ0nlUI
4vYUpyN4froKWUxwavHX534xSaI0kVRqhO72jFFAIuWc7Jn5Inn789lHu/MY5BRC
S9pr0MoiMGL3xHT3rdb4n2KiMD+vZX5Bx4MBN7GXM2H3rOq5bfZBg4MjJoWpebfG
OU06CCLPYASQuuagMiI2D457XW8DLKhYFrDlvJrIwy1v0LWht5TQKBAH6TQBAcqV
YVOzuE0Hl6n9yQrtwlRvXyZxKKrKzGfZuuVWmAhPnCgp/4OBIOfVQqMetwwvsFzU
wsrTSbZxB4/LJf7730EM/+SS4XNkp9CbeyFil/6mi+jpqAGmZEg/mfBYBX5ljLjk
oD+Qbh72XVjCJgZOaVpegGAXc7n0UCuHY4+vWgAOk4Eui8m9OBe21BUOOk+zmgxC
nCCcNVwZpuIM259VhhorNUaQgCFFPpxArK2lNDhwEHIs4APLaeZovSv4yqdjCAkA
T4VI1a0eevNUeOcfigGjWvqD3+6HeH5krYiZfRtueID58jmvmOtdrCm7qr0aZ5qL
e8iB+nD/sLq8qAmk63+ufsIlSPRUJ7T1OEwg9/GUcdqmEzO9o7zgzae9XMBoB6rS
be5eMWqkBOkTlbdjFUwoFdZw2LrpgifxfuDlVAOB+rDW/jffWv6ifExMTVO2gg7t
T6YbIim+XCSenxneSrNfIeTaTDBSBqIlXqJRydXJ3cbDSUV71K6WRRCwVSkVr5+o
SO9SSYepXmpmHPT6eWEmBifkklVP2kC3kzJ7H/rSLFGvEsp5sDtUotXAeKDnPBcP
0XXl/LBrFr0fZChl/1FX8mmVPZ1Jv2dE73wReHBQMHLMDMHh2C9GVBdaYMRYk9Rf
tx2ahzqfgLz64xYQ71lVufNDFCPLNriNMhKzp77jxOUglVxzq+R5MwxVsIeu1lFd
yM9rw1gXsNwqQ9oQkgfiPZoc+GyymgI/ybwZPyJTjcUKBFvm3b/+FKJU8gQ+IxEx
pDmvuMgXisrFvTS4TpiDxwTrmHevsFAwO9tN4pBPJ5O0bGQkNGP9efipTsQanQrx
0xqNWh8kRdcmYP/B8kqTZ7bv17cJS3njY0Mllt9xY1P79OzKFJkVfObhVkZiXpTy
qnVlJUuBXkwMhTzxmlfkZ054UvcNgHRz9n3KSXCFGNonfgSK8O2JvME9ztcOaoqz
nsV8bAMQ9YfVQMTImEn2syam2Ii87JPptkh4n1mBrEFXJfZUCFMFInB8rBxQtWYi
XItOAF/mJzDLKIvqekwNzTTTGFhYEkMpVUrz6mrbxnLPDneFZ59UexcKKIp3OM/h
QE7KVq9XglBBBH9snvH1/6+gvyq4xAnibt54O1I4rETgD+65Rv8i3B6YaTqNqQFo
OZsMwcoKhWS5DzbYievlSI6Uhal35angzRsperWzBhnzRsuCmyn9rT0/UL1EWwV1
++d4ik37Dm0daPOPsfz2aisQaz1vnjQ+SQZZtaZizmfISyWTdmLD9zEQgTFVNRwh
7VYGwQsY9kyptRZKHPbRRNvCupM+CoaX6mp+x5jG8BcaxnQe4hsFyU4fWWiBYqC2
2iYonk/TFoE0WOFKUGYn6LzXRMkQEur0Ts2NzH9s2MVbbMjO+LdzkpxzptrLplW7
d4ZPp9rCz5QwpKEcKmpnx08UTZg1ieoTXO3Ty3ID0KNkG4PWKtrG3w0/ye+z0RtH
TJ+is6iG1NK8EpFX9dlnD2JdDITPOYdEX3Fph+WC7dPzGLni6sTMoX4XlaD9Di8c
6bDXDNHiFc86IsfYzRSWw/3GN/THxcKReIV38xDRzt3GMPA0sGLKT4uUbsjH9GKm
AIkZYURvcQ3XLmj3YeWBhFzJyaM10VYaSfsYsSrGQD5icVZMbqlaWGOeiY7yugYJ
+2MqMTdn1KtIZWDE5hGe2T0YImgo70L2CRfvxcJGO7s2oPgebk6h4LFJkJuAu1Rg
eqvR0+f1ArSsG6UALoCyC1RQXjjDhiLX6rOW09VZRp04TOGfe0lXVVb5cxbRj+R7
TEG3PeMxI1G7q7PsL54V9ijIsm/fUEJ45RGmTpbnh+QGyy3VRB7oTc53tNDc4FSI
WYl6UjntAsJFJMsOwpLksz+uh4/jm6+0q4uke0nw+JqT8DX3xgptuy8kIESXA+wO
7eUO/cm1KyOAvxfxs4pbDqBwsy9+awSFUVmGJgcnzPqoeKqwX6sxfw5vR1Jk9cMx
8vc1nTb5Vd7oO7bk4AjSDveiHsbbEvP2jyY0ksa/QXYXE+EcomjA0nzwNxR52eY3
K6ghldJN4w+bX54hJDL5F6mJ9iCmC6KlWvGNVS6t71K65qEQWel8TheStpgAUx6E
0x2lyWWDbpzX1Xpgf/QaxD8rgpfx96yvqhL3/aXWHWARwUAllaR2AvsPzzZ4fGBm
BlwG67vlP8IwQs+qqP/Q/MMakjmx5IsoJ57INPP4D6725Y9o2/XmgTFqncFeGLHM
v+Bd6gVzK6xLGjLnoqus1RcdhEr+GOLUglkycrtESjUfbNx57zuoPatP6d+oSk4g
HeMAmfjvSyyNtw3Rnk9cbMlVw84JF9TJUrDwBjKy/KGVwooafVKe9CGu2pGA26i4
IYdB8LSQM9iTVp/ZP7E0xa4wN2/pwqA8yL3MNY81XdSKDIkYCBqYCNyLR8+6P6uf
YxdwDhNd54egBr1DruVxSFelYNXxarE1QNlZQc2KmMFKrsonuChZAT/2L3Jtxl3d
Ou7R3Gh3K6X5Rcvc0U5ZG3n3EO7UWXHU0AP7yYZwWWD6kASAS8d4q9tSBzAUrUbx
90wZUK2E9WdvG6LGA5seZ/CrF6lPldqFI4mkgChmTDHhH7/Jt5DNGmuZFCjJ/hzG
G/f0QSeQMfW8+lKaVzAA7SU8gR6asSRVC9CVon22LFnnyASgMGwOzIQTuuTa4PVR
aCadhuX8a9uRQddV+8d5tPLyCCBAgh5D6jaykcO13ncgoW0qs8+B8w3voda0GFWR
1b6I5yOaTNEp72WK5T/jHWbX49H0frIt/OzUEYjUvdtALukyI2z2+1Z9uaGu9d++
F0VtAuGeke0uzuJYuT5jpnxGbpOdH15rySHhLPJSA9pyE1G0IO/RTcIo30+pn5vP
3MCgNCLF/WRSRDvpXnFkwVuO8jggTc5rMnDloH+9GhG/tCIAzsXYxzGhza2JsBVi
iNHbIvuV08vzO61bSqqirgacDmaYxBZpxX/nEpu8NERSWN4DjpWqMr5SZ7P0PRM4
EQNXHoozTwh7E54GZTXcheq1YJqJjlU5uUl52A1TcJfOmgwi0W3Mr0MHuN2On5DC
YJ5rabO+2LauhNF6xLJDE8GO7+ddAW/cR4Rigix7BGYxDliVdgebMKuZzSIFsqJ8
ijsVntg+5lXb/sATbu7JwY3jiqy5g2JHtydcTVqsS7u10GjDHICJoXCv8/Ri2e1Q
MugZWrx16GDDX4DB2J9tWcQjFcuEBODGX9GJbZFQeoqug81Vf2/b6GMefTN5YCvn
vhegqnQDS4KHTgd7rU2UbnS0GNZdKEa8n0CCXGLRz6MdIfZKlv911yfx5KLuZ48s
Lt4mpzkTPHeWbLc8uoraa3R9uMfUDGTafRiSHPDkOqNtnPYf4bgfWGlmB12VBWHl
yELz2+J4exSEXCR6OZrqs9+8up8bXmLVO8B0zGSYMrluZotIzEGUMi0RaRWEoGXK
YlsepPbHqsu/S9TY7iGdS2CcFRQG5EUitNKYkEkyZNChcvE6QgWIOuMV+3V30Y0G
OTrAbmX7NT6GoRvjue8adifVIPMaH1+bWHdZPmnZFiOqhZea1yZ4BpaqJHIc+a/n
kjZC2Zri7sY5hFYA6GhcBrfmKirQa7ubxchb94CkjA/SQGkN6ynEd8LaKXIlXEfF
v2/Hv9DTnFqK84VGLHNnyen6wuRkOhFsMIy3NtE+XIoFip4+1ybjhoPhaPko6oWZ
vJM0Z2FxnOUePhIwOlCQXDKI2mRD7UM/AjMw1ikKSZmckFjME9XLQ0qxvSYZeJQy
MUIrLaEFlwXRoXqLv+EP7bH/hp/gCHnS/TYw3Rac6xicRg7isjOpfOjrQguUQPTD
HSp6N+GuSinwUgFxmvpdsMyPIUTFpb9gQi1ybPrfweBjEZRR+pI2/myswk6YEZYy
YenQjraXdRHw1PJyrrocOZGKd660JKnvFReZ1eg5hTNOOBbI7CwynYZiHIYnOGBM
d3E8vmV1kjGkFaBkR7u/Svk1dDO2p1Ich9tkbLGOLe1QT/9K7eE84OgLe0zgUVIv
riLdkWF7d0rk28YF+05NKZennWBTSaLiCOymXmPAnoqfc/81NE44uZQ8yVueYNVl
+ZKYLgy6M2E+jEYvjoWy5jyMivNoiFJOoO03ahoZ2r4knuXId4ZvAAl9lk+JpmDO
1v2vSCwIw8nI6nkwLCH4qPcvWgo+VtcEwT/TraXf8nRgym2LIfKbKUe2FdaS0eCf
Bp6biPER3kejhjN+X2MIp+wWh30Mib+7MUY5Ndvz5l9N8Pj0BjYv5pVZK78GQxZT
VC9JdbHU3LHklUjVCS7VBpX0NylQKO/dNDFSL3Spw8so1CANYm/Hsab+ZzG7ouZj
mY8uBJOQF7Dvnduxidy1/2rHv9QhEIKA1B3dFJPlF5XDv4X3YorbPkOfW8NG15bf
EprlaTCek/LuB23VS+8II4o5vXBBbsD/jVzKZGzCnrN0EPrmDlAk6iS893CWVpup
vIWXf8WDYGQiVb6SzuA6dHqQkk8KI29o7oyXakpliU/BQfqiMKdYKMwjzxApaepd
SLe3kRS88NMYRnTkWprMcDOJgd8xwMXIc9ZPmZ2y83UB4MOXoWlfHAx2NjTAZdRg
dJZWutyWCxQQnIYeZtyLLHsstY9BIFf+tRKyy0fGuE5UWU/YhE3GothqoWlZC4Iq
r/BdJykOvTwn0WSuWvEzhqaxqm61R9BbXuqM1cls8oPKhryEyJ+U5U0WaL+P8Wzy
+LyffBBRm0suQgEqx07hBt6JDKmGEfZEycXOEw4dsQNqTh1aRm5FZoSbU12A3WHg
oxkwrihvlKuYi5pshvJ2snqrg9gCraLnb7i+llX2zJRVTU3UohRAT0vNcGbsiHPE
p0LrH4pYDJMed4Qa5dsejVzioBzBlC32eDcsEgQancUNSVESp/Q/DJ+zdodVk2GB
N9Q8vCGIVSLzWUtNObX4X04RF6TW67lxyLaw3IHAT5wTadcffxJ4RHemQ2itrMoe
seumVuxpq9ABEuDOyZIb/TLpJLxJqyQ6UnBKjAVUmxsa0Twt3jZk8R1TvNnlIe6O
RDiPTAXF0tfoNVWSCv3v45Y2aeL3YTfiGa0hkEARftMDJ0EEE51C64NxiZa+tLJS
SRl+nuQ2OSPW/CBbWbFLW5uwFJxd93JIun1wSoakvHcHV1xSgNcWJcdFFYA7rVbM
7+LGQZVsVg6dYFBWqXmTQ48tYv4ScPu9zayAQM9isVIzeCJotd+ycC/MPDs/r8A8
Gy4IEfHfWv9PZed+Fkjfajafqb2CIJHEHpYTzm+7eKlRfUOTPfUosLbmz8vd/ta1
AGBdUNQhRzzCluc188CN8BNeUftbT6gaz3ZmUw1sDFF5gkK+alrzbYLeZKJdkkQo
isp1F1Cj0+EtoLKiFiDo1WCoq+WnT6WtzbcNjBLTTMRErdEbL3dbRxKI++FBAsMP
Y2bZoClMe3a2OXqxUel1rVceblSZLgFcWuGKOXmzFEwEcGpAuUPui7BN7WouLXtW
a+Or31GX18g26qBwkZg2D7XrrY6J6xL0JOvWiES/aTSdPmpZ6tUhxz0vicV9awcw
ChG8+O7sBFHEQg/TkI5XyuxkHiAEpBwE9GKK09V94XbNIW3OxRas5onEN2b5Vqat
uLO+WQm1emsf8/zNR0pMVVjG+qTlN5nvPwyEO1NVnmY+bmtfUB0LhylefOoE7NyI
KbJQGYKy0VrSDVvtkHJM9RLlJMPr+PPtx/eyGZlWw/8yl7pMLNuwICeu56fZer5w
7a2UQs1nD+2sGbUBfp/DgmNnXnkeeeCPvSQiFg8XdSzmN1QL7LAagYfvZMxy2G99
OcUTo17jBVHdS2yQ4nZWgh/s2bpFVRFM06fw5lw11WouR4Xo9OX/pAnVnFm9GOvc
ejqFEFcsVTwnZ3CZpjaMkGdvllyHo0o0IUH2sQJdYZXpaJGeNw6SJEZpCcWSO59f
fdczQve7Or2mz/brX0B8PvLflObocrv6usAER5FLROuF3fQjnTKgvl5yoe6+dxv2
KAUh3uVY83d152N9acSy/vZ6d8Z7YMKvIDS2KJMbgIhVoGGS76qL0dOxu27K6aCn
1oe/dJusr3fekl4MW5MknbLB7TmZGkIXFpUhLe04YiKdx0COa1kQOLtCdyeK9ez4
80nTBwdpNoXX30RWUWie1ateIEpArdKWMt1OS+oTw1UjHg5qke9jYwex8ewjRxVl
2wErxAfk/QdSN1oUgeRrHBAaVRFh2gQv2es86aO9rb1pPEAYOxk3ckGbdbmGC49U
6gvNLE2oEU06ZJRlHCcX0sDPqBVPUuwIY7Gs46VyFf4Um+5/FnhywiBNEZHyU88k
2WBxj4kZESzTE39AW6VUVZ6Ul9PMT7NFpyTRRdtGEj4kxxDrzow5aK27IPryztJF
c30ryBqeLRLogpifi9mYh8AiIdtZ2l699MB4hQiWcy64fewhGvU6Vuaec/O1TSTx
oEiucHCEh5wRWl0kiBTWnZAbaHJ+TBY3Og1ApPA7K7Mm/obUGCvookys6tsU5TZd
qmzpousEIK0EcceE36BMXzsiunhJKqJQSlkzlCVLechm/RWdNX2zSwUsHC4eW0qM
4hZMV9bQqhjk4v71BA+FqqjEXxJJnSbIQtA/f/dDrSAbVIYs5wOa4PnsJLMlk4Dk
vDBu+4mgIoGwCdhmnlY4DBmURaGcVdTjvwt7pI5lbTY8H+zV4its0VMFbgkwQu6I
6PBijygnThPKOWXFtNHI88Z3Ak4xZH7d1bUHzW7cXZLYinvMnBeXHuAmpXjsOsss
BEIzdEbgqvSOqFFhj29ZXbNbE+jAwebzVUaEc+NKng2dk2Hqvb2kioBbrsZzq2gR
9U1k+0Bctxv827ZHk/Fw3VkGsnFkUpTmmkZ81/PrJZB77aXPC+B0d1Q7nOY4umpd
o9ouHboJBOyRn/1gRWFTHys97NlYIxPTwykPzF46ok33WZF10thUdXC3XOpqvFjr
gbxdkzQhyoxuU+VnV/Ldvak3nx0V9R/nqVQ1Q6bDGsIZ8OE+v6AgGtm9Jbr2NGWI
TC7dq16Kh+8Mvus3WJTniN0DKlLyydLBPRSoa+dskI9lisqN3iEcqB3gaXyQ83e8
yHUNmerJcLnCUrujmvPIBS+7+s/NUAKd9VhAyyBUaBRGbFrLVRXS00mylOGKsw9u
/KqsZTlYh1CCGeQru5igDl/TKlKV8knSOHv+Ni3+0CjQ+Wo4xMN9EjKnnnIfab5h
T2ZgsZ/C3g8p7IAKtj2Zn+eFRznyxXKjX3nGlerDj36tMFNiN5U2Hr6niIapDrep
DwEl3UvKRyOEl39ciuzacEQ5ApccpqT6x/fcmUK4K/1A02nJks5Dmwdl31hp28Zr
oJuv9tK9DA1UfuXJTqADbY5S3SIzcgxSgHIfud3GFx5RX5Yjyh+FSiOuDb9DeWd6
xxoz6GHMoWebP+Ofkk3AdEoyE5dPnCKdtELToQDhwv/E77eVwHHdYd3+PboVFQJi
oFJxRqc11VSahJF531G2VAbPKqs8beDDmJwpay+/e9pWHFEhZODXiBqxqpHDzTel
GKDajlB2BLLxtAUk6BiDvRwGK8JYKn0c+kEPKQJs47v3TxTASrcih7R2vZq3PxCA
CCOjWVhsR1k059rmuC6ZKd2tnuemODZhB/vnyUC5WQUFTzVJsSEQZceUmta416k9
y/rtiDLcOaQibLKCXX+j3SMtAJGPRR3Kib5YOEEsc/q/smcCFg6A8SA79vMGYTHo
SVohiZUFXLe2SPMSymeoqTLAQtDB5SZVBgexLxAcTgzTH7tFk1X7uUrcfw2DO8xy
98RcLnK1IenTjuIbuQaCXdd2hUtSFpbFHbUYgwZCtM7h35+TYDC8Xx89hI0HLAnp
h1pk0eJwwts+geA393huoWoj1xjdh0xFuek1mQwQXfwqJ62qlwfZJFPjvUr8j5LU
2IgeL5vD/FRixqGCBGWsHhppIBtVDxKXqYdG4Y84SXRcuGm/alOpdCZPo2cH8dUW
B65RMCgBSGYhR2pAg9cYD17r+LQN5R9UzjeEIFub/GIqVWJOgUQSxVJxcKrt+IwM
69D17sICl0515kS6YXFMKtTOTkMmfTYlkLgCLjC8dTdwjLmojhDjTQEW88ScMB73
7phI6YD9JYzalJWKcdSLi34OKvqSPdeZvJx7wTEBdiVnUPXEIo9M0vAB+6d9bKOi
UgyqeuO+WMW/z5L/b1iBzsG/I0qF5MXW78bj8pev26JbaNc32zzJs7Sr2XA+ap7g
UQrW49yTQWCmDBMp18bHKDEzPOygbj46vuvfA2LROJa/VOL4FUJ8Qbi4nKxiTnYd
NYDmKE+kDE7xlqx0wlj04S7w5ChhgWqvbt6r3lA4Zq2LTVvkfF8k23N31VRwlpHd
SVwAOa5UlG5Ufkl9+qUa27jaejU/PHBzDmeIP1451ONSsXwtiyuuseFy2ZYKK/Wg
G2qEaB0rLaBamMicRuicb1HFNDo6/SkcIAAAp222YNavT4S1JvKS9Tble4szqAQn
VQKNQKiCu+VzcZGAIcUrr9/i2KFMzHuej5g3q3nmEvg/FIgWurB8iFZ5kgC7Q3Lf
3trr1ax9g5GRr6zP6VX92hMMDdbzox40w8O+Fk4ykN3YbxlnAr0GMV3rPc62Nykb
cAWEs6Q8ayzw9K2SNBaZDWwNxce9DYSO5YumRHu11SXjqt+Mnlgfm4XSKn/Si/8R
X+XTfvQFs8QZbgy70J/Lr0o+pI95LqeWbAvYbtR3cpv5dlYoIkLva8T9bT/qAKFV
VV9rNLb/kldjN2UVKfcUgrthdFslmQFzrVuzMhIrVmqpkV0ijlAYb1b6fvVo7iRO
TIY6fIysLoPtHB7QwXiTZ9tXPLKgxScyRNFhteWpEqTZdBPFiBKQltkhPimciKu8
pIEujTaHytjF/EVzIXreIJl6u6VsjpIa70wGL2THXHwaRqczWhl1pdGgtzISe3gy
jN6z+1ASh+V6vcLLdtXQoLqH+ywuW0mewoCXKzm6TaE7tHJzUp6liRMYKvtbS+SM
iPd9t3sj6FibiD1FBbIJJLpFm6K9Xop8p0WaZO6rFqC0lTEizyzrj8/6u10h3KyL
VTeOvcxvBhB67lEjqnP8boH00vNGHNG/pTYDQsLsHYFau38hZl6l3O6KlsM7J4JB
fDMofCbJIlDKAOBE9rx1sgdsl2rHCyQ2B20KJOLk7wL472xIyCd1jI1rCJLg0Co+
jwhpCpsZOxE5Fuaz9h0Q/1kCO7WOlc7GyvAB3lgkyH0Y0MxBQ0ullVerOz92GPK7
xZQ+BLTTzc09tjzirWetnZ10BtkS8VK9pyQR8bf/gMK/PEGTlN9jQpkCfBoigJGy
qNauPM7ji3KdLXP61C4m61c/cglSj/3vLQdi6DNwCXoH5NZT0OKMpbCvocljoUxC
Oy3QB4LmIzqLs5JNqcPhPAd1hdA4bnscAjJzy+vGGUjrUoxh0vsxSW0DbszFHG1O
gqfuX6gqsBlXM5zwYLOu6KuwGy7psd+1WEuBFXz1PY4h5VTNYC2ZTDyLeZZKj1p6
P4XWjDPoPf5oIO7AbDlskNyLStu9azknZyCTzk1rUBrSLD6tD4srorp9MKGouCIJ
waOX34hyHoIqjdxkYDZxu6KFBz+S7TSuF2wpeNlnkKK+dMyRhW74QTvGmjOblSvu
2s/omGa8Mk3bVVk+bk/SJFrX1/zg7leyb0yc6qMErFmxf5wrGqAgUqYj0dUxCiox
pvYGtDoQDLuoZlgY05STybxTQjsVeO/5lABrAq8UTFZqAvssQmBTFl6rnNwt3z09
sYxJfT5LRFkCWEoY+ib2e1q1GQq9DRiYjWy4BtyJ1LnuWnkVe1OZHnNmxuo+gg4k
ImBOjCzk0E/CkoSURehaQW5o8GBq7HbHJ8SBP4PiLTR3O/xHp7E6nF09iyPmT0sS
EYbsUBugxz4dONKyN3lVo6TfuO81etdJwsH1kNipnIptmljo4/Zd4y6YMQ68NpbF
dHQTV9ryv7FieuIhVaTpfOf0RacH14BDycQIXuvyxxYi18T86orQE2SagU4YekCg
dfu9ZlBww3A3aLVr24oSRrNz3sOm71MOL2848sxqY4Qy++VahlbCx/2BEpBl813b
Rw/X+6jd0nYZVTqbv2q0OJEwcUIK/khhwvN9W1QCkcMo+8/HwqKhmW9uDxfUcJ99
nhvQGpONl2/SlmoEOHqJykThbDGoa1JcVqmrhoI9t7YQ0sNu0rcnGgpJNO5dRx1J
L/f3AkOYtZG4+SeYqc88vdFoFuawx9u/jy9XZnQ/2SyD2aulXKxnL2JysOorH8VX
FkQ4HvQW1stMfY10lcFLJBe8AzaRl3PF5I5FpYkwjAkz3ad1d2ecmkNuEYtz6PlN
4oXQDJLvV2K1o0ZY/aA17fD0aftDAFSVsFml7X/50HdQas7t8kURVoCS/ZqQmGQB
IvrRgNhhiqoRPlUHvpyBkjEb+jq/iHbXyVse9c9RsyY7fteN6fN5ZyszU34K+IRP
vbAnmv6PLRG3RzzDQGlJKcBXsPjIF3Md7MY2lDNf3QrLteNjRqYLp1deVfwrUrKG
tmas8g0GHJi3bNkTIb2/ZG93C9y/7J362h02SPiolgCp+Qbg/uIwX3eh5Qaf/LLd
uQi4merllWl5n8vs+Ts+8AAXrl9OmKzfAMd9cQjrYRiaAnIRsNCk6UzNzYWFa5bM
EhUiZe3klOW+80J3A7MZNoVIbKgkUxMdes4lLsW02nNUcPtvsxy4sjkNRYZkutmG
IAQSgx508GJx3t9eUNtWytIuoBDuJf0OZjA4HPNopwxqKULYK6F/VGQGLcC6DkRo
+jdDWbVf6oyausqDd0zn52yFvUpzXsKfW6MqQ/hzZ6GDPKnKjhP3qjQ+WmMD9KAf
qgDgoe4kXWglktmmZ/iNaeS/LD2XdWjjXFSSdSYmTniGfL2ZeZBC883MXB4V0s+G
Xy0hhT0Mgxa/eH6wXwOhd9z22SLn8IxbccmUrGtlWDHuo5/hJAFdpj5/8R0xilb6
ue98N0WrmXYAW8BeOVW/TRX9yFSlzMqkQb+0HLqv3NORTn+2SVaVuSK/xjPZTtJz
ru5WCgJRO6QQ7RpffKGw2ab2RytrtRn8C8a3iOGiKhEI6g0L3qS9tkNX5MOtiXYB
6unH0AI42jjpMC4yv/2WQVGrkSlJivmqdv6EGK2+LyP56/s93MTUqo36AOTJSfJi
zrdgjnQ00QwjxW45U8LFHx21DkqX2kn5aFjj1+/m3cVGqjhguVb8L6f0iQ/Xfecj
R9Dl0y4HZJofAhAjHvxYwhdaFx83tEyvdh1py7UUUJppV31GIFXeVaKL00vVwSNg
2+tAK4Z1jBzZWcr3OydZ7HiYPrFnB5Fbfzpw3K2cb6JuLKJ+1u3rnykhtnLJHm+K
NBlBvFsSh5G2YxJzcuECuOpw2PmwOITI5y0Wmf9Rom6b5oPQJo5Xv0JtWrJSTWfO
ZqMHXyW3isR25DIgEoMcy7F4+t+ZPk9PODYM1OBQ/Mwhsw7cEonqVCr7MFJF0mmQ
FegrS2eU+3MS3HWYreXVmH92M6Xgy22kyov1WP8gbHJuynMDgoHYoaUHD5ZBxQ8i
RCSXL+AFC8IukfORkf5JtsyYJVPB4VI16PpNRahY0TZ/XcX0cVmwxIzTq8VXbob6
jxUTD4u9yZz6lBIXjxvnZm6p7Mo4uNt4ekZS3qgRhxOy1Wkmrqlv2dbjU4F4rntv
mXcd+T8M0WNLSLr+FCQC9x24DGB1YRIVMqeyMIVVQ68gkNzBZ07a4seAmP9yuCvH
UZv17MHTefmAujltN2pUK59vz8RwXTNuSIihpHntAEKH53e8bSVcJUwPwCRHoJlK
ETG22Kg/odE65mmO/NiXLjvWqW9RSLKGQ7ORDv1Fn4ADBJfhR4WbsHN4c21ISAVx
r6f9ZllcMacL4guSmElmZy1yH0kTxIEZzrplWoHWhEMSvDbxQYjboiW7gBYGoy4y
JSrkuLm0ao3xjWt0tf84LZG/Bz2AEzHhc40G70y1K8P9FF67Hwkk7GDNJzDGG+5p
aEpYcdnE+VJGszseP4FvEuAzsDAp8Icx9jDRk6x1gtN1HhQPj/FvmYpTh6QWTaTX
EV8Nm7sTeqg0/x9c+Q87ZM/9pLyQzFTSsp4u13c3SU2ET4eBYVdoNFniHZXQk4LH
6fi7y+uLpAVYdPlPZP5+Yjglk4aDHr3s8HVFgoSusoHGObUMUO8u1+MRkyoCU82b
Jrm/E9JkZmm4UjCdRrPPiVJGEOyIQTJucjm2vqM5PgrlLXvqCHW3f15ydc4DAuwJ
mU0bS+vLjK1N5ryQ0hsGTNcWc43zcTIZ3MFLQZQ2ANS3lILbarnCefZK5k8FUrUP
7cN3NkeXNK4mrQsdSzzSmS/O8yNEvv2y4iaYzRDzK4mwTcgAEdRbOz+y8sXc1mJg
FVJ46M5zWcqZgHiAl3rL5b9F0BLvfBH0nP1c6FvqPPkBByEQL7n82ZXe5FiX/UEV
eYUqP02Bi9p2qGlTFR2S4w7ArpRuY/+29YnySPdfcNStJ61zL8nqoR6+HAqF5A93
kiYsYg50JjTB/D722NBp6LPdQxzNdG6i6W6XYlrG5uxx0PMqbvmi5vajPRevlPeh
0jnyuPv18UOPNkfq27Tt0taiHfyeUfRfgtNNqu8NWteD7LEVTTZVZ9SMHkLhMHGD
xWGExU2KUupXkTB6E/eiOQkrqbtHyjrzMrP6D/NxJ/Hc/eljjI/PKkTMVNqoBdMp
NXK/7Jrfqb8LTzW9U5jZcJQinDaheMMbJWs037FDPO4CXKTpY5XUhJtDDYYYXOEB
hJ3z9/SqRbHM4zNva+Q8EPzx5lhONlEdiFD/+X+5z2rY3b7y0c4tY8Uurug2ZGVn
63n5CbssQOxHQsGjYKmFa7UbvAHsxYtI8FVzxAe2+gwkS2JE7u7+eaa30s+oHM2d
doIS2Ty5tDBnQdMNwqTTWtYo1zZqpd0t8YEj9Y3A3LQr2RpjFc1bcu06r04insMj
iTGIt2QP8qIFb9dMq5TSVKCf8ByuI99QzmHjwgU8uwi2ksuluVRB74nA/AtwXz9H
RmVM996y+/DvoSWpvCNnX4/S0NDmeySwBmbhJaggHAYfv1k14UxXCRy1EzJ4jMx3
7GNhJObFR4jLiJ7MioxC81QVHBGnsxB2OGM5NKMK4aqVncP3D7fpMZxqTAR+nBwF
G+kBTLlWDtBlsSynbwJSuAAPUIwJOVHRT+6P9HEHoTm9zSwML71GbQKCum/pN8gW
OXfiT89kGX8UFpz8Wtsr7Lptmqc9mzUScs3E5ydDGBxnoGL8RSqNTsPIi9TTF4AX
ojy9Trwl1tjlEDgSa5vv9azvIi4KHeijOhgWR8rdg1uRhK/i0hFFxVXcY9RWLDzl
yW1WebRsa8sEeGF2l72fUyO11k3Im+ioHJJA0AN/Yq87vQ0qWgVO75d3YYn9XeWx
J/7dfkAwnlGKbJ5BzoUQMUA50eyubnrGPtQpgAnJkvBYCbcvuIEU7EvaofkIqNDd
i2GcFgBOSYxOD9zPsNCt9eCzcDlDYOgYq+ctCWv/h+Nt3ExLMDXV1Fm04sFuuWzS
NEtD1HC3At7YHyPNPTbtBQEqxdCRZ2U2S691KcSrl21BlMoPc4Ew2RXVQv3K3qA9
pp3DAlfspZbcucUNaTh91XPTXQD9JL7NYBH821Uq5PhYJXWqC2R2jubUYnWq7C6/
bqSz9banHAWhtC8Yt3KQsIYnyjOoZW+FZHFx+Tghpf291b0x0hulnUwnKIsyaMJU
RM6Okw6y1B6SxSu4NgQ+T1MufyCssSnGy6mMcqg4AKbtBeigC30jQpBmFDoOVLmH
W2TYG7i8gI+eq+IrfhLjz3S1zy28urT+e4+iQ8qgliFkof5rGNE26nqAqZQ8PQdn
3iDvIk/vkp8B6viu8vPiG/lEAre+7tffdEOAD01Pmj00EZfe7KEmO9lfU86vCWBc
78kQKsJ5awVnhSWYpdF8MdF9uC7t8wSH7pS+d6HyXv3nXDdc+kDx+ZVRdZ2Qrdry
a4UOR8aNAqgpgVnOjWnwxbB/3ZVjcmd57DUuF4amn6oPAnJ7LY2UXOOIsRf3w8Qn
4zne7IGHtENQ/1VFDog49Gtmds8OamD6le25Shac6YlfwWlCPCyeaqEhUkMdLdAm
+E6Tp8YfLtweCTczOooyRIdjB+O9GQOaq/6SS/Uva2tz30Switi2UjtOOwPGPj75
XGBm4hE1w2dfRls9sgEfJZNtu2s2LbbD1N6G6wNgQYBDRXcCGMF/QgqZ51u93+Tp
5aXQo2DiH2/Ek5WLv/RVI/n9QdMo2kKdIuCNSEoyDv5SWVi1UtoS/Edccrqn8MZS
NOgnsz1qp+Axd8GmtqAJ5MjC4SONy5oTyuxLFOAzcEE0Z5Z7oo3DeUFJ6p3OKwn0
9gMQ0izEzfCFWVpsN+yKyXi5zeLHdzORw09VGAzbkqTS5ixq2M78IyiIfAQKYHR5
Zba6nSuAR7RTstLVRwputMEq/7dlS11ObAvC/ywzD0wBS48R3MKrcbopslTLXJAg
JNVya7A+btqqD4q9/Pl2yAEQ3kD08rKvwJrl5bxfO41OU513kZWjGsVMaEvNmlId
qcUzn4i44OtqsKfoKTHjTlR+jZ4Ux9XIxdoYXNzERglkkENolpNKkcoL2+PQE82V
e1nXRK2O9iTrK2OYbdqwpynJto34E1EkH2lPRDmfrVUchyD3efNnoweAbNnkJD5g
i7Mzgkm228T99Ro8FTXpgpUuGqXxpKZyDVJzsUftSY1USfkT9u6SlFnqiJXBTQLr
x7XGytc8C/gSfPxEMc2rq+81yyWtXH5B+N1jV9JNJ9wN+6OkkfRtPHDlOsF6/9cf
Z9VgAZrU+pg/zt5/9ycAeTE35wKVrxw4CewlK0UI67x/a+1rvo5BG+QHzjhiZ6b5
A4R8TThxwBx/jhd0uro1DfUiDMBN6iSLE1i3NzICQx9aXAvbNLAZupPkk0X1nrSd
lcXf6PDdhrXUV0xS80ofcDl+DKdvIsO396scgJEVhLELGijUr+RM9Maa2cC3qTfb
ZuR8lQnbTeecFvhF/zSlQjMAZATt3YExgQd87J05xi8f81n3tGvD1gwT/BIAbw4f
tEPpDP423K2QNczJ4F9xGqvEQl7p6IaiknpRqbTFcVXO5lC5H83oItvI3rGJcZAt
7TbuXMMEU1+mr3ljDn5N3RMAjVMHYKEhwN/Yh3+rn+xCk8/jBSytZz7x1lxhvbV6
QxnjpfM6UkjKl3FoXqYnknYB9GP+Q+0I24LUXW1WM5aEDegC540GqZJWiK8+KJAv
S4K0udbir1T88VYLIBDW9G1D9xeSzCbtwbvSKkZXt2V/Lnbh/pHf5T/9ut8AI2eB
BiYe+5kxvDICF0PP9uEEzCGscqA2Wwu02hMz76bAhnysq+QOf2O2lVaZ7yRfI3mh
T9lcI2JiZByfkhVWhMnwdHCHZJOZC9Bmuv7mdf9UZEChTiaZYUAcovkXUhl0q6iN
ipYT9gnMIQvlNRMSVi8312seylN7Js7cz9LRixALtNcTFRJUbCG4a8q61NBawH+p
AG73D5IgwzYwRLj/75qFGzn5g7uM6dGUw94aWOtWV3AT1tmRWUkjriIoBfZCilsI
hD6hFJtUDcJi/CeXGqb0AFkTDMl/ryTN/ooxbWtWLgieLyCWeqe0j3KY8tEbk25x
kWjJjA47DtDvQfTUV1ee17H1v6qbpq2JWqILgGyHdsmftgk7sRz+h0Ah/wCcM35d
J6xFLh7PaAZXAZpJPebXz1PcdjBRAWT5cccCXyvPiPwE7N+cB/ed0KFUk4EVJ6P3
l9FyhLOIvqEeAwhzJ9Xd8PklfbihPEJ4gawxC5qYL3bpuj2yKdsGoTP9ayLNww6X
unERjEfjPEM96UrJGXajw6bLSz2r1MT4pKV2yXUfe+ADyWNRh/Os4v+gUPmzuJ1X
OkO/a9FfZteRVNhqW+Fo7DrjaZhIdc6HKzRrkP2CcWmYc7X2sMEqsMNKerzAyZvc
XDwI5JU71MPTy3LB/PJ+K4bOQqJ3Mq+2MPdRidmGcqn+6/1ajvIF9lsc1u7SHuAQ
5IRuBODdsLSKP3x6cY7Acnyy1UeNgxxskd+HZ37zWDAeD7HrGlenFCiveEInVT4a
EOOHsED3a9tmInh8p3UMzBYm5AA1hYp3S+gVJGl38+i48XPwbSboCpeGAmPpX+bg
Qe0IH5Dpd61Tv5NCFD7MuSLEzb8wdyGgd7efkIHJl2ko3kL7MaYfzMlNGI5KBxXW
jsZhV/Ul21PgMKhTHWJHVU+y44MMkKWWou7Tft3ak8VMsI7yhKfPK1kkX+GSx5II
6DkvFYK2NjGJQzuZN8fug96FoikeDQifITqoXPd+OAGg0hPHemKrrIWo9WdLU5HM
ViBjWiRRW34t9oa/HpZ+W/aLRbjcXoyLA9IzQp/sRw5VZoZSVCDmG+MKrEoOX8Lb
Gsuffryu9tReM7I2/PHR9HB6xtjXweLzS21Zm07hpW6ur5zXULICgdInEzS4PxWT
mqNTibz/yN/2SOqcUS6wecqm1hcoEy3p1kHZrQkdxWnlbX1EN7Pkw6iGlEXQmrBP
ReXBbdAmFgrywW+L5LsP4ISD++mwe5MoU8Hnbgxalat3kVuuwC3jteavo3oPmwp5
irU4fgUYQeg6brOtamtGKgVOI+Vyf03+0Pp4KMKT5Zlcl0vCdhKVW9n7EkqlB+Tc
2w7y4kyPCVzhgXB7F9ptHxWKk1g56oBjY07+Woc31DcKTqJxBqPHIZIwzxlCLU+J
hUZ8N3rzdKLy8rUrOxvyqtzsFQQFpdLzJ2TcvdZ+uftLQKXl5HJjO0EZ69FysYHu
DL85SE9f1B2cW8kwFft1n2bz3yPB7/2YLTOoZbiCUH8m9+c9sGO5+mKuD0DYaP/r
CyhKP7t1Vdk6UUwavcAQMimJkhYhgyl6/2LJR7WvDl9ZkkiL3lWYrJMyzhIcu3YQ
8n8V3+ReTKHZ2ecDiGmAsorDpyIZnZOKSCCEyfO2tfgEiY1akDvXm4fVo8PEeYXn
KzOlt9GpuVF4ce6HsgiGvZMd/W08uXY2v16o06agTKik8V5EzxJZPWddcjrJPZSO
HqN/mQtsMWWc9+dsVa1PfF5zWmgCLSBLALKeJtNHWMr8vN3lxY/1iwYQuXOyJXSP
RtDXa+Bc4iBoC4y15nZ95Ngzb8DBkANvwedMS1iY9CInCG1a5lP43jGTqvEm7DJI
pYjlM9G6w0KPnc7Fh8rI5TjelB8dVENRFP9VDgM5wwr3i0UXIoQ0xM9lCeMT6BG5
SL/PX9hupVWWpzXz108MwGAfBARTbyQTPUHaLZpM1wplP4Uje7niVMEWuAyhk+Fo
3w9DdRGbfmkLnOMF8QzEzWBhbTKIkdeGXtCHC9LMbiF9Gu7wysxkr1a2Sv1Qz65A
qTAv9DrzBZ5UaVChXDucsu5aGPMRwfuO2wSJgU9NjuojWlSAU70jaXOMxR8k/S7b
P4lrTI09YJ1aurEc9CCUhOTe3uohAk1ZbztkoxSNIp8vaPbCG40qsfwgMO7+4vOo
R6O29/DSul5U9bWyM1s2LuM/RB6PfVaCmWw7Dx1FYzDb0QjNo53DLAzzkTL+nCOc
rMXL7O47Vc0MwUmrNu9gY+7xqWzdlarEFZATW1NSjd/86QLJXeuvyi310a53Pr8u
ocW2HywXI5HjCYtVZsslsj5ItKhjFi2wl9tsDULevgJbw1XkSzle25tJkDY8wjiC
34Hd+cXe21YP1ItXqMznSxYbkMQN8UDLJNTPeLFZq+Tu1n6NscAscsWs1EqVlFP5
pFeXJuM+f4TKBGp4ufZntxO6XYfx35VEyrHct0MYwvkE2KIugoFMOsanP3njqYKc
8w7PI2lKMwkWMRG8qbqBojTtSWfXu5dqF8eBUxoDHPiB2ecaVQ0SR1szcMVEaJVz
2ToTNIeA5CSskRiGUhWAAnaGf3UqM2/j7w7PCl0rWILIBFMgFo+CWATSu6KFJ2SD
+kwnRZ7BD6wExQ3mMmQ0ElfcgQ++MUWLWaPjM5mqTLKxDDp/DGD0izIt12VcqJ2l
hnkk4IRqb5VWfm7X2CfD9PAx2/zfh/1yNBSQOFX549JrI0cq2W/NBs2y8JO9I4F4
TUqX88f3/f29TgtyQ0aHD+OyVqg7TTcHY427iGFtaaCEl8o7I7LgC2l+WcX107ul
nwQVZ1WpzTEVlpeRTzp24cqyxcj9Q5z3V7sEzFeRJKUpWHUOZ8N8wB1m56otXsZy
VmqCt4qWuVcY2k/IpvNjIHW0xZtMyOlV1WYGZhOtMHh4P9LxtNps9Dy494WUcGlW
Q7rC9zqcl6jW7ZjgQhsxmJjiq9fXo9lxkRGqWstRcu+Di8fnwBfMmI4e3PlOj5TR
CpqGjbonXGIEVqEKCdeu14r3Q6mHTTtJQ57DK2m9k8hXPLRvcJXGc3Gem9enLxdQ
iVaZncEmkCI1QxTJ8SBQtOWh7hsq/36sutiVP4CQQnp27NVhHI7yqHosw+d1m9lw
xQebEdAeZZIVf2JTDmkva5ZitL8F8lgBLQsD67qFCqj4vh6fsBAm7gme0GNbsMqd
laKG3aKBv80YvkyN0BP6HMGVNXydPBC6dCCqP79p6wYx5DkSjUXpCUerjKYY0oFH
2Kk2Q5z0VUQSWlNrqNLQzXBSqZBeVdaBJC3dNfXlk7IEhxFQccQnM7Sm83jdo62t
37n5IKWGE3fmObxHbwuzpNQboU0E/DlR0ziTZSDS83aUx86vZzjAcZZdDelSg/gd
Osqn4FHgUx2fIGLUpFCSq2VBBqeraNUHsQbLN2taS16maKfCWSlfLWT+/CboKUnm
X5RQdXqgNsVYyDXpU9yGG2QsOZIQbvy8Tu/pNZK4HnS6hs4Ro+MGIM4c/YUu8Oau
HmsbAw21X+2Bwy6UcRWtAZKpc+eXkEbhWssg9GSc9iPnWaDo8SZgh9hZRckbFPsF
LPCnL/UhVOWXjshZmSjAL2Rv3DrVoghcKm2LS/NqFATcq2J4AQNRJ6XlW6k1ogG9
sAoEQyfABWfWR4eXkKHEKU+BTLF0+RimVmzjSyRmjM9Ho1ArlTeDBDXkK6I6QquB
smSiNEsG5dGIIbzdmKDw+MLef/9Qj6MQgdjHe6ob5AZmLYaoMHSYIFnskJQ62HFo
57qC5JzjUrtP2hHVaNF2Yc9V4utejYR/KyxS9MacFYutOXr9bbqKDD1PSYbUaE68
/tr2mxYOOohWhsAISxEF+SpcKG09U1U7+l+eS5VRsPu2SntuS0U5Ho2WBujp5H7K
X2ubtvviEUkeHOJ8pShNmoc3qo1qOKxh00SmJFaWeOrXQ8+Y+lLasfrKYvaZI3Il
6+fI0xaRPxlaZRFBmX6bIJzCsHV4vptOi1ccjN6mpN4jaUKEZBXp6d9TAnJ0EMPl
ozrLScPXYbZDbvrhDT6gUEH7/r08YCJDuzUlcbbgZA4Gu/A5q+2GjggEZxqwZFkJ
v90v7DhO9dhpWkPXoczlO9A+wjCxeWX06jFn9nGdN8TwaLnOhqs1X4LKm+gAjShs
53JhNQic7vVB3yew60pCc3Atv5zIhQqeIACiwBUm5auv3jJ5brB8HygLa5j0JSh6
9yrA4kmXTDo8LegTIAjjDf6/TeA+nxvieLjjgHXB9aM5Kl27tvQYhpPt9p5CSklX
5URcp1WBF0qasdeKiDLjNTZIDvAPIur6WV/6vIyGG+01++5mrSreTn0MT1EXlFeG
hLNzM1DnpOY2IdEUnLMoUKJahR7U2hT9HFARs40A0qQiJTAbxXIg6H/FN7h/bFUK
F4mXZvLmieJsThOuzev8UTcE73Rg4GasMqHpc5Ro4uu4GfL0EeiULB+F4YOC27eB
NFLGR70DJpDfHXOY6z/UuXomLH7w3UhYXQUYdWL198jigYUp1NzJRwx+Tpxkpz5z
8+dvu8agEYkf46FEe62FHObMmwV1l+jD4zeAQkB5Oeuz6DY64XmxmvgICgmrWm4E
F2scmKooLwviVaS3mX6TUrJypr9hzQvYY6zyw8w1f1i/82C6tKhrBbvBMxc+GaVc
XpcenkWaVkZIYovz+nSj9w3M4hjTgOclq3sYmCqlKzIvGPGkMS6/EYfyxQPGEnFe
JDg/hnnxpKM1PqZsstO2VU6ek1L9aBK5JtlWFbUmCsWd072Fp1qhaQvKdCJBBZWt
g+2Uln/jLmUZvOBczQSuTkriko5yclxww72WPMUUJzy5reGoQvHWeY4ri/EgtROx
Wl+1EOqoI9GexWoTE2JH1N3YgyHATCNtwfjGPkPdNd+NcDcfq1kgrKUkX4qpKAiL
THodaf+LeBX109pgRPGqkDP2Ov67ex3Qu06Fuqkfooq6OOY2DdCJd4oFGXUf+1ih
wMvVg3iSTQpYXtz7T8DYTMEygxnHjTXrQS6TJTsA4cfNMgggtEuq2MLPbl040uCa
0enNfEwhPQQZsnanUgszXWv9aXGCKut6XNDiiPsCJ05yZLzpwLIcH1ok947YRfgR
WVFT6LAlgAH7SbQuY8nmi3gG94JE8MEZW7UanSbz2cXDdIjMPvonTxiipEXaTCxJ
CtNCUSGXGRPpfSL95ahkNGZ4oSWn3RLsOnCL4ZvPm+esifIgTP+ZEsuvgPuenXhG
XqvOwAjRl7VSgjJaVcLNolv94Kk9q/FQ4xyetT1zPOHkERxnLVN2+q9NiR4sz3Bn
2oImFvy/kH3RTu58geuHvsHVPnfuMR672k+CZ29PF6kw7eFesf1oVETqXKzP+Z7x
+4uO/AZtskT4jN9TAegCcSOg+94g3xn+RtZBtAF5vCw9JBHg+NoSDkGITdribIPH
/7WZibn1UuRtdROL97UqgzCQn/LKDx/uupSe22EHPqU9B6PGA49FWxGb1CrU1wg0
t9pDUx6cmdf9+xD9IBqeNnOXkRjRMKunTlxysBqOxCSTcbnc0oSURqv4ZfvDXP7e
dqKFTVcNT/3gJM1DC3NBDHk7iGPGlKnMAOnnWn51y4LHCGKUzzcil+J+/x3SEYqR
vb1YCnJkEXtsAnIOY0XhfYqBVG4nG7oTghs6+K4uvu7AMEsG7j9t1WZLlwvgARgU
S4ReguzZF47+3EcfcibX5/yZ9DRqMlL5glgJwTL8hrL90zyVVq8kYuJzzkui82Md
Ig+1VW9od+hcmVCs3UyXxmHHfnuyN/Jy9tJlUB8Vt9OEHrGABOhiZnoP68RGmFMm
l0/ceqODsMq8QR8MNC4wJWswADPYavrmlEUgiQkzKuuoF0CnnalR4KI1XTY1xcSR
6dzpHfsHQboQ/b0+SPhpaq/Pftzvaqg6ZPHvQTc92lMVKu6BVqHBqbmbg918y+x+
E4+EDKvcJjs+6gnGEnu1ZtIjW25YRj/Rs5oKcORdVoiSVps+P8HkjNIGyZt5w5Hf
a8lxO3hnEEAAIlary4PQlcG9eTMuW1utQcktdxc4V9TEiPdCn+485iz90R2xAaJR
ifCIJHmV6z7iGKEs90OxId3aqLtbrOag3AN34IlVUQm/PMmYBBVRyfmdu6wYwmjy
SU6bvDavoaTOSjQbgrt8yUGrtguHC/m9MBE4gK1tnsDbFU9WmMOT15GasqTWsK4C
IDSZW0TbVcIBgvjY1w8yyOf9RPIH+kFy18/zlmYn1r0obnl6jpuP7ex1XRJKnPch
3IHyJvCnU6w2BLA0x5YvVqfM28VvU9Rb3mBy1uP4XDFyqQn90quWfYuLASRlthpZ
1iStmu6Xl6sFbeYs5Bzjj+xSYhsH763l7C5WogH0gDtAuOTVjQNRJCsSJGQLO9kE
Sc9xe7OY0xigtdiu3+MragJMitA9zyvBDUZsoxZrOdbxDWd9cHF/Stpmuh6r10Yi
6P49iYBua+j2pQBaM1Su3sbZKam8CaG2HXth/kVobW3WglixVHe/xRoApqyJqtAG
4n4h1MzSXOg6XLPWRh94YepGYz7yialFr9DRP+6733UDek7m3rZqgswQANj3gsWf
3E6nVE+PjN3m2E/LtYJYaulDJS8IQP8oSuWdQNflkiWq0RAiWaXP3az+RNvrep2E
c6LJnF2ihCOKZb46oAkxQCF8nyN+mF7ukYFIFlXbNwNwJT9+q1miwn32MTWRhN+2
262fNDqqtvNzAh1k6kukberlMH8kFPdqynZfC0GAPmGK7p3oz+03Vgio/HBCeIN1
8P18xLml7SaLe6Raq+Ra+h/WEOjdJ6XM7kMJ+I8DSWNw78JknvpMOdvpHqrpa7b5
X+hsde6tloqTmzJJKaMoWi2wOE38rn6e4QDQk/ohG8vB5AQNKBacRJ1jry+nFID/
7dWEQuxDHjKnqwjZS7N+QV+pM1MDp3b8jv/zJp5pZPKG4LiZQehGVeDA2N2syWla
wJLgerIFVvTxMNIzKQi8+ZVYCdg875KnuNMaYKlrX/cRGkXyv+Xr5Kbac87k+Pz9
pnJr2oz1y17pBS3LxnpxMZjvs8Tm2u+GNngx8dzPjBRA02RIZUDf6b8VJLS3ba7n
lRQBmPHNkz3gkzpjsHCgwyf5lFwCEp9z5L3JPc7cmI/wSwqWwviKPNF9o+/i6fzB
5EGc+iuEOs0cSNcEXtc+nLjNl4mPtuvUObN6BiYWeTR5B8SrPGKCuX7tq9O7m2jb
jS6uG8rplX6BmJZs4WEtf1L816jeGBx1y8b/cHhjAbel44YTb2WCTw6UPzQhBT6u
PPoPNyzZQZRM018loxM+XfpnK6qETZGMk9ct/v9BjJ45k96SsHnVxUttYcSXkiZs
PHi3glyUWI5R2Hntx6wTe89mL5KDt62QmOag9HGwkFV+4dMiHGJd0Gjc/Gt1lMpE
gNyCsg+CCbVckdjQD/OaZOSxgInx8LOIyffLbWghkLleH1cxIoG1ZfvFC2dihJOr
0G9EeuHMmFH2zPbB17xxln21b4YPTTxNHDzqldFBSuQ7InMIpFArSRobr9GkBNCU
Z6YhkCWiAEJSz5qMGA7pqmJuY8fhBHqOkXjineWYcO3SKITyHmNRcNOXlLbcr5p5
Kj456HtwfQN+J1wY6Ua3G/Yql09ipItGAR4O2xwe6AVKlMoR2T/1quDXhibt3/UT
4O+qZ3XZxFlx+31smzf/a8PTvf2pFrggYXi9tzsX1Rz+fOxbwo1TaYfGAENJ27ef
0dmQxLQbpbHRjf2fDN07FKvSU6wqJ9I9ndPQTvgH7G6hIt/14fSEp3K8LrYTRZYQ
0xoJA6n72LkQY/eowmlwe5E1YZaO5vu8zTLUyE+xja89A09+L+6w6V4tQy/cOV3X
DVLB2igKkn8XWgLkyz8OLMWucbDcAbnMM4gGBN41WLM8LC89tKQiwl3Ned3BonPz
ay1FHz4ufMb7QNsE7Vez+163M5iB8QEsXbaT8YZOQhiuyXFtOqoZhP+AlK5LBF3J
GSmDyZOY+sJqrPsAhq09iKB1blPV02kNVf6feu499BpkIviOhDVoaWUjGq/uQ1zh
R023G7tV4AQKBTS/3EQIyLBa3u0rjhBJgCUKw+R73r+7cpDJbKgQuZjdiYJXRdas
v074ttfn1vQGYooh0O0vKefXp23m/dmrUfuO33M4K9K70DE4Z0MZma/ugbkmrZ4/
tFeMx5k+02M+Re1B6H9sh69IJTG+Suyyc7Hpc4l3uxnOTGE0QNcPC+5mlwFxahPI
oBvuMGAvq4nNhB5yk0fSAXUysTB89b41PFHVymuUy34LVT1PhOLsBa/kD2HT8yDx
MKpSv4c2NPCrPmClHCyzIcfAhzFXzVGfMn6hhQnGOde6u8x0Dro5edhGFKZ6r9YS
vvtow3qb68l+8060en7mnXmIa5cR5tjTv/8MQTgW3fYSpc9gOEd4BfIfQ7+kQHHF
yEPk/njEMdlkfIICotl5bA832/1htFpvOH35pvMEr+pHDlXSXhT1zPNc4epWXInz
ThrxAE02ZmZ6pE+ufd6e+3UiG6q0ol/5X1pjUiqZUa1QgYI0FaJJvGcoILStGUN2
7+yS7sx2rAZwokT8NERvSq+LgbtcL1bXlC/Z3C4EuyMFalJdiCDj6As9xRut7zK6
DV7ClhJaS+kAKlICEq+60ox0DNp18l+6aUwsD6OaZ9QD/yxrabvikUtm9vwjd3nI
K3ZQ8/5jQ6uaeWhDXnFGGdLWJwDz3QNR9GAaXnawqqifWG+QydijU96zQHcL/77L
F3aIrGfpiGTWOkoUIRVLc70ZTiapEV2agNqVFPLF6i8b2XNs7cqM4FMYwtFUvhWr
9gUg330QHCFfcHzHOG7T1qOYdPJS3w7YZ79O0+qVSw99L7h7mkABzlwMTw9xMYSp
xhYNddOF1YlgOL0KUeM4fW2mOvTvAvaQOiDI8kffGQqC4qMEiuY+/lqhy0YVtL3/
iAlPmH4Gc2qNU6fhNISLU4/666OHaqYVyyixxazJQcR2hTX89UwZ9rsAwpQpLOmB
13mTBnMJUyz5vKdGpr59n6S41HQHh50709Lg2QevNz4Nk1OOELbDw6D4iKtS+DPB
O+K4V7Mm2iIdDZ5AZJ5DkcZH8fj1/CHld/n8Xl11wftTRMprfqgp+xw4beHJtvJ4
5w/EBKR8elh67YMwv2IAs0KcdOCZ6GbzTqNCpXVKC7nRDri576WPP4qhYXuUN5Ng
YX9qtITtwPnbhidrUhYnIAmG95mROaiUynKI5f6Bh76eHzOQW1mZN5zuVsyDg8j2
zwagUq7DMLxMeYjR3NQhZaJeFnNYa+L/jkuVaSjJwoncXV8Of2Ufkb/bBAyliXqJ
GVb8zSRl4IltkVgcj8Kf42/v+DXYivoOBp/QOkfbj5hADSZkrjK2gA7sSNf3NIbR
CMbjixQTKubu8p22tjl++YSZndZplbGjFptfVV1/pve01LQyfTx9OHT5b21GBcde
HTtA/idUx851wFjQ2KIf3yk1gOUHhCq1Bh+fn9XOwSArs/vIYzpi3GJFIZmlBy74
FVUdH28hhaoYJEGkuNLsU4wpnbfgBF5M+kRdc2sKe0ytqqaDnXMWNROUROh6knjT
8fnYxGcWKb88HR+L/V7V9Cv7aCz/JvPoO2IPT63G8yCwaZK+62RxJ15ox8oCDm96
GZA530aZMkwm4RNCaQ79UzTRwxXqfFpE0fjwzZFIBomNBaZoz4mRFIFseBfyaT0S
wYLCOUp4gz3aj9XTs82xLEy7an7R5hNWbDZp4QN5MbznkW9IPuVqADowt32jxn30
XJG8w1DSIs3iYYGOJ4Mq6byk1ngtoGamPSuWnUdePZNUmiLFeu08lIp3CK94gFz1
Hd1QU5y1BZ7cSAPQVDIueudrpc76OSFzCX1zILrK5SA7y11Yqo42Kbp5wxl9xJjI
Usip2ab8fVT4gXDixDjgF5shsDkHuDpPGPhKFQMExi5iCJ15pnptEC2gyGztw3Q1
XqLcH0qsEQKyJBtfdlFUyfS+WTJ4/W6aCg0fCu1/oC7hWNQyY/xdIL3u4kRdjMg2
IvS0g7gpYphuBXGlVOYUApSCh+0hR2FHs+XdlJlDgR0Sqkkc9SzQMyHES8nW/DTl
iRH2MCwCzKfB1GNciftBHzyzDfdrn+YwE7y2tupEfkqcXycCAavkAG9hDxNH/GfN
DymK1J4Mbt48NUjqFe7YXW6aS6xV+S+FSMq5+7M6zz7xCtM5gWUxfukJNpw8Ohdv
q5qfdwBt0e0ILicvuNBLfm4exzTdd1S5d0f83PI2xhDwIvS9trVkpyWrZyZe4ebu
dn6W8kXsqktDqCYM4Y9qb4AmBEO8nS/Dz8+USSUq9ITLrjWGonkXy+gZlYgD1Afa
D+3KfFjMlVHW6CN8sZj/tZJIObWWfatvfTwbFD5cFGKgX3Wx58/1RQnGEOO/Az5u
9QN+UPKgJIHeuojtUndRrZ32aCD4odsvInSIhec5H7mfX7ngTLL676UbA8sLJYWl
wvunvAzOw9tKwl7Be+RfqJmMHvCpipaUrbLH+83oR+DOsGMpxzI6BSIhh5ZVkTda
rbHx7O72G+aDsq7nNQ7gghMFJ+FrIaYQb6YQS4k7dhjbKtw1fOHMaqab6vOwdz7c
qk6MJG8B5Arrrh1vyiK1mSa8LrbwXvY/SM1hXFI1pmdUdGKvXTasYu5PvgGIXeVb
3t7+GXIB5qNNTU/gDVzQcTG7a3Lu5F90KxBE9vRTyELNnVK+/m2Jog9hY0TW79Fh
nYZer/M8F/1OHah6i2lS14H37kTC4sQtHiuRcPLpY62S7H7x30maAweQSyujKRHP
awUTvyJISGOw+JBp/4YwzbSknpgbR9nVW4nkEwp5pOd+eRg9Kt4p4G0FzVoiecWv
L5MrWusEY9GaKVouN0tRVhyrkfSaTpukZ1bfLi5Zdlj5zR8Wkd5NtSikZ4dD+l+9
DjUIgyeNgFVdnqtj3b6u5MIQ6plJoPs6+S1M07ZVCXfaRcIYfDA/RQs+I1TWBF+D
J6RdWYHS3eivNPx2RM74QvwWUc5gpVR0N05cAWJefBbo4zO8f6sQzoqdBrU48I8K
evn6qRXJOo+pvA93rPc2sApSR2swIyEnvBONpVK3d3xlmQfe1fIz9hKYGb7vS5bQ
maw5+3LjLVn4xqrY69DJP2nkcBr1kxm4pGQBEe8M2q3pTqq64B/h2xAEFf1S9kJP
I6LKk9+KY6GG4aQoxvmRV2M4Lg5EL24j1cyzmeLxzB2yAWY7fhxtQeUPpMrr7kmL
GEWrHjxhqKyIF9g8G3fRkP8fQUX5PyeRDKeH72Iq/SitKiA7bpHZkfy7xaT8knTb
X+owZ5ujCl0V8NxRjcX/KrjGXjHhK6iAeRTQtx60gWG/yylhHUwT4+pCR0xVhPzl
kPL2INKIzhGMckFdASjPYdwFc7q4Mf3Rk8pmlG/9UFwYHzbGq3CWd3BWTHFoUgEO
XsmbC56lJqH9i3DDbL1lxxhnLYMECr+5nuIDEOHS1N38HYgixolK1Bod2h2mvpF/
Vfa6yLirBpozAhy6ccs2BeMUgNU4b6KJG9moe2O/F5Ih9RUEXDFf0G29hBKKY/t5
AeexTvhiuOn6CmGVh9s9odj63RER1NTrNB4YIOW9CaBvBD820rkOtBTsJaur3IRN
PoEYSLhKChsmiKT7mkVGAceRuvyOoShv2No0NZYihzrShCz4/hwpgnmScW4U8+3y
KFdF8mmHOEmeBZCg3vdkwPM77drrQN3wjxThDASPcz1n3lnSQiwT1N6Tu2UYeCS3
ASNO0SsMVzswzzFHZljFBjWJfRoxdmc+v1+9o7A33covJr1k6qTs+5V4xIr9FCx2
D04mbfhWCuz/ZvOVvrTuI1bn5mbXht7OfW4zPdY7P5cmf982MxXnDVlOVJRthOJc
wvpFaGLNFaLdDAxnS/jdbu9p1Iv6GGyvkdaLV74zxj1m2WrN52ORYUuvbepvqo/h
VmM1gb8lZ7PsRrTTRPzyyH7YPKaOeZMbwewG8nRKbXVKge/BywSPPUXLKWvuq3FR
`protect END_PROTECTED
