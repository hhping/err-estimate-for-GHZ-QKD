`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HX9o6OSH0B3KfBp1A9g16UcFWGGLDHkRK2FtnXNNssFjx4X3gumn4PVQFR/nBKG0
/5ZF216/adZs58eoRMKJVenCPmXaQKPh2oQP+0YEmP5GcxlwFhAFdVkhWPAA9qnF
Prdnta5V556kvI8uq7n1oKSfXmI1bbrCfueFxKIuTadE8XEbgBKeIOTpuh004QAm
K6s6gopIg31Djr4KlkCiRr7Hoey4cmwLeyi26LQdGfYNDLXQ2x/rR3HFAtlotbnA
XQX7gq9YyTdN4lqp3Rc5E4LN6tYMVpgEIsaob7NbfnuzFL8K3QH8IoL3ZmwEKuK8
DzpiwSecscajdt/07Lka8u7vTmP+aDhn6elwj8J7wGDUJe1BELFBrLDsQMNk0KYs
MbJtfTv6q9LQrXuSsXRLDFcPn3sKu5IeoUuFniDwsJ9eIUVdo3HrVxwAFJPfzurz
N6DAVkqXwir9ofI9Q9ZGTbltfIMOVvI+mUPVPVWuq699X1B4eIMO3V4oKptyOVV1
T0LMJl6uE+5MVwM1cyFA2y1hBpE7Rz9MFq8XkGyK1t6pVPUnbNb4vAdyHOji4Dpe
+IgTGXyBBg0geyoSpfkyFsCK8eAh6UNYkLjs4ZWkUnhic7IJVOAEbz7AQ4XlX6qA
ffF60eHBjDuJdRSe4SvJ4Rg3Z0jqoMQ9jznUs4SISC4Ept9lTxIXbwnBYMUMtNED
usp1ZjIGhQy3pFSMss5yqASG9aKbCexHpx2ABwbupSG09qDcDaTbgcwB/2L60XFY
ljipS9/8DnDX7os34OPMXCqSDq6Fnzkx5xJu2lCWgsRpiykiVC1grlDzjkCNgohh
VcZioRzj9EM6dn3NRDwKXA==
`protect END_PROTECTED
