`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mJzT8NIzNXJC/8+7s09fr2ugg79uSarDDHCdkUfo6qLzO2sS43aJRcev7leC/Eue
KUrpULp38cCeKE1sfs9Xw1BHJ3/xSNmdgg41djJgD3ukcuc1VGkeCg3skQcAHlUT
3a6IIHaJsAwJOqB3HgfBfScgIoPcy22NYjJsZstHQbKkbe7mPIdUD3UKTcRulsqE
tJ3h91w8E3QousNAlAlb8YV3Rc02vPhoDouABQ+ybmbHOkjmGyl98WLUt2g5sOOm
6mELTUuRbbGkjASgiCMzlGUfz/UEy9aoZ64GkfF/Ii4JOz2om7/aSFHaJw7UJ8aB
u6SaoJoe4TCMt0WmpeLQ9JCu6LdUwwKlVsVDZyVrmdnClRoLVUbIxWPR2rQmhQl7
8dy/5tAJ4Vu3orb7venVyjkyHVduOce6l3EQSB3jo4+CWBa3yxXq52Z0r61CFVQN
g42j+B2q11S8ZDTVfo3LZL54eMGThlVY/7EV+nASG86Qh2x86VTTLOPHP4aWhND/
zvNuMbIZEhVR/19Hui1nntGVYDZHPne8VfH3zr2c+i5AvfvECQDva5DnON9gkHEp
LaDiPvK1ZoOgJ54MWMaNd7s3FDJH3BxVTUm24YXAGGECMPCQxea1OBHzkCV5pAbw
8tMMX1xKOd3bt8xhZL8+GfqM9faq6q/tb50IKQqFyVtgQjXiMbZQfTmAvJWoC9s0
qYYaKXsis6v+ofFBxEeztyhKFkAwQvh4P1Oj3LT27T9bt6ym0ytkl/9DVaz8B641
JwxRrIJ9cr6GZbZXHejAIMp4xtAp7c5wAq1Rk/ixvYPhQLRVg8U4/25Q6i7xnUfx
QjS5ZkMG7crizap8KLAZYMMlVVuxjxXvFo85veEmpi2ZvYL+KHrB4YTdJLwREVka
u9zV3SUhM8M9yfkORTSB6WTNn/paIcw7t3WlFmXsP8M1/5P8GaczrEtjnErK4qKt
TN3nOf8SQtc602YaHUb1GZptTVFb+WtXIr5KUVvIejO2uSCWs+aMOIyhVX+wXg8h
OlwWFQbPfuYwenJ9lRjjkAfMiEel2Oc+LUP2znj9+LN03pvnd9DmTnEvGlL0ykQW
/PdA815QSFuM3SRGbIM6bsXFkiv2vwSZ+FNxUcAyixGiDWqM9gojOQ2zdy++vLJq
KOVTuab8C1UBza+WQXa3DJx0NCCXTlF9mhpKI9VDi+JM0SN1ucE1J8Fev/jnJL2K
G2jMuaf/hlZYxuG0OGb9h44+C6TvzDst7zS+MngpM92YDdkE8DCCYIEhVpdb8vH4
g4jg8QtnJqzKqioPFdmJh+k80gGXLQQYL00rE/uhM7RPOXL6Wonwhgu+NmR48gsC
ccHT081xGquo1nIc+5EPdcblSHNbTJqgjdjl+w0gvCfuZqfpSPJQ6rCX94uC+rDQ
q5t5ekGgefSqeEbHHluRe/qZiAScTMvdpps/GI3p7nZUCnvXpfcMv23Inhcjt1BG
M0hlgW3HvpRIetriMinuk3iElm8qXaDgx2zhfx94p+6m1FNvFMX/gmX8kqZMPF8n
srp7xvSGJjl/6dDB/9To8aZQQPwVpiQTGAKB+HwxZg2+rC0yjkP08QVgePEYybUn
w00CJh1iBMC/ygxJ65vCrUBqIQfFewyGYfLuZSI3lt4aP4BS0IfJWx22LZ0Vxl6R
2biRBjkgwYXk7bCBvGyTzXY69HYWzkCargwbZWqvr+2/Wa4iMqPTkKkSWxASTck5
8byL9XjT35BL0FL+DJ4gxsWVkuiYrE5ARCnv3a8uq62Pkc2BMG8B2lumvs/fqIrS
6GfU3mLalGi5oNO9wFd2otCaoXKQjbA4AFjLMusLbTRcYtOOXsgtrm0NXObIILOy
wsK6VDeT1fTuFh9qHTaVPuvsN2fbjU0NvuCJjK68bqGvwhmvA7LqlgeCK0LXn87N
GEMEgE378vNVGz4JCnimmNuYbbcYClafwX9fXTTJebgg4jsv0sX6G5lEdnKqW3lS
abeAkdSbICZDHRNZDILHSfUr+O6EuIkk3z6fmOX9swo5BpYwX63c+3fqJdRjWsSN
GeMsvA9tnJjbVJwgznxyVrCy9KVyB45rXOcDbDKMCg7GrMIWXQkta2ds5mTdXFHn
MBiTco7XFQ/bbLTNmb3pqvrWFuBVoE/QxuOIMNhiNbVSI9ZYEZohDOhBUjuV2Xa4
OfZ2eSc2Ds7eIYNPE1yCpENQWTeahHBVx0IXmRBiPNp1Cf05mIkGju2qiXrso8FN
b0EsYh/SJ6HOw5wC6qeMocEHkVxKWo3MYOFWWu5qCjYPhXxHTjK1TilP6ilbFoBe
rm2JiTHmkj60nYMfCowbB2oTFlbDRVInJH7ue+M3p5Lo3XDWda9jF2AJ86krWHUD
VRBGF/dUMnoXTPdnKaIy0TYCthabKGrzzd1SyQikmsVmNYZUOU3Uw5pciRmhhnaK
Rz9dn2qIMlWZIpGFyiuePhhwW+VqFJa1bT+X6a8TeiEldN9zi+Xc6DeP9roJNYvH
DIdHur8wbuRp3EroqyA/14yxgzNMlp0AuhI6G9f0hGsmCW/iS9bvStCcTNfoe7zC
mH78nstu9TL7IjpSKf8TZopIiPiJoieXCNd7JYvYku11Ji+x86mWq2FLz1rHfy2t
97osNB/aNKbR2tv8/NFjRcAdtN/1knNNbOal/Y5aZgVE6jGqIXiYC6IMD4hMwwqm
C0DE0AHI5syHTwyM4NYiiY8RXxR+47G62HcJozhjWNqs71ZoZio4aG8s3kNDcpEW
jKBSWpVaW9iR8YOMviVSq/qzlERwvyBxLvpTzdYIotRdXvtir9HXice7JeilzaNy
bBpnOwdBqHjHmVmQ+8l6y5ryR4yMV+s/tDbGDIji/R1BHxid6Wdq2KLBnCCvI1Jf
kCZLfxUzIyvV/MC58/PIPRhSyhoKXghXTz/sMXYPFdDK3Er5NG/593+9zzTiMcD8
XkPo4YUT+zUQMJsBmEB0RFhEtwsBsRRV5NSF0/1e1w2FnKe7KtpH680SzGPr/3AR
BW3UZ7auJlMZ7JMrDsCH5jIJeK4AKul9b3Ywc78QsBja3VQ5cFIHaMN41Xu2I2o0
LKAhGveKlT6lBcUUenVWJ/C6NzsUOCvpexMe61c79cnApMVtRLgTxl6inq8SXCmR
H+8XYpnlaPtVX2aS+q6pMvTeiyZVVdpR/KQyi3gBlgWk599459iBgJYGhLdZ2qjA
gMrOQQ/i3pV0iLHH8rBozoSzet2wxN1kmck1pX/e6hQUNgHtEMHLwQaehWx6NklI
kd3EJlmtJGLxP4/IZKgjB74zpdE7xFb282GQnA1p3p/nhsH2boWKBlntA80s04+R
l+SapQFNz+77Z+sXjUtSUh2yQ3PjnTMPL9ThfkBuwysZWox97ZBmU+nHDVIZqjeQ
y5LOgf0GkOVbHUtJZnKBnPRyxcNFHQQr2or5CObT3I6L+t6c8d5LxGJD3PCfb3Mt
qXUKgZsLTpM77z+tWZe8qCaJfd2RhEta8x/PoSrsL2vbbwKd33CgDm/A/jD/XNCW
d0DdmkDtaWZvQR/9Z3JJRNdiahUJuw/MBn28w2jbH9X0AZB7NsPKkFIoFOyLM9W3
uc2qSJEF7yiLfQR1RKyQHB4Cx4KWRG5J7EBW4jbqahvx7SiE4JoF7dgdUpvG8V/v
a6PClAsTmKxLZTwXhVOw5q4aEw5V7d0nC7V0gHd78a1yNScUEMDJuDgJv9DltcE8
iywozzKbU5LfT8ecVZOgOJpDo4OOCpSJ01ROkbXQjqYCRwLSa0tk5T3pBvdTcCf2
7zGQmdoA+bKe7IUS7R6v7FVrv6V546wz2mav6/F4UsPuCx4DLSP/JCnTLVshLFsu
K0kuVpnVNyauEeqqWglXjMkTcEsD/sag/Ie2EKpUguHVQISVklcy44l7g44GdGiZ
f/UXwMIXyVxj597LhuhV5TR0gxUswuyIHtanzNetLtlDMwBytBDD5IPElqYf4gBJ
fQmlnQjedrBzdB52QVKe5kwoBG5V2mabOrtkPUodvmVXw2qsBCM6sPIFWWxS7qw9
zsgmFS0/hZeuakHclFTSm76noA1mBoNfjcxuJ/1kHtKTVYXn0yPS8fVV03oPgqaA
dXcWrbDgDiJD3IBeUne5LYcvBw6qWCRznfeoRRTQZtkggtnnxX7y0Y0fh2P1DSO3
49p+URqYgj5RVGnDuanoiHeJifsWsGNm8aVQyeqHG750bQHcD9venluiBQVqHloe
1jQYkyhajPArkOYjNEExakPm97J2ctdiOGG8jH8ATxajeOB4yyLygf5afrN+xXkO
hTwzTf1qc4N6YbjwccTxmVGFCuj0FlEaGIAWn4WzEN6lGPI1vXS8xiy+cVxWy1mm
yM/n4kg/lJd7w1w7rJmTUim53MFGT2ooFaDqj/kUv2FABWypeWhsKRmcz3W2Uenu
y2yhWo8RPjLaWTN5YlDAL+hHwnBZap21FLAaHga6nVeqTEE3cqYb5L4br7wAIjtU
+WoVLQudu2Bg1XEkbpmdl//HENO2+nOSvV9N73bt+x/EMZeqe+x1clQ1M4b0xnJD
ltF48K4LXjqa6oVeDCPMws3Ub6+49z2v40WK3ztFel0+aLupFsw42oHd77rQB823
8TwkDAaSpRNqfquXrCo4rM+c5I4q+uiHT2ryE8gp7IMi/OmLSN1B6SA+hbIdI5ez
C+zHtD5dcvHsvaoodNjlI2TSv8wrhWSV9/X6W4T2LIUbv+RCSZncmVkG6+GGkWzy
xxpwOE6heH+2U0OymMI7KtbHLDprYvdnfO3/93AOLz/wJqULtdT2PjzUCUFGC3vV
t4WpMsz9hKm6huEStCwSQDuNQy+kvd0iabF43CzHgj8rHaCMtqYVH2UAPjDBgWvl
F9aZdqQJmVH0i/cyxzzOrwrF5pFKv8jmA51Ij78si8gm5dmQwW8vV8m+ERzgrA0M
RydUH9cHa0936E/Zp4tR+EfBUxhdZZW8nJjF5Dab4k/fEw9xrdld9a7I+p/txUT7
ddo5+6dqMTikUafriMMcWscnpp3Zwx+4HME8zlSGP4Y5F+DLBPH21TY0iwmbqSmR
d3GgdlWfmdx+8Hqw5dbpHEyeRIBDWMv6nBXrSfwaqJb//IA7AgfdlPFiH5tggyec
8RdlciVTyKlRaNykE8oFqAXxJzZG2k5fcmkWjXGmL7zeFNJN5yk350FJ3uLgItUC
QXFZuSyRUkJXeuRn0JRF1qwbCXlHarPF1CXz70KaitcWpUMPhHVp95jApOUGhP7S
XIkiLOHdpoI6Qb0W6Qbjaxh2Qay7IB4onIkdcNaiAN9958qHCuVKjzuwTz65P6G5
g802dOJdr2oU8vwYkxeNxC1OxVRMOr+ABGwQFolIQlptyNpCrJtyD2AalOb4RA1X
3M0oIPktTHsQVi9urVR2qHtjq2a6IdDc4NJq7gEObFc1NGo7cbWdMzrnDYsqyw8u
8/ITfCxVtUNFVU8aHhywFtneeWZgPJKwQpwNiZq/zEyyfsg53VpjlT8U+idoHMf8
o2XPrIzNk4PlmMhp0+E6wC1BD/+36QnYGmFkXl+8d1pqoqoQ0+hufCwFDTDF5Us0
t6J6vOy20ZMsIgNLl1f12mg6MvowVpIVfQiM8He/k4J2guc/6LbgSvVsKiBdUyuI
MZug61UDodx3iSze1k21p44VCeiv1UdiZ1yYZRH2cI73Giz0OhpcarvEONQzZtyA
ss+4FTmwO14TMwmi9UWfSFYXxSdAg2sdvBil0OOwvCMzWZmCrVmFh4ZSn8up70cf
+qPBMnnZRX9FplO/FGwzkiNdJtt/c1NCD9slDt7mO9Qp7gd/37Ho+gHIqFAKqv9a
f1YLli4OaVHMoKCEysSi1OQlD5wv9ERSedr0U9NRSZ9kc+GHfzWlba3QxEcgEKJB
0R8MICdi3uf/lgeyVbsIHAvOcu4+56i70PrUdOWYbS//CGCjfD6Hfd3ughCS9hhF
K5n8z9qmMBIwtazXQlrxu8+sawdTkG6Q2P5VMxLjc5s5J2Rt612TjtjY1A7jWoNh
iNADLBiKDi19hpqZ90OOCuyrzuApLl4PjTSvni9+AUwyGgGLJ7guxQpfA+Kny4dY
9TLI3PkyA6zdkvgRpUfHN1xKQ3ADidkqwXywYzmwpgOh19zAyZcUGsThsYznnJVE
7QrVq+Hs8pFO5hcUiUCBTO7ZU5HKRJmDJ/L5JwAhcxJFfjGDr8HMD/DTHSy4rNbQ
lPejf370XeNND1YS8DqVMMTjIEZYbRm6783ms0gr92VpyL9pTh1urvyklqQtIibz
/jTlchxM/2y89JsHBJuPxYrMGR+kJV8LkqkxF2VqiPNVASPz3YD5a/jZoj2mT1C+
i2QEnrgpBc6iHyEn0atdLXKtN/QkomgIpHMCfakAGR9+D9ik9UOietbYoMX4BxcY
9OXKCP4eZOEYnHgG8HdvJnkJxOM4ljU1GeooeDJQCP4BJY8aosUosFFAWevYnVUG
Mp+UkvrxxIXBoJM9s2ki6qnayJS49eFaZeVWSPLjbTDaJYrjsz/O287R5tWwZaSB
KD4ns/0D8gIjPhBmV/n2/3JNGhZvyFESbCErSIQ4OuYJXH0VvM7wVuHG6dCvns6E
6T4DlkBVLi3tVTu0sSugqh11XaSGmyXX1a+cEnJMSwNW66MSy1WKECFfrnl1/eAh
aFCkpmXqcZj76vLNYt7J1bgWgDl6LeTSScRBFFZGlSxWfu798fOlLQZ5cjafFdx9
VX9IQF65SFGa6p1qLK97hxNnZTesb6t3GCjA9E1h9g0ULdWmlLSAF1FHF9yOsEvH
H1RbMN1UghWN+pgQyb03LFaLSxQiWvLdWSjEtnwEjedl7tneI42qorjy7gVD0sLB
iX9WX6wcIbRJs0/8Mp7GmnkqK1zdNnOp4iWbEncSRt2poDjN/YS4SUIg2y/mYE02
ELU9UPMKG1SkE8LlHBun5jmlOJ+PyEWBRnVOLYkUb44ySlKTnqUYebSbMhtdOExk
Hg/K5KZEF0vPhP4CQEJmsNJKBODqPzaa/CWvD88VD3h+iaZkRAAZwUuQxfPM43A+
92zS3+SNRWajViQXKE3F8Bnw48fFQqyEH2Ed7i/Ota0brTMriKGuSQqbW1k38rMk
leitoRcOtWG6XoYJwB+aGnBdk8FdQ7iccWZPcxXCqNMv2xxknn5MpmtLICJ4atu0
2ZLI+HlUQdrWW9IcBlUeqDplzyWwMWU1uqNVUAiBAxxmZxp+cdcCBXs8uN9xEme+
dPSa0lODNCvbOMTkcfYhRj7PZzQRvLIHmItG6c86/46iwxq4H+9uTy8s2PK3NJdT
KuiGYP6fvq7g4JXT/suJ1V54N/RUC8k9+LieKahi/qmmn/RZd9V1Kdyv4OfastZY
+gAz2JiJiFysY2she/F2qXPClMRfm55wrDErjZtBTuUwACZWOIcjCxu8XOeCkn4T
s9wSLGrIFEm/MSNCI3LKM2A2ZqVd+8l2SxlU4Aos5JOg2o9cIjnp6ux+kjFFT1xj
cH6VVNFxeCJqiiD8bbMl5QPhtIVLTXoHuPN65uRtkbZ5bfLZUIL21aupKYOjbZCG
ydnAY3wOFm6G+YzbbW09aHjeehgkB/jhkRBxhXSLZhC/K/TLeamy1Cc/9t2b6Ne9
ayAu4aIpP8N/cW6uwkmmsCh8WLZLhYxZt8z8ds71ayJjhpKaUpz/gtT3J6Uo/2hc
UW5/j6W9rnf5/vB18sX9tNZGxzNTe6bj5pHgjgT2I/WJsud6HCwkhH2MwrFpFm1q
0qnGdOG39hIKrZWS4HIa5fcbJlsmthQ07++nDh+uc2mUkYD1Y1MWtBCO3zyJ0y5d
3OueKdPnavviD94r39hhRIqg7cshIEOj+1Qvn/QxQ9moM8T6AwVeRXtABVGh7Aly
R0/xev7YZxWVxywVVJ6QQNhkxmDKm3sffYlQQ/G5Cb7mDdNkIoZAbWW2ooAXJ4mc
heBlR+AcnJVEsP9FxwVLBc6xl1E/c+KSdprY2C0wVd6Yp/IaJIxBrop8pqmWyF6c
R+KToOvbJTZwcxNUjUu1Zi+sR4mVgf/aet8UeExWEjPLHuEM1g8kEGFwKZxA/xZL
L5DxhJCch4CTk5E+oeG5Hc3TIzHyU+SNWUYPz5Z3sLAb5lbuLZYC1c4LWpAaxIy3
XOP85Hd+oy4QXzsKT4xIofx1NSB2pIP1EvQoWLbJPpWM5Whz86gcUdEl19LZe8nl
kqnTeBSjsOZsMDLOBpx4R5q6gH0/kQoA1KJ62u3eW9jBA3nzO0ClNpfZS2dlkxue
c/KPomqEvz7ISnpoB/yZVUoX8lSLopd2Lb/DjzJYgh39av8quEdZ+bt1nzVkUUlP
aaTw3/hiPuwPaH1Fpkt7NqjwUuOACelMdfsHTjCXP27fLEnI6F6BlJd+a8C4zvgm
3bf6TmPUZcoMOjfaDkZb8Q7zwvCSbbZPtGeDf7RVue15OEwayN5Foz2iy3tGhJyf
3ONDpYjilnd8Yr0KFhjHvbO4EQcLuBsSY/bsyY5QYN8m5B+Y/cOqZTY4+vit+MyG
9TmDALD11P5UDDZmOL5uIHevFfnsCKAX47uQzOQTxpWMJklTgOWjTVrYfLKhvu6d
xkEW8kt7NNCro5QH8Yu5gkTl4eZd1G/ha6nW9xPKIK8aGuPAqPSITzjdgAvfSlHD
vDYvTO7CxbOAPIZOIxwh1QJ4lGddnBwb4aBqg0O+8+7VXweuBTe4WCLDDWxMOwEc
Aj7PzE37R9rokOwu/4MJ6kbZu1/41bEs8UY5hWsF7lWPSDcnnrJZR5HHZKWuXhd3
xiuEjdxitYxcCfKZ3LWPTnKNdk+UYFJdBsWrSN2JwtuO4q/+jI0Oqq7HzH/P+B09
r/dKL0w3tkKMEr5rSSkVz2se46k/Ggrh/EQvqnvfbVvrs6Fq0FYBOWhhHKtrO1TE
8sKr8la2tnX4YYTph0Es5CU9+9Fx5LlptZYXbjCxyWRXaSF7hJasOXv5aXN9gHa6
x+N7Be4bGiK50AUfBTpjsSQ/E2BzLf46tOq/yf+vD0Flz+lGEBR8WbaX0jW0lPxC
IHOquYMfEUL/Rc0GG7gaqWU0AOThdeit4AcVOBrDTtTA1tx9MPrf+iLboOyRYPuf
AmBpyuqCMMpRCBIFcW+UuOA25fN8dGv3qHVqLRMmfGO9Oat2/OIi1WOXBfwo2bx9
kjNvYRwmHXi0crI28SbqwjH1Z27SzpAWDlRlsJOHDdUMeYP9AvisaLr5oskvXNC8
VhSi1M6Owx77y7zyZC6OdMq3qQqarN7e3KYOaOm5eftV15f/ba1voU2brYu33y27
tEMzKWXhG0c/N6uTcYrePBD9pERL8rbK7tU2kBbJg59WG+xJYDR+JpLHrsCU9kvR
zqJREt3PgQg5POkZz/w9ctE0LjNr8uMLZJR0KIbxfAmcUCmtdfCicOWOgHSVgIg+
hQBxwM3SQIhffCBSintVSEgi8QCogJ3YEbi0RJ48jzGGrjoi+f8nH8E/egmR3Ejf
TiZoBJhpZ+PonfoVyvVNKiyrsComCOiR2mW0gZvpXz7V1n2UrvdKrY7/Gxwe8dD8
5NiHNn/kI2Z/CO8K8upRbI3XzHuNrM0BkOv9DZUitfbLwX9Xuo3xvDF3IQdHkcZS
+BX4yDewiZ9LKpTtMxsjtpYbwIkMMtigBYec12U3IRuo3n2mTWPoruaSubVejnhL
IQ2P6De7UsYI4G5+VyjJ8JYH6oTGwWYc4aK0n+CSg19j/csL3ddaf7v2pq8TNyyJ
pivwpwtuDzPOM8vmVEoy2nKz7l+YuE2ctPHv52ukBVNJBpsKzzraEbNRrk3yEMLQ
g6S7r4BqgGK2KTBb11KEY35Dm3xUPoDOypmfaHl9rTAE7XFPLR37cWZbbmPOGTAT
AxPe9cB4do6Itb/06pTj7/u8XREV10JbpRwAEOCKApDp4D2rttSnLw4vMu5kCWb9
nhfaRPPh6UDn+xr9hojHLMNMtzrAG/soOknxQe9CSspaDeAPXSQlrNGYfz7FN0Hc
cEa9WUH1KvtOT10/w8rJxMedqh8RC9iR8FLY/uwXUb3iYhXSiQwMElaqu5jDFz+h
xkIJaASd+mvgLnJRA415RTvfH1ClsKQ8yFLQV0nW9NjZEYoIket0kVZqYB8Hc4HP
fdVM1FLuDAZTqJZ2Ay1LsAgWF0L6S64iSPydbB0jLrNQNlOWAkt8eNrs7mHFddiz
G7vmZ/Fryq+2dxT9STAO/ulZdTUCAkj1YmXrM4xzyr6+Gxq2gOTRSrOef11hPugp
3ww73adQappf3wEB6YxQ9jo6S39+Cw8AyrQTTpFPjxF0a09AdJL7Qc+vJcWJn9Nn
QyNayIrhcRtMVu4E+3XkPdTmEN4nhaONURU/iRcr+svLNxUqvWfoYilsBLYrB0H8
LGRASPSJMbi0faI9HIvO+WmI1Cdchi/8AO+fBnQkaNnSGsr4Dfe11Z5zkJAgNloU
51ipPopdU+x4tRYW5EEVGSZXCY1FsJS3CFRzOIrDWB+2Og6I8mezzaYi35RgHKOQ
R5tENTcpsLBCF4Qlxkq0+9zRmSbeSDxQYtf4U0mBpQsVJ4nM/6OvWOUg/W/oPnq2
BpfUqndc8UJ6nW+QpLt/3xpbxb6Nuybz+gfP384B28ClPfe+7V2mGYl3AFd7SWs9
Q8iBPIPeGY1oIDW+iPFSiMGJAkaBkQQUtkwB2vSLNktbXjP4U/80dhORDNMMJ0FZ
ype9M1jIZngg2NvjwIa6f1kVQZDIZzVnvbi7BmP81cmPq7hznQSi7wjOsRqLxWfZ
xKNaZ1DgsCTy8RlkEvaNlXRnWngFgnS0Vj6TQ9xF0vacoVcYVXZKDCaWQm41k6VR
Ek8I/kSRo/7cscxtKsXcvjWnXY6TCDhwlaVkbUxI+RksugQWTTymvaZ0QtaSg79A
GDLShxvbxGgTTEeh3HbCefAhWN5kvI3psX6K6zulUcuWbDdLp0hnMzeclV4OPlnL
e1mDlhs50LEMTmie+XBy3OhxaZyvWkDoiGO7ruKYqiLGNgBkwfqphBeV7ofb5tet
m0SO9QmnZrpy54PA9XGTs4IRfc8qpAe5vFItV12aKxJv6TQU/0mFfKviSL2EA/sq
hmNvwRFTYSQXpCHosssGofB9twHSPL9GNQXbTfzvNxoZEiYUG8sXlySWh61O9wC5
FDftYod04RlipbFyegRWjBTnkqg9HIZdJ/EtfARYLnJtqGozTviRMr6jQD9/UbVc
WHalKVMInynhD4/fZMD06D0JolmCW3CRCbFlz32IImO9MsW+nZc2WbYc2pJzOQA7
8LxIJepL+ly0oWlX794x03BUKViXTURKvQZjeSdH53uS/GTo2msO9BamJG1BNYIM
udNSGMZpkBK3Ucg1q/s+5Y5MM0HtR9L/hjKS/NxtUZnDJL7Lt/LnJLRbh2jTGDfY
Z7ePWLnK/dxuH7MLGT+/JakF3iv6+Os76zAVdEJVhiqSC+XxcXOcPMpvB7qzRPnR
z1tQKHLViOv8kyptbHoU7T5dxYaOnWchdLB87UzmTHizeRWsWuvdbDeJ2NwXLsgk
CUDQllE9o1ZhJX5SrbTJ6Eh8opUX7ROfJ80Mh/rGf3FHeE90paH7aeaOpnc6LUot
3N/UbSQhPyjPWaJx2ONWw4wHW30P7UoZ2mWfnERpI1nPSTFznA9zJrs3gteEsfMW
7Sx92ZeWGYMSmCmorSpvENmZjjDgA5KjHCSP98nc+1Hdqzra814NeasgKGIapXUB
goDbl9J9eNHdKdGBe8ESF1QJZgrTmQyhR0/KpYCKaR6QMFLbOLdaMBg7+rBP1jKK
pJgecy1OZOx/J4DZsoxw1A1ih4/8X0g2v3TehSxOn+e60PlE6JnDjdEWZZ/bGMLg
qphRn8FUWcf1fDdFvCBmaBZdBOLYBlNh/55NZGkSduaJqHppZWLBkj8ge7W0T/MK
CumxCUA9Q9L3aUoJbA/RH0t+uXf/e+ZFOrTvvJyYs/OnUDFU4S5zRmko+lpMZ0km
nVM9bCIOyAWrGXrxvtSNKNqzpAZxQdRsyDp974hUpAZpSlY67tXojFDFjy2dJW28
+my58H72ZoDaEIMaxgHIwnNoDEn1FKHXvbyKH6RU5NBRIzMkFjH4hDwfNXiGB41h
/xa/rYNxKxr20VHuhzu8I5aDAq/dI9ADJv2FQR2lFZVDAgn/uMIi5m37o7WETAVc
rjt7m51wyNuHdBokGje/G5p9tk4+hhbQnfMSD5OVHterL8GmdrzPVPr043Cuq2cS
cI3coH32kjkk3rupMunszgILFwvx8YyTZUH1WZGH1UmiDfyXYLwCqytarc63BTpN
SwHWUES7xtYxSnxWs2hoYlmlQlVLDumgS/MEYhdgruLFAeKYSFfG27goJXk76EVU
XoIFQG3g9ia/j7auCCvyprxtWs0Tqc8WtosJCirMUNxoM0tOYkRXRBlqM8gF87OS
3cMEt8V1gvHkQNv6EShxNRo8XoTaHes62742l3lFASbrSX48XCCDbvkTGx82N+EL
XopVswD3/ml/5Gd19++Nrj6Zw+E7tdIJvhE0hGazlt6g8KP3UCb78sgny6Gz7EOG
DFWtpP0X2t7akJ4tD68We/hp2RdcBj2KSp8+XiDlbEYUVxEXjvbeeMLk7c7bXMxH
ZbTLWRlxsmjGnsUuE6oACbGxGzITb29Tnh/FuHxKsC599wG+mjUhsbX8VgoxxLSl
H+DYfraAXH4aAEhJE+fWeHyWeXm55su3R90/Nu34RdVa4/GRADlIoaAtfLnaxPbU
twG0QIeGYkbyBH1K4KcB2geZHXNd3dJK9bAbDUYGvg+ncVLmjch4qzHmzkZ+2Mxa
DawfPi95SI492l7DG/LPnMQ9G3KYb5tSBWXHzdkanrrf7RS36oOPiQ1ZkOm2rJWT
Dzlrf+RowlmaIrV88jOFDW2cwDlmYEOTYHA8X5bPDrTBHnbhE5ljcfFnC8jshe0O
Ju7zo/1jNOze55ZaAgiszAEpm7PJBg0BjnnsAAglFKZDWS0tRUm6sbrbjBRiwpm3
l5QIQE6C5N38ALyZd991l6bD8rvLy6N46f1uxoPv2FW5YORIfWsIjDnl4PIFyolT
cvmU7GRH5KYIroUbTw8IFNyfJxup/IPRB8D0Z0Wb6/DnkG/4wfXuc+SvalQ6+UFE
8j4QvT/SmD8Jpa3IblEffosOP/mXAAe/1r/5/1rg54/WSSUn8uFykaBe7xFHVx8r
+IMcFQIJ2s4gOwFc3ezmaoBL0mdbbHC7TubzKt11VGXeTpOhusAXnrpxmr4tA4Wf
tCrUsiUooTjHH4vFWj2YmgqHufk1otTM0gn8tuNwlZ4X9hOtWhiQuGnvokiL8tG4
PVhDrsVhH4Z4WIsSicEqoaoD5BHNnRc4nIOjhtnUfMEMd1hXxtA6q5/etSbBT4YM
+cgQXtc8taEkSDbwhh7SeSKRKfg/nyRo6hY62GIVAl5SnQPfbwP9JiA/td4QbCpV
DA5IDD2+sMX2RJ5KxPVi7lDpN6ptlUZP82O3GSVtOUPcRfl+hgPbJH9uvK9c8hEn
sohdsMQGLo7BMcRkPCHa3W6HmevHGA71jaNIlfvE7eJkzeHyFKbFM1Ynsr9WFntC
Xo8zA8mTmvbm0bwYBDqzZB002Ixzp+7QqoChuqC83NdCaw8ozWQN9s0WMOl2WkkY
FVzdkq5+4Au5AqPI0nZv6sLFaoXPAm4iY1nWTo5yKEzYDlsnkQJ2TO6YEoPvhJKc
ixRdO0FJaoTmL3YF+uKihV/ph0ZYOUjrb+v6oNhfgE97wysRweqAYloRzbvM5yIU
Znu/LCgLAusbOHIG666sNbe/9DyYzl+juDUeWwdMLN4j/vyYGpp/j+92k9F0vle/
6cN/3sWm0O6/bsfXiIGz8g7ctmiYg/j5Vbz9MTb6fsq/LySrODn4b0xtFcJZEO59
Cm9ugYYTRSFPQPm/4UJxe5gopZzyyKQzGCMaE7h0Klzrhqwjgp/p2tY0zrC0TMMq
Nw4qJK26swAAFgE2ErCzFCKbFCkblWgl80wd9Nzy69/LOfDHVGKle95DLarCXezo
/FSTBgHk5OU2n7hQqNj/ZIdC5/LrOf7tT0TeHpEfIY4dl9+FZo+7DhXRFJTpN5fi
ezMff2dRwPzcfrZ/qsxidaRbUAC4Jzcca7onogIds8mUBmHOyX23F17PpiCeyOWr
soAuVNz9kIRBo401STeCBUs9CSQLCd8yry7X1KfGvYfp1t7UjVdbR3kRk00Suli4
LGwTmDjRQ9aOJWjHsAMZhNqWMctZ/fZFdeWez7v0yHnyApaaDBOZtuxGdIvgHTjH
YNsQb1mciELOITC30VCISPjcrqnmXjoRd2OSeU50wP5NsOKE1lAPPQBRDRveh4Nh
gPl5JYdN+N+4x7Gyk0CK6pdR/AtyTvSNO6nCbSnHpF8cCNylbzlaoSSUOSi2bDUD
ADIqzWqE1z96qsgtgrF3wvBIYD57NSiqxeT0uFBGmjNiYk36GripKzlQfIPc0zrO
qPkVMfTMa5C0aGEnsSeHWeIkXqcKw1oU00yTeT4yVy3hQNDEeqp2cxZZGa3cL6up
CyJugK1QncoU4pkc4yb5/rAtiQK3AW+IK6G/YXbg+mZkqSDyYet7hya0fv7zNM5v
cwkgeXJmQEkio/Z7cGRXxbVlzatwI0EglwYN1rTWGW3ajgQLvs6poWthRpIi+WGK
WExgiaYYQgG+2z9NtfgLnfJkWvdbPVDVtWm2U15l4U+1qfmx2l0mCwNArvKA8zLn
7moJb1fU/qYRY23Gvhu0wsB1PJZuwCGdehqu00JZkC3ZGRXZnw1i+Jjf5LSa7hsX
2Y2XjMkvsLTy1jUzfF+sPjxPfKzh7LRopLMGrYgaAZWl6ybox20BP4fkESiEn2l4
j+Dlk7Gys2mwc8/r/czZMoiS/Q+CPHFInLwPznjCFSyVPitqFNThNUQETSkPt3p9
z3cwgY6lyyNOpZs6nnHbsFevtRTNXxpELPPtu4NCUAxEc/U2qTS+IvjyVn9IKsR4
FYdfE11YG/duey3sxz65V0FIbg0SLMr0ejDTkQlG5DkJ9cqwwxxpjTdfumlf6mlB
bsRyFgFQFEiXwpd4Ot3+T+SYhhR6L0UnrlXeQYQqiOYpn9+7YuGxhasMRFedukRB
QpAnfTZ1wTIj5ldhoTgJrgj0g+XrWm+WMX5MMX0nYSaqtXcz39QktjuxCObXesLt
PIUXNfYls0uTrA6W/zANI9yW9+OHmjXeaByb2Lp3eDtcIExBo1eTnsvmpa2PLkP0
+OGbkkva1FzWabwxQJy0J+kgsdOdZJdc5a2+0nHmOtbUyxtXTmrpxfWAJALDgxQA
hPilslRhHoVKXqdweIP98fi9CUJaYRyUHcd9enUIi3GYANPpe/SffCMTt3ITO/mD
fKbukw9b3EaDqoNa/QEUwWyB2GyIovZ5t6jDUuXCrgZ6G0gaDZ/3hfmjbaQHB6GB
qD74/aitLhv/9jhhGy/4YcRhjj/CGVERvOI/V7jP5eWikGp3Vmi4+tlbyFAbnTHE
pnw0NtwdZ4Vn7sBT+6WgjuGPunOSztjgyiSvAKd236bcvqut/OVuNUyWo0B74Jpw
I2lKxdAVg9cvcCn1wdlUVg3IUxCh6RFov7e0D6eiRxjDb8yYLn+M2k+aoW/rSRLx
WPNW9QbIwVcft2p7Ye9FJFdWjMOI2Xoy8PgTx8DERZ0OylqaKEzOIrRPv1u5cz+S
dZQaF5yNMEc8bNcCks5jNYJvU79X3+VkCAGvEM4qCIk/wYHDqOGqtmkHI3XdIG7y
bVSaGDEZUrJg8qw7s0fLqkAS2FQvjPKsbZWrdDWaYFVDPkOK2PoNZShZYOuu5Qaj
54ayilReMcL7L4uGmTfilBJT/Wl5SF+JGwsmSjG7FukkR50QaFArlnBajdoHtUh3
INdtYoZt9ub83tX8l7Av8PxCRFo69IUffWfPN6CNKB6zCsgTULwPfhj8c+lIBHAW
IHAS3iKWde62c7+TEWCRQaLS7rMuYNDmrhRhG+hg6NJfd1/jENokZ0Mdzlvfak6e
D+J7taLV/1d3anWUWu492RXv6eeNlf7gaziBBlsrE5FWSZpv3WbU4k0Vk4hVY+jO
bn5CTSeUkG8rnf122x8BGb6h38Xr7gslMoH6OpQ3Hv96GjP/yRaii8CX3jToELcJ
un3/TNPuYNDIlUWBw3VtGeIjQpPBUld5WidBrC+H7G+pM6pbflTkMGIgcVgOYsPT
XfL+43X6/nn9Z64ee+bpDmMBkAr6/eLs5JJrPXvavPUomPyB7hNlW+s3dY1Fgp1T
XFrDLK8krKEgn9ec9EK7ZfX2TWgxGue/Mx2frD6oKNxlCYsXDy9VZC+8l9S/l9Rl
3w8bDgVzDcAgtkHdTE7m69mP59TGFQX66Mnz+nh8gQmTPQCMgpM1Zhfdl8COLUdd
jN40dyBLVtV1yPIHBtA28lpzw1wjwWgWGBsldKdiZO8XRtOajKTtct9dx9rIorbA
KYDYYIbZ8KvqVz+WxoYbHMe6FqNQLK/TDyjL37BDYRaCbdx3bfboI2r8NjkMoeKG
XU7n065tQzSfKNgTfXjmjy2kVaqzObu66XmRtZOpc7t0Ilkyk7FmxdGJSkjxfSTw
cA+PcLwiTeON6iGczLwnqmvXb1bA2TuH9NLghW2lkSSoc+wlQKVdTFH8JpFOTv7+
dpOngVRm6pv+CKqnONLct7Uu8ddvR3xD/Kfd57jq5tcLDCTRIV7+RfMmvD7fsDEE
hX9/5HCH63rONlFNDaxHEtrmXp/RoZBXWMgl6KNlvb/FkEPGCU1akWrcFnA4HUb4
hG8+PKZhEbLddz9z4FhIutWl9kMK72cnnKgWzR4N9EuWmWQurUWyakwS9/GU08xH
0DjMdQhjqPRREg5j388Fl5XiKnY85D7487hI01m5t0qgjUCwzYACpz5D2/pF6qwm
PoazqUYhxfpxVi0t/AwKGEGwmxH5L97t6wgsKIq3YY2654MG1iEdHvDefUI4esxO
dSD8C9FhI+YTKR7efRhZ5SggvXNjOfMFpLNsZHnecuqJfwFn0tUKumAGfTnnWaYj
ZqCBItegZwO5A5gw72ZMxW0WB/gZAt1/e9/dmTmAR+67KLR8nJKK7ZKGwYLWijhS
J93HRvLODlBLinQhxn1179FMOFubfxcScUO8MPVdSKW3KWf4O4ScT0XgvORZ+vnA
9XKGu3ce9xGJuY/9GydZjO3AYWySe6fSYB2lqSewh/EhGzU0/UEqLi7iNVLFSgW9
DYLWrR11RF+86WTtE/LjmXG+JbIQLMdupDWt28dx9B8BoJhs40oWBbY/Q058Lx/7
UcIGnXsBdYvLTQpF8zqGsCpvtJqvfhyZp/utrzb++c9Kt/EMmPJty8w9vdv1uu4W
2ij93TO0vhYRVr6A+Sz84eBcF+AxOwJV1BfIqiLsOvNoTlkesapgZKa4/M+9CCL5
+kCOobeSrfFMVAATI+JOmuyz/daHx1h8PUB5vw++lMwlPXxhNjhpQ0ed7u2Z0O6q
dH9rcaqRmvMlpjlIaYNS1K1cEkP1jw+ynCfTEMJ26ydFurrf4Gk1P471cF8HzLvC
LHu17NBmlDTdJN5YNDoybx3IqrocGlSVIRXHItyTlHUa9WH3gw5ssXWEJArGrG98
7MHxLYd4C7ArD2ZRkoToOiO1+eWslRUPMaAQibkiSsETdNgR9l8rcT09uc5nrGzX
x9Rp4yqq00lRqC9D7hy9mGn3b6CwYtB3hZMAbfbf6BV2OzKvepg2bRkGJB3/7u/A
acc2ybyL1JB5BFvruuKBGeVpdO+QI1Rz7IzOxDsySGGI90AGlmusbhn3rTU2qwC5
tgzsZ7FvRTbGlcBVB/BpKRj4gEAkdH6kqMU8vRz2aEe+Cl5NRHQUpzxtfHhKRQ57
+pMgYLxuIBjESO8rTjTq6j51qwHFji3GzR1eFc6Xuk4c0yF8d01EPeyBMhfg/Gro
7Dgk+Jbs88YUEZ7uDDK+VA0UeuqY/q3QxE3+JFaxTQ/t5jAsUL06kRk4gn35XQeQ
oCGHCKZ6VLLmuwLGLCi7RsKvChZoNRXaQkufjiYjVQCJ7vSTlxh/nVctF7sPSSso
wLCyCwDEkllXTmP/8DRrugoGuAmNZWDS93YlXqXTj6H4l2Ag24LEtGSXiScLjWT6
vnYzsCfYIRlo9ZhyBgMBOs4c39QhkD4LDFUxENvdwV9T/bPkJgpkcpqOjpJyZ5s3
fVJyEis5wp9Fk3L/Fpunxt9QF1Dc9bBCt1isJsigzIt0RDFw4ASldMgvG43oe/CP
cjw4nZpwTocdL2ROLkYiGghwEolPw7e5RwlycvXQkQBp+sE1M81t03q96FRzvkl6
M3odqrz5xEi1tVHlLyM7J4yDxPTIiMSX6TFHxb1NpSDeLinicLdtCBe+o2mIPHzv
IHfvYXVcHRbTlBugXv6VcoIBN5sxNfW1mC320H3i6t9cdZb8/uJX6Jdk1g+OaO1e
U5TvqNJPtKwtzD8iF58fnpn7l8CXVjIzzbKe8IVikpdoSb0aP+yTW9kWZ/FJirNN
j359na80UIv1zO9BX20ftjpoyBMbeTROqyrIsknK8ZkNXxpjJqsuevOyI/2B1ryt
W0zJIv5uo1yEbG37ynYbkQC5vTAbMT6aQSE8QRBLtMbKXwDN0V6hI58FO45TVxZS
ijAieWqZ2+96UN+yC38bqa51ebVPxOW+EApk4wFubMM62MVlqb4bOdw3mb/enHxW
b86tCa4eCa3b5ojF8ZmEHZbJMbxfli1OB9wTs2XyPKUTBB6Jp6NdFgwkfkZdX8TF
03XkSgOA9a63/vN8SIUKqb0T2TDRPMwXl3us2ngRrwHiIDcDMFA1+D24pB/+SiQ9
D1d/iMD/gHY0bg2ZpM9BZHtOJ3pf1heAasGjKUfFb4FEGhXvSNIfrJGkBjW0rInF
qheTqeChKPhfRSddu9a9ei/CFruzSO5i7FB/38mQ2Eztjiz4y2jwbgHfZipORCT1
vvUFaHuIgo2Jz8Ae0079EHyhpYEHtw7RyszAsvl81UnQgE/CsSWJCs+NrP13WIS2
8lJhhLmK3/uVIUl7wbX2X5tz95lekY8wOlcO9r3rAdJkJbnfLlzXRIrSZfM9DNC7
EZ9b7gbXigK5H1T+/6A2qHhMjmG++6YKf5W/14o9q2YaPm7kpOIXM/4OoriK3F2w
UGikIudoPgGLz1UqEsvr8XOajiwzmiVhsW2rmrttJf23D6xz8r+MnDZjFhVZLfva
lsGO4ziG+AJkEVP1Fi6ByPD6fgse+gVt0KTbZCOF4UMz0lMRCT3iAll8Nun7A7yK
NXNTbtM4ajQgBSGlvXJfz003mY1wV7dj90gFRFKloe6aWMYisU0uiCPERadKHT4l
Cc4eMzghN8EucUTT1CgJIa42zK+KqfptVp6U1mekzlc2qEVKo2zDN4NkHOd1FlUq
wMEF3ZvRAMgAsT3yBBeQt3NPPL/8SUMhKjdmsSZE0Aufo6YUTOeW+2v3PAwgw0uy
I5ZV68JnUg8paZBNBc3WCM171My2+5edryR1BROSW0O4BDv+qm0pitxsZrNxwMtx
903qOwv82ESfW+uEYuWhxAZr6BwR4ONVBbRmudR0nYS0JP8QV7aMu+OJrmzjKb4a
Wo33luXbNxABke6kSkoEcWIRemyYhTOI1D3efefuop3ewo5mlOp8+27UznpmFTR8
xNviyzKIsl2ZO/2S/UERhLQlMmCMOpPwBKAwfaDrbgzD1+OhKfgLo0ElTm2MIrVX
5G2mfHh+05H6dhXMWyoQaHXd2Vs0Gnfpe6ov6bI2UF4jFcHyMLNj4my1ISFFl3Dy
rN5o0DHrlSxb2nEghU0A2CqcI5Y0Owb0eKOEql/YC8bXz/30GIszyzIhmGGczd5E
WfzVI9XqaZYze4/vQ1Ag8iTWjneFdInYRE22OdX+40IzqYVJe3RqlC6n91hAVeq4
ZFc6Srizf6vwu2BNWfMYmupqne0p+N59KEK9jAdd3doV1+gX2TrMgpHWtXAZRtkP
tL4o06Wppg2j5voRZXzznfO2CMOkN46/U0q6ez9bvjYgb520FM8t+sUZufIwi/98
0/TeSiYy/zZl9cFZNmsOVJvuaHc1diZRgRZlfD4mbNQz+TExp85WL/CxImX4Yx3T
6MQddIst9VYoP0rK5LZpKSInXLp7k0go6gwgpcU2vZQOIo+zphHB45L2x1925SCD
ix2/Vme0NSP2zhg+DnvbGctAltFqDNO5IndJyjiznWCWPq6N1xTsREC/hcBXegTz
DZuRAYOttCkYCIrs56GhUkw6Qz9Biyr0Xd5epV/qC62QOHTGl3HdFD1nrAEnzS6s
7i519wzQjVsbyyMqUOtCKrfyyPiyP2Q94aYHRnF5ZUvxfZrsufY5PoEMghKC5TAf
O5ihm4CXEq6F+SbCdPKB+8PpTVURQUTHQcLtcy30CHFuSUTd1OfffoV4q1mRlRqz
1LtYp5BcVfLnKpS0pe48LQrVCEDfPw8rxxJrQ7HHJRYhkd63VReZmJOV0guplbaB
iYaeEbSSVEtTAk0UxY1ETclswUpXL2xohyufOvM1I18j0MGqUE5dDW9nkIlSxLwR
rHQYD0ILm91pgi1wO1BSHr9+tZvfIc9fb3Oiw6yVTrGffoQaXvnne3smUuOc87hj
102JqL6Z71ZWkZ5SpQpEyNN2I9UOB96bD4+QVyD5AY9GhFhkKwg93/qhI59BU3iD
F1wNSu7tkyiCuH4m1ImxSzz0dFbWlX0D2AgsbzXW3vFg6jFNlFPhYGifQ6ydFXpR
K0v8lAunGmL70T3Hjo+RgQLb/IPXVGvLT4nh5iDl/h3II068J4rfEH3jOISQ5EPp
p/uFLuY/ApiJXdZiiWbCT+0CzOOYT14wACKZSlLy0bSDHWu9KCigi4Dz1GU9fHa2
uZ32bR06UGbr5ebg2llQpWrO/gydUMaY7Nq5OZPTy6gea2jYdTpMd4E/6neGmJ+b
n5CPMWbnbMT2i7rMQplXnikHQrPBDwVMv4wy1aSx2J3UoZ9szHRkCvlR0giAveP9
1AcC9FH07/D96Iw713yNi0ntdxrxtMgctNa0h/+CXiJf2EDFFQ7Uj64COXsBgF8e
wlJG/oOPb2kU+k0CISJ0ngzDpcfuRPRkqTPHtvc9jWyXnQHkL/dcWeCOhM3Y3lxP
x2FOr2as5bfLDnoJdc7B1t2wTszNj+oVYw8FwftS04aVOSwQrQaXVHzIZ9+O/e8S
vKuz6zL0whYleSi9Ge92W3fT5ucJQwYPet/G5C6R9SYyRHQCSDUnGHyHRPsNIYIs
eTDhWoh1pIx+Y9EHiAY718mmZYMIzsL6Su/TQ1KyYq9Lg4gU0Xl51wTLYTU0wzHt
qFm00KEIeg2qBsLymCn5MJ9KVA6FAZvaGoC6e76fXqThkW54AEFKl8opCU5E/ObZ
I1Q/Zqwqjenp54d6msfSPCV+r15ts7t817Zt7dhQuRrURGwqXG+QkO/GKceb1SAB
4Dupp9FSuSRvZnfUXJU3Yd21caKMioi7B8mgEq9VLOA0+4CEcTO3PIXY+4qXtfLS
J3SUBAgkApLy+VgyyMpE4FPi1ixZfBrHRfAMIck6c1LZYlGEx5lbJLZ8K1egccly
xOu1U7E6bfips7JHRzvtSVr70rsCu9nh1gaVfvRW9+Og7pFvWyWKldBDCMaqBdeS
CspgR2KifW6XW8Jx8L2Sq7KNOwyWuui9fJHL9KDugks0nOh2LqVVctuNaSbB5hjB
gAu3NJ9XKVSlhnlH7agaRXdwOH8/x/PXZnVPv31Ypi8r87pipbLSBd2MBCWXDrc+
Uywj9r3c8EpMQZ2nZ7aOrBQR761qznE/ULR5I4P8abxkE340rxptN1+j52NJKLxu
oDjqBA/Y0vyvq08NnYaSmWq2u1RMaK5tHecvrBs85V7kWcIN/fiqdw1OuHA/Wica
jiVgU6cOnIr3a9GlZeP421X4wdc2qT/wqRQce9zwu/a0qPt+BfyiO1pxPiJrgBcI
f8gmhGS+OrCkiYxoKymz4mm5b0iDiAstvz69XFIW1kozjAGSvIavKNg73Z+wHHlO
X0iT3ReAksi8aIrWhM/iOb+ebuegviT5XED2R88u+4TAiJXtl/0MwvhxfYhwx2Qv
yy/jRJMciKLSp1ZFBDcEYeY+ym07t4AQslU3tDQtVH82osuEPxdqAYbpU8KuKhmw
wOvi1hO6dDp4s7mSt+y6OpXD9uyJapOBV+hw1lwFzc6obIJDhc+dl1QOABluOecX
H3EU7HmFWJVFs6tMORLrGhgjbPOa12Uc10UZp+/ZxA83PhLSDk+1Z2oqVeIQxKeH
p6opx7bhQFh2WKWAN+tF1YuAar2+Wo+Xt63H6xJNDD7nIeqZK4oAHHFXcWWOksNf
fGipiOaC5OYCiqCrSXbDDlhKugWHn++cdiABOkq2uhvgYzMIOvoSm/EeDGxloeZq
UxVTHQiR7cT2TTqUddQV42Y9goP3C1iDnfEUij0Be99ksmsVbSneWpk16k+NnYiV
xZ5f6EiDyogY2pa6oZQTwluAU3w3/rJGyswWYarf/cQOKcEregWjLK9AElYLYrdl
g5YwJP3K/G9A6J18yxgi58oR9KctnklnKsdWp8fKg/4mGY1WRFkdwR1FVRGRHJCP
19oWgXEDv+ebfjZjDKEtNHdLk0j7wgnaum96wjigCFvY4gdiPvytYasrMoDDB0tP
qdTO7VTs4RtQOAZddUMxamkGV9IjNiywVwNhICHLn/2m18yhoxDqhAvTHztDWHzI
y4LywTKdAIxbsAWc98iMNXu8Enx63dZ+EiJStjCkfNxDoXUIJGRS5fXy8ZJcFNXk
KdWoIAy7CoWi16NqyXnN4cKkhmqm7FbZTSR0DunHVO9fm8Zh9XV2C9oDXjZyOpsh
dxSeQXutc1GjCfbWdyT8cgVxWGTmnZHiAJ+SApotFzytLVUPoqo9btB/iyDhhnKe
4RKlmNYtaKm/jeoJkBdcgiLN5u9ZTtrv0HXRpF3p5rhDc/mAiJhM80UnkEHRRy02
f9kqVHUddiILr+mq4aiKuCk9U3pHtEGqkEYk2gZJzrCauAKcXj7YUeHiqktGf/F6
umNv48krg/eSjf9lynjBjbGgytOpqWBYa5nNTyeTRjjUM7DXUhrTjLwahwJ9K5Wx
MYrHhpYwfqaBmdy3rNo1kg4FU237Cg1W6yRiMkQ5LtypGJdCtWOY5zrYFsM7yyzM
cPiyyM7zhhw0KV96iDvPYDxdJZSCleiUooOJLnlie4ZfZlU8jvVUrX4JH2tTOsKR
xNyCEfH7Yc/il8QfxWoenkrCiEDK+fPDyNPS8CnqD3mIcdn1tzpCgFoWaIaNlgD0
VLiM2dUxB/ksYCBJIOGm+jpI1wYwY46UyQnZdspupkjVP8qUewnJ0runLzEqZ7J7
m/NuK7tbrwO79DV3DZKWoUzIVS78YdyHZlUnaoK1OWi0qu8QXct/991ntA/enalh
mAxV0QSOunz8eg6jYMPtt4GaXaleRGBF8P/gA4upDNWCBXdmcqWQsalZSQ0FvOXu
9gVXTVePi1ao70XVyESsd+rg4Zx9qwOyfXTfh5xPWPF7lmSxCCdugyGS6V3XS9SY
C8gq8rSX7g4hb5ut2kSRxJjwQF0DOKWGSIII64XfFGpzlSeEgdD3gIPTmyZFIOlh
RsByLWZtLncQKVUGi3P8VHH5q3qnmFTe0Yl/mYgrAEnp7utmJiRawYX8GZxrPzsl
8f7dAdYgcZ+L3PqDHc6Dq2dFK3u8Qhv+d+/trL21BwT4O1XQxLQMvcuogQc8Ewq5
8ZU7BHkzs6JNQ40VjxvEN2D+lscFYYirvHhB7SEA5sgf7HT7D/+jDD4ME2UcdHzZ
VKzZL05txz8sya/JXzK5OXPn2vE4k2MxCyuFXdAjFOnxwPqCQTdYmhfvDxVo3oUX
YCI4BhU4kiqw0+DHeF2urtSUP2H9LmvDyIioZQyxsg/A3P37pcP/AcPPbHZNM/Xz
4SeR6s/g9sp23VIqLxoaFSLfyHVuRjGctaGX5Wi0P8yOvtCuO0dIop/DRcYsZibm
Njy93v9wYlTZdsUHuTeGTU2xYyeFCodXUY64eQWXtMc2mjatkq3W5+SOHxsj7J5V
qIvrWszoIj4dbnbqd/AVOyz90UI9SioNltk5t3qLzl24Y12djGuuQcXCwZWsEUaP
vvGbH0mSMMBKBjLfjE+CGiBqFoo7lVHLWXpBPvsiGvnfh5d3CKS+9ulNSXU4cUrz
DDIhvggSbNZ9qF/5nwk/IxlC6IuOW0Jk4QYQWg4OFWL/KSIE5EF13z6kHBEDzk8K
xbVFf9b4VadC5rnPkDLPmnpu1AjngHYI94PyPaByb8W5UkUEDVASYUCPmzJ+WXJN
OvxHntNF1YZ21LBpBUebwx2TqcCfMPJkf82zrhLsbA9yLqLJyMNAmtkfUDmpCBSg
qQZXW/Ir97MjEqRQiqVTrvl4dEPsKv07+qL6/ePQbRdHPRTExYjGX2Khi5gYGcwV
/zU99wwnKrtkdG61mT3ftgnLn1muNK1ivelFoqjZEd024gc4E/U7sPJyWb/tyC1+
PfytS1FlffKDT2TmWhFDBP2S8YTepLDWiCgk1yxaPivBbPymVQf6uK194Hk6ckXh
JiIjIFO/DaCBRKEwePPtuw6M3WTyi1j15Ujlr3OtPX9cU5yLQkJCYDdRzqKZgtAz
WSpSRIaiQ247QHgUjXvONJpMSj6HMAprLq2M676b15rwJxJOmSGXpBrrSCFn7iLF
lk0NFfFgxPJpcKzF6rNKIUqoAYoh/hkPS8CeFvh5w2S9M+x2RQS1Ufhz/h02OtZW
CihDAGsjRN7k+vmtswGzlFQeX80KQ3LoASp6B29QQDrdH/6Ey27K0G/dc1ihio6g
NjeQkB3fSfO/xeS+eIMG6gquZE1rKL6qauYkqkNpn5mw+TwjMn2kqp3pXSMuNeBy
l26h8wwrwiito+RQdhVIjImLStt7MWwY0UwZdxHo9PZejugCnydTaTrG0LVTj8/n
H3LwfcnO4XdlxLRkiPs4rtsg+oRuZRZRExxu+1b2DWg22PBDUtfnIXE/HVA29bz8
PPCymbZ7bzVnyshH1de+WhMoMV3ADa20F+o0vWZOjdhsF7dmGjHF57idkiRZ6qhh
X6HtvAteAXFKpOoZpodxR9alsbgwLkALoEsZW+xJCyhnhvRXcdQe4qDUqT7EDDKz
AZIBg1iTZFnJ/nUC2YhA99ZfL64rfKKMrBOWfeklqIpt38lmsbGyGN/cZB8wJ1yW
7DlSoEPoDh/SXCdBeoxubAsU6xNhCDgcwIHyzY8ki/8Nt9OsCHk+fd/cAQuIQ47D
ovBBSLHKM/9Wm7I9INYDNif1MdLGcM5o03p2WmRRBDpRYCS9DxDks0ocKNUv4PWu
xD9GH3aLksg77n3j9/zWm0EsX1UvTo5HILORxaxJHXgyWipBd623ww57bFP3XUgQ
9e2sfbRJKoT1kTcG6AOqwseMx9HYSm3/habWqPcNjUj5fnl4WemJRpqBheP7uORr
8Kv6Vkt8htgq0owWHFLMVq665k4WAlbJ5wbfZF2jyF+9X1Ka9fpTqL1rXjTSrEjh
um/hQW+lzVxWdhF+ZsD3n3afhri0etvyFNBh3v7fg3t7n/lrkFUIIGokBJ6A4QXA
yaaPN/HQTnKGq8w8wC97wawiThf4JCFkD8Gq0t0pU7kVXynaCVy36i7MV1HK9vuO
eS3VHoPw8qhNLmPfR71JrtiIDNc/rFSDxYAWzIpEirSYvvl8iU3tXeaDLMiKRJdb
WGmyXyFy1sYU/liSvO0bHw2APzwyGG/CvxRbiH+ftsbrjwecHiIWxhmRjt/8enr1
PTO3xuMf7/ggf3lk1shUfF98QMD3tIAZDyrh9jA1XD6NJdMyVvTEEH8/xSkJcaYd
uPm1Ztryyskzc5aHrdK2b4y3hn7IW6fNP7HzysvXKxrFN9OZAgPqqN6ZLz0LZ2Vn
hDurAlCedXRBzT1T+vcYiaNqbsVFsrnM3YJ4trfGUCbZuoSpvrz4DHDkjEf7ISsP
Mg9isBGnzh6zxfF4OAC3mxoNMYi9ngBeV272mjg8FuY+DY68/Ola9O/j6oAt+GJJ
/ALyfj5MaHvZ8dV2iO9SN3voe787tRaDuMrf1zI7+g0piM5UQ3fvu5GlRdXF+w0c
fbVj69mFHKKV6ZRDC5CMbLX+5N8Jx26VxBHVon4/mA3FSuYk3GGkImt9ef1BXRJa
KKDPGrekRxZ8OsPTuRQn4MIrybR1k/z9o6bU5jmdYIrVULgC0SHw5lfYoummVEV7
U7DLOiLWOib1PZHZUImRsbrflZ6AhMi6ezwDeuoOTlbbLUSAXbOkheU+vRAQkYFv
6XPgUFR7Cn48xFmxT+TXB6PhfPhYbPdr6Z9aNz5QW1+D+WuoahKZeGH/fol1KekN
KbCF08KSHrk/ldJOjMmGdGHqyBFa8OQewDqM2AV2kAfWCs8Dj309kedbFXZ4oZku
Zu7KpInulz7BDcTFIf+yruAZosSGoHdzZZUw6M/d2qMx1cg5vIvt6AN3dWmv8OKO
6fsYhWynKGD3h8QGAuVYbzy4ExhOVa5jk48XD7nbabfATVDdLLYkE19+psIh3ygu
rtnqid76yGU2yND8BiZheNHzsGCXB28Z6uxOJSVLefQDQPYSGqUORBvSSzjLI7Pz
zUqNeVVTyEpFYjGuRGsoAWGApDXbuQ14L8aJFLyF4s/qDT4lU3SXlMpoJoIhUyer
8KssNDUh43T3q5tC4jLJBQvI1yLiKOv44NCM94ux5nqMV7jkncyFKEEYNVs3z6t6
I2Gy9DkawAScX10ZXPusugQ46cSHXIsV3RLM2wPrvaoZq/jWCeitvVX0pPJCs8k5
gdnf21/jNG22ZXr35+IjXiqWwq4R4cK1jj+MDKWZcYqS18MzSGja9ouzge7lhfiV
PRmlk5Gr3ZkNu0/2Ryf7BPMR6Xt6cYL+GBCzvu4UYa+cqb3g6TZP+Yk85cPwRfhu
tUF4Y5mOpYSlMEhWT3u23TXGj+pUmYMva31g4jWpvxlnFSaMyrBkniBrOU4A2WhP
MfVDT6TXBvy69LyiFkhGl3wAyGtRpBKyJGrpsOzQhzGIt64troFyH7ET2hAeklgr
mdIaHO41sz7bdQq0KvrIIGBHKf9Qu7pDWoIAs0J9nrPaT+QF/tHV/05avrMkSXl9
g2dF+nlAfRiQF6k9bWFhdREJTWtKby5OGhsIt/N4qTSEm/02D7vFcIQg//McM5bA
CC9ad3245nVb4kasHabuFMrurDBEM4smkTO0oSyWOR/Rh3m3fiSI/L6G99zt3XkB
9QIUrar4OhjnFp/OnKhk1uH7JTvm1n0YiO6KvAZ6fdKY3aFRekZ3BrkRuXmshF5r
QwsQVOJOqgXd5M2VQyhsgXWEkaAzqFcwkqPTq8vql4ucYq4ZATHPK1I84z9s7LGA
nLpMpoV1BhWImMxrs81aFNltb2Z6AJesz/ccFogjE8mdr9hYtjGWnVw4rCZRp4Xl
hE9Bv6JOxm0iGzC2Osd/AbBGcWxdkCGqtubxtUey4TGOKUUguB1ejU38M70CSiaG
0bnC7cof4FBbwEzM6DQIF54gSZOtxqfHRwMEY/4FwfVQ7h5OR3MGknSAKeccHMPJ
YtXemEdk+WidNr4mLF9eIeaV6Um0TnDLQB1ZfTmiW5XxV4DnH9+/a1HFpLfGHR2u
nkdVRr35hnsdpMnB/SM/Ff+ZalDi8qrZTeokYfyU58PMyac0ypalu11XsroVUCnQ
pCIMYv5D9kkCpoVazZAVPGsBH5qfzy3br1t389C5Tb2MzYNg8G/mh+2NxWgsYZqY
0M7SC7O4qez/Um1kgUsWLf7j0TaNACZKuM6fgYsq9SMfmUFCrkWsnyMupONz3Kiu
a6Pyj0z/aQRT2OJnq1npgnveYaFJ1PKoffz78ECpTQFtPW2QiLrQJv0DRAsRUIMj
QDH3mcuz4H8+7Jkj4+bxbXs9hGtNhQl9zORTvZmwzcRStd4z7XHksieWHvRCH8Pg
UirS2NJzlGHuk+zQ1Y/gTngytnECTfGg0Jrp8GXeO5wrA10JV0U5rDB52TWSvVN8
uFWFoXJOZnnND8ysE6mbBcOGlzOa+ZPjBqmqvPFjjuAm/XSz73n3HokQ6BDC9e/U
OgVZ5J2gamP1c007SqNauVZZ1vQppgkuM1aHNjKm6l74gdbSbV45LGKIx4SfwrPg
fYJb72uK5ifjq5vPVSlIzicz/5K61/I3pYJ78ppiOeTcOwbg+Alddmtebnn12Y6w
yRktXiHK/kOqAWSlcPYXXgkT4qUu2xC/+D9tdrXRyhdSKfJXTzqGZn4+QMKWT5C7
30d4yc8iFwX9EvvguaPhKXUkBSEfKBA89bSkHsLYMtDVWtqhgirPu1M11KgHJNW7
UYdUN0WjmZT1WVIhzYD4A1ITQep3RySiJHw98vFpWw5NGHdJUWOV6mp7KXJ+nimZ
r1sWrIsOq7V37PXO9ioFTMHlZcuBZrJJHfT2vva68vRnld8TOYA1JyaqE700nIw3
eu1PCerKHgW2LDewO9hkMTtZNhxoFnuYKjCYIv+qayXXxj1nHu6OO9EfxMPU0dj0
e9k0ZtZHLTKNBd60dvUIzdgcUvyDBFXj7o0UDpSgcW6uPHTkTMjO1ZoNE0s6tdYz
bAr/ImlJvVU0gsDh1K0iMvmxNjBqNKwj07ngBs194PLg+IhUZvOObb4ifDC3PifT
y7U1ZR+HR1w/azbbp/QGJW5yQxLuldLU7QRNHHi6dUXZorBrxLLznUcFmMuJo57a
EMrX1KWRKKmZQb8nFQTBSyDSwLe63xaV+p0yU9//oTZiawxDQ7WqlTNfURxNJ6/F
JnFL8mm5q1Fzz+J2VOk20SWKyVPTgILgKJ86IcE/wXpAfW629B+Y76ECy/EhPq/7
qeuRjfaMnR+RyzAOlvbezleo286lcc672sGclRJ2A9NkHyv3QYg9DZMY8aaQ/yHY
+0GrNQpglenFv6Lx+a0TZftdFug3g9sHnpUIYfSIhpJJVCJh97TKuJ3SxERRTC5u
rmnMkcYxuOOGM5sGAmrmq70dC4GEXy0DeQajZ1uT8X3L8dDlkTgoX+Q2bHnS7gJi
PVZ5WlRYCzzpt6tncyL5N2qSO+1rBZ75QnVVTU5zOchJiN8+ab45x2+9o/y8zcys
dodt1RLo7UQUOr19adP3Ce8d9pI8HUviudKrIf9YBxg8UvRXWaZYRHc6TnbxCvJ7
ECKfW/jNS8NIjOmMdCDQMrTCtJDyRkmQVkHJ99AG/onI5cj7o6Y47uDYiDsMUQj3
aa6tGtQg1EtLYMKXG2nuJ6FLNdKlocdnf2HuLa6sACnDezdf+ut/iihWI28Tbzlm
Kh8sjt/gUgPRXfKmjec9Q6rWMFEEGzkkk65OdHsBEwXvGWiyarq9C/lLHLCxmEFu
JcF8DBhm1yVCGqGPO000O8gJ10g2srmJWpwxpD1ycNpWgWIe08aRCMYf16BLwtNd
XoZYaUwKhJp/6gnKi8dhLxN0eMQwFrv9QoUhKJaXNgcRnLSShrP27ucs/vr+aHBV
488Bv20vJAxuD6w0nClx6LiibifYuJnZqXGGBlLdk8Hsgsh/2MzpvvhMvyGLbrDr
i9oJ7u6hDGzON80068P07UOKWvmO7cy3FnsJ3mRXw0pNQHgTFWxXvFTJBTJSgbkj
mp7xMr2t1N8x4ufRtUaYtCdwFtB0FxAj8ixqf5rPhiHi5x5qMlOW8IBSRoktMqs/
Pm2aovjE3ZkDh5XNUSIHE17Lfg4gNTcxCijJtA4wJrEb1wRc9A6bTUxshiswm3wE
uf38SVeDPdOTi8DayQN6d6mjiKER3LUEb9lukJCAiF1GfLTxlkppi9RqYoSWwwOJ
ygQ0EtUgtqh5SQ9IOMcCu38HJMKbJibkQATeJCVd1MygWwH+83iMCNcrvxrbo5ig
s0pJhUEA3BG4y72KhMrv5mMpjVfHebXaxNHsEzrL+kxS8s4ysIueQfxZlk3OHT2b
eI9l2p/01exCYvnR+O1cQ3COU6vnQ912CNvtRGHDgVKI/FxJGKGvDND7d0Gh4xoI
oAfqIP6VScM++IxKf8lWwz5TiCX+2d1/unhjW3NPlFTd081Ll7hC/3n3OmIGHNyc
xFq35+ItcJmHMMCXI+2a9elP/3Rye1vQEJ635SRN5kyyvKTYwX6mwsNfjIOFUxF8
+FhpZC3CnIIj9dSRnk0psU/s/raIbpZ3PcXhZJyj3gsfYWwI9C+SULKbAQvM/0Lm
rks1pAuoyyb5/3OJm7I9SIygXueOIG4Hf88waTL09lFsZQ9HPWb+lPZrRC1d/FX+
hrQcmsG3OUY1tpWpG6N20lUh0z9OKRBd1fphXH9O9mClexRB/Kld3hgf4G6K9tFu
I8vJdVhOlrTqBdNuWMR02AoQUYvenWkOLVZ3188NF+dLb16hVhR4e6wCbGToS8RQ
XftpDYxTLWzNxaLQTYUBn9IGptwFlzyxc4Qqyrm4ZZsGF8UalQlABPxXX6DP3f0z
5m1nfWPjbD7gSP8jaYbe1YWMd6+oc1KuHZA3GAjSkr/nsqlMFcAksdwp14QSz9VD
SDYOElQLFHY88ye9DU0hFOOlJx/hGhHGMAFQixnW5C/MKuz6Sl8oAdtOYWN1ZleO
ECKT7BPRRuzXX9NgB6h1RtRCObZZiavnxG2x2ykRkq90eIXvotgUkGKocfYkQC2r
oThdCFVPDXp+FylKaHsbW32WG0Xm8E1QMip17aydvvid37l0NAi0kD9u/Qz6O2R0
gkCLenCQJocLQMS4wsirHN9Bqi0vCqYZongKHHSdBUrIYS4bxcK3Siivu8eJ07k8
qzu+Lf28Q18AxJU67tnCMusOV8rn3kf0BqYmk+uaYkt4A2Y0sJyZGs6+88PanVuS
70a7YhdnZhW5kavm0QXAlj6Ewnq5F0J01HLvjDWcGYSxEUwTyCdI1LIyXuyV53Bi
mcxwrmUcyzki4P8Dqxy1mUh+9UUfYTK3Jtl2C6+nGZkIMrAqoxGu9kMGkqiKoUrs
Aasw9ttTJrqy0rJzY5RJ7gblBrBKs3PybDoaUVgmmLlDfT+u/SaRm9JkCjsStL22
ieEHcSUy4lrGriWtEX39oeqzISBHRpCqrRQ7XG/oiAx84jMBglfwiq+FDwaP0mci
LmvlAZN9Gkny8Vk0LfbODZbPYm7dr6MYsUpiAtfuqlKXEQ/nNcZ7vzXIANJgrus/
K7sYODn8OtGN9ruBJzg05gDSbhAkRRb+qQaiosdfbaln4hgUGesQBtkFusEhnwxr
QDCmyA8Ti65ILIIxegMzpWTeFQSxndJ6ZxKxbcBlWYQqBptOWa1EfBr3HEng3Jjx
KVA9eE1cCXJl/hKvXnnM68A8naTOKqLvMNLNOFFpHxrjmrzBVCZMF38eeSnviXen
OV3qHRx7g53ZUbwcBGX7Q2fFqu22pV94+asUDPbAPa/XmWG07KpiQL5JUX3jwzBq
mtPG4G9iHEQnxAgR3dm4Xw/J5+9yb/mgguM2jgx2aih4qsyOTXuYsb5NBv9Bycpz
ZCmc+OGHiEEYq5ob/VQpYKlvntBQr1GD2TbVgDygRKL4CHlnWsL3N/JKeV/FCqn8
ePWaqg5FIlhDOpWst7x3bJOF39DqMzJQdjJF4nw0mIj9q5ckxe6GZtEnJ8p07f9a
8ECxctw7sQ2E56Aop2DMefmIU5ujcVctf25j0Ao8Sj3uEG+NqSjFWLl0en4D53s3
W9eJ64ZqX2dM/ijp+XjZlYObne9+wiBAIehSjt61EVUKRhXsHHQHVHht25JrceQs
hDF3v0Lrzv2/94j4+WlU0mhZWTAYlXBOMa/Gajm3Z2X8PmNC0d//p0YnQUXxeta7
53ZyL9V70OdA5kypnEXgprx2hnOYj3zGixrzx7J+MXeJIiVze67IDi+WqJe0bkM5
iRQ00R7ngvhtw9YOlRTQfBz0gWd7Tuoa7AYK4G3XDll/4vQXc049DC8io1+bHIOk
kU1rYuXhuxi9yCUaCC1p9OerpjkdYkX0x3JkWdO2/M0J3wmZe2BTZGAMdRl3q/E4
irxN6Qq/WKn96pbZ2p2T7OsddKbWHov5vg429nKLZe0vOPqgqRgZLEz/KpE/Q4Um
5YpCBwuDC59+/tmsoowbeIHCXlczjBRIc1I84T+uiMO6FTYJtTHugWJF3wpocDDV
ptHSniOtdtLOwvSSTJjvUsBmlotK4rVwz+vob7mkal9PMeQiIc9UNWyGtB58bDaC
a8qLnRrNVrbkbhydcXBZEFX10xMgrofv8fYpXzl+S1CdC6FNJPEwGtWoYq10iguV
V2lZbHck/go4GwpkTluV/iqi1sQfpbwJG6Ljt+7YPjzWQ27N3et8eAX2uahYAyet
HXsDWLjTlaG3fOhrXn1O6KfOwY7d99JgqD0SCVf5oW512IghzWPUEUvRJb1oYjJz
zqRp08mLSMTmsLhaenR3YurH9tdAkKUku2K/w0L80i3oVeNuF4rZijfoPgXHJtwK
Fkti19UD8gkoyzCtLeqRhxykqWZzrGm+5nzTa5rpoAnby8g3lF3uFOMNSShcV0sR
TpQSol+KwUrZq6+ztT59spJca8qFERUGm6yt2l4t8y3Mf9cMUze8poxnfDGy8bcI
X0o3c+FDsMIlpOXibQnEup+GofutWk6W91Gxmmx/8cEHbFk2XUQOzJpuhCBnqdkj
kG9u+c7X1L9W0e3DwS+4fy9OaM2YSYf5Y6vF1cyit4/dF/dx1mzyFAxnovkSudgI
Yzg835lpJ5qmiNIbAwM0MopLxvPmawgLcQfHYIGAWmDA/X4GRCAHCmpC35qAhz73
rW5Xz4jCq+uuWqoSLz2lPozl7v70BQ4zOUmIOVYTkkAyo9aEkEqxo+wYBjLfpGpV
qBkJj1KXpia8MP9kf8z7HZsM4CF3GNEWC2CNxdT6oOfip/uqgdkGmApg2XooBk0b
vOL7tc1KM0rzN6+SOJDm3bmGokNaLQZUMzZ01xyoIophWTdHNzrfrNPO2QSUtQ7k
cGul8PKLr224yCTyWXQ1rDIuhJNh210F888O7iFooJPq2xlWzMuASjd6Np1Ns6Ik
sf/hslODZG83lCTjfSIspa4hLYTf7qI35NitukQX/DRPMbp14Nuwt9OUkDrysCjx
JSf4zjQeXS2xRwzdbXEU2SpLia0xsP+bbo8JyNeyxCZVEJEKBx44tdqfSrkZ8FH9
7xe3drdcsFMS60J9But08tld5RXBS00HScmJxlfhPTH8DwnZl6NX1q+a25XfytUC
0ytKGLOWjB0TJTU23gTdpcfQHXNOwgXF71kEV9JIFhEMHZnZxoLCJ8rfoE/29zEY
N0/6+sRg9Nb25Z4oj32CeDwBfopqoV4eVmxRG1BQz8WUGtbAdRfOKHoRmCrbxlDA
2O5YGDHzBcLnLXUATg59psVIFp39cBNg2gy39Rul7vIGhd/BzpE4TzpDbZpQ2bNz
Di0QJ7gkouZ5MjzEJVOJmTm+B30OqtfqedKU5/qhwR1HXntmjD/QR3VgObeTyY96
ILXmn53v8SA0+jKXFM3/RWsTF6SCt7935qbBMel2RnbuKZ04xztMCdq/WAxqgTpD
znGHToQLm7jqHrlCfBYOV9ipVaREJQRMSwMreiHwQPZo/mdqSenokzkl90nB4ugC
gM7afNZ+4B+acfb7vZFoKicIQuavMqMZMJn3nBPdWiXh4EDebFPa0QyZmtIG5TRD
upCC5JBOB3UHD8qlhTLphzap3Iv8BSwqAygwKpGQ+v0QYrnch0Ka6GUvkmJ5fPPI
61JfHieSldda+4mxu0eS3ssB1deooLKmSSSXlmkB93V1zTORFdb5bsUSUXi2x+KL
/CXY0M7OCZCD1ySam312C+96rRKN5+raOvmF1TSMpo8cEYy8eMfaGyjQHrrcCjMj
GSNcqGWGQssJMWtZK/OYgMlQUBsa+3qv9xUPc0nQA4MweCeqvxobQ7XDppmXY7AD
JbivSwexQppLOtWZ9cMOqktZlIekqMe+oabgECubo4zZX01FnHnvv2qJce5RUup4
qGHKd59wCbluQoCZ4GlBcwQEMXJUUjop1eLXFa2e51XSikM75K2ho/bfeWqvQoIm
k0msbn9z2A7f/ClWA6WJwjB7d+oAHf9ASPk8c5+P4FNMnGMPsFqgOSNZCR5We0gZ
p6XIInQkkD5gsUwoFPJ26WLiJo0Y/EcVC+0z8cP+dpsj8hukjLqElVODGOhbf3Qu
KNFf4NztfDvlOaoRzH+VJi+QTwLecNd5rbb6aJftrSSJn1lb5pzIDSw1y9TCh/vr
cMO+n+PBuFUsT7veCLayCRFGf50EmuN9DXYRYw9W+2xInt/jdC1O0gOlDsdOsUsT
+JKE72fC/bExepd8GD9vr81bWgLhasKG+7rP0VnPpAMg8AzPY/MuUuwBXHLgoErc
DLFuzO7zjOwxKSJDcieWjXkRw6xBH9FhjRbMTbWdu0KqXuqmBaFZkmJPafU/YLEC
CSKG3jyrZlQqHvoM/oS5qnXPZMN9QmPzIu5DJ6H4ndqJ8OQng+SnAxyK6FQF4jkz
KQCt2ZWhKvsifjm6OkgvBGKd4F/j5cAfTKmbHL3y817w9AFDdLMjTXbEJE9CNZlB
E8sfz2PMBCSZhV2xiboDHw9TaNhYOiHp5Gq4Rs7t3nI11ev/LEnXuEKiMkspGkwN
8WUxQx/dsMwNO4Ofaw4ddWC56Zq4ulKOwgq0w6WmDbXDhMCVTTcbjV5RAwezSDjv
8YWmK7K44lwOHAiK8ODpnA1BGJ5yvSZx3J3DS1bnOR2ijzTuJ6ZimTyMeCTEgALY
2WmCyF3NDHEy4Q3dUzydAopG1SQM31wLVBNmUThKt/gDhuv2wa0B0YkVLDohG8RB
EL4SLbZc8tZLhmjDPd4WgZ0Ho+W9V57adE2mzqQn+3ZrULftTSVRTO+hhIXvUaOl
bqtCHo+JMYwBkrxZk82R20BFzoFlfJJKVCBeDjUQ0/JUHW9hVTReBOSpZaK2FWvB
W6UDTiSxZL6COIdgHwXKqpKJzq/NKRakh3OonSbc+Vte2EK76d8cIXncWdwWgwwM
ZAcMy5PDVfpd8LcAg7dl/PM5RaKhC9YBJBaXiZ9//PZbTcI+OMZ9Qe5X4xSyuINc
OzsuBdkguT+l9W56FbESGtLuTRN177VglqMzD5HVg8jkWXw6a1nemFCEZjBd1aQW
7ZJ21BEtsYsAtXN/eH/EvzmEIyk9tWm6+uPSTxNABS9UmjUTsX2Cm2XO61CrQnph
wegikbdpydat6Od8zKC/+Rw8KoZCueVbmUIWrn13VVD86RWxjjHtNjmbHACmveQM
KAvD8Yy2GwWAwXn4VhJ9A3ELdTW11AdmJDHVnYAsPzBk3kPN+uSyw1Nz9AxFR18Z
f1+QOXRM5c8/BM4YMWvV6IG32NlpgcxPAMPI9Bk/Vnj8aT3XlcjGwpc13rOSIecb
2cAx3q3MTK8Llgp8yy7Wbnv5LpEKXfFIUYaI/6js6wnx7IBtcGbc4OmAQ/agBY4j
3XEaJNhL84ocpairRVSsLTUpgtptip0b6cbK+MB8XCbpRAK2RkFzh7Gt4tfxuMmN
mmFUNGoXbE93XfJRedmTR3dUn7r7LpKGYgdhDjYc6Pwyji+18stxC5H/MTvTlVxo
Df3J8aDAuVbGL8SFoWF65Vh44MQ3sEk7MX5SYHzaVtbBTuzL7BofTxtH3Vu5WB83
ai4ssZIeqB94hWhwJHe8znHxGXca7bbvscgiZbOpjGFC20KDbiTY4z6EsEA3arHG
msgZEEcnJt+XOGWTKy+/zCAezLz08rGik88v8cMCyiM/xLWbEol/gnN5J3Beg9ev
AWcJi8P0MtvLK0M6aUBe2Ak3aJ0s5yXyr1pSCdxidmVK/e+8C38RjKKaDYfyPVHt
tlf1LNkg5NpJzj2j3uvtQpvAseO0V9rZSUEvX5lhicxASjfcWaRCA19CjrIt1CS7
0fEC/XLOL8hUE4Wvnr5BMBdnMfPm7R70BsI0gxZA2crDZJFjVCcUyaeF2OVUfhJ0
HkmG/MznThdO6ys1BjUHfRM+eCZQTZXUpW/A0YdDZEPLXZgx6W4fKhGKI2VNLpFv
0zOQJTTOTKuuidmzcyMEqUGkuCkL+zVs2UOEuh6Lhd+BmV6Bx3TjawBnUiyEo/Bi
GicyYxq2l2wEThFmMfygYdNtDD7HH/qNm0dzrst4ma1i9rCq4WdwLwCekVmQHgUj
slsvGyoEHTh3iIKMD5fiHQ6M/i+4fSh5tQGS3qTxVQ8F97Qos26893X1zk9qKQcV
pkSSLBe5mFe5o8IMVkYxFyt3Pj+FmIO8FXvWz8DDcHFRB8oCEeEJ3er366vn1Owd
pcdizTdwKl7SHnacg+nWut9wxrtI0lw+aJgE0hI4ZSCwQsjDrkZK3Q+nxm3kQ4y0
Q6nrQ5+MWdAWszjoiTewC2b2N2Jx4gaYZO+u/uJY+d5u7VupIZOetOlYTP2Xm/Wl
Oqy+YWIv+H4ieIw8OqLwcdcMRyHd3xdzD8p1MuOH6mn6ChU8Iwxr1J/Uq1ob5XvV
C3iEoNlWTpec5ddAIq9h81eqkATDtcJlyyzQZL9RsnMttksmNr+XOmrIWTpochP2
ZI60Rqbm3vk0L7C36LOVEkwqbUypRhYDf1E3cjea9T7gn9yuUN2sNcmGnM8Xy9IF
SS26u034G49uZhCDBtfvcioROo92HY43OH2ji0GpjXgkYZBuyUQdtZyHr3jWxCwg
qtm1P1Iz6dW6GoT74Kmc48jhbGnBheD6RtB8OtFyumaduLaHD9SiCbd1ThRjmGO9
30Cx8oJMMFQgLVRRT2DxPt3jrLuFIkML1uaZ/3hKrxkSztw628MgXJtvPVsbZY87
/fsiKPtyus0OI/7HHc9DomY/VAQkxAIjH2VrJJvMzU2eKONRk4jXAAicWUCRKIfw
yhxCHlbCv9t1rnZvMLNz1550wZmcklMQ4AvDFO7838rIPdMAJy4The5VAVZJa8Mk
hnrXBwnsCzt6ArrVoqbTsI/mk7ergQgrjQbkgVBZh33zJEh+8ZVN6cjipg2poMY0
E+qhcpBDn73zGgGlTohXQhwAliTtUXcv90tExktGU3Ph1qEIxr9FoTJ6ir3cV9mV
qWpr+NALMNCRj73p+231Do6ZpOaAgMJxqTPZvjOQMHxW32RwS8+E9hc0bzLdSw38
DfheKyWlKbVzz/PQgwEDWRVkY+Z04P9OpfhWzynXxXSB82KaqbWifGGs5BRnCMWG
8O69cjinFzxE3uMwEC77UrqRBvwhSG2zClUvMOl78d7UwC6rAUTGML79ZkLmgWFy
5BaPLSSShPq9weRCWnQ3RvvElkqh8ucpvx4QIP+GKCHYXFx6jTNtbXSduyrfewc1
52+VwLXhZefzyxYHHU+eo59b4xVuRx1t8K1wCbnRNfNbOOJNNHu+UP1V+qymkt1D
L5Y3y/mrcPZTaJhnQ0t502yC+/r6LqkcPqJGbpeaaKmG4Kz5e92QVp6UfEiOLCbO
GDFnZqTj3fCXPIaB2FheKq0gvVAUNTAwYB+zu7yPTZvm+MRLB/5LhNtv4jFmAUkk
4yrYgRK5wtKpoMHFCXGTBEBdk/aDojZ4Y8scNsvbhk4X3aek7Yo2T/cW4pQBcWqm
emdaGEACss5uc3XzqKW0uKhbsVlIPZaMhCBlzR+f2lPF76msD/lKT6k1JwFf62yX
qeXlLYh9YZYSdcWmF0wre/tDpTdkEPgfBJu/d8iJJWpon65jmCmv60voNooPQ8Vs
j2McdcgthyaZ8OSNMsA8vBbUaAknImJBvHwCSU8gi24JqHVmrz/UUNh824gk3/Uv
gnWnnDE4X6ZXydNgvgmC0TtLhQ99bIKGIwZ9/gxlkQ2ufS8eFLzgwNSl4Y2+m+v3
vGPL2G1V5qfg+GGqDUgmBPqIfCI5BfaUR5kBBfaqVTEMUh/g91ixedXV14BPBmrQ
0YTKe4qJcFEQutvG7b5b20Al7vLfEkLKs9lKgEsfbe+Zpt8tAFMk3WxWhvLWppNj
JG+3x1YRpWBli/KRt91+sxFCXnD6aIOJY8vQWXkl0upQUy6uDxh8bclV/Ff/BbpK
DouXdSuaJkDVtbpke/KivUHmaikWP10l5nC1D55PuK31b8vIHyt1eu3YNEjJSRdu
ldq3xlY2HK+N9a90eAnbC4UrnxnjiKTOed+pDK+legWgvcConNbJ9HSJ9l8yYApb
9Gh7LXYePXOMUGBpBqZpOUsynfaucH8cBGR8teWHd6KSD6lzWiaOSLKj5mkv8/T9
h3BFwD6z+tjjtNXoPzJIaoMeD5o6dx6BKPcB8on8MdROQ8n4uIyNgM5Aqh+OP3S/
ADY8R6WIrrELDX1AQJKDB1vF0hU+lc16pEZX59V7LHQ32PvA3DLjDiDIG4QurXeS
n6u/Qvjk/WNxBV7oXoR6K0rPVZ1/qX/XqYZH9DyRUiNQDMeBdSfZlNnka97EwpkY
jm2UkeHQhOg9OYwfPMUannUuUmpCWVvmbdhLVWPBkeUA29zXv/6YswSIxW8GppMh
tGKOmVLqDEYA4UuYvi1iAfVK4KGNvdS76cTpPvjng+urf2EpfS9gQ/PiH2L8OyMP
+Hnxwd2ZxjScR2j2zSBR+LCNNEmx1Gc18LtXqf2Nqbqqjk/ReUpss0xsaYmAvxDj
Gny1vO4JY8ZkcF0lkAmPo8Sr833hNdKGNwDctZVxBclqjBAkDvt3//bLBv85BGO/
GdD+PIZ3QogZoPW/5PebGqkiD+ttSU7ZxykiM/RwX2jJgSBw58PfrCr+kva/oG8d
F361or9IUF40PZSi+fn2XbEQ8j05W+pNMkzc0ozSHKG8ZQVNkTZ10jtRNwYIoTJO
uYADlx2zJXPKEpuyV+KiHehoM8L78JrG8IakkbEktmwWa/04O1dgN1hrKDMB+inf
s9ffdxcFnxE9Vfk4/i7Y2C7m901LYjJSF3KUC6dbzb0+Zch3T0RYhUol/5n37bko
nykzn2N9PewE6xgmUPLonJnhWEcjjw/OQXAqob9i7hh1gSTCBeME5v4fb3ESckyb
qwH6X1IZAufxwWHgtHCEGQnGP/IFNdFXcmdbIL1i3+KGiNNfXDv1yRQIQDzfSc+A
gjIvA9J8i/lEKBaLHNpVGsy68QrAKjZTqvWBSDHCsvxWGmr+f31+2Ll6OdISDVXY
G4Rz0guxRDZTHa1X73EM2P0OMABY5yUKCTNNCYDdBJ/xFVh/51DpRQY+ZubjT7xt
/lmwgnZI2QLUcj0vbRnj1JPL42RYwE/K6ZH9dYrW08hz9CF9jKtALTLGH9VKveiJ
Y5PwGtM0xnW1X4YeSDfaUrRqaWe2vsYDhSXEnM709u1t1c2ccwtu407qEzEk0s2J
cE+va5bWB4ku9ioZwa1+2RxbhrHN3zU1oxAsbZ3PhCUYcqtmM9sOdKHt+vjiMR/J
exr8skxoukC9Lol1KH8xrt+EaJAmieHJCzjKFaie+2gvmIUoQTTgiR/k/ndy/mjC
CRdjV0LeQWLYoKpGR9R3yjNdH39aG0FX2VgnFUhB+jYTUl5giPgtcknSnyHvJssh
HT2VrJ4Q/rf1hei002tIM/rqyJS3mtOScsez/mc8/vy4LolyrIoP/fZ21v8FLEfT
JVOvADmDbX/O/W20YDDamNs3R5Oyvq+ZshWu9EmXLPJbZD5lDmrKwQcYsvNsVvwz
w/OisI1hVqcbjMALWMQGWyHBkDcaJbmocFXV4kTIsMQ2IeAybUwiWG1qXwFp5taW
PurrI/cfyaqC+j+YZS2b6/uUwZU/cWj3NvOs5P6RNEeqNlgaCZJqxy8G2JYJWCoz
jBZC7fdXym4zzuIIrzwa/m0awHk6X19bc5ZXVkit8ZJaQ3fj9bOPB0YPtzKk0o/J
0SZdAhldGo4p9hopa3lQBCQIkdViHv6dbsSYY1Knw8Ah11iEYDeNeBud9ByzohgW
DX7r+pO6oxLZaOnWQYAK0mlsdTWfIJLK6PhwYwiSNXJvDvc+5UHMKaVGn3oi9ehl
XCc0/DA9Y4aJBkjHrcG2M17JstDh+woXxwXBKKaOyuU/wDuq5xiHxTutDxSxS9Kv
cg3inYZHbzF51zmnXt5XTRIuw8nyZf6/ij26zIc369JYKKpPUeMv8mzvfC5rVoJ5
O2j8OQZA+UkpY9pM6obYQTC6HPmjm+wBvr+yoJSsuffgyaprJv5iGhjELMw48fGu
D6SHkiJKgKp7QAbep/tEjBmXEOOukub9NI/heg8lOqwJZ/cn4jWXbCryjmK3h1dn
is4LTd4c6OanKoNR3cxmxW2rEL3/2IqSenvI0tTEw8Si/E/ao9Q3MFJSuzXb7tTe
Yb+WaNm/rOB+pRe1+NtPDunFXfsek6/W6RF0fynFZ6yttzbz9KCJKK1oJkh8Axha
wo9bmPr3euPQzaMg3biEfxDitfn50cwo/Y5loy5ZGkuy4r+cDPvkTmLjIhZRzDuY
hdGHRsdTeOnOaFqawcTMzles49Mob7dKhnSAG5Bmchq+z6MCVUgD9LlYoOyx8iVl
EmstansACeGlDhDNTuUzXYQtD3uwKhQqXy6CoV+BdBYxzZqDkRlWHz+nwTrtMQyH
fuuFzVxjuJnq2MapJ021tGAXP81iMliojhN56usp9BdvWu7d+LrgoZy1UY+qaIFt
7UPPEXD8IL+kraSTYAAhI/khXQO8mH+w1BioNSJ47E7VaYNoVJBUNFLCV3CJrnO2
b8LlEIfdc3TLR2J1nkcyZiUSCBpA8DMoZthi1pFpe8KrrG16W0ugnWzoY3Xi4rdH
Ow1NL0sozteJVvk1N/neKwTH1NgflHgzWmrhSwORoI+U9Z3M6rqYd12nx/4omXGW
W4kMa3oqW/lhm7LOvA2TeQpf2+WYpvb+Dxz6hqXFeQ19l/UL50s7sfNVxSHSAE4D
aMUXjGcZXzeVxQgTtEbtqggJU0OAb5+UtLCBvzHFX1RGo2gMOONGfy0sTOGIL+r0
HlkxFEWKqv0kGxndn4xeVJ+JXcerHSG/wOhO3qFnOULGQq/JObd/z/SMu/ZtnU/t
OUvHemyLS2Uu79GeiuYeKjfbma8C3oaVgiIg9n36WoKe6TsZmT7ufQtwhezGyq2S
gXi32er2y3vnwCS0oRc90x+WXHsW25jOSM/GN/Udb4b2GmVx5mF7JhBrbjMGL582
uBVr9nC0yDxMsSQW3+VuVx+Pjpd7qopPsYAeS11Uf+24l7+i0BgIuW/cq5vF3kt7
f2Bk0NMuxClBN3YljTPRWxp8YJDWRk9DAcPmUdQkdJzRT0Xl7S7EBeywBoFvPhfu
AAOrJjPUf5iQdXcga/jTShchHPWBS7E9leKZcB6yHRbE1TtM1E0Mb/KlJM87ZxkH
+tJEM02f34E2E87BesiFuUVRYUBJvrLYLVQINpI+apeFRMJ7PO5RyrdgXSpuhJF2
2Th8AaNVP5lW6eHxiSy2EXtnYXWnRV8mNl+4fgVg7IrszWdWvVXgujkIvkxlhajB
XBdFy3o3tofDtmYCEXDXQgctoPOeFcj1TPNgbU5pqOxDwmkQLRWC2TVG7IHRhunA
q9wDvXVQf5ZFhVHYtEaEcWXOI09ASy3Yli4mQClsNBU2aYDbtdTwADPdFv6VsMg+
tpVJowbLyoTEhlN6PjuYCdeTMlzWIemAEQ43Mpcp3rTo1IcHuzAcUtS2EGiNnNrX
lZGNyi4b+dNOVeOAqtdNzZ+AyqvIhFuA2XRqCX01w7PSmt6XHLrC7WPAFJkDiLAP
MqyZjVygAw7KfJ+8CHS0ueLqOhGVYaveWooaaSK9WWYtQZ27q90XpL8fNjSdMJjh
GEnfoZs2rDSVY6CXHAULz0eKKgEBrK5yIKt0hb9WGS6MFDusJQcmNAtbp2O2Wynx
aDMWayw9pG1EMpZNP06NRxvWukxXQaw4T2VVfL0xC9Pdpm46NwQiTZpyiW2qY0nk
fr8JpNeavewXoNCICXNgRr9qTBPB+oIhoN5RkdRkyfeWtvb9a8X0e1MNJPoQhxJp
63VIOpLU9QRZhfrtSsWtg33K4EY0qsk0lMIpAs3GZUhlZNesNwlctg3wzM+ABwFL
GuzVZLjnpnGw4LonnpImJ7EN7mkh7AaTIIj2J3U1y5CPO6i8egliKG1V/Lm/RnB1
hMxBpHh+TNQenfNadi2yGORS7Xa6p8K6GYxVKkLl+3F3dHKcWGmpFGrCXgNRN/xG
+MFhWiNJ0a4I6J04mdF82lCvagFtBoxe40gO4mOrR7pkAXOzI/HglZ3oQJCD5cmO
cMKVM2Zz4bZI4JPlpRBM1hw3XH4w5ZxKhI0Lgd7em7m7UrKWijk3wmIply2fE+er
YcQzrgXpCSqbQe/vxxzL3Ridfr75rOitEV2+Ka5RNxXuW9ifLU+UI/vNVdShM5Dz
1RmcWpVBiHVTIBvgWqkQCOMg7Dk/elAUtwuohoqFlkHjcxGG5+K1vXhAok60qcnF
eAlvegAmwnxyFILcJbbYx8C99FJ+Q9baPJzJDkdiYVxiiMHiEzg1nxypCAYmyT7y
j84OVFvpNZkDbp4463p8BknkjCsGdqEtuLi9bqLa/uoprOFE4sg0HW85RZfmWg0e
1SPLYCEwc2BEdfXJG+SawN0Pq5eusI2LLoKAS3h/zxXUSx0rCF/LUzrCqRzLPyfJ
b8z7d7nLhcPI51XoZP3OKNiKxXaC4QL6iQmPuSXIbi6SOcZU6GRu5KBxU04BRLGk
HtgegiLpJk3KXC623029B97kMi8Fdr+xsqLSW5EETyYBb7CfewGTp0MxBBv4Wa+y
17agbD/8ZXjNdoJZhUik87yIhq/to8HTF3GfhSHJ78vpLDUeQYeOdFTLPoWfHDPq
2fi+Z1kwC4aLfOXQfNpbB0o9FWpASlMTgci1ZWn9wia3ASmUGT80KrQTC74aKUEh
rwYg+dXjpBeeIi1w8lV3ggFiX5nEkM6MAACwpDEjVIoxKfN5HpLvkeWJ3VCLXv8D
asVUZQMOIb27QrfeU2OjRPU6q5yNTR922KS17xlR2FeRI84DZqc6EPY1XMsbC9+t
b1YcGPPa0hfYpX0OyufoFcPg7HXnaPwEnauCw4bt6QCvca5KiO+Ik80mc6lJxROw
/935BRuXW23WH9Duia9fNTuiWcHyqi6rMymxVfMqRPTYyZ0erAHAy/gMIuaoP34W
+o/61YYsl7Cr5RFhZot10mcbqfjYp/UYgU0Ypo1tN7Derc8o3Qi3wEHymutX/zLB
3jvU/fSDhxGzQ8qw5yPhCbIU5Pz8qJM4VuD7FnMLKsc6MVsxeMuB+X4PYU8J2hIY
/k/eGGliNX6lancbQTUTJG9BNmeRRmhk9YN0TmC80lgU/QpWsrYYxs+2I5uuQMr2
/DJ0+nXqfnFo7XhPw2Nm9QzGxVVoVZWAQSg90nun73NPDePdXn5XZflF8JTMYL9e
W7VwA/CJWAc0/6Q7Ke8a/64i8mT8P9Edh2ZLViC6qkhYs4JSSBVGpbjPD4sQUXK6
RauKBJLMO9EZ1yk9Y8qpV3zEzDE4yTawCi00w/EUEtNgG/YGYo/ZpJrmcEim9fNn
US8OcF3Fji5AmW3Lidt4s6bDhbUgTNcU3hFTfwm2mvgYOVmKgobwAMc/o2vo7c7N
bMs06B9Kk/Mf5AOAFtkMydJjp+pvoLjF5gaFjBJRIfHDRFQloRsv9a7GmRD6nUec
lkI6uX2DPVJmgMQKQOZIxR7bfQck+TWKl+ZXwJJJYcum4kuLoJ0WbU3hWm90/dyM
Km4NDpTy76UTfIj9yEazo7pvw78AkY2aTPfDAcgHGK2/q1ghP7zwkYHVoqQORTVM
bfyMDBpwF0a4IN1OofcMynud2kQ7QAzaEqNrRv3xQY6jLZJ6cdi6hD/2ZxuA65sI
TsNpXOIdsB4+5V+PZy2xm9osI0SmqQdzLNPtC3jxA7kAbSUSqX+8e6JZ1sNYKDv3
0Uk74dp4lj/6UiVknxl4KFMPCfYAYll3Z2gDSlTWnGPB9/W7S3FBcAqAPBYcuiqJ
EP9lYcm2yXtz0psUqTJM0uSO6ZmGMvdWjVF/IEJ7vA+RdD/SWiyQZnmfG0I0ppba
DcFBul1BZ29ADU9oAEmIGBDVUm7yi89qnU5l/ML2dpJDtBfjNIXUoWgPkhJBMoJW
UoijGmUQm0GqHoebpFvWcnyXoo5F7QX3fdE4DhCxBm9pbzurKR77vah6yu5+NXQ7
V0WX7KdfWzaM2GYyAQy4zKbO5kuX7A5liJV8BvcIavmyyc2eb4Qj68Rg2E0ySHGZ
0od1vtlv1EqdNe4n2A3sTjPspwlrdmQ3drBS5rDWhDbTu8JVGdNBItPFRvkL/eLm
IsxtthDEVjaMKEwklJd9yv4CDpYexfnJHWMlR0nRKqTAzmoo/3gZl8bLYUlax8VB
woP+1U6p0cK4dIQEzpL8EBkzarRjlLfVUgM+9V0NgYXx2shzWc/Sp4zjgD8WurPi
xTii5u9qmJiUOuJOJ2wH0JHCNTvy/1Pg9TOcb0BkMheaQ6L0yMZDBonGSiewpBus
V56yCCQck5NV7WggJ4Vl9EyVsWCMfF2F9hezET7uW7iClLqFUVgg12Q+g2/nFRys
cnmML7n+mbW0k+mAlXvhShYF1u8TzAF7lJdWxR/hodLoK4URJaSLqdbQ9gz1pq99
UZfHtBx0ZB6kMTgiZgGxz3+GTCZ8vd+Zur88sEmRWL+GZdy/EPj5IAktaDN5WU+m
PYaflu8Vg3SX5hk58MI9Q9oSK+Bm/56pTyU7jjg4PJgxfCT/hGURXYklg/n3WRcj
FmP99KiN8YxaQvN3GBuXFeOxQqTtl1pbvYxZmwEUHXBp+Er7xEmnWHC/TbUDWQJT
SK/7EIghbVRDSsCofq6e4AG2ugtVnZy2EGZQ3DAP9c0Ql2hhfHXH4JfEu0h487QR
YbCwwx2q0XQYA3j9pkt8l1pJ/tg/Qxa6UhgYqYCgbjbxh3utm4vMXLrl3wTtpiN1
LXNLOYUbzIFhZC55QixDXb4p3vG/BHm1+L8A+/c3wjJDSsF1Ko2HltUZWGR0gSi3
UY4xfDJA2UYphMu7/1TMth1ry4ic7S9qfdzNTfOp/VGBFX/yAAj80tF493RDyRQK
HO5EpePjrWZAHey3vmGyx3B0gB7bo4+4jnAR/Vxxxh+tzVtlnQn8v+lAAjDiFU+O
u5xhTZYDYIowRl+BBI72eJ1XJPXO4rJVKh1NGowV4vuQuZYEWNB7piGTWPU+SSvK
H0uiz6oFFoNJU7p8vqkMbTmFBswAfspz8kYmYmDYgK7hEeaaF3VNexxD9mxdQaT1
4lRo9nCW1dqhC1toQkQD+Aj/HfmsP2YiI2Kzs8WAUWPA6xns8oc7UfvJZeOk3E5v
AUozbzc+qTQDckVofcy6wNHyHSudAkuiWIP2OhKhhR9p5+tPoGgmyV8q00g6OHVE
H3X4qhWVfToYCE1yIHIOBbcyU4Jtm4wpOUtbSaBZWlqusBRWZZ5Xf1JwHmaF/zcx
R0Ipi2gYQOws4kLClZXAjAFkyiXKU76Qz2J/cAzfVS4HYl3EMdF2nJQ+7cNxDDZJ
j1QiTERM92qy1qMBHlGrxNXGmS5bBgsP7X0IsQ8aUKJetAP15nawXEc+o2rG5KzZ
Sz4RZLzGi8j+Y5hsvoUfleldhEclIW/xRrJpdgfqq5ihJkkgxKIEIh5oH0/8gEx8
p07w0OuIcOzIvaAJ/rp23anvh7RqYYJmgri98wFMPzLbHSjKYV9uqYRV63o6QUZp
jOg/yjF090KsI7jYnfUMPMIxtLmokLxkoF5jlv3R8dwXqhltmWrmZHM99h2o8/Mi
JcfVbf6cRZaXjNumu9QcxFyOUtv5Oj1NZBKHXVi5Q+eCf5JPMHPRLgUyJF8Z/diZ
CpHKQtqzkVc2gB+a18DhN5vL1M7dcUHJtIiD8QJ9u8l61oQPJFLI1XDbFPxhWzF8
HvtYjC4Af71+LO65X44ohruagcz3AjATlM5FU1o/30F7dE+WsqyyoglnwCRFLtCh
0fyYRdDezTwjwUxwYygiMWNRcfDeVU2LQgb+1q86ILKW6aMHFOmSlrmWomTFs4W4
K5Uwmh4/DBt2clSXEQgAr4UwXqahJNT1LhLny3U+c2oU8e2HRejYJhby57L7l3P2
rJ8I7fy9AXSJQy6LjZUpWjcyq9NIn5ouDXKLG6WrxZCRl0gswiKpQLrKC+fscx4/
1ZKS2J1ihmVEgmSmNuxooQzx8mi9rq2eA/PCuhLvWLc52KBSw4fWtAe3EEpOzhF5
9FShwKSX3/2YMsRw8MTYVXL4G4SD2Th2mAekP6Wb5lFyyWoJLsf6K1oa0nxPx26u
2kyw1KIOe+ksGmLhcN2zbGJVkU96edUtSdXZTan5kwe3wkKlDq3qqkZOzd4cviwv
UQUoHYpUmNV+EPx9eVHditwPhYXos3kSdSOgpeGoD2E/mhsMLIrsRanAfIe+MW3D
E622owIH+AZyM3ECcWRuE2+DwgXhsrYJcK1JsFDoGjZZtzddg5CJfBly8j49FJBJ
ZsMObsjyBj8otpkeWmo8Kbh8+0AqO1pH26bx6zGT3IaPq+jQVtTnY8ZNrTX2El5q
G3Ehq9yw1tc6VSMYyXV2+dY8GwkUEHbVu7qAz4vBS74whuErQeGdM84rDIuNpSKL
P6jca2cWCguiqBIgCn8pnDUQmgg4daSu84sZyB2Ps39h3X250ABYahuE7EVgm9M8
RFuGJJlBLxXojq2p00u+Vb4dtT5JGOht2zHN6ubOSMWUOz4a2sdMwkTlEgmcy/RT
NQ7yr1z+Agv1bFCyBvEVoPlSTl1ui2yxzp2/JJs10cIzJLXNPMTHxGtWlUBQ0B9A
7aNFZAUaiFEB5gjJjNgap0L5/VHGW0XUi47YaVka6mzhssH4oRf7WX64SYszFcoO
qXpTscD8kRuOlNfNpHpMuSzUjva7sqZZftuybXNj3BB/wRyGIvln6pPH2SIU+XMq
bK1mPChFi4tWg9k4w7BCFILZV9axRJs9gBYDoz57Ucv1Qh1GF70E8vOC0Be/5t8q
8N/2US5m9EO+ZJ+iZ+2BBc04xPSXR+shp8KsTLNp0Q6fdq/GF5IlXtILiUWrF54X
6IIbAAjUhfN8DK/5VEtPnPLHMoVgAkqozx2NAzWGx1VnY5GzWT5QESATPNFo5I7j
kcmKS1E2P2hYJD3TbicTuMkQHFsDNYbqJNYJlsrD8oAS2OjV2bqNKEkgqnLDGWl6
wMUok9HgOFmnauMOmbB9GThyGWrKK1KDzHGyW6eXhXlwSgTDOTzxmsOw+B8wcoMA
LnOMnAppiiPVBr7BRpuRIgJyNPyzbzw0308rUxBArF+63NaglrLqefeoWEn1Q+Y3
2IEtRfGJi+/fKBDeixo8Du8LtG5db86/9YtjBgJrxG8gGzSGIbtTn9bFKeF7aWXB
LKzI599PsPViDmtwlyj6vOGlKFAktQVj2NRnvkiwzO5GXidMDoxbenzbtdhEf+1u
QudqB4Bex4svPuKDIC6UXD1VxJXSOx+lmu02mJC9yNR/flVzbSXh9GoJLtCLfQub
GYY+1KH///EU77fGh1Sw/DO5HfsvDwkU31SewPjYYr8NJgAdcUJms8+HFzUIQenb
ACIq5mrt58B68kFZm2OdtU/azLo7wCkRH2Dzgw7XVsLkNJZJBh50NGuD3Ud1eiBc
DGOMU7o3FzeZBx1neH8v9L33u7JzTqDnWdWMHuIlnXOoPkYx3Q30L/W8IbPPFY+g
H4hbKunY4wgbwkeEtFXaOLlgM3+UxukpBIoP4xW6xxRN68f3e9hSsOhpD5GqLEY9
gAbNn5q/IijWEhdt9trWKp1rN67geziYHnJtKq8uzJ1x1U9sCj66VmfkUV+TJlgU
BcbfM+lJtshSP4kJJhyeykcVtofKpK6SetZqStb4cp1WwOTB8eqdXwwJ2Z/lwF5F
ZbK39kZ1tNTPhFnR0ROdHLb796zd3JfICQh4Z2ILnU7QmCU+BiX2yiHtsP/rzgSX
y+5xl8EXgUbWSJxgBtn7Olf+8hHNvkdrmDMQVmc3RZfnwxB1NM8BVGa8glsqAZMj
XOiZ+e5BN6WYjq2x49ItCAq475xSKjJUYwk6nhV2B7lDwGLHsriBhVBcJ7sxJs2H
zMn0SF3sQiZ8h6oY9a4B/GI+b1ZcFiHt3PJHXLc7g4vVLfOmHlex8pJxR9khskU/
7Fue3LmARMvgesmkTCM7RWu9xotor7aZ7bGcChEcqpo1qyVVWNG7WVpX2Sj51VdV
dSNh87FORSLs4X/TGFSHr7Lpq4Gy3u/Ce9gg3B6/l7MPQhpweyRt0AZkZwmlSNVr
qZQxWh7QeNZ9CIDMsqVbb17UyEee6UupgxS6pDbtYJJ1EJNi24hLbU9gFVG1m0gC
lFBk/DtF7ALB03o71V5lJl8NgpBpOBdF/EJiy1f5fQ6wyLyKr+QLJZ9XgyffL1+N
8RvDq/dZl7iHAxnCa+r7lE27YdqW+ZhYmomqjmmF2dnu6ysJ2xyR6Du4/8KXihca
djk5MIDnlKjJLbYGha6V66mJc2VbYboZaDbiDof6TiToNutlyEW3tJ/JEVEjGY/s
RT0UuCO1K8sru21rEX/+W9PYodf+bBIYrbjZURQEvICYB+qA9ERKK/VeWc/lo1Jn
YPyrtmVhatx8QyGn6Ol4rO62G7XeE/jGThwYCrVfHPL8Jo5w+8/bLAAw0sIJ+UzI
KrWtmsDJLc6GDRkmVW3wnJIjRGJ+QfaCj5JCPTeyPqyRTJsiZbdYGq6THxKhYLTO
i/2hEQJa6MW7VA5WlXzmI4b0uZfs04mflcAqC628vGZ/tsbS7XywkW06nz2+f3oS
tQlU2mWuwe9dSYjvipLHnEclGOvrakasXxAsgOIYTPteSlGq6DZ/lsD+A9Lk8HWB
tnE4RSjiZHfrELk+xt+E8tl85L4TFP9H+trI75W07IoLTvMV8ORGzo4m8mpF6tBi
b0REv0f489v0zfAGh+Ntqnyrgb2wWIlx0B8hatMuyvrwnVKt9m0dVC//1ES2MWDq
31JWRYItDldzokq2O/PxWfzRp0wz/+VT1h20wNX1bxMZG2zyKaqlxFpL4/sAeLJx
8WCu6EstrKhN/5TrRJ2gbV2zCnQNwhqXY00stTO+s4kcsWEJ6AscvUHVHOuszDB7
L67nivL/DRxJcSNqkeHoJtT0QMFzjs+Qii0Wk0ojfYyJjRbMiXp6dgTORbBUHQYs
jJEG+TP8tdK61VDllYVSRnNTI7dBNjEdSOB1xRB92QqeujZTbwmVYzYEhVGvcqqv
FU0UdReLbZVMqpExFp2Klu4uXLR4gkNEfU/CI4dVSJTbu1ozovKta+66Om7krdy4
Ton+er76votnqvw5cDwkoeFnv+lDP5WylicGDNyNiFnk29nnCnOiDYNtU54es3d/
VU/nYXZgi8+d4bKUo+/9TmJhVga44b2rvaQchgSN2IvYdpg4QTimD37ujvhU1Q93
C93JS2+tr3MApBup1WjPQ3Ks80zYKMBVIXXlcnV2T/PHAW45UsUBiTewpQXwVgmV
xsr6Xq2YNcEEp69hSV6IruUbVs5MzasFr70QSwF9OSVQiJacRckXKUbwTMyCcerm
fSAzpDlLLyD8F7ZKB9/wH1vnVV/wjJyt++agakMqqsQ5FktsrXl/fGzel2hvvdtk
mtXFOZEolBqAu2BDAwigerO6X373zmz12i+hGdDcK8pFu5J60jwLysSkLhdbXCxK
82uuMGXx3r4thwbCo+lBAPl/9yfkjr6OuKA/CqPYOuZTweYKTVsSyLkPL/g+4aLo
eQI5aAEg3nQoNlk8v5gLJ2I9JdpOuqB8B5ll+Zrp32T8meftIr9WQX22Sc2wui16
TN+CLI5MtMYB+CM4rC9K5ipCUTPOSbVTZx9C/371JwAKmLhKCPIOX1Y1BET71HM6
Tu9C647DNXs8bQOugXCm5pM8sT08jSSgVl/0JFiQzDPOfPQhYR38VOjDXDayjHyZ
jxoJknlgcZuJNcmkK1gDmfh6UZQA1/fLbDD9OnPmym98TnKStdG7FnT4nAyu6pmX
mBCOPByNH6YQPgbOsqw//e+g926rQuNCpwgYm82DNe+wxiXQBU7DT0+JgldFIjuC
yCnMng1yMqBGyTMQ6AxnWgOLp/5fJIOnQHlk+xM6Zv3Cadbzn2zaJ+xxgXi2QzeS
qJOPpag6FBiMo8QJXb9JBLlLIxlqMISX8+e85bL11/XcBj/fZTPZi75TsG4tEFer
9OI31o8gou7AuXZ6hyPpcNEJfF0qmwMuaRTCBXNI73V1TfHA3ggN/DP0qkialQHq
UJ7v7xg1NNx88ftn3RMWOZysZX3EK4QbHFbVtNpGnrznJZeGEnk8Al9aDa0Z8qKL
kTETWkprjD2k+nk6G8EmnKtXh6/5SvvoDg8ZSBxdSIMQUDrDerp+ulwV0JvaZa+6
8QI1sCsVtxvQnthH+fcrJ6+aZCqAOewvEwg55wIEa5Gh3xsU0lc3Rz621ulyVbsu
tB/0p3EtBcwSwFDXoOTVZw2t/EGZ7PmZ4cJeDvOlcLGz/0RgHCCuEfK4/rv8SlzW
q+WLvowraSiayO6/JK9snUMj8CyOeB/Csq1zCKOZGMRBRXN00umxCUPlQB/pWGUi
9fXq1KcJ/DThzd3rU4F630iBw3Z9Qcs8Igvf5Rp2WTmNoLKe8zh29YJdgzU2sgO9
fkUgq+BioxxaYf5kX2OoIumzvTODKI+LevKGXAbsdAz23KByQmzFk0b1Mt0FAqFC
qaxAmxuy/l+Ub0c/POWGgCJ7PuzFoMtyfDEKpqpdCyEyZGKIUF6oCDfSFc1p5UlB
oWGlhfaJf+fHrvKxhsewAcgNL7hxVRN0KxmUsCi3e10mNyPtr5ytf3DjIdei5WEl
tqPpxN5anjh1Vj0JxOsGP4Z0vFVFF59LPCKJU+TL2xca2mEfZZxG3gODvs4iuNv8
nKcUfUjQ69cNLPyCULVxBOAFy40bhE+qX1rxIdqo+kmXvF6Clc1HY8pXiIICJ0KP
WDbkaLa00+RxBfIfOfF0Jqd99m2ZGEPbQ+KsXxsVwgHN8cy6wQ2WQw0cRelwKzn2
MSZAkmxM5kx8MQr0OwNIAyaRtOqlkMeZUZFuIYpjTYb0H5+crSkVKMQf4ZzUv4nF
2MlKaV2e1GCZ0p2eowky3Rnuu0kKjh+ILf1YFVUyOgaCeZj54O2GrHafHhC7wh9g
fVkskwrdYOK4KT63q5lzzbuzA/1WdVuxjsmCBPbqZ2B8mkmUtR0EzXK4zOfAFQ8D
JKLjNLDwoxBJg2BNy9mEAk92TbHOc9WBbrw62NZ/i19u0zNJPA9R+yW5MP9E+taL
pc8SQ8xI1V+Ij2kQaFR2hqxJKWeQJaTrq9OrXdxEXjNjlbF0k80dlZ/sdznAhn9g
5HlgovOLg7WEjzVPPwSg7W+XXZrxe78qY0MzAP8/CqpcF6eHQTAO7thpOENHBS1/
P43daJ24F9ZXiqwn25NtSQBQchtcTZFx2dt4badEaIB+mK0Pm9f9428Ht+/C1x9H
TcS6JsdCMzQ3naVO8ZJpYYk911ivLunjOEakfzJ405Z4PA8/cI5UVZYBmNLErsxd
uP/WpxwFtkzzfJiAIKBZq69We5a3z0WBhJtrS5SyTHeainkO2gZBJODYyX7iqaG4
hGCqubmQMimTCzcDo9tJQ8D+S1Hls7OtNQpf+ETCT4I+leR/dc8MU1GkI9XjxERK
8KAIGUNUvLXFOjpM0lAg7Gm+iwOEws9+8fW0P8JxnhAM+SZnyo6zvL1NH/cbbBhH
xtewuP35j2CFGGMvhAtfoDZoCQlmSGK15iACAbwzJX1StZ/dQiUDF+BU2MSQoBrg
l2TfC5cUJYvyps3A5FAfdlnGEDfZfXfRRteKytc9B7jl+H9260IuqElTvGFrbNjP
QI9uUDztmUUc7R/msUO4p0nd2eiDR6VcW7tYsQ5KfrbhIPGWmzNML8oZqaYW7B2D
M7Pdj4/spCzWS/JfGjzcznc9q61qGTbiVX0cIGeEQ3NsR09WOWvFJfgWH7KEa0iN
JEFg51rqqGtRiMNru4i7n3zjmlKK0o95Oe7pbAaV4XlhZOJL2aPyOMVIIJNnbKMK
bV7lkmXuI8RAijvSfss0eO2nx7n/KVdkVSteC1n3URU7JOlkD59G3D4qFkTG1QH5
p8/xaAFwRWLlan9WUN9y4KQ5ku+Ko4zJDS0bLsEo7DybAN2GDx5nV1d0EjPULGiA
Fe1WvISuTrAVnUvp7mMVzB6D6Xw1h9iGsR1emWZdXq2BPB8hApr0hNp93KM+5pEE
RPm5gE9KdRCD0FC+YBITsiD19Aze5jilIFi0w2rzujyxhCAgSb4ZXVi/5OdXm8Fp
HFkorhdIsWcnII/FxyBwS8dk8u0X5JpTPRxscSM5cp3TaF4cvwtvPEl4CRuEhilI
jB1rv/NnSRemL4hUU7jC9Z7OaRxkZnvPiopmsHPpdzKtpHoqaycAGqj6Xxac1s1f
uDZTISrO3GfOxv7qRrJHu9ktJZOS1QZYVfwAWAD4JiLMAEzj3OKU5SQltQn68v10
drSW8IzHyP9R8nzaZYINUroOkU9ztyYun3xeryHp2BevG+gC2WzuyWwyqo8YyWvf
9maeyZq+taU/+V2cE5VINH/x0+VijSrP5BUJ+AEUY5mWZBoiTehT0YUOHnTZnJay
NVnNsMosyGRVQFoc5TcffabIO0s9HrlEUgmxnGs2+23pu47+i4tqjuerqSHSzr9L
2H5LvHK8SGq7DqW5vO4BHTViZand6xDeNlaTOvbRi9cBVk9RhNAzb0UfuYQWPhvd
gSwxk9hAB3i8tSIh2nPph8WoGl7zMqLaOxkhsOODkFseZE1v4cQGrZYUm65sv9Lb
Dnfdcrg9GwnH7lepGHPlvNaMYsY3XhqO7GnxND/dSVcAaKl3PMZ9HktCTLCSw4Wc
/miQGAvnSmQ/TwW+71hPxd6S50yPAi3e48p9eoeYrjMZhgaukLznOW9GunWBcYEs
R2SWHb4cRWGn+rhvZnBoaj8DPqe5kYDQ1zEPhEpY4X7bJiTQg675aBrAmLAoyXe7
mSm0lNNC8UgAT3OFokPTYCUctHYol8PFTbDPwwQ9xx9jm1P9c5Ffil9aGFhZ5ZLL
FTj5aZ9Bi2Foqdn02enAV6J92XFnHotLWKeFvlbUXQhLVdHzCSpm7VQQt3gzx29R
HibFlc26cgA2pykUIPL8icch0Nw7OBB3GVE0I5sdPFWKdZbYjAYILNfMC0qXQT2o
fatRq//2fwyku4qqnED0PBDJM2CjmSnCvmlx4pCgVdVWN1+ug6M8hKczi2hwpFrD
WCyF6IQmcFIaG99Gcl87C3uZc8N2dfQE9mpBO4H0PejaQ6iP5TMBMSXZjpxWYhfz
ua7Wu/GQ52fCst2N6DXNKXM2OQzGf1MESLn/RTHOgVwzLmT+S7fhJlZwdCD+XaMw
YH+lbc+44nWDvi0QEq6FrmhG7RjmsPGULjMGFvMqlEVpGzQOHhijrLKIJMe+1lL/
97DQbOx2mLRSqaRewUyf/mJf4HejS5L8snB7YQjRul3dU67EKqzUFPq3dqtJH3Gw
xA9rg9xLo4/qmFnReBAGFzf5rB5SFEtIVMq+3ELDJteC/i3t8ecvf05KAD73pirh
Ix2hMru/fTifLT6nKcTHwfFrYtkyoDiTLqD4gT+ZWm2gkfLSDrv3f3jKDGz0GERR
5tTuYVAzpubDBFBe+MNmlTXkdI/QSZm2eYCfKwHz9W9ltahG5eJ3YyXSz6PqEfLe
3pCDTQXfnvkqNyl80Z54NxIZ6zqrpdaiQGjXU2s1fure0BTWE/Kqotc0lueLI2T5
FOgi4bA3ptSWLuXbS+DXRtF94lZK2IvPaLW+/r5JLcjNQqBCaxf3JS2/PGEGmejH
g2RficBih4xa3oGwXpW+AtiJt73k23Fbn80omWD1lco72UnFBtye7L03tgzcOKXR
jFGYjq7A+SrZUDXjOdDEGFC7j76ZrP1NnKJGBLAwYkX6mSdFL62ThUO8T9K8GWRS
laM4gb9pwa4JX0J0e9A6C/WlSgMSFxNPrMtbLG2hFQaRK1ERLKdTNJS7vFha60VD
1SWwwbwgFNQ1FrOSI6cl3EFuPEe0VzSA4VPElCxvIc6UnGG9pIj1k23cIuKmttsu
FGJaEnCyOMPxXb/mvjOyW1EC4U3WRDKA2/Z+FvUxKckq0SbIve0sV4OZYz3R/SLd
BTBy0OZLsSOouenJrvxHla+fFvUvDHIaNh9MtigKaEesVrhI9rsozli/lBiU8+1D
+GJH6qFuSsET+lcq2v8MWi0USZEojfY1l94q/DsasOSXCi2jRo4qp1AiLYteVpnY
tVsukXVjisaDct29Eqx6SQIe3D9S5+GPbmQQ4MnX/ZB3pDMdlbT6WAQiW4ul0MJ7
ZGWvD4Tg3mDoUPrpPSKqp9wvNMjG4dz9q18S7JbPULP3p2jjRdc46ygqQrUSXjFM
aS5qdnmgQlk3QKxnHt5Bqe7xUW5cw3TBF+6mJ0gdv1heKTf6uPmY6XJTzLpqA6o/
ZE3sMlx1hxVxyepqfJnYesSpJdkZ8WW+mjscPpfjBkw1SOSaB61HJBF2jKpk6BBs
ltlpXZvbd6deowQtcuar3/r0BxA//n+n9HDAAyvj+o4ipj970wlb/u4sVwnn3ccS
WLWMR4chxULkeaYwlvMcjtfpYHDLXKukZYBgIB6ABADagVxxZF9T3QAxfJENp3t+
+ja9LbsAyLmf7ZANoj1oZhXPRZv4mSFEDcwj3BtRRf3P4FZThLIX0glsR+h7maCm
GInLsjUCTQ2uIn8ETcnXqTDofWQtbRWXu3TySqFb+tPzV5xO0B4Fg9gmaTHflaHW
xH9WFKSofCVxlBR7mFMCIGzAqagkXLcEolPHmpToFKPunQr2n43yqOKnxK8H06Cr
9cTUkE8k1XplcZpDTOTCSjktE5pJrkWPKHwSKBFBcndVnrjXCucGNBeKZlUP6h6f
wWdO1DTs+Y+x43uQYGJvAlto8a+DvC3ejCuUpqHfRKav4La41hgJvl+qVH6TeYp9
zk+c9WYnCWHmsNuVco64O5c8t0qD3BwXW1QBB24E0/gbJxdUUWP+sUciKippkNvt
kd1H1Fk2QtAzoDs9WKhBT8xH4LAWHVvTCvuJGIbOD5bYzhQfhA1dpTjzjpiHSUp4
Xo1u4HzqtGcm2YyIDI5pNmh5/d3ev7kvUdSWNHL+NQXPy4CgU6oEuRR5MLBL+0WQ
TvueO+A47lbFX9NJ5scPBU5v0llstJ5FO2iEdWOvpwFD8X0ff07DNTP+CorTi21i
wnzJD42cEL1d0cS7jEpW5tHSNrNp1Hsqkwy8jtACzdbXWbs3OgSaOME4JD+4zCW7
y6GD9Nv9/7fZjvdrZNiW7jhDM5c6gaBNYno5J4M8l5vU1KVAFxf0Uloli/VAgMs+
JOQRt7X0ORMADvow37GyNT5hAVLvA4XNEV/I/wgGg/bEu0zIu76Fs64n7JelC8Ys
q2gMXgGTun0/DomIfc/agmMQ8G+NCy9Je59mYwvmd4lBXG5D1vOgoc41mTUmO9pN
4Ic2+Jl1183LS02f2CbFjs32NvnaEFDst4ao5wmAyRhtn6kjJgV7ZxSuxKZwZH6D
r+Wjk+lWE/JPkoydjjsow50JffnXCJmUc9L2o8asri21jDWZz49UOEOE/yJoRxn5
LfvKkEYPXK+TuM6H3rz/V0JvRkgOwjC19UO/V+4AuhwigDVGCGUMRSRGGn+hYsDv
kMR2u6+zWNsvfZ+f3wjL//0IupUpu9ZVS8cKcY59CxXTTKF8dohiIE4jTNd38/q9
rPuNvuJ84YNm6LP3itNyu7z8oKcOmTGZJIKRRCXhPUiZMikn3CaaZzsVdzzmaI8z
fIRfI2evd0kpbJTqE8Vu8rXNSnnYubG0EDdYOIg8guBbofTtHzOU//KkXg5XxWqQ
t8Cm6hmvnMviVR43Mf8IHM5rXTRhELf2teAF0E6aIeAImzXAEpOYJzO4L1dSJ9qK
ZYZlcakkql/qnoBS4ejXIb+TtI9Fma7IfyUoU44eR0UDvQDQosRr8kSI/4HtOftO
T7zhTTUdlOU+Rz0mV5XEYq6+iFrWfsTKOmJ+jO7VboaCCSmDFfyKwiRNu3PFM9qM
Pb0FGOm8Y2Dd/SdDALkQW3u4vt5pKoiWDHUvJYaSXFz/2nW2BFyrAFDm4Zqlb55z
JzQu7pjtdAEhOYuOINL2o8M+LerCtEgginKATwoP8qOiXyhW5xn2r7/jy6PC8RFw
lJClLC2HWEqP2lWUtGxZhplJmh3zruqhuz+1zLakdisI7kT59drg4Z3ytGmwjStB
lu7ie+jwPcKD74K9xFV7MiGRCT7ZbjO0IguAJlQMcFlgUa99lLjdXwxxCTt9Tfbq
mANclsmLWpK3NbGsCqnkzRawqUiswJicFKGLbD8zaphG50kdA2+kiJ7sAeKnSQG9
MvgjsP7phj6JgJj2eQuNnPh/J2X9mk/M28couDxB4n4PGVHDuHd4/H+R2apVoLc5
rPvG4NBucU69CNHgBsZDjkB6nRYTMOOg5DBA4YpmzPtVQqPs952wCB3zYfNOe7y5
Sn70r/f+2VLbeuu1pb8zz5uVtzm188e55BPLWc4LbFTYF4WaFi3SajPZpPRUGrgK
My8gMGXzKfomuLx4en+uVLikNsjMS0g1CkVd+SiOGmSGx/UNsiUX5EvHXwB2Xoxz
rGAbX1bu45HHsfceLz9qZd4Whwpx9mti5rWeTOhzZcHabFlu0G4Magrj7G6udLZj
8bTPP0wDQ4RuO6wBX2oJIFecC97GHRSLsu9gWg2YGEB+gpHpWj7uKEhhU/WB0A0n
WpybiSw7hvPau05j/H7byF9n78HP2IrNIcW+/ta9LCIMIcjLdkLwWRoDZ0spC052
1bViX9nduMvS87WbZz1jKnZES9OaikFifvLdMs2ErWb6SY4Er03xqmdHTv67r2PO
oLdD+UDpdlrpXHVh1v6PLLlz1fesXg5dR6W+DSL18tqfRbwIQ1k8zOJBNZQyBfGx
Bhdd8PFzALleVlg2Pc52h9ZXEd/aGD10YpxG/zw8Q9Zt2NyJyhFG8lU9avj5WVao
xXLrBXLHOp1ZCoIUe68953AZUy2MeiGVGY8FheyV3xgIJRFhWG0Ih7C8bfVr1p3z
GOYB0KPlLQ+V1QppmhM5FNqd3rvJpH1qMx6DwtGgFlyhXyKABFZ6UJ2bHkvuN6ky
AqFfhrw7aaMmhAS5Xu+9mTLJRk5gvAI9y40ECT7Imgl1zjdk04M5B8de2mwK72lK
tASfvGoXeM26xRVYBid/b1h+Y/ncPBnxFOCwVg2gYPPuxLyjIgDj6LGPLm3fPWGU
sojXRrNuo4qa/fIS1tDIYFugMl1eDqXNWoyw/2+mmanE6Jk5W5HC3ZdKP1DmPyBg
r9eypoIgsr5iSBcrbUjxc0ygg5nEuomYQ4QNCdj9qUEYSPypdX2Q2bOZzuaA1+Tr
+l99jvihGQNW8DAgPpcAJjFYuQjDiPGTakl108PDT84hzqtvNFvXXbyV1zAfWOEk
7gtfc/yPjomKXEb2kmlG/JHKMW7Cm/njf4RStzrb5kKoBQE1RNgYW2iBl3KSwdjt
V99fXCt0K+IW5qdgIDNNFyO4T4kH8ptdG05nl2wxuVdIK+RvaISMcMTkeuSbKTTP
hXrIeHUDRq/j9LhmZj4xaEDGVNRbXCwm7y576hjTGDDgxV3eRzjKYGoVchZzaHef
0qAnAPeciZnB7N3nqqSorEP2xIJN3P7QWEwmtpatWyLwOrIB+RLquWuAjJIkEy+i
EDEZ7pVPjKQS/YeV4bN2MiGyPFqbCHLouZ0LWX4mxEWQ82czbguL1HrsL4X1PRtV
64l0dkybjsfEpSPAsnFK5NwwUeIo1/CpT0GyChfQ6OhIJ48zVIxjdxlzhCDGYj6X
4ka8EFgXwzj3VIZgmA4c/aV/xLxx2IIr1Ud0admBzwhE9kI0JEUkl5sy1wqdDwHv
EFNl4qV8ifZebQfX1+40acIp9kK35IZCLQRtY7s03X/0Q+GrI+3r9rE2W26yVXCp
cI8n0v2Tc8vo5L/NFBbruGmCwwnmJ0oWYBKKIogd9WvVNGqDU1785hXMETkbWlYN
5/C83hU5N4p04cOueGIsTpPufyi1Rr4WEBUg+9gixxNw2/Fb6W6S56TcTSdMUjrR
upmDaYvr05cKyndLSUFCzBFNud5Ar5zxQRMv2qeYByFjgd3omzsAK1YTGYoU/gQp
FpN3oLP+uhg8GyHbzWNtBT3GJJIjDFwhl4YUhqcLL0j6pPHBUF7hwUXvj8ncmQwo
39pr57ZoJwn76KCrvUWkog2EhYTpptIYC4yp4X2r7t3fuVpFZeFaMMwpdzZl6oKZ
JdvgMuwuD8o/K1v+x4KHESLPw9t4UYGnwcQ0geDfGAwa4Sxzdu7phrfrkjouiQXS
o5KsIDCA8Rv/ekGkcuPOghd2Q/unr8THEE0duCCseEgXxxCEeeIuykPF3sZo0bh8
zGek7DcqyNOFa5NdUY3lCz5jhVGwGqB2L7HSdLeeEJjb/O7lTGLxG1XpCGC38iqg
w0MBdMWk1wWevR15skyEmlViv/JMzHz92IrS2Qdmh4ImyRYUJKTrj888I+2SrI5I
1meBTVG7nfZ/Tqh5jIxrbbu/vmxIWnuAEABUY+x1JqCnifnqZ1yMdDk/fypKkYDH
XLQP9GgWpVzX189fa1Bx6EAl9YrxVo2BIwHqmSHcoDG05h9JBbx2ZTpvW94oh+0r
f/SgvWaT+12ZlG/RLKC5GPpjGPgedQ7z0KdckkWW1WM3kkiAhiJsDVvnTPQwe4wI
9OurUAEDE8TqeQOd7G7detyHRCF4AwMyBHX+Fv86WqL3RshUrjAYhHi0klUkK/be
ScttweYYG0uqBHinJkzyaTHKgOcERPe+bZGhn4Irpf/1Fm3u8iWc8H1+qs1BJ+wC
dTx/l7F+YSHZFadKgS1kcWGhdqcvWm8dAFjmIbP+tEV3ebHxWRUVDBUS8ppowsDG
TpuQtjtcWVZhxu+pcwt/3nXJAwqFaFbGn1OlyyLusQPZ8yjqZU3h/2CDq6eG5Sq+
rDcD4iV/zP3BnYrOsijYb73s5LW+ibs/1HZmTA5xBL13vmJWY5BHSd388Lzmhm5v
CQwTihyuPRM8womTWNsdC2etRiaQBJv6G7Cc3AWO1avSUzyEaTyXophCIt1IIkoG
JImQ+793xAYDxZRpdjDTdkUkUVRbhxCqOt+YGMGIT5Mo8j0y4vAe1o07EY4ifsPd
LMsBWGz3oqwnZ5v3DkPZl9wLDkRtw3X6U4ess/P+b65S/PKpfMLVr/i0KlTJta5I
84H8kxcvEIlO7Ffn8o3D30GxCVu8f7vpoL9KuZQrM19uAk1KkRo7t2zf/CcInC6X
gdJEBAq+NqyvA1bCrLHjhB0hHVzxcUEku4zyvvmKhYqiRxqSauoa7ns2DgwnVXJa
Q+uiVAXWJ9h3Jf2dHhrqV8y/ymhWse9fHmfpkF6hqVNcVYqj0dI6IvgQ56/6dWN5
IsCK4tBe2jnm7BsnLV/gyfPVt5XWs+xOjZb1aBfJ3iEtr/4ZsovT6cizxl4XexDW
WCe1osCTBprXm1MOr4bOHjlySChP/Ae4cZx7Gx9pECKwUobCwARwuAGT9i0pLHGf
eFG2xnUuFp0KvPe1m42yYOw/YsH6okXB03DWE6sXMCX7219/oxkL0mh//YMrRnHl
Yqzo2B07qhml5eJybOaA5y7uBOnHJZFrf69mPLiSGW/UlOKkOfKuWh4RG9HVmk0K
U3JVkgKynFLeg9b7aUEDhwGRKpz5Wb5hR2BTTmImpCM7rhqCXjJ97vhVqddm26Dz
fLBJOYHv8EH4t3+Nd61xd4hMUxZNKX79h1bAvOilPrcQqKhVTByaH7Kr92kodwW5
v2TPvYLQnbwPMuuZ0u+KzSEGt3+9LKVnkddjTzx7kAF/WPKiVTZgpw4XpNeK7mDi
ZA0uW66XP1R8vU+HgBVgyGDhYzYTt5l/2PkMwtWn3w6KwGX5yhJzqwLboQVKtKjj
6NimXyMB/0yFA6FlUl+dRc7d39PSfa0O3vYdsOjI4a7tMaeyCqgA0A1I2CfdKYaQ
m8bI3DarfQOaWSpLSVwg6TA1EkfR1OVOrGiXnUvhMcDRVdM2mJUT5qQrRaADr5x5
lMB6YxnSOJ62xFa2lCJ1oC6XYv2QwkdkVVWeMSj2z4fdJdZpIvh6UbqRCFPHXQww
MEFT8BfFtEJnSRe1IwHSvWJP7lOlIshsjXLYrqSps6eQrjGxyjJzkf17LxTyWD14
bARWqeowyIwto4o+e8e1QCfFZxOD03K6FZKXRB3WPigghP1Rdk2WLhNT2h2fVZVk
a7VzjWOuCurJqhWP6R/qngft0CdlDY33skkm1zlkXF7gAOabxCVR5Yb5whkJaRM1
+YPakgDqSWbZSBAbWFyGtBrdfrbZHwBgtm5wku506OXHATVUKXw6IuNEEcwsGsL7
53+DIrIITUkEv8aimmqA5fCpvTSAJw8ml9J6yFyN+wG4wiCbRnZjkW/ibQgKHjmY
sk/ItJfvZAxJ71w5FuKDyf8AWkp8YGHxOitvE/ooW5W/AO0A7NUi9eM/cpFWmxYY
/XgZI5o0liqlqSON6tEvN7FKZAnm86OucFCRbu+FAotckyLQyDMfBg34Cf8vlQEX
r/0bwm7y0m8+vc0UzI1KQ73MODZpEGIjMbnAid9utuYwpdNp04aQHmBv/YNSvHAQ
LcycGqc7ye4pLgqHQL3T9G+F89Cjb0CSVJ0Lu6oTTN7bg40l0Kye5Eg0ksU/lVeb
tA1RJBG0uSlBEHm8ZyAPxJqcDYU9lfHrPTYVxztS5unsgHB+w2VvPD5B/cy+y81D
W8TcMlffhWFCQAJo7AcBxC84yNgPVbO4CXVOvT6jVbrGq0GcN7DQujmliYFQVkbl
Cl2RGBAAnb1eqp/XTu/vN2WJTF1kQH6JsSMsOu4QR1jp5VIr4Qz9bHuC4+Fro3Mx
fFv0w4YN7E44+FifR6zfG34WzrEe4nsI9X+i5oSMCg6Khc3g7XrHRoPj1AT/4JC9
mvL13E3Czhs/D5WaRMBh+gkBXpLOi+MqtQ0Ca0RlJAZqLmgH8xtJ29pTkGf/YuY2
lG/s7L9eAWEjfWIRkwXCeVVFemLO7makmYXDGPUGNtGPQYsjTH/akzObl7oy5Pay
5SSOYVBjPXDwdgXYLzjfi1MOZUl1w7IZ43kugnth+eo4Y5VbvX8LuqW6VbxZLhcS
Awku1EchgMB6fKDyWVlS5OP7kcMLbAb8YDT15rvB0DHFSzJKKtRxHK3xibBoMRAR
KEMiZaNY065QicXudhNcJu7KQwckRmeKotnOZpxangTrIF32n7hanfvLIehwTGet
1cKBfQT3pCFdnx+pJc5Zw6HzLDLXrqxiK54M0GGD6dkDJCqmLeUP7TYYe5EP7cnE
ENkj+5oxa4ltYRJNjQ9wiEbdJcQ+m+sbcaKYE+d8HvP4tB1xAR6OEkR5l/IV5bnN
WMdK1BljltVtRg//mY97ycgtuuElPYK2+asP52p1Fn5WfwGH8BUyTxQGRTnvnHzX
qqvFw8dzekNR1KN5bIkCi4WIdGpCnVFOgjue1Aq5oOy+Y4YzVxjHWXvAjFJRKs3y
mBkuSKWzc4WA7aVmzqLaejtr8x87ma3iRjiYyQw8CTN5b4yghlSbZRXheoxAwYIV
jyRPh5RnBY03bNTogClLXA9HU5we/IQ0MA5mv71sHdPgDKcTqgZfFdROc8oHCjoB
FGX4JkL0uyk/wQlD4ByhTocTULIDonIB+ZC7/21rbsnKfWC5uHdEz5urRhQAzesZ
6TZOOJt3aWFC165ltV+SI4DyVhSZveML8gaAEt4pw7MA+gQX7mD4gM0uwWSYeLG1
8oAZMPaNxExnh5UmPks9BruAX3ja3mf13PKcSfrMD935+GiEJ991S64KAWRgHH/u
1h3cgak7qvXCy7WEPcLQiaHipEeAXaq2eseFztErmWdr8hHSvfUa9814ZcQ5CTOC
XWmC3B+7ZykZKsFMy1OvLceZb7nUJs0mtsNdgK9hB3eJW/CpGRmX1aOlB2OyYsnw
hTZgfp0K9NzHhcNpCk+7vWMQJkYIYlEdTp6q1FsW6VsC7DIIat4XIAdnn54kfD4N
UHV2eDUsOKSZIUw2hnCqRhYjvCGNbZ7NMuXzJqdDI2pe3B2Y7+QLOm/lWOg80Ung
MDvq6IbnnpKkZqxtPy0+RcfD1Po4yn/QEvdql4MWqYzWQxQYTHXQ8ZK+6UVByx3l
RVutkb/GDFxVhNMAcrQPX0P0kvtL9gkSLZSxZXGFXwnG8JvgieVaIASwEZ1e6oyB
OzCk7hA/kFdxgAxpLT3/a4DW+pCukwWrEdu0zz1oLqDUw20IXFTOUjZ3H/VYjuch
xXQNrZxZ4CGoUMw6nyCZ+Q==
`protect END_PROTECTED
