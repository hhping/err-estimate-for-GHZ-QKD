`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oStiEVDT6UCPi+/9uTzgokfvlQkUlUrd2GTmwVeKV40+DeJixJwuqe4UAKPRm2PF
X703lqJLRviIMmJAHXgiBhbX6jIUwqRaNTKcZREhPXoISpWJo0LmirwewcSt7nsQ
YEksMnz5DCjdKOHleENI6/bQV/mM03WNuQajOhcwVV2fMIFj8xQLgEt12N2k/hjn
Cg40UDy7k1YJ0Yr+Xxd31rZzzCp3VMMxHIA4a7OOU+UcVRkF9dLasEOfQMt5VRtp
LM+P2mVNMselRrKj1T/3PLpSzA+jHYI16da3D8go2SmZrNCvxFM1IMMiq9eWqcI/
/AcXDJ0KV8P7rElRAqYt8RtC6dT1tiznUkS7Lv4HKbJX+VgFqqF4/6pIwb6BCmQ5
bz17MFiNhknP0nCo72LDVKs0BiXgkWe4WJ7ufz5ZVWGtVxBPsbxykELJJHKhkIV0
tSy4nKqYaPH83WXxsEvxRFR43VODjNDJA9xMoPgr9XiWtVQLgUnmncQyLXDt0Wjq
lw6hSXq5oYc4ws787zUhS/XNREOypAYpCIeLaXLaytmlZ8vw/jCpE3j7uIsWcoN0
soL93fH4QGdrKs77EyokFOpLXp2xrHlUjLFLk9my/PGl1dMQstJ62GbF8odlazBM
u+SsX85WbtgN25kqNRCFfEsK+fX9KAaA2O3x3jqq5o4WVhLdz2wF/0B9nEKMsXvs
gHuW1E49kMaxndIP8sdsZzzwtU1Icb6j9pUY2a3xpfC0dszRTklcsifnKIxJ3gmb
ewH33vgf/5Sf9Oi46JiEIuKkagdJFh9zoicvEhtwxW8N5COWKQm6isB4oVYQuISD
ruzYgLVJYKlepOC8jLy9TtOet5O9cBZRhXE4o4jfojtH9QAuo3/EvRGJRuc4ihfJ
VtJ2qkuTyK51Rl7Zf53a72veXFzgeVGaN/hpjNloFU6B+wyt22lweUIoxHpX/1zu
s9PpXnxFjkOek9ZMG4OMGu1uCVqFidX10iFOJ43Woivgx+Cg2bLLXsAfr5pNgxKq
VI9m++6PdLcoolDLg0BfYhK2Ea6+cVq1M+q0IPM1/50GABqU25de14t2eTfvuYUN
PLhSHCWyoIHjKqJt/ksvMgxIFXCBldDIbhOTc3Wu9dEISmnv0sQqZ9ZZ1H/CIj9P
6nD6NdrSYpwWvGPbczqANQOn6ZlV5mJ4cd6VIYQ5J4cC+pfH3Fb8k5EVu2ImQkeM
E/QVn7Wm+mgitAUCyXkp0D+zjnOO/6QB05ov7dlhNGF2EqaYRhKdLA+vVXFv5EDO
rD0pQPKdJXk7g29paL0Kpw80aP0SLhklKshwUHcRDphgRzCFYgxOQXsUe+nMLEX4
QL1cn3iG+C8lSyrKDN1TLLhtbwON+RiWpvuXmpKsDOvmmQHJ0Ee7DYuQyqUyf1fm
cG4NmDoeVJfrKVlIoLwDhC7Vns27+Zivi7dLrduI2nIkcLo4dN/Eg7AAEpoN4C4Y
WSsSwnFzRQL3xmsj6csuV2ZpGMfduBKMUsH18IlRaX/X9kOmVbjQGL8h7osolPjp
ZB9KT2ApPnleuIe1hy08eC9qz8sLMLsIadd+uAOcUpKNQ4UczB5cDa+mVs+245jw
+6kDOGKZ5DsfM7atcpkVhOwnDsiMtlkxTem7GNGbHp5DQG6gZNGgsT5ZCOFc2a3F
BhFjZPZHYdnKYuGwNPFVzm3Z3g81uiLMQg61UnBvFHQ/7QCUAD4LqYAmopg226tg
KVbAOA7iwde2R/oiYIxjJMMOhFtpswR/Q3Lfc7NUKDtJnlkf4o9LQgjt97uQ6f3s
DWCJfH6KzVjtdOLxDvTIj3DIPh0q9eeFM5LR5nVgRQBdvt/5T9AzFTB7szH3/4eW
CF2rZJNdJ0NU1KR87WOhigAM32fX3b7+I5YipvIuTZKzqK1GS+uQmo20iau2JzaZ
/a7moYQT9OBomfiAZ1EWIyWSGSvP7gJsLUdpSyJbQk/ug899VC8dADpBZ+F98j/D
M5wNnHf8xCdFVvGHI96hO5t08yiIJIiQcr67tWDErHfVlHddevfjFzgmrxgJ8CZm
HfnQoM5oGv5EjVhTlSZXPvap74tgtEETPxBzNlxQZYAmbyaAmsR22OnX8SCGqAhK
34kprifiaGRx+MgPput2z+KSHqfgnioS2FXhPgOR547qMy+mBWh4b/z+f2rvI3H3
DM+tZdMk3B4NQClsHD8iVBT1nXt85LWujUhjThaYn6DPYWWUicYHLjTPhXyjDnqA
wjYrotLLt9yXhjPqID50ploQsm7321RQ99PQxsnc/2dVIX2gHXqaHYl/DYgRhoOQ
06CrrRe5yMmboSmysJ/7vv5I0dzLcbT9jTbaITIHjgGSgbIgUyrX6eUwsuhvYXFK
sSMLkxVJstTQe9GI07nbpdoZE/Jxv/E9WyGhaqCzjGekwic1Km+uDAfNxjajDzoN
HplW8tA7nDup2UAUESvQ1N/BEjIAZXsma2Y0QuAbYYQWzDf2xKLI5U+U+b8nwqkM
`protect END_PROTECTED
