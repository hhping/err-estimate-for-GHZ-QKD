`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WabBk8PTkdtGuyaNngNOTVzdLH0a5H35vE0kqM+41dGogYOH37LIFZshuvPvCoJc
32ULR36lzeeNXc5nPb+Fj6sMFwVlSZ/up9hxc1Ip4E1oFxUrsaQyr9AzPmyfEJLt
cosC3giHWL11xSskX/+8x6W9Mui/Op5rCG/3QBAMh7Y3MZSq2MPx152UQdLhAQZ5
GYZ/FVJ3Uf/Rdvxca9ACGeuT0/aaTarmGrP4M5F2+YwDtaKlwnVgh3o2e3PtPCCc
QnJY3BAL0wmOvx/8QA5oih5hWI/0Q3JZnQL/NJZ9SbNZbPYyzx9GA8lIFwKvNURx
7RJVfpZ+Pwg0L73t0k+966+FZW7qmCOQKXLGhgmOdZABEpxXGvarIAmuIRAXTBqw
oqEkyhacEuSPrcyyG8VMP+EWFIy40NWLYw95gJfqRLASvcEo9Zs35b20rNtzNKI9
Wej3YsMdT06Ya9A1ojNbFwUkrccNX8mJ6udb+m5gvn3aDx3MZA62YNLVPUxTdkLZ
TDRWt1x+7Nd5QRR+4VHXMlbkuey68iUC3AjIbULew6CRO2xnSVm5qT4129NORP+6
IiJdiflI0NjEQh6jqUDWp+wVh7W1eq3ZxTTCA8S2wG7nOW8sPkbWPRk8T617C5M3
BPOW9ejpnBUHAbAAtIieLUPIhtn0EemV9s4oXDXi/MNyonj/HZ/seMld3alTT6hn
`protect END_PROTECTED
