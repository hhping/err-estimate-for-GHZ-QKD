`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wlqp2sjtqjN+SooBgzTthrDe39FrlnMZnz2FS6gov48G5XJMt0qBuf3Yw0INJjWR
fNbZi2QBhi+P7YhjJ+pVKuyCgvZVpwyxO+KkWKzg4nZgCaJk5pcUUjHiYkzj2VqZ
/W8Tm7mYG/hr+KO3XakkM/DCccwS8pugRYOO3JzYdvJdSveOx9Af7eePOIFBr7is
741H8DTMg/avArKY8opxHfVOyQcpUCESk0fDwaWGPMPFx1UODqjkut7i17X2zm//
Cl/becA6uNGuO9Y7vAdI7Eu8eEWYqctqAOuSQqGfRsontx12dwtX0Choq/Y6pEvY
E/mEyhh8T6/AYSA96wdJSE7r9VhW4Uu183gHvwp7aPW6jQXXSROAQwHJBwUxgybr
R9s+xz2ZJ1sc45DT096Wj0O0c4yOeuFbQFLQSuBMkgsMbpo5KDvima/GAXlhoshb
blJN0n32u5I9tq2Gvk+ByK3NGkXjW45KucERJtcEkeyEP74pzXAA5kB1RuEg+8Ts
EOPBO+r5f16EPllFN/wrro1A9mES1EXCM8wbPMR70SBjoYYg5jfN58IuoUbU109P
/xrwsa4nRzV86YDF8L4GfBuV5Y59K5GinDnZV0YSY6FlJR4byGYuzqZlCdSd3r1u
SDUnlFpiOiQX5AMtjdsSUc/ymEAuT6Dcd1fo3URwGrJd4yFS3vB6bSiwkA0NHGLs
C/lKLW0otIsSBhUV2jtzKHdmYgB0H6Nk08+p168GmoHpBRe7KhLndIsQ4QX8NaCG
b7s1F9WRWKHGbvQBzX7Ttp423blOBWMuZEFBnj0jluf0XVcV50iIPEGxzIhZ4QF4
gap31NrgudyHBMDZ29nIncTb7PG/UCOjpFq8xzHyYR0ZARaH+lgTkkOA1QjTYdAX
XfPYhkUoTz/0Nr5F5D9DwKYcfV+nFt3WtEdFpJYKVCNyANHffyPVhOwsFPfXMZW9
fzRrJFkpO8/QcBQMRgZhgXLVz1diH1cPYUzBJLdy2YvnlM4riRU/HLg/jxCGb3dy
4tsu46q9E4/8V0TNTn25Bx7hiwgFfxz8MDEhSkFDgaLVMX7B5Ia8hH7kg0Iuzz4I
uMWrg23Enn37FQRpaPDagYKB7LEoQO6hRQUV0qVBFNdtdNLhkVlrkz0ifyQ7ikNO
sC1uCOFlhB9fMhOqaF/XSLflRWdUOpVF+WfXBOZS5HtNiHNExcjd14pJJTKUtnoh
wL/gVA9icQ2VnR8rbiwNUN0RoT1cLzXQCmSBvFmsGM9IXyPm6vo2hNcEefvCU6vU
2gQbokDko4mtk/oPkK0T93yVqwhpnf2kVES9VjCyOnn+mTdR9bcgOq3FWRW2WbmA
+qbPLMJoTw+hzKP/GWfkvhB1V8Qr0j+dzskQZqIZf41yjvoe59jjB4fE2bq29DCE
MyVE1QUsOqVbNCNkg5jxh1O/jdPmgNH4uo6f3Hw6RE/jPdV8jjABPe1iFxUcx1M0
5SQ+/WTaXDNLpiVpSXuir6PNdX/X/ulvbkxqsit8SYAJ9xZISDC62LBO17Kz4E2S
vq9SWvZp82HL5T3oEeWcpUeNIEDmGY34vgu7VyxoeN1hFfmZSBig7cQzLazZkfQb
MXxKpVAUrYZ6xNuwG5wxi+YqcwHihNNkOwSKh2vdMSdYlzBvhRD/Zx/HtZM8eK0Y
5N/4XyrtoP7I4RC0sdVydgjJP4+wmmdBem8xQh1afbpc7YKDqlWrTN5q13jY2vIa
EvvdN0wCoEvozy19Gya6g2fcL9Y72eIIMR4uvk2O6AfcdqNGcgjDtIv31+BYulNu
qMDqbxAyPZHSW9iZdFVJeOsL3wepB3y3uL9bzI/d2I6vjAIBKKmxCSYMdkTJFl/8
/JWNiVYxQiILWK4oMzvuAbq72Qe1G8gML9G5syc2wDdD5Mc2+wKtaaRKxzmzfZRF
beAl6Bxtf7NZVXZyChzShsptA/I6qK6PVbJdfyK/U8Q7/Lj0ivvXy4GUR6sv6pVY
of/kiBlMmEiy/wArhDloUWuGmUdZmKS/2/f0UR4vN9acIlHcKQAJe5Bf68kDieSZ
jYK+MvX1QTlhdZ7JSDBmlyzb+2NADYRBrwkiS6JMPtD3hiRkx5LcDGbzv2y8QLH5
VGmqTDD3rkA57K/VVwwbpvUZBM574t5SXYPfQNoF9NqcEWT3w41+i6mTDFKLFQSN
EeTU11ZU69VAGA4B8EAi2t469VDx5La7u94Mbp8ek/mWbQA7OJ/KAaPUGx5nJ6FI
LTFXXuSkEMzfi2PNeCIbTrT4IvNpLpaUbFwMBShAG8iai9ZDJe5XQD1e0kpvZfSG
lQ2t1WWpYGyk7RQnK4xQI+EKKNHxQR7CRCnxCYBuBLXgkUmXv8fsqOGJH7Wy3L8H
bFG7XyqWebFnsyOobRJapKSwJibvoSKIErE8/cuCRfwhdXvYphKNonq/V35L8iP6
sKWcYWHtqPVGzaDPSyV9gTKl3GDWQLTNIq/kk5hNFevrdi8py1cr5AmZbt0DJX3b
8AMAlUHMtKMgxX4tQW1ZBe1U+/P0WeKfKU2IaugTDyftW3V0NLu2cEGjb+qniggA
VYnN42cgHBdLo0Ykd86sV0drTie8ZYC/d1RLOgiuPKsrGPHq1tClCAxK6W4hGl/2
f1G16QLnqRr7/WSAGkWRZKZk3TyaqH95pg5w2ThAZMjFk3Jx8/UbsT7oS4Xi6jwk
DbtvEqpgG9VXWq0OXxJyVObKjDXdb0F/0tEQA4a/cihc2bvDr1TCcf5YRO0WxUbs
W+SIq1yl2cWv09AVVyEOYkah3cuQJj5vZ+mtXh19M7GGhptlqpWyf4/iryY9KI7X
xk3Z/GbPGKftp0oKCXZ7/3acyHy68ulpmPDYu6IMzLmEFsvKCX15dd5oGZxRB+GG
2+NLEx60MAm4S0LQaMaf4kFgtikuYJtg1UiQ89gQuh2nAL5ixY+8LjB/8Nap4TKV
dzIo614agDhPZTmfHW7UTEAShlu/rWXUus1GjyKbf52f2iWUEo8UHsRrm9v9vZ0V
weLALwIP+vwYdIx9u3NagPh3DiGGnQNHavAsWAIusCALTqNgAWWS9uwPTWuxjRge
RJFmxpaq+39s2XkofMfi9McDFTivxnTd+d21iIind4vHwYKHOzmxTJgOTH97XHA3
5WYrgnKU5jAFRdOpW59a66GMCImhoH4grO/CFTfTqJ7RCcvT0LdOo9X02C6Nirqd
26lKI3xYU4L4uJJ2RBRekpjjdX2zMInVpz+aVmGeYNbTZoBNwscUR+ShrNRRaxxU
+vxYlV/SVGzx2C7RSRnY+0iWE15BsTzLH+AiyobpfG1zINIC0nTjtF6Z0xO3kGdB
RIGYfgLLb6iHr9YP5WG2ULcQZkzL5lOnRy/DAygWL+927jKZdMmczxmPwM2GfOLI
p4tqRF2tLDP1I8AnmYCQ5GTBU+mJ6JosjJKIAh8rjJe6NsxtT3bBvj0BbxKCfEIO
2OBiOt4eTI8TQb+lVuILffEeJFEFOfqzE0H07j9OtgLM4NO/z5/0v8PT+xw0X8VW
MpRvNgdIQrkPvTcG5gFLnusaoWbcnaUs14nGoqF8mur7xkweXPJewI6+Hdj+5hIn
dfWd1TroTGbk+RsyFXzZB2VYKfjrNblZOtydqCd4ceix2vLd9VLKCY4wzLEv3IRN
FEDAK/bNOxv3DUCD2RmPd0WAfYLzNn2WeqLjkJpx04DWFz8a1EK35wNfpv9G3I7y
AvTUVzd1Cf7ozTb2UVkxdQ==
`protect END_PROTECTED
