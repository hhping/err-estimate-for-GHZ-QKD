`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZoK8y4ukStK99SrPQw3vq4iKYE7FYCN+u9Qetf5SGIKwGLK49qPqYEZQFDIyYVvN
BLikErQMch3p49/QTa246z6zQm1HaLFBgXvLlbgBFs28NR2yf6HZ1EA3rtzncbAY
s6MogKqFyiI0F6nfbxl6RQNu3YIvWvNE2rfSOffLp8TT+k29SiMAqSZyY4//1dZw
mmWXl9cVKzUBU7j8Rklxeu3Ol4ephoxqsQZp+r4hm/sANf/HxbwmWmZLPS2d6zKX
tBdcbqePQ3UzhPlx1keZ0NmAchgpSulJcEFtuRUXUPsHBEYm7TpKAkWmDXkLzwjw
kYTCpMVdYsX4pCs33dkU6w8KsL4xBQimKxqIoMwbeyWBFXvktBV5sBgAhA4/pRrL
Zhr1n6sHzY9nK6KSP/m8aDR6+hhA3Yukg4lhaEBYC7sHhrdIRIJLMFUMGj4OS7uD
ykTbMkGgDaMha/5J0zzvlRQKQSUNHiuZ6pefP07HKpgHcplf4O1Rq/xpBZ8rxiFd
4dCzW5cKQmCs3OdlLzWVYRVQ2d91XwxdBa38TjKV7bMI0+7ki8v5Zlpg16MhhK1d
okjgVyHUHmgQMadSPtGUe1q4+rnZgDSiJivOipQy1mfSXsAFhktSC6sewLYl0bNW
IPGJGlnOZxUW2tDSn6HOya8hFHmoAV8hpIw5+/c2YxNb6SClQt63R/Pp2zsQMOTm
wKUjrp9jjGZrichy+T4GnuyPFVBIeO2GSktL+Ub1DZo3l6i5TuAt7Mb0cXapRP4T
DnO2csINwL5+IqWYhAMpsBAvjvsavmJkq6BkNnKDNm4YNIPWlKw5cUUqW+wet95P
qyBSKE8YRqrvXFugtVU+HM2WpuefBUt+mxhNQJOGUZfuaW9eri/rCxa8moXBmGJz
3Kx26uM3YOuDiZaz21yhEK45G4E66GE6/ljaRd/rUmCz3HE8U18AoAc9HGgqbWi1
w90oXsIsC1j4CXb8FyRlRJ/vDKGJPsqXsL3N63TxeIJ+L4lUBRUTvDgTj6dW3oBU
GKDdDzy4U4YUtUyL95xbUCXVczaIYCzRNqablaqOpI6b40Nh7HvoOfRm1uIx1jVW
L2OB4bSSHGBgIk3j34xGRDxn9XEGnqOWq4ydOzXn7ugTXpRtlJsBMNZJG5bTf9eu
eU2Z9zgcB4bhMXRDx85sANOJsm/tttv89lk3DEwYIMht9UBqtmH0QDCoE0Ha7ndQ
Ag4LNmN8iItp+zpTjdrXeA==
`protect END_PROTECTED
