`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lLDUsP4nqhic9WPlqMHm4JB8KFZfkmWfzTtRIQxUHrsi3pwowitDgN0Nf8VZ3l+a
Fg7/wJ0pMbQPRtq2F70LRw+VvasBrWf3AoKu4460cANQbW/TZXYP8nRCG6n23V1b
msiLv+Xz2O9R/FExOZ1pd4CqQBh+4D5Dw1IYvABuzwxRN+wqBgLr4tCqrnN+TPUs
NLZSu20610u9uPl9lqwaEnM07SZI7vgJxrwC+zFZUeA8aeySlyOqAL2N4ATzmY52
ujmE2kP+2emJnpKdUWFDCOIawJytOXKLoAuBt6JIJ8S2W+iA9OLDo69XJbln9u+L
yJoVOY8FsSzc0KBuLFYTt7vDQCAqx4+oc/XGACxs60JIfN+Cforn+eLVZBO15cG/
PNWUN7yhoCaVM7dyJFhWbpmJdcAR4xII6VYbFEngyw/uCA16Lg925WQqeyRg0Xo3
HLf4Nh6df6yDhnzi+VDlSH98lrSuGx9yYPJeDrVCgA/850CJZdAHl06+Q6oHnM0O
KghJhhu7cphG/BVt1XuQB3AYGKQXw9EjCCH8lpbBEv9xg+zjqqTe+/ZE7s6IAt+T
1PumOZUo0wA2uZFc00FKSAndw4p9KjCoCq95zVVzHoSQi52uk4kGRiRW0fa0HMtX
G4oa482N/p3qwVqR7nxf1UHEPRVCc8grvTMgYFxAMMImz0mKWABwXtPdBCP2Funl
PQ5a/DQsPbY9YA949ACqWyZrh36cqohmlZimUrB2xkJs59eGxmDU2VPUEAJM13/I
H7zPHnNRDX8TcL7S6ltuXU3ckehEidhVDNSzqB1kct4QrINYY7Jr10Kg/to/7tuw
C5bSZqYLPKFr4tmuzkZjxBI94jp0857rB+Gts4UfDNwjgNN8zbgyQh8uNf76ISV1
+oAwjNs1mDxINapt4q26ncmE1CzGZ5fm4p5I4kZ5oNs+5lreJdaNJLPnwARe2B6j
cX8Wy54RDAnvDf1IgUPb9W3tBiiVQH3TlDjqxWgS/3nfG5TPYVgFab/lWrQtzQug
Mt4AXPpzHizNNDYUVWeELqMs+FaKVkhIzkrbm1JyGVD574cLn/hpzmcMisp8gm1n
Drt4TkFSd/ACbdcddhyC/tHecUGbH3apJuXVzNt7bgyK/DG+O0dPjYELMc96KNbL
7jD1dIw+TpAvTie/XvjCCsPl/g3C/U4cD8H9TkNmUoACGOIesFlyaAq34qhayzvm
hFfQhZ/G98RY63HFO+k4shxLEzedqxG7s4Ugl10xvRCIk94CAl7iONADyV0uKQ+0
ak8F1Xy7IL4DVhEA+V6RrW5zOQzmR+hOF0fIZKqrcEeSZ7h/n81KI4uQLwgLEDeN
BC9sKanuqzim3BMO2R1kA4FX5d6Iyq0Su9vpQbgZ0xGXQomYZIvBRiHbYOjputeZ
Nbw3YB/yh+cPz0zKV02IH3T62Ugu4ECTXlYqNRaYBwir+mV2bxDbfgUse81bVTtZ
sDXPIAHJx4BaGqH5y3GAa/I2FHxTWfNEIkOzu6UEyqbl93tKxpPl50MW2dyDtMJd
IEGUAa5v5zJefhrgCqQzi7YkNhlUjrybXFJAJbfqdyTrKU3NPri5BcWSRFqpfefN
8kxaMeyeXK7mXws3s6eKMXgR1Jw+0zW1pptD01MbxzUZNT8TULluVftwbNT5d4fP
ox4T82YEmryLdreMKl6Hz0oPG6oUbdeyqoZFjOOuyHdlwZN6Rt9MivM+CyNEcjAB
r/XIaRSRdas2FXZ201xLLA==
`protect END_PROTECTED
