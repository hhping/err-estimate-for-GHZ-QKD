`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U2MuTwTfCz4JURniycliQCvTzjb0xFP01M4dWNpwFUlBLc8KB4VaOoi1gM3u29HW
sVL7UHaaPvjL9m2llqap9sKEYyU2R3TyWFrTXnUklO4GmeSf44w4eFe2Mj0qOEHE
RevGswLUvQa3j84dhBctP1vx0fIBjv8Ny7mpYLYFk/kTRyylTR+DeLu/6S0gqd3Z
Mqxg9XD6Opuhu10EtW0b/qdexL5QN0QkzalxfcwFwHz8M/8P7CCxRHj1NBk1B3j8
dtD5iWvTTNEhQ5oLh+XRCxo4PQORC0JSJacZbFCE1h0UCtzqTDlm0A+C2xrY163V
LKjtW7gWVW6pDThtOOD6vR3uyFBCVPnFMY76NDxSTg40yYrdfKGpaJSwlGD7RGzR
kgL+cNHqnZZlnJcrm6ZPLELJOmKoKfz6khLAYbjK8pWRfK0mSY6iFHE+vksTKigq
i/lpnl8VM40HbLff7uDYFHogTpd9Oi/ZrIgAW2ZfRlDDgyT+Wz6NlWIDkCCo53TU
wqlel3monGyPWSzNNBT1OQ6gHHKxhrq1TVW5ell/e/+cqYJo6IRsq9YPKpY+Mmbj
bwpisMAViqNx2lAoNAoPn20/boT3Ck8ueVrVoB3groTESkcY0l1JQ7YHD965HEh/
iayDfeVKfKkT+BGHoO5gKP5rUIADtH5IYfSuJqvmtT1ELRsZ4FvgO7KJHW3WeCOk
Ks81+GPlcJ8WsIP8gL+TKLm5PRPKKANkwuSTtJII0KcveDJGvPBmwL59b+ZVu1hJ
iKHUYFS64PoMM++sI2WoC9nxjV0HolehOjel94YMRDHWSkTZAFHFf6jj0PUA+ft6
HDCZvWHOueOEKFOeUCdz2crGDGntWzY6UortwIx0QprXs6q2K0HkIc5V/5FGTHyv
SNzOOoVYm4WNIT43YWdNzc+Ie0T7Y4njiHMJtehBQ4FA9s9cKCoYb3hN97cgnXmh
p80xoKT6CM6KJsxBEseos0aPDMWmvi4zEINbbplfzP8A5TVOA6rc2DMfHPBxRrM2
N/4hBtfL+mdR6WSkFxtg9ojax+xVpAcwPz5WfZg1YXVVx5ms8/5lXx09Rj0h5PHe
A6aIf3dRYqD9Lp87DB+lTwxUR6SoYoGviJ+nzH+Mvww9rHQIHl6Wyo5uPU376YBL
Tb9pcDohwTyPIrxd6LAXoKM1l3jr79akbdudVBCBhON8T/euswJM8TFUs9tzd9UI
jbRVhfi7qUeZgnuiLtcR78fDRdCieoveYCiOyGyfwf9S8y/SQ9giEua8DNcA79t8
SUPEF7+4GBLZsCm6dHkVGtx03walgXKFiKK/qBFt0ivzIjlSfYsumqcSjJ5eCleq
ULaCbvvHUX72rgF6i6zeKWOEVdHepN+xLR76qHLq3RCXJjj12sZMHU3u0/qJYliw
AOF4RL8xgOz9u2ybKgDdN6VR/GiT1EdI2ZhnqxGx0sZgcHAxvIL5cB6he6ed+5ST
M5KOmy8AN1XFkT2lIJ4dryfMVR0sFsdL/3RlxzbzWzr7xO9ME+Vqnq7BO3amctjN
NC6pENpRLlUDBFlD7JfoCYaJANMF2JvDjmqzCzXQ4RqPaqWT5gEdnqqBR00+TzDt
Ctx2gyHj1FYRs3Y1eMnV1ss0fK5A8pzmplnyG7A2kAWv6Y0qy87daHPI9TrD/KHe
80zGXzzaWZzkoAI6eSciiv9esqrJNswcFNxwl5tu+d9G9XaUXl1hjVd55eyE8rtZ
TU/gHGtnutHRT5ZBpqYP80pEiYX7hxBbNGoi47pD/gVNyZxS8eIF5+KP42rDSvyL
15mIytNG8CCR1c5Ir/UFA7M+lh3K+Qq/SYDu+Xbz+znUySJFfq73ogVSi0C+koDt
BKRyC5vUNEI7+YTrhMQKWptWvxrcw7kvX3Rqe2sPI2v0pbaNHLgxOflWa5Myvn7G
42mxBqg35PXIlZ8pu9K8uGHsCUWZL80jiG1gw7vdvHz8zXhvZu58PHGPab0tReHy
x2pV74GuPy1oha2jbvOuymF33KAjCbvjbb/pnbWgg2Iad/A/CxQv5EWnVUJive5K
Nf1f4DGIjFrUr91wEcjROurS0VyRmpU6hg3mMouumXvpejioQbp6QauOtL7jHgeI
RcFdDeloyvXWU7GtGxdFSAA1sDvXo8ZO6Am/N8/a7lUOJqr5gZjZrBEf7047pm58
jnFDFIxjiDacILDQhaTzgYEy8kLEQVY3SRx3wO2H+Ssek+Z8UT8VggecmVS6zJa4
ZvdXoLNH0NnkPRGXebsJ68sng/5Ch2jzyiwTyzhWopxElZD6Idy1zfzqKOvSv2ve
NWQMcC258kveQ+VC3rYzQy1XWxTv9/qGz6EV0CzV69Jijxo9NozyBndNTRr2xSuJ
L6O2ESLfV7nqgQIxqHyyV1gLEwAv5Bzqi55U5AoUQBRkaVUFj3LRF8YZURWwpv4j
+ADQ0g33V0k+ZFP2WfBqhl/HxAfd3HI3xmedHErdGqTkAwNqi6QfirmcZIUdlfNI
AQlj+a2VF300vPiKbRwloDMZkCukYxeuOapW29r+Sw34pKq3YjupAlSKkuQa6wi0
IJFcLx6APKixRq4G3dlUsn1k3T1gpyP+sWCr0sSfovbbjDE5h5GP0iYEyhjhPawx
4RNcfawKBP50WW4qkethfINhoD0CJ+tXjHSkfCld1EuEUMYVZMiOQFGzYMhXLuLc
wqCWGeIS0akS/rC8sk8PIGAGKOkqQS4nGMa2tSt2rJnM9wv4VAE2C3vhNBy8kQyX
IMSNiab4vlZoyHYPhh2CQXs+B83cKQ9WnxHOSh0tF8ty419frN51AW9bYr/XuE1P
/5kB7DZvXuquBOIjY3NtemzuzQKAHTiVQWxM9n7IJoJ9inOoJf7Y7R0LE0wwOiM+
mIH+IGbkym4zKgjCcFnIWYJ0Y1BqCWThgn3nmlfpzgyzhV7J0WmtehX0t06svxRO
5CH/sk9zuwnGZfHY257VVcvdD2+z+xTHIX4H+ER/kOmGWIRt+41e/xXxtGB2/1CR
DEc+wC3Ixik3xQbZKGnHXvBGeRUyicg+sJkC027L/M9Mm+lT1yxLBb+lCZfemVHi
HmtcHdHoRZRNlVH7zzDQ8hkofxWjlyZleTxc0uAD33xlO8+Prpw4/yTKBcX0z+0D
gBZ4bOogt5QlJOLn3JakFYpQ8NOms6gS3tdC+joRs7uRC1QRMJt1xMutqXR8on95
XkmNRiFyS95BtjVueEVgvbLBynnR+rtLodAO+5GUg5TzqKKVIWT6M4pDzRkPUiMJ
Pj6rS1EZZLCQl3YFVEx/H1RinHcyi2VpEtn34dj7aBPWvV45PBQZljvTgUm0zhP2
pWXhftPtK061urYZQtRvQb2qY6sfqirahmA33eY2jiPyfwpAl0sc6+JxS4meSya9
NI+3aZwYRI+aruEnJKzpSlGBArNydjiWlG4qDXMPOhJsJAFGpUYgHed4kzDggY04
7/auPkA4PF6JxGKv+sYIlLWcov3Y1cAE5Olk7JoYBGr+tAJCGz94I0NCDYpuaq2h
jXVfQvxpZdLilHHZkDTqAlekETy2QUBQeI47eDpV7LFG2fnBwl5njxeeXJOjgS7h
UgJ9/gQaOBLeNQOuOXKBZd7+Og1xHmQsN9YEoLMvJ1ICcAEPkZz5R2l6Uio0o5ZC
HUvHKlZnN2TKtIShY5mxbH/86QavJ///xttKeVfZcNGNrCtEuKdr9+3nXMBP1y9O
Bs1HEbgUKS4QQwSdeLU3Ki3ipGLVldhFAGAK7zsyD90L+bJ6UUkH6fmcC1DpwIZG
o/H6FebRXBc9TUE3OKcAYpNgdnyj3sTnsg1RMZdT5iph5sxKHjnvNSASKOxHSjRM
/rQvFzRaCbhdRA3ppt4WpdmSWEEUfqwjN4dwsDrk7XJnv2TL6q58AEy8EIBqFi8t
G33mcWtMqeB+U3Wrms0QLsrMMK0wzU4+qBLD/kLD1/w/mlDFkMEc/LHqs8K8WagU
8W0BHjW4an81w+ZLHl+UGlDKwkrcpreTlYrbZvIZpilbQpcGJtRs5D6ADJmv/9bJ
ieKjdWBrR32Q4FUO7rRsCXl4kDwu/gnAWXaUimc7u3aF7E6RXCLfROJ8QWEfDJHn
tF9wLkGArJp8VkaDuSjpi2xErimY/FAzu5d5UR554lTpxryCKDzuDPpJhrJVfwn8
M/GKj0P88IfesScD7d0ptsrBh1tlzD/tkPCo2C2nq4b1AsM0NZzq+mB7X7XZkaGP
MvH58FHWI/Tt6AwN7PjF+COjnFX3cQEKL40E+yJxn+gsLx3ebW+j6RI/7KpS7zv7
FjV0g0oeXhXCkqirlm+nVX/N/eMAtWDceToSmh23QSBWHsjRZev68gwRIs6J63Ip
Q7y6cd4z/Ba3lditJZ0SOGqxSXDLom9z6bTMFO8fvk4pQMsQi81JIVKpyMdvL+aZ
a6kHBJJNvnEACiQlrhkP6spZobHT5kLAolU3zUsb2PUFbfJOrSFDP52IbarBD4dW
rmHCNpv6kZ1eCNrqHqVqik+ZaRKszjWJACyzLe2tT4/HM7QEU77Kqr+zWsUfsSi6
5A2lUcWGhg67K+di1QsVTzZrfLf7QHWpek+CuS84/A0l6fTqwW+jB2dgkP6q5XKS
iy6vnY28EvRucBTjgebUHbsGhp4PlrsPRERBbLjJ9JGW4SGtpsIM5+dW5GP42ZQe
5ry3rtjrRg8PhhuYqqaCgbktPrxf2+4ulVnKN/gm5q+tDmi+nKY1Cdx/6GEq+DdU
fEb2vc6/WZH3DuXNkoScvscbKrzsjV/HbX5mPNNu00pgyxf7u+7g5f2U9I+qMQ67
V5xD3OPjVuK43sDxHFAaJ6DIL8hb/GQ46czhW0lg/4MDnWhwu+3fRNsCLpCyZ8zT
T8sUq29R5w/Llii4WTSZzQXElm3oZO1HJGepy0aeF+zi992biGvpTI5wBoWJk+2f
OFL8FEu9MgQ1PZHs67Z0w97iMkuhIcFdySFnfnW3w0FzxibcvB7BHbcovz0+eeWn
JQZySFBBrHEnsOTDwoD9JT4svXN997Ian45LGHZHQv+UdH8GjM+i5ZXUMgdOe8au
0QJnoVDAvajSUNMuiIbT+f2CPqrTrVZ7WB3vr1DxLEycQNoe4l066HnwdYqRKK3Z
L0WxZd/7h8qLixBAaPlrMHup3b8rmzi1mHJ3h0QsaV7nPA/5ZubFb4Rp6wiK6o7m
Iv2unLCMmndtfJF0b0HmetWhO/Kj3EzD9r/BtbLuTwLAn+ZaGMD3lVkqjHqsPuFz
sJm6tskDBJ3fhBU44iU/Q5+TBootUTGQLpWkx91i8gsI3zMz6uxZOnz3rGXrkil6
yoFEcl1M4Nj0HiE/BAfMBXY91xmWlTacvXzsAnkbSSBTvvoFwsCG3c+LuR/5v8iM
HU7QUdnrOc0TtEOw19ColNapfnDTTHwRk4+ey9/uE0zmmN0Nm1RY97/v5b3wmHwl
WGUTyWuzqa8fY6cYBMge8s3yM6jM+736lTBmOlhWVsiYcnQEk5scnT2kk67HPqJd
DkWI7qfAS3dRXbWcH9R+pieMW9xF54HbbVsbCkmobtJsH1zZzLRh6OSVsaUeupSy
b2+kOptQAFtrbZNsAh430pMjhH1/gTCAo85xcghnYLid5MVTqsQs6WjGumw9pHfz
9Z68PUU/7gmVF8ksBG/Lsc3xYeS1znFWMKXmgvhvkC6r8Ttt1WK+9gHKLjW68aDm
H6f8T6R7BQsbV0KBQzmQxi4xJ9XM3vMKP2CsylxyKCe23J78T5S9iPkkWnV3HZIe
HMDi8BGm2aZi8yV8sStYgkFmKpNjFnM/XJC7bqQ4dP+PGtj9jhavVjhWR+wW95a5
b44C3Rb9DA1aU4s4wvjBo+ssAvK3a4nk3gn9uWJSr/tWVrvZNNVGHp94s2fxRe+R
FPayHdOJI7T0zx9/tOFZmuvXpD7QiWJvZKIA/Eb6rUhzOT39Ph8BX0BZdcus03az
6eOmRv85IVGPcujVW/EDzN9TmkRknQ2shvbb+HHQI8bBSI8bjsAkxuB7pBobQhpI
fZOWRuSdqCMcwo4fSu4YsgAZgn0kRSAv6azqY5GFr3WfosmzeJOrj6R3NgD2Ts3j
7f/ESRBdRhTGE2xeJ15bqJZ4o54klWpEYONvyT4CRgEV5swDRgJsMzZtusFq8Kkb
z8Eb4ZgoUVYayFJBBS7xc+pISdbRRZ44CAcO7kwLW1wf+zLG/E8piZquVucOuo5o
oLbGyglMUB89/lrWagIZLNOcInYn9vyjPdwMlfu+WqQ1khOwf2sTeiUehVH4Qvp6
tE3WnbBx5TIdePzsmPC4WAitKQ+wPAcryL1RR5X5GD/6+3yjXiEd3SrsiIsgfahq
809FSSQrJDuFz8vP+NALaY3VQ/hGc+eSa05Bzb//vuoBbhqYdE/FLSrmwn0Qfccq
TkV3Htnqdm3K5ppQdo1RdSOSNJtpOryTi0S+86orYpC1JkyWHVoTd+qzYMZhg7st
a7pWZg0wk61aZ9xAhFWROdzGhbQO1ZcJxeW0rmxeXB0coVt+WYpf964HrxUTB5SX
aHZ9oEYL/5FEqWMMslTEA4as/kMNh+/VVttS1difmp8kfHeKGG2n0+gMv6iCuCrL
Qe/hmPZUMlvWpuWztYiTxL85OlpgHgGpC187L6p25qdvM1EAEYgH/BN1eyb6C0Xf
RI9J9EgWBXPK+j985Niep4SRZs/fP0RRxnmIng0t+S+En3R0519SxppgOoImXfB0
QI/6hhdey5N0sto+qCYUMnGZ1iDRpe/UGxP7Jqu8qABsOu+XkueTSGlWQJAhe5kG
Vy0DHimHVlQneaY0+GEPQrAHG44EE76r60rSdqCKrV8eipf088sS2YXV8eBSE898
/t33IXCaLRegrxBCHErTg0NqTYpUfwdRgFVCZ8A1pIZVDda2ng0HshQZXoTiQju2
OiFoy1EqVyvK0ezZnEl9ecwx4a4kSqPJdj/6+E2W02a3P/KwnN3ByoJ5mcY5ZyyC
8rKydnIAD9g22egntcIxsbImMgxC+LVRoROGegOnSzzddmA+C649UoV++tIf7zoh
GytsjdWUuBiF4M21D0riHHFjdt/h9L0nnhH2fnjyxL2Fg5vprhiK1K4zGpE1BDGt
xSrYBT50GWaV+Y+S0y4kx4BEn9TfBFsRKf+ssmasO/GHXnr0RKCe7JJqIvS2PFgD
emKmqk8KDxiiThbO4K5lHJ3+cydyVH+VZPxr0YS9KYnke29BkpDdygLZQZhqrZmw
IIGOELySgVyP0zaDajhwzcsY+m8SZI4/7M62yCj4gKUXrsicb1pOqt/4AEo6jEhD
kSTGOC44XOeB0iVbrB8i/SW/pKiF865qa6nW1ykLIShZQ+E79Yw8mp6eRnmv/Dkb
bUpfQ7D5QuUi8z7Boax6JzdykTXMYaRDbs+g9qOvxZOoH2CeT1aud5rrbhNL65pF
jUa/HeD2/PqYnWGgwIa6qCBjWnL1MOdFl0sneRE63sTyPJ4MAEiC+km12MJXKNBS
rhThNrkSU7pSBgY/XNRX9MiS36z2wZxfQ7vQbBjybIoPWxrevEOr7ox+S7KMbtUV
vd+QkHeB3O2YtTgjXMPqtTa1pHPBs4fThvJc8Hzcoo2DwrTPJGY3CCDEGqHvwl8r
ZtLMxu769o4tSmjoAH5a8QTSlE4pHfe4bI3kfEjiYDL7qmZ2FeuAgZzlMBISP8Q5
JcdvFasG0ZCZKlXq3PyL21ceLFfdV0/vXkbnx6KSgI4Y8VGlZMVxdYC7az0fCO4/
k+3kix+kqSwwvMKBSRgVEJcp+UzUdhIVZ34ULrDgoi1Y238LB7Cg+/+DxMzXsz7O
B0bxmWToFxnwui74oKk4tlbuBFz8xZUh5UQKhqKtBPoWUDsEcku3d49Czh+gp0Uw
5/2nA+YD4myuzrQ8jqH0jATAMLI4SQl8pUEgPIFrWqFKKzAghO56wTbtGWQe1l0y
ywweISzwHlFuwYStJOzXreMUcRQp44ha4CFqizCqjvcmvrsaJGoTfd+jTm4Ha1Cw
JWRwF3Jd077g6aKlPkMiQzYY6Ip2buuuybDP9pMBHp9VASd2qACX10NDtxRrsSw0
8UHEgOxkxeIEGSkc+FYk6qEv5dkKlxEFIJO3MVZBt/tDoOq1ka5Hf+/w67sdYmQF
il5wBGVjLNFohOcnJAIblF9twq2Nu1vHuOhWexVfb4b15rm4Tl9W6eFvBNGVM+OZ
fF1jX+Ty3mHF4sCNbgb565zNcH+Kvf7wSHt+LiZHAN0EOBSH4Ce31A+2xCNpqEB7
HNk7NvTyvW4ga4HrNsPum9i+hUc0sEIR37rSi/6XHsVpGmQ4TEyM//l0yEd52MkP
NppWtk9Dryju8clXnTf+DqHrO6i5lNsRpJSpmpGW+tVHtfXZB2Uchbrba6K9Qyzt
URXzRknaN3EIi6Tz8SSDHGvHWf+oxK5fOCCifvLBRMhGo8EPfULj/Vuli/oV0AAv
y1IpMPqVj35ROyslN363KRsplyJk48imdtaLl6Ipd1MWwCLFuKSfdmpztwCPtL/P
6WGoVBVfhN2/frBxPGcYCXyV2RCV9pKQxKS0bwDu9MIQm2L9rXIGQiiMflJqhK8A
tA93qMfhwR0wEqAM4gLnTkBKsbA3VexLz0bdoZtxvzAUfjEDrP4ZdJgADmUXkaeT
U7gq6szXZQEyaf5M0tpbNW/0AKTQbJOqlr5Xiv5bvJUFRNoc+KxBHDePuhCgqQxM
pxHPR4uzmIOO8u7TY7Lb+nc+HKMXFNad9mLAlNn7M/pCSwV50OANcvUSWPvm+gQY
1cAux00ayjYattqFTLumVLvMH8e2SVQJ9xdOM+v3JtTcfLqVBl16jOh+5vDBOGBM
fMIDjDUYHE2/cw5y6HEiVZwCAnjCzQYKZc4TdB7HI5c0U9o4aoSqpTLfGlGny4Sw
NJTkVyBHQGnfUCyIpQUV++BpkZHPOlbamC8ML8gi06bNeW1JHYkU8p37E6Ds0x6C
OyQPrmo0W/NLLwr6JXnJcgZyP+uVq6fo2Ncto7epy9g2WuTyUqidXTDHFvffS9+p
R5tmvURZL1VhH5yQBpC6SD1ay6aS3GKYi6msFS1olCkhAmcHCh0XgDzZlVl2n5n5
Hza7DAoHjaCHBApC1kG1Hz+JPWHqRwP1Twa1B4F37j43UqeRVtlA1t5CWJ1IY9Lf
yvt/Un8NzYtqB1mEyA2mKPb0f9d1+kbzlOEP+jXL7/isA4nLWnQ0vsiQ1/sxcwwq
2v/Z3F6iFlgiXqjDZAKQ5BZMTDS21pNz7bnnUiZH7eAnKrYlOQgNLvXnlJrv9hIt
3/1KjCcNEFmAbqOhQgJ8rGYKp8AgAT4r0HpddisviYWW/sy6fNbm+adJIB+5JxVH
ZEHk4vZvUL5Le+WX4BSQKr8MpXR0cutJlZKUgcuAVRgm4uOoZx6uMGTf/FJChDYO
rkVzOSEKQ4poimKGX+tVGnuWCwELQlzKYOZET15czB39W5LQkEa4zt2f8UJiVb3A
IR6wFKT8aB268eGGrpqxqpZv6M6Xul9HpcHRBL30haX2eVYhJYP0ktAh5AqPHbMO
mXXxEnLhjHLxGUWmwDAIIQFMs6Xt2gTNEo73EzgQCqsHcq02liKqGDF/IAOcGcpN
QHdHXo4gVRwRAekiOHB3ztzaeO6nGmNoeL15Vw00hOQD/nL8huNeeaSsudAVOoun
wvUqAwYC3hQzS06OGsZ+nuZZrmJK7JmpwyAUevDNfqlZ7iwSLf3FP7j7SVkZW0ye
Q5OQQFgYcTDWjdL8mprt2KrtrI8BKEk/leTHxOz3U/r6Y8/U8wSIWG79s2iuMgfS
qI7TJ45SACubq9AZL39bQ1hM0livaxVYEb+iZ3njGrDT/dMo920RD9tkFl34dVP6
jPGq89GsNvpFkvT7PqiLCMWrwAx2QJqWcKwAtFCBhRDsqqeImpre8FgwiDLRVLd2
/hpoAmmyuGBVxgsCq/C3o07UypNQxjCEFF5LCJFtDReuo086sc2Lmxzr0wnrECPq
m+CzTldlhT0GTLxJrybZyLsIolDmtNtYx88SRgYw6XxIrW8qZYAI5Keyr53MEmfY
wAw5Y31oOhCpwADuWKv+QuGrK629KDmkE/lCnUXMl6pwA6gB4qx7J6ikXTHM2G72
67mAYl2k/zbI4O7qic+fuDgqmHQdQykOPP+4FNtUNqjytt1XxNthTDXSq/pd7vpp
CJPjWjR7O3cbHuTa1Mr2LbT5HQgjTZK8E1DVHoCjPCqSeKtVwoofuDBVgmL9dQHC
wmQkIMBBID0s6SjbDYGNV6Tc6gTE+ZHB5Zz92mppjkj+DpVcmewrGyRlnNTjWMoy
HWr5SRx5KY5Fi4DBG0HLUE4peUtqhyELBz9hoWohdbslifrfstcIF/0Lfmb3xeVh
jcUncqIrdeCwq4bViy2jk6lMNJPS8Al4hWXz9qItoCKr3HPNYCt+mVna5MjswxAN
Z3MrZJJXCNsINvta5DKnsPVmisDr+Yjw6R8T2mQR4lNe9jpnaV2YKPGw/JW1CWrn
8tx58U1Z1KYaH/okTp1WeI9Ejwrv+74Uzln6t7XmVxdR3VivVHoihntkMEpbR5+l
qvjOlnFU1dknX3vS52XVry01OAIUXLVMQczzAE0G6Xpl8wvgi1jr/Saf1HExxSBt
71NVJiimU3jn9hQq9LmQbdT/AhkFti6V2yfoCYrvRz+0PzuFqq1SXfizJ6UlGjz3
e7Vm20gXmGiMTKpIu+/1TjMBSwt/Qs4cIHxSowT58iRuAl+EMXUttsyIpXlLlU+4
4XwvU+TqRGUpxk4lbxQ4hmmI4bC8mRD7V7ge4wS8ZBvx2XOEm4BxC1L/M6WLP2qc
0mMcDRrjheJZVHrM7GfBh2n2vhJZ/9LjfiYcdqEdx/VSdPCDIK4b6TEUb2yXVVT9
Jx6Xh2gK5B0VKzmP+Ulc57X4sm9sXE2vY/era4L4AvUf1UGyeF9OB2mSg6Fdj0u4
VpAvy8jg+EZreI475eBkQGWeGJscNwFGjsvU7/UHDiACA7Bzw3Mtv2mEwgJBrEp7
hvH/C9JfYxrzSJj2NgqAvZ/+r8u+dN5+MdbrQ257yCkfb83x0ByV+l9NtgW44uPh
bORuY8+Qrq61veTQGDRB9D99JrLVy5T3ZR8aMXe5jXhVyM1vDxEd9mIj5WwYPO4k
JRFLMPKgxmfOYuIANAmVZbFaAxcjoezmJ7BmYZj18QdtGM17TAPpHC7cL0JZFhWB
teGw7rdQ/mmjB9s+8nlZ2x1Z8HjSHMMw7Gxgvf9frfYgd/vxzr96Xocg7LX/zlOJ
JxC6YghlnjSeikcqk1tE/Fjn8NycYvWm5VKFXECwyj443sQVUXEUdS7050VnBbvt
YpWqkQHZpG8KUkbalg1wIHE97go+XaYHlwCeSKNolGKQnGx7SuXwhbP29adLadUi
KMKCbYRtz0VlYXbmtIUV5Ub3xuNsH31DixRuvAHG2hc0bKXDcD64t+qTVycrf+F5
r7kjTrjOQ+CC6Snd9DZtGKOJxbJUNrq/cBtfK0IBz+LFYoIUbDTKJEjYqFPZE2qM
wPRXNLfffCKcGC+wjvTWUeYLMsZidW2hX3Y0U+MqXOKjNtiQd5RgQeqBJGDAGU/l
dzeI79Qci5SpuWTAbLiJFkNXaznBwn+bFtTkvyODDmQIYRqG+6HerxQbjwrnqTFU
GF9O5PgDacFvbdb1fGykUtFnV4JkqGM7Z31sAmRE6UNQoAPE6MQbXWWTEK0SvcWd
WPpIAtvML81idyTxQzVYTAAEOijrTka/3jwrQ9vcY+8KPzJiQbT0WKTXyGaYvUJS
t+G9dew8ivS0loBcbOr+Yz9kI3iMSmyhYOAP1R8R9f51J/Ia6wfI4aCigTE/gAZd
tk+eIxGtxClr1AjHsQA+lh7/vm34F46cprSRFzJzb7wLY2Cu/F7Dq0WdNAuDaE6C
yFaTXy/Htou874fLJsw14ztwQiznU4NGIu4xe2iVSEa7NWr3Gf+MSiAdKgHybmyg
53u5c1i/YfcQwtn9mVBXHIZIu8Q9SMyPmLJA1JxHEbQlxg6KWOhizFRIiIx6lmRD
vQWPX0+6acmMfJ9WiltXfd0IbIkNIVdJY6ASKEuiX7BCGdOZwbhBtp1iyTx5pWVY
B8ziY3Go7XvEHhSPjbCaC4G41eSpK0IzvTTHPiUo+wL3LsSNKV4ea41sedpAE61q
oIIR3XXjvbARSx7nSE/vrb6D6K7rcLTjjbx33yyXQk+3GLAvQuAqn2KWmgwNNF2O
nz6K0XHy6dIAKwfZn180Wdi79IBNTisuVOEI5Ygpe1R8nnD6KukGlAHUmFalT6Ww
wDl3J/enxELj6KMHXuK2evfWInT6mkAAdqjYVXg2KzOnXjxX20jmu5hBT566sGhC
wKF2DJ9TtzBH7iGgMaly20pnLkI3QNhdToci5UCIk3Ff2BcLnzCiMxWEd1Mfbp36
py9NGMeFdtPOKm6Bhr8nnUS1wKYT3EeLic3sSJnW/iVzZKzkkAKS0xGlStIN+aqh
iN+l2shQTv/hGN3DPy6OQYOR4L9TukXXlCWYxcbuq8aMwGY9Xe6qNKkCVY/Kj777
bFTrgTnNxApbvNUtEDIRbBdbyrQr5NJmkkuZ1bDlxS6l4tk4HXXiKxJT3ANus1Tq
bzsLlAQWWumpo97GVMjLgO37DDUxRRiinhO9lkTKO8Ktwm0uUr+REehWyyKKKE8w
64fH229vG9Wj+Wy5L1ySu7Que4qJzgRPGoTd6ViIfaM4ow8DZNkfI08Kk1dd3MXn
8CP5hjevdeWpxd3ZCbdN1dAwvRaQb4CZUDCSzkIUVieaTnJWMAnnERGlKMH3BPHl
uRa81eRvO+xva+WyfRRNAEqaJjFzza2XtIpN2hKOyHYVT7gbzssGQ8NH8MP1cc4o
cEdKKKJf112ccTNy1q6v1p6xc3Gu9vDlcHhXMmaf5eK+jp2iZfXyTtl+lzyl4s8T
uHXJWfevLZHqrt99ALEUznsRqlbq5aHrsmomrk851SpTCWpwHPY+ZRGrcEcXZGOz
Nv6N10gqpJGJQ7eU8QEE5nz5xWS30QTX2VSDgWS5SCOk3RiTG1ibtjbvW8q/jaCv
sbUBpwI9GUzg3E5SmH4lXxneslcJZzZCPvrGuOGJ3XaxK/bE96qLTJpcfkRNOKNF
skCLKwl+6pG4yCf4X5F4UwGXTZM8lxYRPPJoblye+qurS+6eG0CNs1LA9+CZ3ten
XOgqElLrxbW9uwwgF1a+5aUWUjihK7ZSVYwpz4TMBUXAArDBKMgkCGE7SoIwW+Yt
42qoAt/fxh8y3PUdCfZ953Qg76HnaF64iaX0T+Nbwq3YVR41nu9o+L/oFXkC7M/Y
jEQESKA+LR/PO7z59H4de6ITzi+z1j0HBedZ9ptZ4+E86g+tl5q7tafyz83igp+h
aqoNoQdwVVvCByWTLLjMutzvF7NoTxOGZNtZqiFt7fdQAuGSRlJ/4z/jJYfNJ9gr
ZbmmzpzU9GC5NPGblro31e6lZMVi4/Es0Pj9MrF1wFkJluT5SeONrCIljzK+IrQh
I/tkJCu6hgyadKpBUHj/+bAZHKtMLq8CMIUn9xomNlasR/uyZ5EedTgzY8krSIlY
csBh/G7I5iTQag+W7ofUhc4ZjE5+qoAb27RohDZ1FhZe2EEZoDp+gysdvuwn+UqI
Zo39QknFE9hZzfxPprLZGm0i52cwcSYZzQx1LOPqx75LWGQWi3bj9uVp5BotTN3K
miCvCpM4G+YYZ6RLvVzIKpUhpujTFbIyMHJfOBgygzCuB7dSp24oRj+C0qMwh0RL
fpRV3I01Kg4vXLnmLU+w64v8StR9PM5mnIqTPxiz8BBL1Z+H89ZmikImtmtvoZpH
i3JxQNm6kKijB3LmzwlsObFxb9nFzUBGwborXnHpHbAGyYB0rFvwgRZptHnLqBip
p0Vx0aERTEbqWVaN783oif3wgZ5Do4oD5pHSXvKc2c7exGntNtrnvkA74o+orU4q
H950xfBk9+mXnVs2+3G0PFYzwB1mI55ZrbRSDgWe/Ig8ZYvuxSn489XHyrFxMcam
G4JD1xzxMLvucAk+VI1luz3kxNUU9yh293IkPDOtpqYMX5nCpehKTN0XQzQPNQZY
bN0is3A1upBh/heMsVZX9H4IyzeMIjGIvDWzl3mVkqpVC/hUDIt+o9oEfiUrbGYz
MH3eK+cvpBHSV49FI44WZAshnUwo7m6yD/8dtIq22QM3+aprvHCnbSKB5SANgXE9
bH/VQmJzbVkWG0jEWe0Od7E7+hRA6MPaTAtvp6BspUpadDMbhkQb1a/P/RshQpdQ
FcsJmVcXCJnKuosI/8DcsTSuWCiVC2LpLGRJQLTkaJNm3QOttUHrt9EVx5lj1VJi
Ndeb6Pvyz2oQw+AcCLF0oxrsr6QTUsWQ3jw8o/cKHQytPLitQY3//5y7w8ejnzMC
RAsghlXhTCzXVncYHmBJw6Oj7DIp1Qz6gUHNjTcawnIuJNSd83OnU18lpNc9Ziwy
lnIBrhfp+JRSCzwf+NkH3/Lpvu+lUrjIMo7p3wzxFr85N2TBwf4Aj9sJmHI7LrYW
QaPi7JoLOV0ibJ/0ccaAC7a/1lcDfT89jgLZY6Xt5ldBwjv9Y/NV38mCaXaP1O8I
UXYgSNpBnFaX45B2iL1SfCDg46N2pe2YVaJD4/Y7klcEo7k/VQuW2vi0dxkJf3vT
hsfxIj6mKXE68h1PxuzrHf1zUeMVA8420OOyPbIrR06gAF5Lm8MuMPSyIfqNj6Cm
GTfCMwu7vejTueREu8l5wmT+zvS53/fSOvMilG9B77ygoNYgZWOeV5vn2c3qHM0M
O6mYgUX92NaxwRi+9SiBUcA/3dVnisJdHbCvVbR0fiqudGtlFH+0bpEHwIG2K/T7
1iy5OLlBU7imwR54Rb00z0Q5xigHtpVfLtForMyAtHrx23h08nCMvowLynOnAZvF
xKXyZ5JOmwwPtASP+VBgtAi54fBCrw+urdKHSMXBoDPpIGt0jA2E+hpuGsumuCAr
FVxR18TyQmbL5Kx7E9oVHkFEPBC9Myod2AK1DHCw2SekTLMVEs9a99/Tg+9I8ze2
WRAfT/aShNjKNlJQct42dcKs+cpfzDISMcwJ5AJmQnYuqBJ0DxWS9eXwEAyV/fk+
/+WgcrsIpsWvvpeq1aCziw6JNTxmruhGZzkHw5aTuaes2sHDKxJj9d4/gDEkxE3x
bu8iqk+8WYudp+xiWpYDwOHVDq8aCLww/g4lY053O8JC5MV1sxH3m8s9uKDqCXS6
nUU3qWBSuWy+bSf4I0ms0+iMSU/v2/okM0avq62YDJtiw/psVSyiHkxY0p8fdsCt
7mHGZ1/B8kh3B98fnxVcGIihvzHIiyaKw7HVAdrWaXMGfgzOY89CA/Ppgtyj/tpC
+5eGMWbHLB8h4BbSJgotccnuiw7T5iC8nj1PLsUUtD85Dy4NTGNqov1OXqikxNcx
ibyRG6sm1193s/pB7tJNx/+yoiEq1ch8ZWzsM197iK7KDCiClRhQpkTRtFkrueTl
jNxaDJUREreNv/U7Hx6heUDUOq6iMjf+CM1ul88OpVfDpYdVnYuQL15tSNayUX7m
MURZzP5ReD4EVw790KbbKN3CukZFt15XgbjVemhKGUMUR5DYhnYBGka8otT7uYyk
8APTFFMXKbCyRhFxCacLdOo6rku5fnIHWI0Zeg3XGsQWsNBK1X/Z6Ypfn/PED8G3
FrMlLnmbYyQCEK/LUydir1Ze/8sdcbKxtKZDv2iB2sUhWLSAbcVZAvYo6MFN+Y5l
VQoT5+UxIExby30LzLgxkQeBC58GkI0sIJPyIZLiYfsrYo8mKTje0NX0D27mvhEs
hT5rCwV/Lfw5D0tfvM/mn508dKePiCjDWtXgPsgpGnp2yA5jUx6WO2XEhqNbPMoy
qk3yw3E2So/vK4FoEvxsmtuk0jD/GT5icJkMqJl2LGPmGrwl2+gn1OQkA9gQL4n3
/XARtkiNiBAlHRSTlO6PaC9Ps5F2K/QmHHKB9x8qQFqvMrV9TBozVLZ79EBVJbtt
r7ReCCdXggdXW1ExMN5X4DytLXlUdF7m2jikOGvMePi7oMfNFLpbaY95G8O75rHj
ErVKblUvYwUFbZUHdIuDTN/Mi5+I4dVRN1j3WwAtjCSOII7Lo+ek3xMAoca04U90
jlvE0ZCsE6/NqrG6L295L1Eu8Bu5RRK/dK2pJ9KWBhaXYPBBQYTq9zAxMBC2m08N
Z8vFXoQ3V7gs1zj3vHUZMt8hPwEIthyliWOxjV5mqziKXHY75Rw2MD9GskYrEfNr
a/gEkP83o2kW+32P4bIGiJa6Bl+H5WWz0RyPtazBPQ7Y5oda9DojgrPUR3LZxCAp
h47C2yl8UCETQdbn1MjLSBfO/1J67BPwO9zoVgZv9+O7NsQxO3FZUrdR1V45P66r
2zxd9WuZ4xtpatOx6cNXn7ypchsAhZSUvZd5YKTstZ3TG805CrD7JxVhlekJ/fbm
JNrwUZwJ1r2sO+5jLjQCScGcTIfhMmRHor+3dNEZv/os0YIsfLK6p9AX3oLCOyJ+
6uUZJxlVa9B1RFYt64EWPluQKlv5KwxTxvrv/HIU3Hmsrb1l5LNSe4VQWf7dwrHW
iPOb+wb8CWrYZuZdLfjm+yhgfpjzmaEbZbXWGV1dTasq4j1UHQvQCRKZHO8zuTmE
RNPx54srcQ+izEYwabkGWETvHid7q4jZFM2fORR3NyRiR+GLAeI09PC1ZUL1iOpf
inFLvjmnzjvVf8ZLUf+dmomRU9vS3NCXbbKGr+e14/8wR4WhQcwnrrYTYcSJeNoW
mo8nmtUqZnEsJmPld/9Vbp1NzIgcE8FrGLKpn2BczIMpRCxPGNFj1l4CyuG1mPgu
IXNCI6PsnHbfVoXeTTBIdlyS0bKKITKVr4FZh++LhSrvl6d2EPyDvCfpqKpC8SKs
cnvAGQwA4u0zJZkEHJGvAYFOjoU03rznSs2ZrRStWnk8pDGvyeyc8q7syx76Joy4
Iw4p8z1fs/oY0qS9nvdLD3jLdYmdSnbPHqqynX4QrbO9bYDw7oGv82yTmapccuSK
B2FFJQikWIvd4pE/R8W6MazjSMJ+J82VJnEJdc5j3lUq60PmjnEDhF8TQ6Iaqtxp
J3xZdK2Gpd/1ICM+dMQcv/T0DMqMPTEY4l9j045CKpwkI1UHEYJSJhWhEwM6PS+l
nlJHPlNHRF4i9K6DY6Q47S/zCY6buQMy8xih6AK1jb18hG3Tort+Z5EPhaoB1YWr
gHQIw0YHqn2GQO7Qo7TvYm3o3NGj0BqJWbbuEerVIEvFb9fA9xe9wUEFXfot/9UH
jO3FtwhegiWtBUphiIsGvZdzHwfZR7x3RIrBfuDk0jGpq6qVIWb6UqGK2OWpD5fV
Q8j1BIgBGHFGuNvUzrgB8bPMDxTKy6+nAp3ZNrOPtPRbNQfONxEj3TILBjXDllpU
AIsHlLFrfGEJTFEaVuY5QxQTUrRWparhdMAKlkCWvXUu+b50B96QxQ9NL0Fh17MH
nK4rYbGg4/IAmwnmWvl/kHNsdhvjZnqmhhb6t5Lok2BR/+InMQrMI5hBMbZejinl
KwAaD9X59Caa5qDu4WdiLMV8+l9P+iWS6jBoP+NGW0XpBrnSbKqEQQgoc+8UyT7x
XPPcOaRSe35l8MgtMY8pnmdHTF7K+twyK/yslbJB5gVX+d2W+69+cLViE4C8mClK
X9skkqmzXHKI4G47kZuircwNAEmUmoQs0bKyxV9ZQLds0w7C1W1z98GKXkvpVmZX
Je9IqhtJnJYqzqFTRw+YMabWQGbmGn24PYVAsTtZZd2ZkDtGJi9kMOUVX0kC7bR3
MpkqdJ7BeaAEtZDIXia1anonKOCfH0Sn7g4ZyJdz4w3WayyO2CZ2cnwFhsfE6aNY
IPNc2Bv91f/OfAKYos06zpw659ScWC+LG849vufCQcy5INyjSVNSnyKQMsWVxvez
6JkKSoSzt12A1fR5eJPoFupXXclygdRoo0dj5VvQa+v6W3tlGceYxahtFqipD8Ha
q9RIDjMg3yFvosZ7iwTpYwhf6QavUCsZlVGXMzzcAAntkYKQP2Y7AEW/HPwcKync
tYwqBL5eZNEhqAG4SvPSZx/ENNz3RjILlvrftQ9iZtaVThEuhiYxDmtcaroRtzsJ
rtaiEYGeXyebr/t5o05S5WAYitYJEj4HmyGPCdtqSF7qkiaBXxmpeO1zw205O79M
lPtlOCObnJ4wKf+ypS/2yh2zIMhcOfM9O4h3al+Qq4A+Ohfc8Fj6pLvw+Jn5SOBK
6P39hRnoCA+WjJ7xzw7iOTPxJWGjMU+IUk6vaxnQdWQQ1LVg3pKn1YO5gHLzIp1d
lr9axxTqcg+SnGfqR4Y3IW5BHnkbf8XUPgR/fvAYQpJ9a0kYcrjkcnbbd8SjhCv0
0sWMlrHEmh0qhigMkxIRs0Ynh2XVVOEI3EOBeh++SpshLbGbPhh6TElzXUpgKYbF
lNpJUOOvVG44UyjeKHxcrt64corDyGKBpjAzwvy/sD/hbGg2O5BXej0lEBe8KhSu
xvLYsZRL/py24VksaP6Zk9zLYSCJd/PX0xJWl02vCVXx08K0m5mzqYbM+SjxI/lX
gge2HD4M9Pzq1LwfK9qVz4VzYEi0pAL/TH7Qdid3h/2t+6H7l05V62ciRDVbKgzd
5ZsK4bOCR06KgXTpg49SyQA14f7ocWxFyEZTCzvX/inch0dxatBHtrmKYRgqTEU3
ap4LBKdsK6JTqmKMN7FCV8eU+wKaRmaHaGkD+yM8VYq9RFYzL7A6htf73L8WVgRv
PvS/h/FZvxFEgpTfxOTVdQZJgDr0fiKKlmhs59bFlwAR716BzdXI9ye0cQE9QwV1
KcxqFPlaMkHyEBD3EK272I5I/owtwdZFFBiXxNvSVFSKEdPynNd98/okw51E+s3q
bbmdeViakxCzNxk1FioJUxTYBPfxAflPcJABcaH2rLI2++1up4Ksf20HMChZqgP3
WNmadotxqt7TgBN/E1BLebGPh0NbRkVRXGrUYUsRJmcTKoPL24ecFRAeX8BwaGgD
l/L9RhC2GfTS6Y3vokuh662sbTwcvD40xbTJTY7D651FpLUorLyfjEHBue7LD/sH
zCIk0IXQXE99ZE2RrRp0PhcLhfy+CF9FWMUuSe9gbOgM8z+3ke5oyxXU5RApQUlf
bxQoHtrm0agywL1GiJ43VcfQUsM0L8syccu5L3OcWvk80mJfn+0UnoY0xY8fcDCo
PAHL1rqqfTmVgkOM36RdQ6IztPDcmc9lxqn87zBy+kJ681rVd2V/XUpRiHdvmypv
Bfht991SX+dA2aUxjxNbFGkP8NydjWF7nZ6rJpoa3gTMPBVNV+Ct+Hd6ILVV3WU6
h/HoY0PMicTNoirLGPDHAAmd7AI+G8yzh0YNherq5V0A9P4D4s7xZl1KCiJlaVUF
ugkYd4n1paKmneFoicZBd/FiDh3ueSGJrPYJPXSlSq3vdf2432sWFSaEvrzQYQgW
lrvhN2vn0VMSwMcw1Zmaw6mlyiLD6B3QfHOIBPWmYYG+RjQJ4vQ2fp+Pwjjg+QhK
IcCm6LqIdpZgXZ3nUyTB12IDFA9flP6FAa1Fntt/HsJKBYkIvuuLqHghavkvK46g
07TdtdVIpaAulgkgJ/Hi7j3/Ljyh9NCGG1dyRoeHarb48cDDQfFulwr////hyNK1
mfD6F8FAvNjdOdbHiQOeIt/7c6lqYCNJe6LDfDQ42ScUk8YPMJGpkcGsIRP3m5Cf
vl0YBE9zhJYgF0GRPAJPq/kjdZKs7yocsNubHNXzaDEHHWiGGlUYxyQYeshdFIKb
MewjNUwaBrA79iUOFfP/3Xo485liUzuGEABw1CWfLeLdjJ9uVDvIMRZ6EnbW0qqj
duktX+4S+cZTR6Jk+VcAthXnLbVOUjrBuWM7qZfgr1GyND6bOF3jD6cPVAMEF9Mr
KF3C+pW8HSsKDdX/YYl741JSdsuJDNcPR1TDjXpHh++64GQFZygVaCIvdwyT/D/5
GUCotpSd31WgFCyJYDV2HYRjr8v1czBcd527cTAAz1s3TcAvwo6d+pnofiwAPzTY
tmOCof2yfsCNroozd05CBEKnkmjL82DebNVEw2UY/XwNThxHrcVHO0vMXQsPhSL9
SW5V+SpAsNmAWdkg6W36p3Jx+Wr6gwnpBZvQEhiKBgLWAKT/Xks5zVDxezQiPFJW
RNokcalSZivegOuQg4pFDozjD4ftaYDi7CBTIFkwOG5M6/5qFMyjKIMlYGo6f952
M99OQCipp6ByLihCyuz40QpnE35dh2WCdNLPE+YBva8N2got7pSbW4TSUrIajJ5+
BFoxuWSKhq+th2XMTt9kBe09wqb3R90LEMyc4w9YZAFooIgxhBViQCHAk3N44xMr
l0oOTa5SsjSEiDlgBB++FMxr+xvaRKrVWxYUD7bwJsVx5Faewon1Nn4GrSTd7PYy
EQpqAnlUeyZOo71VATKaZZfSEfa9/z3ina0GSeN62Vl+pqiHO7+VKSxgu75cm+Y5
sW4wViwjg+rD7wnnys6EgpSkyGQP4fUa3O17jYrjgb+PSlDtEv8Bmg8sZKJwR6yn
NpXQYHycHxCCE0ZaNwRlte31WIq61qaDrgiJvyMdbirnAWVSpwAapiEZ3XM6Cpdd
iHz6zpl8P8ogauxLVvGJJhY70IY3Oa66lJEMJQRnENhUV4nubJLXm04kkJ/JcopD
73QTQcLXQ1jDmVo93vH39h3CUHXPWv4uh6qr9Fr80vs6NymeyVC68uFWi9uoUAih
uyloFGwhGOwIiSrxEZ6yQkIpsXKmhr03lM+KTqAU32XYGnzPvvzroXaemOeDdrql
nndV6ZyT1dp9cRpuriUGG5ME1ZA30FkR3uOtn+VwrB0GbUvCjdOtexm6q+MlHDsb
ItW9JupfhWOQY3BQkiujDS7ig4OF8aFQU2s4JcgK2EUaXkIK896sFANQ8cFLkv1i
rd5eBblDhSh06MFKhDXQyj60dcE8fkbQDpI1ReV5JJiNUR6K8hwY+RbkTnJz8sZT
yybsKlWK0RIYd6YMCw023cgYYiBB7eGd2wcnyqWuFNatNGGNQQVjnx5JeGw56zMj
JiRy4Xk0COjLg9mOOBHPZHjK7n+hf+nTxTNGcD1nPWit7a5KgScjh2KabqmDrbp5
waJvqDZ1pG5JzpcF//3aEb4NGi6GuMuZvEZXBVxJuzPJvMGc+99BddBlTpEMGXoE
p9JwMt4MJhMBJmADsrZ5qQenTxaI9pELPFDl4xK1V1epw+r4SRLiwrFijCkVh98v
9NO/H8ew4zWG44zopcH3A/A0/XBDnPkMWmGjA7EGHbIYxMTgLKDBej2+f6s1n9jf
QijBAUS1qf4BNxMBSV/lNbDgenkD8nyDqzAROqT3kXX59zBoacsY2y1Ofrff5AW9
D2t5uiii6YBTVEr3S4zVN4I4ZeUCxNVUAiIP6gmKVfO21nx+g41wWyqQMjLflr10
BrEiq2XxFfGJFfOTZWFAJJwgoMNyzxDlLsGXw1HIck3ft9T4hsNtuEE70mox5cQ1
P7g7g8zSuaj32jXU/CFgnz6tQCW5twF2bf8FJ5xp0YpE8nSY2zesV376vOlPMxRq
yrQV9wNOCR+gKVYzTpWTB7OroYQNOv2zKC60wMg98Kp2SSlFfaXpHAExCQYQgkjl
/FwEbcsanZQdUHWqeVGfCZN/cY1xin3fx48N5iOxT6Zz1M2nhqvDdfHruVHx1ela
7u8j5oY2lgleZroQE9TZURP267X1BHjInTG3sIadJJ5AoeSrPjAoJM93+tfOtTbx
/ZRu0Z4jYtHnW5rc3OyaAjaMIPW9CUjbb7ywLC4dJ43J1kjLAuBzfOAiSE16mh+T
lKSYy52D3d0HvtR7Lu4OsShfeYdYBBUC1XF+nLo443ZEGNuwfqNCTc3pgU/AuHdn
AJZvOm2brP/vAR7hdxklm/dOdyHJ7YQAB4JhW+PMP//2+xC8or224OfYz9dMx37P
a09nZHRTb7Lq4LBSaW0wfjlyK4qFO28LY7JOZEp8+K5m96Uh/tvX0qExQLnEHzNu
gZ3NgCcnJE3p+FKWGxCLsKKDlbf/01MsPRDO+/bkXXKhqF//oa2e4e/Xo2fCzQRZ
fbFt5HkdwLS96bHSPEytUoD43QCwzwrME/4sWzRQ63mslXRlczjCatNn2dWogYuw
H0ZWCcA3E/stJ0bJ08Lzsvc5qf6MZLxxtZMQYj6/TPWoB1a/5Gwd/PdzFYw0tQUr
X1FyYnE7Vvd3P+Vo1HXhOypgwZh0IJEV8NguAjJMPpDf99qhT1bPZQj7NgSC5lLS
bvjS+gNfDwmZ3biFsl8gKQUFq/1wsu8hxPxn24itcVkhJdaja9WdjMKKkaCw8VtL
eV/LhC5bDtMGIeaPse4ZApj1saW3jboGgnAllERfXft222fRRm0ucdRUhldPg+QC
9Z1IgBWGRN/SvDUDrpDzS/WS74rGbre81mXGOijZflllW/2151rz7yAJ+AKculko
TdBMWNzHQ7idK6MDaXfv6xNwafY9OVPdHp9GmYt5Ow0DxotspFQePVfU1CYCM6Nq
KU6foxv9NvFrkMQcieCozmeftp2NfHl+8vDCsxLIv448MBWthiUdUG385+2R+iGm
lC1xNhwjQxYMYkjFyLB2C7+L2DxcGPOrKcJ+qKmZm0Q9BBqZlotEtTzp3EDVyyHK
lH3EcxoMeOeTgavI90hf/a020Osd4pD3t8lFyjLi2yTlp69tKcA2YAnjNTVVs4GY
VCP86d2JCC4lEhxGKurqajEYhAdzCDcgwLMbzFa1R5KsPNkqe5AiuJyxOnZzzOwN
5YJhySFWupEYbr71JRMrJpr5qH0L+ZVlF40IJ5PqVQapZgn3d1jZwNUF+/EwGmXB
HljBh/Ed7FkrVjMwkBaxMUwbRmNHJWb6tf21eG1yJhes/OVH1FTofA3t4WJXy9Pt
IRNRw7WK5S4ak89JvnF3RFVB04l3JBlWqVvhHsIfp9Kvnw2VvkU0+NwBcAbh79ke
V3cWxbsGtNkpuWlhUmcgoB2Cketbl/D5JvGLpiJzsOauBwEJxnjonoAYLBfjfpUZ
Z1sgvCzy6dAXKfV9/dI1Omuyqs3saP95ewLAusJVCKmRc5QPXFnKM2BtNpNiRDLW
uFk8f+ugyFFwG1D966KRL1BjMmnTJZy4l7YDT55rIQh/bN67V1LsMw0o1StNnW2H
WqHHuO00UsO5jmSqN1veICntnyJcblgrrccz8jg2dtwA8I+JsqY0rJHydv4+MUo0
xUAf67Kyv2/xGgGXasyR4Cc2gMKR3KK96Z2kGIUJy9SxKaH+X+K8D7C+FRgMWQ3S
Rh9UgJU0ecYxp/Wc9hEJMf4R/AHucmimvAky/4dcJRUOBK91n8zAPpAeQrhtp83k
kh6bGtL9g8pH6UzX+B1rtS9yip6BfTkTN6ek2YMFZ4Jo9EbIlWCD8imzAAXO/22f
RDQDvp4fjji6somYgKv/uOnuGH5jEIPfc5ewLpfFXJDg3yT5xlM07rgYFt78EDVn
W1bX5n0v0UxE3wLoJ5OuymuPCkQT84Fn2EpdZJ9u2Wh/XwC+bedH8nIb8DIZL1g4
suukHlQWIhrRY/KWWDb9vGhmo1Q4qXKB/fpZP6kOeIeUJpBblHJrgqSgrppR44Tg
Zwrx33UBBo3nHvrw6JBSNylceeI18k3rj4EX5ROQud9oO1/JuSe86rYiKXjHFjqj
tYWGhpV/U/6PUskFdIE2dSxT1UH1jz3h3cOJpu2jjoPio8dl4/LxNq0NBSSz/llr
QC0VJEc9ydDuDTW0BFdy/4HGL8qjF/S+AP4niz2ec9Wp/L5kUp8+N9UKgsV3oVFU
hG5SQ7zYNgb3m4Evz4SXFhcgnwe+DWJenOkLUBHKZmzfcKTucP7cwmsg0yAfzpt6
598UVBCFZmN8oELwgoWFDeEVZJst3v8eJdmbm/osd/uQgKbiezk+1GPp5GVM+2Tz
iq8zzgNcKr3NXuf8zTPy5eGWMNoYsyIymIQvPkpp6qzKJpFeq/VjE1IL+4RD4TaW
17F5tBT/rxkVoy0aGda8deQ/qvblb5baByo3GeokZXAnjZNwGHEGY/L1WA+V1H6i
Wztr9bldWslbL5mJMV65e4UXNAABYrxgfTeyaXJML0cMttoQDaHp227WQvQnpieN
Xbbpy7qj27V6A1FuaZTTSZg6EUDogoJCnefQ6yvP0IQuliur0kQT2lbNdTRun3V7
mDaz+3MIo7aQyutuK9daer/SFmKIyysSwUayOwkyBRTwtWXTr2JzrhM9t4Hw74rc
3PZVN2Z5ijSvaqwQP8W09NCdgcRkwVzzud3wftuCN5mi4obkcc6ee1irgKtEA8QY
AcWzq8vq/SIZZS8GCVrEyfu2t+uEjP9O+FrHSkAID+McHQdhq3iWTdQHHQCGlRtD
E+Q0f5tDT2ZLtUqSw2jQYtJaC7F6Qn5McbN0XvIjzh26W2meeJO3mlrr7NerW0N+
fR/keeVIl8VOShP4F+1eCWhgxNeXeHhK0+Qct0sLb5TSoyyAGwVKHJ+dYsuJeTxT
6lAbwVi5HvP3Jib71rDBH4+o++aG3niTjdPKHFvIbkpBYAnt5rfPxpzHkBhRKk+L
0FyWf8gndAeJ4wz+2dxQyx84O7BTAa4dQeqVsBvscQ6h8n3YhtTFk+JE+gZE/VO8
iC+XdkX8rJpx+IKIZVn/gCQXAdQIFVqSl+B2T1k0Vsgp1Wset6WOxTzmB+KqW020
n95cPPbxiLG9Q5/NT4wu3UtjNUzKYSm0vQUU9fQOSuYglddje/OQ3ujuTQx6kwes
V0+HCECVZraokOxknTDFmg5+kZmgjhvM7nf6Hrw9asAWwQ623J1g5DYqTdzI6JXt
vMyKmO8+xYvYneIwajUOOtUaofLN1edqR5jrDlAJJXI+PEcwYA9hwVszBgv72kKo
CvixZQ1AMOvJohkGV4o95WJlWxmK4nhTWe1lDKp4XUiHRvK/Iz2WhPv/o7Le43qT
M66iLSATXunMQN7ne4pHpd2dofQBBU5wNtbyhX8z/pLJCcsqn4zNyAZUjMGrsLBm
CqXYKo7BEGjkElDOgWZhCZS0FhxvybkfbFd1Et3VmszM1o1JxIy4nrfqA6LvaNIz
2ChHNQzMM/yvZxEpWJE0/aeiSBkJP9EaC2ZrnvCbxr975QqeObFMrrWUyy2sLM/x
HQXcs8kg0AVSrOqSiCK3JZrncyBL0RBYf4Ai9Y6vzpUQJi2hCsxJLHuCim19LMai
8W2wqMJsWrvygidpMfRZ3GHq13qduPsCjVJRY2tif+IdBurpM+SNzxnkzDMtHyRh
25zQD/oXuMkP2ahFRGyh7i7+LFfxaViLurEVQ99zFe3FyV58BNLhQczFNfhAhpIl
9TtKj5kNOfT93HdXUx9pf9w9lA7d4RPtUHIwudr/z9omKuEvfCJ+7h7vxTpkqFQs
Cwqp9mSObC/I19Ir6zswAlJPVZodVAp1lzEQdozH5A6wrb3iMbWTblue+pwrQ61Y
OsmAitCfDmNtzmQIhLJiGZlSeNtPjg1ucPC3Jn2wnW8JMjm2Fw0znyU9Z2MT7vfy
OWrotQYrizi1ZJ+empJWaHpppJl3104RitwUg8noufE05syPy2O/Vtp4jDWLUUPG
2ZyCu30km/AQfiUKmwwlLeMnN6azyqpm6ttnUQ7v7APVH8fBtdEagdL1nFZSWKMe
kctLpaHOL1ByPcJ5WI2dQjY4XOWLszwI1eVxHRiX3y2KuuzOwivkDAcxdIMysSeJ
pYooBY+9b+2GXLz2vSWKWJXBn06IfHo4H6UKrwPzI8BT8CasBBF1J1oI6a+s1yWt
LmIqMl8Ns33DpIeNVQkAklifch7zN9MyOIdvM3aGvbBeyS4Co47jFDj6mArlxIDV
B5+pr28e7uQINn/ok9tCDzM/QPCkMMa1BBrp00cbkECTmIUVaFPDCsUtTFDXyYG2
D0g0ngMe/JJy6D8OzLAvscgkk5jH9+0aX3L6ywEMmq7YPnS/R7kCriHfptlUvRCM
YIk7a38UKB6m6mwfLmi5fBUDK30y9rMux0a5mNMMIIr5msUebLlkj9jwE2lCVL+2
lzBJYYyM9g+e7WMNkL10zXmn3udZDd+JxLbJ2q5STmUKPsDm9vDWQYGlWiw3BvOE
NA1eA9wllfdf+xo9LH5GgbhsWcVhPL6Q0usxxAjk1tBLZiUI6svlDqnGkZF6bt41
F+f3r66YvBWXRQu4EXDlNOPVa7Tf4paqaIZ6YfG6nB55YuEBXKTNXVXQ1dgbvVl3
OjJfr9p0TM2L5MBR+/u/7G9eoIAUv0AkvukRiK5Se/sfHli5dtqbT11XSRRs+pYW
nkEcjJADGyssdnSNvrV/lBp3k7DIFobJ5/TkZV9szkl9UBczF3EGxEr8QqtPK5Sx
iozQuwxf0IqG4LP2NYMIQ0+flyWssHUn1IkcTB7/Rhc3XtSjFMBA1bGORPR4g27T
t43wjJnN8gytOwFQXaelDeGbI4uL4tlepyvG9UU/uhChywi5iJbbEzQvrVoWC15X
Q+yYjaDqWe8p37YLinOYC5aXhQgPfPErcihTgZ03PXn51C5XPjXT+H+LPkATEvx+
OepTvdEqlTafMnGxqR78Qh8stOpkBUSFK/q8bdoUvjCSLg6tQP+GVVcYpcQEFR6n
bfEQ8ii6+jsoLvVWKrdsqUnRHbfJfkO3DXbd/nCjNCZXA7mU9VisW3LJOLlxoSkd
FjZF+U9p4VSEJ0vkZEZ4PjPm29tMrvvnjGSQrykOmGyzGMgipFVgAZPf5/WZPwGJ
uBI8YdkKP1Kx12+6GzoeuAdvTDpwd/vrrQOI+pamsGw7E0NknTz6/9mMcOQKerAV
yZ+V14qx2+989qYpaoo8B6xZp5lJNXR2wDcipmu8aSVFe9zZcl1EP6t70fyL/poi
hE7OGL6KHiXuVc4/M7V95o2hP09T9j6SW7CXHfH8MMRiGFVEfltgZFIqn4IHcWUd
BeK29Ywm2fV92VFaVN8LB1JecZ6P5+xHWqgyu4uMXQy1g/59zS11SjQq1ty82n5g
HUXM5pqeYndlIEnVRYZpLWYAcnTEC1W28+QC31Kd60xLhIi31eRXJks2Bbq+2qp+
oSI3CyEeZLYM4XMkeLih/Sv2DjWgBpBmCSq4jQxpZPUy0qrYzR/lcVSy+ryDI5x+
gVHpYMnaXR0ZIcqBVBqHTNG/ZyFRMET1AdtoXgLWv7YtM16YqwMgixADODql7x1g
7hwsSyvh7L/lLyp0LAB1Jri3AMnoLU9qUrDJm0G6RS0Wa4Gqb2kUBPIKqZpVawY7
UAhZ4zAKhTInsiYs8eebmYkfUbTvN9I0jagU50k5Y0eBeve2ITJElRNfa1bj+lDI
I+UwlfRZoOdqPoKlXLkhwDyjQ/eCp+Auo7DcDJMfQf7Fr62oOBW9muoGvH21W3Ej
ELQjZD1CzY+WYiD6i/oxlyJkAuBUzHvz3BGJOj90LVSKBkqqoV4u9cC9f1wTcEH+
r+IxBXo9MUiaXLCOcMgYQ2aONN1+ZyFyWpsQfbSy1LwjS3eO37s5AFTorhA9GQG1
Ixq6BczASQ2I5z0vZv6df1UbyeccdX9JqX4sNVJ5ekJJTAlyGIcl5f0LUA+yKdNK
o2xYRzxGj0ttq9zejnjB8FW7G0RlevI/yR2yK94tOwJoci01dgUcEE6nIMj2KHE1
FT4EzqR+CuA6ac6l7BkRoq+J//02evo6kiqbLhMNrHRrmu9mU+HMM2BrIUm9er02
ntquRNWvsLHjtuAj2dEmURAt9MaVnRdAhTMY4tP0nI8A9avaikvUQ/wdKJ4bWu04
JUN2eMZkCVA6wHhTpIc75wFlPuPdNeAS0GTXFoobh1feR0kYLKJWXQoFA/8v5TZp
oYoiN2oJLlieVhnm8VDSl8S1uU/zBQJ3X0RAq12r4KfslHXYkPRhdEEQz3TIlZUR
HgxwizXmg1wuTvT3+z3JnNCmMrJ59vCXOtotsCEl1r+IaUXLgw43hx/XWW8SUgzB
cPzibBt9bHbxDSxFbD7VZ9nrjchL1BIDJQRLGgaGVbQudeRcIn4JF4ku+9lwq8qW
YiKsUj9HBIgfKp6AfcXGSA5vAikt3Uhf96n7FlVFNChFe81DFPXhdN9eXTJT1aCa
ljV+h7jw05sjQ6BarM1VEKrdsqXK7q00HmuXV8pnaymqiyGfFM4BogbpXT6VxO4I
KAVSHm3mYGBPvAquny3LVhDbRzE0DEfDMIWkXru1Mc9JHqoUnz/I0jqNync8WCjp
5h6mLk3gMxZQc3xh1sMec4/WNuhdre3v7GBgmbMU85lF9+i5GmOMrllJLzLrVWyR
k9SlgHBssnbS1CEE8ZeZdlrRITdiN+EQIE26xpqs33+l5CPbulEZOsVvW3WkuFWV
6p0MZqR7GuG8MxbBxVr5y8qyeb3zXHLQyXHKoZUGdxHa0CNY2xfUM7B7iwMFWhjU
l3cnqVWlV1RoXhFbQHl2qSlz/2KeDvO0VjXbsUywj4GXnFn7LAcd/gPMZL8pBaTz
d1PMHXCo9xdQsBsrIGImAfiEAMVaSvjEbKqmdHrfEzh3Q+1zBRNMrfAWdUamk43r
5cxa3J9o/nWa760zu252gvXjOq0N3mnpUchBjr+DprrRm4Q/mYDbvKGw2PoAVjAi
1wdtA/xt0E9ZU+oqWsAOkOLDhBBK7FY2jW90vekag5E39F0N/t4YIelq0G3K91+U
6X7G4dZMmudU4gOcUhkSjueCiQ7Vx5YWmsUH09JHCt0jDaCOLmotqMOtezLgPpGZ
gKbcYOFoIRtzJaDZuxyy2USvMLdidb/HsSg0oBwnPN6lYJvVaenU8Mnc9tktm2wH
QjNrkOs24ck3NtKyKdXdKA6tzvOXoS9Ph66/j6YeARCv2syN1jZ1RiMYeolwwAMB
hugK6ZrCX9B24FPDGwh85NaTPyLlUvKO0Ek2bJxmqfIzQMBqwsfSAU8iZOoW1hzk
mi7A9RU3USYbCOEXfk6diU9EU3TuU8zf/gOOIt9/1pOwCkmqkTZWMgncK4uOY04F
9lX15m5rzMlMA1qMuj+qdbcclq4ieDPX97vo1LQdUYBokcfuB/Nj3qpM/ASyzHbP
5tPTixO/lshXTBMvqmlVFoiF/r85egoI71GWb+0PXnvdW0sB3yXnPOamf4tjZOzQ
9IQUKoJNkdCuAPbaMFw+w4iK9biRlOQpD9hLgsWOhh0v60kJgOFZCPKRfUUShl2H
qV+2O5eA4hRa47Pa5gAhh50+EA1oTBAvRpnbsuXlZM8ks+REOvqPIoGdNNZg0IGM
deDaysP1mH8Gx3hI7KwAPPgDAfMWYONAOrhMZhCFMXmeefyWfDG5vxAiM7ziFaUf
bF+rRaK0JRKqlokKyO0XCQhgieIfd1lKTqsl0cy4aTAXIET9RZEGPounWyGMqlsh
RIWLKl9plpBLNj4PbKh9O0X6b83FuGZ8rgD9z6IdbRxlsj0PDYO5jsPtmAZaDrib
ANu5SqKk3nWcjLCGO1G8lAQ3UrDYrOHukphHC9kQ74PykhCd5sadHsBRkhKuZr+T
t/dTeffxEGQfTSxwcNwpjKmXMvPRlm0C2qmkDShu1d8caMoDwtGIrWrmA5R1S12d
idfdVex4wW6GcdDMgucDkXEUl7ffzc/u/tHb1bkjA1tA7nzSa2WwcLqTNHe8lMwr
3e0zlWYmZZSIe0VJoh+kjXaWoMbN/Q7pHTtNGK6e4Ni1iYWo7Josy5g4WPzBzR3T
97NzjizL3ZNawCndAcl5fyEoXIobTqb+JkMRVdIp9DxBywLIK9obKAa8y5oYxXD7
icsSngChqoFQVhPYRTnjFwxkCJWSejfo0ntAOJ4KbiKOOSXnpsuleH6E3oWefhGJ
sQyyNIxU3RBkMs+qRQeB76iRi0fCtghCwln2wT7v3pHwkVSNtdHpHDJgm8Tw/98H
HFN30z+6TcZYTXUBQ2CW8MpCBQoOAjoNCzUR5C0sRcXmAmyc7XZpqgd/VPKCA3dX
BFv3Lmh1gnP7e0A+nLi2E6zWOChvzussxXSLXaGmAFaO2s+vsXBV+iXzvfo1RgcT
kzJXOfjIRjIl6Y31EYMULAzha17YpkkLjSeAghcJIE8W9ZWXuH4eZmuH1lcRrV7U
kiVPC8zBmyyrj9rbtYV7MysrU2BHJGq0dwFLtgSnvadHoOy/I7UF/rUp0CIaR+rO
Po6GXyOkAauISPgFj5qN69bZR5SGHpT57nEG70WmlUWtLzPeDRam4VRAZrg0jJ54
TQDtM8+9Oc2GOS+RKee1e1J8tmejphCW3T6Q7+4IhWrUmyT+TEMq3U7QQ/BqG6DK
jEEH5SGikj2p4d7EfL4jBnzbjTPljfp+uMRqnLUv9FF42LiXKU4iS4wQhiuMgAjX
qZmFlhwKBUugAU8AXybDG9iuIcjWDG0Zqkkj6KgmYuRKUqokRib/vhrLYy7abwno
WVDsQB1qFeh0qSrx/IQ0QbF0j+XduFc6eD7mkKTmDM4AqZTHhXTBHL10CEGXMxzm
Sm1KhVCuVtY4jZ1pMVrSYI2PhW1mwoQ0+X2TdfR4q0rbV8k3XJyTODfbRIBbH+S9
KzcHw1TjJ8VycbMXiiFgrMafVLQw3LWWN/b3HHXx615kYD6pJwbm9obVplXQ53yK
duo42wSbFpGH5kqzuAboXgnUEpylUwMIKviz9LpO05IPZ5XAf0NYzbfYVd9fkMkO
5hBa/E9Wkz1zGfxwI77kXo+wXYw2rYZ4nyziljlUsi5lfxUpnJfX9fI573jMSkpy
8lyTlvPGZDiEaQT0TuqvQpEMsg57PCUXmz9e0vbCOLg4wqreaU5bvNJlkW6VpJTM
VoMcp6iofd+w9IQZUvXnHbu1NgZsqTsmuns8nyoFfWrMQeqJ8e5zBVwNh+NRa6+0
0vhg8fFuoAkN3GTyD2L/LuGoZ1h3uhhc3BxyX/hiim52+3lK4i6FQC2i5G68Q98w
nnOItDk3stT7DvsWUYBtXWJkF1lyFgPeAzH08Cqmp6zSgpXxDHuu7kCteRwjYZVQ
QYc/DwB4v3mERX36+tmu+kMne5hifGwRj/WYohkHNhNL4bMCf0sf7slWnUAJkzwn
sECxmdTdAXWFXGpI92yJ13qLFFa+n6cDnNN/jlQbKHBDnG/RECZhsQMotkR/UIlN
Hj+GVJhgrizbAiRusZFxbZabynAOfP+T5BpDIn3W/5+GDtl/V51/ADqagN3tvO0O
R3AKxgcEuCv4Zc07c/IHn4wRWjQQQ6a3R+yLpS327HAbHRptoAc4xZZUdMNMnjZv
dR2vggaWdwdr/nbudmtAc7OnzCa7QY3YKWysVNvcaud8lTukEsvm5FVv1FHowxjb
BfQq1/vqUlK8LrpxmG3hV/Q5WjB+FmXATJnLRqjsEo4A/k7751Geg9E7EZGYS905
Rp664zsNP1fqdl/TXRTTDqVefx45GRFAYp8F3Rdh+EtQmAnawvfw+qoH/NoM1Zw5
oudqhJs6diYasKexSAN6RZ6tMuEG3HEBBAkz2JmTHAhlq6FdkqMjsCw9UWPgNjnV
YrcoBw2CwEH0j6KJQ4RDnXKcWDN6eQtmHaXqiMK3BFklFhiCDnWJEMEiodN4ocwm
Ycb7WMM187jNtGQGMrXqyPogbaPpXtH3aPoToDdu8GF2BmC3w4L1OwS4iPfwB4Zc
8+SyQwdeOgL2V8MIVP+npPvYv8lwYU70eTgasc+5k3epkW/yhpUy4mtAu/eanCoJ
s2QASlu7qAJokicBb29mNy8L4GsJlgfe+GA7J6NRRV5FXMuJcmgtGz1FPIZQOri4
0GfE5ROcCZpKVFoxEAUlsMXP/JmnWu0Cl4wkjLJwUJ/ZupCjXtrM/0XROBFhGmwS
+C6WhnQ3x8L6mdemPNAQYhTedsHT7o/oNFN9p5GBhUqofWUPgaFMV2mUHbJaD3bI
U8E5GT0qRT2jQlkYRHgVwqjks403Vyzq+zGiks2VPEVTxY3gPzzyEs5XsBtUMroI
EVdcOW8r8dIknRdb/ORSRO2Rz2pDW0Gt9iJQLDMW5vK1mbOs9RMHcqCDcIazzxKD
8UHQX0uXPlPbUEV9IFs5V2FghdkBZcIzhmyUCowvCuIgC+tbQId1jOD1/WMlkZ8T
eLow8mPIKZ6C/sBsvmPGQ7Bezal25t3LFmjsWiUdu2mf3wJDp5HIiGDpe19APayR
PSbSGU9SpATuVEpI87aRU5OYxADFUSefZ3G9K40rOqT0k6rOWuH+8b6o/U8x4hUy
DiZFzmx74VsiH1RFClIqKrVlnX3QizQFArpwDdOawIBYTBoMWLGxi0ubcyYoQUC2
TUAeI/nD9Du+GNPL3iuiFzT8CjzO1HJTBK/+EFEU2E8rS9v640QpVJzPtptfyANd
IhPm4W1kIMaW1y5KvfnHbhx+aqx0M2B/ZSB1b7hF5xhZyeeYwn0/waGVLje0gRFy
eaW7na2u4N2LG4mAJeW9+vpKNKZke0BPJ4yRjM5ZJnw4v2XrAozyM8LkBC4YUiom
bmJNeenMD+M7LBpsrxQm9qzMjXcUz1RjR2lwE1ZJ4Zhd6L+IxxGubz3/I6mYaBRL
hHVMdttMRncSbmr1YTLINFvQxcaeLNwk1Pq1EZCbL9hXQ98lZ+YHLuxO3XDjw7ZU
YgJ/VE3ojK94BZi80ISO1MI5WdM5JPTNDsiYk/ADvQph4PqxzZjX/TQ0uCXZfZto
Imo4wGMD6p0RYIhKsF+TGrc6vsrio1gx9a4JdygcSERTcIfnzWxz7KpSmJ+ACN2R
x2pXBAvZdiURpkVL57w7nzl8NbyTubDoie/Yn/ANZsxhCsZqm0lUhYUK/yIgWD1i
1RkNwrjsE6xLEMPA1/21uIudnZ97v7SOErTXQMHPCq52G3d8VAL9kBZyT7+6WSFa
96LmiiV9ZjOOYHwgunbmn5g3WdFMIVz4E4gXKQK915tG+tX9SPQC3NRDONo18T6T
LTi/VacpKLC4IdHfgcwbYgyGl7T2DrgO3qDm1ImAubcOhNnRwL2RQnDMcuoEUuCk
+uADyEKh0jhIH59BFNfAygY+j+NsCYB8xIKOJGwehXBgWeOSXoh5toPx8PNw7HZT
tnlO5f0e+PGlLXhiVFxe10W+0ocxmMaKqTsZFPeWOI+2VUnGM2G06nUFC0okGXQV
Fwn2ZNuj8sVRqY6Vv9dA0QM/8dXpi8gNAIiky4EpCUphZCApmEFtD9x4ZAeIVKfE
UpyOui5ax/QyUFUil2VKPce9Ht48HbXeBif40E5/+D0TRB3We+98tTjyfMg+cBIh
jBo2NOjcv3OjNQwFm5zUxUiTwYYS0H0kHYUq9IKZ2HeoeF33iWR/DU/wNO12dHx3
fwAWcvRaMmV19HPyYnkX0j7/OiQnrbV+P5PYLyS/UWAwPhdGlEeW/ZQhB9548M/x
q1L0y6WqRq00bUHV/cBsVI7PCZRJ64f6EYcPGo2BNmjWYoqLfHkTXRnS+YztBO1P
XSUGI/vbGR1YNZ7fEUpN23rV+lNdbQtuiIlUTOcyZVk1er006mOFTjQ+qbM6x4ua
KdxlYZ7KwdgtY+Qg7bbH53pUithehzDsuaFDmutlzGgJp1UAwHGFwGtircDHXW7q
XOaFO+VXroWDU67mCR/hzuGtEsowjEBbNjfAFBOs1x2qdYXQE2p+C822fQ5Xa5ME
nN8kz4yrEjduy6/GaVLZESqwMUZOELfRTpUZuwwu2I/HDIf1RAhyv61U3Rnd8Wz4
XKlU+ivBWYY3+FjOQRuSTTa01wPVwojHm1TWNqYhnKuLOUEajOLNkcm1WRVmUnki
iZE0JPjbgZLQCt7AtCeR9BUpP8bYZpBsjtuPv66E2mBOFLb+rChFQgQXxzVD9Rtp
w+O5qaGapLGm4fyANURDOgr3BME4vPWw3rQKbwbYGDg5n0SKDb/1RYjtLt09Jagy
Fe2N9Wp3r/0DTgOKkkk8xv+U+9JID5FRSfcKqVremfbqZ03pey4UGuQE4Gv843cS
aoQkmHoycLNb/Sm+0H9GfTHhJ8hcJOD5/Xpp1eT0PnmzbPlGCJunVKXbJQqCGvNj
+WHTuELhkCoKsoXO/oKb2eZUXOFuDbo3pAESYxn6r27auQg8h7+nXYQi3fZTj4ss
b+ijWXCX8wR5tlmqtKpKjx0mZQMQS/+5BwjbJvD8PmjVxpZ5RcyaCM89pFrGTiZO
kgwXK3ydRHrg8YarLqctNSBRXw+C6AmdFufCZL86etWE3T198cL1wlECpo3buWRC
L7eYkPV9mAJ7QoFHcrB5gXf8TQYw6WPDUF38uiCvY16Bv5hpzvw9xIxmLGMTUT5I
hNvBMxeviNYFCxtfiCz+IBv2tbA+ImMTuEI/eEWNPzIQHpaJ4zi93Cs+VJkPGxQc
fA/RPgK4OKJNWRVNnphfiV4Id3OVFXenuk6S5ml4v9FXWmi6Y//VONa4l+SZuRxa
dI+M14Pew4C5QqZPLxzs6cnTv2P1TcEY8noj2vYglDdskxq/aTkp3VAb4O65f4Yz
v5TDJMBNtvhENNfHbztghYncAstnjnzyckC9z4GRoza4D0/PF01jvS870HQXMEyO
7ggnVwcyxTRmMLvNjRd0/XLzA3v1yWyFIomwg+7gCjCF10qYz9ZE9zVeGiDuNt7I
YMPxEZQP43ea7mVZE17RPLcSo3w7kd3bxrN2pb5J1CLpV10+/HDKlUy+c2vzBguk
o7RhaqKgmT5M5Xp/UEyEsrAB4gJG8miNThQAaWM+vAnO3d57zqmq+CfY6RXuAMB9
cyH0XdNI2VemgiQWSw1KmIErS82zUd15UvRq5R8tnnoXoHEh+ZvbvJbXCwf6e8jw
X9J97LAYRD/DaCzeAoNpZkN2uIXy67GTbwhdf3ECPKJgJeJG9HFYdij8Midx5ZSb
zc6Y8ubTBIpvMReGPuzaLb82ey9pADbInynstTmv9TSEaAcXwrJq2Me0wfxurGQ0
TN1FbsWepD+4/s/thajCiYaZbd7xZ2Rco25YeMFmU5XabrYm9okKf+xyXeGdOYNV
Wkg4WRHLmuzUyT/W4ADlEqkrmJsDOabHBTZKNufd+MNkcKEBs+3Eitkr8U+G5buT
Pzqua8rNOWuzKlrmPIp603T6/AJs/Cx1q7WYDo8WeAEpUkCAqfQYXnkVUoBWwKL8
n1RQaBWeflKQI/YoMaFffCTJtuVKLap0MvilgivsJIGbfrsB+M/B6/Syq52df5Xb
pwE8Fz9cKGyT3Wgq2Zz5LpP5olRCA70Y5gyiRl6lVDUD6CoJ8+7nlUb5hfV4VTnT
UdrYr6gKXUi6isfeobxqfGhU44c9xicB8RnXUz8itICWD4p+/uAdVLV34mJK4bpy
z0etDM7FBR5gkBgpnw6LWPakJAdNsbbsS+7i7Rml4/lpWybgfB6bZU4DtLXFqDIA
0TjjGyY1JauofWpJXjTIUjpWkUs42V6z3nQtwALRrh6Y1T9iKJWjDmXUJpup4e8a
vV7aVggd2sRBS1mA+YIxC8yqW7FrCvbUIfQTtH+9q85MGCaw0+PMnnT+zIcZ8kse
dxcJ0FPdpvyfnfowMBFOnmjrtOzP0EYfbEUE7YOhTZYq6ErdvVDa8uruX060jnb4
zhwAcWBdvUHuXqiWNBErR7rCgtFrcmTj8zahuxTa+Hm7EDlLd2v5JNcoa2Tplu9p
8hBMuTq0K7PKMDoFuaqXzZYs1wIBaYUxvQmp8r7HCT58O24V3funclGicsEbDZ8n
V1A0CTaIobtUGZOoKHH2STmmsgjqfKUx2ttBqI4IGI1E/35wj7/0hAPb1j1Dil2I
yvYVDDb9xHHmjSBwIQL+DFmVaMAollja9TyrkAmMlpIhellDNMiCZCWwHBVZ5R4L
BywW5YJ+y6NSTHbu6GIYQ4pv77+0V46P05ERoeVI/1Hy+HV8MuwQNv0HM7VoACoa
s0ug+tit8eEmS5mUEOv5NtwJWHjePWVhQdLVbcgKnmDi8pIPcX/fizc6NTq940tz
kfA7qm8OHF9Y1VnLYMzQTck7htq7jGvHHCi3MFh8aWkD2lUqS8/4QzBocDl+yLl0
DlX71BOKgZhSAm6KcqYq7kthh4EkmUu/TFiC3e1NPDPTZfTkSTe6TmAj9n30xILs
YQmgx2CTxbEDSMnaTprupp5ZRQT4KBVQaVInGaA5O4JE26AGmv4mj1lnzx82HaNR
NuuL8MCDhatytzh9o9tfms3D/51dEdN9T5ddQIN9FUOKulFRuN9ggRvhU7+OdN6V
M1bqpE5ozh6c4CooLorNtIi8onzlDkTBCT9eShbDt8ufjj9awxyd/YAcPP4Q6LMn
AUKRLERESM5vJls5USf2TNzIrzAEU8elnymqDtT0j/xkd1BHcs3kekuglchAAF9f
8tKmq8KiOMet9rusjRB6xtc3p0MvRmG4gHDr48/w0eGei2VzvaifGUbAxNT6U1WQ
jumEZ+NzuoAeIZ9JOd6G8RaYhkemgvGTShTPFN35QqZ+/Jf31hlUY+5TVw71wRw/
c6Ifoq+MkGb9HikDqT4+rwUXfXOOdJaRugnh4waFAr/SG22mhsCl0BEC13gz+BC2
sxwHEeNHB83zGMnCpBv9toUnZzRIfhQvp8hh/SbIt2QJXGprQdzWy1MH24i1n03S
pN07cG1XuT97vHO27LNfMPEFyoxRChAFAqQra4PAZpQwXmzq4z7DdpzZY6Es3Cqv
l11prkTR8m6N78tda/57Vyg7JkKAtXSJdlROyI6CB7k+CmZQm7zPmqnyenFsghKy
XLIdHiZsGx2L9yy4/7Hoqvz4erso7QgJf+wGvZzw9WQS4fz0cgPOYs6xuIk9s+fX
/d1qHwsPTW+/fgaeLXd72JZ5jUD4D+TS7Dd43HD+JCQ76FdS5ZW/+uFeroRMN4yr
Zsj9zHiFkN+rNiEzFVGrM81mucoy7TkGWgr04WUEaUUX2QJ67Z8ZQdgneE21ewkN
w1UBXZn7WQ3vy1/Y1bc2/GwdQWgNJ0wIY0lpIQJzoFoYbizhit5+4ZrFAg2Cm8mN
OYkrNvbCLx+iB+kwHM0VnNl1nvnroV0HgTw/SzmbUpJ4aSSGpU1UerKJsfj8C8Kb
j3yR0F9BKr+x9/Q9F8jxEddrWN/6O5Be5IU4XSgABpjzfhKb1sSC3ABwI3WVxkf2
srIF64syJbLtPW54FQtGlAxDqNM7Ub6/vEwBGoxncl/cZKPSNlXNrTowhfJ3GBoU
oDxMpUeZ0uVVEDI5MHi0WND32Qe57Z3yjiFN0Uz1CvSoxQwG079jBWM8OPWHU9Wx
cAMK/ijjBJZeFmDKf088mPa7Jwp7Af3lFSyE3RF69n5yNwtP6eNOLYbQG0rfAgQR
rrm5E1fDYXNswCkSKFqP8f1StkF/tI3nYZvObpKutbO4xvtmgg4UM6ndEjT3abnA
0/BDI8o0L3aa9p+fuUWWE0LSl48egAuqxpV/X2DtDcis7GgJWqPDmbyq7BPtEhSu
33ZMVW9/SNq4M5yXJenTIZlaFJ4N8SBwrWf8fNqugimotwQ6/YzQkuepaYCmF27Z
1qVeSxjvHPvQZXmqgcuBTEpzTJpo6/26N1nN9QUa5Oreq/DdN76uso8+xuI2duqw
Py+TNjy93cRCdLyI6/aW6M3b6tB9rb74MXsvfaKNeRkR3UhBRWvw6rOQmCo1o89H
Tl2BPwHULOsJI6Y+dtxH9/eXeFEf4V2sbMON9d+TMnIo4vGxpbvVVhJXkFHnU0Kj
Ed8Es33/hf3ag4jdPobjl96+LIaNsuuHYcjq2X4IS/mehgj0roQ5wKZ8e7HJ6L4q
0U+S03tQvBYEJUc8n1eWvywj4fprjwrXT4eYqZsmcKib2y+N8NeZre9kPv53dwwW
pueF8Aijoc1l9NVOt6rt6mhHss8tBfzm1o8YwYoF2qUyrNLfFY6wQcBFnbTYchoP
tVpav5oTz2DbO4g/LmU9SqWbTVm18ca5O6qyHG5O3p/rkFOcnVbJMTjRXGXXoMIX
pdxRvQd9qQCmDReigbraIOyIUYT84hY6Ul8BtUgojkxgyS2GGwwIbMP/Yx0rAzf9
Tf3ZJKytSDVNHWKtYaTFa/VwkkTMQ+ivt+UaaNb+o3Ofv7Hpt5s6s84OCXAtNQq0
jeNCXOy9lttuMGZwF497ZkLut8l9tEU0Gr0CIQbe7ngk8WmH7DvT70CPOQL9eTmG
4GcnkjXvfJe9wY/w1JSKEgEBk7zcb625EGvx654onE8hgo8M6EhvRXasZ+9wZIqX
PE9l7021LqRUQ5xUglgJE1UHG2cG/8lGfKtV2MfafsMcwomtwbMM1It5121+cuIt
AHZngLUtmdPO6wn4SZWBfMHn01wHz6hFpH3Yj8fFeY82+h8n5WN1+sFsC98M6LD1
AsYuNpG+xYblNBEg9ts5TniBP56/GJwTNoZyU5xr0Ej7IEUOM3D7MmHqRrIeTPCt
HvmEhiywouudaogqj1Q42AUlUXROR2eE9lcSnb0afTmii8ZpneLA29toneFvLah5
ftOP7qPqW816tTNV6iuYxIqNDy86imJd/zwDeDPk9O69Xay2SDGcdnvqB3er2Zs1
gmLkeMcrK/I2tsh+fkiVvv4pWcMmM0YuFm3Vf6JT0t9pmN6An5XpPQSdldR6MzWE
W7cFaemllFBeS6g+PYRV2qxPIUlfE9sx2Rv3u0poZMGs/Mb3PSlb/B22XGuyLgwG
keAv2b1PoMJytYSHRlmejfNMAJvVV8xxWjl+I8rMz9sFhd0lY3ZEXLoAQlV6RyN8
3Y+9Gxc7m6P6U2S0JmzpmOui/yDWHgSj0Xauv6YbMeARTZjvUBts7EcRqiuF2m5R
jNbjD8wF7eroT/eh34jEhyHyJhOpSrr03pNRMQ2milIwAAmK0jqIZS19GlQprWX6
GXjBlYNg/xtsPF3p6Zsad6jemk8jFX+htzgsdUYrDfce3Hc2Ly7WyXCUZGDVoWM6
pfAMR2IQJV6ennbVKi7CUjGEBAY30vbUes2HfU0emvj0QHeep0pVZetWph71DpTy
aaAmS/ATQfFwU3u4GTjK0+PSTvuYXY3am4ciOrFyANlG2tMFcAQsJQGDUrbjpeSA
jdJr44HH9doPJjsYoY2UfXHvs7/96dIxwzjjywxwex0U6//ejcTe84IfolvqLfmM
Qa9HDotAbDa+xfHTBQV9WSIycsd+rk1OrbXdxBbufsKigmzyRsf3iHv7xDb1opbV
k4iWH5jSKYfjFUNloqNbgp358NESRvrjzf0bZRogSmQ9+K52ZXELoFc5Kp7DBmMN
q/JPAGgkdo09wzE8mAEc3x+XxIKQHZ/uYCOx8UUItl/QFtz7BaSp2q0pAyx14UOG
22z6yj7NHBoQ9JchaIBkbhU1MebkDAWP8+CQo3IEd5O8RIrUzMGuiCNYcTGkZBLO
n5pQBLEdbzdBD+8e0IC55730pNR18T9Gvluws6sFFP7kq8wL0f+IN3XiYcBwGMGi
DBOgYKAJNcVNlCR2nv31qk4NkQo+Et5RXc4HFnCTvEV0U68rbWg+Rd/8W7O4L99G
7dGiziedM1a/KSuvkCwgjAOdqpV0IIQTksF/ZWoJ07mlaD7ODc3/2mfYQj/7VKtf
Sv+hzJG262iYvMd/Q6cVoT9Xw+aGx1etvsst6c5i3cNrbxaPDPHG/5IJ/YT1Exg4
hgta/bsjGA2i4y0Mon3A3rlyYG91Tr2dGQgAEtzCajGhTonmiNkkGc/UUX9WSuBf
HBqRbW5HouWY1aYhJucvkYaQPhgYZKRe/5mHqJJwB/Lslv3spaQDYRyKiUGvCKWz
qR3+/F5IprVI0ySfcox/1YwGqkS7Z8o1dpu5cPy3ZJd0i02aKa+1axFuQ8hqmbPR
e5bxsYGkhWXogez8a2qSpzXbj3vL4UxlKBiqi8Ey58kkE57sv8g/yZH8M97fdcBN
DzGgtFVOzJhd/gjFxF1YaryV84zCE/fyIbHHHGN0uvhcWx1T/DiZVJF7+WxPYKXU
PVqCmt9sNZXlmFUbebgNjSneGvrGpYIfhPdWj5X07cyUSwJtezg94SXv22f5nTvU
pU6XaCmZ5UjbGlg1xnRjKczIYnp7CcknPbf9hGvfUeh8s0xIa11uYrqBIakkzXZy
nLb4VQI450mqpr8HKiYD1D0920MG/nGFyRFJhVkNBHBenvFXObtfgPcwQGUPrMy6
mV0rWk6ddYA65eTjlAlwNcU5FYve3PJC9F0VCQdU36EXhq8L9XVtOq7dHX//ONIq
km2wI0ikw7ynh+lF/dwqWsCgDdqfvUg8GroORbsDukPBBguxk9pGszrZ4+RdtPVv
2+gFF103DJpSr489G7OZMmv9QUOBU6Fejp2aVcF7/E6XZ6Y9IqHiOBARB6QnFMo1
5tALZMsM8Xiu8A8ttVHV9DbmLw/X2Hy5Qr4dI41b7FmLIqH+2EmP5o0OPKT7qoxO
K3TMRlhS62UruFR2YGjdlB9+HpCk2xDze29u4gs8ZnqtIkL3KDHhVoZ7OMe6ANCd
NdLXoAuAp+5hyCMLW4UHlf5REH24L/UnAGqRis9bLH8CB87nDGY9zfbNqlCxOaFv
I2odT3hsL+zalX693s91VM70B8zCEg44+OYPd6HUOP5PtEoCoQ4yxXoEJr9P8eeG
L0DGgl4MOdSq2q4sxaWkysKDEMYA+sbIAtOdKX9GywpcXUMQW7L0IN6Z5wAKby3G
uEn9VnAwFZrWInyyNiA6FnYLaXWOo5/WVj5vALMXVXP3XoL6/fUQlR7AmUHFaDG/
iJOaMKoGRuhQD+SaFLvw2MjP9+Yh3bfk8SRoW85aJIq4nYs5edm+b7y+/J//BBdj
tag3luAMDFo5FVlGZhRW4VYFbzP6VfaHMouEn5402iLOsB0iDNqUCqmH03UKbzw1
TyN5BhdeB2YjRw9gnijmA2PymwKXrevun3DMBhuBEKpEY/NnyYiNGu+UYCvYY7PB
AhSq+Qar+CZCJDhw2CPrwv/drb0TBc/RzVonKN75pscORch0pxEtuvPHxk/hM32F
RZiqfcpNbYxmCEFC/Y2iewYHvINsP8oYkl5HT5eZXOvb4SsVN/rLDlV7y054gjkm
LEg4pSTUP+YISoLb69PUfJ8z2hfLiXnfZRl/PRvdp1UCF7U1GjeWjgQNc/GVnJcN
GcYUn2k9PSAugnRClNFwIg65ZfjLp7kxKb2pRHjiFMVG5T+s+6BoM8VUx39QuqLq
HU1bs4+2EoGLOzoOUnYkNkMOHailUUdBxRyS8HIKGuX6flSlek/Gqg9Fx8dbgDfs
Q78Qmjscbzb19Kl3FujYO5SC0s0Z7+XTVflPy3FUZXE4MRPKEwOK1tMqhUaNnZTL
SvfZVt6LTMMVJyFcNWdSWZUlsLcrWMf1vNlPdyjEtZeOLm18n2rUtTOTZOzJJrqe
+BGwl8qptDtbEb1TuKodbLA0Nqgy6grz0dhmCkIwrCvEkw51achXLSWVS3D/X+DW
Km48j+Kb+RfdOElas98kJAX9GrRcDCGi0rQedqr0QJ36Dq18HxU3LdbNn3v2Svtp
NbhfFfkgKxm5aRu67+VItkBt0F/JxqgCWKdYIMgxVfgb4omXwxZkBXEAQ1lSY4vf
0oFCxiL2wJN7SUsH5OekxTSPwGQZKG0tTCULZR0odZENW1QG+iRH493Cv90/5eQR
O7dPOKkJ6bRZwy5b/qNc0wYhq1socgzXySo0E+AUdMJQFEWGiiaV2VZucWctxyLx
iNzOEIiMOLElROTF59Y7IEcE4ndgsdbwfbnxvEXY3OprIBT9BQdbKFnEqBi6y0Ox
fjpMP1h4oE5/9Ytc1MxL6Xb1Ls/uB53IgdJ+byEqL0yb5kgho95dSFxlFJgKFizu
V6nL9//s1Rae46SpJr6OVFdavsxngagWorZ1id4YPfE97+O03j2NOy0r3Oyu4Rwq
ahlm1/iE1Cof/6qQS4KLd+jtFKz2afiXauvvwB/nsGrUaAgVY4uEvZDn5Q52qqPH
eqImEkibtZuaB0WzQCceQpzbnfI5BhHiDZ/Y+/LIitUBTP2nMoZgFYb4FJ3B0m3K
RIMAgAEEJlljFx1POs/udU2AY0CNsSN2ylWTdqjg1xN/eACMQ88WWjE9kDtmMGiW
jjKDNR2FEXJJQnKxgiVNpCPRJ2cmuOQ1MrJb6S/2P+4Zvb2qYwv4gB95Ntf8pJmr
Zqhw7+UnFW9v3uMInh+v2HALFCiB+Nhp7pDq0vN5LGiJKdsFtAGmFXmkxB6adOpQ
6nCgZAIdKPL6Ru4J0+6ws7d7PWiusHSvpmSksliI09eeKBm0Clj+krduqSr8eTkw
YGCrEF4sMSaRx7cdayswnZS4oIIhcCPwOopbhVkRYHMcQ2OHIfSbaI7PFSKlLXsc
5mT6c3s0wlwdUlrIEaFrUHBxKPAatPWCDIPCMglG+dVMHib+NUJCsAkBzbyKTfnD
hlLbe0RQsJjehTWOfCEsJ+thnG9SR2NdxePJgunXugEP0cRi8B0+E1PFOMJf0Wjd
qjHqnMZ9z0PXskONT756AgBpTX3zjFMKe2wTkDniwxd9/6QtuNdyuCKS1nbQGwbk
cVVAUSn5MiAjnAqWzgPuLhvPBq9ylNYnfrL96hj2V54tNoS4QdEsBXWHNcP6JAmi
x9GfBzr1oFSK736YGsJhW8eIUc+Q6RKYSQLgvEa7d5nr7IHSutsGKsgv6yHnDp6t
QMj9cFSbgAOBxLL1PvtibeMnZ+M7bah3ypPfs3YvnBtmhAfVHy4grIwB51t60J0N
dWQkKd6iGsPsGFPurgGqWJ3AW29h9Wa47dQkfsuLn2/usX2Z1ONj8r53rB9JCq8i
6+MGzlLkAPSlW2EOT1nyk7QElF6e2gooyhOyHKAIxkJSh7DEjHo5dP+/3v/r/vBr
quq+cbjH0yDE1s4/u362vZK0SxVHG3pbvvIqiBo5kPFHmvIfYHOTQy0aTpRHBsKM
ifixNyZIa/GQvt3h/7acWR666+ufO4dXCUrdbbhidZAnOZ0NaM5/4Tu/lrcv23/V
/94IFW1lC2epw5OCok6BA8onqaV79LS86hj8z6vrwNx74t2UTaepUyrAZ9LO2Wl+
644JenG2KHjXDiIqtN8sQLfkBqkv3VKTXv9mThZermD5vbyJuiGxnbS34xfl6OP1
7eDkPk7JGKnvLy1sRgXYNp/AX6eH3shAU4qAXOImFJHCgfAtyPnIpoyiROpPwQe0
565bny8Aygg4MTZF/95+hqUqJQDF+Nz0PVP+wM/goUWNTtEI21nL1Y3Fbb7gf64G
6jD0HrmTwgXRy7jeEnbsefIwdn/Nq0UOH0c+x3bOZLG/lz0WpIM/dp8smNa+a2xj
Cl3QXxWkw2eFQfjkvWkX3qyvQuI+q15M23jamHQrVS9tXzRS1pyBpXcSOWsajDad
JT5W/KBGFE17DDh1X8TwFOLtzKLI4LbTVgGlxkDb2JHTmX5+Z1FsE4/qdANoY2ri
h5WMqbm/LABXpWmwOlURpK5O+9felrNt5jdcGPU7Iidzi9f7sBTzornSyWUN/XT3
rAgoQueyYZmNHMgfzonrFyyDFq19khCn25wRL+gxAKfqejqItcyPMixqgJyqYwKl
z7SsZ4WxDhcINaC/mAeOyCRGQAckZFPhEJyi/l2A9TMpNgJHAFKSOw0qGGh8+En5
yPS2AYlY/+GYwIfX0OefLCZom1qVqwz2xExyBISwY0gC/BqYHsJGPhiPeqyUijbF
C5+I8vUKtLJeBCVknaZw5n6Jlt9ykmOjBwU4PLiKT/I1xxC2nxSp49LDBsizFouD
0+TW47pnCepTVrYwEkj3vXgCR8hjcdwDMPubb9H+xeCVfr2InWSTxYJ80teRWjcv
k8zlNfRbncGMhiDiBHtEGtV3VAtFQhRlM8V7gsOAdTmebUgZk6omulkkuQapXgsu
/uewJqcveMb0MNjMClW/5U0M9EwLjh7uOWybIEhsd2h4pImrhociDXAJNWHbHwAR
2eHdAKYOeEdTL/o27WtRoyvDklbprAGUjGuSq0ictwxqP+2lfdz37yYEjx1WQL3G
kdxb+2l/F0O+U4TClunGoAozSHNOFhlNx6F+EqFWhDgk6yde0fp5fz5UwULGaIhh
EGPV4PmqU3tq3XlW06Z06zTwCmUBqjniVhzyyjj1inA6ndBCef8POpH9Y6jcXmoT
Qgy+hV/Dy+jp7cAbSZioWt7L84v3QwCV0WWl2pHAmKxz8wG8cjW4RoeM9yikyFUp
4B9fW3WF4g9EP3Ms8/LfDxfERYSgwd+Azmhr9ddjNfPzvvR7qR8wnpkasOMjzY5c
FW6CnMrKgKJF3h9H1DZDw9h8geVf9W2sUqBF+8oJYGHjzINXrgNCAAjD9Ic/rCGB
5O2VYIx5A2VZPl1go6iLDaAyOeE9R1VpM5hcVwHwH1VWjhibUDHumdZv0nEprP93
7LJ+ol+U2Byq+St/R7QR7/eV5yTFo2dmSJLbeByJ5OLm/ZYaDWyE3nd7nO+kWYuT
zbmBKwOJPY08Gu0niNfF2W5h57cqJ5JqFLEpXEe83484BJP75znUf5dQxNJkYl24
YgSxgO6pgl/aFfA2u0tKowfXkXxO42pv+tYwvqft7v0glYMgUBIf6ZX+RV8xOXRk
3HxfTTFK161VyGSWgKMJ4C+xG/qF8mVC6L+wgrPFxdQN0lLs4cOCPZeUKut1t4r0
rn1WnMIOCqpwC/3ihTKOc4zF23krzE58BDltrltrSh7fdNWpHYxDhPWwpbfdD/k0
pGkbHV7q5PdZ7T29sWm58o0CZbyVZDIB6QP3X+ohjtjrXQFtQgzsCkA/Q8B4Lg7B
86E/qs9CafMS9DEvBd9LMWGazjYE8XaMCLfE8DqEEMJWf6jDG8Xu+6z82E3NzMli
1r15JaTllfMO2ChpXqeDdZLRn6QWdkbZZE+PDxbgJcsJpBOIxvq+e7pQPxcdaAZQ
eMazEX3zBIIVLu2JQ+RjXwI3ae6MDa8yyw/i+1vGOVoihCTJEnf70+xDZWp0EGa5
ZQ+JkPndT0+mpalCf2jR36VmigMihpWis13aMT+lL0a4lIf8nzASXfLsqcKj05es
9Y0qzZ9ApJo+/MMv3szy8SOnRRo2jHip/dloCMoPsatcHWFGbEyU49zBj60YPbdL
hFlJXMxFMMmdmoviefpz3vBDTUa1i1pRc+8R7htOgfWRHsWbYmizv6xn9a2wPKSc
nF3xyHGmvTXqOVxCNlOc9n/VMQ2JDIgFKGtUiJSKeQ1oCQ3+F3vB06Hq6Iou39UN
N2RGflZ0YIT3nyRjHxDdkRO+IVP+WbnxmRsrh0aWZTfP3lSFQKY73KWLYkYtrQz4
e3S40i/kxNajEWHvAAmAxpNovGpmllvCFMcU6dod5N4G1dcKpQ6ajsbEbqJnp2aW
41xZYWkC7k/r511PZLaVymwO726yzNmHM7F3Zg9yErcovUfKIGHM0Ne8u/0eJPtf
uj7ETxt3F6mBBo2g8UYlULNqjBd9aG0qCIcSlDbM46I7uCTXvKnDgv+k6m+HRWYo
JL8Y4K+ouO4XuALSbOuRiVKY67v+lZMIIuzLnWkh+nHc3Fm7F9mnUGQ2/mUwoSkY
EaKE0lpnY8QYsSGFK6+fHF3jKGFhKzsAOoA0OCEXASJk1CfvZsqXbp96l72KXNeP
blkn8vU8blcL+2L8C7XfMak1rp58ug3WlUHrkgmhJGOLDhBYmRqw2E7M+H47vGZh
IhYBI/0sLrEEXeQas6oV+ONwZZxJwYRnqMBIeNQmJ6yldF4yLWt4Lw/ZELEEOGUm
+WLKb4Yga8E1puYUDGChm/J7+uQRTmNoJxQn4+H2a+XRhAuD4Xv4jjjSVYwjtk88
p88HeTEkOEzF05atM1mNTamBiKOtBAdRJKic7RlqwPE+pLXlBBa2Qo+udNWpwDVY
w4CVyuyoaLzqnlqIXXpK+RGYZJ2OF69KI6Zjb6y64KMJH8ZgEwtOVbdqcR9qIKM4
bl02YYah/TjLm6MXIdWQVsI+/fAydEpUuvyFLMXCo/gdI40nCpQAlaiZ0qHOWVxE
JCKdlNoexKjMv9/oKMbH0i0mksF8/Qqk4s22r1mdOCd8uHOwCl3SoU/RBbbmEx4V
QvlqlcML8N2soR6fyqvoYwyog8r7jiQ8y5dBatyV1bDE1ERoXhwbHX3dmpXro6Jy
+6aMUsOwrEdlNiZcqNvKblpENm7aNDmn0GaMFaqIaAlPqoKd8+qumBom8SOPi1q6
HH126uU/XFlWl/1G3Q/ZhzbCAiYIYEJVWmJQfZp1NrVZYNIefkRJ87W0VneafKnA
aMMCf9rbqMBXdhz/dDv/MiEg8y1mLpLZ3Lutp1kC4466zFtJKgGwAWIh628OrHzY
sfWgGsKN8oQ3etnsvkGqIDRbn6t1Y779VjNpEm9iRW7nY7nLNIBTlh9wrVVxxrJj
hQ7Vc/uWXqjisJQiFsWZiax6Y9+BzPYnD34ss/gx1nqMzdmk4SxLzKOozCkfXoMh
NDOvbUTjGIq6m+ZUPe6p4EW6mkFfmxOZiIIzeEGZ01hhamxuwnpExmOTv1Wby9F9
G8uFQdbD+44Ivy2aWmEHyiNi4yQi2zHcCVhuPzwB4HDr4XZhyD0kQrBbTL0hZwvb
S+8yaQHH5nzIkcSNF2gc99P477f1h0LTy12CA4C1dqfWSkioh+65tIIV+ultkpnJ
nN+jqY5Nb3xmn47+uSkxPi0+ewo5mvRYtRd9+ubKzjQU2G60luG+I5RnWDx93w+x
0k0TmVSnFyAN5bbmYnNv9l31JmBhYmliKB00q6o9PO8OInrZ3zEQd44JtahOGl2T
KGlRWey6I7uZQLt4Z6PEVQRHQ37P1BfbeG4Igr9cYcGvvC4KEdiac8C0gj36V86z
95qLhyHsBK+eufEAIb69qZCeSHLaF9C95jL6et2cRYomtxN7W2B0s/JJKd4J5uEc
3I9WsFP66EP3yh66OvG2kxcV7j57v5TRU8h+JcqwY9VE9zEeqXsyHkFm4j4a8QWv
6DxQL5COrNqEsPgCU9coj5BnTdxEo1jv/MYf5bU6dB4oVS/fLV6axZbcbTJX3INn
SoFQjk7IjAySSejOyyxA6U7NjDEvSg9KqEPCjzmuu78DDOedZFELrlCz48bDtrTx
xacRoKz6P5nXn8hY2M/tZGzDsHutbA3VqmCSFMjw9SaYQLa0l3Q1aie9XHvaxuRq
XffLIKIIaPi4rVsgKXLNbUyRUGt1fDwAeH+uxsmSfFoIbRDLR/Di1opyl7W+z/Uv
hNxxyc1ln7hKgw6EmqX1WG2EZHkNjZdmJDyEXSi1jCxp9nyupfgG1a/ZgHzQHyHi
Cqoa/4IAKY13ebdjnWkr++1oc3r21p1grNyukCUb4BTnipAZ+R1FydpC17R/N66O
B/MGEPbgk48bVYjS1zk7KuznMc/YtZ8t8KZFpVI8wb69/YaeqQLdAVm345TMIK5j
epNay0hw/6Y2sBfQFzLz+pLzxau5XBEv5I6JRrZvEJ9bdiu6ZX/ADl5+/v9DW5u7
wsk583DfE4j4i1wSF21eB8hm6JYw5nmpgj+Hsc/qoEZXz7wP6bEwoyO8uPoklvzk
plVmHJWbPRvFnxeNMsPgc8DDASuRVMt8wT4hG9ce8iGAas2L+qWTGXBI4+QKnINp
Xn7wHHCvhqIThyZP9YWeK/+dlozdDZUB0NPGrFbcXRO++bnCL+f7HOriP88XBhJo
aCJdLT7YO5i0tsUxvYPiUwZhOq1L1qldVxp3cdqUApIscd+wLF51R+2Q+CK7MiH6
Btz5I7BD99VeXeLUDre1VjclI0OCkqp9Rr2+J/pAgOIHSOjGbxtiWbR5E2WFxLMC
HJE3yDA2jYBGMWwYaexyA7m+btfpkZRwxiEx3UE6sZJaiNQF5sWKpc3OtnigX7du
A30YvwHluBUyJfwi4xUgeRrUC7/YTE9k0V5U9YAxgO7bw+tcXRW+yhwjGD9HpUqD
w2I6qVdJgUmQDaQzzJNweQinEA8Nam9kj75TVoYhm6KwvhGFQqpjH97l0r0836WD
d6DmKeROEgMg3tU6zmbLlmoCTHpXGr9N0mZtFcchOpjaS0tXldFw6xSJAeWST1CY
koM+WYqV04xEL84IkIzF6olKbM+Msv/qU/Bs6/SeONNp4ma7YIj1ytyUJ/F8xFRh
QBiZX947nNDTLfhnYQI9bcD+Ut3Kz+mdWkso8Q+Nb18a0iQeeP1Sa5pc/f4az3Od
UyPgaf8GpRAeqe6F19KL+Ub241+ZQAtKRrkyM8HaQkKm3M0/+lSKzSgDR/hHmFul
BXP+SddLMbQRVg+L1gZP+UsrH5cpXIaec3goa/+5bJMfifa8e+7kN/mm6dJNI7wn
n1sOKnAm9M5W0H813QpGJQW3nTiWs3+hupwrKfQaK9IGes+NeZ0NpfWhTYNDknQl
imjf53eylcGNlXLjgsF4bvHXnXVGjCOsRTyxTur+c/ciVkdANs93f45MdSGWq3jk
AFIRzevHOojpQuNukQpDodlzhEI33yWqm5TJfybDvkNWtteSBCVAFiBGgVWpi+bu
9AxkSNiSOckAo0aoifZhQEliSRSzvbV1QjS7XMBPyXMskxjabzTOm+N5RM0nQu4L
L1ouaKteHowqmFNB67Sd58EMGRK/v9qqRvvoe862KBKijqyTta66WYAFe21vo9fF
YDoBrSYuL5ctF6eJBIaKuUt98hqX4Ik+VdOa8c573DzPJ0evq4YPYk9x0znJgPYg
TmItYYN8J2Z6rQyI68eQMK7LAY1BLV1eLHlBwNj2GXCj0JVQ6zV8wBL75u3VbCIb
WmWU6rbr4lLohzz3pOaB3cQTkHTBG7r4aYBLfO7XiHpPTQ9kmfiWakvTlZtiKOG8
80lQS921gYWRckP4srrt7W19D2wtLcoaGWIku0lUMWp2aA3nM/yTRhGY2KhuXFm1
zqV+LK80djY9RQJbAJCVhMvV/PdLRLnsE8PWRW61sMx8hlzQ6Dx8/DpfE0qZy09c
vDAN7HRN5nAMMxDMvfcPZPyG37Ds+J8BGKM9dYOiVjeKaalH60r25nl9yCVtoW7t
1GIPg+WihH7Z9pZHdcoczzNwy9P4U3+TOlTMEzEhUOm4Rb77QuQkQavWNoUBKo1O
mdfDLocRyuZVr8LUO8P5+ImgVdP2WTYuAtiRoqgaH7wDyWofR5Gq+rYxJxHzFQA4
OtVSl4o0XJzM4e8mo7zWhnfo52Zqvyl37vrKDWa2kXbiQsOQV66+JLXnREcYDITP
PrhrRhrWT1+7mzWxO0L3Szw2bs352UT8/BwFU6jBoCdbCT8RSNkokXEEH9RqIGlt
Jd/mEcWYs3f2C32jUT1o7HRhNwelYNBIDxv1doU6FbhTnN17LleCclRYkrgTbpo+
glaeQNEqTSvtvVPrdpMZMM6HqZeoY/FbzSqVI1ptNoMd0OkESnYUt6D2q+8WDNrI
q754hbblFBgcEzpFweiTr269OqqTKKo0gZt5pTF2MpqWn4b3BM65zktKHKFIdbkt
s4s1y3nB1QpEloHhcAVbSUgRY13IRG/wLmmwTFEWUJUMtKqk37Xk1XlcwFvEEutI
BiR9PTvCBOThBlXF44sCizzTktNxV98vqVUqgzUnQdP9+yLaf3m+qMSOHDUtOQqK
KPYVvGBn3KuaPskOTvidUlUnLTyQeTTF8IVraWmy+nE/19E/KoWytlrNQTaD8siL
lZHogvDSJU/K0bvLez/qApfyGOOL8vOB4ZGGk2k5D3g7cNUE73lVvJKf7HmOlUZp
yR6pPW7gYsOse7PHb4lReStzxx502fIPnpqLXBxQjL3+0o0mMmMQroeNJLvEzztR
xTvW1wielHCHoIEzE8lSN3zNB8VkU1srvsVxWidqgyMcMJ2VG7zvO+uA5borLrud
nhXEVCfzYaCW89i77B55nTm1/iHiNcljAi0CSxbIYtOdmWHYgeZfs10dX/NWmJUa
0LnTPmr156rtsnGmkT1Vu74V8GSnfTeuQXMC+nxLCnEnf7EqzUjOHif0RKX2RS1I
FjoYFkDKZSZlRykf5rHin64pbnhCEwgbc11VHAuh9f/N60xv+vZPofoOSxrd8wwX
FOUsv6dHJoGsqtD9JRgHYGUMmghIC8iwtuBE10h36V2RmmPHRtRb0Jem78czCDQA
LJ87LHtTsCFT9oHI9CZNYOQbktvg6+mquAqR1jZQPg1m0TkhqqsAeTwccmOPIzYa
vbwXEuB6M2+IJOfS3U1KuU+w7Y4FT5fIYnhQEMRHU2hHEPdLjUBuew+dl/pQKqlJ
Lg3hrhe+5/wNvC1yDzAymQwmdr4AT8lTCzjEi1Y66ujE9s9vcq6Qw/C9rIHl/Vc3
SI2g4v+jahOvXuahhjxrjIsXw6DS8TvsSP2CvW5wzXavEZsqR6zMfrZZ9IVwxXIT
eZsIQ1cpHcTCDceOHJeh3AYskhTtQvbaFVPJ3zJtuyJj7sA+jjMs9lng2cwIFy/J
GssYihgN7shK3My2rosNh2dCvLYkfnFUyW9LdW22mnX+8Ioqc/DYk8aGYAhEymFe
if8r+PsjPy1ugLVR7v4wIOClXt/tgFUS//d6xnQLqP/HWoh3WX1SjKGPFu3vDvrH
Y8r2txaJNuIzimxUZysKikrdltnNBaE8abigbxf8iZpqDlW+UIGazDmS5FmVXW0S
AkWYSXWmHICh8JRAS0IWRBsoqvddQcH+TK0OpMZmUS/IfZ6yN3Hp6IXoO3OFzXBF
h5BcQOgRC5fWJPiVJuONrPkFPl0XlOTmjiwEKBluwXYxRo2W/TLu9DoCpVNqURb+
lJ5dURwXkTfFYgFexbmsdTIMkhusj9cdqYoq42V5ZjSnJkkb+MTstdUM6rhftNuE
cKPGiTMIQBVV+sKLjmjjd2Nd8LjQaCz2kW5uAWSF2GKZj38jSIcCUioLl2LnloOt
8IJ3AYkzlC8iM/97kjRMx8vi6z3yf5pdZTBwZrLnM9YkTPsJ0KD8Vsu1/A+kb+Oa
tCU38rPhNCLrmJ0vedDvR9vIl9ACooOKp+OThkAQaKekuuNbBFf9v3g6hUejwxS+
52cZ1VSZLkWUXYuyDsNV+/YXFxt+N+OxbvKAllHD8k28ZQR+7EjcjmCimTwO8Hu1
qeXmj+v7U8fueRMiLlXqj32qOo2DhaX0m3tzMW6NVbGu7oumeRk27BVHtsAqtWVK
0wauEmkTJCVW2OFu3QXGxXuyBPlheKeVsMyCAzRDqunKtEprM/zzJG1QxjDbVaYT
TwwLFokK2EJRymWw9/bgG6OElljZOOswLMycVVlo/P+YjwnEczqpro/HFlcEDDZ8
lFw6xONPwsUN52OIFWkraBHHYLNYpnlxIkue1VEJvzCZMYQsu/R3yibcl3yGet64
b3sLUK+3vB03hG/YpweRi5VnOZe7UMG8knWYhj1zzzlKK9Ddst+tcXxuERIEXR6g
abxy6dSDHCZYRWRojilMzaCCuqZ1pUPDUBif29TJ/XyMiZeFl0JkRBF+AhmEtFol
9a+8YFOeAYDMj3U5mFqXnrcj7TeDjDN1BmrCf32K/ITe4lCeJoOFOEAZ2QqP3MBi
uXOxRp1Q1uJeaKX4Dg94EkZGja38LUiR9Kbk1kC4jsnla61390rVqD+gz6IFfVoN
ub2PQOk0QGn4xL4dT7aUEfANRUIk55H1NryBrEhBGo05vR2GghxDSCOJhALsd7XU
RHsed4fKwF8GhbS+B6pc7cZvFlwMQQTcWa8XL8YEzRYz3sFnnnVqlIAbgEUHA9w0
BmcLzruxkQA48DKwKk0LBis8uX/jtuKHUa1IDlL/JdtphuCKqUk73MP4d1i+g3yo
/YRi66Wihg/UbNiC8+TNaqjU7D4atoWlXlQk88d4rZTaeS8+kS2w5n0lcBEHLHmk
VJi8QklKhESKjQigeSZTjSIGhc9+oNzhMDKcuba8RIQDC18jo/TQLcK4nA15HRvC
rPl+RtJrl6svmlsvpsvpQexxzZabVtRUEgCoFt5dWGM7aS/j27Kdm8qBJzkZ69yI
tZp0+D2RF1jl+ytNM3S/4K14YXNWFcPF+xlk67aunxocrZ49Rv8XsN0H2eHMnF0W
BPwUK+WyiaoROTmegWoGTkKFCDnHE2WUZpk64xR+Ws/sfnBbgBkyOzbM9HwU3eY5
F+onqXXxuGwtNW4fzlBVShf3qs0cEePnqD+2ZLzAT9oiAku2itzKr2ks8wkxNVl1
J/xBao30whY/mvxL9n4NFbg6DBly4JzbMC0GWgkKtNFDRhho+YIzgP/QVU425+Mr
dqhd5zrgRCp6d8NFRKxkUojDgwpFU5rQ7EfPwdDlinZHmVsqKPihhB+6SSHEfkml
sVTffLYBndcQQkfqTeinRIIJcOpVgXDWzcpah5K2TT6p0TkgUtfjH7U2su2UZtsw
qYCf+OU8W9EGOHWvYPJqDAseVdzItJqpC7kvMbJqBFPUuhr1Hn/ZiGRBOKQmA3Ew
PQvwDNOYN1qjoHJkAtYZ2ed/x/NSjjIA49r59n5IdrMtjPKgabxCxE05WlrHsBte
8eIkILS38maXwB0gITDim1jD/Aa3lRibo4buwpjdzxyJvP2iTxoFy0F+EZZUMDvl
xlB9BAPnAb3KVxdmwTSefXTIE08MtgpDbB/9QHxhUxeXIcLdYukJk3ROJuj3Zgpi
MilpwI/CJmdl+aWguG17U3/mne/MjGed6shEyvxSYFm0n5aEFmNiK2ByD42hj02q
jEvv9z+C4URVKPKx5xz3Zfu/c+IHN1QSSMr/W4bpt8Nt9cwfPbHESx65x2nHvKCm
kG854Qz6yhiJkCsmHFBWpx7puLFQPHArVaySzTqb4HmIgS28T8kXkSuAi+OTnl9o
nfpAFdPfmclHSFILJkBA6CBEGQhU7YzJ78x24Yv57YSNTp/PeJiL7kWMaB7nOwUF
1rrPhiw0+cMc/TjyMz6WCHta9MIDydZh21L+5xGIiSyBAq2oK9wJdFhohqyFajzT
Dr7eUjVL8yXnbL7+jN+RArjtj3KrB42Nki4VhIAeW+OeRxgEKjX9OxyWNpSjZ11c
I1VZV8YMmczaF4lAS1bzZlwYxEHf/ejW4vkLHAo7U5OJOML8P5K2LsxiTbjXrwsn
4GzRiin+OZliuio/v55I+jdE0OvzsDVQNn9P2gvRVmia8PsVUkwImWeY086GbKg8
phd2KX3uVOLezTmISIuNwTm4Proc9MYSK9TiNWlZgs+FzG5daEhpfqeBkdwxEf/s
YwBV771jBxE6ua7pTy91SYZFi/9nUn1Hvlv3G9F+pXmIUsQVM1wTPI7iEajT3NMp
pn/LPEYyfbRhfQdCEBcW0XIj8tFCFTtNR9WfGqAAKVvmQni4htFOZg3qZkfLcliG
gvCdH4dqPF4657DKgESdIsq1m4sELmyfe6b5psV4jdXm7W6J2T2PfpCSt3Qehwac
HbcvUCRLzg2oxY4ZEQxwstGuMbJe9LnWbcFq4r1FYg6ddmJZHHnQPr1M5mMO/BX5
7VmwmZ0HMYYhdExxw5I8Ox20vNpSrc6PQVOO5la23g5cprptSJStOyeKPwyni46H
mt1CYz2yEvQhTTqQrzDWAxhaUkBJTZ84DHHMlLm29D6uKzv1BMIG6nXs2TA8kg6h
Z0T5zOKXZCrMj0HNBLHC4W5ybNp6pEfd+QKsTrC4N5CKOfWNm9yPukBEQAJfUvLq
z63CqY+zs70JDc2aL8CKmPNpY7qDIBA6bKoCZXcSe50fG9sBfe/usKxoaMNUlO/E
O9FDgH8oXY+cGsNYr7nVqeyf/tnKinjWDoyn1Mj66wlL9AzpvSjwAIkgnaC5Tdb+
dfw1LJ1kMHgZWiIenqQfO7ESsOkt18PPoXYSO+3dFmmEXWd3yWXt2ITFQJrlE9pv
P4jyU7v4O+kl6aS05IUbwNdZH4wf0ElWrgaVPPDzbl58gbp81SoJ4aaMTvlJ0W97
VPUOv+DaPg+f0QaXEbjmkS8t6Ql+Q+i+GVrbXynzuq2ug088tnyymo/DCQyq5xNk
YFuw/YN95yagWHmrY4vtmN16ituJduoIR7rHVzIfh1D6j/Ofm1GqaULIimPsUDYN
20AkaNiZrctd4alGDLrBJq8h1FMjW9qaRNjp5N+7gy2zB2qfwHh0lYKZXuRRf8dT
sJeW5D+Doy2cKgKamKt4NesZQyx2Bb7yBUrVYG8ut8R1F/8+1qR0Kf3rnkOGX9Kv
Px9mS7BUKQhBN+af4Lqb4K5QgyjuSebs4DyVfir5ReYHdIWnMz/nLSe5pjXcGxs1
R6dz3/dwV8gEcblczutse6T3YVkMhIyB9tIlbZ11ifqOF5ZI4lmtDytv5nsduhJB
UNSJzqpqiqlsSU2pHP+aSA6CDzu+WQQDp3iNDmaEcTM9lPHUCYkpynTv502auRUJ
Z091v8MraRMIhtxYJTqHAQJS/7agAAFzKbaKZOeNpoe+Zr632scmPkgmrRW23nHI
JflWKqeynSdQkgJuXu4r3XHzQXnC2InsMgXrmmMyEEKQj3VieDpTyqLXo24HSV6s
zyIOHfZF54LwAxKeX9Z8RfJHuEUywj8JQlF6yhvEqNU/gwdguzXqolbkq2WYJ1ax
xocU2wOs1bDK+64YaZplJ+Dom1/csH1rB8lNdFezyalreP0eBxLFJkK4NDMBlK0f
HLkoEBfP4gIlJYpvul8lj+PkVim4Ns3cdp8hEjOd7xYXu2einB9jp6ggGZTCmSK4
aR9rfr0ocHx+gAGYKrvC5lRfOszFrIBTHu/nUS4OTrwgoIvBX7DyzqZmbm1BlGdr
TF/tsuNLwCOnMVuLbpwwr4T726K58mb1Rjmtf1baFYHoWxRojOvDxsH7aDiKshib
AVTsBchdEnJHFSaA048/Y1xWLD41z9bccrWYsZfQpyJhbc7Vse77+YP489NRILdw
/oqXLA9qH4xC8+OxOMPIkXMlsz9UCZxn3duaMbEMS5tmMUnNgNSDBxD4ArH6HvCS
4VYt/DmScKafAsZmbBuAodHWZPFYyyQLxBcokQb/sT3iDvAGTA2ldpoCsTTI6CuA
hu7FJLQy1FtExuaBZ3Z9aCgI7RjfELFqFgtNmfYaRIfoODMxAWvntqM4qdIMA92u
fOIrjJY2s3SFPBkSqUni5hBWOb4JBH+0eSy5ByEhwdGy7hJa+uk+PTzo2X8IkFDS
PDFY22E8VAEbrVpBEmhiyp0qyDEp73FYJsngog7sAhREtZ/a3ZCmS69qqJdTOGL3
R08Y6tKMXmw0ZmktB7TL6rqEKRy+gpG/QDh43qAWae79cNAPIm0c9Lfi7IXcoMnQ
QYXhj+4Iu89vv4Y0UIaUg5pcxT/nH4qxIeDoSXMt3YyC62qoPjQpD75P1hQpcOJZ
uP8HLDedlO0fTXjICsm5kSQX5lNTgFI6byKVWvVBfF+pGJhqiWgGmyM1g5iEK4OX
wrvfq/H40F2V13UiOyceLJFnsdkrYAsEFG6R4656h0aQQ7YfxRHrr8aJXXzIYOQ6
DO7O9Xf6i1n2a4eMltsFBK8zQdYN/LuQ7XWwRaQPf8troqYImsoIDRNFLcNQEpy3
QaY96LwWoIWmKDGsMHvZFGXB1B4QFrGjhLOM2JCKOVtdsALUFE/P6mydDX85cZtL
cvV00Yj6200ch9aM524iuumo6C7teNH+pOn0n00MYzlawUWtuL3pUqvr+oy8MOjJ
V8BnxS/2THSvxAGZ3M6xYCAuwvutZpew8Wa4yzbh3vijySopVXfau/uWmsY797fL
4Y/KOFyXFpvKpTqueQiON/QQpy1BtMM0pwMNKN7oK/K4KbbFfb0dKYvGlOg7XSkb
fTN7/B3s0NY5t4eqSbgX74SfQUQirP7+rWi9/j5NfymcI8jG2Fe0/tKP4VB0mBVC
jJv/wG55tv77p+AeEdTQ1Cj6JIWrif8dQ8v7ks0KSAx9y6gynwBefwf+iwLB3s/7
zkY3pTYb0rVjGq3LtLhUBjy9N6MrITSLovoZxEJyndP/hKQq6XlEETjVQyuTVgVf
xom1uhEaDk3KmB9UzyXLtlXGpZm025khVwa5Jp/MM+zKyg1QTC3dV/B9NPUfTXS1
zW6Qs/S4gRNKRzi2W6ZYsH1iKR7E+D/jEkfy5cGZzwoFmhwG22k5MQjNCzu56Ttw
I1KC40fo/9FLLraUkobnV2CRAvjEShYN/k8YdyMBLFzLIRJk4Kj+493qma8KK8qh
TkuTeMN6W+PPp2iCv2utMnVkj/jzrrTkfiyjuTRRNFOgMxLOAn+rJCTmsqCW3zj6
h3vIrabqK/GEw74OfF7OzjEuAaxBje5BAIApi+sBIxBJKP+6sg0uudb5IQ65ifHA
a3gtse6BNK9XvdYx7QjMYlsilQwrxmCEklIVCgQTS5NFBX/5dfE/MMIJsi0pne3T
9SCK0gCfTok3WXP0K8LO3DxIP7Ioy31QllDb/sDQztG9BsnwfdDwmIGmB1MKX78E
0ZoLhaqPW4nCg5V//gWC1TI79PxFNU+1u1qC1OPeSfvBVW/jvpZUpuMVBK+oQaCE
WS+q4A3vQdUrL8S/vSk2472grOH1kImEpH3S5a3pBu05llcFXfByNwqXQVk7cSs1
VgdbzxK1oOPmMqlW1Ubr4cI5i8R7yz2iU+jz6b7b+LucLU50+UITiJ0vaMuk8lmv
exHNbnPTa6b1Z+tsOEhwQtmV6XDkmp9qwK95Rs3Thxoq7RhyrrnMSufkeKwNed/H
Dkwf9yxKH5P3JAfDQ5118AEbZB86Mhf0gcAT9kLGreKn01i+/Nt42/uB0yE+/S3z
Oa602oDf3WERKIsxhVCN9n9dMi7T9Szr4I3dhD5YKydI9e1I8Q2bZaspzP/YjEe9
1Gfeu8boHCKFbYu9wB4xmrOYTVdhAcZAXGwmda8Z3BoiXmMtOntcKudUNbDKVbjP
iyPV/D6NnmOp1nznUBbkqowG5NVAg+sZDsKw+Oz+W9RhzvCv9E4x4nfxDFMjJzat
Wxo1eOu5TDe6efPlWFyKmucY1YxPmYmhrenTIx6zNI+JWx7a9Aqv63VWMIBf84yL
4peGH9JBzv9Dt4Iw7EZrs+daL9MCh9GYD8eM274Wk/lVasygFtnYsl/7g5v8CB6u
1XP8941oQ4Xt6kyKGnBZ2y4n3/m/h329T8pDLR2U4Gug4o5wQ2R7AssFeHY4dKjL
Z32erHL79P9fAHNppStMpo0ohfDYPAriEnLxQNvFNrHc71w8iniS+AaVD+KZdxsc
0tV2wTPqHLtHBZhV5FaH2fPZmDMd9DVYrlCggFKC9iwDQhl0YU+wDUl3OEhv21VY
a60BoiifGfNt82bPCR3LDi5rVSQIKaXNRzjoiDDoFJl/jWztC47kDSZs9yPbUdnt
RqnHtbAVx+EXwMKSjvDzWNAplGNvkfZ4uL8SL83RT5vM7m37ayKfAsHXMM1tnw1G
o4LYb8b4YstjS58k14jEVh1K9LRtp3yGqv2wr2mIPl3gFf7NnoZYELRQt6wUK1r7
cJ73FhHYF6FtsJmHNgG/Llh/tJby2WjLgSjdWNFdMJYwD9lA2lPZ9IL6Bm4mcNTX
HE23DK5xpB7lQf9ZsSMjekxDlRBe1vDcphamAgagLT2MygDG8H0iZcasZQ3iz0CZ
LA/zwV4COBGXxUqFddxqMSphIiC+iS54aapNXJf3SNTt8ip6uj37qLSvFCLhLAUR
f6K0nh2RR7b4XFUkJlXSdxZVWhK0tJOuSykvdDiWMcsdO8HdGSaLiHNVvhGO39/O
uafrkXbWor0LeHC5GwGjJFaYwPpZdGTICBK/fCRECEHBJWWk4CdeHgSpRQwFP15c
NgjB5E/AS/KSJzBq+W+ILYiOdGzBVX+kq6dNGj5FeMOFJM4Pk1apJMdUNGNVyUnD
JYODL1RLRRmghGl5VY1wMogaX7o9XZuwrofxd3/oCkKFY5TRpCKEEyJz2qKhg7JA
oiX0qRt2ibhDQQxDvEIH8chdwRdU5fNKtBlxwNL0ReK1Hbi43j2bUEl18VXziZay
MS2UvHOso1HW4GkvfLefX81g/txjd4ZAC7mqeFbNexCX3EcwK59BtpHPTswZ2K/1
t5p3lwDLjJIkd/+py5bzmskbeOLgk2+COdhdjP52k4pIt42NZJEb5+WOEWGtYgg1
fpTHuU+aaVeG7T1hu5mqOLDM3W1+UkcOFSkot6DEzs8wHVGZwQV0ADnN9246MkkY
affq/XYkMWvU9SQCKSuHgkJBlzVGTvqOnXr5Ka/deJF/GLJ0P5iNerkPxAfTrCMh
pkSmGW7txvqQJ6txfm7zXCfmjv88xWh2Dtpuz26wrx7bZR9o8gkHc2jbI7grSjen
mypb6p5eoPTPm/d5IJhiEAWb803NjXkPIH2aALD/cz8azSJOKCS4Hq1JZMDGbfPU
xWCbAe5305kXub2ZdrZ+Nc3HBo54c9mGIYGDykUg/6wqIGYBLdlg/uNqPXQdbMRO
dM6k4xjMvRRvpGLUEf2URNrKg0vL+82DaMZ+f3HEvrhbePWZusE84lUZ7aEEY5vV
bFVif+jVZx+noqOAc4qv18agEw8T8YTkQdPYvYt28bA1svU9xTa73+MlgcpjMtKW
L7P4dSw/Z9yvwyxYyGWET6d6zMZnT750eNODupSQ7CM2s32Q7mCjkMVKEodmlFcY
kLzOqmrd/H6rO6VylxUfUPoElESknB91nJxLmTopPI/FVqrmDQXO4ZJ3+azHAjBv
G0rY8ACWxVtEOBzCQCPQOdo6IbRmuvzNbzUi9rD1LyoDJZO1ljTN3ZheP1x9cKIq
UzzbSJEwOt+xezZl+Zeh8Yj4239eEGEdS4072ER6psnWIdh2MrNI9Fa6KNqwSQ+t
+PkXV3hxiQp2wkI2K81pjRMX/W2C6ThQRt2nykwoi8O9PP3rTOgVmwhucc/WIrJt
YUiF9GbRxgiXA4PA8MaTxPdpmhIITOG4+X+m+24GALykfli64ulqz5mph+3m4vxg
yriMkYJgpdHVvtoHE5/MPdZpUIXmxlmEpR0xZ+l51UNy4Jro66/WhMqlrJL0orvN
i4E0yQA9titenax71jUh6luzS7+ZK37QnMAY0PsQkGR1B6fzU8enKihuKtuy47tg
V2SCvgTKoCvLLvNhq6cIDltn9GzaRRY3n1y9ranNZ7TmPZ0lw0qxfwG0rQhk3MT4
bUNsi9zlFb8sFutosdhak4EM7zm70G1rOYzzN8AA/LyYCPNXTt0c4PiX3o7+FCMb
0kQxhMOLA1aVVHDeUoG623X74/KsCYe26Ei7UBOuDDnneSiREOhFRrLxZvRETJy5
u4taRo+RGFx/TAFp8GS+qhrDGh3o++WAE8xEGxysc1LfQc/H7KN83yYm2il8Qx28
+5iF99OCktcwsyHSemX5cPmnRm3B9xccN2kfdpRsgmcZ9AdoL3YyZrhzg0RzYuXN
LwqIcv9kzOvLgq712KUMG3ZS89ooFb+o22GbpugMGzAyRooZc8OqBavGTFbsZ9EZ
sDrS11P7FE3uoc8Kq8/mPzslaNq9qP1vctYFz+3zQ1lD8hq+GvHan1oZ81NBJIlS
S5oVe/95NR4vdMClyvpy7up8M/B/FRz7d6XR8Iw+PTTVUjWiJgJ3Us0/Rot8iAAQ
A27acTz+z89IBhDOe6ycsfe4rbP4tD6avEewQOOauqa+QkyK4wn6T9Hwv2qO7CBK
QB4E0gx2sWRAERfQEcujFvMuY10aWuqNFjq/xeuBUW+iCQ5fMiP/WVlaFjEbiy5p
minL1lB7wq5Ok6to8gwaczX36fhC+kuutmGx0b90xpn4jisU2prw/k755vbLuZSj
JMW8YQgWsQEKlyDdM1eLLvckLojh6u6m9Ip/WS6VLF2mBMPY2ErLqgm0xfu/nege
OIdFjvXFDUiV5+0JptXMyW36Il1M1mn8QIICGnTHUFSKMr37gvw7ToWBJxyIVLW8
FOVqlBSakuSz/95MH1nop7NEiS+do3wii+UMJArzI5Ve2s/z6evRc87oxaFpebyt
MsT5WJzeTvNgouz0ZTnXKrQx6KKuQoF0gK1u8PpyEyp0ihJgtmnkWC1c6IcXTFan
ACH00F4zrqjmGWUsLxHvxTBxZv06TB3IXN4FdfmfI/mqKFtRP+rcMr22MHnmk4ZK
m/MQa6RDf921E1upmE1Ol1S0rkiCSRKNdl0f/6rPBttkbNfsFJJCHy3PlmItqLbY
ol3vm1IEWF+XgMeconTW0MMlZVzpDdtSkOfA00W2CG5EKu3TcscZ+2McMk869M0r
4dEHMs43TMmUhqGf7PhBPVrresZb+rhY/OqcefmVX5vvbyqBNU5H2xxCpYGTnPpr
kfL1B01NaDKMwLALrepXayyol5P7l3ORwm4KKzGMLrFMJexmA0rMHKm6Xes13j47
E+E/ovsyZiCfKaikb1pU8LrulRxbBzKsCk7lSOMTm1uu6ryn75aoqky+hzb6zHPI
H2xhwIcllOzU0/Y7x3FdAEEdpkR7rv1xIMjkZm8/Dg+aw2hbH56WH3ecfLuE1ogv
sEGcO6f8Z5i58Uuhc6Itveq860DXLDywWXLyfDozAuaySNC+iOewUmxVj7c8/zjL
WOEwZnPXq81rSaiZBL7h/6v1k2N11Ix4RtWgfT2fxAkeQreazZLTk8YmjAsnJxhI
E3waNrtmNPL37QNwcVelsdlrGXuRkPkJTESWu/89k85F7tjvPUQ0YXBVzbYI+qQf
ncuxoc0KwDIA9aptmCIHRwfU82m6jFuBTaERlnzR2RH2BZrEji+9FeK7L6ydSIXk
xqN81iATAXp+A3mmhdtCSE9n1nnil6x+3DoVNduWRYBmThah3yY8hMfZZaGa9TU+
SCbQsiW7sDoLvABJZ2zcYjA3LMHuvjuc7r/+Dw/eVvHWK1krSqtrFcjfOHaKAFxq
N/isuRAJ0Uy6LtT02EfTLof/p21XUl+y71nPxfTZRWuKBl6gfkofrkRxEnJ97dkn
cciakvAzImq71buVy8jtuAYWFBkj4C0yjiMEWjjzicxoszTWz1XnQm0d4LZDRcZ5
O36w9ebz+XEFdXRbYZYk4qaZegYPT9TuMlJ7st2hHChLKh8vRnY3x2TJVJLcEfSk
C/3UEhq2PQh4hxsUkZZgp5FTn1YQ6zKGrlb5z0TtQlGwQCfx0q7whMDlhFQjtH5c
vsdi0/DfDe8/u1Z2Q7hlY5ZpjPLHYKKW/haRC+LaS0c8qEewdEbjzS7F2TO2OodP
WNgSHwt8rJ19C+wKBFgcwZ/pYWwqW/WgVhEZFbveQRz+hkLX/CuTXi/f+UYeEF5u
6KMNIaPR+Dhis/O3I60EQHJuD0trq0qflQtXOq/KXzMbzS86OmpKzQ66rEleC6VF
iEGdsIpu0MeglOYThv1q2rbkztbBZH1J0sRPaIMq/GYntUn4gGcWPhyzd4TMhmi7
/Gouha+kfkOwrLehhEeTi7c1ifKmwFQBrbD/RyNw2Tcx3Cj37IikYxasLpsx76tw
nSaUzCjzeNODpW4Pyq/WV9zs5qNoNttgNNR1cdhJLz2MO9gaUTJjdVC3dYDJMLVQ
mFUfc2LKNKkmEm8exrVuDO/dusSIQaHLc+pTaUVJ3Yiyj+p6d96ZUDPQ61CeshdB
OYSDTrRCoQR+99ofgwy8BSshzRYqXbcxtTd91vPL9+mLpFG/fVM5m0LBiJHl9//h
WtMU1AQh0lZ2KNdBA6OMy8bSUpYSu+rr99ny7n5Pl550iXe3IGSZJnye2LJx1EU9
xE5DiSxncdfyiE6TmK+dpWHh1IKOEJGUBBTRuUsMqetVzu/JaDkXK0vKBATGWf7F
Ko6aCXp/EDcZpyd5XNmfviyZET86hRDz4SJ2m0+mmn1G+W0BlYWAp3xyiH5z0E6a
uPgXSSNOAaNZdG3yX18M5VS5USCP26OJy/iRxQlZNgriNSVTRyIlQf93lkDirlu9
srL4YjFqxwK6mfzx3gtxDFxuIeFj61W1HV7m0Eg3pSijTTscqu/wA5YoV8mjympz
oSW0CPT28JU5Ryn/9U39WXSKiiPHtv69k59JhmwW1jFyVhs/WBGuJ8EfRUMNk4QL
oIV7B0/JJoRUVi/S758O6Mdc6vNvmrZPsh+FIy5cfgSaXTOvs/s/AIaYn2af15zt
JZ2iT/496DaxuKcdy9J+hJSqAhl5L3FcpaPvMYlbzaSDQ5zqLPBtsapU92q7EdkM
/PebuTBSEYLTL/7OJj6WkIixVLoqK1AjTl+7lvVoWEaCJpjmLR66ytc6KhZTxrM3
n6OwUdxVOOw7aEHEOLJIae+RYQwZs8QUaNRZkMj480dP7gt9mF/UEnkxeavR7B/q
dMqtFB/pQDqonGxVHJeXDspdEIsPpGDlRHvN2LsXIIlyEoi9X73GlrtU3IT8dwwQ
1KbdJI674tD50EOmSHILleju9oqGGOjAV+OUMfLPaAFRIwD2BpIrC7uZY3E9mRRF
yuWqe2vop8GTBbTtODXP7h18NxM8BICVY83wKxQsoh5YXqU0JwWjDaGMA70MYKxQ
1qOKwcRcVOQYdSD5Y9MXjwUV9ilXeCVBh7SNkT9Tr3QrjCNNbh0nI+XjWam9a/jO
6M24gHrvJOx0KEvUzmWvDp3IZ/+yUGpZpP9jTFBazpuuOjkTm75hE9NnnHvuJskA
g/zkKL1PlmneTMTEDROp2mcCQrOzKhg6zw39q8waPbhxBrOTV0YQI0PRrDbtbDcs
w5UD8+GxcPOv4TGnbBJSlyPnjAZLBgLdcZ2VvFQomrFWrJ3OtNvaO9/KnOTFlWiW
R40r4qIXvHbWAI4mC9yblNLX56fcuiNEyqWjhspTujMkIFQAotMTvPa1+nyKW0rp
KHry2g1LX1FvB9ehfAhunne63JiErY1+LeOBLkLfp6QIbkZqALUr/TQU+FLkBXFn
1OLbyryHEixRNmOLlJpG/rO9udYEUXlqmBXCtVJtFwLFT63apJoogpwrY/v2yOpm
TPF8KkDfG70m6qP9i3q3R9lZfkzc8cIc8H8uHkfTM4CX1y4i+Xdr135tGw39Hjm6
shVaqCYOYC/LvWi5+trXsDrRDSYUGk0/a0ZZy2A8hOHzeqEM2Z3S2+sVAudARha9
iUXrwTpS+YpAygD+lc2psBBN7uFI9CKGe4f+++kfZq2hDgp0VHEb8ADHxlOkB2x6
L07qwSY+j6QLj6zzJNxNVoiXqIyX2UL65fOMMhl3iJwSEYXQ+exY2xfs0L12+2FF
aewideCX9OlphdFkIAYvuj3bzd1+GAA+XngTAFOraG/NWU79RP8BCfsUYuTdkxB5
T/iM2N1yqzf5pt7aHQ51QSF9QFLgq1Q4Bzu8wzz445yoZa3FFJgwy8SnaLHeogRa
w20Y2uUSqKCtL2ra3XF0AThghjCXsFI8nPdZNhjkURzoPCESvEjsbwZrKeln/3fU
N8YVrl4t0xJ4jiqmnlxOuMYmyL+iKy2ZEbq4YirknrtzUGtG5UygXpVstTbai5Uc
mA2HEc83rcCO6J4Vaduc0yta0yX6yqVb6d1K59xXbzEZZ0OoDT0e+sIiUEM/IZud
rfLk7dxneD4JNg8nInVfoWP9V6Dp2yhMNQvoNjUtRgFOSCPAAOrkA8R/pmhsqDRH
VGa78WjgebStGefvyzY9Ka0N8uFbd9u9gR51trgU7yAWlExtJpkb9JLqPlUrOZZQ
/fv2chM68AxgPDB2xrUzoi7f3YEPuA41rpRTkz4WjldyoPQ85jQv2yrWc1y9EWEe
d25w9iFOhsnOAvYeepslMtAm7eRbLAea6eAiW51Li70BjyQckjRNJsSgm+2La/TK
/2ly9eV2gzYiceTs/f6iVYzMROiuW6CPJZMjtzXNY7m5hTKWh+wqLBBerB5N0AhG
gYZLfupdHGPiA+KO7d/P/UIKGlAPnrCyZYjJ6cIo6A6AOP3iE4H76LNNo+Gs1+Xd
VmA47BRMVzJkuRy9BNVX8sxMNCZopjAHUIJ3yRRsj1Q7LiBPjt7zS392PC0DojXf
8zYyApjce6oS6E+85DzHuVCi6U8Znw5h+2SPTRDr8C/qj2VP1o3m3SHMECy4b3zz
PhsiP8ceOEQTy4QyWWxCpZk/vqJRubK4sOzFvj2It4oJpkeLslpZRZopxUUnQ1pZ
50fHHptg+OQHUW1zCFCWnu0UcTmf7wEZqBBQ47ers9ejIQm2sBgZ6/dwX17sw56v
bdQoyukZPQaIrx4UqSLJj4Ej2PK0/YIG/XOff3USZNwkpctH2A9hRlu6s2Xzegc2
VxmXNG+xoXi4mooRbgw/HCDEafUrJdhDVwwNkBX5ekMJlV8oCi11S2SGENUv0GsK
VaucHafr+otUEtEfgvRwXtHTr05jIvEz6vm2atlmOtkOb81ZJ19dCctx5Zf5rX3V
9IudFFQsIWSR3RcmB69cHU30ShbW2QMY9r6AGwaYBkM+VL4DyJDXD1m6IkGrH7Z8
fhyw+9rUexaF0J55+qOl28eGyDeXNO/9VrKC+QPgIAC62Nntz8dlBnMkPnKG6nNs
QJIxP6tWM/H4wrKJ1LOJ2seSUiY8t92dsTmWziuEukW6LTwJKTCPDnaGDBYgXR2m
cvll0TU8rDJ0LAwPBqRUPmYp6/xn9+HWop+36PBkUp+U6FIbYDH+fVw88cZ0dzkC
OO4AsHcoAHHpGFELS9xXa2vJsraDgkZgbT9iknPVjoAWs2EcBLS2Gs2bel18znna
6CViXubpqs8hSHg1yAftsmYByeoY0SpFOS9ZhjovPiJrD9cwh5/Ra6tc041D4AgY
aHRfkrDpHmo3HKJm3xUKdk0S89XyGtmCwFt8xygjyqPrCkOB972hOrcmXHxUuR/B
HKjRh8IFXozWzlTou/I4zRROAWkCOixyOZ2b8tBwbWzNGMmPLd8acaucep1WYlGX
j1GKIcPfzZM8k+BGdxNBV/UkOzyW8FI/Zh8Df7OQp87SvKWf0oKBRozyQEaYVfAq
rL0Ljxpwx9jMsWc6AMrl6oXOUtj8DmezCpBpGW2yJBZSleVNNpB8Haca4Wgq01Wb
4c4FV8G7DbzKhU21TtgSaYFMYme2FNtI/3poQ5Y0nWPctP3VaCS4Jqww60YF9KEO
OtVqtT8/7Ge9BxLvTU4z/q32smoUcoB9swyvBeYTMDDhioZDgzeQInjcfkPDoMK3
QG86wmpDSD3mkAXREqYFJ0RsPcOjZMadD/uTaSdl8X5yCc7hkpkY7a3udql2Rxld
blixF8tNClzgjo8YYx3gpl1qtSMc1SZ+MAKpHYUJteyNWjDcrxlflYDiogPftYoI
L5ziPkGO4zzsjf3XMtOuCywJj7OzGuDP1P4owNXL9L5cNtsgBOJmHxi4upBTIOz3
zFJxNrhiSA8xG44Bd3KcrdaOHsnP3DMDzXl43B3k56n/jYTxJAXjhp3SDl/3JZvP
Q/CPDMPYT/hni1asxEl/k9NIp9VeGqNq9EaFfWyX8GS3py2AmJEi8EigBpdaREmY
G2yPdl7+td7XraPKrx5dyLf/sh66f7MWdFDQ1bhAHeKq8cHzCWGLcPhXEbFO34Yx
EbISfNQK5XlQmDbzgwZyuqXDA5dntMsHqIuQbhyIJRjMtM8Je4x5PfoQ2dH7JZ9H
zdBZxKGFNDHhd3Xla4F95gWkyBOO24yiluw4w+xk543wnLnDSyjcXc/78W41ktWI
9TEQrqvD7jBjao+2Mu8G6JV1T0RMyW6u1P2nGaC0pohLbzE76WuhW4qGHSi8PXU7
owJs/7DaZDBRVDYnsvjUKskVBCXXYJlMZ6fLYHd0n22SCK1eLlcQuCCH27E2afu1
sRYkx8kCrmpfm0LwOZq/1EYSXGRZeia4/SW79kgbpaW3MYj7AK5tSAgQRwys7UUW
y8WyhYDrkL+N/MpbOK1mFJ/PJkqgoK9tiq0bdfJZ08FSXtL7lDj0Qf9BoAH9dbx8
hREcV7bgxopJx0ulO3NBLjTmrqgBvaN3JUBZTnsLTyqGKXqaEHaD0qIpX9YUOd9Y
q/tb5Em66To3RjHaNYHPWybIjTNdVajZfFbsNkfrhBnTGRKbBESzOl6svSTDRXEG
Ft59pxHG7jJM+vn7j+lGYJ1KLvnHnLhx8ml+2kTQgAoGHvHvwdztV+2a5B0wtTuf
j4nlrlZGJz6IDJ26E89gQpvkVB+b7gFNupxGezqwYCZdomTA5sfwhn2tkEHLz4ms
JVHiF/f+Y4Wx50MPlHbWJZYqwWznZ74fBsP4Ci51UmGw0Q/A0uq4i0FR0r9keE8y
bus4lrkkZQkzUVRkY0MtIzBSjEYmLdt5H8jAUporKVgPaUjvoewBivG7x5VLdPDF
ue6GmPt7y3Fe5KyQarec8dXyTxELA9klfh5uXFcZvenjPcXK6coYBafmcvmnxtXD
mVxmIABZS7211OLWFBKa7sNLNKefEH1u2jmHQa7OE95lNdkSa7EyiohT+Js/llU+
ESc0z4bohge/1XOPU/jO3E/mOKhCHUHBo7BUhEDLR60ZNVXVM5f89dJKfMD9ovqh
qPp5g9vewe8Op8AQD3q6MFtTPiFv2IxcBJdEe1x9UFKbi3Yt2QLStI+hgqKYQNtE
M9VjjHswIU+cFZQqeH7zE4hBKLoLX/dC4W8PJh8pBqai4MGaAQIJtHgC9oFhJcjI
ra1j1tFZ763LbqEgOahVH7uJ5wNfK9hDPq/mg755ngXfCD2GwB+yktLtUmBRT8UI
lvn+/lvMenLmjLxmJGjradlXq9e8bWuYjcmxtZ6Eova4AUSbjacvIhyL6mtWpdtp
wPANGPxGVK3R3kYR9/lXPBmtvGHdatJZozD+bQpCKJVHRa5cQMjISKkBb8O8a2q4
oVsWaSn9i0/1yfylAxVKkeaH+vZBoWrtSSUzd+gVk4Ub02OpNn6w/U1/GiQWaR56
UOPeyb89V1Cx0wDYb3TnQvSaHVqfjNya3KK52KN0AwMtQlIAu9iP3nlVM6BSB/kt
Msj7gmldO9UfuecidIDJW+1wIfKDDad5pXwWDSjpqc8TOOOFTqUXB9/H3oaNiPnM
LVY7T8pXL0KprVL3FSf1xYywE90GCjepw9KvY1sHTsUPLE6UbaP3zJ7p9dZQHClR
cqYeQUfPxLqouwBTNjqUh78DqayWX6a8bYRTigozSbNBAkGoJ/zoLremYcXNnAEo
GjL9TKJ6hlBJelqtqpINEcHl3Ceav91GDgxwMt5R6GAfHxwa+6sRupbeDZ20LTgo
XgiIeugHQl5kTTJlUcLFCvHAJUPEQnary8neluh8DaB20GY7Gt0qLIsJUP2mmMTO
O8j6mkPOO9fbloccIP88QPIWKxjk9pWf/GkottdsC+MTxlcj2yKVyus1Q3N6L1QQ
a5CUZYeRrj+To0mPZoUJ+5mlKq0m9VhOY0VsaePY6oBf4pI3yGAfEJtviZNoLSqG
xNMWZuUUBKg/nOy+OJaBFZMAi70PzM2uUdFpZdEgbu3gNuwlZ3t2G4SCYzDWrFw7
GElAJX3DzjGXnfaw4YCEImpcEQC079fNu+VByDuouPChOdOgnweoeJ6ART8ImZwC
DHraFDJTJE7yQL/ygAMDbRq8aN/3Sq8F48IFc/kdtLOlTtngUpqhYiU+kU8UnRom
5QpY483umRfDi1lM2IkcZEvq3C+GZzSDe7juG3uYYc0jU6IM7jD/tFkxnrRgXmrC
DZIvYwaxm9rGcePChNi0+BQq6HhV3HO+FDN5jMBVrcTbuRhL32L46sfev22f8tzw
ZUt0bSI85fQxUuHtfIh43Bvzzo1HNXkl0RgI8mL3yEJH96I6raWcnV8/CVd79BZa
n+xxVRKuRxUznf4rmZj5LqsuZohhsaGckhqmBss5ZTVAtDVyszYbOE/wzuKRfkhS
+EIiV2AOfXLrXxC8HPrrSVJO3ttWbua4vtK9gobzD3r7A2whp/ZQIRIdFtdfwhMz
ka7pIoKDACFVI+m06Vi+456L/XjK/BCVMn7atMDujHFIOK1TAqRxZ4Pd/Jwwkuv9
bFLNlHpWxQmsSZWyPEr/mkUwpVty53+kwuAbVgX0USafoEtDxLQKY3Nt/XJAhZWo
ZzXnYU5fNf8olJ01QTIVMPmGxzxHPMq0TCQT3a1L6813qNBuAvdoVGG0gxWhay/E
tj/5B9JKf7HVz0uHSqipVkZ4VRMo5LEpRTzF+F7ShujMyFVbZYF3KXoDmqmUE2Ar
lcafoaXItNnSmLbwTTpU14Rb7iui4SbCWp0N68x26piwmO1043cqj47ujQeOdnsK
7ZtbqiBvTARFGlLvKYdrjfKdO+f0d3ZWMzpunzjeV36v6dYAkNvt/kNxiQEt6rqb
qpSy/TwyFsmzdTxStSs/O7RwXU/T1LFKA8C6s5IeXhrRBEoKSOScYN5YOisoCF8J
x0pDaZLhNvG4gNSE8U5lBvN41tY2vtTvjcP1nt+H2trVeYKkQU+fRYBxjsDy2muG
Xi+KIYAURukF1vKFFdeBkz79+pk5tA/cbNQ8WpD9h1whezpm1/8JxV1Z44+FEXM2
va7C3tIc/JmBR4av78yR/r3jzbEoyNZ/cycDGNDViGa+/7kfdAsD6URzTSy7f34z
cJq8dPuAd0bNU6Uw7KLhsITvk8/sfe8wmKV3WCtAZ0X1BI3DVVIe5vj2J++kqZdC
lDDyhO1EYfBRFF6Oo9eoDOZkQFPiFIywf2k0QTJ2Qwk3eiBpVlIsG8hf2HVtL/GF
eLefvIM+GypvJygLMOLnntleF+VyXmy7barfEyGdtbjetrWQaibak0mgljB1QSmW
OpOZMIW+Od/rD/w3sE2h2AExBf4pDEPYDigls63/xx/UzeaOZD/enVCoty8NDUgB
X9CFdoOx62WJoANZMutZLZ8Kn5iLg+f0nPTYACYhHOyYPiwX8fdP7eyXO9XdwLA+
IfwNsLbdz/NWFn6QqKX7vcmjOss40A1XwKEcH9teU671HvfPVU0MGlxKh3xQ0t+o
56Cjd0lNCUvLlgEPOuJkd/pU0kQXNOv3kpONkDsWNtRGt8i7CEg/6HfNbdZpijfd
hxpaQiSCGU+FL+UE5InCmbmYGkC0cIogVbRog70TvCE+vmtYJCbcaw2M2prNQhlO
uoHpXc2XzMUvtaMblxRhyeLuZ9JSrz9hmSscWO12Vh58olwCogJyDWJSxbscPk87
eRTu9dic9K/s+zz73Pa2w1xe4nZNawtovFQkyrYPATYFsjiXDTneus942wIT6+TL
yD3aFedP5wQi0wQ+RYx0YHU17nvjAm1FjuyLJaSIlnj5i2v/RekbpTs672fbT1M2
WMRcyxrw3kxviH8sNWI/hoM2qtZ1li2Gkfx//cTvbk6mQ7eN6MnAp6MUs9Y44pRC
mI9MmMTDRqj5wImRnJeWUkOB0uGnWxuHBbnxtTsnr97eWVeqNWX6CvzBzT5mH5nB
i74SI4lInttzhml+ZgB8ExMym6G4NV/BaW2XJlqMTeJWmtTX4IJ3VaSfRUVQfygz
3CmYNjSzkItuJ8UeOC7h2MOcGDOC429dri08Yq7eF2X91bRGTp/xJL48O2orruxZ
7WlxsUAVPKx+rTKWa/IgQOc/O69zcjEQ31QpMEF2D6XvRi/rDQ8Yh07BdLX8H3qN
DhlX6Imc4v2zQT6mIax4mDqC5wsaJO0L9mO01NZ7xVdHoFzX6jMPyAs2qQX0Uqx0
Ajo+1oXEnMINDZd9uTCU2iWf0mR6hyWkz1ZmRSM8QkQ31nr+p27CN7PngJ5G82er
B7G/AgzvkxDBAca6IlT45y2W68rAcJzUgpI/SDSSokswxMXkFIMh8X66dUT38Nf8
+p5p6bQcdgYYG3LhT/CCzht3iuPStPzliZ+ENAYpJJoiRniqmo/MwiRqhEUUP9W0
nMlVuZtOVV7kyLsQItouhfjk7OXW8DlgFvMCGz9C9QCIxovjOez8SA/ayGgKHKB4
RZRbCs9Qahl3FxrGIWCQlm1ZmenrBsc92lkICOhJvxjABtswUq0uV4x4gSvD/2rX
nbjTIKpTgJuYO2iZJrVFzmDf9DzoI52iKZEtxL1J+xdRFRSz2Gf+vdim6wY6sbHF
DPVM6R0UPalHzdKkOWR6RpTFa2UeicTV2a/k8xgDeAgmEqIg1F1X4aV6MvqQ6AmZ
IIOJGa6pXrUWzFzJ8f8Ktblyt2XXWmlcWM2IkHGKFXHXLZSPQBcF2PU2bXGLv7G8
WagS5HFvwk76F+NyYJ/sTaK2dD9GfV/vz1k2y4EPN4GWlschm+am/iI1v/8RHK7s
6lfiADjonbNlc5bmLujwKWGP9DRx6wNVFflDjYLnT50LAxyvmsGJ6amXp2h6Q7AP
pHp0vfa2BkV/P6NIJjh0bB1CpIZ/L1L3jqCbfbbJJ5Hazx6bLNfTwXwquYQAJZyN
G4S0TRSDi/McDkBhshWJd8BC5XvcvGsAbiGzKyVQkLNxgMjMzVFp4xnlZqraKXw8
sCTMG3UiWfQBMi19Ft5g4Vptgto76arAldO9IepCgcCM1jl2ucLyoeS0CtMSXzY9
NVWhSAb3E1yEJct12CPJAAiSiJhaDmn+eW1DvFLmm87m8/BJWRQ+4jAGS6Rrujjy
lgnNGcEHGZDOV95t714mks0Ww4whvMIPx6Ip+P7Knvof5KIbdc3y/af3KXiWZVJp
Nfetlatk1Ec5Sp6oCljMwnstksnaA95Y6vVF1/YDzbu+qUYUC8Tks4sBS+KAHYNX
od0Bn/pzNHe2EnSmAMpuXDV2+4nF0U5WD/UqEZdEp0UeC2IGDLj6J5STpdH9OpBk
dFCjIKEjktnq6vl6aszAqEJ/0sh14eitkS6Q/k6kxW0yOOYSzjm8UiUuw+BHHUCj
Q9O6BThyzm+Jtyh2UIey0ni8BU4VBEWsru4RD8MTOPvAtushkNscUt0IYUodQuKv
qtkWoCeFc5BSe/tzmbY33rQDYVN0Ib+efWhYxuE9XkpoVAXpVx/feXPH8qYk/GOd
NC58ojrd5hE8vTIwSN9wN8V1dVvgBtMUFkli/K7xo/FFuCiMcEhPCqs1ChafRXEE
KYUz29Y+1GC5UoFbXVAh1TdeYXCI8vkRLwar4Orh/Zj3Ij5B7NENFDvvrF7eQ1Ml
V2yKQW7nD+hQBDuXnwpTDSRvbUhVMB4sq1WwIuL0WHxfBCEDVRJdxjcNgSGeGR1o
0LHtI6zEhsSMSiJreS8FsMvbhuxKzm+dMREIF5697MzNXLLsAeJCKXh97t2I1oHB
xmiqA1G/w0ONxnXw0RgoR7fmFHFyEzH7TtQfVU3aIsfd0yNaoTFwTfRB54PRqp77
29SSwVppzvBhsxhwXKR0InhP7PLrVhNxG7yZRfNFA6YAW9C6U9ucM0BljdjQ+C0x
3FVj8UTGiDTg9AeuPhDTCI0NE3oY6qMt1fHFItzAGaOHdD26KmDr5nzbF0sxE2hi
bcFhPPUU4Cc1Fpz8tmvaJzbIhKt1NJ5lR9c/7RbMimpbn1cFxoenpIJO8Ax9035C
tIyHT63bPZajOb6GhgvRueRacpRT0V7MbNt9ELmn7eLAchgtNt/fbwVLoVn1KU32
ragRDFqNp7kKzHp4/2Rx/SBTBwdqqJaQ08BmOtHqyxtYiGWhjiNiZAkjI65ygmW5
QexjXncAf0AlxN4jd3+tkI92dAB/XDC4Zn3FOErYmH9ogTNFTUMfDF+EKNvRZnUM
EoTrBtkrj33TbKGfvoWm+zY4iR7ficc/iJ5TZCgXrhHRkI9vDS7sAik6DwIct7P7
nIgZpJ5+7LExWPPs/XFGs9lYEgYHbSWWt0uxwOa/a9PX7/uNgpv3YLJcQ/zIpyW5
7FO9rgZvZFTBlxjN1SA9QcwJpSC2Ur/sm8BIHct2BsxN7FZfErSxL/wiDprI2GWQ
39PY/5s46nJxCT2YtWTKEqSb+X4pbap18EBEw0iWZJ9Lo/e2EpzYAwf/gxUTVGSX
6wX1mapNs2Lq/6kAC9QO3aEV0Fnbncvn/O2M17k0mBa6axVIOgqyf0pzMOUrXGYc
ifLpwHaL93mgfXX88KFIHEVmUp5iAc279MB0tczSufSdoyDzT/uqnObOdTj/PahC
lg+ChejS7IhWKcOWtwEuAXOXeB2BC1Z95jDMqTMaA2S5LF2lNOgCobrxsCJZom3B
kK+VWFmogfO1wDQsgS47JNY7BJPcE8ta/FUvk3NnwTK761jA7uPFDCWfkV5AonlV
FMa6jhmz6RozSMm9NpDVr1hOIYWueK+gWJvVhsvXYjzwY6KwUyIHDUGO97gutt6O
mbEjt2CjANuVeT0o36jUrYkn8eFNQOtqHz45LBx0n/aZZ5xrXv3PRhop2C2xyDWD
l7chUzr7QLCuv8dd4AgyKWrsnB1TBIKny8oppvqToOXMCPyusKTKfRdI0306gU+f
uAjl4VVJLfELs9MNg7EwsX+tQeFyEMbes5aZwiNvA97eENdCA39fvv9vJCtH7Tez
ITexg719u/vTa0Uf+UFVD1XwpXK6J3Ps/IsUQ2Rb/nY1IHxyPKn3MRd4Zb7eN9cS
xjji0bZZi9fX0rd2TmhJ33ePn8qB2mc9pK1gBF5uULJXSF9mwsnjeV7uXh0Np8t/
oqwgTJhlW77fAdkUAqfRqtXIIm1GQ23rqWWEuu1dLF+MMOBw347fl62T4y0ci5Dq
LDIuUkr687IF4wbt75s9J4g+BhEQW2S1CdaJmVdHDnrEq7a+/YZYv/Larxg00eTd
S76lEOUrEEomGsI4bdcUje04ZseTFMixr0UecqmaI0huUu0d2wxL95vOuuKo+QDl
VB8qqR6p4Owxx1ceAqyTIg+ON52V3D2H13HfCyhih6xSQ5H59x2q5sPiXH7yDb2W
8oIGk77coUSk2mYwhiIzyKosGt7S+8SjR8QpZvxaSj1xEn+Ay0Q6nH+1d0+LPddZ
3RHSOQcW9MkRlkSUraiB1cEmT5H3cn65ECZLwmZoF9rhyH3E3t2V+afNrNm2H+4o
T5naDZ8qdprjqNum8AjbDLusp50Zsc75a/S7N8/DryRjLCsswn4gcUe0TrZZDdAi
Adg9xzSlq8Hgqm5u+7wKu3J2pNaejjEGJ+CCgh67Xt4URmlR5C2ieQ9/nyrtaPDz
ybriEiFJCA8PmeOttqRxZ/9yNf1ZluVhX/Cg7rsBzA9Dau5sZgHADEVBe1xHqlzd
7CUqlrJEqStjV1EP3VluLLlvxvHhETlRfWQfyOTX4f7CkAffJM2EDaHdd/DW/IoA
FcqttmaHuesryCtwrJPCwH9EMWpQepJeaPhGvMBa3ZmX9MzMo8ST1IdHWzj8t5I+
HMuDoRoMPEz4zcUhUjLaW617/lT/BSODxBx4RLun2f/EZ/qwghKUT7oeR8G6t4R1
K+WxZrNq7jKYqsXggeJuV2Dm7oM5yt1eNHfYtauwg5yIUTOfyjmg0juzs+avg5BH
D0nhuiO/eGyTzfMhWrgs9YJJX4uIZHI44f8gPfqLJ0Brtmebi3yQDHB0m+axgJGX
kKaKTKjvvB+GN13ceG2nm5tWx0byKF896Ow115Q1Rrj4mk7yxNnxl2iHZuxDw9lJ
aN6SNlVJ3BMRZZibt+NMfVVruFihbyA0Y+S9LedjlYxs3sSmPxoBaodO/r4d6QWI
zLER6su+Ee0ozUEh00sI4l/5nFfQw4+vFs3zxdSrA6Aw8UskfKmaq2s7cTrjcIKe
QQx41O6FJGFhzRk3AGn0+KRhXygIDP89S2S/8oQP7j/N4xyiyCKI5Zf+ggwm8l9K
19xT7isZp35S97LdqEzC1ElgKGHO4kyt7lmrBc/ouA81nwOtYufo4jViuulWYztB
oTRhfh7dusnycHB/nLhuKaOYj6nbnU9zhQzqW7e3SFKpPw1l68pJHNlZF0kpsHZ0
6uopFCOh+L309qGayfpMeQ0XPbw0kVTEV5O6KlaSmraKhVqvHSRYpgVgQwsdUkmb
QD32tyRly+vTqajHQNb1vv9UFSAiblArLTgsXi9m8Jh/xJ28CjnOpwP00Pt4IpEC
GzGz5cWKzrFUoYBqT3mkr9NPpfrBatmdqeVjI0SU7U/0tx7nWmYEsZM6CrKB1/GU
cYu3sEVWxdRhCe+evlLfU9+mc6Aap/tG99ow+wfKIlFfQhJvbIVDmtmb/jaiJcup
U8eEc12oWX2iH+1Hlzga4mG4aK0o1PLQz77kVnqigVZ0pFdwoZCT600Xol+4CcVq
D8XwC4D8m6zcqyJi1y/PQNqYCtER057gnBXECah2lKcH27qpk1w5NsMwA9wz3RrD
PfIZI6nqMgavBgWF0p3ChtIkuTWYLKvS4ZR9cGyELE0aA5L31iuQsjXz6H+P9p8h
YSHWAQnIMuF61qrqufet26awvIoMxe/eWRscS9Z+/uL3RsBbElgM6DNrz6Y0gJAb
yF8jJwgKg0ZQl+SXmB8bNdA24BlH6NQGvrxSxv74eeaYyVf5yzs+/OCfNeejRR6Y
V5RCpa8wxrxy4AslRabCjUHcNGup2dSk9PuylOAlZZ22CgkwKWwblZYp0BO4zhuI
POp6ixr08pJSTmTrWuWM8ct1ea4s1UTFuhlllvEfK+zrRjKLvCuGFT+99G6ZHPZK
/jJ9+YSavikAa8lWT9NQQuY1PT5uGlQYnWtQk6cVfYlc9wdDPmMNMz/XnchUT3F9
3SV+eI8ncvYiL+wEcThzuyAoaYDkdagEy2FnqM47V/njcphDvQtdMdAjWDbQJnTV
gmYXq43Y4v5ZvNuTLOhvK8iERxpkIMGYIN/scMlG2trJdxF24dp5ptYedGQnczrL
+twFz8PH49b6MQaOV0Jfi+ISewB50Vo1OQE+wgPQjKwUR+IHoXhybdpfvUJWMRZJ
URbD5RmCKJ31bq0KRfVrArADFXSjaKut15mp9s/kWoheFXfn9rGhbcei157++oWx
fuIJjLpmXBoko0tb9o9V0iCWXECb8OGz5C21s/GoO3Yi0wO8vFeeNMn9Ru61Peo9
B+k4U4HTU8craGVZeLzJi3PSgtc672e03Zj3UrBmGEv1yLaOXLpCFis+qNW0p6wH
Uy3E1d6tfl3FjySSVTgxpTe7jP0y5cXHiXi3y3Qeayr67Wh9X6dzFu9N9qv/dItz
BAOwRp0EDhgEFe2fouwNBGcRBOSOm8TL6Uoz7PNSzkZ6d6CanZ5yIqRv1iAqqhiQ
KbIYB9KjXW6TClIusUFFeTFCx9CGqgzB18BdoMgF15vwALOc/klDfko8cLip/GYl
/ddMYCAOmxHbUBizNuhUujgnl0SHfAZGZkB0mNEcNfwM36Fm4lt+keDySxcBndv/
9A3yeAvdn892pdluwu31t+yvqKNMLkt9EmHtSDVk3jciNAEdeOD5yp7M0y77O0bb
dko3ReKl67AV/Wv4iXD7a0KMWj9zc23Gtdt5Q7/nfqDvyvHQzS/isYMIpsAfOZwV
N+2KuTUtfbRINAgKELHrJSnxa2dqWY8XOkw8MCrDv6DtfDmqnUiuDpNo8aGvyXem
m2zlJVC4xjOWWToNJqjd6uvQVe24OpK+bxFegsXAHt5rCip2oypuZl3uhhVb1w/c
G6orjTsUVCOoIDzeCczpKELmQ+ecP9Nh0pCALCKF9NA=
`protect END_PROTECTED
