`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yZqG1Ot9zlsqjneSK9ApqiGWHdW3JWw9S8Vgwcn1aUvfYrOgfAxsuN3vTHhzATsD
DNoTOMJXvHyZ5SuZKjZRUvBpL1BoHN1svM5wGhOQ+Bcw+T3bJIUxOEpGjYwd9vsi
SvYm1SpPKZAkIv14yZ2QK5kx8KEOqCpSOr1AhKkmiR8abAw1hHkMC/WlBuKgOCXJ
P/tzhelwBw+UIptj4mXnkcnw8x3wna3U5mpsoIGh7fxfPSM2x87uMkzIQVmjKOtO
Uscct/i5x6zOZceqFWu7+Myy0O0oBR7oCxMLZz2M8/TWl6AmrQGxyH7lod3KxskM
CnuVVvhpEpavRRghO63EdB8X3cof8trq0mZdkWbd91uFEMsFAAi53rKMmqRyyreT
VeYd4dqvRwbBv1Odp+6QdBpOizvZkm/ebWMpfFiKRVUw8Ljj4+lGGgZChFXaSaKr
r2k2Ic+2lDPRPtmk/ffyJOROJeFcNEpL4piopW5Hr7kAhx/lYjUuO2mcAjoI7EKA
lRAttaMRhRvYw6KvWAkjpxcI9UGFtaTO0hyuIMBWeW9uxkNKwakzodF+MkRUhOjW
Uz0hotfAu0QRShoxtH69PHFs6OilFNddfgVM0XlbOqZ1jE7waTyKOVjuhnEEjgOe
SVnez3iHFJpPjjg9fc1XwO2CX5mAQ36vI9qEa/dPUSvoGXLpHoQOtDpUY3iXLhOe
ltp6rkZ6YkJoKtCrcIGoiFu4wq5ma+X3tm35g1jFnax7mBum4QAfhXcIoC3eIMDV
7dN2MdiPQJodtiL2jZ6rAI57s2feZk+cMQr+KHoDkStGbds7doJVvRH/UWWD1N4U
6QmNSlFU+c/ohxCTw07huTwq1lT81oh00QpqUKylThO8DjT64fM3J8yFcO7JqEEI
E6IlUpKPpaf5ASaPZWAcj9g66mJbu7I3WXhF4astsUuGm7M6/ywxZ4hIT5E1nVkl
BYakWzCA50tTWk9429f8QnDfR4pENA2NkcWgySA2XHnE58fr4wkuZHIAQjiJ32lS
srSXkQl70SGOaatUHGpe6OpHgzfJwR4yEhc9UQUHH23i6554XITqCUeti4A/+dI6
UNPzeEIX5CVwCQVX1kspJkG+EOxpHKB0rea2K+5Y3myQxP054UFbD1tq2/MV68M3
kOF0wlAj2iGSqXDbxZS9WxbvrwWNwOZCReptN0+m264oQFBOjllTeCqrQn7rC9EX
PueIN2wDgfMNAgILTDDsFtnehBbEtG4JWZ2R53E6b4TYq+Rmd8y6KgV9OF5CJj/X
ea27u0aZWOxzNuOEM8AJZKhTlya1nJ01/38BFFvqWMAQ/QhRPScOHd7Az2XPO9Hy
aIEh8pVNH3na415T9t41Nkk1v9wCU6S0662LQ+3HgvNwSvAXxL4ruVUsCTnNaUx+
pGZ/Z6QnJb8uo9JLHpmjD/bq6BhwEwB2IExhXm45DzM=
`protect END_PROTECTED
