`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hINUls+YRbG45XM4Fm/9dYHXvBGZfn7r0MTsC3qyfic938Bx7E4XI4l8cRsd2BoT
n9U/DuWFGELTTus2li/FOKQoiGikvMc78DIIrNVpEfKAt6wqMZa7OY4R90BJMMmo
YKOVrNxwFWLqykMYsdV7DttRKvt8DsCdDbWpNVqN05isjeVTnGndFkYPOu11pOH3
rvaT8Ngypb4k79p0ZJupBLQDahFObJtCN0QO4ubSTuwppOAatqT+ORfUNCn5rFTR
HsWrShXO62RRF03KvaQAJBWN02t/ksHaimG6dCVFj7mEDl6uIpo/MdtUZnpa3UV/
fEzpDDNx2h/tJMmiQQbx+Mkzm2h98lN/ldWzdHfiEXlTsJNI04CG6OnKRty+VHDm
BnT70BStf+Btl5vV+i9R/0lafpPFHlNT1K/hsNb4Y3A=
`protect END_PROTECTED
