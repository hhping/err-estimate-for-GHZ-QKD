`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lcbiKiPrZ7W2KID8Ofq9KR3RySbIoeLa5qYQB6bTMLYyVkjBnSAYF2wW2HfigZ0C
3vmN+xmPaBuTLpRgiIO99tGMO1rZeN3wdfvzR4RmGgNNuOZFCxnQfZhamauoqvry
VoJ50kHhwqKYBGE8yrPhJvlhgWHn2ZbavXbL8Nzupfb4WkrgCmqq2ZQsLaiepO6z
o6So4s2INeB4ewR09u8BnACz1RL5zSalW+hA4P80ecyrK8ttSvRjXCHB4PjOzo6b
aP/qXAXxyavwnEW7PYr/GFALhqHe/aFwCKmte8FJPlviSCXKJgBrPQG2z78QEz7Z
XJXFaVkEaX0+38/xoVQAFvXRc2RIbLN4kWKzTz5U5yIDxtlg4Gi53idyMvkjYjPx
KFr84DMGeh7ABTGuobY08oUT70PC5ck/hzjWJig6MkiA99QHbcNmTe5M71OOxLmw
EHRtwTWkyMuttrJcD3S1gyVAb1Lg7YQuANvfW5dxqoDNPS8f89xG/0tVa6A8JAYH
LwWxtAay92jR2Jz9/uZxz/sk+a6A8yt5Bqt3fP5ZjsX1YzBoK7Ti9QJWBWBbsIYY
RDSkfDqyccm58VQaXc/mAu/mbGGUaQTO/Q3q+NQDozvtnq7vjosQ6EMvBD3gCCYo
026RfRoIeEOlTQkIWPzklubQSmpihwSs5+SWQe0sOTIXi7wrsXvhhHiWC2BJ03XV
4+lUAHeh3eWoCQf5eI3m5FX2UTMI7ROtYPIhhmMQmrVEU0X8GC4U3PfsnsvVIKRf
YUC+G2kCgYDcoQA29m7W8C33hM8f7ynUlXBVtPPtuAtqzdItiXZW4CH5yl9Dp1oX
Ewl7tmT0aLBSj260sNJDpX8j818fmM5vHJhr+hhrVETlOUqm2m04xZVdXuhAwteC
A95ho4I7GAb88tqz7MRYNydxi02nagBwpNTcSWauW5DTA+z+TKgUAjH0t4NGXgVW
2OSLWbWDhhLcQDLqTnNIA0d8CxvruSs7hQl7Lcu32SzzQvz1RBJR5miqsXJ+5ikb
4pGg2y1Z+ggguO5drOnVi/yMS3SDeNmMyjgdHfDx9kf/afxoN777+SBPONwYcChb
j6fElK1KBSjn/Ca/1fYq3ABLVLsCUMyIGxgX2zMNZsXyBCXsixhpEiJv3l6cQXA1
obZFj6fvJXPV4gFCy57t3J7WfKW6GvCxel1NXGRiliUg0maJhb4LKmC0b8z3Z3OD
vsy/RFWa3cSIMxa7f8VcidoFKXPV/kTDyMaAvjdusdzx61l+Rf7HTPey1gXRu5Rf
uf4xeeNRWqHx/s94o3OB+XdQWixOOrz9cTS/aQlfiNRKc/j8oJ010CSzn15tbp6E
BlRqVBlN7vY3B0MQ5qG/iqE77UmZaRDTfe4uEK8UuoVuyFiKk78xlFsgvuVxzV8i
RU0L3weGaQ4FDPdfYqsHQwrDUxw7qs2gm8eGL8ih1YcSoJdBkmum6nDwb5vb/p8U
SRWH5m7ZFIac5l/0H/qicj9p1X/Z/bdTS+1W9smKaD1cEMJkBaGjvfJ+MMsYgjVw
xzCkUeX7TXhGXhAkOZWQNHgB8TvIxwhBybB2Hu3jO+L9MGJ/5cAlvWQZm4j8CTd4
t6y5EMYqnYCgR9NfcCmgXF0BDWL5yuA47IRn5U/1ryiJ9wAGGaT/jvdVwegKXiPl
TRiKNaaM7dzLH1o7Zmj8iMqHKBxvl0b4ucp/azEULYmXeUs6/9bTyCWkZMVfdZ7A
5V7J3LIBR65vCPgbr20uwE606ymFrw6QRMw0gXizGaw=
`protect END_PROTECTED
