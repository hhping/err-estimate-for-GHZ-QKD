`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5r/ktyJngM9phhaBTlXC/NJQQcgtQ5i5BB4+OhNz0zLx28FqdX00sLUl+WeejgK6
ueg55bSSB0EwcGwlC+0b6u90cmNelNgf1uDCZHu+Dm3StsfbkslCsHfzdO/n09QE
X/YcLSywRDnBuewDepZ3ogArD7hYFJCdzs/jxC79g86GoonfJEluYO+kzMgwvyVS
e5eHjbd9lIjrcTDNMB2aoBoCgCCmw77KtSUWgJspD+8fZhifMTkC0C1ORg7QkoJx
AJsYiN6ype7jE7nYIMcNlFbUUxSapqqkD1QtPxHkCyXL92eMcSU/JFe5IP/l80hq
H/mInl2cApt7Yt83ie5+LOt5+Tj/+xAAy9m3CViV8y0UZJIdeSvH+uPKdu+LI/Le
1/BCGMzIAoTbr4Sf7iSb6aSKao+gZm+6E6IWFK1qQ/XNAB9YO9QcwdzGve4DKVeG
7fRxTg/uLO5qeHwrY4fgLqt1ZCvHDniirhqACGuyEvR/lIlgjNnxUf2SczIuCvMC
UfvztYtKtszteRyMCJ5rp5C/7umCU764ye6k9wSyRR6IXJ2OxkSl5kMENyWkMVnn
ruQXNdYVeiyoF2IPa3RStfSynC4K8ieBCrdC2UQCYg9AKPc4iySpj4vBNd/Dbu5c
bfbN2HS85XaGSXXX6QvfWZHTi0h3a1xUAGysVDYWt/CEJ3AHF8FyeyuSEwEwUddZ
ORpxdvX0MHI537meFXOmCA==
`protect END_PROTECTED
