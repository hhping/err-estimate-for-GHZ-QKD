`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Fn5s67DjPJuhYF8FmPdxpa77lhFFUFA+9TGpyrgzAIpQ/McPA7+44P9Tl/MrcrN
LiNxeqty2BywgTaZLmq072UgsuV6i4qnkjqvXzo3n52KDWS9I3wv8UCiIRf8fjsz
xINrDik+ef//NzgJbmkU4s+qsrsBk/X+DNO2fEtQdrtM2dqh0Cqth8kt1EfY60fF
wxb9WlVb7f9IRCIAaNX1WNFo2qJdRQHYbpMiP7mJY50kuT1HYZya4LCO08O66bMp
cLIcE3f02hne4ITnIren35Fq5ykP/9JSGlqaMr1bfkttAr5gK5Fv0FZCeigHszi9
qehIbyFQG6CfBhExFplcXCOl9nuj3F8Fg7MO1EbAqd8EzjNRDZ/EIr3W/Jsd3+nO
99Lw/PTiuADpj3WBsA0Y6CygMuxtLl/uECZn1Lxsn1jfxkNZyzkPhfF2y2nw+FdL
HBhSqRz3/1Qakpir7qpNHWYhVDiXgX3xCwoUEpTVHCk44V4SFHdQISTsKsze8gDP
xYuS7wkzITWH594t5GUpP+Vo6X9irabAsL5suUauFdkbtcAA7tELw0FhNN1ZMdVM
MXcZZN52XifmELCi+WHzgUFBz96otewgbWkj3/YAOVLX3NQtZPHcr/vWd4k26BfW
aJIIF/KV+kNZGuJY6Cr76B1nfGatP8Mg4UK5HQaGcJUUt4KpDKVVhc/U4tThmS/X
LywaOCAoLkfaF3tD1K1woJjVhkBhy39JUOdJRPTQaJola2dj0KGyAUAfzILsCxtv
UKkvwlQft/DzvL4TQZrK6AboWTelSplTLEcigCvolIgOoi8Qzy7tOH1duRcTvUbN
4vzu4YxrerL0PGWYTkfmmSQ86c9icbGn705Q7HY5v9MBqZV2RKqc6WdIgK80ZQmO
FRsPDUqneR7lN9cHmEXeN80alzrD+czRVZftLoCrO8gIHlmppw64ninEIUk4a+ry
Ms+1QHfuU8Hloh5yDkoCp4Wuf4C7odAY6Ywviru6ywSb3bVKJRAlUhO5sPCOIudy
oWYOEoi2YIi9iqg/AEwjivQAkSxdfHxjATeTRJk2mwAdh9EF9rvsDdvb3TFWtsNf
aIUDYuZgYVxCkpQA0gnSMWeazCO33CTq1d32eD3F4srYq2zyu7zJALy9DHvAfnB0
c0As1Pp2Xp6NOA4kvFs4RNK1/Xo8zRcGtxp/fQuHDiWzTWPRuMxcDVIQnmBX7Ftk
4JvZ2zt7y4W6hu/rzpGybLwytjdZqxkliwK9GqY2Fyf6SnIQVEfyN61yVxBVpu2I
VzAqYuVx4t+oZkJgzM27F6g7w5IfOA7qW8MC2c7Ut6EvJGEkVcSkwXTxq0mIkY04
NNJfh9HL5TKi1jn15dwNPV7BddXRum9c0jhHfszL8iyzhp0+0LtKVuQWdXZZKswQ
oIRyLT9225GWHtYZ3Rm+OKmU1WjzrY6ILV/EiHS/feldyKYvZ94Sh3anZBdMU6dl
TilaCYA0Ar9UMQ89Nlmy+dd2Im0GoQdwnemWkepFscAy2nm8mQYloeTtvpSxFfpA
LAJJd6h2+kSqlnWMecapUrbCYSfT50CTSQzW2iUiWSpQ2hmSCPzeZbQQaVvODgz7
BfiJD2C8bc9BZ1HDCgXAtAuwu+8i8hP0HuOSpUNetKiNZwtOWi5LqlQY/AYZO/An
+GsXlt9rymnyVGhTjJmsH7pWCtesHZUQkMmUtQ9O6Z8OzZxfWcOksH8Ss6QeNTOv
G+Tl0TnWO0Cm+DYGCPNTv4VfXlOfM/otUNGUkrsxpvAWoy7/Px+8YDpSx8qeR7PH
cuUN50fb4mqztnLeEefZ4DRYsBYhQS5yObOSJCNw6dkJy6SG6mlAH6ywUnY6YSXG
JnJi5ZfuQhQ7tWt9TI2eFsCxx+S/a70smky3NG63F3OSRr6wQyzl4ZT1LKE35ctr
q2u+JrEvYWl1GmzMeLD1QtI14j9FEPK+VWyRTfqyrARaHhNbFy1plm1w+kyPVz6B
1y2cce6sRtUfrtBdCTUh1jQmKFk4j+NtMUTQOkas/qJQuDP5Tk76lbMgDwIwlTxR
GtMzGFHf2XKXm69KvMb9LIluEugoM+9D5YeKaGbpoShg88NmdgySHNgSFUfjjssU
pI0b5vKvxIvWNC33H3z2ibtKXm72JwVNT99J2ScaurSHqw/q0FxVdxfQ4ykn1JgS
5MGHjXHH9I2xPUVsIy18hhevxp5o970q3vrk9JuUdav3Cp2hxslQUYKy187GUEez
hO/wy4mX6pKfde0AMOXpZDl4aI5Mi3+leyArxriwZ0VOgNJQQ6V0+S60dMw/vkci
r2qsPW3/mQRJ1v9M6xnOKNiMoDIoQdR3tT+r9eRaw1stCFsQXx7HvsDUOEpR7/eI
AqklRxPg7yiZuc9jUD9tLoxzfH/eWAdgrXtO43BLyIVgK/Rx3FXkscQodsgJPDaH
DZeL+q1zQ4SUlPpqClIFmLnkHvDrJ1gYaLt1hHSKYJryNu0gtNEZbDM2FE510jJn
pkghK5GOkt2LOlp9fYlBD3hDDF8w0U+Ju/ARvbNd308XaoI93AZklTOdf9oinAVz
aaD2Qhuoh1Sm3kw9kC/lM08c3UL4ZmuVxxvAXAkTrLjoYg+VzMQzxTQZ3VId2ibL
Yep8ijKwspqmBP+IfidXpLKrrsdVxBwsAttGOOS1UjaMm8YEdWIRvILVAW4X56Py
7garPiv7V3feVXCGgmVxtaaK4AQEoEkGRDgH2LexknZ1fE3D1TsK7z3Vi7601Q6C
iRBmuy9BM10TsMnJaTb+RWmeRvjjZhFbiSt3zQ0SRcR+edhOwNbuBFw6q7hj+Sgc
YMcxOAtiu75SjnsvFdWXSDU0OjxdZID3iLJMKjkTVWMqBpzbH3dopcZWV1dWyntw
AhlBlJZLmAFoccYW9DpjL5A8/gBSBMKkhzDhdEbPEsfwhvVNukb07DjefmnMCV7u
BeZnVBFDiuuoIP5M/OmvuuS+LzqHWKOORo1qsW7WAL3Y17u8tni/JGO4WrDKtSBz
hAGk5RaQBVXISu0HEBzHxAgCktTAB7msZhUuzeOqmMZtWsRLBlhCkMIKtXo2tuij
HP226ZCkIa9NQdjd0wOinA==
`protect END_PROTECTED
