`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t7mENImy6CXz2TApHF7k9YgmXXYvNddx9LFjuF7PIENi+uLF25CMa3FP2zqiKtXr
i4DG1xRb5zOO5bbIOiqFxc4KoYlyVds95GpO+2d2I1AbpIhy/2gky69LTOL4nWrx
x3HJGh6oT1xEQ9gAq2bCngIjom90/t63ymNAB5UUkzsaZ7+IbQCvw8HzQEOUXwa5
3ys6P6GRgRaYeYBbtmXHPSHVUeY7u8GPMLEFlVgU2HyzGXZr0RbXzkGpCb7RBnyb
wbJV0RmVSq24XLPCybDVNK7B8atI5DVat6KUTXbS1oVF4I1v8wkFFoCG9MomJb9U
u5Bbw18dD6Lsy7sWsJu+3aZ3/0NwOI/LxjhAaCf20KW3WSEAJSztfNJFYy8lwwFr
QOBqbpMDb+osFy5bbyZ5dPAx7OM1OMvQGNCOiPkaUoqe1qsolxav0bPiUDUaTTeY
Tk+bo3XJPTFlpRktYVNNdByPzBccU0DPS2QExEc3OKZQXQtj0GQXsdt+3ypQf46y
g48vIz9mcG8jj4r29LDu2QD5xRXN7MceCND9T9gZCgaJaEY7gn9v4OByJpoOoto1
F/0eKzvMzQVA2l7hqfvJov3XUeuPE8/nLfHjXv4hvLuhM6mmTYbrJ7Q7KsTFCfSj
JUUOeXpq/9Stz3FhqBKaaB3Kwo5IPQdVchzCZy+xxY3K5b+GLdvnfY/jM044oZaP
nGOL1vc7mZ1wh4bIiy+pyVxzR1ga3oxYc3PfeKCenxuS1b9wrbjejUNnjVQHsepN
IWz8BTGRlCEi17C0P4ws27+/r+CpH0U0odusy5Trl4g4E2rOnf/3VjO/a6FrMeRx
vztkRX13obb0DAqrd8m9kuQ6nOgW4XohF3cOiI5AeCwqNimVyQG4wjID0D62/dOL
w+vdQZEtdbhNs/D7ChTgTiFRttM5wZ9czum2k5NodSnlvXZcCfgPqwwTkQmhtF9A
5uQdETKv6BRHc5RP1OrBwDIY3GbPhTGwEUKUfP2uBXGAHhfn8Y3LVYaiSMW3az8F
2LCaTFlZqBFy0hJA92royRllV7Rd6Czy8aX5FNsE1UGBDFcSUxDtzzXHtSnltxmN
ATIRbNq8+PXMvNvrURDHqldlRlpS8WoSJ/U3HXBObhVrqYfGHGa00E6BWkxdNDGT
tIYaK/plEx1Fz6n9Ub8ZDDn70eAEL6CUlA3ZdH9yvqOWQhYrJQY9Wo9Fi8mYBZX1
4/ofg8pj9fBeKD5cvdc/stL4kO+O8F0cW0BpxMLu54BrTKHWWHUrrwRcNmYY9R6u
/A9NddFdULSGzdvwjZu6MeID6GnYozv3RLgagb8U2m/xdIzlFIwAeKvb3huo/Wfa
5n8sUq5/vJFqKg9Y0ak0icWSZmMSNzLHskF/UmAcq+BRTc+gwehjJ8BpJLdL/YNS
IcNENnNmeFIX/qb/XLVxsbrOHYAupdaa+zhNUQpECeooLBP/0wQ42gRp/q9re/pQ
g/e2qaWAHzkYuYVRd1gQqJ5zZTEF3Fa7eoLZBFqiY6dfTK5TPY6W51Cl/JIay269
xHcA+C1q1M7QwHJtPJUPOHcbGqz4AbJvYmFVraXtvtXkWNPXvvurnOf393tAhHHK
EX4BZRU+9XBG7bTDZzuMVxrLmdfrRyCUWfn5KLfe1KZlJWYbjskyHYzH6ug6N81n
aP2oC/qHqPViXcj42TrEMK/zmUwEQ/iFKjJ1/85WjG7a3xDrvHvFGskm/kgu7PBf
3EvlcYBYnZUeb/genSjYwAbqtoP8c12U49aLz3/B2qlvG0Ar7Ze6/iQ4IhEvQ8rP
xGnTwqDBwZX1IE8UB4RyD7mrgFdmL9NUwxdheX06zt19L2csVA4qvBKah+YbSYdM
6KNGayiOf7agYQQ59foJE7YLjIUoKhlfLs3f51uBHHG+G6USs8aTiX7th1iasYd3
ofH6JPovNVlum3oXyy9CG357C8X5ioPb63ChdzSyysp0emZgbZW0a161NotCnWO5
UWYzWy7Kl6koA02LM/TavpzujovKQxG9lwF07YDQzixQCD4lIvg57stRcgMyt5xG
eX++7+RvGb/ttfO1k1ch0qH02RjOCfpC2VYSYxOd/ltINnbrncONhWNbE70Y4dee
iTDQMl53P3hwMhkasgnyfXYeWNCIpF36NJilHpYQEDF7CStzcMyABHueOI7dC7pO
6K5/Sdo3xlEoLt3clz4ynZn7d0tqtKv/OA/47Jl/jFvue8r3y7FWmdnMZTcvTGQV
Ayozht35IqYmMk+5bgrrpgYK2lMuwx3GGQc67fIdYLMDHLPONJn8WYlKI8wGdL/U
g4CcZ9D5aqwIx5/WxG2Y26SHaTefRxaDCYNCOO1y+e/Ti4JsXMOo9hhPYcGbv8aD
f+rcyWKyjKLFOIoCKns2TPK1lmosoZ+A1SWxaqq8fVtVsfYVzl8YglEoxoEwYuBC
Sl9GLmbeCOejEqsSxb/tUtEIl2xu6i1PFDFZ63z/OKXt/v78ouMGiSwHiNMxPG0+
knn5p/FRvIvasquklNt3Js3hnpzYCx6cGuW8WVOq72BJ+0k4sUMea1dAyWVQ3j7Z
J2bULiw5xhetYPIymqQQZ7p7q9rv9fJL/zdra3qpsqja2dqMAxJ3dVULFuabmd6i
icAHX2cjV+cWbgvdjb4PRL1xuA2rPbIcsUmVo1kQvdtCa3kGhMfVuFtLak1XAnsp
P+NesPo6T81Dljt1Cq3B3A==
`protect END_PROTECTED
