`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nBkdZ/nIgK0lFFVUFBXb2gBtMbgedvdxPaULXkAJZTGrMZ6KvN2/khKWVlr9mHcw
oXH6XV0/oceg5lc1NbB++1mqlvnKbjz7cXsdMzhqK4rcc7MoRXRjvoPmoEwhcDpo
sIvNyVJDVXb29Il97aWEcPOUpuBgS9CRPSVvhKpu6lVOd1QGPIlNMAxb+FNdf+lR
EZY5fFqL4qw/dgoD0/yCY8uVuOje35onMp3qhJvSZ1OdRhFUR3AYrn1CnfVKmh0J
xwA8h0yVEvFrGe54a+EGU39+dCI3d897byhBqg41BKxUuRSjV4vLVDwx4+ibHNfR
9QCKOoTZdtlyh2ZJ9rozBXmBohx2QJA/x+lkS1nI0iyR9Y5UY5Azkg035hnRa0P2
B1DL+sa4raim3QVJf3igCLJGD+1Zw49o4gV/yt04ahg=
`protect END_PROTECTED
