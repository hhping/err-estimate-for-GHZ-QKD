`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5y4WVQuN7jo0Cq/4jDwRdfoEtrJbNJVlLircRNplNGK9F4ww97v9KCn+fGVJRTlJ
3IP7ybhmGAwrR4vYYToU1562xoZbRnF3xt92/V0+k5N4aOPYuP2xUH+rhHOrGK4S
r4bpYONYdac+u04gbIAjtCrC91rtrmefvvVa6GZVaI1Rx3rE3HBgB1U+gpA0Lj7b
9b4bUryYOp1IMYnNEehU3iACDhofkxBGmHqZEg7DNtDGTnT2WcVAZk1143aNy9uo
EMi8BQ0ype5hq9jKQT8QWJljqKsP3pqeOBZZQOTwMLLuDW6TqCzpb2hXTVcJvlyC
7KQJgChPJtFUBX3EGdL9ePPV94ypPG9LnuhEA+juu+sn8zk8iukhiVuaeX7i8kaX
bvNgBCw8W96YEqiaxblQFM7cjrHZLPoyAiyxR+s1Iv4kAB+2uLbESLSBSt1fWakt
rxp8XkIpj6crOaGn0OOzd9ASLbKvIyPZO0KIrL81SbvveDgm5X50uPbXZ392htnk
eRHh2c+UHiPfgHqYSDdFVgjARSA1YnXB8IrIOci3nbfTVkKTCSvPEdVx6FuxPt+c
9rUo5mHEbCHZE3Lwkr3FSjTv0oe6HpFUrvc4dYihqcewPMHHBYokwMnGxWkBAf4J
n55hlmDxt3SG8r0uc7I8Cwiz90yQ4w2v9Pml46cP2vUUkbS7g31LayDip9GvvR70
5fWVDnF7/uhhV/QLnWEHkrEA/kUSbPBnqGmqq48n6TKqVddVcZ14LODU/99hkr+M
Vy/h0IQASYh6apTaqvosbHA8E6z7NHxmFbqsixlWtrvxLFsxegYbD9RzbXKxCJ3h
k/W4QEXlrKZO/yTVyF6J1Zf1Ft1r2LGUrO34oP6j8GPtZWGcwGhmqcmDq71OQg/7
lTwx9krREMrojzP7O6Tz8hTTq0vYYwI8XALjM6FigUfc6IJ6gqEM+zQJreULSzVK
320AcItRmAtgx5Li20ZY8OTdN4InwPqPwlgrswWIWAVVT2CxXHov3vmIkzjck3UX
zrtkHlXnvn1XuJQ+sD4mca70k1n+ZS9djXAORyvho27K6lp5opdDDsXJmGSumZkc
F8KOQQKQ8czt8gg99uNrItDuGnjJjvpwrY3Dho6wuR0=
`protect END_PROTECTED
