`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3o4Mf4GGqIX1WWMFTnNUxazmUgdsivuGR/hQ1r9HAx5OXAK5LRXFjZcjfM6mSIfJ
FnXZcO41kxnH9edLFhsR6bZx+6Jy2+yL7h+qsb8X8XZuiOND8w18beKp2DFeVlwK
Pp4dW9lz5KDoZo/nnhijDBx1jB03LaTRqLqMAdw7kvVDkRe28f6RG91aPoE+L2qd
twoAeH71EoVQ0qx21P6bmi8fcUwDyZk3xya7DI35yvFlGrEGIewnXe9qO5hG4uab
loS05Z5SxT7EhR0rz5lMUTm2RoEiTm0zCYaKIb6oPlJqsj6QCGu+UcuELv8yBwqB
T4/RAKoCXxCOqSPdbBGBE5S/YovRy6SS1GzuXq2cBKr9bmmFPCVAoxo+gNrcVL8i
g6y9G5CI795XQbmzd/2SXNGCG7pIpaTqdj34kNspVGq0HF2lkl3TMPZPJjNgdGSr
C9fionjdWyhNR02lxDPEWsw5eLVFHceSnlf6XFHU8uq4t7lDLgTBO5T9xKVC9HmA
feXhvnw/4suGUdObM0CaLCgHW/HpE1SzVIun0g114Iuwahqbr1KRk3fy/Lr14NdQ
uOG3E7CfyyU3n0viNDE0NsKkr2yaw2EBwybtOEpf1n6Qj5bIkun1ChT+FEMIWsM9
jr8bkhRPyzXJYOUlEbWGqDAKjdW/ND86scSf/dxKN41tKbnbWZqwh8J8+DXIyqoS
H5U/1ED6M8pP/0tV5dR+3yHTvW8B2woWmLEEQuToMEPtlutNjdb/J6Dgm+cRPKFk
lsIgoR56qgw1oaLxd9okiK9l5++6g01iIBB5Djb+40Lz9fuh21T4sunZUZHOSXlv
qPQDY/oPanbC4h9rWCa51A7xce6nDUDheFo7CfqsHIhEILSP3sv5nOCXqv3CO/JU
SPmVKwGtXjM9SDk88F9MiSY2YNOfsEzyMXIvc140+EhPTgQjz1ciYvdPXHHdLG+g
uBmNts+ps2RO1Yyd4qwRuX1FeqejhNXobYBDH93JaZStg5Atf6Gr18wbtRN+ThgH
TJdLEp6HC2JHLKbhwe20J9tQRLfUIas6ZSPUgE1jjguifdNVBsOZnv87dnKlyg2+
1bdjayizolvRH0Z+a8m494kM98pWm6/PDV71Exnn9vwqEAOCrUvgoK9f8OPuUwnh
/2I79LL6fHNYSs4b3g/kBV557A7TEOCHfPEfQw+zTyI=
`protect END_PROTECTED
