`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mgPD+4jgZ4a/YKRk0bAr5KomdgGerINNISukd+kSDjFenlO7WhvfWjv6T/IRIpLh
wFOWfUypg1SoreYO5LZ0c/hPIwudljTUQ7zwem7oFWl51GGgAAmeDw4eUBFZggo8
aLFIZz8+7+FshNlKRxYlHaJ9vOt4tGlSRy/b1g2ifNWaCBllWHgw1kpv/K2h6T+G
nU5hCdt/qYRDUNgMLTDli7izYrSWlsKdcCojECTHqkvhbT/x9yGbKNlVRbF0E95o
dt9lrAMsDnv/OylQKiP+slexpZZ0lJWIOP8A1SZibVHZJbCim7vi7dJSXyBy8ydP
tbxt8mrl+obQYdB1oEgaN/IE/BdX7dGDHaOnvS5Bb1Sz6cYWhfWEfHPYMZ+GVQ6I
9CMD34bwcrNz6GH3lZWlokqh3UoCGCaz3sGVF4geRe/p5zPpFroPEhLtZbIS3UK9
ywhjDzkhAE2TesMvTAohU1c0ig6OV2wT9xFROVFKhEXMpcnI564TltkToCl8S990
/aqerDb1syM1/mZT4ZRGxrPJGA/Ls38o0wv/vqzsszcplcr79l2qqyE4Q/FXYCtp
TIeWJSU40NFwQMs1Y5mM8n1M4evm8xbWpm7dARkllxG30F4osV83GrvLXb+YB0Qc
mA7+81TczcPMs+s3BakPBVWvgeuSY9ONesF+PJg6v7YqHoiwQ4WBSkpZgX6xOpXT
16x7XmgLpWE8OtJS4Yc0Eo5rU7GJDs2LuQZ4QdkKR7E0Z9m6rVVrs1E72085qKfz
H34+KjMaKWPVqdQ/lRjWypR2Ogm2worI7CCkKhgaOC4KvqL84CoJK3Nc4Tg/1Mff
rFPwXo/Ucbjt2ooghC+dRqNWwetqFmgmRJG9BI459aglBAEvf8hXUrtLXXZomGJX
D9i94XdQbRuXOzg8PkO8wXxBdOzg7MEfcPmkP5fGwt8eiLI52FdG0GZKhI5gLOGo
AYQltZ9iU+eoJ76MapLCqPZJaFV1HKgI6xIWbZ/wWEORST0r6IsDYAD05zsH2bbk
b1WOkfz0UhQnNDu0VXy+pucWcjTqAbr8MD2o5GeO4rY=
`protect END_PROTECTED
