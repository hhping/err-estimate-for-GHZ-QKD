`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bf7CzWAOnzX0sFCYpRurtRu0eh75rJD5a8ir8ySbbfTdEMFX4bvHi8E51ZZ/lKz1
G3cn+0c7TusxBuZX2bVSB19XgUe6cjrgrPLajeNCB2FLq2/kyGoIgbEA8Z0zUnyI
m139y3IqJg5QO4cfQhQrqrsA6M3ACqeVlWZeD+vUUvYfKw6+FS54CMCuNwncRsDf
vRr6ZYYkgd5Hvq8/SYcKzTmjXT3zZDnUsUCsmVWgDpm9Qvbe/1XhJSIU4vVbPn1p
L/g01CXq2ZeYCC8EZQLYHMNYKLj85p2B4dB5lDepwficBYEVkoSuFrfeVhyJiriP
zXsm92NwXSFDUDQ0JaJA5nYcm6X/GOJajK+HLpH23m0dfIeNx+g7qELvg/41ri1n
FsFx0F106gP6krgw8tpj0ZgJkdQOAtrOHpIa2gmFfmoHHJ9lMtNTNEoA8HwrtE7S
7/SIF58zA+jw8/U2kLc/0I3h9Yf/VOIRiz926A0mH8BIFO7c/aaID5xA0ePuHfzE
9Gz7H4xlIM0E7LPMNp57HI6nc3y09c7PbCVCot6ipn4btsRNz5kfvfS3XYuX7Xgv
IU5kc6F37m7dNhbt8dWacXmwhOSKivyaLw9LAXBwP8Z9+HH08WHPFkEtBV8E3USO
6hzCMWZ6erlw/8Y1e565XJlTTZR4X+jlO8el7dVa7DmVTK1IeZ/MJYGUeM5XOD/6
f5K4YP508cNOBYh9Xj/qN5KpiijsQ/t54FxOMEuJ6vEGOHfnuobgMxzYvTDIz1yl
A7KOHP9ukBve6Un3R+17F1Mm2vP/R19f9aAmZ9YUHFJDL4Ep8SNq3nM5S4SDWVhC
yDkoOvOtS2u7ApXoVCtaVGDN/zZnevo1eHCf5TujM5NBOQSfmjnfAgzMA4T7soYy
zUaLgu8qOpi7gtFmyXsahft8GeJjgqOG8E6GibE2i/OiXgSBfrqHeO5lHZb61KzE
OEva/4TmhxgyOAN93zBL6tGS64IWV5RwZOJb5/zaH5yWmyhD4KW2tjMf/SwawIhm
/f+T5MVciSBUU4Gyg4VfzWL692p9xYvwTRCVD18RC+aRVHYYrwB49w90Ji4qIw9q
qrYtJOOxoWqNhtPCwWP5Vhp0vP9fDAUtV01yRRjFVqVG7N95eBY0chOyK+5rkijh
hASq2+HplidchLMp8vKjqtMpsMT8p3jLha0FSPtNS85MNf5pPN3k4GYAym1pmrbX
nNYHLvGWVEqIzRuOBQg+4ShpjU1IPD1PS7m+ceDYlZiTt6TM4fOYNp55YIXyIqZr
BK4ltIcNZZ+IVbQq/3DB74MjDccpN3Ube3z0x4Ra1dl3Vz3M+rgOkeNlh8LJkZdk
RXH0J7xGEFT/lUN6pdn2eRqJAVquz6kBFNJEQ/2nMExjqMe85xcjXOQFCKUpz+hc
dwEwmMv4KbDThSnE9oxQw5xqfeiDLAaYaYwf4oSKPesp4irlu7FmmSPJwc1Bd95c
vIXxWweIKxlmi6EnnJ4p32x1LQ51LaRXXvNXXDZ8tE5HBE1wE5F26XYKnqJVQFmA
VE4Ttj0pROto8e2YD8rAGQYjwlCu1G54oxEtX9NgZjsFEKTT4IaX8G4H/UiFdu7G
kthOYc/u572GcnHkEaofib2rtmGQvmtqgfO0JwqsP5HCyYgaMRRAqKRjMxtwsGp0
yA67drxmZwM/O1wTOejtJcrw5u2YNmcb1Wt6JYenRE61HF6RDRRwT60LkXNxu5x6
tsdvBnaUXEkX0r1r+M068esVhm7XsCCdR2LgMnu8QpKiV89GDKsMwVwXJh/deWI0
MPGEOUWAGLcWzJNZVS7vU3pIjz/yytSnxn12aLlhn1bdIIzU1Sg5phdKitfQFssj
MPq8H22RliyyZj4WnRFYlGKkv5A8B0aetbH25nXIemC86ZmgjUIg/PVNmh0OGRDa
Y9cEt9pdhkKJyxZlkJpMtQ==
`protect END_PROTECTED
