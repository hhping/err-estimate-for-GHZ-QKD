`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6uVgNc70gq2dVO8TTjyORNyu5tPcxDDwrYIdJuAcirw4OPhxsm6twK+WoYvb5H8G
o6xYAUD+L83aZvdjYFWH+Utgpyn0B5A9PkZIJI30G5Am3eDQu+xBCrdcwFIl/6IB
vjRQmmEyjkQHRCtoReBwzNJ6VN5RqRk5ABlVSpUjPFXIiY46cn/Ljt61kw4ok4zF
8jx0P/8fK1laa02ertMOdSEVrVcAkRyFw5Kyg2qk3ltDiP6EyxLamAkV+C75eWIG
AOEekOFzJbbWWKFu+don9P/JrlatM/xnCyWtSSLMfhXJUZ1NEJjkVJopqFCAYhcy
uN0p4jW+d99xs/EBeWRxPtW9v5ByE00KU4VojeTewLFUlLkV2cRhbW9yRrEYRsoH
`protect END_PROTECTED
