`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nVSPn32KUt/BR70fJ2u211zhx4UDUGJ074W10EXl69TDDeO8tUdDQHPs4bAhapK0
16HhLdviItZjW7Rzb4BNMnraoFNY+B0aWhJXeuWyDSgfpZFDaDJlZO2GGh3KK7Ro
MeT7NKs6lvuZbajIIWAqSnDl/0ks9hl2lPxbXHBoDwGqtPXKiW0eOz+6/N0dGinr
y9pvzoTNVc5Vu+r+53zwFEEO11Q51QCXYzSkghzwFmAhZv8ownCOkDIJGovjRfAT
sP/OcCgJOIjsfWTASgB8wuQ9iR4UPSizBr3reV3dpxf+ZkxrdUDS9glZJ9VoOk7k
zoWuYY+RCbzCLa20c0S+h8pWmt+ULueKu9hVvEOPuQ8Vt5catOyhNkOArMKwKDZe
JTAgjjuTjGRZLSYNR97AGhNYuimLX57zl5ujPrKyirFT7bOkC3U+9lplnEDTGVEY
K3yrE+2u8qKDRMGerewpCDLuBJSz0WMReFaUFSC0fnvOVbVsw5Rjh1KFXVpse7Fn
seGHCTYC94vopEcPBkZTETeZjRuOUwcUmFL9fXe738K3uoKz1i7Gu+WKRORF1TDj
vMIbiQHqnABZTXhWKPeCEN+2+wa9AM4GXGtmY2yiuD62WfX/wql4iIEbXVHNhvLt
GTre6vcDRTy9TGM/ZfD7nuHZq6GU5N4DiiW1MU//hOqV56j4oNgK00PyQBqI7gih
1VYNmfcmTNN/3aUmpEGcD0irR0AD6Ycei/qt/mp90jL3qOveb4LMgTfPTdgzf9uJ
pFTazFZyz3IrVKqQPmxqp6EtsYeLGNaD00P3VTgvcIyx+lj3QbZec2RKM0Mv/uuO
pBCW6740r/kpUZVIE3ZUEzVKVs3TO2EL33ODwGB7PXjKBaaUTPgzqm2CAWfo/1r2
SG+k2NNQIoqcJa8nEuGR/txelGywjgoN3FFi85AmgbSPYul5x2Frq2io6hRI6d2R
hxf9NCju55PgVg2sj8PmO04/CT1+pxqWa651qeacagW+gclZ1+o0UuuMphzCLkmW
eNPcjyZpGMwRK7FmcLTo/R6NNretZfQEXOyoRYL+EABZWV8OumftC+K4f380FuOX
1UPo0lFsgdyMuSJZ2AGl036jmHmYR8U1JqufQ8BIruvw0VNSaZzmJmoDc0PLMrMR
ZbuNg2z+q1xG6DTQy4whG6La4JEyo4ESdbeaFEMIqKyMD1sCuWcOrRZlR1tVHLeU
3jQoz1esK10Nu/BSx+s+9ELqKCk2R+h7WyBb+WBX8hRzxm5PL0RaokFxWDqsOSn2
/SeCYzN6nY7iAzqM70pbBcR4fTqyCJCjquMJLqnxt1wSqtZ3xBCo5HjkWRBaELCo
9auZcDy2bxsWAV99ka44kR2kYyDlrfZRztD4OuXdhdVsgBvT+5x6JHjV08A6Po0V
W/cTwH3QiUknwBDMTVxiAkmCOqw3CjqR5qoBy0/DRtmtCvxb/Wf0Kfdc+XFjam5I
8dzQYTDhT3lRhOonUk5/ydqIxMVymKime1wrPCI+AyzZ5JUCsnIhZ4fZ18/cvGea
zv86C/8yhS6PfwNBOklyE1yV1L6eFPOKs+lDAad39bw=
`protect END_PROTECTED
