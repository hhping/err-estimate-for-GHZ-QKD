`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iYQruI7uh+CtSSN/eHVnDpNQRos0NZT9IKBtVL1DgXzAzoNa1QNsr4hUqmIsFhsm
gu3Ga5HCbSbVfBFNWUtmTdtHK16qbZkwNG2XLv009CY/zdcbJ/lJJyMYKdLLskCP
/Wyzi0lPeQSyy6ARA1VAQ8LI0UjWLCv6XYPWcyUxHHKDHfBWKEdFTAIRG809VsQ/
puNuKgtvVwBqeGGIiCCtgIGVJC/zDOsimQfFMLYAWFgHkcqtQN9AoTeXPw0FCSQ+
BpNaoyBSc/GT9030AdjFXKl84BubIzQ/3GElTAmzAC+piCchGPiToDvGPUfpZQ3O
OZMbMrRUINjNGKtuYs5kpGlebi0XKLX2u7zd+RSBFyWz3HX236rYRUe+RYyArx2Y
JmTJjX/KIoY3i55sSyjaaWrjltXLXr00gv8pZTgPc/uVDpv8Y6w6zpAsCc0qOY4N
ZZVlVrrkPVseqzCSVgEmig==
`protect END_PROTECTED
