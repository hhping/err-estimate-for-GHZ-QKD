`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f6h4B7qEhdYa/B6KgP+BP7WiLHdtvBVp4LpVvEeFZDIZ3ciXP7V8ZO22l++/c7fq
oUC3A7EE7f9vEnd255hdiTY/5nkix2J8M95pNz7+tvTavxahhz7ASkNbRK+m9oTU
V9AxIzDyBOx1QP71FjjbxOLbefqayu6lCcONe5b09HWnAD2V2ExXNtFR0nGTRCSb
mTIMPNEG1McYoXxUxvH0xIAqyKSvlf2nlT22LRDLxGvHK4guXSl+2AvZQdsECtxq
bYyLU2QJsHkPLLfAqcTk0gImutbxz834H/kMkXLTn/uOf+TZ4ER2WyZbUq9I1cMp
nYsqKL6MQ6R4FCat5QKMdR+a+Tgk6NGtKvbBHKxV+B7Fd77maZAQld429fFmCDUZ
v4Fy2L4/AmUKxevCdu6eiFmPfy0X759703rNF7egNS5jJxx4RfEk6/qhAL6nKf5D
xWdBjBDGy2C7RBvi/ZUc4rDx4UOfB2JnY+qhhgSqX/JA2UbRAc1fsLhbJFFsoD6/
cP6kXtH4G8oCD0rmjY4xlyOyndUWl3kYXSl56U/F49pLkqHTU8be4Q+r1XUONjJt
M4ucyGi5xdLpEni/M6JYURF7c8cOuCWmt1AaJIQMbRNMnrGU9Vi742yY3ZNwnG8V
y/Nl0pA1Qlln5J/YmcoqYfhDIvEVvb2I7in1ex6/g8tcyC38YLE2KdvJw3G1ff6Z
erEzSCfUGykqbtnxZODNORsjW5AkOWgKNcsNYhYp7zo14kvT6sT5GBN7fStJ9ADD
`protect END_PROTECTED
