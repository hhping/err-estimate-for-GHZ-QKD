`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
es8P861mmGr6bAcAklQJrKIxv1rFNn0ZhisdblpHKvlJbyBfKtm/RR8n0SfbvHUS
sMY64b9w1KzSVy3BGzGT8oHztxEPQ6jqQGq4WJ25IqGLB4iCS+sj0np+UY39WTu1
RoOn/U5qs7J7SgpdLM0yc4aJGywttBndYz3sUbbwnI14QMNfXM2g/xjMko9BQm9b
cdCovesEsPB0wezKQZBkKAv9N0eZgot6bE9gznbsIlZAta56qoHVA6FqdyA/S2Nv
RW+VfnqtB6kqihClxhFMryTeqNImT8JNYGiCu7DOMw1mhZEPsrVJuQnjjehCb4hU
hMJj6scZ8xqJ8zJElcAZM0j8jneiijMIUe19OxyU3TGWMm8WKK7Boj+mMhBGKb7I
4dNzE4+pKZBywurnvGA7FD0aEWFnZZ1YQsWuJnz32Wt1jt2Bz7H1+wqXgCPjj7cK
s269lgzV+I/pUz+gkn07rTUUGpaBOr0vECWB7Lskq6t3DRaHeMXrMLfw8jwBOaKs
TxWD3oq7XI5GaCN1fomgs2LAdP6It0khcTssqbxKEnmZu5yncWC8iHYnw0B2H9e7
76d5j6QiNdDxXDEJV1DIFpsjcoJxLnXygvKZ6FAnNAqJkhKL9vrAvKF21ztl8dAi
kMKyE6Mix0WXG29S5ZybbA==
`protect END_PROTECTED
