`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fpnVzb0lQ91oVrvkXRInCVtF7G9kjdjuahUnbEb0ImRRUzAhhAz6j4VP18R+A6Fb
AaCaNwLhbHco/O2cVixwMOyA3p/nmHWldb78zPTc9JI94e/xIkyIQV+pXs/bBKNM
nzxBoC871Tym64in4VOBbS6LlfgocxGhDUDO4Es8U5gbY3dlTo8HTtqS5LJKVzUn
RQe63zXBUni5eveIL2LveEeEWxuqAADCnCIdVcNrguV/3oHAiEHgy8Ns2epXzSTO
Iu2cxx72nJf5Abz/V4r79KCrg4RO0uDLPa6R2/sLbXP/beMiLaajXf+ZS3Q6Zu7L
DAf0lc5aHtAIeyTVOSsmXpV4DPsdq6qp8JR2BsqCYiq7bZDUBBIe88NTUrv1+dzi
fqJImlU8dVdh/jxeOqrh1wF2kNx+cbV03j+uf4D3jANrcRosZ8DDSJC5kY/lOQog
iuOT+ybvJUaSpfFLBWhrZcBmiSTwigUcC5HS4gdyt5fj7jZGPXtgE/3c42Y34R22
2bMBzXSoPngpiC1KlvL7iMUGrAd+kFMmKrvB24kmnGOC+oycLOSPFuGE9TevJ+K/
Fa5M4YmCUOQuRx1X+9CNmTY2K1hlY9nx4cXNirzACwZOsyyEYihfXF/F4wbrYRkK
ln6vSq3W5MzWc3k1XfvDnMzmMeYK6L+VtkR3dZ9SfBC80kkl8NZBdgpxW4qo1oFl
ai/pQ7RUcxGQKA0wqZvCXMasC2jJCnqI32PTuCfgN08eS1itrGOldbbFFPvNMVBS
kMiTpsJH1maMCMHsPgLpCyfQpTgUUicHyTaXAxf1zLnynPNeK2ttGSgwN/BQqq5v
8fBmPRo+UXVUDbY1luycCbpciSC0ttznPvcFuZaRyVCyF7A5l7tgX2E1v/NIw8HU
X1p6UTBzdR/NGcXZV4WEyG3kecGmat6v70WcZx8u2GWojZ3VFqAsBA+9nS5mfq2b
KORMUK3/3C7DO/Aw8gLWTUJXaK4oVBbWlgbDyD9kNxk7QgF2GcD1mlfq5LPZHVkZ
2Hv0+MR/b8+cFvOQ+q9OKf+GpR9kJ/jjOKhL6/XT723cNuUTrUZu7S3o3dMDw09v
TutSJFquuHK6fPyZEMsoE6ynOvsodvLjhYp9EjU38u3/5YoXhx+Baocu3S2icEKu
+4eD4Q8fPLqha77Fi9N4dvPteQUFqFjmFtLsHAGmDhtT5UfIMwkIGya0L9xGhkXA
nQTP6JyOGWYCweenZOjpASLOhBirNgX/2RxoLnwqAVvssg4mymQP5wcLc5bLRGay
vyLV4Cf4EXYJ3aQXqEZizJRdJwg4JQ8CEQZp/F1GXKVOkNHYLEGqiEkhcJ5AkmiV
hdR38Ik2k9c09703adeXQCjpxDzo+1ijfgSQ0JCBfhyFdqSKS3X+fdVfpSil5V2q
cJuTvtaNnan3h98t3RZiggQ9TRnkrrwb2Tx5vSXlh7Sn3Th6lP1ro1Mgsujoxjf7
AucJC7OFsJwZf6eSNt129e+pVr7TmuaMeiF2KxY8D8stkgZTWzakTUbwOxkGoD2W
7RuHoNhhv648+3Z/KSe6oBEvR4M73vcFSReRT0OJYtyUnrRT5J8fBjvWOwUOdY8d
h1QBF/nN4T3Z52/E2J7B4ACWnEuLaOZRDn5livq7bPRSb9lhdg3+b3NEiRicvdkv
KyTHKqeK8GLIlW9SU72IdlmMptfM6gSekDyhbqr+uIFJPUaADMQT5wvrUqpNiTWa
OqhN84NCJJjlgD4C/wvHtbE6yiQR1neO4B9agupuPV8kAfOXQ28MywMTvUBNxT8Y
6x1FFpef8W51vHiITiNf8R9MsYWD5quVZT3EeMqPQqB+QkmUt4AKHN/uuVhE2MLy
Mtj0LmRV8iTCYIfUstXwhgHsw8mFKl7AvfLkny/T0MochGIfX+vTCRKlXUNB+eP2
BcBZokRI3Sp2CpNUrjvmww==
`protect END_PROTECTED
