`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2HkZCZ9DiTyPo7NmFALk1+NbRbwlaVA9PmlNr2M+Eea/ZjF3J2yG39MUa1gLeN2s
dwxFIOkv93gASfRtTtxxG8mJzwcJBo2+MFeGxM1TKV4oZihu4FzHW3k/fcQ9FX9i
BcPwXPhD36dPVh4EQBZw8wFpVlLWnPHtr1JKfSytyzYSB7slFC+GFSYslVBvwUHB
Qur6ggE7Khx7/6Qp/vT3hXMygVmTQtudiVs/5KH9Swz7vXjdk6myJh1d06i4lTMY
CZebeXa6APd4543TpkoT6TsbuL4h8W9LVMB2wgwZbBygXWJLBre0g7xtmflHzsFT
gF5B04v14IJvCNAFG/v5NBkIRUUzt938AD+mA5fUpc2K5ogfEP2F6drM9LO9S5dz
oaYrDWTVX473QbJqr8L+E52lyCN1+3R9cYHkS+621jvhPjpcNaN3kP4vFCQ+VP32
mjQl3k1feXM0YoedlnN6na2j2wSxm4ImkWRGZrSTdyHpAcWY6Q1GprWgJ2hZfSyi
UWovReuTwK2z1syUz4PQBUPCg6HuaZjGkfhBWMWx7Ad16ZJNo1K1E+M712gVZhPM
Au/j49ioiz9n5t9bjPb/S17P54BRdLPm67U4a6yfRWN9QcdnVMrtGd48WSadE4Kz
xC01f1xezGeZA5Z5WWJRSBXkNpy7kq6WGIDRvyNGWgGxgzz4tALBQpEtYE72+feI
jYGilDKaGGj1ScHMw6fOtwoYo8ri2rw9aONGL/2dBSJfdWKTM90ysuzD8Fk4UHsF
FmSO/IrT//mgIolzUceQgDuku2OHNP4Yr/vi8V5CGYv+JkUNRiPIybWnXFmtie0v
AB36NlJNSTUPHrtCiMxYR4CF5E1F5KbkQTocrgD0ec+5ViypJ+5dPorK1//g9yeI
kBIoaR76tNtWcQhgVTdNUoAZ1AqmwKfXZcM4IwFz1/3kpeYM0DChbb/n51t20mjP
ctTFlbbDgyP0wVVDt9MASjZAvirLQg8ELwbNBkl/41uJORhLHse/iTUJasPda+1J
H1jAEgWPSbFKROzlqnf/VnHaZGCgsInYuEnoqOSxcK2V3jXDhwJxdawPwmEEtNaA
Yy6m2HXLlWALdjM1ob/KWdCzWyU96wcpnf2bkjyw14au9+WoWNqROYV4EmwzStf3
Z0LPby/olL2opvcQR3ITAYTylcHYpHOgV1GMK3VQoDQn3H18m3/4rwXUm5ZaU6oq
KdeFC0trVX1ZB2J7IR+fYbBff9pNCU4N01sKiqgbl+dH9S/2963cMFPA4T6IJy8c
`protect END_PROTECTED
