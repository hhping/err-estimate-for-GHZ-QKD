`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6dhFtkARaeucCFWr3DC+iTn87SClHoxiE4TRXyXUzobp9wwBPAwEgf/n1sjgCG8e
Jx2zi6JttJ8iNo0RzxBrUxN0pJvVKTr39IaYpapY/2ekkQ24BHas/EThu4egSYcZ
U5hnWLTHwYroBm54dFklKb9mdCCL1rlIDxTzK/qdjmItaV3bXxiPUfPIMZ/unmWg
fZqX4IN7KwrCSfvPUShB8JK2M9EMMfjY8COKjfNM5OWWSnlgAleA9w4U03nkicXe
w9vkKH9aIvlYbNazlQrmKB0tHtMJBmUfFfYw419V8FknGLNWLIdyXA4XidQmGNJ+
j6NDzDeF6WWN2+Ra79YnbdNAAVuUwx+FO2xLjzyKvhTR2DLCXe4A6naPpgJU2zm/
X8TzQrppMiJ8YlYVUklI1l0RfpG3TVHkVmbR3WSDfQJ30OZJSU7uQcxK4e0bz3sT
4PqKfwM41UNxJYyAwKC0fOhEqk7al4EZcQQtj1qnsfAfC/NV/2lDfvbeeNS/T6NI
7FsOghYZd6+w9WoRE/s21Ws1URkHdKy2ZY39A4ASthVgJUjTXO1hFb+etlwoQfy3
4K19pNuOdejnNklzXCXJwVDLbGfT0xCmxt3qzHZwRwBUd9PvraSFO2CFj/672KZ2
ob0qGReIpK/PjuwZ71ddijpbsOFfQqDElSLnqAlRqdPL9Bp1kDWVH9kwyHMiMFOY
ROV/5Yo7lDytwvor02q2WnypQLx+McrH+5k7dnjn2Oew6iDGWrg7TyRcKpmu0mBM
SkDzW6EszUIC/2nMMPbgxjo2gZfBSU9L17Q2MFqCGFXt/KPz9xTipM3jngGffdwQ
FXMtxFSJ79wsoOAT5Ov41SSpYzfC3njAI3KTWGK/A5S1wdTFIxXLW3m3Im3WnC9A
nZ3KOiIEBwe9J3/RAURuWAApPniJ/6hednl3MNm7J9mWqVD6kqDMWaTIIDqD1pXv
SzUY7395VzI9gVpemTybjtA5rf5CtBRVNexifWHVQz08PmMFPyp9mgx8QlKtAjEz
BkksySXvt363S+shfKqku8QA9m5v1ACbE04D5Xf180JHbf7tGr4dUqi12baM9kY2
OyJLnU6NIf+U+gtTHdvmc3BQS4BbUNjCnPnQ7ERW0cPU7LJn4YaiNjOzdAa8A44/
QydmWWRP3xc1hXA/QfQH4RZJRRYV03royWde6DKxOgTMr6eTM8Wo6NGDaRDp1gxs
JFhKMGQOm6IiSWHxHo/NRr72H1gPisd4w8+s+vbx8B8JYZ3z1VtAPM/pRWWK5Q0X
Ln9vjdM4zP1TXJtQIJ2s9h5fzuYx9emIFUvOsql5EhjnrkyH9QYSiYtyWMKn8GEK
st50HPsjXPA1Ig5EnMfubKMSgET/kjSbOCSnBbVn2zgm73P7aqswQ5hgT2x72Za9
sojczH9GHLd+ehp6F6vu+rNhzMI4q7p7x8pI0QLfbEEvNPrhEpHETTWdn78u9CcE
8H+Ic3bKq7MZYIMMuE7a1Bg5/9cy/r3tjGurJoI+DlqdqxEV+puDi78eWrfBjw2M
hS9P0nsMKTmVRvAoPJvygTBF8pinXP2Y/r4NnuPTUg8TmPhmzrK4lOid2cNLSsWJ
sDQOtjVRcUKKkim2Go/ve5XJSbs9xuGWLeCzysmKXIK47JwaEm0Nvk1JSTUr/id+
ur7X0J0ymrNrLa8N5hsZ72DrnvHYmzvDSyTj7coDBAcRu4bgOVt44FYb8C+X5e9M
Co2vG83+soZoVIM2iifSDU/U3jIV2MTs4QaxpJS5I7MY78kY76MfrDDTqpYcb9Jf
ntKHOpbHEB74rw5cn4ukWmjMj6RX4M92k5143LeZ7Vk+1J5B8mMlXHZr5ZIva3OU
T6LzMDbgsSj/aZijGdz+miaCughTn9J1HUGueZJDd+2qlTDhKmdCm/7C4bGoWMWB
PXHcpyPZ26xOr+QofoX7ORFE1tC6wVSx5QtOcbsbNibKTZ0NKb0pt/jtq9aAd1gD
a6pnDZ5TYV+nNN//TExpFwYtFCEI/kJwCTz3He/NzEJUpeie9b9CVTVWcJes1+w3
9ty1jc4AHJVQWZfH2X6NtOvsEnCpqPfPB+c8h8Br75qQoHMXo3byAuIGv+4GFE+a
TjjbYJMdBQHwKxoMrG1TcbBdb5mgc7Mbu5NVMCbQASIWIB1L8yW8H8QWkiELJ7BH
BLG4K0mCwkqmXvppAIpNDcbbfD6hhadPgU2UZdTD2bnxHGV44k0tpnj3ycqY/05P
cicdFjAfTc7bYjlL1+biib2hWOr8BSyxc/CoGNY0Z91f5nBjCc9Iktp+A+GFZzjv
`protect END_PROTECTED
