`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tsy79cbve9tar2nLN8HwiV8bHqYiUGlzQcacQH6YK1a0ij1iQusqdk/FW7cJVpn1
uFjIzveYjx00/majbRsIORgVkwABD+b3QOUc8n1MBz23EjTuFRgOwwSfwNZcbBAy
HeGVlgBqbL4Hi6AkiG7Ou5XhR1PCKujnSroCVBdx3u0NQUP5wH+eyIelGIa/z2jZ
bcaLfAGy7ppfCzT+mknsdPK8bEA8lzmdJMI6mwRGD7pXtVW1Rdy00VvaalMo0NH1
uiyLOY7JibifdifJtmqcjkJ+v3o1q33qXGxTvDj9xxyCWg9YdvDKZKNl9Ycv5DYN
KYxgtINOSmKAHXMJRkX5q+qEUcV0i9fDpQPT1EyGG5gzeRyn5UVTvEEd8ZLw9cP9
Jfc8eA1muCCbHvlStAm4PbEaUQtaUu3UqngS36krmrg1Wi4jBWjk7gwbOfvnIw61
hT6VS19B6NhXgpepeva8sa5qSPXwB8jedKPhpMOaKf/yjS1fcWLGXZO8gd+UA/h9
Dszm9Ie3JDDTVRgza57H+pljX/iegSrEUALSuEkAp6R5jwbBree81DmjKyX2FtTy
ygCIGP1wGSdOQ9GLQEFuS8TjmZgJ4WjyLAw7h4mB7stC1b1RbPsDtou56suKNcd5
xoQVBmJSbBBGWLtD3QWu63c1zqvIOVhRIQrtkB0MV9Qs7JzzLWsXIr5MWF1Pxjs/
YdZ+B3yw/6ME/TGOy3gV3GX1wDWM2ATJbVcEni/UJ5y1lh2iV/dAm7mgCpgDJI0x
+YknucUqzs8E5swxkwdM9UEluC96x+TMGjS0DJVkomzP4uod3HXkW5YUhStUAJDL
PM2Ja773c3yziVezxVIMIALArFmi7TO2Cf6BOWBh6pTAl2yGk5l3ub7tcvjlsjUD
SBCk/kedtmKBLPAqgaDk+CTgF7PwPZj3h7RzauZBrXxQE+uxIm5vZBDNJKzNVNh0
zeewplSAkdmmN0aZ5Ue7hlH8u4xl8EbPmueBHnscZRz320xGCuvS80WowotwtaGh
D/mf/IuXtk0OPoYPR05/7MpXrQHx32OWpWaF/36fUB2PsVka+4R+GCKYCqR1Ld4F
jA7TTeBSznoTeYvBF3IQuxfAEpEkGruDf/jHhqXkCrISLsgkxA+gk5mJWzSlyHnB
9HaDefuKQP+bfxsPhvDKfKj0wCkt3eBDhT54881Gzn/6j3YdHk6aDloSEOqUfAJt
PvEy+Mxv/QIoY3qBthU22CivhAlDB+L3WxO842ncRDCYMY7Okb3xAqpYGmtNW1w6
PH89mD5waJO/ZTOJ/WORVIP8+hjoTnvfCUWFWV67Xo9hU9NjJaVzL4Rrfabz/ACP
qX2F+gpRDfQj3Ex5g1QeiYgql/QvXIR/RUPEjUy5Qgwru10hftLN6TcAW2KnjyCS
CxUCCkKd9veQSORHfcGQVAheupDZsvL8/LKwLz09vqQE4vJmJ1pAkgOy7YmrDEwx
nc42bz8ZF99XGzSnNtW0qw==
`protect END_PROTECTED
