`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W1UXh+mZLayGZ/50Y9UO6ayCfCk314kYam0EhUosRKexF8VY1tNT2KNnUtwRAvT9
TgZUMkMEskA++3jyRa+70PJmtYY0D/zmgjoxwL5I75fgfWDRpNSQymjsAoAmKgEx
rBomCO0+Ya2biaK3zJpy5MBdGLo06czKeZ/br6KRDQxwTlagnnLcFMv8OVaQbi4g
aYMutolWnc+lQ8JETkEf9HA5iFzk3Zj95lYZ746oepiE7gQPfGAlzl7lj3kS9iug
y8tPJfb1ptKfnwLzXvzgnrcWPRJlsMY+SPrDLjgUyj1nzXJV5tPwxRuaZxLS1zjF
UZMnfPMR5Wg1K+DkeQj6yEGD3e7fPT/w9J+HiyIte0q2LIbnpHZchD0umiI47rrT
19b6HChTmQX3+zuAF7bgBSsQQe+n6RnTbFWWCZq1R3OPSTXXy6lJQ8x8ZFQYn+1c
qmFIXqmOylfzVthYBnXqjzxxy79JkcekcxDQOCPPsptCvfMTKRb3YAd6eoFhBguH
GsuNiv6xacITSSqd1GSuFLHOY6mAfQkX8WDxc9kn1LSLGoaqLV7sjgKdqPs49uJo
8+vv7U4hu6O/IHluCNc4koTAEZm8RdQfXkCZn6/zpjHTHzuqA6Bx+bMXRQ3crFFW
x0admkR7Z/mAA0/e+bg2JwxKVHo76cWvC0m1vSTfgx51SyS9y+poNvjWonCpQYYJ
H1YHoA0XT/HZPHN+aGR+kbosBcT+tjQo7mMr/Yfgmc4k/O30/MrRHCKKdj7gkoEh
ARXzUS/uXi6ABG2BNvixz7ca3UjkQc5hb7U8S+kTP/A3fAMXxyRR90oLs/8w9Xrw
4DdnPzip0Lr9RamZuY9D4daPQ94AvUDI0L4Z7mglKI0cP632FGe5XzXZOjvlhnq3
YQQdaLMbQhMpyy3meLCNbQ9fpC0ohlr63OpAwewSUMRfVl75yrngTrO7fr15Fqcc
`protect END_PROTECTED
