`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w02XP4dGSfhVeg/Gkob+e149snZMptuJT3K1uJetZBo0SabSuHcMgiNhck96O8XU
GKwP4mnNbQOiOlfyFYwmr40YAn1DLaCSq1QPJ/GxWMrBVGbLxUSlGIWslbPcF4f3
CdwFvSElluaFDyLD1HJEm3S/BAPYa/p2F+HlGprwCjhrQ84V6COrLIl3ahnFVEg6
pfsmBqqiLpqogO7BhkF377Zb2gqNlJjWAaUQ+WRYwLJtDzR8D9WoQjkM9tLqMQG7
r4/u4hcPZSV4TiJ0xtRAS8lpQd7oN2Ul7jBpnyfO954XDZZ8kwE4l914W8jiQV9Y
MT9kBsPjUlJbMEWpQ78rP1ITmIkZPNAeOqxfCZ/UfEA1zTU0CkxbG3OQ74wBteMy
ue9mpuo0OpDNPZTB8/SjURx2MwrQWfZJuFkmfCDsny3QsVTgVMeJtkmf/EtoTB5l
a1btRG2G2IP/tTuhx9rKZIJcSQXIPwH6LROnInnFR20pnX7dzV5tiGNqHTPIIa2C
mgSHZ3VKb7Kx7hpCj1W7vexEbLQF5tFAzpHUZpc5wBjS1ebwB13FJAvHR5ChZTuM
dD6AsUB8W86xavSW4eHF1g==
`protect END_PROTECTED
