`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cg0dkju/7hl/Lq7ax0ZNLgrb/IgYMbu4+UUsMjk5NqFSSRvElZ6IlGB7zHGr9RQ6
gnBsmUwcwqe3KG2FhhSHvzEw2qfMI4tov6eyOcvazw1TE1teUx5RyAbkzCuhniRa
5YlOfJo6EGKS6DpUSV19M6d5EAZOeKPnEp9iJSO6JgSalHBA68K8KWDIYuc3BqwG
NWgTLSmma6x608UBDiLXk6IMmuIE9jjmGypBGf6lLeFHWX21jNDMaRuS9dxp+/Bb
03V2vNUuHtCdMtnL3PiuNEx3NzRZ+GuPYaXAIvzH2QJG5A19CkO737X92u8cqWUY
BQU2m0kGcX7CzLjdMzXpI3mkMbsBGaykZLOfHZROAdAGndIgS6mJiNBbvReeyA5S
1Onvq76hN+hcR427iVzw6+gdljK09xTb8foOXOocm7WZKO+IOsdnWAODrnR8JVsD
jlXlP5OLZ3umPD5NX5sXDzgQe32jVRihFt6X6PBaGsauvvUhO4iefhtyyMqfK6t1
MnVILZSbxgG7NNoP1KxMGtFm3IdMnnFC4TF4HZiZz2VIbyQk6jVWdOZRfqpajstQ
HWrw8OrRiuMxL+JVexQnpafi+SolcdSkSFvEz2mco+zFFd0ZiSuFsdmeO/VybCSM
jOFiD6XI9YgIT0QvhTIK2N8b7BhShos3Yh4E0uBHQPQ/vW7ex7Put4hbEDC18r1W
TKC4maJSVsRNUSlbRMG9K1KgvAUxeBgniiqjkwl+LvWpHrY6RGypCtHp2Pdiha43
zfm0oLSlDKO63Myp/8j1HSqfCH8jV99Dcg8CwvtmzRtPM/zYWE+NsmDmy954beNc
1RD/EwZOqKngELvwzuUw3quT30+za9TFHU1hFyRbVGe8wKRzQSeR0AfmQM0hiV5B
6+8hSqOw4XynGb7CT/WY52Wm/wv1cfImnnYEGhxcUcF8UrTyky416pxNJKkang9h
yQukI3Y8Gvt9nh8XSpIo2ye0PO/xmS2VXRoAi2zVtbGZugODE761pGHuD78YAX7R
QzzUFD3OUqSoBp5ZAuF1Una9dB+DUCU3/O53rR4zWIKNv1pRmljClzKHNJKl+QMQ
hqIEjPVadJnfU9IGdshVZanIYJbVm2maVtKmze9wEM71v+lNfsEG9cQ0mLMmNg/T
ttFhe2YoVIfSbGiVbauhkk7URoZreH8dnhvykqpUqShQb2WqEidhWfFwdxgiOCpS
QH7wC5nC4YSEairynbmDixAEMKGUFH7i5ZtugSWEyLvnaN0cY2/QPNh0jsFhylJ7
xBpgsG0+8TBz5bN22KAHBDri6O4eq9SrIoVDGqMRSDHhXaAW5UNNMTiHXX82Y33N
B/4XW7C3dm9ewSESSA6OvpVPZNzIADF6UvHIvW64+oTm94XINsa1qY134TahTVOJ
rnZyWkIgomHFxFl3DLhLg4dnaddAPwz91p59EAFgHDOG/iCPO3neu0F8MeY/Dhg/
XWNdBvSJG7Zm/QSklkDI2vhMKHT3tXeInuArwFPpkXF9w6z65qzmwqrTy6ngi41A
ZMFp78ppJdELjsOEVVg0X3MgmuhsIZgvao+MbCRSetrlj2CKC34SebGonMl9Acmu
YyK6ZbqPZu89M98V6FQx7cl9xvqR1gPbsv/a+JYjsaW6JWCwU08+Tfy9K2P5b34z
ad7f2I+5DfevO6ESJx21qfQxOVKH13q+/R2UfPy03In0TdJtByUugk9OXfMXMOk6
wOWr+ry5D826Q1YniMqB2w4fTJ1EWJg3whlwkeKSm+OwaGvedm5qfifpt/bGI/V2
ske8dfS7OmKotEDDdAad97hGQVgeKs+yVHMDAFOio2olXe60cxXDrP9r4npBp3mJ
r7S+TYw6g4zUzIKjyln6NBxbTXndOEJvipqYG1D1QfzA7SOxxJ/MhsUxaxAL/whQ
ZzTtdWB+rbrMioIYG90v4ROCoIF6M6VMtpbO1ockc/3Y/+LNT4SPFntuotI6nvKN
luJObzVIPeirReELPFSUA8Hr9CTcVqJy4Y7PefhJX9P9egndcz6AWaLsvNc3mAzS
PABRMGW3+OPRNTwTZY5dd/YpoCLTZd6pUhphMsb1xTZ0YjH+5GuR8ZTw6mWc1or/
4uIr2PshRJtmc+5erFIIFL+f8TuKoo1vswGjApQkGcKJlwTyOKzOu+aPSoe0chJf
+XWvCKedzzjCEERUJeic6rTS7t5UJlLcAMyRf/5LcTP90FFRmVEc8ysKYYZ1slNH
t727JxKy8RaDUHT7d+QPlULVVQEycvdlZfD6k+OV5PqOIqdaukbhJJhDktyhcgQH
B40RlqRdtPmadZgwkwG26x+3pmQce3zQdqHFe+WZPmwgb7gU91oSzT81Q7Yf3u2z
g9IaINMgk2ZZ+RZlI+4UVQjxtGJZxDL7zsRne/OTRxyh7xoeot4xLD/7hcGQQEWT
qNdvE7NOZ3XRDj796G9mH/qsdZseIYEDpp5m7RSzQmC1hjlgB2tx6MQge6mtvHwU
y7m+v7gkUoF0LYgfKupwlLr0S6WLiSaOdRG6BHQXhdDg6sESAoA9jxdDYMyGVcG+
GuH9m3pWKK1imFsF6MsmzF0HUkmM9btUvHEs/1yHSZqiIzP/ECXGo5xeC3WC3/hC
TTVx0ElTd69qVuw9Hmmk9lbK1e5IRi74Dv5gMekxx2j/IvWT/P7ONEnHnD2IWExs
luwOfLssQ9sfbmH4vp5XQWfSmxaj3zGm/5D4IKxQjCaLoII2uHDqOit2phZ/S8q3
xeLW3QMesw2d018NQIq91UgAzFRJLrnPoZOtcRtKrsCEg4ldqomRQSvJnW9jPIqX
d9BQ3fMZqf/YZl05H+GXr6FvO7Oo45bzbwHbxbNNvObm2T0RiwexAnfcseIhqUHQ
Bzt/MydfZIFY7vTppwJcgKO5XohfHS9W+t+gg4AHAM8Oh3scYm6mxwME/zDLELRn
VntxMpBkozxaRwxCuOeJBOaW12M+svqBcXPqGFNRXJlAf2fpxlW2Dvah+BIoxEOS
PQkS8OqIiXRQD1a3ZdqGwV5VZTttV76TJQCY+KOJgdU+iEunL6XvxHF80uycZB2k
PnsIdaAmVLj3rDyCwybFGh1IDmcCr7VjD85TCpUFMOsiHIWD6GO70HP+kicsc281
JJbZEl4zeRrZi5tHc2vSwXXuQaEIF8iMQgUd4nnKMA9jPZE9M521MPzAa1ki0g+f
Gfy2GYUhWuIfhT2RtzD+24V7EZ4hJnuUM5On2UxsdkjGfxidYRKxI1dtE2XG+FPW
G2Xi/Yg+Gg+C1R710IC6fDzLHCp4QhsVZ7jhrIVrV0IsyatRBobdtrcev06906hN
vFC5aLPkc4SqW5xHkAdULppSIJW3brmwSRTnpewWogqRaojjpQCdGxhcruP2Npzf
JBZ5ojcN40YH6LTeaFzrSDJYY3VG5qLScZSHoZKwNEcmwhH2+zmky+yW8ISLyVJk
af/18SlTMM2QWOGjJb1m5vJIHva50t1UQ4DvxFmMz3FVf3Ew3KEBnqAf85ji7vED
0xSGcu4K0hKEuzEsPScRakbopGhq5FC7XEbeoOX2C8pTm/WiETGzN5Zrc+kSzOTg
/lt7/z+3QqBLZPWsuX6IHv6VG2aaegqv71foCqWwB3OHnnwL7/wXuBuuiBPXwlt+
HuDv5Yh3g2yDJLD9KvUu9aLKETDL85YkgpYFfaoY3JLaf6p66nU457UGutI0AI8L
DQRWUiUtCWpY/k0XzC6s/i61zxN2OQUIf04Sjnt/SOoOjeBqLZH5x+7GLyuavABN
sw7DNd3qRabA2Y2yQxDeb9aD6Kp2t+Urc9arDgZ/PtwCXN3IMcW9dM2FhwBuVtfH
nWZCChPJ6QoKmWWkO1H62AOzU8EZDtFJRcUxB8FNdzJiaEvQVSQvcIV/FOv9Y4Z9
jZ11fabUIoGP0xHdjSvgkaDV4EIVR+S7ILWdxrggBWztpzbqnnb26bAY9FRihB9K
63BfdccL6n6mIe9S3Wo5dfiZfe9TwkNEmd+YoCpDpDVBByOpSDSthL8x/SAyKsIf
JDKztzIgmRqVgVMjVvDsYZLL4aZQIVp8NLsOg+8LAFu4qWPSGDS7hpjI2qJa+R3S
dfaZFk6ZMbeAmvXkHcBnVTMo0t2WjleTZIqJ6gM7a2DaSErwSa/snn+I2mV6gTbs
cikJffSfK7inGbPpgyXivOeYGNZDHZgVnOAO/VJJaGOEDNvz3BrGRN/mRXg/8R9p
KoPGEQhw7t2dEbtf+F6hkbuMpqFXnPpW2jmFytEeO7IV/dwTm5LDPSH+DeUj+8t9
vMWhKosuaP/ZAvTHdOgMmY+qDmKSRpKOGaYslfxLAaiF98Ir7dtvQ84QmteeLvNB
x98/JW0/M+g99rxb4IJWrKgUo2S0UFlAqlaQjGc1Kewzha+C/BLkrT6IstXMyE1W
6msUqruWGBwdwW61IHgk62C34R01MhTWLqRYYPERpisgMRbVjzmGUn3RLSlgwkcJ
ejULdPkmBOy908ohVgsFO8066WKX5kbxqEito/I6nRCgqNA+Dtr4a39nLA9//Nbc
O+Q23OLq9FplBGnMYoar9V2eaSgAPLTydygvLy74Y90E9bw+pm5/M73f5JhQiVyK
hnyRCTDE6qC5rmQfCJdtBZsMI56pU4La5P9qMWDaSzU166maat7L0HVsACiKwKq4
GV9i9WKY1sf0OBhGObq6MbAMliZwIsNN9R8dFrWc5gbFhJlnw9SepltKAkqljH7u
hBIvmrZznG5ewFxhg5yBHNGQeN8zNXPdAWkYxkkkWiaZ4IdkNGWQlUxs+z/1SObB
pEfXLasr4yVnLvW7DFCMOy9Yt0BOmf4dWRHujBoWjMGSB6Ke8RY6tXzm+qONzAHJ
if2MG7kdrWMr6nZsX1bFw+3SglZ8P7n00+SOC6sC7GUo4SfRriszisgMiqwgTPg5
81C3GSTTmlSQwx2al9Lb/NFA7VonOhHndiSl0KjOgth9DhRb0oHnhPxCDke4mXbC
89dQ6+pJTBQH/UiDbII8xS3n+DXFdQIDzFRYpk6/DHgjb8TaR9GrYAfLobyOBTxr
vKWWTcDQkjxHuKTvmknEbiVNok1Htwr0v2G6hVlgDxFJ3uf0m3ipgRB4fP/6W0IL
YIzxRRpagDCUPC1jZBPA9kvxufON77PGZvCgybuqOj589IQNBWDMMh6BcIkBzrQ1
PJLqYp45+p6AetNAFKnc89lOQshGUd/EUSP7KX9ojfGxFJjGnHqt0sFAtE61AQll
La+WHVcaKt2UyTXimcxsgU+SnB+X/DVBlCfBSKmDxzH7RlCfMktLIOl/hULyJ8s5
OaCGQxNYNavHI+uSxnX04Yi83covNPTPmAv5MH6YRD5nD+aHSL+NFjqC3RUy+t/o
oPp/HtTs9CgqdXxLV+7n9K+MXf3GrpDieseO/9PvnUxM/iuOcdof/IKDo1mqQlnB
GF/52ZxselWTGrfEBtu8lgT/TaOTvb+ENymDa553+MGLXJ8zlOPsaLAvrucg4FXp
vJ3C3lxJ8XXAF3Uc7nkVssrgBOENIVxW04dyeqcseBGHXPrabXv8u41I6voWTeDq
n6GDp7PeG++7tqwjeU1s4xgIlOGucTojf2iO0heWbPpiMeMCa7s8NWWwgh/4dvQv
DvpagNpsj8O02AHVgZYwExhh2V21n66+Yvt2lhDUmCfCJdDtAc7+sgu5MC0ir2Oe
55s4URYEY/M3BmdfriMvlllCdrOQlcJEwEIAtZ6bkHs3UL/LHuPxjC9io2N3Wu7v
Ekc2ssHChRe9CEpy/gZ92g1swREb4wwLwlnDe9xumg0/gbFzRd15z/xVc5jV9NRj
gGBhOyYAkLwtboPGhWTOJsKeVKIOpvZFZqxDvsep1RJm4WQwsGFkk54qRF4PnyAy
CMp9msmplO0frlsIQkNjzqsXCW8FEOWkuCGpFiX9g9ncG78srT5NFArNA7Gxvc8V
8i231bYRpU3+Y6nw3jxUmCw6TZm8Rx/j8U1J8ZfWqD/14m6pISfQqwUAR3M3so0T
F6Vs+q5RE5xq/rB5s0C1bupSrrQeZlYfeqGCqKZJ+QpM65B2ZRhpdgvZMrBJk6Fs
0HDPS8qbbkuY4nANz8m+cxHYwC6sJIT+yh2k8E8xA4dii7sf/BJAcvefN4rtciEw
uqS573heYoyUfNZbJz8bSPMrLqUV6zq4r0Th4lYHVOQpn5DdqD52+cjb52eHvGo2
Aoa7QCpPcXclYobyrzp+ZZOD77pWodahQL6mT3+vt34vm1+L+N832WxHG1E469Re
rzgchTOrZWsOlXgelhiuBgw6iR9O/GcK3IiMIzCmNMrNhIzzFr8yZS44E3JuoeqX
+6x8Nqe2BBEiZC4TtMEUB+/r9XAxGq0vpc3jbzT86c9dXLO1148MTfE7XWw7cOgU
J1pNw2AWYBWCJxWr6rrbCj6qpjdbsmLOMNelRcWF3Hha8sqt0H3I9vlxOiZJm/Au
lve4A5O7enzJNi25SAdAM2agMxjSNNispSlNhjA5T8I7rpKT4jUXpGOB3APaeOuV
sF6k+fZeg5fG/NIfNGVBNYmnW3gZfxyG9zumWKqu7tas0dv8SuR13yBPTKhv3/YN
DNHip2V1Uge/eVeEV2Tp+CbHNqSv6XMmL4fRWWl5ThsZRJ00A3Gy5TSamVZ6s71X
rowHGGFbUBbFTEGRQeMPIlOND5nkSDcTTP0Btmi15yVjbZdouMHPPvlz6znJsxfi
8waz7VAaWSNk5a2Pt9astzKRhtkM6VYwUo8q11XIpEFps+/z1xFwe743W6RQWWMT
fTBbOJaBh5Pej+aDE6WUaYpO+/RjsCmiw+OHiT1neBrB4kS9x7/6xxFhheRcgFNf
lSKD+A/JM7AfiSRs/yxKEbMP1QG0/GVUxExvJY3JWmIjaLfa81NlmCVIkgA/XtIn
AtwI1bwBEJKmQ5kPaQoBnHQTExKyhYwnvQ8WEIaT2l4oJCiyfFLfmvipA28T5U3w
HVTtgTu0xmuz2wOM5ZoOdKV8SL/m3M2EVoAjaD0RPor2DdSP55m6lxYV69HOIX0Y
iR6aUu3Emy7kz9liCbCHvKG5u8W/KnynxK9g5mfCU3Vprp5kRRz/LjtzG35X/EuH
PeeiHiYs/zrav2FbhT839o42dZyelWjZQay+8s1+WsS40+9hKc3OL79dj6cMBm7K
Qprg/u7LNT4tyvhGAkq6EdZzD2vKk19RDZmMX1rAKZOO2c7i97Mxz+4gp6Hko3Ox
9x65jLjlzMbvgVQNnhD/FWy4BoELkP6Lo8qvudRggbLNVXat9QAMhFwfzKnPT62B
loR2miY4K5uo6PbGqiezpxJ2nljY31nP2Pe240dUEQT7fIXhmeDjZtDxr+GFVkp6
kwWOsRGOjrK0/I9g0cbpFqFCGfvvAKoiR5shMhNZ40zy3ae4FvLofjhUphG99mr6
6WAH3NQHOiEU+iTjb2h/3Gx7XwDF2Q7HOG65gxqLFLvkZ1e2WOcdD5ZE37xo/QKl
X3VqiOk34VVraQvG2omO+Z/WwlLs+n7dN024TaejDygJzLcU3I5o4uiflfpLCm6z
q3JchjTJyF6pCJfhGdvwB+zlB2JxE+AHrtngMrbF3M0mYIvnKBGc9OPZ2I9eP/mE
bp+3Z+m2aU1DXCp12VkgfXC9Qiirng3hVg3Dkn/XqjEJapWXPW/7V3lO6ANgKEfs
uN9vNgOD2BNI3jKHz9ypMNUh9/z2zGl/DM36jyYLt6rmbfrkZdYKdSmmETdzmNiT
an/c66n6SVQZM97+sR9ZYixvCzpeslLTGyQm+93DZVLMfdAjwCbAtvNTqhleqvZz
upI/TLi+mbM5bEcC4TW+HnRE1+wHvim6guKagGDZFAJMb2yh+j5Ut+vsKIOsocYu
E1IWU77yJqvSDNx1wMWIGQXYJ/B+XoCChsc34Er+laW2lEDq139rZi6LPvYow0IP
Bh7N2XLCjNfiADZxcuKN1WK1JqpNd2hwJKwnSRk4eo6XsqWrui1DVT8jgmSXd3Lo
Abi1Te88hOWzk8SjiZcS+bv+uuOUN1mNPXf7P5XgiQ9/kvwZ+Ah9lE/+KNEtwOTb
BltxrRYBpqxKQcLiJzA01F0Y57H9+9vQUsHMS435J/Xg3GrdzN2s934mNjNS8NaJ
2k6sRLTKpBjujzp8P+PNam7JPLDQP071ihA/QTtL6gGEblLNmTeQoIcHRrdNeL6Y
WKPJw6Sa9NDJFtauFXdDlT3rKV++eEkBJU/4T2B+3ClTJLtvAsSqB8eEY1Lto91X
8qeR2PxZWRH9lHtzvUYvAlpUJIyhDMxU4gEN3kilmfJcYMAeb6pNfpxYxVjZn++s
wBd62QUX6Bhvyuum9Gh+S8ijBe2wiT3gzCDsxieFxv/6cCi+3/dVHCvPQfbuGvNB
VgsqAUpYplqnz7KDnwE63ovzIWw0Gd7piXovIUuhNB+6fpRvET4NWKZh1jVJ9Hka
pdsLvgi0QqwJa7i4Zjz6JygmVItD1OsOITKRMAwlr60SbuA6lVLB4UqpBQj/XmdV
MaGFqiNab3M2mEzeZLLiPV3y3sTwscvI2D1nt2R9kDC+4fsImeCeb14FK/w0D0NP
7s9Vx5EjKzyqYoc8w+Jbgv4wtilHspuecXV/1l9OKkCfyR3Mw8+w6lnl5FGx8MCX
Ai2gPvaMlE0S54GeDrbx0vsSQ1VTntO0ru489+Eu7MXHczALC76SfKgTow+0UdiX
EorabXuBefJ1Si9jfl6UcIZcg0PGvTOphB4RKWJKwFMImzEPy+RkKsEtCeBJvabR
w0L+QmCIlBR0yfIMP2NPgLWZwaC++ijK5p27Kkh+idWuKUaG5iRoq9O8nhoWQoue
GB701eZ00EuL9jeciQGIVzqAp4agFSSKqt90eTkEv3Sd1IWU/FEOj1ifmXN47nI6
BI8SMfp4mftRf6UMJoiVbi36iykT4SbJrDjuagvGF/qfZnhbmte+rsUrBl0SCeBL
GEHqy/4popPRMC/u5Ie9wERE6rUGiWuv1goEt/weGcA3b5X9OhShLN6NAmgNR9LA
RbBbPw7LJ7DfZLKM/IZ5ROiLU/wzjS5mlOHUqn1vrQWRVnymtnZ96YCkwoBxLIc8
lRz0NyA7rkHR6fahUmjluPgsVgTbr5K3JuQu2gBxVm3cjHm2qZn8lqX986KaX+Rj
9Y7dXoczbc83RPMsLQjvgUsBlYy3G6OlpVYKjdWHUufqlqdwVj5vPe0BbTjsLlGn
jv2QOSVYOXjsj+bjQS6VVQVx0x9npfZQZkab9ixFA6Sga59TZ6VaMfXhdxJjIj3b
cyUhZ42SRhq0sS8T8beJ9VChcqSQ3EhbiqkJTGFdowIC4GrDgL+2SYSR6MPn9g/f
3yzas78WitlwxczL4RkxmEhcwLtQbuskcA2IxkBX+M3rlXfP9IDrltKudV3nNfKJ
KQMqCBqogWVip2y0pB9D413quurbSNRBq2iGfpkvNaW65hEcRB9/Hu/FLXby1g+E
roiUXRDHsmqbg+1I9kbn0X6cDue0kCi5/UQRMtC65Q2LeLIyhdSpWieeuTPC/wbi
aKlSkRg7woCc8XDJphFplyHjrj74Oz38NskakNdzNLyUfnQ5misptjhwo3DEm60C
0J+AacTS4wbvvdQpbqQcmmXe/fOLpfsu66CnatEaHD+j0FBWsk2maRkzwCSneZxH
+JM7QDPxoQEOSea/kXkS2ZkJnul+bXiPrfafdIADuxbORXzxTG/6ZBQ6O8BoDOQH
ieP6YmdAZ7bPYKg3dfkofWNegP7dvr8nPIkVKsUklbsxIu5vmj6gPFY8LZNG5xH1
SdqxigEpBQncynNXs8dZ40QujJ8DTqhEn/c7gpgX6YzqzS87+yaxHY7MN6741aIp
gArJzsAUxwFEHJ1jx/A0FOZwxK3ryCp5Xst7Abm3uYh5yU+U3jvD9MUdouYOBSqr
ghZwPmTphK2W00qZHlnGNAD7XwQdQhnyEY0zyez6Zk5o0kZZ/sZWHYQi5ggWluX7
mtmG0o8OjqZD1tLHRRgoUhc94A6tujyaWPOqyoj1JuhskvrT4+34MHU8HnVKggxm
ZcYIg+/i4iDulCj5Qm4GrSRvSatFQGO+ljaoOo2YiKyEU5T1eVzbeqSTSUheuKzH
EnET4k4O9WKKG2n2EumXByt8EJCJb8Bht+ehgeyCp0p5pMIt/yjZCozkEp+3gLzj
ESdNpkattMv1CgSkiABUrQd/UmoucJA8Uo5AA614IIgEBVQZjT17OH3RmH2GMEiE
OCn61f8jQEC/BaaJzKk35D67pdbg1lXs/YqjXyc+hbGJZoBglLyYguaPS+QW+sz5
Rk48GetsLl/1OYruPCLB3ytgcrbiZfmRviEO9bsAKHQcZzHHlyFkXFIuqGNnzZgJ
PfH/fBM2GQp3aoT2g2DnsIa3a9aAixn4C5cAKbOyXaGoLbazWlAnEwsex5OhkqhZ
UVX6gYodlW+n1qoc+qmsK6rdYCwtPNl1C7lKjAbvtNO3HKLo23t4M5X2nAf05ew3
USU/l2ukrywkoo/2EpZh0/rFctlhHsOyLXoxxM2hgr9Qn2MJG6MPBUxAYVjiBKpw
y6/URQey0/hyXEkev8n+bbKGdar0rJECkvx+NsfLzxvgVOAMxYOZlvQpZzWUzNeb
QqvRua46OdboxJjmpQLZplYKpElT7csG4hMn+Jto+YW2O3kcqOHtpGLGPideNVnN
5DS5miA8tB0St8DlWkDcneGbCgfPqxpcQLvlHeL1D/vUuoDS+4uzcunKrcUYdZhQ
nzWb774W8JFC9JHuVZRSdNfqa9VI012Og0POFZ83lC99M22SrwHWyXpPWdw5lMsH
Of/V/jSPgapwmSgWBiW6HUrDa07UKtH7PjuwltWh/6qqbsbufpsKUH1qPiUEOXaN
GsTFw47IoXzZc+RkHL+QJiWZZpKUlSFOdxwB/zL3ZwaqlJRPEQWbEQDcdRIRWfkZ
VGnaafP2YH6HsDh4JvQ4EDNQ6xyh/oYlqM+Z+L31hiuoUihDW2fEW+dgj31V4dyh
bNp0vNrzaW0f7alAayfbpgp/nYyEOjY3cm41kwRoMJ9zfk+EZ4IZ0zqa9dUsoTpc
hEVJH5keGxtvatLCkQZoGhcG1fZXqd9SBXOCLRwoyNf+Xz1M99nsmyPd/NtOImJ4
bhfXhesy9i/bjcGZylMxnY4ewy4CF1k0WIywPPN2kRT6zThHt8x/XjMozlPpalu9
x6SQjGIznYIIknxEVaNMgwaEPz6UzPyT2XmJLxj58mbCgMoor7eCVFT4df0jMYh6
C8r06w8dNp4vgSkkSdJgUaesuvrSYxB3vGCV1+URgoWhA5fe1xIzavoVlkvDECQ/
wOD0jDy5YgSJRXPonu5HDh2V3e5KX15/Yuq1geLxgDxunf95Ry2DMkpPg8P8jCha
4xS0REtbXeu6nY9/2lXQiIpQfejUfpwN52BxdlqtnNE9z7enDiNYanGzGtHhxfSy
+gDUlsJv8Av3eoWkdOJbJflZH4TsKaOLUlbYtCKRrtYTktAeE8XTBwqup11yrR3E
Uus+6MpdL2Rvt9GlejUMWwsbx2s2ZZ9NC4zOYEXRBVpQc927qUYLVAhs2LxDSLQk
RVceTNTq3bjcUsuUpRinKeH5OLLY2qB1Iwsi11q57IARAWxonYgRRPCs6YIVq0i+
ra/Sgzk3g3powd1NRGMMtWR7Xtwj2j6xwnAIa6W4Bn01I1ZGSXWhTxU3h8SHY9Cy
DlGKT9TRCa+IoAT9pxwZZscf4vMskIGdUcrAoSjJCYLAajqsack03m3EacCCPPbD
+rMLkmVD72SU94qsuH3R7RLeq32Aq8hANMtcnwPWMR16kLJHEYOWtXALpwA1HH0l
udtNsaKj4i1o9i2Ar27ADME7U1KCCHaBKk2d1xNCNpHZY/rcq09d55Cu0aLo7Xq7
xZFaz2NbgXMC0EKFp+q849jp/Ohx9raGtoLLX8608VgOTgEB/mHHbrztop1T+RHm
WMYo43vAdn1ca6w6td77yD7UfyRfiTAlA/bWXxm8EZF2o69LU4MMtOAX21GXJY47
RGFFJ0BAsj1mWeMVQTVGONcJSoQ6+eqV//K4ytuEvQrceBoWTmgxR+Ir0B433n+M
HDawxy12rEuvtKfDEVVNP2kb8Sp+H5i7xkaDLDiR4dJIPLFY+/9v3/MTL1SBmqSi
PLSPYqHaHCx59aBMfQ97citg9usNRk22v1qxdVf4NU+53fee/yjObBXEliYX8Aeg
grj5yQl/H4bsBtDpicVNGflUxLZATyh9YsAhixilMG6Q1H3llHJCMpTy9RfZrKtc
atM/8FAvp3cxcVGVvmOiiHPPOIMmi/diUIu8uyBartcw5Y9lkIlaIyfRCmyfPnM6
dQK+39785yK447Q+yvpYt46NE+bfAaP4iRWX3Ln61UgcCpWEtAAMkH0ZJSNzCCFd
bssAo9CxQW5hHJ5S2L5N97KZwpYT9IMdGvqg2LEtQXWaMtwMpPqm53RtdBb9W2+n
33ur+OLn0tUJePcsTmmw+f7vyzy/HOsrP6BGfxZb9FQcLEDKeYgkhyP4Klw7VlAz
zUznX58a8M02geOtJP0I0J+78Bu0ceo0BP+4BGpLEryWRzPOgwi/4sr5E3zlde/s
OfVouzc2Pee77jyY6K0XzrLlC+OS9jkr2OQjtmd7OwrcPj/El/R2Ed262/LoSFhb
dCgOqPuRh6aBPOfzFBHcD8APlSYWAhxBawRycNRoCp+upPsK23j/3hgj+s+UG9Nq
qMIeyhPV0ofZ31ltyT03Dx8IrXnbfoKypy1rKkYzhexv6oRG8YvwvbuLthMLfual
AnTy0iqEv39wTpkznldNXj21hDL6kotQAT64NIhXZ9K6/iXS/JndSl3VeKTjDYXv
/f/msstop1nyRtYxjHcPARz8zeVtVlT1yKxwV27h4zgW/eip+p4eSeOd7AKWmumR
FCW3eGNKvrjlP3jOT/V6wPIC2lfAiQk2SUFDEwBKDTsO6R0bkeF8LY5eUrSwiEMG
d04dZKUQDSS0n84xeSR51qposcEZnJ4C1BoA7Q23VXT/4XJ25fDYlsZW8PjnNJjV
DSgsSnn6ptJmE0cKvc6MWBmJm7nzqG7wc8e7dqo9vsnnsmPokT59QhQWXue9CX0P
vid1C2jcuVLBc8gWAKMhbCLWyscwYbcNPewKCnN8cXQLisKIZ3CdoUhtHfQD0uGy
eo1m7rB62YGe/FkBUgjLQg/HpMV8OcoFHH5XQ1WUVDJNsb7ePfqF/gVd4Xl4ZB8D
yMVqM8LCxmRO+oIKZzTRQZ6sqENwCflmZgRprvMbCJLC8LQkIJap1c3DeMnABtUT
TBsRr2uPxmnY6n1Z7GyZM64NZvojtjcX6NChkP5vajJ+bgTGpoPH2UusldjqJI++
qa2SilU0QJpVMl+s0Yti6z7JtVtAq7BLqOClRKk1IifIL+8ghX1axax1KwcYXtX2
jXr9zdQSMNBCRg0jc3iNKGxuM6b2gyfABu58XJU3fvRytJMPqfa0CpCpgw4nrPQ8
c5LDrnQcKPr6kkCku++1EePnXs8LUUFuTG/J61VmRsuO+tBDM4o9tBB7Ck8Sg43N
8z2YJb2rDKdddyqrXy7/Mvl5rO/6H65qpiiZvG2bff5BuNChviTexj9R/a5OU/+U
Fcip+oR3ybZ9JZWp2wdqfKB1xq2PkG4RmQdqNe0TEu46k9f9RjnPn687pRkUBa4e
6o4H0Xi6iLONREOjtEDWbZqI7XQMBunWaBD33CiayydtrTTlnFj2NfQcbS2/JQZR
fWeXx+y+e1eBQDdqeu9K0D8nz0XaNaQS/SDf2ujb5jaj51gOVg38oQt7epxkRcfP
c9qDDPEZmFJB7d5hICVDLxulXzkebr9bDN/wHrXPmYSgMTE4pVl6RjRwjVjWk7dC
MDgkaNr6hgHqgiG9a+ZAQ+BSIBiABTD6y/wvMOPwbjWKGLlviE25HvSxnY9v3a6a
vXPs25fBZxTqdHkFCht/ZlWbrU57f9eqXq3RjR4JH8gYlALxqlGdo3zjSvZBnEtb
fDUTq6Vez4JnU0DIoFWDRPJxfHzVnCMYjD/R0zrmuQ9X8fjVJRTdpiqrPJVjCE46
1kHA5Og51kKtVEyNrBOgSK7wetYYbYa7BTRCzfDQrHmWB+d+Mc0cdG5kVo3NUGro
p2TwpfGQ/ebWE/UIdTe8GSfpBNYN0TsKd59fMI+8irR/7SzC4XAbuMl8Ex3TA9w8
YJY5ne3utgT3bsf8LpZsu8irCqRkOCdeNcWrdTCQXFELgAHwE0k38bEGF7yNT58/
WvctyXR/Dskon9Y4qV5azkPjMjdqbLhVgMkJCIUNTPMv94zABb1wZz+1vLcUn/sS
0fJBfx+3ouAHRE9be8w0vUMp7MDD26k2c4TvDtGnmL67hPt3cf0PZd7xTheGmxq0
oAIxmK2MJ84dfm7gmYzSdf1H8Qtha3FMCSKWyhP29WZnz81ttk5Y8eJsMKoTUbl4
MNf/CCGptL5cCszaf6UKC4oLQJoG+1ZoV7f0BYwVSkceYO9Zn7kpymjRssOGFmBi
BPG31AkuYi+btaRKv4Z9rCO23mwrXkPB70hj7nQCq9mJhrDqVtWQlmC/RTByznjn
VyRyOl+EWI6s4teV730EJu8f1vhTvR7rEWkhhsMzDZdbCfULbHFEExgvYFfLp1/e
7roSgQ86fLLJZkWwcEnZQnpHE/duqzpHpAW6XmknxtFZRRTbUBm2d2dVz1VpYT8E
C4lljhLyIy+sNE+fDXqHBv1YFpzEQ9pLyjsbZmaWF2var91c61MNvTFRxLFmhLCJ
C+bk0bsY9qW323OCTd1iLA+zW0sIT3CeTT4hixN663qA4VEKdjVIkRhAQXRTK683
9MvwCx2MHfIO2Qp6PIijqLfbtdfDlRe2Tma1UDCQW6O26CwnvK+uDM00k97EatVu
WoC4HbA+ZIMYuXXnfUvc2VcVEewAOHhi3buGaL2a7u1w/XSoV+uEBn8f2Ro/3OIm
3q4QF+7V7IRRYsvq5k9clgzqQidLrbjG/orye/5pz2gyp+5msbtgmgxkdfyF4LtT
gXMxkQ9R877DdV0cCvOcDUjkw/1+S3AqegsRXK42WHpFdu99urW8t20eaLwLn0SB
BxFrgqr+OHUb5XgjbYoxxyNkMGdsFsksPJ82E42fUiMy+SlKE9uuqn6bwopYAwkJ
sF7A5MWYGgIo+ZI4z0A3bnG3ksyTxwyqRVuXpOKkcIyxAl/e1NRzSoBwPM1gG1Ml
D8xdqEYuUExkEYiJOuzCwJDHF8XteCDRx3ANAeHXw74sri/I0+heY3MME/ptePAR
jnuX+ch8VTahurzaEozMuoMVP8oXt6xzhc+KxsGaOUIONkrn9ryXIAH9ZFc4t6sx
iHLNdg9nGUdHdOixJgFzgYCGQ2Xa+dsMGX4mhqIqvz2gJDAjWI1W71AgaQSNK34C
1nseMqfL6gmAGfJMWzXCSVZKkSJij2R2SY8cTxpd/Y77Z2QQ0raOf8rncc+QCU7k
x6uBJYbQrhZzge7tx5ovpOATSXI9sPf2VdjzoPFNw+KFXASAeGU+xfuJSBnWeZzz
Cj0dNFJ29GSMahdxebrLx37NrylCYysWEce25P4p8M5tSVX1i4lpr+cZt48/mNHm
ljgUiVaDBEY7gpMAzi57yfdMOmGt1IxqqzLc9uq/nH94He1Agqqne+N+6iqbUf7u
Di6K45I78QndlPqoonpchLJnho2aGnB8jldHqTHiMLTAllLEt3QLJZhOTXqGZvHv
JkXokKgCGxGmcM0Hy4t5C3p9HI8SsxLj/55xiZs4U0cr2/lXvhaUeVVEpRsb86lY
4DsP9QiKKHMvAOv4vH6PDEBdwRC5WHuEFVHPUBB2RbdsDrW4oLb6Poo2RhEcAMdO
cd4t9uPMDDKX3TXsQnS/NWoQkaykgQOcJabD2O3dNSmr76wfjnjAquTp4jwAgv4I
TSdS4RAP+/OvX5oo/ErTkBqPUC47DeGlPHZ0Am52zamr81rv0wliGHE/qhE3PG22
x0NbXJCDAItD/SRXn9ak6pTNvqBU8Am6NpirNgmQEJtf07dYQuEi1/ZQcLg5T8DX
ojBqrhXKm7YM62nXA/JUhMh2t735qn0Ay3aIf52x+xr9Ok0pahUuOHYUlmLZZWOb
JvLFPtNnTRZVaRlj6awAlNPdiVzjZXf+ZUbJ+q5VJD790NIJIBKpGDpvW4DoAr2+
8zjLpNHai6xnQRmtDVJkTN1F+CYqxDE/g/MrpfGUFV9nL9O8msK4YnsvS2fb15bb
rUwgeO2XOMp6jIb8sCgGOI0L5VRzycu2RvSZnvQnv/jSvYvTrw0acgaYvUWif04q
iBChC2qA0ax0SFGfsKHfisTFhUmGs96hXPPyViJzRB4jXYPIkVH5dn80EQpYZ8f1
HOY8LfFNWcGUvfgTqVPJR/EbqBWvlJ19RCgTX70rZ9YrdnfP3/mM8FWFwCb/WoQO
g86tES7MSX/2+gfGd7DTaauVGB1yA7RXALkEYPQx85+N5GsQ/0WGG1Y+uieTFZbe
djt8SqC0ICJX2JgbwnlzRzHP5g4BiJ0m4ZJ91W9mLgcY+6IKx6wdL3lMobMqkxSC
aRpf+LmirPTtBZn2NESe3Pu40EvMwh9+GfgH6JDZSF9I2cSnPI0fBFhq8+mxqwh3
O6aDn+jcTX3wXtUECeHdoKJSSx9akZbPHsZJvtiZmSMzZ8qLwddSKZswHmE/Enqv
F7AdhiIzFDn6sTtYDAYFiqoxooYZQfYx6URaBA10EuuWNPAc91mVheUlOZGAHsf5
uk26XU/bYYWgpL/lcOs6BDr0pW4Dthen33pmIsjJIlIj555wouWzk9CRsFCsrX4Q
klqnpzpk4YUWErjAtER+XIGU5xvQr0fDnRzEOL5MudWOs07kDASUfnv1Jwj67E6p
qJwea5lgHfpxw3lWkUJ38iEvMecN1BUHqqxtMyBlOGes865RLS5+MNk4EyQsPXhb
lIF3wJhkoBwSp4lMMnYY5aPOExkIpDyjHurp+MCGudEP4eWQ0QmP5eaptOjiHVt0
KIDATzyF2DStZn6D+PSpLbKZJxgjjw7HfN45eZslnm2qKOwJ2lPknk2Jy2+rmUAp
IQeAKKZd+5HIFWzsCU0du587KDVWmn2VWb2+0y/Hxq7t9OnkYqC97mmCkN5ZP954
6aNlAd/tapRR3svVHre05h/BWzlRptu9Kch4M24wGzfQg5kxURBAMoFGnD2q2OL5
CwFnYzBuUU9glnn1V5penmP8yFafCS0Wz2xijIrjlCjmmhgn5EudvHsthAdjJII4
C4arZwqNTDXa7XuM8jRbjQuBOC//o6JjwQdxJOVbsIWyyDt63FLzgZHd7+9V309o
WS6HhoQza1vMaBYMl/WeZtW7DEhyDeHR6sFRLJX1Q6JmHYLTpvK2b/nFQIglfXVl
VrVrGI/YX4pbJsdk7WKlwIVA8JLgxG+slD7ziaz0Rkw/EY1Mx5FjFzBfta3FGqDh
pnEZPpGqi0zjRunAqtJBZz6qhNoQlygkAt+x2qizJUcCiMx7A+asT4y2mLmtMHq/
nGKuXztwoitQWbB91BtjagiRBCFgHi2pvP5aPq7ktbwiiI5NG13SDj34ExDvLhcC
R8zBuf/1VOHyWIRCQc/QZJ7qwTbvDA1f3No41SCkzTgXS/wDB3HgbFN6qzmqae9u
2C3udNBQ6gsPKnL38e1prELISETef3YfIVxiDeXPYrD5vY/sUpjOxTyrFFsabHTO
xmderz6j9G5dZINc/ZKJlmltffebdkuqwq4CV8OCClwA4cdXpxrciCrTJ4WX3Fj1
nljUi9rPlSZx97mTKpNKWtqkvDo1jDZcs6nHdwQ/NGIBJAJ8q3+R82NyZeV02mnE
Ece88oeB1xVbcSXnOje4TFzEtKenmZwDS+jpyinkmx6zUuPBpDrgRaEiC1o22LXN
rfzOR3HgaNYAkSTKAElgHoggoUiQoxHdRlsL6fNg2l6jg7gSAvk7ASlGl+UFmIjh
wMxBHGiVVPAZPUmDx9fl+sinYIfuDhVFqGonpX+qcXoowkRl97AQ7aUGWWYLIV+4
ZQ4XWOxDT4ni7zLKn99a/NERqE3MDUE2HP1lbzRtPRxk+TDKLMdZkhlIFFpmwm+Z
AXBFul+/3d5LQOCo4eggUIofF14jxbKeJ3I5qbmldzG1fAEBtFwL0qm/M5b5zQ0d
otTBKlXjWzLzDBMQXHeZKTEdgOjkhqjwQqhjQKUFBkyKT8FaaxqUOsYWvlHwjdl3
IHFGTpCli3gpPEwTa7wm2SStW1xSnohY+I2FdYY4UrJQVlFP0rScjtKIC8l1jAmr
/4RrgO61CAA+5lHk8PIlhiZ2WtrPZF8bgKa9Y6qhJu/Oe8KyjMXVHyREuFXzARLs
oehT2+qKf+RBvSh8uL1NgefTF5xPYugTeG6jr5AtObIWyYqr8fGGsn5J8JTS9VBg
Pj2zPlXQwXqO1djFFldKL+xTupjotHWUgsBQaDUICTt8EhyG8TEqBWvdilzK494m
z4AUXZuhrnT75jMtv6QdP03ARiQ4Tbuvi0avrlYgflLMFN2hUsmcgvCD2iJgbU4x
9afFhnmC0weGDvjpH+bvIlshIwnUWG24SFY2TspsgnwD2SnxzDGvYRsKNSxOYNWY
Bn+f8Xdap7z2Stra9YNk8nCkfGvj0AoH3j1xgyXzp+EP7X16ZCF8Ve7pAh+CHTBB
oQCtZ3sB4fJ/ES6c5cE+yr5vozmhFNhAkjmKkfusg9m0rDTXIrTV9HPi5RU2pfCV
Q1kXDOiO7lvcyCSLs85JyhO/wIzzrCAUMs4g1gbg/aRvqIIx+0dvtOe7GwpV4Bmn
8ND8atCmIvGPkTemuDwPZSJU6efVjcnDyTMKf4rJnE+D0SBsdvhRgJlz5d1DRJQC
tiCBzQtZo90rzIflL8ByQIT+8RSEdOr64rqUWuajx7IHbPnsXwC3u4KXN4CUiriN
uovOa3d9Ja/PVuqJynKNp/p7t8iHk6Ul3Ksg3l69sYwXfpslND9wVL7Qeg789Kjm
zs+NM/DImMi9cNrbluDASS5/SPBlCSYKYfbNdYJDYdDmWtWpsunIWsEVh1BikgrM
X6K6DXjLhSmxmwFARFKz7z6zuY33o587V2LJX2ib3N9iVoOlJF1wrn2nc5JZOU2I
SGG2/fc/H+5Aeh2SVsu/JCiVYFQngDFaQ/ZAcWUH954sRXUOUL+Mu5Jmm5WlLRZG
Y6GMjBsgcdVGh3f6+t9SLe2yi6ldFq/2Rqci9w/S7ssSUQzRAmquxU8jcb58z/8K
4WOQzbcypKSnj8J7kRB74hZ5ViyCXSUeqTvGxuUPoWMBrgyejZ0xZ5eFdJCqLxpc
yj1m9H27hSq/ww+TZtJt9IACRiVFia8JRM21Zy3h2u/GRMQ0m/KOklkTJbh7bgyf
0z8FYc1qGgLWNTgS6SlrWreprJO0ayF8MrgUV7/yWnzEB+YUhTrK70aLg5zGomJf
vagPjkhP93Y5UfL9QtlbVB5vf1jVaY37ItqrT8jCY6lWd+7AQ5pOw3qG3ldP5zVb
306EaxETHv5mai/Ivfiuae1rH/HrW5Q+KMSlwVGSjDhqvLzIuTu1iGsrrumnEipO
MEmOUX8zKeBzGwNdPYPBbi8/3FqVHniOy6sxkGKOoNkaCg3/pDTqY2DMFGbS50XJ
5+5m//+OENzSSztrKGgXMnEWCYIbJiPhBTWPeUisZ4VDiORmo1n57WPgr5LQGbSC
K2X5oO2psDgLjcAI0Pn8yhTbKGYUyHv+W4b4+5GuBjoVJF8MJh1xI27bbxoCart0
gCe92Q7v4W/C44kJwdep2ppFVbTZxyE2Hq6gJclcdU8cQj3uR8Uo9TMj7pLGExIf
zCXpb3lSOKJUUAPhK1VP4If6ZQe1Sj7KHGtkD+jp79mcWL7xwuzGEWrr4YDRBWqT
ZqzjKvfHvWMeiTsXwJ6lrvgzuOCp97YXLPoLuDsWBfm4ikd2aOcj7sQbUvsGPMCA
ONxmPv/jTxi1eM6ZOYv6q4GbzqhhjQxpXM7Ci2O0ko227FcsPlG/z9A6PDggT4X8
3Nne81WiTHx+IIehrlCyqIJ1h2Xr8L01PqbsM1AfMBc0FspiVlyVhLZxUxT6u7XN
clNDVwEEOxOH+zGU1TtfJgWw+QyJojMC0iQf+R+h3QOjDl7wKH2zLsOKWIKHnLT0
QR+jj9cvpBUHAFWF0CpLCchaC3kICFE3g1Ir1tl+ZbukKzOdegIc8cY4uspo3PFl
uEG9VIPn7h6iY17kPXnAjWZ/8JYWWXeNXPgh5y+BwScepNwKlmqwWmON7B1lJ1pi
Jmq22lih4liFa6h4aZunvMx37aH/+nYK3gX8aWxqNA+3gpFufeT4qtGTVDbZ97P7
zvf/hg1VpWLffmpR8BZc8E27zwaaNHaL/VguwRbzJkWbZe7PQSh/zNp/RYCMfyMl
O9Frt5vqjCi+V5uEE/vfLHQ5GouCeJhG9KYS6W7+myTnJ3pCIYF8vE0MN2phpToA
alQX5Wh8ae9wfAOiDMKM7Kn1THfZhIZ6cIO3EFj6CGdMhJRUBlluezuYcDANOJbH
zGqy/F3/0OeCgBaXHshCNmtYgbnLxIid3IGcCfW1ht2uHRecXYh0ZpvYjlmASDAy
/iyseu/l1pwql8/oXezUwS70o7Rslf4smHtnmr81hhfZKBhxr1i+hW9Tf36KL8MD
kYgfH2mHZOFTszRGSpc8ax3+mUzlRSAvCe/7uJp+nEn1rj3sDvaH3TGt0JtVliwy
uR9YqwJUWFCO1qiqAwDT7GZbiZuhLrP5HLqcFJhmsRFr5NXya7vbGyd6Y+MrJz7U
euY8OMHdWAfAXTA2QRevCqXQEip08MLVvU72FoWGqo5aZ9Qq3Y2oA1G3UU3lOcBs
TT6p375gF2sdWGwDAUceMF9HsGLrA4PpquZO4p3q+aOldU/qL1GEtXMTBgwnBRcX
r6T9CtJzni7UV75pLratkYcGnsNnGYAAQcX3tBqWiguHqlEBVXJP3ZjiV3yNQVD7
l9ptjwytOd+HV2wct+SHDiYB6s7nSx1BiN+i33TagKNhEseCGIDA4B9TFevB3G31
GzkWDMUyuQJ2m6hsja9RYj6IiIz3grlulyhBea4aDSxHXrF3PXA/hCXqqIrLTuJM
R4G5xT06ioyJLa8CE5QCaGxIyeZp5JeYM5301a4WinAomOlS1CUtBCcAxZFZOpYw
JCsytvPi4FZziP50hg9TXqXfRkLcEnohuh1Q4wEwBEJnoHlCF9ITI3SNZq2tyNQD
p/XQA112aIlZduhyG7Zz45t05CMMKv4eXnhtJnF9hStv4N6WlCrcUnVsXKqgItNB
0y85PGCSqhgQrXebAVmmpjCt8IaKJcWUWHK2Abm+cNR52TlhZ2UKLls8GFz7CYg5
8q0E/51tRV0esETIWcgEV4ZZ3EYADocgFa7vHUGMrDS1HB5D+DacMw6s9LXBetZr
51+erNFqJt/nhEAuMRVglQBuyFQK1MT71T1NzLWHTyJU9bV5CJz6a6Brl0VmFDlQ
bS+6iPqLZ/JEuC9kr+lJZvV7s7eSEOIShgFyTcNCnHaninT9iFFaVV6byLpYqdSb
fIzOphj1Lra1o54X1lfysWlRJfOIu5zF8cL/PXE8lYRPfuTeSIY+R3O/WYOfwvY2
DP8BgCtgmxURgShFgb7zt4yII2Jm9gvfcyCnxTZCDfRsOmcZeSoujNc03RHUwFS3
h7rs8NaYSk5v5Nt1O+j/o/5DjRWjWSfWw/gpm2a5HuE4iCWR4h6qBOxUmMIX3bY2
D9Mqlw4NJjUyP52hLwTrqwHMWqfrzqjX0AULj6yOatpQwpBCt/U33ARATZ7IPSQN
ZQ+agh64i1XKuDldlW8QYlyUS/1dZ2236DXXmkPlQFwtuJtV2NAenW0r2pnWJztt
2jlElfSQblzYWe3XVzXUxQvpbOGvEcrhvLnp+1/AfMgYaIwJWtSXkXIKwXfRogOv
kLW9aGnbF+u8I05l9Z6gDWDzLkjP9RDQqjKJJJPxjqbtI++lqq31BV9aAsvWusuI
IyiXKcrB01WaNHoCRZIepkIQUJVXPCzkZvzrbn4g+RoO63eb5BnbPj7lIfysERlm
btlgLf/BzZSstLZyl2wk/rgxwuuxYL3ZQaLP3EoXxjM21IIoEKo7mzt6k7NSoDCu
T2SAzlNnW4KuUfh9CF+mQrgX1+50agzt1rxUdfWX9YdCLIi9lt9k/LQyOR6a/vhD
bCwSwRnjLMkZBZRYnW7sGi9UCfv2omsV64852rEk75S8W7sD+yorc6+99WDtkLs8
wksF1VjLXBG1/dvJ5b3jbq+RdG9uZxKKCHV6mYYWMp81+mWZkEQg9pfmFucVCBxV
o53FN3yzYCfu5FxWrwP1Yo1+z6paJyTApnJIVDCpCTrg5fYm4IBXTXznWb98c4Ao
0XJTdssr50Nx9DyiLtepuuAufY4Ahc5uNHX0sslFf4iS7iRJcnT/7wZLB6U39vE1
Q0qqQo1qYl6/d/syUgjfzMRJBe8QxeGllfuaVCT26ZJEhIkVJ8FRmLrsK5FpKP1z
cjb6WcpPHYs0/3r2p7Uncd2uDZH9Ss43ssnyDattKk6EmTSpPKh/QiA4rP6dETwd
1zuwVCVg0F3G39i4SQ12DS+/vSKHBPmqG0bsVghAWAY4+LZ17HjoJQv25CiEGflZ
qGk7TTZyOP9KhDjlh+KKCtVYyu/VmD2lG18ZoyqRDR0ipNc3ClQy4X+BhyyXTd45
+5NjYHrAtBbHcnlLKZq9Br1EdhPUQyWbRIjswKjoq11eO45VmJFqkAnZ5HWqDNb6
NLgXZ385toKceNJKSTHKekDL6RAbYZ5vbUWTmPvSfpcKTBHLUrXz0th019YomMqS
Sx0WGKx0NzUIDmGK8Zy0yn4o2J9sGbG9uLMRArQWlJVPImcrfRN/r1izN1hg0Aqh
QAXadWBkKJUcoyZTqJAO0izUpVa/3k1XRjD/t2gvJilJJahic4/kTeMPmg8gdx6e
hz3YlFrHaiw8RJ2sp2fX8d08tQOmaz8zBv9TwWMU/TD6rrgKPn959nKOJBNJi/kC
uhgimYaN5NUTieA16e+8kAsMzyL8SZtKPbpl+TaGcv4rYxIVHbihq9LG/OX11i6D
7EBawAUjxlbuiKIwh30xXcr4ycKbb7vXyPL8J0uGZqZ/teA/to1NW27T+rDzrv9t
5fN9uC0fCcakUird6lZYq0WpsX/tgI3YFuJf7YcR43rgu+w9ziD4o0lhjY07s28j
1Yz8zo5AZOQXYbvTak3FYdX5QJ2Lgv5YpxJUd6F1irrIf4Bu0LnVcFmMH4dgoKKk
1ThSEDl3xRju5xa2AwoXUbPG0J0C84CECq3zEBj/z1c9uad3GAQEBLxhTAMuoHXY
zk49zAPQRpjFKkQIYZl6MowG1jHsqV6gfd9KXsFy7GHA2Sd+NQk9NlBfEm4PfnBE
gFzmYp9nfDSVfvU8+8NAOiOdJCkuZgPE+4C1TGbAaQuyDHEiJVgTBpF429PyFZ/K
SmOsyOIAmLxHAwle13dBhu0kf8o/sfP0+rt3FrCTnO2+gojUTd76VvUfbK1M+ZKF
GrVy+w5yqEU+uN1qbwdeS3YsfDZXDyz6O264A8osSF0nK3M73x7ajfbOQJi8Nu32
Zix3HLkJ9sC4tIIe/DnNtvl4ljr8ioRgOjBgSif5uqsNpXXiv4rHY+yDvIVid+Xp
4nozT4QQRwkcbYFf3jYvkoF0IbAx6gSrNy1MSpQoV74jl8QsnSZ2C8aCbf4UBd1i
dU0tm3QvzJ+FR6as4u9WRYIHNQiXaYivwN7LEXXpCTMCr9aVkIAUQEG85Q/Uz2Lj
lS27e4QCtgkMMLKPOaEBM7U3iuHrNbfoM7BfH0/ndz4qfeMMSYRkW5S3GMedKvTP
JQyVYMykVLzK97pJ/JXZZQUHDjE9VPm5lFX1uT6XYdUl1JP4z5AYPisVcN53pnIz
IzHzWQhqAUulpGrynK2AaS4GauNEFsPa9CJb/bbbK4eOUmGUIH/idkSSNBy6FbyG
4HMwrQ9SbfnhtPY/m9NM9+IdfrZ+MODbbq1JxIrfCUGeJQp6DeF6C0byZoiEwLiB
+kYLDfV6e1jiqWMBNJvcsIA2YuebPAecoYDHICczW1xxLPAe493Qe/kjoptv6xP8
N/R8QAA/MM39K83Td3lSK9kI10ZkUzlcM/B15E5g3kdFR+1zG40LzGmIf73sAIbv
qLn+gRSuw+t/O+SV23WaRaYxN+vYFpkiqveQTzmFHodBD9pXFfrd/5lQ1+ziAL47
xsa0AxrnTw0gq+7oaeUjxYHuZ3QycAVpkg5XIfqv64H4CoQkL5o6GXM+mB7Br8iV
98Sm5va8Wn11FSrmYAWGGhQA2xy2bN40/gQrlcYOeBUFkEZxrBihU3QS+RvhfjV8
9RuY/3+kcbmIK3kFgpPA4MnKjb5bG+iZ62IIvrG5RgB2h1X49oAdUfCzvd3QEThr
RVBniJ6W3+T6Nxf7foD8MV8T3vED2IIs2mI1T0EABn/hLZQ+FnS9khUonLWOPupx
QAgfk4+UHaRH6n/Qw6qjTtJ1Mh75c6wk8lOy/jpHlJFf1eg0v3gWpCtKB6KXdppk
9sZ/m/vhHMkx4odIoGgOuf6zvnMk98W6MM0bnCbUd5G5+LwhyxeBO664/lFBICs8
7vwc/PncEIjUXtGhDIDxUpUoUny04/GiXktBm66SETwaUleYXV39yFnIBYcq7SMk
ugLvCcgflc1pDvM65ir4NsSIyu/64UkUk1/CvlVStvcajyhFKrKjjxI+w13bbvwv
fV0AMPGHTcdhbT45aZnDFW8RGXV2we3zozDCxmTgQFLNSbBpAuSBZOJcGKly4FOx
keJdSYeYRM+L0wNXVJduuJsR90H2iDI9+8DWRhiCtZlgTZQlp/YnovWLJ2qQ3VrO
ymVsUugHCPIey8b/Jhf9Yfvj9jO2JM3lwTjuKTZrRoDsJpXtrRpDdOPJgFSInrAr
xeAzQslfsfC0HB+JKJq9jRc+Siv5A/NBdg0t8/4/e3FWByuHRDY0Yd8lW07fG8wu
2773pWBFxCoMPopgPf6ilczJPTUHC+0pG/3IbuwpD0b7aepOpvcRRvgzS2H8tP2E
kkfAPUKCCtfBXKV2l3/MRPBq8zxZLAM3hkoPCG23ZPwkOgtFDu2wmgnECXOS+bIF
Zhrf63wwAibmP33KFYbjsZNVButOPbFPwmBaaMFaUhmPHCpUVyuAZNBXopElmLuI
9hTW1/qLJpbOLYTyFeTOpXGj6fskP5U79IgBcajuUt0SdKBHFs75ih/lCME2aIwV
HqJlBYPzxDTETtKeisNrGDMB5n5EXxTlNtHncBrsAERyjhDWg1h6F9Ly5MZPjdxN
jEb7L7S+M3JU0u0urFTFn4yWv0zwfBkaLX5L1U3rByP6g8MLDa+L/F0aAF6STfAt
flqreCeu5n/j5EnRBOwU2kfditqSde123yGhJuZZrzS4i0sAa9s4yJMCmPwi6PCq
MKTpMPEMGwJwr2FNHvCiiJIlXePPr619EQ2q1HvKFBgAj86vVZQv4MltPmOUzecN
yMoacmoc1w5DV+Qw0PtvLVr5q3X9MoAK76CjpFU5EA9HXLuLkSUaGlDVwkyS6L1x
YQ+YZHxdapKByxgszO+vHRTl6EoWevtXNkGu65w7kDJOpMG9xhFQ4GcH7FbdinxE
ztPA7oNjo3WdohNKP/HP6KluprqjUqcgE9tTir+c75dm/rZhtU7VkESuE3oR4oks
qCu8OyD/L0mqkdNBaG4cfZmf1lV3Wp7byeQHo40Bqys8MlpxxdZwoQ58ykqHxEqv
P/T14px41qWBQCypQIcDMySHBcZlHHVUhAR6hzIy4gnp67u7donbMlGC/OMTU7XZ
sW948Wc8qa39FsTVmBx31nsr9a9k4h0cGosZkn5260VvecjOJymf9MM71R3v4Wsv
dxFdtalwlstYAVqvgYSghvcq5bZ9qRq7DHNFbDnlg9OKwLnGKJFlbeZseeGM9tl2
hHBIs8Eqb3H6HBXG5Qe2//Wofen4Y06HgofmIAAczlRp7uP5mc9tdhba2n3t3Ki8
36qWqkKlETSKgHm1HRyxJy1GTnGrSdT0NeC0ZFjHoNrFiTsEX+8m8yolfLobLOCj
HrnF4vW5UM19dom/caoaVpeIP6nszBHKJ5pyI/AiWIB0G0biyp3NSnQaBOd15tjH
PJPSy61/4fJn31k38+Ov76m/5Ig2QxsyQUcwYn/czb2Q1a2GIHro23039yG0tz7g
Ns0ppBmdPGGOXmxYFqp8wVoHjCTiYEbX5rVuEW4cCqJXsmD2mIRV+kX3F7/HHZCn
26deqMafQtb/WSh4KfEhGkl5RVlWi5ScECi3s5DCxjB3o02oBOKbVBpJgAKBJsW0
xXDoRDyYm9fFMzxaSnpZH23hXS2GDo3r5LlV867JaS6Jw/xBbb1vJmphDkFi2nBj
5gatl397BZK/PFhrdAHTsdNEWDUPCO/ye3e3iumcMFiedK5H9yxbkPus2kjDs1RW
9U1Xw8n3Icf18Aam0EpQoYPlCMbELWc3jbhhhFKYOpJCtjAhJvgCFkMImEqABMbP
jZgMkN9qezW7BtWtcKdKwbyK2YwDm2Jddj4NEiiHfLaM5/yqYJwQAHMJO5N8alMR
lM0P7K0WlsiY8qPum3iswvIPIV9Y8EtEIf6y9LbpDm0sDxnvBN+uL+eka4VxkE+n
Pbn0lD2Idf+wPD1DbE83dBjD++aTOqkygANFklDMq2KpPHXURz5H17JSg6zcFkof
aOj7NSOPcXQ40DGVfteeKFUKZf/63MkoSm82lhCMKXdb2jhhWtbOLNgOkkNRFZ22
RQC72v6yN/yeeS+q07YeMxkffYOdbxs8w0+GEr6qBIyK1N3zdK6YjXzR4AJ6pDEb
Sx3GPnyurmQw2wYTulVjsH0EBtXHt1Q8Lu8Ue46cqtFVbbwPRGXFW1p/gpZXRUuN
b8uataT8oylJNUGI/CSeUrZThSkJZkzmC3/6VVzPXXYNTCCmoIxTr4HWkO4HXhCF
y8mo/S1gHmAqJtKlJw+7xmPOE/2VDJ2rX4EBI+PD/o24AMLDnKVqSV9zn4Ia1tgZ
5V0Zaeywj7XoXRpFEiRx1fkEq1GIcYBVIpOSW6EdXDqiBXlnVfA3QYXlV+g8PnV3
+57c8nEPiNsoXDzhWtKLZhl8XQy8ZO3uUFILAFjIIWd9mS3UZ1krjSdn/Gd9AeiN
frD/lVPzX+p9l9wXJAwygsMdyiGQDh+HASFi5R0Y8eeGPrpnDOTVRhXzQ79AYVzZ
grqOxF/so26haKoPEafh+ys0VRb5tjWzFUXt1aj3hRS5XoFMxF4yFdEfXvA13WPs
v4QUP3P5MJ2fb+/Oi143MOmxK2kvj6XsAKMMLUn7tKU+G5tIRXysuxXGZ6ayFV7j
pvJqiKiuv1SXyEqLbM1uIFUPDe0aO5C2OWJArbH4KvCegqG+Ln5n5P/F5gYm2EfR
V3z0S6YBM15NrdnETW1k1uWpkDi6XwKaEa580nQ1x+5XTsEP2OtjmXTD5qg+hHtq
Ru4EBLDPmTYZFYEUdrg7HwSzU/D6ulNNVato0WeTnlAaqwJFhuy+bl0/8s4MGW0b
Ik4dvxRVwTtTPWBo/2/OKNme8mgCK8vvTZQjy9nvwxPyJWj1F5pO0o1jeP0e4kP0
GT8qsg/lUJP8k3fNLT/7lqGZXybDSZHPMQlG6fcUP7Vy/gVT0kQDf8ddvm8ENsfL
rtpuqwGC/rQIsMuzrO6SlNtTZlHx1bmWV9NyBP+xrqSXWC10iciNPKvOYWluXC52
ALHyrju+784au3UapzRZu4Nw+Jh029falVZQfduowpmSe5mbZyNLX+nXrhI4dm+1
wUHmqzkYQPnfzb1L0UufJgXT0NbIIA7ywALIEji0GYKAHZ6nNzs3JBaaWIhIDThm
OHx+47PYJ7ZD3qqcDlEUE0QDyZxZbxUgJdbEuS4FccP/Ml/wY9tNK794F4YQDJtJ
x2VHf7Rfn8h6n1AAqYttRi0y1QDmpaGaHEi267pTe3q3lE6plJAuSrxI8xFm6FdA
zulPqtgFO3rmxSfJzO+BTiX5Ak1neR/upZCWdOLvxZ3K3l2VDXQlYEuNc8X8XucF
96XoASnbq8mFGE4lxbwEJFjCNql08rxpCJLnQMq8jyRXU6AMPhnryo5P5LqatZ1e
bOwqKS7dNQRddTLi1LUrU9eKxuhDBqk7uO3zKYzFqHIvxZyz7p51YiPH7pdT+1cN
4px9K9/G0aWGliqO801XesxjS0BdZ/MTgBuNCDab+lb+yIdh7fU1sX71al8xbgez
ufwqiuMH9nlL6a3+wPGEqwR3X1Um3EcyD3DKdNK0HxEemQbFZ6LziexynVYj/Dpa
fYesEoEGer5k6nENrGNa9OPcWHmcrw65DLP01Sz5vsMY8xpScZZrtHQYk4oP8ZOE
53bzVwTOHyotTT0lwn/XB/eJyCODj7kj56KKSbhlPhgzUmVCcsH3ZrRAIF7UL2RK
sg2XTItgLQTqqo3kxnZCH6E6Y/mk0RRQfAfFA2zQ0baJMJ+o0zsI8OobxVlB9PRv
+6URTfuO/Dxzab2wzOpKk9Zh2X2ntKP4l/4D/L26W2RbNJj3WGejxQIGqvJ0i5e8
hk/7GZREoclUN2axUoZDWBaVI44lriAUtA2ULVzXCS0LQY/IxWOQoC03EO/YJLPQ
xN9Pn957mFWCVC68nIrxt+L3/ZWZfIFcFG96kkoIuUYIjNYoH/GaZIDSKqERAMuV
FeafYAvOPyBrt7m/fofDFucNyahrpmvd6YoeWO2A+Xt6nsJ+wJEJQNGHH6ZxWGUm
I1lMlm9KywBoIIqCUDCQ5dMAJL9ERJbyuxHyJ+BRPLbOQwdOLZr/3DF9wcHcM5V1
zQI5W2BrjXyEeGrcqx6GzrpLEA3fQTsWzyaUYL1D/bXeVv+qy8DJQFHGbbkZazq7
EvBWHnYthbImlzWJ9l64AH3KvnP8+w0jLunrhdw2F9qLoGGUmyMweMdu8lJubWGy
3JQTxBeOp76cQNtRvSo2lPve/1nAbDGxvZTwahdRhjQuH7ZqDscVR87XkYRDLNiy
CFwuCutbjJENs9DEOPeMOXEeCQFuCsSuW9Y7BTkpupKMEm6Lm6fzhTnzmSYiSJXM
RuxlgUVMwhArj3EtnXx68Ly/cq0YpXrT0fCPnVrqchxV4gY45gJht2vAWsJMDs/b
bibHJMLsR0ialP++MIK3Qq8oDPddvkHbzeCD0HJuVpwzILUHyM5VXzwJ7byfY939
ZY3dRr/V6UX4yUVv8L1hC8CSrOH1zaDoD1G/ffP8YJbN7Ct2utiuOdKYAbx7v2nG
QQdFhF+XQDgLh04OMeBRqSb43Cv5mmYMAl/T9LR8fuq3IBIoULh5hxMRsTfVRY7z
QQMnMKZrizXaH0qGBiYarASnPZKQEjKBTehkj7Vp/Clh552vx7uFPnUrwMy8s4j/
IfFesS9LVcHbLTRb648WtRAFUgTcCgbvuruVRlIkO3dJ5C741fwcUkKg27lCa+Dw
fXdMQN9xfOkvnyufZdnvx1x4Qm/QW6mQVEktZL5M54y2YQG5MXtXEoD1aglfPbt+
PoGPP1ilkZTHnILoWkCRbbpNUrFrAPAUrihu+b5VVCRG//1NoPo3/m7RQ1kbVKah
GxrYGOkdVWa3/e28cDIW77VxAlw4LHxIdCFoUziJPJaCzNcMIQzbzH1CapFThrRC
qovQD/xTQTl2LnFMkw/v4/PgQUVTiVDIe+9VOI6xgjPfRkWgp3lx8vnQ9N4h3qwW
38jf3fiqbZju21jK7RIRYbWAyDcifauT6ZJzlTbrqAAMH2IktCFSR2IzAFjkl+57
t/ihFxBL6hETxOIXjJ94rH54mROIBuS9VKv1XQeR2qbQCExqUsyTZZRrzll/GpSa
Oe2xcxKijEysj5FeTiy+eP+6vpO35J5C9lNX1lY58OzvSGiRoazSdUeOVfsUdghO
6D18AFb23YoRBuPWkQeztbKVe4YapMCW+oeqj8g0jrjXxpCi5WUDXhhDj47mK+gZ
sSdWO0sb3w2NvUBVcRMsHYSvope+5ruaYlbZyiZWPLc9oldTZaPkwD5/VM1pbJn5
Chnwh5ml5S799mdErZ3A0eI5enq6MJyv016b84VuJ1FRO5GZXbPlU8TDRW+zB2W9
SMXI1/uxm1Z9+5qLOAPUDiFIu6TljRpx3NCjwOKb2N5Ra5e4qDV1SzhtpUbe9eWw
PD9WnYg27D7lkSejJBGjGJO/oE5Zq+WohLQ3nfWi0CPqnBTyQmx60lAaAg8KzoeN
n6OY64H5OUj5/S6mDY0xUZlimX06EatGm7mGbpLvl6cCKBtjvem6RNQJoLRdJNsH
1NxXvucFhmjSxW4lBCg5aMbJAWXzOGwe3efTMahrcPQYaPnnGNRBWLeDX1vDO35w
U4nRBYmZQQAxTE4aY7F4HDkue+NII2mJ7se92z8Gov/pxlhnZBAm1kAB2v4xMV54
QTEKsQvtEOW1qV5SuSt10I94qvpoSqyJdaUzDB+tnSLxaaXii4FePe3z4jhirNUu
/X1LKUtqO+MeE0tzMoJGvr4Vqnr4QuCXxJXQebuUT/XFo+icON5XjB12PnHlUCLi
gt2b80H9l1bshk5tW8xy4wozRl2XweOnwqxzhFfk1V7kuOEg/tVgImRDimHD/nDk
XQj2p5XxkuTCr2q+1NzA+zN2sy95KWiWmwFjmGgjIS/gjq27qqTMDW96T4RL1KJ+
qGsLZC9xkgoKdcZ98LQMSnZKS5AqVypkfQh1hXidHGd3qS5zOLC3azJGkJsnzvX5
YGfonD/ZQ+8b3L3cz/Q7HaB/1kVUPfMC36PrPlO+vvBbpNGuSwKjEbfxWXVLFjLT
OlZ3SufEQYi1Q3rXTJxIKNVRJBvAvNE4EbYz/vvdB4fEyah1RGLk74+Cu4QTEDL0
Vm9SNUNbDX5qq9TQHybaiQEWs7G832qf4EYy59H0+IOfG7edsinqlkdMerifi7yi
9eRvHE3nhuPPeqyOSHE+Gj00OxypY9haB160MHPsTp4GIv1aaqS/n3FOTt8rmptt
8GaqwCRyA5yNxF3a9+z29DxW1KW29EPWj4GF0AyC2FIiXyR+rLMIGoi+EAaCko75
oGID5I0ft+IBoFgYtoEvIEbEJvc+dBQz/6fsMxfx4CbIdPS4ehtQMh1k5/gystYf
/omUZt9K0XLPVAT44FPXWf7OVhq/9qMqm690UGOrxWnHNgYphY8rutE3BHruUDHq
z0GLRZGvsvqp25Yj3tdKeJoCUNORvcrRT4YPk5sun+X1ZH4IZroxUNWpTTAcAEj4
0CjCGiLYrWjx9BXBdbLR8BK9GOzqwhvhJKwUV0IUyc8qMQOHSPTYwB6oZTopJOuN
BB0RROdS/KRu6rckNbT4JcocNIi7FKCtBnYFOZvmYj0HApBGxCDzNdx3lgI420qv
h3knPxAkAVI9nDiyyB5k2AVKUudBcJR1VUx0ag0FRV7mqu3KH4l2jTIRQL6NAmbt
W69RbSjmC0dsV6mbTO6oGgKj5u3ovxFvXp9cSMnPleeRqJq+HNfSSERfzCiVbxm4
8/lAI7IyWx21I0VjyWmafZ7UpXSqygp8Gzh0uDj2UkbiRjJkuf0iNkbEzLmKiCjx
6NyhYH5dErWsKYa/HOvGAjlgi1lQyiCZAUL4UlGy9dlimFALikcZM1JaHNi/7eGt
K392vIc2lulmrcCsBN79THcmKxwZe/BPZD4YpfxJ1XNlZ/OcPprf05WIjE7tp3XR
PJQAZzqk/lNK5fMWa7F14rYHMinwpT0sRbEIjw0fv5mrpOmBIhboCK7BOVHzNd7B
5MuMhNsTHf7F75meemSiUWXcSgBQYfCD+6w1mZO9T+03EnY6C+tuTPAy7QaZEtVC
6d1rTR+MwT8MKbhj5Nl7L3Tl+sSKB4z6sgdWyi9BoL6wHndvITzUFg/FOY8TjXJc
dN90K0Gn5ccgKfQ5qC2KivD/GmK+LX003wKNzNpjzGkQDRDOBk1uii+qhwU4nOLg
ipTvM+cLqle86EtPxGYFASrh3DMCbcPN93kXzPjxxt8jbi8XtcQ5wgEsqSA6G7Ms
MksViJ5cPFngD6bQ+RoJnRXPxGjv0ylaS3TZoGNiY2WH4c10nQe8saNDAa+FqtWM
qq5h7qu8hFSgrastq08A0Ide7PSvHwWycHGtKHEpd/IofyOsvzboipKYSoDAE8gO
uQi5x5jRraEhPLGwmANqS6Uc9uFZ8kozCxTwIOuexTVNzCg9Flzj0iw32yJVwt15
RBCTlIJvjfWIa1wEv3gsuIIlUKOy+UDrR6E4IVNMmnx7ehMCcvmA0Ih1IEZWw91O
DgaxaS3h7EjeBc31W44Yr+8aWOXjngn6D1N1DOdBjdvIYGJJGr0ddUFfuxaFKQk9
It+KS4DKl5X21Hk63LS/35VGVeePfKmx3eVF+XGgJkjCTkT3PSHEsEUsieok5Hlr
a7RuKeWsopsUyEIB4/U6YWb5UoDwVUhXOs9X9425j7gtE6RdFxIlw6Ct2xmf2Rsi
sxpaGUxUiTAc5jPE5bPdCcwvEhFpaKlsDHoutMHDgYhYpPYwG6QxclsAEY7m/Ez8
n0vj00+IxcuBir/1hFAIBdV2Fpi9gbEXOtQOh2sM7JqxoDkQamTOD1+3yIEdecPm
lr4DW4xJDODU0LNNVAMhzZzkLMoSnmBbbLh2vdNUipKnbtyKxcrr/9aSVt9hX0Ek
/9K/5YUe7CbUmszxbnRLWh2I2mrHFiT4+LSC0RhndXtiDywGqySUdTPYdU4PFY16
EKcxRcqA6pRu2CW7eNKHp2OZ9/hAr6llmUF5nH0gxOK0jrFhF8kQfOkw5CzXzI0x
GAnEIteAAyCS/qPBO6vxC0F7tF3brNZDSNfIAQeA/EYcwt6UfMzH0LWqQVWjbytb
kUHTUif0hTrxdLWr0jwvLrqofi8XxwLFsDtYp41qBr93neX4q4ogRHiaId7/dlEr
R3B9S1eVCPXnLfy1TA0SHyPsOrRhUEsOsRRyLD4Hh+zlpoK2CJPUA2Dym+kBGXWD
UvNLdovUX1aR8TvuNvkWomqQtOpFgykw+Vz2Xu2rOxStk8ldrKj35bBOFR2nloYK
Fn4oZNspIZADoYop1WkNy9bqVc3RoqZrDCikwoLA0x5oUttg3R50qou47ZEzjP6X
+8BQgQBMpvrD9zLgOXTZ/dD0oT91VR3JTDLtNAP3guwteCQK8Ex29VNhTLMglNai
BOirS2hp/uP4D9c6w6qsqIqMFZQbgnLLLCp4Z6V5hgXteUafAU6AgICCxXj3e3mF
uQA3EIth/stSezEbNApGpt39B9D24Y2FsxN781WSfAPJv7mzTB1z84CHpcc5sXLd
uE3NkmaMSA9dZk2t7pUfK45/CQmOa0NCj+cu9cNBlkNaAId5+9u805L0Cuk3JT1V
p+CFLLCC59j06EO0VV3lKPrj9Hu/ejirzftTxDvNKDKsOLedPq6o8MW/vIypPbdU
nxz59IgvMMEnTUiNW1Zabaeq0bKPlKn7JZTvaE3urvYnfVb8N+UT0IIfwqYvxZ1S
EvlvRrK88emwUGHZvl8ZKhW1fmh5TwaeOyglcL3jpdHxEqvP9g65XoIe5Kk+kIAU
BZzDoAdw00zMxb/+jiqrdi8kqqMW8ZnQjaovtdqO3DIyQzhWM7b+KPxX9WKgpanS
VKJQbU4k4iMhIRgP2L6eao0lKbCDhpcDnYSzuDdzVR4YBFWuhwuEOdbRED8jaiw9
+wQw+d+xwKY0Y0A3p6Z1pZv4ZRfOsy5dzm6tstYDZpz5azeBIS1aDfzDi5W80Z5t
PlRk6vu+8N/tB4oBmaj3H7fd19qxdZD+mAmjgAdKTtpT8/Cm8RCaMz3KZiYinxVG
LoOujzy+EIVpU+my912/f0b63PJbzqqZNxu6ZWnWpMAKNYvx/H4kVU+VUK1tIA6F
Zy6kYnNjr0Cdbzbz8o2vmPUhv9n8wlnlsp1uiVXNyB8w0DUOjJ2RPg//23tGkSCG
lXgcM2CFpm8//XwTahkCPI/BqA87czE52wCv5UyG1kZikIzs4u+C+falIAacexVS
GRG19ibwqv4lcq3TZopHNbhRDPe8GDvF7a5yZFnEsiSay8wkZOQ8agZTV7trlr76
iSYBiXFvHXhxy4KlUrljunJcWDirCkqApWihgaLbyFz1Xs8cdDOYGtAoezgZjN9E
ze80JuaIfCBVI77rQ/0mzsI7r5gezkmWEY8mjt/J+Sb28zm667a8vAy8nk8NyUXX
IjYgyXqg9yH2mqbC0h1wSjcKq/UZcco6DTlVU12XwG4hp+E91siXbS/Xp9517gE7
vs/TNQd59Xm0uqMnL3LHprVQilaiHblpKc61cANYxfE3mu2k5fz4HB4XHhULGccA
fTSE4ki92XI6F5BRSX05fa4Q40584nVn4PBUGZqIMCnKthTgur6kRtm4xfMK6hJ8
/ZbeUfZtvaxVgGgb4ls98IDcl2kvwbAtiJRLs38gf62SGagy9Fp4kNhdC36YqXfE
ERft+tWPBvGarWjuWISsh6FN7a+lVjonMYEpcviTT8S/jlREbte8/IhfyCIl4q/P
iwFdv8xxJHg25bIh3nFlu3EWS+NbFsr0i/UjwWOkFzj3HQacj1qOLJLDcB8wuwOy
yckZ+2sMkPsWhnxwZ4219A9KyI52oPJquZ2G/gCDmM4iT4bXv1UjvnSW/EQaWEU8
HHg77qbcPH94cAvjO1HQXzzeB7zFtrN1WFfTSYL+A+LbjYVbL438p66GBt2EU94k
JXemkH6mYFXiEeDQ/U9NhYlbbt1rz/PXhpVcOU9UKrd3etd/U4ne112feff/QyLw
WcYaSe/hXMbrRZ0Dx9L6Xpv0HMKt7RvWlIOcdXJGvXZD6/3cJQMr6dlj/P5l/TUk
1fyrgd849cVBn2o5ze6eaXRlxQI/0J91tiSqiwpUbulVIknAQ7OJfDAtGNjBt2EA
7a9Ouyk9OU89dJsZghsI4H3HdRV4xPxf368v5XBORe3tHXYSuuKYISuRm3dqGaJH
Ljyf3o+iJ9G36ZM/HzGA0OEQ6kr7ZlErZiyEfaFK48ubKsr/Z/KBe04YL+b6g/Bt
dTsyANATzKpQgPh30KiDya7y7wI2CHLTQTrBuIi09zAwmVI90m2y38RUwYpJAc0r
Xh+RXxPFgxd9XWqUYxa7H10PFQdydcMNSWjfC6PMxxGG0XqxDOVVHY4gnD91J97z
bSaJ4sRgSQW7G4tt5m+xFlxrK2FafUv9c7jAf0Mv3JXQZrOdPDYEBxIm0K8rXeyh
wDFXaJ4Mu2+x3q+HVwMMHzm7OpGvEPc/WBZAoVsUV8IshaDChR/NmVdv+ohnJGfE
NEIOfLAsj1RreiCRPFAS0/FwIDMuKOUlmYR41SxoXCL+88sSKHbQ+EWnk90jZIR7
U58fstiMjS3DQbqv52jJSNfYEYagBCew7whTKAiYYs+eYvHw6CUWYBiP6e2eo/AW
HVK7cWxfBBqGDnGrye2oPXjTwHO4h00bX5UKrBTl01MgxZJQHIzZKc66XVziCz9t
kYNXWaLPtw+zOB+QY99fHSIf7UX8621G5bW0SEhTd76XEiKRf1zUt9UPcLIVM2QK
teI3Ay1aAvob+14V6JtC+xn00JOrgf3RY4cVp1PWignWlsH73Z93Mqn8evgfjJI4
m3B4P/w1xx9QaQJvAGP3/LRgARoImmo9iBQcIXojD3udLY1GbtekvO1SuF+ZJmac
nlGa503Dd8etdnznRImy7cYTcsAeBOq9rYSLLqAGbKQWbhiMjmtdlsm4W6EXIxyR
vKfoANLGcZplY1vVmEh05Qfpp5vj0lI+GmDEcz2of7SXXT3ZkrE8N4bMpwSsHb6w
VCfn4dp5ueqa1EPRPGByiIpvM9MMvHO8kLLyOzGbYqN7bra6stPurw1vngjfrMJ4
XDyAF51P/P20XF7B5VzoPqVTjvhXQ7Pd+hyq+J0PXacPxPnGokMK4CySIsR1gZiR
/8E9v5a3+DcRcr5JosHv2k/GJXCLKXZFKUzaVDoU6dW0FQR6ubk22nm0YxGsPB8t
3ajJ8xwyKFOf7fH7RcVDLRWfSYE9J/SEf5e3gOTEfE+BYq8i9sdwsaFhLPZ9DpIo
+aU0VCOCJ3vMUurtgjRT+prHDAwjKoe2WcSNjqDUkzlXGmKM2dIRc0XjxyqaX7ec
5ysHxsRnVbkUd/gc0G8sdN1mgXxWRJOww1frLvon1X4SATQ4Jv+eJa0hWylL18bZ
Ex+iKGMRsNbIUWROH/PgGBZtGXXXr77Mx4+OZ7fw/aMesTRG69dCt2A9oeLIPoFV
HWw4PRxrK3UP+QWjHV7GnN4pi+Ipl55c9N2zSr+N8OER415N4hU+r1sntN+ouk8v
xSQzuSS+IKTib4dOgIdq9BIe0i+Cq5ZW2/pP027oWYat2plbKmBzBWAN4vVs0Qau
x5pHrNq1NSHJeG0wexgwehhIsL45fGHUw05jydaTrE2MioBcr8rhntlh9IP/Qx7g
SdR75cuh2hqPCrQ9D7RX11aIYtACbYA0iLy8cxLUfs1cYgDysWMjZWNJWmnh3p8h
cfozfW18rhUfNXxyCCzgJ56IUEYSPDpzoeBPJ910gbeCsTLkZBi2GMV/7fXUuIBs
QCCqZAVu2WMO+1+YdVwGICVxBStDuI90if6PTjv2FT+J4/+31LUr8PCdL3XNs1j2
I6pw1fV4PvzrxzrjMj3UGHO4v4j/EDyPItOJb90oVc3Me1+XUxRASUzyxFAXcl3E
LO17CcFnOF6c/Xte9kzQIbmZ8ReZedAkup4ht+YsG7MxBrRd356KZL3eO0VDSts5
UcHhK3mZTGM9uVVtGqjD3XO+hdkEnSN6/oAlyrOngUuY7mdzbQKVaj9iH4ralOYF
y65n6l+Px2LCuNx+xhf5qzOctz/joWfDeT0QLbk4Ab3PNZK1FHHcIDXYeLmm1nK3
ujqc/Lt2XkrfKNeSeFwbakw0JIAx8+/3Sn0vdIVF+7vq/gpvUupechkV18LUtbjJ
nwyI5BjAb3Hi92r/0CYTCtObYqPV9p+YSCVsEWqbfD8T4u0covJC2eYhi5wqodxq
4WTBAevvC+65XzgFDsWi6Gg7b47m7nnT6do5AqYyE8grTwHegh6E9QV43LNKQm9F
NDFH7t/4c9YPlPFzcr0VjgDU+8oD7vTDjUPIIa82zsnVx1jrK9jwQoQqf9n4jlOP
Z+9Ku6+tk57UYDe/hOYYbPubbHxIU7kh/cnnJSYeeCDdXRP9dXqIADQwBWkGfymS
2CaTy+dRNf/QbusYmy6Eb2rcJ4YEvPIHk7xIvOdIvMnVDk9+kmsz+iYJgKMI2E2y
EoTKDVtehnGEf6whPFSOhQCHMygHDyRHA3b31DWEYbGd9ey5WMX+FePv0K4AGWIn
1IahBrcyUBYRcFDp37fz0DYHlRbGlhUMkm+M7yOVq6ArDus350/HQFBi1tYMvZCM
lSZ0ITy080tjgr8QwsnWXDTxyHIjMPLYnsLzzuPMSJxVhYFoZX45UQqNUXxQapKN
pYI3zZgQ49XNVt6yY0gwQt9WZISaoC9Zj5Y6qV/UcAZsNASHUSS9U7C2B+eWE7or
sxZQPFQLh5yzAtDYT1cnf0dg20k8qnnEdfRyG6KvqElBzhxMsQhlccQ6MZE0miA2
WyNw2unfqD7lwm0PswTindJM+mV0++RuP9m+bSUg2Y5nQAXrY/kjtOoZLbspuqQM
mJSNYeNWDrTeQYNNZTwL2Mi1esJtMMITpG6FNcDFy3yEmTAjujQSk3WZdFnJajsL
ZTH3FNT184O5+SYCFPTenDp87Uhgli0sqFK8fdTW56b3rpgncImVBMVn7W8FMP3v
wdA8EHPaC/BrXUVeTnVCsnS/BvrS6k+X4u7k98zUrdbjMmqdJKFVhfpERx+d3zug
K1ZlMx0GwemuU0xUadDmUOByaEMz5i0IB7ls6lNA99jYj2qMsLOOpcRqa5HFMSlr
SD4XL6IIOvt2le6GMMssNNuhYCmLH63A/EavxbBvkZ0m3M6ixnLJAkCWy2mQr885
M6ehze1v+OiEVpXFzBkIaTowFYLVoPlqv2odZZUwNDNtdcJuquWbBp4ZSnZchpPI
uaY3QZWpKKOPvkdn4NPE9vY+RSDrLOnjQHgA4YwCIZlHvNpMGaOaiXaLnmx0R/BJ
mUslIsJAjrkx4w03CAGKdNDGTVVQ2t4DgNguW+qffWwqp4cwCEKJ0R5S8lw6AOn9
jMrCEMPii5HkCoZZv7eUqgF/2ryD/6FfFpyltJ3Jtli1jWDteTTHHyH0XJCGZX8T
VIqqBpVLazRhj0Dzu0jgHmiv2NJT41tgJ6tOdMIb5l0LO+o0BwYiScQpRHZxEntP
hujKo7jyQRDJCmzzJZjH/Uazjh1Eeyc+zDK7iweIekcPCiq+szPY1ivioVE2UYeb
M7DDU3d1LfJwdh5MokZIiQ/RsKjKdWz9xqSZy7irmkjBGRlG9cNXewIDJ+g7nvpv
jQ6dX9kvabVJliwlUDUQxqEzVi0BNWeeqMI+HL2Hv6wnpudxpnKFDROkLdzFkh1V
p+kyNwRq9T50EyetDGs6NiGuD24N4G8DVPCxiiTZAj0Iwi96WC53gBfaF1TRGJnd
oQRpjCGDbLBGYTeLqhJel+H+80q/hLp7HwT+74le9aQ9IBKq3Vvfio0f2kyyNORT
K7m7pMmOt1M6wkgZAYBM0wlV/x+IJS1z+MdFZvrLY5Z/ZWGhnpXiNsiBo2XkORqm
pbtORKvoBEeV70k9yPtFo3rkN+PcRgzB4iIndFQ8hnjTiGiwOT4mXdUva9JXPtbE
KdPpZMCztrnfa1BCpblkw39pY7+iqcSNYq+556RNC41K2nou8zXoPxK4B61PsvxM
Dqa2q7HrdoVNDZBaLMDBxPiw1vEXBSgPg+at4pHT27fGMxPDlOc0sOZ4yxHZjq6G
5dwgTJTF+4ahZdEF80H6Z2vRmKgONWLAUWHa3mECA31cDANIeSAjCgMqsNtXBFzn
teW7x/0gkfao1U24RAXvrvHWBcuzqcX5UJ1g48lmJYf85M+osMUMNQzjmsIfzymQ
1NSNOUt9iY18pb45q+k6YyllgDK6HxZ4PPZ99uTeS/6x+YnjSvOqjVhIqhO0MfFU
1a7FJuCSrDkZ/4rttDIwzJp/KsIK0kNnlyQhMJ/sw9gAUGa3laS7ErzCLRabWkNH
qHDiw0yzyabddXhvh0ZSzqtF8Kv9OxJ++l5cazjEaBUgoNS0a0X82v+MXCFCStmZ
eMdTgs64ebR2vwNjJtQywjQwic+4KD/R6njwDAzcmwYxRcEhxRa04wQM8aC+ZYXJ
9UCoYJ+Pmzh101THBrmlgPB6rfQLxmsvr2hxIbCo6VtNomksUxyaeuwNZkYNW6T5
xCAECcidrrfzI8Unt+tBChakZqgZSuGc44ifE6ikeMKJSLm++UIUHWWitwQOQtVy
GmDssOwCe9VDfwQMNSkuwJUoGNVqNTmEPQBCSQ7oe3fVLCoFpP+2zgcu0cGliESk
w8cDxXGvrzq/uU9ravL++zSBYZGxxQZAsD0B4h7+mWLqfTseONTckiy5L7uZCleX
SJOhjrpQAHFW6qdv+Lm8p54xYRCtFIVVihqbrUjfS/9GuFuKbQTjg0RYuqXD6e0b
2s548dm4CyKAf4O0J9MRaBJsGP7JdqbvowmnA20Ke6JjaT4LTY0p+dNAcgBnjDgi
79Fc/OrOH9o6YltRpl7B/X0w+v2Dcc4FllKQU1s1GFF7FCaJtNu8/vDOQAaQcrlX
zPydAThi8Ai32NurCtNMn3AtEFZzVTXrg2dTXyB3Y33A/qbmDlAyo8UVDaBD5+r0
hHfdDwlOJvOGn8axY5dqAGgubw0Q7n5jI9mSoZUZAMkNVgr0mxwckAYaeBeQOdLt
JuVXZIzPISw1FLUl6SANtaFniX41GHBSpwWUEPb7hdaa+2AatA1cMMiROh3G38MP
0lHPDd8RIhE1yiKNqfGJTFeotbCRx48wXQCsjuhct3cVhbAp2BaLmF2TjuzXvqNp
xc0ouOktIXz8bi9AzP/XeRx/OWrYAldcO7e+zaKQsS1Qrf0LYsYa1UiI8wkS6Lgv
iUM33awonLCmQ1LH9xgnGDn0WL7+Kk5/AQCcZAnV0fquWQDVV3EVIfbCML8AHyH4
m6NKqJWgMsxvaI2zumGamZb6pVE+LOdJs9ezBJn/XnFs0mCp2TjERGk2ZtSD/UrL
6H0kNXpOgvrEpyUpaVS00UM3bdQ+3hH8ijPdscAy0eWOHC6Y3CGmmZXauv1hha7G
5NqK/yG1Re0zPhtHBOujlXLkOL7Vepxgw8BEfkdv+biSjaHuzxvjEsZL4XxLC/Tx
bkqdYu7rI7IzW9klEmZSqS/k+H64z/Oa6O41iTT1dVS52RngYumJHcSaAqV7P1rm
vv6wGAWt9EBeAaj0h7fPuHlJmX4puIE5djBmxLNvnUffvq6EFXWfpsHKO7FqQPHJ
yc2S85T0hwyirH1EXlu3KrLrLs2M7SC1wyjMecn+JsehtL6ydyH9zmIOSdXuCRKZ
ZY1GfPhr4fz220vyZJdBVpzPxa1ifBmP8v7YSeS+Kc8a00/05PaPMrPJtJBmNCuo
ifahOzdtpWgFroGVbiIQ9DM8aCMxRh8awAvYYUspXUWVErJSWPYyCwAGP59Wp9SX
EXgD6NQTk8zQJvx9mkuogwNgvFfcrA7PncPqv7wfE5OP8Pzy/3PARzrdtAW1Xo7R
Fi5bGGtr7Yd0KXZz+LMSrErK3YJoBjI5YAjeRKRGrCAmrUjLfBNv5gOtUknDV51P
7FNTx+qvQoMjtacHgJ90cWcPdZSDOKcYsrZP7vAjY7bfXjdeTWTSLU3VkT9WjXZp
qEJAq7zOeIrq/Tjw0DknYMOnQYcS7SmT8W6UiQ4mmx+VZCltODR0tq1P9/GKm+Qx
81FC1lv3jIN/vSQkLQ/QS4ZIhL2ED+++kp2yWdeSBlLqjq+kwp5wdCilsjgzg7ua
6v9zlHKeeI1ET7FRnjnOcCwE6NgmVP3CHFF2kQvJNkkbOfW7pF8afZF1unrBFDH2
yheWr+2ZJbvCj/Y/nMFZxf0gwwuaAxD1ElW4Do/HDcPJ1yJuQpK4D843SqW+JqGd
yp0QKSqSyFuG0aBrH9VZl9HVz69i7Sv1cs2zpWOnXsFE58+ra6RSpjYVDu0RIi5T
JVKTCGG07UVwTKvEDIzmvTDNgVOy1ME4wGbcSZGP2YsgGcyWw0pHS3P11uDqerVW
oRjHla9FrfVFcyugzvGKcI7/Xob6SOpJJPG7xWTVO2Eaf1hJyK0BlPjvmGD7TmAJ
d6PXHMXln1TcJrIS6SDOnE0mV4CTvm6G614g2+ecs3j4LCQnmhbi+9vPzWcuL6XL
MqB3Vpkhd0Ik5AsYVDhLEYvQ3tQfwca2kkLPugGzfhIvOglE19yJFz0spp8GhgB8
vxm3eraM93Rv+yCi+iiI+Mkxu7uipFQHeZEJiKePqvY28FUbBWukCtoouidPEkGU
xTPf2BhKHKPiDKN59aN0X44d0qkl6AHU2DwmOPhrDoYuJhTywIpEm2PM6HMnsaoQ
ajoZYC+M2Ll3NNoj/koWHAABIXcVc0FTYTUtNwXsCqHV2dsJg0mvlOOG2+0AcgzC
W6A92HU2RaCtg5ePSVl1s1Xod2lFpCHrZTq0kJ9A+ladVdbi32aebbCrrHvEqROF
v2QSM6CzFWGX7UDgef9KcihfYC7CjUZnWpzggxo5PwxFOZpVO605ExqYQCxbqHkz
fvld5tGKG4LRClG1lf0HjFaneVnw43dZhXWOM8AYP+PUvSWqs0CDJZQkU0ZvKrOx
HdoDEsmOZGDD7udYR7WHqwcc4VhYNz72FBlAv+3TFkxa5mHh3pVyVXiGm5tvh+rP
IZwiIKRFiN+0drdpE7U4zFMn1amCGWznBLMR1+yqpEn8Lea+JHWOrULjmR6erkrW
nz0vupwZuvMYzSZmLPaiVkFfGkXLJB0tN9O6ag3RpjfyKxEboDoyidFhenzgWmdD
Cz/LBSZJfUFTbaYkr/SKKOMoSIW5cftzJ46I3oSbN5vLwSDeT8L7IkzZpuz3F5P3
it4aCcWz0AQm4kZbLz+mdKaydywv4dgXZZeJ+VzS5ZrHVn4A8pk5R5XX7F1PMMmw
nO82+HdNe7uHTSIMFqePRoDx8KcuQ0oowBawmJ4oLXHDwymscvO+qDbqKMprRyIc
BHfSgqB3k4FYtQRImc3v8a87LRpYGE0iy6QlZ2kJxdtZsl+ZoGfjePb/GrdmKUuV
icUgnh/8Ou8qS5ya0TtiuGCOnlfa447BkzXqHDBExNF2O2OpFTg+o5+yJHeVn60m
osi9+x2oJrH21gZVKiyZMzmaEMu131RUfkRV/NPJ/wOO/7SSeqQBfdnRcdKiTRob
sLqwGl9Bt6rLuBv6UgAzZmn5yCEGDWSlx67JrIOug4AKQLYUJtPjsrmv9yTmhH0f
FvSBDVrzG+MPReACmcJHkdl7k0U6W/2LLFSfXG/FoG6rwBUA84OSd6PgJekeWW9t
Q6dLX25ntpmocJE+ydekVHnNmtr3YSBazZu9cNOfUQlJPy9RoquFhBVTrgicukYq
FXDGbiMpSH2oK9EFXFIuFdfIHZ28av/s8na22hyIaP10CMfPKty4gd9TmluwdT5E
pWajmYoGcM3TiuZr71Qz8ct+gqNQmv+/5lb5MDm9AwMITaWNyvdVAIA4zItgNHk6
4qIWhbjpSA5CNKVBrplkDVqDq0tENUi0B65rsycpJHVQtz+Kv3N7nL5+XAJLP53T
L1INQaDOYuS6d6fxIQIM+o6IkFYr8Eq0etL74xqPCRcJnBnQezWWpuwNTyjg1IRH
oLCIpad1BZBd85aFKUtwbgjEx4bzzlj6lFfay3Lqb3jlB9tdPrukqIYwbC/tT6Wm
koS7E1vZF5zvKsh05/oTzs6ILj9eZLWHtYQ8p2YdqfM4hSB24wS7jzR6ZzAheCEK
cGRdl/3p+aSyN5LLUEyPa9hyAkPNg54iZE2QEwsxgP1lT0EordIlpKLFCZ3LLKn+
0ExjUlaXdz67AzLWCoYnuvUyLBu6CtQE9F9YVOdvCXq4NiBAcz/SJggHGkXt6TVq
6WxQyZ1ZzajXpwoTgiFwH4k0ds2Ebpsx+iutoUM/L0PhfzkdVriTiVMlnfwtdX73
9MwNEoca0yj51EEYpaU23Cz3QDI7FxBRnc7lTLaub3bZ6ouA6kvUv2ESNrGN5MBw
htMrGl3WbQCW2YrZoY88G5cF8nsRgl8ZbwXt4L3ovSXJAmqsDEWWMQdejhnVUs2C
YLDCWx/5M2rxv5FdUidYReSwE4TKWreMp8+XJQIDR8S23ABcCPVZydv65nGGc6IN
07DB2RC6kxV5u5EvHakqwPmWQHI4h0+l7SdlabY4Umh8ojvlq81+zbYqFp1KtxhM
97WrHh71snPkNXpZnK0nfezHm/KIcwAadvzxXOv+s3B77U75J44OWkWFg+563do5
0DYo5Kw06Meq8HnltqcA2WjCyc+FJUgIon5hELMGSQjokWSeTQ0sQ8FiY3AKS4O3
4zjDm6dRxSrUVh5NtcIsMAu3m8hq5I1NsWMD3yjDCFEbz13JADkeXnWr/WftCAGr
XcqAL3zvzVZNYzySivKj0KJIWfVyWM0/Z2D+5orhM0o8fx0iQeC+5jL9WF5pesbI
LJIC+b0FXfUyezFxKthtc31fKyVaiH9As6ReAPtjc1qx9S56kEdg2YuHUShiCiXw
dAVIV4w2FCEVC1x+84DqqjiYZ8yV77LsT7prQXh8z1sH4rhcqmNPyYvr7A9YR5Zn
0SYp/PAfiXFJKDVCiIxp+DvATe7nwvlaZdHelMgFTmYx1sOlBAK7PZIv+bAT7kWf
eCd/0qEJrFVrinFy234NqbtgZysrp3eZV5f6537G8uB4su5BEHW1JY8WjLkz4qEa
noqA3NyRJX9aM5qzfxdcf6rxkEBp0xNNC7sgrtXAElxO6CirSq/qheeeb+SWus7o
dxEtPSmEqakZ/f6Y3f0EbObYRDZSf3+Tw0Fzg1v1+RDht9EeQqSv4QYjjCSw+zjs
pclyyXs1Tr/gCD8PT2aOovz5u84pBTN/BYAzI/TILABobc4Yhi7N/yMyAixLKAzF
O94Y/YTTtQMsO8jLozwgQ68bksnUwSCTRwjK+56y3zQTfokdv5BRtvFizGSSSYPd
RULUptNrrA7yVgaKz8U0pi1tEOOh7J30JW2c3b6AwTb7RFPcfu2u8kVveFtAHTKi
V2xWwgkDMiyNL9pmrC6SbiGaX6RuiTQdk4XtTtTL1aw3vYIvvDyCHkWddun0vTgx
DTS4jNZWzo/q5MAT2RY3539upYj7J2zz0o8kgkvjBTcKanerIadvSu5Rjgb8N4hE
S/uB/095rqlGzjapgPEwwbMiq84J+2X6WOcHjHO1c9TE34EH4XwNWjXnslFRlUFm
ol+yveLO/204+Y893qSDoLK7k636jUhKJyYnZU69dvNXvpoPk5UalAAnnvbb7CdE
+djsf8fz1L3voAMW8/riDyBHiQK/0umiiK1Vd3+3Ipzkelw9BZUWcKVL3Hexgs/r
m+WSrCHwRg9SASGx05baovdpF44BZeRCb+f4wGsCV8i0wMQNZuHcNhPAjIDZwYeh
tHr7DHUTRjXolfwYHh8lQcwaux55XL0MoLPWzd8vi6/OLz04ApIu7tLYAlHx/qiD
QYiQS3FS9yxedupDwlfuPP78iTS3eWIt9IIFMOy5f1VbSqy1447HNo889ogWncSG
cgKWHwkqnBnUdyn7zZhrkAg7l0fn4kT7d/e6lvyieFMIeubTrT2YXmx/iSeoLs/7
/VN6N3zMKzGETVjEfPpyD8sXIjlzeSQEAXGYbeXt9jnOR09u32/LpImiQK3RLvQq
rEw8HptBociO+ioEA46Mgns42ZgJoIVnHwvn8HPTy6XjswN48/bAO0D0oyBTKkNF
z9u6E8om+0e94YKvyKzIdmAEyPDTtPtaG1M1Vz9eOq4u4cleXfQUC84Yf0H5eAgg
Fbts/7BCawF4veZ+BGZdb2ppYu+T7tZtzqX+uJmjsl6MlIYkRFWlZZP88H95z3XD
LKq3wciCfRNJsdWWOlhpFCm99D/XB2YkU6w0TOsnc8as8l8uM9CotCfT0goW1DcG
xOHeNmL2cdu4u1Aqy0ppQQbbeLi+Jzv5OOazyFaRlU9pjF+gN0CI1TjxKKdLViTz
oG6g0UMX6cruJU/X6m2dIgJAjMcGr1NWY0jMkEWHZKziDKA0LELNVB4FjYkiyV7z
KZYpz5T3im9FyZ2O9RNw0r1H+Ue9GNvhck4BWC6wCWahXsTgLz951VRr49twY8zH
dFh+td0dqG/7oEF6JYrXKHhCU4qfCBWx6DwakFIOFpPS2ocxdaJvV/ZV/42TPr5O
GtyuNiwT6YunrS//BuGeE1HpRys8aepZWMgSwJk/7GSjfAZ+La0w7Tg1qTOL0pMr
0HcZBskdUH9xIxQVKbsFrRdTPj6Sp3Mntez49LHI7PRxlSyfDcpx14erSHfF/zB8
I8hOqotkyHi4MIn1NHS9HzMLXzg+rJSa2qqKX2InQUl4dgFul7JyGXHCOD3Dh0Tj
kjszPRca85mRUjDj07/FhhiY/nyoEZpmICTo7kOurutME1wL56Aw/lun9T5CXefQ
VpW7q9laXQPg4VDRxW875g9hvv/5LJ3EicsXqOoABlZeifrAjszYN4oOcH++dQ9P
Nqi5N9fvjmpZYlY9RBHkz+p6njxqpkwhHia+4nZnRr5h/SBE4EQ9Lm4ZwibpRtJ6
KFPn+eu+tc/TQrNNnX7KRRbJ+TDaFzruPJyEibHIyZOBmxjWgo+nnLCfDBv58Dnc
8Jv2NZPnQjCqk3zckosihIsU5FBXGlGrYnegi+IC0IKJeXW6ugARp5OXblWYclCD
Yaynq7Rj69l1b7T8dqgxEFCUf+rxSWj1nveXjupRjNR/ifKmAf1gwu8odTu55rei
E94jgWHtvq4ys4/yIhlMFwtgYZ/PBkgefxCP4MYYNzqU/Gjb6YQAZNpWZoCXIWKW
L/AQPGhGe7zct75nAK/JiT4tjrIuXvO9l1T7FzHbm8RPxOA+YorLweJWqsXFpBqw
53OZPfSvS4btm2JgKygihfAmcQLwA1cp0gALfTbEoUgEOw1Smkyum/HUGKAgYxf7
9CkLq7qM8dsZvxUjFXYgvptcEPecb3cutrOhWAXVnaGFYiCKIGpfLESSe8SpjuDh
efwzbFm6CK4jhUsoB7HxF3H7ZfN6ANr3/s0ZIpuptro1GsycvhDVrS44zRh//MJx
0Cil8n0mkuG/T+Yid6JAd/5On95Av0X76Hc8zucYBMs44rdQWudAcPYWg8u5cnhe
GIKNl92QdDN+tUY8IQvgsAsu3tB/BwSgE7wpZVHbpKbEVso27scbfSe/uzg0OtuI
BU7eMvSzZ+OJjHg+47wUsWDrN88cfv30dam1r1HY9PkVaRpoSKZsDpWq1zIYKp45
Nqyi1MvfyWNhQ+BsZy01mNDCk6WlecFVy/dRRK5Q1lBZXv5C8D59Fsr4UvYdMhP5
Vp6y4Goa0Pe/JqDhZwm//O7zyIJCT6pd7J84DakG/f+GQrwzSDAaXlDqMRfjiz4Y
MXXmaBtrDPlBcSYSIa0Z23UEMuPZRLJohCyawtxMyWjynIudIwsoyNjNOoU6elx1
vPryUoYx1BnGGF70ckhnNvzt/drJlS5dxTCir7fSYeVrXoVfddscuAs9LNRRm3hh
CjVoPJb9/9T/ibesE2hn1AMUqnROZbQHsDwAHBnrz0MV7oap0zalXP5c+ZE83E46
4d7+iP7szxgUebgcis+brrgO35av3DBL8QQkjkyQ5QCT2oe9CpA3Gh29Mq4jNRu9
/fidBbHSdIUH7hZjJ877XgEesSDoPhj5dChV/LlJwdaO3YStXlsTckyI/pbDNP/B
Y0O9/qC5Lyi+RgQlm4iOkZv2pxThblmlZtb/iEt5/Sn6mKR3H1FmahaL/ykBL6nj
CbaeBMXvHyL89JozliM0ZDM89qquFL/9WHDMJ0eQLYrp//IWLzKMcu4iwpTVnJX/
5Ibn8jMSCqyGPTKChdIGDtaIddnoXCo00MkfpRfMvOfqTchiB/shKDs95bo5VZd8
1SUnIcdGVPy4Y0gNHIna+fKlOh7hTyD68V+QGUmvwPjtvRZK0lgp3+VhJEwZk2+R
/fae14cjwYXawUdGjxUkIS9FvvvGzk2wteX9G9ruMDPVQVLrM9yZX3j7b8e/lhv0
vsEQfYiDA/3T/aVeySMHCGphqMUrhafU6cCGynOXtm5g+Av+reSk6qtTGu/Mej5C
KZXXDTGIq/EzXm+F4Kimis4zUOjON0YCb77PF+4GAcqMo2WpRjbxJczYMBPQD64t
TWFvfsBx20ka7RSeoq7grbhuDjYx83fRJGyTJKOCmD9zVJ79pJ2JVaAFqKLPcB0I
O7HCS5X+A30zSY51wXbcivhcSLDzoB0tuwIFkl0WsZqEJJGeuZSmTlBePt0UjRnp
4BMcHtfbk/3TZTRpooVO55yv5/TkBH3LoF8rqI7LjHAi3yurwQA0IQi22J7qLn+q
sGPcAIehUpaqmsWYQ18BkOvYdO4JvJ/Q25kbB4jYD9Y/YhcWxvK1l08bSEBEgUjw
Yi5Am3PBwfMFwqyuGYE9jGcZEY3tiUukUz/jmQRP3VTiFds3s+FF4tKrADcnU8xA
a5/wTx2nH6INRsFF6ApmZlPOf8hxoE0+NuhxwhYg+zS0lJrY3kkTvqCOgTSb1xOT
G3YVJv5EuVIkzGlqpIN7yjw9L04EeylwOFtFq+2p+Qd/IFK6Aed4NJ2WWNrzV4E1
KqGPOz2KnKIg+c4w8dF2+iBIost2A0Xx/U5eqYmHGsb+ysJkMxK8a7n0XjnnLWWp
+RgXslIdaBQ2vA3QQLzg5Fn4xHejkZ/lAYI5DgO6YhtMnH1aHBiSfQ2iPvjYnRf1
77hPIcv4N5ztwDbXda0adqVNj1/6pcJTyhKQqeDg7RZiet4XSzOGWBIL8mq7ZbKo
zDvVYewWirC7mvTqMfVfcg6WZejVx88RJpeEPTh7TchUisOcW7bDM8u8ri6bZ4YE
UfqW18PEI1alFnFbEbguOzmQsjmnZYI8ULSLgsifKev0Fl503I87vdcemHp8wbVC
i/IJxVXK38R4eXSSnnjvRplgrNFZ05UQs4MHqyebGo4U45qRp2NBc+m8RQsx+rtf
V/C/tkHIVy1Bg4Jz1+sb6aqK3s4hqRzgguwLBQf4EgEAOXhFO4XvJc5p9f5WSiRJ
z5R+00BJH/WgLBOHUhnjACcmgmCWE9RYgXr6MMjixKWyX1ENB6omP17vMfHr7P21
QvBNz9HFg9WDgD+OTAVO5ymoX5NFCFKwUPwT4WeXZitcJKJFDGTC+LSHADrJDknB
S7Wn88z4aMe+lSduJmuKEYIysZ2paQaHOFz9+pMHpUgLjHd4lVQF92AbZYVm2IYZ
mPuJ0FrKnNjqesbEY0wvm928lOeZ6CAr3WKzfKLmMixbpcPv7P2yu5QFGDsxIjWd
tkVComxOZz3h3OOYdxwZspFskaE5NI2WXDtT7Y3RsuxFhkqUzy+sjHWBW0lLKcyb
o0uHMex+/JYQK1Dqq2/DNjrWAMTOSbp8iDXAN0F5T4IZwIE7u7lMLc05nScHqYul
8IskXfMQLB8QIS4EZWQSBceeoNfmAA7uEepAl9+2wke/770bRphigeMquh+SMTPe
DJBlQFo1FYdvjcklgkWunxLq8Sg3jsXYBVlE1FxAmdTghm8CE9Hgm3vCN7y8HWkt
vDx1BulML6dYUw2L4HDBdSq1DeV+XWHGz3GNe+fWYUn7ETTyHqSkrzdph34PqlcO
D28zA7XqUCidBWVQMMa8dh+7rA/4HH9I5o5OXhGT/7Ch3qkgFzFWuk0ZgsMvAfMQ
fXLF/+kuYX+4yi7GwiKkCitQgc98g++9qH2YJKl5lXR5qDVp4ND1NA+78E0AXCHW
IKVZ2PSVIYRVDeWGtCCsp0L57YjF34SY82H8Zv4THaDRS0dwEmHvLc/bU8CTHJ9A
FOXDkMtptISmbGkjx4i2MP06J1TjFeFfgrJLXoLMgGWLP8fEpSHjTt5GmYbGTwrr
bzCHPQk/M8iPjhW6UgbgfVzOsM1GflGJYJmVXqdeeOqV2T9TrZWBym2S+J1Tzjw3
y00MNwup/DwHL6HzNBUbp3/qEe4y70xChFu0Ff8kJb58WKu5tc4eV6QAWMp0vBFp
2ogGuEARwf9Flo4cTigCPwFSqkVzid4JjWfbVAl43GcNSy3fHtiTb0DH9G6/cmj+
gZlVr74Frk/jpGurX87DgyxEn8MNmuuPnMyGQD4Q2TPI7/a7xzY5uFic+t8CmFWt
+rEAAOCyFTVI/F1gDojKxp7U2CgrsV1jkVOPEcBuUp54HcIKc7z1rfg49ovYHkNQ
rJVsAZSuLmxji0FXz3vIMUU2i6ut4Xyzaev5xJjgM5Dj/8PH+APNflo3PfxTFdh4
jkDHp9ZEJ3umP31cEZPJHeNb+NGjDyxDNyQrzgXcfjMt1Hiq6hDmM36bCxuDgIwb
SlILpJlYsyK1Qb1zQIkQxNjTORwsoBb7vlZRVvN+WtzQOzltvUgRvLSSfeg5FDQ+
oaZHObZ5z9XzixGhxpK3zT2BeJ7TQGtSGN9XB2AU58LPs5NUn9fPr2VwxrkODIEk
OuSCqRu88b8k3TejmTv6FJtjXHUGbbhMTTo/jaDUKchbgP8fYeas6g+/T3fbePRz
ZNYYDmBeBht0NpuNFjdM7hJTdPVm3IPzdMWDv4cUv2rV/ediKDxWbGdmx85wxJXq
hbXCbABsdiVdJdohMrzBUJZvly41n3D4apPzePfzMwifRkQcAdA0EuxH0UTUzo4R
IphRiXJBPEXgMHpGB+rdnqCbmMY6DEPbyHSfpYuL4/0G+bVJdIST0ye/hlRuoca5
4qctL6pZmJlssAGHuT5sIJp3K6D4WAqvSVRDINluKaAASZDk+G3k6qEZlmUceK6z
bZOPXCTj3b55LSXCPST7AVzDNuI4S0gtwL+WjtdF/REwrvU0UwPiTEsYSMArd7e4
iO77yLgRSDvDHrhFp5KidB5iNNuNeYhXWGco0chFvuHuIUBGlwHjIydyOYxXRZXq
uimfb7F5Ybeu5HulqQwLuP2lIygrmbWClvG64QAuTkoUowAW2PpdpsU5tfAsdvGu
j00uQOKM/62P+h6q5C6mdcKSbzS/MBC6HG0rTjM6SfpT8Y/WzfNRRD3ObGUgnWd9
0OTAnTROsoxe8XMhhhL5fl3m6RT8E9rRw4yzvaa/MNQL6TXXQGd+uKOefFW2LYfL
rSCfVJEp5DWjz3YfrHh8jFBvrLa7nkHlrJylglamtc5T1WJdwSDukALJhCnnOFdU
k9QbIG0nQBfBpyGlcVAl3PG9y0brVABZRM/7XHZnXWPWYVLwm/wsJCAjBz0GcSd6
5U2t17DKIDzfF8bR/BHfyfoI7pJH8LrVKfZwz5eN/Ja8kTLdfUF0S+VnYRXOhRnm
pa3HNc5GKv7v/YxiZLgXpP0UUK9e+CTong6DOOyaU8spDlhKnl8AzKIftvuAv1JH
UV4NOScoDLRIvgJsUMMhMbFlZugJjRfGRLpmW1ARoYxfh2ycPUTQw/l9/57Vm/5r
AlIMhulhGIXOmsvYVMow3Pzi+k3hhpYFdZ9uuPyEpgy+0yeevkXJuBHHhmuGewMC
UQIptIw4OvvWIFxBwFJ8BQlC1NPnC71Rlbe8Q8wmHlJorAuEWvNASYDA2y2+/ugJ
UY+mbsGhZOpzIKImxMj5XqwvutEsQftUl+sPOuXqhRG5dHoqmsvbZ9TGGVTLAh8j
7sNQsKvhZzFdxiisyDjzZ5b/jElVWmDWChDMmZN69QV1F3kqBh3Pkk5SckJCVHDv
yPL5PjGXH1H8UkHrc0Epc+YSHncWphvsj3Zj1XeFSjfgq8F/HrrlTUEzMgK0Fcw8
wF2D/axivMy7dFEGAs2CYj9OeQCQs37mPhMXA3Xobmf5waAH9AA+ama4x+DLo71J
dKAvDkhlYfYbtOwM23qO6LFesHbonPtw9vxBaB9er2i0LoE4xG6l9cgximKAX+PG
gfI5NNCQDCq6Z4/FfiiPftQz5mWNuFlo/lxXcbPkLrTKbizzGkVPvMct7oPXeTL7
XdhCechi8jMsyki6rjSq4VpE3HhGdwd2z92kJs2raSoCOkn08F/m/NWgyZ6jVOCY
F6vKFswyeHTBIgD4FfFwZqIphmREwHOrDt5mBHxa5zbkMHIDuYR7IvCK1WtHtViN
8MPxaydl/QyiXRsB35/Vjfdb4SpEOROxtk7GR6XOANg41Mr3V2lu5G2Qob053/81
77WIb5fMNsctxpD0tCHPj9jASi9NnbYgdZxq4SMEd2ZPD/LAgpywX/H/Shahb8R8
GtDQqSzYX4nMbjF/pwONDqMyrXZdW3x+BXZ3MHnoSA1qH3SHekk+w0If4CYAP5a3
A6UBUALeas2KemkVDmjkuNopcxyNdleb+8aQ80kPY180wGuc5mWm5DHyKzzq9JK0
G6WW9G8bsutBvxdDPKPfneiGv0sN+ccA/TLPjKJ5OPSdxja1kYFfxRouAt5wjZKR
e8ptXKnzXgOg3cNbkKeePXExe7bmyys0osIpA45gxpSVS0LfvjbmElZ9qegA5YJo
LP4Ong0r9oHxbamDQcXfihDYAxvbcazuPrv8007Q1IvrBxObocd/hMvfQTO5ldny
G+PzPGgOt1IOy29GWr0uyEbjQHn5k+lH8hD6Q4Hhw/x+OXlxPCdyyf9YdTs+6OkO
5z9e6TQ192dgzL1y2QEvX+OgoEO+4E3Tp+6Km7gsmTIH9AENrghAzAyi17QXh4tI
mYbG3lsFHkb3Nyd0bffHxmJpNqskruyygjCJ4L6tfugbziR5hKkq1p2Eeuy7Zgf/
bvdewS/6Rg1wNZ+zV1yVzCSm/SAcuD0qFhzsIF1lHIS5IflsaC/Iwswj1q/C4jVC
OxaLw7HdD4ErVD0v5bCQMb7JojGtcgXq5UbGJnatQ479PtMSnp/Qfp/OlzNJ/VIt
qumudihN6XLq1g7fyVTl0utC60O7b8n7LrLSlzXcffaLNSMaWS2jJU2WAoK8futD
Z2ohklZvgDLG9znJfTNCWgn/pVCfcLhBV1vgbckgVvEHA+cMT4dWc32y6Jb6o/w1
P6tHtnb2P7hYKfaQqGN/jU4ScYDE1OmIf7xmzbsQnOp41grNQJqwPo3Zq93bvQVa
eha68b0Y2n7EleL9cE8gI5DJBCU9Nmos8rKYJPhEqUUHzx72GuuFvXBXv7LxrpnM
3WJa/qQP5pKHND/mVCWkjMhD0YeacJQPYylVa73QiiMVERwwQsLJWWu1zeyazgWS
RDbSQxuXfti3JTZ+YNuJ0U2GRhm/oA0fyy5wbqhGEn/ybMR60Bk7+ohRAL9aQCl+
V/kDHV5jMu2eIKlGtm5tB4N0NeuAMRMLJivsn9GpwPWqWcurIOHi41wHSy5idbuo
Fy1HXkhJApWAXHktQdK6YhuWKvMotCHCqqssOGnTswCpOmabtsn4XuXy+FL+lvk5
0wHBsMofX6EWNirA6u96p0i8wuXPqZJTpFT6ZyhxpUqdPowB3/wXd0rw8/Kdsj0i
hxVUVtWxG3PjCwFF/489EyDt4fxnSAbwZ849uSaX0nYcnm/nPRKIZUCfweBCEXrM
Olt8bUwEZuMfhy+HklkvZgtkR9OgrJfbaW3g3CUXMmrxoRKPtLVF/q3pZ8BBY1mK
JNNMZTevtWpD+Gf2EfqMl5NMuJcR9lvePy2nYXiF9+V0HE7tgPYQEQAJzQogmb8Z
usKlBVYisaZpr6sLkSi3uyJMrsVdV62sYEM7dnkPaOLkqNr3riEvaXvW15mGPN8F
SbNKwywxEG8KOXCUjjYhgjebKhONHkzCzL9KyLkPWLqaQNkz5V1xo7YZACi99Sf8
2aohlzndX04O8wrzKqOLGSET9p/WjgU3DslJBp3skXsFLTwbepBulU7S9zhl+s90
mjJWUpjKxKi78NBK2tZeo+ThTtk+2QOyycUC9nXpZfKKXMD4p64aDYIfar+k6odR
IRnJAzq/HOIPmFTjgZG8N8NgFJNEbYQ81EuQk7TIf26VEukZxzFkrr5a6V840BqP
leJy+didfYwSG8XjCXvbFAev+tf+tdPW4w7dN/rFfhEH1t9zIj9DceRxlHC9QqHh
QF7piDhAP9q7wd4wAjMx48nFaPrZi1unzB3GzEBljYMEVTBh8z8JH8b1NtkHcrL1
ZaO6X2S8+GUsPcb+BHUzzSwQ6quZyrEM3aKcLeNGj78CX0F2yuRS/KwUzHaxzwKP
hmp4smczBS8F5ybKaqLOZnsdCfbEhhnS9PqzK1J9xFe3VnTNiy1WqXW6zU0bHaGF
eWxyGg372qLjwF97RiDThWYnygD0NqURFtsBLY4F3A9lXhf9VVQLFOPQjo3A+wmG
Cbwbtx39zh8wpS+31g6ZBLAPm2D/rqrgoMoJKhH6TantNcqYTuMZDDdWZhuVoBn2
e2qHFz7lEbm4PGQ5vL10gc96YAElhC7dG8OvM7tm7eVSwKive9noC4iv5ozD1rxl
0pK9MBZye3GXFmCawpBLBW1ZSm9AGxLj/m7oG4Ngdzq1tpprrHAuQ8A/It4A0upl
SwzAkqm6m6swTqMx2ukR5vF9yPlnaUiw7JVJgbnk4tRhSdf/L3til6/H4jdmCQJR
IRnBId+QD1QV8NgUJQkvRftzpYzpcujRqZkZUxFKIPlAMi+Z+yp24lWkgBppZg1l
+I25blZNAFUZJkkS8KGYrNhC0VEE8o6R7Ufu6my1dLoUAK30I4ZE1zPd3GIFjmAe
LGYzUSknui46fUjrlewPRD6s+i0+mz1aO35dfWSGBCIm/DxYLAmzzj7OCCQOk7rt
7mTvRmwRUOTjjQ9jKHcAE2ks3rNorgyma5ebwcUGFQHgWrZ5mbUGgbLwHQDK3hyq
krHWnYENvJCEZGpuiVei6XXDRt9qO8zyQRSD470iUDXAa46areShXEbyDDug1rgu
MbC73ZolIdc+1wZh3Gf5HaSJ8053ND0bFIN3XTePceysiZxsbmhmKXf+DxLvRli9
r7MZ0xsmnBj5QQp5anm1SP0fkcnIbZbSMvC8zlYmIE3fSjeKlJmrIURK9if/X1o8
c7jpzuDA3YbSuYRaeSq9NmxNgCOElpYN8vG75ATKzPWnGY3rW6iMtbV5tOsIJ8hq
uUHBKJ+P1yadFniDQ5RHspyH/ngBzTc8YI2NfA+kP5WP+yeqnXSzo8ONIrW7ssHW
G71ZVvEjBmytZvID7pZMwX+HBRfjEpE7/smYFi6eqO0bGWyUt7GqH2tLlJ/LldM7
vy0sEGoeslDi2Qa9n/VfVz4zwV5cNyxsHbJ9d+36zQwzfPWcglL7Ik0vChg4iZk3
I4OpL+6B+QFICVELcomSPpKmi42sSWWoXIcBLCpELhgOnid8bLudKJW0kS3q+dGM
KjQuF/auKOsyNpQMn/q8cKisOjigDXYt5qXAG6isdlIJu1gj4dUbKhtPt5aWnuFd
LtIzdHTedFyjSA2VuiotFl1CgDJhP3zaVfaEWGjIJSdk3E1XXQF/gJzR1vPLoZYs
/jKbIbGl8Jvu0EBOlNfmvk/wd7cVp/IYaTJRcQitKuZW15D6W5lMAf0DQv3jfKT9
Y1tOEFMnJuorJUT4pWQpDJVeSYG/vO3u0G5xrQw4p6jdn7xnvD/Qiv12OTNcBWLj
hGYx2Vvi42oL1DqQGE1GHSVshqhDzj3Gy9ZFmxJ46I7Ko7aLoZg/ikeuvIW53+38
T78byMquhfFSFWZpT/M6VwOw4Ze8Et9ETKbrZjDvXVZTiX6J3Uq1Zcixyqr8kKV8
KIc9Qss244KMjRWfDeEw0OghNrzz5TBKGbGantSlv87cKjf3scTpEHj4Y0T+OK7k
mVhkUl80UY18XdshqdX7ao6iaNJbqD9j2LwysclTByQUOAphL/4py/ZqmQv7J8DW
IwAPfgHRgPRc+RUFWKZ5/ptf+gBXO3DybnCgTIeFvfXT4QnqUQqRtZHgUFglCZgz
LaS4ruZRkQLlkgDRNqt8/dimnpr7j7t9K7cpLoJZU2XkRRfII0AbRSQwZ41iKyJ+
3mFmdpPqxXIjjpE0j04z0j7sUbno5MuA0rEd7yTnooqaMNm/HeKg+18rpo6bXpQi
3EfbQZtR2l9uWzEraqm4y+M0KX+j47RfH0HYf4eNzoVVLJQ/gGUV+W2TqHxHswg/
AS7uKbFNmb3E1FaWq79mLfAOa3YAXozGNDN1ObIEcLVVLiNqHlbXKuHCw1nTGk+g
5QDfQwEparH5vbnvO4GHOUGFZLgjbjHM++N4pEI614bBm7xddM5l4KemOlt/YYAn
yIOHvHrzIGkvxiRTAlJZ+pB1Gkhz1aPcKk/BZGJNJiYyCZ1YIqxZloEb8ZNKFEVA
OTwHGrY5ikS8o+7eV4NHLNXMz2HJjJ/K3VbOZGyZ0zT3n25OgyZGFoPaplO6gbT9
CvM2rSxsZSxbZ2WjDU+v/boSTNISDy5gFx8H67OhRJ+zbvQyV6l2WUZXCNHKxor3
vXGOBRCeThC5+XDHhQlFOq7cVdiKWxOftLH8gl3/5isdP+rtO3OHhNCoWvNkJ9FH
SV84f8qIXxedMijRbe/cJgAG2DWgoeLJWrqJLAj1N8HXjuBuRSYKlJt0j92X2klH
5iBFx6kTyNd2VLyAonZlUWMfTzdP3GniLIDjgOjWajhduzC2l/ypUSKhvQe0HvtC
6W3An02yiDrLDsy14YR7W+FXcgyDApWOlFU0L2nKqnR7i5d8kqUkVrkRGbhdemau
9ggLbvslChvnaF6XV+ako0vO4nALa0QH+a8cIkZ9vJJaIdVU5TzS0+nfPt2nG3FW
ueVW79G1R23yPnZtsxZ29DFrx4eOJOWTR4nSXLsd3NAlrrPzqbT1N0SGLgm1Hksd
Sdu4WO4UxYa88rLZgK0Kv36XlRiN8DJ/Y4LVDFZAaVB5n+oor7UdrcsjM2zWnZRA
g3T59Z5r7UZUXGmgwivpMH6XlkqZyoNYB0RHjp1CQn6OKYqJ50+bopI+Wg7S93UN
suLZdNTEIaTOQdyEwmUvxB5+hPrCLYYuUulga8r2qFy9YclDtiZ0f8Fp8KW3Kr8K
7T01IwOuVZS64TPA33lioA3DYw1EH1gJKmSTeqU7HH+Tp63v0eDBFCdIscVVmyRY
vTmzl9PA2ZTaM4KdJR5ijRogxeQCoWZvj9I84kL3KIOGu3gBEuTpp43ttdz1Wumc
XQAF6G3rRIJMSs1zZwfNHqdPLtqj935OEx363EjQ1Ls0epP8s1ywvr0hC+Ps+n0e
6e7Ni5sAl8kI2fjRM0cBzkcHlr+l3lG4ur1yFabZZyFYeG4zdVryNr5NDWvsBenW
wahLJKNrR93MdWHCy6leCDG3m9501/fraQ4JvsxDOL615NvcOkPqGZgVxiPLr0jL
e1aeFk7d+/WBKVhgK6rdB289m9kEmy/IsX3zzkPPcp+koMPi2zzhMDSKoZ9j19lf
k9ikoUcsNZHLnHJLy2sxcg9okZc6F0gDT/NUn2iZFE25E+B1TkCgvR4c58JrypBM
6Uhm8qD5Aw45zYPGP/xeOEUbuur1OCqReed/eKedNWelMCfkbQidNMZJAs4MLDy2
KYktcjAdIThSlQaFZG5Nj1+3dVVdaHp3a66XeDAV6ceYmvbELVL7v9L0XRSqTktR
rwky1ZTNWAaemFiOkXRxkotTPFI/zee5d1VcIKDqLzjkDq3zYiokACAT+5NjbLZ3
B+kPXph5G3N3uPtAYln9NhA53FcoUQyBsZJeBKrv5qHQWhOPq5EPXTXAX0Dz31uO
RF1EufTU51f7Iy1QW0KnWXNg9329tqoWDlWnp+Pwx4onV6kDii3Mjzqh2xHpVI8O
uIGVPfKZzMrmFjX/RBmVb7qG2UeNQ7lqoeIC+JE03FaFy2HDqXyt670twRriIJqm
VMyN0UikPJkCIplMAvyPxdodwn0Tp/hWRw5t0u/5/42cKw3bdf+dO+T60lyvCD7Y
6K2IzNhk0anStBJS7Ws1TyI/FuAJNXFmFa5v+5M6E3Szc0fbfIrzYmMeV53eLCgi
T9yTfFaKbK8W4OOAPd7p67Ce3+/GqQSzmMovE8FXXLDg682ugp9YVg6W4QXTZ5va
Vu2BSxUhmyB7fbdPxTOpC88wwSc8Pu9Gln/TXwGYWFu7qqjeU1JQVPV0IRPp9Ihx
LZ39ZleuHzwfQgzBmvxVKQriwq35d9kGCAUGlnTQm2hYLVYyPbDvOoHhJgo05MpY
oOLAyOcV9LVWJNEtid2DhWsb7KytLlEUbzifhRdKj4Dr4SJCBkPVXojOoXopboNe
MvCIeCNwcHh/U5Yqoc6jlkt0AwkccdKBo+vUfoZy2GxgZbuhlG4/JXmZGbrFxzfz
q9PgW12qyFfcb2BAEFJdiHDS0nSnv32A/Jk9qgJwDrDunHPNhGeY1/kWhH33Cm/D
NkFK5o610db4IWQfmT7jzzMH+tdiFw5VqHBKRqbqqQmxhFy5BttDEQEPzYQXAAGJ
cMR+GhkfHD/xR3A0G+DUkAyUfADmvi+QvIQyeYzIhN1J42AbBMkLudbeBlXyf3ZO
wbGzqVt0MjyWvlKvLJYQFFesimZuFuaHaJSt4l9v939VgeNNj4kMv0dHlxvPT5HJ
6GIkCCWMW2s7B/b9fjTVBQXOfN5KMyKHK+knRT/vdXq2fJRH2UuDqTGDmd+150lM
UP8dFMvvk00NebHs94oAUux+pUn+eOdar2R0Wy0K99OtI2/iLguHMV3+nvBM91xZ
fvsDmK1KhZr1v5wytZoMbDuMothYYDrhahqLTp3J7Njhl0iGKm10hpi6zUrrbJgq
px7/6B/X5xdF8Pg9UNtoJBQCWQrUM4tnJhTfiYqFFqdZpNndq3QTwxznSj48dE/E
FYVce/AAEQm5i28oFib96IKPTGIh//QnGrNdAg0VUuIvyXfeScQ/5NeFz9ZUAkcF
oyvafM1KIvZN+fd2Jnjn1cyqTNBwQbehCAOpnpxylGgGmONPyzkolKI3TTtPFU7I
PDSg5nN8dq1Btq1vDFIFBH8IbUunHJ991bNkRxozzVI+9wRgS9zih5mcBPut01Lo
LwwCp8pLmKHoRQDfBJqoK7FaHrx/C3NwpVQu8o8i2m8OOnv8eWa7ruOfd+I6ZvE1
H7RJmLsWEZE40iGw7x6GdSRPmjejS23tjVGeC0xrTTFYr9x83WTZ7gLCfhxtdmwj
0OS2D3iBzq/wxaNi8qDrF63BCWKGy0jJ6KT8CMF3iE0Qcdk4VlNrlrzr+eQ4E1W6
YLiNtS40+McdOC/pWrOiFegHqScLeymIGjKs/Mnfx4Ak1DJcODalcSPtQXdWm9WX
VDozFOmGbENJkisXPlrM5tiBm5YKYSzTjsMmX1376fVy+XvsJYgeFXMxH23LLYOQ
By3NPIXWIgVleyBXpoCeZnTWyBRoypc1L+fdnHwAn5yNDvbLzb0uEmWKrNjHc50z
AjT7/OGz1oiM/aSr4MOccPW5dB/aBx10thP49REDA3B/gM+ljDYuKQVpSIID1OjR
BVcWGIbquohQ6zXKrhzx17sIGwaShcJ3RpKL31kyik5pk81TPu3ernPA7SgMUYRp
zwho5CY6vUNTV7HAggbDvpyOh7UXpusWhBRV8w8BHJkboker/Lhf2A0/ysM3U7/z
jDZZ2Dsu0UTSsgcA5panYa6YqCqLUQO4YJ+RyY12yTFPbnu7zBZW81FYBF9Xobp/
shZyPV6A1FEkNJzgN9X5Khe12sAmTQPHwa1rxzyyvcu4kQIS/IYHGc8PkG2SwzYE
eu4H7+qYPc3WpxJOIq8zPRXzmE+Dx3D5n/5Y4IMX0XodiSq99mHhkyoRwn0ZtvVd
gzV3Cb0M/KitxBLxe5aiRoaFCmpnYCJHpEMGTPKUx+p7g7SiZaAdGuPo/b1Tm+lX
glr0R4gdduFOTsHaWJoCHFcVkrdsiqoUy6enoBi2IQCPZdAEoE+az+KDrA0VBr7Q
RNONZow30nEYkr6IghTjRmfX8SgMcRbb7ACFMUzR1IFI/wvEEYAxbRE4WHOqvNbT
bWWJGA8ASKg83enverHU/HRN73JDLiXbCRkQEY/yMP7OYntXGe9zJ3+GJ2dfPdaa
5JvaJF8SRJnAfz5pX8MJmRJS48KeHCpEmRjGjfLXT9Kx3mfA09BlHJ3SadWkyjC7
/m+P8eS5htdFVEbqjRaO8xoo7fiYOU+5GmzKtL8Ha82OUgwM/LxPEKD7tSypEJII
PyUb7TRc7lpBbtLV9w2yKsEC7A3xRw004B3/U/JJKXHLdXZ4ljyq/LeLMJcvcWNI
zrbd+W1JfwkK4FN5XO+wl34OJHUImKxW/6TIO0LMeXsmbcc5QQMfEUeZzfiT35Dl
bRwLR8QZts/La7Y3gKNlVD2V+1ac97KOKa9DB1ZG1yovyNY9bPDBChSTCfMQbNqF
vU16/eLh837M0v7GEn9PloD75SXZc6aCUrChlekHvUYq03Zv+NhNeVu1b6U8nCfb
YEyF9lqYkArmJpjx+z5s63qjnyoC50W3uVEiB2nUX1vAWxI90GIRT37LxBgr9uzq
HDjtpFUhHaivV0Z9Afpqx7h4KldjOor06zbQqHd9jAUbiVqbjB3NZYlJWqxZN4n+
joYzKQ90uGvseLgw0MLgsJpcCpUOJf8EijzkfFyq+zw04pP/EEnxVojTMgAOqo1h
aPzfJJoK8yUffsMsFm/SL/5Yy1bhyo0Y6/0e7fV81DfLURZRWL/hsDsmhI1YVj9p
Rlh4iNVTx059FZROjf4R0i3j2b+qcRif29cdKyTitul+DhdB4/BTKGbJ9KfWR++Q
b+pXl6QOBTXqMlQ0qPvYh1MbuimDTKQrSPGKSoCCwrZK1qD9Nq7sx8scUnrKR3VP
6/Gh0cbOl/TTQXfoyiLzWk7F1/eDl+HMXWYRKFBJYNGeHtDuOmBw0lTLyR7aIqZ8
HcGD5ud8dAscxDryt44zlIaEL69M895b5J8r2kIyY0fGWwfbjsumeFb/0gpseAlk
pEfZMfvdimFmCDdzlO1aWcSCL600ZTelZkXknIC9aFJcy2mqzcX6MBYIz4UCuvtM
I6kQjvkbMlLFUxdd83ehfixsNoySYJSqzxCjBBcZ1d0FRevLBBfQml/H+b4qDUd7
IaOzktYJDzleG9sd0fN56m1NUvaeOeNJOdvtIzeW96O70rqAcRI4pOLhLBXSUd3C
QHIOox2aqXSAYEll8O7cHoh51ni2n2Zu9Yp8K4oKO3aLn/mDbFmmrh0A8+1QYdW1
5oMagwCvZ/BQZqQ0BpBYOSyakvh5iEcoU9/61SYHyqQZmzG5TFG9+5Bm4uRlbmvw
gKhCk6FQCVJRjrd+ghTWk469I9fS3dileel8dVxdSAz3SdWnMh9TZVefUb00oX+T
K/9NViI/c3coa6prBj9ynKKLoDKr8Mhzv0l9pp0J3fMAvxL7BOmwYjhLJ74eylp+
h+5P4tC4lG9UWziYaPoHjjUUvxA7R0NU2xfhiVpqo0o3ZgOirCIRWLin0znCpiP4
owuHe3bF7S6K50W0g+yhBCn0dtlfhFUmAdq2RsUigtXcD6QY2kc2y2wBvBt0WZTQ
NTnXIHqqApBzW4SRC+rr5oeO/+rNAt9mMZOVHPvF8gLYXETAvqN+1oGfcoSawJPN
PW4UbOxuWRw6Tg4OW3SypHY9Jfj/MihNKXE01pR2PENP2iFTZz1DqMzFWYa8b5gu
KTQZNIZcWX55v7q1W67hay/8Fi+p6vsEni/OCHyXvSc8ildk84aoy+roIDHAvBG7
N7HqkDvMfGSDey9/yVdyHdf9OKXbOfGsPJQvbYHAKTU7g8lkNa2QndsV16pGhmXj
eqZuZ1qVs7bAOTmh3IFc4N1/51kXpGpLizWXQEHjqy2aF99Aa8vwzTwl8Z1mgewJ
ZVyYOz1mMrMFEppokjEpLnH+qG759YCLfYaGXVIn8yWDMIYzVyW8TJWj9bJk5RPb
rYaAblfdSdSOSZGuoUPXSgWYgnC2dlS25yOQh9CZxcn/iUapKe8lHq7FqwQj4nGL
+NnSIyxxvHruBUqALOV5a3W6KUSumWnVnBPWbmbUxxyFSjCTRJVeOHsI+Ov65EDA
oF47vYuebOJcLMAnnQ67PUzHghRes7CgUbxpFJcOMU3ocM2RWoKnzlpwrHDIzmWO
pnc0ljo4Ob1zylKnphMo0k6qVrcOaxxdtYEpqVho2g4k7jpFlJnd8V0f5fngjGPi
sFNI7qV4GT2qxQcM/5rlYl9bFq4OWWq1gxEX8lsuREQ7df6sNadQikH9F0KQHskm
muejgm9Ryt2sqYolhRp53HD9U6WcbkTVbbMYY/iYjIQocs9osvD0ABFvsQq5Gwqs
T0QBlY0oB/e8ealgW59MqWZT6+4gMQhxVNPPfjMvDRTEemHsLUVK//9pE8vLIB6S
pmsXS+bUSu49GD2o/o4opIwV0JPZVxQnvMYE9ULSWjxZ0LLfJz/GjUlUrnpSxnLA
R1fELlnzxTUyeCOLD0ywvWws8TMjdS8LMEpDZFVFW1tMi4Ukd0TExpcTO/3Yyh8K
Z2qP6liXzjAMUBvTTMAEo1W1Y3qx2U9GdBzb/qLtVR0TiZJ9mYQTt7jjKQZfIJF8
AdiHDG5gf9BNs2u93+W5iBVWsk0HmgKIvK9R8zKXUftihafbVjBQYoMAdfaJQc4K
NQLYSwyPBmhrQHNca663+tUya/4qIm9Fr/+PduEkWR9mYBY/yFzePX5KPpFcIyHs
Vu2IGLD1unJc8mPv/xN5y3dhwnfqDQyndKmebx2liu7aokod+go2c1L+cO6TEz3u
cHTTMwjFmmsbylwO5s6mrljPy8YRqfDcOMxJCC4ANNq629It4SUdVIRC58ckw0is
VFGlIjCD5J/F8X4zA86AswD80xKWWvU9PHzFsbSpHYhz94vW4dXv4AZmfZ/rJ0fn
qWzA2k2dIejmo55t7ZTNcmvAqLTjp3SKuYpr1bKE7QUeg78Ko93z6UTHeGEMutTJ
X6LY3tWRMre19J2FKdH/o34KYfwBZzO4wvj1eaJnjA78UAtBiJFUwkObPp7XDK6Q
T6OPZ9tk7gnrfyXgxJxOCTJPXMirdbxAdaff284GR8L5azzh/zMvhXrYoT6Szabx
2o9F134tPoU/PFAxfDbOTbwt+mM1jcVBZjIBIuDbC/MQomUC61+kAvhR879oBzVr
RhmgspwsXjFChFLrjtzNtvWF5uxDI8EdwKgsZ2VvZr1MgmpRuZ+4xf3eagQ4Ix+C
SLmhRM9H0HCCZ18gPW8o2i2i0OO9BZEVQfH3h7xh8un4Gh081ES5isfxVUyHhq65
Ne6XvYyl7boVs2vSE1BVNlQ9R7DAX7pntuiioBlFc31h5S2fbZSZV0le/q5jY95y
GwL/Ne2psqrQK4gaifDJwNqOL5lKpNpjCmQAKajLi8n7U5uCvwNuUmcjiyRO8xqy
hB/kT9giMdR49CgcL5Uow06gkQaB1Zr5FBO1c4OPAaJg3Z3Hn0Jsa5dfY5q6ay9T
zyDEAYd+Zz9hDU3hhbZBtV7KzhB11MoKTRiQ+N+8NCcjik8tKcDGaYip+f+AkHzs
cCAgtK5NOBvYil4r/F6cF0Q5E0ihg8iJAgIIs9w3BUtKTphUjGA999UGAGylxiZS
l8trPN7QhwfKDq5P4J7xv4q2Y9Rq8bS5neyOJSHcq6nNyxcTc4DHWAacuJ/vB+mp
ciUfqI+ii2AXM/6slDvMsVrU72WgXoLN1jrNGbP8Ux6PG/du+Thop38d0Eet0Ath
BTGzlgX1WXQaxXX3ioLtEeCiNeR9knhgspT0vOQ38QNtdjsZDIXuD6mOL76qb1+/
dmdJm6/NSy+2652mVLkIpEmb80JyGc88ru7JhgfptSYJlCVgo3iHLQSec8I4EaeI
a/iB/AknCwYp6DSmOOV/lroN/Ms1nw9au1aeo3I/poArdyjWMiu2sTM2Tg+0f6MG
g/N//ulmowghMo+OTOFcLBkUwj+HaojQ3/u+nF21PCykdGDsBJTbDBgT2B3r+Is7
ArNzl7shkknAg5kHkQmVIe4apaG5N54CoBXCkfKoJzus5aV07UwA/2PrGAbnW7Rc
SJx8g6cu8PgtJU/QRmSKFlz074rO2BJ5lgyxOR6RZFpVU4SlXj7qxiS+uT7KPut0
NvxQDwgEsLT4RW4XhmNhMFpTC+GAXzUqqXB8Sakt942GnD8UP1NKY39HurMirjzY
G1ukLGT+dQZkisTMpS5FLOm1fxSNkSMCrVsxHVhVxx4=
`protect END_PROTECTED
