`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q6wQxC4U2R0VWfjoec0g887iqOtvwcC10voUzhguShWeJcR7umS41ZCREtuoaudG
a2q1d8ly0rCX3dFtV8Oike+/DP+7OYHUqSHae+BV8DOsAaSS/lq83ZZLJF0GE7pm
0kZDMD0foPax/JdY1Tjag4CVPBfjg6fYBTrNZ6xf1TY6fI5Xqs6FsPDQ5AMWCMCN
9XIEOigSbCBuu7Yrgd1s0mky8TLLiPnEzl2XWpyDQXFazsbTKwu7quH1YtFHxP61
eAWbV44zob5Yoaa2lGKNh0gDTRsf0608iwnpfYTqb4YwDyuOtx3CJJjXoIqT6NCy
gFkgeXKW0HGU7fFTef4U1lRgDBtU7cjges+A+7Z2rra/3wCaSsYds5VqSNC/luIS
pEtp0+3XUUduMhBkhbEcTufjSXv/MzHZi3LBtiiMsPC3oZ+M0KbxHgY+Gg/hQ3gZ
gRkxJw+EbtF/ikas3os+HwAZWqzh2SFRYg9TBkvCmx/Az9zRje2w+SOOIvFmLPC3
Sm8gcEmdeJEVVmwuR2WWF0Z+ufiThfzQ2tYU8TffgT3NPCqA1InMpJxFNj1l1V+i
sRd96wuVPNOHr2NNb1+dwZX8M9aIzETNVIC6Rb8/fqA7mcbQskm04311Wr7bXFqk
r4+EDKM+uA2UlwQihxqyDZzJuMcNxV96L8b5bA9Po4L7oW0z0JxHFE04nz6eEmNC
JEtCMhH4uwt580lZM5tHslcVJaAabYRD7W7UJwMn6s63wZsCU+tLJ5TXiH1IdnM6
L8khVG80VNyoKahMcJQlPKvJ0KZ8mSuBNxbl+wGjcEcGnOqlcJRLTLzFxiXQ3vJO
es8Tr9fDTi11sI/BeHMAxjEVu8CHojgG05tO48HNAIOPLTB9DJ8snyDjijvALCpZ
8FiRqbdAD8ofWNc3/m1b3V4LxW/4D0N2ZGisCC559ff2Tdlt9VIdTiaksAfLKbzs
cXWvhVTsJWEZ1MMLHP13am7fJdzgr3E5sE/DIwuIOyXg9gG0A77kHNcwZiD7cVZ0
pZoLyiVuT7ESPdKLA3FngRTk7P4IqZFb9/loUx7kGdI=
`protect END_PROTECTED
