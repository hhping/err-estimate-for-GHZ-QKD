`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/y4mkKsr1LRbfAe0w6Qo1csunR76joVqYQ0Kt5JlEWOCDkgUKYIUi7CtTjsOHKpc
qIt4v6qLyZ87tmtNPyZ/willPABLKKWE4brmBXFP5YscmpJn1CS6S1GadFUOsU21
Y0UnnzI1iz0pVg5aA2a5O1wQvFeNyHqN1pbY5SFE3eRt7t5czxre3B1FT4Rb+5bY
aRAR2CQ4E/op4C4oK1ia3RnsHvOGPTiLuDHxyY3XrhOmrPUXeISrLXCxw5s4EbWR
vSeiBVIqf37WchTFHIccFxt4sg8QtWSXRqFgzR2HvfM3Tzhcb5xhJIBfjxvZ/H7z
HGYbWYzMtTV/WGDVaOHmhhJSFavi3pwF6775bpJlOGGiZghW2bzNrPFmJzTB24Rd
e+3TFM8k2k9PId5byt3Hcuaf10c8bBb+r4ZzvwKT9IXd9dQF+kUNvO4wQavUv7+C
UZ6IeNahH+TuHMJMtdGIOy/yMO+CqtiaP2mtK1vSwxXSym3eDgRQSo+P9SI+Tujw
ACvIuHIhbh0sQ57CrOQ2dCvb1P3R0CKPbtKETVThE6tBKDrAlF77Zor1CV/f5kRH
moJs5pqvFPfZSmkcHaa/CvQxRBrI8MKa5GzmVSugSplvyQzagEplXtvlqQZA3Seu
8+I3otBxpM5U8PdxheOrFh+yTOOpersoNySWcuLlcRW22ALJIXKKY1g9LSzmhwm9
EWd+CqDCd+/QFA5C7q7EPISHRcD1hVRYeAg6+t0mhOFpMCX5wtFo8bbIOIXOQk+/
Vk+F9qb9HbX7+jb67pVFUhrZim6BbSqmHxG7VaDpTzQgJVtPvUlpmwdHzfH+E2Qg
3XHycc5MaZsA+2w1ICcwFPpCAoeni+SZ7Q3queOdZXrPGZh7DrwDOuCHo7i/gslQ
IVhP0DbcrudpymdVt6Kv9h1veosz8v0xTlfhnSsSOBU/3hO9UJrL4Ga2HpHwIAdL
85VV6GTHs64pGh/Op1YlcA5GUv14ZUsmnDmfDcm69mdaH0wwJAJF2OprAuvOqGM7
Pk1g7GgnwyCDu/mdUMdPe8Wr5Tsd1fA5d+MNAXcfN9ZdThxNvsGgNDtnEzJVUHJ+
oyO9SUKAfVMg2xv/UwT9kz/D/9e82l2qZt2kiQ8mYik+iuy5YioHL0X8O9MvNGhP
xnc7Bz/x6g23Gl3RWLoOzBxKPxChfaRItow2ihJr1+UrJk3vBNWWN5JEbGYeVwkV
joUCF1uWDy+Bbuhq2NBQ55+/0lpdm5xuPMpgEvsYR/9IkeD1HMr7t+1aGTlesPlA
kZy53Aslh1xFs7d3izXDpcC6oL8RQXpiqD0bPABSWPdnjQ5Hh1XlZLYbTPj+V3rq
Z9EeoVudMVRKPyCj7uR1Qutmx1MuEF+ixugNyBn/QSMjaM5F++Q4Arxcpz/d7xuT
sAUxcDpdkY/98W1X5bS8tHbW3HC8WPG1tM8dZz9GgUM100iQbCxaPtOtq7wIIly9
yXRFXjEASv7SeyrhSycJ99x0j/zXjEKAeeYj3T4E1a+3MCPYVL6/3AxaXj+ZHmc1
qQntj47dmitV+oSOWPNs5xKxEUIpTxFYqUFuqjwVLrreydj0vSXUqxr8orLZK8uX
SoibfvbB+YcJShV9QT/BBkuiosdUjXCqWaULRsKiUmgVdzanekYDH0l5xzRcoQAq
ktzCYfcoXtETcBn0F/Fz902OA53PJSMwiGVTijWGA0s=
`protect END_PROTECTED
