`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yZbdbT6Qa4uYQqaOgxPqnwSz68k9slbK0VQp+uIag4GUDz9140JM+aufoe9Qb0gI
HzI2d3evFDk66+1k73PfH1biwZP4OAZk/8u3tQdfz/ikrWfPRHCncFm2YqIA04QI
B5iCdJqHdGAD631CHms1P689S/BjCEAC4SvGJsYNFl1C85PDjbgk0M5MaKF3Cl9O
CQ+my68MvNYLPK4roLiUKoc1OJd55Y4IBg+e5VXsOQpKzO9nkgrF/fNK4p0uLJVM
7ezIp0VuFSwj/ks9Kp0/bKDPsIR5FkT26Gb4B293QiKrjb03EGia8ZkVz3S8KTSe
5infq6Z8CiSf8mPG11qowflKB6oWGcdh4hC37wU/iCemaAwRhJ4wlZ+Ehetg9dKA
91k1Rc08NEuO85HwgEvxUQEsACEj6D9L4wmamqiVEe/vfVRH9oPRqZ7043BQnwHw
FF5O+mMnujolZbtnqDLH1mREfPlGGnXLGAM9z17MrFw3fAtZx2IfyCWtvLi64x92
H+MHBcw8KQ89j7IJy/5L9ns9yUhctiQoexIJUjCvWoDsycBeDL3CzV0BNQhFp8eO
wJycK1P7mUYjHB1MMJ7PTOGNvSzGQG5p/9/w1lOvRzHLUrilvB5mYAdpEtSkx1qq
0LT9hhDmR+giVTdO1cwKtZ7dgGrVJUiAA8MkL3tghNsi/966Ztq3OqlpuxLokYS/
hBUQcvyFgpjamrlW2r4Y1FvYlKhjjzokoIcZjzOEC1Ahjsx9f1B9i1IapbliUKlE
bo8Qq0arupi9pJzg5AjxtHvef/930blgMx958Q0EY/NGZlA1kBLfibfWQfdI19vV
Z34SjVihYdL7xKYsn9eG+KKeZGW97abyUW59WgsCtPgYXRahKC0tDyqmmK6TT1KU
9CGlO7KMCwPCdgQgTRWv2OLnWCxJPZP6i080T0XthVst9OLYnon2NXVwTYPcyWBZ
h/px4x4LfIRnQeHqBjX+5OctECQrxsAYkiErrsE4jVvuDoF/cz0Kdc+oi+USXrmu
NaOXH3p+OndDgUdYrlcxb3Pee7o1v3bhSe52Rl7JbO56Yt2uYDli1e2P7W2vYxi0
4m4gsv8/zkiCb2uaOYu9x3YpuxXVnEJjudfTIdDljNyNlulTcszDSj30RGcs6MW2
052ZORaybvftJ6++PstfuyALUZtOaLOoqf2+E3ycRtEnxO8E86ZIYRrn2rwVQpBE
TdFC7/pm4z5ePh7diwQwAeLSJy/4/5X8+2gQQr1ifnDlGaQyO7TobCRmpiQe9reC
Ld/fCNiM3YSwcmYFf/s5KxIyQJcr+ekHHL+4xT7WQ3nyuTU9I1qPgrIzfLyJ8R+A
pB3JNKfPxVOVw9wrfQuPPayLPsE0VVK1QIcDIEHl6ywMGgm7WDZnvH3r/ZeFngJZ
U0YFAZ8fL8JD4qXTXANMlfY7QT/YLL1d3HnuJyYBb6TNfsRg1bvv3B2f8ACBklRs
hni2DT9coX+y2PBqlrwd5wCKwgk1AzCYnVZOU5G9okiN1Xr1rgWS34imh4/dgtvt
vj4N/L1f94iOttfQRq+jlOfTcMSRSboVGE5xL71uDEkOUprgXePlHWutTvLIB0tB
Hp5xvxiHLo3QQHsHCV4FlF15JMHU4SYKLMoYJThOcp3kafjbTKmAlKxHNq+tVpFh
vmnAT/caXK1QnOcF31bc5q1Uvbk8KJbv7JMKSGhdljU7PVMhGtkcCrjJvvC1WOpq
NaSX9DEbg1dqlQXS1cfmmzWpja5s8q5k2eUHTWGqNTLYmxkmmglPHPf20M+gA9/Q
aWuX1nH7X9G8c7vUOgRhSclWjh0Feblzx28VYMC+Ct7UeRd8zHrD6FL9MnkzlDji
s/1HM14t4B704dYJsshUx86YDLVL2hJi1OJ6hQNLLxr58TtKCcDtMyHvC8+kdMjg
MryYg43AS7Bg7hdNnIEiqKXuAryhIhB3gTJuBS8DHxTSBPuGV94RJ1GlBbOk7PZH
iqlrXAIwkzfOItXqOEaUWqb+42woMiSsd5H3BaDYhev0x9fSaKOzYiH9ICpZzYD4
1H8EMTalOOI9IPFdgITW7NOJWH6C/Nhdiq/0ZYqEYLy4YP2BvzmCKdlmTInAB4cN
NuTMNOJUFPl6gI4pRo4zui+UMTMM15iTHdcgFONl47qkibiaxcWHz1Xl4vW5FQlp
qKQ4GidpjnVMf+A3YFgTJHfgY5Dw4cDffFY4m/WDg5bI7GIiUosxftvRqzTEtwiP
vN+2gFe1Irm9hJG8ePGXSioBv/RbudDCw7Tkq3IkXakAD/syz4EWdyK1Wa/YEMcy
V8Nrp+tOmt5AYU0Q85zg28lfS7WvuDX1KGzfj8nf4UJ/gppipPTPRv5wq8m7aBfr
CI2vnVOexUb056gRz5vgyhN2SguJ5h/RrUjxRnFgzBxfuvZHgPGFBF2VrRBS1DNo
imN7iqSOXaKuGMC/V5B27GQTYZ0KnXdi8Q1eJ6n7amKznX/I+8neAd2cKs2pjqHj
YtCBgZMfDkIrH2EWwKmVakuORfDWirhWIsghgmGgbfkkZt3IVW0dd6h50N/uSIv+
xHHJcl1D5BsOLhe2AKpFrYr7HbKD95jy1Ad0ub5fMOAVRXo+Xe8FLm3XrssS2d7z
AeqUZpgY4C+OYYOPvOMRnF9ZjqonUhZrQk0E17a9/FyqKUyQt7vX7H1DeHs3dagZ
Qi/g10+ZU0XIXXE21b2YS5B1c48kNVUKA7UYE6dHUN/kRJavX9KXmqEp3XGiLVfx
iEpuurWto66bl8WOt3aVr0cAZ3RQXUvPfGCqhJqCUKVKQeFrddo8hgx+lvypEDZf
+6Ii2sQFJ++02OJ1ClsyDqf0+wPnrIAgKM5a1hiMsDck4eLwvsQo7/sQqaTNZbjo
hpqfr8LZZ140GPW6kDyZXHzMSyuwZOA1+ww9/0Lpf1CZeeaMooN0HfGesOHuUf1q
m/IsmpcKvqjxoxWr993AqH8H/8H+Nuz526yAzO0tCfTHSIdKLji7AAPSU/9gVp7U
ooIbC5NsufzpJ222E029LGnbqsBLoj60nDkfApOktxH6Q6tBNE7Kz1AfoqOMUafW
jpTDL/9SYDyW+CrmuFCssP7g/2HMpqHnmPyifJYKnVW3MHRo8gYKPKuIZmzuEwLE
77RCI+aYHQkEL9cSbUAbmzITPuAEOsPk87qzaP5S9OJ7eUj89gDFKp3AI3am1v/T
tDp6A1UWgrc7wq91mGCTqMFuTsuAs35KWe/F0X2jCuHcrhHC+SNGjoYynF8tzpkI
aGckxYHPZ5prVqZ/2Xrcf/dsVFCPKtkNHjKHjpoL4JooQoSn9G4FIJGXkIYuM3hn
KuPVcG4mSf0zP2m5fS9tL2bLO2KkCmVK8PJAxLpah+1RntYYN1zaOEXlzP8u8IVa
CVcwDuN7XB+tl5OWwIcxftYk1Ajjck60pG/UCALlA1hcey0cVJ3xd1nP0+slcJWr
+OcCwbmkU5UmK2f7elGClW4amDKcU+sywBCauGBAi4CUWopnNWOJqrcZIz4Ba1P/
XSgT+W3/RuYgRvF7uG9i7sWNtXFAw7mIgqrmTJN4GFrAzxIQrwrzUB7WrbYo8Z3S
kDbUkU+NbKFOAz1blLri4Tjnf4VixIglt7/gsvPqUpinwbHTWLpa9mrJo3eshZdS
46bKuv24WWE57xPd9jeCNTK4sH2Kj9WObiTkrG/zOjvLw+11HOf+HIC0o2YyTn6B
aCGFAnDIyNghAlnrgLZIZG6wyXnmaAocqelet0jv4u8r+0iy2mTHJ5lpwSClko1C
lpsbjhbpm3HZrCahRaXxKpzg4cGFKgDyd6xI1jxYnkI3heOuPQKpwgiN6LY9SSHG
4ckdssARiHokhaPov/BtgW8zjZPzWtqp6N8ZgEJNSLU07yMYo0X7xrjfcRUcxweq
VOrsjAmpe1tJh5zRAXjKicUhFFMz7UMhosqVwqdkj1O9Ap9Ks31Fp9wst1lXRWe7
etp87YUA3fX36/IofjN2T06fDnnOfXkWR1CrH6HOyKX0538Wzi+AVt7qcIgDK+AV
2MWv9KO/nRVYmndjxeDZL3p5Nay/tWiUYtKdFC235M+c+lHL10rDqMs5mErgjyos
dLthLlMnvB6kLHk7utwV1ihqxEs4Pwo4im1rackEOi4r9YfsNsAH/eYvG1mRXWAP
SZWDuH1LooiIHh5rhkadAwjhCWVra+JcLKIzFC7Iun5f03azXcSrWkz74WPv6yGS
DVYo4cbZK44Kdqp335A3wCctZGd0fawlcUWW7LSm3/HbPp2K3eTfZGelz2bxXHsg
3fkc9faGWfKk7ugZqeVUtDCYfWMm7k4i91YT1Jcsm1i2YsM1Tt7fuzSjAjBajOYn
`protect END_PROTECTED
