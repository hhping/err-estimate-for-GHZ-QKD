`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f7ZzXNuDy6JXXqPEemmRZ6tRD0Tx366pEAsWncq+OxPnf0q8YwSOqJ9HyFLhrY4I
0ka5BE6FNnIwPum6VXr4Zvo2RjUxQJE7+JAG1+EcNmrTVatda4PbpwR32s4zcVj5
kUyjDFO9EGhd8ZaNi4Cx1PXV4Glx7N6uv9K72CK0N39TcYgdM/9+yPHdbILAfyn7
ce7fS5DgHg1lVrZn2TgKfAVHriZAYFqolYvcLj7REOO4uadOIcjE6P1cQVbswAn/
ZG6f5dpo0BiltTcrw+n9xszVqadizH5b0vVXIVNlXn5z/8Onk/WR5XrVQGispcyG
q53TMDWAwGDy7I6vdpJutrRA4rfS7PnyD7VJ33GX7HrTvdb40MoGpnagShXgQeWm
IbutNydCXkGpaobzIm1KjECWBOaiLkId01yA8sFm365MXfHnwMVpoUHMY+pPJ3pP
j0SH676XqH+19FEqf4J5pUa05qPA+fQpxsTO6S79pmGBjPcdeCjQZLt9TLRJmFed
Bm8Sm1phNJlT3AXx7zspbcUmoEUSHvwjyQ5lDHcvRpYoWAv1xjKjX4OxsQoJ8tAG
Z7rtKSdt9l4Gm848SJ9CGIZRRs3KqNR1imN8gFQhmfX89auam4rOj0OWEm1oAQ0E
Bqd0WDyEN36wWpckVLMnwfOjlV3giStckVfn+UOK38+WBDQDoBBk7914nvmc7x6N
WbgNpvoG9xAi4bboUBh/BfvN0RQPCHzVfJD7J6M/+9p97rbIiClHBz32B23uk75L
0A6IMfny04EU+uMrzTevOYKwVpJbmivZANqcTDlvE+YUYx+Ae9XEnpX9q+5pJagK
Sb8I1qWjV9ILpH2XwWUYkgO0+IpS4HoNh9+wkmiGCmUPvfEUoXqNGQoM6APT+Rau
ecUdpoChhW+M1/mVw/uIgFqCZe8MvH8rui3aejof9MJk6O8m6fS/y/vSkXehXm78
5EezyA/N6Qm2ZbNoIkvB3ZTqq5Ds15uBfJB9irqF1o97kjTVEMuxlqzDEXhW7pn0
zbxsx5VWWi1xt1P3AlyWlCktfmyDLleyN7REwXh8jKOvOUKibbRCQbJVBKlT09D2
eeWZwY0duDO/TGbldzoAdVfeaHqEgR/TcxieyRzf7GVOKW63c2DaiWDeWIWcwn6u
Cb94tzY5rNQ4ma1DI2toTjpmn+Yge41fWK0q+q946tJNdR7LKHOmfI46MrkBGEwY
wT1OikgrcdMNjkDROpusyCAcYCWqyI0oAA+jjan8bstM+F4mBeRX8HBiYpBWwcli
tE/Rg+tmBrlDZOLR2tC4T4HJPjI7wIpxfLr3DJ3fPiJSxEiUdMzUnlF7WqU5skl4
UPkS14tmHBtiXC1XjqoUK82aSwbJS7IDB+4RTC34WztxEx6jsgGxtZRQezKsifqT
N9Lt8NGHqGxMd0WfmavIDvCbqsEGQGT5X2F/jJPBJgGAxM3ihZFv1HoNt7g1bAkv
`protect END_PROTECTED
