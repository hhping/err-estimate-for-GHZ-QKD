`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IQpAi/3+G+U2CHMIRKdi3DIeailT/V18dOSahK+dGXPrQUEOunO4EaTOlNymwz0w
U+9H2KG8xnoT4+azfNsDelyqjWhOtFPzzYyYcWLfqI679mn+oZhZfsQoxP0sPyFg
yn35Yrsu5jy9AR5kHT372J8Wrcd3MvMmAZKCow4DpkacEP2rDXM3I2GUTdSYQf6s
p/P7hqFenJUwxXbP0yYeJidNwFbRQaPAt82e1So9Hnb22IO0nWzc70JiZmS6WDMI
r25FfzDRIMnqU11sa5W3UyMRxsLtjvlEsVbGxapkYi509XjLfJ9B4fc6uqXGOjj2
+j8Obb5MYbitGocbP92XPjyFnwJWBINtsMjiLGRzR29C5tKY5lXF9Di0uXsnMUS6
Z559H9qsYp8D4NsxlQsotRRBeUGMxS7WeHlSIPRO0DrqXQKSA5xQFXRiwx2eT60l
McCxVbURpSrxu95RppEHlZfhlAaaRJ0aL/6Fhv04dmCpFFcXX0/Q1KKhl/SFE2yU
LORezPoBXx1ca4OJVHI/UN9SpPWvfrzuv6gy1hwOd16qqorgWnoJUEYvDW5PCpmX
yw5TjtMUO+7WV/alp/szA33TmQ08sv5+f5hbMiIYml4UCvnrKECPHMyL8LNtYFO2
nnrI+eggJg+GUElqQEqIakh4f970+4z9xgd9WvUTzHLHe3/ejBnkFnKjMJGTJkcs
JnvJrtaEwsXBhTRKfiI39uBbaBrKf3whAhlaT2XS4T3B4KlgV2+7RWyi4WM9utII
T4qc5jInnSo0iJdtqNA2KL8lJhzmwOCQq4Gky40XQQ/4yb+xaI9LtE0zWVfSEzdN
7oB8y+B24OfMtj9sHTCMvzD6JCQXBCaUtMClQy0D46/xaM4LAh/f5KSNXf8KxC1/
MnZCqrHZVOIfQn7QqUTdvoe5uyo2Ae4txhEbL+/LqqKK2UIlRwOgzDI3D/BZ35or
vnIJSZlrq/myYSmTANdUqcmW8pMiBkd1zDOhktgUG0s8mVv9p1iL8f6DnJrRd8lp
P1lldHbKqOQxTOt2/dxf5/9+zFVDS6r/7PXgYSw51d8s/Scj2y3i/O/iw/SMqqAQ
lFGL+6aWHnaO2PkB5EdOBKIVZVKsgV61j7G4V8SPii0jEvj5gdeBtkVumHf1QdkV
OJaKZ51YyjyJ2IHCjUN6lQiCon2Q+MiJKRG+xXdl2IpWIstX2G2LEaYsUTfa+5uR
o3rYpC8YK7qy71ZlbKmsZQhbhxMW8K9N7nrO3zxHwxI1IdTXR7ssAUHzxTLrca9X
9JC9mDB/cLKa55MK0ltMzcRmnttxwJRfIT8bs9DAVPQnzMr5A+tSX8z1SFIUeCDd
tqQ6vuPQyM97lw+xPlzGsP5aqgOVFfpxRgjX4AzYqJk6ZUqSLlPSlOM3kN1NWVG2
4nEeTZLVEzsX4M6vgjmpuBGwLMj6SPez1ydI0uWnZCSoJbnMDeVvZfY6aWHed247
KM6k/KAuihg5nuS+S8bAZ+aIP0xg+jJSTBT4UwFyRvOBMZTCXa2jRxLnnncev2yk
SZGHaAPNQMdx6tkN5DtEO2MPi++7HzPgNCV0tUpxQRbgSPRfADLpXfNkqMTe84ls
F2R/MP/NcQ/D6bd+XlOsKjqweUSB/B+gZnO4NsrrhNTDQZd24PUPvDsJp21mCpJG
8yZlhLJrQuY3QypFkmSOuOnJYiwqEuVjTlUGTe+0T7gHXnhZp4PpoNoqMtI0u7Ll
XcHi3LYn9UhzuoAGgXVB1JWp2eDVOFu37gQAXw+V/6x+qTybMIw5i6gNPqXLfdCg
KxDgOlTg8MmqIPHRnUfXSm3ocx1GvZeg806mHYnkVVGVPoMRLXD63yHaZvlfDMC/
9MOO5Zna09eKjbf04nApchyw0fgVdhFrecLn8EGecZEtm1PMZW99YkvSl6Qf7lEx
c5Hakpw4sFhZMRJT8sa+5VgH41evGBnkZkUe1tEdKjRCRI4JN1SR0oruLTn34Q8c
qbSfFe9e4fID2ZXhaKP32XVKQRHCsMSR0MRnKMuJzK48g8yAq4NLf5l4Y77ZAVCZ
s12SVXH6fSbtWtqMzEgVfO9aiO40WiEzlXd1eH91zAbCHajBGsa/bkv4BpKmCkOs
VBWDtwolE1VSulKNi/4zD2zPunHMCk18AoJIAfm+r6RsrL6PItzpZxwgwWpHjp1e
bIO3THI6SAfGbeH4ze1qR96k8T68aLlFh7F20Xd4jcWUMGpupyefI5CQHLppHrkb
VyruNMokcNCpeeAdl+JnqoG0pvdVsBA6hRW6tkyDlXPPXufqNI2VD8ZWRqw5NPUu
+MJjgIj0Uu8CZkfvWHobC2qoJTRZoFGd3aTqQ2ZqT3NBgYpnP0XYYslKO+TTqkQ4
3QuISbYC1RQS8+YltvxuEDD6Ff+c3H9pWZDtCEiRQcVWFjYk3sbSITGq6AgmTHxo
Eo87m2AUx+tzpLm50cMgUYaDVtMw58Jgfyl2fxPqYGbxUk4Sh6Lovg8ssyoFkQtf
tZyw7mzvab2NNmw3lg03Nny1D8P6WSVqjmj4MXOcm7NGiuhmlCBc8jx6S7OKSoA7
IEVsBw0mGTSIUF9CuoaiJshSUI75pdQCFwc2FefXh3pOaq10w8SxF+Pr5o+D2nxn
v2ahQVPZp0Qbk7EiwcPPmEf5xCFYcQkRJr5tjeaMmnz1DzrmB2vea4RqWosNFb7c
fAzOPctCwVxjeH1UEaJOtXxc0zCPe7ohkfGtJ0g1cO6TFfo7/an4YYu1ovJzmULD
cqIxYsIAxrWQVQR/MqiPWj5kuOvdUr+Np5O0t/4xPKX4kQgq/1agbZFa1P1Jb2oK
tXhZmjRrP8Z+WADUp1/iX5kX6MHYGbrW4A8mDIDbFPFz1KXok9BeYRvY8Dx5+CbK
AoIkqCGqIAzZ4t7payKXsaQAFguKJEWXrH5MaXttwj1MXRnPJXgym+jsRW2no7yt
v7GAZMvOaIpGb2yU7W0fkHQHd4Ee4bThLVuSEzFCvXK+xZhKcZ3O8HxvDdjExpdu
iGkct8+U01r+7XoW0fB5Bn9oxF3qhUpXwO2s2pq4tJ/EiuV+nHD79YqzKerwPdFi
BcohnOusqFxSMzwnR4ruz0d0oKx5yzKGkbPhukpPFwgk3NkFBqVnUZEQnWaGA2Op
tri/aEzKg7Deomph6GacHDAyuztkonq3WEBZpiY/N5s6ckUwIbBchSVyIwLIwymx
P+GpaZjesuNjSWyjPGsdTXQDUecj6aDUo61KIS4moM5ELoWe/hFJl+eW1ShEtGW0
pSg10RkMuvqTUQ+H7+g/ob5kSXd6oDaskzNpBr8wy+v5DBg/qLiuTsPzS4uMs2Dc
WfCgqIyMrKPR7A0lUb149VsalT4k2r3bu5RRpRF8pYCt1woznaFbaVrEYjU6t5Zk
lzba8aB+gmmU/3MDXfm1eKHBi+gB/C0nsf6KA3uiuAaaMfVo1C+pAGGDxy77Pwuh
suoeMkA2ZTlT27t6Pcx38FyMLx2A1YJJTxp8Y9gu7knHyoxHzhAmeKmsyKDH+Utm
lbFPEmM3ytfqP8YmJQMQVt/WA8/gpFRMvnViDd9L/NJqMoovjv6OXLTDKT5YIYap
jqS1ylsh3GHtJHgdqKiFPmWRFZiRC+eP4Vm7WFoasp4mzrB1JmUoI2UsqtyFvGn6
9bpfHhbFGJPO7RtuDk77MpVJENELBp2TtFe1WkuuMDigvmfm7BS7pd9tBRR3kZ8S
0LaZ7VUTMs8DL46aTtIx+Q==
`protect END_PROTECTED
