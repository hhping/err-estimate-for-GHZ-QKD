`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I3SxTm4liiB1+9hUy9Qp8X9W2+wo5dkfy54dYegJgZZ2solUpoLMKLKKBMkABNa0
suassamBKUPyy15wrTGRpyumdkNm4XnpuwcRmqZaP+2Gd3KI4mmUXiWUpNyaX3Fz
PBEP4KgT9OM1oktNc7bZvh9r97ONqapr6tiVss0mrOl8o8UeYl1yMJa/PQ//wiAL
bArbdj7bx8K/3K3stq1/8eg3MJD08MemGhbf/bS0/1h4VoHmIMjamvJGy6R5BqxO
Oxx9kZMToRiX+DXovV817YtdBeeIJMVdxPji3HzZdsaee07q4hFMycgUeXnmRtHT
EkhmbKeBKcebNbU/T2p+L+tATGNfhvHOwWhijIVKLvPe2CpdLwQUXZmRVeR/hcDb
1NC/TJzpPBZ7cK4pBKLpQO97jrxFYEKs3LarT6e2j7DC6wfqIdvxv0DdZsFh/T6N
arkMav+jySfhLriVf2OpgGxs2I32yu2QVJX75XpmIpAToJxxPY92AScN1REzsJbp
aDGLDd9ckIt2jnRYOFfk81l1NuOeI66r5CV0DP+9XEcT3sHmuN3PZu3s+S+mqgqP
/HzS40Hf6rHW32c4dxiTLA6H1w8wrCIVEqdyCYzZgTHHQ9n7ijtuVl3Ffy8+xeYG
L8HmMd6IwQX2VnY2JXz6TQ9wrGvc9CBXvfUJ0TzSPdaae4sGBv4xN3pp95B/SljB
Q/FlHJ6jCNBTLnqY72FPcVFmWguaDYHcH1jTUdRYdHRGYIGKETOa9FNJKiqxLr61
Gb2urRXc1LNwym5fg1uIhhapCm4AjgmTJPU9ABm2ApI545f1w8phtwpk4omkgedF
su6Un/fYe4uVFntshWCpDW30HQlQoYr6NPH0USL1ET0nB84KB3VrTr1M3rLMzl14
zicG2y/TWFhVFeJQERw4i9W/QdFbMeOQ0CJSHXQrA/IjyV1f3N6nx7tC/NaTY4HP
cMJtKYyAfAsUkPhnWdjxzeh3AkfOONZvIebtDS7ScuyTvdaDIwhArptylde9yXTP
dDQGD2nuVAWl6hW8fWPtdHT7yd7KZtrahuh4/yTArnd7TWU3NFWqEq7vpImbnVbs
h3Q2Un+ih/h2Y+NQ5M4ZTzawhg+F0suLZ8HI0vAm1EbMKxAgChVtRPsNUIM3Pis4
vn+hyqbvvkhyldCjhKAK6mAoQjueSFCCIbVWjmCsqsogV8t8REdF42sxVg+BEFj3
RPVaZ9XZpeeySFxh8fgwfv+rIr3rqm1n9qH8Dra5rLx6HjPZOTR+Na81c3b2yoK8
+S1wTWCfBZWS+koVCI8ML0tjzmlFz8FFm1jy4ZXsyfs=
`protect END_PROTECTED
