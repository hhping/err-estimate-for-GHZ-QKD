`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/gfG6iLmYXM6FDZDNYfcluFxA9GEg+2qa5szyyUzoOOYzQx8HKfg/4Fru9zCaXHn
yD+xCSDQJkadHCuAoS5Agws80M08aZ0Eo37lnaNBbVRfIChPDAlowrL4bZELi95m
69x1lZTtzN4oqHKflmjJitDeDQ3+GkH3mVrZVXzCIXhy1D3hSPNRBvygLFJTfolJ
vWpownENRV3VVaOcdwjsMaDPdgpm6hInTiCQkxvUkDzeGp4uCMSg49uXXhitqD7a
KWV8JIZNa23Jent8ziu2Nt+O7MjjjlflIvn8k0NvhsTMS3pQoUplcLSDFNsOr00O
Cqzo9KX5w0F8mvN724Zs1hcmZ5JnZRKkr05Sykc9Ehx+6uZqZEUapddWJEytuLA8
FxImVMR5VMIojvKihFJ0rQbEgFjmFoXR7TAOCj9svCW5BWz/W76cF1s7MVbNwvhE
ydGyLE+EUoX0r+6GFiMpliO4avXGhwcWE+7cT1xehx0EJW0ZIziv+/6pi5i+cxCo
iiCWoTi5vqmTe56MaFN864RXfnj4z59pvgNyUEyUq8uEiWykrTOWUomlZjx8GbEO
QD53oCFRE4RlOVgX1H1H1e/sKBbjSDtEjgLig+nV2dzHqOoXJnrnE9r0klGdDdt5
ZqfzDcOhNbagB6ZFpi3YtCDMW4hA37750b2AFGyEkPYiFxExtTYXReyysMzKraDl
FHNY59o5CTBkgyP+UjYqg6li63WkKAgC5SdP/WU7UapYlqhGGETVm4dLbxfY3dQn
uqstDMhqFKHUGVuz4D8j/Rz0dOJxRURSc4u9APFyLlU=
`protect END_PROTECTED
