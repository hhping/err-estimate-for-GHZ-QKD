`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
22Rk7O6MIB8AhCXiG0Mf/Oklx7d/8Si0KWwO30loptfUgjLcn//ZwTA/SbbHwBQI
TFG2vRZrSdJFfyWJ46NTyJ3BVIVBnpIx2DxQjDsQTzgo/PuR7zcYJiuSGs+8VU/r
XHRnmH2ofZPFiDY9tOao0SQ8jDrEwbRv2DjKS5HXNa9kcFeSxytLIuve0lmGr+/I
+N1UcpOAIOcVMjNLwF4yqBqtkCMEToYb6XnSTKyfB1wHPY1qfJlg4Bsgeg6sJNAm
De8IMX01oiIjCA0lSRd5/dzQGKFl2bKaTomMaRuk1m1O/tTLStaAGLQRgOUsGyng
9S34zBvqyQTMgejN2MLXm5wg3/sKo+j7Ztc/+i2m4DySBCfojQmhOH/h01G8lwmr
Qz2KcvV00aJikdQELMu+PTLTVaRJZwJEAWR82GUCz6eCLa6si0nMhCU3z4jSKe5G
oGAezvSfs5B5xmLEYQ6oIul/NBSqvBuUWsQ+lNvnAbr5OjaGtHNAlJZsRUmjPSSq
o4TKmnhKaImn4OQxgPXnk0y6oq9RSXvd50HNxbMi/pEBp9EQ6OyPslmGDzVUKxDB
IqIkg0e+YdszKJ6ENZtg++O4biqpyxZQWjAzKiGPmQlKuOHmHvqR6HQn+q3S07Ot
/NCckIT+YfF0brh4KRPcBOTFywYD8ZAIGSJF+0FAuRu2i1Egl/8LTGscAtyPu6j4
xiLNC7v/tzV+cAOxUNODzE/Mr1fRzUMG30JdD55T83fMxhZ9hmeI85qPWc4gn6OT
5P7lVC52pesS+z5SU3dRXoz68DmvZTDDOz5mQfTxFfNneLkOa+s09fpdWkRn1XMj
raGjbxfL43bpmQ3R/zggAqZWD6/nyQjbCkXk8hMzDbAlpZl+R76ifWnAXTtMPJ2D
3WtbbYBPOeGNzjKGAnaOk1tXq8zGee2y7ulzp6VM6H867ja2UXjwV9Hvec1FINE5
9Tbj+TT+VphrF7Alj+cc6CRu0ImYGB5/umsLPB3QsIJV9voi5l4Q0lK2Pk5BcCun
fbDTWe95tVtbNduvSKKdBkBodHGXMeKZl0tPJaF94EWRO758+K8BKO4ba+jB6Rd6
pj4lSRHz/N2CJFstkT/2RRF35PsS39mdZ4Y42wXydFm+HczRlSUHLiVGtnIydNUJ
jb+Mr4eHHjnk5K3RSoU8njKPRxBE/U2iwRCHa7oVHT/B8m5IG2Ng0oIP5XzxK7ir
ok80xImaN95zaLH1o7LP3HSj4SSqNjje5A5Vp38SNjPLprW2cWJGwwMdKbTbCBqY
8k6315TiIrLbWgT2bVWxPIN1fr8jcWatorjA8RFC8QJuk4Rnjon9ozZUTEfnPepd
/qNKEi0AU44FDOr4TDtUtrUCh+0FGtqf74USa8GMO0Gwh8UP84pbYe0K2cEomx96
g5jhmgsJ6sr4/ych2MWgOOmxkJ7c1l4upcrrAs8oIExe57WuDxu4HAlGHz9xyMux
hLcYr2U+194bCkx4u9MkGkPQSDQlINAM2BV1L6lytqzCqV1CN2b7NZTmbDj5FB0Y
l+LHzuKDvyQVZ+7TAmilV4YSkUJyZAIryp2Cd6rIya6TLvcxWg9qcExiSoFDLbii
XeLIblT34vLaoXx9mev3CaxmNPiHWRljkEgQ0gA8dCX6qFv9LRtamyEdXv22vfj7
6AigZV6tnzXNXBg6GYPlUxgE2J+HRbcz0WMzjDD8N7hjCVCjElvzMbK9rjNvJ7oV
S3jL3OQCBugEB2zuJhfFgt1UBqQOLd9ehtmTqvKJkz7FAGY1GUWxcFrwu0ZfzF+7
o05cq2U04lErfBnLZ1d7xlQWoZEfYciM41LPUWd7UgNVvFODNGoanpO8HEZ4SXEs
leNRfYZaCiPLbL/HaZWU2nqdOHhu/DDDMrSgBkALeuiwRr7iVlnNWE1n4fdXyFHP
OHSTTny9537bFO5wySYGTdRWAoFnb1ArvViWGEKMiiw5nVWa7/SN2mCH4m5G9ALv
x73gWLUZpFgSQ8i7cGiZAqJhOqVWsjxzltw3HUPuqUzd5mmMq1lB0TZ1cM3Rbe+0
Y7KFHRsz3HwtTWf/Ziw9M/u1xA718TkezMroE9ov3cmQd1uilnDQB4hhGSjoLhMt
AXz2MHBMVPIGORWjpqnZdXj09sSHxLo+e+SvSm6ofOrIWKtKQmzsk3lG8/lficNV
kuucJhrMjwDa86wVEO6toId5GY4hXdaQ85s3eO64LVmH04h/nHCrRnGfNvcNrhpB
Wg8DXpwjtPYg8QXDnZppMfBzy4+s/QyTdgyUpO/FCXXiQTQS9QCCyBMO3MBTOEmP
/V3TUQdqbLjCmRpbmfT+XOC3+l8/5C+bHQGWQ57PY8JU2ZWTOgok4XI14BmH8txl
suw2yTS0QJNUaJoU3nvk+NY4My0WtH0zTWGWlq977ilyWqi5fclQ0RNBLmZzOIcX
PRWop9gZpx7zdokLbFRf4WfiTyNKGjSBKukC265o2ZcJJsSa0/j2pP/RgUzjCaxJ
LMlpGn7O0CVadaOmBIhba3FVOeJ81HlUycdVaWi+NvT6bnmXHjpPnWq9czsjmYpw
P8VmKnD3Nwsr2xOpYbR+NNvPXtg65J7O+1R7RYpAeYaWlyXVvm0Ti1cgTN8/rsFt
NP4sBbbD+g0w8JcmgCgwkOnpJXesZCJsKCSNd/fyZu5KHHFILTUudzjdNyPo/teD
hmt9srlieEpWSu5UM0p32iNoJ3tgb8t62u9zDYdxYLrmCpyDr0gqeea16HJYdOAm
zxgha6I+qLtS2mRakMG2VGcYWLTAodDlbRGdngNXyAY8llsFGyoT+fsHRwHw3zi3
DsvcTAfPXhvgsnN2A+oUN2ag83oIjd1hLgeHKULyHGyBxdNJn+u5dutU+eoJYdo9
F9mzAsQEcfKmKq+KzOGrta9mHPIqysgBSSfUTTh4vz4CasS2cQW93TdUde/GzlGP
Ejv9v8qm9CSn65YSC2L4O5pCWX34zKUSfIubU1TvoJqRVgJvtOuO7VwfFpwYDGIE
Lafpf+snIqvz0iHeMOOSquKaxjapN0juaQrDCZMlQZI9zwiBXrJDyFqe0uqm8hhS
W+h5XnwBIjYdiRCzXbyqz5hb1cELgqvTDKjTN1ZzM13evovnV9h4jTbox6RL8wAL
y0SdmyAmFfzs/ZN8nFxhhVx0LlfasGEj/GeAaljM+3owHm6bDFbZrYTdsv4ZbjOf
etCLbsaPKchaFA/l84fEd0bE+Fj5zZlQbDAVb/SB8GhysKzw1Km7GBEmbQ805vj7
8Wpc8D9ESj5JFMX4RRUeNMxvNtIC7TZnQx4xQEvF1zM9YSyhtn9CUo6ASrpq6xFL
sFMtv/uHaLva4BGLin5jihdonhHS/F8qEvfdc8Z4v3xm878dE+YiXWsY+ERXUbXB
YBs+XSsBQaSzXur5OIjR7m0bVCKXKp2tYFANJFdzT0qJWzheklp+bYQzk3CdG8VM
ozS8ufLZlPFtJBGKRFLvDPlmgKOdh0/U5MDVAJybCfsPK+QPtfpjNMJ/tvunaJ7E
7ln0ZsLPxXLAvbdA+cVa1QR03lJyhWGUb7ABdzBqeZNUXqQHsuMlju+jxQ/Zwmg4
eKrduEBeapvhOxFmrg3Avxu/aEvUtpnH2L4aE139aexQ1gv3PSWN+qdOINCFqpoU
gUPbdxGqr83tTPkrrnP6eqALoPWf7L3zLGOhZAgeZZwZ+qmKxWo0R1xKjVUNV48Y
/TdeVl1iv8rnk5qI6Jo//t5WogtGpVn/NC9E0wfrtLNjLM/A3HWQyNJeezKmmSMM
5jimM/9ATCydTJFe9XNRZYz+0NBwBoFkx2D4gpmPXxsiS3pH3H41a6WLhBlyofUv
8hHPn0GpGvLMDlxXffFizLgLRAravLbKnmIVW5W5gS/4+r2Ql0Q2eK7zmNoCqdw7
Mz9pmGE1WGaVYIMktHknjlclqnwcu+FL/44Vtgufg9yCswAPUH7TuTSqQHgBG5ei
4T1TrkUQ5YJUh64PoZlzt9XyTgXW567CM8xJmKuEcWiFOmPiQAjnhvGB9CCNCzld
lfZmqUjw9c9VWePQ02yhloEwYqat9QDKTwIDdJfEhJOl2mN7i2wTsz649rjx00Qy
hv/fGMm6hbN2RZhJDGXceaqE7Ma69tUltG42kMERkR847undpRPKZ6pd2ueonsJq
oxxByfXBp5kssiDGMCXgBwVNpMBVDqlLyHssA4SR/maekiiydUX0qLZ3c6an+9Kq
untLRluIAwqLSuoPVOk8oVpnbfE8mwHB84IvcgdWOi/Fi1zDdVJE1CH62qkC72lm
lgV/TVlSBg3jCdijS4l5BPpn+MJgWLcV3fVGZJUCamH4UGUuxYSrzAuUgsuYp9AO
x71YluaHkb1pbBUzmiB5GvV7XFNe1LRF3OcZPvdO85BiV0yvAJihxV3OBlFz/jfZ
J8hOTxHeEjiN+MyqPYcmoXgijZoHtzwqUv2ryVYfabYQTugBBaIgcE1M9McPcIYf
4EvqixfA3YxCjugVzeXY4rmqrEABQJzPYNY3gCrF+5q7Je9VxO9Senr00c/uLolG
AEvhjxwmQ4XqRzhxhhgQQpdJlXj+tKNJ0KJaiYeAhCbGTEwtvW1//sKokoYqzjEV
V5pthkwJNu+4Wfnn/tzP0ps+Lt/c3hHboaOUgEdx8C0QiQoDxVAq/UrHFHF66rKa
8htEASGecIrjtcMfadxpp+ugmo5pF8eg5NWrs57q7v5Zan82OXTM70yC3FQQXbWb
Q30VUArO9V9W+ZOLJKUBkHAwFeuR+5/go70t8ryQtIASQDcq5xGsDPjkBbCCo0uE
Jm8/Us4kTN1Q+pLRdFZXLIUoUV0ci498OOrD9QGf87W8B6hAgeXXRPMRF+8iDAH+
GCDDiwT+hL0zEglGocB9Ss3Fi2Co2ik2eBSdx2xa4q/wF/ubIQ9x4Yuv2sjrZqgj
U18JKSl2wy1nTX8r64dlbmTH2wqxfcN+HgtAvQeJH+Dbci5DZGRBVku/Zd/3RnS1
tquYq81pjWxiEMUdHdEoDh//cOes7Q1PJh+/OeG3/RBRmhySWU4cuor/FcAmO64c
LtEQmNXKe8Ine+ZtbsD40Z7/a5MhLJu1FlPUT3PIVboTSSeF8tCbyPiUFkUQrn5v
YAgXyo3WvtD3WYJf6eBa0Qf8YxujGYSKAJXaeG/fz5Nu5dGY5mUk9bequ/Hig1Sj
UB6s9/wmZmUnThDKbMHch9BHNZhv56qzOQf3Dfc7PC6dleyP3G0wdcw5qLnD+6Wm
H8oIrYjK7NJdARGANIC5vUMoZSK096huMCwnAglNUeGfzJESaPEn8Kus3qereO5b
HxIPUgKI/aE+GksN0wkeKncXdDeJ3HsU2fpg9asX6NUGHRKfo89Yw8jvWDvYCfc3
klLM5Q5qaHGHzUpLT8jX1F3CWtL5E3+bMyS21dQ4cYqp6oPsraQQVg8hznWqa1IO
EARmBxqWXGL721IhFm7mw+Am33D01E4dpD+rbM/hEXuBI5UDlWLxjQjmc8n859pw
VhXtIxCG84Kh0UTncZoVTcM6A0q88kWArLH9BpNINlP4/0HevdMJv/FjE7lEO+Tb
bMNuhqCjXsYNpcG2nfQyXVvdT6VdGTZSzz18kjmcJvzjYCrRSBXzuKXkmHDATz4u
gklzttnbRO+YOeLSOmR3WS8azEkrxzOaUGKxOLCzR7EdHPQBHpU0guN7WZQrc65o
DYqEFL3CNgcDEUZH/D8trLS5GcsT17deKynAFkWAkTXB9tQme5/y4xy1XutHF6bQ
8GWdCt0yx/fG+65RZ13yQm8UWW0aba864tGq6yaDnCjaPipOh7Llz/mGksu0PGxM
dxFkOVRnvmHGTqyhAmhOyxbR+62PHV3LwnGTqfyim5PCjyX2Q3IoUhMt0P2WlMCr
NDTl62EDUztAvaiR3uvObmDsH/nKW5wd5GYJ+UI5Y9S+fZzVzuaazWiaJc/wEKeI
1sR28f/PeQQ4vbmnzmnSDOHdZSygZRMNJ+XdOmXBWXnXb+GHGNLr+J78gsYFAb7V
znSBQ4kf+IYlit8fedgabaU0jikcBFUThOWETo2Qw+cRlOva16x/+LAFKeaTHxk8
kJGvgDDMaYUWCkjKyyA3c8Ol5xdNNmPxAFRCatVZ8vZj9NCf7gDqS4nVyy5LCspw
JX1NJOa0x4EnJvpoxAv1inRfIBTEzG3uN69Beuf2tOO7puJj8ZBDobuzHvE6d7Zv
sLNDfyfOytwf2qtgeU5YWH7RI5GJmuaNuwBDLY5fYxhNfmfVhA8PlReMWqkkBOS8
n0JuLpJXif4huj0rZrd1X89+I4ZjI6OOU9ERhZX1xzcxa/yGzBeecioOMkgjXlhv
u7Onv9FTi83HY7LVJvHOO60nFnn73r56sTYjRNYRgCx2S2PbZv2Srb2Dg5diJjVN
YTD6WYYXcccmBkUGJVFvltfjmkB6NElkckc64z9vyxwSZ+6452JmH2JBszxFV0g6
7/UytiW8FeMXH/d/eJOkiZLtT++58Lun69ZfZRKtar58GZlNkEfBB4TMbH0/bT8d
TLyhgvcGRWCxTrxuidCrhRJAF++scWdhEay/NAdfZfP0evjEupVndc/GfjvTkiP4
LaWdCyme0MGuK+VYtIlg/J+8h9TRaA5+uymJ5lkhwEKOC3teOyTphymM/W0eV63w
7a9TGE1KO17IAWOhU4n1X/y+UgL7SIHBnZvaJnbYMi0DmRhYwko3c/kLdKsqUIqS
+aFGLXQQuTCNC3po785ecxFuhmJaEu1Ns0nX0xakl/FQg0Q9U6fH4smzuuOEm2Qd
Kn8YdXYw6ZfOuMs994vaEXonNo4uxRtBGOiOEB5wkEzZZTxHRbvVAwh+/GPZ5ken
jkYTesj+FMoQXUK3cZVLHBpfzGUZmzDTAVCsEiqszVGtAKYNZwUkL8qHlYW+QX+h
4ubu12Lletq97OChl3m1Au3MCFhLzRNFvmEOXfHzvQ+P6EfjrWIDza0YiVpPZmWy
WDVG8f4/SZcoh0xmlF/AB2280yS8fpkov9tjIBinN2NF4cYo/JI3Jiv49/WLtsAP
kWIEwfEAKOTYp0RXlT0FZcMxILpXxVwdAXA3FWVtAom7Zp75YS0LwTAmWe5NigP4
C/mAriZSH67KvObCBHpn0Wuf2nBOV+DcmzxKcwUTUvgdmOAD0DPD1Vq/grsZFhMZ
Em1XEhw3y6tYf4bLRSqoSkj9Ls2HaHbCobD/ZTxqAGwbU+bgwSLJf7I2xnO58JKO
Mmbl9k2PnlrRmKYs8ry6W7WpnbCIUkI0tTPtl4ffpgzv+j7ZvzQ4FVsgaxLETmSA
IEqBEnv8yqKjrARXEOdKgOgciulQEclSCdeqCpyZ5WgcCUsQlIPAkh0a8scvqfCS
yw31lej91XnfsjTHWrw3LcqL2Fk4OFpfnsTAfBPd1GQd5r+pSCNGphfC4dLiK/S3
Jl1C6ge54bV1MBx580YMtt8j7u6d6axxXxfPAPU+r/W1iYLXWUyD/DNpgfpMminI
Kgty0oRikiPRhXz52t2jO2wAyAU4Q9t2ZayTA2eEbjgCQeX2yuBg367crs3qJT4u
z1JevcJasqXjZTbgQGnuR7IJjbw8Ku7QySDrEQO62jWWWrXEZ1Ml4R1zgshYCunG
E8LjBZ03CrPuAweTNZEHrGSPVfZZiUCAZXWnDtV531l07MR7q3bKwmNfdMgbimIn
SSF4EhTF5ViWxwwXC2g/ie7TNIaG3svOeQhtyh4H6Su3aqNm7Y9iXQG6XsevHjUf
i0/NCghdAjgtBciv7GaseoWvxrvhUfiyJVW09ozCkoMi9M4X1bzhvX4oJiteQgEM
2+O7ktuF4ogRoslL/XCMNhiVhuddTTEoioLr35vTPp+eOjpFblu7yJUmWnefN0lV
C2bYXiopX5t2Nfp6XyDx4ooqZVlsfptwSoTP964E7uaFmkTU66DbvTcDaMvG5Zrl
c8hRJbyAXZDTf2a/SDTbPffKqD+1lDgw+u7mCkD4yschykQY13PVMXSpNHZfDMYo
jUzPmDaPxLlXXThPdw7YkPWVa3h9QOVJCV1CZDnKZ/eVlTG4wpmO7vWDNDOK4qCB
JYCaA2C44r4YIQgq+ahwyJUoJL06lg3CrIoKcyWKiOnQQufTQKwwcLvKRLTpIjiz
riHuzWTSdGBYCsfLCgbsAAgcFIWKMLBwNwr/hilo8Kh62Yp9Tg0BEFOWKkbvA+6w
8EvDxiFwen8YOEeELAkr6uuZqlU5M8z4aa4IRP7ghGqYZbZyGAYd0SXJhzlG9Ow3
40JPkpcMnmkCCMMARV4lkM5TAtAsweLTsosVYFee4et0mLe9Lp+ALwPSFhk90flJ
5Gfihji8pY0Uqz3Xbt3B1YpiRH9orsYN9pYtFrKpOM7S6/waKjqxnTTn6DYGRMi+
3qslZFlRjKnLwdCcKYQuXjEb0d19MZUQm4eT9v2mSxM3MD/pQlGFSHC6uGm3Z4fk
m5zVZhFR4mVn0JwxvB4jCCgdUt/l2WOskznyK9GWzWb7LvTZBnMSP2bdlQ9p1Hf7
/nU6YfYcNrAYeU3GZmfHT1XBZyy/mI+lHI9MSRptTVqmcFj/aYHRMlpHKRd30TQd
QtTw/9p0MscMdeBBEM5eBkO525xYFPhlTmneDBMQnnhb1s19ym8jbfG/IvucCQH/
TSrSIJ9sHEro7HAkPKW9Sy/iHlBpH/wJLFsr3it333EFjTn7Ez7xLnYG1uGzVxsD
l09TJKym/uLxWOT+b9bCDCkD5gDCmJbZJ1VVefejFHnXhD9q/KCCp9qiutzmfYO2
mSqjdr1Psbn4y/mVpP3rW4J6BKXV6nbeKI0fKziJsv7LZnhBhSbjuOuZ9DnqtJeQ
`protect END_PROTECTED
