`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gIPbRUyYm53maRZ5ZiDTP1Ig4tzt/FAdzpNCavdZz8PkHoCy5KpttDQuPO4th1zN
lZyrDCyXpyI4LW4b/YdiQJHx6tM0offE/IJf6Das4naQ4rkBhVpSqsFXQ+63SRos
1wnUbqgyVXfDqVWRl2k5bBh4yAlIJdVP6w8UGHlydy7twliKFMmijgP1Um24lfIE
vDKN5FyyRBYWnJn55hcC/GCD6T9eh0ToeqFJ7HYqgQ1Pf1It9YfF9a+DZ2TsYeMx
+qNX2X8YPMgGxfW9y+3/LOfYdQ9NCEHVh9yhEIVxxSxRmHBXHO9nxMt6DRjYdZOq
zTgdECViPQGz1yUEnUyWlOZGN4D/RNoiNpeG+y3sLzcj99nz2gW2UopZ7BhfkicR
v16UkKxrtaDXUpXw+o4Jz68mGKfw8YntyMi5ctYq2aRisXNG9U+IKBsiF3UApWjs
oWWN+RbRITz90ik4y9g9EQBEm9Pca5jif/SiJuK0X6iIgv0TDetTAyNvD4LEGqHh
rreK9mXGRPNa3OFsUH5dOHsFKq34xdIQ6LbqlrYAsNCKZN7raRcFJsZNgFgTjyRP
OGD/Pv2mllzkmK3iSNpAlDgtDO9qNkKwyXHyZlmILqInoJLy4c9gYuioJI4ABXwj
MVhUKUFs2n/SRTi+/MMiYUKC1tHRKU03IDfKrGSr2uPd4IRS0vUctLXyRMfV67Dg
Pt321mVB6X/E6j8C49ZAtSMoaF+PvRpNr8I6td6ky5/KDkGY4/VatXAFldCXw0fc
QbEjYlKfJ1OrfzZDqNGBlwRdkt2chZXvqAk7TtEXVYYq2vknSny4u2cWcjUr+BEd
q5ShkKpLynSRLOK6omEmqyGHWhs96fBZCsvkjjlaD3cmiLwb16qZ6s2yyh1jhDU2
kVxpGNfXrtZfj/g0t+SGs/QoB2VF9kzPaVy7XqJuhrhWZJxFF5MjUUBNCHkQCwx7
QZH4BWFLBqtOPpoQNphaj83hvQx+v6VztZIkSGeEC0nsnaY4/v1XlttcRdCJ1LZN
j7V634mfo2mvRIFI1YUkq7zN8KPnVdsF3bl2drTu9QUz0NpSOXX43yCIA+Yajq6j
5b61KMguZvXSlR8JKrGHJy8wEv2d5PXe9jMe4f7pWtlNHAj93nSetn7mhb/CBixl
gJcOpGzRqpw70Q4wyWP33cJNGfJqYpZmJC6qVSzYmeFnKrx3VnFL3AkvvcmpQhOZ
LpAk8lP7Wc+P6wIqCy8DIsuzbYqX3zdM1dBV2xg8KS+Qvm8kWYQD3/VzVIDeYkmK
Am0CRATuApz5ZgMpHDWDeI6Z31kPD3XeWY/6kMplVhUPqOpC9ow2E9IfG/NUXHpg
`protect END_PROTECTED
