`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2GOZ1uZW+hgVEBuPWRFEFd3LADODaXmS75DBrfj2jEZNnhL+XNK84iFrJZ8kiTRj
RQ2M3NAtofLj9NnqtLN9tGeTz/oAZryGMW1i7rao82S341r/tf8xU9lS8HQWVy5b
t5q1S9MlgUx3vtFKIylZuN2Ej07V4RB82CS11HQRakzAJOYlvxchYRlje05N57q/
iTtmMj90Krhnwe9vkBe9DfRAel+vTQo7jGrpotbgvp+5h3IqIpIw4HiuY96XPnlF
G9lNwxHhP0eegP47IZwCGun2tspVdJs14M7PowKHBkqZRl1zyiHqpGUjnMLLAR7R
9opw5Lx+YgzH+NgV5bs/eZXC6Yg9sh7ueALlVQYvaXtvFt6ppoNVZQZMnNIHj0ec
loekp1ugC/u/aflgvqidQWLKianeQe8ivgtr1OEPWJVi7xuaTOr48RSBsHBsJgei
zPSpmNeUtWdEsqyuwTZrWUixl05Tl9QNBEKuJNDiaCnXxlLD3yVH/kgVOxtKb0oQ
WNIRzqk1v285ArHtz93PmYrUZvv9RyGUkr5tdNRZTR+6Ojx0UOn77n6fX58lHV10
iBhYVTEWd1xaL+CScQXKiISenPUeeWFF57LwwFDCrPFokojzsWwKcJqRTJjWcU66
xcCAeGyljzRY4TLYCSHAtg==
`protect END_PROTECTED
