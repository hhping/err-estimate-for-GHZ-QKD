`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sIjtLYNT4fuFRmYynQIk4jl0XzaTpohoIf3M34agQ2Sqz1uTk0ZL6xv6Lt2SA1ol
YbP9XuhC48rBzx1Y/TelX8F6HzOw07pjX+cQoBU9ntqyQE+bUjnzhmBEw5pvsNc0
3Fr4oDlb+0yfSAK3gFsvMLqSUCsBjG1C9xbp/9YkuhFM6g7dF2jQuY/x9VhvdrYX
+1LpHZ76fm+P2wDa9vvThC66leUCcou6f9k3JIeHbinizEo3lCzeAetKbPnTkyQV
7Zzzflkfq6gSHpTtPCZ+A65LjuNPE5kkmNYif35LFGKSJm9vq9+axdIXnpk9MNqD
F832zb15zL/GPxcgQYeag8m8qpHfnTkdIFlfZGYTVF994sWhuF1Xp/8L4PoMzRpJ
vylQiVkqznXXulveNC8jMq9A45nKaCYF3ZwEio6vJj9azsA5BIp11ONVs3dzU3yY
Des379Gi4eoTQMahf3nQ/3gVzphJMm1kfpdajy8JFo+A43YGcMOcLDySULzjcELf
+sAycij8YebsWvv9vtOhUwTU4q/eryZnU9dH8mSNSswgE5k793fBJJMHGOf00a+g
oXcWYGaCXC0zKyu7NilRxIMsrUH/LCBlUlGGgnmZzPqvNGcgHNFcbBnXQGe33Ii8
xDaxJRfs2BMWllZJ2xPWzzlZ3KXYS9JtziFjpufTCnaj+GP2+FNYtfr6E8dVu7JB
1v3qWi4WyR70fu9GayKj8Uyi585nXPiYdCNa+ABQVeem5natl6w9K+wyvGASxdpE
90hvZCT/5gMUe6P+VSZ5PieGxV4Ld7q61bW+WLaoSHI=
`protect END_PROTECTED
