`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rp8BiKRBwTCkn0KcMCAn+eJt2YPI+80TRGZyaY7+q4Saty/mG8qYxJoRxz0iU+pV
Jyz2X+xvcZ5eym982eNHPsOJlS2ks5HarsYv6Y0ZSZxKcsSpVx6t67XQUFUoqjCx
88U7lbJyyty7mLwI7bqXLasd9Kx75ZYK5ASnrrwi3fVuvqsr4es7x1F+SUVwR+td
eXJABVJgYJYlb0BJYJjUtcQ/kgqbdWKpJqcgwTbgxSUIVQbRTNrRJd4C15rqap/Z
0j4vJcFCAnxbdteTVa8oHuzpn334qvLUUpFPGmSmsNou5j8+uDpHn4jv1mW4OENU
ZRMb4zdpxinp923WHGy8bKVcY2rmqsa7uarkTpE9ZiYpsDX/W1Tc1y5xXr1L2h8M
W3rJnXhZd+UF6i93e7bFr/S5/6sTw7JBW9FzR62pAt5tAznnE2fA71WWviejPSkV
SBVq9DRtfMboSO9Wx6+zQ0bIhiSs8zZkRC+ele4buAUj+fybRxmHGDFlBHsUhhUJ
u7kKVwAEhod8rzNxsM6dsCkw9kc2WvHwx0W/7YUONLslSKIzao0O1RVLAdEn4DbK
DI3ZY5DsjNVcaf/yuMMVWmdDvMrVICf5iafo/kUx3Q2CZgeVk23pPx7m+S10tHdF
HGXpdnwfAf44JbhBXDHqYyyIUNfYr5DjaTqjorXbjTkW2Dr9Un9n7GvLXTVqk4tt
YkVLQKu0k4IHc9EcFG5bbDdw9Q4segwkb8iBJkWP8e1dJPxq/P5JPvDg8tvSqqTi
YuY3ezgJxb7DJuYkLgp94hav3Bbeq/jR47QionRD1gYbQNQ464le6Zgf2wiZGxUC
ARsFlvSIUQMGB+EPBaqCDi0rjr/5zXM88okMe2gImMItSHNnquMCeXN87MFhwPdN
y0W9oUOg8CdOVHLRxQe5RUQT9s9d8b/fDU0ndBF/NYPdouksGxxAUl1pGvLr7sdg
NTrMn2uyAyreaGdhzWXr4M6knozqPT85ah8xaDFIzUi13XPz0omo42K0+O3rywwb
Y0HPd9rPAXIUsOgcePe2eriMUm732MJkhznhHWPAL5Mg8jfgVSq6L+BK1k+K8ys6
qBn7Y54YLqgrivAXgHFPS9IIIZ7gshKuTS2NDLYTtd4HHQu6dom9RWovPM3+OHZf
0oH5B+QstvB3YmTUI0dnLMQbKAxmCwqPLNO+35yVjHjsSYBiEtJ6ahDPGuoVZi0R
YSZe9osHW7PrtyPBtRYY7FciJCYPkadhJMStOBSx/9u+RaMzfnoUFd5WqnE7lyCr
Y8vgH13LaBJIpiv84etLW/5/5qZMYRfPU0r8mu8AtVBwJ/fTtrdgvbGsqmknvWfI
SI5TMqBJwWQc+dbxblu0hIgEmgOhBBhJObycme7uOnSkGyGtwKIkcbzN/clxgU8n
ozcuIJR9/giw+gUElPDMM/o3XHAI8WHFdP00ZqfZOcYJaQhGucJyidm29OMLRqEh
+UyQ/fnkbPfXPQOQaIYGblGb1IZ2slY3cuwZ2lahlQtgCmfQxobUNH/J3TaAP5w1
POQCPIyMOmJcN8rEyt0XDegrGEHJxe0b6DB4fx0HEFYvUqtrAhKED+28gej0WarA
E/dGTTV7FOplQVPnaPrFYBXAfhuRkdDwHCn1forOCNuHYaZTjOJDUWwNeYpYGmV8
MUoGjCLLHbFqcbMYaUNXEqdWO467Qf7AakjJVP8K5/7ISvniZ+Ald0zE1gH+TS4K
/NixrB470fg+MT3A1V7zHUyDtDogv3eLqW81VDF6CZ6/A85wtH2DVSgrWrmMMBuk
B/b1h3OuIFrfzlTsM60vRLNcJ3C9NsTpJ9Cf6pFv285Qew+MM9EC79IvE03HOU2s
/ykN2rbkxE7X0DjzKuouUyTLvD6hD8f8RCYgl4s679S8x9bYK8UH7rwhZ+SQn3+/
zq4DrSpCQ3o1ExONFIAQCAZsmZj4VV4orwADCkfAdg/EXvY7RORmphqaeoNwTRuG
9iw3ITrQ+tuER5q6bTKnt8HYJfjd/B174Ru9SD7ou8rOufS6G/akwfnCRsUdEcJ8
PooBz2hHRCujlKJMa0wfrNtjsK43j06bfqlmFg4t1H/hD3Nfk2o0rT2zOBc4LQ9+
19JeB/5teYqLhT296iaI0yDxYVITnBvG4SATJrb4gRAPIpZMPEPL2qoIdxMSAYng
891OiVzR9s2deAsj524rMiLhc7qM9sHymXutw8QAq0R8umJamaBK+XBp12zOwUaw
juEALiLVXTKYBw8xUftGbgFQZarvRPzMVk0xrndGonPLla+KVHE6vWjMecBc8OVe
/Ncv6eVQPQyXzmkepZo2SiEeYECgU/Rd/j4d0sS3++YvqChFsnyLW9QDXx/qhONe
VGix5eAki9PkuZp5H3y2BUt8DSOOX9u+XGrG8xQBjzhy0Sk++W2Reut2wDBtZOh8
Frmi3M959VdOZn3+5ArzOQpB7hv5NW3VmLqPW2cOHEK6NLZj4RiAgXHU5EnP8Ofg
7oWUROtlDnOoT5X9xDvPkwpsv9QcmR8mWqLRyW8dmNMRBt3bK6wLsS4f94jJlqet
ZSTVnDo2DO2JO5t+Af6Smlg7jPiu115womSL5JaQlCmQMdb8QlMUu9UYx+yY8hll
4YiLsvLpFRapsO5G9njBLZfkbh6snI2rTl4zF5sME+TjKg9IfJ6HrnymtP0b0JGU
pUm68LyFwrRB+wsrx9rKtamKtlm+8vV/hm/BMI5waIQ9QZjhr04XHInmrBmI7zRd
fu6HFQgPueveWsELneE2uytcrHtCrQ/3I+FsHxxGTOe+jEL8nz2rMgzm8wzNDpOy
p+B9ykTo2C6MoXmrvDFnd4FAi5FRpK4XUFccOiiWpW+xSxiDm8FVGEVw8Dah1T0N
QhWf/fRdrihLfsOtWZNpjtfZEAYTzxOnIoFXAF1FKY2IcRqeV+ERe5l4Cdcacynh
jPU5lSu7T+ORTUdb5d7FrQtOgukGdONoAFAOevFyd+tVbKXQQ+tywBSd3CxzadoR
cX/XLeM7T315p5Uuyt5+X/phk5bzgw4Dm1kBmyvbF+4JYUR7bmHDgs7+s8u8WYKe
gJYjUdWPWZQket92jjQnI1nA8lyyXx5PbrmaFJs/I7sKdnbcvNvyXaa6RSiSyr/l
pWyDnaXOsYKvh+lOKIks2l9yZno8EH+kq1VfdvWDHn2cwjevhoBbIZhMAlLo1h1N
x/8vDQaj4X8ClfyYzeYNi8asx1GE9977HWO980PRetTU0Acv6q+Q/Z5vX5RFk0Uv
F6N7AAiyEU6gfvZUS0rBEAL+yWElW/50nAWBBdcUpx2pzHoCRySsqGBchbP7BGTK
0wdflgmHYMei+m3aWqRpVGXoQjAaJHstu3Ge7w6Ag3F5kfzZ+HjsXcDayOZt9E2h
VzhC3+cdnzNv3EzIkuhA4b0cKfRx+A9BlpasGwV64W9mJA0V3UEQbKKA1UCG+YqE
XhiGTlJk3rBUfqBgYatVJQ0a3Noe4t3Kw+qXkvYJAWjcaK+LJNzH3HgvMBJpFVQ8
MAqTQwbHQE6NV7AJPYDlBTbvYiFOiUqGg+N1HYrkZdFki5UWCOl9Bnqa253/IPKM
F0wUBTtsgdQhBTvhHTlQX/wCRENrEDu59bhdSBfKsLVWdOZ6afRFQUb1omkEFQ5s
r/bYN3Jg+NwrRk4xF0Pir4ihH4VsTT/HsnHnsscuCGNLA4sjgAs4q/VH9LIV4mrh
kDKvnor8gBVhYfDE+ckOuMItwvdEOiAvQ8MkGKdUlXEtyi685BGlI/Fe56Ki/6Ha
AURRIx9ABdVVUjJV53t/LJC0xuCntg8w3hACEB3QDRzSVO2HSbP4YUFHJZaXIbWE
JFQ2ad5GKEP/u7OPboPZvGn4S2w4mZ5Q5FuNyThlBC0J6DDlocGJ2Lqut/eGSChF
xjBM3ZtxYC29P0imY9dBM9gtOyDWPQiH2MqqpieNSpIVnS7rI3O88W97ujkQksD3
104NSjQ9xqppVrxAlDBEeDiOJs1Mjt6aXCuaQg1/k+TJoz5CxufepdSzlqUTabqW
SPx0QdvFmcfWkj6YfMeBkwanmCWBeO5q2rv+f1QAvvtgoEHAVHqJWaCuQLupA1fG
kAgt1Q+QQLQbr2/yGKj6Kw==
`protect END_PROTECTED
