`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WeXU7yM//+KC8fFbrqBImYlTHgKGBKha7eap5lQq5y6776mdoHNUIQfTSnRTY7ah
J7+zibNHwSOktULLll42jWuWaHCbrASUVo9qAMs5RT6TIwordWzd/WuQ4LHZx1xH
efmCJm5prZaWt7nioFKIK5w+i7u8MhfbXSJ1vD9t4i5tkB1g2P9R+eih7WhgVZaO
v5GRlLUJ8EISvwhaoJESJRI8HyNhpZkjOaFJVgQ5aSH1+GfDQ5w897nk95Tn66Sc
ZDg13AP2T6hyq/ROawyJJQIspwOc601VNAFmx47HXChCBhjPuZwumpd/ci6PSnHp
wVqQ8c++oOpj2tKumToaYR+rrStt0n0TthQTahFGK6L2Q/UJQGKlGOow4E8gTgsS
RsCEql06GeQNYLoC8oVg1Z0Z+oCRoduuV9j+lg5iFDNs4cvuzeIBDBol8TILIeAi
RPiNDSaRlBSvZ7Spcm0+yBhG8Jm83k+mys9QXfKgzoTnWO8PNsjsA+Q3jfMrIlpb
oIvTmwyO2mELBFdFS2uTssZ52d3FAwq++H9SmMFE+VBF9cxsMrv79q2/FINfM+5r
kQOp524TWdtg9DPli/LE+8Vrw6GDSZW2OeyBfvvhz0JBVZzFJ4VVQT/IIVTBxF5N
9U1/9GT3aZDrS8KUMCxUqMOT+tQZFsavvHyLs9dbxbQhEVcW5UZSRXZi+BmUpi/+
5ZL3CSA0lJPjbIHer/HPiQ==
`protect END_PROTECTED
