`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WJqJih5iAVd7S5U3eZ2ToQc+l4kFTbQ+GWas6CEJwXej656NOPrGwGfuSpnLWHwY
xRizEzNfNW2BDubHjFStKMRVN4UX/s77iZvIsXyDdeLRJAlZIkoXqhxmzzR/wshI
etbXQ+qzq6JQbxZzE5eovYWFjlwsthEQaK8sDEeQagztWYi2nsKKfU+4OPUzaXwZ
ETweM4B0ggv9wfGIiA/Hzw0j59KFeCtRA1tmuk2lALYkJdq4eeDSew/TKeg6HZFF
VHpjc1J1rJNlMqLdZaYEYDaOPHWJBgnuBorkInSs/7fuw0wRvLBLII4iHpf4GWj1
8oykPB3tol7HbPKoJOCf5az1jKsl9n60hLwHnr1o/4Bi8lcpfeTm0f+nlki3ESpv
yobLJRUyzLkTv8Fgf6vYl0UprIFgwLvJvBuCoWuyh/Ch+q332b+qW6FJSC0v2l9o
bIlqP9nRaInX85g6OLuwK3s9WE7Z3n7qo/TYEdDFLnl2FOHtV01Vt99XkvSy+NV4
ftuXu0MW7b10bleuDnFigd39Ox0tSSlzK0bAaQPB8uOGNX+gsFzKCquJN+nlOTqi
hjMHiJXoJebbnsTHAXRkWAtyyY/+oWqHoyH+23p+NDDqB+Sb87inQnByAlfsHDGd
CiKoRVUlqV3L6Qd7cYIRBdk9QPBNnn4/ND5f9ViRp/EVesiLFn6fNuy1lCK/+2lx
rA9TWwviyhRKS3nYt+ov2hZqcAVc9EZxVYyQ2dUX7NmYw/cf2gCViI0jDwryJvlx
HoXnL9l9Qu3JXTKh7Lpm42YQP77NFO00iV9mtkWhnMMCmiUaOIu8AdDtRTkqT5IE
RjDP0poX8B/vL8LJZj9NccDeyTBPQ9XCixRdyM3wBkHABuQi3Z4fI++8snHZJtz1
5/NvLakhx++Ja2sZE6AMW5OgRY1rdOP/CY5HrPhhl+deroLkro+rTk5TZOay6H1O
j1H0wMioxNkHMjsY0lnjZi4pCAVNNs1llVE372TKG/RIdUA98vOeZseJjYvbqvSJ
55tRp38CcgM1eh/ZF3ftZfinjdRfNJpiKEr0fkUUmdBjNVbNl+Lote4yYtaCb2eB
Z4uDXjncFAzZh/6jldL2WC7i19v+F27b5GfYILouaeDk/lHJzyCs373ttpOhGM8O
PsUF73V9RcVyroQtR+7v2XWAMXP4fLgRDWm7dOSTAfegX/i07olQd4nYqm+9Xj8j
2Q4VLRb8XynTZZxjVgp91LQ0WgSTfXYEg1dxpA1UhYSOQyCCuOKHEd0uBMmYrTCo
mpngppEAc56HDRudydUe4O0n7nc7BhCVMa773jMEuTXmWvSpbMGBW62wD7gBJc3J
zZC/ezWDMPIBinvOppi+tKN3IrTnsVWKTfIZJjTpe8xZhZT5q0g/kA8mu50Ie/Jg
XYjBzRtQiGpUF1OON115rkscWdfhOVEfbIbJ/PgC6zoN7Nn8I6kN+zT8vKiz8F2l
nAVJb+/zduySPU8KJswL/bWXtCqDGsRWIJfgwoOMHyBZ5enbdlR3gHUq5Zb2UyDZ
iH802sqV0guZSbzWRdMWdDgD1GQqXA85GAsxf0rpNw8g4H2eqSZhj4gewaQXY5Tf
oX1nztgFSWnuDDrliWLWvEnSMGklENo7iWVeOyM+DP4JMZRAXEy/i2EePTNPy1/V
q0ywFN/rr61fH1QnJwwgl6JxAXCwNGeEbyXfBRZ++HX+fW8GthyFhDxrSRylECdN
HNs4XNoXxldp7W+7wKs4rrBry6VSBB8L+VSBRJB2we9MYx3oZwQbMBtAcGMQbYmm
O6sD2yEzlbd82e6TpMa0eKEx9JVwb7yc6E58sdjWtjho6FYHAgqIKE93cej3ICG/
Rk03vmZ6xKW3sM3eEOk+sy2iLLAsTOo2aWfF6O91A650h5oistLi/JYaSgOlmQiw
9sG5XExBm0co5Jk0SD2B6oOqPENdsLc+8VMi/PgVX2ZV/sUEwPhR0wGGEEa99dcZ
vp3nOa13NdtSi5bLv/Jboxhc8RiKNXMwFCFWh1bYh0QSk5aDw7kUc+IslGoDLIXg
iwzY08CpVRsstlK6J/D4xTTqgYeHLHZw9Ni3DlDciXs0g/E3WsF2M/CnmrNZ2uUL
FsI+QmqbR0wKHsfZBVSNsfPt0yfYMo8Y01tvEEAAj3aMsUBKynDCpt8rDV0ovP8t
OS9UwrdLsFFHpxNuVD28NoQT51C38BMEmDK0tO+G/Crpc6fqJGRkBxXNpkexhHI9
drZxTR3IdKgzEa6fl91CeKMOtCicKoF0iFX6X/ApQpyYDREjR0J+J+42Qf1hi29Y
aUlmaZByORBoZ/koT8tuGZDDoYndjDrUY+VapgjhFO6gn/JZ6UZjAmeGdL5u91fI
wa7DzPNQbdVYqO5zNsmCDjEju028FrX5ZoKg1rrrCuhGSYMCZMlzBdjhiRpUACX8
fws/Jta3+/QC8VP+bECeUOk4VdoZ2u9gUQnz4MlY3WAoxbgkWEi5Rfci0KXkGNvr
ky6ZSVbcCOZIbC8WvhZ8i5KepMU14YWhnW+4hTERKB5y2svZILCfWvh5UeFIuk4F
dDYxAC4F/381Tf/qSwfxLpuFOpBWINKdi7GsocMauBlNfUXw5Sb6PO2Bd47zxaAi
EyRftsk6x3AYPD51XbhD41LPReHmw08RwOMCEYQMJ4V7ubPP9AhaplD9saebkyTR
GHI8Umywx49v+IMN26NvVJd8u8flIGqwpsCTLJlAlI4WhmuNCUOo+pfFEZbsEVFY
ufmA76UuGKOQy2cZ3Yv19R51HLZ5cKPHcYgKqPmp8KiR2gGR6uJfqAjMaHXUgzFj
bSK37hEaRKCmWI1GPPb/xu5QfFTn1E6HFWq5QpXcdcMZDHAy11Ky3JlXVwk8DAXe
dDyvQLwL7wHzYOr/N4NMmudCTb5Xx5TG7t6prNIp+Z0aejQeChYNf0pyrUXTVT7G
R5fUJgyS/PiGp6A9DSGt+YUfnH3TntEnHguGdErAoenggd0DJi1TbWkb4V65JEqa
xWOM0dTNB8Tb+ohZgseKSUndCkW34H/C+NzX7kaw0PJgcO2grTCo5aI9NHQqLNNt
ZOa+j9N2IiEnO/emA31+mQcDJDeUzdAPgf+XoDQ4nLOmT8wiociEKxPD5AqzLW16
Rpb6GHUhVzs+o4VBnPJ83USsvSemItDJ3sebKWfN8wbCqZq+idwbM6sT7P3An47H
5m/poFzADY29bH8aJ3oI+tUCL1SjMjSsd1bsCFeyhNdeu2GfV2GpIOiO2sv+O1+v
2D9Xh3Gp4YvMLUwqsGDUdjDDAeGTe7eFAlCfjnwKX0KjcNmRr1JnOCeLC8oPZ77o
SBUcfXscen19YaAV37YqkBoZOU2wzXq7TwjkUBMersLG8eT4mPE/jIuP3+wj5eMd
bg8irI6E+FeiN26KXMZyFikYFu1wepMi0oY5tvY59HiTDIdliCpOQLiLef/fXcMi
BVaC4q0DevTE/6YxDcwM7/OEiR57nI1UVa77RAqmMLwRoiAAR+/mBylyl65Cnwaj
F953AeRQq1caSlG6KLzvfEyNq3Pct/82+gmYC1aHBwQXQSbiTD7PkIYMcp6YYx7b
vye3lTubox7KjJUoApsr/4pqLY5ZJWlV8/ZzsgOJPdf6Ip68z+Ga0oLVtipeugfr
oU+DXOwrTxCvaQ3AjxyiReRScRS3AS5owKLz2fRIX8YW358fz7OtkZELlkeKVyUs
V1tNFb911OxXIfMg71zHQmSDSaz8Xbr23X2zQGpQ4hkwDQdqtE/Ad7Jt4ohUNWOD
wWN0uyGkjHidZFU+fiaVil2ub4cWDgrYJVbkgX8QKpwGsU8td9Dcoru3jxR0BCC8
kp3GVV5M0jnQyOVSzCqogey396uYSrywBDQF5NJkuWmqeqq5s1PzLKRJYXfxZxFC
7Th2o6GvSOZ/tEd0bSs4tFww/p8IC8pODfUCbqrzNsDNgP+IQVaKOgWa+ShUZvmu
4ne4qemyMZZiu8iQ6q+w6XSrajmHmRHTeLLYl4RjwPByUtXOpyvKvYo++p2OCFul
2ajaJMkMXRHeiHZF6OqojPMLoD6KzcUVh4T8O4pNQKwq1t89W/WRE/9pCJKuMSi7
d+02ApbikmET3uMEY+aF3jxxbsDqZbvuc1OTmwXeILVPFW6FNE1S+DXLTzO+S3HE
/r6R6cw05ueXcNriuXhpBanI3LOwzKqyEwiYeMNtMZZz3+UNs24gZO6MBCqGYObb
B+ZZusD78dwp//PKqr38njE8c6nUIL94uIQGvN2m9pADmlVScB5BxuJcqpi3QtKk
KurBHjs0VAxXYWgG9mCqy4hCNm7xcxFAeSywdwYjGdRoPFMhcZvBrJF7vEqr7+CU
iQfadPnjr0sSVWNr1QfQxcv3woSW3JaMtjELLTUSM4IrJnGaCkVZhzzR+JhoUwkr
MWtHx0pytgMBSD3EqUB20R3672SHTZgyPtT+MrgANnh6gNqbGOraZRMcFKwtJ7y6
2SDlRZvJzb2bMtnTFZTLtBU+1HjUYurZgNG2shXuBgovDPyA9+NBZXgw1Nk0YRC5
WHy1iJL65cskFPmx4XSprFmTQm0Ek7fpCzzoxmmdZ+0fChs/XDQLa+PU0MymG0eI
Qgx5cuVwvlwbTBOwMvPs2FzkR+moBZTk+yb57bA+ap1erDWStQ/exxY22CwnNhai
fTwvGskPgaTc8E20+UsMcyRaGuzeSYRmaY6Z+pE4p2mYSmNv1PlHn0t5xWGvjJRT
qiPMMdfPRBaZsUSKhj/wHim5WgrnPQsW9Dheb/lMd6tl391UySAhPQ5GIv6vRUUk
MVFg/RfAN5qLDGVVBcF5O3uRm7q5ldN8cFaslOA41radp9OZXJgmbQ55psqfe6M6
H3I6I6vPLCseIsFZ2DQcu8iXIQQKuz44S8dgoRGRQ87GryJM6M1GYVJ1KG55Rsmn
ebupKvd1Rc1czzFXqDEEblFWgW++YMsl1tldpwJ57y38rfyL0RRWXZkJGEwtYKzF
vjrIlK9ZNRziGGvFM/E3vzAmRAsZ7INds7e5oPQ3pzMbNRxUlD8hCjTqQ9TIh+uW
I5kqxEU31jIF6nWbBT4ENiWa9hp1jutPQwllww1y+LsuqIaaXaokS7y+ChBWMUgz
HSd4cWfMYZvymF+8E0QRXWJQpU+bN1E1PLmv/nvPDGkRQjKPdjqQQGxBHgf58t7g
uGGiAl1GAetbwjpatjAz5yS7FA5ISCXGNCqstFgAVygaeDQYc+oG7FDzmXg2WBet
/Qes8shrYp8YEkuwdKOXpRDUh/BYeOWSW+9f/E0oup4+9033tq0C0TPHvM59OWDj
cJyYN7cX0pRW+w7wiHf5iGkGcOrg+nVVMz2/CYBhbIFrjnV2tjedWGFVuvvEN2L/
cWi/m2UwIy8wfYZ/NDKpBOmo23FcC8u5kxk+MpN0h6DDv/Q0A7ZugJwQS/vFq9kL
9PsS1Mo4ePyh1bgR18c50d/dN1heQsLKaXtEzZIsGYWfEaD7Yo+PcT7wgvl9Zh+U
U3gBHMW8iQxNhaMl4d6O1LIZOHdSTLMWI3Pyq5R3HUVmtIM/tWjyWgOXFSOdbD4p
Zx6tdeuCQnkVfrY4StyBpKYkMBbpEPUwoThO00d/b5QOTils66Z5fk0lcoqSMV7g
D7U0POcuetauu8dYRcH74OK5EimPVTGcuGdX3H4Yh8ETi+9O1YQPQLryI+4OeA/j
x5hYBKbrGs0ZeGElayMvJiRpMhY1Btw9swYsSexucWcwO7exJyyCCeo9mnkGsJt9
WF202QNARaOXrkNJEmVrVmOSeGZwcgpFUb6EsY+UIAaSRhHpzcKgcjRAVQk5DCXC
iyGzSBzPNMWDkI2kZRjn2TZrpAnwl2DP9u/Nqx727AToSkWbZ6dDrZSsqocl2DAC
xzTWS2Q+UGqQ4EHBl30u9UDwFUmX8Glwdl25Ji524zuDFL2IAU6xpm2z/eK9+iei
CX4qxS9/vDrCNBSpzTCXb9MQH5UBKeM3hKf4grzRZeQBbmLeIs9McxDufQiy77yY
jpIpAv+DyWzAA9ttxnDATjvXzA6VwA4iy6epyaaE+bg2s19EGOBSY2um+HXW2Cdg
FZMFrE8U2UK82Iuwl7vTnWIggh0umA8V+EjOdTXrjUcioDLd4b8OUIxujmpnj2Oa
fnz9wzvBlWxpO3aMrJWnCKT2t5BRktOC0edq975z+mLweyikxHV176sMMvk5Nony
BNOmEKCIruQZuvMlHq9pWhnFYVvjP+BF3Vw1ImHtdSISkwVa9c2USSFAcc/iauyx
crnZLtqJgOz0wzPsTqhlVun6bb/zezmQHRzKh0IkmuXjVE1WKe0lImr2syA/4UkO
22KvPLnlz5WJB27tzUlMkFH894veSYTjBBNtlT26EUqEphWdf8NVrUmV7ZNk3Fu2
skoKw/SYDAiKrdXmqjZAshfw6tgCfefSUXwyHw2puDkTma9MupRojB2MwQu1xYuF
ab/Qu5okxDszJpq1zyKKP7XnhB919oejxIuQdySfSKlaf0jak7DmzwAmICsM0Nhc
ozid4gpDrYAHaVQNfD3eDhkAGOynIlC35tbWb9PVQRTTHO8MzH+ho0EneaWaa+RB
MK2pVUdMxi1a+YHCoYwVpZ/jb0bk0lUitRyKjlKCK+v/tiVDLjtPeXgw2Kd0qAm5
p6V+aMI15MPvn3s3AU+yNlmLk9b0pQ2ehrYrkfGizLyDxr8JdER0o/ZmXU0gvofo
fE0G+WNbSWfaeH97TiBfmFMDjPOuQLBvhKgxuBeg58YfRHCLW6SmskrRiM5htMcs
1UUbl6/zW0+WAoPAI6L0UT2hERGriP7t8eFrgX3PNWzsgLC1FU6SjcdVjZb0FtUe
qVTprUl5qIqI/SPei8m32wEIJdzvUKa5jKJ8XRD2auCBRvWp+goMmzRcSgw5ZhMj
e+aZETfo7SN8dHaLResJ2q+0m9Ctng+K1W/vjAW6a9Q8y49VKHT7Y4c+E0y/0Red
hYQbC4SsKr+SaltQY8btzGp2OmYzPJJuSOLHfOaycig6qS7NQPn0Ve/Bp3ueFOTK
sNBXi+QPQ9/uESr5ykDrZ7TpQypBCmijD/ytyh9e1AGgV4twu2jZLRaD3xHCz9k9
UVvvpVKWQnvQIE8myhTD/fmK1V8To09Ns424/5swtqmTP2NFuV6VDgJdNHM1a4bc
ubhpjcAbEoJe8n6WgkcWyE3UiF9lsgk9H1czDQj0RXrrWoEWxBfc6jzYia6BmPA5
EmLC0f5O3dZn32ayHCRqOvfU6iXX8jiAzC65qteR3y7gpx2e9yiiE3ai+RGuu+GP
LcZyCxgkZDvaFs6E8EPGglbidL8S5Kg7NdFqDw3Gw1vY7LD7n6ju9fyy5ihz+uap
b3mFeUXG47xw427gmPRr1kHPvEPpQ2647KyQLPHCYeETkjz9edoS25ebtiP9WXPS
FB0FpWd9pD/SFUPmFtTuq7djdJwt4Lbsh/x1MB9dKcEXUHOd66CyukF2hCpM5OMr
f4zDaa/418w3QvNq+Xh+TmWI8d+0+5zVS+o0OQh9fF4kDo388cTw3YX6fX6R9DXO
D/bJdZYatSkwz+0iXo5nGHafkK46BEnLewx/hQ99PzESU8jv4IhHqpPZVd3BTibn
OWJzCEImfS7KRvwN/IIYVb4nQTQ2l/geQzp1K3VWp+wvvHAYY5BNkrBXCNRWYw9u
PDbngtOavIIwXynq7gOs4WJE7vBnCDxNOTli4hSa21so1Sp7/ASNSY4NBfey2ruD
GzeZ/0UNdHn+fu6fSvkgQ7SEQth4I/18lVC0hUufrLflqLKoqvM1+GehGtxJk2/4
9pkf294vuSTBIKIZeAhng1zxlaAaNiF1fn4c7Ha/8vP0ZSzZNucJ6b/TSkm04KFu
sbaARTvT/5fE23j+futmvxij7lIc7Bmw9B/jP4Duocm8syUlKkyNnsHwBi3Ts9Tm
j00jAZGIojer2/Ag9kthyIBti078TpcXiv7O/JKBBiM6jKroT38tmjHloFikPljo
afw2EryUMIEMCBUsXUjl4zewW7QrMUSvgLKmBc1FJVZfO4QjjUbP96vWnV10an3j
T99n0zemyAsbWObTjF2+32RrXGZxxbEMmiisccQvUPU8aUouZta0SIE1Q4pdSj9D
ahZpimRh9fE6uIFQp2pbu9cMeOBYwY2SAT6CHyZmny9shab5TFCNHKScDNz/1fsR
WZE2TGKuzOFUeQP2diXIsFxHRV/EDrK0HHUMHO/4oj8ESaQtI1RbEURDrniOzZ7p
JzT2CVswSRwkc3kh25VNJk+aGSiRCnKO7Bel670VKznO4HVpQXXgBCLSrhrvk8Qb
Rp1DQmEg7ky+yAZtxoL6KzRMTGzV/FNjZcroYEFLJoM7/KgyyI6NHsUwVt46uLeH
MM7sEp0twmhHsQNuATC40o0byo7teLKTHbBKfGdvZifSOH+BTl3iB2TySakix15r
CacO9zV43amzWL+AaFbh+EBRYwC4dAANk8C8DZuoHv67t8i8m10rfgI0vXHnBWPh
vnFTHjym/oRTyFfxVlqvRTUGujfis3516wPS0HE3EQl17vYcHbf6pOAf3A9sxK/H
nD9uAp/z/OWA89cPQjWqRk+h39QVBejKAVNZWHJ28oiZdwcXxNKfe4cPtXD/CM8T
4l6xznASiSUxdwdERS3wbmlFUY4dbkRfsH0Sy9XtQZiUDoEkwNB4WOY4Z4uKHP9N
dbxGVu9cxOauIVkpwfT/xuzJEaTg1Gf3jfRcHpHHngPAl87rUdcdbmdsy59DN6UN
CxgZ8gZhpAD/6Wx12vcC9z3ep6Jt6GkMw7ML/WwfG8s5d2IF8indazAO6wKAsg6z
NwykgEeZ0TkuXD5wlNVg0mWijeenoL1+CLzY87a9RVMUU/hNFZETGOdypfiHL9oS
gUZy/zB7EvXRyA627KsrrT6DMqcjzdd4+sj8eI2qd0UNoNefTO3pkvN/SCMPQUGn
A6JIBjB63vqSF9nQrlvNnSxn+5wliedC32QnLT/zQspqDVqumFTqpyjIwIvupgoj
EGqL5RjvgijNkLYa/tqbQ3cTwwhBz2Q3Dun3+cT9rVN7SxJ7Km9S6Wj+wxRvh1PG
6dF9L19b2VPy8wQx71EqxAhn2z/NNewIxHcD5Al73oRSg2P/IZbVKRKuyviYzO89
Uh7mZ3UDCwTMS/1m79W1qkGGWsxIJu0eiPljJqCBe49lyKpQdNErzokObfquVFwo
Fa+DNlmTJC/bJEqZvVR9w4njrJCqHQ0XPzQ4tk24/QBiQA3vz8ARMai+/iVvXBOh
Ed33xxTgN7UZrUxK2avvdIVAj/Tb3wPIN8gKc4ZNisWWfjwV6opfRvCvtsjSX6Ib
43fTXeTM+Hl2sOzxVdXdFAsydIgJOd+GD3eSVaedCbN0XdsOem92QMehq0tUCaqp
BUsBALuUFf0vdQt5YhwLHpplCoyGYMjZVmchBYZzPfiV3r7a3sjG9tlTSAz7XhMw
EevbO65e4VLP7sEUdpIsY+ucWeaev9GteBxCXrfo0QyDvJ8/utOJfkNLl7JALSg2
L3rp2dIl3gTC4K4cbDdC+hpChuN458PAIHVznY3BlBIGh76cZLhBA19PUMjeHUYy
faukmRjHvEFw0YjWhAYp+0RVxnYxEtXArBSZdZeTERgf/CuA0HUad9hYf/pO67NT
eF/0E+kcKieAfM0xYOAV08/dGHeZvL8xOE8CFi42/Sj20MZYC5JTpwstJxBy8E2n
0Vs/LS4AifU0KZk3KWHxaGO6B2MK1xU8gH+dyz6l36/a/8psCt8MpPStnZB7wAYd
WatcVWPejYW7MIN8U5YJiRRA8kUiIyS0KpslUEcflJ7UkGRnX1gy+1oXHE+UZ/8B
zZmwZBrHXr5/asj+gLXr6c7znyD+U1gs5DIQGFMghj1GHQyrE3VJ5cQkbYL2pJEM
nK8FKnR4zeikcHMwh+Zhk8e++zmSB4BKEUBnxXaQXSPnQldVUEk77FbXWOoYjWM+
NnUyxWAO7AP1eN2toPCoDN8T+CUFZlZK5fk+vG7OtMkEE9n7oIB/cEoacnIVBJHt
G46ayVXbZ/8cFKN7j0t/cqlIJ0bgWbCqJAaNdpC3IIuyVlkA23VsfWLrMqTfk+L7
oK+YAxq4E2iVDHIv9W+3cail+ZFvuJQL9+3n/GEzZUvtOZe2MYyn8l2uUIOwRShJ
FwJfcjHBxJBL3jx8sQ+Kkr60315LFFmNSVbTUoyc/Yn/ZGB/zNfOpfcwndWcv4Dj
m7Ol9iwtBB5k973tumqyDj9Xuwryjali5Foew3vrCU08DBfSLYcANq72fKqibfhP
zOeu57qXBygyp/xsbzP/y+/mQvcmnclWFUElNw+W2NI4JeD7RQCEb6fQQwX3JbJQ
/LCgTPTNseF/iAe8QVyufmdSp4MokGYbukkPHaOGrm4sh7UyKnnAgHUQpE9pQ312
qwNCCBKHI4bK7lGbNBBp7+oIcRnMtacAeZ98M7FowWU+ZFuiT6UnfWetcjht2M48
xvjZJQR2g7pW7C8k+Lwooj2KmS1002KbvsnCBVKeo8DLt8oEzz+D8Ag2r2kcA1sE
VgPlXCyQE45JNJ6LZ/C4ZJ5eJwsjNCbntf/DATNTdrn+Mddx5KVZKYdZJQytkROB
nOmx9pVGn3ZWVEgCuGh88aSoljv8Fuf6hjU2aFfiePnj9MOxW4QB5zbcs6nmI4Ho
rsCL7JsN4BKPLw5iOL6XQ6q5af7iyLFetc5kUrqlOBgzrDNhM4O6Gs0w9YAvBc+x
5e0TyKO1O6f3SiaC3O8JdP/9keYfwiRkRhNlhETwbGMZARBqc/iKPyKPSMLRv/VL
kvKETVr6WXCCzg1drkYLxCdbl7CvCvbbKFpcX0Zmh5F3wNSx7MGdv7NIv5cY96+7
IW81u6HPz+xPgSxM6ghhMngO+mR/FsQOTDm1iwwR4z1VamSX9Z+X42NPqNqjV4eu
sBoAWQBK2KhBaGvKTJ1bZfqfdrki/XKnhaYVlqylsktbf4Fkz01LfU+gD8MKaTfr
8M2EYn5gVB4x2R8EDx8ao/7uQHHDQ+hoyamcnQ4NE/Or200m731cB/hZVBw6AAHK
xux2+sEmfmi2zZsxzggUq0lHPl6ljlwRvQhfxGRS22ep/n2dixikrpQcwmlX+ApS
z6HO+T5I1+3+eL4ImHp5NHUB7LBwW8KbAX/r7usQ60v+QePUBbGUYoB0ZKi71Pc4
MAzE5TN7O/XL2gmONwAZgCvUdmqWV3NZKWAKzKL0v26yhu6BKn8rxmyjOGtnWpz7
lXUSsI8pvJxPZJg9vDcPgnRaYE9lnr5uWZbGgMrvnKp9ZfqfcAyk3xrgfMwhLd0l
xNdYP50fC6Y2fGy3VsbcoPpSEnzNm/h4iObHmWvPoVfzFe4jbKi/aq5FywvPDBjT
Uhe45XAaeKv5BnrNP08XoVjrwcSMLxAYXAFyiSxiy4/PANuw1uHGRfPoGco7++kH
CrT0O4lItu+jkWljoI2IseFi2eA6W6iauWPWHb1UgwdbD+AKpWPU99Q1IvVDm3OL
+Ekqb8EdC/VxSCPr3n1aFz0anozHa6WlHnOHrVxIkKo/AVOlo/qKOid31r1acuqJ
YzfJ13tpFeQVv5586HaHxTxAfe2SBwu/6M8NUKv7TxV/ft9aH4pYjM51JeqV0Pyr
XxH90b43s9qdcDaPB7XKCPlBiVeCug8yck5kxWSQCRu6KUnFa04iH116stDICQal
3swNpghH66Oi0GgWVswCEjgrgkUzvu0HtVjn0b4CKFSMhWuld76z8sFfQqguIz6/
U6i3F6EikAE8Ve99F2Nkv84/iWBHgP0JwTT+q789ELnKSAEZzS4AVyByVXasSyDi
ePWY5KaZ4v9y/iy/R5f72ZFWZjwOIQSVqAdTpxtwqPo73Qv9m3wFVAodoVMRYnbB
gKLN72gIAc+UMW00d8e+eH3ZSqZRvZOCh8bR3qfDXGarYrRgRKvVfmMwxbuqcIeE
K00DZvb2uKScTNxXcnV+JLUaUMSCVWs1kWN+USCoYsphmP3qA47sj6wyZk9qnBQc
Fkr9LT5H5bvgqSV2wp4CxvL4PEPRr3s06x52AF9UxOfxIT8R7UwQIl/pQEXaMuKm
94a1m+QyP3TWODfj+GWeJbKajt+270cvgJQIHQ9XBZafDq+USS8GwOlPByz+fuqO
MSnY+bySG3ntqFa3WVjFVHbDFt15RffYyoJmM4G4XZN2TW3s3s1cUY0iHwb9cEHa
uMl2T9nDsTgPrqNypyI6f00ZK5nWSOYOpa4DbG4oRyK2Dptw5qGHMBaQVcsnJydb
04s8l8g42E66MKhx1WNNjRG7n3ML/Nth9tnmDHt+2TcMomZwccn+j88xOXSByQtZ
dDh7R05MI4fmLoDPTI8W8ah221kLtpa9U02xHiNH+WUmZ/nMc1ehDeP2NzW8XUtH
eoFJ1QuuqaFs0OxXt09h9ZpIUko4Z3YcBDPa//KNKbxjBze4DorRzfYUU5F4VMgO
cw1HZeb/Az0qN3RWOlKlhGQzd/4C1EbucbFGryU3XQALph0+wrY3DopoZ47ukaIt
nuZHGA+SD4DOCt6jhAUgP5EUFWUC4Z94TZat8puuGsRLeYJ0XslELe8lRExM55t/
H6GdZjB0P5g7L2Fc+on0Dl3yBu9dv+6JnQAMz8rj908SFYnWrOT4idI7b7g7f8wy
uF38F6F1drbXtTEDkZkyej655IWkILPs6o5w1Wc60Qw9oT/kUDIAWIjoNFeBic+w
w8Zih6g4tRCJbJDHQdN9+8shQqFa+Wz1QLovnXG20R1YJIh4LsFUThPpsl0N6VGU
wtUHlHhGW8IAWBedyjeCvHvpOG8raqoqaO3IQ9OCK3kkjz5RBBPhlXH9KjkGSwON
0uT2haYcKrr/GeUybcJOZ1lFb8uutqSa+Yz84vd9ZD8RQ2qqbCcxOplHqYPfQKT/
+MTqaiTAoJoLlI9p8NpTwng+MmDI5AZs8qWL71oX771fNV1I3rW4MSAJhovBgxzz
v5mo6amQc82XTQF5qS57C2iAbwEFG4n65VMoolsTaz17INpzf8VXcZAdhf3x0rni
DwKC0dXPjHzhgYDl3XF+G+CkBQFSU8t+C2NfpwJbD6EyZXOQKAkWWlZiGgA/pC/m
hW82xseVkI5EN0L9BcItWLfijAQJ6AfVCCOR+Y7D8trYHa6EGtyOmOo9AlAmqBIB
V+D1Sxsj2TGI4d2rIFCuQ0jpQDGV0/ad/WPY6+aGDknevGFSLGMe1ov0hDpjgYN/
YLQsvMvqSM3C1UkOVY+hKUFRGQ1LL9nG7+udfBr4VRN52x4iy8I8lnRNDtCqDBNg
tt0JrRVv3uzbh6pDbfF3tSPT7zGZ+b8ZXN+VU3AoszJ/sq/osImSyYjWFh3Nku7r
51lSHYreInpkvJfiLcW4/IAXi39uiupWdbsBN+Sd2NA0QF846J8n67bX2fD2hODH
+aDxFgH72fgYC0q1BwggC8TQgF/xUaQIDm6D6hJyVVyXuMRT9Eb8prp5mWo6wS98
KvgI1x27vSLIJtytlwEM1tmSprBARV5aCQy9J7bKt1rKZjnijLwcS3MdH43cv7AJ
k8712hIz5xz3F7Ru9IhBl5DDR1TZBpKc0D4iZmWe9wBhcmlXgbaW5H31A/rcwJtG
3C3cRhBwSY0OoMS3K/mgWlQLZLw1WpN2Ir0c1YIgn47hLTJhxHW+SrzxpgIYPuDb
iKOd4Cgj8CKLX09JRzPizMxebCLjMUu6hJwCCw+KfChtjzHSAEi7WqqBCLaXTOdR
0/RaXj1EqpUkCKf6rOD8etxTA+PULsV/iPORyOqp37u6oBhut4mGWEdjgNFNwAEr
Q+top6AOcAF/hly8t0HxzdIhksmNLha45R8KaEQTRa8zTAPo1TFM/BDmpTlQqPiU
ddq4d/eyaT+M5WJ5mwuqi5fwQ18z5qKyCJImIJdf9hsvz5svh1APQ3CJaYC2N3sC
7ZzANdMw48/+fIcR73zYQa36BMcRjq65HcOlPqGtjDhlMhp47RgTGTjN5lcgTktu
ybq44taCiRzmKlvFiMLjH6OByJkXMMirlXdR/blvjTFEmtkw7t72Xja7dEjmJrM8
fwyItyAs4ka8e9ImPYUjrDf0fjZjN9HsQbJ90BQl2juEVA362XMJAOqdDKtvztIA
eg+fG7RZqlPCf7G7AOxZ8ox3GWfo9t3CxKVZp9ZtLNDGSGOfbnwz++SrkfgG7Y/S
18+w39l88eYDPuBtvr/4NTuV2AFCSYEth0N72zjtPNmN58lcB8jfgjAd1nF7RDjZ
KD025FKi4kkJu6rrBEE0RR47nuuNo6OWIbOPc1MxjmK6HEDLuvbtXoz+tvGyXPqH
BFvjv83GrcUkvUaEfp2XJSYIT76dGYNMx5vFszkDDI+QgwmH8P1tgOHvLZMTGAYi
PAWhWqhub//xM/tHAYCmyIwljHJzDAEKEAIuhx3rKPiK0ByBY7o1JQZxykj8XFFr
X472fB9kYWoTYdm4HeXB1xztIi0+CDYScf3Yap5O3YW5u3zJB9Q+mE0Kv2gBFSk8
o2mhtWectNyACeKCTLNJFThSkk48voyzjriAj9ZL1oz/GSr11cIVtkGkan6wBzOm
+r5Y3gx0pvLIcoaa0FX3ohHSd6SK1+EbHX9f3FmZ4/MLkYKNfxWDzfT6PQ66knz2
lUtsRmQuvcoNkDGZikpEwWHxtw9kQwUxqoT12Fx3G7zrJnZH1nRIM9e7WTs91meM
+/6XBPfzaFfZC9F1Ranys9PpBkX3Ex3IOshs0tNlE9907lI/nR9jcH2kl+/dhE1b
BFfVLrI4fWNFQlTL/lh2S8fGJ9jr1hMUJi5fI26sPvsPxYjNdE4flldc9jDIEMkZ
BwVqVxWTOx7f8RH56avErkodWYbt6fZdiel9ycH1PdvdH8KhTbakRDhtsW4Nfe3B
diH1UlVk55eO+oM0rRNGSei2Ing3qZIJGXCPvE0Mm+ItHUkO+/PiPB3ocIs4hnlO
hrY3FughSoQGLyxXXE8bc/ubbdYQMQClsGhJR3QRBY7xtpe6IrzuNkKRi+Wug2XZ
Ljzqcs6zWZkALOtaQJU4fPuawrGJQ6Y0ga7r8HmsBm5eI6et1iaix5BsBnJWLTJP
WWjKRi6DzMqq4GBnXD2lIv5HOacO7NqmivaSrQsT3pHFZqv5zH7gDrA9HPt42pHD
GFe8duIOBJiI2wL0lDditQTTsTGyDgDIpayVoLS3Ta/qfP8rPTvP4MzZWa+iECvG
u55Mlj02/UrcI4A3YlwEUnDHKBbrMVcUY8Q8ggOXYKLQIcwtL61lgUQ3tV0HQWq3
mbwQjpa1L5uFSXAzNLf1O4/D52WteON46IwUlglHCOg3tDD9SNIbyLYYbxQZ5kAe
N5rWoHcOz9UWirkS4I3jbBJNdaWtNXGji4N7bbxER54o+pjgUtn7vhmNGdFxe6Kt
ORZ+OSyZAHNRXonm8TZ7d3GWXJvFkxM06Jy15e3zcu7z7eIAvHVRb3HZ6a9UHxKL
/lrIzka8xv3egKARpOcYUbD0Cb/m/2kmLDxUcwhuzYv5oMmXECPG2fFTad1Wey4N
SbQLdkX0sQzScGO4gN+/CVVpN5iqQ5K15n2naMD19Cyt8LskBRWjKUz6iligTYJk
2iQmNa6lf5l+I/mICyoK4WL8yezEbzl5GuMnuTD1huEspi2XD7zr9Jp+7GFly+6B
k1ZUs7JyDQsAFp3edD0twM9U7FmiKfrixl7AMiGmFqzD771bbss3BYOpOzJdxO4A
Eyjsr8hnW//sa+joFybODBArUToa3O9XzRkYT0o4kJRGflWqAXBKmfhXuT1ISaAR
f43S2NbHoizEofo16KS30ABN6FKJ0O2hbY05DkpBh+KkXE4BSOUZpMD9y3KazHHD
3YgIo72wY2FKN1ovfnWHrIK/gsb1D+gpqol/FBuqz0N/Wcs02BOB8dvRtwRorfI3
mCLB5PZcLDSgXPwYGmGcp1F1ZoEpOBjpyUpuDBUyQNClDvov1u02KPEzITHVHbG9
xe8Un+UpPEyflhAz6REQ8gwSPDwUhlWyZaCr9SYDYZVUmZZCgPgwiA8sNYAmt1LM
s7HbNQgl58SCYu6x6mquT886rF5d3E4XqLMeqTRfU7z/lcaTfqAJSw9VKzdAnQO2
tsHrI48BIvOP85VVDHn8nB0AqXfu6HtiErumE2u38bDgN7JaUvEagxXysX6vtHX/
3nyJDYtGo5hgq+8PRz0ISTFuMO4+ad9J0J1Ah+BYlI8YWYqZyo4CD7ylLV7Atpsz
DbZr//ZCs3dToGxWcsfdSjPwhfmmf2vaFXpHtzBiNjIWGT6OrA1krfqitGV1blcq
JVAl6l3Hwm2noaAjTp0visS/vwQ1UsZph6Hf/QVQ9tN/VGOhm+9Q1ZZ88+L0GdVM
65VQi8gtGyDkGTSnHElqVKrTljk+bPhXrCyqMPfur6Cssob7Hac7rigw3LwOJFQu
AYOsRk2YVjYMRN5M6rgKI+JsjSgKJ4WyOxk+ZN7VxtYRTJn3BGu2IWLxORzp/vHb
54cEXQb3fiXAAkmaifMPDqsMCg+mtKPjWcHdMRwAgoJf7tbY9fAWN2zZ9W3taRet
3dFPqCs97Qb1U86yy+H1c0L7RXERWYCLXiD52Aao7aOXWwPXqrKl3gSKxaoLhu/j
STEyUNzub1Ngtc1NQ14g0JKtF3k1Qp3+hC2+neZCYPYsUN+6QdNMAPaxKDtAqOdL
U5XsPAZVL64iDAewQ2TzGDEgym0hM22W95cb6vrqASKtP5MGsRFmTsrI/UHbDFKg
N0hOgczkF8cFLiIBqN0EMvQeGR+9+hDbkTIpHvOxAu7inPbmmlgDuOePrGYQ7Lkm
AWA8Dx2xe4ive21oH39iy4r47McQ1aBhAHvAiEV9akaIwiQFvPsLNSKX5atL7YPH
kn3aTQrxPGPYrFtDKJZxHpIMlkLTHxJSPhkx4EpAAYdicqfXFCDPWq3l5NaeTlKN
n8beKo84x78uPsYbNEvs2F9TzsMC5e1utLeu3f9q/07DCtW8XihOV80cTk8r3mvD
Im43A1AoqTDnh9j/mhYBN3D7tYCSIBS3JzI/LndRSVcf7Byg3rihm/X1i0Mj7CFP
C+DdYpysGegO1FSYE45iNaI16oqEDFJ7Yh/Cr8sjGzYN7oKbEmmOus/KiYKGziwD
Gp1VCEG3YXzOPnuuJt/hAX/DQzY0CT3k5GHSrmk4YDlGGXwYND/we5HLi0frkggu
s9TNXohg4gbdaJpzcJ5HS5eHf2z1/tBDHcUuGm5M4NC5zsSeKu59HbFCDNYUD93K
dow/v7Axkqk3MrDC13fUjiZbrk84O1vX/Y4dc622ntt2T5ntxIlbeG2jo+nhVr+x
JVpF6F9kWZWkLuGdIY3mDkF0kWCDrxoED2tMZfY2eHLbiro73iNCg0y20DXa2k57
YULZ0edA3400xCTlOlMoAlS+C3D7qDhoSFL9EzhhtwPSw1bMBPklmBvdAU+nA89X
rM8kQ8tBjmX2pBCH3RCdvwNZxYSxyKJY/UFM8cmMOThLdzImGKByoZZ6oGKJ+Blk
pTi5wgIwb+svNpLMGfi2psstIz/om+MVr8ZPsu1O3wDSa9S0Gmxa35JZfXVj0AAb
BaBiUPS3D23ITzuNqEyRrbYk5vr5v3jaZVqd8NlhcJT/K1OcYjFX9y6xEsVfFY98
Y33mqgVMv73e9h+++AwsE3hsj9zufh2lbxqcnPVaKcQZiHozhUGosJ957X9XOe93
UW39kiwiHpfWDLI0ceykQVMHoC/Vbh4N44GER7xsS6wkuTM0nAgaXRamp1ov/Gfu
XMx2RhWRnB9Jcv8vGq1TpHTkN/owIla4BnTRzViMOarV5R3yhNH4bXz7dWxist2o
frtvzMZH/IUgD/p87LJYTEAJPXJ43N9zRqxGObCUjqAMv9sFdbtGajh6h7xko+NX
PYeX1P8TUhrjsYWDbmCcHmB4ksZFajJ+hoinF7xPxYA92ggxCbLkmMatKgymCkca
3eJkMhADFxbzdsOB30gbv6P4xdjOT6uwXA3DCgRC4KsYOaPQubHNwXVjFQ+e6me/
1zmg4FIoqjAs/TwPLuwpJKhnYwzORCd+lEtZ7m0LzCbaO8VpdVToVu30rdNqiTd6
66UlA41TY8LDeStmlYfAskFpLCjp9P1pZPxKo4LYuWHLAUp71pkhlRtr2PgtwjOO
DvOqo/iihad2b26g5pzLH8iHreF5b5vh6fWQrXY478EpGwyvlZWde/TXN3VEhEg7
U0noL/SQVTFpRUWpmgvSWHC8OWU1RT4z2psGO2l5+z4JKbu/x+NrMYbKFiMr0Tpa
05ICb7qGHzyJPLkiSbc29glJpeQNU4eOf6MLZhuB2IWmb4890Qg5mu8s8G5cVaYH
D3fDfApxqXV217q2+XmDXHNOv3f1+6/OyQlaVbXDIJgkt/Zkh/pAM6QgFgB3Tk7/
BB9HwEQgbfNDAE3Hgm12s57CEFEonAnQmKLJ5+GjLEc/NhNjbmGAde53Hq6StWBw
x3snwc4dO1ThDBr+hWcMG9qi7zl7FuL6Ag2jqvfgKwnDEz6gsHZV+6yhJLmKG0zA
69KAMltEa2j/gwY8OOKNHlqlbeYE1e6a1bZYQgfOAbLR0Vxtu5QWy3jPEyzCI/om
wBY8oKFXjQL+wstXWoeckTJ5Qw1Ip2va6YtiPExaIU+5+l1JiwIBR5BTnZQrbvPQ
9WpfNMS2vwdPvi7VKL+pV0Z+aj9KIja6Pax7Hq5FVkmNRCwV51viiAGz9xrw+VfP
A9JvRGcpXMT4mvY1i5Rdy1h89qgiDq02gE7szYxuUywC0bDZCPNYG21UPZFp0IJV
4ZnBr2PTgE/sXVt6NS0CXIbaXDaWfTLYONlnAHaksrJuxa0WfKBeC5FgS8DHrVfW
xd3omJDY0aUqNGzZ6YajU8FHAN8AnX4nVZA9Y2v5/cIRKRNKTAUj29x+xWIjyHUT
rLKdDwtmodsXr8zg2lRcbp/wxr26aAQlKgF+6TeD+lOBe7Fobbl8U2cdNR0wa1F/
AEZdsnZkgaQdbmgDo9JUcG7LukeYmFkAZXA8s8Lkk52OGgmARkRDIKTnMjIfhnYn
UuYIelRDxPgyqmMWevTgSco7STUNRA/7ccjf6UJx0jfUngjRY0zl8MZX//ddHEUA
uR5YwZKITgY/gfTdrpyHH3M8yecvPbrqIaY+9H7iJslgBoizVfrQcWpLh5MAohyE
yhb3/LYXPDnF09C85OFz9bd6qmP/RSOhLBDYEkCGLbKU9cGfmm7ZUCbbkycXyxFW
WQMvvVMDQOAHODN6kRwqbjVODw+HmqYR7c7UCw4nVQ8zQEy2HtQCBCktIkd9/S+L
I0P9GTw7rs5134aQcYKLvwDYQYUUmY56rTxqK4UqQ6AWOxfiIoSUhcM/CI0y0jnr
sDB3ePn0pzXBbqLSu4d9F9qQhx94CaweqcCb6DFwF6H9ts8HU9v63gaMpmxxw7e0
6Yw8+FceZNR/faERX8GuwhxlDkFcZb3n8KOq5jrWGWLG6OKBUCKKHfSBv9be8CUq
GBV27mq7ZVs8WgOy43vKaULbggB3YFBNDfPTBPZDcX2dy+gh/XscfD01vZgKXW+V
VQI6prtob/CDK0s8Bj+kClGAgIthetNaMX2ofTDWC3UkXOJm7kCl0sGngqWgaArk
QiGipjtLSeSBPG1fKwb0ZBE+fxgtVoHIoHPSC51SmMuG8v2eQXpJdT2d30tHAZ0T
kJathv6CgBN0/ICFif+yBXHgOXsII2IZOOCjnBdtQos9te7wkB+sZNU1xPgRFW0y
bZnf8N61dfxux8ce59VbfMaux8cGRBTnzb8zBiqikpqKVWSaGnm/L/6Q/MyuXg7D
9GejpXOXnAH2Q0RJaYKrXrRs6NzEou1TPlgRS+hFGzMqZsUQ7mur4l2eqFHvO02Y
WrFfPV4Pg0nk+r7IPmOBuE8nDak7kKdbLgbyUd/1t13DqbjlTuOg9/BWQtCAkB3L
pjCB2HejpuH74Cml4aKow0rX15wp/ffWzmTvmrVmtWacgw2HiPZMvP8C+9dDkcnb
c/1DtIHGVTERz/xm8VfwJ6eyZ3cxDFOQ3qulQg/GDSIh8J8atJ0eBG3cMx8dkPAp
9SHeB1Rs5YU1FcCZQOVq1IokmRya3OykX8+0MiNvpRRmpWAL59/36l3sZ//cXT+J
WlKPyw9mEgnph3+Bn7sEyi4Fqc2itGatjIUt7eCsTLA0LsMndLauNcdkp2B7Er3k
7Hm4sLzzAEzWRBZDveGHKOVwwR0XOuaX+9AeeiSlCOpir5XYTCKa6dJHZbYdGJLo
bg5hnsJk19FB4PrautE3h31lVkRxXZJZk7T2BZIqAervPch3TpSHtbmiQzEslTsU
VenRLYkqbxLxakceArywr2n2H8GLYN6q3i93lxAT8Wfr4DfjsUqS1eC9qcDKJM0u
HV2d9ioSCjXhvMeCSsezB2drcmKctEBCJXkI9zuiQEdz4rxLhz1oaPcrvu++LoA+
asVCRUYgqKvrBr9Wo/XBL31FKB8y6LD2zvGAoxsu7LZiQrnPMFWj5eryPXc5l3nB
FCD8i0uQwH/qEToUIvzibfEBkq3tTW0COoXO/0A6dz5uG0d5JZ3s4Z0cB6bUaVmP
+IylqOYdpxlJ2S/M6k4odaLfsgJmRpsFnp76IEMpuOrfAghRkXr6oZqTcZW0/RAL
AgzzElRKZj67w7QuzdDH8XGVJTBVXL2e8ucPcvV5r8lGtKm+/gd0eRivkL9git7G
xXgXNq9PrDa28TpNQXT4j/1kJumBITpcJjZFTeRqrcdk0o+GJZqEocFUpZLpq5IF
zFs9kw2HhKi5LvCCYgVKkL30tXbHmTH7KHet2qwm3e697hrsuVzG599ezyojt/lr
BvQdk01tefxOrzPJGfx/240HsCgjWi9n1ObN8MUcUv7Cotw4wYsN0FAKsTF+8Azg
O3IndC6Vj3f36sAynnfrH6YXmU+iMugqXjQ+fhbQRsD8e6hGJf4tdtIJxc+V2TwE
U+wVMs32K/psbduV/DQc1+9Ct1dbjLXUxy63DZ2kpRSt9waH8DxdgVxcg+1Tr5SS
lLhzJugwypdtzf44xBfEuY/GPtCYEanSjpBDskmVLVMwkrIw3wQmcoDaW82lhTBW
5Yo2XjjHwhuAFDliAyi+3gPV2pFFdlaIeiAU3KQHfWYY3BHjzUb2U+d1Jajma75w
4uudwTj5Aq0YTmjEFfH4visZB2oskfCR8dFz/+GTqEGbKSfOCySR3I6hAOQDoWkD
bgJQA/HoWDEuc1wBvlym8/efwUL/3bmr5IaB1NQsxK2vXosJEhjRnJfnkhAWZNyx
4k9/ewykKO8J/mzj3yj0W16o0FjhNGlrXbgVTcKWrS5+VCDcse5sVCQObJ9hs+0l
YM/P1VPeIXbRe90wYQA+K5Dh7qs46yYgrAQYc/wyEYnK/KZzRWWh0t2tYdcEBYLY
W1QodX5d29GJchiIx5RGson0C1ixoRh2JKoGALbrGtrhPenjXs6Z4Q994WMiU2e4
jjlGjOkI3WgwiUvd3ZeYcqmakiADSYuTdiiR8dizdYqVmVUtB3t5UBGP+/KVbXfU
g9foE+yCxiGY3QBPVhD0d97463gXdOYDDh1BZQqQnK/Efp/Cdg5ssJvbofgq6qWt
9rhXQ18dIC6QNsMQlsSuAGeVD0mft2/n25fTq/u1dgmq2UrNbO5wwbZUDig+KXAT
CIXyPK3VsyyMcSq009iid/kytyLjfJUPaOkahBwZyF82wKbNAK6HbxMCQADPvxdp
3YYel/eONA/Mlr7McadbfcG/YYl82LWm7q1TakDKwkcIJw3vcay/umtpnqZFtsdH
w3Z97u89+x4+045zcEQ7ssSLfuhPMNhCfsWJNXAwXlyn9sk1Crcmrrhe3we+upMM
WRaXFML86sbcd2yteZSS0zqpAGbQfbO5ggzpaj9V/NkPgNoq1UpYC9YBY54Tr99k
SZy+qWEal57ACa1jQL0LzQJJh2c66vVZxGYVu/p1IMkR6Hq6Gjn4Tu8NI0Qj23yt
zAmxOcqck7+N6HBvnV6y/c92oLgONYZ0KUwOENNRvNwuvaXYbDfRBVsJ5fvdI8wG
jhb7Z0FPrKNseY7OSIV9dB+SqFeS28kpkZzCuwz7X73bc/RdOcq02e6DM8cFD8dV
CfiV0fezU7s0yXwhibRu4BpokAj/EwCE82hqzSRmIDE4bCzcLy2VkhbhWah5ksVo
Z1/m+vAIp8i/of4T2t5CaxpATklBQJ7Wb55oAKX3ovvM0mV1SjuSKjcod7DNOO26
9LOrGiTDGrBy9Du5qWZdbai1c6g6fPPTcBkE2oq0VgFSpp+6QjVGwB3c7vM17XNi
U7toyyLlvwgfbdP+1kNV4i+7sAOyse4ON2zIuiUBksvHOlfMlaGBgJyDeuuyX0pK
8U+/1mCLxLeGjlpaH/xsyxnE/cM3Ta5jupRuZDNEmjZquXk3O8yh/qlrQjRPAzfw
/j2JVAGG0lLoGY2nV2b6/fqgKFtI2qMECdCCG1ddEPa8W7dVApK+eoFsSoEGs+Re
nQgY7qEkB5+sdta0LO2TkShmbkgv6oyfdQ4B94Oz7D8jsg4HT/5vEems1rWzZGXG
fKkzscktAKx6FdyfQHCUsjnw6cXZUs3vbgSNS6t5bLOH0/6IzqwH0JXPsW57QYrt
R7qUFbEEMiuLaQGr7ZoV8hAu3JKeBr8UnzcGhPZuSn0wfP9EoXmnF/ro7dRK5dEg
2A8uu9HT+1HElTmK62ClysH9e1ISDI/55qHum+GvgVN84EKhdOKC75O/BY903Xtg
xeoHDZcKDnJIPOLny3267jZsyD9JdbTwhu5TV1PSEalcjjSp5XoDdI344G1ke6n8
AO8RSyLstc2YVrPWfsXuvPzCJw8se6Uaz9YJ5J0yu3eahHR+QX6fJ/Gv2UhPFwFR
HgWxgkGyI4VaMgeCfKHvCmaU4KkYwFimjfdoOEJtX1V6Hf5z6ruWIHOlE9NoYcM+
1AwcCMaAh18qPIRcHx4o8bFj9uPS9jU7jdQF6rS9wxGltiNvKAZ0BV97ksXN1JkN
jN2njhf6t1ArJF8n0674cmYwN1Yi4d4ZuFyZPPKSE1yq5+TEUQdfsGBEtH1benH+
uy5W+pPaU8Vanul5WZ3ndOC3F9PR44+VFEx/wd6kc9E6xfLK8VF4wB92g/SNoImc
1E2x+rsshLVS4zhMLSAICtT/z98irh+Wxd5ODEwRc2pnEls96f135+AYG3NTtGDl
utLuzOz8o0DaUVs1E7MSy8PNdkVn+LfTWgthH4uYsQPVqVfYMkwUlGhmoi/JG4XW
2Jy0KN2POyuf4zOej4bnX9r2LTdeLIH9rWhUOYKE4dgxNCsEier8TcCUX4MQxrQL
ZfyRgP3F0KplTcvfLbmF6QMgkfsFvib+RHeKW3TRvw9GW16gOwWZjx8Crx/VBIh2
RCPcpx6jFBhLmxKx+CZ0TQglENm0xUvZN6AFke3WqYBwNuCSJeWYymxlGsgYt72j
u1VVn7UUcCeq6I2i8q4hYQ7557aZc8+EU3EnfNop92JXf584qt/3w0yDTSp5/MYE
OCcdDk7wZTMdBH79sfebHEI54rcgDlK8nqy1R/aqxwypv+BfcwRjnXh7EFCv2hNa
4mezP4Mx46LBY8Q0nJYBgIQIVHfSMoMgRZBqlvaGliS5pCBy8C7GmLVLNTRcIXRt
NyZT6Pb+nXary2dtb8+OGRSlalSwdVc/jL5NisE5kXc8SV2wglBp/PN/IDj6XlD6
hvLDye0Gq/EUAGk01Ahs1qrT00Ycxvy4KKg974F+f670tLS2GXuDTtWUaVFt4HrO
8OLHG/dHFqF6y+C1/K7xzbEwtZXxrJMioSCaxVpv+q3W/1yScmMC/F8RvwWeG9cI
DJ9D/g63U9Nev+C7dNxXqs82wnfxqQgjFknljGaz1kQD3ci6noXoxGWWNNqeZZr/
I4zytSiKJr9txGPIrikEnXWiUM7qxeU8mh0rqbNoR48TzoomMdWMBBOloRPN+Ebp
lVooF3Z2w0/R67kJq+qO7+/dtECXGwSFvYwZMwZMKl8cc9y4gPdeyvnTgI3IcDpj
VJvMbWTepX+qYdcxrpUcQfXm3GU1/v7jnNyb4JrSlzauNpdpKzaMMRuNI0mfBq1W
5PFpLMvHZWgnno97mL7S8fDgu5PEZ3cYW1/uQkxxFA/N6Yu40kzlZlunN2/Ca82q
xuMSKh7XEc7u70ji+TtQQUejKRUcPRR9D9m+rUv5TsmiFy6IUFbVfyAtRYqRJL3q
k1/BQ0Qq4v7Qb9EPZoqvDGoLYwpNhTqem64h4HZMQ3yv9R34534CsaFZw7lelA6c
6SQpeuCwZ6iEHNi8T98qESzhMfo/T0PlY1N0BABDcREnPu63e0hnBs60yXlOzpZn
s4cTTIjn6yLUzWMBCjNSg3yfjIGmt4NgwpyJaDKRDiLswt+co2s3hpjiG01wZRNW
VvVbkjqZT90sUhpuVp+FoWnBooRtoQ6p+k2qQFrw4MMWy9Z0GFuEMdk92dqgX2jf
sWpgOpDmBTbYjfJ+FC/PpVPxvuPNNZZQPF3Z11U1ahkgEi2WsbT1HzXp0PMVR2aO
AimzB6qlFm/AEHE80oc9T58Z5PNfS2h1QzqnQoaVyN5cTRwgcfLB/6BgFHSV4hH6
dPfBTLalL/5/C7iU+u4+slLXu5XNfF4sWoi42EUnT8oBslgp+SWKNg76bvDXKb+w
IeLGVK4L7X/7X4LE9GpOk0DeblyVMhsEqnPR2csVUUQmA1cBy90MeLeNv9lCfj5r
g4s+teEY5rXMVt4YdTWZOHmBgDaTooSXl4H4q22zONcwUgRum2vZGEaeqnrIGL/L
MK3DzziEOmiHnOGco7Y+woEm6JdqEci+NHgzE5zKIbI4rCF7BG904xi7gh1a51M0
vAJOTAHJVSmNfh3vHeD33kUjwm/ELB6p1AUz3KyarvhGIWgwHQCQQlRD0QXoCGud
4ggVLN3F0bTkz6YyaL9pZgp86XoVmDEQJIxnTPPDT8dGbpGeGoXfLYorFB7p8nQc
XKGSb2yNwFbIihD3B1YbuC6LFLbozheGUL2RWj+/XPBGGNSWXninqnFELtYE35+b
lwT5p9toIDJg1ImEAZlHUoWkHV2nN57NGMd83/Hhn1H09MlAiVH8kbgeZKS0Qo2A
0BtZNyQEhhYHrUbF3MuucA87GQsRZbihxSPndrYEph1/zD1L0Zby0Ph2TudSND+h
AQ+m7XPwvEIEvX9RY/fRIVTU7ybk5Zav8OIDpfPZY6NZtXaheLMkT9joL72os9IJ
oBXqCVnc915gYgYaEyye0DWWFcHaBb7c9DE8e6rnyMVk1sj7pxaqNfPuSRtzv0uV
mDkgl8g02A7x9NDI2eAlMX4voXktlXbaTiu5d26bHOf9v0dfdq4sETqGtjwarXLR
8XBAMQYBASA0TH4Ql8YU5YNOyo4+RscMeOikML7XzFcXUbrjf5+wS58szrIq2sK9
5308WxxkWHnYJ0MDTPI3XoKD7AyEtP7zi9PfEz8lEYKjGhFp6SiL9a6hS94AlYd1
zUicHPvPrMogDt7Fz7t77dM3bWz7/BrRejhg+DNbEQY9sNpNmrNa6HS2BlUkc8HY
AAdBfcn0Ulg/xQgkAnIPN22t4VJ1+upBfjy9dj/tgtwB/43EGiju45/jSCyudg5i
bjWKtVHOvilrN1MjYA7tL9h4w3LBvMmgKJ/XAQyNyHx94Xjm0z7T8FmZgb7GfK/x
MAkGWTElpPHQs6BcDaPtVUAZDIW2ipBUq5UJfyVt2wWZGwvX4tOBTuOfv5rH+N8r
0XjOauJBVPM5XgEQPRNw39VWW0JFm0SPPHhJOSz+4JXySoxqUqiz8ClGVVTVP/kM
sdR9CG/PAfIKJ5tTueUmfVz3BvfhvX5aWoKU/dM5TdR5d5+zUTWOSeersPEuvYaD
PUbmJmEpr2rJRg1ckje+VSJ6L6W5lrDCmcBuS0h9LD8hjpWFp5Pc6p0BxVx1PEk5
qlkpjyjSu4e7tXt1oOTI2ChD8nMHo27QdiPAf0nSoEkcpQ2kjkyHVqc1gCW4mtC1
qvfJMtHCfdNuyggGVp/ve+/jAMQFiJmXEKBAraJAMHflAY2dC1zjplbwRoDaiWQi
rqwSteEI+5/CLid0lihMXPliDA/2SNFx7OTgFcsRwke2w444BasUhM1CEbDk6U2f
K8ybQqLo89toXSMYaiEDykhx+drLyOh5lJhinOqY37chOwOc06eowZ1v5Xfjg1sk
pwy85pMdH+LUS/CiEryEi6UB8X+j0Xl4phRhunW+gKR66vc4bcsftvjgMMn9i6IF
5X0Y/IX/7ZaiOjudbG9PpnVz2HQW3yby+xtv8g34XoSLBzF29HXFcNtCGSE7zHSx
rE0yr62bZ2iSyOyov7rvJRwsyTqiETw2x810B+sepHy4P9li/Ajg3MuIhRln/h6i
LkIQFhefRsgXpgBisgdiEvgUMzU3IyGaEZ5mO1y3792BXxD0XQVybCARgYxDSsgi
c/7nXuHtwvF5agOLW2Ptr9gIfFVn7G1nKsA8SGS68lt1RaOOnTDyvEfUwJ6+3CoK
vg2vbd9A0tAJBVnhodnQq4+L8LV/MokAjLeIFvgTnrIbN4oG/uWfopPSDPv9Rzj4
KrODcdJwgzMR6knIvUZO9/wb9Qs8MLSQtf3HLRRg8XZomNExJk3TnggAy1WCumPp
bhoGSz9SRCg96V1i2fcZEXMUjvh/xD8ZGNU1IOnjc25QRyi69+HfnVZ7lU2t3NSK
MjMk6RA2v06Lvb6WfPIZr4vmpKvykFgDsWCXEwcrWyAj0qOU03ST0etEbVsVz8bT
AbRCf823tLLHFLc5Uah67II5JpUByYR70SPuXZ9azUkw40uWpcY6Bs7jDd+zCpxt
TEHNVjOCIRkw9L35Rfj3S+kleIKLtPEbGfGyZadecnTwU/vvIfpeJdTKGEnlsRIW
tA73KistYqewtnKnNn4CdXYOO1UUP+dhwhuYS1e3OMpP3frDjwax73lQ25/YBcza
3xQ3268ZELzkSbheGaZRxpmCZfI25XYPW/VWzCHZ6soUP4tF1hlShMj4RKRpV852
jWA9+22iNjAfoTY+9BrfOyG56PB9wRoaQSnfbfumuw55Ck/LkbPOP2Bgx2PX+41N
FJBLUXrxOqV4MKQTR5kW4gI4kpcPxGs/OhiUqGOCHdZDGGklv4Hcw1sBWKzxvRH3
iLu4jlkhClJ4czPLSOsmWeFTBaKi9iRppZCGsetP13h+xLuKfMp8Dn7z4c1/OYAI
d/FrczEN0faC/W3kOV42rm92xh5vpiHGtx/7sCqwqFqj9mDuvWk/vouLNoh6mttL
1QTz1yoL+eZ48ST86cUt2+stTgX5YvvQGKcHEEuYvHPrEKWgWwxLgOzhsm8z9rm1
vKWMAmw6GmuuEjlBa+YkYLVcKGyfArklEtn06r5OZdvcK6YUNI5NXxPQHM41BLGQ
Gk0sEvPaxXDlsFk5ZV9+aS03o0byv1O75A8L5385fVjixWbyxuTvGpl1qDjN08ia
Mj1H7kDYUPNxFUK9o3krR31iea5tydKikgA+fsAG1qfM2vdDQmHF96uzSj5E49tA
+h0Cl2u2AAnAV7ao7iCsMcym5bJTnPd4ZdvugvXbvOt8O09JsPy0W5b5e0l1jU1/
QBUoEjQUuaagf5K53BH2cvLbuMvYi1CVefvvp2s/JvMEXc2Up/SGygpkMfRPxtw0
9tJASAFAxzELLzOAf/cBFNDkpwkQ8ZwM80z5RjItdNRgvMXuZShGLNl5MKgLpbNk
Vs7x7HCXVGR3Xkl81j/vFNqROwyEIPd2GCZsfxbssouKedOlxUsbOwC6YrSB7bRL
lSXHDxWWWhnpGR+clgsaD2nnQ0uQeubWzOQAJZZoES/XpG0mWB9IoIYT2peFkO9k
t8/LyfmlsE86L9aEOkaGFPo277jRmJvF64B3H5xgI4gFpetqjJucu/McoVAUUmEY
q956Td7XVnqCdoM/P4Bvqx+RBzOR0SBLTPQZ6zKdfg3+jYbc4ADbnrznQHWiOPZk
QZYWdrCfLsAWV0vCJImhV6SWMZaFXiBDFcHeSDgtNIjzbs6EJ8N93IaJnOf2xezO
uG8piy90B8OJ9ldRuOQfqNzVjTjX/Errwr8Yjg9Ei/sbGUaea26tXv3isrntK3iK
m0GVDl0tXyAbLmtsvYhMGwgzYMK0295zEWNllAINeMBygCKXPU/JrTw3i8JOACQP
T1tMpjgQ1jNBYhRZhhGQFkUVSVTBQyRJCaaYgaUP1yJL5lnkmAc70t8zORblUwSB
9yq3bx6AUUjqS9bhWh0vmxg7N6cToY31eXVwJ3fYScwUNOc+3Akugk0+zUW+SEP1
4vbxVTHFMvZNvIhT7EIZZHcPQQXMoIk4VHlbKi0l0U/8BAXV4Yb7KzcNpuejNK4O
L7Tp/Pypjuz977PYlWd8rQvCLKQepddl7t/ig0sSsLpx7YbU3Rc07Bd5ygZbpPW5
WFWxs6+bo1b2dkG92NO+j3oHpe80X0mMFpDv9W5tRN7ZdQU+0cia22ZunHornDke
3Eo5EF2ZfZxXV1vbayKPylmWKX5AmjFFwnIlkhOrCw7oJaJHzAzG3QMdu0YVzYEb
BTfZk/7CkOEv/zzuhlcid2c7H+bZG5/M9I9wCtKfMD8NPf60tGoyUBt10sYhsSk4
3XL8Z8T8RZAA/EHHvKn16fDt4yNXs5+6/E52G5hPqAW1YIwDHj5kU/XoTwUmaHS5
yF8KxKsKsN4E6/yAbOXJaS6rHfAkmQknHCFfjLt360hKuVocxjW7D9dWywBAwm9I
f4Hpu37Am2GoOjjldXdg8lywSvYc3l9WpCq77R8lsK/+fiMAGOwjeANAg+VrSy6n
Ym9znECETwqvKMNf4xg+Hr49SUW6ZmIX33JlLCSky8+isU2hqs1UZntthW3tfVcQ
JenKw9L1weJPLfhY0XrAmcHlKZCSHjJUOEl9cwVd3Ew4IAe0cfZbCou5ZR3KFOjK
GiOB20KGn8iW1N2EktJqXSTYIeA1O3fBtH2WkfrQxIcx+QVkbl/CqNR1+wW3e8oz
0JGo8UqDPryFhUVMFZ2C9aDG+GL2FecQc3aortGxKVghAoWEKNc80dTstwwWUJNU
AsCbJHM72vRhfoRCVTQMFt6bZOHyo0Nv67VcCc2H7LYTjw5iAKgJ+dL8nXvRkDVd
kqTkd00yqqQXZ95lxoJyGTXStWlrnc6Mo6R5SSph5genOPs3JBcgxU5y+ThCwb8B
bKw9roAMj6Se6CjhXw95uHrh/LiopyT2mWjz/xcBWw8rGvcBdEeueVCxIWXX38K6
KsUOjUUHrxwJ2XLCgHVGweJEYlMH5kLt9jjGHh1VqQuiFgmcB3NiHDrt/k4Ras32
HCcMhQC+aUIr5yyoh+55bSDhKQ/xn+v/0z7QednoFmF4ekklD8vlyUcBoazJRKa0
Gx+L8OTJinht1GBNV2Wesli2zuNGPSnmGZu0DpWqasmUJfoZHTfCyiJ4ZZkFgXuA
tcwIgk0O+cnhT1wLEajKzGHaY32Wk9nktg9j6XYcFPzRP81yc6tpEmLO7Oson5ku
770YdhSpR/YC3jJ4WlT+jeg739xuARzZ6MkN57munqRHVLBUlXsfrV5q6J61wVpI
loHd4KfNzcnAhfnsJVmkxn27ufJ8oyoosenV8Z8I3LJonkLRqqwzThhmBUO0I1it
DtIsopIZFwYEkFuYXALqWmECm4iXpGrVhm5qyt4ZG8XG/V7dvUZ5g8DNwRbQIxQP
AcFhCIPVnKgWJmenh4dfkyP5pAIRmwHeSqSzaGTtmMnlBgPzPDUuPK8t61rgH85A
vVfB7Skbol7VRekk3xfzZz6ysjgZ0/KpQwGRqWJcXaWsFnQqEWlar5h1oxJLxEKt
bE9Yo6k9RmoanRAwLm9b+rkAlpH3zC3oPa2cKtTivO0otb2J50pjlDrgnv6jHKSK
hc9qgJkSdmn6zp0ZUccMD+IyBivnGfhUsPrpW840AySKnktaJ0yvjbDlI0hBN0CJ
/gnqpzmGfe7v2IkuVyV9StVn4LqhpOAYkvc1RAaSWueUw/iL5qAUAiuktJ7VuzUD
C1Q+j0dmdwj/pH+A5AfFPG2f+KX8BCePuThAeRCcBKPK3T+IyCLh+BT/aC3TrPV0
yn/KL1jqLCWPS2AVPyqzVl43WgXSYpCDLUBOLlWwTWN41j8z8qwGL/6ste1zhJQb
Yj+fnkW1XMuW6k9Qt0FPBP57WBRulJyGgPikhTXFWn0DNBr7J5VRR2VH+UDNVB0w
sjjv4vu8IL9YR4AdF5kOr02k5rJ7K+Ng/GX3ByP1oFDyyI+4pQbo+FJHJMGNA0Pq
C35wVBCIXDHeXWP0906SXwl20Xw8yWmVXLdVx5b9axn5uvstHZerArc8ep4kRieC
Sat/Hfl5uhAOHH9uSlJ4j6Bnwz4WOm/RBvkg+Xk5tl/cf+frq9Cdo6SZr8bLOKzL
1++GW2siCQB2OWah/D+aZ10u5u1DdYNTOnwwFodl5Ut0gYQVCQYradUDZVlmXWMy
Ze/CULZtkIF77uM05WLXLI4DrDhvwKVZ6S4robwTofbb+D8nG0z/cQ/pqho8EQ1S
jbgrEo89/cfK6oX+Cjanthc38zQkvvNSOZLTH390SSxJjvljuW68/nUmzYnWpO5w
elLB3wPLIz7oznkLRp/Qasa3wp6hIRm4lPMhn7IMMbZvkmrD1t3ShOtBMw2YHP2d
m6Tbu1chNd6LeHNlONBBlliSt0kMtCQrepp209+dAyKcLBqfRYipa/WthTyOFCgL
jRDvIAPsHF2Js6tHaEVp2fBcR/A2JdIEvsjm+I2WdmKoB7eTIDuXvJbM1sSg/9Ni
QKUUUhuwOcvpZSs88yEnfWmwzeX9nK0N80AAs3a/uddvq6H7wRxYwgbkRj8/2U61
qnjwk/D3dbI4Yl/cYAwDjhf1iyoDbG8Bsn7WxrtUluYgFNnW3SLS9nBOMkWgY7y9
DiB1GMquKDtIvG8972Tu0s6Df4VFTjtyCUIQ9PW/kjYzCV8MaBGgUAfnUnOwao8x
DLgHIFgQa9Dz2Zzrdrkc0ArmdiLnoBwTT3JYb+wCXLbHeAr+s442YxGUZptBHakQ
G4RptrxaCH4zU5cV45S52K26/wxMsrudm8QE7IFcoTPEAM52kunnvieqTzEPp3rW
vgWiDwdB3wE1YArNU3tkhyo5yPtZRjyCtOkLDn0c5KjfGj6sczoTvA/4yRUUA/D0
b95l6kQLCtIXamgUxO73+o7DLdZO3A3NLXhA3yDKV3Kv1AeGXQ9UTNDCMKMXbv8K
3RttkQQVu+3qoxEuO73HoSKZhF25qlVrgCD1rLas9PqCVAcOxTcw5XYVqqZ0SjuR
JxRWUlPGb/fi/cObkfl3GWYNHzls9KtZ/eQFcf9BbxHnHKVVTEMAXc159sVohXWb
ToZcPnESVAHbF99DrEgM45m6ZgS3g7jrLAoihjh8UKq6PRPDrLcYAmUNO7oxflT8
sTnl7ubXsRjFGsi29dvfpPggF6QS4gmFgjlI/wU0Bzjy+ugxVGvGgsIKwo1+9mIZ
Oy1LPqq5HlDitEHQF6tMY3IXGuN5AQ0dGyxbpk/B6MlEzUiTA2NlQcTCaOWlB2O1
xLTCkxtl+UmWjYqeYSl+e0dLacvztGVTuDIwhQQudp5Kg16lHdbs5J+E+lMj3Syb
SrkEQEcD9mx0G34F+flcF8UBonUYcEROnsae5ncd4K/EAasSMQ5dbt+nwk76NpTh
k5hnKKZu/+EeVi9H9FIUUs2yI+OrA0T3Y48bjzIEYJ0YzxQWKgAc9/oEeo5Lv010
rEh9GuleXAA6cQEKHOIWTc3JStbYXbaHSXaXgeU+TgtvtIcEgofVUoULxgn3/Brv
AmtRV1FEZu80tDQ32wBRMaeYx0XqjO6gwbg7Mqz9pwwC2O9xGIi1Z1uIFfYDkni+
gYdUYmlGZE1DBOO3yJS8262unJ2Wkg8LSKCDv8gdhxxWMyGcEJXMrSkNlS6tbk/2
R5EL+jCXJ+xnBdBRFxBEIjxG5feqvwRouDUSHF2CA1LEkDQlRp9zy7ADKd065Ock
OupnzNsI/PyevddW40FyL+nmL5hQ48C3oBs4z9Y5ShV/1m8ENWxaSpKxzE1PfQl6
6RDio5O0A0BVGusaddEWIYiGnc3AF9Jwn+MWP75XK4o9y20t3jUwDRwJaXQMNzJa
/ZHfkDw+bL+yBaAl3ZI1FsoTErG4JYr03P/gju9Y15zgVbTCYf4Rt08Tj6OF/63a
PL/uMYY27kKa/9Kw8eiahgwlq6fb9WOTU0BSbYO6qKZxAdKSFd0HoRN/sJEPEOXJ
VqAatte763jGDbg/sR0XPJPPgiDg4a1N+76fqnGW78eAir/6SXsgqQTts+LiSuBD
wVKqJjaw0ycqVmBXDqiIX7PLnWXHasTggK9ZgGr0BT8jhI3aphH4loE9oTjqXcJh
AMxdLOidhlnQFbz3zL2i7FvKLwSnb0lUbhkEloX0yWG7gd2yIkguxnZJQ+x8o1gG
kHol5+5+t7PMHAn6tarzEsahDbdPVR9ZrHMNHmPl3dfr9ese6UlUltuxDX7n2cjz
7rsPTwV0xv3ujnfqt1/Fz2sYd9ESzseL5lyL0KUj2ZrHFLKavdacOnNJIoUKo0tJ
nbsUmvmYmXXC0s3UpMWsYDgiw9Tg5KHYIMb0MD5hqqrmgXcaIvvDKcxKOqQ8Y5ec
z5tekHBuBFtAsYTu52seQnrpeRUxQdPzK0MhaSpSXzWXOHTyA3eH+40Bz4to6kXw
1RnVCGqE/94egE3JRiDNgWTx0R8E9gD7IneacSB642Z5EYIfeJ2S9Z4y6g9vJArC
2QRXvzp6sxNwZdV27RX/Vdwyb7OT6LBxPm2qnrd04IorfOZI/TWUgvSnARb+qUX9
NZNPCE7x0Hs8UmAvUbDjHSrCy4vZAkvq2QCR7SrdRRXNq2LTJ3eiPP2EdFAMdtwr
gTob8CtTkNxWC78G6Fo21QNrRZdI8xHu7a9LdXbit2RAa6uD61dTtdaVx0qSwoXa
Wk/JRLm+OQkge2fK/BI6+44/PsbHGWH0cGZSORqeA2cF/qgJPM2EcdYF/MbQCWUs
Bdu9c8reWWQrW486wGmgWewn+GpyXq6N/Qs3i2Dx8t+5WWqr+NGUmi954WaVxk1u
KAIHetJ0PdTFWryTPhEHV6avzffhVFMk6ry+4K5G+OpVNvvpi6iUiLA8ZhcUAh2E
ZCSEwbbvrYJZpeXBoqYbhYLD070hZ+BXe4nze5gOryF7kuA9Qvs/6ldZG+6kR0bg
wgpbjFM/19EhY/njgwmcfEzEgo5mX+YFf4ZuxQmvVKXtJkD77JYIlaJDsqtQBmKa
O7hti/IFNpBxN1KwcXKXJiwsU05PunfttctHg6Y8WvfPJzlYWHu7DfJPo6CmNeNE
1FVC2X2fUpBoHio9LSvdh1RERAUC254oj0ifGpyHGgfS0uS5a+5hvkKyrr5od9jG
RhZ3w5TZYlU0d6wOqafDrGQMZMIh/jlM/8tULTP1FGHgBD87Ptss1PDV2hzhnO/Z
QOXn7feQkr475qHQgpZPznKEvwQQbhAQ0V9wV5Qn2lXw6VwDMzhpqsUIKf19u8F/
CBGBa2+zaR0tqXGbJ+Y4WoO/um96l84FHGBlG3uMnwZJSle0TmVSiBxlkjilTc/m
8UGaAThYx/vryz5vr+OYzwp/jrG+/tKY5rgMV2oFGVEGPm/tf/78zo8B9c0VtYk+
6gTqJ6PvCaaRnSlx/fL7nt/r9aejK1wGYp/paA1CT16t16AcB0TZ6ohqVt41JaqN
Pu/L8tUUgqaYlmm8l3bRwKz83QpX30so7pkNT1dYF7pQ+JwstR++g/AjxD2NpMDT
ymt8/tHn9DiCrr9CirUwFaeIP5LsKcMtK12iNKtMa8QvnRhZezWP1sLH+/dtWT9v
s2qJl9gODBbxXEDy+vMoMAvlmHkRDJSyexTntZlecXEXJ3nOB+dK6ASRN3ceHy67
JjyxHRxYZxdfMItQJTs8MY6MuvdPAEOg6I1CbCDIBBEG2nIOGdrWt7JpNUODO8Hq
QoOXLNglDPTRdDm/7hl1ouqsE0zd9ykqE5BDjfbOKBXmqQuzFe9QVGgtB4ZatatO
STR1snXsf92yOtOkcxwygdxvzjmWH1o4CpHjs8/72VORr2F0km5aQhaK2lSsRJrX
xtFv0igwWbQw9zHwGY+O49Z2AQYTBzGQDyeVQw5X9R97NFAULd916nyHNe7XwkoP
V2zFGM3kbe2Pre3dnJi0pJOHRrnEHZd2ZB9lznaXvvfF2F1u3n17vItTiTaDvgOW
+ScIZq3hc87qa6B6PJiE/EO9Nvmn+SvwKvuUOqRvq2sjTGPB6QgFo03MHjYMs4Yt
Y3huTSTheXSIamFSsk3+ntfILZhL91JdE4zmFAGdC2pcWLZkKgGP7jC7afMjzlUZ
id/BeqcD/16sEsfwlaLVD1KRXVM3PyeCh3MPetA4dDDVHa1usLeppKrjMHNTB2yn
WhYrDdl3IPTBm3heMl7dteE4KpFsBPHfTRlzMCvXCqSwkLA76Rb5FZldiX8gXEpN
Y5kS6wxEDcRI5ObWHKoufmh2dOj+6qyvJ6DfWoSWcxcGNKJCyWNv+Xe732HUPx/m
WnWeSQAeHbpYOpzNoupZzTWhS99ceHLl92ukHDQ+F28N1FxT+mmOQKR8dLgVpKs7
8h0t7MeFRpjTYtxsba9EjcpFEkGraNuLknsl38dFFvPss+pkWM9cs66Ss/1DTHNa
F1cZW5GL/btuqRL4EKaYnQIAQfNrn0kkmYxTUamqfctHyjPb3LYDBojCK2z6wjJc
FAO2kT7ffebyebXEQVdkXKd+1hezb9Hi2gpKf3p8WGncRs+iZ1Q1gzNo3D0RFj+/
HAIGe7NURzu979On0HOmp0m48myvKQ3BQIj9uNqa37B3Ijd8CJS0VZVXV2HYap/c
CdzFNtkhuGypgUClP2zMZqJwTpgzh5JD+LdeR47HdI9eg0eKgzrweFNm1XNy6AK7
2kMJZvn/RlPj7o4F8WYMIZXkSrsLkCjQDDo+2dca8jeACJyQNnMjg34zxQtLhrCd
E4C+MbqtlXNyI3bR4PxnrXWLJrohDlihqUdMToO7KFqDeAWUWEQPz5SlmCdnWngj
Q/amJL3e4ucu0G6YMJHjIedSxy4vm9nK7R1zrYSUBxZ/B1gmf/Os9QfwG+gM1Nsi
Aczn5OGvblIekviRYr+99OH+axr7UvCMn6SQcItpomxkuKyLyeWwNUJB0JViMPJ9
dvUNlKr6s2YaMdnEJji5BmvL6Z6DUeu5Dy0wLPqtXEyIrEX0ei1BJ9TDwZ5qVd9S
50EVfKDpVBu7g37GOpx3ndDgvEVfrzMN+NrfXVZue5L7HuZuY+qPvMcwhVdcCW5V
sVWAdDLitZzA8NVNeY1zXuCrMBxzOw69VawFTRo2cpToezIQKO2k1QM1+7mLmNv1
aXhESOrb0X44d1ZwLhfqzKGXQBskQ4+7raT+nbbLTkBELATDpgaFnfrdkEAB83zY
cWUCD7dqMaZj8PKZzSfJpwO7IffVX1GSoczcbFXaHFUYXZUUqXM+OtduwqIx1zVp
Xbjp5WXwh59npg9SnIF/zdHp+WRFiMhlLkxXliIkiASr1QHPwzicD83hEOk9MMpi
tg662fi6ygcse1/XW3ewO5OxvA8wDIM0OPh3mhC87sXMxub5rwCD46Bh1lhNEJtX
X0NF1lqqfx4TvAQzHXr/o5syUzk9HSdbWPW05mL8a6Wf8xqaNlZgP2GYrD4R8bDM
dvaABHReGXNpQ8n+2AoxtbQhrPms6qR1M9QKC9WJhF1aqU6+2wFUdIgfhyAx8Bhr
+UsU9mKYakkUxG8vxGprFW21BsZ48rBnDr7DzaomQdmU/yx7Gm5y1/jLGvDFsxf2
L0uETWa433KnaQsmKjwb5PpMa+MCTb5TU24thUwBp/2d3rojrL0KyaQmVgJXnoNF
gOx9UY0WDlxaw5JIgpXwpNiiOqp/UAFZ2LljvmTeivVcmcJAmk9uuOEbRZT+f42N
ioLKsGCHfzGsHYhb5wNDdu156H+/M1Ub+Jezyzy3vdfLR0sbTATApQrlxUAluhRc
jTLn0H/neBOysRlsKHd2gACFTcj3KgUONNXukjz89TDycfe0zF38PO2U+0VX3Yh8
zeeUKgSzfR1QqkRSkaxAvMnRMyWK/C7M35nqjfEooz7IWOduI3J1NJXANSPHJMYG
V+tvDDMEDWcigDnFfLal3zsUkV3pI1dboAUbU4OiiwcSI9djoqq6+hnO+jk31vsb
SNQaoRsBwCOHso4wX1GIliKg3hfhoN67fhqwRCnCemGNC6f45oCo1RUTpWEG35Xc
roPAyYRkHrONx0zhhBfX9BPlW0XGeBi9/Di+dqXIIR7C5i25AxA64gpOjjk46iIV
4wrBa1uaLx+vMHc13i3GFyCjkjZtB6a7XzXj9dM3W8/GhXthnOgTmVhSMOyu5PXq
XvYrgUIUU3n0Qp4ctGlN8qoVVSw1S23/D1mHgICN2SucqWzLl/vE18LrHI8CRh6O
YJaKP7ATn1kLwknJ1WRRLjRP9ude/sBxKplC5MpbEuHSOE3+VN0ZFQ/JPlGseqwD
aiEdCuhm2eIiDokjpTlJdPPUsNdgHnBWCP263ERa9Lv503LQtRXA4bRdUAIsOO4Y
AroFVTKcjehPIm+RPHYrsVbVmM+kNpRjjz/oG4vnpHFWErEV1QbcuJEJl7NnX9hD
nS2g3JuWt4BYESWfNCl5jrXtKV3Te77pAso18N1QBODjQc9lWJ22tTDZsam7bk52
ynw8mdY8wkjqw+9UgHvY1x9qnh/7peu6radHSSwYLH3ps03Gnc5JcuPwbSCv8LNu
BfJugBq0/Qryv5mqAag246KTFjnz+HvjnGRhgWKaPU6hVPCiGVk5jkYJcLujpUFt
ug8BwphZA1o8lqLRB7EeCGAPWmF+sLqG8nMOJ1bVnA3uAB9/6eqKtg4rz5dAGl6s
FN/37IG2hcp5WaHiRM0WhNfDgwc4HM3tKBoJjfNw5VrSqHSle3LZL4PCFXEd6SHk
lV6Vrb7iE8nUBniZ4XA3gwnz0v9R2TIf0mjNG4Y5UJkq+Q69Bq3BjyHlc3CztKkB
2uaKlD9VxMQdD43255OPWLAVuJN/cQgHJxXSreDgRVWvoF81mYQ5fl4cCk7iQVPq
O/LRKWklZAKQInwL53SQBBbRhPA76i9MEg/uwiISUAYkeIdPpIzlHfOLQEWsbEoQ
Yr2bM8jfG7Mr2uawDLsgleLEDK4Z4LIvQ5l+pR2WVTjwBfpp/f4urcTBEbGiOqZI
3DeITPo+q3WJ5LVxajPPJXIJdPboWaZ1Py29cae5pjbYrEUq85WPyKkNrXxXanIt
d9DfW8hw+acWA0N0g9zORmim9W8Pfm2O6SVA1CC4YI55pTc09yzuckEk+Ik/0GD6
ZGCz1i3JSPOjW+pakO2ek9nfCqnseSRHhPVxiNUs6BEIWeqIVARbCdoGL5T3QZ6v
m7RJYeGJa4jT9Mxxy/wpaeLFrEogNa9MCcEwirmQtpDrkmBa8kD51PxdxdNgddlk
SSwOdzo9vXyaexDQ9wI/EiXCfkV6eFizCVYfXIQZfZP9E8jLsui51sAnL17jKcjS
lL9dEKSfskeXKkKSwMdDeQE8Ou8fLm6z7ipL7GVfprfw70emYnL4Fm5LNbYQOrCr
7Wq6/Gtnav6B8MegsjTuSzcAbPlFBQp6IcK8FeFCnbqdsj0OyHIARp91xYJcIDD0
ScjoSwcb/ZybvyHvf3ziV7Oij6cGPS3E/q/BMi6xdP0flWSl9chb2xMQPF6pSLZj
jVQt6L2+PxPd/csiyA88Q5ouNmfn1NqSCX13EuzL9byERH4ODZNmzdTQ8Jx8qNf0
JOzPosSC/XKNNvsilt6/mBkLMML49jEXqfl+aOIVLDJwNm/7dGIZN48vK+NPreA6
43pgiSTV75EFlXtTV9pHr50hUPXakCRd/FBpUP6s3v2Hg24Ths56ZlY0zEoWxs/1
dXcRcQWl9Gmz/kOEBb+ZZqln9aPQOFSGPVU6UI+VeamhE+N/X1rMOOBq9cGJYP+C
DwguPajTH0pkIEaoPYFMo6IJjevL0INfpy4h3Yw1918PN1EVCwA5b2b0MJuWngJB
aL8Mn2O9qlcWbYgko6UHGMoLTUc8xnrmy7t6ywhp1we3pTbTUyA4NK6tAnibV8cA
nxdC/QKd7Bnld/oS9bxjfSnCCRbO9aPR29y/yYvwcQzCxzHEN39Wa/Ix8iiej136
FaVhSUGUjtVtHYUcsWWkak4DD+VQ4JwLHi9qoFKEcxMUxDm7ZWx3R5BLHmUUNI+8
DOLbVIRewby+KmfL7Ew+1v0k5XUywSTHISSQOJjXc6QKSi9dJziWTC9vr+I6L5QD
XFAoLVTs1VinB6DR7ctpW215XUbqXYJvcEvzoAxbX8yFAEAtZgQZCdtmWJ5BLA0F
1tAEu3D2xn/ayWx3O5F/bOEfRQnKLsSYOkNXEhxUEm5OfKZTwagXIahBixTbn2sB
QZha4yXTlB8cnaJJBJgenN+2w7uga3TpAXho8PzpxZl+Pk8fD1rAHK0poIu05SCX
WnHZbI+hX0zIZjhem6rgKa4XLfcsTb+H0UMlenK60m5Nd1YiPJ6MElA6co1xXOz0
I9ktpbIBdeQI77tH7uvUmYGtQmIF8psCnFKpVdFzMciYMB1ldYQuwve3EXIfRDok
61LacjiL4cO+kZ7eGYUe6bEzFJ2rovdseGOIBI2lRpnXDoutz0MUrTbY4On0qkpz
OWPHviXdftundjUpdpytqpEOHz9TPIC1E4n6WEzxINztLoMViKnJiZZQMJUDazUq
exkc58iiDhuAiB/zeQM0H5wKAV+hPDlBeEDWT3ATI/dB18DsY/bpTn29qG6pbJs3
XyeRO945dZZlyaE8mq7H91dU8vamyKpVMYRa0nOwqLNBAwYZYy5SHF4zVloDBkf+
HMLnIckQtgPU8mjTw307Y/RiaJ49Hj62GuPlW+YTZ/YqljcGZT+qgDJEj1FhAhuG
agh4WZdP9xEMKeoPVl/eMJNsOxyNMI1mue3sSjWU5n4uR2lTd5iixknrHKLSF4dG
k/hVqK9xttYZnW9760Jt4RNfvD++xToHsM8001gyDswVgwq8QzL30ywo7TiedBei
CBW9IpcHvKPLscHVTazCVG6vC1gJjZzUKqODq/fjQUilsfsvXHiGQC3BHsGsj9xF
/JsWAIbUD9sp5RYYWnyhFIA2fakUdgnbOwYH17l2/J6AvWcqPM+vahlF7mO+ZNlv
BulWTBifodW48c0snCyICSvd5w6TZrjiR1JeAa1S2wSE7RJ1M21cE8XeyrjuCEC7
Rwi+AkZrupokkNubdiyk2GBGtRGe71AgaaTDEhepBZ/hvjH3oibJjp5BzPrnUn77
8zqhxsDNOMf7Z3pfXrPW021pImKjiJL0pAvGOLATOx0/ato9Xyv5q/EqpC/MXd5g
x1Y5L5fRa9dZrQAvWoH9UA/Drv+qNjEMmmjeUCrrvHNtAbw+zqtZMWUlg1e01qKP
BD0Rl9YUPHIV1Ah0nBB4f/6aDQD0FRlXdvrrv2E8CejE6wp3MEmj88fc5r1pZIXr
lwDFSO+A+07KeP01NFE0RsQpaqYVAZHkR2qRrHrOJG8iNeVshcVgQUz5x20Dgbal
PAmuq9SFJBAiJQQDym4Dh+varrFScYgJX40mlZs4IG+es3C1serFmsSu+1c+/f6o
V0hyhbIna7nkzt/Q/beFmPWEKyJR5cvB5b0qnHUB5mvo4shzYksqK1jKUBue5l9q
+FSJ3IpsnoJo3yXROOABDprdROK+ysb+M0VPhEHIobd22wlqCsxuPxBjygn6P8qe
T5TQnERJUAqWhtHOK8MY2Gzm4dQSKSeeL1c3InAX+XJIuKSOscnXTGOKItOzaHVL
UfZfFJgt5nOpdYFtOaYeGcCHSB2fXdf1KrPraZyYiNw79/6poNXTeYNfB4b5Nsad
pJiZVdi+DDtTHw/qNUnRr6VIodPAuN5tJmmK8fFgphVSCSLUrDW5PtU5B67dlfEZ
esT982oJtK0DFIe2UieYGCBGOL8vFoYRPFSzv290Vc3s2gxxiZk3iIRCI/RfhZpK
PKm1LHssf1cRzIJMUD0k/TS0kHx2N+Nk3ctXWUqCiqVpnACGskAo1+2UkP0OS4Fc
iJgnK14ZmUf1lFP/uE+OrriXnfL9TZqHOBC4CTseiJ/8QoTeOK9zckvfWcWcUKbw
tvI+8U8zM4uOnuPTeZC8swmS3TEu/Lee/V5e9IN3xg/CdhJ5fLZsLJEgjYyDCead
CRbpQs1lp1dN6sV6vOII9+I93bGUYQKMk2yLexer1W/PUm3z/U8MFeyRpGAtVOo7
+s/iA1+lPcjBQXt86DBCUJH/tmCvOIUFrlnE0vcarlpBk25IymX7qUsAP39NrGvX
vAcCZI2ZLaC7jNt1Gni7QN9ROL5nWZd16QoQqEqXuIkY6DX5kySeYlk4fPkD5VL3
GHsJmu4pVe3KRDnpXqA5CH1LBC83kBFSAKx7AYT8M4VoH/TuYaY+OHTEc0LrNVuN
s9ZcK0ace1a2eiWbE+FL9NSLSLJZUGgapEmSk19tq+IIV1dgAahGGfY71V12ugZX
mC/A1lAC5ZMON7tMFqjf5X+OF9y1qQgtXYmIBZqWUMcBicqvA1yGLxq9WDiOaeeT
EzmkVhekFTpVYC79ozWtdrwfoA5hIiPXWZVOl9w8DYmltf6qj/lZd+8P8zz0BDQK
SNIDlWLSe44H+yEtS4aOqjJeN2+CBIvYw45jrYn8DqMn6Y492UZ56l/Y/fVh4Nhp
/sBb/24xvOTUjQs5F8+rZFOrmIBUmKfnXo9Fzev+vBa5BNoebot4sMzQlFRaoKRM
tlmQ/pC+g59USpSvrlT+1oM+c2NSaPLcYHY78MqEmbKJdpUEVUoNFGIncKwEyerH
ChT9HNUKMxjorJ/MygVQxAjzpKtoNOLEvRXykLeT54xWR0gTymdrRJfFfIhNhTFH
H5qG1ZcDveVw4F9M5ifl5/5BKcBFAtUn9nw+pyEPBt4D2hSeZaVrSEd7o2KGwjFn
7u/rgapVzsck5/b+5tVO+uuVRZej87iVM8kHxUBEN8FFUang/dj3x9NIbY6/Vl2H
8HB3OkSoybTGqXPls8Tk3DOOlFukPEfShcDYQTx9AaOZsBkNr+iZ87LdvxMNBgMd
6sHkVQl1XGX7uaqEG/lSbH9+RHcGPD/C3YMmVVGIOY/eYjozwOBsFkq/lcp+gw8Y
DrxUubwvYKvMXFzRtmevtVy3+b7fwwvQdF6JmnqMGIbrfKer5KFQArpTlUe/8hCR
5+cmsJuTJyxRy0c1R/kAgzRFwft+qaR1fjpZyUrAYun0JQOLA5SudQbfVDJU8DAI
BELqApAfJDb89Z1uLVFthdWaHpCBrB08MhweSUssU6tAn5ZAhLLgRq7rWllE3OGD
I8Bji1vr6G1l4KtF4fQk4Dy9wHdZ030nPZP3ODWRl20mGWaUn65P2P+Mps7vjWUC
ml20NTDPo2XvCSCNRQ0a75Y6xZaqXBZwQW9PcdvkAYRCNyiKr0Q5p4C1F1Iqf4bT
QfLJocw4UW6sxZZDNOBj+fj4PHr7uMhTRn4xLug75/PXeYMcMhYpM0kPLifSsOuH
wCFv6UdIzAxowCtWncrcIPtffjbFjXgtPB5LgxNjyj30/zCrn0rTcMFBnhJNI18n
R+Sw8ohOwzMfcPsdo5Y5Vz2V430roDsaP/7KaBhD8ZjvfR7f9lZxbn4BJ6Qgk7t+
yr0lUIplISXKWTlbuOhPj3+6ED0NaVnxeuBZoq/z1V1EOagT9HUj9zsN0xzqemVy
nLccCdLLXZ3S1Wlg1RXn2D21fDPwpgTYI7ccgFhjCFcgfYnrPqdS9kR3XcTwcgPO
CGgpfEmSHUaHC2LLGl4+x2Y5Y+0gqBcQclVzVR0OuSF+6YpYuzhYYN/hQaKlT4AU
iSD34LZAQSBix73ZLEOelgvrUM93ZQP7kfoktvmmaPS5akR0WlKLa2uUxM2qxxZI
vFIhfwu225Ewy22Z/W8uizsRfN2DrYt909lZxH7mpXb10uIXEk334GbI6rwkN0Vu
JUHv1YP7HZ7KcbqwNH8s6lO8Q/p8nRGCkDJ8AIeszEsUoalNaTM5A414OCi72AMS
SjIfVIyzsCPUZ+CupTBxDrSBtq6FeN8y57UXhzSZ9Y3ZQX7W7HvcVBgEu6q+/hZJ
A81CHOGUn7d4Qx/el2MDSz4/jjRM1ysUa6ipZbpzNGNMIPt80nPNY8Gb+wbmDXug
nEK3yjt60xzHq4KI5kGYn9YByyCZ0bj9c0Sprt0r469WwQxlyJ+6QLLGJuiocCal
J1qbCgBjHPp72XXSbAr5NlOZrXOfqd36AG/1wGyoiG/JZtVb6YKarCot5gm+rb1M
gCT/5+D/F5HgpEuaxVFdNP/E/O3f7o/7p67+38t31dWp45reO/o+ZmLRsgYhFZGF
8YDd5+t7+dNtAFxNOIPr/8Dt6AMFdWQ6c413HHGH6OknevW8wenCJPQ1oroFNOo9
R3zoYeiZ9VFa1SpIdX5w5QlgnRnHUEHyTzcRnB861zaElcWilIbJvQTJXQCm17T3
J9NTvnWhTgYNk5BxhrhtFG2a90hBYOu8pxCdS3AhyEq6caqyKe9OzJsiuhIFPg4u
lHyz+YxHgOOys4fpyIqlP45uuoVG6ti5zyjlnQTgFc0u4A+EgOxYlA6bzX4klRc8
JdAdbOtwt/jYmwyANEKzs7ItlKbfAQLJ6nc/YozJ/FzJLO/0+PwzAicoVe6vr8+g
pq+tt+/E8yMhY2LkaI3gEBWkhwwwaNaG1H5k5n6W6jHWWeQslC9l3iQsguKy8l6A
giO9j9DjFD/7cdm9oYhoaZ/BEqXC98IRtaAES6CSde3/I9w0vCRQ5y2vxy6VO/YY
DQXeGmzkZhe9NlBes73ZWlgxf8jaEjDDEuJzcjrqyO4C6fcDBjm0xqSmSlr0zox8
FmF1w36tefZedOmY+IeZnnaaCygL0gAuOImD3JX0BCBucaLAhemHLByd8Nh6UX6i
6eLfOFEmQCP8i6tEARUPvXCBWwLs+1E5lHuImIFqYHIP8XxqpRK5kZZAV2NpXryL
A3TqiGFMMcnKgm4X2sc9ELZH7a94263SXtircYqNdJu66XP3LgHYFEYywdr3n1jn
CAO34FzQvWL04RNVa+CQlL0Qmr7U0vIRdW3kGjo8lhTy8Rw3tS3vq9/3x2CJnbHM
Gp9Jpsi8NXqz7HXSivK6DxkYUdsTLFjw+LBNj6erTKTpXlNW587LoWsdg+iuzaPz
DrcenoF9M+84BidCVgIhZlxm2R5f9E8JnwHcYAiBHP1caV/Kg2G5djNtdC0zEjLk
Rk4k8zlEBhfXkgcorGTS1Qu+FoI2JYAleaQ3SjB67cEzH5otK/zfbaEhaF+XnyCL
BxBBMay+sCStWU8FjUyPIt9JVaGOqVq8bOxy2JDiS8ZR1G1POajaTs0sHUvjm6fP
ayDkaYTUij3Yk9hbNPvCPMBl2PAkQHvB4Xe9JjY48jxcpC6XxzrhnYhZoSD2ZI8o
4S5TR5wEGc5fHsPb46kOt5d6pxKfxUpkplIW3/E7v+E76IZmvVoARIQsrrgQ/6h5
uZxphNYXkPz6LI63petD2uklnjgM11AYJ/FqDBu0GVOJISWr1eS6y48wpJgCLxmH
1sISlEzhqcxbQa4swrYo4J1YBYG0f+ppTCs8WC3VFJYaPRO2E972tKYdSUW+6bag
5OtwSzYT2CUINQD2HPzmn+LDo/GZeX8xUQ1WRShl5ICkFGr+WeNfJYvGAgQ+EklT
iA+C90LXXw8emqViQbr/9aswc+goOXTfD/BhiZe3WHAR363IYClkNjObtiSgqSrU
wDbAS//o0vuUy6giffpWQ075YTTxC750eev5h+o9ShfwJ0bpLLOfIUKv1RKrpuQo
oalTyel/1N6v+yG5ndVYa7rSklqFT5l89dZ9eh4Q1gpbdQeLJzJ/OW2OEJp4w9Or
CjgUkox4a/Cmb2fugcoKQeH5FuWyXOZzdUIIu4q4oizgu7qEEhQ3ukNjgIS20zqU
itBluOHSslf2OU1SjKB494AJFM1oI9R2YSS2/0x79mUys0yefju4ZK4k2m3q/dL/
Fp6/fR2j9hiGggzWfTd/O5XhO6ah8a4z0nx6H6nehLgMJkbDWdE8NkZ1kPwrpWuJ
ZVUg6EYOo+EjHnHcNTCDWgbbJLoQqq3+fMkGAHeqgRCkeaA3OwTxuVmRvbluwg/t
JwF+EhlbyAxjKx/mKGBNyre//34XH7d8W613kuTBdjEtZZEJftbC6j6goWZp2qZa
SOhy62ek/VDNlB9lYwoo0A/ZnHUvFqXmKh2AIfm6slxIHdNcJjZyzV6zDTSkcbxA
HtuXhIIsZm9AJwhCLXd8asmrQelwsEGEDyY1tXXU9jskZ8cCz528DmgivpxVstow
nSNBVXlHF8HxuZIV2wrDr/VljaNGX/Tiy3Kk21LesqqbQ+dHDgG6S7+mNhRjNrpe
kmdCXsD+P6L46Xo55hnfztmpOsBrpYkeN1K6PoC+fC1EuA+kKc3nf2DYmWBfhPdl
XXWjUjFw2IFwg/1GrmPZWoBt0ZZjLa2tGp/JIgGpqHzwGR4UomZcFcRp/X6SYb5e
zB3bRrjG/K692EvlBPNlUtPmTMZ02AFECr5lML+tbdW/xuXu0z6Cfc8SWAykQJNM
yXOx1egGTauDj8ycSpO8aL/n4K7Qt0tNu4NiESuRzBS6BThvFYxEPyRb9AONfmap
cdZSOkaSGITClzrVwrs+BGho/ReEZiyGpTuB9qlQta1VPeSPRqA/UrQySTHmIgGQ
GwWhkiuvu2mzdhCahcsSJFxaeijEfP08cAutyY0Rb9J5lTik3hQ73DOvU940UOdV
qu8KoRHr7JsvAEAmvbhxN6ojl/a7FS2te9xU0zfy9QA3gfRe756tnjfT2TuNzAC8
wuQczfdniMQz25+x+Gr4zHnLGXDJ4u8hiO0lVwXRJsF7jXNmxiq3B+QgzbeB0ZM8
i4ks+lupt+LcaRvnHLbmGJHc8LzV7hny1pE183UWyaNn3PVEksPsnMFY0FnivHgI
RFGFE02AGgBskQidJe0fbWvNnhRANYqIsdN9BRDHEBZiOjW2Ug5dCLG3ttsk43y0
J7LNB0GDOJZzKZcfh8wnuaZZEsVda+r3qirGcO6CvCD0MkB/2IPryxro5bMiiLvb
8p4Q1/VPRMz2Q7tohm0dWIh38Qlzka27aSNriGfnHTpHOvaX9o6NUnqnlVBbScXz
kZ1LMxkJo+kEDB8Icq2ltDS7RjQYXKTcHdHEL3FvXsA9ocNNQh/InMffaCEPaiFQ
N+mvYeHZErmEojZ14r+G0ujgLEYuN7I0OK67X+5PV4hq5bWk7z6s9g1ABByDZxbN
48Nd5sDK2idtlHSa9sobVEm0UZU4XKpa6T/7ubGfTEhRukknsoAgILzgHFPZKPS7
w6XK1eIeFSi47CUcglUJ+zjKfg7aM71Qt1CQQ/EuZlRMGL+9J5Z4sTnawLp2lPpz
l3EjthQjQhNY0kwElDMpj/D0YzPYLJK7j0+LNX85KZ9d9gowY9d1+HaPWOe3F3Yq
CyEB4zCgV/atJQGCqoYhrLmbYwRKbJW3+we3az3b9ftPoERl5EWVlKwJUwF0OKTZ
kF7w0dmeO3fMKdK3JyohAYN2N3MSdiMXfeRMEyMQ/DQle6YeHq4jAbWOrj31DdVG
Fz2y5nBuXs+nQ+tF2GaG8pzdw0XmbayjHU3AevfFU0CJIt/TYS45tYE2lELOVR7z
xaQ8+xPkU7y4BJiHHSmbmAdKzvDRwMP+kNjnX+++l5I/wT3Ue0ZJSRen0Lijw+a+
HETSvDowwdINRhdFTEljpnWCzoQ3WFzqBcwo1oG4w0hN+w6hk1rYG6150AnpFOXA
xmy00ZiRphmg/cWxwqerKgaGX1EnXYogVJ9QR7xqUkDhhQlPdlFulDHt/H/X+2vF
/HWVnOP2o6F9pK7cfAubMrUA/jQmWPV39S69LAEkHDvtdEsRD3FG7YOYmvKCEKUg
yYnjoRlOJJs8jH6j9YH4ZUF4M1XCjdQq8jKGVT1lrTLIPxieT/y6+jxMHIIN561V
b5w/0tSthV5kcSps0ETLZw8GzIxgq8hYTXg7u2jd3R45Fq2BNvAJIpEMIn23C5V+
Cy3ZADCN3drYtGmM+bW7UfTL57hUeScDNul+ltguXpAn+R/Y/aIskg3Qa0gno802
Ay176AGP1CA4qA4vmkIACuyGkhU1KgcBbT6ckDmHFNJRnVDKKbUs6gZ0ZrCShxCc
IETw9HZgNL/tO/AJ9gxbuUrWP67x12l/+176s2ouJ83bwCnmN57YUhAaKIWV42PT
h0VrqU8ZYeTCd6Yqu67vDQOa/pmkrTmJx2V0oDqQy3/UZC6cQger7zYHn79tjW0A
Qk6OxJxkg46qPiQziYUd6UKmRF+etGIWN1yyacI+1TV850T0X2zNx76CQQts7fAp
/on9chxIvMZn1W12T1czCTjVk7h7vc4OM9zL/9AHOtgnj9e8JbhIYl0fxOuc2QSr
YbCSAuC9r9Phl3eSacVjCbVAqQPmqRtnVH/QrERuXWgKx78G5p1pqUWlE4I6JOK0
UPWWLT0V2Qf1rLlmTkalEosMRss9VAN+adscacbkoyIg5lV1ikJJ3SZsHDP7lUuJ
4jUHyTXuHMvsLp/7aUR1VayRXdRoVSDrKNMqmVp7UBIhZNQG5zKOsO+sA6hEgZgb
Cw7brkeT4m85mIdv3y/h6s18MtiIri81MISKiLMaRCXIJxAnnmqMf9Yg/uI+jGP/
7I/TWpeIJlW7TJekMfaw9/wY/Y7tJgnhNqkIrJtnrpQddWf+13hrXIpLuBLplzYv
/QV6TtSL8eZDXi8awc/d6F4HI6OJnThbl0iJCHH11Vmw8EOJmQMIfwq4OQ20mkqp
lg2wfSYmDODVUPNa1toemj4MbQBIP3FRwwYcJwENz64+8cD6oZDfb3nCr1VtDMum
aKMZAt7jjadZHQipuRS4PN0UpA60CYGzCG/q8Xr1weEpji4T2xnG6xqz4BDgvbIO
gyjt/vKLKK5HYE7bceyCpE6FU62YR5UhrlBmF36l0c+ULLU6xquj686Jw6/ygaak
AtyV7guBnNasg5QiUQVyx2aYf7PYQLDhCFPr+ywAe/NqZbnTsQrijWWSXbwXggz+
NQ/EdzjS+nvRvmWbpD40RdGNfCgBxvsdNNrHwOLhOdf6OkGKIbq2JnzdJaDFUtMN
AoKrduXFH5yBLHOPkdJ0Xk04RzoIlmYiqvq/2SNcszM2lxi0D+7J7Kw8ptl+6q6i
`protect END_PROTECTED
