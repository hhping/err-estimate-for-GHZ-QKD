`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DE+KBnl/1FmF3vESPYz1A9vzQojP0mrEUdURLQeXWMzilZISkW/m3Eik97lh7yfw
2eQ/WyFoqcf/W5EmUE6E47BNgSqjfvxgeGDcsGd3Q7BCG4kpx4lxPvuKd53dHH7I
gNtYxc5R12DbZQQr/73ixn1TojIWohWkPmLCb16p7eQohaerUVSTWW79TYMMFrOM
iRfeNAVf5MOUW6GHLZ8cz3JZrO72vZDPhKVMErBF6cX2JaN3606uL4m6JvtY62fs
RG19dZyYu4XHDJGWaBXT1LDNtoKfYXnB+3gBAcpbqzDSvgUjuzNt4d/Hi8Hh+wUF
9I65LiOcS0Qu+SFvCE0qeAr0LYBofoY+dkU9AU192mGfZP3RzRAYCrhmndA8ZJ0n
+gJ9Hk3+Isez5rrCRDAx3w5imoDY2WzjMAZATtfn2cKSPMjw6CL5HT7mLv2Y2RIz
XrT1E26v7sQNDDOZGnEANTU6dzUbe8SgTWHTHwCk+tzzEgyhYdQO0U9CPMK7Scah
blYWl4s4lzri4WkPvy/XL37zd1UqnkXLp7JWUDksa04=
`protect END_PROTECTED
