`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eG/gpdB2+H1LJDns39IIEpQme7oVen6H6k/gm+/i1y4n0rMVnDOzI4gJiQkTUXzi
h8jk5AwG6tFBTmtVNV4PauHhem2EN6f9dmsui8pt7k/SwlxORrlvTf282tFh5PQV
bacIfHAbbt13O5wGBe95gfb5oFC2ZKcG2KuxjNkYq/ca4XqhClD+nHvSHObBLWga
FWgDoqPKyN6XIYQJXRaOOktBEs09sNgALlqgXWNu39TR07GT+3ciA0uvqYjrX2pE
7KprFKsXXkgHr7t8kC7zCGhzVyv34LmwuAAKFyNc7qMAu9J1Jxiq+jhH5k/rp4/z
E+LALwA+gYCov9EbZFsLsEH2OKwuTgJ+MONKOO4oewi3T7Bifzj88iKzB0uAZTUH
iuT1L5NvC/TLBh7iOORc62EbR0gF4LWrycDpiHICJAPD9d3InfbRy77KnPTZVcxK
TY4RAiXbMeUFe+Mik6JaaXsLkENI0Q89OyYKVQqRtRPedAHZ3Czvj0fcOUK9sOE6
l37gf7z4jYkbNgzfV5wBYuUzR6ngBqMxLzIjsoaP9hHGhPdiBeKQKT44SX3B/ahX
1eAhHeCF1YIxYq64GNoPLEPHSWGhmJtkCZ1znCTkNdy8AHvFfh38jDS2fnXXr/n+
IF/rUQNzUk3JN7ACcBeQei/a1TjRotk5EtqCQxhNAzSrfNCQlOyBaM+cu9f6Q4k2
Xkj4VqDZroRPqYT+2w1XmePgAXbD5U30U74+UeuC1aZAPGtQe2UZ15nwBuFcZKN9
k2rst68wr89h7OEzdwRIQM8jBR3qztrOzYYXJf4qxXIRyRKsb1p/B76EYLGkkg6M
sMyK3v8EvEOe5Z6hbzTMBqTUsxScApFGbsK0E3CL/szYTjkJJMB4L0JThmeWLro+
I4uvEhDehLKKXKix0EGHj2/XF5mO3aylmh/B0gjrqS/yX3c8jdoJ/xNYCHQX2YoE
HTWX7h/1I1T8mIWk4xu8fDUIy4CN0S6lBpjogZqp9NVH19EqKHgTcenfMqGId2Op
NPb+c6EPlqSntuZG4504leb6dJmcn9L+O/5QRfkgpXOsBapokIG09xi01E1tZyaY
gsUTSXNhtxdLEVrK3D1fNi4SI88jbS/PbZBJPzLJnBvhM44jfavJ0OzQ1Srixm85
Xii0nFCE7Ru3v69hfLjbzQbG6ZdmQp/Ll7WCgHLA3mzfWTFMHHBkaVnrmyiXj6dB
cmjE3zxM5+jeOz7IGz8nQo1NeB4vRRlciCuSC0v0ZMJeV3IHmQh4s8PPWow7duL3
laIZ7ViWOpHUlM3fB58rXzmpYiWw8bSzyeWJmH3XgEmmtrcjCUZ6XUwHdhulwMbX
C1GefxylGMIE814xEWjlpxtjnatbur72QppLxYPgDORAflQcEehhV+T8yfFmzUH1
Bw0lcssHRgdD6j8cUFQle3DyTgzAyTN5oHicS3ygZ+ysK3JsEIJZQS2YX9Y2HIul
fVhe1UkKfd+S6cEuT7et/LYU2OD8I/6MY7lbUo5D737LuSWnscMadOdze63/bv5M
IBR4n+pBo/pphSd7a8OgsgZ5sTWP44HTKdM9eLy5KrOHNCdv0dcDOAZ+3lgvR6A+
hWPSaVyuddXTCbFRhFDgpxCbSkQ2TynYEKyO7czrHJe9RNuSIxMMuBh7sb+OlvqW
S/37jThgB+W0yDXmHPFXQjWAw38y1WKOrghtqguF1Yegb+GfpR6ixk/DER57RBRh
622Zf8MzNXpkzj6CK4McNGkhU0uEYCMUOzZsWiDqlFQl4LQ0gIVOKYaVub77etnn
ws+LSmKNwXVz6ksrkYZdZCmlXv4xHDQ5l2Lbl6mQs177JTPjiSDvybernUP6N1h8
xS1wjxgQrcWtTtn4LsXb8geIFQOf6uANXpGuejoteAhX+ok1Rg0IxmBnR8iV+uab
9oIrBWd1ycarYqjoRqtJQN0WKRxZL4ZZrnSTyJ+ZzgyJvZS0F/dqUSQ8WR4LhEey
Yx8UeYEIAIXY62yuCcpEdI3Th5puoVS65pBSWi0jj0q3oXxEYshLrNraLzg2ScTH
fdy1xsiRo2v4yIde7B6I1sIuPVFGPH5+RIxqw6PdigKkvaEDQcblZsd2g8SulmLR
k1aqT84HLeys8ntLGzORq3fgux2zkmYe4A+9l08PvIWy/StGHhOYIVbBDXg0AaH4
jcZ/IDxD6j2CQOnbQP1duDv8RWGHff/ZS7UNmBD3xKZn42e490LAiCXxI/waRiSG
Yzo6QVOx882dTmTZ2Vyg+FVZGWVLBCVVvSVwZGx1XEuUnPlP0yw9s3R8xoone7t9
czJsYISnkKA78NHDjRdLwKqDT4BccDaAzpo8s3YC4hMZOgn0mzglM0BFG9MCoPy5
1d1i+stSJYzZZKCcsPfnawvRg+X66+FR47KtNQ1jbz9wRYELgzcX1ehrSZKWHdI6
op9NxwzUcBXTE3qp+j6Tld8DaB5vbuS8m/7VoreyIv6Apn12SOzcZb8XiQAbzhhG
PwryQbcoo8RIMV+1fOnMLz3PLWw35LoJ4jmExy48grCF7ljhxmy6wVAJDvDiWLcy
tZK3aEdIcl9K2TWKBpqoh583l56C4HhW3t9Y2Ci3Zyx+NTy+/XaRJ3NDiDjKWxd9
1KuLz2fDiUr38NOPcGdKFwjWr/2tUdeOOwDeJ+77N0Ze/aw9dQ9eq9HbEK2wg/Sg
oVQqX1WyZHogmZdEZAbUzQfSRLvXTM9JNb65KJJZZjlPQMWTGG1zPqvPejxC089I
f1Mw1KY6LYD/1nXpWk5zvVT0zRE/XgkwxbM/CAY5sKbr653YIY4KbNbZNrsptjmS
bBv5P8surMloGPQRDJ1N5rGAH8qBIXSu9hmC/8PCPSYkkEVlKZnz1lQD9RPAYFJS
jQcUChgP7vPWHIBU7KWeLO/4dLRiUgaw+0j4zvfbT1QtrtL/H6K03bYW8Yi1W86L
wtya2IzyWU6erdLl5+OlVyr9fR/iUdz1Vtv8TjEBANCUJgwZ1ZgFNRKO6iYeZvnc
Q0pFNhJZ2HVzOd9hRLlXt0cO25GpfU/hHQFbO+MQwqBAJiOlniHYxVotyYYPeVm7
o3gy6ITnR1GfvxKcaFTILJgYJwJSB2MjQmik9XuvQo5Xw3AVUoBX75NparcdMRIo
i0BSLC3nroZk5Twr/gOxxDIQ3hQWD56hB5mjxo4k3gd40md7vqAScWWgtE62WPbo
9T6bCnJHsaItx3GPQ0u3vVWYo/5NHCMfwiwTzeg0pEVABqk/aNizV1N3CY2o2jFj
0JVbhr7ykpPsVTtyEgPAR990O67y/+F9K8Q5W/TlSYsoDPhNskwAW+aJxKp0NAGS
WUAdjVfuDvydCkh+nVt92fFGnybILb3erJyYeLLCMlyyN9ao+haBKjnYefrfMMJ/
459oZiH6QaBFWxN1oiRPwrwq7Vx2n5xaRkzQJH8uHZZFFaoY/ND2cCnszo2bkmdf
eH+QTUn2RwN94YA7G2G8k0J84ZlmZtvAUsDRnhgCqihNu6fnKwKq8cJxqr9uPVl7
60ppwjAsR2AVKswrHSZX36sPLVEQzLJcAYFuuxLqcTC92SEwvq5+KgGzDvecmsCl
ixJpNm6NdRWgeUhzesFWxmR6WGyXmBacGSXDfXkOB1xaMghK/mp79qP5gweCf+dJ
UlQ6UiDq5++ddd3P+2vNZtihPN+XfZFH8Nqi7EA7lEy+7HKpYj2w+4/dNYj9/Kpq
zDgEWk3Lp5O1tLdL2SYLa4nGVdvZ6vXYc1QJMmFrx9njUJMymZ/u/TA47c85jC9b
+YwIBWK8GJGZfYdrSMOiYmGEYnCk8NOdg27lcicwhqiesHWg305VbmsB26PCr6mN
UVaB9EaN96HJYpk0FAMnC3bFFsZJw6yS4FhIK5sxQY3xjhUrybgLSHoA9mxxvG+4
Vs/gPBxsKBoA+fD/jbu+5RIHS6DkC3JFQzZga0KgDxivvi9FwIfwYp5ANstYLK7X
di/e+lfLnBr1i3Q3V++n0Mh6Ero2z3oCVMJl1v8eNm4DTj3TD4vYN9k3CuOgJNuu
KSKqv7OH4HLZiz0aUq2VvhlhtA/h+XLN1uXo4opEJwd39SaycrIVGlP6W/Tk3zKW
aQjyP5DNo0lIvkhbElR8NEynWF504reTxZCNsEDqPviVyrJXIrzK7kqAcAoMah/i
Wt9bdzrAv/1+m8oi6Evau/DIqAD7wWMf8mrGhumyo6CuvfmyZqV4mN5+FDOy3ebx
VzOL0pCdftkHo0z7fpj0MD2v1hvgHSbdQ6cVJ9PH6fykNjk31rcjSBMRI6CBz7DU
MpSEZvcvzxZUrzLd/kNCVPoKSZ8+j7NfozU93pOnmpBCY6zHN34y2K0Q1z48G8bh
2Fe0lkZ/K+eHUKZjQmyN9bFYtnM+PZS4OYorpP7h3QVAjeyhvYmcYGq8NpzP7+ic
DcUQ5vBBQzpT+LWohan3r49+r1U9H6Ohs3jRaxM2YhHdVfn/vbqht9QAcfzylv2U
uz+u+FJ/biOZ+V2P96JNTJ7J8fXTCBrsto+o0+QD9u5Bkq98YHjVL+yCLWb4+E6P
EJ52uDn2DKh0RaqY0r/WCjDa2BRFzHSm520AvJNzo27uN1sV/efFimVnGFlx7Pag
jVLw4sYpYs5/vhwbD2QiuwGUSoQLXmj8/2dnfTq6HtroPfP6WCs3KehPHasllbAH
HjPg+FjwUPAi6Ruyr1RO6lza4Dt8RsXQWVGsnSzQF9LbKzw94EKPp5n6sX4afmwG
ewoSWekWrtBoMMBs2Z+3ipZqLcCBl/FTrfeuqcOjmql/wtiK4Qj0daozNCTnTBCQ
DASX5tOPh5O/evbWM89JWpiXPoT9pNgMuFSVcB8tkOj9aCgDYW0ibDeb6jrKVfs9
/TbLpfRjfhPopKr3AXlenlj5LLtQ+eS5v7XFdFM8yNjBpCstIIDy2PfQ9ADlq+aF
2KsoLurpvupV+bj0TGGAKQw4b2Wld1r9OisGD0JHwI2W5As5lzExHRH/WQahGU3w
DVJvQ267kPEAsBfqF9FzTtOoGKnv982lBF4odl9DHSZMRI1nrOv0zvjt1fx0v2wU
cTl8JbiNfTkQ1yHDS5lZMpCE2bEuWZTQduz9a1HuFf7KPpIFzsrb/0njNXZwqNRi
2KVC7pu+IvqeyAPw2cSajKOp4UxEFPBvIWhOI/wIOgVkv6h4eiPT5henAwjD/3eB
0bSoG8kjmLAxZvOU1x3H6KNCFEg6aLDaWIcmy4s9+gvdeVOgExt8jrUPaATv2JgQ
bEfZ18Qnku+gejfgmC3IE30n7nIzdH6f587YvNWjOuJ/B5VR0pjLDzOsYdoOiaJQ
tHIIEwKjKyOgUBTB9bNMQEmzXyIwytef/ISiDNLNYiA0qJ/oUBblXgICXUgJJcYk
fTnYvLkJHgGCEUniBWymOvdHLuejPskraxgIX1w1IOqcrAJhyHp6Y0QpysBOkl2I
vtkX+NA+mPmUL1f48QJJSiH74J2c6rKvhOthtfSI/StheNEQtZJJGsjyMp75pZcN
28DW99coUdBzCcZeSDXIDfePYq9GUUVxCUDXVaw931k2Z6Fvg+tv8d35UYKaXwtx
uj+ZtLmzSUPSXVP8IP6hK8N76ieYENgW44Y7R9TSZsvQikaohvr9lOyP+irw3WwZ
Hhuk2GAk0ZnyGGz4qo6HbdE4P7G8bYHq+y9NSs4mT7/z5PD0wBy2nZZEra84dRGk
6sC2Gl70qQgtu/x6stPcuGzSbARlduKvKtyhrqI/et7s16huthSnwZZlSfjr35xq
FVbP7v6mOG982Z3yuRpYPxZCv0NUbZos31e4MhvX6feepsub8YlHmn3TpJCorFjq
WxQ2E4eTdDXsRR8cgwVleIsEM1S1ymYtR3hPUzT/Qjeuk3J0uAmrLUh+3z+C4VcA
FEfVkMewz6vF4xfr3KLLy/l1/z7Za88ReNTe1WYclM5gJjR0/mwh1i0oaaJU+36b
H3bdlKifmirYmKew//5fC2yJICK4QPiXiMkt4vLq+GM7L5bW4vxO32SkDOdMVgdK
mtE8HkKBgdHbeJqJ19mgBs3otcrF4KRE/lYeCUlZVaOv1waDw+Nnbonj9jg3d7gt
Qc1nY0nbYR90tEt2zFut52k6C58bv39qKo/LFap54py5R7tANXtGiUHulRv0xBay
gjNeHeTTCQtAIdTQ6KpD0r/+qd2IWCR9Z1UCepcsyApHY5G61EXNQ6PxN6FokzBr
4dTq60d7/hAFuVttQjFO0PmUeuKcQ390khxKh0HBDn9sQN3lFHxoB551L1UcY08d
p3Si1fRSzHmtJkZ6oOsdmYE5FYq48pS3dvFWMlQ8GkB/5wGhi8tvjKxVAZbagyJP
gqpgRq2pTIMELjJMg6S7oaY5RGxpPWp+AahIWmF8v3ZHPAuljy2enG75rAqOdyeW
GGVWSweTSse2aJYer7Wpj72WbTJ9o49gyx0gSQ/n6/YfQzKc0KkoS6xUIJKumDMj
KXLRkL3sB/E8TS+Uyx3p1r9IRk60wN+CH9Utnfn4VI5oun2GiIWvMMrMcjm+oitF
PoV0cDYDE4nO+Ohn6oP3+EFnAOhJSpCpCP4o+5zwLEd0XjjO3HwufmZ028ukhwo7
mBXhysQ5F8Q+b4Rw1tnfEpV6mnObQFSXXOqh/008LhePL1B6lg3VOETEBjW64xAt
UP41wHsT2iF6nW8pwRdTSh2yD3oVBbuR50cAgzTteEw07RYJCBOSRNQRxpDcW0g5
JGfIz4VI1QvwP/k1YP0STgvrwTARt+jkZ9FSOTgu+Ff8Iv45YmKFpL0L8YLT1KpV
X4ELbT7Y56meJ4x0/unD6FgR3OxPFr8cUAINwq7SefDUHuMG2VuCu1xKlhHRY3Hc
`protect END_PROTECTED
