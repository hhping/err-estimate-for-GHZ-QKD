`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xecy+RYVZMJbVM7RpEnQZmgx8PrEn+u5/pnaKp+Z/JZ88TypZZVcX0KVQpLfUb0N
HWSjMHBD+t8dT8nCmMXCDqGCwx0+pgrMBFDig4fFRUR1WyFLYzNlddrsYsAvvLYz
EZFXWnyRi6Uxi0z5oXryBtEqivRaUaZvcQX0k00N/235pbw3CwggkWUR/eu92rbU
3eCmaKYIEge0l8ac0gQokyRd35nXzyYo+0jm4xw04oLKGHUgZIXZEB4Y4bxgRUfK
sf9Ows9wrqqZ5jtERqHybjRcmMEkItr1D8DJnISGZEhfAf+qchJMWxq/9MMBOcV4
XB5Mu0+CJo4jOO98jJMFY2Rnof6iwOB/rK1e0b8UXig70WKHW8DVGQzsT9gGUOI7
W337tLzeVy4+eh7xVvxL0ucnOzQKkzFRuNnYNffEI9EaJ3Z/Uekng2GKvlFfWc+D
FZDRh7643RoQoVjFNrxxq/ILDNNoJetjaPjn9SSyJ1I=
`protect END_PROTECTED
