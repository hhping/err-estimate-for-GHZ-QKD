`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7kwa0YZaqArygzsmkHZj302YtDM2Jz2E6nfjroc/AF1b7L0x5RZ2NJlLkw1FCmv+
uiSURNU2iNFiddw/v50zPqKhD55ejFlUoJMbPEDwfJlBzBmw3Ljwp9uKJRvONvqN
QuGI+kqU/aZ8+rtRN77rEE1saQgcq/OfDOxXKSGr06OZKTQoVOcT84Y6xgVfDfig
8I4eLbeVK4A/0Dm49VO5wjgq5wVYhYm0FVFrIyqm8OjhCcTFJaIA3tdHaGNjsu1c
g8+jIjsQPkxaWPLgKQPOT44ECaE35wVEfSxbxXrZ+D6h52kK/mLTf7Pdqj29fW96
pauxNzbJLeea858g3BzegpXA0aHGHvyURmFLlKTexF1HeGl5FFkbJg5oQTBlZVbT
TKPCKr51YxBZh/g4Xgg7EP5/OcWIC7W7PvFnzkgyIuxhh4F0nbtPW/acPhv4Bgf9
D717A3rxKoocVGkF7VCzt7+q0Mzs4/uftEfb6SB14UmA1Gh40ViinkRq/2ANrbbV
RA8YeuSqS9/k3wJpL610fwncrtyqaVPDP9anJiyD1lepXj00/HyV8a+CzFOoxJ1j
UAa0BnbWdAeUJC9mveQjUNtTADsv++Zp7FfNID3QrdU=
`protect END_PROTECTED
