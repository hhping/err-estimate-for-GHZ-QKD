`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Egc5PqKxZO8jClJh7UEa/2MNKF84MpQfrVTC8cPKrbHxV1sLAI2pIbQNzcvEP6LU
QqsaS6H/Mn1aca6LuaNnHKFROXdTz+O7dTURwmueloI8/wLcvNXNoQx50wAI0IK9
jHFIJYiTciVFiq9I9Ut/qsrB9ePXrfvOca+s+uQZHZyDHGi4Jr066kiPASdVaTDe
+fRatiHNJctrLx/n5uwq1/5R7AQA0UBd8zhKDF3Iaxb65Qz9VF78a0M4qhoO7yHI
gfBjsQ3rgIADUUb+UsrBYArIkd88yI6rYpzazop5x1tfHD3SLVx4P3vbfc8w11uc
AHqKlVLTLKLuannkLyEoaTE4YSjMg7hgYFMDtb4MmkiXlPNz0kVaQwuiwGB3IITq
qosBBIzWxpEkYowk+ovwZd686cqkBwC+tb5YpWsljnd66FbUHE2DC/9JliyH7Pww
/N2LD93F0UUJF9Dpj1HjP0I+5eZ98fiDlUTm3GYm+6sQ9+Z7YWf64zWT94slzllg
5UhrBB0ePMURVrxHJFhrFg+FdhCPLKKVcYGzOrI77iyIv1EfdPTmEGYMbAKzkERi
8jzkLhe9vcJAGkNwsCcAI4GlIFHzPUbV6dc5QgIWDeK5IcWfr9Gop+Qq1eUk3/db
F7gRoglMHQ4LJKq2v6XAGgfcXPV+NlFbccceSu2mAJMPhXTdm+OS6UUpncySIuTZ
`protect END_PROTECTED
