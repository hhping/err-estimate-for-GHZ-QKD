`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+pcOQ1HScsGsBY9EArUv5WqbjNDT2V9G0CFG97vSo2vyu/3ULScyRPoE2VXDDokM
TwyM4N36In66cQROeaKnIhgeOE2dJydw/cAtRtfE54fuFdQwwsDESRbUQ/H+uDQO
W3rd75YkFpZePxqShhrHdZNmjMCOLWbNzXx4MCAd6gUjRxm02Fncke1u18H6cvHV
DtcaTLDUUeULI1U2YKN4U4/PX73seOvS/HZuFbNBSnRue+xw+8ffXoedZnBNbOC4
kK3PN1mFJLxkZk1MGj2PjldAHVGZX/lBIWdljhVa7N58xRYpUj/mXO74Zyl/krWM
WSLIk+lpq1xVROL+CQouXASVM5ljKe8GCHGV01HkhYVSspGEW58Jfj8q4+hbyTOe
2DaTOocyj7HWDx9FHrldFgImEWGiMmgWBTR4u/0DNzSVSqpOPa8wNNIPB8a0AmHg
cc6EKAJHdFEX7nbF+yMZbiMpHFKe6G+PxqUNN+1FAhzATwWpROXEgL9U8LCmZsDV
2Kv0l72KGrNjcORpvDkeYCTNaPsEdadvwfDXSNPM7j06vVInFD3Pq8O+ZaS67m4z
CthMHdo3AnjWhv9FZ5C1h/dXdLrhXkkS4E4/Co9/1hCekHoXlV4oitsATIIv+acJ
xgx9aCQdI7pp7NSSsCHLOh4A5uSlctYtKLV9FdS79LknsgtlmnqPUzA6Sl79pfLb
Qh+k7eh/E8J7Z29xOiP6+auKnS5K5TYsZHmHRLNh/7ROvZltmOdjHB681/upHarx
TzqRLMY11NtpGms+jiJSGkNN7oRsd1KnleyWAK5AqKgQ2gtnA3g+2VvrsoovROdd
Fd9ZXoh/EQ0yfzfvvMYK7Kn8uKE8HioaCUv1Hnoc2Mm4cdUmX7hJaZJ4ffvmYpcQ
qZESfFYFe66Pac09Ak/0F/gOCeJXNkXwd1R3kUXQZ93mowg5+6FcII7Me8S3DvPj
x6GqnZdRKpVNqMWVxDbeK29JuoZ84Ub1wljYfikW4zTzC7/C2+z0YvVeKf7g3XpY
zsmrMJYmX6dRgmkRuNCARakHHL11ejqdawoieiv+sQpupU0wwA06ngFwg0Z+1f4h
ZIdn/+VTVkBqd2BQyVSd/w==
`protect END_PROTECTED
