`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F0auVs9qWmlhHvMcGjUGuyWlvVBkSKUkQg3RhU0U1xEpfqlsg+1dFfSYdv/9gEt/
6OESW5Vbb2Z+qpt/apZ/sA6bvdWHicxSYkBywxxJz4cIC0U/qQAUz/tyB7T/K8t8
k6R2k5B2vdD7pvQ8qRGThshEG+5a0Rdii1wyg6Tw2DmiRgw8mXW6n74vtvHmwFQ6
1NrG1tpyxctdSzYdOTMwVzH6I16DTE2KYzwjBaOa5bxVkZPFfAAnfIZl4hTHF4c3
eDhCGjyuN2liOe5CrpZcTnJAoerdmxorS33wWI/1Sr4eKhqXBlzunVANEZTDI8wv
tkVkObu/Etg8KTLRdyiqVR2DWP2ZJtBpM1bYbyXrhYOeuj2hi7Pqylg5dure/nD2
EXP3UE8RB4vAkl+3rK3LEZ5Mk63UPO9AlkUEvHaZXJiIMdN1brnfcXFtneM6xvw1
XLOjN6iI6F4oRLR6te0GZ6+X7E2gU8GgWF/F4+oZnVBDb/ZbAXp2E8WOGy5saQga
VQGf1B99y/xFeiK4A7OO8ZDG9oQgQ0vRxznPf4Rj4TMBghZ0g7DxaxM6g04yFA+k
odmuuRAa9Negds9R1vIxwEHBZdS18WbQ8wDTfdFxPhqyZIqs4Oro+IETFF7u819V
7l6WoaJ3keF1F0SYfa70IaBA5xQx780/TQKoqRVIIp6Jjl9Y5NSEu2bdUeEi/3EZ
CggmsyutDogKP/jdXB0d2fv0XfHe1jGPjnuyhP+y28iPhVO0YqyQ+Y0UIAHZmkMR
5PEq7bWuy4dNbwL0nZfaTDYzCI2Z5dxOD+X791ky6C4NDQ85AL0wdiONAzBP4lum
Tst7BFStub+TL2mhzw9qmxPM/3xrVuQx1HWtfLjOHci0rXStXnQY5Ma3oDbI2N6q
omFv5VEGRFpZjt9Ltt0hiKimfVxWfdROlpqb7WvSK7txhOFifvjn21iTZfoORODs
xYh3kucnt+YvW/hYNiOZ5FEPIMJewIfi585W1imC0h7yzorOl3phbrhv2Y1qqXFJ
bmIEEy1uObeoih5CEKhVnySUHC9kwupI/4tsdlKM6oLYgXVxkRIypCvSVTLOf41p
20c7Ku/NKlkSZMA+SrigtJaLBLGgXSqOG+pgRJvoqe5n1vbUNx99j/EUMqNRE6j6
5P2OqKB53/YMxuGbcPcLK2hwXQfsMLXTq+WPTRe+P6H1ahK5aBsrGMabF3DRfgF+
TpWyE1dTGG7614XHmRapInelpcOEhhy+fLdfPEoiasSFu6EKrXSVduitlTj6iV/N
yDzk+3v9OxgsKM1/EGDBAqazQBdWSXJ7cDmRvY59K/7uHzno2JuiJxS4BdCxqQ3B
LuyfSlH1ceEg9Ao7brT/C3UkNKOwEKFXUZE8SZD1pLbh6xwZqWVNRlHgZ1j4z+a/
qdLC4IFhBl9hJVvLcXb/sCEWNDIu7adjsf4hC0WeCeTHkQwleLgzqwa9BrBOX4gS
6P/u0iUpMlCntEBOPVZyw0fFyp85yU7SKlsR8u4fDQ7kTeSHrsd8Q7YG+zaiZwCz
YH2px5tGkEEW0HKO7lbrwSjgp3F13KWpOzNJjRdmV2KuTZ7AReitcDtLwSeyifJI
r4Uc96VkA0QQHXvzk6FWNeGG7sYSDuJnMJJtOk+pt4UHaS8HWx8r4R6FIjZglmGD
/YPSL9u4FJ5kfxJi254Hdu5TsFVuunmaJMWhQQjRgWXD3UI0DXTaOwx3dg1myxYs
Q1bZHTUDKMLzt+nq5qJA70iNFi2/ZnR8P+tCeEZhBMvInQ3WkZlDK1qgFic0nEu8
1foHY5iJJCZZIuqTHBHOgatoz4mD9Wbn03xQjCz6S23LroS3hfRar8CzVxIjfwBO
ttnO970JdyJmB+QIS+xfZhnrL4RF4SpL1Lsr7o+JUjPZRB8OnHoNn2xEEFTB7dXU
b7hBxyXeQxh875GLtXo394GtRilgvBy6SjFYXexp5/4h9htK3UNOiVqkmbBqXwLN
/fC11duAfIpT/QApz2P2TwyqlDgFz7ZfJ7ovDKFiuuJGzh91wgvYMMO7lZUVJO4e
MptsE8nfal6Qw7AqZ65f+9vYUvnpwf+5wXMSRSejDyaQZukxN1WVAoQQ4cQIA4FE
hoYTQrtTz+WygwBgCSWFEr0UFGJBlDv2bMgVapVmzagil2skVKQIeSMdlgkqoakM
aV9HLIUaBppDVuZl14nqEfRsgR5b+otrXZUo2jO8mi+JtKYoM3Qz8aiPF1dv6dkb
2stq9Y8gNU58V5qb3kWHwazS9UGptXPES04TT9s4fzkOFSBoaEEofIMkfjG3/1yw
px9zuxPWvUx8svQNaVzRro4PYZrbrxKClt9RD97lL+ga+ZPkPm3MQzr8zN38C1Cn
rp6hNkBpTO/hEMpFBd6ltfwINTVacwG58X/d9pO7+k9s6QHw+lnkb3NzAb8id27j
3ia4LXvnPgSqac34dtgUYE5jQWd544ooWh0ggGqH6AGGb5qjRAPJdKiFdTWa+vOv
PtmXP/MzGeBAWVC+7Ut5YLUxi2nxFKAsBjpQNEIXR4VoIirvMV6KpHiI+qYjqNvC
dcCepEqvgf5SttpaIPjXlOi03oprdewTs7gNz9tWL+VYx4ZucwNG9ouPNf0ESSj1
THRxP/e73LaFWg2VXuOQtx2AfyZFfc6D1SorTp+NnzD/VcPiD/JUqb5t0TNb8/+L
xCpaxNHY/V0QWMQ9NPgl/iqLuY+bfEZ+QJg3CqouVpU8xQpEbBG94GXG2qB2A6er
wMiGMhSQx6kAfoaOWq8rvSz8RKNtpto2Jddxfhny9Mj9eyxQfD5CHkDDVFEMvL9+
sEymE+F5xNrLrH4iTkaGIBHTbopp4SweYb7B3OJCPun8g3KkkYwF7vMB+Tu4zN/p
/DvTSvY66m/jrWpYxgZ19rEuNUviHV1qXz1CSUtD9v4gQ9ikNlHBpWqgChwdJK0J
6ZOcf/lQVHJ14bgsTnacPfFlsG0MMFTKNGlOa7/ryvmFyXANHVeuDG5VBDCbhGKJ
RQizc8+sGWl0H/dtFC/L+rBpOiCBP0hCo05EXmp/J9drFeQ+IVnTlYMPJaoMwJxo
zwI+gmuCb7NLR0RTs6lbmb/yyizyaVRoRJoZNzFeQz/y3YVnaEc3bLieTe1pMwCw
yW9AQ4E9Uy0ccX/ufj7kj0ZHmOP2JCuSXccnj2xQK9897v41UVG8xfdhGCBq0+/E
6s6wlZXBGGxCd0BE+OZAaasPR8lJGNZUoW4mWXAyniMgennt3rSe/1hDn23UCJVG
nfaJUOOerIKTryfoz1E4qATYHYVMR/7te11TKlSZqQe6igE/mX1CaHi3nyQbpkN6
LE8HbjI9NvfO1f58eNNj1csPrbwRqInCUSQqhTJydKDkrWR/qsKh63TPhHgz2LlQ
uPpZzDhAldVtXmi3NdMrC5W9kxLhzqX2aeqggYA/96blcm+DB2GpyW3+GCbmdCWs
OKf3ZbsudrfnGtHQy7rIx3euXLzsvzVmgX2EbSurGUaYgnldzG3kjt2dssOXiffT
5kDlw+/lK1LNmlkSOVN8wm0LPZx7OCwCY1+Jp/33vA53yZEtlt2UwTpvPpGEyQdF
DfbAuMVR2Z64Qq22kO3Q9ndLbbl/IVGkyUKI1PUXwSeAW4R4avN04NSo8ehi8fst
TBi34676BXIPn9eoZ2+mUovlC1nFzYCpufX/gvIWRRBAwJWthPFdtPgxB/KXWOPD
0ruqHOKrbwgb9a1+UkFPI2v36j63KAopuSmmT9fUuG9nVU8GD7ZjIZww9/mv4cZ4
HHTa9mYER33IXZjbd5ayblOBzndO/1Xx1hANks/9WUFgAe8mpdlye1HiQpWl7A+c
3ijQeavFwJp7OniH5Z/hGsTk7bpnyn6eOS3R2YFvriDGSWAIw9Eg1LFxHptiGdcK
fZPo1T/GZXL0Zmcgn4Vtc9obIx3KBmumneDPDXmBzXA6o0ie2TJEDC+aDSVUepLX
vGO2iSLvGcdci3EvTOwp6RP74IIoAyptYqin/Tt6zNYlCcPnlz6nfOuJrQAsXLqh
Q3PatpDIMbzfBatugA2UHkopgGvaSCcLovXLuzSPc5pE5804/K0jOgQolDNb0lY7
n44VgDmJztjn91/2jDgtZ0lEa5KzeDgg+yrQGhjQVpxcG9ve1WDd40P6K1NToXtO
f59+8dPcbPwbo85FzZJgwcpy6yY6/cW9LxZHs6TNQGsD1h3Kb5DhGiSlS6XL8kIZ
hjtJXe0J7UIq/F5EDVqTrx6Bz6U8z9OuOUHYx5SQcc52vLvSkU6hwev2iBSTCdyu
h+MQWoUci9slrH/vkBo3Utz+GOOMTvzz7+13la2wMHB50NgOi8vDdm6o68BRypWo
0UjgxjAF4d4G37tTu64m+o/+OWRcSeOgZUcTepx6emJ/3wKCK4L8vxrzdvUWRYob
0cMlS5Q/ojvPx3esJ+dyAAeDPdHdziJc2iLejEWp71dlCZ4uOA39r2bDbD16NMaW
EC3lcUZVzdmVxsdKUgNeD7vZNhr5+IDOcUJ2ZDq5Qbya3s7J5sV4Gd17CPXD74IS
rl7Qlu3oxeFkln5OyKSitkOUsL8N7hczjfMA3f7E8AWD58icyrPGoLipQoJZJaC5
9Pd1nznmWLN2v0TRcdVD1mfik5ls6gDtUl9ZOkeGXeHq06y+i1r1fLtTouAlSyxs
Pihgfu616DuXJxbnhL6RNpJnISveWgf+iOatdrRSHD/FyFZjRgHbuuVXBFGbnTjx
VkJNgHE0CPpDyLSs34aSwAX8Iy7G8LglgfsjFoJB1+I/1pNy/UHteVCcEeREdnKr
4eOjW7zbOhhugS4ul/PcSbfilR1bswAklxOCoXwGc7k+7U4czQdIIQws96roe9Ht
xvZ60OZWC2woJwzh2aQg4ExvRXl0wYdiImZZFK+nlKwtSMJM412reaJdwoGmdGDF
AECBdQ04WriDmhCaqpokK1hpWqz7S4GP9ZiqtgB9dDh7Z+sMfmoQFUT/EVw7yvDL
5A+wx/THd+a92AzufrDH1hWGz2e0SCZ+5XeavJT+Rj4CQ/P8ekGSTaEM0wbOIKdL
HhG4Iy2CucaJX2I/A+YxexVQ/J71DmIm6tnHzSCngtNnbKXlvvd7Yxnw9p/e9+s/
xGGsZXIj3+Yn9rOuT8jlQRBeu3tUPhcQxT8gNpNAJVDqiS5ZokKKPodF74acLd7r
mFcUrIoeJPnQMqHPppkjxBqttJyUIy2C3WBdRQ6ZL1tSrLHAb4G6FnMtTO2qhmyb
7QAmvPnG7XvKdRq/HcvWqbp6XeUUw0q1qcit6IBtvh+Y8ySj30SFzln9SvtKfqrH
pMn7qJ0gwHbWLY1gt/w+AkDo7uKnHFVQpunm2EuBArWpuZB9TunBptM6W9ZPHlhN
lCp6Al7e1h8Tns3tiZTbuzAhxhgyfE+HV6vaz8u9PmZUNwzNZfPTiSb/N5KZwl1R
3LEqAuDNZgyEIcv9yQp1n+R0H4OoYj58UmX13hB7SL0YTL31CqOv5/fISCmQ45yX
6Yf/HjhCjFFL0k9Hee5ivq7f5643Zg4gG0SjTyXkvdLQC5WzojMxHwvm9/11AQkv
u7XWhDB0WepYFEeFZn7JNGiM0oilgOYhxNoxfcc1nR97SwU68oYWkBPSNMmsOnyV
J5EiF/cnqrtibmmmkUs2AanJE8laZ/rXbQzulmOd2pqUzBcZrvtaoqdDAY/hX0vC
zVEmkF5dib3Ib2k5ZekR2c/H8PssN5Ot3uvZ6/esC2YoYNGOiuzR+cCKNBifXA/K
GQxZFj5hRABMPWJFD9xBlkaozMm3sJa5T3CVx9ZoN7QTvVoSqHPm1DEt2NswVa78
WPd2IijFNFLplOSeYjR1U2Pk2QwYVCxewqQr2H6iPh7lQXPdS1EW+77kRrfp8I+I
XxNDxwFFTnaut+joMiPicvTxFeSU5rL/HCdKu6a/imUJKiylN8/9WOH+7kSTanC4
12TODUHIq0O1RmSNSVK6D7ZS9io9f2uusvo9BE4SuDuDMVq6QRIZlZEoHsfwaBKq
W2JX31eL2zVR7b29ncrujrLIeHwtZ82MIj9yh7YvSJSUAhycJcM6eqZym3xhHAh8
O1LXdIJA9qZQdSgVullzZ0D4F29KvqvZkUddkR2i9ln9OoeeZyJsHRC9czkHQPZw
OvhoP5jx7Y+qOaeebRicqzATDI9ZS25QwCUfckru3mQEGwxKqT5JZJqiVnzoOIwn
9ZE47aVJww5ozq+gbTnxkbsRs8rq0FttcuRVTUSEHYQKLXXAl6g9nmJK55Y6ZruL
T0/Vgc8bfH1o/90eJehoAPBzVGhMYzMWt9w6TI1MVg3sPzLyokQ2VV02I8FVtEeF
PEvYb2FuDxmMZkdfBk7g+tjC+LYBEXMof6/Z41aYHAXDlNbfZw/PT6ff2XTtb4td
Ifg093abeg6L3p8+dm7JtKvXP6CqTl5Q9c4rhBKwibgD//LrcCOkW+3TkLJ0r4GW
riLNf+aBx4Fm5TOXQGBs/tpPy+YXoSH3V6jML787/aVPU+gbNZV9dYwRx6PT1o71
1s8SDBx16e6BZ/jICpf28ctxlJwLQg2KxGfxpyjd1Rbv5mFrqQVs3ZV5h9Gb46ah
LpWR87aO3X+j7vG0FhLZghSOhHrh1hxFgS2sNfXuoqKijVYdjIIXqCoJWjJ4V+nk
EUk/L4eBdK8MwYbtIkqoqwGbBLZS4F8yKpwmvauxgXCTmitS3rgx3o1ZWxp6+mwk
BN6gfNhaEwWzTbDTWofYyWYNaDz7FgMmX+HupNf+U18Ds4Igfc7UXt347uJGWu93
xnh5nB1QcnBBZWdx8gR+xii/CJCnACG5+nxE7VKrey1t/RedaOQ9l0hT1saJKlTy
s4jMrYBMrSv/Mx4YUwmoiFY19TR2Gt7gAcF6p6hanIVLKHfofySYk+wi87dvkb72
WGlfEzEiaHxh42H8B+A5bJ012fAuqvTOmal3It4DynokVcE7n7xLx7IJoA0q3hBv
OL7HvusipBuHHh+VzOesv9BC7wJxFcMRwBDZqvQ+r1jE/wdp4zK+PWfh8hzhRMkf
oNOt9Jk2zffjj1VeVYSR4trBTsOfdai+aM1nqsilrpEEqdtRF3IShYz+pVL+hWdX
mtFqLs5AP9PKaymqmeBCs/aaGgR+wNoHTW8xGAA9ZPa8QmJO1iYzHznTK7WTpenE
+hP5wsdTy0sh4u1RpRgvF1RIXz/dNb/bBdY+7vjjaAnzZ8iHywTt9gucE+Sat4kD
B/1AZTq7SOuaAqFj6Rhy9G3JguaP4YSBhxv7JndE3Fnfvly7+E3VMYNiV1HBkis8
oeABswsxiwPgheJoR4EV9ykWRNBiSG1k7uHJoCpwkWJBBAhxsqM0lowneug4mDnc
wUqBqAF8XbzKU3YuB5ZJ5+t+Iu8AA1Si90CCG16MLA49uhY0ycpIiBAaunIUewEP
fyDqm4jiiZAwccuf93ioA1ZFy5eX2AO1qyvLyWy6umXC1N7gthLz48ZtmieA/wSY
puV/NRpjf2KT4WYyxzptkZT7u8REOsuF8SEK184NyLpMZ9hnnGcKa/lS+sDlQJPF
0gQZwZN3o9P1JQFHnT2gIwMXeFrsEkBvG6xv89/Pt23YYaqwZ9ELJAND2lSuLqZU
bKkDD2QCMg4UfTk0cPJlefWV2Nb/xaC8/x9to7njangSIgiGk15FckfmLa5Midk1
8diGrYvqUjtj7/BpdZbmBszkoDxk0xmQQh6SGednKa67sCBBv+NslEW7ByH0asHS
/upusJWIZ+zgVY/CoE94lTnYO8W6LBIfa4pKcoLi2wGVUPsJAoCSwumHZZYiEUdr
SMvkwze6yVDYnBsVJ3n5P2jIsLq/E9DClwgsJUP3dN5SelzElyJX9LoHr2mleXkr
kFKSCZjE80ZmEqa+q/qDQmhHV5QrqTxVj0ODv+B5ZW+ybAeH6nFuAykR3FYgCDus
IMyToEGkL3moj1Vov7cq10Q81Bg9bFkpoEzDniv+r7wBJGGCKuZGAv6P2wa7iYwS
QxFxs3JzIAyw4rmvMfbBBFjnqFKAs2mVd+N1Tb1fo8TVBTtAZuPXKR4ccbsekrS+
mqEXxtp+AngiBX09aD/3zfpn/SWXwEI0lZNdnR+RO4DJ1WIRVxt0CnZo4jRZ700u
W8A2F3rEM3j1skoijxsK2yWEHFv+eQjDtqw+kon4CYNn1NRbCA5r0B06MZzu4vcs
WQrhwRLzmuNmOj95Jb6bpRU94KjzBU5Vkxjd8PIo3j5gGciq8puW62l4HV/l/HYO
zKaN2KEk4DoMyHra0bykB6lb0/SapmNZ5WUHd03rEe3zITYs7kXg57p9zrlwFKps
j0lSi5nQwdsdbNWLtn5X1tj0+6SsIio5iy3mYsb32eniQXkhnLLnIrcV15yzRtnG
PLC8rh0HSBqQSSvpU/SLGLJVemteQXMD8JXhnJSuCmoYkET1R605HQzz4wsm/cB4
9OKLB5St/6cjiDFMdqGP3h0U4OHnQhLENVAM8GCoE5YsmOvj94uJbhliDjegva8u
lOF2wyQepbYRQrnZavHE/JPitlYGweHpnyU8Ct/l61UyttpmNAItXKsznsUY2Hvk
Xrt/8YKwszSgc1FQCEDOHsimDT5XJdvUzpjNK9lR6TLPtMinGYNXJoqvUwUsy8C7
lMheuijhowhIWGiYrsp/FoTr05gOWzAjMw6ZgaAsBw12tCkpVwToY9gzNPlt3Fo0
YP4VgnIJSYsWuDn5O9DQBwEiWBc6d22/+dPsGsyOn0L76jNEvuRETou1TvfLFLju
ExjrIsrpTdQ7StjL4APsGOrbMoCnzWRKZXZns8sRo0WfCxqc/RLcIxK65gDrjX6R
3VJLUC9rv2AIYTGDxB277mWIy6ga5E/40ppqdDn3JYbJlJyxvuKkK1BJh2ZqfX5v
PZ/NzqWWWpik/4CTEfcLijFjbZlGDm4kg/o02vXHGKd/UEQ0GMrMkZP9NNnuARtw
Sdr8mOvqIcYG+E+fp/R3/mUOgM10pHxtKcjupv9VRqhZnRk+CIRxky0Bcq1fcuMs
u9e3UM9KOptBH98jjRfT7ULw8TWzWFynt5omF2Xa+xJq7VqELoA4vVwswci3JoVu
sk6P3y05RXBbNapLX7usGltRAyS9YSc5fq4IEd5foeVzwzIQxeItqPO+t5kR3T5t
2alyf1/9aQX8NSkqgvf4AFsRYCj2ipBvsTUPPIIAzrvS/7M3thQBMnLVhyyjJOEj
6v5rjyaLlsI9Iuf9X5tLu7Ima0KUsJfOxMdRTcZUfKq2ZBoG/jZJaBgz4ee5Aj7S
jC5wz3E44kR4In6ogZcKFmcD+3NVzSxID3dcO5992xw1wpFjlhlWkz2IcFXCrP9D
vbvO4ajtNMbRTK2IWRNdl6Tj61uWCWArIxlxpDrejWbWkKMnES6mtNjCxuBXzjGO
JThr5DAcdBRdi7bySDM0b69oOAG2gIPqQM7gZnpMm8znvDJ8aeMYgO7ZJUmddzvN
3uJBJ9SnOyXHwyhVnRgGReiqnBrQV+vPZnGX3LaCJhxNIfhtT05AxVXACdjixUCn
7gN/FNhb4bzxtmoSR2RWmGcqAfQUoZEywmtdcMuT+GmmMiQQSvAogjhjVp+mvAI6
UuPGe3bwAp0fAqdZCR/DaeqE3W9IH26hFTw1UdyFVi5raW04hzTyySVhmw52x6ah
YlGRo174w4IfgPEKyahiAv/I8+ST5yTbJe6nifgyD1k+nAl0jW+Hl8gEyinJ5kXK
fYc9OsveBHGNWuUG1nS+qyi4MeQn9SaHQjGb9wCjnEYgvePPsjs0MDpY3FPEB2/9
onNxKsKs1wrR3kXiPusQVMh2AQj5qKmJkYIxshR/dlmY7SUkL8oAGsrldJVllH2y
9x5umrYgNDvZRv2/sRJBfHdCU+llwJP8w62MXWisy4iGf7LpuSueCCsgsMLeouhk
z4mjvQxwyexRs0WChG6fgqNOT7EUTAAwa95qF/DeY8IfsVYMtorxvoutL/73xXb0
O+U2MjKeySm4YVIeVB8fUyHBLzOVlzRcBeY8NSmh+q331ksaxPjCjInErIsMERtP
FQ+HREI0PGCX1VNalunj6KjGWgUj2ZHRD5WA99dapjsuZULEPnkn5DyubUM7rERO
p6v9XHVeLKBpZJwlx9iNBKu11hTFde4MjreZ++rCRJSRADlI/PQeAi55KtNvNeOe
6trL8fW97ramprlR4ZmLw++XCsCIqNCJ3pGQoMUYjeUtGUvsLXpCcItwfBh6kBXP
9SdOP67c9Bi95ZNRHvuu0sfhB/vON4chHsI06FkIIffWflFIKE3KlWBo1SP4Ar++
SyEaltyt1Kv550mT9V3/6QcXg/RSLUOxHebgDGO5Uqk12KUWDSGqHGKORS1TcAWk
NMknoN0jPqk68vV7Np8gMkJQHSxdZAfNYvagzO4ecmsdp/nBS5Es3kPQKEL2ruUU
rOvgJZoffyykRBZL+JP6D3PG9rIPwsW4PM7CfbK9rNlrF4pdDk6l1x7P9Q9Cn62R
5p84WoppQZd9iePN8WKDKpOyZJjGnl+zPUn0pDp9JWxhbmdpGRCcSqIeHgW/G0nk
isPtaR/VujhshqmI76KLaz8mRVVJMTY40wFfZGBFrpmtebt8H/pFk82DbkU1fgrc
0AMwIs/wojxYwdaV8hLPnlH9/cm8IHTXG+Vi11ue85aohkB/SlicabPtrnvtBJMB
0Wl6+YbtvQJQHMWockQdeNL9qMEYvXg04Gg0UEIYY7nfh0eIDgDTS69bblC3ISpQ
KgV1PcJi+DK1cIOriLcll5ZO3ipbe74fz/zL73i4nENjSwmbo+q1Uuyqyshc5Uzb
LJG1AwN6JcYabGovADyU04qi2yUcx8mUTl5/1FfcRYPXaxHCwQHuW7DooLM17FUd
HzFGOCX+PbMbQBJ8RS3AapvEbI4WelYSsXjqp8be41V/aXEr4JD1K8CI2NB12jP8
DXn0o8Vr8JMe87/ee5tm/9T6ouTBHTtHVuo6dhWmi4DtzjprgVgl+rjdUDDnVYFI
xt9nImG5T92jmxZJFLyUmSjo/FQ/ebIEls4aG3qFqZdRyfCgkHpz1ziQvoFFcSpQ
jfynYr5xqNYTtMls2YQVaKo/a4iq4jj2H1lul3KguZjxW1Y3Mp7UVQXUx402c9eX
y1rF+EtI1Br1f80B0r9G7n5acfDXLFj4HpKGqFOTq/0j+7yPjSxohf0fNx3bXJW6
vnJd/eOMinZXd07t51J/o/YRPl9K2U/A/PKwDAR9iAgO68gw0a6n+r1VVC3df4NV
tKuw6xYhQfnArtZA9eq/JL1Rw4GkgAAvQidmwSToed6ikiSkgvxYU8EUuRRpmMxP
BuiQZJJsOTFmI3Adci8FEIcfcU2ioM6JLFXZikt+S3EXQsE4lRNstogEK1hkEbeg
QtGMfFQgYV+O4DtY1y7oUVTyR3jhf6bhm9aLNwG1eQi+65Gxmbm/k8f8Pppr6WGo
uYThPFjoKAZXLFgrLnWlNVJvAHvLdCRnyfHha2qjIfoWfh7m+uvpLDZ09BJb0uKX
/Xa5HmBoQ8Jkiqx9AAVCqjUUVvws0vHB54A83OklkiR/szjAIeInFaAXloBASAgo
q//dvKvwjryCZiIZtEZfSm94vJk1+owuscPp4Dgf1P2vpOAwQ+1VQKS34pL8mUhk
cxbqK+ojxqIQGskgzCQEPoRPmqON+KentVxW3duHkpve9qdCzfh+TNA1XWlQNHBd
0FIXmCHwkyigHBf79AwmzTYt0uJ0jsfyrSCWGeD2lgd0a1lF14yUMNiDDOgzShyM
8qwN05VHkBwzTQjiIiSNRkGRHet71tVQJJIypfH7de7Hra2TPXvIANUL9Cq/o8Nx
x+eVUjMOZUhJhAS/nrFPDJ/wLTntGREE1SKV3NeLV81J8K0ddcpNTrR2qyFzfKFy
U9Q6JISCXoiKeFGvQMAWaCGK9zSh2yYbD+BojLfzyGXDaCPPcmKUScd9oLWcOnur
mOJrCJRY/ANVKv5snS/eaUmfB1V70gfnSLv13hSw7omqU7QaGU4+1CqRYsrYi+wr
JF+jC5h9tgxpNQGlnOd/T4xF45x+c9VFmWPDOFbZz691g2NoKzd34WBB0+b+xjx2
0z3TRCz1yy+NZGZIBKw+yfR/hMCRBZlO056+dLMsYDHAVbjs5f90TERLepjdP56c
xvEl6UY2la2degOT5oKqGtLMBMVQutmer19DMYaOPzbqCZZvPBmjcJ67qSSYSrS/
+eGptARvPghLd0MvU4s3rR164/dCW7Tss098LxnBeTmGnddQJ+9twDXvP85KTymo
1e19uE2nuOlkenGLVGaEFadbGRqQwEMWUxk4VEbM54RNCMDVePgEiqa7U7jiTutS
XOr9xFP7KMCXAwA0LlEc8ofd2K5G6ZUwAdONXmPYWP2z32N6/A7tNQUDNzBwig0X
VrmSTaLCz55QWHn2lF8QRtgHPKK3yecJzZM8q9cionAPGY/nIsazAZI1xA7kQuRf
c8l1ApSfWaZT9rbIU2mqt+eE57xGGe/pAJ9oqXqv+Y2ybPFBnZi3Wm0neMEj2cho
nOK854m+LvhkziL+5ji0s3f9GLmivj1e9Hv3/NASIyCpXS+PQd7XUVvN+R48jG5z
/nndb6pD3XlchGpndgV0ONhtHcSF4rOIa5Y28YtbbUdnO1rWUsnSQ3uZg3gnSY6J
5hsaTyBksGjHy8wnvsIv7Fx1Bz1OdRRA24gb99qp4aMAGFZYyjcOG01m4OFSd8xM
MyA3FetlHUxkGr3VGVnJqF376Tqz686dUtl8WlrWeAngl2GWDiB6CLgJG0ZnrS+s
ZjDCJsWLEi58BT2xkg8KC3ief7tB4WYbeKomg5knc4vdYbUBnIUBU6uVyyIAKhZW
4ytazrwFIIvkQ8voDOuU5XkERCKw5T4DqQ98v3XZDUAcqDzmR6LpL7DO0Axydq1c
8NMbkyfl8FMfG5PBKmkbI5BRXesEGEyOzDkyyCYdHlcypDtM+/Cd/dUcz3zqwI7I
cQpAXPLaXuKwdaKFRt23X5oMKz+gKXzjR5spg9NQycO1uiytRYUOsBmruq2Sp5JI
drLWWACctU0nh3LN4dyRrJQ4mwF1nYKnsP5gNxNe1lX8Z3n2gk5alcAosIRNuVhp
6dS/dL06551JnFjOq35Y9IGd8O5D1+CF+HACX2yhPa8r2+V+ka9K1S5YMf6vRLVR
WrhzPLQCIwGnf1fGbBpz0OxcUlFgqW3Ztb9wsXbV6QBH6T3tW6/0acZWQrXj19dS
Jc4j5UGAkW6hJ8CTwKb2nj4Ex0xuV2j3/HUrETxJ7lo8kTFbovYGgBjxCjrGIv6i
yxOXZgnE+VLuQu8VEP8HJhJe7NQXpQQPGri3SRqf1T9drfCROSyp+YYvoc15P2Vc
73edSefWJ4/3+PaoF4Z5yeXYIwSndV80597ZM9fgGj94FnJjoVJecTiCGQGyCk2T
fOq1kwUXE/bHnkIVatDKxjW9u0VRhKToZ6jq91P3d2oAwTdixBKx4zoVBq9czpsT
WrdXhTYLeXFlrkMdBERSaQTNLNKrVKjVswBc+pI8NeZXxC1V4v+L5KME9qPBXF0s
RN33Cq+vC51qqyVBVaFQxfXELrNV7PMl8IY1vogMq3tQe5eyMHEQpMBUL/GHt3RM
+X+n+nHwNsdA4urAM6MyM+Xb7LqMQBdhddjxDNvArQBDEkFKWiOrNIUycGL9zuf1
IZd+tnZUpE4eMtStea+xGXojRiS6qmpOxz6RU2gOSHQW8VvVnbWYcuUZTHSLncdm
okRrE727cnDZWF3jv2ihbOquAyFNSfkUC8samfEnZ1lOtY5Nx2jYH/+z77mY5jsH
vOWQBJesNR/0GjifPD/AeMqObulime44eFT2FyvWr2yJ0Mckxuwum3x0mHX/Il9g
Nx4ES4YiPZk9GksUB4EFxUTremVZFV/mgqYwCsM/yxBIxo8+heW6YchbJy21H6zQ
lXvCvUOR9qgXljUaCwb+xDKKuhWrzfTWnDmH84xYsc5xOba6yuOOev192BOfUtwr
8teoZb6lfyc5AzpLt63Scc8lq3iUMepl3aSl4iytcPLkIhlWiWMwrRHddMk1HcYG
yvzN/RBFqbiWE9G81sZEnSTfx1aCQ6td9vLav5OCitOiDjnzPCzUnnmsk6LX99Cb
QIj5NfdMQ1jcrwpPnzakt2s2H8qhuAiF7jImf/yAnyy75GFko6sGWkGYi2A26a0d
FV77z507HGLNTISMfDtxkpJPM5lhw0clWDwufhLR8pm+SIazdnYvEe6dL1sZssTn
R2Rf/73spF0Nhr4qWlJx/dacugyhuhSrOdyrlWOfN6eEozeEkoJ8hs38tKKocpbT
Rtb18myMYy5hUA5S+DGfH6jXItO6RSPzbChWyLM9qfWebyh0d1aiOWKdEfwc+7f/
JfFDd4/+yxhvUa+IWmEFI6zjdRfKwa4ipUBSCxaufW7AW1n074R0tJouDEagov48
vgT5v/2B4eOuiaI48XS5scAWwsbJpgTJDUvZYN2BMgmixyZWUJnmvdZOroWhFBWj
/Tt71JrLkHYctUGVuBKaEGOKC+S2WHuqlXOsk4eod2o99S9kdkCk3V78povg7O6M
neTKbTdnjyKxZUs7qxiVz6NAusHgAK9hj/vAeIkstr1PLoJ5/dIlOgzWVK4DBsB/
AQcmbgc0z+nrLlNoNE96xkQt+6yWbSvJAyOoNRz4dOx9TDII+un+niksgGGmcJtR
nl+QmqvtiFLsq27jdwWSLHU+Z04JvXesTU5hTj1xZLGXJZyy5kqNC+VFwTE/YYTe
ssh7V7DZPQl1UfmcoLEE5PWo3TBYb34z9QgHHwZn+/NBOVi5n5jzQiWk6YL19ywe
VWqR4mk9JkYY1FgmtvrbKzvOIGBZB1IHBYXciPxm3xtnHf46W82tmlAcitijF+4N
DIBJYhH5ZbNX6S+PrHhckkz6xKiMQ62WP+BJu8z9tvVbJETtlpAUIVveaNyBgNrL
FOuOMMxyHN+d0OAExaTcfw6hE6oTfai+UfW1k10OaWBUI1Qut/5RNeKSOXICb/wd
BGKlcnRmLygmjJVFMS7Q8mnBK3uP1aaF+EcnrfR8FxHqcfz35vUJYMpJKrXO4gml
42Fv83ETqdqZ15qtIjv1jWLn0rBfLnC/riKLmFsjEl+bYSibFONUcggVXj1DdNgl
bF6kLFTYyqH6Ud7DQo862C+uhGOppCvYoCjWSfWAin3Wr6TD8fQbkiXl4MIte1c5
hayn+4bawINFYqRJjg0FUm8j3Q40MfD+KZ01yj6vP9jYbkAgd/MefvWKOdJjz+1D
6VsB4yQojf6HClK3JSs1wru43KOTBXTHDoh/aQZ7e7K+cvSWxSTpFD5Z/sQp5ght
fCm/2kGwZRKXKx832Qga4pfLBUp3epyuRWNTMSoHrIh2nXPRv8iuTSueZ4auhdOk
pnA3fgawXmk3ECJCWVygWECSNFFfB+7gvyyexReOd/mZlMOHW9v2njyWzaKTiV6x
riGJVW8cbxNE0noO7BlJQgwxbh74tke1QIrHgbBWdP8m9LdgOcU0kR3u+0qrxoJf
GTjoptJsY82OJd71Xsh0gRy/h9d426ta5pihybHblNqkL7f93JnutbuEFvEFraPA
1af2FFGqZc13aVPkk3PlPrptuI30ICQUf5kNAtRyZqDSTRn/f8K/PbxN6hmzuX5r
SwT3VQRbgHuGI0W8ISThjafovO3Izp6Qkcqkh6ALlJpMfaRgpYaObXqE31pRqJx1
hW4cxlYFzt+ZORW7DQujJ91zpVBogTVGflkC0cFRaL7PyHgujZNzhTZDLGj6ot4m
unFPwozBAo0pFfGflcMvwROC/XmHi5n5FrxcD8reS8y9g1NOo/dR6UNATnJx5Dkv
C5Jc5GOdtX+nSX88PSW68oXLgOcoX6/5fqPzuueGgYgsMIN49IJS1G++appsCeOt
BMUG+IzxeXun7VMipLCeOu46rSVAL6RGNbX91O9ePPJ519ztREOXWaSC0hXXBYOe
CuErO58rXlb2cSb4/lgTXcMC1Z/BrAGVobC+SNXhApKeKM/0tkz4HE21V1pv+yzd
SxTHBCrBbZqmfqErCccuqBxEFZbzUYdM2LAIALtyp7V3258kmq8Bush5PRTKn96l
37lq1SIQ6zpMGxZwQapMOcI+qjKzRdncFJkyQt62i3lhajDMNOBDTAKGicDsNplI
Y9/9q4MwhdWlEsY/EAKcssXFbZfujOc4QjJjaQDxRhsQ8RdOt2qMZF2vlb6YX7yi
PZVh7J0tPpcC+Jgp2QffGbtFXrFdKxGqChOSMAIZlZbzUtsaA1zYPV49EyXEDVf5
47i53d6H2Kr/qdZOFIFEeKw9rmhugQjP+tst5QWNLkztX9eTEcXesTMiFaBiAOlW
VrdbnGJONtyqFCg0Hs7jAP4q9SI9yNMdKuBi4SFfAvmmTe1CS5FByDT5feritwiN
RCBOzm+Ih+qtux2tmyiO2+fJ5v1t6khhE+7QOqtrSR4KDs7gwJOJVR4TSkWgFqZ6
YR+1nqsPElGe1Llq2uZV0hqDzQygb3sJT8FiueD05B3S8IO7KoYo0Oxz7+KHGoC1
qKSqNEjyxBSX/paD3JN9WwyeJOnvRfqPV/pHQ4/6UlUiDN32TjxUt/5oKoomgLPr
GjWK/C8sO4PfZytwBgcJaTYywP1vOZQsCwQxF3EgMP2ZdAaAMq/6F1VeZMOrOVnL
iae2as0d9JdqdA45tbKMr6roVco/ZDmmYlK8aAFhfBIqOePG/4kTAQDwNhxNo5PG
4iAjxjDTyS8aUQM3oa66VKSoCvtruBQL9Zm0gnt12ILH2oXEDYriMotsLprfbx3F
2/OhYN18oL8zL8ET4yD1WRDindMMuzDP3NxK86UoMBsBa5+d9nYvRID0VwosxJFA
R/H6segKNnnngB354kn75/Q3QgEZMqCuj2+7GF40IGlnT9xhqzPsvPN1oNdIcvlR
Tl44iUZ6LvBwmNDi1qX08W4w3C6LpTBdKhES5v30By8LLBg0bKeIffs1WvxopTRt
M8gNMJfqaBQAWxwNClqcFxLXbbSfFdz7GUsqZVChO8s2lt6+94Anrl14rBPgC4qy
u7qJyWCJxfDCxwhj1a5T0cP74AQLKJeRKUhdjFfBbUgNvmpLsdQCz4yXUOvtFda8
3uK79CUS5iHvMDx8QZ9Q9ftdT5urlEYtZ5rAWhbitOEN7UDgAL8S9D4Q4jGd9e6B
H8InL+je7OEDIKEMlUYcqeRb7MwHoJGFJdW7dMzturOlG3bpVmw2Sm5itwgHqEfP
eZlzSLaI2NXlspA/8bYv02rdYzLqb4YLYp3Vtk+fcboSUswjqi4iQeXBtcoL0t/0
hYbczw0TThMhjNggRBLxuqJJvgoozUicObHA0dsQSoJxrjupoveMQ50nxDBPMJ/C
Dxkl7mL3XvIay2RSSJOJcB02Ij785zL6vsh8VASo1L3TrB1v3P/d8m7k0Fmjvci4
W564tWBf0fEcz0w47vz08facGz/koQ4WtJzsrQRVzOWWXhgq7ftnzRbqQTOv+BgF
qnAOjHccllW3bFgWbO+mqqR0EDLiAWLImiWtOeMYWbjJFzASVOfUVjtM1YhFi7E1
GEpUK6y2L0ahu8GM9DnaqyAyzKXB+r5YW2nT4nnl+5aKaCDzQZJCMgvQHYUnWNBo
oTkhHolGuKs7XqmQOsZfuys+cOlifgk0jOnfBpupyql0HMVCDqDxwj+kCS34F84t
BgRRs/53uas1G1AnZMkEzxYkfa4K6U9WtUldxYlI9KmIxNM4Edh3kknx30h7SaPL
p11mT7FmYZwo6nzEVFMqjFamcs0Bf5yviv01gj1RMw5QaxBIYN4QkQYdcmmnwkVM
q70184YcNulmIZ6nhxAO0ZADi2hl+HtctW6N7YfNQijnNP60kL00YOdnBn9pG+74
WIJhqqqp3BHG0nYlOkOESLe/C+mKgQyjEt/hDVQ0W+ZpkBJG/gvMbPkS7d4sh3Ml
3wP8igAbulZnPFGhNDu9fpkZINNV27JeIo+sdVOt8/8u6NirDI5IRThj+KYRiVOR
eZjX1OPgmf+iFC1KcOcbiMwxbi6coLWCdCB0rN/C4+Jgr4NWy7endE8wlIFtmKuz
f7GNp/E75fY9cm4ruESvsmDopRpelY8she+f4fW/rWo9W4tmPySg+1wK283mhOp7
jPukx0hr3bz0fJ5MNktWrb8LHXDmXrrIHrWmDi8TzgSchTxKCEv+fYf65bHT6M+4
axm0JJlVfuqD7+gGp7n9GN6N49FqFvo8lMKM4zScCX0sHHmKitBRRVvTUKDUYBR2
+0sgRQQ9+QVBHTVlTZU5fKp2FCq/Qej1EXJywvCUDr0G+r6MdDdzet9A/yx/nJkQ
vqC1fKfCVgP5jP8PYe3VuGGc55ZIBh0d7FlIwrtjMLG4/TqJez8HEUpjsvb8VoJ8
ba6j67K+QXJlFfFVz2+FVqZf3cyTYv6WrZvsQqz947LDhZXru8NuIF2FeRVx1A9O
0pmpmm+Zoj4tm3YtyuVW8wzvRI3V7WBarAPoNYMcDWic06qkqyOrE+3Jco0gWyI0
YMb7AwqERpvX+zQ9OtBL24m/u2rMtLNDneRGHyTO92+mV7cEcW4yADnz0i8DSs1T
0/3/SRXnyPi6Vd/0pQ3055wN9T7i+rTp1EE8W9GEh41Hk4TZuYjC+AZBbqe4P8cJ
ewPXOXLABre9oKw1Fa8sGJqoTfY99pfuZ3Zb/8ldP1hBzrdf9jvaGlEmLOGFM/A2
rihWG5W+Xnxq0T7FQ1pof1sTKAC+QGXHBtm1uqnGJ1bmsaXbQkEtLuDus4Lwrwir
DziSOMF+E01CDv4mhfUfEg2/YjgbQSAD32lmT62hy2jbqsSx0CdMFB31VX4stPvG
Miv3PUdq4cxxufUYTFM8Yppw8+bb6rNhxWZtBtXLytDRWumRaWl0cdrn05JEX4TA
2M89JnHv7w3CDisCavZXtpynmee+WhRq9CfqsRK0tOG21UQOX6wAAHaO9Mhdv27I
INpmHueZpbheuE/5VTRgSJIEQMzLwkMuA7pe26osUwZOwDlwGpRYcFldwTkgfnth
DZ1lCK+8cuBj33tTZqz6JRy6CZeub7UG8OREozusHfhX0C3oZ5XUue9ZLYZ2SqOZ
8RdN15t7SGi6majqO12poczCQAT0NRzCVNfH2AN91ftc4f3QegVVb2foAM4cvxdR
NBWyP/avTdffLLx2h6CAIVJoMH2seyZmxZJIR98YdWIR/h7voANLQwwLxAeGm8kp
xBiCHcooHCR/W8zlZSpozwotzgPeTQ5lmEmSB0nTGxpKxFLmNXwwXgivDYmIVRoM
uw9vNx8q1bG5BM0TVO4NEAiI44fbg/IFvc/zOsp3UzPIObOMumWDdYF9KrEzy0vj
V3k9D8C6Z6x3k7QKPOeBfO07K9HYxDYymjCVQ2MN9JhFyeQiNPsDCyKY4VnGRPD4
XXQoOd6g7Ad5vABKhVEcD22xoOJGIKxqDS2syBFeKTsuAVfzdehsF9eG1f1c7kaA
uZtwQTFTB+Sbynec+m/OM5HSl6MRlPLlSc0CyBLs2JtEfZBeEDxZuwzeunMz011q
5c3aJbNCe72mgqDC672MYVuGtObsGFjsp7TgVO4O3KJJl6vPJacM7eViwNx6ejtV
9sh483q46lH4BlS3pS35arg3Qs0Gowl9wzKP5IFczNrMcbwDStUfewb1dJutuZ5b
RoI/nWUaLRWIyFLgIZZSK0rtQJuSv2VIs8qkAB6k9bGQ52CPbCncb8VeQ7wq+no2
WXIpF6ZqtSSWtw1aqwN5jfyNPqoBQJ57NTapxSOZOdzCEXie+Q4bKaUVgWZdWAUy
Zu70/DSaO41ixfEwv5ULOUPgPHiqT5JzbuN7TEaB7859k4d7GCruwh1CRxoO98LO
HJFFCPG/vQiI5LBrl8ee46UEKqCmhGaNdzKv2VNa0yni+72DMmweSYNBz9lThcAS
I+sjfc/qGurSzAbz/pfdNmMSnqdpHYKtYCoMLKvqEHqmaQrhMdvG57A8BKVTmP0I
FYRSErhNZEE8g0o8RHkql3mq1Np1ZXhDmMdaxY7vUr3JKBku3/IHHukIiFjf2YDV
bJJCzVPu63o2AZrUeCIX/zD7N4ms0z/KtVL4VR/S73MjWeK37RyEFzL+QdEJj3O/
XiDgxJICjuX6GiJEXnRv66MAOMQ2KS9SzShcLRpqMgl/kWjBnt2KLPlX3yPI6mI0
QfBk44ad9MKig+e2wn0Zx53XDx4NIAJrBjHy2/iaQVhVYICFKR0oB9/o4VoaJUwU
1BK92xtEJLwU3n93XW0L3Mx/BLq/BYBAZFVMwYztoBFBGyXx8CF8eAhEZWD+gzdf
VcCRw0NbcA2O30z2iIm2OYqxjmZWU30v6iWuOE1vdE7lUIUlfwp5n0cKMVSJQzvJ
X82gvhMAsYQCcdck0YetEn7P8KK/lyyGbaQkFBEFG/KAxdhgyi/BVxoZdqVk8CWh
X+faRY75QkofUw9iPRKn8jSUf8W+hORU+GdKHxlzxbOOvypjugsHE5AUDJ6mvEl+
eA06JNQKtM4UrXCvNghisYMmgRDgx1wj7hcn1cFnubdjeQjKZ7AtNDN01/UnWeAO
tc8h7dZz0esLeNg/VeFfsxPFf6Yrq9lYAkAAMaKc4RDHeDXlhpqx3ntslC4z78yi
efbKSCabqLy/otgbS8q5No/9gGbxj/6Xt0ftHUuLiyedsRmcw4INqD+pOw4qqTNa
AzmwCn4qkBH4BY39BiQ0jxpKnGGeVkYR9RBK0/BEulSHz2qSOTD8VLSnJsLYUT4v
EqSk0GsU8b8aI8DlI4fY4t/Rvojdqv+gJ5f/9vuJrrzUE/JxUi2yMwpjMplv8OyA
gxuEed6ZNozzBNpQ4FmcHDgeKVDD8rKgyHE0tMbUhQA1qXXkreqLQDzXuh59+afb
U6aVshak0HWPcmrwVsI5pEHyl+wvQKUjuaZ4ACeZlLpqYb3pOQ9Sv0dI6ZbnX9bc
rwz8vuTkWXJmFCJyjCkyd4YKU1VQhCI4rFfclLTMu9BXYXVoD5W6AGSZQUb1NgzD
AYxXJBmCmZ8keIxtqbvd3LRBUBXNUcuLaBEnEuyJ18ahd/zBPHYa37izV1VBEZlE
2jBo6nKQB6lVQbaSJ1cduzxn2RQBI5EqKgJNt8UDgKD9LsAD47QWggY7krlE9OlJ
ZlZx98kzInYGjidTowDdD6kHAl8037bcViIBQJz2JPzOXEk/rkkR9sEG3O0PnMaK
wYkXkqBtkRst5b8oeflANGAUFJkNasyvWh3aXnu1ZxEQseDtD2k3+HGOpoaNA1em
/M61PraIq5WpCGckBcfF7osNQTyuaG1uVf0PSXCqcQWqmf4Ilj3+HRFlDtqcKUAc
s1NSP+4p3Pn2vGwvoxXxa7cwjekj5VdAdczKpgFf4SrHjN0c9cJQTWywth5Hvj6B
yxerMaQAxI0IEgigYuZwiHwERI6zYP94hnfhxxe60/bZ/alOr6TovNNqgbTK5/uc
ypuZ6fkeNd9dJd5gLP0vaO0ySA/BqwDdpcdph8g3Ey/Gvu1UQyysGQmT06sDfYWK
WZgKiVi8OrQ7JtrctL6e+DejDkMg7sqHS+eYdUqgJnbdwZ264ybImKqicH/iduK2
OANPvGAxkMKunpdDPPQYGDUjnmNNMHR4xQCPH0RHSjTntyL8cmkRuzvrFIUWyKtL
9H0NkJ3DzEitcWSCShOdXjfN57XuzgQqlVlrnvwfI/QLczMug8+XVtVuSVv9l1i8
FZZLOgC5yBBvBIqmnhxk6vbjWHE51kTTNRdXlfiUlKGPSOcS6+haLblFpnzzKQkp
WPAs5tjtgmR4F+9kYrrn5jH4TfTmZpiElLjG9Tzq7JRAElJghx+3JR/koFVjBX7q
Rvu3b0zkpHuxt7//syz0hZFLqqg9JR7+RvOgsm3fbI5iAfUYNXQa9KkZOEl9eCJq
bRg3fB6YNRJZkhlwBxt9ZTHMbGKBHENxgdhkXNelCIdgn/W9OqlIkc+2QHt5fksz
+2sgccFQhvrrELU9wworYsE7DshDMvzLImXOGlciiyzTR91BS35Egy7obS6g2XJU
k95bi9N2d/2VeueZX2PqnZmwZZ6wqjefKQKW1EdL0oCHD5qsqp8WrlLsmqGCLYw/
1ZrSj/E8nVdP6FZtjlGCh+e8iYzYb10bdoaLxYLs//GmAraxS/MILPDwVJrRhWcL
LtcCCrj72JwAq1AfSA07IjAwqvI4AoUy8eg6Y+VhzwnTdNQQkAwy+f+cLsQhvNJZ
zBIx4rg2AjCUUVly5qIt0ICPhjdSdgpghzJl+WdFXrXvZoY+Ee4wXsnmo8IKF+h2
0enoRpyx5YOi1DmwNb0Xoendjlm40y8EB8cFuZUNXjeqzuCSuZpnX7i4JCdNlnfF
N3plqlPK3NiIiLevc2nZYu4cvPnzbps1gCdXZKjaq6rqKoZzIDCGQSjvYN5eTzO4
LVoh8mrP+kPi5uz5WzHsGnpwQ3USsrzGSpkRcuZU2Vghd+seZM2Pjx8qNFVf6img
W+zh/sbOBNX6TsHE2nsyi5MdCVbTlOzyEDTLh7xESNoLuP8LuRyHrjnTN3I4tLp0
hA7RHlmXGggFvTsuO05u0w1is7jPzom0OxeypyMdfpAQY4osUPhW8juGn30VmKPX
23UhS9uQovZqeihBuuNjoaXZ4E0Qw9VjAcVKlYDYWgao8xVwnPCAMve1RdzeNlfB
kCwQLwd362e8G7iErxtZ9zKjrLj6tlLtjaBXK2tF0fMV+xMoQBR4qFsmeCOkdv8R
0p3e9x6mwgb8o6XpWI5GVkmj6h9PONVxX6N4OgOIaqi8zpwNIs2hZEH48imtBrAH
OD60523K77Bitu/L6Lb0Y+bDT/cC+QA9J8PS7cBamIh8vrXUOhWopohdyWVl3U4F
tUhkAsbcV2H1r4NU8qcVJdWefZLAqnRA4ArSp5UFWUlnxWj4OB7CSOZjg18VTMM/
d4zeOHNf2WCp2dabUGivPwPCEjxFQ+/8x5FR1N4sK7GZ9n7gDMsbhfl2RB3jTrdx
reWY4fDZB7PMpX3po8vI02D3nb7ET2ZBAQmPsx2kun/GjCrp3nywwBgtLgA9gNCu
1JzW+QqmwElpEaOoywdRvQeS1qNSU0ahce0ubR27+HDz3Q6l0IpDNPCmFcrJoWsg
+Bex/mY+Mbq4kBcKRPNm2++83pcBCHus8xIi/9nzxh5z6sVK+iqEBetCtXgnUJAu
Op+YpkXZPBr+oMgkUYSGVIs7DKnChFBwTn8fHpFBqqBuNjW83Yhv1dcKzAziMTmb
q8xIToG7yH07LnZ28C6YQUMt6SNxB1KZnpU99nDdyxiW9qllkeB77Q1VjyJsQttd
GxHN6/qBEQ2xBoa7FiHvqD+b/G3QsT2Xqw4RSh+RLmbJXPrjTfJR5Rw7tvyw6Ynm
z35ISrpaWpBlDQsG16ZV8LqIiDVWPo/PooQl2qk1ILJz+f/iGR3Y0q3bSNCIVqbA
v/nl2rTUn8d2Evayie6M70DwNBMcgVIKv3k5vmKc2BBxrI3FXUS0dHonKVx00gXS
a2D5dgCxHFBA+eCFecanSyUFNof2ltpBqY8EPDiqS/E9t2d/M7GaPXNfFC5MAeqd
JE1rHgvoI1v7ArlKnaFp9nb27Xa9qjCjgB6Gb9fdySPrjtRWvhZBVO8psIOU2FbJ
zbGYhEAelaSQsju6p1mL4fzfRldE4nllgEVIUhzwmDfDmWZpPVDOW029nWs/nqzy
o271v6mzA4l86CBF0Rwun+3r+RZj25KjtrFJsyEuiDLHa+loncA1SO/WI1dZQdWO
pIyw8nh1wkTGyyw1Yzi8w2KoRHWTsyQMQu+Viz4Y/r3MvdQYxwceuVVX5MjazzmX
JjKc/BOfktpAMiM6HET4cBN8x0ntKRrDkTv15UhB6wPnGiuCZYQE6o0zIXqL1lrX
zCFG38PDPXSPGDxUR0V/IJrsPdCftPDI90PZEr/qHpgrf3N5hccHzkz6wQQYGuk0
bv47TqpsCt+4rhj3vBNqbrsEVgrtVfUviTGujwDVnyF8Syg5XGDay5yib9ZX+ZFI
zjiPGENX4Q4UWGvkgcZLCOAdNB59efpuayeyboH8Ve8DTkAdHu5iyHvfXKyBOypD
dSG8mAA48zNcCXqljLvLI2ErJAPJC1UPwwvf7OUEphp5Vmw8B3wvdKuD9ePadnO/
hWb1NdpKaVf7IGdLaagabx5LUt7ch4NgrQWD5DLI46V4WR5A5Wg9wIknuAbi2oue
S3lN4kmJ8VbsPj4NNbuxZTl42i+cjc1TnJUdK+GH1LlDmCFPHlzAWnIhmuwcDWhf
erzUGzocha2y4mdzNxEfuzMT/hifvs71QH5eTA1Hmply9r80ISnJCIzHvPRamSkM
2i4ScVHM9A+WoQNFzv3YsbijN42kTt2voyHyZ0KSWH0h2mFYN5YyNO2kfShmYWkD
8w70BccVh933HflVXZoN5BBhQsT2vJmBNnAen4qBFzVoclrf1eGn3m3tIfyODT0X
RUHaTieVp64uPwhDTlIAMnOO4d/8t6/Pirs2HRf121mA9czjaz+uleMfn17oayRX
DDIWPiTcv0ElznaSLpuG/DXjc0g3YOMN1Q0GWpdXoxA1P9ZzW/uJCOd5TGK1b8Z9
LSO+U6heiwXLtgFJokq80xegk6Xc0pgTS5JbLVK6zZpIgAx0U2ydlbKN8ldROwq7
za1f+EFOxeI+I3rQjLRwxIUnB66IQzmlD6g5v0TC7rF702ALs4ztpI36PXFKpBmW
8eMJyVMAI6QXfZgZgFXcqq/LMvzNZs9Edzo0lVOvv+q4OMOfC1fC6c4ymxwV2eX+
EO04kAWI4gPa4t4WhNSjE8Wb8nIvhzpBsV2pu0ulGHgTeIdAGZ4Sli8yNYxVkwZf
vcWTzNfnku+zLPTYxClS1jvBw1qMfGuRlKcM7b5VRNK1ZkIqbYqxWcXj0gcZeCnt
K5PaUdVTijDN9rJrSKiIsyIIMiFGqD/m6L31Cz7UnMQO/qIZ8wKphNzbqb6Q0Da4
Af0j7fJs5bP3m+prY6RLEBsCH7PucZ6LJ7tUtXrS8qDeinTITHMTiyD16Cj8mptA
gPo9gzJWY5mD+DzQBAINVC1NZGVg9qPNG1BMTZNHJAub/epzFAe0Z2YGtpyQBa/Q
PivZsmMsCT1lmVJjwCGPf0oIl8xlL7ZVirCMl50Xwk8C7KlOcIFejrpAs5zNmh6i
qBHYeiQ21nhc96CJLysit9uMMzXilNS56KsRJB8S5Nb2XKNFfR/W4nwp5/tNaCd7
CZLxTBs66bAfcryUSYUDNu6Ql7m3vYepssfWP9nSxpwmcami2PPMsr0BCG6R9CS6
VinXViEH4mQbqNxkXi0XFOAltrcVGBl3QGLoETT71OBpLfKmBTDToJswMGOK+skt
v2944m+6BZ1Ltzi1QDl1owQqufLmgC98JiGBvRxUWAMzjy/xFZhi6U5NZ3U1ug7C
swyqsawFX+ObXt2N8ubyyeiLmGASCboaILS/ZS40WJRCkAZgGjoZAUIea4aWAlN/
Zw9EK2/V0rTbQ6PAZuba8p/eiWfTo9N+QaSsW8V8Sy1QEY5ArI/PQp6KOsqgVb5n
RovDkdtOVEESbj3nP2wxGyg1Qcv05wgsBvUuHW15P7c7uNhstY7ghRhPZVCcGQQF
mqjgMfN7s3LlHlwHXnAF/SQFb8UrH59LhVQZICBwVkqGWXcgjIfyG9jPWRKtSuAm
Zqvjdq0gWtA7Fo77NVHSezZw6SlQoJL+daWYQlkhJAiEGmmc/DF3GdfSkcUK4NZd
y18y/gUhDulp8Qzbl+3WOlwh0ni4Mkwbg0hxFOu/nSpCl+vDQ8yanhZc/JQ8J7wB
GakLWDvFeAQ5zNdRt8TtKvF4n26kY1gSJJpSa3AT3E4/nNy/RpXOkJu1VJHLAIiM
qpcqLJzTuwMUlBAEtMRSirhCjPEEhjOvYyex/mcBAlp5Apy2LYmhVMiaGza9BxyJ
kNns46VY0UmWeQY6WFclHGEKuGtE+XbI2gSkFHbATMq2D0ZBROXouP7Jg7wu2GU3
FE/7oaOrjX5oQb5UiezAq4DjCj1f3GL2RTj4woxHPQp8zXA7jFLRnSJxZknkpENL
F3uCHA5xyONkfYqQtw+p0P69RPHTlmKPSlpO+jdy10oHE7m56r5jnc2k5wp3IxTN
10M/iat8J03wzGo3tPnmOc7+fKMBByrYVN0lPyWhmv9B5fv1+6ItPaWKU5UkviOm
jVlqtQNB+Asw9554fPNZq/zTRGqtgh0s+1brBlWFZy4a0ZaMM6CXxzhwgQEanE13
SCB7LEFcy3RFoliKieYahS/x+rEgz/Wb6eUKUBralFHdn3nKNNL1Pem3SPV8aK4c
jhNf9/1/EZzfJfUeKaPzfFfCOVoTJks3lqC2JLrzYa7vVSa+sRfS5bC1Y2XZqlb1
z9e0tGUu/NuCj11E6laEYDd1VPtc2zjhpr9abTvIPdZjk2dKyelsElVqs3/74Gqi
sTk8kTqVTmqLYj4Jr0zGPdge+QMRJ0FUSSmIPsBEBEqDS8KOwqFoQgbyvFdRegSs
nAO370BoDAdKyZB7wdOcxGyh9cygtmcBBAkBIkOjalMeIcN2sA6G4fbMCG4ahvKT
2z73ZA5ef3BSzC0cd5/jMYa4i6AYPm6cQTLbCkQkBM7GOhWsDizfUvcph+XCWCM3
z/+Wr5MLDGJkaRWWsl2tHlxS2lNs+mDiNnuaQhtbL5jnYisMw0CcyoZjMMl7CAUk
QyfYwJ81x5va5ciXXJdRxmOJHVEsroksaNx4kyKHSgaEiIZLVzJab2WkLLykGB0k
7SEvyffenbzCtRmLqi0KWq6JqBT4bO4XWHVKeMuQ0DOrhSP0OPPwh/Ul/L/VfbMc
4IjvkL0GoOlqHsRoXeDy8/4XmwZUuF8wxLRmA+t2KoDSvznAWhzuJgIQ7IiOaRI0
EJ7DRAFmDNRO2IvjKxUgbiAq+eONWbrGZupu4iq6Dn5D2fEYKMFWOmdw2aRMJ2Vn
uGmVnr9i86bGcwjOi1OVDT6dpe1gWw9wlPwKrMIX3qz2uoxmFpXq4pACgUkf7wom
nJsU+bbDRIFW+SB7ms6GZRRBopVua2Ektz2qeGsELh5dbFLVNRICQuBf9Xwswno4
zINQryvFTkYnRPYezdiIqusOXqv8ZHwqeeybzTeMvAfsgprj54eooHpGMrkNsMvn
1zViJtdd9GOO9RbIHQ5FlGaf3d19FOmUaRPziAWSShVcCKja+hem6P5i7LDLT6aV
Nn+/PNbH8fFftljrW+Zn57PKavaMPIDgspSdzj5d1EdWwI1Exayae5ZDEtweWJ4L
7Hwi0f2DAsoRfr9+tByJt2LV2LcPnCPhwZKJ5xHlgXzKtbxTbBY+uNx60ztw1mwe
dT4CYB8MAOc98qmBIfeHQfvAuNjGW3OWdYxiiUBOux2RwS5Aw4g8DBZZ8KazIroM
bak6Ny7zM/2w0QFaJiZzcZdPfsiU9SbRPQg3lCUfxgQFgC6jW6OVHFx0IMDhc5lf
UM6KvAyV3dlOLzZW8/HZ4C8mwHbImWnPqMVyO3+5wH7fN4T9xTSDUGJ+YLNTg9Qn
dmkZm317o9XIMkS5KYfG3YgQXJSRW9JyXvKtoq9naLxXjIc+xhYWuJeU0gbEJBsg
hBSgXH6cfTgzr6DkSs/MtQ7pJmcF41oStP6/Bi4BP+GpPQddh2sfgVSTenVL307Y
Ui9p4Kow3W+1omrvGbRSoZXHuSquDIQoHLrzWIsXLPF5Bpi3DdcWz3R5oD6oBOj7
2fe0Gys4FeLcZ6fBjyXlXreAZSVaSVz0phLIYAWZAEb7Y1OqXFry6UzvzMcRVDKB
91zDFjXlq129SEcyHWC5IcoLcwdao1Y6er5yp9kbS87VTtkT9Bjg3IWhPXGF0rIo
0iuIqb5ce0ifDVdtkJC7k3H4yLFK1tIRuGtFtFTqgWGftdee3tKV0Or4NqVVs7DI
v/yJtrwSA9i/NY99TxqM+Cs++q5nbLYKDApZ9VFxgYkOhpoTTcrYfabQWzMN7OTq
JCuFfcLpmHe0X845aLRdyTxLeCr0/CFvuDu5oYLXAgik5lxh3IYIIaguQiwmaisC
5HfywjuBY5Yk51kCT/TqpswaO8J9A8D92JzcvtpaRjiQspWEOLfd6HmVLdEa5iUg
hDmdFB9B/K04fX2UtCs7oZOMoRLwzaaJG1GZGNj4NY9By5Lp5IPhFuDOAy2oM9hy
AaC9gv5OPCdZpm3Sh11UzLg1gyFXSA2YpiFiPJI4sU4VvBJiXtraC29+focZukXj
i+rqXLDXy5J2Mi8l1PYbB9uJq2Bq2VYzGwWa0AdFOrBR88SHvQ6Xc/LamCrCW6q8
1LT2sFLCySsKilyGKY0dc7VPnryfcGBMYpLf7MBTwQXcd74d1zDfHcN2eMw9bN5B
upZ5ToIkBQB+e5jJeEXUY0N5+BMh7tj4ptf0RMWH0U6K4iAFhFXGj0VPdi/N6uNo
E/oTNWD+iJESKDwRuAiR9JmUGDakRNAB/4KZ0isCfAdCeVYHgeF5Rc+wpaVmQS6M
zNML+kuJ0pQbB6dzhGcheFiDh/Qo8dIaZo979YJ5AuPJBVefA8noi0+7FE198/a3
uZRRxApwnWtKhxWzNIqdOcZsrX1wHBGADABwR9DyWeWe3gRSVQzJzJ0B/EmujwkZ
Qfh8DTks7r3PJzDarywnGyyl3llkkvbGgp2uzBwHxatdKM/67Lq83AcDIvCoAPcx
ROf/gZjGj0HmM9Fd/zXZ4zHYFJISGqWFIQ9qNFRQC+nAmd+BoABkqxdp8v9JG2/e
R+RQjR0VOl7mpDqqSMVsVleYsN48jTyHl74DtDxjrErQ7sSQvuFSpqLApw9ZiTaf
xTduKDYHN6aFhZ9eQ6/kTkkeHfZso6J67GuLKEyLyhsr/VRw8XVz1LLVXPH74zn9
5pfs0d2A3kwJd/s3b7th2uzolsAsgYFcSb4grIQd2/6vdKVBSCMqdBTYVeF0qFiP
yEVmQbAftskdMGUDncr7Ig6U7O7eg2OfpQqKl39Ev+RtcuXt7HNdM2/K9GnLRudX
5PkOL0bSOVVucjSg/cYSwYFpgYG3EcdYBSWMXNJsKCf1MId5vZihaCJ5m4LQpyBJ
o67ZPN4ZzsS8fGpsu1jRRjCRYbmt2SImma4e9tDGsznk876evsW1M/mIGWD0OBic
Q4zK2y+StR8pGMLU13WrSDzu1lU05y8i/pXSL4dqJLbhkqeccbsD7oCVdKpK0Mqf
XCv4bT9dHKRPlGgcDvn2ZbAYlanzjyrpvw5aKF+IaPy4botRDsnINDCmYkx20300
jeEuu61Fs73DXlQ9yROLsWxztwfgx9tLaRsvxc9FsQGIPeRDLJCD7+srY9lZpBNm
yJuaeKpZLIzNwZgYWHlRhcBSNer4Wj5CPi089NRzlSZ4Zl4CjbzPBV6AUsBKsN6G
wEcCBg5cLHPDoxwT/wtlAmc5wWPBOdVrC44lw7u9VRpBvxhdoU5RWk4kPdAHvcsG
QXqBBBYmr7CCe7Akv77MMNPq/VCVw2EKAsOZPMq3ygDipsE/7eF0upXcBgeVqx4T
BP7pSyHzs/Ui8mCj601BXIgoJjbaFh4Kn0XIG53IWGVMthVnRAH32owlrh30IPEv
aEY+PSDuiwExpHq7IPTjJrULczuemIEVbDiH6t1w9Ga6Zvtya4FhNHjZxQ4rvJdN
znLq3BBla64ynlUPhdv6rJGgoz+yteTzTSWKepIMfqx1Jj4h29/jiscyT8jAQ5Qn
l52eHPGeN/D0t/tks0AIY7wnV70xmiS4RjO9Mo/Bp6jTwIPTaCcByBYTfO741LWz
4VUY4RQtkUf9eY77GRZWidhNKi3GdPopS1gWqEdpCiyyaDL5MQneSVgCu/Tf8Juj
OkR1hZZi1sbY3ZfHzZxxldiBJp8jdRvIKRV63tI5izn/WPYHvZVtQjrzdrADctoF
Mv+Sr/0P76Dpqsq2ZjiAuVcQ9mfIabUIbfnL45DgS9B693W1V925UTlCmre3SXmg
19A9Y1fpuvEP7+d7YwemQCkPihmLy96nyfhX5Nrt69zu3QsCPnsSo69VUbReXJez
nUEk41PAgYgdcXtwQCSPGQyRwtz5VYlwM+rkvr3b/PCytGsCfIPYPPqH2/eBwtrp
QIO7YSDwAitvHvS3/bhzxVFWQSNK+/bdNV8z6YNWLF/8XIyseKoA43Zbsypc3J1S
yGgVcRx1gIkQmNZqzWViVkPC24jV91PSq5+3GT42Hmn4M5glNFsR1/4h4jhClYIp
D/ka2QMoeF2vOSN5CuPeJYQVTMBdnr3sJb6SZ8vbm16soYFqVYtlC5Qv9O/W93X1
Q8mzKU1odONS/wIa4uysJfTubyUoGtaDFxPA4T8qEtuVPZBLWFfHjpJ73/hbTtd0
qXyI+zM6oeBRn2w7k6y09b2UY8NHZXi9FP78YNI1kwzJjCQFNarORvW/Lqlh64Xt
fGbhkyHARrcuB3tZhTi4qNJw6Rj5VBxmw9LZudx0+PcSyDwc62XllFp9Erb7i5J5
V6wDe5twPwODnd3nJtYBE1DkTX/qrmsvjiyRqgef1Nv2S5JWADzNd7LmijCs250c
KlfaTXhUiKOLVK6JUWcKNziYth0Ry66FxSICj9DqlghMuvlbqGsfoilrOF4lqey/
Ogm+umiaj0zbd35Zrfj0kOdJ6AfRRLO5c9v+7Ex6+fBn0gDOfYL3Ac0I8+7mjXvd
NwsoTMVi48xAC0QMyoZ4spIQV25Drrzo0INw6VWwtB4rLuEjJ6vZ3Puvafqh3K3Z
FihqLY6DqSR4oJNWoPezKEaCPSnZuw+WiFnXRHHxIHfZ86LUmHvhV3JmufJFuMVv
E4XhsKC/JFZmRY3JLxhz9H+p+PnM0ETSz601rw77SgrsA7HogXzv7/qf570XPu0U
85KDHz+H/U3aU05dVPnLad6twJbJHoBjxGMFD3Bp1yfV21Ik7+9J+lxJ5PCjgh3I
sc/4VLqwny8fFRUtCrPo+2OgZJ97YKSxTXLZ9HS6hd9Ner8xjZcqLsDYkMEc9sKX
YzbHYzOyRG1Li/NhyypA6As2aivwdFiEVjqcPZQiGuG6sKeBgWSMOmaUMGfUP+lU
iHPTsho5wdiktAZkt0ZAWzXpyE9LaNw4WVgEK3Fh3x11XrcLP7xPQ6+gU5iTnoRN
ly6ugq/lDaWKsJItSe0Pfp0hLM82FIXDohC7BNiRDktKW3UIITpRF3hxDe3zyrTh
PU16U2uuhucobwuC76725jUZ7ss05otV6zPPpPHu3+Du0vo1B+6yeAp/sxnyE7iD
WHFzCwVxkvZefv3Fts7LFEerIB6XHSQyPlHjmKWk5VNS+dFim30G4dNBo0xYjzro
e/X5t3UR1NLhor/bC7/QnleuOk9Mj1RaydVbC5yn+6sT7rN3DpE4JFtukVdk3xwv
LgEzZUd4nbpzvZ2S6UU72T3tLsbiLzVifzqnAkj6CXosRPuMUWYWRHagzxxrR53M
2GF0I1OQW4XPK0bAMzXNlKgkZEbmP6JDZP3fgc3BwoTG8y1cZMhsjNwYiR1Yulnt
LTxtPDM1j6Da0nkGtelQPdky3TKB/IAPIBYPlvlrSjjd0RTiE4oYUOwWgsyw441Z
0f9SLuFZNU4e4fI3BTy+SlmxoRZOYD3XWizsHVt7ixDYBGk6lVo5oDjE3AGPRMlj
r1OQLluQM19EMiR8SRpYDaAN5Ymi1Di54JMlOuIl4s7NSm++40wVfwNPpyRjVK87
RX3iXr+N1yvSu5VBxnO1XjNGSSAMvKNuyx/18aSFSHOGiMyxQtz4ZRLtOUZgidCX
+EJy64FdBLrtDatDVWilibURfN3oyR6fRumDSsAl5UeYT+AEDRaTkGezBitRtOPW
3JzTuf1iHhhfSUcO42xWTDKdUfMpw8m6mRxubpYbSxgJtWbahaB9iscHgN/CBLN3
f3hEN8cdSenfX58kBMlBbnoq+PSjo1+fUF5g4N5Ip0zhzhHk2vKaAW+qheei7kaz
3t/tVroLAMJ8Yz//cutsSJoKtpIaeb6d61PHCILnoQ1ns0uQdJQHVpLsPg1/MvKA
0KEweS1ArCNlcIxlgWy9HZRMPWni28qWPH10+4prMt1XqSruyBuM74H8uuSh1iNz
uRtPpeW8c6kJ2lk3EHqAPFPDk8UDhp676kfX5tV3k6cZJZqX07BwyTMKp+0i0uzk
pc/sS/utbS5I/ezgmvbgsxaeo/Ge1AmsFW0klbrxJtNUBw5a4oC8peu8EU755R4x
L/MooH3MuMnF3Hr6Tp42YpFervp24ALTRChNbYF/E+PXQLcjfbM4uHZtA51dKZoA
FU3Za+YL8P1BACaepy5UQySWdLCGpiQtls2stE16+YGVGx8CZtqXMZY1euD5ZTvZ
8YyzYUTLdwsg8gSZH1y3ycAJzYB3tLw8Uvfn7X7zDy7fOJiFeNJ+lb3hgQNA9CYW
L8xFBp6fTyVqeDBcd1gKl4Hb/pmdK1CFBNu491XxvTBG6QQGhuCnARXPnVg1Wr5Y
I6L6kcARt6UHSA2cAO/dvEH7to+5vasjMUw4RULLzfgIXE+Zc0PN7LDHZReU22XF
PYntFQEEuKzkVFD3ii7i96VnEBZkw81l8IBjUEfWGmUglGDJi1sEf78UQcZl6+zD
Hi4X5S20vQbaJJsnNx8ZVOJ0lCaX/rwbNwp02gWnMYge5zeY/crk2r51ooolRqRR
GK4pkQoD4p+QntVfSsdZoyoGo3je0QLnq1JoxavYbpoD4vUxM9GMtB5+qhxubgs+
Sn/vuDv5BN5qYnMu7hhVFXTx341WyRXfByi3dxefDeywvcu9qYO2GeCgxHRO1o5t
Tg1MY2iZFS8irTx/+m2LZgCuMGZAmFd4gBO97YmqaP2psEISvGpBqJpakmSs/GGN
KKhZWtnf4E0WwjlYXjg2HKfLAksbAFzgd2PK2ymrwfRRw5W/mTjIy2311bTQk0Aw
RjZKtPL+tB7c/nv7hvGqN2ZKEn1iaNyZDwurTlsnUNUW0swkvaS+/MtU/lfLV48d
eL7aWmQN1uL8Dw8S2vJeuwuFWjYFJsliA0xoLRPELh5FVWE2uy5cIHp+egsuVy+q
rP4hk4mlcryY0pr5214ENFcumIBFBzlZHlh1RIoHL2fWQ9Fx5Y52lFxrnswkQndu
/0CeBEObkiGdfsmSNUKacZcjgpLi6n5yec+kCtz/UuZPpUsI9+shJu0e9xdtwqZ4
5AiFTx2jo9waJjiL2rjwDZu1sM0O1DIbAlHadyZstlziOpcZ8qwY50KZCHL92OPA
RtBLdA0wJNHS8MJC5MDrUPc8ewRigiLmdEdoPrAc4Dgu2IhstcUHkt8TqpMFyO9A
KjRch8/0E0+Vf/2VweQRNyckE8pi69J/UuRWCl/ytgy1LKYfhqm4GvgQDA66d4Yh
CPc+lfXYLh+ba+MhZhq29/XMjhuB9CJ5Az20IaTEzDtrr+UFYbTMTWHwZmIoCw5n
N5W1N5HhO2znQPG+3UqQq+wqYXkmOWKJe8B+56ZpUxB+Kb26ojK99u6dgq7cisSC
EdzO7By+pThqIdn76IWgWUW3SmHexVlU7CWEbO5v8YJEdmGk1EBWyJAPUaRRQ5kY
ctRIG5TB31oBE2IV3U8m5Kwtndql39BMqJweqVlVY3oPEEkk3rUYre68a9/S8y4l
A6D78UzIv0HDj5YoBkIoB1iElJJn4GOiKuv2h631lT139550tp0iJzF9hJT+v8Bu
2ihuH7a6wbQbsCKteh/suwDB9tzg0vFEtEIKPYypVE3qLExiXNVM6fHzt3W2HRGG
AfRA5CtEkS3XqCQSa+ZWKmzmTPt/X7j17iZ8ShHuSuglToxEEyxJewvUFNvTpan3
/aK0sgLc5bcTB8XD4k7yS/NaVolQq9cjxVH7Dh495Vy1lZKcZ5TrX3RdMfnh8Lbs
EjPpcv25OvEiH8Wku6Fwsor3CLVUzqBKBhrsTwpWABO4Icm0wEQ98T/JbJ8SYIsY
26l8rCFw6qSMf/p6LcrV3KYAZHnMsCM108jIhCWB/ywebeTInGiGTVl7diSlJEE3
ht9DSpTFA8SJRV21YhVNgurukhL5IiBi4Mv9qyhnnsDiGPiPWcTUziFtCvn8BDaw
F3ToXfJSqvwStBBdY9pwrr9PI2eQdFX4tTcljPQHClWkl4yRmHiDgzTrn6eW3HJB
VMsQHAXfVZdNKW0prM8ZhmXcifti6EHLxzXPWDJrgtgFwAJW757PQeiewXKRFSpY
l3P6F+bnMhBg0E3Yt+YqY6VBBlVd1XIoswYc8PYD2GY8XtuolAhDpakiGg2tV+ht
Sg0DGtvzqJbFm3NHTvQb+nzKJ03R1802Y4x10kHZLdJ+SpgXXwqGrHDBYcLWKOXm
UoD+Ohuz2LrHCTg5B9Ws6BOL9Yk8g/JJPP3tvWXi+EB3nubV+4wcnARsBhRpmO+n
2hE+nZZrSJtDvV5xPVbGVHRWT/9LtJdVgC2Lq8FtLGpa6E4/MQ0ZhmCeKD8h1tLu
O36QTph8+MOnMFdl/4CpFp81upOLP3T4ZbBPE49Vs9L72e6Ad0olhx4ornJMSUE5
Afx6VHJuDcL84CwA8JSsr1sA4G+OjcMflADXKcZEQNXk5W2317NB6C5rSke8GKuz
+EvuaMM+xAajy9cXmpux7M+L3f2OGRouyldCeL8qdqHwUWcogf2aMx7kjxR7uaZN
2aSnK3SGwY/nIai7U0fO9CpVM8Au+KQzrXhSc6PHHsJhpuPa6gwYKGttVGI2G4bO
anGqVp5fD1m7p7XxbyJU5YvQHJnD+7DAQl1oRtDsaxr82hRcsLc6Bc50kt4zADt7
HfmhQp4EZxA8jsffd6Yb7jXyPmBE4y9VsAHqd41n/DhJOTMQX7Wg8xiYLLUDU7Rl
3dVLFNDXmulwOBfcCWX9C4UPpAUFtG0hiWhJD4h77wj4ZrXrGoUegUFE/YwQrhS1
JNdBS6/AiRIdZ2QXuEXrVtuGB879W25qs+9KmYJxBKP/4tV5EKzMhsL7YohvqG5X
9ycoA4PvJrrv3YpaLBlBXNh88XxausdPLD3tOGibmJ3KmtxwG/7SACFRIb7lX66/
DeBC0KWBkjgZlfD5jroiU6Mw5KXNMRmhgRbZwzzfkoylQIjeCnjKwQVVTgXFq0ZL
l3RwWiNMrAEbH9f40mxUJS+p5oAhSNO/7cnvSOYkmc9wZ9MCxYdDfdwYm/95NlRH
dMIIUxHwyZcDq7Pljhny5eXLTdDnlHozgGAVThosLp07gkZgje3EjWLd83CIBlya
1wCtVR96OuSRajKuqX5QQB1vRapKcJvkUTHXdv+v/i/uuomH0Vj1jmiXYfn1IrsN
UCcJh3Pbenc9tx8KjV/FSPf5zUrP/cs/F8tXOIUeQZOgRbCrQI2fc4feNCNLiq7b
YX3LOCJUebQTT1qeuPERdlvttmuQEQbYjVXG0JBBqLh0Q2Q9fK/HaZ/bgQ40yqj1
rZZEQS85oRoWwfiLt9BXi1gJQw3VLB8/zQfNh1klqY+lxqrfZ8J0AGVtcsjUPMio
yNriruk/yVaSoeY1IooL39X2q7larYk15ncod6OT5NG3ZAFRN8Q+s7IAHblx6nNs
5sh6Y8cf8CHeE0XQ0l/kIzYg0v9iJ4WWWkpSUtzZ7JQg37n6V//eQeBdN6au60rq
jMPlMfFJOy8E7gA7fRvjrORtX5mDig55mb0Qu2HlDK+ss7kGSPE6RgCoeqhfOtyf
6eLja1YaMj4exUPcg4nLc6U36sVI2JLAeUGHNCyUOw6Ymvh2ZlG1m+bKlpcxm/3Z
Ypem+YobbGCU3H+IG76v2LhzyclUP3WyRWh6D8K7TjtPG/lKsUilmOec9NW5quhd
/IJH1shzc03aKVbowAqbpBW6VB0xvAPgQpNTHmRvrL44hTgJmN/z29Y1vjOA8m26
j2YyAJB8fUj2TgMLk9nRCeqdPBduxzuVVNnJ55FwJ6nsGZDK2wgUf40nKvkQrg35
ywx8eJ8AVQ4Ql8oi1Iz54NTQtuf01dHm6/lgbH9Uy1O6FUcJkW8uzOlAR8OCqDcj
ap45krDh5+kHk5jMHRP7c4MI2OvDSpkkNmJyiKVYHChGJjjjq88XQKWG1vsdCN45
HsXBqoQr7bdjxG4kqKq7DAtKyFq/36mQ/i72SKjiog/BHr7KNEV97htQ7Lsbs0XW
+BarEFSgaQJL8KiUk+ZRqiqVfXg3B1ZMAo5Qpb53V6ynz+eJUWzUrQUmjdzgojbI
EfySkulVUEyF+6q3vjidmHnQui5o/w8MBmx7+kt8YoubyYOFREfJ6Bzjs/Km04h+
GdmAWRdwZSSD6D9/qVdl3Uj2ttXzlVApCgEd2UKJDfVVIAghRzZLnyPwb6m4zNe2
+ye3+jQpDTYg0CMSZB9v6rNBYooSYoD5J8Qp6pPmeYh6BrkB5tEo/JmdXTbS6jIo
rtpTkCHIaBEXJJxBMyWJVLUWXwTVwOVMeK4li8mMw+Z655DW3qKy6Tq5ytwr1j2L
sZCV89rlTLZCT6lVvFOLtqZCWPcxqXLttLsm5YPOIPI92PDZhUcNwMBa0wsWp1+A
O6TH6C5VYV1F8KHsHAwInd1fHtnM5YF+07Fmb+M3Sz/NiYzqkhrmYpr7G0fylZfO
I8lQZS288obWOnuXi5/9oDvrVciK6gv0UhuF4pOfSkAoCMvkrnMw2UF7R4VSOYo1
RS6+hGaimugNvtBuyp3+7fb5lnrnBFi0OHRfBsCE//yXqFBdBnF6aCv8qf1ghVCz
GsJlTcNuxFDI0jjiiw9XTr6hW7nrLKnzKFJ/6YDf5+CG15XllgjL+dSuECRHKIE9
+aJgNXoOXnh2A3Y73G7slBC7KY6NaB+bcqZDmacSlgztzwxqMR60hbsPbDHGZzQm
SIM4tve6VA3pC/xuCXreAs7zygeo57Gt0wFo5iGaiODLJJzqH3gHSBifOJ+mZi0e
IQ6gbFAEA9m7muz7pgYPk2+/dagIBetI4M25oHKwRYAZ1TLheAoCSOTURa9gU46k
Sy0M9i67rFvKJHPe5rx61oCdnEbcjVXYhDWZxZggxqk/Kh/X81gUASoe3FdxTpbB
yEiNz4Z+SwVOc9KRbZS3IXob2VIK3sGwWi56dk+AXjDldCSPsBaFxVcVh9qRAVcN
PWjwDoswO1Jq+VT4FbRWOsuDhUDqJISjxGwSqxI4eGSxxKQH4JoRh1vb+Vd4Y7+Z
l3xy3AWa0PlTjGrSV+PCfvePEDQ/Katmw+HZsRzQz4SxM3hmQpk7BXG9cKPE8q7z
UKt89G6Bpi8GtGPwiN5Z9AQzc4r8FxzeXMAvhB1Z+ySESP9Kto/0r44L8gQWRkfj
p8iNR0oX9Bnxh5nlpt4+g7Po9qy2tDEe8rRJlNKYydd9rXheN9LXDkG1EX9dV/TL
F03DfIi/2QLAO1u3WJGida3ZxqYsA3EhrAwoUpyh81AhlQOKOj28Jqzya9W5fBnt
JjlB+T8/T+tLe/c5+8n8k3X+6Js3JBFkU5RG+d5BW+1e7demMLsORZAGA67cGxJA
h01z50zewS6O23E/fLw+yXKm6eljsLDg/s8wylXhbNusXtkErrwYVNgLjeQGk2QB
fi9dvW8DxMfZZ3I8r2+iygzZR7gAmtKVNfRcN98T/8YdCvyg2FipjUD2U4jgYQFr
vImawCcip5DEtWLxBySG7apvJIkiYdmMKBOV93ZcSzYhT1ghfdUyoy+G69zjd8QT
vUzLHGcq+b8j/w1/1sRoB/bbVLDf5Fwx/htejXIXfme6l6UnpBiHcriBJ/wrRfNR
13YdCGWn7TdEzf/Rs5gLsB50R4Qj0MiyKC/acg0iOumzgOnES3My4sGBwnXk9+n/
gc0F2wzg6m3HzVaGTLRdFPmFyZ7u/bcAGkF/bSSxvnNoCLYEYKwuP0pdvmme44z+
L8c84G5jAYNaFnfYto2S9oFq8WwxfgQdtmpS0EXynEGtNpMVaXb5uW/mr/3BnT/K
qUihdholFCbcdYgO1IUkBh+m83u2fwXvp2ItAYPAAssnCbh7ofTCHVbWcufUtZIh
E1m8fPKmdaGhNiklyaABrlOhrNbD1PQLsC4MNnw0TCOQ/1F/CRkdez9RYZ3Iq3Ko
/6W7yKnZcVMn+1oaP7si8+m1S57A08pR35y+e0rwWMmtw+tPTWbs+FvWKmo56UjL
WJHToQ6P7Clf53P/uV01wM3M5bH2xAsHWcWWkweD1Y/Vdxw+fl377mTSFczRODyV
UbfnK1a8ryjGcMT9HTfigH0tl86PDOaKgibqBNTAMaK5SFuuISpnqt/+wzDt6nSQ
f3kMsIbXPO3H/yOqbZNS0PlkfnyPKqe25jrBR4fYJo2wrCLO8fuNXJIUh5wYMcpX
v/7A1FZdUx37iYrVX33WSEXTyhjD8K/4N2/F4EFzJT/4VqBHwHGwcTvd9IFk2zbR
26ilXC+iU9+zk09HSdH+80f9XGinthERTYqFrgqrOph3YLFPWUTUkJL1O7bcVCr9
ttHV3VWh2Ygitl9f5z33ccX4BWaFDj6eCU5yAFR3uNpoFkPDdBiHcTjKyUSPenEB
MNFkuM6frLAWv0AqAG5tyX9wOZ9FPDGQIYpeaAp4IuDmoWOPTrkt1aNKJA4ufOKv
Jm78ceVtC8MwVVo8KKJECScfq64ogSMOkQZykWxsGbc2i4ntUtRnRKy00WC/NJJX
S/B9tILcjzv4uNK1MxrapwanA3iVfAQdq13Zo4pUVcUDYt09LRMGiWfXKVuUakjd
P2QcQMnm86PZE1Qwlos7DC/PyK5quRxAVOx44cMclnEZdF4pHfasQcz3+sY88qh1
WKvKQuO0Elxb/5JZaWYFCihxfpmlgBxo1O0liWkUyl6BbxviMbJ6GB8V6bNQt7HB
6068MjLI7lh4DuZ1lEJL2hetOxvRF0x7tIDOxMqR28UiUYyk1HqxfsvTZYvKKmeh
RFUQlaZzW2+ejOQy7kjUpKFiuC61vEnh2aD2egbmZFbzB9xY402iQ20aL242AZdZ
OgAk5LOb/gOPWJFFcQchwwv/D/9GGyviMFsVdoSO2gUuHw3K41MknzZDNbC4RrC0
ksbj7Ldthb0pkOSQu2I+U1Ec98KEdva1WJr0odXKXbwAQ1ApHCNm0AzcElQ1fRZ0
hMpz9wyjkd95z9E45bVh7Sl0eTFeb1ytco+FdYk7nIG7mZkZWvhly/16bY5Ndd5s
PfLEZPLNQHGV69LGhT8y/9oyYhEH1oHHD7TELLxP+dlzu+x/hHd4Qxb98JdVcpKq
2oClXdJPL1E+TpIc34s7GpN7xuAqXwdVcuRRaihVK5wqMk1m2twsNPHkq4WzZmZB
zb2/DTgetoaQHUhuC+0HWv03J9l+1WvWUh3oWVv5YE8OM3v2ztmYfh52xyrRrvyA
H0eNrVD9WolhFNR9MJv1Rw+oa0xQuhGlvgu3dRZwQtnqxX3NoH0jFBeN+bz54CBN
TVSzL1twNKDvSODAWekJ6x9c8R69CvWu655HOTMrl2Ys075N9ahmY1UqLPCBcCoq
LiyU1Vsdnpa2B+eTHci9XSKf7HQZaiO48csmVm94heUTSJEit8a32c0U9g/WKKFk
37iSpkEVDPGNZ21ZMu8+SWbfu6GsF4z50R1csb3jFHU+Rxq9vQEHvZ5A290ypIaP
cRoMXm5KwYkReT4kxi8M6eJZPgTwhvUE4ZlISJ3kSgmAcnKM79nu8aThti5jkyyF
vjhLu3bqFktfQvaOGxmoqTtmUWBkTFfwMK2uVi4RmrXwRlirvjCAsToz+mLe3QV9
hpBYFjhNLmiT6wsVAdtH4aTb2zrpafVwFVGt1AmDUDcV41rgUmvfFeV2CErR7gMX
4YMpE8WA1tpPEeS8p9KjE+d+cRX0plZSugzwpXy5VT1zMFXf2SRDgz+Lz2GIMWrB
otsT5D1CQLBkmkzhHjEjZBnAmpaOXx3F11u0wuuZD/gyXVbxPo7c+oyVUkZSImoa
SnoJAeX4aBgv2ItYPJpA27zAvHuOrbUt93EbtuhhqTJsQWOkftn2Zu3+NnRQsuTa
D/uSDMP0iofU00KwSDm0OU3ZhbJuNNRR4kpZ4vn8F4lg8Q2VhveraKA2kk8fVCEH
i/PKgXCllDKPOtmnkYV9bHYQTBkJ0a1K0yHLuPf5K8XQPAI0pJKjzOhOGilwd6OM
dRW6xHidvP53mrksQd1bpkj1E9U+DuTOvJtbFVasd0SKNSBRufiRkEhWVg70TJSE
GAUO1xQf9F4fvxCRtFx1gKCn1J9gfDqoHc1nkGMLI/0kRhw/Ulas/PvUrTzTtsob
sdEznQsUMVlL7wO4IF7eBCUq3zce0RfiF2cBbo43het8K0nJbnvFqQabtE0ulUIQ
cZDuvu3pNZMDVdvsRZH3j2QqgQ9lvWaJ+Xh+vq+r/R+Q85Wf9gaRB0ahk1T2m+Sw
J/zSW2pvqZoHkuQz6iO0Hukt2CHu7j6LcyRM3yM+dASqNnbPqQLAFpc6NKYlT+60
rhLZCKO9kLH1Fg8D970e/FPfaM+Z+LiezOBpvRHerPDM4Lhve8ZPabMiRBn33JuA
S60cd+bD8imjU/htmszKwnfF9Spzgye2hUb+fWixOtuiTQGMoFq3DBV2Ujvi4LvC
d43rPCTh03T/B72l921/Apw3koaLXUa0mvBN6bKBsIdCFGAvhWrgNcmQIpEBqAT8
QBfTToi91sUf+Gq73ms3Azx5WlViPrVvaHiekBRsr+ZiaUL/V0dPh2mfovDa2Q6z
lBE+84Ar+CYI7Fx5i0pjpoq/TF3RB1UVuv4ljiT5x4KQOaPbVBki7/UTJDr+R1qz
97pDRbKAU3a5Lrkg7ybNJdYOeUr3HIOKmtO7AFnEWeSutZdDC2Ti2QOFFo4mZV/W
cczKH5Nxh1PZ9YS+mQDE2OnA3nUNCx4ujb16vu/2O05UWZnWbSjc+bgZWTajD/gq
VF8vToE4XIITPfGSbb7xSU9AYW1rKnbk76SUI0x2z6F9DVxfKqlxl69vTL/rjMLO
HiO5zPji1UbTfYAurrTPsVYwdBBBqLquPOA9x3W3H5LfacMd+AFfQYiUsaanjmtU
7rv/6XQ0A9EpQcIy7jAQd7JNMKt/OQjCI+QdwtAB9Qz7GbktKmZmcjLzN3pE6wQt
kyEws/c2APfeoZu6IWvsdZ9k4zcSKXbW5Tj0BsWefsFgKwCH12oMgbp1yr+5LdXq
GIJI2mEpMOgMYWQ0GZZYvaQ4Yupf55Y4hLPHDE6HqT/esAD82bjdmsK9lVcCoHas
evsjd8VNjrv9uOpOZPTVfQnzgZsRoL81K5+BrEdzkPbftowGjtuvDFd6by4GRrtE
x8T/D1gLlcHFB6WHf/dNDPfTugld7aCi0dGXvI+65ouqmVgOkWL1BvEGmQbdOvge
KgN5tXZdVsC+pyX0XF/R06cnmUs3Rs2eDPD/DQ2w2LBSfDvhyo7m+p+AyQc1XF/q
+yzg0EoT95X67KCy2DX17mVun4ixkqn/hnOqgsNgOAq/puXVabvz61LGSdCI0ap7
JwZQrf5UipzEZ6Pai+BYjZgNUcVB9vQ7QjZy1MxSxcMgUz3fzzigoL5dIBekKNwG
qXCTKf+o/kx1pD+EAXvb/aTwr/z8pBjuJ9gTLKd7aIO3wRW+Ro7N6+XGa5bdrvCQ
w3LllLYXD/A1i8u3zx2WICWP1lIkkqifSxjjYv74t2a322mN42AkdKQRVL/87w+w
WsgQ/tBDwi19RO33WbOxC8WzVpbKBdxndzf+YOkpZxZdtiA0r2mVBu4VmzX8JMKE
xjDbBGRZQMTt4OW/D2pHrKSJTd3aom1SCBCyvJqfDPicD+9o2u+tcovoczLa6Ac6
b5al4u/rqrXLnWInDgQ4pdy9t2I23nCJcezdYDySaHgOyC0cthmgzbi6HAoFpaDq
u7d/zfLvYkref/pZhZM4jjZjKfDmoLRn9QJuK3vsoHnYSfz6HAfruNwloifbLafZ
sD4Q3CLoUH+EFzPPWU9HsncStdizjlHss0o/UzTzM/dFQC3YTYETLYvw3Eg9h5cQ
ZbEh+cok5F0Hv/66zrB7IDl8Hogn7sKi9Bh6fTxYQRIJQtDJOC19xn6TzwBWWEzV
9TYBJZIJBUpmF7ht64slQNtq2hjeQtLuGKHlM59fWXJOZYO75rWPfSc3NSXjuqU8
7DWQqjrzlQffmrMZQuRJfHXalRTQTEUYjgHHurVzPfLXEuyZu84L2J2uVIk1+C5k
ECXPTpMutCLh6Fj9OIUhFzPfujzb9uspDrJz3E5jSpnrnoGu641+89LcDLwPbIxP
b9/8ULmZzmICRF2+QnxN+09uwyMQqpG65RtQTAqjdpx+VOmc8xRq6RcxbBNNBAzZ
Kex+3oJDscTNwLIE6L8vbwmNEhdc/oSAIL43fn5QHTGd1Yp6C3lpeZvYN//8iXqc
pBlRtdkD6JUv0BUoarFxhzcpPpyq9IhH9gNEObt5awhL40+lyI+rjn+bSxk9SDyU
f9PbJzI+Fm5AxOU6fHqF6b47veg8AhiGp5tQ48yuk16N5SgZ7IqGZ8f+Njd5UfmP
VDS7s7Pnlk8h3ONjMsu+ZlFGdtDvpngyBTzBYJLgZgDpR6+dotxyUlyuoPtSsp16
4oldPDqgOpMjVgCMzQ5KJ7qfaxwXOjHQxOwXDKal/78+lJMrF5GBM9NvALgdVo67
EMDaoLgAljlkGz/Ibp/Li+vjDTuqLUfJP0SBRWjcmojKwHYrpm2LMgKzcl+jQyLW
UfSjol+eMCmP8cY0WpJSQNii8TCHP9ZXWE8SQ394qCJkABUQzAlxQcWsKpScOj0/
FvlHzuxtVuDsEio3HJFtdXALnmdYgfVWe+K4DwasuzuPVBrQBM4m+KY+ef5iw2WS
REtR4f+LgLcSAVDvwkRStmD9ZWJFn4/EAVpPrF32OeAuRZsrHktw3fYTzM3K57LU
1OVa1A8+jXpAz5r6SBiQiLJQMRpb87DlCF4HBpFkr3S7s6URDVPcGX7dK1rYMP5P
MOcnb2w4X/m7TjLn1bSyDTKBTpVCga23HeJTtT6cYhFtOKBEOGL8qbF5ViA/wVcU
NySG/ZDHzMvih+1sqnvJOy1GnIdRzL1LNt/XYed+eLOFlLZSn5bAZLIPmqBlfRXK
TSiBalpO0SmhWAn7VNNoViwbUQ5DzrbwBfB7dQPfuOgAi8KoXvnRak8IJLWg42Ep
d2oT4xPQnJVR37KQok1yu5LwKkZeTmKBYgPNOJ5uZCvci/r/UOekMHhPUI3p2Fvb
h7UhDnN+5QQWTAmmS09FGULunVERgv7htnoQIxzv60bwXouFIHjhDkFZ5NXyUoui
EIaz6mOi4HBFipXnB3v3G3ePsQAFtlWyoaPKgQvisNf5NEs/B/ibCGEQRDjnRK2f
lQgFhz4HGzYZ7TjEpih9CgcZSWBXAFNINMebWDnR2NTY2J/yUNIAPTTCod1qKcMG
Iwbv/rn29MYSdQSY+2X4rYibVvnrweyNIhAPFDyS6u5bJ2SB4YX1JMMo5JtTnGyE
3kV8yxSEEKywLGw0aYu/maWscUPyh61dF471ON12+aOpkj8Z1nohYNx9EELubsqz
jMkgsI7d9vatslwdSSJmaDkCWwloEnTBwEfET/M63M+BqHDYpPYIKpiTRxSgvNgs
fMANaMmyIXpIuDjmOnoKJVkh5ioTsqhH6mw880ylnYvkO7wL+sZYhCdZw+COdp+E
EIozYAyaEsxNm4tLLj7Snz+zDW/Hvn0rwVZGz4Se3Nsw7UG0vgyvEjEiHjw643eN
BceiX84t5Co6UmZ3e7qzBTovbtY4OVBE4H7iFAAmEMcYMWdlrLCnqHszIQ5BH88R
41UAK2r+e5ynG2apqPFqACEDo+OHIsDkLpROV6W8vvxmPI0NV51d32T4Fp8rt6vu
tTi5BJlczAMrzyUq6G2dOcH2tDKpx1BbPRiFsVgIYiJQB0zI0Ki8V5+08233bgLl
fXd2sZOBNptg50atildQi8kP7tGC7nofsTjPQ4hcWjLGW60PjVCqSDWQXrmtOvIz
/PuGvl7n3t7iqLL0gnt/VPUwgfKJWRO6JGhTzvm8pTIaP1JjNJvOJzAlH/933tr4
r7/6piqWhVgOmJwxDRTd4fHtbEkyB6ygw1vJ6XxBt0G9CIMjlxt9s5UgJ3O0mtsZ
ZlnvcNKPYS+pXV4iqrX/ncdxgOWNYbO4vnaNv1LrQI4qCz7L4o9wSiEdWU/moOUT
TMrfwEfWNOyQJ/zLc6u/zvZ8DMmMPzqSsgk/73a2dp1mEExgOb0t5Lu7V6GLffsu
yxnt5Kd/+778DgCYeeY+QnMDLab9LXX4qam8rnMvnZTy3a3ZhbO7U6CZyj+9dT/Q
6azfsO22XFi1YrE/oIppwi75DeJBoQQe4lfglXZ21+SirctalGx90zdWxPZM3RBq
rd/m0GTe1Ph3KHajhlGClWANc6JUlA+ssvvJ1CO7Hvc3GNrJidkpDadZfy2bNmWg
hLDuxnYVqkdzJVYrpGYc3MAz0ubQRx69nYjxx3WVP4/ZP9SzfqivWXKYKmgBFlHf
Ehd+Rt7fJ8oiTJRgt/sy+6eG4fxRs7A3H4AEZIkcMBJ7vOCFPCmk6OIKtNRpIOVI
GDjyC7rr6w2stKaD/h4KyEU50jo+rRW72BGdd85Yo5F8eySCWII96UvAuG9ED8Xt
qOkhGvAv0SII0R4qswDjpN8TebJxC/33e+1eNb/knX31V/uu4HZARaOLSBRa+Xfh
yfuTkPylbGis0RHTYZBoFifW3QAtH+OYySi1hyLJl66JStXOH1p++1LsCFciiYFP
ktsKnMASH8pamGe28Qjb11wWIL6Ie3XT6vNzEcvTSk/MS+t3LBDPvVdQU+1TJseb
/aVI4d20Mj4anfjyXQvsUTd1fEldZUBSLhDoUP7SgqU9BgdVuLpF/SE5YjtgSTbc
lCBq5eccCSB9EXF5zuXzn1ZM+YTtV4lDrqB/EpIwk1pYCqcZJhN31Cbyqc92GtZU
UKkLeL1XC5Rj+zrfdRkwK+A2A4xDO+G3ysuzcIWtVVvKacsWGgtI+EttjXK4cdsS
YXKLfXYi8NB4iB2pWf8WMrC5hq3ym5bFNRkM23tJIis03FD3UbfDs/VRB6pIMw0C
VrLVkAEiJ204uxNg2SU1A9kyfPsu74rngxkmD9IEecpmg1VdOFwD94R9lbjFd3CG
Cu6EXyWdUztdq+1aue6bn8IXKEtLAWoI4kwRnHT1o1EHank6VPH4u/FD+Lqywmdd
3rm1M3g3PrzLJ8gpO9W5TuXY3tLlqmRkp77Knwp8RSR7X4uCYi0WZnXGgzSqE9/R
z9kavpcG2aD3WwUWpkd9zoCG7AZOKomG1KwuAPZMldIAEs04Ge4YPmE99U5vg6v3
ylvAlrVfToGhqxGe1T1ty3MMfceTZ2sqhPnhEjVCMsGtTTY4D7AjXq4aRfAcibpE
Fx8fdOvZQz4KidfGiD/0yoCmv55qgtamDGAS8DvtwNqaQnSwKTk4Iczkpdbl+9G5
hRWnBmbz3/EVsTDg915qoisHMe+yE3ogGd6mCxtWjTVhFW3mk1o9Le4FuLNxasVs
lCdAYWAq6bYwy8D5Ax+mqH22tRloZGwcCNyX1qlTJ5nVspiyko8I5C1GKSoIufu4
myI4TtWQTe6tVgyzM1cpzpSyHZ8aWKVseAgBOoT0Gy+R/3mBlN7eO3gEYpqELDwa
rk2AGBvlNgBzhLtZO+iUswnRqmTIsFpNG8FAJ3YbZxUvxv+UMHklS0AT61dsiuYY
1ejcE12M1r92pZS79pdPxb2htVR+fXxs8m5emgDZiLqTWmoN/dktTOEovgNN62Fo
OIUtln3WuBqk9nCF06ya7Wloi+B4DeD4TKiJsnTVqK3s49gF3YQKaG6A1JWbBn5N
oCrXt7Yh5uv3EOyItJwRMqT+dQGeUazOcHmshXdxDkaeGML8UTObTLxkW6xLPB3y
73Y7neNLLWan9Pa3nilzhMYJ0MUibDU6B35tLrQaz9zxamd1BCgaUUPVWxkvBMZE
66aumm74FS9bYsn1TNcIcNx1bhfkzIR8z3Vp4fUOn2dX8Yx1TjGsfwzt1p+fXCmd
rv0KUNF63bf6w/duGaigIKJC72o111+a0L77+qtWQQbbGBH3OGTrKq7iOvaD1cQ6
GkVA25H4zCXNx5phD0xEqBjPuUOqgfMalt0UhlweMDfSNtixQw4MM9T1R6eCzPAr
0ECfz50RT8TlinelP/QECidzQk08Qc7SjWMPU2nhlQOI0xn01u42JeM06+x3PE73
WoXCF+zSYdC7eYDve1ACbhp496iiRdjgEZkBXrMchy1inmwRIiCG2eGz316Ak2ag
qn4k9GWiLZQQ0AV/q+N6YEwsIEXqBz3ZSKiPJqRmdymaUMpAwSEVUmYOCoGixDj5
FUMwGARz0l9LEK3aBT4uNYVRtCJhmDyRI/QDKI/VHj4QOJC5TF8eqG592x56IYCj
FY9V+aIOlYnmNGxGH5kqGAPdkpGovvy5AlKJ+90gnedvKEC+3eAliYZwFwlZgef0
OqqR8HgUc0FG49NgM7jxA7K+V+6ZSgzthRLR4pL7Z2pF1x4GXCLK9SyDMvnLo1vb
w/FSiyOSHN3LtIs4ai78V6T/P3Qv/7oepcKbkplOU9sMKBv5useXt0Zzh+NUj6QJ
jRkpcXCh2PIUGwW8ntVy6GrejNPKNmgQTYIjmjMydg2IObhKwFe3RVngqNN0b3uV
PGgz/wJUYVMQn1erh5T6bvRW4NWPYiTUS57Mp5pV/q3+XYOeO3xGBt+nHOX0Q7l6
hNo0IZ/SlxZZa5my9vHNt24PoE5I48pPe3UfHYX6/f5Eo/T1DGyMzNOuOs1V1psf
7mXYgQr5ucQoCn7KV2yG+c+abFHPcwEsi+hsw9Ga2BAIoQ8Dxz4sEh2nh+AAB4pE
b50UDswRpCOQRabFSG0ONlkD70sL7G6iRdD85RaaMQfdYt4kwqITEW7UsCT2RPjj
m111TJ3zsjrl4qo+GeBhaZJ+GYi6gSWSDlHZLPyZvY4pYzsNGXYCNvK2vOqHv8mT
Vb2QRX212Cf6Tru+toUgqhBHU8sDOtFoWi0X+9bcrZe4nJCyK7uMvp/EmONNF7xO
UqQpJFbIj4jjZdkVPS/6qgdHzYNXr1cArX88Z2M2U/WO//aAkk1DL/U0jfNewU+u
lh7GBDHA+6ZFKdaWYfpWRMy1fdKS0z0igYd+BJxUtm7PYQpCg6syrnJAbbjU6x2g
8Ofp5nwHTKeOKkIl3glJpitQzLB9ZrFU+0wIS217UBQ9tQDDOaA4+azOsNsi7p/g
AVkcdIxmOXrdZUPxWEv+E6MYHNceiRwAKbA5zxvSO3cTqMckVyFMFg//trbizSx0
wKWzxuunEKydcHX/CLV5uf52gdDINl5GxNxWZbeqHIGPiyb67AsZzlEbgRuCzVgn
ebm1/QRW/anK2TRYe4bJvx419xUxtGHPJdyeELzcn3ByGVCsDYl/Bq7o3/QvhB1S
rlSUIqGLF5o4/Bo2SiZl0AuQgOh/FpEXLwyGGf01xnoKS+3jj3pYLe/DB1b6sdhE
V1oC6LIjCQqLrGYG/UjjJXpUdGoBMQDYYAvDxVQEbG5FBqVuk/tzI8bD2qZrIKg0
ZrV2sR1AL7Mx9TfG7ikWXJfafnNRph9t89Z1ZqSHfmuJqIRY6wacYpR39nrhA6Fx
vVysDP1td0zPst7dOZTo3B9FF4jEKmiMFsJTJiQQw+vaqDAY+xzbHownHA1I7hwX
Ar9apzB5eyQDsxr8AGWjyBtNSoGK/tGVe3h30dSWh+bZfQcrFKHdYac7qzVIdGns
7HunqP0U0xG8uvGYc5fyRfgPJkuRBb5sy4tNR3N7wi9PhKrOuBUlS9sqfJ/q6EvT
bOQ97bk7GHekTEeHjnRoqKqJGzXwDl8XPh7fWwAzP5iAVANBn2crYVIrRmT+cwCO
7R/is2xgxQMn/tSktRk4YJlGNNWuL0RxIXm/r2wCJz6AmWBXM2CI0pSkZVUlBOka
4wRN5iiWpDlklr2zoy362b3TbYJJJLGO6Yb2qwXixSpW38XRanNyMS6glAkZVcbT
9Zp6nJYXiyn9PGUFbp8s9MkwlRmfnCZZ60Dw8pbxZJihqPRc1rsPOOVyhnizl9Hd
jgRl44qwvwEhcHVRfDc+etDTWe5IL3r39gHvJEiDRIN9BqSoq47rUjNxumEOq14g
49uePCx4X9UTFV0TVy1RKxmHc/Y+a0kXrFtR2VIMXY8TNnwf9Ypq1ZIz9A2fQgVH
7ydMQrtSqfSd4P1imA6JCy7tXQMfYjr/AMUM44fqcnqx2CNoR3Wa2naa3PylqThK
S7MuOUhWNf37xnhw0NY+sESuvjMYFvWB8BZnahOTNInOjTMdRFE7XOSu4SmfLlgj
xALiF69/ljhePBwx8WRShGbVrbEkLFRCCOs2sk66FwV1m1Q4YV1QPI0HyC8u2G7u
iH1pZ7XFPsi76wjWl7HolARQyPKHHKSaFaB2vOqm/mIm9D2PSS33U9F7fs0RlU0H
2JxYKeBG82ylX+z+rIPSQh9uFC/6gwfy2Ek3XHE9TcGFNsORSzE3/+UHB3Y0Y0No
WqYK5QtOl3oOhVL3sIctG00AeoOu+fVgMwXzoQkcaSul5wqauDbchGo3QrXt2vD4
UbX+C4glYB58nChPUojb222TQDr4sUOKbGgPAcc4T2OCti7TsCXBb00wY4/c9eLA
cVjX7SwtdyznLQDD/c9d3UOySfrqk3EiIJMy4dJfLUws2QZWmNuKGBjbm49I5KSE
1f7x1m6o9DHBwLWBl5mYhu0TCMxRJCYQK7x96B8EPasWjdNOcNBhC9yy1HpRwSxD
tbD8QGcFKEdrWCrOcTuxBiTMk/+NiZDONOMrBJbygrkPhGHLdZkVdvdwN/uIWFtg
yS4S0fmVGAtlcnIHCRV9cwVFx8tETRN+eeE3ctgNtj0ZlfGVVd8yPdZZblniGxY6
9LwPw5q01HqyTJ9q7ViU98fbRMyW4AWe67ZE3lWp2cfC9deVJhgSH8ao91NoLtqf
RiLqnb0nBD65r3S50nkQYPWX5ebNSfTQ6Gn4yTxSyXpx65NyF400VCHW9GWp3JPQ
+NlWsMmLMug3pA0UdaYovwtrBwzT8qXp+mBg9A2RD50i8isskDFyk+sVuwSh15WO
CpodkZARpX68A78RqrasfGhMoSTd3NKxZhd2BGUi0ns8Ae728dYuGsCCIMzmN/E2
u487pb04Jg5aX4poy7iAZvrEk0Hfk8ioqFN8XlbjKNTifUi2T6HC4FtUBfRnI8f/
Ma6mNg3U9U15FOWzfQOqtWu2WQhStRHEWCK0YbEg0JlxwO/IvTroq7dpbWFmAMbp
Lw3wDGjIKvVqcweRUQlZsDoV8a4YrPtBDk3gHYC8rq+gjoK/SQSsoBeTqpFAEcsA
Y+D/G5JsmOZ51F5dSxjOPxWWhVz6K4s8/3rj3rTNkIUTorvn0QrUHfV+rbGEXQVu
V6i8Qe1IgL1khgOTyf3uu0288pgFlDQYZd1C6aknlLl6ph1rhwGUXqBJ5hvU9aGP
YgTUdJ65LaOAa2C/mCUGQ1Cco0ROK2TwKQJGJDE4fc5LybppYFqB0xd9oegkadE3
B6Wm3CwwPaxx17lPWairTSk+k7hf4MwrY7r+lICzdZF7L4KMC0mkd/99f1QJOqPn
0Uy1OFhqAXXxfPnbLrDBv4k1wm372PgZi7BP0fZZ3CQr1AFsAp3ZLcFkAPVV3o/y
LwOYJOoQoLqAiyyHDGdUzzshbMtfHhRWnsEMPVwf3pyJtTQqD5F29RPbKILsJuIC
rruniuC3tQKRZdamkNmA4+aHxoQQJeQVoYxq5A+i5zDr/bYdnmf2MoxFn8vPOiHi
ZvGMGpmIY0scLimz9pz1HMfCONaYNcMEUUDpHuvz89FeudRJBezKEdYKs0umLLRw
SEPnqkYay9xTRChjJZiBEy98TKyvB+w6Q+R42DKc5ZjjTcharUapruUAm+Idt/j9
LLG1ItGnpYRvduvvYmnp3qKFHuIUcBJpU0pKpGeQkbzJZE1T6d/f5/QSixf/P0tz
gUBYbI5ZHkLGOUYD2EW3k2XL4jdeW0yLaOissh7Qe8gxXPm5RY84cSfdkp7abL6w
sgBI3/z1XRQKHyLMxl727qNx918OB9DfZ/ZhUaPRikZ/FzXEILiG4LAK+KLOnpxF
yB7/m7mZig2hT/BimscdZ+WBvejJoMjBlg/cAMkx+hVbRZNkORLyGfI08pN/kfJg
JSK2V6SoG4yIqtgXQ9g1PPbgTuEYFQn1k3sj799e46aXftzYL9kFTlBCXrydBy0w
txN5hHj9KthiBPZUOp0Gc9mgUGcRwxlyddnrL7fG4kf/8UIAxHPfwKrY/+alD8xx
R2rMRSB2mtIQcy16knoppvoc0mJJ5oSVBJHpwFDfhDtM6TA396A+wabgThyfi+of
QXIIVn8L1+3eSm1sVNI2f6b5xIgP/VDpAimAKwThSZYOjcMwGqOKsF7FLnP1B1hF
doE/K5FBbTJaOLxrKwIa4nWFxiXp3/i4QQyLdwOnN1LdR6DBJiRz5LMdk+wnJR/B
wIrlbtNaaf+bpY0lD5l1g/5/PJk/Kk65EV8Fx3jxfU2BOoRh2UuFd5qYmCdzQAoE
JgXtowzzoa13+QhRQtq2/nalvmE96nyXvzaETX6Cyxq5KiL1JdsNg/+BfWEEYtJB
BbnyQXoHlpDsOZJH2RVXdyAxt6KZ9Bi+/T7NvQdcnP7X9zRTjscT0bqIBxetXKg7
khThTHtQFxNhQHSxQINx2xWIjFtO6Eiv+OpOYolSb9VT1tCIDtCxmb0WwSySmTUp
GCuMKb3VARcOCWl+tZxKDRsASvjuJD73ih6J5tq3c9MG4DBgoN9QL8XcdUFW17my
Cyy6LnzXfRwl/Q5kXeSlA09u4DVdgSvlfpzholQXm3JP9eZNUMBVuaKxMtJdgUoT
EjIwVqavnDnhiHer0+sSwBPMcS5Qx34GDVNDiyneAfVnzGTEH+jEwjU5NdY4D5Ko
1XwdGNv0HLp1iE/Dwb/sTcwhzEbbufHXbwQg8uKZh10NxRa8Qwwm0UAULvD3JsVb
pVn2W4/YAE9jiodNMSpang1Pw+EZh886BgfyqkrBeOmicOoAXTuumZh/oLSVRu75
zEHhb9Xl4YOYizfmh4/U/wn0xSt7Wd9nTPKCxdXcRybfeXzFYDOHzdmnO5X947mo
+OOimp2auEs7kyXh7z/JXooUtWmprl4wkVWgVByroZvfl7nQly+v2gQJ/K00A/GP
j9Sq0olaRBrZd5HBmG7K/huWVP0EXFd72ZtBLDWJrdrdR4G4N5nNHkunWmpMBU6u
Cr42tkUQW8QcE+9DdC5KQt5dis60AtrGakjKhzvCzCfqQjUZSoPobKV/Fm97gD7D
0gQw+R8zHrqeWE0cHDtCh1qGQc78Fa4e+jAv9OsR5IJe0ApEgH5h93iENTjwmAiF
bUQDwZqF4YhENb68biCg2th8EVLOSWMYhlPU41vixBEXbYwg6rzXsMaOaAPo4jQk
myhmMsITi/ONUd/qHK+Kdh+rZFdI75pn7ccRrc1eDfhOH7ztkFTBnhbaynWnVIS7
a6nOIP+4P+fog57FnpOmqvY0kCPon92CUDS8U+LIHjLmE5X1HffUEc9eVbgk7ONR
qJU4l50NE+fIRyf6LpJCADvrcyQO/G/FN5YbJTY7z4ac0zENujs0oP6+6mGjsR3y
KUWD5hcqM1dx7GZE4N9P/nETpjTrHaRTuk24ydqyRdD739c93Jc4l0gWJ6jZssXW
iA/jtEHH1QiUoaeblewBRquNu5MymsA8oGvxp9J09p8InH0CB28pL7kmAJKWkQWI
M1gvghvvu4k34ZBIWROcb1YcX0Pdtf1mj3DYTFBCEm+a70+9Rx1U5dLx1c3OwqeY
FWsqljN5iMybaCqpb1OmF6MqgpQTAlBKPiDNYi8fLGn/8l3Ss7oUksOij9RHb9f2
Vh0yy+j4A8Uikr4/LV6FR+L4H6PejytWakeDexR7eVmADqWri+ccp4uIL1wwqFl0
hv/K2Cgwd8mZx+wNBqweg5CzWtX23Nm0PlJONnbho8NinnntD/RA3h5r3xdcsC4H
L588nHuFhwDEWKGJV4Wclg1FhM6XvfPX6x5GFvt/GqNAS18iQgIdJftZZt+yUXED
4e3OGhiTXnHcQFD6ko3lWjjyRzn0fBaXu4ki1Qea6w7rw/Jh1KRr92efyclQnqqh
1O4qn9oZH0u97A+Pv1gs3MDwGnEi8fpqun40VERhjKKeksmUBez89X5tANhnKfJv
2RtdbfruKdEP91Lem88NicpIJlHgt/eqBqEZKP/mYl+pN/kxpONUIeFAPWV0WeFZ
dlXzwCMGw1zJ8v9AX4iVH9evCuTssJNwnMfrvQ2FgkF63rK4ZSPYfdzp9qtS4yvf
mZXimDGEtW1yZdq88JeBupcYMpkxd/5fW4XusvYuDQS4ljPo1i9nCWGdTuKLW761
Ej4eaJKWVrxnznQPKjHeX1g3TpMa4RC75raZIxPbqq1T3FqX0q/VF1P3bwi5ts2k
6pcm54HprRX93/XSUJW8n4VLjJ8b8r6zETDlvJSE4gT0pQG4/WYJk6ae9kk41x2M
I7OM2+rnaKrkB9F8eD0WxdQb5+NumRtTOTDU3iqb2JKL1trEuKD1xqolxbCHcgoO
8m06ea3eG6cVCKnTEIOI80hFCASRiKGhDqAMECD4m8dbPOusYu1F4ldIQ5QQ/jFF
fF716aUDHNZDYX9OlW+olnc/FLd0hYllRa8kCq8x9jDY9eGVaxYkGtlxdfIMtPVu
xvvlWIlrojV2DIUvDWcBo/0M48YfCzptD2lhsI0+YAAGK3dKonaBO64KV3odYewO
SM9I7BFDW8Y6kcbHiFsT9pZjIOCARxHaG86NBGcS1Zsxhc7JSIU/p7+dhi1OBWWA
fh0Dq1trnitbaYAw0z8rmW2iAnG05tgcLY+TC5YxKfpMIRMpXFPhmB/8iE/tjAlQ
562NgWXDbKlOxlyU8SL2a4ScYVYa5XZ2FFc42rJQK/EmuJhmODkYCZyZYP01FLVx
Q1kIiWK2uc3DMIFnIfVcxCL8b6Jy8EdPouMjYaiSBYa68VjCfsu3xuaCt6fcX6Gg
8nqoIGemK/k5ZkAOXVuBJjZrsqKOg/av9jhMJuilX+qMc41MeOBIOiANOjvoQTt+
uyO2Cwq+uieLKxWMo3MWwgkZWx+qZV4TMZ3NLsgL3uLxcis+T1cCTW/cJ56ob+Lz
HZlcoi8o8BYU9trNNDyq0TkBtMMLj99kZGQ7041vXqx7GGt/nt6ZKwweVCLKU0Ls
QucNA8l5nKGtvcBLEz7EBrr+zxFGyUzaFQzFGHHigilrA5JraVaqe971c2GYLxvJ
afFMM37JXnuB38x91gnL0/YSjQVlz1NG5TDKONTCYj6R5Tgn21GiMroEjUPcyA/C
6N5bSjv+x63oqq352VYewluARiFlRWN7FS7QyKnXki0D1kT1+c4EZlvnTYbJaTiJ
j67i6x3xyOsOioarRQRFIgug0EOMsanugSTB2mzfaEeH4xDHtgfGrVYlX02hmvp2
MAUtinJ344/bmB2vq5Gu+R8z3U0LwR0XMGEs4JmtTFG0hCT+U15Wtypvzn8Xq5xe
vcmLuu8x1dnCnMGihZyLHz9qkL7Ritlq6jK1tQe8SLop3rkdC9eMJArhOTBYj2b2
dLXXAfS3gMnde5Q89/lfLYkTiv5Q34Vs7EMO6mJMxVT3lyHb0lr/W9qTXTEAFUoE
1Ia3l2/rooDm489Vod+sDeYmSpE3LdMtIhfcVbaKO6InasfY1kMHX7iWu2wh4NKn
6WHusemGA4W6Uo+UFTQMtPIqXkDexdJFbA3BEv08nyzhA1d9KfJTrK5K/v4JKAMw
SRInT4tR4/vwMenNZeOw3/EwgrD0o08p2iNSGL+/xDmelFKwV1ej5AR2tsiuMRvH
ztV5AdH2IPTe4KDbjnhzCgI2ar9KQl0I5hJwKhJiepm6D7r0Mt5Ik3nOeFLleD83
etVOgyE1kAtdRe2jH7EzWUKJON2Cbf9uwdogfyRuy0tzT8muW9eeCAJV6rEfqaRz
iEPWbq+yB7uSXeRmFACxLSvmKGSOZxkguUItDsJt5r6aBkQB0LeFbhid1ma0/Ea6
OT39PTfblAvTMgfq52tpMLJKq2Ay8m2Vbwk9QbljRDpnI7M3oaHtPjTw5V30bClM
tE6cilud0/+31dHZyBiV+/dzCwEmWBbwOYE41Bl+F0pRrc3gwb4tWreYG4S+7QoU
yDSfjMGBG5gtUHiCtESRSQ5mxwhKZcjhUqr0ZYBzbHpGI2adhQFxLltqedb+1gDh
Rn1jp/SQ4+yq4F29v0Ih/M0CjZ1Zgw88ITwM348q5me9S5TFYWvErtVR2WyQiR7y
YbmCGxPlD4DYNm7ErDsOq61b29gEaLdwTW3mApl/+hiOMAMN8KcA2iF4s5kRI0+N
fqUmnG8K+VvXwBHwuzynHQPFLwf7uJXq50m9D9QluGAu6nqnAl8J+Cq/xYzv+n05
GndLBQvoxBj2wed4XRzAC//o/zor5bH6kttaiNkPJLVFV++RcdwX6VE8CGktNGkj
VlSBStjxGWK3rw4+Ascv9EAmSMoxnqoDx6gf0XyF/hS6tz+R9QfR+LKqiG5ZAwTR
4Yxmnpy+xYIdL/9nHt402ykUMqO3tckJ6o2U5zadwF1bnEOhAwz9UAWDCxRoztdb
crSrxNL09ZvXjDn7vzwoN2qvHswZcIsrts+gM8R1nwEvhX9fXkZrky4sLQrE4Mgg
OHvv81rd1kOQLRBRl9nFf11hYFvRKBfMDEqVXPvf09Gp6Oie0t7u6E3BeXey5HE1
vYu+uAUbU4Y4kfy3TXvoFI9JmYj7/KJC+iSvq+KY6g4J5RL/KvbDHCyBQ6J4N2jX
PB/XXkGS8iFG0LWuF7rDRjdjz1dZCoy1m/XsUgXdKOyDHR7t54WwQhX9hJLQbWJ6
JSf/YQUZa6TxmeFhr66SysV+sF7oZQhauGIj+l472z5CpJnp6MPHsavcqMd4QNbs
qaAfM8iWOFM0WLJhFa3nqG0uil9BdX+EFaqSaeGpatHDFJA4dWVXh6PqA3MhSH3q
GfLZI84JlBS5Vg4O4HJd5iGoB3mWdo3W23cRNgPQKZKgJp0wUx/zr2w40NlxAuU9
oAx7nC9X/zdgEdK1X8enqB1tuZxalgkhXAwjtgT7Vp2FD+w6nRgUMhv6VewSYpum
qjFqFW0LVgdTiVGuSLTroiIIuIWeivHOFaSwf0vXyfFqLSHsO5kQwa+wikZIwyA4
ceVIL08fZgNUk2sTbJXDB/UADqYrk9hkGKFNIr//w86Ejf8BQ2IAUuiCVhlOBBFX
sisQJWcOeSHeetn5ZI4kqfB5XxUyQFDMZ52QlT+HxBYvvxYgWhkWD2Uc3FJTtrwI
WCNS4bpusoDb7SBHESBjaxp4Ro0qjZOlZhMYBGVuNnpxKdA7Jhclbz1ihCMlL/je
ZcvQYTzv21twiWvcfZ7rLT7snEJQ6YBPmLY1TdfPSLx2stPzjyHpg87HsV2Pc8nT
WDRxt+93A2npZiDeXwt9W0aevJk4j8Hiy7wJ5Wabbo0UWB9zjCFjR6Myk30HYieM
Xw7lHYlwKDl/BMAkZXaNo22W7MS9Gy7Qj9YkJHCIXSGI4hqbr35YPwOKuRCL4RVF
pWDdH5D9bL9AZRP2wpsM7iZu5fEMW2Cir/AcVM3lifuM5HsDO7aa7PMKsbHZ5qfG
1TY87vHRc1C5G8r4SEKHCRYYsMB8ZP+esZ08MnKn6eTPj5DEx5CgfMkLV4/HRx6l
gHvRWz8UWQqhaIlOTEVZexgNw10kJIzvStGOBMTwrwNPbwDkVhPq1Jx5yBPwLEAP
STwf17/W6224LiAwmJkkBOgx0tSiJZ7X11x2w2zlthpP+fBDg+Yd8+0NAkH/a9Us
2JVEw4DpvzuDUyDSBO747RmiV+FX9fzv99ilaxy2V0xS5kbFzg2EwLVZrVHec+SO
I8NOMnUqN8ePFayzZBwiPC9JN+COE2Cb2OKK4sa6PHc1JtCU/PoQBcEJa39nBgVw
ehtjM7ynSpnlkxdelWpFtUdXuUpIl8heapO9zSOnGSIzlgyMAI6x1R07+6CztMdd
01pv36xPdtEJarZ7vdErHjb5V0B7+PMhfnvjnm69qDAU8b2yu3UleWvHvCg2fx54
u7Qz+GKrmUaklygS/dNg55ZPUZJSmyuFf75A+206Wq0uJRB2tfqiHDAuAUYJafij
gtWSwX5jQDjrE5FmyX6mwtKmC6y1Ny0hAVVaneV4txJJsAuabrmtMhlKdc7MyG3b
3PuP7k1XnBKxIzACAAhipFNGsGtniuUiiZbENR5Go6Q8fmihWTdpP7mnJ/YKOjHp
ShhihmicgbR7mbCD8APYn3VM3n2w7K54meVTFvzygFcR1rCjEu6hrneWWe75xYU+
TYGdXYGaRpGuCw7LRuUjiMxc4Jtm8GPGxY952fXW/HIPD2xltUcem9XVJM9ox6ih
6N2elXh+VyRDefsxHTe0cYZ9VXtmhvbYRWkrkRIxmOQtRuFc23p89LYfyHbq06XN
EztDCqHl8nuGFbkERdZRpod+C+YuZcJu7+XZ5kMKMJMDayOwR34zrwLGVa4iOfgu
xrs2hQHvVfLoW8PMmqe6/7M4wcqjk14OjG92haJovv8AfTjl8EoPekh6M4B0VxqF
XIi15fD4+UQZIF4Z4zoMSgXU4xATp/7DFNMXjfEDms9h1MCvsUDY4a4RPHJ3Snwc
ZtMHvLgnT1HM/kYpo9t2RT/cQBce7EicAJvawax6I28djvRSqgrOXydwZCKeKbHn
ujD03iKZkhUcrUPlB1VbH/vu88j2vt18CzRfg0GNIa6u8hHC8p0/nlunLJKaLaFP
snbF6T1UjqD7aFfIZ4gehS/dds8G3g1rbSanz3cLUGyglfloW2GXwBglFvSuiWQY
`protect END_PROTECTED
