`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4m/b3DI09n+PRAbZPouJIZSP9ZSAUbAVAuzQBYtlUStYJDDECHJMJMCjD6FCQt/x
QYPbHmiyHkw2zzrI2fxUBxfUywoqoXbE07KclvWiWCZszdzT3s1DRMuWDxeBrIv6
zrPdP66dw/ARKHJB34odfYwg/sZTIfBVNbhn51HPp+3mHu8KKoiBkL6rHmmmFvkq
Qs/0Q/4rxkuDnmUKCNo5iQ7i1gZx7u+C+eNGdfmh59vf171KNyBWl3vXmU9QLGX+
asBDdpk4N1eV5JPc1y+dwzqeZQJ23440JkvpvFSlolQLs2RZ3EXmDS0v2ipKbYgy
d+BMGRU7BAMvXGwPz767ecsWlgikNDm71qCUuiRKvJ1GDYZSph1f3zaUZik9MBaL
ADS2IO8I6RFSFf3czi8qiKrH49W6Rt4Ai+mSRDN2mIo+lFwLz4UoBsHt7KvBJYuw
X8O/LIhERR8yhSO3ulNBPWicBekQ4u2Zni469E14BDmdVGCYdFBzTQkuPV5rd5jl
iEV3zqNsni5kwuB2zyCl3gJp13JKWKX+KjB+p3U/aNOwMKytFA1L0DXi9D+Qbnas
vfjJ5fkJ8iwGbLkZF/8ZRCK7clGBAz6Qfh/dSE3u59oy5gmu1hnN20KfDOyiuPjc
wPNN/bbS0qZ/PMzFXPY3iHDgR4bJuExUbiJE773Y5ZIeyEjpjNTc//0rcuVkcjBc
DGM7PR+B20jcb8OXFgKYbPoKtqW2yCbfUYTcZUh6cfBJIsfHT/03WNaNorAT6lGj
7TyFD9tP467IDNBUzjE8++KQCXPcFev/iiue6zKPASD7GRIjn/oMijFvhq8dsHdO
B2lRd0apoXzpchVZ5YKPDoRrY8HfIUFllCrBiSPVTaRE8lE6bl8/sXQAu4iCMeMv
Wvgi4nUjoHI4ncE6xTYw3uSzN8ezAgVoXlrQkiI342qRF0oN2JJ8EMM/SQpi99cI
yaR4li2h4juc8hOzUwNC0JW/bm3oHZ/3h0uaTQQ1/0a6+mbxK2GpZvKAeG3u5of5
73shn6F+w/pBMDDm6+mLxENtfUUOCfVPJeJT6VJ6FW3Fx6b5L/D54SC4/4eBHAdW
u1uA8YcIJ1U3VOMPRalYRH+earyLKwfiokVyuPjDB5fnCJPwIl6M3CJQbhd9A8f/
PLm1x3iIJeteAHdbi8idw9DkegdQEA08C1rT0pMmbfN3Ds1Gc8vf32n2I4cOLr9O
JuSwfC85ilRu05EkAN0+ZNDJ5n2yb324D2dYWw99wUQMtIkidkdZiK70viTlgMyz
XAB98PzVclK5CuQ90nYKtLZ7kUUiy8KcJM07+cMKI0ii7mJJ+Z5Mg5hG55Yf6tHH
VbDocgtM4s3HFT/jN4fRyw==
`protect END_PROTECTED
