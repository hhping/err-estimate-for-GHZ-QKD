`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9PnWV42DKjfMEQx3vlknMuNGoQmqtPLkieiunKk+GThCKDSAq2tBn537RMo932v6
bvUvsGFQAfhg/dgO/JRL/Za+3iPSHzMEODaVL3O62LAEDu7jRZIlshUuWn3xxqU+
pFe6gT9MlsRA5MCtWJSE6NalyX3ZolJZ2RkZooBG5oYUooMx7r0G79MjmUCWxxHa
5ds78vq3V2D7vEAHk9uxJziR6aXYzSZSSMNCmZP1ILA/yHaJ0uBihNoyfD8MBFVe
KMyQTXD6dvheTiLKf5HRWNj6JFts1mxDBiGGjp+sOWMfuE3c9lsDK+J6gjgBfvyY
H4HBote1/BCw4qxXXt8ZrqzxUI43drSQWHXTnBlGmFFcx/z44EX9V0Jzh0DtZHvd
AhE3P4Hr2w3pFPHNThC83dwgXNHYir+OzmdudHsYgm/RwA2ZrOjXHvLH/vOXOBt0
A2zzZBX2Ta2hYnsTxTYUeYV6Y6e7vJsJTK98nJsoR0nZ3tg3eLWiTBHjCvNVr60g
xK+8ifer76SNmK/oPGHGzdBf7nQHLDoEKP10iHazRh0oxmbGeoEygF3VZrcq0gZ0
AHDgVIuR5ep6MLJwfsIeUXghy/xATBbFAqfmIa0oltYg8Kffz3O73Rvqwoc6NAil
DhJDezyCtjnMtzKkhW2u81RlCjQrfEEWzdb1QQ0yHG0cq+z5SczYADEsYf8Aezg/
DLJZwYsFsS14qwxKext1zCJ01zbiN+Be9941Db/pGyT4h/KlTCukX31owUarNz3A
gCHo/DktMNiThjS3N4i4Xh7FO4TrPNKd/Wr0GfGn6SObiFWJ+JCZzmXJ+Q476hJ5
bRDzCPXG60mmqtsOZV8lbttOzBDiuxU9mclxNSV281oNtopZPanFyPLb2TTp/x9H
3aZphD7C9/iZtSljpEw6f9GuwCGGh11pHBRJm+Us4V/ONlwo0vhR9i0f075bqH23
aF5/Crm+fuuumJPFLQiqXv+M6/AgYNgcaNmQPQgx8lpggvMKwQ9/Ds/wmPoGLswV
l9c7DeBxoylkaul1RyVPpZHczOlzZo56Quaee8F9eSygxWf2wTRIARrFgpP5Drp4
A1M/6TBRIaVygLrKSvm+YfL29Wl6MD6MtMM9aT5rHzNtSnp1ocfKhfbPKl8pssqq
6WEtxNJwJ55/I/zTii5vEF2MJadEdCHgCV7xTnAECumxYZS8d5h73l9LQcpjqHgk
WPec9dTwEbQnyEGCzAXHNLSJJK6gg1SD0//h2wVVvtkb3+9j52X4SoQ80mADEJcP
YZuwEN4I1i4ZTI0wuoxK5+d94bbGYsy6/kY9mqhlqF9IHxmxBopD2lOKAhvK/JbS
MQGNEL6ymQ0idpLXHxpEf8f9aNk9RLXdgO9r3P5DT/+hq61xhOZGXUmaIBxGriny
ze7+0QgSDA/57Rgv6DXL/lDYeJRmkqwWSMNn68MeClB9xUg4+ipapOKxspiTCS4A
vo0gwTONq+fimdy85ugM5YlkQIi1jYXQywSX1CpedTEGq1o4Hb0ATfukk0EUyl8s
buHtgeSBvkMYCMlzIrN9zU+aZA0aBlWtg0vPmSldr41eKkPhAf9eHUvmm6wPNt10
9zuilWHFDNsSQXRohIxcI+gzvJiAM6rwylbdpEX/WA14a3LTkzjR+39Jpl16ddSj
jucUV6MdMla2uBuwWlpTecyaLmI5HHZR1UMwMix1NFJpeMuZ+iBS33KHQjiEofsx
xySR3cvNRHOROZ4Zm7VyOrzmny5J4EwvZOnYeZWuULXEg54psY0E58weuHIFAalG
q5yWTZUAb3CE5AbWiAqoJxGe89l+EwtJmfjpW9HI70LJA94cJiOsUei4Cfc1vMKq
AtOAyLv6eSn6l9OPNfFf9es54mNGnRP01qEo79hTpRss93AfElXV2Gm4QE1M0kiC
yfhNQcHAAM644Vpwy3Xo6A2X9WrpSt7QJsKDaoLgtfWzOBLg1KOSDPq5UAIxprz0
nWCY7fWj1fR1nGl8mHTsuS6VQkJAfRG2pXXNOWMcUXnR8X5Nxlelpyva4t37Dyzu
Wnr05AEGIb3NA7Jv1/2VRN0j2Yw6rQJM7RXIWMUwnBLOYuWQkxV1ZIsOjvlhAqVr
cmBgjy4JIswzn9xcrmR9JUWJELZtRKKfx1Ucc6VUngGyMdHnmiHjzoQd30z3Hssi
sOhm+TS/qWMC58YWCuw9QEpSBhhCCURys/yvhxO+7Fc6QkB03VW/jcyO7rNA7dak
IYyoN9vmj/oOINMVKS0OlgcfLv5VNUVZKoVWDIykYoztqewOlL3jc520Va6P0pmD
ma/3HM3ujpiWj012sQRyXgCRwVEZsIQtWh/rM/DDJIvp/tJYeLQ+nPsSZlIrWVIW
AQxKziRmOu/7AryFX2eUENGFIgtduJROqjxZcepGMZ3YaqHcpc5QdLr3ktEk2yjW
XBVxk1U6auXL7UsZawV4ygfF3DZnmM7/1Kvne9KynPjiD564a/+e9TcmYszBhCNT
BPfayCtgInkWUIf0aTO71r/yGVoy4TfJ+JteGtElfHlKc5ZqvMyt0h3lGtYPAJVu
nI2yt6RIXoUQUg8FpdFQBDwMv2ymmQ+BRINB0po3wx2flPiv0B4qR2mSr/J+erOM
BR+e1SJJ+TmqUpTV5gZtF7tfvT6uB7Y/+UXWEHx3S/aSqxgVSGdtR4wlCPmwwq0r
TUfFHrfZ/WIgznOQfigTT86b8jOfu5SliYUTEhVXmSi4j9rxkGra+d9kVSiQCXDr
3Dhi1mv7hT1SjyifUM+M7Dt0ukVXe2knziw1oLPHtVOuoF+XK77exqLDy8tMXmdn
jMNs4OGa084D4eHg9xC29e0jgqosqytE7j65eGFiTUyzFQKQ+77H1MZKLjUlztJ2
kVGOmb5BWftM26fjZun08DtfyMgo39P2oSzec0Br6msVkprIOBAtS6TF2f0skS+a
imDFV2ihPVx6S2frApCJbLczPSxkBFrVRGwvw/PwFn8IZP9pqvoTQ/dDCP0cggG+
YQOkxf0GwbdQxg+VzWIRpgpW7pvrb8gNUaxGKlNB2EdcugsIwLaApgkLW7bMyP1Z
GCgVxp1Q5CeQdr6d0f6G6W0ryA2LehbbGyW6xtvclNI35tWjjNhZxkVeG2Jr2Mqe
PHCOUlcGNqPms1gadiwCFTEGNXbx49DwA9VWkWaaeMYk5lvn0S4wG9IBFO87Ztd0
vtXLmM7wEtRu2wN4aLdRzNHZ6JEBuaK4YgOdCeXFq91aJM2VsUmmH8DCJ5pwLrQX
hQo2xtqaWnvM8KZ1mQLATBQVHI5TXN4R2UGFRHqopKriW282uP8QhCTqq4EXsnpO
7v6LhAO6dJxcRj/o+hCpJjSd6Xjlbo2oXS7lIV0VFEWfEuHCewMbCcXGcONI6I60
JHuwyemDorNaM6FdvPbmxW4dpDST439bWWEtktwZUWo6TIuzIr/e77lObTEOoQBL
S51Bm4ZvtqPsa72GROMnWir2otSU+nKTiKmlMmDV5pA0ZPomKQVdvNdjMIG4RPI/
QGpwVLduiXNPiZYgB9tJTeMDz8CV1sokcb1cvqbT8G3n8OMWEU83bVDTixl5rtGl
eR2nHnG0hsIcjpnXgnvi6gUCRimYXkjJLvrpJWBMGqoKbTdBMmnnpj1JiU8Dlf8L
kINFRYI+lkBnKbrhps/bNDEwv8fSxvFjG4WI54EsuW1UP9R+tDSE0Clgy/1N/YeU
jRhdDvmXlrW3xvzVGHOsEGlh0F5dFXK35qaI+ZVfIyl8B1NLUlshAl/C5XKMUSzC
ma0R5vgMWsf4Vg3yN1YwvMU3WX+rp3YNbV60nsWrKibzUzYjUe9skRoiVc80wfqv
WKers5g2Bvh1F+QAyLrPrvwL8L6z1ljvUsgtUA4fOQcKZAoQaGUHJJsXTm4Mx5fV
HlY2MhDeOnPrX9zK0ZT+gTPE3z5A/YIonmClNMu3RuzHWkx7KrUxlD+vu0PCi64O
Gut6dVioHBXLVPBCeBZQ2bKVh4Uin6T/bSTCOc+P5RCkvJZ2UfrbksguKHZ0M4Ek
9jMepBuKkgq86J+KD4vpEWsj3o3bkee1ZkKDu2QClwJEn0CxjHYHQrvFkbdhcXey
MVtPc2h8qSH5G5NBCiJp0QH8UNqL4owjc8s1K+7z+vwAn14nWQVJxfasSADvoCLO
2ql6drHZAHLZxsRe+OSk1AH/mKKqwhuk/Aj0baIH35h6GpG0OLCh6S/5em7t5nhf
lxG2e8z7N9poZw12neETlx+3uSP4rSoCYdAEH4pnVXI0ml87gncd4okenHD9XLoL
45looKBjZ+UCLtwdNys9NRZeEWnMDPDjYepZ+0SRDVOQK1J+BJnGUyG/9wOuYsg/
P1Jk8S0sZEHYuivtVrbjOwpvwXaZ2KRcw/YF+6nS3/JIqrfzhZTmEGMAHhmO8exx
wl8sO95RHfsQ43OfydCCzW+r+mnJ3/2evR/qzKF7Y+P12v1ivT6+ZoOzoVPjjIYg
FqYuXe1RYdt1P6ESqScydsG9l4hUsd2GncXCdMg8TuQwektDg1gFyvuBEvjoRsrv
ZTKijUSgSXH3DxXNwaohhD0/t14+Tkmy+xpAUItV9qyGn04dLlpQpWdm5P8D/7fh
gIy+9zK62e2x0NI2dg5YOtXpsIgqkdaADqmGvp8YWJNlzE8kqhkWo6GJJUopaG+2
kl2zBYDT59f66tJB3YdXbYiDL2AgHe5NVb6nISxPU5juj9bRLVYfY/oAQHE4OijE
alvfyWCXBOTKeebvgpG1hmRXLeh3eURzdzxuzpo9KmUDAOG6H7GyW3YIAvPFjif4
jcRptSO6g3mE7fA0u3Foa/C1bm6Ia/Gu3wm8WqUyUegX07FK9VY8XcboqHlrccay
AdsUTsS1itGLtlm2GI0q0zLqWfUvwTg69fBHWXh5x8EjmkbmeO03tI7TWosUrBSv
Xbwc+leOQKNlVAWtO7XCh14w0YUi0Pfxx46n750zRMiZE3Y2inJM0B8biPi2Tt6U
qaxg6KIVPMFfFNeeOFbY8FH1AgLQ+PEhN8zrUlMBkTUSxeg1IPISaLhrXCa1anlR
6b4TatYOCEfFIF2EtK0v/kZAvlhARIBlPy0gou36G1KzcrrAS+/q4yFchcZqJ8jJ
aktMz0JPJoohP3SeH3a7c8N6WrcAiY9p5Iq58kOi22Ct0KpA6oyTPQyVswuao+N1
VMdD7xmd7HgRPtOU6oT8eSexe3HGouci/Peylqqniy+Ox8oC/QBICmKwBLLd7QdX
KVjRvDajpDjW/C6R2rpFe2M6Lb9XdpYAYZOGtzN7XE+Wp50Vu0bRxyieILURSdHa
f/YN07pbN9Gy+SeYDf1hzUcnFwFZ2h8AARdla26OzXMCNVPtl64oFKaJN918s7M/
7s9JxEfzlcQafZyOwiiB9bzEcOLEP29nga5FI9RL8cjHi1EwkAztncvPfXSU4M7P
g1yeSzZIg2LV0NPVIpGoFztKBduhtr+d3LKgQ2VsevV69y+0JJTgJyONif3RwioJ
Aq8ZEe0d8R2Qr6Exk2SZmmMCuLMcyT4WsQ0IHMZjvzm66vQwoATK6VwAggxr+xTR
tYFFVa8uROR4bK6OodqzH9YnM2Bg6mOxcqFkWyH1X9Q7ASQuCHyLw+JWVHqyanRH
EIZE6NsTadISY8EEN8kNgpWPyvwTnhHWdpTl3kCwVX66BKsElPWm9d3vJWGyeSgO
qttTc4jxtaVR61LNaLU54iClbHhm17G9l3eupwVFpm1bhay4D9W4gHAKWx8bsZMt
uXEFc2i+Y6hEVasNIiWee2UqF7hM8lB1WzKWBTPV3CE6GkZ3mrstLHHi7Ue0l+5q
/3p6UxAr5v3nn4b2FDzSLJxrF0DtmfyfFB1bXibgrsWQ4FL4YjETcwO1QP7fB0XZ
78ljrTKu3fw8SFgSgSXkEN4aYYlZ0F7CynfOQez71HHa/WpR5yJzWAMFvGNIhSmn
5yogvnZYpK+RgvrTUjYoFrnikHmS1mLrhe+MgswIQqDphb0x9WHWc/+J2Yavodi7
NrKmDpBcTCbBg7NB5ybWFEMydqrN0unwd+n83fGEEyMyUbD4C0tv5kDBgKJeFN3B
geqxEoeLjlpOuGP8Gobhs2oyhxRJYQ2nhfzsOpJ6lbCCQ1V712T9GmM+k0m3WBn+
2nK6dpVUDdXORZYNYt6PEZ88mw7QU3vpD8XElflrhQtLTGlnk0pcsUCgRneHzZTt
wX3aOYtI1O+THV04cAZUDxCAhOlLqT63DIXkV+Ta7Y5pRJf7dBeNQQEJIG5vWiJx
NkSsN84321UQNcW3bIeGIFla+4Hch4J0u6+H9f3RajlVr8jjvQgKcuUKxNAYyG9O
ShsazGDqZkUgj9UXTKLYWa1U7J76vmx9C1gwt/2bjHQJe1gftCpeRf/p1eOeAiVH
UjNiqQfaLP75cd2b+epHMDZXddnOf5rM79xMJqHXZomeqT3kqOrvQx/sRKqoPMiV
gVA4Ag0iBSHP4IvIizvk/FAS4tnFvR7INMIBHYo4kQ3wFrrBzMXSxLEuguzfdCp7
15SS1B3Pu0IcDRdzq2ed+Awwti5fmCqaPD0oGds6SjTmpr68UkOJGKKbUSk2lxih
ZNfFwlwcEJqZcpBivBl9OB6ZtDO64Avc8WpTKpSkpEAx5HpR+kfl4Hsr0zFkCkrZ
QPTdP2//EYPbwCWbRjJLoIj8DwZXqv+/8CMvSrggsAAEoyyC6R9XLeBAmW16Xfq7
TpbKIjJseo8ATWH4MOWqsX1b79l0e+SmqfQrCV/gbQ5MP4g60j7wNVZLI86iFfJJ
PPBwQyue5x0GLwUDyA/eqQHd2F7y+fC5F/2oiRQ3Wa4J1yE24Yj3tCBux7GvOXD+
QOOMo1+WQzqXj35cTpWzeXSkKYY14WT0eDcOIocE2xqWnY1ao+icMcu7yKSveNoZ
6N0R5WTzxl/LJZL2HhmE/KCxu3nSY37cP0JeCzH6jtTnSTyu9KFQm38/MIZkUtdk
YI+tH5KtD60mf/eLdJkFuFZm7iS2XcQDk2/GBGIvpQI7Qeww++nQGJDPhewq0/ey
wWZwY0pIN/xUksQYLmxXAPdSOfdMFz8WN+I5OqqFJDE/II8YJCoP3hbZjA9aj3TA
VrIGWUEYUsEAiC5bcW1rhsuWFZ5GKdkAJ5DxV7KEiOChT1Wa838A8EHc92LTyzO7
CNBPtQkDX8njycGr82FDByeb1Pou1r/PxoDg87a9t0FzmaM0gmcvjN+/drTXLwVX
RSevCZUkCW9yOiib9pIyQWuhnGEuEAwb5ZqFnt+TkvPiIjBslCMTtEZS8eSIvnUs
7H8Mq6XRJVHIn0nexgLEyLXN7VusjZSGofG8zR+yCisPvQGc9o+CiFsFlpdok0xh
CFJQi+xtf/64bRraMluduQ==
`protect END_PROTECTED
