`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bsBi6HQRSg8OL9bUlwCCMMCRgkF8CfU7kwoM1VYgffD3u7+9SC8o0e0MGvHZAwf7
zXhaMtW/WxsinV6DW4yT+ADbjMvzv99gzRt8k8f2MCL49S6LjAJ4ZFjHEde9sbCD
eVbw838y7NLTWsw+1gBky7ra/W36mIwyJ7PW2YDphAqmszKqCwmkI5MHR7kYk6sc
bwSliCciQuhaWqDnIg0OKP7Lj44S9XGb7zgex2R9+0ziJapYbsKlKlUlRciKD3k0
HRko/K9HhTJ/b3woYW1HnPwyZiFT6L3iYugTfxHkH8bveeeJn8jtaxuQ/BIhTsY5
c7tF0lF4Gv3egkVeXqHptjmfV8jt7ukFReO0Lg9D2Yt0d6s6PrZdGu3BCpvJHRQj
q7BsXWASEIDhFydlG0szTmiVo2aCSFMuNXOwV1WSYigJGaRZwPY8uP6qmSbRmfLw
73SU2kS1e9SVhvYsYyqiqzl/sGKKECE7ELQhL2OqFfOO59XnfFKpQmHdYles7wRy
dc1ADaR0ZgN+UkX5ini7crFt3RzrEy71ltE2GzMjRS5KFrqCDRyWcWZq5FIJq2P7
VcSU/CiYe7oZyzmtuto0G8KL0+92M0ISwEHMofw5jrWbqpxA32QlTTW3V9yAQlWu
fKpmqH40ySCm3Qv17zwKIvc1YLTsebEAYUu362KAoeotFN8IE1NQT+TTJPypmnto
/BktJGeYl+wFiHBw9zyeJXmhok7TUvnjdtqp9P1Brw9DqZZ+xyaSMsAgGHjnqn1Z
ebc0pTprj9D8hZRaE07ajIAwAieNI93scAaMvssSY1H+5+YuWOyAKkCFPd+mfOhQ
+UaB+FEu5fV1Fx6DaYpk0p24GlptQtKA6/KlbK9NOsF4AYc2UVKZ131DHX9MAaG/
PAQ2KBmbg7oYKNMVBGWIrZ0zQoXmaESZABMtTinD++zh3ybJdSYH0WrgxkK0Mxmf
7j+nUuDDSJkHteXMPgNX/YevG8X/tfJzibEQh+UrutHUKOfg2eQN05h4lQemu62G
+bv/uywERgwZLk8fIEinZeF7DULV0phkN/Ecrey/kePWQ0Kpow/91DmU0bxYwiAP
tOmFaCGzqQfp9+pinBi4HQYL05Qu+N/eaopW29FPydhutEkzrZOeoSmxx75SA18e
xNzkhG7MhUaADeFZHV5X0AR23xKaMWC9IwCgy0lRegu1OTdV1cOwmCJ9nDV8oB21
PwF3GgvMIiXoRwhdkdbBX4C8pQZqFYE6lzQkCSyGIngeuVVLiEYLMBRjprYQJ+sL
6Vk1+xPDtbAeySY18OHnlWw7XGQZTwuZRmF/zmmVxk94BqG+VXvwSJesC68GdGyp
A3vVjLPKhJncIWCc1ELW6DsFrxqPsGpLOlPb16csRDZHyxpZ5NApN7CSswoWTuNr
jWMooGQjZLPsrzByr4SESOGR1fBE+JeUYWHtnNv0BPqLGeKXayIzYw7tjJ9wCj7J
cA4ZO9Gb5SlFW6Fjxx4tuB5LC9jVzp0QjikYdfaWMCVH/qjOLMw9wugxsW7zrNYw
KYvXhHTNUBtjL+4XNMfjb8I4auHHpmoRL5thPC18OsZIZDdG9w8LxrAlstzF2WLc
L21Ez31u2zilto0b2gm79yIlbz0z6n62nXefYs3bBFOpghZAutl74i2a/8Qf5jj8
1fs45TmFZINo9HP+4E0f0u1EdokxaFhmiGfvp+4vg+2nJy96Ivh0BUbKr+N7pLNS
F7F5Aq2LN8Fss3fkWjfGIGqO9LgFhWojlrcov0yLKj2twa8QtsJTtCrMx6i1FG5q
+4eaR6yl/9GEVIDmZ6w31UCI0rDAU2KiHDBq7jMhVgnakVNxAXVBsR6pV7udrPWy
ElH6WwdzWTByyuf7WVioQrPWYJ2cctCtsn+ceiNAZaTLW4QkHGEy++2ADQa5xOp3
IkRs7jqcXeISyd3fMahHVRow5esYw22Dy5th7OcII6pzhQj+as2eBy0SutWHHsFP
OAtbhTVIylIOd7ltMaG1ZJGkPuH0WtatsX9L9V7A72mYlJHMOwgZYQdKQTwDlMy7
tCq8FtS998D7zeMsu5w09Sv3GXQ2qbUZjgK8se5SdUVmPDkZs1iAAAWSLRWp4J1d
iak52gs9kEZ9vQgpGmNG9x/E6+JjygoAb9Xp8cqJq09yXqorWoLLZ4QkydqBlYlR
rsEym2gP/g8XiwLdth/hqwD9j5NHn1CNQAZNvBKesPtLlrxcVzlNdWvj5a0cKIF5
r4L0WH4AKOSzfLhOWlZCcTXGBRMDQrW2bD9C0DFr07IvSqQ0go7NTinW00/Dw95X
K+TG1PI99Q5q1n96Qfw3Hte4Kr1ZmG0A2xmUTluTrAEMrY1KHrxsXnyso5Ga+Oov
fFi2jk2g4XVILZqSYGJ4rkCTK9GVU17XLxGwBEBg67mRYeCnaTMmEeC93+Bpd0CY
pyW3RkEl9rlgI4Fh7Y9C8g5lv4tARfLhtr2/zshbzKZoCSSzHMPwtV+EOzmQHsAn
m1wf3hq1oTHk18J2jAbOyT4sxXexOeEdH/8IOW9ZxlhViIUgscCbVByDANWXuRsm
8hiTtb1sRMWarKIqaBpKp6cR0FQXEEq6uGgS1M7x73mPS4m+FOupIlerpaDTfJV1
MoGWtqI2pVZaAiGolfVhz4Txzrxe1Z7Saobi/dDa6KxC6jQPQ4bIv17IlNDqTTXm
jSti9K46khAe1kl7aE6L7gwoi6fP/Hw5SXjzwzOGBgI2Bhm+4jU+wm2D24lQ00IZ
ByGky6iYFVZXg7WOGQewoW+xSMsdxeU6HdFKv2Y+0HsNWbO0YQERaA682dYEbNwd
iWM/RbrTfApZWtJiPZBkZDv5oSNfAP6qyG1cZaORtjOL5H2hacQuSRpC8R0qdRpL
9uAucCtaD+cLb5NU9lh5KXWL2WfzEEEkk1/Jdf8QRQms0qF1tuYxCvBHSGstRhmg
bXSohsE1Ep4Yd0Sfg0YNcAVCUe4YbfYTQC42+6mJk/5t9y/VAIu5zla0VPI+kyl7
CjAc0giZLrchE9Ac7wjipqxOJINYrnPCKRF8EbqDZ+fmPoaJqEWvnb6hE1MYi4Xt
/sBs14FtJwpRU/iOvUBcmks3qiiLfTOuOYTH+5mwBfn0c6w6CA9JaUPvwR2dYbhQ
otZdSkI43YwFsot6f+yb/t5mVQWyKAI2OhxKuU9w2BDWkLXCI6RfN0TKiq7r9nOz
vB7t5OqX9sa1ZAM5RXTmLA==
`protect END_PROTECTED
