`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h4OcuugVZxUkgHdP6JhIsEEcDnfU7MguuC5NZIcqovSow6HH5nF9AcvdhPSERUzd
YEN0CfKOaV3E64/u6prPviE5P4bXMV1XhLGxC9vsCbLvMushpLFZWvGjBZDd2YqQ
BdspA9Un7hVgQnkVabmSctG7W20SytyvF0aXCY9yoj9RQyloG8Wyv3g6Yj+fO1Xc
LfzGI5Gtwrawy5hfi/X+hDtJqxX82Cm3u6VfowEfYHIF2K6hVBESmPNl+15Dws49
dixBJUaczotQBw2yQLA8c1snOlskbFxhrD/FhiEOQF33CrXqzpH/EaOzkrb6VBd5
Z6I7Z22wEiB+B+TviF0hQGZVsZcO+fG2XgDG1vUUOy7KtKO2NmBGhM+2/t9R5HMD
RMe2YK8d95jPn9HkcfzceGhNaG5AwrjEJRAxZeZ6KW2Y9w1TN5LSyD+yGrxYvYBE
NL20r/q8OWKf55EtKhG9n4QU30ZOOmhoftQ42iqx05IZ69sBflGJfqOjc8W3ExJw
bOCBt7fEVEbK+zDkMJY4b3NKdwzcCpNT4eiOpl75tdm9mVcsewCatjbEO+UkMhb5
bKYBwJDHcMUwMNS80ZQpovm/y3zRqPFm99Dsr2JtIgWRZSQkoWuzXOppvWBc2sm0
XoxrFH+1lXOYvvqulDcClwektzGGc4rVr/qg4Lq2nEzYHdhjYUdzD9K2LmaxTmcK
OXyFUZi3tEHwDDSgE6FR5Wwrs+D5uaxWq2Nmeto8+Uvyc27Lpc9S7zHHqmw5V/xG
`protect END_PROTECTED
