`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pmCADWqz54r2R6SlvVTrIj3Z32Id6/Nb5OiR/XkkZgkr5YIoNOLYmtw+ZbKFZLez
o6+lNFVvTvASmhE7ODWgSMhXc1TTrrayf3JXIiCnNnH6vBbf2y5PZVJW07mWuinp
WKNeWmZuEsHsr6uW0mHN/O4XK/1Cq4JBkxazTemPAljciQcbIU1LVySXLNHzVddn
HUwscQFktw2o+b0W3+k0uGaJ8GNk5vF4gMFVXotoWTGeOZKR3+e9DV96ZluXGy6Z
Pj+j+A2E1VbMSOzuOHsxJpbIzSMNa9Kp9JhIua3l+QwTKtN7FKeyTBUOemTrJAC6
EUMoNP/feM715HHMs6zH/X6kNlS3OtHbUqZBjcazGG0ZY61JWxTOFCypcb3uWFEl
9ISwXlWWbij9ysfMWQcIIoIC4fUiuTMA67ona+9y9BTbaA2i6EbiXqcX6mgnBlnW
wETQfzvG7xKGvghxtRINJWzeLX66WNAjCTstkae5PU+E++afG9Ot9Ta0KTJC3RBw
zBkKOPQ94lbV6sftYN5ws+3YfzuApyksuvg5bPiNkBRXJNwrgt+bnfUrZSuRZf7C
tuR44lhmjq5ygs0NfzX2+Hob/NenYfdxq3KREUiwbGZuY1Co5CO35qejw1U0a23N
xp23I7C8KxkD6YySntY/0e+irljRrbEqnAN+reoZEgv/Y7IRcyn9cx4Xru674tS9
`protect END_PROTECTED
