`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wSV0ZyIeH6MnrLBhGKh9y5UCMG9J3t4I9U88B0NzdER8iCHY3UcuHTmmlCkx8v+9
OJGyvETrCJybyVz0Fe6c3QMFNHly1qadwSMnMzEEn8Q26gCEMgXbR1IP2Ut2++2K
mjKbf8d0ljIdQkBhTgTpLG+bb/dXr8++LUICMEzNUgOZudi4tZhOI0QvwstjRcu4
pk1qkZI8ZBCwdxw1ThUiwowLZ0uD/01eY+X0J+uTApsQzJ5BWiw5IasbGzAMJfyc
zYuVJbJP69v+IpBv52u7hOIzftacVurxeCelPz5m7xa19OTAHiMkM1OxnXKeCox0
K0kdsJESl0azkTwlLgwutfeBa1JWWox+qZEWeijAQfc2DIXROwo4XR4bQVCkByzu
dD7aT5uzQCR+rvJIh+PGRX0lGJK8mzl0mbZMOxySLF6IMfs8u8kdpPt3eNfa2Aey
CMpu4cb2ojWwIKynYXBkgkNpZ4vdtss3LQTAiar0wyKpNBPPcwLsemPyHB8dxd3e
4xaltiXZq3qafWkt+zHx0xySyH4cCuls+aLYdyIdSgx4MoJbYwBkobfIo9DejLaL
VNKWzxo76ejbQ1FdFYzWOT0cn1DEsBuZBpcJInphBVrWx7TRugY3780geFLmW5QB
MKnex/7aVLf+Idx+tOnu5q01/9uE5pi/ApCjBUka4T9MQc3z9iZBFCZPL4tR80Gj
yd+rcSWTRuQRPE29mmPZ9GdH1z+HaeCfr6D078sy+wz9oAsyYoebzkQrI7sjDi4I
Xwhz5g7KzXfcgB8hMoRn6t2fsXNDjOK126lsCKaMEdVR6tZQr6aCEIqjlz3OcRRL
qxQZVQWJTwGc/3ovSxAAxOB98jCxB/A1TTRCjVGf3owCqn53+mTPp6OYX6xT8KHf
X9uX9k1w1qB/JGzq7QAsKd9wXgdmZ8O0qdd+/ih2pOaiDoG74X+KJAofCcO/Mp1l
nZRtZWUpubNgcjDlfyh1bAM/Qh90658Bxp90Xchw0rUAb9oV7OzuZ+5wnz4JZDJC
WPkoOk9RzX7xZioZwMGFps6H8KC0jeQU92dvbp6lEC31x2oC6rMmAgyBW0qMW0LK
ZFEifnIKUaIDRxCvjhqCyQpXp4M6wLR7p8f2dd6Tltg=
`protect END_PROTECTED
