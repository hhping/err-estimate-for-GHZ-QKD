`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lwF2z1Ji3psl6VE+i78bikuhBlTeLBiIjGcFwyzUr7zKSLw1bCPOr+J3PPqIU1kB
PgTtn1WEBiGiywqe+2NFTo1G8rn2/s5ERF1PxABKlLqw/2AtBXM39Kyv/v9gXwjm
TtP2Om+Mmbd3RJpBDnLDLuf9xvI3ooiIdIF7481UAOdzdsFFifL0PJyV+fkslceq
1U9PUU4szJj1fZEuj5BZ+FzPOtss5EhrgT8MrEVmacwws6hPxRRQmLRmhG9H/fBh
0WB12YVyB5FJoiVYSAevAOeNjroSMPELvbuQ0vcNPGritliX81uj25W60u+zuyj9
rx7AfYl/w/X7b7Ecrgj8ssUogQj6qvotMhuWeY5rwJ0JCke78bOpEloURWPwgGE7
ZhlXtb3AQrw2a0SY+hjx44q8nvyMN6HP0mBwR5hRzHkKP4W2rx5Ajn9CCXvAKxKL
DXpdB9N6rWEvhyZHq6mkhTjWWyekTak2qudK04X3DPUpOF4w4nlLdD31cSOrrn2o
Z2L0+YA77xgwBJxaJ0ki4b2UbM+XX7Jd0Ui4yAiPomijBe85y40jQBjwSFXSUwzx
mXxcWbfQxiW2AOQkpGS7XLuc4SQN5kHLlXXjKqQkEsSKmb8MNmepNy/zSnC/Gvwy
6938BAUvOHnD1R1DSo0SLF7VVl9Xcl862Ap64evW4ZEre4g9o5DmcatWtjiPjIAq
5VKFMlN+F+GDzYYDYpSnij+C+HAh+HOBECaAufFJQ8pipIa1+kFueLYQyYZJrZDc
bVXD3ZBzHZG1B6ApcVHDkzpMmW1Y/MiQLoR1LXE1N0xyfvC5vq2sg/pXFcR0/JIP
MwSdK2mvOUFva3BQfiruF5CnIyZTppHJuFvf6pgG8+jX8q3v4Ry/ULGoJAyhCbi+
K8irgHf9jArAl16P5bc6gwxQC5xdxvJYpDMI1gPgWFSWgPIRPLEPD+1xcYi4RbGl
lpdo/9oAnqT6hVnLo8L+TX2v5DBdK0zGc+tXN7pn5R96BX6c7HjBxAjThooEhtDp
lFd42ayd1kzrq6H5bAru8I88eGQWRcXhaKr91jfcwgKF1/3cNDiJS2GNFkTCgwuO
Juws824ZegNsOwH5V94qiBOiRqHj3dSGJanbdY+0Mx8ctZQ5F7mpLwtW8M2rVwCe
c9rIbenIMC2mFvPl+z3MxcXSn5j52tsX9aVfjgJtYO/XX6SL2Or8kIo3ZZ0X1mw7
RmOXtp4cAcdZK6LaFj8e8QYpyi+i6sFcw1e4Gq9Qw7alXzqu8ogZ2D/lB1nMbitU
AvOvCK/1WGfFoybt6lC5j0imf/iiSDe+iayb3/ILPXlfrkKZnFLrKOvEoiM+9klL
S0yti7+e1EIldjCbej2gQwvj97JaofpoA5qOzpj1V5mUSev4J5HlhxQjvgQEMnC8
CfxrzaqwfSstuyGyGAOZhq41hrhJqyU7OfluYNQpzMNpOo9HIzMYL+krx4EhzWqQ
rUdcD5gH9AKCz5no4hI+HwNhmNj1ZpGiWpKfZTBOMHfV0iQ8KoIPAPSTnWZnOcob
0deokYjvtNj2CryGvBCQmyHMGxSlesVDGE5ptjMLFLPkuURVkMg/QA5TSgqKDDqR
rQiX2pFhSeggH207GjU+ymg1OXw4E4HUuCQdAA/XZwgNa2Y/sSuFyCBHbOFsB5dK
+fr2F9/0qZqkOEvCV9wElCC/XXxbH3XqYaFF7yG/x+9KwNantTf2tzOw87OOTGMZ
1bEmBOSkK7hBhlijtR2q4pGTOAPCZIxSSF43f6e+IwZ5ND2vOoMakv7/XUMKAPkr
C7IqvLwA4+XLOrXEN/ZU5dVYeB/Tdmo5zLoNSD9GWGfKnNCj106rWZ8o/X15pOUv
1HR6emh3iBhW9eeF4YCk5xyh43PbcvNvd3YOEK6APXzt70ihsUZR5YuXJH776DvF
G8nXqfi+WUhAGtBS5nGDiiZ1R93kER/kHgwG6wEuYrpHhvKC2ggwJHpLmIgwMa/o
f5RwjIKgi1TvBr17NmWeo25C6JEQstYknnSDP75jRC2lyUPEN+4TXYQAewuxO5BK
T0tVN7EmpSmowF8BwTeStw8Qu29RXpvDxyEteI1wwRJsNOPU1/ihNpy0z4GmMxLe
LP/UMovQmAqsAHdToJrcGN6fnpgO4FYOWFiNIKQIE/F+fp/Op9/NlgZWmkflniIv
Ha2pMMHtQKvJY9PXtlv8WYVSlBGIOu2A1N3t11++6Z2fTW+jZjxPiXwJdmDBmdMD
Jnf5sTlnJQ6o45uTOYwjqLCPgKUBjuPKMDm+q+o1KQi0jNQUQq4ZFaZBQ59+NH8c
19BvvE3VGSsY6WCrc+I5hd5wzcN8IWiMe1aF2+FL0uPFi8OC9Yw3n8KQvUgX8hK0
g0BjGvdhCWwRGGMErGSgxINx0tXmlGeSb4sbf6UIO9CZ1XI6lucDmo545mkWHTQB
90YX9QaGxl766kYPQsOToNvl9oUlTtF/2Ey4tAJ7kPr/wOJaCA25nYixaEVbAz5g
cxAKN10MDYN/AlnJ3fErWFeYklLo1UDu3JF/HddbthK4Jykd0h3n44UJ+upxF2Rs
ZbaXB9ZZyk90yf7Ky0jk/vIjV0dDGa7ZRdRLWY6iKjJSPzzHhnQiD0fszuo/HKJe
5zO2rQ0bT1sN1FRsyY9bAkuuoO0hUMI9q0ful3UlPbxrjmnRm4bbBKXUyFkc39p3
QhHssNORhKQTWlEo4OwxCz2bE4TmWqzVHY2Yi/CUWh577AtjNNlXkqw/LHe7dYcn
eKJNIxrSND+XzxPgR/YrVd/a3g3dze2fSdnMLZz7gsorV+y5wqPuYPYwgJ9B6bKM
b8U1puW7u/f4jQfAmKtS7gmdmgHjMoEgtADcA4gxnVAq95Ve4oJvOdeuQAgArpWD
8ULXEMRiZbwGH79wmr0BvKZSn1kVAxZFQn1nSus9e2VJsk7JPiMLt8WBtGB123Qb
Gt84TYoThjNo0vOImaBFbK3qigW/NRY8v37hccsaSA/SwQlN4rQ3TDUE0reQ44oa
H8oxlNVYfqORPQyPedwsQ0P7dZXHj2qEegCSyDBPq4QEY02Xs13LLAVmEQX9V4Ns
7egVh4o5DdoyJuzRi/jFdRF/yatYb9hJldAGGKLdguagAweCfHsI8j5nD8/34uiW
31CzoAb9MRGCVB001YXO5ArDFhgxOOGqC1JHRAFqEGFQOz6KaerGr75Lm33W653G
y6NsJZ0IXd4R0BQIxwuqOqw6Yhx4MQMCFaWWaH7R/t06uyeJ3IwxR5PmIwDoHD7s
hLJUWVavUaDXrlRYJzRHJ86c+idyoggCQkQ6C+4XdYMUpUq5cQygWfYLmTLtZ+lH
A8sS3wWmDyNh7Nka+C/8MAfoyFSAc3OtNyhpxUxYcqFEmUo5BxekZ6pb9y5tiXFn
zsZCfrixjUeZFKt2Ih0d2pwyY2FFVhBetNn/EQ0Xi/zb09S2Czktv6uNsCMw3GuD
c4SczcC8TMqJfqwkeyA+UbKHo6npwaTK2Rlval99fVimUci2G6zBrljeqX8WnF9M
/rvwatezEkMd8BNqXAb5v+O9pQLCf5fG8n6QAK+fAofLcHuWs7SPQYyLEXYtazri
zpW4l8JTWh7o2oKRjIAwU8r7cGBsWk3AUgXF3OzNC2BaoPpBQ0mAdYsaTYqR+AiG
NdyXi4U1AL/uecMzZueaqMFFjN5JMp4HraAYc3/9sm0kg6cZRFZBZcuwtXxIw5jo
EykKVBZRnOsvWnAtaPPQ5SzW9g46kQ2fzXSwCsHVt6mn0N9lwRNUVNER7kH9Rg+0
1AarW5gIUHMw6DQkMuakIlGSM1tFbO0ey0RVrzJl0sWThzzjcPJvP9PksLhTTxvk
gjuslV9ktKfqrXRgBAZ4OrtMAE4kWkHc8SbbW/qyvySCyqBZxKOgdxavWr009vxB
jkehFHCUFV6VK4bqs/05SOfnDwbgtV7GgnQJPYktZ87geKUy7SeeoPt1GD5z4yic
VPn9YubmbWJr2e247dL1TE0T0P4JyktKMhAzeGxiWsz+zb53KPL4XsivC4OTpzFF
MxxkbuaLvPWmscKdOASKwy/zyt8wfpb0ftsoP3Blg4cMp325p6DcnnSHnlca9AAp
HMIRsllTjaDN7nB38vOaZ2CD2TpNIntR/DHCt/v6ZJKUOPgpb8CwFlvvw9xp49wu
8jK2wrjpA4XfaAYU+aJ/pBSaFlGfp5Yqcj0Sbf3mwkZTfBzuurs0yDY3QJsLPy6L
i6XFA19YRby9yXG4MqFYMUc+CMbR9DxiEgo0QDSEu8NtuQRM3nCzK4aWuWTFq76I
O0CDiiVY1e1++KPQ01MCQ1r35Dmgkhw1WWY5tOBBDAAe6a2yszE+qmvzTI+UWSiF
`protect END_PROTECTED
