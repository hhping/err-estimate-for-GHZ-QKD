`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aBOuekfRn1vk2c21AHXFdRcLutaYcqlhzRM5h3trSRPsCISGCL7wYcW8K+qJo5Ug
OSoKzvDE8w09yq73NEmWGwdvEsJoI+CYMhNtm91uNUrglwP2afb2NJmBZoqTicEY
CAzsI6BtOjgh8eOxUjWBvp4yGEAjYrMMXQNOD82Un1ocWOgxOfB86AII3aknkTQq
9mXyHH8WjT4g9isv5RBEICMRrlMjeX3au6en6OKbEf2U28TatxezH6YGd9modljD
kAj78mznm+NyzzxXix4qZFLznlw3UM3C9xUeE6jgIqzJKboGtdvUOr+7jWXS8TCi
Afy3zO/ieigx9hut2Rc02t5xWvDyEUNKgfSiDGtBTcr0ykotL3/pkq0hmXQjK6rA
rZbUjrayywWF/6BFHJr5oIciptalcaozEGlEOAReghl4bYPa/jx/5JR5UXVAMg54
Kr0E9BrsnP6W6pGwLqnNS+mdN2wtyRT0RfYyCot461uJyShdF/5qtrzwDCjD+v+x
N69sRwtP3vx5O32swfw3Tt5UWH0Axg3B050U8XJ22fDoYVpWSC4UArJXyzkyPdnd
uYWU1mmmldSNEhUCgz6d1DO65dSwYaW/0E01ZODfrqrDLj8Gp4jkBBrTdmMsx1Dk
Edwir2KOzRcUVE+XsOEnP5Nvh8tMUswQeO44lWJ2v+vIhDrnyinywVyewUq+U5Aq
kyby562GYpRx+gvwEYYxJkS8nXUoFlTsEzd4U+hKfb2kdxcjQA/Q0B/GRqvR204p
I64bkmnwX41BlMEV1RRNxvIW2ZzBw39ClsFBhe9m/dzpnB7UB5vCaK7piCQr97eK
79pg+r6Nui/Zj9dTn07nbZMt4QWlxDWa3kG5l0giztGnNPStL8Xg3WZhH7oBjZDD
TAl8MwiV9b2i4hjFrY5/01Qlqx/ixDy7cU5+IzHXHGdaLwHolLrVMgeIgrtohb+0
ccBRTSwDZN8aCO/J+0dTcPlpAY/cV//funuObbNjGY4E7Rrut5hd/d3D1yTKZoaL
moK5XjJDyvkiW/z6yWH/V41aftT4M69UR0gnKlc4Q0WZtD3wgJoAT4GeeOJapN6S
MzzYQaeDoYRk3a79qxL+tZ8z9Uot/CAYAxvP6zPQck75TKo1JrwgUVB4GcPGbGU/
UDCr1lvds1tXm0sNUAs/HcA1OIqAviKJRIgQqSrJ6rGkyMCwFqW0pX9gP5hmmcKR
nP4vzAW4LgGe4t9201UU812Ugie+OpVwBkFK6q4069a4Q29mwZajADqY2/B3Zm79
iFH4gzqKVMaRRD/tDVqT3YtwpW0firO/NDC85LxlXILC2jUK/QYxelq0VpZzxURI
uUmLEbHC9f0b7jXzd2JfdGltaJ4/VyIevmY8jQ3+Ww0D+G+em0aoxmJQNW6Tf6PW
2z0CRXJkmmFJUz5uphLCnH+FZe2GOOUQlWs80ZJy611qWW0rjCCbMIr27wXPUuzm
FaxBBICPSyVSa1bMPTdtZk9GBGzaPzNqElFnn2vaOoYkAOaAAIvJPcTPNkLUNpAq
XNcsAdV3Ld5OFOX52lXpzYXO5zdJ00iVSeKf/v2G0y+rv0ITDczCOjJBrJ9h1+pp
U9uqMANwFHGNqjT3rMHVtQDf9/4lBSRDIkbi3f9Ek67bZWFepHjC+8bi62l9p7BO
sqK0LVpPu4HwAKrUvmU9mHvhE1jzeO6W92BYtKm8NZ7jxmEHcVXIoNu4Pm9S/rHq
FHQXx5kwkUZA+0QCPYerAYQO4yzMkseN/eXrVPM2C8z4IVc02UnsSNYBT2oLV2GI
bV8hTdqTh/kZnj2mzgukJeIkZRDNxdBcsICuSxK12wvIg7g1H6RDb4F4LKL6pAmD
PA67EWcq3vfocmoewtBS0sWtzo0gJesq1+451ciwclFlOemhcHhCAtWXu4DOMGY4
G0JlST/itXm8u6ZxEGU4/yC5kS6XdHMX8/WfB1GETTro/dfwElEo/lBqFjW9VGhk
zNFL+DBH1DHgH2JseSSvPMxInLp4RzxV/1WGJ2ph6FK+mVK8XxESHHY6h2AMvGqf
dQBMUmgMr5x8bn0pUimuY3B4F0m/8+2MAnaX81p2pckoGc4I5162fOKoIms1vmpo
nMYnsQSELdrzxj5nbpGDUTUi0rkhwuAb+k0J5zzgNRuwUIQg1KxhAyHckTIYVE5n
+TcUB/TYmRoSWVXwd7QgRJMtLTHBQcCLflFSgt9cCxTbgZhd6Ni76Epp0DxVE2++
39pv87kQNUr/O1azaI0W37PQ3+rHnea2fQUC5DjCv27xk0xy6VOJ/4ct6ozgDO3/
iiZKo/9p0SbhocpK2qhcka6Id+Nh4FOFFi/n+WzTH/1u1vlCrWgQhuiWGMCjcCTO
OejUK1q0tNj4dg8WwrRqJ2D1R279qSfvZVlC8oMdPN5UQ6q7adIxg7R3W5ox8ojt
MBp3ISLnGTSifhOHisrsC5pCnoqsRXJ5OG2Z/eH0zYixmz43/DIZAIn7qNIhRhPv
B7yvytCAqFSulb9HZ6t7wAsKnBAYRh/KWa6qUKGTsi+PT9QwNdmpxhGbbQjlmOiW
+3nypv7WJbDHXYWSXJEQz0VA0+8ACWuJeKw56fIVOk5JQgRkbJkHtgB7yEsm6yMC
tTrpa4IVncU6ZRf1XoxE1vl+DLTzCRV+GKHvUdfasgTylN1JZ/HgTnIdq0PmCfNb
NW8iiRFXhbaxoIWcri3ByCLCD7woVg6PwjHOg6ku1tB+9r2jOUXag2KPr+ExtnEF
4eGO6ZrcF1gvBOyyGPf0YHZrM2XfalR7mZIpovsLfGWztUhuQ9j/NVDBFpqEzf3E
ezhruTPxEGmPjUsYeJE8ldyEFcYdigs4OzRgvx1PNY+0bKJFQrPwvlvwARbJmwR/
wuWv+v8PgNsiNf546f3GV06kcwtthoLTi58R1VwfXmswiCcIrlBSrH9xkAjXM3Uc
63LkhQyWhDwENpJ5G9jnumNklsYIJv8/vBN+UWL6KCqgVwFT8a0067IkPA6Obdb8
vY08nXlwHequKUv0wQSDCCF7el/9awNJ3jfHnaFbtvALLU8W8yH4EOWgu7+W8QJB
s8HI8vod8BXOGv6JefVI9x6QcWSPr9ORpUkp6IZeNjRqx8bd4jQPJW0qXX5X1l6s
+lchK21Yid5XpMr0wEDcTKUHScj6kMMx235lBCcGXBN6Wg8uyq9N6EFU3QxzIFcP
UnosHzOw7ga0OiGocTdyMNHmJJWukIVJ+rrf2m/esCe77yvAzjpEFROX01rXOwfa
5tdwnLoLXF/KhF9eudiVJ8fHi6tsY+qRJRMFnlyiVKZxSXFlknmNTknCaj0TbklY
vnpm5ciiTSy9vyR74mD71m9rjtMRTHJBO3QrcBVQt++bg8S++zujBsqKfgJQatzl
6canDO61dE5vq9fEHZMWEUGPwGYz06o/MhoAStWGEFqNJDbaL4YUD/b064F6tquY
6b2qwo7EpeS3wXU4V2+Y8moThT62z35I7eWo5+RgBeoYABGU5Jj1hSXV2Jjw5S9z
+O/XG0+o+flqJGJuIGxWAtKjN2oow92YiojZG5QYbLnUcY1e8gIc4QRKswdYWHc2
Xc68iMskKhRq4Gj4n99qzA9FbLWd3+PL+WPgkV5+nga+GVdKLdoH3+q01tx7QkF4
4XhejNAAgyLfSmMSbOC3/VNH9dOWphHR6223PJr9LejZgVwo2uftTM+GrDKxZ+e2
6RQ/snZxhiyxNhzdLc1cyWh/yPH5zalL4iVRhdbbvSafzyz5EZyZ2vPJT2fUlvAT
kKCtzzV9BooSaCrGbh39wjMVZaXLMN5O0R5cr9S+3GD6xgbX7SsXi+yJMeZB7mcM
uaGx2P/h9/5VcQ6OHbRGGA4dye/0XV3A+dNYW3bzRmQyGTygZKWv7c1N4UH43/I+
z0bTuE9kWZGgngoPsL1NTg6fJ+ghTtCteTbcIjBl6q31doskXdR7bjsYfbfBTjVc
rFt2ByPn+MaayvQGEs3EQ/ros3K2hrwaLaUsPJj8znBlxX2OpCD2zCVaa898Rw2H
pNZo/t8llumt0B7SEtGT4NkdrEU7VQ+0e8lmozOQs2MGKnLGjSrwXag4SESpYPy0
oo4stzWC7ncKwezSl2eH6Vt60clOgZLBZE9O2MeJ6OZKB7FxTs1kveCeArttnYfB
ocZfoen0W+5mxBumRYsRYiDbHQmYwOOv38pdwCpJ2M+vJNHQ9qi1z6z1KEa/uUqB
5Kn/JZ+Ie4AyGOd87sW8Wfi1LEfQCutLS+6pzEAtrg0yQzqgmWI67FerdY2cZxhK
pT957Q1Vh7Nj2rJRdl6R/kha6J6tpipak4Lp78mGjiR448WRP1uCZfzxoE1nE57y
RRCeVnlfHms0EtNU6cq3gcd3GHZE9es2X4W0yd3DU6GVFKBdALvFqwAoAVLc03P/
Q61DmXVJ4wgkhHURy89hWRNj5CqnwCxEyofCmSTZm4nc4qDXuAMrZvdbrWhifjVJ
YQ5WOmbDuW3iIIHLH02nQl5BVhxWD1cwru64pk8/A8B1KzcAyfOGJgXepqJKoKCK
MpwwkMsghtHdtbLM4ZBikTrGh6G1FFAfywNKKjs54F9hNeI3FMXsl2Ih1G8+g2hQ
qne0SMwIjl07gO/pchbo7Bf0eFjPhehF1+QMhlWezDuCdm2P9Sqtj/YwTgILXahz
j6I/Eh8l9p/SgGBDvkAEbNKqzmvixEZL4wsDTwiexenBlU+ZjZy6DUa/B0lNp5m5
juVrClKlcdR4SpRcV0+OWUhWiMRKZwWe/4e6XtmiH+IM8VWL7ybMYMR+9r7+67RO
3jbkkciJsjA8ZIAIYMd3zOJt/B6h9deDDtngtYe75RRVksEfhvjF6R1iLvF5+DP/
jXxwP7CbIrWk2gAnojRwVgH8wanElQCzbOHugDDl5iqSAgvje/ZdKeJryAnyI/EQ
HQOx+kcZF/7tkNum1zjgW8CKo1RDcTEh6GfqtBrZKruQPpnLvgugdlsfV7IKS879
vipMiHNaOXMV2ZfHCYf9HnVlvaItiufG9ZqizrMquGFVpBAK0HYb8jfMO8fCK4Bq
Vp6Uc8cjQFTdxeevkl/Assq8OTkVPvWVlpUhZcbpDJxTBMu2ojltwqOvPKMklE2C
VVMI/kcczn2Z+fi0SdyvU8MT+uLZx5GRNpFMCAW1TSUTBSPa7Apyd2oEy4cOOekq
G8JlpjH9H2gfwHRzeaAnC1gEwn/KSjBhb+Q0Lh+tKf0gFyd5Kse+iiRgkJeITL5r
yskFDMA8XbIRbNnnvkYEpIKxkwD9sXPV9kKAYe+qy4NZBZWokHJx0+/+pAbFAce8
ni61kWdi5clrKAuv8w6x6W7Z+WJbBFXJsd/ZczKYyvQgMUEM1mDHYj9x8dQ5zddQ
oxC0N7xcU/UGfv0u7uu6U/IUdKrpwkvv+4SoTkxpcfPwC4swvI3cGOSIGAXnQcNC
uOvzfWSiXwiQCk0pQVkJxqL4sfCgNpLuFmMhPrw+csogjZpJ14WJYhW6f8Pkrd4C
4XoiGOlsIziJAIPpusK/AkCNNBHk9Pycn6FM8lFaNdNzgq0M9CSGm9caURkNwweK
6PZVGxDu3W64ImgtwBKCeQR/5DSipnSxkmpb9bz2gTy7kVQRwo5IV6+4vUt2fbez
o/rKlKo/hN4j6xv7737hu6WeBtk16i5kimXqTiWVW5IxHCfv7xMMppXzjc2eASYh
6cGWTQVf8qStN5WY4D7WHqdp4qsxtCYfVO+hdn42TmGb2QBJKUEqUEFqp8noIt1y
RKcl8584NHnULSHpi2Z9vHWK9yKYqgdFfFSltB+d6jF3ULQFcoiYH/w2ME5ZTf7n
P1W3ilChn6sW8z02FF+Xa3WH0qdp01LvmAAYcSRV7E8ujrkQNlHwoerQxscUTVB3
4ankIxJzVB/WxjZFSBfDg22S3F1WirPAEiMifxcLztOCq2fz70jWv4P9RqK/pz4n
3Iprc8tOt5FMIQYXNye4LozRKX0O7V5EL3v7i96QC+AwCRMxqPiB4wNk1LEsBLN1
8Vjihj6ohh80l1Vw8y0MUbLsz7rvA+bjAdue0Gp4BOKHGR+QzEeleH8T4Tl8Kypo
72IpVclUSM9AK2Fn/buAhy628UOucFMuFyBW1xqpGQpJ/h+rAKM7Js3cjTk9qYEe
m+liaNI0MK8E32f2KjEYQMcoRlVfowz+pTrdshr2ubTJB6TTaIM8YRtsPNR12Tzf
FVEkWuI91azJejIkVPVyqIK81QtHae4FUbGVA36GxGDLQkjI7/jsotrHkJJvYS+Q
kVW1jzea+6AI8vrv1/7H+aA94GYAbCrP8tayygQybEg5arslyjKQA8YOJQUwqY9u
OHLysdxEFmG/+4QWgYELSOalgvomEdwjbiNkA0OU2bCUy6lZwQmrysLteFwG7T9S
mjbaXNxnGuscEHP7BVZ92ud9+y3aTeIgygi7udEpfZ3gD+F2II/STl59w5BsC5cK
T+Mkv73qwaLKqYRAZ8kvh40veeBImTZqaw7Z8TgtNABgyTdNplmnhi+kJYYQ7yV9
aypzwlJSkvydwHyviVQOwAqOMYqId/93EUDmHlbRDzemia0n7p5sqAdgOJJCM1w4
Cml9jyjSVLp8R7L0gov+foBTYU3yGyE9DEJ8unnePm8rQ+UA9MhmZgO8QETjgojS
T2mUhoZJZE5CVKvQzJkRsXXbdSJchYnOBfV2SoQ+Q4Hf+gA0fH4+IwedAmgh+ZIc
W6wu3G0beqg/Xf5Z/p63TsGrkOoy5+4xczF35EoCLmuOHMIJu4qdns8TNlLBbZnF
xLBMlXgq11gC3tWjJlFzJZHNPcDuFFPkgZiUA6FsHzvnOLwuDj+wY+VtRYQcpfwW
+PTstboJUisspu9wSCLzRoeeqCFY5mSAR0UtvxcxdS5dkEEUR4NVqL3BRCuc9kBm
ANpCZ3dwjHSr1OSwDFqQxluFPOntii6tpkjCJWOGQo05ev7XxOeWPEwWqZfKrF+c
G15KXD8IyFKlFY/n5eg44H6KHiCfCHWRaCiBRNspCVw8cx/+WLVIoS2m9pXy1NOm
Wp7sg8w+u0INApW0i1g5AuhOGlcTa84hRxmSK1i0bw7d9mrUCTwSHFANboKX9aj7
nOW6GCKzEO29I4v7p0KV54f125T/xiDFAyUxx87YGsIVPfhursD5xabjQ4xWj2Sw
uF3aQUSZW84FJGGeQgmLTWYJXWFQY7VWvuLa08f6otrJVRuE62jkzpZ9V1H5YvE/
+N7n0e+BoqPNG9OiXNSQbICZKP6Adliw9ko7nlf1vgmEn1Rd6RO20tMEFJAx8KYf
eeY5jhJfY2OcpLzfYl9q1L6QHlk7fk88/ZiKXd0hm3lzKLLDuNRN1Rr/YLYCnjkp
n50ipD76dJrI9jgqWfMnlaucUylSOOQBc+f5BLPd4PFyQ514KpIc+XKA7Ta11Uat
Yrjtl1tOsZUX3zRhWebBtRklTEE7pyy0n+qY2W4knZvt5nF/5cVuc0vkvucURjyN
AVx9TFrNc+/dJz1R2CILqxLIgP1JcxsjyjVa20c0/uCxluJbMoI7/Mavo3CpUOUy
g1K00ACaAPkOPGnk+g9k/22ZgYQteBEwWO7oWJSNgGvcQ/+x7bSzFAecjFYPWCIi
ZmexCVulgejeLZRa6e6YwtQit9aPIF4/sQhaO0hOatmCoqjDa2QaA3+zZxpGrRCQ
EWYSef9OmFkNmWIVJKhnLXLIjHinoYBgFuZCxGnYXy1MukdWvC7kfIHxAwjkNliV
E/2KiosOZ405JNNbKIRPGYRDNI/tf3SYc2ObNZz5Y69UsIX24EfxwRi+WW0hkYeZ
p6kAuWfS+XQyVK2iugoUxWspzQjxtRfW41eL//vtAKk2Eor2oOeACrU3QvypFji0
7g9yXhfULslsjkCUOLRon6CTtySD79kPELZFw7jl42vY9wSFfdEw3X69ZIrs3R0R
XmjMXltmDqkKzbW3r+6ZLcU+FYOsIJNi74zFuwS5mLAVq6hIUmZO7qLgL02vRJhe
Ywu4WFGer69WIth23QiVuXKQw2bYlk02x9LhkCobW/JkUvdwtY5pODnF7gCjGZO2
SC6KrKnbjc+Jzxdo0Fya+WgY4iSwFHzmTWwhanBm883sNr36bJT4W5Ib9AV2p+97
npvPK3yp8Ptu16IFHjBTgjBCuIhtQFoXuSPnKMpQE0qT4k1lPv8KBL52gossxS45
W/WkAh8+/aKM0xJq1NKiSzvUOLV/fO/m2ZERs1ZbWxQsh6CEOMkcujT26UOQt8ID
9IpUq6ispQZCBWKzASPC3py2U+O1DM0W1CNsPBKINEoVWS+J2aRelcXBMcQXZlSN
brnSdIJSiUZeCoRwMszwseIv0Dsdez12rApNrpK9EhIPoSxQSXVXX/yKBTM2ae7s
zo60xqUacErYMd6pv1rs+2fXqUErLTnKfGZtAfiKeq5mTUdney0ST8F4suFi/lTN
jUD5xBmusV//mYrtL+5fGpfqFXY+16IYRwX5HBLX2sAGERuiQ3bFiW4GPl6xfWkr
CyhBQxMTKw1cbREN80HSy+kvbnINd4PqwAs+loidIXFLclMuCvDg5goQBXOk2Mfb
uEnXeG78Ic0flGZCFIlOvFOcAR1qmWwPSr7VIoWJG7S8Jt7p8E31SAoxPEVzj5G0
xvKiQChErpV1lVJSDkMS+RsZSTnBYQ5ioaTLohpNei9kqAlatdZn/VTdFc+MbUWd
lOUGdYZsfhVTwF0Jt/VfWhFYm56xQTKJic5G1GNVuTR+u4pkfZk71YBujb/9dMhH
Hj9z8r6pibZe42E1kARorp6TgOWpZDYrtQ2rbdyfkPYgVdYeCubwcTxZot1Tg/1v
UdtS/Hb2T6kmj3/a4hxz3N8RvOUdNpSwhoQTIJSHA0cdVgNxTyW/KlSwRkIGpMob
DZJ8tf+NS1EXwXzjSALB3/mqkKFc1mf9xJm5zfFcrS91OsMRLNpomKiQj8w6lrVI
+55o/d0fZYnWcw7TYdi4GHodLLX+vA9QZFS1WGgw6jel/sip20FjMvrIk7neWwpM
HcsFb0T68R2ugg+IJ7Rwt/VfSa/ByVcB1uM5/N37x8LMLwlckFXcz0BH+4MRocki
3l3ngAiVX/L3Ay2m5DbpyxKSbtYJ8bR8kbupqL2tCuGzou+snYDuNbHuDy39Mn4x
u/FyY4xAOl/tLCh9e0cNi6p/IGfAH7ZKR9eYEpZBZbc6H+vuenCXCI2ZCHQd03mZ
ePnNlx3fwgOMvFDbRpT0my6T3jFfxeBlK2J4z2QfAKUh/3BAS6ZS3Eoe+MM78efZ
dCafst8blEqSDSpGePDBXpYS7jznIJPO1d9q/s3AOuTaSsmuVBupHXF3EW65WEZf
TnUoCprGclQWVXGhA+5lgCrWfeFFOyTKNOaIEYBhEVwgXC4m5q6K23weL/Ba6MJN
L1+HVJWHz/WlCSV2dvOHTPMAgz7Jvwib1ZCLfv7lU46Sb+X2w59xeYvami2wiLh/
MlDC+VS0v/HHcp9W7sbB9YABAS2hEyQjvve6rYYcvuU4o/FcSX58qpdOrRD1hRpB
d1F7Z8TRWtNr3M8mFVPtI/dktpwlxTGCe3LohlQfBRAEINgjTcS+OWRfjdT5hHxC
9Dn0mYh6df/69kj3s/zvscEcdXMQVuky1sfCPRcr/Mv6Iuxg8h7HIJRGg57JmHMg
K9yQhqiLoZjVXIrbYFg7Rd969479I3EvXuutS/xXKDeF6YdVKK2vGhKJsaTGb7c5
TakE7jKDJ2ZcuU8J9RhrubQL918A0R6puyTRnRtYahedjdqcb+WQVS0owOaKa3PK
Wju6a893i6HkrcIWAUmHfVsUo7B0OOCUVSuZogmlZcGIzOuV1Vy6vI/Zd3ppawHC
dKPFtE6cZmehcTBJwfghp1cV0hyvmh+SFtgtNIVfPdn4tOSkoWdzeFQeWrJvrYWG
Y1gFQky2PtAbPPJEux/Ci4Ijk8wUiDYdkmECCtg6k5BXknkJE1p3K0+bI5DPiXhK
Xo/qSjdua2tXBmjTBUf0Afanj/AfNHj/NG0dz6vLCjOJBoaT04yf3/w5SOtUFgwS
bqMIQIW5sEI7Frp9OrCVxX1cop6fT/gGnHh/yZ7XaIaai6a8Fb7miSbCKbjMtvF5
hdh6aApXjo1T0Xi/PVM2KGUWHRtBpOOeqH0xZvhZertvI/ewa9xoEM/sWRYF6WvW
4gKAE6/DOhGDEMrqB/jcV6K3vfq2JftVMTWjnq4ysNp08EKMHss9EtjmKDvUg1AO
1KBis2pkqdYuE7oEa8WjjXd9B2i7EohGd1rkkCvH9a0=
`protect END_PROTECTED
