`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mbS1eVeg2VTdSe/xxL/OaDgsVMn7wRZt/Xu39bjPUlDxn+T+qixihePacC1/tUMt
/Iw4vZw12g/aP3uxRUGrxyoGctHNstJZ15BaB3qzYYReXduVL0+lJ9ehc/iy5Ew3
2AHJIuIx/8/brWavNUdcYv2dxptTY2oszYif02ayRv707lvM1RlsRvY6x0uvxA8C
cClVah/GOfYpoQMZ4oApjIQoVosPUG2Bdcv06b2yG7jf1oSb+ypj1D6mYC7Vh0+D
laSGO2Stk4epwuJHiU7R7uO4NkpYxMUV900K1abQIXFIdxiitC/hsCgerEJh1ckj
XfzyJddDF8zHYu5GLcJ3r6wZrhg+cfk1/dLHfKoUvmfWnF/EGR0I3P183IzlwO6B
qwm1YzwgECsJk8nzPEudYxQkSuF1bobXvFJFCxNScEgvTiy7eKBTixGR7rHFfsQ1
0edTmiMqavQ+t8301UEBM0J3hxhrYAvMigzK/zhQ4iPS+HgBkemFJA8jiNy5scOd
MX2BEJigQmd1l4BNPXjBXMbJLepXAtWYCJUCQKQsKdDSqHd2pme4zjDa/9AXzw+T
0wu60uA97ZG854cQF4rv0W/alUGiI2OUOf9kzlagc/hhDT90TWFSbTiSCJF7tqP/
PpD3MgD5cEi9nWATtF9qkwB6TSSpCT7ShQzC2wpXo8jPu2kZYtpG39zfkSz1gy0F
y52bUvbWJBSsVjmI/OStZRQtrMm3zirVwrh9O/na8deeW+A5ljDimeNOyFSNR9+I
VpUJ5zIULzUVtr+ixHZ4yxYRQmjJjrk/OWlrN6GHVi1elAMpByxlp8pycVOi84+b
hiQ0afNiCnLZrWOy+6p9uUlIM7hGrHACBs+pFormJALY7EJHIJDZEVhyffSM4vVF
ehDqvfgzVJzMzXep3tBIrqSzNjVJjWgOHRCdfylU032KCJzrEAklQz+l1g0vHdh9
Ma7Gun40bD4wHmrcMSUTCeItCXtU9GKvG617VYlNyrOPbiU/pUHtr61/6XQMff4f
q2T8d5RFiAplys8DEc6ovOMINMWCpkDu+ths4oe0crturEdvuAdTn3znmLHSelYn
fyDiXuCWubkI3b+l9Lwm3yFp9ngL2KlugsgWE914noN/fxbq6LAbgTdl651XWtoD
O4jvnAKfMd9Lzqcds2xJV8gPk1xt1p+utef4E5CZjh4XPic+XHM1QoOIekADMQLF
xc+sYPA8DjoHB2UC1z2Csvm+KFfVjdkaIbWmSO5eLkcilvVYtv5vHVzF9j7+BFhQ
p7gSy/pLfhkPEpA2wwbN6/1KjTs+pHU72IeFAYyD1w2h10+NAu0HpkuNNUZe1FuI
Lq8S5EMM2G/UUvCjMxVnHBOjmaSElvo3dwjqtt3b8I0r2WdnkN8vZEg/zWDKMG0m
6TEt4UQfnRAG5iDGwcrsmgTNcTl/4ziGsx3zMZ0wx93sRyzFs9nMNmUY1urelkt0
VOoxaPEJ/39amicBdFRY/zzKKM5CqZonrPDjppHGpGOkiKtU2VzoOjBMzzvIV53y
gXBv0H+WeLudeonEsyzzjRhcAFCiCXrsCWWWnbV9NOozKbc9GixYHoqilocE36y/
Cc1Gn+nbnzHoV8d697JTGV87eY6ghWLKafEAOGfrD74AUBfo6JYMZSE/eQA3+9sW
WwuU8VHQ9IJO1iDIgu6wabGasNKgvuOX/FKlgkMCtHeJlnrKP6k1k6Pfqzf12bcy
zKRaWwgOqRO0/l3xjQYwL+GgE+yv32uKEvBh9LvMIXoIuKVqwX7iaGaPZKOPohfy
ctUD3O+4WoS2B7ty8Nj4518kgGL//HlpKaMLvbU8OwLBLfSECQDl36KPm+4igtr0
0A6RGrgeEY+oOC/+a0Ithb0DlzNCw/5fBhmIs+LYxG2W77B2pBTKOVqd/Z3kH1rY
BAgCV+gipLzAkaqsuDhY3VI9SDOlPMCCVj4iJP54bZtgSjeIsyskw8KiJoPyOVXx
8hZzZtLYPEaSYuHbgvnNTDI5VcgvXxYZklQALJ9ZhG0f/EC+gC3pOWLkiJHEucSU
FucEbul27TYe1FFoDBt2H8ThMNQHUD33BxKQL4CrvHzG5K34TOoCjyCbHFYIM/zn
WhSyytGQcQYKnOARVUBe9QzPcTqN9hEotqDBX+cX8mOTIOHJeRoH9LaUsMWgWAnN
PCnj3GEaWxpK9btu2BqlZm60Luw7p1ekYbpOEr45CbnQ+SzYkcV3GcoGiNhvQ6Eu
zblNibLVOM1HPIFUKEHW3Q==
`protect END_PROTECTED
