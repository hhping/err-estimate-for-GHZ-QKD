`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hXEZCmeK/n4oQlQWdjB/KRLkgaNdu4xDgJQpBbNG90F2GYMBSwsX2yPX3lY1MoKD
dlF9Ugu7zlqEmbDY8/WPyKqGgbvnUvhyMmYysmKaRR31P4lec0yU/HvYcZoEH5Mw
b4odNUxGvVzgrhHtjU0vo51Ai5i96A14OFaVbMh4MVDd+IbuISGuPv27SFjYH0mh
5UX19YGYvoOisWb73AA4A5UD1lwtd6JHHAAVngpOfcjMLgGP0ZziHkA/ZPJ75Fcb
sxZgPCpzMJyO5xtekITCMcstG9+hbXZr/dKsQzrm+vNf6k4+vDrL5ojKGnrNSh+r
S3l7CAnMmGqSBvcFZ1sZuf3ICcobO8iLLJ6/PQpLOTD9iObJILP89nCRmaiIYh2t
e6FvNWdHA3ah4QP5t/yviDFmAVrIY4fiT52KEoYfkmDGOmWOfu+Q0NxsPOx2hLmE
ic66tvoUtjnAjYrroXuURt/5KBH4yXYCiV+CJD8mlRTVHTdd+4QRh3CxyF6rivPE
fQ+AUVYx8boXVLwyDa2mxbDfz2VF8XnUaNxa0nf+3XA=
`protect END_PROTECTED
