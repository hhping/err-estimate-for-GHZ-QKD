`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vmz0AHue5NV6avYq/uP1bDza3Uvc610YmvaU2zt+mTfhtYID+fTGAvtPhBxRue7m
dgsRCqQhDg8yj6snOcqARR5oT0ed54RXw1Yo/GCfFh25mgShLX1DrJKipR89s7mb
kW6NquyqNuEvmlpnr5EYn8rDsGEubnS5VNIP41zPKblReXaKDQqlC1Haf14KNWhI
nWuiVHrGuseyLihrAckGuUdLQ8yTU0hJPPCGuupWW+Ws0MtkuFUNlb5ZFoYeghQX
y9B9TkMN7KLYSEIY0bBhHRRt80LqqTEK+Mb4Jax6HBZ87/u0M6AB1eFyqtHKQJ4J
24X3ywc7LlF42m1l2rJR7GsLC9UQn5+eIyXRJml3hw82BZv166RO9bneAXpBxYsJ
USzJhG2y7jq+cQGzFMlki9ROEfK54h1tis/HEpUFxzdMGN5y3mrR6dwZBhHNW+b9
e1/T2c1mfjgM1LTULLeE/PVNYr/1vq8Q35XgRjYVnfbk97XW+0LfbJDVMq6msUfr
giwLsmOTCymV3cmfb2QYm2BO/gP1LrYrHCjP0f2TWrlTCDnpjhtnMQEBieEFy187
gnuXPqW8EBaxL6Ekc4wadJfhp53opMmI11OAWe9ZSIYJZki3FOqGfozzYlwck0B5
68HGDTCotAQQy4jh2pNsXdnWWtL1IcR+J17/bXUg1y+tOc706CNYpkpl5Ha15+kd
8lh/zpTgb4i+gtaZ3ijbZZVwsp1d318DH6NWaUJqkzdGGo2VrstOS2JUA4suoy56
/H9XJKl9znWF/x50Zzfhy/Lq8Gq/kM4Dw72ZUeopyqC8pOUWUkGi8NKFnkmBd5L+
ed7nZ+Akcr6H3QyW3nev9BpR/oynzy7EoU1tfKQh+memMeYBVFxj+WBbm6YOdEus
Ujfx+yFb3OhQMz0LZwlcZ+IA6feT8s5EwtK1+l8KxDniCkLa8rMzT++1AyCyvL/l
MCLiNQqAQBW+6DeDsPUBwbCr16+ep0UKULWZBZl2DT9JbCTq7o8F9vOH/uhTv4w/
SszbMA7HAg+bWK9j596brFE4jZAnsvjCafyWtVHXWJCC3bieZyKTNvDBfQenZzL5
KVYBLQOY+FSDPEfho4T4e1u00O8P/Solr5kGI2u5sSZDa0woG+Tfn6lr/LnMX/bd
4XMotxcdIr2twR1pDS4/uF/uAI8xup9tFxjbIQEeklfbJbMYeA2KP5fTQnWS3XLy
WO6CwJwVZPX/J69wo+E0qfsH4wbMMf98bqTj+MQSGZL050RTJU83+flPjzUsal4g
E6YenPiLLXBdtMX7wq15qRZxgXoigw2XOTK1orxM010vTip4rsODulqcuFhnRYT4
yJXIgz8HGIn4p8sF7HNrTT7gsw39u9u8aNMtIXWnrbQABCpO1F2I0Fimf2qO3Lj7
iTIsAbjAfC0VFYicquVQVRtHnrTcgkIXG7eMCQC3zGnBcQv3gSDYRs9QbseaeUxp
j0gDr4ZON1zdhEYnLvWWsGm1AiX51Gn/8Bn5OjlypCBGBwdsEMu2xkWwfLVGoJSk
fe9bNTCNLHdjEYJvBJ7CnvzCtzxbxPoX9FlSgoLiug4bH4MGPxbDeV30UYVdaW8i
gSfGIIFMwPJhgBoOzq/HnjR7VJGqng+RHhzA4AXAN8QM+xzcZi9HyU2EqCQ9FZPq
wMP32J6u33GK6Ff/UXVR6KwOWULEquA3dQ1PBcS746hozOB3qhnGdP3uNzUWXpWa
FF02cW9yJoYY+xBj93wfsqkWdxHerKcirwB12igXTUrjiUEYecLTON4DJFDaiNmI
YVLGA8WYkjyFcn7o6IzkW1HsExwXqk8El7gO30kc7u8VcKGTUCEg7SooHio3MD3V
L3S4fCnmnbV4rU9+IA2d4dtxI6Y18YUl93DbGQogPvWCYL94YJ66ayR6SckERzxk
dZOJ3iiiG7FBVia+gySFdKbtylQNs06f+wqB5oZqxNrnkyBuL4U8y2EA+yb4BsUX
2aPM+YOLc7NSZNMlGeh18UZJoVY0SJQC3/Ffe2liEo4v8mMb+Z7hHDcRrceLcBfl
xZteYldltRSgcTqxptyZ9SQSPuSXSlvpFbT8ivGgGkqeUdtMrbpVTCW60kYADPfz
iSz+bJkL3JIGDi01y4aywTuMAJGdTwU8h+rUHg0iskbiCJgb7CHxKoYXpz190y+J
S2pHDmQsatmBmh5xhQMCYnX0IgSN9kN9UKVWP+LepNnKVwCLL6Bi9x9mZkN9Jgrn
sjq6hdpo+FAWQv3RDDE4pPlsjO0dP8m0lSWUOjgBxI+CkgQrflZLykuZd2X92txy
ZsUcOSxXWNR0JutgbKM35zevwjY2j4qAkzXqZTZua/5mI0wafTOycO3qH/8MlGXQ
aTraformQOsJ2ULogJ+ixXZB6GDO7pjwxG40wTtMJM3RAH4k3mPCHgLjrVyUzBcQ
Hx/NXygQuMNtju7m57/Pnh3wf02dVf5hWIBVkS6yO8usET9FK47kF0HbtgFIClP6
I3skO+IJdAWqLDGNY/RpF7H4AgwM8I8YaedHe0azr5LJZrtyYln0l76qixzifKg/
xtD0z6djnXqfEGUbGtHUOhIbavvzo6MZ7Jr3n2Sr7jibwExh3qXAZdLZ8+FIeLLE
5kS1+Ecz0JifSwOSAa1OpbnDW0IMegTl6QApHD4ktbuqULILxawrIk/Q3FvcM1MP
hDTnB2ktUUO6xoWMDpmrNHhMSGiL6yx7qBUEeWtXj1Rmy5GFevi8O6A5JZ1e2yOr
gsiEzKMz1Hy7u4JQY94lmy5tnLD/KDGRl0JT1oqLgW4oXilo8dYfusB5v63lbrGL
xZ623yJoLNBYTWMP+11k04OErpqaK681GOxIDo/8wfazhSmPwaib40hEKiR3bvIJ
BVb77/z8/pswPxz0EsFM7MjqmsK7NOhvUliBHNMxg3NfIfQvwrChsEn72quz/5fN
aRFs0PD/9y0QnXESo4OQcNW+VA5Ztu3PbstlPIvMgzy7TenTBS7IcUUJH4F8EeZa
m46M5i9QLsVXbq2F7uBFtV3LXxIXwUCesmZf9zTnaOI/vn0y/m4YrwzZFMLdOjLf
jXlKwWmJO9HtlGzD9cBiguvrauq2iKmzIOjir2XN5qWrMMbOYrKF8ApZb26oNF3g
ueujRfJ8gWiisRUz/3c73eZqbq7Q6E+jAH0TYMr2b5W8BJ6hG7ADPF6i/SaWw+6D
itsPiyZyNwrAJELGGoqPhjgFJqWLC6o+8M4+WyAsqaviWHlqKV/8l59hOGcnD6ER
PpC84AbIz6tlNksqox5P4v3V8xOPCu4Ix03zxoAIZmi9uKmPa9HIhnvsdJ0i/S/9
WkyuwzLwustllKkddSfbcE4RFNlG8JAKMCpeSpvL7VcMjk3lCBhSag+WgTpXI5je
rr+q1XRXcjJ/DyAmbqvdnwPWRbyr2JnR1VEBS7mZTk94QlZADb57ZKKqPmu6vLx/
mp2DRqN7VGC7iigNym6plxEs/axETjpYF4aE++0PMD/a8KdWSDuFUz/eYsarfgrh
7BX31e/4N5ajXmVyn8tXgg==
`protect END_PROTECTED
