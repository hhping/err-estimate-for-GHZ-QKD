`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6bwANGo+XDWPe6G0TV4MhZ2Sof3znCmNgnvyVfYwAypLjZT8ATNd23aZj6SaNR1i
9MYY1A9MUkQXjtBlkQZ07yJv6BS4X6cHFJAjjttmrVIZOvimnutOQ4T06rFByaSd
4VcDmstf1EmcpL55JBBxwKLELPmM3DBridZlSyS82MjGT5LCjKDKhpGfZSkVLCs5
o5ciMdl0n4wMagygrxIpfntI5yBqjm4eALlY6DRwkRCtAucFu89J+IrobK4z10xz
iApfo7YMdPBULsMGmRDItAUL14dKXKn/AoIyxFqGKBVmtGIbjvjCb7H97+VtNR7p
6Bdo05ja8w1Nf6wB68zZCMGkCLAFlp4oXzBbQi+9qUPDFaBYtN6QqUVyM+IrHumV
hPzWj3JH1PsyIOGk1jrY6rGaepWyVQTaD3rX4KgDZ3mIIi31bFQj/iCZ+JS8u9BX
`protect END_PROTECTED
