`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1+lvmWZlJB1oo6RqP3JGpnChf9rHRVy1s5pUoibUmM/J1YxRApBhvSNfU+cagOVf
iaj3A1a7ZbM75VSk0yOBiv+nQxP1oTiwCFey5xLNJK4nZJomtXdAxBHwIPRau9l2
dH4pmLX7iqGjbkxYVjkraLot3En5/8EbjjaMpf5OnbQ6ikamJxIHm3z8uKG2LAje
J0/SyBNNUdER4lrhDQf/NZCOOgIEnV9K1I4KHAwlpRXCVCfnxL1RR4dzzp5ced/E
Nz2Df+Nlz9cvFlWcbHqoBVjWg/sEYRtsKuJxZYlEpclsGQrEjGFlzUlR/58XwUSj
vRCnISxnvIM3l6n01JCJc6nj9eJj02kRW+BrAgWolaDFoRjM6E+TC8UIzcP6OYTI
X8Te0vPQr6yLhVPJ6CeuVt6K5SPSf5vR9iOAPw/E3I39FwOnX6+dX09WOeHRGrwD
kkP5DKHWtMpljTbFcmJH0dz+bU9DhVrutt+uHbuK4SaU7ztn4Dtza3PiQ9Bb2u8S
iGohd7Fpy3EDpGrx3eiYysTAqaTChD8kwEbmgXSHA+hKUgp+aGKUr54Az1mawhvd
YItLf82OA+xGfy4OPSvKO/8dqZK3/fEjQCzs4Yo89SWTaELjQDZAokfmu3jvmfdU
rXigSZuxp2BvyrZ3Cf5mZ+4BS+aMrHltO4LL4KsTd2IBh/LF6kk4d/x/FvDS3ga6
qoN2YMZFAioJuKMQN+ykmRcXdKt4qIGgqInvIZIQDN8tfPcq6hVg5G0tnomkBXbn
ZDWKn8Liu1Lzlr0PlPDQt0xH6rlezQqOsSsf+apVeDC2Wz22O17K3fXBTexBIBIe
IEE8OCtD1nasptTd6N1P0ATJWglIKC17KaVLJPzNHvCrDuAWJNcQ3sm2AKZNe0a1
c8s4fVw7JYsiBI5/EotsgUdOgN0Rc3BTFl8YH5Ea/W18YK3RN8BIdv7ejjYFw+WN
lil2pkwPuQGvGOgYL2Z3ptaBc+WjB/ZJsQo6EAWBLS8fpmuHjs9rsISk+au1ogKw
0MzfzM0+KIB9FDmOz+QwPiYfIQAWUEiTLaHHIfrN6WQ6PNULcIFvf+HwZNMPvKoe
PwVn6YgBfubXHBHFJmDc2MbL2si3Fz5pVa4SiFuOqcEayfXRllsv3QP+k2ot18EH
i3Fskymidci2nzOAeicewN4fZoX+DZ7iPr92ZYqG3NNcbehl09Qer8fHKVsn21vk
S4BbcsYKJ+0ZLiZHAcUM1vNVPPvqrr7HFrYIqXKutk+0bf6BjV/qCjskDaibFd4r
qFugo31UOEr7zgOnMeMJaRkIfNDxuZb4Yz4hMj7g42zG7mX8D3uxa8kSs3IDRJ/f
YlflGlb9SApcziuwiHg4RS3PuHD2CvD6AoMl5h+W8iDWfH85x+cycwpc5INf9W/a
vVMuW8hBIm0WK78SThMxxVopNNPUWIgaNAw6OX4vdUcFGPx7UOnwUN7r2wvNabLL
dTXrvkoKr+7FX6bz4Sm+0yvr6UoLhNLOAjk8yZguCTEhsjDqBMNtnEiBHLXQJCts
2tbAXXO6G5Iizrj5gvtbfWTxsku0bqiVsf2qF8SNNstZZ3VFg+KdcPt+N3acqItX
hby4CcuxPDQA9RmVOxxfvyzfZSm0upv+9TTudnOHzp+XJFZFzoJWdPKqDc/OuXD2
o1FhwA0/MO96OFs2lHtabosPQB2PZBM/viX2qQReRnJtf4ZlJ/ptNhdCUGxInvr9
JvPifRCCmBWoTzUCYwhhxmKSYzr5W0LJlFcCpaHW9pU3nzR+FvSNIuPrf86KIi6b
xVCPAcha1w0zjHskh3MrUDChBvUrdLmxa9WZ084GRNcc1Qz4GeUPU3+ClVj+T+Ma
6j7RqaVca5i6tPaH2DVwNFgDk3DOkuQBqp8zwHpMwyzyTIUUebRINiKPj7vzHM82
Md6EsnexJ0GAK86bauIhOvkhmGmuCMvHuo+D+ewZs2JeVOWgtYVqI+sPQZmhxJmc
+QB6Y/xBNLLa3MtmRklVdXnwv31WoG06fj5B+VoQ6d+t5WIV+Scs/DtFMRpuhYWv
ZERdHYHdDcF1ABXD5ZVWrUxV/9auzY0xl6vWVuE8Ko3YbM9my7dkuruF06y/h8YQ
xwmujB8r1mIzZyG5/QH3NCo+3TC9Go5Bga0Q1hyV0k2ZnIxKfhxJ8RIX1kdztiqE
pSBiAu/pltyFdQDNp8iyA1wX611W/Eiwst56JS/wGzj4CdWGHzDMUAh7q5zgRO8n
qrJmC8Oq3sKD7L3zGFp6Btl47msF1uTa7V7yvyJ6k34YRKoq/r5QQ2oZgBBjzTac
gwVgat0ZiJbomZ8LlzOtiztUO5AZomOfCvcZynadRApFjUieiJ4Gi5wJm16l3n+a
xNQY0gUc3y/k9f0ldy4I7UfD7+/PEygk3KE4xmXMGCvP7cnqUwD1+yIwMlgxF1O0
TGeogTTUznn0UnxyelKlAPvWGM6FrcNe4QzPtyVogOiRH4u5XgjMouY5YBfeRsgx
bGWJSH9iw21gotGQvt3dgrGy3sUxNr1wRWIBRGLUfEOjgyg0+TuPIvOuumjXn1EB
Ui/kdSsIkdlp0xToM8O0vMYBSC1yt059BDstivVjXRyCoLax5CIHO8vsCH7PS1Qa
dqZh0ypW+LggsJYxC+t2DRUU2bdDTDVYQmzVAkvspuB11vIXFQ/RgLIiM7krDSnE
ypIL1tCJEITxUZ/gh52Zq9lktM+iM1AbBiQ9MiuEYB0CtnQUuleMvs9vMw9HCoNh
z7KmZZl5hNP8zu+vf2YeJV2G21tWPAHsc42aQIIpoIIotW3s/fCPOYBEyQoagEsg
OeLNEuzpbM1dZOSyH9LfCI8tT9RJiFR15ulgCFqlN1ZV4/UXfxnWLaIvVtss5K14
Xpg7Ba5CmwIUm7isgSHqdD4q6sgNhcWjpt2YdE7bZLAFaXqqRqjToAtl+Wmmid+X
fjPuY1zTyczcWVuTUTGcvIZ0lJ5XFd1bLeN+ZUkSPNxWiLuNxHNIiJdbi9jyzQz4
xOkZ0mXvrGnNcFnzMf0p/KrCObRSG87nm32M8sUuc/AF7kv2FGLorVss+ktDTUMg
J/lCgaU8kf3gwFmHvnSYOikiWckDvhg0G5VSEo/qb8sK3vVraGTZNg4gIvmPBicB
OycKFjfTFNrHX1HINrbUzxscWH2KYqM4Cbgi+R7TyBoIsYYYxYLdRSWxzs8g1wcw
XJfJlHXi682CmwXNH/nkKGt5SKg7QWz62fSfHpHFsc0+JFghjmXHlKf7LAj4Fwsj
oq+Srn+d/tZMT1xoWXytVdkuZCPxnqakdHdZRRHZhTymkPcR+2pcz+AN5gVWWCab
2sVjB4PtAeVNEvsWJKMbB7spV4mzriZxIqLwx45HytzQiFjbLlhexPWG8ytQxWFv
OEihobMmhOuOV5ct2TymYgbfK5gypsfrxBEuDOQSUGQFWHmRR8CgvGI6uA6WQtC3
o6KXyTW5Km7Buml3JcUpf+vOIfojYYlMs2sQvsGvCkG0KEg0DNR+msUt1fphaE7a
ca9s8U2WXo/dZqPqwDHSCnqhI4xRP6C7GwRor0HXIcfOzSO6TXuG/jmTmGCgJOdD
DgA0wwfEsLDpzE4AmzVBp1zawzwlkCJTf10jG2kRnhaDGakntdkOf0ROZ5j5shoV
K48AFTCfvFrOoE3E6OxxE39tU5M9FUIcZiVgoNwqG1lYiq5t+/5Xb7rX5V9K0t1v
72ccCa/rDq3My0D0j4nI5/Rj7TlxGaGk3UmZXmNShUR9Es5uWOCs2EExZN38GRv6
6ijqOXMytpIdPSthDJEfsqukMjaZvvZ1hVNhnsfSXVfD7N4JkFp88eara/mfiAGx
LMFhNB3UeRoX3TVLRUCk1sV/COkYWYnUh39NyJl1yOjzoc8kFQGwUmxZFIHNXmyy
z3kOGlObuMp+nbl1hECYm+Yxoa88Scg4TKNA38qBNzHbzfyMj4kOOsecg0a1Szij
2AgkZSSY1iT7NTFBBZmmMb8u6l11MW+5U2SMqctqbLApexr6i/mgeTKxJjpkf3x6
JVBhrHP7+PAFB5xhQrqy+Dug8O9OQfB4vVthCTFjaV5I9wj3xpBVJ4e0OsppBiKQ
xLGPopenP/O3/GVioena7FdNwLRzr5ydO0kH7fX8ASxv7p9ObHlp7uyRZDNdGTXQ
VcUpQG0DoehD81DaqjsTzg6xienFngcWimyqP0CBbJg2YvxdsWoeCYTFyIz7Enuv
4R3KLKlKRGnvccNgERLzjMoJYesRMGcoUfZJVLXpnP+xJ6Wc+V34IDhh+IJNKKyx
5NJQFavnOdAR0th++N4nujk26rf3Ph8Cq+IsIskOQd9o9Vtg6XMGAnxbmoAhf2+w
qZfgPRt1JhMvKdHkt/reLtmQH/bi3Rsa7MNYBkm+mmtWYGXdt3XQ1q1BTUPdsTHh
58gdFFl/aFxjqKDedSKaJOmoY2bmUCmZgB6TwSxGnx0YBipGgeOqUafukuDVCrKG
bT6iHlwgGKVd279lsKTA1FlcqACe5kY2Pzg0py1qlOUGeV+NpyNQGkFFche6BPe5
ITjwASuCZAgIt+ST/GwfomCBFn8rflOvc+TXXrQCftXYngnnkYHYQz3XOvef2o2U
grTGA6aNDCOdpxh727Fv5ImzhwamDQxucbOvIBjAsGgJCkh9v+yg3mlSDvP5NZgR
PvmhmKJlHo6RR/XkTpXQj7TcYq91xONXz2oZbt6LtfRCI7nyOyb02pH+cIGE4DTq
C0OFjwbTSfxCEv37AkIeVooPz64rzIqvz5qz21wiydmSEOIPnY9ceN2vWsYfm82K
bjhE/xOJxWeizhzcb2vwENyX8zkTaUl3IKY+e4uVRcqkc9PdyJL3WlXdDtYwQSLh
btHLKzwLsgstG9rvAlusYE+hSbFJBVo5JRapqykZkXJOYCBkzsSmYS1hTq9SwVq/
tc1EfVEPtCTzpxVVEnjacrvVhCkIJ4Od4pemTUccXEJZRoqEevsBOmkleD3BfZn7
oz+2bLimEmurzrz3hBuv1nKykzuFhDHHEGlb1b1r1GEV6pn9oZbmdEhldMx48HBM
jwELbIA1toyxQrQ6bira7ZqFh8dB+A3isZKjvgmxXLPiRwxr1iChcQeAiTgaP+W4
j1KlTJLeTh2UjqDEYdFxYJttfx8epfbZka1dADomNiwftjdxjKHPgSZsUg4sQpX2
QJ4mUB4XMLG5pXNOMRPZMQiH51J9Se2xJTAXADcZZiQbfgNxa84XxY5AqN8JkND4
PlY8t+hsfyTKdKjd7q8o0xvTDdWBsxUS27MO12bMVzR8Grxq66kTWQUnyZcZ2qil
dLNfIzorGPZsnpOBX03N/DW9baiUzW4b7xezCwBDgdhkMVAHNqUcALw7SWqF8to3
NcvS0fMJEMzsA4a6oCYILinp7Qi2k+IM+PzIO4a3uQRQkejZw4n8DYOp0JJo5QJ1
uk5dvqaZX9LYKjzDyMLQHaLbGEdwdcySBTFHSjkgRvHGwBMGp7XmYDx/39zKcDq9
TJ3Rb9cHadQu8jtbVQoDjnlB27MtDp+i9d3vmmao2u7Xc0d7ud/6RBISlw0bSIDU
pVqU4ElGu7ud2hoBJ5EWV7V9xzWVuUj9ilvp9JvTLWbOFmSTP5Fi8HLpmPX070M3
FdgYqN5+9LYaDx+3JVhOug3+To/QN7rhSWX4IUPkMV60eCKYE5+WpWujjS7Ls/6C
3jC0QsyNexwntOd4DcXCRM/L86nrPqKanFHTReOGUHtH9HcDq4NbBD1jcSVeXXJc
NovoCPuepfsxxt0vagVrJf+sJFi24oufvWQrBx1J4kGnGFT1eXdDftpnBgu1e9Xo
i3pgW1BIEn0sBnTtXJakW7mwSz2FdxEV2epCesuWi7i1vC8tLCwZUI2XpkMB+Orr
iosOZOLZodhoHtbTCSbBzYd0ZNW49q2oZBKZ053jp+TH/agoYMD0EsO5VpBFnYev
dkDSIPsdqeI/4dKlTvJ83cvGu87dCvSIyr/qXz1jHAPe5mqsXM5eflxVVFXzGcXw
HzFc04AjV9fpRhJg332AzhV3T+FY8Jiba5i4J/MkAtrVpmyVhqEmOyEQq+iSfvv4
m+OFfQkWuVq+PEWeyDnKw9HzMpFop70RDCmkBLqAAiyqOhh6rQkqK+otWJ1XsAKy
8rjh4kydeZVvdRcLRn8CPPMLcw7tWnFW1pmJ2WraDEiQDWZuJjzIZcQ9GUOaVIay
v6lwKtKLud97f5MPG7Cye0HJ8dITYE5MyDb+ELyvPVR9NQ4olEs5BmCMd7kjax5U
c+6YlTTCq19KHO1x10tqUIHEO1/dRSTTppTSGAqYvPabrtJfPtQipOLkcDk4FNWd
3BRzE/K4y3N/v0kszr+t25BVgRvj5J0b3dWLeQ/O98mvQKUi5PzvfmUzZnWXlTXp
38vAugxOSROkCIGKLa5/HTHrbv/JYmJf/Fn2YSXhhf8Wso9u4jm9H/JPEjVrpahV
ZX0xipbludzujOnk21NHXmL/8ZGf2xVJ8Z+69HQRJjG1TESyDGU8bTAX4Kj7sw85
iIGTNgYpWRvkqJeAlwIFL9T2d120cTfA1iEAkPGVPIxjQoObWzQAlQAdQPcuVF9+
7xO9Is3jhHsJE0BIdMoPZheNrz2+wKcaRXdFAUKCqJkvc8dIC/Zkzjr85Uhzq7ZH
DYDPSJVCLmqwZjgtkjlsQkQ9Kcrq5HkFqSTZ8vKg22N1bofPOlPydfHPy8ebtRit
wHzDQaapl6PLA9dU7gMsKKQB4j+2aO0Q9xHSJPQUDEvJIDnfGVDvImapjScuYRIN
vQ1kG1jBI1wvhQuk2QFzhS1QIVz8a/zhaqmja8D84zDIGdSMFq3iw+iQuQet0gS5
NinUEaon5tkLqjWcXRFiW/rrn3C0UpDnUX8C1xbN3rZ0dEiT3+c8EPI32JPtFJxH
wkqG7bZxOFwrnw20EYBkGjiqzivcv18CRPBLQFW71tqJb+wFQWRUE6ed9koY68S1
TUbddD39lhyJPWnSauuNDLXP7e3P/PP+hLwu8CquC9hpMQyNjWbsmGMLCyJYIkJM
YknXcj/jq+tfUcNbs0zRNRpBv5rf2hcul3dhip4lWiyexKT/pD6455NpCzdE6GMS
PSM41XQEXVaoZiTArHlyYiA+98KGHjMDrNGo2B4yRqg1OzOkCaVoGQMI4NGx4vI5
3HTJEGDOTpFySPT0L2w33JzP9Dd00jP3uGZW701zAbKKa6dCOVqBikU3TvRctZU2
EYV/Ye10lb901xrJym6YpYHIb0US6A8Cf5xNeuOHoJDkgfaWMiomGOENNoKSrPLg
XtjoJ0K+reqtowprHz4OJhfZfP2EcnIvIkO45xJ/5bYwdYBuBCy4ohda2g/xvr6Y
8lm37/ejZKTBg3P1BeL/6L37xRhT8R6ZT1vOrvP0GInXZTillLz3wkiIYcCKcAQP
HpKKNGVpeWUQhuLkaEUNm6SLoEKCgXjfCZkABtoho7CALPtKju00j63IQ0isBJnl
LINnysu0eKUSShm/5fwpWKptgzo2fhXhyb/HTPb9RfD0EyvGwKiiA3yqJEeMJqFK
JYgGm28UdtCMBS7wp+IXlqJvV635GpoTV0fNwAHE/URBAaxNpD18K760NkOT0n2p
zMLDrqiSozdKun/pb+2CW7phcnw8kCGXm19jVqrsaKeHCgorVLf0oCGHRfvnkgBY
IWv+wMW5pBnHmZYb/lBffLGY2yPFznOZ8Ob+RKZyCkRMsxX90+NNPn8Yuma1I/3A
RLIrd3GfhVMsv+CIiRINxAfx4XYopbZtR4LlF87VPtpCfJfCatNGTeeDlMK0BK6E
jiaeZnTbHu0fifSieHZIpGIDZp2x77qXQ2JAceJPaLVJfKO4rhe2rCSZ2uQcbpfH
VD5fAzlhjEUeQb3/PSe1kYyagkvck3wvv1unRlH5ylMsxQ1W8oxeA0w6kQ+slVsp
fdID5VK8jW1mE20bjNW5h06IZsAIOj9Byx4wru4vU1NB1LV95NQE79p1Pi+nOkRJ
KNw944bbkHTVq1sJgz6bixjUKOm+p9CIe8VCysqdCNILNhhq9l7TE4JjtlLnttGd
f07OGFf1sI3Wg3fmRkI921tLj5ElGQyLSEkUv+87gawapxVyurn19WDYAcMgc8tc
tTbbgDXtCBSz06YlW2PzOB1u00Nd/HLMGaZcZFLFBL5HSfL/79hxbbNC0Dq0YAe5
TI6K7YlNTrheWz8rdMblo8MKc19n2clBSPmUoNhH83f9nx8Jq+pc2THCPRJ2qhow
kfuHPugB/6KwoD0PkG0yjBOQZFhD5vr+JNjqpP1Sa7nHOZfkw2b7I6DbLe0HK4NB
wiES1JOMX6S8+jjhKpbRqyWIxYHPWI0QwKwQAhPf/J3hwQyOdQ+EcXwAIu8EPdW6
4QIoSqEJO/52I/PFreLPutfowl7TSdPlViWQvJMvMOWTeuV8q+jYgCjV7Y3k7DnZ
8itJ/TMMPiDBsoU2F0T1p2rrw+5rSA1WFGp7X/azUAfRGwYvzMnhLGiMeTixzyUC
gDWCmBuw3orB7CyV+puzfDtzlfLr4EX3Xv3UM74jPcOlVjQhM2VQvTOvKwOGNIbl
Tp0HSkL9NF0EVQ2czRu0DxlOfJ8+bdVKhs+x5/HvOo/Sr0etLnlXnR0rxXv5iuzg
nnQoqlcl1m3j/80gBqoopL4mMe+g6HiZ3BMroNnOns0kluD2+iOjUuc43txZAjUh
LUUIe3UYaEbYJNC1Q1vz2oc1UD5Ivpzi4sT19LSjaotLb4qzC+FLz9LucR7EuK0C
ycaMTYHF4acDTz/qyCgrtVusF8JYzZnqsJYyxj/z7nq5yyYNjnqJZy8b0k9xMoZa
0R30nqsdIBnfD1q/N06Hzn25cqSkDdjhMdUaLTCCh0a+Bi+h/PuqSV7mdFYhwoZ2
0DSnKXI8Psl+A+cuj6UkzEcVXOVGPuXjhXyX5yeXkm1znPZgqKASt+EhQrEx7aOo
PkUuuuflcSEIO30x2j1s3H4TjwbHJNMK2whcfqhAGc0Xge4kUw8g1yqGRuItIRCx
Y/x9TfHMlrL7Kjl/zBFwmb2MXvuWBB3VyT0pIPTXa486Jg5CaAGpK7SstPWM0Q+p
6PbYgrShhxjxsBEKDmLA0/vFmqyp+uapY41ps7fcjZEcCniHZwzGC3HGL0Cl1PEz
d9GDDhqrciza3d0D4dwbz8ZFSOeXbFhbk0bJ3EaV4Pb5YZG1QkfV/e0W4F4T5KXG
IUYKEuMfEtS3kZjr4qMZmjovIdDyPDfhEsCJsTx9ZwOU46YjEQIQhckWWH4DlXjf
F6IOXhyfx4rVTEzHG9d+Euf9ag6lvR4bg3g2529m78iatsZsWA/19/bbjZuje6Jh
y6bpiepjuYDKqI/p4HVW94YYndEU/At8M2R9d+3uruD4mXXm3APDrpcRxtz5DfqS
H8NlUYt89vhiq8d0n/aT7tQzu5zntd9kBrl5YL8cwixZkmmuqsxTbFVpy+kZhE7n
3gtPVZtkwdLEAkPE3qM96QH35/XMba50QN9dZTj9Xociy8a3Y6TCkQ5Zt1v5ZBfD
TK2yJtFx6xEuwDkNtZO06GaUYoS6rEyMHDr+gjQd7nUh3ErJdcyl1fwtu0ehNQlK
z0WvlwwrsIB7fhT+kboIyeUIsI1tJPalCEZbS/eMjsT+5uX6xyugptwDf0s5oymP
YCcmuQS6OMBZNH8kEgMTxYTqGKLS+Z6x8VViyDTu/DGkKvNBSheSTssuwKWXQqKS
N5HJtDXK6e7ja9t3Wqms/4J0jWDgfspsVCPL+6+JKas4X6kDtb6hRT34wMbAblC4
GafurHN5wRrU8u1O3uD8JmONKtJIn8uXkaxEI6fbK/egrEb98fKjDq7yH+e4YlHI
GjAe6MNaDnJqooJAderBlYt0eyb0Sm3ZNhKdr8HiY0aUtV1R/9hw/HTumFxkAWi2
343qFHedfrAQiAMbfkIh1MJsyP7dv85bKgrsi99YhFMcnaupZPc8lgpY1JL0jlrI
JGNtodZEkNS98bi75Oky4QLceXd3F30IEWRo7FnVy80ngytuJwMSspbxee0n9usn
uPmMFhdkAdnYGCdz8ZprzoPsSQlTHLE3uBYy7jPFVeyXFX0wB4cdz7i6nvE1+5t/
p+28W7lVhMzLJSFr+g2BXuZ4I7issST0DAN6W8kJjgNFHh04fzMvidCfkeOsjMgd
+s15HsdC+N5y6uDimpNgh4x9/54iNVKUnWipAR6d1ap/7+O4BtLL+oz8YRKJO0C6
gjKP5VGIRkT+jlRlADfsaHsTCD1DsjZtZqCc6Fl0UvXTw2GP3t3VeDaOQBGw2b5J
dFX65xm2kQudMT/wpj00bmCTvs3yphKoUf10lnD82rpoTnYr0j01EYC8DhXRr3Gg
j0hn8GdzxfklfgSKsI+3A5KaumZ8QEqwAIuepuC9Ssr4lJBiS7k6B3gYDRa2k3WM
pWC79qFx12SZGWCFCzYifdtqo2DI2cXvAGfVyxF4GegGw96ubVvHO0h0LFtV+jzL
mg9MhtLT1zY4im90EdYYo3N2rvp+QAqkoNrNJ4UJVuA8IFDxR8OKgltflm1hExjj
Y+Dkzp9sfhYjsh3N7OoeoCitzAaTy177hU88AiX6WNVF2o3laAhi2ZDyO3+bvP9R
phKfxkSWKPjy96CisqmS5YV6Elr1zCTmbGOG44rrlkoSNkEdVwezAIyf9g9j1Ae6
hlpKbSA7Aw7w9afvdcXR5HTu+qxB749F0m1sa5NowCYEOUiXVih93Q2S92bzDU+Z
yI0PBzrV5PqHFazSts5SuTev9lJKf1gVBkbnnloHtMuHGbm5U0/Bpjb6hivsgOM2
pgKq/G/bCvicrivVi0VlLo8w3/NM94l8Y78xGU8SswoB3dGeZCgxsORvKDG/yMDb
KrK18dtpiKrw5k0ZZJ57fpb6VF8qqcY38OSzitXJiRR+bnGgJHuzQhn7KNEBz6G9
DXw38am6fDXHSeMnB8v1t4H6FSYjHxILZieNoWvl5rpuCZhl2mzMvGkBKcm1dB7S
BAMMttTBFXoejeb67nIKkCn4Q/cxhEcyfpMmxt4Ro3Kf/X7jMEyRbHimJ97TjTiA
COhT/u7PpLVice0uxS7ETfrMEPiRteD4YvrtJYfkmk8DiedfBTw4JJWdi0VomRRO
j/3tcUobVQxR0uImoxj9eKb+SCkQzEemv45qG4BBI7iVIGim0/CUf9XCnFrgTSIz
gqFMOoba/iSM/9H8fBRaeI6LR9jRsb0wA1qYTCssTHvmuou/zdR1BtF7dWU5msJg
XyyL+AxZt2xz3l6tTrdNOKGtjWWJqgOWe/Qk1aT0TtTIkt9qeP2NOrRScXFNqPEn
TMRihGf4qzyieH70Le/n3FiefcVJwsAgRf9ebDi5Ja0MV4i2Bza+U/T6u4kDyM4I
J2O3TKz6Nc5zT8qGCmrGxCDKg9mW66hINYQmoGw9eyC/rLQ4r8iiQtbAKRdTklbF
avm7W9gX2YW6MUPAPkhfbtYt69EqfkzFX6NCzaYs5I10NMuAqgmiOmIcYzGeYMoQ
kO3LPolg2fkdtrQBKEp7MlrZI3iBOR1RWDGlytDqdOiMh9ZvP7Fj/XrghaTmpiO+
0f02apYGaCv7jX2U80SCFOaoyfe/DF5NkAkWP1GkiWoONg740sXC7yUPPICTjNca
Oc1N8ejsIRv41kZv/wOUpm4pKFRfMMqSUv5JXOa4gJ2Rwaq0m8NaGBXQ03k4TUwm
7Al/Q4SgGBr0EDrTZtcJpkVAw/L/L+dI4FvGuINEPfwnCCVgiCI+ucyMUnuNUNNS
9g3V+BXVtgL5qwDWCvZxWV8lKy2YN5onJKpiAGV8kQ6hXtOwT1CqvuxBd/wL4jvj
5lpaPK/gz/I9hj7FSgu+wLNyoeTN2gZcCAL+/tA5TwudldhiSxw894nwT3kk7sIn
XerBjPchvicOO3reM0ptObNGmsRgarB2CXE+k1hk6tUos6aj9esrjPbVN4aF3sjh
7vIBpylewyTKxnkVRbmT49iezMa9GjA9dKP/8L5HNng/dIADLSMORXGxZ9YplUeL
yeJTyyEcfJ4W6ZOKfZW3VgR6zw9zgztoH8J0Eyvf//jMR0ZQNYIa8dGXMyiBblF1
eUaZPk4+AJ3Mm8s+mpOHfu8+79YJMcRN8N0ZeEs8H8VjPnFoiVopd2f47bteaS/+
kc+cYz9m6A95S5XA57Z8Pwu6AT+dlo2tp+EMSUVCfzXNW5Ks+Ntz09ek4+TIPN9I
8nYHG63kfMGArWTRPNAS5TfRcXiB8VjLdBwTQ9nlIsED4tkEACuliUsXv2z2wHKO
8pF6J31HZd9mgs1qtAlKKS64+oJfvvfBEr5hzqWx+1DhcsVD+y1/q8+L10a/oMci
ue3cCEi29LgjbA52ElbAakg0mEFVC4ViXoTA2r+GHTPmxzuKW+Y91l/jnOEYKxrd
Knx7N0rlW6io/2xD4+e13AF/AFUiLKVJdiAdnHaBLyRT0fCrfpQf3rHYLr7sG4Mc
ZAr4L753lNN9pW6eQXv7k1hj9Nu8p4u5UucCGzkg1ftTqbldFr7ZqcFwKKeKE0Hq
RxddGOfV+eLDyADkI0rkVku+6H3zs5/4lq0VMsKQaPngkYwkew4hqYlRkL7JS5Wk
65TK4Fawd5rt9sQWd7WCcQKor/59WhUsSOIyX3NF7DzWmRecl256dAtUgpVUrfCJ
e31jYfCmADf9kwstJHVAOwyff7fVTGOx7Hbnp9pmBOshi9a0wl2Um8TNTm217bJB
4436xKEUx0YviLcPnTmKRNclFdyzMQBjNXRIydn/IRjzhCyKmy7m7klFMCx8Qlgq
syB/Ggg34/LILjhNsqMYlhCaSKZk3k28Gpp+WkZOLRHJKr9AWBtQSGss1YH5dMF4
ydiQeCu2uclRBLRQR1fO9bOrdxn/XRruNo3AW+L9i35Pe30uwpJyIYB9SzRdapnA
kT3WQmrFMxIIu+YOjzp4aBzNimzD81+s0IlwqlGNlr1i3cSJ6oLni3IBa5njCGCy
RTLlCLG1+gPehS9eNNlq9wS5pA+p+W5gEiOFWKOVK4JudcCr5KYS6L3Fl0rO/OvL
gldBKHqmS0W/APCh+j1xcP9sm1y38gSbi5ixUMsSKZ69W/NvireQAeftA2LnPOW0
DIPzsJBiBq+6aKrsrviCW/RaaeNGnGqKDrca9sIZliT5HaLtmrIlfwWzQPQIosbg
JIEnHrC8b5WTcCLR6eHkmdu95hpN9Y8SMxzZx2aqM7XO4RAdKirAn77351YuWJY3
kZ/Twyo9wtRBxZPLkuxM7LFfKSa07gI/v2tT+bqcHvRRYWOSCkgEXPD7UEstbqQp
PcsMzQ3AewMPr4kPOWtudFHNusJCQZ959x1q8FL0K5j9M0luVQyI9E3XjRIvq47z
OOWCHtJ4hSveMxQV6pt5mXOQZ077pE4VLTDCGa31ZeEC8krizwhmSVSjbGXvN8zo
Mn/UTr7xN0sZiWG8NQ7buQVFP/0NLjk06u8P7HnZ9VmyiXFfzFp7GqICLHjz8oyF
ZudFoSe+sCVBkW5hpypriK9YsR1DCmwj6bORlp1hylW0EwcMn4TURtR5oRO1YX/y
UcVtrP3QyyBq9cXBTIEUWt8UdGJwbzSkfyg1nxobH/HTkQV9UcRx+K54OEGKGmxG
TvOOgomV+cRT/tOUfn+xzWNMAoh6C0AMoGhWvLfbj0YFIYt/0GiQiBJvP14+OdZy
Ix35WjWxbOLV4D6Xw8KcHBmeMcCTQAANSPb4bgzlNNxy5w7RGaj7OTWIo8UFxVgW
GsjmLzOaykslXdtx8mQPb59uxb5N2jqKjpYc/i+3owh2Qg1EEIMQQPH5l226o0DY
+wFRmY3nuBOao2ZT+76qdj8agbC6zFvBJAztKHV3OmtjgwcDgY8Fo0HNxaZocAZd
XqzjDDrmdm4GawO6S4oyVkmuKX3IwRMhsQ/CHl8DdDkXa7mOIvrvDB/v2nTyzY1N
OzMzfYpH8MQedctxhr+cIvnv2qCOz8667CjLE7rMfeME2JxXOpgK8QsmkH5SedVg
8f2vwh+pmlu7AODdSeviqS5hd+5hGaCtSuqC8JTiwxaW8yuM3bwlMDZ7DucogSRh
KOmdoNn5SkC99mIIkiZ+U9JPp8G56x1oXx8e/xlT0K9w0qxFPT9IimAZhoFFccQB
9ZDOL/G0LfuO6G5kMbuA+dBfguXArZ95Hvom9T+4TqJincjA0U1KrQcHxJl+ougq
H8aWoJcCQKoqwp3DjEkNQ9exmm4OtJ7BSxih8LYmhViom597gzShie5nQ8VjB6TB
VoPjefmHe8GWuJCw3nI+IxZagOXD6f26kP6BoNRb1bPpqSZzz2D3KN4sn0iIqDwf
0+Ddb86wxFs1CRan9Z9+34OjcWw7k5UPD/egau/wlxAQIhLhwI5i4KzRp9sqcMsV
bAg9BQ3rHMNIHlpGQgkSvdqNM6F8bXPyEKwxNwE5erVSXRIZk+F2zY3MIfV588m2
XskTI4tc2y5hPh0QqwRC9PufEoMbvS5vREWM6eqmzD46c+RIehl7Oamwt7JoCHF/
yA3kOsvQ6jBxb2QVSbZit18rrjWg/oiWkTmC8vdV4ij502EPGKfMFtH2H4/QiFv2
OVzAVhP/rJhYgeDM30Wxrblp1eYeJSv7nXQSd9y1RTjS1Xzak98bjJwMry8Gsp7u
Z0jj5fPi39Dn7PlV2+uHqREiRcJxDh66lvknLudSRHXdapYASBEX9PSBCS3bh2yh
TS59qi5VtZNBwaQfNO7yhbLae2ZaeHI1BxgKjh5jk7vBO5rUPnd4eKcG5NzTkU4g
DqiG8ghJW3tvCduFrbVEEFHiS2TvE+z5r9l4qLSLIfsENsboYCbtLp7xHEQi0g8z
+QSDF2hSF3/+5HVleq+a/oPCWOM0nm/Vo9EAO53CoXVYGoId5fNIJ0qtx+QRO3CX
92wwS47PpbzQBJvJ5QW0aqeoGedF+xvOf0NPYHurqtOLAI1OBu7QlRSUf4yn+maU
8819gacN3VHXfLMOeGE9RgnMX2nFPnv3rp3yicez9oPuL4HO96783WAjCf+MgChT
4S6sZECzzf8wwWb6fdSKp6fNcqRgvRshly8xhNGF2J3V8EPuAkm1SezN2EeOpwJ2
drqWscz+Ik8PITuFMRMWkR7kGlf4HEqFbbHLlKmHjG2HU2WQWjXxD6Lla+K0zCTa
yZiOf/ZRe7JWlJcPKz880Nx8b+XF2jFpE66ICoWy6RhCDe64tGEeTwufcR7C2PDo
xKtwVG/3FMrk3eSIFcTUNHjVM1XSV5dMYHK5AlqSIBGNwcd9Ty2KOBe28EjyrHQ1
RWJGCpPidCtoa3JstzDIIY1OCgN0opole7V2U2JtYFk6h5uKsP8c/27Y1gcC9uuA
k1WTl5hip/GnJzf5kaOOmnKUpTD0zYcStkcIhJLNBxSxNIvN3L91Um4P0eaH8h66
0s8XuDTiUSLbvlz2BDTxyGeF3jgr2RA9/g0p/Am4TlSUQTWDbeaROXuac4y7oLJi
6kDmQtXOPiK3e+9/b/m4G3JQRkaafLiFubSeBhVph2IrRRbl3DmFjseJtvpESS/R
UEhQLTnqNEgUuBGiMp5LsqWW0/LkLKhketNvmY5H2XwXLbrWZXPzdK+U+3DjEjOb
xFUWehQch/L0tcxL2TzWTqLJMH7roj71MDrYMwQvqZfOtkiR2vTuWbnXNZEetccp
3vNWFcrOJMWV+0i2s2BVu5JGtV6X1Q8zskzjpV7LZ1+KeA9ndNd3GNnhLJt1w+fc
iLpvw3+RvJk5fYJyatEeic5YQKdlQPzbTyezeOf9ljKb1V6TP364jKmj2K2EKxvW
+tEVI4p647Pwd+DXk4qQRffKnzDhmmTeEC3/emhT121Lnp9hVrhUtblaSztYbrr6
sJi6W///6zpmpJqrnkob9PBdeVqkAvuCjpNkGhkP+YaZQYDzpF/FzV9o+pmY3ir/
lEh1HjrU2BEcZiRY1REy/UMW5YAQh95+vNVF11VsvAJ42rfckXg/rEjHTPBKAiF8
XjOGVOSmR122qKCgOYK7tIjCdFhDjxTRn2NtitH9zzXeZ15swyNqJ10bwHGW94He
J76v81rWpc/CzoVPzoBYmQH1XNyQI5pTHy8c2NCjjCMSHGeOuZoVEwfKIVqPsfTP
sdmkI5rGS5vcNtR/xFr9qy2SDnQZwNatoRtbVSvxi3SfLYwXHu0A3lSXtOhP+K6u
GWFIvQ8lYWjAFUvLjdZVvTqn5BLisNiWgmM//Rf2/feWJVyGln+ZTHs2R+CB6LJd
8fJOJ7CGLpOyPjFBjgTELXsWkOG5/R1/xeTMKCsxKIA/fOz+lAj0nz78DzprFfx+
6vR/9xNFXgdFU7XdD+77EK+/GRvtk0DCxTRWFxjQjJLF13qDLE45x3tVUvyooU9i
uYz0Gi+xkI6zOXNCbRyQdGVNcFljeTBWkyrJQMYPgwUG3JmmRgS49cyOMQFvhwdY
7AIttyV3kRQjG4hNglgCw3sdGpZ3a2oGSaemmX4yo1EwtaUpbBcBHdcv/3xqxqZI
48yBcT3+5eDnpAiOFochf6dxUhzG1gTfXZZjzF/V2Q99d242YYCmus8/LmWSpF/4
WnzSMXYVmGsYCwc26zKXPUBrEdX6pM9WS0Zqe4euVMtXUsWFEMM194EOaPV6ny78
Rk2SMllvSqP4D1Q9pDh0TEj+98P2XnoPEwU14I3Gb394yJezPsDFcQl0XvgsvBJP
AKugTUxCjbL21YDWVLO1SV6cHamX0akLuaCDMKO4D8IfHttBiD6J3EDTIo3ZZU2I
hflFSy/FkRrf0fG91/8VHWKz3yhQudlUHMAxF5sPk5J6H3GM9qp64rp2/Bcr3Tps
z8JV6JO6h+vX9LszQxmA+WOxh1GEHYrGEjTlD3tm5dpm6FwaksXnPQfBcu8+tcXs
UufOCZWH60u8VL43MjP6ZEsAcTcZ7orhztbEfMR7naNFRtYZ9LaPizYE17tHgw/W
HTKKC+tcbeXn62NHqmglucf5L4BlNdLRhVhN8u2zk38Lkfcpe7qoOhmaEt4c6ITR
qC66Ysr5LgvqOluJgr41PebUzLj9TsHleHzg0/6J+lCQ4UtMKinj3SpbdH8E62+B
ybobQ58az9uZJg9zNCjVhs6EdU4lDQ+T+GRvwHHw6Rs3mfu5PxHBAkYhvkqWCJ1g
hgvQfKW5gsRuWMciJWpUQBl3w5oajzkxBj7owPDHUOssuvipkUK/Jc9lb7mjkiUi
IDMxcIvQMSBVoR4mHTPDglPezQyvk2sncanqtZj812MAXhE9oNmT9LBbXfyMGppy
aXT6TYVRkNKxqQfwR92z1jASLsNukGVyTYVzvvBKwogrO8oNNeLb4zo/9g2xC6z0
pSf1KM3J6yB+TYqYMmDERMiUcovFbwZaT0H/A2QKb+HUHs9tMeutX5LNkB91CBXZ
lyz1ih4FJG8JAuVzZ6lWXyaEhNkBC058DxAdSuW4zzhncLe24TqJ8QXpL0L4QqqE
Dwkuy2L3UlKDVyv+D5WwVC/bDaOeKQPmP/32HMetkby6/a+ajiKx7f08gNOh1mZR
JOksItDX53IlHcqj7O3izZM3pX4Mo/6rbxJdJ25UZuCQXKUpDOoJO+tP6dFXNac4
MiFpVWnduS+tuu01Ts/rhJpshn9zf7Nqoa7PxyLgypKHpdAi7Sxg4W8Du1l3vdZ/
HbAT1D9874ZWd7SWMNk7rPn+hlOD3ak5GnIOVWqXHo8u7M6B2IARhYsRWm63D6ln
DrnE1LH7IHie1w/ZpsD7huTSRV3NdAAdP/EGttME5EVUkI1dNfnVD5RussoyUxua
JpyJfLkq4IvFQh9eCeBQbhqw1+hQuKTMaIrwnF7e43+K0ClvIR5r6mxcH32k/UBB
7/BInVZqXPkv6/qxMILRlJV3M7ZpxdGcZSMKKYo0NJv61B4DjdLTh8sVg3wYHcaW
ozTDbwRDYc8nMiJXNfKfMruNVlnQ0xfCe+XxY3dW4r8m4t09dQhksC+moORT725P
T5cy3a7TvvOVmA0Zpxp92lJbKhIH9Lwzhq5NE57Kns9qrRsAU3xbPRAnnIBHNKs9
9S+xWrX49YPG67MBcTHIAr7YIo/msIFMaHSy/aGfF25ScRRbPOYHsfqr+w/o8o4X
ysfj62ywViZVUw1K1var016tLskLLa0IZafASS9we5WxzKqchZo/9ei+/VCfJ9V4
nfPJQDAcaf8a8f+W8pEBLlyDy0NQIhv9NkwP17QU+YCypd6fCNqVZfw26uFPj+Ac
bjZvvoeEKyWqJZ3YwD1ocZLMmkmACLhEJL53BvsLCHi1TNw6PTGowFEqKJ+jkR/v
YV1vmsu+Ht/l32pLY3ZJFZrRtTCS2HkjpKNyDKwmUShQuVWwxnEWxR45De2ONS42
DW+NnOeqsvtnNNDnDHNQki0TKEsLDyH6t/0PKoKbSa9YRIG/8Vgglb3gTqk/GBlm
xRvBCoAXldXwYiWUW9iVJMGpFfJ13gLmL6kRkI+yks5P8v1O1KqtBr8acyJ8UNme
Cld3y2oLDok5/tDy5k10epC3ROv0iATxCHjAWY20UsDRLzz+ijfS8wq4eBNwn4SS
+izNH+C5Dnlju0hFNqKcJu+sQW+oqJSJjuLqUuR44wK7h/pxzc6HD+ItS1ZiIZuS
pCpveOYkw0Ncq9kOfulbelPx1yKRbPpooAP/+2kHazWHOmrypkYNZZhmclCI/3Tl
3fXVOSZpLPYw7D/RTAY0qa9nbick5bj68ukhPBaL+MEz0VAICTpEyex+wcbm8T4y
pHvQlO3DJPOSK00tdw8DTdEzEyvtZbAzQtbzdFOz2adNKw50bEtpl5kJYbRvcbd8
CNegmqs3SS+aEf9txeZfgDhh8yr3v7Rg97gJPnc7GsS5MAFLVbV/2me4wjNOKfF+
82jZenUtI5uPHiKe8U8AUxkoCuYBVwmwY0masyEPfmPsBAO98rjFPql5DaUxHjCl
IlrxLhG2WQwxP4pK757xFH3H7/wymymTnf/h9b+Zw9T7ECd1IC1u/TxLAi6FTWT/
oRFkitMaa1utA04Ub75Cv9oNRqwQKqDWacpbuF7ouPzBg7dPCcnD59T0tY9PvzvK
GHB+k6vb7Y1W/dZujAn7suDCJGBN9kYZ+GHKm2gQM7vQuT55m5EMsSwdJUcAwWAn
mM79iv238UP9U94LfxMzmvaUSKAe4Fz4omo86A73s8FBrIfj479D15lR1Gsi/2ml
yNvfCNfQC/0L2hs3SamIE7DtG16qSaymj59WByUG4kiyRcJSPldHmiSuGCLJ65L/
HfnWeQyVvBwuNPqLe2v5k6fQm42q4h/b3TFy+VkRyq9TTJYFibUL/+wInnZ+/bFh
Y6Gtjd+AjJfAHynOmRCsoQw3z7mmjCOREvQtIbQ8wKQvFw05NtQ79K9Du75BgScW
1ZZ4QxcRoa35mbsQlwjPWx3/uI8xraO4DY+pfxELL1JO7QCc1TGMKDjLCaa4MLP+
rr9KWgKr5klY6N7uhv955BY/SQUIomwSEY41rZXeXf7/7xbYklpBWS3UgRfiN5yX
0s3Yi2omtH0Jd44qaXIvlt8xCxJ6w69VQIC6WYFsVclkYCZojD/SnagBqvBAg7/p
ZXwgRF1YJJ3ZI0LJibSk0tU5bfPRLpmK5+GN5Cphj5C+jzBrFZI4Z7QD+6UT2vh2
X/XMblhsKH41yYvzOrBD7++8LiO0eQ8rdWRjwQgeWH4AEZ3wf5aON8MQvmAd2I/7
1hz7ncsjtdXO/61/Q00CBba/VwTsPU7KyjMe8J/PxkYqa1QtAvrLy0/7KJBQ5zpw
LVoXOgJKbnnD3dkbxiHAYghhGqlvVhluY2VaryJFZKUN0iDBzyp+WyjT5I9PScS3
ydriP+yuEBMBGhnGg0NTmF+1MvIcR4XWTG9+XZRtttMU7wRl7wfXGXApIn+Gs9+k
q/Qmy1136c51ZhwfhzoL6TZ0kP7IPFxyEWL0uja5UGkaDkxIjT+ysANAr0WFMBYd
pYd4PC/6l4MBY1ZKSLlr93iCFcL9x06si2M+7QPW6NvdPL0IISD3nNjtPlSTyKwK
IU0GP3HfbWPF8OZXTw1K6JEs7Ee+ddhLNViRq6Bu0XJEMD03B7CzkGy+PIwcMOGx
vHVeu6lMFjYkrL+Unr6E6H7KPL6mOPzlzkhENG8e3e8jr6CFaiQgW6NiweNVg6yq
Nes4ZSkykYx54kC/jIJssQ+nDirtxqD6kay0AcwSjPjXW3YCBJArW1GF6iezFfpC
WhJstTrDBkMBhAn+WZFYxL8VF0jYg26tLW4/WRVtPZlq6eyiEks7xnI0Nsr0i6/3
xEo5UKz40M19D5cWzuGd34LEqmt1JANe8eo3x+RxuCznE/7dnzIJqt7iryJrlFuV
ttfxyK5QwZzw3WYfqFIrzUziuK+VBTLXEwoUhlmKWJqDQebngiiejBL2/1FvWb4N
Sk54FJ6kB3+2gAEE4zVKbkkmg2fvT9k6wQCH9kpsPBTjLDTclW21rEzi8sioq3ca
0y6WYxfS8uoCl+OLT2Rppt7UKnK9sZUMyf+v3C7hQP3pncYUAG8iDsHKegg6cdJt
0WShY4qtTPlQfq+GaLMvN+hxVSyDW4qFHl/LxILq/drLpt11kYmimGtWaPHXdE5j
eVrHIkTP5tIzy8cG+Go2Nli7tSvVAGfWe8f6p4uzg3mNnvA3UJVKRi/nacBZexb+
/GMmeQ3qDy65Mb6QvWpadZ3WbaPQw9G0e/BaXNfH5RnqvJa/7f+BvuzHjZHSHim+
50GlFlz6c47NGwC22RfLW2VTmgvYPoctxDqjrm24FPOf56Gt/ELKiL+jdRQcCRt4
AQvQOwxtJxtkynNM1C0ZvQFt2//5A/wpAF8HzVML9Ka2FJogJ/Elr60qgVhbMC0l
1r15vjB8jhgn0Sf1vRdH8z9AaW94UIlWwY4S3ugrs6K3AybECb1/KTFmkgjJKcq4
k2Fs3zPG2xSeaECP+d+O9HIMcKNjp30yZVnPXhegyaRRELGpVeWcWXbm4evVjw/X
dckJCpsAJyfwhmtY1H28I00mlLZyi0ai9tsm6U9vn0KW8yLXStpjYLNV74UcdBUw
WJc6dqLA/2TOF8Gy4X9SPG+D9gps1+0c1E7ADlNG8/V+CkiYnulr2UESwORRKr+/
ktdv8IKutUHe1S1tLJ0tLIBzacAKpkp5B1nP5g88IzGWTur+U3yeSDkF5BTyOisw
hHX1GSXLMDCsxtUrJD89PMLAB/mdBiG4XukPjz0TuZqulHNOT+wQofM/fh8J0gEK
WAB9KKDBivWbsIJqtnm4Fo1CUxbNWcLtgw7/9uw1mnzvNNVj9cAYdYIuIyAzO1we
xEAMUT6JOLZF9jKiKyQV7pJ1OUFRsFcJ/XHVe4Rt5cBJt1QNNtDxpkuC9fKAWB4k
zDvr1vWqQj5l1xDzo8ZlbB+rkjA7tC86MRQydpPKPw3s2FtzpXbIx8BS63afRbUB
+O9y2IdrK9tmPPOz4gxEaezmiWH7pmsMXkMdHnZ+0+jvvbVHf2jbk0RFn4nB1cwd
EjOze2PB6XYA55wlDnxTlF12LrOlIZT/sKpZWjAqStrFK15IAnNmVllbjwp2SbJm
7kEdqzFb4rPPGcADvuHh/SuBpXnU2k0EnxEalR5MWO0hjVDq7UVFuDjJ5m3OfJTr
EYArMVoPI6lF9hCRVGCDkz4T0qCPT59LnfnRwrBOD4r34c+SswRTmhywqYK+/1XW
yV8Jl7Ybs+8WOmwLSwCZjHLbUF2GKOh+/L6IAVjfDDKoXk1dYUIcfl6a1i+rZQwA
PFGiolz8jcxpkmTTm9fj/INyWkiF3cSK8FKuu4Cx0FsnNlUUDVzGgHVHvhnAQNz9
bYcjoIrYDMzbc99MuN7AAChrvoD5Y6YXGiTHpVjq8COGR6eD12m3FKU1rv9fXULY
WJ7n8rTI2+msTro/eXHoEmxFyuahklBHVz6BeguxbVmkm06rZIYImZHXKPffkcma
5CRNJQ+t5NfCvCxSuR/4lXSXzn/CcpIfPuBHC46hL+ptVaqf+gGj291tsFPHRvPu
GaqBm/yShuiLLU4UfigpmKm0wuEgp+jBw1guYwlEDKPATqTDZl0owbNbH55PqmOU
L4niooBep4+t6BJPVZLpyWBgO5ld3yZVJbocGYjn4+nQMF3QyBYzRbsEXil8kQMU
5xTt8p4nJINdko9vyPwyq/gTvYmScWHaO/xssGlXIFswI5D3BzbBU06ED9ZaFdSx
kgXbiZJ4HiuIerWgauaWT0hNS93FzGB0FQ0wKn2t30cILB9nlf5HYW15HdFP/HG3
DgfN9RtUoj/NBIJqCEQKtsUL9juc3XKJdJcJLLlzmkrz91OJcYng2p7A5REn/etN
wegL9wUBVTnwC3YMdsYubj8cqR8DwGCFrseJjz3Ka/dxLRElo6axz7E3d2x9r6G6
PF0VsNwqZ2Aj6/Eon2fpDNc3ax8RnS5mfMBazlobx0/ezLiUumvEVI9EaoqgghRC
ANhFGnG33t28HIdh3siAc79D88sWfdzfqxQqek5b4KhKylqEnivmRCLOZ6J6VGU+
qrk0f0LPDdccFL7OoiwZ02T5ezuIorxlaulLQr0iKqDtrZiGDjT+tXaByYuwT7+9
lY882ulO6yW5aUk8dW6dH7s7Ozf0LvYZMAISb1dL10aiH0aQWFlnEkOhLqkViTLF
yn8FMRMx4dgljlEPB0oOcaZYb1VDsBdHcI/lUXeEEKduA/AYO2Syrv2SO8cv+ijY
JG+43jboswHPMsyjDSbJULvUGqEycp7ZCtr7ma9saFbVCpFxF3Sm1U9R3fKbMWZ4
OCw9BFLeN97mcXeuYLjXctrtp6Jfpx429xJwcKuOwM1BZZuRijCxIbJLRurve+y8
RuUJX7yFU9wRy1xMjXYFvv5OoaIeLazLto78Q/Eqav5gWAMaCvCROiuMdTFxweqo
L3+OOdTWSVNBXNHyTHmq+1f5OLDlM/jWu5ge36Gxuag5jQqQvuT3aGw8US/7TVBX
/y1CDOseptcVr9Jm0t0eot8Ew/Q4P0s2zTFKOkNZdCaRt5H4qUaVGAX2Nc01l3eS
yH7ZoHw7imDU4TkGBwIrBvkgjaQM3FpjzZFKIBfV2nCHdnoXLTTHBJLbf3kd6fTg
i3WL3R9Wt1ENR0+Sh00WBAgIZqfBMbCw68Zwj+h5gQoATEWe5rN70cg7jigMdSSb
nQ2q34NJxvfTiuhjQ17Gdj8Xb8DwrBi7pLwHDEIneUt7lgqsWaMw8zAoNZXjBMSZ
oRR9ehxhx9SdI38mdJwXQKDe9EmJQQ45Y3sTWEHi8X+VpsK3B8nN6aqG4MEvJUEB
iyRg7PKawQPNzqeZrEif81M7FcoOUu5pvNvbGMtt/yLKoRbfmPOJlAXdFZCmZFSc
dQkHnWpt7BIHr+QNlYYHEKiMHfnxGlqolcvIHSQmLQgyUnCMNVFkFuIZ+AuC50Xw
2hWkeOoGF5VJWgNKBS3KebGukQxV2xcGZc4rZTr8RL2vmuSnuuO/MKNVTPnLcgvR
8n/C2z6GbnnyOBHsqo+IGQQs5a5vYCzYuovOB0YDxQEhAQSMz2EBQfizym+NLDZL
bpgOeyVu/kca5euqf412tp3e6YPZ7vhX6K+rLXox68OjMpGNyYOBvPOCnr+Qh/YY
oFye8xtKPuix7rg+UgUbAnB0tID0shAPLuctHE26gpBdDjBAo3IWQqZDHzfMNt0i
0ZLolhA00VrRR9xYXx+lARNt0PMySYbmrDc309nzoTCRLRtJn4ZKl8vksu4DI2Jf
YQ3AvjzkUrJOOeZCcqAgAJrw8GGtNtrYEnyD+OO55hlnXykF0spO9VUe8OGNp2I0
WBASrHJFWccPhB+kvUojiJblYkQxzkzdcHLhbNj7hcVuwEiiijkZW+/QUV/loHRj
fWJmn5ftCHqt6gqub152h1PUz0lCjluJ/Baa5ShhjHk7uBeYaSynQ8SO7dh4YxmL
Aha9sMVCvDBtO6snxgy/NAjxEI+DPD+6NQhi7ysi/Os/m0wH30oDJlfNqu1LYF4H
oERPHyswKcOVTCJaGTXit4iI5W8celbjvbYyaKbHEAls1FYbgNjyKVhu4coajSfY
X5K/L27jD7dh9UxAst83JnuN7j0PhxdT48T47jpeV1smbP59dSVCo0XQhT9jBiDb
hGFVzm4ck5B/3d12xnRxrPbUd/o+PoNJyg4SELSHvJ69pgy4R2yz9tOznTmBI2Xs
uZTaljVpLcrotS+0AM1Ni3CFCRIWlAKzXiEOWOv1E1ikcd+NOswtwBrOfEYkcttm
v4kU+3F8deV1pUig004gvBDUa9sFDSSzGlx2/PlifRmjztIrLSo9LQZVL2PCls0i
YHV+TSsD/ctlYfA0DAwlx+6oyPc/t4UL6M6suGp91rCikIGhvouf5KpUbxaOOzf6
lfMJvSho1q3CvNiTSpUoMCtT7RzGCL5Qk7aKqNYUa9HI6gAae1gigCopPCd4cwBB
GYLDJkVs0+ug3Q5zG65zUZTlyeayVFulpOhPdGs/2oCq8FGFjnZ+SovLIPLHCswG
rmERo2YB1faxUs3AUvV3q09PYUJ2EyqT4PeNFX/r3Sr4s5ke3g0wIhTWCGfb+enS
N+IMdr88L1vvk0+f7IkbGtOx1fDx5jQPW3j/Edzhg9nSA+fFkYk5J8PFwOONmACO
uUP8zO3vBaMgNPNDIsKmiUK4926EEn2KsYisr1dgdbim36SstRpFfqTjWxMB3qhE
5I1P9PaY2WXa48KO2Mw4bNGlk7lfFWIpC47jnLRA3lFv9gxCLJ6GXG83I2qE9GEW
26idMcwWa8lH7a4YrDH82Qif3zXtygAy8b85X7QgFRH8TLOPMVVgXjPD1o61B5WY
LcL1z7VEj31J31AFjLznwjDkCkxRiJBy7XvscizD6C0huUf2wgYbZhzGzc6HgNou
FUDCA3kzWqV/mgWD+SBeK7GZmvlh2EsfpSuAtCnpypF361oQWji2SjOhVISmQ8EX
Vk06b7ZBvuwEEoj8/mWeIOxwGkhJ6C5DJliGHPiZeexNRp6q74mdiA6WUs4wumUJ
JR5UxR9XHFgkxgVWCF/oIyn1KBXG9sBxpFeLO3ahCr2iRjjENjBRYK8MZZwyEF3B
Ruj93/QAjgWMPZchxQwB473OW5uZJYifiT2fnDAAnv16kRajaa5FLswRhwiAQh7q
tHHxXXcPnxj9gcGyBpZprtwZeqkFDDjWV46ZS2+WbDN3/lhmMtQXPSYsVJlrYIPX
z/tsnmYuQxgCiZzgw4ajxKsh6DY9BPFmrIWqHismqIOeWVqH6DsD62EkIN08uPp0
TAd8KWWerevYpZvdpXFAGz2OThqR6KOzzM2NvQkc0+RxeRiSUSfJo2MTN1kwqT05
0eBM945DMInG9yo9emRam6Uad5Nq2HNFjKxXL8X7AOeWwlfnc/FBLNn+tiNYSf0U
L3cMVgkXYaqwtO8vUnr2uKeo3Rxw7ez2BYsTLAplcB5RYxUj4q8w2MYp9Kcb09u4
QordYiM+in67C4mwO16tpLHzqAk5ThzpcKTGsgYM6HAxGjBerO5qVpboN7scnTDn
dE0R+7zMcLjhsztImcQ36cCJ5W0+uy9jo19bmEYgLz4U1+LTPgktdSFqvMKu/MCC
SsyHNnWKFwpNPhkPmiKgxwUo9DPJDcT2JfDMuAqqStrQtXSO4rh8JvZ9oAIK8kAn
1X5XxKNi+EibVPOc2susI2Av86Pgeg9qYrw4fQtIMNENw1O9NSgtENClIja0WWoR
0xJTHgF867PQum6WXyc6WDTaekyxtdqBJr+1YEj5Jg9BPrvWwQhbSSGP0yFhNT8p
r8pDCXqpK6aWeOvUQoPN/x2yXnVIu8OqF93QZ2SJ8svs2gqrZmxWNCptX9RdExvC
abHuBVf4US4OrPblONNMBsS0C0uF7kgZs02XDv19zwqrPd01l1hiZEOfu7Hwmmp6
BDibLRdA9U2H5LmWusS4kW/xHBR1mHDb4njrZjFjKqNw7uxg6LPLChP0JdzTFU+R
x0DdMxjDDK568Z8H9IFAmgOW46ckOU1yUjDGGslv5CT7J6VnICY6rsBtc8vIlN3t
fFc7b3Pd5nyyvpfnp8TtUArYQ8oRQ0jNaRn4pYa+hIsEOIE9VQsdm2/OOVqIgozE
4qS9OC7tyvljE5zLtMU6MjU68JTHvhQFckykT5zu89Cj/ixkf3eTjebGf9A+g0Pa
8hLx7JKxXx0VVBpmLDOkk5uyBkikJQn9oLpaNnE0qr7hKyAj3YFdKFBZ3Qt29Euz
9Vqi/SMq1+rkw7KLNllEY7tEiEcI1PItrsw6EJN5N4U7HCqaoxYvqR9oU62DJ7Wt
zonrdZ8/J5dnLn7ylZv448hmAMV89Jv33PHjinIonRosOM+uxfFyPkQV1OWm7dac
JqfPZwocU+s/Zm+CDL+8RaBj4MZknoBy5GJZald99/RmoEU7cVJBQoaUmcvezE3n
/zbsa3CRfjn9uSgAnmNmg2vDdwOhXRo2VT4mkM6PX5QNBMPQ7aLGm06XtCOSHfmZ
UR3qgvulZsHc16LfShFUvz00e6I4nM45HSshDisubx1HjINRdzazUCMfisH87mRO
EMi7pDh6u4vRfxGwiOgw0cKlSjIAcfv0CB9BiTzgrKXxeDQHIxnYr4DlkRlohsdv
twqjqrgwZbJF2OWw+/Nq5qcNME6yVEnNxkoA9ZzXVpCKI5bdklo62/MZ8STm0358
rNEVBsPRY7ebNmxqDWhi9+cowqh25ZcT82W/8EpU3IhRBIQ4XYKYbz0mlydpQuKL
4a+1xEzFSxf4fMBs6td3igYAs8cf2x50ky/jMLf5dr2ZVUDXBVklzmu03VXM9sEK
6nZWB9fW0+al6gh43MfYQ/NrOICc3RXlh995k9OWpd8Ujo/Pkh7ngpMIyT1RE8b2
nGvLy7Z37hUhjkNeNvDRZfVc8tyM8PX+3BOxDRBWxwEiSsDenL4TNR6Wi+WDXXQc
N+mBFqHcHeqWQf/66V9BdJ8i2LoLy422N6v7NRv3ZOYYRsTwL/2IweTm5+3E3rrL
rA9mJCicTDjMJqnz0Fug+zYQwE333zv8LetrxAt6ffG6iKcejOEg+qVH/2r1JSmH
FHCaqEgx4YRiuNVkmetu2p5oY57XdZ7A3r21jR6iVNYBQPFhoPEeAUrPEE1qkesy
4P2c1OiuWkAbA4QhfMtArmhxNyLtLuTS2qBUQCdS34zjYAltdfpb003UgDNOaeH7
T8FsepbsHPqAnk6ihjdE5+FNiXBDViIhwGeX6tJl+IRB1eZZgPAwLmkbrAPYkYjm
cOvvM2vH0KKH2asggTtU+dMxZ1fQvEtnUSSVFMm0Zqwr0lqeJOIOoKkNhZiUsgl2
uG15fClk9CWMhU54E4hvmIUz1pcJ4mNCc52Fkyv6U+kNCkEYfvef7ra1Dfmw6OiO
qwXcSQx2L/GKa1Fac/RXeGNaBUTK84pb5V5bLwRSELGvEq3a+cWpVG6eDaEEggTu
iET+2tb4Unoxqwv8W8Hq/3zLxxkqKmVWfCFzLrSyNFKmT4j9luE1YCHLNkJiQLRU
PCPywEVgd2blOZymQu6OuOAUpqkPPSPy6aClXolC45Tg6JyA9MiqQJdq2foyUDUt
rLoqgl+7WiP8PmBvx7w+6Q3MzCrHqqiFTfp3u96s9dIZGOAKFDhI3LE/x9ypqSQV
/VPAq3kppaoDZcMnHucYqIz/fmim7Ln+xKSwwSmDF+hs9/tCncVNS65PA8mxwO4D
p0eItMJxtzSMQwybECzfF+N/779uSGUQq5MucVJwde15s2zTDx1LYe8oIpTAh8D5
f0GtpbE1wK+cC+/lo2IaOVaf0KUoY76UqEsqncIK6COKnhH8nXzbHlVY98QPQHbA
QiEfAaRmm0iuAgI8LNiZM9WMpcC7KxS6ghyw5HrobFkJ/2UFE+tcB5D7M8OR47NX
Vl2iPv9BsF7/vFEopfpLPizcf1Xyf3H4JjkN7qQdKm4qDSXV3w0NJhk6LEx+neVB
GE5mlXBTAMTNe06jx0GEgOEZBZsJfM97EcJl9EDoHgri0HOwMqpT16hY+R45bGDa
tlId51fhQdaDal3wHtFUnTYROYFq48qIbCwtEaow2sYtXDak7VTzS57gW7rh/y36
VyqLExySyPp5SSfE2SHbcpfPcYoZRdufICu0FhSz6DtA2DrKk95CVsa10guLGPXW
RJfei94utV7qHaKFmGM/xkW0wHJrKBKC8pvWdWXKZ2g6hdoSx3YC2mw8uMh0o6uX
h8IaNt51YU/KiUZ4/MAP6DiJalIt3US3aRzWocDIYxFhgMHpQBMUTh+xyPGqUd7K
L8xQ6fvR8rmdNA7CwULfV2sR9pu4ENnyCVQ7k2AdbURSgvFAV1qLeRuIug3jbeQj
dnOpPF5OUjcFGHTJy6hROwb2EH8lb7gUgHjYCJoYsV5HPGjm+YhHk8YO3VLwFlTI
TiZcI9pcYx6Mcnr1SfCM/nbTNfW/tYt2Yb1bgPPi8uwbS5iBBvVtqBQ0khaJ20v1
n4pmruiFjsiA0i/S2GlHgRm/E6m7XGaCfS2viHFySsp9l1K/TANJc1mOx23NkOeE
78bYjoz0VMladkLGjkHyy8yABBHF31RX6zm3j/n5NDxDboPuWk4VZdo/G6Iq9BXb
VIknCKC1lNGK83HEF6CJnBTviy3vORo7ufVR1xYvwCG/aK2tV5J5kqhruqsuTvb8
xFh6uCDv8d2ntgEKHLVyrVltdbYLJp0TAvFOjEMK23lncjU1kn3RdqEYOBvd/p3D
gqzyIq+57+JCuUFSxW90v3m9JY2JqsJdk7Lth70RjyAxfMa3I+QZGoPqxexQCqzI
ee18oUakqaK9LAS3Q96kEtaEM+HPW9VgdAUuH7MHSdc4xQ8YSp+iJOyj0mn7sqkm
BIh45XgdhUQevsh/PsAAqjE/F6EWvzy5GWrTuM8kyRvYMW9yfQAObbcK2rdefkHc
5mY7b1iIyb4uNp90/Hfs7Jc+uioVEgK8HgJK5WrV2c1KUi0jNlNB5M+FyieKXCq0
3QKbDoxqmUewcQhnKDUmrmVx3USf40FbGJQSdxtvwvuOm3DIkSmZpwjYjx8ZsFad
iehZn/asgDsc1gZdxrd26pbVepkz0IBsBKdBvIoZTI+ea2TgYtbS8totJXM3cmnq
HBRQqm0rnq7siHXpGwPJzjuIQ+7qWo0uQFYJljJFDvaXEEzcdiyxQNo2tPkyb5bp
nVEitck3iB0u3nqnEmPB1i9SpzLsauN0dvqmRncKtl9gprqDdAO+ssGo9VzF9Dq7
VnGa0w8z8cOYPGKhnOPKrUeDBLwqxmGYKDOsYATuYPh1DOtzNH+aAaxdVhLaM+ZU
xrObSmBkh3QkcBQ1DQZTlJh24s/O6OxpgUqvyPqjMAkZV6IHXvu29cLiD9S0bz/I
VZMMY9XEAW2LkM6D+33rRKFSHOkYJnQRVE7fqdUQCrXTXudfSCaADdAMvD0H9bT3
OCV6o9JI36YlENKJe3JCsqGqAEYbOtektjH8eVWgk/69YDK3DIVkUZvudaH5B21P
Fe6J2vjDQTZDmOIkaKw2XxAX3BTqh8w5aif1DeF/+nBPc4tqqALL2jkt8Mlz/j0a
yZos3CI0q/v5ug6FrRD9qmkK/v0zOYDwYSJZRfeZ6yd2qUcy7hsVOVzu92r1bpET
D+L+iCF7lkxW3ej+NJIIGKmeltydvhCClWYISdsx+8VhBHfznmPvZ+e0SeDqIX01
o4mauoBHrNWoNCgpwHFqD7qxjXIbnk2F7/0lk+bZWMUkEIkVWH/j0qJ87wax01D1
JmeYQfpeAdjLBbdZVZlW0bRtojqSL5Ou+QdyowN/YV4Wz5ike9Uzb+k3hIOb0AZH
BDQfjZ38SWFzxGXrLsaiFV+2FRAktQO4/whr0FK1tsqeOFbXYjaqR2I93xLSm+3Z
7sgov287/Xv/U5OdGOivZrxEqi4LIZd9vLriPQ8c20rZyjO4J+Sh+b5IIr+nBdv2
phh1EO4TeDocMrtLg1JNXQSmmQIyrn3+yA9spzAb0yE2yDVBP9waeisLqtisxQBz
X1adGOZz1+cpknAHWV9tbayIAQKZMYfkSnpISaMglx6o0WsFuN/c7J7i+aHnIBeG
OmeYnFnQDd7C7KYpHUpjR9Vq8qvhG9HZfHWBMi0MFsZxZKo6l944xRpeSP44CMnt
woLNwGtSUyH7c9pinVmGCxteN43nyhlPu60NwumRdLxtQl9p2mJKiKlA61CqwJXh
IQNf8zdcEi2bUDCddc3z7WrmEZ4Qe9uiLeMkjnW2W3MrRbYaWcAUvLnzTZ5tzapd
aWn/fuB0vISnVmICJ4u8FvNrso3BaIi7D3cyVMBwjFd9XQK3693evOP+rw4/nikx
haSU6eDDhnN3lG8/cLa1+Gs6BJ2tmzgfEmihYzxzXteZpX2ydVraajII/qewRG8B
vOG3q5wGX4gD9GekHwVRXMXJzb+CvIJp+eKgSrMLlZ0e/OD5Vklc4WSpUKyMlnX4
85xOvFBEwcZy1VJcqZRFcsG7BA7Y9DOoEiUUFqINCtq9dh/bvpgwImG/ENK0cPF+
/6VZzrLRRGX/5BoUouwY7DZtjzDXmh5hDbao2ADFZM0wGbiw82P4hNzo32QP2OzF
GFZdNxzgn98iyT1bCGzAvgS1r4St5/5a7TZotSW7twxfSXiHW1UT/oRI0g4mU9i7
6wyVVmbZWE+4b+ONeLrjnNjSDhRgfXCqgkYMwZBxqhnX45NLbOIIotgPl/g6PAUe
3bRjC6QxOX76OIcsNF6/0B5oCWA1t1kEWaA4/PiyC+wVQnsMRZtuZUC66l1wzLKj
aoIPIs4cU3fNllgUhHWT8Di5puAG/t+v4u8gpsdniufjgLCJuWQiq7j7kP6j481c
aRMOFpdg9HdO41G7krL1XSc4MZ64kPST+813iuIDSJgLEo8WLnuasSr1peIRYRh2
c5L9OQ4ORwit3TlJdhBW+MKAFXJZZsX3xtWEKsv7lN+gcgVfdiDqDWJ+2gMRYNRD
KMH4rv/rZfexhazTnUizV69rC2HJXeAcFcruGK8SIprEDRjjTW7xjRE2hcaaaO+B
bMEdCbxLfkJOY/b3yWzj/yRdvrbZHplfgWg4sh5oMuxSYvjOFtT7J9ma8LkrScn3
WW3JHXRkUyoOhTy0prKfNjNTzUM6T/YRwegi022tlInRQAe6BpGN989yeHFV6UD3
B/J6pAkEuScN4gtG96IIDl+o0nyE2qzt+Z69YvbgC7u3jk/RAllGun7SdyszBYJN
aJN7xwUEErHFltl34FvwOobW7EmQqEAxrRFUZtVMbgzJMtsYZxQjKtpxGZJGy8n2
TUdSFHSFMCOJpSIJVbfGUM1MuTCB4tYL6WUjE++kALJgpAIzlPkGfRgR1dDguUIt
AH4kSfD+hpgYYYN71o0YdATAQ3BRWqNhBBoUQG3ElpSs0j4/hAm9e6zCM9UymXwX
wLl1iYPsjl6a3afWt6l6DWeYNPPaxDN2UsSTj+SIFzooSmLRZCtoiQDVRqDWosD+
U/1mqbgNJzThiSlp5KYS9ywmO5i0xBWG2zFVivVVhL3u6xcnCKFKPGsygEnvVpEB
uBgMpqUoX5O91t/YdJT2mg//xD0By4PYCNWkxMFmuKjB5n8RtHpc2dSPw5GC13nP
A4UD+m0bUfgaM9l4dX5z90pjNLUa1cyoR3m0rINKTdonaQCQ0M1B6yvp7jhgwJk2
/FECFCJo7Q6TsygLiLP9cNm0vh+Ud2B+a+2VBhKG9dd9khkhp10V2VieRgOZszrf
LK24GWfGaSr33LKfP+Fhgshk6snpuam9PcL02IQ+FgVfpcOrwe0rY/TntxHEV5Lv
tlFWcPEQ5DFlX+Mpj58xhp+bZ9QEowqF2cNQUzhoEkDYtg9NfS9uW8DHQrJlxG5x
696CQ/CaTowgYuuHAFymQ9MNemKoHF2Js4xM0Q3QRlhnV/KaLiWVPIU+oWH33oNz
ow7p5YGvCO4F5BasaN9MBD/+JmcPsKyAaHA4eJ5XF9v1t9v13nUQMSTenatMMAZG
LwkSbBZOZZrJpMWj0blYDHvgpUvLU+w621TV9+3s6cSvXTy97qZyWzA74vhL91qE
0QuCpyAj8o3o97VAhUS1XmnSfgdALITCl2FmpEFVggai4E+jNVF1YprVzDGQvZsb
AJ13lhWt0tefURqOYk6zxabGiMc0DBOKsg7pCGZo2RULucrB3kjnOseU8esWmkWM
9C6ebxIIy6QU0PFoS5yV8nJC9vraAapbFqUbDJgFVVr1+22ke/fENoaydIDOp+Py
qusSVmsZqT1a7fMbaAQYoZpEmwpvrRVFgSsjA+AGVliozZJKAKhsS2eRz2TgmCPj
bDZ94rpjuj0asptk8UVjn3/PCLpRTDk0JuGrTWxgoQZmye1KGWAP+X3ZQ5wmOFFe
MhXg9nzLKOoRBjWl51NTfz09vN5tnZ0OW6NdjmyCt1SuSd8cUkhmm/Q/EeuCWPSC
zOTvcz+UPzGEWyAXy/bnX3ZVptNVqEeihNAQe/FEICsL2pWm8eKPBNKLDRN/hfqn
CjBmwZDO1FsRIi4ab6uQslYk9EOc3F5uTFSahzDwVsLDDkcsZ+/vIJcg6EbYfqlE
ffEGeYur3i+iJCXz7at+k1eN0QfHBpm+3FSez6xkzd3ejNA4rHL7w64zLy2widgm
/NT0SqNNomzBwR3P722QDrfi0DER0TU/hzRb/d/MnkVkAxEYEhw9+Qfn9cGS7f0Q
knly6iNvTFF8KA9db/9lRlsz/kLXqMgrDq4k6AxMs3VwcELl6lxE+4a7e5Uc8Gkt
wGo5XID+TsSILwVv+c+8Jt2JwFfN/N4XPWhzFZ9GgaA/iuwH5zLJFyULZNpZ9yQy
ntr03rZY9ssG4lxb5pOReSnft6bRwbMovZ0pJfjPVVE5goZUEsBpBu16tqZiDXDO
7XnycE8zSFqnflke3l/jBj1e0ctqF3/pFJ5pa2uTFlfdjo54ncCPwX+UBaIFAkg3
efe3Ju4GNAFKFQVVWhjr1Ovow4xj9o9jxss6JxfOyF88vPDW/VFRwTs04w8f183l
KVFrELQ0YyLS0+8BUx19ZvdHeAIsKHsIIzlfDyFGfczWilBByYVuW8BLGHEYn0hW
AfDPRqBpjvkWligPgOJg/y0AbAl1nRUlZIBP9EW7rWBLR/W7N38nz3OMlHEYX2yX
2z9C8634GQ5MQllEnD1xXVotJBlkvCn0v/L/pDrUadg1+LkKte64AKMf/L2TOf+n
NpjXpA10/zLRyYLOTVYJZoRc3UulA8B0b6oehhinidPRwmCz5JrG02bF/YjAd2t+
NjU1e5Ql1dGDEC1GCZYHRqlwVBSfvgcUwhm0AmmZZLp6Dv0KqeCKRNVcVq7nNyxQ
sYnUFAsqtZOCCus87SK1fX8Xg+AkL9LImCON1JEM4XIMsgY91zyEMyB+QHuD8set
G4mVeRgBXRa8cQHDmgWYdyGFIdY6KLeTwaj1ztghPhCHv4cTx4qw01rtPV3uYNjT
LmMsx4UNYUBXYjwP81oqJGBaqxsgGAMk3Drzzo7ANZ5814jhqvdSMN8xNaF3ZzmY
I9UqyfDjYEs59NNcDIeFZR5mbkcOWtapi+knluKAaxAng4rQB+knmvfjgdx5oiFC
0ara35ryavJwgDsrAfLS2+1Ark1E0ZcuZlUG7xC3eRIIkLX38FgWi6QFw/W4mMk5
7V8Ea0GYSwaVUebS6ywzrbUVDu9rOsE7wVlUhiYs+FLHoepXo9sy5XmWAaVDLh67
U/v0JJCe+13Iut4p8wi/oAmdzI6+WcBr97PFaxbNFMRLM9t/1HRCN6a+I9MGKf3l
0J2ZHC7sjvexVYjLTSxf/N5JljXxRq8d2qe8uxRxGI4I0NLnrIc1fJS2SWblri0m
/ogsv0CxzSRlp2xDdzLfAr69WGwLwcyQO60fYeyqpdoyoCrFn9JZP7zEGbLeBzXi
nBLa6yvcqh0oOUUjwkAN088GsSSk1C4fdycm4Hqc1MUw9kU2jeDYm8gIzVnpL4/Y
CKZZcdLyVgU6rYrc7u4jUu1f99z3ZPmZ1eQbp0iFKgGkhltu3mStKaRAi1KU81IN
qOgHcGZ5uTl+P3fX12FmJ5jR9SWZ8xH+KiSCwWfjAXhR0AbNpARQFIUSxMfXXrAV
n6xAqtKLMSJDX1XlGPY3e9fBT+RqwGMQIY3JoNIx8MRlFN4iyNe2VUTo+lUf+zBy
bsfnp3QfwDZ+mOdHoYZ7aPPN+iJGbtV7Oc31yUegp1bNNJlNz0x+TZA0LLaW5cLI
R75/MsYpl4zVxKrXpsgrlLeWMS4tW0RqZSccRwbIpOoxe5rJFuNaDU0xyqKOlHjn
/0oS1onkdvoJe2ojeDCPkioYdmAx/4qDd9+28lgWTHEMqbrbktQL1JbO0QjGKovp
J1n8YEaZ3BPb59nrgpF5VDYkhlwpBKQoCjv3IRAXulPpSu0aZrpdJZZvLU2cXdZa
mBE6nUY7fJo3YE97Mb5FyMSq8xd3xCY8ny3htFqejH9ZaM0L+TPotC779ioerKsq
wwZUE8o4ClM5TT8zbbJR+PeLZrKT6EUi32dGvjLQ9DzeT1cuUVVOTNBmu0XIUKfY
15/vgpuCFvfP7Bn4CF+KZjCkjcg9gnl0EDoLdWyrHvImgDzZda8BE+xZhad4L3ER
xONNhjvnOVOnkRD/h0xv83CU9sIZoe9MDxtVR6WijuKaF9PtPVC/vMOakuBnU4DL
qPuA40Mcx1NU/NEugPK/ij0OoMzty4g/n8lPMG7K0eNAe5OdGhbf9tmlkaLHCind
afcEWthvdouxDQZRSETn0TxUEWqFNYCSX6DOdUlSRZROW5P95yIvebGWhdTPJT1Y
whBZ5F/BHYjOArJ54O+U8/zdEnEBtjF7jMVPqm7Ju5oWGKp/oWqx9TPlOBdqLz3z
qu8k0JRbBVZBoo6LWuIKoCuND4NczHXJTB1xZyHobRkKS3UZEf6KntgT+uTCmY2k
8pAerR5fI29ducITU6YcII941Jch38/8hAdHe2ueZ34+KtohplbtLMd2jkYYL+ZT
zJPov4jOmS+4twnDxvhMshet37V4H4BKa3y+Nf5GDrrrI7P8UuBW+LFBZqW6Fsg+
WMYvmzz6h+o9vu0rfwrGe0oLCdGvwOqh21BUEWUgfLTqrPPDX3PjG9wz4+6d2YLE
K8PSMVXxVFIPgW989SpxHCAUnAZlSR5Qq8hQlHsZeXmq8TeW2lKYjqWP8Jn/36Eh
HAjsXHExLhiV2LUF9OFOII57wcKDsSeTr4oHU8ccCQlcUOvL6XvpLPHJD2JcDhii
9k79A/rPhNlcvAu+YoGhEFwh3FMpnCHTKVxvsnayjKfjg1OAkYmFMFnSzg/jXt9c
jdvK783X682OGI7NvIZSBKYstEJjrFiufl5HNex8uBMQ3F/a4buqhDfjIG6g6LfP
WIY/oVHx+RRuccyPAdtF02nLIcLJwEgZuLmsBSw+t+XAnOD4cMcDj8+LKOxRoz/O
vxIWjs33WItRwW7AFKxitR92X8L5OnxKWTZgF+L/i2FQmjtBXqT6Mxn/dIbEzvik
zeohKAL+eLcajFHXFvpxlkl1ckUJeyYFP3nY2gZPty2DPN6eh+ba7TUyLBEsK5kv
L2MBRGf8p55aiwHgE8LRvBUjdKmc0FThxgaGh4abemKugEmgou2+FPhau/POTLoE
+X4F8gdBoq00yUjfsSFX17VZAY1GFUrlOMKvvp6rgkwb7YZ7yEPZwMBjAsiiD+iE
/trRthXTObnSlYLwCkj4O6FrcLAQl4PWfN9+VZmh/ZcAti0ievSK+Nnh0V+/s61W
u//Bf84+b3bFUzBhkvooT+Wxr3bF2QhH4zjlRoaZftETYNQ3+PZkQvI08dzNC3p7
BxU3TYnvubVsfS0RoFH4qw1FJly1nqtN2NMDtq9zK8h+BLsn0M9GK7pAZmCfPNE9
PdWDnolO4xhMGddHn5wxtk+eTBNqL/FDS59/Xi7Jmd2HDDDTOF4RN5EvM5kJw2/0
uzPhB4pLoek/FlPZuFXMYlrPWGAzqijSiCcGzDwNqho8My3Zy66hwiPAvvmSUp1s
Kei056/7wtuCK3nuMpJ1dYUUvrhAJDMamEnT/6KUWT2fQpmc0BYJS4xeL1qv/U9L
8yvq8kvobZ2Q40OUOnv+ssqVLzop/ycrA0J8t/Pb9NdS338+U+KdvOnffZQ6wo4T
Xw4dIYYTqc2cEouLcn3jn0dWBHzFB2LuTojp+e7nf0EtTgZv/ySRt2WFlB1ykf8F
13EvSIcle3l9EBDMBpCHkH1oSzw/RTkIS8tlC8VsXWBysbSTNuRekqSIn4mBmGbD
46cLichNzgBNhq1cupeRo5qPUoWKyYFOxK36j0lKrrpH1BQp7pYFT6o89QUsHt5+
C29dqh2t57vKbl558uyBe3CT4b+gcCh6D9snJQ49FMRUjzgeRifj/vsUbpMk7b1b
3fjfLGS34HIrzuFo45R5rzBFLh17A8mH6DaUmTg37EYcFaHbusFARSI37Q/zTcfF
ozoIOcqqYPUCOLoEgcPZfbyWQy2Vb2mkb445lpAanFbf3bWyo/U1TPnP4pjQTQh7
k5can9OmmTF6I7QVl3BrOfkBy3xsyTT0Hc7fkKnL480HLXT6exCHj6YYLfr8aSpq
6qHQOyNGL/wsprWI/o5nV1KC7EyCESQIRne2KgFvqsI0Jbvxja5518g79vp4uwjx
FkcD6z8Uwn4zzm5LGAylEwY4hYMG5mLYn+0ttVP8/yugMfiqaWkWIVffEK+sIZ6e
EH6uF4Tz1UUw2nBTKxoEWFXxrlglF40BRcjYKLC7gXS7QAJ0jV2pjg/rvssl0+BQ
Tw6AzN0NaDsKwFdVe5d03LVQgMFDcJlHo5/OZ65KPsDVA0okTAdVcHVlrehgMFCx
2DxiO933u3kyiY/8/G+/3uQU6sgFskqN7kiPUB8pKVeKrIa78ai84yCa5SypikwZ
pB9HMBzrKNNsXpzKc8UNKSwmM20kqdhhirLIaq552b6nxP1U6fZLVZZnvwWB8xeK
XbikUTN4e7cxZVO8DTCsPY/2Bz54N5KiQAG0etVyrpVCabuaDh8Xdnqb1dQgpsQW
GQOAPPhPpE7o9zCciTq0xxux4HFMmBzy6wWB8CvHS8Ub0j1hZ1Mlynw1TeGNvOTI
4EQfAiFJ0BMo4xSPif3vVT0V7oS0qKkVh+UGzFUK5T2vTv6HLswfUXS0ACkWKsfd
LGm8tnVPVjMogzXItKZx+wHHq2JtpWNXRezgncm8pqT2zIvO1cqOcJF109qPHyF1
LUoY+zmnhsvM7fah15865eaV+504hMwMMPpeLcrDkxBeVNvwqvymAy9nVNaVHdk2
zyUL8zUuRjIzj02ztglXqDZNvVMaB4Kng9+W7Gb2D1V5mNj3iJXw1D/U/BlHW5PE
vWYXC6MYwwRYUVSqGA0kc+oGaDYkSGGpXqPDmrbsuqFjvSt4Xr0/TsX0k2STz1IK
3HK96Gj4KvUMv4DPcTl5J86NGK4RNtMflzrFqj2e+OJbvhZPMoatfuceoJy4xLTl
Sziio9Fs7RwcJ3a7VEUSfRiTmN3tdiayX2vCmMNGcIy/WeSMNeBwbGpbaeWC5Z/V
oPNUuth84dHwTLy2cB8ojNfYKil7xFkLdUiMv1obanLM1K/EicvxCu6fL1wPsqNN
g4630DRRyfHsVX46c1XxUIdp3XIfh0bga7yVFR+VN6w8V/fOyRqpMMjNLnD50u8j
VqgptVdqnMJJdUFmI8hqmdLK1ILVl0utCrAQrHj4zsQrIL2iuhmKktjE4qtHegby
1Ydty9bjHHb0I5VBKmXvx8p4PNHgn187RYQJI3MZFzsu+TvtmLhN9rj9GxE4z6rs
AVCo2f9hvjuDYVapjxK1oBPRQuvQj4mMKz+jEUgj14jH+9rT4CpM+PL/bta1yy4j
0gDYXeqkP/05EDdQ7eeLQfZbNMa9J40uhjTAUzPJxG6WI2/oT/0KezFkifJHfDOM
MU2Vtgjut+xT+ib6/kdS2z2QPXlSy9rki8rW2lhLXnXpMhOb1LqFAMvnVKp/jhzi
T63CE0298FC/sFKU/nIniidoovgo2vY78jwBHOE8FVTisXVvCQG2VegKpexmgePi
YwH/S6nCZ7m+h0B/0ARXMjxBo/8p5g/nF+GPwVWtA2XUSRAB1/O3EdxwK6hF57Bv
fdAweIC8K67h/rVQ8Da4zl48y7JRixZQYKwScdeifFk9JhWFSG54y6vnhbU0nODI
tfo9uTAtA9qjw3c63afC9HtE9kiX+9E6vFmWAVZsAmgDqAYMxqGJuQWaQBYHMsD5
VpeNGAkZxiApX+itXF3kO7xVE1p69MYfhkGn+xbzTatB88vwFGsSUeZnB4Mh92mM
lGYjT6sXxL+aNqTVMaecWrhWetzSmmf7CvPRuAcJP+377ofacj9KxDcArU3Cp1Bd
KTKuQ6v2U9DlvIbmbPbe0Ge2ar7KLdEMwTBUV0kDtA/AX0XQuogZTcWvjVbsJ1cc
8DE6SOAOpaSSxjTslOY77kQAO6a8EobhacfEFioF5ZbFOSZZSht+X8zWJ+9hJXw/
RVQWZDQMco8xE9z4lyS1tpBx/NImlNmp7UWmjIxFBTka9KYZ1tnKwZyTzW0lYuBA
Xpyb1zQ5xmqfiTIssEvjiBTcH9Xlh6ZyviqHuE5qeGK+n55kigavafKQ19fxdVQR
VbPLQqLvgcoZ3NvS2EzObsH8Oj2XcWyZbzrqzsN7aFqmMu3Kprmnk3CTaV7PC+LG
RB3ESQ/lKuqdDOiuUhq7KfWTndqDei9EBNho/JurZqgS4kp0/BV9joz9bzbUdE/m
sMDmgprOcaZC7l1ySUIBLsCe8mUzV+/14iQEKG1AgA7raGpCvgH+9eOdwULNleNL
80GXtCxlOa7ckVhllRwiVXYOiB4m19O9BL9b5wKfPnIZj4XWt5J8QGjZJy7E87LF
RmVGwnjNdEOrNbXBtu2W5viYpfSbbGGvUuj4O0DwHwN+1aremwYGSKPEprD/Wyyt
AF3xQ4MdhNBR2/KYad9TP4G+suyUp64cOGrNh+8QyCWDTuMisUq+17aFdjWkOeU/
oK/gyQ633Yu+at7+094a1XJgxBG/VRb4lvEqlfm+oVuzcMbtdH36xDgL1I5RaHSz
WHuJyT+SC2iHm+qJQ7rgH2v7biF4eYmAtlRshjUs4fr68lY28CSN2+HuKOyvvaux
V6W2tu5jl1xiKoG3IHBea++YJP7QwTe+8wd+zKmW+muagJOi6WE+qjUHBko24v89
mc57dAAKQURGSRxE0R4MGtukxlKVw4BOHTt8gspe5VX/WjKqFjcvFhATxILknbVh
62kA1rvjHrVBdOmndIdrs3rpN1iJeVhS9Ud4lSSQuocXOc0V25CnjYJ8bf/UG5wz
E6M9mrl9chz+Rei9mpbh/3Gy7ZZohHbw46BbxlgcL9YLTGOg8YiI30Ie6GxAMmSt
qQP11NWiu3eEKP0IA+C0L4bAQ+CdeG2o/W6woXa1QjzQBhZAQ4YkkQ6GQlzLQo21
zLCCMsbdjU47aCEQVANBwKRYnv4TgBNo4rkOME+mp76Jo9N7kRBlitwF+REGFEbK
gsMG4inKpzsIVS4v3mebcXj7ClqtHCHYW4o8uuJYuWYZem3+mhUkKbPKzNuFHIXB
syfdKsw6glwze3qxUw9dxfvcKI/XXNUDZDi6C7W6kKap+WHlOi3Ill1r7e5HpFFy
RFl++IrUIaTJDrJuLeXF/vLqyRQb2v9JssDoQvmYL2aJAHZMuJKHLz83H31g081M
kOUNW2BLBoX7Ya/oXCwvxpiAo+pIBRYmcPNXq3Ypd6jq7hVGoRzDjHqQkdrTKKtC
aBk4AjOKQHuZE0DMiQm+KnabpAVpgHYcKiU9zb4RtODOTehDXz7403j5E4Qn2Ekr
KxO9vOt8TNg1S/DPYmJ0an0CYcJfDl26YRLsG1MyfAWdPK68tMnnWjOXNuLD6ivq
9scJ7GwQtg1aCLJJJOHXa2owakBoXde97AtOusP2aoYrollUpfN65Qmw+UID/aRc
dQoRiBDNDBypNDO+k81VaXnzJoaYb4AEkwSIrNTvC2IYIK72d6NMHS2OQPdEfOl4
cBpZ72CGOPMZTtO2QaUb867S9x8Lx0tALTkY8x6tgarzXHFXxlZNGtFFqXVyV1XJ
LocBbLQ0Q6Bdl0ctIl66e+xiEhpIFbCkaEiC+s9JkDFGZgroR726CU7/0G6O2nJK
YBQC/LnfPU4E2hUxjYEanJCsFLm8ljc9egSwbXqLJa72IBA3vzK8r+p3CNRlZpSu
Qx38reHXVtMrZIgU19WgLIC13rjgkVPRVD94hWm/LPOWNufSDS4Xb8tR3ImNLtMk
RlyY6cS0YbnCNkPnOfbKUJHxM+l9eM/WjEeS8xYexmb7ZkJDaRdJAyTOe+EBgHEA
Xz/57ds4bbaJE3oBzvwlPb/tw8YpT0saQW2dj3d20TLKHKmbojPmOmhaVKuPlIw4
BThqKHZLJb4hnrrVrDCCWe0Io6fBxkIWqA5TS1ZV58ib7bmkI3XtXMTHDt2gMO7x
j8ZR2K0cjRMZyNr3dql81K453VDY/eC7hynfyNC7X2IET2uEhBVLXCNSDhs5xcOF
gKpSb8+JKk3M1zFuHNLTuyrGAYSWbHoK/6GcjUjbMsMSQ6NkFAW0Fco/jnsPudEj
QTPgikTgj4M/eEdH9C/BzXGbiZ/o/IUUcKU1b6eo4fWnLAjEjcGu59uoHoy3r/Qf
yEkdXu4DaOuJW/qnI7JY1RbJEaS1fFXnxu9yL4tDaWqp+hYCLAXBqoOrzcxCcvky
X/OUUToLvK1AkmNQI+7OdQo1kcMkbXfys9TLOnz4GKwq3LsnwdfPktfwn7zvzBP5
N4fiXBmUg70f2zAsbwMm8WsdACLDh/IKDHAGTCASggTRGeLZsMyZUSBFKLhRQ5kJ
Qy84LRpp930lB5Ned4FkualPvZ3j+EngSSEzBnKMyfUCDrWL2I1xbuIcZsHsdDwE
Lb/1n+kIXnYH49i0fYNYTPpXNWgOuJulzNLRwCBjulfX32AbO3XyidHcNjFj2rql
IAMZBJmdBJy2Fn10wmGSVaLpteXGslelQxq5snOYG/kc69DNRDRcPzKstYLaxzmF
Ka+RXiTT8CSzm3/yDZCCwaK14TkF8BMb8PBOmeLX19zT5j6zZBz4Mg7LhN2m5BH7
T+gBYrfipM2mNDYBghYB9zU4/Rhp2oNx5Dob2oK/ZCT9yczKFbNnzXZAU6GHndwH
XjPrETqTGLdFdhR23AcGJGBNo3tiEVlzsIgsp1B6TsRQsM2MY1mm9paoClQlCstF
4M4dwsv5j8axoIlP5Aru07rryrZCKNhV6fwTw5+M6hmEdMaVA4+jjHCg/ydYrT+j
lqAYWKK9KdYtOJ4Nc/9aS/VlgDp5zTqYsP9M9ne/Lu3nfajZwtTR1jVcxpV9ea3b
rn6TUBPeTAbxJrE/0KP3TVyjcLG8WKBPTo3eq5LGjcsbuoBe1XueuoTIuB/aJBmv
l77P34VAknHW9h2rEGUDgv0RDFjqfy4o6h40ytWTTyReWQNBkc2vJNABIwhTSv8J
xB96qWP2DHRBwfZr7KwfwngIhK/zTJwn7oHGiw0oQa6LktDJ/rKefvpE0NedRFVH
dlAJoz4r/xNZA4syfzFvzbZIXhLKoJ+vbn3yK7Tz4JLos9wYdkqa+DZGTCbYa/a0
Nboz38I4Ixmhu6l6yHKTzmyaYdkUVDkki/YW1StV1Kg1HzrnhmyU2ZsQsND/0pAv
B4+4BFDg7GHUKmUZogvqqxv7Th286Z8nFFJckDik96UkISnQ5RTjr7sD85ob3HG5
xSpTvVOwXiP5rmJpqXM2u0w8d4bvUCFuojxRbPoY8MpaMhljuzpGoimSWdzYCOtk
kkylApkg19HarJ9T359q5n1inW8zWi7+6aq2+5JW6Xf0p13FkYZ435FsP4vx8JB+
wNBG2ldpxFCo0BKtYTXOQG+7yh1wqprQajxC4MV3ivCOF1t9iy8I5Zrqg+/zlqQv
KU5h74YWZPVQ9mPEuJWIgiY8VFF0aJUEF/KrSw/ZfXosVRivsh3+n2Q7N/W3breE
MN1AJ6q5me2pWZlbD53X0sfGT0lIKxhILagY1Ipn6f7vJSH89Dq+pAP0MOm2stIq
LvXve8vErfGp2P4OJOSqnFCjBVW+ACCirS7p5txzfg3YPXUjUIAd0e1P5+My5CRS
RYQczqIN9UvgiPeLevJewwnWMXevtw5bcbPrzxIGtYvueVuaZJe3kldtYqCKLC4U
AHvZ1vMWEJZpHrYGya2GDTHyuQaNGfQJPky+4CdAVF3V4g/EylmRoKYLfBedRh1U
2HQyesx3DgDi8ydSYe6LNXFrgFrwOK4mbxgV12F3R0VPNA1J4PrsLltcRbpXyGLg
N6vF3LXCgLYFlWguTwyolVvipd/nk8Ykx+PbctVJOBpPD+qqDVj1MbK/x3qtYRIF
ic2ylqq7l7eHtOf1tWC7J6QtYFIGJuYBx+fSK4y3kesU0+kKzQRvTiLHA1teMQJg
VjM/RMk18GN/sPGxwTjUH0bQGQKj6k+rn8uhe+jZ09QlEwBhcIga4TEDVd7k4o2m
0nPY6t6TlfXx4qeiu+wRUxCZx444efudMZ5QNhkZzOquYX3RvnmAEdaIdrS/M/6G
NVee8uEhLgaAKoA4QmUs6SP/uR4ejQeUe7PSm9ob0b9ugVjEK9yRyeaTfAl+3PN3
SF3Hb4tWVBhIOWdoxEYVOmZ3xRpSOQCULe0hJBdQcFU8InlSKa3oH8RPf1CB0anw
nYPJ+ZNIYQ7wDrT4qN2gCJsxFe1LugkufG+8GfZeof4iy+6Zhi6ad/y1DfkZFqKI
obZyKCv4Zy15uKTFBc5JRE+2hA0GVGkNbOl97hJVQgzFNPu1gv+JD1gRKbqLp7aK
9spZo4/KYKHCCMS7rHyYDy4JUpymuHmTvTGwPCi+ulHGNTndtCSYthDKVqaXU4VF
aWspc8u3woqTAyeFY68/hhYAM2HftNvBGLyoQtAlGDHBSkNOlY3GEPv+28nu/24H
nzms4mLMBZd6QaMy/JpP6tI9bjO5IYEOjufmXCj/stgLxC+SQPDakBT1XrB62jX9
m4yag9WMkela5xSqV5xXHRU7SnPwr99VX9bfDezXApJKo/vpd8n2dEi+Vz49si5Q
kTOklcuec7L1tIJ2rVxR42P6qzSl3bDFGERC8akHEfqPLJMwOcry5+yzOo0TbRfO
S3FIV9jOQ9L9DWATNZ5DiiPAqHQlGwvnlUB5h4ycUn3evNGJ2ukfHoFe5tgoL0SU
ogwl+TY7DAYLikPY3UPvhQAIaV/FGtWWoOY7h8HQ/jpg1eNrAFRneCTxCFfGI8Ns
IFGLsjwUaWVfiLA8oVIsZKIbvs4Hc+MeOfHBBgY2SwDr3UskBVSBulGIwzZbDkZE
GS9vJWlmFIGuagYnHShDOoNpSvkQFuCIOJm46+PS1OjpL/p/07vJPD8AIKOeTKfV
H2WRSxdPZfEL6D/WQo8h/YhGiDPBPdMX1tB59+SwvYYpmTZVDnnNODg0F/oXmn2I
vQj7c24hydhmrS6elnxgo3ZT6TKY4DrNpr1Jn0MdI+ssKboEnRY8ehU/uC9XqbRc
lQBiuu/lcGd8ay4aKdsJpNgJQCzS3x2IXSmDkwFJDAXb5GBa0SCT2lEa70bwu10A
t4pc2u40y4Vg0TAJpi5R7ZJNZjX7qf9Dbu/O+qGC3ejLFPysL1MCJerF/487kcD1
/wSB/ZxDTmXrdOaSmc3Z9ppa0iIBkxsYbQzWOa1corb5sADyrVVXDhuXvTTl3tNA
niok1YlmQbTkJgDQ3i1LZlGgh1Y6XJdXLzrCxO13KuguH0FxTp17ccLn4Noa94+Q
XS1nUP+VwdkCPABXt2u7eM6wDMbY9SzZDMhefw/vIPSWRQ8rNyY+uiSDquKjtblU
chDG7DWKlKzHuTNsSEnKk8TQbpVzOrBaM3guXcMHCgj9MAJG54O8T2/r3o71T5Fz
P1vvAtOYNLBeCsExHVGIQRzR60J1s6FEyaYeZ7lOWmLn/bRKlc0M4HJWQWu14Bvy
CsX7onL8rl+HvQC6mhGpJ6IrksrgV05SsgDKNAHh1FrFBmL6JdZt3AWmTsCBBu+b
bJn5OicNLpUSE4hghM/MPG2y+AUXpmU1HwSQanPtwtfYtIbrlEBiPvq4ds4zDsoF
gLd8yRssBz3ONr4oHlb6HAzZ9cgj8KGJfSrZ0Hg8o5klgqbCmMi+f99/KXicWmUx
xkcIr4tk2mmKWRio31uE6o/Te5kMLjxNHvMCfIr11p0JTfpIfuCISvQm6Ig3LHrA
ryfzOa27Jl+2hmXCJdsq7S8sSLe7yWPrnWYxbdvBZNoeDkRervoj0U5qQDubZf7Y
JCwJnAuRVx3+sCpspO3n12aAh+843k37gkakRnZaTJz1Xq3jST0baA3Tv5hriJSL
bwnpqgz+/OYI9ic+YoYaL5rbq6K+4sGWMMWqTsR8BERawn5ypVxmaTCb4/pc7A2E
FFLvKl8DiR1gEQUwlrWb/Edvb/7imaYQabTQO9om13SuyKqKhMPyA4CF8slzBKHY
xS4zQkLDoJcmDDGk1aqB8IAOGTxVdDfGomHncM6r2GYC+B2lZm/uq3yDdVPRWZxT
/KLYa55BUFbNIHxi0fdG8eWZIIXFw9AKRsMgenDnKPO3CcGhnKuLLqK/kQt6ChyC
uR7Hz47mX+6ScEgGbttjlRQ/3/66/Bxw9Qk08c8HiiUAjFmAE67+lBcTwgHBqTHx
ec3ZKoB/ZyYuaI1MOgrTizmgm6KFx6FNQQjLPYGWJQm9/Q3BaUyBUBk4y6uMYLLu
n0+19oatYpGgrTJ5oC46e5LWa/fYh/r2lwFkjTgJOZAL1mA3lLlTfsHfMtEnq9aP
AgbBGEy39w1hpB3TdoCMPaBjCN6AaEi2RzPfTja45x1vbXJuk2jEY3IfpdNULjPG
eZm3Q87Mb9FrYdCO6sD8bLegfixHWQpSUTXFhL98UJqBn/h0qe+JRwZYl99OJ/Mo
DNxm4SA7FOigFyde4sTArp3Rpg4MxwHreEBRbnHP4s1rstI5T+YkXgCIJnWUIMlP
wR/ZD+Y0q/3E7zRQuWHyv7H3KNraEPVwdFlMhm06jhd61U1r6qwpe5j/jvaaC/nV
wKDeLh8tQYXTSTsSxCcZUW/jrRlX1p7OioVUdtPa5XxOYs4Nw/wDj74FFVAMIYBh
+k6oa/YCojBVzCpFfSXzqUkuBZ0BxJMNUCwTxic6KU29YtuT0fsqjl275cOt3mFi
1Dl2ff8WdzxJ2qMa66PIODLajYx6cQLw2VozSMVemAHKE3JVsTmH2Okm2ctBlOOj
MlDMvf+rI9YXt4fStirR+EwKHzlck0xmAtKliw+JjdgPKNAsASWx63Bn4+hp4QhK
bYGghncqzK/Vau9xYjCfdouAtQajjwLPuY6/ohg791Z0A0bL8Z8fk7xi3XPc1K4h
wciiYIHHyC2ytfSak6BSI6zKInlp1WPp9jdwWodNlLVCy05e5rm5+BQsJZ8DbaRU
lc3ORFfVoFxJVGqr16Yd8A7FgzyxtqMdh0mXjW1DLZujo2BAJlAUR0S965FeTJVj
DyTDKoHs9iRn71Ug1JVkWNEU5RJsqlimwn865S8XC43oAgYIWI0WTNh5gjisj2sy
v5g8wK60tjaCG8amEQTZ9+UYeYcAs6K1NavpwxaQeanb6H7KzktcGnZiiTX8xGqz
dxpfFEWYgUn8qTMyc2gvFqDdeU1jtSlZcZ++W2RwtjxBAepgdAVr5PF3SNA3AXz7
5foXnn8nOw4bNLlBfCM9adOTCCb0K5yh0bjPrBEwIVKBWERvlO2BFIYeyPCzwnXu
4pK819rG3MXTBRgDuLPV0OFznHssZ2RCxD7Vw3CRIDAJfdR/S0eZjmF9cAKHTv1j
NXvDEHAWm/MKcKSlhqfkGn6U+rtGiCJ1UGJ71Ib/rwAdlqKuQR4ysRV9armARp1z
D8UxrOrUWRk717GuGog/xocsTfEDDVp1rVRp+yWlfNIvH8115qNjN5+rgzTiWibL
Z6kM5jLXJKstC7dm39sj8uX6SqiY0nDbt0pGzeMug18PR4YwFPLCINDiCDtOa2IW
jhEML1q0r5vOmqNyO04HWiZ6izLZE9sVqS1M4BcQSqnTf6bAqHYRJi0tOxbgN5i/
p4EZBjSOFBqH7jYN114PFe/D368bIfO/cGIDNuKLI1Nipjw1rbyBdH2razz5iGNE
5LatKIUY7O8+vTejWMdkGa5rUyptgMVU6dEHRKR6cR7m8AYBfEW4B/O7hLgXZpYd
u05vHv11Y+Tk2DRB0dGN8obwlI2H6b6BIo/hvS3tzTJB6z408vj0n2JJoimmw7hA
j2pY5yhzBju1Hiw8mmCYFJm5iPrad3usAtcGFqnsmizln80EsDOMELvNCRKH82it
/tB3wRaMQkUhqoAktE4CeEE6fyF39LsKFyKDm0A3jgqD6ediqh/F/lbX2AKdrlEj
lo4kB7Fss+hZK4FQ31SLBAsQpzm5AVGFmQTLjvvMkMgp/RI5iFAhJOxyNU0V/916
Zyhy5MlP2F4mLtYUIfRafKytUdOzPJoQA8bLYRv6mBJkCZtQPfcOhLZRR/wcXMwB
U2FWIYyKZi3f8HVfKjNpdEokUG02LhvinX/pdKo/83Y2bala4LIoO7cdSg5KXLQi
uMX74XtNwfoBfRL6jlEed3z5M7ylG10uIZd45iE7T/DvvmDjKhJQ++uNBoIJLSxh
cPRHzoTus2wZbMgYXQ9LzzVQ77dhaokZ5i2opcwhQFf8le19I1P+u8XMQpZTHHcv
9gUNnDOeFF8J+ldgF7y9lex7l8r8vedOMGjcaJc7XIBEnZl/T+pAgwZLX1f0MQN3
DYmeh/XKjmVUpT/M6sgWgrfBmwwdwE1ROIcsnvbxKdOkWc9UfYYbqPpO7AxHJD6K
fVWAP9ydfWFidzpyZZZqipsg/GBhpX9apr8Shz+ZjhI2nkc4UiX4DB0FvnosChKz
Yd/S3HBSI8Ce3CPHZO1GOqgKB8mVn09IxdqJ0436OYfE4zhjyA8f6s1I69/Ym4CE
WfrYOu2mizXyEy7IhLKLdI6GhK8sv34eHDIYcV45vo9PDs2HET2evEUAnbPSqAuj
IjiA3IMcTVBnUn9m5mREpQaeqxl9pOa9TclyEmGBrjIr/fMwf6j5eoGnQngOpNTv
IaqKtEwkIhwWRdP6n1L3sEYMOrbZ4EmYBaoUzZbJGS5dN4sxp2ScupwWhxfNW5Be
HywyhiIv77ZBCA6G8sEbnngSUK3HmhdrpM1nCTkVTryaHQNiFn1OgHsS1GKFAP7q
qIZni5XvdT9pzm1r4IC/E3GT922ajF1FnduLdHgdEzq5yNYD2f1b4UHAvjPiDLe9
ShzcXiv2D/trgr400ZVZwLjWzt0Slynwazfq2zpMZPgGB65InGRQXdHKE4KL7tbE
vXw3iFzOPSS2nqF1Ch47/B9qF4b2LpTVZwEmcWp4wNzvgRrTsWBQAU/5yzIMp094
/kEWnZoNtrFIveQOKpX6s8uSUC1TdY6dFRRJfZHK9oN/DhxpOxASidlAKYNrfAF4
E+ezKoMHilUWwASxOcZY1Bo/CSIUElnGydp1zL1nGZzlIHkZdmGAQgTE++GpAFyQ
OfaVuNwsEtQMOJ+z4nWXzL4hZrC6iJ6l8Ia+SdP0bIjEw0fC09P/QsPCMJEwJuVw
LMn0bWI97XXebEBqenqqWYS/qYMe+s4+84S99YmHUEujsS25AkOANoVV1oAUlI0E
wpGGZSYVZ3xfgXn0yBsldcLvTU4LKRG325OIn2VSDCmtyNJkGxZcY1l2WtRaznl3
Ws2BvCUtGaCfYGdQFqJOMe2LzP5o+DNjRAb3YjuNRj56MQ9Nvg/SexsVZY5VE5Xa
WCjzJDzxtR1Bn4G2HMkCzat2497rXvfeZAPUVfnDAH5XnLTMmX6V8EP3liZlLT7A
VAs9ATKpDgahcYsU+jOYoDEfTPdc5k0BjGBIHY/hVofaKZVwkDr9F2Q/8v+Jp+9i
P+E42bx4GbHGi0uKCZatWscGclmaQPQczT/z0mfiLFsg6gKqKjXbMhQV6hFZa9Qb
rF7Mf6G5owAg1AUWKKumSJGbdozzlPLD3Jd0/ny0H1ojDlkW4ECmVB6PEexcK/hA
2uF8XFT14vA6I4u9ek7vwdCMnvELEhIHBKtpYuFjBQkGQrA1eD4re06MXbKgePI1
ICMwWoNH43Q21+1lMiF+8CkmANjSV6IPzAwQUqClt76VriOeYUuJRtJ+mLKHCxS2
mf/ajCMQbKmesGZI9UgUT9f9QCxXYT2ITTznsmD50vudIR0lkwI9nsNRsx5IO8ac
sLtboVRDrlqJvbv0eu0giz1jKViSSSpTro0qyEIMWt6LkSVRTZl0NOciuSh4NF77
oPnmb5bq/PzxZYiPwuDWg8qSW+bV2pDeer8zA2s1cIAYSCDqC3dJib0pSa/srbdM
Z3TTOFdrwekrtet/Uphp0OpTKhKmUIInwVi2BWmGB1XpGKtjLeY3iMJfHb7CSjx1
42PjMPPL+3eFopqA2pxhefp3/ID/MQjmM5n2DgCpioPY9TtvaitGcz99J9LKAbwl
+uetmoif69onWWR1KQE8ujLC4aoMGmNIcbl45oMN4yGdsTWUcbNl3pIg2djoRatU
VEOd9JqXPNlHYL+3q96ked89zRTcvqtOuyZ4eGd+HoobpriWjQH4hXarzEmYn+tl
MiGwEGn5wY86KcvZltz/X2AQNCf4pecgdRvO9XHV2xXV0lPFwMppIbP+XEHtcrr5
J4nOplsrKlYvNvyuHJ1B1sLWtjN8wihPeK8Pml5Cms5AH/NAQxNrUL3BRfBv3BAL
2Z3w9f9ylt0VgOk5vPyQvPP+fBP6kxOAHJY0wB+6uR3QpSMyXJjZL/Ird3epIdFP
L2vKLkOFm39ILCYq08qOSd1knhouxmTx/ClggQAcnytThDxVlRtuoh4l3fBh/I5z
uNzqNm+Ey2R9RErihmXDZ/oAicDFqQ7JwYcWsrzO+R8Ovn3JMn3wdL/27mV797qu
Tj4rcn1CdateUD1uT+YBflm67EjT3jTVq1+IT4oL0UV7pa0F0HWABNrNd8kPh/mk
G3t+e5NBN6pclE5LRG08ybKTq9HV8nwQaaurPTHtR2kvig4XSWvD4C+LDPA6j4ja
CKMr4MhLdJ1nKI9IkE3OwxU7Iww5I0fsh8ZYXkMDCHwuMQkXtqB5x4KL09pvHEKe
KYOZTGzl0u0u1eqDPcX6itUBRNdAlSghjhkNP/29jabLq9U7nbn9ifzDWsJQoyaa
4/6dkjoVcq0Ub96WH15pQdAN6F1FZLiYlKwCmaKtFVC+AUSl8fSN5SGhFZYClrWl
8jOLPCacg9Aajv1VZtEQOqfYqWGYGzgo3WjZv2L/kj93YMyOsv+jqaQLmmftL9ZD
G/3MfitvfWcVyTSRO4xlVOi/Rui9bUUSiyztKK91Dz9wfrHo1ZDWG09LVp6sqqXM
RA9VYqfZlq4nfy0ddeBgkFLuaMQF1aqnS1c6+eZ8Ih7MdhYMiTRnkc3CHcRQXuWn
qvABy/2+01BGy3IKsPjgyERAgnr/ewu4pPKxHWZ7ZGJwzFjBaKt9vRFU+aT6B2Dd
Ib9EOfNIggq85HIFwR6hkP7B8xB4srWeAnWe/7Gl8caYlSCrR76TheqRpVzvATbi
OWjEMIklfHj3Hs8cQ5GXlxKr12fyx+BHRJftv6pN/J03JJkIb4y2S9lrA2MDBade
SxeNw77BRW8t94QWUBqq1SOHN0sc2D6ImycUwICWTvqMJBCvPsvpk/hiLTeHgRdc
GSoVjo7UKYDgBXM32UAkdZDnmBKfA9lySskqoapqOhwGIo1K/2pWshbfK6jPbEVf
Zw3AxipXnYysRWiwDij59fS+w+8c4jmwg4Z/EpRZ4D0Q4TS5MDR4N4Bzb9t1Jg04
8nRYCfqG6QbNBdPatmCkPViWHr2Yi+iF+axk5kBOzmvi1mgKR9xwFdsRYPS2cNxj
iw5QVwdO0sL2TKfBretUWb6CuAWxbdlsNYXbY8FmWCHHYaaFKu/N3lvtHMUPgjUH
3w7cfYMLc3XcZRP7DSwYzIPN5dCG+SxJXiE2Og9xVsToKA1TYQLgfqdl4D7Julq4
VMu62BG2KioMwmd6QpQF/OoQm5frjrilD+/rCIxtsgUJneFYmFfRc1Akdq7I2I6Y
4w1fJVI42C8p0ygSISTR7w5rArrG2rgMcJQj9zjMUYfs6TfHYwe/t27I0bLuAV8O
u7dw4qDe8vff8qTRJDSDAZh+QubA6yMfhXA4r4BoFkUtrKp1qltW1cWb6L/klXHt
bZABmm0Xvc0rm9Q6CbQpmUABjPVX9Kb6tAi7Ds4jU8cFQan055p9XfmCja8wnyym
yCyiC4TkUp1V6COhi4sg+GAdS2G3WcnNGzzTJlRlNlMSAI2ZwTV+AHBUoSBZnm5r
K/ecD8uSG/xsu7TYKz3938CIV9aN5VlL+L84tVRx3X8xG/YWA49AKhsM2kf9tMaN
Z7uuDBdvWl+1TAPT7IsFViZHUlJvpEksUHNHcKbnGZZqr3ijq0KYdSsj2kYfn1nP
YqpZZ/MmGGmiXgGNSNtHexAWHOzMrBmpqmuFN4YomQu6G/rjq26WplZLcuNhPPcm
oPXPY7sRbo93xig2g4k1Yz/tNfhTNdK8YyZkrh4HvGXrUTJKT+bB/UIwyNLExISS
34OnbK+v/gXVypydt4wF+l/sMyprF5RX3Elsw1/pNbrSHZ+3tUy+Dw74Ge86FeAr
lZADotU8oqqHQpgnKbVm6bojjnDCv6+JMOe3cAzBTS+Yb7hFYEg8ucWg+rb+9ubC
G6R8yTvJVIED7pLtOr51DspMok883dBsbkD3UWCubGoV4QJJ7mWbtu28Pa/s3G1k
IEsaurUVX61CTIjrjjP5VQCwJXezSFwE60UbkA2i8tai3ihEHJIHc/5zXo7vPlPY
5wthm5PGqrIVHrIXH7+oPorUgwWY2msbU5lizTWMJ/KqU85eFVGkHH5NXKrcVY0R
peOIPgD/KAeJ/8ms0nKpkAc1sfTHvnuM0Tyi9A96qtlRacSzR6Z9vtAbYa0n7wWT
UXspjI/d4QCbsbG/fS2YkDSBk/ivw2b67OZqtbVzMkjXa38LNInieQ9EcME9aIaq
3nhNbAG4fd5cExkn03iV6FIse+eXwjcBHu9IuUNZXYvBppFV+KorSfpkFYqFKw9v
IOGqWtUXE8JY4HhcGd+AhXPgE2REcODNCX669+kqG4OKewhzKsEU7CTWyjJxxXhW
xKYcvHg7Graju7Y80YQcK++G08iqZYQEoQf7bdp31X0FcYsz+z7ciJEKtjplZcsE
6snCTJki02yEoPVOB1a3WSQWGqllofcT5HAPOfsiH67MVGyLfEahVma3O2dn1fEh
mldfCt/rOmfp7GxoEjM4T9pPNAnAID2bxHk/wjgBr5JPNsYt40z0cM7tJ3s74KZc
YUIOlb8HZYkvVronQx/KfoBgCEL6l44ywzn9QvGG1Wl9FdjlPId50kHhCvdE4p9o
8QyDkToDfUkjQIe4SVJH9/dcrSs6TcKA/yssjTljBTJPTJ9ov8wVSJtRzsNNHb/L
5NmWxBcSZv3pWYCtTb/tvyJ4o4hwXkBiOlqX0DBjRNPUCRxynk5MUWXt8UkDyyho
6kZQldK0mFlhiL+VAcgh3H3ItPfJowt/g0ww9PeFKmYmg5Tu6fOmVpVmXz7zJxrr
tCcre992O2XsKK5xhiBbIsWHj2yPQN4BkhuKzxyYf/bE36TPTu17MkBfR/USSDRs
qDSN/mAlApZKzOvUfenisz0kxksS+7seW3t5jSjheYJ7EPCsrjqHDZzfCNhrFC8H
kNqREUib2jlZSKL0YSqn+QwjkVB0xU7vvNlFdvrjFNZZA6DgKSZw1T0S5DbV9394
S6ab696HyIeTPvHmBOJTq3nydYdvB602ywghJ6CttLo4hXsl6R+5VEnpt4jlI3u3
S119hXnD3i2CzoFW5wbmoYtMhz/mANRZKKxPnDCPZOPcVKRJ7tak0QfQPJr5SvQ2
f+3dNZh5SWGPg0/2QiNtOSKZ0bQE5aGqRf5mPdM4MZ+NkW3Sia7Koh7/SszbZKwy
8hL5zebkRM9evm/tcMznR6eHzCK/ZbZyy1vuZ8Q+yHrhL/IB8aFgEqme+qBCiSKe
om4gnczDWwIV1oFh67Yrj0CwoJBwa1QP9lbmOMQdIHWLWnpod50Gie0No9AT9A8k
v2w2sK7UjQlFwbzng7l9FhMY/rCL1F2GHS9jFj04yu6n/emICCwPjaSFPPBOvosj
h3AigSXdTJuO9TdS3q9dRzTuE1No3FmlMnvLGPV799FLC7CFH9XA3dyas1rVsc4h
Nn0PN7JBWJR/8mt01n92fb/E7SlPtkadF7kxD63OXyiH3gh0lbgL9CnC9COmaZ+w
whpi0+9W7gPpmpZ3V7KOfiWI2ifjwb/GZjuH1gxMR9LSrCEc6AyShum0Vgqo3WqY
tHByft39VCxy/5gsTYgZ38ImqqtKNhCgvWxNiBof7B4Jt1IoaJLfbOm8QPWwXgq5
9VwX+Vm/6YnMFo3ZJpp3AYNyEnJMDMW10pPNgecxU02uXDS/gNjGm8pZ48JYQHNO
6xsfa32t8sja/p6d/VdtNgj3ex3NJjNJsiXw8R0tmXLdkyNiqp6qEj5I8LHtXErX
gxh4X0lNMcloPdeVxpY56y1ncLpgf8xeqhXsnO0rYFa9P63fjGewQtJunV/A+0iu
xIgfLJ+Axoe6GvVULIqoIoUmjk+FJUzUYikywaY9IMVF5uqVrBVNu0us2l+0llOh
vD1ktdv7XgGQ3/B8j1WBGkXQQEpmJXZiMhnOmmWHgXNSy/51j2dNA4wB+yyUcK9G
5SREfRthAJC/+bBdVR75fS9Nu3c9+lW/ZZ0fT1A2UaPgUmktTTnWzOBdf1r8vQKT
jjCoCXcVeaiMxHdYlAK0mXJDwxUIpybdbgM8CRqrrhLGfgUUQTrpDZY35IFwvNtA
znH0Qg3GN16Z1pEzjwqTw9HlFbH/5sqIo5+Al0ISogON8JYEjYaDlLUz7UexhKba
uqPtV3CiaMOdzq2IE+h94HecH9GrnRBLtZs5mRjEhccx+SZefZNLs7iomoyZW7jQ
gZk23K0C/G+Nt3/8V1lK0D+ZqRaaCWpw2gUF5eHunEd/vdxPxLA5yApAg9FRC3Tw
Q+yp8/vryQovJepiraOqbFhggFK9cyoFsRkhkwCaGSbavchiigHkdYbJRD7vRs+g
gFgXIXEwO3PpCXPFg9SKv1XSPveQFwfI4+pWq5TxBNirsMCxjVHoPRrCVwXziSxP
V/4L1UKKKil9faPZ7dVeoRKVJM4caUF8JnAXpF4S+/v3FQmHhZYCn56A2HLoRe8c
CqBzCTjG8Pu8+AoVw0yBGWus+p3j7BmWiJjDlhlE0ZN4u2OGiu5c97MmK1BhMcbo
oCPft0QMtol6+2sO/KXNOQ4BhZeux9MWbxG0MiNGSFN1tRJLsIgB8FJyyrheeE1T
5y+WHOL1zdnPIVCuiKTD3at3kSNhPSraNjlVRFbV9ll+EXjWv6ExYzT9Rquq+QTF
7AYQOYMRNvUZGxQAkUnpI5jhwfHrVGbPShFKCYv0Ha/4b+I6eNOE6TgDebND3phR
voWx1hoDfnNPd1WEJdlQ8b5u0HSTvWjDsn83fiCp6LpMoKgvJ5lY0mAnTRf/nd9+
biKwT1iAerKNUVAZO/rhneEXeShEOlpUTljPENgYPG8Nwq59tdGVan6NB4i52Xym
VPeaW8ba6Ao8y9LVkkEjRtOwq5V3s9ziP6Vx0TTPfaAaVbbYQqW0ahCRq3i1thiv
08egVWkRAELxJTdLyGiIG2s58ga9PqNRcVlNSBwtX5ciFL0FPqiKCacPJiN/lv//
Jz7iIDS5iV5q//Eumf3cJ8CZ4iRhITIaCUrh0dlGJ28jCjywMbI/yy3eY/8Qgsee
0V753lmTlJITbtJYrbrab7+l9umjv1AtSJRdN4m1FJvwLL9a9yyeBMfRWY4LJJ7Y
0hR8Hm2Ne2aFYo6ksQsvG0BKYKEHcTjpb6qdKqfYnWG66YYbhp8rz1UJJOfbB/nT
/XVe+RLT12kIoeGrUE42v+2/RVkxicGAyfHi1Tgx+wG7YclTCJHlR0Izhysg9bU4
gfdzA7VvuH/2zoqhOoA4R4Uep0/02LsVS6Q9kpKXmpD+bdDINI2pLOjcJqxvfGDW
Vt0MALzFesp2J62OTv0RDTB8Lr2RVZTsYMUzyOzZlC/+d+72BK9toaqnuTaXyADO
+WFVqOq9vnQqrkoQeLJOym7PsLFw19grt647rND7q3aSpb66o625vD08FF30qB60
0C7n5ClU+1swYFV4d51/kPB0YPGRWSFF7qBgDCu3sTnvnrgFRs1XHra6v9HXBjjP
MFFyle+xUTG7+tedJO4zHmzP/XgA5LaRtcIsCP1eUCiEw/jcz458R6dQq9AU2OC/
NGvq15qbO+JNTloYLzev8VMNDvlPug6TqkUJfKU4TTKM0nPUt7dY9x9HHm5c8TvN
HFd20QY8wIHEkmS9Dv3qolLSfhATdJSZpbFiOrVBrzVvA9XWZHB/muK1mkCRluwJ
xq9ZyelUNxlYNRnwVN9xhPJNPxRXC5l0bVBF3oVfhqhtw4IaAPUV3LSd2wAtLAwp
30NAIuhCwWitoR9jPWxTPbGnRYPs77jlSp7SdsK5i8qfzWHfXAgWQlvyErs+VN02
S28sFOiCwCeXmnL8ghC2gqg9M92FmDyMolTaPKgZNlRUn0mi4doMSGtAnHdYQ5tp
KfLUy+cOke8/L0RtnbgMCyfkX29RBCppAIdZptdzrvYtx8pXcYT6C3EV/nd0MCnX
Lkb0nE0qEDhpR4xqXH2vdoVaLLLjI8LoGVfY90jyC2kl0f4X/v4YHs+8kzVAVVvU
mZ8FNbBksOB3pWA9r7PTvysFmECs7DoBzhmyuBAZBsbHXsueLyt9ZIQKZBvOFWE6
YNNB0o/otghV422aY7RwSD38WX3at57FMZFwQ6f2OLiA7ZW9jGQq3+pwUDqlSfkD
qHvdwbfRJ7c6W9ntq97+h8/7+Jrg2jiXwhHYL5rlkHZqhjcCHPeg/dzYY5f7q5dj
9WTjZFtFzHihvp61coxtpryfsJFys2ot+EoNcTXzWu/oEZ+csA1SQ/YagrbFbsrM
EvFblRgHGtRJvxWwR6UUrgNKU/cOYudPIwnCJ6l+9fYaQBHMWIxY/zImwFM8NxKx
1At59LbvhkX1ol0QX6LbF3CK4Da5ms2wM7dsM6f1sHcqCKx14MQXkNE8fKy8Iq8A
Rs9e3Afn9P4+zu1vpID5GY53MIN2TXIKmaPxwyGgzmS+6wYvou+tX3csQMnCaYCn
W7ZlYAqvSZ2midR+gQM4ci1itCw/jlN3wogarkM2fQGHNSDkIr3E+gcEZ2iOjRAU
5tbM9loWBUfybsACItb989n1+L/cwhSz0DUwtKICgJ5kHxQbWeso2QSb6gsqcmmH
q1JLVs4Q9ZQdU3ROXuj5G/grwUScYekaKJntow9IisvxspA19tjTYr9r4DpMN1Xg
+3We4EEYzaeHK3qdVV/tPkCaYntzdb+JJQdowzVP7F9koleQfXzglmLkvm+sJcEu
sWT1fxCBAn9KDVdfGYK0eQeQEdYug3DIi6dM4PN5Ms2y9x8vkzWbIYt27YPY78PX
1ysPfWQIXhZd3OKsB6yD9LOqxng2B/Syx0PsRflMypi089OEpAAXekoYher38A95
GMiIK6gL/58BPAk5i0XAOeVhuH+17e0W3JKE3MpEiBMEqHeBY03rMQo4g0tIujGu
g9TjY26tqMgVuqq/BVzW43+/A5S6kn3rPtsj/fJzzdVC49Fl7IpAw/rrrg69Fahj
s4EmSIoMNFwnwFl13+JAR4GmfNsA184XwgVbTLZqvXvnDrpNBfNVBuZAJ1z5U7nI
t3UYjTzh79Qu1XWzL0Zf5UUMxtqjhruknuUhhZJ4dLlFNvC4K8UDOkYf18hPAO71
fkfLzzsO6kdsDyKJ5tr7yMDtkg15B/YxsQ/F2+ygcwCma+caZTB8tta91Sj+JoAj
au8st5lP3SOpkNLjchxjYU191Zv7DPpqdUFPxgPueTXjpLhsiMXyWFA3totk9t2l
KsMDpFavc9HzHTIVezwCgJ2bcRPDAsLBPcxqgDX6TxsPC2ovjqJckzk0siC35Y32
RcwXVgNECS6z8IW8wKTGg/vHmfsm+GdkQxUSRobdqWstyBlwjmvqeAyL+wSvxRtE
AvgdcWnMlusTVd9eEa32s5/dVIxfWXP+IWzq+bPxrEKLzu8GDYbD5yyolZaT/DCw
aPKGlF9Gr5rt6nZS6mEQB8HPp3W/IGpN/v2Q6J/u4y+wF7YemAKAx5RJFgSuWTFO
nhCzVePIAqCkLOY9PWee1X51ugVb/NTQxOlQij6Y/8q0jS/zc+KNDPoIHFH+V1Va
dcz3+uIufvsOrWgQPM2Y7xPg9frpH4KnOjNpcNozBaLuw3zX3bKW6STL3JCg/uo8
bmHiqWYnIZQ+qaB78Zy7lONwmChm86BBYKNpFZWq/LWvgqcSnKH7eRrSQDi1Z1CJ
2Rn6Y+w1PF/BYPlSYy51OeT8XxoQSkFnUJ6UnmWxaKKVi4vIIVzrG/Wy8OLbZuVX
FvfS5P8qgIplShu8rZzCQ1uw7euPXlZ9rrCDJocc03cR+DYqIwXNAe4BDS/+pEvk
owdgY1NuUQ+xqKxWpPh5iYhNTkF2sfhtl+PzzM2B9YBFwYM7Dlf7mYI46aL1fk7t
eNrZeWbLlVblyTIk4Xcb9k3BXEdLjtDUKxJxssrI8eb0n0ns3WIUIoYRVgyQUEu4
X10F3oClJ6ZUXuqYo8VRU1OmNZA8AuXraYsTBayFSf3CVhgY/Y+58rU0oMC/gC0H
0GxNbuBntNTOdKR4Nv9/MCsTzNVcWQ1QRmN37uBrVhxunNy1BBsmEBIN8Yfw2z/v
kLpx6WYQcmYXkwaduIGRJu/CYFqcAsEMHlQeYhFECLkuMYTfGy0IRNNu/lmimJCF
qliSmDjQWwdABQYnoA9IlNKPftRS7av4f3GsCPzvcExoQrA67QClRQyPxxA7MraQ
f7DDhab1J6Kfw05C/bZIdgjmVJcdSlL6s8bL+jyqUk/NVXYaW25CdU3/06Qs2Qin
BNypUq10zW1MOGAD064Re3KrHp9W6OXkAqnWu36PIL9si3pol+RkNiBiPOj8jDb0
j2ghjcmu/+Q8BRk1XbmfWKj+MZCqunNTaa27Wx2LG6w6VJl0/pqLYgjktfFwXcY9
CQefGSqtVPvqeRhM35cb6yF1Q871xky9etumoZoXswSg5IiWdAzb0N8uNy7PrTiB
zqZMDv/0bNT9QnpymP7IFiVXoKXZJKTd8HSAjx3WPHjnZFP6iRXOZCDZDTPFa+zu
Y1TmubAs8LZrQla9+XjVp4Z3RQO56Oh2S+F2LdwKzoDIRMXl/k5hbAHQ/C5A10iv
5t+7L7mUJquHN2grQDi1YHTkkgHAcmMU1x6jFaDUGyI3x94R+tE1k7TqItl/2FRc
S82DETTWbaoSg54VOTcFPEs5mkLUn19yoZljzenLWr7NAkpg7Gviotc8wyMrDTeX
i0XIDE9n218x8asnjY6+fsdADu88nQFrUGNGa3dyXG6ZRbKBtmY8JYbL2cGXVeCY
SPxLBeVqDm0+GZdCO3JRDVexvDgSTmJCF7YXtYcTcpT4mao/5cmwe1DWpeKSSfeI
07e4ppHqBnFDrSuWfPpY7THRBmQ3uxU9Wz0Rzpgt+fz05EmtMTDAUDmVvKJKJLwK
Ns8pkOu2aY/rhe4+3NbPWHl8SKSWQV4pCJOBMaAcYAzrVUqn9LaAX9+9cHmPjnob
cXKoyV0nHUIsxShmZJ0NLHyk87QbMAAcHaUGUkEQ/zdyl2UuTbe7MiknEj7domDI
cTxiBkAkJml70kgm/j8iLM2iZqPgTRQcDDV3w7q4+278k/j0umZpwxPfS2pethof
bta8UwB0iZ0Y83OnU8wZpXBCgW+JRHCLbrD23BOzxDsmsftnNbJdod6aVVqXi2nB
D4xtYIGBieerbNG+nU6Pz/XPWoyIXvCnULP4S1Tir05yfIT3W7S7H8lhiNT7EHSV
U/15mxRgbXFj8wwXxrIoLbNUFvsnxbjszNvJUBX7xuB8/h/a45u3fKUiJG31ln9m
tbFAGLmzRklzRZ1DSIcy9MnLILxWxbpAbJKFRcd9tC0tork9SIlcArh7NoxLbKF2
Y3/1wIzGfIYoUoVhtNpFCgN+YzSbVvT3e6S69Cd5yehlMLpTq5dzN15sem9NuwHH
KQWjGF/pOc0lliARZom8sTf3BI5iN3Q1IPlzy9Wx5Rr4AbOYgZFqBaw0Qg76kIWe
1ya2K9odk+B3fhkLtx7Pfdism3Cm0CfbgYcydXAbrX2N3rpwXXd/3DW8TVISwyGA
V2bZnsHzpSGBRAYLMAG0BEqGlOBkcZcDtgVQLSWjAlO3bP2h3G80m8ocJSFG/Bzs
s8/va5+4duODMMk+BRV1kSFzodH6IJl9/WfSJOmEh7TjGrMNRuax2QBG2KmWuaWa
3ExVf+tTj+J1qVjStAHc2Dms3jZaxsp6etMhk+aZs4Y2ruxvFooUAwWORkznAM8I
UsYsyrOG8+lbLvpCVres0snG5J1uIbAPHbBJxJa+61SLcniQStx53wzXW7vh+/mh
B4I/fCRxFGu54ztITE79b6CNPDLKpFMzIdKU6CHBOCvUYP/SO//lJEV/ENN6RqhC
rbZXwaq1DZ/duqB3DMX47n30geHRiZho/zTScaqzpHLbxzwHhrj9Nc7N4QfJmtYh
WjMaSTIxSo7UTihGPPW71YUI5DSDSLh/G0nzbdN3o7/0EH0UNDdkabIa7Nw1fKu7
Wl0fYWC9owEF0RpZAGEviqF8jaSpu03NUdztTrGT68Qb8HYweiXFgYbNvau1EMcV
i/2R0rLpgdPFyW5tUFx4NIlgMPTKEzKhJxRsE9hnB1vj1Ozvxl0ue+fLU5T9VFo7
49ckfk/WiGYqsXIQ1+NwqcOe7XiPRJzrPXcYzIH7gZbi0kQ0WU+YD7WsxGnWo2it
tyC7BES2QID+VwWWTQAPy3YbLjUTwuPMAPNuqlwiPkKExMcgBopcxuu5ue/PJeWI
k35Pe2KaJQFDOnHinQ9tepKs0Hi7A76LWk/+gE2V7epvydxsQHEA1K/GYDb6+b6K
`protect END_PROTECTED
