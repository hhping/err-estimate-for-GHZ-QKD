`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t3dQJ12T8Dx81ZJpUR50CcX3Z2d5uk5/yVG0ZEObfd2zbOCzvYH/viDB9VLbw5Pk
HGETj4by23Jq+iwji0sh3A643Ktxmw9KFDJbgolz4ct+4KF2nHvzBbA59iqy2TRs
bHmamVqC8AqO5vdgvXHVaP/RmJGIYgc0gdlSsr7WW50K4sPDC8lQE3kYeGPJJ4Kj
I6tuM7aYc2Z6UfsLAUbxNUdJg6QF1XjKaOvl4CjGrITbTOX93j1l0IcVS4zG0nbx
fj1KOrb2GidrH5FtWCeEco2eMOLG+8SgZJLtUgB/rCmfjItUHD7LGgK1nJGg0lx4
m47ulbm2ig2Nx9ia7Hy19LRa9XZir1sChGjYFeau+ydAtw3SJglCWm+p0cozOit7
vdoPXiOLLaK3SYBSJaSuWf0CL/YycMz/SktLESHVW/QAy9vx3ucvnaS9nAogF//3
EkMsweC29ooe9K6l7z4+0RUKm5ZvRMOuOe/1yiOdjomWZCxquuSlNw+K8tKo2EG9
XryyWeJnpTodQT+q9xgKakDCwKWkrvJ/fzIVfyeYGsOA49JNu9YJlGKAsuTN6iDu
JM17VRypHReFaX7kx9wCDNwRbQK0SE1WnZMq6ZGoiO5oRkf2TnxjKIDP0Ig1Uvam
zHy/ZnYj8ATcmIc3GZXSmiXIMxOG2reJEldcOjVRw2+iq4Rlgo6lZd5AAYFvM9oQ
bEhYZ5HEi5UHLrzONTIYVdAdiv4kYw0WiIQvpk4yz4WAI9OSzPlbM/p0jza4uOA+
yFLk94afZSoFoIUZ/JAmbT3wI4hcz1+Je85eUk8gcJ7yhvkMJ+6LBHQEuD/XoJEK
/8bAvv+oKokvI1y2CA6/8LbZw+56zBYcJOru7cvG/9euTfYzyc/+P9JpNBtsigVT
w66eOv1KY+OHmzKavb9wpPSemmWy6C9Gjj31Qvy69QajWZZUEwrLyLEZpo9nOGtt
if3NNeMo39koQVovQWQ5LJlhVFVQZnqW2rcRGjjP53j60YQlDa978PQCQfwB2IJq
sCc1n39gZPIomzP5nYejhbp6nzE0Rz5vkp52kLK6IdxSMFr33QpeJL5PoHB82Z6X
7OObj96s8Na72/5AINKWaIL1pc65CO9q2GCh6Zq15InUOiDrbBXsKxBgy3l+7xrE
agCIhlswgADErMaX1fL3CsLtqEu42r6dnFvwvnWR5AWpXJEvAo1ryOjWWqVK8iuL
1839U2s0G1Fo2lJ+huLQKGsK3VQ145vgYdelUeSX37HIcxtFCiQFZk6NzS3iIsoE
7zddFbhyTwziGYRpvkdyu+K75X9Dm1uscjVj3djBbwSZ2m8z05INN7UhMzlARtjC
MiFPgzDRnybEwHQcEagFTLJ8iC+jyyzzEkD/OQdJmkGg839cqWCW0A1J2kPI1kdd
OZeblu3NM1IayiCcR0Sv6IrPqa6nrUdEUx5TnoD+SgkR1u7D++QWakawx1Mk0iET
q0O7/WLlEeJ+hHFoKoRw4yCUY8iCO5hhP9BQptVANqwK1f0dHE06EpjuqL3wWwSD
Xu7Q1m/tQWKhIZdOZ7Qa7UHllRHFBFxht5jV7mHJhpHkdBgrDWnuEQZpqAPCJDxp
dugvbAXmwubUF6+cOHLTORm3eW42aveiafEQceDFMRNvtUOtD5gWJkz8fJKXbXPq
lkOLbkCQsZF/lxFuWF/FdSbuW+aOsWH7GTrCMbMV2q9+qwb7iljRQyVBzX4CcLVJ
Ol2mlI5k4aGDhNuB1i05g/Ukas1BuwT8KlqR5vb2jn2IQav3OPG2uEBIM4kKJsiS
g3XrqZ6AFnVM0zhXc1g3+vtG3NkJ+KC2DViEWMbAHbcWonVk2PMh4wPaBu/UIYs2
W+sNTMKVe1QcMXk+diOp+9NLoORx0Ep9Sk1oC8z5boWrdT98PgZtglIRY4IMbNFa
LcLF3WLKpMmubBq1vT5PZaqanfdicC/ZNPydws3g35iSSF5Cu/ZY8/JBzXQy96TB
4r8xDHBBjmtaWB2VApbzSbsA7sm5FPNz4FBllJPh4klv89hqxpqPXHNYivIqRUoi
M+Gz0xvW7Q7iAInHOIJwJcHsLryC1Mvwf5pGHF7JYf4hjZjHtKTWmYd4am9ZUD9E
69iVKnAoILcIuqCyKeXe0FjdDnj19GXMGTquwFhRgOiayg8uIK46+mqYij/QxC9r
V5nYhVUg8QZ2zKzMSRP24AlP2CP1FKbdL8fQiza0+nygsJooDIdRF5Rnz9CnrQun
Ngg6+TQf9aEIuDWGUJ2k0qrkoNr5yWHKcoxJHxx/UCXs9Y7phxgTmbv+Hl8UWv9h
Lr0uWfrT6a37tLhzi5MlkaNDgwcBALeF+rLXzEniuIl3RMA868NxX8YQ+xJN6Wx2
zkMoM2bm1BX2SAc7DDLg1tQtA9+OFfym/aRAYsBexk7RSKF2UbMxW2mEugSZIpS+
zIJD3YI9GbN6NXYxyEMxHF2GBZhA4N/qY+NeAWQwK52c2OKiSN7NYo3wQNQR9v5W
8cxdnBnVgb1KZ94kEDYMclxGXNnpFgtKI77Pns9quVvX+xvrVc5vb6RWE2zqhcwC
2TqwHWTF73Hn7VYvqSl/wLLPPa3HcVLryrdHJuEhy4jYONUEcnKKaOe4Zwf1wntH
fUng7+TAW9VyZINxh6VIHEG9hQ6RDQwUetUDNA3+O5auCIVuJQng4Qj5PZADINuS
EvLvHM6nQxjPz3BZM7P6VgYkLn7qnW2K+pdE//xPQsaT1ioEly/fCIqhOogxXwYX
O9jAJF4kk3x58v02sAJTH1up/BL1mvru1wuoATokUvvBPXJ8lbKSzjkfWd4lMYym
MORfqzWahtJ4UpviGb//TFy0aUPT2uJEOJ939RTNFBgC7jmLSgvunSJrd7IFHF4L
iA+98hphor8JYIKpQfgpzo2AExIGDwBr4GuIjxk78fDGGNjVAnZkfORoEUtDg2iX
uA+DgcMxrOaYGHrW34g6dFCVfbRWO3LJ7EFs5ozh505YNzBwgWL5xDS35+8yQuVK
fWMkyeEh4mzk55MI2609ZbdwDI+X99xOHIazx8fcbfKDV5r5Y2K9rMLDfVuTc82T
wUPfNyIJx1CLyZe0bm+XhA0TWmQIL0zwJvcTrm+J3UhvN+GjoF9dKeHOeXDxfWAf
0wCSIF6gwf/KiPAem9M/d0vA6sfrjpy7WsODpmZtyMW2fn+23kzAR4Ni3EpVFKCD
CrTjPR2Y4aa6iK2hJ9JzeObFSh5Z4pxuWptZct9lrRUtXertFOz43z4VZBtuko5G
45+Q4SnyHoNzdWdVF7wMwjTDGbhkoHIKUzasDDg/jAxG4fVl2/LY/Uwa33ulo1sh
O9Z12dprbeEIMPNRrf30Ue4duWbb89BoOivHKbbzJVgv2LG2FNPmdglDhVp1ZpYZ
nqd2xxP+Ex00wptID+rTCErrmA7nx77MFP7hA7faIpoG2w3rkIdn/S+MjdbOmx+v
XLY7E1a48rhe7AIEa9DUcUQ/npi4/TuTpEjo738YEylxX1rw/ZXigIIuVnGS8waj
apBVTAXBKonY5kO/u889D3fgx4aGVBnBrbM8omrfD/8xfX5FZ78x8P3DKwQKlabc
YODWrjb4WMr0Ydxbl3X67y8ozPin6DJKqAqJog1PMvkVnxllzBVyecsateoXC/nG
Dw0mtPfKxlPV7CYCZ4aUbaE54eBO/Jz2ALzWNdx0ki28LzkDK65BGPX9a84n8IZP
0Y0FilRocwkRkp4Uqf7iWcEnzIVOghS6bjxxFJI0Tpvr6AKXWleWXmHNtYyk7H28
yP0vAxt4DjwV3KdAUdhuHlF2oPwIRSUlto1G1Z3CIgzpdY9o/P53v86NvqD5IOTZ
`protect END_PROTECTED
