`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xR6pCSGGpvBemPEuye5NlObw75kcTJ1A4HIMk4+daV4MATL6todOF6Tt6s4PMulJ
Gsr9ghXQ3b8Omg6miUDKoMlw508nZtXUlJmLqTAQ0WdgDgl6h8ptczMj8SFyEJeE
+v0nJpyOR/kTwbgeaoSG4OtjeQQDBnwM5rVoFhtXI8aJarmwL4SNrjwbvjW2q92r
DIZb+6xo5Wq/jXBnIyhfXqokbavrWvx8DMNtIdfDM9QVi3d8v02VE9sptlmcf2wn
eLaiv3oucb7b9tFa659K83KHO+rz3ZBjE5cvArgymk+/Qn9bwtJ/enRRcxp9/rh/
E8hpsnKZ3P0MaveoVKFyUihEoEbXzaP4ALdKnDK/bq8Ht7yfVOu2xHxnyFdCwXGz
SpXcCv6DhUKum0iJusXzU6cltiqc8KMTadHbPu3vKYQLR0sKjGVJQe68su85xI9Z
hD3vUfzQv2zHTWyQ6aSeZeXObiZtGgmyuMndoBGKC86AW5i5OaT8WvKWb25x4IFz
E7yE/YaoiPZNl2H0so+Pa+JfoZaa+8d5AXj76Z8igFUBaqk2lEWii93NBzQiuR5/
gPtthwTfVck2cbMlxEzGTviRKcVWEU1G30WkK4ewqcfRBxDdAB6cyKZZXMATedw5
4SuOuNODruWgYyGW9drlm7N8/+IaiV/GGmYAP93Dsj0kHyX2tsVfRgqLOc3fpRrk
bK4iAzGov5P5Sj/ul4WepvbmDxHgy1G5+rzxIEPGuWKCXVUKV6qP1q0069f8wzNf
zgm7cgCUJtPU5MTBuM+JrQEvyzxWmpGPY7GUErmb+x2Ed4zaZ+rgAQ5PVj+4uytc
2vGqQVb6A8PUzWT4OJ7QV8ozBMYzLSIC/fip7RsypWzzIMu8Bb01oTFkEHLkIQCR
tubdI1nfYbcaXTk9caD2myzqS9AWEvS+nEHsbDZXSbWqKmQSPPRX4133iqaeU2sN
lPt9fQUgxak2z43oLxawq+HaWaiZW1x9at7Nd3LJ2CkeV5qWk77UspjKo4EFlxKf
/sbOnJIKHZq83Ozed+MKl3nsfPthwptDfFP7lt2PgrE6df0J77QZDf0miluqiDfh
c0fikt/f8AZPBd9Acoq88BXTsrgOp2UbuBJf1/rEKV4AS/5T52Xs0FYYfjk3AOz0
qSvBJH5eR6WEeKkQ/Tk3Pik223gNDwqI5eSrKI73wlwTVYiyNn0zAW7L8ti91xXp
s5+ynkDqkqQR0eyXFIWvEpxSkdBynX8AlkD+7C2IDD3bGz+eRRhFv4UiOEUtJXzz
SFyzmcEk31+oyToTJnJCDz0d5/B8oTxn/jv+t336YsNdVy/RKf+F+PEfrQcC91LQ
W7dk6URFvP4br9HU426YtWSbXEVsXXcr+CUR8HhHpogEUlCE5pkO7wwQy+xNF79+
clBGlvNa1VNIw/VNq/3cJnACcRUE8E2NGWTU8Do66wrz+Wk6jS6MyPJK+S6KV50T
ryIfTMRGqtFTy55Qo29be6CZ8WQSYQb2s9YNuPJ1r2/2X8/Thu6WDh6MsPWwa7Pg
ZULiDNf6Lvmy7cUbW+eTIPD8Shq9IhTENJqKRJ79pMfEDCj+r29WyAKX8ZLpBu2n
4DFXY//kQMrZFEhxCN9FExdWISwAxWvzf/N3menHA63f4M3PgTAMppv2wfYtYZCv
PzaQW4rZjFNZJyxqrMWCjOUgMbbSzo8KC1r/Pk8UEIf0RjqVbCHKnORbmhYhjW7b
gXHSdxxLp0ZUeSRKsVAnXWd2ILpXEVFqajf0YeUbvI7VVJg/zaaJn7hvu6t/R9AA
G4RETFZ0ocF7AE9T26TgQ16o3JB9rpOLPgwbpBRo9q2UAcyHTm8sxnbbdrv5J4ZJ
ssbFQ7ucDlkfkphUFSLU+5rdKaIl27xh10J2eVVFZk78cahsmViS5SszwRPbAyJ3
wQXxJ6fwJRM2wOhMXylqZCr+6Nzb1tcf2y8E4KkGHqsLFf2DnjbST/emQrKM2aY4
xewu3Ro5aGupet87jAqjznMLeT4NLoD5AJtsck8QCff6ijIsRoLB1oV0fl7povV/
tOp+key+NuHmqIIGzudOYhQ0orxNwmA1zzBQq2tSitP0I/k2h9+hWDZ3/vMzPFyJ
pTyP7/i3mGaJM5VQ5B1Bln2o5RjrmdiohJSZkqSWir2n0Rq1nRufL4clK+jhH8R8
GXx9Ycd8Rw5Z7TOvtixnSyfCPBPvIROwmibE5TaGPFmv58Phx6M4IPekOz1qz0MA
PWF3FDTvQxSCKecOCtCfngJ93PllOMYWHAWO1D/fiI5Znkioii72V86ONQQqUhNb
pOKKnVmfde0ze+3AqG9RQCgzAT/Si3msbCkoYJMO0iZ2N0VyXrqT99bbj4eh/x5g
WciaC0UX8LkXJs/egRehdg/yq8xccAG68tjk3g4w2QGkTu55S/y0UfhjV2UFw43r
qGEYP7eaIEScc8CsJzYzdG5Ojg94mocUWH+lxO83xFV+HA7QT3XlVUJm782DafNR
hmnrR414/K43r2GeoE5Rujj3KJ8gf3LpB+b9j6kFZm3p0As4NSGBJvvM+Zk7EFLr
bKS7vSLyOVrZrLvkSj4yNm8TvS5lQ+VXOTu4I7+6MzTjakW3XPa1MB3UYg8jG22y
oBJoSnheWruTVdLS+Gp8o+gOVzPTW1cMsbPpIHmOVqz+e3k5IkkoEF/5vq9gBaYb
y5aWViDy6Oq9k9BzhJkWN8Lgjr74G9zYEOsPkWb9i5YmvlLyU26HUp+iJrgVNYix
VmZiYVmayVCx++30O18AU6/erx8JnzblLX7BRezpK5h5k1hveaAFG6e2KWF33CZ6
4yrw0aWJP8/s5CIdN9puErLF+8pvzsOqRsKm2eiyN+lDhzKOKtKX7y6TkN4o5GN/
+5/DhD3ET2IkhpnxfFZUbEeH6YjVN6vcEUD5wWO+1CEFOA6teub8TBEPK9qaU1kv
H/qe5TmRHwlQ77rBY6LO6bkwkfySkJr4bd4kbVHsIZs9QGyrZnq6RZZCB6Yh2ote
z1JI3FUzCd/ciCh+P5y8ieXDRMRnryLX7gAPhapGjYqIGK1ykF+gSq2zpjGGjnM1
54bjZ5Q/ZDLjjVnB2Y3Rr462Wvo3+Gch5OY7INaPLSFL/L1Mw65hT7bSG74ILkB6
RAJj5RuJhSg4HQYqbPwdt7aDhHZuYVpWBMQmkgWFjvUfojyYrKbDtqFjkwM2xoaC
q6jsX4A8IdEC/lK6khMFVieny00cEGeBMQUmQAb01P1phN39orL6pnCZj0+YNF+e
PBqUN2Ha5lvv5hj2HDcC4/O017tPvK7NarRV8CuQPupaAdBVSAUUpS2itSzUvPRe
X/U/YXqzZ2vLSswGRp4GZMA9K1WqBzOGEr28z5cHKpe2kssy/1nRtmc4s8FyNQvy
pBKG6LCqkC2Z1k0iRtIx/CHceaFu0l+UmYKTwakjkmkKTTFAf886Bm6W32Ztr5TC
FG40GzP0Wq60U+qw2V0E9Y/qLgTntqSBYoLsNFuiwEjUIjco3Fr6Cf5Kd+jVLJOV
qY7yStJXDRx+lNs1d/r32JuvuVODcucFNUoiIEgzlrNejv8OB1vehuAPk4gOmtfH
GS5xbfJE6sAEJpecn5Xy+uicGQ2LxfxTsJWO3bvD0hkwOeXvFIRHWjYF9IPG20n5
jWny9OTT2T8QZ1yst5BLfnJkZscFq58z7ug9zdPlsN1DfjohD3FPXpt7cSBtKVq5
AkiYxm7Zcl6k7L6nPJuh7pc7tKq/bqhxpaVsBNujf92B8ThcfFjV3+9tLseSNLjQ
+LXB2M1QVCAPn6URs9MBAMWfH/UG+5RXLk6RZnqXYyhcHs37uNt3KrOTX4KtL1xV
j0KZ2LwDweq2l7slXQAb/0KYY4aJsPY0kvFdCURI1Rsy+A82Ig6T4OKyj7qA2aR6
sQOJe2Rlw8oqegDhb8ofiky3GgKhPx5f7MXITRUaGNlsjcXEEMR1loQkxsrCPcRk
gBYrlrbcbLCbiPfX04G07EtyDxGcZwNHPt/wpowRMku0EmzEuwXmoYVjlSTZNAdR
QjA18jVjE82X1ehhlOtwmCi79AJh2Wpdmve3BNjK8DWJnhg+VKtTVhrrQassP03v
z3vbc9CunJiC5PltRfNWQfsAifSe1zXUElUey0pSEg9K/SmsBvBf4zii/dMBomJ6
XDBMW4bwsXRQD3wHaW6ZOBAzMAzHbR+ZIuNJn7ZjS0IQ/xIAN6hFYhVvirepSTI9
St+lsLrEdTriZrj1jeGlsV2ztilJYTWgy2GEc/AtITMHMCxjQwLxVzik0oeyqYVG
bNnluZd1UESLEGT0byX8gTqWM45IIA+6+GEDbpXlf4GGV7HVRoRd1DfV9nytEfwc
EF7F8ltyfBy9oILlJgQv6LUdICHfrTdPp6TCKYiImvI81zB1cv0GXdzzUtT1VaoV
0LRWaBGLFoJMfL4G3veKlHq3wiTrTnlwVg2lOz7e36DZSgPrVDbiCT+PZ5M3ABjl
RmHrwO/hF1Req5/A08bkj3YAlxppFfGE9aUfbvQffD0m0pXbVHh+1GysMad/7KrX
2VNxYUR4v9wcN9FWfPT7uHQGaFiKJNg4Vj6zWOomTAHFf7CktsS4ChWRz9b0B8lj
nKcoaZJ+9TUZdk2YVdHZX3WUO+Qx5u6XJNv24y8dWh8WWZ2dM0A5dTYmbSt4BLur
r1l1VqVHaixKlP9oDpiY1dN5XILDhNJfVXzB9TX9HbDKfPoejm+kkvEhf5mbT8+t
C/Y8lYWNNu4qWsc4OddsrXBQIO57GnUpYAmhuXSxDpUaqwFQDsD7Jqbkh4LA6qIt
jLL0XMrhkYQZjvwi6NpRhrYonWFY4rI0xRXE2ig+tJnpXbL2e2i6TL7eIygC9jtr
OXca7LkYPugxFqfFMBgiCErXo3D7FrOyTAxahRj+G5VRZe1BpkMP+RJ48espaGzi
9c3z7+lpUNJMeeHGZeFhfTisq6QWFKvpqz8KMMtUKoVp3Hpb8DAjQb5aCbebu7+O
1L0bIDb2Wa/W78Ldiv+CmsWFzSpsupkrC/UOJ+ODUPsI8L3Jh34E1jZU+UkEe3Kq
jHPdp41J+2Bpg1jyIlUh93WI6ndDd/EcSRIMSUIo5Lx2M+2Op99u1cBu1trT+X8W
Q+5s6jEzJ5ubpdIhGYZ9JNR5vWT4Mf6I4757SJWCKEgETrJcU8I4vEeVQ7Yth7jC
1j4Ok0qFTu8Dboi5BYUbC5FalFwrkWrJ3VQdMVVDTlrGibR4sY768sbBx3yKtlHJ
w0GyK7ODucQYv5v4QlOFTsOrlCNM5y5eUeQFsDV3xsIKfmdRc45dCThv56o6ed/t
Fl8opYNzp/qha+VhGZbVlLuc4kxdzUd8My4R7KPXjKylcN3ju35IoE+s2IYkETAX
LjibUtcZSKsJ8X4RD9gHlBEYfWHclgBxvGRWvZZkk9j3bCJjc32J9y6Y6ShwLUov
TH4sJRZKWYULfmQFwHdOz0lH9+DTJtSfBQfltLijHhOJ/8kxYWPXz6fWFlskNuXF
JNw4tkDlf4AR3YvcqJJKLfQVQBd05M1b3cLppw/GNn4jT9XMDx/dFVqfQ9ePHFPy
cmhC5GK1aqplQl+CTUobPvKGe9S4XDRLVdstFjdX7pmrMI7H74CpvyvyCuc4oula
Cq+f+o/qhfJ00wu5FsS8EP3I1EgZe67snC/ssa3ctTEZP0Kh9Ws7YT8cC9+fImuf
DGnhOsrKdBwaU9jr82czzHknc+LgjoQQCa3T4O7QyG7YS/EBZDNCpezAVYunQX4g
woPYtSNj8GGsdsdxT10gInk2Qg20ux5O5U4WclwqQLcPjH6Lq0+0f6VmSEXNFEBV
zciZxOcSoCr3JMVjdXqEzU0mgKIsQ4oDwIxh9zgujQ4T8/O07+nqP/gl7w1IV1RD
0eCVDRCC4Hdra734IOORA/+evIkFGmophv2rbaGnFBB1fy/lJFVLNqGDAI9zDAv9
ET0ToYrlKXnRGs2YS8voDRP4Ea50bG3MDYhmfz6z0HXCUwCmP/nlvWCcuQuCqMGr
NnVKcYSSxQFkdjRAOwBIuowWzJS/qXQXRN51XOPP8oc44ao1kDDVo4ru5AP0DGKg
dBqA03riM7Ars0JUgcqeL5Xvw2cUJHTZsXrJW+R8y9NGyZYEatlQ9AwWjosPi9co
Tx7DKJYkjxD9FyhM2Os0y4wlOKXGlgCe5ZsvQTZ/gipd1P+EwXn1NYSpNafGyB/x
QoZ55I+tSCUHBv/mM82f3VWe09NwLPKQmSyNT+RtDjWQM1sLCq00y18sbwa2Bqky
ju4POrnomtAN5OzAHF/886Cez3R46SqxTtThmgHDH8K+N9C2UA3s8UIsvo+KQWvS
HtVZduzjb9UvVLCRxXTHDv2LbrVXaI1azbN1oXXthpx1UCTflDcsstq129g0FPR2
+HaRg3VZF3O5X4PD0NRaaPZOY3DTeymD7iWVqWLauRYKLslrsIbZJagx0+zSQNOG
tBcM8jyWOyFj4kF4IjDXcjUV72Wo+lXeRSqv/KclUrVF026NcrmTsax3wlk1Gfbq
LIYLP0ESvjVGHcgNEtSTVCYf6BTMKaNbLH3X9aK1caDNs1CHYxgdnSFvjn6riLXb
OS8CR75gC3uMZgd20iK+tdXgfd/kCvkrCkO8Xxi4nPzoEq3h1b+fZ9Ty13qGJ/bl
/mtTKX5Hdvv8rL9ZrUrgwAiL3mnN5KDLLcthayjgUExvrtqW06CnA2fC39ma3rCt
7t+yW5G7QQPpm7MQJT4BCPIFjpwNaVAx3aNb6KBrSFpqbbp2D1gapBvKr7Oe/07+
QcRCWLHjvRdeoEDuNzPg8TlR6brvMjYjlqc/7DVD4/OJYLFFM6NAP5ndYmw4c31Q
xMXBCmNtnedzENqpxIiqz0cPD47Y2dKCyvb/j8DnaPf6MQmmA/ZeCg7vqmR4TY7F
j8ue7Rw5BoNOepwacWV6FXJ+ge6Lg1nn1BLoafmJs5QvxunXBMuLTin6IaQI/u3Q
BIW7p5wpNd49/ejepQ/ye2CepngS+cENxxyKCVVO+xicw7T2Q++IW2i1i25fpmiN
TAgriRFmhqFFN0kkkETqzbadvFcGlaVXa4g5sL/562mS/Uv7K3o6hHCioDbDaLs4
8EVWVsYgiomFDu8Z/2pxsRdg2qOc5jvGbmSrkOlwtgACvxquRQw+hpQLoGI3gE4u
ptbuiJgIFtJm7jdjBLPEfdKiIhxX43Jrxd4JmTRmDutjpeYG+dcxhsroCT9/6ota
6/XmI9XANNeRPSpfYns1bUDAw1egg6hGrAFYx+UFbIBtv3FnRZEKV3NHE7Otst86
rR1tp9bQBh5fHtmXY2XQ/CHcIuYdsNpQOEByiBN4jj4JJljFgba2SQfE+vgIeXsS
b9nmGgre/v9NorrAmNr+3QtOPIMVhuvSP+CGri9qvI2kON6AgxfBtQ+ZQ3w25WMB
xCHvANgMRab0JXXT1GQb0oEDXQDcnwwqaww9DzCeik8S11HyAobjdyqpv6Hg87FT
x71Cqo0LeTHi9qR/LyLZGqFuE2ahi3EY7vKvp2E9ncxlRAtSA9/aIBQvPScV5/Up
f578uqqrYguvIDpuMguIW0GuH/OryhoN70znv+D6QcVb+xrywADZzHL3LKsm3u6l
B0tFh9PfH38rDdZTVnn02ZBwBQQhqNSphRiNuTz+lX9LmQXGpRUcwxArLiq2O3/q
YbnR3phbyehJH9rngn6tmy7I16P3GCrdSz5UTrLUegWFq3N0rnkcweeL7G2ZQAGb
YEAa85Hx4ls5ItDLSACIoPYs2ZRc4JZ8xbRrUNzY7j1+A0lx55Tcs7ad9lxGgaff
y0Jf5nNAfav/7pIFDmjQtZiXu9m0cPA/Y0cdxC6WfXRun32KvzyAmQivXyI1XDEP
gPGQaVxuoXWPpx/6xSMF+5H47yER2dL0KHZZ0FrFpDFmG6Z6NcuaBmg+PNFY4qEl
k7yYFLyax8+JF9BhdiOGTD3MJhl+La2frf0HYgEwMuCy94S6AR6y5spCESiNQcPS
8Sv125cakwKmxgR4X5ZHYgF6B0YwREsmXddGBpITcGPBpBjGqu1whsvXm9RI01MT
V2TbEMTdAUPOZnsLoQaSnnOpTqIyoy683nbPLYegpSLEEPYwaIYBd28DaYUDoTB0
hU7uxLS9ed07/YnfIZkLk0W3oCzURJA+tMKTxjfqGs/oglcG/UdCNup6FwpJK7EN
yNv6X6Rs4snvpQTZqWJjYm1Q+e+oYyT722cGjM2dZT8pw/TSy3LtvtSLPo81LdrK
1g+VNAXJXjFKam+XvYkFBmcT2+gQgtCpBHvrEPqCpolxxVtykCzBbGtvv7Y5tv0M
dX5DWVy12btJms6WqgjMGr/CrjJzOpjXir8W9+p/UGGG0nm3OA/9IaZYJUe5ID21
LsTaHhddRAYD5gagOFsO6+IoVfbe30VyO/Ea8QLF80hO0ZLiBJS91aVuapARgIws
zBCAHjLgSwj38r8W8u47JugJiJ+ChoJMycGKaFmvcq1r6foSYwJHpPrY2xetewvP
gsADvsnzOkKn+XlelnMuWKkIXQmR7a+mP3RZ10xhFZ6/7Eehrlrmx6du26KztR6U
7kC0Y3h3P1fOOpkUIYOuean1SxybuC9s+skulFv138G9TQukwSYJNola4cpgLDDJ
oEWRAhSJruAHCAP0VdoZnd8tdn7S9pLaufixM7KbOTqA6oQoJKzzHIijBREXIuKj
x2a9fYzb7G3rK0fleeeZwBckIRhdwK4eqNv7I1O4Id3NGale3vTtihPD1Tz1yjvg
ftCcXBJKAxmQOZHxILFWlc3qkQyUUH5cqerIK8s+KNiQaNZ7ymsGazJ0lGarHra5
0E4ercOdqIcKRZKtfd/StHj2h2aKh2Wt9b/viAJa5EOku/WNj1FSX9tZR/KrwAwD
2RkV3O8Fz+m1honCK0KkTyVIHJMB5o6a1efimzyyJ5gy1qzC9JiUlEJsyULHwKhv
5hs7ijLOJIa6SnRqs7yMTme+aXDRkk+Jpo2qV1s08bmFZBdq5KLQxjY0YcUM/1+q
0lJEUjs8Ulea2DCgkRshxnlP9mU8xMOyDBkwM/idA3DOP3qv8p0Y8XNs1ob/jz1F
l0+V7WRYPJ86UZdgnEV3mDClJO83lh9yz4/unFhRoaHppU2u9vdQs5e0TFR0v3dY
rMDOTV8tgXSkuLp37oR8rLSMdtmrSWidBrDTuHJ9YB/Y7RAHgj462/lOTrDwRLPD
2DOURPgyGcdqv5CqKolINjNjCBRWHvZjmVo6SN/U/r5/I0MKhmqpX1yXtqStoOfd
48J01wM4xmWrHDefGBvcD8KHF8sbvQSfxgiQFICE9vEWQaouGzmeW9maDXwnhJbw
RjCVOD4azsTOeMAQLJiFO3XseG48hYnlmqfD3cZrHUI6yenc63rHINc4RSO8WwtF
LItpPEG17vFr0ylyB7lH+Dl2lBB58BcQIJVr6gxj8wTBXCsYz4w2bkB+ucn7bQtV
RrN7rq8h8D4HUZ1lDzAN8OVcSkkluoKKFNX0JzdcF2cvJB4X4PO4CwWIXTZb4zo1
8UE6flYuzqAX/Ir25PI23sFo327mut/LYmuG544sdD+wP8qQbXTIYpciW66lhvaU
FyECfPGwXG6fwE93NE6HnhjpF8AEZ2yYF5p8AhqgY+TazWerJNTm5SBy2EkFp5I0
JTRKVrDALcv2fPX18giTCM/ZYiFqJ28Eei9MpnVulTLGi7ZEAwOFBJpDoIGOevgb
/MlwUyGSzFfYRRQ5jwHDGHgUUs0OR9Es+7ke9b9cjMLSWFaWZrLqu1FUcNsMfMlj
rSZns/X8s48zWNx9FVED0KBGa2GQ+SS628vbgmi91LiYQ9Jj/QhoVTx1JO4RxsOg
dVhLYoiwrrMH1hHqx4p+Kz1ZkV5GUI+jPDqvTZnGAsveF2Si7bFC8WwdkQkWCBLM
giReMbYDAZv6o9mM4cRnv5W0EYbVxar6zOFV2T3uuKT94JAYERx/XSuiJDFTvVB+
Oy1o9zeDzoxQofICZ6KrwJ5p9L+5e2hiRyAgcy03nF6qFQPN5QMCZdpvi6WcYIlM
r4AAPJRJZecRBqBHqXgqJDFSHOT/XMCK3xzf0DITCmMlttHzDKmKaKzUoSo0DStM
+gtLTEe5EsnEWxr3xYEW/fyPRncFITnlrZCO8P+YyM6/p7dl7voPIWwDv9XB7gIw
AvDvUuyjpToviQjFCDKk4/U9C+RjLjX4DMPTBhykB7Hb2x6xkp27URVqGgQIFttw
0qgIeu8PfqFam5I5WtBD5gEdIdfrkqcQs1JVthPhHNixPaelZkoEwmILcbC6bWX+
pNUJ9z2P0+sJTYFJUyX9aZeo8nGETBYT/OzIUqZDRqg3opdB2r+u6/X0gJHViK0A
lSZ8qlI0Os9LW+vbZDkFPdYiZJfsJBXXaNBEkD8b/u8Q9v3/OsV3HpuURu9rvvR2
3CyR97aYdqS60TN3MfnwX0Qusc33rn1iJLMWmPVhb/EM6xV3OZT3GWKmfAR5XoT3
UWYZ/UTSC/12O3tCF8X7y6J96DxO0V2dosB153WDBtfCPTwb26R1hxbkOKKcpXJn
dU2Zl+NjfOKFyml4M4wOYHhNSnqTCDEmp6EB+Is9EuFzq4uthv52tZBBPpevlxGZ
116nCIYaHL9Kr2zBGrqkXi7aUiWACgz/2MzvxusLdiKeAnfBzhCGr9KDCGuLHr5L
HBbq9IBtNby1rbg31qix97kfl996+5WpY7iVe5Mq1DmGh3bB/tJ4uPKxlcbnqYII
V5dr9BBrI5Ah8xorq0TnMCyroUEO40CyRGZAU/gIL9DVdnLvXEte9KrhnBJpwCVs
kd69O/ZBwIS4qFgpQb0ykFNetZVfFT7PpYpBb4EAUqh9RaBhrCWH23BJdJSodFcS
D8uH0QXv2CIGzSCCBC3d6ousQZ7eondakFxaPHTu/TM9TdIZicH2EFhjjhvWgNMX
K2zi3TCopEN3hji0IITIbi6H/pVJUyYGZY8IGoPNto8qSiMGO1n8VIgbR5j/tC8K
LS1PQkmfVyBPTMpxGTdBGW+qbX03p2TBxMaA8rs1DVRiIhCJgttfxCsMYZvJAcso
XrLAKf5/ucAA0tAPi3QOlHJJgvdoHU2siLB8j1fSidyl8HGb/KIEi+PWMK9wxw3a
GOK29Na6NCrkBPUSuGJE5qKG5N5AmX0prct4EWUhoJAeOx378NmztGXVNe51+t04
rGWC0tRGimyuzBwVS/DAdYcMSB3UDNlUwRDeajmaNlA36DBDAcMZXuRk1+Dq/QiA
d3tvFaFrh0s1Bz6qcrGAhY6e2R3U7PKj/IsNOi6hd25KW7O7xtLzI1J611fgamNm
Clqw3z1o5M09uCkXxlCM3n6K3J0yl/kbW58ZQRF+qEacb+OjpS1+WHWuKLcfniFI
N/YdrWlhNvqOepOzvQWYEDXjzYzl9JfaGQNnWGJjPZEVjuRsVOnpew4vArgE9ZJR
C3hiFhrbjP8QxXcIWeCMRjv1oDgs5MvZzp27Qnuq84qXrL1Q9Ee3kA4gTtM1oNZH
7hR/Z5suGLjzxtfCVS6Uu2LSUMk6F1JGclNaGkhui7XxKZotQ6Xuzh7Ckko9+uWC
rXRKD9Ft4Lgte6mOWDSHD0VfYDVnNv9lZk0I+82BHpNxfTK6016VrdDgbwj1DiiB
9ysXXIJp+u2nds9CqIACwWizN0EmSaPGrtXqSve3a5B9Qc7jMixa8Filvu3O7RVZ
XFN8X4eRRGBK3VvfoINqOm4T4Cx8t8Jr83JCOCWXPzC0gggwChO9TyxVQ8Wl298L
VFnlCuBfO9hpH2j/Oh+n9RDgMdexNIrjD66H8rUHJ5U/LeQmOew9kHi2Plll95h3
o4wmQeBgy1sZXbOjSKnpWwWI2/DHLuWRcteNrNQpY78Qn36vVFjh0Dq5Qj+O7IHP
VHL3HFujxwkhdZc6sS+nOo1KtdhcK33Y+6RFVJL+nK+lLEF/zRnNaZED6FzCScbd
BNcVvPNdEXVJt8heqSMfxwLZPtelLEpWPWhlS3uJY0p4DX7M7pwu0wJ0AvQzSf7j
jfeyuuUsqUoDiloJZPaBDrfBBh9IvO6LUVJ2+9kZ1VarX2BbDe2hYBqMA8/CEkMN
Mh4XHN1kiqw+i6anRypPO3PMrAP4o7kDIe0eaRZ7ZURJDVZ63u491sYdfQLdfsub
1NIEvgnhebBCnNcxXwvS2JJuoVGbnPNzie8oy4BJznDMGGsiG00oGkevewSQRlXk
rG4rYTNcywst/3Magrnem6YVxLeqLOOidRsyZef7QPefB6ZVirfA6l+FzMm5GLN9
9/37OfvOP/Pahvg/Qr6T0Z+1sTlrDXCEQpIbolDxbu1a3W3iVEg8btNoWSO7Bme0
NJ1l6GcJy8hXsdgRnMzSjrwJ1R0yHXzGemq+4qYBXjCMETSqsyIxV2YW68Autk+P
vyaKDHzTTTdtR4nzHoSq1cUg/X8iMu1MVlrzNyRF9w8XHj9MdGlnCgJJyQoKxwAI
38ahBV4/deDa0Z2fbxhdhUliU0P1bBuYFBwRLzZjmZQ/QfGjRRoq2E8HQ8Ed0uuc
uWsPuFDuzNtTr7c3N8cAfs4qY7RLUwBnB7mUTsIRo8cAj3AnBFSIQ4+zr4r1Y5PJ
2Wli43mcSVnEvUmsR4wr1yG0vYLCycxMPsQyg1+pnx7EvU4qNXHq0JRn0/LL0XhX
+xo4se8zAkjRufM+1ygl9XCTADJSFsWU2+tkl+AirLgzv8N3uDmFWAhdHfi3wH3i
GRBsK5P2tsl7SxTYxxx8D2U3lA2WiZBqhGhdqRLrPvyl+ikk43J2AyfXR5wg7n9B
wcAJQ5tluOUq48jGT/h9L5Smq/x3yv4CuZyJxCuOq7knB5jFwzwu9Yiru/cu/NOT
sza6OcsGdh5XCCCumBIma4XDVF42mwk2PtUwdOfdLlcL3Q40jZ1NLVJXzdlvfXij
j1IPYja4deg3/AEhYbHrAO0mf3MH0adz/yPvuPb6p68d2yJJ8toSjg6zqPZNtPwT
XvhLnz1NE9swIeU+aUofCGjTi985zxbBtUHWB7KLUy128tRc3MkKCbL4JFo35GEy
Rjv5igxoCER3gCThfGvD96gTekl6wfntR7x6Ic+VXuJVvM2ikzV/PsHVe+4pcFen
gh9JUTHOVvKkptfF7DwgbpL/HBVisnviLBn7Rp65r6SGVD50RnknUHoU81hVvqiE
8UlegXQTRgxAy7CBhoI9Rme53fR2owvQTKCtXpCIdiwgmcI8Hb3wlU2T3lEYFoOn
V4LO5+n6vmXTTsB+HcpJ8dMrpuwqp8rJO/Q2Qpn/C/6jmVwusZ18gsytn+dmKmjV
7dOvkK5QhmTMI4ExErGwF57ZHezHrNB+vo2bJeWds80hmfn6Z7YmVibnDBDk8qAm
SBDSs63rzz1IOwU3gOuxDrcLv9Ogl7Fq0D1F93+TLnER+HAfZnF8TsJzclXx/6Vw
ba8tnht6UOMwRmhdNRhRBfQXgLheLyxp2VwDpbbXkL3Qfg/OSQORQpXwdytBxdnG
Hhw2+vsOJLmbXmqCNS/z3MyvG3/hQ1gu3ecfnz3gAWraOGdBQ7y2gi259+TJUjZ0
RFWASnfBaHdL8WpHeTN3ZpwG5b4TYAyDNbfD8js/NCdMa3K4mqip6kIU/KXqYITZ
hiMXThvKL9ktznkIWhoxCoL5Ae7dK6hr2o8qOu6BbhbSxAgodM7sS8PGe4QIFteE
L2erPJ0N9CyJkMP4l+NyFdrUHlv6z2h59IGE5IcJgSgBHjVFWddMQ3Y3sNvin37+
CgTzxGEXWyk4yZKVwWIyIelP/NmsxjoBTkZroqODDbp69dAy+nLnJHL3GsXrz1wF
iZzHhMZCZhj8qLuSyi2f+LAD40Vs4+GtAj//9kmBC85I7RbBDLyNUgA1B2KzLXWV
0RUeEm1bpR/nfXET+zQc99o3A//utwpNSkmu21kI/0jBxK/q06Yzk2217C3K9N4R
8HnU+jRF41EmCxLQRDzKCG4j/8VmTh4HACTMEc8tTUZJrXwOVFWcYUmYYLHMQbVM
PnehvmrT0Fuj3GGGF3IcZYcHgAY+lA+ZHoGfby0BSKJDxuBs5PWrS4GB/6s13Ccf
g4OeZ0ViX7IjzfrD00YSE9SZsnLcuVzxRXBl8hvmo4tpqzskMQF2Tb9gS+j4OIfO
JFgl0b21VmkEm6y3dVvew/zpfdAh4BjmogYWo99ZGJZZVP+ZEKgKli1dplr6ldBP
y1T5ifE6pJIi1xNsshKKj6UYte+/fdru9B0PxnD4Lq3KmFTsHY4okhsNBDdtqzFL
avNfB612RgDa2J17iLs64I84l1JmPinZRoc7GWcBoJYwCVCgv4kA1eqAHxFwkjCD
xNChVr+tRDGbO/RufgCV+WDQKrwHaf6W9kmObo2FwRiY0FJGaOkKHF7WCqmBag8e
AW7a886wJdIrYlAgoeGpbPd5Y883g7GvlLmju4E9JTfDCdAwnW5yiBhsN2QWZmTm
jSYOFnZ0tbDM6ADakyAy8PLF6DlzfLLE6manQjTx9jyCgtyL0HzlIn6Utr2V9FmS
tRSew1A6ANtgamwyJPv1xokIRFMJvHOe6cWG2675g0cIyu8OPjsDHPhvGo24ZRJf
qXe/4M2TStow3/cF1npMCz0wH9ZO0UKelHxyNG9LBZx0Di+hxDmNCbbztLT3nZWH
n8YpO5qGyx3NYx2AOyCDPwGmaT5ENX8JBEPy+TER1Dl0WBPMc00wXxxa/9QAPHX2
c2qRszByUl/DF6TD5KC01hf56KXESocWAn9ESdaTEweFZ4YE5LxNJAgViMpsanIW
TqaisMDDzpQ6QU933ybnv/VSJCjnQwjMx3NlsEM/clOKvWVAi72ZxeVEHYwGctxa
xRdEaUFOEvw9lh/zz5/WbMb7DkqnaTAKOfVPilnmxwL9IDJIoLM8jNms3Bx3LIze
FnZ3svRj+54NBEPGxCZcxdIzy1PLbEAewvTVjNShL4cEtUhd0RlH7QHGDnh055oD
n2TcGVbokRxAtJwSukQhbi3nqVkP+xzfIw+k1fZKys5fkFf68mjJ3m/o/B72wt7y
glyxP0Rl77sX3SKNfLP7Ee1k8UMf+jHPnDGmqxonO++EqCRaf/rawtazlpcJvCry
dDYB2xYwV2YZ2sZ4IiA6qRESKhSKG2Zx6BvqCpb1txkD1QdamWaGBTDYTH1TQCTK
7kw+0onXYZwI3DggZHxh5iA/9ARsfSXDNFW7oX3LxsqZwNbMgi9eHa8Zu6NKDYFA
APiG/YGVNBTn6SGgqYwpVEb74MFBYVcArN9kJ1fEHoBF7T0oEUGg5niVq4DJ12b+
hwhHnjL4XeWPbyxJf5GWoDatST4aIq3jecLbbd3b34qiGXPPMAcfciEr5IH0XqAP
gCjDliwzCOOLXQ66VUsDUcTGR64JiUkL6s5bnkgus2qsHxELIoPJmqNFI0IUu2WC
w9jKxBy15DJVdC8LxYZL+OFhc99OrLsJ4fNCLUzLw4YzWphPzfMIL9Pr7socplTV
tXCCD1cyW5zQtXhNLV4dAVI0TSFleFlYnANDDCIm3v1W2tArPwljEcQe8tG5CELd
g9Py0rCE6K1slPg2E5ca34JW07Ra5gMcggRTsumEeen0+uskuFYHclIIhZUO3d30
F/Mf4CUiZQLOj6xnZPbURABSWivPcTq+kGyMZmDiDwq8i3N0+Yr2hXxlWPjzGGaz
15Wsbcu3K/Gp2WEzXmb3rdU3cXHQeaCZoy7x18NcTo7tnbyLTBna4uvIRyOR3jZ8
sv9k3m8q70840Go76rYqTzJyUNmSMW/ChSvknhKNJs529FxPWqK9bsGuGHq0FRO9
Ts7RNQE3q0AVEU+/ZMo2Mg/k3FFBq2ZoXJQeBKdn54cyT45qoFeN+8m9nzZGglw8
mP5V4PevaSf0R7iAWzTZCJVVjmUb4sQfHXBK1sB/SQTbLxtqi2iolnzUbWevIsLV
dvSMUCE0Iu9N0plGuUrcKYvY73bgIXJdjPs0Hz3YPTrPWVTdVoSLHAtKfv23Qo+I
Z2KTFBZNKghqQ5A4mnWXiw==
`protect END_PROTECTED
