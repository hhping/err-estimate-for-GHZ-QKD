`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3Iw4ONC4GYVwrOqjaFPya6J+nu+RPxzN6/aDoUWjHhfJdwuvjMVCc+ylITNwd+qL
ZeTA+3JClCHSiytS+WRnFgBZiNAUja18PFRlg3idte2MwlbIEP2R8MxKgfc4koFF
cvdnuSTOI7CRG/Ghy1Iwuovi/NP6PS+MbMf/7c/duSz4xaojwX5Zk38fKRBHFGBh
jJWgNhJ7WcN6hnGYMXUbo8DhWWa3rl6/lNKOrIrq85e43f05IQTNNMrB/9OwKgVO
FjgtlzcbudLZKvcri0exxlbBH/sUVYn+qMFP/Ae5o7Z6lYbc0DZPdhVDmzbDgW8Y
9OULzPdCAfgxUlElE9qq+r6BgtehCvS6tLxHZ0rMfzf2aEiXmnzU//NPrKbhH4ml
OUG9wfvW37YvNAYnSlSJ7vQO/lh/s4dMcl7NM6XkyApu6Kg2GtprXfQqI/6QxJzy
fIvQqHpM2FVmzi4zdfcaAhWdTxkq/Fhyme73ECPlzSxv6GpJYD8aKM+fSchFllAS
dEi5wRHTAeM8h8JiuSFSRNDVam7qPDXUZE/Qi9UqfNuaFFg12fcc4WxxMAOFcbIE
3kkr1nxFHYQ2iTx8P0vlUjHikoZbqbNbNL4d3RCuEALjXONrGilMNYBpAKdAUtqc
Xq1kRA1wGd74eDH0/EyV6h4sSrRlhliIzaltRQVPSLOI+lWS0XmdOJft+h0n/FLP
QRloz/Q7EVoSU+fhHxXoTdG/bkrimoJRYNLI3sI3tkj77rraCKrCnbsdUJZs/KIl
srfmfswEI3S++DVoHNb39cd+nbAvyYs/Eqf0e6mX8PPvkqrzAqFLH6EheWrpQ85u
`protect END_PROTECTED
