`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iezewROVHqnvSAYGOF6kHs1LCeBh9j8MYYADVVmZ2t7lZ2rRNB8W/7GVU3+GOp+9
FOL/QQzZ9Cv3Zd4JE42cKH+jQSvyIyQJxhlezmqa1E7uJkjYFgKjL7EgO/MpYq3t
/UJoH9g55YWqSygybozD7whIKcwNJU5YRYDZVwABYppMU307+uwWvIjtmbPb90Iz
T7khTWpUGsssyMHAOpvaTkAqCnoMnD2NGTwdQSD52tYz28rMQadCuYsbh6l7j6Sb
nWQaEPcfxZsiIWaQ1GWnfpqrYwxulyTqcqNX3OkkeY24LbgnnWFMu5rpx0qAh43X
9wbK3XSjlxnxJ1TaKom4lV4oyBWK+Hqptq7HB/SclVKARQLAJIUjECSRX6HG2aJx
a3TeI8j1WAicusIigeKnFh1alTLzqwLYSXXHNAUD5KtnoQ6H/XAIdmJEY7cSQtOz
jAgPWDga10Dr5hcFjPtLXIC7TBgBWFhf3a+dbGEgpLUR/YSJkua5buFjJuFqbjgh
j/pqaG2WDSKhk42SqWXYTEHMLneJWcADxp2xEcvnfz2aJPU4hT0Qiizn8QUr8Tbk
ODGxFkR0aDhVlCrX8489q3MoGjb37/OQ9Qz66oJXiNQ3upN7vw32qG9iP87Dqn2A
Vlnhu/LnaDLOBGjSCzSGUQrIfb1bMQvgBksx0agTygwhn7gupWcL+abtoJTZMhA1
clsSHBiQ8DJoY9IIRC79STQ4p4O5OvH8uMfeFpfFKNKaG1L19dCJtycQzjIqrqAc
vqCIr/Tee3sW+VH0WoqY3PaofGk25suTcMHvxyIZwotORy98Hn5UNL26bbh1rqp6
Vb6CXLE2SxUy71EnMDWMI394uzaxQqVolx1Wv3l+cSn2b/BSXSweeQ5BZRXqqsJ4
IeaVyqc7RPYGXvqRbWBwBQhrcceMoHgkhFX2pCpgJ9NTYwA3ziWbrpYSOLbEn19K
qJp8GeeZUD9xypRnZ5IXPR5vFFEQId6WtRUcxUryMJcvKOTjXwVwXIoc7sqBUYSK
lGuMG7xDV7nbJp3pH4o/nWsqMjFQkuyoYolSfPy4d+f5PeOvXyQjc15HWRRz65kp
9MTZKYPI7lJnmjbWRkm3o7fqn4lPWw2cqRwVNeEL0FbnlUrk8XGjrhIo0EeVv9F7
k0ZDsy53wuuUVTdPN+3kUHKBNyAUPUIk+dsHk9bgKAcGUYVnmDRfKALJVXVbS0e7
CF+YiVb04cSllWmhnbuVY/TIQ5CHi5uxPM61L07MC99g9vdB+31bGe1vRy1Tx+PS
yXnltUx6Lj/jm8n3IsgWcYBvIKWtTu3yN4n79FaStyBzAa1D0s+hn55RlBLthlYT
N5o7XjOGBuzLCFGUv3WV+7YwAy0ITEUEY0Gau46R7cETwkXAtWuHMENjpkWvUn/D
icQR8p31WDgQq2fL/eW7adQMOvb/VsrV7rouasNSrLPvtqL1EH397YF87GWJH40+
TnLPRz97AfwGBj0sEciA0w1XYooovPS6LnQAFA+zdp6RaLZ7bxg0BLNnZZsswnBR
YtuR7ZhWJsoffHFBAHyAob60bcc+9C4RMc7KO5SARLNkCW7mkXvAfsoHiOdMvn9y
0TkB6wCUKBGRNLEILDNb4/ONaJvB2c2eydGnKeCyXNXew/AnQVf3cobnvZOu0WFZ
nbQlflwzmk1tyDInE2y8zHc+DNKcMgEIbxMvgqKrouRrQg3hZbZi9nf2R2hUBtgH
TrtwnpLepn/WfjzBgSnGU2IhjoyHW/XSbDWVr958WNdRVD6gEcVRPEIGl2hEAFJa
0Xl+6O+8Ez9BpLe3Tkmkv+M6200yhxDYC8iCW5I2kUub16m+MkI/XT3zAx/3zHYS
kRQSujiFpjjvgzNaqQmZ0iMI2USsW2Ib1OyYsHiQDF3KsFAx+GgfWKNAs5acJOKF
FiqpirzdyeP/zo08qpRdLF4ZPqEB0b0Onx1nEu41RLx1lBxBsvnm/2QNgX11btTQ
oHo29rI4Ifn4YGAi/ex+kf1xLYNMLehYwXVqxlWzV9Jk/hA0n8ZSUfur04m/2u2B
taNuMH30ztgWZfzZEG9xEvDBO2uSeglM/uiF6/WA+DKdPytLaz8sJiBOUHxB3xqv
gVpSh5HWKI6X5UHeLtb4p2pkqdYNGONX1wouinmZOW1JzLosr3UVHKxF6NK2elOS
ii8sC73YzK2VZgnQ2VXNZPtyESKoGCB5J52lwXRj4VhnHwT9Wwk3PVjo3DsYd4IW
5Rcar6wBFajmtemWDsjTY49HFWivL2EY+9WzIncRC0QXd3dag5fn3ALFCuLapUVC
dda3A48c9WAbJ8B1JKqAOvxSWJ48NauXnXAq0lnHT9FsvJtbrX+NUmU1eq4XK2dX
tVhb+/pWXMwWVjE00uKTkhrgkISFf3h7KZYz71CyrCQR/MlF6G/m6GgrFLWbClHN
d2GQQUvgfG+VFY5VGkiOQ2Vl/ijMmjlgZX6jkyt101YHhZnjmCsPOfNvdtPIyeCi
jgcKHuOzXoZ5GNwtR9pMnMTDzYwHBT+tcqSpijOkqTeZCmV340Zi0iHxSAu4qtPe
LAQmphkAzZT9uCOVh3LS000j+43jN7lgedn3wSG/a/MtE0R8vggDWjEtL2I3+d6y
bIMSfgGdjyK5l5vxJBob13tTnZaqZueJoSuqQwmxAScAPljiyT1L7OTrFHDm+6aM
amt+Hd27FdqvMGqcUTDtsHWBDcDmKHf2oSVll+WnzzbMvSBA4q0qIdRBtF2GoCMY
7UBMtFVx8jpLrIdmU+9Kgj1DSB3JJpgwvkxYw6521KkOm2YQf7IEGigFdX7GR67f
nCHk+TKKvGWCKNfGyvrkGMEmJatNoO6F3X51tta4h6voJH+r3346LiwQGQujTKh0
qMnmBoIsW2l5KBEk/IKDHk9IVknRvqO+gZbpeArX+ELz2wD+wZkxu5rjXhZs+zVe
I8OtpcVcIAIAWaIlMRwpnpGuXYn8KwyxBUgphlspq6jiWquvgM8jex0Co+3n1I2a
6Pu6b6/bY1XqeI82YvLXpn5o8gbJ9nrsH9QQkURrQk/Ee4MA6LTS1cZevvDBuDIE
SRbMJIvIbp6O449jo+ixo2AYWYQY9j7XWxeF7uyaM06Q5tN5bKeSpxd/EfSg+A1D
wrfEmztsODr8OGds0ekzdSh3Np0wfk21A580e+b9i8QNtaRKYBqF9nYcLNQ06vvy
hXzwGwDXEsVPWiywfsfPzci7wzEaZtZ49bDZqP0ckPLyntTiqAytoQgLlJJ8w7na
zBfpZNWtrjsG2iVUA5qqPgXn4cyw+kc3ue0NuyFpGf+Q3aP/8Lyi4QeI6wZExSCw
cXeJGDxxQ6XyBK/9RAlHB9KtvDRsfKeDyD9kayelhBczIZ0o6h7YWj52wkQjrs9/
dSA8mulReCbjaqnzfJ4TqM/EGcEdVRH/b956iuleM6VrjiPa6fRJkIX/M7Gs/LJy
1g4bfya0Wm+DJ7ln5YsjJPC4s/NGG2C4Iejyr5u6oKusm1KdfcS/nVaUzxeu23P5
u319hndGWtLUlaVbATbDQ62XZ7WHVb7q8QagxfHdFnYO0ViaBSeMpAOCiPJaEwqz
bguLWBazLnQDLCVKR4ePG1eVzZ+R6nCUfNuZdEBJ5L7rQvY9qmKTOsImUgvgIZK9
gNP1ydRR8+pOr2der148CcU4DrfAAA/AeWOSfngbG8xPfwn1tuXLClJBhs7lR9iA
RUvFjvbmXAyI0FCgIQETVltKkY9S8YzJjmuOlRd+pUNdtHzn0QmGHDwIRGRU/Rvv
BQ9gtz0XodIV0QSpD7tFLC39+VJO3zsqWAc8+YnUzvg3c4maD12WWheqLkjAKSQJ
bKJiQc/MnI5TNoILDQEO84KZKqj+BQp73kY87/C5vazzZ53qXRURDobAFBuC1q2b
VxGkYGa8eIXKKLZdy744WfVHcTgT8M8Yxd9g78LVFx4BDDVgWKiCvBRDfFlbpa2j
VCANP/sRgatzW93J5mUJyeLGPc78qfPAOkQqaeW3hDj6bUpnzd0kLRcruapvc20M
AzgwhMMuMLzn+4ajJ5hl1YH9no3ZvredINTN+mGFg1rAlWSWD+MfcRTXgPmuqt94
Ll58gWytijSnaweKoUXQEmEMXl9p8VO0XQpt4pnhA3GtRGMnApMoPR7hlkWv1Y5H
F0j2iEjHYQC8I3+nW7aXV3GfrsGT8yHr9MTmjsxSdWRUYLStBqu08dF4mEjMfHxE
ksgRD5ZdjAwfoOm2EKQf4s1msUoLsoLciLucMXV3RHhdU+iPZQeQrGCQ7SnhugbS
HGEvBwM4+AIlsmlJX7J7gS8Qes11vqQdT96xYtqE6uD3SA2bFuPyIWG8iat8QY6s
LP0rvP3vlxBewv/LHQ3+2ijL8W0RUBtHVpzOElgkfsdvIvOUxisSn5M2njPLXaDw
TgSDN5beSu+cKeC4Fkk8Gt1Av6gdujik799YVAFqaticOZzWWarO3TlP0KwbJfIw
AmiEM6EUG7dromR38m/HMPa36RxlXaApt1GVXU+XGvkaUVP6Vg81sy5RlmW/aa67
COKKUFCj1DOrsld1csFq6NIwzOoMW88zf4/JH5bvplVaGJBhBL5o2BeOYLWcRuny
fBxHcM7MvawOp7TMkw0esgOB27VynIJucvH0W3F+WR2p3tMET6Q0+XkhFHd62yZh
XdYz+WWSKaLiRqU7oPAWi0hbNV/DohdGKbn/5A0J1btQRT11cGybaLqetHRO8nkB
Wo4Hl+7olPrBSJKo72csQHe31Yf0c+iggLRjalcQf+w7Z4ZsQ0KPQG5z2eGM6rGt
4NjkQ9ZWYEbNPBBeLzxp+w==
`protect END_PROTECTED
