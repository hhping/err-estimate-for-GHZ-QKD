`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OQ/G4oYzTdDi44oE+oP5oEo6P+BrJYWnHN7N/qbp5IEaU5VzNprWFtQwhTIDvWRk
DiSaXANFw+JvKOk1T5+bAZki3x08I6cxt7H/UFAtMFQtwayWJoLpEWF0mqSA9CPp
dJs4n/MbIMMZ3RvhDOwSG4YNUt3wYfDwdTcuNgtY5HQjeRCKHe6GMbj+sZp5p5ak
V6TRVuHBu8p/sybhggmDo8tU88uQu0XhvOXxqdqHWy3ScF4DtaRGI6oy8j/m+r/6
2CKSSJYXiMs/erZ9U3j6FeA7zet25a9xj84YZTXp4a4yncZPNc6Z1FAuDbAql3q6
xK+s7R/WFTjyyQ9KRgtJeAyLOdx9cWzTCGk1MaJjRaXbII2xD9rbdWpLUw4dx5iw
bwyRLW12Zc55cXHW/XiKsVEJezayz5THyrciJZk9r7mSehvsQ9hhkousdD4Ya4qF
qi+/mnbBMV4LjFibOGGZxsgjkmrjrP8VgsJHTEPhTEttRz61XiF92DR+9Rn46mbt
Nk0r7QrNKbg2JmZmjyw5fNdSB+h3JRwA9z/alTP9012laai6BozBdlVCFn0JT7vX
JTfjSne5tkiKu/m3K9Uxg37XOt/dneG4rrwYbIsAxVbpdaPFisR5dNrLNbZK7BEk
8R75/I6ozMq9rsiGGKwpb3nDmUGJy6L6ukqlCGC6BHEQfoZuUbZOEEYtlLHM3QzQ
i58vFxNRkvY6OBycbNKA2RLj5CV+sLNl3In/pXs4yfPE8spM8c/JMtuhIBg0M9g8
k+gbV5jhPMXUVfiDvBoeGk3weCwgifAB6ZE+3yHsSzcdnM1bGW6xoIK+hzYHvfC/
hdQ6mBTeZh62S4+sZJYV93OVgk3bjsXjYNreTpo8ckbMc14g4QtZgsul1g/jKtfm
8e52KDgql+qM3e5aHGBV+fbrNnTYs/RAzVU4mBvAJs76D/PI99saBQs3kOzFtEgZ
VEO0PoYLOLu+DVCAU1y4U0AJCxuIayWU3s4pt1946cVilD7OWs/GHnFcriMD8usY
QA046pwPr7wmRhiEdhGkrumPbjSep5G4cDyManhLmtMcVCRSkRjtDTULGm2mSHxH
p1gDTkRdey0zWYUqIegg3i2vQt4lMvSANS77gZC9ZQ6qw5RSZe7o5t9xCiC1kqpE
cyYhEh8nOkuDhAycspcPc/j+LKVOKM+8i+dYpcz55oQ12a5sKyMXuiDocb4jj9WD
Gx3GpZXQCHjWwh/+nCiKcxFumU5peyVIG2g5p2uifs4=
`protect END_PROTECTED
