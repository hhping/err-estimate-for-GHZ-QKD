`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mvi7npwx91Vwpp4ZasRajhB0S6b5nYQ8JEPnjEmId+7BbHVQxE8h9ycCyg3Lt0Ux
FYtcBuoDXNxVOmujYPn35MV8JgZEsFwJsNFHaUJ+FweGX6j1++baY406psHWsd41
GWekfo68+jm7RS1jmnH8502jSEcA7p/8MveNO4ZPwD2lZcVvCOIVv35MSl2L8e1o
DdYE1uhF89idw6NeJ+vXmwbctlM3c+tstOgM3MNnb656sqqxl11uj245bGcoSeP6
6rZOoiPrefl0txqDYu0LjWjQ7X3B8gSMt1pbGBr6NCGDCrjUmXoMxmBqmxA+AWMN
zasvQjMyibUAAfEHtWfEDLH4uisLE3I4yTrqiOnA505n2wFWEtR2nY3I/r9UOfTg
DPMd0j46ZdAzNY3nS2a0YHhAtTO9oAmBX23PTylVSBIcwBmOPBTPQ5sauC4WCyxH
M/OtKBZtAGUd1zCz84jC0JB5BfxXIYuVnGdBWGI28p787qmQ85BNeCCl/9cm4s4E
gUs5UxrijmY2K5aZZUF+tsRFm9d74M6RqUKf1LzKEXjB+WhsbEOEmmjk0+cbrZgO
hgEmYJT7CGq9ETSvfWseo24qVoRsRuH1XoAJXq6uf15URBcn0tT7oxqNKEO42DcN
qYPtnmm2pywOmkfEUH190ii8B68lvUSYkSd+AAxiT6FZB3q5xTwDBlvRd3wGQSJv
IALdH/FdCyBEV7MdNVly5H8LL6q+J95bVsxbYet8dLznXB1jgoOXGkXv1qfVpEWS
bLAfx4/7t8gQ+Yrr/DdE8UVSjJ6xVmB9cI5gxaHubdAX37ajZOPxw3S26sfMck7D
9sOnbwtQBXkS8w1d2aa5VHDOQpxMuDiDvLiMbXMVM39DbHp6ZGMhng603ERVdYbz
EIKces7hAGfn76A4TjzLLrb3APTN2N1jwOyaSA5/xNKjtwXxaiVDMXBTSkpQtQQ+
zc0Q/DZclFX44GOOiQy6pDKMIc7Heuh/R/o+JpVSDd/ii3qEwEzHNv6n6kPbFqu9
MvXtqvkuyxWc4VFrcIO2QtoBoFRRCiwrd4LwRqngvJ8+UwOPFCA0PzMGyaiCmsIh
WasM63K4ytXbEtVvEubyXGROYPaP45ORtO6mM7ZxFZCJiMN1DKJ1t8AthksyFP3j
YS3jq3AIii/ySxlqHZtbG2QYPdc/nR7NgzGDMMBWW1dcBFCvFZRLZKMU1v0856pZ
9RlUJ0u+/uJeyanMlWcuM3D/N24JSEmtIBO+0nKXKrLpsRxUUxSNaB+dA9jMp3pm
BTMAHbAiARiGhfhzXPqyFBvEWAEx67C+8MD96LeyvaYzukJbBpwCYmnZ/ZM0dAva
b/Sw7K1x/3ROY+/BbqoXeUjsZ4TNfj6fLe4thotsfeyqJuh0PrZQTDLZeUoORznr
SjwtnDH0cEf/6ULoYKlys7sJa5y/8jzwUiPO8NqjBcy3JG+/C+ggareZ+nCHq3DT
8i0/xMV1L/pMkM3lKLw81w==
`protect END_PROTECTED
