`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qIl3F6i/T/4yDz0E9uHahUduNW9SkxIVGW+9/aUd7DVZ4K5/pey7N+Oqs4Kpj45f
JTM0eifCi37r2VpBgw2XCK95h2ZLYqRWzPUNTXMHYrkKG2nU0kF/3x9yAn62Pv1Z
BRhikkMDCKDrH1O8eP4KuzHVpfMZqJUqsBSrZNczGSlPmlDRGV/XJSHvwpVRzFSN
ToKL0ukn1A4eq7+feoBl1Rlawphs0WkpULGmprIfiL9T7feUZR/Dqh+DcKu5H2UU
u6tg1WLxZnOMD+OymmZIRqfjXnGuqdKa5ZfQSsSoZHb3E6CVHMr9Xb0LksYFMrSA
YFBFXclbG9r7SGGpW+REtP0bH4+hGAcEGSPu+8hQz4uEA907OEJDkTq1kLaFT2+L
y4bfMQ30DurR139PgBWDJjt2SAvRxtrnoJb896WAeC8bzT4RpsPbB33zsrUAFKLz
9I1OFIaJqHu/ejZa1iWyCT5vkcRa3cYOK3RI4obqy/0xeMf55B86lKaRji8JfPQ+
GmGQc0Zi1Re1C/SPL8yQk3WeTFgHLvuuWSC8tsAXwJ83rJZsUDmGQ1ed4nUD3HMQ
ikuIGb/XYi1JA0uGQeLFsZ8316z3oFoaBdqxJdJAiRLn2neaZlnCPrD8E6ziSJA/
C9azTWoZMQ4YEvSwq+/YHOV6JnhvWd5+2m5UnCnCu31DrdAaBmUARkdn7VWL7lXm
upGJiAKzaNqSbtj/f5smC2M05eg6wOZ9BoZCPZYoV64nnKjmzQgVhX5sl0IBlZJ6
Nva+AB5+syDX+RpIhYnikcv6Ecqmj7i+Gi5h90V/B21bBpWFE89Pl/0VMCv48Xw0
cBTb/tDsaMvSKoLd9ufByABigGSsO+q395yHRLzK7I5uoCQVmtBLjjeTjskU5hCi
i61OBqD0hMk9thHXjuFF5eCQx+NRr0tUuB5rroe6Yilmxx3K/m9djuBmKsiWXohi
I5KjbuiGjlZ0QH8/zpYC7T2IBw+N8eHbtfZkRM/wXuT+vi4efPdQ6oqsCfR0tlal
xGUCoCp6cfOVpIZhvNNTHlBBXbOvVY+QLTaO4xmMRdrjVOGb6+0ZpfcOsaMguucK
6VADQEuuGdIjJ/3lcJqiArNll0zp4C1C+Pub115mP//bwhzt4X4C9xa0mHChzznY
tzmKA172EaWT1rZkS0gr3m9hRIPLmO7eNLRpSeC/i+YUHIDDxf8sbSEQ0ygoKChI
qdY8atgI+3VvZy1gir9VhqwvMj9eKpjtN498AzWx6IMGP678WBmQVMlP2Bb3jyPa
NpRD3cHg6Pm7MLI9+fbkM4qPSV5sX+9+Gu5/hq+EWRHMdAEstEsN5k9W/ES1Fc+2
UGBFKW584e/f9x5FIAWWLYx9eAwdDb9beQ2kcjsRct1n7D+roITam51bUJdoi/Xn
uzU/tlXKZGbxErNW2WPpUBiBulg3NKDdlBIPVAVS5eLYQTT6cePhw39G0ZxN5grt
dOQEYMe1M4lW6wqax7IwU8LgkrL5AyZC6qe4qEpLqN7fKpbHGpTQMCGeAJe+9GGh
nF+a+fYD5aiEkG8wgMVLbqcGTZfU6IcfZPL0e0qtLs/26FVum/HIZy11AGyxISmD
UNGMqVJ2ly/dkFjGcwoGOphGc4TkNFtnVIFHwpAoPvO7rigm+Snt9QQmN9uu8iFH
LN0d8x3t6JUKIGjBmvbjexzUO0BUUopdbfh/+Z9xLD2bsowdbrk5BzaHvYIgB2yb
GDHZ3udk9XkzP//+VgxYL7+17srwsY63uc4KbXyAJo5LlBfErYklABLE9cvR9rig
gV69e89neuIQcAC7TNL8E0eNxbbflPdELQOMX4U1YY1SRwMbZZwYNU5fkMYSbiTg
J61bY9lZ0aQo4ZlCCBGmew8SYUs3io2yCkSo/KFdmWY1kEE8MzNW0x6VA+1RZHZR
8BiiN10YNPDrIIwRMDOS9sZzR+ifVqdB/ydajy4xT2TBlG3AQQIPLPGRklNN/3A1
YQ73Z6QVh4AXPSwHDN1IXdfLTuTwPiEy4L2KvbjVKs1sc37BapvlFPnfKvOF2T03
01qmhdo1sEi8YyqELqiDd02fiYyk9eM2wtbE3Lbf/Akq+PbEclJNdSXOq61vXr3X
TD2LiohTtDQ6D0rd0UNuEKVqB7qZ6TJjU3yGBWp/f+etaRSakmE4x0dfCwod3mMc
DjCaD6pqW+aYOsx0XKVD540WMnOTGM0vBXpdGy1QV/p4EmuKJk/XXNMkH5O9H1+/
uVGtQbpuJaP2uEdzeqhhIISiWmiV4FMxEJC4EtGNS3Lbnhk+h58QkdXNYVtVVNGc
DIs0zEtxR4pX1hru0x7YsqnjOsX1bOnT1VXT9AtlqDsB3M5x7YcLsNlwj2wDu+Wd
vaWfD1s8MHuCU6Ev/akgVYAfHvKwgDHH1JceVHmOaJNbPv8L3YJY43tFvNAsPJM0
jEbT/u78iHGSHHu2pHmZ7/qTUd1EKU8UD2YgMEAdKHxUnrfpiWWVn3eFB7038/ye
e+ys0ROa9nJXawpORYL4LWwEX5tXso3srZm/HgXlCnZBTdGqvfzcRljOoRJNy5W2
KuBXz+B11xZrt2aotU7sRyidRlFfU72S7m1TRQUFrxoNsBZPR1cD1Jn9XbApdka/
h3Mnz7rz4+RN+qSFxKxBEv0WxOhChR8qjEcunkyIxbQp/eAdzMrUi/oItKf2uJbO
DQjlFN5wXg5ekVLhP8p7R31gYmjDPwkrKuxn3I8Wg7dJWqrv4RE8xG4MkxqtnSnl
avsNj+4KhQrSwLFXDL9clYfG3HQPnkWBTXVYRElZhYRJk/Mg2y44V6CLKJ8QXe/F
yJ81TDiwN6mxfytw1B6mCpvHftd2jdJ73aDEXCF3vHtWRaQbvxCNFSilsxPkzjKN
4mAgZPO52mlgiEmuqAFYhW5xTFyC4tWOVKkW1Ccu0xcxHsbHcnEXpWi2bFoBjF/y
xOdEwKk5PYwYSA2w3EQFoM21c/oxK7EVhkpJouEoyrbMK+V1m62pxirIzuotE728
cL7ZLR6FETf42xlxBqhsluX1yDWvYQinbII/QoaXbSgexMN/BU+7XT27HG+68T97
s0rSBqt5E2c3CgzX/EzvfraBOxJdCzkcE0NdvvUEMiV7okscdg6TSV02dxjx2EoR
QTCibVhLr9zGLgmXkHSNiX2I1GbQ0brhxN+lZKAhWQg9j6PMOTX+rLxyZP3pULbd
IqX3Sd8AFxhzWmuqi+Bz85fY6F0yTUWT0MTwGRBNB8E1dV1Mb1wC8f07MShvn7VC
pZwrL3bLZ+xYa9hEn4nR9UXsjYZkcIGpG3z8iHm4PCjMxhF1Mdz2Vf+pO5Cu9TT8
STmNYfhNAwElIAYiW2FrGdeCS8fXc3pHm9OEC2xYAON3BfdZoFbF+jb23UepIVCV
Hjo+KHlvfGHBTHygrbhZDERRab64TuJXr+N0obxcbJcNYWJiElD5a6MRk09dTLxg
j1TCOyCOVqqDWH4OfDJoPslz0uUxslXCNMwY5ZxDyeekPXAdP1tuMCRZPk5I/Oj5
UG2YDbsdYPw8ucSckpcZ1bJTxK+P2ghh4EqJk9T73dYb/vqCbAWFkQIyW3ggrYu2
M3fbeKo9XalH4trVHAL/2l5qaMQUZeFrh+/ewspaFGEXIUzdNrq6NNtDLMhqiiXA
pVDFZkG0XUPdR0puCtUpLv/7EgU0ZhkWecCXBANuJrnDf1QHno8KRaoxTyPIcBR7
P1bn5YbGOeVhQjjQHQjohx1sLgKfkGeSnyxAlb2xv6HzaVoooWXgjx1+7uqTFXGr
Z5idPRBJAuRqzsNxzzxMJDXS1WG+3ki93DmjpkpvYnqukubBQohQKMUi1k8OkAXq
PoF9IgBKlpAoSURvH5XdYYNKqT2mHM+LL/Q5j8w+NCxe+U+YCXZ7wP0y0l0LhWgn
zma7mXz6pmmJgTXb+xv/86o7n7xw4AdF0+XQ+7zc/+akzln7g82p/5szx6U7ky85
6LfRbrCWKmheyfIdbgw56jwQqAe2TBsB+6ORKGjf49osaiIMysDJSEF6TW9BlF89
PKeFOKABd2/lOyHhvum+xaoeh51kQ5FKqy8nFFRb3FEo5zoqEtGMpDtzyU9/cbu8
hoZJq9JjGAUHEBA4Mtn4DAJe4Z9xGun9WbYm3kkdian281Dvzayn/68a+nS1LBl5
ZSrYDKiODJjPQajNbcViUQPRFcuTVVMn7/Y0lY/iagS6EPNMC59WqJSA9JA2Iq+Z
IHm+15AqLJXtCqzSabE+93Uq3BBVwRxZHMSys8APxMAfPth6zojZe1lkHdOoMIQ3
NdWNsT4TQC8zBo5hDwB0Z+wS39W6s8VxFhp1Nxffqkz6BZuMaVCTBcLZ0q83EnE2
XYww0vBbyu+Bcnp4EpTd+hQ5uLjjojCEsI6oz0A45d295lj7dz9UoYagr1zOgjvr
Bgli0HXi4W9Ucm1AmAffBRB9AOQWjahG/Kf70gFbBc1zI0OGgrzRuI3ed0v2QhSX
dhsu40eb7zns7JzQj4A5RKy866fH/cn/yKyj2T+ugYzWlUl6Rciu87mv7PnVMnBu
HRYXGR+wGGpkNob++Or7F6ie70spnmyw8OVgyk3+/yxiWZqCMJR8DJnsU+krywnR
0mCouWE3Rldm0wXQuaL2Y53OQkpMVuapNELOsTlHouarDMsRhobvb5OciFEOe1gD
414uWcBmPGonOrYGVhq2kHNrxAEgxT+SDlIOT0yKWZFEKO6lrph02Y5411cnuLxI
uB7wSuwdYb+AMDap+feUAvxLwxjPBuYBiUjI9lpyvz7MQTsIyiGPD7Z88e8wbnUj
MfwtHl1YE6TUH7J1mbkfpfYqVAvNnFuE/eBls2oq6vSz+pOkDy7faMoSeSVxHvpV
dcnjJAgV2j73Pl176ni/S7iHvnNbI+1PPWmxn5BfWIminflSJA+YCkWlAX98wIc9
mzKzV7X7BYUUiE/gVZJA52Nl/+1JaTbfoZNBvQonL43KnWj16vVM9s8rFWrLNTau
fPbK+Li3IWwZGmA6nTQcZMmq3YOId84n8oLqFac7O0PYAcW0HYPMz8i35VhpjG8r
/vGWTqVmUUk7JXeeEZKvU4ISRFBV+heJ13ayHYbSgesLebv4ZpIPg8xucxckXN3Z
R8zbfkuIM+zRJm/Q6Qr9BBEoqzQc+OFU45hjlRIB9tygYyzC4+SmBeZmWKQCK/tk
WUUGPgZBG//NPgDu2HPMr8pRBBKvqhfqD702guU94FKvLdS+w0Ns8viaoSx6kESx
2wiH1sQxBVXo2BMLBpRzM5tmat8m9/rV3QKs0vH7zKRhOP1hovd0XWIXgn7hkk61
i4vcFuRSunX21axxOAe+uJbzkZLm8y6XsjbeyopGSH78HtK7S4a72UQ5I7EbZv89
SIh03Amdw+jQa2VVbPfSKi95vjNd+nigsMUxLGB5wvhegpBc0Z1QdPgRnXv7s2IQ
n3CxYz8iEHWhKuhmeHTTa50YnhwBLZGwVXh3NCP+pqb6t75lrQR0KN0xQXWWLLN8
kdF+DEWiXk+pGy3IFFawHlFDydoER5sWNH0EJt6FjWgzmssYZAh1tWyyh8SlGlrY
bQTAcx/t1rLjCsFwHJouBxo7rSyqL3gEpUr7Ut4Y1mGriq7NWYqt1OczJc8w/CN6
8D9rqLnKx5BhznFO7zPnRBwIGodffyZp2wkfTSxfovy3ad3L2S0INiTv9NryNnzJ
hEHm+CipHcDJkvj0tPtMX+z2Qa5+rj6R0oUVo2QTBbjZI/7g/PjZhDTkGYiSpZx5
4KwD2tFGZBFwvSGaqTQy48CimYWpCWjswMcuFXz2RpPd45tS7mNhTKtZ7IUFTD5Z
8CgzeUAmiaattPuT6qcX2xTpKPsrTV0LPryAemlUFavHdKAu3tXKQvrYEX7DG62t
Nk0OH5/6FGCxi2NQKRld2IzRQgOSVv1Hpdfw+Ut0jfRJIutPTYh2hvgnaGIhdy8v
bc11WBRPDzRpNeA/raj05kNUiErNbuV0UZwNd34A0WRznn1QbVWrpoalGhuaPbfv
0kCvWIAvVcsnSe7PIfBSMbJdoigeSJeruZR5NADOCP1rZNJ7N2xmGLq9+2c3o71O
XLfpdzKWMflfWtElF0Qi6dNUwH8Z3JAItMAET1xNGTMZ15au9fwNqG64mfTyD/44
60qhUjyv6f9yCH1AeOAmXUaJRlHSRONyEqMKyWKiLAhOIchqtKASUwwO3x7R9H87
Gj1GhmlZtd2SKaWRC8kG1ywX//5WbSDA9IvPwIY+2FC4Ybf65umcEx6kSvqF5dTJ
kdB53I4q5TS+W5gcNp3/q3DN9Dc9VsBdqAPg7Cm7Zp061TILXuUL5q4dAP77Q2Bt
7y7YEUrJSdJ0p9iXTR4lM2oWCeSX6Vm9R7wQl+BYISVuMqApHQUKtbifEeDJhpAu
yGKD/e2dv9aVfOawSvRSaFFO5XEV57F+hf0k2NbSee0t8mtiaGqrFhI/hY5q3cwH
vV9QrsGEAdE/3UaKSlPrp6Vt292PoL44quQCHldN0GZfNwIaFCXD0fQrla4jScOe
rv7JpnL5BdYPaWCplUhGhGSpBohGnIlpRd4couFVo/1w0Fjj6lSDGf4SJ0wRAfzZ
nqq8w54ak2lJkNLve+eat14I86PNqRsMTsKsMHzvqlN9MEstf5iOQUNT9Wn7IE4W
OW2VtSe46azrRnsG5msmvG/sEZHjHgIqjXmCFNTJxa9Xtyqaz3J5LxU94E+i+8rq
XlaKnXsheOSPTKS7cKaH653sMRwDJ7RlJFBF08vfglNjFcg99PiIzFbLMWgwf8o8
YRD+/uOX8hTKFSEi+/Tb3mEHO++XmHWfugxdN52zrARwoJ5Cqt/P0cBUWikcmESs
zenOO5X2+BQE9oRpCNqJ6aT01d6h0Jzu2p08ij8Fhs5jDAKZPS3goQF+gm68f3Hv
lW9z6d6HJwW9rBDULX8NPp31S6SQ2vjm86MMH755+P+KpY7W42Nl/Fmf6NCMqDim
1/KKUnT9RJHC5xsp6w4iTcbNLwI+AOgjv58yphlz2yec8PL8cUe9Y9VckCEncwqP
ujJZSXWSrhsLgvjUJUQrlQjbICpRo9hPbqrTaHAy9iRCu0m+NaCYTV3efczOnd51
EVUFM8gMvCtSYCIUt1nxmzPjIrTv+nk+2COFN87Ijof8lKaufAnRJoiddIjJnUfa
3XdWdRubYf0q2sf5XYjXvjGKQCTAawcB/bqju5YFk/cWXNuWZsZa4Sj6dvuQ19gC
5kaG7Q3gohzS9skrMI8jIuHUsqtr4al7v6cyytWwZAETl0ZXSv1luxyt/SqJt4LN
EYiOzn2BYajRLNWEPrZxHk9CNoFp6m+TZ9tbFZ00nOKvKuAKRw7sZGTjYTYzkuVl
OohvpvgPihOcRfi11K3nS9UZYBJFvgbHXKvSmNcP+B+tlDaA/Jhw4NGKo6MOCh4L
5fJY2MRz5HxL8MVkDsJ7bpKdp68IeIYBvRxuaxwcu8tEy22jsH4qOsCncFRhCd6m
2eDBdsUPupg4mik3Nwut9Ey79ZqKGZgfW6RCyNomMpRhb2AZ34L4kiPUeS/NEGtW
jRIyGHXRZ5V5CH7HrdE2+lzfbanatZmhL7ueILbfKoglLOnm0MNdg/+cwjvw2KJp
D3l6U/Rlf6DdX3MPbYOgtdatsbnK/kj76ba/29MqPAwUvDt2nBlmcmeAbwSeyZBd
1bBeU1WLQmCaL+cW2lFRsqEsqBPp9xAfxmGpMYSB5N5Talm8Mj/KiLZKWws2ltw7
acskh4HFgrSRryC+IhUMRpbXASE6ZJPrZBn27rIAWwXfVLe0HWZ7tGcoaNHjQSpG
WFSW7JHP231JFs4wYUYL9wH+NswRGam/YZpyrc78uxzfCWrBLz35R7hdliTOk8fy
sk6dqKOrdCYZN56h04nQPaMQFzpeOauZr5dig3mvwBg953SkbMepZvMqdv6hMeZD
1imHQBo9mPJoFTA6nnyQsWUDcpfB0LJd7OKp26Ab2ViWZw/7sIS+PsbJKW2sY6q0
DQLeLLKEvqO3w4rduSru7TXsbZukH1WWiVYkD6hyP6ozcVV988pUxUemNIx1HlUi
Zrd6ovq/meUomLIS/pjX4IB5u4wArOm4pBs9lyZmzc294NshekR6qEVBMuS3gZhc
X5C7r+tnVCUHSw5Aouo0Aznd2E1lf3q46c3PVufBMWF+EpHlzw8G8UKNayzN/jCY
Zrp8adR1KcxvYR9WXAQCtkTL902gqucxJcl1Z2DyhlDQmmvflysXT+Icj8EOuAPT
U+G93jxl0R8AU0N7gc9ui7vsSxYdCx0PXDY6RBJR+Pq7pUiXP/fmFFTnKcanMYQF
nFfXsWO3ljoTspBR1lMKmdBPVPA1Q6rUP/WxT6wMcu4TvzWrrdHOTz6hsjz8JMk6
MvMxbgSOkyMKsAH8SFzLbJMJgIstMKTOpYzq4SU2ukrVG082s9FPyC3zsoF6oDlw
KT2FvzzvWK4DjzpZ6a/5OBXl/MOD7jfJGKZswNPZ/3tRMy6SV5+gqhs4HzuJm8gw
6HLwiivvPsPK85fDQrX+/FGwbs6wcN8OndBS7uytG1ZcONwZ37wb1tdxf2QGyrVB
bxa4EeKzA79EUlCSUoxQJ/x8wF00hySabRjKszwQWdRgI3MzfKvs0azaRGuP4VFc
4rNvqirxubJnMKArNWl4FoSay3NC6ASsDaEfAcTCzjoO6JGbGa8x7MR3EqtRDgqa
tiii7ua9KN2/PWQy0/NlM/y+8zkwt1AD0ndU9CdZdS+GnkBSc6Lm/eL/WgDeeHvA
0Miq4Yv6LwkNxqHatt7TcbxN5QLXE9XD4JF8m8YzUVajUu0nJuGxgDhC5cqYL6T9
TP/unwDmC2gB1sQsK3yhENMIzLN14C8t++DlRqnXhMw8sEFr4nbnsQfG2ynUhR9C
eL/P7nPyLujJSJmU2HSpEWjiLi2YdEII32yCrpaqRvO2eOGixaSK49l6mdpvUvW3
8Zn+Lukq2e9moYiBJS/KtSZkJewuUj0iNKeWyE3z/+2Hv/AGchdLloUgC1y7djw+
3+KIUiSUzhiTbjTPlTrhBeQm1i8/BAbC75Rgp2+05TbqIE/jjELaCaOEMwj1a2Fg
lZKTzqjsermTLsUvmUztl4zMoqFYHTfiQlM8+4fAyDTl7YCXTuJZA938CrzD2rhB
Pwk3U2NKViUWp1VrvHCJTHS5uozwOo+Ty22nIGzUbPjXpSVaAtMm9at+2jSx7r4S
MO9pfei5OWMjifZZRk7GycdljCjaS184dHStLn0ay6hm0IG8mqGdg2HEGV+pLE0f
snKDkwfX7m5ERr3I5JLaEJIt810sYxeDj9tqVrUNwjPEh4ruR3GIE8s2joOXtDO5
qEquUirdLCfKZptH1KUP1ahCNsqj2Mq3HQmkDmzi1gyqUyUrWWI03NtQjjJumkCf
lSpKq3pDqKSvlG5TQwmlqj1SmdbYRhJ09l7xjGpsetlTZ2GbKdgV9dNly/r2n8RS
eQBg1bD1ReKNA1VtTEhREg+o36vmgarFQOy122so+TlmKRFTElJ7Pl4alC3ul23V
WXOyyCNSqOTK901WTS/yh3r7kcX1tOU707W7JsD9IgVRYSSqymJ221YWNlH+otNV
+ZJBuXIq5BSY+lWT+sNkc5SIdyGLtG2STMVvuwOV6PHPT+VfE20dKxnijNCEHg2p
PMJuoUrqRCpd+8DkfavJ9Y5f9Z/zEvGVzh5itRnAmdxXQ1HQIzalDxblimbgat3h
2VXRMY7i9D1O0cwKHFF16NdukvaGfB/WAMBPNynMb9vdLllHfCJthQ8DBlxTEvSd
y9fJLm2w4H8h+WgvqhU5aCRUcn1QIXERiwJmpf4fPhDGEYhBK6e61wmJhzo+t/et
3J9B7mqdJVdSvIlGHkmmTS5vxzTUdr3QvTzwemik8YLQ0U2/D2sI4f4H4dL8xe4k
S+9slPi5cucNe6+CqUgToEyU9+QB+5Mlsmk65Y3RA3UM7T+DVgfpHvJP/jTivf9G
VSc+ECezZPyi8wT8sgkidq2Tb6D4fAPqqcQxs0/oVEKxHXJmlUsrcnPDZKS7vb0s
AMcduaCVZcWbNNHbB9E9y+0sJ6rNg2zAwgcJn3XreFfXBvf8vUKHCgWinYBOR63W
a02PuEODQL1awHIdvCkxjEhVXUcC1YcARh/YSpplxE1AnbcSX11BL0r9atOg2ckl
fkAAm+cv10AyJdPev/+IfgbWVXv3K7O0Js8tRDtR63xTzuZqiSIGMfaO/ybYjO23
0KdbLaIequiRqf8QcHo/V1t6TACE8j3SO/IZZLcUP7VcolQOt4THxSvB2gKbfMYN
lro7NsSKpUiwsuE1trerfpAJBp5iPG1p8Zi6lnVKJyOfxLx45Dv/G/PjEOQuFfMl
9jAAfmLGym5lUCCfuM0slxQzVkc1wOwmPePFFuQLOtSWtWjQtZnt+0wvMbboD1g1
kMcylyKBdDkK0ijFSfJxfqHJDAQTWWji/fUlH9vOaEAc4x5a8oqRIBJgbxblKCRT
ERGOQJTeh4t7E0W6Z8vIVP4WyofwzvB/frbfPg9gNq941M9pJTnNTE8phSlHy65/
JBPAPj4/uXdaDks+KYyaMUzYjBdwwcicke5Ot55HDbjrEBTEgdq99VvqoiBGMSQg
F8WlSyYKfBuBmJqTAEFkpDs+QNNIN9IEOF/13pHjV/MVvnesiS+wYVzQn95kkr8r
qu09Zp5mk76JZhnSItyWYQp3tCEoiDkiafN54E3FTeoexaswcaz164RQDsGEAycF
JOpJ1g5uXKR3CMtZrvMFcU1bUG4NW233n6ijlperod2ipBgulLyUhulq+mcxVE1n
zvFM/molCZlX4zLLhgV3V0bD4k7ztb0ZoNytEuckUVpiOweBnWtX48uxYhlIdoB6
3ImEZtAgrQtY9pMI+ghecW9g3jOtX4OdTAsy0sTlirmodhcVCcYmMEOAmcFUU6ti
qV8sIY4hSDusbESPB1GEY6+DdmUOZT6viQR7JDUd1U2g+p3uBHH7tk8Z1yTBi87K
pdc31v4fgZhIFjaMeghnQHXyf/ztP2FMC4uE14J9xXgw3hEBlw/UaV6FzMPeoGlG
bbeClNuB2tOD/DCoYKRFSYr1yngED2qQWQZefvzmrhiuS9i7Euztt88Cn1B4aXUP
KRrL3wXiWqG+9B867AeDu5Bru61ldmBqkZ7gVEWRYMCgCnZhzOiRzY53oo4bTJrH
Kx6GK59qyU0zFelesB0Gb02d2CnxYCvLkMzAWyoMpnh7SiX7+Y1J1oN43fUoxVfQ
y7M5E2a8KPwfWWsU8EOUrlQOBojYIXZAPmzkVclkGJ8jO6byuQSFIVD2hoq5KUre
BYBQM/eOeYhgRFdYeCMIkV1Km/IZo9HPVdaxHXBHaf9syDSzflwkD2BW9XfZoJRQ
+kWlaPZxu8GywgE3S66c/Kg2EjEzXkVmsxzIJeRND5BTYi7qZvoHAGoI6v09JAfo
WrtV1s9MCbVrGNRi9Dm5dmCX+7MhrCRwTfaa9T7M9jn8LkFkJVuF1IEX7OXf0Iso
hQ7zQNjePBzUN4D0Rt9IOgwr2xJBy7rPz1fuwMeeGYKKGNW1H+bgdATjWEF5NtJc
y7GJdO+AnZ+rAO/NUYUqNZYwdzZNRkbTHvsy1tI7zXYi5lSiPyAZoE12Qk6HP2RX
LSBiWdipb4JooPlDAlcr2UpnC4ZpTs7DYbwxG1Ign1mVKKpfvxAzXYXZqiREw8E7
YGzdGsLunYW/rArOqTkL/cGgGaL6QVIX1tOFfXIX/H+cIVheDphpnVRq3jDYzyH7
EAPYhsj4zt5p4cmXsg3y2dn73h9yyWV03sxAOCAnm98lyw7Qb1HrjC0UWymrLeS4
TcEyKK+kf8ke+Y+DUPzzZK284uOSA+t3Huejpreo9irBmQ9bzS/ExcwtUOz9jwJv
DvZ/eTgfAMkfBIz1yVyCGgABElXqupuHxROkMXMAiz1Ur7/r6OVZDFaFx1ziIacY
hatd8Z0dThpFI/7tTqCiRivfhWYUe0w4gw0zUpPiwTtrBVOJOkhZtlp1KWoGNRP6
TiKVdVIvPiZcLnYJqP6nCuq3xemjuo/fTmO05AJJ+w6WyiRmXCaJO4MUZDigyniO
NrcOr81K0EEM28pUIYCSWlUz84s+nqQAco8rXxNIt1QYwl8KG0i2VSqWwOsd4eLi
zDkhwiMENvxbyGB2LZ9nfcR3+68dGmoePEUNGZCyojdsdXInSNoxWLKyK5WEdtBt
CYLEvAqOabnlItpxr+8/Y5Ro/9/Fp2fDi6orE70uiUlsw/ser3zTxY0XisU/4T+0
a0zXxTNW296FeZKdolV8VtURFA5M6xdpTgoFqegXDSFTHdHafJC+8i1dKqJdxim/
vuqqDYerTy4GIES34+YTEptnXl36+kbTz1ttZOq7No7xFRb7CKeo0cElsNKCjRy5
J8lIVRrBzkwofGekkpehZCudc9kD9fwalWwP7Mb4KTEVzQsYJcTtNHyj6nDmBDVt
Rd+jdjSILS4anXrMN2GQF76renUfKJc51P80xYtlLYfW5Q7sCJ9RAaqHTCfiBSdV
Wq4d6LS4ZKOw1iiGQb1kv65sPV1RcQoKuaoC1qnwz06L1uHj66RRGcMKJ/REHIwu
+xc3eJ5xc0Rx4J43IwlHnc+E0y7XdY341I7nu8mP4jPnPdqvp6LFRJCWpJ3/Mwy8
ceV4Xu5/1Ntq3pffYb1xBB0LmstFuwdZR2zeD4HSV+MVDC1aQf3P0nwp2Yeus8UL
6xuqN8LOBW7DxAOyTi+bIwT2N9j+48lzfbfH8hmaukughNP7aKyyhIW6R1bkWPWx
72JQhJ35dW4G7m7JiL2DjAjRQq3ErcK3p6bMkoKOAJlqjQNKZ6S17jZeTvBamwCp
qA7LX9Erl5zowTewoMxOb8Mt9kPQvfdksUwbelFFznh38DHiOfm7z+TKmAmo6ih/
nanzjf293kqiAZaQiDJZqQ==
`protect END_PROTECTED
