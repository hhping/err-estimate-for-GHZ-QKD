`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aKub8nRY/98SvdS+yBxHvqQuZi/Blx7NEof9ZlJTnEwO1qtJj/FnJo5BAAFSXBPP
5+6qkLifQixcwnii/nbUvIN35IotzrR4y/pBA1dUDvBe6wffW4W7Kzf6HpMiD60o
StcvXhi/Dt2SE+r8cpZ56r79pAL9TxfqFpcoQHnlJAg1InwUduQ9qZWkbB9vPcuK
+IJGCP7lize4cFN8JWXQmHsK0NbMsR8d1O8+7aaSRLy4YSc5BYXZYXmkkkEJyWoO
8ZFDB3WN85c1OrtbI++VAlV06SgmikVqNAPAGIvGjHnAEFzjY+DfLAw+eAHpF6gb
rXEFlIC7Wk9kaeEmmR3EJQb6uN3mohw6ulDjljXWxQud7MglOQi3LMLoswTBZDj8
ZbpZB1TJ6nVFLczGCXoC2VcSgIJVdbgy6MB0jwkkn13SRec8KqS+ATDeTUyYJydC
io0f7XIpzNsR2sixHwoKG2z5NK1CaRkj6IJHg58QQPDGju3OaR67qJInxTROzYZ9
4C61ZzvW2gd/mu4xjKRdTZFtadaUeGP0hDiPn0r7qExCSAfnhUO8WeeFJsm9oRmL
hMfLUnI6ZHdU/uMzGT+bG9T7jh2dGwfpT5YWEOKZfWxIQpQiWcsqvH1nVHYvrmMU
XitzPyH1oryQQBZG8eIxWdDGY/XRKZjCWx8Olt+/sEHtDegvrUvCEnAyxe+R6tpU
y9+L+qmYckt5HjpW0x3Br/mYVy6VF1gVEJ/S3Gp/RA+mpuu6hIJuEMQQQvlktCrK
7/3UcCeVLGf/94/HDvF22JREmoXED1i44WoChCUcACXp0mr8Jgy/Yx+RO87QJiuw
diYYhQue+ErRcLaAzNKVRs8zpCouJcjN/qdb1RwIcnjLnZ0QzrUwS8WO4ZiVax9l
BijlW9J398Lr5Ia2a0f4E4qwpAFUxkZ+rYZPy0ogre6b5u69iFUo6YvWcFuds/Kx
7utIdYBGglLnbBEMXr/k6MF0UESOhRicd3EKopMgNCIA7YJIaSZ5uBScnoTGZ6vK
ivkMRCKavzcjBgropY4gcfQoAMOJTXUGrv7wCWYnAXfeBLbdu0+R8Fy2sSG3ucZo
w4aPW5sDn5eDXJi9iD1PfCW5je3nIF99rDY57WfObh0740rLQ307tCv2B0Tr7KsH
IkjZEt6vHT9UOUfWJY4z443E7xcn+Krc4CNqyY8By8xHg3bfIugwWZm35uWyzS6l
0gS7tD6NGeW1NjztKnvKdxf+xYKWp0oY9ZGW/Of3KcdQ0z7EBx99Slv+H4e5HfIl
2rZpJl+2Jnttg/KSHt39REkWfv8NiCH4VwNbCmEEDKuF2Qd9RMlpx6O7fN0br12M
rEMIhxXlgJcd0UQg0Fzgp4CJ8Ha6np2bnKq5SUYUtovF0iaTWNTXz2FHlQjs9Si9
H3x/M3ZRCupahBhfY8nmyj4aoTeo1ehIC0XfgQ+Zefq4Xx7/OuDeDrDctJTmqtIx
TR9EaZ9xpN5NEU5CbPp2E2G9EmqPtCDtJAXKmPJ4UnsbN1VT5aCgClbw0lk8yXDc
iMeGW9jhYCFO4xZDLgHiLDpCNaAUHd8w97WHTjva9tljUO0rzig+E+9cMbX/uLTT
jtHvIqrOSkE2jOeJW/D2/gDwuku4smmCnJ5ok4rXV0hyW3wXl6KUYKIlCPdR/f46
W7cxkwEro63yjuphkwVuu0LYcpXnWcR2eDoKlGiqK/XDzIZcwolIT5iejiI3kPkP
zzvTOdiHs7f4MtLstZxot+ZPLSWwu5DICoFVfCwrctUtWqwL7gl5uYmpWr74HWs7
WZwaB39Kpo5L5uu/9xhGOqKJWJi8yfv4fYC4QRefSrYIUePDZgBapnjotJSMisQS
Eyu6ORwyT4MHxmHdyCRj54fNZbbLWGjukUEuWFeAxyQla1Eg7JCNqr6EbzIOuWbr
/2gNPefA7Ccve7bbfVhFvIS9WHtKRgOn3u1KIelKTPkaFsFpHJTgfM6vdDXFaMRA
AaVgG6xZl88iZBT3wldboIkYMh0QhCzuSKf+i7ugnrmGNAyJz+oYMSdLFMj3Uaw9
ip9SZTZhLhmhVMb2tqWwKX2opLHUqpWtReeV9KduJg6aJdPaAI6mh/gid6DZg9mU
UgkV5bp8ZzcpGNz6z7BDhAF816DUMf2vY6PhSVAxzw641ANducJmpkU5i6lNJxO6
8TuWoMrjKNapDlp90vQLlrFZF6+QgOLWuf6stPzyWAZlNpmTnMJBK1gdQ7TQ/puS
HEEwqpiH+Ly74kP9cSkOMXElC39ohK1AVkzZe/sUqSfvWyQTBL0kDDYKM7HW8g7m
OAr/dH6RkXkvfnL7aZVYCdKjz3Rypx01oppWxyU2KYuwgnU/rRFK5N2FWpoJdR3V
MPnIBMXpxlNlsY4nuDB9Em5fC1Y4QhjVDJrni4c+aK+sjPg9rUtw1H0IhgHhnAi9
GJG0SeRTDsd2PwPdQ7rL0ujaMHkvWAK1X4XieWwvyH7AcbR3vXhLI/4EKmEbuN/b
LWaV2BsTrGidRn1Ty8BaJBAcazwbFV/UF/O740DNwK/mHbQOO2ZFd8lUgRH4Yc4r
RRnYleGC6/DuoVoURPQgngbZNlisBFVZjbJrupxZG+YNLkgw1dF7Ptr2WkDdWHWp
ZRz4YZgkrahA9jjaTyDO71iCpiSMbSTqrM80t9h+pLvCSOntXauw8tQEExkkJjt8
WqvhvBJGLK8CGd3On0VIuTK/p3keiA4SJ5mwOHaH/EOG4UDahksWrZvDXNOih9hj
rMcHupzGIVvNmEDJ1jsFarnYLYZgowclkY9iV99xeIQeucZ3PuLfetGp2seEyQVO
gPf2HTw3qGVEOSlBQUSCuTNxV98usBViEjTC9UIyoh7ln5sHmnw3BkVXKEa7vXLP
kT7n6Yr69EByI8U2xePwdBJuRBjU6Y4olDp67NeHbSwH+hAvxh7/mPhUAAKB9IY2
d/nyLW2Y62NLAOqVEZ/ZUWZC4rM/yRxWT+D33u/qPFbUFOmMiqAY/MFr9KKe/F2g
o5LB/ePN5tRfb5zr609HBMhZddF6ZtgE1pPRSnii2RNSa2cXPg1SjVkhYLsCz1fz
xutEvHu7PuTs21YOLWLNEFhUp+Ibv6CSV0lhYkCRz0XTzD2Lxf2mZdtpdn4VJbRF
9/K2RCKFZWyqqZgOm9e9ow72z3XOQ+KcLSssls+eDA2GGj/1gzYLZNXEEBMr5UXZ
4zegwDknX1jiMwBBCNZ/wFh1U0A/1hjR2sg93abgX2Rr+6+vqL22gNLmCG1jIEz+
E8wd6ClMGd+S7iQbCORp19g2NyntULDVin92kJaNhRl1npv/oM9hRY3X3t/RPJeX
TiVcJgEreQbCC5xWT8PQ/gu/0f9WefsOTH7smNjGGce9pfD6gQY4bSt0Gyfb6qyB
BLnWdvgVr1s9D5W7gQgk00uHHvyhNiOBo/TbOz09TWgyF/gv5+PNf7aftPV/QhQ+
978spT0ttDL4+9P1u2ttELQWdiBOI9bReNBY69xrHhNbjJmB374yNMS0tRifQMwS
YY4IubftrjAKcsiC23HMAe6aExb2k5cb6xTPkLJFyXjP7j21zhXoymr3w2tycqxf
0FXNZzoca30Q8uKdPp1IF2n+9jF/sgcDp7BKJezc4vylrMKGeOahZs75Awl/MOn8
5SY2mfwuKaVeJJO8nrF+T3MeUdi3svVM3iD/kWw1+RS51Diz7qPuznlvaRDFiK9d
838Z7Ezq8SSxvf60YELFDoNvmLdK+DB4TKHoVZSGvlN9JJ5zGyZDMBUqZk5OtjBY
b2UAXy/hNavJixLUb/6QDfCigMpH6CjDYsDxheGeQMGsr+pM88BqEdbUGsEV9Rxy
pBXjkTYwMmsJGsvDzSPxRjfk/bHLR1QRGgjsBPB2Ta5SVMxDbnpk/Yaycoi0GjcV
lzmbpr+9crA0k65DbGcMvZnGKa3LvvyxLzbIvQeqphOpS7p75f1yKV8TwHOqUpcM
wssmAYhPussXxQqcjvgwmMmVmzTHpqk5ARQWvNJPYdp1LtSWrZqTV3lj5W8rzdyp
xRR87lcMfLcuSF2sVS8U9FxKuGwV/kopqb0+5B4nbdV8u5kf7huWrw1mpxyojUpD
kW20gnhPuz5o7UcAJWhd+F/21h6WesMff9UyuRNwCbBLKWeIcjnXqNvQ51Xl5H/e
s+gLvRBl+Mj6TOuCJnN1hbWQRA1GDEQ+8q9wlVH/UKmDV+03TTGPMcFdUvgaCYVG
XUqTP+plwvJ5fmC+hL2zc0Q2Kf4th65JIyyHEOjMB9sPzi3WTEWPNkHqkmVTOyCB
VHDUwvJbprd9VjTPAPJW+0Vb4AUirN6Hug199KvcziWUq4iq2Yy02hHLBDhwYVG0
BhQjzGSlI5V+XUho1yNnbHmK1ud2nonmpGatltyIVJ5EiKiLWAc2xteBFFaipZnE
J8jfwXbTc6c9hpn4iDLUnZ/jcl8cUBYaIkGAlrdvE2xP1oiYeKG6t6rfiDOJMv+I
5t9BT35hsMVmVOQOmeIthDcX529ajzmYjlhwGZ0MmrN4cEVhgufu89uzJo5eBdWt
kyMSReheEywJMx5FGIGkCP5ILbImRGj51j/0tZihoHZA38geJjSrl0w+p7m2UqSR
+SpQYwPgrii5OZRByPvgUfwTP2AfAubLSj1Hk+sJ7sZM2zeIm5WPq+0CS9GdX3Ln
yC66dlO0TmWAH2Bcpyom6ABGNdwBKTJfmOWgTI693Ru74wzq5rxrDy76wG5sTYXD
/jqyvvnQTUB7cXJ+vBZ9HtEgL1WsSYTUF7l7VQLiKw99UI9FnbANy4UUoPwRDB7n
I95XIMO8pTLDTZnpsZ7jJSvPZoSAcBnm3Xjyal/cwf/oaVIPqLsAEFsiLCO4ekV2
hwoK+l806V+02czE52PHhDD3/j9xaMAcLsE6HiTnRqPxIhcyZV0SSbTu2dRTZgCC
j73Z1gyE5BOycf3cqlsK6Kqup+kzpsIEfI3VrrqhaXiRUXHeiyjT2lC4FYolwo6s
nAGAkSfS+N8s0z7QPoOLpIAM5SjqbPPPHIMMD59dG5+/fAPpg6WKrFajHnYHaYOv
QjhknsulA70kN+VMnMmIvtIRIx/OP+xft8ahPLZesY2SooLDkST659SEVRnpyotM
hRiRoqoPY6ofqsuYJIh+8hdovsMI/uddUG7ZqW5yD7eLK57z0spQc5IXBto7SDdE
UZHH3UlqUIchxiZveaqxmBdLkNu9w7KQ6IG+JxjdmpcLngIFBO4mkBYXJoJrhPCQ
3MCTrYQPQDap8Ru9n8bV5O+MWbbwR7/mLW8UTcuTIeHE/ouab6YMPhMc0P9vXxKV
p0v6md2rw4McWOlj8VU8VuMvnjIDWO50JD/LTIXrdzN44kNIAM4ubjP4zq07zzIx
pF6wbyr2a0TtfR66xyWPsqXYoieNWoUp4+SXSWGnB3t0lrsSUkb0nu0gASF9TNtH
Mo2IQKTmgoR2ggZIpaqaSRF6dx/2dgOhcRXF3I1lIQyUCa8qGQrNGzQFoAFfkSQg
yikLBOO+7X2dgCdl6cBB2iKDdYkoY1uX0du6q7qsIi3OlXdjHKz78ssI71pZ1DwO
NO4YbKZBhzpI+Wkk0CF/K5qvuLTa65pDNqPJ8gGAZN0C4AtRmoXZQfyLnFs/tqgO
U+hIuwm8DzTgCg1R8YYR0TALFuCTYdGgpGkweGbXuVmGVuZFRMxIDFSlfJ9F4mwn
nNygB+Qpv6553ARNgJBLHLBw7wtzthy8I4ICVpFC9wu4Zsp02vOMOtmI7rDORotp
cxkxrMz3j1VK4vy1YtH1Z9cMPUnIQCkXMCXkNKDKCseZtMkHXPKh+LIhHlg9d9A7
fukUYG50cc6y0nTz4OKplq/MdBED2CYbaMFTnYdYT0ajN3knqodAH55de9RXE9nt
n4qaMdvICHmYDAu91L8ssz3B7vr/3FNs9F86QPquPBJwt38yvbCzLb3QzSTUHzj8
wXqI1ik+V2nnst3q+xw0Nve2Yl91SotQ5f6u4KCvKIP2keJDtYWY1Y9txzzBWwRG
U7gz7GKZbzGm58E5pVBTG0Kf2/r4e4XTWx81wabA9R9sBUAvhWC8L7rSpgEP+KBy
Im2lrAGt/9Amu97LnBC9ddxwnAGJ3zBzI2oZ79+BNTzQjomhpDYg4SYwLSsU2jCn
HHUZ2Dd3SfOJiSKqk6UVfGb4+z/Ld5Xcupn153ynTpy8MundlyZ0o+Mnpzy5med3
J3ZM3yM7rrcSdRe+tsGuXC8gP7CfbXGv3QR+v0WIEx/WPLrv4YgCMB1lTch4h+j1
Q2kbk6wkfhiumJ0Xcc92AOUz//CPaMF3yX4tku5WIX92D/nTiTayAIy1+Fr3AExZ
FnfYqMR2pa8iTJ/fm8yAGOUtGJZBay2E24+t02ECLS2PP6cFIe27om7Z90dKEAzK
DNmpcX8FANE0MMNHl/EIgAbvsEi2c3LXMxbcxfATggXH8dCwDTFAbSEptQCA5rSm
VkVYuezW5nv3q/CUl4wMznRJ2lF2qy1TNJbvl2A0aCSZ5cKpSJn+FAUTLQ8m/SIP
w4SgG+qOOI923Elq1OayETgOFEg1qKWLJ+nG8GL3zmjKaNiWwzeThzK+Hhh+Ludj
758N2+e18eUMMlqDpTCWxnIq3xPx4kSD7UVBgjHSbLY2fP+E1CTP2BJAkQQaSiRz
sISdl4wxY6IxeDVtjuCY95PZYtec8YewA5yd8YgQlDOyW16NTSUCERSMwS5cFvRU
uZvLKGJXuOPC1o+BxVvnAObF5Z/E4Lg42AT2Lv+twBITfMrQbVMwKfmGvZP4wNYx
zb6Ol4wXOG+Fjz4vpjeFjOjrX+YocMCud99L+L5JGB4tAjuJZ4vDQlw9RpsZ8SUl
OvHG7JPcL5L9thRlZFFKa8/I0cJRsvIJbM2jU//6j+PHRGCPvu7aBwOHyrFpZ4UD
4+krD/rTsOL0GHdBULwZ7ZlgGnajThdKKLDVS6lbplXjq2Iqw36pF+bEw/LW1TXO
2CursUC8jte183gkukzS7VVciKDPT28vwf0QDqOpsz4YGguvaBw1u/f6vCPoHNVA
2WtSHVzOry9OJQ9h3ryGatvGQF5ZdT/G/zNCFqMCOINtedbLPL2+yDjm4nLXmdCG
ukH+je7rxruy1jzTs0NK0gQOU01kT61juPlI1LK0kkinHgYHQh0Csb+CwNU+EQtc
6ZdkNLcXEIRCCBTvrscMywgw1pj4RQXyHbTB+Vq6+TyQZtNAiCQwGVvJ20aHVcZ2
pjQufyo7voul1QDxEB74Vw41edoO4ZxmWwDVrHEmKFYhnWI/vXsswGMr/82m/FsA
vwd1ShoXHrK5MuNxh6+rwTuXqKG9gynjXBX6VCJNO9jmdx5HMf6ggYnIlg5rN3P/
hHMEVfrzoAl03rx0HrDjVAqCMPviUyfNgBJAUFAYffMK8WltKJE32Oex/7o79jUy
EZBgyS8KZe0kuEVIBwyyeRBHTspGNFnDZTf0qs9VbTq54cLsrqWae2b4iUYmH/hp
JgfV25j3LKuQRlgQqt1ZRX2BVB6Gemc3Pnyj8Ki9/4TCNf8jPgf37yOY76mB5KWd
6g+oERhUtNQ+8Ef1Gjpa1kpreO5F2hajQFrnraskb7JHOmZ/ybNaN+Pv7Ukpfnsp
rR18rVKHQ1gBpAYlkhA60z13g8hmzXApOYCvFVENlQgJjDFoEccaiDjmPpyMOXeY
488Q1QBorO9Y39YfZrVnVQc20jXSqk+qoG4rOAwbEa6z0MMULeBpYyAQZ/DNu92/
nwbsL+baDWTfq7GinCVKQGdrwVoTahNJBICkiTMgeTPX2gFM5rDtq/ll4JxkC0H5
tOuMjtbxztLgPNg6j1zwnwEsJ3XgtNHfjJbTQ3EL9fckizF5qFuy0A/nt2UXLqTG
Ke4kep7qehbeR4B/Y4rWYtZ08Bx/PO0GBWhtNQX+F/CH+xqYHzPr8F74N7IeP1FN
Ml0LNdj7yas2fHXiJowrCODXuzvJaNgBReXKtkDKiY3Ju3uiAOySN4XI/ZAnhpvF
Kr7cH8buvG4tXlr3qB060rBdTseH1tWW64uvINzpuBMymvDFr0ubde0BpgWljOoc
7sHaZjTGo20uzygmqusT9YTz18y8YZY22zrGrWzpinP8M6EQBQ7tZESCZOXP8Upe
7iQ6194ihPRhcgVGHfmXajjmwE76rCj72IEau2xm2Td9p2UpOQ9I38PB1WTG9eiz
2h6L9MuGMzkv5XSTEz8E7KuUUTRICUWqykx/kMfKf95/mW483DU28yYlyMLXE6aI
Q75QyP3wRNqGfxsHNxfxBFWpcAgFpehdgwthENcomIOWCWiS8Sdrl8R8Ljl+tsxK
Buh3tdMwiYOxdxH1uZRcxvb2MrVAmynfcyutU047gMLSvxeh4DQUz4nnKmivGbqj
6cCxE4+TbVuqrszS4gYff2YDkcLHXlZo710Ujm9VhwKgNpLJ+eeB+BidvP/0L9c3
wjJDvoVpfXjRg+dnMo/Y+muaTSk846wWM6oj2+4ic1HvNEBYP+JzOxlYos8VFRnb
p35krG0zoZEurKXlSbXug5WhMqk8Y2x02od3Jt2RSjvNMYKKlNjV1D9+pKTzQEIc
N7xIEXnpZbh8frjpQZt0JSr1Y1n2s00m5QMAVrj7cNF8zJNhpP8fG66VrsrcaqLy
eU7PZiTYAjirnmRw4uLTBJot+WDzs3R1048p0XztqORp9JnLKCUajYoWpgxbVnW6
TVW46x4eu8F/+2VOa1DsSAGqCdahKfkXS00iuGpkbGc2gOHWSMCS4wHKix0ey0+S
Q430NcZI0QBAzi44xGSbqWgM2QXVzC0Q6C+Bcd4W9E+JV9IzV8PA/UajhH3THL6h
y/8EwWeHbiqcxtP4tL//vJ/xmN6VL9PwPuwiO9SmJDtl+qM4zCh61LzJxKs7eaZf
xewqpy4+8qMNIjc4U/E4jSVP1aWtIXfhqwLD26+5Y+2wKuV/DJ9tvVpc3AZtDK3P
yGhKX6AmMhRdFJ7TNUDdmClusIJ8u+QTk1LJyyYOdIqN9FRmNsUNsf/O1aRgR9Vn
l7WFRED2GubUm9iiGffYUHyUthhRBW7QM1gr6D17UsPFyd+Qx2AA3cuuBij/+McQ
TTAs/zJGVjwa2QPD2Ina9Aj9JaGG6BoAnqZRA7rC+1QDHsshN+NR9YVqI9hJgKiN
hcedrMt7L4ByqyLHlbeixTj/51PSJEuEi6wgmQSm/FjdUZMgF8NvXOTT6tJ1R6mY
RW/FEOfe9r7uuCY/XpmAeJ8NGI8xsknQGGp9PXdThLawgyb+LpHJpJO/0qsTrAGu
HelhJrYPbQHb5tb5mI3DBJZN6fh1r/JV7BGuGjQ7jtBoN8NXM9Kglmtjcr7I9Mma
KuixmzFcJxH98rLAuQa7mErIMcP907VOZzcKNYQalxLIFFlvqccbIDzmFxlJmFkw
fT0WWV7Tn8V4hkBOVsGwkdNH0ZetrL+4Y2/6duRToHlfzv5Q8auYpNoM2LC4r8qs
PVvgnZCctgqBMKuS0DwFq59O7k6wDTX7sIxQ2O7Ga727+hbgoADvX7tDYplWK4Cx
qU8fXY3FNGq7E741HMQKi0a3xH8Fu8abGYEXuXk7AZrvx6DY9s9rX6IR9b7NkeI8
oxz4C6YXjETRVKIDGMVHMwBzY8AjweOjJbIlOe7dcO/HPojEacx8t1kb3fL6ktni
7ICFwyFPtbAbQa6Bxx/qBKVsnHv53qnjETgvO1QiKoRNtEaexmFV3FoYJk21iyDu
alH3tj5NBG9E15RekZ4a63+vKxuhm//Nubn5XHcf63bkP6Wi6uBJ6xTcQG3C30Ff
PJTwKQuePOePW3m4OfcZdtrbfcBV/iS7RtP/C9UesjAmGBsquu3wQ8JINK7lZQFy
7UFkuMvIWxMkFku2BhSL1KuE3SlIV7aE4n/VZ+0wy+CvA2L+OXo3nuhC9DHeviBY
jk6/ntW1+IpMaYEuC0cF0uxhKG67z2ChpWl1l7IMXGoHZzHdEJBgloeAxTCHqqpC
cLvHLspjmTqoMHB28LWy+1Tiz8yQ9VHJ67xxmU3Rp7T9KOpjZXEYYmsXyGNJ1NA9
RLmpePCPTyzyaDSXrdahcsMoKSHlBySMWqyb+TD1EjWWtHltpachlfOADnfAw5g7
3GZn8v3goVbdvrx/4cNGzWJmaqz5MvDgyNa8YnJ/Etnrsh77Yh29hTRUB1xvATHV
78GBoBvS6gq2S2LO9wiENsk26wKzu47wNmBdC3zj30Sk8TkKbAzntsg/C+FIUrsZ
EaeHzhzR9UZSxcUPToy68qapMJ6Ia52SYplZ1IBCgDRG5eZGeL47cFIHsyRdAaP0
8jjl+DgNtjHLRtub4DWbtMqiLL3UFUZawb9ZkyV78UhRQerz5rjf900jGuQJYPSJ
F1dbAsxi6OijKSlxYHlwosd7Kp5PgREkQEA5+x1+wmsqf718Inzbds/aAuOhT1F/
X6c43XCL22wDupV4HicrMlg5w7rZdyqZE2qF+K2SkpWT0L7Hkvvi1g+HPP+4Q0Xa
DdM6+4o7PoUrnY9du1SiK3W9vUhJcmCg+1tWrD639q6rHDPUtpohRiLtu5GjzCm/
bNgWMkNKK1iQpgEm4MwSQ2GKtY80og3U67S9hTMEnT4HPorQRsB8PSfz8SyW3vxA
55Vx+S2hBX/gCJpzWXnT42PoNrD6gnWBBtnl4iTxL21qA6keCrSfkip/OB+00TtM
dFBz0Run7KR/3M3PbEQd8jWeZe0U0+/Na0hBGQ+u0iH4vaVB1yLgEsfGh/vrR4Pz
bxRBMJU7aJbRuWSpv708C5Z1JykmiNTxK+p6UL19bGjgdgb8zU2nRZLYvt3RcYdr
rOU9ht5soXloQGb+WdgL5Q8ANJhX9NOgaccb6fUOSWocWwj7DXjI0bMpcC+yfKsV
fQ33Rf4Kl7O9Pmp0F5mwBud14MxW9Wur8pRAVEF4fqjfDNx86Ww5I3rsm06Rq0I7
XKADbCwHPj46SGfe0YWMfrykwCcK5XHCpNm05l1AF4JX+/Wq7z7nYONsNjqk2l5Y
QskUk0LEnYiS54lYYsekMN7rlpXVMusbjr+JIgM0O5AkbwGBo2BJXS/MyTKIrbWS
owuUgfXUgBcU5t7sRcQ4NBI9Leqw/bniX5GyvNc33tR9jBNXnEBkIjsOpaUaEgYl
AZ7WHOL9TDPTDgd69hVEQa+i1U3w57Xkep9v0/7xOLRjCeFchyTboNn1fQGkB+gB
3Ce99DpGvM9DDUmV9F0kMJFnhqq6KJJh81l2jqX6sNnbp0fHPDvgpmmEbughrSGE
TsgjCMaxFED0rmHxBluA1IW1eTXjWTzyVGh8xbi56iTAuUoTDYFG2vZmatzx2xMs
GexLaCKRp48P+v/xuZCx+apKVaSht8Eq9p3eOOr4ZA6mxoNo4OiL2xXfWYNDiB6/
bf81im9Hf1rBKq4ZJnhcie2NQiQItfaaIV0u3kaq1WW8sgqqgSXGxdMYTfp26wRc
8/0zsGCHcqNWEnXcwkSlU2e9JSIvJCBdU7pzQuGu7f9YixpPOeB2iJnss/F4iX0+
vKjnEhiA32YY7oZ5Uy+1PEYjC4OHpOHqJo/QdWn0R9Z/p8T6pdbCKiNc/ej5cODW
8Z6+hznp95f8qObWjDTBuj6Pj2OLkcB98IwCEr2ZWt7XULe4d6A959XkApbGWCFY
9P+K8RZkxK1fnKUm2Wqk/Qcak8Ik1RklL3oNDhjgabpdHj8tCfyGVaXmNZAF43pd
qkhDLqu1+uJ0xcoYENq4rOtaAmPOP8nymzJ1HKBEEYyoyWy3WK8BzS5bE2OJXXxl
Lm7g1bX4OATXrxNj4parvAUXolFg7ABQGYhm30/a8KldLIkE0X7XICLOZiTbdCD/
GZ+VT6NNmYpWos5+tJqSe1p5JlrOsA87sm+dnlGo0+/Q/GLh8GmFUtnvGy/cpmvO
MtgAF6PxQNH+hRbs8U6iBJIpN9IALyA0v9seusOEbbGVcPZ5p3/Vd5qBJt+07Wbh
JU01bBaqhsTTTRZ9kxMF/xIW86ufzRa9QZTS1JbudwjB3BJFt2/wOI+CugQ2uD7/
D5VnzS9k1FHnyjWMhk5p/tu/KTu4at08VigzDEEiMhzauvRKjEYaBQgZs5Il8d+i
TPFYt4JlDhbsTG9V8QIyQWO7mnMBSIaQMZWxva08AXZH6o9RP8ya3bzb7qvuREKQ
4cV7D7tBStE8f6GSPM3dNIpc/hNkPcyAZCX2TY6Yu+kIq5Z5UmK/Rs4qSGMB1Wdh
+h50mmlJLviQCAPQKhimqaOfMnh6Bh8jy4LAFmDIlWV2E+l2z42nCO6MAYKiFgWj
KkTc0BpNVdD1vFzLcwXD1+xhPJWq1oqQOE0l9zFAdOFZlgUa9WV5nT+PlpTy942T
yg8RWkBiyh6X4JLnrhmf/fyDGODZwyf3Nh1XSKYP8DV6JOLVeJQYDanS8zNyNU5m
wNgopoLMmksTy8VtlLwBUlD94TG2A8ue+5KB0+Y/HvTQGZMbDp8Q0/68vv75wglo
6Cx7jpNXn91ERWRmWkFUmQfuA+Ag5PVWIj4ws9ECcVkq40NnOmYm+hxdPdgU21NM
VSCyQa5JeuWeCFngo82p8wvW273MZd77i8tvVcd9DXzOawWPaqTIo6n3LdE2yo/k
N9p81ubjWkIwL8efs6W3SYbdLO5TzbRbAj7QagPGQtDlF0Pt9UMGtEpFx3K5eHZd
TaWPPSWBoHHo0k3zIVaY2izytzWbCSSTChxg+AfcpYdlC484dJc73LWWL8FXbNzZ
RKFDlLKEsi1zXRWMTTtFmWqr53riqI8nVt+UZ77NVS8voHi93jS+EubNbqnXgA5G
i051cWNz39l/cDa7XFQF6eHVwDbHkTKWOx9N8mft4cfuaRlQOmqmhER/aZc+Ivmd
PTDBMgVnVXf+trZsmSPGDkS352TWRFOx3Hvdrvld+C+iv9F89OJKVdfE4Vlo+YTT
iUMo1VOwpzMpspO48fTpoWhUHdHLNrkcNBCCZPF7L8+9oNeka97IzL/znuBrHwyg
wYKl+GegavNQhG5CO4hzvXW9HIv8UvdJDXXqfh4l0Q/OBmam01Oxme6I5Z2m5lE6
jGgFprbgG91tyEpuRq21sbzLF0fETuu2VsF/rzEmxk+uU9DoPUj3ozIFYz5Qcg4t
G1363Xij8Kyjpmpi+3jb0kMu1EQZZvnyPI4Gw0Jo/bVqV6bzasPGJWt8HMNHqcYU
uh49Xv7wqihoIc9lt1UFMIrf/xCAjdkpgDPTmAlDe/YdrwSH8Bd1RPahhFAcqq1+
lK0sA0XFemAArigwLQzhAlYWGx4R026d4WetOhbJ16MEdwIb37HVMJhQhR2f1hxt
WdDwbmCu+ZUnJbJZGSIdiY4qv6LI+iT7I+HJdPCiG5Gbuh3GrqVyv0Iy+09VBUyF
aS6S66v2sp+5CtXLIwIfhPqLL4CCcA6qvJvGAU08Q5RKwkosQ0OcII49LZGNJxR/
qeXM6KfjXx46AFE5Ya7ovmGNoVuPXxxYSwGh7uO66rszdExXqtCSc6GCzegunXHl
nNNbwHjBeEiedkNKyMWiql/H8ZmEV5oN8ABvQnzTxq1lycCs8ER1yO1dLH3T2EVe
87GhJsaP+qUBK2jeXvLGgIcWGu/lWTNiIG28zsAy/P9mP1TvyY3ZfyrL3MqJP7RN
msbNaIrTbrn7YEJoNTwLe9p6IR1bNOMCLTU6sfatH4KhnXeSV3R00JE8EJN1IRKY
QA+akpbVhQpzXAR4UJIMQhTRVWaOAmXxAgLTTSRRkmIOuJyZacFAjv46O9Ijem9b
eKe5fhDXd54zUfMOpprTABzbcbPTNF2w/ZRtTR5aDA7EWXhbGGgcwy7CLFRwcThu
5K6JGoe2Bgwsg1VZKwwiwlJ39g2ejU/Vu8DUGkvcEFH2nCwGr7KtqiOVH/i529NS
SretAFbMedw/jHQa1WBo8SnnAdHvBAJf14Eq0927szCQ4FEWhvNDBJWq1i5l05np
gFBYhS879/4s4ijn4vcvfH3E0xL1pnj4uMd54XOQ+Bx70wxJ6rCReH0zPvehbWSI
gkArCtgzrPxEekFYd+wi5EnS8l8rqcoCrMdDDPJx2eHSx87etR0bU/tY4idQH1J2
ang3ldqH1XB7tPSxtWYUbNkfcVObC1dA54bZvJPxoKGjKtXSeaTCw7PU7brZ36OH
9go0sKkNtlGMkfKAVXThP/77ad1hKHF1vbwtOPZH4fW84lJsQDI6vJoCkVvSL0DM
bd+S88lSCJCdCK6F/tb1SjZAcWztzcDVMy83PA6TlytkBC0s/xNu9EKc/EvjBAfR
iXSPoHdGJ8OjoQHB8XCcgVS43XcM3SLQojr+OjdSdX0Jk+j8We1CUvnd5S2nU01x
gWFn7Hd4ZV/m/QrovxMMkcI0Jeu6oDNkYrSWUZ72v9V8DS8Oj7CenrWmf3cP0xJM
jyR/mjchiFrGBP5Iy3XzkG+BpKaQLu2Dlg5woj8WqOPF5j1qcA5Ed5kii98KOz8U
hvU2jVBpfSEqKiClOXiD1ritqGUVIAy6E59PKVK0nj2nRxpAsOBNTkTlIPiXSMJU
ZknJp57ogRonY88+83LUlxY8OBmq/vys3PZ+2uTesI7vptdybzq966TbQ7SY9xaG
3KB1+9A/xxnhnsXQnQ5sTwibrnnybpH1tXkno6QEAX2F6RwZTwot9JcY/ZOOD6De
iKHBd9hlf49Ug3mHhPjJ7/gzU7omU0oAV3iQ69wXg5TDLU4N4F0jj1ErrQXi0m6S
tiHkzq8977nYPSHS2oF6JirLs/GdhmKJIQkiinJNqL2Dc9Mzmsbd2/5IS/6a2zk/
6XkKUTokatehDcmSBrJVV4OZC96N6DEcla7UUExDyjiNl99nv5owVuk/+KXYXdcB
5Tr32brv6esZZXBompHgysOvlC5fjmO8VLfG4NsRwZZyaLEqM2ahRmreIo2PDXLN
1AdNpy51MwIxI7Xv4RlHXv+3dLwrRowsB60Lk1dRlpePmCjR+tjT+NZwwYXkS8to
3sALvqeZYNPEgKTGJATdhkHaKyQdzV9+yCVlWP5OeSPxVeadPEVeiCmSetXkJY5H
D5HKkVc1oZFJ6CzGDOpuiyo7thDuxFlDe0wnqSkpp9DapkiD7Q5atHyB+v7ZpTcL
0nS6/41CkrJ1lIINi7WGWEWFVDa0J94uH6QB66CkcXD1u9vIiAraDRMT7SG2ta/C
Q4VXnQypOhzT6Ime22rQdGheL+4eazmzDY5UKvRB9tBto5CTIm0XKcIqlIrrM7TX
hb2SSCoovNL1ByCZp/0+Y+WokgtausPoHPhop7m9Fnki020dx5NO3I5L+yPAf3bL
lVOF/icEE6ektuHh6+fbat0a+vjUAXOxc8ojmOO0Ib6Xi0lkAHPwuFRpM/KERfiM
CD/1tjQEq0NCq0a7OHZEr0rat6ue3UrcUJZh4GSgVoBJIXSjpfEt8bRt18wRmoC1
5jEpIeaY4MfyCqkv3zZdvTgb9KcmUHAtkI4RZl5GykoM6P9FHfkpLC1+54Q4S1F+
0v0wzjrCdtfuMCUjMwC+k5EQZKZkF2oXaTmG0D/vFm6Fa65s3EJXTjfJ9YP8icQq
vqkYuQz23jfXmJyFm4rbFkjwWO6nW7Zz+4sZ/HfNqVfqI6e89kUsWqPbfR/rZmTl
TDAfdxiKq/bUZTkQ8JLwCu3zfy7kdbX5u5LzMsF9wVxgDxfuPMVqsmx02Ammc9oF
x6UUobNZinmc1YMilzTeYJPiOnpnZzbPo455w3YPz2PhuQ25dzO6yOgiUOUbCdMh
4iV9ej8bAuYhKX7ZG6eb7CuhaiXyGcCHJgGHk4F/vl+T4C1lIfs53b2x+HX3ysrv
185MiOvc+2yQTBVtWkwtVZpZfUnKNmHJuqkm+Hakau3bBHS6Ti6X1HbYV17rEVzF
djEJPuE2L/olZQrYQ7dY8C3xV7IAvtnI7sfcV+2/KCppaSfViafWz8mGT5a1TeyE
PHCaYDRAOsYOsIGe95SGj6FDcnJUlCfDgVpKkj+OBQx9ZyI85SQByQpYiap2/LO1
1O9gQFVTiEZq2WicinhoGdQ/gUObW360rqi7pYWRHvMjkYmlYHNrQJcF2dImj9iM
6it+QQ+GievajEv3cq7gJJwgocWrpDG6Nn+jPzQR8nB+R5vlbKlnGiE7KMXtN2dh
lzXkvC0rrbBXdE+43NmbAk6hvzBodl+N07+TjJ47fhmGkAXP2iUxVutD8ZkLoGpm
VcfqounFMpFRJ2c6jJvgRzB5U5Upf2/cLzybawH6uh4mLb71cGNmpeiK109PPiSF
nThh/t74uWPlCd2lWQVsv431/HnU2yTyoKiBy3mZiFRa4yLNB1GH1TUci6TXp4P1
tnf8BvEFtU2elPxbS7SWzVe6M6VhkgaQ82IwVwRiZKoGhnoe6PE2oFC2qaZCfrnW
2iUJo3ySxFx0j8NgVkveWieKDy6IEd6+2CFWfPgdCgmRlUwXjjMxIMOqeGdrF1ld
mvx2RovQqO0dXOplQoZzM6jMDHNc/xhONsrD7rtpFuidW6IYYve19JiikjGfnwRV
cQRmdxbfpP1WugC6ll9FMZ3djJWGIHuducpO+Y0kMaHE5AwB7HXWennEphGcob7h
SgmLI874ERbDcwuzdfRQRCceQp9hquq4rgucAYWzmmJ9OC7+spYQmqlNXwJRXKoR
X0nKafs/08/0t3GbxoBYEvS8y6rdXTUORSRrIqXj4z36knNmqW8U3vmFSvYy8i5R
jAwcCo71yAOPvL+PuMea7dHF6AARA7jHIZjRPcq7qiPfSQA8tmNybBrXfPuQBK2d
5hjme9bmml+HA1cVhGXYMuyt/rbT5XsHMmHEZaA6/MfAjK+C62Ma6dZnFtrKmVYU
mYX0Ue7WWW3kREd9JhX/s7yr0Rx/xcPX1AYyguv1BqyD4C+4skkJOM5PuXRUKNmj
YfUqN6OMZziIP7YleVkLKZUCCO8jWRkQWWr85ViunD0qw5C8sgHfAV7e0DRleLyT
FgJGUmt2hhKtt1KwturYeuOY0Nf5J5iZqlHhn5CumANOS4jFuRUlCNO60L1ap/FN
mEJ9XYthAF1CGJQaD163iqps++MKQefdLol8OBmeDBtx/2oJvvh8yMLys7Jq3QFQ
w9KyDZ98t9nul+G4p/s6CmxySPMkOi/RvWqu4O6IY6b4yUFxRpsGERgdrCiZ6Wqp
zo+staHC8Z/LFMbFKheY+d+1mzbXn70NzaFHjxbLzQBHpKn+2tRLa5SW8N4PH0Q6
4YS/xSQSULZfUYZUarcZJW+hE53a/Yq7iGXyKOnwKaHw+GgQoaqYuNcIqyGh/Tv7
NistoD3rzBsiwFgAZOMMYcx0YKSke+FcNdXj3DgTGMxzcKLPzUWYKb9beBauFOPY
BYKyWQXMiTRXJBdkWjEjEhJsgAVAW+l91IFr6A2btj+HZO5QZQvtoZwm8uEdV8Qt
mu/mnmSW2XDMrpUChC1AzddXRojXFiWVZgXIz+L+4h5b4UkffS2Jx/j+Zz6qgGrT
RunBopLpa7EFVbDLLiICzKd7XLgH+2YmjDtPXMqiy7xM4B3X2UCSByw8GSrBBoU0
NAtXUHeyKEbld6tu1ekIBNAm47GAd16gRvtWJp52qwW7KZmDwMT5rZS9YBq69KkI
CTShgu3jo2Yh5T3SoL1V3BdRlh0Fy5E8Cgr6/1M9pPMORbrzqhzNVrWnxKBNU3+b
8F9NdtpuV2GkQx0gi72ZzRb78umCf0txwXg9MEfHJ30XtiyYLv2SzkC5yKGrnusN
Wb/eVcoJRFAvtRqTmU+2zVxD/dDalxMXQ/4OlIFSqOJPaL4IRECyZqVmO3rZJRsS
ioAPSnVQyVQq2khP9EtcEn+wL8HGBr+xdo9X/xL5K4rcY64wEZwAj9g3QPSGBwx+
X1PykTKqP9slInAPXx46vpzfB5LKx7tgtZtl1eW1gCDPkc7GZgk0QlVpNOKvOomT
yoX9UJwtpnrQmAn4fy2IheTLgzBiSnbglT9gWeUeC9gOKBC1QaI2Kez9Z/diR3ds
81PF3knGcaSzZuKIy283R/Z57bP4VdNpNAt6rojFG01SHVVVT48TyLLYxV2gKUE5
sCQiGjmIW40hjzZfanXvaNEMdpVA8sbpYrxLStUSIpL559h8XUgPh+ug4Nvc5cgh
WLuNwAaWHmg7QAoy6hymUgyS/gatlHkzgTiNjEm6K3jFuWDSNszNc4PLKsodFs+W
SLSjs7KseneTw53YXeEW4lKFB2y+j4f+pl9/dFirWla0Y4WssSOhPfdZChjCOyjZ
+XS0tt1+PLAcKaLiu9yxRzS71siZpzFldYuuljHfouncsBgiJRqrwSxAAZe83BEi
ugJKGjbe6/MKfJXNG/QXWnn1PzoXWUKdATAPiHdqzJRmlRiG+R3Yy/5a45e/jmyq
ply0zvqAHJDtrOfBk4a5WXxseh2FIUYLCQ2PY/EKtpis5vLzVPZodWrNI33O4rU7
HzFbaI4zs7LDsYxsQBilQMZqec0y+3G2Va9Gqb6D8QmHJRCMYMsmSujvjVDp5rEj
o6mExwGkmOLJNABDW2qtcl7fu2+kk1ZSSoMlAmp63+/MtHK1IR+5Z84+tW8XPtAz
peeXbdqVAbzM4K8mMmQ+rMvj/+nuPEmYhxVFSD89kvszV/vC9d+atoBZjVQNVxMo
zuwVmYMXaBKUHZjl+e3R2w7aYhV6xbztaBaVEbl4Vn/lZ48Pmd0J1Yn9DGbhIqX5
wg5eiTcNCM0j62H9PlkNIBs1WtAqM5/plofzo9BXz8+1/Oxp6Gj1phwAOBvEvW1A
K63nUB/QesTWPZUT9uZaNPH+hblAy7D+WIzf6OY7zecpKUY+5CPaxi/sUK5S2r+t
ebTYfqmXI5ym6hf4YljE7pIoROIvbYEFVUCUo3lFQ67WmPJ7G8oX8pwuIpr9imOy
JAZMq2XdDZDkJsaM5WtZ4TVg7a+J+eQZs5W6Ij9nr+jOkbpgIGzTdAH+etiZq2eb
a2ycdQl3v0v3AWAHZe7nhIdSIIsFM1eGVKEK3QULNRtkiBNm3uGg/0DepPzm4kZT
4zrnGGilDC47FRx2OZcWrb4HbVrCN4gaSqIICi61c1wqJRkBHWH9jUfpSlTPUBDq
vox0WIaKPOuxbVeGjcOwc/UpcIod5yEy28Rzaec83VMvz2NOA7qsDy4BepgzL6iP
5im909me2iPuzMLue67UskItuxuA7j7U6ClfW6LjRX6AuWBdlXdOWco59XbIM2Rq
wo29uoXeq5VHE/41tRTWUtVKf1j/3v95GQARNt2ilzXo27+Z+ViT/PPwLPHbxdfk
9+ErvBNv8QS0aOfhSns/dw0SZu1aDEogR4IBKzj/+gPoAuVdJyrEMPLwPvNEJTzp
UwL99s6BbhcIYhoVVOYO7OdV1sHUudXX3U7asnnMb5jNuOjqLvXDsECV2Qxvu4lo
KTEFToHrKyCxtADNKsMy1dyAA9u3tg7WLEnL4LSqftn7YFH/bWlr0glZnxNCfVx7
ZXEtZ9RZJ0/Yy1Cbf3444iZucDBF1SRBcQCSDL8PlBXZX6hmmXCWiNTOVjMRZpRh
J22BRXkvbvjrjq7pO/y1mJmxQ138l5T6ADe1VO00sutqQ/7kpjoxvGTMbMboS+p6
ETNU8g3+ATiHa11rudMoyFTSloOqDGZ3ym8E4VgYF5jAd0C8buw7KxPzU1qhB0Qt
BFwKi7bMfs25aEQkvL9atPhLiv52NLB/J3Ak2Ie3dSn93OTM+T0hxWE9dpdp4UHe
QBqIqdpEGErs/76UvoGaLy+I8l5/KktX407UhTurzU0ZMCccFHpuO51WvUGGRyaw
IHDgi+ht7TbPRjTFHcSImXzhYZuie/0rF5x4ePMpLixHjzAvXj7xsLOhan39g6LX
LfPucLV6Q755hXhMVABqrlSGBhKNpAbW3d4k2x7xqx/Bw7y9i/1hnbH5knnyHJsq
FRrz/5GA18oUCP4r0+u57FKr670qq6FmbuRbaddHDQpYZjdFr7Z4esw8HQwb0g5n
wREncB71D9am449OB3U2SMMUWUMBvHC63krS/e0GD3rsuQpUzao41DWGCvTf7yxZ
7hNs6r3rXmVG3Krco9bAa+/kU/DgfgDGAJxbb0jppg47IhoSWj3r4kNDq61obfxY
jRoArF3vM4BeS7rkuPeMuUu9PlBu3qlO0xh6IYaF/pvyu28oJM40nqwxAUxdAGbA
vAh09IzvPLyzUu6IImsLLZeSA0otq8uxOLGTdgsGad3dyoj0uyGwX9C5v6K0UI5X
RYzO2XVqGs08G0t44Ow1e05/AYY68XW9lqpPHEpLLRAFZ7TJOf1FkCOiKfF7HK4d
89GXQx2m45kF6HpjFgM4+AmofHkUsj3UEgHogB2+HOJ6oKbC1vZkuvHP5q1Tsf1M
U0HfxYlGzjCFAKGHtoCFRALr1du2Q6aLFjhzk7BkK09iV1perrIYhtQoS11MWw2h
6DAZTbtWj9SC93P8S2BSZZIRRYQyFtEv3iroZytJlPVZN+5Ii67kVrS1ir4lpCwP
gBtwcRCW8e4jzllFanekKvsxxxcSTeljkHSLyzqiDwccnvUSV4i6REn0tMQqxEIB
w2FDntF3VHzF+q8chDVx9tl33ITD7P/Ngat6NOAFlDevn4Jv2ag1eI7EAcdEhSYi
/SJWT4tm+iWyZf8FmD9OsnAXXAVV82ci9Mh0MoISSZHdqrQDvlO/kV47rco2ZlYT
O580SpZpaVwPHpASanhFlVuqP6M9Ya4YtiUbTnMVtLtLtVEBrfFEpJKIMMYc8lgo
dAQ79tOH+4QdFUmt3F5zoAyysY39UAk4Jv9K/ecxtOPy5UJd0tBC7ALnHMRDHd5Y
xvF2i/xbAYuJquYSyqVRnXowJVTOmo4/D7prenMjqRu5glCIkvfJjlaTI1Kg3B8i
o6WFGdjh4OlNF47d+0JnOYkHcqdQduwUsQZbfzWdWtNRy41UpP2pO/2TORUzvilo
YwH6gWZJ06PpHNWKXQoig4XvP64Jt3L+8NW9nc739Zx0reUSAuLaSloHRpge2jfV
3MRiPlCBWO/6cVLCOwVDhPf16bFgdo/5lbo/WxGspZdSPL6J9gN6KAyYdC121OZR
IvvrsVfMHZTgp1abu5M0ONjISRA9wkEEaZoZF5mwwf+al4JFJ0k1oJO3I9fhEti4
2Q+1L9rsHCNX1kURunCrNYNRN5+z+1q6Ld94W8P4KeFOmuNM7pvdhDoe1lEZUtYq
20QXWq0R/9/wpxjV0pokCUI5KTse9KNir74Jtx8bRBgc7UYMlYn7j7PPj7uPRh1L
HDxUAQ4nk8pbknS4BYVCqHlKFrA6k3yGCtOpyNHNGJCTROxM8rtZy+kJVTyW9NlZ
WRfZhf3+ErhDD/87PZm/e8BWQKSdB+Iuot+tMXNq+MAFxPgF1lgxRdaT5bHwod16
gkFRVdPIWhKxN2eM34/Um14RCwpP0lbBNHU81LGJ9vzQCsvW8znm7uPVQLl113wh
vSeY1+bKNRHSokvCj54FoS0DVK5jS43Tr75GGR6g68J8L9ieKo2E7Z7f+mxnT7oO
LTQ6Q+n7DpZ3U42T+7qT4WMSg1rAP7SJz0lSwaBAzqMjcGaF4eB+SeNI70zwg9+T
52GCO9YS0Pwj5Dv7+j3opzrjcfbSKc5OXjhyyijLoqTzwjXsMBQZL8ZXlzl+F6pU
uqAB4Vnj5vR9F7KwW95aYdyGn78RybnHftDTMyb6JG7euvbkMzfCQP6X2Hb3zJoE
+659y3dyk+gO1vMcSyXuwmgEOvELPMwFZdy+i07235XHckfAUYWvS1jJrh9PJZ9p
e+2ZaStoRSL+Yb+rM14aYQIPxS142KRUXvd75wsrc/FRwvVF8gfPEtqWfX/jw1mh
A0XjFbCHWKFRYRkACfIRBx7ZsooOBdfzK2apgkIF0fhjWBCBJKwASOupCRNSFNmM
liz4hJDYNa+wDyLYMSJVqVRKOtZBopoYga9PlNGmIHl8RBMZNoaeFxICjUIumdkp
51nYDMSDYomDv1JZy3gGel0G8jwSws14nHUixIevgzMeuNFOsE3+oY3jqLuTXcGf
9kA/FAQaJAp5W7qKb+YP5h90+IKjeQWrdNI2D/HUUFht6nH6JjHnOhLvurLcZ5fT
jOc+hsYlUtnCwXcmSDQBF17QQP1K7lY8j9Hu325ZMaPzly+B8dTpikpd9Pksidji
x41Sx7EdnC5RzSL9OHITNFT3mfuyMWoMHNQW9zjFug7IwqUYQZkM9XLMFX/CBFLo
cdr9/pzEZFMsHD4aj+yBA1fQ3CakRwLhVVq/4oQNrCF3hJ/PyZs/zqwwo1e9YmBu
sISK0uJHfdTfChPFYJ3j3VBFyXZbWlOghAdR/UoZMKoz3YUpQ0q6P6FTJlh4XIKG
E+rNTVWzT66Xoy3X2jf3PiRT2c4mjt6ZoGWXKbe3S7Fl8krhcGwe9BcubleXBALa
AHjc84RDZ4CdNaC2ahNr+9QK3e+7sNnMcHwMxHUqYs2OhpJfo9fU3NaUyR/5jgJt
asLyiElmMj38vGvy69o9xsJpYv2Nic1tbw9PShvbL4LJOvjxeqhueZRdPvnHJj/G
K96DxT1wn73aCzn2CqQdmn6nhlXCwRoOT/dFQmiZXbbmzEtnjj6PWzSifokm+fQo
UNn5S3D28BA3I8Ci4r/jb87bOV1UAUw+akEKf67DtMKlLNu09C6hNUy0sXj60vjp
toA2UAGD8L/XyX9/M4SsztgULTCyHaUndGMNUkI1IsVHJVclVAE3cGkuds6j+r72
4A5L95x9Pb9bWcl2nlltqp8iLVDLhYNOtQVUOqXhTtR5FnSh2ukSgsT1FuJNOWbe
A7Y8ujUJHE3MOZJ6+GfK9tSfZ0mWYP2XMdhbId2z68rLAki7Wfl6YVJDdsqI8YhX
IsFQ3FjJijtxjMH6eVY78JlzyzlQXF4OXYJKJMyhZ4eVGMmuVXPSBNaFO6az3WHw
MKNKaqoGXz3HfH2J17uR6E2q5POcXefLDFS6tQYE7giUpATusOMWZHWnPOc08MUb
FoYMd1sX1DbA7F9SL1s/Ucpxk5/hRlBD2vag6jx1qhBISP1ydv3B1MEjCFX0QN2K
Cg/Y7smpCEWgFLCMof4xh1XGjiWSemTWzXY4mpavETMrhgAKnJ20TenFK6vxEeHS
oQCarN+ok/yBObbyMBiFEGSIEYf6o5iAQCX97NVjOadBF8iXKrjK3KQPKqeQCm7i
hrxoQopJa9J9ampE2F3R7VUZvjqPlqjMHB2uJVIw9CJW1Alvls2D36/ZOFD6K7Tr
qoN8MHeMD2+zw9Lc7QEyh2InhU9Ngg2UHeYYHEha+Qcwid+YFJhaJTq2COP6skJi
qkkDHqS77VciQ3eWl/QedroXuaj2GZEDQpZHTQTO1pCHgdkoam/rv5mXR3OSrccB
PxCK4Ukrx8x0KX+HktUl97z8AMaisCNCiuXQuM3VYT3z2tZP+SwD4W44Q1Vsksvg
fMw92OJ+8eDqkhbp292W1tfPiFJmn9Zhq+ts2z39L5wSQ9tB4NQGPbg9O9RCZbyM
q4BD+xxcm0JlgzkXOmMXPu+j7yObPMHmw+yHwFMJr1n6QnvXLf5y6IpMQWTAtSKN
TqIEiuAJgElcSldyqaM8yHqoKkavfM9SFCW8bNfna9R8iK8jRjzD/lj4OvIgVbBa
2T3daoC91SoC+2rCzwfvj3NdeUTQrPMW1PuJtZEjeEnOAkq/ORjeWuqs8mc1W/Ve
I+/QiX1yCPkYCEczZtrZX0YeTx5hd5yOW7eXPOKWqkxmfplitk/21iwejXD3Tj+9
oZHT772pde7WCZ/oWuO4p0L85bSLIiBmBmiCHLp5fkt+nDWHzObyjJvKAv0OktE9
iTWiqiWyo0Lg8REg8ScI0YiBkByC9T00H/IsyxSdR0+boCqqyv0PZxRSlnhaKwv6
wq3qebxYVyh6WwsCarHayaV8XvO2B9HyaEL0f1jl+EYxUBj3fzovUnqrl+NWlVUV
jwNt5JnhwI4AqnKFFcR8vK9w0Sc6k3yFvv1sFQ06awKsgchws9+zjh6JXuXSPFu6
mpyoxWrqN4qjKvAzLQD4Phc6YjaXfbmz8XNBQPN1xD5baTBdik2VHy958qS70qI0
jwWQtcAPNaP/I+rG/3t6UW/HSVITTTwI1hfvkbQ+PViD6CLK4w17KLXD5jXnbFZt
uxKTjBfaXbWJdFbRLFjQKH/SEsetLJzKM6lL6M9h1ryGmYaqlnIPqgIPS1MwYaso
lOkhhMDO+VdmeXE6HElwudNujzG1CTaNnhgXYtzu9fSvopEpVqLoGU4CtzPYtXP3
YBZy3Q29Eg9Tt3ACaQo3o56UtfGTkrFed1ElCTa+2IzmGoTUUFrAThBpe5dSGqqc
hauGmqdbGPEzclxrSvpGOpsad+IM9utemOSfbbT3c+WlggWvjfc6+S0wSCiPZrtT
TLrPZ5ymO4SqQ8paJMd8MMMo33ZQGHSGLJx4aezA3BWC78YxExrkwX4aHJ7zm3Yw
wNb9vfCm3I8JoQxyKTPqwxfpcihsQGHdDSr9lt4z+TNR2OaCLu9A7Byh/sBY0Vzy
mAwpFryBpKP+5UtIfjCaokGEjgdO42pcyMUA7+Yt9VIsm1SZjIB5ni9LBs7O3K4u
o/wvgr7BKkrUVe+N4Fj6dLFkT9NbkS5D51GuADLZe5tlvq948Wr5djAFmudXDCQF
Q4tUnoD3NN85AmtgPUGuOXlj7t8WAHPfHKLPef/+Rr0rIY4FCQ+Hp0V/dtZNDsUE
5KnI+gPMMii01twd/gt3MrPtZOruzkXcJKAOX26BkTJULn4gGkblLZd0xFijEm/c
6F2ztY/4vlDlaZ5nTTe6AFFP77CYte2VLDYwlpoPe5Y8CjQRNK46zEOAA/TetQpw
ZeM0oWe1Cazmdiw0IgKgAQUwZaGtRSngB1bea5Lhg9LEolqvqUYrNiqJt0mtazDq
AtQEAfruSxCzQ65r9FmFnJLhmaNNjGnbeaLPfMAa42oTO9HKHDGO0v3rjfdceltM
e3fJD7IJazy68F65ac4a10QW3xjppVsXjpnqzA3Xk+s/CMdEyz3MEMpFxurxD/LZ
Lgw7tLW3p7NZlLUPTFRLwuI0wLZJjusVoDjowikybF2PoHE5F6vvZM7cjcEI02OJ
8t4Ej/0VMt9Q778TZWoOtp41Jl/mONXpx5KdTjt3vexRzuLSLFWhLdEVtEKnUPl8
tzb01d25tym6nJPxcUH6o5VKqZ1SNSCndfRIKCEWuPhDaSvVIUCgP2FqPpXd3ZZs
puEtrlXm6uM2fYxcyYyoNJT7u+3Pg9wNT0c6ln9wqOUcE9jtLN3MlgXVxFQe/Ika
eqK/Adi80MB0mTK0qexzD2+tXXc7a0wz0ZTxvldTSboVroSZEZhPZxD1R2vHPJVc
eufQ2TRSyra2SS+elS05tP2pCjXF5MO6T0dcOqwvH067BBJ3vwgJRoAf2Xzqi/vx
fpAEqnIVbszyew6xnuULqGBuEHXJbuhueU+tWmoZqX0w6cUSqlW6M2RyZg9Rcx9s
k1P6BOjKsZFnni6DAFwYHHY7MdJlUSTVu0qOkpbL6crcyLRszNOEiiK/qrK/trZw
eU+DWLudRIOT1ayJgYkdmhkLf20p649yB6GlBA0M0q5QqgYBm7YkU8f3pCv3ewyr
soH1htYixUylUI2spmtq7Kyq6iwBSJdGvBBSTZdmRXMBoMynTwaKTy6NKaqzt1hp
VUXpj7Dch8PZe1ahiwwgIPxHRJtSwoeHCuaIEKlxe1a/U76mmefvxZOvGuEiroSl
zi2NUQCEVC2zphMKjMJ3XMManeY6KWCB+z/3VHiAVHWARZc/4CJ0IiEJWSms6Ny7
0D6Ab0vFtqRQEX6b/lXY34pK7dnaxgkKDvQ+1wPzTjk4+TEV375goyY0IMZTNyDn
sjbpcSwyluqzUZm3QESvd2jqarSFOcwTLqutYaG+PNuGpt/M99q/aiSb9wIb9Hmi
93HgZCfdFoBzmbHp5GRzC1wyCTMOFW9n7MZgeVFbouzIh4g+G0DkIFxGnaNFvjhb
mTx+tsS6hEd7RZcW4KVEJymcF55FDbnvuqMz1AYFksPb7UNCogSfUWKtbzqhQ0OZ
7pQfyamviMhWN3vAnXwBRmKcruhbsmu1jjYZaWReN7vvTiQYOlpGaJYusehr9Kbk
jivHYUvaBpjFIBbvi6ZYc5GwH4e9rImJH8wsO/5dgWcWhQzHHyTYjSdnIWEQsFAn
GGR77jAPrtmD1mknqXqxpwC1GXR9cDeNGluXnt3IC3a665Hb+pGKulZOHb+Bp3aU
HZNP20W8vjfxli/Rx6h5p1lKvGE/8p5FzZIHzygAJkzeiN9zXyUvmArySJzVC45f
J8BtEjuFRKxAaoTInjf4+ldHj/0AAXq/9DrcrVAKAcfTtlhzUMDspCycDNZEGhr6
CsVhJhnMAUNWTNQ3rYXGAEDRAZwz2RvAxgyDh7js8w0xbgkxxd6QR9doKVR605Jc
HkgIYET98MhMKateMSW5gt2Eu3m29Pe8ClrNA+Q7g/rfsW0HR2Yh88yWsxuQuS1x
l7eghjk37sorcJCPlL+Sxelb8leImEHUR0wV0HxBa4rbyH0FRoeBBFagRvL2ccj0
MMOERw11m0pFypxLzce2NwUQmBH4xsyjg8gtr8uDjw053kJf5wEfzCTOOxRQbfJt
mSpJJsZf9vIFhXruuBLMTn9Kdyp1IyhE1Fo/l5G4mokz8Os1WJ6YWs9X8YLVYrQt
0iDG+FaD2QsMvGEdai3B/LzXVAJHXcXZJxUdIl7SAFJjHvxyOMXoC/xj9etUDgf7
8la5D7BGmgFocc1vn57M8y6Mv4RJCjemS7TBHoVQS6JyIfa/yNcpP9CTgpNJLL33
DImz5D05iqTVeRWFtFw9hOxml5BN4Mklea9n8rV8P4JpwGH0PwoN++PeXAee5/1e
4uzSJI0/OT0hW0xdIyxs8XsHlA6n7gYvv2C2Re8efz4z3a8PtXNYpordh1D8VUK9
7eBghw5aS/ogH/T/KedK0MUIu/+v4Q2EVJCdE1RW1OvHdLsFCT4X7Z9/gw7/fbJw
thxn0ha1lrmqwxlLU8BV3AOsq7/dNrsNVtBo41PGYY9TRmM6s9ds+z0TbbrzlJ7B
6PWZGavRyYX0CF+dv9VVebPllKc+nLQUuh/FrxB8lNLMQkr8wSioKgDq/+FJIwyh
/5J12cbETxifq2FZrgvrJ7Aj1M1JxZXb+LLUPxZ+whQA0slsmmT1Kw5Fsc+UFr1w
BCy0zFAa+CrQ69K7NNjt+27C1QctMvV+r3N5nPnThnpKTrVcATwqbqc2hUNBcndy
0cy7Jpn6RAxrKHch0lM51lWTgvacilzD2IItKp8VhD2Jq7Fu5+MCMIVpaPEL6qfn
d4fpAV6KWYbpGDkxiUwFfy7/uwVyLLTMdf0Qpf9+QRS/11lEx4cQ7YK3Dm2i3Lge
p9MHzHpta0ZX0NycbPcplkWpSzI91DmGXK8pWxjUtB7NBOjE6q8PcloHDu/K1F/6
zAlT1D1DqqN2QSKs/9Cp0cDZbZ6UPKZcqiK1zYYT9/B228Tr5JUNzuzj4xharKeZ
L9LrHEh9ntezWQntlNMLseaLnX8WHJIqZLJd7GWDNyVDGXYE4b4c/9uu+aBVHI8B
y35X/S45AIoglt8YOj6B2XNtq31je5KX7YETOxdb0l91blhDIOw3Vm4pMWLr+KvM
4C9k/6K+jOJMV2JGLZnCIALQc1nEK5wwpr9oEDngrYNQ2hTezdvzNO7ZbIt4OQEA
2rR3qXNWehqVFvPKrbEv7fe0Mm9mchou2ENvU1n2oWTnZlfCtLc/4l9dzsOSsIBg
iEHCZAewBYYE5nKu4jVhNIR1QdBgGoRI/UsfYrIE31ipKluiA7Dy8+uPZXzBLfXK
AaYTA4D0yREC8kHZz0iu+/Aj2ShLttzAD3M+JpfGp1QmxCiSO/BGZRonie7LOa/m
TUeuEXyFIH2iXbYTTradvFZH7mb9EJ6+KfrDWHVLyzd22EOV7R53wtMWl8EDjBIZ
cUgvJYcRDRLnRgDvsqRBDfkR35Kpbw8oJcxINDj0YDLDu+62FCa5s4fJu8CN6f0z
rcDNTbNELOn9zAcxVnnj23mzz3KRyNqbwnOm6wY3p95gCKHjKauQEXzx21lOPSId
N3IEJqmyUu7VREiD2qKFnP4hTYWl8Kx7T8jbtSs42nCKnfgXnoXKoPgaxNZYNeXB
CKioGUqBD8Bz5ON90z8YjgG06oWSqulzKbL244Ena5sLCMPbWnOWsnaziTl+I80z
M8zZqGvn9wYO7Ve4LNR+BlBYXanEYpDFdTqv63dsP9emfff98D71YeozMUno1hlt
N9sEngmpgvGHpOPCjVwHvuChhBrdsTXtNJPbk0FmQF8UD8zfQn4nkP1RbFeWKPyh
90MED8Vb8ct6S+LcnTRRf3EVv49nv8aqExty35ZcNELokTSkOafnfdM8drzdTaMU
Q08U3X12RW7ze35Z5KUgR1RaqxQVfrMu5fR8dLYg9YsY5U32IaCJBu9O6qVo5PEJ
C9A/fQkiB4n17wxJJjanCGEiANKcCYvAw6c+TK1rELfZYs58cTo8Go3cP2DB/RY5
TAqQ2S1fqQEhldOZ7RF5MNIrMzO5ONhOHCkRS13TQLyfFoMxy3JRh7lKkPuXCWDc
SXBYu/ODcHcnVK1GeME6vV09a0tiUgTBTBDtPoBl4dSx+w8I/3fhRpao/49sMmAY
5tSjQSGQm2VNCf4GgAWmp38BrZzXSDm1Zv4LHO29UjotYSjl6GEx+4f47fg/XuTp
WoYpDaCtJUcYjje4vbBLwkFuBLRqSMsOSHY8KOQ8wr2WDO2nEKG7IYVFULcCGo1F
Dd1d8uaDiUMoNAPahiljFlj993/u92keputPL9kobT9NNXO8fM0SYfxigB2Lww2w
WsqRlVOEMXlAY8VDrg6ABskLkLWsMuAgzEVY5sJUqUPxdhc7LobqL4Nh0BY9B8fd
blooYrNzQfElsxpsWCVIVW8/yFxZ80ZdAyoyKJyRQZEcs+TB8EZMLJl3vfL0nHYZ
CvTiSroBxxrzFT3MVQY12594uWpZhjEM+vnMyM67nWNs9QIg690zj8o50mp8iNGD
l4LJflm8pwx5+fV46gQxqZC92Z/d91ZZHx4sdArnaoT9YhZWpY9o1mck+7gnNEdj
j35KGY34JPhpdGbDdl564Q/kMoIVqYNBX3hcWyiztXeqcrnt7mu9hCy6SQti5lkG
u2NBNOfzUAaiJuw36Lz2l4ep4ybm4sP8ZrYXQZ/046+lD7RLI4oCw6U13Uh8+XPV
08f40Bu4T6625P9A91VjbWl5iDC/wRiMclvirYAiadwuMKjGkgqlWs0KvuBwMS4x
/Bnjsw8hpdGuf375Y81Zl+vJjSQXAtpLxhZyU9qOocuKOjQ4VfYcyc7/EDAfdvai
4a7xdGhs/3Su2QkznSLrP3ii7yRa+Ya3V2VARbVYgtoIOg8cXcZZ9TLgVzjz1572
E3rf4jobnlUWTghsuoDsT4GKMiULTDJomxtzCsV12teqoKsQNlqRQLqb76tqevA1
fpxGMcaRvl7p+n9vzMurlyyXm0AKIgWgFcqdij6Uj011oE7gUhP/66BCKL/0mmMj
3kXnTyXhywvJcgIuOYwEcmdO/LSDAxuEPOil8yQDkejHVfmlafy94N0Tia3xL/Ly
pAg1fcn8yqoLAeco68nbFe0BZIbQ8ip+LaAMgBhKKNkhp5XLQaUM9mtuAPnty/sM
gke4zTB8CvpZwuoWI+Ut9bKm4RRvvhTKrmMAbbXv1NSNAyxNlnBFMpu1Z0MlcKU/
z8c5V5e37ocXAGx91VlqT2lNpPf/YwDTzGbAuuH5m6Cgd4GNlkpAxZHTBQjtfeFb
0da6pvM1JzR2Q8MkW9+JH8p2JzD0SF4XGFk2MsMI8l2epdWTiX7xTmNfQ8GpaWtj
iaAGYBL9znysYtQKpikz2mg1YglnFRPbGmKzn7mw784yRKMP6srbmVUAC+LsAwtO
fIhewjuXqrFwgXvgS80JU3rC412aHD/pcRYxLZ7ch/hoKjDnYSqFIdBLO1PXWXc9
JMvZz/wRZZZtEFR0bFHMcWN47S1joI1WrQMglzu2zid801+BOkLmyz+yxAk2Gv4S
oCJRQg/7MPd9iYhOyzBnR07Cp+Q8KE51kSiXeLR3x59xi9j2nwT+7YfaYRPHNhJw
fasUqqZXi4tzvB0tTKvw2wvdAXJUW6jsut7K2S0NB88WvMSM8plryNIPM8udipV7
fdu3CLLl4xlv3S4kqjtp28L+VCgCU/YobtH1xapsHzeQd5tzETGIJ7MDqZS37VI3
4TSDik5gfxt+aenxxskkbAbPcV+tTb3DRQBSryc8wdU/eCkr008DLotMWGmHlJbK
g+7IX/m7FvBfJhrOokDh+FlwCZLElSxilM4dUOI4B+9GsLOxaO5HYhScux0GWtLX
ddE2xW06uQyzIAv4YtBHvvz5MUqrtMj5uCvWEjKibW1bCsUAYgZprOUY/DBFETLF
tNl0DRMlEdvEGFupbFTYSXz6qlOxD3FMjqhxHnVdIwH2brNh0BI8v+/afykGR2R7
pO7jDcNdb7p1nKf2v5QSJNLA5tisYK0KIgihYf/SoyyBnnlaxHQRwtYUvNgc2wBj
Yf1v3LFc1iJ5wE/i2JTahngxCmyvV1Ih3XQXDljro1aP7HtCjBxkALM/dL/LpqcK
lAMqC7SfMnotkIa9yS8m2HldLdabzScdCTLMN2Nlauo71VCnknqTotGlkjqF5rk9
MT84JNvDz0WcPNH3GN7dlu9+IXOP2YSKCU0Z9g4L8Y5I30kiodjLial22K4dt3k5
6rJlskJ/RjimtPlNe6/Q3qo0KVV/Y9ZFyNbXuXIzvskPb7gFEFAPRy0pr3/kpOUk
I3xb6Q0Ts7nhJOO+AZWP0MJHnMDdQd9iywRvTiKGR4pCcAs/grqMrH0BLm/SoYPa
uPYd9vjP503l+jiNm83fF6qyx9a8tBqd8oMdHuTmKVfJs2C7rh7IWG/gwaYJ1hIC
GTJODI2wiVY1xs3loM4zDl+4dtkTBjyOYDAdBo+kcY9TcpVYkQoUF1MDaJPxBBj1
naxGB8rIQYgLRSRE8yzJD+HwLyZOmpoIEIcMSQcCqNG6VIyC02ObAqMDHqdQl7RD
N1wnXxQw5n6o3ys6NOem6ZinrqDLBMXJLzn+cfEFrjH7SmeanTXeAe/PLMjhHHvP
GgNJTDm1b/fuFARFQP4Pc4EUM+b00B76ZgBWVSbgBblYGeI6Bhrso9SY+KbchINP
geCIkXg+LK4v3uQlhIM8SNgy4yoekrqtTYoR9W6iYh6M+JJGM/Lwhdji8GEFVv8M
FqALkOa2HeWtFo7f58EG79E9mYJzxtZRknHhBjUONoX9/CLVkQCHLjKGvNW7EbKP
qGY+xCXEyq5le6dawveAQGCnVV5DP8NIQvB9vL0eYwsg1yp/P4KxTDTiLk7ePSUb
tY4DkCd+qxQZZBoyutwka19f+oliljkRY/ln5rt8+iiVpCQ2Jt/J4Z6RgNxV8knl
sjbk0GUBVZ/Io4PJh+iSsqzEXqT+//N7x0QqK7fKxjZc0Xj3eiKyuu3hoPrMYttX
5Bnh6+W9GbnwBQiWcxXekEGJgrn8nigyG1DYTHNAXur4OWD579UCSU2ablvafcY3
Gp5TJRLmvNg8FvrCSsSax342xPlf7A2IlGwtWHRg5yw3ydVBU2U3PNLcW0Pv3XgB
GxTm7QO/bQce0VOp0SSdQmr84MT7AP5MRQosKLFq+cCyDXFi4DgOwPSzgrEjUDM3
V7qwNByS1reVyHbnzVtXufGKbdmB0An+Tm1LjYuVyewFeXGZs9sYhGQgv3w3EJwG
7Uj++BL/wld/kv+o9olS8yPkI4dudNMvNocDTy+Qhy077mciMYNDRcDhbLA93ImF
q3IKwHMfvWvAbq0j5hnHNxCTKC94cx2YaQT+9mho0u1qs05e7bpwf64wdA34iEO6
dW8eRg2PrD3feUNln2qpKtttBeP/koux8qJbhTCDYkaKm64yYBS95yBwuX9U549n
PfOOCE93lvUbJi8LXFp4X2wYeCVD01ZHQiDpuScjDhUE7jvYipiQp3cEcDMmldkH
Fq+08UDqMdaUBMJwcHLH8I4c3A8VSvIqeG/zzboli4hWMAai2alg6bFNQgQMVzey
ECirHRjRhTE0FEE2UGTD9m+jcO+SGJWSU4GegR/7GWnIBOtl4FOJXBSCoB5aiva3
gwM5aQxmCRZM26lrPXCgtg3RJaVr4vf5s2QuUQED12bhwxtO+ATXPrV8RBWq6tST
GrK5E5ZvSJuDVw1w3EUStZsxTeVjH2ixsfZ+JPNBCuBzQLRFGlrcEItQwUuczxg3
vKWWDftDESOecKFgTUd5Nn68tmxvqP/uO1D14ImdEwewTl9X9xLHbuRZN5zBRI5B
4hQKXl2KvjwrZ2g4+oYiHOK/bb9Lo4K6cs9QgFcMDYtt/p2G9FpbHY3eP5bPutTx
SHz6nNO1DBkyi70EKWOGuY4aJnOI8HUPSTddfKNvdhu3l9IFjlWQ9b5KTNgu8Dyt
EC/4iuJkNLrpmKIMIIsFyh2kArbLPejizOKU9fkHGQ60r7Nby6yb4m2b5W7xrOLb
No8+CGTXNracs6RGdJJCR/pV4/lLB73VmKHlAjWpYoeEi0gH/q+tEUJDk1kSj2gG
RCGxsNYCpkTdCQPWmB6NZkPB6Cy/kYD02/wZHPhtOPU0yXPbSdxplfSMxU6rq2HL
50lxq1Y5ByvQDKUgicrs4Ceo66WRIu7sms+uzSfXsNTC+snAKthq78n1zJeqPOKo
ac9J9VZA583iRuILCswIPKJiDruvYGhvbdn5JMgU7xgeCjRMu1At8/vnBoMTq7Oq
6ChdLSpyAzfl0Ydmral/f+st/+va3p2oMIC7kYJKhYi7t2Css2fwxFB0RVYPchi3
f4xzMuA63thZoVpbGooyd2IKCbta9NfUMhTXh2r53HF/JHhJPy4uaDFxlFd0FqkL
lOfNx+E0/8qH3TpC1fFKlO3a2C744sjg+UArdtCeer/eAV30B+vRQ5QDMh1sDG49
6RJswD3WwShu02z9q3MDnA2e1EMe8v5T5WIL+zapv9m1qWy6moFsiHhQJTAEyC0B
gPJyVUcNPnhQlDA/+XKE1Kv2qDpgiiKWmKYcTEmQNsevaCzO6NKBw3QaMraHMfE7
OroQAHFlgapuGM9RpxZymJp94XEMMMMgmvTP23o4Kyty2Ot6dWvOW5pStfE1jRyM
0Yv2cSoACEBWEIXmaNDvqgmVifEZCJpcD4CuZH19dFer0d4m3FA00p+xsas7WC1d
5TlUlZpXw9qVbNuan61FIftPidZpZMN3xgSP4JnDHonEtVbKxzK7/uEKOSmJ2yij
RiWPFxI9L5QQxhCynqxsCRWxSqva2tv7t5XQLNRbeZGaqdEcelxejN4KevAFFQ/o
NoYd6kXd+3azL32CGiMadNEKd5XY/9FLvmO6yjG3wOh6u2cQ0mbp10fu4Loh//E4
cC54vb81eyRADOkpNY3K0VaPc7AS5iHkjWn8JZsMOcTmXgHXJvirkex0QzlW4/VF
BA1qj7QKywaoiNOM3yv2SxcLrNGD3htUSTR/b+ywUGZLlmUxnFIWatxCayvLXuhT
RPoDWuWCiQ6FPiOfvtErqOhbJOD2rCnMMk8B2enCi4G6qChZoY7o0CvuWV2xBqCV
vQu+UaQk1+Y1yGamTkNPNNlo1Fq20vz0TwJuIFJrLEyHdhAhe16Z1TOcHwKRJPwu
Vj9B4n+qOBS6EtzpD3rZ7XT/LjIzGyCgSaQNBplMPtTey85XJL9Co3lxnXgQezT2
RHgIo5S9Jq3nv3wBAHcFLOnolR3qVLe0I20vp4+1VNJR2wpaiML+yJKkEHzwA3lW
sZkwJGcZv1yvW9Imz1Jj5uiwqgDp8LQrojoQN7awxOE2wmE1GsUqzUw7/Gxf9AJR
AvlH9tKNwyC7z26h+/D+1Dxd3WYlMQE7sA8WTlmH6LakrRu5SEnvFKjlL89pJxMh
hSFOpLGGYgFOT0xKg0n1/FiiyWoT4GzrpGyDsmDUzY+5k9UClzjWoyzc7c1SWYTk
xH8Cwbu4IkSQiyjt+8A+nSoxZCa73HZbxYoe8QxdU4U3UcfOAqEzxDONyK5WvgpS
Rw4tydsUtbErn1z/E4+1Rc0jk9x4PeMmTabN0b6pZost+KeRuTvvvLZUJYwOQT4x
Fee0IAG5dXgdBrH+xfSZcDMVzrf4/ptHSNeS9xTdfTXiSdCc0L0JzKNIEcm0gwBJ
QRuGYIeQT8EnIMyWIusZwvJD/0+T1vzTYvevrT8yJ3vrL2yIq3kkKB4zgJhnViEl
snZpsHl19BZQGlzXxszWVYMLxjqDU++8zT3wzODkqsce1rhzLxkgwFI3B5gspiFQ
jfLsOPuQV2rGDlFQvyTyP2snIG5nmGUZ5PsTLJDnIKzxl/+NWlyNK5k4w1I/O5so
bakFW6YG37VDjaa6azg6v/9aSF24VCOKzBUDY7/e9dwKfg/0iDjC/Zotcui2IVVZ
/ucNHoE77Mb2fckg7mB/IkeqesR+xiR34jrRkC7RWkcRbSDoo5zUMBgzqs1vFS60
iiZfefteeysA5/k2dQLCvXPGWAhcLdLrv0e1bayT+hOm649RGJ91lWXMhdagcUVg
dczz+tiAnDII5spLHmD/5ZN53XN9zOjhaFPUlWHQhKgpX65YiF+usWcwohSOqli4
81msIIY6VU/F8Ux1HzSaKxfnsbFznKr9HRbfsD2rF88jxOi8Rt23YkhYrUTORTf4
akMjODJc0hKNuOKYeUxJr5o8XlK5Rsygh5QzNIUMSVQsUqfKZ9Q4I//niDhRvCMJ
4YmAPMAeyW55Dihb/M5m0T6MW9ZeVxCtbqw01yKwx4IbL4NXTaetsa6w2c8aRB9c
Lrj4818GyjDRIGP1BhUAlQDBBWEyLaQ92dj0b65rOtNgMjFvgbKoBPKtPJ7muF0t
5d5mbmfaNQtVCfiLEvEXVRsaEjJB1iOka+zGapjqS/xCaDcoy45rDf37tKrc4gat
SRncItWmptzwq+VsTB2J56FiZcgo7Xz3W1dQfa6flxqqvz8OJnnFfNBbB5UwvOVr
69rtd7uab5PqrrQm+nJ+734jrYGW1XcVGPyPDdZbugYhj31PxyQRGE0C9Aq9vq+P
xWboCBvwLxyUr5oFamEBuDIMUe7mPhl0jKcpcMwfAsaAT9BpSartYIf8/RdCFD69
8jXGfS+GWJdCGhfF+0ooFAV2dMGjFXDBxdOBgMtEsJCPdH06ERafH/F5dIF/7gOb
hXXoa7ihk9F+otnUbtpUNZzdoTQjOtaObUkDCfArETgpvHB8I6GIzZWporvlsue0
f5X8/iIYqKzhrNQWEm1eHm6WJdFaGSIDhON2BwN1k4VA30ujiMJ9cHtY85Ha+GzA
xb0jeHvrtNeMbARyFCpavZAT8+9TvngMmi9k110CR0LVdJLT4aGOXimi0U64/TUy
XScnpZoRX8ljlBbVwR44y0eQopLlqA0Ye1e4DCG0rgQ1dHdC0UXDdCMpgkUvdCtH
7qZ3U3X5Dhw/KW8mDGXFxVSPaDOI2wWvmUsp8i/HQpzD9pY092XBmbuvmw2ErEjR
0ctDJCtbWfqg1DfXVjU1+pjqKr62MXqE+WKK/aEwM1fUJYC4ntQK5SnW1Zvb4501
dVX8I/JxC7rT9Wk11XNFGcT2sEHiE1+rvT8SGNeEeQJOO2lx9Sb4s3ohNXLYyeTT
BfZV5z23fXVaAeYfRtu04ZicVRiPDUTbari9yip6qVDlci9bFkt7XoD9C1uIi6/d
t753WI8L6xBhVb9F46MDV7f9Ns9O6PZdBBvgHY+jKMtvg8yta7o+WfqA5DCUoN4Q
HxTQb68WCIrjlNz9pO7XHpVTqHhf6lD9G/nv0UtWmNeacOywzA7H0anUktX6ACAY
xdM4L0DmdWNidqKR1rb/WlTDadBBEV2u1D8giupg4Z9hXdMeXEBY3NiCwxCCQCW4
J2WMiI6wA16K7OMRDe0I5D59TuFLsPneyqNRJD+NuYfcEvsN/7TPTeq87AGPTl1q
/qH20tZYqN/UAyILdiG85yYtvnEKTD4Ce6F332VZFMMMyxKWftpyEWvpaClkCo8e
ySTtHmSBllXiU0VYLxzI5qcVyI+5BVHmcWWjmtCGcUtjIISanSnZyigIzrfEcRna
FUTifzG6yVR9xvPKe5Cilk463lKfQZ4+qEWoCl7lbI2KFpZqIUVIg5GoHkDGIFpN
xfT68hyaN5Ihe6sJfAsUR0Sm4GW+668ouEOmsR2+sa6EET2kRDlHsg2hP8P/tlJt
ezeZSsgQmRQq2Pr1cHlt8vr2cR4Auxps+mkOHzzQ54nseTJBuBH+NRW7vSp6z0mq
hWzYgTBwn7xUqsxi7lTiRv0JEXJprGKCGJlvnYcQ6yfws246dYOi5Rqu1HBiQ6nz
YlDFScNbrGMQpzT8PNV4ZSRHEpLyQvbHk7dX8YT7WLvX3kvp89QOg5rnZ6QUlRBw
ZpkYhuQx41Vb2Wl9P0ahw9ChkqKKZANEOcoHRdIXFqXOF7U1AfL7+2PLLiOLL0fs
hb1k0WFZ+PmiacAJg3JoMB2nheutfp1VXdMtnFYaesfBcZWxa4eMXge0n2qUZkJZ
sWSuAUMOQTOdLY4ZJZDjDHf5AZ1HhI9epXapTnH05msV/4pDm3oiXnCAGE2QwtUG
gV0blrUF5qViTFJswDp/lQFcS1xAuQ+DktPwyVwN41+wjLWGQz+UT202/wxLXM8H
klpm+U82CFs8qvw5OTxRm/mJ8EwhT++0seLJ/kYk/rVUQcYXx7LkzFpchynRsU1r
Pyuk7ApVk3iopavMi5IAJE9XKjnkvPjmldN+gORJesJEkQKuXl1l8NDJIWaY81eo
9Eo18N9kyroGGZ5ehjXqBv+ufo+a4949MgGWVPEXVmtDQzoSoA7b/FmL3NOqDZiI
5VTKGbGPnqg+WtSP58upOdPxYrd4s4I9gV2N2XpaZekBspi2IDWnxUx2xPSPfwPW
MeDg0IJevLs08arQz7Hb7ueCdtFrEW/g9rMq7TB2DV3JQsWXTEWDpQQajlafB/Y0
fmhmw4oJMLv0brW4mGzYvAHLwm0yAYEQ4uP11TOSozHUXrk+VMSE3MKmjykZkjpc
9LkDc+MFDK7QfJMpmOvigkZlfFAzAj8RpRCwBcAiAXhbyfvDngbMzKS9cqtWUrv1
ost8HLpvXybF+xKyaUx4m+FLOXElES3WTfs6xbRbHl1NqrUAPezGF5HfjCvrM/2+
O28Y4SkNYsVn2qgD+mSbqYC/idDD1+j+Od2bny6TW5CZ0eN89CLxx5nUl4idY0uG
s8E5juOiEsqhkQdqAwOn7byM/t5yaUMOuvexyYDFP2p2J2PONh4oy+Uu4FBbMXVl
IxlFgrjRKA4hQT4j6kUCu4V2fpmQVprtGWMcSqF9t5rXTj/0sAz8gxFQkR8ZUFnm
GlvrfBSEsn9kn7A1Y7E+OoJmgkApY43NqRNBoh2g9bH1iTQP8BAa49R94Be6G5NF
7Xgzla/ePA/SU8KX9DiedHnIrmyhoYoV5O7DyihYG/SeYD9vTmR9AJE6qjQKN+js
ZM9S8SRqV0GvClk5nXv1baW7ZJY+1mzG2XjAxQL4mLaFw/JYf0pG45E2uO9AF2H/
ZbJ9OCzxhMCZuthriEjIWRjBuMHJkJvbltz1VTH2uTj3MHgaCTZPOmN9m4MHDCJ9
yDT8Ak0dIgVP+kUK5QGLVZF6+48Qp3SJm1JRuGYq+GEOk4HTh9WGPG1q1HDyxsJ+
zHxS4OQkj7hTFxTCsIY0ACbkfFQBBx5s6jvNcJGJqjAWg7HLQlBzeIfNJtOTOwCU
tT7L4vP0BCu9ZFOQS2l9ZY8Y7xMYOAGGPXSRz4Dd2+7fg0BQLWYgBWX9ktT2Wb4b
SwOZXaf4ECdVQA6uAVTm5bE5adag748VeQrFZIdyp9r2NNomfX47rHZoLudk/BQl
u7L28w1U4WGJppyN0NGIEe/1MSn5QIg2GpXUsgXJbvQJoGDSHkJb7A44oEIoJ7yw
vOgHgGGrSxK9yAboyiJsSOFqDtFO1qTtXhsFYYcQlXjps4ygM1TBh5lhtVGJkE0e
V7CsYs/nhm3MRkv7+0oVxQ2LpVD5Eh5/1xGFqQNFSBSjOgAC/sA51F6OS24KrX+e
NQAjRxfkgdBEQEgulDQfT2jDjR2edl/x+5qjrFkhR3OlNbAj903FLafoyp0YNkhR
VecmA2boqSQoZYxns6A2/mtd5CVIv6S7aPyuF939NHGsRgjpEvmq3FpcuwNB3xeW
Cf0EmrviPt9LQW0CVYqLc3i2OJma7B6DUcb26oT4zUCOF/wtPjEW7nND8d6jT6Mk
P4xF4pp7/uUcoTSjSkMiI44t1Oi95A1/46PYztub7iLoJwt1B0Rb0HXFXwdNe/OF
NH9u0ln8MNCh+s9+1XqJ+NP0Gt0MCrcbkmt6g4zVhLWP86IjqSrkdQQKcp7bqXo4
LQVBT7NwmW+T6RB+NLRcnqNjt3y1oHSnWEsvvwPr9n9eUvHP9s5jhEi74Hl4Ldr0
GGMiL0yc811+ZdXban3qn5p7h9zQPUY28IJLYkqCD0+7QolzTl5RtOYbrEhnBxoN
QRhLowB9W5dQs4cZOOrzHOotZeYNZKAeLw8sMpENtPm2t/lhKySxDZaqcQwffDk8
mwgf8WgxD3v/NJxz5hg+91IsthlKwVDfK9G274/0ATCPW7+9OHoXXbwq89pWt63F
AkadR4l+zV44m/4OtH8T4aSHxIzhqyKZ+uoUhwaoVd9pa6RYUDCijg1OZ1jNY8Fl
3mvSOpictht+hLPkCHv/10fha5VVfspUPPFJKIRKQAs0Q3QMkiBI5rACzT5uzBem
/XKeq4v3B4qCAQvoKdPviNdHSKCZB2akd1AaOmsKu64h4zghxe47AK3ggzq2TpDq
o6jhC2M4LMxfPaBUVoCHB8vb8B99kHk9wGnTDqLJ72KhSCPK78cE2Iyt8Sz7Iuzr
XgLDB3Wgx9Ikpuf0OjG6lf5bwAwY5e8mbzOBMz0JKZg3VDMBc88NdNBrplDrJBrL
Z2Jt49O8nOnOgdJ/z5177Nh/tJ0NyqjtU9C/CCEqeKGLO0XcInoGN19jOu4iXy55
GKYMmtF4RkgPMQ8dYTwn9IG2opdAfWoSLvTcKlJ0b1mTxe7Ll9vNF9AUKfxAcwSg
vZrzRwjZOaDNtEn8iIOHsnvJktMeMXjx7JcAxBH49oonzvoh7rjYUzJBQavz4Up6
KLWyaDgtUj0BS7Fo/RZVflDcirNT+CxJx8y5iEpyQP43yJJuaZytpjmLqATX4xqy
VAcnHO0WSfx4JMbZiPN7UOfMka35rzfiOrxtLzrv8axNHo7jFPtiIY5t+vzxohdY
OFXSrw4vkDWtGf5AMt6kOOMFil5BoCiC+ND9xZcLVAIQ9/odc9Hus0Bn0pqKqM+p
co51cRKSTPQW1g2VBCmESgjZq1hurjSb3Fcl+b8dPzW+UrIudiu2DHPjY7z0vUW4
6R3PlOSu31E7hklkmSIYW4y3a7OBm9SXf3vXJzx8Dro3x+G5l0y9h5jantkkfljB
gaN25JpcCtPWtyh6bMCSmuVyonGgykuzvpOxIr05MTZmHd4Lkb7NtJQX9iFRSR/F
X7ovdyrmFDF8jnBfhbAfRCkNdTaDzx60St/LXUVHlt8LRIxbXrHuXigKD6o+XSpM
womsR8HxMnTQcNAP9MnbeLYZz6Qt9obG03JZgule////n/hmqZ6eD7UoCTKbyX1a
VmzsDbVte/W0/eOPOWySvXpIvnc+GpXWJhfNUb6fyJtAIAq6p1N5lWOiBgUk/Fnn
WX/y84DymciIxQvffV9mefugpg4SFjnkyZtgUozUOyKKymQnIK516VIcL3Qmr8y8
U8Zt82Kok40JTajSU/I7KSr0T2NN8QV3nG1wGki21DNVacHzZECY+CAI7CFFf/3t
bWjCgZ4F2niIHfYymOdMRv7WgAKb8lL62wgDsl4urKoHx2y7EUXYAOb43SzwqpA1
jjQQlZ0XY8MaIfXO5FwHIfTp7D4IIkhr4Zo0lnWjNeTf6Wohiuv6q4lavNH4v6Cn
0mBeHWTii1dXZEXOh0NTMMTnaSVxgGU5/nKxbntbWEdIo+mbxUaTKDRE5mEai4tl
3/ScbJs5ObBCz3ywscLYblxBJ7fVv6EliB6f7v0xRjcoGmHRyLw9vUBODifhY+M8
vg0z3Fo6RX2RsjMB9S84ZgMco2j+1u2H0krEXpl8tcjvASeX0Jb+2kS/Xh72YZzi
9IuB2VgBx98hIiZCgFWdOiaHiZsLbwbL1ifaqd22XECu/7QlvOfJFQ0YutAsBP7R
aDZOF/fK6XLbX1k4IHitQUtadIgw8WenTW9GtgpiNX3qQAl+Z3OVT/lAlNynid/D
YCJPunlwU2PeN36fdfQabznJMuiniS00Slke/DhuiXAMCpwZl03mIyjM2Rvho7/5
s/WxStN+e81NVEkOVytdmQnE7GmBTOD/XQ/0VPCcT0IKEna9H5+hhrfVEj+sNhSK
qaKB2tOQSTX4+RkBl2NmiIqcuhDmBup9YXa7dZw/SeIhaEZkFbfS2061iVJHrSwT
GEkcJzFKvKPGsx4zxl/Mj9nAeA6RFfY9q2ErDTGO1jrmqzEFqNCcqBvNTB9G30pJ
CahNFBlUzVmxjDq9GG78h0hSqOrboMqTohE2pM3D1//Es2EPQYLzHeUanosNzD1v
gZtPz4il5d2Te+Aqv6dhaoDO1Swpcbem/dj5K2ySJm4chF9gUAWlAMHU/NJcKZGH
i/5EpyFrXqfCBW3ATQiFB8FfhBEki0d2GwnKQ81lFPSFSRxpwlnrrBk4wAtLrMyd
uOoOZ5dvW0NIgVjhhOTY0Pc9wcQgohEZP1BuOimVVeyHCqrYUHmy8Qu9XRdVzwUo
nPBU4xwKfij9f+lGfoJF980o0srDycQ9SXabmAHK/weaIaJ2R1r0u8deBFnDb4Qa
10Va6yP+0P41kzTXQvqRpDOB/RskV7nySiBpvDeCvK8d5Pj9QWMYPTCgSoj+xKql
86uJDcUAPT4/cNXxw1vupJGg1nRj1FLHoFstO91xnx7V4nfbmJqWZGcrL2KHUz/A
kjOaitrVbu5jb/kZwdi43WO0dLh2V0vJisLnbYLpSt2a/gxRnsNfxw5AEJ+/XT9t
Hz9Wmu5g3aV+BPERLHEOTobwM2ftA0H7pNKadDCWplMkQ5nmCt2DdH4ltiK2Lmm4
sib0lSzRaEBRDZORBwMAsihIZwqnvAgLIAWYnZ5ZKqcyrdjhQUGEgAUefnEcK1Lm
1+7mWmeXrRQkLd1XAm0/t4XNmAOhIeU5Y4xXBuJKmnAFpBiUStbQaW6pZiLk56p/
HwbigY7KSHx64zXIXJfa7yOgktUWg+cYCuVOIwF0x4SviLNY36dnnESycX21w7N8
NhblI0rjEiukoSfeF84XQXEy4wpAROvdz+dpCLGgPzIzGR+arYEj3p7CjFNJPiWZ
Ib/M2qoUh1Re1Soav+CrOFfOWXwescSxDcu7rIVRX79veDhLew5U6UlyL/P2Dg8n
8WX9WX7oXBwh8FAbBKS90Q8qjXwLdseoTV/Oyqr1fdwpgKQCa0/VblFApArJJcaW
L5EnfMvTTjiiutxvWxqZthYhnchrzc9okKinevDIowuQWimKRL4mYHT1W7I0ihuY
Dyi24JQcF2mCnx9BFeJAAHOJj66SstZZZyih5LyTUETxuIjh3tFJcRVrVzwMhDYq
XpSC6IT4UbnFBteRkUKzLgS6Ns0Pb217seDXfTbvIWy4IWX3HMatwigCZR1JIstS
joFJSyZRlMH5R8jVHgxpKTRv+dIgegRmAOEKCIgB0uaPbvg+HE78YqwXtzPBYqx8
g+cebK7rwTbOrbk8jmQctuIoLw5Ae7rMvec1f/Wufc++b5xXdwRKNP9LnRrXgt0z
aNOSZYZofeNBieopNnLL9a6l/K1l+kLYVBOuG1D6hC0J012ax+BrKHqFoDtcnDzd
XCi4AHoWnNSxqpLDFSA0SOm43VMEZMfMvqtmmoqvHsMHMvOskROiIFx4rsxXTJq4
KXr9mn0oBLjI7l8w5Ehwgt6Hd7l9Sxy2XMt4PyFEoGMD5Rxb8UJWEy2JiMPFXAUW
QwHZr0MvkzNBwztQEe5NN3s5wBJhSQalsz+HKmzdQc5MHX5EJPrNam0Nb7LQenae
ZJ2HwZea0vHBwqFOWLlGrGaGUoynI1PCPy1/bAK6R72YWJN8w3yi3J6S/JrDxlQv
eb+2Dk/6c+M3yJS5kHzO4ZPaynU56Ygc8L6JXlVMAXZ3BQWlPezo2lZlSknPzpFN
GHqwk+r36/ck/P0jIwRtPIec+iYrdJ5aHWWAXaFOmKV1Sn1qkOhwDP+WBSUQc0X2
cX2+crprOUiUPVtfmI3mLnVss0DnSRIPe68riW/0cm9KNcWo6O2Dngy+ruul2FcY
yn3XcOX9gPZOclwhQ/mMS7chSumJdmed2RzQisJeejg2dmE7tas4urOIqHMebT0X
SvHN5/eC8My/vj6bSfYrNYSut4BNYVLWXCdPQ1dHPsRYdw68ujfS0fH7I6nrZ6aQ
yDkuWScgJT6kTx3oVDpeVl6CcJN5xS90k8ABTKF3IVwbaJXVdkWGhnO9dtC/yX0A
7dzwj2CMf2fwkLYkb60GdRCQNizP+ueLn7YymEf1XSC1LJC35mDhaUHQ2SfzOvJ6
+prm69RKAXYLAL7RJ6yC+nvtrMorFphm4CY4usmJ+rSfBRjjmbEy33NOhHnVq49P
JfrodOTZjWywqxNR9cDhL1dE0MW/ZV4IHqhQxtBHEhSkcnaZukEqSY5ZsLT0xLsE
FlT8x0JGN1XohKlFavlFdb7xlP6m/ke6SLknBFp8S12uli+TU8IipRH1gctccv/B
q34Xce4MfEuyKnQYXOcxlecWXuIB4vzu7mHTblKiiJ5HJQ4ncUYRnK+5v3GRcseZ
sgFVLjL6iufn8te5xrCZJQl2Xn4HiqowVKwFszX6ZS1323QUzXXU0LqPid8dxfqv
/NeQcS9znn0opPyGKZR5PRgz/s8CkyYLzNiVJnyMFiS2xPlebQ9PbaFIgW93FP/p
RnUJBg2hoRYJYaJjzpcmQmuo3Bdaa99ygNUf099ZJvzyj/+i699EuHEuKI19Hv/W
8DM5B4pV9WaXhJLw6xmp23ddINpCFTcquKFR/9XHmcU2AAkCd55T3AhFSOL0CHA6
GAN/1D6jgNzxt0dRfV6o8rLYGD1Enf/aOyHZxXie69AJ/WM+89L7nAQypRDAEVIN
CbqdReyyw9TZGFOBO2nr8Uht45QtTrM3PmCG2+tJ5lGNmPy711gxUt3WvLg7t76E
rQaANZI81P2Z/rcQL7fIRSryEZp05sN6+PWSin/7mMFIShrmZl1JdBjejjaRFxcx
t5XS67zoCx6sGBZmnFRf3G1Inp+fSzEH1CrjDgCWLg5eq/8K+QovDYcHTZqTJ3kJ
JOQOWSG+egXAa4STGQUae+58eODYhiUDt9ZUxvlFx8aGin6Et0VnlC9exCpAtF5b
gaX+xBTqSlhA2zkJ13yd1OoqXkCuRABTdJQG11U7hJEryEyEFW6R6zm1VbOPQX1N
jeVS3ebalenTwccUgQOsIUfL3ErOPcl0XG/epcKwM4DDfpBV3OeRWhwIURBVsArB
nVdVp6VGAGdktq/TZ8XD+BdDA/owfLNFHHznAPgZj6AEMqQc3LsUt1jAlbVWOlfF
UDY1qPpptPN6A0vCnYI3WXGOHE725k2lQfNNQpC/OOhy2jj1ikkA+D6DLnd87CLw
/fnlQYp+f1fAZGx1XZjgVHTCcuDXgJ17Or764s2zG6mh4Cxwr35WSx3iAL+W7oEv
5zHAJw9CbpOAUtj8EVN9oU+fb8pm2WdDiMhFcg+23GBi186negXOtF4NL2n0VUge
LdJKiQ6L3if2J1agXrhOwqcraufr9jJqXdg5T0MmYjw6zw78lQ/8Fq0xchi+u04o
K2Ss57xgWDA4zXYegM9t9PkOE3MwK7JSGESrLaAVQo1Xgjp/rhuaMtfNLaiZd1uh
EGn3IP5xzzgscBNieI3eUBY/p/Iz7yp3KKw6dWwRCftJydHNLePdP8cCzcFs4EX8
CCOOvaBYVE63mTQn8nUa6yEWnzSVoE6gzv0R2qNjpGAOv6S1Zp1Gb8IIF9STmVj1
vyKWmSecHqqzpqg/6FPaaeYEZmSfwJstN8EyMuo4YmeNxPVRBThWt8oboL3Xn2By
PNh4N/5eQMyYYAF+SYczlsm1mx+lUak94kLmxe1n58bSEvAqQ1kUnNCt8lXopV53
xv4n5oTB68ch0MD7uaRN8LLxl4fnk6kE5mmteKF/yoTBLJ/BL+s2ROgY1R9eBzBR
cCE5xzrlXjCmc8BOdKs0p7b3QhtU6U0PK0quKEaM4YCCjtkXm0Fy0e7iph4k1YS7
v98rs4qt+B9p9fOaZVuA8lK359/mHA44NTSNe7V/MxxR/mIxewTyfWcflxNLPiVy
d2kfgv691UBv3aRmbD0zQmQlYH94NAgtpcXmHPHbdfkMSeh3tlJ6jXoEP678NrMI
b83P/I1aBwnCEfJT/73l/1PXiWzPCtb2WElmgxGGILWJ2t+msCyyKSPqtdOWTwgA
D/Olz9AKKLc0Oh3GYX8hhqzt6Mu/pD7XgSB9QHg98HuVo5PviWG7kF3gF1fq2Gxr
ixA2u9bqrhMufhdpjzpkQyTJ5UscPuVgV795CxWlCVvX/G8HaJl+5MmJJ7WcCC57
13iK6Ld3reWEuQAXMbsfaoZJ81FoWHHAwMPzxaj+GBALUsSqXhVXgVctrK4D05ky
lT7MSbUeH43ro89VD8ndOGK3G6H6quvJrdseDTjbU7nPArYWMmVsZ5IaN/aepBC3
PydCpp4ihKIaiwM/iobt3PCCQBV/ND+NV2bwoHE5dtUkfvnalIFJ3pMT180SUXAF
qgcPhOq+rKzqfzhyoztvA8NHFjdU406j3hgflbAWuO2Ugr3SRcN68tI5EmqTeAYO
pMjATfPDm+6/A7d959ZDl+WeukY0N7ZMy/6gCPBInne5Iz0jccbP3GS+qtwS+2uZ
AMUtzY9SFzYuh0wnSnQ2J9Wg8zx6/eE4asKdo2uzd7CAFGx3KrCZyV2O+qHQyArG
X/SfKYuu9R6hBOqIj7M+12H0jwNk6gixZRJg804CYApJIfBwpt9eARMAEfYAFjb7
UyYvtxjiBT5SNjEAtd0yzO/82HxPx3uIvX2+Xafa4tQO3uUN4qUNtk0GWvDAMTX5
BtV5KATwNFv06VuRVVstvl0FmoVBUlSHbTSJVGtpVS+A7J8PBtKk/gLlxhRWQivE
drjTKUxo8xXBRDWljpedOVw4pQtHefYH/RCUx2uh8ST/kVdtnEA+GKWhbjPNsN9C
f3PSbiJdpVjJalO+zswG+2FJNAf6On302xCCmLN9Nm5nQd2a8S2++TJhV1kHEsjL
ThaG02pfOY3IUinW/gkY3ELpXz+EWgjG7l9GdWN2STHKU1mzeBoKJu0omYGt1rrU
dVbOihafGAbbCY8AVHxHBEja+s1EC1SlhUhAzjkVGpuzUVgYsYnyuWCVikw8Hh33
pUEoq/h+95aCi4840wdLeZ1H1DTImAAqklgjJKATU6Psq5P5N0RTMG89ttkbnjBO
IPFrbo2VynOX/MD0Qj3beHbvbq/NL8kiUngiDB+0c2Sc108/ZrBmOVCHzvrkipBB
r3qBTjKp9vLhHXCn0CjhPfPcRY6YBzUa9+k4/hfgZnEuoNQhaufg1osMZa53xIIT
0k3TxUYWql8/MaLkOIrXNI7Blyco5gkvoXVaNQYL9kRB2SFRWQSKid9TeFJ/G03c
rFDROGdD2VTDMk0mesEMKM67qpR9U3ePSQmWTQvlgOtYPEXSrRa2wGEc1NSz5YGJ
x6bYMX3pRQZdPuZ7F1EXElSS7gCCq/WEglEUYKp7voLT5Es2NBsHV1BAGNd7ndkd
tv3mneAlJTMMRmnuoij9opwCxhqAdWsx8VHfn1F+ozLJjATkTvLm/gkFUl7TwukA
ZooUnCYBj0CgukLtLTeW7oc0apguCGT/2tg8nYYGBUfN1Vvzx4HOgAz/+3iEfpUX
RGYTR0dKqtTiRxT4uxvudYzSfcw3LWb9u4qD90ntXLe+0+tAXqGvMpLa0FrtPUUQ
z41/0znZQ9N823Gi+DFfqRzel4V+iMKPG218x7NqryDB91vb1mR8FlCJ+fZpSk66
kKxO45+B9wMsfrHcXiDdAmWdWeRo8Lz+SpzVnaliaYrPkRQW+tocbbrG8sVcra3a
+PmDZSU5yLYChrnVpNVyqwdCcJ3dCqD8xjNZ4QH4Bn0Cxdkq8lJ/odNOdq6GiXzS
GF7Crseo1Fb71jxr52keAd56qNQwAYEByFd9DVPxSoD69YU6lp92sNMC8SzDt6nd
YmJYcTtvBvJV2j9GJAPtnhHD0OwOdCmVUS9/0N4ZS1G3i5l2yi0Havnh2+/ELGQB
glgMaIrSaU3VeaXCYRpxJ/bKcCdl+uVfrQib15XyBSJTn4Xsr2c3G47J9ZeDUWi5
xd1wZZHgOnl1MfksQr3mH1MYsKYnZGDlDI57gyQC+HmNU4knOIn9ztykO7Jylifz
n7rHG90GsrinPskDvO/Zh3xYIEZ4sQmCZ9xuiZgRonB8JaTRKgGnPnzNgJq58BvB
53zUimpZfN+WKUpVLh/INOy+Vfe4X9QfGTt/c1l4r/A/qmbSHFF/Q849oHN8NJTl
VT/wrvbkI8RE9oB44QZK1xz/p5pTJmHob4VdbuPQij4ZOVUMB761OXZ5bV31i7Cb
5jn/jxQOFm7o1iR6Kt+KEkMKBDJmnjU6YOpyc+gL3rGhKbg2NYDmVF3y4WrzYyOM
PCy0kmefXyuG1bB4aivzJJNT1mBui4yeGnGN1P2jGpcncf0W6iTcJrz/kSxU1INv
RsNx68IxZqe1Ax471K2zm3npwFmsWzruSQMMx3Y6VicSIILOXwQqlpIVJXwOBUS0
3RxtUTKxnaednjsss96/9N6ssjmh1aPm4yOUR/1Kk1552Xv5N4F827Y3/4mTl9w6
Fm21u4f5zEN00j5GuExEpmE7S3AnLuIxc/CbTEWN/HxzRNvEVpLWdJ3WTB/wPbj8
/lqZKuSpSr94MmTvK6JkKOEV+o5zQHHAugJlWKWPd3V95x6pwC+kBGTRT+K4kx86
xekU68hVz+oXoKY703h3AcLmuKkC6E1xFV68B8MgKYJ2n5G0qLzcLU2h24cVIhiO
SY3hp3nkoxWU8oKa9rhj1/926aH70PBsF3uVIkbVJten+mtpojwKh7yQnq4NEttP
WTBzHQgCMKJiiwtvja6s4oNopJ6fgSPxotZm1BAkaaoNbafPrANh2hYRrz6ThIC2
Cezj5cPXRzlTF+/hGD3VX5bkj+xr6653/9Dhcui2OusFe3TR2il++ZMuMMlMv/GO
hhOAlFhLvl43Ggb9ss7WeSoLfKNmbfpg++A0MLhjxrZ/ndhL7s/a4XrWzMU0nc5j
wSkOaaGunU/3ayNo6KdGMNHTaiu/BnYy5eY0SsymXpwbxcnCPSbjPPXBvABQqKAr
dy155VsxyVRc6rDkGRl7a/L8ldD8CTZzQWydOJNRxTqQp4k9NcvP+5VprhZurgYm
FuBI+0sb4MugyH1uxU/sPV80HSX4BnrN6jDnd/UB0RpsCi6sjF+v/xbOFjRKQyTO
zUYycfJT2vEFn21ngn+v9jBUmkcFbOXF/EFPbzZ4l46s0CnGxNFXOoL5L/AzBuoM
RmpHIcL7zJV77Rb3n25ZGykxb25Pt9nLNIv4tSdWIK/PjOf+6SgCl2xYUrVhtopa
n0nyZjehbpWl7hsIZybanKeHGdh+MjElH43NZpjyK0F/PdS3V/lQSSClPYRN4XQC
/ed3lFh9e6f1PTZud8DFHKuMFoqIF4RFv5BTTzsPwLBZRrnW2/i8es4Qs6H/y7tO
PwHlxuj+WAUDwOOmNMJZ6lOj4MPbzsBqOpYr75e44V02DEUFsp+/mhgmkFO8iN1q
3vfNB1dO0u3Mjd0SzF3H2HK16yaqmxyC0z77CEocNpS21UkaLmjl2ksxsYqylpsH
xFncxlJspwTgdZ3Bghn10SrzLgHRKVeKEfcQa8ujjFMaRfAnxpmR0dV+hZcC0zR6
VkvQUaO5Em08ly5PW9vJdOgQ3AdK31OPiqaw0VQwuISPwEvOTTD/mzpulW/w8H3x
ne69NiJUrTT9CS646efz6V8g1Mdi/8NAUJ5AhC7oqaBdiRbP8LX/hlq/JMvc2be0
muiTs/BGUtMVdK/2nH4LYjEP5WeYJXnC7GduonfbHuax9/y8IKmB2boH8ojFCvSe
J4wm/wDgHjLIp6UHzx+jRUq5iUIsT0vj1OG1PdFkoWekcjo97heYDVnbEZUG2cBp
BLR8ckng0csvWEQf8xb05/FVcj4Rk7Fp/cDTTllvKytGRTUK1NGPI2Q8QBqLGgCU
dXJe2YyKe7fyaks18ziGms2Bue3v+L29QKvRJE9B7vrIvO9fsBv+viEyJGCy2dGX
TRxrfY3AMhjZEyXVTl5G7gbIAvQ0SMSMvch8VsqvcXIxQ6z/2egy0SnH4FBJyQiC
ggmqHYfhVukxW5I9Wnza6CUHEbK/K2620tIQUV4aVXvTJ9F0V/vWEVrBnMWGUpf+
FCPfgGrptL3pAAy1uviPQ4mRSk6DPw40I0NLzZkTLQhmuTNWFElwRVC4xq3Y6dhJ
GSD+UR/oQel7O4x4/Fkke0/T5oOS0BOQXJKqf9N6NtQD8AGfkf+tSUUCwDfjvgqK
S10SciNrL7HygP9zu5FUZ059NJcVwATtwt8H1SlG2ZEpdN1AbbCc8xD9qjUBhjJO
TRGZCIZLeGhxnrY9CYkmJbmOlyF1zfODgfegyni11ltZH1BAuKfIuhy+zcvpGNBb
MuWJEqH2qKAOXQTxQzYiAZUeSLrj+uDK3Moz0AQzvBwYheK7T/lgGy2QP+QPNBAV
G7Ft5EVJKYDZVpvAaPomSOWig27GTGkRymIAXCJ8cEPUENQg0yl4FAZLdOq/F8xd
sy0dGnC7gWAoy9PVO9IQManlj/QrQTIib4zkRG5fxLjKtqPMy9I2rHIMX5GAinDl
D7mjbuX7uaGh7Tdl1Y2TemwSU7F0orN7S6jl8oQPIOvbnNhCgv+PO8YUYDyhUM1I
iPIsK28o+dGD3zbeSZZ99/r6WTfblK4M5MbyqdgVJktvHis1pUHTPIQzX9CWgVh1
xyaxyLBt1w91Wx5kERuZFIEj8NNPNzdnrybrKwXlsAbyB0xyNsiB0mVq1/yP99sE
JihuE+kygza4OJK0FgrySZypilaQGRWTJMT4BHNCMUyxhJte2YZ4PoYD7NT0a26H
fH5ECBSy44IBL2gINE6JTgCGe0toOerEtdyp9zFtccWJsuRNZ4FAvsWiRUx4xMnH
QrDJKazDCnc/A66Kg+zzwPIdOZeEqCHdbfKii6SLSTtF/aPn2l6AYvWtqpbeuuXM
4Rx3qge4xjNV35/A0wK48//JHXN367cCsFr8hcx6rJOG0rq1bz/Bw8F21heZVLFa
A/44P8NplH38xoxd/ADEkuUocqXzzzD+jgpH/BX2v6FFjMlRbYmFmHsrtxznEfZq
DEX/Y/120tleGeEgH1qPfWU8FUsEjdMrCOE0w7CtM20c22E1ToSTxq8XkFlhsoDK
MS3GdfIdZPSyWanMjY3nYan60uwHJVSxkii7q62o9BDfG+xLOsupaUW+aF9ucvZF
T3DPp6PpeDUcyrSei01f1eCqEhGfXwbP77Yu03MIdQCZdFzFeqNRA/YTUVImzV3O
L0KLhy1EmhD4bSessJw+nraBRwwLQXoEa/vXhgNZlO6ubD2jWFr1pEQVw2sttWo4
obNdtTfwPl6zyMC6gL91n5mMY7w9RdJtJuprHLxtJAEt252+jRUg33tYSLbN5Be4
MQScLMB1RCXJz7uCWlvtTVSXO8zNbBRQNnMIpJOKXBepumzdsVDyLX4IRMG9hqVE
rH7/IyxujyXcqy3qqlNXWh0+v7loK2TC3vmeZ1elPnYbX/PbccR38r58bOaz99hX
Zpmkk9g2b8Z+GSjLP/L4NU6r1VWVB7aqTw+LXj/H6WdgmP4SXhfkwWoKrkfJoMRY
afdcxam4wEzg4S2eJG317SdREbt3l+2WLWAuGSlIHIUA5lpxbilGDpwIw12dEC+Y
m+/Dh3bLTKqjzgnme6NBp8gQvyDmrbOs08h3+Oe8Qeutq8nWfunwS7ZtVR1Wuwg1
tFfThlZmY8Vax5efdcdspWvo2BPhKE1cx55fIjxxzI2sqGrDIflNYv9ACo/vlCuT
FVfkd2xh3Mzjfo9avvZAxa2iTjqy6xIkKhumQORoCPjrcixJ0jYIVN3LtSQ9kmhe
sd33eAhb6cPxe6lhEWCRL7NKxhtGA/0tl2ebEewes092YBgJU3A7HiK3skODs9VD
JkMsGVZBYU6EcMc9BPs0qjJac9VewVte2aG/s7cP9fnD/qnN9VBAk/Ibcfxv7ebP
OCNfoJQIX9dTfS+RI8cSZieg9LGLBWqlvjARfWY3pvPPv2LYXqNDKDbi0hkbhlDQ
FAu6bL7Vy8p3UOUZyydQxowJnKuXJc3ir0nf5VjScrQabKImUOTI5T7K4xuMDZVb
BvZ+Z1MtYfaDXMn75G0km1X/sgpuuuNwiKC17jmJRmuI/gmD+Nroc7scL5D2DDr+
53/CriB99xJSfE+HUl2XibvL0WkooJfuAf8JJGmM3yqtjxXhNF1/mbw20DXVcmGF
dLYyxRglYUm9YS34/NtQ0McjArAQKCEVmliqeSCWkAPKxaFwFr+UE3kaj7r0dFD8
QGCn9ZB7l1WBuFzjum5vCg3hY8ozCk/LOyN6FEndAGK1O1HkRw79csDqVCo+opNF
gDF0MZQkG+Gfp4ItRs+MAgzLf4HuWD7BbsNAKTRA7BtyLyv7lK4xUcwUJIbmDNAV
XOkiDGzFtuk/pul1sxsmf6t25Hb2idV8jegJipdpBg7FCMeeKpUhzSUPz/a1JGTS
0/DKXxAVavYyMOy63swTjyh84LhlvEQjyGaWCKWeWIQR9gzaw8ft0GL1s7MTjf3B
7E5Omi2cTqOMxNzBvezPVBxPpSXNwK5pEuljzciz4iOfolcgp1AY2Ifo2M94D1Tb
0tc8JXapbb7EIl42bYLggTGK573TOmYbsKjIP+VGCILn9ToCkq9a3tqaI3DHsqNW
YV+JkR1QAAJUg5rt7bifbpnIbxcVFkez5jaI54b6atR+LmLXi4/YDA/kXew625+M
wUtadVE7kpxTIUNwKgJAyisbX+irI1yEqfGDJU8kjfz3Tzh62QzqoE/TjkvwSqDI
cGfuZkvM5JkixXCMye5IsFbOlN2Wgqkp+7kK7BpDiKVa8cglP8DtBAJFCh9OHoFt
R3gdDZaa8Ti/qhLgKdkLQlpcCEx+nUSy4yEZtM36kfY9eTYoQFuePWnCE74DGUx3
11R19HC9DuhcuOru5ttxntHFPJBGVpPDzcud4HbaHcJRgXZCNuZG57u8jIYDnbcM
/x+hWLVnyl6hLPNHmxFXmbVfVsoexCVy1rK4atsCGYt0JizoJy7LvmN68TaGLJsg
cciKOmv1/fe1d3UFkw7kD/HtAaLscheQW5Qhr7+NA4pIYf/ViokhNqP9ubWws4SN
SYFYtE4PlHGAJGJE1tmKXiV082xqBIiir9/6kntvEyAdPIg7aqMWL6Vq95AdAMKQ
JAeGCXzYGKk7DDzaSSUc8RxJ3aGtHfJ3Ox1MhqJhsNeGZxNpS9yr/JyhAn8TBLuk
Niyrz/yLciecQVN+KgmHgdMpgQYxZd2YtsvvPTfURih8m7h2R4AVnmmhjoQkRcMk
jPoqtCNlGulazuqxNE29LYM/qVb6J1mV0bgxbr/C7eGEcHFx9leNpVrTAImGU69j
BgBRCJWPYJPEXUR3bVlqZ8RFJl4ZuZ4u7k+5pIAJAel7Ws0pvrKe+lGek9p4jeI9
C1ZNETcS5/rEdAna5Uhio7BzJ444A5zG/O1PmHaZjLx6tf5/LwTv5W0j1iLFtcer
nKONy0daiVOEtlqJXVFNgD7eTcGfgYlZn2DGYcgTTfQaI86Tkz0AJJgHTdzhrf6s
J/LdikeCx64sKIfQHsAY5rvRigzf0slLDzcFKqXME+z4KCFayjAXRQrpQLA7Tn/D
6uzucolsYA/TbDDdKXcYNrPCyibHZYhTjrTilfJaWzgOu2TrYGXdbZnvr7Gw2TG8
zYd01WKZcuk3FZqyF/eKFpEYtQFDDG+mYGVaxVJBkDgk9w60XNYxrxW35aAjZOTZ
8bZX183VMgCebpY91QF7HG993jDfxnx9izBLNfk00a4ENG3H0jirkB9SPC+1Kg2Y
6qhzWrkR5W88oAcEE/ceV07CL0CkQ8pLz/oRQZSFB6KoDdjCYJ+D/HLaO5VG7eNM
rKNKb6TrT0pVBu++UWNjoKd8RL/EdHHfP5gbIeVqPHZdpgWtxyPo2+VAOGz/pvV3
kJrwLXy6hTsfvYXu1aoAw294H3z1nKJuhxd+C3U5pSt0K5ciGIJdnMAAVOF09kOl
EophyxR9bvNUrKads+ZtaxzlQE1uS24f6pFQglEEe4DKrt0J6uFJs1svXlagWiyd
uKVdb/4cu6OQ0ZXD+28UbHcrXjQW+KVonZvNujublfo78pH3RivJLTs7/Ktgw6Kt
MlwHxbj81hZ4+U9T1sXYQ5Mb6Mf9gP7jYs0ZCjIR5SuaggcYbm8z5jHGvL+BfxYY
CICPaIqSmqDwJYZNk+ju5vVRFjiAXaa8W9jqiS+TbL1kXhUV0OYcoCe3PJLppIVh
x/4SOg1Q8gEsBb1trPp8qHmyzp6IWbM4+7T/Lx3ams0zHhJ/nfSpY473ZH/CZh48
yCbPdj9v0l9Y0K2HkpH5b7zKdopf0B9yUH0NzsuC+qG2hOLanxFVyjdbg0cJMGEx
FSoFehhZXlE2giqZYuLLGLiGi9efna2RQwgxFhtJhchBmBpRRPo95rDAvFvl6Mwe
xcRkQJUvqle+ETzfaCGWVTsQbV9xnZwlqbG7ETQ8JZlq9vxiP5tQL/VragVYXCvM
95nnsiQhhpw+V7wiSrDy0RPzAIxM5m9L3UwUPWwcNZIlPuGySRyGNGtRCYktjlFO
kA8vl/Ps+T0RWBL5txfKvy8V3A71ogtCMo/0XtMiMRHZIbkRyiGPjLqtpS3nUO5x
giaE/JnKVOYJShLg1DtNxNO7NTMYXF0mpKetcjqaUV2niZg4xvlPpCNSMZ/5Ro4V
qj++GUpQHYPubtXfXplLHDYIyXdciUNgMyFIPaa8+zHXioDV2Dyh95ZqDz6vm9g6
jBty60Dmub3QCrrmfm02k/cdTNy8ESWmuRWN8KTHXWK5eezklpZD8hIqPFzYTMEF
h8AbZm0v0tS49med8Ycxie2N7Yu5a2t+t6oC4Hfk3jz1n/pGBmuINrmOr5lRQ3xD
6wTM5T6+tFLRwyE02WE6dDHd08vooxPoYMklmjLZerr9uhsLiuyhVkqMLCJ4jtSj
UX/PrO5vQpYWhyAfuqSJ05Xxts/1kfIiC88svfazsamTrjUwjdYDQzFFAQsbZnaH
XUK/lAV7LXkLM/C4MD6HhyBYTrrU6umKNV7ck8eWNlWTwLOkp89KzkJp0lWM23Sj
hFt7pp5QzcPmDp36hgOCju9uV2HqL+Cm5CdPqcT3HEdFk29XbvDKKFKIhgXEJjxL
guZ3VcYveoHmWDoJhDoVQlanw3JDBygfknEZVB7XsMpdeW30UNNpdjOfRC2sxjOB
xLThm2h9FaOXIju9DRoyDvWdGrE8RZbYrVa6MiKEoRZeCIzukk8GZdO8LibkhFqq
xjuifZjtMGCcwDqYciCaYXVfMxNHL5AWEkuaDHqg+yFXgCM4JC3ozAavbnk/0gLT
oT/3MlIzHWruoqqvNK5hr/vUZylDuNSt6TbebiRrYQy8nDYoY7s29KEtJLKfUHiE
60Mc7MfuqM8yIiGRxfdvP4bB7YBFMiSgMpVOngW0yistZxS6JHoOjHvLJCXX5CKh
yRgGv2lYZRborthhGNSfWbzuH3uDQ3hFgq4QBFbr5i+JwrDI/W8Q0VVCMRztP0IS
j4qldfS4tDVskM67Iwrr94A6zmerD0x/pLjKDGmJlpD6c/vInU9sHqWAEXueN/9n
guvag5tXz2hqmja44S5paf4EiTNk5zYlhZzFfvobaXFRnlc2xHK/w8CBOT2y7qwr
lD0WsclMyLVtOQTD1JYyMsr8D5dBK6P060h36+7tSuotqqfLyyMNZWEbhasakqYv
2N+qz3TSQxyzVwRNWr+prJ7YG5xfcdWIHscCiiWBMMT/dlq5KFF2dliHTVa4Ex6g
QZPW0rqJEARETNtM/QxMOyKHQi6XyIhIN1b7W1e/XtONEFi4kkxkoUHO0KbjAt2q
NGyCfMMWE4SOlCKz3wCs0JkUX5/f4Pf5WJCc6qHz70E7DujdsmKY9CtVweeulO+P
pSsK4QKTJHvBelroexQFyZmh00beMIDNs9WDnp48PMp6HTe0We36VhoK/sMD5l7g
xKrRmSmiE3+rW/lYq9b5OvM7kgmQlQ+iSfOKUEL7jFvHgE0J5CnweVxpAjvqTqjD
Y/p7w26pIvFiuZFrTxT/b7ubJyi3PfZ8+jaVSwUTi66yIQMliuu3/AAhJxG6d2k8
3s5nWC2VrYkVCqeILA7EO3gSqDR1543OT89fdMzHiyVReU7/eeVQxTfXPcMToosn
6kjkG1pDWp75gcnjgmQD67+PYcqpNNGampWCs2M05D8KZ9Rn2Mh3SDQ4C6LzCBr5
LWmJuX9vNrjXpjudEds85eDowzkSMRAtnCLdAIMkJIPVmjh2ZOI+wU3X7BnCjj3V
oimPL+JOfKggQeKTgDHJNajZvZFNLVgTbSXN95m+tWC92GPPfEUcXWK+LpWMUATD
znIGkVqWRKnBN3zWntHpBT/GGx1EBOfszPZSIobWPtZAXndpoWNeFHTImVGOChHq
NoUbXQqn0Kg2ijo31ja/mNlnAn22tgLUQDSRYAzQn1KegSJUBMfF+Hg88HAwve9t
Abz6mZUfk2SZuFnUWySVQ7ZVnlC6bGbmtPSO7WiNX+6ajy4972zBSpdczxU6aaZ4
YAZEI23BRpsOL/pD16xuInXvIybrgdQZqTOw/w6D2ICmJdMghxR+pb0iGsIeE0/L
574OE2mJR4C45S2t26ZTzokOW40N6JfFTIBN7/lNLSKnC4sI/mS61LqEF3Sg0JUT
hhl6SZ4arCHMkOwozZubIqoxX4f6U+SopPpTAFnQMDhTJShUs6OX/in1pD7bdzTE
GvagSlMuyDoCpnsTFnbFqftqphIcbV8G9hlccdiBriTQNhdo7Kr5UCDRM8m9kuO+
8tmbfbtrTTQuBSC63QiCHZQl4Dl6MmcomSqk/rhGD3czk+jRXmUDapEslXnQwLJF
LLEgsIVN7+XRzIsU7hqokRS88e4CAvlevtNDTcDMdyVvu02ZQuVSZrp62pysRM9S
lo/ucx3Th+dZh0s/nxz657GOjKBjcWGsw6kyz01fzhu1MAUaPDbLzoWG6/uaF+D1
AIbfPIWGZ4JiAlp4M1Fo4/ZRQP1lFH2juWnfhYO0oRs6Jk6rGCaEKnH7Q9/J94kp
uYQaPpCm0c7lK/158aQFe0klHLTTpsSVGOKuiaMgep1pxHmt3+n6GvNjA/gT3p2F
1EAt4lV0c+pal6RGdJ00m02EneLZOTwzRtYk5EStSAxUgdXypzLrsVC3XwpX/P9R
hRCZnXquRN0uuM464/ybWz2+4yqtZ0Wxm+A9aRa6PPk1UApX6eflwx1UyRQumvLl
wWSPVxmAyCQ8PIvbUvnuxvQ/Li33wsS5HEvhjvU8RaqsQfAN0n3wwfKliYsQTxtK
NWHZp6lAA3kjlrfKole0KVXtG1swx5j2OUN75wpZKEZq5oQQOJidZ0olY+zx+WHe
sIQzHzBNkVcYCorZ7fuCqevc/Hyx76/wt1i7LuynJXpLi3bqwvkqqAsEupskIqOf
Y08PoH4SKVnuiOmehQvVjEUGfBKT9t4XP5S+FL67eng5UoEykPForu83tAdfMjV+
alJTWzkLsn6Zh+YmQdM2L8wWqKgQACizXsZst0bTTTFae9JEUvmswcrhVTH5sgTz
DBPxDhaCXKTIAm4YMIIizQYYfcNBwxKvR8it5rR1KnYxmprZATB6TC5vYxT/F/5k
GALs73+BS/2ffAf8ZBlmF18SYToiD7Aew3lGroZhpgtLuUXx6faBEGqnfbrXe0NY
w0sbEtsjPfu3HJIL9Bh4kb1siJhiD+4oCUwdGe8JXZ1G+rB9kklKY1SHnmpflkHH
xhWw2Nt3mUrkXT97+NApL07S2OY3j8cO9+/a9+cb5Q7D5qllQCgTvS7TSL510uYr
zb9+gplrLuVgudGjXixUxRmILquHwPBK7Fz5HRYNFW4GZKjC56juoc/oUH7hwk0Y
d7VxkLYykyWdv7O+6rIiSNec3zCYMCLTJ5cnvirg3INnULb+FCddiLDbJ9YLGjmJ
ay/GOMkH0+GURzBA3WzqDC/caqU/tJwz4djAtyZAI2Ts8jk3CUoUcgflmql9bhve
a/XemTBI5omwHt9g81XTtOjx+srsXZQ0/1+PCLsEuPBZgHKymOXQQbEDoJWXXhhP
b9tKlX3PCMK5EVx4u7HnUUeV1LD24FDbhMzRmSxfHWw4lWBv0orzzi0NVbBrmBLM
De/iv1hRvyU/cPGLvvQQb3VAN0oR6RZQSmhxfRukYrlgD7BNjrqoqypkReQDXBfc
zlRQOnWH+IzWLL6w1xI3fFq47UkEORKYuA1L/CcjohgXP9ZnDRIKSdxcVE3Lf8oB
ek0BfsiMcw+tY/YsorzTXUFetvHbNFLVnowg3zfamZiC68W/jARY82UaxtzY30/b
QrZJFH997LCO2iPM4ySVvFogLiCEmZCoLUWT+HCNj0Jl3zwl7Qgr2BZdKsFpGmVw
xHItu7Lh7XmRQDCo20LwAYbmHFbVeJ5jhxuBl4WXWWeGkmNgXYy0P8lWs3ZENT8a
dvkldNET5QIh35iQgobcdN95REo0N7LBniIJHlCxwrpBMTsB/Sl11eDWc8unzUZB
Rfe5ZZPUoatB3sryewW4mtC3lh8eE1ZL/qD1WO56mXnO5Pjw2KOpeGj8yo7zochJ
2wQAYWkg20zi4aB+boetFxef3udKoDLcug6rtU9FxgqzIOeDfY7xqzlt4r8SLyK3
zsXwIt/1VXAjGgqjI5Ma9kFkZDEgrfVVVPxJfwvgC7jBXT+QUUxUVshMWcoykXaB
YxWJQ/uqNYZAEWHISyeTrr4VxGZl3/zWzLDLdqdj0ploco/zIolHXzpnJH8eLy9R
98gPDGIxkBk4FoswyjXLaqGFR2AzLnwtpsE6D2ir/KGljKiViLMg/dU1h3d0SMWT
GofQ15b4XBBn1wK30XptZXamqRE2arqlsjDzrNb4RZCTdG6fc3bkSWs1IxJIgF6s
JEpN832kG33ujY515B/TbS3Zz5vYFN4/6SvXkK42DfMVw2CXlnuj2JqkYoYP6oDf
yF+A/n71UX7FkbJHCC+30pc3mXOjqegRdUVkvZDBpwMVxtg60M37jYXAF+IQV0zw
GfkFA2HjX5zkPAH+MpMu/ERIlcjofVYb9DzK20gY3eqZfSmLnGfaHbB6F2BBR3J/
LM2h3oWcA3JgK2qGEiH5dLMImE4gXlRpan3DghCmO1M/qOlw0LZCsh/i7wuBYjoS
Wz698plyw8jAjTGA+ia667o5CpjW9ELw7J3F/lUmkYgkuA0HuwzG51G3V+ZLJaZy
6Dua8//jtC5wP4GcHXt/whnY5sQ86QnARafp49uHXUIt7VGhfAPOvg0zZOQEsj+5
WzjvzYnEHXePs5r67OPy+DQKlHGPXFqsLMtW/GMiiEEGD20yP9D8MCqc/jGu+uuH
05HdUV7sYzSMcKAGyJHr4LfiXRdw8xmTzhOD8JJ2cjefpqjWP8b5iB8AUbdHsoy2
Ku4q9t0OoIIJuTNJD7szYwESE8lLWD+/4pZzyLPyvuy/MeG8lYkARHqJ9f3Dbbby
oDJ2BO5XP6os5oYJ95O6BRLcNPIRXj6WI9bqoyfTigst74YT9N23dETuSN7/1c+h
DA5/5kmvbYw0fbBbv2upj6RhPVg1sZcGZKxzICA9c1C7ADp3CdAP7tq1/x7YpkQB
ZloTL+Q1oM18ZTtycY0YRkpHVvezFvYbMiIbmDxaUjTzm4CCddM//q4Rnh4TX8PO
kop+qf86zZGvbsPdLPGBw1hNewJRY0CFuqKcHmn7mg2/uJwEu/svqiZvw5wbvQlL
KWckC7nXPfJsexPfGTWDIBBYqStJgazSzd06qNAbk1b6LTk/CA0g5XNyl/7fjBo1
Ya+6xvDmi4Qrv5YSpTiBHaGPXE52EMytRz3Q6VYzWVg7lGqo5kvtjJmnnIP0N1ll
OKWsru7w3lXXKRDV9M3HJml+YCn1RbsBJncmHtswbIWOWtviWfCQ6ftzQr5N4cbf
Fegzvrhn+h2jeD8cR6yPp3qyT9Zvets8XSRl3OhUql0ip1oYqJOiemOIJxyXj2l7
3fd4+6xjCvzY0/2seYYisMZUXtSEkcTNcleAxGJm+ukFg8L87wAVX2BTvk51GtxS
yTLBNGfCjJD2yJkX/bLIXFcWRZe+W2LQi+s4G6XgNwskwbo/loRJCXzusD/J0iuU
hcIPCtsAhSswzRYh3j/Mz528MZFGADzZDhuvqoauP+wO24MvY73wCX51WQLHqlrz
vvHcXZvFuUztrz+WB2m2BczyJaFWB7ryIaf0WO3YafJu6DMphkfVuA0NkJJI8rGF
K2wk/0Rox2ccfhji3qqr4xucdnB//vNqYyVFpTWlbTw0EGAgnMztkcl3a+4nVStW
NCm1fcV4W/VrX5Q9rzIhMkS4dvnGkK/fL/0WbSOKH2as5Pv+lfAZIzvxIRFt+dkJ
bqk7/9m7xSaQOAMfK4l2TOwjh6M2c15j6pLxmsCcMdpmXbT1jnfxT5n4T1YGXCJH
GPhcJjJ7eDKaj7L0IxzbbRP8IyapJq5lNsyLv33CzU33TyGYz/lGQvHYa981s7Cg
SuIhNmGWuohiBif0T2KQcdozLCwLD4TOmFtc+vVLNpzlapC5BvjewC3gUgecBGUx
x+DngMcuQ3J++Jro8Q1w3r85NYwN21FKY0gVaJLZ1Kz5Ny9rQLMVpYOmv9/jpxIY
lPiyiHMWQsJ/fpkOZtZGi6YkvBQR2Tt0g6PTOD75PoxYcRtpLFauh/sUuhqMg0W3
FzkrX3X9SK1SbVg7cKDCjVxS4P/3y4B6RQOE4ljYTRpUkXHadqPPp8q2vkCtotwg
9S8dK98wm58+BcmybLFxnoZ3P5Mso2opTD/V3/dw3h3yqCL6hyK22YmeU+I0lCVm
pQqX+dzbu0Kajy4P9nrugTZqwL4YYTH1zrJgQAQyomjgmvj7kIAaipRSOMqE7Yr5
+V/agJXSSoX87oN9FL6ilHCznRjhzF0JfSQnK9JQHA0OBTwHC2C7Hrhvdezdfe/i
BuePNIBEVfL2hS/mh104sG1NO16kER+6+LpeCDX96lAHNkpwzlMv57Te+M2+W0YK
tNunb6N9XHPWmafPbJLZ+DIrM0uZ1X2v+cMb7MKLGSALTvBvCD0i6yUdJtb/sOrh
eBfz3PdkAnVQgnXRTM/YBMTyZjUrWn+j+Uw58cDcTEZ+F15rTx8sHBiNz1xNq25i
DRYMOvO1uy8giCcp1GVtZAO36lcA7bI1mLnzyhzuXzjldo6TgdAu5A5ZGtSiMVJm
Fjr+YfBtqYEpuskXP0H9FORVHDNtvkya4WGY1qgR6OgFDjmg9SpTyPC1RIctfUTV
KUqS7b1yzFnbi91AEgFqNR0VxPNF4qSTgQlWK01x9eZbFvF1uEZ+Y0HpgMp3M5jN
UdJsaRKMqD4jfhWWGku+pkX7oBn8BRRK8JjURGyFKndDdcWk9530cQLXGQEv+Xc4
C5faVh5VJqaS5FHFpsUQKVC2R92XScWuI7XsD9uMF743Tei8mDcs8yf+AFUQ91Q9
4RBnDdpn8kMp16c50lLSMmuQAabqLuBdBrPrG0ukdcsBD7a257734DvB3ZlNIYZM
4y9QvHSl0QSdkh4GwbYx49QgaqmrzWR/kseb7fned1Riv79lA2fh2hvEYyA1JxUg
`protect END_PROTECTED
