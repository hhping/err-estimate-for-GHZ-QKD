`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5VrWdVBrBUKa8xb0zBIDxZN2DtC5BDwoSIDoL7KgE7xPZagbt69QDiBTBd61t9LF
fNoVrksTa6t19IzXas9mvcDhyfubCkpv81/K2/ioZPYaX0+tiYNpj2vDmUEYnIDD
j9AxNJeUKi7w23dHfXw24uyj4xMdUQB2HjSoMqr4Wazf4pivyc9Mb7EQy1q0dfWs
mz6i6eZtgkR/yBES/1nRCuEFBoUQQgPUeuTbZNg16BCSnlCcgW+H94kU9LQkNpD4
y0WfJyS4KRIJM5K8Ontydl2lJFcuSuJ/iIocsBoxd8oCRu2jDyE15gFBoraMG5Su
zL16V+fIh31IT4bJdq6AQ97UNBqx07CgMqWojIHvCuXVD0sX0KZ1Af6AjAAKOb1C
5ujR8N9qXxW2Czol/nAliAlQCEmIpX2ISVpjjjFNngtxaBUcqqIV8Wj2dtztTyBB
poT2yYTU6BmuELKezvnC5mdmIv61bUUeNrpoY7X/OG+81LfP8jn9cK3ie6sfw+Zc
xFnsUWrF6uUGxe1EjsowditSgULhGyY1rcX3HjbhTh003uf7DyIQyivexQRdAOTF
i6UjWAiHDegX+FKGhP6qRhN8jyf9RTvPxulFOrNuH4o0rpi6PE5HQNjDu1jQE+pW
zqNnh0J7JsauFr1nWJXFyh6RmINxbP/Rdo+9y7D1MFyf/RHXVsYQcgQNJOHpMuiY
cDPNczI/2PYTaIavKdEGN4xKFIBGWJ+8heaJG7F/phDQPijc9/lHQrleMhJ5hBf3
iGwa3k2hxtoqjYyY1Jr2+H4MBpTeOGAlli8SfcXe/12jEu5SuA3yZvvt919rVw2R
RLeMr5PPNkZuSW4qMNjtMGQM/flJBZyhaFYOklr21PUoIbYb0g92v/hsmRKARg+w
IXGnbq4ks8bAId4MdZl1DbobuCdT64vbLF8+MVfgQH6zmaxQkVGlM7aAOyyZszzH
KuAdV8EbjNWC/aapded0A4s/cMjaJW8/MPI+0dEUHKX0RJQ0dB6dGc5LBIeNnFsN
wKOGV0yiGJrw/BhpLL9VEBUxu8xjD+IKfpiJMTu6ZFhTqv82oiVLq3dLtjn0uiQq
NW8FDlb5fT1wNXcQuWIumP/vW84vQERCZHFElrqpql3sI3gKL897Jt8oewrGb0aJ
+ap2l0JujnwaP2ivudZMIRXz3j1jfCW4M9uGknp815LHLGrJuiybly4lF7xSGlyJ
K15Gn6J2FLtF9LIU4BSuyEz7Z8Exy/heJY3+DII8IOQilacheSrVFy7nLXmsvMQj
apk+FxPSa0vjSDfA/CMAP7U62eKb8VVO5eNJqu37vHPD1z6z8ribWow5mIxT6ndA
Jie7gVg7cJVDS8Q+CRajil/VywXai5iiknlx0Hinnb86b6v2UtM9lhck7ibjHwQG
StBDqHBvwDERoWtX+5HMLZFVP7u7Z3L14ar/Vy5SMukiBumxkOYkPo7V2AQmJEcD
Sr9rALXefYF2x5zxn56GoKs9mEy6QPsx4Ty9pjJp+gCTEFpDqbRXQUK/HV+WX4nd
x7ybyyRku5JDV+pXUZUP2Mer4btr8uI+/fDfdhEOZmJ6tx+OSCOFQ7PllXAqYauO
XE2CmIbQVE/OOYle4aSEwSZd1xHqGRamrph1akVecLl17q/GC3W6H8PfpCTr7kzZ
Gdh/LWuYNwqOguRhse3ikqzJeKo89iwqAvIu1ysytzP8j0Q3Kkt56p88DZH+4oim
a0l7LRhCxqNH3QTjdBc221207SBd2Q6sruXHj/J3A2Y+8UM3hCCtO0P42S8u1L1W
QGHZNTbLcGpy4JV7pF1nnuOo+G4n/8JHKQQRIByK9AfeWh4DMo4DeYOyW0mNm75q
Ty1rElSrLtpuxTWTjlZXeg388i7WaPDvkv53nryitZzB9tZVS4YE/tW/2lqVW09T
FSI/2cR50X6ztn86pA8zaszlvVgrlo/Y+/Gi2Qjciux6/JlfPbLXAxVUZchJidZ7
hKo8I/154oi0c5wJNPP9+X6y6ygekMY2pjOjgsnxOmGHTybmT6+YfXuEoQv+6/lP
ZMb0z9uVA+G3Wvxj4Whk2Za90+JqyMZmMnmG5j7qzpnUxb7dFuND6hCd0bZ0Gssj
Il86NczrA9r1zH+pps3Av6+l8gV76DtfOSwZRYQcQV/2pMVb/qMgicYHy/4WGKUq
ySC72FnZVhtoULpqs3Wa6uFWi4n6fTI7RNBpsANm597Qfea2igAR3Dv+E/RbE7t1
vYmmvzaJ8pa5hMasWaxYUXX65xdJ/r1oiKNLYYZqARN2+SA07thJF6cByrbYX7/G
lvw9nS5g7ZB/1/OIPhsuGv4zR5+aVMoZKCK6wr8WcdMAsDCzelmaXGa8gUgDSMFM
M6XoG5wi1PpMU5P3EtFXRcxLhFQwKSf4oxWHC6rvSB12lvYiIVLrIId3d5DIa07g
tSGFuA+fNqenWnUki+yDIhPqbK9CzkbXL28hSOn8DAGafekmeeg+PPQzWqj6Cw7b
a8AhYsDu4h9pfl8Tr+azvGcEnsEG0lyLJOk5UNcNaWSB8bC71msWJ8+OAJV42rzO
kA8Rx6tfghZoHCr0TwQTXRHlcLmYVV5OHXpE+d8DIcFu7BqF4cfi6w0pSC2wUvzf
nEC5vKWOeOejjl5/kpzUgLh3fTrliQ90FkhdcMuO23n/Tse5UdEY+vcTF2dAIxlR
mwq0E4GQKIaKJnL23+rSr6MWGKvjgk/sq0djTMPHSq3S5+PGHJXNdhB4Z/p7nc4m
pVhEbvOT6Luvs/j92izPTemDsn1VplF7Og2k3b3mtAjkZWvQOhfaB5/pP8/unYO6
yFGO0JW/yn81q2l2JwulZDenF3VuhJYHC0X0ySv3aEo/QA/4ke+htcJ4w1XdgzJt
p40qCdhy9kUjDjFvIcHzIaDU4aiGDinkUZ93DH/GzXpQFHdrstMSYvmmFKKT1+Ly
Q24cmDzMH+0WE7FgSe2ddfbg2MeFqPeFDBYKEVBgMp+o/hUOQRy97XXNfXE88txP
+CMTaLNX86DlUaRIR9soAQemU8VDSAS51yki6o2ERze0tQrKSwIGc7dRCwVbxPRK
WbY0DpANjUX+v5xJD80sSoivUlB4XyBu6yoYKrudx0MGSlRbjzKzgig/YyjbJdjD
YPS3om7nEA6U9bsF7DGOHVoRWb9ikldqlUIQdUl+An3RZIFARheEL8UMIxsmpyTE
cPj4vTssYzBTdYPE2AJGIiogUFKXUhfrSlqhJQW9P1Ksv+J9jt2OXDBGG/F0jsz5
3omgvLfp5m5U2/HslnSuyZ0o/UNq1EfCyOzAJA4kHmuKvcl3xelBFi4FPoicNO9J
KoAsicRBNCikmH+oa9JRmPIVFgz9fjujCmAQNDtlhJAqnwV7McFTrtqixro38D09
xPT+yLkp3iQ5YH9mAml/qxOm/75C8+iTUMavfG7CUUCFNrs7lV8HQkpHVellQYM/
ZCJphtJs9Mb+CTDtHURUUsvUgdc8dO5UkXnYX0w/pOdNteT3RL7lFBC0+sLHSYpB
kITVT09MJvJWFAx37JSB4LXNHkibhuifo8rD2irIm8DsmTTjD0nDcWOOoadXUdGU
krUphWoEWV9ZJ1VsQEIqjcsHLob2wInrYeA2Mj4GDGuUKB4XJK+As0OHbAM/pb35
QTSHSOmQBenKu30hniQi9AEf+s7ztwnM9I7pRsNjNzv+l0tJEsZqoul4bA3TRvlS
cmofd9oFMELEVwPUuNFz4PcdpXIza7ia2CJVBaV5PiIib+iIKBUgN5xCUsAgpSBt
4JfR5LChk7Yn9EKIh82YUTqmurcsk5FBxnkuJgNCsgICNJKtTRfpjfoZchuxcWKJ
Lq1I4tsrlRtRRpuHQygy2KgvwPKTPXsSN2v2RwfJ/F2qCj9r09UBOqjNcPF4VlqP
5KDohCG7iv4ingIhVMkAO4pXfnWCUMOoL8J7YhEk+/790zOGkBm0AfQpnI9f6QcW
vdNjoZYSjaJU617Wv4HkoTFzxzXIwIjbzNgHjgWFeCsVzcuTvcBCA5b/hbAX6t4x
uS/jZYJaF7AcBOy/oVqGTHo0RokssN5CqGYC/AiG1UBu4E+l2dxilfsgr0+ZzSle
V7RizZk5MeBpodpAKqHUB3++jY/ZpFgDH6ig0GIt2o8bImB1byF5tEpOm9l3sxDO
IMVdku12CInt0reE0xnnMtkzHvpQMlXsiZH037fNFHDiv04DvZ3yjsPHOLSLDt5b
pawGC9Tgs99E4IyzZAuzzRoOgvwuRbuhnTZNlw1Z01jd7pKKgacW/5rtSmkEsmmq
48d4Go+gaGVs95s14UjELLMHdTDpYhCyKjli0YMB9RG28XMCJQgplKkcanifwXee
HcYGemKGg/LUjNU9JmTHRmU8btTRQzklAjVG+fAXhwQq0M1HRIoxBda56SbgJunF
uE0M8ggPhech+SBSCkjNkg/NBovLezH2whGERUWU6C23n8tB0fdLF0jwGPV4z07e
Y3LM+68dfAGpEN3WQaqDtYCaZaGJj6Y3Vjp/QfAXcdl+7zlgjyA4v/TkX/ekSZhg
xBOnHBX/YlVj52BWj6me7KljHwDT9rxWGtERVH+oGyphK+qF5tIJB9vMfzd6krqi
b3jWJ9UnGeRyYjw1+TSZ6R3KdathKsLyGvgZ0k5U9yDPdNWoIe96TBhlLUa5aASs
JggqPFVZGPXaMScRm9pTqHw0yeCvYCub2mSRty3SP6UvzQYtwFhjaKmF8928QIDY
zuIE02/2jiTm5ZdiPtp51oyUI2m3tyCKeDOZfXKV1s9Oeihco5/HAHmelFY7L8+R
Oh6H7dDWNJKaGc1ts1Uo9xk/UmEsXNPYY1eDQaihYGaADlFKZdY7XW288IdV8FNr
tTeopjtWqic6pTLM1GETpV4zL+4KeydXJgR+lcajVx8lwUQrM1dnrQHQSqpWW4dH
EmBTVnfXNtPay9fH5Qxr/NKWywttkkEr5cyJDIo8Qntt3XUP6J2dimEsiTSplFQE
tf08nCV0G31aK95i0A/oru77ewqVpgmOrToPncm9ooybGn/Kyjf48MJMcoOBU7Nk
KWbqLd+Nn9iSsNGQtx1MSMrcbODD7Dc4nw+Ub8F+rHA5rsiC6WPfVn19IDgh/bFE
zUxn4LCZ3LAWjvNirz5oQEiEbUbZyM6UlQIGuGQLE27mAITfjBt4MzrJJcklLF6O
ChVA33xdQgUjH3DYPfMzydrW+V2jN8hQL9cKsX36dk+Wj5VJt4bs70FeDKM9fpBa
NZ1YQSuBajur5WL2yhq5WRScx1XvMiZsYwOqbpYiy+9vhzDY2BMdzjZG0/vLg/S+
So6yRsZvB68ONO9GY3uk6ARjBMfdd8T9/aX8q55T84WzwoetlMG9Xb/FWmQPwNVe
vEE+PWndvQQtAfrS5LcRYrmmKpgsRBsb7cdjdiYLLJ/YSVymE/Gwq2RppuwZJK1F
RhlSdPmOJDTJlJq12JIh5NYN58SuBHFSmjDzIK0SF6feRtaUIZhy4FauWCWEO2AJ
siV9NEcWF1Ylm0+47timMdnkx6wP/QIzbRtr9s1mLtF+RoA50Z1tqTcLD5zExmIR
AycCKOGcCG00HeSX8YMamRKtymiJDLRGDn6lo2Ob9mbevkHDJz7i4VqrAPaLwgII
6xJZ/VGmvhEcVaIIKcoqALMSAdegk+2N8PE7ahTagPU5xlwpMtH6Zo6GOK4wV97h
Bdwgnh5eZKWRZHLMZIQGmO6gqQAGP8DWEGCHc2Ee6Xa3exd2QfEJbplamxdaMcL8
BWf/QvHLOIrGpejg2pFnQux3ON77nWWw+hK9BzxBzJYi+62+mhxNVuIyqrh8OoQt
51JUi67vL492UwDqum8U2gYqvHF73uLWXfdxG53BpZMS2KHhbNX3lni/i3P9mV8I
DW/Y8+GckbnDt2j8OM7djcLIvdSHxq1zaoJ1gqn0sinLavkAqYckMDyYuQbSE+Nt
JUku1eUaI49hKNyqz9/KUxtWd6YRsH+GHEQg7DlKGlsn/8kB+jglE8wTKouAy54/
k3XbdiIIFWiw7Ux81GEh6/+hcDlHhqtjBb3qkDbPwra8Jw4tGPNK4kwLdJKHzCyb
AiAbEz0/MRWDNrbI+R8IppgpQBtmH0+idzbCih6ReXt0Okn6nRJGDAf/jgzGNINn
s8l8ng3TJGa2qomboET9tTB/Jqh0VSKevPliMCBIH9NBKF2tg8RHbVz/tC5Vjb/B
om4A1gAmQQA9BO2pkmLMk/d4Yh7GhO8PAcvHys44v+YUqSjP3/yL95VezNdBkXoJ
XAm0kMqEx8yc6lPiSMJNPDnxAOGJDUlgKPN0II69yrdeqTOuLYeKC+kFudUec1ko
KZVbVfXPMK1229gikswCjRMfPd8HHSNyuW9fXymcecLd6el54RMAWLH7/1Qzw3IN
3EjG+PDhtCRmiGbQaurq3dmn3PEndqGjDn0i64w/PyM/tTRsh0BCljEWtjgRLvsW
1EMVJ/KHDATq2tE/YDehrOWZVzWgVdEv4ZRF6RWFYhMaJQJm9gbe408a+TimPv0R
lhvbafMfgTMUSiKfm1U7AbdgnCmxskPix9oSPl5NoPWFb/TZoemw0Xiz4rxhQ53q
CsQp7afDHFv41CZMM8wh3ertp6ooC/qikaoTIA0yT5FZYhYPD4HRG7LYiAQVmjr4
`protect END_PROTECTED
