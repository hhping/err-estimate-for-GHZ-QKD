`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z0eEhupqP946xUCKUjnbbenC3D19/+bojZWmNgdnj+yYracE5NZWxZ+B1tHrMWPO
cK6G6fRtcyOOeoDrkTpVI4y0hnRekJcvIIh1Ts+3l7CMITaBtcRIv4V0INQHwTI9
ZLiBiY1vhTywL1YIbCGr5LY6p6v+zrZpQI/XGiZ57KtPYJ1M3a57ARfYYN8BIPeK
J31v5hyS2JeAkEETy07a7dQdVUvndvY9847hSa9aYgHS1YmLPjcRHKwjaXnnYX4s
t77Qx3yL+ReF+S96r1G/WegMIKRdJr4TVSkHANlYKVedMVhA72etcmdpprJ/defh
GK/iwhj75mFeNt6nDVZfrsckDjiDhHGJcVkjFfpxjbsZJL7mOF5TNqHlYpXCEJWf
88JD48azDrGnaejaRDYvTp1RB6Az0jGRSmIoebmW+pafzF37cuZXl7MmVOUVQMpZ
dWOUaEdYeKNK5k6Wn9hhX4SiBwHImhty1ZjSkVfAHAv/VZCwGgywDZYdxjgIbGqL
9qQbt8W8dflc7fEGdUkyvQ==
`protect END_PROTECTED
