`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/V+cr+KN/2zqHDqEXzhGtqYxdNE+FqmOeAX2TMffjOH9mEh1H4V30/a4pTzdIwkN
O+scpssNyFQWhA+joQ6jxIGp+zi95u7ExJnw6GOnj/v70U4mLkcWPTw0yEQW2Lsk
Fq9p0fhNdRyfjIJmpE+32HhunET9TjWiyOBY8yIxYYiXrBkXRs3LlFDT9sCs3cWD
2hYMQbmQWGbHYcO0j+yHFB/g/TBSRD2sUGTbhKC81ODQpBNn/DchGE87V3HvW/4J
HQcQc8udSNUVQGg0+lbbejHVWEf3ggpJ6PWNO7dDxhQ93lsHws4sOYqHHBZ94GMP
+7C04DAyRZTHaTDjOB+REh2s5x7nuUGGdlcBA577fsSFfHXKsNgzy4TS8YXGZkgU
Gsl5k679MQQTL3vgVzYumJCZu4bqxu8vMmPxfirkvJ0PNBpfw3mQsGdoGtX49END
IC13/gR5gOlGidBMzcpXngRDe7TCQMduEtHslaSLDirIRm/lTQNkajCpJZJvy0D3
XOD/2wq64hnWw6SEo9ZNdd0cL9hVCcKCexWrogdXvtBNpBgNDrHJYGdDCshgByfB
iJ2ELh+V7WY7ogXK5g+p61FYNS6y65h0xZA6qZBTnjIGY0jNUY/uOnw6woJWpsaE
W5E5NQR3Xi4Uj63DAYI2h8avhCHoxQ3MKPhHCd93NAkZptIKLEi9Nf7hqefWIn/K
ugaBEiXac3Q4/y95URvw6A==
`protect END_PROTECTED
