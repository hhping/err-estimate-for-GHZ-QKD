`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1/QxJ7hGeWAaSQRV62lO71BPuuIXpvQDwWnX8l/z5sGi7Gx5Qyl7ZNBFpSjMuRxS
UAAnIpohWhkVuyo/KoLa8gyGvqHdVo2VrUEsNuJxQJxSFmHDcY4gEjNE5SRyl2lc
cKgSKIaDCTeC3foaum51oVnKah6FMpblpmWZCRtHAy5J4m49iMunjkikpRyDz/ss
yX1aNEbk98335jT2pgIWVfCZvEgAswk2Ssh74Z7p6Ml8bw6wwmekkDCGmTuDDTeT
FcNnoN7fYm1T0wqIIQ9vX2kFVSzFxfRjNMA6eWJPdCggOM1Doe9pFCVlVjSYhtuf
Uw1/XfezoM8n+x/qm+cwjHQj2gqan6A4nKLNl5zsS3XaaykBQfzR9CfJ3CZCPHOt
zZrSNJkYGsVxS9MF5YxWd6Ellh0hpIqLQB9bbCQVaSxZl+MKK/2Gj0RAEIoGSM8A
Qb3dXr0W/1mqrKEWZAHoPYMcf/eGSvpRwquOQJARrUY+bV/aSm22wHQQajeg0a5x
PSmCeJkuu5e0O8XNSND6y3hDGrAzMIVBlxV2y68B8VVenkrNWjocmRm89CGXcjqy
kBrssrugtiGzafBTIzHCSJPznY3ZTCbY+y7V2jFPnmMGYPPWMbAkYbKvlupMyste
LHNC81tD8RsuBr3nXlT3Mr2XwduWSEJlBOcQsULAo7bxqdp6SoEuBQbJvMSYqWai
YCR0P+Ngbm/vg8TUTvFTbffD1tdcSG54x6wW2CO5M/E3o8AeH5PRGDF3Zzyc1H7a
NuT8UGonxwaDACYzQuzDwnMfzPGOK8S+is5LLIXcJSpKabUj2VgczFN2z8CwrNfL
022uvV2uVo9egaG7lhjP0ghlw9ysiamMSme3ZYUbA4Wsgt1eBeGewbFwdE9pZOM4
kFNBAjK2sK1185YZR9XVYRC+ZwShoOTbhMBXvNllaX+LXcaNSw4CVOaxo3RoeT0y
/TXp/3NjpsTJPAbvZYo8C6TJNuqVZphzUyZazt0aSTuZbfnf77O0DQ/eDOWT+dws
`protect END_PROTECTED
