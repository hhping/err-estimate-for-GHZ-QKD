`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IowhH4bBXet0/UMmhR3gHLJz7FLNt4KLKypUT/z2S3j1pOEiQVmKyFuzh8w43fq/
BpGAcQL7o3/nR3FbLzhq0B9XLLzt49QMQQgivzTB5kRlc9NAX/wZ+Ugi+0Q2WIN1
HzStUkdR4ZxH8T4ve4cbyfQQiE9KEUKXmzUVJL2XRA92CQRv2nFJmAR6CYpYBAWw
053OVV6UbK5euq4NN+NUXJCZW12ZV68Iu+fAHGxzW3VqLwgLuAQEuulGkKFiQr3r
m/aOqTpF7oonX6RIN6/Slqg/L5pRO0uVe6nIzykHCy4sAktnmIh4SLgkIp0eF9sM
No7EoZQyjCFq8d1xlg/dMbfth+YOqCPnl76+rZmWTLQUdCLSPXmknKCWXndf2gCM
JBcKRYE184Dt81MBDDZi3pVOaOsYTiYjoqMO7tGvxowEv4AvyAiv54VJ9enufpgW
IW03v+qK9fNf8paDn99G1KL47AT8RLFJ0cSMQ07IYAYkk4Om2UIrurmOPtWLJ0mJ
7Ro/bBRTx3IGx3hg9br5bC6ejisWHiItFRYhkywA/kZ4tPTPs8nEiTqXhRf0e40a
d3YSYj7542OB7Dnt3YaI2f7CYL9IeP0ubqCWIZpA72X4oWrMSdJpIwuUxmLPl/ME
pIdi20UnbDry5pUAibojQgqQux03rRTSFqp9mIwp5rEqWgWJ7luMzIGMffb9r3O2
CVzfD7BjZ9a/iw9brAVbjkZ5CjPjTbZEh+PtyctdqoDRfxde+AeGmL8kJKnjR+cw
ZimSVe/I5xoeBGVicrKs3hUyaAZsshta90t4IxviuDwCuzFAohJQ24H5j9c0WL00
PLay2t+ZSKRUdqhqIMsA/k4MG9J4Bug4ggudTH3daEvfAesUbNOd2H1sGfKrlUni
zGKcPQS95/Mf3Fm8ePN9msbbZ5eY76puMoC5A0RM2QAk8OlQTZSXsGjbapTOeR/6
KkFZKJVENAaA1pW0ckeFxiYc50AUNULMHmv2/YQhV5i9lXMcCzv8P+QHv8IqD8Hj
N/rkfA+FZkAeAY0dOCZ+VFHSftZwp3eJKHZDzUE42prP8cXLl9aQK9YRHu7s+xYo
78jJhr7i8xvxa0Mac1RaA2sGGUwxcAcdgBEONTMyNm1kxiNvy6nlhD2p8y89++Ef
B0z1PJDdJGy14h/C+SvdWgRAGhDmn8FDMiBUfKH4Y7VDeqSnK5ub2YuOuAxxDMJs
5fDkjOiyF8Ik6TsxgV8o3zQvCjq9rlQJS2HnHppB75gdbTLBQXQt/FLi8aOMUsoe
3aNU8D6lN3tTQoiSw6LgAayxoAlxey4JFV4hyGVneXkNAFDKniT4IxgRCYB9aMxz
66yWUf9He2zgYUquKqjSIwK47EVozKyYpuT3C89YG1vC1wbT4Htj9DfVYaDCdSLM
Bs3h3kqmLs1Su+yRIi8HbuBQ73WHKASms2sMngyn9oNxpsJns67eG4e0LvUC6Dsa
eOIguXBpmthhVYnNUJeCtxKyaR0lm8fEiaQQjzv2r2cyzcV4xz28mvOnqAmaCsu9
+nnZCS3QWRPN9fwjuAM0xDF6+hpMrFYlTd8QdTp3yrYKHsG55H3341bV6B2lfTgq
sy8F5xUBrSEAdpjN3HPpTmf+oz6WZtH9zXYHvcZu17UILY+gXAa+qsKGkBNg0ea8
Q+M2Ick3UmJwdC44eS8pyt61d/1sXyrYk/SrqbHqEw4s6fG77ESbYNUc/wX2G8rg
W0AOHvxyCRtICyN3kyhSQxD98XhnLSK+pZB0GAEfwAFuz+Dho2+wjzb00pzAPzJR
FMJs+lG0SSxeEqlc2vBs6BObiiGVxPQWkg/zjqjoyMnYfNSlSjJv4CcB9IznWy8B
9PgV27M1oH3+DoBcBHL6IFddX8NAGsfn3tBukN+IPmeoyd1+Mqjmw/GnzhnV2fhH
nM6RQ43waMXNMmLemBGL3vXBpYFzT6WkZQUoSno812tnTBaBTW9CKdDpU+i9RzD0
hAum1PZxD39iQPnc4/eG4lZcQszZLquTZ4WPFsYu1pK1YfwV1byymRGl8DxVM5C7
eKPEKBJc3boJP5bYd6YVka5TJDcmYKUbeCw6yxTr2g9SzIK3eqNOHTLAjwu6zMQx
AXVH8C3CITGPer8x4ajvWaVyauMqbeRY0+BRcwK+8QkWtnTciPkMZtgkB8eUMGXn
hps1R37pPUE63WvmZFlkE4ycSjajQhTesThcbfjfjPTf6OgXV+klmIYS21hDzF2v
c1MeLT3od/xibkXWtfB2bMf1nr8z4XAdNnh81UDSb8HJRR52ldD0d0AylHXnIl58
0O2TMZXrAw3wTwCb95I0mIgJNKcfxvlZ0fMDUW5OEtAVO1c6EVWDNWkhYytRGdlg
btLK4tAGUOTG3jvpORDQ+bzLf0/QTsBMMBtsl7z1Fa8PrquCnbD4tXoeUFdFgQc0
3IOuyg8zVwQo65yS7ibeF5KFdxDRxgQCdXXK9Ir4n0kdgturU+b0pJKSizB7GP/T
uqDX9xHozfbP8qRFVIffm/eBra3gns1t30qkMQIOxT3D9KqevovlYFswYIBULyMh
NnIjUB3Uz0Rg8Rf7ZE8leGH6qYUorPTG8ir1OmucSYVB7zHwrfHnFpTkRD+WPEzr
0N69lai43xkARNhkyJWw5EcrIYIZWmkj+SUzaMxRi/hIQwms+k5wO0Oh3VJ6coG5
k3PteW1SWD6T8wKv4bvpYFWfKvCBmm0FcpOuTOYLmivMPkjFNIWdxkRwVS/ZNbcs
rxI1PRov1Hw7gS5FZPZPBZqhF1owqbBGjk5NnG2S+EfM3zTASBsmE70JwHKmDagU
EbvME1B7MM0VAY9TTeqZcQn8ptElcQ9rtaEFykxsY0PRwv3fehCg9DdhCgWElW9S
sIf7JXElvpqncsxtSwzxmOQ1lTuARzzU/OGJjKD7zgdol7VNXm49RfgCR2QtEdJH
lNPOZo31Ti6rnX0mSxCTBvNQjn4b9rcpCNTwkGT6N44=
`protect END_PROTECTED
