`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cHAzu7RT2nU/N7pPQ4E9x2WG6LgoyY9W/5oto32xVtB18Jc8bu71+PqgKonZzx3c
gbTbTqe8GSUv9WDC6GEu36zzKZCYT0Tipj5qyZNJE6cMrpovATF4ZAXhiuqGmpwB
LDpzH0ey5aNI4q9Aj0tAHD5bzLBExPHOUys38Bh5R+IZdE0lYb6A5rHK0nwPLJU3
sTrtcuoZYWIVKzcw1wDmmaqxXdejRa0u8hD7gGVCn+OnFNwXPtPhFuwDOU0FhV25
OxI/5Z0+Z+mC5ESKAiSaEhOt5nd/A2RzcnS8NjieU5vq8vrDCn+Hhmx33f9FyjN8
D5aDI55go9I1uwgI4Qkep+h716ROX11U4qWFYydgIFrhwCInM2HlnmSicQWJFyBB
JIGHAgoGzkBvY0f4CzWW4OPtEJHiFJr9XUXisBTMk62+CWOf2ov8AQD+Anuu/5mY
ai1fXITL4zfLmkvQKS5x9zFECnDvgDRBkl+7Yj+jKE+T1G+QfxwUAhzrbuJ+pMkD
sgg4SXUoQbYQLKt1UthLMtQraExkRt/rG/6NtP0m7o5bNXIHc1Aj/fiDwnBub3ij
I5IyvZYSzofr1fukDPLlW3BqXkZSlfkxhmCrg+XqN2HoOTWpBN2G4zhxLjh3U/jC
Tb185MLSQQNdc9qJXoP2UFhIHHm6DwOj+Q4wFO4Fm2UFBlxCjhHSU9khkf3StiMh
K/d8bliAWfdQdI2iEx8vJk4AUYpGcuWo8UJcO9jbQakvulGOGeQfbzb9iEpSbul7
71wDDjh+EXcdr6C77tRsZh7Dpl6oiqplmnFfhv576dL+nV/b90J7Yhn0MbHXR84u
Qj3yC4H3wIJ6Gc4ZEkDao4pwjqliyCPCNr6OzB7tBir1gxn49g+XplZ0CafxGM8d
ubJY/xfFGMoo2gokjYlzTR0t9n+cooohtvSJ4acOI+cXYYr2D0BeUIreUAI8NUNO
cUsEjCT2ePVv8uSP1DGfRUM6cmXK8s5Es4hB/CcdqJWx0Frd7G6OKQ50JVzOoiFE
2hCNrqpcAH9n53YA0mzEfSmlsTSQHkn/ja++sRLseWn5W5l8xmf3otxXjfeoqxvx
qLys1/C9rqpg83rv2sn/pVCwG8iDDReug+TuKMqEtts=
`protect END_PROTECTED
