`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nJpO2G/lB/nhrD2AXii3emAWw1vs3f0V9no5LFKtxdhfWB6CEH8KmIunEqTqtU2U
nrB302uxdKQfbiRTnpXppkgzpoqluo8mRs5I/J0Otp2ePBFAKdoGiZzKvqq8yeMJ
nkyzpsTZnh6vEDyojH7tCraaXf8CLc+j00jWJRFundFGGAaV3jpw6Dtzb7pu0sX9
AR8YI0UpIxEmPRg0kFVOezzYJjj/M5I2zi8beZeFAHu1m9YEGGCvTO76fRIkWELK
sk0ihzZDz+qZ+nruYSBJRtNeLtr585fjvzA1cL5WD9jYcOG0cDBUvC+i7Rs8QC2R
0tlMwiz99rIhJ9glQYG+AALxeqio6WKLCL9JpZElbJ2SDFHbckG7MHmfGt2hGv/t
+osoVDdrPRbA5mvcgSHiIggLccLja8Dbrkfkp/J1e+kiMgaSMFIbZa31gzo1TspW
vKooyPyP7+q5pzVlUQW0j6+vubmUxZxxG33BNdqSJ1PQZ0BwFLDdIZnoD2L3emRZ
+qZX00TKrEyqdHz0By1gxJjhdkdY2vHGqwSkkJ3LOM1VXZDfaRUSdxItqCJckHZu
ZITRXT2WBVTURMxVOLr/Iz+0kCWbwMO+bpiRG7FLd0eLbPkVgPRYWCbbAD/6G617
pePv4FW/Iv+9XfjzXbN/HzHDYLDjRRJS0I48UGxSIcc8LYz3ZNEpCG7mkm95+zB4
vdzf5L8BNUMzaMOnPkmK2aMrGVHuy4zQ20SS4BWfy8TM4nvt6GOgUjfzreyK4j/H
ir6ATG+3rCD2oKvweAhI5Z1VnKYRipQvQd0YQxbFuCQcrZP4IAdJNJdMDTEjPLAB
cRP0pV5WmGI5hp4VcZBhJg==
`protect END_PROTECTED
