`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OnlzwPWL/MriJ3uIiYhXAlhhiiiuq9pBuYurCoPOUtn9tI5TprKPibgpfzy4ST7F
KtgylwBNlUN0yJEljmJhIFqo+DXu3KGpyOhAP0QLrZ7y4EEmSUu7OLOmxD0Yxm4l
bvQu8UH5NOa/fEa6HcLV4zXAASStvmSEzTQjYQ7K+8DmjKNRquyI53TSYCCNbaco
9aN+zd2Zg0wnf6fMnOruzXr38LjXPOu3a0o/irpwVhqYdVt5LCaadnmnwo0Qdm+R
njI/OOXxk3XHJSKSPPORHAjei1DGYj4XsquyaPRr0cI30h5o6p2eiV/6VA8hBkr4
0nGy/jqsV5ZFt0AF8sFvIl+eHgW1JuwWgcd/YAtXaKybTg+Aw3NrEc1x5pIDTrvc
XzY0izS62IkpyPR687YNNJC0uv3HrYvUBv3/cVWZVCPI/3BqAEidUqEvjxHpFMbc
KAa8CyL10+G0eMIICXVtEqNMuysoUXA5pfG26mFwrGY3wNwS/iDsLzGSAOrx68Fe
aWNH0+eEMbFofXkYQn8L9yOis7O9cOZSQKCcot7spYC1PR/2Kul65ta7vi3y8OFN
LMjpoVe95nkdY++yo667v5vCr+ofM3zkuQ9aPYtHtNL9PiMPWhQGqZ/eEJ0Fv6rc
U4ncmXT732wb2/o8APhjlklXIOWF1rgfsoJ0MYDjZjsAyXeYu0lH0G4iK6Znorwi
ikPVtjDmtOTVP3TAMxObNrodaVNTsG7NRk9nofFABQZHHhf7bynTtdg1RBnhniMI
kN+9stALD2PZ/Pw++MM6bRoGsejXExIGc0Spaho8H2ZszCx0nV+CehzDUKih5iHm
wQyKCaXHqGfaRKH9L1rqpUV3fkveXuDTyBL7M1eqSi4zdIRu9fnod3JbxS7Df+D5
XpA367uS6b9F4G5i+bea3uKLfTtjhIfiYP9HPkXn04jkQ5Dv83rlvUxszslNNL89
pSr0Ps506C/wOGbVT02Kz4dYVn1At+PQrXRi/RLIHB1ciJCA/s5+DeYxrv3MtLrM
RCQQA+pMPmgDX6bVMIl1TqTOFf+ALdIp3V+WAgGqKkvRPvRqsmb45ObwabwVHLGb
4vn9droKGV4H/vSPW0UP2wKVm8rNJuKudL2nNZiMa+CT6Z7SwWK+5zXZAwzlrYFh
w2g+IthKWqXP9cVLG3poofHRs+kyOU6CPRtBQOmlzUvVh+jcxI7Yei33Om8RszJs
kQvRgJiiZD/SQdwJ/rfoZ4/cAk7sfz2qPKXwcienhSoOv0eHU8Bkp+ERwGH/Uokk
Prbq5/s+dj5Bk9Veik9xGRF5vH9DKxFN75QahQa5bSsjtxkKaqmupzX7MIGSGZxY
EVxDUwRhBl4w4VaEZdbZNUMBvoz5UjixrBkQfzBaj+0WkPZyM9LQ3y3WZGRHMQLA
M5Z3sPbS2mE+lLZSEdLHUn8ZwkwCRwfpZDeyU81vGHQ5JaC5mqIitIFWxCPhjm2x
5ArAh0cTL5OxmHXSS5HYGxgug18Pty3iv2loIhYRJT5FthZFg1q3xX3YeYMIz2xY
p/HW3GBUEyK9ifDv3WzZGcczwVt1Fet0nEiG332JvWc9VibmD9pgpuNGm2qmc609
9LRGHDDhp82oCR8QxFxNvZBGgD2JVcReZuvCzuS541fWbn1gMV4fcmpsClXhFQea
q0SZHjPsvvKgNP21X2IjgaJMioXMBkFPP2o7VdFW8NWkscUUiQdGwW5u77tQax1h
xXDzAmKDpctWJQfs09HbsCAtg2sy4kC2fh0dKv3tQ+aYEuX+wx4xoZUcywrJX7hL
`protect END_PROTECTED
