`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
51xNB5HUxTRU9n4Rx2ZGHYGIyw2xOO/yVDqdtYg42/+JW5fa++ebUX3unUbH3BZ5
Hg5IbNisPwDczdoiMm0U6PVXAuf4SKzdrN3fCOCYIG3dDsoODIRAjlSZ3DGKRehf
0LwXfJpHUVKZTSbdpql+g6IFk00TgPGiavaSJNqTuec/IPD3WgJNzFRwpRtjq07W
nk2/pwvWkNin1s35s68KlPijbwRRrGac24uFCJG//M5KmQVvJf+BY4phixcmhESC
vmxtqqaIIqQ65/8aTYh3A8DjCit3nhKfWHUsKKl/JlBxpblubRCActWBrrSYW1XZ
+wIDTkvn4GcpcF0l0W9QlcOcVGywYquZjtAvkjtd0hv4p8rLNDh8D7HDI2Ko3K4Q
GQvqhhv7feAsWNeJE+dwh0R4P8Z5lV0r9iNoRQW2tw29OQZu4YPr5C67bfFnDhUL
TWpkqIu9qz1W6bpn+PtLn+8FYbZY87RPCFOn0H3ieP5XdXrhhl3EqgqoVxyv/4w5
9jc601vnJFdD8xtwfuewVvCPItSqr7ruMxOBRNpnS178WZqxHctFxOmBsBM+OUeU
4XxMXV/eNaGpNY2hgR+7yWYoUQyny7aOaBFn0grb7fXD9BlECPioCXQG8+rrsad+
MW/Owk4rvdj+6wjdgbrgcaiGAo4fJYpkzw9OoNHaWdLuBLmOsFnA9824c9wten4Q
i+hWORyCz1Jhb3Cusp7rNXqgvvaIpAPMWr/ve/NyQSRA3fl6dYP237u/8mZwDPTI
tG0Zo7EN0pgrwljB2hWhz3prJz6RIHBZqfGdivN1cbX/BeUv4NqFZcmsELROGIMy
VbOgRJrImQtteJ00zNUgaCk+3vP1m7j/wggRIPJym3atCe6TkpRkOiE6O54KCRzz
9EhSrfWtpfFUMPvbyNxhROUwYXwlJc4Va3hCzeooQc8173KXywBvugjRd6UJhAnZ
AF0UoHQV5q4DHUrx0wNJ22dqi0fqqEvPC7/FRuGVeOr+kg/3KgFYE/GaKexxmDpE
ItIlqebOPHfpgZBsDwTHlq08Iw3iGOh0gOiIosGyGga4PwlH+t+n6YeCs/4Rxbeg
ZmWpkSEExdHX+AIc90IY+NUFnDbjOVtJWbkb+NTzA25s76hSspyrvywNYy7waMQZ
4n0lc/ktWTF6DTHCG4cipArRlkqdjYU9jkrFKCaD3Sh73Mn8lOQW9kBkZ4MLNFpe
T3w3Lai0Lgrc/EYRq+mKmKAOdJiYOxEu/oGftr3IlxIlif+0bdhkh2RCBpqNItRn
0laP9tjv0Ri0/Y2CUUmasmmH0C9zQQ5TfTh39CXxJjE=
`protect END_PROTECTED
