`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BNqEYBJTwQMkD+/g8AhvFPbJ/7GwYbY/DbCVmY+sahQM+LZ3QKOlIQ/5CG+gdifS
POwV9T29dZKLpI6eS4fHhEIISracpFXGKz/ssbfyIFQwVF9OHg4wmPSW4rqx8uL6
EAmDjV5XpxVKCE86tcrTd3jPpMCIoQYNVPbvBDrpzfxnKlpN5Mqv3zNgvbkAgDiH
DVrsAnty215osjV6bno6nbMP8MZQqWx401G1bkEiRC66EXQlbinyuSuF3n7hWEQI
9Lwp0obgZHF0KdfTlaz6aZeO7Hy4fvt4ycCV1LXqC85Nk044cSheaP0UgEX+wzdU
oPJfXwDmycm/A9WXO5ZMHWfRMBYl58532xE/hSYB3ZlbLI7TlU/MrNYZJr16Vc0b
khhPQAm8/NSkgOP7UJcxZxVJBdjP+KolIjnPwRAwv49p/IosG6NPY0E5W2caPzeF
lHpHqDTiy0qAz7cAQ+qkps+dB1hz/hNYa95vbPi85CfL5qnj29CbkGAGVRuMQMg2
e2KQn1n3UAvb2qhsY37NierwbMPHdjVdrRKf853zx9lEENokwUwqW3zPCcaVl5B7
0vhgp4GZwrBC9fCMou1ThCIpX5vf7Cvz/PupKJOf5vFQXThr1eDjmPHYoqJ11IMJ
BuTMWFhFDVhgNkkLusSpI2OggbkICfd4UWzgLyX1+fKF6t955nkrQwZwAUqU3Xel
TLDUkIqQCvGmGFeOND14y7MPd4JLMX5rs4+VgUMOo/ZtVCZhoKYfgFKnUYRH1Sxc
Ozk1bLIe4BuZGmQJT9fEVMjqateMoMzW/3BhUJb+EdTV1WNnyJ8aH546RhYyMC7X
8RQnONCVy0adINXeSsV/3lgkiKzA19KQlgNDbiyX58i8yvPE9qee50T/XOsnILyF
P+VzWBGfcwEGFkG+7nwmJmil6Yrrrlb+zym/KbB1fNemfzJaKCJ/t2Wmvm13ebd6
gyWQWhDhV9XfY2HUG2qGpM9cGR/JfukRFMT7NtUFs4iWqigjI4H2zlbaWglMDPjo
dABo9D1ZKFZoom0XHrCCzosXMPEpmEjAU3lfJVXCaKpSJ0DefD17Y1UR6BJAcWzl
kamq4J9kbIoSF2mpwtSdnu3DwbOvGtxr+LS0TVmQjqCLnO4EfKveln8a8lH4HYBk
W6Lg/bZPfKdSmRt1l9UOIh733JGujj9QDTMm/v3+mcZ34xkeqqCLYpuEaX70mcac
KfA9o4ynGbXaGeX1Ci70l8FYGQgurIcXSBYTDh2Urt6GbdjsxINmzbbmBB3A2x5n
ndvFJlAROWV1NQZhTXjoHTaEsMN1NRfzG6wlFxUkxhceSEb/jeYkKtFUEvgLhepo
TFViqEs4MNB2LzXRdATzdDJ1cbXaH9o0mgUcs6bQcTuYVgSy2NWjiAwj2OGZ+rqo
+x40WNW1opYzudnGuuw0hSMgoNbtBD2WhnlTwOXbYESeWENXDe9/o5hoDcW76ZKM
1OnA+PrVoaym6Hiv/Ap8xrj5+CyFv+uoRe681RRzqxSoHXPyxC7cP4PZO/FtliZ2
2MuCrMRSOvk1u4NVZW1U9NuM5r2c6Ix654f6/85v9SISBKDDf9agljfBmeqDGu3q
2NOC5cQfqN7opA8hc5LzxQuiv6R/9IG8E3XzGQ9Ws9w+ojQupJEcz2gwhsmp59oj
Il4tmMrg4hYtcGN/tAT6KZw5mht43y7O5ULeUzuUcAupGe1t+d5YjNCPjAE3pYQ+
3hc0SEErFtFw6hcYJsPCD7JgaR5B1Gf1+cNJpwVYYK+PeCpyL5xhOlM6rio7794H
SZCrnvyciTdqs12/SBqL/hrZIHRyD+OA1irCXU3S8p9qIKPpjRfp4YjMg+q0+MLf
MG8l56/ux2e0A17bNzGwGQZA6yDEjMyfM2Prz0l548lL+mGg6mVLkNINaIPX3hwX
jNS6EF8RlCQ/yfbSOKxoKg/XfKGNVWRVJ9x3uEuvKBwPxlFVmFt+Tn54PoN3of0q
Jitkv6KDHUHhVZf2EbHpkSt3qlpFl8Hsw7xqIVF2I/ot/kstRmXXc+XCDi6JcoJ6
Td5cJ7GXxbCSd76aV7z6J0g17SafGszISuH8W+NKXdO1p02MeOugUsKWAH3PN2ns
kNI8VGhxzs+WdWY+H/GraUYg9r7dxXH+2FZWcs9j5dqtkoUkAkAypnId1eS+Oyl6
4PR8SbyF3jfK+YgFdOOtdfSwldRV5iPdifOhT5uwKoLrRr8344VS+Kv2PFW/i80c
eDzwh0Xe12URaSFeXWKVpQZNThoMmh/st7YLniTopVX+iPKxi4roJfga0PulWKwv
qqVNSpfWLMR7OnMt/8xL7dmi/JDLDRM24LZUpp8D+ry2zPGyc+GmQP5CVlJJ9wMh
ACX/u2f/jj58PfCy206np9pLitrv8JSXCXZiiFhA3UG+cwT+w2uxK4NDEmtUtfLk
y7BGdchk2MXa7s1d53n7nWiE3jqshMI3iGvX2JYjKuUPyr7fYc90Dud5xvciE3d3
aXYeaafIIf5DA97QtCJUUXLwf8ObLIKaJYvlPzhEy7R4jQWYWATjaFy4L6PvBTLg
SCTOJaMvnJLaBo9f/Jm4Xq51vwLDh9sfk8wfxuQa5rc/dLUTxgK5RBaBR4XRoi8r
LEPZ0CV1XXae+MebhdL2vH7SCDXYB4BMn+KGFVJ195I6mau68bACVouUZfwWAVK8
pOcd4BGp+Yg0wYsc2EN62XhVaxrtsva1IqL9xZvAkUSv/FsV5agtMj4FzWBHVDiE
10aIrl01cMc/N2LTCfCWc1Am5dW4yA5EFgCSaz/tc85DoUs6XXXxDGhCaOMdneHn
dtsvU+pTnfVaMWbO/HNEm22OqWX5xtORmTY3zTuTD43IW5XFUrpnyC9jEovBuLM7
6UQv2P77/sNMKta+Y5UD8XHWUwQ5SETvwimlbP87mTib6su6gFgbrtDadhzBv81i
h7YDRvejYhPqjkl50HWrUMhT8VCRYMI/M1+Vj7nVDyRobpXRgZ7h+vFyWLypHgTX
LXnX862qBQYBaqSuuk9w8HvplMDvDlU1fd5FqQHVb47RR5dqf5NExziqdtVtIp+a
O/+bs2/5KJQN1heWyFWkuJ/TvXn2+ElSG78XAGt7lHsH78G8vomTNUvnhFHH3oWP
8eflOiYxtpnXLk3kMpC0/P5/Z+UalxvUTuk4GNYJ2JXyLZAS5QKY7lYa4F3rbEat
keD682DXjt44/TBd8FYXeKHy8+jCQF4vrr4lGdUyVvF/HXnyWfQ1jtanN9QJfJ4d
VZMnLL5OowpyfTPEW1K/k0w4ZZlfA5rlSfFnINoEu4nqd000LOPCduz2ZmJ+bIdi
Bg1I+ZjunfoZTls7c1lelLEYXZNobi5unIOcIrWiqxA8OZvKycZxyeAyh3WLPR8f
+qL6+iV0Ns2moPeUuf4mFvK6sFph/T/OXNoHYL+3OmxvjMGg7n+HRXmml/q9Itaa
s8N13FwVEu6KzPuxjVOphEmeOAGXF1gCkDoKpyRV5x0q3J29SxT886avd1hFbB4D
/PlqFcX5iV1wGeQImnLtOKU+bUYJh9o5aAFTqhznLYCuYyh0/wQKJFldNI8bRxwf
GEwYXIoQWBXeIDDoImsd8tEXES0Va/+p/McqSPwyveGmjCAPEVACoyzvFaGEeZet
HNt+AI2O611thKk4OfxPURkEz6ozj5q60x+RZM3GHk/k2CrQBas21mCWfEsei/Qd
WFTUgn8lVGQBsJvGaxCZ5snDsjxWqSuDJv7uSWCZY1oexGogQbL1UuQkl+5rMmlw
xQhgqX0zalSOYPXuAh6uVgbxkm0mepxPCkgTBFDDkNz0/OmY6Jv9e7uxWaEPrROM
oeGtDG16s5YqZ7pNJeUjWBWrMFgw693dWhYgvu8zRcbbeH7ONLrBJbtbwkIshtXh
x791ShY1UV/riLv4Chlg5YA1joCrWFohu3xvF45PbcbKXHVT0o/xuC8sfpYN5K6U
ccr5HYCapw1pll6JzhLbeCAIMLqR2k/lyOXHBa4oPTd+Xe4F3VMNp7T6ZbqmGmFN
JhCyY7625HZ5TJabj/wb4BRNP127KHDs8bEOMtgpa6FTtx2uNWpQLqWOcBuphKbQ
20/eAbg5Es6qELn4eZFJmVgUAvT4uus4CGytLhDBnUzAF1NQVe15kTqlrkbjSPHi
Vvwd8rPG2yk4ykP0oTqmSUekqVjiN5FNpnW3kEjiRmkYjzERWXJEw8K4LZmdqjPf
jdS3HkPdb8rAGvDb2buX5nGisxp4fS8QealcSMWNbN/s6HT5+sNBPZoYiGONvTA0
pMAXKD0R8HD3L79J7TYIIfEVGvdA6FHGOxYPoOVzaKYZphWJS4im3fA5fqYW746/
sPhWpcSEy/D8ivdUfgx+lIia9xZq/ttQBkJ5hN1v0VwcQ/GbhIxoslKTGBTF6cNm
flaE/3lMPyix2nqWgKzcSQhiXuYNm5cOKiNHrusTx+NVtYauhbFQg7mIhq2QNBNf
jNWjJtu8JoE2GR/0w9q3Q26jtFHgvipRJ4zRh5oxCUJSijJCHs5b4tmULLFTFZE0
aLBoa/TTJ1KncMtkNnCn+SI887CScP9Pi83tl5SaVTCF8JvCZjzmTJ2csyDNHr9v
m6/bp8pp32FDA7g7sKJXSeUXNGmjHmKJnOw/kwFAlLw3fIQ/3oOFsCMvY9auWp+E
apOr+78Pbxs6977uZhdf7WgGOK1Ef/NxUjWtrlJYNeTDsD2CrU/PSKczP4TyTmUu
W0WUnOL7XjZxm9rznhX1UIdGBrP1wVkduiFzYULxvI0j+8u43ysTwW+L8sWyw/nX
F1YgnVUHzEXILAM5sxTvNVM9zFtK4+dKGWTHGZYJ8Nvx1jQc1MdLIRsJCsibEAev
XVlirlj/D4+HEEttixQluWYVr3CPGhJnsE86x/+jviUPxMH+jT937/Q/WaLlFCBK
2H5HNC/MPD6OXQIPRZZlm4E/XB5mqoyuu6nngZTzgFCQ+kmCxjlG/o9nZNPYpyrg
126DzP4NKLQLTMD3Q/Xc9P9hLwfiWQdZz7MgOqvMwBxBRSkc5gzt4sMSVGj0SOr9
PSotramVgJrC05e5yQvxIkzMuQxU4OOqTSw7mQ3osvtfokQXDCGjpDUQTsf/ey5o
9/TcSlqIpdFU80sA6IY0j+wWhcyea0Sr5sqNdSJiuApyIXkQL2Rio9RxIKxpoWj0
`protect END_PROTECTED
