`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+oLdS8UQd7o9bOdaqczd4RGSG5Gf2Doh5xeQOyZHxZImhi+49rzgMffIjcQFrOgf
eWRfi3ZXIbACSOS+TO87P4Ok+gRGd87djPj5L+PpkF/Jmkl5MnALYVyy1XvHtaJa
vIUouty3wgwzSBX/U3XoAS2bkbCVRUIEwUjd5yCzI6npREBjq9C872N9nf3ILNK6
tvZQeF1jQNQBBn/s5kb5pKaiYrqPzRAcVlO6zyxFPZasEHDUoTi2FxfYM89nb/Q9
hbyjyTIBF6ewarFFX43p+11xLxR+9Qkn1WAOrK0kVOpJ0s3Y2WhGoczQEr9tILrH
6kon1OpIZ3JGNkttczqNeCtfYzPS8R1odlDlzP8WRJmw6b9EWSGjeXRfdU+vSKgf
1KoLFM7QonSYch5scIXGAfNQ6wqXGR+W8WQWy/gKNOEzoWZJ2iBBFWhDoytHJ/d+
KN+CDE8Bq62e4TgJccObC//rvWPGMF9za8bcVBq790k=
`protect END_PROTECTED
