`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OfOGx76VO4FGdPNPcqLVZxk+NaB6YD2mqFCzVBPlxzDQumFAIuJB1nNtlrsaGOgS
trv7XJgXkjkiei67qTi3NuDPYxez0swBWbhgHXhyROFa8g//YL5PI7oajQvVR7p0
VtFTYS13gAQXFnA5zLJXj2Zo3aoXWcj/V7S+pz8nQST+Ox3G7JWZ7QawYaaSSr80
1aL3HdlMQ0Sg4YWBocZi/RmgqqUsVKzSf1ifBOW7lO1PJF5xD4QcHx5sE6+soh+8
GD0j6ra7CEwjdqanhVtNhiEIRpAUZw2gDeXyT5PEI4K4P4jVHV2NCcDRhZpBygOm
/K3VdyKkZE6JMGlpIDj4nbimynfd198eXCd7e5UPrn3BzCQ2xetP83DBSmf+rHl5
uP42tJuGu8i4a5wZEfLuW2L4LqFrjlvD9xuWYucp0OGHavS25LDymKI3O0tpNAd3
JwRrIUE9aZUf134ny85QJ6eze7wLoaK/DZyFynhaRjBw1irleUPCop3KqGoRFFj5
Mcobp5ztoeF8RSFdtrG6FcIe7VIxq6P2/bK326LsVQwCnX9ghouWk0Znt13JXunY
jjrd3WwhrPlHkaSskkU0Npk0znKpca01ps04xskcmHtET1Bc5wQ7KsoQ4YMQ5Scq
wds9mOMZ9CaitWsX4ikSaikJdNlCuiARjqltA+vx/TuaJkc8f14CP0eIUOcOqgcZ
fC40xLwtWqu0OfZKODlGRo6mzp7NvFiGGhql+uE4+LWAA0YEccCJ6F1X2MwFV0J+
PtufHjbFZMWshDNhgMAtMY5ST0s7+DbDuetgZRD+KJuuD3FM/DoaghzgJkBpiBM9
5ljdFcVkgcA+WThjB9ELVcSY/cBOVFBIhfHlJPsm28Y0M9DXuzze8rG7Dgf0C+xX
0SwztvneFNAD5lgw0QODy4YV77Z97HOOXi48O4bRd65o7NdX7XLJni3qdBpzCb4C
s78B7lyT3/AAdDxnaERZXrwUTQw7d6xkcL45QtH+13NmuS0LEjO4IboYNNzLmMSq
`protect END_PROTECTED
