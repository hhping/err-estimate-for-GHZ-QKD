`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lt8kDKvZOpfq+4sRvjJpkFIaGydM42ZVD0bS9SeJ0masNkKzeEls5lysg7LJ9/J+
OmM3TuQkjoqEXrD7HY0FkecxNufIe5wlq7QJCXFIjsZstRjJf14/F4WLTsQDciRb
sxzgG8uR6MahwePQlk+mvvcw91yxLwT+EQ3kjGKPoYcUn0b/qFXD3+OaCyGwPbDL
aLZIYAL6rsXydMAUymgr29LoDUSIOJ0WCjCKCtI4pxf22V/UPuC6wahKeCQgPI9d
HVsdK2mPjjQtRG/x8ByDRfa03NkrZpeGlz7EyM580Ne5SgJ8vb86YKPH/hX4jviQ
P+wCIHkJF8VUJqLNj9Kv3OXkTdvX8L1nwS52HicDNRMbY7RAPWGfjbGvExJRuIyZ
zcAL04GcRPk6CwuczLYjQwyNmR2bSzhnV3wT4/ILl1WrQyP4FsWPJESK7D4M2GH+
GaptbRiu0xUVN03LNK3srRCI0M77ujZNxY4Hx0/EnN/omyjwo/IlQEjTe3MyEuc0
FQ7MZTNoIuvXemmaRSVER03socpiBy4fYxKAEq/hWqzKHeB9pMJ/NaKjqVXdU6tQ
EMxs2KMZdRo3P+g9vPdyFjcO3Zl8aumrioaDSWS2m4448RtxhcQbbBH2XAPeR+RD
2vPZ3BaGCNFZaC8FJyzAUZeI/vy/8pv3x/fpsAbOk6zyBq5wdKRJqqOSdqjOZw52
HSsmYQBYXq8mtisjhBSLxXUsMBNHdRBZG8l6aS1N64SfS/ydjVY4wqFN//ttclSs
WV34vPB9OkbqlmVgODKZKNKwf+CvdDsJfA24PHPY4JbbSPZDUHJtFP/wkbHcfoE0
J1oy6q2Q/M/r7rrojfrOuFWkbbFjw+54ObekyGf92qhfk/6LlANAwe16LqtAKQtq
4Hraro2WXSKffemmLoY6f6gQov2EFLP7tQUKexLzrlLnmcrYCcf1C0H1N/PrMlEW
ZmWDxLsv8iQ1gMOBdIarNw==
`protect END_PROTECTED
