`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D7HgGcooN9W8WaSLmA5z0G88KWPJEMrn0y46mPPUq2GloqSjz2c9GFM96Z/u65kB
9cIqbQShM3Tp3qVVJtak827r3vRNlTFJtVJkbfn+Ol5o3qKDHqTTQ6RCdP3RUt7M
rswb5nt9oOCvqL9Rl6Wgvb0RPYx/aFXTqfLCF8OVbk3f/wXwck6n+uYk4mCzJUAb
qoNCLPYT1HHt8MDUGU8UB3z4te51NLDR0SQL1g43uobnXIfTdPLD4fBvJKTd6a9k
DdsN6VGeX3YU7tu7jrQtznwVqX6Rf9J0qg5GYLfZ5SUVP2HKnfu9F0oVMlWpeYoH
XGafD56IZrEHatbiJStAqZgAvgDW6eDoQyjCeeWZdH6AQAv/SQ2zyGqflmVg5plM
cmo/L/GOyRP15pvVmoG5JSS04rqT1YVIQrzS/PD7G/j25fufwhnviwsqdYvIIU++
4QWmbNYWVrgGuNDNwnRVzfTCC5OyVF8Nnb1HUjtkyKGjHeE9nK4VdAGl6EwMWEUk
PP3JxJ8gyusF7bVV9eH2PZ8zJGoXf+eGcwDNRy6RKCydVpFFChLJAPM3mGhNnr3w
X191S2XfwUcAPVbXQaLLzpja7ZTnNF19kiJtGMzWujOGKLfiQmQIb+FIzYw3FkSF
1YpATbHkYZERkJBNaARob1bxOaNtywyLIW4LWMlQhyUPCa4qnlYvyS5LtoDf8v/e
aI+bYAPfRhNTZ7+rjtLuxwwSewnQrZWOGRPEjEYFZsWwUSR0W3mP6qRP0Iiqr8sF
vS/YnZJtHR66k8Mm7JziaIRbDuAjaueJQ+Pv4x7Yx1MZlXQNYx2c5aiylAmm/uBo
xQVCAYiEhwA6f1voPuX8FKDu+Fj98K2rYEAJ/x6XEsoMbluDukBD1JzJQxQ8C1l9
3ENMHLOhYkvCBvb6/ZFJuZ3rK29csbrH6Bm6tTYt86j/lMzIlU746k2iFrQ/FgwZ
ws+6c9gu7zF0XwmqS9ntknj3DMlqw2BQk74AIKMB/oyhgOMA0/cnfYgqwWNvfXD3
a+u2I+DW8RpaXC1Z6LwgCH/wYFbkmL6U1f/sVZBYcjVdkSeNLL6AKLsnZnXiWv1d
uDZhgUDy1BA2r8X3mfzHxqUJKMBqqkj8K4kChYliFm8g4x+B3LSMBh+dR0FHAEJT
0YXcTISZJiOF2fKTEiTiJsXb6Td02lUqgJ88Iq0sV6VJ84RJk0GXPIwx6jsh8F/6
Y82VyeV8KT/GXgw+fl6hfMFOOFlSMHsbvPGDlnqZ1+aBZO+3Kj9s5pdDuH+ynWt7
0RORSo6+S8bU6VLjs1/fl/G7f84FM/zEzR1szuKlHizbv00m4JyoryYam6WXPA5i
P+1vstEXmMBto2Bhox4rAeERpF6r2zbk8QoPle6YlGtdU8v7/hAD5ZysSinsQ25H
mkALkjchP20sr11t0Iif5KXpRUyDkQllx5t+mDU2rZ33/LE48iO/on1KOjoTDJ7d
Aen3Yyf931mXKQHdaf4RAM+C0hFPwa96nhlJ7/+Kb7IpqrmlYi0tPWaTN5aN+nLQ
+sJVU3u81EMvK8rNdfoFUSAtyU5b0zb3aR7hI0GicajaweZYgwPPvUeFQbaRLTgy
BwJaU81ssk5zyJvWhreDYi8dhuC07/5WSh+1qJIEaF0yrNpRgjmtpRd6suK66o4B
6whuG2ydHYJe1Y/zgm3w+n2O4Aq0HBAI/1gClGPjpN7tFLUsPCPGu7F/GYB9MMKb
s3jygFR7YBkA2f/FvXR8XUTrL8SabqKhiZRaW0lZoajTAVCsD3PJQ8LMxUVoWk2Z
Zx4tuDXIlB6pF1YWgzHzHajhJ0T00GPgWedVt79g8TlbI7r99UxW4+PSGvRkqJP8
wI0ao1UGamrqmJX0wZGVEicuyJi4V5WDC8RC0zwZfRDDMIcMSts4eKrUPaNd+MTn
X0kHWoe69k6xX9LTPmruwvpWaaLttuJK6g+SDPTnfqzh/Do/xiA9/5jrUXL37pod
tfpQIDRVfLgjH2xnMh1KmI0VLfNgX/4EcT9KYqDTtzqn1lAwDRg/Px2IjMYHShlW
aPBb1VdDOpPMT+ChkGIjWCzGlVhe5ODYbCw0M0cRYV5O8rFLBgCekBpK7A7DxDdD
TDxJXdjI/U+xpDIXi1tZI9bqlAYMAsmT2gawUcNLP1v/9ZT/w06fXH76QNxa7o9B
pVi+eytEM5g7lWYInhGizr6XGxUGC/98A+oLTioFTSB876YnPvUkofktGuiTEBvL
6CWTpwxgW+4fs7mJPaEThISzqcsFjx4GGWOjTYRA3bfbu0h82saDy48HgLKnpRyp
l8z0dZ8zI9tSOJ1bAZlVzsGQ7Pr+DVrByNVnmsM4UGhKDfqq3XxvtBKMOgGXnyJw
SGT3giBqyvkCA77O9SA4ZxsCegdSAFJNTJQbS+R1tfAUQYAeTMLpTdAciCkWB6Ei
WLJlJArg3rb47aJ615d62JBsSftsXH6hbtvfT3yDaYnIjRO85xv/JLcCzESCpXYr
rWnEQ5u8sCTFV3t4WySe1Y6PFDpX1vLOa0StMY2STOkE3drksF2Skx+dDa+04qhd
zbxSLTJVu2CUn/f550+GYbEDvEwCahwmxvwdwNFb/OQgUaJoktlS8+WslcRT0Ee+
cqrNVUzKItOAF2zc8UxePGkZPMvFYF/NZBXLmWJTmMfc/RNqanm6vcHdRYqLSJBY
AmJeyEWXBXRMaOm+TYWb+3uiedsiEeTTu6JIBsEB0cPLU30SBX4XiYxCkwcnxkfE
5ZVCSWIAwZIZkSYZZlKKyRbodoNzFsF5CVtR/dWPCjwvDgMuvQ2MCJA4bgetu3oh
YwTvFYB9Rh2YrbaNAkKALzuC3M/qwD6vr96orq2aefP5uuxHZZzIPxmw8NAyJj3F
+aga/UrOfBa92M7qxGW8qYclXOzCQ6cuI4RuH/VmT846aDjq1mnyA1f0o7WPDANS
qUB99+s6XevA3ErwabN5ujzGW9+bPk/6DKzyieAEQ5oSx4qY7rCQ+MCslWPM9+PT
MKieZBrhgCccppX22e7wCTju3mQDXMxy+IQGKa+BcjraLmpWv3rmDyK7ofDj7TAu
WbXnJz2kldaHPVCbls0nQoLAlDNkwBEgLrfhIKp+gnMshx6gTCQwx+pgYM01t+3x
t1opRE/H9ykFTFj4TwRTcXqSHlAlhkULXy4yRgRkApoCj5PnhSAw3etTDJkzYfby
xFhDv5Fa23414MCa9H3ZL71bs9fw6aelhJjtYEKee99tDyVLNJHMhCsuJtaJBmZ5
9BTIdTjfRupDB47FVyzJ5PRTnbxbb8v+9IXCbwBC5aC3wLD4d5iWU+nypx+z1GZ7
+ROcyI6yaKUzpEYWyCETqO9QHDg5ROPyKov8Sw93SefLxYGBVt8ETnJd6HQGoyo8
VszZtpnVK1hAlwwH25XuUg==
`protect END_PROTECTED
