`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a3/jU5u0OV5jtLNu5myovtFXh0y5ZzbJGOtgXRKws5+gtUEtcpDoRXiUmzDkd6Dx
MBkPPF7LMty9gGCrHRoxY/wVUF+d1oyHxMsHRnluUkN2EK3oDtTUYtcqc++F1aU7
VEDBUh9lGzoVohcQCNu8XISBjaoh168YFocQT4UO+i05kUfzMqp9m7XpgGSL+QZu
u2ZBnhDZyGBqJ1Yiwec8t5My4d4eq5NJmssR9xkHb21zAxwMdzjIP4MVgq/fd3gb
IifM0ZEX8zf8R4EG3/WsfiXWT16jGXtZoa4+vBooPsEuS94q2FN0h/q7H3ewHKYy
FUx0bJyV3URqMek4BxDzttXkkjl38CpBI2IALA6QOH5YH6DwUaad4htTie7kaeyb
ZlvHvwUZD17GUsd+fH9NwSKF51r+Si40fUFJdZeMUFs=
`protect END_PROTECTED
