`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qL0CIYPHSJANDQKouTg7+p0l6Pe/bHVOSlP8n7cLetalzXmNIXL0Z87HRrbiEzIq
yltc0Ybt1mx9PvqszVvhN3Ivc+/CKXPgN5qq4/K5Y3LTNXcaI2kBXb/xU2SadLS3
wUai8zbv9zQIcH5QPiEsCKTbcRzDQ6/zIfB/cCLD1OykXCaCn8Z4Xobqumrh5q/D
5q+wgrJSVSWDANGH/1ZrF9HI9YOBR7OCjx2I4rTbYxxJFCS4mDOSEu1SeBa8YXX0
n4/h6dZqCP1zBUt/iViqDwak2ymol9Gx1rjJ+O/qQ+1P6VknHjup2ttUEmDruWQ0
y0i1t5mPnFvdFYIxm1vKOgwpLZOmzVWlJapI1Ebgmc3/+ngu1an3LrapZfa8PldV
HIZNQ5X4nG7g7jhFWc8TpyPorLUDTqp8d5eUzO4caWthcOvfIW4TaeKJzIMcg4if
zlTtRuHIW85JgnWxxfQeK0wPYWgSXWl7ofbzqoEGNUdNeZHAPAMlMBiyuu6oIczQ
nJ5wnK088g+i6NfpQHlztgJ6e4wwEK7ArSHk+or1Vz/eh1pXwo+1s4ylgtMN6R9j
fhGBVoZPGB61zvum6GwLyf5Fq5bicmN0XPMlMKBhXEJltlAHxrn65F3SmkeYigyD
Hmy257h/8m4HEcMwBXLCPwi/r3SPwiNkuV+F9EcjlocTflAVyc2T2E142hXcyqI+
l7yHg8NjE9gwdH1naFNs19PCPDGiqvCLsqpbYaNZ34afrf4E2AC3icighQXbkZu/
5AbY+znxZiD/nnWrfvKclgpMHtFQkDG8L1oJu70lGw+6Ij3q9OYRk5AUeoOslZqI
55xjdcr5kI6kRcMiDjCYwu/XO2IAhcy+SsvFInsmuMZ0YPDsT+JzhGQSyioIM3gV
JhekT9gvRD7iGmORbKHZPQO4Btp8NOxSw8kKn86qd6dbkmdX4/Qwob9PYIEG6V0P
Yk5C52ZtCBBevwLLpOchAyySNfppnH0KRwBCzeqyk7RtVh68CztJLCw12wAfwCPY
+3xzV2RLf3OONRQvnwdpZkZfhVr5nyK4bWu1Oog5KibrX//eo2jAdMvNkA+UzXMy
GHH/vWcQ0VJGDj9yWaD7dM4wAR2FyL84LT8UuZCGeKN8w4C1KKjohLEHr8mNjHtV
tZeyu1iiPYRw/2F3KodMprBKcEurr1awMsVmanlJbz4Hg7S3Ujg2mfdQ4PVZwDfN
5yTkBUuJRwfQp3RV2cAcSJ/+n0YPgSz+26EJPprnXJf6ZFWf6nCU59p5EYHgeGDp
uh+8CBZ2N4shUUvHTkpygwNvcFiEBxNIu5mkBEaQ9mCE7wXWiW+siR3bitDgJcV8
P8ZeOoLtg0ULhY4MyOqSOdFpp0kuDu3Jlo3ovsfxWY9U1FgqGscd7PGfOJSpRPq+
ZaI3LOXYvk3bgL3rFMOuZsLYISXuIRAjdC6PgVIfB5hpjXpNUeZp+ckyMGVUczjv
Q+McuCanEy7BCXInj3YKhrlC9qDhh14t9TVTFytxW5M0mFpW8Y842LPig+yKxaXp
wqlVSlBkEGxIiHQeDPz1ObJgfcBmHR9WLRwMVws+b1B59zKTm0de3M688rpUQ+sC
Nto86HFna3dqfO7lyHMCqlqSFGi+nlMKN6C+5lR3QADNuLDuA8ujNlGhViCq2PVp
UAYMV6PDYS+HIBnzmDlWj9r2vDwCvGKVtMLAhReTLx3ygb5emBzCGNpQEbX9kn5t
2SlPkSLtkQk1zuO5iaOXgyo3Y4o6h/ZORO2s9SGiOuyrlyFjmWI7mQ46Twvc08cF
AKDbwKi9zEEg+jPqkR82lBZWxYeQDMVBmf1q22QDPKmWqy94vvRrMEb5NUn6YsBU
umffKR+0v4s3V7fvhCT9INTbwkk7Ln0ExH/IiOhBfTVXhxlqfkhl9pAq7sVwMv/U
spHjapSTGxh235qYwjXK/bPYXEA/UapCK4FXDJsuCE/LYTOv8w3lO1ppIIoQlaqw
sd9dvmMTY+AbBtIlNhZWokKa2scAI5IEjwiQnmLFrZguJIXsV/DBVyzVjt2aYH7K
DdyEZDozWlSZS7rfMivIgqdqZ1y5AE0w3LN+u5kLWd15+6e7Dd2WQj/m8lm2Ww2Q
YG9KCOPh+jWvUPZlMEVuLTnSxrGDfKXuYsyCet1ALQqfxIXvkuQl8ez5TIq4jC6E
groOXNyjkJ91w1Hj5xkyBfW+0ICeueD8tZzKIFeUejyblUFLHAQXO8S6Us1ilLtx
GntlhF7OuA7vQmtrsNXd5QyUOJhiwMC74cofA7/UCRLRYNfB6Hd8w6IXAZbO6J6V
/BuH1IusiJhEOPYkH2PSLw==
`protect END_PROTECTED
