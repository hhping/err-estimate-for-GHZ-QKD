`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E8inn6g0/Ah01fdKmdtUOYnUjsBosTmXnM1x8H2Hu6A4zQ0XdbMOhZ1osVLzVaJz
NUIesDtvwsC7eNFhBEzTn2zQR3I+TVnrnU2zVEqCK9OWcat+Je6v3TlA27gD67wp
l6aA4y/NEPbh28ha7VvQHa2VRiIpIBX1s6tJFTXooXJKl24pAIzRkTgxMNcwhzbU
2YWPNKimfRZ/jvxK3QseKN93iW0v69wCkl9x0KhOmlgY5oHlW8Upk9mkQl+99o3/
iNhZW76Q3LUIzIQWrT9tlIqcE3eEt1cX3Z22kfz+g9413m7QZdcvkAdEDhTm1MiQ
cz8Oc5TXCoo3LH3q5y+oAfL7OMdtuxyHlqXUiNbUus5XS5DMNq5GP9/PJ1O/eomC
scbLzxdwm1KywZ4kZ52Y0chWnokZPmVg98bSpEifBN+POcmO18Gh432XCYcQ2npf
AO+9bHY+A4D2crGFTJtJnBaeg+Syfqr6f+6JJZaf5/rmoMg/MkuriIj6WGKuHiId
3NCiW07I8+KznLkjg2xsFYdzPg66wxEOy+lBFdxa1ivhK6hJCov5EStCsbRrxUVF
jdA3Peqfyzr/hJW3u5f2XoUTr6H594/lh3j7EFvd5lk=
`protect END_PROTECTED
