`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HgOgDvLi8nifRx8qnVTnPOgOnvbTUSyNHh563Eb6pwYpqGf83FTL8ksQdCqvP9rs
bwmMG8f4yZRAojXJEKgRVjgopm5cuynrbU5AQX0RgCdwfaSFwWMizifasVoQJvby
SVTI2MUmD2rH4DpWKv8UmnYooqXNnqyGew4rrFFqvrsp6M0rKD0NDT5CGTTsYE0I
XcJOTit1saIj7uf4KM40yHcJUxmFmr2VU6PzPWvBVPYf6faPPNJFR4KvZqyu666g
Rz+4ME9+htyPOYSR9tznKjIm9GetPXHe+sxH6Xnti5iDwDANH7gZp/CD3bUSDrFi
lAP2xm/ASgRa3if9NeDqoWl/qOMpGDyDe3nhCX+5yu6L9IjKnCyAUf5XHWP3aBxt
tvveKY7D0w6xT9uWdXHOvDt6R5sYiGx53nBF+5mFUsh/YtZojfRMNJ9ujBpHjy0I
ULtLRoEnS7TkEbcqrsWqLWqJ8vHx0JB4r1kXDeGjwLQ=
`protect END_PROTECTED
