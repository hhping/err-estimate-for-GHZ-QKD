`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5kSxPGV4jWItO2hgxEJRzl0yCx/l26l1QvN7JPBLT/jVLp9brFmWW/Va2CdU7eHH
4U76V6Y8aPFxkMDifQdCvwdqiLd7IlKpYnEwVLX6LdPpESq4GKfCFw/KdjxakoJX
I4BPKzh+Oj+YiTx1IuUphMbfWxnTA1ba6D1iGmXfopE5THBbb5ZxyEpYZd2bhR28
LenkkSFvj6mVcVEhTLUVqK0ZcpA4WAort7DNPN7J0mY44EBIa0hPh+rDx6xqJmYV
Ud3imTnsUjIhHfn9msMirpaHFsuZGC6Ig3hJwXO918wO1iGnHf9nkg4+e/pwwRow
W+Vie7QNmcrR5dZKGpYLT/AziSttedXuQ8yAa0oXk3dMXsLfKZmcHo9mF8zmWNix
jhXgOpRR09Z5EA0ocV1k8gNAjQywIT2R14X1DpEmSzyq3u0CJOzfIQGyBGt3MWRV
XhZxTOq9DScgXSQvPXE2mVp/096w53KJzlkSJpmaxe2cyjb6yWUKjK/q9Ewl/C6F
AUP368KTH+rKwnRsLGqx+Ph6qRX4Av3Y5Bampp+YRC3Soviq4bwnWWNn9EtdD0vn
tnmOey1/oS5/JpIjhm7rrhYvz3gzcvLtzgfGf8mqIgSEdjr1MhMN2y2mYWrL9f4H
cveij1pXxYP9EIvIT0QiNDuDyFKFmbiLmWqVnY7w/lRlsetRaMwi060NHeOWvs8T
n5n6GST+isGOACEVSEpiVTxTCfxjpnjZvk42Qynl3uovksEhxIlL13cAaUReHZyC
PBNj4QgXCqWuornh9xbxJiEaijxyZIe10iw3PIwVP0efhudgNmQA5YbkR1FsoPNy
VJdyIZp4T7Ia26wzij3w+5VPYKdD5do8wLzzCySpeBUx+CF5tzicZSUwkyH2agja
zoo4KA8eJn2RcI5+P+6aMkU3yV5qOYTr4qSiYhUt/8JiepsO330ee4ouVKoa/4s3
ckdWxTz1hr5TinBXde+Sf2TboKbnZXrWQsrfc5xkoiUzfDPP8xwggSKt8FWYbDwC
vC1ZBtOsi60sXdlptEQqqt5CiMICfGnIE+8FOgY9Qpr0dVsX3eMTzFmCitPu5z60
tqvEqcmwQqtX4sfQps0VUfQVttUqUAmEERsFRhZPyQIBvT053naX1mOVvVSF+wki
dI3H/IHxZxLOM7NnrzgrtQIh7lRIaEaNWNRPZGRFb3HQb9mMbPqUzvIYEkbIEtqt
o47mPNdr1t4QE+6rRNy3MdvHXV6zJSyAoIfX06OqIGVNepZ17b4FtXhf7QHV6XFI
ty6i6QggdQylY44RqIDIM9tD+ZNQtgc6PNCWcSjHuXFDWkbJdqNTtaZAdZe2l962
0A7y0y2o7GsmYDwnyrYPvjJQ/mr8vnPq4ORLqpC0Yte0dOtLvU9/kBuhKc+Vuvw2
mMVRfYfgnTIWky01V1eOjlnDzwzOjdX61bLulDFBsOIJUkHSR87NkJERwjoAEy56
sfej7LgFE4Qk23VMmJcj0fdBzdrVkssEw+BM1wwt9ty1JFProH9fOARMQDj1BX3B
5b+VBQBthzzHSUpuVl4pkxlHQM0dZh90msBmn27tWrMvwtQh7h6hG9Me1I2xtCdn
UCo9oGDe7/bgzYtU9p3bP7rrgmO40zShIghPsOs8i1rz+n01loc+YcDxBxQVy9Qx
reNmQW6/yT66pwPbI10Weu8zjyek/rEF9P6nbwfgA3cguJd5BfTdto0EywqHStEz
+SQvEXfdJb5LW2mIfOtMbSQ8MBqCN7SphAd3dib+6Z494GIDLODkRZaYXK+BjV23
t/wlIdSz4ZyrldJk2bXObtQB7GFMLepk9Ku2B8jB2qWdDm9Zl7H1ZNyEJywlNiS2
N32fz46G4QDuzxyuD6a6UXbS7+GNJP/V0wSkLF1rGgMxxIFLfGztwozHCnXvEdsi
Q64XKCbjp9uXNHPELm+yoGFdkKBp2pSW65GC1ELhNgNjivN26jgMJEnPG3NS9b4J
A1WvznVfKHNdfzbax7zJeLt9aJ5vnhNi/gumMdhnE0HiEAKf0T1fUyJFA3zuafQl
mZ8n1Iqpl6RilBxUOCms5rpBZlo2CZcCitMnTtcMB9OFQkvBgGhjFGjOnXED20EO
0oJY0r1Xztc9VTBKVhvxOMxr7dgvlrD6odgkGmizZBYjpVam6lr+S10ULJM8vfZo
GKQik2FRT8qHT6UZU2fZazPzHUoDnulDefZ2GOGyj+A1iz4XVt3+JoJQLtsmkp4k
AY15Jtq/2R+bqeTEmvtV2CZfXpJclV3A6Bd6SkLcmIJ1PuLTvubDbcwQgjQcIBcG
+1VZvIbuPAxw6a6Z6S9Z61j+p0DMonegAo0UcO7Bg9gYnwNr7+yvooRqZi5AVcOh
sFc3WxAdaRd++4rmNz471xJtDDGxrbBgAHGfQ/lB1Z6jRPP3UD4r0Eygb35E5z8b
75vqkRR2erTy0VOTdNhRS5Xv6Y6CxFEIZca/p/7h5I2lAkUqXcA2iIAL+1r3psgt
O9xrIJhJit24LVM7VNOJ+RFzbfl05sRWQkOysTy+veHe70OLAbkYRSmEIRrob82l
lY7jwkSwNpCLdJfXIHgoQGY/o+qqUnx6mOVmNTGLDxOFnf8heIe/eEABtEob/4zC
GPY1nwY3bQJujd/DjGZnSly2hmCC/LtvAX3/vIuTd3s6Se2D1kltRXkSfL0+0fUG
wuq7TnBHKlGWs9hcdIug1GcVV3aKgeTzC/HbU0NQffvHAl9k9Nxbx8Xir086ObiY
Cg68f8ZNc2reTjxOd6d7avsp75DNFq7E9xoKonOreniw4ul+KjfH1NmEuJgVJA95
sm0qJKFBxfJWGPJwUkznC1E3aa+UxGzxYFUmAJ8+xUEGDGnrt2ZAcfMNILO8xOIT
KAsivu6ltfJfbHArIJ73fsIpPIEPLstioQT2phYBME2aqGwfo60i4zb0FcC3rxAw
GdnXixHyr+5h+FJhZaxzgtunu/rLi4jznodMb4I1wjCJQNQCMJinVEVVSpy4jObg
OXUpWzb7SwwRjMe2AprrRRBruGQUsc2OwFv7S0CwHVXV46JqnrWOz+WQ5t/n38p7
S1fP0CSJ/NxQyihstI9SPfKVfiO9vj8r/lS6EL0gpyT4eYp3GEw9RGlfejW/fEqy
oP77Gt3VQVohzhoRMZxW31Y0177f/RZLDp8jGQzxUClzELU+z+DbWIT3hA6LRnAU
v1I/5/3jX787yjHXnxxSY/MNuaZZ4THhsqRDjrdrjtKTv5T389JVAAKSnZg1G3Vg
6HpiFAXSxnsirrVK6R2x5FVlbppOmVpAEZvaQ4B6Yw3R6dMI5lBhKo6MRJTQbHjR
ex19JNZ7z/u3u6MeAnz5ZcYrSNhBmmwFOeZddhiBZ/U2pNyD0t8kjq6OKq+o6YTV
/S9OqVBLUHiiCxYVAyX0kJXOASiTU1WL5SJ5Sz1cLvkOrIUOt1JxIn9thUXydrOz
3j9vESc82Mvnnd6Yv4XSY5UCfZZ5Yj4Adob0isoFKC3TK4VR02KDSHndxpA+a7eO
laE8aZiAV0++zgG/hvm93b+a0xjZram5+WDG947MibtJoH1zKtQHtX+DBOY64jZ/
DggVLWrChG/PWRD9Mg/dZMHafoFmAif8PDY+BaWJ7fptimc5TsECcjU9zD1enZh0
0/VM9SV5N5j9Ax3HrcSucBVkjPYG+AVK5kXY9qHtCGRyOzA79C8ZkTOiuSeJtsCN
+r4lQ6QptsO1r65eLA7PE0sbor0DubhDHFlH4GVfo/VzbeczaqFSeV5uJ6vmkFLo
GxO3zhjH1syiZLF9AT7p0kY9XNVdnxGaP8FVuXGcExrZAm6UdwpA9EWuvljkizQJ
m+vzrMaNUoK5Jh9wEFt4VdiripEUQfFV2loCTPkN7jujb0QmQHKT0SBH9neRuY5U
FK28+Epjx3FvnNO7sgN/mZUhSsHhxVAdw9dgKRmoANujzFNLCUrzU7vZgl8wuoOL
o1l63qXskJqm+hzHiuqpdOllAzXxuZBlNXc5aS9rAjLXovgrZyYGpmEfWZiSTN4A
KLp+ef8drA7TBZElm4wGmi7uyP54q+wjfLRYGZr+4IE0RqKaRPLLggbv4AT81zl7
ATXKhs+VMP/WsfShcf3BlQ8K4Ag3HuDnzMpz9NogQm4noCDeI9XEnLJrffN9M9kF
ZPoZgoyfAQ6E5uPS1utRqy8KVP9fkogK8Mcxuj1UysxmUUNlvnxlSQbHWKvo8AFv
IgQGyCNoTKKv5N8A0mQlEiCJCBbQZppkf8C5RbdmyNSJMH5+Pq5d1GPA/FFhzpZa
iN9p639WxArkR1VIRy90qGT6R3txkSXCwEmCcjWd8hXrm4Kqn2LRgPWcswPmt6F3
+1uFkD6qrRjin2mjrcKGgoomQ3+68xA9sa3H87d8HbnxTvmKHoJuy8fLjndoa/HP
mm6RFrzjYlWR1Zr7DBlirfxap2Q43qudYxSA6NIaZPBU51ejXEUj3uqjnqz3w995
LoE7mRIg9VA+ZqIDv/5RVoZqJYHiTx89sr5h0NnhpWCMTynXznJd/5rwNKdVUc/h
dSGbXfcwy/s6jYM8AA5L7MO+UxkVzUty7tAMiFRvrIcBCE6DO22a9iuwdy5fkI4q
eX3FF5i5tS1lZQJJRDB4hGsdQllBD+QGRrgyng/u57qIKQn8B/5/Tw+bFfjFicwM
y4W/8qviKUvl5SOavy9TJNYKSOqEA4RZfdU4WNKgrY8cB9ocyuhc+UdajaIWxwh1
4XVBlMUiRjDDET2rLs23PjHDa8LZ3LJyJNjpP0Db+u3qo5vD2+ng69W/XuQkFjtw
vJ+agvtLIJNEvw2DP4Eh9bsUz3QtCFbKHg94r2PMKD6ZwX0johERDPGYcyNS66Qs
uTS1udiNV2Toe9qeytuVR8rBLXqMTdBLZ3GJL/5PEylJka/hee+pPkkVO2cCxLea
NMgabYR7KV8Wxqc86M/aAwLTvzJvVEWcn2S2mP9AUjBgKkHznfhKxGGYpqB9pG65
SoEU0yTSUaZvNCs4JMU/spRHqMgma/7TqngRBt15E1ejOmT7KbcPYZd1Y01SVVae
NphDggAwntjs6U7pzqLS10uosnjVHS87LjtJRbSCR68h75+209gLBQgZOEft2gbv
BrUI1huUuLmjhl7vM6LgSjYIaeh/iqKa1nCV48vBPqypwyIsubUzOuRee0MksRgQ
GIH9/B9utd/iFbyfgQF61FOAIm9RF4g5OJID3ine4ayd+H4BsDjsc6Qi5EAVex49
oL9kAV7n7s8DlCFAV8H9utsc4Wfq6vZwjraCL/phkhVjICVnEIx95/LjU9mOt/5d
h+mdtFu1YNf9FPnBi0HFPOMjTZwRzntfC9I0GxF9gjvtCtniDmvEiCGznIYy0jmP
BGtwbg7WePn845LrQ38LN115OqGa9bUCAuY57bBW71ky0lPeBx6BQZbWo7dUP28Q
pAhgPYArbJNPMHzmzHRP/zg0bwO7K5HMRcwYJVD+7uMFx14VVdVEcQpayLgmNMS1
rPZgsR1lX11aHO0uJ281v+C6UUwxWc31g8Ytfh6K9URhgy//onzqB16QnyYjR3kD
AWzQmKrnWdSl9ZJvZBAX6LXYOnf+qfu8Ozl4m85IR9dd0tjF6HXeCCpjz++kawhS
bHHvFnHEXMrT1j3vSLRBHfGystVAAzV0x9yB5eW5Y2kxYa+GbvE29FMhHsk7UxWh
WdqLQobgU2kasiL4zNdC6fqkfiDXSZNjcIDhRMeIXwGZg/jPd81+yaDXnaflgW6Q
nx6wySxuXXEPRmd5tVYBWci42IMDpw9IK/FZKeHL8Rjbo2yoaIJxYWEK04xwyUy2
D+vXmH6bUwftDceXlelql4kKNeUjcFU43LyL+hIC2p0xxiBZzV18h3JAVqmFzsU7
jzPKdjtnsRzW4Z04FiCgRO8ueoEuxKXbP67cJg+nKhvtfLOEjLTkb1+PIP1DG7Q9
GCWHQHfxIYqOPBIHpDzpp4X5/rwxnONBDoD/dSMdGpz3i9h918++rFMI/aQVJdbu
/DZw1H8DUog/l5/YaZRniSCrjtsOt4As96qqVnndyw3s53b5KIdogtdZukK1PLtc
Sh8y95q9T7vH4BSCtCCrJBWxyV0jfF8P3QTH6/FwL9E+VCs6lXAZ6AGlcwLUj8Xp
HVyqELBL0+hBw3RzH4fazGALtQzo7OlHldWPS9yBW2Rokz2rJiawmY+uDfXlTqhR
uvdyzeuvI7POdrJx+Chpgh4ycnsq4/T/SUHpYtDYypDTgG7By7pEAM5kZXnO0E82
jDwu25rz4DmcX/bYMdxK0QoQL8NfasAULzPcp0chds3WMS6ZWeuBxtQp06gn20Hl
j79xRvw4plXmh9mBSrnYAD6cctZ0oCLP9ZOyCHOHhdffPJd8e5/r/dDgUqMmnw0i
Sm30mdAJKYOLF7dMdgyvyJVdP6Nf0m1u5pSGuSh0zBout8gpoTeNKs8dhUs6IwwI
37YQedPJbQI/Vr0Z3jxY7bzBSbbp1ELyQz6Aatud3GYTp7E5b+nm6piNr8S7+tg3
uHIfeE6t4OlxicLvvRSZDqeQoACVocMD0aF+WhUcqKcOGdh9USEJttCbzZu+Jvvw
GqhrOBFJrnEbBPqCypHpI9cKu9Bb9wISZuDN1zZgy9zSBCI8irC7obd7jve7nOVN
wo6s1YQsVaplNYxSDE8h0TqXbgPQaf7hBT6AOW8LGKGS3i0GHP/OZxuJ8AnJlmWW
3WYfiB7irOoTd1goa3O8aYCoPNr5k0Ov3ST+swFqloXLe0XCOE+kuMFqw0JHdnOB
VyhedfZNyYiedzDHh42Oc2yAuP+xWGncOUdrK9vzRApzTh3cUxlqQRmM87J6eUHS
Ky1psoiYDVoSRYX6FQhYDMNAhhqfEdbqVev/0CU+RWQKkaU/y1IhKhIEVE8bo59K
wdtDM0RVdlvxNQchA/qVlLW1xE6yUdD8mT69wU70La9Z36JzMIqwTxum+cMD/T9O
UTKtHu3U0FN1uMf9k1CZsC3OgZubNFgoNIF8DqT5ZCFoZxOvoQXJMiPmY2DeSXyk
HPLCuyiPrBMYUZD669ttVqeIRhTWfo+AFKvyntHX8QT13E8FVLP04+3U8py449vl
RQGe9uNkqJz1HXa3JmrLKXPuV1ONqCY6uXuwRrjlr3HQCxdkh+VLavAuOHMdgQvl
8Wpag8QKGS7DK1yDACwDZ3qqFNQDlVTI+HZOhvkvPApRt9Y7oT+mfL1YXHOxoT6w
x6eoEUIiZq4XTlIS8doIFsiNf0OJ/rdiImAorHRcksWd1KMTgwXoaC0Mu6soVwj4
es2d5aF4q+GADr/8sh4QGU82+wC2RVdt1VInHvbjkTgQUYtRoqB+jGaHCAkBW6iZ
tH8puRuQxlmbEqHtAuaysnXWFwH9ZLOcS+pHqyJuXnHlqPwDvU78YdRMESFXWZ5C
4ARqR7grINNInQK4ZbOm1u2mRq9hEJCZjm7mcXJPFLGPtII3Po3iOJdk1v9rdoKL
NU2ANT1285Yczog67JD+khmhQRk4AwJjtat82UgSwaghSw+zDkLNAkgh7wbcQ5aI
iBzrNQvjS9qKb6kmuDV+y4n7laOwJVZRjKoUJg/aatTvorQ8ujthSFsVKAskDF3w
jpHnyQDqVlrQEeRVDiJMgWJD2LqZo4XeJwQfdQaGC0xZAP7kZvhqO30wsv7d1RTv
84vwInYFohAmqtL3/7sqXf+tv5tx0oBRGDpEb1uvjX8PtE/Z59/5du9rre8LueAY
mvmw/F9Dn1kuPJF3u4pgsAm3kuWkV/v4+ZFzkJzGu4qXpAA+KwmeYi28RzKY9txA
jCZ0OjA86vc99sOk2LnXkJzVHjn0znD4GNJdtC8C6Z6R9bAMixAmhlA694AWuWHd
rA+x//kv1ZnqVKnDgLAZllyFHuP4OzwcebGw/4/lDE0YC51gV3ayV2ECVud81D4s
NaOE1Y5Vnk5/ribiz9I04UzwBivTIw2eC5fS4qVAGsKJjzwRZQOVN8VwypHxebgo
KwFBRUAbf6SvLbgWefkUmfv97YIuxRGRFpeZ/P0CTWpC6hEkJEZm4ZUt0kHuYCXv
7kHtbIREThv56icps9bs/ecvZ7lJeaSe/TLZ6CJx3hjzG/cOcdqsA1r2kIYG0gdO
ouLIt39x/EGcT7Udvoshi3nm2pHxMqyIN6OtxPQDOHSzcj5gCJnvvfK1oRtWjd5x
60d3cDwpLJUXMTpUO3QoaTzx88fJNZftklEyW3WEKLv+HN4jLcerhxlGh7svDOwX
LqPee+klDXZxOI9772sGLiM8MozeHdj1zJbsSFyaAQRJS1dGbIpLkUqWD0Gx946V
o+PxxVQQvj+JP2+HCeXO+VvRl/ETj+NsaG02MhrmhwHgzwwL/UpS5mYhJrM1FvlF
mAlywcoUMGDjcaXZA/eqF5xEMjofsC2MP3ayP4haJReHT/fG3QDnvq/UHGt12d1h
KV41faBIclDOcVi5joGsrYEooOjv24/u/CEhmizge01puCGhQV2aLsb3g6kOfOiR
Cg34ZiM4QGqOBL4L5i36ECI11WR5czxqotpJKJCK326c+t7z+xvTIIZdGRSkJd0R
u5Q2/UWAy0PxqJrMzVyL0uMchlmp6EUWVIdkmvE6aJjDcdwS4WX7nhMTGaVIvYnL
ZF1Id3nImZfPw/UwWqNipJpcwaXYykhkInSXA0HtuZe9zMAamymgxAAmNjtgHJNr
/j8/GGaY7+f73R4ylYxGRBwztvbk4kN8+NdjG2F/1VRqnoopfBQ0vlg9AuXcdEbw
+n+R3fArjT9htKGXzpqqUW+y2Fydds9Ai4tCFwvF+QkYA0hnwrPrR4VL4pB0Zyx2
NMO2tat0UW99EhxqDsshQ8Mk1t9KIcs5ert9ZK2kl9MYfvceiSHR/dMKZJ+NZnzQ
0x63o2IfGZqa1Kip0Xqo/4KBv75aBl/2NwyQ70jZpEjCuRrd5+GhNZyrZz+D/Gxi
aEBW4WIyzo3Dy6cMqTY/2jnR7EF5xezeXVCN4emZ9x3WNIysUUXqzLs1i2sqmH2/
U6KJ89zsJxu1HzBUMObAXhSFsyAnWc5t3GPPtSXui+TrjRnS1umfk38bi8fMUpxp
ONW3P4nC9oMqooSQd7bCnHL4t8UY/2pFYKX6+0ynbMJTd9uoc7su0elE7y0oPJYb
sXS37wgDcVweTJ9jGzbupvmgizHfrvGvfeSXnhfjlWbKevfKSSkdf6nrzya+TZEK
MqPEubUNYQe+GbYb/6AmAWvLtngHpOk+uhYM9p/ZBk0mEprBesQUr5WaSLGu1ABu
5wKH/Vmq5RCeS6q3fdTFdBmdVbFepG0tuZJzAcTZ9PWfcOaM/WnY7hvKBA6BpuuF
9bXxNL3eLrN2unk9eMHadDjmRqLO23CqtwEm49Iv/4T328eZJ7vADyLcio2F6p28
jhX+H+E/J/S9aX/Fh8toVxSxtFDteOeYyGe9GoR6rIZX+THxsRJVgquf32vBc2L2
syFpg6aX2VRNHjdnJfMtXhBXvOAe4QHBYg6FHR4QC0h5uoPFzqQX5Xq4f9lAvmjg
oV/1JLNvKJGkCtfPFbj/CSpNI93FNR84AqnwU4SEzMawFnr7rW8YQWRc598hBuQQ
tVPuiGgvPUqEtT0r71MGMSV7U5nrqjFK3rahvbTghn1PrpJ39UP6JRw//qu9/KVF
VgYvUTW4ZEwVpqUszBm1nzIlmvEUo8edWPFa0BsthcADdUyhXququJkTHWlj/jK3
m4EfsqqRMPebYX542Xczz7wvsD6lW6UT3YSR0FtDGu1Y/c31Ed4b2ASEDHbCXf8A
v1G8kwznn5uqaBkbDsqOS6cFyWImjsmoHnLUQvbfENwVJKe3VUi4JNSVBsFiFdJI
ruU4M5WxB/0AXX86BdW9HbN8ojtiTmL49Iry41iGo3QRLmb/Hlv0OIg4J+CE8olG
I/mU9n7xTv7y0naCouRjxcYc7ksyOUOP5y1K0Z/0Gnvd7KqUWhNfECcVFSefw8qr
8gg683GayQUwD2B74C6kHQ7iF8jsNLLKOelLUAg4UDsVU3n6VQlvH8wxqGzAE77M
O14xdGyBE0h/ZiP+LLsTdrRBL9g0NDNGcOYkKsw4eyT00JyQVEYCQ+u7u2zOwa8H
iIgRSqaImdhJrACxWRROKLgB3kctmppmA3v1BHyVpxJ0AIFauGme0Y9DO6QjkwWq
OAEmu4Asqs92Of7eF4KBG5ZXGnECYCIoJefH509QyayDGrkeWKIgBTe+2iScf88a
56DVKgeEKwUEOEk0pEijC7rZXIZ8LqLiixPU9jV26Jmydj5jBDROu9qa0bs/E1yZ
slR7VTMB03+CMMZyOrbz2ur6UUFM5gHWuNAxklNr+D8/vX852PyddXAJ+BFlKN1r
pSb8azR0gHaxFGhzwKP5f2kQFDJBeU1kbdUkXPAn7vlJSWGldw0Cj8rmQFiUSBJt
leiS9H7484VR0ADlcYLjTczFZUvUWup+P4k//E7EvW/E+N4QztcMCnXckBzKBZHw
uAfkSfVK07wFrNFnxiGBrHD8zDggsutN2afz1VXMhu7hARdCgSstMUW5RhrPBzj2
ElxQ5ydrCUZ5gFspe5QfXQC/G0uuZtrrjTnzvsVuDaOTfIweKT62aGamonyA9VtQ
mUGyR3pLpC+JNzyLC+9Cyt01p2caoTY3vTedb2044AG7UX7zXLE+cFxVMoIPaSK5
X1xBqfOT/1FLmy7y676AEaaRjBlIm76Hpr+i7X3sacHRlnZQ4eyVCbyEbj13CFn5
cf8wsFHu/CVAj6BSZNaSJkURrozrw7Ye1OCQjItcIflG50xRgimDnec3MAyDMI5j
oHakmx+Fm2UYRQ5w4BXTGlV79iMa1CpB4XtqIoRqGZ29Kf8CDvr9ez1mMXnD8XQ8
YuroXpO9jF8Iqd80cRYFTVEpUktIL+sTGDKKBrDJ3mp3MO7Ya+BIF1rCOljVJirB
eUCTpAdCWLnuR0CrQArYquj9Hm062GUw1Ggu37lrCsbIAieSeeKY4ot2Z58t6xqX
w7SJC89vk3xiKwRhssUK+7RDr2FPTwP8AFcPPSw0YEu4ndFoTFzssXB2NhNcRbGB
O2ab0/8b8owSYBOw7PXUEgXi5rBGeNdXNvU6fjeCsa62Yzab8llhuE7bzUALm9XV
l8mm7s7d3G7zPWztiYI6WfX7zbn8o2EBdlMQxO5YvxWD4g3EN2OYgFyBU+E0xxOk
RrunRegK5C91YRcA/lbyYageCmsxM0D1CIeAhqDEE3tUuowHOownDkUqhmNnMZ+P
Sh2IIUIUpRWCXJqhwPVSCnL1jrHAeLYuWhguLrUS9vJtNJOOQ2OwvoxE/GijXlYy
OL4d21Fkk6YSumve3RgkD8ob93qrVz4Kx9nGFG4u/4s5TnnJYG6ftsO5kMABEDeD
4e/KZM5cP6iM8OGvgEVyrI5w1lUEQhy7LJogV3dBVLK3dU/HjI+ebjpYsBDJyFl5
X276PTvIr8hmJk3CvbkAbf0idMgfBiJIhSm9UjsArGJB8/rrc0e1tLA341Vsk4OF
rLAxo/t6MSUEQZqEdcoZEM0HeiZUMxrlJ8EGDb7gbBU0YMo9Ax9se/Qi+OUa5Fvd
JRVvQvqsUf8RJoOf6m0lubbDtzCc3506XJ9LvG50oVAvywADjF21RXhBygEsiwcp
IAyqGopv8OZciGMo/09jSLngPIPAKpLDHXFn4jL7fd5PsG79zE1t/2HBQ0wky0AE
0uFyguJ1VWb6Dqq1ADXdUPVI3eNT3sM1xcqjxIqSP732KHiQFBq1vHqQzC74QzhD
+nyF0V4tvzRQmSQ2FhFPRaow0Bkgt7D5UDXTk/+00OLc4gjJPGo9xqEO3kH5QeJn
JDEdGq5hbkdYKnVYZ5VkMVmqH1rz/j5ZaygPlYy+RHlCfFuBDq5sMPzd98XAy8z7
iBfaKSo77RYjlZb6k8Mfazg7bXMODtUOLKVkFm3vs5Zq1J/U0lCGCjhpLoOXhXjF
ek4y41DUMP/FhoHdu8cQLcwleO9jwA1GdHypCIfCbMrG4HwKYcwIR0NVd20d8mOw
aQBJ1GeQhynVEZWUFzRXxECwPgEkeL+tTuUQoLxS11gl59OZMQ21dOfhbCwvHdQE
MjqtmrSntJO58O5g++xlBe5ZNLItBqvgyP/HNeD8VUHEmDraM69eaUnTJbfZz1aH
KNkG/PYi0fQqfJcq+RZmLedajLBVQxpwYJf/lAsPzzw4KB36fXh0AUaWAQA9Cdal
hCz06W8ufavdxfcQObxyw0vhLECvJpRhIf9tSfXVrPdjhsdjz6tOFiwqd1qDW77C
sPj5kL4Njf/HgTzQ2XlTb0Hm08P02oxLtP83nBvXhE1di8NUxrWK6Ur/kNlUK6lT
PmzV2gKPJ0PqrsGZRR4ZKaabuSAZFNp93bCMrRCl5wnMH42D3lJ+iGzw898u5Lq3
p6sE61GO85p188maU3YnO1h4ineGjWATe4U2ESNTRtlwiS/ATgL26FuqkkAIYUtG
+WLUCE+oTeVFLrIANI9AxGaxtrL+5PGJovb7ruuIgSFflJw0d+ELpA3w4/+oDS+X
Y+jPVFt5LodSXJ0NAtamtmNa4tN6Y55LYeKSOzocEs7sNLjBBIUFUo/g5fU1UJ86
v5X3ABN5vqv8f+dPEEY+jYRBaX96fN/A/2h+dn0raLPfWRBgbuXvhiU1FXthjfGq
G0gdAcOh/+wG3l0yBEbIRX7RXyBC9dXSOzRv/aSP0qEoZd9laI6ZQW7WzBsDT6ql
iX4tKAsUTJJnbaivM3nH1w7jv4tNGwIuiyf1E3JAs/yQLBSOZ/T9t/mfdE/IpvxZ
OSC3ZVpkxoNKmsBFx46TGfLIXaktngaD+W6DSzNbaLCOlm6kXaHlqUYxRHlgxvP2
z5AF6dN0gEjubsSbdXXxcHCMrBAK/Dy2kQYvDrdJw2RkOgWjx+Zu2SiTtAE0OT6Z
Ug6lkP8MZtCTqlRUVdxo7nyNBx7y8fcnMvppr4ehJUYAFsXHTReCW0BAOyB59i90
NQ/SRegz3iB2iG8IZD6Xfhb4ytobh1Cv+OZ2o9dmzcDimrux1TI6T7Iaubq4SwIn
vusWApYahJY+yrGLxOvcAUvu+6JLetDZhjgYJko3dQTLIo7xG/e0w+2wR2pdmlHr
8nu0CdSgbeGZMavuEuLtgkTFPrXgXUQ+12qEGNqnOWB2jfG6eA8pUy1pRsaFlbn5
axVAp8qE4uYxrwoJ+IOigtR6efwXqcO4D2Hwz6xu5eD4Z4xXcdBG2nFlX0ckW63a
a//7KIhpwZPYhemjVrJuV6vLxyjut9lpZf5dHlt2zZj0dOAXn9b0iY047g+GqQNW
cJMUaVo95HKYevo26/1Mh/K3Dj89jPSLgVat4exSjkp8SgoKj7wwJeyhn60dfQUz
0FMNMiq1qUDZK+bBbsGLdTXnn/QoVq+SZnPfAVYFesm4D7EZiOn6gzDr4v7K1EMu
LS1S3fl0fm6BL+DaujqYqQESbBXWMR2H4gKWHLIs9gX4eh5Wwmc5dlxh46X17rqK
tXbesOsn/+y17MbErFDUMbI6hchEs3hX9T8azvrcfvUjT79FxRivUd1Y0PAzAq+y
jpHQECOlVO3rWOYS+yzxm0OZT1wZZiJXHYz7Ltyn0MY54KBlyH62a1fx0UqR9abh
Af1T5xlzLriqx/uUXny/PYKUBpSk5g4bdHH1jaEf2Wp3cj5pf7FLiT28MnaankaN
6RLu9PleI6uDknRKR37YLq6inCEWmDqhH/5UIQbjiLKUTamachGt6+HZNFQQzVK2
l/ZNzxj1WoCCuJuR5uJMwhOt+bD6K+b3Th0zPoKdF0WnuVtrgnKE9Zfvrr/UQWgd
ledsdHpmhfzFG80rw11O0pXLhGZLRGEyduhlzhKRDEGTYRoCVrLb+tTswB3MI1s0
EmEIqYJ+7VuiCO1hx4iDDVqRuLv5ckrnIlQvLqql3VJY+5bCigEzLMtYqf+3Kmk5
MDztsD/0f6mtz4QJyVJkZaxj28gZnnPA56YjxgVGkeevKAwnQSaB7efW48CSwUwr
dVD5lO8iI5bCUD7kX6gGLIoD1Cr6I6pXsqWBRXbVoae9js5weKAECPFzvJHNjYkS
IPAGhtR07ypf0OBi+o8F1wQexky+wrdNzTPE5afYvqZpFpuZI3UvkG8liIhq4JU5
yNIDHoSw1uHB4qkP+claULMvh9wLwcc12jQE0yBQv7IuQDEVHA5rflFY2pu39gMQ
2DN+rmwhWnYwg56RgSrVbZG5NBucHCFxdESlWh7p7VRgyW79zZLZbDnBKY4uG04r
6BeiGgUWwZZB8RK5BSC0YNXkT6Sfi1b5xe4AwrQH0oKfrx6zF4smL8vBERsfhq0M
6BCmuok6VfJ2GnGHzdeh6bsFtzlQa1iLVysiYb906pqYcHRArEwI6ixIPgWZNL5l
qiCPkeMQp2zDufe1HuT42EPMMxGH09Q7HlZXp4q6ltm2XBzrJLDU/1Q5iVs2i+bb
R65hrRNetPNiPkyoTL1OVhg0dKGA1z5NCOTo4dfa0Q0BinqWv/MaaQ29Io7eY7ah
Q/mVdRXh2S7NkdaBMyPuqGGizSuATipoZ12mS/VmKeAxA9wirkp1v78W72Rz6QWa
QzZ18ckMYrwHKQfKngA7jfvpoOvCs1CekzrY5HisAXRk+6V6l4UZtyB2rfF1iMNp
UhN/7dNupv4ybsGUQQMK+LNL6rmizDXNLARtMp3A4Dnrg0IDSaC1FzAArZq0bJB9
Tbp1RMMysA+ivnr8sZmG+7XYXBMQ7BuHnt7RvbtTdEnkBkM60Pqo4VHTeJt7qjtw
mKCFfeSIA9LQuLGIuznh0RES6bJnrUgXxiN6j5y2xk863y5T1BP8gWaZNvdDxPhj
XQQWj8oJBy2uoDd97+pY5dX7H1KTWVwN6lIUoBuzH+El61kfgOnQnRYGEI+N/9Ho
1Qll9vX9AWKyVwdw2ggTn4qpv3emLYLAaHPniqW4oIFBh9vjbWI1JoHOudJlcLRg
VqlQYo9eNlsP3SmFOMfdSCyip6wX8nOoxdv0OzFytSchD0+0k1r1D0aNShNPYZ+4
OtGXrh6f0pUVFmuIhJ+2eEmJSHMMSbo/isnqsqHBHBNxguFftVUfwj7ycjt55yEl
Sazr128oPi5PE9bIHp8VILlYtnv3y1CNXkAGyd8jPFtBynC5/KzjKmPyz9U9XdpR
I1KVKcozY6xK33R+cGjPpdsU8YaHqRK6Q4balvAeUqdtoqKJbinYJT1XUr3MIes/
L0BUhpk4hmrHLRslR2L9JkedYiskASef1u5/XrkVXJnp6tb+0kqi2d2NR/Pg430g
X+ZRG9JADdAT0jCDRL0Ok++m5kdJDRrvB59vtypk1wtw8hO3MbZVNyG0t9sitkzw
UV3r2eqIaAFv16aUIfCLmOX37n5Fe6qYohNJiSP02fX2pjS08SHMeRKnuBszLxY7
DfxbAj9q7L1irwA5WYaO3/m+TR+hiviPkUsuud5fQ1UK/lnY8mQQeDBbH41RPJS+
oIof9/0yaPRNVRlq6tmAEax2gkwN0kPYTZ1NOE3gbiArgPH6WvIg8LI3OL1+4kFp
zdGH8iAPEVsAKXSXIjjilF8Ynla8rI71zAiNAI/8y/Si2iy5o3vsuCTT3Av3CVr2
E8nLGFNp3JDt+9lYZD5FI/OCvYHT1HaLp7hpvhlLqEfqZLlkm/UP77wXMNd4nTaY
ArCgoh9MoqEmeNaqlTnb1ETcl3hsokqe7wjl76BjWs4fI8Q7WIkWseGE3fLlBEfO
DBRd5vDRZRawhsyNFpGerRA+IY/Qd+8j2qQP16+gWq+PZkaY+v2UnBwWUlfRAhTZ
0eQ1Ffa9r8/av7Rc+G6hAH85OnS0wBlK6K6SYPTLKT66NGWd/TGRZL5af6S+o/Mh
ZGfmxL7xyY0ijW276/juwc/yds3HIytyrY1xcSg6arxhMqo7L0LLbH6k4Aro6jmJ
Sj8/r52zOilQqu3yKwjwA7mZQK7iWZu9xEO6XrPhvATTqHIPyO2wIZyoQyWLHJzF
yJaV7niUvqE5mFDWuPj0XD6Nx+pcLl2ApNzIB3sPuBzJTE8ltshuJA5IUYqicpfI
EhFCxaKn5TxatKXfTs+/PyMJ/W7pxSCg9kA01U4moHtXpYkFpgTnjl18v1Q3dHPo
VhLRzcyLm/9P1591WaEKjVZydPMbybfnNQhXsA3hwg3EGQKYLEKuBVtgG+/PYfu6
8XHcXzlNrLfDCm1jwR3pLOw+2piIr30julfR8+nrLhJJjNqhyzSIsu70ijtAaz6x
BBkdgxeVRDHz+5ix7oGex95nZPtEqSF/e2gtLAHIlLE5+T2zqJ/rfcG5zvmCZRi6
PptoRzDp0r4bLDGZWNdwuH0GuHREcrioB50TnsKSG2pG3u1tSoGk1Wq9gGeCoEKj
1vxi1cE0abcMurUmmDPHL1b4rk+ngz7X76nS75EFayah7bYSoPEzraznFSJYoi5L
q9CkqRyHvWFXJQq3R0nTjBs40FN7k+/avyFofoC5SPn27ghbHFV4oo0tOn7IWyoh
UVlP4cGx4meUGaQaWP1sAO+3JToiQvdyDd4momq96Mj7bRrqg45WhvYjjGJ8hIMq
8aRnAsqK6Wkb1P7myrlKUUS9i9DSeeLVaO8G6ZEkgl1af+UmfVinD2EuNk5bujqI
qNE9aNqv/FQFJqTiIb8K6axhgCSjz3OZ6N8mOKhcvXw49TO1++WQI3MdE/XovEoC
+N+7D2Fcn/h2eThaS1592VQhFubf/Zcc96AEj3olwoi4ixrR1ak0qF5tuRMyGHVb
CB/gV6bTasllyWHLepm7AorQPMvFtKdpTqLuEjZ9yZuxNi9ClkjmyTo3HH7zt/JK
y3EA5d/GsqEddvkONCPCDUrfixtpdH66UvJq3EIqS+Vwl4ugS1hP8L5HPWwxAiRu
JPHbq8TEs/z57ctn2BmMHLx4QZgm51rtzhwDCVGolzSOz3S2xTwo2Cpi61SkMN9k
/mU2Srat2DVG6OIutHa+Z7SiiWf7QCu5h7UTUrpiCBBmLriwSQdAI3phqw3qGCtV
rnt5y6E/mEzEk/tI57xAuVv0cM9YGI92knJ84pZ0sM8km5gfDFQYsfR8yyQhxGTD
SDeLP6K1VHuWMYcBTUr6hq3KadpWwin7to9oocK5I7RvJEF/g4Rt7fGkVapFJorV
mgOJ55sxXVrrLrES3WJHs61KCfilPv68XkGZ+DBiBH8Yi/XcMTzdgqikR0OG5EB4
gMJxclogJ1uLLemfMzthRvLtnPqqx4biD/QQ9s6uBZZmD14JU90PvKHBCVKB9wZo
UbCV7w0TUGC2X77gN7m/O1aADX8Yr60tpcdQH+mcsziQoPY9bZlR6M1SGn7cptah
oF+RTlB1Sd5PHH+g749sNgh80qpx/+sit3r6Xd20ZqTKOkOyG5KjvyS9KtjOWIsN
23C8g9ZwOnBJYK13ZduQtsyJL/3q9XVuMeQvuS26AdCamoiw+ygrc8uMQidkbqRC
wF5txQoITE3Eqdxl7Gy4eBd2znhRv2aBqACid/XUnDbnvYtwSX8fQ6s3XeR2GrLm
/S39NVb/+SyOQ1YEhsodMayS+/O05L/bK+Sfct+vs/1tTfM5NGDQT+VZMaloq+AE
uqvpRjnx10wqADuujtJCydl5OD02vAjesUM297tUrtp0yRqMhpEAi6r600hxj+c8
Y/wieMjFDo5B15BbBuAozkezBULxwjjhZRW7pjCj5eAZt+46LnE+7IUCXlUuy8pQ
QnnDw+oEsKrDk2rClG4ImT6KIJR7u+qv9RC8toOdqzI2jtifKPnvsmD89z6iyrdO
w8GldGBwEchiobpq5IjmMePgIeLrAeyOoQ8062Hat1FWahJSBIgeB6jApCFhze6K
3YLF6xYNgtPnjp2R3GzWn7DPUIYWXkm9l2FsiM1+RR0uqR1h03AnbOcZU6i18FJO
ow+OD2TsXVjO/axfqW87PPSQ1Izrl+GVwhBROHsGlS1/1POei27i1Ojxfvls5nFn
F6lAUPGuMibx/28D/1g0ES7clmdzL23SRedV1CZ4WOvY3HazIoWj1/znt4POqnIp
naScDeX95VdzosBs5gYlPS0FLojYuoKn1mTU7+PqeFsGxbGZ+HHfTafmQfEVshpL
UARGA7XTddkz6jsFUd3TL+NdjS1qRe9XX9hAxoj5at5uWs3AG78vaLkfr3IbEbaq
U3a/4L6EGpjfv5KTDr16haJXKqcvhR7s6Wmj4OZonZvvlvCpj7iodA4I9sgx4g9B
nAblff1BQ0uuyhy6npTsp6yQj+u9woIkvoEa+6/gx09dFf1pjkActu7ezLLwGvwL
3ZFxZp2FuERBoBihlp0MhzBR7rcc19xD49XqSCm9ftYqAkU504/wp02Nc1H7UKZ7
bBvHc0JqzpHPzGcyFZtQi5eTBwciMRuQdHY52Jw8/fbhW5E1OmBODS15kfB8TdSB
oLYZvv9RviPkGqZKEUOFvql1WdF/WzLhDgD2dXjPxg2YJaBINPNsBn1HndDZzpNg
3GHR1CxxzL/lXkS5y6zIrnmjs4eLmISTEtdMpUzmAXV3tosUBcDWxDlq5sItH5V5
W9txLN+DDtDfS9mckNt7dT1O9s3EHujcsww7LVwF8KCmM1WNsFiSOBN2/fQPxC1J
TeHtP0D4roYmaKRfahEMjxFX+w6+EB3S2ZPw99Yhd3lzVzb0VtJR/ehbxh0DdHWk
HRzpgI6ofNWILs6IFQ/MGJBSe3JQ2bbqEEzAnenDR2ZVvevqHV+TMXZWCK4PY/9I
10cSjg5CVi8TCmYeIjl6wkYUpkdgKzY1Mc0S+kbzQL7Li77yZrvQS5cApC+aUkWd
0iWo7cI0JZ4wot8QPbDfGUYbCVDrKxIsg5vEs1b64Z1rJUR8+5Ac5acBpRx4FQNI
TLeuyt6suVpKtsuV/kJPByzIF2j0MdmVYfUhqHyaWdSXzXked6SzPYgddiYsbdkd
62yMdtp7N5o2WeGO+5/JPmNHqX84cJdAFAFtje4f5q+DMiUJIScC44YcuakYlsPh
WYhqopdZwOR5gMhy1chbLGS/TRPTonkLF9jCIErQw7W0JCGMP1iIwEHOeAD6m6hx
nQCyHlGAY01hSRM6uV/wNk2m4XIHMgBUuGNR7JNB9iCXsQ02Qwfaa7b5pCbavUBD
e3oapITQLaksu5JpdoLZIKx047sg1VfSN0r+jkaug5VJoDCC2SFBIU5KjSLbEMS7
0fS8F55CW7jQ5lMtYr21MNtJXJ8KSbP6f9JkTiawG1vhwHj2ShMedXB6mwadnt0Q
+UO9WlUU7Z7bwmoFiUwljZsgfpgZfvzDmlvws+LezfOSUNxLMCA17dqWSyTOSdoE
H1xh9sq5cXtXr4EYLk7PqofXnjNhhvFhV2t69jMo6LYZq0CP0p8cIg+GlsrmIRPS
4cDwRzH9VE+Tt9XI+yP9Tw2rND6xxB+2dLEfb36m6dw1vd59cem6F0F5jIlYGzxp
wSBUp9zOtnt/K5E2iCwLJdYYn7GptamCH3ecwIHy9jcIKEwTCWE+R5BKtRiop9Hm
U8cuDbU8kny1tAzMj/VyuvxYHVq0oBTgbwCh57hruWV/1t9Bo/z8xLoCxf3dtPGp
53H93YTBFSwE7xJCiqy+DT4f2d1PCYoQnfd1IAzXzttu3XOkm7wXMUgJ1TcpLykT
ZJldrDb4VaK7mBfjCLHmHwhJSwHZ6L32zyBMkIF6qeob5joqh5TszqTefitk035a
MveCdoeSdlksY/Y+Fv8aq4v5LJs5abtB26wyDmpjlWtTmLJBmI7PdnJXkHwnVNQx
jJU1ZRNRJ/HCDy5D90dYi4LkJMkqeE+c4r08u3Hvz0aDOpKPd8rU0M9zbtdQERPn
LXWeo6e8g+sZKIHLStkDVLMrZEPpmugv3k9m+k8GfllNLfpuBFTo7JAfdRo5h1Jl
Sh1wP1JAwudoxA4OnVGFo/mfANMKjv5L+FnXK2D9FbiBcPTPv3eT5K9C19sQLTXg
vFQiFeoBBa1ZLzHJi8ca05a9lElPVBepttR8JILXgsnpLLaBUevikv5XlSO/wpJ2
TAfmyce5KBiPTxDAbQt6vJt5R3LDztv+Hjgmz5cUyr6jKIOwVI+FSGXU+pnB79EC
h6MtbqlmvUOdyA+opHl08zNexj5z4UWrs5j/BqPyhEilAm59tAwR4ke891j0dSUf
vKZ7iO0wxlZxSCw4VSEMakgoaNUpBhl1hXyEH+F0Amv8WzewxZs+0GF4DXiVzYNA
O5rJpWTHwhQWF3VhbAKP+BHR7HQeARVVignCZrUVNfJGnGyKCNODXqMZ0Y6miZWV
MRiaWOVsMriC695y4CObiEIHRumGgUcHUvhLsjk6lGN0iABwco3sOWJcP0ZMR7RM
2uJaX6i+nYblzQS+Vk4nzHV61WOvAa+/y7r/AAR9/Pcz8aNJPyTnDAOPQ1xfhyTO
I05N00Up3CBXUnHU0R9j+9NgAat2BEFrNlono2Kr5HaPtGUBkoWUhzCu6R373TC/
OAb3BTPboTLojhTdBk9o4JmLR3X7ly6nvyiU+5ZCESVrqW18a2DZTGJrSY5ENIud
t0mstoAnUk7i3TKZTf3om8zyMLTqCHswxxc3StrPFxXDAxsRDPEUxxMEEMpAOC6j
AiGrldnSm033u4WwYFBS63CIiSNLR/hJwxry5WO7Jo7zM1k0K0hhzmfxJ6DWZTLk
KRwiNy2HxHJUUXTjW/kCUP/fPbUy68kEoCilLUj2mreBzapAbdAMR7BLyahL+Wrg
YocP61T9It/GLJLxMoAEA3avFe/t5HTA5w/qP4VgPEhpDrGgU45OWnaqE8Mxyhxs
dJJjhBoQFQinkhs34YCETzlSm/k9FVMOwxm8A3t4tx4xfy9GROyrbRL6vVbjsy+v
+zZM/Sv7vhbv7rNcG4SdPuClMBL6xc5TAN7rWmP8bQ39ZIe3LJ66dHUiyrWOlwqj
U8Z0CJsx9COLP+Ejzl5+6FIiXMr2a8M6SBTS1C3SM+IFftlS81ESpkouRTilW3PB
+PewQY7HAQMIfZQxtLE23Q5FfxKNW1bOpewfStabb0SGqXMjKhO+cpnf/R66g85+
6KlNNztYDl6v5KFvNxxohkuW3shXqYBYP3nzl8tGeYk//kN8OEZBUXm7B1TPutm9
7mlxTmY0Jp+yasQDFqQK4de+M9m+RCdYggNV8V5Kj62uSVaJlU2uJ1hEz/VekJ16
5Rr7KhYAH/Y39mx4wXnRsbwpjdPtZjXg4I/sARd1IvzwurDcO9lbU9tf+eXu0yvK
V3eLz1QFG867ElsIPknpxtzkoLy2E0k2AuqXQJKBRVKRtTw1knaUVRSK3ymQe1tq
wTWSESkhbZttC/Hb+aMObDj4q2AasPUU2jCmRjWD6FLeIVcy4DZ1W2AZq4/q/9jO
b2bufIWxXT1C57rC3bBh3B1vJ3It7cyYthkOS2Y/S25V7LHQNz3vy0Z0y+ONIUcM
MAfiU4LsepKIAkNRii0h/WXnxSwDOamfLIWKSlrS+kqgmCJi+IE2q6zOCqJF+5tU
suSs9RuhO+WAXj4eYTUe1oqg+ifD/Phbe2cDPCaTR/UAW/2qfnhiM4AtfHxyEGbo
TPdEVBw3DYOGuWJNEasyt69jPMw/8r4DAbfZaDKfh70RJlu1hWb8aQZpxhadw14W
ii92wGU+XYJb9lcdMjxMo3w8Fxcva0X/JnTdv1p1enrmtD1obD4pPej0u6eLivo1
5ZrowOWYzR+bQDQ2Db8oju3MvcmhD9iUkB6X/nVO+rcJi+kUKQzG2Ecx53Zr9YwW
oEw6sneIwuoWy7IHwkqlA2GIAnemSY+mqZz4y6OoQd20ip7zC+ZyqPTboZpMLZne
86zuYcuHLt5m8oXQnYXXVdiuN4LP4SIoli6YcHPMrF7NMmAzOA+RTCIu8HCGuPUr
uoXdNmVp5VaYZNjCczj0oRIQRRnd8zkpqLXEcj5zDwOP3C51cMujDaYRV+Zz/DSu
SZ/VP653fd3edDKKXYov+Bj5SEYVTojj7XPs7pKz8u0skkf3y/iaNL/hhxRVhg17
C8Ry/WfMPOWRuSiIWFBA3wrdzALm9K2zYhCU7WDtxKIqK+3EHcrqu/wGbR2HzDGd
e31fQtbDPFhrl9sOUPi+11DUydX2ZlbKwCpd4hw6ZbdC/bmCE7QSB+nG0dI0zPTn
LQtlmOwfggrbVXAcdo3eKcFAzV2DSAPQyMtwWbk13ccygZGG3NyxPltW8D/58F9H
AdAhwqUIefvtDYbnEcYFapnq/0T8RgzGlge45W74Ny0TigUDMagGFf5c20cQMdup
HjjtuAUUqfcQAjeaY7RGgll7Lh1lJRKV7RpDKFEqZAkyw8MIYZkik3udPHpOdnF7
xVKSXTzUO91SdoozX3HTuNvXaYc9knXAZpvuibi1JngM4CcHt+o11Ll4jqtDAxo3
u3oAkCuUZzETTe7XTooelB3cNBkud3Pl6tBieUUXHlerb4ybdrG+7T6/w0AYEtVC
K+CkwJuYkpZM9quidIacc6SoGopoNUBZINQOSxAF62SBoJB/b3qY3fXRJU8rk8nS
mkESZGXQoksIOVxvCQYoK6vj4OQ+RKqKtX3XYG9OWwvXp0VKSoFRPeI+bI7ojkZ3
Fo4KGa53eft/XWLpfErYjlPdEOLD06uG8ybo6ppYKFb4Ing2JVAiHlZsQD7Eyquu
cJa8MNxWyU4qnVbHsoyie5NwscF9DZZ2CpE3KBL+4LirwMOy5Nw80KPJO/q4ELOf
+P1MwUUu+p+T8DUBzVxDut1PfK4DC5ld4P7jRiimnXtDXjs5rRK6RXaTlkdgroxt
xbdEu0q7pNZKZuB7H0kqj0IC+5UAlffCPTI7Qhqub7/E+3Jkv5k3RD0flVvL/WiD
8eqp5RSR0a79w1ZxvXJPyY7aS+Eb+8siYXOy9vvLPEiUU2z/01nfEjujxpZ2E8lU
yvUuTb4iUOqiqJughVD96c3ay4SkEkx++yuZohQ8HVRnMYXc/wndNcbhNKU5lZGR
hcjozO9MIUgrSozgaGThfDiKZZZ2G+VkjjVW7r/+3ax/WxTbNpmsCgDWICuSY+dA
FUXB9n56sXuQph5FG09DmpG9vw56t4aFWETA0Zvi1KNYq4lNAsZ+3p0uWrvG8DKU
nYac3RyFc8E+L3dcXm/mZvrzdCyCkOD0QfgZsuxgiIWepOxPEkSYRm73vFTp78pC
v51cvJnejkIW36uIbV6otk3dyc13cuQY4V+nOarUNGy7AeQyxwqMd2ivfSUedn/P
AUGPNpHyWKXxB3Kt64GJq/QMjLWMuF24cT4c2H6tJ+5mdI7zMZ2zGYHbCEhQaFtL
jvmXgkLt0YI/lMziLuGIZAuFzyEhM8WZCOmc/EmzSoDIWCy4CIY8j5JFsOIKgGYj
x9vJImzkCktl5vSH9qz36b03ZNt0+fQRE6bT/Q44SfLHH6ezm530e6nRAfkySi+J
bjbe0kaH4592NP+O6R5pAEc34WV9Cb5apIueJ3dd+klknT7cI9S19mBBj5NcmOjh
dZq13SMDYKLgdMwmaiEb3+tsyCQ4LU2qh2oMp7PIYur/qX8lHTFeZBgJ/X/AlnZV
Kq6IgDxZ8LO3FC2rmft2Cg6jWYn8BuIYt31w1BqcTdZyfwp3c54KOdlVQOJufejz
J3yoVjXH4vPaFFwn7TfHX62v4F061xNcUfmrvUprUngXkTFXyUqhiHNrtqnDqIg5
xR+g4uYwnFWifV26A3E2nEfw9QFs6D/D8jIFJm7+85P+pBzEMxgjEZIKds5//N9z
zcFk/OyiUS9QRH/Bp7V6ot4Dz2fdnrGAMFNl2ygNdL6InZMpKxpGhX1xH2mIpCcd
bRaomTBzME/X/eMTe8OBWQzsFNaMYVGpsSL/c5MyQu1iktAONOTcCqg8L5ydG7Ha
TxGfDfNF+OPeHmjoIgCGdtnStmVQj6ZuWFLajYdhP6Q02sB0kZe/+LtRkT6R2AHs
Y9RMQdoqyAAiV2zkooit5fy3pHFsJztvZKf32O0enySkncXFx9m6nPyKVIfP3WjV
nHElYkMIrChIeBzH2fSjPIc3XaXvjtUkIIUfHq/THnX54y43QcFs5+br3CHbLmhE
NwTPx1XjOA60dabMzn44nhMhehLJIlu+oC7RO4VSK3phJ+7UdR2KaRAQYz7Mz9O0
aM8hEsNy+iLX37qnMx2LJ3mYHIdhQyUX1sf/o3mr5Ooqv6wsV9Yt54WzdDQ4lOQM
EX1McHt1rwbeJJh/vxoMkKjTaHAcDvHZiyrDJalz+YDVXX0hYYH6pBMIivAGls13
Po3Gvms6rJdMcZhiWKI4KC8bICmcFNbwcQMseJrhhdqdzuSUg6hVIlsqiQJKbRlH
5ATF3PNW57Z86ZQAjv4+I6tMD6f6NDXrqCr7e8Hr/uxlJo3gRMUZybcMRVFDlmqn
I4KaykVXhQLzkB194+uwYz7W1Fbz6gnD93Fc+TEoYc60qSJasAGc98IcnfXV1CJu
TQtJYgdrEALxXbGMqF42NpxsNBFIa90RC1B8yiTEAoREwMRgpuoxvJENMk2vLjZB
BOY8QVdyviGXI5hwYLQ5VOB1K5KTxq7eryyea878EoCRi/m5QJuKiAdUSIL7BwTo
8/GzgKwDwBsc7HiJnEcnwxdVtJEspbfcL+/5NewJwf5YOnoC5Q8hGXLCrG1/YsYi
PmlndWbBOKZ//eaRiu3aD++3Wxpl/EGWpNd8Qwxs8b7fy0khShG3lKNG6MQNWLzL
pJ7qpSfQzvMUMUWqTxlKkltbTnCoskqG4m/2ASA4gfzD+kQjw3DQdm/tylCVQMHY
vJqdGzBLNnOC2DfN44CU+iiQrbxDhMoPMzhn6r4GHNYkv0ksgeDj33c9b9NpEZqJ
NvQ/qBZskRLW7rIqaDbRGDSxHCQoAeTPrX/953xATy6qMV+YWWPJAn6aCYtP/Hj0
2zluSJtiR+f00b3xi6qjcW0/Jm4uU3NXGcIU8z/9CVOXUfKqyhHUd6Ig5l0w2EGi
icdE3/D437t/jAhC98yKXfFzTmbp/uoNxzv7vntnA3piQ9QG9E28kucC+e4Iz07R
5rkXiazpVhlF3IWEC4KTCZOLy8zyz8c2siK7spZd8Hqgi1utg8TgP9uXGwS4iGA1
DPTdk+QP8DDPNsNch7W0z4rcTJF7LHaz7ooozVo7HB/QR/kkJxPCu0Y2ZtHZA5mn
sljhglObce1YIcdIbdHe3SPzy3UL3/61eUz7kkgDm5yUi9roNh9/DiuA3ZFGkR11
rj8RS416QGGlH+2j0OD7jRpjbD2F/QDs/WFknqV9TW8KksWy2RI/I6Pclp8MZQ1/
5xlfxdpboS0TNgfwXd/a+9blqnDrfSg43lLsxD2r9qRCcvWh1Z91FGvVovR2RyzH
Ur4F2n046tgEuWxfdXkkjHOy4U+jku+mB58z6606hpPL+he00Gs89QvYKOtg6JYh
I3NrgbmUM6EI625g/rfcHtJwA8R7u/fsj6AvhqzXxEvoCbYYkIRiciQedfbVobBb
hdLdV9wERcmxrhR5M4Qap7kzVLjuM4tgvDSeroQfNmeWSAeC0TB50QHsZQ/nHDmj
4gMbrQeFoxuBoHPT9oPLesDjNSLprvQp9joIuBLawxwMAjbzXUwY9Jrny2Cvuzz6
+bo2R/IqOTMXBHn33XL0FRI1IfEQN9ItHrjk5DRjKQgJJgmA/Hu6fkRaHMBxbeLl
PadtDtwAUHU7Z6EFNLnfiXdznTFNKs/6ckf4U+VACe2ff8FW6M5xMSnYaTIHrE7y
NQTsiA6TdSPzi3PJghQDX/LfTDDLTMEnX2Eju1Vf8pZRsELGlUjFmmOooHnumcS+
C4y+C1BWNZs9PQgPq6NElH/Ej8XxHVEUJJNt/JKr+2s+5WHh62LDSc5o7WutKDkk
NIG/AArLgXiesOR4uqGwxJkQjunyi648BWLufCe1FRvhuqnVJMWIJBwaLhbsQXKZ
8KzBgch/zCKgFe5fDfEz4EHudRDG27sN3hHcyPJ8zlOyVMvRgNutzKqPELLNjzFQ
jJU8mnaWw6T5DzjSsJIlIf/RFGudDuSksUQmNP9Yo5XgOPkwrbAg9+emNNuRhn0P
RLi7kREBQxfN0UpXM9Rg3FLKnNx2IlX0Y7k6lIBz44463krSB80o1LXIzboNMRJX
kNDaOrNQTX5jS3P1Hct5wDZgt4LDQ/aBXayQS7tlxo/OB+MkLpMILn4po9Id8fsT
giTZ+v/w6hv9AAyEQNEvus8z4A/kkS6pSaIBXP9RffdmJx1BY/s8cePNimnfNSJ2
cBQYoF5rOkm3AUX12w3KtZ1tklbNLlJds3kPqugzeNI13wFd2Gqt4ORe9jXcTRAT
mDy+eekbvEbEEzAywqoMdh6QQHq7eq8s1kKhJETU2ji02m0areS80TuBzf5Pn1bM
ixtjIOAeK77vck2ZMtwddtOOmtvR3YjOxy15mwTO+W5qkZfOjUwIHCushA7nz3OS
xQEMnOtXy2kFHEtPKr9Myn7LluxS662V0PizM5DRZSxecqbNzynLFm6U0yf7yE+1
Uk0DbnKPixEr1EzOU/X8jR9qTDTbYgwL81CAaci8af+bFgcR4rH1m0dmb+XwrWHg
xSGH+DWj8lTMMfnyRCJZlAH3UGpvZyrNOU2njPXJPjkB7K6lqh+OzgUQkdzwthaE
uzJ3KL6WAGet1VJ4rxOKEJ9D1WnAOVeXtAt3M61hvII9w2U09YNKRfE6yrIxUwGp
PU85rkdI8/5U5F2UjSn2Tfd0QP5ri9V96LGCZGTtYDSpfGoqiwX/9xbsPYaBy8oX
8juSLXZW6EjKp3iT0Kjn8rc+LiGLr+uyVnl3V3qwjvDIWf/1Tx7tOgDtqwwTyPTH
rFcxxM+N9IBes+tR2cMMIPW6cBqV64Iebpsfl73MeNCX5CuwLeiabO5PbYtvbyNP
Aqa09NR4KeZkpBXE1icwpRCPIUY5omtcbYcYj6s92tJjt4auDHlGxjBNEb43n6PM
PdRiSljqLOFTjB2gDmV0U1AAl3C/hPKUoW0ibCm48tzPqstum7oKDl66/VlFA+YE
GFXBXq7dImhXkIBgQBmNHioHVZFga+oJesglCAPfml9rGgt+4mERUzV7vRIwL1b8
InhovQl86MoPw+uW0sPKOm9Qg5VCZ8f3oGDFRGAx/UPo9sMTXW+Q/trna2E94iRd
3Nf1P6NqZvndzQdIskF5oT+x7+mSeYoBszKH/jgD/2VVj6hZsUkUF+u8I1LRq11r
GvO1FT3WgPk074ttFI1S60TrUbo8eDsPJkIVg4KdklMm6fkov/j8Xqg5VYkhp9na
tWYd4N8GyLgk1nfHfh7QD71R66Ansceq1Bco5lfhriX0kKj8ZGdnYsSqyxje2w0U
/Nfndz94shvBCw/PG3Gsd8tKYrWvEZVbFnfjuTtr2J8uhgyddd2LMge1xivhwo30
CN1tsjtoRmMgl32IufbKtiRK8+BP/MZzHLhl8ylWC7B/nrnN492zn+CrHs+FbqDV
/SjyQZ4leCD9DO6FsntTslukksNlLmZ4TTjpWoIZUAISnHWO/gB54iATVVTKpmJk
ft6NQgf/4os6n9TmZrjUt3uDOPKi9eTR+H/BQ/v/kbVdfl6EUid5ebnt++ZBv5wW
dMSnC3uJvS785omNqer7Vb0oa2fnZnPOWXHB5as/qFeoks1PFnbkcUodJitkIxFe
t8UjY2UCLIR+loZUgVZPXEjMbO15WwC+GwlOPt2HzoXwgL32As5TUBJR3loxxjPr
eI6E6urSiPE8n0kDfHZJw9MSRfo6OnktU/sOtNzDymHomhtwpaplYnv+w44vXu8o
H+v0EF/V2iedTLEQOo8wh36QM+yWA/9bU7838WSP99nOxuFCa2HKEIiYGxcuVNVN
fg746sIxLSP4pz5WGdMfdEt90Yr/fMRFiDBlj0FV8ediBLRDmE0qPlmi9f64iRN3
qWdgtDX77TfvnT9MHN1nvBzYUeUcbxS1FZ4/WIn4pvWgLkkgXeQwawtITGOoEHut
9DFJgYFZ1e4MYNqnopXp7tV8Q/OH2HF2lwlbqxUxkjBG8lEiolM0QXpe8bn5+xl/
aKmXTJECEZhDhnEHinVWLy/oUBB4Kw5hdov7BTTZCQ/SUpy2knQc019WU9RMn84X
gx0X4xBJO96acqtIkL2c96uZdg1x39E0bAJhS+xoFp+Asu0GwQGS++V45oMZpZbE
ivqwPGcL78VpeLphRF0M4WpQFSLOE8GK7706a/EMIY8SBu62nM7eyX+GzJHK3a+m
aQrgvyYnWug0oARUwCWL8u13xM/zfy88rNKsYWzikHhHxF3H0oGHw0RBSNYNbYj4
4u2GT7mNQnj5P3JOpGeYEPk26r/O793gUbzcwFoDfSdw4ckkIh09eZQLpk0fCqtL
ULl770l4AXo3m5LzTwct4nlzYGE9wfVsrDYfC1qoMCIvWQ4MlwsoQ4dXeWyOWpK1
zpf+HXmZ8+krKNLdVP9NtEELPKd6IZI+5A0Jr/2u7mRmGw/nOg05RXB7dlmAacX0
BO1cRm2OyId4rBDdbEC9mtVRlpBKr+vylPRV8UsWQFWr3JhyNjau4WzHBLsiGLX8
RBSP2Ui0vyhGntXDALgdY9sXifdmhGFu9SDfrnYOzK5Zilj+Go1u2f4FFqDM5YDD
97lEgXboNqwVXm8WSm1gVjyc0S0jO2G6vAxtVukLC1ltXJlR/CE4fSBkTrFM0TTh
neFxhPYmS2Yt0Pq54rdP74Qi0WcUuYv1VWihCYOb5ABxwckKwxQ7beg75mmBM5jy
YFN6xC36N9YON8VVDTcdQP6eF194EQuBtDTGzWFtb3kVmcdGiyUS8cP3qDOB/oFS
V8PxFoGM4+g35xTKPmB2ELniBRy2kxZdzs8VMDUCSMQN0DlryY3e4wlnXZWCO58R
ViC+NCm0rc5bz2Jn3HyCiluEV5tJXMfA1cjmXlKgJ3fGlltnAB7tPfheQR4L23Yb
CYxNc8zzRggvS5FI0Bznx066x1TeUgnahU3bphUf0hI97J+DeNa/mwYXd7Aaa2fa
93BnlLz+yWL7An/yVakAztxPwGv5cNisG18AOXQp41DLq63f2zSUl4C2d/i1TJ7v
At+cfbYX1fiEMMcJC0QKV3GkSOIAa0B0njMaZe8hV29Z3YpPxb+cSTYrhhl6dLJj
uFMLUruAMMcCv/bojG01+HdsJxZIRNNR+pV3MzDxptEqJpd2YVbGg5zidl+b31Pz
mc/jc2wJE9e7ixChgjGTrQkPl7Xb0a6PjPrmMAfolMJrHwEYJqU7rLInlSYMihhO
BtcKLazY8PnrXXg4M5+3MFh5+xj8r8pl6MS0U9KyYjskiFPlJR/oeA/Ve9JAem7s
PeZtiuHPIWrT8JoRCl1Fv7X9l40sRo5mDytV3a+9vYVxo0uTe8jdE9o4ulnXR4mv
OzUkiik95yZeabhxolT6nUXkA0gLgGKeXHpu/mTynev9sV6DouACOrESsB8X+QJn
yQcDSc6mvuL7sMo5TS3QDyuz/mawutz5XoItpgVXnHpp0tGDvXcIQrXvFa4sxaCC
bsKy3gYBLUcO73grD3N+gDBlylTg7kjny/sKomceLtGy0+vnCe6HQv40WmIu9/vR
3BOAIELWkVPEaTZseWyV8UAZGm1+zBpt/QADtk+lgSQ5yZ5WQPkFObOqx9DfGi0w
ZTglo2YNGnZtQOMa0C1QNSQeh2Gyld5UlCcg7CZNMFUHEJfbx70Gph6+t1kSvPxU
23uwWo+ZPrh8w+YJO4tjwHyQ8qVWyVo2FOgm27t62rzeLCMvZmK0dz62QuE74jjE
lTnvyLoxEQE6bG6Y409uCPH51fWjkVDs5Rqowc1lDMS9DbkmUgI6i+AEfnIcUvOe
33PO22Yb1c8W8M7BbOesGFpC7IQf5o24+2OLlhM7o0KfKng6bEg80//IIMrUJhVl
xkX5zB8HvoSbvsx5cjZqLNfRgULZH+yvq1BCD3Mgmj0k0ySYj7IWNC7SmiezsxWT
qy6w5gmI6iNoBo2M4rcYKwtKBkgA59PNgpijL+M2NkXHRJm3W4tuAZE6A+4BWfNO
O25cSyBgu1WeKZccqMqGTaOpYyV/TjT6rKGfphQsA9C56Bx+7KbelrDkXlkfRT8p
ofh4XBSvaAK2UVeMPcwrdbjX/Cts+9f5In/7bpKw4t5D/3HC7j42HlqPXsRiXdEK
d7x4e55oGyyDpqbMoDRvH8Ty2o/Z6bHUziu/Q2kvbczol7kV0+iB8HUQ5AmSm4JW
xAx8Ow6mg0tTtZZrNfinE9CGno7M/IUOq/Iyl16jPkdeeSwA+Zwgux/4764mms8D
gDPMVL6jQ/ctHU6bvQjtRgBFayGjz+lT6yV9cZ3k/pmT8WwlE6rpVnFLvc+Km41n
vyWhNrzJf7CkaG20RJOhe1U2aHjhhGEI5K4Nj7trondk9sQSvtqoCd6aInPeJgNV
jkBZ8LVOI74HHnJ2zOHLZH/5TkAFyqT7GJDIfWpFNrBSAbmUZFHkn9mISY14BI07
JhMvzSdFF+KP8VqqUqlTNq6sBgbVSjYRbupM8Paod9D9cDKTALY7ezrlORzKUMk0
mRmteA2dy+NY4uPB2HOM0xVptlg6Xh3zhISt+6LXnT6f14yZtTU5/Cyb5VHjJQgP
wsE35TmTB+weZJ0ha3nNvRidV4EjRu96+gMO4D8feEe+5RX6RPNc6/DP5zjdHIKz
o6uBgVug1ZYD9a8jXlZET+Mq4gox7wUZnrwHBzQDF3nTEEAWZoSQ5LVFNBL80jEo
lOYeV3ypWs/begGY+my+ZlajrDYJtvUWCmJglTa5j419sqUzaD+M5JLvi+piG1wK
7EahCwEYuaq/WKvTQKAGftMvw+obz8oBgCu8jXe1xz2YAfnzJRoO2p2J2/+fFZKr
6tNV7XmHqaXuvF1CN1hXXQKZe1GT/h4FouUnS8DjHRgNzseBrOQn+su9q/ep63NY
wkUKvPjLkBWx3oI99+iUVtSVVm/5o2klywKrVRG3XlmATnhLZQDPuwV3xEJA/5Nu
fGZB5rh/s/ksBOLpaSik4H4myRnDUCllSKUO5q4JxV0H2u+/fmtWEf+/JZ+5DZct
qTRoxV3lLeguVqyfwekyyk4g2T5/D2ZtQ5jY30KMoHDaAcUHVOnVl8YsdF+u58FO
lShRZXLG/tXsuE5KB5h02Cj0uV7TP+ucYr1nE8F64C3YwyfxWuzemYj7ve65S7PI
YfLPDMWOW6hY2QRPFYEhGvL67MRiNzeGc1BtbGa8ZnQDW7/Hv0Jry+TumD0J7KY7
4tYeGI2e1ZHnQ5egjz3of1K2WDj0CtoYHHZdgqNxKxXOwCpLPCgopX+CT1O2rmcO
HgXeTwnAjn0s+p4HRFqqXdCXCLX7YJOS3CFA+MAEkKFi9AqgAXS5/y7fdqhgrHRY
VRpyJOEDDZZa+YO54kcYOvUiDI1Q/OoJ0L8y8SMQyj+byRq/HlqlS2WDjKMRylxZ
iB9w5xvpvMrHNPaymd3PIKzRVwJENEeIsTB7lnUw1O5mCN5kzv5JGjx/rpSbvkQH
osPx10PyGx9rujGk6wVYOqtyuBOrGLoWeFmQ6cWjEwKUhgAXk4+nB8iFfj+IivTG
TmTxaqzd8H20laKpBCZmgme+5vrIpMyLCDQ1h39VqzG3gauIIMojTs6SAg79wS+v
nFYv4bf+aRIeFnbhMpOTyZu/4wGl/bUbu0OCvJKV1Gf25k6xtGNjoJb2h+feWI0E
AEU7MjeemGOXcICNskJPPvDwu/+/3on8e5hiQ3YRJK/yeL85BxFpFAtfJ3V18qiC
yviIYTey6Flri+eKaIPf+mt2hQgWNoPFYnx7w6d+8B5Bl3siRYJvd8xABbSfi8yq
lm5fU7F9q8na4QxemRQUzTgwpynAFEWBbzlZSKNzwWslE5aNYuUI2pWaieoqn98z
jUd+YcC24Psh4CTTVKeKM0G45NHGzQwGzN5suVdRftXsRlmtXzbdDNQrU+c10IlJ
YatbKNRmu3eA1mZqxj4NA70VkVrF40sqA5WtirKzN+sRkBteuwHg8WSUYgSItHTZ
R7/QEsEhEGk+Ji+mEAkdls4zHrHM9W0VyMfHWL8Slcsyrjqoeo62i00KSu7UY9Ay
GaMgYXaidt/WjyWWzzGVLSl2rK51lQrgqiw64o1X/TqI2q9q26HvKokp96lNet/P
rIu3rOmJlU9WFW0BMHK+E/ABJ6wjg2fCamGZW84KK080N42HIOQ7i7llxrF5cBx+
eBbF5zr5MoR/Ug5Di8ICIRitEokZUNu5eqAMQs4N4n66/sLP5eEuGh412izSnWmC
JIModP8/LuNP6Xj8irTFsHVl8u6rSsK1DU/LA7nzWnK5lfApr4wWZIUJzp9527yf
P6SY39r5NxLOdvl2yNUQjNbZA9aJnQzG4eqxohqH27r4piebkIr4CVdsuFXYaWqN
6o9UlGdYnGfPm+OIM2ZsorGWWf0IAY7NAl29QjmRV/LYo8XmomzlXyMYByS71rSo
LHpCTpLEI2rtQbAIyjWsTq7Uk7kJF3Fj82H/mpVEl5q4TdnBg/iQK4KGNWjLdY3Y
OBO50aGHMeGzyJmbB4AhE/TQeU+rngl04wK9pS9PJp/S+7/0DX1Gcn6hQiumTJqE
rzb3DeSg0U4VV44BUaJ7fioW8/cvHdIvbNZK9pfbTBBJpMiimcGeASEir6boUvRs
Ne0FzzVGVt33uNarhf0mYZ1IpbeaLIra0X7XMyoIygm+JN646r6VE4BlNnBQhtI0
L8D7WYQM9Ov8QgYrXge2kujWXEmIfkIJLCJ22g1TliR7d/DxhccxLXzGGG2lJUHB
kQy4eLMGupYKBsJIwtBN9gek9H5W3Uler8SMf+p40g4FKw4dn5wnRtZcVHXu3Vhl
nZVFUiNx4R7qy9UPw1Zq436cedS1MnXJl47Ie170oHhrm7i2IrjU9JT3H99Rt+o7
YphrxFeqse1tYd2aXUWsRyME/2mZU+hJCFZjI2G8C1PCCTiB5fAcmqapDjEkZvnw
IaFdqkTaVN8+TgZ9EAbHPOblRguDgPYHfOGdpuuzJQzGf/PE5hxKgYFVjGzyBbaC
SxdStF/kbc5qx+IDKK8eu9oT+a9yJnGEKnT/hoinR4eGUFvt/lHrlkNBs25rIhKF
cgY0L/p+H0fONc1TWpKbiYFgH4PT/6rWUhIZ01dZLV7t1v/orARdCkuQTbACf73x
SuIBUr9q8KEUlM2Va3rVMaEHuXPfB9USezNZlnet9hSk3R5hC5M4wcSHmnLSTGVv
z2jFRmdp+kMNS6tRDaajNu5KKZPciM9q6tEC5jneYQMPJBjHbmOW45zpezy6K3Ll
tov3i99pH9zOqoYWCsrcRArbB/ALxCWTicQfbS+rSGFxO6iRfoboWusTfNjN+Qau
deJHtF9OpQFWFPH7wwYvJnASMgXVjifMdtHLeVCbWbh+waEZKy4hNBYjCwBeDC6M
cv9XK3a2oLN1fjSQ4KaPM5ay9knH/o7P0wmJ8gI7PYOUSxt55VI96kHgofRKBKLy
6BR6FrQw1uQEhbhSyWi92gkWW7WacTilNAt9+ulRWSY8FxpLXLVLsyP1R76JSnGI
2XXMEEg0v/wj5s/cDYV99Qx0gVtJ0ASKNAtZDZGpyDwwE3Osp88loyHwNteaflx0
umMQ7bT3BB2xe7XCuno3HNg5a/feTt6MNWLSZmNd1IBJdbDBVw/HNYRF9hav+Otb
wJU2PiMQphfpJqpNqIWjlNmXUjNASv5hS1j1K55fF2fwJ0+RYqVE3EwVS4XuAYjm
eq+DJbktj81L9OGqEhi112LpMu9JK1z3gxGfz+1QSU4HiJNeN66Pm6f83Mlf5eOD
m5p7y7TKGNrcROJGAK2DPaQ4MUvV8Lu+IiFjdk5qNu8G7PmXCrqjXVgl7hOzc0M6
r2Pos1V+09hGmFojrZ5SIfAxS5j2Fytd4PHUA2/+dYNz6S+E8HrCDpky/kftjklT
9141JbzYTchHGWhpSgxnIU6TYfAWlmk7jG1RYdnR8lIHwUuDfrNtUWD/k9C2wtSS
ci8ioGCgAVbyX7h+rsa0WF5iQF0NMeO7bvVO7Bk2aPv8tMzRma2z9jnZiRDtUEKt
JdjgPQAPO/cQ3TZJwe9uVGbu4hfFdlBs/n8g9z1zDaEAU+HTmeB3rl29lT2lnvQ3
hRzPIj9j86otSA0DX6NDciMOR8HUO3vtFbaWzQHh7SRJBZS5xjINwSBsdJtFMFQT
4aTJP1Q/OmBq87n2QYiJFngLbu5M0rvO5AVIl+Ph9VVjmWbTKS7GoQqdV5MIXJL0
1xauJ3mt7pLRnA5GKtyae5lMHWKENC4LmL6SC84Ur0Yd4gKuMdW8eod2ANwszG58
v5AMDQEoYTVtp9gfe1Eoxge/7ZJu1Cs5uQ54L7tNLxw5hqnmyTc325LVjCk7lOg/
ET4UTqAry8c9xt4/Z+7Bh3ObvMK0uc7m7GKc/gznQtr4v59sormYYbTjHo2gDY21
609+yFDtG09Gcvp4I0OVHeAtuK1ioUbHlY9fQw0j8dwQWk3Es/cyKa35HUp7ciez
/9k0ogXNANuO79WyZqGmx4PFeMBpR3/gTR7oql9rUf3dCquQodlB9NjRlho8LpaI
9qtSmwj47O8nA4d6CmJ1A9B9yrVmPzq8BHRSygZNMstJt7BNzQQrz7oCAo2ofJAc
4DLS/ii4Y4zIQMdPVcXqSwJ+7eahlBwmQbT8NikNL4bCjpf8Px8hVXwj4Cs0M2py
3uAEFrF8B2HdNFkwmDdYMPXt1THf68IYxqJm+dW/L2VoiZtf6P3BTf/LH1QPs9gl
FH/S2q2mYVAX7MuHGEsjOEOt1dmUhHrWmQG2DLCJKRBF935plRB17b/q3++ZXRgV
JljBaR6SKc4vFBCL1oZNrrMv7F4k0NeunyX8QjDrifuKNi/rrCmizMtRT0pbiD9s
aS1wJv6Nz3bG0ViK254GqCyOxR+JKZKQLtkkX+nBpR0cSAGLrG/Uba6d0WrzqXEB
MBwfv6h6jreyJ5M4Mjo2ZGQcwtNOgJsORm95MFzpFwziyuJicRQCWcpeKojBEofX
dgPf0HrqnMj7V3DGSLWly7NWjfCfLmBFqeCOAqzog6Zpzwhb96I7Uz3+xu3EZmoP
GUelAJAU0k3grL+5XhdCaZWw8sJB6tA4vKlqwhSALpknG/IWoeNuxbyWeIHGL4PL
eJRxIcyUjrZSYoX+T/kmtMjuaG8sQaUIvdETv0jycXZft0zFEyL1zpDRDshaw88v
gdpr8g0twrtmkc15EW4MG75Jg+iQ4nDcREgOd5F2CAVqBwpQGPhw7EtZDE1uz9RS
OdDA2A9MHfdb/AlKpMA8HNjaByP2+gtUlvm04Kiy2l+jZLLSqwEtEd+knmZoHfuW
zdOZIciqhOEeYzYy4fLwIGz7KqAGlFzyFuniQX3xhz9ZBKT20czoUgkUJT0axG0V
VQB0OooOvZx70MZd+nIiQcmGta444YofCiDg2ej8Yo1ACjkDupnRFx2qXK7C9Zda
VMoKNkKeKMAzMMpm+n+tINXFlH7ePAkYLSBBnX0Kz4gOIVHf84SgZ7CFT9T6bgWq
sbVwKHAi3xaVxFdMp4xUx6X2CqWuRXrKnSqaqfQQD2M4zObmW680HGslslxLLQfD
7CIuXEDX/JxSTsbdczMev5SrXUadw4DQtm3xDiHvOJ/U+CJQbx4bwWAtu0CsVVBI
rG4SNA8wz9f1ONYbqaY1KAPHGUHITOzMzs9iWBU0ixMpcsf4jFCEuWAbErzeKmAH
2Mnx9LK3tv+zR973rFj2dT41xn7VC5N4z2nVUlLuOMDHTnUmB++JkcM5BPoPn4+9
8sr4I1QgUTLtQR4749gF3LuXhA2jWoGgYTXKTaz2WhV8Uz/mBDpepeuOx5GZogyA
SOFnWxLsK0iUmhn5U91THJQb4BbyPnpR2Xl594AwnwDq65w4plbk9ei4lnm0PeQ2
D6qPVM8NmBB3IlA2YGvPKTA0OawcZFNpvDtMl4EoL0dO1MwrJDpPmQ3udEubayvm
4xWO9UOMrk83yek2xUTgENl59agmzhrDRcQtcEvk1YJmGwVR2Pro2etiqbY06Bs5
YkG8at/HYGd3yt/w6ol8Gb6nPzzk96aEaQ6EMhBBbP7gupvsFTQBaBq1P+W/MuRv
uzsGGV/UYYGqZn3pH6/yNgItQMZVMWjRTJWy1DyuLfW2au1vnkPG2Q0K4jGy/n1w
aDcFGX2EZbr3jWRArK9pQZ7suRZlRTyDkJxPs5ifrbV2YyKN2VfdI9s3mA528sKe
jd7tJNRR/79Z4EYXm2yScOK1iolMFtAt9+yrtuQE7AdPd/Q+UbHOjUvPFckvckg2
4Fi5hI04Iw/aSZQ3cuJi0VMxIJW61kDks4UAeoq3VWaw8yA7zbxHMjCXkQXd0rm9
inWIjeYeKFT6lXHrXHlPXTqSZ6ckI8ZOykV/hyrZimIL2ZK1kAdXjMeLtStkd8L2
7XR9AubWxr+YOVcITMTK8i5SIX2JboKkG0Ce7yR2mx5/om3ycWZRYgJcWgK4gip6
c1POSEbiRLdf3q+hvr+R+D9ch7Ghp64NoswOefuxLUKDcLucedC6e4bkodS6rcyK
1S00tsNmNS2BvC3H1y8Ary81QSdieg2vXXDWB4AiAKonAYfqxlu1yduUCGurQv0J
3fJpIlgzIm85wZknwvZmq8IxbdW2U+KSEcN3rxqez5VKCaTsdHWYeLeQt3ztamX2
xYPmVXFknwsmP0Qn2MtRLII24TzYo9IhhsxTrd/yi2N59OnYnszEK4dOTZ4Ex6bz
sj1wAJZuIutJW+OHn2MJN7yyAzP51my67XHtZvaoFOVdpL2xE6vzwm9csvrSNHHm
eWuMkWDkxHqWqEdmIo1IJ+aFQr6S8B/4k6mo6WHkGjkphXiM3iGsGzyJqlTl+BM7
TpCw6111e3IHG0h/jAOOa+sSXnaZnKhbrz/gVQrvz0qcjAq1X3uX1YrWV1KoVg7J
5PA8mrQ4cFmWCe/l/Guc9CTQHHKplBQH/aBYmIcNCCugZujpky18++I4YuKFSeRQ
xQ3bZt0yVIOLjQpr/qSaCZnqPe8ics2+jAwutOpbqi28jl5Y5oYRNKXkwJHBpFkN
XQKOizR3jNggeWyg/RILZx+r2pJuDcODFV0K0Xnpefo6kwXAiHa6xRXdohhDchup
RBiJSSZAjhCbC+S1K/UsOuRo7GBu7iUjR+nQCK+Mc8o4nwFPxOrqPJr5HtmmoWbJ
dpPAY1G58pN/+Co0nll3uDGUE4g2HQacRx7fI33XbnheGLB/SifiGubocSkS8u5Y
/E4lYrguoDoSEX79JHYaAP43ra53yfVKAwJ8KkMK82c8msna+m6gJRkjDV9X0t3M
sbT8jkmPqgma3zHVAJEg8Lx8WiAnkvsbkxaCNkaxncr2+43a8XN88wbqfF8hHhln
O+gsoNnj/ylgscCvtvjONhcSpgUPrRE3pxGEJZzP58lbEckgUoQscEdpIW0zsRcH
hI0QwB/Ha2hKcXKatwcKiJe1ZtpFUnYzCZ4IM0jwVRJt6GCYqUq8ol8PYEtKOdG9
XMTWVg0KM3+emx9JoTimL7Z1YGuQI2CwkUDmtK2+8MFpEX2lWKer6ERP52CObP47
dYbK/JSERY7YsMZGTCAZ2Bz07BVVudRVJokXnRz6D5xIeK/dE2dNknN7K64SXnEj
L53gDqffL5EwkbrGEbR7nRgWVdJuTzpd4WeadQjGhupth5MGJhS2hJ/MmlvDwQkg
WR09yHWy7SIBoar/ciqR7Zm625Ff6wFVSrVTx1j7Fj4JSbkOt12uobgwxKmATb1p
2JKYvRQUFD9SIP3XgxMGme0ubgMCky7khjGoi5EuS1vC0SNaSJ4nAa1WpT9FLeJe
k9WaNJJd6sJx6G6jQ0m4/aIfl6uHwL0axpAB+fWqAZrQIfzQjVsvd7UGd+nXNMoC
r9hAAF9wzXTlxGLyvGjQ3OBKnRTMn4jdeKUliYO00Q25VFKl3PzPLaUsuH4egc1B
nGHHGCV0Flw11EWPSArmeFL5AUU3ujWhk14Sr85jnU4vc+cqt2rR2V1VHb9o96Tl
tlI9vAGEUkK8QpF66b6ElCd3T2Qeppvkd7ioWObrA7kMYhgi3S6jEkBIrTSFmi3C
ngXdC6d7HmVB2gCu4AWk189FyvqlGhijRUdfWajs8aQ6RsDEs+mN8qU6uCbky0yM
MXIVVCmr4/iL4Z/X7dCWRFdgPEFgNhCshHs4I1LjaJuDznptNC2drBmLL0Ad8Guc
n/sK7i0+5My7SkeM5GDWpCZQqdcrpc7qOOUAlr32ds9/9zE71vk6rToOEPgs9ZPq
ztCMQjM656WdWxwtnEnMA+fMVvYEMuQxbJ8/eaFSPOvIrGQ4tgLOpTySGsQlBaQp
a3zst3Wbf4M2aUFBdT7iaQULM5S9RHC8cwjUu+KUwSQol0ntVl7Sx9SC4ouBajoQ
pBQL0xPFnYqbC0ntnBOX/Dgd0el4sm+4VqTQnhxB5eHjyc15OqDnWg6ZzIdksnQr
sn8Mw3priZDS6s+//JC0RqQOfN3b4ZZkAEtADQxkhO1J9jb7HOboHin3ATzfYE4J
nrNQRf55y9VU60R2P5yZtyjp4xOpaHCJEGVTWxnvvqkG0Zy4xX2r9aeatMYcfgr4
eIbrzN3W14hmzXOhxvE5My7Uvg9I3bKECdxeNcP+MynipxyG+zHYRtJhipWI999v
lXjP4o6jQFc38or93lLo4zO5Ssa1VuGjoC8w84shSyOYJoXyhKdf2qrJyrtKw+1R
170Omy6RMuX8PQ8OpJWrI4X8oYk9OEoIb8muKUdrNYLnAxJIrdvfwX9QqijybAvx
TqFKenWQWmzTZMFZgN5kn065+sV7vVLbToUCFI1Nct9HEyXX1DivZx5eDe3XtKUn
Il2Cce6/8FqF63U+vLzUQA2udx9F0fIyfg4mQtYh+iM7J0c4vZUIsAUEYXkhp9XV
vbO/zi7M+k67jmIJDT+Nml3us0Djcw/0CXT4A44qxy3JTtZjm43PBLXY4GY3FWsQ
m0IAwixSsuqPFWnNnJmGBiA0daAcT7kjXBckqTlK7D9QjXoBq+uKo1v9GMwBB1yx
tFNHCF3PB5lea9dtU3v9TDo6XvLMaiuhuUMjs0w5ayjioQmD6G7YJEMNAyhmbIWt
4wQBlYkuB8A3790W37RcUKEtqLyMq50kdCnV5gL7FBr9OyVwVJuO123687H89xqA
q/uh6CQvPlVNC5Uqir6Iyc89C8dyNx0Je+wnR8fcxjHjdRxzI0Zp26i6Bd5D2ckM
9A9xIRK4S9+5YnI1KCRW2/e/V3gWUATS4OFNwwcOllFceIem+EvDKASYHReQFoXQ
chGbVtyxr8JIbNhXZ5Qry8tXyR2cexHEiftFbyABE2MGZ8MbLuJsbWamP4NXf71x
aUPQYxdj/LlIZsCG4VGH8q3JDpKbGOl46S2nYd0vikdL8iSA0tFxuFxmnz7IQfIH
W3Swev7mm+ZD18Mm22hBA9IzEoP2dyuOGwe0OCxHGDYmoi9FTQgPjNUUz0AL38bL
sMHBcvo6j9ekwIOLAtKzsb9JYgNM+kXTgb2XQheCat1ssx6bJNd2VD32TO511Hze
nVUz01dNRhTpLANQmLIIbtZ+qBKH1/wiVMxfoWPRPf5NNpDU/5qGcdWWUV8gZzRa
DZlfj3/VpNVlIGY/mTXY35scPqYtKB1EfAzJKQ+Kh3T8fwDs4eTT3CwoI8kEJpAN
8RyXal+6pXmZSykL/Zdi8JPJgkJhe2JJnif720iDx3I0UWS3xhDe5mRh0r6jadM3
EhCw5hNyvf1plh7ARqkgsN//LKWgJNXFTZB0vL+92K32//cQ9IU2VhhvHADk95bN
avlZgeOfVUJemhCMiKvPysjN3D/M6GKN7P14HSkGUrDXnWLoURCtjcrexwchqfQv
G56gxcZZ7S5V3Xkqb8Ers6Yy20hHBnqExNXxnm2SSF9L0cZv1fO/jQp1MXXIemAd
xeZLWTkhfgPtnEKCxgKdgthqpgYxn5Cp06iikOmf6QUgZLRyDg74Xic0T3jtoDiC
z6xanEOEKVnL3ga9W9gpyEV45+EvG76uJMA19j6tkTzEdT+ZgqTDWs31MhUxZzHP
kX6KNBpysz5dYY5GzkYd9G//XechFVloGH5A5vtM99qBspKMfNDbKxAy175qpWGS
jR9uMNkZxJjLKyZR1Zxw2X1jYaRiRjWuiItDnWfAVttw0TSeq+N0dH0LZVaBCPvE
Omvk2FNbYDVtjhZ5ds9nVa2uufuYns1YCa8rFttgsHtpaOOYjiqXiP1tJ/JGWB0j
Z7ORfU0XjerkEARJDJFhnEVwjr3V18+0FHgCwKo5g0Cn8n6EKVoPhPbE+1T+/MQd
VDnCWyoymL5+3iSE3f5U7sIsYtE8DKXxDhCWA0LFVCqMpl0g45Tx4pZN2KQqt6L4
V1EdzN7kQ/GR3Gdb7aT7YzwwTUWPALHKKdKdgeiCMsoFJg0uQYIOUjAb5xdsuBER
iVHqsolzaLw3A7K4Io5nrgyKGSI/vWu3SFCm+rmYJVtT90alxZovbmFVKMD54FWT
7AwpgK34wR4Kq9vT0Zuzr2YmaUQ0PwxjgTbxagul+SlWkLYItQi7xAuM/bHd7DHr
COtG2x7RZgbl2hFTc3jiXS3Q7wFjhfra1StmbQ1ElmTzb1PRtimYX2A19EnQJ2QJ
clMvCcF9DBKlHDcH50OcRkSCs0kxBeGEF7YTBp5tENRgRA6ykZnO7NBvvWaVtEml
cwmFQuY/7f/OpuJzaRVZSYWSmevSedTmgCopo2lo67yDRdAyWotNs3kBHfzuU8Oy
2KJ+VvuC/Yod9J2Fbs+Hu0egMx5SGTjflbYBPAdEpPQC6cs5mvkSzPttYgDGi0WY
O1RdPZFlYZBeVtLzVu7FUcb+rwiPz3l5oZfuSYonewVe/l8KqO8gRW0SI7jCyn3B
SfsUyDrT7MFRkuLyr/8qWhiGZ9qY3p0QZ6ZEc5ilnlWRtNKG++w9DMQE3n46IiNW
aZJIL2nr719D4EXXk8bKASkulG038SAwrV6Yk0HhyaTuX0sHXClVuYqm/SFIyG2k
yTRA26QcG9R+uSmjvIUkAjtOg/2fNIIL1Q71gFfMAhpNd+PWXrPxrMS3pcpasZq2
tvGXCNsQs/k6UDOow8GY5BUxtcxpfwHGuCj75TAxbuQlUsuxU9r6MrsdXJc146NM
xPrBXZ1CaPVTM+/9b35wry4tDUXkMb2Uu3G61V7+sNeiKcjeWzVKheYVjejMZG9w
Aawe0Tx7ZEYOOqf7XQzevSbNhGSpDQzHWjd2KXnQ1rOArbGFJr35sCEhH4/FjwZI
GaUcmzHqXj+EkBwVrCmpbPeOU3OVT2K3C9XcwEBOhUM2kyu/ztDb288HE5qNYhH+
vd5CQ706uVQH8WqszlxZpZe0Ocnj8ix9r40Px9Wp2OWQiNa1CG0b9tX0ILmsic0Z
NLxuzHr0/mZzlH7EjS3D6swvh6Y2hXKViZotIxJ59nXLyGg4dnBosyDaj/IIfgUQ
orXtAlOusnfF0E+c8723lKjwY5CfMo1ZTdKzPSHpWKpwPg2BI32gfsXUcnXWrKVE
sFT8XWpkKex3p4IEgtLfYr5VOLf53m5N/f++QHVhOsco/d9Nq8QKsdBldciKMRV5
hu7jsYLi1lCrTQ351Nf04inteUQvQscveONjAQ7uPF3njiOQOVn+rnBIjhiYQn5q
YurTl2gIL5k8nYny3SAjXxanlwkNt6xyV2i7WFyE4cwo9+7AkKmlX7itTjfNQc1P
q2yROuokS+6JzSe5IV3qgMOHEsrPAtrM+TAMrE+r67Md1/z6rFwVkxgi/gWRUcS3
DOx53sI6SWEpMxV52FGEPBXhstFQuR2yoB4JoYiL/56fvVl3xNxJ6f0eATykWtDr
AY+Qk9j9OuADCCjnxF4wgFB+sREyFJrcnA/U2kVhSX4ZP6C5m9deMvnCX9ZzP7e2
8d/dP3vDkB5NpkqYtHKruU2EIXzrVJH8jKqZCwHXAWtF1Q4l8YkfFxY8ws/R46Y5
3KVc6Wf79fVpWEi9k4Wgh+25FHLW33Gn11dwsuK4m1IIgLR8du3fCwdf4YbCL2vw
SVmo5G1WajTwjfxrbVfGrpNQ+mLq8vOE3jc2Hsu24rKjVKnjuJeh5MthvEe+a0h1
7r4nyW/tWHLMf9fPaPz7/EDw8kyyeXSXs0I+pfUfiKQW2i8zqc1YK1xqDZH//PmT
21036PM+SsmTqUODHwW6TCMgHBUSVYk2pdvkxkG5t4mxeWNGWZtEiGPc/PaH7R6g
nHyybaFDOPXfXOHSiY1wFUQD9YvNnoLsSKcAQUGUn7uUeTHTEQDQzqHjG1+Og74v
edXBM0eJRoVffohi/TkUf3q9qV7QIrwnK0tGYrlb2gOFoqGYP9CQrCw3IkbJlB1J
TSHSIZ7BRtG1uqn6Noe4o5Rim3KelMpZ/x2b4/thvXkBa4Mes2vRgCxsNVJST3sI
W+K+Vr7O8ZV9C5Q9BV+25xO0cGqf38BuaSRSP/5hxYkFlsm+E8vWQv/klXTh58sp
0JGXDoM3zVvZK2iQBYGCBoL/saAr9XaRCTLjM2q5dEF5Y3ADQxv33TpU4WHpbWwx
7/Hcy27fokQhjFy6vn22h/P6VkMJQ5wC0LGGthR/Sf+530TkzuXG8+8eAZqVNCDq
yNtPddLY+ajEW6WJetct/z4ViqiKlirUWkWbM2OPo+yWAKLkf7/jGeafjELH1JLE
ju7cQ45edWbJTGFm5J8ROS4vtWvH5CB2YaUgelkFSRa+zzinxFzKgNBW/eR6zzoq
Cc6JltdglH8iqZrz0UmGgsni25e3XyTmfx0fy8CLEKINwT9GGnlpvrQ36kcdDrrG
XQJvhj4CM2se7JEwVT+PSRrt1UcR+ORtXca/f23KKUxyevdqbQKV6oUyuOnAo51O
vapVMkJ/7/MZw7lQqvEycGFqkvJSEnlM44yqDz2vpBO3HQf2QOlNrIijdg0Vap7q
0hxKuCKPP/PAIWea0fnH+NYxWiK0uZ7a7hnJWqY5je2jT8x53aIPfK8TZ8nOJ3x/
5CJ+2PrBLVs9yUCCKfgAF1WE+MAj5gufLKmiAG8mr9S6ZedHUNROrNMp27v9Ssdb
SHBMuOoi+OGuZrBQwvzZzvBMGrP3CYWAji5z5iEIu1lT756d19CQnlG2gFMcrukE
KX6/TgpiHa/+SLl9i1ye7qMqYMvvMUKKuYPWx1qsMCYNd1pm0GKvjwaESVg8E6O3
itUTZg8FeJZ7PO031dk+juFUgl3mkjgdxjK5d0CvgpIyxFy+VX411A4+K2Hhjqfg
w2p4pn/cOnjbox99+GYcMTbiyW5uCEoa0kIa4yV5eJg8RpimCs0tkveF2wehHDWC
7bGa2TDJcP+Nc4nQla6p8aDrLVWD8eep/l2EiZh8M8rmd4x02AAbbjc3enJBh7iq
ZsQTpCunZEhrdpB7Vpv1VFmZszxQv58SsjYqhoIfXWtL9Yz0nYUgnjjTyDHb2vWj
vhajwQNt07aaSjOMDsjY+q1unJYVd6z8xlDdaTF3tcpG72aypeu6Ps36miP3104x
7rttqtCrSSnM6U9utq7pB/nXur5gT4LErsYW4uXPatrf3M/JPut+XVmaLvrI1llS
AdrqPZpNmxiIc0cSPJeJA67x0hMGI7b3eK0bgev/IKFsrpAFMZBbvU8LOK+YyV43
BeQJWRqF091mQ1INnEPZSk5qkRkWx3Q6BWM72mqv8oXgtCvWXpTOhUJBkSMJWbg7
4eMASN3P2PFs/vGp62ha9qYiodsp4gtxX37KV/wehBBqMdu89H60Wd+y6SIxyxPl
4UzJOX13IPvPmrne4M1cWqpGntSyprbdy4Q0WIc2Zc0i9xhLkd/b7vGTg+h3luze
DZEHnPmssNjqhwlBdj/kT9rMK8U/BkhsvrAsOgvJ/Fzk84j3vL9unTpkKWtTZ33M
AaX+LK/g4vTPJP5dwJA/RblgRwNo3sGsXyMs/hLtcaNgzQo4TA8ON3Uw8opO/alt
f7PC/9dLhG/0nt0pIFTB8W6voQ53mj1aCY9UwoJV1Vy1Fka+pWA2qH6/0I50HGOs
CQtEsF7x3prHzhW8Gi55B/TZ7YkYk/qcSr1LIKj08VssHjRlYOAsMagxqaHEzzIP
EWbGgSzvb+w7zK8R1FWPJ16Wpm4tGoG+dqvzGrX71x01MiVwF1kityWbcHBFHx4j
KoDHN7MaKjwthXwlC4vR7Vq11s5/eTHcsM7W+3NQMOiytp5I+K4YVG7rHf7ElvQI
FfXjgVkIbR1gKo/ApGwZjvOPnO/59l6JnFUUnMwXb6jiE8PUnqmJP+um9uis/jhv
gzqRYmKXa1gaFafBDlVqIZHNMMaCiLjFHz8iXCJmw+v3eYCbfN2x9s7UtbFxSOok
E8SgA20gvr2M6t4nZ7uWrTuEMNv5EUL2muBEqqA7LNVxKO5yYaWUnxIVVbHNhoUe
IN0w8E7PNoaJMFd9TdNUQQoxZu00LTGHMJNXrA3T8Uav6nzSqf6xWJmVyYL9Wxxs
pKcdUUpspZNoqqyalS8VSO9mszQD+WCl2F4UXBW6uAvEEcjqqflDrEkuRH35Hpbc
dE68K7s38u/xHIf/dd03/2jYE6D0yoNWpjN4pR+pkfrozLzWRr4Pr+ALZG/YO5dv
ApWa3tr2hQRHvsq2T8Mj3k1uyClqH1O2z1jhHrxgIsaWP+lv3x6e2qCuLKtKslxM
ak0A5WQ3AnXmpouD7h2pPZEYMBP5S2mks7PZfdRAbMwi6coxWCO5D8OdwZxU9q5h
zG6pTef+75jFKadmXIMEaLs9BPfv68xcONs7XsHSN595rolQAyOGgt7bhiLsyRhb
3Kd8puA4NzpRZi37SURVP9QM2UeSrDB4lLkoT+cUxy/9GJkDF75MB274qul1X2u9
xTlFXIwqo8MEYDYxoWM+PWWe45AExGT+BPIOnUbLOrLlVn2WqndoHHngKvaAmArK
ENJw2oGzJfn309Wjxp5ps87SEt3UfWcJje3FSeNwxPutnCOwanF2qN0eaisItyUp
yUmTJ3+/wQH+rQ1l17mTG2/a1jdY1mBJtzmFtR6GOB/F79snL1ae3L8WmIQZIn0n
hA+cccPMW5gVy+a7V3HRilZ7TDf796pvgOy7C4XCLLdXEKEAax6qNGaOK9KCfVif
LpLw8/7B3iLYtA9SjmxNG0PlbDzpL96skpDBYDoYWrOBp10uBuuzoo5JLo6tZ5cj
tQuBq4SgnUqIdNsycl7aDqZczjC76tFWkTqmsHhAHR7PGgqKEcVPfyC6fvdD/sTJ
Em1v0iEO5gCPSu0PzUxc2oGzrqThlwcvTL5MoDXJwsOptvmzzZ4QMpoZKSO7Gka4
XMrgIifeXSIRHveQfNt6sAdEntsCHo6xLpQduDGIMaAFU3zSJ4aNovLQX6C6hs7f
sR9tJji1ewrp7G6YMvLQdiM1EDLdigfj4CpWE55en+WVLKAg2DZ0qj/KqKc/RUrS
REqwVycXc7+ohItKPFvhrf9ivscCd0BBRN7+yAINvIV9/lWKO9a53JNpPDvf2YIB
6qO8N8GrmBM4SLSow9ZgpVk4Hsbv42znq+QOuHkIztCalqHVQNHsBcjVC9gYhUJ4
+CYCrw9Y9JqoZJduZAaHUu/fVFBwCN5bAOAvTbe9M5VwqC9wSy/AKUaXZR1a+x1i
rvizxjdUc3J5coZYX0+v2NyylCMe2jLnlIbM3b4HODyFDcgoWPIplFnyVkwmqcpy
Kz9JEYh4hEvq2j5oxwCZRDIMq3MHYNEr6BU3KXb7fNsuA5Tyf77KOywvp4xOzZPL
wfXoAowvwh50YlD121CfZmmARDHV4ALfqIxdtb5fUTBZYsqA7z1XmrrT9rXv/Qu9
Htu2db6rMBDhYICi3P3suezw2fAmPz8Yao2ctRxPNdQM3+LaexJqynTftVySy53y
E/hYQb3bhX4ni5TTbfjJt6jCz+azHhcCVoSiC5TEJpszGKBy6set+wp23eCoQmLj
eqTd+9YsmlxRvXaA2cpSu0s0DejK+B2az2TLLiVoxWxnlwvVT7xiC85E+xCzfMXv
hWu5vM3bHPEayeDAN1Bm5cPOV25qzgZtHOl8Czg+fU00GxBU4H1aOukNWbLWOgyV
ag8vccZbxQARzBC2Un5WPDNDXND0C4Y5RwNGywuOhA9l6ySCl0lJZKBvsiYinV+o
crqIax6WATJSAuEF1v+wQjVUfx5FMHWCUlvtdJ1GlGUjcNfgCCFWwfXhM4KNYiGX
zoMCL1TBreGrT+3m1DF1XpdkLxrJJ7IkrLzEjq15YnU+z9CxMobaRiC+X0TyvJj6
CqXXsX5QHYFJpl60vPxLsLoEsuAxUACQ9uZ4ohlGAHBxvaJhYsk40VIxt2MxSrxA
SIleW737cjz0nZAc4jcY3X6k2W2Z0SHq6HrXqQCzyYRuSirXLlJnFU/rblEXmPy8
5QRcdmIS+qxl4UDiXt5+fPGJjsdgz6q0KXug7Ds8fXIy0EsrkRFE4AhcUYWPnx+/
xF6Q7fExMYngWIV4aVeg+6+PSKQKHnAKQQLuZ23UHrix6nX3X8Ip2Shv+jhwil2J
yGx5EuHh7IHdGEFJXWLrdi3443F16NL71CBKMX31jdxEhCKokRNEMgQouFFjQTU/
jvaGBvEPsOmTv27AXoPmJworny9UM4blLPFzS2vUKERaJm7wel3ZUtMeR+EvgTjU
Gim2ycMIBzxE0rrLyXgH9G9mLUrxAHzgiKC5tZ8BGAEw77OBHmC3OfvHnZ+5yPr+
xUS0xbc4e1lZUwQjMh/G8atW2MOVTeY/Ez6u5+Av64nk/hCrSufx2EyN0TBVGKEY
5bUf4vmrf0hCL0kkzK5jd/RGNDUE9By0Vzfp0AKwvN4vQfF3B/TMazC0eESziZm6
iYiymv25Sl1hZGihpalmzKBfuSfzVTzYGjxAF6uZlrelcr0tJvDF6t5Uxx9MyhzY
0it7hXfKLBmEGJ9W5l5S+1LZPmHOwQVIC4emGxbZQuOkwudvHOTMTrW1HsMEVyQ+
bPSRIZXX+N2m/is1AorRmTk1D1Ooa/8wXzRmBwopyy6mwjkaRdKonERacQpj5CSZ
dBlT3EhvGEps7p/KXsE+jzPjsi4BdWluNDuzTtzMxjprkV1Xmu5bmLKt0tTdKf2E
ohvwvk4FSnLQlR1VWJE3yUHsMYmVraX/tCo7kQ7R3M1jug6eYp4iv83mUar5wITE
dfvZQRT0feydJVlblck2VfmYV4uVuea+AdaD8ApT4lUKw/a46VwKhHzvhiUPRuOc
LQPk6hzFgltuJ5sSXxqMIkq8jkbTJ57ewCQiNduP0CADmi13tngtoTgkybaj1DMX
n0/RZagb2FxenTc8u4IcNANU/0O6/H4LB5jfL8Mqq0e0FOW9dpdNAM+AUDi/Jnp/
Hh0pTBwk7xWDkQYferxJcXo+wQgJFCZ3BtlghwDc9K5wtGIae9kQOKV1CPcQtbqx
qP3nO+dXdwCxyKotnVdC6wn+hFwYgAVhuSxjpTBLa9FbB8PeyP5hEvGisemc4UY0
Z5XCfSEje6/uDorS66laMU6kyedo8ngs/sz4VU/AqjPCLdtX/qoHAr/rs1o/dah+
+MM/txvEPIAu6Go/ynq3sl3RprEME12Y4XCi8axstO7VxEnXh3Z2ETwEpOyGJz0a
yBRYN778Sz3G25C1/gmpJUrltuLieS8P+cC3M/sawtc/edlu0fPbDivVKdXFxbLY
+EZFA+eTe45t/6aEE9S+OFWXwuEp8t4a2nyCwpxMoRDpUAGnas7bR4QD2vAGqS9c
CdrEpsSmwSe2zxhOHPnOaSiI4PsOr2w1s2OTJ4W06N9SmdYrQDjJqLww+k0AB7Fn
oKe4MIcRyE7/wH/5o/AqlXYk+SfQv9tNWwtGvyfs2d1L/641OK1YZrxgU1hDVgad
ysiCVdQGsVWMQ3ciCBh5SN8QhLqBrYGp6LZbXL7vJdlDPbN6xFU0xQIN351ImPb3
/mFkaJ2o8r/alBGuUXx1LJN0XBEosA5rd1O+SgnMeJSgxaLacE3BGVW6pFYMFdpO
IbFp1CdIJB13vc2tKmXCDCdTby9tVXPOu0ulji0084rRQfi2zxulN1/OAd7jpaui
WamB9d+dZCI8He2edVkfXoYx0JNkXZ+932AASYjFA7WGMCJtUgWr3GIo9IZe1dY/
tj0JeIT5BsWtxipJUS1hd0abaRxbhvNmLmLsVFkmUMAdwara3DZq80Yk4S0vIYva
vnY3tRbspN7OylzvUZQJSg5cYWAsSSEsiXlC93IhmG03c5JHhyME9AyPtgpS0oC+
lJrKsqLQgUtAmkKTMdrdJR3Pgw8kcQaBfPxr2tMfIs45rBWaSko80kk2Lc6RzNVM
VWR7GeF5YodZfiGIZ9qXfnDBVN2B7LdVTKR+grozUKFm/XYWAnrAql/6JG7beXUO
Enl1TsMzFAVhr+9qb3cOiAXHNRfuUuj0cWSRL9TU+8EiLIZ/FRpzGND8ilVwsF0P
71K4fd9ameDRvEpD9i5VECVWcwiFMpqckrBTlOkE3GLAYg3L5l39grQZoLdlmi3G
iRK09i4if24O32Evth64T0J8wK9L0Czx1UnNG0PzrG/GU9NAy0QWa1YxaQzMPWRh
n8dKinWtuo53Vgv+gHJc+DcdUn+vVJoaQYB/dNzDll2BqAxpEQo5+BICN278kLJm
QsJvZ6vVEFhQgqV2k9PycItl/njWMpRArTyIz8szC45QP6D5Imn3iDjLi4xW+Tk2
oojfFj9GR3ijj8pZpU5Ko0CChhGPpxIKk7xUXHoa6cIViZayYB432OL+rIyGyI6m
a6TnX+vkDNO4QM7swpxJi5i1/nhKBjDtOE60ese4htKZlXVut32T1eyHOds0Qx5P
2t6FaREgNGCLIctfNmYxAl/jtKTH/h+8XaCReKuZDqOuP97owppo8dwv3Xv0sms8
0LVAOIlQEm2X1ZnRJewshCTZWJQmeJzYC2w2vlunGo9FO75+aoSS5BeVez0PxupW
sZjEuxowewdjs1PEw2CM1/MR3tpTDREUxlywQU4yJclf3lu9XPGdnP0ZBqoRodPW
2DBOaT5gWpZOSRBPNF8m5RK2bFx80tng1t8U2UbRPNgvNI/yrimVP+eug//qVvW0
U42TqYtxlaozjgol59gsy+Sv0gAZ0QhUTNOX5IR3x+rIZd7i8ECpNBmRLjm7SsVr
i1ceUJ1raDQdgb2dBFjwoKzSd+ke6u9Bd98VOdvfrc47deh3wWGfoNnZmaRTQZRO
I5sjizS1kqNac8BTQLQiKVcyFOPcWrBVqOewBTNa0ZWEV7EPVAkVBCUoih0ppVLW
4DbdiIoRYik91YOWU8VesxkZW53y+iyfzZ3VRu8/QzxnB/R5lyZcF9+uOrcuRuUj
LizdqquYc+pNg9YtCCUu9zq9g0Tw71e1cagHu4xQxtrWeEM1RemFR0Pch761m71K
keziqvOQuOCrD09Sy2rJB8DAb0hbOYfwkXItZgc4j5sHRnAYMJqfG/1nGWKRJqSB
igazNDqtT97Ef7TitZ3LkP9Vu6D40klDPFT4jGMf7akOZnbjM7/oDb5+u+OhR1/H
ymKdSqJlknMhvzLCjM2/S4esKVSkwGDGDd21iA8Ajy/e3SbYK3nSCClbJZ70eQyd
2GKaMZIGfNMDKAmPwSkBGLo/b70B8uotlQqs0tQXGbvhtbXXRCCz2CNROoF1VMSK
W2bRNUv5T74XDybEM1MqrmM/wB5CCjL6n3QkQWbFS6IM9rL/uuH6xoRUF2L3nXB1
HINpmnTEjEnMnPOzKJoCQInxQ8GUCrsCoRN89ULqhOtxgFwGZa43GBMb5atyYq+y
O/oLPY5khiu0C7d/sJK+e6aC2Q1mJvggravahcSJ+xFy/CKXjXOiY9+nN6Q9YqkQ
719TwGVNdK/qPLPZbRlp7qRzn8DszfSDYE7dfI8RDKWCZXnsfupoJA+I4whqksJe
EvC1QOnKO8uxZIwQOSjZWVH27O2i9IVerE9G61Sj1RfBh28k/8dTzCkROO6B6GLr
ZNbWyIHJRYS/y0FV5Pi5X/tKNDFKjXcsM2xGXI64ya3prScxW3PRXbcWSw9GRkQ1
i5xYfJ+ooPQe6gQL2OO7Jrk+laB+4ivO1f5qf87tUYW2Www6MfYDlx2T9yQNlYY+
9mgwrPWcO0grIzX+SwUNEN8tlY8oKklGPFmg69HmVqa6F8vTi7LHiYlF0CxUVhTa
uxMvmzogieD7WqzK02WMpa8VOtnncwfV3rDNsApSgsRUZr3Sh6kopE7jWJWKQfNP
RTtFvgzCNw+tELGOXJ0Z/OcVUIHtqLlzVSK29iRBhUwAmN8ER1jcRjUZvCWuG1J4
Rsc14PX4TVnWStbTO68FPiDEMXobdQMIznBRCJxysRGvj57OKhub0oS9qKMD132H
b5tZQP0nDFUEtQBz2InEHl3g1Bxv4uKiMUXjlAFPiE+nnpKZKvnqcjPC6KHtoTk+
8xkbyb/DIm/QeMWoF9UqKFnBttvIgznvtMJqN8rShg/rNmgFD6BLMcuBMhOR1DLz
fX8FJXSQT4CBuEVsXxzLOlYfwBC2mhoJED0HE1e/ZVA1mEg7nu8kf5SDkmbL6bla
Pw+pf4no58aAFPvt7/2oke9Swh0FfVpWl7ToyxoR7U3pAJi9G0Osaa3NHicPr7/I
1Sc0i1GnmIukzFhr+MwRogpCpPrhc7HrBU4SKhuBnmaiVrSGiYDYwWHH/r6kUM5t
tD4sWz43jchhTO49BOYMPuW8u6fgj5gVZRhs5uRgV6D+iedSUiXnbeXVNxTYaaM3
m2iRyuGLC6w7V4KRbytkZpzAyIkzFulAvarxY+W3SuoAUOVVBT0QQkhqAtuURaJB
N40QrM1CjtOeOVL4YldhPhgP8ViZPcDioXmp4Mt5OOdgp/WmmvEod0epJeFM/SRp
HXl6DHvidFsed1iGS3ZJs5jLSurIjtsECLyHH6vc7KO68jdlO/0KXk6pVPPYTEJ0
72A2ySP78Mc46O+IDVHikVasnLxl7odYa0jEa6foZYOuCiv5aR/YObC/+YF2NdBp
37NoIEakV8xFVXlQmvBiL8U25dtWalcc5Pz3vrU1XZraV+2k4St+VHhhboQ8dWo0
wyGrEjU7F+mRAN/AY49XmZdH2nVl2+1Y53g4aK5gx0WWAazlpha4L7ZO/DYu2YG/
3XrQToGAkhFkpmRLGpM76DSQmfKCK3/Xzb9lp7Iblv1CwmVR9h9cTXSbaALO/xhl
M0rWILLyba9aiWcKFbo/g5XGzMi3616Vk5fx6bNSv1jlX9d53slgWgmN8JpZUPmG
g/DkMmHRmJw4/7Q+6Jqk9Xbd623GBHM8QRJ8msQVqq02TK7rsWtkqsoOZxCRhuQO
FxdCxqMo0/cMrl7WNUnYoQ9T14foR33k+fUlI+z1q5/VwVEXrCuBZGGFFs3ck93L
Fnn6/wIhAWHqbiJlk1kvOp1g1Eh0OwRJxmTYooenAS/w04Evp7dcokrRkfMnlLhj
HVV3+dNAa6PgKRIeFNGh7UMqkkkn4mvCVAFwG/Wi9sF7qOWs9e1uGlD46FhW92Fg
MpU+PHLH0bYYIPrwuxmZTpS0e8WFitU8TYa1MrssUHyIYYjwcErX5O8j36EwuUHX
PdXrDcC84SZ+si9S11+RrGi8+i8TxcuYgV6SfDL2500IAqTR4Oly7x0hDUUXtiKy
mSWjcUAnJ6BFT82xA+CGqq5fQj9VNpUFdUNLJyGj7FfXS5P62Yhntah2ELg5SQJS
NbU/sB6r21xdisoHlUjd8U6JTyGADKuWdFUJdtoE5bp+XljkziuTrjTJFa11hTZw
tQ0Y0gtOU69h4xS71gmhfEmP90uXQ2Tca3Z5Bmd44LaFp8wlwG+ZGDa3dfBr8HwZ
O8WvM/BVXsuItRkd8UvmNhKrFHCJte63WfYoIFSpvhONECXiOCPo9Q+wB2GZy72C
yogCCL9FvuzBOOZyEFf19qq3UjNzbOPBOmnyIXzgL03eKAbS3GyQ7dVJy0TWN6Na
K8iMFUBCHfLyyMxDyH3yZBBOYjlj90A6yvERTM5vzHz9ReNQaSuoBCuLFO54lSrv
2aZoIXQMcmPi5bgzSphWGqp1gsB4/7ZVKUi06GGsYbrBuAlMHgLhW0+I/zcR9IOF
SzaXHgBNXb3pWSQX8cFKanx6WkqefsqyZILtckZQ7ukrnq9kjho5WhQnR2yVdgzX
+o4g/cGTW7Pw3f9ftLCQr+7Q5JidpUbV3wSkuW8aHwkp0q0YXgz2fnSxFvLFoIdL
tB9Er7C4ISGyzuPD7sBjyYt9OL5QBs8HPfbPeeK0sBDCtaE7jS5RXLmLcxCgicL9
a6G0wykxwQcw4OXbc+qYa8s1Zz3ogBNGZeVY71ovIxm82Tzj2MMT/RkNXG4C+LDd
5lLrW2K1tGsSOnFh8R5CAjZwSWMS0hmb20dOAkw8OIQGkEpPw4RLWqJBgvpcN7MT
QJ0ZVPE0NOqkAK+qqHAUs8GGf49M/1XsbWxgPLJUOCJ7YFYRaw8JQfZdLgyJb7wl
jJsSnLeL47OtwFDynxcYw8T/DYAKd5yicEsTmFDmbt9IzG3mU2pdRiCHmpoFNjNG
WgYHTtUfL+qbI4lWTP+T+erOCJA7EJmWLPGYQDnKZgnkWreUjmd4zniLiwjp6qFl
17HK5xWKGnEWO3p6eg6jI4zOaLlIiLvlrBUS6xtFB3lYerBskqP8eyVKGvtioVgP
nzzzL1LVIrfFJOaei6Mrk00F15+2Nb/INcz6/uE9fbqC53VV3U3iK+ufZulQArkA
4vaYS5AIobYjthnl1yuUBDYZJGGRisOe12cdtaIN1qwShPA6CiNTr12l8AEy+rbq
ddpIAmm9IyFIz2Z+jfcpwfw4TmbvUNYeXoB1S0u2JsgpGQuR9I7gC1ne/IX+sMMH
2zBlxuRU9KyQGyUy9oeRHrGCiOsYdzT11evYgUFpwaZYJaON+Sl+iViaGw2qGym3
IbUCBMQf8pdx/7qMyq5IPYHEkpHxXoxJAAuff1Fqs/r6J9u3JDk8+z5/yaO/KMan
rJuTJaRAf2LXnpX7LehqgZ3BKRLvrPi+Wq5QU7tPZl2AEfHdXiySKBZV2mKBfVrM
IB2ENIw7yAA4AlJOjWjPOtO3teJyysJchzzoFVwa3RmtBD+crcyrOTDk4aKqNPwD
v7M5/OoeF2+v2paWoCIG1E+35JzfQyVQoQ9jevwdNIpcwFI7qyXD8PKxXLgFIfCc
uKoWhkp6Hb8lLucOPD2/gUkbvBUl0KAgqmGKiIM5MngNUoZtb06U8E2YfWQbd837
eWHCWBLLmIKsxH33lWSSQdPP65GypCk1lO37pCsWEloAVdzeCjnbFXRfElUKOrmX
2mwUa6ebdp9R1tQmxPA3wh0EUlZj7he4b2Ga+9g5vt5Cl0cH/TCbCp4PIzl6foSC
Zh1xGFuZISdHvsNVSGKQjsctaCEuEf69AMnONYnVZQPPLUc3fvuiX8myA7uCR//8
q+Z7IyxZUdAMIMuUizqvS8yMopYfrN0enza16g3xr+GIccsoUQ09MRXEh8Foy8j+
f8QIsoR6P9/Yr2nmNCiJZDBPwWjIglNTBFsbi2UmZ1ynRWt6bMhRKpihHTyqx99h
yZypQH3kwlNuJNj6qDkV1lGRmTiGEtQH+2x1WSzxFsaXUyX0YvlPHoRJtyvcv+a1
nKZeXH3evhzPHyrPDgVC+gh6jRRsKwwA5RwFx5oN9PZ+B3+tOQHIx7Y9o94Wl2xl
WOCDA3ZLDwCq5//Ri/L1PJZD5g2FTx0SMgarrzyNOn1mtfygCnnom88VDd4HJIzB
deS8pEIOwSy+BqTPpQ8RbrOELZ7BA1etKBjK1/lgmB1hFEM0NtmfnctsrGYkny7Y
ehAEiws2v4Bi6Og2QpSKxXRVb0G+yPHZIFEkzd8CyU8UOBVFhhjywPbZkxINOqni
foBNPgGtaRm9xoC7fnaASg6dh+Mn3KI2ny8sNKED+XVqCIj+lA2xcxFJLIXqbUns
6NTCtRZy/kx6/Nf4IX7kI5qdegDD+9nX2Gbv7rEbj6Lmokrzx0VCBkWXH+/w2Bk+
Clx+ao6E7hojmzSfSJRbVN5Q6icuX7iACSSxKxnrqrQpR/y+Sv1b9cy5zk3Xuheq
yaArskMSIpEwOFNT3a+eBelOH1yjQ/0wlN65L03XYTG3T4RdNRZPW1LrfXmwd4+e
RQ5FZAMjd4SJQ6CNd9RWjZHAYuNXTeOwGqzXXJVJWvuO3+6RZOvosUYVkfg2KyS8
xDvr6CtzcEn2Np3REWtYacz/6eRNDuzvdI7jeg7/3+y8+x3SW53eYJ5RxY3HujaA
miEyxLu17V3RlNdIZIttBhX5ruEHVXl8JX/c7UhkQjE3f9Vf8rMcnPAXe5YkWxlI
R/0WSC/c1zje1/v/RZnTRqfXqKEslMzl751kjMxwGY7KXfs8JL86ELXWvyq+7x5T
1+5NW581qQsKaXNiQuDbRz302seFYp5TaKpw2Spn+yhPPgN47JkqFhOFy+pcAFpY
ZGtFGs6VWDgIggdl4t0VgS9l3Pn6I+PrCgCHNliGbZf7NeQCSarrCjd2YNwc7G5D
QFVEHxRiLdUb+2s4pk2IWlI9NS4BvQsJ3/iiE/h+DdwtwomIJFN1mJYsut89D7jQ
VKFmp2WVKIS0CHbH/naChPiYAKHV9GrJRpLJFp+D0H4SoLu70MnGPZCagz1maoNs
aCcUd3lYdYCtmBOQqpmsI6xTDRUhcd2h13srYN2q35WLHayGZaP2m4YjIj5Thimc
f1rIspab2qO+bCf5zjr4nRpS6+BBsD2+Vhl7pxBMwsEYlalqjlZJqa4qnvz0CXlM
mhRrQRRaEpd8VKaziOmln3UTz0bFiCnosAzKcdWpE2xDEclP85qA03firHK5J8yM
PxMHIGCpCk9hg5y3ajGQgL9gDrn7kAhh/SZs3/h5tol4zSc9bqB3DPp2Iawk2fst
6KmCiFa+d5uPdsOsGmyVnFM3+DjhyiyhXHaxtlyukWH3gwpEfvBvOEggs0TbNJxZ
lpBd4WUlZSaMvtCO9EDld4gxhvrsN8mcfSLRZ7jup7ulwbv3qN2Hw9kErm+RrN4z
QbFP8utYptyAmKOTQFggIBrOMMYCf8WLeoVap5JUhTANHdmicpcmqKaFegBdtZ1I
M+hPKmAKHJEUWQI19gItg9nPVEkTI7u0v79VDJ3+OZuC4NKgA05cII3qnZPG6KHL
5HzsVlF82AAaIM9HLvWe7JHdQW0feCSgAbqSdFyZqiagvI58WjypIGNesemxHuti
T0ygMx2ES3Rug/kiYE4EHRXyhcsdyEXA9Gd1f1DNFYL6g2L6F2Z/wl5RGAnRamFm
OIVZWD8/+6iiGHexy1U2fuwvRlk4dfe29ngMmfQhPUZKafSrAZMY/ZkvYc/CiiIh
dy7SZdehaXBW5ehvw1/XAtc44Oa472bx6vg+1MBs8UWfrhxqaemY0tNl/7O7Q8/H
N7VQb4DsIj33P31wKt2iA5+Dd9iyoKkohO9UQFScKaLvy7WDjWYlFPFiHMt5Zkhv
lSYvsYyg1h/8pELW1/bUrAZOR//44/fTP7DPeChVs+z8XfZOb/TxsqSuARrnhlAc
HTO5Ntz3Qtw+mM4bVBAJ2F1oP+yQlabXAtUK0W3FybokLmBAEggrpGyfpi4nMPY0
PWHUgy8yz4wlmTALK3jxyKTEJh87UPVhhd9aYusSOtORtHvZ5DhlNbRwESiw3mzV
upcxi2AlBNoXurLgJZShSPlVj8KLn+Rye8RiFwP1gYJpEEE/1gQ7tHbaKXNJWIwI
UMGdliJbl4JVWPEW2mvjr9JitZ+r0ZoP+yULFjfqyfbHtTwzJZ7MkSqwM1cZlU7D
OdxdknIC7AtC3j8NXpL086QFO4sm9XlOOvT3f4n4YHrm5ppPkz+q5TGsEoTaaZYo
kQqPkk3WyKrqd1y/lOPyahJkiBpyUJHBsS3PSaw0JHNp8/8NAwIxmOvghIc5aj1i
Y90c9IOY9pdaL/9PHJIqxlAYsl0R/lqZg3hnaUsWwog3fNgXwsHbBMh7rpJSh5oK
SARQ7cK5nl9R7M3yTElsHyliaATh1923gcN7BDu2cKZQdhnkLDg+fsKyZfp0z1qM
j+RQku8ZGzSzauY1wZWuAfpsaDT6eHET/lYvLgRzEhoQjc0YbdJXGScEhbLnTf5d
HX3meZhZMd2zuifmR4MHORz8tQ6J9hXf8Wy6cwSph/4GRxY41ZDTsmw5KOxe79gJ
3nm84g/do9GDoa86nxX7SfEKPeTrV3w5MORm4EQi5F34d6sUWvrC7jRuGCQUuQ2V
bLAhoAlRx9CBAmr5rzLvi8xE8yJB9tAsgTWpQtN/YBjEObZWH2LsWzUw+v7YX1Ar
+ziAW81b8NHiri+ZaeOp945/fH5MHREkR9KNdwggmfNHtvFLLiSMKq4DbeT2UoJV
2IxWo9tMDy0RarLRCo4uiDvtcqg6k0rRne+QtKqEg0TwaBmZA7qyIStZnpC7wShb
ejRF5ULFxUxkAdJgfx5HV4c9yE/yTUYHlqU9Bu6hzYv8TigjNPuZ4+HKwj3qwL3R
0qHTTdONMt8Ir8oB5hk/nGVX6t8L5SohfzEM1jFNWMjCRgfhEkQFcGwBPM3LLjy8
ktH/Evi/NzqdnYYVElUUe2UagTv8Yjd/4g+osvrzLp7I+wfokTS8ttlFkk6dKUJc
EDmLrHfmq/Iwr2y412mMPIIfrUWyRwMzqNJL/tUho3WEprcVRHw3nk25tlxSIO1y
zqTuzNJGhzd+xgq1k9XB4e+1koU5yXACxUn+og5L4W1tlqfocJGsK3pIow0hmzyZ
Rig1Ft+gpySSVv5X6gAlBO/c9mXhJ7FGzDxjkEBXxLqWpaO/xNZ+JhXwBUQlsmrL
dtnbMtOwUFAQxKctpYI/fAtoSWaaTNYeeZ/qlGaAiUFHyAI8K6Do41wsSucWaJlu
DFJtXlYIO/VQDk8zCAktN89rbhr36YOwhbnKRWhgBnR8CrEwvUdSApGdhFUyVW0a
c82fCCYM7idnoo/La40vtVJRzzCF5Cobyo44KwCp+PkdpH/4P0eH6P4oeQ78+Gc2
BIeO0W8gbe+p4FE02teNVHQvO+Oyuj04NX70fdfJHTcGoTOeT483c3QfRvj2BmgW
glhNU+v7cEwSjABibzDHv1Zzy3+7mRMI87O9R2wkrk4cUNINSuZ4ABpveWFLhTiu
9xZrLmhcrIXE3NeUO1UXtQhDmtMJva89ReEoZJDRLTHzJ4c378SsFIoIKhAdvF00
sDrlsSkj+PTHiEN8QKJpBewZpSGawAqlmLA3uZ4GvYU9njyLxziAJoY0gKVSrWMz
enFReuCkCJPYAMY9OXio3aLyeBMn00HhwHS0bTcfZHB+bKTe/iiN3kZ2yf2rmSdJ
TED9NOTfH3d2RPWGAi5ZWXPnKmvryCPr9zO8+mxFRd80u4rUC21TF7V0pfc+RQvN
2sVz2TwQvUKoIq+AcSn8DfvYJsEqVJxbPATrIHfh1i+0+R1Vj4VgpviWVbwsP2HK
TZlFeQrVAIHBowuLoODJcjoP55CGTEqdEVWj3qBADRZ8e6lH1yeKjYzLhVYPCsl7
ndoUhnUPyp0op8B77pmA4Pj+RzLeyGJ3oup7V3XSMqAuYt6xci3oiC+Q0WI0qbdK
P9PnKJ9+DNiV1wTBbq2LeIqSaS+NevYt1ef4ZZM6T6s6RH2EEbrzq5zS47CVaHwQ
21fZjERhpxEAX6YRSEwDK/+hFfefl5QGG2UK+XfrcrZzdCRJN7Q6LafoUk5c5Z/E
f0Af/xGwPk4+l5xOEhid6X43HSQxG9nWZJBjH5rWBVlfyMw1D9fXkEHaV55M6a0k
y+eW+rNR1sPz87K00D52UWfysg+5pNSJmZ+bs4VW8Jw4GFEcq32MD/mSfLoJg0HC
StelpuvFpTCdIt8E2IbggywOs/vEYqAXClj/FG2862GH4lZMLz1zk1eR6dyQZ2yt
lU3fISJ6VKlLWZvkgmARgJarOa81qUK1dcXSsTC21skvbvSAtDVhAbnQS5l4+6/b
PChQaJ9CLVsjhQreu3oQIonmnaoztjsGgWsBpLOpkOOx8LjuEWOta7+zEU7YhAMH
y+2+VvGYy4Ye9O6HVK4GW6YGraGoyh+Qr0m8c1uS/VFdpyYMF4G3LNiybjutWEXx
CitMRK2qJsgfMe1f8wY0XrG6aaG+hjueiLfdWgwRJtbigLrHXOXNmnG54zS1ebuS
olutqBvR82AHykMvo7iDhB68PcCrawwLftcV5T2Z4/6hVsSXITKJc0e6R5s7GoAE
MaqSthj+sa3wzCp7tnOLKlLShe3O1logHMpG/H7jYpZ/RA4m6BWTFEsTzQhrPgcu
0ngsfl2/ggCEDjiTNBbXfWZoD5DneU354ZmsM4wwQglBoB+rgvJFYHv+DET0gChT
oVqBIgiGloDsrRvust8R9C5jgDxYGKD2kdXRAPj0F+jHZKvAYP6CoQWAMpgKWnhl
NClzH3QYkVi1NX9iXyoPloRBbO/8aF68a8az/wUcPn2ai/jj1JfXhpGLEYayGFpB
WdAMYrB+XwXr9Op+Q2IauPFSGQ8L4kJIz3HXyduLMNEmuBGBkUleVp9xIuUkdolf
zDIids5jMWQZ2fD4o2JE7o4Nxd0dxQrn1sSp1e70zy+Hw/+m5McDECHKvn7qBZTh
MU8dgSp62rZ2cXsZqaikZDZX5bRL7tFeoJQfJAGjdbnz598QUr58WwmulVtwUSVv
F15wdU5LGaC19FPDMpU8R61IPqHg4T2G3Fve9pVl2nSolhR53V6YVau2iMacnOfB
QhKVFGWId/z8PElPFE69FEhU82Tgqc3UUJqhpACpf9jR3MT/2N/tyNkRrPw06vsB
5X3A2hh7juH+9tvVPsV4UMnqHwCsaPGyIPSgyLd9H9rdADDrXSHvbgRqETIZTe6o
KouuKgh3zLriYjNtuF59k42UEOa2urHk85gxWUL80V0IEJTM/KUWrqRiLuVEEq/v
XfHg4oUe6aXSqLl5y91/cnuv43Iia4Y7bhzQ5rQR7u82RSZ9wbVZ+BuOMRtw0BPu
u7DYPrull6bR/hwrgEr9llvHrb0RGPBkBQubrB1+7KiXgBwFYI/hL3XQm44jSSWv
wik2sCswiSQzHtZ0c3NIU9NR2AlWJvoAOLKMIcQ4FlBcsaxDbw5+DmpwR7YK0kLD
lEFjCx+Ulw9FU21EeyLTgwrp9KtHr5UZLhxVSkcvh8mxvZpi4zeX/zjt8Y+JXHmP
efX/e/z4ZO+DsiNv5yFeN39rtdpB5f0v2nuIf49LmnNDDQ5Dg2M/GX1wVbPfZTYC
TQIyRyMo6GuYuZePwzYxD4qDvCKBkgWheK0C9gTbAvsURyosFsLx6b1bqDZH0nRc
a33303dVsTyEOcSoInw1bBvZmVnx8LRbhO0vyqorGdkUCUp12GuNxRsuf/XfMBYQ
3cYsKgqyLMS+d3BKBR7VkLot7Fb+bCFnduJqYzrbytEmJIdERqb3mXZFeRuUssx5
8ITlyfhdOuLsO3l/mhM9llxCM9La6dwN41S983PVfsA0mf5Ltyna71JgofAIW6TF
6iMH12QjyND4LcPjlioJmaHY5SApbGJjzFYzXSCEG7Z4AUjBHDXX1EBdOWeqEaIg
mDpQHVvBJQEiRzgH4e49fR7Jgggw8JKJ1BPKMfayTmi1S1Tj3SWt4H71lxfkW8qu
qIfXda1IPJFsPNqW/+zAv8vgHQ/pSVmom37uRg1BLoKML9iEjdmhGuAMwEJMJSul
UeOAQmxpWVxCFrj4jHdoIlHk68Zql7hTSaOsHxcnCrKPmtTJ+zze+LZQ5aWyDJhg
GqAwDE5vksyu2l+pwu1Cu0JQdGoO04W0u8Iv51scXXQsxiG5NdaccBqfWpiQ9eUP
6lcVdd/w8wG6a9vCwCcG/12bAMJ19DGn8DrUlkKzhw/eDQIodThhwSGC2kSBCI4S
KbZm5BWmOhoTKGbBL9R8IXRKjx0Q3WE+fT3JNtVc2yGh8973DmOvTUxf008uhoJ6
nBJq3CnjhOX9e4vLdi359x6/Hd6jq5SIWW6bAu/sq9l7NejBRYSuG4u05vcZh+dc
uVMF3IM/j+gAW7YO8FmM4eQ+5r+CL9tSCt5is8kA9JY/7PUndBDRW3RUcq647Rhm
WpKbotKSdmGskKxDvyH+tCbAGOV9ICPu11FPvEbP1+nnlkLakJkKrCy+RPlAAUPJ
ZDLnvvsyApQzyrGu7CDwe/BQfcDMhPjDnNrnCi7oFBNKfzIKNk5tl2Z+bEcZwWUt
TIbgmzT07xlPW+hQcVWx8YCINCzY9BGCg40Thuewi08O8mxsUr+LR+QCnbxt8/cF
YeBY/++XimUQnXmV20V4pXLi+Y/df7m9oeL/wIBP5NvrS6w6uJGCztyOxx34IFjZ
DN/ZVUn7tgFsM8Bv1q8T5lO1WyX68X67l0yOM9U3Dq4uEplVkJyXAZOOA4+1kbYd
Dz4Qaz2P/3Vd8mdZSc59Oo2YNDQsWWcGSCx0Pr/pfIOxREKvJbtGy1R7wCqq9Oyd
FF44RDPMTPn/5hF6f7ZkVPJt9ziHwQ2ujj6YDwEnT+kiJPAizQQE09tAzyfOtgh/
4Fn83xOZ54JwWMkynjE7J5EUnLv49m9fFVWKWVX/6th1S+I4R6BpEVTGq7cl0muS
qNg/UDmtsIpEmPhrlgY4lBPgzDrq7VNl7ZZnoik1hiJ4cziBnOOc9KlGfjFqVRZl
tjye7vchqRL8tGJbdd2qFKPJB+icP2fLnGcpFKIwBiW7urMTXQZ7Y6JoGdx5cFEQ
VfLLrwMg+b/CHd16XxGXB8UqbPy4lQ8nB2mognNWokGXeyxcMMcy7Q27N3XZNZYy
SDWvhlWls8LqYCnQCqFhr0jG8WzzNVhpUviVGXtwXnlpXyoC1TkW3ouHXG008YX4
JytFsZkJP3jsEw5Yv7joQ+/sQFv3XdJfpMxF6oFfbxu3ANyfWR9FnQPXNRr1DT/5
1qZYT76S5r4zbfiSmOUJD+QSTvCsl+bBX3MavOqUPZSdcSPE60Q0bzqPzW4HkWeF
DGQMWeMapjored7Pco9kAeLb9uGKMKglpNCoVyBAfbkbLcx29Ktft7eb9q2tErbI
oGxLjmtYsnRoaES/3VQiNJu+yS3BMhv3SElYQNe33PecYEHzh7qX4UGJ3dJrk4OY
sOmHIKH3Sa5UifdleDddlcoGszT++53GNk/RL+WEchI0+iRlxn9AsGp0xIeivbd5
4zHMKc+wYjwp8NP19eojXVGySRmggxzrWtA6Wmq0dxEe9CNWjo7e0voyqwJ6RtKR
7epsuDrD1ywjKiMzDycTOwr6ww7tpsfBAjNj5AaC/8a7V6HAkK3d24Wy4pHUMCld
WDGN3oq++55y/fOjGWBFQ9S5r2mQaIERDpAH+NWP+tFuNZSfpZouKObn8/TVjV5y
9J8r65iJeKSkwckqYwWZqPQfIIu/SMdndfOCLNboJr9Ng3UjVLjnxengjeLGameT
ukFJH0BaPUkiiisMH+kPD6nyXbeqgPokHJI9Z3FUcWui5wRdrW2y+MwmnHMSuueA
xfv5XJtAaUprAZCFvC2zwc2MYoM/XC3+9JgwObT9EF0RroxRDl6lZZGrNjKrIZlv
n2w5rX004IWFJk7tuyZOSVwIL1DDLKpEt8TtrL2/VP84Y5nclMhmVcfVbIvjhr2Z
D75QjBQltZ0led/bp3i7i+r4YJ7gfwojU1OxExTnPihu29k8s3ESdTLqnG7uHSE+
MZRrR6HUr0GpdTJe039H2JN8CHx4eTdF5eFzJCbyfOFqhdI9wGf7s2fuqtgb5pSv
mHpREVdEcW2UMh6c9wtxr9JF6Yxpp4RgIpduX4Xf9h7Hb2/sa5abV+I7yPxSnAU2
1SBCqSqF6X23mW7W/npoEa27HhLeFX6FeP0zKrwTxsdz5a5g70UkIcNYt6aoo+pV
tkOjnLlZaVBQ8FkMycOhlW4bDp7JUHwRffTismKsrVRNbYykc76ABizryjO1y7fJ
ZSZI0aVKA1eZ2Qu/K/urjvrNzkpqTc8LJLK7HtSY8saLUQfyC7dNl602YW+xXEAX
6EcyQv41E4VYH3mq065UVE0TMyvEcdTWdJAFTdQe3lazI9PCWs5KNDbBXeCn2ZnV
p4Cp0SMbgjawTe+lVNRxnU6XCmG8gFeUWWqAm6Y5GEk1lGJDMATAjbqr8YfA3wyO
GeDIeGNxzmTDNTniaZHTX4KOftEflWID7EXfeaP3CHDJtYCwP56xaLELp7j4BOqN
XfDTEsdyWVftar/DZmEs0F0ZyoRRMRG+7H7z1ex9jTWDG1RDX98/uzt7JSK+GqJn
kynuo55D+Ed5ntukPdeLlPKoVqumLye69xivG0EI9rfGLr5+IGM79sa9Wpe/Yt/J
B44akGygFR034escjrC8iDJPA1wglBdJ/7j27DeoNUsmghfQdRUhmyYwcpZewBsa
AcvfxAB+uqdeAL5NiNFNb1hOt6HH2oRUBx6fk6e5KiU5lY+xeMc8ogJY0xt+58tx
IWQB3rTsgkcqNBtDUg1sf7PjmrZj23u3E3nc+XGL1sYldsksRGmmoobUU1UWS4J5
W4Qs2TqOhWAqL571rg0xMapk7JZJcQ7+TDvbvO9Dfz0eplQLQiXKEr0WPHgPGohD
qLM1ZGPGUd1J6mjEPDlZh9bhG4abJcIlnTYqudVXs8NDsF+WJpVRPIJ6CC3yQglF
+B1leOt1MllWLRKVd8LKxTUHJwMog+RVt15wbfqcem+H9RuKMAYoGIMca5oT3IxS
VW90pbi07qD9Kk7U/2pB54s5416O/c+7ug6v99+BAsIsbe5XI0UdERjOfwGt/EFe
bI5QJDku9LbZcrWPG8wlOpzvjVmGf46YRETqy9w+Cic2++lTreDRswwzCYbMaav3
QSutI21stEFiLOgAziTvMH95XtUBn7LTr/cN6DTjjFtFdAnwrWzttYEeUiKVgm94
XNYVT17VE2qXiXReKb8vUNFkG8+D3B3S+DbR4KEQu44b63AQsdlJ4HbNhnNr2Asx
/6wSnqDdwnhYHpI1KUn7ROaj7qdoUDigTVcZc5GavaYwx9QodBfv06op14u0CnZc
jc37G2J6ZXaCB8L9ObB58ULwQU+3GUKR6AzaGilq5KRJMjtw7iwWHwJTmG9OuVL4
6nXayIKLQgtJ/bBHTLdMdz+LQE8iWVbVrgcyVjjEEpKEME1Dc2ukKcDQEzYvA+0u
T5uUN4gct7e+CONxD07bVd9cvvBhuVz5kGv6g0l7ZuFeA5ps7hI3/McSIquGScH3
+E4FyFmqUmtqQ6HmRYUpvpEiy0ukbjac23n8j96Bje2EZN3d5Lpqn+z0HBpSqRuG
wTF63NTG15jURc7mK5RlpGthnXudZReJsH+RBn7TkBmO8A1rRn/nfPSwUBa8UAZp
LzUVNnjKudR/xi5vM0kAXMjJy0efBNB6vVr9RqhKTKN/bXby1pvR8LNyXa72GBuW
Vd4Cd0Pwr2S40mle5dlaUsOCgm+N4MpQ13WC7lIHelotNMHk8xSYXuQYTlGztrbd
pp2ctRaR1U3oK0dp773/OXuo8ylqY5DVujO2ivO0stGvLlScDM63tH572gkFpOGF
Xk8FGS+qF+y1D2wbRxZyGSkX9wxxiIJN+lA+H7Ck54iLAXwW3omHeUJX3Uwf1Dvo
ZWS7hN4B7XLibFj83DDSJJ9a6Nk39QYy0wc32Ztxc9LKYPcpFPKQ2zw2/dTBIKTy
Aw+bGWxLB3ZWL/DRNrFIWviWgymB8XN8PN8JRULBjfQZakEQwcD5J6gSj25DTP8B
h11m8JUDLOOQH1TIzFUYOmZDsYRdtS0QIxOu6bgex0Brt9E0z9jGjLkVxg1wHGXr
fYHinGRis0lmfB3utnxmPIaha0KgGnUnaUVYyeGFlQZRD0EGnWYbj27PG/e+0tLY
0cwIG54G2WRIUnE6nfiZpNCCIOZYxB87IBjIj6Iei+njWmoY8EeXfyC1zobzTsJi
MxAwgCR0QTH07xSvWFENuFSiaZVumSHc4njXellN0wKh3TIs0l0MzkY3oHpvvdhs
JzrHNFh57uZDIoVgNsOmsdKm8J9ptN4P0/QDbf0JBEZjv8FA8NhJ0qqX/hCnfJdR
rn+4A0kkcR5dL5eKmdLin9Kqx+/hB3/CeZFXx0znVR9kn7yVUKPrioxxb3m1Mz8y
x5gq6Q5O2sHG6GBkIOjXplkFoEtt4C/YTIwimsEFkUOgcptTByriPCFHBWuOsPHJ
WtNMHyybtqBZuFGcSzEipLvPwkRvh+qc+oqI0ziffP6pOilQY0/wmxWMuJhrW/BH
0LRje7FdvDVMCMQxeYd8go+WdCTDO+LBULGPo2SBUfCoXYJ2WNHkGpKSIdVP8grL
YF7AsOxx77+L+D2Qunc5waXLKcfJK+Ym/jYLudzI1azWDfPQqsmG2vOmGhKsXn0Z
ISQjzmkWDZcwOmmxvLM6IYYZUsorYEtEYdrnpxVL/ZEynWo9XHKdccM8HpjK1+DW
SgsuIr9gMgFFOTm+gcBIMxPlS2CmCbdvZgPKFFHA84EX63e4gem8ZlMxOteF1VkG
CLP21dqQ18rU0b/AsHAG7gaVFQPKDP8dSFlUy6A+e+hcSi818otsngD1MFdT2WdH
89XNSEZIWwpY/bRskAss0a1TtBKM0dUo1/A7ZimnLSrQdpbUJeEKduhV7K/o+o09
KqT/jOXiqkXdDFHvhj4+vjCbvsNU6N8rK+jTdMCJ0qKbiZihOWiMfgLt3YH6MY+q
o+BMyX/o/5ZW6AV4dnRuyzEbGDhoeJFurVPl2j9/W3ADs0xsyA9zJJ2w5Pm+UEi0
Sp+trAqL2wwbxUMKnll+gFnHzNnquYSe2CQrTci58DKeau7fH7gnoLmqGP1B0Lv1
r5cSu72g8iIjYnlq4Qc3R6NiJt6G+L20nEmIc7mOGB7Tp2g2D/PX8XB+lB4119KF
IRKMilKve7CayUVhkHV2vgGuokD3VddAK89I1GiEp5wo5myp749+Bvm3Yc0xHsO6
a/6rf4YOib5+FWQy84zV9dQx+8ZnSVonh1uyomNcvRM45e2pfC9ESLHVzcvibn7U
1gTlVBs3iWwBDcf9qOtQcdJ1TFf6LoeDPxNIBmlcHTtExkUc+BVb3w5lK009yphq
VrtW1meIj/iRlC4H/Vy0nggAkeH2wk8Uw1EzzCJNfGjnRy7G4O6n6WrLl/zmyOs9
rgjIZqGmAYHWXp5CggOEVHQVyecSKHMVXL5jfoM3jpB3JzvWjC7jdJifM2msVsra
90f7xBAgfqZklgnCOax+mpQK58jxzpEdf3SM1UFvLsZmhcPdlUFx1J5ne3roIIsZ
W9cUR1geR8dwRj9p6Of8qGaOhw9K99OQv1pxVRWHhoVZvF7ERvztt9J+OFIVx577
EeMJIduumMsz92/0YQWrhwTJm95VBgE2wKHCHrv6nozspqKSm6G3+bAyTKRuofc6
cAhGpJtIrSQYPniLSJDkfffc7xnsw3TO5WuQmlBZGbRNGmnz44h5etN9/X6/wnQV
mNJxxG/EWGoFVdLtisUJ2hMep9CTxMPbezUHdAXsEkPE3iJ60cI62vc/+3ZRwriJ
DYuASM2tOTUJiuaR6OsUFozIE87r2l+J0uQk7pWun9dkP7lSzJSzu0mbxTov8tO7
HB1MJdk//dx92kLQuX7zPuY2qeYGzSiUqdFk2ESmDg56mkOvqa9+jlvzPS+QLnEY
H65uIo/LIKqGUwDQdMLPP69z9INvjAUQ/9fnIPjC4cytJcdAuwFpePEjmzZjSuOp
q5D1HW0z+NTrL4pzMAeRDwh31hTPiAaaye8ZbaSacRWTCt9R6drRLrNOUfgJbayx
mHO3D8jX7UWes3yhBB/1ZusMRG9Zi+Y8VLDiajKDtjiwyVP2eSkQOUEiUYiwg2uN
+RPWZONcdoVINY+SzFcABjNGrwrkhmLLm0Gl7Jfsptt9MFNBPL05AWjUQYEaGggB
Gep+f8woSTGUo+6L2MHfMY1zaevz5S/5Rar1fCCzQ5juSIud5zehs+HI54GoGzbh
uX4mU7VtD+Myqyg84amRrb4Rn8yDg+/KRFrc8VkkT2hps1cvxhg58KnqytlbrvYB
d6/Y1rquSyG6/yWe+14mszyljiCq3yORPbGLSU17U17EOHIOzuO3AAFoeBgVuZrQ
zaV4XqFFBwfW03soCEawWU5f1nq6fY/Sd4n43NodZtGNkSp6AGrq8pfErNYnhWaC
JMSNvX8XybuVQY6kiJ/uPzR1syCOuvsSsprK3sCA75hgR8Mwiki26wl8dfkSu03m
x/BCDbW9OFW8d97bYaUgdF9As14/mpf9OY+TSvSVcop7Y1WKNYfk9gyDbhILPTcx
xGDm7ObU/TVaA7xZDcz3As5emhNLkH2AszhYPFU4t9W+TxreQCwvzwj9v9doDE5/
SphuMpEEz+TD0H+lcYavJyX09xVivEN5WLzC1TEHCPGiM9nHt9YGxbMNiPahEsK5
jI/agwsNjLQOm+ElhWNLi45CfXV8DuK2dfusA3OGIgcYuEL6417ahPSh1MrOHQY+
iuxG1OPtY9hvxYT0MCDGXRdOiyJnHiNCmG/iGFRJKCyfe+Na8d/+TC5tU0n5O/yv
Etmv9uMAftARepWELmMtL63pU+OR7oveSUvYlSEs+ECmdYdVcMEmX+dTBi/0g2Y9
mWD6wgG8/h6Yb+C7bMWJAJMwguwtFjJw9/KZlcBeUyMKaiBVbsDp4Inxam88tPwG
5WZA6X6zBZ8rKPt/TnF/3FnM16cjRkTZ3I+zND++nBCCnPQbvkFC1dJ+0S7ppc+2
VHfp4C5yNNcrCOw10Fb731m+CRGzXWSo0sFj0XiW3nL9PJP1YUNTgWf+pekJSfvG
pmCLTqfekvIShihtIIRH4sN9i+jHhrASv1hbhmJYpOEmTNlSOEXO/YmxedsVvy/V
wCT1UzxYQuvICk2mF0zeNSxqzTRhyGU04GZlLPTk4/em4FZdPvid56bznaskSiuN
McZuEYKOcrQfIcDcJw6B06MsrVMHEYGI/Rw+QsuIPe5WNGjCgHjTHBylX+mkjgEz
v1zDdAQJUedLob6wKcHzmz3dDELhZ+ONPAGcmNNXzJcJegol7HVJS2JEQKgCDios
mjwG4C7eJMFQZ542D8m8M3feeeR9McPs2wXw3btp8VDGj/Haz+729j7kT4WUXjml
5qezVFXlae9ZMpj92wGJFP104AHLhTZ49BRsPzoQVmqA4O0kHC7f/70hFUm9sJB+
PwQC6W2obCQ92WtqC97QqIzL11Jb+SiMscn+QnORd9x5cl1D/bHZJX5e3pyvkJry
QWoNyULjtITacz0LWWA9UnO/Oe6lf2f1o31xMFM45gb0CSUVTZce7oAYmnnEH4Oj
IvtcYYDGTW63cb5ca262oSnmXXqErdevqrcGQUfvE+D4c1+4Emz85K8RWD/tsX/Y
rgkYmFV6xhOZEejONgV7gjamjAGPlBYYNmPIRhYSh8o/7ludgPla/wp0dxGxFFWq
R9EPsMp8m21JnaZA4b3X1MzwzJqeYT5IwfXnJrSLUd4rbJ39C8ELF0Ln035G+01/
3bBlV81EZrHNjRSyIzwXWJ/I6lEF794u0YaWATbwQoMax5uI11Ie94+A7dIL4Znw
cCGlEJezWpD4P2+M59+T3BwoCBPH6IEbgHrHaq0dMbXMHCREnfRdtjs7wwo9kIey
RQvcs7VhkcfqEyM+5txikm6WrxfTPoqbnspdb1+jvKaVFUH7xg/iRca2Sc++Dj86
7ZdBJbrNqeiHWsAIqGvtx4WpIhRe+SR/Tmz3bWWmBNC8b4Ea4lri4owF36rt9qAQ
BJ+/0bAbWXGqU/u86zh08f1sifPXiBEX7RYTdbPpj8HxdVkyjU+RqWNEpUZT2kNQ
xoMNKUDjRy87dFWpCn760WZddHbCyCf4lr6y0VFHiLXLVL8D/QNfqKpRnV1xNfla
gkLaorgi/LcIVW8I0IRaapvR3dUJVnBwnwv8X4oCsy3b/LD45Z56zh4ttBrCBQd1
bzZNjVuoNkC/JG/aSzI+2LFY1uHFQTV08r40RqUg9+X1s/YjLAdh7zKkDv5oIJ+Q
YfzTuFnI9absrNTXaG1aJ7fYwUBYWixh9uVwLcvB7E7sBsoxBgxxrggZP+eUlosd
OzjEBe8hDVbnrNzMPJ9USBgsrI8Suqun9L8fOKT18VDu1vk19FLwjOn/eAKHPrhh
aveyPDPpzUUCe2Eg3sZpRu3J8hhamIkz36s2obb45nLpJQ8eBkB7nNHZItny50Ok
n/t3whAv4ukIFruJEWQplqxAGugw6b3MIOQy1oV3sMCsLrNIfFaQ6vFXIxyrH2Il
Y+Qn8TSwNWG5pZ6W3gzABxIig20Z5FL679xnEwKJbmWWH/qBjvTaROpoaSTgBS/h
afrFfRJanP+YD+i0uQBqM6xmwV55u9Gce41OgZ4AqRmvH/LxvUFevXn/fGyvt4Zg
fdfPn76iKQMIJuzrftBnhioOUJOiw9zEzT4b6CfFYG1VYRja14rP6IBwWk17WOHG
1u9/3QkiZML9WUi4mP9i79cCQLEskULiWpD/yocXwfhhO5+aXCqTJF6jsZ1THXgv
0SKMluPpUQRMj1+VcNsEST6IWivpTKV0iRc7wH/E31B2DRaWQdsM4gFyPK0MMBsn
ree2Up1dPb38OcEUXqrRvJkt43fikhTlmw0swXH9yWoLwNTKai6zFiagp62q8mY7
PnieIaWhxiyu0CbWURfEumDsNW1VpPOECRUbN+j0IDC8yBtODbj6sCe+iHztSzsw
NqLf4K8zcPbvf2DzfmJ5ql8fnxSmgYUXeQNcnI+/9XHhMQJfAMFPDHFxIPyP1DBp
7HjvodW/Rk/JRFPd6JZolpybX3rHDDnVInjLkbCuRvAG0dZkzBe6NENyHw9AZjHO
RTGelHoCwImKF8X0OuEPYPLxgwsqFCj94H67DZhKWF6fE7LORpELXtjrf09HEm0I
Q5bqB26I8E0632CZaG6nC/ANeuQkzIcpqsgZiDJoR34v7F2bA9Hr4T53HK2rkE2E
hVRDgDP2RdpGLVsuhNeo5DKZcjuME1E5dhR8vk+pj3LCDEQeQi/fGnol9cqtx3Ak
zb0O2newsflIF39x54Se1MKmMa2Oo3r0866UqPHVku2mJcKvKttOvvF191jYHk4E
U5DiBreEVCmQRQAmHL/VkReIvPvTZFEh561K+WDqGzqll5xcpf+6A26UijYYmu9E
Pgu7SCO1i6N2P6YrQ1ufd08a0WgUYPvO1o8vHLI9RGzQ0aQ+Wg1CamW+8lDsoGBT
s3/kzzgYscO4FgKU46WpacCPHs1gkYPRy7t5r3k/AwWiaPiW+DbDpkzh0R6YD+Ds
culaAzs1fl5DrRXAcPXZFmSyLP+VYJb5L1MG808IZGb9hVXH2sRJpPEOKmMusOPL
Z1DfFasbHtIu8dS8kP9vFEpNAfE1mpF9F3GU/vYrYnKBPEe4SxteOlUgENkjJM8A
Z0fi/Gw0GAiGmTZS1hHzpS7cDm/sc22XSl3/9DyQci6u+pODqy02FOEnQvls/yPM
wJbVwxwOGOanx9PXeVXQrz2QLbInkihq8v4cvzx9Kx+7RORaUmVTjcBrArZgYprT
tzLVhSCoUcpZO8vCHtdC0ydkn8cgU3iI76bRKA/z+WdJy60MmmXLX8HFZ2sZZILg
Yzya9M/2OF1pVYbPORPTF91zbrpGn7Iuaoy3lbyXzFUFp9kDd3qh5z7fdKgdhO3C
rmYclrTqch0h7XmB55aFE196KzHqm/Mev11O0upDQNU9Pi7vr5v34aDHvbBypvjI
T5Bb+29KOezdabKMYWefoUkpb10WWMMrXAWSTae4FPLVDtp3cqJXGUGwgYCw07/b
VwtYFtdV+X7Jf5OC84imHNrCoADENoIjDzW7e4oAowbbM/wpoEZSq618BKY3ZwOp
ICKlnq57BcoZItBkwWarN7WQkwPidqwE5iG7ooHB9Op6uNCsP6Bza5yEZ0ytgIWL
NPOaIGMMDgYbe6IcrHrkMGnT8nECRApY5KlBA7sx6HzQHrqIONAzOIbS3G7GC9e0
zwZV+W9XP3ROyhJJk6aYhiGqLe6/BfdL9CSKdJQLArjc3vUyuriA8qW2Bg0l6OMT
uPESqh9JT1pBnaoRiSl7lBOUiuSj36BoynneHKn87H1fUYcoMMfa56rqj4kfSc8Q
EdoDRpIoqfFAx+DFF7QthxXuViPEq15UEDXsTseUNPTYaEzVzIQiOiZqcVK7StJ/
ymHO+Gw4IiiO8AzhskNgvu40x+YuapZBck038N+e9AEtsMxsP5+JWlSjwEybUOsU
EYRreh5joza51WWgdo/oOtyp3z2kjLkhRv4auWZ1y0nb+bR1ESVliWSsMSrm6hRd
H7JaPwPFgLGrXJ01CceNl+NcdXKzekvFFvaOsORvgoHW2ZLkTGcSTVDpsxp4dCs6
aZFxu5xoqEMYqXGvTt6cp/Z40CBCb1vFxrGcWpqqz0OepcrVXZYSQ7XUg7ufzQh6
g6h4aflmxQs4FJdBfx8qGA+PAN+H96Lul6gQNTeKIvS+rBi9q4Bzy15maFrdLUaA
cuR4Yf6VUGla4/GJNU7RJzPZcpjskCXCy80lONatEukj1FbSNRyD2OKWmKlqBg5S
vhQoixEgIrqZ3uPOZ6IPq6M1rGXBAoaDEwiDk9r6xR/2bJYKy5m7vX0+aQI8yh9g
+VeyY3k4HdIWmUD1DlqfbSwGJo0WvIO7C5PxQKbo1J4d8DDaMVu9EGgSnRZ4KWjB
KagY8K5QUYl7q0YjWQPjX3DqPj8E7Qcg9KQsxfzj/nTbwXk89wkiHGabwNTXXDRo
VlkvBy4Y4y5TY7lBgcqOSeb46IkJISMgHMMazEN6bkVPlKsxnta4Vk2ZGuZDON6w
wdR74EVaVedQVLzcFu81I9OkD1heIiCMGUJB+cY/L51VC/fH7dR9Nhecv0c37oq1
c4cPJuJyymHXIciR1+opidnz/SVfWPAX6JH16BITZ9806qurpEHB/2znpSFxejc+
tA0/1Pe4fLwr5clTBj3YLnWv67Ksx6Uec0jPbbd1/PrFsFkuHi4hkqiOzCZIOju1
ZwLbwlVs6Bo1fLSEWxM8gsX2hpqPaqMvGZBz1asJVwzV8CFe/ONSEPBA6N98dcNo
3+8u3szE9Qg8isD1EhA4L57hrHyC8HcFzjUADxoM/veUbfQiLU/XfKvYuMGIuLat
QGDsmQCHWXOHOm/fmuVWkRE8sHwA+CFLFp6UWrFAc5A+uBObRNGIAbu+mnr+WFlo
OWGKu1BA4EonVRL3KeGgcY7hmJk1DUbIMNXlzsi2cjkSoP73pWDAAF/CmOyJ8sYv
gbLmUZSWL7NKR1iiUcXizBE8eBDl5QIKjqCwbohJEyiVNm9arKwJusatRF79LZQ2
DFaUU/kvbYNSMzo0k+Rhc32+q5XHEMoe1XfdArbuXm7c/buK2NqIMnsLgOGCXD/M
rdhGFyQ3cP4gylR7KMX19IeJ+E6iH2WQuBYZ+I9vNh23psCssj7XdTXMZgiOQEyJ
uwstNrWa0wciEa4Q1wXzTK4L2+pyOuGhk4OAd5szhAIoPm6VGAiLJBtM3dNhMHBP
fxFZi86ZlUmgUT4kgWxpo3RMYd8ZIOEJC+rFYoKbW+MX7dHpjufY+4cVtmhFQDEE
iV9WlP6hYgwuSScP6kQU2e9+nPXggX67ZFYvcD9ffLQtydQv4ucIu0/ww7Ek2azE
c6CUcsh4idVBEADDTKf8N+jd/HfxWudMHWARBPaHF2IZTfaWxYKQBKZENoi/EbQ2
fvD2nZpQfsjrFinpCwOt9qO6AwVIYAVsVD1WibGsmD7UJx+vML53EypHmuyaVGGb
1FIHELatETjLoXQHmYdRCP011yBNaSsWfa/gEYiJ2paAK3sP/dSqEOCoU48z8CgX
MC+LWfTkp3e6F5yEVxSoWYX3tDrxR3awR2iZce3JcViVtHZMkLLGQmpAvQWmv1r4
8gT7wjAIyTwgGm0RTK4N9yhVC43XgpTA7zcy8muc7fx9m6k8cq45MEgVNUjj9+Y3
P5tTEw2gvtE+rwfwRwP3DspZfPDFswIfEXtwvAB9MCG35tRBc0SfWbAtUbK8wM+m
E3lXC+YOCLntjQRJxT2etP3Goj0aW7gansLJHgc7Qa9mpBZpoe82snBcqnTN10Sd
Rsg1Zxp3GhcmuCmhXvPnJpw0wDh/XwnLX+QflGqYuhlGFc9rL71eaOaAgt/csWsP
hYmN+1wldI4MHuWsK5JStRelYRa76Ds9+bPnuiTQ+FKiSxzgZF8FUgOacqS/D+VC
/m1IelQPi6APQzGkdiDSDPFbXGd5luweJkFHOLtEcBt8fIuVHmbcWpqi6x9SQ8Ky
H/vbgWsxzl24iuQO5gmmMijB79Kqp5OZT7vt+GmCygkncXJAVMfwcMLu7wl4MCmE
mbuxOcKfL3CcfEJbMoWxhj44t7ad2UWV++uXqh+pNyicw7IQV9XXTM7jbepM6GF9
WfQWiOZxGjGUlhFvHJ4l2cUETkoANMrYEX7hziSPkd9c3viht/h5irICnypwpHih
NtldVKZBa7orzCLeEdyCaIdEptC3EvlFLOAa6jKYxmeqDKtL4jdI6EM3bV7Kkyq0
Yzw9z0BjZxfc4wtWJMRk8uFGoPw6ejVIM6g0V7lphvnBbjXmPRBJ1HR/jRqBGkXP
zQ2THMdoy5i/dAa/6/4nYXirPkqyKneyNkffnY8ddMrlcErFJRopMGQwiLp5MPfk
CfYP3Mtjh+woKQPa5a9Ff+grEJMFHVmOgsdgSyBFobQC22gZuIsuLpTiWxlZNct9
Alc3GHmAEoViOnciivLtW1W72H/K3dr10LYkKvhPj0aK/BgeUgNyxtwguPpzo9v2
pTsbwaozKBT87P9qadfD9zi15+9DRnmwL/IgqzdyfKggDh0Xamd8IBQUM5MY0yeu
9cSmG++LWlvggKVkLvEPKmfJwxLCqMYK+XysZpxpmsSrFt3Rccj9i8Oyxp5yyWXI
hLDgWa+4LQhc0iJuHGVrjVcjQe49UExG/sq9nycN0ZzYL+xJJM/+X6bRBF2A11K9
YSTo4ZvnlE82kusYYHiw6Z/tzXlnHQsnXVFWI6eGS0DI3aP9toYqm//g7rh//UCC
Z/q2CuOIrzWZoKXLc1zekAhShTcjNRYA6xF7eqiVUZAWgIlX/2UdJTO+4I/LRzho
4pJaalgH3KMlO8k9gHQi7xukVgZ01lSPMAJ9cAEin6SDp7yfwyqMfvsYQwHr+GNB
6G0Pp01y1fT4swoUl+PuXlfROllxQUsCwEruzgekLOsTcF33zzlNBoZjKy3lBEFL
r29ouOsWvFCJZ1HUGe9cRjkXPxvdwsAuYgEqxuNVqaoRAu4tNOxrBUYPP+9n1Fhy
jG1PvPpj5/ghe6ETeJUUPIja0HvrN9fgIOLRkvmVQUlvmZ53QDZWBhlPYq52gSyN
Qts43o3yFOrrWkvKsDAraK7x7onB4loIKlVjPfSPypWU/NmqmbC5H8q5qRcd8U4A
pHMVC3kkfqeEtLqDeOAPNnJ1vF10zugGyNjTVCVf55Uow6kKUp+MVHMP6ViRDojo
zif0rguwFi9mnyn9gii/WsedNV9XRB7bHzXNJej+s6/+Vl1Ptf2Qx0NbdGWST5XL
0MG9KeDVIZZai8/Cw/8+Pb9UM6QvxPtOnnxdUG6o0ye5kX32boEwk2/07fLppkFs
XwSj3ZcWHzzJswtvAcCOCbqfkHIeHn/aiufjZeJ4BuiNbOz6lndwHr/nvo921tR6
ivaGMILqPADlJIkKKalASje8iNpajGYYMf4tqB2frtF8fFbz3jYO4V9JxcQvItMM
wCLMGJ1fR3d1fH3A/D4cds8spnHB0RwfTf5aoEo/kl6sVjImXNoqjSxemDQlOcPM
KECKf+Ff8WUMVlmp5Wwz4gGoaFhCPsEjBzS6k0/Y/mBKKlZmn+zXS3b5pKny6f0e
+frS5HOT/c/1Al/th/ZpwElywZvDzagsRnRPiFNVFn/k7mNf6WHjT50hU4xhcB4b
jKwzlgPC8WWsZK7t8oetYvPiYccwA2pjA3+Yc+EipPXNUEmefNBfxyEGP3+f3wtN
72dKXbTi2WJ/FW2g6of+xsGhOECKNC1hzxfXBSydZAnMQ/UOxYjM+x7AasrUgCY9
SW3X8XDzm/+VUMo0sB1rkD7z4SCBheDCZW7XlAIk38lNX/C6TauvnV+qshlzYjLJ
tNwGvWAOBuAZtP6LTDC0OAXq2YiLmeaGUcRXgXqpMWZ9j9CcDONbsXJCuKz+cDKz
rKOtz9jqFeg1nWTWQKkdLQy32/IC/8/Fejyykf+3GL0Mf9WZlni2LBm+5jCkVO+8
55q4NLIWfaBehD284dC2UmF1dh0/S1rFQxg2+OQutkE7mkMSiV32ln7R8ZiFyqpd
ErCswBH2NF7ThDumTmB/xwHXwvjrNovA40UtOEHaOUKWzG05cIMTcgDAXvU13K+r
IbrVaCBWMIffL4ItVMUQYGB7+2hMelkCAs/9t5ClfdrsrHUIejkEi4rNWxvY5V5U
/KYZkXcr94p89Cq0gVXzUSZvmCWUJh8fScJwl0kx0pz+Csc2zNAZTfVNBSj7BvrP
6PiNwxYZ2VUJmwoqaWglAqgBS/5X6w7xs8Vazr+08bwchPlzyyjNgrkN3uz3XKfP
nmTG2rr6Oy9DAM2OewoMeiXI5RhOxEGUy6ctWA5PVj4YArwGVG6bzTf7tSfDL9fZ
VektPVe1L/1DLFSZNc1YvLIorejAEsAr4Dlsg/VBcL/YdroUjvfgWS9BgWNBWwmF
oBa3oMPXGQB/RVgYD7zfCwLW2WC5wPI8rnyTAJ4n/EZfwZKok97UNajm6TL+dyYX
HqUqopkJB022bZM1I2czEw0Y4vumjuBSo4V2aKw0EpJRFiHLyhHrYk1re1Pkr+M0
BMg6W9EoZ3/Hp8KWQgrVUy9S9q2c2C+qw6FsAw6rkPn3CLLIzHMvHt9xNRUgJFs4
yjDmyQIdU9jkgRAP6rUlzCmBIZSJB2Er67LCUPsc0PdwVqfA53hYJGlctkJat+7j
Y4nF+lz9CWTvUA26lsSKdA4NRQJimDxkddOj/bJ5EwX8sxqs7gQ7E4+MKQevcaRM
k7JhB90Nf/96MI/EZjxlER0H384PglYjmmQkXg606IV4ztQKjNiYT2l4Mj1oMPSN
F2sk4R3Jks/FSFKWI/Yheozg1ImqczH3gHPOqHNcL5ikCglpur4nnHpAEcSSzIxY
wGsnQ2ZHGNjbgErZE6mh897ykyC3lzSaxSFBExJ5uk3ggl/z/DGJ2P1H1UOvxV3G
QiSeBEgZpV/jINRjAd7W2IX/HKpqVsS/kpYAK1/bkEKfiZ1dTd1HBupP9DTimvM0
NMnM+aFWSZV3VHuD+6XDkFFmY18yYK20uOjswN4KD3IHIvYHgHAxnwnEM5AHAjE+
4CveApaYBO+Mmeh5vs2xtaloKK8KKQuaUFOP6MTirwZ/rEkylTZ2Bcv50KhN7ueq
G0ZjYiiAcb4NMixsunbYEhFKST2pEqLmDP2wuyKI/gkz6o1/8H+p2bCPDe8h9/Kq
3HYqj4wVkY68AVM5WoZruN6y7PhJ5v33lwQufmTqabxbyn7j/UxFVQPRA42Jk0gI
el358IBsfGQsJrbOtriSI8gfmfR8G8/YK4782JE0NlLJN2PoB4uo/Ot4S8CxMAZx
VIrFw0ZGgxUNRi0eQq1UO8gW4D0T6rHKXTn+gCatTD/hF6ahTMJOHVlTKp7lovxh
auAaA+93Psn91F+UHEZuojimHBupk0+iLHMZ+7HJzlyQRtrAYjTaPGVMM+0xLtjV
zS+YJyEtL21qm1RQn4zvtJwMgD0N/rsM3ZLoeR8qxFVp4lbEqIBpViCA5v8RzdTy
gbseWKiIDm7nJFCPOY6Vj+hjKHoquH63ZuXNCQQri4SmZxB6MRHoMy5HGQumbifb
xyYK0aKFPEfHTsna4STSz/0B6It1wo4keA7lpIeLj+qS3b0wkrYXdXRgxrYXDma+
voZVOQirWosX+x6K8dcWqC6/hsX9CyIdDXCGxH6lQ4JunJCPRLZSWzn2s2JXEgYn
PZ2O8g92v2D/9BHB8ZPeFkWg/0IRWP+axx3EAjDBHcSdMFPPUGus6gi4DZQ0thiJ
3io+vNjfd42R0+a3tJ81YFr/PI96BtnLHKz3hCRZ8iTl+mPB4WhUHFRlFzlybOjc
vjldX/ulf5076IKgXiDJ+ieCu76piw011n4lZOv+poSnlEFL2hCIGdAF5cw1qzRz
XsVY5z5m9QMmBfMnh6WAyUeob9zfiq9sCpm+kFb8GKpy7i0UdqigbmkPZ/Qei1Er
ektojxs26/9Stdta1usoDJLwc6gurarTKNnbgnq9jjIzjfACCuKD/SNr+clVWjnw
xvZIZdD6ifstEGW0Ijk453/xjzsqX46xpGZv2ZQ0XqeSa8IINTehIi3avzgSOY7Y
A8N7DLnOPSHI4pa5Ag4T57ZUJSlevtkQAaP2PVAKjpDqvtLvRb/QfajU2+QjeCf/
KaCMoVetX9v84yIebpdrhuFtmAttDsWWVvwImV1KN3YExusJavmWhvsR2b49rcQP
jnayo1SCB7ZNnbl0BTgYjQy+ouu77RCuBX/U20aAVBJLXmm69/89smTNNLjplARf
w42dclNcUcKKpUJaajyxKo+HMmeYdKMmrnnSZx+zWnX4XDHgwQ5FT6TtCO9REgfp
T9U69udd6eTspCFyEonyhzaJOxCdQx2+4bJK82i5LKXf9Gwulwtk70SpB2iBNXKR
WHnMvV0cDUlR66uVkAi90EavCQNtP42zHnZ5Hqm1ovCYn9ZrhlgWvKWW4KvgLZaF
b50As39BUyblt9JSVRxntxJdtR1CHx8lweZZ0/ucohZYbNd6bLzNuP0KxpC1FShg
sUqX6qzo0nN7egrQ/xeDynswp1vVe0sBxgIxi+xg6fUudA4jwwnHt4ffYPy9iMRG
pTZG6cW7Th9DrFOEGS0BJPlVc8mmDpL7+46u7JahvFfxC+1Y4SOh+1+IUZ7C3S1L
rUqo2NPJi46MQWaz7QLGswmqEGfL9uZiDkVI4CHXM3ODJEBjjbxOuNyvtzo+6YwQ
z55ohOQMf5AN2gWjeUiBrbteSYz62p8FBWW9YDSGrGS1NUy1LopZq6nv+3lKNwiN
XEeVSr1SHJ/ogfj0BjD3i89TVRQq43oGVP26lT4RpWMI5C+5JcO5IBUPTQ3fv2dH
J62r3roPJL8ZdBqro36kQdnVaVJ+K9HltunT4GnpeNnIhDd5E2DYI+Ok1eIfxyHM
tmfa/WzjPDvyNS+dYjpxbmxioOoqhKg4VSidNiENfIthK7j70u5qlKVEK60DQm7b
0wsH5ium0aEflS9XnIdnwfywhraxoQ+vVn5EYhK2uwigdg6sBP3GQLnQ3QbK+XOy
78vATptyXvCkzLNYeLW7DaohB+rdr3skgxgyTq7z32pWU57b96BEkJK7ISopk8+J
Q204c7Rjjpw0DJadU5Fzg9znX/DN3F3l6YOWA4uoKOSdPjb7ZFG06LJXUjFheSyg
wwyuHwOheVqayReIWn4xCnZlvD53WpmHLsYva9+oHKXdgaaIArpEqTRDHllsZZFR
eRNSJJ82f1IIHP7ZOlqUBujI0fyEQNvsXgwQJZyOb+phEZ5bd30ly0BAL2j/Rhi+
CHCwDMYObzGExE+I44eYe47ebRKXGVoN6chMoKcfjvl9UZkjKnpk/2O2J7mb/ZDL
1jrNwtv6PPZXitIQUqHYLfxd3p5qFityXaI3wivjA8G2c1k/PVOT1zQ2oz1c8q+B
ouR8NsRGyJ05VS23lgElskEHATVU/sFQfbtxPfORCyVJrELpgNlb+rQeWD5b1iMp
26MiBhaJb3+7CMNK/TQe9VI7u/n6wo/zXQ2DD25c7DUzr06XG3oM4zibH3RE7nRm
nECeBK+27d6AKxNIKVm7cWG3p4ekIEe86QfEQ3g/rxgXOomAyIXk6I4/b3v02W0T
lk+X+wMshEM2t4GPEDUi4b6AWxYF1CrmItOSSIEkk9hkmEe0OUxiw4s37W89PDoJ
SRoAtMFNszGmgYXaBVfVysxaNLq6bMAPL5UV7ENMl1U81MovO5SNgscmybeQEIbG
tME/8VXu1XxxBLGHRp3A3D+BsjPJWgt89TzV/fycaqXts1TL6MFDG4nTVCfxvptV
QVZ7Ajj+7KD11kFTH5u3BgZ+v+/M6iJqceDVFbiFZSK1WWj2MgAm/VSrzKiugq7W
aUUhUA68RK4RCbddkVReLIWA9mTQ68dEV7e2iO5MH+y0xYQTHwqa1839EJiGqy6P
W5RbWxnRInPvOUk4iyGRxRnxEkGua79zF1NhYX8SV0cdYbRaYcGXjH4s0Ze1FS6X
WwTp5108zbtPpRIkTi/stwkRHZcoKiHhN5kacCHTCTyEfs9THp2ZiWSeGdjB4Ez+
yiVK3e1XwAw3Fgi4JB9jE0EBC107XkNtDu565YG4KWuDLgx1BGn9kmHWg9blk2TN
LlIh+yqiHoazJV1Pi6dtmYEKFpFtb+155+evE3NtxNlxcOG5HAkqFnfN+hzTaJI9
HmYKqBZMstK+EJK5hli8qGwCnIfJYz/jvNEEXMbAHkpBolEhWF0UoQWuTWyKYBpn
L144gYeBuX/kj4HkVXyAnc/TPQZBiZjWmPAQ40xyaP75v8Us4W3uWKevhcSknIoR
vJi4/x7Y6b3XL3FAEyj1Ce6bO6JvXHaax6x40zfK8coMa09afbpYy3tXDzYnZ8Nq
Rmn8hL0SHCSy+uk7Wx0YAUlDKcHE9Ads9jYTs5nofW3nxM1M4sF6afCjANn7Crp/
NcUIBkNbCE8QlqPtug8ipRSM7AhyMvJXOgwU0/RAwojbhrgst1xeWvXRkOrw+XO5
6aEDK/eHIer5+vUom/vHQ+4pFhNMKDTXjABp0iZu8MflkkSwKGPYONotnd5T0z42
ov4o84N3ffoq/uy/WoDFmeE+xmMXz3tSLiSQ2VsPGgi8MYbUMfxNg4VjZTLQWeUK
5K/iWF0QPh3CWI0JtAgOe/oRdmFc9IItJusfl3Go1Shfhpwi1wS2Wrom95+uZxkE
MOsllM2WWnjD4I8jzHGZk5xlrFQxkVxH0Kyq+uclGccx7QRwgOULuoQXkdUWhn5d
A9vZl55NLjblzECg7ObrYFdWB4OfdG8Cu6CnRtdzd25jxEjvkmQrPTZh5os2CXwU
KvsGpUH3rQkToCdCOZ0JnlcYWG33w9DNCvUOs4zvMH/xb1skMuKt34nt9p3/Bggo
y0c4fZs3yLHEVUxTMZYEdkPqz2HF3P9Zc3uSef9/zxEm7DjEMRSetI4R/mBw/Fr/
V5RFotBluuumXL6ZWXq8Rh837780GUsTDqtuBYVhsHZp9mmBjjRmQSXIh05l5rUK
eFcAJY9mdO1xqmQlwdu5V3teAy0P5RMgMyoMUXDb72psBSGEVDbtwsKYHO9mM3ao
rQ/SjA6EQJJWLBWzkO/XJBV87GXXfW/uhKtbbkciAmhgQdFoWsD93JnbTuPS7tGe
BisCRD+TZJIGzUuGYu3IoT0Xjh2Jf7QGLqTxM8ZpRbpoghS0Vh7FFwxk7yb/ezOb
Ztt/naIQll71yEn8tH03vYxFo/y3Y0k43IPio4s11MPsM9LObPujDATrgD7Khizf
DcAfZKoLVPqNKiU1znVhowdLyKjgr4Dee5wJ5Yj3RkD86pi/trWxE7TD/sqFHaTe
F5DoLtUjDzx0yXj+QuKWUujhL9VsW73l8FyWucFbDSqnp0WLEEkJjWd64BVYQgWK
c0+h1X5KY1DJ46SCPI6dc4JY7Lkg1SmbELyQqAGyt0MeAvIY4OzwSCHqdX1uWoXd
RKwEhx586BG9zGee+X/6JFLy3Vgf6rhyW57t1lZ2emg/+mQ62rmDKUd5FXl7tLjv
49+hKcUhp/PPOAdU7eDHVfm7vhPy7vVwW18yl7spvLIIgoctRU2aEH6BcD15JkvP
iwuCvV7IoCoWs+a2Z3v+DAZr5D0Vo3JI/NrHomy9bCs/MJdgaqyZdQjW6yXZMrLS
vmOg45qdFRkCb5mlMG6do3CSU/HvuKsFPiyTQd0S8dngeyOYknnXzeRfJuUbm68m
acez4H+xRywsRoots5BV4Ya32UGea6CxiaXb7Pi7znWlIq4PbyzRit22lLoocTq7
f/xlX3AmXkp8I/X2+hfpm2LegA05tWLLYtGOTPn1R8Lnx7ogLnWcsQGGbQ0XnH6y
eh9P064iO47F4DSoYvfen54QB5WpgzCGGTYN3iOy+3Hi9jiBlKiqChe2Cmye+5UE
1w99ZdLC8eluiljCmma85EHgT7PU91Dg6dTLv4eWcT9BTWfPFYJCMRG9xEDyDEz2
NwwOMsp3Wg2VTGiAnSdsrAssNCYiqJZKLy+As2Ik/GuupcTfWlHUSDkJSYWh66SW
tpVVeUfNbZpOhbpYkbfGXcOGNA+xegpaoOMpkQTRNz6ioR8kOZcIAmP45IGI4IxF
l005kV9nX+dxYQqHOB06nAuC/8YlNAU8bZdhrbxSVi36KfNWEHQdFBK/d7e9YNuo
zM1RD0r++FWYdsnYhzCTaZbzK5zxhhU/jim3Nuy/85ywT/EwmrMyt7QSW0W6Dzbp
of64kNDCW2Ba+BxOR3xTU+yWGFMIGgTYmyUPeuV0Xa/m1c3D7wLM+qPpvAbOJ7ug
sZRlukJoFIBVyWHCsaKxSCi7HjzJ68pvZuvEFSs+fbpSLH9hdWip0L+QfLn/welk
JgPgW3fO/34RmWdVL/5yRUPtYo275NEZpqk7FqZRM8Tny5CK2trqacStW89PAHrF
EvqYp8neywtN1a3NtFsqCDwiHbMu8XbzXkUTMPRDSfOdzCJRQc9FcgzJ+Utg5M7h
yXNUgkPUcKXqNFm5cgobarZt+PXxMLx8jHAr/kkfSg1PzjTxX5QLrls7u+PHUxJv
I+yg3xuoLO2wMvVrw3CFXZ4B2i2Q8twJ7hOiwAB1gxg95sEON58mfJKkoaaTKcte
6twJrUZEMuhgmVTG6vWAmfgfNvnxaCaFSOQcV0jHMB+nqrZubnFGmEcLWj+ibiA7
acjxVweDA6oGV92qF8HSv8ixOxp7GiFWo+rWPGEKNXik26cpOiBZhgzmxk5hb9Gv
NmuXYYs70vefmZvqjkZu3CvDHH2Q8LvV331T0JVshcOSxVBABqpjueFrd/OCfZXs
Rb0xiQGoBFZMjlMhs8g8KZRsv2k5aW329P2jcz4DDJqP6/6FM8Ska0rDjEq9q+km
SjM66zj82WbQmnBOQkSynZtmd84N0erAt5jD0zqInHqwV7z0V4FYlom6MeBEFl1j
Dl2tF/aA19rP5SJAJzUMeY5f5XTlmEvjDt77i3Csoz9yt77YdwK4nDuM3R77Pl3+
tMj7f8n1sPlo4kgabA/2xpC+Pai6gZGy6YTY0Z7CLTEDcHqK0nt66dOXZ23SFLZd
TZ5KWJy2bkw+vpFxx9dWxzjESGKoMBWmOgpnZNGLvA18pUTlrwupvwe/4A3ulr2U
JUL+iarTkG2/0BroLb88bk+d+pNFF8BhhA8z+bjy8DPYrrZAp11ipTLBf3+M9MbU
B4hFZX3JSI+8Hkl32Sm/zH02Y8hj23vR3zgKhwKE3QNa6/b7h0kzdLSUGQi41Lnz
hTpd8Y3Go2rMjOECQ+WF4s6g22ECtvm0mkETN8gEctQ/LKDUCW3MGbwInhcMv9WY
IbvNQkmFK/LKQXeXWWGLzV2jWWhLwmEEbJnOzW3fLUhyFH2rdPF5t9Plj1hfZPC5
S/R6lTnX1UyNNjgHzkBwS3GjjpGSjtKYzRcN5PKAzd0Cxg1pVgAP6GWJ9Af9ACFj
FGxoLa5FNPMoILdF59cIWkxMi72Z8Q5MLcP92pkT/8CbmVh1OcqWzUQu3sqnDJ40
p2WzRlfk4uu5+TFQxfwqw9oDlEn3TfX6GdRnF002nw0Z59bPe6e14L5zoslKSYVZ
tR66c2MKHKuIqwT0dRD+KT1mOsgJH0eAyFdLrjhV/pHuhLnTSuBwFtTscXZkgY7g
Y8ltqzDZGpuvQlHEKhEv3zwIT1azVzwt5Hu85YBJz5THkZpY3L1goOWTcaL7IUao
jCEQitinH91ZKp4YdvO7WzQWy7vMyTZmyC3/KJn8KxzjWHvFHZ5Coevy6Q2LNCfj
2C6n5zCJn3f7A+jRE8imtcL3aw2EA7LMwyi5nvbD+pwasJRMMbUM33vu0+p9en9K
32CKPwouq+KOqiaVILOVqQP3cGRjgKqvKmaVKnDJLCMIxccqPiyt7j/OMYQENJpq
ghrrHoi13bqfZl6KpbTghHDWpS8KX4Y3Zcnzb7qm9DuSz/RfuljJ2N70ZmVdXtm7
hRU0KkjJYNvaj2q4jV9SmiEZJj/YziU8EsMpiYJ9Opo9M7LJi+amvhrU/ZNOkFIU
8KA8FHxTIAd0VGdM6lotYSWQDM9Nu6Dc2nNTjnpaI85vKbE9CNV0LiqtP7GL8MVW
UHdeyPFkyvKmih1qAjD1spbSjhfxsmr1hbMGtmf0OEIBLg61OTVONtCPM0rTR68E
wKtaJtRARiJuwa9OOpzuQ4Ga+Q+1VMumea/jtp7nKYgl7GsnCzld6jCYa3vDTVmV
Tz0x6/klZXUu+o6e88Y0vJobUQWOZQkmVG/EA0vB1u9T/PRBsSqlFZEcG9FFPDwu
P1tKy7D1jSe0AT4yAph60j86BjGpss4gfZfN8wPL5tERoq7hQe3V0pKqzyWQtEYQ
m4BT/MplVrUhnftVvy4ocWgKNJpdz8Mf6Poyu4g1a67iUeYdR3RtiszxCb4VxSGt
R4oK/HO9xY8qjK0JAX8Q+Eec9vSow/DMTR9l7UbaRuoz3PBsln3EPbjRoOXXGfnN
cPFxIDDnlW20y9s2NrivHWaUkZb2yOAH79KRax3UUVJDtANtTdTB3IIaAJycHZxJ
uGVBnkP0MA2AZN9pgkoZaMPLL3A/HDt4F/rJNG/Xeu8f2njTP4cDkbO2vSLjTW8Q
UHq/8L3kPTCGjDSTJNkxVp5MXOyPvJXI7Ja5b87aHFbjYWXvOs7lGxbTPGb26eNm
rpoO212+kKrJgFft029jqL9KqlbRMohlyPxEpq2mH5dKSDJ97nQ2a+srWRQnDDHc
3YpQjaYCUycYZUg5T92V0V7dcmycRUaUOgW+NWPHv774u4mJgnBK9rG/d7NzeYBz
KAK10qIfhX2+h1oLg3UqfDkJfeMAcilFA5TaT34Lzp+PbwFKKhFCW3c2JrdvRg2b
Z8f3P3bZ2oQp9jLd48eBEdE9sMgRR3d9gVchuDYvWfvy6q13ixw7QME80tljgzSn
byysPASqSTfwXuPnK4mUCLMZEATRxDeLu1XrP53NfSGkUrgE2UI4IReUl2o9Qw1e
ietp6NlwhKxUTv3NMTYNcPW9jlWzlGeZYg9VjvralscWQsuReUqZXCTduyC16BOj
DDdorHdU7blnUoZqIw5t1DOsD5NDNtScAcbhkBhdXae+lDFyVftTw+yzfcGBUHre
CO6mABX8KaO2ze45YoVsMObxHxaXjWowu3xuzNtxp+KFvVZUKBJfNUukpPJy6ddE
GcIy9qIPkC2eDXExCEQ3Ht/QHeU/YqwE1/nFggdMYXrOukKQHz0VLljYjHnhp6s3
FX4dtPQ7s93qJTkkMKuPa+lQOkfpnHhbMDwtQjZqh72x0SNt/gSMEWYnwKv6ueqF
UIFd1ldr00HsQLV2kQCDVV4ulq+fKUIQb0NABsVxypkQZtfsbQZmLSPyYVkE1L33
eRn9/DchbXTQ7CazkXCDRy310XpWKlwtbyZA3t5otujmERSB2GdSejnytYTjIvgb
5nt+c34YRxQ4cZMq5wlki5/AVXXBqiedpJ+WaeR7QVQDVnHudlnxJROLG0qJFiPb
as9RLSjhhRRGN7xghXLpR/NdCShoga3axzgAg4cMr/IZSgNzgO9RXGg+PByfSQ9I
P78+wciwLQFzx308lhpWB5gzKwkFbaPLJWQkwtlNoVWQmmFgrYNeJDtSKdcwxx/r
f3OEl/Kk8i/+eDA9gYx3Yfg0Z+QeflPtgU6RSJd5I+joszS7Pr0IG2LV/TC2oqVk
2zLMrLRG2ia2olKPFWBcwCm9pVZ0TZSUA0/GbwnbPR8J2BSZ/FiOD42stjHR4E60
1Cn9Zp8dndllXnIImim+NQQJuStevlU30LFa7//RfPFIIUi4dUoocXZJXj5J6mYG
Y5nUFDj+rNjyH8xkK/Sea9S3rSpQjp4Mci5RxRSx7Hgs8IDUsoZ6z3lSUl64tlAe
Mr0zx2e1ecDo6DzolTxRcecc5Ts7oMnQRWjJV08MxeMdutIkjpCSjB84a3x7wnFT
9LpG/ZgJuoAhZyd0tS5oUNcuk/Zh1gCP4YRhibXqRSqF6jcyLm23nlmFuc5lpQ5K
WA5OUuSNDT/Di4ZQqFprO1wyfxrWdzAKHSodZxOZIcIntqwB/yUFHQ5Ldd7oV/bm
Jr1ykDZ5LPwl45BAAgA89ElouP13Or5E1dd9GSc4LLUEg0puzq8ua/CcMT3k93j2
SkgCbodPakPFiviIxwvY8XQmNE8VKBY3rtYwow0VXzZQueeY1nlR1RUulRuD6rAT
hb6fApvNvqg4BLR0ZXV313DDsO+zZkLyfoCGznoUPwcz6IoKbGjbAtWic1vRkCcJ
X9wmcmBxfXjDnPkPaZYQ3ndIJvW3YzzjWvWZqK2MHm8xhxZGmwcaynrNpeneTxWV
SpfWIYHj7rk3zDZ1+NlCddfxCfIo+NJ++cATtxOqMe7hqfeqD841WCM1xX2TGu7K
fMJUppeEnsZlc+zxVlx1QBQXQgyazZiB83A4ZROB8iHEDF9UjAMkiio+fPF6b6TQ
Ahds39tqtt5wJjsSgbp8TWU2Jl2z3j2BTjcMZD/LybXXUYstBG4EBLxsyq+X0xi0
PUwSu7w4ZFZQ/0NrnIHoi+Hu37Oy7mz1sCcd1nYPPETHFV3Ih62CMfvYsoijpb2j
7FbK59WKQ/s8qEVY/zV1OzLaHKkpY59iwtOdjnKxXKcOq2pQ6knTEJ7v/KF1ZKmQ
w5DoSIjTRJDZmsCiFZKcu7KJEA/3tFtdpjCTMaVJDdt3aq7Mvk0AQddRP2i9fHIw
tft9RPM7H9NH4mlsaCZLkXep/TcZBQKceM+U2L6yk+XvSaOT1hOrn121rtOIT797
ShQmowGRo61REQITtAw0TsZ07/fHT56Z2OtStg0NDeBG01lUsOzxMz69+DW4pB6i
vSkET+6bAX7pC5boOX0zUXMVn444lYKr8C0RxsLuC5O6wcCPw2cS5T/pxfc8qbMP
0HM2dhFtQ9QHOpTxFVz/GyDOyjxzdF+zIRqDcQLYfT1ROUOC7/mFaJZ7BO/Cdvqb
5Z4LyPenJSJoWh61C8c/TRmv6XTHlzcCmcVM0S3vbDd6R8XVVwXdgp1k2OzjwFRk
WeaAe9Oel+vD7lqAj2ljoNvBex8Hjc4IiCGk/ldpxvKQqgU/dGDhc2ZaN6qVL441
TCBfV8Rdvy3fvtOPksvVUnCwhuzU/1I7R0kiB+o15VRZW6lFk0WeinXlH+0iTSzg
Vz1RS7R8w0AwnY0PvGurnAxUqxdh8pd0mftfFQAzaHn4oTMvEKineAQUKpsWL2U2
erSYGR/Co4FN0lDS6s0aTBRx8X4a/XWmQ35IN01spz/GokqUEv8XvzBbwvmVS9UJ
Gk6NiVT/sgAbd6sh9JUeM5d2jwTGIxfWXBlQ2lBRlQGflFdGtUJLJlY3gr85oCRS
8uhc3UlYuL/8tUs1FSexj+jvP+Imj4xSxxiixEeOo02CjoeJn0TSYhqAUtFJszml
lHWXkSldtbPREHeKicC/bY7PiL5I3TTBcKPjvT2kFWD6vwe3jHenUPyK2469a11V
kla9thF8G4yiucnW1M+UZ5i72hYJYzm+PPJap2C1kxh3FgaA78/Uln+RH4LhLlsx
LXAG4yi7yWPSNESj20o/FYCfuWHEHB08Y4cPrA7nTkvxDEUQLuP0aOgtzvJvfbOR
sP1hOTIb0DEJ6iAg3UhXv0zdtk26yGtZ3gLJVIzflLB6YJG/ylkJMa6g/cVM+njB
Nv958AzwVcKAeyX19WvintlaimvUhLvUwpUxaUj1lWZE+iIzUeHnEydr1rGKGq7O
Cov7A4AyLt5wIw7fiaa0hIi4pWXUrGmhOBc3Vo9fY69zVn4gK+ncaIyNOTt4VdFa
f/JC6aE5bJn/4qjLitwyZbZEBSo12Z+c3nQ9VX/fMnWNsl9QRSBvfQ40xyGVjnLY
eQsSmS1MPzQ1pXC+OoZ1/6F+gkXaSEYdXMuncfr9cBPeAW8e7DmCr6vIFLVHNF8u
sYuRP7dssNnHQ2oWmZbjmzS/KVX+SR3WXS0mE+3F2Fupmd8sqI17wucWmQFtK4Yx
WvsI7qrEi+0RwJ1mJf/20zgaag3g0fIkDwF3gU+69j83dp7q8StEWxXBPo1YIP/S
Ctej4MYFTnvnCKOPxYv7ORP3C0u19wk7mwFNmNG3wYLRb3cAlzSbWnYjyla6JKql
c2qvFdxV1RCE7r5wgJVnUfhY+dsHbay/L8BNZpLm/QRK93Or2Sfj6KF5l11WLopg
NbJrc0CCurUkWruPIJbEtQ2Qd2N5RP40CXm+sG/jjMh4ND5vITJ0zmccRc0BoHaj
c+ZmYjk2NXlRK8YDCgsNtDzc7nYgMFEUNqg7E7Y5W+u+qQpTAfAcYdoigIbkIia+
WDpNQbfDOexZTJfdd3/ooTR5tZcu/DQB6ayTFxfotQlnkHhehzUdPZvsuO8P0XAb
V/2uf00y+sWPcXHQt+UXDX0U6s3cmOyE8V8fJxTwd0A4pe/Z4DRVYuVxniQ7ckN8
568mDzzlDXJ3z9qsf0Qd0VRipaiUTyNXadrjCvC8tdFbBk0eK0DV2P7f+4L+32L8
gCE+Bbf2tlUtsXOS5fXXIlLa6Hy3RWuu4X+Ac0A/ChT75eDuGJxZkFB4qpL3fa4u
2k/t/k6zgt0+k37DhViwxLtpcXu/szMrZRB+JmmfjEd+HeA+ruwFDLdgWHyvMeHK
/KuZmKYcQAG9erMfpGt8LYzA7c9UIZV/8YmaWKnjoed2748zZj/55Nkgo5ZMwHPm
wwZE+sjHtacQD3Cy4b8X9rqyQCIyySOoKUwNCtFUQvIJMkGAX/IOFDWeq+Jh0vRI
B+6VBzC/w+i7EMEjDl0+tLGQ9p05w4oayaKhuUOfjr+YEGrqvRFusZm7XPl/mrKX
CuHNeVoy6L09SV8tUDh8zMuFvm/2pCeH4+d4CgDH6Xr/YCZlckMve0Kt3j6YtrSZ
TPqBwispHajPncEX1srelkjQR6ixyyxJbLckwQeYYvCLFPcetPGvj76VQAfYkuP8
Fw+62OFgeAUKDhZyFqAqQJuboeCNXph3fTA0iofpgaBPgfToZsJ9fhk2yhFgHp9M
5VB8pVf0mwtf6S8Ht0V+pAl8EGpIT9+eBznO6RNYRBTmCqfC5pr7LZ2p/Rf4lsT0
PekitaIZf8stVYC4qIoTRo7kN4OHL3oUlz/50E7gEvsjlqYCs3hT1hBSyaKjPpsw
a+E23pq2PeotpP8rFCXotel88opvcjQ/8mZIur1Q2rmY6xtsXq9gzadD2WPCWz3f
iyC1/dZbAxmlQDxKxkBZqKmuPJm6zlA8R60WhiyDXntP+L+xIDr2b7BUJetKY//M
4+6U7zZ2GWh/W6hNy4VW5IsUTb7PwLmHIE58P1NHyKkgXgVf44PEejrXHsf3WB/S
jvdGQrO0QJXF7VoDjOI9iPONbTZLgEisKv8w8a/M20Ut67VhTPOnV/xcMVmKfp4P
4xBtvD+6+OHyNZIQSCxrNh2tK99EJkf1KYxu1E3UnloTUBaBnKh8BSIksC5cLWzd
/QPV01KYUzJkQgcCWXcrrNFlAziajqQmRgOPa9Ejj6aGseeK5kHEQCJ/Iv0QrXBd
+cu2gOYJQdRFtu0y4eD72AWgtiadVGxCWqJaROeKzHHWuYZsblEU+DmZBddo7XoL
PyVCLNgl4cLLlLXn50LzFWWopD8gpl3Cu+4OVA/P3gsStypgKTk7IiEa0y0kXrGs
v/pfVUojoJSQmxckSJ1/Mp23gXulPEHN5pT7+4/byKiX5NFbSMcbxVYc/7TsNxl6
pCAQSQ+3CEHt9+JMTB+GJHNa7TJGVbrKMJfsl7GW5ijovDw8ssFxpD1LbO53y43a
+RbiZQ13kl3jGmhcte3BZy/y+ixlwiP0t+OOVKqJUo4gGv2q2+FJfYE8NtYkJKqk
vY64POwpc/sBFcLUyHws8YXNAvUwaFJoJtDBkj97fzGzLEl62Sn1ibMpwlkCK9AP
8PsPWuxd/xh2Lp0IrrOkKDQvSgggytPAxC7IhOd079bVPYmUyKMfYLJQ129fASp2
D0Wv+EbGRjyHE3Ovj/kk7QGoKlysNYGRWt1FH415kjvC/DSl5dzM+eND8aLVrqJ1
jWWobOs3Ctr8uLyjhk/yPW2Mgy9CgLfo1kfPKpTGRXoWW/MBCBuDFt/BEZJpw206
FQsPqfmbEx0yAVX0lZ+boN0vPXiiOkYdWgHEZQ2Vc5kivJj5ELixqV06HNwQsHxi
2gJwDNkpS7go7OESYJbpSdqSwr9iF5amxvYTGCyqLZTHIK6OwRqYUS4CUDv/BUXf
Z4zPNN4GAB3qEt47SwXsht4R/e5wqqWv+WZss/5Mn8QNW1qFNX3ZoM7hRH390Two
RvhNgO7k9tGlbqkMuU6GG0vkWF9SYhE3+//gDF68qAAcuEeNxzJIrodZlquXlc5i
QSS0UFnasbdDppCC2rO9w66E5W1nTjBMZ1GkCJyZUKGqxgFSk2+Wx6pX77oazEpy
8SUKz3s3WkRgtebQqgYhWZEnE3FCMP1uHc2i9DLnt9YGkvyDpm7GbxNeCbkwgsUI
wErFBCTOOAeORtKlu0wBw/APc1ejD2AsjKM2PqUdqyK3hmZnlZUnI67PNAcFntj5
kWh1KditCYihrtErgSNIMgf6A0vDun2ATbkJMIRCeS99A8JJyGduWkpgYExPBxh9
nuid6bARJt8WXh5dVmLWbEfgU1kLeZWNcNLng8w6UEaUebo3naEmf4C8RUx4Zawx
1zuao3mQCCVzeuM0JSpHsW1I/s20ZyE8gGvqBmpcPLUlkJ58O2+qR02s4CyBPXqK
/VBn8P8X3dApaIn1qchlvl3xknIgMfMMAyKjvhgvR6I1IBQqjXUT1E8bxFodNLFS
SwqnDzi3hGn93f9W+alP465OQc8DeVe3ea0vtcEvKOCg/H36CgcGZ/8ImYhLqxEl
qG2FCIUZYRGp5whCcRgWTtCCCiNmlGA9LQq93kwiZkjE4G3gEQmE1Ld3MnJoGG4O
e6Zcg2rxOhZR94EZmHfyOZzEHJL1u8VWvfFkW00AlZggrHRacDSWBdmScGAppyAe
PW4yBcG0nZLq/pjp0iE2bL/nZdyZjP5tAiDIgIzNSz6hlbt77JKzep+EUsE9SywJ
68DfdruchrRbM9Prv6tLZyEBqFw/FeMLHS6+Dnlw17V9lW6U7D+b1oS7gvSBLsLf
1rRKXNPcT/wvM9Lqx+0YUOgjXxwC4t98T1B2sdGfp8Cigt7YAm+sFhlilRvrs1Cu
hyyoG8HsCcJbTGnTNB8K4GeUT3c6nyz0s2OtUyJvKVL7mEQAWxWJJJIl/zxhOIbu
S+cpLEk5PP7B+2xSM2KPXx8dEx1OSej/NddfBO9gnwcWUWHmY9TCd14SrtjU0Vb8
pEcQoVSSkx7zig29OUWkcPdMW/4gZpw1rRxLDa7iUqkSPUrIHQcGlYDcVh9/I515
zHgDEqxgyRQni3PD3Jjr/si3NLuMo9KlAXL1au82ZDSDgKLtpKe0Isxo/DNPPhZw
XQDoLqmpeDOeJj718NPF+v2irsIZM1QkRjQE4oHV0uGQH/pt5MJKEaryAk0030P7
n3ec8UaS38MlRWEbbAB7aMCr+2OLObIXRwsJjPjJJPTpJHK/9eimS6oXapz4cBBH
ibjv/+zKiuzs2dsGEOfV9gcLTJuRNVHugJiP5oYncVxxaW6W7YNpfD+kL3sBirFW
u/s5HjC6VO5d+w0wrv0QtYye6qgfks+mQ/7ywcJ0fd8rVmdTkznqzZmWULfutydV
YkH+BvUtG1CTSB2oBhpPZPJyvp9dWPIkfY1bXv3sxkMkZZO4swFuzEER08uA24dI
YKLyps4hY1t61vGXm8gOIn2MEdwvloWkdLzQNKxm+62Tel4IGx8Yw8LS3JQLsPEU
tixKX1GeHXgor3m9SKM40w3ZwD4aRycg3wZpdhODITKfDNuog/eJdDkJeoV8kygi
gJtZ4XvjE5gd7eXHjbVTQXjURnUL3D6ROl/HiYrilxPYQ9gsRRPRlkRWvM5JW8B4
UMkykuo2HZDk+Yr+4uJVuxXMrP2607vQTekqdtE0wVbnToP+6eB+HXL4XJ3H2p3l
gcbzJ3Q2IhLy2uYNYNwUlN7Yh9NSDELO79kHE+PXrXDi80iq82E4x4qc2rf5dgBZ
kuD2dCZiW1FpCSAuu/7ro1OfOgnM519V40baQQsENoniZetjcI4TwAKO0EDq5Yhs
I1D3kErOHdCZYRHhvvKCW1fguH+rZUuWSXU36bCJGumPQ/QgEe4RtIFJxtclDt1I
vACOUIMfr3DjIn8p+YvBb0le4QnMHXLGG5L8EEeeDqV/7UxwrPYjm+NkKUJ1Y4+4
LeKiHF9E3fwUiacnxFpnST69isZKkIhosQptp9evbKjugiAKP6Q4MkiebmtuQCmz
QQwsZkefHcYTOm55fYH5yb3pznBM90r0R4javwbTtJHqjyaJF+sqJrIiKAAPlfl2
E/Av3Ojp5T7m3fs+6zRv9v9H/Bfqzo2gdQ67+p6iXojdKng3DiK5Qbm2FNMzbY2F
myDsI+D4hNqTTTEWDGBqY+K+w/1dy69PJEjFdqP51o/WJRan8KSRb/z0itdtoqfm
+y4declAqL7S+xDXIg9yk/wYgdzyRnIrliJvwkeE8D9kkVxelMnaGj8bQRDjbg5v
xAB1loAoIRLlsKG3wZSfIZgz6sX1z6GcqbOmJJyvVS+nZXP+X9pm9roNuRzmbCDS
bHPMPrapqaXLXpcYqBChAyTjx8NqaDVOc/bwJ9AR+zmhuYpLvuk3lGgQf5Yh2Iri
74vs0LKRCqEfiZ9DCmzjJYj8sy0k4AwJNox4GWsyKmA2bkMc7f4iIxLElIw4JyWO
j93AO462l0ab8TnKQTfkfkeSsvV298C1L9akN6ypAVMKLq6TV8kLP2nax1dHwuUo
lP7jGzErlRLMPsvmj8qjBWsN/n/9PWe/FEVwcBqy4OEC2fpOo7pIiG7DIeWQGpI/
TIPGBe/C/EQkZcw+D9ORhE7GHLKRNGKalzTAQt+TFFEBaDyWYvboDTtzBIbB2j64
iRQH1oC64BK2LJ2JLPUg8tiY7kHT4QfTIvdg35XG0fPtL/QPLfq+Lorxskse3jOe
ksn5iMrsgSx2uXW0bZJuf2hOpHHLXhH9v7nBduW8HgW9XAgWh4aAlnkA6sC6RakL
bRwUubZJKVKkD1ASiTNQMhKQuozt6RwUrWGrABccJShlWVvZ+cup2sDm2k4InTm8
05HtefTgApR5+0eBzeHPeOHA9Too4g+wz/u7DYRKkvSHp2Peuteq7l6cOd9L/dcf
Z3JdCMmW0maoKjRgM6LiM5fQPkAqCHqcv6iI7Q7V4Qi8hVkzKOECe9S2nN3Oszt9
9TDZZKqDFyxiUqA+nWyiu/PuXh60C1slDxNt+mxhksr37vfBt7vvjQfMQPebzAFR
XG5eb2ZnodF/MIFiPI3ff34ov2EGp+4+qlgbSvKpHB5AzNEbGMgLcBYL0gEUvhdo
AhakX8FGjs9gFOdf1yvydBJ0beKVf0jRQgmZIdfNkn8hrWGaiGvMOIm21XAJzB7p
eEBudS7wcprfw/NhBYCoSJIwMkCXsbvzeDCfzUYW4ywFtwCxZA0bV7AqXbBIvrlm
xs8I3FTS69edWbea7EVobp8/P0ShvODM4bMbuHV/z1HJeuZLy0s6ch0KDLBAouO7
Wm8VbynZDfCr1g9+iCrjChgBq/+70FBhls0tOZiSgYiv7RdbbdVN4LeoPrEYf/a8
dJUdJsdhIX+k3K0esrc+o9cuNoSnFELbKSjNxHq871WPyfQlQGHGygDb2FQV0gor
89bfoU0HUe4/wG6IQAjViDoF7Mi507/E+ZFfZ81+YOMH8zTZvFe3Z18ZDWx0iO53
DIl1dtdeK7y2uO0wMhA7u1xDm8o75BCzEvKRUHJT5x/xTAWnjZ/HlLFNTLleIva2
2/DR83Ro56XTbMPpoZPOwEKqxc4oCmXK3I5071gASXq1Cv9DzABoopi9vtrz59S2
UdJwf2+dFmUNWPJwyP5xXaagM6n7bwbmxZw5QWiJQphJx5wRxSRDRwyItnbz0gLh
eYRYVEHyX6H9CXbcHIJL8coBYV6yvbq+qLpIu4xnUfPOVzso7cBXr+J2+5DTmtHD
nXzPIP0SKlr+bdGHd8JPfjXMQOS+8t8gYzyLh+e1d+TldBcygr5s+VI+6yWCppFP
rLDtxLKRXhKTBiWpMT0O/HfPFJg7yj6dnZrT0N4IicXndjKqsEz+7bQIxM33URsQ
096Mlu3NojDrQE4KUHPm3WebDU5RTuCiiuPSe2/tqspF9V0Y73Cq4GFdP6mc55g7
xMuTtQoUVad4UB1x5/Ypqr74tQq+w8L8xSYUjpKEwjxy3qgxDMfcxFKkKiz09CGS
AXOdx+uOHId0V4lJD/A2/kJZR6Mow6DNY5XgOlLS21YTz9p6DHDES6oqO4PHlkm5
fV7cQ3ZD6Nc38oBar8siysztRHt8KtO/g5NOUNz6cjDhOwTNDIG8dpmqrnlB+70u
KtdpywK89JGdT2aLY1xor3I7kShnpaxRgZdC/XKdsoaGqV8FT0m54QhyqI5FpMvp
1quu/gVOp8fpIYN5M/JU0spL/12x9tbth4/ibnMoixQCQbKdC3Y6GkgWYE47Hi0I
5xHzRWId/9pci6+OrBUXC5VMXx4mkeK+2G9d35Y35Pjlc4GBAa5bggTK5qOl4TZJ
KymZosrKjJ1Drw1AuPG8cSUsAjySQIANWHjto9yaBDpRp3Ss486m3FMHlzrR4Blj
1/S4gXPI+/wiwEkOAs78yjLLdEVelJo0hXED8BBwliPXo8bED1Ik7POcIYGDT5qj
Hy/EDRKNktd7s24vqZaVdl0yI2NnqtsjtLFibTUjvORRc8HLuwvLpy+b94R+Wjrq
VhxDU2qM0dohCZ2Pv3QofAvryhZQsMyCNsTGvwaQA9DwUSKtc9Qnu10y3NtrcKAf
iWROMZ8Lx08EoxViLT+Xn0mLvkyhawONjQAKcD15OrRcEyxsxQa15QyfetA+eqfq
0sqpyGddDnzlCj2u4N8pGpn7knNNELSPtu35Rkdn1Ue30lpQ3dvQi6+ou/rqv1Ds
d0olZ0oc1dO16oRyQbr5UHAhxsbR08XEK4phIZdb9QUU/f7Wn/oY4RunuFWbfeow
Ks9I7BGaSdRkc9OuIu6dZ8dtlYU+Pk3clkXVosInUlBOujWMQYhBpq5abedhbH9Y
YO0pJoaLC/4NVVxTmZNPsmPIkY1QZlWVXQDt5xmiKF+4TuXC4KZ4mSli/FgH1lQG
7B58GRgniC9QYi4UKD2VKnl0lVpH2g4eOQfaIFRUQtYMXZFvlcEH7+vAg4Vuf5e2
ADbtHDqiIhn7+4XpSzJS/5UfpULi/ah0GrYIJAFBhCjncJp1L7YAVJf9mb5XYk2P
FNXEnQGslpwKDRWR18tXdRVfS0kZRNoBeVM1Z2zeQoyZ0vRcaNq/LMr4QFOyWB0Y
u0fmoUvCuaD2fO6D55RE07E0ctu0Q5TqKb8TokIr2xu/LyR8R34gavomAmowMNE4
yifhzd4WoTkhB2OEm7U+b8KFoKjJIrNb6VlWuMIeUSznz4vV8Hyp+XAWvllhgrVF
oexUrE4LANgD+HZhkhCH+La/Rpv/eAc5ck05dLRH3J9xtPQz4OvEQH350Xep3cIH
n3HTbn3UHgMCpAdIsY4UEDhvTgeB9kNs7F3hpgzcVS1+XWvqMmiy32Yccb5M5coH
gl4/FsF9SOcNCLGqxYEAwLajryMQ0MNB0HIohEsikfIK1cLgt1ps0jSbU9xt57Qd
YB2KW9LSYz8cBuMmXuAih1lGPX35E22b0ipdQuPqI7opVMgBknPNhbfEErGQGx1g
E1EQJAel2Gpij9a3WW0vlGrgf8BaQ5QvwqqSuXnU00vnZlkViw4VojZy8/T6V8jY
5K77QZitoXvDDEoEUiU/jiMMwB4SBM9NEA9PM0CE8ItQmjczjkX0BxmUV1tZv3gj
zp7akpsSocHPuOQ0/ZNVn81xGxGePQJ2BQxveq0T30liJXAuRYwsdrIZMfGLjqEn
xFxV8Knb/ZZLgmmlt1ROdBjRhUZfb05BUh9ixCry0Bh0UCa7s/PPDUdS4p1IOHRA
g8/JlUDrL3+N0Xg9Mi6Exhm2SsNJMPap0/2h5ksHw834Rj3Kg+hm4zAoMHS9y95a
6P3Yv8Gy7F3Wc+aUP5I84Pg4RHrMuQJ105NM7LYeFvTeXcOYKAGceXyVgiRsXjKr
UEw5x4v6taFTA5TgzhofAIq+POnWnIiaHYW9pRvud4z9Td2CwV0qDZ8vAUMS6vW9
+XyJ03E7bRyEY4BS9hjUPZNrjR3nkAQ2YaF0UJxMzvngzjzoo4T+HDZapErYJWbv
QJi+MlA38PoDhYVXMB0ji2xBDKyTsEEPPo7PuiW3vbkqQalZYY1j/5ChCt/U6f3U
WR7U+2RE3z31dKize949lJqHM/kTZttwWp9ecfZ/4PTx5coNHEU+JKWixq1nU9Nt
7bz1zD0rXmHMWTri9X9WX7I+RgXPqH9NzEilyaPjdn6aDMvTwJBwsCFoKg/FGT09
Vi03uK1BGgX1VWQKjOUvm+WskAgjgCYl2VkJiriMgsquUAvSCpY++EeR3et+yK0c
jSDd+bpmT939KpQDfqman76pVAyr/gbVEe4J0ZINaTJinCkqN39Wl5hMIn2Srb1O
k31rmLf4jWZXqy4w0DPX5Ypa1g7wlcAUrTiWfN/1B/VKTxVTxUMz3TNIdPCSZ155
5InooBNbgfrTjS3TwFOh0eLWF91jbfmCJdb9phe8g1yFMxDpvViWoZ/yQI3nEXhS
GZBa0oKeyapgSc/rzEO8ztePW4rQE4qy5Qk4B9amXAKsHdK57atyl5br7A8O3mkH
UNapTpcUPN5xE8zDZ/VzLxI47gm5mJXmamm2KkSddjc2ONWVAwxbFJAAI1Zji4Bt
59+9zrbV0Gt03pKduEie/bMuMG75TGNAEwMC1pRLNlJemW6Mx/2ycDV8WZcAp+vp
LpSdEmlUqQLNBrn8+4MEcmZJAYe2CmiazN1fdDpCPj94YKUMKQaEyQYB54JYvAxY
2yhVSnMXPfUN/4lU7mpi6zXVGq0fP/dwKuns7QgWeCdUxKMrRygucxEjtG5onZfJ
KkyXIEdZQGHCl9AsaUXKJSe5Ve8U3WK+lfq8czbxqEXD2mOkpvJAiVRxx3Rxug4K
9bHeIIKscfwgRob6Utarg43Fz5Hc3fqrmvGHdISWkJN49+/319hLiFk7pCSocwwJ
eMgIcVQEvITYjWZEDKFqKq+1ynLrpgnMUf6ay6Ak0MHKnzi8fKAQwA5cvoA0nNiF
7xsO49Uc6MJcgzqz7kO14l4bSXvIac1OR4pz+LpI+mKK9Nkd411IFNjZRUb9W7Iy
pa4MN7A1+kJQ11DzonkTHpq6h0BEfkLm7MDY9wodqt38cRO353WeIfC3XGsJUWuK
ciN/KZttbFbznqhkXVl6gS39kzxh7+CXNtm5RkoQlFgXdhV5FWkSs3kCSrEZ6GlP
7rwE3gYFYHk5MIdQgfi7nKROoePbE4XShGT96ZqP/j0RGmN+BoBZxiWJBcNtzvlW
Fuwe5OgLeBYz/AMyDevP5OlxCkWEj6UEd+nCXeGhoHpUaCEiL83XaBt/IPzs8vST
ZhSfyfvhSV9UsVizTYfGSFXeCgkqYK3BJC66otjJ9clutpU6WozJ9JEPkaA7e6sr
aMeVbruimpGtwjO/GjH0/6hnSn+icx/Abf30cmRjBibIIeX3md3+U9IpAdUqrRno
ODYKD8dgUPU8JaqnGawjn+yxRznBpg3OZ5lBYN5T7PbthbKgRaPue2SULf54j7Iz
MpEgmKZD6GdE43jHkh/pAzsnzWRbitetbUnmhJkxHA57CFY2o4K7vqjnjD+TNNKO
WZkQGhpwWW2I8ppiaHfZHy/osdEvLsiGO/XHgXibnALsMUvWuIEC6cNSKjMNqPue
a1lRjCP7oA+CHtpUBQdUYPXf9tnZQYmAZNYsdg2zMhKgkSH2FTTuA1tF5u9cBQrs
Gg+JGyJBCsl5E4mCPppE8hVUqezWj0VrQeyUtq+i9CwwaiNkkBlEj7Q3S813eWkp
CHuiF6AuQfQe5c6ftnsgTQr8FdJzBBoyJQERBjXW7Mog3+3udfusDhJCLx9ljR1U
qgKyUMqsQul/CZYHD0FUvz2u5BIZJRzZaKS1znb12zi3qkwK/J6TNXGWsVtu8Gcj
fVqwBcEW5z6K65bfZCc10b8liFx2XI7cd8AWR+bkFAm8NwlxhaaOMpzip5eUXwN9
SmEu0xBNbxsS3QMtsRX/W2skc/DeDZVvUuQH0rcWwdjuulECZay6ZoF92B4jH1xa
cdKPS9Q5l5tJomEYj1hcdW5YvqqQCzKKLciJkNNqyr2Dq+JOLPp8dU92RmNUfMc2
6empbN9yFrSw8AYAinzXfDAkWwmQH6zTdxSWXaIjYMU37/oucHelD9BCyUC1hVMe
ck8gls8mCW4f7+yzBgf6hYW74/lB+IA2W944Fvx6OZLSbDZp0hXbqX3UwWwy4t5S
n5MX+pbK7LUDZ6bPxm0aGyYN63xGGm4QgU21jbbw0nTLXnQ1ZLIGGKoIeBk9dUp/
wGw8dO2v2r1qVn0dImvE6yABs0FyT3H6hBppA80yw3eSq4Yl3ZpA3iofjhj6R6YF
NARM0+4dhKZ3OCa50etVoGPPlRC/5AaZurn1q8yu6n4uKwM801uyIXTVVrHFWA5O
FKoV7wVEU69iSxnfhjZHhHozUbc3EgbEWtEN5n/OESAfl3lOoNoXt19TKOhUtKp0
pucqs7YA/vOS0KR+qsWM4k55fudVQp3jAA1a/Fy0iSqsYVL5D/vdE00Xluk6hKOu
gBUz2lslhalnnLYWL5zBDaFG+7AdGprrhFgnwBrToM+YhOlJ5Lv0IB4x9YXcrzG9
YSI1xHGabgj/Gdh1RVBSOze8z6CZsiU1BxrJNxOdheHFakxQAifqXwVqKhfY241z
8DBjwjsBDiq4qyVFbGbPEmkjcyVkGvAJCeECqfMf5l6eM/rpdeL1jgLe6A9L7cBK
d0bYrWxCkm29rdiX+aBmv/ON38PS21LDXkooEivOdziYK7bAiArRHZ95/0R4iilD
vS3ib9FtFOyoY2BT6FAe9/vHnAXwqJLxtCWW7llwlLpdNioLysSn4wEsUMczJ9C4
sjlh46srP4Ic+k3vuk8Au18bX4tpjKmdc6U8xyqQELl04bbyyNTNOtjF4TDB+1Tw
iTIqHE/LDNKzJ7fn33jgDpmlr2Qg7uZclswyxJ+4rXUjtaqNhT3P95W4f0yKJDlH
zc71qnq9v5wdvWKzeP+mx3lYNS7slMPXkZl4Upb8GIJtZGdeotyVgWU6ZKgbaIgu
DYQlhYEqjwnVaDeNAfEdlyjQJNfqNhIYeR8Vxz1pgRsfNnzirY1CN3/372y1kAgz
ARwz/aOLO4lzzAMdrtKuTDHHAy1l1zn9507jLhZXxdzGAJZTrq3kcfLqcC/06wvs
L49F0wZ2PXj5wg8L2q1egOw1HCnJCfmgRnB4e3PzbSFPWGfd7/QNXpUyqBjxcOeP
cYLLzFVNgKl2/EHnrbqLv7Kj/QBRVYfEoshoAgXX3Bf60qFAzu5hdn9n9CEGLbgp
fqdrs4mJ1AXkSFD10kQ4ZSEnirefuVIPtK04SwLMLmoIt+LudBiCR3hQGZoaEL9T
Gpaia6uXvXvoYbFa56rkBVi3VADlJ9+9fM6f+pAPzqRY7c74KNS37wmQ1VZXKN1y
X+5B7RIsFHjIZTKU45b9poa1Pp5Qd8B656CXKIzfm1oj3RsQ62fIVyKLYdOtDgIY
1jlIGwId3/o2cfB/lGVjntU7wGhj9Wvoshpoh6YifXNLgXFo2NGUwDIzm1F5DsFU
Lpcz365tuB5SWXLCPAY79btIePgg1CFE+hxSjP1RyBQVoRyLFETlsF5L83qoPQOU
3pML3ZJiqSObZ+8YxvixCyHT+0KtGcejon8SonScHbhJTTBkPKVbniAbZYzqekzv
Ybxdtyn9h5zOUpWt9C/O4Kg5HhqaKgabLbItv8nFjovqIcaXH8/ggevzf4oM3Q1n
S8+4BCVKEg3aMFJ73DdguI88PLtdZ1Dl7OGeOgBbUQbFdA2o7N5OdkpgFGpZWfrK
oodeoUV8bwy/mMmjUbx0IBpHUKSkH2kxnmGsqrj7epdPjrSP7THJFj08gsZhfVhh
NusIf0fL4PK4uffopqaCvvjFlnZ0l3uS9g33tBzovUJm6Jx2Hf8k6s6UE4xMNcrc
anhUVBT93fA6nLl2Q/n/kYSndXFlu/MhtoGscIKsIc9vQq3mGPvweuABHNhognIF
6gt5588PVwzlk6rnItdUMrxZYzaNXW1PRUplj/Dckwha/W7LfLuLQ+qos50T7RYs
JjaJd7YsDKRyxh75Uk5R9F5cujmXhCYZqz8RupAXbXcf2SscCvI00Cl2w+Iwix8I
ej7/4mLVkjCFIsCPbI0xyqwr6sDSmPZhOJvTcfBbXpM4TYbetP0Xv6c7JdGxlTMr
UahM9vdSd4sfAAVoz3aOcKfOtJLxzWlFWMoHfrSXMQTkfLu1pXEur8bx1AZhnksT
1Ntj4IE+N9Mlt4IpjgHnc6fAt6241Fad8GPbbsw2jcF5JocpAgYp36LibQEYeeR6
01bOAotfYHZS9BPlmktHUID0KioekEaoSc5SInJmX01wf9e46Z9lKnJAHKihL7Nr
EGOLXkklb7ne9cK9vYismwpoJTKn8cZ46P2YgeVVuoCE2BIwOOdcSDYPusNUdCpk
8SIPL3sVXb6cpFM4IUdYMIGtcNZMOyMRdhj6tduIlDXXjqlktjPq58bZRVSVoLMl
uE5vfEkVUFvGMg0fGmYECmP1zgmcXY2EDpX4DGoLQLvjzJiTm18NFwZLe1Mur3AI
fNIZ4LByn+cFp1CCZXBPksNm5599BNypT8W+NhDDvTzRRPVq06jombsEy08312ME
K9YY6nbmANrfGsGswfXvegHazJ13QynSG9UEqZSPrAbAWED7Ekl/jDrOMfwo3Shg
fTLCdb2mrC83Jo4ySgJ6O89HdQZXE8kAKaqVYloy1VBAcmrgsSV1aOzK7AW3YcOv
e+afXmAMXfhCvmnyJi+Mdi9W8Gk8MvZ6yV6qhdRVrkYUYwATNgpn8Mzep1nDCQMq
ziAMAr8OlGnSStXC1fAIOkXElQyCBW8sTEyTllztbd9OWdgUyWoOsxjWumxYNcWq
jm6yMDHmou8C7bTJiQD4kerOG067gTT0Yq+QS1H0VFrUm4fbQfVbHLe7WaiZ/Z12
zxySK4zPKxD9DOeuz4mS3PqP0VTNtoNlRGp3NCOINwAqAUiXFfYDtLu0UmlST1hn
Rf2PhS+wGBFTcHOl99mCU4UL7rbvM2BmycFIVYTMDHwCONcU9hAGjBZQ5mErl6c1
V2ZafklZTRLJ0ynfsiknlI6DTlyV+M1Aq8lBMyH7LIcw7C5lc2HMTK+yTzpAzxLc
BrAv1HTfZQEAD6ViW31nDtTPgSiSK8rtvE8xvtNgAIq3f9O7ysMqNfz6J9vXQ/P9
178o+73aQcKvURGdv+6nkZenZCeIlGVHpoEdXFnGTZqCTnGTGcINXoihPySfr/8c
gIV3/OTD8Lh4Mh+wjzMcav2v2ppn4iwfeKokB5yqmcnyycW9i0OLuC0YnrcqxQVI
enNgWE2s7cZ767bEkbvVWoePLDtJZtdDe1fKMklIPqRBblhaBFfG2eYb6iJzLMKR
uLSPJFMw9j6itFHAI8pEzWE2DvtZ7wxz32I13sTgS7Fj1aEgRlsdbzzrs9dJk+4A
GefABJe87SxapUT6oxsgzUwxZcG6lkxvewjM6JjZx32R69WmnpCkoiTDC4q85Cfc
Bv3QMU9C1jRiWUmZtnTdcNXKRPti4wqvVEBkRjtdJX4RLMI9dW7UdFYISfqJda0L
wHtAaixcBVdTpY4RHwiZ+mGr+99bAXsduntj2AQ6v4yVH1ykHEfgCORovAJtGfny
ZWyGt7adhxuPdPJqF+NBkjT660r/LUYGYUV1IPAwd9zg73quVT4SEHGG3IypyGXA
2Fq10I+WWnGTFN+Aa6SADAzZgalCoMVCcG/+CmCc5LdEM6//KosIgcmBQVbKdNnV
KSIEm5Me6KBP+AL63GNms3j1nA3Z6P3nw0tz5Iou38WWEsYvcn6BknuHxUP8/jm5
xVzdmtf4CQcZDXJq41l3xmc+U565nur1x0z6zRkbBFjYdk+DL9rIA6dqXSnuCdu2
bioJCOjacXBWkdlV4zAW6HuvULb43U6IGf5pmKdb0gtxMVpLD0ibFyZqF7pHp3Nx
fp3Xf+wC8zyaTG9vIyke3CNwkigmWNXuQ7bikDFPAaI0wCkvxw2oiMvfzNEya04Q
xaT6WtWz0T31JbJALNHOGwghot6Z34LMaKHlcs7pSULZh01KU4KetB5ay9PqU77i
82RljG2lgC3dBSrbZsxLagXxBOlHAn3c0ukyEWq0mZOxdBSKp2OCeKjlThaK7e8y
et3XSh5QqeU7hNJPEWNis96UutiSrLMNz45/hd3mJ4UyfwDrC/H1AK1Un2jY3eak
8FYAUIM0UlZqYWyGmtLYJmDNZXYaozodICoUQlEMZyJhef2w8M5/wDvDgM+RLHhs
u9J7XoY0ypxEH4vsirQzV3WdMZL88BiLg6yFJcSzEEKez6ytYm+J4slWwtnzSDkd
nHDh1e9ZOpnD+bunCBLqz+LMUUHkky+j3LF/EXI840bZoMMo6gbelW2EvK2bn2NL
j2z3iYPAY6wD5oWNKZHsyQe2DpwcOidh/uadJHHBM9tJTnVwtTI0zaS9tDhkupou
u2Y4x39/UT9Yfd7kT+urqCbLXcIigdnAzOonaSilArB16VKGub6NOGqwnrS2s5dz
AnuStKBtbpA9uEODSrrT97nRQaS9F2//w5Slz3XjmY6OiG3jQK0O5AcDg6ZYzk8E
+bllOF/7rFUfjGZnCvjYImAmhkgpQwPugVtXYhfYsaAcrD5Vzr0afBDR10F+62pj
UIAI/sUaaAsd68v1GlN2O/MW+AqltLXOWzRCohVs9aFUX0U6kNE9w6zQWDKxIh4b
eKSW2Z40w9xgwdnIp8bxT2Ho+XT58OcZvT/GpS+l7zB+eyB4H/zdkKfOnmhvTua2
XIdSkwFLs2XWFt7vHvJcROokYSPxkII3wZUlh6OddCyJBvCwQB970mG01hQ/5cUI
rD1zGR8H2TbikSPPfL8ILbrfT6d3p3Bwt5tADKJEvRG1s/q9bt7Q9OaUucWQaF4Y
rdJmJqpy830b2BoxyE7+uAeHNuuu0OtynFMUZQMrQgPDL1yZNXUetPWnexdjxiXX
4UGWmLW8VQhRgyo/CTi13R4u3rnyf3Xf/pl9SmCKpyWjUO+2XLoLiwpWyKBj5tYx
dFmdSXx9VbrUF/JkBTXQBbkT0szHIgAFNAo2lDFBEaLwTriJ1MGkzJeR4tAZych0
xQGV4yIc4YRJ5Vg3C0Gf5fXoVdbcjIcmdW1zDabvEu/MsWxD9hvuHSufg92cxB5g
+EyW59PNlYmsd8LtwvoVVlnpGUVqugMFQ7GUtLWvDDSG4tdgchnnDTtyq4Hj6SUQ
MgtJaCnuzeTkqdVvVApMLFR33i4QYX8aU1kCTbngZD0JXZuL3KJ4YKQG0P5psieR
e1/qvEqhYF2Jvng0J6+lqwjdkuVP9mR3WqXwhW0lwWQf0rWx/dsek5u1mlJn8Kez
DbUrp2zJGHz9fwK1MPQnNA+4D1GHLHHpZ30PDyTjR+omVrPwKEp8S/1QoZWEVQ0n
xyenNCvbaxNyg/cgszL3ghiIR5ZFK24hrdBdtGvbYdUkVsI98VZZ2DL1OQ8IdE8V
548cGsznfJt/+1JllX3Cz4EeScr52ui5fvk632LPZZqigCGNE+C+F2z/7iHFlWvY
4LvMQr4lAkmbovaoVzqXUoGyzhEqVWeqxijHXhPf4nmQQ7BP9EpESYA6P7aB8e2g
BJlO4qOXDkjjrjYenjarHSq40GJ3PeQwa14UuF1H3HSoEsX8mjdQx2Z8JGYxupfI
0y1rqsFMvx/T955V6E9Pi/ZeaG+SmOW5RrA20M4kFEIyx67YNSNL7eB3uCsoTTWe
Fu3mdezaEJFO1KgeLPiT9Vch/9dwUOjEjnjDe8glIbJOE849HdPkUqHJ+IFdqFZA
8C++UobW+Vkm6zUnFaOtkn9v1HxLyguyzwQUiMvVbavFNm55gkTJWmGsfPzu2h5a
g7S1kFins9GGvuFVtWCfxc/FTC33S6rVYrZmHwqVB8rocv4+NpsJTg9H6xEK3iH6
EIRggUFGOGgb8Ey1mZjcu0QfqyozV7dBA4W4Y00c498oiVrnThrp03GngPMPLJx2
ZmJpv5Hgtch8K/tFNZ9OXYbN37JqyGmZCT7qI9E+rhfLXlBJwiYiL2eeBULqx2aF
YgTRxNomeyeThS0BMXqhg1fL906jaqKUd+RZvNNcnYD9Mz2PCeX6DBOVRVcQv2jl
9cNhzH16dLqhQ2tgSa3zHEmiymNc3Hp+1YtRgAgtWkw2VHu2v/OsuPjV6xh1rzIG
zHTRejhNslRWP0ZTX25OiQMeI5JqO+LFRUgSl1NsmAQ4qGa7s3fmGFo4NFtLj3iz
XZmX0XCc0GVbK2+1EmifouSH6jgBUECLddBNOX7+BcYKqDLktcjtkSq1qO5EjGbe
lFiU6LYf6amCXOCpTyQ9XY+vfa15qtPbHpI9vy4qfe6LwdxiZdCzoBmPA+g4zxqa
NpvrVysn47Rh4EC8cjpVZ6vzcEPm/5q886EQE1cTlgacmIOL2OnNU1EAldcWkz/S
XrlUf3SZkq8epNlVaueRBLC91biTkhlMF0KyAsVE+4CW2tB0KPMzHFPRY1WwaDUF
K+yvCz9JSzW1NX03UwRRp4sfBe6Cq4906fbbGigY7nnqCoRRN2G9vnUku19b7vQw
vGWqjA9NQRSBQD2BCmYfNveptNDjdJgpwMWjtAsa2BbdK6Rh0jDsbXSgq4SSihrM
5tpRtIiNerj6F7lKk8eZg+N68IZBa+V70oW/jvotx0FMlwQsFNsDNCQUK90pNHMB
qKdyiFpco744p1QFQfOsVatoXZXUQAH10WoD9UGc3bwdAPsX+DNtN2iTJEY+FJQ+
+0JsWZGYtc7tZm9YuOvA5D2LgQQtrX7Q7UhEIKPxUaAUfYZus56JrUzVvBXn7z/v
221XOM2b0UAbAQIDcJTg1u7sohK0bJq1ix36UxdS2d972xFXeZJvRPXI+ceH1cdT
xVWdXelC89XftvCcAoK99Hy6xCfIULBTkWcxDSn3hMWLOaGr91Jk8sysmNtldDA+
JkIBET1kMd/HAgt0ydZc0hf4kvDavGSUYvBkBFqzu+UD9/hVqmM1vVc17U+rnUMI
dNHKQY3ilQ1zfDJ5Rcuqi6ssx5jVpQJJcM0RxQXyWJ2/D+quHb3bdKSGPzLaplqn
W7D1REQF6HV0Xw0HGOQkyEcogFYBPfzeazaula5TV741bnvfHAmqdkvr4igZ+P65
qKph2IHXs7YGgsknQGduLMmNCJkI+GHLa+Sy48USmT7uDUFsGPkOhFYdTUCpzFB2
V75IO99Pp7l791HOc5ql1lTvP7ZT17gLN9bKICUM/O29rP1V1xjWKl37JqQc5V/6
zOCowAjfvSCqGGJLCiDLC6E2XuHaRWBYJlN4W4LpWS5MbOruIcDlNHYw2VvKP/sM
kSIkWp7GxYFVsHOgt0RVTeAXP4UzEPAG4aakPCv6LQgXqzWvTv5tj3chvXJOXyYO
HWo9uW6Sao7DKjQztNUrxX8u8/kmXA8X4alNO98ZNbLnwksi41Zhd4uRVxwibfSE
68iOOQvR6WRr0KAsiUlSOukJ7yV3W0pDLdVIDIWt4GY6RNDRlv/rDHhDr1HS67ej
muLMlwkAxC9JbU5MiNRwSpJIHSgrdYSbHdeLs5ZXjBObCNyYlFKfxC34bezkQXhv
fGXxQKORE+A6isUfpW+0/RdMxChydPfN1vRbRE+iz9biH8klT+8Vm9JBIg2she8W
bGaTbSsaW1vCIiPmTJBeeXyNvOfK+9x0nWTkX/MBIDlFNsB29cD5e3idGWa/47e/
Q/bRetxC+q9qXCbDlo1wQEzvYIuUnkMJskKXMZa0Mtzi/IxFofTeDahFo7Gn3tLO
KCx9oXK8u+jim4Q4I/LXc4wsIkNpw23trX0S4Y5npA/aZ6K+1HxIALjePn6/UqXJ
xvy1RcncLyFp0uUPC558HPxu04tUYbS5zIwMS9WTeI+sK6zwU8xkfrnyMoSQPaZ7
KsgRFMxjQj/fgcSgYEAa4QsO1EsKbA9ePyFNCF16ZarMYr9fof5YZ/W+7SZzX3bt
u4f34YVHgnTAirucQjrU81RK9KyrWXFWq9jtQCEbrCNYYbs1XCTQKjrPG91baRDp
tsqT9x7+X32a8z/t9KjXE+bEAohgOeesJ+ZZCLyZk/HXYFqxgyKzUaqaYXuSFBjY
/3rnbMTt3MwSYeK72CkrGi8+nfPM63DixaH1VA4DMjQJ/PibfK+LcRvZ8s3q9m8S
o7x492JUgb/miu+CCYgT/pCOKEofkM6Lw+5KiHxG+2jPRFConimMDE4F9U6nHATZ
r+bNiC8LPyYSOY1vYeiPDjc+jtroO79rr6pu4ApMZXk8Q5MpjtnMH9brawpsq42D
NYsTTY+Ryjlfb7G0q7J7useLn7fGXeWW97txF/meXfkztX168UUQEdNKSQaGYibr
Ey7GR0MKgcN2kDbzgsmXzOksj8aM0rTt0zW5CahVGwXgHJX91p7Ami9ZXqmSwMkY
7zfut/LIEX8Vlwy5kM567kR95I5nLJWBYZligwkzqz0RsEwSL3Yg6kNdYqEIEs7M
PzZAEnzCwwZT5LE6MoRLzCsGkK/YXw6D23lP9xHIakQYYfTG/V7z9xOAh8FAbqc5
+OwYno03Ry6sYL8UlSbECJ5VGHTV7n/tCsG9GHA12HrTXWcoiz8ZzVLGICdRkkwJ
LY2NksGfgP6DaEtUzcZaWsrAIccDO+8u1uUel580t6n8HPZa+Of93BWIuOjpwDJH
7u+gVOCatm27Nj7/vga0nQAWR8RVopiEE11awZB9JL98zU4MZb+Ye7CWms3MN8Xt
EEYkpazbeVXSofxp8Xz+yJW9GNMbwSs/xXDevx54O1IotXbP8jLp1vW4Us7+Co/p
9DWuA9vcw/HBtFCeL9tgWAbT7ZDxQgB4WBLlW/SCC31pRSU7vi40ccOOR2blzM0A
BEy2eoFtsOz/FC8aNk7cv5mq8ojkij00ToILCOz756xQioqC04Kd6tXRiqCkHKg+
kU0on1MOvzUctwXuz+DqX0/rQ80ESgQNq6tYDHZimQA2DkD/K5VeljbGH5IHB/fS
YlXPOMbYwPYaJh/YjQewejvg0CVSlwMBNKprQrfnURmcBicsfFuo3UudXrDz589n
ZKUY2kYKgHpv+tlkixesGMr4AX0YPHd3HOvDch1DKYwnQYGg8oiINS61RK6OGAOn
PazLDqX9VAs+QKhHb2rHaAc3Em33ijI/9TqxVqeUWZRaMfDc38E2Q2hXEagZ3koV
b9plNTDhetOPHASFYpUPiU6c3DXlrquDe4kzshCnG6klQtXy/bVTxJ9BMxQICgqh
jTJxbscB7O6SvUZrOLm0MMODOIMvhuLGyWQjgNr36EAhRgQv8U/+QhKbA/1j+9vX
70j9GASIXs8IwC7yFhAsXDKc2zwt8qJ3fp+bn6te+7rDwImQOmcnuiYQuq7aF0Nq
xM54YEYoc9Vh0ausGDexzVk9s1Yh7SNHTuTzGkdVaIbZtnTBiackjKjBLUxSfTC3
l4P8dXxeeE4QMh2Z7JS/rqJv/6guHoTNqnwmgV1msRlMhn3c6zwUzqzYcxiixQc9
myAavN8enZzIMMyq4ea9hAKOF4eeIfR1sS3+h60tJObTmr0U6SFXVYLdsWyvaw+S
UcMNWcb8tp1IKW1DtrumjrvzRiTP2BOynLVX68Cz5WTpwe1Q8+0qKYZoYYd38jER
3A8yxGqYVEizk/u+JYLnBOCGFTKbWxUIoQ238uLvH2EzullY6NTHlsg1f/LEWpWx
AmjGIUyynQ1U2nvwGVMOCsNon73y1hGpIfWGY4j1XOmltxjrNzvQvmG001wyeFmq
sUixdEjxe4MLOmYmCNQBLc9V/h3auuDJyXquBZ6yT+CUueRZZ/YSMMNxvAhbrpjw
38r/vYw1PbmgaOnGxBczv7WIAxA4ekuXxksfrC7pVjWRHtZyJartfxvY/edmQYki
2oCc0OjUGuaiSwsQs+JODyNGGaU8klCMLMDHw9seBWJ8XSKRkBiw3oxDKnicIEhj
Foc7mvd+31+y212TbPaYnWie6e/CnbLJqLCDtZ3uL4W3c0qJlALY49topPzOQ4/m
FT+l8E3ia6VaKnGb40Kz5uH7J1djBrkEX6WlfG5fc3iCXE+jT+OcIkc/kr2avFIg
g+iSL1o8X3+D+0qx16nV0rssNW/h/iFyevOlUyvdxZaiwUTQYqoUfG1tuh3DT5IT
N29M3Zz1RE80oPKnuFrbzm8SLUeAhS6rkDo3vA2N8yT+vG+jBbQ4fn9p8Yfv85Tq
wRyWDOdHAxUdeIhfYII8dlofABkyPb6hawzLQqZ8UKnP9tlSUMZgZmnl9oSkvrd8
7Hv486dt89SYLDdGbl4EacaE72E+zdST0czRH9mLM0Jef/v105CDXOM3eI1rqFEk
XNeAmLgdV048awW5gnVPBwffU1OxSLCBlOYyzrm7ZLA/bAON+tq0R9jEP3LWU5/h
zJmjyVR01ExSUIdxq5Ml7PbjMYA1M3bf4ETuP0oTZXePcfyMcTVzUDZ9S+9O/Wk9
76bIzscF0QUW2nG0qcN6v29gTLkeK32R4gnpFZ/pBHJ2/DfXabtKvimexKWR2PEv
xlIf0OtxGssBG83F1cfxBZzPKnD23jsoXl77KC8ljr6qk9GfblSey/y2ZozUcIAv
bpKKM2c3GCzYNTs+O6uxYa1ZKO9PXBs+OsQDzLT1IiUfropwb9M8LPSf8Vjd7xwb
LTizdnjZdX9GZ4UkYy5Oowvq+vBV1N5IPfmjlI77ppagXwG5WPB/YsRoC3d1GX9+
kgDMSOREZ0hIlc53X8/TQSNFaoD1DBOq7w+7AlfqxXSD9IcFTWOmWUo1ATt47XHD
9qnm/x7zM+r4w7MsmbAZYURrDE6DFLKWSRuDGVlw2yOyeW95R0h6UbcUJkyfc61/
t4zGgzwnLUSJU4mDDOjQ7WoDfSTNq4fauF1hdI+66a2IsTWBolFQwFs5aU+MYFDD
5yXYII+yYU/nJe9sNvs6am399YV/1i9Le0639gAqVWI/GWipsmlpBeF0t7EvZ8RA
wVEoMoURs4yyJ68aKmmUg5l8RlWtC56lP1OAs3u2vbg4AdF4OgD4QsMS5A9ZzEwv
Nhfw7vho2WVYah2UdqNRB1FMKVs+ElpzIsaTpjfTLn+rDVzd8rsIdfdG+OBdSmi+
e0U3KY7hC9yy8OWivei9Fb4ijXs9XlKgTSHH7Uja96zapU9SzgdBnr9aeXRIzyzk
vNggSJEAz7P6Chf30dAYVzieN2FiQCJMoQ9k/LGGTLhDipjOBiuFqnRT8PrphmIZ
gwQ+YAHiNfCuVJiyniGPJ/24V3TjLIT8ZP3lQo8rLPUQ5wJFmBYJrFEa0cdksxwb
Mwvjln+iRb7Z3g+PzXdJNOOLb8HBg0F7w813Sl6gpPdWj6+CCha5wcwbxIpiY05x
R76iRnu6bouIAyCOteQvVkQLQDy1XTA7uWB/00FmQ5OCb3Wrd/9PkOp58jm5zzIQ
17fXwLTop8eTNyHxl0vIUdcxxMNsIee9zvPYTQzyawBzw3v/b8eAahnxhlVChc5s
xk6/UsvtRmPEcOE6NbwcHs+yYoNXdOvnLy/oiV+U4hW5xXmMqG1GQdBiXVHrd+kY
KD3yJLVniT/B4U0i8F6Zt0V45fdTPE7ZRwyb+kPj8To7U9zDzRXdXIiz/SrZR1t2
W0d1CRc3HoVTOs1P8uIEwb2uBUnQad8jUjM4RhEgaXW4Yj8Y6wkOpulTEpsei8Qf
HFUcAWSeGjso71wXTutxF7+9tZhmIi34yWjrOfDxXmzNnvKRsXCCIlo1si+DJjmn
va3C8ZIJJW+ZAmh5e4Em8YBJ5NtJeALj7H4q1QIboHRZW5lhMseoedFzU5idfSdF
HJlSZgYSJvErclEU5ul4DOf5usWaVRritfvHfiOKS6yzHvCZ+fmwzefRSM3qQ0I+
3uMtboLA9LMuh4sroxfjl49AR1FysyGd3d54t7xFL4YkOXIqJuZWhCMZ4/vgJJQp
8rLjVOnTmEsTT12Prduec2/p5rJD0yR88WDECQo0bsveXwfUujlMHgtIGU6AWe26
yo8TTJ3CHz/ykrOzxhcRUDGSvExQPywlUWay6xkCTCUqAuCc2JV7tJdxMOPRMVJm
OYJSnAP8Ui2ayTFjnMcQ+bbbkUOn7OhU+eOhO8J6Lrkybc6V1E7qn81e3wqCEChk
Dndfg1OprYhCgV71xgKDaOV+RxWaL4u4huvlwgteIIQ6wCNnoawVMmuRzEmYQouA
lPCAs6kSRuYOs1InzFh4ROoRQxPYM0+BT2ZFp2IufuNIQ8cRJUmUTi65dBAX9z1t
WFIEs/ml3cHJJPUVrUC9Pbvi+D76Rm8lwfXjt0z+yGC+wnR5N0Q4OgwQ1JQH2HiT
Y2yJHY9tOVuwY+wYGpO6PeI1sWZzO4N5jq9YxeslQ9xAZSk9HrXHKFvgt5Ew/Eu2
X0by3eMt+yhh9Hz6FaXzxul17TtzWFyA6BUsHHFR6Xo3zasa8RCBLN11zNtx8T4J
xQqUvyB5eD6OFWujBX+ZTp5z7FCAOTaobXyJ5n1b2e7t7WyPmek2CUiSvb+kQarx
HsHdYj2ZP0ZE6OZ/U1D8z3MdYuqHRwdiG8eXayWc0/f7xWeHGscNyCmKGCDOL10i
GZFylDE1fls7eX4rfJmsu4t5OGI+lhEeVQSm2cSJtE0sosY2SJ3THnBKAa0lrPYT
ozga6dN7VYq8JD77fXjSjvgmeOWKva129i+IrsvZsrctfuA6xiNZ1ci6TKfC2Yln
kltu4QtwRpJYrfJpSkBbkHDifO+5w9Xcy5U/ONHCvDh2cnYotMQIumvRxiQREoLg
f3DsOR5ZLcFg9gjlUN3KNtTiwlu1DMeoNKmPlC0nyquOwpXsEKgbzcSEO2AiD7DR
eOlC/nom7yP+kw1vnJhi4fFzAf7nt0ORLVm0cTrpb9koZhTV2MuaxKn6htXJmgVw
ZyxsbpzxlzuYSLMdRT7Xj+9kWmv7LdtZxHXlnrwWGZOszSOT8d8/8IDna6oGLJDI
Gu57EG0OJLGJsGnmWmToZzocN9TkF2HqGw8Iz8DqK8LPfE7EboRAoWdSvZjLTFN/
jSrnHbqio5j3APafxrH5A6fLExtZal4VToOVdbHeEuBoOHxnuVIqB3npSHr1igaj
FcaIPiF2WZswOLUF/AhwjVGL3DqIfdapyYVuY/tykxt34zk7GGSb8zOqpv9rflNM
s1Lx5ZSg2OLO681K9DVnN4GXl/1xtqd3jAekBVBosV9sgUhBSQ9ZBXthqs02YulN
UEYk5Yf8DA907KG5Rm5aVXJ+Xb3zg/FsqV3GhyAzOY3hdzAytpUpBRqGYvkwgxhK
TPLEj5YsVmKjKF1pd0lZ1anaX8CyScFYJsFGXGGvOoOfiWOExcDZCZ0lDy+DkKp3
LyUj0iKp6aTwvFxVdOKbHkxNcDlOH4E2sFaclff44/SRmyoDaAugAXxoOT9d9jUV
FVnDGy7/eZG1nuelnqYzyWmj1gwjRyv2vJHVPvrGHQbGbtvPqNkveJWxwv9C5IXC
z6rZSuiLmzGi3niiTk0UnWxHlWzXQNXfONP2l8WguRZOwNUE+P+1crwFJr5pH90E
hLunKYIZUHZ2LXkn6tU0m3KruCCkHrFJyP9cC/42p8y0rzOd3ZdCXcCcZ3BAWKSJ
UG9o3WBMAr8qD7Q1TUzx8yNM1mnIRBWCYmxutKLveiAJPTQkWuVrM+LQ3+FANJUZ
ni1so061/hhPCco1TbELAeFVJSzgVv/OzLrTb/xsumnsbTW9wa7RT3vlIXEhfnFZ
H1xyU5T2QlaW4du+VNWCONeOTPaEXgPaLT4Xrtv00v4mfMFxkKRORxCu1+a3q7Ts
ZGm/k5LkKwUHKgD7ADH2hH30NcBKhruFUQVFiVHpmq3gSunwyaC8/AVYH5eSzgnf
ZRo8PLxUsi8Q6FSCykOCbdsr6w2HeCgSlf0T6y0Xd1jq8E1UeqrfyfKmqY0D9IlH
+BxdNLUjueb/IprDan5iMdTGdY6tCCO/GmoMBjZIJA/wR5CBxEBD/FL2lWpQ5eFM
OxTv8BYAlfmVW55rTbwsvBmMqk0GL8Inm2uG9nBKXo56t3sr9cLY/BI9UXnmJoQe
VKsi8utmkjrC9LYg8DsN9w0BH0cUwY/gevSSHzAiPnCsaJX/fkGux6n3It+aTPvb
L8AbOGNQwyyvs9+82aGv7YzcHWDGfRPdvZGSQ5FI5ZRbFiqeWsg4EWvS8SWcqTa4
EHE/kk2S9CrTp7Sdypme3o6akXNqavif7bR3bdnXJqi7rilyebksS6ySWvmX0jT3
fEH0ekyZ5oLShSd3qh5S2RgquxZlFeRoHam456syTMLt/BTrPjVJRQyaNu+yh0AF
VMOcFk/bIEcg775S7vo9WNONUWbfpJUl77cJZLuRqzbJgJL7OYvSLsCuD0pEXZKe
unNOC4KbGe2HQptyka3F//15itu0SBRJkmlM6yNd7G+U4PYWyyoZQ5Jcw0YG3vyt
ysdTeUPmbMYfC/SVxVGmaGYpy9Erb/bnv+nIkZgc9rbCAXWwC2tC2coSsnGLPPvZ
zr20pg5GIFI08Wolt/LHyuqFU4w5Jjw5M9oTQirVLzH+X80q9dx3nWTwSbI50hfX
VXQsWF9n9GzIipwJ7AvIV3NoikZ/Gjn9gMHPv6Y7FzQUkq5BY4b49N0ByoayQtVW
gv6zTh8dptJyT/oy/NJoODRBcokPqeFYsmSaaP9eq1id+sO3N3pBj9EkVTRvLsQi
rNk+72x9lIXY4RHcaEf9MVHmzaTeCrT0/+t8ddi6kYmZFoQ2tyIaYCoawSC6+66l
i6/2uvU8/GJvpWk3TqM8CpgNp7Tq7Whh1wM/qJYbBRfLscS17MepiyaC88qxxFMT
DNU11T6YEK/rkdtwAfJQVnBzwy0KZDN7FGoWJ4UbBsZgDQM8FZ2othJN61XcQvsB
U/bnomojaWwhSf03p/I79vEnvkdZkFUAKEUzmyNYsLjtixEXlOsmL5wr6zc4kjqS
iWuT+kHwJ41Kg2ai0xQSGQgfOOWnVYmIB3lMKC/w1m4xqAmi+4DlsQB5eZUjHCRE
NF9oFX5N8tcInSpqLQeuaNyudUd4CoWSbktwsNg3sbEyFqyR/urUAv8k37qJoIqG
a83dFRpxiPPt9MNCx8VctMIlQtTy7wEDO37b/Sifh1LkkKmGnyiPfFAe4av5w49E
soY1681wsA2s5Fs+vaupIqMxmhikodpaZTLYsab10qrZ5JHIVw6Cxy0Yg6jnTOKC
e+HFciMD9MCoGz4RA0B14357SPJIYmh9/TI07fnGV/2GUQ6mpvNQYVX9JHFp/BfU
eBhZz+nrYiwO6d/VCoXnQaeQXg08PcKne+i2/GeV8MGjUkvUpfmSdsUpee+ePDgq
JUkywuEbSG2pOKSiLuP8sXh+5RPflxVtJWZc1ja9t9NZ7S12qFnos8cNAXzvAUig
eSlzBMUoZzFy4No+ZBMGQTvc3Yo1g12YwtOQiALjpsddR+IC6AY8yin4AS130kne
E41fZ/MmFIrjQuwFQDiRwYoETOY4Q2KmAroHER7CqIsXt0mOg5BuLMsptGmRln7r
If/4niykb53/DbrajhIGK6tlumjQ9fcF2tD8kNID4tyZGMk0p1c88J5y+JXammkm
CRIzXmmxXWRLuQPufXsZ4L87Y8lDD7+6to7zVi5GKCR836/d33J3oQa8GLxWsKb6
1g577L6JRxSrvl4kOX01GLJLMi3knjUQkLSxAGCawosVWbHJVecwcUM5EPMJtpIT
+5NpyAOeK6WZNn/5G8eyI+4PfmbYG+dL13rQ8QgiH1P9wInAAb7PFpcdxb2jVupp
to+sziId/ATKxfIdMCG5hbO79CgtaMaylO/uI6I30nwaNuP/cVTTzkZpnW+krGf5
hxRhRt79fHGXhpGReIuHRnzLdWmeELyTPZ3Uv21sHLcwDylHJbhYwZWtG4VsCw/F
L3VA5YG4K7kXWDsXidnJDKDBXD9I+xay/pUxNGj7RRp6IUKmRWnKxjsCZKD5Ztac
HMKzYxo8OlEyZx9b75zSDq7k12+ALWZNaT6OuKboUhUJURcrtsXyfVc/VFPbtTTq
zHqAAMZ0I2zzvKUjzrmG7p7i3huxy23JTHmggNgbai7HCQaH/MJLO2YcQiNsjy3y
0wijnQYrWMncMH/sPkMH34cQSTi7npdzVIqQOnuTNzEe3BpTijnDUA6gZMRb22d7
+yoBa2u33uu/0JtBQcSSRovHHSggvuJuAargWV2pJML0DRx8bZ0aisR5kTj0YV24
wDHQ+hazaYKWevvejUBoE+wcZC6ZzUfMpkSG9ydWjqfvGWPz2IZCL4VtObg95qWA
2hrKnWO3LPsArCrHZ9J97YmK3YANT7O2Z/s87zh7iFrJ/OE/gmCI+Jkx38qVmnws
2mJV9R08JSm33E8HSLBNfUgA3SN4MCaP5zY7x7xZ12cbok/MQzuSJaWywOu/4ox+
jf3QGvr8YRhFMZ0Xdt8diigALhm6WFhx1PASe2KYZY9nJizK8l78Rhvru2E7L4zK
L/4AhLI07m7LGz5msjdbI6U252FjJ8APAkM4hspFEj4as8DJneKXFbEcMT0N8uH6
06IrY4h7YOirHOTEfApr6SpBAUwBwG6JyXpRTYYrCUWmZIvsXu2RSPSoiuKiwCNN
mLxdd4M5cMa1SrgBtZHhsa+w/12AfAVqYHEDVYZHTNyTdMyboARFsgcPWT9gvbb8
NZYyCNbSlYr1yKpmCLjt7VoqvMOk4sNIxpkvxoAvlnwn2wl45oFc6FJphkWoSU6n
gp75+tu4BaIym8aPf9Sy+yIL0MSWX/+LBi/XVT5X9RgtPhmJo0PYzosj9TLV4Uh4
Rjlmzhevjdy3r2DVWg2/mjNdsyrK7EhkOrvB5aEnl00eMtgX/NZsF9dkrSgV/P/v
BId52fWaXhvjn/nrYoV2HZ8e/ETUtEngRk26/c3zi7qIQDbq4IjjzaQjdzYEXHTC
M5iUZwLBW+yfm3lf+g9yOCxjFHpMhBFBVsopE1iyxVVNEl/keA+7OgBCp4FvF67e
vDtTzh9lVW8VJ6EdFpRPI3USB9gKz57Clfg+DThZ6bkPeK75DR0kXjybCb9eOTMx
opQSKXJAbvdaIieWL+9etxgbfmtYJcidbIUD7oYZGioGUJBrKNgu/X7LXAxHx5y1
N7OaeTAzMY9swUjOUBX8niPLNiIcidOKBsUIhyp7nIrCjmG28eQsGPkyvjgb8bnC
ZEgq7fvbvNp3xtE+75zI2t+qcvZjNTzhArwrr6SJjqsaT2lzLMNky28mJk0++iDf
Lm+c1o5ceQtDaijuh1ZWunH72e0AYgzuy4aB3IFRUTmbQ9NeVKW3DD63bFHlG5Im
E3rmovDwm1m31WSrbVqGNK2P9OR3xn8Bo9vJ3AYIv2Xim1dePLNl6iL5p8dt1HO1
2v8TpgYRBSbbEXjwmeZCmsp8zVSqNoynNZlxwwaWxbpvwrq8JknsdJIDQrC3iyWC
ont09g1dE8MXc8nmh4yH8EfCUr3CJGywisIM82RJpR1vRvil/9q3dfB/Ka8xbK/m
RP2SbrjkYKiWaz6k3IibG/ZaSddfNNbnyYTCA1JJCZYPTncv7SKDK4bQ2umFiATn
8vqSviZH71oL++7BEliB6fdhU37D2uY9LuX309F7BhNJ2vp/zRHph20Vnvr3UVNz
pQ497nmjOOzt18u0JAtB9yTA0+EgpchLzqtcxTytkB1aTrVGWxaoQGK9GtRvjOOt
SHPtBOEImG25QXvECeHvB1uALi7A9ukCjeKrYF+3gyjqV4mxq80o/If0OiXxGiCL
vUnIW0T6j9EraGx2H+Ns/OM9t1l56J3xVP8wWzUy8ie+2lP8bTqjI4NYsVRCIXJA
Ra+r0DWI4aHvi6sEBGfK/Ls7hQGXZsS2dpVaapkvHvnfG4xMtmQyJQQc+DdCtQHK
ZP542W5BNyGFvS1G7UQmj9IDzfrD1mm54rKuBPB2fAYOWneBehIbgku9NclAZgb3
7h1sylp2FIIjSfY5mgWahX+d46kqqSaN8AfVaShkA0C8cc7AX3dQUZ/fkF6hXb5j
+rQjpFRFzgk3Ijs+yt9znP8V/yXHhhm0BcXwZbkrs08XZM7FpO5t2cTG0+wE88yT
AkkSyCfxjUpek8ZobHcFWoZs8yUtSHOs9Wwbn/prxpGD3ytAuFDHWcmzdEY9GRJu
nA/N9xzjN7GyYyvtW2PaAlqrP3fjU2OFcFmvZg8B9syHGCwXlRBsx/aB0fZU2DjX
zMdHX0/iX9VUEyIfcQ9gn5cLfCJFb1mdLAiO6O2KCk+4k8xD0JqX/hyrAhPpZM8k
XpL92QNlfBHm3QSJxLqnLEVjX3/0gJjxV7MZjc1bGWXliYd7baJN5QqmLWNLuA/v
jOdq3HiHfFbqE/wh5a+uuNrxWq+XOSjUGaYdMw7kd86AN/iS3+PlixYEXkuaT/up
5HLQScHFwcwTCgl0QRbNgDdE1qZpw6Qzz1oshGyJ9C6h2WhIcPJNInCiaKYjoYRg
AWM0Nh7wDpcj8mZpBfA//7pWH5Y9LlLb4zFYL3YUjGZZVFI+/hr6IybeHIkRW8Tf
Npqcr9cy84VvodE8Ix48y43pucczU+b4G114/F+HJcl8LzUXcVcQe5D0/M8ZPTos
Io2aZ1n1EQHuIY14+PquskW3E3QZpby0SQDAP6tsFIR62MGMVn0JNWe6EL2RESIV
indqAMrmXLqthQiCjkwHANPTcsWgmIx8qeEQFTc62j/gAsXLEeaUf0LPAlf5OuuV
q5FVu8muz8FZmTNEkmMroKSaUYuCeGh5JUgugUuFGQ9iqBs8nrApLQydaaUY7sBI
09CJC9AMqopjbKoQD0wmjVTeXawEtl+EYB5THYgIatn22lai5wNS4VOgHPLI80rx
dlM/BeAqME/ilO7gbMis33ywbwFaNbF3ASgn1smFSwUL2G4EqZH2MS1qgjOD0UMr
mDSzr1gZm1eKdMeNKqLENIwqU5+B+7Q8mLqEKZTwIZvQ3t7mY0TR8Ne3x5FEVNF2
yrTgpiIvPoynIIIvbJnC/4kI2NPVuL6xZKcRhl5YCKY4bsI22aatip5eyfZxYKAL
lLBamc01aFyGjRQwzxTvml0HBmbjNache/aUB6nLer9619Rx4dBeT1dDe8pD+plv
A3wd01FsyQWbw8NRIDi01X9QS2dKjwPjv7deJp5sJhV5q6MtWdqpb94XuwcO7F+i
g0sv4xObXXMiQkXIZ+hagRLmMhWidpAS5VUf/tyezzsuN2IQSJkvgN2+dSVNe29E
Mr5SkExa8TmzxmB9wkcTDDNEIEdgr0TU3Koj0Xc4JLoi5vWUIare+lQyfNJcVSBX
+C16vaOgKkmzg1/R+iQ9vvDQnLu85aAdjELR76ZTwMsieDRgfZXSf1V5AwqDz6gc
vZjVB9dyIyWwquivhH3girTiY31equxMaTWGSBPX2fYNrdfJP5PflysNSzn5rFI8
t6ff3ikb1Wr2J8/eR1zZNvEkzNFJu1jN+3dih9f+JzP2j+gCM5YegNER9UhVB115
QpBiaPWbK1lR1vcBmh8VXdvnkGM7zfTMn3nyGQw5uF1ppA/Oo2Fi9DpdByDjR/WQ
KFXKhkgf16ZL0HdVTK8ZWfAE7uI8MPwEYkonsOZPLGnf2iiY59J6fBnmKi3X3SNB
73PeTwBS7+3W113jWasNczppG1QHhra/VQZZN7c+aAa5XEBcpPLeE7YCUZfN6geb
S6AEbZB10llWMNAVYT2C/edIeZXtiHs+AxD8xoivayqXr3AfxoeBPWlPodIb+QP4
ngen4Ut4R/Sp/jdkSAd00M25DQgP1EmywF2qhZ9E9Smp7oeJLe7euv5qeWZ8kBQT
n5Ca4LWBhx3Y+TQW6fZWsIszi6rUjApegDM6c4bMoOGp3+dF9nDhDgdFygeGAXuF
p9U++D0IGJ2XDF802irc41nlUhCb2xIFjC+j/10ofcnHg2IHYk3cBia0OyS9NGC2
68MDs3oMvTCTRmqX3ZnfiA1gSEB03u4lRkH3aX9U4JopgBuaJNsakU4HbVlWcpU/
kCM8gT53k9/jQNTvww2psvGGwu74x05R/Q6ThIoM3dT37v7hv/OUD3/Z31AOsXEK
KXl3VV9psd0wl5XICxhTb16SE/tSMa9rArd95Z+jyHewsowA0Ttt3Ls9ipfxKGHK
oNwIUD8YP4zqZNZ9gYFjDPxcg6gha/PisDRoqxyf/BSscwBYp3ob0oFaDLxHDp8c
W0l/dtmuaNY3/s66BEpi0CpVIu+oa0WtdDp5xOsxjlUXbMv0mew+S+VGkceSKH9K
Sohqlj/UfLYHunLUwriLCTGmMXRSVp/MAnL3iQlAcwHtqtlldhFP7xOnOEf8eDM7
0luzNn2s0GMXDpzYizS3JY4VpBgn/vtkI8DlWylpWZ4lyIMFiphbIH3A5tq2Re9N
SnY1kdNO+0l260EKEkhbAdkgV6kTnvq11xGQChXOq4gqIhK/PQfC6ergb3C7gTlB
hhoykmyNbhMYnu6IF2Y4hKzG0thsoJTOiMPsBLQzVATMtsLkAhSf/WXCfBjY571n
xQz5MaxU3oaGS6SKWcs8EXrAU6L3IaUuscWyuTSB/36O6zQQMnTMEQUK7/20beup
7oXj/d0dAa6Crhp4y1slcMQGxkk4qMbIkd+5g8HVUtOlXIBCdMLALB1tcUmMHam9
5+ti3M8Biu4lXzcWtiT6JeiY0L8rXzNuO34m9aP3k02zUG3KuBlMNtau8VWDd2JU
RzP0ibShJxJNii/CeySY9DBZq73MYNGW/NFx13dAxpbjQ1v75i/i5VJAilg3NpHz
5Tw1Xc97opj/llemdMnJy7JsEOA4Aky/yFjK0cYO+LpTaiV/GSB088hS24CJTv43
2i35PQFw+dpAHpEYG86wMshMC6P1/i4k+mrY2qRzIltNsxekOz1REBWtcVJlbr9X
D6U/6OlKTnH/XH/QJDEmetQ8EEVuvhu0q+9eqd50Fa5qt8p9azdL1jGo/vc8zR90
LeQfQFIybLqLU7dvLcaPIATdtmzfKLf8Re79pgDe3V2Ho6P0isDhgcpsrSAyeld/
QqmUI6UloDokccM2cBU2l9/Rz2ovwXcBCR2hSBObaHjGEhrkfaDIBjYZ8JgfKmXh
tEsyEUP11JHl0/lrabKEIyC6vbP8fefKjldlaiB4Enn5xzKjGDWeRgkxKd7FeeTk
ze0ypsh6TC8Fa+1mGSHgaWjet2PomUMAKngh0fKNJSGKuAuSHPQIp/5TwbhhXBSH
PakCJGaOouISrFZ/mVc5xE/SuRbq5JVv/0APW+0R4Ecls2BS7lnKYTeSCuutbBzL
v2zYdEWfJywQDH4ICAvaX5sWKwyKJ1LigOEySgRVP0sNMJA3Be6G+E6V6XHwveE9
GpGlHIveGWAIG6+JrWAb2qTF/uZrZvYnMyNMNHLnmt/JPbrLpb833RF2qeUKG8Wx
/Mp4LFoBRwnentrrAdmwMSjl9OPdEVrpd+9fDWfv0VReG5zcxYbQDzUCgij0im1Y
5cfa92pvom2pNA/KmUzfkMcgkR6H2UNhiDpbPYoYjGhz+IgGx5h/tblXia0MxmLM
dR8WqsUkcoUXVG/jPHWzhJPSsie4OYIGmdnIavVG0WxqPhiFKGu22cTntgAQPxYJ
bY51pqpkYL5/fwfEaFyz2zvaM1ZJE3bQOZ+TX/70HkflW8bXrioaDFiVM/nVXmtl
gvE/tmfB4wtbv0lFV+6KCA2/4C/r8mcyDqmMRchGtYYYT45hVYxVqfj/F95uxXxp
IFjLc6NlMzom6ooArOqsc3HLNX2V8dG5aNPfftRzdIW8KdyKHh8YsOQYGZtHqVKD
CklLvPKVFoB/j63OL6+ZYEFX7mTuMfYcu11SKUyk5BG3Zw7K9cDFC7L1VPEWTwJq
FE51k25fxMA27m4AMTAgqjPaxk6R++ImCRWAs0pmc+3ROSzl7vhEe0G27ae9D5uE
GPEOXRbso3m9yZvdJJQaC4MT1RKrYEVXrYEewm5NNlHtGKxouv++Mq+96wxSxdNt
5gxmXrrdNUsWppWcTPgq58QuAiUgsn8Niz6+bFeKED5a1APT0FqlL1bR4SlFIDDY
3+wNAKtcvXCU6PtVOVibQeENfLi4gh/xw5agyXnHhMBQo0vAG9eUIp5t4If6O0Ch
1Q9+4YBTbXbCnj7dChGq96qV893XBzUnGQATPNCcH1qW2nKhinHDDcAYjo+XChp7
XP2kQ8JE4yfJOOz3CyIseasOZ2iMeY71o3k+fBS15SwSw7UUHvk4FmizaELKq0Dy
rMYt0TL+CbAZuwkTCtcIlmq7/IWPdRkDLc/6CdrYPXeHi6JAGLzKzaXdHmcmOW/F
Ohc67zh4udg8cG8yPQMks5LGkm2u/aIlt7w31ScJaXUYGHIJQDyHJd8YmRsFHl4m
6I7RiAtJH50T4F3MrC/vsgOwvfUOLAeiICp5uHsB8b7UIt8hwCBj4RB1h+CE4GL4
QIs6RvskCtJ+PcUbIedS4D/23l9SwY4tpVhbJMzkk9LSKxy+DO0nXThY+OMYHhAX
v5hOZWJJBFZ9Fd93xX/deYzE9DvKvnK98PeXDdCnCv2U1o8mfEQdsQv21Ao4A4+T
7k8qJQmkFzK5dp+ySEuJ4Jd7Eir+z7Z3INeKIR+NIMIUO81lhHBrevjtcotpnlKq
BLlWZleRY1grsRwINjFV4W1wyCWxRo1J44MEZdJDXipxZDmqBPM40hnpCnHZpDZW
Ikc1WYlV1ZGHPcIC5q77Sbtyj+rgIboENFSyalO5lvZ5hqgFD1pNuhqCZSMTuKUD
4ZFL+MEw99PfgP0FJrwuf5TvDjO2BPgdLVXBH7W2QH1JFXoHoHTC3d17J22NifQU
mv1G1NowY2kc5re8QZ46+BSvuEo9avZLg9cQxmXGbfxALSWdycGdtdNWnGtLRj4D
OMaLddLEOV6ard12rIIuJ4Ppyzhob9gIf9cuq8PJIcXfBXqth9p7e29MoyNqxw0g
I/pzefhANm19dI1HpopWhtDj0X5FOixneBYsAER5l02nFe9U6pksJBNG+ryucu9Q
l21e6B8Qrs4X3zZ+aDCUEGXrNUT831ImfIgxStRnIwqK0uy49Iek0T5Cm/a2nKki
swLaxODlphM57tQlHxqzA9C9Ukhh86hNVSBhslbYHBYajtFCZTBlKcMtFxfZiw/t
91zqqnCps75PWja/vZznsXHNb3Vhm2cObF4/llrMFdTzm9ElIDE4bZSca9y1tebe
FYhf5uXaMsMO3SoOZ9PByDUGB2qAJVghaR/Sn/t51qLsYrGSWLI6cPrnjVcTY+K0
Et9k64nOpCSwvjTcxL6fFvzKEn//veN65/klQHOUsnf+kujZDiSkmWuIPVCY+aCe
AEwOYQO2dhZZB3EkKAYugbpCKZeVQYathn2ZMjxzyoPf9mLQo/FGCGcWrjO4x6ln
n47GQC6JaoZr0qY0mINHBHiscBgz09BQcpPoeh0AS9GQao/rlqLqMM+Jn8SV1JtG
B7YhoBbD4hLKVp3f+xjbQtVg+/4DWMvXCnFuRv6FLASgLo9FBu8/wd72gQecuvpB
5WgiXu9s9QpNTdRHJVl/0pjx5FwBmdWvm8AgwBUglDQ0eRpuzkVmgcBXOfsntwyc
xbk4Qqw3rPLsNR2c2Iq8q8MCCxeyGII35rDyxIQ5v29zUryJgMdiUCDcygVnsapD
XPTMjIi40PwaHTijc7XLKilk5B0ZpVfPslny5NxFVgRANNq/HIl97o71CIUw12EH
zxszHbtaEjyOlYDRyZGn2uV0mOX5xhBdYxZ5EeoBgU0CGCD0vzTy1k4e6lsoQvSO
4bHj99hf4MCe65LrZHZ8W60I4Yqub3EJnjY3tiG4Rhyoo9aQOexXqd0x1WpDOZgP
aZoHBvl88NgOmZje/y8Tot8ZdpM1itEjNnAGvl0KHFlNeGvYmPhm/IkUvKAoOt78
niOsPwIh0fSz3hKDNamKgvT9XMobfI7L76xMRge4mbjuTZgCc8cnXOHNIEIMnWR3
boCu4GtPG//ndG9pOe7NHUj4yPlNfr9817tz+uTepe8pwaUuP1Qx7XetqDZcKpVl
N2n1Nxp6r9KbLE0Kqd+n2dUz0wa42XHfro+S9cWhOmzBm3sTI2D1DqLk04yOrrIY
xbcLMO9ui/G/wiTqGxJmRQLnfqw6bt4IOcp7+El2U86CA8VVcwPxjMh8RRVtkGwf
dHNmuzbRsTO7OtwBxG1wrdP2x1q4QKJSWp1jlyegxAx/YniwlWK+Q5c5v3WwyUNR
4cLxsdSJTehAHEWMttMk4SmvQy+hdpUMDG6aJrZAk0E3qsOBN3m24pbc46JMTHbr
ZNpntZFJ7RQAKKgV9BWdoqc4ZvogiRWWQM1awmYgNy8qne9eOzDn5RWCLLfY3mIL
BSTaiskriVpweiKrdMQXjgBFXqtGsagEAzqK8waVuDDtf+JKjgYH0f1tYoOBp+1N
SEBPW/SLVa9oTuppH8r9M0woJqjEU1vgGJ4WbzUJCQ7B1JgNMrhNp+Czksfnrw2G
rRpfqv0eAHN20iamxO3XPVEVBM6PylybmqleCUSWQfSwcBrGrcwiLY0LFrwcFICw
Q/k/aGZNUD43esRrlFNULHA2u4A5dQS/+HQhHWBunoNNQPfpef4Fb+a70g2i0jig
2cRjy96GJeIonMRpKbh3Q9gxsaaHnjNVPWSRhe2zoL9nbbow12WlYnJ78gmism8/
PUMOawnvy+MT0Sc0m/vsrD+5KRLSQfWqxgS73umitBP+VCr/VJIrK/rsiosX9rvg
14rB4wIrzY2OcQ3kAoaYiO7IpTy50UNJX0U4siZdIr7XJLA2hx9Xw3O0okpDKW8E
MrEL+fGC/9m3xD7L7cpn8JlPcaPVyVkasDwYsRPXl/Aw5Wsyv/H8ku9Y9Hm4o6tB
1B8f8fbGmG3WUux6kFoAOsdsfTuvMYNiM5GXqcgfJQ02PRYVDKIDFvCakM/c0E+B
bqdb2hlMch05BxmpG44Kb8qwK0rGn7p/ImXAVrs9v4a1sFWcyd2lC0PsemmLPMjO
28bU1/bvOGinLD+BF8lVY+rpRQzj03QIVw8P172yjOMYcMpGq+CMhact33t6snHb
ipet8FSOXv0Wmb/vKzeg++2G4FzsycRXYn4yLTifYi8giTn4ChO5aIuaMHonXosv
4su7KNWSSG06yVI5E+oLRFCnT9Sw/9Okc4fd2IGPLlDwc8rvFEl4PUDIK6V75hP1
xsJiQaY19PdsPCIaDDIHEriyx+aIT3+DolK6GVEkYAxVhsCXQNjT57nQltHxgn1i
l3stSwQJ5L+U7v8TC5ac3F5JAtwvMmXtbcy/P7N5sbwJ9loid/2wRcEMPeE5iuSw
VU/EcEfDOus8wyeUp+FkbTrzM4POsQmnUykpNWv+5tBPxKz3CckTo/U2zbzLbcWj
amgKRjasrnoXlOZMV1chaX9khyVn79cTgDvgfJBdbDtazQ/vTW4sN0aeoYjHas59
EcW1vs0I92VId422mWnywtYKHQm5AsDjrRmj8eyJrHL64kGEcm5gJaxhQAbHjBBA
QHU5TkdGymgZpgdKkRfsq6yBiSpVkIOpXokB6sK94FEygrBfnM60CfJEZqXwIHuW
RqE4SdjlGKW6z982xyQEXah8c7l/+UxYDt31r0nZdRA205Vvcc12ct0WGxRTy3LA
nGkVw0O+XIInC67syKz5DdCaCXlb7KGS8M0/NnbpqCRjlHPj3W0vQkowtGZjFJzR
/HcKK7X9KcTT87nqZ4XyG/DM+T7GdTl418DTxv7ZZpnkJE3Qyw7vyOuknAShDU1L
/InMFE3+uTOoOkj6YZQqexHaC5rvMYddDpix5alaTR580oc1iWrZkCpBgb/cGntF
ZyXJZ4+eAX029sJUHe339Bi9rS+Bg4LKAvgQiD32CMSnmZfRKM0tQwqTvIQG+CDe
spL2vGsPzdMxtPeW1/suA7RC85zd9bOL5sDn2eKNjEx4AqpYy0AeN2HHU+0GMgTN
Ojo0Fa28EXfoNj4lzRWoK/NW1fqSoG94EsxXXTlKsv+7fa20Sm/pLwsRQIIcjW2M
neLldw55lubKpI8zNkScQPjxtL5GdOvziHhuPyJLKfxS8fo4b3LMeSYYwhT3Fm4x
LUr0K+TnVY3GnSh3WjSo0UAs/mFWf7HYldrZSRo6aaw90M7iDXk6wZD4soelWmCp
Lpr7cGg/1tQQty277cxeoCgfqVyX1XiO9Yc7tfHLMqleG4Cs0IOlV4PJ98BDGypg
ua5B6YzYmRC60BeXi4yuABWQ778U+BYMMYApC5SlAOO5aDVCzPQ8D5J1bJlpmo08
SYpBE70uviv54pijI/ioMFdZmI4itRgzhLTAAmLNqduHq+5k8l19uKyi6FLKs7V2
3OankZ9sD92FgJFkt7aQO7ELtVZdtaHt1T0ceZuyLq2j2W2LpI4zMU9y4StuTXCi
mvCE1hUHAc40AOYtht84cqSTgRSEXaSRp/0CQW7U+eoOb2Xsqy5lgXrJFnkYFfb2
zN14GrBoxmU7xm/4n6iRhBRXOQHEUB7llxf5+RK5y0okj+pmZX+YnDg/le6K8PN8
ItgidVz20PwqmNQ27O0p7Y4T1lEbVcumoGOAQyeKGYdJvl49SHziXTGCxBCCdILV
Fu66C+WUhSfaBE0c4XV1bTNvuOXQaf1+0KJ0mT7uDv+RJmgcrsmKyBaHsdlMngu0
SaftXS6lBWHokuXBudegq46gQskr3+b7Ca61BnCGmNUAWuglw72/OTCrgB8OSbji
wYrupLkBQh0i5oTSVd+wsCvMZ1EpEFrC6qTe3LbziQ9TlfuLkDnJVSXbxmobm8+N
uz1pMNp5XEx6IVc5JO0XQGNdaQsThbd76BElWygC9SvQXgUXcEQ8RENeMy2vW+8g
KD2FqoGkdNxywUNvHnywZZwXcOeFA4wqb/nDkjk8jX9TAu7pnvb5mPLpNS5AQWwJ
Y0vaCTCaEzBZkT2eItR8FNoRYyZv08cvgLtvCqFdwpgnVAtBTrc8IPvC7/MMMe+Z
ULSvAA3l47klcTwgjYoWGdqCMfS/TzgkrMRX3EDW6LloU+AxkwH0awzYr+IngxG3
wRXgDg2alDUamYDrx1oprclUos+EmaraFKDipe9f4jLDtqOeu8/N9yRQH4Bkk/PO
W2WMUmvL2pjtUHt5MnQc4q4JlcPjcdEX7eNfYIjDPmM2cSODKeGzzheCw5pmX2OY
Dl3mbtfmidQaIF/ZS27+y7jj+1767sWA3CtNEpy8riRaFAmrQgrP1J3ao5VIztEp
HpUgAao2rMvYYS2rvNzaLYJ0PuhLJObeXYCBAjg6/QBSwFGEO+N1f+7JYpy1V8Wr
nZuRcQ8u8Go8n7SXg1q+0ZaEBO1AH4vbkOOUM4Mn/lDpTlxYM3Vz6kk7JaSzqBEI
PuT/qvgfL9T0KaqmSJI3hga8VONTy0ArWMI1d4U7SIiiAPO3cO61EyKjYt3T1+yW
ZDqlzcAjT2lMjzWo+v3zi/B9nRFnHliHeApQAOZg4AmzAs06N8OcIFXs47U+Tx95
6ug8I15kcjRZWKkeO8V7liugfu3q0TGUgng0RyOw1omCs3QBpiZmQ3HRP9bLEjC/
D/LJeHHa4SvJqA4hlp3x95upuViPa9/MQ0s2qop6DBBnhSuAYs70U2x7U19o675w
iYsf7S9JqqV2z0paKDWT5NSZLRc0y770qaz8/IaBQJXZ31S/HqEf+2uzABts9xkG
xj6SNCgBvL2QMIaVMMBrKrkLtw2Vk3VBBiUAn5hWLgoIsnVp5O1ELrOmS6QM8Iqy
dz/pK2agG3gNuyIpbiesqZ83a95lBJJNVPG1IqzdTrnWjpO9mh7js3EiKUmgnhLA
wLyRxlziXg4nBPHoFSIjnoaGAQDRSHQtqrFVq1zeFKv7TRlOk/WokPT426ERXzYo
cjK+morhjVPeuU5Z2EefXT4b3EfLgBvQI1QWGEBiRsSWQus6ck1Ubym9e5ED0aXt
IDniZDQaboYbUs0kIatlzPXS/rK8tlWyM0UhchZfZ8eK04aPq+qjTqtdk5l79kd+
mxf8iwRGqJcxEpmXxjDe4mcvjoWQGGuNsdwKxVyykUR0eKU0N37GSxPiZwJfg8lY
emdgE4eMLavn86WBbro5giv/bJE2MKB5/QsA1doA9bxw8dYWWi7MtS0mIBOZsTqr
Wgxm12V2/85/ypzHrJwQUMcPjTWZehf0ivt+IzBRMFo3fgGNOoGh64ZjPbPbHwPL
wJP9IxtPlWgcH5ke9zH8PppWQApzeAeGyaZ2r+v0k+Sbx8Am8UizsNg6CgmEgBcX
2lk/ysZ7wUd7LHaIsykulo3aS68MeHApVOvmaUO6QqzR0PNtQaxEe3W4IX2SovFc
E3GXJ3mVA5YzgP/4NvTsABg6xbfs4ffLWvTeL9ibKmadHJ/HXBt4erPf3cpCP8RZ
Od3RVYEzFNbKcKfGV8SAmm2JvWokVZBGkuki+qCzJHBNyDUB0C5VGLFeLwE8UUYa
0+OdZKYHpJPoYzfuJY+0H6rYg9K0N8yRdk0IdJYlghqdpMJwM+IUBBRn4No9eEVq
g5n4PW9VPygIocdpwzJzCHefLLG9tYAg0YslP57V14lWRnVmeetPHa9N2IbhAxCa
OiFuiSN6eYoYVPObMb9H0EWEsOcSBbs8JK2HSJnMTuENqj90/INul/moNvvmw2oE
ddgSFbUdFbomjbl7KUIne25XaA9BV16fLyBH5+qwdRHelG+7JvtV7ky1pRP5F42r
K7z7+EmDUtTAEnzNMW1/9ti6CkR3wsTB5IkZEHviMXd7yMV68GAcBHgMM74x72GY
0NIkFUtl8bzRc/k6nvj8PUurDV6dYkgejFZOi4SPgc8ZYsjcO8xT5NYk6PmFA5MN
4oaQFVZrRSVfPYde8DxxZfasUkpPSkJmZvZIAAWN1YgZ0V4tF751vPrMzCUdRNL+
0+oK2GHODa0dCYX6YtiG3avyYvQRDY9nRuqMZT9fsJupXs68ZAi9zoUvGNCAOCoq
NvjT8zctSblVu3RGfInu+WWLwv/ThSgbkufec+ySY07mhqawTn/f8qnC1iMeFb95
fvDF3KRW+VOWY4orkg5wASLY36nkZ18uodPlAxELZVP3cOL2F66jCkzEFbd5Fkam
dsILQuyZPOh8EG/rHwNBPajoUgTwzq8gQCfGfRu2rmYwxXnDuEAvzIfGfpqW5Kfd
F5dfGvwVPBqu1NsMbhNjttA7lNhD9nUWljUjDf4Sv3gc8DvdA0xyPyqoftkEROTL
fgDa5pQ6J68sNf2ep0LGQMYrtBZarqlozOk5tMaHbq1QJa7swbnbTb3Qi72Sh2oM
b7jrT6dt6Yz4T5ChaFLC529CPhzQSSts0PjMAtFJ5kdXv4Y4qwILmUG+2CEnodh0
ms4BtdeSy1Kn0IH0eVCB9PE20lSkvKF70ReBAUnVVyYOVSD0wGdg0J4IDqqoHjq5
jfxWEtU6BVwRtpArhMPr61Vk5EO4Qpgl6jp48DH00XrugHKIFIp3THn4vbd0Bdve
mH81Kvm41Y4la8Rxd9W/GVJLu0Yy71vAe+MtVRdW5L9zQgLNK41tVupaT7eFfrg+
WiOLlBEWOZPnDK/rwIft3if+5fbhHTQQ5uY08OqY3wHdzmbOFyPzIEAWOVDPtdz7
9337KDuBBobwZCcrz3dxb4GvYCstCjBEca2DpJVXOBVpEDlRHDN14rMQjBwrAuy+
t96GFUX/bNpDGFAsLBP2vVvRCvMeJmCYEMIPe6bVDr3r6rGD2Y6tyeNRltk84CE8
3HJSseXkogpkAcKMCpM/olg9+0NYvNrpETiLuwlQ9fYcFvTuYMYf0oL0KNfGeEwn
rvclpvFVMToqj9LM6TJDV3laXB2cJjFk38GdZeqLf34uUqYv9vFG6HWbvbLWH91w
7igq0LBMKiAfvZ31lxDupou2Sj0REYRy4AEXFNHYL2MGyiuKn32nkHKaWO9T5AdX
nN5R5h41dM1ORWiyR8cl1mPMcLmke6vOKfL35P2et9iaTKdpl4DkscVxDj+qpLQZ
b9UtCuPQsArb2D/KYC1AguyEc49iFLWrASKYw/5OTtPood9OBepTDdeAH8QdPvl0
A66iP0q0MxK5RqVp1SvUfFVUb0WWlJajnsZkgnjfN2B7qd9dTGBJpGm5oVbPosTd
kJjyeVEj09ATmUsRwewnLwb9N4KhqqJEubVIYfIRqcdVyuyxBTwFn2QVW3rUf9z0
RlE/7yISVXZcpSru5KHscSIFTeefXVc/bGcj0tuHSgAVyE665/Ggw9Qb0UEP+v8l
pgB/mFmHCMIZ89xixryh/kREQm08PRdTKwqx+vxoaXnZdXb5B3bqVjBKlKlW3Lvh
dI9RA1pI8yEY7JZcx4XNvFgnNp40Nmv70y0vAPN1tuyd65EFBKM5LsTiN25FbvRn
NjNDZFT1tDy4KsOKMAYmtWj1TSPjEHa3gIqPRcML5/droi0jwRk9KfUteF/WfRZ8
CBm0WH1CJIpaMHOe/RtYZNhh0H1FYeIcqvmO21ixNnfumSduRdGAE80EivNrEfOO
3ajTmRmA6OeScNkkTtKqpGBWwOPccY9i59jdMu/XH5iG+RH3ITuHpd/VsdFdAWb4
2bl9CNeiRFSk8WpmXI6lPHXjqZEJHEl9TqKZBVmvImJi6lJTpYi4Sr0yLj5TuyI8
bOXe8iK4nWPxl41hVmZrcQlCbbn4FfGR9GAiN/rv//EOdpxMHubJslJycwyGAFPB
gcQ4KME59DPIDxqT1Euuahqt5ziulOZejiHi93/0NjZyE20os4Zy8hSvwYZPV8cQ
71Cl7wrwCcD5X22lG4c6lNODvcQkMGXlLLHzOyxph1aRodRC/7gUiLZHoN4Xf/x9
QtkbHKMKHxwCxnfkAleiz/nxu6soMvquPPLvGTPzcUyiNWWWffBHboGr4NdHZb7c
UxGEygkULAFVvmN2pSi3CyaKMBGOeFMOY3g5UVt0u1PEYtR+GNInUC1a7CvrdwLX
tiwXD+xIiuxxssk373gsqcFKjBYekdEMvDKkURavCW5XKNqvIcnTQkcLZBHeyBta
c7z/0vQk+o/sCHILMTK0M/Nq4KfJZKEzcQFCI6Tfx6U1kme2y4Lt41laPYluiWTQ
rg7IG+i394n+G3QN579WiOY5WWzCO+fFBKRAEA1E2jrnGgUuGrFa2HWSdmIrrCem
YPuWc3yf0jzbNEvUoVT2ejk30rehyLjqxr55OUpoy2xpEwOoRJZMLjp3LyqVCd4A
bsv/CGHf8vZn4DYR8E8alt+bYnIjIzFyRNy0OSm5u0ClZAvGM5i7mzVHeZ5WFspF
A033IoybyArmr+F+8dmFFQmgp+n/UPCxbHKxKMyTO+pltewMbDa1wBfUxiXb/wDg
mP94BogM2/HHw0aoNf+a7SZZAX+VWEBQimM+VTWVCu7RhLlSbPJD4XX1A1fitFHY
U5ag3g4LSQX65IMOfyD0HH21CARD2NUTTJcphhwChCs8F3Ejfgbcaebb0YamOQlC
GhuhULpYX5v3eubLw+Rna9XObVK5plgVvUshf0la9huLh07ofTolO3fjsfvcmh74
aU4ClZQ3asx2S1QUe4+yswzUlrD27EGLQfnQ0Ao3PLkCmjZVXEWXQLSsQFvrKSpD
LQefN50lnz/7k7N4GuEDHSWqyKnZ839Er9/dx0mXSsQXVRdKOHV6L8HRkKhLipjT
DxdMUiL8nAQRNTXXarcQunfQSDPIkT/LGSwqDh5bTk2pz2S3dExdtQlKEWRcVDhr
Zk9t0lV77r87CKR5gtqujd/MSgZ6+gSIJ52qhHPXkW2ffK7uxlKBJUkI8cjbxrG8
wxfthHsoAAmh+0yyDDRBV9yJPY8HF5kI7gV2D2ib7Gn4hemN64a5e0BNkM3/R2Zg
hN/1CGvbJCrw2RLU+CLjRtN5X93zqzAQRNzNhFZjuQ9R9SF3wzMOS5IeNSyGNHRP
qIiFSMVusNRYf+idJd4q9mqo6gGiBXi1V7Xgd/If9nPDwDHMp7Aj5W5dnoBrLziK
uH6lS3GZVVJSn8LTYAI+ys/4pQI6FCt5DG528HEKhgtW4KupS9W7rzwG7cf32i9n
u1f+n2H7ZBvJFK5xlQkC/63wQcwI6z0Ve8rn6PU3nkDZ5eKCwNNwuz4Fh8CzJq8b
nqY0DYEbpnpm8IAEmNhdnjCP/6wiu3wXIZfc5BVchUFQUrIwqBhuEIjTrvzd6oib
K7qxNc//LRXOTKzbLu8SD4C8eU80Vh3hdaDgLZMqXbj1AdVQ14Jc/+Wu7I7ywDu1
bDnpcZrG8oq0hTOsaKYX03Z27BkyEBqqY1RDG0Z3ycNIlPb2JmWAiBsXPPLGveS7
MZpVXg2EKkG3KHvnAbv97UjTud42zqs9SiwfkgjItuMJ8YuapPpd4duOsDYz2o12
oB4X7JLHg4Lvw5kqO3/wKXUZ98PGIogFtkaI6/LYPNF/VChlXmWMh1ji7/n6Gl+C
pz2t4A8GR2gWxver0XXpl+QXMWlvKeWJdcRlU2zMrwpqvYGr2gISab2toRTRpXTL
AWPeEVdX5OzqCR9EzL7xMI4hh+f7J76l+l78VDr5OeyM0N8RxBABz1vLl0Y7lKip
0htL3HLVcgDKFlesDHqA5RTlIooZPzdcoknuirXzi+g2vSO9eNrqi7HpKG84Ui7S
ABM2dJkoLnrSBDvHz4k678acw6mD20vRmBoZEorC/+UE0E0ZlXjxNRrLZH03EKVq
wUpOVE2BFDqhfu5pfjnLos3rRL4eeOq10EreAGvpryaZ70Zz5UppurxptAOPsYEP
Huo7vL2QtaObKrsPv3S7+1YUG8pm2zxalpOlhZLZSsDojWchnFyT//giNUG/vjQw
klpcL7jeIxbJA5f+g3P54Mygp/bbw2tHbePBXTmwk5fB6di8bP2Fh7vY/xCx3qWq
/Hfb7GIPT/gPppG4yRPlhxfN4ZpcjFr4m4XEpCzU0veNBAF74twYF0McnP0QZeMA
QaWnS1+04vgyuNzyXhG0Qz106Sb0PlEMfvEp1f6opW7cHOg7LSfdL3bd2xU8KMHy
srJhLx894RocTEB4YunOpBMlhfGk4Ectl+PstQgoS5Gw94fwCtjWqJQ06fZ6r5cb
hRbykau/kFu/+VG6MyKG/a/ei4waN/SsBd+IJuoGGxV3eV62fxxblLEb8tMyzX8u
eHzlubxGCSG4nlOD+2u/QqdPJnaxNN7/aAZn6pEbPsiO30WM8D8kGwJm7Dm6/etk
oTYpljoZoXpp09YoG3483EJYGpxSvF73oN0EnDXB5V4HD1a32FNgQX+H7x6m5umV
5K2vXMsAUGfp5fGZj+LASLUsyihcNOSLSzLVtfvJKo6zTJMm24m41dXKwaQzMmrb
TDLbixaGy1YSgMZavsdl+LDnWu5FBL9CXPkeoWkv6C6Xkq0ILF0Khgl+jHwIl71U
HhPxXXkc6fHyw3emNE7jGcNe8JoQD4o2zpV58XNrp5fOh0hVCEOigZm+8cfRX94x
zYRQrYUj6Qym4aDUB5H6INCM3Q8Z9o9Wrsl8lKJiJxxPupprO/w1AoAb5iY8mhss
A81OfpYzz0R4tFfxgMl0Nk8PdEf133/rm6oTWjNJgthhnXodV+GRFFNH9GWYMJLV
WNzqbUYfydkh7VNbuWuILI54J8hi3481RVOg7gY4THycXvwuKRA8h2mpF+/rWkDq
Hd8Oy+RISFWWPmUCX33eNXKgDnGC1V/IQ7qcYYPNA9OVOIKqRUGfAw9j6nbkLmba
LCnR9jiMzavvziKz3LadbYrz9OvhFllHzS7jmRL6/ot1lT4XHeqrb1Yj+lrWges/
v9Qe0tChdgi7X4rMpdJ7KB+cZ+PM3Pe9D5y7M1/Z1wTpDRpXoe9+Z2cBwGlv2t/W
LC6oIkbwg3BBodyc0zwcpbNNUWq8ENAQMQ+3bBDqC4RWG68KSshUJUN9PNRiDbub
IFxGXQ3zgPD8T/5GeMjtcTtXEXLK5xdnFCCBy3VavzB5UklOyT3DzgOn/wAr7zQ2
LC9hoeuE6kZ3JeTtfPDqnG+kkqYpDFimzIaP/fQ4T7mnsq91Z/dBcRzHbHqHqqdk
hZ/eILYXQFRvNvZLMG1Zq/2a77ibcnO3ScB6qFCT5LAhypock0ZBsej50G8T+p6V
dzocN9WZvw1JCT+oiOZCRHnXDVvnOQrSg1369XTkrtI4NSjGdQzRIe7u74lAciy6
4NrndC6H5YVCigtttbdEatd/RfYcUicl4aakta4485dkEAKiCKRNuksMrYlda5uQ
0TAuyKAJKjHaCuOaMpfTt7csm/sJzGCSWO5LjWvBSUxMtD75LWvLihkj3qgY5neD
3Wyj6sBSExqYunykTEuEbLhdhe2nKFJz8nnmNgWHdwjklxQ6+XDkVyAeFdGEWJOy
OpPMv9yVgvaIYJjW/09PktISkgdl5sDiRLXBH7+QM4iLhgUIwcCEL5WeZTbd+oLi
d683+ho3TG/PsR5WwwsrkkwP4yoRL01zIVgJFO8BMVa0YMcxp1AUo/T7WtrID1Tr
SHl4qEY17ci3Snz1c8BaGg4ZoMIggayMjXVThkpIl5q5jHVcVEyX2tEki+qTD+Rj
fzVN54KYYcGinm7qNBrfYvscHoEncatncgh3sqJ2/xabjKU8O41qc5W+ituq73mY
JhrWWuw9tRrVCqkYAIZ+eGhNsaskmSRZG70FGY5HswHUTce2sVJA2ILZYVbKUdjx
6eV9ndGQGAkaINXRpWsWvV+yat6y2LWD9M4KvSRrwQuT9eUn1QleqIZvSq4KZJtc
1DWuC9Bwda5iT3k0kqbGu//5zScNFrQwp9VQD1EEbo8xKCX94LpPW2cuX+i39/qB
LzxV05Qu0wkSpM8fvDp5I/CaDib63jHDBkwyt72LjFWNAJ9bPaa3S0BlVUnOOIIL
fDBlMGk3Vb7Yd78o4ZMIQnEHSeT7NdFup1v8aJ0m1NZaa/qZvAJMre5Pqv6MEqOm
rwRKh3c/p5VywYf+8s1BKn40j0HWIoTLmSCuyen0Jr36Cg24/oo3F8fGhmU6sY7j
XJqSISnp1QwJE1pxmCb81qTSD5JJuYidJBOuJSeJ1nyTIxU0aTbBvxijPZRLL6Tr
FE2Rpf+cJvseWJCmoef27/Bpd1Nkfw+z2W2AqdXTz2bAMvRZPob7iD4a8/kwA4eF
9ymNC2qEMd32Yz1HU6silpUHsf20A/kWqh14k7NiuB//JrQYy8PX0IJ3AGZKsKh8
zFFfvyf85wVzB+bDQdGqG640wrsbZv3xYD5L4dGnlI/Kp0GcFuCA2emRZgqZ3274
IoX+CBwTL3P9vb6MH2Fd3uVSMThGov+zzugG5Ah+UhsaTEXmCk8dwrhathojcWmR
g6oOWnDH7Lg3Fi8gKGePh0LVdC6rqrvoluv5vc5pG/cHjDZTj4HoWzqqQOgz4Vzs
KHsv8hs7kgqGyXdZSV0ksGMwFLRKKKrXzAkKWcHEXDOhwSBUBLDdz6Ghwj3e87r8
60D8ohKKVPvXQCxT6+EqG5xK384CfICYvk0iu5I28cRiaoVhdPz8qtdrcro67Tzz
c+gQekxd+0Q9XcYFWS3eYzKD7uchaRTpSD1YwYlSIupejXN5mE2RPI/q3MMd4OSF
6AvE6T+n1UiyBlnlia1tIq0R65VSlyTKTF1qGLO/WY1+iyXuJABPWutCDkEA9sQ9
BjaVKRwBDs9X7qet8E0KY/mNF3Rw3/kC74eM08jezVACvd1F2fFj0JaU7L92emo7
7GYjFKGVbFyvdnBi+mG3kz6o8yRqKhINdHXbua24yjeZyQpIRPW5XicCuNmh/YLJ
T8D6ymOb0ZtamX/v9LTs5z1pCPHbvt3plHhcqrUxEatOBW+olpJUbJ4bg09tfYsH
qXhhs65bONV/jT91+r7OALie5KyLWCS0DRUziXed4QDGB38N1hhbsj+rJvIrYsyB
fKtkkRDpuZc/PgOMrWkpHRo5VZkv00qTrhxxKllgg6cqt74QnnCOCtWDwCqAF9nA
2ICnom6UTfI5wH6+mUEXhf+H3v+asDcLKpvfdRNu5KFbc+Zx4BXqqSWijLYrSnFg
MS+rMOTVpZVObsTq3FSG1+dfBMbT6Me7x+Hu0OakJ64Wop+ndipIdhjlbkxNxoN9
H/k9DZdaikCmq9Mmfw2ZLYFFUbJs3NTzZZe451NKhep7jXGIBmoAuyK2lChGx3J7
GRC1FnheUU9i5IPJ1RBHKmHhJVodiBADqWm68R9YJXt32V2NYBk4Mm/FFIf08lLx
zTUTwbw8DkKsgS+RFZGjDVjmE4oGwKVCwtgnkDEKR3hNlgzEgIML/JirPnXMRl7H
KrkKRFgsQupa6T+KD/DpzhdHi1JLDTINa1gH6b33hoTgB1iyqO8APzdu37/rsxuP
MDJ3kWbLxpZJqLcN+0R/+LJrY1+yEXDVMdGiTLIPrBlXlH2yMffPyEpohn54n3Kb
X/PS6r0jneNCky6Jlum8CkHHKzQlOZcttpEFJ7RnGpcgIiA74LOUvqx3Z0jJ6PRS
sJqqZZEhkW1Tpxu9bKD35/8TBZ4MiXVgwoGBcAAeGiw7ibP9GvzUutyAzvpEQF8F
SgDerVyGQ8VE9OD9BSHxKmRGjPXpcyj3pv9BoDPkJR4OFb+vCBcyu+f3548dEhRW
ACtWoKT7uV6eD8wCluzSlSLWhY9/doMaPGQ5dPlo2b7CUe/LqlXq7mo1B4V7Z7kk
AeSnhaJpCAVyZx6/4IjwvKvnHBlj8PIyC/YFzbmQfGqjm9X19iI0s2NNCUytTdGs
y6PhTmP9O9KnZ7Vhc0srhQA/qICK5NnFhKTZcQ0hMa9mjaVwAAQAkoD96/K5kLGA
Iig/em+h0inIErHTlS0stO37CO3SoJGy12YG4C00SJ+9WrByM9lQSv0ryRufHOOw
ZW9lsfuDQE8JgQqkaVaDyKKW6MJMfHakYJVE3nKGYYfFfXoXEcXCl1h2z8Pmnahc
8UGOF7z5XPflKI2l2Cm6sGFdJA6UGkgmvYGHXhv0F65mp4raNc6AT5T2hEzwS/Mz
qG9Aff2iALi6yRIyCdaMNa08kVED9iNYFDKx11iusF2t10glE39xYzSL4fkYQRdR
NJ6W3W1MvdJbX1VEKBeQnVL2ZQrcgV7putHri9P1LrwKQuly01vlFAbmTIRiqic+
meneSA/U/P9SAPe3JldyAFa+VG3mJ2DClYHXgfT/+ZGli3myA0f9Kzro/XBa2bN5
nRpiCLITS22pLLOBiaUnk6kCxLr6olxaqeGnjsgMMhb+abf5KpyCyyuNSberQdl6
g5lPE+tzmJvohvqAC0O/Zz/KGnuXlOPeWf6FJT9QJDRZ0EHPl3MtD3EtBvdGEXMF
gumCIfkf5KJ97xxNN+3Wb83W4KGTmgt2fr3U12m9keBiM1ys19RA62ONumouXkJz
+m95BgIYSFQI/yTnWcpVFSpLmEoCZ2Cm2+dKRb/9U0heCud3VbvrZgj5nuNbQYVB
CUcBeOrt3WMDCkCkRjd21DBJI8BqAe3fOlubbMADMgd33tpom2vDmXzYoCKtzqYs
/1e0DydMTq//tp5n7Ok4TcnzkWmUazN2pfpxgYpfwhMnZX4RLbznT/G/CNjZvB57
mQ5D50jX76uuTHYEwkClKWhFbP2ivKxQz8SL7+3L182Hq2Ou7WCqJQuBunp/aUEW
hTozaU7rsYWC38NlezxycxsrPMOXkXKOhjxb3g6opnYcuon7+C+qPSQhL08iyjn3
pujlvopXAOw8Xj7Kg5tTvO8HDwCOZCAjj+G6ZCEMCYxscGjhiuVp4AUg3vQlsAsx
6XOAO/NxYwzv0lrV2pQCZ1NsGorqHzKRYwuUy99lbGOWU+Dsd16moJS284v0zI40
SZC33VLXpxQPe83EicoeXbe6KPmBMIysXhS41tu1N5lNHDA8hQMPwIUmkZEoKrDJ
31d/cizaM63VdrRSN7hub+Om5aiEYqO/PJGMKdPbHW/m6YLXhcDUuOVL1r/1cTw2
ylEyFEFeYOdREdSANm2RG+i+MzfT6NCmFXCw0J2FJ6XE8K6ddlx1FKjPMB50IZOh
WUWm/jmISsowc7Bcxmcm3T2hJxvnlhcRkQak+44MeLwQHVQ7vm0euvr65VJHhpIH
J2sY2g8uDyye6xmuFdFQdGLWsJlaUFhH4gFl0AlD35OQXXW7UKtNmua0ybwimDvi
3kyuSU00xcrmTMA/E3GmzHsWrFzeRbUTb5Ov7Fmibqj/JFjB4UGa+81l1Ho2qz+5
Pntv/YQF8YzWV4GTh050ZYXn9dUn1Oe4AasXJM90aEy71b9+1l9gcElIPzz5XZmH
1pFbQH/t1QhD6+yOHOXG+IMjELRf8YIoiQfW4veoA/c7U9PqQaeqvgjS/gQs7mac
VWw49R+95R1icLzAzjCjBmJgMkjm02HYE/CmwcRIMkcZCxFCJpkGuoEkekzS0hnT
fGwLo/l3QPM/59dgKsx4+FCsIx520WovunlYYubzJ0lDzCodMKrIlVyIC0gX89JE
dj4FPuRzvgqi7y9wgeTm4sbuWROfboFxkq4yX5aaPqwJzcpmnPTPuTB6KEDLQLwt
2M6XV65U1Uu7nSqgWbokh+1+snMR0xTRCN4qTfkS6w9CH6tbtC3wVUSGLjW/vag+
ta406jKSbaGJYR8087q4hAUHT+m9+uiZOuD136Wp6+GJjHmhTWIcGjKBizLl89EW
rMP3nET0I4W1hNrZKLb7Emc4F8F9RcUi8Lhj4LSEFfkpFuUjrR7C4bQLd/O1JRU2
13oq6Kr3bV5ac2YAIv7RvqkkejzX4POrxXY6sqD/PcglgJ/d8McAjptx1MblyszG
izAWAQAxBRteyYjlPJQCfbY9jJivVs/DNwbf5ksROEwR08Zj073QBuAHb7NWU6+f
57HoycGZ0Yuia+nYK8dI8VMXZ+6CCjCRPnx5Y68VGVJR0HmObh6J1Hvd7wg0L7uZ
Z6o7T5PIkcqdV8wxCrdfNKjuHCAFPqRhqHXIlWKTRz3SHtTk1XaonOHnEOEXzdrW
iA6E0Muoo1QBRP2XwsKyrlgaL1cAUm7q6wBU9AYxs5YKrscAqD/xWv6j6/0iam7/
1wt1fja+5zJLOL5SYFIjF5BwlhLBGzOc6njRJ5/NGXcngBdwOOwRVaLuSm8Jl/Ls
ffIv7ZiRRWTCXeTI2NczdxDjziOIqRuWd74w5eFVrzj1RXsxBGksSyM05T4VRwbr
sEowuaIH3DLzu8grcJ+Z1/eP5l103b8t0bfWvLSPXrnPggi5qIGgFa6GYYmnwUMG
gsca7lQbEuw2QERoya948RDzR1TkhKAMxnMPnTyiIQ2O9I8HE0tXF6OusQzsTNBs
LyQYkIu15OnA0S5/HoYQUK9eqc1Q9bFqFFm7cTaGtf0cw6mcLoTdg2XX5+MD9za8
zY3qML7djhLL7Q9Eva8SKgEwQgDU8Q/QXT0wo9OV7GcKks/sryWuNfUeuRN4mg3d
jE1aQ4vE+/6dl459gH0b5V4O50TBPcL092jKuNWNm98oR1c5z2vRfA/EwpF/tvW3
9AleZSpyCpgA2f/HuyWvDDT0wLL5J4aFKFzojjhgj/Rp8StB+JAPca1+FzYGYYM5
ux7YRf2q96j7yEZXXh+/ORskguIJdB1H4P4A1CcAtCp0R7E3AI+T6/F30c3Kv6dM
minZWUfcDfIdRxZl50MJ+Z5hLr2qR7L7HOwULQeNk6ixZmbfNm4XSPSzbCzbZaOt
Y0/tClEAzY0Nlp3oSZesPnfFH/+2upmd33qAmZqZ+E0Da3Y3YUpIQKGsWOH1ekEx
euD4QH6ym0Rt0TEm4hpCbWE53PWlbjtOoKKS8+HDFiVoYqMGPwZJwIIf9dRIUYU1
O+ZFIxBxOi1l/0xc7Z9dtvlTrlv6rIYF2eTu226vEbRurafqV5QiNWPRPLC8NmoK
JYtx5zxxC1JgV5pggvEaCdKPh0ynFm7tuIW/CSyuO8Majpn2f+4l16tKEJzIkZII
5mCPQIW8srk9QOsgdvCQ5UgoJU5iON2JZKl09cNcorBnga1IDM+ytXb2h7J7zM/K
eUkSILNH05eN1W5Vh0rCXWojw/3Erz8jWzrLZX944Rrs9Zg/uRrMG2YCp2X+w2IF
z+UFyUIshKS0UjO+qd1LbBLvSnIhioO66r3RyZdZvtXhtudkeyWS/VPMPe8q+0uJ
HrT59qjaCT0svTBGoIst9iXdyeGVfrUT37mHjFEa/mywp3W6VY1GaVplfqchJoCU
p359yRrcPGG3pWec7StEKa84n/A7sF6aLD2qKKRTEyM5aI7yQ3KktwwpiD2m+xmQ
8Ns4Q6iVDY1sLegIUJlhrQj8BaZ+m7tajK/KMLTsF5nxm739IFQ1z6Qx2gUxF3/M
OYYtwJlTw52FjYyRqAcpuJZLe5q9hMQwq+VIqUwt+x4zLO+8R7XSlwGwawXjgpmN
gqZffaMQMvkuiZiUcs6yqvZ2JqIkpxL3MCaKCY+4pA/uNITfdeWkD8iH9xPWC/9+
aWD4awEOlR/Jk30LPj5fCiCtZsSrqyFh/Vifl63KFS5COOuYdo0xMtfb0FKhEzL9
aVo6plG2OMuBF3CpqsdQlREzZTtinenFqthXLzCNCqGCHX2e5IThPHM5FfLBh1vk
ErMmZi5SQ9pQ7LTBbTmh731UyEKbdrA3cDhFC4DDLWauftrTDVxBdo8WzRcfH7Nn
OE1lhC79oDO6yetn9cNm2s90o28p9iT1CWmWc49JI/a9XYRyWUahwFHKUNgKEPxd
hEgeVGQdjMO5gSY6JpGMJgilwGIixu54BZKGDXhvNFDrY9dWv0kXbjRQrAbWl7Ab
ctUvpcpky4i/T0X0eSb29AXM5CHMvDbK+oy2quTvsBhun3RQM/XoRgwbT1aiC9gf
eXZwmyX/fJA04z9ebBNEk8Fok25E9JQ1S27CR5Y8osK7CD2SakTWOknIFsnx2FuY
NuzXLux0Tmlz7cWgVQYXhCwwfpXTr4/sfpBTEGi1GDzx647SADIAhadCjLDK0kg4
mU7kD3eCaWpn5jYZ1S7PrJEG8yGJ4b9Q0w5bu9u0VhpyZ3NGPT+eN8URHTpIuRu3
UaFWlXpLswa1JuUPXqUl5wds3BVO+6umWBCUifVo7ugCMwq7gknGDUvVdbCH5I+0
UP0OgZlWUh9YFJ4P0GWkCV4mrjAFqZa6M4i4KYQ94ym+x1DNgKEvrBs98CIK74k1
1EdQhblOD2LDxpfKQUnQ2T9V3wAwt3bZAZCcVSiWJ0EKg/D6QYz1wOytp6JyYykE
emEbmjtOdsj9oatMjLTJ+EZnUOXCjYvvlxZdC12ipqFKWtlM0mgz/HGXD8XwWkq2
wuZBh8VyGDMpWXGQRUilfRfelJloRLSb6gj3FBnxzG6Nw3pUeZzps6aYtGfj4KN5
L56xMkaifcQcB0ekvls+d0w4bWDN92t5j/TnF4FI71On+nYYKuRq6z3q0jNb/s6h
WTknuFo54RPCu7GmzcSUt4Jq+Od1ANryUabUSWwPkvcRG/rJf9bgUdOLQzxTzNJN
4L4qmopNm1FhVhkIMxt/WiTlvev6/0ZcPPMYORz9zm9zo0JHFoF8cpJA5qCqDwr0
VNGAspGM/vLJC8huTIT/2+syXeovJq7XsoQvb7VidP5LHJY5ArajxVYqCVrOC0OL
rXdbCRx9wSKDiNZ0q7Gtw9cwfQ7kKIPmIuDYlK4QtmQZe1A9DJSN2V5J2QeNzasF
0ptRUR44Pm1t0gEm3du9lBsCDafNd6lTshWisp5LShbOTi3xgPOcQrs0Qf5bq6G6
y33rwZKho7iivZ57Mc8BOwX6/3zfm3bvkth0nkDd1Ua3IiNItZLOBEyri6UMHv4L
J0S+lhhGKRx7pZFM/B8IQhauh7C9SQF9tZB6j6N74TsYT3xsVupTRHNeJbfmYgLu
wBUpDEb2dXkiEdbnYYkuzdgshnfCUEFu6/vqe43zqGQ35zlJzbxTySbUJb0GghgD
0jwgenIbQIbMY7NZEsuT2CxQlZIyD6JnRXuWAJHRh2hr8zIDtpMlu3KKF1yG+Wug
Vgw0vGUkpTrQLF/mf0hThWXKL/tTlLN2UugJDajyHdd95K66tEeIO8jVcOV9mE1X
QM1uZNafSMpbh8rDLLR+Xw8u8ISmgJHAyhq0k8femw4n1N/jLeSPtbTkxu0kWYEg
n2kgd6D03rLYYKJeNrey3yPGYpfTOR2xnaRf8MMEp9hebbZT5QFcoB/JGXduDTwb
JVUcq7AjXyXtSM2q76s3y8lbJSIHiLm7IlMzqz0Xc8E6B0RMF/ZKOn5yQanRowjO
CnJdDV4gKpZoQ7vMzGid4p3ppUkCFNHU0elMYkoni66t22+Zgl0jPmzum7LoH9Vt
YXBEh+I3952qX/EIsok5qUWFGpffotbIErSQuYvKuYplclu/nKZiJW4AL16dvJRv
beAOCJlAVzsmvdt1flENbsTtUnSWwcV/b/hB+d92OTj2uMjeVmrZ39MZ0YjFBNig
B+ORjJLe9GZuxO1TNmLcx/y7DytcHQjwdwpMSUP8cFjnr8MsOUEO1AazVDJRILXg
JIuXGozBKESm7IFd0xc5OtDztRr2WbMgypu68DOhWs2YGb1JToSEAl4x0CWU42j/
gfQaT8aNdpCw49e4m0O/AgvVxNopK4QIVbdz6QrOv+xZm0J0L/XFnCmbcUggFDOy
j0gAgQjyBeeLGX1fMPphEwKeIJFq+JlSv2HDGYkQJK2dTTMcuLIVysjoSpN9ytIZ
kmkB2V8ZrCCHO3N0mFfmWtK5zF7IlgAux1aGFpEhkKmhiwNDyHNumtRo65gzcQOu
/jtnU8wprv/CGGIHHKd+BkP613ShBG3S3SGWImTmGdi88teLHDP9fj+GivyGm2RW
peYtUBeQ5Mx5jK3myI29JNmVHCXjiywQ5JsKrYCs3MRBPAqHsvpe3LTNn+bI4Uxa
ZPoi+QwN4vXPGkYp3av2kESplpDd8Axz6ia4wi5dKqPX0OIhEnKz61n4L/oq7U/x
Y1maUpKnmLIA6AVtKhPys76d6FRjQWGgL7GwkUTU3V7j/uTkfE25B2Z4RSzSoD2W
GuC6QMabAjYsGtH8Ejw6KE01jQcX1yryEUf4Eh0RwZNS9PglrxWsDCA7Qgy1mIVa
1E3mvqIdqeNVHhh80fGelhYUAqGcoGQmETJ844zAPpf+eP7pKhUuX1zp2DEkZfUn
yY1wXMBA6lgSI1s8ahL4k0ZP2WFLobJqXQhJSzVT6akV+2/pLqJxjJVwL/SH1eW+
nOOqSwQyXCKyTipt4qmp2d+p6K78y9eN2lDMonRpl4lZqGodUCuKejgCqxTPB0ud
EOy+1vHVM3l6t6+Ph26hy5B45PNqe8dsatEGE6C5+/G+alqwZwAvHUhSf0yTqrRI
w9Kpo5M4iud/WcW/nztNjAHYU0wNgyuNWKAwaidUxVKfniX5KFd33ToZ0PuN5Nhw
bbmL7Y+Tf6CMjCPjxQBlgEhNHK91Pktx4KP4auVPNhmDzCp1Wf75wghQgMluaMBc
+RSuoKpdRADwPjthmUa0clpHG/yb92NJkU2wCgvkcN+iwgDbhXiOWmqPA6utM+Is
CDEp3EviIDe6qxft0ewqo7PHmm6b9LxH4YJsJS2sXFAaOtayV9mxpXi/Zntmdqyp
aqDYmI2WD/CFR7ZBSOCQryXflmIH0SCZTwfqDRukG1+mJ2gGIgQnavQsKI1+tytW
uX6bLJcOjyDR9D76280q+whvTPywsNx+/i93zbBTERnSwVmY8XUcT3p3DTGeKa82
Psm8ZOOyvxabkV4CxH0BpOYVV+Hls6ifFveJuNyqsnbAnHWgoW9ArSIJvrMHkl5M
tqDUtZx+1LroOyiBk9gPVLG449mwZj00zN4psJ3XcnqRW1gHoGwbSNsB1GYOIKgt
J/SytPA6qUgD8795S34Ryip+7eBjrPbOh0+A0HJEqAs4cg65Bz3galKP8ygteNX7
YC/AMKMWjtuADf5SSvWdjy8PO/qJMkY1ZCvwkdGMVAj6J//xuTJ16NcT5hDAQIMb
DAyOlNAhrq0Uq5vNy0wEsvAjE2hv6Jve+Gwf0UvyKLcFz0oYVajwkWQNmmAGTEcY
vtnfuO4kGMgz54UYS4RbP2rXr+IOJ5SCxBhDiojA5kayVmKLD9ptsZlZmhYJmrbG
GJU7pXuaGRx6DB7fyVAzFvdiYWTvybbFWV55jIRaDR8naLkA6N32d1KALjMHh5DO
0xDeor94VMWGM8+YA/aYmXtQKE2FWrRiwHT7FEad9hpZc8FOu1rxYQmsgcq3Gi4i
UnAcXR9EM9Nhzrbfo3VdOM9qziWoHN1ATJGQT5W9EM7a6Ou8zrzjIr3Y5KmU1YZk
lPzwHDeGNoipv8QZ8TRFtlJqUXITdlUCv8hAcyWWgXmBIVEcfYVqN8fVAXpfWDAt
ELRY8+elozXfxRQKPFmQonjSF9jKbTWE8ig1h297A7ljJzB6DKPwbbVsz4AefFIZ
0K4HV4DOZgGWEwfBmr4CHcLwI172J5gINkt0liQiNOpmSi5SX/jSCbtdRh7mQW9X
fV/pR43Izou0cR1/Th5wFPHiCRkVoqkKTOndcNU4UNEq6N5fBQpoP3pAXcJzgJgd
SCb7Dv12KUtml8dZLtCh/yBlHsNUOoAAzF2BtzBnU66VSb8qIFlDV5yXj9SP2v+X
aCS3jr321CvgfVIqfRcHUoAV/cgHHTyb8OhT5pe+uJ/d/to1TO8Y43VJb5Ys2FRc
QC5BUbWZFOyZFX8+9YeAOajUz+1Md8qxS75JrKFcj1H68qenVzNRExRubAQCFfMo
pbbqyvWgV5VetazIOwU+3L/rd1QXZPOoHvS9aJJLOSWlrwphLqa50WN0IHGHswGg
rrBjAXoTv560NC2tRh9siPw/RkAJNOjndnoDgMlSs/jwaYMmuFYdt4oesOzBlYnE
C6IZcguXTd6Bw294l3tM7c1OkkY3cfDwAPglz8GiOZARpmIF/BRLvgD+i7dJ7DkD
wjODFaQVL1Poj8625QduBjwo05mEOxe+pr0CIQcsXT+x0irxeyhEJqN2hbbbNXza
WeYmZZpm6sZwSqY8QkyyulKp35TZXRF5GNBBZKXfv1l9fB7dUA4C42xg6LcesRwd
28EfRiAw4x9R434YBES9YJ6mnMrsh6/aCKJ0oq0miDn9insn6vHiMyhrpO3ARZW4
cuRQ9EMutFh17PEqWXREHb0Z/5ELljsCdFyPcqjlGu6yoTaTTs3f/RZEemnxSu5C
xJd0tbhlHgWMd+IOaaxCRAPc/U7N4z9M6SLgTgRf86YpBEWgAgJ39Pp8U0ipyn62
92Gxpo7PigSfmPVDsrSEFYIhRIkqdLgnXtPfZbwUbHZRvHoRz5F5XIyrd1KDh4cf
9Ye94+K1dMMx/GJ4b9QkSRegHLEQB6Wb3nSlOE3lxZvKBb5TPpeytEMrPncQv1JK
l/T/ihFHFG2RZR47SpPPQ/Rwmc8QlmU3zckmy/tJV6X72GxUqCAWHlSn4no88j0T
wFMt7GZJHRMpMhGl1E1My/0w6xNy3jgoq5f5sROgOm23sISVcgbstVFUP7U2nade
c44ENTztnAAWsFEltHHAuy6BYKLo7bIVKK81YK2cu+CaWayRLdZ8kzPFH3mkZcc8
dlp86WsnxykOJO1s/LFtqlMPk6qsbGzLRElS2O6sHbfmEYCNNVK3LoVsU//ik/hG
BTFd9qLWmugiK3XQS9t3CH87UWhgUK11K+l2RDDA9nv8Bl0fSuZMQgV4pl+aNYa9
C99iI/MZCYR0SpAdnM6zD1SEqQA1laRZjxkdkEoJzI9eYhsPMmddpP22aZmAGoDG
5Gzyq6OA5AifHZl7vrP9qV78kvC1aPRsECOxgLNJVawrx1Z4BfWSiFAgLsaqfVOS
q5w0Kb8nlo7Ti0Yr+bxeeHdCYCn3PfIB8CTVBTHdhtIvyBlPP3o+RmGIjEPvOc1b
RZyKYI/VuUKyhCvk9gqlNdgzLqKRf9Iyk53pjX9AIlFaIxXCXou6K98CK9wj3RaQ
nKavnItFGffDnzyndmlT++PC4igHVs4cGNtkIHttnJY2oQGtChgn/LE08QeDYkm4
OEqbxbMf/bZrc2uQtJhXm3MxWe/R0gX9Iwb397scChWUyU3aNBGH4eTZdcFXIm34
9e2lHOr3xmh9V2ch2rptmpyGNc1TrOBcpssvpeWNYdH/3V9H6sCwj9RZDDCFo8+t
r7l67TRcv+QpJ7JxowhneJWpp2tW5YgcacjKxBMay49SkisV7CRg9O+KuKdHsaGJ
SG6EO8cqF/XsBe6gTR8oxJhG6vk/Th7bmsqgEajVAHWKq6CieLLxvZa6Rf90RRPO
9pyb/SjmNZyyDDQU7gK0MluDuaIkCTvQ3O7VO+ho4gZMUQ9A1ffh0GoqCePXStNY
uklaKDqaMdaeEVLJiQJb7i5xTkrZFx6YbLq1utfNhthBcMqKtI2l5siLsfx9B3B7
Ekk5g4/O6a3c3MgAHVLj/WQD+oqaIjQ6u2ImoaUp3EcKRFP5sC4QIh7zQvyd6AkG
KFgz0WOqKRScfdIU7/wEwM7Q0OVSHK9qtQHA/rn24a4u5fWzv9gBONec+G40G8b1
t5rQv5C3Rdt4bNQptVUxo7vxBDqtZvOFOlINFfB5Hq88PyN2hpgxGbabMsfzuOit
PHhX9HY2q4DOFfv1eBYkjOK4Q1atUrAR44i7btpNAtviNsK2l+jvN5sxAvUics0j
bshFI5QgmS2JVGkY/Ef42+C2lKeXB99/v0kyoXN8PpWrwP9qPavGqPATvt/TR74i
ZG5OQK/VNMntKnoEIHlJ0TDypQ1rQ7BhqTib6K/c7T1EYQjFSg5E1TEx63I+DGT4
ldWMNmksCJMs26fI26LDa9jqvMJuhfNg+aRYqFfpFqBmhEEALBTOD9a9YHjtdZ2M
bmzBNDB7KvRcYI3WNWfwkkPt41BvaIx+xttNvfyTd3Yy58T38Dfllg2X7ZRjp5vL
WA15wAXDd/d+7XkJcF/kYWTZPjZ1pQ1aSamQix589Fyl5nw2Sghh/fbU5UgEy3v5
YV09ZR5ifxcaFGOta3q12HYitnoJRj7jNK+2R9V6C+BjD4mWP4s5QFIebwuLGWks
fwtDRu+xPh5FghUHNTBWJLZSiVlyf5vEI6uSU4n2daDQfh1JD+BKu16LQQQ8NFvi
jDsqT8WY/SjRnQOoB5qCBGid0ylMpl+OH17qhyKvo59UCWAQS4UVGTtAG7QSUbtY
LNTe4ebbe4TRseKyUdd4Qo7/giGdAdb1RP5YIA1a2WriLRPmZt0aWU14yfS2SXHA
kHlLQ6M2SkYIsCKmAFjlt6Z7sDXgtj2yy7D3V3ZQavmKmUNV/LJeTsQSUeKtAUZw
sbIe1M7Qx0L0wwWwAwYSWSWZsnGIamKNxZougKAO+WrYGEkSl50BwEv0/lLtdFUD
GszGdXxGwkH9VDTtbRuguWAmJIpabOUPuOloSvg3CuFyMYcLHYEJeeOxG/WXlFQk
nWUCaGjWJd/tlY+zC0AkU1V5M4ohScmfQgddRQup+NzGTJCrxWi8U8MSaTADPE1O
9kvIaX0MMdbr9uwfGe7J3OtYHk46M7CpMV+WPBea4EkraCYhGuJcdbvRyylcBs6V
abs0tj/mmW4uyYOf/hMi2Ps/iUUD2yp+I+BZlGoCzrzXiVFw0DJbX5WZXrAjDHR1
euRe14rwCcmTB99KD0CLAJ5MBppbovNqLni0qGgcMdrzwqCwMF+0kssgMh7B0ZQF
YcjyCty4hvijRsP+oiEc7OIKszabgVwjuOjw6Q3r+VYY5LmK/EFMbUk0B4xewrN1
9qHMc0/6/j8kl4hyDiyTUg6CAglWp2qz/ey5hTssnKTlgZ/VQ9Qqu6Ycv10izPxc
KVTN/TiCtogHBclhbMThw+6kQM9bFur0WF5rV80zvy7uWyYVkZ6LEpEnQz9HC+Sz
ysobPNufcQHgYywDOa3WqRG8X8h1nG80i3N6TDmWSupc/eEG5f5oiCIJSqLIxmkY
tzyG1gOPtAJhoSeknZr9x2/w2gSSzmLs3hw+VgjMK/ZkQT7tRZ6apt04rUbIpdM8
aO/ewVSsv8kYddzBvpXpGQisMiGtTh1Dh3C+ZcrhooZJSxagMnz2hKbu31IdbSMv
kqeaDNpMhvyOKkA24QM48Sh6s5TxJRVVk5jd8NFafsLCNCOs4a+e7pV1ATj6V5sI
PCzrTXRqgLXcnr07KmSzo+qtLmNDo6HgFOfeLSu+KWSOs/Bd40TNaq2lxrc9QP9/
y1wiod/5rUigCQQ+bpJVuolvfprL/V1x9tUDZsG4jsHih22rvgc/0/Cs0IN05I1u
mpzyTfgrmngGRyCeSAY+DdqjmAZugj2+Pyqk/aDtkUWDPgozAkMhI/hoFURdJEPU
6Qc6jfotrI7cllQMol3ozzUcnYEbrTVNmUi8j4D2pph8/7soEqQ+H68ghpUGhuRH
jzr1dNuVoWD4Z9fRwCh7gnQJryvgoQuedKIiRDToRhf9JxCYbVX6YAU2z6wQZtpX
m6a4nUfF9Wk200N5Kqdy/8liGEtnqirlzJ/B/C3lZvusJBA0pDqcfQMPsCbcdOUP
qZCUW34xUZK8z8RcOYGhAfHF9yDli5CZKgsT3zlaI5gZzprdnqucvucJY+gir6cH
r8xj470gljFKVJbEe81wIMl5CXKB85U3BusWD1el+dEO0IZeIA9YCtIYICCW2qT0
VyG1x89eeTwEzVUXxbM9367Q2u3Cz51Nuk4rQWXjM4ZPXmkTs/UO87H9vNZaKtl0
j+bOxcfOF1BF83iag7SOUdvge17QhRfjaYopAoxEF4kKiNa0Oy8AYExAx3ZfnRaj
n9NwFhbDmcEuHOwp6FnBAKCOfT0T1J+jZ2KPAFFKe6XC8aohN3TCu7PhRUkya5ak
gY2vCCvN8VrSOt3oup9TMsMOdtELyYry/NSyxRcF3jQZyfaMT5KYg+eDtIqXRhkx
d7G3vmXC5m15+CssdXYLelvXCuKS8mdsT5K3/TWOdKCs7840QXYgT+Dpxj4GR6Sb
W3Do+m2Zy2cv0KRKnuURkYGxh0sc7JjsNi7GdzrEr/jA3fzuDCi1mjpw598EQlZg
pLv98j3RBECNlLR5fzsXKlUO+WRlwSycR1DJV6E75j1SYDHrBzdEb/wjzCi655OM
axHo9n5pEHL+D3unxhgZ78Z28wa8311VGkRKroc6pYXjgnLxT2h9wfcGF/PDXq3t
x6ImxUWTBA0Gu86G3ezQ1OCTSg9wuPJPycvtmeC7EFCypfKdQUQbrkFWBMWYycrD
lDJqtQUYG00RimWKL7siUg1LZqAlS09gaJ6hN8t+5k+d3gSfYS389swzY3xP4n8j
w/xGUhvjd8ttHMs5pB/1Ac5gN/j7guqDlp1vEOwfIKssHaV8KS4j9i1fNgNnUwRW
XA5o+A/t5/VTXbPLuFLkA4YC7iK0Y1DcNS5OYznj8LC9iG/qSf19geovr1LXBr6U
yuMahLV1nJdR26Rq+dMQUM3DCqc75U43gqpFmDuOGDCzSmJQmnM0ZfOY7zj2Sl6P
KpeSCidpGJjUPMIMmMukiR5WYdp0kWVainl9CulFiHHhSh62gNNS9Qm8+GMQYmIG
qd+M2tcP5SpoN/Bi7obnFUm+7qqH7+zYNdR8v45YSt/sBH8Do1VBnfVcreqobGXj
0i42sCgKc+4Z2vlCJoe8UWb3eGyDcsIeu4/L37HBy+g8wmuevd5gL5rdDS0TBXuN
qTdZe81BrOK85zEvCJ5sdWcq4jXkMVoJYHLL5tWWo0s8NxKkG6aVBXgFuzzroJxJ
39BpplbK++T71Qb60ya+NwAyAMQLsI5AhfjRTQMnLJooaIidtYm4feR+71raStPr
pOenmeivRaIxv+zYvmXNXQhPKjLYCtv9jWp0qSIbtX5V63qEISgtH82GGLAdmqvL
Z++u03C4UyCr2hxoF3FWLkv/kP7QtcYa47w21px/lXiJ1EpRhj7WH4hArGiFkScb
2fm9A83bo3dh6UT6zgX2C9b9WpYiK9I/p2HBA56UoXolj7xypvSAFb1m84bWT4iP
U6FsAZWXPH6I7GIWdC2nyEmm7Rm8QO5RIB8v5V3D1uLXN/q+bVYjaxyhMut/O/Is
rJK6zZFZNK2TIk0GtWsmEComFDWR9Z6cl9Q/twRndLd2jh268Ur9edJoi3y4NROo
JPGdN/2QaNYiE7cV//oV94EnBTiTvcLyw9UU4zEwwiJaH9lj8FjjIgRIXMeKa+wL
7Z9PWQJO6psuZcGBoGV1NZRp2qObgYa+Ff5OiZwLSY/A8MZ7olJqJQ5E+KP/DH0l
bEG0j21qLJAtytL29T+Ig6cjiarWUDSTxbBahH8xJujPFesNrFPackLsqQc8k92K
HCD7zuhkOqZAXfzuqRdIo5Po9NxdktkLMfi+udH7lR8WhaRrnyBk+IvffgeVa+7i
forFlXcNYIGdy940cUoz4oghVQ4jYsvRtV/tRn+6Smc80SobU83PDvnueX9b//IE
rhzX65GbicLFGxlvfw6sIGzKYhWYxR8H7WlZx59zNTASgFjfCW10cof5y2C3UcYX
7zX81rTpWG6eRBeJI2CRRPseRCzwSjBTZQCKeOui1C9WUjENHGauO2TzXdEsLlBG
9KaVFdHw116ibG7GqzdXK6Vg9uonopnT6eB+y49fjrWZrdqzL6oHMbTpdEqZ5j3u
kMgNDRhiJhL+/E8N1qbl9SK9dxOyLJg/0z+dvKnhxPcjGEXNDBCzZ3Hm9PyGOOvo
WU0WClvZgVpm+IRQfyoXr3Bjp0Pq+gQL8SpvuWW6dO575zhNc1JggmO0tenizF22
Ht6A1LvYWVJQIdDTdCeIWXmzU8/gkAbnw1DGEZr1OAPhXjULeN+bpjDtT6f1u5cY
agkh7mrAZAbdYKQRkh2ObL54apXfNU6eWNu+kJNkW9SKdsNhoJVYLFrJGV8XN6n6
wmLjLA5pFg8Vd7wki/HNzK/1lhwck1naNi6W1cm1Ee2GtRCZTkL0hXsxzsDEDSvT
AYpbl9toTWKl5TIh2fzmmUdMF2za/zwAOkFKsDDsi/mP4EHG9+QB7b5/3b94m/Hd
AII4jWMfrJNwq/5VZDKGFIMzeS+LdCqrGFuk5bJ/nQmBFJHD9O6NIa9Pipk2l/pV
aBpHw6QPcShtt3DqloVOZPLM8atSLSvn0G6SKlgDru4iMKcXfcRKKAy6EldCsT+Z
B5JDoem9SMQEU1CS5qOBdV3umCsbiQh0Ldqpl2qOdxdimUgTggkhwKMnFd3S9DXQ
9onBc+WdMrz64W+X+E4FPvMbyq+tWnzPZldsbFAJhDQtRXNBRlUJx+E7WTex8ns3
lMK4fNnJx3xyK5lww2ZB1vcHoon7QZLIHZaAZdPbju4MTvN6cVS9khg5tKOWWENV
6e4erxc8fSpdpxH3kJtAdyJyM9Qv7KkNq47Frecn1AsKCaT//o1oase6E2h3g3xk
mTsBrJNSToXoBpI55cm91FW7A67UeU1Iamh9x4WYPfAIr1II57rYjYS9SlqHBZ7Y
qSTlbsIVmY2e7x4mIycbGNTuwRJl6rQSKku2omKAdnj/Fyupij62tS1XZxprZO25
8Cap4EwLISX2LLLndm3eknFjjgEO5Jf6SulAfZKcKkpNVsu/2qXZj82pmwcRXpcI
a2sQjG/PPdnT89ihYLlBgB7TdaTScf0JDrXNZYmnFMIYXN/jNWeg6Hu5lA9Vtlk9
QBsCywA1dxZTyTUbP5+u60tY/jns11CVv14CF8DN5+o72HJZLZkWHJpAq7+2RKwY
ag243jgxOz/C+4dDuiwU87yxjwe8G7SZMYtAo9YsGvywHX9RW2BbB0cGOGsGJDap
AAqFl7KdyCh5Tmn+c134nkExmgPKShCzrSQrCcix5iDR5dbQdpFSX8tOYylIx2F6
lWt4lrKLKhrVTuHa/aIjNrcBwImVHEzWeX34s086PsDPLo5xP/I1b6VN2oRoOssW
XO009jslqU98XGR3/GXqfcC7JrBk/B+iBuUUb7sbtbAfQYb9A3SCZQ1zAcrFY2YD
LZrSHsC9fJFnC5YfG2MsdvyoT8z2yPhJtt2Pr6KGkAsORslY1fJVW/evsrE/R2xN
BnLDHEiiejMnbyjqVgPd+M2Dy01GhZEh97Fjx9Xx/lvpjKATJ7SeYpdmiBSM+DWP
sJvQNdtYuQXYFkWfkoypEUHJkExS6WXOtcg/OW867uUFEZ6q/Z+Na2t1+NG2fQz3
3sbUm9l1LFu+XeyFRWDTN94g9cpY/nf2/0tuYSrwr8DYVBQ+/AbZ1RYIHu8PK0+P
ipvNcNME13qMIa3RInW1vRIy6BIOVXCBfIa58gvShsbiHbQvlMjopna8krcuc4pP
31EjmtwfP2cNipHEB6s+DHKu8XGjSXgGY0F7uHIwditI5hIZtJm8F5FNmdrzjp/P
6RVVE5chdnMIIUYXWXqTvjeHzy+uZl5xMYzbAv9FNNdPdVGFdvOGhXxAxMvPjVRi
zkogMuof/8CCCFU8wDnjOnUA5G/QY1fQcuj7hXtRyKwHicTB8r+8awSizBwqWC2x
TdWdkJVAHEjuE4A2ikwKfAGeMgyBFLRtPORO0ZaB4ARSS8xAtJs6C8glM/DbzTiG
rW9VBpSOtpHiTL/4WvH/b48GBbJOzNcTavaAeTWVelcWF+M4gODsZJx3RNC8GpzO
0ccPomGpnHnBuw1pzmcEuIYNy2HGjo+i8BPAXILFeWuKASuEdlRECIWZsxCSxaEW
1xbb0+dZy6zKLPHX8eVMeD082vlGePnAq3W9pwHN9imr8/omvCtPPxWaTcTsMsG0
vMsjgSWWsVZAIcU5Tyc2kaCAfMsBPFoac90b2CiQuhpBG30O7o2GUr/kyPINvxb6
x7SQweNhPucKZM8mxaItbko4kLV6t3yGN6jR5geT2hXBtGj9WFp2/KbJzsT+3ZOh
dIIgdveJe3dppBL8uAuG4eBJYKWDzYIsLRBsSwXc2mSa1N+mF14GA1ZwaHJvDu+5
LDG+yU0eMirIt5Nj0bBPCyBr3wORHcioMfrQyNtzfHyKuRBEge6GLg7m4Si0M7xy
5B6hbPKrNFrQ0QP1YLi1I8MRJV58ejaa56Xkd2JvloISVyTDzoiuUkArCk5BEpz7
LBq/Dd4t+thlzWNdpBpZX/BayQE6y8+DEzs56Mp5CvXfHt/RTKihWLkjk9tTDwKH
ydP4BwBu01L3zH0L41Cgp1aeDdMUuiVgdlDfIlSvdwm+PonjO4LcBs+yR0SK4lvB
sF883/xqehNKBdUjeCne2gLdEC4Aq14pTl4VwBSn0AeF8XZe1uvcbdYTAU4eEdqs
28wUkPu9yFmtOiTqBZBjVxTh2YV+PCqkwQhAoHFwq2qX49YweUBQ0R/t//a+owvT
Sz4YqMbkC1y0+AMiwvZnWFc8X1WG6tVJdP69qdt5GdALoQIxfZowNlNRoREVkTpb
mkaGkXglkTllSHCkXe4HtthHUe4IDulbK52gEMn6CMt0VS3Upgl7sL4K2izXK1jm
2zmlP1uGVgVNKQz4/Mz1FomGkUeVsW3ajUDfhpJJe6PcpE/NQgVJMh+mW72uHjPL
vF9UZHO2XHB0yMe4PIN4YViSjYq8X6s9Tel4E9Q4H8wMDJicyKWm3Nqw2wqXfAXH
UD3F2LNIgoB1MuGZ9JZkwAIo+yWlzajHgsrLWRSoa7dfjFDJNdBFJAOftPalHfN6
ZkvOohcZMAY3msJREIpHhP/dRygWLtz/5fpqw5qEyJBnlHQLoGwoMKDuweOhYtNj
Vd/6HgEqrA0FKh5r0uuh07Aca/55JK+WU7A0Rwe7XVLr5VZL48V8Fqg4zQZmBrxZ
vjOqxdjJ8EOHV240PuK5SpP5TddNstX38bCi6gcqQJvlIDTCOrsKIJIF49n1Xg7k
/2yWcpJveUPIRi7+0VrpSgRrhD2SyIhDiIbWEkP/u/9wrXQ8udP5enD0GREeXyO8
htQZgpNmxF5oYsaCbj4cg+O+hyiWKDqSOfNpmKPP9cV25Xu52vkoteupIwdopvGV
4O+rRrwH03RaihS9Ft9+VdXU+D1vDx2M9kuMU5cB2zKPsnNL7m9PIVf7493/WAsB
ELtPTUTFlPc7iim9rARqGU+Tv12WfEBzjXm44XUBrIKmh3x4Zf4J7HNaBx1AtkpC
+B67XKHV2GTbuO7/99T2u844SeTt7PWckME4OuFnY3tF2JdNmaiseVOndU0XF4xH
BqvxOd1uxFntxYWQ0TTtW3A2Pjc0uxQNXoIYawsD+0RVE4AkCS2XfA5rzQVO9w1U
i/HBvNmLUgwosEYZYV0C4bl209YcrqNWk9j7E2gHYWAF6YEgyVKq8g3xSyUgp1o8
3LQuppKJYV59KnX/uRavAKVN11hI3263J8HwPs+XumbYFqecXDoqq9uhCw4qRADm
8VwHMg8s5MRKieEDkaygtiLsBAkI147MZevXtf3gMWaJiRxVW/dHmUzxtJPCl/9O
91cyeTzGXXW/3/FukTF3/P6xHv6ai3HjxJv99p8AjvJh+Y9eHJidh6gWJRGp7rN4
VMUgCScXG7rmMZFXHW/CqphEdBlHu4EB2lMlMIcSdc9iHTY4H5I+TGbuLKbcHElI
Os72+/lr8M2ZeFTBTvqJUaWjqE4/Jo9ueknRkz+LAcESSe3sjkh/rsdKGf4Ljfe7
3igKWo2PLnOGv+nHOLY09cYQ02Ay9a1NwRimdwZElCqCHutJMD7dcvXG3rXNIZGI
YqTDGUoqlUWHnDdBW5g7haaU8NMXWFNrMa496TKyhZ8gceSutS+NQdqwYM1Ete9K
TDFhYNKU45Etamm4Bz5v7+Cs2R0RCHyQ+3mX688nqcXO4La0hUGkx3nnRyX9hJbQ
01B08ThoZBfiB0qxhHj0Mt46drkw8DbIXjHojnEolDUPRoZ5kFSTBhhN0utYyWmi
m6MnKPr7g+MTzmR3JxEApNyfVtlcWNaNUydQ+1LuNi/y6fe1Ikkh02uryoVeQtCC
TrCaONLf8h5hkQ+zqdQVZ+33YW0wdni9bX9QmP4nOlLxAsR7VzBUAOSxlK/fZv6q
Cdu8Eh8lWgSjFC8rnDUwkWzNRLL1Zb1AvnshiPgXsHH+8expxZCJ71HRuyZmw4vl
8N0DIODMfYeNk9RVPkVXOT6X8Y/O9yV1YgT7DeyAWKxyl9T+JyAEdaXRa6Kl3xIi
+iWy38ajdi5ezAAZ61ez0NySg7CT+tZ0jhjYQIMybq4BWVSrN9KXG4CE77gxdcal
6ST29+rxnqbwWNC5GUqlcbkcY1Y49T6UKoYQGN+rV0sjEA4h3pmR6WnRoCiIRjRT
5NwS1JJyDkW+ZzG80zDD0w05Yb/ePjFLAKoVTAFkEDU7OKIwPC1ATo+8ISGMkrrd
SNTz5JwpvEMSWk4eWVV/RH1odhnXFYP09ky1RuP3BXotwDjG/2VvFNFhqwpXsjQS
kGlJKy2aP7AtdOuJ7qcScFCchRuyIIISsP5hQXDrlCllCq6OXlxpjHF1Fr8Nkv7w
/+wiGk+wnvKPj4C4wXDUA3ajMpJQSoxhrucxdBULKChyv2GNUX1w0d/0IGCAaXCV
V2er8HmkzapbM5eYlnyszUjkUX0O2FjM7+DhWMSjgIRkkpLrl/Wx5HhBr6z8iWfF
Kk4pApJkB7fM0/2pDtCt4NDRN436RB43ytOdz0XwQaG3aEuJUH+2wJeB3JNr5Seb
BJB/3e2ziJO358uNm3cC2XabFtKQ7HhcKHo1Ys9FzQyR85+PgwbJ0TcwafXtPAzb
vjdGa4Vc0P0JCQsyGfXWaSiV9cQDes6nlljiyTZYHQCkmPqc71tM7rArX8thKzxJ
5/36htzc5PAluVYO2jbwb//yAeqgXxymn1kXrmtV5KO8fjzILhvy5IolfdAjQOGX
QPbbJ0B1jvdXekDXUE8/KeuCZJVpDcZO0uOQusS9pwv4x+Y9FeMdaB5bqZxtU5NR
tTUuZGZ0mTyglQ+35w2BJyahpiKRPrejOSlzqZY8PkmkvSLe+bFt1j8KCtuqx+TR
x78MbJsW4DyNq4cIae7tMf1NMMF7swFUymoGdvPnTK42eUfpYLIrwC0NSekx4oWD
0bWpLRPneVvCyAq6tHXAh3upfIdwu5x+MobiswJ/vhHyVx7bRU5bCqHH7Etf1Gh7
xal6omFWOj2LlxRddSFJ6XlIcelbv9q+nZTokHHu/Q9nS3UrwxQR9O+YLplvFHQy
jWJd1rpKk/S+M0pw4X2dPdjO8nlPRh3VtQh994BXm0CwHRjegkSd1jXa7XG+6Rrw
hQhbSMyRcm3oM83jmVeo/KV3O6SCLybUe1/OzFEbzaQ8W4mXF5vYIxvB9Pn7sz9D
xswJnEwmUnoEMasPtwdyKjd3jWL48lfLdjZA2q/J0XuHBi1BYThrBrHS99LKKY5t
Q2461U7j8gDSMMofyhhNpDpeokH93bPMmfwDN1EE3j15b9eh0yv0rOICxGB7xp2T
c3yaFJdNSCAiIulxZCLPDcU9UOkVHip84B3xB3k/zcY5L1I6p/hmgNKO7+C6P8r0
I6psVi0UaZajItt2LF18C3fzWcoy1y8q8m2jlizswBWVnaZbbj05ydr1VGJ+J20Q
0eZrd9tbEU1XLyoxpDGUILjpvJNtR110pjln9NM/PrNIecslgh7CzsBzvYcFPUia
Sl/FMUmrQV2Bt6Ctjipo4vBKgKYjMi40RkOJY6BIVYFlXyCWAxvHG0thcOTFb9v4
WOfsWYo5vCAH4ysesrSBwxIkPJHpMOjvvNBnG5mFrNkXxGhM/9az9fwGGxr+oPbr
3DseZXGLVhFG220JCc9e/WKDTnHnPiX7FIQTIOAsTlAwb5HWtDYxtJwPJSs2mIP4
WOkwsJ3lFl6Ib7qsfd353p9ABT4wlHkLOhYNHkxOwA92MkvLBey13/QT0PIwfNss
y8FwCxCROb/ap8BjpufKnis1tnitYyLdd2WlvVRnYxWtXXdDnjHVC5GR9fAozTlZ
MFNbhcqRYXXjMg4B7UFbXgTNH9/yd8hZrHG+DZDeOQXtAYGmP5gMbRe1s/fQerlF
HtkE4gY+J+FdvG5DzsIzzIFmlUSW1yVwrdQp46AJhKw8Y9qDnoQQpiSVusGrdIei
SbJlDvnhNMibKfoeFvu0fhTT3tSIHl1d7ZKNnnFHoVi8atyxDEHaKTTKNLGFrUhB
5lR/Jj0qE7Wa/p+xxLsGqQvfZls/i+9M7EL9zfSftmKwamhDFiQyGTTxtO9SqKzh
gXzYqYXMCjeubliyTuYP4UO7DVU9cYbaTilTtahrkcSz7pRfkZovT4Z1QNopDiaA
BHiTkK5ltSWjpCCEK+SgKVFU+1bkFuwOz08lPnYESgShcOf2Ug8C48lyXEybn3ax
N/Fgj8qffoQmpm3d+ZCZKD2X6lZ75GzgMuAAQmvC65DT6Fp0CO3RwogCuYT6XxDi
QlOlvZIE7aNDmkurKt3MLC0AB30OPG1FQ+Vshof1rFSrEm8tHb5MC9UO6vVf3+ok
0YwcW6C2KcJwALRG1aI7LcGpnQ2CdL/IH6A9NBePygWnGVliqlviUgMFntwleXZ3
8QKRsydWFfO0pSlCih3bDUZLK5fm+VKUp0GV4rAAqNI9nsC3L9rb9TNsBt+FLPmn
6ndSP8NdIVs0mzWGqtH6rHFf+3qHRRhWJYwPkIR6Rg3ih60CZIf0L/a1c2ibC8pM
9y++SKx5ZwF1bJpYvBWI5PPbc/2gw6z5Q1YDRKHPvLaWzymh2Tjt0x/JCnHjGhBh
9jYYPrM3RG+7F2r6qdvED8AEdCUeK2r97Ah/e5DMmz4WctExMsXQEqzm5/n90zlg
+Nc00hubyRJ1VnGkpbGmM9bhlkr2Ndpu1yBglUfsIqqbtz1sQ60RhY1ScsSJRVsj
stRr+nVVw+2uPKmVr5RxmTBVi5S96M2Ta8SsOGPYur5cNCMBzjr7TOPlgNpnxotx
+enmw9eT1yzPZSruweYTrQQzbQqfrbWna78x7wctOqQJfimLPjxeNq7LDvZr3XEu
nFDKpbqE9awHxa2FsmGlJJWENNt1QQmfsLq1WIAVHbsQjK0DrbbuocG7b9iLfKR5
wKwlaqqTNfMXTQ58kjowMKMWIehhj7G23Jr0rEUtOHTnTTroYSPjDKA+KlID1KtA
0SV+1eA3FjXxet62O+mVeVgyhCH9EnOvrWYeHr3AySU+mmiClhmcIAZUjZqr99Mf
XBjKicaUzPHqidDI+5uMnjUXTObhC+JQN6HoLrFRd9OCXxf5aRlX4rZ14PoUBpHg
IYQKqVutRQEZICUj5+vO6jzhtBISNnsUe8Smn3Wyzwsh+Wutlze+XSKtULgaL1Fb
QAZG0oNVLeG1AFVqqsk9ETf2GRV7QyNqWjzvuAnXdPiLudEtArOepa9rhS/eAOyK
LNWGZGkjLkV1KXcJhf/4+9RSOKrv7Fxy5n9AIzVNkc9UDgreg4RJNN4am9lULhWV
Jft5MJ9pWjOyEPLYDjIF9XpvOh87S17sBnDgcw3CyvaAQuXzP9gicmJZ7s2CNiNU
eKBUNwTsU7xKpUNvLIh4A2PpYtnFSRUL7q1LY668nY189NyZGVFu7FsDqhUySM5Z
KhXUoBIbYNZZP4ls4u7s5djlsLxlEFmyL0o4jUKGWPgcVXf/8QMSEUMWGRIBdJ0/
WIvuh1xh6mns7jQBIQCqt0A8sSIZjgBlxzC7ukxOxP8sC0CXlv6KYgF0Kfc6J7n2
zAu3HW0typR9eAy6vqTH8UWnf+HjItk65wOfce03rfHF8iKE77jxhLNtbhviOMvD
NLx1byQ3FfuNHbY6Jf3XIwgZJLNIasFv/uHNnih630P0JJLWcSZ013qrIfNIoK0P
6QyE+Sn2n4L2pYYYkpDayS0nv2sZNYqYqqKGfK8rTHtCdh70/Ryxce+3qXFAnGRR
36us96E6ZD31M9CIbq/Gv5t9rNkIll0xMukmW4+uA4MFk0tqCY4bLhOA/q55e7Lo
UYaZeN82T64kz1eis5vy43HIZDcf4gWL6o3reR6/3BcdnjdHNaIeZRx6aMoEOKd5
T4zMMNsQG1ySTWNBA/0wlMUkpz95EkMgcuRjmCCBcP6ttvVLTy9SJZDezmd3QicH
7W2smpRjTE0iNUSIP5bfUrGPB9PcfKeSzvNU24Fev+WB/9psWNbN7JYYfDfC7vpS
1PQfY3lsF84Py8b9uTy5YfbOPKW6yIaX03qp0FnTMgpFi8yNPBao75pLNOzBYE1s
33TNfiZIHuuXZRa83fYPkuUWXwdpaastdzD3WyYzH/uBcYE6IbqgzrEVfxJTXK2N
qe2drXJt96RCij7IGlsIVb/+r0pZoBGdd5R2VRwSXcauAuX70eHAbekKSsNUxFOu
uH5zVfZbV9WXv83NvU+rSvqPJc1ln/ASR/8TPSFnkqme6n0GJlGw7rYUBjNv6R/b
G5ezIzikacRIKoPJiTmPMxIeqbekTDIPooz2fsC5QLKIVhaCjvPyZHg66M8C+79T
S/RJYf9ma7TtAqgVQfJ/2gZ+RjBL1Dfrbl1n7DxPDAUOvY3GvlYvo6iplpe9yvd3
s+FFu3u75osOgLSFBQq667QVREERcuciYVjn2cSM8/GGkmiIRuiZVO40S4KY75FV
0uo8zEXJlEG66ZIXCPsg8XrCSh2nIod1KuYF4J+Sz4t634TGifZpOb+qEjHoRyxJ
Y8CkdM1T0+tHIev1ots0w82U55NJjh+Y0i48YRDqCyW9hkfcM3l5yGmbsrnkTy1r
Jkyy3BgEjImJgxUtNDEdmetrfpB2SA+LZOyBs6XJEBB+i231S1HvKzn/g1TvJtQu
n4TtS1zQmKyLLK0n7J8Hk0lUEo5vlS2okYiO9cMRD3jr0gWVi7x1vd+GmAgHKEsb
P7vTLbBbbwsgbrT1QnSvYq8RT2xHM905g0b8+ETxli+/4ombY/+I4l+3f3uXG2Nm
x6fSi0sbj1zqkkP9HzwDvDS5ti0a8bRqbSlqb48CwLiwCwoYn/5ERgd2Ow9yMrLo
enZBjF62T+Y2z76dqD9X0U4I19iisqjrJN2jkHSIXofkXdXdqPw1N5PK3fmOqIiT
gTvTt0taSkEiDI2f7po68+6jHVy9Zwee9MkMUOE8hy59SVp8SoxnCDDG8fdLX+0u
YzfR6Rvn4lUoLyUzH3x6UPuQ7Uw5OtWRDu6GZ9eCyk262c3u7bCM5Fs0uchN4Uj7
7bVlrj9bp3W4Hur9a86Q3f2bk2BwQZzhFkmcwueeveUZRuNfkO9lF5R1aPJRH1Oz
K/1YExqXaqPIN5KKauGN0mUGHpGf91WfkPDaRNecSHXV4TWKDu4HNz2JiQ+W//0w
Xa+ZgSFxozboq9x/LR7b6vyF0aujif04yJ/5LQbeOkpCNnZcgVSxJ2tvTckUE1QI
qwCyK2CLnQ3apXdLlzVZyTGw5HVwiC5FUyxCOFWDoBQoNgtbfgFeR9Rbv7wvpxiI
hKqF36EzygQMxReNRISgy52FZjhScYMMbvH1IoPNGcP+log6fq5ieyvzjS+TcwlY
xIdF72IKgl5rPcHPOVKsO4AWXH4Qn+NBMxOY1yC3ZipSvGMVqHdswfgruac44BN4
tTSA5qxNnvgU4ahlubj1rUqVBfoVKK23ICXfRJjXNLAic5YjwtG1JeaJDU0Oy1Ti
w7rJ1mCYUqMWUyljOiCyvGZL+gRW3ReLDmotR/tgORniN9y/WE2BER3H/hJn3AZj
KbHR4Xhq3+kF5auC+9k6EccGT1+ai6loFTKnyWykNa6Db3Jpism2Z01le8b7P73L
tZ1ayzoWI+7RoaQnlj7nEd6aC/33TjsYT80BaEFO70+e+EqyawK6z+5jkBPPYT5F
JGQnKv7BlRJHHJGa3ndp21hs4BR56CEL9uyyM3HWKs3aA1aALyrlwILQGdLIRzYl
2LdnjsqSJZcZD1riD/A610NJX1alS3pTHMTQiCHDSA636rDaK1jxG08Zf/XYM2+r
3V32NJ421Pmk4JO1FkWFQeMA4RjPtJ2K8F8xS8HaOQTaf0aSZtSxZKfK6U5xo2Ba
zzDrupKk+CelBitnNjVMOlYHvbtKHOOm75KCq76apG7g7vfddzKhAgvOpNy9mmA+
n+ciBqINqHG1ar5JcEWIE1WuE3IbhU3q/ygwwXPr57yxl/bcWR8TgcZAPvgYfdyU
6eER0pLU9KllatYCoOPwiqvXXs7et+ox3uCLDLoMnrrSsvnkr3O0c3wTPVcdCwAM
m5qX7Xppxs7v7yd8yuVP9e12PNjf0WvmOvKGSAL3//Iqz72ziviNITFiFDRABAa2
MnHWNSzlFzc6ZInr0KSXrf9STNJnCX5G2fKjE3w4o+kvTGOUTQ3CsDFvB/Ok3/U0
MiDSB6q9NRKtfmy1hvgR0OrRTvjhte11QIlqQV7GUEyfvuAvniZJfaRVuyOupaWV
Iy8P9ebC2qIYfpQZsbVC4f1XZoGVpp7idS/lc74+i9MDANYlwrU7GIK8KZbNtT3E
tzcM7N99iQ0hOzaFmJoF/xb/QlOAoAmuxbvzCUuiLKPsja2HdCYdnpAEY35/npNa
CTRp9JTxG2ocTjZDeu23V1Kv3iKoewez5yqQ5PLSp4kL1nNJ0Uqi8GTW9WxOJ+on
azX7ujzfdJsz2sMHJGCmp+b2n3D+ZhgVaNhT6YILPdCtmjrtW6LjCK1oDnY8bW92
nw0Q9q3NSS0mBNo2l5i7QDBd09m+3FR7IViWOaN9DdH42Jcc6HiqXD2/Cq3DFz6t
sdHtfm4d9VXRDd/njCXTyKTV9dRQzYPvTFaIyqC3Ynm5aBPAQ4Baq2vqLTE0TFch
PodKpJxFWZtWbPp+kavTc6rHsxmmfc8+Y8/b0lDKuiAinyCI7gND36CyCE6FgR+d
JmtMvW/bUe2eH3FTuurOO7ukfjshsOFLKm1Lf4qo0avdzkyAivRZIuJvcwG2Vviw
3J5SFDThklaxt5YVuZEO+3qE2NztcYbr8Q5XHDWYqUAlW2eckAp4Mq8z5qQ6fDcu
CdSo/Oue7cMCi4cMCFjr5gPEzQnh3Me9g+F9Ry0aZN1ySiieMjOx8DMfAuvRc0iE
7KAK+Ippu7eiskVm/rr+7hD+OOItfAsuEejq/kjl7w3+VOylifmcJbdCi2ZAR2Pb
vMofyd8Sz0pcumStzYf5137BdiF5ILvSOGb36pST49u3BuehFbnbr2NT0oB67uFV
PtR6XfP37RjjQ26NHyliinnbxfbsTV5zCpoEMaazHzNgoiB7051gQ2bBrtJd7d16
oSlUQq1xptcpGSDSxL2dD2dhVOQzfdrhu0aJa/zYejOXXqh7GFcJeA4ZXZq/qRof
eoQE9ebKrMQNC4AHtIV6gKEo8Uh6ZPu5ebyY80M4/Kaj0NhgmoRGJQmG9BuwR9Fi
6qNyjnD5bjW4AqZEh91p11eXeLTw8Ed4Bmi1Znld229ZDRIg1hk2iY4X3wktLv7b
IpEnGRzFA949SlKNj/ZiRuSfKIrc2G5QVgbPEUaGVsC5dUuFL0dhLqqftKhq/DC+
Xy02GECTFMcW1CbwFb8UbhST4Mydrlq98RCL0hyTQEyULhSM29ldJBKAh1TYTtz7
KWUsxxfnpR6G54GVJ6VIS5x1ixJkEk9pyJStcQbDWWR6vYH7MCf8a9tuYWZFykwS
yLM2B4O8GT1+aKKvH8meeR76zWjcsG001d21FC/oGnyK6kc97HLkzstQ755LsfSW
lySE25rXiCB/6uKSY316VzIrMZXu1tUU3ElfPtOX5Ei3t9KXFf0kBXBJaSkh7pIJ
QXVPpwiA8JrXOexqQM6m9tp5r/tnzVgmJ+GNeS8IutLy7fTfmljPRVVuEmnEZe/0
PcnEITrWNkPdv85bO3IeJwb96Ekf2EdaUp2aIn5T3W1o1Kgi1L07EnnfexbRQioy
3CsPl5XAWRzb0t9OQ9N0GjlZqRGPOxKVdSzkFDypmwxfhk5weC1Xwp4QJ5jr5AGo
Dm7ZM4DC0AG6BwgPs8mJrYKCttxpdsfOtEdmirzIKR7U8RbsfxujabuvLo8e6/py
LbRtAWJgdMsPFA6cWNa/HLXJuRwKPGz7T9q/yE7iPF16+PLWnhP6N17fMiMBrpwM
M+Bw2BXdNg5k9QoGKQWKJbo2BW4mgxoP3SUgBUYDJASc+e110wBq5GD1cWG2lDtj
OS2xedPn7HbDJzCutVZcIvwP1JPZsKlptYSGbj5wXiHe8KlDb6Y6l9CedMo4JBPf
zbJEw1/7OLagv7taTZbk6dfceC28MHFHr8kXAFS6cjPSnh5s7zQeOJt7Fb9sRAw+
UUdX3RGs6a+MY2n9vcFXKZTIR0LQHkRFR3FxbuTGsEr4yFu4ak8v4led+nxUNZQE
a+xX3s+UtGF7SpAiiqZJdqpO68Gr3OLHbqSCP2/q+8xRpQ7nflTNDUpSCL6xV1y4
2CasKSR/O5Muypm1EwcrdCZxMXZW3yiTGKbAl+wh/7OFMn6v5/jellwCzSLOZsEC
bao08zUD0x7FtKbdgejR5ZhfHfrVXaqHjPNb7pt4+XyV24A+XbEy1BFIDn3sPD+E
EWKBQ5DYdxFJl4m+iRNhB8Qig6ghSanDZwnm1E0nVpki76cus3VOtRnno2a1TCNi
4bKk4CljnDYIaszoox1C4cqPzHlR1LSU1/IznhHz7saLue6z73bM+0CBrKMBcwe2
8ig5h7H2eUn21cqzvZS4hOZJYHipwfbA0xWM8vGhzSIVM8KJn07TBXtO2pWM2Wko
eo4t6Vwxz6RwQGVTPzxgooarwZ7wLneVBP8YiETWlVnIFIUcBNkmElKnp/+vU2iO
UHAYAc+ccjMQbblZhO+MY9p5oRuxbArXckgtBpMcKpzyjlAoAQiiDIIqtZiqOcK1
oiJ5VG7X9TJPZyli3ZewT+1uBgKThthaQqB2suVk5mTWrZLiMQYZrIDMUCMBH/Y/
981pFIvEG0Poq/DQevb8iALAiYcAyP8M1CnIS87X92fPYUkEtJP8BIAXN8VpwYMO
p682H8D7+d5m4hTHskjzJYm41xxAIofIYkp3dUCeTp5Out9n+VvHFvpxFuthYOw+
S8up6fnjS3d6Xp0J+3xg2ZcsNOEc3s0ZsNeJkzolbaTIgD6amoxnrgO36LJ5NNJ6
qJB00UFfO1ZCg4UPopu1UV9tPmHAMaTa27rffKboShb28AAC+kVSwWGPKmG9kInu
GLa/kD8PwUXAxOyalVD0fHKVUkT6V6pqhgTj1O76GD2linCna8AVZ+oDjEOoYkSU
MrECfdmUPHKV1YBJzgb/isFr0DWO5p41MYqqhmpdcPk8iZZnG9hZDDAjjGGB648h
aYNi3dqXIAVFwPxdhuwZVtqWOw+zDMQte01ZD001zlqVZ1Rkjd/DTHpR0xuknLSw
wZUa03BZ33QWlZp541PLYsxcwWWAIAIooCMuFzbBJNAzaj8wmkgTN4FbEoVuYTEq
vMAjpp/mKwtVCDcuBG4pyLc+MSw14kLJx2IAnEnPgh4EnucGFEPFNinSHovOcknk
EQ3KPkhvGoFAKZkqSGWGY/2oryAsf9P0IL6uiY2bam0EZZssMn77zGJ+RblHpGwA
4pDeijH7jJEv0KQMHjOErpDtucfCfTExqad9j2EHmFQsw9Y8GVYp2fR/RsG0abJ6
4qk8ynvd4EKjw9JRUPQuKyfnxUY4su4YJI+1LRdHubTlogSDqmfRWIwBoVNdQfif
CdbipXESTw9hR1U1Ptj18MMdw1y4WfNXd6XlVTAnv9acPs9UTCsGjBgHmgfUQ1yF
N1iFv/aoY27qzJa5y8n0CRIaafbRiZ04krh3ft7+qPu9kwBX8LDshRFp/E90ofPC
tq/TQW3bP9BmFAzxgA3Ba9uKzI4KxGzXE1PAyWK5vVY2Ek/ve3if4jtO5IXFNj/d
etqTUah0/veBEYN8OEdD65NYdUPpEGOkf0T1wPldN/km/T/MGl9Lh52dww3ieVcO
YbSOkTLWgtzGgN4Pk5kRsHbdZ49duWceY0lwMZTSgNM49r4NqDV7Lf4SipFOKFeL
bEBiQ4x0++8l05iFaEUpcHq3F7aMHFhLeaPWfwZhX1Q4yI8jTWEoMUrf8ZuPJ3cW
GcwIbwzWtGaEYntVNtua7EaqmULXVqE2gztlkDz6BI8oei6yGz2eBtmUccpHlkt6
qDSHjLa9OUQOSmwdmoCIhCzCtK42vycPkj6kyCP4rf3jMZ3kHx4M5P/41wGA5Knp
D/rAp4vHCWLCSxCJ+153dNlul0XeZmc5sYVba9cehnQ/x3AaMBVn4fb4AcRVijFe
mjnUnhh72DT0jNxE4caZPk6yGUE9W4zizRm5bB1kyBnb2YxaFU90b+brImbwgs2V
CIrU+eYeFupUgNFOouulFEXmElOX4+LLx8ujtyrF11fEF4OsM8c+onOjmyx77/U1
GuPcRIDFWy3WyCbe7izUY86zRilSm2E7KbDx7Ud0YXYGOV+T4RpPEVyulCRKnc87
TEJn7UNnQgCqtrhWWCDIbtCF9/VSpmn/Au+ETQo8wT3LXqa44UQ95BPlSWRNnAF4
So7QCuiiAr881KebmoCSHNI5fPlozzHu8t+RuDOoYezSLOAk33QqEpMH9m5dSBPS
IVzWZF96rBZ27jsfbYN+Ft6NEjFg0kzgToIls1r9xpubwkV1RAjuYBiUOgtUY9LD
bvtVUT12fAd0fAaH6da/M/0AA1BNblZk7Ruto34NA+enpW8+/0vUsoUD9HsWALzk
jmf4EfJUJ08GqjqxzynfLUGKQGZZqAJDd2XfrVqxi/WQIlDmT08/8wvHk2Amz7Q4
aRQuIDMxNg56oLGCfHPZoqtP7RrdiC5JFYflZhOEuM3pdJaJ0IRPlupVKl72Av5c
QYBurR7PlPegrwL1/ajaX42oDCeIR3fcLPhpQzkgdWcu9AQxevRg4HWuw0NLlASg
wQIZF0HZWaywvNs8E3jjFr489ISDbCAorILQXkjyVAmNjwRkNn/HKQBCjV3A0bg+
Hd1J/zo2afAtCAnpdECDDGMKSQzLezkkGjGKmOzBpmgYuix7DG2bo6Vagf2F4iEq
RCFaZBNxkqsbAh1iAzAYimYNurVTr/lF5hKdV/qqW7w7VJOZtr0nJ6d+BpYOhmHr
fbOOgOgLXeRRjkQNV2t8fJErX8MMU/SAGpcOyPnQEd5reHxYspjbG29HIGDJ723K
A6Qdk/5D4O1DeOQr24zkrROl4HRAI2cnHO9bWBfxlaJFNYSS/O27UGrB+zwZt0tm
suM4bWnjrjjx4xZpgar0EU3tLO5BBQn8r2fEBm2mWV8lekQIdHZNqZBNBHXum+tg
odAzNybKvdgLTRRy82fx6BsAM3tei8712YW4aB7tY3PdObKx8GjIxRi2niju+u2c
sMrG7hnfJq+9K/Pcq49PjfHRPkeOFLfGvrb2eH0JcJOGNrPk5tiO01JM/nI9BbRY
gix4fo1A4NCe7/kPTodPAVPJ+ZGFxKq93iS/cuxbXTU0qUo/9/uw3LU0St/PtOqv
SL97eiHctlCz4INKLFf/96f7JwnUUEfKYaIotIKH/GkDfEg5RdWEjC/slIYWZ9PQ
ToIVQ2U8Vdp+ZEjME1lmyBcRAH04ZJJzDmazmjB5dro/9WKZeMY+SMDEzPuoNrZc
ioz2aU8SlZfEBCXsEBeNCFV0Qwv6QloXlGFuHCt819C1QkWU1xFwgiqEX+N06b4g
HRqNW3gQ4cBNw/GJkNWfsIEO8gqGBSj5d4axBnJ6vfpwN+7+DAKLW8+vQ1mApJin
tXuE+ZviGjvGBO7X7a+w8PxCtB6RosoPOgIkRO15cRlkoTLIB3ZcIZ3VKyegWe4s
Zh6JXhaHl2sGGl5uyBHjxg0cyuzb7b/rsOfx0GrHwnPjx1v/TSPsCnvgInLxaa7y
rT5qe0S4NbznArE+6weUg/XGUdWtyexmxglLCvuJ6yvMIP6aYITR2qv4iw9XQTpn
PKvZY5psIHSJhDWGtHnr5trczSYeuXN0U+p4u0NMOKr7egRb3XcHa6Iv7fr+4LNj
ibJCcyqBU5HN6NbBtRlMStgXGT0hIpdQN6AkINofg/ymkyK27K3gP8tPrdck+HIE
AUM/A7XdZjwVk0+xWdXk+jctiJ005q6PzSi54DMQa+6sAvKcDbwEnmfjpoay2f+5
d+BgEo52g0hGYTuc9TWo7K6nUOYfH4ax/nHzI8QDEKKg7K+2Kq3Lwo0yIvDE9Zbu
DkOxUORQmKxb28gLZr0jGqAXUTQveYUKjusEXN1gr42DfnxodkPvtQgG27nRVX7X
TIme3T3zMaN4yxDtp39sN9GxGw6vWg0tHLJh8iRIdk1+SFdI1cqm9hfuJpdAB5xZ
+WuaZ6gP/ntD26qXBsj7vNvQlZzs1qGZ9KnMcZVfULxMdl/hpPUCpBUdUL9B7VPu
oe8MaxwbPTu/HgMKv41dpUA5MfVB4sAIoisNaRAKAgrPxkzW5Efuh5eMz1mccObg
fCku6VpIyE5+MT8Cc9ucbYex5N8qwK3xP8zdBV4+cHnK3V94RzRuRkpyEE+WEKUd
hX9eD9EKOPEuwpUb00SUr/gPiKcVPCwDf+ZWkk+QnvXgwzb4gpz9xuy+/4GJ3Ybx
VA68rDGgRVEmMxtNkroceqgKY9r5jdL7GqSJw9AdNi2rHIqImL34Q3TVTC26lQh+
MUwtpPTwYxHxS9F6+Ft0rHbPVOPbv8F/eJgVnBv8GeNpk0gICXYYYfyfOudd+1Nt
3MZ7FuanrgiYE6rpQyc2QrO8QD4JJUGDvXFE1NAIyPD51/yxOm3iLFdicZwK32gy
YHsdFOKnijKPOeKJfMHnFID+IwxLshHQ71s34VUhLmYovmQDb5fnMp8QeHny6KUw
73vP/n1M9BX52cTr/LnWvB/YNEun4/OCvKbxzrXOnfYN03rDLjj/m833X1iDufWE
0AIWX7ks36qec8NH+Ky0Mo+/kca6puhkx7O+9LkFU1hvyneDMq2XzZYJgNvXH4n8
RY+O4uWiSaymsz2sxikD+ICI+YHyxORdfH9whdW5B6YiuIRn+2H6Uy11GtgUBgLz
lOZ8rtdO2U3kpAPLbC+CzN8Gs/FJkgln7G0KyPW+NuJY4fb6Inf6N5wd0L7e1ZDd
G52UfClMBaa1ckh90DapR4IDyubfRcmm9yDZfRlhXo9sWPjph6UZ58wWUzQzjwNO
6sHPxKCRDqlAVlWwIFqM/FIfaRugthWh239gxnu1do3Z3uBPFwJkvXsxfMLKzYl9
/CVDtfkc+Z+F7ZNXrsOqbiTnD4hNXT9kc5icY21nlg9DMahmOW2C0+sDgx9I4pMm
tHen32R4MHOe3tQvazfjeYIhkCQP7AD6e/nghLtPo+TQr6OtODJ2I9YAFHgm9yWQ
TJorfgHk++rgyp63e6cJbdpKVlbVGqf80LcFIv8A1xNdeba1Uh/OIkAqf5Cox7+k
g/sUb6TfyjNtXfAoKcYjdyxhWfNDBsm7lnMHl/zoSlrDKXNesKsM9geNov3aHh0V
QB0Apf+bB60saYw0vUrItKq2AmjOXNQFvrQ6kIU/xjI1ShakBg8U7/27OKYZbKv8
kXsF/Zb95mNYdDgHW921aW86UNHixQ/GMSc0RY+c6EEMnR3ld7pv0TNNRQod2uhT
37Vgy9LFQNuDTLvocKYYyGC15cPRYL2vztGe9bVg2LzGcoW/HrW9NaQTet6kOArv
ex+P1zYhr2Onz9PIOoy0aEFkM2hffkiweox4PIXqdc5WJh7Mm7wpH2ryX0y73dvi
YrEe8tEXtORjO25RUYzzl5WfgqS46kzC2BcOnZ5zFxc6gzjeovs5V9UvJFhMD6IV
r5JkdMb09uzJ2fAmaFgZ6n3Quz10hPshSzLO5Udz8YdrUMG1uvqVouhbzlyTGPcn
1TR1N4KaXgBHCJGFolE98mBXBl7nJqYxPvt5cvQ0kzmXVBLOxpSQcVA61MLcaxvP
C7+kNc5cml0SKLBrfnONPxsFFhDZhBd18zlSjh/LgXyFU6diEe5EFgLmOwxCAFS4
mtCCQ7Eezm6b0P72y+aksYYKOvniHLYkAnWoHorKzHFiIlZqN1lpKkTv1H08Peeh
kjBkAlN+PSKII9HgWEuCdG/TvYn5Dfp0pRERPmHpda8kf9h8/ybD4gtHDYX7nDyx
VNSMAdEtKH7ft3Dg1F0v9q8fPrz83t/exC+XzZBw8rX34rc3gYq33MY7S4ADp9EU
+fzpuH/ECEKL+Tv+WCR4tG1E7By426/O2izv7u1cCETwQLG2guV4DDENL0kusEIx
TYHPPu3Q69qRVipKbtKegCKDNpdTCGXhjqtUemRxiUeNnGHUgxz1pdQzyBWT85+v
QUCyewpDth/+CGn8YMe39Nw4yPEZdX1vYdlCHj5E9e3Op8D0ls9VJIMq7JWpPwG1
wT06Hu2qv7bNYSt/3vhVy1XaxQjq1qqh+2v30IGv69dqAau77wi59qeHmNroxuRh
ZEFHlkwb7tj/6hWczgl5u/Z6lhUhFUIg9vR7wQg2gCmT5C4yRjvoim+TdVN/hamj
Uit3TQfb/OjQ+NQ0qQuVe0AG+njtGzW1VNISr/Tm5orQuwQznw4i185GqDY1FyJp
W5gAtPXo0EFtlVLKYQ4jLpDpSIwQ7Oi7QU465j3F8tOnRB71PwqLrjRPRdoV0c+q
h0aY99xa2br4RH+gGbhge9OSiz+NYAcc42ANIrvtFEtHJ1lft31Sqfbqb1InhUCO
c3TpXuQnPpvGDPvYdCxMHWNStEKCTNrNVOcO2dRjlkvtUhLLyDsG7Cox0BwZ9BSV
mmDGvB2uedYECYr+QlSlcCz6tFe2rAIZhO5FHOe1+i8t2F26Peeu/8zwd0e60QdU
lYxRhJxiZyo4a3C3GWcvEI/hY3fFV6nahKXjjfJKE036Vf0/maVsDUsBiN8LugdX
e89JwyLP2hyIOXnW+RPeis2YPYBY+qGW4lIdbAWYM+mHBpK/Z3B8DhEqHCfvN+MV
Pt8DNNv5Ce1WnHjIBVtioFTTpLqGRhfr9UUeow/Ty1zQSeWFy2Ra/pCbCg/zQrI4
hDkiuy8GeTbh+ihX1sCYqCE+EH4MDSIzAlpeqTFh3Fi9Y7xJm7ciGU9oTjQpslfv
Pt/eYYpXPqTGDQzTiyWTxHZxMxuFsvGaLufZYyOaJKbYrMnPVJLvS4uCpxGH15aj
ie2ytMyWTylUzmhgrPk0XMIrLyv35d/gnqxBgXC12I4y1FPOeysMdEABl+lpA8hL
dJQWCck5pNE0EYgxMa40wYAPgS135YGAvjDaIEHZushld3Qa6iLN04cVHU7IzJY9
pZeTW6OC3ZMCSSNBhY7Xffi9nER2X+jMp3MRkiJk/4syYJ4Kfb2mlHIO0s/mffCs
d0jhhVCqnQrzfzo54wj/ygnwgvOli2patqrLWq5QnsUqGMe0mpj8bHBipM4QYJZQ
mn21QL/t8t8laht6yW0g9Y/RiGEGAHJ/7g/N183XZhJR/bYOfZpvVxsqJaO6a3St
nnlfBIkIyvhblNxcYIldPa7/2KkBXTqn/4VXsdvjtYFuPR1TwQss2uuT4Vbk33vy
YM1lJ2na2sANOc8jfiEtz3kvcnr/W1zaUauGKV0Bpd9tHU5i31x/TBWyjydruzqh
Fsi9LeDCHh5U0hSxPGZ9b+GJsdYMicvDvyjQuIB4QrAY5XkmV6A3UhcQGCfFWvBy
5RNg/AzivQ1FHt6su1VpmPVzs3PhUp3954mcqqCmno0rZHcmJJ1/Pl8cBDnFtZAM
a2ssETsjTO8mn3YgqMeU352LytFvF/Uv5y1qllp85wX+byYOUiBFo3kP5kXED2RA
fUEoYVDTTkSn88CiuCSlPVo/1HdRbodETaNGufkFe48uoBS0/KeB+4XhocadMtfe
5wf8A16ojRyWDC4cq3P2Mp2grXRT9pgjDvLlnEsK+x1vMLYjwC4B7sYoa/DvBo5D
yozmxUkl7tNq8df+GvQk0Ps6SFXFSEaoczu56YG2Ff6MWscXYxQ3GDsJS8uZxkta
rB9bXSvKVvxBQspGJLtIZwU8MH3QMuESl+o3RzZ136YOaYdGd8pIyOVWfWj3LJOp
7q4YjXfvihLS4wWETnOLkugtB9HvDLusMnWxrXt+SUcaCpkOraeZg36S7RnsGCK2
FbfE8NIkqKWY+WngBKIViIMERqsXQpY4QYnGCeHGy1H/e7d9vMtu626ExwwktZpg
O87PZg/avnCFUjojJm23ACG/Su59moXpDzF6woaY0uSYpXPg/x1v2Kxq6iiMeLvk
BCoZH0hvXGY3DDqi9YvFqdyBTNcf3bTxXycz6hipnlLZ3dMpxwhnjH8kXJ/8Y67A
mE6lQP//yaMJKpq2vZ588XA5OnLuTiOTGUv1zytaWonewbuSSlmWaWoLab6gy/87
b48rur6SELISDjR3IwcjfH37MIphq/eUqD37qBDGXPR0W+bJtgUbfLZZHZlIdQB0
gsXvv+kxmxJHrOg+waV2jACJksHgLdGqL8fmlOKZkPHCiexBC4j9CRCUtj+o/IGb
C1qGFNPdEUDVeDA7Ah9m63HkgAK8BBECtQnKd3zT2RL7Dh31Kmars+gDC1NBBSoF
A0MfvbjTAK4ADD0VsVenXbZn1SdpAPEn2Qj+QaJjP2XGt6YnGBeCWRZRlwIura4D
+pywMANXObhFoGYKEzs9qwvew4n/dwdNhdXvoPRrp3ke9G7LM4VKiJaznvjpzE0i
JNAd42R56QkY8NYIxJEiZovtPEbJ6x06nOb6qb9U+ARfPOseaROUogT7pVrYj6NX
Q2nOqnmY0skG77HcQKTVE+02INmufXNJ/XcwIF1y+pZr0naJJf3UcGCUIunWnRfl
tRF+3276k2DJRcZos8zOlKm+fKquipP2snNaRYmRtGAodmlhlFGXXpSwDlBVmeVm
3AwMxS5bc7xmLpMEhbSpi6hnC3tkKnqm0dQQR2IMFrSVSNxebK6yKYxrdtUOUMuR
J3h/ZSooAYQbHrFvX6Hp4ctC5pGhJAmQ8P0vGrycY/ECH2pJZg+c0kkaAO/Wyj6M
EUqBsPtVR+hhE4raYqtuHoRXwaUSZbsOQ4AKnhpjfOdG6MFf0Emt7g1sH+k6JAna
Nrd5TmN+GFsw6d43rPgPVQWW15OlZC0svvBMIN1g1erKv1PACrOxoWbmtuVoiKKl
HxWw3hFSaR3uDV6h7sRVikZtklQnvvOwy3VTdZcZAV3gVj/OcAgQiUo03G2TC3qi
/Ddb9SuNPB9t6aqPnWxG15DEHkYfjq5XqLi1zT/0dt+9e5PI19wBFUybuSOJVYFx
iUqZPnvwQr4FtR/5Z3r826auh1PUwIK/Emfs+NBTQWwP/G/UKgnOIbbmU/z5AJ/M
vlRbmgvRE9ZdaqH5ab2lwSU5o10YTYNbdWIf9pR0rsQmnSa6DFpr7biclGCAb+at
ZcU3Fl0q2MZgxJCZHAAs2Wu73fjtc5XgjQGKvw91llgH5tfDc2myQirmqk/d6JoQ
o4ZoMGeddty71OB61QXVKK2DiJ8y+u/8e9oebaspCOqXVm4/9vY8CutDBQKRQ/9O
VUdFrNba0zBLqIz5nxm3+Zzxyk4aUmy3EJ87Ypu96JZ21fPUOYCzNnQ/0yY5kMZM
T1zkHho+S+KYklkfHb/B0YQxf5EXLugOGjekYZCgbIeQtdn+hS9S0C9mxFnAR03v
55EQPJ2S82NTHnvbeOKGXNS6cTszUeMYtj1zVbU9mM0FVATdgVQyXPWiVp92Mxb/
rkYcPmrmfClKRP8m9YXOVR/FPuimBdbZhTpFQNNsb+2DUEwK/988BDj6guZk+H48
LNwiV8KAI+vF5QLjT7mIMH0l+1WN4EOJmoxbCQnRyOWntPtXWMMl894kmHd1+emL
jbdrBmOhqNSJOlfhLu1EmjURhR3/wtCoa33JqBku52SY+vzVvWGje4jGIpVzNPgs
nww3Qen1pSC/sgK5lUO+SESSe9stAscMma0lApLvzZRsgDbsUdosI/IedOJY52mK
5NRsaRPTxghMf817RH9d7+slejCar2jr7qrJp7poVFcvcOsHD3XtUESXgr4ryWTk
nO/oS5xftKiGZ6jzDNYlYTol7wPlcQVgnS+vGkqMv32ObkqHwoW8kP/RceI/tsVY
VKChf4PpeWzG2KQenDeM2RireJ3MVn2+IIT0fzqAtyeGt9BvFfuIW+K8jgGVLMIQ
zD9x1W66uPjt+hZoKoNaUW0GCvTx7uec4JvvW1MMOJDnoxHKILn2/wIhnccLodhp
St33qEOLczzlNS+AU3M0RWxQdsm+Mqj4OMSpVBJc3CuGks90DLaOSOfLHwFm+N/2
R4lZERdy8I8YbEHwJcaBQQTbf756yRFqleqcU60XZZIrfuvo0YyK04iWd2o2TGTE
PeVz/eCrzSNrVDHkPqFJZNkyEGkqGfNgC57UGbyhhVnaByWdpA7HLbeTVNSmIEm2
dk1Wx7cd3EId72M1sdDiMPytabR6pnqydTXcexA22HYM6WwF/O0Ngg9ZpsWYJDUQ
XRt5LLae+oWivXDJFCcpmMz+84cHs9d3zMYtmi2xf1GitEB+S2QWX4jANAydEdtx
mnx6bph7I+j/n3nQpWcC8oLjexhPWRm2R97J7ie9aAYuK7rI67+C2U+FeV5+I//O
AKpM5+MPGN/w2/ebJStQKFUPJKYF/pm5uZ/upyEwdL+EMYb2I/8cLWEAgp0bWJp9
/A+1DPUt9bj/nV0G1rUz3PmIozhsDGtNtKwEQdgZmSztJbCuxCkNZ7MTDVPwYWha
lcrzQOj+xASn9CL/Z9Uawl0pTznaEBhhFGKdWR8Okhxs+7ml+5lZe1nnpZd1gZzo
WwN2cR3PlQcA+LRjF0sac2mP0hoSW3YyqA711ZSLxoJjt9awoRcT9gTyY+6Ybt7/
rwNdvkOIkX/d82DpdmtTUMcScZE5ScJsfd66NRVKiCR07zV9BoKz5gfspcHWRUcL
UfX+RvMIGV3EVVwuiD+L+q4jEZXzrl5c2Acch2ocsttViGPT/MjBtkOweKS1T3bT
wrr6hJqTpPrCQLKgpSTkojQVmi7ZpP91l/EwUSaQWDnq1BtRTKbCc942MqSgb+La
XpiKBqVvj036VNlapJvz3Hb3b8FphneOsDEgs00oxaSNpsQhtrLUTFzq3R2AIh5b
WLIN61dCMJ1TuSrPHn2LMQuQibYlvnMTKXNKLr/vi+NNAvkn8RMPOe/E32I7t7bN
uExyK+hqSXVrpDVRv+A8/znLKDlvjZzafZhKRQNYInNMsDlIbxAaWOTbjy9/zTLW
dQ2NtRk0DeOlMPgFdMls4Ur4BS7bEITAoWULxMjEsRPyPm7kMKy1QlWhZxABPz40
FzJ6rBaVtzLhNmMCP+DxSRhdycmu4sLTS2DUmNPvbbWj2K8L/1eNxu594D8WjfQZ
ZtWjxnYCR8avS9fmwJ9MqJ6ds74l7+E9C0JQlnZXJK+BL6eNxsj11PUjhpd1XKqI
+lVr+OPPlS3gKBKR/9rIoeGyv+0NZkwPmJNLJdTwN3N8hII1oqp8THS4gv82RXmv
p0Z6tteoc+VK6irfUMV7RcbWCAmbFtQZZzG9FPDAAeSaBhtdYw1gsl/FejhMh8MX
/EN5i9PsugS0j6Q1HHit71mm43XtfdYnjKrGYOjIBQCX8RxUaS8xy6K8931trka+
lw/LcipfnFUYFfGV7NoTTzXWea/FFUbVgV1tRvbk9WeYtr/tWK2/n7x8ffymeQUG
ihu9RKakI8Bk2YjKEsUFWlROH3hKaIvc6iPhuCIQmOej5UHNvg9iNs2OAqGy1+2L
sRGlvlQKbmvd9KGiEWYJ3KtoDbps3DFpQRgmXrheRGMAYCnFyqGgSl8La6wwgDGt
crvkOWuwfBa+MParQ9t5U6rZpdicVFyyflvAFSC8AB4XmWAxgJXL5DXVQ0ZIa9qv
P+B7K/xUkQ3xdSaoGcqc28admmsH1QDJ3WUG6t58bcjfb+5pXyID1f0WiqrG+ucV
yug/zxYDqkdE71F2+zEjrtdMTPhXDn6al6uC27zmZO7HZibkbcHutZh+9FoFKSCl
DjJdMdrpQNIqrj4O1cSYAt0djQsIbW/tY1iJhIBoNS2YqMNJfWq6O9xgGfWHKyWg
MZC7hxO4uekBb9t9O4rCG5qq9buNcKW5cCbgUIs7I/AYFBtc/Ob6t0YQ9SOXRLN4
2aaAJ2ngZ5F9gWR0vpv7G9fq9or2vHDtLlRH2Wn3/82OzQUF4I8I1+yhvEThg+D3
tC463paivJRxXdFSilJtngde4joTi/T1RdWzlbkwfc8H+H7xvVdm7xBEn8pQkEf2
ybHZEdyAE/f0PtBz4NPx8vcr2IeAXcNmQdzfEIRCBSItEiC1DR7iy6Mv2+qWtLFo
q5DNAljUJcpfOQQfa7M67jevH6+QvVniZAImXqx6L8wrO+6dpxWfhdtvpyaKW8MV
T9fPBLQYhnJxRnhrr0bKf6g3U0VBuy+yPt9XRqsVtTVjvqu7LBkUjzOWq1eOXaqn
J6jeUAlKCA7cgQK3MoYxfDfncs+eazEkWmwNt7kwTf7+ZjVecK8EcZ8m4WF3JU8a
Hh7oTMrfDnC3weFZPW1X3CBajUZZNBXM5hzIBtsfK0KmoV/H/MTjdHs6TWl+U/BX
FETbsd7isgZb6qcskSEtcZbuqttLczMOw5bmrCe0DLCqNRUXKfqwODHOMheR69Bc
OaSWxwhOj6RFX80YdbR46WB0HqC6DBmv9nWJ9T54JfxxKMdShRYXBis8sLZ2thnQ
UgrEUauYlZ3SObaOcj9uB16RWy1u9sUVDQPM/O56BdmdbCtStaCLbZGFe7otkAqW
CvQjAGLalkbUdx7wKcUuEzsRXL4XUzykL4Gj2hw4bQWu3vuE59nXWdgAU0RIO1rW
yBQvFThNVU9ln42JQUqwp4aOwOOQBZn0yT4QOrCL9stLx7cHbD5S8ylVEuGecmjL
YCEeHvDic2+SVb8AAoDkFHLm1RUSxorsO+z0CRSF4+IgoFDAV8gjuYK6hHgxavXl
LC/fKTaiRNMFlptB/3k+IckyZrXvmLAhkNs5l5lo070pBprepYkhrkrhZ1WVrUt1
oTxvh+lzWr4UnwcvyWKTY0JLR0XBeLIA4TXfp4JuHXLd3I533lYR9MZyTZSH36Qf
YCKzfGLLcmt4KOCqvwEpsDR9ssDyya3yJScAH1If97TPwpbcRRCtjZ/dV5c+swlw
gnby58z7tSFuO3aBirekiDxe8Zyessiq06UTbMS7MKxJ7SLTWE/pDq0LG1vmuuZJ
5OzexvyMAPvfkb6np/C+qkDBea062MweCqvM71dHF2idxMVCKMziaozJh3qK++t8
q01QVpi1MAsk+itUaGWEfXozxPbPFSgyoPaWC3jPexUH64tERRZN+PCVlhkd1WlP
H4qv8Cz0N2mcv+h7oW6o8qhUA1W4zg5URrf0KrX8FlYwTwYdVFuPDq/Q1+KeC1lo
uzFI9l0pRs3ePBHnnDuXFUWT9INSB5i3DPLWsOc89JYiri4HAjTFuH8doYi0RKE8
rTbV5StvSnABcvoaTfDD2kTik+IM8OybAZHqcVeraLMepc1Lv6sy584eXwii2ZLM
iGB1YKpP1/SMIARst8fnIk7GQ68vxT354Hwkf7KtiBJj5q/ZOMhDW1AgWVVmnax0
dr3F3GkHYXXoMPmtuKHNYSj2/Sh2lh3jZ6s+2RnFWLxaIeaceb9ke/z/QveZ6kgH
25imeEEKm1dgpIj+HhwVjaBtRX6yByhY4nL/T6t9r7P1F4vIPqIsADaB3YB5B95Y
SbamcLGvFyfnV+1rEAGYcnapg7OItsfcqHZzn6m8z6fLp7bdkdyqO2Z0ITguHQc8
bEgK72+1xeJVX9X97uAsta0kjV94HV6xt4z6ph49+tnJ8rixS0F8goahYQifxIyP
S0LQydHwHWw5p7SHY2Au6uxnYX1NSFemrDzZ2CLN7rV388RdEMcgG+mrYiOCm7le
qEWZZdtzsKAmwgIospr8R+mGy1z/gXUx6ca2qxNlp2k8BRwmojCdIavh4AjmpxW8
OBepKGnuY/c5VGikCeRiMz6rkhXnz65JGpf9zbiMsPMcd9WgfU7Yo1SAf96B4SbH
dRC/QzA1QUEAmHoCuKbG9SqGEGyvvn1R7bLGEB5LThrAQmOPZXq/cQTKhIGCA1+i
1vnzv0ylHoc+c/Awp2ZftcfPLOjYsgpv/+Kmwb5VrCkkp2orMl6Mg/U3Joa8bFj9
BvERBMH5DjHRNcprs86Gto/kzrCPr+An1rRoeT6lIMZ5dr7Vk6iJbspXE1CDfhIQ
tn96B6aYGIl+bRjo5CIdHggx/wKAn0cDVCN5JKZCJRQyoUUF1OwA4AtriwjxgFTZ
lNeopUumawYkbnDvbLZdtfWOHFC/SLhyA9lFcOVpSmCAiaEAxpUllK/hfY5ysDT/
/Hbr8hW515W6sYgQdodI3zyjMwBawgrda2Pd3eO4FAf1ldtyJK40KIsJWEPBeFFB
zRbo8qs4XmD1vVw3eUbjX4LiqDp/V+iqL0i85P/6nkDdInjrAENxAm9HUqCz5G/A
miom478CTXSWgC1urT2frYoJq9oGyQ7gbm4KFZvknQ5KvfbAkLrZkt5umRf5qv/I
tQ+nBQhZfkhF9c05Dr2YTBkwOQF9kTmdz5a5XAYF0e7xvxteT9XtZlCZXGTE5RkX
os5VcXDU7cUitHwrF8VSke7J66Mmv2ftLs6yiqmTMALzSlQ2u6JOZ4t/hvQfQvAT
PqmpYJ75f1sAWMnWh40SqHfUypyGHHen2/sTXLz4vNW5dcMwsJKzeDxD1s35motV
lUZ/h8nip7JUnYn0VradKgCIcbv2BR9S3OUsI1+rrMFfZaBWWtBHKwz11y4zPpPp
PH/mudSikhFc+Ieo4/0FOJEEAN+e7G8GghuPUaG2Th1K2/QblLUXvHZd1Y9mLIYD
kCNs8yIWdK8EOvoiJWB1KOU+J31jWnuVJpwZTRJMG8Z70ydQCFY43TAS7l+4fmpy
cxKxTrtbHrF4765dL2leE+KIbhJaTt1ehgVoepPd4cNEj5sbCbHW1C0exFGbm32y
+Lgzo8+05DqGR9r88jSLaMEQ0bf+GivYQgtS4GPznW/bZ1n7z0pEOgLkyW9OyKQF
Sj1bpWZzuH74B7wTkCN3c3E8ERkEs9tTzIkLsHocoBsyXx1qrSOBkiY5H8TxvbuI
PvYtz+x9mamD2wONHzvGAk9TPGnNnh66Y6YKOL1w5rKKpvZFsF6J+dMg+dytAZsP
jG/0vI19E4enoYz7+3WhflSanqIbNQIMaXenhDvLrtRSBWGQXFuzeWue3nKlRRm1
uKjDgkhoKSyPBQh8bA/ZIFaqXrJqra3nxxelhjaQCn+LzaDoHPP89L7rzj9wri84
8S8zJkFMtJ2tOrf5D+mgKj4MdVFE4P/ImvtUZK/WiZRogvDGkU6EpeezZ9axDdeZ
FYniIvE9fFkCd6lu5PMW2iO7HpM9Sja2vZLkZnE69BEFotwqLwsJf4+f0AbHbHzn
vuuVOgTH81jUySGnzMoAxA0r2f0pIbhXEFka89Rg4P3IPmFQ+nR8oZpARsv/QjVn
SvBRj1RHLdMtuzuNKDoM7Z76TXgmeUOb65yHbmC0ckDm//0xYHuKzi7B/unSs6Wc
gIWIsx1fF5okJPRICi5kJhfZsJzwWC0Glf4TTqrcFbsijVsuD6BeTgmXBU4pdl65
lMKEwLZ+V979UbedthHkg5LnL24sahlfAzEJgwWArxv9ygHu1QfDG0cZ+bLDnDoq
xexIFLFb8J0YWItzav5XJrga3T361RTRJPoBgQIC847x0S0Z3gEhBSsUPFwpxjPZ
qxAIetqB6JDIYXOSVW+0SmWLl5FWQF0RY1RSoddhOluGCy3YVnTbJ/5V6k1jlN9X
yfnpreCXeMHeIDE15lOL4G6OArWafdU8C8xbing2s+kmA8TjSOc1bgSs3vDHncPG
LB5EtmofrupXvIqbep6qveG6fc41enPOrcc5eODhuH2yyPlmt8m2fGc+r2k//v2J
j7LfdyuL3qgSfdX/BOu2vAEL3a2O7xvrAIl8gCwJeE7AtU/OV8PGjIXh+QQzLPzk
R/8QI7FaF/0Nhy5Y7lQOeg8tJI+6i162Zg7kuyvBUZPTGBu78SfcrlNz2iLMQFBA
ZrmfJvB0JGD1lkb8YFCcFY2TEOjDZhVqi8l7t8XPw4l47h29E8pKyj1PHw3QX145
BTd4KNnV3njhEWryeH8OF1pJS/YIbs89l6arR1E56reCJ/ltcVF/F09ISKLxDBvP
y1/KAB9r5zbKZDgUeEbTSo//PrmkCyyTic45HOxlC20T22g38vib33ynsFAF95K3
CwE/BjKODPmIhS9P5ARWdimur7jsixpQEDbenQ9c5JdpneXxH4UsUGWCdZkUr6uD
jnL0qO8EPMraevl/FmBbx4FRWh9RrJUow1rkkUNcrPX6W0p4Ui1MmNOGaXiZ3ZKK
aNTnmk3NAYQPo6gMSOxDwB/munLKRw6VjS6pA7PiV9yapgkPCHj8WtI0T04+QtB7
nVGuFNoFqp9Sk+2Pog42ZrTln579IZH8RjvLmV+B/62wo3GtdCeNMFMDiGr3zzxP
PtCCApKosCWH1EAL/DinENQzz03wFkBRSfdHZzSHTh8ku4utea0OUGpRP2cRqPit
0OIP9Uvn5+cLcS/vrgZR7Z57dU5AX1Wbbj870d10QziVnMjduvsaFzckDivP+4Z7
pnYGyZjuous2quhnSRer0pJQLpCw2XRO4PJmgd5+6z1u6hh2iSaNSs7F/7eZpe1z
JmBnT9cVLfzb1wbdAR9W7G1O7dkQOA9xni6yPTBhWvShJhEUHBIxFaf+PGITjjYm
KOT+PLeJKIM5Q6k9n6StVcd/5PBF92um/aYeNwuuQDvgxJG6lbBLg0Du5w8aDa6m
9G6HSmb/eUOAUTCHc1g4vFygUXVmdbQqZYoire7jZ5EWNWWQ1qPVGFOrmYgUhypW
0huVJ1sX1PNwplE3NMC7NlCApz3IP2nzwrR5QmrrwDkTrdx0O2kymLhquYkoGalG
sF6oPjQKlWSpC3vISfhdJTdL+FnLYdd2Id3xvQV54g1jD4w4EicGqTI6fu86UYE0
0A142MD71fs+ivZbIiZw/5RwfNWa2bJOJdYFP7UJQXAEasB+tena96NCKKVsigvy
oApxdPGO2/jivEsMm1OGyaaoMLWyotTnh6H395/aSsFN3YYrR6qN20EqrTXTG3yU
Ch1CSWEvyeWCOEbztJUWxt0sXLR8TRryK1eTsQzM3uD1ivvIrapvhPF68Foxf4dS
qW08dQFxg1l3Jiuk5gQrvpg9i9MWveA0wH0dkZ+7LANz6AbOWfTQSgg8D9qhSKdC
SfwQhcTYmcikW92255eTTLVGCSuYS5Fot1OjLaQLG8TzlRztDGDp2a8pVqzfs1gB
akXJ1wewqIrHmCz1Ygudmz+ChkG3apbprasnQy3uEHj1RZSb5fuz8DWQiBmF9896
SaHsn5FiOXDMPZrMeSF7FnEwCJ6zpC5uZs5u+hTzaSypagJVBPz8fnIfGhoquuyA
HJFuNH/kwHaMxC9vULnj7AYpqxH9EYilA5veNE0sLIzP8lKHcoXu3hEbxD1s6a68
SGeHG3co5WZan18Qav/Y8r7RGbTzGzQSjkK/omfBNfWIXC0eTbhJXjelZGwHe5uw
rIhcv7xoQb8uMADytwWYjpxKX4E7aCCEAQQdYU9hhhTRPhx7kbLU2Axpt1jkwh0a
ZeTAW9hc/X2obOTlvNzL8ogZHChrayo1u9fP6OReZHf8wdhRAEyCoGgVpTGqav/s
TfSTnhF9R3v/1BFGwcKAWrG/8lsWHJpdYJ6yRwDlqhUDOUarjZDe4q+GG9lNjDvn
9WPueOLAJ25kp4aHpaPyiWrLE4ibksqGMC/3RKpGBfn18cbWI+G2aRb3lzd2Wt9F
NUHmVj7+YI65eserus0zJE/0ypxu9uJx1eBvRYiMCKpEY+NXqGuOv37Iwkz8TMhu
xFCBkh1ZGsX2qM/NibMpKlRKEawotgoStEjk+f7+3zIYx+CmjIf66QxZ03xSx1H8
KKRHZgXFIWdYzJR0lf+6eP8+6CQ2y3jnJpdlj4FJ1YS6MtpzsbvRcMxqsd8c/5wu
dNEwUcoLAQCLoj/oQTbP3ye6FipdEI38UCaLM8smEHtf8uxVhIkLYsZy42rv6u3V
6/NP3pu3SIoO4xGqRhm8yDgWl+T3UtnbW1RZetFJ/XMeC1X8Ki/Z2rxbreF9HbqD
EjZ9I+JIT9TEOdAYI9H1IpDdwpM4KFjC83v8jofUzuoxkRCHXlpMtIezFftSrhS9
m7upDy/+lduhezD4G4nUgHaFSdBR8tgnuszXw1vIZdCeKCJpuUlrwaiq9/pThN2i
PrhMsXxBbI7VPTKqMbM19bDMgTFXoEuG/ORLiA9rHXl5NVW7HiNGD1lvNk4uAM2y
wQpmfSx9GFM6eMS//rP2jP76hW3zilcjmS8VbgYD6N8JA3apwjZ4cSDiJDCI08Nm
mV0fTbrD1NiFDnu/tIMdFOuYTZtNiud+eEgHMzMTuipkPUKVD7grLzc+u1BhYnb/
/ny13eb/KhON4z8It/8IU3hIjoX1cESlguGWN1Wc/+N2Xq8Rlr9rA1ycVQdlpn24
XNP1KB1I820dGxKPdmM1NTf42AEf8oZCPfCwl/LVwGDfSO5zpFZ6A7hg2ULNm98z
sO5f6rp0in4+uXnIFulzsAutqAj0JN6k5Rf3HZwzH0ic5yM6wDkSqSNucgK5kWlI
RAkkG8t/2U4MmKT+Z2TYK0sHOwr8jdZcUJslrHtTdIgOGIjSfMo8S02cP5XyX96h
FAnkZAR/Ayn/ydxwaonxbzn6xIuvzW/g0L9Bu1UaqEXjjVBxdapYc89p0ezZtB7j
7OXMyikpnwXUxu3hgMl9Ow7IbAf1QGaQbnG/mNXiKKGrhpHCBcaDZb8qJHEOmzFV
JNCosxTpQkKfdSto1meHcVqkGlikuiPXXqByvxgmZ6JR2LcdX+7SfZN8Oiha2Idb
DaCMbUPMTWT8pbsgGtqbfrvCd2ueRi5/TwRtb32tvtG0d0D8wbQc6LF+keY/x7GY
KiNb2LQ+Ner/5hMeTAvkxu56Ba83dHu41n0zM/DKo4Pj3CEzOPz+9CbgoH0LWY7M
LRuA5/LIh6Y1TE+BfAx3BkGSmr5BwAcJMWkG7NPzPq5NTzAn+f73JKvta05NBKH7
0BFGVbItLpw8vbylGdhmss6YOE2KeTNOZYjoBb7upaoBisnuQCBUXYl5URjhaipY
jW52fu1qWGP+D7GB8qaHjD50iLtbgYBNlOIFBN678H6+dijRiLz3hhZ9HAtLvJhV
igc/EY82gjmzv2E7OE7jbbx736TGRL9+7YRhZhj1QXKNtEEaqGf4dXV3eMaIf8dN
CDF0r7W4XL62XPG/ZTbPzVqp5a/QWCUqLb661VKh9Bt2+vBYcvf5drMR7QPdrU/C
9RT7W+ai+FNR9c2xlmQtvLPbcB45+dP2idOTLNXpfM9P/Mp6xKu3e3aBC4Dg3ZaM
oP6ui8MA/KSeZmEm50chPrNsbHXNgz8HCMmDydLv6N530rvaw/UFsGeA2Y4KAQRg
ididIYYwUXaF/hJHqN+SPWQ/EqC5QmHsqfLUGmnooM7gN/j9DkGx+3+APGGeFMlt
i9Ov62sGrdfz8zTytIxT20YhyiAvr5XHtUilbL518jy4CLHC50YFWWuOkXr5s7tA
sPQTh5qg6ooX69/9jKdSE8VeOjkiw/RMi3HvyezZ53u3BVg99IY9GJEYYHMpzxHF
LahHjsddazR1Sn0XeZooMCr5NpPZX9hGtDnFSl39VQvwiDOaoJejmC2U4JQCOnwB
pejmwZjzBNScM+i6kpju1iWVd79eElwjFXxeBw16ODPXIHBjaqHaWhG4Qd58U0nH
RlmYx2o2EZ2cr9eF9HGv1fqvzHpUjORIim3aFE7roaP0HpZk3A3RBtWSHbt5ab7q
UwxGjsv5nhDJEkycVkEhlRR805CxWcJ/3tNrqTQmHm/+c+QLa8AemrgXDRsoVSgN
dDfDc9Oyw09NqNDkWDa/EzH3fBMsYfrIjq3N5OOvdjT6k221qGuoLGA7OzSPY2/N
TQFl/5ckgZUhCIb7tEn/gT5EWleovVfoTyTteCFRY5yO/IkCScxr/H+myzGS5527
zgOGFFtLD4CpkP8VwGW1yaitqyit161kebPKFhzVr5adMlb2CjsQewW2i0N9R86g
tblllNFzTTjxDo5LM6L7Mqc4sJcftLmWwetxjtjri+27LbMiWQDCZ74sE7vCyawF
2tl1sgG6SAAxCCNiOfCFxMqOXGQBTct73ghLRBtLhOLcrxYvegRSbjYxV1xAhgrq
wL1WRboJS8+DAH5LZU39VovlEYafEtp64akwALW+Ieh8zQFKuIZITFHzaBZmaQO1
eMLd1BK42PviHcdIkQeVeJvyZqH3uYYrH9GHeyecbrV5rFEiF7CC9xdHBygm6D8g
HUt2UE6DJDfjiZfuA1/WdtEtZvpLU2KbVMFAgn70ynIg5pk3P2c0QVmoYPzGAkjQ
LupErWS9iX8cHY1Bh1zqUC6C0qe7hSkQWrFDZXzx9IdF6mDzK2uxEGH9Xe9TIe3s
v0lYAnocxMwyBCK7CUENCEnVxTTv7/p4G64L88PhElPRXMxqsyDiIrT4nJjTAHTZ
MO8sYGYier+Xi1PrlWnbWgBOxwOyKXMv9XKj80UO1qZsMtGS+ZshCTSoQUFoRANU
NOtnjr4C18TJ8BheDpkrCRVX+UF4H9ggs3SZt38PkuHC+ERzSnPwJfmxciGKbQUW
VYwWyisjklT5AkZ2kZEoCOqacFLvjWhmjEuRfJh4cwCTqvBEPR4vkNS1dxmiOONp
ZXXsSTeBQ5vecyf4j21CJca6U6KwKg0Y8IEToxx0x77v0fNRc4DFGL2EzXGlHuuB
VBc+ispgHp052V5sexrBDzHo6xMrcT3lRfS2poSMa6q1XolFb+UY2oug8Wokk72B
0p9p5SxMYJVJdKBanTRzX2tFLNUpnI4sf/e0v0MhKOcGTPKg1vg5ni4P04gRis9/
BEzdzB7ZYpaPca6WSEWVto2lMCHVjbK+622kgYx2JtW2Ky3/+KUrZQgw9Pn+y8a3
UoUdBa9+KekX8ipslT/J2h1JsUzZqpmo2rXvlcXiy/UpwG8RN/PE5PzQ9i7Tqbb2
5x8kmj/hL8EWPRnAUlf5JnEJch4Rsw10wHd/ih0EDWgtk3VmxaLPCFPdPHE9t7HX
BN79iUS7adaPB/kru8G0zfpirbzP9SGxJbhQMGtPOomG3WHydN5EUjMA0f8o8B85
4w5MfNDsCLqXdZ/+Tw69UVRLRyO0jKmn/CqLTuKR+wEuKWdqbv8jOBQYBWbswkua
z62F/i1OenkIT8nxm8mvp5KwR8paVutzaTlq5MMWDqjdu/malJGMaHuhpemEtDIk
WkO9a1F/130p/fdfqLoI/cU8ADR9s86CvUVpuq3pxBEooL5xu6fVxVVx145TkDKw
LDaDVvbHn5ZfzzNbMk+it6jnJoCoEHYY2BsWc8drtIOvbvcNolFrL1EfzCTQ2OZ3
B8zi+xmxHoxgA0/lIZ4qWCsvBitGeiHkPLiVw6gTgGgQ6p9CvVvDLsuj6X8mnakR
1DNCF0LWcC518bzIAYe/XYQhcea8d6ZCxxx1CxFU6/tKr6apck9CkbYm9fADhdPF
VcBMpHY8uC077EDOV1RVxHXJIQ7MAh/qpX/ab7xdq62aJrKDy2BigZfk9Hxy+RMY
LHqIQbOwVUhrWvVZA/R4pobs/m8AoLvjYTUr6rP2sGFNbsbOSON65YRxZ3LrSlCz
tTrBnu+XhQqrNGTrkcKpM0zhtXd50cEVWQMNjsOGGrPPcmWjyqWHhF37FZrTSwZp
PbwPM883wn9pLGCZnW+3eTlavequU34vGZ9ozXBR3B0PuDGb4g9HrnPanPP2Zt/O
rn15xLzmmM6lzp8pCm8zmsm2qrfLvPc+Ghfl0MO0EjIH7j6V3DU7lEmHvvq51pvh
U3cK+nyFsrBVvqTpGJYO5f9iOea6ukfbPtT8bgSTDoHHKOWig6v3esF1tyPXRchy
m/tO4o/l18x7piRsJn5k+DS8i90vhbxBUiF79KnKBMgoqA0NqGC2ePz9r8JLFlkm
EmKFeoTdGavJg9MVd9LTPwWnrDrAh/TQbMzWQnRXxPOuGjjq760YGRIZCgppWygp
8Zmx8p0WM6hJGojusVGWnmPIpg1l4wk0o8xX8yhQfEfP8AavlWGDteWlKOdbJU/6
w51svAs0tmtmsYZGiMTDJJ7eOQU2WHwjNKrl/hjtUmHR5ZkFVeTvwmbJ/DOGryPl
a35F2i8M4VMXI6y3cxUXW2e195CkBbQSeSsZY0ErB++COGztCWkcLRgNiDn7o0R4
62oGVwItHcXu2BYjxdsRttMgEciD2uJG31i/kG928WwteKgNvjF4OQEODYYnKAR/
Grh81bgb4NqJi+ROnwKYlJo+A3K3vaeP45m63jxQ4ukWCPTgZvjGC9r8RMEwq3Ug
Jfq1PoROkZt+WTIVBMuZutCOVc9vkEZOS6GEfyx6UhUvAgYDNuB/RQJ9nzcr82e+
mIrzEoCwO+c+G97nGvtUYUy+fU8QqEZfMYMi5XyVz3Rl4Yp0GZjXdaH0oIULsao7
h/6kfeDKmDZbdOZtsyEpGOiTY8+qK4lWC1Zl0UZ4Owu8sA0RFQd+sExIqAonbWFn
Z0ybo6fs3D+iCF3iJdvMymyJkOVJ6HqZG1xkOTYQVVJEDRENIOEVrYnwrX9O69ni
RJp0+9BYl0lHtpCgwApd6AD0qYKJBziB7vlZD2FHhT5gbw4VaDq1JyWwJleJXZBU
4xuXjnI8Jlcnnt1btyHNB1qtrUOrjGUNhIqvFQb5wZJqS+6BlCCP7y2/WpY11NYo
5fOXaKKUeMW4WB7h3c9m2Dhq4WWGaECI5piQGpQWIm6+0bgkHoHYVrHB0kUAW+xu
JK+qkRkeYMwF5PauvLSjNmNWc4ToJNIn/ItK/TRWMTubqdKYVg1d8defXw/t1qPA
jGUHbpT+Nwc9iwRuZnlewu1pkhpSSPzwf0WUYivnGhzFDRtqHbPGJL6fAMYEwkKo
Su8oVgDsspo7UTpSSg5vbxofPxD0EP+5gm+cFzbVrFIN+trx/MbTVOB973UIRnmc
Xzy5T3Zss1cj8RS7JUHN/pd9B3GX8sNrAEQoMzsWERYTnvfjSpm8kKnXfJp66+6E
gCoFprL82bvRXSiZJHP1Hi39XmeFNvm3R49gAA/PQLW6Nt4Sc3RoRLSzR55+F+wN
RssvuHUEejB3/7cvZwB4uvxArzc9Vs+AWKHCJHflVR06gJa+wGp8eJuQoSckR/3H
ALrJQ/qZ54g7lqRWepnkrfdzkZ52sezGvigHSvHikQI5DipfEdUzGhoiEDkq1YFi
YlQGQvrGSciAGHGguwYyJ0tKwNTtL5/ZWySal+nmlSyJsukR9UsaDI4Qr/vVKD+e
J/d9u8ZBs/dG7UdTNkZfdRoO/2YwCfstG1jMBZJIHN4Z6yiAFJuDxlh9xCZCBqvF
XNCU/CpYxdrjeaYJTLgvS+2vXq/6NUse8WrfJVF1jRkEx9Mk53yKys7nDs8It4b/
o2mIBHz5rL6xukj3MQEeEBUwRWvvPId2kJZ+EydbscGfuyOVm20RmRh+9rquzqyL
guhs1hj0T4JLDlHNgQUSbRKiH41FXUgggkm9G9BtjJIDpFW04YZ+SVAtqinKh1Lo
erU5GjrvPuAcVWYEkrpvMTNSuCMU67uONPWsMeUBaAuapWLKFus15qBuiKRqZCzU
q2ySMX0OvVAMTTggelEMFpbbx3SAHg1qImYF7gYtPwAR44pEb78SRuJ0LW3Bich0
IVjSgeEb3gKxyY8cP+nv61u9DKrYhVzYxHzrcyMm+RsGV6WQxFtaudaQTQN4edFh
5bnJs7ZzKMUy4gZqio33M2znRWgJyKlyFZPwpgevrRRy3jxZb0Db5t6/y7YSi+VE
PukTU3A52Q3fOy8hQG4rsEVzA8k/kTilGnM6VgFAU4vcXc4j/jxwnvRA725S2ukz
xYPtFnpX5Fxu0uvRtceUpN162k7EWHHXB8eDf/K1xyMMxy29gcgPtdWcqYWNfNUN
VIy8C/b1kMsJOXO7W5J9+8Atdmm/cycsfxoWgQN1lTtiv9Co5RJ8/SAFvNbyQhoz
mS7ntXZPsqgmQRHNMzcSCCwXDizzq4opgECllL8pO6AssvC0jNMIV3Wgf1/ATH/U
/9UlWtluUuHt4SZclUrTtC0hY/TTQnpiEg/FNR3NElG1+AQKu+PdG1NaH7mfn/wJ
XXqvacCs+FZRAJeQ/Rg1vAjKu7oGLhGXYxJLmjdzTTwuC+2hUOdNQUO8RPpEH/d7
LdY7rXcfk1HKsEenWF6yrjxpKWnFtHji8EEA7mM6/GZ4tmcMwzfyeuA589WYkA2Q
7dq8oK2yNB51e00P58WY+Mo31ZmeycO2apJRioQhKN04vgAn4X/2TevqxwVJpt5d
lY7MaWbt0JspNVsOr40e5vxE+jYGWFHLWbjSdoNYBcxfXqYqAB/tyirZO0ZDHHTS
YDKp14IScC7XMEPGBA4ZLbdEw7/ndplVpsCBRzAuNGbx250xiNB1/zppBkc7BlN7
8OBxtDx7X3hVDJkwl4ZrEgPfjcI6sT/YS1KVirdUh5CNbiSOie8CyFDtdszzFOIE
NmjfaDYKOBPo7n0/Lr0RL+FYgHCbfUznruIaZs7xTOxpfavcljUuetEEZOwH0rwY
cORRsnW3F5GEG5OjINhQ5vaJfXf0dIvFGlJSKF9fW5qg8Lo2YBD/eOoIsRpcMiHK
rt9uk/verd67J3djZWE44lAzUWbcZzLlGjMjIUEJOAJFxrOLADV8Zsm/BQ09sGSe
ty+m8YPNlq+v77CkEGkpj1bcWGGdV/o+5ENf33eecw1tTM+zBxOJWEWWAEcBKEJG
MGF3/Kh50nH/1NXnVEVt9mXUTNF+bUnoT24NKpin5umnGcAT+Tgr7UmnPndrQfG8
nryWxD4uzKKcnUuq3aEoq0fYfz0KTr9MyElZxGQW04auGSXPzoHhRoD+RyIp+h+P
o58eOA42/6Fst5hFB58C3TLtMdUqPRRW/wvA4b5deMpIGQ1Cy/N6lbomnpQ1sFpj
jVDwLavKelIt00Inxa9pl4KuGHB0qgWhxspGIY/yxWwaLHbiyYofFbQ7EP2E9neK
CMTfumyVlCSjcLJ1eDHqmwSqggva3fK4nKV5KEaNXEhVKGN3/m9FsODu1DlosbJv
7x3UB6nqIA0KA+v4fF9TVnHXqiGO7e1XJtZaMr0FvCcvy/2/54dX8fHj/Ti65I6y
Dk//8EmeloMrHVzy6uaDChSTLso7gvvw5bFTKUUsQNmyz/4/ZDEyVLuhh40blD7k
8zwtuPJpYUgmWrUlBfGtrAZ+Gy1vvetQApqEOnB7ye8/+sRgXwJXV6J+KxJtJGD8
QG6758A8DCQau6tFhnXuqspUsEMfmaAzue/vXVQhMK8ZusJ8XHK+aZrAS3ZfGVP6
k7EIrwKPUzcsAsIkvy5CjCRleixrBMuUm2dAH0jjho5ZxdOHpEBGfOl39BqY0vPB
+mpCovhONWBVQnOcr9bDZne0QPbTrO2bNvqw+cwYa2BxX9X4IN42wtflKhElFfaQ
b1ESW++mSyOvAVKlQvxuOHq2arEQWcBsgy9jGUHTRaAA82RMEp1D0rjKj6Uf46QO
9uOiLpPGE1O+iJQctk8IF4wabrw74U1KTu4lR3FAs5pvaxpyhZ/Oi0RrGTQLiU4m
FiYvSNRAwIEJoeBTRvO/xN8cAywuBYV68riryNPzMGhMYWNXMAUCxj61X59LydcL
u1LVyotZY/U0a8m32R+DY2lBZpkVyhU+0GJFhfGQiAohcuVrbBedsli5UeXY0UYC
rFJ4Fx01fWzvjq0AyzO0N6SGxulrXLzWVVKG/cKwBhpCTwBC45FnQhdx7cRjQJfa
U5KRXXYamKeDuArB2IxHfjRKP2Gx9+p8+1ewDMyD2qMMJdSMsKT7OwZzqZuLzb6V
VrdWwJgmnYzfa4yNmlmHcPL3mjSdazzD3FSBEulZAVkpZGcBQoj8PrO0Gz64rXhz
XLK3NdsLeloDcJ2y/Qy4zRDGvl/SbM7qVEk6eSHM6vMB9wdTNPoCMTIHAOUDVhuf
1wP+ar4dAslifpmyZhLBkLEt0Z18kTwt8ju7Wmr+vhOvkaAch13DsLUdVb5s1cAT
inPu3ynJZ9YGquY7PP4t5Q7edqji4NO5uiU8h4wNet13kuQoCeXUwziB049i6kxp
DFpdlioZxO6kD5LUxrQ1l9YO8I9Qoj6MAB/2X0eArK7JGYj3LBw0eyvrgISgGvni
NS+4yPaNOxlugL0Aqse+1maUSh2QtCjemivE+ws+6TCW2FOqAEhyvC/m//Q2SptQ
Zv1pBCZ/43IUqWJaaTwd6gmLKMriHDUsFy1sK+Y2d4MPr4ppkuIpUwF5Ta0PMW3s
Gq4exWjFe+eiRxOJFN2Aiq0vA+IFQ7CJP4T9jcXPX4iG2OVwUYvSw3JNKWjt1KgT
w9Gcp2Pz4W3bGzIFe1Qa2DvdQAFrSRW4It3TvMLVEFK9NNrHl5+AiYitrCKjS2lS
/GnUu78DhuMH/+MUi1RWigLiZG4nXXNy8WeWdg7Vco1RrSgR6aDhnum+srZVXIHr
LHucXVgIvcbsGOfVlDOc7H/G4mBIvdFxabTDSY7n9QrQKcaPSy03/B+MHEjXJpNZ
fik+6bBhBElQc+EHbE0reNJfBWXB3cUMBUpagJIzdBdmqRrMGGUR26qNGaNCWONt
g74ld9w4y0i4MAL8T5yFNRjGR5osHCUfqKtEIrBi/tHWUD6nHOMvKGFCIIBtbIdG
5JWsxsGfUWMRLB/7yRyExc+N5Qn2R25hkYNd/CGqExsqfrHIYWuGl11LC6EULF/o
SUwl34JACyxQn3pYyQ5YWyjCaLYNawURJyK2R2Tkh8pMCINPJG8BS8Fv+eFwGg/z
nXP4kVhccmXvThaBI4IkmHDCU2ILqupKX93ZA9XgyB5GoCPW7eVAcS5I+tLDz13d
kQuZopi1VCIkPlG4vlVbmui0WLZ4gv/P/7hE9PwkYtGMceDv+bDkNQG4RgnQSb1f
ZlZU2IM+2P19vzktNqpqGEP3hcF3DSrtpg5CO3PEk9R9Ua/JIIGMF+EEOJf0NiTK
O4SQ+b5rQPcgb/KZjDbsKRQT75w/Kaktyn/ekDPN7sAIl1QUeDfg39nrt4+aB3i0
e74HLVUK8UpxBmxnS6JseiuVXXfrXTYSWGO26UmgZF6NpQublEw/FNRjJ5eHTlwN
owSfDQ3F3khu4tGaMBhACAyo3+e7OiugoL19J2p28TIf9+IeAHGv3hoggROxJrfU
pz9H0pYxcPEhjIAR1gsRJpTzwQwPWdDS7jt6Ur4L9HU4IrQXT9/00H35Retkc4kY
/6GMLLfgzl9EXDKPYcLC32io9lEvDLoDApFajFhLsPRqBX3wIzO1JU+R8CC3Te2x
YMg3++R9ZirxeQj+/fpDrhWRQRJurSxrIIfuHuX/OYL/vb9u6Tg/3UY8uS9mboEZ
CpOrXOVfcU6YkeaGyKvvCLCyjgCxG/Iqm9HRzzj2T/5Rc6+3olkj+VMOoADkwAPy
G8ngrTCB8K9byhIbDwDnaQSBQcgB0Sse0dsiuXf5IWeuzxOZ7SQujpgxsL0QEjWx
uldG/VV3SqGpTqHE7g9AQ0AlRj0Qd3k5oBpXJS3GylqYL2Td8kG0CKwemLZMblrL
KSPgwjEc17PNyF3hF4uQ0n6O40TGtiMpFd0OBz4Z063o2fqMlwEVixaeWaD1pOw4
61HTjPt4vDPyh9sx67md7GsYtvJYg0k6VuF301N8ru4wuYiL1XLrmr4/DLl3oXyv
jYXUkd4WjwCaafYKJOQ8CSwdILGVYSQaaw6C/NXq/L54nxPqr9HgUtBrX7iYIdcC
XOzNiVoU3EBn0SCIHAFtD3PHq5yh5gvegoSwjzUZUNV7q0yDAIuE8ROZh2u/Aepa
uulOi52fRzIO8v+3MO8C0dxj82P9eA/5H11hQxpD5s1FZJlPb79do9pMwiqPwbtP
5jUgabhtudMAkV8/tGGG2r2lU7/CVwzW4NTgBw0jfrivM9/VimR9FlccARSc0t+R
lq2umq6htCLRXZKz82inGAcOvCCTeDFfgTEGXfW90rbxkIQE5iqsdp38PLZ/jdUX
4drI4gidzogs8Cdys3pV9pPhqDPgHStFnU/6jHiJdLb39yF0+NUGzlDqrzBC/GB1
BzAmMdU3Az5wwEcj/K3StaharyRYEyEwGpj/mPzhIO/XlOh8grSWCNlAGc8W/3go
ramBTbJm0sP4vg5n3sjI1FOpPnj1ZIden80NMxw9DEgO3fOdh/HiFyn1ABqQ9T1K
AEVwJuCTZc10XzoacAp0uhqxjNxIsYVHuBIIOFdJ2Tv/oRXAMn7/12fseW8vmE5a
UTXh1gtIOYLJztygiftRxCjWvolo06PfvqxO+v1UhZkQCAnHEXe5FGUyQm7n8wd1
XKd7OKKpSR3vCR37hLuBPs5vtXxSAVFG0YlFUr9s+5+sAKV9BZar2+7AgaS94nDA
IM4zQXeQ+qfs7fMjTv6Q4q/VWVyKlGCKulWYNZXQ48BZBHKXcEUcTyMBL2XVSYHj
kCAObxdeuI6kHKLQU9PLxmMEvU3f5Xjp4UKnOMcT6I9Z2JlI3QzfyzlovAU9awEn
P91Qdy1ILnHmgX86IOO/LtpJahBRPY4gVUsOdlQaG0rG41VRVt7V23f2fHTw8Wt3
p7ItpryJskv4NLqKPSDhYfPPfmlThgiwqj0pGV2uTNiF/ALmWutIJipMdyJmPMY8
eolc9di4oNso06xVRwnuhCKpY8KVKNVhCo15tvehe4jLJw/4VM8VBcq9C5xm6nKP
Y3P28wWByZCebepc6KLvTd/bhdGrH2Ltaiwgfo6jwAN6Ef3oIdsg7VroH2hhqsUH
iOnANbTtkxayKuyxHegqwW5O2D2xwry8xKraQb9KheSsYgNr4K4zPKXJF3W+7L2V
odjPVE5Jf9gkfSf8ngwXcLQNSDmPRvJt0FfrYYs1o4Kte6mTEzP1+PVtSpbxODpv
HzH2VR7KLk9hTlejjF4gDDOLuNu3oiOQNCzN6MPGM0ygEieJxSP7w/DNzrs4AHiG
wf//9ktunBfkh3VN1XO2cJXrarz7B+ILBboFLCgk09hbhEwqMau7Lk0PPpqopenW
JIRLk+T1wHQi8O/U7uVtjL39uJGi7eYC2j0OhomrYnM6XIpjVwMVJODqyRkDKG+f
WOIbhX0J5+1B5lFOt1emh16tndsN5EfASZjm38OV6a1JRcCR9kxtbP+emU0ovP1x
LNUNjBJ+Z3IzKwiXpzfbMQwa1CrzIFtLLOg1+6jnQfzRrTJD7s/4MTho/SH/gSPY
UlUjRvUVb9YTHIgjBEfSXqAMMIyofri3Lzf960CWKp7hlOaagrLISISEVXdRtLEq
kdtNKNzMxVT5gVmVelCD8jjlPUNttyzHGQwldwlT5Au2SODZa6j3uTlpCI4EHBMv
njrGziQhjdAGECur0FI8FGTQI1U+kMQoDbIjVN86OaAj8ovclTSNJO69pdAUceRA
oIjzw9lcgpYYZYxd0bwbb4vLjulDlzyXnPHBzb1L/vtPNlN3R5OEckHxKsCWLbJj
FfcMg8CoqRP43sJTaWJm98hwEh9Ahchded8vMVwr+6wKITdhVER8vUhaXt92TuOu
+HDaw4UxnAWqWaD5s5+dwi92h1zhESuwaLzNs4QLA2qMIxwP6dxXm9JUOnTRZGbN
el3gZROU78LW6Ol4Ah2hYVt3kFcBYDlPVXA+Giz9xJDinvj80WX2cHXVnNAh3Bc6
Duz4+ey9rMTuDBmnKhNXNW2i+7T22yyBW0hpDZ61m8atbJwPSDsl9R+7YNtF/iYh
nePCI3Hzmpj1j1czOYQ8lsvLJ7FzrnoR7n3vbfpGRksel3ZwjI4Hhh7ITYjkS9TW
H/mxkoAuWHtbtF6//RvRqX9tS5bBRmSL/ES2oVm1CpvsC3aEv82lLOZ4stZ2Zta1
yM2xqYaUwGbEoQbNGgdhxInq7dj39UFN9qbwgfKzoXr4g+Utq4RXshSdv7d+wt+a
cBNRIAtBlBCh8zN/fVaVsrnCKHIC2+MDuSTOJp73nNctfiAJgyFzC9VDOPkOVolE
tDXjOAvLfU+duSHgXgbkuWSBL3rKBhG7XIO0MFNyFPjy7XpVdCf6WZkk6lttXYB5
W6RTcdh1i7J+LbNfejewBpSXN12ejL06EqZXeRv+bXIqRQ0/XIVslpv4ScNP61bx
qBUYmbuHTZbIZVSCh3Wo/3rKtwSTxDYNiWRihyiLJzuhJhDnSDdZJvCm7Z2gJfPM
6UGmUyhyabgwrdSrnN05JPT6SQHXFZR8JcRaNVw95lXBWONj07Gk0bgZlX4Nw/4l
nx+yk3tYwkIVk4dSGsUwQAtAo0hIY7bOoxRxO2E3ABqReeZROc7JM1dwVp2ytdFm
wCmxuSNQ9yceMxrU+wvRBsvWpSqPMuDjAnjZ5Mfpq3ckS0Vm4yjY1h3z+gt+aSNZ
fgFmOlyhFZTRCXfLME02kq/RpV6vVFuzieTcHC2ak7pbvtG6DJ9eX/VIGdLF3ee3
ZDJeLhUwTM190PNkAVpLVNkVVUdfsGZZQXjWiSuFusL3qnavFHMkJygATGmnQcvf
rHsYClSra/mxRJhcQ4zPMorWfATqGtsw9wxzPlCXCRSOrS+tUXwUX8MG0GhCUvl3
hMGOvvbsdyGH3wL7sA+oHqHERj7qrTRITGcV2Qva1H4DTCBkJOok8LuevnabWdyJ
TSEQdLFCPkVjj465ktYMjLVzyZGgyQqwqzsLn91w3pJWDzvE2FA+HKM+PZWJXUZZ
cmiXkEXTMM6ZCekWhuXx6/06HEmtprTBu8oU4QNaY3m8uQlhKTQDnr/L4QOMZBue
jFOA31If6IYY38zfhugtzNxv4zSzPMtWLmzqN6cEoUbYO+9VCIeTFw0hdLV28pWV
t2taEWfbm2jzGW6zoDeFytcxqUt3qckHxcLi6tpElv/SCUUc0zx5LUSOqpLJKq6k
HkJf9LJ4ufUKNQl4XKfytxYzNDSlzZtuNH0DN5jfwaq4erC2TPtQggKtkSSxDXdV
BHYcXCgp8ZUdASw/uJqvIxRDESf1NLlcQFOfG7QmBk90PIiDijYRaOfyszdm7wWH
ra8F3yrpXiPZQ/7R16TEOE1niD1pL+8WMAvXAqw0I3mhxT6NSLWY8W/DSYwS9oaX
jaGPU85R85RDC3zxgMMWblW60imPaA/yRidgwVmboxwp67VzjGx1YLoHIu/v/2vY
KvIZ6nkVDEdlgLGVFu2KMD7MHhgLDienlQg2iWBDZko9HcZPScGdMWEItTuec1M7
F4Y2orrJW/8OGZf4qvVC2kpgvS7b9b4KNLnODl1EZ0YiL4sC2hf5UksWThE74Yfn
w2zxc6MA6spvU7R7jumZXYxHEeLpQIeLHXnxOEvZbMFxOCHAe0xLfu6L/CXsnalu
4p+M+VPEgTtg/+3VKcE6wBvY89EUzf0/q2TKZUdwRxuiMVR3baEq8uaGN7hfIffU
fOFCkONFsS1AWr4ta3zkPqYRVpl3RTe3o6tzz67DswQeZ9AUutPEUSbQj3uZ7l/R
n3/QDxjPWm6czEfvWojpTpCYpAQicZb6Yyux6tGp6YzPv2LgQu4HNG0Fb1Tl0uo9
PAAYHLw77CZ4fIYBE1C6O2yyduaKPqLDxwhznzb/0SIdgV70tMPlHTm+aQiT8jAW
WfyHW58C1AKGUPDhEWOLSVTSISM37TQJcAdY+R9hg/xcXD+BPVCMav7ezNWBvQc4
J3X90SjUG36EiyjkJFUOU4DPTFgaaHiTTPAAHvi8J011xI4dwG7nI2B4g03Ejm6g
TxkEW6VepFL0T2nm+2o4jyGN9f8hGmopR6pi/F82WSXd9RDNDuZjAXS6AXwvB68Q
pFqBL+tSNVDrdpY0bXriiUnywO6RmbXLjU1oXaIN/OKEVRv2wRICZBWIvrhWoPRB
YBITsvAVstuSVAFFWSRg1de478UZgqZc405+sU/irscLkWEJNF98MfLChzn2zwWn
JBDolwypddLeLZ2MsRWe4jzlbkIORcMf07tTjOacTUy4hI88/nb4MYgAcJ/P8rrO
f4QJsEPM3ybZ0g/jAj6wzBsG+qrs0WjPb6jSfHf+D+3TgjTjC8aFLaz9v7RmaKB8
+qn0mlzsuRMcKKX/VpwifjHdq+2GLdDLZ5q70fUagXzM8m+ki0H77QPBYDOmzhze
Z4Q3BXzNwsOjR7UxeJpGGBAB7lw1BEB7lqyDLaq+bAgLF+Ql5Zi1tHKHif5TAAJj
hFtXFmVGFtf+u3dAo/T6MqTsvevAfLV2bFxcRt+h0Ozmh9xMYDYQv7nu81J7bTPQ
oeJKzY5jbc6EAWCyRMAjCNbuiscJ9DI8UxWU8E1Mv5S2AfEqbEXmUAp5R8wUefdp
s74kcvR6+fAQ0o0XJm6RBvr5Jdcgk2jCPJ23f2GP2KNcziHATCgj91kXk5fRzt4g
YtnPyFkIePTyeAU2IHZQ1V7E8KsFgNm5XVWi4ZUVvMz5/1iaY86NBuG9WBhBDjuC
+CaQTaTxdMKPakYvU++R1Un8xnAfY39w0Ftho0gh8g0LX1j5juCzkcJhZCdG6TTW
aTlPC+2PG5pidlidMQQlQ8i0aZuvnOedX3wzM4uajdACL9doxTRDJajCZpRDl8OT
ZYdym5Lp8122aJP7QH7c0+JwTQeWTkq8aYZcVMjjqlG/8Ij+bLcphP8KPpDDfWDo
Un0R8Z2nlK8v4wojN1JwNPeXs2Z+oZZ4HD5q31HR/qgHDfI48JFZXwohRxF3zQQ5
qKLvgFYz6RDOnb7DohICb5qrbnL8iF/6Bwa4UnHP7v8WknuG33py22GYPOJ5fiM8
CrXfcHs2Mi9FQYutKK4fK1sX+Jw7Okp1dnvxDF4qTn55SI6qVmog1QLD/zGa5NGv
txdMmaJn8SGCS2dcRKkwU/KZimGSRRKCtDdbE5xUBns2p7VO+iOojnEfZ2s78VJn
/TpzvmVipmybt5P2GnZPlY2AQ8m1zF90/NZpdIWOrdXkVapyeeJAwdJCbEaDEMTG
QzllDGzy5AajtFVsK6HBfmDIqi0y7LmFvCwBb82cxEQkSow2STecprt3k9h1q5q/
FYO5KGVxTPnCDdWfbi94nr8OXn2mxb2w1R2A7ZW56kIlxeRVsuWV9Nh5Kgh+A9Qb
3fDHvrgkFE37mzJ82ujvmNoReyVXjuuMQAIQ6Avwl+QRzalaR2DAvSwprJZLGVca
ZFzVYOVJc2JERx78wbRRuxWFhkMjSE+f1uLRdeDcylr7U+Q7HMaCKV5SbB69gque
ofIl5ejO8hzeJBObhLnznCExVxLXBIOroRV3fSe3TRo+Lv7htSztYTifP7hKzrj+
cr0+TaVfZcXxh6RkY9lcwE1mPwIDcT4K0+mYf7oeCBfF1lgPiU3AxcLm+kn6v2DE
JPwXnvgP7kDnIB+ChaIPoh72Uemn5iYBtjpGSk+HkN6P7jzFroJBiof5I6KYHq9J
W8oC4wMOi0BT/wVfrW+1ZmKOzQegJgNWo0486qhldCGns+gmVFotVz3WdNW0dMdC
xA62H86dnjR9aCz1TX6S0/IvwQ0jdS6TXLPJ6OnRVZ8y/3QMeo7OzySFmd8pGQFD
ZGkjOjTmDuGDnyXCoUpLb4dPjr/9qnz4YcMjBPyG8DLBXlQakegqU57Uh+7FcNcw
hTAHsif7VnHJBkaYYMTVt3tfBiCwuwFZ9bIZk0mzrP0THI7JfYIGHU8+xPxbON4B
uDL+XCsroNqxhnR3ZsgVB96KAVTyiRI9Bz9CsNhRiz6UC1uv9bSywMtyDMZmdvyg
FJTI0hb+RyKPa2gCE5Y0S7mHflquY/+AcsksHJGoSSZZ03Vg8ZZ3F9bsf5Bicwew
pjILSmcCKPbQUBF+POyUPheSoFyCNYGm3eoPoldXGAM+UaunskD9/lmfD4MdQav3
ALW28K9dfwR62N0TqCO+21crIEPr/E+iGPEe+B/YOaeHu+Ilowla/oBfpK80Fpki
5zHjpNd7PJhq8rBhh1rO9yiMsVscFzK7Vp1UKGgU3EpZ1ZdzbnCgoQfvS4kDAoMK
+Xvk6HFVPOv9ZNlzILrZGI1iAwg4PzsJJxe7FfR28C26Ggqj5/+8eBmg9QKbNXIh
En5WL3pGK9CpuNPE74XvM9ou0Se0Z0F4OBEZgXhFUTFwEDe7NoADFL0da61+TcGC
FVrYkU7Gbioq6N+ueeZsr1OnKNkOvuy1LYAEFxueeeN+FBv2oiTZNExfz9oEoRV9
qes0UJbmwHpCwkCfkzPE+hPXjt8IT4SkWUodCpUhuIcMuqYRQv9jMSZlOnS2N9Qq
X46TKx74PYk/5jJy9qeqCux6OyWOKB6lCrx5rjlpsK94zg+NbOgOdIhdnsuBnWRZ
I6o8umBZrdcmGH6S1R1PWXTYLHVVo+IEmPnSaSPOd66CTPO4EhccmT5vB7OSLLvY
HT4GjLEmSkjnwKYWInKFFukrg7LRf55ATKRTap8ci/IL/zzeHG6A9PGieULhD7Vj
Y9ip2q5cf9JRbkurMxfvU+WOO/ohWk4PjXn0Vg4PCgJ/UrCd6fH2SlZ7B3Dwzc5+
ItpnBwcXxJci4p5luFjmsAS92h9ndCTdY6IFJU7vXuaqr5SvjiNaEm/nIXAJ/D5Y
y/NrMzkV5aPkfVnCEl3j0rTrHQTtibYueUaEZETO6wDXdpgETmGRj/LeV6feUSwT
tfIumhsPffiAmh1ZOh8WDuuEewpfRMRNwL+pb4dQGkRbIRvh01d1RPaS8ZId/APy
nWg51Js4InGenKbgQ7tWUrNoeEcBw1JBj3KiTtuIV40kCdkFBgod5T9ISx5K2HUJ
SzmX4Q7mk23ojmPcMUTPviCZnpQKQm2RoVXWZZx5Yw/j6FzspcIpd4873HJcD008
5Rac4g1TihQR2ruILdSC1Ir1Kc0xdep/nRJXzqiP/t5bzoIEGuCeeH99xocTlsKA
ifRxwTaV22cqBdu57wcOl1qAw3AjKuOrsGiMdUDG+fQ4P7bYgi496185Ip4WNV2k
ihHnUtQFrQlESeb67d8DIzqL4YN9/Hw72xt0ASuoguKtbLIX0c7aWVXKY6nX74D1
4yN+nmmTCucnZjXMPe9cOGvHg25zVM95iWWzrDP6/F6S3jPZhmwbAMP2VuvFkfVk
el7sblYNiqMzeF6/OgixTv8qjRt6bAQJbDtvRpexo1B1NIzFJoR+Gw1Gkb60/OsN
Np0yaISJWwsAlGwCnxiZwxoyuwXgqDjTyLcgN4tdeQhebVeSgABrzekzUtmDCwAc
g9yAWcBz0DuxWYIhMtts7J5SJPHMSh3yrnYTErkd+stH8t+auTBHqS9idQhhr+9X
iocSFynjrMNnz12fE3NmuSWIN6zYsVcKaUo1I6bkCgyaKxAOoGO7RsEFsEzi82/5
lDkfrTGEemcuWS8pE/c/Q+bmY7EpsINYGX17vFXv8YcpK4aVX4u+WeT8TQzMsSiX
Yvg8RbaHMASDhQdYSJivxL7ocHZz4XUSg9kd99gxMjknE1teVtp9n64O05g/+XYH
eBUuLvrFne1MehuI7n1u0uiz1jW7Aw3LjoMNPVKpIKMdYCH2XuMN1FTm/D5kgypR
KoM3eZN2qK7YwKpIp1ESqQc2yBYZKAxXmG6dPdsWxFR0nbXufBctb67YEQxyOA2K
uJiur13rYdeS+LwtQsqL5RlFFtQ0dEJ6R5pAswNg4X/J45Q8/m84TMiSHNkE4/o2
olww5X0b1KhQkauCxV58zJOd3vrWP10engFOhALHy9izp+8pVKAw0BlAxFIK02FJ
othnWkZNxdYPodXYHNn+7lw3Owi6pJo/9rT99CLFz0350wMPWYI6jJpNeHwyipyo
pPcbOlZlr9uJnBjVuXMDFkIyCM14KxfN/W1rtNnVLBNcO2zyKhhhCKzHTjd/Nsm1
Jmkr+O1YlhJr5wuFwEAUwn/pW0doNhHuXahDP6ovTiN4WmQhnfMJPlDLFCf1t+zt
YqqBnSfPek+1WWcO2sosxSrUundeWJqMR6JokbscfQSr/ETrbnTbJCJufJdZfOZ3
u29uk5OqLCS1JX4CSP+SBE5QgSlixRe1Od56hs4qxie0eAHDycwzM+tg9TFi0//b
Kk+NuTBDPJeE26W1uJrWVEB+2JMsMESW62DgiYg1X1ZQold2lkAnRvMZwXEN22Fj
f13I7h16nu/biXk8dAa5zLpCkyCtVDLUVXIHz7YmDKxbhAHR3dfmKyXIPNt1jSq/
ZcVuY3IOvkIO3BYXIeYk/5/TbNfmV4JISaKVn7T5qMmNlix8fjqIOOdZSoNF0FPW
Ze0IHb9JCRmXbQz8X+vdNEyIyTrc9AlfMzTrqcnTfEHUcwcGU2iRJNEOBXyMMveI
0oQX8KgLGl7zwfghikmHLlTbQ2T2Ox914hFmovK7yzcDhrtQ6/eT1qjqbvKq8pdg
+IC3wqa+O4n7qdHT4MILulRQ6d6vbMTaNTGDSiA9aAv3eMCbXK8fTQJrotTwBKsg
2L8Kkzsy5xw+eLlwJSBjL4ZTyAhk5Aw4HCHUE9YLL9JPXbYfbPIE8IzTP42ddMDs
+OzNBXBq6lFLZVqH/wYGxF/3v29jdBuqUReMlSny1tH54Dqz7veNTqkREznr2zrg
qmqOCkDxdXo+yAjVQl5sZ4OCSwJTN+p1JaLdlA+vHs3gcKyxbnEBDjmpBu6+eQNY
AnLRVajIrNDQ0TvXqDo6cZu8GuFAdJ3IbaUeHmBMIC33v7Det8fXSMqtUtJN7F3e
vtSDE/saRcewUs32AYT/dY6ZSK1gvi7PLZ+biQ6gdS0ur/fRmMpEHYfz7e9jaHZB
JbPw3e61hpeBfyi0atDCcbmer/6tciJatsin9yO9I9V30mGDeNg1W7b7guUuGbzn
1kKXH/dRMG+VNHZ/nT3tLMRBApWJCR2/GRm9JDStj3NJgc34WybJEdJe0MhSVBQJ
oVrzLHfuFDg3Wy6W4HL/jeroua/kvFw4sdobvS9ejceaHIpW6IoM4EK+0glt/E5V
UmCRaBaxR9PCsHJE7yi5bezm99pTmbFrH9UOsxwKOLxCx9WlYJf/Rl1FtvdylGc1
MPpQA1U0LDpU70nTX5JXvzbIPE78l1EyiCQ2JWmR2TOBhrltsSCSYpI6ai/pSuHl
mZicfVCYGv06zjv4wgJ3G++NB+F9+JFbrmwhk3xNLxzmpBoQo98rQ29g/SEhRRAB
NmmLz0zGPQB/hxGNXTjJ7xwZxxTDxLmwiDw9N4ew6PThRYEgFiKlF2IRlABpU8UR
pgL2t/yRHep3+yuZbX7huuDgJ8hYy1G6CbDwxCha9w39v5T9g5AKSKYlZOppv3Us
Xv0wyjhxK5Q5YmYjahBWlInW074UUydPSGf/zOtiGHuPfDPNmIvlqhcpI3FFTBkL
i89R6sYly/K+3dGRGVhkSkl61s6vYg1fAwmVABOhvTU1WWoFfaQdmm4rVamq+QFh
3EjWOykERy1Wer2LcCVr9UYfONynrfsic8k+UbLnH/iftjsV25UYhF0zBQaKh2uF
WF5hq4+s+d5CcmdgjlpKngQyBSX7HjvkE18RcXU/mzAZ8/Hv929p1MSLzTVQejxu
DEpfhMb8x7h6Y94bOSg5OZGTFbZ9wwxuo4g7jw3W/zbRiI5qJZADmesL7nDdcPLa
q47OcfwSwedYtwp1uJQNXE6C+P3m9xyMx9f0Ndj8Ug91AXrJQQHEOSIQGKYyRssi
bSlDrGgQhK2CNUUaaglTi77c49b/bUq+Iu/u+qfS/OkwkM/IRItshAeitpl338nU
bjG33u9Z6qFQhCNLB39PJEMBi1gyByhr9FF3VyZcJ6UkY22ZbDnXCR+He35HDkIe
xvfn5uaJGeoYXQXP4Lylzbp3/XRbFMfbk39my6CIo4GEdcxy5bTGr3320YzBYM8G
gTvLjpNM7+daKYOPzw2RnGbUUx5tXhsZj9EkiAp4zQxq3vca4QvC8V9URGu6NtxY
fvGpEwzunqjyfCMjC140rhZ2ceiNHS6qQCATVVXv5UqRJ+mRw2dDR8zFIdocDvQ/
DEp16CW7ERGmk/B0NHG03MKLJR6cbzK5LH/UdYRma22tISUXVmj7Srfz4FUMoP75
y3IyR4/vFs3MDCpJR8hCk68UU/MzWAmjhR3jV5hQM7Zeqfl7xSkJgs+dh2Aw5jyC
VoX/GrDqCLs+lKA0GwrH7N6rJ6Vdk0jmAK/iNILU6O8uyligytAs4voA9LtkO3C+
0c5nzzCr1I8dyCqZrIQKfR3rwY3R3LYI9Cob+dJFcCW5QBr6s3rvdNBENJn1xZ5b
A32Qpr66Alh56l+zKEQuy1Hv+lclKnf6YEaqkvmvyYr/+lnYOpxfirIShmo+xOUh
wIz2hjbrTAktaTGLtuue41lPwFwOd5fbMtVR/w1hEaG392/AUH85huhIjN78iMPK
IYWTDFpcHLrF1vEzVTx9PZ4OBYP134mrgkom7nQqsQlu+uiQoxvCL1wYn+NHIWJo
0KDzC71U524Yl+gr0HxYpSHZnZ9Z9sn4gdLW51JF0CzaRDHmrQ1poI3Q7N0kO8sj
2ekiDVfzxTQ+XWjkqx8rTqIeUz61ykxhs8b0W637xDpyO10DEJh8RjzlTDv5gfdO
+SQ1wPZsptvrvpBk9nFCtx2pMrzHkBke+PqBG3aMq1DYs3rH8sBxDLNuIXjZqosI
y5sMN+iSI50XKPx76hL5yXN4UqrmmIkWWt9ULAov2ZzK4VzzzAdIoxKdviMoocxK
JsxxEgmx//G3DGkzqGYa0p1nr3WNxqvG0zlR8qR1U+DQ5kgIFVcd/swNt27O0EPq
hD2au8zbjrK/GpUBVXtfPet5m0RYnn1LqJrnkP/i1m8l0tJ4i6IOGm1OI6w4XYEE
SJ7LDIY7CCGGzL1PeuCF5llNqxcKidDARIeYOnrBh0Na1F9W2eJ4T+TtVgelDFdi
4dF2htX2R3pRTXHNiboENGKekkZagq9eJR5ZcDVGk8XFLBVly5c+1uy92AXsXjB8
W6IcuSRPnhkGeGIa34HapCPvU+2gHSgOWNzQ3AxoIv00WyzPk54aUxhYHuhYC1h8
Up0H4VCLVToABQc4rVVXPl1wo5hh1eJxAYg4qJPuqIJE2wf0+bEU0mtsHM3/sODz
HkrzzZrGszDK9A82VtNVikyDkfoGHV0jcL9GsMZm2vFcBT0brCqB23xRGlWd9AUp
jqktT+4Qo02MbaHS52yhzvxS10q2i2AESqcVM6a1I1zRMaNjS+wjn0yXeUn0VchN
iWnu2kBUm7cUnjW8r3zAQTEvKaIX2UGhw6rSOY9DlbmnByDRbTCP/3uwLR+CV23T
pvHn8yveFWze8hcF0YObynZxPc2O6mWL3QqzmG1ThsHs8+hW/RMVJrzu+Jd+Dkqk
JB4H2EF393C06CTxJkFI6cg0GR3/Gy0sNc2XRUCQ93bqAuLtxmHwsup2pCEdpjgR
LKgczCUPr/rB1GUb8uKmoE4KSdrVWrrDFlj3bWN435ylRqexF8IX0dQI0uyy0CRL
NVG3gCHx+IU4vtl2Gg7hiDZsacFrfVnxddf7ovc1LcZOdLJEIT+v/UdleIKaiS5+
Q8PgbUSNSmTA0jYlPUVanENtdhBdSPYDatIeCRlreHSyTQXRD3kjXlFnWZdW48L7
0IcRTnpTKBXTTfam2oLvaymZLfpaOBJQo6pTCQ11kI/iqlgsBgY/io41BbpdsJYM
yts/nvGMNRojGWG5szrhtr6h9u4/Xyh98dSrxmXeO6lWvUCrGRUjxqziTHXm5Q7k
LcLoNLhdYBKasEXFQXluQB4i2LxJC3Mvy2iqEXxO671gGw91Z7LItPTNTqPhkJiq
fnpn7Q4Chu46avSkq4SbXBt+rOjAa/sJoRa7hkbGl+tQjTFVc8nU45jHGemvGQdA
lbd2BgcZ7xMeBjGTg6TpDZB1Ut91yhNBNWwfsM8yuZi5L4fKEv26KuPF1Zv12lWJ
U6w+6MySe8FgFNcQ9CxEssgU3O5VxM0uV17sR9pB6PTtEBhsqhoWGAMTjlmuMesU
sNVhsnISHzRuxpChgjiP/F8Ko7WzFP03r32toEJslIjhJwNhdQRrzQO7LDIKme7A
q8Qm5CcK0Jv3lV3ZEFcELFXjnDaUZDTOT1sslcZYeIA1ylxPGmvso1Mk2/BbGM/m
mxqUSzuGZLuOweFT72vwvnit2galvE9Wl8+sOC6ze4M6seWiFD7gZO1uS4DZAS5Z
g85dhJ5SyY7IzpSS4yusakfbh90rGJ2yqFzfEBBGnSQdFSQvWgMA6OJOPVHPNV6k
T2WJNG58sxAjj13l8Owhi83/u+7TNCJ5pIifTC8CkmvlTNK5pnnyJST3vVbyqrGv
tIX1f6RmWWTmNVwRIRsgbm0ibkXHenQ4NrlEzvUIq0GLszBONPd0XuOmlsC8mIck
/cwMpcGePWK2SFI55bdFvevAshSukWytH199RC8rS5829uOqfFp8/EXYp+nSHHIy
DgrytNwA8kM0TiuS/MdqYHEd9QP9WdkKty1tJRRO9mljh8FjO3YYjrByswzyN9GG
itT4hw1qBdDvOzXZa9cx8RnR2jpfeYbhcjrqFnS60BNmHmCSvXe8eN0D/SzDWZXk
Xx8yE0swfjm6F8T+pjynk0zSUyKEgizLw6jtbc4gLuNjPsLwXQXLbquk4s1tamDB
bfba5Ep3KzeNU4NohYN1o21hn23UHS+j2gulfCluc9Hr3brAdov+VEbEJKJ02Gav
jjkDAtA0RB7XucqhnhIG9v93ltSmSHfvwyxe23GrlUNmZnkYgBiacjUpupSly8vb
ToOsBf5Lv6+fb2iBIyXfwfNKPlG1iDst/WuLLvS2lWwzryDPRbhHYDru/LYvMNgv
I/ZA7zzfmDWIMAaM0NGVvIPjzv8/2DOIXmldoTcexvfBFnOx0p8Reg/BLatbSkIh
gLVLfPGxOIRnnJzPC97TXhS/SBDYTX0jXFxzCsnp9Bqt4pEcv5B1HM8Ibz255u/I
qwRo/M1jdZ/sVOIrAOZWpvujyQwzrkyr1GLMQg97QD+4BPfI1SDwBiEkCBXI8HMi
RImI0bBhqnY6f8+QGWSTjm7TGGaYKfmz1absYDFRKW3HCIUZql0PZtNjGLxy5jlT
fRhCN7N3rQafWsSMneyFQj6BYCr/T7BvdX/uu3zzE+3vvrpJfykRRSxN0zj5IQX1
lxFKG8A2uynFVGsQnob/9sxrnkQ5uHngby3jMCui+w+Ot+KHfiFMp8hzEcU7DV8s
CZn3u8f8p4SGwsnJp4V0+BhTBNTm+RkQFGtGqYtZmbfRLg2qCeuhvYJnfb7c05em
djXQHUwx/bcAw8N2w3VhVpvRxElxb/sJamz5efzl+N467lsYJkIDFff0w0DgM3wW
m/jbOG3TSCMh4XLAfSA6JvYGjUvePPo9W0cUBznQlKZMmrjcl70NcGFdJDb44Ltd
4dfLoEEuy+0MqdAlNuIsGVVpRyy/n6Zt/IrqLRDXdUO3QEW61nu7kH2dyg/A3pAI
IhMSw9snAoHKlgLFdW5Xc9iSwU9PbD39PikEObmp+WB487/9sE+IxqeNGbgHuzUV
pTG3Mz4FVIGDDTa6mShkrbdFtxHPPAIRxXm1nfxRKGa7wS2qWGyb5b7kulSqMCvw
Xk4r/0dYJwyvr0WliWulEsczdGfJX8eyS6rJMPAnVeTfwaMeQYDVoIG0I+J48Adk
qvS/xf4XdwvdkdMDttTuDnuoRm4b/YST3ucIxgqfdE0iIw1sR/iSnrWiB08L51Zj
ba54p2ebqjDdtXRgjRboupxpGeK6o8y34yb4JYhKGgycVSbKatE6ZiaW3pQz28G9
2jU/U7aM1JcGPQUgy2+2kEN5ErkNDLoQ0CGksSo9F6qBw4l49yokeBHVHtFqHLpk
S5YfluZqeeAc5H+TvGf7V7y6BXDaGreCDNYj5pGGoBEQhkaWL+PcxPMBU0tkajKI
u0aTqka8j4nFLzQhw35507abLltH9HNhLvCcLSOpE0jDxLQ2Iv+XvO3WiqH2AaSJ
LYZjZiczAFwZ7N2wZx2UscUl9ORNwxvl8Mu+PDMZyn2nECuoptxV7s9MwJF7fjq8
wi5QlmM4f9UaYDto4HO4kAoCtUUNaQukZDdr8Clmzcc8zk16kIV+ceJhHBwULcgp
k1kuDZsUvuLaeRJlk1BVH0cXcjH68GYkANnx6tFYOGziJF0jmnX9eiWjYGKG8mvm
20a7gU8gOqaZs/FEhxLPNuuvQzd4/wWBH0aMxi6GXLR6zanPN6nDEW5mJrWE2//3
/UEfRpbWkyFIqcD2wefmymGHOfxUU9wBVxoX7sSHGl9jSbd2gmliWEDTrV8CY1dh
/2dk4i7r9SM6eZ6YFn+8jwPmZQwCkLBbXD3bu/h8xV1iC1Mojyq5f9E1pOnkV6Ps
c1aNMc4R43maC85EEkMY9HCpaCWp+bnqssMaiK2/ON6NR7BBMBWMZQTMhaIGU+Uy
bMHAmU4gk1KXUt2+C9BLKckUGLE0czZKXllXvViaEBW5F1PV53XkSWpBa8/gwKpy
v6JPfH2VkiYyeznxHikzDwTyPESz+qQhH36lYZS8kXYs42MZwwWeM7ljYURy7EzD
7BP2FifLRGrmBCKcf+PD7Zt3RQPUpzI/Omow4wIqDIlF8WVDKb6ObBsx7Pz7x08C
MP4CVNfDGenz7hfnO3YyZw9P7Ft1Wsi3FHHiypVW5RobUqNzrha8LrBXwYaCEkU5
f6Pb1m2Mj7vNULIYQdOIjvSZOTAP4t0rCxoxhb2YyTiJFjbwoPzEmEAU/7sir8l4
68KcwAijxhaVdqCMk0kN0215mH42LW+D5AyhVDJaPszzMMQghIoxV5oprBHRiMSF
jPa3+p/5y4c7Le6q2lDLpo7fvLGxChY1Y3BWC7mZhRc4FVY96HSXQ6RiKVaS9q4c
FT2ov78sicIMs7LytbpbE+QuD+zsZw1frKjqc0WOf2tpAWyGD+YTLt6USmKv5uBW
OmnvsE1HnZX9qG9jOJ1svSoZyD+00c72+8GYyEhflgCNBd0m0fl3KFO9RLip9QTl
Wh+KTPdxDHJWxfOjhXJeZT2I0R4178j8qnz5MhhCD4iujSPbIfpRvicR46E/Bxb9
Qmq6tM11NtDPr2ytfh5zXjlegHsg/JCICNFpb0VATJNeEM/ie7QV9ChJ/j++Ae4D
T5rJWIwaFkA3rZW8OrNH5a+rVIwi7/P2Tk4nkd6sbLTvLnP9nVApTsfSMrXdy2FE
n+gF0Eom9FOywoTL61UYgzIIuEq3Itwye/ofgD4CC9WYxukd7H0lEC7X+RIrn5Fm
eAM9cojXli15u5I1tbhkIE+mB359/b2/fELgUkmvN1hvko74numodG2XD84qKdfG
MTDG+wECSI/vgPsGwiteJti281YJA9AjmfnQxnIMKZo4z3GTXjcPAEHtXP4geAOB
M+eJkCdGDRP+AljXee8tZEzv7icrWA2r6VnozlxeXugQQ2+HN7r1M338NMGdI8b6
wTpJQAodHXTzqfay89J41uy7ibZTKOM46Ztl8gqeSfitLYrNscuHu1XBEZT6mqXT
DOIiEHxF/prFKWfUhNnl6ZaN652dTQAV5J7y0iZ46D9zbLTs/AiycW4bjiyrF4Ml
aDU2AqKrGkFvCM0Sk0cAx7073RLc+5vsD2CdEQOG6Un27DKbk7qw6JtEnBBJYQgo
bzMZebngkn2o5A3HlhI9Eo0sfg+a+Kg6KAB3S0yMrb9AuFFTLpnbbOsWwjh0rUOo
i85u+fZBB1OMInAsMgK29+WSR9i2u2LXHt6HcSQgXSP5zLyKsulfFrPDjkpRc9lC
tUmxvo59VTkx+c3SwJC5yO3B6zN32qCER8ip+Xp1K2zhMFeM4CYcPxHtbLi2lkmQ
d6ZS+Emkm1yHoHe3JNpam3bDrFfxOAprB/0dXVGmc7P9914cGSNp7jbeeme02ZCX
7AAa4VDhko4j3ay6ra1AJ+ERuOHbmIQ41Q8kqmC2TwNYm8yqYLVF/6MABQE+/VsG
G2NPfXbqMlFwg9ioc+Qvb4xI49+tpIXIlqiWtrPl6tFZ4sSQobmaExxxQPrHEwZu
V2/31d6lcYcMtQPRbICf1VK0qZkbbAY9UbSEihvVosFVy7pVAWC35CGRFKEb9q8N
vWjUW4ydqVHLdmFgfHH+8nBNnG5zFZytFPn3gIfHcL4Edb+WhpScvHZKAhpOKfXj
4GFarKm2QuW5/G2wdYoYN7nFf9PKXIyOpl2euZAwy3+IITY0ik2aOTD0KK5f0kto
qSo8ef4Jdt/lgQUMw1vuojwdZ6VVkzjjKegV0FkjI8i+fgF5YhGrL1PLWnyyqlnc
8cgSAtRCy8lnFhJ6MvNoo4vkTIF6jHj/d66FOBFvoqom0FNAbWJ2d6EdhWrftHir
jovubuMdiySEFwdMjV0nK0Uhv/Bgk31ABPzwAcE7I0SfoRHrPbMyRaldiWess6wb
PieDwQ7n4bF95nU9RVZCXfQUzI9dy7mLrHyW43nN/up8nT7BKvIZKbcAawFPnSjD
WbRRsnjwsZdPHMHjErQzMvDfTY6e/MzptMB6aQOZ/rnzrqRvlnmsAE6unqEnMQiP
XVnFBeWCtQxrWdWIX0rlGkhXIsTxVuNU28Z1N+Eyim+60BgPbncQPX+n6CPfWeOv
CEBmfJABWB5FXRAIbweUxm3x5JbQwud2nJmOv4OwAxXO2EWXvwDDJAQuL2v4lyue
BdeKtZuWhnxA9uI9vejgfOfNmJHQrQKXJOeD9EZwSEW+Za+ng77qzsYr48n+tvUI
brUDd0vbPkoPzJCh2sOMYcija3eNlRrcS1W77AHNXeP/QrYt4r4N+jU2X+zbiWn0
Dq42tZIHf3aNlcJpxAKmzkBoo77B3HgTFTmGDxDgbrtlO+kZUmImSrSAJelAnDkv
qGhI0b68+voPxmVyDE3Ht1iDmyUEfTR89rBECabqw4ZiVTAwpl4VRic7XoyzH+Yy
ruvGzYORSeuEHc01xesIj4t22/4JIs4h4gCM2jAJ9RJaCEZu39HTYmIypGiJYzYu
1b6TZpiqsUHuI0EHKN4IQbQZ7RvUiOO416BbuDEZ/g4qS6JCajibLSLfp9MX4A+I
6btKhQTvA2t5qtbiWvzddxVGVDzQ3NJJ8B4TVpeCBgwp+1ZjF5XKa4F5oXZqyEXE
SE0/JLJi5n7HrtWcdG1Auf9UqIElVkaqtn2OHeBfu4arj3s1P/SVBuxfbi3GNYIA
O90RrpqGbyGGeaX3J3EdDd4HMfKYJamVBwqhl/ufEZSPR6i0cH2XQjohH/xyxsdW
mUtM7s3U/hAD7kP8vE6jod+EUd+lSJBrgfFWVRKW3cvkEjcEQHtT/+1gSMWECdzU
hstMdss+Hb9vnGPYeZe+y1Cfh2o78pbOcnVjzLXuaFJ2NY37+ER3sChFqBRPO1J3
6TejSyMVK06qqWlK6pq9I5bRnrUTuTDdSOh0thcNNKOHdUMRkjqgQkGRBVsUnBCI
OkHCc+seNungk1C8Ed3NsltTiHMhQZ5UQCfTWw3qZxgWlSBNIhDKG4/dL7e1PSbM
U0OBufU0HddOK1DJpEx+C5hsVFZK9LL6ltvvCQhZR6k5qMfXFNCfGki+9zkHbXLn
VffuWZa4vkXopJxXZ7AyHAfj50YuIlOKt93jfAA4RKdumroJ2u3v4ercCutaXsBF
WsS7vjNKwgex02e4Va/wl6gH8Ge0L2/pd7gwPyWPeUqlPxVEbseOkmgzBy3YorSv
Gk1ZROEbEARPudHjwoY1xF6xMvFHogUXYWMyn0dNEyehbCC4lU3aizhFMLZf7lo0
Y2ctR9Wax7QPPtQ058EcySu9gNwBDL3OefOvVPsgWKfD7aca2LrnPUF9630Ftfz2
aiFVOkG4pAQaLPJtdRqaLC/PojlzSZ7RJBf9Rsb4fPqCCATsx16OHFwBQoJr6x0D
srEw5jWhBvT78kIk+tIOXUnRTfMqNGWIAcINPK46jRTqkhIcCDKDUZgg7zQ099JW
u8W6z95Z08gUP7aYtNUmp9bBv1Z29TCX4HumV+XNGNv7BzMamlmBKbz5ejxTi5pj
w0gAcOr+GaGXr7YgZP0j2AHqawly0OjE2jqQMYkbgfq6SnhcARNxyk1LuYK9f0f2
S+QAgP0dOWcPcEQh8qGY3+yCktPh8fpWHygDFU9+/mzF2hu3NbCuJ4k+CZ6hCbSY
faKYJdOKQuQVlD0GHwcQES+iYENvrApNfjJsGPOqfIqa9/PSJD9ftZ8/kfQLldoZ
Bfyn2jHC5IRDNbOky28vp7Z/mMqymX4sklPpdNq5bR169WQ1acowzykPFLiDqcK4
RNtOA/UkZQP8bp+1mWulS95cTXDaHrNyoCouceLOcFsdlJMzmCLPHtN1f0DY4Uef
XOmfld4IcyrhHYGCAGPvDuJ0j4l6b+bERi6ySmwOuBtUWOLDugXNjQ3btRPy3Sd+
sYqCTZtiWtI7JYzGzUMYSW5kCHplHquMZQdQo8MbKjUA+SoyOkPPVdaPuSLsf+J8
mjSebpafVdxy524SyglHERCKlHCVensGb3Z2y2KLRCskUj8nOaWucrDWLZt4IzFI
PUGL8hLcrgl7/zwH50p2zxZALxsmAh3NmTSy2Ul5S6PMGYdm7wWVV94app1i1CuZ
bR4ove8kHMXvoRTpB1Fv5mqItqO1+6wryKj6khD64hQXYLH95f441vblEPj3aWe6
LkQt/JZUcdQr7rvKR8P4k6NqVmpbur0sWCibsaS0CLUwmA6c+zUdjBxQMaWVdmYC
ooTxr65UpTWQYGuznUMpvXaTTaNqr6GY1DC41JiUc6Cyzb+yLnkM1BZAc/HrjsLt
8VXn14072zI5119UwWNMEetVtTDRd6aNTSjPTl7n1IWvA1GTP4QWHD1LR5684iK1
WvdFReMQ+7nEZoK3QbV5tedCKvoyzqAlsJbbUhBDV2tDH6uhvXAyLbGOtYNv8Gz8
o8/4+Q/XHKMIVS2WXPAhW+UYO3xzqGaujbhnyFabAeAoFC4yKA88oYL6aCh8UFbY
w6aOGYJznf6iSjgwAYRBWA0iouGN7Lu6NrhyH52gvvEvv9Ghs72gEtJWUsGPg+MA
gmuZqPC7I/JoD3aQeEqnc4M0QEg3PfxWljNpNCbFD1tfqWXgCZMaTPfr3ONhv5u4
Ay52GlUDF/lMlQQh/UjqLxJtQfd9AwEluWja+joftLpHDOTqJvsxqfvU072d4PRM
O0rvt3e7WwEJNqwZ41e3B1h/vLjpVUrV16uvx+yg6SzM2mhmAPYbHb192TVZTC4j
DjS4LJ5dK0yekIEreg2gwqigSH2odsYVneSiPl+/U36mjiRk1i8qRbEtwlB9/o/S
Y8jaViD1Kh1H/3YIe9FQJtMd3cyflhnEsqYkTOSF1WvQocfVSQEJA7nIVc019XM9
uxpDL9AGCK7Gc5nOGx10rOz4f1oprGewCet2XUah5y6OlI8NJOZ9Negl+oG2SZn7
6ZHP2MP+17o5Zm/8eCykwtrn7yv5IRnhLzIWorafjmq2xjy2twotABBSOGmgZJJ4
+TfcuKAm+Ht2+4UFWh+HenXz/8n1RBVd/rDC/CZ32UYxbA4lyGNlzUT+8gKludla
sIP79bmHoG2CTMJu/vhXHPISv4kr6xNraJqO/U0Rj/YqCElu8RgnCCkx/TeOgorJ
Wg51RtMFYS9DRkzggwny/i3jzW+bLzGrgjnlolnK5alyKGoJ8u1njohWSRo0d9ea
wsuJxtYGM9M/8Z64PLtXKPC+BEJO/zjei8Daggk2WGAaWsfz8ZOjSiF7oQ6EGnUm
mW1mGGAMyQArDUeBkSj7N53VuZCWuBEpYKfFy+eIPDU7rtG3moZO+dyij3vu3syb
4sCRSJdgS33JOXdKBz61tD7/CFzzNvU+BllCr3Xx2SiMSyNUV2u4UwUyK8VKkkyR
BVTQIp9BRyJ4H009I9a5w5hv8tdS024q07QGN9Q35tTeQEpfM6n6mBE1CbeMNfXB
xOIkiAA8HXDXd1Utl++PfZBBg3twPwm0UEtlxM37yfBrHQmbkcGLjEXyS+8KIH1V
d6Z0dL3R+BoGX+iV+/SMDnJJZN5kFKco43jmVJ8XVkvnF9efjY+dmmagKKaBlITi
T423b4T9JSeUjHl+XD9rBu3ZWUMNzLCRE6M7YiF//fbIQ3ZVU53l8pk9Vu5Kary1
I5ENh5L+8cFAW27yhrL1Opvvc6eBRSR53awZ2jpDhusIiADg8tEWxPBjmGM2cy4X
WocigCOarZP/4ju/rFa031ulFKXrVm/TvJUJE1hbqkEPfeF+3suyobkhOZZQ5tZC
+a5j0TwhY/bYccMle+OSMbtl/67BTVRhWBXOUzAZNqPumixgdi6SWlgiPKSBtJre
PLNsXY6rIIebv2UeQ9R60OSPpnbvJzupMXxbVkZrbiIVfCRA/Z9bG/qsOkSyys0c
rNa9KH1NWaKQ3d5RVyxPGGmapFwgwxATlC5997W+EbUjDX4kI0O6ulwY6KUhsW20
Z8npovyEGbDIFqrC3M4TptlRuRgOz+FPeIvpg/8ET1pzS4DVb89g40b6zfa/5eoW
izTmiGT3fsqIlkJjFsZ+k72P0eNfO38IQYvcCkHnZprTLng1FIn2YH1IRFpSpAl0
ohIzzN6qYBOTDU1gEgvw7jt4RF8kH8rkHmuyE1Wt7+UJeA82qjyjFs/r2De2H1Pk
kimK0XJX8shop5AQ4ebsLCk6h8v13bzOe9s/piZ5ZuBpoDKYnOQBcBYH+e+eNAIi
v3ZuGwtJ6wSzhsSSCdFAeKno9N7MZ4djYdsbW0ohbkSR/WZ1rvdRe37rWdIlVUH8
igdw7fJFz+YZz9SklHM58sdTMIA8sYzImh+E8dMeWczbcJCR5J33nZN8tf4BVEPx
qt1/c3oB+kqADge/REXL5S0RGruFJ92GCvSicvfjuKQnzuB8V/uNOguI9bvV8A6A
QNq9g3UygvHSt1MCmjneWlbsQZtNEw9UA+dSAwcTgtNBYw+baPVZaz47XuUpgy2b
8bIxsqMoxUEsET2H7r5GcxkWQq0ziKGiNzBIfIyT1RFPUunlL4BoQaR8EPx5FQQZ
HdiFFtdnjnVtUKjD4pCfQkuOzIiIB5uG9eJhdT5yceopr2XzohpKGbmefswwGCNb
/myUiirZjM56HEDJTSNVqchEDzbhxWNLEtGYXJpjMUUvugLa6tqXgFse/eCLVqMz
RJvqMJglcYTOijg6py8WosPjsBLlFkmKF7TQDmAXhWYhpPw8Ok7q4o4xgd0QWEtD
BSrmzctKTGBgdN/15CuaP8wIMz1UXsxCZ+9Xc3J+i3qbz1k5LuI0YInSGtVmikva
z97FCEd5m6ebWEnMGsqEf13cEjBwVbN6uJCZN7KhuVBgtM0LX99ClGiz6wt2mGIA
iPX+nFRCGW8KeM+bU6u7PpJG8Cg4fG6qe5JgEWKSk9kGQVEdl34dc1OClCHvUp4/
FbJLfYaOsbmU/HeX+M66hgO+3BBRUHpqoCCBoI/EsBMmw8sftCVHsF8nDvCdBpEc
NJbIqCO9/fWnVujvaE6jnlITLkbOwsYMGX/F1mUALvJeYVXpyHrHEHJ1FOJnrS00
xhLqkiXotCWwtz+q2C68Y5hXD+Lw6eLunm20qV6GgT42xS1hEO0Zg9SOs/g77xt2
hY7UwtKc/5M6dTAlhxFKinNkcD59EezY8/uJHgVoNmjIcac7j3b8KNf9tOmm2Wry
Hiz2SfPVtFUce+ETsKWLgAz1prqAKZtnDKfl3QoqCZ08sVEqCMT17PYsxSgWs5EF
/yOoN5VQEg2TznuBABY1Pkx6hfhZBcpQXwBjc85WlZQ1iL3SGHUMPC7AA6kPLD96
IKnooRtaU1x1O7bvJUmISFI/xezzz3ZqYiM/w+ByrKLEtfsnpEumZtfwU6KcG4Jv
4pi0WRG5skgx7VnmlnuKrBZo20N2ZvZfafcMwUpeClbdnmsOmp2KqKEt0aW6kO8D
OlLzzVKqRYuwULtSnSB10+uhbO5UkUdnGYCAHHzNlgoFVDBSV+EN0du+VLjzYFP8
7HRvpJnS9J1+k6Bu6tVjyTIRcEOtiEBF6AteNLiZn4FLjuMLIspBfce0XtMs7XEh
iYG8NwzIhAC6i+L3+hjjxRiGrfUN2vmzdMtMoHnaR1kjK++i8xvdywGMveUCTlyA
r1o0XAS1BJBlsLdBIF2/B2LvYLwfc7KJDibvMtmWID/G39JL/U4CPqTpf9Bc8Sx7
fRxcuJ0DwzGpeQumFCo2JLZQsGDNkl416KmqNWzj2RsfJCDp1D8kLdzGa+zB8wsy
HNKWBqvpckOkrz+rmkxj186SHLLDx0/0MQgOTIXwASiEbu44aLmf5VZDE9XOk3Jn
eWvZwPeK+EhT3iC6fNqu4esAXAbElfZZT79JNUhJ4Yyk8ZcL0lcAgsaNMUk2C7rX
JTwQSJFbm+120KB+ArXVXnQDl/443goM5/UjiQLtqV32x7oqtS76sGRyyF91HPnY
dqeLCYcHluo8vnNcreoiihK51hQfJ/rPq0WgHeKX+PidH7A0sbVvAUpFUqZt78Yq
+pKWORtNuZ594XcgHnMfBxhAueuPGglKbPwpZe8OcvC3tsQ5vPjTY4H8y1Up1hfy
tJUd1Hhyw8dLVtnavM4jtO8R8FdfJeQgS2vAGCgEZx6taf7nEOF7ZPgY6Lt+Pv3J
VpLyDJtoAEdYb3qzXYwor7V2kqiOwuEF5VD9wYdNwxQgagzdtKAtoEKfYkfvnFuv
S0UzJWy4oNH8+rvbGoGcceCVL7lXRz3mqwcsijFyCxp+rBxjsAvBZBTRhaAie4Y/
46jZhTX880O9ibX7OkI+fV+TCxlShoufvhTvyBsuoDu76ztEw+SdQw56gs9OwUDP
5T05FXbV+5KqxPrS58ewZXe9IR03A6kGoIuU8wgFj/lJalVh1crAdcy273MJzo54
TKG5wHMcM7hMUCBKQau9pW1OI8MoxZHUkWSjoKyt5OPOkDroyaA/BqNoMubcW9XU
L1odxpFSN/bmalWeXV7oeJN68S9fkR6owov9809RYOAY3M73AHs2sMeHmFX9zVIw
jqkpO4wOJJDKChA4FPjZzdBqiFNCty1oFKeZdUS2Bw1UEfuyI48MXF2iErN/cZC2
4mbWPrVwBM9q3kagTyYEa3jwHwUFjsa9CkHDp975COsVkZ2hXYyZkV77K7KEOfSP
I1nh9tOK6CzdFKB0rVPoZ2+RfUs9UTKOjYpNiSmFCxJfHi4/bjKYPno1hcKiQrFX
LjpRa3oMZFd9uqrpQFIi4XHIeDATobmzERUsMmKDSU7dIJKyddKbuXBWJd2XaOTO
MUnyGGu5P45GA+MyDRHv0l45FHGA2HvQyAd4falDZ4SYYX1MGmY3ApEMbldoY1D8
3cgXWvA5mp336+6pDYQ0pAo+VQ8Af8PCxf2GboTKv05fyMOhceuJt7bIramw7Icg
jzaF9AH/jxI+wJqeMiCqRJuCa8oAtrbZFEXCoqMUg6sghSIbTgetsiCTUQXdhWqv
shfeKJWBzKmgR9ZgofkyOE7Jjm+257PkcYseSE/kanlUx7blIiFITfXJXIK0cXZ9
CxEgKGUH/BcXOPx7rgnYiP/4ys5B7XkKyhkOlHk2hA1CJ5SQcWrdfytbPWZVpE34
g4Ll0fZBjeNrhDpYhRV/NpvQ3J/hBEfc+ULMO9zEZhbZwpNuhyapk8aLHhJksarX
jg5KQkFaP6l3VhFqZaaRgq9arIhVdnaWBVMsoJloS0nxWKKprPsy3TdCEp/NF4Ct
CvYayT5TsjEec0jvWKPIBN/KSfT7nxN5NhDJFJ8WCX4aBWFPOwL61sGBBgqrWB8P
yV5btsVZfHRM2/TH/ESXwHZOA5Bgb6RxOPe+Mhpp2daTb99iK/ji10/A74ZwFcMQ
lSVRaH0+wLkwdMcXvsAxnETaTf3pN6xnnqszjIPoM90Cj/ABDmc1wvFGP7DwH3Zo
MYqdCt5kI8S27tBEDIhzpCUkGVqoWGQOxO7oMhDBpmzSDHhWbNX/k+aYfnNfQ7Az
nzPaTLt0yWm7uw8h0zi8brzgSQkld7LuHUZcrD0HZts/HTdCLRu/k6KPokzkHjzl
vPcXxViG6dA/Z2jZVTCdADvFUhAfuGL2/8640C/FLJenSpyjugzK80jhZVXbuOCh
I3Jq/2C1RrkAR3WlCr904FOvghA9VITHVgOPgKLCxEWo63zp3CNB55QgtmKq73zi
ol/acqz1fSZ0+Tf+zTnl8EJKRdrFFq5DAMwws7QBraNAJGBIrIzUMTPBl4ZPfPbA
+JNpGmm5TLvf3VHAgytkDespmfB6wJG9XYM6lXBAQST1uxdFUhAKo8Z5F6f2Youh
45edjx1vmNVVCkrg6goaP+M55kF56TRN0pyCibYpnP+w+4JpQFnl5Hshxd+WDAVx
Ul1uXPgm/MxT0IH7tkNVmlyr0wsbQ0RIqs10+1U7R7uR3P4oG1GmnnUbiVGNHFLq
k+9kzq5c7TlV491KYPQse5jClTcvDTn85HcpInHg6nE03ebCZpb415vWwH3t6hjF
LuL4mQhf3wMl19S3/FkpfONdA2pXZVtkAD7uDIrU/FPcfEBQtz4Ds2jOilw7mL25
ldWHQ4yEYyMpBZTNe5/cMruJappR4Ry9ikg2ROp7edcPYv465JqkupinV9jBBIIY
JjUOE44aCRdkshEx7jiqUnSpJ0DjPtgW2ZFR701FiadU+PDvBlWFloaUAP0MdnV4
yPfFnqTYbtqKouyPr7LeXjjn5wp7x1R3xIuI1j6hRd2VmG1G269nEzRKkE9tRdBU
2mnEwLDBSTCLgr+J3tP86O4RDi9QKw7UZZW0I7HsF5bYbcZtmw8l83AyaUayd+xX
eDTM3YTZXnp5B0+psNEXrh817d8M1cKYJ3jhiYoUfDfI7/WPAV9/yfoRU3lch4oj
OFTmP0g8MOyQOcVCHxX3XyMvBS2hccPL0tJpCJ5VAYEF5xjgSroDZcvEEBGSVImD
Jt+lDtWclCcx7F5NxhspuNF1A/lrqGR+KiRMp+YffmslmJF0lH7se9V1DL32t3aC
tBUXKTFdzh6MszeymYO6UOq2NNGguX+tfiH3Bco0tzN5l8MkiNKc0IjHxgN5mPEq
+4XXEQP+Qqc474B/kttRUYf6X6nJPr4uDEF5ZETtPZD18Q56bzOcTA06rtiaLqTY
b7W/Ekii58EuchIk6EhxzdGJ/tq/G460/Xa+KBbT+dBJeiJH9Sf2nwqqfcDvYKdb
lF7fNJn45nDmS5cYYhGgSwGsfszqAtLFLwT9qfqzztnyH+8l8Jt/ifIMALFx03Ks
7sX59VXx8apupNULzlIrijhhSmQE28+hAk8tSv5FjcKOkrnH8yavCn0+9/P053lt
UhQgRRRG3A5fVfIEd0TwY7tKo0Vls9gKYv7IlftGIzt/U8+hYTEUpF+aALw8vLut
BmvRuMQC7t2l5uoLTnKNNFs5PX+7gXarlI53Tj9xM8gD1ra9dCjWz9bpJjlFSmJy
cNzCcWGYWVTG9/cnwg02UlMFid43tW0oEljCu6XCHYXZkqEAylQaT+ceEJj5wplQ
0BfQ5ZXXiOnBzvyF+86GcDlwpG+wVupypmsldT7fa4210usK+WpT35W/ATF/fUi7
badfvtvvDbyXGMUVdLws1Uaf9zbwkzWazKiVdIgwv0jE7v/RNfXmbh5EqxKkibCG
ULcbL1pdbxGlrWZ/p65m+YG5DYuOFtnEi7W/UD5buChek97pEOxYk+CP9zUuoKGw
lGMANy8U2JA1o74J5kUX/8nEfC69CGz9eX0Kjw+g/iplZar8eT5S8uD6ertXTczf
gU2exTURqfSNsIoQrQ2cUPfgWwlVyugrHYlCKX63FhKt2tqvMs3bwh1qqlV6js9d
0+hmmGG86rz+cjqKiLBwpnBSuNEtNVlW3B/Rx3R67UcDJLCSvFtQs77H0CPJ3fKZ
AIg3L6olcJVkhWhiKolLS/yEUfCXQnqWwDMdOPyXBK1pBO37fsWjgWyKvWTVEcwj
GLs8GKveU/MmH4ZOu2GpdFA0MyqPAw28GwN+3ykFC1Ax4bjZFwenb0Fww0SEZTgF
rzw65JtIXO+NYvvuaOb95hdWjfSbyZpjbOdQqtOJnnDWiIfGTQxOyPfw1TQq4BDw
6vhRm31igIYFrUXGlbfyi8WJr5SIuwmQvNvG1vaGRibqMvzWw0as6aX/RlXFDgtF
8atOG50wkaYuvhmsPyhYUJzO8THn8FnZVU6NpudF6J6SvQJhFVN8U4tTP8zDQWi3
aqboH1IyrlX68ehN39VW5y47B5ZZFd5ZJFht1+y6bmEmwH439/mNS0hwF66aLmH6
D6o5K1KPO8Ym5FN+aV873YnDumB8ttSrxaHjQpJSpZ2WinfqplMfi2FsdbLifWuM
vns8o1n8Zqy3J6dP1JKE64EK+1TR38EpqyGLAtKN0cIXYAfE0gMjB2mPRfQg/FIp
keNs1F7qC2joXGDpJs/Y6GKoBlGB0bQmjCLPju4unZ6xCm5UkiymoyRFqxsdbOKp
Q13ux34xE0g9bNMQYvh3S+GPnTi9uJbQYqleQz2uJQ7X6mSnjRlAcIrFK6Xdg3qs
gXZRiq5dUg3WBXj9SvZISPIN/WVfoNgKKM8L+3KANv3ZyBOtF9R2RDfV8+MByqqW
kaWQSZs9QPfEOW8UgHgpJGUVZ6/N7btlYWW331Tln3M4G16Di8wQ7/DDVhky8Akv
Dv0iru0pNmcw+KCbEreCxuY9Hl8bQplKeG4q/jsK+EAI8s/rKH6gzCZpnvDH8nud
+G7IQtlqLCq2NkOFRxxM+FSZpEDHDISMnpwQ1rkkTd1S2pjBxdtDFd3xf7l2JSsi
exjliJwU6HYqppm7H13uFp6tG/HACAaHsS799A2bgTBxLB1ZlMcWMEzn0RVU16w+
RHR2V5nOX+N4zT1L62kLVVxHCZ3wJKDrT4NISrwo0/TJHLYoNAptjNAfXLyrdkGM
hrY4SJ1wd4IxskJDu3C2rYe9ointftFnxp0btuZuleQOGlyHfhLqVXITDIwgFsKg
unGluGzvrg8VtZFdzTTlzs0Gt/Gpc+0WJZ9gwJ1DMysfZ467N0ZqrXma5R/4tB47
rOsx0pEwk0Ya55uAT3gJ0kbaggguD1fXARbGjxhPGPyZRCXYJjpF+VMrGsz1cpOl
V580YS2DaSZ2Or+UE0U4AzxaIkYZVaZVPzX5iolmsRuhC9TD17tmQO+RXVjhYF1e
/vk3VaNA0UuVBzTadR/LPC1NFbcA2ZjfwsPgOBS5718oDCO9B+uIgjATKtaKESW5
EgySpL9MyAsHcvg4b2ILnmvfuEFfXqVcWTMpBqxcBUVaq0PNIu7igZAo6SkZAXEW
ltn2031ifObbwpepZ6tSO2jiAvzib/UHCdZTYYLxPOW/exTeBBfD3xu6yz0Rmr2c
tvlAkbrj9aMvP6SfM+Y/e1g1Oh93EJYo8Dt7cyrr3e6T6r5r2chjFpCwAcXxFEMH
wQoF8lpqKPpYNkRWiBQuAPnZQR5OgS9PjrkDKA4dVnAfSSI/FxFpEUh3qQLwTGuO
aAjuir4NkttoOFo1sG8nDk/lyJoizSMLSxcl6fMiIQSa8rAoJHgVTOEVo52P68MG
2wWHxTy+6EWxhZq2RbqAcvGxzD37eBl8hD+LsWecxjpdP5N0R15Yj+CHXxR2KtJh
AotqPulit9lG7mhB02FAAv6WU50Up7FjX0tC7sDtm1W7ncyTz2q78X0mubwW/8qo
dffPxYbF72LP3ovLka28N4KZ6hrCEGTgO71tiro+i9m8+XtkSXY1y1DJfgsQUtKl
6Ks9j748U9JIr0yRQKcjfv7hkKdJxb/CNbKORoQjF+nzoDEFJfje4Y6X3WgLtxgg
EaaUFWBLYC4gK4SqR5ishxFRHbIYvZp09c1grbGOuTGiI8rhuh1w4B4YWw3dIGc8
xmjcTXORs5l8He912YQUloiQwYiItIrqYNnpOX0cUNouG+2y0rvSQHmQifd7MNW5
+YOQ9R1gPmzfOgs0oDos2xX7bh7QUcUqT5Rv8nj+UWnOkhUYYR5l9sPZLlCFWlmD
O4hAvzh9LNbBWeLBwIGpcocc6RPu88dorGcGnZIWgdb42lRhFPqjEWO6OpdzPU3o
NbvFu6S0UJQG4dKRIWEQ3ZcTpSEnsoyc5SBbOvOR4uZFa/p9JE3TEOv5ijZFEANR
sW+CAKrDqhRrkB8Uuh/Oss8h5ruOfO+njyLUlSyT6+T8NKozpyDCri3tlVEeMQYZ
FVOuHKJF9HqrEF9K8CnXkne4RLF+135onGDBgS0gtEOI8lxAI+QQm2U2nNdKiHyE
bQpNhRgn77Cvy4Rx8baNq+PDzCvFj1ooet85nam+oXSe/5qv1NA+y/ZLI3ZEG1Vf
nr3qBSjo1Z8o6uzgN9aWOWqYeT5wC05t4AIVlO36BTHkZ+UvpENDIfwWNLhh9ydH
jWd7QAZLNeztOLQF+xHwomte2lHlaCnseHnlTdQ9+INQHNb+DVRiwoYd42MDgNS8
kTfr9g6AljQW+9SI92mnH8mLIjmjbdhNEi540QHwiWl8+Ed0MpID3QjYwF7cjkrz
IAcla0pkW1+uw6QjtqThby0fMLdKNnch+NGJcyxaV7/h7HImrkjwXJiF1jWBwMI6
t5CqsTp/scTgHf4Q+hwW52db5aGOqew+RJYf+TragMxGv2lLIEIpssspFekr1APH
++EGHuw4pxjbUrcBWPfr4fpsAgF8FK0Wr8tSHsSqqX87NvgYG4eZCE6X/5A54AeA
2M43/qopx27PKIyKu76XC8OC8dYR8+FqR/9RK9nIhK/fMwCpawu6AT+pQcTgSMAf
j4NDsn9UshowZmSoYjzhOocGPEjThoqVYL65vbGaqx8d+CYLVdIemphBr2t3W9i2
hnWZ493HFdkY+mF99LSLURKFYDqrBUTu+fiak8Zavhc8ilaDQMVBdRgKCoY/OVeS
VR6qT84PehrCvLHRpdweojYpYjhgrYhwNFK8GQ4SG6BQSQf09jzeMDXSlD8F4CHM
8joQyhqqLSZ0c2oWzhbbFGXN8Jn1Iz6xI9y9w7k9pHN5WS18LdGtTxknWHkKFZJH
RIpAexUXRyxuwhl1M+M/bkELj5VWVcyKYydtFcTJC+3tT13PQRiOEBdN7YPAfX3H
BmAiU7VdUlp883bG26T4gwSFXlK6ZQ8zJQWvLVohED4vRawjx4Y5Jh1O0N+0m16S
gFvkVX3weLHqbS2htMIX0N28UbnvmvxSN75rT2lMeSFWR6RJX4ZhuERGlVDwzXkC
YVryL4SlHny5QUky1JgrPNo5pISl4eMWpAUoLPIPoALac+7bQv+ef8lGzX0UdxSJ
kolb76gYcbm0jtJe88G1uv/zt/ydjV0qhOLcoXxz67dl7ST7X31j/UtR7R2KQhPv
IsT8c0CFUDm2uiANKJkKk7um6EV3BYG+/xgK7l3FPHQPGLfrl46TriZ9N719ts6D
sigK0Tz+1S9WyStK0UxPgRMKT/M1JmY+syymQ3C2x5I88cvTKM711vTuuOyxn3uz
yUojIZZjLUtYMCJXrmMlvT3Vl/tTXLUG0woGMoXUoVXlJi7C0e97NwqXqu3oSdHx
Zk5jBd7CfB03+x2pZmJV2YBfzkIIQkN+z6Ppd7TgDIygn8UbNBF19djafvcFGUux
R1Q5vd0GiDCBUl6pxW5f/ih/nIMxSSOvADG8qqKtuE3ORgaCCkI1yl+/8JHeZBYz
R2pRP3znZWBo5k8PjERWYHQAUhoXsdERHCfqvMqLxmV86NNGRs2rSr5RHbV6L1/O
Tp8LV9iCgWoZulamEd3DfdpS5J9PK21a1En+GCwSMBR7g4XdlOnnkwHLdAosPdY8
bY53bALcpzaeeMWtMaIbaJBNmvH2UABKT3t07VOSvkIrCW63SRDiVttlBKP3LCd5
ZpOWUDXcT8aXw7CJijYcfsnw0I/XoPgMHY5pCL1QlMlX0A68CFOKpAhPzaQRlzoM
EmxxIj3HxHCLjbvI4rzM8Y7/4GjdvM+fw2RQAR8GyBUUBVL4kJxFCtS35EilXwjC
TjM9lHfiacob3AY7W3DvfedVzFG+WUtaPDSc6ZT6mo8HiXgEZvi/88ndFwiUC28I
PnykZDuzF5atrB1w4DtOqjTB6Tt7JjyChHDPiUzw+a0Pxo6LO47iKICRl2/8oDQx
DBMgO0RT1xG41MMVBzPsa4rXsPhD3NeZus+IyDOazdFYlysWh1/r0M4lyu1ArjhK
uUPCjAMBOjkx7nNaWO4HKN89IDXmlOlvrrKRNH/9owLT9K0CWtQ2r+QlCrh3aBKR
FyFRqRvSx/g7oKRAvvka+bmT5CkiBwfY2Ps1kUM/FxZ4LWHSdj1Ur+13hRgQg8iM
i4d7j8Vz5UF4zCZglBlAEdXpltIeU0jywQ+/YrOsXIwO8KNkC5F5oHfhJEZfLTkK
kphxLqE69b/j2asszzy1cM3dfdxpadMyS27FOlO7rD9cIxqA9rWWHLtAiov6BEXY
VsjR8a/T/E9ap3pydRVGa3erQ8tTwtLWaitAJA9Tuzks3v4CubikRDgEVLZg73PI
Rw53BGts5vD/I+m2EXWar45VNB5g9nItJW3rxniKE8f+XodZI+lPTXCVYMan6cbb
6GRiFUjFnyoIvVfRQ9iYMtVlpDIRGfkcZe0DYDqGg43U0yMGp4jcNtG6R3altd3Q
/Ry/mpj0qCo9Oa+FaGKgvbHXFJQuyIefLLCbl4zl88xPiSbmNCX+V/rYzcUO5lGu
I0+rIwB+cVHeqVXrKJABxvmH1Sr1lLRZJTt4kvmPJ0wMIYhv/ihVHpgnvkCT/iNA
Rf91ReXdGXsd1Un5fbucWQ9EekCGR+MvKmSEj9PWy6v52Lan+aU20llv6RYKRicI
DiAH+cqHtoXlb463h9zL7juLcr12Kt2SdgHJFw6FYdnil4PpiejQMbv1GKeQHnxn
ekvomgJFMvhMSRpK0T9lDdV8QcS6alQ5pwE4mwT2k0QLRrLVlK2r2J0inPiPBgZr
sTNnqiqZUKdEGkupHlHqufhuLeIZDvLMcNvJJcsIx+rhCadiKbUmk2EqtT7HJAmr
jHMOcd7pIbfJC7MAx6EtXCPiSRG6pFNAC6B7M770PYVnCtshwaMdKYJgAy9Oh+0C
Xs6+bnguAwIzPgkg6RL3iFFq2Dspfkuy4+euZBWClVNvFkaUbYc3Lq26cbF4ZFZU
V0MR9PsGzkPLGmZYDaPqZUgJvftKeQCcNtcRxoDKsIDsfxWpI/VbvLLVf8Y2I6BJ
JRwW6WAzu/Y1fkevxb9OT0NaECOG/BWOLJ6B0YqG4CJ5d3mMcn5jljSNwglONWPD
XXo4VCW6TVbMd5jxKUZvJn13BrDfhtwHkND26ZxCAMdDMijnZlCxlPG1YGY8+YKk
4xBv52Zm5X72OSI0j4DHigIkeO5LXZStdv8Dc+FnSMLb/6JJIQOisqjvS++AxtwO
mut41/IA5u6GXdyvaDa+mq2DOnOmGAQsgvfzESkTi5YX07DQ7jo1Nr/OcyNC1G6T
1xiq3ogw3Bafq2P6sokS9JsVptAhkjUlt/bRrJgx/5Y2sWmpZs5LiAUyN8eYXxU0
qjVUjLPIGSr5tx19zl8iAYwu4MeALPjuvLl+HKMfpOSVoUZQ2D1rnBHbh6Bx6z/h
pljgggd0EfeY8THLT4kycTwx55Rar6SLIMp8Mdjzk9urRG+9GNN7dv4x8kUiA4RP
X27OvmUvI/d0A5l7fsPGY1id7nbj44rZxxrIX+WZz1mjpOL0Wa0X31Lz9/2/25/z
as2Uv6esoxSA9DZ2qf4EuJodT1Aa0EtOg2u6gLbQzv5Ss+fgmSZ4Pi4G6t2L7jQ+
LIlba94BDW0GfdscOthhwKyMFBlQr4bMNgMCHepNrIoTQTDzRP/erWurLNleQguH
0H8syYL+UeeJW/hqR4wMaLE7A0mZzIjYoHvwsNXa0FFjGTEFn+zhVuduw0/3+8+k
zVNVy0ZpYqqkjYysRwh0KMTj9AvRR1EjYeyccApzgpYzJ5I4ios1vOxR9Du8IuuO
Mk2GjlplxjvOeg+MkCQavYG+oFWPTyfwQQGb5506v18O715LAcHqwnLPJb363DIA
YQePI6iiRtHHGeParu3aYYeAhRWBmfG4fT9XKIWLOl4ihR5SPp6/PuOE6Hw77eaA
aWJvw6Saocvr3SMHLqxZq19net1wttnLiJH3E918UfQWpLPVPhZOxpMrL2GuWXPV
XA0ygcG2Ym6kbfB75peSlKbUkuh4E+/fKBAQ9+zAb2U+N/zFRI/PowBQuUI1R0aF
J4ws67Ock3QpCoyMcv2PdMD8FFE2kBwaTCIpCueAty42dEeTLu/wf6+N9Fnjg97h
xBt4fj10zlGsHZStzsJhbqAO6A5i0BxWRobg6MszRJufUZ54vAvUR3g5kUb63Ruz
1mBZNmxUrMbghHxz64LtNbOEbCsPFY8629vPLUXBXOjax/7qzTkCwp0oxaec4qpz
XmdY2Zm2xPRYUOCD4b/p+c0v60GdSuP+8NMB5Z/pIXZk7939MUrI3L758OoMEyT9
+9X7KxG1T6CNyWZoJ9Z9IezYCStE9GlKLFvrzBrjr7L+BVyb44hVG5BbMvGr1Pyc
xdDBPG2+Q6dVPq1/wBmDchHOgWhcJFQbKLmvcf4rFZkyWrt9a2BVM1LvnejK3Hbd
H75cpH70Iohwr6u+wj9BTHOeyhozkXe6EPoz6sx0a89FtL84L4hZj0jPGf9hOz4W
FR9tk21NhJ6vcR4mLCBtOqYwgNenWFFMZqOlfCD3Mcfoor8CKnKdr22f67qTbFZM
x2MYeMOAsyip30UW5D0+EKabaa65cjH1+JOf3nwHEsp/6fbJriJWqs5O2+9CAVC/
FVHV6/iCCKT8ZwVeJdPGIgtD43S+qy8XbwILqqUXqYSw3rEFZtCDM6Hg7O9J1Xp0
5k9muzrV8jB73Ghs0F0cF7sbDVSe6Z6oIxoFBJC6pFtg+W18uOZT3ajVMyuWj8Os
FUSuaycxdqcAj8XbwZxs3UhhNvMv4klcUvhX3S0fKEn+j4BLB4NUDl6Sv6ooOnPx
PLCW9Tsn2aBtMCOPnR4n7x+gqBYXQm5JQNNkuu4qqQR4Ov6TmVzicSMABbFSqlOy
P9aKEACEF1e3NE444N+bzNSqg4kNMmV99pzX+TvpzuZfJrCbkgxwyP8SG1R3jcQB
4u3SC3Z+786HK+Ls+HmeEn+qHnpilJa6+5aBt1PrTFBIDmIOPFjHxWgN81TU/8QL
WLCmXPasRHXnrUAJS9MizQBiTHZ6kPiYTP7/sh4Ff1cnlv6uCGhLcwZwPxpIQoQ+
e3cGpNum80GwqtwpIOsYEMJANBYwot4dZp0ao+8L0mL9V2gj4gW2j2Dldyt66P3M
EJ7/7URQ30GVRBRzy6Jr++EYTnVV9T+f+FyzFTkLtUXnWlWwwyvJ3dKfua/ox5WH
ShJjlJqjfh+vh4/Evyt/aUWh0TFoMklHPOScfRlOaLlL81rbxJT3vmLJXoYryUW4
zPh0I5ZFlpA9GZKAxKHBhtVRil7OAjkoFXchfb1ryJpMhOPwHORJfm+GJrq75UnB
QKEOBuWfuUERcRD1/XuXU7KMV05/CJdLnEklu4JYmmS6QUONByQTJq82vAnmdm7r
pyPRxm8Es5ga5cKJpTypy48STbsnEeJIx8/94NpQUgiqsjQr/qVtroFAJcxInlr+
KhdsCXhYF+4LZrhbyZmAlllQIgpYvhjuysFehfz4i93MXo9ieFzZAIdENT57SBZR
A1lJwZ5sWe7e7OIVFhmM+TMSXAUNb+6f+1V9qrvN62bF580DIxCPsEYLVnf4rr56
h076LE+RjxB26JxgZ0D2FhGqMDGaoSi52HPbsDgFDjQvLf+ApjwnEyBmhhD2A9Ty
AjC9geU+0DPo8QQJKTjtxjujCuyH0u3ForJOlcXSaDMK3KotBZp8ahaXcIHnjkLf
1UChwDWR5IOuuZlNvQ3puGdlO2EKsXyRVVgOMHZJqvviehyOkrGbhjZsSXYF6ZB0
n4reMwgPBxvDVxhoC08wExwT6lbzcjYQCq5ASOuovBc2NCsBygfo25Z5mtOMm3jy
jTXiel7vCNM2SLEK6qiniV26Phd5akU+gXQR3P02YLhPi94l7iEV7uF4FGeE1pmg
h03+pvuJI5aRDYhPazKSDk/fS68QNAwPiTCLPxOyWB1pKdsM18usNjEkQQz5Q+Wa
N+g2sO/ZqxFJ0mbh9O/VpshzpWUkik5jKabfkuVB/vBpshu2ww4WaCyjyLpeOcTq
TVMGoPBinN684dlNvkfSLE7nc6aZiGPaHhag6VY0uq3BUzdWR/sj3fDxUXQHuQQT
r69zw6JrSySM+2dmA3FV7ofjF2z84fCQFNiG0q7fnQZEUQ3Mw9xC+2xrFPdhpXFl
4/iFn81qPpS4DYuohplokTBdE88RR/iIsmfQ/3gLpMBCqKxR8rKsGRgSjuRoL//j
CpOqa6ywSfU/dKwKZcBcG56z/XjWuCRT2U15ewDUCWdMDmlSdD+B1S1DQuhCriIJ
x/iy3NxNweV0hOCNFsVMfaYOuPVEEAs3fDESpVSaWuyaJgazwV+BSvmntg9XCWAp
5km1OKD49Oo6P+6CZhluRnQ22QIKGUgX+Qah0IaKaIsw1AgqV88But717zige+j0
E/lVkc0e8CSefHzQaU7lIiM7udaNxegx9/xH1EvqUNA0JOOWRdGU+b/Qs8lRiOKk
DXZCV5UQAjhyjM7IbDnmG/xC7f1Yz5k+NIPYZ/VRjG/RBSKOfSa/Lq/SejLgpnwH
s+UW8eStLxptonCv2dO/Sz9bN/IUxIu8nH4Qca+cj1VfEWaV53nJOSUHuFBpeuDb
4ijRD2geKlW1HIK3GabFU+dseJ+9ot8m5Iflc8OytgyYvkKNx4JkjnzhdZzhDvSr
FVzVtNUuITKNbhCdhMDjsAmc/7vr/frVu9gYfZowCJQvLRSfKx8KFgHCWL/l037R
rPmdX+OCJ25Fs705IQuY4i8YRHxb2V9LYxOXAYPhsWbNHQLyVsXUQ8wWBH/uDJA/
iPOehWFTPZuL+dXBlmyK/pAXbxhKe6h6Vq5g/1tu1mQcKgKD1Es2SvI/GcuIO6Sx
96QYEq8mHc3Qn0q4JXX8Orari8LXmTtD74/eo2zjOTsUURF2Utv87m9BQ8pyHLdd
a9Hi9US4mzYB47fZTlMPHBfPJbiybEKJJ7b9dg5E6lZHLNx5R1TteYhcAoVdWfn0
Z7ddfCJodhouPei6cp6qtpiiVQrlBSCE8Md9q/yGqYvLD/z9DaxSq3RhFvhX7CWF
+O2tweZGcFjGaAyrjQriQBl4R2xNSaJgeROcQTbnhEVYrlYRCpiBiQqEGZUuFUXp
AqSSzmiHEGkehyoKnSLE03Cqt1io3K3ji6xziDCSEGfKzCUE+BIkkCea36PpsLv6
X0/AMbBR76p+BjlN96L6s76a6+/MxBUJsNm7wERX6V8h4ekriOK1h5/ZbYn5YbsA
2DYBSuMotDmvUg1RIVK5PyBxRstlp4GGzoeJDWCoggTzyAP6QeINWZM2HMP47BYG
IrjeG9mG4xYXBC3h7fVtT/EHXsngYs8u2ekVohSD9GObHjjeOad8Iesn6WCO4Jc8
HdNwB2Pv6x230Ek4Q4KSUpBfwjbQ9Nu16rzZJvOobrmhk45Nu5uOSzppp1mBE7CO
72c+b+L/zl7aa7BeYP8ZSUGYh74Aadho4hmv967cle9b97W1TZDgHlti0+KomwCt
CBv1GeUMnOcMMpQnTmM0vmHXafHOnhsOEnlCG0f8QnYtzo4Wo3MtNIWlxPpiegP/
XPjkV6vqkrzO3feXHeuZq4MVAt0nAW//CnVh61WLoCCAJ9zTzrr046rBVa4Z6HNj
SJmOzPwGlN3UCX05K4Pk9R4SOt8+QRRimVHGleFKHnnnueCWRTUzJjaQNNkjs46q
x6gKAVUI5zbDmFpCUxAnWCncy44nnNxAZUolGP5y4nHs/GKrOIZwhAzN+K+J/FAh
nl0VcsQ+PNvOTyW3Bg36GJovVIN7HhzF7h0+3fItnX1RE48ZkrhOhqZnwP/Fx+7k
F0pOVO0C94iO6gzmbJmE8v1XvgvJ26M9D/MzO7TlvPqUWp6Yn3NtS/QXCBVB0e9/
XG1nM+87Irj63DA1Dy67S8CVVUlE46kUfcBXU2Ryr1RFvt2zpd6CBNaMztl0rxmc
/X52F/OhyBPU/GZ+mqaQg1qTPQQWsjo/y1x74E5zwCnU4u7hXSa30chNk7GsgzMZ
nR8SuGT8OBsHqYPD6iBQfPslidCt/VcDI481Ghib6D6gyg2m4bKWp5GB/GKDjPA3
p5FWochxQGKh/NI5XK1aiu7cvTG/EoAsThPbry+NebMhec91Z6qZitnpIqts3+YJ
iLMWVDLGZGzPrIi4udlZmp4SMEWLieAvjQrHs56g8qeipJcBxJJ0g5qrp8RzX1eQ
7yU4A+vfNlwxrRtkS1ZrDLGKd2mCDSOng95qBIjulViIYrpeqLzXSZReWdclNGZS
7vNG9Rr5KA6I5lRq3Vx3NUIkEqK9aGqOaffRW/QXorxrNeiWlQHYguWzX6ABUEbC
TKduZmINHHr6vcQOvIiRnI0WhnovnkllCd/ZEIkawdlljG15oYa1odXQ5jrY7bR7
TXYBvCjAO46jLicLvTONpyekrDdakMtld5nt7/T/II6MFfxX4vMrv+GuOj14vEH1
+uGIvMY1umHR8hBbxjW/ZYIRsaHGek3nm7BNqIRfSWMaMghS1EbBImhwKFL6Km3V
OgS549TESPyJtJ43mP2VdmKCMzTu6fL7fgsm432HoHYZtujXeNXvJHd8HsNXjcwt
t864WkW2Qgaqfl41EH/aTNW66QIeXI3CbltHnmXKmCjgqAlk3Ki2Syo9h2l43JUL
7kWQ0IjY82yzgTOQH0hpMODFMLNMe2w7ecC+JoGNVP8wz589fyPb2wLdKn4PH0CC
38I7cNRzDD6llCyMacbqw0F/SluV5yL+fOrf3RHjSLk9vxCJm2KsC5Zb0/ETcrpd
PB9VB0htsntdhjzS5ainDrQSPFWckqIAlGgHHeJcPSnSJhuLnOpQJD0VCoAh7X6T
HUSQS5g8xcTMBZrHcbnXw/PGIWIpfD9XSGf9sf7vEKqdXhLvDiSVrZlVT7K0Z6Hx
wZA256Peq6hlO3azv2SbETIeP1VTgPPNn/wN0U7thQ7YhkHwtAUcn7vhlF1a2njN
zkhikxpcGQ+wC7g8R4sIEDK5vXZ9qj7B1yVemO+6cDSKwjL3w/JBYpfu11tKLVjL
cGD/BMYqxQQj7QHKpoj5pX+3s92XnHBhAcQDIKnbrEKRF0TrR+mpsaamrj2cmAat
TEk3jeUKpwpEahrYDwi12G8QmUUOxgxYc5zbljcU7gVMFXMyVQgG+Mx/3O/1AHAP
SJ00Kf/nRsrnxKM4ewSohvdZQnfc9abLshApmcM/in8QXZTxyiiZpHnZbBdihKCN
+9ZRiwWZXWxtTT6TJo85iC4+EsmhlL8VQQ/VSU16mPIj4+iM4Ggk9LQnG+KGcCD/
OAHSK3tNklgQp/U3uBMhjgispcqeCsGePgB72LbJDrFtFf2xtePaqUKauB1hoYyf
+se4ArYiQr6TBH4EN3RSfvJ8DdxnQpYWFtFjH6xXMbdGjYFTdBa2SFWvpJW1b+JH
rM8Nlt4I+AGQ0/kwZCijk2HRQr9kRXVokbOKs0C7XIFWPG6nlUVwRAGVfoNnk3d2
7mCNYXmKf8srkkGXHpIxdafYK134katQqav2MZRIMHy1a7B0rIA1R4bhSa0hSOvN
KeWgrAMzPlafKi7YCWvvVuFDbnZxGslvvLKh1kPk6+A14DShiq/oSR8XQwjVg/q6
JAam11POGyA/a7itKE+uxndIgf5FS75KSaeQ7tnxsgvQ237v3SiezWTg0SoCm0G1
k6KMDL65uuAl9ooXQsBoOv7ZgqFXLgl6cfYp4CWuZwWGpM9rFLgulDnvPexCUL+p
sNd3QnBckeOHCSrrYN+crkN1IQnrVRa9wM5CAWT+70rsZpQiPk2SNEQvO3Ay0AHs
aCM7FXPkDNa7qjdIAwiPxNWHH0Q++ah/WZ7pMU4P9uEZpyoo8bf+CVNrrvhyLXiF
kpKvEAoi7LeD9VqUBKatj0p8OJwMgrDFF0dp5rOqoiIRkzCWGcVgOXsagUPIv3Q2
CwCNKp8c6LXqXONTcMx7uh1m+bjbP9E+VY7FslwuW6ol1EpZeFGQsz7t/+qCK6W3
BpRqcaNZJxlzdVa4wULCKJaPCxCHV2ha1pvBv1HpqLLLfa1y44smo+1BbOpq7Fag
jolWKn9TGrQjNzyRez3rldt+SNPJOyFvEgxpy8v7tTOd0wAkCBdcdEZ3DyF5r184
SO72FyOF2LkccgGL+O6tlRDrFWgHrY5qhozGur+kx66GQ/psy7DOZpGl2Cbl7Ink
kgMrSG6l+UfgBCTpH5WjEYwRlwtJRkKM6NiBH8Z60urNhEY1ZPuYm1cQRF/ui2Mo
FYjPmWu7VKEeRp31yHUDB439JAjLca3Kv31/8RH/ev4qxqmhfr48cJByhFQ8VQlI
zwktHzE1Q8WsENNPn0DD4hwnoOSiFXlIXtxPStBgfxnCXmeHg3otzWF8oJLLXMaM
ws8fuGmD4Rg4yJAZZGZswAd7T0zbUyFuSr9Jvw7TmIaxauHJYkXUnbI+SJJUeWrz
UZTqyM09nPZf0MZlCytI7TsOZ3odRrskMAgnhP1fu6Jjzz1KHxPlL6RkwPZOYDl0
cVeS4yx7aCHfNqKDXjjAmjhf+h2B4+HOEkYFX4RkSscTgOGZEVlCWWeXaYb+ZAqN
ojjrpXyNfEWmCS/klf9BX/WDElxWSxLA9K50z43IzbtAmaf9GW51saiWOo2a8jgm
QMJTRgNbRe7ItKIREQi2BbM+l8+B5WndhkIv7E8MP8nZOspg1sNsvFp6bMpLuG7b
xfHXJziC+92S/y7U93y291yfC7kx/gDBqYLVggfJ3zOuwpx3683QMbRE5MeshU1C
sM046mP2qkEkQDZJHBRSVrm/9h2+FWk7VRVl5uU4nZ0XX2scLBcVQm/zvsdW+Uo/
QgMTnO5kghE+EVyN3RYGIXqerWl0IC3ICjnb7tXaondxe7HfQNog/y46sdCiGQkh
RaXCgSlPg+p+WbqsWOoRfkOyWFPgTsl1hM+/NCPY+RCcgR9/zWF9Lhw7lOcCXlpl
gwf/Xs8Ed1etwaWlmo0vNZcNl1yRp0ExZ3ZrqYTwHZZhLJ+wXYYPnmXStKL1mg6Z
FY1V+6UAediy1BUQCzR81cHP+tbCiD5gHvw4uPj+uu+xya4Xqvh9/8AI6vwUdurE
8p0CB+Y4tdMvLX3b+a5yRG2h1V45zJMHJU47LdVXjoUZafLQZS5x7orzHpcgmi0o
3FuHhN/Fzgnih8trqQXYeJU7adrM/Wu7DPGMZEDOcfH46ZIpdIH0HibNG5dHznv8
srBAMeuDkZYTbjLi4RHy4J+LOa1qgpJTFPsHo+D8oNXB+XCQBZnRqJ0nZPVcpI9X
LCgWq0H9L6qlVl7vpJPHGZPQfHvuvdOabA9DPQOA8q9IA5lB8mWNIB2h0lRCzJMu
Pmm7LGFrK9nTWyCd9lUFrlfLtfPcEwKkg1CU8Y8p1LMYFVF4+pJpgIfGD+aCYf57
5rF++XntV9evEkVu+5L1zk3yAxuCOi41VF8Xxr8XRt3xPdGzf38p1e5pXrAoFHXw
DgF166Im7ZWUQfV2HS3zcAxdwYpo3qcrrPjTXedAst6JDcvJnEtEl0HQG30K6D8V
0peBoG+0eltdibz7cfeg2u9/1kItaJOUGliMoJovB2wpHgdIjXmYloP/wUS2Aoa+
fXR5aOH49+zbHiACWyWB71mZ+JvA1oJUZvVuwOY6q9pnm94Gq09mKvM0xOMyKGD9
zG/GlNq53H8WQcjJ8f5QdWAUlxr9WCj9QXX7HB0PPn8jf94EBr15aoUQJZq6nyVf
vPCLH2tq60Yx8XlnU+yyBxlMyiuGlGhWwrdOenrFQBa4XzMWJh6HB42P3q7eV8aV
NtiLESU7/NpOQrF2y5qb1gD4sACrdITtHYdhb65qgZjT/b50R+Ko1SjRT6nrgYT5
Or/MPNgekkt+AtjP0eIKJeitIF9Du1qpiFiePvTGrWddLcCf7OQk02X5hnjOu+No
rIUgqDx3kUwP+l9IicBGRKQXBxhfZ9SgIsg2HlXMtY4jut585AyTLbUY2ahoW43G
qsrbiRIrzGOIjjMPl50kGdp7su248pYD7Wu7Z4I/QjBae+r9C5J3lZ5PhQkNj4AU
Fq8K2yT4xcGzu06+jPlCWmXUJdNYRaOHZt7xzJi0rIXQKZQIcKGNgq57O/1StiwN
v6XcITUEMp3N20eX4F4LfKLZnwvRUjtHXG1sTzCsg9jzx19r7TfddSnXiQJTfAOk
frfLIx9jVnuHnKzOaxIvMWGAdf+cAwq/p8HPOy6yU8/M1tKH3awzfOOkv5X4GqrA
FOUTxF2958MzHTLDZ0mPv4kiUbmF6Uoxyl0i6STkX3litaTV0J1ahvZL/E87As2m
P/xTrTIy14k4PBWbB3dtJPzbYEAvIA0MnLqvO/FuIHaeVVTG6TCBab9AJ4jmDf88
lvLOvTmKXghUl9wX70iDSud4bat+rWUEC2wbpUp90gjjkzkJE4AqDTUAmz7lvff+
DXBFnw4B8sU7+cFfbrnKTah/GvEYHzT/P50BkENMcvTDBBCGCfp894kPIRNwb0H3
PyQ9E2sO5rP7olm2QhoKxrM7KFJhdYnjzWgkOXd/ovdwYdKtlwXNj23myhE7zKzc
2Nbb8q4GzilU7wm8PqVG8dut8wVGD8JeIUC0M8CCnMF67V77G+sGZRl1uRW8zgqX
9/M0Y5HFpW53xG/k94xdEr5Jrgg36HOZXBwIGnZtHt4BI+YUs4Q8VzUbwMVMfvNZ
jvnFYMSyY9US+UMG9OfZtVCW814pYZr9O2AXWxxU92CFj5rYzKqx0DxftL3KtGvT
5ijMxbXcBBpeH5YSynoH9rji7UKSsAvtYKfEdREHJkq24PoDlT+GeJGTvv8GqqYu
o3evbIwRraJWnd5Ke+16yxNz9jfQaAUqxxUkvZCVl4AZBTYtURzGIDPZBMg5aVel
vJyqsg3tBSON+mFmCCwEijskXhlv8sCCZ7ul3gkrL13B73G3qzRcNyCUGT8reBCk
i7lBwlw2cQV6XdeWTtwqOpDhkvoLbaLF8q1AtHs0x97ZeVUyE43i0IR61zJEAYGa
8dOgGkQHnNdd4SzW+fLDD2q+EXZ85sBU1y6P3vCke6kVlW0tLtwweCWZKhuldA3o
qO+ptuM3Fwe+fE8LWVZynxdPhkfrWmeaXz6QlSQxvGOykUtfIPTLvUA9fWB8Lgny
dseMtQHeqvarwpVMJgoL88ukXo+YQXmP2ZImgrTwZqVbNHOAHiazTF0AkklKmUAC
MWvWwtAVJWBANON+9o+iYttwemfvjaNTjTebgtB2ZnrB9zQwpeygCnWfuZ+LlBTI
R+bwOR8Si5tGawONl8B1gVmIu6dalqgaK4bk4p5hM4iOB3Z4NpdxDBZuLUjrEMWC
wMKo3p+C6yW9hw3SGviFdcZM1ebtBGcxrEVcoNIMXjdj98HgaebvRLdhsdtAI3U4
QVSz/7UorctD7G9bBDWVseJ0knsr7h4ECgIXdKSVC125HX+m3OVO7Oi27fAtAPLq
N9821sZVlEJVzBmeE7Krj9ZjMu/ox2YQTvlQVvNXIR3b34raM6Wbdg0f+ujGU+5C
p+FpTgZzbaVpzUy5K04iOBan3loqmcSwk50bJvNENgJu/j8Qy1Cf1RN1tum1rslW
nkzIW3xuE26KGKbziJheO7PNFYSEWM7ZGocIgoF/5Y/K959SFG6gfb2g2IRQE2NI
sdk9nlSgQqKRUMMfyf9P6iK5m/uzygC/ORrDY96RPLvVsai9Ode4XjZoYzKWCkBK
itN/gg7CylORjPlGTbnMWVIvXyj+ubVYil5BnH+VXIyjxUhLEUNz0VFc0qrKNupY
fkbzQi0wmYpdm/JTdEJd/Nf5gYgDaGa4XF0WQWr8D0PICf87xk02HEMYjO8RYyJe
C2h3CwisRhdmuFWNwPKRhn4lfkLVcCkjHDaXpRVn05ri5ilLsRMpJtXQ3j8DJ9Ym
Cq9VytrTgmQ/IvpooEeEzlOXun7w0Q5W5/aXfIKc9QQXaZD+phbTE6PkpSABPTbQ
6b6WLXS0YytFxZUowiacNqMVfmONxvKqU7IMU5E6TVNSuVpovv/wcHINewqO87TR
hMIWT06w1ziYO8mc/g65tKsOGDHYhbWEIvgN+LqWQPm91ugq2BfWrO2Q4NsCOuC5
I8eWj6d6yTR3e+nn5t/iqrOoeT2KQW1fbiAjRXKu4uFZDVBhe5/vJmvznSAKu3I0
J9dzK2Oz8WScin/nUiPmrPIdNvLsql39bY/oHApOrSMuJcSrFuitY554Dzo+fc/y
UhlgmG8cdBF38dS4/mJ/sXz3R4q158YBhRTCtFdAc8klfnHqG/xmkSDY4N23yrnW
ZumW7jLo1QZG+6QquaT8jFTDmm+66EK0vx90t5V4/+4mNbpCbIa0NqAj3OZhqdXl
fAbMrpIvPTkBVYzFQImXkM7XXyEyat5ij5eDplSm8wM7yOeXz9TgS5mel0uOUoIO
2OAmoTmY9OzvdLau/m7lShcl1CMNBJ/W1czXUpLKiR4xIH271LNK0fairAT8FxXN
XH6pGaTMn8MmMOZig0+fkGYSSFjy2B1g9kHzpzVm3SB6mLyMt6zVBlqyzDcp9EkK
OSYSBZmILBM09d4Wx5+zdT5sOq9m9zKe3FUk6rCb/3PiebxVDuo3OVG3S/3lqHpI
G1AvyKUx0Hi+LjMTc8hL35s6UTHDTx/UKTE56ZCJhOUq+/jSir+SJsPykIx8LML4
I/Tgb/HcYga5mxyklf+YsjgsMng8x9momv019ffY54i76NBUnI0EQifJ8Hm4rxn8
Sn8H6zfB4+kngTTCRxRQc0F6oNQEjgMxxoBDRyLVsqk40vKiMV6vbCoL1PLWYXRK
m6zE6oLyKEdTxdGT/QQeZzV/H2apauMrtZX4Cgm6eUY9x/bGdMmsPaIrk08rb/QN
EBEiKs+W7YDrtzsQzCaGZjKThDPJohDLliVDJVq3/amh6UouOrebxFlDozS5cDnV
LOfQn9hx8Zytl4SRjcNvy7ljWSdGmOP4C9PZvxhEnx9SnTdqrgaXnWn6HA73n9en
kg21zQwTee2C3P3q9/dB+fL8mY82FcJqm17heMY2EoSrv2ifB21eqwTzDyCj8iow
58V0KrLLcMvHcZR3W9bkplWLYUf3xQbL+fMWbc9TaYAdBzJL0R8TB/6t1CeNqsIl
DL3uNek3sN/3J61PA7tedwBVV//OROT+DHgIDb40ixbZBmyRL68skCeKdq7MRmWQ
40CBFKHz28ffZUCnyIfBX5uFCBQ0uwNGSBrHQT3XoCrHh3HKLJX1/dY0DUgvdUoD
uqWBK9pQVsUlf9yRc0rN59LutCsiMIdLNfUMQln8WsH2KQ9Tk1zRYqG7nBJqsBbV
xZW4ywEspVShwaq+PbmQ2X6FTVIxRc59GRHg3D5XijaIx5soWWwjW0B7mdDVNbBf
dMqQ5wZ+UoPB5P1W5KD/QYEoacYAQhyGrUTUPwOahPdnbHxBHiNbhlnRVSV1Oq/t
r/pInFv2m4nXCosY87ZWiq52uA+jLWaY/2X9taEoRuACXE4bSzFIopFqjH3/8gcO
txCvR/Cp2WWHmSA/ztCtvaYoHJWQNurQ2sucLhxDz7cy35OCQvcT0WYaE53Ph7q3
TGoPIRjhMRo6lCajHJ1hio+mR0dRoXZY4vQSuJVbvZCVXj9xnHgUWMLm8X7DKU4v
nW8anev7+xw/izc3BPgXQOm5tzD2JsuAN/GJ453EFa7MkoaTx9bKM6SI7yNlv7+r
e6sS0PNj8KANilTGdEjyW1r8PuXMVCix0ALZQy533GE/5MBdqThC1uyf5IQw41Mi
THSJJF9pl9SFAg0oGQAwB4IqXhNX/0T7NwWrXCjgO3EZ5PkYYFN48EBQvo/pHxkZ
TBem7oHYBTN3kUYIRST/w+7o18PXVzdJIUa0tLM+AlrzQAE4v8/QwRKt0epjeHIx
qp9xrNIy0QFhEmSFEe2v8di2qOSzCA+c/I4d9U0Q08QXy6O2RAJL9jLbMPjDvzlE
jvtN706Lt+FiOuGt2y76Acce6ogND0Zfdb21UNxi/7YrDsmEyEpqToEOFZYL5mS9
sS00DSedJHvfLjozAisN5Rgs4y/ToDCeT8hevO99y9R+lpo0gzDRbIcqwN2/LrHo
OEpBO81hs3zLvh6Vx82u8qoA6dh6PKazwV+19+2/zCKg1MhfW1uhGrxVxMaZCDG7
FY8zvu+XW4gEO/6u9oaAvZMiM97eR4dyTpMPIbzAVduThJQJhcKBUJBVZl6R9BCk
psZ5vHj+x83bje2aHVZYaQqqL9fG5CYKM2c+e2lU3XUI7FgjqTk1yCNWGVDiTVAd
+8GThkiWn9HAfhpC+95/VIDgx/V0RS/BmCoVJHpDVBmtIGCWoeJF8BZHsBTpUtwI
LdKEc/233tPoEXcvnWjBHoZ8HLFtq5OuT1IjlVNKnE74OVxTBeOS1abMf14qBDj/
UHiLlssjBCbn6c0bXyIbbDKek2mGyQslHaI2gOmBb42s1nEOdk1gt0f6o/C7BI9Z
5rv0OfWgdiWKmEBySPGdD0GPsVi4TTiXPRr6CaYPlEG7c7andEaC3pg5W2P/8IIf
JMdYr+qvma20nG0x7WBEY3pdAZN9MDpSbLrdlR253zw2M3CMV+MoJnEjBucFs3rd
2JcV5YlZvIeR1Gdoh6lvPP/eJhhyGEhdptcT6lPf9vYfSd8FdrHuEsPq7dfM4KEL
GiMIC9iDHrOoOrYjxhcbQt/g2ySiAJ3YdwcRpJ7I8Mmz7RUUgjHbcsVFra0fsm/O
Y9qgAoAJGYIDJP2dUHKRRm25vitQjwUgdbI5VNomvdFqAWoUmJ0J17Y8+UE1Dv5O
Jm56q0ZGUFlszY/GTyj0NVYQFJtSGknwfNTQs2imyPkln6OW9V2ET0OrFRu9mw2w
Yf5gPReTsQX3nRu9hLliJ6f6+m5YaFDeZSl2txV76eaSHQnlH1RM0VTqPu5HL2/W
tVenBlRratCYPuyk8y+SVu17KunzE6mEwdLBqM2OTz4EZHyhrLcOhHC6rxPeEXRJ
S57jT949OdtHx8DQvlIAi+qKpzNGW92KdFO11Wokru6KR96++cltoTE71oRh72ux
vz21+FYl5uqN7kpO9R03RvuO64ExLR8RdZV0k+dIWlUiWJz98uywGB30MboUd6ql
twAceOMEE8DHrbE3oCS/XBdzzDUOQymAcZE4i3Q6uDzBPhCpjGjmQdc04R8pTybI
cJ4rFIn+kLedVp8DkYykSmygRaqJkHmTCumTarWfgh+W6egac5vmVhC2sxCIa93h
/TKofl8DShKROjJOCn/8SwcczBIcXVu4v9vJkYlTPonux5K0tOQ7PQ+t+5QFaZzg
bwCxeSATYpLzbpxGO4ExZHF5wRNkRxpmX3fuvZVsV5Y/MA7EM2PMVFh+0l7m3/Mi
GxFCLyvVedW4Qo7FBDtcy3ogPI23rr27Rca4NjVjpVOGpSImJFoBra7G44R+khn9
ppynG5VAXfXiix7/aSjsPa5m3nS0hCA/RtggWV5YSr+INegtyQdaznTOVoQVL5ja
cIOKDjv2/s/H4yYWI+xnDSWTFkABk5Xjt0bwEtEEO9F33nH5az1kCrwUqoQP2QJ0
M1DcpCCXgcYL0LMRr3OTZM0I/oZPQkVMa4O3oPnAOlBaRCuC5M/5iDtMLu7oYmAc
aO61dGNdMlG16SGNdTz+ObQ7dnTVRt3FEwwivg0ru41YUueG86mTJMnmcWeWntYe
oFjVtX2piWlALDfxzwYU6ifYpFPRZRM/R2V8airVk3gVaToJZVqHuM/N6mxsnV/j
IMIVd7gn3f2RQ9rtTrR7Kxdd8ZhN3NkJz+1v+I64/alJLnrYrVLIa6xtA6pAaFWO
3c6bqya5zydxcpbslXZcFyHJOCuUNhdnNFMCchp5eUymfPwOvwzMOoagzQHem75t
RBL9IWNMHXIVlJ4iQqOCDCtCEWuYwjjSQL+0DmcpCchMI9V/hNUg8ksqHqTvXQxp
9aXCNFkvgFE9fMxx7fzagoRTsvtRXZ4vDeMRmNxlVopjL8Z2pwu8lVd6g8fytTos
Z7DtHzh3Hj9bJeKDJGsgnUDgDuakUD3kwHWGyp3hxnO0D42sm+Vz6hB0gj6zAOc+
yd+a4q/Sxb61lGTp5RJtWmaEzXGcWH/crS+Q3/ACLhrqbn+HHphMi/Bo/ePrqQAs
R6hb1oDWM1ltTpyK6WK0S06i9aS6Sg/jvbY/Bniyfz3UqYcpPDnoVfS5JFD7szm/
/AwPaEIz4ABb9yRSs5ueUHMJLeVxU1LgOJhCg/GWBgHuWeo3QnN9nPZ1eSdiwBCN
SN60zWxUIts/YxZZ7o4dSehlL/CpBx2k+dhyZYnDR2TOyOXefCWsN7QAIvm6w25E
QyMuLDQyTZn9QrE1kTkx7eR7mwOUNlalPp4e9oGzbWZ2wlhgRvGJgm07nndF8p3q
HvjXGXUC5B/Y+3J62BgO/H5y3y5uPvYWxmTkSJw/NUv4OWV9SXGOluZihLL1BxAA
RO4jUQgWW/yQKTYqbx4RmM6vJ752zOdojulyGWdV/jG8iHPZhdLbMCfBMYoR83CM
CmJQJuaB35NVKaM9J65SZQ1/m2u1aPJMJzpniMWAmQaWgb4Es71Iewnl+eels+WN
V7F1/CYyAcBQvcJKXsQvyzDBHEkn+eIitY0jdIPMAU2uUVmZx855cINulmYC1nKE
kmK7Tr3jvg4rh7iH8SLMZVhiA5z95LcrV5JdIkDdhiYpxtHDHcWdYx7zMK7xtYRo
4f6Trud87O4G/ewPULWpOXhojleFqzZtmEF65OFgcNRkTch7l4F79hyYylLebgs1
8aVIJlBFN/m8S9hM1vJkQZRQXfqOYhc+FiuukVBIIaS6vN8ZC6Unlu2648bOZLu3
gyyQVZ93FcBcMpn1e2ocW8L0H437TZ9MDHukpY7gQeeLcQY96tdbpevjsxBF1jGk
/bAzVeXSYxqDqqVc+KSaJyDM2LYD/pIm4a0kPy1OPdjy3dGKZn01qGR3O85UZXnb
NiH+TrqPhq1N6l5m2Ge01WQAhkSoBhsAlA25ExQNSflIyzHqD+5wbwVpUVprenDp
LdvOGW9OBF9J61i+SYz3FdUR95+ZZz793Y8AUE3kaftXvkL44TO6S47Jyb2MPqGz
E3oWtxVy5Vry6cF/MoFFHS9cvaiMpLLAJ9w9dLjhF52VSxcGwNOOzigoFaHl84il
EwtNVQPu5WZkaF/5FVFM2o60a5xzWuU5btDW3YmvvF2nBpIdapnI/rv25RhOxULg
nmdgVG2OL/e4RaBLrizoe9xrRl+bXddz+6BZ/tEcD2uDJ1EUHJ0SvHWUZSFiJymE
jBQA+5AU6vMXTQVDPBHycuQ8LV0jVGWYf+NPaDk97J9u8lAWbZgPVaFxbtjVAClo
7sPrPgvh/4kXnTCAloSok9vZgZxoxM6W7JtCwf7v4NoYpYjdJr2u42UvdAFhK/ns
RaniQxJVapIwL4uq0jhsZJnZKeXhZ64u8KIBYpsiBxFJDo737UfHe3yudVvnLk00
kjxqRyNcCc6Nk1wDYFYVHDGez9Rxy4sZMPx1d3Mdg8pYy5xw4o9GDgKBK2qdIrFq
MA2e5GLb5OPBojGIagKzR87aHMbdEvtqB0SMrhzw7QQU4kR30wUI3ZfzmAoJUrXk
gM+JN1QS01pnv5Hy2sY8ppF9DPYWAS9M/sqMTOtiR8m+K+gNFfr3fmC/tM7M092N
VLlIpn4Vx2yNDJ4gdtCjtmIR+7z9PS1JNZ+9KAff8tmgnAaYSwGBgDeOdT7vJe2i
hbzasEXHAckN1sf2SRjCk9aqUurxdJXQ09yY0pSxZlr0RSe3AnQ6WoNfO1K0WuvL
yB4e7glpqm8a5nSqj046dLvMOWNBTXSnboJIHtsC1/ficsvfHbZzU28Gd/a7nvwf
1MocxWYl/IlTASX/ISvKiy/kuibHmyxpUka+WAMH04CiovHe0rOSvHnC6ncrHwgX
A50iODADTd3aLKc+ZF6yHDoBclab63QpDgGEc2q+1BL5vyfET5t1qi7+xL680OFC
aOdB2sIYP1VgF1yn3joXFihOhavf/e/sCOL2MtrZGb3DdIrX88jMd8+DZ9meI2Ok
khDt44BipZwadRi+ufaS9GUpy8CiOmRQfqIB/8x3pcy0ci7SmdvZuDDWriuR9gHk
rH06NKZ26SAUJkVZd++/TJbFQMFXt6j9WJka50USnQ8L7x8Cprr/1Jg+G25WAy0M
3I9CaWmW8thS0CGtNwHqhEXbpi3Z+B/N4xmNWkJMXFhp9ZhSr9GCJtXCHMDpCmiQ
Tvz04/IN7fja4PKHP/xBBHrxQDierFZq5fAd5hrFtI8uscpD+qL1c9lfmUJNBIQe
AQvzlRz+ft4Yj+rmgXZyJ6GFOkp4x4PVjX0uEJ1VWtPxKPShyloaKEbl8TIgmDKY
xdg/WMJkVXYOLqXCkI9CaxRaTa6QHJodqG5XsrGe8aqFcU+2YBH/5BA4vSN1F+BG
0qswkNgdehvrp8AqrNdVh/Rkf7HTIOQMmQTh+ldQHxhfTMl03mbCisRf72XofX4r
J9Xu3HKnMMUAw0UjMq5ueaDWeJz6XwIQSyEuOix4stYOVGl8U0jmUMKEGIaW6rxD
EbMkXB7atAv5uXf3MCLMtECUNwyHQ4cnbTjrGQ62E/Ud9kiJG+cL4s1bHE5xxhR7
DurmP51PGlBNfsKnSqljO1jXFOUZ8gXhYSSPQ1HH3Nh/bGtP1w0GkIz7+Uo/HkuV
98KK3eS4Jil/hlhY82k0307+1qe0kaHZfBnAMtaqXuGZ2Z5PjnXCtsc8VPxE38LP
4RzYTA2AMqXCHRc8Pfu8IMilUwBO1hJ/obm3HVK/rJmala8pxxVLCe81GfJE3lUb
sLmWpp8QM5+c4Kq+ZIHQU0v10TyAOnXF72a/oedHKPOEnXSgwbWUepS3/uLYDilo
QcaX6OU5uXoqrFtbI9Hl+c4OLdYBnm9ANohf/zTWmP1Hb6sIcGC5bvRI3yxMuMba
zMUudip6oXlxzkt0/10i3FnuiWOnOY6dvyaGB7y3N91FqxJmk0Kwm44xIqGhPGNz
WJ16NCwoafHc7ytvyH/EYybT4R3fd+td0yktyD49xM1XAbzBIIz6Ti2Oz2MfQJN7
KRQvqPycLMLnDG5Af01mSulfoJyNuwdNybpGN1+1Q2MiVyLBxP7SqTQ4IlI0NGQI
wg7DsQEdPSaK2C5AKc2oyc/E459wmSEEJ2tdobOo4lNcYxLdF2MsDKcKnjfpeG1a
dtKHHa4lOEdYe/17eMcACpcZiiRRx4jVKBUrCkkvJk5NzCAG1CHJDgJHITPnqGaO
Ert4JLwNYEfP+LdVBlNf2q+uZz3TVwyLFe488Z9M/SE+NZnYGgUHmMRfVto/FAUY
CKtCnsz4COEe61Ga4+2vhvkup8tvUjYFFAH5HfJY2s+3sHpI+/ACLP9v/VTdXtpr
00ELU3FnPVHrc1WfbSVE17qYTopVI/s7Lix+1osgtTkWcxQV/7UKdqaua4SkYbdA
ej0jMLA5K6Y6tZDwwYPsA34foPpbbi0crb3rojwkkeRr7B0ziT04I+k/x1jG2HEN
yIYXrurIwpQd/EnZ5nJBh2p3gIKLIbDtLrUiMZvZduHcAiJNwO/VwANS13UckRoW
CEwY6FQvUxAkm5jM6Zka8oWWvHDx75YCuHbZRz9h26O6uycg0OQZdG7K3YxBpE/e
gSbMwgb/C67o03J7nmEWgq04yYIp/x1hiEehzsnWALFOhUvV1VXXT2/44+wUPd8z
vC4Pm0yIzxOz/fs/5Bqw70ptvaNe/qv1RfaQSpDJ3QGAOfX/Qf3dweVdvXlB9RjB
t0KFYkx+ngBP3N6MscHLdnENR4JthOnLkwPdBqkmTz6bn79J1lQK/stNwyX6/6O1
39tEBlTkjIClt5BgNwLCq5CuWTsN4rikQQBbORk003PRztpajFNhNsoW65v2iVOu
aF/B8O5DzCjeaER9H/fh/RV2KdHcPKJSAfLP+e197o1Hm6hkvicJ7bX6VxtWR99w
+8OR33AokHjunX3cmhiOYxfjA4/3UlARaeSOjDH12Oj1eqPpyHOtygPax0weh6vP
435m8LUbRoN9yUWeBEMGDSusHjsLHEHkjrtAuQeMtt/sllqjeicQqVWTEEx3qbuv
M9OQhDHkaxRmxaAniBZt2X1oZPxnD7lwcJf8MCJFooBBhq8JqEgv6+xMBLDJDagl
1i8i+ccoGDEAqsxAJEcQOiZBsRkq+9OnPk1qH+r2dYxutDuNoS4IZ6DVfV1/UvNj
QULzpfJZBcOblWRts/5MffEu0NqtTUBvoiLyQ4nTd/YuSsnuPaSmGYb3uX7QcUZ8
OLG0gQaAhCum5y1m+PE1kZj1GBmiyyCk7wo1GdlpT8FIDHwt0/Ggy+oqGBViciM7
TRF1j8tCCUUBOVFRvdfL9ZQv4ahdeUg9yriMw6h5TMiMZ0HKr6WzzzH5mShBY2hQ
5gmZCocNsHUCm3XXOfw4tQFA0E+QLwx0/353833QtF9hDXKUsNDA2UH4IjLgZUUo
7218C6XYbdG5y1YwpjA/W7Pqv3mT61PAgGK0L1bkvY156dkt+iY6b5MPn8PJOVnH
M8CM+MbMdWIrc6daPGjb0B2BE8R3MYTbw11al14XEgyO6iUs85fnsyWzse9sQJVC
ZyOcL66G6R4vKbYFNtkcnhXMmPRIW37VgHZNWcIod2rL2Ql3+oi0iBh8ChO006DQ
lW2W0tX38QxP140xi1ug7KYldCtHmLfKogyFeyTkcR0xxYb0OAoyhhVfokApb/5n
xbVKV3iBU2K52Bx2qYlDtZ+K4JHWJ/salRCOUmPGUnVxYa0tWiwVLQylNsv7QuJ1
kEfiSRE3oydbOyP9CneWCYGfRkBVr3RqRerge30pCrAbTqbU/B1Ozglt5Oc2HC1T
n9lL8HBoCUqiciGM0JRN5RsGBXDajiy3xIqipa01VSTn3ofqs/2ilC+l0c1ihLEY
Uy+3EvCXh/DP52IY3TNzElVr/THF83CeW4GF9j0AgdLjwL/vjK/TgPu96n/tIL5k
Z5P6o4APnbns5B7l5x7hsgXXWiJRuc39EVY26J1ImdGkwRKAieQk/NsylkGUarAq
7nNDWNa5IlDuis99jj+GWnul71RNqUN/15nvI9ijVwe3PBv/6gDS22thGNLb4UB0
VdYY7YXnh8eTzgc4g75wH1eR0K5Stjx2W97iq6N9hJ96HROTymlMQH4MNs4gmI0C
n6H1Yxo2I8ArnJtagcZYjX78q10vNe4ET+QdwGLYNOxXWiR3ey7OsAowLkWq0t1g
wVYaOJxZ3O6NIlREL+3P8IZYFTJGyJvpUoPoBxsWEyhkAfmWHq5rx8ASvpyoL3R1
QyeaiD7ISSVIrGjw0+pfDq1yNAp29FxxUFn52wTcPi2Qckrlmunm8tMYsK+XIF1I
OvSRUambA3mQPkIUuQZWjvsY+Zq3dyvNw/U0oYQTcO5PZyd9MyPivooerybipR5T
fFKVeWTwDAyS5EpE614y0dW76OSTrFqXy3Gsfhm5k82TmVCnwGW6dDdq03WEl12f
M1tHVx81ucZdNOLGAFc/lAlO3WBEHi7tAg7cfCFnC7+pnGPYO04XrEvEXRQTiCBn
Aj+Fpgi5AFMATJYAD9PVkfxOFQPeJd4NCermznGRZRVCFUD/VWCG1tIJkM78Bq/l
ZuTxtfnc1tGq4pl0yD4IkAIP6AwvSQrrYAXx4Vd6w1cfLrx8OOMGwmTpnW1SOe2n
tlJMVsGgB0WJFZYMMeB9yOl2d4vUh67zv26ksqWSh/0mcdnrLinVwtt6SUbadiPB
YNTyX9DSrm92LfxkD6Oc3o2QaLPLfz7UxFe7Id4W+FHJzwkUrqRJP1545rLE8xPm
YF8PvkZPtRkr47+MPjnVEps+syTgERKn9AI0XiFKct/1tIXQRYQj2HLaHmKJbYh1
CY96z6xWxsifvS62Lw+FY52RJCalORfacVbM2ViouIkSrctZMOLvPXoahw+OkzMq
Ej8R1koiA3jw7pgjAOqESAFe5rCpvnjNyoug889KgSvuloJTUNI3C154acdozKGk
DkMuS6/7cxM7r9ebFdwobeVcHG+cg7zNm42OhsUWxBVj2WPFPy0/6NI+5S9J55dz
UY+u7wzlvn39cQb4eSrrdz5QVkhIbwiO5NU0ejpMfbX/sZ4Bz/2loR7oVHkad2En
NkHW3lb20aY9wuXWinzsEF3+VIG3GxxNWpme7htlNLVNgo5zAGfkTJXgoFOiYqHG
A2jeDJTHYoaseS5cVhaH0E6jDooIQmJc4EQGPWK6RWus/o3Pp6H95Ik8j6uTcKYe
akZ6bofwYyzXePSnVldyDqKiyJijRPc4YDIlAJSPFAlpK2COxq7p9kXJjPvlgB57
1LiTLoQlBxwR1B6n4E27kJ294lOjo1OONsKPARxNnsJxdERPYovze2PJVJJ7KSZT
jgOXGVNOlNALOnrQ5kyFWXtr9gelns8fIXvwNZGNW1qauZpzVGokKQPiOP9kEUir
rOgYszdUvaa+t8JqU7tk5GH3IZDC8mXofakbf4RyXUYj3OwAkwpVjR4Og/pGrM3f
/o8/N+Y12pye6fCvier6QBkMK+vWWv7QGPTee5KGUHNOfqoi2opAYAiwtXiQLKVB
mhbnnKtDDhfqx3ykXvRxkwuWdd9zBfBBXtR6iDjj0GcBcneI/mPhRiUcCOf0jx3s
vxwixIlgx05tT7WUXCPmaGvQMYiaZGCPNQFQhX5ZJhtxlk6j8xmt97hV5CIfNReY
kpMaWNZgfy1+aJl2+Yf2I/69sCXnBLiu1BrmVRuEJNSCdCmkc3gFSESBymTz4UoR
OgdNjV62caLdcfOp45eSAFFgJsQIIIkoO5F4ByBWafF090N2sSOTJGHkYwNZJvqe
fnVV9tHp5ehROD83CK1nzrxv4LWSo/RWJIIurThVWvTSzhgbw47a9qABQwnsibd5
SU77d5XZpDdxk4+zLKwbit4YV+r9COMqxKiqHrbogjwgy3UR3fcY7FORh0+hHAhS
S6ujf6u/LXWx8gMQPJB2d8igwsWt6rzQeKNNo/rWDOVUhSN2EKqZBRqW3DXPvWXs
p5XIeBuXVA/vpukqm/8nmN8XfKHNxd/2MdkdiKDK9IQs77dkGOHL6Fkugboa4f5B
Olf4hDEun18WdQ3AYh/Tx4FoSwqTsYfC/owadf/f6lWRA8BccYcVfAc2qOigVLgo
KlXhM3eMmlvte5gJGlJXTDjrhm/yP01WpTJWLF0eU/7kt9YeA8X6Q/fZFbAWdd/b
sJ8U+YWWt9wEBqJIDrTRcxQ2Xu+taWHtRlknuWmubV8C4a9es7oB0f1riXwpSDxM
+RieQ3XmhjJm0sIkh20s0mG4YrdWPNkl0Y0GaPXUTr3othseqDKubh3BP7m0Kz4E
JOk2K/AyAaD9nWKKUiqmk1WymI9uXimnd1mhQDBSkJpoY5OcwmBx+v33OCkYGYKI
lb7POu7MOZrTTRR41xcPPztH/oN7jOmH+YlqojIuOxoEDHKlauWzqcVFjomVJoLl
0N/+J19XrAXwPZpEEARRRr7j9/BFwz+6rzDrVbc8U1AdquxUiOTlD9G8+gO3jq8k
MGUhvWunM1qqjn2nrB/H85tkudoxanBZxqBYjuLkQXNoLF+iQoWgrnyteIQHjkGK
b+cywRGBh/lGhaFkiHg3mKCn2XYyOY6N3/y4XQnXuuRTMlvaPzawtwNfIHjlHP/A
9zQsPL4fmF/I1SAh44s1vmWxRhus5+eHVBl4ZCgiP7cLszg7lsqimyznq1u0t9iM
VtQpxASbiTGHfsBifsn5vceF4Wpn2oNYYZmgLTRhuBOsPzsiATg0RE4uO9yq0uX8
vB3DAC3ttTyOJp5czn2yACjs3F3pw2RtimunDiGhBJVxiIMPkq5gk5/mXdCwf4lA
eB6kmCLF3QBW1nYEqsrG3cA+U90p1wI8rQtXw5ME3u2vpdv0YXrZBG90L9Ka6n60
mrJBvvWmkAmXuhpbPUYnl4510M2v9RZYbFx0pkMS4xpfrzih6uoJCgHiGXz5y6iN
/GDrxrXzzsHHBNhkWLHPvt1Kh3fNTTcd+12PeSbOUoA8a04rm8o8YrXeBuv6RB1a
29DiqyyJm2rJEQjP9KVJMwvunkhefEQoz18MyizZyvmQlqOdjF0rgZmkO5O9EMzT
fn/HNaGvL13snifWQEoxIb+ePY782VSy6kiImBGdUPXyyqTd9hzPJkSyFXfYpi4p
c0OMAI4vZHeCLtZm1bBYlX3KYTOdZ4ftqsMfTMfr44epQ640/XbTjWCuWsraBaMt
iLMAAFtQwB1mg1pDNxqsPGNkpdrL4AXhL2WjSopviYBJKXa/UOlJZa98pxZHEVCy
YLIJiea+fuUKYnYl2gaepp/CYN5/oAsHeGdALVKcL7DBuX70LVSSp/lAZRh3ihyV
T5ZlLYZlKhGmgHFTF+DmpVdKeaEenQjlAawrL5E3FOxgU0xvpEv5gNuNYvGdkXxS
nXtbl7yntJTqFPqB+qOw2yZhxzJEEHMQLxMBG7I9WgUV6h/zYsoa/qYGRavmxSNC
2k3e6SrlW8Ox5sWWODSZr7pjBrWgqG9icp3gnJ45s9c2ncPFqyIa3FAnRLrQTJkL
MHQylCecd5Z7swAP7FeMNhwIDtWLEbjfOYxK8zYO/kT74nNKi8N4xNgW42oagM3S
/Gmg0L2QjQNjBOaNSowqUToXNdBUmf3SoU8mOS6gh1Otco5fEI2o+OXgyp598G9U
OA6VGfCWTcpFB2bjQ4srZCUFepjArcufH3TOB973Todc5plJXYcWqb91tL3RVYyr
9J36V3wwLtR/2rjLdgq/vpNlnWIx40r1jECwLZT+QBRMS55wfEG2+9qePKsiyRgQ
p9qTRfLPaQQUJPLrXIeGWHtHD+D5Vh+SH32viSYlkOKjx4P6oGmsMZlS+6ZCVF+T
Axnnt8VmpoXACNfA5KXVGt60eNutZfHg3mA43B692mxNig8ZwGTJXHmXcShVt3p9
yhD0E8OICp+mzHCXHvhMkavSI0vqFIx24H6HNGxgrow8vCi/mwVDxQn6a3ng56Ln
iRuUc0ks8b0V6YsYfwIRJR+anEXDoh6JzHLcznK5nd40cS+2Trk5qG7AMesygNNq
wYYdBPMqlJDYDwuqDSGcCCv2oznPpWllFxZJVKHX6ADGXRLA2tWYSfH6IDZen+Go
VUY56te4JrZf7R07vYFWtxrz2f8SkPacd/J1YQrt/MYIDxPhoGYfmLoYMdlG5WZs
5pzwBkhPecF8rqwXvHS57noQ/D0V+oQk16cVo7qex/hopgfrbxjMutUwaZ0KrkZY
lkLpnUlkU+fCmHkWA1Y/bN+jtw+KO6v8l3voFpD1x5kYUKx1lAbOOEaf/hGG8l7B
yN8M41rUo0+KQ6sWncEG7QdooxCytURRJVTVU9pk40piKxvumflYKUq2WQ+dvseT
dKHfRq4ty9EY+QQyLz66YI+YL+S5bknavbzr58lC8ndgPSElHiJyLJEmDpHxmz5h
iZb4e9PdIC9jtKMTNlKIg6DVoGNzMDcxdSBw3EOEdRg3Uc3s/b7GL5lQ9gmXdL8k
b97EEb+gQFTllMH0B6LKuy9ew0WuPh1iZCJKXtePsqfVWDcVwHbVvA2wo3frf0By
w3OIoTLqNl4eSU1i9fcCb+0xciiOICNmTaeNdIw3YCXO+gv1baCT7xkQUFDdUUeL
AGtwJDZBZOuHaUoCBNJs2GxGUIp0YG7cpEu+Sr0ZCwUMjK2V40OXLQEfHu+0/l6B
/gmsEwLImdnS0BvnoMMh4Vd4115g5cltXUqWO/yHPYyJb2WmMJ78w6dDrUhARI22
L+4RM0QgH2hdUbz4Uj7cWyxNmZK0XR7mA4xTXxG10Dl6oKvhW7Bn+im2btef0HWJ
zD7ipZ67l8+gt1GbMKA0QcAnGkbn09xOs1UnGj9mYnDVxpZ6TSVZ502whpvu6oi0
uY2FwnwpdjsxXFtLT/BCmiGSixK6Wjcqc56VaXIjG60qdSjsNE4aMg/WPloj7DrT
OtlGBue1JPLtrKhC4IsQ3DRPxVEW9UUG/1Ygl7ztmF5uChYCbdCcLH5f/wj0P0QX
Ih/EeCrEQPlumHUTZ8fN4d9hV1fVeic2E7WopYJ2fr53+vnwEU80Ul3s7rRe0G6w
TweMi22rwxEtoZJpvjrOkX7BX3b5wiPI0hmw/tVNRrWMx1aVmP/hV6rpioGRH1aU
fT3nMt1fsdTmpoTpI9UEEzC634hEEk1cHhHFnlxTULib87NxKHhv7ri10acJCCao
Xs0yJ69h/PssojrDoAmp53u80H01EaZsfiMBDqs2z/gq3UbYoXrztOplhUerDTGr
+ZQ1Z5Vs6fcSR5iItl/cx7LSb5zmURrWUzPatn8rAwsWRV25nvamuiE7+ZSgAVMX
d1aY6nAQ3DAFm7ze/vo5ZZp+SHJ1ShRF0IbVOQ3cyubLaryW83R1s8sE1q1HBj/T
RvQ9KIiBawelhFOkJ81gpoSpWMd8Yj6ccjKxuSQ6zzfyX4gKn51qxGkQ8nUr6MLo
x+Rfdtr1luht3iWTesptSEG7dOZy25HEc7/UBXnYrxp9Qoep879FxF0uDMEYFqSf
1xu6qlYcFZ7vTcLTVxAX7dbkHyQR09ycQxUd2iwKmoucC9kOKXV0oMbZ5hPjyyfc
4Ap+Voyqh6ckzEWN6hl4PeIkZhN1QygjiGxRGPkv/YP2HQ7t1pvQXOsLDW52djZj
eoHKp85cwo16SBN8q5uF8MiZ/5eM8golPTpz0GdAbi7NZTg6Ji4fOWz5hF1aTb+t
41COmIqHlxCEtA0i/1T0STEhv6jJ8KMZMn/rceagdGUlwPbhM5Viks0+gd1sARcN
MGEDyAYnldtKFSsHhYtHrR+h0i2L6RwpBFvQHTl9uX57jiQrioLfK86RYxaWWL0k
iVlRVuWg8Ylbw8i4f3ui6rrciQOikTSIZOl1Mk2/NZdL/dGPj8yaDn4i4c2Uktr6
ypuQp4WJ47GAPCc/s67lg54j5U2SUbPALSei0NKG6U2aIXXzUHZNC61RnehsiS3X
/tUGGArEWH+/GWawP7lEtjo8FCNuvvcAM+/MIbNE2zbDt7xUm+Zv02MS6p6X+NvB
J9DxoujiPh2P2F4QdrGloYbek4p5OrekxAurXk7NRh1Kq9cxEWDvp30TrvNZOZGO
88NaA5q/Ayl1fyMBtT9Lmg1EqL8DmblY3A2IXKzw1C7W6YUDlXmNo+0+EG+GULFK
2ajexUag/UCqHFi1+finlm4cUzH6nCN3kmYGU8Di8Qj/u5e1zBRYzX4+jHpM870F
/Ziw5TK4O6Gp26fOmVe6y0KmucksiLmRYEjEw7CHC/7KLNHwv6xznaNkBLqR9FM4
VnYDa9Vp2F3cSUTuxcptC4XVJi671J5mT9+qHPLFUDLLp2d0xNCn9GowgOGjORJe
55wKwdoN0XRYpA37v71DM5CAgvnBAqdpesU5eB81QA/F1gshiCWSEzDWdoCWthjl
9u4y+3qDsQetrfn9uVsrhMKYSlGPgCUYA7+uiybCxwUdtM/NMG3qk/8nO4Q3nrfx
zzJzrfC1jW8Uf54ggu79lyWcPirUYb/r0FG33u40SfEqSv44n+EG2N5OtRPLSsXy
890jowfY2rnv97NTkty3ODA0valYcnsmLb+AYtDTvhxrLqSCArAXTtTBIJf2McLa
OPjQr6XHS1ku+TZ2D6ah8xmI/xFlO7b3zbO4m7IacW+u7oMTHqw6gitti3EqHeEk
88lbqqbGnQOYVqFchnfbSK5ULnizFuM9x2thr4Z2M3DxPO+uCnmJCPy5r/XK2hJg
eRcRG7Rcq28C8KwgeGwQkNvzngZ2BhPegFSWNN6neypn6p477p8CmMa40/Wjzo+6
MwSByHhhAqf/Hgi/lkT+0kiHTk5MmJgjnIrk94nEELMGUiOWi3FqAtotVClLRbhC
hr/dEqHFEjsrBnt5nzyNn02PVdfDVCyRJ3k9lCYrKHBk10xGQMjNwGD9xt/nEgZh
YwokaDYJ9gjD1yx/6WgH9K+7AEa27Fko0Z1PFUsZtAc48JR8CHWB4GoQmrrfKSSB
Oru+jN3uJNE2kJFVCa9lObGJh+37jOY2da84w6LTF6vk42eIrTxUTHd0jUvz6uY/
Na4EBx9k38psq+wtsq4lDThkKv5cHQHytxND6IpqNDXmCOMPySnx7a16lASP3DNP
A7yi8NNAKZ191CSHepFbJoWr+02S+whU6uAOZquLXjxoKG+XxEwhlkfaULV76bLE
A5i75q+tlHRRgZhtjfS0yebPUJB9RQZYf4WRZbwEGPMKKcqTTIEx+vlXUh3/yHjW
T2eczdi3RgyINQ/1r6XZ3ksucFnKEWqM7AYAFOs4owFeE0YDy4bnJjkHJMqtcv0o
iypMxzojysJ3fPEYsCPqKoDQQselJBSz49YKVoSkYDYVBSuayItCXU81WVwfePXM
TRMqpNw701VsyNHmq8szBtoQ0sjJO+4kBoOHgkkCo6VPAk6tpEE931aPAJjlOHQP
iWdunXIBcuNbE8jlyD5vZi1eujL5Xkt3vixA9pSMg4m9oq7xEVPkQ8RtWvDECceo
Y+szXHJeOUN5JOqPqSj9sFeYFs6dBNtFOA1J6zhbAdQBUv5O88iArSa3wctwmWL9
kEVL+JjSFoHNvGxRnzksyXfjpmpdpxDeBF9oy61tmO1XSveNqc9p1sO98A6fLM75
Gfmtr5cxr3fMddSiVC5MdPekZ/jaVvagEzMWnd2dt+slTY0j6gWwHHs/xwhZ6XEy
/VzAm/JyisYD8XjycP3Y8ohpIyqgHiWV0KsJaXwDAcwtn5u9t2c1M3/ZjGp/9usV
lx5zY0dmasnh8ww2s9h91bh5ZJdQiyKmCxL7L7T4+PIu3jaOkYrYv/3DZPuQV1Xe
sXAREKsFo5pd78XtvT751rQhnCG9xO2uNHcUDnISfb9xwq6qp6A+a906PuBX3lCU
IVbqqKwTEBrtfwFZR9WYvqGXrRtBSDb542k6R9/tX38d5oqOMlC6A1e6ylAx6pvI
fwAcda+/hjER6rjDshcz18NQioSMjXL8MQz5m+ycOZmnucPAKZ03lSPHCJOEEcKU
9+/WDc3QBmAA7l8nnRx/EXFIK/dW/0Dq2lAxfIP6m7DhNmem8TbeIL6ARTAHoKao
XM39tU2ImXyTQCbupWQY+TrGwvLMZpsd8M9eBgRFEdsyIVGqg5CKE/lbrfOjfUdC
zk3x9dE5pnszkzbSGBS8xb69MAGPgTBnfgODbDWgCd/id4QRqsJZwyVhYsTS7QVX
DMsqvoh+S5LXmFy4kT4iOlvUIpQkUJdi7pO/I3LzX3/0yMPe1pCRgta+yGtj9lpX
2/RhkiuG6jt/7VTUdjkmHCy9fUgUAyhmmTRRSIDYzWiGao7dbp9UbqgW8GcTT9b2
hKXaTYkxsKDQUbUH7QNtH9Z2UUFobr+Q3jDVvgIHa7TZyxScLqEyMRq4AjPOELM6
37W3xjEcwnhlOeB3BEJcDvzy9jo8Zp/GJY+zsdhY1ReTHJOua5LJxgD5ubhza3W3
5YT3TXHX5kBYmHdlXcUGwEsYgJkTyBaqAN2ODJl6v65IJtE5mu0KIaieahXcPidP
oNLH2bFbXcu1G2mdrnbK81uysasIUTDQXwmUOKQ2RjA1933uRiuRY3/u3f7A94jQ
dXdCR2/eknmaxwog/TwqECs3lI3g+JFXnuPIjEf2ELKDIuwkfY1AQH7Q29DdNqbi
RM8dWPRITHhulrV80CigJ8qrndAa9PY8G+ixY+Cb0Y3Tv8xCkav43rwwrSiy55fR
Q/w/G+Qvx4A4dRlHeG3hQ47uZUNIqAxNixh8lDNoY1aXFSTfasnDBhqxC/8Q9L7E
mH7ceKaYPEF+S8rrTSsZrXS04ITg+MeGnT6RWwFsjghJUGOv/9hQqSsnTmKyKy0s
1drA6KxZDEtT93yvEsbQzNdndPZCWO4xK7gSUI494wUbao6UTi3gPQW5Z+A2+Ksf
Z72IbgyyY0wICaQcog7fZn20FuRTg0VG8OXHvmCLALRy7LjBldhPLK3Cg6VWza/K
PVinDpXnBwVgepbeVbSU5UFlWqdzY1N7QQmTfOpxDx+pvnLCN7oYrnoDIhLiQYVt
m24Ep/asDP2SG24SXOSOT3/64TnJ4NMTl358qOe+YC4MENdnkCAUUFmkolj9tFav
ALrD0tsnCwIRTHsgm/RbAChLVtl1wpF/9n+9deo4qJgRjvVnOoQO4fOgGkZq/mch
CHOg5/gLrv/N9WVI3K/SmipXKtX9q+Uo3fWUrD+9XKdHw4SaMwLKTwYGSh+rHJ+5
i4eT0SBZ6rHEQncFCG8fAo0jRQdf8N162GJLTKo09UsuGWHpwzpZFWd/csLGXa3h
WzHUYwi+r+36E3BjT09QpeGBOMOgT1t+hohJ9kOw5wQ2JCPr00cAaUiX1qNQXiTD
OHWaLodEAbWUE05dlSJfZ9qe/Z602yAlMhtG8+CPV2/DzsWIVEnghctmcRdB5Omx
YMiboaFiHQguLFYll4WbBupZCiMeY1R2Ak1HJWf+oalc+L4db20kj1X8B1556AEQ
8J2ad5uyhDfWYHMCz2GdggRqK8R+Ol/m+3e6TnTXrrVOFAiCevRyatfdV/RFa0DS
uDKJbLwKeFshrASV3PqSxg1RWwqGQCwvnTXXvK5nXHObuESDA3pz+grfVMJjqVGn
XxbinAR6tyilbLVgr8sLIcAEunPWqQ0ce9FSKx2YKBRVCpUwoXQo8daUTel/fma/
pl1aTUKnYJdmq74ZDHWkLBgpIUFyfCACkwjD8hELfDMQiJX+YmkTUmdHJMNIQZnd
i6/coupPl5eieultcgzBeHEd0snDINvsAWTHClRG6KU0rPCmxqdmUJJ0A2mDZUsU
MBSIBmA5/TTr7Zq3FS5txijSnTEUXDQVhz4KL4YLc59FPKgfHSsSPr89cX5n9bN1
iWsx/bXjfd+rGYtBBmqzS7r8Jot5USZD4Ji2B7I19rlDxYi19IGNhhxHvQkIxpOm
tdMP7YCDAzpZcP+m7HP5cg/tBiRk7Ri1+fOVOLBguu6bw+dsb8obnsfpDO+2c5Pj
f9afl9fb5zaq6rHsmDnVI7n7O1NQOwK7wDRo4O70ZV/6Zqil9LXiZ/+uhEuwgMA8
zoMMYjsuqe+WCzUdCwx1ESYi8AfxvNJoG1t1Btk68/uZSUdkhy+l5b/7UXjl1DyT
yGRJWG36XCH8AEjncTYKDwSJYlWF208YERKF0sV5vOY+HjsGaOA1QxZ66Cyz5wC1
GzOAkr/RSDwts3ZfCmuSYMToVSaxcpoP4PNJ/loHthipftaFqUc5ZiAMgAa8NszN
lrhm7gVkGY/06Gi70iID0mh/LsLUzEqyPaafmehwELCQnLGl65rrobJN1z3TkRZH
ydXHSEsesxqGMoiyz4BNS2Ti6k4NEfGxvyYA2HFwcwfePXebyPaVNlirC7K83rwx
X3nev/tQjSeJ7oEMimxLesN8stkjctvTRNtRFNM8CHv+HmjyEK1yTCRVgsvH8npd
2+SOGbJt2/MtHpKT7lBoT2nempkiw4BFuhoM6S/11/82ZisDCeSDMUqLLMQIb60E
GrUKWuvV8eTIgBfj7LCdinm33e8673g7plCv5ea3/MN4aMuzC0RNUUfshWfJfsfa
S1xPLNtljMRhi83ricEX79hhFaglZnt7n8h4PNUaGWCeGuOUgti3UTbNjbZzKr9A
lks3WW5+XrmGkhy0GfbRGk8s6y7IoUHaSUzbQwWsb6ILWU7eKa5pw/i0zq2FKocH
hUmfhb12c1xcN+P4rIdHbAw/bgYwrKAXapHXbNnK07YOegIrVL4JpkoCeFTTsv3f
Px4RIWHlKnx4N0itFm8m9z3zkRI+pOU1HLQ/x7OLCu6JqQEhZDa8y+b3HmOshrLF
UKJi/VvC/vaNd90T+dqmzwhDyG2WX55kt91igiZsUfss4sutYWcuWLOtwmV5YTYs
zX4qNkrs+kVRuMa4GDb6CTFeG7z6xYTt8pc/unDhYveUuES3nUfGrl8EbWZhDB8W
4xb3kiI8sfbKAgm9pghTjiKy8nIg+lyu2YAjd6+tgC6CuqNLOT0PoRSSIfrJ4ycV
vXGWIoGMasXvLmwklIDKsBBMP6vK0hMGgu4vxVpQ2FOfnCHCORVvtXj6WmMC0JQN
oG9Ox5J/CS/HpWerfcRYJanlCqNBvyXYYQE50YKLPFLzW4WSDhBR8r/twipQX9xB
ik1ItJC5SUpaM0SWgD+g6NXmi6tICKErUHWJCgkCsAQcNvMnrEketA20bLMRR2Ey
cG6L5iQFdWs1ZxORnbxwg9QGTFlLBEhcmT3vBrzc/gFECVdk7iJXDP48sIhL8ieL
tFHeEmHahaC0vI1aHnZT/UL4EUF4B1p2dcXkbKyxLVBvpgBYa4lqWR20iMGIj9KT
0gkal3L3aczv6k6NGWXWxlwsc9UzRFov4GWnmVQikfIymZi6DRBKDbMqcr2RQbmA
9mEXqUDLdKeSPtLhd+ZO6l8Ix2uX9SJiG87D1bxSWn76FU1+xKmd3BgBFkI1bEeC
LmjYJYeLoq6XBEDsQKHucrQ3csPmrt/JmeOK0oyu99tXqHMMFCv4xmSIyOtyMVCj
Lm0jAqbd69YYJ0nxIKGZItSctfcRc46n5Y/Y6Ay5fsWn7aRvyR8CXkjBEurvc+6K
1zmEorgPEZqDokXTZytdysBMnKLW3QAKw2lR6VM1s5AOvg+m92S99UmbMK3rd24Z
wZOreYBkIzpTIINlcxrVVj/fB6oD+9ryxpLDJ59kmvA0PNztPFSmKpAJbX4Qqhvw
yZBf/nybtiP06+rm8qULtgHBHeUQNLEFBEBaB582WQhbs9S6fdSyH9XCI3E+ll84
aWIigsa25j8xOH001CtqYl9UgDdJl7BrZT/coTY1cNowIjQmb1QPjZ0ZgE5esZSu
vczmJWwXkAPgfgsrZVHbERiHEslxvadMhRpz9VqqWsseiZIUJrBpCG3c/x3r017t
A3tzp6cmtdGLN0j9iFOTVYrRW9fw+K2MXz6BXroaXksc3Cf3v1Rjx4oNcjYAePCf
pwQgUpUUmwWdayDyXevz9blY9/yAgm8rdTnw8An79khjJWzaCkuhcRjvpBkXNzg9
dEcRUYMJWxCwGDUlJbOr7LeWtW0Y5g/ZVP+SoyItuQx8arZ+eFDBHaFxdjikottc
fFEcawa4pxOZNLsVuE/+bx5xDktPG0jCAermtO+lHPZC28JZWjQgtitdqqgF1/EX
V0fM9GmE/2vkrhCqif6S1NpPDRYP3it0QGEC2lbkxZD+72xxBhsaHZYOKQujP+Zp
a8IbmHJaThTuURBnqxOQkSfT9SoQT4TWJPx9EKYWRGG6D+jWmpcIB6MFNaxNj1hs
rVRnbtnTP53r2KGxZpQzdm0fZbKEBhYlFApejcfT/4BTCiEIRExdLJ9LOxzVC15n
u20URs1p23e1gX/z4Obk1LEYte0IiRYA/WVJzs6q80rpcHOCBwcWnFWLom8fW2sX
gEur/hxMH3uEjsZNCKvWZ+tJ1kt5E71YAzjKu69xtiTIb3duJFMtgWo1uRd7brl7
0hmVJHogtt/3m7BtCkvCq24UaW8llnNbxG074d0d/kF0xUyjvpkxQ/P3GPLTmaOy
XT185U01R7OZEJ90Dyv2Tm/KriI9GfDCUnISvkQd33X3q0qisCanrLEKPlijCSPu
J5A2cuNCyE6wx2J598DynVghSWeDU7GUl0b6old2WrygbUCGMNh0k/aPku+tm39W
44tKnXjre1Afa/MYbaAYf5Qy6tfLHrYTthXI2TQBvkIAkku1aPi8v64QhlTUmMap
t8UpfxVAuaNV6Vjd0gsbgsblNybkKiBJIqYx3nZpSHqw2dO23kD4/B8ltTHXr/k1
E2brdp77BGmALPE8iUGfodO2qJK6VZ7WzPy+UGcry+Z3KSSybndBpMKQeOofE/3s
nEH1bQmUwoOSL3exBcEQgF7YweJVjcXfb2Hv6HlVTMk65/bAfNHuRE19CF1fgoPT
mmUGs7e5jwSZPsWdl5/ZiH6YRsKbBtKJBgrJfMw+ZJw67Q4P5wIDP44YoXN9v50v
yvEICc44zE/LPsp7C/R1lee5YJDDSydNS6VOAQc7MTGBw7trmKZZOncPU/Pjg6gr
86V6Dbfp7RHBkeYf8vjInOaxfzKXVLyI3eUh7X0k4q2a8DXafvij/pI+kUHj9eiV
sHV6qDT1XBDH2dCr6QOX7kaZSBJ5m2ML9qPxPXrAgA8UJW3PpmBAi13L46HcF7WO
5Gf5T6bN9/UzzQjNWdzgIe8wSyEY6unRmHn1nB31nOcBqqvwCjTfUplzpOeskqCX
anZlkK2fVT2OjLye9xo1ukKPGt7gFWfS3ucKDdGKctvJTshtUB/1OS/zzGGhkt+K
+0kiePExQeNmAHb252X0a3thTF/ucIzEPzWNZrTKfITf/NZCQPDWaz2mP3oTlKAf
eUF5xpOMuT8lX0q4llqkfUoVavRMGdEqmpiKO/WZ/gQLcgh/32ctaeqCV5PHNB2Q
9dDhGRhaQsJ+ObFCwKhqraK+6vwJRU13yuhW3dXVO0bTF1qAPjTbbIeCfzhDEJIp
7C0z+Sm9xmSXBbz93iAhoG5eTj/IVnjePbm37w59TybpE0El/0mrJriPpFi2A2Ge
W1cV8thMHIE623whh9/gvlHIkBzTy+vxC9C5VYMLHrr7eZ5Ml4uqFVjnBtK5qvEv
H2FSTEo1jXGYR/v4nXnUVXUSzHHZeZxMDW+4Yl+2qSFs8rVdzUtS97HALSjieKzq
MpaFenmdPRSUf3gc9NjvoSTK37WQRHjYBnzbxt6B9P3rD2VosdfaL/bvWdc1J0m7
VwALk+4Soru9W6ne5XjVs+ptF++yCogObJmremYzf2WxLkPbaiECyxVVuuNL+Ig1
ku9FLMNdc53eoUBFWklCg7xXu8FHFsmDhg1oru9jw6KyByfXIAfOne5BRqH1FpcB
8OuMZ2YWSDSxbo8cK8pvERgM0rSFXZ0U1d4LdxTO1lF+UJUN8EIOMYYWP6mvabod
biJzqy/2/V7WWDnbhX1w1K47XpciOUBOelBDbaJcB8Y9UZBI1PO1NlFsYHFG5s2T
Y22uKIcEozK//TPWJw0pE/GcPZB8pJSzj/QZg6v5s6abCOT+jXnUNVazIMQoc7V3
7O0Y+p3Wa0bjgW84zGY5AA/H5sNoBF1HUaa/4DqLeDUquHO1FW4fejXo4GX+Gdqh
QRhBinqoi+LVtgxUPnfcefz+4igY3DnlF0/GVaO3/ZV9Jl6AUx4UVNif/pMcjURi
rxkR3ho4WWZvTmaWtOk1NZlbkMMe0FEM3KtXFAkKX6Bgmuw5jI1fKBBWkhzUCkRv
yGW01TNuMEQyCAZcCkKD6WClD8tB/MhAUQjXNHreg7SpmQmK79nKQllj989s09rj
uDPEYMdco2L6BUcRLp+clbvG/hO93MvDsjzUj4El7QLIPaqIdBdMKf4fLO2GogbH
KheLGHADX+JYety96/6gSZNNcOzINmjf7jM8S63p69l3NvolaLw+ZEwi5GS5JjiZ
dEI+yHotQxso7S95bKsfqdThHcbZL/3fokvG5BDjvCS79Xcb3Wz5/hAKUZwgMOdS
/DDceJKHyxpOc0X4WUmM//w0fdEnVxvkEviPQiDAcJ5KoxB91rWlkOlTefCaw6NG
ITCN2bwOhwyriuF3EVE3m2mZKuIeKxOcrWhYpAbjZ8HNC8ipxeaE3aaFoYN287A3
d/JOx8FB8+w8kmYHJ7YlycQQkagNotlfYNBPIkaUBIUT5yRSthc5OCzQ06F3G8JA
qvSp5uEQ06SCLy8zirDdWOVfEzjk0XHOJZaSYX94UUTZbEWIHOkY/hV5KD4Mk4Vj
9DR8Q4HxLVdDdCwvnIhh0UnBy922dhAEvcCdAHQCEmfuaA0DL9s+zJv3vkbylJAa
aJe5bvMrL6srbTlhcRXfaVCqv1caDnjfCphQyEgtvG0FHvb1Y0+gwDDr4tu2Yeom
qeJRjmPyXT7qU3YcOApQsIQ/FpuL32xG4b664BSM/M6Qraopy5IVN8pSeDhxPu7F
9AdKuSSrEJk4kaSFj6+pP0kzVzF7i5hWRkAvPaarNGECooHTTHN1mifo6Pv65Dm+
tjV2+rutSZHe2z1rirmiX7/9LBVCFBJRwHLqNT46k063e6qbnUpRgMEkLDc485dz
UMWBgCyIhgbp1BSeUrTP7gYoHqvGwiLyKQwdri2xov4dMP8EizxwogrI7pEigKka
PbeIpK0Ek4mhqp4KIbxwt27nD8No7Ykb9Nz1BxFgckfK/yS7Bx/+v/QlFV0nwCM4
c/mrRWldPAHtJJGHd8Aj7C/JptxwYkAu1m2fXYTyN44SMST0weLh4IPGr9QNyDvD
YaDa6BfqbRwvEHS9TybhEVBab2vY3QwtHboNlzScB/lXseejiKw58CLmR8eOxXrw
v94ZFhxSaCYq4DIwHGn17x4SUuYGBOmhTlu2DfLwJtAlB/ABB/ImyFC1c5+uAoGw
ATXzTl0rNOQUzgmnZWFgziAl1A259hPPcnjoLBqkxGnL0hS0kaWvcqW2TN5IUlbT
wAHhiQPv0Q5fZEaaqIwdT+//GxHecPN+3G8UzztcOBOumMVl2jDhqh0LpXVC/AYA
leyoyWb82pTFAYtv/SxZUJydlCFuq4Rcu6suXkRHTie/Jnnf/FXFxVIvtXosix1u
RJ7xibf1GrXBVpix3ggRs2TUVK2qAlfrOuv65vyk3PcD/9h3FmzjJFj6L5yX//Q9
P0VRFCCwhhkOZFXuDTkkR18OYrrCwSrf/pXPIcXf6iuBBYwXg+8AHjz1FZJ4kAJJ
PkFbSd1iqLk0D1Uyf9RGrbg11eahwixOXGQjBKke5cDpbWJJQlYkPt74NDXgaAYR
uIEj3y/n5Ah7wtqiyUcH0g8vgcmKQknSr1K0ypCerkBIgBe5jP6HSLfm65joQ5lb
MTd2uCtwrRPGk0ibuu4DD05ZIFMBO4rK3HQNju518rCJuHO+OnzMt1bFLF7+LDrl
1ZmIDvlqwD9XjUD3XkQmo6xgpzYVQLmjYTSrw5qMvbNzMZjv/A+Ug+gx8QZ0hmpZ
O9hPaOUzjEm1HVovtUkBxD4EflYkwZjObXuzecmxB4d3Jq8UQ0JkxM9T0lF+HthS
oMK1P5pEceZpUKei97rfc5z+QoBwGWkGf8RbgqAcajEgbGK95NWLI84nO9Pb97Wy
B4gCHBEOnKPbmNTMDIBGAXOgnihc3h8xHdroT5e15DK6q3to+um/iNGB0V1ChluL
482hS/hK1EFAh5yztAr/1oEwYkyvu61ucLnmpD0OXW9BoF44/UVaNjL3jD5kbFVG
aotVGaf1SkDNnF/5mGHt1531pB0xlZyMld19EAH0aHgUZ4Klu83vwwh4WeR7BytY
qER7XteloWIN3G9PBeCc/tD+lMSJPKjoaCgh9NRUN/ri/PFB7vsVfb7RqQTowZeg
DyO7SfTThYqka4LsaGua03vhNJ2AGG6ruGZZ928Oaez7pL64xCYF37wP3Kt1YaUR
qNGCicxpihV4ENi8vNcxmT/KVuSnCG4oEB1hxuzNDw6+W4GheHi7yXJwMJPuA6s3
Njj29dj1gunykF3xL4DTRCsxg2Tbzg1FGnrrIB97RPEHwuf3Sm2tGz0FXpRCDqIQ
+UQmkDU14xzAnF/AHjiLebwNDw+v7WXXyDcXVM4qVUBMY5HqkQJD3uV30lvK1PGv
qIqBCLidHnBexKo52+c8mpFKdyxTbgsTxMo/v01jwEP5eDiH0qkOLVpTVS4/GaZP
MjrBx8EG28+I/FGQ0Qoc2hHcLt9WOM6nmwT7nqoZLv9snHWy5mFbZ1dFot5mPwMZ
mc496bizgRJf+gXR6Zv0FxzEeCnJaEsqEynfpeUZvKDOTGJGT1+RfQ7ZJLAeSA2L
1j9mbxUQUBCZQrzSTwSTP50izkK6x77fiJx0xHr8ecqCvo6PIXp9VT388xxPSVaw
/gG/O6h9q5pPMOmuUC9AsiydoMhnwi7+9ZjL/AjqlQaHEYk2ydx1cenBNZwqR41S
wjLiSoCmUdhPJT9byJAZI9KixIWjkdiWtFTMT3aR77IzKm+t6iGZVOjh5jrsH/4S
369TdZsG4uZ/JJv+6qKkW4wR6UPlfpQWNWZVo+9ImawQ919YS1EwrdRLbWmz+E7v
sSidjcMUWq/iCk037vnfWHy+VfXr1il27Q2oM3EQIapa2LRaEEE9bqlQrEiK6LJy
EsrHyr6qAklN3eLwT2rCYnYwWfPC4K04hQ7syP7VSqJWGRO4LhRmOjZ2RS6udf2d
U92joIGY8c9a0Ux5k4jGlMaQ2WRHar6tbt4K+5NzPHNQCXr1jMrMFLuGg8Ym+K10
cyZlWYLTjaCiIkgkHrE/3nFB2KufqrITvMNNWuCJHzZW9xViQRkkV7MH6s+X/dyi
yUVuoqGVgNblS5GApKG6LIqWjz7sZyv6i6owHXwj3eGSW9VuTe8F6ajAnQeLkvYJ
DsU4Et6ERnxT+YnTGb2ycvcr1VUcL4JWnPAzaRU39lfUj0JxXD+wjcyw21Fds1eu
cy/Le/cYaienR43r0QFA1ZYY+DhdGJjkD8cwJGSZMJqSqgdS3srX36HNJWSD5Uwk
rp9Ru9Df63hP5LXrFDsxotCybOfvaeP+L5+yQSVEuzrYToAv0Rd1qNd0ccqmziDR
aiU0Dv8iOsgCbYLN4M30gXW+0qksDh9XpKvfVWW6R3lHZB/hjUG30/rRnOz5GcEN
dYrTeMtMxZRUh+PzIdkDsPr2QKWvzdU0L9GW0RB+JSh/Kij2zOitoQy2+ETJ/lLz
m0ls/9CyGBjenkL7tUU49iTOYL1PWnRiHWclpUY9G0/IfH3NnfHV33k9wbVeD8V6
ilQivQjCCyBM28t3vDrRUUTAkMNAXON2kgIdyeccRsE83fmKZRhcHHEoa04yMV0K
kW39jsbflyzOH7TG8icRoVcfIQ4P7XKpxemrZUJflgg/LXXKDazZ7IbA5D9E869S
c1LnxH9OtXd3l8LkoSP9aBq2m0ZD87Eg1fKSJeYzJN2j0UdoW7MwetnbbkmygOrG
o0MMERGRLUP0d8m4KOEQt/PcX/D8taDbFZzB2bqjfDIHlnJGJRoEknjjgowIsHdz
tmy1gzbkc2NiDdC12oA5kEanRr3BCcqOZblV3i+0gEec//Hbem7baUHLyufqD38+
V9Gdq2pjYA4jNr/bZ/TF1VHstoe2Q6PLicpEEuydmypBg+COVV4LG8pHFfzINqcU
dSYjR7zlAy3JMz4Jv/c2WpFN4pk/EpHJVoSNFh7C+cJVx0BSwved02Ijo52Streu
RQK+JRaGW9aCTXoQh8lC8zI2PDOriCRtH3lCsbVkHuN7C09LOXkzFFSZ//VXcUNn
5HXfeTmmk7ju2rxEJtNQI+Voj5gTnOucmqhFQVr75oBobT5oid14DVh7OatfEngs
Y4xr6wrQkAH67iEwUr5hTj/C20Db0Ms9PH3OA9Xxj+dsx1rQbEpyPunc0MbZ80lJ
THfZNfjDX5kF843UjaKyB8WMCSY3+xq3fnoU2LzKJVHVnGNKG5AUW1hLYcCq6Kny
1Gtxa3pJapCmRA8UGXgJP5CI707eYj/22DMxTpAk+c8/wHHhYUnTDi+xCswolmje
tNgZxAhy2yHuyW7Djw6Y7MR+ycHGu64K52OSSG1xZFpaG7ZJQb7UAjc2YFOic3OQ
BD6xqZpmtqajbYq7O7XvQ0p12m+grH5vX6bfiYfG5toHM4f1x6bmpaldv3nfJHZQ
rb6m1kNlUsUScZPI5DyqvIbJ9DUkaZNd0N7ZcKHpQpF3W5UrFeDPLdbXuhZm9yrX
SAjEBwKm3NVh0sAc+JHBHA6OMpOi7ARvmm5amFahdL8ePamdq264+QMnAQkZQlZC
oL9yGCiUS/TVsFUN06H9i8bmlDGd3sY2FZ8ppXorZt+Y0ZPFTVJ9u8Hz3PARDnx2
97MA4JFabou+vKOSPfIjNuKvNKzBM/ESxKmlLEO+i+O4mlN2fpd8IAPA4OXwqx3H
yUODscvNVTnAnEnvPvNv0msXWWo59XjCYAmhQ4tBKrJ+WZpeiTbLsBYDIZY7hzby
nGpbfptKoDxNo9mwHAHjEtkc1kNnHzHQaMQ5tA4BDp65+2nBuVUerN7x+L20IiEI
yZDduDd8Ts9efXztb8Rc9P1VBcExrFoymRzaFnjBclBMo9H241wSozCLxbEUns78
1U1wVX/PlPX2W096AzuQKV/nJb1/u7NasDpMZfcN/tPB1UL2CAZOueuvNwEEt3IO
WiDudnbdoXGuQ0RuRyUEGzr9Wgmb3LMsbhMNmgnHMATMiMfo5wOp3yCbfoYwaNoj
HkZIB9PhHOBFh7w/ulGR9GQIwmZpwMjwPic5kqebWiXb1jCEEfdIHrbxvxtxI62K
I8o6jL1nuz89SGs8L7eNA4U32DC4YWULzxKrA287Vs7gMxV/RTHdNP4kCsS9BE0a
ZRk2/+G1FJS8wjl8QjgyLEUu9hqai7ZEXctOta0n1mKx4BzsTLGuuLl/CZRl3dKk
Vq8W74umYsbW7FSltYm+Im3QUtXtUnlOCgic+YvAFYo97i02XMEafweZo25jAcvJ
WiYke9uJP+d48EOJCdFyapQ35wfEY3MsGVTz2BFO09D4CRmTtq5C314wNOiZFhR4
xcaoq1rspfLOsyE+ZnG7IwmFbNY0eRe47wJPotjhBLkAIP3Abl6ThHUiTRLh6WKX
ibocgMO8QXG6zJhKVATS139Fyy6UXfWGztGHhoqdT3Y5ICtxQxOklR//YPsQdWLB
WCThw5kbVX1wI2mYUXeSJ9ndyMkOBUT+EFTAhThM+J4FJN8BZqba+vtje6KheuFI
3q/0XXLNPgOx8+ZfUrGnCazQf/mDfIMbVfFRDOLQpKYnScODqWkf9sE17VLay4FM
6SYC9RAsXk+HYOuyD1fPX6UQfrKX7Rn7D8+icA6rtWsIGr43FurHNPFEg8Acu/Pk
GcdtQtu1+TtNEIoHMk5FTNDe6RSCWnZOqMUtDPVMMT/zqpmbsobuwro/tQa+3yg3
x72QMTruwJww4Uu5vrpwRwOa2uGsCwFh6YFbFSNTvXngRE8mNWgTHevROMOhl5g9
JKXMNBx4T/ERlHWluBFZzGQlrIYvL9GxNAJb2GFz3UZHjboULqrnzrRLn3GcAfgY
VHMuM1mbOMNgA9Zu+oiIrsv4x2wrPRyWjAurfic2jGTbHf/41IkgsZhLuXK8rjCq
z51AU+7jZAR3FO84I9S9ibrPUCEfnmuOnUdeg/EFjh128kPEzqS2bL7qEsYQx5hv
He3rGTxsBtMgKniDECOM/xRiuCMPqgViO7l+V/DGUMPiVjwSTE/oiCXcHUHT355v
W5NJSZqdVGZfdZj/UZxy80O4vBh8Pi4zYlFVZOuUhLN5Sry5e3TVkFvq+J5YWKAX
rvhORwdbSHs3vbzjWAe0HrxCaL4PIsSDVeDqlgNeE9p2FDnzrJ8iPmgAyWCTPQjJ
GkUaLiQd0S1fFBTlA60Eywn2sbU8jVqkS0NMRfOCu1587+/lZzAtx5HIfY8e/5Q5
AKLDrNNesFgLdiS0vsl9Rhid/zr1LWbn7fnbGhUJawYSLpKFND4ewf/LyK4gKDJO
5Qw6CNvjthe2Elh8BX5B/+80+9tZnMLFF/dSOijOWHAefyVRAotxRDa8FTr/Na3u
NxkTpIQnEdyKF2DkxMbaRvwreVZGvgkcVzdsbhu97g3O1uOLIXob7PEKxPoeMJJo
9LlNzIPPZNXYZr7piytD25xjog0O/jDim22jd36dXZCWBh+8vxsBNGwj3geevekM
v+7nwHmZi44Uq8mq9GkzZlYDWUNcCFmt5BUaMtLmj03s3VSLEAQMV3HLn2RShzJ3
Sr3yfNhGi0aB9a+1LPrnFyRzVIto0wXkEjeFqIatdokX5gKmqnwvjiK42H2OKgwt
muAVgiYLZOcPO3wmKmSTlKt6RjBvceqX5qdCA993Z+3n7+vOq4vo3b9NOjJaR3T/
DZVYwsnzsgNEC2fndVlLU3Wb2AsolIF14wf9jHEsM25pOsWDPUvLDT49d8/nT7PC
qr8oruoQt3gB9AHUm1xMsSY7QYDBLM8J/1CQox2fg8uQ0NJ6NlY2QpnnAMblbzUY
z3C35curv7aUloRle+heqoocAQYF5xBwkIN0KLWf3OOiULCmpvk7fOugAe0o1VOP
h6XA6IraJCkmAvMeKisBaTG/ymzv9OXBmSRzIMD+ULskiyB0ayQoWyD3njuUbaDG
+RjL2Z87Cg7gRL2K5SrSpkMbwUz5HR6ip2CYk2T2lwoOocKtqFssxP2T5a2ylAuq
CAQYvu2H5kNhvNz4l9Wz8EMfEZ5QIyAd/861SzxOOUSkH8cxV6uPDzwoK+GbjFs9
6O5B5afCJ9twJ0GM1v6X+SHx+JfPwhQ8DNoiJSQwYGGrxsp4RhBxaM1lZXt4vyeB
NsNfCp7D9BEFjhLbzJ+2DPDaD7qQJrzKHgjBS11+Gdn5GsF9oOV/xNCj1XXDEtm4
0XZbGjvgIBwIqZPsVxGivKi1svLMNRsso+XcVm709h/mT3OBsYUwwcEyOrAooMdz
8iRv9BZJocd3Ir+8vpnJb3QAPNw+0grONldoWgAUtZYAIXh4YktwnPi6AYrfDVus
RjzMaJQJicd2ngO5e5sgxug/LBs0x2T1bomhKwnADMqvdB9QAkySV5yTXHhcf4yf
LsXjzixpy2wmyaAuclGN/Krko5HeUUmusNJkDilgwTkZIHvOk8hrCU2zLzLspIFU
KC6vCqVzbGyh3cerKtkb3DB+caThVQE7JfxNURQdK5PabwBD5JnDBnq+905PfNrq
I7wkmLiJwlPOBclQOgWwltAAnswjgt7TC97z+npfPqWgHWbm13DwlDCvWy1QOstd
v0H8WPvxYcxDRQTbmfs9zHFmVqF2ndCd1AZTwpXxIORUm0+7RRCB0zgtelARSvCj
eORAlQEJdNzIVtHtELwuqWxcwdUomT4jvH8jMysgidHDXvgdNIMhwkuIioAujn/7
f49O0XyTU72vSMradJYr6CpQxDDltygVVZwU2koV3S3lFJ4aOMZprQw1M9MFHV12
DoKStJbmDsPf3VKzm0MsUiENvcvey16R3QAKufiGakoYjXTspPXudW1OrQ+3Ti2z
B8ofjSBG3pHhkx37tyNlGolEFXEvMDZ1NPxfSG0gvUvMAsKAN+eI6v37e9/sS3T7
Xb5UqNRwQPQLxtTsq4Ynuex+l7spCBRdh1WK8owiXnBf5k9S+yZzObLb+37WqjG4
I59mjq0bcMjIyioYdz0kvdSdwvvqHDsIGKtHwr63y3y2gd4WjNhNoayNIH0qtAcI
WJvtR24lfaA+R3nhapmLhf0UG5J48N+WOJnH5n61+bHdhurHj7l6UGEyvo4IAdUy
pb2Wuy4TJTe1kjyags1Y19CmFy+rHweGSn8LmL7QCzf77pCFCub8hF/lcTmAiza/
B0QcfiqVMj9bS1iNjwit+3I3yTi4nUMUAO3iL4fEQk+1zhA6NntAF+jtDZe1K83e
cgR2OzrOdn7qYAJOobdsOHP/iL4T5rwKcZPOiNH+6tuZiQWYPY1QdXgB2ImVo3nm
Du0U54aklkQJj9RP15pExMRLlGFrj8XTODJMrFXG6YO21NBCAghWXWIoJggUkpt8
/IIqc8KUCmyMqgF63UxLjPwhu6oafw/VFwUsNqz1jykCzVpiMG/cuRJy18lJTXXr
wzpko+KcLUh3aa/gABn0aO1Gq2gSUQJ3piOd+JBDrfwFa7UTRikMNAC5R136wia2
rb9zUtj0kFn1F4yPxxk6BIXn6jI7J85pVnp9ehgAyASr7Pq9tJKbxubv33bMi1IQ
X9aV4ehZYXsiquDUSIZGtA5drk7tR4CiO9CZHH70fXGYf+FWM3hml4Ta0A5EGLdD
OXWCpm9dSAl6DOQkrAD1y1plvsRzD4NY8DImIRqBALNGK14EwibgnSZaZwN6QC/N
xVh1A8zdVpsmIeUpiNhUad9TdnpMEo0IMChC7MSyPfOCgHaZQsThLZr5+k19yHgB
c5l3xNFwYU9wdp5eCuM9n7vo2wYjdE5qA7k7rPeSofSkygLD+i0hKN5LOFtfHDbk
Kb4FTrH6dxeX38KImeUHP/vlh4EmplN/DtCuX8SjKAlORgcM5AyRef/HwKBvGD4i
6T5wnWGX/rPwteGuBhjH9Vs4bU8sF0OLy8ZDQL+HqMQxWo1dtvDQSHZbmquRKRP0
HCMqTxV9VgHi95qoiKZjn1asNpfgOjBR8srlgDG/J/66e7eHq+u1gzVFfCcr8n8L
pzW03h2t0bnhp4bjrgHorf6pQk5+m50g3E5FGyHneXKjjxwAWT3EiIBfWCsGdQpP
JdV3fgK1jV3Qd2gq4CIC551DCPjL1mIjhbNIaWIT4v//KfTg9wIS/m+vvIrkh/a0
+lKjsOhvfz18TR3GFBdubNNRYwrkMb2FiMqlSB3xek48kwC7wYkNHtmGNSa4c3aq
klSHcsN/LaH4ee3JpfJF/SZtJJyCHuWqQbokh3sROA2L8KjiJYMQFGUTT6u4KLic
2BHm0L9I3mfpauljl6SRU+BDCR7tltey7rMDyjGV3LpPsFacrbTrlz6VPuvSS69R
wZg6hKh/0RJQRzTBWX8Nn4c8tStAwGlgo9VXc7Zmr6b+1yLhhzO5eZDGXUV2fbtC
+GIy/bMbt1viv0UFfh5cKY6xcJos4pXF6v/WIeATYv1OaRMqYaO9jBgTcKVJxbSX
ZDmAAoo9WkcXYTVuPuMh+hVCMWC2s5BGoybJRyel8A3ng5jb6N4Da8Wk/e9LCETN
dFWud+TYfbC7TvE+D1Dw+H8ctCzpzcgxzEItgX7R7TiZBhsLACu2Lmf/itVjnpYn
FD7Fq6NqhT/m4WnL2B262m8Rk4x5x+dzApt7TJN8oReEjgBu48tWw2G6i+xWNlu7
pnRpaPGHSFKz0LQjaCuchrvYMUReVDp7VXd+l4h0qbG4nUfWdKsk6FLA92PORrtz
LxUEnapAnEgmBKK1IGHU0v331zQ/XmuF4Gh7LgwaZoUz09jw9wyBE6YdJQLeVQ5a
J6qUAN2+BFUlNPgbD4WTDb1J//CBtTBB+axLCV6tiPq8T3+ogzit/5VB+LZfXO9j
VrULOTigOCtlhGozqCCebPddHWHWtSj129+usSJybdl1abRmMhLsJ160tdcp78EW
BNT6wjVx2i7rzcq7qHO+9ZuLLlUOmxYM7xvQaxQqQd9MJJFvB+KTlZbz3LMavlmV
22MZKOf4ISO+DLscyy0YLCZH2550OY717IX2Nr7XfBPE+4D7kFV3tcBsjO9V/MDQ
SHi91bHcfUHNTaiK6y/qlrNV5p+n31VX6fr+gQkTlfQXdp8Y/PBcHfjNQ8n2uiMY
HZII46IdWLCItAu1BnodBHj45WvRWWaray4+DRmrui9fq0GeQRDQBiC4bp//RhtC
wz6+bsoeTvKX52ALhaqFRXkbgxEmB2SmdkJKxusRBwAydmtc/Dkgs8bSHi72kb0G
jlM0d2QFzP5G12gFG/HwvU/y2rAvNg+PPpDtJAYG5z7l/X1Rngjg/62SwI/nJDaR
XKHC1KxdifJbg+1pQX0c33TXcrLrqbYINY1xfZ2tSFq1fTUcIa3JsYZWZwtPgAVo
bp+vF/ght5Oo/AJCguCaZRbePpniNiJIVzuz0C96trclFwjV2t/AVmFLNOW2HDgE
CKnM//MODz9iFZKTOqLF2rifaLsMB3wBGfL4f80eG72jC0M557K1TF6hYUdttUJY
2vfSJSeeKhW8RDj3oknoDHuU9UpRjnd5UqbQYu2Y30jtClFygVIyhoG8k6obyU0l
TgvAkFUBBoErbKxe6vlsWyzt+TmyN5hZ2zD3Has77nbS/MJV2/tO17sp5EvKHK3m
WUZy/7FWgb1CdsJOyelYPyesyPJk+DRNgOfFXTSXxteKWVQrRgLQraadJhhiGBDQ
3DeECE5ZHCesO0T3/Kv/2eXsmJHya10DM+nM2FFXWN9F3oq1qn2qkLUG8sxcyWoD
zF3y1k7MAhc3JNMxow8G6+5ZcmodCgj2OpuqRWeMaA/iPOxDCGhVQwGYuko4Ds5n
TEfqUIjsjCYocZDOeggeqWYA9tf/WUyRy1MSufvIW0rbo5ZjNfcSM8p00QkGqyaE
V3SGBKy4ujNVz9wekblGAigXnDIlP5f3rzMntilcbZsW1kHE9Y4oPlWS+evm4Ibj
cgjIedfEVj0Og+kMwuYHuBI8cPjqjQM0zK7Z2pj22hiuEwvsXaqPnG+HSRy6Zz8M
n1aO+9JMjlitzMtjGm944rq1PD6cKChggRSI8sVVRPNUKrlJACDCidV3FAkhtrJM
HUY35xMhMPZfgT+myZpARGs+al3MWD5TbfhHQWj9Ec+NTJooN9/maHwUofwQdQ55
uohhW83HMLOygJlFjs//pjLXEGukoMDjnZU7jPnJ5P2hWtajMbbiU8c3ooH9vYqc
yxVocaeUsXOAZDz3LlImruD2DIaEgmA/4TKhmYHVStLX9dzaNmiiE9UvE7bAAk98
3T2wmq4da0JQ7bWEVzMGkNCYu/2WxpKlCngQjo4HG4AJBO1tFBhq/V1ldV7LjgD1
kR1FuRICPtK5ZYySilLAoCWnlAOJaR0MGakhoNAQL4uH13FnZlvTqQULGx8Y84ip
WHJ4mHBN1UKSh/oL7wXt04cwUDRl2rDGrO4tDd1CXyBHfa09G3BavLxvW/q2dcy4
1N6ab/buZna+mLjK8ch17OFVSKZqJh/T0wD5MZfyouvb+ARhxVnbfAMGvnPkV0v2
0R3x9Pv927N6VUsvfKeI/pnC6mJgrO1yRZcj9oaGbHDMh0LMurIwbD8kaSsiUsjI
MaqPfS0H7BzaVtT+K7A0P0yzBBV+K3Sjjas7q+nBRN5tH0Nft21Z1zlDLYGyghLS
AWzgh+IWzrPz05ygsbohPpsVp4RTy1UcJ/dUqlr574rp7DrfgTz47B1NbfAXtten
dta3Qmf/8SdJXaR0Pt4A9C7zhWajR531kAG5uH3N/rePVR96W6cm0bwocipa0ox4
4jeflm+Y0g1/kMiAnWHE1xBLmLDphTqqOtXUxGd9AVL3JlEl0+cipsubjFie4okF
4IB3iW1rX/5P9l0brZ584w75v1T4vduCHe/x8QxPLAApRl12YyYR+kdP0O4AZFO/
j2dVn8LHx0ri5R953flhvPRU2uE7ifqWK2uE5F6zX0zF4zzONN+oa1dkqGT4tEu5
kYlODUWS/wdLRPJNl9z2bkICKjV+aIbNQZhrzSWMC5tnGZ339gwJPrk5eqAciKvJ
Yzjjzrv7Gh9QW12hF3nvMVFqZ+gykjAoqj2DSsbZD3Y52JTso2z4Ch4vHymak7V1
hkUjxRXmOYtCPhX8f4jtGkG4hWuT2HG1147RQJJk4/tuFg2ur46fHZ6OJ8XR7MJ6
vYQxVtQASpNaz8gMLjEJTFCM/N7NwyQdYf/goXUoOyxLwJBF0HlxsPia/VhzPwPD
lmVrV6M3tComlMdoojWI3brnZzz5CCd2yQ0dJMLWwL/PGQgGB1mOdXjGw2Lxmu6M
yVwQtsQkLgDoqK0zBSPVK1AMvO7OP2hCpccW9HAhX8Fl01hjVR4FY+a7ILt+7DmD
uOWuhwhHuypLB/zA40DoFOpzyTPv1tWKlxd9tYATQmcEOte6/IACjJQQumrOc108
bexiQjBvKrD8DSh096bawygKEZq90/MVnEuv8y7eNjYEpqRmLsEqHRIW1laGRq/o
LgMxEVk/MhulTZjpsvirvXcIaTE8st7GxpVtMory3zb2ZKIMAm3gn1e/XJ0WR2ag
3dVYYeMqpOaxVeb55G3cdDhKQLl2/5h/Btm598fR/rltAM/rFZAygc1Q9zSM8aYI
0kkmyWvYVKBAwI3ENYte7VuEb1QAVmm+nOqQlEEJzvH9GRMi+qPR8kASgLzDeIQ3
KlyEzbc7YQceNUztu42sEHIxu7uMef5wkEdyUxxtYXR60NezsIFWRYMV6MhUZ0wu
KYCnjeEcrI1tczVsZjS3AYPRAEVlLLo1DxvtdgtVHZuOeGCf0WREWiAE+ffDdpSy
ZGEyM0pcv14dLPK55AZ5CrVelidgPxSWnlFEKpWu2zEs4ZUuGYjWrfMp8oIWhsZ8
oVVyCQsCBwbuZuYdMRRqqEXDNNE3syrbRJFNskGqxMDVwjiR8kb0IyjNU++n1xvX
qkFuJuvlnOc/n4abLYsWeYvucTBJTCRu4Qp40kRfF8TiUPMwT0TPdlvWof0glqgS
G0Ttu/uC3iQ+zF6/PWYw6CS9SXFuz345PN2zadxFiZO3r+0JKCjivV3tsNpBIV8m
I8IPXWSwlALNzFluw9pYjdb5Iy4/KYPAVqub8BBROgd4lAwHTreX15Ssc0XW4IXX
PTru1D6GaTgehI27ig3LtkPVMEOL2rXrLkI4Gjq+tIzxrpWyWw26yq4q4ZPP1g+s
J04utveJJoZVUkdxvx6rvSOPZTXHxTNkCrcwTjnj6eI9oOIMykWzwgiWVHxBLq0i
aTvHexpMIDdVbEdGhzv6G1sW2vjfUdQMYeuB0lp3+AXilm3BXzqBr9iRyafDKsdX
o5Te5kD0+Y+yrgcD3Ez/vYMKXcrNFZevAbVASHQRP0HzgGMTClyYEwfaWZBVJS6O
0jarZaRL4GD+uiIrMcn5ZpXCQN8TXVZCohPyrHKU0Yo0omFFNhEdf6h+W2Gyv5tu
82q6DV+S0KfM/mC1woaoxWJs7KUSiE3ioTNdgMXJOAJ545G54qeewh743wom97W/
G+r8kaCKD87YoXDNul1RqfrFhhW1eJMXymVcPrntuY+IwMFtBF4+ph4JZr3IiLjR
bVKcPklC2bAGEcr4GUf1EFrLnFlBX/dm9gUE4kOlgtRI040fgJH96Y7ZqYeS9qHw
7nHtK3sF+yLdNj99a0GyRKQdLFObAg5aThlDE37wHi0a+3BC7NYmXggCEjZ4sEmd
+S0ML1H7wyTtD76DRIC/LFR/td2u7lt5C/D9cEctnQq3hvm2KenO21dMv/G7O4ME
SrK+2dxxYreiFFA7l8Y2Yeid3pr13Z07AUiNVf/vPpZ2Bbmd8PwFwkJ1Ycy5X4K0
W9Hfs8cEUwMnx+OT6BmINU8xCKtrZM6z/jJrc2wgUsNu3mOqUMKoc+GIcRnBfoj9
dMiJIkmsNq66+koHMADlX1PgJ8y9tb8+9cOa9wHv6z0p96kJWIcBX+vq6Fd2ugyD
2IuJENxRzZ5ZGAT3R/A1RIfPoHuGMS5uKagxeg6g3EbxU7MbmjG+W1uzyJ+OWTvp
IykOG5Zgvh2NooiqbXTDT4fKoMqfr6m76j6Dy+U7uk30KPwGN/dTz8UqXxzG1nRa
ub3GGNLxN7HBxzrdiMabiXy2IelRpOc0IP+zXxmIUMWFMG8jRN7t/sRhbdZVVBgL
MfoBxikebV9cflBALwd8idIpWjHN6HmWRPMCgpKAm0WB9VGLA+5fpnyumGAkUzCc
Vg+H1EQ41egPjczL5GeYbROsLmtILqnjhgpTAccvr/kiqxArKK0cN18OmTmDD4wW
fvfoorMkpZAlJE/rqyUPYj76qEf3VzBz/5bHqNnVWGrpKelaCf5/cIIUZDNCFFr2
nz8QI3azVNbcShqOtA/YyTCCAjhre3kz13f+iSAjugL64uRA5SmhBJ7DUKaF95Fw
8hIOlvRlMb0jgujsBGEuQFxQHIUZuv3uZo7259I5QVuREejmVbiHevy8gu2v8kfQ
VuyT16oEzHjD8Fio7SzbfBoeM0/hhbetWZJ6XA54wTyoMkbAt3NghMI2+b+YWeGm
It0Y4klwZga3sKV2Eeo1rfsBy0euKWSx7FJ5V7Nimyk5DnCj+jA3FNwCNOJi5N+s
Thbn056dmeV0bKIcpxB9S2OwbRDV0/vqoXNxgPszf42nj/F0ffnAs+Z3iEM+1zFP
tdSKijcVtdWcNQ6JcXddjjGtObi6q+PMJezfhrtqV3tSvlt/Q71iaRSxXlpZl9yG
S/Kt67ix4mLDQ15w4cZbxiqaOjK8aMj5ug3sq29qcyYNkxVEu9jtLsgVx0xFTtpE
bGdoIGwWi9zwRn5frVyXBgf8Ip/yXfWjIpcSLCrWyfNQCQTmbzwVdDTgW5bG2EkN
s+NaS9hwZ1DYI1XNASox6Jx9IcLnsWIzuFDxCv2ypwuAzffYdnvN1SzTf5//7p08
PsiGPrVvu0F5zmzQKmef7zFmZIKFhkQ8dV5CxKefL81whyrUavHwctAvXlGsfrwS
TZwt2Y+hCDDzZ4QWPbYX3YcajZZouKIis6nikGgujA3fjJm+58SsPMSHjRLqmTB3
Kz6+gkYwsGCtasw8yh4oWLnJpMeeXGrO0cms+hIJj5PMmgHm1GIvyxA1e0Fg14/Q
M5WRcHH6FXbbaC8yU7BTrdjIpz42c84u91GYETfOypzCwN8KVdDBJXfpErvaVpxV
aCJRMnFOt1jlb+0wlhHinn6QVQIKdMqiQMjIZ5EqlIeAaos668LTj1x2WMuripSD
nom0ScbLbVyOH97Ut9lNfjD5ufz3gF6mAX/Am3vbR0JRpZaFw3kaKMq8YM+6FnSv
jCpsMyJ3w02AuqT3NE6500/RthtSf8M7WKut8AauezWnX8Fkvn6OT3olf/1xVro7
27EyODI3KS2O8ppVdt6hAMPdhXinXONuzNRNtiTUZFK730Pfi8K51rTjQ71gtYhD
mtGPBojlboaJvvDWQX/tW1YQWPI6Zk8BJzoOggLl2Rf3E4JK//IEvgMeuppHszX6
nWLZO9SPU+71KFhiFuAO5XzKrZMscaDUgjKJGU++VLjXIn+WQTe1PdV9pO1MtObj
bAH1BIAgN2BmeWGaPdy7O1rC90eZ8Mj/5I+q8+bmhR2hOgsnTxCzsgfT7RHUvt/v
ai5nTysKhb5n7UYn7k9jOxo13zZldCSDnhxh4ymyu6epW3LmnBCPqI1qkW7Y9Jbs
gNUP6inMyTH5rkMT1gWMO58aXgZA3jwon79fZtRUClcWVANOJfvh27FpzNGPPkE5
5zIHfxPF7A2j8HutJYH+WWHXVrIldt0mG7WLNeCAT50fc+r8iHHMrjkvY/QqmaLH
G1SzyfI6fHCPjK6AdyjxAki/HSmH7FSplqo7Te7+AK0WK7sST36fhRwNpqr9G1nA
n3ZQtRCdvJpYWfZFU5xCFJunSfPWA/G6iY9ihDswOl8ec2JhF3hFZuCnwLaFx5/K
zFbPPgfMBbeSacnQyTRiZh8Mw1Q1UU7poP37pG1Xi3BPA6H1fXJv9syILtDsvW3m
NFE+52lkhHG/A6U/gbziocLmcFfkLribwJnxEVCTeTjRfw/jO3am8XW6cUAIoU4u
yt7+bnoGdIVbjztWY2fUmfwKMjsYXAWs/27ijNfMhLLIE/V2CDi4nTEj1FjsfwgD
AJu1bylyU3zUhvyJ1jHHLyNkImulIyCQ4nPka1FXwRNUo/WF+qBMKAgVpXOn6zXu
KFcQBuWR5rYbbZSRnFdtvWFrVhkBYcCeJmwUSZCNmaLkodElpL1NiwWjW3krMIn7
hxShpzBch0dPGok9mJwHBh1LVIUvT7bP6Ni3hlnmRhqCaOD5mPs43paZPPfsq3Q2
+i7XqR7W82e6hDydIyq6L45cgEVh030r6z4mhz2a2Q2rDV2mDOCxqwRJouo31AQb
JZpk9U6j/7eIPBtLroHbrKBMsRwce3pNhiUpA7rPWuthoRquyF5wsLqZsp5I2lHP
ip7vEPm3BE2reANqstLy+KoqhIw9lnWN1Q3ww87DeYf6QxdBVFdBWcmbLzfjqOtU
S5AUC8OU9SFR3YfPMoAExs9JNeJZ9LzEdFfy8aDHnjlbXXjWj2pO0f/bgF9hJow0
JoF1BYAsYFFuzh5IoBWbYyJzIlHRB5REJAJNx114jF7zH1qD/vfXRtIMnatHS+AU
dQ6gc8S0EUIXPyEDSPCltGjIyQjEd6zSq9TJkGXVC1Oe+gUF0oljhkGtmsyKZpxU
9MtATaiQUfN+gp97DRAsUSBpC6V2mehYZr6rE12C5gj42tw8SE1X/4uKXJMCmAON
26gLeyi1/ekxYd8VB5RweE0B3xj/V3pe8N4s+U9ciXZSabFsMML7UiN7zEQzfxmb
SI3ZtF5FVYnLgDOxFBtad//L/8ZPKzs3mcS2UiP6E1C21KQaL0f3Vf3LyxPihhUq
pwjXaT9PrWZ8SvhPUxuVxrq6bIT5mSq3P7DJPaoZ6zfbwUuwNlCNboEwXcioWuQG
ZTI+4lvWLxNQ8WDy6uuC9LhCAR9ptwlBoTp0fpqITXr6Jw/ZyysT+xOJjd32uDE1
C5g+slNQKUkfx+pxft19tXtFnu2/SxUmndm2xOZT6/hkrzBix1GhAnHvksJSmNOk
bteWojQt2RK8mSv77bg+p6YROle1yRy/LCINbB4yuKaLwDSo8ReZ6cJ02wU/q2jj
E8Y25SFVZ4cKglVAkMA5fPk4bczjW+av0nF5DvwM4Js12q40rV8Wresp6fJGLJet
WJVNdjyTcOfGtazhwoqOsL6w36w+lflP98rF978F3sT9x1gip+ZO5IMoKC75FivL
JUTWHHxZr8Z+DmrojJWPu228hrifZSLF6AmnSekEkP9yG9msH0tlSw1M9invzxij
JEby2utdn6HMIOs5wSRDEsIPKxDL+COBRoXblOm8q0F8683JBtJWcgt1SMPNzpd3
OrmZGv9egFs+hz+oam2aTdm/wyXTfyGMQ6EJ2MNOUkRNRGROA/jxL8HNd4CzPhl3
tOcZit9L3AgVhAlQal/RJvm6eiIILJL5Jln8X8+YLhnUQawIrKqmg39ws2dm3Gi9
DdaNoL3jNLEBB4K8fELRhNSfNT9jvL8hk2NDThxMdCQiIXad8oxEbOiQPxt7TmxH
I5EyOnt03VWV181wGOBg8OBXjiKlbzkJ5wUKKHFOBcqc5/0dS00W6lGWvvyAh3N7
BKaeA8ZNTz7p0xPBR5Zcyrfxh7/fGnCSvEiP0lbDrzIWKhPCCXswMS0Q+u7XpxtF
3JN/10ZuTI+MEfn7BifYzSRtWv8yZRkVodOA+9xY/qFi9OvuGXtFA0GRptQIZMpQ
qX7X6L+nUCKFCCeUPKyKSjsY/DOR4klmSQ+2c+0wbpWLYe9deAVHtOsb2JUFsIrv
wy5zi0yIZLx4PVLQ8xRADMdYNsAF0/Ffkf4pbogQMg5K/J8bY8dD1KL2hZdbwiZY
uBQmLgvJ3pkbcIzWSvqaUsPiwqQ/3C8BLL6S2n5Fgvrgp9PgxtYGRmh8zmSQBqem
oZDSp8aZfu4IpOHoDwiJUFmMt/AkQs0BjCLX0v+m6s0IuEs0YAOhiopntPgQh9jx
Syd9aTeJLE82Yx/hYthY5gRQn4em4deujkD5qjWBV97d9MEr0AXWAFlN1FRmyD8k
d35207hLjteFCs7g3BAN3YoS3tDa8NmfPRHPZBqxqrN7N/DwrErf5dPrj2+Pptvb
QRU2xDRb77pLC4sY+YtZMSwnsQoOR3dvrWJxaIzwPmuXlo2O3BWb/MedpGc5dnkS
WrXhGHVY07Sx/dkt5wNp+OmpQxe4lC6y+Gy6S59yst5o1JiE2Fxm6sZYo2K/o4Ub
+aNnjjQ+jsoQWwusQsOHtI5D1uEr1F14mb0xgqTgzXV5A7S1P6zl1aggZCD1eMrE
ouEV7SdI56eGuswCRIiEwFw124/xGhUCXhFmc0I4eylCTxRcc0729VlzT30NWkR2
a2NRY/0b8lBfQB0Nhievf/cVo9bLelZC1M9cLyrNXbr9DZXoEEm1HX7kmpgdKKC3
24N8zYojyahqxGCIluMZyv9Kn795bqaK0WUlyjSrj4GeOmsJ0jMl7m18IrwhRYnJ
bA4YBUk6AoC72pY5tzWJotfJpV3VFH1u6bTYIRrjSI0xpMpCE9zbh/I9wZjWedMR
8k67IOli0pAOSn5BDnPo0Wvez7zxHhwixC+yhHP8s9sN9zxrznWbVBNggZ02bzn0
7Q6FV5pH72bWimEm/sJBkzetQy/lR0AgHqSeSuZwuXby2hBWDhhnHxTadRJVT5gH
kDJFr4DBM9iOLJO8jdzlrEALwfe4E0f1+LEgW3iFRwHScsN9XmBk2IK6Hr2bAXiO
sOkxaAgT7/EbSXscfANVNYyxTzbtk1JSvOATQRZhJ9YlCIfQn2C0+ThEkFSUu/K7
T/SmTTf6QSA6AjXJAjxcLsz3FiTsaK0K3uP1SCzVkQ+RmSEVHlrhHRDRUfb+iveL
EpLlkOCKIq0gT6nb/X9BwnVZgHRo3tcmKdoRCYz1c1nnPzR2DRtFKRLCoqicqNJH
8pfKyeyLEiKz+tHRoKka/Rh/UfN+Dy2krAZkCZBgz3KZzhJX4S2ZQNiMxy2FoaDS
rixmQhdXpnSYCPxklH20RTQu/mT6A5DqGLF4LDkjINUuOKIF43pnOj9QXjxE5M/w
nE77PC6kJqvKoi+stj4+Jg5zsvuQ4g7ym8zExp9LJ1r6xwKtGZs7w5U4s45fVENV
NESMtMEPhiJysEo+gr3YYAD0lH0qaO6W2PZQgPO6Qri5pqK+m0mGz9Mm8IlT5svo
dWLRjci+Xy2DAB3fT+YmgxHtnixna6caP0ckI2u0af2TXT34+vfZZ3GApCQsRqfm
+Bt/SoSdoE6PqMYev5rFWYWn1h5fYumnQXoGubMiL2oj4tInIEhMcqHep9t86dwp
La5EVVARXDJvyrOwj4as40yIxZD+UA2qHGpuGI80jojOELw/PY4KF5spLbfWnQK6
nGh+vsfKqiQCwXcEft855cGCKZCENhYOliZ2usKEMX6rfKW4Q3JvZjWy910cG85K
UoFZPHBBiamzZCCwzXEsVWBiOULgiBIrviIJp80PNaE2ne8B3DX3BcwDukdCzqSj
y/e41DL+57fnQYrar3XpEGuhnBdAUmcj7w+rKl8Lv0rmeAY7KWJ42wrseZOG1MW+
nnjMlp8v+aSjVflViqlu7HeuYH/aCkF3ELINniqnD30EZPrEwRC9bZ/7rycEAodT
mj0dxd1f+nBbj5mjUGrUExNfKXbaPBeSduK/mmpvAn2+cJwHppqzjAKrAh3Z5NnJ
jL5hrI8PXAFI+DMG/rpfsD9+vKJB8AW48a6sPz+oIfZmlCVeKiUcAgQYgOY5QEAm
ee5aAWWDFT1t/g0Q7BqR3KHpR/jgzqwFeNvqbF9XHZs91yfwK5j5jHdXPfJKuqve
q14S8fcpLKh/QoQ5NQDV6GwXM/X7FdVg6OxTZDhC6Q7P2c9I3OS/TXGn1yiMKt59
ZNf94dayTEzX+JqecBNuRFMQy636wRNcvLIJ89yvyqebVCe7ND6f9TooOYfq/kM9
fk/GxuYydrvMvnbXTb1+39d5KSCB3RHCIpS869yj4jezVAIQqOgg9ryCljkj46qa
+bMSVPeUDNuISdulS1/juNxt6C7AOku0RGDWMPzdITU+57rMyKX1bV6tNp5s/xOA
ObeB4AShN1D+agHdzkIBDy9e3t6atUYmyJfawQB8jISXBk3okO+U5nEAGromOGje
2glwko2lYOfk137C/s6NorfRliJHkD+ZQEs2xhQ/krs56UftcEucniTBQ28NUaE4
G1oyLKN4i7Y4KlGimS6JrWxYkX6obeMeDCL9JY4vzYHOJD8+ID9J5Vn1/R/6PZ2w
3crB9Yoi0A82YtEg75r2vgmGn9dW6/VHEmbJltaTuJwjO1JBiv7msv4UHFfvRjBv
O5MYW7nV4GcAXtAIHbTuOJ5ZktJJPH/a06KjuSZTa6g0NkPYgG2CZuy3xtLf8+08
xzjoOSg1ycvUoa1bGE3775tS0YYAm/fmKi+qzMi70C0eMcIKVbKWxOESnt1Jlo7R
5IkaaaTCP1ChpQTzMCTHtCCbmU8CgcNzRtSnl83zHN52yzmQvz/t58jWKsu2zg2E
kxXryfoAmrMPY5Zy5w6esbvQgBeTSeyvWcAQWId7VAmY+2SlJs0MaPFbMuQsqgw6
P8AieWBcQs+64nkPwoRTvluiJGhSGXRhXqh5bi0DEQov4FNqXlb2sPS1gfoN2s/Q
8xZiolAE4v1rHNp0HXjqsyeQLnp2ACnXXyy87oxuomI6iokSHJdhMP9qo7u4ZEr1
7jRSZX4TmmcRoyubidV2gse2wIM+d9nZKBOROwlGE7s1QszWUhwuExfJqx/4hdLw
40hmFsYWUxqg6PrlrROYiU22gM82TX7kL/p32VRhvzotdt4yow8AUdVTYbMaKgLw
66hMFBtXl8y8RbxAp3wl/G9gTkBKzBosFtlCi9sFXr3gGLcq1YFdrvr2K2j4EM3B
IbTjKi1NS609wPaPfLgu+8jSfgPIMpGFtMgX64JCKwQepnTIeDGRqBjnP74gJCYi
XDWWIWczz2s44887Rn5Ql5KrOQxGDpenWlFTazFgprpT9+/MP69340FVdngJngRG
opeo2JKBkxM3QMT3xrRpmZSzW73JDDM3XHMbVPGv7Me1Tzoest6JQH9ZdlL1FapZ
/wzw2R4+5d1tJziVIyzOw1plVAkKl1b5TU3LYqeX2ZwYUvgo6++kf6QAgrwgpBZK
fBBpQ/5l027sdLWelJraVFhQqJEILxnCWYq1ReBYml49c68bWyYszQ383sVyrCjX
t/Us6SMIF7WLklRRD0vOFmJg0Xp8yuaamPgN5D6/fUPwZD7DPTUEoTf6mD5QHBBu
+pZVXIRS7JgmOEmd/lJPr/C3HEu01XkDBWKJWEBkCuZlYgPLGQrJP4aMgwvF7PN9
KG3FInbOre+eblMBfhcsiNO2phEsxCN8DrSxyGUDnnMOFensPOVwtb4a0GzmKtgv
qW6dZwx95EYS9a3+GM4lMU0+WuWRfRLKWuzYehwcAaWVuTxZBg7I23C5h1skqygZ
llfTySOhl/ofUJZM7sXKuBmp0h6/juvAYdAqjN7cfOrhCENNiX7KHhlIt0cb7XAg
XQ4/zjrr7/iitjSG09+dxeTZF4IoKvciGjyaMh8om6r0fhm5mvwrzduUELRjcoNz
F6DSF6bcBoTDZK5vaUMoX0WCNc3f+WKqhfMJU10mvPI9iec/QvABh7jBw51CdrcV
yjnabfk/wbfZoq4t4GvSkI51vnYdLqgHd1lkocH76wdCtlNAw5Cs5FKG8MkKqkrt
w/W2hK4YQUaBjfUFkWXs0y2gpm6w4O6hebueoAZyXOsJ4dBr6k7tnuqFYgeZ5jGQ
s9Q3Ao5fW5jcrfBmnT5WHm6vgFEapXBPYVLJbgttP5x2OBOS1xCvC4lhV2pCvzbW
qGn1t9xSoVQsyc8XISA2LNjfUPoD91cBpMfVybFhrPsPBTSaV+XOtbBq2bFytav7
NnFjRAUYASrwixhUT9MCNZB3lBt3CxyFIXnbcsNOzwqtyP0lLgMEeNElPCObN7+n
W+MyBV8EtoEMbbxJUCtlH5JiOLaebr4e9Sbo4scyLzmkX6WO4LM65PAhjgZLJbCj
95Zj8rxJJvz+dwk2tpWnDsUE/rgwA7ClaJ+4q7RF+v1fpFNmBE/PiZXgy7je1l68
VEPvFPYx4v911JHxU3Zn6Sjcawz7Jwe8HAvni8/IO6K1yOROCbM2ESI03UR/gdqy
RPXg8hKMYUdGAapQNZ+OX5wCQszPpxwkxOSM3KgBKiGvrEkXrG8v8r0m7v51ar/Q
dDPZLKm2zL8gx9Er7isFcC5G0eBHbaLe2chTDHg3xdvDVTdcFyhYeQofi086KMDh
cVJZIzENSHH7ItlRlzwqg4QIJvOm3UdxVC+egVnY87NKcoU90CNGXm+wcetUq755
vcDWBSYm3MDf4gHin3m9Y+4B+qI0DECNJ8I5VpLVSaHtP7hZsji0GJ3b4f496rfP
tcBn3Qn0Q+nKFUaz+4Vi5HHHGbbRnGAhTYN2GwWUN00+ebL/nc3jFQbU1RAPANpS
XI+2HTu7vQYDh+pW3K3D2Wi0zPnMCOvTDhARqCXDrvcaQSlSQjAYMwrYkADF6Oyd
KAhQJ1wLg/h5BLFOLwIooo96AEXwWOtsz1T1VlPatErLzop9wMG6LD8nUFHY02w4
aJYdh/435jmiY3XeJ9HeK3XrlvjfT/U8oAoxjR6DlDZ+3nHGioVd0/wV+quO8Iyg
jHTUvP9NAM1nb5XaE1nLN0oduEKwRbsPkLf8gnPcC4Tcz1gVVGJ2IMR349MaERCS
H31EHpUS/f7qDh4Px9ZAtYByI6xpDvCh9V3hpnN6ty+Ckwxij7qwydA7cCmFwz8O
RE0F/OuDZWoPxu8I2MfASrEYn0WollLxtqsgt8IIPFoYDDvkbzcoWM9OuGytGT+5
zhVsZRoTtqVBj/AuE4Owvt07o/WsgPkfyPzLyr6ZHShemS08FyCQ+2sgSi/9IIpm
a7tq5NtYqX5uZyBLmJKFdXef1wRxJDsyI8Pqj3jwtmfgZZzTRrO8i1jb9S18j8vO
t21HeHWZe2xI5T1EM/QQlPnk5rtKs4bfHfjOzbKWXUBtW/JhWc0VjbkW4GcTou8G
VXNVDoYmWC+o2kUi2U+rfyRCgFMY+WSAV5qID1AIv7XceTwA1c7Qoy871eOayETy
PJEMkafGxwmViJNS0vxPQ/sOp9dl5WWAQKEsu7VNcoeqDVvam+2BwKa3cZmOvPpk
fYUzjo29yFUtXJu1Xbca/FYbqJXKF14gzdXOI10aFd7ME/Bhi/j+mXGugvWrli2J
sxYysz+ghsY74fzSZ0kCkEzP9tTJKeYqu3z8jRyoJz8/Wb6FXpi5UXnQl6HUHWjU
rny+m1LgRR5A5UWDj1m/3zHrwp6neYw1Qn3ZJO3cTAvtOoBlfEyDB73r2HxFAol/
XOvAzf/z6U2Ta+J9k6Owr1cksm6MMbJdKlRJhrZ0UQ3hg5/BRbfbSp4SU7dk7WYr
p/zzaCgEaaw97wQaSH8xCPvgcwHqpo1l8FfcpdxzSiz8xVWN7JTGubIrI2Y8d87B
uuJNiy50iEmQkK7kmricP3SxWiKimQZNk+8SGgBtcgab79kW+In0B2zmxSiyzCBG
NQIxwSSi3p8NdREBk1uMZsjADjwTWPmpvvRcCtnFNoxmPLvMsprm2WVGhSysTJuR
FMCXnQm3M6Q3RZ6D8wK5cxLLo2VHA4Pj67DzWnQbEkN8DoOmY8gXsbDyRAdVX66X
iYOu5yG7zfD3g60VA8wDg29yJ10alfhpqxzaqfSn6YlRTHqnSKlEypiVz9+Kr++0
PMYHjEJk806p5V0UyLmoUuWtK6pZjRnsQH67pOIDITwkmG896oEjDgAPZeu9xz0i
i3k3aNMPxP5NykhWmOp05JlPi43qb2GzbOevP00TZQaDfw6YlEAbiucDlGB6CrGT
yO4T7CeObyt0hZ5v/qQYb/JIWJ3cBrrheBhM5dITXF/aQe2b+dVHqfmMOOP2Y8K4
xawh2rZ16WTcInMj0vQRUY+1pL2NFeHmsuqZL8JsT3IiR7Q8VA0Xjuk2lMIXg94r
PgoKD8D3KRVu9oCyjHSSp5DWEDNc3cy9LweWam5HKq6uskDcp1QHoef1nCNhEh6I
DSbjvqeppjs7tigvde3KTmLw5wA7bRUuajFULoViEapIceIWuM7SmmsCvsebm2Pk
er7e4/R/+kOmZS2tuZRLZNFR+7t5iBYsY1vpfOLm987Rx1RNqMAu/V3TzuFZD6K8
6xFFP8hm3KIWLx9xlIgDxMk6hbYsiEA0FHKJo1EmwMFwTsNKh+lmSs+riQIXKPkg
eUoLXfZkxZ5CaPQGbRqVTe6R7TdTHjjiPUbWF0hckHdycuen9jtI5nYS7axKciap
cfwcMFiWoh0X1/dvEfnsNcRjP09KZTCupBUiOtO2w5Gyj3AZnb0p0XQtzDq/mH8e
tOSrq8jNFfS9FxBX2B1oA1Wpz+GzDGHQVnT0km2zFIKNNtbtH7AzMt7Zx2x1nGef
gSKNYUm8DNE/BrCVokca9sXn7VbxOdGRDiKd+DW4r5qLRGihPzKl6LCEjPmwSJna
v9lc1Y/FHa7lH5mphV506Vd82KdVq+4Uz42xuex7mJARtd2sbjoKj0OIAuA+7fsI
hSR9mS0LJ0VsqwBIXvTNstQGgp331RxpVLAmUwMn6faFEYr0Q/5KIG6jM5kAtE3L
hj2U/eUYKy0ByGnWxvCULzz/+7PaZibbHazjl06DbgVS5sxr/qAucb6xAIrGUPgA
HBk44SWHDZcwlLpKZzzkuFnnl1ILm7XSk5Mlind1Ui+q/mvU5ssP/hDtmg4khV7h
F7Kpba3fDyp7BY+xGeLhGRvap/+iqx6WeYpPIN1WP2u8MG9phJlZKvjlgjUB/a6G
qEU2KITzAZwTDihAD3Nch+LXT/THrxGSeRv1tHsJ9sIjLQuM2O4Fz2m7aRwhdVte
jhGjk0jcW90QFdV8v1rqA52OQfjIhr6yt3QRPNwNVdEobkLrpOzeWlT9ctW4BkfG
KIT47IaWuznzWrVc58Tb6DkKAA1MkqRd+zZD3UtXPSy7XoxeBt303mbMoQLjfEWg
+dPwK5K4+8zD1t90pXgcq7A4gFe0WC6w0PzTv3cytZK+IAKwhwXW3mdew4gYfbaw
QozrnBNJw2iUI/ApJC35Vbfq1SPZjloheyDUGviXhHpEEciTY1lZtlVufNDloDSG
9DjwZH9NWOHPbgjoAo/CxxZnpnOGP13XkrRCNm2qVAr/f3J7mlXYEFc49LC/yE1b
cdXLIJVGP+CNWdMXoGl3wSLXm5oQkIBH51Jp6f8R+7PbcXufEqSmi9vAlnraOzGx
3Ch01HoY/Ml/9cMbZRIKBVO5pzKVgRagYWePz9v2Qw12XSTk+VzBu8KsjAn+M8ao
/s20bZMBN/O4zBzYHAnN0kx4J5WiQw4UQQ7TPLZigQzPkIsb8RVJ64dsr/i1+fOv
oFLPksiy9m/d5wZVYT+lpF5grf7W/Uillu7JRKz9AxoMixUNQyFCPKSOPMPtCgY6
KXntiLDseRxd/D+2wqf9ZUUkd8cpSm7KvXbPAgGMHxPLGHWqdsr08IEgA2Kob8J2
69u8az4W58u6bBL5gu5aky4UqjxCdnEAj1W3bWjxJ08HIVCXacusm587jlqkFwmb
Ny/fvj6Uvgqxr0DE0Y0x1jzOXMu7zdDjXUnBTEXW/2Q7yeoFJWfmHvTcI3jEdnw3
gKE3k9lVSBfAyvbvxVE3zmIFm5nncT4NstTiUvxlQCfClaN9iOtxqMorce1/EPRz
BXanVj1ZcdmpLYd6274ww6VAKkD7dtm1QUdd3uiWMlGF68I/KiNFC4nJ6SWEpPsO
4gqc2N/isu4pBUnuxyLHYwqO6DXt/TYRlm53I9HUTo3LK721gqIQB4FqxvPjNfZF
S5gRDkX4Ez/S4cHbqG9evOm9WhiFX/oopdpEcDBU6h8QfDpc9UIdceq6NrfYACa8
VU/UWcAJ4GAKVlsXzn3RmL8WtNbijpCL8bSi4Loe36Q3xGrzCYCmE/VMnIILz9eH
eQZwd/zuJVOuJ86coDamlJGHO7vZpV0T9JKGZkFpBp+rvT86TiwNTogpzvGlDFs4
QANc70NUfgGzxuADrbzlljJ9BUJbq8g+hsT5qjc9AhmnxbNqeQovKXiC6wmhQd4c
6oPEnVFRX0gHE1XzN0PvvUypLF0hI1N7ajgZ9jyElby7e0W38WA1f3fUxiXl4IUK
rtdAzh1r2eMi0wpCPaoi9/me7Ys+q3cZu4rALbMI+EYvgwJ4N9w543ZEUDVZIaQL
KoJ8KCYOXXZV5of9enfoW7RrVDz/bwlVYS+Htf5sadBA2jxSLOnJefrGjmjSu8oq
SYQRPLHx3SbCu1LpY+k9SXjrYxpz6/l6aQBkdpzHzPagrhObNd1ZqUdnEysJPheB
YJ3fGgKu5DQQsyHwuZijY/NEdNpdo9y4RkZdDZwSEGNsBji9ZA9GjrEvYL06YZM2
OYwmcbL218eoObRsl1i5uNkS+5/qWbmUNTMG0sf+AkYmV1O0oPDtL90t2ZC/+TaC
caqjQVJ7RTjVFTb1wCphA82Z0PZCP1jxXMjcDHwN59jsfvOJxrLad86z0BfHwf3o
oCwcJohOkvjsTr/Px+SXKNDTGwUbOGQDRvGz98eOirHFwTSCv6ysu4d27AgWW1h7
hbcNHgz7M42owzz8zrFWYlmb10emsahOdDs3j4WlHz0Bk3IBuIn+qPAsN4nfwutw
gc7AbtBu5nnXX+tF84U5PxgCZG/FemcVrgbpoL5mB/ZGdm5DX0oB0vWRPxFSX+GK
LGrGwwysnbnBZCySC14lZc8lhHsJi/XKFokRoKJCpdiAoD3dno7jaeAKiTWoJ130
00V0xQO4QT6874maqBfW2kPgrn/RYp5HUeIL/ueLpuEwyc3dLaRWYaKb3zEZGtxK
3FDSDVTZ2sByQxGr6o70VqvDbIk6nVwlafOXB4tME95aXhycmKVJ1N2Nz7VDk3kS
nTE8nXOavgGsEx3xV6MyC+j5S0v4ZA2E+cp5N6P89axVO4e+bQdAXQlIqoPOGgS+
MKmImdvFCjxU3GJhH3pTnjN4C5QB6X+BvZTvaAV3wX129TmaunFWaUfymq7R/k5a
lABYidkRadchx1RWVTeezDiZ7JujKYrTaCaY3k8keI7I+3jJ9uYfVbnWJV68MN5K
DN4ar7mLEdinJHfzOgAIICPqDgOlITVt8M8LF7tlcwSffkIGE4A8qay+mZLpxVj1
io94iV6hrjIKsuNGueWsiGforVF3fzdaBbQJZU4XFSjzEDNCwpCJXUXgoeavtl+J
veTuyL0ETeBePQqecyJW6sJhyrB9Zs8AP44hdSm4oCG7jgpAf+XBz8n+xwMEEhrl
t/j8PeiPkuWZGtlljZxgkilrNfqZlJ8RGkDG/jjU/XL0e9a4dRXuBaoxkX4jj84x
amM5CLAYoZLa0SApC1Pq2oYEv7fcN+50CntcixEQXA3C7DTkDTjVO3xzZjFqJAjm
BEMrFOKum9HDvvk0AZxpXnR409lTa7sVcPQTeSR42inL9geZCyZY3LTUWS0dJFg7
OEGqsyOCxt29m2LfSIZTrF2G0gpTvLCx7mkTpkROd65c/Ql7hBGkaDwDvi/HX0d8
M40GryI0WiXTN6uG8Kx8hOyv7jN4NRl5NJQ6zQzjoqIIKkkpQLkzs2IXY4VLI7eg
9SUm/DMtZDwdBm/FMPI5tQcgjXJJWVcmOyllY7kR2950umzXGW9ZuWJig3dqAXkj
Y4xkabqbhdv+FDJYH/baa4bS5mQWYkBKnJwEAN8+oKx7uZuqUeOFN23TftOrNHwJ
HDh72ivVIu2Gi/fQepHhgXc5pYU/5P3cDSENXESY7vstwug8VUKevGno9r36Vc0e
Pl2QaFN+204aqBgCVGc/gBuIc00T8bhe9t2vXt8naKF6UPzsQ/pSJMAN+gPQGjkC
YpxF2qRBfy2uD58CdneTAo2/TsN0/EW8pm8WpV7rvACFiOn5daOkRtak6DT7t4G/
TEGRY+r86vnRYYfwuoYUoIgxum/BnIfg47r/xHQUx2XoMdJo0ewIo1uKycJZ1jK7
q5mkrWjJZNgOGs6Q36BsZokvDkaQhZ7JIF06CMXl8eQitZdTFbWYjK/5yes1SgU8
vz7Stq3hXfeC5EX95mSrrjZwmrAWMmfPUhbwS4W2CiwJaCVjzkZ6/0k3IFlHhtHe
OSvcSEGNf3NwH1Dn04GzmrQJ6/Ysw7/N61SRCovhU6G/oaJDjKw1neDou1nVc89t
5pg0H4iOsuPX/lQ492OTYVGeBzSIWWcq2jLd7cr45oA+BNswAorraduNm8zMdNkg
X1Y4wExq3d0AirTPOP7N3ozSoZd3jPfRaIAzoGBdQqF5p2JVfuaF6ae0nBUVCzLU
8W5gZbBDLe88LrwYasMTWPmIdM4hec18gkXqXeDfO50V89nROSvQ1kTpw5ApT4pE
BVQJYu+kjNO6nV4TGX1FF4es4TPmgwLZie2Z8mvDyHwnNyy7/QCfjqq9WB1NTsKp
kdB3XUyM+2rtcP2OsavGm3ICMnMUP0KNFjwS/Mf7cHDYoMLAK6JpmDa2P5c+le/8
zn9E9N+oGO+qvvOcrK37yentMFi8MZg4n7pisqlE44+QDst4N9tcitDmIvpZYuw0
6jMYDvyD5QzDuerklA5JPCyAvVI8w4xxa5JuqceRKXeBFpJi2d3Wg77c3K/JnUDe
sMjd9+O3UM0luy7oRT1bT80jL2eGSckybUn/D2POWBZWuLdlrFQAa243vBM0anm+
oFHKvMFUT513Dvf7/uEyM6q4PEUSuJKf/hVnyyR1Tg8YwK+42GQOKBxvEzNfcuNV
DIyfX5AmCvgtGQj4DXyDjb7pUtwRlSCfIAn7HJ5gPjuHuF4l7TE4LDjqHOWui/Kz
tRCVrxUsFleTpGitJ329jgJlVAh+Fh076KkvhyZyrzt4hS1xMHq27drug+ayYq7V
7W/+NWgsbNuXNrWgrJ/dmmlQk5I9gu/3bXwxKvUN9+twBrFcjB2ohB44jJ3SihD1
p5pmplFaNfJvr6Rq8cEUhNZW52JZj6padH41pMRudDTJd1PSZFs8jnZc5FBMThIT
pXzWWBTXKVTzTTPEYLnWm9yjTxxjnPQyIspcqAlXT26uLW6kGxq1vq8lcuBmwcSV
6vCcagCnDLb1lzOr4IO7ySJ0n/MQh8Ta9isBxE8+AW5DdcVnzMA6sBaUhLcz6sM0
UpP2VMNHbC/QGbi22LvnGsL/b95ysHG+fCR7WPvPN2m5VV7v0MDqP3w7YTJoKegY
P+UgkTmSm3s+fonOQr9+kThocVpEbHRYvpQtkxheQxib0OW6oZdq5Y7Fb8+rb6R1
sYSnTtVBRFcUTkL8fkwIUxtapWAXWVyBRqbWYgNRFK2IJw2cWjitnQ1ZVkFrUWP3
W//GT7Ip17/ROGkILKuNyvBAP/YLVdyk1z56USJ4HvhT4OKdIuujuk9/YmBsaZiR
4HHdOtJRTsAWxhs3lNDNL+lHHvvkPWldQiahexPwJ4ac4d74uAYFHGAX/QUtCvV6
4erNkieKexAFO45YvU1jX+UlQ90ahqQ5AIimMGP/lGCOn5naC7I5Xaw1/Fr2Y7wP
WlI3IOUpeciLq6E9no2xvxU72afzAMhN1aH/4zewj9koyTCoBh5LgZ/+PSyUHvVZ
yLuRpgp/HqNZ+kVtJYlT1f3GMZzxE6LDDrpVCXDTu/TwDTkXvm/pkNKOOvYsQkJ+
E29VD0MgDdW+J0wLDFRb7s8JDyoZPHiVln5iCM64XqV1Jus/Y52hPsNRzN0+0mpw
Vut8LUIQB3hbgcv+1GqYOnGbnbwFT1LKkmJidWgLl86l6c14FgAEeDL5tm+waiSz
rcHU+Iyws+xU1LK93kpL31C8+JvBQGWOMLZ2MIlDejVG4Suo7mCf1erxxFVoW2G1
iqgVJfRl849eojsSfnR/IXj9YZeg093cGFgDuQM9AyYt/ayG8B6jpsIACNVdHzsp
CwKszH/MABkWCQNCM/Q5qHFWir/95LTbyZ1iEBBge7eBRVq0qQ6Q8Jzh8F3sM9+f
c5KyKylHJ36v9IdfQDmMCPhhdfuBfdu4fuEGck6sJB1y77toBNVChPl1g4G1Ljn0
rtk3fXJ4r283zmSVdaHaBHNeGH5SG/DHT62hzfy6DzQikjAZ5fi/NvJQV9j51cC6
CT8QU9yoHQkkGq+cKaoHKtv7DsZRQTil6IycQ44Bm+crQnOqM3S9HGptgUzdGrOJ
y/ti2oCl48776jYe/mRX8h/sfOE2z4RA/+mGPjScQPjdkzoYlMpcRevKyqb3f+tf
/R2hT5sMEal2JZJCcKL2cE8OdEnNMteyhSmkdWSuLwu39XOKWoE2phpQfQDQ1g+p
4S/bl4gb18EF1rynZVRrRdPkbyUjbQ7AWy1t41zfmM5aY1dTsM7HSDwVtZMO+gIA
TfP22CiXewPR0/4/PTcqfJW+txxdMPdl5IWPIj6q0/Ikp/qD1O4hWSSKM7VAY+j4
98na/vBjEmvLF2f+PRYPeXyq5ZbFp4IKGT7yLnr5GTuHIFFmzeoQPv6tXGEsEQHK
7415PDn7HTf5OX6Im6f94rZX7gKARm+Sl7dqblWP2sHiQlEv8qpnZUCyb62g8pGt
qChjHuQCIgbjtplEAYTMHqqbaSf82R0dOpW3dJestETYUrCoRpL9cmxOVRnkmRw+
7geKBKn/8ASROGXvIQ1VBQMeUMK+sUQ/lvakei0ZNemOa7E7iLg0U4pwmK/cUAqy
xTXsmK5Dib15q63a9EXzcgoEqTWeRyFZRjY/bWWXSB6pOr0mNI9t0UH4oV+7yO+T
g+MvM97bJWFGCnVB37TodpmS3NfRmuRTUftS3FeZCka5g5LMMB89z9ahaCfyoevl
LEnDDFaxANDAIy5VH3Yv5bsBShsm7JTvG1VZ5ulBtIIx0bBR4itMufeS4D2gvozD
a3VltqXUaQFkD7kHMFzYO+lw77rPOB970MnCIuCuAPEfoumyI8bAFncSoFtjGzZ7
d4QgLgCd4fT3XMtzYid1lm8wVrdz39rRJ6mKkVLPhwV22UcIXIi4Q3MGDkbYzANL
1ZtJIGKrlahtR4sdQD8ARG7PXV1oZqnr5UEYBJ+j0+kfZdVt20qlvmEsk/RVQoG2
z3QLfq8TcUV52ZBNwq0Q24tfgnI1Y635o9r7dYPDebIDwmnhf76r8QQ0N5F9RvYV
ri2Z3o1h1SNA2vU5elYMiwpN3gP1ZY705KQ/glJuXtjub7oZl3yT4iFsL2noM/RB
ayqRlGcIRCYSYVm7LMcynUu/wBHUrYJpfh3fAnVfI8vGb6h6uDYsHa9Z4W63riBZ
5MPEYbj5Uz8zpET5+nUdirSrJlXGxrWhxTixvPJ1xRd9GEVg4e/hh3j+zfuVIV1v
m5AWQD+qmd9Cp0iClWsDurRGrAvIhjOs7iNWxlzhbMUnf2PIeMIEWaIi80R2Ud85
FkZDFlFdOUOxie87b3mBEb1R0yUWr8+rhx16QbIfRmWs/LkBF6lpFTKqZETfT/bD
kxqdO99BBMhDQQSFB9dsUHOoMzjZMW9G1VxQtn31k8pPWyzJI9MZnDmFYsvQDLJ/
kTe8bMH+60QMGVOGYxpLnxKiZxNfEfHkFh47eREeqFyPPmiU+BOLfrNLjjs3fSwF
kvNQ8Y72QbKovXRqYR1UROL79IJn5m/vyN5zjDYeJEXSAcsnLPIRvFrWFAFb2cYS
fVeZGXIHb3jJ3hXtm5iAB+esVK/ez6vbaUrJWnqsoEtzsvZEOYHC2gsydrH0vLf9
J8F3la7b9XEY+tUyKmaKM2SrkHwi+OeDB6WfVRp9ZX8Mh1N0Injhi0Cdd1A0r891
udTGGYmfRXsZFo8no2hz2+uikR3D4HimbXb5a5V6xF+//XgA7TBERUr2hlm2DoTb
BTFlWdcbGw0+j+J2pySDMADSWtxMtuRZTg3MOTgdEJBJUVS3AmxW7O3SoR07MjMI
eIFCGhQfmG5vYw+DOnAxEUEpEC+hpfaPnDSdkRYbUGWGHb0KkY3cjG8fsk1nnbq1
IFXLZcu2Ln+pKYD+m0mL8YlYq1loDOxNimgle63MrlDwNUnUQ6PL9xVXL8VceZ2Q
9e5ts5obeTHzmycEEe6eB1x5SCxqaKPnBG2EDqqa23uL17C9AZb9jwACEUoGRRd6
WjSOydDU7qUFX5mMMXPbnI+ArFUWUkYkcJ6pijRfbp6eM7AQr99wPtuzym3LEspe
qIIWEYonKO/GAxkK0dXpYK0mTRIe8/beJSvLYxb3Jz56NUaDVrRLdtSbLABmLvJN
Qc/UeHjtfnkjm9xxvUHfw4ukT1iMXfWZBkAId1H1gUcxQ+k2SqMCJQf7USiUYEqv
kTInZF0JwimoJdoEXhUvjWXrot5WXfjxMgcilT/ws4XTB135n5RwsYIee4lLjo/7
6bK7xGbVd4x6+HjcE1kt99UhuOvJXVeP4x1T1LUZ8/utnHhWuLfdCzJOIM5MJ1JG
RuxefaWWOgoNEuFGuL0IWzr/qz+ws53uVRF47OLrZIYGKS8BP075BqUVwo76G2HX
MdJLMuMCAzSnQ2YxI92ZBz7WdF860RrtphjmtHGfxz8ggmIk6DIZK2G59UaNKzfb
qVSrgnG9caz4meolaTvlqovSQ/B0Hbifzz8ZH85i6yKjz5JCFKFq7oBZGO6to22y
77TWta5tBRTuWe1DHxq173I8IfnLIvAgMa/gPdLQUOp8Ktk3SRxXQLzYLHPQp3G0
lsc6I7Nhe2iYDPlGDmFNKgVs9cbY5x8FXbOkmRCow+mBerlBKoOZOp76JpZGED95
PCAK0ymhRHLmyuxtkuScQgGRcPm9zaWsL78JurQCY2JVSYH1YFWXDjfCnS0MZbtI
chRqTNvGHGptmZ5V4Fae47hDxntAsfZRT6ACdGIpKwEeT/BV2ey4B72+08Fz8XiJ
1YhIQryV87JXSJ9fiIOL07egQ4Iwwm6pYCifFyWc1Lc90ct3YUbJkO2wt3REsZta
rLYcQyd+Qb5QtdvUVwoUsEx/OQHuIjSejkC7y8qK9zjtU7cDP1g6g43NTyQfVsr1
RecDHDhalNfoJ36Ce0buBEMDaJZXH2JHKcmNVDSPZzLA3XGfPwYA21wb/cZOZknp
M8aj+hyj/vbTiH6fegVg0NQ4n7yLqLJ6BU/dkRawh8LPRF1M2QhzwB78vegErsTc
d/1AiPoZh5CG71cJTPq+ctHhL0bDMoexK0tegU3wwRPQdtVi+tk3LTM1wOyxN9U1
lLBvql5Rn/WN3LPKNB58aA8xNFaMHIqtUCpUT0nuz0D6osG7bGnmhYpINkNp23aY
pFhykvkHeTdV+ogQe9Q8SQmln16h8cnA2aA0GvUfBcXC22mMypfbK0pqoIPyNNwC
QB3eSjFh2UWSVGNAFg0YT48nAbu6viPx1zcuYLq/Jgl/BagbD0ylMlN3eXUMFQRk
D1BFXhR92Zj+DBzb7zejlyKMru0I61Cgxl0OY4YY2QmAWj5dNJarWnxoYvhtHzpP
NIHyueGNMT71ysboKs5vLGUX21r3yccOuO4lQ8SQV1yByAGt+kbNsjN24mDtf1Vk
pbQq8sE9qcE+ABVAFM47IeSiFCrJhn7Na4D7ddIMwuJBKWyHOc7+oNqIHwtKENvG
xx+KaR7VCdG1DqjRCzV3Cx/UbasWNLy4xc9gC3ThioVFBcMNoXv/RUuymoxkK57j
akzQ/o3TtGHoDLVh7bj/YvUCNju+CdDQXXLtSM0QXaQVrMNk8QLkpuPIZnLZLayP
2yPB72+3FvWhlf8OTjm8HjmC1zTOWBa0JceUGUWl3nk7x4R7j5Mwapu9fduzKjbn
Uz1D/uFo0YJblsw8kCA75Dus4YiH8Yg7iTbORisMmeui+CmbL4fjUlU1JuehfilF
dU3h99br/QJAfcWYoVNP5hG5iUXWY6PnbdhiSLNC5k+kJbVZVvxVdZgheoDkB8MB
ilX6zkswwxnGlrnrCRyFwc5lyGdrIHHTrslKGxYXTnWnc7rzgY0tpNFtMtljWXbV
5EAsT9U45TXb0XU3R1+OqlHpnjOOi+GeHZAgCvtq13RzW5E548T4/keRM7aZvv1C
UpjbGbzwdiqZ97VjBhZOuQAJhvm6zxZZOKVYGbEZEb1DjlR9g2hYQTz/pako5zUq
oMX9zOot56aD+Juhrv/OSkKaX2GPmpf1bU4j2jdfB2OnjsBQCwZ2eZJUNx0xXztV
YxHbZLPEzBZ8XuXxBRX1woMf4pvRO8DMtL6/d1mWWhHkcNtCztTNhjd4rPLIGBag
QaXLWhoF/llPM2yKB71Q8LwvHp4H0AIatOJ8vyPnxjkTvFXNT/IqLMP1aZWN+CZX
Q4glq4Rg//YBTbH1RojJbDZNgxJohLvEuvmeH3kS2Ry9Md5hZa+cNIywmwUJWZbs
5qhMpOnizsPn3XlO0lHEStuToewujCNAYn1vVo3RvcdydXn7/NElw+d2ihtgF1yy
HhZDHZPesicICPCYJjhKJUH7HA+W+Koq8NJSMdQ9PZfDPGFfJnOiwLGsMVcGwjAH
U1gd34Ojl9P4PlX4Af2wELxsBcwSGY9qvR5d663vUwYUXXrl7lYci56CYBLGlPx1
SdT3i4t30J1PFEL0k5h8+pw3V9oojUQqvT+noGoymgxqG15rIrvE45l6qJ8Bgxga
HNqZ2Sa08rpkGiNYKbiqbO2P0CudBe8lZvbAT0dyMMQnT3APE3kyM8nMzvXl7oit
J9isKIFbOUGguUcXmaS/BEWzC0BwJ0SGXR2ut6TkZdE0kURzu5r0OeC3gyiQKRGB
jCfOsrIqekbP2yDq72I+sL5kTR6RuWqlAZSur9g1VjeIWdQFokiIAbwYCv1NmKyg
CJLtRrtDhP916/WBdlKHYbAi/qsjphe2hZGn1QXJZtoposMf3oMybtNXvK8fy24J
zUZPpLgv2jnKgg9PosL/04aa/3uwps/LPpCTTCHvnZ6Yc0QWYpKpJjTg1MWte2yo
UjFUMVUj+H/9CpyOUkbmXUcAfaD51JdLsQxEJwdbyF5pmVUBEQ0NDnZsHkoLqzEz
3lY3mZFoQiHOyCxWXW6dGJ0vvJwWG/LXTox49sc3clM9VZL2b8poQ2xzm0wXuFVP
f1lPvYPFfasfawDXXDzrAAVOOSjaayQMd9XRLwYem4EsOsmAfjSLg53VUSf1TO7P
sLCQSpTobpJXH8+NJHNgpJxpP9xstbL8rcCfONCYJdsYX0xVC7AQE4O862H/WKEO
Hflz9keOniZmVqq3ZgN8KdYECx+KOrjPpr3XWUwkBfY4KknBq6Ipbib5Z5wo5tez
lKTITNr20+hMd6JDwmwwqRuwCcZ99Dkw8B9habUdPLAIB1QZrrBconppfpEH+S+V
hAKu9DdDAbk+YXiF0TkbLVHfpHTP06toIacYazFjPQM+yxaqkBusGrvg6PGF8cQ/
wzkZQqjy5bAfTyMqM+3m6LAOQc31MXI3O93j/YIawnttdWhZo1sY9LUXJ7C3yvNK
v2aIJOxFeAdZEtkXKLPPnXPGH2XZ/Jc13xfYS+o0Jy4RNlXi359+6H0SrXLQOHCW
algMnfqKkgHHrn9lLuJX4VLQ4gQpyo/e3xQEOhZxIyNSpYfd+5kgwuf/1A/46AVm
PwTqRTFuyo4fPTNR5FfncVMUNCPY4juZwkYL30putJqAIfNW+6/6T1AhQgvwvK3t
TwmsMS6tc5u+Vtfcc2jtsUOYco8L//jA65tlMSQv1zy+Lc8oC/k32oHqClqIv8fO
HJBKuTvEywwjOhmUSjIPfY9QVALYzefJara3vvG/StgZv2n9Bu4IOhwM1BeFRmqf
lS6FsiORTLZRc3Tlm/HsrBGaBsd75qQ294fuIUIlz4OenE9pfFwXnl8kGc5cM3dU
+Op57S7bgO9+0zs+BzGwPgGbN3+MruRvefQE74lpfYDskcW6tDUfas4aZBT+hOaX
7HnGfFPrnzd1PixqfDbzwt7s/Rqjq5yLGQruTlDk1Ab/SjA+/Hht/LLcgocb6b6/
hFMFfiKaTHRsEZ4SXgXvVkpcaD52jwt/1h6qo9jTIy91TDcA18xCJcHaASogfLWl
vgQsXJ7PQwCrsbYxG34SzyE2WYI2lnpuCMdPd4R9DdecanWnQ8V+DQAFs+RsxkCA
GKX4bZt6uUB5LxsLyr0I5v56vm4JYmeg0nqtCNGcpn1P0lBosXVo+Obvgi7zveXP
6gqWKfk2dSQQv/TuaLarrcbkF4FiPumpYcISiom+4vvxBKqPulSa6NSy4piSgbyR
XDjVY4FKOqJp7aj6DR06rldpHCBb0r3pdkpMEWVzUnP1x6WGiVQK4qcEdkQJa0Zc
h1nVhCmzsJR1rqcs32I7QGYMnbbT5r4QrPUL/MphyqO+6wCylOtmDeArn9dS5fgq
WY4TNoirjjhllQD11xZFVxWvG8EnGeQEY90D6w9jaocZWsns0abTcZM1dYkGbCKx
3hukSZPKUg2O+AvdDzzAo5wbQ/a3uar0xMs6Scu8o2JibLBJs6/CkO1QPtkriKPL
8vR3DHRmoOg05frDba5FoQiKsCw++1oYofC8Rg5phet2m7E4CW/k2eSNEmTqnC7i
l+0pXdkW74TnhSJqOZpwhhNs0x2sgOlFsuOAfDA75e4baXtoTlWlwDjy040gplsz
lS0M18fJj76bsyjanVbJWfR2Ui0J3glXmK8xZL75PM6Pd2SkkwFycDuaBUE5XF1v
xAXK+wO30EiI/Kdjq/bJPzZzOeqj7RgKTr+JCoTMnsOdm3SEnrEKUXq0LksKOMqV
rmQwhHZxlW0Tf2WsyA5buJof5SkwSIsLSLkCIQHMCT43lg+uO7FvzXzZtFSi1v3u
19zEkxsa1WTtqEouovQv1w2RNLbNmfgqwdBBKEt6eSiL/VpN2yaQg5Y154zc0STE
1FPKFV6Wpvy5Gn7SbAFlDpF2pd8XnBaWrPf31GSahM/n0paym6XHHUCWTRkky9b+
gHYUgo9FpUlaIbX4CDf7MxwJvSnYiili79x2pdPXhadWCUCqrs2/7XOa6ttrCLYW
Fn5jOhn/Rme+2QFLtIzv8DBNQgR2AhzIXPvb8g85eMRP/YnorNZc0lU4XZr/gJlM
sZLHvE3qxU8ASFg9C9C+nBs186fNj9ORuv7II4hZ5jR2oxWvg3pcVuJbO00N3F8u
oZFqwICBXaS5/rMMGcu1LdKWPSLStClNNXIHKK2xgmyNG81gVBk59QKDvZwGtyTm
11f9s8xef0rkYt2ZLQ12M7zHiSbHbqVDgDfHwVG1t+VCpqS+lCGWNhOZDc/qyKni
UJgh1Z0F2V7sMfavNcWBZCrEc20VYIDBTDMjERoE/tT2uvOdN6ReLjySKPo288rg
+rvPG61aM6I1283SZtlLw6CAYW4oJsjJQqY/CD0xUQ0w+VShU/dGxDQqPNoqDzVH
AqORgGxCwUsYGhog+hijExJi6F5wAoKGEzS5tajvj7llROvfsR+N2YdHd6xvATZi
B3ucX43yBhKBDl1oqdWkRpvKDds9JOmIlU5TvBk/1zoUBLgCGL+Cg6isjDSQMifQ
9NX2QIxW5Tl6qW04smJtbo3I0uqWzDQ4EZScbk8WeTS4ew687Wm18lHWR4xEiBGk
w4bERMrO6Dgfv1+5zLpD9X77R4EgjbywZXv0/VlTdzURAtCX6nJArxatr2TrbkHH
gpKm725ZZW8+2kHvCA1MDQEhwRKJK48YCWNwOON9VWCard5Hi1vVZrQ2k9ac3baU
7uw7qu0GbfOb90HmpHNc5Omg29spsVg+3VfhgEqg/z5ncGTRhR7/YIQuFazPJKws
qK0X+FH99+fp1ql9AH0829NhJ7YuVKEYNB81iE9R7dQWbNljPCDjc93qF+xlSYsM
/9ZfK5fW3rEK+N70MO3A6R8ntBBFsRCOxw62X9QcvgKIgpAtGRav9cCltIbUGvVf
POmB+t/RV74MOM7KybOgEezbX2q7GuzmuxqE8S3FHIFghqFZPPF+/VEoSPmNMW2R
jF8x+A6mqjGibQ3yCkbqMatexKLKBwH5lwrPrGSCT1TbJS/yiVIhX7JqORTNFrSE
C/pqtYswNXBLN0ZX6adw+EVUq3hB35uPWf/thcmaTgRC4l05yqfVSfNRTBClPRvS
30hpyHO9VZ1ZNPfLsHErpJk6LRjiuT3VJCIs+Ws1lgTT40bRE25jq9ODQGKkUPSm
QKnLlVo1QyGyp3qXhdtxXPlwX56EWCtA2ji6eKo051kGGMfI6vux3E19nBKvqUgg
L9XjKtSkszgAzdHfOAsA1gOmNCnWFOKatb09I+vRDtwAnS9E6W5zWh2jb72L6WI7
bLbd6IyE8rf9U3e18IWVHtSr9ZOHaNi1RsKNNWWT7A0tNHDHKhxHWeWGUbSiHWRK
+U2nT6+mGzW4mF/zCC6j5uN96UWEFE5BQWucug6Lg9UbEMVj6kcGly+5g0d7mwsX
uXydjjuXrVvdQ8kmBGKskF2wvPryYOac4SwPPC79+pUbatVRD8VScgwcGEj+6gGG
feO6zY4e7HvcZiED6KloGNZ+63L2Ay5+IJxvUmYPDylWfWVGgXJ+HM8kEh1dvY2g
tcRVnE1+xKYAnT+UYisezsL0KJxWgEm2fThhM8rJmaQ3cSfPdISfIvFZdo+UEs1/
wmLRpoB3pQGZ0r2p4o6kWl1twLcIk35db5CkIVUn8WpbxXiWsNRm0YOC1ceMqCIc
Mp3lyJxhLdv4MgJLHgW6RZqOBJ8HrydLpnwRubbP8/aIK2x6RN3YXi28I9wgDxzt
qdCfffuTCYdeLJ0VrKlUYGwx5xisUhyR0pXIiOMdo11lP8nAL3mLUH6qW9gIFiFa
b2tf5UG9RsjT9/ZzYvTnp3yvVpTG+H17kklDsyyKvLkRy89+Fr7RWeUT8mF5xt3G
O1oMDeeD4wZhhwAVSBP/l9TuK5bp6tNcsfrsff3bThC2pDgeQnef36Ix6s0fALnM
mhWc1ytEQ93GaDqhfhAeSiJM1/ALuWWyliNAxksT/TdBzNf4F9JzSbDQwRRMq+wc
mOP0vF9e4yC1uFDeHtZ6ulCAKpxY1iQ1YndJVlXKrklbvG/uz05pe4LowTAOmk3w
69jzT3fum7uadyXK/SBKX/ZQv9rIEeAkSd8PfHem3ocRSpOTf9ZXQGeLP1DOqx/k
Evf1WP30wjkiJtDol9o2XX4JnEOY/ggzoEabOBUkNS0ywwvJyaZHCJDYXdbT7s+/
uVy5nNLoz/zblbmaqp8l4yOsra/DCn3lAh9z4LHWg11KqpHMs57SCbw0X98Jla/b
YhYzHxE8Y2R90WglF4jr4Y/8HtVMph9FLfcUDYMrmZOExWeIZM3mmN7z+LrV0rqd
Ex4pyFm7t2abC9cFyxSzVALpclMH2quqMB1CzrBiEUJfMG/ydb8KmZIBfBT4YoFg
pleyOKbuh+bk1xTuKpZUHlUh5tnAeHUdJEHxf4uCucj8y2y4Np9OgfgjCu/xZRNu
8MErpUtqkuASHU1o/qobOBIjHQy3gUmeOSmkGatOjT9CeJwEXf9i30jliuZK1Qzw
+2FBHkxC+VJ17z6CR6XS3eAJ5kBLJV3d8gVXfodKPa6iD6hy3+XUPnd5M2U8ym/r
i5wIqT15SzAwBVoiv9jBn/+juBIY1kVXl2WBZnhkkE2lo/dIgDEbUSNv+glRMGUm
kK5/Ok4ZA+158gIHkC9JRU9kbJDtyZtvRhhAFS1GlqDUUPcgjpez95B+XvmAD5LF
Jv4kQyLp01l6h7G/Zs5nQ6qwhl6FOm0tc7P4w0Z6V1isb6t9vCElBC2GkiQ//LGk
3oSpwWnRoqZ1gFjhQ4HQse/nz3Wbl8Ml5H2VM2Y8RqcwbxkMWOZC6w55S73buzfb
BDC5rzYeY2M1XpwhqMumY6WkJ812sgR2dqrd1reBM0tW3wwwr7TK8QJqRa58Vc4k
Hsz3kmKfp2vtdFGKILfJ//I0H/8H+3yQp5PhnqdPPa3ZN1wBXNtC6YGcnvdq0YMi
K6D1e95haWll5xCAnqNnX32PcLT0iqhgDGfHLGt2lGa1+/jCbmY87+HyCqwA1Hde
mpCp4UP+VFEZQHn+IHIJUBqKi/slhts58p6ssZnfQ6KgoyOd8yomL5qSPjGLkxk9
CmLNERM1VeVoT+59ltf2CSQF+Yi19+5wykvZ63ACSffmPo356iaol4h48lcwIu79
hdvENouFYjozBmK23anmB6gzgS0lQUgYfS3bcsXxZbLhXUThJFXnlz7qlL1mkxLP
VCUihK9z4uLfKtqJ0xxeV4YrrCqcG3xMSyiLuZueF+AGZvHz25pUFbu56eOGiCMe
UIlyZ8yabKSJmdIJWtey1giDbMehWFnz8+n5Z4xtDt0UnAqksBFkLMAqcGxAkXjb
XIV34QLgF5xV9WY8ah3CfcnngP1z/4Hd0bya0CVhvg/HES7pQu38O8X6F7bbBJdX
I4mP7YbDmnBn165vvgkMHZt5DxcIeH2jfS8rXYkodPcGQtJwFD4nChicmovWMB4a
ad3GpkGo2GEoMARFPNS8ckcQ9jfVd5a0MG+0AqmHLWS2A/fdI/JycRsnbHRiXwQ8
vWLwthy2MeCjOdPHLUy7zNK9CDAglRkgR5D0vN4ri3SXEVrLEd8J2VA9ann6GWwI
gwfIdJECE17SaQ7xsoik4RQQXJXlJwli2rmD6miL7mZczadMGxFmTxz/2UdWGaJ6
Qm66NXdRwNeGd61Rh8pjSKNxEl1h81sT//LurNo0OebGRbd0BIbR9ZZxs7+UeqUT
iz24ZkshZTm6t1qTkRpfg2okmPPnM2S7a2SjLUF/t+eZV6WOOKjPmGlfy16BHjKN
42ae8Msx6JrWsFI6M+J0XxPEmjaMajAt2TyJd6hqFerQ57La0OUA32qL6WUTQIB4
r5v6MFI0ey0HWhBu8SC7WINYA62mKMQxES3aKYKlVAtJKHcwRURBANnxCmD/8J2q
CmmsDD7aT96vyY8ZH6Qs+xZeE3+ZVPTchkLIhnSFGYLaKQGaf/twZ9y4XpjcA5A+
tacSN22x05SYUe+kvFRNiycP0svH/WQdj9YnSvSBRgyfkbeYMwtJ3A44Ghdq2tYZ
FLEw0zkUdWfmmdG/nT1EgLG0VbpuPZgIXcq9bdqsUrPiawhoGH7cttzBWb6V17o6
qCFeur3dzBoLBQHFgOAnMAjxeWuN1C1zeFJYUtquxS4oqRgMPY0ituLZ+hljrUrG
jisIBrkP1LvAB/3YDCMxtjjyPJpW5qQSOiRTUYpqqmameiRcsNpOX2+EhWDhbHLd
f7dKc7AsSDh9nkyB6vt7HLnIvGyHsfryZHXQtWM9DgHqHmBFabTMSUhSc++gHfY2
w87KnchIE6R/fCdZT91AAJu/iDwQ5+oZiY28n+G07iHVCWPn4vPTmKjKSTfT/tlF
sWaE+fBV6SdCcLf5+KpgcJd98+zPDyNDXNtGbbpunbNkmUQpi7rgNEGkLcU+gqtU
N0fNwWQnN2UloBwavD+EzzMZFt2mSabCrsk8sYWO7/0IiNf4oxyuSBOwvsZvxq8Y
CHbZUp1C2+uBni94YEFG+YiLgd6APlu6wPokO6sdISWSufI3pk4RrKgnyYpnmrH1
rJX5tcb2VYEqtBKewXPq0xjv1vuB4FYGbqpvn97x8yP9bj7VoEA4bU3rInGaPkSa
Ula0fb5lsSBPxFDzEmJW1T+igzwOzMwEUht4lqFoP1F9WpiL+52OX23i7Iumda6c
SDLFicpWSnSDdqdaGOZmKn2z/6opixn2xqxqEY7SPILsOzxQtJnPVu6rEfyTI0jn
vwPzQEqx1bsffeDGfiItWD60kKyBvfLJY2vspcBn7PI0hyN4Lu00agWRDB/R6Sik
t7Dbg5ZkJAGJJqHGycrQF+ohbNjpGJ3Q6j+st+q2RIW7IYllvhAMkJ1d/70OGkM0
ITOZE8hOhG3Gk+i382so30C62pfjS5GTXe2OUMQ/H+JI5SVK1dVwzgVtaguH37Rg
QMoQMPJRfaVgBOclIFxzNg8cyGSvkLKTOrKCytNBup5SZmjWSQl/ij9IQBSm59ac
ysxFjKQgodsFgWFLxpb/UzzMCvRQF9nkVlDTyeUlWTfZS6nYeQw0PJnybnXAmpAk
nY/2/oPBZpdAXG0FHu45R9yh8WYNyAXp2YQny2QVpTRwIdomvdaqw6r+GDpQGVNN
LFnQLI5sLkYlrRh7brYFqRWVor9wgO3336ZgcvlLGFwU7Dqd0otH67Zh4xFIKwmP
cQNfSCuc/DM0AJj+k42dhZf8SOEDNqDUadFEjpim8GWt3Je3CWfO9QeNEyaxZdwu
HrBI7U+uQHpIs4QDsr16B4rY2OPgOQ5Mr8ZvIaGT5t99j2mY6wSCv6IQsypokEWP
OEfgLy0z2d5fD+AT4d77twDyKRFykttrpvSQECoPDvTs1D8EH+pwWR3gFn3yiupw
kDYUqHn73KUOX40IEsXG0PR7RLVLKa5LW3DNOpsgcNMbg9tt776+k3p+C1c4Pu/B
AuFrxPI09iK6jx+ESBg6B4U8l7P0hC5D9ug1AuaenFa0jqBkGZYELnuIcwvZ79Rp
aa4MW2y66fQa8nCMvgLNq83YI4xqrvPZFBwf3Qzc5XEPrNhyHXsZIueskplA02kK
rd4DV3JWPvWxcrbYQn8MfPpnOegaFTe2CEe9rquEe3+Nha0/Xvy6VDhlAirT1i/j
kXk1d6E7MNCQMwS5YGAFZsnmsFnrIKyOV3W2JpMkYePHivKORLPRDjRNtPpQ2GT4
xnuf0AAlw8+TJfJkHX+Dqd+geIUW2smpj6y0aeWvAFnJi5PDPzRvHDFCooExapLN
BfjjQwMYviXIMlPhElaB01DYhc/gITtddRGGocHvPvzOklyn/cq39V6COkLMmpLo
K6Nuq42OuQDphaABLSt6bxDKluGn9ZhRniAx0IIFb+WTnK/BmVteeB6pR6WFZkDZ
Qlca1WR6oCVMVu14DLHaDgKAtbag/pnX30aQ7IILPZWno3ByB8bz5iq9UbEEPf4A
yY03oto8jCHUx7KQ5r6ValBz+04fwflgWDTw8fHtaYejhs0xoSWQ3REe/vHy/jN/
NjdLcz19U3+bqi6GFKkD98mcP+XnKSrREAtph/zGf9hcA89k0ntl0fHIaQEQgnaU
LfVkyM8Q8hjgQf8Mlwp9rNJ0MUxVygAo+/slHspXfZACuwSsJ0/IV7RXAhwVfrlc
txPfH5tmd5BhKw+BSniuAkdKP+DyEpJ4nVq/KyNcuf+Md4+CngSQe6Ac8GZioQ4s
2zGoJb5l0x+/fZnQiUFAdbJ+Zs0eOSESBGdyCOH6mcQujm5K2TGyyM/lS/ZFxXth
H5ZJ0GqFx07PTa7uWelm5B9HSDvqQjB5dduey3NfKI5pHAh++G9naJBziSvsxOmC
pLJ8PaKA4AiyBVxI2sPrPdH8323YfKhHYYlq8OZDOiF8GyF0ZYGo3Pvz+lyL5AFb
a39bwo9EzIV+oPrPqfgNDhTLr1WGgAwtV2pRR1GG809z87k0wblzT/E0SwOwGNy0
YEnSoiMIip6QSJyla6pU8X385yN2NiItY5bRzkI4ZdaLzdTrhRF8SCV4DlIcJFWD
IugsmFF92AoFO3RfdbU7qXoKEfQEbAd7VKogSugXLvmWEtc4hiFbWDe1WR6tKW4f
bvAj8TtUbmvrh1m7zckxtzqSJ0aAJl1PB+RJtSlHb8kMahEHqVZTsnSH1fZh6Pk3
aIhdR9nNWSbHPEwZtL6IMxT1f+1a4LlCXHsyLHEKzSSCV5fF9Jx8WO2AIVp+jlBH
GNajrhacdfEBLoSYYV+XfMAkeUVouMPamvBoXlZHGneYuFqvU2nhfE32Hyie+vIc
5c4pXGCRvYH7ZinYYdYshiy/kq8mB4NNjQQlLWVmoJkjL4UjIogr/RTPfKBD2pUz
lbfu6OnbmJVmIHvjqylzQm+osiMRHb7GiNcpyxCO0P9L/ZWGkwTquqHM2Qh0VHZ+
yaARA8w94r+MB+NfbihgWr1ViTd/0qJkujulgEChwKc/9THOjSMz6l2inXJCeiuM
nUPXPnGU/cKxjzwUniFd+z/duEanGKU3kwsjY+gtReuxsxXj6HwmxYekqbMMyw5/
X0LajqiBnnHI5JqNHNkQ+K1ZFfcwH6o6rgMcmkPEhACzq4bzGibMHMp6utsyffT4
QoS7dSvuAl60f4i2eYhIbL7KnjG9gabinEnVgBPMul2ZYBaxbe+/S6zMRXMy3mzE
RtvGvTTUnVALFiz7AsNpY5r7EmkszPP0k+LsfomrzuSRiizQQXUzOxV3gRHrl21y
1YQ3USvdE8Ttv8WLhfwsPk8oKnBi44Zfs9+wmAqpcY2ajGgGkY9+UASNkEjcdQqm
peC1RtxH89Nr9EOQZJwLD4mIBKFvUYrHOo1lVOz5lhTxRB8r1sebi6GIijIKLuk/
fiZqHt/I/CtORcCaJanp3R/yhOcGXo7FFPnxEBih/olJ2Wl4zVF3/G8kZerqFS74
NU0bEMFbh9vTrnxdRwg40NbCqqTvxddcgN47mczHMmJGzRWxEYcG3xvVjDNwDpDe
jfDy6BvhUEG65MSKfwo7Fp0/Z2EcQGstj/A5JpcJBBpg/BY5sxnbsDYuggCgTiSi
DDbCytdoDLWIh+H+56pbjXnjGz1hC393NtAZmb6tSta6qqTyIzELpM468N1WDdlk
KaMaECUnIyaJtgY/XyPPg5wRJNN+evc7ZBGvDj588kKZ4jR0E6FEMPT/XyWtoMPz
eTjN0JSm4DtImntehWDxffKMveNf4QzLNpGJhezJYJh0FLzEWKscBnwT0TTSGNxo
v3MNTRleSY82uHMD02r1V0+dYI1Us0VqSrf+DSvBo4oEfNM6DtIPqWvxdS634STH
tQs8IpuUUehKZ4Erf2+ckjrfYmB6UP7kFaMekPHZta8pcgc6+RuiB8i6tWlZsKN4
8jX365XpK1DEg2BRsHjDXRFP+R4HVV3oZUn5j3qd4oOG6Y3l+Lz12CjewP5zlNZB
mLCxKID8Ium/bTqwgCz5Hy36NrzY6SBmia5ceS0i12SUWF2+AA4Q7+DczOFPTAEd
p8jEIoOJvODsbmUQSiNySd3NSdtDgh/eE6IhJavgJ+gDr73veOkHvwBU7Gh7LaU/
y2cQ55xmyBBSVdbRfFgXq5PMPJ4AW9rymShyN/RxgQfLbuRoAObRlgBcTa8tg+4J
DZHou89BhfJyK/cLZVygG9+QFwAdpY5jmbfIJi2oiv+/fQ6hIuIR4iK0wUeL9Yhh
QvVHE4qL6UQRpIZNfVh3/xmw0P42evByMdJd5fq9Rg2yMa8WYCAHJf7j4xSdsq/p
2OFEljgxUZPUdXCDqJ3Kg9eZySuYhqJ6ikC/f7oTMu++VtnAOr1vhpHV2Qe2uFTt
KPc4IdPaOj6CbKQYKTerAuicYZKvDc0eAwp7j/u+Rw1wP2CsNT8iqE4lVNyTDhJZ
MhK49vhByd7nKCRObHD/259Qd7iUF1m2GQFMtIUNSC6OsQyzbWxEd+e05RMHmXcL
7OosKci1PW+hu5hD2xWwl+kOjiw900wpGlhtX9qEcxNd7e+3WQ5lc4lXiXkKAwdK
Q0ccJ0XyxpQ8+e6gqYPZuSM6UIiLAK42SdSg4dFM3GrRdcQWZXx4J9tZeffuk7Jq
vLGB2j3Tm1jol5JJQUE6Dzi4Lr7O0RKCbJgWSQ7tzFYID7Oj3IF+S60hMdgbd1Ui
fEAJJI3CR/b3dDx0BXzK9xmlI/mesI0tx472ZeWm3V6reT7GBHi4Ww6g/gMBmhQC
MFrbwbCwFnD0X+4CrqF+v8DScsGjamtJvacicn0IW3JlDSntVuEruxcfu0jO3moZ
GhluSIreHlYzqA+MM3BPfp4q+6sXjJVq6DA6pRvbydjdPngQXyg9yjzTdOAXE4Te
YtfJhyABhUATLRe6dUbg4CfPYU7xGLqe2l/z5oE7yMlYqoH3xXIPWbBkbb9srR3a
vmyQuCFAGrVRGdc8I4Kkm5GEOiBt0iP9MxwOyd98XtmFvG3L82iOMzGSiLBLlscm
K/hIH/Y9h2aIge4KrHlaHzTmUuFhOOfB/6nHuo4K1/G71W1U1r9cHDUz6ogrQRFZ
kdEyoKb7vntT5G25xhbDJRQ1HOxjdGVxsQicA62sZh/C/Ht6IjLNeEiT/s8asEK0
jlwCDsWmK5AhafeYuQNsDp9/1Q1u7spJ10UFaise4aIVxxwJdBEgrmBDal5w9j8/
/9ppWpEhdHOxV3qVPttfSpL4UViXR8S22f9N06OwtgiV46QrUc6VxP02ia0NnXjB
0Ns0Y1/N5phjnWX9GZBYl+kAXF2F0tYjVJkcDoMPz+A5AbELcYU28/uEs2aBZgDh
5PKK2wrxpLCQA5opyhDjkbc/uZitwEq57HNPZmwgCk0dZ0ijjQgUr7wXguI8AwzG
S5bHc6WrC9JLjbIzl0qHpKU+lnrx94HBIsH7uIp4gf8qzMqcZyQXmxMMPRTyzGyK
gec06ezn42T0QuGIX9UlF97JDmGGxpLZeGTqZaw0XnItptCncUDaRbG1NXlGlTKs
7oOsCdjY3zS6dYJAvnyALwqCi1g84N67Us6re/awcgmQO5lb6Ns4Qb4yxp1vxsaw
Tl7TfqaCb+/+COZ+NQp0fAz+rshag7WNfWqGg+dItEHoGomzjssrJfRQtoifeHWC
hMwh3FfVVsmz0d9+uE9x7BkSMkh+rG8sO50Tpag6rVO9+l68g8fAkBkuX3c/E8UT
dUzLje58bHPgRhYIaIzuDto0j+x0eVdlFBralZRTLnH3LdB8rFncpGSyxaZfkUYk
7e1x7/clMSEnpDrRzWmtNKTr9dY9lhghL8gsZBTcHvCAf9G9xoZ9KVkdjtvXFZHj
D4FrNF8eHDDFtuM0hTLXMB1vigrm4JwS1oeishxSyASteyuz/x0WY8ucxQUm8wn+
/LG+njM35VpBrKV8F0xDK+AtEEB0AVeWi164jHOdwMeDzgCkoZ70WozygTZMWctA
E2N5KYWKkiDxDJ1xWPh0ta35Yoc2F1/kQUn+JHTYBCPF8zrFyYrCY6EKbhXHhGBZ
iukW4Eox5IvvCgHdPkWdBR0L2VVVY+n4ZDBEipkO6x9pOJbyOfMV7TuRawA0dGWc
9rB2Nq2FQfQpKWWeY/0hlM0S+g14nG5Blz5XRvY/Jg/2fy4PhpdM5Ph+5s8y1ZpH
AZoJ57M5lQVw2thU9o9Se33xMkBHgtbRYs3aZZiXRbkubBUcHOqgnSYhFp19dqTs
XU3D0g+qniroli6RI9NE+1D5J9PHA95A7nLa9yIWx0xeavccRccFzbKHbGs9+XlD
7FMU59yKf0XQh1ur6GUd6CdiAGxn9YdRMWobv8fMh+QUjmIf50yGOkAmuDY//6QO
Q5u0l+ux9CFciYYB89BMh9N0Oo13cyUVyrkxDnSlVeLr3LcA3OscjvcquUL6Wq5N
Ua8ZBqKcGYjUBw0TOqmcZj78Jj6Q6ABIuJxlzL5O/Mbj+MwS3kQWvB7sgURa0RP9
kLLQZolkGolRMt2uUJTcSCI97httF1GIKh5z/MXLpCHGJTUm+ABH6w6l7NzFPfU1
YcuLcgh8Ld2LrxwN3dYJK06LD/zK7ylCvOWmOjDH3wGOzbDyT6S2dmRCnDKLCI51
+mEYRXMNrSTkvpZf6dTG+WjahXkQhw/f+MRYxjPx4QSejHkWlPnOxqXs7+Zs7yJc
ZJK/6WyB6i0vd0YkFjgpCffhbkKHygAslLN2PEpNjzQI9B7vR2yzDOE3RUxk7fhF
a9sbbAJr8rY3ZN00FB8pcJjoSw/p6jCl+AL415gLQo7oBCcgZeGo1ZUI+a4Aw6IY
3XyefECn4nwcU4Xf1zIMNJjjcvetp020ChBmAVW4nDVK44iG12/KAwzFjR/9my0K
Ui+RUyj4XPkH3Zl8CLxOaLRkyL7SqjxN76ieFvao9kfP8gGPldXiyuhvoLmkmLl/
051EK5zYKebEqE3p5yK+uvUWjvq6iB3l76yVdB9GLuWQgRigX/kC0E87YJRXMD3M
NLNTaPtIoFK5eGed64XB4eBipEHFidGSBQN6JBlBT50S47IHdyc/ROqR0rkGwjeF
dVmQHmePWH/wisq5kQUMFtBwoIG5vGWD4xgH9d1CJ0n0MDsS4O728VbgVpT5H1SI
4jyPE89GZEFJmHkinj97KHV+8MpKiKq3DXhDrdzQWADHz63VZNKfmYEGzrBHDY2p
aDGORDQAWWUPvzTg2nkPq2ftPgpHTmYWtpX5qIsGX0n/pllOZphWrqJChzW8MTWJ
TycdQ+fvgVfiEvMLbDRKUnNtUn7MjEoLZaYX4v74EUJe6AHRYFIUEQPIfA5ovtN/
0RSztWJn7Nn9pc5E+ZtMn5FHLlCT3ViUs3eHYMRe9ofXfrp4nd+1mNZlnQAMf5jQ
BbSWX8XuxRFc93C5iiURPkUZSP4p1pGlTInX5yYYDT87NjS15c0Hyu0pZA5EcGSH
aZv2f7PP5ZgKfI0uP4E8rR0lAG2z5XgD+Hl5Dy4IgX14ZwiOdniljkKrxRZ+8+j7
wrrSsSqJqf4Q3iMVZjxoLxkhsCrlYsOxgJc9Tnq3CD3ouIprkOB1stW1gjYOLQdw
xUIpytKD1s9/sWc8fGKCYteGfd7oLrwCrNTF2yBLccLqgLb6CmgwaG3Lc4GuGH5J
UxnVKsBj8BvpaT7Gu+A26xClE1xNMWqeNqT/AmbMhKHtwzITsBZDQsNzAsuf79ev
onBF+rJEXfqeDnMzsHJXDkOUjVFO72FG+y01618STDOM7CMROkYthkfb1r9CUhpd
ZPPS8Zd0mkd3WGWE8Y7W97FktoXbQtewX1wuw0nsfbthrf9+fFJ1/YmEbvSS6qUs
AMTzA3tBorgGqaCzx3QhOPFddHK73BG6V/mMBy2iy/AFvh94Sbc+E7I2Fr7IbOHE
DV2dIXaxLWDlESuiCHQfCh8Yt4GqYIIoEhygIP+UlN7miCGJwuWuKZVb1BT0UR6+
oJW+Wy0+X4VaAaeW6A3OVwaxYS0zCymHs4lmf57dPBHZr/2kHfJ5+TXyWXD6LkE+
aaV8Lg5KkuwC4eBJlCMfk2e+wPXGRyv8T2s519atMeFckq2tk5+j2wHe51cO0KqY
6jKsji4uTe803SLxOX6Xu7gbDBc76RFXvqtKmGJl0mdY+aq5yk8MIc9LAOLLQm2P
u5ePZVv+awAMmSdXdyRauR3JDjpeoupIdOWjOwfqy41DLdYvqROO6kVhr+4vkd7Q
wR6Td1gnFaCpgsecbmViCunolRQxNd+HsPuxancM3I9JQPaz6HduB/E/2iRDGtFB
R+hcZ1yBgME4CkCcmKjBSN0ciwxMrUoFSeRcnDf1G1bfmQmZ0sJLffAn2ZENU3iX
vy0f9PDDXHq6svq0nMxvfGnoeO7VPvWDAtKBAkqp9eEhLOZgdImesnMkHt8a5CFd
JqzFU/pvfzsNKYK6JbCD8Hk7Lrv+4wYMfZaDftmfDFF33RKWu+MRsFUBmKVK68GD
AOIHw+hPXLGF0SFuzzu6K8J1RGtdrnxq0Zf2cCBr+PvaRCjF08RpV4fw4aJTnGj0
USzVOlzDnXcpAMAjxj2fRcHPNxeVHA7CouUMcHjlhxgYeWIJ23GyQXhEDxsmzqiU
2F92DNIgFm/1PqLRMSAuILbf8kfUCtsFIxIexl4OxKgsce3zaQjt2cADbHVHTLNI
vNTyFkoaQWewqI7H5FW00WuJUIPmBhEE8YEpgUCJ7hbItuULODULv1N8MkjMomHN
BUyMx/7CaqCoy/g+Q2HrDNfVZPGd8xS7l5054dlItMdGtvGuvkyZ3tk9j2ag6Dxo
sMDgrrpdrViWFLqAk/9UOWNYJzsbUmNnzmPZ9EDrwxKSMHKMSVa0kwr2VsobMkHS
v7gEcBL0vLWE/PQiU6sPO6ciX3QCoDEIq6AyA9LJAI/HwTNYHXc7DYil+QmJaMwj
q4dNK/lH7NwHCqIdl21O2OLj9bHlMLGpJazAlBnf1OSms+nOh+yw/VyAtoQlLI6Y
EHofty5iqZyKTr8gbqxIe6Fwj1i9DeXU8R8tnIIEGEpULtMSzTD61ANU/jN5pQ8f
gFP7CxjTvtmFDs67YwEi9VL7ohPoFKz5PVprGXCT22JuobxvX4wmDaJgTYFpuGb6
99nqOfMU17UfqkRq2wNfk3BwKogHQyXKupzCiykP2+cRV37DKrYRwwewROuVe2Yn
FT5osbyduo0jqX4zn6OOamREP826bHQ5zzWKJBN1Fr5o8tasCFLgR0KGlRSA03DQ
IxsUOrWvGYoNYE3nEEtE87NrkNkn4q/ZJ/QcH5LOftklrAZwNIZgLN21PujbcBP9
oYz5ayKjX4lqHCrcmXe+UZiX3a7j1nIKg3T5wuQODlpb8pTG/ntTycaf/i6l64A3
Sba9aIIjL1p6JLasGMxaLZSHuuxkpBTIHpjPdTSFCe/nsPsBwoW0L0F9NHvkTcmk
4yqvgQSHyaXsYrNBHXE0UyVJMil0UL+nhssbnLfqfZ3qgp4xoVZ501dfdL3qwhgu
31uL/xX4pVcEIxW51dGEqoNleI+rjkX97gPT1xvyQi8Rb7NHzA4DHWdA5A3y4OEi
vP+8xpYhJni3oFT0qjr5Hu7HWtrl4y3iJAECt/Yk1744nNS3iR3f5bAEImySU6Do
H8Ae7kbY3JgewaflGgavf65+xYJihMCJWY3kde/e7NicPN5rYrSyuEvzTg53Wlt1
We+CjILUkJojNj/rMqYNWwBR4dr3v0VFUobAiuEgktZ7NnEDUvWE6XQAxjO1D6iB
XVvyNpdBSuvCApIPXdvpToETpQCbLfqz2f0D0erQLen8Hojqj8EgWOetps4itf9t
oPUNjVPN9mogCHlOOD3UMc9ayjNjf1TvzvlQDZ/dvxfG7NDRdNniUufRq2X5Kn86
6JP4u04WpocQyePrrnTwjqaeMw/7nOgBg+nuuzPjMS3KRY3K5yuLgzuzriJyxB2B
Y/1n4arINnYFSgXiLyL3s4MzBjINr6VU5hY5CrN9t3AyMZ+PXWx9QU4t7Bf/nstd
70TXHWxxj8Vv/dQLtuhQgzYwMQ92XKo+l0iUotgHvoT/xupu4asq22WL/lGXeHzm
A2Bxs1iGz5ru3fJhfepNpRxYziJ2uo5VUpYkajL0wohcQefVILuOKqOVkFEq8icf
8AqeJr8sowKM239VmBUHNFoAmO3ONiy6jOYg58OdQ1nK/rLbJpseo6E+1JAZw1rd
FXIVt4VpdZL843RjHiGP6PLwgpc3jA7nmPjI0w2rNfIKstQnxQruy71mzgZtCo7u
x71qMYvp+meeg9WzgY5hiZmwV0QYY+5wYjUKMaJk3xibH31T4/89ZG0zyk5ZWhb0
uAORS/l/eeWHOl9nHocBLNQRE++fbTpGru35+qy8sEKWEXkkwpog2Wp0DTHKUUzY
1Mcq8vj+nfk32ey3hGayVB038AG/b97QeB1BI84bNjXG6tbcNP8MEXaWX1Px3ri1
H+KSwxALCqgy77SfsdgNRofsoEHNR7HAbo94usCKDCEhoAyKFeakt4qXuzSZpJEz
l8oMPwLKX8+sBNrDDToDEtI32MkXGoeiD+CCtbREl2/A9nLp+wmOsHa1rVu1LqAj
weO8vxIexL02pAUXJZ6d42Lev6TnVgZaYYdN6+hJ7hhdaJnTFVNYSjsEXv1I8E7g
zK8B4oYnbQHFU/kvbI7LxymWAoDBEgbRrEbpNqaBzL3wVH2xSea8ZMnuhVTbd2++
G1C9yZdk6az7/PaAJxQCx668PJWIDlzj2aY3ivS1rWcFXWSZOns1Q7ykXsVH7vqs
dfwYOXHVX0vAyiq3xg6jkGoSxpWn5ymeZNCyFhwwKI67MTYuZurnCZJAPY657Ne/
ifi81YEHJoL9E3ll6C95UA0upOr1NSbanqtvOQbgxPCaJANZjMnExb6pVWlMVdou
Zdz7Pf9BqPCKMgx04ll7zCQNtJdkLUC/DgtxI2lSH/klska99NQv4apHXh2ovglw
zQHkBUk2yVKW3IRQ4+JoCSA75KFRa5aaOw1XbmhfaQkTGsoVn0zoCIRSl8bfO6iu
gmBb+cQ8Br3tiHRxtG+YqeUQGp6avOGs+m0Xnaou+cMH40i9BwOsxe21vWEv0Mn2
/o9/6jC7HN8/xDqLRfKxWl0/N5B3aUn2TKsJk/dKKmnK0oqp5BAPXLdGEqyV2RsQ
ZM+UATN1gTYsXEj/UJMkfdnClMNEfejZiIIeSxeA0kF07+y4xoqKxKjY2+jmtzfS
ADOKuk5Q2HW1Xan5xZRs+GTldD9yrdZz99x1eE/X7XZDFkGdweUqr8yv6G9dtCjD
a5Nn5ObnOXytlZYataP4cGZRlG9Jamu4+B571kQMjaPxlOrGHyEXYRD8pb53QUfD
vQWZATI+Rv3aRyJlcBQFdwvvuuQh7eQHbiLqL7NzHvf/p7ytuEKLmT09Mcdc5rKS
2vmp4YKvC5JOrPkbLt6Ms2oOFqfTIVgbzvHdfz21FXE27VBrzyHz7vUEWuJk+bMa
GP7hiBFuRk8mStgvcG+Ujep5PUVgXhuiMg0Jc/uWVKM7cbsUg551pkdcmDFbksm4
dbsOYUn88aA/m4AZzxeQdzMfhZ5/fA+rSCl9y0h52IoHOrn+mCyF9EuZwRB5PMIx
k4C0+3FRYjZGaVr1me56bj6J3S+K5yP9QVcEkFiiIvycfhtNQH7weZorhLNsWd14
UXvhVUixKAW8DRkbK8spwKsaLyiJvXYWEoq8TYTGUpPLJ/gghdqd3cnhuiOJaRSb
n9WE0K1EylwE+qUE7H47qoR7s9vZCSpq7Mresd4llmTV3od8ejlG9Sr3+GxrehXh
jF6KAe7zsnXOxp6kNkatHK89u2PhMWC31PNxoPCiWy30u89Yyj02kDu7hUZLJl+3
J6UA3SGMbC+w71JqG3hWpS9ZDHVR1QBia73l9P42sTud9ZCWlRDracGBWuty29Kv
ZO2/dbpoHNekyYDCXlmNJ3+QTN2A88sBpItGGwv6E77Hig0OY9rlQbLqpnfpTga2
2f5soT9Iv56YTBomOa1fby4NRDgpbysxakaxyW34+iqY9yIgudTpmVKxHH+6lRpE
EPUBdCdlN6pmX12SR/hcELxxdzNbI0jP0m2TeS+TEVwJd1VIVl6740I8Yz9R4XlI
FDtYSiX5fkc8dlf1SHsoZsuT12aGMNBVWcptJ/drx6Ti3tltxpDXAd7erXrUMoF0
+CZ2K6H0aaquKsLYJdZXSS2y5WYslGaKWu4CcZfbPDKGn1XFqdlhsCOfd8FsxS+q
mhpqf/eykCgDbrjJKlacJ4k9KrAuvdXl7TspKDkcPRSTxBC1MEgZkZtwWS2Z9Shm
CuMkTUiwiIByJz0RU0Mo5EIGHnF3NO084VyL3f6J7Vv2RROVlaUzWGIOrGBldp0R
vT6dLZxx9JWScvN966oZkYjNfeqmyu/EnzBJ4XqmoNjTQGYFp5Flyu8q4yDMYDmH
ro7IiiycyXINxqE9qD1BcJEXvJQXOV105XDswcKIQZG78N8d7x4y2t4jGt6FaDOj
UJpGMFW52eqCwhyiCZlH447Gm7nD3Hfbb4alpKnTelovY0YdYpcCUIHOOXAzU4xA
q6tfvvrvhdXPXPT+5UaUcPVmqGwJ5agOUXcGavjEVzk+LhqjC5hbnsvOOxZ/C0r6
2vScO/mxZyCwZ7dLvA8W47oKGy2jvR+o0ZYrG2cZmf/FTOoczBUGclN5obmH2I7A
Y7eDJYr8N9FNyOAgf/MVODaBQIgaPKGghEHt3AMfeSNqXx1yERxMiM9+lAKrS5DJ
CNwxkdEatPiOWQKkDchVkdIp5ZCYJ7RcFpWv4c/8AvfW9wvoPH6hWe2+Pf/wuTWw
bwd5WP/dXPstOBkzQdmaDV0PZSrHcSnY0cZX7aToo1Z0ocnHFEL7HQrWrymDQHvU
nzAWv1dF6odZmdwcxd/27/NZpNaQYzU5yzIp+SLw5a+g0S9tjVkvAAOHRRlVEpEe
F/L4Lfm4DjiC7o5xXfQxFoQPAcku76/PisR53LoEJnINS1ZK/kbHbvEX2WZVE3EJ
tRwyDdO1y6OPjuXvU3cbjEZeco++pD8jARVK7mf4kiTgYJOq43kcWPk6lpuChKB6
O4f4A4CrvzLOq/yJUoQhdMqVTgSKSkrAoP0MDoprM8Auc9L6WV5fDGjiWsAgQ0Qx
3/y+w8B+d9R0jy2kLwZhK4GFyMR41+jEVdX6Qyu+CVCROeTbrR7yKWObcixUGbOK
9xMljYLtUma3EceLoPw5AqQNWBBn5BRd5YeffI0x9twOuEcE3fzHAURm/hSHMJPT
qGykW/qz3HD8gbX98nhSkweLb70shewH9VySqWuXE9lpL8KGHxDDeUAhgFnE9oFs
RQthsofGB7jqrA1Z1VcN9eA7qOisW1+3k8uKGNVWrYfAAdKaECtmnCksgFge27oI
68g+h3MsBhQ9bHO2e+vAF7uks6hkXH7J/eqrFzbqcX3d/dlr0WWyG0w8TNmYBgb7
923vG8NHGnaqrRt8qkirndRpuG/7X5azH74+kdZC/sjhFQAgJT3xVfd4f3EaQS7S
9yIbVapECTPlqrvo64geADDkkFpIA5VhywV/kHpuJqGB88hnavc7LAX+LpRuoPK1
K4buKP8nnMzwn2XCwWpjkcJR2odLpIROEipkGxc2vrG3R2mnK5co7dt73M9prAG0
SaVqgAdHrwEzPj6dZHveVCSQVZyj4483codTK0NLpiButzDZaDzHSQpITDA4hXuH
qtiLkl4/3VDy5BFOQkNNhr2xNFSUMPL7z2A9ZUA2GN60oRj+B66UAWpETPS+syLw
ur488zfSkV1ZWDg2XoDHYbTtNUJ9u4rSeasdvEfdwHCHUCtpSoNLczFFH/CAyI3a
4wXv7gqiGSJ9XP1JCVt9L969NLWx4AyWPZQ9cqa8juYSb9PoMAY+YF3Xbgx6yul7
lrzDoEh/OR0ivgQ/e6uG6RRrQEm/H6Ejj8PfS23OLmEBD3moXeN4BS1QyAlLEhIm
kl0Pbb3EbBepmeBqKqQexL1tY2IHO4a92jstJIKArPcqcE1a0/C4A52nVHF+owCO
xUv8214VB2uV84mh81ekORhbS6plxbalIIOF2eRvQRuKNsVn8JWrGMuxWFvPM9++
qJd592QyCr3rZ8eMo0xsjNkyRP1siLPFhIKByclRaI4whD1k08nUpYt7OX4ZrS0P
PcALMmuDApQyW+3AD90DZpYCrex/6i8BZqTBwgZCokSdP7XdX3RhsIuz+lho3j6R
YxPjNKvW3FDL4KsS6PTYlotdEEY7vH4rp2+ZHRhQIIByJTtOWjl3V40xWWVDfl3Z
1uAj72/DGJjvKCSdE9uM5V5EQvv1wKuroccHtrg0dG+nt+rGPd2H4N1ljmSUJqKL
+EOP/JykCSKqb9Ya6bwz0Cl9Jqc9VNIv2H9wfOrI/U/tzWuURLgQ6gjGf3kTkNAj
nWnfqR3SR1juiAXClRWdBXwxbOZ/PP5GDP6QPTM0X7WUNgF84b7AlOO9U3sGz+dD
AwKccul1OcVpbanb4XaXy+VuoG/btCyW1B5z+MDgawDVFQx70TQrYlpk8Tvr9BwW
6O2MG1EH5OiUqIz/Q4+FoAQFJY1uhe8A8gKXP0U69l8wJvLahGuCKY6J1OrSvqYD
/KiIUTJH9cBTt0Y26/wcviNmeRBUfOqdyf/9dmYuMlnxT/1DuInNIqY//7JHcI0t
IRiHCTSBU2l4aUGcNX7xZ+jqqKlMR65aRknE4EhoMN9kNXiCycyY4GCIbqcnTOVS
GcYLRphunrTQDujv3KC0G6VJWcl//U5GBmybLKtWK46iyUAeiFXZxeBR0kcx3UCs
8qRiQlGiui3cNaMr8l0/Gc/eBSP62qOdDTW+c/X0GiCUFnPyFL8iturIb8jv+O7S
RBCeNVZr4Ft0Y1CGSzonU/Txkm9RT2PKcjh25b9wXFHZGb0qd1r/6q5EPFt3xc3y
1s6p7maxdsSu5/KOoD/LrX4v7epqzr+qvCEeFFaM5OytNRyllqJkAxA0/q8DyfyV
oasHpRw96o4g3pfNdNU/gAGhjOlatCSY4vABALzWpmA4LAYe+TFgTVnpdEwtyrSC
NlyTTLmnwK/2IFnMZSQYCZ7Ie5XxoYAMt5dih+GEa6uVflEHRnS9tOb/M49ZvfEG
4ghPW22wnLK217Y0iBmFZTeLf8wO76JMF/r982OW02qvVoJvHRbHAdbTYoeP+6xR
XztyKwG8u9/rwKqlJC+W8ewhWyG60jPG+Nrp9kmddqa/bJjyV9mfkQOj4bGbBEsR
K6w8RCIKzGKrPpKupWS85p5iMpzVY5VT/+YREjq+bEktkyiFo9HjWZ9PljVjP7IJ
WGfZ4TQOhHLmw9WsQDZfnqIyictOv+0OliyV/xqTiRxV977ke8A8j2lppxU7tuzd
b+RC9NahMiAer11SPZaSA6WBnRxsppBjrHDs0cEfVgFsXL6qYYFZO4obhs3ZMRcr
2GjwJ2MFzWmHUKXSB8OLmrWBpkCe3lrKGWIBEdphzP/TTscoTITvel7COHwgiQbJ
ixXC2Xy2T7oKPlkqkvd64JI+XD62Z45HtCzo3mx1a+FpQ8mCfyuvb3tD8TqBDI/u
TiK4WAxJGkeMmITt7XCloYxGiNFa908xjANN7spFviRYPjzKagXFOSb7mpmFQwn+
TlaqKSLVV2D38QHm4XNTBqWcqQ/0WhE2UhDaFQg41GsbEa44SIQyXG6R6nAZESKD
pGGKfrAjXArKSYOxQnoc3TJavnt+zzWN0eg6PsHCgBaxe9vgH5rVsiETKIt8urW7
q54qq1X8L5FQQMuFR16PftLI7AqnQQE3ceZo0YlLIq/AoEMn5Vyw4G9F5dKq3U9m
MJ76llmvKnAU9RGgUbP3idB7szYKQb2kelPZ5C0utS7LVHAc+MXTNUDUkgNP0GoB
POKb9+nqfL0zMV/wdvGMO6JBib6ggkm69OO5kae2yKmycMWX7Sa4HmYK96CDzrEH
VmlXmmpoBQi4z0vEdX6fOd20VS31lld1Ilv/pK19yHRFq0sKgpnPTF9PV9YisNGJ
pujvCstd153QiIHFU4NAva/alSsd1IYTS2JX+swEqSqlwWbNYREw0mCqnlvOMt02
yb8XEivH4i3QJO0EdhINzanepM+r6wEsV7zzzlhHxvMDkPTYG6JiB8Hn82keRYFH
qaSYPxY73jFL4O3vksb179zEg1vbZgfp5Kvrj78wcFznbuSMctp0q5Ho9IBvJtI7
w/ZdaBqRHRPfPEHtQZGyqjdeFANmcHFJb7Ftxjt7yphkKAPLDe9p2Ruc2hTxIqlz
GS3cX0uby4LCjFEpsj4VZmhnjY8BDLWES3koumOGOnLZeYjq/Y1TouEj9gBXI51f
p7USYaS4vw8mhJ7FnG5fIHVkG9K4d9PfrGXn2AiDZJDCVtj1bLWhceFatXp+wjiE
3ZEq2XnKjKYQ2y2LK3I7rfHWZZNCEGa+aoymI4kvBs+p3JUJlGat/3YjMdB5ct2e
KskFrfy/phHkkJIVrsWpaFBwO47lbI7Y88rgvxquhvAbXXSu5UjowKNhAI4HGVBk
RluWxad9C1W2EDpKmM///k1mRRw3rcuJaGRHqoJhkE4xah22E/k7nwn/1is54OPp
PMB46hpllNZjpW3wj2vp5VW31WJYuoftaFgXWdJ+k4VSBMLfhxRFAqpQu5LVY4qc
Y9MVs+yYt3QJdQZFXJzqm2FxkEybVgLxJdp5sk3XzWyLks0fdDskBtU47Pe9YH79
1kb3FZVVDwahsr1j0S5NLhAaEcLnfNhyY2dDWUkXPAGyucJW1ecwOd7cDpMCtsrK
xxnBgOENBN7xAEN2jIHMSvE8QfUo12XEv6cFKXpz2HET67LWTFsTte6gwGANiL/P
zQz03RjqrSgDLF4Uw503yUxAw3ozvDUbyenqYRsDyagiadkD3j7N3N3Nqv7jEAKj
tTLewHX4qLc2IneNSTigQWgMZAcdOobq7b7u0rO+n+mCaSocahVWANsqf4pKeWAy
zG8MgRnu1Z5s9t3uqo7+jzpj8Wec1IZKkZ6pth99kC2G5Q4g/5lNhAmJqPilsHvY
bEofL1m+MSB66ugtX0VulQps2mSu+QY5tc7Q/SKswDkejgHeT0T4Bi0bCjXuyYSb
vAK8h4ip1qv83p0Zi9gSnhIzB0dnnB8o1ft9ddi0p/7+CxPze3QYrGrv5Ms7ksEB
tFH9qJqfJdSstA80Q/SlTlTc4dL/ZDXZzFB4iyQEQZXUva+Fn1uLwdxqmz7dfnfz
xWab+Si6HPa/WYY+QeRe2tObFG5AeZ+5enkNsZ+sl/ZTE0QEeaITIURHYSFaKZ9n
n1XIThNfF6WkNglRNr3CIzHhmnPInJ4ZKqnildda2YaYMSi+hoLsPbKbLSJQcDAb
/tacmt5zNWOODDKnQuaCttyo5n1KqwakdZ/TqS24apc/xUNB3USn9i0ZDdOmvG96
5rI57n/AzKWYHnnwK7eonBBaYS2Wa8gFTCIqU5ly1GH2Amk49ZhTc2dpJnMWoG1u
5MUhQFf2wM53vOD/ISvLuRKvoRLk2Gvt5PS8sULXMw6Uqs5zF12AXIv52gbWTN1c
LBxKghwFNj855rL7MZ6nQBDAkuGxkBW+18VtwF7w4d17Q4OjwuxUklHVb0dr/r9j
7PEg2QE9xR+GXYLwNq6O9eMI5M6c4KnJ0wISbuMx/PQdJoHY+swemK+3pCTcK0cv
pAX9Nt06pGGbBvENGxmamEetYUP9yBitmd5byPxwjWq/Ln/s4oeG5kpw2/06WJIR
Z/mq3M9qxWEKkfJWiPrzosOgvVZg/oy4Zb1iYCzCU7MPnMhkCgqf6XwCganlK7jH
WdhqGjgD41+pE6hy0AqzjZ2kYhFTsGGcoTsZM2oA+qu6re7gJw0uzSeNMPXO3Z7s
tL73yrqdnXOK871yEX3/FJC1+bobd4nVoH8rrlCTAAlfCT2X2FR909pkHDiwUycC
mJg8en5PgQmifd7RVfi3TqBq9j4buDjv1P0S134/xpaDkcsXHGP3NTZAZBo63K6D
dvNWSyi4AMG1wWoY+d59QYn3q2wcngs1HVgO/dM5FGn7v1q1oq7Xt8FE3hqLVUlc
V6kt/cEhjFq02ir2IikobmUWpgKvoJs+udEWSZCBfseQ0Li1qTuJu5FNd9DKLAI9
sQXyYqTh+2DHQYt7zhNpcX0xZHIpXU2RoaBHhb1PPy6TUigpnQDmOZl48yy1ugBX
3szP+J1YICCBu2NNDLPfKO8CLeP3UOU3bK3yImdaR7hxFoO/jrpOYEVoyfTapiAF
4qJWV91nTnWIyKXeTsQ2AmeyOWOHMsnWHtO0BX+hqfBOREWoQjeYlrNTPny9UgfH
OHTC652uBsWMgeO0SzmDlhHacSb7DtBAybDF6+5CXJIfdABQLiQ97yau0fsN2Eed
iV8zr6ibtUg1GUxsa+aQc9iZy0v9IrHPfRJaYOznLjnDvr34RW3WpmmEkfciGDhR
vU7zWJXzfHh8CwKdhWMEHllhHivaHp2hNP7WuD8bP7feplZFR6PLVGl7RlKBNZ4J
R1a1PJIhtDE8rcMT+VVh3022ANBGnSI9WFuUkanWUku63tzdU3Hd49HNoWlzU9fd
4j3G61K6hs1ywsToE+Vx7vF82JDTHbndaw4zb5v37LNe/Dru7rU3ScD+n/6lVF8k
FjNwkv1sLUlh8BpJ0HSsb0JfGjBdm23CIONT1l23eTfcrQ+6l1H+Ukuby1UqRBGW
8j0sHHiQAb0H8LCMDtajDDbGK3UC0/zV6KbSDcznNTWU3ZeFy+tsm1D0dzSl6FZt
4n+SKBjVDDWMV+bZygfrAQu9gk8Hibm3OlUEIjTtOZe30jJWg2ofoErCRJui7Np4
bv/seidO+fxtQR7vDjwUOoydC2uF434T8u4AiDziIinOxu1FX3DO8/U/eWH5mo24
sa0IetmZQQ6T8g8GGvPaEREj9Uo9+BoVkeAq/27Ha1+OQuoW95robUHvSzjHorna
DCnhKoJrm0oy8pjBfSND1WV81Mgx6FI+sY53xGdAxg3gpZmn6s8eCbrtYxhC8nKo
QIEAPhi3oUSbtOPwtlnPBczX4rQ1D7nC7CWwdtDltcbyBMEL9tZEOgis7H/AcWbJ
RF+5rBYMbwPLeGFHaz0j+J5WuSnfFNEiS+cxX5e4P3KBT8bVcdvi9TTrIPe6WUR3
Wga8OVM1LJlmHCc6kMaKZWD3j52O0S7e8SbbQTkUnqxKsUPKCI1kU/CObe0Y8KdO
nlIv+EzPrzY+7shJXmo8AIF1TBy/F/MhlKfJ8x4HV+/bCjgV+oHlLCrPxK4scmV6
l6U/FgmORHZb2BUJKloNRcxPTkfy+ivnABdwASQJHs9uO+qSWzQdXo8uZ2tuhbCB
ccux5HLP/Ne8CD3KiFn4ba/8MHtyZdkkN0fu3gbYRhGVCcqqT5/iXbl5OcEHyAPa
9CLAA90p9WJASHVR5vCpKIlS/mBLE94lUrx5unW7PRhp7CPa+XxsA6bbGP29je7e
M28YVz/fqOqH9/SNqhG8q5yUhnwEgNwGizs1QW2Wow1+jtK9mKYyndjwnllu6PgW
lQHAc7oHWpoyexOn1wvQBJuZV8s4YZF6G7FzWWcgjlpLlBfZm2SrynsifbVooRMU
BO9RMqTC9DfQECk17F9ZQKKEnxzXcDn7cku3ul+EyXsh3Bs1BUCEJhzL8uD9o+jL
sWdQTQuhP28q9Q3gh2Fwm7yZNc5Xp8ajRV+2PXf7ZI+QgeksTe8v6lRpBOlRrwR3
3eo2qr5/tINwIC+Gy42JWQdFaaC728UxJyKn8uKumCaOWtmMxineAsw3onN5Og3y
h1eHBDwO5tdBhiL5LHVfcIz2l7zxc/b2IZBRzFTRGIKXgszQ5eCMVo/6rslTjOQO
CVr4FP+FcejmupTcCmIUgGlzzoM4YnuEdlVbM+A7Q1l+plWYaICUG3wsiw0VQZpY
LKZIHqnc9MThHuB2LKEINQ9gSQLQLZihECDV1IibxIfAIljz9bbZ+SPN9gLJXPiy
eTQmm96Ej2Zk93eP67xVb8KtgSg0UgwbR22/0ifIV+CzQkGdUBn2bDCX+plJgx5B
XREpxnqp1qsrDD+Y0wthzzjUbW8jCQPEm1/ZT6ooRHZHR5eY9jjJSxcgZKhhOkcr
CrGml99QBfktOskqDeMIZ+J1SpP9me1dlvVRxvm1NyuGJo8ia+s+bzjKOmJ4z/Nw
NdkmQYv0lXrtH7GpfViYrc1p/Btk/GdjBu72MK3EiTWUkwpUr7n714NwcNi1HxkW
hlY9+DDTrrNTl1OI/mFQ31i0HmKDGECYI49KtduOO9k/GysjL/y9CeTV4swWEAeU
kblFd8UT3bpuYNZ7lhShvoKqi2kQf83Lg5+rhJ/GbQ3QHj1AP8jjlcmkJ0jDgeg0
50m0IanL343NvDk5Lwdc/PN6/u8x/f4+9zuDi2WjmAryoOV3pUN7uTL1HBJ4rouB
KWsC7SrZ7Zavq95syJH3Tb5dibZOr+NctBouv/9tvreKjOz+qedM8zwRuXVPMk5H
DoA74G+h22T8SpacpI64j55ftmdv8LK1UDlYsPpEVmNLXix69ImFPvyvwkDKkkYY
RjBrxIPSXVFsyJdQ0ExpvLSk861ZCvW0T8AZDx4JT7fL6ykVVjAqlKBXv+29Tmcq
olv/eGq2wf0ujBXjDqksP8TpcAq4CGQwOMeI3uAsGaE7TgT56pIATwl6O3Hhqz8J
YgROO5MNRDyrphrEGrKwG0/IVMHPCf2bHbxm/g0IcUfLjor3Nnf1ZGBBWTME5HN+
mMPn1a74qxooqfD5lzdTLAlyLZ37fj60sN2/2m0CZvbApAC9aYPFAd+HU8+LkYNG
U/7gJsPaMUG5zSOwI/PnZWyPvexWedgZdglDPB4jAtTFh4M49i72cYGfJ6zCukW/
+fyUSLBxNp9olWWoRLj5ARbX+5d+wBHi8K8JpLjwvk55XqYEl+eypQa1hvWkL/AK
aUTUFD6Ofs5iTZ7XXSC7Ekoe0gd16GUb+xiwT7I+6ErteEkeIakFcV4tQxPhYSMl
vheks3S+VWCsjTYsCmusozLAlx6jHhFATHtEIDvuvvMwV21ObgIL5y3cfua4R+eH
zG2fdUT9LQxkQnscaIaEOku35QtI+orNE+Bgw3Am6Br8wxPE1yM9rPhXWBsCWi1M
OguC/SpvUb5ITZ8Hcmi4Mki+XxDRgGyl2CQLIM9wP2TfXyU8KoppIYcrfWAYlX1c
gcZSKreHXaw8qZ6tqWAZ0D6V+sEFiDzSV/VHkznLI4U6+G9NgjwLuCJqET9tCDh/
xtQHtoIleeeO/EoAsjt5J7h4dK6LtAiKTQI9gcVv23bYNyKh8JKxDtfxzhVWBQFN
L3a+i3xc5PLdfiClxGwuJ8JccU5KYLvFM7uUQVzv5nK79TtgO8B2Lp6X1qznjcpE
1YgV/SAprmiVKPzqGciR4M23TBauytsisVU9UBnK03LrqYhwbiitHwYzG+GgF8XU
GH6lG6/McNYIjG/8I7QCkt+cWi6u+haz9SYZ3fBGRsX8u2tUryAm4RwpOJg++gzy
8NNqQ+O3r9GIj8BVk5P4MVSQ8+YeRPvMp1Aw5+gESCoJWXWf8qU2xvymBPCX2QQy
hlgCiqWd+SYNIJD/pcE7T1b9i9Ohrm/SNqmyemdBsIDDrEr3Sq4eD02M8znE29pZ
AAPgRDGxXunaCqTZzqA5heW4CmuUrOU9kAQbCMhZYjPEKNCZpxPCdwajnCcfEWdY
mALIvQL8EsIaTDKwfI1xP8LThro5bnga//QbwRLboBvzCHmz7JZbYrpGyNeHpxr2
PN6qOMWm+EOLotFoGSw/W4XsZyX95OiUAhGrgskvAYAjAJjWoiJ1o3X7boDo3rmJ
GPrl+Zj5OBTgi6CkViPOdmP1XCuGkDZDEtQOYZcj97ed5GRwWDNVJDapq4q59RqC
R2NTQSjfd+2z1O0VtPkrRrb3HBnc58nYZrdTF0w6rXk8zSPoTdDV2NCJTDPg3vMm
3Aoyt24MrgQM7gFEopmhhJBtFjfb0s5e3McMnWD5I+5HvycE+sfn5I6kCADmARwj
18PNvKnbThzDkfjlsFMlQ2v+6zaW9GHwu7vFRWgYY35Bz+jYtZafKFo3xp85BVrm
JN1D0TD/EZzief4AKDN8XtG2oz++MCKTFhMEuaqR3Xd8HOSSn+paUiSnhznGAAtc
9QAxGt8ZsM0N8pwJHXRFbCDgYqzfDxB1BvzD4xVfXKPUzvLPOey00vMsjCa7v4j/
SUJcdjEcswIdlhizTC1CtjgHiUyhhAaRxV3s0s52gH6yZ/BhVTzJ/lw8TFIGRbSD
8ZdPk9aKnPb93JUecUJFlHFww8a8CzmPPxI3VBzLyPsZkXrpBxL5vCIaJ3Mr+3uR
qGKgxPFhX20VJlzEE3d5QdRmZUYafS3iyffcxsSaz2V/Z34VIdpmp//2Wo740Woc
WB25zCoGkuZwdyhodP7CrcXs9urp/rO6mE+CoxDgYBYvRUHvw2OYtSFllQ0wIvJv
w9vL2xCj1t6qUYRon94uZEqG4NxJC8iph5ENi2K3AD5MCLacqwoOEWVI0rQTVM89
Kwc5z1mKnX+EdgwMDyLDHWT3nMHo+63AfjnDKVVe9H8JJFL+iLwoNKbp2c/gZAtm
spMMZBzV/940Kg0IsI/J27b8OzglwfF9M4lnczEo8vAav7MU+rt5f3obPofUA2dF
mT243iyqgAvNfmc6wLmGvNHsbiO09fLjpfBBmTiMWD726drZ8bkvHeY+XLDPGewu
k5LF2ey/S45XX6d6NaxVU85buyjcvFupXF5EluUbESfqNW8DjbERF+BlbSC0YQdt
iJFM28ZkwAeMlQi9xlKZ4ynE7MCZwA6OiN4N8Ut2FSmGrv5X0n2LSf32dPeS0Pd+
v+sAFamV9IujyfizL98kvHWdZEl54QWian+weRDnqu76WtYHZsj/yI/3YiKmXemS
K4/ICJXdUyzxB8hMtBGAUfXP68hVA9YHJRLGHu4uMuCrTGM9te/WHOsF9JNnK9kX
JgoSodxJ+ELOaxxCPTH/M3OlgIolkXkCyPrUQjqOfEwE2/9ysqXzKPmXLDFF/K9s
nrfmBHo4+e466BdclopFti9FhMCUBL2zhg1XdSeIYOqYc4OxLVvmG0TktIStlxZV
m0nbgULm5VbUS+6LaXqjSKgGMi2o6iJfzqKxK/HuGpVMh1uonvnHff/h4eL328Jq
AXKDNwSAAqOHR2l8FkS4+l/OWVO3eXxkpsVP7jWo3nfIcmOCE24qH6U85/zCQW54
wdHRxp2jHhsgzrhESbbt+VlJb53K6WjEMPQR2waHvP5vLjB/Hcmo/Rr4wn9emM2c
QBDmdbHUfJo6BIGA/3tfb9jxe+BqkBLPJ0QwD4dPSX0TWYCNtDTWuqJX2BrH7C6o
mRqRKGpYlDUbK8yL6qWCRu0THTxoDhtXRFm8Cwecpd8BIaoQc6tz/gS2A1U+VH0u
WLKSV2yedQhqI/mM9chsqV7BWRg7LzJ3lVWoCDentOn2KCnXnlQ/BaUgKZ8kjWoU
Awbf2qFyzrryhXczpn+OhCGljy9d9tfd+TfCbi32GbS54f63f16wghG1xd+gAVIw
adKa9ePc/WWfMjVb4meFRhDJy/lvkC8ayactU1gsR0eBhL+cJG19IuUfFcAH0CKI
m7lKpJSDmRab8g+8GpQXrAUrce72G+7HHJO0GmjNPc8g8in+PnnEJkqX52PG7P9T
bCVmjsJpkyNmDYaLVwRpWqZyu/YveBpn2kLctci4KwxZydzcF6Sizabv4kSYAvFb
77/SDi4PqdEvo1zQqJcj44kdl5H3v+DMcntiobtVP2DTw5heCU2oZ8bKf6U9UCX9
Hjy5hUn10m0ZBParyJLVdh9kd458x6zTSYiv99N4BV6SAzMTu9c61yVFopHeSDAC
thxebvh+61Om4OX3Bk+pqDQ7BBYP8eQUCD+F8NlKUnRlhxzF11u58O6/EIHpg1aF
Qq9XKgS0pMCo+TRJO4ymEL0/ro9wRrU/LClc4zRu4HAVXCsQZjMAc+yUxiMLWAUM
XXgb1qidLmrpWY21djUQrwNAq7aTfv+F9as/ypiaiIczOY9RD7ckIA3wTCbsA7wf
freZmb9f3v5OKFWoGIS8ehK957mx8DVUDmiHfix5QvDYCrdGBRx9IvKsiz7q2gQr
x+0/XP9Weqv9g/59Te+sckIYN24HGI1usgCkG6QE/SDKcpcWAEPtgFSdsEqwUZOE
VdaCn30q0SwDCanbAG4QcUPeNrly4d2HwXrsYCLJo2/GEb9DOjbs/a4aFFXrBgA7
rB5q1veyTofxAymYj0HwjpsdRlSMvJjat48PGHVbkstRyg1vYjwMQtb6shTyvQpN
+UJ9KqPxozk7QACC4/93BPVkyV7204qJ1jhdSxULlnGI+5UWumGluEeFKXkidmgJ
lBcD1xZG87KmjfUq0pJoM90G+5R+/3yk6ojIie6f8V8MUmz4Y7DWezcRwav/NM8z
ZfclglA2CfcuOZb+39RzgptzcuNKUMhEEx8jP7FwOkcca5xWwFj2Mmf/cBpWZlcd
GBA0h6wQX09bfr/8vo7gLthkx8zleAJA1NYgtk2HdI2ae0fpLwh1csAb0gNkMP/v
CvM/EBtMmhyeKkJ3Jtav5IGCHaHpZcG4vLnKA+Kxwnj8E25Wjjm5PLImT9Y7U9wY
6KWPMAmgMqzxo0AQNSM3VT407meaJ23vGd6q7RElMf9z8nV+z9dL/uo+OhY0KFeN
dnoEzLeDq2RSc7nmA2W/GSuvA5m7UZdW36CsRuZdGhWsuecUFqpnJAcO7CsgyZLF
PiL6wti9SPTCwXREtIAOhgOfKtsxwTmG9bcAYZk5/7dq2ddpxaNmGqUmPJASj363
cJYUtF78kpP2iyYB+u+DJ5O0BaL2BbE9+ZkHhgRoKObEPGH4KGeuzLJP5NjkHrne
B0mPKOWP8TwT2zo43BeQN8ozqRdvX8UuzddG0WM4hNWeW/fCODnuARcDX6houpZI
14UPn25XItsa4bIHNRNnrXsdsEA5Bb84r4Zc0u1mKpU2z67pqx70PqRIza0djhr9
skAeJhnCIaqJuhah6eALqNIQqnaS1JfUULv5jF66U9DIwDhvWv+wAtxwd98djTq8
9GBV1XS1LUpR/HOZszlvhqasZxmipsURokF2eUJBBgzRxbwCLpIkxwwYttfTF2bT
IrQQ7zegd2DHTF7wRcbAOBtCzCADChU68XWo755qME/Nj48gN/Si2+gH0nmbtJbp
2KcrkgFcKa7OeuIpTVfjrWyu1mt8k/SvCyi6ECq+H+c0yyK/zsS8rkd/KsjnuzTP
zm6noz2V1A8pJbn3m4x8lqVi2Hujp+0tNz9Ctti0MdU56jukDhOuauzhQiN+lFpl
4OZNVH1FaOS2j2tye5k0d6JziSOc1KSMygAouHDCxXN/edi5TX4Rkz9njoN4TFQY
G9kGXpBXdCRYvLOpQEE9ffBc3zuqZU1jKKUZzlBWbn5KkFfOCEIPBKIMiOwLhXUO
9Qh55mHF0U0xcYH1ue9IvOTBfOkfNsPNVbFCf3QdTlvQjCVLcj2JohpbCQBZA+Fz
nq9VJDF73YqaK9K4oaarpIY68lob8c+lpoO/y+sfIQP8gGS3hV52qiQyljmtUuPw
bDr6LURTZVVPXcFlGjzljpIhcJ3LBo4bOUQ7mNu4+cvJUzjopm05wlLpRQ96NA5A
Amu1eWmetrMvtJw6B5KTxCP3CMqvOiPlKuBhq1YwTEFrKDAxEYxr86SU8RfUvPvs
71kLvzOn5fZhfP8azqCkQSwo2LIz1UX4WfIzI22G+FGOg9GSqUPyMSoZADvxuTWv
Nw22IF2FSw9c13T5MB3cknvsDUVkugq+uwKbBAPCcXH/ESTffJKqougQg3JhvmFu
vBOGdcKJP/l5gUwa5d2eKZ5Fh6J5H4qtF/7TJS4xm4QVD/ZS29OZUkWXbAdZ/RTN
9wPmjgJu4ovmIGbNOwKHdHzNSEziyvT/0vxUloc+jMGOu0AEuofxOECHH2ehH9YT
AcbLcf84NAt/xfjizPSWecL+RQiSgpiMJh3deJUIwO5FqWK3+uR8mesEZ9Xjp3M+
4BVvB+vkw7q2nOLMOSsjzFY1cZH7c10300wMZ7yXyZ7xmuiX9fgmBsUPb44mULmV
DvLSeAnOUgn04O0CR0zwS9D9Apg/WfL2lL8zMR3v1+FKKpoMNSn+LAHhfWX8Lt18
r0NmQo6pCmVvp+dmjHp/LSxEc4izzGE1at/TXo2dwzYZ6+3PAJlFdvXkKBnpE4Sp
efx+HEmdkF7FgjRBbbB+3SA8vrSlK2FG8rdxUWFZurzLPjpmqJFodCgJ5awAI2pc
VsY7oQ2ca71u9CKNldydK7xcC8FXcaPStd1S2FOiXVJiBUMHKc5/6evupS1W50El
qvfMREAx3T2sxvyIzFuBxShpznbsLKjXFrPUyXWkmfJEVZMyC6z2I4pmWQ/dec/s
EQFMvaZ5dqF0f1RPfqoNA0DLBlZvzzLNBP9Cm/B+pHHqmW/8psVRGJE8DVERh7Sd
HBUtokSnbOBGZhw2Hmx2lUtWuK06Y8kYbJ6TrGx8OyrzYRSXbIk53LzLjU8W8EJG
rEWhZdQbdl8htLS+ixyGuT6UGuX51Zb2frXp4PbwJJ0yER1falAxTB3vAolbq8PE
spqbf/7CcBPwiqhGCZsyvVpk3HXeBsBpwyzNniwo6KjrALDgoJg8VBxK0jm34y0F
cOovyuKc9p1DRNua+CfI1vZHE01afb018bSNsthydn37xbvvdPLHOYxz0e/BXXOw
a2Zf4/XwMYm09eCdDZ/pbIjyr2qLaovh4MR5LR9/3zMA72DhIRWsSO2MHhujYYhT
j+/yx2H31X0pv8Frg8Ii6htTtVUiEQeW+SH2+mxvABZrIkyv59RUCxi8JA0g8uRN
qzKPzngYxKkYf4PWga6dFVp0pIaJHR4pIAZV5h9pGKL5U8y54punLwGJ4U2Zh5da
YpU9Agxjb9JHkqtqGP2iIor8ESHItDqHHsHj5siiDqbpulOupEuq2BfeD7dG/tMu
Jjnwa4U6+LD1TY3lm2dBEyJLKP3vR3YLqkRrHs7tLAtPHryENSeA7FlQzsWUlZ5F
Q6+kxYWhR5wQRySfrGLtQlF6sqFbHIsO4HQSKq26oRF/CaUmLOKCic5vQ5s+m11I
ZuNfpB7g0W7BSeiiSjxUK8a1NfaPP8Im0g8f9xjpt2xq6Yf/PpZWWAzAHsst6ATM
f8dz52Ptdjb2Bz97G4r9zj27lHZwWZJOf9aXNxMftvX/cy6caEWw5jeNR50isZ6s
VqisDT0AVLYeP6ItcAErD/ZInsny3C1ox+ozRMFvErf8ks+jhXRn/zhwV9HuZZ/z
QJ0zDIhCQu80SyOn4uNH9AUAyfAXSf4RYtmjdhW1adT9xAd/r2HLw02xWsxaqiTJ
FoYylato3aMESyR/i3OKpHsqMf0utA182bRNuVEC+fRIt4nwfYRV71AueB2EAKls
FHfYp5o9SCkMtKdeNnyJeymTyJDtiqRF4wBmsdjW19UtwBf9Cbv8+nTBAfd/q56k
d+IyFisbQQLvwcdYVIkI+CpUjvqWN8GzDKIg4KSoLI5XOg8sHJqonoh+84PO6+mW
KHsXeEvCSKRQbQfhYFMkZtt72UMi/lmPL7Qtt0kQ259uUEOl6IRyib/LKx0jJ6X2
yzUTzRKcUY67aNE2dGR1zRXIu9PIAmGP6zJ+k1CfZdKIfHCJuAcVKndzeEANfCPn
alc49kA53cGaNUk4q0ccUOItCbsdMiY4ZmKYUkqrXgLhrcHENfo0c0vjJqwxHNwa
F7MClI47GFkG5w63ZYD06DV6TRoDJX7eRBm6Rcaz2bWMn3YElh8RjrhCyrog61pr
HiBoraMXWuItCc6bcTqmb89hM7fiqn8HDJzVzUq8pQFjUluZMTPu7CbwUiE7woBU
5x9K8sV4W7TTgHj5yfmDQexXFfb3y1OGJGd/5URVP8p1tuJxWuI2EN/ejDvTkFn6
L5HPtDofA+yIFhUhMbro1UBP5kTcGcg4xquR2IyNKLW134Z8ksvHJoMoGHEfV81q
WmsWZE0MYjj8kGP2quEQaYtz5gQZdgCTHDAlaBKGKXDpRUg8P4QIhjlJtGT1WrEb
BT1zp7n4uPA2b4EhI2jB9C9w7OdYDfYhnI8KcXEh+3RQKaIRc4Z6eaYmahGNulPs
x+t1HQ2JxN67/IgTOR9KGtkBY+YQjHz4P3EnUus7MtWEIoSDcEIA00mK5V6BcF2s
NFtO5X9gLZtvU5GAkeINC32bXKs84qMcleI3GUXgL5GfPrDE1jtHo1XpudAz4njv
cFkTSirxOBIF/KpMDSIfKD7WVR6smVcWoVKECtXUmR8ApOxJq728JCJ/fYDsbpmE
lHydYG+Oc+Vn7y1G7bQPiGRyz1mtV+9kBn1eQoQYrvUi0GwTHoXel8sdb+sZczI/
onHFLoLe+KuvWQDAKZmjtzuss7god7G3sW3OkqATmIn+AmoHMPr5vQi9bnAUxSjX
o13ty7Oo8mGYnlhvcvUsgdjonpuabq4lIN3Sz+pxUhJ2El1h+tW3GgkjZ+jgLxDI
da6dN1PU+YU1GZslxnMQj9XndDOcKl7/1irhVf/YSx/DvUn1gJe3NN2p5DXalWpO
+Nv27bi15y6bHgTd3eDTdeUvO7G9JU+Ys0f20qG2qLyJdgiyZJ0cLThPFClsO+0/
sVgBW95OrA/N5BJK4wwIH7wLqS4ZRF/secA+zrEdlGNj+D5OpblyWXjKob4vK71m
/tk/5KbO2lh65RiCQRJx3eJFNEATGLT4gj6pvb55xCRCrABpe4FuH4EAeKu5Uwas
5VnYm2ZYXd1BHBiWQHB4o0HByf4Va4HyqaVutnVpYqcnevX6hWh9uXY/rlLtMuIn
mzQ9OfXoJk1no9mTOyuezgbpsZIHD2bTF6zshrQmHkDCx6zA2U0W11u6/1rk+szI
avh22CgvOQa9jn5Yh1swfZLHQOgd5qn39SkTG4BukaGTWrotoJF1IcYxVYAA2oMt
Ro2IKC3ALXB5plG6D/wllC8iftg+rYIUZFqxkrAvRzfoKYh/DKj3yuqetXUJUEPt
XJT1q42xMiAsyN5NNCDohHPfDzBCZQcHrLiLlZZOGhJYrwHD5K+XssS0nSssX/mJ
85KkM+GEMAkF5BjXbQIz6eeWa0S2ZJVLBjPytkOzJBO4tDV9qm7SaspzR2fAv7dV
i/lfAR1DFzsDoIHQbWiI+KVDrTpe9ryPSKkOGq9pJZRBSDVK5OlZWKZzuV/Ysinm
E8jX8L30k0UQVYptvRueOPGz3VjtGkITcvfghFzqC6flrTbuAOYnUcfu2qsRrGD7
v3lVOOP+xyYH4m2BbjZgJwCLWCEQTTilw2TSM/aUhoFwt8ptZJpDG59ed858GDEe
0++wU/D6p0lf1yHl+FXGuw3ADe1DsNlfqa/23AveSN1bsmNqONDJ7wbK3NwIMsY/
+43OLAh4+3yv8TCFLDt+AfAs9Bl5ovhUL+4i8SJ9LJQORyv2n8he8YOgbNMWhOnC
zFTX9Ovf8uANoP49fYsS/2zo3Z+JyiMwFnZdFUtnTjw+T+2GZtHnm4gLFlc+H3xJ
HkqPnamHxPg0qCi/1adRmeOaFEbsHw+/MQ6uooTT12unALI/fbnXYPMxctBOkRZu
2kBfK/+oWFnPRwae+YgxNqzMineJPLZq1gyzjrlPvI7hJWdohfjyNdDKQ7lx65pK
EO+o3pvTwXf9MOvMSKoaLHSUUbjnD5VmN03C8G1VVdKS/QV1A4ghcUDPaeF1Joj6
V1m1n8A+YhFoBEpC2HNSrYR241Zc5rSVO5eqpb9d2FGykTubB/QCtoBFThjtdhmK
lL/ChbcvVOwubtIRMw5YuFNijmvTfu33UiNE4yqGfBPMh8uWeQ8jSSN3EXuDnAMH
1/ylHvR87DBKprzinCh4+qPlSPFdBpJpfuLVGj/Xfnak+6OCo4eIoePp0fGB0uX9
52sY55sxTO5oZnaUxQmG0j91Ckjvt0294O5uUS3x85v/8aiTI4ghhow9pJPhOY6C
HUNzWqpkDHXLSYkYvIwffiOlx2d8AfyC6ODYVI3R60Y/p/o7zhB/GwAYGcsx4Du1
YDGYu5pv519K7nlZvf/Qz4hBtJCGhUW7fr5LDpkfZOpGCBhjpyOMd0td4FV8Fbh0
blNCOJ0a0Jw+GJzaOHiRbgpV+AW+iQo0EGm3b2pAi/RtYQ0HpZ5Q8gvyeouAy1fL
6vgtOihbtO8+SurJIwP/kdRKk7RlFApklnaDKjmsHHgYGZYJl4DF2932aNjhXxHK
eifOdjESXtyfpD/GryxOTm59KEEQ8f6hbfYXLxm1HZkizZBh3pYUOnasrJywXN/v
Zkt31y4szY1UZEmS/FKhU2gzmTEipQKEmdXt29U5OG22LBx1oqNnP03i4wSIi9zU
/iNcPrklt930cYjDfkvN+rVTqYBV2n/FWstZnftdFt5oLKDHVZI/3EMpqBNf2b21
VgYfBpwv94EV3Dr7hy8nj3s3NUn4fAtZXW9Ac6/9FW/5yAB18aHhKRQ7fsxJFxWi
rgudAVsffHr4LkTP+ciyTpWYb4yPgNObNrasiN3+7slv+yfLChfyTQ7PqZXlKfIP
OOsGFODT6RISNORLMigN3KT3Av6WGsjGbh/c2P4IEyGHL+3/W6KElCAy9/+F5mVG
K6ZpZB7U/bn55eWmEyzUvXW5PvxjbUYanAU97FcvTp5oAEJkrvT5T4b1U9ABPb9Z
55ZaC9hzszjKgcZDAYv4Vz9wjIURgFocp0gYjTNM7Ktgicq/mAo1W3M1KXz+NhWg
9A687zZ+Arp4rX9HxFVbrI0DVxgb2PNF7XoBAPpqJ8JTrMdGiu7nyQsqGWP3+7SA
2j/UInY6kBKh27xeagfzkqu4hyBM4QbW+RIpJgHLDak6v6Irog11g2sYRBGh3n1v
1Wg60GjAR1cSJfzVPx7uxNlHBcV/CxfGOGX3M1mxg1AmTIZU7owdKeLkxqr9FfQw
WKKLuJgnEDqEuOTgvJyEJkorR60Qe+X8EqXC4HO+IebeGdm2AbeYZU7gnZLZUeh0
zpAstLqzwsm7bE+L5/fPx6py82cdDiZK8tk8hFa9SGzuiidZhn4jfUCb4tffRAUi
Et09MwRfHPQWj3ziUSJD1o/EHvXKlj2dOulXSZ1fTzYRoR0ghpiHXKRh7pQ8lGpB
+MYJHmtXZCBt8WbLyW7ZsZ4GkvbZdHRgge0pd+OTlRmbFDCDCVTZbdgl21sTs/HX
v6Kp15h3BZBfPcm1cRhg1sfQKxVnN76crVHIIgoyqLIOuElQ/acyxZIYdSfXW9Vu
/G/kUkjoNtKGUReVBWBpJ4pucAyl9figolM5qdjCc5gpdpYodkrPEQOeWWPpvbeE
rZx30Bpkd1zfJEu3y3MdjkUzNWRrWxe7Zq0KRrupi7B0gjuY1FAFa8HnMS6uAUvy
mOHT8Mt0rulpRy7RM2mCHzrNB8ChqyRXmDXpjow+p56O3GOhiRqXnVzxL/sMDQkb
qIxYrp2Mx1figyuASCAACdOJm1QyP6bhJRVsdmaTGak2Oqobb/q6y9n3s4LWaoYw
5GqvBaiPJds90cfE/lzSmItZiOck0GImB0CczvOFsW7XSaCB95IlOUIrSbfFEfc6
RVz+4c5UhZ0AdNWZLf7LkVfJsXq92aYTgvovyvoqSz8cu/FaL4AjPYP9BNWGVpp7
IEHvvZh3XXyRATlwR70vtCVupr0I9pjau5jA2LMIS9vs8jP9qBrTHdBQrg4KObLt
BsOO4y03ydeWuKPy8KeNJDA0a5MDHV4VCJanKagURfe9edzBPngsESNGniLVM8MZ
ADl3b7yDaVojF9raaUg24FYAt1hNO/Y/wVrCXHzc6Ewz61P2xatAAQbJxdZJYh6d
kgZ9X55grlg2CJa47M3nZluCRGoOKd9PqxqY2hbgGUwNM3EAlM7Ie79bPYZ14cZm
Jm+bTRJhyNyQ9cKBojnNG9LvJ5A6apdtOPT6dedGbzgp3eoG4IhjYZXzbMYj9KV2
T5X1OmaDpUVRLzzGe7P6HDp652VJlsMbfciphU9r6NKXxvSP1RCN2PesswkovTld
99O2dQeElBtAeDQTjm/prsgMD7cXm3fKepGRfdgvCWX7bjGZZ/U7Jnhpv6ur2pEf
dtBOCO2E83Or7YkZeSL8BqZ7zp8vpKBrnElJA35jJdJ7DrPi3UB7t15YCXzvbZaT
pYZ4dboRFGvifYIn+cDTdZwvWpJook+90QDJmuL6u1LLxK99CZwfZznnQweKsx89
djOh7uHxI7l44Fb+wU8pVI52vxoQwyG7StAX1HfDiqY4QkRIh0KmBS/ccC4JacOw
rmHmUB1PXEHiSb0KmxIzZ85AXWvI3jwNwyNsRUTJbqv6lh66GAhbWCKW0Yjy3OE9
c7suuARGuotZ1PHiMcqbzFH6WgIPN/JY9KaEQMZBi8wjYuRKKl70G+FFvWrwb44w
SkBYHkoDUPYz6EBcA7h8x+KxNQTNkFWJND4fYFG4CFlmwSvMEy71t0QnU0Z2KeOd
zMnj6YRLkZVmXSDa8tLVFRUATHs4OBlgbkAT2TtacnARk74/v2YIgVAEtfWgXfXu
08VGkGkXAEfIYCbVhMu3d27rDtqo6Ms3NLPEFisOMcdWnkO5kOdA/Yf7eL5DrcAh
6yxjpFpBA34cft0g7yEzkLPog2OZKUdUG/r6mVURa7ZMFW9l+FxVgVxnAo1DdVhg
5lWpi+5Qi8Q4x1TQDJ0r9yCLuPTJ90hpBuV7reuQH5jSNb0FeteQ2Y4HqdMJ6qCX
XfohvVwESd9FHVXkR6iFHcfHeef5hQ2u9Lu8bKXoIS9I2cC7v/oTt9jdYjFxwYl2
WNtSKUzBOjIxrS6Xr0C5hKDedPBWLpLd1MUsiMDRntxtrRY3Dt7vo9I+EUooszHy
jxmJcU4kmXskhKst5zbcYZQGwdZjm4ivZukECOi9Nv9HPuEWWp8QctI8M6SY2ka3
XtaRvfV07BSs5CDgNa3d6OE1M4L3n7Q4VDuyIPNbfhBeEn/0Tf4aJn7gYiXxmMUu
OHmhrd+TXol0P62QynVrKme41w/156GTaVxTA/XIEmksz7FFtPqiUMu60ImtEvff
VuI/vs1TmbhzvsFmgrcWp67jcCqqyPaRTj6yb88Ba5dLXGjgKV3w/fO+Nt+Z1Kid
3RDDEGxQertMQ+6LuwW8k5f51sJo7TYmaY8X9O0q6UAEWwYAF0cVKODVqrLNCqty
t4SXqva0T6cG3BwrPxD74sl9IZTg/cFJIQre6C0sDV/G5pEPL/R9+AvDwY5IQqJf
DlqofWxqGWag45YGMzgqmhz/2YVNPWMVjYWERkeYksfUCo7LvKYj3KsQdkKmZsjH
uetn36dKAVuLIZ7kawNuVxWpcqfTepCYU7jlg6E1qQheIua8rxqub7DbmkAr8BIB
nQ+hfR8GV4BfR7EmUyER8C20wFwCes1SSMFi/NDkUHV5PLKCJOKbtsGYZC/UDm87
7iu9Z5E9hJ59ngMailKppraDUVqDGG0onmc3t/c6uD2r/YjFLvWCaLykz5dUmE/l
K9vNbnSXKT2iWx1Bamet0jvgJ5YouOqlFlmiwOQIMbmCMQ60mRIyABSkqGUcnFZ+
/i6MQG8diEsfnfLlLU9JYgkjFyzuEjw7pRoDoJ+U6M+gj8cNA4pBsgk55wxAa44L
YG6Jo3ug2+XUBzwztSAHtvvV4iu1tdD49DQQNEhf1KtOL3o1L3shE3wmfFgzsX2y
S07LNo1hrenWtQXWpoeqncBWkrhctTqFywm6hFh0DLvp72WUF/MMYqryRn3aIM+1
FZBxMqtnGZtm1Te4a/EVIrj3OKaK+C2FQwsY6YdPX6gZwJ1LQbt2g2ZWFqwtf5tF
XEvhdCJqxWa+L0nEj1xtp0f+MCvcTVJ1lrLFs2+TV1IfNivF1mvzS4i9Eel+UGIF
gdaSQ6cHjlWioQX/8FWtd9hbySB0/tXVZ8rTCt+1ZmoZkm0JBwlrQE2wptBiA3Hf
IJgS8VLU63GVQGZ7uyD+KkJOLHpe/ZK645yQWtcZpYIs/2GXWJdqWWNHKvtQfJJ9
dgBTg9K4bh32/P7zT2BQIgPNuKDjEN1RpzwkukButsACnbDgckCELRQ+2IqU3is1
osd7qvYkJWeg9hIDEZAkZ7NJGLyrIxS8XO1llo6WyMXIJ/0UfzIs7hKpWShPZkCS
ggNBZXmrkmg0pJcbslT+qHfA34AoR0ynv+Gfa/hmu30bd+Rd+0hapTpvlHoCywno
VAqrziVQgQ6sHyFCry5UbxirSetnsBHK+/0PMRi5zH0Il0seWEr30XWYBs5fbF+y
3cqP81uq/EmOPrOOV3v7Ttn5NcCxRz3ER4RdeoKvKcmIAYq5urEcVy4MkMWrawrf
De//thIkwU5z9nGhQgVBYHbM1mehmMkG6UAjfbU46w5PSC9/WbadfLD7hzk6jLZv
jjja04SQjmliK/jZhsoWme6Q/yYd5MLLimmGWGU/qY47rbmVAGpstGrUwdvpwnFo
GZSfBobmR+xEstI9JahwyjZwDC/2dhRGqSK0UT1fE2zxOrGpGIuGqos42ljB51eT
a5pVPgtt/RnDOvNTwUC6EqcRwVpA+QmufJqOHw7P84Ys7eoG+KK8tymh1zCrMrGJ
xpYZ2cw0NmQkE/iMPFInSMJZBdctQ7hggef0jytA/ADNIvir/BZt7RgwybeIzA7/
bcszlmAKLW7zAWVrbLFjfXwXMd4aU9hsKObynJxW3reSReFFpFKxSr/pMnS2qO4t
alpGrBi/Rn0G85e61cy8Pu/UCwlvvWbhTF+I9ZMIb3aZmQHmPF2hF9GUyH9Ntkta
C05BrdKFMRuZ0qEQbE1chOaMppIET3gNo0eOLqXm3amma91IeB2Hr6NHMg5Zhuk9
6Aqu9igdMYlw5pAyYt3BrDd1tq+rC770S1UZKBm2+9J93f/b1DqhycjggNW8X7bj
u//2M/YHGsule1/h0t9Qh1VC3YgsU5S/GX5jcO0f2+t0AZxo20mluAd/z1Ai6GMt
4oahISM9vTNOwdUhZvDkcV2IDtw9v/PMQ3ioQJyxgP+hxYe0gAT8mbHbMErrfcSF
ZDce3DcmQA+xLTdQ7WuIT3xzVdZ97dZVOEJG0KZ+HnpT8kVZnDq30BOFDbVk2EX7
jcu6VItsEyZWpTZLHesJdCzebQQIUuheB8FJdyC14QNQmdt947hNoBFVnj8ktNYB
OZRWAoKtaUHZv0hO6qX5JWTcNntzKHszEnD6z2ejDPWoExPW5zzBeTKmTcOux1Nv
NrYOXzmro9hJLFWOrqSvW4kn9bfOpPx9m+Yyr1ou2FJUXTtsMowjI2Yd5vRWZ0gi
U7tu2DtGpvlkHjqWjVO+v6Gu3m68btjjMJogeuWBAGAqq2Hqf8hYz3UbVV1AWh4y
T/zCJUn19eP88Z9fT4Nu74MA4QwFQduhqbLirQJ0gLpVi4slV6PcgbE/z0jwFTEk
fd2uy0ycSdzKc1p/jMq3ZXpUZDZohC0vco1bw2CmF4HpbAPi6W8hPfCQ6jk3hN3S
aoFPAYmRzcchLpjNBV8osqyJe5GvOrBt+tMTCV62gPy/71MAUX5SYi5AyoPkQUlD
/QrGbr0wyNuAA+7yDFbBA+103T3cysNsxunvtPit9M64ufXT/Pd5kxRMyU4DZRYF
VgAEAzpnwPklDBFhroeCqr2w1PpeufxYqggb5jsq6z7gZN01xw1+qpXRmZkRhRSa
wMmASRO4wP8MoVjG1mxp/LvmgdiObAbB281KlYzo2ISPlEVw0F2rWu2n3PUCUQ9E
MCYWHUPe34Ayx/uAcYCDwQ0MouBxRFriclu0/rxO49te5WuqFLQ80c/W2kZH5KOS
akPPyudIupZloE4Q2zddq8eLpJN9BRQH7QfffzA6WpGuUZDKavlQMTt1UEYTmVXF
96LohRttk8Q7+Oc09QuqsnLlLCMMl1A8APUijuPUpRWX9+sh3TMN48jC8X9ooEXk
Etp6YRkO515HboNI/mST8zQFZiiFrUo/M8Eza+Y2Vzl3Z/PBon91esP/zAY4GVpA
8MDoxZ0lfLI7XV/ffdHFw7Gec4MXdbadGRrkp6cE0SAhc2x1Je9ZjPGjdzpaocLO
nU2m8Q+TDPjoSp27Gncz8JMSoC9LEu4yzacNGlIcuAoV6egfcEW7cUgediz5IjN7
ataVZa4DB+bpW1UY0f44vy/+clTzjgQat2BXoOqaxDjahQFz68h4khMdd1/MhWI5
7bD/qcXmuJB1miKl2l6fvu28KhfbZy6xLFBlDPpAYIcrM1XQ5qTMUTHzLE9YYAzh
etbUJBefpu7GhAfq4nFONDNm8hYq4dNJjekW7Udct/cBf9nKQQR7U/Dr1mSlEkgb
EJzKFJMb0LLCZ9pokBIHenXCodOve+y3Ds84RR2DKRjEGAr7Tdc+YD4JwbINU42I
Ks2t59B6VXhQqh1WD84RKpRV0KaKDVjj8L0gT/o47lX8b0uKJ5VT1ZHwByNTzDlo
Ma0/ouwWBlHhouqXqQsgjUsAmqZVb7EsJ1vtoNL6iectlo1NtKZMdVhb6+RIL9Qd
jyb4Znf78XxurJ+CHebOzYI92oKRbDba1EXEKs6dGe0Rn9ywZKnweMWYVoScVbZ8
tdguE+VCKRTTReJhtvCJxt7/R52xhKi+/Lr+HygjNNAre31TEL2K6zqgw6R0wgi1
ynGnGbYaAMGQaAvLzKfW1zQmfvytv8P6mNNEa8h23g4B9cyVMDazaCqETTitDkus
l9OsaBmXNHycUhuULiBHrgi2SgZ0DnCIEeh/2w+W2TxYiWz0RaI0RIG0pZvH1u8h
a3Lj9meZLjIKna3N4GjX5g1Mt8IlqRNKrAJ4mXY6YsYq6IUZofpbkmZTnZziwBbj
7kFErRbJffRq1m3xGXEaWW5zm5hff10F9dLHlfbZmpq9E91N58b7l1ZQdqSjcRi8
D+8oMdlHKAe/zfYWtsq0rvkDvNuv8KDysdY4SwCrwAgLsinr6rAA/V6E+EWrWlAT
37/GBKGJLkHnbGEOrd0DPbAsZ0r3qqT0eym2tWfO/zulpAMgxqeT9VYxQsIvX2ji
PDR2jPZugtjSLOXnpyGFKJbhZgjzNvvktzIDv4/G1iIWf6C/QDhjQPpCxuX8Wxbo
iwcVd76vO5M/9ogALFzec4OaH4007xdO5IOgeZfu5K3rvmOT3aomA4bnye0NPYHn
C38sEIXZzlm4ELQG0RTP9XTl0ffExQwaXkLTSZHHvSDnAXt+SdVhrsiK92eJn9y1
cQUcfszBxL4GbDheF4mIvCDYwxW387gvWOqObOkL5wFAIdgsZSm3fKUQffPEAV/y
1+ke00va6EHTPjmweKToSVv64YCk61VDTB191utr6tRSTIF0eMtGb19I38CoFz9L
X27M8J49aGgPyq529FP2fte93Lw8Z80qJtwLNnQGsURKYo3l+iZZiW37yK/Z3IgR
WvdROFR8T89n3r2zIihTS6ng9eTmuzLAspU6BmOSBJQ06Sj8BNMisuwUk6NbRNQm
w9yseTa5c74Y8jIS8uwxaJ02H/pB4p3Hl+jLslMBz7633J5G5f8u3DBUIoUuxMQb
vcYJXH51pr301zWDZv5cVrS2cgFa4GVuJYL8FwCbHgNGO0+6pmjFBlmQGwwL3lJC
gu8IuhxsvsKrxbOuRGURQaJXx/opFII8mYXUCbvZHWkynmjAPdHMB35zfNYYCVXJ
4o2xz6p61Ie1tcif4zOzmicfGTLetKmYEAFTM1XCQhTewvOK4FONqRDeScqU83W/
Apn04TBg7h+DRucCpwLnxccJv/Pcah9hPbp/IQ6D8Vcj3ZClWel5CxXgKDbvQeOH
6oCqwI68hyfT2SQ53Ve41Bd+rkJ8DhEAqkIfbHgj0UK5WRg86tUQ6YEnmPudWkId
JhENCoaBC/WuT0QAj2IgyiTqnse5diROd4Oqh05mP9Gp1WW1sEtb1u4/pXDBWUdN
2xDIZiScEdWDaHn5LFTxmbxFWOHUwbe61DHZzNvbMJ3zdR2r93sN9Hu74b4Nr81T
gvWvGup18ejDrImbpDZrjDrlHLfnsMKODztYmwyG/VxmrGXx6tYQp7XNPJLWhqvu
/qqpeCsO+SMdG8m8oewGQSffMSiO8lafZ/ONm668ZVxbYvsXrM7ERR8Fh7+hV2uu
bN0qnPcXnnyAGIFZmFedv9vm01O6842lO8NS4HQO4bc8HcxXleWeu5rMTLOtxZw5
KEbLG2V9DpuUmqzzGUEJd1i2MLXPk+kY3Lrsb4k0CvBx3ED6oCH9U95iMsBZGGtn
6NcvZZQW9HgH0mCTOm9+tHDVvNZEWk6P+DWXtD8/hAufggdJqdBGtWwL9YBkXU2x
6+TPXquTlW8lPyP1GWapXOdJTQaI52yJArG2q4tAgI/d8TuiRa4QMLrMz3uMwkir
3De/sEhCQ6/x62MkZnB5tAP8CBJyHJJDSszsUfgRa7NrIFs2hV9CanGAGv0YY5+Y
icRHbhb/YpanWf2U2vLMwO/li5Oi4p+udB0siAup2FXghooQG9QxwT8rh3epyZpo
E3jS9+oYFuKbB6LTqZkwjXND1cciueer24C15mDWMBRepmLNzZaeGZw+Ex1e1mFn
cou8XTh+grQ7b5aXdWSphV/j6UtlKhqzqknm1gzu3cxcGbLC2mlVAL25VL24UInD
KvKVblApbVYwkbLuH2uBccldC1yH3Daj8l+m3gq7GcAvQxmq0/CixkPmsJhz9MY9
1pVCZAaYd8qDrNinoThyuvlfYQ3ECK4xD6Ir541N3o//RGzrOExl3ZvnFPQN135a
b39nT9OL5F2HZOIt7Vka7EvLZw+jlCjYfLueqfw2IFSnJ2fHSFabp9Vpgci9ewUF
73u0UOreDXSPGdlx4b/sP1+uR2MTPvo/OrfS5zMxQfXIi8eV6TVPXatrinhxWemK
Ihq55RjiG94hjKaSGFYjBXNp2JTNTrNno08P6ZS6cGLY8a7GmZQO4yd9qkPTrm1v
RbOuhU77tr25ym6MTRcoodDKyp8qMXtSRWl+cIXmAXQYbvICdSHYE9hXgyhY696r
ldHsswQpK1Rz6ee4A7Y/dzjIYai4SpnGZDJSmkSQavzlZRpu+9ScRmbM8fKc1O7W
QrH+jEAm9QAC2yY4BWXW9S6ANz3JvWR9QWg+miI102uX3fHJHHBVtVlzbuH1opV5
R3oPR7iMdCycofl1C0d7kvQT60/EPOyOgEYBIOycyMC+8OV8MA7Qd0H2382F39EF
y2m8ZoUzh4Tb2miKxquRzkqkPKeH+c8fQl1rTGPeByA5iPBvNiTnQkAbqXZADo5P
abxHfoUJkyBmOy7m2OV65wG+l6puSyMVT8LhjdRhxA6+WW8xWZrNV8iurhfmhbSh
HPsVmWFZNNNmWkCFZwHzX/u46aYCnIHRI6X71Rr5UVyLxZhmV1mIlD1mZfW7/yBS
YEozHNHp8Qvzllv6KsMrL7+Yrqaj8oC0Ym/D3aSEl2dygZTW4wzsM25fjG9VBM4q
eb3/R+igdxV4KD1/petL//KfbOhWc48qI4DjEZkIueZLkBG7br926zm/H0CxIVjU
ke6gRzfictu9QNsnhEEypjTda9qkOFnv0Ka6BSt7d/f6C8bMkZyWDiQo0OXag454
9Lp6KJSJV6FXvYQwclo0zn1R+UpykPOYE4h6s1avBjnL+QZV3Xqjou4c6ViWNQff
9zpL9GxPgLH2uYkXk0ee/W82/fvA9bJzxuZi9KEKc55AciJqiLf8anIU7//2yniq
54v5D5gTWtPwyADcx95U5z2lC9Mxrw6i2CmAp0tJqgtHr30aLGTm0GLsF5xGxzHw
p9MXCAvU1iGLWEL+lVvGJGnL72VayHfzdE+lRq1r19wxhfmDs5Bcb9rXOWcuVcSD
LLFW1Hv+kBgCjv+zJyEam3Lc4rzn8wYI69khUehjy1C8AubHGruGjDeyLuNxbfyl
gUBee0fKuviTaa17QKJy2ztZkbUXamo3MEMNOX5Y3JKrPyQ4cCqJsBybsSL/uzrA
+anj4fekD6W3XrLxU26+QUCyKYiIZkLu0K7v5DaZKFyK1ikqWGd2JfmeuGxHz3ai
b9ZW2W9i+hX/l8TDSYp0kpmm+0Vn4bFmUzYABDHxWela5vBspEVU60yMBmReTYVt
7mXPqpXZj0ID8NwrjrJJxxxkGdqRwvKFo+k2gCmAkz+9U58vM3zcWF7P+BupRtMz
EQojbtQt6JXEmeS+k7bgb6qk533cLLFgoMfOCoknJMDGEL9xWRHpMlhVxIGYK3hP
sJD+IP1YuyvSLKsasVyXL5QHukA5B7/Kq+9oSdOpBbCPXuw8MKqRMeJ5WSJdKU4S
CaVMOm43A+OSDwUb0ZXu3ouRxCpQ3ob1ULiCfPwiq1gp9Vp+xD/4ZJY3BHA14jt1
cf4HaYSYJcJ7U5HZNMIDgbritsE8oGUZcyyazO34D0K72TBtYu8SWWg3mtiZUHO8
vzhGXPbGP3TiIonWRPqaRi+RLQS4aATJV1ejxceI6v6ECva5/KmuokRWjvf4uyTX
iSSx6om+k1hSqwfSD/jo2mXRKf8KxN/oNOvMSw9zMF/ocbNAVm9zJW4Nh4iBY2aP
TnAwtqGYi87Uzgh9klUER2rT0CVJgGg/S6jVI/Nrg1jknqpVyr1QfWuVkKArZTB1
tgBCdhPbiFx+0M+7zpDumPoXXE0ZQXmdV8xMYHXTIgvCAF5SWnodXwRQAMLR2KAL
P+GHnMlNt3IjnRjQJanKzZslrAlrd5BVvfPhbfaok+eHyQbIkUfKNY28wInJKNmH
GsHc8/32TYjaJPI9y0nH9aNDVtvYFS5P8KIr8B+md9W/wqlCmJfZvIvOeaINb53T
QxmFt6mAU2NzbIGz1U2SIIu9dissD7df4p/evw/tEZtzDRf6QnLbbOkpO30wPBUc
yNqAmPXBa4ErlfuyqLwiyl9UcvZZaJjvqDyoQtU2VFbZ7K6sDzhHDiTUfvPM6XDO
7Uj55bxXnVatsTo9bkYhOZ+Qua48L/Ma2/HHgZcyooC1lUEpac0+ke+HzER9JUHD
qAo0QGSLQCSpDHMp488MhB/jrr1N8VeutLxgs+QMgsyfL/aefsKd1qUj0foWvevZ
TTfJsf6kAapYErk8iax2Eb/O8HORMhfg9+iXnwInqCkorf0Bsk7dBQwhSyhrCzc7
Px73Wm3F1bJMLMeiPVIf2CdnS/v8egVSTRA/Yu8V90FnsUhuiGKDvsQn6ljWOerH
rW4lw+aEvrAETVHvWioh11n4xIsHaWDVMYOjJNymnFKg2jpWdCNW90+Q4lpYRM2p
U6QCNxQ5MaM13FUc9tiEwqt0N+8OIveZ5j+w2+lYBO2N9d+i7l3LtG+zGutvJmqb
UOYmwyGf/97wMMV9D9EcMl1j2eoHBV7fK/Vwchr9j6ekVsybFYAxztR4it2HEHDj
lngrqS5LV5603RD+cCxcaADylaCgvF9vZl45iSTeU3lM+A1MMu3WAJrp2NW/hBi2
b7nv4lhC7/rN/hyezLWXP9zpVUxiQ1kh1ymajrX49EEl4i/nwltm1/jKMkyBclud
W5d4/LZxKG/PvEydxiarZ2A/n7hfvZ4FRu2pZEv99PRruHYxjO4iJ2cFATNY7nEx
8bMcE3mvFYoYixWadcNKFlYpyUczn+RAOdKGBsgMWtnAsPSaBedbHhFmni4nSUmt
wXFt/dRUqWWl0YYnjAqw8dvXTQX7eSK0ielDlff7TYjbrs/SQyLqhED5K7qIFq8c
bobi3Qpyn7dCgqcRWfg5o8zomuL7EyUWByCjzul39yWZpg37viq6s38V4AVbdX1w
Ls4Qs1Mya9soZvvfe4hNiUrG2Etwj0YJikTvmFMD96FMZtE2egsYkB9DNbx1cBAm
IHuLXPzFjwL3DH7ks3girSHcnVMeAq8PVSAlyrcbJiaziNg4+afxmFpG/c1zqFjE
pg+hCg1ZTFx0nn6MRNUrREOBWtyGULzijl6pmAIYLP9HSbNAEzIvd7pgYMjW9obk
0DslTLrBg1+pZ7tQRW7KoK3CUNUGD0rQd5IVH8ditjuuxiIWHKpf0B+GHO4LdZDs
gPC5pw0Rq0sabZI9A3A3DzdHRd0sdyl5d7qjUxDjGMi4EzhpGaSfAH1mDT6XDhR3
yBNmyaLRfUioz3lmDl2ja+61mevplEH1HOSiwkKq+JBCMWhb/2hC+NjoTAfFDnH5
dWlr2R7qGSc83bGOVbVVdNo8kEnpGR6EqOGysa+4uNm8XBOveV6xtNZh0X9ermH+
zb5esxMLX+KCxJiHqgNs30WYFV7a8AioAvLr8PQMI9VFJc9o3LCvPMvdVdwiqIQQ
PdE94BVR+AHdnuYSsl7fCJg//uBXT70/D5CKQBmR1T14eqFT+EiePVNaPS2k9Wak
PUPXqlFIJV8uyb9bGfXc53T2++5FqHHImBRF0tOIDrerPmEdBptj2TMb4oSpXpuV
M+W+c5C30R78IoN2OG/lBy4A67Yl77HmEsiz6kvIQOSl2O+hOyRITc0LuWq/XaZk
RcFafEY8WuIt0tE2PDtLLImF8QIX0VhHkocpciqbGblCCcrVWjcYovQggTrokDQN
WH51FKzL1t/2tfBIFgXt6hYEOGlngfn2s/9oDlAyuR8Gn/FbyeDR7uthb2KQ9Qx1
ViWZ0GWaNT112/8KARxW/VPIrFOOJmuWR1amTIMXuWccZPEjoUjwaoF8truPNWRT
8Z1+V7yvz/pCjnyZfXoBV04qwdn8QZbd4HkozCfwXmmx5nZi8jaBr76Ayxrx0dTf
m3uREY/m/m+aWS6g16aySh1HXm1xovOjg6EmBrQDDUAKv4OTXI0Mq09+DMXh0KKk
nUZvwRGh3lNy6m0wfQLiihjdtbqc3qIyaOnw1DIqcWMzoG2XeK+45/QB+R60wf6T
hzVOUTMoPpVCaX4t+HpWkIUAAan56brtXoJTQMbneLrnHPr3kAb1rrkQJg/X8r2K
oR2rPp/y00HvgRNDLbFmkIeSk335A6T33WvyVxkDiKyV5yMTK6gYOcvYNDVfdh3Q
rubcFMA3ygJVMbt/jZmHyj1p+ZSJ/P+D0Vc3JN5oUKX21Y2ba3bGfadOAI68jxmF
Xww2B41ggrtUdIK++26cRPYqu7Sy8giboJUUdygJOnCsfSua4DYuF1gfMJmjqVv0
vIiPNSPf0bUTLi5dN9CUe75wnUSIYeby3CUjODYLQPN/pweMTc55z1wyPCQBszzf
PLgvX+3bFydfMxWyHRqynLgsXGY/Qs/NWnfMZKw+0VT05wnfYf7VbCbUT+ts43N7
HldbmZjihB3vHNLermPz5IoGn2utA2+0WsQCqF4NZML+up9L1ILuyTuTZNT4qAVx
velCMy8i8kHSj8SDep8D8f1Ia/QTSPlhMZq1+S+oRjyUM6TRSh0gimyUCr3NwLfe
k/9AfnS9yaGY0nkOFv49YM8bij7D9UvpBjk0t8cFmXBtNd4w7BVmKpyGNie+xcQG
1D3YYPRhDWyvayWGYSrQr0ow9JoTF05s7smuAQf9cuMn6gcUsIW4399bxX6WT/Dh
wDx1hNXUy+RzG1wqCdcFV06oGl3WH2RMDz92CRJYHDEgAigjYwDjRCDAeJka6EmB
ADtIhAc+CK6kuVpbWP1nmtb7wZY6JVdsK7LbhYL801lkI5tFpdNitKKmhizDuy3k
apo84rNYEkH1jbrineC8vE76QN2nWkLcRlmOP2aqxy5y+WgMnNJ2A+gFe/y6krii
iDqrSuDAZRUsHx/qyBDUK19PBMIUTkzqA1csGOfshrXEVZ9mOZWIVEvgCHKuG1Oo
4SmNmsPup27QeG6ebv1MjCsBmV6TUtv/GGcxq6TRix2SUjMX68HYrCTw+Qx8donA
g4VYhrfjafRon5Xf8NwPKTnV+c/MpRb1dvAb9ObGv55wWemhalrp60VrBIQUPwhU
WjHCKcbbIZYu6JrEoLvBQ0w35YR0a7Ok2D/1/xyY7oP4mc0z8vBauBVm2NmXr86f
bVvj3JLq2odsr4lKgZVOLt1cYV4oPGIKxq7bYJmCCioOjDmu5AuK63kN/qXHPi2j
DR+kTaRwvdMfY292imVW9/ApRB7W6FwkH5QGmzotGZqQSE9bBW/XDW8Gy8Y1ctnP
F0WVbtJAQSzOSAyGWVlj8sxW4msS2wj3aek8Iy3Tv4YwqgvtkOGY3kDilT4qDGA4
l+h8RG6Nt3XH92XtALun4zbIWF4EOVQQ5ZhNKB1quSQRy2ou55Os3Fwy20yNr1fL
Fb04vx4iHssiqFu2NsnGtLf1Mgp5i/ZBlOfVupWPuBnoPBtqrkS55q4CSUd1jnNT
Qyo8dZwXlFeb3GjRQXs+k3guJ1YResxeYDmszCiBahUck3MS7ck2S/qbndqT/GIG
348fF58h/KJGRvqChBKsL5FRDey8skaBrhPxJy4C8TPOh6yPO9u11yfLHlMO6H4w
AaEJGb5BYpQbk6+lr7ORCGrVQNAhwCk8K6lcZr7I6A4yJtAbWgjuLacropa3u5kG
YBK8DxzXECamEQEp+XLV0fHWMl76vexsuphH3FL2Df2t/DF2ncqadSBlD5PetLXB
6u2c9WK9LMere1AqA6aRxKyWBFHdE1HSGGYE9dVYn66DRjwXTEFVb8kUjGT66Gfg
d0EgJlwtntLHK9MI9dAlBfm0gLZtksewyueKZ5UDmonQ1efugD7q6NYdPoSOssTJ
/6CS3ArI7hXHluwS0ev7QTfX5Fi4NtCUr6sWeoZLYaBf1IA+X6zLzORgh5HZPlet
Ss+F97ZPDDDSoqiHP7JkcXbg2SZbvwP4fpxmb75hw4NAG4/0Nn5JxUTdYmm+dK1o
t+niXq35S/UeAmZlRChBZac05uVVNYXAs9BfR1SUxu+0NnFD+nLx4i+/xcmrXoMl
jVWEcunZU80QyRbjAzQySkoZkMcowWla1n70VsB433pLvNSbXd6di8Irs1XHWbSq
ZfsMTo3ordKEQFQGjG30aOU44QRoGWilYU4HG6kEBDWIOf8LPxNi8TRO9FixBHob
Cd6Kz9jHvSOEJkkMJiIdPL5PHvz5s97ueEvu3Av2U5KrClHyP2y5VYleCpwQztm5
W4QBPi/dMs0laDYzU1IYCrrWBTPweM6vcfhIExN0I0X+/nie7H9ZwJl2hsYOQWfO
3ItjPNsCv/g/lE1180ZkQYj3Qle2IHKTAND8oLkLCNMC1loO18Tuf61UXe7LxCmA
92/PSl9ln1ocHEk0ucl2yMy3jOu4lI44CxqBTwZW/vDRwrhnjTQGYHii+otIZRcj
03WNTql3i7G3L/3dyykFHCeoEjkLucz5VAGgi7t3XpAvpxvYkVmGHTGT366vDNG6
nFfGisrnFz7oQcNBLae5+X9IiFR2vEnwDowIt20PetuEe74Doc1Oaw3ACotd/8uT
Mfp0THVWKTbhlqXufuiT6kPDM7Ezv8wV/2Y7OhbBBA6QS1Lscsm1q7IUM0Ab60yY
C2VOSbgaFNUTlTWQZEMOzemjQVEIdi9wz1hy16VVgj3ufic39AtkQRQSZgldrsKa
YpxWMPk1mTht/YCFN2Yg7xzMxniVFoIlm0Ps09edI4L7maetc1Nu6uK4HSqSB2Hk
M7Eqb4/7KnghvDUC69QxXRPVYzf02r4dmlInqJdvJi801KJbkNtxibXWdY4ByzPt
UX1feVFuh0sM6/334W0Mm25vKCg+oW9p/HDtZLv+RgAXXhFTmOEaaUsEOjJlf4V2
QevtCbM/Hi5+2SWiCf6/HN9TyvvxQigd1QoLgqNvbEH5ThjDekDnWhXbFYz0T/x7
g3kx1L34BSTNPVrGKG0LIi2570KxRDO29/jjiay37uYL0AY+EJdT6pxqQXwYVMTO
2CO2l+i7W3yNHlUWdj8BLsgjVEJV9rHGc/HQDuMTKItOhUvzG8rP/P1LUXZ3OPHw
b/oeq+mOd4y8bqVb2iPTp42tTeVPaIb0BGEupLU7i+QuIj0Kbbk1jLkShZfrrMJv
vYbZY9s54yH+1COX+wbr/1e80VgFmOL01q09bxRlv/207OW/0gyWDanF5HnrEOpU
oxs9cWieHT8II+evi7uFlYULsGT40QchK5JPieARp2siCGfxxyRE1MSk6ikugEFa
nGvSfGEhJIrI8AvvUTTqruGcVe8gS37VeMO9BI9QSAh5Moc7o2PVt6GwAGfUyCPT
9LRvrEPxcpV7V+eTgms1EMO3ZAKmt1H9QKKD6Sh+04uS4zG7SJF/ozQDrrzBAuWT
egHyhNUsd3fOtPD1MVeHoayZzYxVOVswoUZyDwFrXwOEZKMF4mlKRyz4fjgscokH
L23KQTIy5bndJ4ddYIU9+FVxTodDG9zDnrcM4Ooo5i2Gxymp6oKoaPBcAHYWD41E
8hy4NL3FS9+VI37ROUDgNwoPdXhScI+B0ExGtFXVgPbE14BXrJVF60mrKiF6RAhQ
bhb/hzU8o3/i1P7dhveHfW1aSeK4YBh71mAkhm7E6tON4Q+GOA2WmvJojGEzprqL
dvjuREbs9gL6mjfmE9IDf+6aEz/oNmCPNPYnptQhK3JncopKAu/kpy8EkjsWeWde
ZH3wkx3PhNUvHPDB2fqmm5INztRheM+uG7W8C/qElEiyNT3hc3eQSySNbUSZ7zmF
8PyKrPLrF6ZTKKMs2QnmKT0eZAU7gcbqOySw4aiDdYznadCd4AkU+a8DADWp5tKQ
Cz4m50waeFaXcAP3Gjlq4Pu18sT+nZaE70BsMxeC2nuyImql8xivXHjAx4kDe3OD
kZPr8EL7W0JsptyJvOEG9qsXaqhq5/9WJJNLge0rXjfmZrXShkAcv70z9ODUurwk
Kwfzqas2e5B9CKh5VTA62yKs46Q3Gx84PZcWADc67iPshMpxqIpXa21X8/xlh52S
rzblrJ3Pv8x14nHaF2TPeQJzo1KwRWJsS9STazZ5e0/xSuwMp0raBMks0NaKPoWh
QGDyKKJArBVDpyCnmIfypW9cpEdoXtIe2bq1kvze/tH1FWiA5sobQxAGYF6l8Mc6
DGnjZFxSt7xbMN3L5t/RitXC/SHh0/MG/85tahZZv5mNqntrWpr+y1TYfleUYISn
YcRVDcas88YJqhtpP1rIEOr/WEI2M4zds26VRkGaVAsgkZgVOmNtjJHG93hWpm3p
1B5OLSBnvXlG96OVH7okDsfRKKUhK45TQd+HEu9VywCu/6txE94GW0SFZeDmILMF
Y0f6EU48AF7diLccLDaJTQvIBmsMTjt2n/0NKDRFy0X6Zm0/a4Rfd7OfB8tioHCL
b1rQuxuxiWqxfNTtZv7wnQINc9OQNBv1gU6OTbrA/7qaiIlkRC09fj4Mm8L1NcPv
mt/Klqqovgl7ZUrQeWs7lN8bbwGQ3fiYOJHwmZX7qij8J+joMlb97Meyhvj6ASWM
jLZUhzItaydxozoYU3fF/mwudyXAA6wGsE2beoY5CBCReCLIJjerrkrFAAgNK7Oh
pTfw7RCcFE0R3EV1xI+XeJHAFIRkOM2hFcY0Y/wqatq/N0FArzRkPrkY9tPPdpid
TOINYcroIJJPMuFAwIWiNjysMMRG1nhHXYEqE3Vt5wVqzFPdSncRwIuHR5qRXv/0
/8kz+QBh7ArvOwETbh9Rb2a5utghEYlozOhcQhSf/VLdo70ZjDEUDKyfFhE30JyL
P8uDUWs9g6uDsLkQoTcxvFchrnQWReKc6itPNcyArLltaxuPCcVTJqbhZvYlWm1v
OItylc+SbwaySetXN0ibg/GPpEMKDzIpql7BDzzo3yzrLzHgCXUUMjsmuLAiY008
doht/yl0sZiR792knjeGt9lVYp2j/j2H1IwTRf+IhrC093kK/FQys1cYhsvj6DhA
E23anqxTZfjKBBW9+ym0FL0072KumneDbuSzLJr9Ni0aKijjP41KpgRDE5tnnEtz
+Cdc7lR8lM57d4y5OF+OEfRpfdkAucH4Gxtd5wZG6Pf3sYk0m6yK95u2N2ytA1Sx
V5A3iniD0z4JaehJxh4oIzzdaMgVkN9adpOicRwmwFmRbo8IOPAPN4xnqrNik/XQ
4QUi5fA2Qb3MDAupuKKPbrkYHdQglDfZxaEttTTQKldV5dowSsl4nqrBThBXe7de
0oqC/5yWvbAdCEPQ9G3Q5zT6ChBybSkMDtR52GraOlOpwoMYt9XYFYZtMUT2MJdA
kxiVw05TYylUMXclrWKXQx4aXofVaQhQD+Vs7v0QhSnfW0tyieAThXAYzu35nCVO
j7xljh/A5a/cRoL9WZUX0eAldD83Agleucio+MIMoafiaXejwDAK0zxpfbYI1Y8o
gDKnI30mySjPsZBB2x3/Mg5J3659gWgeqGnOqan7IVAX1oISt30WzYDq/ignhwlP
4K1K1PWEsGF5KCBSBiBThGVfHjmLSvXgieoF4j4uaiNqAltchcPQeiAnHU0rhA4d
eI/thb6kbwlXYGwRuL46KBYm7B2m7CDKB4/j6UWzW9qOKRj1vR8mDuMnVROo/ZV+
nAcmkKn+0iRl0pYbBXkmNFBo5D0KDEsAQHy+q4z2cux35GqCUyFfAvRp7iOyvv+/
+HFn/bXxoe7pIFvDmVywxOJEtKbZviWaFiQMex0Y+04/25B6LD/1TwzHxvLSmThJ
XnUZ1YF99f3iRkDbXmu3MXHyN7jDrqj77DEcH8iuJadufuO/Hngci01UQWz/oiP2
d2Gy9pz+b6US2WVpAgtCvkBpze6vdoBTb1SrrdA/gKb5cFwPi/YolEMoLzLuAZmX
uc2Yc1VFGP/vIck66ttXo5ydGf6/0THMc04ZPgZAlu3+ivCHwNEd57IZ9fZNNvDa
QNXoojcmxDAnXCh2ZmRuQEzX7PWXshi1QZ5hw5m3WRswd9DiaNRj0aJZz8jmlVyN
+pqEfF2t3afwQ/1+aaiQosGJXEqoNongrfyV3Hcqw+tFKcm/gHEFW4dRs4Ykwhyv
OEHr3t5pa0qX/igsOlVbWOTxaslflKlM90HZ5mi4V82l609x2dhO4qZXX83Hrvw+
HKlzD3oXs0iQz+gooxOFmLddCZIwGJfI/bas5zw2MgD6e+XjI0nvCRYcvaEKlVTo
LpOhsFJopX5J6o+GoF6gG9NeIf6qLVrU4wBMAndSiZLW2hmocRVEmFDl2+KOFy9T
ZTMk9niBI/f4Cb2RRE2U/tC+slHRv9vnfrYz7dNgrX+sl5dWnX0oluSKOQQYOSBh
ncaP58Sr94PCZCU0dF5llDGk4a6EiGDbOb6K3F2K9HLcK1vHl/z2wIYYt1JoRDIn
/fBn7OAITD68vJrTjI4RrZucNoBdGZUPV9WNjGB9J0AoUowrpB25wzVnfvoY/isk
er6xyf1gLg9VYLEDeXADcoxyvU9l3ZnD8LU3RWXSXiojn1/Z31kFuusjT4y4LYkU
WCgkG0g/LP0GUQNAR5PqV4LQ+XzQ2xZ0+wscVWWAE0SiRj7Wkv9isxo9N5qZy0wo
qPrIk5jtl5ttB/nIE4eJAP+Z6HQsRogFya3hwKh+oLPFWLZdVXQYp5np81t0GD8v
VsWtaAyFgTDsjW4ABadZlQ8H3cm2R/ae22CletEvgPBNHqqIi7oNtDoxoHSaRd44
oazlSzbEwTvwZm+DD7TNISA9eyR3po3Qvr9vItBna5Nja12JDQcxJzLm/DaBl82Z
Ap8KcT6MxVwNaq2MonVg76Sru4dg+tK+Hxg13chI3O1w+5pSjruHIVuvBiqp/f7v
XZqrtc/QwFjrXbe+ijR072Q7SdoyVk8El+h5vR/w7FPKPZt0U2H7xV6kXLgs6v2S
1jz4yf/sIjY9Cqp+NZzKoLrBKkv/PcNm3jgRveJJSPu6njUSWM6kichR7yOXEj0+
608KhwvbrRFClC9UesT0kmHOoH4lts9n9iDtvkjDVpfVatg6iys6YmQmnpVSRD0S
jLie+baNnNclil6leId07ExRl/U98G8TQBBzsX744p3/yms+ciGICakQSkdHtBAs
0YF5NTFab4fjfvzWjGc6Gk6QRSPMvW/0uAuC5plPMargw7Siabj8ImaOfmAYxDHe
+qaBSR7u3lbk03Va2iWtcD9s1M3y6seLM/LksmmYs9KfD1vSqb64GWiJLtTrCQ9p
03ucIL7XF472Ukkaq9fyTG61HIjLjRbPUDecCyTnAosgenuKkRy1orbjAeazZ+KZ
aRRp9huI30N1RMYqxt+EfEjsWfMRUDpNdGC18CmPsIvwZocS6ngjgNSnLs7fmlse
lRNp+AmRcYaKsN/zFzx/kgh+LyDHoJFiKUc8LzrmzWusufVQAePBhbTtgUJ3rIzd
96R5hIwgh165u1DNCDD56AQ0tAdavALVRUO1yFe/RuCytYF5i4aFFGmJBOVBtxn2
fEfqYsdAtQE31ppduhPFQsjzRYetOqnyr6TRF2K78VGj5OpnZqxHgH3MZ9wOXev2
yVfYRAPBAJRoFpEkqEGvues/7Kl2qttOf6vr+lyzP3fFuSds/8pwFrzbPWzpPfFO
NaKzrm2yvlymaRDN7uXuTXAIxajXyiTI8SkV+OwjEjVT6q/bZgnCP84RuaCPrIgH
ntLEPfxtkY8oNa1uc01HXbfqB5LOna3A9C63sRdIBnVlvPBtUkKCVpZT1+qFSC+E
IOOBENlfgQAA39E5dMektXwzKqKDncLvjITcrw4MvlBrWyVHGIBwdsjg/hT/NF63
f0iQQW67axBiOTj8xb8zR30l5CBmBxvlLZ4rRxIs8Qpo51bYZwUaktRRJcDHKE1a
frtjq/UhWFeiP1aKgnN5w8MhfEIsfQE5q6hAAUDv64cLzgfr1JWhC9VR5qzImWWl
xZMjCuwg453wxTLcKd0kYjczzHTYK9RJKB8TxeQaMTnhsKMKMs8fCnzO6nKcXj5t
x9WOAKjNaH0n1OmTKHgB/BDWlYnJqDPOpZ3PFy0XqooTd/Kc9etlWmdKu/G2sH+X
OpdXallIw3EQ+5J3L3xFyMwtvvqLXD+0FIL8e6kYi09YVdfrz8SmNwd3zBVCORNE
iYnMcOqygCiG/AaJsibmQJRPH6ppDE5Pc/fqmdV8hgx7BGl36RRPHj5TJzd/cEJb
kJc6U1nuTl+VWnk9EUK8c0cFahR2gfGhYqYVR4fNG/264RbY/sSEP6Z8V6RVOXad
XPWeTRoaheUkLqjm6HK8MQX5OBlL//un0Z3dUV5mmuzqVvESM8kocvsvn2yDiKqu
fbSzaX3f4VP0Ja5CB5d6iQfqpipZwlyITIog/ptYLQqceWGZ4yIakYixtOF2awS/
zMN64WeZhNh+fKrQ7bC5FJYSbIwZKHmarcNgUTKRYTvGZe8vi12ZAx3VPCITLruO
mN6OYKLXZO0zT+bldLdE8pvdusO/rH0jbF0P6ZkJadoCjHQTSB6LgIy0i3kMEl04
imNZJEf8kE+yIcX/5MUyYpSRBI26ca3eXi1VqXSVcf64IHFTfm3v5Hl82yRcRADM
JNhkoCXM0uf5NScKU0ZiiY5E51kLRbEdHwC/Ghml0PMAqaWUwg6UIcl2zvmRqCht
T4QqhV3qaGb09lOcxAZoq9/zggRfTOuweUYriXieVxZwK24SoAO2IadxX+CqpGiV
TNvuNsH5KxER8sHHQJXIA18xz2HGK8vO/cWxgeQoBH6jVtrQ3FcGD7K8YL8pW8Jd
9i6s5rnHk763mT/Gy+KQVVdVwLN5+sxruITAu6zcDQvjIQxzli7QljcmhNjMd48D
jk81JjyLECGr40MMh6BvSD7bnLAMJnUKW8og5HD30qZLE3bdOC7RhMe/gKu541TZ
/eRmXwHK2cJoICiPoUKuzGF+6/yw7CzROQ8kXznE0bgx1+PqqCHsLGXh+Soqze6F
ar6+ZhqwlPbyfF7hDaeQJUVeI3r1b30Qlb8Q7INIlqr5zbjvDOKnUz5a0w9uDCYq
VEsPnGZCn/PImoCu4qEWFzVZ0u7WhE0jveN1GP3vAug/PecnuOTCJVmU7uhL6qQJ
jdrDVgrXURHlzo/l/wow3LIvmNy57rwTliWXR5SZ5a8DpxbKdknWhVuU5RgUo6zK
7ruVfRDVEC+wGuXRO8VhWKK/gCyc/wy85pkxIcjqwXyx65r+TqLa8YDjv9aZCjKw
2r/27Gsf72UV0kWM4fU1RFES7BkOlccqIwmd5CqR7RcRTfyilWpMqlbv7wts9LS1
EgDzlDxOJUg0cmOYPmDgWbEUO2B73pJRVWXN9R4sAG65wIz+4sTzPcXHB9vT4ZOx
qmo+3GIqdM0x3E94GbX2pH/sV+BWyD/JOHd3Im4vtcBNXkcq0slB9J5qzgbKassP
omjv99wUl194z5i0gHDp7J6ZMxP5SzFh9vtyWRpmZZiAGwZEU7tZhf+v5vsVQmiM
kjhmzMNqGS2Uxfzej7NhLBEWoC04Cn6sl4VZmY7Ck2Pd/RX4q9hAnXA8BAGF0xX/
znjsrRvhaOGSh56IRI/J2UEX6fUFBPrCpalwJQBUf8P/92mj+MhylpCr9R+gyiJf
lP3NCUzO7JaGbhw2bHDqneF7wVhwnzCOyoDbQMxa/oBtIuYmCWcZFJ3M4cR8RKr5
kfCiBp/Qs8jllVKI/BNcdb48wQI+WW1bZ1MXccucFslhEOvTLrHZbcfq3fl5egqO
7qq9qfNsZ8OzhyY5HryhcBmeqYwEys6LhVaXYPWNYUXrLYQCq+m/cHIBav2sMWlR
+Bk8S8r/q+UKpIkldjodnZt7VWk3diKpJcQewAzfuprZuHL6QEjYhMrTVb3r6Ohs
Ernu7NWJLzOfzD8LsHXzzfmpEVs3ZfJBQqPdLy+juJKTB7Ll+cRVztpTZ3XL7MIP
8DRDksE19uOUkfFnXfgGSczUxditvP97nABMI7eCtIZUMghToE4WxD9teRceyzRH
7xER3CzwsyXbDXxFiqs4VOWtsUuzvdZuO72Iok1KzikcCjEa/5sF55t8J4orlNro
5ikGMaRx16xqpqWNZg8gZUXatl2IOnW6Oph7Fk9UeAhb9ZmVrjFkaGRVy+HAOqAf
IQLyXMxA4lO2K3bEMlq5cUJ5ly2Kd7Zps/7cKHZKoVDOn6m4V4pY6l2vMXQKj/S/
MsdsWz7pfg4puKB9LHeMinerxI4I+x7f4LDirhe2zbhPJs7LZnPUHt8h3a9qcL89
crGwKxihTkGm0zXaY0xbUmaRlVbP8GdowsIrn4Cu4W+5aCGPm6x53UjvcaaSC74u
1YTVrOUJn02qVeQtGDh8X7bxwDQhp4nvchPGugaNPyUIE55sxMGMQ+KtRa3hrHOm
gwc8CQucKzksjvCzkk2sy1O0eOTul2gRCWIhpzIbjHTTPFYsku0v/ThZQn/87l3A
f6OS3AYt2KzAaNmbcC1NhzifF8wsNslshOh75OZAQ3/lBVnBOJlFxJIwi8fIiut9
iMNOAS1l+IEmzaYaM58vTpd63FYIJ9E+g1LT5tF6cu6gSL1Cj+EosJphnKM7KI7K
v7MMjYgcjAcRXNvWlPSVFkc0WZtW3LBkEqbV3eO1zwtIR9WfJaXOk7NZg1cQEmmn
Ugl+jEsxvpBj8pHSCfUXgy7KCeR59BCpMRqgrFH2Gc2K/VksXfOCJl38WInVbMZ1
cpbq92cRwX6CK6/09kbfS/22f2lHJceUOL1DXRma5TJFEw4o1X9PtXD2vp/Be+ez
QhJPpapVUhhAM9i0H/waQMbUgS0PzRf8BpiQl9ESYNGwpBgbehd5cteRwewr+8lo
/SEHkvlnHkuVh2eqoY47yU7rx4atlD2tkfguOoeoc1wqASjtUDQhK3p+1djtEG68
zyPNGK90z1S3NVHg18emOf3H1lmqzDM8j9pPIx+cJSxzOY2e2JkaKnzqi0KUzt42
S2yINFU3zY3ipeDagahKLC83Rz5oG+oEGuc0TwrWWmoAl9/rDiU72olGjNYsWH/m
BXPjBYUd3My1fjbR9EaijhJjezWp64aycnx4SgdEK0ZMk+mWGMKW3oPIRxm/aefP
cuu8iDV+jeQCxvuKMgIief8yNkX41AFzsPiOd1KplCo+EIvHzqXVC9+TRr5QCvBZ
bxf8aH6aYdTqKtyday/aCi8TkCPdbwqMAluW2IQqBhXwc+eaNQw7VzMfcCEPRRmf
h3aijCya1yS3clSas0r2JfOVjKFMky0AFbks5oflLtrVOiOQM8et+voTxfc63VHX
2OYjCkgxvm+Z88re7z/jOX+CdvdDGIoYr+CyC+JeAjmcrCXyRhXNm/Cb/wwglYIM
MZ6t31JoglhvhnaFmhsTCo0FpKxRr441UymWHLttlu8uQ9TVJV8qi3JWVqTfmrFs
hpRfUY20unwCbDbLbKHasuWkZIvEi7TsZb5XKDGLFaGmNnINdddH4LE63s7qv/kB
6pHZLgS3ldkYcVfiBskzrfKmuxy2V5j2iNvExF6zxrIoNRsxQUvsO9XxPM2RGSyy
YBJjJJBoKoUCnLKXqZubdMOAxtuB08m3Cam+4yWJXF0ocTgLYhwhW3ApgD6eUHtg
cTWnITu7+9YaK4qQawWmngE/kW0/r4snYENCMefqAe0ivEsVrjLd2huNgjfz1ujG
zvun70XfTVxctDJdU2JvQ9+SFY90eidSj2l9e8xP9kwBuaMRZ5uPfIeMgtKTHM4Q
gOFlnQTrWOFdyazlON82Fv2A5PzE6E+mtorPEO3I9sImBtB3NITUrB2LIVdaFMMI
3VhKV5eU7+g/MXaAyfexT/gGsqyVeVrUPQonSUYDGHPD+5mb4y0cg/rZ4IWVZj38
JDNEAmNYtZGCAi7gWQgRB6WLDxc01S+gW51yDRo/pe8LNo5VytQqS+el97gjU0q/
FHS3fMNk/x3j1Ah7HTfMPFKfWJTCbkUbgYOC1V9X2SWXz7Bs3g9vpIpUe33AlKo4
nSWpdm4hmg2l5uL00tagFG37onkMyvWBiXto927ZCFGc4oT2aBpgtm0AXfp7J5EM
tYYDSvhv5EGlRzhZ7FJErAdGVkd9o9fZIuUgywOXJJGYn1b/3QmBdAybkc8UMLd7
i+OqqjUYcLTZocdCc7Plw2Q5Cb5J6kmvvViNxKmj5l74Gezr98km3l66L9JJR4fG
OpfMPVKQpHCG4TF12Sn+zH6sKWbs8h6cRCCFrdaWjy+nX7EhhGbPsJdVr33HFcwv
p/JLd4i4d031vvhoyw5ZhJz6iHkNbzZD7y5PbRneKEK72siEjgmU3lAIXRCd4gOw
kShkndSrfsSWFjB+EtfWF7AZceLoE3nFpGozasPILV79OoLiSlvsl20cTRcmh01S
vjp5ASemzFKrIjNlI1oxaFTMFbYEKVpfUnXcBQbNONPhXKsppxx8y/5KQdbjcr+7
8iD5rc6Izf244spJMY0u6/qYN0lq+9cfkzHIfsdB/F272uixSh5kb3IIJYLRHT+c
PPokf1OOq0+PSj1u6tGW4Hms36TjO7tFVO3Cj46b1MOys0WC8giVAe6S8cTInLA1
Djow9ghjVPPuM2na1R6yGEpub1hViWqt+Fu2Zj0rJtrTt949F9JKAOx4WtJ5oRGk
83xxmywbSSdjznfPknaF4zdeuGoCl90v+QpyPKPGSvp7fHMK0b5V3sWIGt6y7PxN
ch/E3Ov5SXS6oOLu9XW4wAaav840GVV5AJMgSd6tr0BrV3nwaHCAYuTm28z2EjoZ
m+4cxmBl892mqarA6BB+JjW/J9BVEO/iiBYW3gPKjUzxs7s1Cz82P7ypD3HQpP54
K8K34PWs5GwKTjbHjun4SOSEPftsspuBg321RYYxNpzNajLOFpseGeeAjjn/6w0L
ZK4x6cVWFwO4hcC2WdtYy75BkKiy7EGEc33hqOiIB3OGzf+JB2UniZqWcbJZcNAp
Wr2zWAbPDynGvN1zKcjBVhdWfGoJjOFmyKvybhzSS6aEgqCqP/2s2hOdQfkh8Q5+
3nA3Z1yYBvvlHnD6argeGZzFpetWAh+zDrllhsZUFYlSO95OlDFToDw8wB32NHWn
Wo7MNpLIMrSPvuAKiGvnsc7fR2p8Rw7Au5ynAuds3nnRAnWqHxd+CmUs8QkfSZIz
V8Xi609tooIu3+Z9+9RdL74nyUGyYLCIgJwB0BpZIIBF0LNNw06MQAR3re4HnEms
w7R0ezTpepB9c2G11cIsyqa0tmQZUKTsKLOpE6rPu8my+acW7ce48bXxVulkuqcF
a4FSml6tTQBwmknyqI+O+9h38BSYZX6dDkMtVbTRozF4c7vudpAXJnphg3pSAsw+
5gSI64QYDhc9xc+b28o9EVpetL1BOjb6nO8N/71FKcUs7Lzs+WoC+UXyiw/igSqh
qys+nEwGWItuAvgLWjsGaC2Pq3If3w9e71Rbl3xRyygUDZ7YSjU9iW9Xt5jSDiL5
LVS9CCKqq77NpwaWYrgVy0aIIrBul2xX7+IDQ2hZ/9NPbIw1tzC3GI0EYmncszf4
uQWs9eBVdM7XuVlNlkJVdIvs50Dy3CcyrrTnB9NEogihfpiDPA2S+bnWHHrlGmT4
yG0ZCOj4uRSfUJYqiapK6mVsmIAyGZpF8oPXHVm670Wfl2mhxrR9pVmyduUpjmk/
blEAOTCMkkpCEPCPRYi4FCOb1fcg+Wq0O6H6E3RVl2rAFPW+A+aviVcvGOyAUCVp
gWlMkUHr8J1rbpb59jein3MEXnXmemn0/lE71v/Stk22BjyM3nVZNTf6De8Vuzz6
4iWYF9umvy7BLpvs84sHbbwNXcJFW39urHlRHxg9o7RCrPO7QF68TV9dhqTh28pW
BRdAXTzGVNtsiEHm2KrJ8oPXZS6IwqsRIV7l0frjGkPXKbU6wk8j3Tl0wBzT5Ow3
xZFddGtaxIJOzRh5N4SaHGpLPaku2uYIiWB0aVdZ+QaeAa4EOkvm3XJqLQlYUnt+
JuIH5q2jxZSRRCvCJMd63+h6lRaDpSWZzl5Gel90tfeECsb6Y5sKEUaxIp8L4yOa
jbOQ9Q2u01jfKM72ncEF9373U424XC4VQQZfoSnnBOR9hg/6Tz5oNuUU+8SdWcSX
UQVSTARQN1wdZrz626aAby8/T15Ox2XXvrLhh6bkNM9+gyUyKCPmyJ8VUG5KVR38
HDuUmEESBHhBPYXTGpOsUTjSNTTpvwXNjpF5yc/hc4evC1L69qLaP+zVaJ6DQIDA
P2yhChXFNGWzLMD9iZfAdH9YPf5y8YblXiY5/0XmNXRMma2zLZyxqc4j224NI9vy
qMLyy/PKQXWmidOgHx/kyfidcmhqCbzihprc4YDLa0O0gbuj98Wu9TAKg1fTjmtN
hDBhasy4YMxs9O733wAwIbCtcEYdrcpPzewIEfPFWZQm9hJKbqnTJ8YuBrYEzvZ4
DmmGrzlBApowVI53O37qyyQtwAq16DuBCvlRknKTa7Vsr/5OI7JZkWsgril32jwG
fP8s12GJDanYpQge3086FXNuyW9jg4quw6UJgXJ8/hy0ESE972j1OySLAMhTbfHh
kZ1qNqkEEbpru3t5nCyyizT2304xY0h2qriPfiZipvY/yy2YRdQBaW4XPi2+Oanb
+Nk8nsx5B9s25Fq8bTK2piJrpel7AnD7PrbF8OuGuVcN88WX/V1UgRQth8USUfme
29UK/guwjwbkGigMtOqBLrwjmdwoMd7whiSlxHwd/RYFMByiLD5Pq2K/PPzaVhAY
w+DJg0lsOClFr3I231rqI2vHi2LhFT6ukVfeU5cUd4B9Umn9lNHKZBgoooNesuhK
9aB575Thw5mDWb9zxC6GIyejpvgwQExpPkdo7VfuMMNH6zY/1TlQ2Oi/W18jaf5e
x7i5omE8Bi8A0OW8ynvT80yv1D+RpbIvqjXAWvs34nbca9Sy2SMFr53DhGTQc12S
DozKreSHvuhq0ZCsaQS4UHDxtEeIhRRVXSNNG4/XUl9WKKchlybI2u9sVChjqCC2
4Tsn3qXBkeeobbCM5gBEmE/Q/JAFgbysGK6GXcFaq0CURZF9cSWHkYVlRSpyNKUC
/RFuK/2roDbewP8IV+fGPRgLpZbTcSewmEkGnNW0bEg+6wieiEC4XT9rvduSI1jG
8zxXnx+iQkLftlM6udspPWRHgYBk5LTicFp61/M5Yu2CH1rCwQPJqMDUN8G1LZKQ
ZsCmtO5LsR6T4AaG2Hp6CEDMcts9hOM2twM70JflSWd8nqVSb6yWwuc8rD1twKtc
WHeIMg6Mv2JJ2Iywjkr82F3qkdowbqzS1SL9Tvnj/hlBd4w6KksXwEwc/Ps/vxPE
zkX4h3LpT7upOB9dze8gO7t9NvvspaB0nWZTcLNq94xvLAFb+O57PSnidW6GMTDP
q+Nlx5WayT5dLYE8gSCvBzHCK1qdgKpvfTLc9KPSWsI4BQ28IKuO7rjCVAGqVR81
XCGckPpuhFEFWiX/EnVFtoKPFVQYO67dEzXhK2xT7LUeOSbCqPaW6SOQRtOCHf1Q
Tmd5Xbp9PVhAnWu0MC8DMv7Ay0Z4Z/pYJe+NLvU74SEvC+VXpPTmCFZFTDXnMdg6
TYGySdjh+ZqcqdMUWBZdO7UoIbdx7AvdBXcD1hUK3OooJ8At+rBhwBxOfl3Ze3Z0
SrC5MAw1PQjeVzx61YPIkwvUBWkGIlz0nnwJBYGr0MzQrO74ONYEcIVCT7oJPLMe
AjcuJtgF24YQA00OgNHbUP4ulow9oFh4n+9zNYWIuIWYrQTF9Atz3KnddUhOKOqo
vmGFrXi0IJ2xw1mLyRTVchlMZWXwnHBHW8dFbz97VJsw68r5iJA6CFZytPIIr3yM
90pyGTVwua5WV59eLqj2rxry02gj/eRput9p+UOQ5mVDHx24Fla0usSJKiIQxE/O
s97G+LZVBs2WWRBD5ZSCNTjKj8z8+8TsV2ZPTloA+G7XPCX7NKZwGyM+Itwv8pHr
TWs/AJJikmTIPB0Vkt33KwjhZKfZL3MgeMgEbNvMcO/e7L+RwxaZdKxcO2C5bqOh
jtor+z/BpcAWalTTfRmz9yXMntje/A6W4K+23PB2kzcizRZEG5g2KBEbe1ev/FY6
+7z+AJntOr2gA3HbDK1GWXEw2AT1K069pnQZBN137mVjExGBpRTz7U1Z/FMtt1IX
74S051U4MYvqoqmExtznLjV7TTeqSrplwvymUA4sWw9tYuJLYDBlPUu2/zJMceI8
QPaKg/6hCxHEDhg90xnojxxipDO3G4rm1SPhE3TjbAZhs9TR65l1q9QLL4w2detk
h5zWYnmoDenKqShOXvKOucN0iPrM6jPq+44M5tvWm3Y6+hZWsg1EnV3S+MAxQsaF
CM+wBcJ2P/SblaMWZz32F1IPVcq8nkNUGCYEmDjPXdj18TJiCmjhlpXdP3RZlbjZ
DYUY/22eD65FT0vU9IO5sAjUT4+RCHkIWPhx3TWfB7mHqvKaYlrA3IzmJaIXROnF
ibSyOo724N2gNAno7oGPGxiGJ0t8ms3E/uHwLWwcCZhDNoY6lF/bwsUCz9Q3qbxf
7+mEqEddpx2E4GL3OTlKF+5jXL2fxZvtoUZCgGH6Rg0JKJ0Xu9ySSTlFU+C3OPU0
0bEeMb53F9OXr0HDMZg5xy4SUkbvR51b8cxDBsLzmD7ejOh3mZUSBCaJPU3Q8bIU
6qczjbK3JebaPVvN5hiymSSQzZ2CywQxFsjuEoUuHjXGxMWhxtD6Ftz9NW8F2KfX
JmDKKQiIVUHCZEsobEPldmoi90QAcAqIYP5STADRyuKjoSEB/e72erEaGOn016DF
rc39pmVbAMLXA6p/HnSYcSiIbpa9hi2jI7WOTsg2oHuXfIwcvRKL1tNtCBwNS//M
8xRJ203GzewLwxEILiWFrDNrgSL5wMPJ1OsgcKdZ9gWRDsMk2en6+keCiioehR21
VDPZ/SlzM9ry+Kc+ozdUDE8Kq+uHYEX0pG2CJEpkQ5yyUWky3sNJVTstwUenNz8e
4ow4NjtdQbxj4OiNYJd5q/ut9rKrV7YBtyU9bxGEEwqn22sqt5kAbwuD3Me8qgsL
Who03QhNogR38ccJG3Ow2yYu2NYXVSCgyXReAFZrni8jhhv5FxwkSQmkFz2cjIWz
9MPfVsKWZoC2sP0Z6YYQ16ZBq4727fGf+PMavm6xHu4NktveM5TAgqVMDR80YM7Z
BJgSKexJ++/IgOnqGpaDi2anOGlX0hcC/HSphG0f8gOVYlt8u5Csh/mko9/3GXpj
/OfJxU63xCjfYWf86kge7c1VjgEiBK7S2zAIfjZnF0WaH9NQ93UMu01AWqe20D/z
DvJuRGdzbSKEmqHA1ffGNSdT4cMJUreKtWXCY7EmNCDFv5BYKjOPW3JflB1fohWy
O0l2ycrm72JNVt9h9nLI5IpJgwa12Uq2Gx6hYI3TIi6oFkQs6UxuYCapOMB7QRqd
fYQug3kRChbFt9AS79QTjV0UHpVs4IOp9nyc9JoAJRLeIOOshKM5jBRTCQPstZSB
YX5KZGoOPIr+9irbPdPHz+k/nmOTT576MAN6fvLNVbadpmg7yEcQlv3Z4gQBREIg
P77xQOQYVaYG9jsuwtIcQtvArJOL2QldfOqWDk6464N22kkiG8NVhWEgB0ZAHvvl
dVXFKZf6wHQGQYLcdFy1UZ/6UmwTW8aF3POweHS4vLvFql28GAv/BpKEWf96+XiZ
u3BoMtp4ZMhVDeiAw5B1RvzJJUix0Ak3rGCNHcXP/3mFe889+7XcH1XHwwNlMJWi
LU1NeQCWvECm3L4p/7U01hUQRUuJIIgdYBxCQcHbWQzw0RnBHHIIi5x/lPMFRRIK
DEAEziy3dsVYLE3xlR5qSpvFHK7rYsWdvCbkLbAAc3Nelpfe/T+K7U1e4Nuaz8Rr
vhUsvxyqFs5lEG4aj/QfMm0M3KmGuADsfR+cWDV1Ulrc7rgXgsHKcrtpYkQZKaT5
FWaNLL0HNr1R9TGTNA9TEVX+0dH+5OlSTupXNoQKSYG1xpRTHeze3+i42Vi6hXOD
nKSxrqOl3r6R4wVgVHwAZ1kMk5tYoOLEZadGd5vV2Uq1dSyHtSYPD6gROSMMXdNi
2vmpw9VAi2E+limZk67ZbsaazKY+pAMElPEw0uTK8PQ9AIhe2a9/sOrYKTPJ16EZ
lFvdaWaitftsmSsOUCxqgAUXio5xvtQfUJysQIva7hHXsQ4CG2faX2+6OjMYIkhe
b1kxSFl/P/jPNBNVHSoLltrokxNIN5Q3b3pf776CWMUVBG6VAuETtLK17rFgz80D
1HBmeZh3+oxzjeYqOgGxWdZEsKBFf3/nUl+cU2z0X5GvAqlRqDq5svltmIN9NASg
INPKQNNO2W/4/oWBSaQBcm1tj+oPxk9O9hGFxQmC3W9LU0gh71/Naaus1KJEni45
/8RLNOK7xxBQqvn3FLtvvjGDP7AUUGJhHiscquVEGmNNCBqfcjOpxoYYQTgCARUU
JRWHWJellgKaNwjTzOfklr7VPA9j2fI3npVVIG6H7OJbfACuXppKGBwktALaziAk
bQLeijmAb4Nf6+VxrNindanTZwg4xIEi105b7U3/k2Fz8WXHZr18EvHblDyIvms2
brpe22H98EAAc7qRXzuVRW1jFOe9JPLSH+MC2b+nUGP3IvzQRZsDxkGXauz2WXn2
X3CPJiUU15gw4DFLutxGv/DkfZIuLai6Dxncy8eGo+fvjbK8RQOW+2mOifZFnuTw
BGEZIDT3/fYMoIZeUcHtgAmHpWNDtA8HhH2xYHPe39lkTX6h+5caWvaLuAuBQJDd
Pjqxr4x44wC5hjBVyrNczmRplSMyCYrR/bONqycsJMNjogv8cYl6L/PCYQodgGWq
04jE0dYXMK5OVMtK+gnQILHeysmglTFNtowRJPUZmzBY4VUmBTmG+bsnSiElA1En
cnd4E+WnRaTfZrv2ulPHwSKnesCi2jGTTtHZDc3Yv7phjylwupb3fx1W7Iw7iNRN
GPiMeISOSHr/kdqxVvCzI8cICtAcIEeYYViSpYN6wcqFQk0HYPCc4yKww9PGNb8+
yItiEx1ZYvJCgz/3grafLNAJf8Ssbmpvv1J1yOHwsO1iM2KMfgaZVe5oWCJk7K10
ybUzcviVzEX2mBU4XgX9ofYp1ytEoXafKBQxsbMlP4b4DoNvthfsnCWN2hjjqEzs
J2UAgvDmWuIpt2kkjMp6TIN38z2ZQC+bBX9ydv/2k0IHGmuitVg8e7R1f/s708+v
6q9bkg57k0BuKcVtGw8DIRyanpAZLGIexzsqwoKVUnID7j9utpuLDJc3y7hpKqzl
BlR2Yioi7afNOWqnsidHXvqShPFU5YTZeziTJ9wjDXWp0fyDX0sT4CK5LKSPKhg1
7QDvO3nlGtQM4nVIy/gm748mSnl+8GFVCXT/eV6u0sq/l6bJszBxLhUfT6K84TGW
8zjGu2ReecQwF2gciOU2q+01OhfiNZlgyfncSebRVIgUt5Geids9rQkpVdclMKda
6hpO8umHUhjdgYgOGW4J5NWyTpIyQdG3vin9t8rrdLOQJVF4eFI1W1Rw9NHFz1gS
Y0QWvODRkuJYetx5g72U9t+4zyzLc6WwZSVz5Rt8i6y+qHAOrek5kujDhk6Mx0ti
N78VE3OsLNA+YczbNW2WMFgKHaFRxclyOojOlHVUFBLbqqE7DXOPMS1nInp7MhUT
kiI5KKTDaZpZAQjQzLVKWqDbm6y4szFt8ZUBU3b8bxc242Q91+m3I0mxZdQ0L6AV
htEy6nxmmpf+gufMPmWgbuPheYSJjrnvTls5Y3+fU705fjXttFPH6jkkZFlz0Msg
JvdfpcHKq0mk99ZEKyIIzsbNjGbOyTW2Mu40tdjvWvnXXzFLh+I+Lb+51keo2eAi
7e6vUoYrFj6i31nKaw+k+VS3QUpBYz3Fa/ZtFJcqlWTWW7o849ZNEUDgLfoRTc6v
bsZHhlAtk8Qy3ht45o1I7nFImofFtVEnH39NM1Wr+eEhbLOKWNzMZy8dFdtHUPI2
iq2zCaNYjrFRrHEjX/gawsqjDL//RFPbU0il/MgoD6HGinwDEy0iHzZuEdPK8B8A
NNGZI0Rk+2NjikzH21Y+r9QrLeu2POaTckHhiiCsxZ5ltOwG5ZjfVdG1CnlFd1Jj
JlTVr0Zk1JFATLfMR9mzcf8x6xvNXNdRZwOEs0FWc7hMag1x5kxe3wSUE/KZDLQc
WCU/CukleZEYWdv63StsygKOPzR8/4SlzwAOvkIIJby3CUdVYoMZL/lW+ULD2SQY
LGf+qXyMdcvZAG7+4wcU0/10B14guDwHoeRoSjAzrSzSHfWz+JSZm52RZ7MyrJ39
yqbssXQUIn9F3XpcIvH/wndOcdDphpUSerhHi5dDH37pmZx05SZqW7p0TaEDWKGP
+q1vEi2gpz3kznsMSQFM3a4DZh1bpxWXoIHNeNFUVD5wQCh6OOAAIkUXQXV9Uxnf
2/9E4zhM7ZlIC9fBzQivjdG57wK2xv6XqY1W67XWBLM2lw0ZVVxGRQmYvsVX0gIb
h7QBH4CzoPDvVo0kxIphFUio6dh6ACewivWQ7gDaft+P7TB54XhtTfnD94v1fkv8
YjavddwGlRiDd/+EOTs41kb66U8pPC/LYj3yMGk6s/UCJElZYdx6Us8Bg3332xQB
N16HOiokJq6WpiWb2x7fnjYvj9dtBhHZKaxcgbYOOiFjt3fdX2ezmiQDqGEE5hyx
/b1DgavBNQJIjClZaRrBay3hHxHXlhWqEvcEpNJ5hUFngL72sz3TeUxpNMKesIsE
xUAPDjcTzqAegaJlCrzZxGdJQbfQ8rfzIh9jsZDGTiQzWzlIq5ln1mERCUInu2ZX
L9yjVbcWQdRHr4wDxX24yMv9BWVQb0O12Desgoh6oWTn0XQ8R8wngQ7NnyzweWet
/Tq8pC7/9xvdw5i4qB4v43hiwmeiBfuxVNwZST3T/UIrhF6Xyjw3eHXAdZjS8LVp
e57GyoFQaghJLbN8G46AXFXVC5JrqY2x/morJDh4YLIGpA40C67uQ1p7K6gm52YW
IhIyTLoGdA6ewukkoWlkwwchQVTmZSO2Eb5jXaSN43eQjs+g4R7WdVcBydV6xdDP
bwV++jKEQjuF+1n6BNZrau+pKBChJelhJAzAANXVLmyVMVoFEDFu9tSlv+DPBRVI
BbI86lid+lPjoU4tVZ1jejG5HlxS7Ai6gOAEmt6ph+eDRLudUQ9k7Td0HyvitMDt
u4qz0/gom5Az8V60LPAIQVzr692NL/Xr9eOneVqILYG0hjLv2taZqHAbB6rfoh0x
UsHDte+j83dOt1M0F4S2M10O8HTJkaqtDLanZsbChCP9B8AHYSga8jzk1ldGsJIo
PFCMwSdkkUROujPlNX7Hy0xvntR0lYbwVEmMM2KSIDIZz+IYGSxiL7r0IY2K9cB8
a2dK/Qc7AeuWy6tdoTutmVywgxIyYVQO2nzgAAIBCQL+9RliHuXjNfOCHzxX8/iV
RKOwgJVPmy6/lPbQWSZAZHI+DQfGCtE9b4G5wGMZG/UrmuIDKXkq6tXdLfqb8vdI
a6BoZGhwveSFDfBPYE1Jwb4r0P9s0e/K/7AhEEzSe2z4cFM6yKONgmSUAbAMpJWV
pE5whVA43fm6GlNk6ti9QoNgVDO+8GSTHo6oD9SrjgdinitVwB6OVSom8XRl8zBX
b5Xzb035dCzI9ZLcgZnQqQ9uG3El+Tg3c9UqYD63F3up7r/JrGpEPHLRLKFRrQRo
vuqassDDBq1RoOj6hbmHVYYQBS7A12njnxVuckS4QZEiv5eFyrxYERt0xU1SPV0D
weBo49i4REK6yn89bH1jtm2eBAPCshk9rLHLSuRTY9Efi/EGCGpItEEn3gEBClek
etu694OEOA/XlJTxqNxtcyLp4d0yB49hpFLLxtJaJn14cgcgTHV2g9Cs3pwiO385
eegFMS7AuVZNnTlZw7m61ZF0weyofch2d/6/PDKFyy5lfEV53RKqZ1rYonzmfC/f
E1gxyKxGdo1cl/1MlcO3ozss0BmPqZGzoYVGvMD4/D5s9qLr6uje1KISphMQxLAW
pp92HUh9AclDzsdkehCS/RVw9OGPiR3Tp2gy7CnfDgoRSTlckTL9EELyWAyo6kGV
UjbJ63UIDzrQMMMT16L3RwiOFE0BDDMnQ758rWK8SI+ej5H3TgeW3bTMVxcoW7oE
0m7caZGOCy0ISyJ3g817VqKmk8b1HmN0An4usKkAKa4ec3FsFyPT3TA9hAxYaeTU
sVkytr4EDTo1J8mjdF7rSB94wgT3e5NwlXHGeuNQ5BIAE/XH15Z/jlakFMel/ZTt
4Lu1Adfj8wpYW9CKy6Z/Q4n320BGSaN/rVmPy2IjSBC7LNQekGG8jASMvh84bMXV
t975Z5HBY9a/UAF/+4PN9ErveH22I8R55uGoV/7epkgdAauFafL2S1CyE14OzmBM
RrTId4iuK0/PsJ91AJwZ3a/G/Nb8L/M2tKDdSnBA/4RaitlXUk4lvz41iNNy91cH
wNZ52SPweXz1l9uUoh5qjpUF7vSX3jXU0MNLKoVoUZWOfPv5CL/96caWqNeKJaVq
tdr8pW3Kmkx50Pey0prc7c5UpTATmLFszYcbaLG6+w56Lj5j5WbV6m7VhO/ePVXG
Rcs+1pIU2ETLXsWfcOQ0Ccel7C4VPRoiiRL+ies9FQE3c2ZUc1zatJa5BIWh3QtT
9Zb9ESDtyl1OmVoto11KChIjEfA2rL3v8Kt2hE9FO2hCvcqmmQvd8GT9cRjztzPZ
WD9h+gjye+rXszq0rQYlmwYZYBXbFI3M3F0uyy6frPPh2y1fNugHOnn+4uZIjpar
ynCU+XsJONPYpjCczsTuNdHyKk6rf6NGZwYQ82pbApGPhLgvncTJUVC5YN57MBcq
mj/CriuWv+YSx0mkbSAU8yrG9rZQ1AN51bFuAO249FHKkRBrQ3y+1yE+Cvbsz5pm
ZmaEP4f0m3Mx7PkHLfEZt9qaYVmkvFtxXThQGd1XSURDodX8dOqG4klYb/ZfjmlX
GDp8+qdYLh3xwhQHaUg8gVkWAM89HuBcCC9DjZxddPUJqnWVcuGEt37lf9BCzUEz
pPz6wbzz52ZVf6nDpKC8cAdhYiT6jBwjhIzllvujt+RrOvgoacozDyI4KYbL4ISJ
sROnlNqntHIvScZRKTa/pBP58/hPSbeu4EALgM5G1kbQ3QMEWT7SG1anC4F6kr/A
3xXF2u3qcAh0FOMcxEnROlJkLsHShy2GQHLUl/12ZNRpTFER7zNtfF97R16ulkIm
FEKbm0yopStBkJe2vEfrvQ2fykJ2prdIA5UsAJZK+159bQGP8Ebci9avvoPz7wNx
WTMRHJtxUekn/LOqyZogmv2RN2F2y5jZ9+1fWmgBWowGbkhivTJUJF0SNhRCXKnL
gDn90G+bbNcFKTfbTTzHTYKqg7ddWkAiLawrcE52i5G2IPFD+Jkx3KGYiaNZWuQw
yiaDpuKTMTnMPh+BQ9rlO217eY9D5hJwXl0IVAoFJy/15KLBe8ORUL7egl81aASR
TTTKZ5bwpKx9/gjVczJl6f64gNwbnDBwCQsI3QMx0r30HSYCRLb3lhVfYNj//ALw
V/oIilc6X7EyEntbzVeyQl93roXI25S5rOXEQKEgc83tPrNZFLL9ZmQ35HNAF/6B
AWDf9HF7/5tr6m0m6OZRo8bW9XNYjYAdAha3D/Bgodcb9fZ8sLhiOQXKI7m3KWyR
ylmy43VX3PahwdalYqt3HC1mMA14oMQoJlQ+9tnRNNHKcr9kz8dUUOIoKB8WOPUS
xY1Y4RdDrdIAg9ukoDJi8nDtUi/AySaOv9f70Czkwhlu4PATijzBiO9Z20jHlbqf
zJTi+RudgIFg3LIHE5eLaEzP2TWO0kl4DQzKwB5efw/SOprUM9xpQyGvipBIrVNg
Z7eyUiE4/NkD1qAqIWx7xvSht+NpaTA6+oKqGj76POv+ljwbyvg+u/EkC1jeu0j8
MdWcNjniYI+M7bQ0EFwECoNENILMBDryGlhGPfIs25J10eRkOUoBzKspFjYcqXu6
zwruP7d2uyApj5AWVIHFper6FnxAWKE9R5TABalDUzh7gvIwx5dbNQjAbXmSW3St
bSTO0CQIYep2ubpbueQ0wjYbMIJvmI3CQWRu908N22p1mpMhsH9wGKJQNGkNs3KZ
XeqkediFCQYvo3oBY8eCvT5wvPbJ66pKLkuKiYHSkT26lvi7ON8pMEcUPC/ojWln
vLp/hGnSZrWEjtGiYMf+6G9zoeiCCmhS4A808REBKHtJWgfFmWz+AeiEf+bZueiF
EQX4MPYGBu4OpHSC+M9tRsIrTJP4W2PtLyMUle9K9XxxRvbYN5dbfDyxIiP6o/re
b1SQ33s7CPoat6SDomrsIqIwR8vTtW/USpHpQxalBg3W5qWY1vk/Yzdeh/OI6aS8
ldGT7svsmjnQI4cQjD6491IItAUDb09f9fBGieo72nAKixafljUopfvJ+x7BhwLS
Rv8S5781nvbs+N9i15olYLlhstZ+YEBPyYGXImbyn0CqcGmwylsM7aMln90F+pQY
4hEigPrLgCyy15T1qS8NwV7b9jotXJ+8OXirTlDrLoRH/m8sNw/P6Igpb6C64oNu
Vv9y1Uh6akuP5g2U9ZGAnObF37Q6QhBPBbuF4kSycXCkSNqgygGw6kIDqonhnu7W
24HDwmXBJhBUQ/cBoHEeTG1mIZCFRex88RjVjk6YZNdHj329zCnN9SJtxZ3os274
gjTbn1+xAFqiBw2GHeVwmbjoaN1MvN2v/NUaFjrJbic1LSKi0MsDKHIZ64pHct0q
c61cMQiAJmRN0gJxGMcsz6AjOve4ogRaO2hWBVKgzw3bDIU6BCqYETGM7ACE6MkY
kiJAqWqMjV2E53d5/F5fUgc03BqImuOwoLfPWRe7f3p0ilTitvRCGxXDBpaBZsX+
NdzQ3jcK1jTIflor659dFqdIC7xtRNvm7A2NapPoqf+12yK6hGuaC/4P4mFsIpJp
NHYJfUcLswZG8tMLL4zgkK2iJutWG+ToXroN9aOfkf0XmfVt3iZzzdplr77eoFyP
yl6NfbJtBGxgGZh0WvR/KrPnPs/72eJ2ndGTrSECm3cgev+lhP4W8xei+peTMVMD
UasrLwT3hmLFwfRIxSCt51PiibSg4hakwV5o1pbZb1ZM6VpkTVG7JkBXn1gL35QW
BzNX0fSucwwoyBqMo4B5hDwgf0rYYk+jVhzYtyBL9LcnLFwkBljgvYT8FIBMIQFG
kJIgCvabbSKbUwTshZGbvTBnAbcvxKB1ddhXMLc9Rhz09x5isSjuOefPQauthzYQ
+b16ZK/kI6iHLrCe9zhOPK2FSLtZIWcbfRKpmOPERILKodEheqTlGcVgYQrEFzE6
YVxjDwhfODccdxNPp9BDN7v4CaqnIdcpIz20Ql7SiCFjPcu5FC1U5L+AbDXoeREW
H91dFZtDuoRUGCUmB9DkjbgfJxXnUbB1MXhcQ+vMT9BPmwShe19G1HZeuCrp4xan
ZYqPrae9K2H2jzmYd4LYCHg6FoUcIkwC2bwgwudlH8CGe1HBeqbBZ4rD72LMY5ki
/Z7ncwuI7cFP+m04ePMuz4Gah8ukuWD/yHRK3U9zQRY5WddUF2VAnDItcRfHecYO
1B7zMhOuWoyIypY4Kjq/Oa3n2M5VsgiOprPLkTlxIOog4/+ZpMAFqx43zcH+StXs
h+aNo2ws/wDezgBR+XnvEc+Ijx23QRJ18+UUYcWujXpb9f1KEPTbYYhNnyHxt8bj
jgQJu0KDSUBBp9NPPf9fcvDFVAg9xiHgBIQWcg5aGHh2Uq/6H8NSx9Tb/aI+ObN0
MwUHcxs1j0NuTZyy/pkxj7lcbLVgmJzZG5EOVRJZeUiBQ/ew7P8SCm6T0r7OkOK3
C2naPa7o6k2qfyqgWTrcxwDYUw0SfGvsB7ZJeX0oXZsF8YUb9H17qsOPNQbNocak
KikarMYEX+cPMcL6eJvKms4kLSLJ97zAjN2lCjODNLptAig2WYtDg/Sn1UB1GuKZ
oq9LR8eKPrx/EnV33/zzeYGPKcIrQFmKFCsYXjCJwq/1umZdiW/RyzO5dSNCxxxT
smjJRPXdhF7AhErJLGmAdYT7YteCv1h/sweRRB1EFvIxJj+BXbUrvub5a1cvI9qj
0UlCdmfFASvztSeNSv2KidHNF8xfcRpI9rb5h3ZMyiNiWw3X6fp20HdDH5Nk2aTX
G7Ym8VNztO4tg6LEhRRtWs/VTFWyT/5o8Y7XCgaFIHw6VpHZUCoL9s9JTrdxcyzl
i5XTpIG71Y1uJJCE+qPWs7IV1z+nBd5HE2u27FIQ9CUgghHC/UPFFMg86/UcBsC0
Foyxh+zrLM1p67uKF07ayQyf+r7JefRXPi8dcyP+Emk/1hK/zvPt9aoFGg/q5E/1
GtCpcN5yEIRkKVqSn2mzx34wFnRA/L1nZpjRAl8YnM6qCgygmju0RvpDFAFOTgR8
pNksXl0RGiSc1GpQjOoUM/Ukt+PvyUMpLwM9pgXjN183cdyjXtohuOmIJkQO81l+
WqlxCWyhaljMVCCq+u1nfaF8g2VvsEwspYC995uxiWGsOJuV3NxdtNI8BjZ5LyTS
+vJ3xgtFnwuihDeOV3MLqRlv4Bd8DCnBX81B8rVy5Cvv2KYKLI8o+5qRSjrsfMj6
Hw6i7Z0A4GVcaMxzWmUV7c99BJ+fH3XWX8eYdmTiD31AwpZXc2nO64scEmy7INS9
GvhDd3+f7GMIRTCaDB/y7cyzKY5f8tcaxViDNtSb/JNEBS0o5aUEmBVtKciLq8wS
d8RPuJiiOuJJ5CY8GWWhpqsTS9tqe6bDvW5ZHROQaNht3OBm9G2uNtHc47dyk/3v
5ozh0lvjGJLNPNXr1cgNxHG3dS6w/Q3keosgsbK5yeH07UTG0oENxq4nU0+hDBbI
h5hjn4ykJchGO9gdEBtJt3PP33+Nsng8k5tnnfy0qwECDREVMMU6/dttar7Vj3nt
CSTIZdNcVPcZFeJFLnrxgV0m3SHtVyIs3A9iIrgsrswOpMUS2crZnVhoYMdwf9TP
psplaNjaza3k9CR0usCdtlQcdaXqkrWPPgPLczSnrF+iLdTMhC2XhnshwmvshO2N
si00W4k9O9/lMebb9nFPK+60aZDexK+Ow960U9KpqeWk4CJEvapZB/Zfi2MlQQQE
u+ZjFQTDFfp8czU+OAk4mD0II9acKnLgE0v0mhtyM2eShjkTLx3Wo4ZfzRmpe3y4
b8WtIYx7Ma5b/SmmGnoRk1WZ8jrCV36df4uHtb5WVB0XYQa1cKK52/mWhQnjdwor
YKsgSijtLGnDs295zAroP26YARtEUaV0xUtmX15quaFzIqiiMg4rpRThUegpROqy
gQ7OpIyKrC5dUtFSa/JWO7RYFtRpvYCh70//fplpi+q1YZzlBNSCZcRuZyBUuSBN
EF6kFHlrapvhZMtYGhyYQZgZ4fLA8ziNsCxs8vGaJ6OQhl61pcKOJkveRyuasqg3
x9vAmXVnLGSUV1DX8FAZAsT+XuqCdp1yXlljDXwq2FtJk/5v6rQbCvFcQqs+MknO
npM9qTA84sw6INKvIsxejHlSWMeXnA4Nxf6mBclUpGN9lwYKcFVWJrDcGD6NHkIq
sDqdV9qcA1khQKUEfuUwboIrCIzNqc0/+8oKu8tH/2eAC18pKngHt5wL9AcHRFVL
bLaKYdmOPNRnep0u0ZLgaWD6nT+7Y2Kn1zlWYRIhGP9XuStwKBgCHvyl9cHy3p6A
nGGQwACGyuSFLxqEN6bh9v+0jLwVae4OUqMc9cTVAqmz6iPrm7CWW0HmvE7axxnq
tfpQWeqWY8TsUTN95ADbkmPcRi/baJ547M41YpsTQwj1jyPV1tPufdnfV2Md+raN
+hFqMS1yBSJazHmK94NSkb4t7kgOaGkTslnrFJPSPkKWZ3ZQwDeLWAFONx6S2LgC
IETeTc4zXCX8XXnQk6OcchTLQt/oS3KCBSCT+nN2yDz/MRdmzxkBzV4F21OkfVG6
Q3v0pMA1dRpvEsk488DpOiuUUi0YISYbCZ+NdFdUooM1I1RN1BTgYf4350ikIAkw
8qMiHdqNgoUH/YKWzDBoLroFrz4xiJ+i+4dFJZ4gDUHv1Nf98fx7N6BD9PRVFb4y
+KtyPZtyQrtZgdLA1uDRD6CZnMWEOaUolmMbaCs2nrfvBwO6d9MpLdzAHDiQnWQt
k5qYjY28/EEhG6W1IMxzwEyr0ZpLHBtr/qUQcHjSkg0MHjFX//r4BTj8GyWgKFZc
4knB7CAhTPfd0VfNF4nJBXXyvGkbd2ocKP/WlpvREx5mn3F6wktP45JdFRb5Cc6A
ovfFFfbRqD+zy+PzIQS6WXWN8cfF9ZO3LP51+2N4kmG1MJDkQ7qI0sXgKAKoKdX9
IN15pdwP8OgK/taI902sGoJF3E8veudY67HYqZ7siV88aTgDbb08EatSLHuHKA4p
qwFpJdA5O9yjpljbJRYuLwY9S59DO5QV0ujZlB13Vw8jZpAAy6UasqucVpkyeA+y
t0uRMnSnZaFqrdgeb65sZ0fpmuhSzeKGLx0Fasg38RNXG20WfvNHt8OAA6+akyqP
9f5L8An6Ct6N0VkN3/lB4unOpTsV8hRICeb+5Pvf/BzbQQtGUaSlWRZqj9t07cCS
h4fmjpnEpTAluf90JY/z9EC+ZbvC3T2jERoHisugKcjNmTwSg+kN5B/Jqu9Qg3GG
C9X/wlZFa3P7D08A2tSoxfPB+FXeBPq61lazB1MJkj0Did72H7IdGP2CbIkbOZ35
ABaMN5Ccmf8U4OlliE9/CWqU+0ksg8JiMGARM7NdbVu4mc2+ma/+tezgTxnpMNMx
hcdEiznIbrAMshGNM0SBMpkf547/GYVZ5uH9x/Rh2BYCcBgoQ/0bfIoEgSsRTgxk
7A6VSA7A+/q38WrcJitbXfMej1LCx7Ao6dVJS2lR4Tvkm9w+sl8KI0XCJshP5bPj
qK3PKfyPcE1SwGntC1GE+oRZONWzgiHmiQy2emNqenMpS6+F05kXJ23EY2qaOCWZ
UN1GqCnK+M0kOvokOPe7yGhHY9+FkPRtzSLhvZyn29tik/8OvfCNPsUacPuY1bML
RCcjhsD+c2Pv8+OhmnUKQBI/Z2BlK1kMbC65+FSY5JliN39jMKN7GOt2e32dYKHh
fMfefcDhVXyGn+8CAxVz+cmbil0EfFWgLbo8MWKI4r4sq4wIC5msCI0O/y5uSi+W
Eit2sM/tdd11sU9Lv4+tEH7kOjXj5FXcPR+7lZJlWlmCyRpJGIppEVWeyQUgXVn+
U5ihR2kqpAWPinBZXu9h+/WJi5kLPSMs8eS29/037PqWbHU5O4cDyaGPuar4f2UN
kEMkvjs9oTQLvX9spZazm9kqgOGz0ijCzzDIS0dyLVR7SddRTVNAdnlYYbHB8eOb
2SBXXTAedKBd6FEkJPGwp3bo5SrLE4jqyRC5TkATHzAADLfEif2n5HN3l4emsYr6
YYPovXRrKDuSLSC/FWBZW7dB3XoZDCGqiWe0ehuQGH0gXUH7sQB0opdWjrEa5sQl
dT9XfDPSGpgQ2rSKTt1LEm/PxtmyWOqQ9hr55Ft8w5TSk9LKnTnMFt5/tclBulE3
2AIiH+MTTIsSvx/YMbtfCmTyA5b9QufL65Hl1GeP1KiNvPdZVkyl0+lg0iMfV14v
jMg58Ty5+t7zoyzJXtVbcq70LWfcs9ZbRq3lq7alosxodz1ApqcuyomNhJb9xZmi
b53nCrNsjyJ9Fm2E2EjknITEyLNcawt3GKe+0D8UoI/n7H2WGbGgsC9w7MqRVIvz
tc/e6x64rOWLQ5MC5b1XEzAeYZ/LMEe3tXwBnU1g8xOOzp43ZJ06MH+bkGfQQxtJ
5Ae0TxxNMw4fpW8w73qK5/TrbQY5ULeGm/UOeM54maFwOz2CeKP/YnLKwDyhnY4t
Af0SCUqYJ+X46k4lNzmcENdHlyOGPp4GfuEL9a2vhGJtdbABvBVxlfHFRqabkFcz
Dvyzlk3dHkbQVNPac2lceFmkjiRVrbV7w0sWUjiCL9Zw919alorrRzjUWNCJujVn
6Lq/ZNQEmettcFlkpHCLHkBQrygk6Dos09waTkrZd2oPgIn2TjBueqrlLd1/RwXH
ErJDYXZn4Rsp0sm9Qn7f8UzcgF8KfM4uiauW8F2otF2u/+DVrJHvUnSUpLkkwLtE
OmUBLQJiKvhJ0d5Oy/fDH/AA4bDFJqWDDBp2u0Y6pwmBuWWgxWtMUGrA5ayRMbx+
ZuilR2DW91RT3yTOVjieTRDxDjKEYf4DYNZRVtrGwb6cUA8UDSKvTDlAf1uN7x/n
sBf62cdagK6FTcMnnAmWgR9CScV9SvmjTY6vjLp0e5YV3MhdaFEUQZYn2mGX1Yws
9I5hInWGTZz6tFGS2+3j3YV+bLrxEl3e4AMBLgeqLUPYfnyAj1xgWrP2Idj4XOQN
/t3P+ZEmHGxzz5gLzL4pjv1ogCy1c88SOmAjgV0zlGqfZhrrLPqTnPNrJ+ActylV
GjZiEVNXNELNDL+QJN0ZRnuFRQd2CRrFGAFC4u8Sdu/Rvmn9q/6KT4hBFZpSkyya
31FcAWPWAzKxpdVjgQfYgsONP+NmA2OSNYzFxR1RQ1WeDwhx8yVC9q7pGDNdKw5C
EcZd4NB1UnFnuQtCqfNaP6M6Jrdxy5LY0tbtQMY+IxhEy2M8BJw9rPDryyAoUZOx
Q9Hg3vo1LY/iqbQ22sEcdw4wy7MBnUeSABojZ8VJBTczPCKYvorPscfpst3mSd8v
wpdG/eTjACPZrYacKrZy/tKyuY3c63tDI35iHlQjDbQOLOEy9q5mARpPApqwSvwq
d/51Y17gZGGQNp/PC8SXCZyXXIkUbgsmdtd6nsmA7hG4oBMr2ndE74O9cBeDTZ3h
oCvaaRBBTKMkgQR2glWtTxENdzDLx0a27YymPH48YTRN87Q9rwnE8JcUgrH8Zuo6
exh/XqPUZeKUOHe0xUnB09lJtr0fIuvJ0bYD1iCEhFALTsz9Yd/Ldcfv/gvS8ALJ
2EYapYZnSDRxvLOSIWnjtw3dWs3t2zV8fCuh9TMZ6pu/++cJ1C3bOfK3FLOzd3jL
IM+oLJvdV33vxOKnWszo3jFM/MCuFVFShbzFqbCpu8etCUUgSAcdh2UGfv9vFo8e
yTQ5wGFNybUu41oyM2dhtDotEIaUeegkpgYiEXnCY1Qa4pwzduF8tHR9AXZlWDFq
g/mBT68mAVwkUsUoYIif6kP/RwEVO8B5SN9L9PjAoXmZOAl4A0vwFcIdsCtxqwQ1
4hgf60M5lKsqHrOPJA548YB9FDQ0tGbPl/Z+Lhm5EVjCPVhNQKT9H0KyGGQd2vtE
kcg2Emoiqf+/AtERGgqS/37fz5vswmi1WDn+f2S6SIf0W2Bthi03OnO8huc/ehwQ
tV1ddOZZtn6LuomWUC65FceLXZyzLTJBWTWcz0i9MMr6GCC5WJPZiN9nI6tiWZR0
xeWc+YfJg89c9AA1PFngoHhTdWaD7HzJY+nHxbekuNDhyP+q3Bbti2ON4va4dWvj
NOH4DCDsNi5qBvYl2nrkUD3cXjt1JdIf4S3R17Gxah/hypqHfgVt8renRyPs1psB
6bCWF10u8EiJvkPeySuztDWAZF2/gB9wNVZYbPUxGt9PXucn767capB5AH8y5XwY
0qkiDxqG16agBc10l01yWyxcx7zWMU6uMIfDfsbDfmsRrpuM7qOx4c2FvozchLDt
WH4pqaqujfgl6qhnjpocV8LgPpqdwgqLZsplnIK5GeUsaFhfPbR86THRk4ZG6b1r
kgwWfxR0cWj8oI3ZQ5bXpyUBXGLWkJm3t7D2HGpR78wwXEGdUmdhBAGeYMngEQqo
aiC0iNblK3+AkVV9ay78MvBj1FKpYIwgnBNB6mfPTGzB69Z89wKuey57bnlKNoXd
KOMmnz5wYAO0CPQITxFDHKr4bRB5oEUg05UKe6wvpHdasxFslWRi0p/gEGCbg1iD
dVFLFodQj6nd1Y9AvunVxQFZJYZfmdCVdCEuvVuOE25fLEVYdqfe+quyZ9Ic/gIl
wOoFD5OXdIhK72eUQfYIDDX5B5KCnfHRWBbL+g8TyH2w+Bevfzn+bIMUBYBAM418
Vfsot38kTrzNXRQWGvCPvh7P8Omed/QEKxtxgtZsqQLseaxRAlSviGOnOpYiM0Zp
SKYr/LWw22EfSmIfIY7M+O1YPyO578QVka5jXBnAdZ0kfT5iJPPwEtaePMpumk3C
Uhj69BNyVOkSKXLSzrArL/+silAv+FXNYbyxOxZLSZEKa3eSL2ikS+SSQUImqNj9
EO3M+TX9geyA1Qm1MUWC1bq+S0EROrWKH54YQXFumA2EmbCcsMMEUR2ikS+B5phx
hJfCnU0O/Zfu1WdfmbJarhcLHfcIcQxnbCVVXPCWIInonc7Ip8Y/eaqcgBQj/Xcc
VpKH2uEUQDoOxLacD33XT/vayFAtrSKQDdcxqytR7Xpr1uFOfrG0RNmr3i71FAo1
DG4AcguW3pbXxK0X8klc9ru3HgXRzBwvjuDvpoogF1SoAYVGD2a5yorCV68kvtFb
X4h9dCuk1AC5vNShyq38RfCMPxrmZ6urUgsmY5OjPIW5WaY0+CUbSErBwHloQDxn
riZf29cJp20t9DI5t9lzOKtzMy0sgjY1ICCiVDZ6rj+hUzoMQj8qMOug6aPGxpMk
1sute0F7u/G4+zkLq6Y8vnm497t4S/8rzgboDCj+NEmKjFDdZGUwcluSsYQt1/lo
TM0VB3i/nET2XRLvftSpFKn9EQC6zA2fxYpNU6F5mub1xm7SYkGKslwgJUEAXurd
K6jn80Rhdnqh/Zy1ZBNtzarN8ap8aoqwx/JOnE5X5MUNjqmKxYh/zHsQ7h9dNMG8
NKL9N4x+Zyu0v9dIaoTiOcSGbpvhjpjxX+znmQKyAyG6rpHpCXvRTNlFJng5Wyrb
qPngBAevy2KGAeSydzPr+SRT6X7P3L6tWA74Y5raj3XQgMCwke0+gwE1xkph7c/p
Zmwr/LtJRbyoCaaOIS4l84+l8vy5i7xV1BU1KBv0jqmyWH4yFsJse2TEjjvHEt0q
E54xB0jcVrznXaPXYhmNmjANFI1mYsFEOirFbYnw6JrJ4L0G1sMdsZlR+Rb0rrgD
sGbGMwvObYurdBgUfaQREt2D9yajdbYPhgOdqsEEB2Xt98UuniuKVn7WLCJlYuBU
tHp7FGmSQNRAUtgxYMT0yI7CatbBaFx2ZP/nV08O0tj+8ImqMSr/rbIPJsXG/G2K
J7cdythYM6LTfTt4mBvj3O5wqFHWD71y9RkTUXtr+dZpysXcE3Jh0RPudl5c4PsV
Zr3JXp2h59zzmRrLDgO1AFwidd/pFoHuRPuqF4GS2XlvKoRwSPBy9cX5NmqRJrj4
CmyhSQPjFpdYMe4iX+kZJPPgjxLFasIS3kEq+LoxAT3Ho/dPOvAzmCsrDUfeeNgC
4y3BTl4UgpuXQ7rnu+a7p1ARPpydd3TltbDsU7XPujPX3NWbhQwRq+5qDVwF4jKA
e97knQFDvE3lRFFAfRfesRLLe5VvTxVy1+TlSfJ+/gyt5pM3mf78yRplxZWBgIYK
+WXxL8tDU1x4S1F3MXzwsmoXTHSpKIE0YiKw74KKrdQCIwYrbhJSIkp7QgMzs/iq
qjy5PcmaIvitlxLTJyDH9lIRspgZUqAhG1elhFTeQrVjXZm6+agWPG4xVysNYCtg
C69QwS/z4Wq7BtvvUyjQKBq/Ajfh5aIEy7JINHW2w2w30ArUaGEBCXnbMXLWCfgt
8U6mPPcdIPILD9tf0j33zqC1zlF1TN/trBedgUZ6osy5ks+aSqWkTeDJjDgUuTED
YPu4BWbVeQimcIMPl1U2ceLoLODBDQONU+468dWPPAAhC6VqMsw/Xs4rvl73HsNv
cLPHsisIzl5S4TwQJlxxoy0Fr5bcKBAblXsTaZBtpP/HGIcF9fKRc/+HC+REqL3U
VtFV9UwYf8pNBdnHZXGRv3Kbt3CJZNjxuC3it8cPO+jWbFQ+ZaAXfTXfdLzT1t7b
NqwV7y+ocqP6rm7lqsaoT5Dp2ZHs1vnX+jFAOZKCt/jiqLz1UMJ7o3a7Z9KOE07l
XZz+E6LcxPBWtBZcbMXDruoZJpfW0zO5L5LnJLX6DRmPAelsAQun2A1FtJBPtFDR
S3JThNSFrXcex/nFcCV5JpDUHiLaQoz8J5ebzNTrBN+Uh0LVhC0ZhGZbquKO4GT6
YLC8BUacZivKElBaJtMUbfu4Wl7XoXDIBX1nEW7DAoltwCyTmQiq5P8CB14crUfF
Quts+Ko78kTFG+qIBeaj7I1nT1GME0o2LEUWHOfcEjb1jwp7Ao5jmiv51ujnHBvT
PfKXppWBTvZY/bpkSxY5lPQxKrin8Zwc+kpwSUm0/W0R0HU0xE+7mPuEDRUL2dj4
lm3Frq5qIuBwiEvrLjK5gUL6CfZDI6rAmUTIYOuaInts4Oo1BrGW1HoOrPNfKAHl
WYP0iMEjgGgZsUztb4C06Ttia605jp/UPfSzVK3Ra30DiyRE7TlGqHOERxMipi2w
7PTN/NyHzYLNnHDXhQFVYWnBXEAUSrXjtu9bWeDEHbRx6SWJwrFRtuwQM9byZ/v2
5DG/EL7dUk42SGCtuwPVmm9TnrdX1gC61SEVTwp24V552vZELMTpMoka5ghqgdML
XRh39ygK23ZvBsq6ppeucy1LNhcajczdxcTc6PAVRjIBWkLaDPLtuBgfbsXh2NdX
2Kx5LtMmVq/sUaYBUcHzpMvXASrEGa48MviMbIpFTXchxeiogNVrDEXywTOqRv4o
3FEJonE6/ABVxLU1+FHopojxl2vwYDSV3rWZ1YcSk7fDO9/AWX6cesqC5+HdZCNl
auzc0MgzoibJd42U57rw57Io9XCj7dKKdFoQSi5HJ4ADCO8Qrw95mk760FY/SQeD
TzUr7XkLzonUmhh2/e03hilqwcUctTw6Kom8COeQ28rjBQzsMs7VGkmZ/jbgK1lj
d+i3GdoHhvK+NCGmWZDhCHYVD9s5DKSUasb20/IpWmAvgTsGL82zIHYnSA2SdX/O
beWtZ17fUmcOv084xMo1wQB/arHSrpJy/GS8d6lfmS0NJZfvwOYgYwxTntCPSFbt
Jpbajio3e5yKLb+/FnrWN6Mu1lEjmLI7oeB+OysiaxxniEKPnHQqnXRJDZCi8Ya2
y0+hihX/wE8T00mP8PdNk9F+ePOCv4y88ubiFLF2sH7FpnSBG5QNSvJ4ZWpVWQHP
I9T5Q9ILdqKhoa0nR3+rgdzTYkD2ZN+sz/bmFQb+dHuFDAhqHcJCSBt29pOE7hB5
fR/1hYSZiqvXENLrlRagU156OaWr07S4OHN8IGULiudIN3niLynKNORTyPU++OaL
kT0TaeIgHivlL3T8/tZW0zI7i7owy1wLAjbZkNSW4+OIt8l6VDU6/I8wQ71bzdns
rwxkOLjtebC8AhDbqZPeeqQPqc6CGO/HDIfQbugaTHVB2iUoAMoQRrINwJqW5wmk
VWlanSN9sEuxSE+FIvdek568CC/uyguMZAplsEp4ujhjOsc6PY2xhpxMVnuQDjXh
+WpusLWbzBj+3H51S8/OeboW8oGd2GoESHWsJieCvQRxwLZJMbtSt2gQei87gSut
uwa9+XaimRsOnD1G5LHlm4e0E5dxfQai8nvvHPnOSyphS8guovhL82rf7a+An1UP
/49cAHpSSzpDAYV8yo1fxqZy5lz5Sa65g2SkIc5aOJIFXF+y/mxKBFTM+RYvbtK5
SdtSMjwkeDFqsaCyIL+6FJYnrNCyGeaSojEX1POc89ICpuPUFVgEO9wHEqb717Ob
pKdygTEPvq39GwJHRIyORlYfEdskUvrh+vLqHH0/hjS16vO7INdNJxYCG65JsybT
+YpoyZRrlQOQRnClRiqmjOOtxvT56TCwvzsLL1Dwd2UcVb51fdHnzFBui7/u8xoY
Wh5pmYKiG6wEDLeKPxyX1rk/a4UWZRWHSxdHxt2RecubT9PMxX0ipdUdGte8qF3Q
NuxfgDVV29XVqiF7ipOvBZG6f7tncv/RwMXgY6qXnsFIc7+qCWYQoBFCFFfGeHIO
a/T7v2VbrKPlM0VHy4MeSulnVt16v6MlHWyfuwr6ofBOhnhAyKtNHPHm+JssYJvh
+2jtqoOXgYlyJ5HI0gfV2Io7cswrJ1xN/kpq7xv4y1L3AKR7pUR2Ufs6vCeOBA8q
dtPS0UPMPLDhp/qJtbZa8HPmzMbl2hKk0ZZvmUeEfA87/8wfI7Oho/QRtGx9lwqs
Tfz8m3g7CukzyWcduxLMreeclkajpMqw9qX17/iYzn+BV2xbbZ1IT7Ipry3jkdUe
/0uJkSpx4K4iCPZxwC0R/ynmuQZxDOzE9vx/GPn7WGnFJGQhKI3/sPRY/0uVQap2
/CZuZM7M2rQb3933MECVXj4l4I23iZiBrdUsCv4YB27povt7gXpeXOHAEr14LIeo
M/fu6rhtG0AMLAZX+L+seW14dVxOOrhnmEYZDBt485AUOcN5hZ2sG1GU5sFYuQ5V
mjEjn/pVHy+Ju+vw9EypvkkaVg4qTKzOgcOfureoIUU20GSIhAH2NcIE8UQJCigT
B678NCDgwOYCGE+jZ8KE7QYyZdbL8pIat4Y/KnmEGJmztVP2ruR2DvVCm8llS4KH
d6oJ2dJEZspY5tu8d9hbPtS40+vkCDNXtAIn+wMIwofYAuFmk3b4OQDP43TzF5y8
DYnsIcS7aqE/Suvan598lQDF0DXtRtZGbZCggtim0GMlYbD+W3eMBBzMSoVmDZOQ
W6+bIIFi2O+PK+y8spRtVchfp69PgSmcep96tafUnyELiA9KsnxB2PWzEQaDuX0M
RGa1YTxjhIeAJzpSvcBKu96XvNlmW7j1Qexy3sDCLTXKg8ztCdCq5lwyiv8UPcYS
6PQv/9FRp7SxhmtSpyMeCazKc0NcQEQot6yAGMCAwN4EJ7H7hUR4bcWB6g6nvkJt
DDARQqbFgVFhnNphgYM0uFI9OcmVALlz/GtQOqAQbKokLvxBUU1rKmgFHSIbEpP/
EoTUq528gjIMPGjy/MDpK+GvUKeuNQjSgqpoxklWYK8h0KVaJp/enyagqLM1s+jb
WQZhBDC8Lw/1dc20VCkxHG3dwb4GonurJT6zBTtJ1e1rlS49VM6fjNEwpBlqnlZg
dSR4l2W4R4IZua6PbXXR9IcL/H0CF/1ifbc6OqcLobEmg8riXtj9sKw2yPwLfO2Q
cPT6tAMQTMCfHbtUK3gqTaqmouN0NlmGElNpb0bfEO1bjDN4gxLmcJeewU6aaG7R
GqJF4vrCKOrrzOnln/cHpjsNmeGhIIM5ZsGYs41aIyWfa499/0UcmWf83JlZXX4V
vsv7ItK6PpTfL+461Nv00VaNgJaB6WlyaG/ktmniSqzhosWtc/rNWdqRGo/9XZgi
uAHr98P4YqhuX2kRAyWx3G0QSAlBsjS8wx6iGqcLVo3giPWqzRIaV7F1xJ8YJJBp
LGhPoZpQDXJSs8V49ZOUxcejiGTBS2AC2ZN3kbyX3SDYxKNUIPmwGGsgEeZW1TGO
ucdLd2DQGQ8yVofkO6ciOl2BmPOmVkettAeCR6r9D4f+hUmZVgXJPgtzDCxklajz
WMf1Kue3F4MBSEXbpnylY0p5F7ZCQvVx2iBIZ7IXpZO0LRxsxKDlmcMO1GN/Ji1M
ZOnD05Eb8sZ8iQs8VghCKgbngliUU6QYDcaNPWjxLaEE5fzalSY1ZMy1nSm/0zuu
d2eBlUMVCfE718Bh49Iq7XwVggxPOgEmP407d0exSgbodFAbSKVT8ct77BSIa1Sy
G8UdQtn4dvEGhfHztDlqd+owzmQIdS6j4v/v1YWivpbaq31e/EXo2W7UTo7BWtb+
JyWSy5DeCBkRwdpfMarvESJZ6s1HB6Qfe3mjivO8aQKK4rWq4ZLBbnz4d3/QHsna
9OorIsM4BpTH2iLgsDVlEAuWBTORUPUumplP9+a6+LllQtIOJFwj3TLDXcJCJjL4
rue3CMT7l0d6+r9wahrPdGY5DKMIlWqUzYWyKwuteBaCeLP94R69ofD0+Nv/sKtP
TYMERLo0SMAxutyEFdfv2hk8/stgaqfjxiNvljnTUMsGFqnBmJF++ekGeiK5Ysjf
eh5yckSkYh84ldUqeqzHMWZNUyP25waJlKlyxwK+cWXNbWA2o+ZEXt5PnnORIjEH
iqGp387BgKicVDnc517u/e68hWgDZwRNuj2NwUNQr4cxClbW2875jUjSFpgxh62p
xNpCsYOCAgZsCHkrKuFFhQLq99Wvk9iFq89g6faV3YD4RhwwFgrg4g9ymQN1s9hB
UR9yjw3ZhN/6lwywqHVIwCBH9thr9f0EzLBXHnBgGrNLc6IrB/cUe31L0RTBbJdv
ivZf4THelMMrqcnSSIxlgwELM8Fe1bXl2O2ErP210C8hke+l4dAv9Luprra+J4wl
tqcq5WdcXSh5y0MmgyK8XmFaLY88wMqkSFpxc8Pst0PSLmSyXWgjOYar8veV3iZT
5l+LrqNFpQdTvoCxDn3w+QRS2YdCgYj/hWfjzE3Yl1tkQMcKjroXQd8OHyO4Ibtc
IbKvYIHh0WKNeXhtfEoTmKVjpg374XXrh6QPN0M8/d5M7kYDJnNn1x9HB1g0BTXX
uBwU9L3c0T7aXda1ZVTVy362ZU2p4Lh4ZuJVoaIz1CdcKnb5B8pEhXeQvLu4c8uF
CIlxGa/EHbkQCjnXEnXDfDyAVV/6FENGlBnT8bNlnwtrhYCxGSfMuutRYsE/L2vu
b//weuaXHa+2x6Y0JNzJiF6otDG27vS+HOJpn2wEluAKs88Lf4wVpiOszdZk2Ryq
1WkTB0IOAC7837rLe1hAou8f3rsoY5L2P+700QAYQku91yNxnbaiSyhfjX2e5cjv
48R8FXYe3TAM84+mzu+xmSFu5Ppi7+KzM2C3FgmBI8vejJJyGkomxoPPec+Or6BG
hDTf308LvZnYczt5R0SCrYIQGeSY2FE8X+Wvarb8n8LdZLRDfptY4Hcj/1epavgP
0OOelKtqdIfV/PYU1vww3h+QNG1dwaHzPtB/i6l0yJk/qvPgL6u+pqYsQkG9TzQF
ibMOMqOYzOCna35bTSIE/HJUXgEWjiHtw3/aOteN4kRwfRYfffFp6orDf3uzK4Ut
HWMx34YPOBWwjg3PAX78SAd5+EOBepNsiTAoxZ5gOcDOxzom8TBMeGW3AI1d5/PG
FSCMJNkWQUjOvjaOOiwz/fMd4uLShneyk3PhEWI8XZ08cQy8FCHdGCgOUAz3TWBc
LeqsEAUGy3nGGKPxyQmEFSZ0EmxVCfg6MW1SJSv+EnhbLgy9mwaDX1FaofW6ZFhR
5CZPIH0rjVbdM52aQ3j+JLa/8vfj7qMk2YlE4NYYvn3xIBHCI4hBfHR6JuTT12wL
2jAVTyoURCPR5FE2bkfG/B//Y/DGQdT8IltS/pOSYEbYwYV2OTToBe3KZI8mQpif
zzrmMceW/mfFL+EwXAXmLopv9UxouegjJWEuUkmlWv50I3pvWI2SL3iA6+6wySlX
loW0d4b87ea5gtK9dO7fANe+AzKA2a9abbEMFcZKJvB21PH2P4Qtpbq2E6UjQzeR
gMcalaDmDzVwzWsfCF9VJr2CRwlEBaHUhsGaI9kmiFIGM4VtdqjSiOBrODTxY+zs
RjXIQKbu+Ikf4XTLYauUwbZ9S2ac9eLqUHKvTWdgi+pYdIpQNUQCNvpnrmKDKdF8
/4lSvSIoQlpWInyTbIf48jkgxbP9H5XWEvHRryplxEt7/unrVRrbV5DbLG6VQvHH
qLEwUtsoDZPh+HuzR1+ihh8xYUXM0VaS7lsWWT9YYamewhdpvSoR4pzs7+0UE9jO
SNvUP9vFMc9qsXFZV5GZJ25y4Bw+d7j04gyWuJytKhOOkSUgTkUgeRTb5DXAO7d4
SnpMc+DmNEte3mpG08YSxs+4poyOj3aY6vdwV550R93siJtNpeN9FIAetqRx27HI
NWfgTNDAiPMbuRI9wwX2+w5o98TltvjPRm7FwN0r4Kcj8Ck3R1GhQYVf4j5t33du
qZ3APAVhFmiyr9JPDQFzzTmfqhjr8Lh9auzsZ7n2WXu2Bcl9x/O92WyIkDFoJNP6
hWiZWvBQWKRzC+JWbgzLdC+1aUCTaCNTLrKus1BtolCIi0lyYa2rR91byLiOatm5
vOrAmhID3y2pBRqDCEW7Sq65ch0l8oTkc3edYe+kxtyW6Qpw0A6wJrw2Nz94tLQp
y3gMY0EdHg4LFtE/xst7OHeOt9FG4VFX6ugT/PLu5W0PoFGaLTAwc2Z7cXi3jZRh
XRp5x1LomdldddxJBG405jUe5Lpm6y8kfYKpo6fO4rky4NDXCLJNNpOPraNtRwnJ
2adB2305WYJrO9Y3a7rnykW30dLbSRmh9n01elTrObQcLYwnbve02kQ9sljjepar
hGe6rZfuJQeziaZlo4ppM8ozsuTCUX4HVLKF5Z6HIN9y1CsA5/jjsUof6yW6KqP7
x/yGWOYD6kSkHlhZ3oak0b4GBrFIBVdjUtIFd2WZtENjvJ0IVeWT+tsDNbeLmq4+
3lOdbSKAFGV9giIh7vJPnskNinQ027APic///gJXcnrd+1DmIbGe6ms5VYa9bdab
P1RIQN1qZ+j7L6G7TZFfn1bozA+zh/SWyRheSX7cxrcLgMcVsnhJAg8iwuSApgOG
tVjs816A6t5SOVCj7/61YWybZ1dDyqyRFvIOwhmKeSs7vUq+76Lj6CYUd7Rc2O2u
jIQDH0eZpN9gW+DScYYAiHkiyyrC1trZoizfy37GXpTHb33dT49F0fy9i/tXThvT
6me4LOmIJIKtrePjfVcc7zX7qYBSBthkgIRokubLYZiKdIBGt4mvOHw96QB61rdB
a35t9dRUlLxrAo/m9ZfytcKM0MiF/Hwv2L8rzXfUfvPaH+6kI872GlKy/th7MZKJ
KdKVMC+gg1IB2FKSGjNv5x2Y4IayCQnJ/b0eSFtAX47TRDvn0MMMdYQ6LB2WCrrw
vwJQK3MHInXwfQldT7eAfmIJAOPv6vnq+4COgZQeefMcci/vWL9SFA4GAZhmhESe
Dk+BUuwj7JlMofOFgevJh94HMy0aoq04VTMQDeknjGPZBR4Whsvc/FP3l+cWc8uE
bP6+YSNVy3I6r36ht/YFXpheKqC/zjnkWR0MtjZ6upOZRE3cAjeyvxMyfjcI6dDn
wmB7qWDFU4FK0bJ6GvBMYhBnd1xMvVZchP9bDhw9luoahf7VYJ29n0l5boiSVrI6
BcteJ1bguSViGS/be2Cy/7/adGgum7jb6RLhKYM5nZWFfvCaSvgBqlmKMm6ODnQd
UglZWGKJPJZ8bFYAZV7o5b8qUEb302FZ77mvMQ9p98thsghLp+C8jbwHa2QI4/ah
YojjurNZo3c/OI9v98N0Nq4nPRI5Buemun6IWBS7Sexirt8JCU1dSILXaq86gUQx
834ALb+HUPk7SKdFPxUN9TPti3ebyyP+qZIEjd2HyZ5JMs4SWNg6Fe/xc+PwB11d
cvn31SzENv6rKYRaiDcEH/qTTviWS3DXMc8nuGDzeWVWndToTFdJHm7oKpAoTom4
fy40PeNBDeT8TzyZCTS62p47H9sHseQv1uyBuO2vxN4jHV+csq120itPno5eIrKQ
mSQE7YC0OMK1gnuHDuTvleLQtPZjUSITDBTz2x+B3baU1oMMj9eDdxylYBb+7cZV
NvEZzIcm66No06xuZVazx+WO1sIqxeNbB3YMdY11HCvsgAWhPjD9R+FtnGKz39qW
NUDLbkMF5WiXiJjdsLhfDfBGzE+21vJ+mRaKurX85+OLDZ5P8Ozksqjiq1/PmZWH
cVjNpj3XtiAFqlwWMUsNbdimtwn8DEwjwoPEKR6j40wB31kvfVatgdLtJtv7DKrq
IB1gs5Q0/l/cofMwWB4/FgXxmGC2ihv5EP+9NgFqL/Cg96FtmrXst06Oo08AYBwH
BuYtjyzomqj/Q89LncZO4W1ZFFkd1V8gFww07Epu4s/Of/ZfVRRa31jw4HClyTDM
mhKEuI2kyPuvPlzaj0JlZ56EO26C4mwywGpJhN0Oa/b2do0/4Km2lRnTNIxzwBqU
FqKbihLvb/yTTFcAgAI/QNyWg/xK7HSrEGwA6JpFOaLcduDKMqADF5AWM+88AyJt
mJHkXxm/lVI1bjEgKTRlxhq9+lKCfwNVojKCsTkSsye6LuVmWpP6YUBwiRRKrBSi
ZdaCLBquVsOgXdnkaU1ellGDb8CJuJ3CTE5FijukiZxwuVawYR8WyrcOqzhVK3Ba
pKiruAFaCh/IWFkBbo6cCXLqIT1IutOUVAKtSXIBXvONCf1TGSU3MhfWgJFbHDhj
bRFgf2Syg39VWqM5qt6x2ClUsr/M3tHeYKzcMjGhNTU2UtUCiCjRiuiGRs5Jv4DC
a8+HP5jiGyaS+oLOdvTHBNmA/XX9kHvIi1IRKPCin+uM4muGSC0iDOBASMgbWn1w
IyD4vG9c9jxc2WykPdjp2dPn0BO2SITntL4iG0dAR2dXJeHXV8d3OZbd1l8rPxvT
4qQmhMlFe0R73CSA0ijYECNyu9E2oafXEx9oDu16+p3urypp3hgCcAZxYmdS2ykI
mcVN/yMPsLyi7W1Zr1J/cegArjME5Zpfv8hpO0BYfa4j2cPUIJ+LYCoQmGMKtgpb
gsrdr0+inVd7ZDch0dxyJ4Bw/aJ7k8n/avvjG0IzOXl4wo3KItG8DJniEn62cF4C
mmE3LgMFrAKW9oqTRrVRmhZRfzdWrUMeGBrAC5uaOnC4R807rtndynjjfukyfWXy
s64Lc6u+wpcaVr0P5yOJgkjvymk7Q0i6eDfMz1eTahyxMTQkzwvsd71x/B5bdVeJ
MbU0Cv4WBaeWHsno0eSxpeAshkeo6dcM2vFEDn4TWJheb2+yXBbMEikjCi3jO0bv
OZKNftmvTwguBmLLdnfOTiwj/ovUqttJoJOmRCpHrkF5laxCIpSEqbIXQjNhC4Rw
bwxmYvQSazOid/pYbYl+4ciLkasQ1IDt3cKEgJpwUVE1TYg4IcLYNZ1pnGZaPMBz
mfjbMtymxfwS6a6fVo3EI/WPWaSTkgb7qruCMaaAxbpCRyC0zaYey7C9EPRlv6o0
mf+37YJa/jBvdBd+4ENXIO+vPmWDbrKfdJtk8XVQrBe9EzCTW1v55MDHoo1P8pqz
J1sk26iWrfSPb+vr2Oh7E81EuyepdqxcZvyEyOmfJVj/YbPWaK5oeRmKQ9DCR7uJ
JqMqkrIwRDibGRzgIhehq2fdzPOjUzkFhtH7oj0ISQZD30yzyK3OBl9vvqz2/rc/
V0yxP+YgEjw3FG2WfMDjW5CDBiHnPR2tSFEaoOc8b+hRtJ/VYodfU7rItD+E0TQh
OAqc7lxgre2wpo8icwoxvi82I8KXDsySneQCfUfqdlm3fsocDJJir3dtz43IR/gX
J4QF9GtHXqfCSluB2MGSM4cjen8NhXOnVPfZ0au7vcygv+sgBnoH6RhdqRh0INP2
optEVWDdY204KoSy6OLfS4Ju4zx4TTyOAn22PHQIVmIBLStxcUEGuF7YSxi7Iu8L
i05leJnuXJoI+Xt1TWRmpp1UEcZyCYUOKIBEJKmzkN99jjYkmCo+MtljIlhgz7rX
YcSXCtoWIAkGukQg1PtTd0EZpeY4eObIHv5w498h2k10qL0X5SZPQ6etlGPf07Z3
d25dLogu8OFWJY0ZJWcKfvSPf0BcVugAkpNvWkCCiZNDy3iC87FL9QW4tUS3EpPk
nfRj5Z3aTDfInvuv509UdRX8MX20hmUEV3TJyhTqmFLiJ1+IL3iErJcMN3mh+ksf
n7Jpp0pBiJuLyXWE8mZBSolPG1PBKxKlzc6K7Ji0mTtgDceiyHQDPqmuL8Cjf+Ge
ysRpLjs0/e15hDiXQhcfjBx7PNKJ4VzTgZrblJxlD5epLtO+su5VNxrfl7J98/pK
w+XIj89JeXp+0k+4u3ngrHDz/iFBqLgfnxH2iKy2OxKGI7I6wSAUKmjAgYNWe4LR
GpDpepVeUpsoBbs6AAvDrqdYoAcsSvi/tDm0OBr5a8/yNl4vJPYgEDbJC2R2Qj5v
RwIDJbniXPL1S3azfzBzcow5xIUSa6Blw2iW81MEf5fXeijuA7cpF1GiD55tKGeh
xo0KXJ6pOZkbC6x1iRnZMuJuZLRccA1SjeyUibA3heaDndLLnC6Irb7zDJ1sE46o
KPerZ1wZo28Qw+nbkk1YqBr+IugHVWfCkhk27YYp9O7s4aQCqidZSSkjstC8Ay2X
nd14oU98oUtVkNE3ZmnekxuKSsDhSIbFNUCk73IMF0MbUMp1m0McsyBqVrWX/syE
3+QOjaKP1qJ5SRW1EMh1+zzkg1Z6nnxtFPz1Yo47nJGGEmOFWYKp0iQy2LnAPJgc
wpk2PZlonbQlPz8BV7sZpJSGyOGfWyrtwnQxDnlrULUlnSwALsFdz6AoatYkFdX3
OZOQq2lJknSW08wvgonyNqzoyNQQaeBT0Amo/Wf46aSSpUdBkgdrbBvpC4PYoHkT
1Z/cR55RrhAg08Q+oHjNOV2VTQCOMRYOqDGbvu3WrOgWiW92u6wCRQikIxfWyGRP
q3tFl24jutnoKDhr851PM4jrOOh1K9r1hUIPr+1gJ1HF9Jn+11mH+s01AsytY/RP
UMVsDTVAxaumGkUHADJMNdCIgNlR+XlCp2XMam/dk6lsh4++R0piYTYSam0Zcjxz
56zQ3mRGrtYiX4nDor2Zi0/13LgvBPAJGzPk56vPG0Icqlav5DENFUVvLjEl4jSS
8c9Vr//rP0bO69F3bdURmgaGXhW86uP6gyq3NbBOYAR1LOm1aMUnIzggBvUtpWPW
k1F1cfYZDyQKkgPpLwCJ7WHqYw+fMCmraPVPrNrCTG/k8ycwh7ka7yxnECfygPdj
AmFPEEsMviICvBIOX25JL6O136D/TcgnwHQfBrYMvd1Iti0iOpL+tNvuiKiwQ9mm
ehq6+q/WAucxrmPTzDlfrwJxlZT4f2863KtRyWZeBD2n2B0feF+cb1xwA9Vgy4IR
75vkKnEUc/1P0hWH0K0bMv7DsScTM9lGYzEycqofErPzHkrF16dezxO5DoRajr1/
sLUtpUDicRyAGskNVafWeldTA1AmI13z8dJQtdGIYftfWp4y3zJUTh7zqiImEsUN
ZMY6JMMfHD66WedaM5OW8oKViV13rUeZjcUmARsSNqQ7sWay4B83pff21PeYwXYg
0MCECmf79Tq9ivcNZHLP8ZoLqfAYTn887mfLP/ci0TYNwHZ+ciZsdMBLkTNmTz8v
YwoyFiCpo3Onig6GMvyvHHIbgzUE2mNXI0LOiG5SAydOiVUVRxrLZoUACjT6Ht5H
GPsBs2fVJaLxrCM4b303OWxAkqdbYUhbG6yoI9eoj8c+UUqhr2Tbu4ia0/SZwF+L
Gsw1VWGaqM7kK3KR2uK6DEfy9kO5KaAQ7WMr6nj5coGU5PwbhT1zo277+VWmUu7p
Zp2SibUa5sDeXtzdBJ5xqTSH0uHyc0fPQKE+Tdw6Z2f8KD8dbovDDrcB5e3oNos0
GlyVGGeCrxMdlDURvtUcEACIt8JtD64wtyVquV5X/3VdbUcAQNJUlFRQNkjJcpSw
sYMRkLBjN5YIK2veb3C+loP/iFEagVg8XDvJmQwM+neBtgpsBUi6wwe1nf1LBjeU
cZS0S1csEofVN6ex9UY0E1YyBEHafevmR95IfEjXc8qvHEKmtGRSY0XyFIrECLer
49QONiyBO+dsHtr8RWwfVD+x81fF+6GKIqPGCxHrQSKBkP7FLKqKX4aXRN9DvihL
PlcdMp38EEFL6WrP7MrXwZvj8qxIadaEPWE0biJK8xM+dl58CHIw33ueVCG9XO3n
VwyhNRVHOLpYA3lMmgP05rwDebj1DbmsyNPdbc6v/sHjSQ7WN9F/62queJS1ZJ3w
0VjnrgLdz4xUkqHSSU5Tu2wI+2dmA5uMPM75GIll3lHHkSjoZ7K+QEvdBvd5lA6x
FzK+xpib+n7NHueMKS2AgSKFFV9bTJsbdLfU1mnk4kkC6M9jRUdF6Bd/pqL5Cs9N
iJ/p3gic+dSO6WAOh5kxrtn3RxaMTsptuo8Y6Qzmj+wIRs6MMMCnG8l0XnKCxD2r
M4YZAjlK1gglSLM0FEG6tc4tVLdyDTIZ0OzM2N+Ya5vLUuVwFJIjOx4RZgl/k5ZS
AmlTxhJnK4ULQqA6hcP+B5q7JpKyNVeyxGJWfhqv2HdEjEeVCf8X8wmKKfD0wmHO
U65XFwk2yXzCNE8VXCmpNmuOa6DJTZQfE7f0fhSXpvC3C+7erDV7sTGmiP9wiVoA
l4Rgy2b8I7CHSCM09jT75HLaT7PyvSvRlgQ/PkSLDEQsl8/toD+eqDBTqLXUqWOv
3tQqkcr0TRaXJDAr9kVvkhm2/MFVY/NPe76Dta7WB9Km66aR2loa9RFEgW+0ss1r
eYFKIRekfqR3n2XGX+YVnT/3bopobHgtlNjsJ8f2UsuiK5WWrECLaHqkBz4dE8r3
nHZwW1JUERDKnmyNu3+muwxJe5WeQP/12A+ZksaaXLeB9BsgRytm+beYTWLlpIlX
D64KMOim/erpUG5Ihk31I3A2Ag2EL6elt/skbWAFzX/jZA/RQ7pIAGbwsZz/1zSm
z1jAz5lfk0o0zaqp1iGrtQthqF6JU8yX3iSCYRXQwGwSXTaa0RtEw+tCNqGe8y88
BK9T/X+bC8zaGuTencu0ZLcm8AurdLQJetr9XYj3DmDlH5cDezC1dDg0jSYA5VFK
/mKfoSEr0XeP08Mi1kYgSOIJLQEQaBGyvivUI7DUVDnI/ET2SVO2wWA8tJ+Br4e7
saRimWH+a/sW4YxM3g8ds9/q7gCxjNGpjZ92sJX7ed0/n/X8UnIXggqr6QslE9yL
rxStfY9hDYnoILwpTuoYsnF5uaWujua6FR/sX7yyXoZ7NaHq/s8dxg+COe1DGwl1
z3duXIrBLwUOslOhgdK1lYFGuYnJYpb/33TnDYeYzSsF3TfT5bFIaxEdDNGoEFfF
qHnoWNGXEcMq4uoc+f+mfRRoT4X5vKlDJ6JeaFscHc1A4jtrrvJZryFMz6ZtXV/y
DZ1CIGKs8aAdCuSscVSY9AekH1EG4MaufB0F17O/vZp5vCT65GXEOxJe6NsZ5i6b
buk5yAeOoAe2u+OhlWI9VE2r3uJNNb1YIUTreHw2qb7EMtCgnpDfo/FFl1nybipC
J6eo2ahr6lrIFyfn0s8Y3o6vNU99XfSsfBkf2waMew9wh+/2FrQYgZ5suTLJ9LYa
f4fwxbCaIeLMid2wZqJsXqlh9yDoYuAfdGgBvZzKrec/+Y3xfUcpFbruv2QPpcaX
Jg1DuP2cEnBQpNlkyUqZ45QR4QAYMFRuRaPH0ux26YzPTBfb//cAGAZWrjfZSu0t
TUf41Upyj6Tfmed5wXR0iHgrOW01RQSjve5Q4XupchdFToJYdu66sjITe9LXpn2Q
xcDass8904GQsygRcR+m2htrN58FzUjpWdYGOH/dAEtH65+pCkS9iKaAWhf8Cct7
bzvxgoE4r3ql9AJ4aAkVbH8ndYaySqFVoI6wFLXYRgaX9kq41y1BrrTYoqM1kJUG
zJMGBsNFjZR0CSiz3BYU+PDE0qdfkkECGnH8LxZFlRM0l0mC64XU53yKa58KtF6f
h5OydfDpQLpHItXBdjoSKUyblXCQ8WzBXDm7PtZb2OkUrXcAZ7UDY1L7em3XMCLa
rnx4e6Dnd3ds4Ea9yWBGbdG3jw2bnUGY+u9JBuRrK9h4gL/74U8qmHwRYdn4Cm0Y
vRGFKK9pHDC564E/VXdBx7rD/KcpY4r+V4px9nIyweRvM+DGMM/+oZEtxbqtf6mJ
bCWIElSBK61IWvjadoMYBiWPklBHHjLKQSqiqnXAxMVatdwpWOBkBfyy4+1gORqQ
hZM6naR3v5WEknTVq/mgzilTc80e+lnAEetky60iGhSJnQ6vCzw9I395TH3PuhsJ
RQwwYfRsy5TzMBiwOTIS+Qx/AQu6EJ5i4MXsKGlw4gN2KcxsZ0Lgtm0Q9k3tqO3k
IwEXul8BYNREAyHahWWnmoi9/hiji2Fdyh0DDE+CZeFzFTslElL7qHZJ0MxmEhcA
PVs55VecYXXqP91FiyiKh6cpmmmMqLlLVJOmS/vzw9Rbzw7klozLpze9xVlhBGlV
QzKZ9ularh390FHMj6H9yrIfHQYhAg/mBHs8RS8Dh1NOQoDZHx8tzWrofQ6BLN5b
XOvP8aY6bxxdOa2gzKwksh50iSU9nqwQVoN71U/4nuonNfvlPDY0+mOHaUvkm+Cf
Q4SYkfPV4roKPKVa38UcUQcLaxLUuKJH6r7GRyscqKOMi3LKv3oKJZ2be+unphM3
5RetedurzSpBp+wNBbP4A528YCCwRd4js/c51qtO4x8ntH0y/GQ0qVHHL4cX9FJR
g/Nlt/EoDgDYJ0U9pd0BYIPBgfph6hMeS0OrVfvYYNkTVfVH+ICdVs31gweWlMFd
6Tj80aDxGktpjBU+e3CEAp3NKWmf1AyFFNIGt5QAW8LblZJ8/f8S3SW0xXEumCsw
cNDAAwAiCkD5HiohtCv5gKyb1sX/yeVZdjdbkWd296ZN7IrqFueuHom0yrSuvuFE
geUcQmHyBQ88kpusxjkhm+E5yYHZ2likQmAHZnXYaGKPJs9ciIpqM9B3rFpqN88/
DBOO8WOLNPrXQqAlnWgWoHrvQkii8CStfNeZsYh5DbxKIbQtPbiQJXz+fbdkVgeU
5GyXMfTjwj8Jd2IHAUOLpzXkhEwP2tppFVomYr/sAxJXFGvE1Npsd5SJ6QDjOZ0Y
nR2s3tqoik97Gmjp+Yv5peeoBhH0TH36KTIg1GgTUxZd6/gvAYPGn7E88bj+OR2X
DNwEa/BmmRGT0ZVGoSsOf/XT27l/1HuUdvpD8Mo5Hd4Q4XWksvz/C8M/4Z4WuhKe
3OX9nzyo090E9jOIwAyJFAbDlqwsNicisre2ZVboIzLDx3pek9hhRc9PiztL0l1r
ffRt7DJzjiO5QB3QdEihHsFfEkkoRPTQGrugKmrJohCLekh7dbp5gRO/S01YrtLF
mgPdI4WpcO/czykQIGKt25qNaXPVe0J5qgXY2KZFnQ0JzsFLcs8SV5zLvQpK0wU4
M/91+nIqo+wJF2qUFxu4TG/RB6TMQPMvtFjRXhla04J8jUCjwxJ/oretPVtNJJrF
qhaeRtwv5qTzA/pYtaJhK0Z/UoTb13u+zaWfx9vPwrmgsCi/b2J/RBHpgJMLZrM4
JPx0s/bKfvVz359XsZC3NJTwD6JvRDq8Vtgq3enuAM1lDU7AxnMmWovTNScS6SIW
6vmFDeunJdHDg1L8oDu2WHWmS6ubx4IZIV7MYdMVm1xmGj46A3H0vJVs3rFxu6bf
jBJrmy2sH7kn8ke0+ZVvnyhhdtAhCSjIIh+nWzBwycGhl3oFjqkmtXRc2ChBHP90
aGJbT1nIqNux6GTzJ4XvlaeIAOQHYx5pcC4N8kfdmLOCt5No3NkyfF2+JAe1jXyv
YWSPLldhNMd8B2JPvo4Os4sDcUQzsH0QU4E2OT9azNDZ1F6o/Gl8z2xt6NWE8OHT
zcCoPoqPCWxjUzWd5mdaS4G9ysPz1XWypjIAs/crH44bUyUhQYnQiB7sJ1iIVxoh
pEPucCYnHsfDbbBCnomrzY7FaGlTNje0FRvSl+x3YJ6FsidRvYN5WMPFJjFDqjqU
MtiG7Szvk17gSd2bU7RwtJRnVf6kzWIC4XafU+qdAo0eIDXXVC6EUWLbDrX08ig1
Nd1mR2783bfp8HBDRzxR6vyFn7GUwuyHfycpLoMvo2bdz2PFVzLuIMUeGKYTOoB7
gXo4mZVT/yQLuq9NtwrgoOj5BeNc4ffEolr+xqXrUzm6h5jxGoxB2zBpOhAFm1Sl
/NxzH4+i3Foc+5LISyLHjsXsmqMTmTgLQU/f9Kv24NrJUXszwW36bn02GOtCQTHn
7YvPvkrIJRqdREitJuqR1uzmSvRqRg6brHFL2aReXtt80+FcOn8s3p3mxy4atx6l
bbkFzE+Qb9kiy23ldUsfon4vbkkkhhRVIFjaLhGw5nRshbFbnAM89cjRptySKyNt
/ON2ahVhSuaAgjE+2o6M/BffYU2061/lgnRT8OMgWKl8CpyASxxz11h8iczLy5Jn
uwQ4WI9O+pAkyy8hlSi4TepXJflewCA67Sn9J28s/f4yu44qy1zQOBVnq8DPQgNC
a37wV1AptrNk0BeVQFJCf5WvIyxrW1Fp4O7H9/5oME1zj4ruyu3is4nmK93KKCcv
KOrwQymW93OkcEGUCNU6Ki3CYhjs5VYML046RNrWIxlPssTouaFp+RCOHXFu5HjX
H/misSiQATd5ca9N04EuxvbSGc55XTHW2ivEm9frZQWX8Xasip1OmH2hjOEXVJI4
lpmYLS8joT0FB8MnEKAb0m6kqLjVbmfEcOJMX8q00ImQqIQpKpnP6FiAsAx7YNIz
qbfFrmnHggOuCcso3Bp0TkuSwa+TqdLl2vxVwVY/5mjdLnGOjslHFAibw9e5BkuM
oiPHa3igONU/Z7nKKpZPsK3+GQzeNvX7xTMGehEOiSV/fAejuO+UtAAo3oPDPF6s
6wwKplFsqYZPU8UMP401TmsFfIiUwrNUvexWynlhnLZvUGVVcU/QJKvNcPoVr7uz
vjf3Uzo1PuZu6nr4fZz7IwfP2bPVFMxsenbBUMXdnTwT7JoyqfPwB2fxDjOH81tN
sPRRC8jiBwOAv3lEoT8g9q5+U3J5sZPfRMFZHKbP4WNb3Vdp1aV5FrpBOKYCPchh
Vo8xp/sZQxnKhhveyWePwfRjoc4BX4hYcXf7+u4MR4Si/dQh6ptAc2nuaG/SADmF
fWHKHKib6h1VGoJlGHtqjn5PhpIMSObqTbDpkIJOSoDmvEOKNIf7Hmrg5QnSwugk
Z+QKU0DpwkdlMKysGiyCHeCfHDPUYK1SryHYeWckRHMhiBXoE27jxKPSY7/zhdCA
g8FBFLKRn/M9o4zi9Knb5JiwYICsOJFVpGAwuV4glqpSwgjAmm5yroEg+ot6B5jb
x29lNL5dgILGMgczje1LF+gVY0jLSfUT0pnUmQfUKABkkDJwrFiprcFfEH1IG+Do
hmE0DbBRjHpB+xrFYWoF+O3usIK+jeT2SsxuEKIvRyosZPfbkqpXJvKnvZYTtkXV
p6a2OJZYcm3o4ff0U2IiY5l3tZluDWBokuBXpajr3eFD3c8cgUOFUEoWz10ulZVX
yx1kFXQcCZPfmWNShWf5RfO9A+OEatRGw9GEfwR0Elys8rXyBL2sp5T5CRwL9lN6
ZtPd3PSnz61BjUJiPairLmHhNs/no/AMHj+0P00qdly9Xh/oFTphbalkf+Xi0gNb
qs2QAYadl7Z1uYnKnLZOq+N8upVeoZr2qEfG47w5OrGvu71gYHJ9Mo2L2X8GWgWn
baGGQoC/9H2QuqF4BJvV78wcIKYeImrAYJYJl4N4aUXyLi6jItTtd4T+GGu1bkta
s0ZypTtIULtds7I7M1MrJ07qi5KJuptE77034AOhd8VRtU7n5QPHyv7KFtEnXWeD
TEsu9WOvGTCInWBnV622Po4XNF9akRIogZ9w2siD/k0fxKHOKZ4f51bas5e4GEuu
Ym3oXbjYCdom4LafuDVkq/ZWVS2F3L7oeEM5sUzGXchXDegysSXZUjOWbYrywST+
kHaJ95ga2D5+G865wkAgUjKJ96glhI7jQAbnUeLYLtnFKMqzg0suyKOHvsfSvVuW
DRoCzvumJUgtqnoqVjmC1gy5vp2qYz1PwzVC2763FuToB5Ku0iuf8kLUxfrOu62K
ZDK1qaZ3xedX7sIqY/bFgM5nCpID48IMRNg3ZW2RCza/rRgEgBEIWat7eNMqwM2S
lCgckNRMV6gb9Unymxf0TekYtecKYZ3D320y61eTVTeF0QQqITOnrVxQ9Fbq9oaT
cDUZlP3wNiCgr2oXF3AvKlVXlAKlzEa/5nJh65QLO5NVkwhWSQ3Bb9StWzApCnQF
RQ38g+6NyYeV13brj62UCecZst5diB7+giThmhl7zxoQZWwrC0UtRFIKexgg1g18
GkaahSiUdwFYYMSizrLC7l9LyuoKXqBpFBT9Xc2cguDQNYnzz2v35Xt33I30Jua/
7cifOkFEFw/P0tOx1KdnDjlbismHEPhiRhwhjPPoRqKGf0tyyidQW8ixvKa37GzD
8kVma40sT8a1AvL2nppomQEjZmkjKggO9wQkrJ13axHthyHrP7Ieos4CsBFu6H4u
8pKwMr0tkfqL2eJBApkD32+Qfpn8zHQLQi2Woq4VXtFS0FoKpk41skkx6lricIND
/mgF1bhNehrddDwUNLK+fRrPId1zt6Hu/gFPyXRYDFZ6iLSReAdW9KCdFZcG4ysO
wOfaCNovYwI8IB80T4wG47yXSC8M2KdF0RzCVDXJ5ox9wy7eCaw2l9HRzgRsMDHA
J9K4m4HdNpK/tYmXFOf1Etnu4GduyPkAkdXZa9dbc4aFuT68if8oqJGHWzDd8vGa
pFB50z0W/QPpUZCcGcFFdj89tcpehdUw/7y8JNUQCBa5Gl+tOv8erGprxsnEJGBh
6CKozf0fwN3IiP4anUeEKjcjFRb+VXx3vpKZaG3ZjBwkU0SmUmntTZUpuwjxr2os
08rYnaHXGRzJiLH4KKtcFoNv+rGhtNlD3RLVBKENT3pU3ywi7NCDTxw15J2Z/XJQ
z/nl3pjfl9TFY6LPudpCAgldf87yFKvkaK3TgTPVxR+LlqNHNOLvLRMjImENFKLS
YVX39yc9VMKki+qVgMaKYQfS21P0Lelth3kjg99X6i1vqyZIyo6KkHAZr/UHfkEm
lUJdKSVPWg0IMPlVX9SBUqWeIMAuZFZXqqSuLHThrcvVCfqFbn4IlGIK20fxqayz
3dGY75eyJrwZ1x4vUB5IF5Fvl21J6fPDJ9kdnVYmI62iLWECrW5RPfyHP+y1+I2c
J9yLY13ZxLSl2dhb4tugn4YXVCsCAMcFO/IsM38Gb6ZddVKrGOInha7hcU1o/6hM
+xucxpu0+6NNbY3/NWfOjlC2+uHqB45dzhDY/h/Bamt8iW/yMOgc78rvTxKZ1O9K
1GIPxEneNczSwrL/LD6W946TLZImb7HrWfmAzMS6IYHN3FJdZY1G1n/ug2YSoe/l
vS+rokz5AXnm2ZjDKWgSJ1srl6ymq89DYbqBs1Y7GqedK4gG3wzM8x2KcNkl+9LV
6k5eBPz4mhEegcVpANfFJkTJUide5SJIHkfVSOPACN1v2TJjcAVZNX52S2aPEWF2
dh42zffKZyKiSREj1pUv31p7gAOC/mCs6D5Cd5dXUvz2OIDc9AxUK8w+yYZFJfnR
iQ6w7hIQxAGiKSE5E4Zgc93rDRyd4GR5LsmcbbaWxUj/C1fKUWfVdUAdHiM2lPnu
aMtQ0eaNOXExhROvngeZBxb2oE8e+d6MO7H9deyGAd/TVhuOeTWqw+2SN+HsaCkX
yP1kILj4EqPfIUf7Yjke7PyVmjU05mXi5G4Yj9zIEvE/4Z1Y4QRxjg8kHh+BNlCn
s3ciqk6S/4jkn/Shq/C6FexWL/NtH0LV81daSicjtNBn+dcrRhGVak5hG15kHJs8
Dkr16Cd+wvwqFcQHF8mJieuR9ftCO9cE67cmQifBP4C/mwNG+ie/JZrxe2aqJR1d
ZGTjWdPIx3fin8Cp7kX1GYpo7fjCdjPCm/YEYRwELJJJ77FzBtPP/+32p3ZGHl/g
GoQiTzsMPLeAjZjDoMvonpOFHUbex1Iq1xuLufuVsBWc3lyK3C9ieLpiOIbV7cux
gi4vR1RGDVtAB6vEpBKyyPMCxPDToB/QzhLvRhVmECzBTlsMQdcUFt5tmHtRHBWx
5HsMSvENVJwN2PN2ce+cAz9qCsO3737pwiQxTWBcoCsVTWBPfwWqVbdGejo5bv1J
hvenwJhfJiIRWijAC+dFGsV7XP3EQmWcGtj6WUAv8TjKCmSOVYCJvjYOhjvYFUmq
QUH92kHLD5ccleqLGXu4V6Q790uWh/gquYPfpeT+71tiWNU/Yc1FvPU54w06z/rs
1ZFt0RrZEHYkVz3MuVN0/LAa1APvoIfFQwwRZM/JHNd8zVYtVKBDiyEqTgp8T61Y
1OXO9sp+X6XWRurUQ7SfrNwh0irKbfJD15R9aIAUksnC9uRRf1ey7hfMHw8kzbtB
3VVRdxS+1Z+dvEhGRqa/j/BiwZb3rzrUTIWp7w0/9ZsPQzZqMHMUPvEdvVccnXhP
vtiGY+16xbH9aMhXlZ7uC3G3HI1cD37dMHpvvWi8sfYJCqb/rU6EGGVkg3gwQ5i9
RTzvQ+KlYRlCmIeS0ptJuLadjHa46eN/gSbqYET0PaRLee4slUa06r03nmRZ6Xli
9hSck5hmb0M8A/acuC4r7be/UwDCedfdz1bJC1jiT3+296iv3BAMQT+KL7t9sFt+
19mYAg8mT3LAIRhanlrwShJLOmzf2EVas63sv6OPeFZFjq83LkR/2yw/1ZJsiXtM
FWwYOfbmiIyZK1ZIwO3FKb7R64n7f+bSM97HrmrULXPEtKOPbKW57bz1b0ejjbRE
CcZSqgABi2mTQgeDwxFBESXmT1BkoLpbiMphaab8IgJ1bQn0UM5AvoxkVeLo4Ru4
mMycGb5n3S6HcnNXmkKBvnofsmpJ8Eghv8WTYb/3A2PNhl8aCHHmO7gZJ1sRHpl2
lMM4qtd2ERWZG33Jt2I3omg9iRvhHNZbJftQ16FrJCBtUXNuzOG1Wv0mjyeaKaZ7
Pb7JD/n4f8QJhZCCDS8ebxIpn+US4Y1fWC2lc/vKxbnukL9t24KeN0WBtBHJlJ7Q
lgNK7IQKOstmyeHeK5APvHm23REE05EI8C0na7LMXoqs5Z78GXOsvkXF+VwaZxqi
pLJLRkYy4jUrc9LdbmzHTULZq/rWk4RYcoMRw5IFOnJiMfyjlQDnbs6Icad2E/3T
tq4Zy2e6t9TEADMSdFjNMYvaINm6JA58R//9RDxEWI4+vVIRgFKUwOde5ZoN2/+S
A21hZycfcWQvLTI74vu+Nerjo8CuXNZ0YvIzjWK+v7BZ9jixBcwgEM1afZi2z9A8
tn468KrT6vBSf+cIQPxA3RV0SXV0rdbNpq+ai/WM3XgF96VvKwi3kKeXGITpxIYk
tmus7w98dpMJG3M6jCUqN4WfELpErU4L3BTBBL39dk/F4ssVLxZ9rKXY3d/0QmB4
RUCfSQUFbOvyCzKec0Cd+quNsWu9OIompvUeCswQuvepkrhGZiC43JTOwvHqOp30
BF5MXGuylmAh3Y4Dn1jRzYm75xuniIZdybW1AulYmSC0ey2gq48wqp7RkZm6vynG
L0x2zPHEasUv0iEyUQao8SjhnbdVrKDWVg0hpSY+85wTmyfJLzxZOsCQgUPNFF6Z
78SDgJjjkSzTM5pabVzfHSe7+eRv+VdNahpCdjbdqKqkK9ZTXerMS6qj6LC4BiNs
PI1ThWMkXvhgmLAYwAZLVGgpLIocRy8PPi5x9thjwefs8ecXa7iQOVkidaufhFU8
sOf/yxRKNK3k9A9wrkPzKZm2Ws/wxzpUnIrRSU8mS8o7z1Br+LGtdngemnwBS7xI
CNZgqYMBYgjDq8lDaKwG3JgrYgW07btk+mi2oM1bDEBWuPR3fy9RIHqAMHnWEwE+
ur9yvAvbgfzrEZVmWK7sAAn6LjhxTZhhwQdQTddJu6tciLm7kBAMOlgf5//XEX3A
2/AF5+hN4Fcq44g6Sx212vqtkxUcVl5WpbxDY32lU0CUWUpLKJLVJ31hZJ9EkMvL
vffUkrESMFKMrjZXgyDemCKgpo21on8RoEJyh79UqqOVk6BOENcl0UnYNQ2/TLIq
lIrWs581tV67oG/PwRpTq2hP2bV+noysMdJp+ZtR8IJRog7vZ8eDUUq6Bfbo5lN6
f9zF9bVkksOjeWUuhju7yb0pI/aHJ5MhBappOJvTtiVNYyV+iPRY4nkf0USjhrH0
qNOF4rd0SgyWxfy6VWGm2lvOwA8T6dkhZ3y5uAjvH6eXuThC8T88tckR981dD5wk
EcJHTyQ7Pr7ezgnmj9QL25TzyBquicL9+mARkB3EXng64PimxhIHGRucOyyhREdk
GBhXcTGFv1FcDp5HYWkb+ArOVe27NqBHIoBx2nokGvf1+PWaxzSOmwmYg+WUNWZQ
SEE25hHyJkFLfDDFqSXk/bngEKgYE7p/9bMq9BmSSzSuFc8Cr4kkHNgU+DGWW9OX
3OIn/0cs3yxM5GLjoBMfJiSFyytm7a8BxS8pF46bcu7h6FH0lX21vg4lD6yJIITK
lGNl40MBG6YskqjOZL5g5/aeVQ1TxQiMQb8iPlIdNCWKtLqGmY0HE8fJu4f6zkMv
2tLK6Lul6mOVeJ4IVP4wXMFdkupT8bIMSczyiSXl4IdXu/pibwPFQw9QOKLLPuyb
9srkXYxuWWtDKvU/PlNHveMBQk+P4LTw6KjZbG8nr+NfVlDqhjxqGkmylWCwackw
RCHjCB4c0gQFVWXRHpYoydIFfv8h34RUM585jHo/gBo+11oU48wX1KC+g86dDOG6
UsNvda2KvZonk/eIuM/C0lWcDi8DAH7kFANihh8mEu+ltwsy4KuSRqc36FaOBLrU
9Va6BQiMBigPDnRLUD3UglpfaGej57rfEL+ffvnyGAbY7T6eXAryGDWbxeIpu57A
PtPkeNBJNaZfpSY7kslAO2Nq8vIVhcgok4/FqYnbWia5OhS9/gHmjIq7KFyTNhoO
gNOOcknfDsBKb1KzoBz8uDAGuF3wYZFB8V2g2tdPFkpkCvRgBqGX69qklRtDkmQS
YYJEDOk7U5SejtH/jLfcg5o4SzA+bDBZ1KpvMX3smas/9sgfpMDunOJANcMa24P5
RsAkkanJoNtdGlWvn3tT3opTw9ayB+/64535I8pYkv9FgnvVZinMZ47WBL/9Z/+J
jggbdPPwpmbqyE47UcAgy+6ryzx5J7MJ1XD9aGMFfZbkNzJ95rKt/Dx45Vo2LAXK
IiG8Dc9t72bEAAX4S4MLA/Ej0hsFI9sqc0T6eA1DjyQeLHuHWvH9rCWvOt9WDcg5
zdRxWqpQXaE+rOreBs8do9u8UpcLIvCAExWTJ5RbgCBQXmq4SHmms0plFke1bmgu
eFURR/aj8arPo0a/TBiun8rNY0YLSmpX4aXq8yyUtV2+CgUAs0rXwQ0ZbEe8Wm6w
C8vHwQioePsC/vk32UHEka0XWAbnSuu/dlNxn2vbAEYhWEcKlFcga11eFP0C86Ho
6xy9HI0IMnjaY1izBR4V+jC739oXyK4uTIqpUs5s4g9pCxzngxjzTuFGYv8c7iH7
X6P/FZTWfCBZetJrq/EzMdXooqELbWEw7nS8SBhiRJtG+cpnvQ+CTpQpjKbTTZdL
dksL0NDeBuW8j1LEdk8np8rIy1TgPnQTSDXWEg2nsyNawNqWtu8d0//Kc4uR2Fzu
eEM8pwyFrnRP2RVzkLRaFWVeA1fCvp67mU5J+RUbxT5t7JHieJnDVPKkWl2QKINO
6dIMMviAo+JXUSHHhtk3cgyskxbk7ayBMhZSShOcoNstntqwfN3p0XU9xd0rw3vN
10ociYnPsoCHr0KYt+GN3XQJR3E8ws4ryB0RzPG1JynmMOB6Oj+I5W62HdCeX2EL
4QU3VmwnyUGKe3pT8MCON6fZkneQYyYEF1/LeztbA5UdF8I1YLNg+CSCSrLR8aZI
cczocWaZOrfzAZLIPAx+byTHw7yFKfE9Iu3DplQEiw0qGqi4BOUXGUb1Sdlr0Vv6
LNpXI9QVsB43bLT42zhFrQljiyla7ksgXagWaoPFLgCt2cUXqy4c+sEE6rZqJ1Lt
qbtVV8jdp9oM1ZdyPsir40ShI6zbKwHhWMkf3VaD6o2yQ1FOuyGiEWUg/tGZQfS5
2JmKA+Jv5FtEWv6plQ1oDz0iGZcUTNkVj1dZ0HBvcyDwh3wtkI46CLI0GErdGzTW
sqGOCQf5KXDFt7DGMU6hIZ9mjQsiAtqwfZhasWoubIj/BA+Eqo5WEqo6Oa2lns2j
Ee6njjqNbCrkkGq3O1d62o1mmdQxhiF1j+08VCOFOaBJPl3QwiVojqcuuqneZsMu
3Rk8PoERfmBH4U4IKHjEIytwXXcefFeL/rnh9iO9deaPJavNNLUh7Uayn5xlFQQh
TUzDuLQs8TOaWZA77Q88HhOHniMmtyTP/B5EwQyktlVTlFeiQ/GkINbz1g56eLqW
POEJOiismq1ZdHP7V15J1ShZ804BmL2hfTiRXwBEaNpeDvtFoYXddrEyBrlMfT/Z
8OgChBM+wEJ6597dhxlZEcTHVXGzincmi4yEEONjbgu8SKLMb5S+3wL/vqrLvjDS
pBzqs2OGargpyLKyuiocadKr1ZXzuxsWk1bjbi0wgJxSN8BZX6eOuFHPeRcpVxLK
hD6swk/zymy/v7O/+KN/6ncIF0HKtPP1EeWA8H1uoV1X2kfMrdFiz/mxoGvE0Y+k
aLkjZ37IZ6ARpvx2uAscHFw+iUDW+0ZMdWcJJOFnIxN36OJSkPUGlHf2uqTHZPb6
EwcGmNTwD5ohKX4wTA5UkGE2+AbefnkK3nmKMEh4oJBsb+k9x8HxIUttonNp4rdH
Ae1Cs8gtEHKHDPPwW93vAFzIh/hEn2CFmCXtv5HNjCoM3IOEA5aBALLtKa4lNViM
P7fmJqW1DERwTTkaKhRGioLwMAqWZFc7xpn1jb9vNwIJt5d4+2cSLD13hpxFzaOI
HLLMTYTAj9Upp4C7VVRA0trSkCh9TKZTQT0yUwopv0PRzV4OC6BSpxvwy+gAT0mH
bru7TMDxEYKddVXx7j93Ky77wPHVMoMADqDtk9cQ2bOfEPe4FuQEHiBfeuLBllQc
8SEOVI/dN5O0wMJo6JL4WBrmKRedb7VHuxlN4rSyABaa/PbZ9UDxQOHDhdYN6Mym
aZlXee4wP6onJ+KUqcehnbVO36rZxhz8nuT8Og1cmbCNeZtY0wz6awuGNbBcbATA
gqoVqU5FRxiRf0Zibv9Nt8WxeIrRBgO3y18kLRb7H13PTK0cYScDzB1r1hSM2AyA
NchBtpfvV7vm5AphscnzwbY1+IvmpLrw5S9jVcwZoIMWtYMcmGkp6PpxcGcIArLH
cygUZR8oL7aUWUhOgcq6CW0a7T9eVKmGNVQZw7MBqS3/OYKRmPXeLWOkROxqYEDW
2jXEnyAZZS/nqYz9cLBRTc3k+4JOZdrZ3zsE/qLiK4P3LNuq7EsXGhYuNR0TNz4+
Ttk2gvKCeuxHRWnQ750Zs75XRVT627cE4Z+vK8VuSJtAhT0dylHwOhvMie34XaV9
wLtZOBDUSytVUyJk21wsX/p1MRAWZ/ePRynf6C2F1OIkI5Ublxh90Yb5yDLrhVMr
rIqHRrrI476/30MTxQkLs5q279ViQp5rtFZgTJzFN8/feIag/0/qvIo3HOwNw2K1
3s+0WgOtB66dS3VVCAZDNa8SC3j1szniqf8Gt3iipMwCG5Rb8B8eeF+/PlKLuN3/
i+I5JDF3ICoqsPxDyh+CTXDwZXgdlNfeZzJsO0msvuAvpZJS8amcZThq0aJqqls6
XTByjFdFFyvWbNFkt9lOrYDNeN3rpdcWr3DptnjA7lRBuVC458HrBr4NLz/LlMJt
NF5UN1+XSCciJrfTVSDbzlHl/OFT0KxGK4MLHyqXOnLestb1kBu3V1La3OCXaliH
33akp3rLcROz7Nt5ojgO22wa/Zir9pS9VfM1M5khkuusZ+8kWrKzVNI0oqVlb54S
UypBqeI7niKMJxPBxzxX8ND4ZlRg0EQXycIgPky+MEUDl4oSyKFU9fTg8r0V6hRd
n8o09NMmBd500LKCVe0JyNdMHT9BQgEQlwsA1ibTdjwb9xzXcs8tFLPKxCPvvUxo
Bl+7Mq11KQBeqQ6QCcMyFbvoMF99Ls1DOhvfFMhlmcI+fGW3X2Dq8MvorCTGs5O+
+x5UA0il35MFf1LSSf6OaXDgyOQAvHQicqrUaf7jvKO5M950+vV9Ug9xjMwn30ET
KJwahfmQ+c/xfmrXOo7sQQjzwEE0o21IcYGYdNDuxjUQeU5q8wZ1zvGxpU9jToDq
kPE/oq3mdXysNqpqMVGSNRWFrVOdU88AMpf+p09BWnCA2RVyAr5zP2eSOeJ2BFPz
XM/UpnZpHDJVWXaT6VJSjHEh/aPULercsScyN5G0yWFxuA4YPnDWi0i3/lJ8DSlR
11tYJJ4eEY5cq3bb18aAmr3d4P/C96gTPLl9jlAW2M2ZKSRUG467V/jr8JMWawYc
3JoYaVboobX1A0y95BZ/dkKnrKczL5TsdrCBjEY9Sl+/9VXafOwe/PSAI9jpqgbm
f2E73mGvgalU9TqA6ic2xIXcROdxrIBS3Zc8Qd61wsWjdF6FKSSPOI7dv5NbO3o8
EirMhYu/rCkMWyn4kcxNVeH/nWkERi9pk/qeUmPbZqrrR3BbDZ1aoL5oKc/9Sz3O
5bM8ZmDn0QpoyVBTaIn6d1C7M1v7o6L2iSQOOxuJ7D9Ivqy5Dbl//Rvdc4casT2E
HTbdUM8jvjQKPWSGMPzMUFc91tAk6j6KEmT2qWNa4IX1NeMGN/hwRZloyttZOhaX
Lp6PrWCYS+fA/CaBR13pX8BHrqfmSGrM+eomE77Og8oQaUbVZI6eBRN7ZSIeS2mE
9ZYOaat9hLKLs5cZKs9QAbNhe2duhAJmH11x9x2FoRJsgKnJQRjV9vHWXv2stXhZ
i5ynC+/Xthk1nR7UAdRQgqgN6wIc/AF6UITR304M/ZGgmPzRA7px0cRmpXrLmo4P
meCQMO19DmYqmLWbKdyJc24nCuXa+vQt1N8zHMy+45P4zpeeFSYR1Nxleatp5xIZ
DlmYPrS0DdEb9qQtu/7WHjimNUVGpP6XF2V/zeDut7wDhX1MaJ3KoTHXdqqSj1GH
ioop8pVnA31LQ7IQtsnEic7ejQFcIk4DKTTJKHDudjKL7ClZ5PNngCU2Hj6Al/4X
q5NbimnFH6+I4MtbP6CKvbC8PhvGH4Smy/PKxhlxG+vO6xOuE3Axx5+gnHHUPpT+
+7XAurpMWod86rHhY0sIJJG4sMJPvKBbkhfCeTmw3CzI/BFoTz6CabvdgAG0GUkC
xTmfmcF02slGujBOPO6iNIZRKr6G2kf2av5TeTU1q2zepFjTCnJuhlAur2+hRm+r
FKAGek1I3+vxgfqjo/I3VDXvmyksfV9xUF+uw2t9SYjswEwYiDjMWeGLKfMSVG6c
NjnIc8Jh/O60n5hsiWhNpYnfmkHgGfqhqVXrv5OurUFwhfQBvgoIvKG5e+6t69R/
0/ZJrQD1VaGhSjVjnfM8WWn2DLYby1F/eAaZx0LOOt5sV+7gCQ0vXAuF/SerCUMf
GlZw7iLjZ4YEcg43kajfgdcD8ymQQCcwLOCmE5xdUumc0nGzBU4eJ8Y4VgdPDtlX
2clCr2tk3D1nm05cNDddc5fjQz64ePYZoU5KMInYKHxfyn66IsbrvXknoYoGyBM1
I6irpR4U1q3iNPNTpdhuTStjOdfhyyRvLIkbx4O/tRs8wIORDHy1AHC8PwuU9zbc
OrUKv98HNDy29H+IPvGQJo/PBsrRpsIacgxZhnvM6vk+pYXOE44vzet4A525zVFL
JV1xbIeDNfWAB2W/ZRmW21kaRyo3NBQ7ybGAU+Cb595W0so/1/HSvuVvYvuKwXlA
I47s0t992XeW6CVJVJ5yp2wnGfUTXZpT1AEf6o/9VjYphVjjJGAzRpdeYj5OAU5P
1npz+teC2F8ke/67b/HcXbLnUa+41jn6dff/FS9IJNLKwCEtelR2T9KWr7nSuBOV
VKEcqcahQcXRUKFujkHbhC+1w9C1w7VFQAO1hEzuXV0JSmCdt0furWav8jCP2dTt
1pPJL34ePmRxk0c2Ok/4hde5SfYChkhNedHLrpsrNy/5F7Ab0wFdOXndKm5ipIBK
zJwT+9TZGLsrHNR5T/vXNDxFmy8pnuJvwtn2+B88vfJyROTAPu5H9jp0Aih6MASE
6qK72RUo1XGjwjcP5wbxthANVxwX31OzSjsZaqzO4a4wISStuUIE+cYZKrmJk46F
FjmvSi8fshq9xgziVl5IdCdZsYPgsS9GVw8kRrw/zt9/itOmFk/lG7Of1w7SAXPs
oi5UFTxwW1Iw+k332V+lIYLkk0zPcRv0Bs2XNCSyHcAU7Ab6kwaPfwd3+AoHB0hd
VhkZeA1UJatd+L1x3SGesO1TRXHn9Uymi2DgnM2AyvnyZt6hy5KsBpffjD5IyD/7
MBq3QFy0hpJhb7rVweh5SPvd59ZUUIrnG8/6ArojvoxXqSxcMePevCM/4be898au
dC5qHL+RbQG43d2pKpw42yy0S/VBRj7yUAWxGN9W0u0s9piRbiJ3/heEnFUmEXTB
udZBma4rdfEW/XADV8+mmKlAMdF+lagNAhgvvWpNPMVwnW8LKLWhJ4O59H3F7X2a
T+L4/ElIDtfaJd2a35PoUQAgcf9Q8wM5W5b2Wz5HtSTKG6Oz1rU7Of4sIpeWTwCl
3eYtq8Ggvwg7i3MJj6oTD99QE/OiZPMUj1Jm00ncCjj69FVWj/1JtnUTV6mz6n1h
uVrt8PHdCJbyXQE0dfblBVVEq6eHK4HsBCSrxMh6BWUU7NICYk0OCvGl9V2okhmK
X9S+WhCkPTxc8eARh1Hel0Uh2krDA4Uii1Fkc8dJh72wLfgfI0MwSChO3T5TWio5
BZmRZad9/IDSnHKdiWgdgFRXWxqjS6MGqvBa5vy2XpueCGGT9ksrFbVd/9zdWkk3
3LRsbcKW8btLeBPbXar2/IpwU82HdJEZvBQC5fr1fxsCHIVbwHg1mklF8RXu+dLg
wOLH9xSPTiuLzvnQtvNiyZQ7N9F2lxi/H3ohDLyaokTCjAJfAtlbOciINJShBfSa
UaABCOBAAYay2TKp7mFnrr0eq3MOD07acJ4oyRxQYAT/Xy+5FuQdo3ekSOFshIp2
4HStxJVY/N4kuHkfZHOy1LoK7BeQ0KU3UEM2cTW0X65fLQmI/dsFY1TWUZYuUYGF
pVJD9uleJY8ybwpckeD2D1E5WdfKNlL5fJWp1H9dl2+/A3xW408j0AYCCHAyqHSR
aU/kDxgf9ZpEvzN0tYMYKmE7/RgLYMh82PGZV2muH7mBEz0aUOjxqCIDYy5aImKn
8PT5xuElqWY0KpuVu7jqJlSOHWMkNdPqOYRndhaDlmJUPBVZsbP1HGbkdR7Lupu2
qiq2LMhVI20lxCa4R2vXXapr0q/m4lG8bzR0GKkkzQb5X9FNQFv573AMnV1iHL7s
fmss3OlNHqLsu2fC1o3oX2zX8jYwMCu7aQgW08xoqAHLCmxK+HMbxwtkHLJm4poI
HT4wtP8oPacaU+qZ4GetJfsuVMW0C7qTASIbloSryL3911XUbfSXBIYbMTD6/BQA
xFUq1H4m9v42gX9zI2JhsPIkGdA+E10ySJM9TbvFzMv5ktMnU9aFeoTKelzPFZ3S
UtIY8FgY/voUg69dHyzzeXExGPO77lUojqB8/YYsjA5yUqWf0sVSdRmfZ3a71UT1
/Hvh1cWib0I8PLC40Ndk3m8nx19qbjdRpP5PZLbB+Hq1lWHslKI+f5Uy/953YpRZ
OyKZmw8iI6xqNxZRVxvhIuSremNNNFDw92Nul/rChzr0gV5n7Volv1p2wP5DlRKh
fwmDQcwfGE9wY+4H6rDt45I6yNFOPQUXgaUs1NbjORdYU/e9QjsOsW5Wt9fd7REU
zADLoMWeJfYgNb4bs3vtRS5rUSleRbfIKRnpHY5SohsrUDaSRfnJvXMpS97/EsrL
uIqy0RXqzNoc1H9t/vOwKkzcKJDAveU2UFc3oaBRXAU8azbVCUxfqNnbvHadgBf5
CWFSCrNejYQPAruFHbSVLhw5bKHSBgzJZKpldadveitwo//4ImQcVx/WmOMaYjyK
q+Mk7dKeMU9fd1aNPtCd96hEZe/4a2B5TBRgctCWrFsu23CtiBixP6IhfQRmsHkD
hnQKtOYoHfojC6ft2XNeTVhRF4p8Y+Mf7vR3nKGqnmKnPfB/wUDrxAdWUt7duF72
YRZNpF+SpEz2j+9aTwCHSIN0Nt72adBL7abIQz6PXixigW7XM5GW/kfKXTtgmr1C
t6e1uZj7rNRSXcKlwZW0419om4RX72LfR4lC+0qi/Mn41//6TpJA9Ad6KztGDTHQ
5c1IJ4t9zKb7eNGPTSz/+JOVv2q7sDfM1OOwj8E3nT8kXEO0mzLOzX9Bp3PiQyYd
wMpmk/us2pIkh8kvlOEMNuqqIUvXnFDTEjELkkV1wg7nOtX3J28g0ZpxZYhG37fh
n7vCtSyaw+WZ27S5FK7gm7Uobm+8oIVmlQ5ltHtrl0Zor9JDpVGAVbikIDOqR+ee
oazFpCDRY2FGahd9DltH5OG2IjbjwieHsOf3XBU/oxr1vOAS5YsCLGPUyKGm9GDE
YxKi3m2Y1mRJD7r0l0oh7Bjcx5nOCwxOL7pJ8F5xmsVNjfCkfQp/IWQA4mEnNqeH
s0/RTzpRewVa10wqkUJaFTAwVgoFKRkwNEiMzDJyLjxtrxB329AsFDRG5OtFNm8f
iX8fhyCg9Ce9+5PoWGuyndmln5XsiT8axFrMMGCqqr83c7BS2MmuIlJx2/iM6zVo
BXPiQ7Gl0so/bf/q1w6lX9aRbiNvK8myzI1TRunkR5QpBI58eQmooH9T+4X72VG8
gzGT4gUjXwWDasyIF5gOYJ1oBbvQE4N9nSnq2GFKyHajJ12O19EQOMF0cyof1gYF
LM2FPZvncpcq2XiRThCeDI0thaOVdHd5V+m/XsKmdpgj6vc/8b28u72jZ8aV1Bj6
L12Sog7QmPufxI/jyu+UdKQZ8RGi+cs0eKmRDZynumRL9szhSzWdBZwMAhFGkDb/
FeKSmQNjrdUSTk+ggMSp/VMV4/kbbnuCP8irD2Bka/nYXJgSab3jAQyh9elGjGL/
x95/wJfLbeN5I7wmoTqoTS0DAdOdIYmF65u9TQnKWqdqm15NW/E4Melp0/9o5CDg
aSjLI06E8FKe7lI85R6lgmT0ATv2PrQWLpbHkCRu5KjmI60Crn0U3n8f6H+ATALV
Sj9HT2V7IU3qOBD/3i5ygWhBt7wEcfuRQrGATSV7fvsNbK9W5kKjNKYuF5mH/X20
NgvYBJIyhLsQgtjBokybdv9uyYRNbREnld2FA/GyawsJTTwgngLC3yMsu26vmQO2
H+xRFVgXyBVeeN5vA3GMrmblB8TTKywUMw1T7vJ4c4+qTk/Kkz5bnVUTjK/7XIiN
WVo+4kLiO4qP16oXAzB/SDwZFt9NK+DqFI4w279NBtGVM4UZRK5+coyvbK5vb8dj
uaGO1/0neo/NOEvGZue55KtkT5HDxGHHY7rBJCVG6+gGymiQqDEqo5kAUyTKJMXn
Av2thChThA0HL010rpOnJ+y+SErm9cPaEW/TuIAvbLjMbMEsijB36u7vrUhee2Ei
tBKQpFeLAAS72ijFkjAul/boLEh5tIe17sUkFRh5h1ksFPJ9hgFb1Ls5ypGpSQ72
DWiCXB427FafPkBnothsst1cjJ3b5tfqOnaN6ZlQ7nRaoBXOP3vHkFHgd90R8gP0
ke39hLueZwH2Cy3Bq0R3lDwn0VfZDEd2R/DhzF1JkeaEF062zMDzN/zeHADDKo+N
x5+4F5W6tD3sAW3EGCoBXzll6n+0BS8n6e9hXbuPmSbWgbZxh82C28rBQYoDjZOq
WW715+dXtatJjH7hKbaqJk6hFszd3w6BZKCCp5HThXmb0BrHtpVscvQLEMtnxtnF
6qaWCmrLDgi4C4cYs9v/2cAuZKnakAoj8gRAFgF7tYjYfHyK2emDHd6dpvORjPw+
KXBHmYR9PQtDtFFdSgx9ybZ2cYdWpmT6LWtCgIR1ob727BlPqQ+tgQKOZrdyYYpx
L6sVU/oWeU02RK11luuVaKxvqs5vgVWzIOiykMv28us2kYJVkY91r5PzQHb5fP9o
M22J72ubeKXbx67YKS6WvHPDJeQUL9YGXbc1Kx9XnLy5qdcc66uaqHvbJvY+aQ+o
ybId6BWCfr2EvvixYPHTDlO/nEGxes97QzMu7gfo2T9HwtbIovBax7alHc5TdR6D
Ts+G/oSoQ6498li4piGwh4I1uuuB3ab5xdSKO3kpO22+URrqYEeoPFOzx2sM2NtP
a8OaF1lbSJ0rEe34FTxqzqUlQo5EanAyIM3JTJ/Mu8J6mqZGV3PDA64S8ZM9ATDT
A28yeLXbGUAjn4ontidDWG/TfTuIBXFvUdY5YAvl+7sHnWAmbKrEaEue+HzNtgAu
RR+lUSyUvozFfLo8vpAT1Uruc/oOR9dDUpZ4wFfwFlJ9Rkfv92ByJv73j6G3Y9Fi
cjQw57XZXt01HoeNtV9WDsQDPZKxN5jydD8p+60tv5U4B8itayJTR7/lFPzS9kSA
S7bbDHt7+m6qnGAR9flrXqaSMNMe5NDHHUam7DIHu4PRRHbJ6DcGMleuT0FfqrdC
RpeFic0aV0fbG9Pl7aQQL1tNeOA/FfSD2f1b97PuUJm68g3XzF3A8lgUPbdNDWRl
2fknwoEWWyxwEmy5kN6qumR7/H0nw8Jxiqnw9mw4GdujvondsI9T0/wKkMQQiqnS
9d5xrnsKHLzMoMEEFaQ937GWvEV96sNDyLvd5d8Pw4zezGExrtMbN2sG6hC5wgFr
mVY5oqqHFvAC7p7AC3BBtFcNeR74+RHscceuDFRP5DY2l+iv/3WkZfDuoG/3KM25
tDc+tj0MItLsngWPxb1YALpspT20jnkKkCJT//oVV5DE4iHrJVIMlm6dvizIP8I1
oNZ7NiVQY8DtyI2cZxt14EOR3Im/CGYYv4F/BZ9jNBYZ1zLWHOLRHQtiHCGjrGZh
NBAdAG1CwqTRx5zKSNdde22EoTmzuVO0pwTjndQiN9qqrbaDf9xMpcnc9JVyznbe
APFvVlHT04nIb3LIq4cp7/TphvXU7aHEjZoB8WVfrPSvehZr7eG+gSDV7816/Te6
YZcK7V/+d2AroAIDKvk/QWMtyk5Mm6XrGhJr3NYJztp+MVgOCTgCbvuWE8aZbD/V
rlSLjKLGmkcsyjkszGxlJqgzpO+Y7vhUdlC6UGeRJrSFhsMVZJvjqkMwH988zM1t
4pyoE3sVTvVlfmjlFWLTAZDvWI4O8dZcrs4cTCDjbgIIRG557s6ifLCAQIFAs70B
jmI90hCUlg8qHTGkPU6vE9KVGeOJ9hXetr6VUTa8X8qonlsgLhTNWTmHG8Aqf2HI
yxYPmkq0NySkf0Ja98t1+3eG1K7zhtb8xFa444LxvsDx/VLUHai2teE07icEb7Jx
EGZfqgwkZRicaRWE5Fl/2grgYZ4+gdHEmEd2RGaNwNVMCzz6kGBWWSFSXnm2BDz8
+W9dUbSAiGWakC+UBxxzWbeq/DDZdYm6NjgudRSEZiRhySPoUqTyz3LA6mLFlr8y
u511qHLdvQOwSUvKnomtlMDrMTxu8IZwgSixUbvIINQKx/Msg2nL/oz+D+HxZCLi
tuauTP6lzSHqYaPZfyupJ3ySU+WwOIoYc1cFEVnVwAkduWC/E7ZPJ68PDkUZ4SFj
n5jJwMc5TAmYiXiNSmdeyf5c+EmfE8F9f1A/Z8eW+QmCbSmfgKMD8MrbVcWER8m9
CPdQkdl+8JevQrXWZ7EH0lzkO3iX8NaRXIQx2yj4LRLFdt3KhQczO+67oPeIzaNa
wK7exmO2YeMQJ4OtsS2Zuwgkvw8GmCZ9s3nuwqYCwSX/jjmexqxXCuN5i//m2+Bp
BHrotMN7v5PKoKGlAXkDidPJSxuT+vyOfszfHLQJ4Hg71DqRv3fHB2/A7SLSRxeU
Bud0pr2D7+paLPOCqntiSSOjqrPCL57XcmdJfWCgumL8158cDO9yddiHFz4QSXyB
8LDXPwB3sI5wVWEVqCbrMTjPvECM85o6Z5OlDQqSWeyVIk5Ht/8hFcJAY73Zh3pS
FWLFk1uqBtR2u7XsOfnEtGjS+2LmqQXrMmph5WIb8IXLZZ18e/I+OMnXHEnrWmJH
Ik2OgaaBRJKLYT3195slsl8w3t++NuztSDUSNw77uUyC2rV9QpAw8drAtbmCukkw
TaLlKMUxaLlExPS3QPrI1o0/TlBozJmIPXvCXwOXrX1rmOmK7I9ZhCRpdejH1jwG
9Fp8aOwhU1kshxUTvWseqyMb1YW+DS2mSRm8jWErqGZpjh3IMtb04uxBIPnxXb77
zem3mQZqP7t9o5Hvf51oDAATl+UsI4k07pMd2mOuzYNUYKsmEK8EwLsqS6w4UpK0
vOeDPk5qMJduJkYFIR4eEQB9Jw7ZTUcbOAzc3ReikeB7CH7XXRaLpfCuluPKipHP
5wclWtbPriCVW/BTFKLTwXP8b+1fKs13D1kcKiLYVucxz9NAzTu5xFaTUNKj6NfB
41TOO+O4IKET/UkR4JpQ/yTqvuXyPSz7qtM5y2f8qgYExbBxEtnYnqKbdvXjIR3j
MdhpKnGYZC4qUMnlATmkLLWDbqgXjr2ejZkbDyvVWf4x4kFjW8uaEd8KgfxFyLkx
tw+xpfyYnH1ArsWHqCGnGdo34mtD4KuEBn3N5CaN1+5OT1tOlbEpluODxcX+Hv8S
YT16/c0iqKttDNWQWQ4r/LHdi+5tERalx43kl3TC5+9V3O6CHSLjoZ0Gh6VKRUM6
+pG/lf5Cl3AwNCBXqw/2OfmFUFE56PqZOy53DqbxC60EonjHckb8BOBIqYFfgwuH
XWF32K6tW0OZA6dZ7Z1U5d2j5l+HzEMFtO6IVHgAA0XSM7s1mXrGLasco7KPOffu
vxhXFCmkgdVCpeOw1NGM5CO9bvR/ImIbnpxPKwXl7pagC/TBl3g2uEjGyCyMo6RE
M3FZMTH9YopFQR7/UGefMcNxJqYQoBuVmpCim5nXP6JEuY0OVm1CrclVIWptQiu6
y3dhz8PBvZ4fZyIV+2bi/cwLDDiWepy8OTgB20+u8FU4RBU3MefgPU02H1W8KSWS
jCM0btwXFHSwGMCK6voEYwoRcZkfTEblpxNjjX7xc9hxk43GeA7J8iFaWBgxXyOi
pWKUQYI0bRaL303uElpiiIczcqz0A4iZ8BoHefCOUROh47yLt8Rlp/idVeyYqDNs
KamAwFsM+UDlnudUVSjEA6/TRrq85+/fD86Nr2tt7jofBz1eNHj84FTYOQSIbkzV
1l9CbcVqKxUnXWV1HYmxr2OXFwRhGexthzLkue+kV4c29iT603BlX7Stu7MMpU5e
snL9YHX4dr2vPzk/O0QKvYYPYHZmlEeM/9Gtrw3afXSOItcbcMYJT+vcZZBzibBo
OantMCO3Brta5twe1ThOCANSAqqxPBCEPSBO+o/F0X+Enh569WOVA/fPuNlG5T4t
Pqfz77Fv1yCdCBUwMoOZIZeceaoT5IS3xh7vFc7hhJ3fdKLNEo9GikSMRh1eBGO+
eEp5O6EiXnEzvjXrHV6Id9Hyl+KARBxWRabWpgAmlwJfxP2VyDVdfu2+O7geXDgf
tnh9D4kun9HQMQjoIoRDi5dcFoLKgXF7kenFOg278DEizSuq67Q/Yplwevfl3pxL
cJZut4Ne88Zrie+jXYUFDWR0KqiGYqMKkO/gT/sbbM4j3Rm0Qt26vFH+QBgqj55A
40Jg4r9+CtOC7Rn+uSn0jfFLduGjzCr6I6LIYgL5G37C3Re2n5z2QImBOwJEL9iC
UcMd99jg1bBavs5WB0NFsi1IvVChwn2K15B4VQL1d1HM4PpJK77a+a4FEAnpX1eC
MurRbcdlBECvlqinDzbuOnFQ2JRt0bgO1Py8aB7qZes3h+UZMKR9mPv4vrO7Cvqz
z0svVYdHSxcBSVg9rL+uKBHRbfJBS7qHO30oxGLWxDckpvg3VNPBIxNAHVUGKmwU
T2QgkYt3ucStmLXg5uYieeiN0toRqFd0xd9qLwNtQwuUhWn7CoJy0ZrQZmKiSQ0C
ouqVl6SuMCxF1LwjFLqnKfZ6b+91k/E0QS2Lt43DAFBPvwRWSWWmB6Ut1vmRhTvn
8WXLkSHiz8HXr87xLts+IyMul/9CKTNZdN4lTn08h97pDaZZDYh4iHtrIFw96H/h
2KAmsFcxpVrRnbz+6IVKxn5XHcwU8uw7joI4asonIT5GLh4ephGyZk63AzzxzLWk
52WVUftcFeJc4Eqe4WgQ5ZMHPeI/MgZ1x61KaB5im3e5tfzlTGLSai68VXT7aadX
uexpErltRF7dz4arqvBscr/0eKyQZ8hcOnXy8vnOsmcRzqzDSmzkIHzb0/sJRB0h
NsfJUt816QbRkQSxkfPnGqa/vWaORogfeNr0hm9ohlBae3jgzLmk22rTzgYmDNX/
6loywT4KohU8jdsiu6HcQ+ZHq5aXaLBbaSYbxSRzR2rPCM1gEnsInwV6M/p8ol1u
dlw0nhSNjZnySjTBlellTrjNUdYTDoNTgcIC4Fgf7qMSBgTLp8vuH3pTWyiDWCCg
RzpsHAwu36fhFJAyHxnUPaSr1fatMP9aZBJrFmJaGtxNnPmszTejcqHWEh14LtCU
TY/2jDf5tjYCmoFYAE+GkZ37IFpfnvWOvU3nDHvL1Z1UWUbSBQYKBjVJcsOn8cJu
2wnWg1ZlJVuJfrjioaMBKU8xQwKneGWAT58sF2Muv4vGBp3YWA9nF64dpbvnZ76I
kKbbjylUQHyIHsmO+XW8PxxiCvnKB2AANXE4PHxgGoL4SsJqQkhFJdVMbTniyUCo
99SoezKHou9CNRbBjDr2qtaCSel4R93Ej/ig7SO3Zkq5GVEdFSCthH6JrlhrFf/M
eJNuUHSB4qDmGtOjRyl6PhhxZnc1uCRoJgUwCHGwTt4M7CFrBZAxbJmbqWCDAr3t
l6TmJkWEv32BeN4oIj+UDYtTX8UimKAw6p/XrmWkt6wdwH7GUV8P9OGQrjVl78LS
DDmYcXlbPBf+wPdD3xcM4fInQ4OvQMkSpfOEj/KTaL30lFnn0e5Z4a4rGM+LQ/yP
dSivkfh+QUDA17LlkBZl06C13Fyf8Ji/Vax/ET4Fdp3bDhJ+Qx1r1tEmPLWU2dtU
VW3L3glaK7VeBoONuDDxxywBOhfdol73GjTvIZzAyosfe4j+5mpTmzEZbEvZ5IlN
PoBUy6Cwi2b0UVTj+jfzp6w6Wx3B3Ed1JiTKxyZEUu6ysNg8PbY2oX5X/iACCxUS
FEZSSONz5foku0kRERrnw/k41e7/NnQQf2ZPZje1ZQJ5BuuAi/k6lDTMpa1/UX9L
7ccsf5zS9aP/1GuwCVibyd5IhcvzVP21H6lYPLRCZaLjp65FSllJYfOAvkTfRsKf
STwo9FKLuXMalWdJhGlddjxpZEAy8HxwTkWKt6twYeL9/RS5LgSePKBMjP/exS2y
vVpcvTMiunvIz3GYzuOAnOs/Gq6VovmNFaUmF4hlZH5KgyhiPEE4xgcce5YZfBJX
GsSsF/GP35hlzwLf0Rtgvh9KOImjoWUrxF9V3pr0YBCQrFflAs3qJZ6OFi45sbaW
APXAGVk29GXzeOr9S5DS1bXJT1KgESC/3YvamCDfSZwMklQ5Li8NfsI6M1ppPmY8
28SGs+dSMftKYmefhDl/gjgxajPRNyMa7JM5J2OfiHs0rhuvJXUUnqo/pvRmRs+T
ok288lx2q/wI2Jvti8XjmPgdeNOwxyAYFdXcOlj5eKs09umWU7g0YizMEpag6oo+
zAl0qyScuTha6aRNsBccHbOH3fMH/AYVWq8JC2YAnIK23uis+55onXA+y95hVpw+
y/IBnPnKpplzC6z6rbceOoV37Ao0M9ts42l/IafQAjwtDBztjNGL+CPnYf8dIxN0
PATKS9KJWocIdz6YbcUdXS7r1CmjmTmIN2b2Y2D8V9GcX85o0xNtAa942MFuF58S
mFdKKdIYghczdxzXzPa1Bxs6xVOQUXm05ZxK5zNUshq0jGFc7BABjt0PwOO28CEh
m/j4p25j1KD5+RnxSym1+bScbhe59C7pjbFQ3EeZGCQ3evii5Fn5+YpyAy8ne+qu
E7upBVfNJpeBuducvoaTMpkQ3a/E6UPwCcuZWlJyB/fU3YX5g/fkjZNmX5w/mYum
Q4FXQ0LAeuxlqoIFWuzd+hys6tstf0oem8v0L6Xr/W12E0dtZ061HLsmWKSEkT3w
s+Cumvj5WHTuldBva34/rwoAYfAKyStlAVIUXDyiSepsX2HpyIWKKKpuvlCWLIuD
ElGzZUmwRlUuC7Kq4s2eK0cIjvjAu7+v0Tb3krT7RNn6eFfGWwYJZR15PKTQBczS
5HmReWQLrp9KMTqHzLa4ggvx8kUy0VP7E9GB0tN0F0tWVJnQuHUZSxc335B1thvw
oq3r4F/M8EOV7kGWxWUWIp3PHaSZ35+59PlJPz+e78F4838yHDG63Zp8Rgp+pQsl
duouaLQ2HH4OSRZ4/GHmQrEDp+psucaefoApCQocOcKO34GzeuspsqzlJMBkyJId
NF/qNdIRfEeVg+MGtnDkNUV8bt+L77ogsyRYwL8qzDRbf5ISRKKA5/pGdXcc0VKn
Hx6I3169qJvWuqOznODNZqgReBB+uf54/PXnXjCWyBemdunvvjUj1tQiH7T6mIqF
4B3Hht40rgUsoo+Au+GqzB9TCdHshlvkOuJ45dH+9F9X6LkCwDbV0uAocZs6CJvZ
XDojO0rc/ukLUNT65w6DdnvXI53JLlsKwezNAMx4ObkcTRSw+46Q8BMm88cYM2kn
IBbBI9MyEK+hLX9mjkBdn/cpHcQMx1gtHvvKsggIHDf4Ai5fe1Cl8VYhkbjdvvjb
eueiT8zLn5bu5NiAQsBwoDxDf/9EkfTkWRu4QJfsJBea6xBZ63CZeBRkZvHARneg
xThblmIb5x1rHkrwm0ED24kVwPw8BzWldTl6fOEiVOeIOktHJblNQljneKTyfS7t
IamR5DkquUmt2yNQivHpI60ZZQrR1GsaCJJQmhjStvx7mOH27LTrPxaZ7HprCERC
gt5srXHFDFpcbMp6VXESd6+7aQxPEMODkGaDg/vGB6QBdYk4Sf4Q4iFZD7bL3qhh
xiAdVmKLgVd2hg8MiJ65n92qGU6MS7T5vLSKr4YIUDlU4aZ0lVORqPmyiyTtVowi
ygSTa0uAzmwAFdxQCdqVressSTV7k2zdWt2yJUVzId6oeKMAOcnIg15d8JWbEKt6
MKthm8EY5kJLibasBZVw0V6uQsClMaRA+60CzjGc71uHaVdBfGZRQAddzVqIdsq9
m/rhIqzpB/lB2bs6JFJq0r9HbHphOUj8n9x/ogtROUA2W7frh/S0yt9f/ckbQFEC
hA9CkxAMxhPnU1R3TTzyTGjo3H6pyx4oEMCm+o5Z/8852aas3g+GWiNlXi3MVNPo
coEzUn9QD0ONomfYnjr4n3XWmENFQD28wCYj4/6fPt8oekv/REZgvR+HNEJjb/7V
VVzvTV+BeLRRMSe8vXj+8wJEDJIkv8K9MVAAdDVCRdpJTQbiWKZqXbg6CGae0imR
E1i6haxGQ0CWcRge2nKu+m2Jhd4iftJ1rEf8ufIzhF8M7/EwX69os063y7Sv4wPI
VjUD5egDIGZZeQjKQPSNcg2LztukTrWQuop5am4AfUFAknLLnbs90I26ZC7v3Eo8
J7clmpQM3SohxPo3xwD2XbWK3CdVm33zmkKwpjFER6A7p3OP9HvgWcCQppAvF67U
JGjWu1NDI4O+auHU6m3G5WSKO++aABTBypF35TvbQJ0sq3bz0oHuHnySPXdqnx7V
d60GPET4vuUOcyPnAYL2ywh12OQKX8DunW7RzwQ9OOyX65hkxzKcmKjmZLZOL3Rd
KYTUOSWhMniDexeg+ilwqjDSa5gKJM7BZLiuLtc3iBYTf4eIa5K3CpB0fe60mUgS
rkzDu0gWZ9/r3ek1SFbgHb4+7YiYCrzS7PFobGDpHt009YiHtxq0dcNwAvjpYVEg
M2bqq8hTyuWPMewOIlJB8uSBGlMB7s+2jjqUINrsDEZZFxmjlVZVy5jA+Y2XlcO7
Wj2HH12vjvnqLWBZlLB3AdpIDl975N6MEBu/Czs9jbtGLG68H1QPbsjJrYu1yL7f
/tyqARiMMQhahBCjPqjyOjsJyUUvQ5XSsexHyZM2zUP4ZNQBjyvSeXBKmQGthYWK
bk0Ns+jXdm6g3WEHYkN7Zo8XVkgczY+v1ZU9LDVgxXFz7wrgQx3k3j2VTDmYukXL
l5WJgajVjgGvga20ik89iFm+ncgxVUeELBDtGri0STM83oUB6+2QnB+5qThSQykl
4xtihdv74zXXMXuXj18bxd5MsOwi4OU/VPd3WOxqkG/OxiXRdsOJ+4TB6fEt7uXo
QJns6cELZxpEXLohiDHjw3hfk7zfuJ6ZeNMlwLdrl6sQXfWS0EoA1aVpQviGnapN
KJc2EqdqJNe7yBsFt9utfkrLai8O+A9FX8JdITHqtJRHJpzoow1EkH44R3QeidPQ
jj6e5Hso0IZj9fdTX9ouZ4mYv10lBAQ7jUqPRRvnQZFutnCva6tYnGfvAsFZZGRw
uq3NGuvcdawkcBQ74rm+84d7xzq2oi9VhKqX748JpaY4eJh4jgBt3jff7S/Q4NQr
WgfSzm5bDe4NFw1psknFfknRWWUmYiinzE1YlEFxXsyjSjtQ2zIAowyDRVJD4uLQ
Z5sm478vHXwY7JKaaV1kXRRowo2ZyW/J1AE6uY1ZxHCDal5IXTYhgeZZlA3HdaQO
+Ztvxcms9Xrd9PjYe22TDz0zXvPeS7B2nE8/LjpbCZAO9tFJrNAFZzYZaTkZxf/q
GOQF47KtljjlZF6bdSM7utHR6eD3m37aN7OkdBCV43kHgbkacqxNt3scsgAkZ7XG
+DwQnuDFhKcmf7ka+9rxNJkmD/Rc99WK7WGGbLJglHoj2B37rCDvhPg4ArYxGroJ
QtLGzZHP4ZRMLX+wM/ML/P0Jxa5c41AsYQQipE8GisvWP65KgK993by2VtyMf+rT
w58lktfOw+GQgriRnvj8qlt9TwKBVMmC2bgESuI7rZYwNa6GcXYNBPUd8+a5XLxg
DMpAHNQXzBpmrb77MTGqr+jDTsU+zFFTHrMz7jIOEKqavjfYSa4qPY44b6GdUPup
+130D/f5IPidI1feszpfaxhZqa1nOfZGTwyMkHcmjNIJIRJ1K3N3SujBRmjwQw7y
frB5cWsysn4YwXg/k9hyf/q1taA1WKYR5RSMk97U5231ZruezGsHN6ZRU2NlAJTQ
1Yav6ljiD4gXE/X31KxOmoqGhMYAIptvsRfO9KQsnAavlmJZFFPBGA3XhuAgRUOu
SFU1jvXhmlBbKHk8XBd2AHFyzQyHyEDodwoLLdUKOKXXJWFO548MVyhfGepE8Vtw
3PWw4EJy2NomWtpOPjZV61dSUW4re6z99tRQr0uSCfHFzBRv4AORTnxB/pCgP9Oh
YdhWdEecb+mcEOeUL7bHqtffruQDAnGUICQUNvI/yb5iVqAnTWIHnXHTDipH4+AN
J9ncJW8YXLIftTlnKL1g9wIxAyXoOMD4WrP49sJKFEh1RmGpN3O6jRX7hq3Ym36y
3MJ2hdlfSOdkBtwmLYuZ/fK62bCxSzAP+NvmJ4YevBIB8JU6oBBeiNUXNOZ/o+bv
WHQnq0gxdq9wsJ2ePA7OYV/kxBDdQpZV1r3Lk4LRhgBeREKyUdf0RI99psHROIbA
5QJu2rW3TfyGVPzdH1PvWeXyCEQdG0c/KVosz7G3jMiJrrVoDO3O91qispit7XFH
I8AqFvhD0c4Yqzs1sd7HtWG4HTcfEzykUjdTo/XR5TD3RFU2FBZdKwh+mgLeuy5h
97A2aAm/ZwIFbofrtMjnk6mVh+O30a70bR6nU1uzm2uUggDKfuMjz4Hr+Ku239TT
h6EisCf53+dH0I76CyLfZuT2rlzEgzGANha9K05F/RWPDgO7sHPY++yoo5ukJnhY
oA5vBxfoIritU0C3d1lGcReKpVICsKFjf44uZjyHmyQffyf1ErWdkCwH0WeaMguR
q4R5yYLff5Jespq7Da4B3Op/6Rqxk8YQu1oxJCPHS7DwvCqlBXQjwXxxXcvaeXqM
GWr7/1u3Tfy90Db3coeolctfoSejL/brOIzLiPHUyfbzl+GhJ0qOFZt3IZKwkE6U
e8Ee2wPbpGdJPvO4gzNcJPR+ze19wxuPSwP9/lxRj+9tmTn2xb+4z7MYRz78WkCe
NNQUQoY6oHxpiomM5GLUirOxb7SOnMGzwIlmEjC2UXfz1W6Hf/bN0L/HLjn5cpFj
/3Uz+/dEDboggRfOR7JwEy1qy9TBySlzwyqqn/Gvm6pJ3mR3sNjFaAbcrePhqN90
plJq0WbJ8C5gAQSVBUfGZzvZu/wg1hoE464eeI6BOPvljB4PnISyJYD9yNgYgU4n
vTMXpLLwf+dSWUTf8P6hpwfAUvs7oZdNwmI4nN7fbaXSiMKdB5FSpXctO0eWmABE
xO30tQDPYwHo/cyvijdtC+/dxRIXVio7EMros3AEW87M1eZUoptE78UOpfXI+V3x
g1aD20BL3W5Q5mti6VWwJzfICm5AKc1DCG+CyXJ0tDmuD/PoAU5k+GUjZAv0u+UV
Sb2MRqPkQgTARu67hToG3R/WLD/Iw1LFkwit6jfVY3GyIY/KCsAu70mCTx1tJQiD
oRHi50pIOutU7oIN8hyuHXacHKeWfOxU2UHgGZyBs1Idu/hk3mA+ngmRZe5YAJ0J
TD2E4wfSxNlroXryG2Tr9LhS/rcN7BdayF8kU2XxYnPsr8YI48x5H71wwswYK5ew
969D0ooQibkJdWJ9sttl+Wz2NGr0ZrZkIREtkChh8khRyqP8QWs7LFLW/1oidyVD
E1KxLiCQdTKF+R+DZJ43qyzbaMy/x910WXLe9OihaIAmikH0q5Hhxa+Ez9Y55S+l
4oPOlLmdwv8i2IUupUI9r1ISJ9xmu8n5qRSnbMr2wCIzMnfThWrQt88ZpR1wUv0j
pyloXCxsK/yw4lv8vtymLvtNjcvWfOEaAubJj1eacGs2CU4KaLrqqyNQtnXmMxG0
zsFEkAHBriFvrB0kwmjRPN7Mi+qKsfQpCJJnXBvbLV8Desl6JLmbNh44HFE8tG53
cxZOhlIRQlcHcdaemtUcFWajzv0R1csUHLYvd8WxsoyZu0UNgW61zaiALtAgp2T5
A87UA89tUHgZn9V+iMlvYikuhwbhJOkXd2Z3b52+OhzbX+1ux/960qaaGBVP/KIe
uhdWTQnOlemP5xIUyr2ZYazRDs0+H+QenqYEeBp56o1MxB4vdlN1Y+KrgM7C+y0h
gQ/VBSz5jFvuM9GoKfBLnZZy3YIkUIlWclpFT3/akr5s5zoQdmrGNaYT8PhM6l0W
r950H2F2CRrOd48KxZGvEm+q+jblUWQjuXBzR72DEVaEXFVz8U99tdGGoYQb4VIW
W4kzGK7Y/NubB+uOOrka4W86VnmtIyUW/FLAOcq+pSXM4Yde1r9wv8kvna6r7OSu
AKy4f35mcVC+empRQnHOC+r6xxni2KymGjy7dFibUklhWuYfS+tJQ45ot9lIeI2n
IHwLkuXv6LSSbFGrnnKjD6LVFynzpERta09PEobP7p08FgUFE/zzmMlbau0Hc9co
yN7HTZI6yqIAcXdPUiyK5jB8VDxI/r2S3ouL/tCILdjcqGhEsiYsDzCnY9gpooi4
r9b+ecR+hxDxu0GtI/ujnlMadCO1M/79cibqPw350VTNywauwdxrWW6mFzB6Kl3p
0qVJxZkkaIbdghiEIz3D/pk/oUoX2YLAew+iVGdFOwAOTec4DRBqopHugi7BE1JN
7uFCuYRIOucTU56Y0OBVLimkHrCl0724RZ+Q+qsYG8KrmKKhYsC26hQNFPEn0GSS
ZdHLjt0K+Jcmmo71QavxjQxVS/a+z+XzoFEqDbpaKNN1p1sogvce9x23/yONp3KP
vEIKVnOLqoD8Bg7cpiSTh9VENkPP7U30Bpcam9zWMUfukk4K+5oXaMVHg6DpEyrI
A6KRYJxUtJyPPz3APL2ipzcWaOkQnnU/MJCInE5l2wsxeBp9EZTpBEkAk/FKl+W9
l/RwLVEqg8QqJiJ9Oq374mMad5mM4/aMh7rDROL2pGI238P7VgPZlXvK9/WmRxg/
DHdMXE24t2b0E6OODo+Og1ibmORfgOK27r/17cAWQJG3yesFCmGFAMJ4wIv9ET5k
XXGEcGYQDYUDD1ea0HiP2lzKSCf1VBP0k8dn+N7JOF7p6gd+3R3pwh/tmjfe4t+j
bFb9vIMbW3soFy9tkARrNIt+7fKGGGXcSSq7ApiSmXowRY2D836fS6RC7AoER7IE
m2LtWXhuW0Tl1I4agH3HDSS/8TJLp4OJcQ2TU2C6C7s3jZXY9wjszmBLuEL36m6w
4+hiPbtk4c8OAhziB/nPGF1D8v7sQGEELcQD3wVTl4z0uFmJgEIUZRboKrJJZzAW
CCNUku21ezXZcdMKPi2IHrNGZCtWVLo6ZIEGCeriFA9Y9yaj2kBrbGPbeMSyH4zC
U3vzlfM7eFN6gqtdtSt1mJnYiPtIoSB9eQA3qJUBS2PwkNcFr8pgODfinjX2HZR1
5/6UoDLs/feE+LLm7IFY797FvHYpLZ8ZTbN0cBoAOA5bvT7qCtN+aSy17cc3H1fc
nk/2J03Dz1CKdzNJScozDKlhaed0UTLOKlgFY30/fIAni5NrUMwEzlAiENsLID7e
GJMFPzrqBzLLD4SGQVlQ1NegVl5qTgl2j8jqcADe1//TzDRuAAelsuBgZZAJI4CU
hOgOfui217EeQPwSNYfY5XyV7b4vuze89YCC1cKLr1nWGVVwknpmXkjNtmeHPSCV
BvvfZoFggmBl3/0G25xRZil3FtpL3gibRztUmf+adjhgGs8Q8uB0zsL2OgGiLThd
7tBTM0HQ4PCz6oT1/hjjsqPUZUZfRIlJT0pKaILUWUm7K7TOsRVucATZ2cL1s5Et
mOaoLi3fChlJBR+/rH9zW2NM8SplEba1PYvzti1Yrvk6E7FbEkRnAiYtEmUKlhfv
PFqNU4G1EJEuqltA3szUUmZ0Ndrt5OH8AFfaKFUBu0p2b4Vd4zwbjqThU3i4zejP
CEYcOAA9Gklvi+/02lsTsDQ9AkD5csKOwx1eJ4K59atUX8kA3BGLxRs04oD12XXn
mbVr4fV1u/4l4Jtb43+kXk8pNThYauPk/B/C1cVkBG5zdDXbOaSi3XffdSNTeW7o
ejo5Edb+dNbOWWw6eta9Q5HTgMgc23Iuybm6V/eq7yDKa3lrknEykOsbyv1SpDuw
slwvCnHfpzWtviEEq7V2bwExDiEN3qtZZcjEauRulb4Ve3/U5iTCspcEcv4F+aE+
/mTsH7RlNIXNmLTLXzOsybL9/MsG/1SOnD0uS8hxQ2ia0s7qyqEMcWoma5XgWmO5
A91xuVUvvR5kNUN7AmI+3CZqpWZGaQx3h2KYAgQNXyD1hSNBC+mr5/8542Yf3iyY
yvBUyEv2wsu7hTzsdj5v2qpkCEeV5tt040Oc1JoWJ1OVg2b9vHmmAulBxyEapZX4
SMQTAzPYJ6D8PTxojUbGyTR+t/CeVBwlKs8TYA/eu47AWM7sjOQUH6uCwXD0E1Kc
Ix4tnkIN9hLvlusg5aisHQEuBKaShVlx/ujQdHIdcXyfEp0MRNLX8MlWrd7bSqGf
l/1uUWVBOmUHOIM15NgR+XFdQfnUhOd8oCSJalqmuVe749xOjAZavAqhnS61DVIU
ztqCf54dZ433pVprh32csWdxhML/cJ/XJYT2AJPnTca38WmDF1AahlghYHjpHwTQ
WH3vYUgQS7Qeq+tohgUYkvjLc8wB4602ScydEQkAQPu5linMZS+VfuvELtyAVUva
RBGfH5S8nFRiNXIEjHfC7O4Xu7cIAKhqJ5YeNAmntXNEOt473tqtPp+RpRiTO5GH
ytPQUrl7KbEpIdWk0o5oqb/dqao0X/zlJm2DhdbhD9AAua8LkRFpfQTptzIFsbgQ
OLOF3/MGittxAuRxcwTke1iuTTGDl52xgavpenNrmGdqaWyga9/UqFKysoIW+7bK
2946ZEDk3AQXu7vk+osriTdgn43BVrD4q8VmKdqU4Ei/uZQxDyXyfQbzMkiEwb91
u/kDCwubjDfFEk8VJJIjv2dndQBYsa0Fg+JtV48QR+NHztqn2xVe6ObX/NGfNjAb
hNlmhX2IqxxOoPwi6IEAG1aSBKLGsQuJVo0zdauxMCUT5kqMl6SOKQ0VUhp0PRuX
dMT/EhpVx3DUZ4/JNYkzahwH+7U2pauWs+Y4C2uKikjg92vIp8lK4vZoUEACvcW3
qTLKhJzqYORiVfOJJ78OeX5+XevMDoBY0G+eu3nyb6LPjbxgY2shPDjqgIVVF4UM
ckbhbsoQLwz2EU69y9daMqWUg5z4agOSYdSIJWcri7k6Usm4HHCXXcK06AuWHq4m
qzTyut3SI+B1vImuRAdsAePDdjSM/klYTbiTBOgc+jD40I0t4ggOlIH2MJZLKFDf
n85HYtCVLwflkPf0V4QIMLrwQfmjmMeo0exhp3hMM+sQqv2GZe+GevesqR7hd07R
00i3yf5hLbuJ4DvIELyf/t2gaI04VXn3fvMkOQsiHUyliJKyCZrcDMyolwvvGEkB
i97f3lcJpoJNV180TvWk+HMaH9KfhDVPo4I7q2uwu49jN68vkx0bvLGr7SG6APbh
TH598NCvmLTCXi/NwiqcV84mmspBR1EkEQ87lIpZwRUeHfdbzFhpCuUxhLY+av1f
6aazofP2+TWGYjyYnC8hHyARyXEXx+ZWe8iaiT5ClcsA+WE8DWLB/mc9iCwUoV4Z
axtZJwBoi+Q+MXOWXPX/d8ThIEXcP4cVoXkUaYPiBILHVXwRweyD2ApwtFrsE1QJ
jSMaC3hKQWu95+oDR0929j/MZEDAhzAMUGegIUzcqkVOx0I0jrOuM/Om5AU/SKk1
SFgeprDljNsQkOfq/7Ll8D3EX+voJmyuxI9vO4Bgw5M5WZUxxxO+rp9v+gyZfVXF
ApdjbU5GIYamhiJnVFINQLho27spREppICl0Q4t2BChgqg26fYxeEHwrN4CWMt+8
R6kzQJBRvIWmy2AjiCO50HoSyXTYbZReVvSywCd0ILaMNEoGnEzr8KYOBB79ViBb
s3gjIHACLlgfCfkwnWxAkFqAIJpd8iIYtPoawnKPmyXnx4dxPSV+LWgZUT0J0Lgq
0+5VcgCieHjPaIzZlvuKsGW2WcKbLOennURg1htN4wshGNRpitk9RKBO82kRARbH
+cwoTYe8Zm1cmmnAWICpSwWlgXACJln9LsPxn2dgvt6iUjpp8S/PRuyOwkDshEmX
4R5WsRDkwrZCu6+WFWag/UKQjlDyqQKcK6Ttf6q8G9LyqvLSRemVR23xrnmMfCvo
l6K42vuxTkf6vqrST0Q3x59P7vCbwpSzMUchoUi+47I9mODA5qTzzzMgu4wcIBbv
zGnHh8fJd/ZELLfxLbtaAZYjSFN65Ss3Tl6b18Fvt53gRL/dZzpLJCs+jmE+tmGd
WquUi5JiauXI7BnUiBGyciLFtdaJS44pg+5xMUGnqfQOrsW1Vx1mYm4wZfb9EOMV
SygJnCtp4O1J1tdXB/MaN0VWB+XpzEOHV1I90HcXuxoGAUNhPbJlkDzYYNy/LDKN
4tp0dM7Lxf23i0Ew8aj554ettGsMoLLM3w0wSSdv2rd5tTmYu57BU1CkS7cNlkfc
EBvsFcsDawRiNgivs1Jv9LjyN93Alfv3FDsfL7penMf//niG9qxekDXgNpJYOM1R
3iR+up5uKPUse0jZmyxeI6XSRsbxhSqU4sKLLhirI3DyWY5M//8OTglRLfWOY1iA
xSBXlYg17hJtwVrtcff8Vg7LmZKRGYyJ8xMqTZg6O/X4bXdb1szqq2dWanJ12dz3
pvs9HV5oflLW6Rnv1AEGGgYh3/vMGN5FRuSdbKTjejTq8BOO65hzQTF6NqHqDLEs
0mQS2nciZzd9gNapn+/lzggBRw0sSBqA/cg38sR2Z3ZDEuqJWf8IM3vUQanOyCEv
iaqe2gze58LHvSnIzeTsI8cLXWBwHZ8A2Ve/heIhnD5CKe1UF3lKceQJ205+7w94
zzLnciDyUfbQZji/RDyEe5IMgmSXeBBfrEwQ6h/bE2KEKZVW+leS8GWuzJzYUkfG
MHQQk4U6GutTp5QCqTvPZKMc8gTZzEeADjKa0Ng6pD5d7kTa+JH/HRjO+3a13+GD
nUIv4ohpAuDsH36VfGzIdsmXahnOVHcNczr1hyBAEsa7pGXWV2oHRpUNmv7FIsgY
1b3yxgOscNEOQUYKiPRA+D3JBfeFuD2Y5XPxzbeQeQs43gBbdHZhFEsoLTWwWSS7
4GgJXuR8zd8X1phgqzc9hbrb2I0HFYJg8si88/RKhzo2xfzSPnBSy/I0E9cpVtYJ
r15UKxQMto1d2oLzforJG6YvWfAk2+/4BSI14DlIj3i4R0IowOpNQ+Bx14+JMar4
z35JHC7z7EeRH47/NDnORHpInQxAuWowenMu89j10HypDMGkcRoW+lzJSYzBa6Fd
VG6+FM4j7dqMJLoWHDxO40Y46L0mZIA4pCxrRNnaKzV45ooVhvLLJT1StBtJwHL8
PysrF9L9NEmy/+KOGFYom+QM/D/c3rROIX2DAr6Me0r1EQHNRdHFD5dKtRGtrm6B
0Ec5idshmunSZKG/AbsANFAGmFzvtTfRSkq3ouJpZ7pzk/GVA42uRSvErhaB899B
1I+H2/mvAuS2/avmnN/wTY3UdQtAmUsJFXPegteHleO9TCR1gH8TBli+SB9U7y67
txBhVXHEQdrTJ/Q/jUkIvNnAxoSCIXTX5oL+oAInGkkv/J4jW60z7gPwVWCkrz6v
LnG92pcIantpYv8YGFlMLEDkLl5ze2xplY3s+qi1mNMJ/t0hJoEwcr/7Gc6vJCI7
VNxofGOK+6fBGHEe3L8Nqco9EEBCFzL8VUAQyQNxpE/51dK3Rvb/FTmyIS9eMl81
hA0LOTZHu+wynZOFwKlmUjR0w4dQSORuLNTeyKzqXBxMPlLR5n6RGOg587uqCxVo
6jzfwTYyrtV9WwO8cnLuVkgptO3Hq4Uf/Xu4+DPzWl/R4ZWz+fdXY1/dGpTCpZGK
OB3fgEETOsZXlfB7p3czJRzarNu+ssw8QW2KO9SrkoHZc/aOUjFQClq8kji/yNTO
Vrx/6LC/Dqj/ljdqynAgFamkhLmYrdyaLLgwi7RjxYQgma/RDj3bvqr0ekGZP8X6
LR+oEl9uuE+vFxhf5sKilLHLqJbDt88BUi5NEteFqfXumlJ6jZld1cIUsHQYW7CP
0oiQ6u4jEPaaQ2aEe2PGv6FNfvQ9XiRVqW5KPITgbHuUM+gjnUHW8qS5bUtfdIY0
Fbpmqy7K7PwSypU7frrP+n5wPlgBBQsLR1FW/6TDafycnO+EwD9OtjLs3dNR/LsK
YejUxXsrbTWFVRCHxkaIrptLU5nxIyoJ0aM41ZN1clxTyPc1063HkwMMkzgxYGYk
l+6vMFbXc2myI8/+DRF2o7uNeXlyzoPx27jlBDqzEWC7U5lrRO63jw+e3+zHOzpd
tgDaCGQRTRbog4sEPYm57Y2LkbeN4jNNgVWa3NPvYhvGgATXXI2qXWl1qm5FGxok
x4W/IAo2EGMOv0IVTzQ9mPZdWRwdAs4wt49kdjKyB7mYYhCzi60y1gf1WhVEdWjg
EBwMZRBLeOubWOVV7ww2n5UHC1pj+4/DVngGI8ppH5BPdiCGGowUWlkKl27wBZ3f
qwqScAUb5UXMv9NhT+/keMvWODQt/mGr9TkgsOFqU7tnpUPlsAD+Pu6JWWqkThVe
+D/YsAVMzkB4w7tLjOJFclo6fh9DEVq+xZpskKxxofdwbvNZwhFmlSZgdClGgbUn
IUOgGbY4DDbVG+poqj1tA9FjiJHBhF8Lfvics9le1O+HsXntxXBcDwIJJnssvA8l
F4oUuaXgBQfy5agGsJEbQXdILyPRrddBMWIZeI7iIUaB2x8sL6rNxfVsUVGmS1FC
TeTEhBNaLRV4I5Z0Gh/bnpGKcqzEoitNEKMJYvfTdThzQK7yj790fD0XYOSo4Oiz
u+ud4bY5U6sig7QPD+/XaipNXK9pZNWq1dc5EKCReD7Zr7nbQ9r3Vv5ggLXc+Yte
29BLc3HuvG/sdttIezhBXyPu4bBUeDTl5hh6A5Upe1RYI9rgi7HXIdTVFIi08WhF
asYUlimk4Kplqbq69c5mzDYSZ03SOpdLQBNxYLlkI0Q6WBajaEn7Nn4z5np4M1dZ
1oTjOUl4pgQA3cS89Sygte3AXAagkWlofHb/wPKGEP3fas3vwvIuCutts772h6xx
z6ZHKFzwIBZ8ZayylJGJzbN5/0Pd2oGGKT4zqSJ596LB6KgoFfxfzo+60tZDGhv2
ilEfu5U56NsQfJO/wBNEmEK4/O4b7cYKu0e100E5oR1EY92dfgUH72eiZnmV9f78
5IISb2ORlEvZGFidoZan6o56jruifY0IZZfZo7tujajp16SGGzdZn30abxw9EVaR
siTSBasNa6ZKoiIFbE5U+CF1ng1vi03Pw/vMxn3JU+TxDEHyNVKHJ/6vqbXlTHma
eK//MmL2EZzuCBNAoH6ITQdDVhvJeV26lMi3pVE2hD3bUl/2BY0AFyT2Cv2VXakb
EmDnxS10yuaveS2ddOq/UdbQ4Nqny6uTUAZyoaQiIatT8ZOIqD8bHzgVb4XialJy
hcwdqpy4nq7c7xqdHqD/7GwgFKFXT+PGNfpWz3MIXLhMK5qDwOYH47dOMssoXqpi
yAbciMm9e9SC378+kdnMzT5hgJP026Bd1NiBBwHcPEn5Ug5CjP7wmuJ19hDkaMWJ
wAM0jvPpTWM7D5ERvDzFPwJiocKStj03jNW0EEof+KdUhfrvhbK/BboHymGDRhmx
uPYFCWjO2NQf0R+r/cDdD5/BcLo2uyUlmPMUMPKAxY0DCy1MY+9Pu1kThg3FEXSh
I4m0rr56JL3B1DA//tnPXSlpfuMR6h0LJSGMLdxA7yBhhyVUfqpeR7glrWH+w+JW
3BMbkUwQ9CixmBZ9CYldmQwuRXvKUIFMViYwT4CWvQB6VY3QiytlKnGaCfGwJnaa
te2TLpfN+cQggH0WqzYn4Fq8jsjLi9yuxL0LUsl5glqa0gEoZb0AhdheJtWJDumg
DlI+uXBsrJKCUx9uJL73MVtZMtaY9gKc/WqwFgbEjZpu8YadytNnvn5mWiUX8CHG
8RskHfUzYAUYrgbG1/k4mLdle9WLNOZHLGfgSOC0tDcTw2qEv7ErxLPJN8ofZNet
5COzJe3gRSE7VmrEGqB0VEvvbDifv+bIOiERhd++POHUDTxzFYhy3gADWOUuIrBp
0VUHHRJ6OVxnNbO0y407abafqk2GFWnIWf7yuxX6GXpl17b82pPSMyEeeI2iQ9bh
YiRfexvhdRgA41xJnBR8lax/5+sKOMsewYdoDYxizUK0JDSycVE8l/irgK43qFBy
q4wLamUKen5jMNxX8GJKOokTT65Mo6BADMHTU5Fs3amJcDL9UEmkrUFF1EuVEOWd
EQYlHhtDNNj3K8rP+PheFKFIHcA9nt8zXEdgAjMzueTuXdSqt5Fd1ipQMFFEK/i2
D2+IdFAbeudL9UDMTiGJaNynrcVIFjv9BVtEqVjMxCscq93SfZ35CiznpbCM8q52
T4muIOwpq7SNILo6ALrLrBK2geAUeFwASmU/Q1XZZCVVSC56OM1QER6xIU/9NgVm
K0XSzjGfCsw+E/aX9ZXHWCcGkUtHd62w9fW/GBwbTziY8Xri7FOkZfTYMnL/I/gM
qZXu1WHACq6EQdvrh8HJqy7Sn4rfeao0GYoNPSxG1paniuu76oEe2Zn+ZhT2nOr3
ML4OVxhW15slYw7fr5ebEqXLaj+cCgkIuOHANzBjHOAx9xn7h1FpNQMqyOjfuRDd
fM3FUnPXsiK/pOYYH3UAPVKYGoqOF6Jeb+uQiQCqNyfErpmyO7+nF1+ToZ6wEvAU
/aekd7c+/Tgttt8nl+NsSqccmhz0Dce4vN6wBqmDe3IR82Ry8MFRPvXTH/8E8git
8PZVe94WBd5+RNlbZM/bAblERfl6q7ZXHR5g5KUCH7YP5+O/IX15Tj7eijwR4EeT
fz2lpSPDqv2DYhK4GhqpYJvz9g1EvNCQSAYIMLkgI7BgaY5xUgO4H/pO03yxpVjF
nV6hjYw0+X5q185b0QEXkRZ0KhllOm0nI8NVav5wBUDqR7S+gYzeiIhex0OZjdpo
rGNM/NHySWczCpCtEjrrVYCtEPjqOZb09oEPX9i+ZzyBTuxUg2KqvEjLIkkNb3LP
c9TW+5D68bUGGT+QM5Yg0N4jkDRKOz291minf/EH+dBP1REvMf89YkW141TratzA
bY8RqZV8C/ADPvuyyrhbBnQHWwX+TGlVKbxgoq9J5mU7VptpuAeqJLoPlQKxmmtJ
etfSeRN/Q3NHq6XfPpNN/dyGe6EseOfYLgtBnk5M+ynZNJfW1XmPcZDU8m/Hh48g
6mIdY76NJDH9TXtm9yjQpvMBuUiyK5mNVTb/K5t/bfh3KLT3D1nNJZgarcBFw/jI
ud7NKIZuiiEHw4E7IK7QZ2sEOBzTPkGLmxw2CwlN9o/G9jhEXs/2msCkHLKGPWAQ
nl43sHEBaGucnNleyPDABafSHJk+DK19rp62On7o6IYt2yvme52q/eO/VymXJFVJ
tII2g3O/kZ+szQTMNRHqvJvD52LwvFqrlVShA5ik4HIuaqFV4xLmx7qH4u02U9zO
n56F5VicSRlzwpLrrCwNSB6ebdnnrxDsURZbremW0nJZRrrgRYWw8Vhf5ZV2Mdd9
08loyh8v7ecBaLFm3Q9nqCeimoXyUNG71N0VnDhcrXcWbmbEJWgRLGrTiumptWDV
OP2JaT5LHYYhzw/lIdVa29aBsg2CgHu1c4SHdfAElVlBCqqG4iy8uVbHC1kqE8yc
US34dE2y03u6+XwwUZpt1rhCmGO444/uEPhOzazjU6Sg1RsanO9m5QWz/SnlGW0q
gqLytqdKuqaukVAqG5JbvV+ydpn8OkWEYTjsmE4Aw47FJvlMd2BFYlJb6WGYi+nQ
P2VQVMSUV/NOUD50xmekXUS3vEXeA5SpiYjNrZD8SYRzLY2NCPHuFtDsUWUa+vfy
7PzAcw5sclAKBNgwe+GovZF8yaHU0iAs8Y1SiXxpofm11Skizx6aFfwneMlbt2yj
NIjLaubAd0++Be1EefbPc1J5viXGTLGaBmxBs5ag7Q2GfT1wbAV3m7NFJqM6Xl/z
medueef+RTVitu9WIEfkQLcazAf5TgxB6h/+Moc5kKQYVk7gkwpD1CzH7/5BUy3u
SCof0G349afxi8gThhxdWiwLYFe1ReUtb/m/7oDYfgpf2ieZH0NK2EZ8sS1C4m+c
mS5mnmfgnlANrm/5TmkJdJU0T3Mo+Wt83C9kUHs9MMyqh83QsXAmeNXzNu/yb8pP
7tUm0KdMDG/9lE2czLqsz64yAF9rlYfbYM/0ZSD5dsz+rf8Nql+fzT6oNhRI1u/j
mV8puY0ax03Rrpy6fFDpi/foloIKom1+YNaD5GP3XeEC0IE4r7PscVuUyMRhek+I
toDCokiSQUQGtXxHz0uo+bLscapboC6FlJkXc6sVFGypg1xoAyWxsXBFaxCXwUs5
7vnFxo8GNFb1uSx+e+bi5OhCSF+Mf15rIoCAwi06+yX67Anx3WMf/cIevQelhKhk
F7U3slcmDKsJLZ1jFHVO2X7pdByi4IpGcE6/IiKg5O6mx6IkTd+eZmbmjaINYXRI
HGBJPuYkhYF6KfwH5GtqyaN18n8ubKJkuHRsimTih/jTz8tR3At9mmxBanL0QCR5
IPAiodF8p/ROcW9/KFQ0c/V6kRiiLk5msGbxMsoYXBHIMGTvCqW8dM6JsoiFIWTf
mL2/Usvu7AhEqOc9fahNfHO7YppusnuXlz8FTFEBJhp3DH/Ml9VSlY2Ww2zMM6E+
4UJUO+ujkU+XxjSSrA2Ir0jIhgHTehNmUc5vZ71XGQ5yQ8YRZhAdkrqbxqd68ZI4
txpuGWOOxP8rYKIl1VZ7yAxOF414bLruLVIsOjysNI6BaY2EojDdX843E4ENygOK
0xfLj6wrxEDupN3Em71YYzODLhvGusE8ccNaxpByHRj98K7DcUekuEy2V5RoEarF
RFZv9CSByC0h72gFkFG4WfAEpzd3+KInMDdqfmhYP94Gdwhhy1xQSAXI82UPHhgy
bIeRP3GZjw3Lk6FRIJI8wbLTriTRqAmGAGkiahOqm0LR6PK6asimULtTz5X5SJeF
/oH9DEepSxwuMICXJUeKXT+F+7vsoPwRImdx/5Hc2MPmHaZXKKB34JdIvZM/1zU5
gFFGM90fz9w5GS4CWy35I+FmNj8scZcZ39+9xSln5gl7q6ZepJXIZX+O6084uIdo
nWfrDqDUQMVcQj9r1Aefn/xDSUe3sRBIxXp0MPIMFuKC0zZZigSm1rOhNFG0ZnxW
1YIvPziizqIywZrbjZ8zV3E3TIg0gwddQ18GX/8jMVDrgcSqoT/bgKkk+zD0BWJl
3Mmvq4OgLh1FW+pQlc3ivNXYgAYKKxFSeFVJTBV+tWnuE1XAIkoydxyZayq2FWUn
q9AiOooZsnW8nFcWWqSw2rvAZc4e2YibOSpYZZkgHeQ3zihL5jWN7b7oxONXnO5b
0FSOxsdFVkZ65dkMB6Vj9v5sGYhVtP3jjVdociaFGhFlzJ6y79Qs0LyoZhaj53KK
FX/kGXhF1CnU2ceu/1EOm/km5NGXWM/BWzL+Qb+smaqMgKFdT8Q8nM/n2M9ZiAh/
2uMfL3MHL6Qsjgdro07FYPvjd5Rh7dR9WcxKWJD2yZn0eqAnwJniUqlcWHvqTJZ+
VNlZ0key723GFj4vvVE4UYwOjVG9jeNT6CUan8aprOBsmjpq79SPPRMlwbcsDNLz
RiQItra7dME5A9UJ2Nhk1nnDK6/qtoyLB+XjdkDEYLaBFpFjurQbC64LFAgzDELL
C0M1wSIx9siPTwP9OZFdJ9PtKCDF/kj9wCfzsysVzO2lgeQ0XOKe7slLTHWYHOOZ
amaaiaKZUSn5VZDb8eVa8Ny4S6ucqp2tHTpRjq86rnX70HleSi9FnosPySRi1U7w
gX+TwwiGfjc0NxXhxoMSoQ72BTCustNpI0f6JQsPuGoAd2cu43X2D5ggW2h1sbbs
j/1ighCTVKsUr9ypZ3WO2Z7wc5XXZK3CNQbRJuUFNlBFRRHw9HLXCLfXgGtg5NAH
ueDDjicJbp22I9l+G+haM+C/usZB2L3eh5RflTOxvwNNGx48dSphIpE50FBZbKGh
tMYu/xO7z4RQ8HDRp+U9Jd9sgr+8SEqX1ZZOC/+JmIvmx8CmqnBhknVV+qjTqtDD
xDI3OiSZN8pvbBbSKrR9bj//mQadsgPHsNcWP70ykUf0dB3hdO7Hm7YPYhveGNaf
yAERJGbwZ4jwAZHG2gKTYSNB5NF6LUxDx20GEj5IlobOJt3a8Ffg3sfDKsZB49fr
lrSzr4C+75hbR6RRTpQ+Y4XP5dhty7gJNpWBJndphpxx9aaow0iKX6q3lnIbF/63
dy3KpXPs0JTjNFG/5wJ6wD63xdPiJz1gi8FOn+gQo7QtQsWly7OxLnu/zZL8rMHu
gfWW6ydMbzes//ZUNF/bdRwWqkZXrvvoL6Lmm6W81IvcCm4f5ZjxwUD9RHPFvBH+
MnIHPwoYIVp6s1owYFJVlIgPftPddltGIlQZLpA4tLuiwX1+40nJ8AEtiBcXENDb
5vKSLIi8tjNncb6FIRP9SOI5bWl5sh4/9v4WIdYu4TKnGpzB8titU+NbfohuqFzr
A18SLpvXkcsc6Adh0TfBmeHVe1wfuwjYcYS4bwQescDEEmTzoMprzFLsEMQNmyqk
JkgQpW8Kjl9i9hFqXGWEWQj4arQorcL6HLyCv/LnjGd73PH1du+lCUTugGj48GTs
9PONb5go8jo3kiKOKT1znwAB+p62vuf5pT5ekpwYFW+pHupN11tUgEc5Xw4DXIaR
6j1tDJgdbW4HeCAqegdIGwTDjmZLN8E8LuXy4dBMd5da/TU10yz4Pc1vVD/7Y1UR
r7NesN93uTrjM3aKIEf6suDV97F0JtDRwbejjiK9GhiT8AFl6twKO4qiK6aeqJ/3
tOIctLkwDOCsgIdCrLxQi3+IG+4CSeRiTv70wa71yF6ZR6uJRNnze+okAmx1QBvi
ga1bUgSczh9B/AbkXq+EchwRFquCP1GeU8JBDDI+4iHF9Lv8T4EDAyafTPhm/JGw
KKHVUbaBOXNNh9ZLn3PvtByHA/SzgC/chaUAwCfSC0S15Ylkk+GLRTZsIb3wrLlo
m/ShsapeTvSmkJNCKQDnOfGu090RjeYH726/sgL1DtkvGnc7P7bVbYTybKy9zZPv
3Lrj0Ttr4Qu9/CfSjX/4Ru+bjbxLHEWHWmykk8eG8ot7R3LonpqtRq6LiuxPy5/z
Vq+n4e4Yny6UWB7La2gUbGVxSx0XF+4+NLwKvPbZtBPCOBRMaqLpnc8B4eujp8TN
qwpQuYoTxLDr/gFoKRdte8A9Lhtfg2XMgYJapXxf2CKax7skpKgu9k3ElQLqTyEv
786Ew1q7NWmTfYdqJiRw1i7vCWB9ufpM1Lgz78RAwmmMY3bx3mQTTavq+Q9gUUbB
fZxNfpEc1bZpzmlXLU7dRBrAumcQ7DcigjPmKFKlxS8i3k5ehNH4bKBTZVhOnQBd
nwEcdjaoWRigTQ8NRPCqkxVQxW3iDBRxKDvg/yEwd6eqEyPNzFototS+kj9Agpn7
fE++1qtkzykpQh4AQMTCCkKUUlWZMEHmRdQrrm1viBnSLULD+6EYBTMt6f0o4CPF
o5YieG/u9JgqntGr0INXkgw2otEfbVOk/7rje4DLHBqUgqwTVbaHzpGVWYT+Y0kb
5qvm7Eye/Kk6+Hft7xPk2HlatIBheKi8flIv0cTo2t2R/BOAGiSnHvjeYTEVE/AL
Q1NWSplLbs82D14T6TenluailbfqEayX3bCfvuzp+hb8wy8odf1rBlsBYcFC4aER
PqPGiwCpgcOJ95GRuv6mNN8Evvi+RLOb5168FPdZskDAy/Ec68iH8lptnuf9zeAr
dv2+f7Ym1gvjNe5MCGSMCyn0jWykJirxcpKW6L37Dfre8iwvuWKxECC6sf1fCoS3
NG6TaiTW5tu3uoT8oNTbNUulmDEiNGHKfT/FDbWaTv9H4YDNI1Us+hIa44TlQ+dv
f9BKEbvr7CZKzyEymxr5qdbabma/jxp1yuSdXV8HXIjxLHkE5haUQV75lBTOXS1D
t7cFUpQRWE59730oXahz1sacZFXpPISsiZrELNLI2dEciBRDSVUgxY2cjy5Nsqqy
4izZESL4CZvBfeDglZ84AGBilrn+WiPhIlLb6/4mT6ofmohaoow9krRhHFs9Epib
asVQk81wrrb+J1GPwYCYOeWJU3mQJbDCuHZalnf0UZChzzfNcyIuWvd+KImFNZCe
CKcAbBm0hxFRGLHX+ROEiXHqdF1NxaksB77ADPHTTm6AwQi9gOoKs58vOwIk5i9o
PH34EEfcYolAZaOUhK4tEE+ZK5ehYmnmC5lufD7CrQLvpdtna8nubLjZu41QGdbJ
wnWsxgBqiR8E0s+IV45mySDnulmAJ3SZD9WKVtOmgzcKItXUKYCLo6CSX82T341L
zdN8Rf3yja8wIavlD6WT0xHwyCK+oh8/vgNUL3WFYGgZBrYuxLmeOPLS/YU/t2xh
XBYe0c4lEYLwroWRJzm5AflK/vLsdQwDryzqVDDXg189J/p7XwN3/kx5FISQLbXU
JN4gYwvML7zCHz7xHUHbhuTUTMIwFOlmeO3uDofCO+rUcfj5E3zsVuv/faspmpXb
Zif4X36Iq6mDB12/dAvqyqSUFhi4mbzxB2KxLPpoYQ+fW25Sdtb67hg/QX+rW0/2
b9WIbeVSKsl7aRW+UrNavTaTSNI+WAMp2IvYIJpHdBkZwc6tHpDe8WLEnJoJzTRC
uE2oU10RIm71Y/gDhZNpAAYsABfX74yPHxyMqBknhTdNwa+O04JTRJQZqrSzZHRj
ee8RJgsf5bQTcfVuk7TBV+CpbJGx/2RMkibK3D5mhmmYaJaxoPDf/zegPbPdwI2n
slXPyjRQnRGB5uHx7u4Pfc05xxLkZUVkTYGLMoMsrUPp9y58JZ9czcGyHMA5TWGa
GhUU2kDltAphttK2qbzfX0UCihstMZeLB8EWufLBsdRddsz8LWH2HZ4YUxcypSnH
Sy/yOA5WKa4gy0d0UGuaYsPkQkQFG7rmqxQRgDw2lP1SWXRbIXIDroL5enmxFRoG
LAHQrkB32AVdq/UeSFPnrqV8uSRUNnCW0jS3B0h+U7HxqYsUI1wv/r0xO6oiuNLS
ae06+4S5jrlMEJulVzuamGpGtPpe5HmE+HJYO3XFX+wgZUNH2VTmgtCdRP6QPRbc
eDPPlDxj09dW2Lu+apVclTcUPRyjRJCW9R8OlOoEsIjPEYbkaeFSqj0oCUCEO6nI
4RFlUnnqJHFjKv/dNKoPcURvH8fKmZEowgNpwEz/W6E3Jwx5Fv8VDZVouG9HQxpO
ZbxOKNWWg/Rtg/DY3Z6ybsk4gbxcIcUJzUcrGaK90jEEAoOrW9+A6mJn2a/NOzFH
UroOto5Yx7jRmb+LgI8sR7eaMbneq6fCzjxmYXcYYECAqhUDE9rjyLOt7NGOiS5F
3KhKAkqUyeD6wXOYdTySsU8bqS9Sf+r118kqzW0lQ8qo8eU8Avn+QJ6/Pxq2mBQP
eF8w5nYPnCF2tnkVzlfUL5JxfPDYvXq+8eh8ypdJmt3LQK++sNAfnmxzzofXC+jm
obrwrx3WZBpdnEcmkX9sCLqJl1n+0ot9HLkVKf9L6LIxQt1ENGBKtvPSzRTRMa8N
gOjYdxK/5t5J1G3ng7tD0GzQKSLuIym7AZ7WTodyV13wS66F0ubJeQo8RNX7xyRs
gYhl3eH95Hqd8GYMDMCEBS3ADhbnqOCa8/hmMdrKLJ1zSxBl/WD3HbSl+u13UuaS
lDQxfChmFDH8R+PIJoBjanQPN3OXfB9MnvmYYF3gV1M3LWptw8LqBlyE0LjKGkL0
kmhOju3W6SS0em3AkzUOFyS5kUjTxQ8ZchAyWZDfJcdzPBTkIE4ICWVGqjfhqoGN
fyk6bHuZFKHS29USVIJcOyTBdzrb7PousyTiSWwORzDNB6AFEaoImX++uZNekQSF
XOchlb7Bv0szGYoSPhMg0JgSkI1Miwu51in1fpkq8MrOiIE0jJyyjpH4/HhjcyiW
5r0XaP7nvC6fzppfngwi6NENCHt2k3n47Gbm07U2Euc74ylXnTjgmdukuf0UU7UF
Uom+ex1xeaHWDRcI6+80OjHC+eiunOrVhG/Y1r+ddevp5kXvP8yOQ+TrpauQMd3l
JeqTfPzlceJFms7s1s8187msl3aRZkl6SsA6wi3kyFEgDtbUK5v7qua0QdcYoWU2
ckHeRKWJ18SKVF3aD3lX0UeAOqD5lKofqcfHf6ItinHVoNQlrbF+hCdtueJWUxbK
qn/jZnFCF7obgYD6H1UAkJWsJqG898I0nCiVeus9P5cxloSmrla3KfHUPt+0Z/pz
aRnaXwgYZQ2IElw5Pvs3BbyIRTLKbBxIkL+UscdIQFdHieerctnJcBBiyDUs4B/s
RYjL312oJkal9tS93z5KaQHQ8L8iHErkB/Hwyf8b8pqZhdrPOXY1RiCDdNh9OSD7
id5vBKxYFzHTXvLKcSBQb5OnKYTCwkjxf9YTbYnukCjP25pRt5HuJPP5TcMjj0gx
Ekeigr6LfRtDSyQny/zV3hpDGFHN3i2tW9WrTrao5VrHg3hOiC8PHuF9xoo17Rck
1idthkEVCVRqfz3PA/IDDzblCg++tX3SQ2qNF/zo44ogphL6allIqrVDvxGdjKjI
N6nwDwZYNEcp7jPlZPZNM9HVlY4Zi2SKKyksjLo9Cda4fVu5JqMxcLURn7Vq7aDh
yCyMo/XcYRkwLxTzB0AVLOofi0fLhM53VIWJ4lhUW1X3HPniDNdWn+vICVrlwQg4
cx+1RH38De+gFzf7/ldLlwxr9Wu3G1bbqNHTVTOiLVBQLb+F2rTvbB1h8Qkp74fc
M+7O+c8YtkvG1oxxCh+pVE0oiUnnPbKWQVFrzS3SgFRm2Ywmt0k9umOd0KC5GnmB
uOti4/z3e0tQSu/X+Qnm2mjW5QuB9/qqgrAbCTzqzq+qjWZaCLOJx/FRG6f2rXwH
1reJUDZaEt40aOQ3Lr1w67eoy/f5PD+N1YMdvaArOCW4wBJC1nkbxHl+Czg4a9uo
VLEyHijrkvBhuxzGyL0JvWFmpOP9KLpgUJxNqcQh9SjNrxGyoEz25jhi8bo5frb7
rCecQdHfEUpXBvq/2PnYsXcWaoiamHWF/vxt+2XVUKuHTY+7KcYd8O30l1Tdw7Uj
wNjOovzaXARkdtFjBCuA8PTg6exvvvCRC0cThRb0P5C4WQqx98lBGUVC4xu3QUH5
cATnXt5BJCw2AL2EjXOhWM5W6GWIcsHzyeiQXYz3jfMCDbY+u4iZFb0ZnzSbdOrf
tBypY8u3CPag9T67aQC8LzQ4+GOtlTPCDkJOxVSQpP9KZZ06wYNzgSAIK4v8J9rd
fMyh7EfJEPMZHhrV68vuCJZNhuzrzKB5Q9JN7Lsk1VEXQ0NKiwFmk58QymTea+IB
GPtQjMn1wl7+BaG2iORlueTlV9aLqLOfuwHUOHtHFvL+CyzeOo2YrFzRiY3mZ6rn
VI8e9l95ZZiUZoNqF8MIVY95OOWh1FVhcBsA190o//VkJo9wRJqhxDu/OzSr10fB
05iGRyYQAysAaBq2vZV6BSGj/3jYRBy6SgBhyDZL+Nw7Yd2+N0sgCmcVfwE0Vaab
i7n/d4Im0VMFVzpL9xd4YzKH7/t8Njl+XyIAfu+1fBDGZCwRKmwLlM5iDCWHa3y/
PImsE/mEnNH/TqxVxSl+ZLcMXyx9kRAANBr6WEMZp8JsaegPOr5NQ4l8b4DY9GXd
tncyIThTc4rFcLLjku5utJ922LA1oeatWwmuxKCJoxyCB87bCMlsCkQ5OpqlqRYu
6QV99MgERryA8JmseD69NFFX79JsDt0iaEmWyv0wpkIdU2fircrYZzi14DKSd0+H
lckclxdLxps3ktmoirqp59K1UqiMDIxAuKi6Baol7sPUQ9A1sauZ2jnR+5YsdGTO
jf0/632I7XHSkDHEWEXyv0rphPIdzMoSAHc6/9q0aHSgVeCi9ncWcyUJVdn1gUGN
In/fhgXZQ83WAum3L/sRUdraQlkyz2h3ZR8WTDaHiePi+uPAlHCleLcYoBfEHled
mZbxw2i7GhComlZ6UGHF1mMcGOEny4GBvnixTmQgitK89YA/ywfROz1zGjLu8yEs
BRgReTKUgedkGdF5Wt9psvYeFdtJH8hMvkLm7FSU5Ue3avpXvMfNbcY/D9w++wKO
voxkF743jCCA/SphFt1DCNHoHi0KzCDCPHjSgJUJ93c60d/Jwk0LJSK/rh+NElq1
RibEZFu0JbWLqDqaGjQFHyXDV+/bSrUO+dyujC0BV9eDRLofvL00lBj+7NF1hlQh
NuZvnqXAv8bszkHt5F/KwDPpbZk1tJsXfT26XCdOdRSxDgwu+Dhr591VOOxd3TD7
lMmoEAt+Nv84GWB/jwnxN9/tuC+Hq6cWtu947xLqf4OInZoYIcG8izeyxVp5qSHQ
Ln+QFzyaHABl0C9J5HN7CPuWyCX73WoHzc7FgZS0eUiQQXVuR9VxqSRP2JXIWS6m
9wagax3lRxvvVu1/j1h3GGqJoRVFrOsjc7eQABigrrVplI7FCz1Hb4N+3fOn9QYt
mMnsDP8kRM2nvUTVfPgZxsBP6e6ZfbKtWf+/ppri8bAkTPXeWvnCSI0fgOrqOC6X
mKI/J4mcnjbnulxkW4cQ+i9rNTaa+BbieSslmt+GkwxYub8+AVJToxbarySZgyUv
GrV0i7jXkyNkgCfpG8CUpr/3cNaOYEVcjJH9/IkFddqBA0fe3FffHdr49z/GpxUV
If1krxOUAmhJTole+WzF5g9MDvPhGEn1uyKZaa3EyqMf5z1iWdJlYkJGxe+29bPe
RL5hCGD6R/EH2B61ljBELpAZF/K/5RfASAZ2ZarkW1JccLNRtIu9fXP7lwq+pnj9
G1/4b1FqeWwoEgg1xZmWfO3jMuyN+rw/Xo1LvbwxVOBvaX2cudFYfQE2Sqdv+JJz
QJc8W9Mr2K7BVUkaU3SNpjySBT91MdCrkZMPI8GwDNDqSKai8JvtiBXZSeeGVmFr
4pus4gsyFnstML+IgDrfzMp61cYhnVXZNkYzFD3C3kZ2rPyZDHgSMmllkqThw2OP
caG3S0nKE2iAs/7wXpehxKWZLLmdxB1/Mrpg11RjBUsgBuOTUEc2jPLDBkFBClWj
dyiIvbvmi99bku5TYY/Lvjk1YwcchMGr0rNdRRA3ItQdayQE9NBPxpgDFj7IDuj+
UvQpRoWsCcCXReB4q1iIP5YeSrw9cUNV22v3Ty0EFo8fyzkzoT/eRqDLhFWJOAI8
Vb1tHGsV3niBnSurW/8p3COeO+U8Hp587/jnuozJ4NfCwtmSxUEE0wWD6joZ+Ra/
s8W+bE5Bb53ZjsNjqRaJYRz7hVh7BDqmCf3b4Do43AN8HFZAmeaBDo25pedYYt0w
e8Ddis+MMnkQM8tBsXniIM/vglnNtj1KqZPbj8KgbJCN8+20LDm6wJDyrV0ii1Ot
dMipaLuUNaf2He8TDxLrHp04PPzW2EagGUTSnLYmVoQ0OqZ8Iv0rHpx+Yt1MIEQv
P2z6GuB7V60iQiRQMOGnIiorkH/jFb2YuOlZBGiZQCxsZHTAT8/l/evw+wtJQYmG
odhhWJmbr++LLMIpsyq3q8fnXqidOCzn6cWZs0qbBAv3EXJzVo+U/fsigymObMeK
DTsZLiVKkvn36qfqGo1Xf6m1xEhzB1P4w4+E//UotnWTthGg29vJY1rAhOxMk33P
8Zjl+KTDEuOfhSrYgmrwBOf88S5jHTyWN3Fw3eJ/B0n62p2nT6zP7oXNcWyA9zU/
CnoVjUSelMUutVTC6Ikj3qOWHGyLU09OKCfVh/F8APd+aAxaV5JgK2rD30XnuOH0
PJl5xdw/M1NUb8Rhk5RfGPmO90F7VeioJbM7FE6bNhOAB7dsRw9xEOdMAL8YG3fg
a0EV/xH1Cw0prCPfeFoJQGP5eTngeTUWWzlvcb+cdFO0bJY6V4FzxofeLrx7j99G
4dmiznNjMwq16i2EJBdNoAftIobXHj0C4WPkBnSrSnokNY73UcM8dyjYtPg/DWY8
ubv9ujNa6dN0CeNzXRsBG9/2/zKwn/QSMZlAHoRvIUX6dXxrYd583e9Ul0rzcGf4
5wKo664W+HsyYvGLDB4O6q7hoTsYwFWEfkAQqQ6H2tz4SikSPyaj3wUNvoyLL5d+
rsUFJqgxNqj12Z7j/G7Zmt/LVHJTgah1rLS1Y8rAznLFg2XEmvnZuwknt9VqNw5S
YekequCzNr4tw7YbI5Mpay+cTh7z8aN2ZNhzAWAwraCoBvCagQ1VGu3fpTviFQ/w
XtKtPOMwBMaQ6VWd1MiGWaMWzUEJ5J9c/i/4AAbirWX3MqwUMicRpAgwAhFMgtFD
kOhkEAp4SJSXgJZc4JZLUVIGWXTRWJKDo0QfdDifNJdvfbhzsJlNtG6CcirTd+fz
4NQpXl6bLF6197Fmd8ibE2ysQ5ydZJPWJ7bp2OXyipV8HZK+ZJF6KDefPuQLqdf6
/8rkppvnO5Yvi+6fg6jqB4GZfaTKOyh8fyfvbF8NoYUwfAsHOuksdCWHcjG7Mspp
mXkftqv1nnX6ypUjvCd0r3ZDWb/GW7knkwCj0Z+0juziDBivrkn+zWTEDEwa+I+S
SWbZLhnb+vzNKVOTBWbPz9KcNYDaRdJNjwRHEzVs6mEVUjGvmnu6U5wX2ndaK9TS
uLBOgOE+Bp9JzF8/oGUPYOYQNamZjb9S52PzPUHZYbMYy9LUzOw/yCW6QcrqQKQG
mjc4j6YHGQtndqKEOG4X+7iyYeCxSvfGNXgCChrYPzfvl2WmqyNDa6a2rHV34VbB
dE5+9isbhUSOKWu7Ig18BDtqN9DH01FKXhWfO7/ttHY0TrE911m5VXMf1cewbtj0
xrsGSITlqwSQvK7PfL9UlC6XbTz24AKbegzuqf7R5acdDm5XNeqshDPjYiUMgvAg
73HoLUjoIZK0jXB3aSV37aQIVpbEve9aK4Gx0B6NVDytSi3AeW3YMdEiLMytLVEr
0yQtGkWq3yTNzm/kEL5TjBVVAvoRQ31BsTlvXpoG31mtxH5SXto2JvnpySo1uccC
g5vAEE2ss36ck9CeUHYb3/dwi9N2hDaBeGHQE+2kpnq1IupOdcb/IBLFjNoXJPQq
HWcm1f2GZPoE9bWoTlaQknadmUK4bdJ/e5lWNav6r66FYE2bDU01OmZmhoFXlW5z
LHlkNpX/pAcbq1MC9KiaJu5b3YkZnC78jD5xL7FfKP06azKfmeqvp2Aq5p5LmusZ
151faTHN+ms3yfyfQPcqyXGBQ1Tmsow8vsxoNqZjqtiy1O56JjiYKap/JrPmGwsE
4rJgTZavlipdiDBt7eaB0Z7uGEV0T5cZvsXcZIPAQZ9Urc8XK6+qBVAkH6lKoDI1
jUW/ZdO0VmQrjW7M/hwHBjXwEHHCCinSL4XoWAB2TGW9/Wb98cCy2SQYemPv4ge4
4jMvskaoBxl1Bm7rEQzwA5F03e8dkxLFFzLm/n5X8gIuWiU+kkKyVi1/fpNg4AWb
1zD2AQ0uvfa1vh2ZOinq57SDWKkR93hvKfwShiUSgiZ+xOOFdWHR8Xf/C4RP6pOa
scCFN5KAeWSENxU0GkRX7V6+7Ya690pPW7zHhNUU1jRdoOzhFKz9nb1ffAUdD8rD
y3p0CsOnE/58SRFsEYVCosHXN+qtus498lwS+8bkOgi0oxP+ZTQnT7K5S1UUjpER
0AI1/529zCNHyYxV+/F+B+1wTkfzNbkNruq+oEdrW6P+BjgbAxMlmdtZQk9i4qOK
Cua1FH1a1bxSHcqtxmjcwa3fayZ9jpDw4do5bfHRadvCPGlSiKSxDgWlnGXLBq0J
y72B5I5NR9qnN1RIoikjhnMBk2FOo4ycFoFJjbKgmf0pZfFSd2H6MF73F/Y7dTim
9+HFQJKt7Oy0eArroD57nFQcgdGzSunsX2JAmKFhSitNlEqJiCClUaNpY/g5MsJ6
MOYWtmjYp8enGvpHGN+Az18rKUr33MvQH0MqDwcn1iU5OHFEhtqAvvtE/Z+caZfQ
facSJMk3IdXZ6laB3amdYmYjehdx4RoUmtAR3VRR1xtFITpcg4xmGUF7MgRxM5Ik
EvrbPRV3GI5rLnuhXkTEkvRuW3pidPQBG/w8KWVQg5ygOJDQWPBgfYUjetghnwo4
9L0aYwSVEWAxQalmKhUdigSuSvqv2DTFYooskYPOs1vgSq9dLyviFGBrGMF9vJTh
tNyLfeGvlLujNgSffz9aS9Y+wHIFIH54wD2tkfGjjXOzB3FRMVSpxeh+9SyxRkKS
3gmW/mMl7z6lB7n5xSryU2pR4/iukK7rdZfhtqICJjEr4Qy9xWdskP2/C7GefH/n
fo+D4YEOgow71V3+r7JCr4OPjT2hPR/2Nj99nbmWiQJDvRpddq2fh4WaX5k0rNA8
xGZNo4yLszy0U/W+e4DQR3DALFNFzZX5+A3q9NEfTaD+5EFnLl20sd43SxwHWMTb
rXV8wfbKeN1HnZVW28rlhhIN/9D+9ij6PeuvrgI7Nsv3irc8qex+maZ8zxDrnx5/
Fx32yjKWtCJJOr0ddSdliK8jjxz9hAOsPrRWtLYvKfcXNrVmwAeziKu17XXtVhf9
3EbONciq6zfHxw3o44HnzMI4atR4NQ01jHUX87owX+wNkr8n8iopDypdiKeN8sgj
9rhSkCn9t/clVo3zGRKuE9uMXxDlXLCfYtIsNGNeTukOcNH/cMFroiOeS9fu8ILj
ckRQDUn37mhSVetxtYLGNf8xDpcskW3XfasOE6g2ChsCrebyRecE414UktQZRtEV
4EycPigYRqEEcck3MxXIy4vGaWLIWcoSuZnyVv9MtCNeb37duaafoMTcWwgsdwrC
2pedmzKVqmQ95SKbm+D62OFSTeVXNaKSAmbZphQJ8ZgelvMZ8dr9QPYhMUNDGXf+
Z4anV1MC/iovE9eSd7PWaJizct+BMjjLUBevEO0ZYvpDlqBzmcPozC/epEMGL7Eh
tT8Mugy20C+CLPyJjMwDYBluGmc4ezSruhHIzAvTgTZRLbOkQN9Yw7jDSvBAzjFu
YSNOHLXT/85KdtCn6MK3PgXrxHlM0HGTleBn+/VdnAiTo5wFnmnv6sWsLRljIV8Y
0KLs9DDSBucJVh75pNLT3fOfricgVd+yzKvx6ZyjvxG3k2SY0Qy+d2/NT+uh9/Nc
ewJEDuMec24CcLwoa2OoOLHcqgXh60bkLcxc+UUvCtb6gRbivBjSb4Fz79zXySZC
9PINebZtIA8XPwNdP38HvMlMjGK5niBPQkv0CjXqnZn33juf4KmWjzXxr2j/1h48
pJhiNPtOiZUMhYvQDKQQ0WvDsWr9Et6AQHpFaEfA5yWKsMvGlKMmHo3QbX55SsmR
IOsHsxgTr97ffgPeJZ8BX6MQ+E4ipnHSxBzhovzj4kRTktI9TdZ78ooLXPMSu85T
B09Nc3PGiXltyvKkBGKe1Dz2pgsUyWs2bKiVJGo4PegJb4Q0UmGHpd5Tg8OBq0ht
+SJQKLq4po4wq3wyD+c8DFsio+3FX+vOQOKuiG0pGC6oJUfTI5ZMBWJq3vnAAGe/
4qDOK2/EvrB3D0dmCpwXSx0lIEhiLB8cS+o/rw0YmEj293aDEQMXEcQ6PRd57oup
revGHr3C5aEdFW0lYHnlF4Fweu99pH795EF1SZvVK7e9fQjTkru2V51e2BnaMDXJ
jCEvjLCDhOuyTJHWyF8AvnQMn0EBIoovVm0H0bqtTUpm5mdcBDgVX+uFIR/aOv+C
+wAdGJ+f3GzB8zxeBZoApJDU5n/NKBHOcv+mfd1FdCv12jszO31Yq0BeQpvtw9tn
9ySqc2sg3aeMQzBSNf4acg3xpcPkhw0N08kvoElIRm4m19datNk/ve0Ym6hUVngF
kOhPUHcSNg5wBEMIhhK3+ELw5oDIcWGPVJU0POht9gh3SpJmE8KnWo6mc9MlnVRJ
RqA2sOt6mfHIgxt14RPjpTjjrVRGLdt4j4H3/xioq5GGTOOVpggIHd4v8pcG9KBP
/ppoY5/A9HU1wb51Z8uvrJw1D+yz2+Hn3SmJBcaCokEYgz1dKVqnp7iJtB8r53xY
V/ljQmSUGkAm95vk8oXFVhJ6mUtOzAwF/4X6lTkB329/mwGdDc8bwH+vJYSYxdl/
wGC9BgM8aupNtKbWc+c5m70xKvxSRvDjp46RXspx7TOUMo+v1GJyfkzDlvOe8cWC
SYFS6ugQDMioqdnPa8cHnckEIxC3rbgNiVS+Zg0cplqI5cWlsRJRwTZyr4Q4J10m
Yot1OCVqBtyoPvy2N88kt/z3YXgxLB9qqHiJEzE4CCmU1qR18Bdi11CqHtjCAxFb
GP8hPlb4T7Z1TX8hmIiijFMw7NfJdEhWrXnqP/OR+XRgavXUW0xdi80zdCrmQBZ7
aohLuh3RSqb1euLKF8aF05hxkzh7QiLwnIND84/j36uuDUJk+dqtoj4yRHtQr4Z5
3/6zvjlItYXG6VujiMY02mGwfNmbDSQuClcg0taidBL+PpQIMrX42qybk38AxtU9
20HHd1r+PoDTUkwPVEBgvfSIwLWnSq/hybKWXA5ECMZdJhvVNntEROz608A/o7Ed
/9DEQ34n537EpcNwKxDZgxrg+vtWV17aZYTim6GEQRIYkLHXs6qGZ/vExOV3kFDv
UYJnqs7v/yHzIblHWiOKp2y3IjSAHngnexCP4iHhT8g4GH8HBOFIWL0Q/pDi0G4s
UXJ0ZM0K3gAUhFeN81eSvifuUUHmOK7MZVEdvhIJwOkgJT3ZIsp9dW3m19iYmZc+
ZcJN01GihuV5RLszyJVg2Vqn6bATVH64OKSMijl1dH1favIgOot2hOiB0jHKc//H
hTuJKgFHbFPLCf4XxagPRP3l13uIiNGGhKLWEGxHOhSSthZ1BYQKGa0nJSfq0htu
e0T1nZw3UfJD/GFPKwo7mpNT5YGxpVQ9AHV0Rgmebz1a8/Agi3GoI1DIv/IFRa+G
3yTsbBZBC05Zowa0z63PuP8m9HiNe6MXbA2vTu3BMdJTIkpuB4bgTVirB0aH7wF9
1ziaPxkLekHxKXg3ktKB2Q2MF5QoS5MfWIVpjqHx/TjbR1ATcGFkWVBIi5vhrkXH
lBchbNrv5zLi+20aowXZeCQDBzae40oq2uIWcY0EM9NFSYnU7AZImZqq8CbZhAXG
fpFvq3agBjhnGD2sDQvSFp5puEuvheqXjT8eaRDi3lWCKct0xLkldDt/3M3paSGa
k+p28WfedvrdA2QHpE9cHrsR9UxvO3B6HFhalx1HySQ6YOCl4rEPPrVaDHxhBD4O
HEwhwKYLYMJftB4ri9iNyULbJEVdtdpNH1QZX38b8KY6smmyF89L4cjYpyE8JiMK
xNwIT/f4/2BBHkOANi5P/XOHNgHTVO9K16bHzcqvcrwxPadmlVKUwJoDco+hjx0/
43otMtDqmZJF3fkJbnZ58d91jp91BhBkJrkVv1ZbFPIXR3cSM+kWFa1DrGn8xbRC
SusSFnmfpvDfHxp9oT1s6EYdjoagmiGT9ZLBvAlN3ea8Em9kB/OxPVrpWjRNerxS
lVzqSGnWi0d/UtPT9KEAwGlyBjXQCTA+26tTu7El5XjUevVOqyKJmpBoQoZcD/Ky
FMecVA76I9OIYMHfXSKYX7HFz8rx1ypbY83V/3G/fvjqvSTCDi784YInUpZ2aQDM
YJ3yfyOSW/uEc7b3ezy84KbqP+Borowjy3o6mwuvedLxM/qXF/rnOc9bDUMFntCh
z/uqbQjPIAcHnjm4xZPqOkAdfIQ7mBZP+4lOgGNIJznBJ9ob65Z1pA1on/lBUg9l
Xjd/vx1s1WGqo9oAhHbg4wM6YD1ZG3hHQ9dpTCBbJanyIfwxfRoPTsNy7c1jNBmv
+JR+gCuzO484LClaASeFyG2Z35DxrZqfGR932AG3LtX3jRCFhbhgHUX5rZdiAFVC
nZV7w87nLSMV08ImLEJ2DoT1csRaG02VLyHF4njknhDaRrmU/Y995h9m/EkqpBH9
uN6+1QyK+4H5YsiwgCFGcr5/ON1nvSCP+HQjL+e/e9RJb+v7B62mzalaenFUhp7c
wYjb5WJnzy9oiUwS9U4Nl7gWTabHXwuwgLatMpIlPXqtsz+puA2VJ1CP93cddQhT
D39RjzHksg0HA8xrXAIA+Uriljq8eWZ4dYa8gIGz+lJiP0TzDEJ2ZS7AocwCJHQy
lIiSp2epzW18c1bOg9QPoD2k+2lsa0ZEIkjgYCp6LqA7hBdvfy0wcV4AxocsJYCE
QGpEWYRkGcdf2SrZvInzyDJqBv9nRPpdqOZdGsfglJNdKmLyU/F6/WVFJWtDZHxd
YRW8LexdZZL6K684an5220S/qWF5Cosx7vqw/tr6QU/qIaHXdkWlIsZwbpy5sFPY
9U9iIpcueqIMh6ZGkILHhtbprSNlj0/D00JW+vOVXx2ytBOdvxHDfhy2ZLacTNwh
GO2htaGYmXN5BGNhfdpUEZqyz+OLCgTtj5O4YOBmRH41tQfznX1sTSIbGJ0v7c3I
V1TnaljWixdmKcqeDlUQZRVQEEp5PC2BvIS6SuBXar1Rg3ofoyo9Niygn2A5tM1I
G8A+l2ENqYYPyiuCJ+2EKc27uWzr5e3unfU7hfdgf6GYb5G2vepHkWhCmPIHAiYZ
0VxCOSNj+efbjA6rW2FzSsnL9132xJLq93XQ+ORMAHdvuQ7/CBPGqQMFHKoqqXw+
r0YlzO5Hop0dhH4VFFvfCG8aq4NjVasVM94dhUpY23LEnYWy0laLwWtKchaD2a8K
tgpLnSf8aqVshp4NxZrSiqRCrkEC7eZ9jc7BNIgenALwo0YNw9As3QrdIJu8eVj9
I7iJIXAb2b4lngp8gK00sZjTXcDhWWlhKPoRmHGSQ0l6+dEoANti2eGPv6QmtmuY
Ls8yGCn5ArJ6N/0kj9vtwm5nEjh7pELLkELTWp+zi48bBK2N3TGHohnSYJqSzi6X
K/Ll1HuRx/1/JydtiWO0/Q5hgpRalRuuPjbamjizMtJbMkrjLhpSUp+3Q3V/R2QZ
hM1RSfoS+k5OuuW0NEa+n4z5Zs4XOqWBINq/pfuGzKapNkNmXZlLhBhfUoCP+mUJ
A+W1DziW/zujChZjinW71ELETE0NSLBZrsyqxoCNs2JnEf0dQo4wTfnLDgfxW27V
fOhrosSM23PW7x/P09C6Pl9imUhCGhOM4DNLlKOU1OUpF3bdgi2RoLQrZ5SkMZb4
zfwtBYFetHiWc2deBR6je2cq53mJTwPbSzK6ajPsluLl6PvwtAoFnuyznBR8HSmx
gkmTBqZB9nSkwD+NM650yHrGsd+WvHXizcHc/vMqSn7HKtq9TrWR1P5DJgusXGt4
CZoIbGJZ70QzX5/rNZmLGY7hkxF7IL/dwdB+YeugZI3+J7A+GHAHscUt6W6CwnRd
SpvXu0lgMH0ibmCBCtYhgyXk4PYSt/xK/Ag0M4+85VmaVnB+cHRLaz3SAGT5tYoX
C28df8oGmTUTRMIGfZba8yXFOIeyEscHhuvrg5kfFtntSHSVC6k3bgzx6iVrAhhX
Ur8EVJYhvf/OR+v9yb0T4aft07a91XQKrLT/sW/uthxXJI1GhS4Fe+WzfjADe/NN
er/VcER9M3minD3lAS6kNUH4qXMcOh2TWXdLFQ1ZTzxazJoom8z83z20KpgeY6X3
qs75rgGZWjDeDa+B4Ffz7lBR0nvzjf5EQ6C6Aqt1f+Uq+0mJ/ghUyoeHGGoTmLEq
NuUE+9DKIvybA/YrKP8Ty4jF3Y2BzVjgmy1Dcwcop38TMNjYgVe9RvQ9sMoHJy5j
NTN9TZFxpemn7ePsuyhTpnDZbRzmn1UCpT7KulK7IMcVApQWODBF7Mu4OzeCqd1A
WIb6njwCyYRJdb9J6xmlx2/xXTVRxr7vYEuo97OAgfCvtQszbvri+M2jHosCmZya
FjsSQ00AS9yhs60zc6VS2793u4YDoCk8wlAtwt1c3ttPFgfOhVYkCY6diliYY99c
Pjcg+KVYzATaAPOX5OQzj+xG/NG6d0P5MFwUDUc6o1rOviHqOfLSxoS2mEs88IwH
tfen2Z25YTtRNvMOc7pbJwyQp5IIVMKnhQaH7mvWd+EbZ7EyoRrikZ02ZQom2Xjz
hizcmtS19jYyPUcAqRhOxqJSzfnDjUV6VAzPLRPx66+5spm3K3pczLDUp9NPsKkR
OHIzyhEMo95yKnsJ/m+e+fdmb82wvcTL9yA0guBE/BS72Frm8UxTwICdFLIpQ0N8
tju3YD4NsTZAaQtVIdVkVtV01cythpvhh4eovYuZq3IG2T6B3ihOgdGI36ncJJWV
akoGfSwsbhecRbzqPw4Ax6WHsEw16BzSvVDOi60RHxbvQ12fZo/Gq1QVqGUqUGMm
DlIeF/sHjBodX3DLHCKNYZw1O9rACWFLw7ReBjEcf/Gx80+ncfzcTUV/8yPAEWKy
y6PNWp+JAsYkhZOgF1Ix7DzWY8or7gok4fUxamucCmlnXoPZvkV5+oyP0ibIn8OP
WqGKdOpumoLvdVHkC8GIbDE/tdQrMiCwxAGU1Qp4HFFdRhIHAQlkuprEuNJ85aRw
/z8snle5DGBga8HO30yadwuDT2eWS8P4ugvlqRkFKrMl242mtSYDek2uDh6UsJP0
r+r55hXNxKho334FMnlMS30pfAIaVh82nLGzzAbGFOfeTq9avXG8sMUaTZySC9Y0
pZ8BDiDwEzMlikAe4Mc0vRP5FVRNXtQVOxryqrk7QNPyNOLxidjaGYl6Jj+jS1yc
1qSl4ZLq8ObWbszswxuB/Cu00rOo0DyXRDtqSHyx3UVNdoclTQH0hqPGETcCaDtu
hNVoNNIbxy/I/fetHwHsRZEWluF04sKHcjQbfpu+na7jmlByUgxfJ8AneaMPmaA9
Obt5KwpIQRLoq1SaJ1KtyK8kA7CV0SBofS+x3WG3CZj7NII02A4apum5dPTP5aHl
y9U2jG55e5tdWBubGFVwsa/4CHuNDKJOD4AjA3j268uljS82wBPFBc3s7TxW0g+n
2GNZ95LL6JAqJlTaIQpIjScfLYMay+4dwiAS7xtqnCyyXRuLFmCGQTaxdkNmePxM
RnhGNVlpx9mtF82U/8L/Uc5zjvb4QLGBX9MaIvy9JavxdOaqUHlKlk1Ljycv5M+I
gdRJiULvKKPxAhIyM7nz1Z4RI2iN37pfkqVmoCQOw/dJQbRMK5tNZ9KtJL95QIcd
W7bikfKREbn32UV6ypVff06cZ8In6j5zVuBRer9Hl6+PVVQxUvc6Auzo+zuGBung
hDxPruJySA0CiL9x2/+ol7+bVyJqawrWN3SdAFrYMXOFRG0IiNiMBInI2nHmZnXF
095deq21EI3lGB4Y2babRKnbD9kkgNhLKjN2HRawtgWpTgOhDtECcdT7e/7lS3S3
EHsjh5o/2LL86ut98UOvUAZK6zL/yAsN/Wi9ID+p02wOlOBPu8qZD5fKihKtvWPa
T7cVN0i50TTD3ndBWQxEvMtdPY93Jkm3eQoy72UtTRtozKES3qO6biiTbXGY1Kcq
bDsl9V4jnbToe7535EjQZsPUvNwzxQNZRqh1BXlg2NJ249LkUJRX62eJnN7RVGLy
2vYefjkIjJA3I3JKph74m+okBHLegg8QDCWp9SdiOKKR1P7klQ2xt1F8MN7qymgM
h1+y7b/lTxiBtd5snlCeLaziUSL/qKHwnnchkCQFEHUmZ5vwQZyuj7wfsZPkFWN4
1UoEifbQYY4uSjM8YzuYdMX0zaKnATpJtXnunMnTtjezCREM2k683LdFXyXP8uHf
ptQM4HnLMEoa3H5PfKoeEffR2u38qJ9wNSfUwQZrP1vdChHNMy2nIW+9/Ie+jomt
bQ7D7pKPSqP3xzkA8RAHIWAoqAeuNhLGUjOkFYSZ8S4OdJ90AhNpVf+z/0kHpdiI
bnwK4ty2eqhikq46AI9mvEQjpKBpV2NUfpIhk2NeLVpY+HLfUXZbDYD5HYkSE6PS
Alnd9a3uj/gFRUC2kNMzlQb2yDCWzra7q0v2eHCkQR+CDTDTWDjZb9UboApHU/ia
PEqzNQc3XBhO+83t1B1pZvzASbzeqB60tuZPI90KA4dfTX8O5b0OBajg/MROTHh5
QjPQmzeDVxFRLzWu+/7fksnTuBEMg+8zOJzDxx4VP2fnfIED3mz7I+7WI71w3xp2
PgF8MgPwu8qBLsaJsCqnNmnoTUj7Tijte6+dZS1RzA06uE/wbRc4CCYzH0gzyb5A
gCTpW65iOlZZHhgPp3SkSHs6tEssZKkqBIQ4X9ZSThCLjjup8rynEZwGhkPtAPkE
vXGQ07k4wVO6zxZsEO8NkqsWjK+0uuAaEkEYLYpmr9h0SzX62bAgyKsPmF4NtpX9
9haneEV3wZmnrN+5nzCshhSp1MC0v3cHgFVs5Pxc0OLo0sciNn6kvJIa5fl80YRN
JuULhhSBbv6QZ+vyie89orka+ngSevdVaUwP+i4VhmnbP6xbxtHNYpad9ID4OX22
w4EegwJJg9RNoszCzG5cr5I6o42SsX0wRQgWw9AXrinND3x+XPAoLYsC8q70ewu/
HvBfVpldImxwgqmm3/CDI/yMFLdFmhfNPTku/HLr8iAmbqzXOP0e4xqIMau+LcGK
FpdqtKcpdH96/uXq/0QyOM9/VVZHbZMdRYLiTEPKn5OQXD22aslWupH/zEKEAs21
W8B2sasUf36+SlyQ5+QrxTYYcNc7nCNPBDSrsCj/yHtD6Flo1I1rWyVwtodlbFrO
E6vRGv/35etSa1zVGsAwTaZ+WGuE47n3DI1lP/qu2mShrLn83RtO5q5jdEFjHyqY
OyfRSrmkA1kDYzxiK0qKNsWoDfez/gs82vfeVSMZh34YZUUp4jQHDBdutrojXPdB
er9Varef8RKTtTcLqCeVQtJmEwZZjjmolcTUKX5jMHcDaIAuC06LVU/6ziGvJDJW
jpfcR1l6LcJu4VS6id7VJcIoF9jK759dH2DBzu7qzMOP8/UB102zqk7Xi8Jlr0yJ
zGkaPrgfvB68ZfcrzENbt4PzTppMHquY16dg2sO3ULpHUIopqm28p+LIujrtv9sN
IgvOTuRfT+h09QcYrwhOSKVO7/7PxUGybLNVGQm+5ra1dlOfj9k7/NaEjqDwatma
QEb60r46UxqbefZi4wOQPSSS9FMmTTrA66OFao1zLexrPW0NYkyRSgsuMTmRfknW
qg6NBsEOteZpqA8AZKzOYvheXpncvVcINuuOHGjOvtY63T0dtBol4cIipHkkBngG
f0WyQDxuAGizYhWhSCWbd7a27FjJeyTnbvrUYyPfO4Fc3RcwUQj3TPjPBapoP3Am
AmADVAZeTRImoFLD2zzTyRxT5M3F/QVFmnGytN0NqNNMzQdLqwYSKVit2HdMiuR9
RRKf5Pf/vW5K16ZGit4fV1qOcK4pMHQgoRmcjjh81qK4gY7Hhz/0VWnrwcsg9PNe
ukYGKD3rSvVxiuPnQTEUUyAkLk2au7qBSIaR1FFTE3wQ3BmPhZvy7sLfLFcyQtD6
dhM1tfcE+3H9em4pwFtd/ZTkhcrXZNOJ7sNY1Xwpn6sWcAbrR7Eh2c1OaRnBS78v
eva2ZuPUUVSLgBCrAEuJOTBFacNgtQPJ/1zOPSVv1ANhfqzWzt3TATOOgKoQWxBn
kr0fgX9TTJChazhogOlcA+2PfTwQviVH8pVZqg7Dq/YN+qy5PFW55Dp/oLy30mc/
bxvKEGD0DIDIbN2yxegH3Su+QIRhrW2vBp3FsE3F3u/RRCrw1AykrIfMs7QhSpDn
NgaI461gremH4Q+J2mA54JOGhkprk3beeHb+64N1fGP56OwVGociAZ7/Stgy0y1V
B01eK1uubi0aX6rHG7QdOChDZOZkfBD5Kq12IDzuMQhqTnoVYcC0b8+meH+tCKBQ
d2+J/U0WuUDPS21DGb+QSlMdDubyWjQ1KQhqiplRKgcLIFKTWFZT9ohVtyaePZeF
F1QswNLISLkZhLmOzGYWdx/LMUgcr0o8urhNF8Q7j0csmk5+v38wCUmCcBVEt7Pl
mVdxNVvi0TcQVf/0DPFz39ts1rXCO3vHF08BueRlGJJzIazEhAm7FH2uu1HBLIZ+
cKVDu0Drv/yLcLE4VSNIARvlp85I7qjAy/4s3YLVdgF1U7lwadNkT3v1m7/QC36N
HzVb4aOV3vvkSnzypHKcVUlzmGSy5Zg8FYYBbX4pM/FABD2j0hYoAVgFJcicpjh2
wXOG29wehpH3fLA2It69bBUnlRnRxiFQn/vL6CjlLgci3QKJzh+dTLzTiN2twFML
qAFML3tiKokRPvzBipzBKk+3ZSV9Nt7a9YArw81oqHPg8ucgeV+89d5V7VA/nGOc
uQRikq+NN8120qZ3UtEsPsMmN6FM7w1ddBDn4Mt7zih8lmyI8RE6A5ihl9zXLY8r
TrC7zE4UnCbK4yDMEWIeTtbmdkmMaMqXybtxOFgtcsMv0PKRdmo0VNNgCAAZ9l22
i00rkU3uHXElSoM96c9HT7RW2ZC0893FYCCkg4pY8RsUwJDrdUm7eVbMWHtKhTc9
5iZBGiheUQhBOPEsk3z+jexTJcOBdWUwOXfYaOYJPixzAJhwQYlj5MEdreIN4EiF
lzo5mut76jgd+iiU3SiH/cawbdgs0BVFbgTVano4jclWjzNQ5KTr65mlSEAsQimx
sxUIyaKOmbDofEXBfZ4huhfqoqx6AHbdSpOhpPz1OkYkIwqS4ppXiz+BtrZud4Pd
hyAKMQLrLHhWj/lbWDbPh7xbw3I07Y52sCCdrOR7x2/dS/PVuKPqDrEQN2O3fc05
9XHl47C3VVw+Ewd8aG5Bz86ywKHTEwXc0jmJn2MfmjNrKypwuXpUPL/3St7lBf3A
bqK8Zxi63K6C7a/HCr3ZxbWVAirKhrlXco0CnEsrhuVtSD2l6YzgzyJqYTiJEgTS
6iWWkbYRnGjbg896pGHeRAHV3/ukpqrtNo3GgbjeE5DvKsTaKIPp88+KQo/1UBTy
P49O9fFgEnS1Cpq1C8phQz7AEzxaS4P7EAWqGzGiZ8yqdr6iU8lUZRTR4tjpw5Fo
itGWquxkeT0JMMn8OkRteQxJSBnGvlL8MtLScwpQ9JsOmPy59cHW67K8j4DkFhJW
vWQBNcF9Ahnf4fI63EJtd7xzVJ0m+nLVvr4xCt8p8SFqa7qCeMIu1SBbGp0r+MIq
eWxTNLgELQhbGxBdRBOv4HOwcKvYQ4xqZCbCCWvJGSE3jNYViMm3ol+9jagQD/tz
cu5qjEXbyKsAuHApHowOsSwvsQQddyWTeScyXNKZTPgbEkPfsgS95aTy+03jjTDx
EgCZGQ+nSdBVYBwQFUForasYHJ6ToHgf1DH0wZD7wgmGa+mi77VHcc/GRnd7IOW9
SHQTwoVhScTM+aOMDnO4L6qzeO7VIkLT5rhS4ahRVrtzSVA+HZmfw7GM8xpawf25
1qVLE+PzxrtHMGXMxULM+wioagiTj1XmvDEH9OPlbpWQmoXk4uJ2EczUrDKooBR5
kInHRRnYeYeOmOzQ00L/I6rwdZfvDxFR7PhD7Pjl46GJlJbBTofyIZ4hPLtCQXMF
nUV72NQo3G3vL91N2WUP38UX0Kv+OtdPfCPMn7wBWBtfQ+4dtK26cCd0U7/lnnol
2UI1alKBi/dGc2C6zVEeLZ1QNBgrhuf/pNTzOE/OVPLDg3uKPGoDQTK6EjnMGDwl
FMTteqNu3MMBUPX0hbjBNruCZWXGo2grRqA/cq7I3lJmh9Z/lFiJ9zi4GBm4JAjg
DCoeEaV+T5HZz7L4qClyr4r9TnteBMg6JxZzgCkgQCvNyMLmsrK+gbhqeMOVdCx5
Tljnz6fSXgVZws/+yOvPJcrXwnUmmh6GBb9bIzW0i3VXq+gCVG5xRnfGmfZN9khQ
3CA2yHJyHmYo0Cl5xPrB4+aOtsx1MB/P8aTX6OXurJdsN3pPWuJJmLIj+91ojPi0
bC0ou6L3CqlU6S7UZAmXhn+y5n2dPQgR+qrt9mB7Bp8epfBhMAh7EG17+8a2s2e0
5YRjYjSlOJsAu5q4cEZd/iPw6ZOUYAM0RzTUeywEh3feupDrKe81d+W2SqvX2wYm
QhHDfr2PsESPYpXpS0gKs2iQH+sX/WO4fsz/h28cP54BaCcVqi5moB9kcs/eRygs
00AXovtRibN4tNPRMZwzk7Ls2EhcgEx9FlwVRaPTMKUxqkTzhmjgVItqyIRaVazD
mb0hQnRAuUrgBBNWCh9hedbvJ+XG+jUAEo/xYRze81mS6ZkUYyF2a6rmJYqgJ9NN
I/1M9FvHLjNPjSa6Zd/uktWBX4jnIUIn/ZYb3r/aMToX+tdUxYeZ6tEOq19LhNRK
rLrhGuCBDxUgWpLdruycj0MX6EC+P4VqR3ScMWg8wXsZXeyYMkywIq3TihrzzZHR
RREZ7jr1nyDqbACSmEBendNFyat/kHiuSYSKIVztKUg1FS/tieDa9tlRmGsjoZJx
alAPdkagJeVyUb4mpQllkIdb0Iyh62D3i8rR6KPFbbd6vbzXkpWLLn8lOP2xK9k+
1wkySwHAGngZjaPVC9ikcDdthH4rr3KpalcPn8ZkVWX91gFeqWOcSvHatxBXRNG9
tSsGuC7CmdwFUsJrgEXgpsBPD7jxLuExze9b/CeauGyiRlN23g7f1Mz4UzDC5Ene
aCdHHCphUAFTJvndhlSur5gMFu0EQhJT2fT0nVXWqSkaNjyNLBPkVzfkhz6wJEF3
/YUg8QuPW8k3Lsp1oQ7pMlPHMfa2GTrWg/Ylnzp0H4h4QgiL9CkkwJ9FtN0xQhEC
Gi4kEoSNCBtwjgfg500gGX2aUOwFifF304ifP31zGzwm7Kibs0eQDlj3YNcrQiJ2
hxQr7zL/u4Q8AV/Ttm/4+rAq21BtSFNaN4mT4LVeb6ngBeNIoXMg5dPmgaVHwVww
qiBmtFfutuXsD+TqawPRXGOvH3YIOWFti7rceXPt5nvnp0EOwDOvxXF7gy3+auGW
JWC0SDWTteOF1132n9GUpI0ehfhDx7Hy6D1Z12p0Lj3RLqcuo40P4HCRhYfHcOHv
yyl9Zh5gHFqf3a8H7yVFy3fEaeWIZmCMXAElWw5sXTR8VOmHZ087z/HKVl8yYEA4
FTp9SD9vSp8VKuynQ2buBUjflO73ZbzwuzPy3wyfyxnIu/tUrEGrTGdWxGLB/cYF
BB3ycks3SdOFzTTJZ6gIkxbXAkXXDu7qQNFBzsNJ31XgwSP2JdBjf6MtGC/862Df
WGyZTW5RKsBde0Pm0ooioamhK8FDwNm+EEeZAIIKs+zsUBRoCpLkZf+NnBLdb2vx
5hOyDYdZb441Fd/1OhYbi5OXwBpULT7EZh+n4vDkSsPPSPQx9RLDVabVnAJcXZDz
t5zgyXf3TAHDktFhkURRsLTTkCARQzK8vNMjVmJ5iBhCc0/AuLlbnm3riAjLlEDr
bCFHASQVsGeotZvS3Jn6qRzETCuq28hcyqnJB2FRYoB7cyTPauWUvLYNz5tjdw24
B8wFCWq2/E9lMoqgJMrHwy3iIPBFmHfcdKoL7XEqhNaDOmFJeX5416Rh5XgNvc1H
R15bd6OhPTLACMNF5ygVrNQYySG1GcdNV/woQkV2VRdkzSVT4k1sGY+PTNjUyLpA
Cso2MQZrWdvkerDnieefwFAsH1zwGsN3m9NSmymVM9qPPQXyMZ1DakOiD/BiFV3j
fip5Kvd6zBJ/KOkG10d44kWTqukm4zZX6iv5q9rTrto95flImuoOFwzQXak/cbwh
RkjAMcgDWvhk0Azs5cqta8Gi7feeKPClpb07VjKXUO5GT+rS487Ujz3jtPV8gxlu
mS56tvLRFPRjuKDvR6klDF1cpUYdKNwkkRVczbraNf2AzDcUpZmWhXaoSdjH5fU+
idrhlRy/jgeD20CR+oqQuQ2+MuIxxC0w9lGiRMlXmLMGLrJVyH63VnPK7l6x/c83
qcLh+JNHcwkOYfo4eWWQ8OqaIIkOnbNKxgL5z9DG3RYqgqMOWlVhIEQnktsJlzC0
WI9SKdoE1ePpkKOIRkhu0ZCQYwoD7col8hwPnnLNSlcAo+c/WpxDEuKeheYMbQLO
eYE+HhkN2gud3yiwqUKkX0N6EyblIJieQoMMERsa0LSJD2BWIGsxtswUW2Fh4dKk
yhGfsfGsXsSCqeHXA2dlXIG3PCKVjYOgDUI/giRTYJBR1BLVTZPvUEeQEeC0m3HC
jKd94ZcepujA9FFWZ0X53rXlfPwqQyZ6b0jdoR90QabIP9mMCPmAzBtJsObuu561
bjCYtem7meoBCDGujNXO95sC1oeknJNfzboBXO7WRqmwSsE84tmybRCEnOf0K26W
UKt9mmfbnVOT5pYUYNhLJOIFICsyn84z1dIip7FOjFH5jAzK9oXHhGlgk0xaReZY
2BhYmfWS0TGF0ztxeS7F3EazppEqialmu78VbLR6iqoLIDG9ZydAvr8H/Ufd3ltB
WQVXgMxitwU6OdVa3q7XinXvkyEwcJcUk63qdPcn21eiwTMmd2Fy/KJnUtk/AL8W
0Uceb3mKBs01KTtxTv0NVh9I2TwkQKtdRWBXnc8zVlEYdlzFytTPbKYqjNWe7jSZ
kVs9Lw3NJK9navX75KimNW961BJ8BlrRZjqmEJIdmS+Z+g10snpdURYH7d5GSJOh
8iqpzGMQpVPHDw6Ay4OFHziPBZZeQRQfBzVqQAZbY3VU/TyKZLkNUaPxuJipKydS
UkL99Mocoe202rg0S25Ymnkh0psO5DcbnACrU1vJPUx2mEA5pM0uXIpnfcGHgYN9
IJAgtu/gXUYBPL7o0PUTYypbwf+e9m0emx+ggmmI7Bh1FSnJsM1UZgbIIYC2mqbD
wf7eASWIpLl3Qfwka0lJWYoc+jGGI3VJyxi8VeY10RxToLg5jkdY3NfgAutVHXsh
dJlzo/A+hSV6y5eVnAOtx/ShZ6YU8xyTCLBw7nUbbBKrwNglzkBG/HONjwvMU/cq
9gnjgyaJQsBpFK4cYJqr4hUkWV7L+oCvb+39h8tNr+2V/cTW+i4dMYdmnsaqzdqj
xXzUEoXxSylwegfsYsFBzGhX3MVaxfLapIXD7dtEUwVnliLSYM91mI/OYRnqIGb8
noNBGN2iw5rCCj2K2auw82DA7gHosec1/nGmJ02E50iRHbMR6pNWgN9M/WiuePwy
fjpnljhn2v7SALJw6Ff8+cOPMH3ZPkhgCDJAs+ndYsezVeQNTHqi7Ye/i2zs5R24
k/D0S9+DSRRixzJjpbeok2kCzviyMQEDghYrzoRrRfqLXJrHvvbsZL4T7/WFLgiG
Y2lj3/GqJZPwq5Um7eSc0uuKqA4shW5BLiprpR65Wo1xjoaKfDgwdpGOo6W1i9ry
VWb3J+/16fZMl23kkvODlIcY47nB43KW8YeuQJBGlPbOHPpiGmYavNwxHKyuaQQb
zL9oT1z8AqV5viqYdvrsKFW5WZvrDo5MCQj8h5vCKZHJjUhdoZHnJIxSwFcDPcho
UFnsXTUg7OeVeT4rPTMhf2IQo3vsped181QJ91iDEmHGG9c23IZ2bf5Ik9vLpv3L
+OPp4dVqeKz4STlCFIuHll81wmf7YvU/q+iAyUNsqtbVudMwYZ4fKEbZZ36y3x0G
jkpdZ9Jntr71tgKoqiBvBNTDd8puBEn8/JcElgLtUI0tskkhtM3Xi/Txte7LiF99
I5EwiznHP0YZ21orA+z90z2nsnWvzaNDcI1L5c7EWCZ6f49CIlsbZ/Irxmt79EH1
Al12flUrvdaE0tW//GuLncYUkHa8rpxWCffbAU2xg/Q/jNG1q3sZXjiawimkPwLa
L5mxCUNvrl1exWRHnRgmM6LYWjX9Ywc3ZxpV3myLg1fvxnBRwWwz7M2euURJ1Ib9
uv/lCLKMcBOuwXizy+66fzjDPRSh/WgguZWmSmsOXR/WBv9lyxnvAWK2RPZDQ0UJ
zBwbfvTVY+DVE7r/+PAtgwy28ioOTLjDmNWGCM1Q/43DoaFTCtiZyt9lCBnxlpFI
NwCH8ef18hP3N3nPexlQva76FjO+mcaK6El2liN2UHbPpaDUtQzbS8zEpi7EPaNA
QpWFI6NQCgaPO3GYiHugJ9gNgGba0fpDpAreWNxDdkWUjjGEQ/mEW+tEVy0KPk1q
yCpLh52tthxqOQHFBvPI1SUTnQm27mH/LniRhDgepcOHVFBDUf9+rlHs4g4mhnpu
9qClI/ig/6aUyu3Ix4lZcGts/zHi3pjHz8XlrDbpFJpHzLCG44y6+RRvmhgx9O3h
iz5tD9AzdQRidAqQVUdS6BB1WqybhkKisgco7RZyQ40jM+5Nrwz/C77hepcCaeOE
PlT1wHWiIol5jzbJQzA/j7Fx0XKRfvW6IcRalwjHwnbZck+VJl6ok0Si5m5P2CCp
j4cv/QRp31wDooWThOJMOE+4y+nqICqJfha0ONghyymLJqIX87GXJo0uryo9GYVr
TbutrpmY407SwsOvl9xtFKPvCbko7sVvEFA3gF27YermI2jOp+PJTskgGkvPnwoD
eMst2ZXMI9B3caA/CuonftqPOOIJsKjohLhD40VPcxHQVMIzWrsI4rcHeEFybyDj
oTa/chwyQ8lAeNGQIgTPuhYlhHdFnWEK9Rd1a616/2Pb8TvpxNAngh791KlQf7gM
IvjXiyCq7ua4iJbhgoqtiLoR2qtLqSoEKl6sJeTwuI8fa//EdpnYVQCGOvPiJ9tk
mGnNz3NJsaf0+3Z+lcTnV3TesCNIXfSZhmYYDKaqvmyHHi7KpnlhwuDO0mxSF58w
p6/xT/MkJplvUyZ+JisMisfEXVNOKxpiwKjqlXrIacLPCm8+sFatL7xhcliW8mTf
kHEtsZLvZPxuRqLsk2xj1IuquccRnE5Uy3Ah0sJwCAcfd32EDr5NL7pnw6hSucmF
L3ySxD1cmOIzscY9PGxQ1jw+3mho5QFRUzXEfq/MmOyIf8XmCScoNW/cvFvVWE33
TygXODDm1rB7TDDwz2ow7QgZ54qUyzrKGbV7knIt5bGzHgXCjWo1W5m2fuwI0xbC
9HWCCirHiLq3+hVCoyb8ZejH2unNnOnMwS+UVgJYoNwVZXTja3nIkx/FDjP4HZ0A
N3yPedQIpQmLcP9bF3KYSqSvX293O6ho1B/Kn2OHvp3mUYQsY1RZkNR979XrPlkA
UpD4zU/ypUONVINhwkFo+zPYs2JZE1Vj5vlQocwRxNzy4SaAt2zir0Waltp9u5M5
n42MzfATme6/0Ru4NTrkjbfQN+1mq6obMigFgalDGtAuAmwQ7DpNdKmWF20AuFp8
DYXm+iS2OwfV9vsU90o4uQZns44HHr8DcTkvTy2XWISfafH0qWTNmbEzv0g0jqsJ
gXd83Ktbb/X1Prj14bY/YeZmVeqOexr/msJkYuKDDjRc4zPocFuC3qRzy/kqeG4w
Grs6Wc4nGg8fLk2jffyspYYKuoj56Ww8Vvb/YcNe41GrQHLi/+vw1SyKbEwLV+Y2
hjpv61tcuO94E9AkbD4vKu3GcC+nnagqdKeDgC0G26n64r3AyeRfCmHJe1IqbvqE
gXEySKHBtb8efr62h3+e/8FSS2fyXtZyCKmHVbH3vRxdFiKg9JPY8wIJi88n+p2c
pop1e6Sq1mBFrlssUUDvYSkGNH9xN45qxjoPiJ8xaozWIE3pHcW9nxq533mN0IBN
50YoJkCnac2QGoFqSeFh0n2tuZ40EwukTwG1hjPRGLYnXuBbre1MkfdEz2kWtJ6l
dN8vion4dTSt+tSyX6bV0VQmPK7fyHE3TInLRB+0ikh+CgtSonYOYPNh1rhjS1Yy
mCAELP/umdZe0bJSCP4SPHhIC8W8KTyRX0lmLj2fNsxifaO944wrhhrpnalH5Avb
8KraBuD1uuTnr+UWbvkQDyNRjjjj74R/2Les1MP4PevMkl7Z5owiQ3DHUjHtwDNq
qMGB7a9pw2Ud1yHaIlXmiKBlxs1iag8ld1qaxi9q6G5ysoKETtAlCPV5sFHdZ5Tj
lFCwvTYSF3p4Q0TKaufR1V/qPi7CQhjzJST8MK6VriTkIhOMyTPyObm+btYguVCn
Y/wpK+EEWefTFBR32uCSs1ujBwKx1FQROcf26ND4zlpXVbplVteyN83jtU34pDW8
MdIigXHXQDj3SB1t61A+HtIC9aGcDIgthmfAwFFYTYCjMBoFv35xqhJ4jz9BKQz/
1GI7WfRlKngRZlyvw6tNgDjfsnrpmVN+llQ4ZFbX9uzybtX+CEZ2+WsvyI9jIZ/a
4Gxu8tEaDthkFQ1fYbwwKoTNh2b3U1df+g82UzySJxdPTKDy2dFnnxyCjtX/1Y7Y
BMplDwj/hPuxpOlxVfg/WQ3VSC/LJ+PABpySmHXw3lP03dGmc8VuG7aqEXtPL/gB
bz6TAcr0YojrF4VfluZTzXquZgTKFywY2r+z0p0pMKLMDUYcPXp/Uje7gcGatfSi
8HzoAfuS+ctkiC0MaskBd7PRc7IDpNiXGzPUW8vrAhiydm7XyqDio6TwogAqJG+o
gQZ9X8MjbadvCJqyhCbCV04BqmeEj1aQv57l3GXeRw68Gq2J7lP2K4gwC5/MWjMG
0iyLuRqU4MyTTd+3BafajQOscMieV97+HVUYHtAU3Ag6tLREEz+FKeksxqDx+Iir
xDU+3pqmT0TSjhSRwaXlUe1TZFHhlg9KXXt6TLzx2QfqhtympdANxCadsAcLzTw2
b4pSUX71CFpumkPIbqePvVDX49BPqibF7THIPMrl9sjWorYn6myxiXPtmmz70GyK
18IRrHM+ZUfh2hbcmMNT0sJV6+WRVLbQPUzc9Ey5//EUH4IqNSjmkYVfrh507Msv
IQ0aLQ+ibqRs3yKWj/M+aqsnChM+VeKkfjqvdLjh+pE6SHqiTxMLrvXdc3kBghSm
96327CrYIlmtUP/W5Xx7tYdhQtHONmO8IqV1h7MeU87b0YRM8IKsYkUjd+6sqlKG
JEEU1apve3ndSz65ulSHfMS+1JcHJfrZ8QMaIaOfsLr+JNUYeuSjaOsPxi9QhASV
MTp/9RHo1QoahYsgQTTzt25MglwbIBeCE9Bzsg0gz/BqayXOEhSfypa3ezO6Jix+
a8+MQUYT+RkbKIE9XVGfGv59Md1/07aCHwDbT7cS+uSif9VO2HZPxB5D4DeXI4SK
k5atWIkw4vAIPy+BOse+U3qpYsjRjl2ZEdxnBIM7ufb/RB72Ot6gA/4fSqlbCpr4
tWmTn+sZaqLliqV2vfnYNOmBoEuZZCIa9sE9UU7S5+kBePsaN8FKN1vKNzh4OepO
Bi5G6ER/l3O3UmQqlTVAt1Bm79q1v9LNBb+PRNQj9JSHERB1SxClABklk5bed+kF
k23aeAFXnMsZUqfVSRvs75yaFzdmpQSXq0P91NgfkIz8y+998Ayl5+AyEI+RdV+a
2x22Zniotk0wnB502NyuWgI8HiCsByUkSPiyH+ZHbvPolIUQr7ZIWPxMj3F7r9u9
tCO4k4e1IhUuUY1kxJTI6syQCaBxTm4SKbTnkv1t0VerRclc4f/79TZe0ae7QFOy
tG2W1LiGTvPnyEFNDtSqDuJPj6gQyNEA4I1HpKeR5ppIQpC7yNHvs7FVhXRKuSxB
SSqaRO/gK6aC9Kcx7NASqGOxfH5Fo8thFCZIE0lE1w71u7m7lYyj2OdFbwZxd2S3
RZLLTL2FLSv+mbgRvBwgr+w17kwtuAnyi16KLbna7P/fuQY4K3FxnbjAFEt65eVM
NMDMc+Qw7jDHTdoOJzYMEDEDSIEv0uvb7vpS7t4GQtjwxMUFZQc/P3jVlKGOIl9H
o9ICv8slBiPMEy7VooCkNR1O2sG9OQb0UDQNfXp6O4EfkF721b+WKey7V7XEz1Kk
M+LhMtJpH4gROO5w96u5F6m69PoKeu+eDGR3fTA95zdz7wTnWbfuLMj0sc5qWEjs
0K+TdNKslBZHrloD+KQOtDXaaVcQ8/pnI0LBxp8X9cpwxO9GFTGM5gxjyvVnwL3S
KmeSkMMTJNqUX197kMY6ag89DndoUwGbHSzhjNAmTuUfzFPu/4Fa7yf8N0TcF60F
IL7cJVl9bu6pXFzztoBwie3D875YGnB1Sl+gqG1+qMFBll11M14mM67KwFJ09pCC
5N5oXdC9bFdF4ajt2wsYMju0AnaX9RjQ6nCMiM9tT8RmhLmf+lwoZ/TnLtk45akX
o7jqlahXCZzFPfMvAAYEqJ1ZjqzYTgfK56nnXz65/NDvSUZDNw2zcwgfxFb6JE1N
3hrpTULcR5cWOrkCOq1slcb+zmnFM/OB6ZsLUuaQpy/fvtEwMy0b8oGQWA9gH+nl
1wJ8cA4T4PB6g64QtJKRD8t+yYFdT6fXQf2PX+lJMdTYPFMSUHKoQ25tT6X2agaD
zsbXPr6ZhphaGFw/e6BkDG555XTHb1mAVVxV9InJNITJJJJftilGQmwvRw+NnVS1
xBEuIXW0co1W24lmxI5L3NegFpMhLRIfB7tpBeEjkXKaVLiTq96Z4BSdGYTG7e0H
GmPdyYjFPZFj21JrRCywR2hNMNcHxTyuIBg8K/pzkW7W7cKtgcTdiOyzhIDwf7VI
3F2SmdhNERVbVMj5FVOVSjqpcPYuupqccfJLdDH4DcntuizQKlHWb3znrGMoZqJQ
WOBbSsU9A5LBCK51jnY6nIocFm80GA/Q0XyStZ3Rw0KO8dABWplvwyDCQm10d2/i
Vv82XsmEiu61xpNqH8M4o0FgTT3LdSjGZ0ZEN3IP1Gady2pLKTdVvFQfhS7nSvs+
LzP1lU7fHzCE4mrQfwkK8nJGGQ+aTgfGlP+dR/fa8rkixAayZ2evqPukv94lF1AV
S0gvbzN48qDKbxzTthrGXDB0J3D3zHGc4C/gDxsGKqYFNxSVAT4bR8yk0xK4p8A5
4+UQrRDi12cXyKPPfOhxkCiKVVzLMaoIPdEt1TulzVw59Zkp7JAIaLGpizYHHf6N
R87RC9pQkym//gNU3bbmisp120acKTANpD49xC5zyVjBY2Pw1YPwPZEeXdo+72Uk
5ipz9Vr+H3hXSA1dGZXUZsPJ/7U93hOQkV3WqsG+PHNT6gUSKdOgOU6qQ1OHLP1T
lFOG6mfmkSOiL3/jeJkOsKi1mQqDWzw8vt0pWQZFOcgCP2Xohg3lB6oZWCPkYQuJ
0FhzkFYPxzHw1lNYn7M70/ytNkFVhZTBLznHZtlM68mCA9Bjt9/jEXK0m3NeOOEv
KUsLKhjF9K1tSu1i+VBwT2vy0TWWcpUhGmWWl0biYzX/56atrtM1jX0kH9XOmDx6
gfAC0D/ddeby93TiPu/zYgCAsCgZDH0/0PG3iv8EVeyuNq+Wr/s48iOYvFUIfl99
2yHacF+gXomNnJKNHHMTkvICgHgIzVHuwjHUlHhaF0se2kgyKfg0L+BVihBYdQNE
a/AfUPueggWKn8wcAdqadc/JmUN6jvrR/l7Q7HoMNIRA9U9oEOc+mhsK0bIS+xnE
nJ/l0tU0cnhTnvkoMMTMOx/18IrLSAMnoz2o13kP+v5rsK80xFi0cnMNzKaE3EnZ
Zw7bQqYAPU76+58hbag6711XPuQdgx5BUD50dMWcgEf04jFPMTQI1mk/tpXnfx4J
1USR0TleG3r6WNR/2ecskdeTPRPtiW3DvbXF+v1o5ng6SnnYyjbXaCczwAzUzA76
tTA8yr6pzY1IoYa8D+Z1xll+uOvz82ic8/EKK/4aXDtZNC0wN+vI/hiZnfwm9ZEr
9IlTEEWw9nzbBl+rSYMtR5qxPUplTYcHiGCVHvhjd5M+YPs2qKT63nW/7FbOTsOm
lcDshQoLRc19hbm5PNP6/f0g6EemIyMCxcJ/CM6LHP32xkWc2DQrCELWNnPSRHkH
+InkWV2Ou1aieYnBszKLVp8H68o5cjgOwNTix8nPwQ5I6bLEyG8wgodZeIlPs2W/
ajjs8c8yuwkGHaCoMz17dvPNf0d28L3uNi6lIIdlE63D9s0byHDvvyj32mQdbGxR
be1VSafiwMthLkjIbj2UjGpSCT+jvvZUNB1nymkwEtMNxbIgJvqwaMg2D4r+sQp6
zd9W/RjhiiPsexiO053uUhPtXC37WfI53vLY0GduQY4Q9/mLFMGPcB3UOBh7fxI4
PZXnYYt+LHoDmcgq0FXZZ9uoshuktEWwRNO4sIiQy00t9AVXipEaHXoj0H540cN2
1XrGI/dW6xYaLfvO7tt0tB1v5e7ryULfol35ePBxJYIo444bYomXlQp5wfDS/RTJ
WndymoSfxwGrLNh2Dns35tU7DpeusYi21sMOJXzduXyuiGAV8VK3n5PVoZFohGbu
LfCaMN9dlSFCJLMEkAcXv50IDsOJQr6cz3gcV783sss20BFjVO5Y/KlT1wEGyjfy
n7eUuplR+vgUIVXW6P7wWJTOcgXFQXRb0A7O9F+hp9f9nAZMJvWFNrTkJEvGbGNB
WNZmeNd0RZixnB6+cM/L+t+/KgY1HkU7RtPUgiRCXB7M+sh69+ECE+k/jwcOrKCq
3gUDoM70yZTdYHJcWkLL26BKKLF3mZ+56w/y0RZr9xo6v1ovnNU36eS+r3G48pTC
btI7WbUEtYpg6gSx0tYjvdvS95N39/7LQ7ecFEfeLvw2jayl+xBJq/6RnamgFcs+
s/3tbwmNhE8TUBGChr9GmIqFUUmDI1M8oZ+EzSMKrQ+DaMFzas8MIohBDvmhKUDZ
x3taV2xnJkj96Ku3BebB0yaN8L8tHWKp8qhUFM37Vh2IUQ6FPOj7BR/5Wn2ug6eW
vbdptc9lddhSs1hxB4NDH5AtQMnCdRlzIPd+BOutOcIer5YWV4aJg9EdHRNWbMA7
9ibBCbL5ArYEMI6Vus8LbnBUTF5z2D+DTnLS801C92lCq3HcqyFevKnwKvBxY1nv
J1iYJkNGfEDFtJk/KidqXeuks53CniJNLZqyNOyLLkDZPRiALsU2sVO3SEZOe1kc
y75/rSIvL6yiSAkRyvaQIXtt8CTk1D4aBJJbMGdizwtiF3hfah58V/zq+TxrSbAY
px/PhYzIyK1lpHgPbjEWVLFEMIUCNFYU0jn6H/E5B6k+PkUtl5XEOJ0lcdnLWt92
j0gkKS9yQ5F9H7feiAVR0fgHVS0dEdOlGJf32O43P8eYxXuZbRtNx5wPYBsEOsNj
tXKCgH/kZt6fMMMjii8T+t2sSruabRSXG4zFhuw9tPBiuHc/0GY+6r4WUmbTbW1b
tuys7Ywi2kMmPh0TCIAYzMLvoD2ESNIfBi0hg3O/dnHC6YEntyaiWjkrEYJrcQYR
0GVAa9d1gkTnTQOmGZJ/gC+CARG5iZu1WJgHF6NHG2XI+P5zhdnFZO/R2Of7dgXI
gjQe66miGm8vBOD5s+6pM3Fqz+pAJFABUiMMWzTi+rdPQY6TDmuHl3VvrSZ2lu74
lR7Q2CcSaNUFfmrbtmwbAaq2xmbCM7R2ekG4QGD2jRlxW2wXEdL1l8R91EBnoyC5
Dg4SLjQoqpG6mQFSnPQcH/MUYoF0FWcZpOqZwdYcufExC3jRq4xVg0ZSuxSxZrki
T9doaBTRKwKsjvlCWmudPj83IDI7z/HSk5rdu1s7vB7KIoLVYOoztk7AR0Y0vMvL
L+A4vzZMWdKQuiyzSpf2LjjxaBFmY1wtph+U/TC64eWjlktllRAJcpKrgHHbaDw3
dzwGFO66ZC2ds4feX1tW8W8ej+JvPV1EwCl9rEFG+oTsrcEzDj5soCArZOpzcRF1
fyPiCehkFWmkPB9fF3bRTwdWIUy8OJn0p6sJ2fpeNi5Ixf+cYE0kyYJWXEpCq2f7
uCIy/MwAe5TARSOns2lU5HBYhx3nrE+PiBk1PCqHvUg91Yp3xYhCkxSvNpG7evXn
pvHJiCD+FAtZP5Do+G5pv+JIB3usZMHuQ4QyOeFKn7aX3qWMpS25ZthfwCc2b3pT
sxeupKhxx3Z/Oy1ITrXZGVDZWp82xEezq7yi3nW6+Qiwh33MFqPgFMJFXvdFzCIq
zORmX2K4JpjG4Zxj8mSTNTawIQFwp+1fp0dtvE004Bru1Txzjo1Yug+TAZYm+kmn
DR1NgvEdalI/V0p4F0Ir55FqUJ37RfuT7HuA0ZZgLla6Y1iPU5/SSW4Lom3NvkXe
8avLTMXCjQWIAArAKBSgJQdv3tzG0Slqly3vO60kYWjQ5aroSjc7Yqc1A8rFy7DB
+ObhTeEvxSI+zcgXn0CIN6NtfwdQBI2ciwhQ/ttYgolFwidj04w75XSMyrLgM3sr
7IcuMkM1whge20dI/Lmi5evIbhc3FRt2P88mCWo4qakMKkDRfz++PWD70LbOkK+e
nUBrk0BOEvv2odDnlVyI++28fHRG3WzXGM1lKcdRxKS0OWejiXbZtvfN6X4+3ANz
hwA+N8AfxpxuuX/rE7s+OUfZjwKVidB5p8AFZFqgylK35fiP9clwrWJ4XQ97WzuO
ZBsXw3XKuF0KRrN/QQzLGm1iA0aHLNt+J1sDzpFNy+7zusxPWSwpMFTz/q8fNU46
FR5G0bTYE0oZk+5mqef8R/30I+1WrSHKlOlaA8wng7E+HLYbnHkunUtqmW9HXaxT
KLiYCe56Ip0VU2xM3bmMThq7rbi/JZu5h36k44SwpcVl6dqPO3+PxT4lFZdRSHRB
tCTMhDyKrAk4A5oN1njMDvg1mJQJLcduyUaVbS6h8CAj5OwU5NFWmtLZf2VZsdKw
KFFMUEZ8983Xz9eMvwXGIC+hgnulLWH+/ysk7DxO7B1xMR7B7HE7k5yo46IKwfRG
aXI05gVeeGyB94B6OvLtweDbUluU50vsBtcdRxB9jCYe7AszCHJN7GfEEgt53WOi
6G5/8ZOwq51hbOmteRWrCd0HKwLVn/MZPw13CaZD19/9b75yGhm4IPlblp6J/jHi
/4iByTxEZAihpf6+QRGvrXciGJ05E74HLLi/LWlsQLMXSaNgf2rxOO2VXtu/1pqc
nvk3Riv8N9KMpj56WhvWOm5jAMfHGLhrHRRPgE15e2+oXPbPelkBJewwGl0u0BEi
TTfsv0R6IjYp0HC5rUxw7hoTtA0Tj8kFItSniXSaVJjmCXfNTwFpsA2OK/CRo9U9
fvPUZBaZar20xUADAXtZoO1K3GTHe2MkJi+qSBAQM60v4cKw6zD1rHnwuBSiMKEo
F3hnh6RzG9QvaY6i8/5dqa7lC+8oi3XQjWHhdB1SP+jGazcvnE6beauxJjQ/Lxzx
FsjHexrnSOagBXDK8bzWbtrBWyQBUjyEd1WynXgmvLANKs12cka0ERp+oD8aBc7z
m0ZkLTRXAxdv+7NwyU/2zN+5Xnebir5iy117h4ItSxqwI4mzHrOGJQx3XND00YBp
JvjS4FKbVp5rBuf7hjotoR9sgNJHmQriXvExHg/JJ0Ricp2sAvu2az7u5zWtbYwx
uCKDg0m+gvUke4jcnkmNaGZ5NoMh/6LPTTBSu5ffqs1CCRAUXGH9BOUQOd9Oyvyu
fTxxP1noPLD316I7bLLE51EgV+tP8TcJljJOvCoRHNHjqaGb9EeElnSzojkZsllM
J0lRi10IQnqbL3ZRt6l98a2atzWdvsb2IXNgYH+7bUS6NVERkrLjeroxYZLtJqCz
JnKe+wUbMQaczso/w5V+h1C8cvPzzQE6kL9sF9eTYYfa0HHwwHEnwO6MuYDH41y0
/v8HRdvem5PG2dZzHfN+NIp/UPNTaKnDKlTQNGS6evaU+gCsyattQXbrB+vu+oF/
0IAKYJsX3T/Aj5Jbmi6hLT/Y4Uy/lXkBwGanV8XP2yDWD7IKuvyxek6tzpFl1Rla
g30hYpLNMbrxhN8Yxjlxof+7b8Oq35+lxL94FEymNNDo7zQeN0qV7db+S/C3jWZ1
6YxMwN29QSRk/tlgCCaqxfFUTHBCjul+Tij0BZOpfxYSIwweML3sG5zqbkKutDLe
pwbYNjhm+6f+PemWzGwi2tcaMhJh6Mp2XzEzLkYF5rh+k7MECafzphGGZpSEpfRq
UlqnKuuNYJ2B/P4/XtMydnx+2ESNGisTtITYjsg/mjNC4TOc5euKHkKVcKreoxSU
rgmnLDB8O3L5tviYdlUlDFy0R5L60enmZkCkZwYvBPcaJpWfvUn/wXdK6wREh8il
yMNqJyxZienRrRj2+ixKzaGzmEYkAyBu0LGNqGu+hHuaU42eai5GYuNxrhMmyCbO
iijaU5Ku25nsmzXgePlCZaIcc4VwWQEaOqBCLtg/mMhjKpsC7oz8B5WQXz4/e4wf
DSiiZnSC4eWcXID458kNkQ5w7Ik20+v0bIahKIhSx7uK5fItz6txB+4g9dNYkJi9
L3liKRKbX7j+dTbJkDPXRzeKs5XTSJyPbW21q7o6tKAvwIZ7CBMyh3Ifoj8KcJk2
06W2XvZRjytiHodT3P/ovuFNflwark+oGaqq4ON4F/BGsyZmbm8k5a1Y6eVwBjUY
I2IvVqq6NBwWp556XKAXdTeZbBQGP3eOF7if/BxrelHNgW+dSzFjtsuNBTCVGuL9
GaKXlMLzcEYSLzi2fyxW5ySfry/wUAm3lqPPYXsgRiKy13FMCcj93lpQhdiBw5lp
6zor2QC4lMFqQVRpg/Pmw8JayWdD9Z+c/RJfORQpajrPjEPXCCFKqyAKomIi7XiI
wRS/MLZ5ezbeCtIGwZOAToEYoz5Gh6h5iiOYRqGhvJF5qy2528pZ7ZOdRj4PyIu5
UVEfF3FZ2laEZ1H3rRmyKbgwF9A6RK4exkhNLBBj8h+9pmvBC71EkDu/UDBifTUt
Nto8u5ZVAsMlpIjiVZY5bfyYqihlm0CVjj2ex4VpEQiV52m4jjMY30Ulr2/YREoK
BcBI7rXMWOlTSRSjXkkvl4r44NFBg5m8LTs1GOkmRYOa2d382ksdONpVLHiylwhC
sWtFhmX0i2unpVTy2PctUeTVF2Zp+EtphTFFNQClmH/u+eHoBkvxQFk9zEsH/oop
Spv+Bjd9agYomYjNWghEGvjcdLmcICYtlqRQZugfSJdX1FNX6nuN2QDxjgCbNFkp
Wdip4n8X74Xh/52mzkVkWQleX9LKIBYCq9Q8mqi2fhGIaeb/CnltPpGHIGyFEmTg
roc/rJs8noDWPwznuBKPWiAFUQHzx9rMqQtRzEb+udo/nhn482MbQeREbHi1YPvw
uEntkdhTbp2Qvwdqq6Yz6xhuGL8ljyWlMJNaXtm/AmmtnmJFw7H3Z2i0d5kSGrhb
RMRSMDoHwz/ug9BLQE+GO40RM8PyTSmnuyNKsvZ62MjLfNHnWVU3UM8MWLzGXLO6
J1g+k1Kbf7Bm3aXMIGLtHVz5iUpK1vPAX9IvjQ9wsvv25nW83Q6c+CrDPPduuUcn
2ciyWphkVa8Q+5KZ4YgnEr1Oae7i8HvGGHsp7+OFg9sRXRqnZQq5XN7aqVk1smLi
afvblIM8LGUhik50vv0o6z2wzx2r5LnEjWp+rPGjVGfAS+8RAqIWiZyQidy1rt2N
XjvA9KpynFS1T3q73VJr2GWRHRMESHtJuKeiQNO72WQJc1fJ6FUGKKIApgyBnb8o
GCsFa4nHKTGJ9JpgSNZNWNpCE2NOSClZqzrQhSoy88oYXRW1EVPlRBJ3j0QYUXMm
+iy6kJxuwX5FA79i1V9JGw2I9ofkJfer8nMyDlwijJXDPp4NJpRfCVHH6M6i57n+
PoPM0Dd0x13Gs9Kw3n9xSjCseAYtYsd8K61bpOJWP1TqmUvf1jm0BCkjYeqgF09+
jCe+fcO5kgavhIE6D/4wMVrgEB422DlIIOW0jR0niYlHAKseqgyX2Z2DZn2aE6G0
oT/f4lPSjyhPE0zb4qdsPv2Z7dlsPPbvWa+wabeX2v7IsvsuVlZt6G3fa6txpoPy
Yn33G/+ZwhIU6/DS5r3JUDP0w1eShli446I6fzbtOMM+qpo/z8tEr2XOUdZGhJFf
K1rYLQ1UWdWpwSJp3hspq8+ab5pY4IeHYZb3Tls5Y+lR62DJsG/r1GZYG4Ya//PV
/dCNEPh34ZNIMWV5/VUS0mR31uV/Y67ujCc9oWJCnj76LRU/yYe49cI5kLaGFZH6
mCUWDKQW3DqGtXuApn/iblPYQX4YZb8yKdG3omhhizVoF7opTkXn77CKrc9gHIc9
47XqfLuAIYOJ1nxueftHPGT+hjZ2rxBIv0Q7NT82oRryc5z+LUCxliKEEVC9LUto
JBiRDR9hQnsZw/Uy9POh8aoZe79ddryc+YUkUCQoJX5YnGgSm6C3HqwfWZCI2HIp
DLpJYU1d1U/L/rgo4TA3KWVjVGYib21cQqa2/Fw7TKqZFDOpXuMOxoMlFxhbiFlC
DAYmsl1fCKsmonyZOLMkxwm/cs6DSsdR5hI5X4J1676u8cNB8tzOZOhYwDNLrvDE
vkmEPPnHdQULfN/pJCpNiI4VPF2VNo0wkS/nU/XySA5ar/+n0QmIkansPD5EDM/0
A3wwciuBMPOGq5Eh+UP2/ETfzXorYFH1hj7RYBwIgs6Ky8F1ip4tM/F4kvgYVxLI
mnLOJqr9c48O7BLsQu49xcL04rPd88/yNSG6BPVAyAlO/sJ0NP5cuPa73yGG6im8
5e22jIF7XWRpY/rLhaYx6+PLwnDVkS4BirMjD8VpLBB8YFFjIcEhxFhidwuzbUPC
Dcp3k9J/aF64pJmoCTxSYYbFgbCxICeFtiNG0SjSRkHhgpSwOCi7fKFlgZQd0yZO
lmydtYyBP3hvEzZcBwbgd7aKe7kmFb+hDphLRkgLAKNcRAxGLqKSCqFR2lQ8deFf
i/q1xs8DjKLYdozzb12+WI5CVdtTDxw9/q0DfyWrx7hdyvj7o5TCO1gtp1VBO/tr
P5uoRBTeMhFT6TGRbd9MmSbOT1Z8yT4Ms/WjPwidvyaPLcgbwLpAZyeDjF3VCqGb
IVL3NvLmTQjATKfcGXsRnt2f9uOZXPpQOC0usqvAuzZ5DxQ2ZmXV7Xn70thc9oV6
WfV1ZRKVn67xqVJAQz7gw9f3oiHt9kP2tp88AD0x36U+pVCpINs6V1dNfUvEsh0+
MzPBNCdgg0jEGnaURtt8st8pTxYKTdQ68vOhc80hQu/AATma7rBQXKedDE2Kybjc
z1jEtk5FYsxWyRe1aKXfD7JIbqPlQp2EXj2gtMDEKd5YdpSsLUf7p7+DYEg1rzxi
0aqzppvC62BEc5lcCXm/onI7aqc4W2OpS9hWIiXSjIdWejhoFGP63xxP2MXlu9kr
sEoTzLayIExwpTHumvzT8VdhaI3osyWiA2v9IwjJCKERXBfUWApDElLRwcHgHkeI
8P9Uhmggu3uvCU5z2CGxKgtfiX2Fn8fBPb+eqDxvznjTNqI3FLzcMI3iOldKgFzc
LCXfXs2wBxiZO1effFq3WGzOgmy6uF8v9W0Op40Mxg+Ss2IluqUwnzgPf4kGmPFr
N9zQ2gy/zN5IJf1kXhdXOsPX7gPl4zkrNJsiqWkPn6/70d/DNd9m6hqhN6qEqfn3
ucJtK/evtNTTrqpu9Nz71QjqWvS2eBTYrhGbMREt4ZTDVPUKBQ2Ry53ylVTJzM1a
Vtq86Qbd8189tzL167Rseg2uiPc/B4j0yN60g1kUOjUAvRU3CFPUlf1jr/aajZps
Mw0guOiXMrc2rJZSFbQJ0IK0TxwOpzULwxQquza2LHdaLPxEfMMjYkN0vBdVoiLa
KKg8Old3lIfzuXxf2TVAOqFKL0QJ34cxH8hJsBk6Y2fRrWPVYbPUR83UF3d3rfB2
6KxVUUfw9i2TuwjyqDh+98H1MWyTOI0G5oEN8owJv/lXp17Lgycbf3RmuZN7PTsD
Bmm4e5fInrwWbdQD9eaB0bIHIGODfAyMbdk5VwkGOon4bwKZeGvU5faiTO6QSHe5
yP5c+AstExZEgEOwj1WuWpHL9YLgvNhBy2P3kcSc5MnaaYHDikM+/freEV5DmwfF
WAKoBO6TBkMP7fvTakODVZAi87LzjrlrjP/IwLRT8SFhIbjLmg0NB8b5eoimX9Hj
S13WrtJfcMxWvDo6r2G3XmpEPDZvYtTsLS5/oXIPv5bMM0eTIcDY49T8fDQk0xRU
rTVK+7is7wEmm12xZ/LXVmAZo8o2sMD3er3RiJ2N0bqbF+r208ePHBEoe7zTijii
SXn93dllEEfa8i3dTs8efso8AfEzg0i0PMuFI9P2FUFkzAn0ArU1GBCH28JUVHTA
PI+ncgr9EtEkHYMLxjonz3wmouKF/cgGVTlCDeYZWPd302LNkoL1RH0Kqz/pAXzG
K8adEGrdgy1wySRRAbEMX5cnbS/NAsUzut/spFj7I2VpJiQ0ut0p49WmiNKz8k2e
xqDdodI+T+abXhqWbv9/V3DNv1v6QAK4ZsLuDlByaXH8U2kXNLm6t+X2KvElaSZ4
Cj/CxNer5weGu7WzmdIZMxxLHRtU/iNYsO36ntTEfw0tdo5pnj+3Y88j5IvrUoUa
cJ0SCeF+4HP4eW1QDa04QBzsmtZF1KmEQrGCoEoBsFEw1vWUKgIMhLZSxWHVvBwM
mPJo6XSmtN2m7Fu1OV1pW/kuzrkZ1milLMJCRJYuMIANaKumBTJ+GNH+83eFve1A
IP5aFHF/FPOMo8iNGyMRD4vjzBF21yQrP/dKC+7D8KNqUgRqpuhBLpvDs3DnFBTr
TD2xKRwUMmFRRuOwcD2P4CbzIRXacDWphG9IX9yiU1H1Hm2xMC86n8LdzfNvCGwE
ajql3x958i+r4ueuNeq3Rm5Vz/U9q3YE7yQ/wkvvooUHwKGUljgAQ6P1SBO9j8Nt
3DUEJdrX8gl5Bj4cQN5VaLj4SfZP37KtNu9KW2wxzEelBixZ24ZsD4Yp06Tl+JSO
nd4ryomZGpfi4XaF1kOZLkNMRdrSV1rpi90fQuVljI/YPv9CZpG85QfEcbhJE+2X
V/0D0s9TgnURt5vUbMgZjHc44QveZAiIZKU2cVWceAFOtGg173baTcxhp6x+8Vp7
IaeKVrCHT8ezcDT4n15E2lix13EcVDfLh23EkVpbEx/Y5U5AlcX/rZDkisTSCFJK
fOttrMgj5rNJqVFjf60ecFt4PN+Hp/pT48I+qxXGjBJukXlPGqWKzhLgay9gQDSX
PFUGlRkmCaWW8zqVrVTtzMDzcW982MNA7fS1Whd/JtcxdQYjPyqniQcxAE9AjoAe
c+S8vW4OHREuZKk4+a9ewW7LCC9M38PHUHM+Biftr8T6TDrvUibiGrxegDjs6BIW
UOvXg4qN82y4WCVSd/LA/aebLi8TOmrqnhBXdUL++oDsdCTT/2A3foOiNV7STTR6
ZqYJnqMUUZINagAw9+6zQcqDbWD78eMqT/PegB3Qy+1nrSet78xn+4twDkZihlIT
2hmd+M9cwKPh2LbOycROYUAnaEp1hyWAH604aP6i6MU0rJAJMS80vtQK/PJsYjZP
Y3YR4pjX3SQAQHHth19njiw3S1Ec5RU9bvyTb08WTVsFbMxcAz2C1YeMG6sKLW34
XzUXYO5ZfG80I8S/2uzYclmDALLYHUlSi5SbgRV4a9n5wFQHz9s27hiZopVaOsxO
nFmy7YkM4MiF5hN1jNj6mR6E3+4nqvmUGeLpP+iO8U1QaLht73uijtlkqboatWJq
M+faeEL+5CZ6nz1mdfVdwtzSZKT5GxsuWzsvj0x177OY3FV3257nmVwmYyj+4u71
D08tHR6eyAgFIBzDja+V9AOMRHM6MAx87U+qSr/28qdVxD9PEgH+F0wbXZBhhCiw
6+h4YcivE6CK/tJxW+FmErSeA47YLCroVh+Bo5qz2Pf6XROrp4EDGRYMyJzjYAHp
QkN59gM9vZeJwFkobWMUm6aKjEhrR+0fpSArqrznSNAKzosceQHSqhwVWtVnqcP8
ATiHm3BQdz+O8DrHLaGvFijuz39iZiMNhSHFtVruDWfJ/d3kFwgniR7hfkG+7hB6
ddFq+InePCgdY019rDLC3Lz/UenyGDltrzdPtltkU7KTtkZGWdRn4Py5SZ+UCMFd
GnYjtWOpsCpeYZtSY/1jA/qncNiBBkfXL3FeP4zbIV/Jygy4Ht0ujr6dSh6IshCc
EdUpstHPHMdPgjGn6GYPESGL150qGXB3IDdt2kGXljyMnyLX/Ns3MJrnDUzhsYDP
ttZ+dmMRDNHnd6mkFPnMsHPnK9JnekqvdeJzvWzNa0uTx7a9TruA/wah+xGvC0Kp
w/vFBLe6GmXMImg3o4KTyRL+EH0rgpj8yWUVFIk/go0gNqSL/yoTWQAa+K6oX8EQ
wCYmeyPPm+jY4Sc6+ID/pg4lun5FxpB9VEImldkJXS4Sdj7Ni9NIrOv5vNDxoUl5
Q69AMm/dD7yeMTJ8zhrQr/H+5rUiGhapbSAC/dHMVY+8ASnOuY+8ypjIKH78Nkx7
qmVGaaM0wiqffjC32TA2PMH0eAiHEuuUclHJyhkErOtLbsqne8U/mn7QhJTuiCDg
jS1DNdP1TZscR+5aeYd4jOPx3TE1V3AQke2YzsXtFjw4eBcGykrsqiEWIiyRNQyY
KgqS8mq/L/H3x+alqtKSHEOnuVJOV5hb33R0+HrZKilQCGM83KX8lMfltfxx4+Wu
kveMOXtS1081V+jFoa9h5NJYq1Z1RXyMkkq5BTOi8rBlB7zMNClHeZlTF8h2IF1y
0gz3gkHESSmlhfJjOM9eA6gPexFJUJtJUaBM26zp/LlMTM7L/xifrAn4GjAlkEq1
8PIFBCiPC7EGFhWbdnluywnV6FCe4kVDTykkjbYs/XRzxZaPAmp7rM8JTXQkiWOk
gjNd6fY5DhOWHblftQTZLLTj6F9vp7rfzvdy/7KKjfwi70K2aPgef7riYP08nlkU
WKmlcJlbM0U/uQcumK96j1R/qtBUx1onTmyYQN5sLLgyfOojaMvqJAVBfl05qTqA
p8DsXWUoM3Mi9SxqCggt9pSHdqTczv76mG2LgGHJfUASN622TAUzX9uXIWpegBlA
nmclz/r2FO22jsBXyF0o4bw+SpidpFQu/MT6hbd7d1RSAX+JtFysFfQ/tuuLgLvh
R7hofHqIMyZv7o6V/KQ98cWXkK2AMnQ9e+6ZWalbC2Krq/F7t5z41A2bc0+xmTCh
KX7MEZS+5M64bJa3oFfqMmTqdUMAEVYcNIBAOJ6AgHEi2E+Tm/44A0IJ0sDTNpmB
TYwmb0uzciQipwvsAI9tR7hyaklb11sdCkzFYNy1DLdazGpolrOuYZDJiwEu/OT3
k0Ma2z25h/Hvhoy4F218mhcm+6CWXJc0UPSyExMkJ/9FDEFnmlPWOiW4xZoiDz1C
6Sd3CuSec3sf3/R5LsKpnK44kglTrlW/whey5mJWSX4TDD+p4ZrOF3ZOFo3kTFJz
NTChvwj5kO7q8ZF93W8oQVekGRgiULB9dk21H+MjrX9Z76LXWfc0q73qxw/P6EbP
gQgfyFqXiqocZALe+zjhPNF5O1QfzTXGunjrJPnCbM8Jt2ogw0QS2Jr8KGcxJPSz
KiCv7Ssi4MorQwJ3HR7uy4iMLjCBt9w9DWnxcIY7otCg3ah08g9x6iWOSFHvDo7s
kaFjnYDL4JZajzW/N3jEkUC6P5GejcWDnsl65NGJF1v7EzoH4Q4f29LmXGc57tGo
isMISfISr781qsB8x8iXLbtJ86PRtgplgrk9kzJOViuHNkxzoextEj/7m7nXqsrN
hhFq2DGE8rf642ZkIlvDYRU/J6Go+RCqYfHDViHZ/lBRya4IqZfn+D97IVmbWKE3
ilbekBK1OClkhQ1tUr4GwBmbUk46JhR+QH/AtfKf104c21VZKp+90Y84vr1yHbrw
EvSu4zFgeJP65PWm53REhp9wU2n1RdG+C2lWHosL0QXKkQWHO0EENmm6yprerlJF
jkEEo6717AajzDGeW588+PrrDsCX34umWJH1maMVTV1w+0dPJ/CFSj5jcTOZysE1
xVJpntqjPm88346AQcID/U+hDyjdGWWLSog/QKcAmJok3IgJu9i168i0/a+WW83B
Fp07FuU79MG8btlKkF9SM5LsQi5mXDbfaa5PNyf00/yg/fBTOG8acNgQVmzJEcKP
7sV9Ja2hTf2pYgXGawKDdWGkkbG6y3Xx122jNCwmVh6o5cLewsiC5VYZynbXmMBu
vGfP34A2Uc8h0LWJL++ZCMgN4p36l6o0xDUebdO07cixpAnX3AUPbPZeru9zF/Od
48m4+zYaAuMSI0Dx/u9g6CNxKFbCUOOgjNFDqaK4Ch5elgLmLmoW653UCAWV942T
31bCPPYMRrEyWM4MaPbmecmbNKvtLDLJKeHZ5wlrpUBDa22YQ9utsc9Qp+h2nrgM
Q1yY9WNksiryHZm/4NcZXkVH266KEgdYSUB67SR9T7BZN2qU+HppZ7UtRTU97OkR
kA/AwVsQFP1F+dLS5tQ6ndbJ4yoCt2cQjhXWCTZz8j5Cwdq8SE7CZvVxWa+rgxg6
rg/tHBYt9okb+g1nsnFXsDYsH9Kv0lz86QDirxDHeigNICmd/9vHPh7PzqllEhRq
EDiH3F4vl2qT59Gkqrj5XSoJa16MluUCV/txO5OaX+98vVqOyRHwmXkeB68pkY6K
7Jx6omKflOADZJ58t8ICH3ouvnHrkLmmPcc6vwvBc4Lt7OtcyJkXDwsT8IIR06ww
O4/F5vulimW49pxtKptiW/jRT17mKRkIvCRQABA141Lws+hem3Vb4KyX4xavPat2
aQoUWtEoRi4IrKri6l0cFNc393q+ebjJoEjJHa5nwANzeAEenJ83KGP193aKB7nU
CBaP+kNkpwh9umYm61cCnfCwR5oJV2L6pJGcQPKKSzlCIvytkN5ne5FjiCwRC06B
lKm2DCJACgHdInZFESwuKman0L+HVEK79mREqCDhnTjQ9j1Lc1zJa8nmsBJnLn5t
EF1excokmhGIGkziGUM4oiZ5NGNv36fG2oxuNqQmm/pex0KIXU0P6Ek92YEFxJOI
U2xqp/02fExlH5kE8XaCKBdVddMcVkB8XXjq6NIsanukdmy2cGXxwlxjd49d8GTZ
yah0cUynuZ8rqdshhD05cPGmJG3g5djGzk8c08S8NLriR/+EvYbel95zhFc/E64N
T0kUfHLiCN0bguZ8++kPOxMRH3+A4bmMRIl/rIo+GhW2zEyDrycNNc59tSDUKbYn
bcggcfZ6S98l6O9G5ZpnEHQ3oj79PzUGFE2Ja2LqkKvEyA4VergJH4C54At7f2X2
3X44euHA9s9JzDCPaLOVXei6Z89/J/2h+22f4ohohVG3zp+CfG6QThNVvJKIylFo
m9Jn8wnVBhEujubjilV1PFoedg8l148fPbuJU6OEbnGN8oijQ6+i4ncPuQ2uOPTG
5sg832/n5bSyQwJrXFbQBkOYFKftPVkMR9qCt4/aQTwapYxWrwZjFS8vdXa6+pGW
Gr0AbF/q5vW7wVFnJuGk0A1DSIEUrPjDNSQZECIDHxFPtkhC0UG7+JFuYXFCuVmv
KIKaEwxbb5rt0SbyvMoJR09dJra0egRhaydAD9ptywrCNv0ib8GGgJFiNZOx78SP
39Q8k+uHDskQAdbQwzI6/PFD4xf/2DzdUiLq6L9r71Ey6MLQkWVsiLPQbzWs3lB4
axBCqgoQ/OJIwBhFFrcVzb+pHTUHD2vUIpNiSY/WHvnSch+yKrwdg1eKGifTX2RS
TL4lsk6NNdi/HI7IO/+/KRfuv1ux9z46UKuqUMRL3jaX8QNmct044ZgXWtWEww5y
MfNp0AjY0dl7s/IGbugaCVdWOB5ephpbeSurzbC3QOLfhDEyKvUQEv3NzPhO/PsT
0oiw95gXfRX00OUiqHVmjTMjARhtnjDmjvc5PAjap05r88EtevY4qQQPOX2TEYvZ
qPzigjIh2VJc7XQXu0vBopNqsR2nt1pYzjLdbesqeZy8n+8Fu9jJ2DQNuNZA5PdA
buVg1pecVOnHYCFc/f5unYpszfStv6RHYxDNd8O6B88nH+rqNcApntlE1YavyEUs
Tw1WgYmsCjN1qwYIdzf/wSbgGIjVexDfN4DpiYC9VxpyvSScjP3avrMNEzhahXjZ
JQ4mMz5qceJKHxC3ELtJxp3Cd9F2vvzxxdDrt5fd1pMQvtMMDAFwoiN5rizPbd5+
AF+L1Vfdj57+1X69X5OoYRTIqGgZsca1ik6C8jhDq8C2BVzMNeBBnpJlf+nQp+zK
ExU2F55Co1noxcgFyiB1i8d4Q4N0oDsrBz2AUNpfRYe00j9NEadA7kKwewz8OGEK
apMuxSWLF5K1fo2vujtL3lDu+5B4lSMOl+biZspQ47+ZnjrvaJiNObxOxb0dhBxu
E6qzJZx+0MRFDrpL16SP9J9+Cw8n9TXtOWFiJA6K1bukQiNohZxMy5LroqJykJdo
Ht2e6vCZqLv6RNIZdnTpSyoxhAv2cCEqSt+EtIOKBjRujCPPInGPnBYBUd/h5bTU
psQL38e0NrBLSQpqiw3kera7UVqJ+5mXaIOKoyq0bPYnC2/FuBMPdi8LpxSvFlM7
3keUIXigLcEQZAjUBFpof61WM6ZfUz2Onz6V2pEsgidqovHShqaQHcS62nllJZTj
ZZaVLMVlnJnXvFRB//7m9QE3V0YNyb694y6NitjLstgXPlOJK5r70tAfpUOBCcB1
6RHt5JlVvNGIqd6umXjux2jC9iIck/7dCzGecLPWn57iBVZ+iSbAkAT5aSX8Alhk
ApFM22d2coFu6CGj7erOmDSK22F8+iOKyq2OlfCO/XTNIjPUM0+ZBlIFaT+f2Evn
V/8K4zbQQ7sUM3YpYHn4a0sHS/Pp/UTdGfzbBKFO/NHqXCrQb1jknRztyVBtSYzT
jJuFF9fuHnxW3m24w7jhPIoJUfsI27stNpLw5svzrKBmlKbsK01wGPIQYQasH5xG
hA1vYtoHJKTg+r7QQ0tp43p7XxYNupY0ym2JAV720MYVd6FT44X6/zINRro0Cde3
pnjHl8w5JNAL5NxVL1CAowGV3SIA+DO3jCVBKNVp+BGV91vu6rDrTuc9o72upEgi
/lMGGKCd2d2+U9UiJbI8cOwV5zl5WFbsdO9fS6F/dU+Vs9l9JPVwxhQ9jKyHcOaM
I50rRMZmUap/HgP/gJ+QkuX+n5k6Bw8MiKaOOAjFosI2G4YRyzhTp0RwU0L+LagG
B/xVjoZ2JLu+po9TBfYQFvcsC0MmR6ipXqjaPmrACq1FDspWzA0nmFM+/GgHftqt
QyOdC2PXwCNsBZzxdDA4q8Ohq4daRRpYTlruShzd/i+G3h5clSSKtbCwua9OGNBG
IczMxI6cjhL0jdKRuuc0XznJSV4ctU/PPM3QOvBOQddcz+JtqkZIH97uEKhH5EvP
F7ZsqQW7r8UGVkYaK+aGJdc6YXtT70kLocjvCU9bIpmKP+Nlf0dRPBsTHl+ChMu0
8uGn3T/mxrc6KqSK8QCYhviLD+wJ9vxvljOhIHDTfoAdFo6Lj+2fpgqI70V//rlD
KEjuYl2zmDfA7OnR6c23YdxW7VjyNHwnCk/7WaqrtkT93z1xT2exG2Cp2VgO5fIJ
f2VSF53gmLpq2p7RH+auG4lVeZv9ZRAs4ZPLrGlpfORIsDE5atnPYiM74+Ka/VAF
249ULJk9GIsRfESYckIUni8d9bZXCgJGhf/Zo3YeCq5hQnJAFt7r/hImhWdP2Uz6
JZ7ZogAU2ie3gMD+TWAmIYBwBgkmc3tphGUtCsJejNwmDLPBoW4lMsxnmt+vIjvG
KRvArjGMePJvUFoR/X7yGG6Eix17RDFyWyE07c3YyZjh2S5aqN/xuPKg+e+0Oers
+dM7D0P9A2Cbeb+ckFQBl50JiH86PamK1baDc+RXAUc6OM3OFi/DlJ/tUGO/kVlH
1SxDZyl8H6Av/VYtXnniIIkOlBzRp34wSqXcVkvD3xOa6nALJH8zFtNzT+QKRBZB
TuyIDqSs+T4gm3HU8Pd1vFstrvvBXDYh0W5r2iOXRbso7asWI3/kHpZ0Gc+aO/p2
wuSRNj0a2F9B52gycebhjASDRAm6q/L8vNdWbUxbbXwuxAC4UMmFjYcghzhehNS5
JYNyfX5HNirsLze0sMq5Tg6CqwyOoGMMnL2uqpwm9bfY4Wfr62p/krkepBCel6jD
eFuBMzXa5BdkUhWbl77TOH3Y5hlK11oOacQHDtsvXM9oi7AFgT0cEA5YmTUV81hE
WVgbh2/93DKtC79jWqcO04PZGGroaEK5BbnW/q0YwEDQycP1sSnC2ozq7hlhnn1r
yFbgJ7sSDAttu4amlUzHsU4j8XLxhMhKCCxj2TXPmYLIvjbBAesbEK/Ga+Vg3Ek5
xrZxuBOPgMUhYRfqVoCLJ71rJT4N0PlYNiVyfaFqLQZ1eYxmkTtfrgYoyuJ7+g0M
FmzLQQuhiC9+xfa4IJy/ZHEGVMKekTZTEDqjDxKQUR3F0pAj0GVcAyPKddL9rwsq
1KoxwPliTihII2q9cWJWH3iw2ebKltjPgVpvXBRz7qdHAnzCQC0IBdWJNqAqOfUe
AaCsAwEv5XY3+lL+xR7Hgd5t/JgbGV175oD/h9iuBfmFZjgd5Uc4mTa5vsC259yl
ukhc+0ekCKsrsUWPLgRN7DwBRZWEyy5Gis6l+hhUAKT+JEwDuOSPh3TdGtFMRZA4
WVNFSDdic0wHB05rc+Dtk1wtLCaWtFGn9daRPuyZMl+uZccSHtDgRhLQ9ASM3XFX
ycBMK/q6lepyE2iJpWbRf0Xal0jbhTQvQr/+epHd+hc2vzQQS3EBHad3K7HIOGB6
ZUb1BW22ab3KPGFdu0yDvPBAu6ZSeCOT3s7iiqnBGPfRwT1MVVTf4ttvxquLJack
J+YsfyLkx3xS+Mm76kPPbcNmo0fAdN6dsgoO4BtzG8so/rRuF64EUgt2/tnJ8xRi
eUVBBcrdYP5ElMa9Y79myhsrXTCu4lhVabhZL17vA/J8I7dLookdoNeU+H33R46I
bnmIL4bdJcPKAF2PpSahvp9wx6JLPtEHdkUkEtHQekg0yw4wpwnSCRNfyBpCLTQr
0WLV+4jUNamNf6AHwY8l3rZXbJQmR7XjiE5kEOLxtUe8OiGNloLeFPZg7suUKiSZ
UNnpYcRrcp+wC1BxeDwCQq7wuIZk8F6DbEtH+8u6kHKOkpSYOzHEgZYu6PX5kV1J
p53emoD5Ar5KW3Vb208OkPgvzVH7ojAxBbCxHYl2tt3201sb4aLnxThXPK3mbCH4
btmpWCtqDd/vyRt0XyaG/XeRT9xtePxcmKWOH8gNOB7uDFPfJQwdwPHQdkbtGHjX
oJCOIgiJ7ltf8ElLc/NDG6AxQiU/IUSqVOsWCauKlbr5Ez12oOdSFUuWLMNw4rHc
HJEetjl1g0xt5iURJu5Wi+uEv1kQT5dsvHjblGR3KhlnR5vWGtgwdCBEOwh6tnYg
5WOCYN+vjy8aqwp7NEo0nAaf75/Q8DBWKXo9BIFyTT+usADBtmTr1SdYSdvZ5SWq
18BCbn7se9UASPJtGZAni0R2QLhZb6G9O7M7j3pTAkmqv+cXMrmniC2lEIP4q/1o
YRE7TbDcZQXLK8NkULNRsp3S/Xw9z8YKGkJvWHBZCzkeBfRWxO3jenKQTwyyagS3
AhS+uWicSxSMcQ/y4g8GJaRMBkJg4NCDDrGl6bTZ11yuORWsU+UXCmDxxxY7WHdH
jHWCYc9QaL3qVq2JJmHfPoB1LUSjVlSZ1Hc0NnvS6Cte4PBdcLNx6z46iWJAdeip
lUkMVAgp0KJVfgXYeVzthB6fet6++wyr07ZSpUz85nIgz4nFFuv8jnKePrE0Qx4E
s6QdkUk9USGJ3VVR1/qboTKElF9ZcUsLh2iL7f2eFHdQfBAJCLJsq9uAc/AKg36z
rYN8L2M9gLWwV8WzMKLajZlkbdPEvTRnonStberkBUTP+MPLrTnus8kzQxLaHE9o
PlY0lgKMlsx5i4AHzqqQ+h0uerqL1Xow2wXobC1arSu7AwQN3En6clv3XfAuhG5z
8eXzmlpQyYVhkVHC1SDXu5xQ0QLvQxXVRHg2pH6A7PiZVWoUYZIC+Kfi92YoKShG
6ZAGxsovkZm99mzwjAy3axyBjVMs/2kcOIwRjzQah5iD1XyExvhEar9H5qyaNBZ+
xEECNere1s3mxo2fkYkitpastm4tWvCe6cK1uE8bNUnUZwRWU1NFupgXlQ4Kq0yf
l1/eFuMkl/cezOeHQFvdZx4HAxPE9Y6bjEnljf5LdooYrME64Krs+GPHLdc4FxMz
5wRkbCzY9St231Pxy6V01M0BRImPT/EJPMtpsOJ63IJPZTi4sVQjanFWUES8G12Q
9JlPn1vQhv+g86dmwCq4NX1/mNN16Rue1+Y/IODTcvHS0jOvi2x741Qor5FfQyMf
+y3RTff3m7Ufi/8VdV3o5YefuOLh8z6NpgPR0uDAEQZ96DG157k8NlGvFwmZYYGg
uhCGpLEe53Owluyk4Bu24DTHhxrnOuiROhqrlcZDkh/VR01b5uun/o58Imcdvcnk
fWzcjDiBtr2YaCqdo81mqvveodtvI9caIkcBALgKOdvkh5j8OaJ0LPBoNJcpTKZw
0jfgihHg/ox6ET5kRtOflmtGzN5e1jfPIE1yQOXjG2ml1S4rmG6W+5hM0sIqQe4f
462yZTUHSLd3AvmCvvwB9GTQ4UFJiNkk1LOAAvgeAJxkuI2gPGddVwph5AHPoa5s
IuPQ1epqLEvsgxK84tGJfTzvtZN2MwPtGeBgRdrLysncAQkCsa89AJcVuSLjIwbf
AKMjjI+ctcICJF97mG+OSdl3dXg/j919w361AHOgW08GtyR/fUbnByDk/VAZmmn1
fV1muV39MmGJUQ2YPxSXU8uqETtr8j0ouS0nXUYjBK4TUXoJM7n8WfjUd8lK/zSZ
/+tnQEv4289vCJGKSkmdwdrn1OL3amKJqhsERQJDkz9qZb5wUWqxm5Iv3tB5Xks+
4G8k6/mweKH4gw/ce07D5pmhaj2e8hCa0D3Gxr9nT17cXH5g38ETZiXfct7yF2Qe
NEtumJU71MyffDe9ZVOGDdhJSgbDQcuu0hioz5t6lU5Cr6vUGS7awe/jEEVa/EFs
BkhTsRK8HKTtY8btTayfGzkbfsEedfFMCRTTQAHDRlf0qjSV/gXhSNKR5OBky02h
5iuNhtIuWzBh4iiEblzg1eWG/iSk+9QwcdEcL0ptvLjPR72wA5olDjoru5EuyucA
rk8ey4qOqvWPRHZ/p9juCMj16Qt4xh7DUPl7pVVeEnGfezVhKYmCQuD2Oj8n7nWD
Jl9bymVES03pHEbWKnjIJo8ipE5V+eYubWvRQxZj48EpaEGEfP+PzC5jdnq3rn0S
nXnjbrXYm4WNzxTppWa/GP24ZASNw3vgJHS7N64KHtlmON6HZvow8boYFCHOs0yM
9f5VVn1dOElutHQlBRpTk8weHXBhlWz7BNMdDoH0ueA6HIufbi57xsFxWz22uyeu
guJlITA+WClXEQ8ZrF4iTwIfPQ2h5TQZpRVkrEcA+UcDt1e7PidWeFdBF9qa2dZ8
agzG+9uwuG2EuaC/CmV6SLHNvumVpRYEJcbp8o9rdxd4aBHhbh9lY8XW2pGjNL+U
EjYn1OMDVdWNZP0fbYgET0OxnJYQea3mvC7NGIWIrXcVKpcEMOnnhaaA56CkH2Iz
WlNTWgdIuIMYzH3DpH+xfhYaJAFl0YLBfhif9UQRl3ddxgQnkEv4tKljxkYn8Sis
MPh/EpkwspryBz+TsPzrFmgRVeaDXgDn9sxRrG5KbmAU+fGf8CnY1sOT4dFgpdoD
JX38zgGODHBzX/Gi1XpYtdTdha3Yg9OYyejZmUZ2L1J0WB5FqgqWn/eixMuulOLb
kFJ0+8ufzyKpmg0vzFvfHLqL/UYH01YpCRONoqISMGGDtaIBCDtLD+CStbJ8favn
rAFtctK63u8x9ydLhTqZ12/JI8kr9QQ9+0KlzttWKUcVcNlf9PUPw3sHG2+ZO/5M
sPXsE8G7hyJPuvvFvZo7D15I4V2A5e5FSJQcrSgB2+tWO7R3XIQmYN3fFMWQ/jO1
CVDk2ZqJmJxnxsBq2vlXw2JP1Yt071gFyOX8ONVpLOTlB/81c2GLWyCKNi2BMD9T
gYZIsJztdKR6pJC+37QL/7J08ncAZCVffCLD4B/yoJ6uSxUdiLt5h33VkFgBXhas
K9jCW9aLFXKnKXE4vC26Yu6Xjo5fl1BaKqubzsZFKrHC4/VEfLu2WEziRs+Loh25
n74ZiVDblrVy8z2JEPTRx7Be3PgRpoBYCW56iw18LhHV2CuBluIcR9/L4EdjhvSO
wFMhdjWESB4zuL7Xoo9M4xG1K0PQsyR3Py4u9D/39TYMLj5K3gAWsfAFRGCx1Gf2
0reZ6aWOJlynwoZqzMcctirI5uL1xSpBqnDTNGLau//larwX2tcS9eWt6QxATCT9
ZqHflOliAXDKo5N/e23nwzuNzaS5BzZ7pNfkdKEWASdetGbfi5+u7gCb6mfhv4a7
ii6cguwNRZqdRFoOZgjHKmZqtIQhKk3xvhQB+gvh9epXtXRgGvMSg/9iOzhMg45h
JcagvSMkf7HKvbpjXl6DEsMJS/G4xeY0cug5aaYfroWyapiBsRkozY6+NpMt9wBY
ipGxKXP4SOTqdecHkjRziBwjpcdKDsr6x+5A/gQ1daNDQT6jkwpRBAOt7MdxY2Jp
xSbXtTvqV7e1Mcxw8IvHeiFwYgc28RFsCsaX3lAQ3hCWpLKA4OSowfkpK774CWfQ
lwrXpP8qKoTo8BnWlxbdjHDbOPxNO5DQduRup7QPYNGofaFN1Sv4LSe8/YsKzYuE
DpgkzpBSyTKOXTALuHAq0HlN4ib+K3O68ay9SkqyCtiIMMUIMvCDM8CtkA6qv9R7
RzLNHz0ZMLXbMjXV1S/041Ouqfbs/CqgMILC9DCty2lIHCciwjeFg3zDo/G47mIn
WwyEWHCPxQOy59UQjFKham93L2xYk/TOcDEFfKOwba7uzVcrHuULKOZKiFb8MzzN
UKcvmlkLSUHgyMpBD/u+VBe9ut62rda8/sH256kXG1jMhjb0wq3EL9/J6Ab7espx
KWahpV+ykXK6z8zVCmxIcgiH2nnTTwxpO/dlZwPypZSp6hc8f9gu1IEExr5lB9Ir
7e/rAuwVM9FvD6uJ/guV0zQWHvCVRaEYCZbOeEmWTL8f8Ps7+Z5pzRQnt8t1NFmJ
/hyGZYSQeDuCazPMB/8Q02LwqpxBFdEqlr4OqH1pxptgqp6a2oNDP++kdwmYjsK+
xCMoYyMD1QwX3Spf6XYVaSI6t84bbEip3iJQMx1m6y9/b5kZDoEJzScdbYys8Yzc
J+4M5a8lV4ibdDCM8APnNwhPGSJOpO1Q4qayR91NfLrzzFF9SVVsudWmQVGMXWRw
dTXiCsG2pNaH9De1HPz0wxcklGZVhaME0IgL15tti3lecdkVcKfsEdbOFMfTInvg
MzKOLHcyiUbC9/xtSCSNti/FD6SkPkICP/vmua2nfV1tmX8DUWTZqYvk7LrqJCjq
TK6HZJHp30A4fHJAnJolUTgbgPXYhybEa9g379x+BHjA+v8do/dvrSuw8nzpv8j9
KzfV8ZVeM+JJE1w300rjaMfRZC5ZFHM/6W2y9xR4iZxirKAJ4dW4bltdZ/O8YDdr
dlQ0yAJaMctqGOQEl/qff9kDYUwN9HD17a09mhkT2QgbLiHKpqi9T7f+W8yU9Th9
hdXTEcJu2uStEEiMowbEiQrd5v/Lx/w/fEXcOXP2ii9RknJLNDfn62RAAXid23fT
ElfjC2DwA9Dn4MpLKtNe77Xzl6TE/zUJEOgTNh6SIt7bBKlyyRcckPCjvgNytqoW
JL2Cj77Gp5yLs/Wi82oCux9BIdTz4DH40aWBNDbK/rmKTKep1FHJ4hbZGkIEhPd4
/kmmdXfmdzcnwQiilJg5EX1CgtiPRPG36+oY2C3zKTWYajKR53AoCCwzl3+iEU6I
nSk/HwFYKNNeC/TIk3gXI9Zkl5MAIMIeeJx9ico/Lnt7mS0VqXaN4oUDX5UJtNSF
iyXd5wt5bz4Ra7f9FQBM88nh8Iswrc4O3gwourfQPqj3kyry98Wvrb1QgmU7b5Xp
NogG1f3S8d8y8PrAwdZEGryvuRyzijHNUVQ+/Y3N3caoJ1jXK0dCrO93Xv14Q+qo
owXKxE6LQIa4QGYx5yA7T8aUyOGp3GPu2zOV0RlvxtBzys7wLZn+/vRRoL2uQNVX
xkUGuvnBtUBqhcS/Vf9q3g10LnSJv1KArrea7ZaClL+nWhElaKcEJjZgAcM4Fd+5
kKQ36FLmK7dq6chvugeYD+DNprFRPOqil9X9QYRWz+dARhGr2e6mCP5cyhm18eoc
C0pH6sGNCQoz5i1WrGqXuTzVhbXe1Mf1KZUz+qJyJHvHWnf5lmGy8+cnh5AUkHYN
lVZb8KrQ/UeI4SJIEdocQ7drdXCHHdGYrZfLWul5aGm4RDWztvA9OFb7pGytNLAX
/WS6/VgODypfWr+68NEvbM9k63XSqu9l/4To5TF3FU0XphwwqoSkfn8GbTYwA5An
Yyo70Oc0qWUX3xipdFm3yJJt4C5ryk17Bi7Piankbzya5dRYSAKzSBQJfFpq2hpe
CzDViZZuhwlwkR47IAOwnBt3TrszfI8KVqHQGwpTizOYYVj2vPIj7721PyEB1dNL
InNeDShDIJedEnHP1YXV/q8HgZfp9M1XiqfqsmPRkEj50iEn0O/qWlwp8MQmkAqn
AWSsqIJCNoB3pFiSEsNT1CaXIP+Ar13q/1S2AyOzO1Nkc3PM8YI4N7h+GTM7ipQR
FIrp3Qad24YrSFZoyuA8aMvi4TdVzEJvedcjEX/Piim9pPPXUIEl6a9AvJZzxwsi
y5dHRW8a3wNO4w81uzUxn2NEEXddxkK40cAla6Ef5v2dg4uxfCUzFZRq6Uoo67ja
O0y1qAMkUern2j5nx8uQeA7Ri/5HOWsKceElXCvKedvUGEMcyGnswKrVSatGQALb
Bzu0zCvOlG1ZFW4vtwxg6A1FrwQX4KwZ9dsuFUBPCLEhGG0Qa48nMLwCYc9EPfpf
cVkZjlrY/CdRlZKPcTURK9idFzqJi8qURY6f0H5CzBr8ngOJ7kHhiKKZwdCikpIN
4hWVpcg941qRRHh2PGItU4tuLHCPnxypNIZSPpWKaeAO+X0zlnmlYN+pxnCZ+En7
nM7h6e0McB4BDmNGHDP0fLZz4BNaMgfYCAt4g2rnoDLZSoqPC+Ij60UOv8UyJiyb
ET0p7Y+FY6kvAVw4uBFCJozfLR2ZIFTiXF4NjrPU/23qrtnaA4191hKsij2WkbeH
so8EHoOd5U+0vaENBW0iPIitxrmSqsrTr99XehGJYApBMazDqYFxPARlyTLAyP6i
jfORa/u1LRgF6AZFZuMJ2ElHZdWJrrw4niZ/YwXrKyllqHmC8aPWexYtgtEpIpyc
ReuIL451IRxFgaNgHqCbzYMiSTJ19qhldhRum6dYhk8zGw4y1vDwN20fkND35F8K
bNqMJCMiyVel9SdTbLPsfxzcL2hD8ogybyX77BScSUD7EI6e/TDfT3tMYovOL8OP
CxBTLIXPzS9k+SihAg61dXcFFwJVLXUTvT50iLTf6LKWOakExDNxzVuYNWIKvWE5
hsGehHpPEi14Nas4j9Fn1T1w9T0/cQdWsxh7FbBs72Iyn5WFmckRa2wrdirk8W2N
CtM5U0o4GZ4z+CEC+36n1yJkQ29lNJh7BgmWL10/5uPqvD3RH5EuxhzCoi8oWrhR
Q4pZGm8KlkXbLDx0mDAGsnqZAXPxP8un8lLf9f79lJGeXWk2cudSkYJ0DgZzoDB1
TUoz5pqcB837T/Yf9FoPH6/visgMFlHpnIsN55ZSYMu5f22R3gLbmN9KAWycoblz
lV4bBlZRduHdLyikQT6PtfOrDSaLv8eNeFrfRm1uI64/fMFv2ei+C+yTyOVSmjrH
5zzt/p81yVn1+Bphkd1b7MEkk8rJo01Dg3hyDkQyUI6uFYgi6dQ2R5pyuVfkQVH3
Cu0z94V+WnMMNJuLCsqwBDrob15qvwrWYwcMAcaa8ae3v4Ip7Z5ro/yKWC0ktamS
bbxQlWeaxJ4C8KCoRv4AS4fd9+FUk7MDiOC0JsgIuLwqzYovoWoiS6Xcev5C5KxP
5wUl8J9XSwtKuDiPtj8qxBJYAMO+Qb74+T58Nm71fDn1ocw6CbwwFGHKh9Cfp/2W
/bewMbkvXN8viIKumcwaU5cCqkZ7C9Ac3shcf1nhO5jc9Fp1I2UEtNp9KlNqZ3bx
Pmkdwq8UzdhRuQ2nDn4kKHVs25Ut19UAP+PlwVAT6AyDaRUV3EuptFgXpjA29DpG
clqjjljucuYqaCqFzUbriZMx1Y9B/kgdfN4TDz2Hi0IJ/m8WTjCptktLoqFzpEaG
826JCWfD0EoA/0KfC89sAGocZgpw8kdHCF/TxMRzixW5ikhv40BCD0TiqNKvtkcT
tE3JnOnPoRlv5UNvLCgYm1M/pRkVuWpnoz3hYvDnE6ZYtTBcgYX1AXQiNmu7815C
JM63Qg97Of4Zj6+zfhP3qHax6syDzu6KzoccI+6o11qYUYyfivRvi3tWnZy6NQek
T19Is6VTPaVyY3utowHhJ+B9i+I6qMTHoLZcUe2sZoVxOdjp4TtkCAJN8rVQb9Xv
Lo9kch1tuKx0uKYfFgh/dRyEnslStR8z8Ow33eg0t6LY97vXMA2kiGh4MButD/9/
T6vLJ459dkbHoeBH3C8c94IE9AxmEHZkT3wkdxENqED91eTNgUcOrTDTad5pbMop
LQBcQqk0V1fqTiUWuCXowvrSC9MaTDq+wgoObyEKAvzsBoNzp52Px7MWEWi0+hTd
S26eM0RrYv1ty+qNj+EZAT/TEMgIX7ea7Ti4RA/wBz9SAY8ELjoWrmidmzvpaJX2
xV0rZK+udX1IIMKL/yUQvvS6pC1j7l/diMW7f0Qg4x+bjvwVOkTJeMoepKlEqPSU
fVqI1twbc6mpBw6UYeC5W0bNScHYd83tKuKRqz4kk8Ru+rTvSK4lQdPN189xoXNl
/LOB1tgD+PSNXb0V4udPW6yvEOZwoFGQJJVM/LBxEaN0UZLN601k7PFEuXJLVhRY
60kRyetB0kXk0ZQoOYQOgySVexjqyHavruNdvX+xiqBKFl2kNadzvAbBRjqdLn1d
MUQkhdk2BXT+xMWFXUh+Rsopbc7ixmG1Tk09KTtzSAa14Mv25vQiW23zSL3xzzyj
cabZyXQSKbpJ5eiLg/F3cVOyENN7ksUmlkAg53sVnIrjU5ZblXInfv0z04aCnkiT
60i0o95jCnIqNoXqP3OjWvS/OQrW/zY19fP93f2r7b9tUNDIUqGOo6qY6mSYYo+5
SSNBlSVDSZhaS5k6shEab14yh5Bq/xYEx2NSJ1p00M1nVoxwCErlZuBB5y27uB3t
Xi/ZI4Cl00Xl8U6myr9psASUTWsKoFAzM/D+9rjPUvc=
`protect END_PROTECTED
