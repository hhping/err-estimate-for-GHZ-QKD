`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
32ztgWzPO7I9Bq9tiNqWg7GFJIJpwh+I4+/Pt721SYz7SjXF79IMqH8Bpac2hUkr
WcXbviwKzke6IqelRqjxFltZPlZpdKbV4QfCN5zzkrVDfEFAU1ovqhvPBiFtMKbp
9HvNXwM9yoUfDP1MZym5wuuDXT8qpf7hb9dm340PiOvvWe/XaCOxiI8gmMgroAXs
A595f0CWYe0nUOlbJ23XkIyaXwiKmHlNkLaod3AMpI0Rgn6kfi9d+ZJiR6cbqkGL
bg9zMrNlxxYGyjUYLs+ayIEA/890VIcsNOgayjoRAyDIi37nH8Yq5DLk9yGmSGTe
BRJ0Z21qC27oxLUSJUBm7oleehstCyIA2621ileJk2dELRC+ggmx/eAHr8dj7nVq
eHqdzYY1llzd6E+xV1gG2A26k0pPod/dflMtbGnXz1piFLyWNvP7T2W2bXEDHnA/
GJb37RGaWitoZN2gy4zSXNW2jgqCXYDt7XB16C72OCZoeVQwOuxOMYTPKe4X66A6
MyS2Zw6wa5pj1xvfrDJwl4pQX5gpijCn/8H1vhhnSBEXoLXy4HGPmMbyEpI5FPUW
HRasljY/tOSTClB7M+piAKz/wJREjZad5SwLH9vzQN+6j/ZqnmnSdrEVCMeeTMZQ
XNphqN12bl2lmtyO2Cfwn5S+1AVp574m8r8CW3R3ZWTkkjo+pUv6q2+DvX3Xtnfc
vcv3zCvdJwjJ/9s2nVt86LgtlFw/4AYO1aA7hZAkZm06aSkzivTjF8X6FobyveYJ
8HE9nAZ3FmevgSJYK8KP8gbVnVCN+ELik9JxUuY7sMCKJRa2flIIcOQoEOgu9Sq8
BwAkOJvVLI2LMvbJ/FnuXuOuMH0DIjpDQrs6tNzx3/6gATl41cDduU0Z9M4cKiQU
No2Bp0uKK7PmN2ZzljrFQMki84cGNCYZBJ9aszIWPuaIsB0FGFPjboYgv4NNJ9d+
l5DPQRIoYnHkG9r+IdKjlNQaANzE5fRx9qb4Qh+k8/1vL9JfruwtUGcsiiZZ+npR
kXbRR3VmPCcnslo1QiDh+Mc74gBMUjwWgX+/808FfpElRs/dK+PcFjQtrNRCBhfu
yzV6kfMD2U5y8kuY9/vLxg8pOVuuBJgfnrEkP7TrOS7EaoTGLx/OngHDqjeWedSy
hdVHYcVHTLtUfzfGuA3ayQMnHoPYLyAaYtfaHts0+5UaPC8pPTUvLUhEO7240ZeI
y9/XaAcud1r4JPhfObAhbNfss+9o36blnT+CDbdRtb4r/q51kpEvzbrrkp0rBwUe
fZ1EJrCSrkqBxINvm2aOg1YEjIg+jcvFV4Bsyt8syrSVAMYZ5g7YghjJepnTK716
mzNlu4zvTwRtjNs440vx1dc77C8fbhNSSSmR5pcQPcI2Ztv3g0dWtfMygGImvTDY
yPIhF97qfP1bud/+xOGTotX6uXf2LDsNbymZaQbxBkJOwK1P5DsgKBuY7VHsYc7T
wPY7APtvqIgNcKyNdSG4WVNs0K6/Szgu85RLy7UAquu/1AETShw5GYFIAUTPr/es
mRt2yV2x4xvaqHM4yO3MMa7mEXT7qVY6JAI4y6hH7ehcqrJdkU/wbLtJT1cl9vSB
iICKPCu8IJO7asEDSPoEvDjmb8XnUkkVckdJUCCqtQv59AnF2H+lIObjs0Xn7MHp
rwUHT3Qjjn9ld8QRyxA3d4PbKIrdBKcneqG7qlMPLfIabp6EHNRrqFvQXfoJ7h31
I8pcaRK53XM6sVpOxOri8a/ip1luQ61kCNfMxO/yodrA9UbeZp5Vjks/UCbPLjFL
UoxG9FW+twHnrfGjji68D5Eq/Adkib2+ywL9yRu/1REXVWakvVKNaSic7nrU/yKn
vGELmw9FJ4hW5AcHKbeqcyYp7oPvdjc21CGh9T066FHdfcIKGuOuR2+jt1wJmyPV
KreZS1MCIkK3KkBa8Z1LiPZSv7Zzul66WJNni3n1tlQld95BprlHu0t3aotUSoKB
KS9Q+B+Zq7nrZzZuKMNKPJY/nLQGuthXNuW/HWwo2ZwQOYbcZn5RRx3R5JhPyX4r
AJpedKiDv42DE+q3WH2zOo11kR4IcAL77u3M/gCCdqimz+JlqPi0HFEpUdI1WzSx
5E3rZ8DLCFDV5B3SvEJjEXvoMfqYCfDQJts2pt18LM39IG4hbiXJMOUrofao4lRp
hQB45eD0Dy09cckc9JfN9BRea22bDDkR3mJUBqJ1APCtJJ5iYPBpE5CzVtFnDCLk
p4zs0tyiyQTwev33aBn2ct0oL5u2vG6rcZeIihASt+/lAnEXlDdRBBhvsb+1yO9k
OWc/S5xeXQ+qncZLYQt/ow==
`protect END_PROTECTED
