`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
scqDxdyog9pHhb0fuNVHjXCCGwr1g0Qd5QPqx/unmXcGgDQMs0hc5hwn7aZ4A/wN
QwrYuZiyRvTkI+PvjJPW5+eFOIgV82nEN4TWSZ+L5iptQ4GnPIpnp0Z1dSt5lY6j
dnkJ/SCbiJF/Dy52n1a9guUsHlki+qK+9aQCnLoluhtRSy0c8ng/qHDJA1MKJLSo
ndCx519XGj+K0aaIGioqkOLd76xTWCun/Dk8o9kwlqIm2QHf1DvTuwKUM8iupERc
f+JHGv/45/FveiabjesAz53tIPCQsx/n2y97P3xTIS7ZjxvOpmN4Twf/3wIq13Bh
EG6nsSe6jA4+GGQSox0zVCkGROj21g7mjHY+IFIExfVEWYAxXzOP/PSwrONsHvrs
3Q4wOFY69iflrI5+ZOYiDsC98n6QaKwU6IakI2cm81oge+2YPUdHgcZEVpPrT9E4
P+Mpxalu1FnrCyl3OlSC7h17JwAubWyvQLZB6QAm342ZwIJAs6UOTxrQZEHLPwst
rUnzM6Nb83AWEzoxw/mnbfpnx9vsLGCiaLudKZX87S7yfI9Hzbhs5v3rx/O8w+HD
q0DCA2jnx62pXQNFR0RW80g6SX6otDJ0IYHpJxXft9eTMuuf9scxqaJ5qtrqNUSQ
+EtReTerX3KKNu46He98sogTZSEbDZI95e1zdqBRFpmMSDE1jW7UsLYvSCf4r3s8
GLYIsTPKeTmIbuguX6VrsNgTjA3S09MD9j7AeVUvog2JaTOfNNAWnUMH//AiY6EO
hlQE851e7/V+cr9Zy3AaCWvA9E48FrAQc0nMaJBMRLexZD0Jtjog7a7xcCN5hJf/
/H4siVA61CZ0OlfN2m/qXPWGHyOYtm5sUvmewdLBbBlW0xuscz0y5Cy5JxjG9qp1
8VKdX+dQHeMFf7JciNcEapLy66q/dtY/0GpuBByjaBtWlpBk7xeRo8lJzr3zDuwo
FhItrOe6ydykk6g+h977kZh00z+3Tg/zaCfrMeZ2405H15OaeNBBr0Qu9lOMEkfW
N/9kryDuLuzhhOH7MdlVkftajeZOHUJKLxuLG2AAKJSNs5ha7tPHX8dxGPfgahMX
c3wWx0hMwHTV6IXC93gdPukZ3xO7z1XmkFv3UEE9IsxOPiH5pGhttlataptf+fFj
s7Pxa2+1jUov1AoWnkHTGgwR2RYjvF2chu1hZFyBWhVykp4+VkJxr0WpmbADLcPE
Utf/sOY4IZK0rkJJupY+z6RgM9ft1CXdGiQN4/zrNb3fTuk6E/kxP9YgQzK5EF66
GnBs76K0KkPpu6YrUxo7+VsiAEexpk/PJRmrDP009FZd6OfNMjKq1KTIW5c5R0OY
Trt0INn795CcyPgsVhOSTh3yv9x9EIgKFEYEk1LJo4KEBvN33DM4G2BZ/0oDunA0
ZB1SCPyDaJTxRiBsHHtyOSUfCESs/iJ54NY2mkJCVEkCqYhHLa2frTg3XOdwlgKt
Jq1fdYYbsqq65ezk16gayq3rWs7nSjlMyVq1W3IDtSVmefvsOm8u1kDBsR7ZCD2f
nSS6s8G7PAwbOX7lA6Tw7CzTefd+NFtutA0ZBlUVww5Ypioqdv2/ueU06YMXYOc2
gPPdiFtBOzf1UKH7edPCqqQMdR5wM5fE9pCBRZUWew4YBM245xEi+u/XiJlyr/uq
9eoekqKnnjfClleAtv4C9/Uo5hMR/NDg/XX372e3pco9wq1dFOZzeOaRYcfqFJkm
EJ+L8rQdH36YwIcImAE1qkpQFziRRGtm57/2Jhg4Ph8UslpjqhydYm6k9Gqf/Qer
1bCQpfvT8xURZPb/FPPXDfId41nSsCIeVhXYiIF7ULHc2y//Qfm6h4wMsywDoGZv
sKz0am99TyzSUmyoNl3Sr3gwdGAF2cEd8sIQ38YOnVZjgLUO461gj81u87GGIBAW
lLPTtkPmymNm2IsC8VdHd4u7g3QfzR3AdWXJazTrgAIh5qiWN6njK1vCOcgVwwZs
6PS/AwDzHNFdhloKNc8dhrJhp6XrnMBcQcfVGxyeXQu0WVONEUFHocJwPB+1AVBX
AYTDRV36DOwwTpb+TY24dMSjnpOxgVjidwozD0X9iY+3R+CzFhK6ZYpTEaiimNDh
7tkYml2alzf74ySQDycEL0CrTqbpI1Y1q9EoBh4UbXVH04AoPbKjJyu91e0tKsTj
En94lBcyRWirEAh3zjY1ydatBWJWEVRHEflK/9YYSVUUE252ppCT2JPJxXoWPkz/
LZL0vIVdCAiy+WUtDkhcA67kJEJ5mP2oLXz8b1a1Jy1y7fS/Pd/XNy6L1wJ94C21
p0WCpG7b+pazLdkHcGgFIMxRVv9RPDUMEJC0i9UFkc39mxTwUsZR94al9zIgUrye
Invj2K+QJ07ytCsDfZyEfYa7ddU8yLk7Jv5CCgnZQjupHyDWijdKDiVfmUMjkvZe
10xhAb4cjSv6evr1V6cl1Uj4VorTJdgZeWDR/zudBYzJAqdUJ6UI+rRRglIGhK8E
SbSLXw8F62WOETS+68PDJLRB58i/r5b/MlrZPe1f5OQF7VmXwp1xaMQY0tewdKTE
KLu6ffqUZlL2PjMuYT2nG6okKPw5Xm7PXQtjWCkSbrS82CBgAUIELBwq5v3vehvd
O+UMj7eWQ1VlL1HRyWC4RddqOPKS98b/QSEjHVi0Hvqrz4d3PlcDecvn0+UyZ79Y
m9KCW0hG259DAMH+iFWtYHeONEoLcKbu3XDMyzOLE9zv4gVXsQ2yjLYbI8VIa7T+
FiNE1a/hXAqNHBz/u6KCx/7egTuQr0s/D051LeytPvEXNNHzIS8EgiXotBHzO3Bm
TCJPrRyfkkgJnN9rWTSdV0m/qEscYRiLtf7ib5FsAEypYHe6fFmR0BJSS6wL1FXb
sK6TlwKnqOH3Q/reK0EixUl7c90jPrvnuhMJ2qbhnid/JKJej+1pNgehHCxlpZAV
fj/KmVSTQRReyjRpmOaPOxTfZn9DwizezzqPB5lsCQLlg43if8iSY+MR5Pob+4H9
XG8YYyJJ89gAJXubMxQHzwRB9N1eAtLcDs+uT2lAFV4wb0aWHQnbbYAIEBiI+n3H
wSRVtuRMIgJlDhSP7N8Cyo9YptSeUsm5w9u0/uU6u0euog/36iGCuxvb0vQOeBE3
LEfONaxGoutvmVWQJ7QFX0cexnA+F7T3W6kSKTG2uiADYPy4rZKoSlruzS5zSUMR
83O+ZjFJgwM+ukiZT9/O5rkGOGYLOV3kqYoinXceI3MlGtqTr52QFPdvp65l48PX
AH/62uPaS+1ySBZLkVvi4rbpnmiUL15G0Kgiql0VAc2VNOmCVgXVChrK+dgU6D+L
ymkB6/UTQ7tVIPXq0Ej9JQpuk7lTD/iENmEsKsM0HGPf/214FLO5p2rUMVYXQcAU
LibC5FGVOe734+aIDwowAB85vnkgZt6HexOZgalvTqczJaGuP4IIRr8GZ+30iXHE
zM328YWaubqy0rAAewIWCeutrS7j15lGuT0vS+D0MSA6WtocxSjSQBay7YjHE0HG
pi8e9t2cyGZH1USYjeuuMwBRZbNuLfxS5OxRKW2ZZIqT5/156APaTafGsXtOTGCK
WunaCKI6bBmYLodxL+5WULvYaizgWKk6sVPv2duaQd7Qj8/UuZnH2xgaPgdMsMe8
VyTQeDPSKrRs1dwbjBMjSKNAnHarGAtWGmmofWBwsi02app37y36yftXHAM4KKww
ThMHt1607sCTAbzzM2/F5VkeGyLnBYG5oc8huIfXaJTy0KwEd8gJK6fkHvv4Bo5n
/EjYttZBH1hZiGQQLWEwc+wYdLnmK7xvSTnceJbhf8JFdCdHpan3B/5kLtqwaAgp
wf62HyncF/Cv4OCYO0lpBkxf7a0QTUEaj/gqutbB/F8jdtJR5bFE0wk6ZPF5/v6D
2HcrxBPBL5wxBJ9sjM5aPLrs/WBHG02QBuIFXFV+YldfhT8soDklNl7m6M9JSeeI
TlP3P+S3qFnNGlduCKfxQ25f71oiNgnq6rlxvyKoSt3r8c4+zYrZ/wZm0lKLDUnH
zGrV/2bKrggRRSUtXtjGb/mFZ0XjbjWP2R7Ad5sh4y0S3j7e4wbMYV5QCPmVJCXQ
KuHhn9EMdHeDOqA+giPJEA8Et7r/DYgs2STlonZKxPK90IRFqE0EIk5bbUWBKzAW
5XE/Z3ezUll3+l5YXP057WDNX3FtGG3avL0RTvdi6nliaQsrkl2KzxeO5QjSAojp
6v08k96HR1S5Fv4rPuEygXqxwY9fBezvlyGxlfIEBAA0B8gcD/h/5hXIoXyHYqOA
i4Ie4Vmh/6Ne6G7pbAAQyKapM49EtjozH42rqMrLV4qus4WnOkzHJ0Sda2uUjNFZ
j+UJ1FYSLoDCVEEFlolQbZ3PPjg0dncGZyuSdSp6Cc1Gg3AuZnE4ampjl5Hng5cq
c4k87bJvQ1uhXZl4qxR/B/ur32s2rgCU2J5EiDxmmoNwsNYUplZyMMkMGrDkBX5K
oXofeNySiIDc6GxeF9ra26Uua0Ur+LYjX9+e8qyovIQjwZbBzk4OPlOgCsWKdAgZ
utySbDrj5qQIiJdU74Niml1HH4GhT0AWuELkyKhR3Z/jkON1Lv9iaQdbgYj+6s9I
ntz7gqhwiOnnA7LiiwbRl4E0DRmb3HbnHgqeMrp/qoq6CXb3tyk6LWuqI99usTXd
VLWfqqC4XkHhqlWHDhHXyCadYb7JnbIyl04UVi1ADVAMx7OZWYmqvX2uQh3Mjbbp
7gbuz/QvAc7sM2Z2dVgY6tnvd89cH6llXLvhMCOI4v6jRKwZuE11SwY3ke1p8WNa
8RcE3VoF35Su9f8Flkmr5UP8T8St1uOOHQ33XCeiyIKUqMrrKEKnmhqCQRsVoA21
AIaQnvwwO2mwkb2DVgQjX6L03POVUW/+WAgELP9qLo5U2Oq69HpE5bBsrmYEH5l2
mSLybmiZnS1i6rrW0CDpPgFqkE/BBJL8hqoIfHu0/cEBXymf3VXs6Kl42d/4V9H8
Pdi0nuLvP7GlMfVjq7Bnzoi4qUP8edoIU28j4nMXXakrD7VHrw0aoLZ5iHycW036
OSQwkVrIRfQXOh19Nox/GnNk67ngpVwJLxZY45+ogmnHOnNJkLEOpd+Syudxe3qy
hZf8mF6LGuCWtK2hkicoWxky/selUFGZT0PjENKwo//q6MxTIFFixpO5vmMgiQrt
FeG/iDxYL1WzOr/T4XZeLMhk+LP/HQ/7rgOD28MCOwtO4eOVaDIhVF1ahuWyxVZw
zedK7DbY0fwAIL60z6aAe6yFjqH3YuUBx+CEUm6hMHSRmWQ5gHUtJWmtpoEyPb5n
SsgKOGwArLRwbNDj32jUzLXINKGVLQsk9Yyol61+cyaWvLDmIy5kBtkFClzYv3Wv
pi2X7cX9DHuCA/ByuiF1c2RoXQ93IIyevZsPexShBH4TaA/nj+iZ3YfxYkiMRzR2
Ex5G95c7j29ekYBpBTZ2SnAAayAaJv6kuMkDZbvFv5vRLFzy40JV675fpnELtS85
bcJnWJs+wIsKDKla9agntEGumkwRiV14IRpiceeTsPwj6fTSRH1txo47ALWYm7hq
qVZq/ME4HAifnb3hs3mspLO7FTPvbq8VsRwTJaMoqH856Gl8BbanIddCDeaOGmPK
OVAEJ7ujiO5TClu6YUJdKGOkvBntmGPfdXGIRXBtXQ1hcGz6jW9z/2nIlTbik20j
ybaAY8kBRPlPbj9YtS6O2t57mmbV+/mtvpIMThxM5pJIrCoEgMpstUPRB+U4UNXC
UGox/E2Z+YssOdbJOnZ3b94ptV3MNffwZT5nOR9qvBZKws6R0YTtrxXntUWa9/G2
PriGQ/u8zKhvL8wWFFyuE10wGaI6uAzSkRNhtMsK8N6t/fT5yzINLM4Wg5quVSnD
ZRNduMFpBgZrMkYWdGYhtbdDGWehuUFg0u0lZ5/rM3Aib5BMtFhGVK201MX9lad1
Tnq2/vuTrddxCRYByoXQqfSkweus8gYv8bSOHpPrC1RTtCFL73Llfaci6NSPZHqq
NMm4JSse+sUTQgTQqExt6gz5drCVUR8BkV6vPdSQJdQYWuN9g64sQ67H/wtu5nJG
kgdxnMduRzVhsV+uJLf7+dLcyOht9PGylQGLotSTpvfJ79D64DXRtbpFvozs+ZFz
PiuE4LGuypw322dnLBnrQDWBCmQqlj7gYQ/+KVfNE0o99cZCe+tXfjw6+OanRw1Z
hF+dnixNZCM2rXbbUC3YuqpGtMV1ONuDPlaQ62SQWrKk2Czmz2VBi0eFtmw4z/Uq
ullmZGjYDu0ig+YniXPntS4NxgSmzfjiiKz7lpL1zjevYx5Avo1pD0K2oyNEcypT
fqoXOD0OlmvW4vokh0wUIJRRAjvjtuR+JlzJOtT2doxqnm4S3EQU64cV4kcFp06G
S1rw3+MxN0FDxn4npTE1NebVrgrzpk/9NuIxSVrhVjov79Jqv0ncdQwCpyfH2K2H
ST8II0lIuc1IYdKA58bgm5LuUmFcSedZmusKRFFet4cdCBsGyXqiKEzNvw4M8wj6
OYHuCFZuvLyMSVo8GckyanYgqDotBGtKaSx4PgX6i4k3SEMetuK+25D1EzwiZJ77
3O5sxt0G0ZFtKDeTHB1x9RzypArF+2pDrV29rQxCi9osxpZsi+zbrH2e2/bS9hnP
nyHvnp6qKTB/8lNq1fTp6rAy/o4OVWixiR5Tx875pGAfn44Mt3hJwsriVDcyfeZ1
T8y9dfst6XLOCKVCKm78UHKY5IH67JQTJufh2k4lTN/aSexgjjp4VBkbAkKRdDFv
xogvLMjgdFYftugROCyx9S1CqwtEjHLEI/I5tIpXB2VBemhaAwqaVc3BLFke3PwE
Z068UYdCEQcbQs0FmV8BHJ4mZtyo+++pvCmn+RJ1Qe9hidGjNOn7axzoKGAigeOg
LwPnNmTCvuI3JadeIG9t8vGONKFrom4Vn9VsXGcid6l4funB9pA5O//UqcpwDB4Y
NxnDYkrJvnA5O2VRMMpEet8Ds3Z1elYXmafs7ai6yDR1g6iX/9+fGiqKiDyWFlkb
Hj3qQkl1HxVDLSQYfQH6NDevIpV4O/NabfG73tae5IPcwYqeyagZ1/QhSrltwyzS
tB8cV2iSyjtqFWLOKtr6CrQoCT/KvNoI4ibRAenvyRmN4LPRpCFyTCFu4XjeYeg+
w/jhMutX1Z3y9QNCHypSW36CqTzdLkrhe9Ut8R9Vz6xibEKxbI9TyqW3sGIWgtV9
iZtNbtPPZsrsCvz8Tc5mdXaOlrwKO/CaeTxB9CbYjj01n+ZY1wczptizgID93OAI
AyUiXKM/08QV87NezWk1u9RFG71m/WQrqV6CS0pIXrSdiiySRMjTWtzBlTgnYMlO
kv13BhYDxkGmuyq51PZt4bBqgrmPhZCgnANWMrvU6ygvWLAr+28Kot4P3oZ9BJo+
sQS8+9mzSCnaSTWvgTUpThn/SFUUhrYQopeSR27Brnd01Bv0V3gRp5QdEHu/xG70
EmVac7TtK887NRblVfwHiVxx3ZbQMFq4ahCGsGsOYXjuXuuaoyUe5G2kLfRL3kWf
4QCu/esloF0TSmh4cdZpqNsH2FKy4cQqXI1/Fh4ClqTeT/37Q3NcLK1/Jy9f7go5
uBQ75stasCZffh1hb/KmiMmkYQeLw9btzVhYae2GtOn46LOQ3mxdrZMfzwnRNMOR
iF6E5Ewb60sVvNz1DVKDSWZcoBXIYC3xyBTMFsumJpHdj7PoxLfawZcX9ar/gD0m
5c7l0w9kdyE46i8sTGo1WkkDYglg3uT5MiVWDRwI86RAYOo0RcZfTEzScmWBFgKo
I2IFPNpjYzd6IPQAfgcrbm1Y5XzbQNNBb1b/MY18p2sR4O236ZmgL3Nxn/XqDpN0
hBv68C1vIIwXbPDepZ26PPfUGwYO7MrUpGW1ojYbESQzzOEjleSy/sYr1NYFXGsB
3urkm9y2uHvAYeK17T8FFfuEYquML3J1V1MpixtBIXR5DLD2PC5qagOZcXDL07Km
gZNcVMQ4WYpiRfXAg8WbU/eC88NIEvUrPrDFaroteJt+6ISWoTEEymTMgkAtO9W/
FahFpbU13Q9CTI7t2We/90PlLVN2oRymTsT5ZSFf8H5AbgKJRqccaw2K8kOj0SkF
HVi1lXlafJGotiQ3Jaj7rb9Itiy/J6WKk6WdG/tvcSNtXB1r0Y6YwSjvHrOjSpnR
nhLb5hSnLFoIoOIZcfceEfjUvrVnyKAm5+MOE7cAHBY/VbfMbkTETVR2ATEZ/gt6
+4V5O6mGYlmwfDhOsBHbvJ9IxTLuN/RaiPXvhFTb4Qr3557L/AiauO6wQIGYSh2C
7/23UTKKaoSsdpHzrlOWege5PzVzv7nuLozzNtbV1mNcyYE6kt0B/iq2+5c+12C/
Ot+2L7nwNqf8WwawCp6pyT0lJYrlKnuwTeOub/4DrkB2cNaHzu2FfogsDlwXRCcs
mbkfimXt+dv3Vkkst+QGmxv0aB6hLeoEJCmSAucdExgn06FNpKDhvOE8yKKWxtix
mI55XJ0LZdyE1oDQYYdSRaKdxlGLNtrudElUUPAdjoDAqew83G5dkWd3AuvRXSYY
Zt8EPWLe9bZQ63fvbcbh3bCpKtkYEIpVagjNTop1ocW2XY9egEMiqGuI9i6SPYWi
4Dr6SFCcU2v1w/0Uxf6BSNjoIt3KHiFjdodjOe611AdcsYnsX5y3DaOn5/edW6br
3+xSfoerLeThlsKPO3ZdXMWUJG2aD9pp3+y17O+F/sqnl33SSWDnW1ypADgsJ2WW
6orwB7wTvc+Qj2sqazZdsBQ2H/5is7aZ3lJWKM0xEbBiiFjK4sKQFnaBa+/cXRWa
8hIWbYgcJRf5Iq3k/yIOmRjZxHjeH/wmuxSHPxHmqwR/Bi7EvxqewOIHePs3ovie
7h7XRm32QlLh47jDOSad7ZT8wJ1xtTxXTU7A4lI42qcwWTgp9Q0HDUZvqnnFeWhr
g9S4X1v4oc/hMeOVaCBFvIOX73BAIYBj7flXGAhfivyNILsMq0GNjjQAzgOpIvrq
5Q/J9Zwq67642DbiPsinpDdrFLWlo2jCry1QjCj8crejADyoT08U1D1i9/5JmszF
X1SJhOsVDKFVyG1RwtFqJOYKtVk1XSIDR/sYaFwZVWMSvDBpzCrHMVik5vgGfyml
dIHPblse186iZD3L7u9PAaFkdQMSHdcPrUsXEKioocAf0UiuK7OXY5zS63n+Qcnq
hrFxvqCjSBkSnjQVUIyYMDcCf1+pvqgPYRNZOCsd2pa2capxM05f1qD7Xiu0s7V9
mSdkQGlYAQSf45Sf9rPTxLSMqOxELMf6cXSpobJBy2R3b8GXmJ65W6C0HGL9Q9hY
g+K5tG+r0p0XldOaBBNjd2AThqx1co7EN9sgXEqvMI05c4JxKZJ/IhNMvt1V12El
/++JD8GNCwrFU5hUT1IiR2/UBP2siwVdepCXyxuohKwLdyGioZFTZwqdIfpORlSC
Nm11EmSfleJBmaFmDJHF/CcL/zwNQW4Q9E+z5oc9bDr/LcImEMPbQBCIacMHp4kd
D33IDHmEnJrFSwKP+g+tJavFD1SkrJDQthm2OIQOLd+2MfnsMmQH4N/srhfpsFtg
QsY6wwZdVQnZM6EJrLMNAwvFldYgiJggdS3YN60W0ogJh2TGYYJRuNfaTeaOMS21
g3JkF1GrYTVKzWQpI9hLYFYvtveAq0hdJAX/snLkS7erWTTX3whikE2bt0phH1er
RifjJ+hOqW3S6GaqkTVl7QgOKAtJnCXOX3XRoI4ICIzYLTOZo/G8WSBf5qEQCdRG
7gkApvYCl6XXP+t79mXxJ0dgzDnTS87KsPwH6ZVF19L5+SSNY5VvTARaYeT4fN92
bPHVyU69j7b799hqRdRhfkHYJ1UCkv+82nlqZ5iOIe4i3aI71/M6Ud7VX2UQubTQ
849wYR+v29XyUQB4OqYoOJEB1scN9Mrg/5toyfEC9DgckDmWyft1dkhadEZZLLtX
8nq94AxXnaqBsOcSrJROhtttjKxRoFwhJcNSOClPNcx/jkW63Joc982hdsV/FEwl
vUzFHQfq93g9rY8P0c9g3nm7iXMY2Z8o2fObHCPqjJqcBka2QfJnlDDihvtv+SQf
rAmjNMj4DfRT0LdLfm3NqofBlHJc+4Z/ERTY4llOOYwuXBXQxDP/oDLWZDfWLKzP
DeEdxiJ1fa3Kv05nzYt7lO56B/TIpgJ/C3Yezky2VFZqDXqzPPC1YO1RwkR3yS8I
WRjTeOoHD/lB7g+dMz/0Gs26dcp5ijeykolDsPf+e8iAcTd2JC1fQPdll8U9mnQo
t++DXO+y72xlXveGN33WWPt9NAaJyR8mOrvxSVoBr4adqD/DV1eSeTcSHnn6l8gE
OSvhEA6l35xTW8f2xFuFd73xHeFt4OKGDXnOxlVy5bcGDapBrXy6xf6kXbLKjSli
IbO5l/APE0xotDX5IxZPYbSjb7mXrI1KuTivThWjxvrInUne0Gy1qAwVHH3q87xD
ViqJylWfOuC3Wnb2LXfrKQMLrJBNC4uMY59B+7E0UbPNKrGBj7ut9tXGtsyi/bh/
wLUK5pecG9bUr+X4DVmqT56Bn+B/cAY7W+TSGItsa6lDncujlHpaFPimpIM67b35
hTsHkr0GcpR36c8M5mJY5BrHnVAWFy9r5Zypyo/8Nl1oDkJfy3F1fYDxmNelTMy/
SP5iLonJdB47tVtfZpUrfZVoM/ycYZPWmeIMs+HxmAAt1AHJONB7dgN1gFdwIfIq
lEnzqXKvJyuSvZhOAijaiZbtBDq51I+Z+Wf707AMHPHt3oAbSrI+SeX2gcrNH0rM
gRvuu98NLmKk7Lsyw++77u5fluIEV4EgOG9HJ3otZr2S5D4b9BaR8oI/Pi4cXM1N
TdVauSnW4B4T9oc8H3DTAVmK51xkmN/7G87IC5dNgrX5DuOlFuAjNmL2NX8ZrvNS
8rkVMza67wP1LVyH9GpxRshoEJ61qNhFcEv8rYRvtLizzznFxz80ZZqH6drbseHV
p8Qwf0HuWMVU/p7fYHDin1LrFKWpVzxND7Q4kxPiAfYA8X/KJRdC9csNlGhcfCxV
EAGoKpAgiXjlQ1gcvNv0eJ/Sqn7m355vAn/vXMnRzilebYRmFhjolgKvUyVvmsX/
kCdCQ40pUCsQ8KQEqk+wRO4wBGeEKmUCvmlmwY64oQEoT/TLnn66641p/b39R41R
6tiwJRaHXDqdz0W4MOeYKZSCtEsOSV/xWH6RcMXD9hy93n+maorITzsrG/MwEzYv
PucK3Dr75bKQ0+cPuObIJqPr/cy24jEizYpO8RtCdk50hTlPDiAgrA1IGl2sKHBK
tfrjQ6Xm0S1iKrrsBVUJve59T2jILE2tmE32/9ILHvF6OqcHzahxvMwSWWtIZFfV
CRVf4pD4KZX0TtQBqHmzZJrQ8mkZ/hxbnrJpKwSJxUOeZkJuE6mLHeLNshYc0Q6k
EHAnL0UNWdfHhCZgjWTRh0R1c51b8HepSoKqYTksP7UVhYsgRi0kWcIqSLYvJIOp
o7kt6jeFRHFkvWql6sO3hMk2mZfZrNcTQ4xm1xXTKYDKgkd1eInlbibeR1s8meLj
8OJWfemxKf70MuKZLzs0cWUqE88cNYOh71g5p/EsQddzIQcpe0LrPS7+hqcPOiDW
3x9UqnzkqK6Ntce7Z59LJGiYb2ECzNgjXzqx9cy8uGBthV+WOdX+hZDuOxt0qtav
BtGpccXnl+gqLb3adRQkGY74xB2kLmQzFRs4jWmJWYETWoV24M3XVsxSuVNbKwW6
h6mV1/bw8DXJcCyeYPLrwdOHMxdBYu323oajEIF+E/OU9hbSBN/nCsA7GGFtOXbl
C8EbymEhmzpfGhGmhywsifFvk/l2nvx0ETLjAOq6BmW9pBJzbs9wfQoYxu5yfAfA
Mi558/fri0wrNvyax9wqd5e85z81pXPW0xN6qaOJSAKBr6sz7bRU4uYIDOclOMK1
llLCVDpS/cCCqKlUzE0JX8HWvHw1bnk4+JoiJYC2Urx8XhRoXxXS7eEvru6YJ0tu
Rx94ZQI01EtPQEecIgpP4F40wEQRzBwfw5bc/WDrzvUFZTYJpjqtt/Ob7tNVuHDE
Duop4EN3HSoMdM6py9H9I96X1SOWSismx5mnRhHiWIMCAJy3Ld2FM7sjv8o2rAlL
x//odEO8Dv2pgxezUd+oxQ5JUSJsfWW5c0Ncg1nfkKsIM8KFR4S/kJeUr78f+OLm
5pfLEpWoSSu8s53vYHOrfYNCQAfrZKUnw67l5bgGIuOqe+qq8yHgt1zl2sL5gZwK
9IMa7jnj6uf4mlDwnVH7Lgv6KNysO9ZJeDIkUpP9oUhfPIRdJh8xXweCwgfc0PhW
dld3LJT0oXtpj+sn7+ZVYFchOuglnw22t/Kh1GRIxtI0jLGjVb4QytUYaf+laDpc
gvVBggXpKlT1o75ox0cLpadlqAdr46rf78XVmeCYx5W4aysMLo7wI/zPGG0Y7nNk
rT1jJ1rTQCKTaqqPyjz5PigP2sGihPRQkeRdFvw9VC/VaT2T9lNRUMeIe3GJSxdu
9kfv31JXYDaTxahxr0KTAapyifPm3DA4ho8/4VSmVoH/BxgVaZxL1XCAcOOM183i
MTxsV776t7iUA31Z9mqD/IB5EXXJaBf2KQMpxH3RfMqjeEsN1A/sN+XbIrABk5i4
S12XbNSxxD+D2Ur2ABCf/leSrcp+iZONH0PVvc0go2k8Ws+9qOIV/YB0aGKCaeV0
o3DAGhkPYvmqmEGQoFkhPx3spvBVspygHF7aUJgjSY4SJccjZgrAXZAmQ97ig9+5
uJJTApl+8rWf0+bnIjmCuf9o3IyvOII3OlETTUhk4alcd2IiCsS4aXgxml7nxNar
Qk97mh2gQ3a7dHvry/sQu1seZJGl9MzHXTpwhw4W2qTYoCUtTNBVCe3mYToOLGAQ
cChUIGUmpn/9KxOvSd3ZAlv+DvpDGRIGfn2efK4DD257RWiDrJSSVHiPdeER6Q57
ugR9D3CZdh8DNnuPI6chPbeN5hLJ3zVf1a1p+AtAkptohoX2Ttxio67kOhm5jJ7P
N9113FVx3+c69JAQoeB6tRtBd25XbxP71+VYE9tqsLDFQPuAiUPeTrWBGv7oUgOL
MVs6+yYGJ7IEmBsBHp5I2vOwD13nq07WGaewlEm9XGCZEUgicP+A3KDQbdWoRxPM
IPtCyHzmO472dyZPtfTIykYaciq/3AzmJahpILpFcWAluUWHlINOWo8WM55Txu2h
MdaNOHlrqswCGlEsQDi9LN+Lj3W3ZQ+y42ubmsiAvMDKUWyYMVB6xyqAbx3+75Xg
+13PXEVQvP0JtWHoLuE/7WcaFny4OtOSoT9xU/4VULqpBm4eIhcr6Xb/gc8RoY/a
X7mfqzc1GlG7PneXwHRRVrXtn/E95du8xgluoUH/A5OAhscRQEfrKBUWc/Q6sPZB
sQY8huQC1zxPLyuQV9UlQtF9vdhMd+6ZXt8kito1ijaPp0RUYGmu7kM4pG9kOuue
+WFb0CRDZnjZKu31haUNotSQqofQXaWLKdC8dsFUJ8M/IngGdj/2MTPFYFEAZi1a
JV439NAvX/KzmQr/vvzHzhC3kZZD6NxsQbBDXC3P7naKK3wqvJm2awr0/GE2LKUL
r4vK1Z0nAVpwMxoUAFnfd5mr4RXtvrthmlHk9PDvy5MZL9U9L1FKJTbHUQAoT0Zk
mnNyfzTsINyxw9jpSihDCOp/Dqq6EzQa3SZpKK85phnSvObWr9bN8g/s8KkB6gvv
4JlCimkvJXB+StJvnMRZCF1DFMl3znQ5Sam3m6hBeQmQFBCebrQyngB6WztUhphN
amR0c2tdt4HQkJKZ7MyEPiyfFyH6sxkTmEp7P8aVRbMWHh0F/dtaHnNQG6A3d+OX
eM4eF6W1P1PAbEvSvFFF3HAgnJmurKBd/SDfN2XsJgwrI7I6oXFRN+HnaTt0i2pG
yd35NnrFWPYlFfIatNTVAZb07ot/7qJCgP152vsGSM5qUbcd11hIUck1bmTrCwo4
G2WO6lkZITtzY0dlj3ce5YRVXSFC5YO1UtJK3aLblLcxpoCOqL5x6C42nKvVcvWI
4F+aH4PV3BT4mtMIgIB7apLOPcWZ0LcaKM8ojzbnlyUhGvT4jDM7xLc5oFJqeCr4
FrX+3++m9LgTnLmmvpXMviLZpM08Yw0S/efP6QogRnSX/ikJ9FhdpXDyxgv/2RHz
sPKQmuMVvwqpLw8ZxjkOcCGPy/7rbnkTUwWrcEPmKxF6WzlrTC8P3DFnN0SgGtOq
CYx7HWW7R6q51XVnh2d4LWVO44OTqDJdd4ngehqLaqmcOd7wb9Ak9ByKP0PImhKQ
KKjtC+bf2sp4iLb8HMlwCp50J+VA9rfFxB+fu6QjZUxqUjlGdPcJRohzc/kDm+G4
TmY6eQThDSmswIo2CW/QAevVIB+HDmGAC8S29Rc84zjAYXs3QLyyVHGAdfDAh5F2
dypdJe9FS98Jv/9R/50tPCoEA0Wp0xSNQM+2vMuyN2Py3jNQ2jjdtr/N4BFJDbnm
1tT4fcn8iqjeD+TalhyvqzQ93XuQJrVYwwcNjvBYpeMLhu0PN1NMvYZqhCpjEBPH
OhzxnWQRtXloexs7o5qMG36kC8KO+eHqg8rhQYM0Pu0pACnj7cRVEkluGrmuJcRC
sd0nYM6JK5k5k990+fKB35RghadNXLUGYb01MPdIhAK8lVdRlFy2K6hVdMESvXyq
3h+cQDlUK7Uuoq/tPMl8BzUcF9b5zMGGpGClgeMOk3qexihWb37ha/oZruTcgXKO
2dkeZkB6QS97JiFpzalq+1P7zu7qRFEpNSXHkolERAsEiPgYHl+9aPgYxtzTzqfp
NyLh7cavTDAumeNlQCOG46e9FN3pprOPkyyqkHvGTvU66Xavp3Ru3/4FoWhwgofd
ptSCdo5tqqyqZVHGvaZjAOoi3cmMGZWN9U79Vr9TFCC8Wwkc7/iin/tGt1nbmB88
RK9eKq2bbazSJF0MGq+92lU2SXPBNnsHjEuPcC6MijRXcrjyabmbn/XJb3/Eq7fD
r5OIxGc8LbSTcre7nk/L8JeyRfhailyZt3NGwjJGGtHgLb+OuoetlrCyvBdvPRh9
baInQAOm4U/PKwugSQN4GgsCMM7euH7ELTgaqLFQHzPH9CqgRK+bepbaM2Dq1IfT
w+Wwsfvs1F6HdAIM8BEwbyLEGKOSXQv2HfeYZVTemHiLr2aXvrRR+9he3vBciVTy
Qm6GXW5xO6kU5QQrBhJf3kEEWvKvj/uEeBkQcWcxFp2F0U1RCUN3faK/7BCf9Wqw
7vmV4uYWsQLgiRCPOFYVsrBBdkkKN07w/oJj11LfhENhaKm18fgRgurfd2wuPUSc
PPZ3gnQ86ZzFQucKCGzCvVVSDdBkMCpHjKkBYUGGvRaldyZpe/cbZEuL8Eh1YA91
WDfXhBGBySepvHCyroVxBss4XPB1gzLTcUJuM04/LcPKYnYzWR6PiC5vgVJ+Qc1o
91nvL/Y2Xf95omYAKGCDmQryshwsp+hGBEGydA1/CC+0fctwU6PDCcGbFHKma9H1
czI/naXHpB+C1ynyQu7sAoN4Uld8OUSczRyIWojYPgRPJAvYjF4+KWHk+jiGBOww
DJ9Y+jnSl2jpAUysC7WKZQS776FC5xwu8rjxMBsBVINve4nAO/4NH6MwNp1Q5zJU
/p/u9pRlRKSyq+XfRqkMBf4AS/3skrdADhIVfx0rNFU4uiTknXik+yBzJYJZifvT
HJTquvXYMnlsq0UqqrV1edSssUKComg9loRVe5lYTez9dwVP7pPWX/E9Hq+0sCOt
huPbtn6nf/WMohMwuYxk2EiJFyirevwzfujQToMb4Q5lQIa4kJcI3VsI3vJuPtip
B8TYaAeNw9xz619ZjecZbLhlOI4EJSUMw5N3WM+YNwIbD/9S60en/ewnGtOFcUiz
0/xidc3QyEdXMARp41zrMHlhXkg2J0+eWLfHW/btFqo3DGMIgXO96MWEtJry6cgF
T+ANMuQg2Rkd4dP80GOyjtYnBtzDb7KwGa86hyuurs5Z3CFgfNGKlfyTRCbVvHtj
HD6mVUQkIin7CECZvqy0nng1JsJIEuBj6r+rsOGm8fBzvNw8kL3hP0aWyV9elW9R
Tc1n+MB6vuhKsK3zKZFzPa+E5Jrc+T0Wyz2TuxvqlMnmjOqhjLsZHtBrr2xkpZIb
WaMHze8e2uRhOu/707hToF/ttqSHFUk85L59phQtV+qt0+d+C1HFt3+eQhYxoizb
5GTUqZrMs4HhrTnNTQJh5cp2fLOeGNh+HbqdVpAbHHpgVuWa03m/cbbMNWZiVWci
/fX8WwadwwoXbpdj0udh6GaL7Ci87GP21tI27Sj2H/zvut5keJSxFo/7pUn6SdTD
zxn16WgZmn3jw+vG5qsweoouMFlyJ3Sac0oQlWum6JR4N6jWBTDlRiDi6SRG6f5s
/ydXzZI62ECrewNLfP5zG+dXAt1XeYdrdZFsB1glN5fuEbSsycthVmmINJZgZY32
ySFa67KQdzUbmAXfUBsUUdv/oomVGahXCOBVjA/uiDWUbKrPnHguo6+JAZlIjl+p
iNXD1VD7AenkyglrS9qkCf0sSmx4teKiP82Ogj1GQXpw56SvHTBNWTxn6uWD6U+w
jGZkMjNQzwt7xiTBxjBJyGOElap3KTfMUD8LFzdcSGCmzx1joljhcizhj42Uf1dy
iilQVGXtDTThAaBzahCq2rKyhOJHCErZHA3O/ZCRn4/A178KYd8tgQaV9PS7tBFP
w4ACkviXBgu7PsTxB1yz6hFMmb0h3YSpPxpz+GXGiqAjRg6y6zbZdOq+oZAsQQEa
mV924kPeOGBSK6C0O1+DJ4UJPmk4l8zCvY5HYBxGZqABO6fMtcpK2cHQiu2I3W99
rCiPRlc547bXKbK6Inx9cnYs6RFDj2/olX1FCtREdp7u+LdKSwLHIMORFmhxunim
UYpTxtdneNzPXqOzC8xouPGpGrMZAIy4gD2Zwct41oYgbKLlYjpg9JlK/NjJUT6d
60eK46SYxTlBNJuRlBn8JlXyQU0IIQO94puClT2+0VvCwplyanAFHmrnwg2dv+Iw
PLaQ0jmnuNOt/Yhtb3CAqvhPTZy2FSG5sUcAaytHVx2N/qZH0T3xrNpbTOnwLpkl
VOwNkmr3BVOVC4GoLxXuc/PvGizBhvbTPWVglVOnH/qGuFAdjR36IRQ7KZ01hiKW
KTbAzo+lpX6HXxcC46V/vwjqyXHsfzMwwoOR4svc4YNW/XJslXZrDiKSu5U1SuVk
D+CJEXgODNxciNjoUs8XewK/hW/VJBNAKMFaW7SSKdt3G//ei06/WLzy3SlJQtdo
6g/lqCjyTeVpszHALc+wmVxkRwDtYqPobL480vtPleqBC2E48VqgOkriapIGwuvD
ZOqweIosv0FDeDQ9qlbwuEO5IaTHSy0S6NEzZQo/0Qd0JLF/73e+f/LqxhZeSR8A
jl1EUk8qIaDgNM3HATBnJrYmufgs7n1aa2Vbf87S3uIoiwcOXrva9Y+3ZJO3wP5W
2ZDCAZcsloqkvSUmAJenUbvzmXyuh/A+kDofXIM1P2BXY7kDpwX1Z08Wd/LhEPbD
IbM5UtyWok2Lf+q5ZPXk5fNAYBI0ugjmyCRokFec1FIrHPrvLXMC6Zyslx07N9v3
YxohBUqb7PLS2SLo0ZsuNotwCcyPJ76ooNdO1QgronZFRiOMwv5ylmUqgDZAKisR
rVfs2XGBe7KLNP1OtNaF/ri6xaKACNJsjG6MK6d1jQM3AMNSBsYkUd48ySq8RBSi
8ZsNn0SLhs0FUWN29Efe9Q+n4GLi5F1PiNtHVEfkH+zhL+XwTs0fgcHgkJSVurQK
yGJaNS+UpU1+4I7ST1enjiU/QCwZHS/FhkK8zb96VieNYqUXIT9NWWeQ4HsVNzJQ
ZdmtCKrRD2b5sPFtXPZHN+kWz2kQei0pp+jNG9UL+HOtYpcgvx4Oh9T/EDEQe7sv
GjR7q15GieeBMa+YFuHJJ78Yk2Vqwy9mA1HPOSrk8kwTDs++RxTWqfzjPtF2LT8H
GseV0DTTGndaR5G+o3SWmMm5V7cB2w+4KK8RJawUUz6Mc5orDX8SqrgPH+ZVeK1K
fnIPGiYn21grXMmkhvfraRjnkfYaEt3UqfsbuU/WQqb808aibOvvmiwO75beI+Wv
wwS4NgYUH8u2Sk02yiCrOnEopf30s7dl55jdbHh/k1vsTYn4NVCZmI3prT+N2idv
WbJcT4ziiX/vBKDfHZWCCCb5hQSFrRKD83m7vwxx03yPjno3ESLC08xKR626JGsf
+12LUqEYDiGa6yiA/oo5Gv86Ql3XSTtcsvp2Z8Zp1rx/Ly6HqndHrj8EdPlCBeYC
6DNuNcZ9xn9H9nuE2y3YjuBkqal4yU7aCGDxKs+VpMXnE9eg2WEZTxTy75kJrnTc
uGDm5FCFqKsCP0z2tQ7wRNsMRVl2YgjaSzXd7nGs5qDTqc12qs+8nY1A/Y2L505l
BxnaQAXHj48GHJXa9m7DaF3z19yc8zT+wa4l3GZu9EspjkBG7TRP6k9wpYo3Ae8B
fYrhIloXf9VT1w57E0RPrd7iPSgWLEAKjIvIKkFzYKbNSVz+rbEr+lpBNvAPXFT2
UQa21Kb3vnSTY8qQMqhBUqBZfwAEUALDo6LAba+dn5Fhtjh/U4qKpjwefxh0Jywe
M2cMdbFJAtSjKPttLN4bVV7/mYE+C7iTsOtTErO17SAObN862sD0yUG+15SiQHZU
YggEKMlxF1pwKVUh0rIPhW5jm42AZXPK0BbPxuCEtwpwggRTb00pGEtcbI3Axmla
Kw9bFWqgzgFFsfO1h8fsw0lrNcQJwaZh86Qf5MsZA/Q52SdjDFYBsmMyWufwxl2I
3fy2UvokfUr26fL4NpWENNm7D/3/cBjtkMsxy3/l/ggLr6POvvTNH3k6QVh4Zh62
1FFFVq3OQ6rka+KSAPp+OMawTNjE6j9zfbyEaVWtr60lRle23NF0TxX2IdGegflt
Y8G6IX1qSLdaavDFMkfvUQagElXAhwY2z8Bb78jn9imQWCOcwc/+6It+4+nGjr9N
Ld/hpjk2S44jV3+OJIbQPg1JINYW+QOEJz3FrL9WkSe/J3naWlEfD+0ZBo1bpKKi
sv6jRActqEkK0oca5PHhgu8/N3ZgtZ1argmfmGdHqX5XTVp0LLVdXMGLGpXZ4kGU
Cgi0AkMD0iEyJzTzilHHGa4otz3yThKr122MONSpOQvhpCNs4sHh6tpAZKsvKVCC
hMqpKVZixYALD95LAUgMq6tV5vE0cL9vDby+49GvIH274nEaPDD6OYpp0RH2Tn+C
s+4N2czVDaM1yZ+wwcfTpa9nJCp5LOf656xCMpQdFu0ghXfPvH/cbQPPP+QOLKH5
VszZZng3QDRniSrzoFnvRrKmfZC9XisbpyVRxoZNzEySsm/H8JsbsYHXvI9zm3AO
j+YMRQTC9M7iOQttg49FHlBEfpjEpLLn0dg45d0u6Q9hDy0vlNfguAGMQ3zeqfLk
z8PKJkv7AB9suUJuQ4gKtrKSeHgkj5Kix4uLC8TlAcUidOcVOPiHvC2sM2t5Y8qN
vpNaE+z0wL5qXESxoV2h5NTbaAHKPRyEOR1cCbVOacfen8HO7Xs5MMlVGKXGmso2
hXpMDNfQdmFjQT5htu+alf/NsbiHWq1tuIz//s4H1ivUldKOifdPPIgZg7FKoJgk
XaL1YgioqmN9pxv4zrptWlysQvHhMYyJaBz7ffRM3da3fF7znRXgtQj8KM/BykXN
BK9VLs8o/BJtJwp6nkQwFM2NRVU2OEvWI9zbBPAesXco6KJdZL2DJxfFylt4SDNu
gDNEcY5uxvgpmChDwGpuypzfTtdWd72qgmKsEvsZoCwgiXqhM/GMO5Dd5BiZ7PAr
94chL3aXn4JDPg14Zey8e/O9xi4uSd8XVtZhhPPY3PFY4vZSHGxNU4Zc3pqtEXja
VoxeX2wTB7/xwzYqTRVNQvKasb9elU1UXBctA0bUWqaeBiVFuNw8QHPyKEEJzCCm
QFMOUeJ/IRxqgbWLsuhXngEfdggaq7P9NxN87YlldbQYYBLA9CYtaRm91pYs7Nhs
8qjdk5AbQDMebXmx+sCdbMIHBZQGD26cK65GZsHn5Jpl31Q7xTr8P3f76mOhGEfk
Rc5KWSjVybfqQjWPAa2dYwMsRfeRZwqMCYXs/sVkCx8Enb4M4wfCThczCiSS2FgF
2WHVcrkE6AuxO2A/13nY4D4c1N89ZjGEIhU292qowT+0e674lKOifRAqIIxy1eQf
0+Tyzrl99ZxbDIBZ77wcexQpCoD5ZXgZG4cWghssWbrLMRbMK0hpSy4Xk6ZOs9xM
2jiCkOcC0SBcelDIX+1IvNBUZjFChSK4t0ecpcivFiJm7akHYHO5KnurBWWFXO3R
E4vX81wDY2SZmzYI5hl2GD4f5tyDnZl9ngKZctnQtE+WMIamshegBEX2MKgSgCo3
G2mr14SQOTBoRTIDPcIYxDgpBBciocAbAk4RwRM8uCQ5GZsC+KQB/BBLfcoN12zA
sp9vgKEkhUPKL+WdUTvdf1tY+B4CMZFEu3K8zSn0aClgXou+62BxQlY17uUmpIGu
VwUFWdCoSKqPZOqCy9GxCgfMSuqD2mcSZeoQshbwXnK8mW3rQPsr22YtsqDBBgoq
xDoDeJOaYwnDI+YiRSPs+D9TnQMoPtgGJfLfLYLbo98a8QjAEGSiSQ4eF/OGoUrD
EDG9a3JypFA9NeqS3WkP1aPMjkGBYEpeAnaBIHgXk1rJRmkVxR5oVCiJuXPEmpUo
MeiHYbTayVPNECnUr/03cHtyRCkLKtYKYFxPf8SCgqsR30WIvY331OWqqBr33P+n
nFd7WWS7BE0MFE0WaCavNvyR8Ld97SapJlwOqCUvon5aiCQBHsOhvKmFksPm82tb
C9nuhn7HaEdPEthp47xKmoV0D6EoWZcUefygvy2/4qaFRI5bnTLSoaUkIezpnfmR
FFDmmFSlmdYAV2N/k7JS/7KwAy/QLxDDoqsCvCQU+i7XK/CngdpT0GNdQ8c6o0dp
eaBU8YgV8ds6OpvjsMInqyoRgl8/nX+1LEQRMQ66VROZhK5uBbSPRSJwHsipJq0U
iYnwTpAmyJy5CLf/raWp5kVL6l7471lOuXhA4cPmDqZKi38crsPDDRnKs2jN+oHU
Usl9PC7fiwXKLuZyHWhZodHUypFIv5nABF8DyJ8KGUhdfEdzbeikpGiodbxAZPZy
2G68LQpRmmlCYobyKAJp8EDIAZY4RU0XBjZcDMSbkDaLF6pvc3EIi5QYUrDPZoj5
+k2auX9g2z1LdWOKSrDUHR+Sc0A/IyITxXGtrPHCf3jFUZUO2u/AbWkKRajMLFsV
XCiA2qrLMA21sV4qQWlmXay3rmLgrRb7H4cdNNcRK51NnC5aPhmdU+p2R6xjGeaI
LMv1Dq78xaGfe07LcVWdur2ZMVOP7uv/Izc15IhA9X9UOuAHfUgfksB/Q9WAd8Q1
3dP56vW980qgGQUhWaWqhS5+Ou12EMIaY8fTBuPt7ybWn03JYSW3nm+HqYj2gMG7
4v89kNewz+ayzibhOqUu+IqcVPEFWQy05mEF+ERkJCTV1yLD4zVZ8Kr5dkIhT/rN
HVcOqipZWJnZbDxuVz/QIcI0evxjR18ky4Yy1tujo5RC57pZEQCC/S0O6+cl5Dwn
t7td/s6OBqoXZazY0/9w77cgTg9qrkiJ3vlp3wzmpebDfKUeQdsVGW3lc3c39QTa
zVzlZYcoCby5Nf8xR0Jli/A279bDIY4rhmMbpKDXNC9ot7NZfJI/2UeOwMBusHoC
kICxfn1Tpc4WvdGVnKcBQ32rnbeSMYiXkhLB+hJ5kubNT1cJnXJ+UWETf1TQFFht
LYAM+OBOamNunx16kXcEeuLrpMCh/bNbEF5dscf9eOsbXhfmFCcL2iFk3OUF9A4Y
W8r3sxGoxzjuCL7qf4dMMzzScpkQ6pv0qtA9ukFgDF0xjCkHfnsUhdPmTLAchooP
2BRdFYeLgsbuf8wLk2IqnfifNItaaltY8QOxM+u3RMThVZc1tCRH668LWrIqMLw0
mZ3QMBtljAN5ZxozGUs8ALOZDoe4pEBPIOA5G3WDU1xcaKzbxoQBKUE8yNW1sFw9
NZykCH1MKs1zQDUhiq7ysmlwSGOeM/3fRPwRnyJkhj3b8bYrAn1S0gF9gFqypFGy
URs1AGYri2W4Zc/nEQhE8ZM4abt+xtRgz8Dwl4WB9pQ8mD3AejUGqcbGtKAweXUK
VmiRcVWzJTTHf7ig6QxMaQwc7nuzbDIufmRuwheu1SFBFqYaLqfywDRhNCh06qOv
yJoqJ51ZXMKPpY+aH8SfoAM1UT8qVxrhuMo4r/BoRvSTgBH2fFtiHUq7IAZeTHvN
AWMZeCZ2MNCFHSL8l5sZ5XvRP8+gr8moH1h0j0ZvBPuNbuQV87wINh/5NRLgnGcf
BK39qJqsop46pg6reg0b3XF1S9k1PwHxh7WZEX1sI+6L/qSHcXvJsBN1ROk5XLmx
wnKBqLejaopaDmRQF8Jqqcv7TScACfvMUWDSeHvKGhpN8Eo0wzzOo7HMPdjC+isF
MFLxIjGU3l7eFz7ebK8IFIp3fRsNfIXRqKyOhjY3gZdjHh3vNDxnWUGccyfEmQw3
tG2+wXgM3RTwAkjtFGTtLZJLwb4zOC+KVMNpSLddhURxNUe92xornJOB1s7mG1bZ
jozpPxVpo10NXAQ+S+g1Bc+FTVKW4/Kh+V6I2UnoGFqOJAIqIpNXZLD8Tv5pAx6K
BkJuDtuIfJgQcI0ecFf5/370OMxfbKZ3uhRM+VaXdN+Pi4BQsGeH90KbJYpsmru6
mozwqTqpYEohZ6CYJ1bpwr5dI40plsbH9VbDQZXNAGxxLqykV/B9yMTdhBXagfSu
ddBoTALOX/BS6N4bUB0AAB8oXbT/0TSui5RpAo8TIy+n+CcAIs1T1PDMipzVG6hY
keliGWxvPzGMU8nbLRpu0N714R/pPKUyKPf4ZrnK507S1um1kO3GKd4a5Djl5KJX
tZ2sGSk0N/Zl/jYIiYwUvSHw9IYehJz2xjWc031so/h3EFuYYK/sbJCGI7z+DdGz
pL9zHWEOZZ9s1it8/v4iGe2ag9OGwPSRwf55fWEhrVWoIxiIZyKG8LjSsvURMz6k
6lVcNfcIq6O0X0aHmF4z4wVr3pWbLX9x+JNWG2WXDa7xEg/ho4YGty2Dz6/nYY71
aycBz4WvjEsZ3A/M34RWprmzTd2fOuidBNU1jHvprJVmMO3VD5fDAdd1UEEu8v+k
Lsdvsi3riBqi4lfvVgihD5PYC9Kg7oQVLPrCww0u8Yo5LmGc0+FO3YsMbIpAGDJX
q1RLtmcNrUM4kDMGZqfCqMpnrnXmpUhcbXnqFTeL0aiTZhOdYcBrZ7STf9Re8ycr
2Yk+Ie25paD5JopWdIgdtComZF87s65MXN1eAMclEn/a2SkiJLmlG6LsaiH+hblJ
SGXAy6xb2seID1syN0CaiBnaOfIw0cOOj4wN5C6CRt9F22BQem1Lx9HJC9RIVgMh
PQOF9XEdRZU0rjbf7TWrlXBu4W1DpuSfJ2s5Vu6LiCb9jsTHOVp8QsNcBZCcikON
45acJTJKWTTQg/Vk1UrVUMoVOMjg/m1rc7oQwRyhIwi5N73qIxSgjLF2ATWM13XT
bhZj7KDWt+zmbZ2GNDyD03qoVJW7pBXf6VrBxSXp633NnB8IClZbYBoKKG2qrUPi
tonNXIDb+dB7M9gJVVV154M4XqOpRcWPBXLTMZbXGklhIzausGd514LeoQBKravM
N9+O6/Xb+4A5yZ/VvvoVMeYRvlHzZqMTultMbp15/3Pa6UgTAM2ShXMg3l2agSS9
SC4U54eBO/7caqpcEobfC2k1SZ8HoRTQgo/IO2yu3WcwqqvKoKr5UUcO4ltZ8y7x
mqbphOON3eeZduPO2R36HXCwoPii1YUpXuy973SMXdLxFuabdfGF1aqmclcevpJN
6cpw+lxb1e1X0zeuldR6Mi8KxL1DYKiklKr+ee6GYbErSV0dDHxu1/Myfeat5/iX
UmkbsK5qa3+jJ/c6wa+p5szmiXil1FuKvz7/1tlmr7nmPjhlpqKRGJ1MDoshdrGb
gXBbAgNEBpQm+HN4zjvnl8SyIIZZf647bQlZj95RQafyZvkm+9J6z+32F5Lv1SNn
rnWCAM6BHCJKeLyhzRviD2ZPreBQ3BrU9T1iwMo7rqpTcH/nYRlfnmcmMjpIEfP+
trEdO0k49jxPKIr4rUeh0sW0m+i/MterIGo+VV3NzmcmXFTs5DZunQO65b1x+dVT
9EOHqfpH4BRknDLsROONb7ivv+m9k+3/VlkgVO8ZcW/K8TGKG8/VAJCEj3BUgEHP
c+qqtu6Z0GHypMDwqQVrlbONsyFSAOUaP9q+nPPR44pYycd4OcareN3TnTPN5uTX
EEZzhyCSt+xRNiwQgsHhXclzfu+mLvvXcvqZXAZxwVvX5qiCu7foQoiykRx9Yxbv
xtawEi2oPtowMuyFjLK2zEJjnkOBGlwFs/h0BSxc5gAjK4By7pEg522rwUfpRHcc
w0xbXloyJQ5A4K81J3oe/UXy9J2pxfaP+AOK6yL1vMVrpGmoBMBkK/RnFSrnPyfF
NxjKe6xKStbciICs5d+K2rhwfr5nFm4cSDmCWNWdI68uNo/+TeQrSTHDk/o9gdwY
n+tsFhP26+Pcy8VqseFIQwJpPnEnJE9Q/XBiGqWK7ngYWY/H9pzM/IdEOvfAocVL
tBkaG1ZPWFi5vkNqyMHXNDxaAuKwSJ9+Po2cEESjCmfRbw1QvbRANZ0erRlKModt
/cutcRbpkCTDSRSqcqzzJEvJQTLm6UiNUcGsWm8kkF7rJSVOdzGmHQn77M+xxgU8
Pw1xuvRK/ByGyaXGIg0850TCUDbO++QrjneCTIQNoOB3lTLnfRm/XERsUVIxyp1h
OvyVauwcYGR0MgBLyA9ot+f7Nvyiu740Z3nWBCaURiQlFPCvkYTNd+NxkHg18Gwp
Ve9J7ootFGYJyyP+cXynZgBZah8KG/XFRjISpV7TADh+3XluJeotLiwfGyPaHIZx
LIklCFFv08ZQnDBHJB1cTBhpBoxohIgunnCP03lWabS9Btpr1gdhamrP8TYf3Pgp
+tdeN1AExasI/4aM63xOmV7axKhEd8qJ+NphDV9piljPEkhP+gcOwPwktrOiPWd/
Umu90Cb7INcf1rr82h/P1tUcOFFYuXLQ/A5XaJLZhuVvvb0TMLMJnPpA3iv/yGFX
S3yT7e9CoTkut3TqAmbg42XYiCWIB1+HKrrZnn6JJUdFonvyvvSOpxCYUmKTGIxX
5egtzxbfV3ic4prJThDyrJgmR3btsKlcrLXkEuCtI9uN6XPBuAG0D9Z7KZcM8FpX
hf2u6xuvoo3IT+ssXQOUmD7WvFUgHxuxL4HFCv3KWGhrjnOEydY5acxE4lkPX/9B
Ca9O4ELHYzpsKbn+2KwQFBug2FjRSVEve9QMOUfiiOeYvm9JfJshHKskUNfRKCWW
pSShHa/uP10nV6P/zeTt1PmhPH9plL/AUme2oZ5Bj1v2XFbo1pa0LeQRtLbpNHM2
omFzFSPEkCn0hnuyMrAX3Demig7SK538yyTzdbv/pkMmVH3AHmlpl7JQOQ+EubUg
2Ixp6vIMzA80ssIuLVtTsn0Z0PsnPVDQLNP/y0BPmpVFSFhgIVoagPizs2+6ZJ9r
yJKHjkO4S45B+S6MoOhzumYIM9ODXM7TpJ+3XbXda/ak99BPwgzi9ix5CSj+1j2Y
z/R/Irt7NoKtHaxonO27PJ+zZ2Jc2BTE75415P04eaG49sJRWjo0QWK0uve7y8Pe
ZX2rGWNsh+98+TB3eplD8K1hdLnWu4e3hbLIQfC6NPXEbGD3OCiqKfXLCAiHyyq0
txIa5ElYuwtYJDjPgYWwyny/o6L4uwAcQTR18aP8kAWhBPPDY9FHIKE0phJ31YJ1
Mr4/vzAtoHXeV7BRMJ7vco5ZUWJJJ6f+63FKBCP3kpqz6xgh6XMJEP4Y1TOEmPe2
5pf8ePcSE6WI7B25Ad/Y9gTBK2Yh9h7m04GsZiGV5CKnXZzu//wc6Qqjw+slIH/w
u4HmgzWK+rqlKDymObPU8d2g42Z0cxJJeTyNf4sKUTivcAvs8LqMfefCOCi9xeLc
Qr29tcjEChlpuHqi/kkcd4keJmr/4K2iKzdz4OxlfJgL2rNVhuhqBz4a050fUsXl
umQKOCM7LgucbOfhPp0Ic972uCbOTKS2jYro4tFz+2FsBiscJL2BZYtf/yGW8dBJ
WyRqDZTvwIYqDNTMV0Q4UyNrzDX/J0AeKZ828R30o7rqzK+CO4J/ZYw/BsO8uruY
FUMKgjhLCr86FFg63alKQc6qaYfpaP0HtKWJGgsmfYUp/KslN/MvY1KXOST5TtTh
d8WC5ZEuANZ047pRqw/ehdgZrhlfqIlu/7XEPv0gsQsy8/DO5mIL3hMNF6vc9DBV
PcnJTu4HWlX+pf2iIZQTnho7EleRY3JdEZrkikXkuDIjvnvuQ0Af3ggZl/vkhUWd
e+/gBWArdR6b+HRIB0FM7EAaEsrB+qBt52H84bfgCkvM0DRDuIbxfVuKpHwGI7p9
nMVZ4DjJJswcZUsgC7Vcb6OqTzyE/JeetVbMc/ZbCMa343e0WPJUrxuD08eX3zf2
8UwMnZOal17OwEONV3UbXyLT7S2LC8/ebHiC36NE+P0pN0nlkU/OJQFEubxCKQFU
VT5FMQ2AvfhU4GXvBoGTJ0Q6jHXf/ZxD5K+ONtLsdD/PsXHpX/fPdYUtyEImDG0n
1DdTyqQ29yet+CKwl4g3LonfUT9uJewBBBwr3WEr0T2zzzcbmJY8KeFv1B3F4kOK
YWoYr1HAoHpvltDGcwIXNmNDYZ1z3CWl1whobFDXoPJc/cgO0eaKIFqC0MVAtpCg
NHm4AxGyACIkig9UydNT3X8T3JrTwQsAgctHANcOVH1FO0cF6nmT0R8F2xN59oid
oit2Etk3a6yll60HEAF+Pt9jfxa9a/+37CLC5/n5jeH1W4mv24vcvC1Eu6VkngbU
JGqjO108LgIYRcsioM+DgLshMNUoPZJY47rQUpaYGnsb9eSn/qw5eYrnJjH3OIPE
9e5p61NgTIEz/ELNbDEfi/GeVhiWbyU1s5YSjGcpd0a89dV9zfJIh+n73724V+6d
ST5Nsc1U2TPka0ptf1k/uZvSKpikGeGdFcd7WPmPzqoNIzeKP4NePkSJlMMHjuYb
ROo5pbjd3a9hHwMmMYZNvsJM7r/YOliC1deYxThuZ6UQgGYOTK0npLGM18A6zSfc
3ERpa23XUDr5xbTXNLruwszHducyjTmxTA3zJxroMQxgx54awtCVxRO1RShGhUEk
/4PcQW/s2ZEvd9j0WjWKagJhbNhtegLej3boDHJps2+VuvoUuDeo3iAKBc2PI3HA
IOEqlwi7egWFb+PL0tRIPM8Lr7XevTNfxh3Zf6Cst7n67Yzycma2W3K4vpe91hpw
2yQYyhBgjmL0j8L7dvNoQIIvvoXVNvYoC92lf1tZ5Mws7duDRb/aNvPuwe/F0SoH
hBN8KbXEuqxI4ty903iT/rwV6HWZFG2XwfQkfK9bNqmiizLnOlbF5eND/AftJC86
rKXcqydRuliKII3lGe19MM0DTwIc5ieuxPreEE561oqMRAgrcC53Qmb0YRnms7nK
bmYZRCEKw6UPZCicT1x25cQ9VzXUieJFW2Bo1v4ac1MxEqUeAv4xG/UYBrPXAZsm
FTjdz1z+YZiSvKQxKhyOr7sF90vu699DxnEcznA5Ob7n6z6Xz26CMjOGZlRQnpF1
uJFLo+H5+CHDPp5yYozBjQb8QWOeYeWwoe4a4s6UMXqykR+eebBdpWyxU/QZLCda
mQ9aDT2+bVYRCsLnALUbiFD845CgcUMKcjHbiLE3umVLw8ocGLCdlFJT0cmL9wQi
agUAlkOVHDIdq+2BKwm34CHr2wHBxFPVLE7SDXvzSfcxRdfJaMRb65wJiwzkKCgS
DAURao4LGcUDSylS/q4cX1o6xXXlqPCDsgJVCHd0/qkJAqX5D8oNYOZdSTOvsRC1
3nAqWi/FCz5WNu/JthLb0XSqumEaPjmeN26rU9E8bTey/tibhE8lnoc8W/0oVHuR
pO9r8q3A8myJT7of6ZZpc1ncIRkF/0hIy+8Q+OaFzLXiR/WRrkjJWENO7aM9eicQ
/DNFBqFczCROlIG4ODH27M//R0tJ+fa/HDIDaaJGkSf2giGuhxCrHxq/7Ix6WJvm
oMlKu7PsowUF5RXFf2XPsfKA6v+RDChzLOWrB2XZ5WITQr9tWL4lw6+SP9W64Klc
EgBDyXUgOb4xLvBS3u4vmlA+4LBiZZ29Hnpd9g1SGEU7fRWqowTCjaiYOXUq2Krd
vx3RloTAp7yfLyawBSFmlZUpIqCD11Anxk1qqdPm3ZxQ737k8O34pCCA94/BNRr7
iMV69VQA/Ic0AKisRK1+zbGzz0APNINzN6a/zhOndXmapbjmVC78hzUcL1t8zGI5
DfHUu3EC6QZyDIqECBGHvUhdFLsmaQ30Lezsx7nOoDZeyXzeD6poh1ADrt+BvUAx
CC/TRQofrSlhPmb0/wQ5ZCHbE5UnUwfzfmDsdEzDldvJmdrdKn7sWhpbksVcDr87
WFr/bT5ws/JRV7hH5iyW28rU3+yfSelr1pT+JlTaaMXN6Csrsm6sj83zOsxynOd4
eNKnPp+EtHwUCS61r/MQGp8xwsUpDjoHpHPjjOUErK2Af1oBs9ucUCRiIIeZKPGc
FVwuArIVWOV7VpGxEInsUdDqGAVBKj8vChb9fk3e2/mRB2eWKDra2Yxwa9/ZGDdp
jkhKNcXH7dHY50DybKpR/mpieYd3fnoam8AsQTR7vrJQkMNijBYiQG+ZB7toHCge
CmNeZZpuNrg2vValrOaTHkGFhNyQ03iaHQ1abhM6jzg0IeUZkLNP2bRceyFtHQue
gNthY5ZfUOALay7R5BZ0BW5/XI9pUMfzzIQxh6mz3k6g3FSK5qtwzML1v/mItU6q
CuVNL6n4N8gwbQP5Md1mvSdMOQjIDb5ZuXXBJcrY+TYvwwIwjsyd+n88m4bbNOlM
Y9khaMpgh3MUMHb3yJPRbd1CbBzSz5UAxNj6GiWUtJ3mHOOtbde7KtvUrhufkzJt
ut6RbXEUhKg4E5jwK+1eaQtlQM2GnriKb9G1whxWssZIR/bIo3kbY8UUg7JzzgE0
Ih35RrFuBj1YrrOJ61E+PymEgsKl1Vu+9IT6SQoG6ppb7F3E23tpXmTMv+d78wQE
mTWxvOUmC9aH+Hilna7WoxCe2aNTc7ecBbTs0WuGI0wURrCpYD3MQH5MRwCeUmCA
xuVR1j8g4Lt+GW7K4j3UkUxwTDUejbZomJLEufW33S5JDPP2PhtJe1deyXgHiKqA
G6lswXsrw+nEl7no9nqqD0SNx5EK4qpjobwrg7qWK4wF0rNlWTK0Zo+tlUaWzvNf
O/QwwVEzolLO3WW+GwP7jpou5lundtUA6UadmQmSqb66tY+763cOaQc+ChDZKcuZ
hqLRH54mYrwLVmm0bs+EFnxgfX+fqM9EEUjSp3QrvJA2MC8fZQCBHvKvr3vcmnAN
2+TEnmgv4CuorQnj7l+YIHEqDjDyyZ8+sHmnnFYlfXfTiG3DA0dzPiZYbN4zkhNi
gqt3nBdlqtiw/YaMLHHhd+cKdXXk661WJ4AIxFoVPFy66QJX2UJqqy4Fu8q+wYyI
nbe5GEfK7YkxhmRpJj6sGFu7fvv8ZZbHyuiQ9T1FODYnxoUSY3v2/5Y92LB9RLLD
m7mFa+OWEABZhk9nxDYSmuXSgBxmZib3yhMvfBgHsCutZJtyPAKL4BS/H9CiqgAb
FpM3o48+yhobHJgGnY5iTP7ohOULrnFeSHXzZI1bMOHhNv0HbzI52BLVJLh818Ha
W59o1YrODBlPBDI2BKsSPzZxAuiHT3jPhQsyaRQDpGLav7uD1XUvpX1+BcFyD8HE
7T7ZLryywtx8GsYXOUSgKqyGTYPj771uze+L4sJzsyibtqOePvZGdbHJHtJscx28
Gj9MzIIWhs1W1iWftYPla/ocGOEkuTNU0/fWSv4Eo5c2FdUc+jSC6kS1zik794yO
oGMbCxq23j5Vnsryw4aqdlcRKnXu8Mn7Fp9v7wXK4b2EAyMKWyFwQ9H9JH3x+1QK
96nr9vDomZwpBaGBAN4FnPCif1Q4PAA/56yCzaa3AdNnRtb6wWo6UBPLazVTJZJi
d7N4mIvgSk36dlQnEyCfkzMfydhF8e8TYRhi4g4qVlyYwordMUZh/ForzdkFUkfe
2/XdtOsxtQtHScikBpxwXedxaoAnkRRL7MkIXWCPMN3n9J6VPVavjRjs2+vnKJru
mp3IE0wzLHdVQ9JeR6cGbZ53nszmF5nK6J2X2cFZHy7RITQO8RKX37uAYUOONvi5
8hlQBMxNUJwSJA1gxwC1YYLIQmx1yX7id4ELXxG4+e8Uz479UM5ieQmJ+BbRwLd+
kDmbxdp439LeLv+iFJ+Hxt8F1oAfysbYuwvi3mIMkTGcc+A3/vQTestjSBSEg7c+
+LyHmQ2b3blo5M/LL2/MwsIaFXuGyIfMCnPZMQNBW01yYoPVG/PNN09fB3A5n/o4
NNChy69JIEB+xRbTSwHPVPPqV1ZcaABs3myyDAs780sy85rOHxQeQUV6hD596IkX
XOri0bhz8MDhYGtGhMIrh6I1T+JSpYvhLevbF+NtdQMrJ9k573+4RyztKGl1Hyf5
RILiDJdqhDqikkFlDI05rB3cTd2Zdx/vaC/baFGkT/TDJe0XJRmzRC764deeAlM7
jhMe9OQT/mvWoiW7UTdW5vafkGD/FHGSdVBjiJvXCSVeSyR6BUZCZqZ97FBsYvYX
362VQT23JL+Bs3rYhG6+gDq3CkfIeytiUi+QVmC1ZrbkLETt0rxW4qgqHXWQgLqv
SAuCc1UBe0V4WbplSc56CHlb5986n5CXRonjBfUQ9XCwN3xOjDNiV3lpgSTYmuYM
P2b4BehpbQSMz6KV87TwZUT2FK8K8+nPOZPNQ+NOsY6a+61JOm1wnLBgnuXw1OSZ
zVrhxSkmaEPz/iYfqlpdyBJkw/nR3Fr/Jo+q9Bgd7ges0yv52wsZa10oyYUSp9Qs
En+/D3xwwiUxZtsrzG75xXcMM3FupzpPEHjunl6AxvJ+eLDRHuzSt+KWMT0VJ7BB
ssazgwN6pdEna6MZ8rq3l5Z5SE+420/xv3W9jc2T0mvj9UfFA3boYK4ArOVDBpGY
b6eGxwXNKGsz/yEWyNUFWVkKKtcQlyo/LK3iiLkPZSkKSYxnk3hsEdn0YfnzlVSS
COMaV8w8ffxLrlUTF86JsQ2OWZisYtqQCaU8k7oUhPAgtQ9AtqrMgI5mRmW3XWVW
uuPjUG3NI8pYahahOjjf+vuJoIUdUnsQ28q7DsOK3k3rDDUSSfZFQZalFU9mRSLl
3YgMWswWly6sZ01pnrDm5AOm1XZ0OdtWnfdmznvqqVD8A9FkRsbXgABf2FVlzuZs
fHgNzKfCzE8UamLYnWNc5HRkQ4sgRFkf2K+UHCH/JerQEA52gLCoC59Tk34hyU27
0xOdugCc4H3Bbrn8tHHvX1AaSXFIxFCfkDmEFSwpYU2jcfPCunZTVl2AbtRXoCEK
wG0ixF0wY9G9IGi8q7LjRGsCpyoQuhbtinZnZrJQ6AzyG7Avcmc5EOamT+rPdfxL
mcnU1Zkqpa9irPPLVz2FK+6Q66QdRRGBnigoal2n/PAKFKeOmkbbpFCuHHJTa3sO
QEqu6ZU44ci3My5D0nMhScdLL2aMAu391IAHMuN5e1G6Rs/ZlzOT9aSoBkVNa6lB
I/H8wshRMaWFdEcBrZYPUch2QbShMZt0wa16T8ctzpQ3KjfUuP5MXjYGbU9UTUXD
opShcF+vywf6Gwva3xe9NMTgKzjt0Aoq2Mg2pnCp92rg0pYsjgTc1BB0eQbh3+gl
LtwyJsh8Oz19WLM7TYml4XdJsV05VmJstWf9OMN/lmqap2KJxt0U5yt2kDJbEPxd
opj5zZWBCtXzFBtHMq9VHKHarZkOETrkSL8A3hKld9bd/ps6/C8pyVrck/jI+BEN
rJiyi3shsu898GzKySULnUyeJp4zvwaMC9VETBC2j6i6J6QyHTby588RVCIu9U2/
4peDcv/ErCYh0qtgk5cempY0pI9IgNP4toJauptEBmOLKtcWzxplXFr9eirwN5P8
MWF5NxY7C9GQPbQaErUVuWB2ua14kBc439qbWqMM+oHXIc76E9mbeTgCBvML/uqZ
jmNH6R7LILmMuG+F8M9svPn7x4EGNHRYi7Tl32P63DxQmuHxc1ecs+H/La67AP5R
O05dt7TAiYlsRZZGECMlKe4S2c7IXidCztT52L5CA7aK9GpK78wJRojII9LjjCkG
vt7in7temiwuL1I8iQ20h9TNLdYVJn05Dlu9iynJX85Gdvpa8CJqDcBZcX3+gogi
QdMF6gxtsT9EuYyYtgNY+sgOV0SjsW9moi/tt8+IwG1DMLx+zem9q0X3Ny8HYGW9
TWK4xfVfINxsbQhEvjKc9Dl6AP22aQ+hlc2Aj+4dPcJz7FF6B8A5YaGYmmaeOdQQ
I7yCJJzJzL2VfTi3otfoBYBwaz3QeGtU6spOTwcPcrw7bgshkIAGJINGm+Dq+yes
ccywX44CxT+qE754L7h6lMCcJIcIkEkG+5gqniSTsyZAolhtKpPP9RTMwwUGQr6h
W2RkkWLBY7iFuJ49N073QkhoheXgBe5xT4drV8kS4ukmSLv1xIzksqoD77/+4zb4
o5yB+jWNVvcbYNyDjZ1iNTx3YSXK1o20IBeF1yaVJDGJ+Frrv6gcR/n76QJN5GmM
odcB8HFTfZEpWlD508QgsM2j/Yip4qxFSTpJekAf0GdoQJevRoPsRS/0j0/PRNj4
olAhQ6YBmMCqIuLu2zoY5sjCIVxI+bcGDklXDr5Ntxepr0L5fWE2uYpsSVqv1YEg
qP6yKy1xP9f9SySGbQCMpYhGoFToGn6P6XeKsy8Sc4KQiQTcO9pZeuocpTf0su1o
WRVCHwP5Pv4QT+K77Qlj9ohBx5Xpowc03RmpM+QYC3edYCOmnnY5BBu8NdmBF8Fn
NqXf+5ct6jJ0D1mOoORCnUrt2NIrYA7ddUJYK68Ugrw1fq2aextmWezDorZCzcqH
SpSdHOMsQyCh86mKMZGderYjaNE9hqLXhoJpcylArJ1769kzs4DWNTGmlY8OnBXF
wS31vovyDC+HGt5V0281AhnkxtGTf37W+iMjNpo3ulbICGM5UwZW5ig7IQNAqrFP
cBqKFr8uGWDgv/qfv9veFWhO5/fpR1ipHyDEEydZTh/rdVxCn1GdOmfqckhrqg9i
mUn3rClEjHtLS36AqW28jAiGqv3SNe+/pTMaOkRzPkZrdClvOL9tKZxxELSb4TVT
pnBSIDyt77C50RlESliUnPmyVMczusTRFPuT81l86vkBjkyzXFFX+qYvhRrXRUFj
4XQ+M1QdZl+xMOCuvRCnzfgeKidMCGsFhr0X5CKsY93NQEKDy0ErgL8853EotT2g
CXxF0knyv67JCAuJUIxjr0qrH70A+Pg1sllxjE+cnutpVtGWBJPQxDkIJpNAuDOR
J7LjNZ7cV4UDElzH/REoJV0mN1EjitXH749v6R/EhBvINQy8/o3zVjrYP9Q5O1+8
FAeZT+XZXuy6U6afTQN4JpdSKcS8/qBfIw67TitsH9q3+CQAFEP6ddO8GQaerJyz
vCBORyMLLA4uEHAceFxVaSvuL1llAlCqlwJjbalpv5CxlykfB74DJw4U4b3gBdsc
vxzpR1NvoKGSnbqvwPX5Pu1nm5pXR8jESyGdgPHQnWF/E0C6Pv0durqXC9KKRCOI
Y7TJ5s7OjDmFHt3OjzJsnFy9sjtuq8XmCrlZ1I0JEP9Ouja4ThptTyod2DuV39RD
+XDF9Hj5BN3WnpDxc+r705hPsIsgW8/ETWb/EKhgblCGHxg7wXMPZuM1fs5KBNjd
eKsjoLI8iKREjM1TX8wMqTAMHYOQfiyDEI6pfFAATCO5MaWu/3bvfEiPI4/a5fGJ
9bEmTfqHJeLPHGmmlmap/yMEV8Z3LSdwwK5fpqM2uLN+Lmexa6qqxup2o5Md9nC6
w8oQaLXFHSGs/ZKMwdJe9tT5m+yN+vNj8iP0XP28D2bzkvjT361Ma34KMYqTiwR1
S0YVwUnNxhoreCk5n5CSxkU405GUlm7Ol0pVn9odXMXfUkcwVsoykyDTO0Y3dYwo
GIEDarnTARO1slPfoBIsYUtAGZPPF0oUMKzerlfVfd/eJSa6gLL7NBXWZeY2HVyc
roCJPNQVt3MEFf/UOQvZlJX3Znpl4lvC2P3r9Sdx8esvdFdgResyECyziBr1oWi6
1cv6f9dWecsQs05vdlOMtjdwXsmgls8klxlvnTz4aJokYfB25TblOeLT+gBhPMLh
Wj8lPAhR1o+Dcyhoo2Ox6J3LxikbJMKssrR5ljNCJTUB/g2/QcnjQJsgdUTkK9lx
yQjFwWt2n1zNmG8DYHePjzBYr/DwgpIGfMx+B6saW58MTLIyk3mcqYtRFlB9IrVn
I/VJ0eXLKjtpbWsR6Mv8i1TOR7RdkSUEzeTPD+KbXi63heIXxmQbhkemTv1yMJZ8
TSgNt9XV1MdvpApEqh0PjuXQmFhNmeGD8a94MLWG+U++ZTCsDlprcNDoGh8f3evr
IpWQSEcHZdkYZ7ItJeZbn+ZjyvR1lch9kJTIVXFn8dfQi68NLtY45ijhcb+vR++U
8ddncXx1prQrEEFIW1IwkPv53YlEhcDP2k/b99FS5XsHXp3/wqR6Ii3Moc7LMDrA
E4sis90RhSG50VJ12E6C1jxxy29aLUDH2up/DeqCYLTlkLllfTW/ODaJQ+NLRgJt
wJcEr2truJFeGUYlq4HqAZH7XjjgK2cF6M9n3g79ghIBdAK0YRRALIXR0VpfT4fo
TucMr04gJMXjmiSCIj/+p/AzQ2BegwFnp5XfQNR+656DRI3fMI4k4nwPx2MEdsFO
dqP0fToa/Q+NHAzh7ol325ngQyi61cnHudqXq8JGGC3esr7z3UfRUoz/UShsV1MA
YTRM3OKQlTUXL2yR5XvsWP/5DYGBwM8jJvDtZjw/C8r7tDB5m38ONm2U8qWmheRw
n+gzpYQY/czpa0aamv6nZvKGHmFTZRdIRSub5w0CseUD6E1EVY2MRco1Cq4QFH0T
fxm8SQRYegy2nSHoWwtEruMsScgHW+9BFfQkXyga035PCHPnpLPhc1cZpAQ4Gp5H
+1vNgGXK0hSHx1TdSxf7NrZRQHotjis4gY7iPZm5ZGm+4Vv+4H0Vu6CxpckTr1ex
oiRsbYJYlQjt5JR0tQiUFMS7Lx7Whx8kzwWKQQgDlqFBH8o5enejVV3zayKkoLY3
fqz+vmV+5oDu03K/1Oy4ouomEIk4eBUomPtmaDl28/AmCctaWQ3It2CbkT2TwcP5
Dod6U/wMFnTBATF1jBTtpFWL9/EJQ0UkcOSVz/EHJ6W5n+PpLuoeXsKB7v4S7m2a
9SXHlbwtmxJ+GDxKRm6v6sGsBqs+h1mzjTa3sAjvL74bfKdPBnIK8/foUDVbgq9B
SQRxZpXE7YBzbOahCdyS1KEhcFDtH4qcMIyrLHCsIRHRwpu7bQdsrh2Dd4YGlLBz
vdkFClW4nTjTS5wbEY23RbRcwSgrmUrl4Pc1FECMNFDhygIX6uP8qQUqfXglP9if
Oa3TLcGzqOAQHDXSMuTbdI+9ScgNhhq584pmw+Czy/Mark+VFhm7UY4mn7Ox85nV
Zeutwt0s3vJ5I93A9TZyQnD2TcEBHUIBeT8N6ZpvqUJhIGAAq3qin/N3Unjr4dU+
GP+tdv6TPOa+oOQ5jMdPEgn+P1pFA0epNRHPO2IiBGtQxGyk1KnQSatEKGlJeQ43
34sh1ua4N5LJ0xiaxvJM+pLOWSkAhK/8isVl+r5g6Bcewwpn3RQpezqbT8isxgc3
n2e1O1SbT/mGQyc/7VExUUC7HOwUoqepC0HwLyZTgnX5ySHoAVrjOdUOO4YFj9RA
Mao4c4z9P1DktL6U2SwSq0kkOaG066YVsWi2W8L/8tcCHTwn418nUOUhLVaMLYaS
olF55k3bcljk7kA/w9AuEB6egzKYBkhUErVn3EfDhKaSqdhVlXRJznMWK0hREzAq
URlx8Nyr9T1Rm2WK4cRdsVl06cHoGNFvcyjGvn2XOCUjAaVgQVIJ8HOG8HYjU+fn
NH1/6HUZCn4IK/kZc4h+C4tPNqkPlIOGX4XeDkjzC9c9JF3Jhtvl0AZ9A7JzNNh5
DAjRhAaADi5ys2CAY2ONLaniIhM4SmbEDKI4hh2UOQCt4u0kcn7gtfbdiPJlLs+c
imbvi7kkyHb5bEO7jsPEjDPyxFL75wAH+ryvBiyx4x5Jovl/2m/gjHEgatWFVplz
Q16lQFNqWgqhK+I2exo2We4a0T3hCr9Xp2iZcBz3m331Vwu3SAz0JrKYH+bh+8i/
dNmXzixuBsAVWCtmDH5OsQl+t62f5g+zolDD0rPyIReWOSdZQXHqnJsPXXw4wmMf
+aX914rK39s/fTNxhWraQcsVaLgAvkTa5Ril3JaNulCqxLMwzpfXnnfFu0MP0zvb
NyaOnt8zKtZeLYHeAUvYqrWJHLr2MBlbSl9YziFtkxj4BJpJmD9QHoti4jsfwuEw
J4Q3H8YA8mpkAj1CU5/TmjwJXSRspyOxg/hIBLVqLrt0mJns1pPyG+Y5rXK6J5cR
FawhqOSyhbOtPf+0k4ydpapJTBFvAJpfPMioirpz9nuI6uUSl4uGEa2U2ipbp8Ju
E4bzWKQGwIumvGozyL2w34QfCDqiNVlRCJ3qrSxQ9z3PlrKD+5M7YKRY4GYfEy6i
I5snbgdBTznxFAuasJA0Q9CKvzMKgC8h9MLN/0Oix/GmlTTaAV+kMoK6DWa7YAZh
xUKw/eRtUWsRrTisKQJoNz+LzY5ZfpP0ilpV1IesBjCy5qTPUKLJijRJrZ2+X8pq
52kkgvbT+sicdh9sPLMv5OZ9FVccdpF8sJAJJBEjig8NdqPccqt/JWh9ra8iq7CU
9NUEQESl1YAbvytjIqtORpabtmww8cAo3JpsHGaHrjnuQzO5wh773qFHRA2KyQz2
nn1u5xUYzHBk2CVte8lNPbzIfdTUd0UE5iUNZWkgjlYRsuYQRHSi0qUObnPwRZfw
CDLrlXsyTC3ML4llsCVXUl3x8xqtH23OVv3dwhBOdL3b00RCAZ0StjoRhOrwrY0C
yb0jm33ipx3Qm1PQ/0zIUB+FkQWo/uviiP4kdWMLEa64DA+QYjP7uaFVwELRlimg
S83vdfx21PY6XXjWo3ZropFbyWwRpEZKCuzA+fFJ0d3quR5v15RYFdX4zbrzofJ2
bnimvI8U9+5hW2Uv3dngT/v7J725v46Lf6mlsy2P5Di6t4LAJt+UmmFg9I9ZrFL5
mpNgrBvMYW0GKdB8x5NUAnttvk8b2Zplpjczz/wx3Rua9RytSLuf3WzE3qHB33l2
GRWOWCPulnFmXNiW6QoaAPMjoJ6CmVeZ8bKtd6bYBEvuspv3rn/6N88oqxJPWs4k
lVi+ifL1/qR30O4Hr+k5+nnVj9PQtSE2RotTiOuRf5+Ar5gt7/4MGaK2GHfbnuI0
/aY7/rktQ1MQ3eIHxlNzASCpIrD04qOzrFoBCTJbFlCnVerbkqMNyumAkiQ742er
/tRFlzcPPUueYVzrkSwPgPSWLzyHaNSiWZKDDppMylaYW0wQsy1yaUKXdFoYojgd
e4xq17PO091hQlYlTIZAvtKOjM7riq5b/bi9rJC+XEQxpVTfFwtYseptgKekeFPd
mF3kwQ3UVf4QG3vxOLGzOw0vp0kY5tRaX/QSQmrtym/Bsdp/x1//mRu1O3G12Q8l
24Z5ozkjCHW96wafTn/BxTF4fGKwnltUC/SNTORzzQnLsWvh4SkorKIGC/f6RVJi
39UJW+udl9PE0TSmp+/Sp6+nFsk8ufiQvh44o1f3Dt/F+NtY5OB52/LBTWL1AuAU
/SogEXWz1Yu/DrsEEqOIRsEXhG4K71lMm6lO9kEeHFQSKsmZ5TpPFMySzvpECG2C
qg03cWTVd4JHwbddgk03Ai0owVSyNYxSfxW2uWohEkL+kYQnjmNdMEVmepIAcHfj
V9TVsFM/0UQL7SowMyXn01jSbmPkZyhAQNIbXw1vy6hUenwy8LltyTTmc+i6tkpO
Rmphf78HXhpmMOlWBWrPiuTr/Yns/hmzfCfKY4nNuIKe2UVPZsFk/OGrBQRNW4Vo
H48dsyt23fO4di/+e7JubMo+G/hDVPZzXFz85Rhqx8rQBknkPg9Q/b/7wdDnM1S+
PYByCWkFTdoabKKvpCeS9It/UpwjAuTApmp9hzel+pl0maZUKI0Xdo8xXmiwx2i8
GIwENLekUzG6JWvrD8UnxEfwHnxCNJOlvGilFSMqOBmsHWyLj5D7TWKS6mul61ON
/SL+SEJogCsFGuFqKDO/6g7gtmz2BfetI+IrR3SQQXGm7EJCwfGaUpn7alwZupqR
XMWM5DQxTb/qizqBrc03uD7l3B2qD5YZnuI5+i5ejXHO/kQo2e4aFrArDVIDEKnB
3TkjQwER1R9yNPz+8L+ImYqRua+OLCbF022Tvp9/tEqbLGraBkaw6AihBwUaHXVL
zxTQc+ZlRa3OixZEAIXbp8i8jxdfhJxUaqXtj2ZaTxhPGbvrv5vcUSBztYpKH3h3
4KvP8ryCplH0VNh6HWEbI8Zs6v5tEBjzR8HGEkZicNLfyQqgItAHJpb8K9R+Fub7
iWOtNy7XbCeD/F9oYsZsODnzsCG/dCw26l3On46jhdrz2zWuO6ObSl3SlacqOAuU
juOoc686ihCIym4qazyQryV8dIwXjaLPQD3t8abeDkU6977FL9IZAJyVw9GW4qgt
a4sg9c6+D/mI03a0POyD3UADsJEpS2+i1pE2QEHTkGXpepY01wNP2F6mIxa95LAO
k/iySYIyP2GEjwYULrwlNLgNK4S+47a7iSd+0Sg0CTRUw6yvC+/O2+Hg/M2mQCkL
gJV+uF53hcF6IszcYhfPnM+urzFmTqqnhpOh57PYmeqWIzIvrFQM1DgSkq7ucjOV
nqgzoeN67DtsMhHEfIS2ayazMNwxhoOKl9aoTQhlCcL5CGDILcQF2r8WeZyaeezW
oObZv0JRIuo0pB8pqJfC+S5dNXI8GBUzsbjqmJ+K+EsWgQhVrze/MRhqRY8nuseQ
gvbHO5+Iy8cO9k7hdo2Fq5ioc42szWhtRcB7kp5BAPyz6l6D+zMOZnDB8ydsHIq+
tCcx5EmWdNO6nQpM3Ui29DgEx6OAaM6tIQpzYARDflI94SfYKATkfiC9IedJyvga
ougDEgbIehU2fNn0IUkyDaVV50sou7PrwhtMF+8c99lPPRWlJnUH81rGh0I6RyKM
b9V28DxZnV13k+Z6JTHBW4pGhdDwczby3JPuiWlZeGU33h9BxtNUOq24N2M0bubM
VCAmhJPT0ZpVZvboCz6W2LapNO3rKQKNkrWMrWuzeXp9TMLPbDSBrQzgMsMBR5mf
sHInJ2EWzC4A9maGlEMGZSeGOFoc4Avj/LroRYcM703Y6qz7F5bHohK+Fm7uj13G
nN2AsT3S38a4LVph+qDDuHhK8mBbeepfmQn7g3ooQ49BChQsuUnwNz00c2Th0tPC
XRQ9ql+BdlrCFGScZaEg8DrXuDVici74tKsJowjiqV7be1SriCwiS5xfWjJl3TGe
0jLbbB9DedA+cpAUrrWkh4ND/EbHxHb7CQnfzYy40c4e3vojRQMOfbwKvSxyRjKZ
feCeogcWjyod4WcJsXZrIhkdKQ+JGlEe1fytlvumKIU4sM3akbbRj5KkrZvFpaDf
dgI0HPXQpAWKLyFTDAghTezyClL7Vjul3k7HLf6tbeEcwA8Jz7CvRkTNiQVPRXa8
3Ud20mTn/RB7lnwVd+NsB2+TkEmc2fAMISJNzQX/DAfHDRSu176Fe/oNkZ0KttJ3
Nigo5QBFj+OWjWgn3u/4ueQ8bPRhh84oWYEPoBLe/3awgsrqf5zV8pEVbfzS1MT/
pkQgYc6P3aD/4+ZsBRvacEH2dLsM0Wsr4Q91+dQJVRcVjfAG2NGMJ3x+OmNIHNb3
ywSp8uYQLOQChNVbi/MTftqt695PuKmW9/9aUXNvbOyBM+967zuA7jRRUhSgq1o/
C6SpWY5cYPQ/GAOcCAJfkjThkLh/YFF5PEUexT8ezCfoMD62EhAFYwVapParmorT
4apcT9yGEDcvZ8Vf1tYMlomDQ+s66rjIfNHKRT/FHbagVxGlsrywxfgvhkJdOHNW
cIvDAhwTaBSbi6q4aybPS3awYHN5KJ319EUre43STcMx67ShT8leMXntG1J3mK9O
4TY3SEOBptULxbNlwXbqp/exVscNyQN2qXxyhRTfQo0+zKIy4CXsPH87aZHDdGdc
kfqcFwtDnhPwTeDps88NJnT2rdSdJypwoMdyF0TY6KtJPxBLtYV2sEMnJg98141O
5+TBrUm/IWcBmXp4fUc8PGC8CAnVAykGRe7wOrr0RDoUYigDcn6ie52iWalLiZNF
DFHUvvC0XGeUqJarrsYeI9HIogbcwq14NZgWXAoE76zTeN11RAHXUQKMiTPdYiSn
NVvIO76jhRnn2NSxE/fDoEjIzqvitZAsOoQWj2ik5fC28E+gtPrL98EpAz1TlXEQ
UOhu5IWT2X50QLI9wHqF+pPxYWqOYYY2xyUV02PlZAqE4RrBXLC0YfMvuQdtrjVh
ay2bTBCdzI3Dtwj45nVQZg9wo5N7mvAsIGsykE4hwa/FGbv/Vl7RAJqppsfv10ZQ
aaATKdyUvQhuLFGyGzNI5gk0Mq5IP4KWYCtqoMTKMvJLhXWabe0/jWp8wicXAKwa
HMiQNUoLmqHfLyi+UKDLgfg3u0uTjqhajEulaOsRCtC/o1At5J8ym+MWBtkZhpOV
DXHm487++YS4He8/ZJD+6riEzPJ7oxUy8d3V9LdKNLxC9dAFGvpgJBSOWw/13vRI
ILpYr5ltE8KAMKm6LhhP6hkp7FB68Yip41TDhOXOXQZBvmNAPS/Swz6aZAAd96hf
BFV1Vfc88p9n36B5AAZnxPF00mvoREz5xgapRmWsh1CwgGUwp7CHRCtKaZJ4ORxy
/NYl03bAg4HSlo10LgJWOe04j9uDiJeDWyBPSZdEly46xqtjX9sBg63bVWBKjY6T
Pu/cGVFcfDbOCrlSlmOunHLtEdsKvxDjBuIDV66fKUFgVhi2UvH4k6EKAYPJOlPz
3PRFiq0Z49pQOoold3vwaBD11T3o0jo/txYNJh8a/DnK5aotsbfYJz3YoMXZAcmZ
GSVftPFeB53M/DUXYBncKbONEAlByKRcgYNaWLrHfO9SOhSey1zH/RB523zQCBkP
gnDlLr3PT8dn5D95wkNSbxAVGI+PZa97WEk7hotmUPf3yc79X+eWvHfE3D9NxOHG
U5WW2H1igYHhswVBv0+UYJjdEB7dppcSHXn8Uxug46ga6ZUsGRMxNP6ZoZMRqeCT
grh58WiJgjbiiV5pfgg6GDlCgTJUAfmFM53hSh+E3HaD+Jww/+3RRn9ZeX/3D2V/
sOuW0W3ui9Gu6W+L25BtNGblYPUmO3OWftYZ1HN86dX45QPSzD8aX9GYmwpPzly8
HfYDFODN0IbewGA3PCnXqmqVnBSgYBxravuUhLwEFdyTpfsVGUpAWKLj9Qqkkk6l
/Miz7aJYTExri8omlWRD7GIZoLYjz8sYQRjzMVcSDiFoSZ3eg+LlxyQD6Uc3JBoN
ZC91eG1aTPJXEQm/Jim2POoazqz4kG8zMJNFVc1r9/imbtWKxz4d7oFUtpO/o5n2
e1QPbE/pTRg44plX+Wmew35Zj1thxGBljB8B8bgLknbBZ57rZj8wWEDRoMxsGC5h
0TZAS5poNIih4+ge3YtxlEt5MZo6iuGpgMChgaSGow07iLf+YhlJHHMSl1myQvku
mM6rrKGBvESi4awmBbDFMucUOQEWwLuMdKJGoKjyBwKoGT1Oth7OILXAt76Kz7OQ
/DQ+0W44NckQ4gKAEQGFDMi+sCsI0WiNqXQ+1uCGYNFPiIkqKhIatghyojkMH2Ls
44F9Pr6XIVi7+0oJCtzo0TMJORsgiNfZD9Rjjtlew3Zp5wpRMd3gq6alIpjGTa/6
raD3RvowTCU8KOhSjyKnLA/L8IaQUaIEfZpt+VVarbN2rb7tjGLUWUwNeU3W2vZn
TTJDtU762SKw+XH/1PFVVtGbF6d/NWDsfR2va+otdd0uvg0n5EPxthdq+9S42J3m
oTpkToa+/g1h7GIGP6pOapb19XRok2yEYalk/Qe+MhCbwkNrCNQLO/kopjOuySJg
SXkcobxj8qnKxBXTZwkDIQfWHJJNKDHBH6axIYlcm+ulaYK2nslPRdVD2YOaEt3j
QutnpvgxGG5IHWN2byEqjV17JEeFgIr0eWPqZ2LDDiQWROfqYuhLOToLxirvH0IP
Y1t+50dWuRv/pMGl6IWdMmwgSxO4kAaYyKChqQd78x3aKTb16BHLXJvezj914Ubs
dNYiZeyZuOzGSf52JLwPoze8pt+ejKUHFrgKK0TzUY1GgoUrnWpPalWAMMhhD5Wc
qYa7FHwGLS9P83Glj0NR6g1kD4c9/joS1uBVcUwDGxrA3oa8LlnvT2GuOwlYDcbr
NfnmHkDEUewspId3UuQloPv31wuy9VIFdCwpIeh0zf3j0ZnPBvuooEgRl4b806sy
c78weY2AnlFaZR9nuX5L/1cZJ2/PekG1jSSPt5ASe5DMeT3p7v/fSiiG1TJFI7FE
vLCHrNTQSVakb080rH71AZEE3V1AjIsULgDkxIbqsChBBZHJxdac6LvTjM16ZQec
MddnSlhIS62Ki4YC57Devj9oZDEs0yoRKyzf+kURcJIfIgHGSL6RRAkWp4gr7eHr
ZFRDPfXc3n5qa50e1HUFZChXUjatv9emdQcfVW9bwJkyLCY0awXc7ZVEBe4EHLkk
r6FLvT2BZxZCUFl+g0dRq8sKjB5oroSqeSCValiOZasUE5NED6CKGulozEz6VDD3
tQ0CcDjDkfrvbwExZ4iB0ha0GxRmXlVm7gAtoMFZ2voet4qJqjkfhb7L//xPo3x/
Q/suOngpmtWJRSPamqCLCzf4GW81BFxWJKl4Oa12etyaGQpHlEcsOOxZz6IOTaAJ
fQ8La4+XDC+4r+yEFN7WDOPSB1khPkUUfAwvuyE+ntNl0d0Sk9mWDTAAwHng1xQE
jeJJ9ukofOfG2vQv0Zya1rxoOPUEGLEV+3mkuUAN1ntLC/M0xihj/ieRiKbzX3D6
pC7IcPOE2J8ZKuI1tfw6AM9FtD7V5JnaoW95WZb3EwRscX2jJIOGY/CFRICS7BOj
tmN07xHtLbr33m4j/TWqfQyBKsszNDwoLuK2nvoE69jPKsNvjjPHm7L5T1YIuVhG
OcL2kK/x2fD7oKRTCrbER5GlA7TvCYPkB2+nkOUk9DWv1rGzGe+EsyuAkwbTXUBN
G8DvnTGOAHCe0ZWtRymGpU2ZHVgY9E9ntZlJx4YAWt8wstfr8PtAgBMS1iSox4yC
sfxpV2L2saVN9oeRsufjb0XbY1P6f8RqXHWgGgwDzoZRBsc/LQgbQxMC9WGYafCr
AUpsftXmVnTBRzP++nNP/WMV/1KaXGao58Eg5YWnjE/DU2rXqkUm0BP5HgWqDX/Z
FrmwhaxCQ3aI3BzzoS3J9m345cHQYeQV7rHt+bL3E8wVvg9QmeZwXnDuIYrRDIg+
7jTGEfV0wzFQw33QDk1dFk4HBdpV7Tbm2UUZhm21n9NZDL5r1Lq3kk+PCbQWQqF5
i0N6nnY0C8ya7PINlSPbCKJIb6xcq587YLOEIP4UlIETs+fx6Y3mYIVB+HvruNoo
99JCmnV8BTPcMXxpyRTZmyFuF1xXa5nSQf3LK0o5ZznORtLg82v/8BPXoi4tUj5I
8jFJ+eA8RndTaNIQkFBk/4U8NtKTH4/fN/4pYCdF/yRs4xROyEoTDVrYnR+rxYph
GgKK5+BOg2fgJBA6YE2gOpQNhdATM8EUhF0QQ8r0talnvn+3bv65Bvrg124MWlQW
VP5312yVbnkbcHWQi7LmxKg1aB/LPQ3OIdpeg1YnM3BE86MeXaLXSRTKGKymxUXx
Yrg9Tg3XycIFoClLBIA90ywrPvgcxntuvPdoqZSTi6hQII5aYk7LDMq67TGxpMYY
g6o3WM2w3vbN/Q33TDOE7sgiMx6M2B8siNmV2Rb03y+0o3+y5ctzCg3CaV7DWxV/
pegoyY4Fm1quD+Tm6NCWNxparTiknPrEbZqmZLP3kCPojPKC+CpdjUEp720OHBoo
y6yBNK4I5dC1mRH9bHP8tRR6Ks9WJ7TTO6C6AIbZ8pb+/MCtV3+k/OaPsmNFwvAo
PMsWLNLiiQLcSmQKuoALCf9qSVJl6GLkM61eo6RqHnFZpB+0HfW0mIgRclGBQDae
TizeLIrtyprYBSLqQec8GaTbbm6tFZalVwBJs+CTRdABtLUWJuBKw4TE+6lWpAF3
27V190vo416F63tsa7MX/GJNMRGnJbnU8xZUAz4aX7MyJrrcBV4J79oug9d/C3m0
7iuKAM3+jHHkHSADpfeWgFybgkEhzo20sOsCCVeOSrQ5Afac7UxHnlgskH33+l4+
QWACD4vB3dhuo+GCUT0n2CD1WyEt2Oa00fAJggVojTWLHIYZMWf7FrS8MbgzcCU5
WBrGWRffxFGj2s8jYvohNfQm4ZXE8LH4qaacbtASqXuxto4IT07/42u+AgMJHM+C
/VdUQSZwKFoMr47PV6oV7wrAGSMfLEjFONMTu5TWtqHx2zLmNLy01LAr0xbyK7U5
2EP1eErwAdRegZv5JTjNN2+rlvPXf5f7YuJx0Km922oZRe9YMs+cKHBJ6WbDYahB
s6BdnO5grwfqhS1sDEleqr6fDQIzb7Et1exY/6sT2rZ+uiN18qqrqcXwKX6k2ztO
Y6Wz1y+Af8OPESuUvV01caXJzMMyz/UI5+jU6W4qg766TRLaZCLj2atfntpxswMf
RZ35LQGgl3mSzxbqP6P8uJ8+8v5RpxKQwO5PCZa3B8l6wWOuB96tK681iq2Dx1z4
LN4CM+vNsTaxGdRrqOPUiKziMg8uNCqdVWTLa3kHKOiAKNSSFRxMxHnM/Wmm/dae
AubigWNPi227ZSQ/E15CB9HI6qsLU2Xoi0LG90znbL5Q8WJ8h/K5PcDlELVz5B6b
dxBrK3U64ft6aRcGIhV2htP4QvafNrleCOJqbx/u7myuFqLBPbO8t6SCUvNfpg82
QQZUANfxWFE147s1qo0tMsJs4iIgijHE4x3oRPjewdb2N1vrMGZEBjOzHhafnRtG
mLA3nPV/IkzyYdkn5+wp43lu0JWbkvgd4Rqv/QySDmIe2y8lLU86eK6bV02DuqNz
sN+8DqDrc5vENIaY029HJAiXUGq2QbYo5oHra0NrosvIP/zSEwJi85oxm+XpCpZG
W3sgLENlAWuSeofnKxArMolT6SwX5XZJWJC9Ch9osbhJeQMwm+lfsughG3L4+g5g
IO2qZdfRLW0iBzyjE7Bp4Vodhj9qp7QMp6yFzlhGX6lpLumZkYAk3FX51cCFs1cA
w1ngYSF86UtopiCiUJfrnt/iJb+h9f0VA7h9nTLch0eYYQCEM9AWoGnrZ9BNm6j4
BT5jL7+QU0uKg9v3h3loNlCJISzgSvRTuUrP7KQyVD/q+TswReDgM0bkT5nc0SBk
i7q4KJLxD5h7JVfaLEAVWNmoo/GikiknclGVQ5kou8LZcaupBosGasITUtu1ryYi
r+snRP8goRngTRV+n8lNy9A8u2VmlhLrdtUl0JPOcZpjigLnfi6LJQYPEuPtIEUz
Hr1UKHSjiR6VyYC2phFTdsdD390NfInvidBxITJi1OydukrMB+QKXGuOk6Qe/R4B
vB08oLygv1471JU8TitMbUQ0DWy95PxYtzTGgKS3b33pnlRjn6exgbugBUwY/WIN
pZDHlgfapaIr5xSgqQgHkukNqIfWB7ZPao1bY/9wP4PJezaEq8XzLRJfkQwKheHI
3b6SEMymvIxRGXVNXHVQpn4ypDVM4ML0p/hxaWQZlra0Kiudc47hjpFhNv5x3NeP
Qei+Jl3NN2m34HWsBp1RU9HsHuzhjp2viogFREjgwECc0UkLZfEQgSZ5t5QPETII
ZvE8BTP2p+9NzkvGyTLDgHslrMKjvbdVeai+Ti9nuIEHFcZTJHrgmCYW9QevH1y3
S9zY2NSl1gDSs/hRPSH2nIcTDwD7ycRzWYuXT6z7FwyH1Tn2QDaASKbNCu6oUN9K
o3s/mdp8btq08yWgkXmNob6v8iUHRcqJUtbByoQG+zEzv7luL27IJPouqYGIz8ho
oEankJy5/p1E+8U9A1LnW3DOiVH3jnPFGXCxfYlj/J8/DVAy4K+k2a4qRV5ipXxc
1IvUX6TSEbl22NYnM+vh3BBeaXUcfP2d1NkubQy9w5xltL/KnL6whXYzyBA4TAD2
m7gBw+mH/mu0LhjF+oBsLzC8urIiwkJbdFwPlzC+cMrjTQjdWlCxmXXtllskQxSK
vmG7EZYIsm8BKEV1zXdot973Ci+VsPxPHM1wPpasZvlecTRZJW3bc6DXSRWB+Q44
M8eeEplM8BYXNibU6H/i5txIv+l+BNwLKD451Fk3VIvlDCQthfKE4g7BnNY/GY5H
BTGzDjZ4hBfdzFx/4NOGbDsKQb8pvwG7P2JSvo8ZGTBmmROxWjltaRIdxs6Tk7iq
W+VB85mEtp+sy5NLXvbY2YE6iRzP77JO34HtQ/bQd8y4t2r3M9ERYL/UUPjaXLlz
L4oNu8wzoa4AG1S7HIdPFKDiZXY7C2E1VjsKe7sFVC6SIm9LxuLtkJd6OwO/qIm+
q8wO798a5w5deTTv2VUu4MFqoCP7IQ+ufJwP/XXZFAFo6WFRaJHF3wJmG5gk4iVY
xLRX4GoIletyrhG2C5hBm8a6dmO0g5txEpQoRbhSTURP/GFsCK4Ex07L57Jgo8hR
XzjbEuXHU6m/vpettsK+SP3ImFLUaSAyJLnWOTUsZ7rXB9EhV2Qoh4buvW5S53zh
XLNwAZEAMfFGqEFKwxIgvVjPuY3tMt0vlRtSWAoqA+ezgo7iHWqcn6oeFXB+9CLw
vGshpvwznJYdMmAJfT60HBjr5ZiGRbFEfQio3Yt8Djh3ZkaJeDMbkc3RY43g6WJf
4YR+Yucc01aM7RMJn575BQJCmPPKL12OasX5ILfFhYF/UgDOAAA5mdv2W/J1uInh
WCQ695ha0ykY4YwCpp54i4L2jgKRlu6oMOnEJ4bb1NG0IjYEv+htZX7lnO717b4+
H0f6fjut+QJIQ/bpBlcO+2Wuli2MOk+O8/dNQxf1ftTD4skBqxr8Ks2rYv4SawD4
ikkDBxcZxqaTAI74IXrI5tzPALr5MWsRMBJwOUmPi0aE3c+U2ly8qGaVZfsCGSId
RRn0vRFT86IcbOBizklbYK7ByJqvggBCcFFdnguPyLo1b2YUgCZs33zHcRPsHAR7
eUgYErFKw1QneUi5ZHXtQNHtPytBPokNEyFUsexPrMj3RDRIEnHnOJvBzyy2SOoK
u/npzz9WcTvUtHou386bgG04jlrk2UmHlr6Hf75sz4BwgNv7a5mC7SQRPv1Aa7pA
nQ6r1tDRhognU97pkAdg4mfUtxoFI8RDLdNILu2MstpU/U0ygnlyl2xWKJURjdo9
9wCatSeqrCTxSzy9o9gGNwVz8hFsLWSb9cCOVUrNDFiILHn5ueVT10IxLSUtuxr+
xJNrHxxQizMI3dumM3pyDD7wubkx05K+j8P+Nb4iurWATuvqbUTDjQzaO3Mm1DWX
d49ZOJf9S5Ei2jQXV6/qm47TwADuleAzBYeRTeK4UlVVferAzvkwFPzJXzbDsNTE
ZS/HlJZAmljxtHRK+FTy7aAJ2DNveug/Vg53y/Vg/EjJN60Knx4uf/pyL2NcjCnb
IXSWlOPUOxxHFQAMCME2BFBY2XAVDjAgi/r8zwqBy6oFwykjXMdBDfefeoRuvQRL
Mc8rSyMD5otEKUD7ETLKicOSeQQ0006umqWI6h3DAmZECV3auaHA7O02EU431xmH
HCPo30Lfp7pNAA6hQ0EZsyYiQV0yZMmTTDER4WXQ8UXIF8vLyJ8kCy+5DmjNF1NQ
yeSO8k8YYOBrd/p6jNSZsdtkndwA68DqEjJJjVJp6WFZ0ifaQzZfIYhm+rBWUeGr
H3TY+/+l6XpmQ1LWj/4ibQiy1+NTJp0wwZdxjirUGPDC79tVlb86KtpybbH5ajWx
r6BloBsYh7l1/Ui7WrV3L/SJRtFgNIZYO/mmt4KqNqZw9F530hYtoSdQGYdLL+31
I7VK5W72+cgoLSnNeaZnfp1E9v9UswIw+1wmn3h+CH5GmAE4Iw47BtYDu8WJSLpj
H89fjMwNXJqZeufI1P9bJCltxtktLHyogA4V9a/LHCh5r48xA1nbp4XSixmkIGeC
Tyu6XHXtUSkd4V1ZPihgPdmzlf8vjRzujsg4yM2CAO5THdz6tJqfOzjEkmwz06RV
OZX6+mzZ416TDKNZ+y5IQLbbT39+YouQtUbYnwB8Zjj9Kge99wEoOAqhT3+R+1WX
RWyqGAg9jCf4uAnaZRqYzQfO8NY/14msPnSV2GzjpiK/3aSn3l4ujCN1q5IxmdVY
jB8E77cNcH1L8dDaTUj4+k9c305ELNufo6uws1IZcejqFJK9xJxLIwHHEGbVeLa1
hkyctYXDlr6fDMEEVJfVkcw6anuyqzD8+w0tP777hsTwQtwq36jOLfDc8gaUOisS
iRVkPqGUwQgwimyUVEjsFrV428nMPZR113TXC22yQ2l5171AaNCMGVssfVS9Z6sz
eIn2riW6hwGQFOBWejA52QLH140VObvo1emB5NMgyL2OlFgBdcznZseS6A2k9j7u
qPP617IRghvVBIx6RttAgf53svcfNmN+JCJWoi1wkS9er+XxisLCwZdroBEPf2Q2
Ud4pAyTy1B2BxCL+S8PrHHY+7YYgUfgBEjg+wBAT2IxOzcKOWgIL9IeChQDqrev9
OgbkQLtb+34WvGv6JwEtveKGuezUJ652rB1idW/HYsBTXZRdC4zNmSsrsLlx62iV
FHAUN9fElK6hoSZvrs5MQKHbPZiucOERTiL5d4g/pPStjag4nO41VL23whXOCGeS
f0SaTLJf5r9HIeFxb/vf3V0POxxXhqyw0lttgBQVQvY8UWS0/PzZCIWUwd6KAVto
XK8il/NYAKEUrLe+IjAuEOWQHwgZd5BfO/BfEJdUCCV5iUTkZ3hT2z62hSQ7myNo
GJQTRDZ07ZNWm7daqOownxHBUUGN4Z1vH2Xup+KtUlmnKihZLvVWbCpdK68aH6hL
+Udx+A4vw4ABWaQXggyLBSGPESjOW4NcmBRwQ8dxYn6mG9Lvds8px9b5zH4m3U+1
TUgxzD6y5LJICQVKB72EQ/t4ZFGa/GGhJ+Af/iuGjBZFlKUjTAMyC6m2l/beZaAz
H/toKVBqIphubZJQNmWQbJbbQahQmlc/CCbXtXU8/6u2nArV7P86v9Jh54NDb6ws
BQOAfU6ind5Mqq4r8hqqGGaRaPXh5DaA+Bdmq5toDW55oKp1ziFYzApg/vEHL3pO
kJGV5zmPaCiTUOJD7P5LnDUEZwtN9cXgg3piKhZVUcvrgnX6qgC5wXjnfgUrFubm
oTjDIc0ijz8cqUTgZ5pe+0O9nS8tdqRGtlu0yiNqjyQbsaCZGHFP4xvcayAf0I+C
NvRNfzB/V7AbHJgbH4DZfDDY9CqipfOsKLxf8DH1LroyyXh0cjR8B8WZZK0NnpSD
MYBY3erLrHOXLcgbAyJeJBEErYpiLPkCLPBv3od2DcqYzgtlQMxO/rssoS+SJADK
wgnjCI2chmKOhJ4nQpSx9teohf6w9XhVhMViW3oncXQ3KTMZWxgdZ2Rtu5AJkX0Y
aMdjAzb7GTCKj10eZ6Pta4KtJ6dHbfh2yIGWehPA1V2xp+72BMF6rn8Vn2Xx67dK
4M++7grFOmvqFRrILDgVQlwuxxv3p2FeJ/9pAUMbiX1XYvgAs/E9HhWkriHxJbpM
iDEOIS/h1TPqB8xIP1l1lqfEDPK5Lfx9iHf1U3I1l7jDmy5cGpJbFYPCuTDRDacU
9SzI9uGMwJNKNGzqUtBl3hD8NEPbDlEdLp7WQqlRlyfF7MsAjn6XUdDPoZSc2V+0
Gq7PPHl6BB6W0Hu3S7oPv8G0JvnN/a0TUIB0naLyKx47fNMBlLYH9rfZ3HNoEOJ5
oPHtXpEkQjN9Fj9EoMefsPfyKcjwDr2iWEDahXtx9JFjyIqTfWrFaoaWrBuC64Cm
1jVGqfjgzy4k9D518Eaq5z8Lcd5sbaVSh5OrSCVRQmQRwGLbaaiq05Oh9XJWccGq
FxzWZC35cS6fCEe4+ap6JVzIB7WwmkGsNaw5ZIWjAcorgAtKN2G56s4BupJfg/nc
fSl5JrNueVmZ4dg81HFVS9kEzmHISQ8yhSHL8QSARTg0afh2dpsx1peNF0YfOiNm
q7hZer/tr475LSJj7tVqen4ao9F2a3SgUvoJK7vSMwxVUpSabWWl8LS9aJ7fmIbK
UMeCbdLjvdR9j0kR641+oP+8PuXpxo/c/g7qq4kgFDnhAo7EDIjH8cCHVpDi8aaT
Xb/EFdj9/E/k1PIPAhrl+Q9+yr1MbHNJaDhfpLrbK5e+TMcxN9vgJRERW1cDVt5o
MfJD4XZ5BItBUPsivAQmxAfHJ3QqDP7wVm6Nh+50Q8nbvNqnj/aoJtN0kpknAM6r
o4lcPN4YC7JtEJr7HWZgSJDP8/qqvESTrjPIqwY0t0uPB3b31U/3jBlN/YRtQbZ7
SBhdiCsTmD0Q0r5ttUX+AK4D8/1mL2pp5CR+F2ydqsRgNOT1+JRSAsUK+Op/b2md
7NPgHDOT6pZStniqIMj/93zDdyZAvdAZFKNVAiEDtTok5eVDDkSGjxLimRAGBr7H
bRvbeKsFjxThpx4j13Wy05u+9cwKUpVOf7JlWbZjvV68FvBPtqDUgx5z6q/SjPv6
QAB67fM4HfqnNagsxY63X9tK9lCUrod46Oe1sbezVQvaINoMA2c3UQtiqaEyXPca
4+IO5Q6aC/+zB9ao3mPoVbqXUQbvR6vhbSIGbjO1oCYjer0QYOONvd1Q69xYnOu5
uCLgPrPq9p4qr9AlpMLl5BizN+/UKEdUmYYSEBj3seBeq3NvSXxUpvciwg2nMjFH
QTjDXA24HiedxgjG/mYpbFqq88xuQIAnrH5ncsUzzSdr5xIytTVWyskw7+reZf2j
Y2tPORSDVFhNWSxuUL5r0AeiXFTjXrxtaRSjLPiIkVfZCVXhSjRAvOqnm7EGrDLu
xAathxoRzbBkP9RSY33efAR3zgdidFNif+XygChZzD2OPy3nA+7pPTgxz8KGV+9/
t7G9pg9zkiL3iHWirb8I0nvUuSMIC25syeN6X58eXreQZkBtXpnHxNTHEAcGt1HI
G8kgEPo2LTQN0zBVHduPpAiD1AtRyKExW4d9dvIQdWqad2S6VWUUeKKmRpIxq26X
6qEnKyy2I/df4i83yl0xIK49DF86klgYCeX1YNayxypF4IE7oczPqcfAA+ydt5LS
t1u5IH/nI1hJBhhj+9oTZ8Drp1FbGeOF1+GUO+y5iAJ/rhw9G/MU1oHFrJUxV0a3
jYMe69OwMYy1CUYwqPzRybSOD1F4MXsgsqlOwh+nNlns7qOo3yb60Wb/WXf/XTpL
DiJlowJ+w0OwBfcrcZ8q/FYo21GBri9dEh8lVhnFETe0OjyaiXBufxIxSY7gk5ov
AWxxEocC9zZtkLsmKGKge7kqwM5nJu8iA7Pu5+/WVymU266EShYRYEuF0LDZvo17
3QOMY+RLfsSW0tveq2WY0100NyPo+UxFYgQOa7Vsu9Vk3OqPfhPwNl55UXOy3adR
4/lx0UOyE6Etgex1y+VsHArtAFItkOCxeNovlh3WxWEVyYz9zIpCLNVWyj/KZ46f
Qcs2o9aQUujsak5D3YwfYCK6yFpYK11EkLMqJuMWCtxoRGRxVvq+4Y9nBZKxAWT8
h09gN+0dUD6oQ5tRy1cFtyf9aCQp2kD2Nq7H4cT5FkZDZEnKD1asACWWk8alxvZp
qHT9p/+RW8XUz+D3VcvJbZOg2smnnNHOelYBgcM1xSf8nIzAlhvQ1lEkDFa+LaCG
r8hQUmbvBRE/yaKpYv2bYeSoyCf1E+NhhrhLIhJny361U+IxL9WxsZvGtVg4jVnb
0qK70nC455D/kzlxvXXrDOughQlk6T5EiKKaRBGlYFJFn1zu03S3QBY2WOvi1m59
2MnYg84P2CW+6g2EwgWoFywsGQcKeBnmhnl7kLuE50C+224b57muRZo8l+iNrM8g
BP2u85WvKhBiED3Bp4cDEVBAEbdBE6nsGfdgmR7IxD+twkcRqr9ayGFhblbZdEf3
R08KpwxMn38vHKzJs/eUWqsoA4iTdIlGgUXJ7Hl0OzMBtb+H1B+mXzlTxfNvncg9
XDRC3UdO5JFzhXdtOVKZsAMYKAvf+Edo1DWv1KjQdzDhEcsO0DdogNh/V6x/c6AA
SceXSsB/5eb+3IyCZEde4/h2w2qIo9l+lQwdJ6lvRYAtCm7NAbEmbf+oFjW3KG12
DJ2E7BEnQ5gWEYyvU8R81tM5glAnTlNy2fnuM6tInXmtPYpb2m3D8+KfigRJczOm
Oceu+PhARJJXsCFa00X0Pl+hE4JgE3nl2p5ce8X90Fw1Xjxog7AMp8aGT0Zp2iYY
fd9eZ2VDTu6MvIDo2AdUFZxbOadXaEDDOz95fmn+XydhaJEvBnf2qSuA9EMi7zDg
wwpTZQ3SJTh7j3jgr+Qgd4RFgo6vI+/qc0jECVdRbq/rB4B/2dF/tM43+utTb97l
bfdLMNTY2DfzXdncRhymiilWg64pum0BiaBIYFG9LgU/iDg85fqxlRK7HQXMkrMx
12M2vhI1KBTCUowJhDQ1P+s8mglIXQqQmBva0Wh/9QvXLwbAXQRQra0wHIRLTWN2
hVv2h1P67ohynkO4JtElEHHDfZgjkqXpOvknz9UBtzwB4uzL2rDs7YeSFxRP2DVI
+7eyasceHdjwFgmbgHpydg7bPSFf6YVRSZM+GRAsChrS7ktiVABXKvsACh7IuQAF
QOrErfy5faTgXUlaSJBy/KQXCzZPYAq9F01suZQ1bbipf7XtDIbbk/LfNtCf0fbl
O2UJDmrX0X7EB7ttG+drCp11sy7heCwJU0xVIQMAv/NNaOxL3IGKxxeCB2GnvmT4
skKdKlg9kFf7ihLjabjwYfSWOr+taC10dxZ39pGwZB6qIiMBrGs9B9+ForTwSqmL
7hbWkDsYWJyaea36G78ZFwYQr2ywgFOTTf6eyhNzwe1iVZEULpNpbNxiG7Obh1bh
U7wkRf7jBemEdf5Rx/n6vqETpJJuF7Qh48TQX16mT3MHtjVR2hz2ubl2apBZntd4
qoFNQQIjmL2lUw2FOX9N14Od90UnC29LIwLHf865CiDFQ/6CkLRRwZTiHx/BexM9
VgaBhoJmuUEMJq6aBOR1gmnFBupITzjOgsMGs4uFo7ToBWvNTxDFGyjbm9kv8LZ+
VMGZ2R1YCI9YRg6gyz/eGVoU1y38VKeDt5zcXIc0qZuOo8d2hyU/EK2tKyGZwR8p
HgY+90Ff4qikcJVvMN6HY8k+EISe0x+kQHxlZio6uhqAhpi/fszRRfprVFVTNO3u
cKZ4kcfbdr2TInItpVXvksIGR2YbZi4Akmxho+4zbWSs3n8K/s+el7XV1/W/PtY7
1G5M90bAlcV+5YunMqpaBAGHrM6pQeFOqDhNESaGQtSMTmjzlKlIraZ5mjLG8FlB
NV4dZbiL5ERRszGDQAMcU9tlfi2R/kiK2MOx8sgqFqKeykirgpedEHciGtGoSVtC
wHM8JUfFk1lkwrCsxSpGukOJAlBeMUVJqb+hZqwNccFstLxaSE1vdb/LJxVFcGCs
cOlNlwF3WNoh+lbLuFivKKRyHoY9A1q4XHr2Dcz3lSwR8ESp/TAc4DBZTy8RjFTp
RsB25mXp5Tdbcn0NJjesOIJ6/isBwAwR+ny1HhZMwGw0iK7iFRHl/RsTt2uEY3i+
DIJYDiZoWv/9ZewSqpoKyhw4WdAuv3GdfeUcsPMq1AWDTAB5aG31Uz4oNxx25o4g
4P9LvSvA0Ot3tFy01phZAeLnohOQBlV8mHIYTIjlnyoP11SsdHILTm24EFFYRko8
mRq4jiAuZUf3WK33Gfby7k5cfcNRaoRL98s73TmzK6QB4SEXQaKK2Y7j3nv/acDA
0AKYPFDTucE5NR64mjFEp7PieJs7dl3danbYntpMGRnHFHV5bqnbxbmJeht5hMWT
ipZipYQIF5ea+wUMi/hgNKEG6HrZ4kzHtMaKecvVnWuVqpscKNmbzgp/iMt7lCoz
7c5FGLliTmZIRYAgI6We5UaKDeb+QRwbTH5W5XiEri4d5XfoQBwDsd8ETJlJkuzf
BU46CtLwTMkEruLh19n3mrZPJDGL51hsyBt1Xj9p/92pQtoCt6iI/uQflTuXiZze
G1DJy1xlklnTeozFdGonZUL+HMcyb51bvLDUWDq7qoHLSwdDzRHhQaueBAuypWy4
X5rWaXAeBbCwfzcPrQPOdm8Dxc1my5Cn7wJHZ4TF5JLMeUxyKnPy0I7dGbAqhFzT
OgEoJbHCN8jaR8PzkWLhrd6yIBV/PHE2J2fb5ExkT+dvJNIkSkAiUg/n/jw1ek3b
qEDgV9VdkR4qMYbyTwejVF4nrWPnUq4a4I9vdY4XNrbqnqCOLxMlef/AnqmemWFG
YzwaadxcwsLgZ+VmK7LzRYdGzGkbM7sXOO2x7AiJ0R2WS4wDi61g6bXUpWAIcWUQ
a6IOgY63JqiT91InFL1SlOuwG1bEwhLwX0obtg4dIFoMQTE/782TiF6ZaF0ogT1f
kKpCfECsQt3DSN/avcLUVn4FzC0pJobXRzfcS8F6UTdUccqipeksNCm4/X/mfee7
KGuVNeDjNFHiZBtB+hPIj8/NBsFs33LIeCNmLqmaHBa0hWGjg3TEXMGPSHCCutdK
EKyWCyQm6oK/t4poz9YBCm/xYn9rlzKKPks6toEidvdCoa3xpBDm929hVWVC5yf6
/2FEA6L19yV86XTDoaQS4msN0FQXTbH0sVKfbeuELdEFq+ci08DzHQXOzC9yrXU8
/G6qT0FopN3gCiKUqsKIClF+thmpcylVjuPo4VHT778cK9Fk3DTlltMcgVg0vdks
Yy2TnPp9f9pP/ND4aaIv5LSvLUl6EEY9nfUpLKta9pmL2qzZZPQj+Oq5N9o5wfWT
1r+hTQCtXCfYnPofCEbO6QwQvpV6Y1osINLk0vYys46z1BB79I3CJsTq5N26rbuv
YcRtiJ3azyyrf85ps2ucz7jneuL+4H2TP07DFm53QCRe/+T7rMc26nZI0FSRCWx4
c53k8C1N0xJy0y8r2lLj0lWTKODaheTHqLTT0lxWqfW+ENBuK5hQT1RRm7+vynX2
h+L8U5Fv+RCQWFvyXGRh242WQsfjzYHOABs0WVr/m+R58+ohr6ESlrc7gSpLJRSJ
T4ldQfnuMFUjuODbobcntqK9LAIy137RwcTVSBoIBSYlIwLqMiuKUqvpcF3I8GUJ
VlP3kpkCQzpGS//Sghle68Xo7fNVrcBkvLCn6R/jMej5Z/cElRPbsUcQCzaCgGcI
v4O44taFypiQAibAoCH/wj5zX3fadeh5BbylSCnx0cQcLrNwKe6c9eWnwOHKaeoQ
wmPmUxul99PeEO08fZHHXypNIOwoHDdlrAp4gOmv1sk2v9YCk9u2bC2eu/Ct6uuv
CKT6VPr510deZ5j6TJyoBza3cjcR6kuLfOBXwQovBdcuwmQqCjCCMQm9tO0h+AGy
2B5oWuUt5DebWSV6mNX3zzr9rBzcN+mRJ/jPxCR22ocpGy+5rho3u5dOENERKqTT
i5w+TiMVelPjxSFjnbDIz+W/5ahPve46R5HdqUwAvFZjZH9Nu9nnWsm7Qv8Zwilo
pOyLe9bU49gWOHStxFcvlF5/BiGtK313FqS3z+EA22AzlV+LJtO0J/pPSJ0UzDp7
ls7MqYybeSF1w8J6FlsOYJW37qwbfgbQMQBMIpRIRQRuRku2sRF2ulNVEoyopuzF
APqwMJKoZQ17sdjBtdy9p0hv/y63h9nIk+5IHVsH7KW/tMpBmCgBphf0ePXGMB3n
KsS3SJpJU2hb7S3V5bgYLNe/EvUdpDjZKriFEm5Ma2S1hMte3YYIlYSBerRGQhAY
EL/ZVZwFGTyWo1t5A3uDleQWTwHiuQeDd3gBAF6iZ6R1ozpwA9WrAR71cM+CAvmp
eWu2dKU0W1s/R7G42Pxtr35/7b3kjD6Fy/D9z0qjY2n34i6+aHphWQn6m1UIOXBI
0sbT3ioiy+J4JPZFhkMebx09D0ETeO2oeUqVRPeYnPQrJBOlrs6rvkrFhwXKN/4b
LNmo0YWxRm3ZJ/SEhgvSi03elHMUKTR49NId9PxX7nE7EZd4ThDUcRVex60skevG
tjJP7pBoihH4KSuSFPoDM5rNbVK5Ze8OPoDyyky1LAPsUM8UwvvkWO1nDiqB5P3+
B2xqqxa7OhSy1Yz6qMT4zH1k0uMj9dZsI3IBB+Ed9hOzY3IX70u9kt9UubpCox7B
jYbj5Yak8k3R28x/CB3e+giHlMV0Atb1SyRIcqEg+fIBKcdKIe41lPHpgeaVeWXy
s4YLpLQeR76bXEMz+29XPo+YSiYV9hOA+oT6pvtVOpIHwBWGTNe/b5NWvtHoXCTa
vUkSApDOG38lQheim1NbGRG7f6RM6DoQS1KzmUWypy/DEdVmFaCtPfkdRR8sEEHS
Ch7yAXqcW87D2d2R305hsu3VSRW5a1mbBYzpNFXt6LFAauWEuUoJXPHjAV5Jsl3l
RaY8mfKZQsXvvlQ0VVBmCzVODBzxqH+U37m/NFTNrJrlz9cSZ6AFbYbytlpKcObY
WbqtffvQEVq+/jUfNbpJVjB+iQmzOxHBdyKL5RWZEyih5H3vEHWPjArFrRksO9q+
hCe7ZbMz2hgtp9cWgGCUcB8F77nwqLvJZkwpGYzxDLDYYunhR4+iiG67KIGiEmEK
kcYnXaqypK9Wgmf7IL3b5tbq66tbo0mMkI9/lt0amczbm7J5aReJXNrrXKwsvUgW
PWCiJ+tQjS+g6MwhP6KARK0vSgpwGOLwo6Z0qDM7JrGYWMOj0V0NHKZuzt2alw7+
ifO5U3Z7/lq/hNCPlIMLxK+YB+a2VRMGZjnhgOjx/jJgqUaNXtWTvCimXX/G7wFb
yW/HF/lQGS4TXdSgdK3+4/mRMJSYVJZ0tbYQck5gCRqIKhAYnKnUy2SGO9e0DF2f
7HBO1f3De9UTym19jocSE0d6mxDYTiOrRDP15HswbBmrMb9Y69kNqNDnH+UDw0ek
RTbxWRCSXAZAy8P6Nmih3fKl++I8C+bLRywT66g5MEpAirPnO3NRO8QIu7YmDjsF
4Ht059GOGy1ceT7B+lOvYpqGc00ootrH9UQ/IsVM/x2XhlN2rE6I+Tyogbl6pH5F
Coej7/y5zJXTrYihjh5VIR56+2s3v791hYyQh944bYu854ZhCHqVB6iS4sqFcGUz
YaujlSnNqQipeEn9FKfoypKbgPthibN7XraKyRcBw7SwnyB1u4pRQeP2EAAgQJqb
sJRwl5faFzoDaSItpOf4Q4QYy5iP3Kcntg4IgMT7wfZJoXuE+ZaNhSMmCBKzhe6B
CSfUKR30kAN9pLe+cUueUzDlRhYQTfOV9ayCWFGdS+a+w2YwiFhDolXXU+w9hfcf
ikO0XXTQKzehWr2y+NCZHfthZxJ7Nd/OsnxMkoK2MzK2wKsl0G7fIO4fQ0r3OiNZ
QU4hL1NqWbBKVrpM+wI1Va7cW093zXkm+uJP+KGVQJ3j875+n0a3NAEcvNy2ITEB
Ywvocv450ptanE03m7O2FB0foUym+PJeOyzXDdr+SEVgjl3hB6sKeklosvaavffi
mOeMYRYD+81p+cxYF8HXKxjIylqIfEvx8tF9Nrt6yqJo/vPIFm/23QbQwW1IiECo
On/KWSXAVYEBIln7hFKbrvHu0TGT+z9nmU8/z/AArN8ZUtDpT+YM6IPir3Vke6aZ
8NGOS2AzgQAFTU5+353ptYE5hz1ZNUhm+rISzt2v4g5NFk3ZXBUSZ6wXwuDlaGyY
yeyeY5uYbw6ovdcywllRzJLdMC6eTnnhIX+qV45NH5FZk6Fq8zAXJH+cHvJXQI+j
+Vs+tD3kJS9Y+NYlZ6XTlMMc+M7+AX+IAKD5C+2tpdVC1HjMNaADiG2ddaSbGBN4
ZaQ1iSFreWZ5rWUuysh6WBTMMNKrafb4lE/mXyq2aG0tmzxrddlqparHdUL4ztUu
frpR1UPZhIQ3V+b3qcjDQcRYwK6v6n0W9fkS1fu4spQNI2RN6Cy8yYnNaiGT0xYd
zdDzxk6z3wHdCTr4gljoCIYEXDfFR4py9IkFlJJt0vGsHGbC0IqMZ8xCzrGrJxEl
De1dia7gGpAHevywsxj3qJZkwM7HnRNmdzdmM6PbISFrJ8s9KO547xf42FiZ0OPN
dEcBpd87/L7U0aLr9GeTtCZ0W0QNaeKVqEUL9ogOJUOKBezXQ1eHwm8lAsfZkIDu
k7DoZlPM48L9/M+9RuccuTo7dTV4zKIfzKIx6AdUYIHIm6kSVWxgzW3VGw8H8V0m
LCDBQfAQp7aS/FKLk0EfS+zYFqRL4M5bYm8nN5svAbjdhs7DlsuZFcMEMlFcv7K0
VbBBtI7NoXyYsiyup04yYZcyEgjTUElM+Iypmn6WEF/Ba6337Ko8Xmou0FBIo4rs
xBdubl/wLR9mJWTIaoT6JxpbfiWv92v1yb33Nr3+Q0Iw+qi1kozP+Gmb5WKxVqJq
fpubbOLS1A36ex9pZKNLRfVNB/4wrJ4yT6UX+mBZCZ+ZVAJS+DLhifysW8ileqfC
tcpfiPYVzoxvidxMG/jwjTnQhwxaQMRgVGbQJTp+fxpWeN8PDbc/U1BkTBWY1tDb
yl2UynVfPXseTDo4jHUIj+ZbE6Ko2+EMBYZCQ702CR1rmvDVGid5bhNLwG+f0e4e
Sk/gLoipq4CUbGSsFmPwbhZIN1w9ScV96iw1V9F/haaqeu+rissIG8xyvX4thkx5
IQU/163vPzpnY9UVcE2JTcH7/beDb2omuoNxa+YHSDjAVPtlCr2yDZ7GDyLI1eYJ
9LJp54zgm6f8Oe3ayodyjE8vigMn+rgwIXFn2Q0/fqxpLt1lFD2/zcJVLCou4aL+
rAkfPnKT/LTX6uBFQ9TqZYrK2Jn7eEu0L53wtEtuYOqzXhiDt5zYGae1xHJfc3GR
UlZt5VIPBTIzzd0dMIctxbsQTu0nN/lZQVoWSJfszXOppdCpOqFXhnDB6KvgVcT0
RhD4jwNQ1yzhcoZdAeQWicACDNsVFa+kqhjkQ7AgNKBZ751XgNw8Pzga9DWGRgZc
FOltVYLTtmEse4+hfQvzDhHMMr3GNT6zTJCFkObszPiYoxzly0p8UOftFcRAfsTs
vptQxpGeWtlnDJx2yqgl4mhdCEARIgkujymW7pNcRWcEcY+CC2kPim9o1bjjDHyt
NQJkSpr29IqELuwvFex/5V1DBBmJFGrTJq7jcsOhdiPeyszo8mMuTKIT7Ao6YH7N
NiQaDFEMGSytD3pCzDWQ40/fbwPZYKiey1g/p+6ojbEpf6FKjF/zEJWr1U9xF0Zn
bkHQtMPFh/mO+BhzX8CtBGWyZ2akFDm679UlL8vbGmVy1XWYPT8RUyipk963vFDz
zySgGXXIW3bEsk+zTWUp1NIgI0JQjAwE/uOs10uwQ7kqnKuUCs6KCYJVs2O6oTJV
i2LB2HuOtHag49UW8kHz+RWU7l22ERvUR2Pn7VN8b36mWA8fcmH2RdUx262azGoB
3aUEMUdpq082TzeVxTOHgoxCGRnPzzQj8l/0pX/ul56LsRZjOAf76KCsnFjxscHn
BJeVUKudss9NGfEBPmCDyHOT3G96uXr5qgqRUZVGN9rIY1eqj0tVunJQzdybgvoh
6bg3a2eUIV+znEAPtZl05RynshBmBk4UvL+ZOSmnCvN39z2+fFzokCTD2GbYKflo
9rnYiO/zkAeeGsbyotwBWxF1644ucRZZqPlECAVrStw3XV80BSWcEIam9cIA+HQk
rd6Fv/QHPGMQiXSFAKxHqTYj9eqQxeQRoaT8t3z8+Wk139i7mv6ymE6dwReT1KHL
TyEWs7OOokIIlqGsaMdTRl/KIgqWkCjiDblxKqcLbd3iZFy2fYKHrFPbViAsmR9F
3I2KXrgDhQiBLHhkNHY5Ofsg1f1ytic512qo3ESgmpeP30Il/syO/eCWpj1otmuh
f3VAhzgBZsjGWPrfgokQNe2Z/27LkAy0q3j8ohWBEwL4yB5Dory1owOIZi6e39o0
76K57c6JChFRdmz/tW2Q9NJP/ojBAR0iSCyUpLb1RgNveL1nqRCmx0Nuwh7mlsbL
mB6PDyR52MOKRXvPEag8hsRnK3Wzo22kznpn7S2+ZBjlRudaUmoib51QYJmbcmwd
Lrx1mbKk0R6PaIpHVv6dIJj17qCZML+LE5n81isbzDVebwyLltK57HByVKhPEOye
UjzSBQvigernyqnz88PqSE1W6aVRK9KwOTuhhWv+CWx8HC90/0OZwe8l2xbmnD7S
I4J1PJPldtZHFwkj0+H6qDoCMIy/ohl3+W1fFqStLjCGKEbgOXVYJnIx8lF/Zlqe
ZpevN8HdbaGXUOCtUwvOg34kB3IvI6Oq6/W0ANxMhLoo2p51TOEMHfKcuq1CQ78g
ObYhWQ7z7HNt7cFLKYoBv0ZaP6NhB/m+W68xkitTOOv569Kdo/RJj1m1Fy2wAcic
oMpB11glAtzG/y5YaAKnKOfNC5YBOW7Jzt0Q0K4lQAE7QyTbsg93+DUnBq/Gr+uH
muuQ7lHqyUCYmxPVenkAiDcq8gUd8vBbAvw5S+AdqUK9mhfs1IX0xo//kRgPFHBv
opqaU3tj9WjqthPW0GYwESygKKHKgdBzRoOdnqXEbVjxe+rr11f3FufcX4WTubQv
vBd30MjhNvhSnnefmoAi26RfEXJweXIjVeABdegZEhoXhGI2XdJQz7NY/lFSdOJI
5QnwUSFvSWBhmw4IM0wcObC9BTYw2tWWin7LuHQQOUwXTLxElydD/aZxZWW/cq28
jYLqFIqTwnIB3SjpWwkHNMKmLfowerKcEHScUyfWWgmf966x41NQtZT0QA/l4jAd
BfhFuQx0Q9PzKjQKL+ME//CKCLOPzhL5Pb/Ms6aKGpG5bSOUUYs8O+wxyjy+hb/V
8YCv1ol9n8idkx0y7CNaByQhHcZ3n0MWJZeNeUv/WmbSIQGxJwHLvah4wVUhZyrT
c+wMG9/GOJqYjOuiP05QwxHSCt4OiyLqMH1p8qYc3s+jyWPD0aP7R39YCn9p4s+3
mfueZpJ97mROPM2I5EY75apq7eva6Q2UsGTnnKEtn6fdd5ya8b7jS45K0Gg89/nv
PgN4ndC/6x9o+hfGHoRchKEFXM/2SSfSgUH4b+yqaN1GKlz2WIxEYx8IGpz97W/Q
Mq5u0i5oMsXbG+NqJe+5oRka/zRK5UYrMpuQn/LvXwskiKvKIyZi3/WgAVcMRS1/
n+y2XhcoTeNp5Ki/x01eFFHfS6Jf+9pqYlRLzFFBp6hfpBJOpjF/8g7c85C8SPPq
oH1Zz1nnHYs8TJ91N5g9h6c3/55lxqDixlc1F1b2DvZoJJ/d5UMrPxRfEfzdp4jm
D1tKC+EsnEct/zH3xXq6WxZkm+hCecjzJxEGxESYBFE71tSny+2OId6QcW9jrTvG
cdkqzdAuN3c74j6zjDonmmUDXdvy/xnXl8w2CfiovBhYeIVanMFcoiG052bdJEDY
LcDzRDsJRN7vk5fQUxBA3LEG9fwBSLiEzky6XXFq5tB96exdfsEL01D7ADw5ZMZm
du2IsLbfCDVk6OlGmwHOUXc0F6bpbTIs8err0fzT3GPbwMYELvOBy2J5ecQAuP/P
h77ZzENbh4+W+prrMv7TxjHHy0gR71JqJhM+t3E6zq9VSL3bbqVnr0XB2o8GEGa1
f5wJMp82960ojQfyAleppcAuBSCspZNRscurT+uV0BIJ7ufnY5y8hk9eCotzdscr
d6qzSsA61eLWszgfL87/MQ==
`protect END_PROTECTED
