`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hE6+iv4r2RcULmxZYcDJWkdCXqKpDR0VTLNH2UchWXVd2RWJUY5T9M7WD1SUcO1v
ToqA1bF7Tmkvqf0Gm65YwGy6/TxdI1hbpq45w1OuXbdyEhI/8raLX1PAQuN5VwU4
x3v7yXXFIJcoUEyuG6FMg/dej4ZwuPtuTbe36VllZ2G7/4BM1o/JifwGRPF+1zdv
tUwWuAfwCOEI9BcqtBUa9nRKoFNkqrPGPf0GCunFT83xpZ7KyKFXBdZK/f69ORh3
+eoQ0nfWdQndDTS+qVtmDrZbP/SqzqPNOuR3pmDbIrtT4H6ZE5lUbF7dpN1auZsu
UMsxC1SQQ0ltOv0lhkC/h3ZnCIQi2tC/W3I5mLH8eUK1O+k1FB3vKDMC4L/o9Qq7
9yaKrybWgDniiKQD0iHcyknzElBEcqNH1HLVMb4BIcla76moEL203Gj8pVGjRSSI
tlzRT/LWD44WUY93K1DSg+iFlAlo5gXhfPcT9BEvbLwW5tKu/yqRwffhR9FVIjn3
UuMp89ZCOjTSIIRLBDEPMmCb+CvLQ6NHulTg2FY4F96BhLu1Yve+KAMS5aUw6/A7
gUsOjaFumqIfEQQh8LSRrLjb7etuxLYfTh7Xsix56zfbUd+7cx0ra2mi1iVTZyNl
ttf6wTCcUxz+1QAebt80qn8oKECqtG7pGPFgiiWbbVOmG8pZNxqyir0srJy4+fO6
KY3H7gYFgOrUduYLYwNzWxTbcKvvs8cZ/hOXS8BzIMs4f1yEUm+1Yz9cV5SL/aUw
JThVfTCmu7A/XKik45WpTszrSKmXg2mnfjLaXD35s+sHX3Rt5wCYSTbwXBoR1zAR
l5x0ilr6WY2niXwIenHIPr8GXa55p72Z0Ax6IH+1lqKq3LIupRmW3KtOt+2DvAg7
flsKGwkSb0MMUcEKD0dnAkIq+VWEFSSW61IQa8UMqcUpS6g2muxScxzVXNG3+n+2
vIUo5gUxDRfvBv7MiQA/wPMF4AG43Us3l9ddRVQdN6/8PgrEoJDUCrjNz8JpQ2YF
XwAi0u/HysgIBtbYxPEbL/Kgpl3J4HmYW4bxmtiq+rZikTjQ90XvZHVA5np75N/x
Ax6M0haffXiDKSAOCMmKGft7c1hw6DWpsqk1g9pa+rN1cCk7Gd1dFjkXMUmig+UY
mrb59b/V8/fxCovalW63RNq+wWRkxRZw15vo7wdOa4eI+ZSvFJpjqhHTvYdVPln2
N39j2OTxkWkxgAtAs6V0J2KgaZaJWh1ZSWbxqufQBHbntnUdIIOMtCUv1clo/+rG
ddjvvVh+KyUipiEtE0YpWhrI+9c6U6YJsP6JyevIjtvcUWm5DRwSrZ8mEzAGaZrP
TJrCwcneNWuRblITqjIB2qYAAtHIamZkhyeqNrrbKiNm+6rrqMko67ZraMG+x/TL
dPNvZNjGULi7kSkVutzjks0hK7J2nqvJxfx18+kquB27obQiSh9FT2/lmwaQR8uT
oRGAk1yp2Ljn7zLqqEdxwWdUO4rMygChEDvWoZi7E3GnwoW4hbZIowRUCE5hJ+Ty
Mg3PemhTMkUjEbm+vCiVTgzF/Ou7+f5EEyjj0EL6bWOv4SulUhE6RMcJud/b2CJo
4nsT8cVrNjyO38/Pfv1gu7SXJ62kMMKUHApdNIwcR6skpjExx4w0gMHP01r+pBtX
FNKLFl1WS/GoPMs+M3FIf7YyUlkiC5gZ6sUT+EtkTZ/8DXLEqxlfEmoh/NzSFeCS
jIfAj8b/b9qe2LgHLoxwe2XF9poEtwyYpYFN0tvBzvY4Uaizl3a2sDNGELGICjLu
S+i7kltIqi+rZ+f7Q/89YVBW6+Ht0mkKM6uAm47NDv2dIiFZf17WqiCGUp2IGCtW
gL5RQbfFKZXamdjxknoPAKJpRUrcxhAE2aznvOsh2H3cMJba88DPkfCd/Rsqgsdy
j7sm3gpAmToPUOd3RhJqk3DktzW7OevAc4klKHcRAgFBn+Rc5ULiyxRD+eH5GbJB
znMX7D379f3e+0QA9uEFmoa1biSiaAE89ChA0ftLZU9nym34a7B2hEi/sjCCxhd3
sRdT+tuOZ1f502zdGp3ycaZzTNlcoE6CzZDi1wT0g+x1TE6YiFwqaRjMcdVz39Ok
ehNi/2g8/flalUyvSv/n27+zozan4ZpvpOgsK/mqmRd05EcSB00jToTwetTqqwQ6
8lH3rP1I6ErcKDfO0OOddHuzbY67kbb3M35hUi7EquRWmcQ6fzIhV5176lmYXq3g
xZeWwjMJmGgV/t4GpCZ8UA2SMxzRhWQH69AsGMYA0A+tLpYZZujHwk9EdAnXunwf
mUOSHNvOQRImygX9N93iY9la06ubgygFyGuGBO0N8U59bCAOvRHli8aQtaW9c8Cf
l6u9IYVQxP8BL8aKC2PlsrDZLsVXkO2+hUEyj8PpbUKZM3MfgPMsx3v0YiZKbDHC
Bbofh5S7zc1swBbVVTNMl6/MTv4Z81jHxJxK/GxrcZyhKtt6v12wXx+9Q5wpBskl
SoJDAGZxxhx3mUzwP0fnRIvDMNfoTUZ0aqJl2b2I+/NOLiLZdoQTGNZrEr0a71Fp
XOs4FOicxU2mNz0Iyn+tKfZ869yuqyZrTMdFaY6IPRkD/d4T1UrAN/MU+Y7OIlZQ
wddrHSykp2vhSLHVW1NfIGnrvdl1XFL/VnBmHQNCW+4+kOWWFpv2J1POpq7K2Xiz
6hBgsQ6IWBiFCrsvQohXBBzG7Vk5IavTNeysraLSIWUbrcrc7JyB2sFBAU+N5Wqo
B7yHjk3JiAFKlQM9nvoHMNQD2F8r2V/8nq3BA+D+bvawKqukKipgr/S1dY52eK7P
5J4By/nPQq3VLg/q3vUaCIipTVIlL7uxIvTWTBQtVZlGNPMsL/miI2Zqj6Bte5Xr
6ERsDBtbYvXIInAYz9eJbgqzAzIUCVwieWFk/kAVAgdB/5r7rlt+k5miiV2XbP/Y
wLfJdNTD70sWemRpIXk5o6my3MRvPQEGxu89PUPvVUpfDHTz6YMUZ+VK/xXZOk+X
C9J1JioPYGfKWC84vRdYD82XHDkpd1RUCWEwqr8YJO4TWvqAaZU7DW7qUY1VKMPg
0+oqxLlfru/snG6rICAkqLLw49XEoJT4jYsyvvvahiOPbKcETlvrpWOckKvKGGdD
ML7atOAuP6HY69TwnVRwxM8PJjTswEc6cSc7LUJB2oDpeDFizcYlZpAcT7UVAr3B
TjrDusmX6s/wu0SDsFECzJ2scF0uC5VeW24OAxOK+ZKAhvcag+iBEAhqFYFfuvEm
FhUM2CKL/riXma73SnyURUkcQNW8Ni8k9mX5H5vaf154rudVlfNJDbyd7qygmdYC
MBBo4QwF4iz56qbCQYUW9qhu4vFaJTdPoW4TSXvJpOdtIo9UWyBK5HtxuTUHfw+T
J4asSJFXG1FdRimY5UjvS0LAW1c3XmUtXivoOs1sDrYQImvklXDRTFabqqkllKWh
65rsdRDt1XaIaqqQOvBVpD99AP49mjOMfK+ttRYVadpUpC3R/r/LWsJavmZYkUwA
2VTGgwE8Lcz1aO9cEY/JPYNdjY4ruRYQpazzZ2SYi+Ame91wjRBFsmXQphGdeYDM
I5LK06O4Ofu/+107Qb4rCx4Yc2c1JeQKpRw/jL/JeRaXLKqWcP0P5aIDoVNjvhqq
7giSUkJDX2tkDwZILtzSvSyI4bzF94VDnMRLdqcS7W+Z+uQreuodl7fqWiVSZnqC
ajJKJI24uNGlZu2NbxPwFlQ8gZa0IMyhLusZsctf9co/VNLxGOZ65P2GxIYarm6w
81bpZ0RYqdvNLEo5Mt2T4Ziib+5Bpu2gDUiv3Ym1SqiBCSY+pG2QXPxQjJEG+Lsi
/HyWJapVLttiJ+15vQMItl3sakDt8igKx51C22CsKOQYLvKKc0UoieqqaTi0Thx3
Z4TmAUJLUuV848tQmUq+cKNGyedMnMNsVXHuY4MkudHV7fJ8eIDoRpYUmmpXFR0z
5SUSDkVuQUxCUyyZYozKc8FEyTl3AyBv5DYEFaMnrl7u1e7gCW2JVk98lhpwfaFJ
ftczoff8Ou04mPbPl7efb63uZo9IzXREdliMaMfxIXOT1cZobqLOWD5bRleCW3Zz
9mnU75xpCB3/M3vrriUqAgKezPDD4MGtvTLqXYvizFXw6BR63D7kK1Dle2q7Eg6K
FmE37GyksoOJt1FT2l7OuneEz6ovgvdLp1GiiClJiCE2lWDhiG4DqL7lrRRE90ar
6rigEYz/LjDd92w42hIQufPfSf+aLvZgH6iEREXnXtZ2o4doQVz3LH1Y+q0vCuAF
DWSHwLC3Qp0P/Us0b/WIxRoX6zu+eTStz8OJZmO0M/oZlIowjv5/mT3YNgrULmOE
ulQt+7+xCoCeJBNXe2WB36nPUFqYBT44nU5MsnBc8Ue53k7sz7ZkCjLf6h4hTUzp
xl6jAKdv7z3E2396ht7o7PE3lVQhegOmhhB6PlR9Tv+7PEZgBnujN1EmZVM8kQIx
yy7m+HZLC9fHVub1wl5ym9Qs4bxvYMPzMc6n8Lv9UcoIm3zqJE5+GLW9pN/+k/zZ
D7qsQhTYOhT2w0lrayjkfOCPsWdOqR4YLvM7JcvX0CbARUVc4Iob/ak9xvkuDpAg
3oArGZ7I4wWGHjs/MJNKUPVCIkf7TxAtp26Izrdw0NiyOt7GQMDlg7F5P3mPAG6L
NHqA7DAEhyq9LnDSuMF1bavjDOMh6zdqxQZzYFPcDSPcWeI0w+bKoWEeizMoVhJ/
NGMaZNwAExTaBD+pMbrBojw1bvl1S3v52v6edukCD3GgxWw9WDRp1lLfibNFlJQl
aABVhTBPLZ028Qyc6gWan/6gE9rvIL5m1JFtuqUmBdgfsA5R851DfgA1ICGnECk/
CCbcTZST+06AD5EL7mMLk+DcAS51yPDlnxWCn6ug8iooXlDe0fxzH7ZTpQj11EGd
tgJ3AYv0KS4FIRU+MbnulBdQ5LKQcWlcFQCUD/UeRL7Gua4ZetOceRw/Jo9XCCyK
F80omR+YehoZVG8+zQZhGYqwlrQAoVM0MNg/drtbY7uFRvTQ/2pdCn5owVWQNKhB
aQKHSHLre+tvYP0BIuKzwCBt78p/mMbhSGXtFd6llTqh7paUMedOkiwILVzARO/6
CFXc3HmxtU9O3GqnEoNicWcMIx1Iaup8ua7WoidaFOuEZTDutLcARbty6pw+qMdb
WqXauQklH4lk6ISbNVIT7H4qOwdM6LcoZzT7uXsU79G/pbCCV7IdM6ltFbIZmDXL
Cw1kIuYHi4l6VNnKVBXxJ8Md94Yq25iijC27X4UO80kF7WH6k4VaV5Fw+3SzyFEA
8BkTtWUQZoMncfRcZHhBGx7ErJm3jPy3c4ai8UsZCvA9MIO88KPjqCobSDo3Bl04
lbwVUOS69cHOf8rXN1qBse1SU44Fytq8P1Bl1yoSyys8oe05KzyqaqWahbDXHV/y
m/6g97H0JRvQWSvy6SIkIlIC6SYfFHMZKVbzMyjFGvEQeKUY1JttaHiXiAR80mOy
9fhVqnOrzG1XBtDHWAecwuNxVVhfO6mtd/mia/Ah5ooFy4l3/YT64z2dC9k9vnfD
JfNOx7Fk1ArnfD2vj3+nScjz6xHHWF4WjufSuJmsb/IP4ruX9z6908x1yMmWpRPo
pzXzmmdmNpgOxCd+ekNxN0LNlZIIn5uc8+2jIV9McRhyk241drnXQy0mw8sHi38y
V+rRz8UHvHun5bWS7/mUCd4ZLPhB169olv4jgFIYwFzw55M0ZvAVArI/6ZqZTD01
X14itg65/3rfos7M+k57HhxGqqgL5PiWRq+JhndI/nB2EmTOXtrDfnrBNRgZZYiD
ETqyuFceogdtLo3oq0NjyhnLTl0JsoMkdt6kpP+h1dEfPhBbhDTLehEvURh/wCWG
aQfNSLt2Epp4Xof2N+hN+KDjjORWgwU8sqRcwyrDXP0yjO5nkV7qLWGRU0X5jpfX
SrBkZZwEjPcIp2GyU1XT53ucNRUI/ujC2LsyY9OWwsJoxw72wufoBl/L1JD7Aigk
mVR9xMYcOITzu6B7GttXTCCV9l3syr/T++eRSmMFNMI5gZAEh+T5FArHdAWBfE70
+X24+/BbbNXRXarNEdeMhyiaJuDjR19Gz7EU8rsjvtHasKav3Khq/Cl41vy522t2
NeYN27fpJ1Z5fiv7p9LbX8mXtNsSzJEtu5g4vtoGtZt5bmmerhMRXPXtFEvlKWzA
1MV3UMmnqQgDTGn0j67FoccXezlsYpIP8UVZtt1axfJuDJnPRN/Spq+zREaOq29I
X07EedJ+cfOsUowRQHR0XGafNspJGTcKJOlfzmN6E+NZeF4Vem4UC8+tyYSI83lC
BYm1aq1CHYhA/+aJjfSRJrgTHTnwNquBfWkPksDzzeXGb1BKfGBPycmldfhPKEZ5
F7RtltLe2T7QlyDVInIW+QVOffk1/MUdf9vkuGs0GodNcLpFXHINrTgdJ9/YLhax
FxAgg0ZZGCJQncEmitg2wV98A9/WDpe+7oqxBv4tdmlG/uMzWOvN3VSEAO5kWDXD
iR9HOtuaBqIUBwkZ2ux8tezWA+LPAYJ6SRCs7xj5WJX9cvv00sQO2vXeermIW5X3
BU0EpACtYpIx6dGLhrjkBksoAPaFE07tSmhn/X28x6N+ugrL3E0h6+qfmVRG2oPL
ptUprMDVH/O0HqhdtXQejxKmfMlntL9ozIiSKRYNvSTzzkOTWDQIkJjvL48Mrrnj
GIZXnlx5xmd69CnbRH2RvnZ2JtJ15W4j2OMClV7NRJovWpAy9nswx+XsqAuRp3qZ
N3wOX3PljnJZrawQxZwTQKrgx8bgn0rrh+SiSpNj+LfPhuYN4MmbdDIfvLPCYGlh
O7ufVQa6itwdvpjWagHMwx5BGnKWsLoIRN1nX3ia2fX5djCa5bas0AGKxXC+1EaV
MAvFp1BP9YDKLbPlR9KF1PitjtjQaFi3cCRJ+bZB0KLX7w5UsvRLmAOmdeeyhNBd
5JOyzyFEgp3m140UvUdJBezvEMrbmIh5rH/zjofCUU0TaqZEp/eirDFTiXTX/4Iw
KmSucMzsMhkxgd3EG3LXsqIG3MtEE3n8tTu3Z63/ev8ideEPEi/CKBRn0/dXjBDN
9FDnYiiRqCd5mFZopWHT+cqi5zEf5GzCgHBlp0GKtrLmjlPxFoGT9K0v+/dAuLY7
11hTD+JgUUEYXPVTUmM0ohDz0CDsDk+QiM8MiWHJz1Rd81lxvu2SM+tuIFoZLgcQ
1P1bZZpMoSinTqt6tanpscKRcXhFg8RVvtDyUDXjwntwglDH7fJ9dvOZzrkwU9Gn
JEUHlNOlVJYCTf9h9YL/FvxTwtYtfdrlDPKlFu5najXk5MbGcqwAwEzYCDrefxsr
Q27/4h5VB6VZTxQJsMRcIPZ6+9brjdBvKgGJW8RkLTU/UUsEfJpIHaTNrP6nU7JY
I37HZZVe0YYNEpoxTBKjF5mQRysHx84b87swfLl01mnOrpn8dXKIkWWFR4xLroWp
QMz5S0WQ08c0CfJo27Q/YLXUwDRdX2ErK3ubCKZyCwWNksm0GBBlyBu4aGIVWmMx
PDivzSGQfa4vrutRWW9yOFCVuzylEewLGromRurVRAwK8HDhLh2e4G2tD//J2u0K
4Ilpho3VdajylB1pY0/Cl1JSZK4ZynWkaaoex3a4vS1lDezrEmM8Ri8/VGH6tnLD
g+J6YOCWjS4O47tZaoaawLpCoZJOo5YVe740CpFrH/5OzvQ0IflHe/qfIJ09dltt
P7mPnuB+OB8ft7X8qpwLlUf/f9CQpspgPd7IzMeEwxesEVxyTnOwYe3E3a9yTTU4
WO2YDT3Iioe4kIY7r6KrYIGGVaTOkB9b6gC7RVDh8FkJLSDm18EwuU3I17vs1m5Y
nRQx5FNtJiQsMDkHRTZ2szV+F4GGJFlMHkEjmNbA2y3Erf2IyqLpT0r2dN1Ktt85
z7qddmfkfKnYjB94JLOHwMz7DG8H7DyT30TsIwTOgwUqC3+E/53HSjEJ4cbEOILe
XsZsXEXJPdIXP3LOwyPMgjrhr4yATnqwZmNlgtnAibY+WYHz7mWX+htDwgx7Ltgl
FhAusmlk8Jb4OT4Oxg5k2V633X0BjlQPkH+dPG4XZE+C6dAw/ZvXJIhhRsDoXtDx
PKgxLOyDmJ4UukaRKsWpYLrHkMVDE4C/CQDBH+cFSjOuWqOu2mf+8G55CxiKTbhO
FWYb8mvxcSEMQaoXbe/BIzcxREUa4eXyg9lnFbMxPNiVO7XUgtrCYnVup4Q/Cxi7
rTl5ldkThr2lIcmpaIp0wlo70YzfUFi608ddxJh44hvkO4rimuqN6dNCFyPV3pHx
Ns2GgK0POHsUBNmReKHmgHDFo+0LhpI8OIFRnc+9XgJZWC8GspDO9jHWusC6dGyx
LiGUODBHwa/gcfHaZ63DtnSHnW9T5a1+Q/HnrtOpNKIVzFXW8L/qN6WRgpdF7JlI
JYKJ9ZiXpN7cqP86JVjc/znKkZKSfwU7HjYrXmN6CLyIdWDzsjTHqdtO9Iwlovxz
TwBo6EQllqJYI19qiCY6WKSyCi9f866/Gsmdt5g9LuKXjDG2yiKF1qe3t+LtJHQF
sDN066IiYVyuhy+0e5Jc8g8wjQEAG0XUcdGwH1Lrjtkw+krR1Eqd78BmpLmIDUO4
VH3AWHeHqrRnTDmIR4hLRoxneydBhQwp89NMFkbImOyaoMZpArMrRQ+grbTRMCO2
+QclF+UTMij62KYkad6qKqFBu4HFHPcYGRj9iJiIUwPKxAP9axXqb3v0DzKHoIGO
5oqU3A0qhOO8LFPl27jZEtgGgz8Mwz08d1JW6v6ZIwPmAn/ZSdnldJoGAGntRfet
EfezoeA8Qa1+kvK7btsaJDKq1j2HSJlZPjj5s/W+zTIAtisJY5cOf0R/zthwBxx/
wiRZeq326ivwb+FngERIfBQPgyEq9MaD6sxDjjlMEMatTmXuWNPrbj8H1Vb/DhJD
ogVB6QaNCxTjaQDCqpmQrz2dzFXmpj11I9TT309D0cO97hZawREJ4cUROVqxOKfR
oleKwMQrvhHxQRngnqDfhUu5vmYStfNezpM32+4nR1fs3wOsyjGB2rfXXVSX4zdD
OCBYZaAggfhVQMVsGIG6fGPHsv2wJ0J0IGwxdVGvXSEtoHtAcj5XyirJRW57UgVa
QnEdjFrtmT0+VLXJRB7zpl6vQ8/xmYe5Cc7V81XnNe0DZJC3HvwgSHJz/kdvm/1c
oiSb7v+ONyJrREeN23BdZzxgHm62WHd+mUTEeL7bOVNDKl5KVONU2yBkdpiLua0y
vVHdYIoNBVnngYN0D+JpGwdAIA3dyposk4GeEyKW1Tn3FvieijwHoIFWhV31DtaJ
IAv5ULWdk1FpZyAfgN357OG0mxjIabcvyq5wwNu6tIP+tdmNmlqrNX4R1URByHAM
N4dIPt+58hATmihzC0kJZwSbG3tcpXVH51G2vqD9dRT2CmkEGnBzC6yxLnq4R1uu
rajdrKTtCYlDOWFggRQnnHzp43iwxWsff08/nWdN+5OaIhoRXZjf7za1bYpG5sZk
ERlNXfUOG8yUvwABunN7chihVwDYrZMSGx4PjVrT8JHTnAoZodVBD0qDOfb1WgBq
QoibxPN09E7v3pxYMOkVBy6VhNJhmKeajaXaKPCBbx89ZBffEW62ZH3vHaK0yMbl
HmPes7FuPOB0RPGn+6B2lVZO9jA48PXIeUveqV+pjfbidOHakMKBO6U2Gmr4U/ED
WHhpOMMOj4tRFThJ/vgAg6GGpPUeq88FxF+rsnazxjIXZncDF0iarp5UheS6mfOh
BrB0UiurTcK3G2VcU5ZRmmdsYMDyX4asSP9SxyPzK5Pg2p/pYOrkW5jaqMsT7lZe
xQJKbgEOf3v9gAi7yTgQvlcDakGyGL/SUyUVIBZZb4lv72JxxJ0taZHHkk9ToEaT
Uxg8n1zQ+Yj8Z2tNvGLKswk2/cJjG0wazr6yqCHGE0zyqFtcajIDLCqcM+C9TbsZ
iCns8AaddqtH+VftoNLmsIO/4jSGanltlBQOfvpt11qBVk9qeYX6cGnPchIwA/Yg
jTrV+0JD1tr/Y88bxH/HxMNtVa9CgudqfFCGqwTcbooin+lqNhHy7ynBQDqJX+7l
TRU/2HDe2TJNjGxfffqfJcEzPQ5HWOzQitckC4Q/Toq4q1iQ2ntsJPzX2iF8X9Fh
JYcQUqNabqlkGkARwLjo4Sv5SE/vZvh7zEPZ4W0unaUWe7AdNEi1XJBx4xfWpQZD
erwzRMwV1iRiJ8PCv074tDM/hSBoIHbxaN5i+ebopG1w3kTbbU1XJixKHuX7Lm4D
EkTQYOioVah9i6HfSJSveWovMsaN8jYBeE7FbbWgKSMOwaR0jW1xUQJNy6NSw0iO
H71ClHtfIxF/mP3N9q/TdRHtSIkivVSZ7BGfNll4H0od8feKyR0w2nzMGevsxupb
0VjCqbSnWXo7LV1PiJaHQAHSY3jdARc6na/LIf9oHQS8kUYJEaE0ozfcv6+LiVc1
hzOgYgu5ePGiYu5ySpKXb4U6snSzRBDZZ3lpc6AHMeW5/BPKjIPhliQlNr00twDF
yS7Nc3tk6gXYjQxYsuxNpdjvlSKKEQxOxQbqEDskKam/y6NkGB5Oasf8VCWeH5iH
5ktRjQjHOsGAqDo6dnTvqVMxqjNEz1xgLt5T4tTZ3RCMiGWKk4kBdpwvhk4WO9IK
B6X1SOlRqLG6zWCp99eUdBYr3sklgg+GhZqj8K+S6XxhuMXEKK4pINiwNZaXADXt
wUglMoaVs3LMgy/Fyl7+6MJ26tLYelPbL7GLrY4f1Ka7P0qzBIwh1KkoaC+DCJcp
m1ZAkR1Gp4OKllpCtGtnSll/Hfl1H17hEkDNCf8x7KcCks5rKvVXYGhQWmM1x0Rs
/vOAFmSVmtAfEDO796PIZHmwDaFovB+oImnxdeZ5fzyJL+Rue+XMoFf9kQ40pyjW
wZNSE0IhvbaPUtGN+pDQMPP7wEtCxaGW3pUmhm7H2KmqvzDzcn2+zhe8AZc0Q6eI
t7or+qdhuG9Xkru0ZVXulqMw16dc4k8af8vloCGkbRG5DGyc6rtNnQu4AWh6EUel
lPQjBV3mE4g9JgBSw32az23HFJNatMe6tpncp79zring0+UVIiOu3WQCP6Wfk/hW
2Ampv4Pg+3ZKRzODfQ6W0Den9+Pf/NRBjBd9HA+35/b0YfMMGp/ssd2ExZo60WQe
7BV7X8xLj2FoUKeeVACTYERCinuw5t8ZKlGkZdwt5bRxRbZ87RUCRBP1ec3vWnZc
223bLve9sIx146FsFO/yQvWSQNciXsSS5DyTuSpSnwdvjYusNOk2ccc2WEqE+S4A
e59R1LTKQz0YhDvsgoKhr/CLMG57cxc89NkRKs+U89V1fj7SHOomVPZIQtry37ZC
TuitpZ97QPs9ieG2F/n5y6amKyeKoosWGr8+cuduQkuYT/45X5ixB+fuEIsx3sFn
TNkKU4OixAse97XsIanxUrGMKYhxSYpVgm6XeWpl3w2UQ1pJR8pL0z755pFqvScL
ofCbUW5JqOPmJgtjxFLTtMHYSBNTyCMGBzQr4rdYoGunCMDoS7QODJ36CkB8fObN
92JbuDFBkikwcIAODQejtJEN6srBDoyLg74Ggsgd5hhk2lcZ20rMqeQIkev9XsOg
GsmNt52CBoQflYTqQr5Wno4SF+nAIZkM9MwGBVecvZt98pLuOYqivD54zJqtC0kM
uiRLmr5eIVxOZY1Mt03hzF/kraYPKPnY7/cKEXJXWnJpfwQ3S9yxN6f9CrkhPNbR
vm75ebtx38OGt+GaVl/XuELtZFdpfYpD0MErunaUjZ5j9LGEu0EObNlRjZaZfBHb
EIp7qlDZh5u0gD9Oo/352ZMw8tbrs349hpMM3VwrJs4MezKLgaGNnKGCqIkxBJ9e
uD742Fit1LW151oo/k2GcYwx8NHZayFFGVvjpMCY4Ntf//g0eSiCLaTZ97tubroR
5U2DST+Zebx86c2Q9NGPUUnHbkfQLAUJiljUcUyNljGJWBamSDJoFqZygBeUUXyo
Q2jHSl6C+hod0DIMc+XIba1HRJBDyDX9l3mhwsi4nTcQJiSo82990KNTQLo7tgb8
MEKlQC9i/clMRn1C3EympLPTYeiItagMj50yoD9hbDr0kbbnuG1V2/grm3vPBoQ1
BlSHbn+W5NeLces7khOBpvbZsxdXwM8rlGE6zpNereQ7Z6zJdJ7v95b33uAufHwC
8XNIW63PwLphrXfkvV9K7DqxPgoV0aDoRWQiXPBU1tZvL+1LHbEttuCE8Mh375/j
bazUZdjHaSyKSQs1mFOeu6FwFLIwTUNJ2nBzI8nS1mKf8krDVFSM6phZcG9cA9Yk
F9XDFk0xem1F7Vc1eJrwBDm0yekV73/3/kff85/Y2SgQM55io5V85AKm985VS19v
CEsHsxqhPJ0pOvu7AmzdhoaLSsjuhESxHXaFXSEzRlcPc53XqmhM961M5BXcsHog
VVM1/IDhDBiwJk3hrtCCerRYUkxPOb6pLaO8siZLAtCeOqffSd8g60/v40t6oLdb
ENr4zAlsJ0uYshzgptmlw/SkqZCpc+yg4Ce6iXOmEdly/AK2oZDR5NJpip4Nt/qo
BOdmfu9ItxkxQU+LovmgQZAS5VIX79k9ZSdgQmFsHzal7pqW54tOhDFCzxzaI2mT
H06x2yo2ovB8vckgdmMO1LmPl9/WQCafQLOHYwpjW7ZCtExiZF8Yuso41trgx5wG
EmKFLCpxQyCkgHetKCdAoKHMlAOkcgbR3RhH3VuspNhWBFdKFh0xPeQYKcuZ8RQY
pnraEhncjairKIu1BJhA6fftUmTKUHBrCxOFK0+ObHef7SMKV3fMKHk4NXIIBjdk
g3XFnwR7M37J+4qDB5zrEABuNoNLC8Wnol8lLrKWEC3qn+WaUKZytY0021qpj/Dh
95gHcQXuepV1UuZjoI7HkiNISKNhFHE5Xt3WAHLIM650zWfvMAw6ERneWBKsx1xu
trTJo9C1wH9vTT3dgsj+Y9uIfX3vKWpV1hB6UMzfirUsy1vJ0aqCjIgKpqg8WxJS
N/dSuSxQdVxfQgAd2AixpnmrxFVZ4FplhwX0nDahQ4q9q4OBwGynIBOwLkllwNcF
FCrreJ3XI09A/5HKbXzyJOQTtaR5dOF9M7sXjMMc75sCIBy2pKMezeFOz8WVAvEy
m928e8VXPsyfFQqJPwkXSOD8wgGUylaqauT3LnEV5CFrIZRq+4dV1GCMV/imnvgY
gjb/uAmM+p+qtyTsyPC8wAjwDxJg76792HbJn0ZJXnpcO2gSnpAf19ZHc0LPa3p9
ZjQ9gkNbc+yfVc1x+ggElTWccmUmKbe9b4TERQfdzLeSdXcncPmwRe28eaPNRtun
2TYFSY49Lh4G9GbkI0P6G8ODTFcijTQfiORBrlQCG01qJw2fKMb+TLSieqhextDo
Mmj9dtrrUYWWAY+ecRfdZwZCw+g29Z208OxGIADYC71a9NQdbEVL1mRdXIZCULh5
GZqpbim4YZYszlNDnI81NzmSqRnscPCg7mYGlrqlopwDso73vBl8Sm6yU5rlpu1Y
e9dGEPOl+anIyq4HHmgCJc/9P+PE35br6xMXWSxq4IZc4OWu6fqzlFcEhitA8V/y
MrlitB3zj6vKcVHKJaufFhI1IQ0UwOYFbWh7GmppYXqJaRopaGQJX821sjIbCjHh
aic3czVpRUslnuv2sAIHjk19YOyrpBpJEGL1ugYwhkZsjor/JxCmL8bIumHN5umh
8qOY1x8xTikZconJ7rgTmPaQYdLfLwBJW/+QoHULg1dEBCxB1Z94wM3L9B30THa8
HGI6Q7Ww5a5NTKCHeiRQOtcRbq8TGAqaJKAWfWGD6CzgEYq5d2dYJ8zZByS6IWnY
zIHY/IOhNi797VSvDJxgvuuZ51b0HiSe8gIG85HZddH36RF8ugig8gAwZLdzZfG7
wO1pJ+MxeOJPkZQX92Plr+UvJVvxdKaXLMcWZxqzY3t1lgME+0h17OJs98gfh3sc
kiSWFF6k3t/tM+ptvK4t1rL5OA7ee+dZsxHC49GFQg4qXXhoRLWRqyVLLz5RbjYp
jf1eWDD76Sp53LWH8qvnPH0XptvKFLJpq4Jqfbu4eVaYUhaAkHItiFaE9M+Sa0wB
aR9TWDmz2gP6AYezhnLnZt/RcZ3BnaSH4R5hQ2pILgc+8ONYTVKfMRO2FOGE/od7
XbvXJL2X6NiKF32Hr5qPQY09H4+5+u5eDD7qB9+dkYyqWdIqAIPmDiCLHcIMP1yF
3TFeBPux6tWukvrHQ76O9+hnJuU09Aqbub1+sJUcsxDXHL3QNRQdHZHFAw7KdA5T
83le/d6DDI6YQ+43xzy28BP9umECjMVOXudAk3KgI6jCLna7VHPrgYWtZGLaEPhb
wDtCSiqr8zb6jv1hxYg5SCiBO8xhgTRnG9oj1Q7N4MIiMtJXLFtFhdlKf4Ah8HF6
5GicCpulM81jOyy11NhT0KBfj5by60Z1IpMTHUzDsXbb1sWQO5wQQiQOODkBky/P
NxqILCiwXI9JKAaZBzNznefWkXn7qWGlR6FQ7MKedteXidcPPgnDG/WgBD6vfEv7
sOPWigtrr/0fYWlJrCCuXHa5DbpzcJGzH/mf551nKubdgDDe9FOQKaiTmrQz0Mi1
tN8LfId7PxopuMlfKqZFDXmn3mwNHU5BVHk72wlFa7UywdJPuSjWANUeobM4xv0I
iRbIKgdowv8+exdwA3udSPvnsEQlyfeF8BDS5UltjfML5tRvSa7c1KCTjIkzEJfc
kReY0K1MS1FY78Lpepofu7+m6G9ARvE8EqLHYBag4UBoFHIkpOk+JO1W1tVOUrpk
1gZCGhWVpi6s5d2OmL+zo4oXwz3XYMPcfChisdSb7lH9DJbhdkf1jlfbwvBwl3gR
QwMGrTO4fn9MOsSInO0R49Ny3UYVmXV/4uovNUPvEsiEpkr3yy10idtwr2uW5VFN
Wa7jh+cSiaSWg/2kfqBQVLHfbkvPf5NpioodPUva1fv2A15pxM9jEEEdyi9BZv+v
JBGLEgrFSXWGrEkPHF12RiSsBde8dO10lY/UZy2DvEkG5z8ZXI/36LESd8h2wkv9
KBzDNahIaqXR/6awVBzFDFJezcU2rUIb0oZM0grGjwRlJJ0+bcK4bT3v9IZ5ZzRJ
lyxE7amvmDlT1gys84sqsrNo9sCtwWW/nV7W7poaoueYO2WU7VbPyeQ4AHiro9i/
dxK37EjBcSA5IhZAdZfWtqj/ebdCKjDSN2U+eojxnB0R+Xza/DvNqGnc8YZLl/vQ
YO9YPhL/fWkNMn+zT6T+ADn+qPlb6qH4tSG43gyW7QlxseS2MOLRyZ6sKqUsCP8K
HciWofkQMuGDFy5TkWpI6xYoF7tgbSEMhSUgf3xkU5flj60sgzpMnxBvecroJGsV
suzEXPq4b89KzogqR17eQOMf0bZ84lQWm4x+qOMx/KrjIY8WGeA5BqDbJRQKQ6ao
gl7S1IS+VePCMcgKiUdnYzTJo2n0qWmKgM3LKBDExXrQt0/wj/btL3Cbqv0I09Ww
UWlMsjqlrm+Rr7j+J+jKY7PVkz9OwzNWrDqEJnNwyC3aDajiuc97wusGmyiZR9Kw
EyFf2KJ9Pgex5gn8fGgyYTfB94+NWNksgvKyLKPCDo3+GnCY4yHsCwkDof4jOrvQ
kk5gHidEB+Hh1ZM8zuRmQe+TWTqeSRGJu89ZWrLfcYsICYiO/KWN6p/lfJ2EoiPV
qrFOQkhxOjg2ZzKmwr0VDf+08em6yia2Q4FVVFR1lBt8UYtY9RdOx+H9qD1WYWWG
OnKpXpc8HZD/ZFk+EJ01MPNMwmNHORhz4TQ51BmHs7o+U46sKeXMpdCxAM0YYPE6
4WUUtsqj2wag0bJjZVlKH1smDQm9slV4ohukDj2mZ8IqUQ/a5DF8BBGwVahZmGRv
6RCEqOmnK90/1TsWGK3zuoodimo8xTItblg1/ygddZFypaIOsUo+TRZMW62lw09b
BN5apOoRpSCnM5jJoq65q4pD8itDYStjD9rjM9fqaEE5jmsxgBDhIBUHlWxUW/kS
quPyH6D+O67KbYxS/9JElA5FaNmXsxrmFig1erRu+mWn5PvxqoQvRs5jrRYnzzpE
D5WxjH26hjcIn7l1w8lHH4H/1jCNx9VzlNVsUmqHYF6ioXg1O7sVU0yp1Q6JL7fp
33QGNLDqiYK1opg2Bg5507mBPxNcZKaUwyMsS81jRN1WQ5ILEOEGqXtdYjor++qH
RmhQU+HgA9glS4FiFg1JOlAE2wDqzQcLCbO7hf9puRoIvHMqNeOLDWkM8VB7EyZS
ezksiFF1v/RDccjBt5YppA/kb9laygoZJngapMeKlCd1M1/pL2ul5oabFeIL9VlQ
/3HaagEJyJjbiPieRG81fDl+3Z8NFnfGIfqNTBJPz1eKB/G1IiHbOEqqZWWgIE6d
9iTH9QhtCS9OHfpvLSTf6kDUTI8LdUDqGwizxJElFDbtxWsDFHJ6miOBQgwAYLMX
aILkSUS36oep4WsDNIc3e25DvaBN2CmybFHkIDm4A8xvMV0ASXnyHWG8dwhki6H6
IEWrq/thbTWMuWZN4kCpFfXm0x515THJMbV+bEB9bjwW/j6HMtKYqbltLUbDAisC
HywAp+Ix2Kv31C/bjBbKvRToJrhS+MdkMfoiTQoImaTe9jDwX7SwVg9fS1RrigHX
SUZgeW2T2Gpij3c7OX9Ay4Z0Kp0g3lXMng3YC3v2FB/gtVZmXmyOugRkgtV4TBDJ
mx+eg9nhXWnerKUw1FKE6yAY77aK8/j8Q4A5X2Vek6G/8QH+vN4w5vBHlSLC4OWm
vCZfVwjUsMNommv2B+j8s6b0ewx5fKrNKDZnPTyC2qVZ+PV/4DZjeu2/RS0U/SZ7
lJyEgaeeHoqNBT4Z7Vf3xXhSpbw+ht+6HsFfVYTVoA0/mNMcI9yzxV3YU3HaYzc6
GjxgA6+PsamMkuGEYAp72FZMuh3XpGN57Wqr7z3mqYT3yIDHn7JhTlR63SR6FEbU
MVsCZHuadDaWt4bPvDTz69u2KHyeMrO6QI027ha9tw8SK9GRFTBbYgG9ePypVf8z
B23JwY0hd6N0vB+sV2J/9By8S8wXLHNHwfpPX4Lm+BkpiD3sdVkCjQqpev+BY07c
vmj7ViJMMA/2w9dctLRa4ao+or81fctby5MCzZ5AHiaABTwK1/8vS4tIMijxq2gW
BMGa2wzqjBcTLNaZcYK1BRfWmn1UpdIUpmtp/0eKTLPf18ypyYbc5CE5Mxn76/ki
aFi8Dd7BV74h6IzqsqEP/+ZtYwJjctOdgeY9Hr8BrhCkcVEzyQh4DVSUB+6g5jA1
UP5IjgzT/usWMMymEknmOvFDM3k75NaPDtoJ4Zw9TF8tlsq6NnJjqrKhK+gK+TV8
vvc36OLRMKN4Im9CCRsduK8xOO2OJZMQ+E3EhxXf4+LQN8EyIfft2842q1EK7RJ1
npu47n7YIS81owBUlmUfdm+I6h4HRNFUu3RB2HBqvgN1TkRdHfYhoB5DfmYsauz+
8TLGi7vLwFRA5e0/v+vLrapzyNzF2yZGMOuVqB3i/SKjBhf4tMP/uQTj1sTvrvBS
l5SZUHVib52Jr1LdLQfITLqs/9dTKvoh1g+jCyZtYQFXhMcbIDGfk2NFQa5/5KYo
UyfIEhc7UIT7wUF5vazzb6X3ZojNqfJvTB5KtJjNrslGkaJ70+DrwsPPdXimKgUu
h9nw5GxqtY04jJyisI5y/Hw6EgoClx93hOkeGFb4sGIR5PfNDWNIhi0C2jPdtgDJ
02MFkZtQSaKjE7NucoHbtU6gZOOpMt2IhBKGu12rW+jtUxxe0ENWHcZrlaCKYJAG
NUWrRYH0s8ic1tqWa4Xeej53dn8eNTvMxMCZFH5mz8eLgfogztVPAJtkWmEH8pUu
TG49Q7QmsINfuI3Jjj7q+3WBS122Z1xQYbXzI5qS9Zj9DOQK3xupGyj4czetZedZ
DG53rZo0pu1Z6T9yuELBNGw9nZTj5fo5Ki9dM8q4kctKMYCA4/9tgvtJIrRrXHhR
8fBfLHJPNZetbRJEj7P/BQEOAfqcxmIvXF5/ECkwBSGila1sn2cG+ZwKn8FtKyNZ
MH/WTj0wFhjVSOhIDYv6+KSbS4cYdq/2K5jGqua6CwOMLZqWozkOyk6WsDhCMC31
6hSsean2cOW2sjgwvD4w1YkquKAwRzfAXoAyexTzGkLHGmSDD++iNfO68Q77Rw8b
o1M73su9K1V4yqXePPv2q2arJzlfUuB8Iagac4L19y/hNqQYIqKEU0p4eZOilVMk
0nsj+XAvRCU+J7o4XRhS8Xvs52BIIF+Ocelh8y/GPvIg9qEXta5J/hjVPs0GY4KK
LxfvwYGxDF/wruNs0LwFMlLJhwDwGlWXKmVXV9DL+Pb+8fp5dnkLIbmjmHTUvbm/
1zDRqmZG0uPM13G27IYCS3Vi+5LuG6YWDnI3SEGhFlz2XxZjd0/HA/vCg99y+KGG
IoPc0nzWU/YzVaEXNZeq3gSPJVhAteo+teQFf0bwXiffkQqeIIo8CVrNEhuSegzf
iND8TebS90ZXy2daeCaJKuCqRm+lmtLOsSfMJL6JNnZzdJCQA/FYHQL8TXPKJlcW
7EEEr4hfsIV1kaakqRA6JuM+dGdjyU8/G73i9q/JoTtEFWX7I8UU2BhbQ38zAwks
RX3eS2jcVit16NgewzMXzX4pn6jJFMONxPS7RUC4E3HP1q8D0E9z+RN5CSHUYQny
OHabX0i1ypDd09kF8TcvjD0DQKuYSsbXviLZLjQg+z2sV8XGklFKD/WFk7bhigQH
of7zKSV5IqCLSreyWNxVNM34glE0Hvf3OwCslUryi3Q8b4geWxzpN4DWWW5gPZGG
PZyXlN/k87inUBw8087Y3F5cN/WKhhwuuSpAwKR3UnJ4cF37qWV2q01ts49Z9zND
Tgt2PWmu1pSqmV60arkPYgCbC70yYEcJSF+4dLMVq0z7hLK3hxrEDMrN5/RcO4bC
BUg+mz91BaFtKxMMM4Uu4DTTNhJidsbHo6xZUCgWxe1zip8wmIjKI1glwEmyb7ST
B8ErgX3Hye6SYiv9q6OCV0OWQ6nIurBFb7zuWxMZ9cX9PRjjCXRFjaHae4V1Rd+j
5Rj35wFUDoNMqnD28YQyYYQqXcWzjUJGMmrVMdoxtPLW/FKmQ38wcejtXqoXoV3w
+346m1EyIYpGavn/xWtrNYfAMW8Hfh+CFkzNx2H96IlvQY0Y5Wnz/uxDmaEDa+Zr
/A9FhIBe47tvbgUBa9B26qhtevRydFEZvkPcn+ivaB60kqvWWKLN2qZwR3u5mj5A
xy7zXwsyyYrLy1VpRfvxrs5I8kBue2hsrTv3QJeX8WWIBkqjSqcFr03O2Qfnpvlz
EG++gjKlMd6tSTlWBBRyqskMgF70XTLVNYCU8c2JNBcocEKtEQErj+rEXlnq9tK2
3+HZagqhvlcY06kLGvX4hk8Pgrp4f67lasXH1FsOLeusc6LjlfjgeEb+n/gJUSMM
oNY/cBd8DaHdYdP+oG5/o7EBBxOv8n2l3Xn5QLgSd4iQ5QrX2Efhw3WLOItO/SjK
n0p5aU7lhSwby/vWuieV7LjC8XMRog3WPDt5kuS+m1lcVs/eiQ2IDJpIwIAn3gMj
rv9sIw+nbnkKHP8uFKrRVBk79cSLBWxaESeFCiXaWogrF9EB4sEnpItiCgHuS08T
L+6y60v4t4oZ/sbkQpoLaxO/6TkA3Ga7pSertkbmaGotj28AoqVk+Vv5D4AnpSFN
4xhIPU7FilJFTKluzEjSuChJy6RUp2Pg2jjJ219l7EJhjc2LKttKWCaeGXJN0WDL
I4ixp3ZNkhcZ3ddnBKgYo0ne4TW0No/3Y1+MBVnPurki8n2s/HIot3BdmFAyh4GX
OMlczrvN9iuQfB+A3nG3xFVn56VASQ+ZjblTWw7+ewEAWkqsT8h0/qfH9VkarfJx
PYuvHURSLUesogD9Gl7I4+o00TVp6I5hU9zaUo/pk2HvmqauYWZFsdi/amaWjHfI
TxZ6eO6Lkk3/LDFMq8DQ/6hX6eCUufdRrYYIYYFKm2VnbzafZxC+4zb/4bqpg7m7
kNnLcZReXUSbt+//rQyDzSrObGUpVj/UBkr93faqWN/kBkPZIm2WuHKw9f9b7dOc
JUCOMRBsEx90lknK/5oLulziT0YIJdXd2s23mCtLiJXZv+TdObqkIjQRSq4gTQmH
MzVd6ARyt8q4rnvyB8vxTQep0pkr9L/IKaX3UZsy/fn3RQYn+bdb7NL2F126kiTz
AaD6EvjjjTWksfFWcD2ITyNNfrmE9HZB4E80ddcYYMlXVDQB3GJeYRwkwPbC4fhg
34kH94iqxOl+kkFqr9PRlN86ILLkgT6CmQau7aR8IBrf+1zNNAkmV9IJLvZO68bn
LzbXtdhvXOj0YB/LlpFGAqcdqT3ZK7psSi2JIl4gUIGJaFjbPbWiBedHKPBzKocS
+Nj0h7fgS8LN/89SSyBsiW0OPSh78Rtv3LynNK4bFx4wNncfNjmTiAmCHJ9wOLtk
5/6iblzks7x/Qmc7nSInf0SugaK6CZW7jyGwHuJDxPa6QPfhjzWIqHCZhLThC8v3
uBnVHkBKmqebOxt3RdFD6J2SsU3snUMl6r9X/U0Y9PdZWTIPlfFEak1+IZuzwsD+
NEPqeNoUiAfUenuP6LTJVYmTdgKeZkN+6WQoa2EwCW5BESrQVmkw2rhrf8ma+FJb
amFQ+g6v2ViGx9w1IkOYdB1sxFk4JW0E0vfV6o4fGzsobPFCQ8PJSM05b0Gd6246
wqFUWytAQz/Ts2yD+9Dwn7OMsVLwjOvNg+MW4FD8cmy/yeP7BfC7rqvZyNeXm+KY
lyLeWeD/OwXj6Hn3HW+McmVLTp9uoA6f4UsZ9EPF2xr0+6qv/eIWkPyGhWuTZX8y
++oSrX4dS1sAirbNZcQZdhV1l/1aGP2PyM3ZB7jsywULJXkB6nPlyUNEki3JEz9B
UUAoQtAS2XVIoGUjaJtYxOklQF/c7LskkV38oaSyD7BBEEk6FsDL3Om64PT6q/DP
1MHubxLh2KeLz1H0zkBJ2ilSen+vHX+6sunfD5HSmLQxAmZ5BoHqLRq5SN2Vq4X8
SUEJ8PnidCYnzGZWcwJo9rp6gA1Z2VHD/0dpnnpPv4yxILhi0LLa9sYa0tXgxg5Z
n45ZPXdxQJXKrtk2HmasFc6wAUKWeaWJ06WP+tV4AfSC8Qjf92ahsOpGQq2Pvba6
5sL6XmYCEFd9NGwNkxy+jM8t5GT7fPuuf0dPodi367vsDkLVxQACIFDRBPH2xW2X
JbHUrzn3N50n2r3aqUfQtc+ukWxlHqDhrZI7fSGet2uF/Tru+KbDX0wv9r/ZM128
tLwUTMLlKaD1Mu0ilfpmOSYYKB+lxRibju8jQdSHHvaieWLddkFQv0Q/8nfl978H
OyXoBCUv/ejanxCvM2Il18l9R/AL4QtnMAM/78XtWwEoR6DdAKX7iHXOypswsM5M
R0CInMAc7wVgyjQAq/vvQ3djmUZ67Xeh2LXaH6/KreVtRvJGSR07+B6vhLDtqpGX
I8/X2Ws0wkD60gflOo/7OPSfRRdVYHIR9zjUZ/vqsSsT0I3l0wgiRaRj18EtwFRg
UaB7AB+N6td0JglHyvSLwbLdANhN3W0sFrVJVfQ79wMc+c5hol6xeGmnlpziQ6or
VXRlI/Cwys1gHGSzNDcD4QkVWvWyknhwXwzlABzT5YJdQlFP6sM02cGpo7e7SZtY
07quqbE6w3DGC+o0/eluu/6m4bt9Pths2PpOA05/DJHfsTCEylYIC9a872Izg4+c
pAH/kmBQwpluar2lRJCZc9QjKMYjUzdwbZxmnuVmlBGWG3B2tA+4BzzBtGIs8LS+
iHFlqPfGUk4LlLkU+GBZbZ1qw2PLLX60y9nYAP0lkSatD8RQSw0t0hukYNCD2cTF
vMLP+4hVZ1t5HAwQcbWf2uCq+UJUJKJJ0TlYcRHiKpe/p84iGZ6Hx47WWTlZJLQM
Q38fMPYRVDc5BmBWV/K43hoJrL/mJjE2f1Ypg1dEPZx+z6jNdGBSw1/T8CE9vxA0
ymXaAEQk26HnIEFqka9t9FUMuJCoq1tDxWoqA5raXsOx8s8SQfjCQBcUKBaIaSmi
Ske5azeG6+yypjQe3dm8pbMf229p4tx4jRHKq5Do1ITUHvOjXNeCIoj7MmaljhZN
VMNsgrTwvDZi2c83ONwL43xl8L/nA+ATy1vy0uFJctR7CXi9Jt1Et4XXYPKxeENV
6cp4WHd16ThO2n0P98MN8jCFYZIW/IwHdLA4N39A0pZ22bG0PFQjT78wrL1YMmrU
dGIRDgpHakRtu2JIyJ7k8lCxssad8L4JBtFYYRyn2WJfoIh3fWC9LXJZAkn+q+qr
xPEar7a6/mR6ycYExT1unDAh7KwccG7mVJeJEiKHHi31UGiJ6OwB/qt/91/IXKCb
hu/m8ke3DTZXrEeR60TkukEmmxpQVksv7lVT6v5gxzxvSn+Ux+BTPrIAO0BYaVPH
Rxorr3nUkew0BSwFVPbuOdlX3EVbJAy7BlK5ehEc3QGe3AWHLi00sMhC77uJrXwu
RpTE3n0/yUsxUDTpfDsThVSEpkYlLal0HaueYMbYA+eU6R7jh/3qOOv5SN4NQJ0V
voX1Aje6Q4mdkPKQOiEvhEMfmKvVWjz+A76qSfSLMpV26KAVn3/2QLnvzZ1nzi3o
SzNHFHVUfyF5upyq8cfILR+gp1QrYY2xW/cf9Fd1uZ75wljv6n+b0A/alt2hJJdY
6uSPXiw4A/Kvebh/A/I9e8GPLwxiNC9eZa4bNNhnbCU3Bq0ZPRoizgFgpR+fGUAT
JOcyXMVnc19EfNI8bRJlJxgiVgMa9Q1Pg64mmRase/CY6AKRmUzxSJsi5YM1JVn3
dpVPEQtsp6Kho/m4Wslo3PDXqGndt2GqzxQ6Ga0Wb2YIa/8F2q4qsmMGOyrmSm97
4KF39oA/dzoZH0uSf9760T54itBQjD/wOYdtvjknHlGUHY37mCRxfu4fWjBQVDSa
Av763xBbCOFfkqMbRssTUBswJo0sogEwDYka7Jk3fx/wZKpLHsHmS6AzqXh6AVnR
A2MRtfkZ1i4JszU216SqtwCcz4nfJyIrlNFXgco5066Iullt/Fn40IlmOVN5N+pu
kW/4nfsXSlDPmjuvBDx159RTpAE6ONaIF7cHxclXXLumGouyX57bu7FmTJ6oZY5H
S+H9v8Ul7pQRygOtIvbTqjbEci6L772jmDPFsLcDThfXbHnGpOAb55VTQ5HYFlDA
ES5S5+hFIR8g4ABhvDDz13ApsKCaAQeQzqFiE0HJMMIiLB7M97q0MK69uI9JOiyt
jyfsajy81FdfZn28XhswcVmv2TKyr4JSQFeE2rByLNHy3Qj+zi6FxN+n4VXnTlNy
kvZu+YvRSM8z+ywU/g+XW9mW0g/4IIzUL9ZD/p2B2Pi89GNf66ERZROiIvjRvn2k
pndEXEHYaoqfk83/Z69/xaopFztlLt3C+nu0BQPWsW6ucdWrkg25oAE08xKwKlXi
RM2IMnfZnzkBCBobkFNT5prY3NX/vyH96For+Q5m+FK1byMYRgyunxXkzxhyTdfp
l7gKXwkIBdsluUjAk5xEK9R6ZCkxXA+thu+ezhhHZ06LYO4a+HNXTfrGMhc+79ly
AQADJFDQ62H8UrCaDYEA0aYQXjr40+honlcGCzLKnj/tsTfeN3ix2VSvl+D7dosF
oznyDjbPftY/c0I8+RudMTrnoMxYH+y2986HqXupZcoZmN+n+5uWIkzVxX+a/yEd
grjIsWIlwy4CyYEF9SF8d/Ae+ap6mPKggTcB6W6TRUsMXZNcr/jhMWEc+6T/rxWr
V3ZGUyrPYZ/WPDBdjhVGymu90LPwbDz7fssVG+c1TFjbeaRNydpwslflILn7pWSA
nl51gdDewbch9CoFdCoa7vtcm3PZ74Zwl4oQGc/4U3KOa+YCEhjxSGh4/AwWaQZL
f+Seo2e7F/ANKCzCa+j4m48X6eCSdY71rcOLV3sJOT6KwvhGVafb+OSegtJbvSrh
GbIJt7cDa/SK2PITB+fNWEzNWJFPfOsRtxy1mwolj+d9R9BA1URQ0oHkp1tDDeg6
va70n5qFQJtR49O1NxgQRgGfdlw780I9T1xQdUef0U/urdTBgySTc37S6Eu76nY8
HWVSMxgxMDgbIiD+613GbEyK6Bv5S30HyCzxa1hSS/eqfN+7dukGoPYJ1J/v0KPc
hXJJMx0WSRQFFZmZHIaZQJKuCo88BK1YtxNKACOAApibw3d8oE43HuZrw9C74MSD
8M2UwDB/V7hQCPS3PWV6WNgyKN0WwpzTuj+U3AdjaZ5xCvXhP+foKYxqB0PIx9Ip
PEEjbcWJiNYGwXAsdRz/FvFzWs59fZnf/50q8fkLZPeh2hznqopk9ZjLY/wAw95v
5Prb5u5lfrvYN35PBWwcVU3fdrRdSCzO6EYMzSDW+ngofGEyCBoRInPMkiN75wVl
QwRrOrcdH11UUGFQjq2Uobs+YQrwEJjTcUZmcl1DJawTH6hUWFLSSM3enAGeKhPA
/j37h4Y3zGbuxW1Wsfs0RhPQ3qJZ1rkS23/LT0ytDXnm0ziNX7W3/kxNzqJK/W3P
msHKvFnJuV4a29wyCUoMVCFEZEQVCVgA66qgZXO7C1zmJ9YMm/sDff6CS0UoqH8V
YlPZgoU35ZK6K3Vn1T2SNfNCG6s6xAt7X/9M4vOQNWXIeYoHihk7EnzBENDPIsKp
6NlbczBJ0Tihft/HpA04O5ONiZjK+pzCDc/u0iAuvi3qWZ/veiIjKrW7Suy3ggPh
PfXSrqhGps39k8NFLxCCtOWYVyX2+98Y4o8LZubxn/61nyMc0oPaSZeILaATWTvg
QAdLSnCe5wl5IQudMeR9GOUDzLpFGPQWqcV0H50f5IxlS2ErF8iRuK4YqqVAdlX7
UZ0K00Yvuw/shLbdmHNdMJbKyA33Poidoe+0xuyD1/nF/trI4CbW2RCieVFgkEcW
qo7JSC8xU0wNiu3AV9JiOYUarXv112Qlz5ad2FMV7GnIYSZfqfHylTwSWCB+7XmW
x+rmXEZTqMrfBx047Uoj9lGaeKK5+Ag4jC9RHwt/uTyHve98XbYUst4k3qD0B3AT
csq6wK5Ep/Ls4HfrvHwTZsaNmIRCm4mHfZA3nMTjqcuZkmjvC4lMmVV+YIJE+yNV
fjS2ra+VRNsz4sNP9oF/EWHrhM+wUutLwY1htNgiADI66aJR5pProivk4k3Qz6jz
yqqGgB9FgCyaK3+WFi/TYhO4pqavCoJNrdInBaaJXEwfAYWo9rqMsORdkRINv55F
3p9prt9DWem2vm+R0A57bAtAg5f1HJ+BWawjzcvBE84oqfNeoCAIMnHr8TF/goyW
QjoLYm+u7TEQZy1ZjkLgdoRbml8oq4nbwVyZt0BAKMXlC6OjOig2YajhnBRqAuuo
Ty88NwyL1SZL2izt5Lt43SS3BgJu5t0DdeYDIoF6EgAVqAel2/E1OXxxs91wb+4G
l0Iwxo54Gv8BeFASPQsl1Qq9jd7vIHVMgtEzwvdhSS/6VqrdV45aTFMrkEG3ZMhQ
97nvckjUPamMAF3GvWCQVyPDuRyT0sNIsN2WuFuVw26XBoJJKOw3Og5vkpig/BSD
lpyQSz4T0VGRq28CYI4jvBBoBtKuTnI+4uYI7pe5pE9XpduMoFUmOl5wLoNucVLC
+UZMIyU6s43vE7y5af57ES+scYjiwAxdoLNDrW0RHk+fSUZ08NOcU0eECBNCT3VQ
lkjFfPvwxIgfPXV4lDeOmiWIB2TyhpJFgwDaxuHi0GTIvqkHbVmXZlB0wFeBSzaD
G9tmUTqU7nnDQBWbDW3zn0K21zZMglEMpadm9SUKmJvmmXFYy/6isSYRJpaiwU4a
riii7V/h48ZTQ5r0+s0tBVKplJY1WhrSy8Vcpf7ByGqWdx9/sKum1DqR8wR4XliA
A6beXBKMK8MNzJ8B8jzMxnuqs0M6A/yFBHCBhnRuhiPhsJBoMnlILS7U0+aYTdIM
3y+T2YVHFUOBzMygEKlFpHI2c+xtWBTJABVwkIizzJCHVW3UT9O6Oh8wGYE+H7HP
sDEyrgCLwxvVI5ATcyLFebXqQY2kOCkp58RRia5JIfOIAT1N730RbPKS12ZPPfV8
nm9Ot5BCx4WJ0gVdjoMb6CxZ5PjWn3GSRMcmT27UPRw9VZv99tBM0+7P+BPyy5o5
P9TuQ3VPFhFSAi6fOxEf+m7tsSn8eNiNQHKnoB7ElqAWoGxVWJGYYnDXPVAMVq3T
MnuZCEaoZuVUDJhZGZg+OqlIAi4hhZhmQtEvC2E/H/Epby59tFclpsWcsosBA9JZ
5JP957a2IqzooJKwIS2YuiuzqSIsfwxvUYcKB7Tk+L72UZDmcqheG5yQ6Kjdml+1
kcSmpkLUzHsWgrM35GhZV7P3EVq1rwdwSHvBp21faso3GhwLdb2Ba4XzWIYRL741
QZhJNagOIenVYWsWvR5SY/MN/Ls5vQhPBV/ysMxMYWDALucnK/UuZSdp1NCaQr23
l5T0n02jlw2UaOTMGGppSkNfU63YhbPFiAwBDr+HZMq99aN5qOj6WaJ1NhyQO58z
tD27yyiJIC6tdqG8rOMt17pBR4Yg9e8oMXZO/2TkPrcArsiH6glzI18Q/wZzlGFB
yPCA5pNr6gS2cLc6AF0gTt58OHA3DlQIB/Jev4a/hQGfVVis2Jebwaqy7PATU+rm
Mq3Bn2ZY9Y0yIQ/EwfBc4aMp9iXQqR2uuRRvBIlKffeeKLa+h0kZlIBr//+3fUXH
KdDatOlMuzrVpT6EnktAkeWelC2PKqalLA+uYbjXVyoEpQWSX4meNz8AVbcJVono
M2RM+ekWv33MBzMfWEOS0faEidGIg5Wjyqyz3VPcsZ5AA1+7x3XhX+V0240R8QQz
cAeqJS/pWhzjKfOqwitQGO5YcG/8iu8bd/+vHvB7rh8bxccXt222lWxKId9NEZvQ
KINhxMbJfwRNiSMNsWC28i74skmr2KWCb/3Xb5mgTl1rqp7wehCvRaXCXaPebhMk
CLGNiWD2Qdf8BOnDXQBMAVRVXw55804r0bDO/zIyixoDuOkohTcMBiUu3ry2yE9u
2oNjS3hYvSSl9lZl2MZqdEUEkG49fGQbf2u+wO36LZyQTk5G51K3SIAyN5zlGgaC
YrbdyIZ08whNX8dG/n0JU+Ke3aItx2SNqAu/S4+uxt2j/ZxEvncOt0Xh83wyVyy5
yd9k2oNlSHir5r4gU2sXRURnLHIbFBcYshUQwxet9WGiaZSTSOduvUZK/xIxGNkD
pLe4yHRGaTaNIfTmWmFF9jTz+wYXIFhIFv9anNwT87Ls93pF10aunBN2MupBmobj
j/nCTfoGQ9Nd4vgiMKwpU23cuJzEu6qaCiq4XGygviqhAriNtDVFnoRn3UgZ6UX2
P2EaEa08r/e+zXEMbs6vxxuFlaWSkeTIpvNqxSxSYaUGJEaSZCV5W1/jiEALxRb+
oFVTxUqdkJWDU3BIrsa26YckMxvc/hXcPrN/KbeyNNDsunSGuw0NS5Ie+OEZu0On
dgygeQmpGk/J5nFHTciwbj1VwVxTFNEBrTGXkALindqprXXm7fpYw+M9RDKIXYoP
JZqZtjF5cWmppBq5NoGBvhmReAO+485KF14c3XDVq5UIm9vE0gf86SrLL2C6RXbN
eel7VCkgIHwBx50DOR6vWQk98yhqB2txuKWCP7ys5ZDPNNixrdXXoQ+HU1otXgQH
ryw/4vBYmuZdDGn6l9nwsUcM7E43nWGfi3FBDIqiLWAyYZHtQZ27mQ7aRVppQo3t
8RIZxF3H6qBbtGJlBECJCRCKMrt3ABpqr2UOckb+b6M1c+6+Aewm5onQjYCQY1WD
HuTV5NHJdwBxCS/f48hTJz5xK5AiojL/5uREy7NDZXIncLxpXb9D8G9/pFsr+fLj
eTtjR0U4Di12Boe2zt107ZwteNwqAmT9UaAzyA1/J/xKddwmPE+Gew/UvmABdi3w
pg9wIiXmLrCQmSnYzs0v5ihHmkbVmMJdLz0wjlgDUd9LjOZ6su1h0MuXzgd4CL5V
Lp7ysloDEAcGTmAYT4cYWlURdDHrOcKPDXzL82yx35+esNFqfS3C+ezCWywsOvlW
TfmSJxp14rYU/VkWn8L7WNMA0aIl/21+fRAMWn3PUtEYTd67Dtf5TOx3EIbxPWx5
XLQXsNXXj6mzGPV4B1GHlHhmqqgWa3cZjuQmLx23XGYTQ0Am++qTtJrrdo3DR+Dx
ltdP9UdJxRyS1rnUsnp6INRJpfscOKQfj8oy4jpCu+e6iFgHgYZs5lH2FUqywpNO
r/ofoG7tr94eqapujpW+1GtyAT8+3HwPrAeKrwIlLGuv6jkTz81Ag1iyzcQmd3Qb
oblmeGomTfpzWkwp3HeojB9qSsJw20Yg8GK4GCw9k1hzM7lUwmbecFmXw1jWQ16c
MysYarlkB8x2vl5atCI8IJv+45lef5GX+hOfr6m84xVVmjIRpfyhgVE7SJ86qNlg
hwB7JYKMybraIVti+p8Uzzvrk7+fdWRgtU7RsIdu0hnbt3QVebiHEZZZ/f4xp6yp
RniHtSSqdGOJL05wUiI+gpG8XQFne6yKCL1J/LCFvUS3lRkVyEFSgZoIv8Ts8oK+
M+fyw+jcs+k9k+9K8ER6IEtuaYcqPyTi4kNgo8uQat+2M2AS0sG1Q4NQVsi3XPy0
GITxzGYI7nvceOyDl0YhkQtOL+juOaY1lnZ9g7NkIbWK4FIdFvT8RHiOhJHnOTWm
/8KTNcaSAHMC27SsOkmwYtDsa7UG6xEVSKVrIoVUHcZGLakUELyzWMznttZy+r4T
/G7wiLRWYJo4vorjLW1/vOkZlwPLS1tsLURW8KgcvoytQKCtCLJLe/6kr2xAHVIW
V6Dn4+YXpIMpkgdNj7F0DcgTgsJ25zyrXV2SF63qPYkfHrE417EbCEzh60Yx8qjl
xdSLRWvNvjEzKA/TuoiS/TFSa1tJegPB9f5a/98Wo1wHOiZrO84X37ecsdlCG6iQ
uWhNUbv3Id5dE9XC7WTk5ccLcKRxCUFe7Fnr5vUIqO1MC4WY+2t23735LZM8RE3j
jY/SE7BDAGL44F9FWC3SQLMwQvpo+hwtt5/quM7vRvzZJjg4pfooJSBIq+0ejQ0O
+sLZXPOVY21CVTnS5QuNKAAqhkEDMsCyyirJOe0g/ndhVw25jKYb7a1mTRalHyy2
WrO4M+mZofcgKxeP7PPi4XVyUOf0A//sdzY9CvyjBRQBO02n286vtDFBYR9423k3
FI8tDcIjIWm5oNq98FLtGR/l5CCkk4R1IKddRUWsi2swJTpJ8gagEtAV8xR0c21F
GCiyzkxLV/u0SM/u7wVTrbYVp1u69w6cBiluERFRQ7dHD7gwdq0YK/8KjfYAY3D3
jj6o3YyUQ9uz1Myd2MzTR9bXZ1vslhCKecJ9Uhfinqn8f1P3gBfS72wW2zidwj6X
ja5zWLwTKpMi0BezWZLcGe60/IMnbO/d/+UbBBh9ZHRZi2ojNMiL9GbXGgkIdvfM
lTHQHh36fxrWc0QWCV2/nO5F6Bgeg/nrW4VSJ19lWcqOVQmmLy0MTv5nw5MqRifB
dL/zOjRbnS3s89fFcEZBCSNCRufcdwn3qxr2czyhjcTkXhlRcanut283jGpkFe0n
3iJxA9aKIbSv51rQxdhRLhJjMnoZR3mo3lCa5j707KQW2QqgMzzTsS8Gg6zvg0N4
ltAQHkX7PBAgwniyjoydxZSgT9jUSNT+ogb5dDfxb+/JsuzXHRAC3go99+5dlYJv
mMgEErwFTzTH/AEk4ae12xCpW/czgg7UZ3OAA+T+hMKeQUyMIpvNH3PsijYD4/Tg
GfKmeJAT3UoCfdIfEObDUjda8SrsGmyjgtxca1XamETTfoYMK1G1ndnf3Ib3RSo7
ZvdhBuoho9M8BAHfH2mwNZyIlwTwpG/H4ndDRrQYWCN+45VcPp480GcLbQfeYo6Z
FFBxplNpXBaRHI58YoFx1yoPP4nCcM0bqLKd8/MVX5Nz1NsHyxf77DRBwfsKJZV5
q4uQVJAQ4hY7agxLjSOXeT6FQWCu5cls6uWN4w6lgSccpi0wY3MAJQg50Ll+sHiP
K5hGKldqmMSCwmYk+Stw1G4SPuJXoycPNxZzW0/c/aUH1d/45p/YNFu/YsxW+D0N
NKrKDSLc5g5v4dywm++B517GFgfi7vp4P6gOrahgI/xRuH1Zycgu0TINyGPx7cpe
chSQ63XAT6gW62sCDhCw+fVba5BUtc56F3fymXhIQd6yxW34sDP01cv/dgIBeq20
yTZewItR7UKfntBYTT3qFC/3z3jVK1A/Ge2BV9YePj0BVbta4cOG+sEGbmLcFVgx
Z2vpLSPPfnf4sT6CM6f3ggHOeds5bA+rKQQJSg6pkvMWMCKpF541Mir6196e20tM
xaPJ1h57CcbxS3nKUZ6cVKvFAKEDjvrIhE4/cSqnjf+9b/80Rr67em/FHFcb7D4B
Juz8/Y1NE7KDxd3KNffhpm/HV3/w77T7t77Mgc2fdO1dM79P381PviJHQ9xDrnpq
6pOITW8CnpqRdtn0b4VMy3OtxZ+cg+f+cyZOwTulr8mHfAXh0r6akkIJZllSPCln
99h3BSy88eC053lydL43dkCzKhK0BOSBv7FF7A5zZg5uLqv/vzAZdhEyXNOV/Xkf
Ce+/8nnq1tngMC7SWCmRDfeYzJ0C8HW1KgOGE4UEonro3HLB47m97uWbicd51N5x
6fOsxzumQiX1OMbhSUKv1JQ1OFdoaSMr6NtlvuO4+STv8pfxnGoS87pRkB9TBCmQ
5gPJbcjaF8IijGNIS2JCPiZHpsy43X+jaeRkQhRRMrQca1E9jrUMeI7pDgfa0BBV
Y062OVHIxvprxkfLmK5oCh73oNmaznw3Lw/asCNjTbYp1te2MLq4eH+Io3rv1b16
3DqJemSf8Js+I3k6X6f5lhm+FZvCXZ3l3T38Y9YDlHr/2fNpOSinO0bW9cgjMCHL
pYqGIljl6+dnHEMXPL/Tm8jMQ3Ri8rpeJQbAUvBkMlNAEULOBf1dd2iaiXsKBJiF
E0d5KzlwFnBlYYyR3D43fSsaOcbPzu7j8ajECkF6dw3YBpgNa8qdNE2Mwu/p/myV
rbuNj1o3PWz50FT71bcIys2M9aFIIl3ulBnGGaFuPwqwqXEdhr6M8K4P8fLoALvF
lCTsWRWkji8sITx9QDy7AhnpE44N0n4kmjfSI4JuL7gruD5T7eu9WzF23oDPiXsJ
NGs8zqZg3Wo56tIYwYU7o0K7uhhILVSh8Txpiv9ehy8dx3LJPC94lCUhcdPsgUdV
G4bLqvzJdzEtWVRRakwSiNWsPgE3lY3uejcV4JcnNlUiEpcsSeQGqkVJz+kMNVD2
eXoruwgBQTWehcKpjts0nhwhO8XTncmF5sXXeUe+/+GioigiiNehlXvaq1lC6YgI
KiuDWYkAFXUuTuSQAgelRfQ2JIDiprmooa6HmKzLPM3CImPG4TCXaxer3u+pVgJp
cbJBdkvbEEnwvGIYfSWYehjcjFAXXENqHrgnPSFEHMKWvw3ZaiVyMhnj/AGF08ni
svoIvq5VO03uzV3KZK0y4LT5c3mzJiqaf0KHbPCv53Cev5dcYInPtkl1rtV17oOM
NrE7zbIi3cAwv9sZq16FfHPsVT1763DQx8RTVc1x+85Tt0Bt73Nux5CPsYC3TMFi
7JLcW72SbS5ePzpSBH6gJYSCyrz4CIW0YxSn+pfWV+SSzyuIGzzkx8kRUHCGPezp
ilrL9/0XptarF1Tx8EXavhCZK82kgJuEKb42RKdZR3OKQ9VNp5MAJjKFJbOEIxDa
9CiUBJvmWwL0JPadoNKdCAFEEspjeiJnlv7Ncy2FLQwiMF2zFWw01mk/Pys8z3OJ
YACaWeSoisB0IyIL7QGqGl8a3qdoyt1zI6xKtn66BIZ07KW9fe/LI/nn7HsEyDsU
BQptj3VwMXKbQYMm+P1B807OHMASjE294/JQZ/4wG7dMtfgLTrS8Z43KiP6Z8m0d
owJw4Mbjy9ldkMiGe/+HR6xuAlA2pAgFeyPR79bm50KPM21+OR8DQfLtlSsYOf/o
KyyeyiL+INhC1MUc5ahgDz84JRc/RTUymNkz01xqCM74NlJs5sC53IdIAh2wWO8L
jaLjOKD2L3+IPzn1gYPmX01dEr29t+pI8tB39r2M/XEkOzyxH5S8mTRJJbkj/JRQ
nNNQPoP/2WtlP0hW+MDGrwrkfxSOWHtVW/hKE3f0wfPmnpc37cZZ7/KJPCya+trf
of7Xd3NuAyIdBmbu602toLvz+ipvKQQ6OUtXsBlit2GRCsD3DOGZxQrHwwzVf+9y
+BkF0Je7c+zHpI4Prb3FaCZ0ubXj4cQ2rlZCaCqareuLlP+y7FWuCdxOb9mnM0/V
oZXTYvc2uEETkzO43EQwDNESuX3hGU4cjaTHavP8JpXr5iIbSqCL2EuqIk5v/ekH
zFn0h0jQYq2ex3ptMBeb+sBVcBkA+wMqehgHzDkHdtDjH0m2FVBJ9sRW0Mx1zJuB
bzUvFVKqB3j8yuyi8SYUyDIzeU3n7PxOlzbUHnGvez+bXMI3PbZ7lVwfn8n9IWl8
qblhGnYvAGfGJtCxk0X3c7UwyBSSz6TD769oOpYVv5QudIBcnjXYTPc7KErAMHjo
cN+il8ajatKI2vtjyl0YT4DA9JKc+DVgP7G34FhwSkhikw4X6NSKC4vXDNgZscwQ
2DpUSLOvA3bTQoE89qSFl81w8oBWhLGMqdFFIgiMWTS9uXZIRbYcsfysUJRQ+CLH
3cB5dZ/zehgVLZwlAym/6x99EvHYVhz1UB0HAR9ZQuuHSmE1kQifW93dq7fEpmFM
RPKqJWn7iD9861JYdSsrV2r7RrCXlqmrqg12LgAzkG9zYt/YOizHCM2EwIzXZ9DR
qXd1yD8yyjZwHd/gIDbHp33NX9A8ldcY78oXifKWm27pFoxMcr3uazaWfSctzCPc
dwZS5ah0QaPfFUeF6p/GB6GNHRoptDEjCmHtkDAdKjEmvS6SQwfK/EGdB8Vb/bfX
KoUZC028GAesappai8plgzN3zvVy0y1VUMlPFCzMTmS1yfXx1gULitCeqMv4jSwf
y2D4B8mQvUthxjhFOrKSgNz8/Y9jrlCduH0rvo4G3ttpzRIXBwNg/Yj+GoUlYAHw
NNVN1hBKHOG/+1XWj7OLWQN9gouhyjEO9M+iolUEb1HTOt4Lr+rGFxVBpKtPXH+m
cRKsdyWVu0XeKRNZ7NpQ6e9LlY+1NRp/uaujebUA5+WO2mMJVDwS4NRB6/S6r4IR
zB3uxLFyyFVeCVEdnxWZCbHEupxxEf8nldFm1B0JsApVhRu3CTYgcbsYx0IABzZD
pfkyYoXOFwJ7LrfWbgsmdb05o29xrJzHUSuEmEG54CUB2c5t1FEiB2Gup0oLJssB
u1RTTgFW93ZrXguhWUQMgn6Dly5Dx4PPc1X6ONipD+AiiHus8+J1aBRkirIPy7+i
WeALKixKs6TeuG7aWKMJA85B1+3lasIb/O0Yd6muJ8dV9OtitEgUrU9Lbr5SIH4u
mXQKGbsEqjo/XSOG4bNv/X9au61kZ8XDhUe3MWPITWLuB+kmAAj5rVYIn3EzxEJb
KB4ZYps4PK23a/uhG0fO5xuR3dn/N/347dqb1fYrorPjUqj1T6qkWQZhCPOmN9Xu
at8613sc08X5fWuLplo0DlnwMGLu924L1Ic+m5C/22Q8CzLh065D1d6aMa66CMwo
eCGp4pFYU4MWDosmYjfwY2FyXIhWcPJ2L0w2wAXS98IW/l+XfMQ9Gyc3dfKKpvw4
JslDA5lf0XfDLVZZmZl3j1jbkvr6lHSv3nze40cvnhO++1U7DOv9+BLycPjpfCDW
/SCSlpZKTgtY/UjPyQnYVO/hh4fKk1AQxzOFnTj+cK1MKRoBu38Uj4I+h9xkDWKZ
9ZK1J61b9+sLh+D5a/DX2NsTXQN3+ikxNrqZPtUGAdiI909+XiaV9WIrK4gbfE6P
/oAVJT6OUWoVoGvALlebXGePFm13xQOvuaOvwtg05QYVxVhqeyj1qRDhbyeQqyKb
CG9Lgqekdxtaq2Zsp4jiALASeFwTh0GwgGOm1Kz8DQkrkLP3rhQWOqoeNAJ508up
+DBcX1Xw8lfNL70Xy6V5wDQMH3rd3qDg1qf2zTkh68Fl6iqXskR5GkHUBGyAZq4I
1w786T/qAfm3yhe7vm0PTjFUr149BJs4v48lsCJ7+LIvMAVBmvoa39EfF47RYYMN
+5ZHRFPCKEAiQbMXtJgWHGT5NmlbTowHW4XrI8r6aenxRVRWrnu58gZIsF33ZE69
Bi5V3jeAzd9bg0qu7VB9j7au+ImxrsmDg2U/iJlkFIBYIQnBliXNdryKvy/8QEAG
mApQsto83y2mkqmp2ca+1BKWyubVM0upGJBS1HqtG23EDgeCekLbJHGCvpJqru5e
TF8C/0PzTS3UJnSysjF577oZJi1qi8N1j4WWA0uAk2sk9athPk8APXlrGxw+69Q+
MOC+13GzqNNhWcggirkurp0/wT2tm1Si7v2uOtMtmz84FXT3Z66GPvrASskuoRHl
lI7N+/zN4SERe0q/be+J7ESog3g8GVEzgSzyJMQFBiwtIfnFojxVUdspPYyrneHK
QbSxfTM3+s8oRZinNUGzjUmC+7f0MON1hwizWmobrzGJFZhi4eOTVqJWfJYbJZ2c
P9mMz2+DOyiAnX3tWcPRKhM2ZeK4H9GqixaUqMPPug9b+OgHBADoSb6K8tsvn/UI
Ion8onYUr995Kgn0Z3aCAKGg+uLZzj3NpKGeMEyZBYs/443dtqIOamh37jfECBPL
1ASgn72nC/WOScncdjrkqO4SaVRQWkz8yoy/8uTOT1GWMHxYVKP9TMxksM74Gh6D
jgZly+sQPI8teyGnhu0QLZIzJOI5YAVaHPjMActPZM5qWBORf8IyGHMh7LIYMTBU
1lbeTftQn2WgMURd4/van6/vtXbLvknHAkq8vSzL8KGDNWcnzUFMvVkSlBHyzfhp
pF9iP/+vJJ87m0+hmyBuc5+wtgx2pjfqbh8A+LS+DrkPCi5b2XoifYrOa6jYEaQG
9IZayQzhBumhgARkgYaR8P+3h1OPc9I7VKWOl388fOA9iSxNozBebEkqptHGnuDV
EL9LgXVG38Stuy3UWG1ozCXQ52HRvrC61jvokwzM/LoHsPxJXP836tLG+oNB3gJL
Mb+UnsVdjWD7I8u6E1WVgg67VGbXtwND9NEgMOtFZCxVgYRqewM+5JRgDIdcy0l/
+mNHoTlG3lcyn9MtLa8F0+Uu64t3JJYPqOiCO16bzKEtMevbCpe1IsyJDCqzZU4m
GiqDMw3UsrdCRFQp1BYug3+rxM8cOwjIqHNRzqrEFXM5iBbfrwLhW6HpLK8iADL6
Pu9CPLJ/q9KL3tEYmU+IUv6OpBbaggA78NqEz8f0DCSjErizJWuHpj2AISwXnyKw
ILQ8/geXX1C65wBkNjV+i1PjZljVWJ6oOY5empptVcfS4/aHborhsIxNNHDMvevz
504MK+z+F0FKRc+pvgSTWuAD0VNpdM9J4CgAGpcak7JescGkYIlXh9UwQ4kvuxtu
uj5VAqW+nBuUjcUEawLzuCldzRrlA22c2/0Yc8CO4W1W4/uHdP9LH+Sop5FhUH8z
3ZDW4NWG2TlfKsXQ2RBpcLaYtjYU2JJytqYP4gN5ZKoDbBQB3zJ78AiijCQ2mSix
0lpf07EifrW2NpWyLOE0GOoQl2ge3VbfGowayl1K8eTA2n9ULGZs9i7/CkIeHWve
qnMi0XhjXv89vGz1RUI5E5runDDVQvrbGSe9GAahhfBkR3Xh1PSm4dXNg8dTyK4P
q6uumKZ7BdcPuzacOCD0ZBF2CQx8yWZVHsoioG8S5qrL5pl2lxFbGdCMXY+jwVrS
6bIv1i6UuMqoGWRVNgfPlpSN0IaK4Y5rSz/fS6LfP0bclcNrs+MEtOCbPNil4nj1
+92oXSW3B3rXZG4awJ8e6gWuTDroD55EZrsyxnmyr6LRFhUwE1fBN6mZN9gYzSFd
fHRuUNMEcgErfkh3rooaDyttczCfIc/yYQJRL6dUwc3Xtl4VLTm4hYBg6mICZ+Sx
fpvRXVReIzQbeSmdAwVlx9/yyVU7kPyYM6QAo10DsAVHtnnL1FlKGcKWHGYytBZZ
Zj4RcgmF3fAuFypiLq1vO8z2v99IOgwbxlGLBw0xU9kahyrMjXIAkM319kq5SrDH
QlghigrQiNTXu/BtveMda2X0Xr0mtChBFzqCUKdMHC7+3Divw1jCqutFyIc0hLn9
57L3ePsGJOFJZsUDvjuQM3JYgH9Ndjsm6lXuLU58ctXF4ATvVTJGMF8EJJwuGTWp
JrE8w7RGPmSbzh4vhU4lEo86To518dBFTr2EIggiH/zOH3GpGSAToNkvtqdngFix
m4vSsnP1IHYuZz0lITwJH7DxidpZ6jsi/y+JVZQxFlH5/+vCWsM2/VyhaGQanhHd
0QPAQ0cW5Cr8XDSz0oLxyA1EwLae9i/rjAmFuz4T/9Cx3EACx1hRNmGn7+42O0BD
0cZyQr+JJNAzWRlw6fZ4G6a8Ud81bgodwNaX/yIXSKH/NKXfIMnLtQW8nagJDLG6
dNIGybX/YFk6Bx6LVJSHdz4/au66VLxwuhIfsq8m3x955krDkWpxuXDdYA8wTseO
B2fcD/BY3Rqzk2rF1rjIUk//w0jgrpLiBfMpcWYh4uoJYitiNGYCbp/kgwH/PUjM
2oMt6UbrSPLHxnIUoKOR8558Q+bfgwtghtiPoEbPmZ0aTSpp3fzlZQcY+l/G+9mm
5trNI0gaK1WUy6GpETmc2iFHMvBbHGMuhbi8zuf8chu6JaqhG9Mz57O8oWjhCGwx
B5EuZYSbi+z8F8KkX21NunSz3tfWrOXX0W/mwkJLVQnoqtRkwMP1QP14TWWBFEk0
D4TyUZUySPLDzJmr7U6zhEiqXBQwMgCQFAFG6tFF8nPR6wufk6jQhWE/s8vPaOSu
rRl0BvUSoEyO+1CJpI/9SAqXmJuapc5obI4GJYIJlGDfOSYoKbl+DkjO1+9hjslV
eZsjnc1SLcnRKjvjPZrOLxDasDxAFrPzCyzE4i/3O7mxUJKVLDv0yX4uT9A4DJx5
iY6bO6of5Es6LszSaXx1iDdaZS17VgumLEoI/2dXh37WdZ8Igtm7QA1bB73cbsCC
+ksVafWUWg3bhIo1emDX7VakgXRsU4oiIaNmwolGz4ekv/vTtT1D3HrN0yS0ehLw
RC7qwSTgvpTNha+uteol5K84Ky7bAt3OUnAcB+HPq20dKJlT/XfmuyGyKPx1T3zh
0yRL8EQ8D8W+XuYmeDF1F70tQ4Svqo14dsyFnDLRONrBixAUVKCg1FAQDSrEIxEz
Lo1d0mw7LjrdOGFJNXB2/CzI7m7UmQCBtxeMF5Urp3NZUqTJ+Q8Ft3dyNf0qTVvt
CFOzkvSIwhye3W99FGFcrBdBb+4DdNbzdyMVnpnhIerF2QaAntxVAqUCzzOpVlBd
8ICAMmgTINIjDPU6aC4NotI4V7v08tr246twglG+YRTN+4P5HxtnmYO8vlpyeGoH
J46YKXySKUfqQjI1uxsAPTNKk2oLqpLGMRNckw0u8okEdo50DCeS8yBVz/ccfdof
WmZB7I5+IHJI5w8SBdJkDSKbRM1AzDMhQ2MUp/3/cPEbCtrJb4jS4zGg1lsSvlsm
fWnOouv5Vs8PmrPM7HJTU9SR8LK5fA6TTW8n51wAkLPrUxKqzRZOia9qfdoshGLN
YmJRhntCNBErMOSJDaaIrZG8wHUrc6NdmxCSzNAKQ+jeW+8hFSufiPTZ/plA/MmW
tZFSNM5ggpnif5gdd/xSXxO2cH8B733vLZ/+Nesu3Xfd1D2GRWxCPwaCgtiUGGdn
hDI9UCYOIGoBdClWiGcEJV9OgcCS5PmpuALV+kBTJCm/4Ss4DqPz+Z7IsGTrpoXE
v2m52GqYTOBpZa/fz4cxyhxx9AbkWW1J6J7tpio4QQw1xJND9tk5uU+BYjh+Epja
msiKePce6J4nD/K2whBf4TV1afDqQFazuoU8VvKMvRJtjuWxrOSMOJQPcYUPO7ao
Pw2Sj8nR6eBgsd/QBLgby9qpOKiqemrcrO4ruQ6oxYT6+BwHVNq0dGHokoBDlFVT
vYIRQQQm22UKLI0P346okntBGVOjrGVfQaOuY6KJz+WgBGbsLEv1GoR86rLxoveK
GoM49E4Ofewzxjvq5dfmrxy4XFVCJxrMpDVEmUNsYvRh+PiAECw3gxigNlTkgBE0
XOVQEVNfj5Zb1B5RZ3dGLNPId13pGha7NROW6F2uNlXKgtv3bGMjZiTDLKg9ESgK
igxvmGAsLvVwl1tPa2YJU95YshIWMsjdV//3Ga8kjvyqlQITxpCQv5Zd3NJGbo5e
dF2IQbEUU9/cyEd1hG+HTYfKLn/w896amex1WXcBLFi3RP+XcPMEabCdq1QvGHho
oZoVkEJ46UMnzCmf2Kpu6aQBs8g2Dk/XvTescB8nH6m8JUibQnHFq+8YH28/w7L0
TBIzxFTNcBOSJ6bXS8hG/MmqSyG/r2MpTnIG3kXCSY5iv5d1pP5uzOdgOG0qkTaN
xEYKRaFKMbLj8QhCd04oXgBWRC0ICebd8+mybpIj/SG0rozqHRZcs5bSMtHPSLtQ
CiakiCTiRfN0nC0/9imW02DfiMaBVSsPzD/uJywLR9vGD003C0KwXuQYzvPidiIC
aa+j6LY+WWUtGqGVCYBfk/Mrx4k0Nnfy7DA8dHt3ptHCkPNJ91Fi15FKM4WIykoq
KsjKVBP6mtLud9rhEfJmHBygg7dq5xfg0/xTvO0DsLgxJzfLosEvn2Y2AX/wP3uC
XXVnqkbvX6zvSFwP1+Ae9/yqr2I/gNBtQyooTMtUxtHwExPRJLTXtnYw+E5atY/b
k6XILxCERDrjve4gObLrhgzb+Ec2fn+0ypv90T3/tzq3Ar5LqOQ4XyCl7sxu+Iij
1/sd3rj8aD7zYOQlESApPg8YUrMQMUfJO2EoWxuJ4LHsxlwxloYpxQFzfbNc8xyZ
R5xUn0etEYtbAf3lV1mLIz56mutsK/cdmqB7ngKCtKG0CLGYrRC/zsiWf3y0ob2G
9jE226x3kghBjF/UN0vg+Di2BMtlK7K3ljUBlJoaZ+/JdT9GTGqTCqsmFeInFcfW
Sj/hRP+8yctgC9TUAYMw6uR0QbOgUmIMArR2kgiZu7X5hmL+5H15eQRYgAhIoj6E
LQrUYIw9+AJkkTz9OiZo8Y7c3IcC/JIQDHCeQMIajo6yrRPQ2tqBEBFGW0oq1pvc
pTemHCXBNn2uBUtUV8ACerSvMT2smyDaOfwZp0lihUh5BuJO7gGDoM8woeZGeraH
vP6EAMDhCTznNLCDloJXF9p0hDbaahNHpC/62rMcciaNwGgJwM7a+6YZadOSO+HN
QECctLR/77c8CpGAfIiU0eBiNb1hH0lj1P4R37tg4fUpCuhku7rjRljHWlaxXw7L
W0O2cNlYruksoHnSUs7Tg5c/ErcJjbhNAEQ684KS+IWXeP1FXsEWrmMfqc4+GeZU
oqmVR2/xnUiS+zYHG47RjYemSLlYvLlCDZn37lQ8pIaNfSAThqN/YLByuGZNOh/A
GQxuWX644dCrvrb4X0G8RS7/6TKBqa56RoeyTht5kRBhO5TwNRDKGxBGWoBy7aui
47DyowwPU8SdkIeJA7v96ZEOyLL+UhumtU9jHdrYiBdaiM8K8NojvdxkCUjCX/u+
MznJYFtFYDb9Pitvajjvy49Atfc2evvM/yOTCck/Ep72CZIksyAi+HpqPGb9djx/
EpvuQVcZ+R2TA9suAEvPsxL24I/EDqT1fBJTnDt9k+hab0XKZ8hd0SuvuCbO/1Yi
/PsF///Q83usUZ9gMaQkM7O8KF3Z8FJfr2vcc+HwgPXgBgflFiuEUtsNiOc6OR8c
sGwopYSmhIqHwXtIZRLOBVIvHKQhZYvt2+iybAk4FSppNxn6H/PpU2Z8Sw6o/7Ht
2enytAkcEdzF/vnZ5AspQ5o4Yp/ySdWl2ytM1DXGqBbnTgBL2AXY841AY0rYpd2N
cBPYR7PbtHjof0uzR+ZkSKUhgKAWTjUOfuthxAcztr789TtfgrsQztqAV+8AW+gm
0v6jNQ93j09EgrH0WNLOcW6HmY76IPf9vQH1PzCYd1BHX+a9v3gKWXsOyX9gz2WY
Q/+ohrzq9of2s3oPfo3WUAgcReK0+WtQ8SovZq92v2CrvkgMS3tY9iIq7GVKdUiR
psCrfxqwQCdiTLUn3/C4oXRmcQXMlbn8lc8BeRxv/eXNtchm9MX9Du9eDhvojDn3
UAdjbDN/X51nbyJDtJoDFnUPI5uZkAjf8LWophZeEA+T14P1vKSgmc3IpP/9hJp/
vAn/Xw1FtTZqkfPisZ7PM6GjK6ktUQnhNSY9XBbXRB9C1l6sjjdtgh6KeGaa8cZC
oVu9TraZH+tz4QLi2YA9SCoHHeM4oSDaCiBV3PFIr079BHqOv+NarLohC/3N3MO9
cZUtOBhuIXreSTR5D7tVHiNbUaWBId70wmhkT/3ReY63qZenW42YJsvI+6qYdMd5
nz9zeoU6Ce6tNsHbFRzVvILRXu4L1sRRIBx9zo+GBVUYCUsNtfpHOqkw2j2Pi5Ug
JAPRvEv0LlHv9DLo7lb56mQsLfUFP/VeCgXmlyksLyjB3hLgk0vrEXyfSK8nX24N
KBM1tNhS2lWSmIf5z95RY+W9ygqShrWZap6SCx0PstxW/p5+l1EjU2/sOl15+I9B
XgS9aZbg98rAqY9mBBPAdJ8L1/eZ+lgfx8akB5bWs5ixpy7YGX03m7J0hlM6XA27
RzWSnp91tFLLIQot/Hdkz7cP4zMIQtEDiFkW8lpP/CwhsvMohdom4y9f+TDJTzzD
gCIniZLJUwrPN20U6tIfwNfYx1uWSc5fGv8Qe6gg3XqmYaEusgZ5ySmatcepRrpe
tMD0W0wwe5H63vtPY4N2DtVUayA6gl4FgKqwy3IhZsS0PYvVvC8tCDRrpvRGTz1N
UdlkN6HZGr+Avh9TpMj2nHbFDekxAbu/kSFpH4PQv2a218Dhqo7031FRK+8M7Cof
iOrb25vHC5pdeJoNwKFBNv4UtV/xmtGcdn4bhhMOuymywuEG2P0VYhYqjydflFFP
scTsraK16a6XWTg5QdFq53XHw15ne5tphaBrTXMBf+5aV3FGPafGFhELnkNgaiVJ
v6BWxnAWn9hTjAQZiIj8U/xpu42NsdeZnNu0C2I6A0DXFHcaIfBz4yn/hsSwiRIZ
CKmK7MktID8Ut+rymT3fBMKdH7iKAcXjorzo/HkqXP+t07oLHezBD644hhZtkBZ3
adIOn4/NQMGaRvYMNtSUu8crw+dAu/xwPASidC8NVZHJ5g3tR6PnYXNdYRJFsZIv
j16NmjHt+FWQqd69pEGJ9mB8Eyt6MD4yrrChfO0bJ/50pK6DkilaXb91IjWnGlEF
AvMvdKxmDNBstfXfGaGAAG0vnwmwNpGdtX2HEC/ZhAteMlA4YSKsqUXgwOVqmOHe
Sw4byH6qNS+9Xv4i9o8fOgJ72HSTB9moL2PNrj/Tvm3vwBWIGN9OhH6V6AMTKPXq
qMngLcAp8YZAA1cgCJcLiTvVwssxLQqWXv94WgVO2l0vmaFe5AlSKlWOmR0jZIX6
m5DwLJuEIb0qb1lKF6H2ly+I308vbPNju4k3WWhZFpuf9w99ywE9fBBFt8xLl82u
vN5dQLdVXxAIQkwXpBM3CoxrzbSMLC1ag5wtdRoYfuc4UTwwW0g+kQ9rVg88PF+H
p/abw4fEnblJSw43Oph62qTiyUfWr+zYY8m5xD3zxlGljVLqcr1oePQAPSVs7Zkl
fzjqDZK6nvLCOuQ1ay1WcJucebCMqCSFcTt9qsmNtWHEbvef/GrLTaPIoFNbSRNI
2USLEnyc6RHkaio89yF4bfmZ09bZdgth21NAcuOqHjlSYe8scXhON/VnPz60wvWV
cHspUb82AD7LkUDUHzpc3Jas7h58rPT7GZAKi7k2MSdvKKm3YbcTsZ/fuOlk6Or7
hDUJ8L2Yvj71lX9sQ/Yw+6EfiGO1l0ciumce4aFtuuHYpIIznU2Vek57cYIfiGyi
Bp4DWnlePYkzgRepNyUqRuVXBcXIG+2dhxZczHj7jMb/2rQJjjcapzk+Srrm+c1/
ffQEverdUt5y9ujCGDHhQZUQnO9gDvkEALAD/sEPXIFu+jSIDISmzHFHjqEFxs1f
Fx9EMqwlzISjaffebQ+mhKJPPAvyAeDELiNNQwm7SQEQ1oCZxKUvbtZmXOlc4ZTh
IVGhoNkxA7m7KQFlN9MRVrMXiUYRXwZcXMTHNnB07at0jCDkzUA1vtVIEbMReyJF
sgwKQ5WZB69fOU5KHMAomM9ijZIP9EY+CgJQZeR3fcZGLMmzxzCd6eSax1ykwk8n
KQSUlVeSiYExcZ0K90mrd5VGJGvTkSAeEURfcbM8csKcc+JQvToEUN5q/ibsfa2M
aE4Hni+jE6csG/lLZseWMzSFkdYI+fZ9rRqzkRECRC63cqirz6lpFUMqNpR0Ff/A
FQ5LNIQUhyKq7MscSXb2QuCka8Eo1p6yVMM0FUsx/H4ZbIoI9SPESCEGeoNTjQuO
+qWcFnkRyc16OTG+nmIiFMNUO28Gqks3+43RBgeWrBD2qxaWALj4JX5XFiL2oS4L
J8C4IdbFRGKXghaSF9slGXqbwjaidpPt2EoBvFy9NuHPUfRhVIwNi2PrtI/yJXac
JMJQGz9ADJ639mPCu0Fi5f8ip52NYONWmB8BJIrU9iJrW2DHQjniVoNhkZ/h97aF
qxMdo8XD4jkS2HiB0YeNrmJf45LAP4UuH6mKrV9FJurVyu/Wh08bnSnKjRRqYxNI
j9LkfkzXzqFAZiWr+k3ue2+SFfSKEI6yBvy0CVQV8Nj8Z8o4bFCLD12H3xAKo9dn
gsOb9FRJTRG2a9A39GBmZsjg/ZAINzyrdvJNb1T/NDICjh+NBCWDYu9VaNx1Ht00
4xHyMcUvyGiVNJjvx6YkQdAaz/KevAKzm4LJBExxC9cyeTpPM9eR7YBBZLMTgWNb
Mq19hemd7NxVmdn7Pn0TYUrCXmfVYCNK90I4tQeSBpgunjyJTA/m9QsmeyBBLSTA
BKzC0fsYNjCccW/+36ULVnapKdTef6L1C30x9zn23x22FxORDXL7fUQCcBJ8kjIC
CMSlAmFG7Ei9Lpq0zfWH1k4ckkaVActRN2+lQnGPPqAuJXmMnb2pCfjHh6geO0sC
UK4iM2p5A/nf5Sl95HVv6eKKZDCTPRrh1Nj3RtJPplBwX7JqvjWDoPRTP6PTq+es
IWFaQiiBsz7wxCA3Vl5d+mkHC8DqCZi5gv/NQD4ZXnYP4uq4J7hsu8hKPm3KS/DE
0Z5dcHlZVGE4Q5YiK0e42nnwVns5abi31MAIP2IgXrqtNfxOw+AKu6kRN4moep2Y
DynsBPGe1/2E2mLdwLC8RAw4tX5CThgg8T7sYGBeZi7utxyMZVUnzwyAqDpfwMqK
ITh3sc24Dq0kkHSlshM0T7jgbfvlZAl0yNiJPYvI/lea4jzdOmnTZ9xnXnfL16al
q5B36+MNavuJWE8xakxgLt0sClWI/rnXEgd64HNnLhOQ5znO6qVjVmRQR4yd79eh
Rd9iWMyE/WdXw7DssCTDIC2VJ5cKuNFsYmx5jeG2oVyG+XtSUFqIXt/E5iDpbOIQ
1SKGCeyg3eOiZTmX8FvUHvRg2Qq4ZwGZMeix03SfHjxkheSVsEXjbdiLToPZjxKx
WoZ5DGm8Viv9XrGYAdaSJO6eIScwBbCbFuPDiJ/vwO9qHhSeZfc/tfuLrioXwD3L
qQHsKxfUtbedT2rzHa1sIu1TDxZ3fo9tZooKlE9IwbGKu22C4RHjJA1zm4JKPMt3
SeOkkmTDDP68YFZsY1EiXBlJ0wp+ECC/vRIwzIw6r+AeHdnU9kT1P8SvOaTzYNRo
/03tA0J5YKEpzGtqBa4/MRf2d29JcpxxqFJiHM38+gILvLtudevZQj6/uDQicxk0
0bdVRAA+n5YX0hI7LMk9HmYzPPxVkshsRzyzACLKur4ok6JiItT7AAa6xd6q16Jg
I9//AziClqitNKD9HNpCn/Ow48pTorlmo7OofOMoax+1pqyEblUf/sWnxQrqCu87
Nw61WP6setnbIB9ZaGANrVvUEPlUmdnYcmvMMQSk1RYBmGfbTrNTdLv/xgSMH6EZ
odI8Co8lKwMlrXK0yCgpoY1XNacw1YthDPm6O1lxGg84MtMHNYrjzHL6OEboWvCe
LxyAXfl6Grua/uK7htzs83Xgf8W5t4cKpLpdh5hbFdrnnZsiPxsfHh6LPIz1sOMG
NdivK4cmGDbvv1ZW1lQRCHeOCKq4jN+7/6XZsAaOu21+bwtFm00xJDrb/JJh4ZSx
MUbvTW8iPHNZhG/XPCSGG8Ec6TCkXaNxIj0Kuw3s3VEY/oEvXi3RpvHG+4ZgVTFK
Cqgb+rV/hE+a4IOuHz1atY2x0Qiwb6X+6jgp4zZI2li5sNp8TKu23IVl7CKiBeZB
lNIansU2/oznknyeRbHQPRVcfDSB8/NRD4d4i1QunqxWgLLduCmj3v7ihdVOU1KV
8A6uFpmX7OtdKQzCbtCt5EoI4gQmIT/AJ6hlOXQVjYA00w8Cur0TohW6Vh7+E3+a
O/nNeSnrhA3g/A10NN8lcx1LT1+MQolgSikadMcenaN9c7V1JygJ5XtVibbrzWoW
gfyDAXNdXZNVwXs8DEZo3cai5C7imtUqRETw1naq7SxxkIwTxh3tuYX6vWbGqIlx
LC/hqohma6OxJRUD6hS5NQZjLattcr+SPRDC8jyM7nkQKa5HblDTpdZ/+o7Tp2o4
MOTFtrIQMWaBIXJ5gqbykeFvGvK0Np4CJ7Tu8Y9p1zBu8qth4YatET3CPsFrrDVJ
Sf/Qj16DVgOK2vwxGQPpUFRuEXLZnHnZkPqEbXd3SrZmB36V3KUVIwul9QfdxEAj
IHa8dM9D/pSQhd6SvSj0y/Nnozbogmz3dhvtbNLiQE5W1z+cdqlpB9H4Ggi59Off
VXldNz4v/TjJm9bCHh0/0TwbUY7xPp1eCwQ9chXxLchIJHczZ/Uv/2rt6hpMgcRP
greCn+B+m0el1adJHw4F9BCUV1z8wZS6UaVq7+L7/ZE97/0GVjy7Pu5z5b4QXYNZ
7UNyh/Y9WfDpeHqv9hRkalysyz173BHUunaFEOR38LPCmg/zB3sPe5aymlJrzlG9
U1herS4zrHoqSXIOkvdjpNbXB/mZUtrfLmCUmQgPIw94EpnqGkSCNrrc3bQkhp4c
s9rHXWOqgeB3lTl5Lc1B786Qs61lOwOBYLZ9zC1qgudTxp1UB4pwx3wYGS7C1vf5
czG9j6BRJX7yq4xlF6KeUWvtIg1rBdu06XY4TN8Ru0w1fND2J36bHsMmL23dd0m1
45/8gwnt7YPpO3uPzJsMTcI7bLfXlQY9aF0WQqUosaO/hUjODvOuV78NQ/11rgXW
zZc6t83UFkiROZzv21jsHezKkBGHgI+F3uKgpmlf3Wzb9/r0eQEJBinthSpKB5q1
jfNEJMxK0cvil/Fx1GDKK8FW8Sc63JMoPQU9el815TTf8R+4plqieiuSDaxZOylB
psp9jhk7o4sFtonf+S9quQXiAQSRKtZs86nE031n+d82+UO2F3qNOBgLNkfrc2ay
Qoh8NSRvHFt9nznk/uKsMNwXKw3wSyYKxsqgNOa3AKg48qVl18kC7SsbmdGhLs+c
c0F24nXpLEvIqb5FnkbI6a6K9YQELAMhzsudDgcqC59HwzeUIU/6STf0Ufl5hxZ6
0guD93uQcXMxRrDw+icWVi09uk/ie9OaF3KqDrSDm6wmyW+dle2+i+lgCbQJ23Fl
sVnQoMTKHC/dyEfkthTxnNTK3fE70CmXMSOEoZjFBx0tkSs8xto7Uu2gx+5GIVEy
Br2fPkwYXH8icVRNunYd1CSK2xEYMD6RWMnfledJ/xmNEojp+jE3T2Ng4pxv4nUV
HR2GAlHQ1TLIWWeSyGY5/VyU5PZDFxsqjJZ7e2hW6SWAzdo8l1l325RNKcnNtp5N
cDPifRAYRnvAHgdMmIL02zO+aHrCafTnOdwsm64brqDNNQQoPer0AhwWLztwLazk
VWh3iIFhIhyT//rb5VL64vSYVh37pb6WhgyMdXjKc5j2HsirQI/1Kl/Km55B7aKR
YS7aU3s/Ni88HYEtJICHeXh9D6rVShhxCu0kcsfRC3v4b6ZDiEMDQ7//caY24/KL
i235ATDpy0lkUL77x54Nu8Upa+oU/pxt87XGr0vBchK9lDHGBkqO/NkDx0xOzEjc
dbkjaXDVzvcH4kjIhrli4IMW7Qs9X52kGeFx8xxRwDFmpzy6imfactZfYmZ+g4ky
FWQrlJGaK6SoNS77chhG7Hb5sR8/iikoxNWGvkUY9L9K0596EB9D4KjXBplS59nm
gK6p2PZTn3/yMMPKqqaq3Er+dMuNXyvp0Xd82ACe1w+3hiHDKh/TaZ3No3WCzT0K
Ih3Q7C+uYmyhYk0pkveoSb/ftr7USVMDn532jl1PH1eN2cuT4M2bun8JFv0Hw6gs
RZdMHWxPphM5sDk4OwzNe/49sQcRUcnaTpPhVq7YvDP59VRDmfiAXVJg3gdWu5q3
MUncEQngII+EmhhiopyBQiQd6Lc2Aen2am+RexYfkfpvVAmAy9pKuJQ7u4E8ukjk
Pd9FbQm+vn5GaKgf6iV26hhtTbWr5HFHMX/qvHq5EVLGxz6uZqB29OgG+wqAtFJb
WMu38YjhMtf8+5G5wOKGfnVZrq6lyGrqBnjWU5FAr3EvGWJVqtCKzTJ1FWuh6pID
VQoEXny9tYRN+odHf2rIYXvQlATr95FmE5MCb42mW4AWisu0gL73fXWQftHUDaf9
WPAyE2KTljP6xWDDsJP2qUBis+Lsb4TrCMhCT0OaxfrEHtOZvKOuPwAiUJSZYZfI
rV+KZAZCkWFT0PyKp/h9IJTg4sQwb0M54MJH4vsKTCxWyaAX6QOtGH6hMKWLAJdq
kdMaWi4PXcFtXnGI2TGCOohe90lUFoRJGA3Jg285gKSCubuUFB4IzDUsYaKCtit3
CmwrhcZnZ+sSHcdOxnj93nn8eBxcZmIuutQWJNb7ED789ElHE4l+8gIbB1f+z7FQ
bgbqmRtC1Fegt5a3OswgIV17Q8/yBimDJipWoEQGV4Ops5mgHfOrJzm3Z/HwG5La
L2DOdRjh36USuRBJywbffjpUNl0UDZyFpxAqsPxi2CK4O7ui+OxLvFrFqpZEKAj9
CnvwZzEMAzMPvXPioUGFepVTfH6tg1XICTuZhCUWwvqx3tIkFibuMIt9y0/kPIZ5
a0x84uiO5SwIvZiCn0zawkPlZC6q4BvgYgRdhPGqJOdmLK1UK8cXql2c5s9znKAc
tYgMQ/l5vrFAE79oSq176bKJtXv2w7aeRu0EJHoWzkZqfzaVUBUodRaHnrAmY0lF
sX61w+Sq5a1ytP0XdXzroAK25Ob75mKLmqu/ijIVfmUX53WMl0wuwuEzagoFXpCX
NvfOgtULpy34GcDKEV/UuNh7CdG0mauIng5ZQ31I/gKJ6wkjQ1nOsC+ZaELLkK3l
k8leRhrgS9y4tIzPMlnOgKabbig7UxAh9K6KJUdqxNJ0VCjTM9TrQuL8yiLDnSZT
lD5M9TdFx5ZCf7fLynO10kW9UfriFKzhsGTNOP60OP2RG2nq/NyY7zopOTStMVfa
YsYqZaSfFAHdJZbgPLZdaAfOszk4/9DVpKCcbDKl4mjSlzoLevibOQPSKnYgxeGp
Oi+duKN8xsTiZxdl/OIczfHKrCoU+OzweWp/srQXEL0DQsjGD7cyfLmLhzJm5XKf
Z31TT31PUKSUBXtAc4paq2g2edOb+OZxRT11CLEUStuaHMPmgQSd0aSvJ+bTPOQ6
erG1DVGqC5w+x6UdGUi6J2Nno/+vAIGBFjkIP2Ygpsby/fpRx7kQVFp7SAmd6S8p
YCUE1yyyyIlm8OpVMEWgQVvCeKujKX5N+W9ELcJ7Qka5kGywWwQKrSCeMZR2JBA+
qgLKcsmsZZJSUkZQ25tdS5XDBxNnVTnNgVxMpHd7iwxXl/E0ryJGB0acn2v5wmqz
F6o5E/1cq9AK3uXuQAdvj4tfbzY/Y6y9MD6qboILt6QW8O6wKuHxM7A7ji626+Pp
oVdlqHOyCzNzcQ6JlYXW02lXFzsgl2RziQJNqdkoLWo5cV9NBjhM/OhJygf8G1u5
TbWqI46O7iLm4GEbIOHylwzlQb6UlW8b497FoYstWcroFwzHWLaM7r2bCwUAUaJu
5PiJRRBr3UPlKMguSrpoZzVkKcm74ChwOVUUOlMyREGIn58NbkQgw9DJFNYuh2eY
YzgxSnjVAF8FSDofxkDLvhx9/Zi6a59Oxkce1/g5lJbbIYiA2tJcQxXngrbJ/UbV
/nr/+g5d3Fd8F2cey5iscocPsiR06MHmZ3pYuKLiepEUMirO+trcShTT+qn4WBzp
L7Ajc2RMKP5YHKAcBAWw+nDqQTYoszzo2o9etp5WO2HkWax1nUauQnoj+N9fvhpv
jY6oDXtgeySQfQvwVT9Bh9MnjbJ/YHw4ElFUTiRfyYDsRvowqK0W/KDRdP1RNLOe
JB6W2350mJ5XKPU62ctDUBW0iNVKaKFimhFbhBtynmNuZcFrTKjn1K90/R0LJpWP
Sa1nqxksyQYq55dnQ3ztAsZi3TTtCVM5wFQp6fOxS2xoIW4vZ74mlaBZBxVyIdDp
sGeenZYBeraovkKsAHgBijYgh9ZzyolCcspj7I99aUSszZM78rNJBiB5TdFoRKnc
FuByrg7mclAMZHIWGUC4Kw1a2teNcuDLbzM22Tlt0JFoW/yTyb2GmpVGAmOcE+je
6v4MuUy44EDsNYBzXSsp15m16NoMvBUyg7QbWG2BjyeoTHBuMiz093nE0EFfibE4
Q31vywPVzRyAWGr2E31JyXvJdAsROph5NPcXuwND6CV1jSNM7FNsmLlExIXyMLr8
cgWldGLpZn48UIMr/UJIwXbRyefoVIJHw+R7ggjKHaOAvsRvrpQqy9Svqp8qk8vd
cn5R0dfk0zRPwc25V7hpXoOevIAAzahb1KGiFSq2CGxy0cse5Vtqu8dAqfSJHmGY
tbSpClbyDFqV9mzgo6FPDZTYL8E9Q8sa+OzXgeddKiJrESWhDUcRlcEYHgvPyGQM
QwUz9JJlJ25oMeq5ACoBzeianpxyhOeLi8LptDFrS/5CUBznpPK3rQZZNmHtBq1w
YjexHOzO7ho+AaHqpyWIzbqqNwGAKNRBdOUxadN1e1dXwd0LMUCc07uTYEEW6/aw
o7NBuBfZ/0UVEtwVDMcT+vLlnIX4e9dUYoH8X2wzZ6jaFZFxRsjSNBYG+75P/p1M
WAf07zcRpbJ+LQWcnns1WNCfvGwCPRWRKKoEyVj4VvXcRM/32bEhgpJbxVybPXng
sYJMziN+DnGoIgaGb4O3Hq9lNRgEH2dYButTHGA4TFW7L87Vhuog+AszzhI5G+R4
HdYBCMLrc1RiN2EfTOINFHG4pCqgOMAVXhnSVkKen6Ps446TfA/ZSypy58tHDYZ7
tIRjEkp3GlTmojsvuhr3mWYLw8r3bbOqXcCG6dzN9HKZtij3QAatlZkJIewvZMFX
c77WFG3qJwOFlOtKAc8nxdN2+odKyimpuOGsbF1a4/nUS/rc1K+RwfFBVHxqUlvD
x4Kmnv1Zbsx8UJt3g66BybB5j2tnn7JX7VNDOrBan3fAcbAo6p/mTXEnn8MHmNOB
06PH5wY8Y4kry3Cq5wP1hLYwhkkGgw6H9pQvgvAQvsVSKCZY55SdZ855CIeH+HdI
Ir7YHG+iRl5Gs3K8yVjn3ZFlX51a5wWIVxiDPecocp71eKWdEgOt7BplRG1Br2M1
Glwhzh0awpJg1O90L1GfT6unU00REyo4T7rchfVNdg1NC4qqgLBj3kGHmmI2cSeo
EhCO6lNP+jpBy5342WdI2H1u//6v5Oa256vteKodBmp+EGBhQmTZORZkh0pJ6L+N
MRRuxahMFk7rY9bfZbBl4quMPW1YsxMze7ZP2ZClWKRMDty6Hd7desUgU4cmUC5h
rHHmVJwU7urZgt82V1vodhJ2X/q6Tv3DxE3K8Epes0M9/Kevk3o+G3h8QRfYfCfc
pNe1GXjnvSWf+Sv1GPRow7BbQp36W28xZup43ssuwYldrquYRGmS1qb14+7DAu3e
J11JE8VIDFwGVypSd12JX72b3iHpc2LXVyQoFRTnr6pMNyy0QNDMuepo16EGehTS
DAqTWyZY91YX3KxDlBFXHlprpNln1mDB11mI5LrrXRf9b+VuZKaFadVZHW/8ycDR
XjETdPGhD9go1jn9CQjoGiAJcVsjr3+svgv9IiERNsMVh850v8x9jvbtgA7sYMwD
IuydZma2Hw4i0QyL1xaPpMo4yJXKAOqy+BWxlM/Ku/tWdt5iQoyhFkK1wIaX89q2
FwPwoW/gVWl/Iiz4n98tHSDrTRGwCw4NhlZviHZ00vqor7pjxkLfG4EzciuzQNkK
6hWxr/ePQW0ng9O731OaZ1XvC2PQoPEzDDk35D/8jIYmsTmWoO61AHp7W0Zm49Jt
mOS9MxvkAm2pNq5cPFvQS2ARNRYLGru4DHnROJlD4NX72yK2bt9/KLmyVblhPzEh
AbeMR/S6wIB5XlVzJO0q6cFfnWZ+5NAsuTbjddruNWFYWBI3YsE9c1l3Fw86xlQO
KzbyBSat6GflTp9uVRksFnn1GdMxZt/WArhiqW6X+SNyYKxu+S7iXU12lQ8YL2Fw
4l7G/djJMaxyGSnrWTR+avIk5o8qNK4Zg/fqGv0z0+80+d2+BLRnZKXcxttv1iZP
UpwnRzakEQr3sh/alvl44uYBV6n7Faa4bBpqE1DHlEWUexDu/WTl//iMvlQTYonQ
NWxjmCvlHPTjuaI1goduIst9zWKALna/Q9Sb7bP8xKyzxDJh7oZj4Q3EDDF4Yf4z
gckfRsAZTf4+HtsCv9iVNygGgaX5LK3MvotHhuc74XYInP/E0FKvXqj/7gj+tDWt
DVsVwuhWF5uI5XaLCYUg5O6a8W0b4OZgY+k7ObwKsea2H1NlwghlqyyeTzNQzizo
BYE/Kk8+mSny4TPWxoe36gx1vUp+l8asxM2Fl6Min45ujC5QTyNlfizPxPhyy0XD
aOJTsVIwFY7h9jlZfKXF/sPNXG/H4JEiQ4eiRi1o7tUNAE8SHvi8O/3sRH9D2fiN
3khs61r22xzybh0r/W5vL7frwzySKvBG3VSZDoiLf+c9Td1OU1cUFeljqZz1S8rL
FE3h/wsKtTRrzi3SqbtpiIw9jGii1clQ2/5pyserJPtfHd9XgfFh2oh6P5Y7CHP+
nFebo6Yrke4o0YsthReESu0YgtqEsJqyUSISeqbD5BWN1cGNfpVbNYl1rmM1lOhB
HRJHw+EzsIUQVRZy6rk2zucGizxEDShMj4XLSlRHRxypSMHMrit3f0B5OTKqEj7x
/flJ34dRh69ksORQwB89daokA99sJ3vm9u3ks9fs3sXVwdy5uraKuDv3R2KdoOZ9
Ln9Qb7AxCR5thpRIVhytxSgwDJ1bniH8j1EHcqo5pPy8pNK88J+H2xHcIsmuhOy5
Ja+JwutgRr5zF/P3jejjN+6WJHa8qODvleO544xqW/rL3EBOKS2ho71UtoanPfoN
PVCxOXkj9ktoXWv2jrYddkpcsBnXF1YfUM0i7/u9yUPQsmpwgtmuKNSXryMWdIGF
7zPM+w74WuI+9EjpZGhlRv68j7SEH1aiO5O0Kb2XaJNAIi/0g1Ust6VtJn4H4PDn
jOdMJiWKkSnPOIg1kYoptKrmbWMLayhDlX3tYPd8uGtVZD9lIxfOkLGbUfZvV83m
R1Itawr5jRKNaySNrlXxa0PmyBg+wqWjoKCkf5GBgjnQ9QQbtod5RYLmRMXlDpip
VSPO6mkxC37o+F84Iu9mltzmARDTaIY6b3FjKo0YXlNboI3j/m5cEM/K7L4WKPqn
9H1eLoo1qidEnkMuRamFrSbJMZELMKPYd52+3toJL/3cevJm+1uwpaB3//wJDMlf
N5YmuqpGlDMC1q5U0b6Qd8XKeHriCEINk96jfECvmrY/cShU2udg0wXs3V/BTENi
3V8VmpYjDFbewh9XwJRNGHsJoehpb+q3iWahIUY8fHQqZsClJ/o2J5CozHzVRBkM
WpwFGHbeXhYjTQdeNG9PYLP4DvPWDCXTBmJKouYWX8jQutaoCpk7IXjbW+D7waFr
yUmhS0jVBI28AOZvbx1YV/J78XuXk0Zzq5c1bwas6xG0xiIjVwDXRmTvT6aCebog
TVG/YGDuXwgbSenWIJfUbpGqs5HpMq39cshh+AOgVd4Jces9R7bBILObXhSMCch+
2pHn7LG37J9/+2OaNhQ2NO7HXjoVA5U4JpWbrr1unYwh5ogYmdqN7CdaYSBH8Lp4
f0BC4MhDD1mdhSZ8Ti4Ylk9gC65npUfe9CeeoWOJt5einx0PDxPgcyHgNcbKhWHB
Lx7QSr6CShH7RBYGWceluzuzmV9vE/Sl9XO/eg1rLxXd47+EKHexCu4/kPumWtk9
znzDPiJ3ENfLxr0bPcUqGOP34HFqbdtSOsUr6ILihvGTcve/bEhaQ9DEnkNlkUZ6
6BGxhGQC4COehSmDs58VCBqA9O2g3aUVylv1TCQCOhCr0f0HuI6E1RAtk4Cqh783
suwlB132KHaS0N98lDZot5YFhMsCQk0kTzJzBF11EA84KsSXsMLkYhNWWvRs8c2N
wiFmNDB1Gn6JP5fhMBfTou/HrHOEORxQtQG36gwTrUNz0OMJdUC09ZZLXzUusRRN
vzvgc5uovg/Gf3J32WWrBNSLsywxEqgtMKRs7ovbDNxcL60N5FKEaZA/RhxvoIyY
y4ZeO36ktdhWAZVPcvJCz9wuQ/3nbb96Jtqsjj4jPfupfRw3uw5maZATq3w6VrMV
uK6ZL+Weuzji2oE9Szsiv/RbXr870KNxSg9joUGu3TICtTrUXd0MDEDya9YdGKt3
U+dlPpDYIPjG18kBWV8GshYeyJxtPDyDoJcqW2RNY1HYTwKckX/Ij6JNNdiIWIeH
TUgNBrT2BOOlxzF7DNUafHLcjPLjT+xvW6rQIt4K90cbj6eJ084aMucEL/TymW+R
3LlusxUYeekg4uFOWPWiC/O9CGXtc28tV6pSfG7NWuPUl57OVi2JcDXBSJHUG0iO
l0xBRbmvdu1QTXI4ZTC4XcK3s25MBRJsZBS5bAiJVW7H5zkAwgQxQ2Sf6vBV74jj
kfGIxvHCrdLPnEakO/if6KqZz5bf+YRusg2+EkgU9HeG0CkclgyVfr8zcaE0sjHh
39u3LuDadNGlsASw8Rwx7O1wl1Uw0+7nZa0N95hvOX5tTGMY0Y1qGmlK89/CsNV5
MNe5FosKwWHwjbHZfW7NZMt2sBCctBTC2XLTPl/xu8Em6Al6GeD15igDrIZJ1pzu
m+8HPC+pFI749Owdk30DQ6uORh4DDNvEM5pOh+4uN30DlrmBVjcQEoI2wPCzcpPR
0TQ20FyjLW3SsK6tMf+YnljnYHLqogDeZU/C3Q/6hnzzQxh7F1uwwP/l3dq9u6aw
x69JtvncDxPqPNwfh1Vl+psRePZirMjQIB55c5cg1femV173+TCpCsyP0BDlssAd
kCmZdbQoMLUzGJl5dFuoSsjrVjKE2r2bEo7r2t4sZ/hPxNuLqiPLMBzEv9xHgI5E
2vJD/P+a02MXbBIc3cC3lvFukhP6fzwzhEQmE6z9ZnYwHxv1OOA7fjgrU4icjqtZ
Qclggqy9FXOWolg/gkI595h9GN4jM9oO5dtBDdNXVnWmIXh9bUnDfBE6qXLVn5yL
6flouOWBy2bhqgU/FmWgBXBCaExMZrSIcY2f8MfDKdiRYoCRX18Th/K9Z1L2Xg0R
ztaPtkRdnYZhu2N9/yg3q1ZB/XyLxZ/ob8hftq+4hvhq5bsnWIYHM23P/0xqBrVh
IHv23xUg/sLYndwzOgHc6Sp/57sSfgE1cy5qJ6hsQElpXuxdHggk20jlhcfFd7E3
oghyzLaoKlKW4vxTIAcibhGiz1lkW+UjSZdjQySLk5a6ex31iesZKUVrSRDJauM2
6YfTQs2N+AjnvNeXUnnbv6jwnoL92FV1N7hLjbxbu3SMRiO1zkkzC6n5B6HgY164
KE76PhVmX5gTmtOWeFp/yMvGlfuCJuuyTYXTE9V2BF9N9oIQChFzmJh9RTrqEbSh
Coo8CFWo6CsqKw/bYRTJQ74xDvOYJOD0yPU93Z0NyVvuqFwZwNINI9UzokaQEUMA
40U3MjSkIV62R1scImIdV5R6BWG2WHC2oC3imSNxnBJ1DfeDNmQg2OP1uPyhsLP0
uVCy/j1USeSaWuPagZqS68OZc5BWu92q5Ry88A1VITRRI3kFTolhYDKXC+5pC9Bh
Z6ZCAI9QSaDFTbcOw1q1geA+y6H16Q1kH47Vc+RcgY3Peg2DGN1vzsPdLMn6yRsa
jHEsUEAD9RDSwlKhkazmNae1wAi6H1Tu2zkGXdZU0zVqvaQe40yG3H3+Vc7y236N
UJUAG9+OADAssPyv14bfvf0vcJv//m6ZISwMUJmzm8r+kEsXQkqrVUq2fUu9pR73
7CxeD3xyf2UGJXvcZU8Befuaqi+D1SMg8VECniOsU18lhXnKqEb8K+10Kd6x5pOe
PA45Bxa/E8MVtOkpMzb25Czb7iaY2hj3zu9ntSEHbfJ9ysU5IPwdED9047COqBU0
5VTYuYVT3DWYdXsTEUVwItMgPB/VY+EV+SsVQSqfaC978Y+4Wk7Z1y2ydchsU2Yx
CTUYQUDYQemQUSEZj669oi3FJfyV2dG/e+tf9Y+ucd3GZTjrphIofREzKxXu5g8u
nNEmJh9p+dI6BZTDXVJ7GKG6sPhAlOPcgpxwsMjb6JMGVyPHCD7eJA+5c7plPIA/
+0x7AZD6pgTYO8pp3zAvrUBbaXeDbg+uJwWhLWLU/1gYxGRAHJqQ/wOv2CMGMeTQ
9+0n7jt+HOlROI8o8X4wU9+TffcVsap3B0hRJq8Kt/GTqq3WH8jQ3Wdtsg3t/SG9
djsgsagecXEhY6CManTFh2ZeP/PfRjrL8gxnlrHpfkAWoTHipzx3YebEaPPEAJE4
j1LkCa7QaYCo5AmBQ7Td+cSe7nEpBNAfXcfaKyQlnkurClPGxJfmeeBmMAMGtPHT
LytR8Velxeq1MVpLR6wGlqG6W0YwtURWuW5zs+YWPtvWrtYhQcBU9mMHR7+RZg1/
HFZjxnTiscrpbu9gkG54t2sFzbOI+peAqgdof4mQUtZZOK+qhg9ED9di/I8n0Had
cYROZ5ja42zT4dFT9uMKAB3kjWBl3MTlv34/AKJU0rRSrkSL+HfK7jGlsbrnWyjy
H/hR7ijLMEvpzY6aMzTuQ+O57op7B4ufbGGvsCN3NR53HcKFDrVUoK/mJbyBds87
ycSeTPPZW6g0wm5AzULsfyyHoaehUIG7hhgGW2XCOsncF9f+Q2EXG0+KyT7z+quj
u/IO8tsa/iMQu/dc+sV+U4csxb6ZaMuzWqkgRBW1xOStAQf7JboPRbixO+3WnASQ
43z1aoAOgq3FEOX7wThYe3cRBmWBgupOYDvUJ3xkRyWSRxe7JvKjLv3Nt3DncnsM
lU8JlYEA+yoX+yApduLceoK6Ziu6legXQBjjNzp71HQHkAsc3HeWXADUa6y828nV
mcIgPISyEUgkLS/Pg2uuBA9W0gvorQyYd7j/6NF9aSjc7cXF3oO1D8cIWVRFDFzL
fJYqEREW0W7blO5CplDp9TEgs3T906Mkrr72WpRzgsxI7Aa+J2PrZIu6bzfNUcaA
OiRAiaXbxbPP2JiVhl7ioxFSFC64w0Zkt2CO4+pJADk/fdDR9Mu/yUJ2YuVIc0bK
9QXhOv89hs4Av2Ns6Ej+rNORFduoKyycm6rKH6BExQm9k5FHj8nQkt3g4UvUiAdG
TmH0N8BvcdAH9eiYDJzQW1aFNRnSicAzLiPRgMizGQagGP0GGO52+rBQztVOxssm
flASbE5/fO74r1FK3vfncPyET94+KFzUahXZsqnpi87PWEsdaELdAOLW+KJ8MDQ8
cwQhiuBo4awfTKbROyzJV1eCQvKhZYOhxxGx47yBwgMji+geoqFsc1LDg6BaOjyx
TklW1j/BldSdLH5S7uWAciwHFNppXWXpfF+IfRZlQOLLYF6kKjXFjgc891rq2WlZ
xcDOEk159fOf2f1LX0qGyWq2h0EMcrVmFP3kD8iPhvtAQHH73VjfdPQvPJLQQ0LQ
JFZgxDTbOOrL3V/BAAmBYv35z4XUZObxbEFfIfD/7PcoQ+vmVkKGB7htBwdzY4F8
KXgGmL7zFM2G7IHGC+qA+SK+d6jya/ja0upmMcFFgVHF9eMPYQ9Iy+jMEIFK8+Qm
BGnsjMvOEggw3He5D0Q3LVWM9mf050G7Ig/0v/kyENSTFI4j3JcaZKipU3faLFu1
m3z2lqVGPWJrXRkm2lLsw22fPl5pOu26XtI0q1mF9IymWF2xh2y+qUPpUkDIuDvm
ZoN5KuVPpIVEpwBATtWRlng4/OQ8t7tDjEOtMVtkcep9EM/vfmiEjk+ibdiwVUB/
BjnxROW17G0eRQ+AlxJ/Fywea846wjpdkUFT6sWZKXIC1dC/SJHsdXL5t3M4PHrm
hNWHwSbSR+kekjO9nzU+jf8FgI9mb3m9XLv2Ndu/J8PCNBQkQndrYkDI4VlRJLTP
nNDVdTQ0Ppdcqz+RqlPmyZwSUPsRgvQOpyczxvbXUM/TLVUOOt67qxqOgc1R77KI
Hawtuq8n1Txmz5ipOdcecsGBgxwWSCd5u7swihLTqfWQYBHIcvDpo0at77Jlg5li
`protect END_PROTECTED
