`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nslROr42S6N1vigWeDc+pAawMaNYvMSdx1rplF4e6kUmFoqaKXgVPklC3WF/M2WQ
6ddHjsMgkDWyrytb0ruu5FrmdF7ijXnvH0A+8+09yBAHkPRydEJJTgfEk2ky6kyZ
Lf8Fd6ZdEum52UAs8RBFELop+gV7wpbEuJ0488NW1s3m5DDpwD6ajWTn8aHDAJIb
6FlEyGN5FsafJJ46fkBS5LmZQacjqLEadGBxlv/L7+eVlD+Roba0mNqBslFbMAM/
Z2wKX54Wzs3CTe9oEwpJxGEPx0hlPOJ2T0c7iuwire2MgyZcAgZKQd56S6CDZoPe
FV7pAhMlE840Xs4UA2DmGFPdmm3VUF69myUON/OgmYvrROGXku47E3NvM+oabQ2v
OBJGR5UYwd+Foy2kEVY+S51RHSkzW7nxB+RaHJlh81LZoTwc+p8MGjM7UT9jL2AD
FMFj7oRiKz1iICPZrktJFihxe+63qAXv0kjp+SaN2Z7ZD47ZkL+I1rHOwl8TC8NB
xdLgsglvHqDqbZ31tps1vTuhwygLgCxcgcEsFamgoI7bwTlPaLLpUNevd7VoTWwt
8ZmawSp6CY/OiCDZPijaVvJEVoGu1mhFrb66lfNIgmTMlY29/uF63NueRYdSgT30
wzGYObHKqaMcsBHLBo3ycZrpnzttOaXQu9mC7E0igAtH1DEv1gptKGH1CU1X9DNH
F7p6TpNGJvC0QN/eSl0rC/5UWQ6AU/jbDCz0pvsi1NqJa+C3rgRwgcmZDbz44UkV
qQPkr4fbeF30v+dfjlDWoto1JSejHwEquxSTKMF/ctDdxaavXNSqRQwZ38aoDqOA
YdRiytMM0pKygTIbo5yWEkAtcKruU+COBpBcXDPGuJ7CE+PqYXTtNYQOp78qsxSe
lR0YC0yTDQqP8C302S2O2v8IpTjb6DtPIi7i48Otu6/lWJ1AvvYTZQYhlcKXnxez
09iuzJlMlgtKEcrcOfLoTBtW9IV026eKzioIIMW5QeZas4D7A1stsGsfLBRWECvR
iIn8ySncUqUQdGkco7X/qlecldjtFzqA1WHtchr3nezPA3mYGxoVfcgBMjryVYwD
yYLBpVKRD8G2fqixjS6s9xPZM1ZMCT6Wx/k59a3ZnumbQtW5wXMeF3j2L2kX/1Nl
oJXJdop4hS3uuB/fNVIZgFpshV32QBnh2qmNcXyJy1jkusSn4wdFnX5qvXvZ2NFF
+O3CaHmjC0NAaRhpHw+9lWC/l02A786zkjp+byjNM9A51yWfnydD7J4s8op6a5iy
HE8aougy4nHBVM0MNLs9xuTUtCORdHYcF0iCdWKEWTADM6axabwuY9lQFPFswVc3
17MGNtRouNncVMFjaLPLc1DUrCnxGimtCw1Ky71VFCFjMttCivfJNTee58W3EoWh
JY88e75QuU3cGNP98WEBiOrr6/VTGesNeBebdcU9yWOarg8sfwDiAJ7eymCas6fs
r291krE0tsny7DDFVuud3jMheELXDYiIpuR0ztnPGe3tYcBKUZg87gmUKSK0Vbdn
rLu7qlIH9PuTWrFB2cuzOTFaw8LRgLPKQmJYvaIz8E4h+uqDrsw1D/Y03ckZNWx6
yT684xdD13DNkt+YPd2h+z3S1TCJ2/1kj9BwgfnLp1bgtlo3k6fDiWnNDulF2WFa
wH4I5nt5RXoCKVlN/3xkWhGW2ZTGW/TZXyTU7gB7I1UGtXfB8dGODmFbLIisI1iz
My6SaBmAFAoA4cH76BT00D8xzvRFBshhtnY134qOgkyEU5JHKoZdFMI9syZKFngt
Pywpib+FWm/p+MXHSgTu4iHZLeNupNNRdjW6dxNK3QG9hkJiL5YEJn7VIiCcJJxw
WqkGCSuBjeL5xMS4U0LvwqpDerCYaQcnHp9+vYG1kMcvoxA6/rHdJ+4JTuepgP1f
yCk35wDAJDI59hj1+qmzSLfEin2qdUiqqSV4pisLknc3NPVWjGhoVPs62k5qG+Mf
klB0ClS2iDtX/4o1Rk4/EaPnG7YoLNsj06HO+teh7wNx/7zL3XhvBPcREkZ4nBrh
Dhw58oGL2nD4SYQWCzmDjGfFxx0Ffp4znSQP612yC1+54pSs5zDg2B4mD2TofVO+
k/BTAVdvy91vFuR+zw0JBkx2fx3L6GTfbuAwAHa6UuBwM55vZCy2owET4dGELfLn
LelLWo7j5QqstBZBBPF5ppGSJkzKn+0tRUoUSMo4X6fevf8OSWy11Tz6jfo1nU+n
fpqfFPEXHAeAPZew04DoZW+GgzyQAsVeyKchF4q/AXmDA72tcRlRuqaAe9ecALfO
cQOOkXKDyEWW+WUPA73mrd/aIbimCQG5JSX0uscPFuhER1rSLhbmr08NdGp/HCyG
B4IXQLIpaelVsNsqL4SKczbzmMyOqmlC/bmLQFQaZwH0U+wwl0Hojj4WHbb16iN4
o2xtC5/T6z5ouCi7WeAckIaMc3eVFclyEP5n8Z2IDBqga8QxRv7j943Td7lVuJ3K
fZSEOzenFNAa1QAZllFsGavK9/YgBCJSmMS+y5LO3YzLuxPoLE0BMadAr9LDINBK
N9elDVZN8Uuge5voi/SdvT67ObUdGrOpa/WkV75kkJSWFNPbS/d6Lo9L8GH/Up74
u3x5JGz4rQet/+89062zqhWmko/dB4ogTFfELjndZeDgdaWsnceEPwwofwoSc42W
SO1kp5SeqkRmB9b8+SEC4uGMMCusBJkxG4PNUlnQPVSoRkiplG6sUn/gTp9qYneY
kb4qwjbLAH16vj6e92ZCYtSDJoJTDLwYR4+MPwMgDywhawemxFgv9afcRp+1CUYc
SzHZQVaGWWgnzJzsO2Ttv/np8hkEc3MLWUDOGFFL1YSuxekRWeNLFW1I38uKOZ/x
isHW0uHv3XzlYYZJjKy3K2xBRRsYcrEEyIbpfo4XoYaKz5ZyVA88voSfi7ru/JZh
kLMpU6/hqUeEnCeR9Je4rbBVL5gLsbRQJyYr7CcPK0hzcuvlRMmRdkTIwL2dZ3C1
WagI34DSOy8MXeN6MnratQmS5ERrkoBr8yD1vTn3oGTKSeK9X8rI5MKrP83nmyy9
D5nDOTyAmHywkVUJwntryGY9iHNjbGbwKAF7pg2Iu02TNcYShDON47C7Fjc7rTFV
526ZCS7F9FE1h+Y8Tym1x1/QLd/6DH4R9sT17DMtaqp/xymHK44gM783iqb3EV2W
RBb+EVTPVK+Dl4mejrlthwiq15xaa2Vu9Ob9goql2Yvv2DAyqxX84Zc3dgZJT7CU
iggaVMWY6y1dfh90fvj6aENHfI2HT/1k1tz8HxKF1KE06gD/w2aEQIh5mUs/XdVW
1ezdkm7bTEptKq2K6zsxN8/3FhY2YBACtCZ04IqYX6gfBJ7X37SfZaqLwHh9HpG+
w7ZWU2zs5LRLIG9+P8ycL45fwyz4er3yZcQ6uGOXb0usEpmzc1h+0iGBpgviJR52
i1a4NkQREtlqkSQqITwcg/o6Zpunnb1M+Q+QVPtOwyFRteSY9CgY7iD9AUfwJdk6
wuEv3MX0O8H+PnC5x5qNSFjmdbKG1lN7w+CU1ihWlvc2JWQSIoNeZhHcNnZl1BIe
5xr0OsJjtjrT/ZBzplExPnYrDENg8U3/bnFJhMOYVzg9qZJWKVI7+744Pf+34iOW
L+xiC3kHdR4ySc6ArMfsELr4XoUv+ZGrvLdqNlLm3BXA8D7/vwWhP+fP4P5QjeZV
2OJ92Tw13lo0qfSD7b3IwHPGzu20ZiSy4toqQaI3dWWQJ+7MpNX+xt0NWOdpmwBO
o5ch0cZf4bR6iChUjQwExTRJDivGhnDDUBv2RBV835DMyGf8aXmWQBAp0aYj79LB
DwKLZ7K7ghbif1ewGuWYIBXx4OCPH92zf64WXWI/KyDomYZHF/LS4FNEEQ9BsTht
jAgA6+CJBAeMgG0ZYFBf84sxkXcQscrk6RhIdfJadiks2MCTr+/86j4Yvacvhf1v
wK0OgIsa93/2BXZccZ6gb1VQxy7YcXMebZo91brAyNIGX7rMBchNStgom682kYIs
n5gAoN66raIa2Q3zp78HgZ3Y1Z+Hm2V7DJ6xs1PjTJwuvUZ1MRpW43UK3Yce7aEu
bjpRyQYlY6T1hZdPvUQ0qWRt/Lscl8qEjnKXmlv21GdOphc4jvaGxko1LtywZBW2
h/htpZTE7Gek60YZnoBS+jz4h5v88AquLrsxs3mcndPkeXSOGNbKLwMRHLWlyxP4
Y+RoqCtQ8c3UyIhNjkFEWjF3obZOjQqM+SQwLx5Jr+l8fSq9LiupdKWqLZy4kQS1
IeO8QxHAXg5fCPH4I8wC5NdFqA2Zso5j6OXu/ylrWUthjQ8cKr1CZRtubwM8j6sO
C5c1PiFWQPLpnuABkMmX0uMf+iLi/vrtx+kKbU4L76OtS1nHETwr0t/LT1XdtuN4
Iw3/Oji/k3fHB0Bi+qFX/1E20KDUyBdtf1jU57305gXQ4QlTGukdFCZqRt9sXSvy
K6xLFO1JkdBjEsOT/Tjpas2Dmy4oVOXoeEJjiTswwNvM4RhwIkBnXfA6bTdk9o7y
6eKFyzSTKlQnHhy27sLSPfJgy70gNUo8F4W/fvrq3RVBG6uexbos2nPNTBqOBak+
VxvrdFAuBRI6CPvev/L1Z4HqvNhCoi40eHljMaPQBEVFWiyVT+uebSW1HNv0jVdf
RaNkHk9mXFiwFEqRfqpIUsPOGp+On0Fz9/CJxFgbUQAicU6wm3uQPDnurI5DfSqC
9q6C3JHphDzcX5mfSo9c3jZ6joD3J5QJPpm919tmJn0GNy/Zv0v4QSG54Od1ovVt
BwruQdsNyT8MwVSwprE/Ht0uK/+rC/os0IY/FUpjgh0bhrax6YfevTuQZ0sQInTu
2+9zr48fCPPo3e3dq6NzXS0k/Fy9SrBpkrUHmTs+lekOhZe4EBcmxQ5xF9zk4YpO
gnY4J2/PjeI1yPIx3jp4RbEvBCXJOkc9aaa9bCsw64zpS66rkIlXs5FDxUhvppk3
16pWfaj2Ulg/apBrpKBSSxVYBlQOw4h0TByVHnIqB3+OHbO1gQ4RqLV3uqBtAibL
SMzFxeBFnyMwhbtjCKTS4lJpTe/KuGYr2iX/saLul2CAtBasccOHlmwQUlrlMnfe
CmP3K+P27wGRFVaT5UYzMkIiCt8rCV94oQ3WpRaVflXhlTrzqk2YIKlS4AS4nes9
Qfebv47kiypYUBjty7ftCrn+29sKcGsq4WNPDAh53xqdbZ93HsMUKGjdvcHnrOyu
xljkpBM0tUgERATd8k6ydXScPdCHfzIjXYsSTbLqrFsBZn64l+pxhePNYp5ADGo9
ZphjEVkaD23iRYk/va1SoG9VbU4Wn4HU0k0KKhSFuGQXEn3SHGUlnOyCiwmBa18z
nqse6hsAQBcI2tp+Q6oVPZE5C3bDSj5mZ0j3kogP4UgrqHKyN5zdtbvRDY6hiq61
NGC3q9gx9KP5D3rxD9BooGY3/6oKwRnIDakAADTysBgZz8jl27wnKFFMC6s52P1C
/OJHxCv8Pd93TmWbWhHoEcaiiwRnkc8SgxE423wiEjsu3mqzXd/BZ4ud4C2micVn
UW7QmpO1Se1b2CAxjVG7yUSaRULGEtUoXrCLrlAyZ393SgwMtVOinpEsnLUs1mDO
SlzimJFrHJ5G4yTqGxO5rKaimMbzeKQ/lYsPia16IxUz8ASTQMbfqzlBqjMEVk0I
XgiXti7Zk4UVvs99O5VkAWI2kOaISnhb2jN7usutMpFZCtw5M3vlRMYuFtdm8cie
L8R9jdy+5eHVGwtjuqICknNOMa5klm8oe1c0JPv6r2mlNRGMsG6sOXlZdFbuFd8p
7WxU6xsmaClHaALQCt9Iu91hLfVTdJr2XrewIQFDvXIOlBri0wc3/pEwrUO03bzO
aKbhyXgrmyAfbiU9gCkW1IvuV4lQvGT62PUUc2KEiwq+Xa2kWz0OO1hcVHlEq2ke
bWZfcDIky12OkrozlUUrJR9wTvaNMladfy1hD8v8QOzr6XDUIh/aiCH4sm6HsKHU
cxf+Sr0eXohOT2lwMI1yoElCyqJkhB+kJFtfT6fuZcPcGBIGKm/RcaXI5oC7IfBr
Aqb4+v9bUfxpeps9U647AmO2auFxu9EZJrvLjuqf8d/g9lE52iXR1O9dMl4nG2Xc
NkxHQiU5NhjC+67geRQLR6jbmn/dTJoLJ6giAKSz01Bva/4+pHHEL44H5U7VM4NS
knluiIaJ8rVW+9dE2lr3R2bwk0Rt24ps/aAtE8dRXwro/70gdq9Iudww5oLz97yo
ZKh8FpbsgWD4DWezUX6kg/6f0jTZcJj5gDP1GhBHhqyCokXHzpGVKMKUAWjSdDaO
b/4dycPr4yK4/bxlW6t6YMfyfxpp70q34LfshA+vmjU2sl+ELAxQGqN9Bq2Pe7XK
4ic6/DtumMVB9a8VEEtlTTd7PgYh6ZXYrWF51w4IHHAUWf8VwUU1lmGSFo+pDnVI
lqDIsmaQipc+qc5a7WE5OtLhCAZ36kaJlw0o6y5DLsxxFcs6yK9ChY80ZVYop/Lg
SskRuSClZ6rpvdvdXUR9GsZp2bVWY7xlbhF3cFdHZGwTsgbMQzxTGk0YK9UaeyaA
P3JuDCrtI9N4WnBM+Zv/8CwbyuEP31w2fgCHWe5pML6FX1KrWMCCyR4tobKAdbGW
pKMWiXT5APa76HbcJ4L58Ab8FkESwoQxi9vzVDP74wjtlC9ovYvNBiN2+sF9I+0C
PM4+SZlTjrCcs6U2fP3C6ZYR2kWGSjWYtMVWHEQrC3GDTo6+bWmsqUQaQQnecJa1
CpSSwldHAdx5CQosI+jj/U9soNA00ci1T4gsBUSNob3TZawvpczREGCwhBjZ4QZd
lN3gwQUIEvjvLK70v4ld9txwaofevqu29y3AQxpSoTbvtcg1l11Dfr/KZac8XZ49
JHXUxXiEfnEE4m9yY2Pet+3nQC6SCrPa8OiIs5nRlJs3Cn0HLveeQlaajj+nrWNX
UUNRjhCobUCotIX0sB0M6t0IMa5X6goAJ9VyQruiQLSiTfV52Sh2rU9iVCD8MhKa
q+qEY9gN6AvsOfx2xR9Dg1HOrRuqiFEmvoPiRAd60mkztMCZViKpsLnoi5u/MOLZ
RAQdUb2VMGr4+B9CC74ljnFDyl1HZaDSaQXznmS+ZEDJQqeCfUymL1gpPbYyDR8Z
6qgbpa5MF4GK5ON2Vh5Pfcuwe6MH/LmxJWiWo30c9DZQ0+dRMc2G6bqOhchqa9XY
Emby1trn0xw0EcbO0NqRXzKIXDNZHeW5NpKxj6nV354Gq0EPwRB0dszJYpwMdA/6
6u4qocwsEqWBVzUNhbj1c0VkLOok3S881oVESTcT/ypVAFtKC0dc2qsSoSMRueKE
9NX9acuJxrSirZRrwx1WwxCKwV43msog9IfXYuPZidIAik+22oRTNmoMxNSIVnD/
uarIGTxfe0m3h0k7wNn6ymA5zNrWtE8U2P2bITSBTjMd5c/vyVoMTy3pnmwKigg6
QvR9G5I3AyuvZhsLtWr/5psUzRU8sqNrLyBu9Gy4vusDwx3PWqpQiw7Ybgvx3T3W
HdkSlL7FHQDmxkPXUvbYpggUQuUmZ9kiENOlC6QHWgjg8MQF5Spwc1Mh5eOlXCq2
O8KggYSVlsG1szzJgQ6Aapf4x4i97G55+84DhsGJzS7wA3oJmyeHiZ/SqJMdzYgN
rON+KDcq7FsSeRj/e8Y5dwCSz8+tkADYR0tGumY736OJa5UDdRF2kES3mv/oU8ZE
BY2t2SAxXK8NL0Lyh5JYavTuTgxjws5dOeU2EHzbrW4zurIyrWwvpk0YxATa4uFW
vrVcbjnY3jmJiWQA7tur/WgxghDnjIIx1H2WquQFlU6wrrzA74f8/vb3eK0WzNb7
I8fnqKV7ne2DJ41ApWLKpOIB7VPsnBvkEcIg8A4kNFyx+nHba726tJLzHOVqDEp/
qJU8PH0Z5d/fXQiEjU6jMjjJq3yxA3sv8iUREk7NvtVV7vzYKGFnDrSOWIVrAap/
xegyIGOeaice2Ko/Q8Sw61vQDOemkdWMOTxrM7bXga0/HDX1RaCVi5v9+SkuCzMd
/bbj+nOYAfUEjk1ab4Ecjuema5PlcEabZCicP53gusN5FF6XjpQsPQOukNcj1E0y
rGswhEJWReMI+dvxbPuTeNJw8+V2XJBj0jnTLivcB8i0ecdh2D+rAIpYiFFRC+ov
pdFOf9iMbiGR3WZEueEmjNsMfvbPOzbF7LxsCQIpVzXC8qon/s256dHIvMJVH7mU
SkGiWqb10gOOxFhX76k2vacVE9tnxugdr6+rWtpVgS0e/gi6lyCTd88EPG3BwHmK
3PYXY3WM/4uqz+wa+fD49Y3sfeq3buyw3Kvn8ttaViAmQC1hP7AZqRwxhUYu832j
WoqexxheCyarKPvtvkZtGHrg7Dc5l4BPmoo8BDVIuuz0inrCzySfG//H32mjV+nn
NpMErbUOdqnRxl2mISAIl2JWXvB5P1xg/y6Cm5uGWkJ+zMglHUTxyGm7uJg9kr7N
oE0mLbTC9NK/bUxIY3Ly4+c1rBiLGTXQB6x9JYM+PaX0pd/nvCIqzuUUvKNwrhFr
/qpWCv5X+8WnWvKITgN7QgzuajlxM55XI2ZsHH9jKBMoMl6I9plgBuVCoOJ+gz2M
dGSEnhd1iJ4sMtf4zhlppCLNUbb1zJI4EjkJhiIUDEYhugB2KYRloXwDwJusIqje
7GZRgee0Ury3WEDi5Tc1ISHexHdZfyAjVEZ3qJ2FInJKEjRTzgUyeEa3EuNGOSdY
ugVnKCf70p5e0MaAJCAumpLOCU5FKlFxH9U343zK68yF60HdxJ+lpcSO+VbdnvHy
MA7OH43T3bb+sOWbEb9DX+f6rBEg1O8OThbm86jpGQWqAG+lxEG/+mBRx9ACy3MU
tzgPJOFR0UVOzhN9Rtl2dH9OpnP840KdF0d2B18HiyUQOvg1Ay+qjCgiOCS2uQu4
bOtwEQR4Ohi7rLiN7lrpIDHv2DtdnjjluZ8FCnUaD8VKV2HepvYNcKiniPvoqrII
lWks+NKiV4YQgQ2EtY8Iv5JXINIE6Xvf1+1IAeAnJkFbIYHSW1iuaQ9dPCXH7Bzf
5NiU82CnpAK3guBuIShViuudPrT5S1fOGUNgMHhxKjA64WrGXlInvK+PWXbGFp1a
92zFyZJWlbUWTdt8149jD0QHCentd6/JPjDCzxlEC+BMBUKHvMYQapT4J/i59iuO
SxSY3a3DCslPnpLE0TBSfVOKDiLR5m+UJ7j3hBdv+YrP9vptjsAKrBsntV0ckYrf
XSDEvtrJV6thSKGvh6t5rOx1L4VwQra42+VL8ndMpzhAiYaLWM0Fzosez4Otuitv
fjHC4KxEhKNwPBdtbEPixvwLYYmeZYSymQx0VwoVf6sghSUceJ/a8thTNXHlbuUm
tU3TBX7x3tYGZNDZTfJMVrw5nZSunMp+xZfPHT1NqVBZzx9HKKlNILzs+GeTmKmp
8364tQNy45oQY+naxgKn0zdzkER61fnTX+OgRNxb4oVw4B1JvbIOKY35XcE06WyJ
ZrvwRO6XhjCCCYVBTkhQAaXxK66XKKu6ROsIV50+CHK8H7XQ5Cxc+efeLZ2GEDNE
AjZnWJ3oeVw8T+ksj0C7bw3+ltwHHuqTj+Yp1qCPRJX3cCK06+NsOn3y7bGGOWqq
sY4ch79h2txb9hz/v8VlJ0QpdyWkqh1kkGozd1+lnPHYh3uqLjTlCFLXE57FQU3o
ikLynBaPxDwH5HDdfHhVRBc+oqT09s53UmvhOkWzZ7mxcutESZi0QWWFheDGUTsL
GNmjG8TxCfYn4wOp+8K2XukRXlCDKik+3j1ALFzAU9EgeUoleyLeJKQML6aGPT3k
FyK1042DTUWZPAe3zM1+gTYnEVKp4ejAzzNJCNjK57jWbw5+UhcjuoJ9WuXn60se
WTEuQthfiH83Ik1jLxvksk5C+jRfoycMQoKwZYawcY7YL6rPRXSnXpFqOcxzm/NN
5w58ivErkhXc9Grqv3gDOPABjB2EJGRps0QG4i1Q2h0ugD2TQZwQF6WWvYP8SFkN
zaLYCwJNj8dmM2o3PybnxDc7CMgbOjhgGwmkUVzkHu1qDVpW7DLilCqPWuo78CXj
ejZxLADvGIQBbywW8hNlgQg+X8D+lE/F9gj5ACh9Jtr9SExYj5FIG9yuUBV24bhr
56hyxo3K52OOXPRnwkbYxJP0K6wMgR1lAvco7VEHCMRbveXzFCTv7IsXONTLl7fF
HNVeGbXQ83lS5KIeXsDGw+9UB4Dts48M2coH9JMWmEm2rgxhDpPPdF/NsCKH5upQ
OXU5DbEuqpos2b/c/YwHfpA4cWoHOhXrCGb6hCKyP9iJZBIu+KYbVvSXphKnrhQB
K+XCFiJUfPwdbRLc5ELv6Zwn47fUirP8hkJGZ5pv9k1FixgicHLlnLwcBCr57+RT
oMiAMSvDqhEtJk3y4osh2Odw3odtHvXnLfBuAzFu5KsN7kv5alhLEZBypFWwlz+T
kCEutuEddnqdA4EHFIvOSiKrtuikpj9Sf+MY5uKi9RcI8jBO0lWW4z5xZsEOIVCb
/unZ4H3ZmUl2YY5UiISvAmKkqhxpZsMbki0SHXHjgW8gV4uaOiJEVsu9HBvXaqQj
SYed1MgkNylwtqxaJ9GMOH3uNEFKn/OpRrCkQ3u/DzAN0CUMOENQqOKSTpMuWgdF
EWmSXlMMSnM6aX9VyIgrojDBeuOMABoczcbLAPZVVrpP7bbsAUKcYXQzjbNo+JuV
ddzs4v/0pMt8exhpMtlBlllGsgXoxzEhd2I+2TtpmRAM/7g9wOakZqeb/r+P8HdA
Z3pngpjczH7eXYHsgXenvUDHU4JMDtKc/ge5vExH7JGRJ4g1sxh8nBD2c8+EjA8O
80Rd2C0iiSNXf46wz2Q0p1lplzVEIy6aPIvBuuXG8YORYKCKKYvz0eG46IEX052M
DoKmylmSOzleO1HHq7o4KMqW6t6PD+9gLmZOQtBfDQPM+FKX/+i3dPJb1QvDxmbu
BVD/Jm21jMds3O1lJ//9hZtiOrK/9TPENTfICcPeFSc+m54OcfXaQMPOOJtV5Z0f
bTOLZPMuW2aI2FGvkXz2S9mJ7cP04k6Wk0kgky6MaAMyDA7kRpze9ZuYwaho0PzU
Zfs1eONQWRCCAnZ2o76wHDhxGD/twf41n3P+7D1QrihpDowyTbCIn27t7ODmtYJN
Abzkj6icrHR4VraDwJWP2vkYzJ1k2chuQ6fSJuqZ3bYqewOcm4gkvOX22Ck+ID29
idIRqt7VAT3nqXVQLJKcW2DgWq7l6FqI0iXaTh8Gt/yA7ED5PBNh7VV34qrnYVZB
b0Tczu83kYAJmN4SS1VcMkF75PgTiGs8xKR10ztFPvq10kRfgBK4phgCnTPhpjqF
d7u6/9la70AIMNJWDNWOu98Q5j95N2VJrPnBaYTXp/0FJYtoUIggHvucSbPOPlJi
167WyTaa9wssYOCtH5J1M30pyDMkMirnr0sfYuEZrJNOmirQKcMJ4qqvXiXvwFUi
vBHabuX+TDosFRBgzyUZ/Ewv8BrWIQfNY17JE4w+LWW1l09i2C7pQVD2zdWNadtn
tAvouUIE7gRj+TLGDHUtQEI/t2j206ciampRsnkW45x4woZ8sX3zmoKs9uMEAVNB
uzH3RMy1U6skcTLSymC9RoPfIjdW2HdqDYOUBHh+N3DKJHcvzh3nKIhhI4Ik8nih
Lny4XB/dqMD/Zmdew28m5upypowA5xA0jZxl0UigFkLESF/OVjz66h9TKykIIS7O
u/LZW70VOXpCzDmOHl+gkTw4C+YiIZybEPuE1L+ZWxuhOnk3S99rxLs1m/Tjz1Bu
DAEc41Lv0T8l/IbACh8OGj/BJb0fxN0qFT6mCsLIZvZHznAvvrz0ZMxAKb6fsLtU
+4d+bF55mKkoSHgcoxNGBmQf2LEjp5/fmCrdY7VH+dUrkfLXq45jDv+JT2HtpY20
nWAdTfa7pBf1fe5wtd+Ych3ngaFNOdqlh4yT7Svfe01O3Y/XUnr5ERGzjMBk311H
JRfON61y9S/mq5YGvUentP3zs1TRQ8RNAu3nZo5KRGV1GgFs+Zzl8vCEOd72lqhu
Fmr9O/VtWUZpt83YpNW2ttn3uzBRCSsFNx9m5rdhTMnIwjTFNQP02zwH9c1gUXDM
mwrweiNxLv/WIQr2swZiFSDzmdt5ahlUAeTe8tQIRhTzzfFgDnhNHWkv8YwQq/hg
+C0JL84THSxez8Qdib1TMi5pY9TAZHT4iXnJcQcAGAIU47eaLFAiU4e3zcPndnLs
LODdzvDWW8KPHSZkVnift8Zt6PvqDFVfV3fnkOKifdqKy0Qt8Gh+tqwYcmSX0XFN
Dpi5JhzZ1w4z+ADGyBxELCGMncN7hwZPFBuzDN81xdbVXmekyaeqiwEw2vzLV0qZ
X8Q0fiA4L65NmUVUlihJKka48leZIF4vgtdxpvPmVHcnuvl27uBuRE0Z9alsbkD4
4Vd4Zv8cR7blz9D9RmuMi6Ae1yDsFWJo0GoS0IUqb52GYQXgoToJjJbZoVbfIAfE
zcYZOKbai8C14Ex0btclPOzxHjVYUuKLTvb1O17gYMLsqAMoiODKZC8RNgFezCBZ
VhqdcIDXZdiiUkAncvOZ8TgFHPSu8ff+PDIMJTk0aFv/fV9RFP0kZZvTdKaENJQE
3sywzZjBBMepFpV4xTinkkcneHG0QlaIb5wVvSsYlTbaPf99DIsEi8FT6Mzqh/9c
XeTjsbPVz2gKVKU9aC/eeqcL8PscHlK7cltoTrjck21vE091itij40oEndOETyG3
srbdnm/41jJqwCwnhOHuHiiBqZzfMjVuva1Ke/7FJlhgWqbE5bqBU6Ph/YFJPc5f
KLDB2Y6b+s9NtyXg6Z+RLMfL9hr5pDdYdMP/L+wlCiLNT+yu6+El0cbSEpyeGyXe
k0w0FrRS2OyBlCdfyhsQueZDqM8yw4TCHzQp8Z9TTdsbEmP1onw6Y1wTMcm1Sny4
lbXkNixfDoTqYtGgYXYNv+IyX/DupetH0SgEMmA6IUjFKWAS6kv1YG2cLj7ZTtJp
B+buIYH/leegz1xfmD0p2ChIcnnMOUvE1pIHexgveuFeO9ASHL89jpPLve/CTLhU
d+vy+rRc5udyMk8QhudIQxjgEiXjaE2Bb1l7qMQt2Uk2RJ82oWJzCOhZBYtucJqf
RBgUKLKxkdN//OheiygkYy26XSl2f2MjW1m4EFTc2QFlgPwHJQM4hqXsoltFErW1
Fp2d3O+ymmEm9IvPJgYOWkA33n86apZ2aYTSveuWxI9hxj++Z4ZN5tNmuO3pfXMe
BrPT0RIiIBeKCEM72IBVNEihiJANvqcyFTWGCM4s1kvaZtEvulHxBdcEoagTYelQ
oH7/BIDG9FYq1OvA7ZnZ/8gAyAdGiRN8Op4GEN6iq7bW8EkyubtHbPgyb6Epjgy5
jC+EIXf2ZisBraJ+Vs9zfBMc0LaVsFLzTrkKwuj8/Cw9JflKojqZKt+epMpdyETz
c/obgJZ9bN0M0iTt9NeSAayaL3M9S/E/S14VjRgNXiDZrhkSKcaLfWf4NnJuI4O1
HXbftyFdoED0x39BfDjWmd3zLVCcxDfucU9nrahCSgaN0d1pptrCUH0H1cBb9nqe
TOYUTs7fo8mbTAo30A53C4BRK7C+YMnHbhBOZ03gGF76ie7vXoai4Ffw3wF6daKe
x2gSg1F0TKPek5z9rh/E40GBrtfwD5CuopSPxFCN8AkH8VjKghtfeDifklktPegI
4fwcDUSzCqmrc24dOWleR/yqYORmXKJtgMJjZLM84Jyp7PQ52xa0DZgi9X7Aoarr
wgoShHdCHXNXDB3yLwYyTuAjf5YJL1Q3zbh7Gnuj562teIBMe7KkUUV0CsKVDTu3
TTTkc4BYlSrSC/sqigPt/j/yDwcrqWX2R1hoyUAw9CHODQHEyc6qOFeABgCIAIgB
/n5UpNEFYqH3DjZ6Mxd4uP7k+muckrM4WufUvqvsiqXjVH6wmXO1uAb9w+KIk+Dj
6KvYMlfLvo9bVi0JW0Unuf9Pbz6rog4NYdhFyCAk8EVg/lauB6oLwHdMLyaHgQ1l
JHVmMZ2akRxobgCdbkF+PobtS5uHAHdB5viUqm0/k75i4M1NbFNF6ChTg2/1iU0H
K4GhCQWzBUPlrMcRDIBBKFK/ZF69NI6TKCmX1aPpuEeQ3d0/bO46sgLI9WcwJLuw
/LJ8bV03aB0jH6/jGD+XPSL0hc2vHOQuVbTLMHvG9hniZ1UCYYnj+OS8cKX+uDYE
EkShunMBoMdsYhj+gy7d+xd+MKPSkjPBdNDX9cfb8WLgwP+9BBPgGcoALk/6h2os
t8OuNMyp27KyQfuQ6UbIvZNk+9iU4MkjdW/aeJHTC+y4wfUBr8uCz4A2R76kowef
lmlrKWqS7YNb5QZ7OD4kKYfFF0BiPk5Wxder2Zs85rfTNZlNYxUjuN+Uiqiagmtp
WnejsMz4tWzAJM6w6hVVWztUtlWweHjHigp85NuZoNyPnz+G6qvNgnZeO2yxCkBn
ocSKS9tymQ/S6ezXfGEdwphzHw6uk5aA1YHgR3AGiBuMy3dyIuG7SG9r/KZgSjL+
CfAsrbZuQHcC5nYpI0y7i1kxQ9g35tnwAaW2lJPSDCbuV3GixakP8M2vIyVBYRTP
PtZoQMup7yIed4r1AMUXK0d7IWCsqIN0XKe8p1AYIAFGLWSYrzfnCD5/6wHHqM1K
CMXHVQYjvHuOBU+AEVmaHxx9/REE2Y0uqOk4BcbdCNnOUrBVrxRTv/jwIPW3rPcR
Esf4cQPEX/3P+yIvC/qBubw3nf/ZrpRNKf5n7Hiiko7nAMTi4iGJ8QfHBYa0n6SX
BhDghCjMgDfFb6PZQAz9b2ksexrc8SanE7ilK3o+lUJ9RGucKWIwTjToshRnZDr6
5C4Ng1y/BRyZAQkwCdKYGyfOzJwGASO5s8f3m1Xpgg7KqTOUEiNDLV/9Fvltutml
Z1tJLpJHSBEkiiNnKn4H9r6pcaNjoV2MZCn+jQ0T3YelTQFcQiJ5Pw8W+xqpOsMJ
ifJLmYbDKUMi5ecOj57uytTx+j3MCX3R9X1bE1bSdAsIQ39XZX8f+b/1PN6snAfD
ToLUVWHwmSAV6EeHUoJgnzqz7h1bsUh04Lc1Gm1veBoNmm0GNKm11AvRVkZSkRt9
G0IHQMLLyJUYZL4IP2tvJydY1vptK3IpkBkH00Z7C4tsOleBgqggSEKF/alGkUBV
Frv6BK6VtoUFAu3zqIQD7jD1oRiYpi8YwjP6/D5E+QNaYROMmZBirpIICGPENDpZ
bi0JC0WX6AIEGI085kG6Teo/yVl83lid52BSgvTZoK8CgiXE3MIqEL9MNN5apHDa
7RHv+RZZuJ1Ki45wIN01s1qhvJerNzcKt555ndSChHm756uoa1uaPkCURp0fAo2R
MOa58J5sQivAT71VNAl6H6Q71qRva4ZSBiAnDwA1Wn3eZt6FY72xlFZoUOYLcvSi
hLNcL7V3SSvrJwJRPsZ2gHjMS8OyuJMUYq+oz8I+ejmjCPE5WAo+10jbIpqXIXPA
MRH9FFR1QvOsTrcHOW+AAzDGQxbcBsoqA0x4PEEYKniuoI2srYbUJj0s7RLtGUrs
TzHZi6IgGFum2fmk1qIDKn/BFVc2ACaJKS3WPg5/7v6YjVb7q/Fz9K1iu/EANNcq
2fXy+dAsHWHwVzTYNMb9UtJr/KIkov1d0th7hqYbhF+fgaAlOt+fX1tov/hBGYUg
4Qf+yd6FLCevYvsrYbgg7ho8Pjxbw/5CUquOObVEs6Fk2vhY+X53SsXjftY89H4w
ATMdkBz2z+puhJgPWff5i+rzEstdKS6RCAX60TzsEmVQonJpSUr4k51/pcUlgTVG
SQQLDzZR0kTitJgDw72XA2dJAx/ZnPzRSFFrTV5/YPG4IuKH7vdXD1NNgI0ofBcT
fzJP5L+npnQVtQE3Jd5dcqk81FcfuizhZxxVOigro1eFq6gzzn0gyFikZH6sBJi9
GATcFUnvHr1DqtZ2CBj8dmVrXU7aq7+oObdCSqYVzLvHiprCbmHFDB/A1IXkNR6w
R7QaHkN6EgJcZlpr3e4s+jGO2KNjWNgtDhvk7U7h698JpJHRKyO390Btw6UJZXBY
YFtXWj6PWObUzvH7bTEtUc9avtfRytR4Jk8h+YrZLfYhBMUaMU+60U38GWe+c2eo
7ZcE+dRU7uqw6fDE31huTg+Zqo5ejQqxBzCrmn2F93Yoez0pLp+zTs3nh7SQvInq
hEUwfGjwZWGQTi3BT4B8O3A2/3xzAMyI/u7dRmFYQLQvyR1F97+ulXh8GZCd8LGz
peQBp0L3qtQsg/60m8JQVNyOscOB0dyh/i1usE0xuP6q9/7jab1qCCUms77nKWec
dOQND4wI/FpBSJrtl+BUaghEg6YEMlUZJlF9O1T645RnXec6OCWQi0jbS25j5Cq3
hirFerX4Yiucow2VAWk+BBkdJKdyKJ/f3kGAb8CNaxBU+FtKFh0vPFM1/+ga1ue9
zdIjLb7PLltn52T6W3Y5hw4PKyHOlY7gOW4BCJcGycs+HZL09J3GQ2oJ3fgEMbnv
24lFJ8jthiPig0IysXoK+c2Iu4n+hR5iedQWrHUHzOPTA+PpTP8gJ7UUe9oI9mUt
bOYyVXCDmIhgyZe/Dz3mnkvOvYsQYL93okEtjvdz+Ht0XJdcNWZQLK2+5Chs6pYd
v+zLDdDZ9O1CsmLgQhN4OL1xchqY0GExfMB2WjnfMjN1h3Gjcafe6bkZHEGQ6lCk
ns0BZpRClXAL2gToqx/7bgwxJHuJC44B5BaTn7mBXWNh/azwM+EsF0iTG9ibQyUb
saogh3SV+564gRfTOwVf7pSAIVwTdmaPBl/qMnL+2vjqY0z7nRpXUyOm0I+0W2kf
UvdRse8kz7+SLAL6+v0+R/ue0Gnj0ujSFIbvc5LPLf1ubOaJ3tZ5oJJbik2Zm/Jk
KS3W+qhcYYgk0+QjKRr8AVfICZlMHyPMgW+DyhMo7TXRpug33NgkXyUQsoAjYqsT
qvfW1ypy1lnIyjmBKw7KFrkvK3RKlRdhjikn3NBfhaAZqNQOq3Jl3BKM3fJxyI4L
UlA3VwARsJ7A0n0hxuPcVqmtuIZGFmGz1fQ5KanSdxXrH7hcBnNDNPnU7TFM8pHJ
ikGjxUz4VxwD/MzKKEVhGUtSfFyTY6zP4JuwwfZgej9vDFKw0vGbsf/uil3yewwV
up72vmNJ2nga235W94sxMv5gaeKZgGnoZyvlmwWJeCUWrw1NoY2HCknraNuFdKST
tKKrhew0YUizT7KEXsKcOw+woU9vsOk/9HSZWP5KdCs7P9ua7NphsYn7O/EiAgR0
MGHfDYfgYJnnDHaIJGBHJR5+dHh8SRzA0BWoMUCgxpVZy5F//TkMxQanmyb/a8UB
rC1sUhHJwX1JBep9at9LT760C3cJEs0Dci/6XrFHIdpxZCXY1XN8xp0IHJglYVhA
6pcK1cDpYNomLQ7VzpmcIng85Tf4oaw3WyIo7hAyPA/1Ox1LeYZ1yF+Xzq2Glvt2
x7XcJ01MByorwqWvy14peSyi2Im0V+MU8/DIYNtqHytBWyfhU8Q4g9pla87JdNi3
WCcFDemAhfEhkoEihFB7uftk8RXjGvLGRo3HSGLs5pAtnu7vF40Fp/zjucjQ0vI0
A+tzF3Vunr3eW7dWxzE2456Q2W5Bc51xPYqZAm3FQSRFR3jy9J0LY9K90X3feV1J
8pI9fz2HWJOrPO6EzjB68SXzbZnNpK+UqggOs7b8IEwKQUlkeINw5yjTUSyBH/+I
b9qImfBrwwUwTU1lT2+YBvonJHGArsLw95BsYTyfXtOsOECdLlGen3Ndf7zkth4M
S//wIOr73rYmCmamaUk/tOvyebDkzq/85tJcIs24t8HksHRf+eDR2DJ1szqa4OCF
Ji/d/SfX5e9KE74t5xs46Xh87Upj5cGiCZbmKiD77uIEC2ok90P8koKfkJ+WAMyq
o2PtLidgV8br+d978vGHecev6/uMMnKOX6b97Yl9tszErkk0mFqoA6ICh3ULFsun
DCcXKY79tFOKllAzI0NsVz/u2v5ndePhCfEgITwxRbyC5lfdDKh0f7VMh8rt1PWU
Q+v/HK+XJkLrdZgB51juOLRVgF72ZPfgMdUcuk+KwzGAasUnWw+ixG521gtCxuQZ
8paTHpm34AFX/i+bjlNLSAEiyPGUHpm7X0mWg1dw2nZy6u0NzVfkTCTqoXocEM3E
d1FkynB8/CP9AEYqPbhSZcScd96JHmjqvafHIqFt27zKc5Snn2AKHCp+CNsqxN9m
8bWRZ54OzU5ptAmIWUh/mR77CxgoLd2mJ5+zy9NA2X6oRa3mQi6gh7Y0SvH91UlH
5Vx3RmTRMyQM0NeH9sYxARolPI2f/cigZHCfzObVhbE0uJ9lW1A+53LO4S6C8nBR
2zXR78B5XvTZo7c+Zmuvx0HkG3NpJ26GCgeCDc6RiJObC0BnSN15bpmeRL65qtmE
UCKl5F7GKrPlgFNNOTgTNTyk77vY1i3cMKVjXU6v3VqAdNsPzBMEYYWC6VUrXJTH
PgMD6TiwKq8oBiSjXLS3uIRkPk2EFbO1/CjqtubJZU64PB93lwyTCE7rrxseJZnP
LGsB+vYYhpKQnn3X8w90nCmN42hDAwjW23i0+tLcARQ=
`protect END_PROTECTED
