library verilog;
use verilog.vl_types.all;
entity twentynm_hssi_gen3_x8_pcie_hip is
    generic(
        enable_debug_info: string  := "true";
        acknack_base    : vl_logic_vector(0 to 12) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        acknack_set     : string  := "false";
        advance_error_reporting: string  := "disable";
        app_interface_width: string  := "avst_64bit";
        arb_upfc_30us_counter: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        arb_upfc_30us_en: string  := "enable";
        aspm_config_management: string  := "true";
        aspm_patch_disable: string  := "enable_both";
        ast_width_rx    : string  := "rx_64";
        ast_width_tx    : string  := "tx_64";
        atomic_malformed: string  := "false";
        atomic_op_completer_32bit: string  := "false";
        atomic_op_completer_64bit: string  := "false";
        atomic_op_routing: string  := "false";
        auto_msg_drop_enable: string  := "false";
        avmm_cvp_inter_sel_csr_ctrl: string  := "disable";
        avmm_dprio_broadcast_en_csr_ctrl: string  := "disable";
        avmm_force_inter_sel_csr_ctrl: string  := "disable";
        avmm_power_iso_en_csr_ctrl: string  := "disable";
        bar0_size_mask  : vl_logic_vector(0 to 27) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        bar0_type       : string  := "bar0_64bit_prefetch_mem";
        bar1_size_mask  : vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar1_type       : string  := "bar1_disable";
        bar2_size_mask  : vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar2_type       : string  := "bar2_disable";
        bar3_size_mask  : vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar3_type       : string  := "bar3_disable";
        bar4_size_mask  : vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar4_type       : string  := "bar4_disable";
        bar5_size_mask  : vl_logic_vector(0 to 27) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bar5_type       : string  := "bar5_disable";
        base_counter_sel: string  := "count_clk_62p5";
        bist_memory_settings: vl_logic_vector(0 to 83) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bridge_port_ssid_support: string  := "false";
        bridge_port_vga_enable: string  := "false";
        bypass_cdc      : string  := "false";
        bypass_clk_switch: string  := "false";
        bypass_tl       : string  := "false";
        capab_rate_rxcfg_en: string  := "disable";
        cas_completer_128bit: string  := "false";
        cdc_clk_relation: string  := "plesiochronous";
        cdc_dummy_insert_limit: vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi1, Hi1);
        cfg_parchk_ena  : string  := "disable";
        cfgbp_req_recov_disable: string  := "false";
        class_code      : vl_logic_vector(0 to 23) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        clock_pwr_management: string  := "false";
        completion_timeout: string  := "abcd";
        core_clk_divider: string  := "div_1";
        core_clk_freq_mhz: string  := "core_clk_250mhz";
        core_clk_out_sel: string  := "core_clk_out_div_1";
        core_clk_sel    : string  := "pld_clk";
        core_clk_source : string  := "pll_fixed_clk";
        cseb_bar_match_checking: string  := "enable";
        cseb_config_bypass: string  := "disable";
        cseb_cpl_status_during_cvp: string  := "completer_abort";
        cseb_cpl_tag_checking: string  := "enable";
        cseb_disable_auto_crs: string  := "false";
        cseb_extend_pci : string  := "false";
        cseb_extend_pcie: string  := "false";
        cseb_min_error_checking: string  := "false";
        cseb_route_to_avl_rx_st: string  := "cseb";
        cseb_temp_busy_crs: string  := "completer_abort_tmp_busy";
        cvp_clk_reset   : string  := "false";
        cvp_data_compressed: string  := "false";
        cvp_data_encrypted: string  := "false";
        cvp_enable      : string  := "cvp_dis";
        cvp_mode_reset  : string  := "false";
        cvp_rate_sel    : string  := "full_rate";
        d0_pme          : string  := "false";
        d1_pme          : string  := "false";
        d1_support      : string  := "false";
        d2_pme          : string  := "false";
        d2_support      : string  := "false";
        d3_cold_pme     : string  := "false";
        d3_hot_pme      : string  := "false";
        data_pack_rx    : string  := "disable";
        deemphasis_enable: string  := "false";
        deskew_comma    : string  := "skp_eieos_deskw";
        device_id       : vl_logic_vector(0 to 15) := (Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        device_number   : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        device_specific_init: string  := "false";
        dft_clock_obsrv_en: string  := "disable";
        dft_clock_obsrv_sel: string  := "dft_pclk";
        diffclock_nfts_count: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        dis_cplovf      : string  := "disable";
        dis_paritychk   : string  := "enable";
        disable_link_x2_support: string  := "false";
        disable_snoop_packet: string  := "false";
        dl_tx_check_parity_edb: string  := "disable";
        dll_active_report_support: string  := "false";
        early_dl_up     : string  := "true";
        ecrc_check_capable: string  := "true";
        ecrc_gen_capable: string  := "true";
        egress_block_err_report_ena: string  := "false";
        ei_delay_powerdown_count: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        eie_before_nfts_count: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        electromech_interlock: string  := "false";
        en_ieiupdatefc  : string  := "false";
        en_lane_errchk  : string  := "false";
        en_phystatus_dly: string  := "false";
        ena_ido_cpl     : string  := "false";
        ena_ido_req     : string  := "false";
        enable_adapter_half_rate_mode: string  := "false";
        enable_ch01_pclk_out: string  := "pclk_ch0";
        enable_ch0_pclk_out: string  := "pclk_ch01";
        enable_completion_timeout_disable: string  := "true";
        enable_directed_spd_chng: string  := "false";
        enable_function_msix_support: string  := "true";
        enable_l0s_aspm : string  := "false";
        enable_l1_aspm  : string  := "false";
        enable_rx_buffer_checking: string  := "false";
        enable_rx_reordering: string  := "true";
        enable_slot_register: string  := "false";
        endpoint_l0_latency: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        endpoint_l1_latency: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        eql_rq_int_en_number: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        errmgt_fcpe_patch_dis: string  := "enable";
        errmgt_fep_patch_dis: string  := "enable";
        expansion_base_address_register: integer := 0;
        extend_tag_field: string  := "false";
        extended_format_field: string  := "true";
        extended_tag_reset: string  := "false";
        fc_init_timer   : vl_logic_vector(0 to 10) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        flow_control_timeout_count: vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        flow_control_update_count: vl_logic_vector(0 to 4) := (Hi1, Hi1, Hi1, Hi1, Hi0);
        flr_capability  : string  := "true";
        force_dis_to_det: string  := "false";
        force_gen1_dis  : string  := "false";
        force_tx_coeff_preset_lpbk: string  := "false";
        frame_err_patch_dis: string  := "enable";
        func_mode       : string  := "disable";
        g3_bypass_equlz : string  := "false";
        g3_coeff_done_tmout: string  := "enable";
        g3_deskew_char  : string  := "default_sdsos";
        g3_dis_be_frm_err: string  := "false";
        g3_dn_rx_hint_eqlz_0: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        g3_dn_rx_hint_eqlz_1: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        g3_dn_rx_hint_eqlz_2: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        g3_dn_rx_hint_eqlz_3: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        g3_dn_rx_hint_eqlz_4: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        g3_dn_rx_hint_eqlz_5: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        g3_dn_rx_hint_eqlz_6: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        g3_dn_rx_hint_eqlz_7: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        g3_dn_tx_preset_eqlz_0: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        g3_dn_tx_preset_eqlz_1: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        g3_dn_tx_preset_eqlz_2: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        g3_dn_tx_preset_eqlz_3: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        g3_dn_tx_preset_eqlz_4: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        g3_dn_tx_preset_eqlz_5: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        g3_dn_tx_preset_eqlz_6: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        g3_dn_tx_preset_eqlz_7: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        g3_force_ber_max: string  := "false";
        g3_force_ber_min: string  := "false";
        g3_lnk_trn_rx_ts: string  := "false";
        g3_ltssm_eq_dbg : string  := "false";
        g3_ltssm_rec_dbg: string  := "false";
        g3_pause_ltssm_rec_en: string  := "disable";
        g3_quiesce_guarant: string  := "false";
        g3_redo_equlz_dis: string  := "false";
        g3_redo_equlz_en: string  := "false";
        g3_up_rx_hint_eqlz_0: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        g3_up_rx_hint_eqlz_1: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        g3_up_rx_hint_eqlz_2: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        g3_up_rx_hint_eqlz_3: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        g3_up_rx_hint_eqlz_4: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        g3_up_rx_hint_eqlz_5: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        g3_up_rx_hint_eqlz_6: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        g3_up_rx_hint_eqlz_7: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        g3_up_tx_preset_eqlz_0: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        g3_up_tx_preset_eqlz_1: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        g3_up_tx_preset_eqlz_2: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        g3_up_tx_preset_eqlz_3: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        g3_up_tx_preset_eqlz_4: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        g3_up_tx_preset_eqlz_5: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        g3_up_tx_preset_eqlz_6: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        g3_up_tx_preset_eqlz_7: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        gen123_lane_rate_mode: string  := "gen1_rate";
        gen2_diffclock_nfts_count: vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        gen2_pma_pll_usage: string  := "not_applicaple";
        gen2_sameclock_nfts_count: vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_1    : vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        gen3_coeff_10   : vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1);
        gen3_coeff_10_ber_meas: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        gen3_coeff_10_nxtber_less: vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_10_nxtber_more: vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi1, Hi0);
        gen3_coeff_10_preset_hint: vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi1);
        gen3_coeff_10_reqber: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi0, Hi0);
        gen3_coeff_10_sel: string  := "preset_10";
        gen3_coeff_11   : vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1);
        gen3_coeff_11_ber_meas: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        gen3_coeff_11_nxtber_less: vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_11_nxtber_more: vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_11_preset_hint: vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0);
        gen3_coeff_11_reqber: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi0, Hi0);
        gen3_coeff_11_sel: string  := "preset_11";
        gen3_coeff_12   : vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1);
        gen3_coeff_12_ber_meas: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        gen3_coeff_12_nxtber_less: vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_12_nxtber_more: vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_12_preset_hint: vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        gen3_coeff_12_reqber: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi0, Hi0);
        gen3_coeff_12_sel: string  := "preset_12";
        gen3_coeff_13   : vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        gen3_coeff_13_ber_meas: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        gen3_coeff_13_nxtber_less: vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi0, Hi1);
        gen3_coeff_13_nxtber_more: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi1);
        gen3_coeff_13_preset_hint: vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0);
        gen3_coeff_13_reqber: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi0, Hi0);
        gen3_coeff_13_sel: string  := "preset_13";
        gen3_coeff_14   : vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        gen3_coeff_14_ber_meas: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        gen3_coeff_14_nxtber_less: vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_14_nxtber_more: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi0);
        gen3_coeff_14_preset_hint: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        gen3_coeff_14_reqber: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi0, Hi0);
        gen3_coeff_14_sel: string  := "preset_14";
        gen3_coeff_15   : vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_15_ber_meas: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        gen3_coeff_15_nxtber_less: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_15_nxtber_more: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_15_preset_hint: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        gen3_coeff_15_reqber: vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_15_sel: string  := "coeff_15";
        gen3_coeff_16   : vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_16_ber_meas: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_16_nxtber_less: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_16_nxtber_more: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_16_preset_hint: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        gen3_coeff_16_reqber: vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_16_sel: string  := "coeff_16";
        gen3_coeff_17   : vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_17_ber_meas: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_17_nxtber_less: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_17_nxtber_more: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_17_preset_hint: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        gen3_coeff_17_reqber: vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_17_sel: string  := "coeff_17";
        gen3_coeff_18   : vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_18_ber_meas: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_18_nxtber_less: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_18_nxtber_more: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_18_preset_hint: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        gen3_coeff_18_reqber: vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_18_sel: string  := "coeff_18";
        gen3_coeff_19   : vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_19_ber_meas: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_19_nxtber_less: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_19_nxtber_more: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_19_preset_hint: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        gen3_coeff_19_reqber: vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_19_sel: string  := "coeff_19";
        gen3_coeff_1_ber_meas: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        gen3_coeff_1_nxtber_less: vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi0, Hi0);
        gen3_coeff_1_nxtber_more: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi0);
        gen3_coeff_1_preset_hint: vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        gen3_coeff_1_reqber: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi0, Hi0);
        gen3_coeff_1_sel: string  := "preset_1";
        gen3_coeff_2    : vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        gen3_coeff_20   : vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_20_ber_meas: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_20_nxtber_less: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_20_nxtber_more: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_20_preset_hint: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        gen3_coeff_20_reqber: vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_20_sel: string  := "coeff_20";
        gen3_coeff_21   : vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_21_ber_meas: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_21_nxtber_less: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_21_nxtber_more: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_21_preset_hint: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        gen3_coeff_21_reqber: vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_21_sel: string  := "coeff_21";
        gen3_coeff_22   : vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_22_ber_meas: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_22_nxtber_less: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_22_nxtber_more: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_22_preset_hint: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        gen3_coeff_22_reqber: vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_22_sel: string  := "coeff_22";
        gen3_coeff_23   : vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_23_ber_meas: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_23_nxtber_less: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_23_nxtber_more: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_23_preset_hint: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        gen3_coeff_23_reqber: vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_23_sel: string  := "coeff_23";
        gen3_coeff_24   : vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_24_ber_meas: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_24_nxtber_less: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_24_nxtber_more: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_24_preset_hint: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        gen3_coeff_24_reqber: vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_24_sel: string  := "coeff_24";
        gen3_coeff_2_ber_meas: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        gen3_coeff_2_nxtber_less: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi0);
        gen3_coeff_2_nxtber_more: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        gen3_coeff_2_preset_hint: vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0);
        gen3_coeff_2_reqber: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi0, Hi0);
        gen3_coeff_2_sel: string  := "preset_2";
        gen3_coeff_3    : vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        gen3_coeff_3_ber_meas: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        gen3_coeff_3_nxtber_less: vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_3_nxtber_more: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi1);
        gen3_coeff_3_preset_hint: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        gen3_coeff_3_reqber: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi0, Hi0);
        gen3_coeff_3_sel: string  := "preset_3";
        gen3_coeff_4    : vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_4_ber_meas: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        gen3_coeff_4_nxtber_less: vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_4_nxtber_more: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        gen3_coeff_4_preset_hint: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        gen3_coeff_4_reqber: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi0, Hi0);
        gen3_coeff_4_sel: string  := "preset_4";
        gen3_coeff_5    : vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_5_ber_meas: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        gen3_coeff_5_nxtber_less: vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_5_nxtber_more: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi1);
        gen3_coeff_5_preset_hint: vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0);
        gen3_coeff_5_reqber: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi0, Hi0);
        gen3_coeff_5_sel: string  := "preset_5";
        gen3_coeff_6    : vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1);
        gen3_coeff_6_ber_meas: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        gen3_coeff_6_nxtber_less: vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_6_nxtber_more: vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi1, Hi1);
        gen3_coeff_6_preset_hint: vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0);
        gen3_coeff_6_reqber: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi0, Hi0);
        gen3_coeff_6_sel: string  := "preset_6";
        gen3_coeff_7    : vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        gen3_coeff_7_ber_meas: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        gen3_coeff_7_nxtber_less: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi1);
        gen3_coeff_7_nxtber_more: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        gen3_coeff_7_preset_hint: vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        gen3_coeff_7_reqber: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi0, Hi0);
        gen3_coeff_7_sel: string  := "preset_7";
        gen3_coeff_8    : vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_8_ber_meas: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        gen3_coeff_8_nxtber_less: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        gen3_coeff_8_nxtber_more: vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi0, Hi0);
        gen3_coeff_8_preset_hint: vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        gen3_coeff_8_reqber: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi0, Hi0);
        gen3_coeff_8_sel: string  := "preset_8";
        gen3_coeff_9    : vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_coeff_9_ber_meas: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        gen3_coeff_9_nxtber_less: vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi1, Hi1);
        gen3_coeff_9_nxtber_more: vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi0, Hi1);
        gen3_coeff_9_preset_hint: vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi1);
        gen3_coeff_9_reqber: vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi0, Hi0);
        gen3_coeff_9_sel: string  := "preset_9";
        gen3_coeff_delay_count: vl_logic_vector(0 to 6) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1);
        gen3_coeff_errchk: string  := "enable";
        gen3_dcbal_en   : string  := "true";
        gen3_diffclock_nfts_count: vl_logic_vector(0 to 7) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_force_local_coeff: string  := "false";
        gen3_full_swing : vl_logic_vector(0 to 5) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        gen3_half_swing : string  := "false";
        gen3_low_freq   : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        gen3_paritychk  : string  := "enable";
        gen3_pl_framing_err_dis: string  := "enable";
        gen3_preset_coeff_1: vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        gen3_preset_coeff_10: vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_preset_coeff_11: vl_logic_vector(0 to 17) := (Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_preset_coeff_2: vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1);
        gen3_preset_coeff_3: vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1);
        gen3_preset_coeff_4: vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        gen3_preset_coeff_5: vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_preset_coeff_6: vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_preset_coeff_7: vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_preset_coeff_8: vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1);
        gen3_preset_coeff_9: vl_logic_vector(0 to 17) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        gen3_reset_eieos_cnt_bit: string  := "false";
        gen3_rxfreqlock_counter: vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_sameclock_nfts_count: vl_logic_vector(0 to 7) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        gen3_scrdscr_bypass: string  := "false";
        gen3_skip_ph2_ph3: string  := "false";
        hard_reset_bypass: string  := "false";
        hard_rst_sig_chnl_en: string  := "disable_hrc_sig";
        hard_rst_tx_pll_rst_chnl_en: string  := "disable_hrc_txpll_rst";
        hip_ac_pwr_clk_freq_in_hz: vl_logic_vector(0 to 29) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hip_ac_pwr_uw_per_mhz: vl_logic_vector(0 to 29) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hip_base_address: vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hip_clock_dis   : string  := "enable_hip_clk";
        hip_hard_reset  : string  := "enable";
        hip_pcs_sig_chnl_en: string  := "disable_hip_pcs_sig";
        hot_plug_support: vl_logic_vector(0 to 6) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hrc_chnl_txpll_master_cgb_rst_select: string  := "disable_master_cgb_sel";
        hrdrstctrl_en   : string  := "hrdrstctrl_dis";
        iei_enable_settings: string  := "gen3gen2_infei_infsd_gen1_infei_sd";
        indicator       : vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        intel_id_access : string  := "false";
        interrupt_pin   : string  := "inta";
        io_window_addr_width: string  := "window_32_bit";
        jtag_id         : vl_logic_vector(0 to 127) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ko_compl_data   : vl_logic_vector(0 to 11) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ko_compl_header : vl_logic_vector(0 to 11) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        l01_entry_latency: vl_logic_vector(0 to 4) := (Hi1, Hi1, Hi1, Hi1, Hi1);
        l0_exit_latency_diffclock: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi0);
        l0_exit_latency_sameclock: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi0);
        l0s_adj_rply_timer_dis: string  := "enable";
        l1_exit_latency_diffclock: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        l1_exit_latency_sameclock: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        l2_async_logic  : string  := "enable";
        lane_mask       : string  := "ln_mask_x4";
        lane_rate       : string  := "gen1";
        link_width      : string  := "x1";
        lmi_hold_off_cfg_timer_en: string  := "disable";
        low_priority_vc : string  := "single_vc_low_pr";
        ltr_mechanism   : string  := "false";
        ltssm_1ms_timeout: string  := "disable";
        ltssm_freqlocked_check: string  := "disable";
        malformed_tlp_truncate_en: string  := "disable";
        max_link_width  : string  := "x4_link_width";
        max_payload_size: string  := "payload_512";
        maximum_current : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        millisecond_cycle_count: vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        msi_64bit_addressing_capable: string  := "true";
        msi_masking_capable: string  := "false";
        msi_multi_message_capable: string  := "count_4";
        msi_support     : string  := "true";
        msix_pba_bir    : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        msix_pba_offset : vl_logic_vector(0 to 28) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        msix_table_bir  : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        msix_table_offset: vl_logic_vector(0 to 28) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        msix_table_size : vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        national_inst_thru_enhance: string  := "true";
        no_command_completed: string  := "true";
        no_soft_reset   : string  := "false";
        not_use_k_gbl_bits: string  := "not_used_k_gbl";
        operating_voltage: string  := "standard";
        pcie_base_spec  : string  := "pcie_2p1";
        pcie_mode       : string  := "shared_mode";
        pcie_spec_1p0_compliance: string  := "spec_1p1";
        pcie_spec_version: string  := "v2";
        pclk_out_sel    : string  := "pclk";
        pld_in_use_reg  : string  := "false";
        pm_latency_patch_dis: string  := "enable";
        pm_txdl_patch_dis: string  := "enable";
        pme_clock       : string  := "false";
        port_link_number: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        port_type       : string  := "native_ep";
        powerdown_mode  : string  := "powerup";
        prefetchable_mem_window_addr_width: string  := "prefetch_32";
        r2c_mask_easy   : string  := "false";
        r2c_mask_enable : string  := "false";
        rec_frqlk_mon_en: string  := "disable";
        register_pipe_signals: string  := "true";
        retry_buffer_last_active_address: vl_logic_vector(0 to 9) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        retry_buffer_memory_settings: vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        retry_ecc_corr_mask_dis: string  := "enable";
        revision_id     : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        role_based_error_reporting: string  := "false";
        rp_bug_fix_pri_sec_stat_reg: vl_logic_vector(0 to 6) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        rpltim_base     : vl_logic_vector(0 to 13) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rpltim_set      : string  := "false";
        rstctl_ltssm_dis: string  := "false";
        rstctrl_1ms_count_fref_clk: vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0);
        rstctrl_1us_count_fref_clk: vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        rstctrl_altpe3_crst_n_inv: string  := "false";
        rstctrl_altpe3_rst_n_inv: string  := "false";
        rstctrl_altpe3_srst_n_inv: string  := "false";
        rstctrl_chnl_cal_done_select: string  := "not_active_chnl_cal_done";
        rstctrl_debug_en: string  := "false";
        rstctrl_force_inactive_rst: string  := "false";
        rstctrl_fref_clk_select: string  := "ch0_sel";
        rstctrl_hard_block_enable: string  := "hard_rst_ctl";
        rstctrl_hip_ep  : string  := "hip_ep";
        rstctrl_mask_tx_pll_lock_select: string  := "not_active_mask_tx_pll_lock";
        rstctrl_perst_enable: string  := "level";
        rstctrl_perstn_select: string  := "perstn_pin";
        rstctrl_pld_clr : string  := "false";
        rstctrl_pll_cal_done_select: string  := "not_active_pll_cal_done";
        rstctrl_rx_pcs_rst_n_inv: string  := "false";
        rstctrl_rx_pcs_rst_n_select: string  := "not_active_rx_pcs_rst";
        rstctrl_rx_pll_freq_lock_select: string  := "not_active_rx_pll_f_lock";
        rstctrl_rx_pll_lock_select: string  := "not_active_rx_pll_lock";
        rstctrl_rx_pma_rstb_inv: string  := "false";
        rstctrl_rx_pma_rstb_select: string  := "not_active_rx_pma_rstb";
        rstctrl_timer_a : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        rstctrl_timer_a_type: string  := "a_timer_milli_secs";
        rstctrl_timer_b : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        rstctrl_timer_b_type: string  := "b_timer_milli_secs";
        rstctrl_timer_c : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        rstctrl_timer_c_type: string  := "c_timer_milli_secs";
        rstctrl_timer_d : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0);
        rstctrl_timer_d_type: string  := "d_timer_milli_secs";
        rstctrl_timer_e : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        rstctrl_timer_e_type: string  := "e_timer_milli_secs";
        rstctrl_timer_f : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        rstctrl_timer_f_type: string  := "f_timer_milli_secs";
        rstctrl_timer_g : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        rstctrl_timer_g_type: string  := "g_timer_milli_secs";
        rstctrl_timer_h : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        rstctrl_timer_h_type: string  := "h_timer_milli_secs";
        rstctrl_timer_i : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0);
        rstctrl_timer_i_type: string  := "i_timer_milli_secs";
        rstctrl_timer_j : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0);
        rstctrl_timer_j_type: string  := "j_timer_milli_secs";
        rstctrl_tx_lcff_pll_lock_select: string  := "not_active_lcff_pll_lock";
        rstctrl_tx_lcff_pll_rstb_select: string  := "not_active_lcff_pll_rstb";
        rstctrl_tx_pcs_rst_n_inv: string  := "false";
        rstctrl_tx_pcs_rst_n_select: string  := "not_active_tx_pcs_rst";
        rstctrl_tx_pma_rstb_inv: string  := "false";
        rstctrl_tx_pma_syncp_inv: string  := "false";
        rstctrl_tx_pma_syncp_select: string  := "not_active_tx_pma_syncp";
        rx_ast_parity   : string  := "disable";
        rx_buffer_credit_alloc: string  := "balance";
        rx_buffer_fc_protect: vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        rx_buffer_protect: vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        rx_cdc_almost_empty: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi1);
        rx_cdc_almost_full: vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi0, Hi0);
        rx_cred_ctl_param: string  := "disable";
        rx_ei_l0s       : string  := "disable";
        rx_l0s_count_idl: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rx_ptr0_nonposted_dpram_max: vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rx_ptr0_nonposted_dpram_min: vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rx_ptr0_posted_dpram_max: vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rx_ptr0_posted_dpram_min: vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rx_runt_patch_dis: string  := "enable";
        rx_sop_ctrl     : string  := "rx_sop_boundary_64";
        rx_trunc_patch_dis: string  := "enable";
        rx_use_prst     : string  := "false";
        rx_use_prst_ep  : string  := "true";
        rxbuf_ecc_corr_mask_dis: string  := "enable";
        rxdl_bad_sop_eop_filter_dis: string  := "rxdlbug1_enable_both";
        rxdl_bad_tlp_patch_dis: string  := "rxdlbug2_enable_both";
        rxdl_lcrc_patch_dis: string  := "rxdlbug3_enable_both";
        sameclock_nfts_count: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        sel_enable_pcs_rx_fifo_err: string  := "disable_sel";
        silicon_rev     : string  := "20nm5es";
        sim_mode        : string  := "disable";
        simple_ro_fifo_control_en: string  := "disable";
        single_rx_detect: string  := "detect_all_lanes";
        skp_os_gen3_count: vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        skp_os_schedule_count: vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        slot_number     : vl_logic_vector(0 to 12) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        slot_power_limit: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        slot_power_scale: vl_logic_vector(0 to 1) := (Hi0, Hi0);
        slotclk_cfg     : string  := "static_slotclkcfgon";
        ssid            : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ssvid           : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        subsystem_device_id: vl_logic_vector(0 to 15) := (Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        subsystem_vendor_id: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        sup_mode        : string  := "user_mode";
        surprise_down_error_support: string  := "false";
        tl_cfg_div      : string  := "cfg_clk_div_7";
        tl_tx_check_parity_msg: string  := "disable";
        tph_completer   : string  := "false";
        tx_ast_parity   : string  := "disable";
        tx_cdc_almost_empty: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi1);
        tx_cdc_almost_full: vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi0, Hi0);
        tx_sop_ctrl     : string  := "boundary_64";
        tx_swing        : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        txdl_fair_arbiter_counter: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        txdl_fair_arbiter_en: string  := "enable";
        txrate_adv      : string  := "capability";
        uc_calibration_en: string  := "uc_calibration_dis";
        use_aer         : string  := "false";
        use_crc_forwarding: string  := "false";
        user_id         : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        vc0_clk_enable  : string  := "true";
        vc0_rx_buffer_memory_settings: vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        vc0_rx_flow_ctrl_compl_data: vl_logic_vector(0 to 11) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        vc0_rx_flow_ctrl_compl_header: vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0);
        vc0_rx_flow_ctrl_nonposted_data: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        vc0_rx_flow_ctrl_nonposted_header: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi0);
        vc0_rx_flow_ctrl_posted_data: vl_logic_vector(0 to 11) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0);
        vc0_rx_flow_ctrl_posted_header: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        vc1_clk_enable  : string  := "false";
        vc_arbitration  : string  := "single_vc_arb";
        vc_enable       : string  := "single_vc";
        vendor_id       : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        vsec_cap        : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        vsec_id         : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        wrong_device_id : string  := "disable"
    );
    port(
        aer_msi_num     : in     vl_logic_vector(4 downto 0);
        app_int_err     : in     vl_logic_vector(1 downto 0);
        app_inta_sts    : in     vl_logic;
        app_msi_num     : in     vl_logic_vector(4 downto 0);
        app_msi_req     : in     vl_logic;
        app_msi_tc      : in     vl_logic_vector(2 downto 0);
        atpg_los_en_n   : in     vl_logic;
        avmm_address    : in     vl_logic_vector(9 downto 0);
        avmm_byte_en    : in     vl_logic_vector(1 downto 0);
        avmm_clk        : in     vl_logic;
        avmm_read       : in     vl_logic;
        avmm_rst_n      : in     vl_logic;
        avmm_write      : in     vl_logic;
        avmm_writedata  : in     vl_logic_vector(15 downto 0);
        bist_scanen     : in     vl_logic;
        bist_scanin     : in     vl_logic;
        bisten_rcv_n    : in     vl_logic;
        bisten_rpl_n    : in     vl_logic;
        bistmode_n      : in     vl_logic;
        cfg_link2csr_pld: in     vl_logic_vector(15 downto 0);
        cfg_prmbus_pld  : in     vl_logic_vector(7 downto 0);
        chnl_cal_done0  : in     vl_logic;
        chnl_cal_done1  : in     vl_logic;
        chnl_cal_done2  : in     vl_logic;
        chnl_cal_done3  : in     vl_logic;
        chnl_cal_done4  : in     vl_logic;
        chnl_cal_done5  : in     vl_logic;
        chnl_cal_done6  : in     vl_logic;
        chnl_cal_done7  : in     vl_logic;
        core_clk_in     : in     vl_logic;
        core_crst       : in     vl_logic;
        core_por        : in     vl_logic;
        core_rst        : in     vl_logic;
        core_srst       : in     vl_logic;
        cpl_err         : in     vl_logic_vector(6 downto 0);
        cpl_pending     : in     vl_logic;
        cseb_rddata     : in     vl_logic_vector(31 downto 0);
        cseb_rddata_parity: in     vl_logic_vector(3 downto 0);
        cseb_rdresponse : in     vl_logic_vector(4 downto 0);
        cseb_waitrequest: in     vl_logic;
        cseb_wrresp_valid: in     vl_logic;
        cseb_wrresponse : in     vl_logic_vector(4 downto 0);
        csr_cbdin       : in     vl_logic;
        csr_clk         : in     vl_logic;
        csr_din         : in     vl_logic;
        csr_en          : in     vl_logic;
        csr_enscan      : in     vl_logic;
        csr_entest      : in     vl_logic;
        csr_in          : in     vl_logic;
        csr_load_csr    : in     vl_logic;
        csr_pipe_in     : in     vl_logic;
        csr_seg         : in     vl_logic;
        csr_tcsrin      : in     vl_logic;
        csr_tverify     : in     vl_logic;
        cvp_config_done : in     vl_logic;
        cvp_config_error: in     vl_logic;
        cvp_config_ready: in     vl_logic;
        cvp_en          : in     vl_logic;
        egress_blk_err  : in     vl_logic;
        entest          : in     vl_logic;
        flr_reset       : in     vl_logic;
        force_tx_eidle  : in     vl_logic;
        fref_clk0       : in     vl_logic;
        fref_clk1       : in     vl_logic;
        fref_clk2       : in     vl_logic;
        fref_clk3       : in     vl_logic;
        fref_clk4       : in     vl_logic;
        fref_clk5       : in     vl_logic;
        fref_clk6       : in     vl_logic;
        fref_clk7       : in     vl_logic;
        frzlogic        : in     vl_logic;
        frzreg          : in     vl_logic;
        hold_ltssm_rec  : in     vl_logic;
        hpg_ctrler      : in     vl_logic_vector(4 downto 0);
        iocsrrdy_dly    : in     vl_logic;
        lmi_addr        : in     vl_logic_vector(11 downto 0);
        lmi_din         : in     vl_logic_vector(7 downto 0);
        lmi_rden        : in     vl_logic;
        lmi_wren        : in     vl_logic;
        m10k_select     : in     vl_logic_vector(2 downto 0);
        mask_tx_pll_lock0: in     vl_logic;
        mask_tx_pll_lock1: in     vl_logic;
        mask_tx_pll_lock2: in     vl_logic;
        mask_tx_pll_lock3: in     vl_logic;
        mask_tx_pll_lock4: in     vl_logic;
        mask_tx_pll_lock5: in     vl_logic;
        mask_tx_pll_lock6: in     vl_logic;
        mask_tx_pll_lock7: in     vl_logic;
        mem_hip_test_enable: in     vl_logic;
        mem_regscanen_n : in     vl_logic;
        mem_rscin_rcv_bot: in     vl_logic;
        mem_rscin_rcv_top: in     vl_logic;
        mem_rscin_rtry  : in     vl_logic;
        nfrzdrv         : in     vl_logic;
        npor            : in     vl_logic;
        pclk_central    : in     vl_logic;
        pclk_ch0        : in     vl_logic;
        pclk_ch1        : in     vl_logic;
        pex_msi_num     : in     vl_logic_vector(4 downto 0);
        phy_rst         : in     vl_logic;
        phy_srst        : in     vl_logic;
        phystatus0      : in     vl_logic;
        phystatus1      : in     vl_logic;
        phystatus2      : in     vl_logic;
        phystatus3      : in     vl_logic;
        phystatus4      : in     vl_logic;
        phystatus5      : in     vl_logic;
        phystatus6      : in     vl_logic;
        phystatus7      : in     vl_logic;
        pin_perst_n     : in     vl_logic;
        pld_clk         : in     vl_logic;
        pld_clrhip_n    : in     vl_logic;
        pld_clrpcship_n : in     vl_logic;
        pld_clrpmapcship_n: in     vl_logic;
        pld_core_ready  : in     vl_logic;
        pld_gp_status   : in     vl_logic_vector(7 downto 0);
        pld_perst_n     : in     vl_logic;
        pll_cal_done0   : in     vl_logic;
        pll_cal_done1   : in     vl_logic;
        pll_cal_done2   : in     vl_logic;
        pll_cal_done3   : in     vl_logic;
        pll_cal_done4   : in     vl_logic;
        pll_cal_done5   : in     vl_logic;
        pll_cal_done6   : in     vl_logic;
        pll_cal_done7   : in     vl_logic;
        pll_fixed_clk_central: in     vl_logic;
        pll_fixed_clk_ch0: in     vl_logic;
        pll_fixed_clk_ch1: in     vl_logic;
        plniotri        : in     vl_logic;
        pm_auxpwr       : in     vl_logic;
        pm_data         : in     vl_logic_vector(9 downto 0);
        pm_event        : in     vl_logic;
        pm_exit_d0_ack  : in     vl_logic;
        pme_to_cr       : in     vl_logic;
        reserved_clk_in : in     vl_logic;
        reserved_in     : in     vl_logic_vector(7 downto 0);
        rx_cred_ctl     : in     vl_logic_vector(15 downto 0);
        rx_pll_freq_lock0: in     vl_logic;
        rx_pll_freq_lock1: in     vl_logic;
        rx_pll_freq_lock2: in     vl_logic;
        rx_pll_freq_lock3: in     vl_logic;
        rx_pll_freq_lock4: in     vl_logic;
        rx_pll_freq_lock5: in     vl_logic;
        rx_pll_freq_lock6: in     vl_logic;
        rx_pll_freq_lock7: in     vl_logic;
        rx_pll_phase_lock0: in     vl_logic;
        rx_pll_phase_lock1: in     vl_logic;
        rx_pll_phase_lock2: in     vl_logic;
        rx_pll_phase_lock3: in     vl_logic;
        rx_pll_phase_lock4: in     vl_logic;
        rx_pll_phase_lock5: in     vl_logic;
        rx_pll_phase_lock6: in     vl_logic;
        rx_pll_phase_lock7: in     vl_logic;
        rx_st_mask      : in     vl_logic;
        rx_st_ready     : in     vl_logic;
        rxblkst0        : in     vl_logic;
        rxblkst1        : in     vl_logic;
        rxblkst2        : in     vl_logic;
        rxblkst3        : in     vl_logic;
        rxblkst4        : in     vl_logic;
        rxblkst5        : in     vl_logic;
        rxblkst6        : in     vl_logic;
        rxblkst7        : in     vl_logic;
        rxdata0         : in     vl_logic_vector(31 downto 0);
        rxdata1         : in     vl_logic_vector(31 downto 0);
        rxdata2         : in     vl_logic_vector(31 downto 0);
        rxdata3         : in     vl_logic_vector(31 downto 0);
        rxdata4         : in     vl_logic_vector(31 downto 0);
        rxdata5         : in     vl_logic_vector(31 downto 0);
        rxdata6         : in     vl_logic_vector(31 downto 0);
        rxdata7         : in     vl_logic_vector(31 downto 0);
        rxdatak0        : in     vl_logic_vector(3 downto 0);
        rxdatak1        : in     vl_logic_vector(3 downto 0);
        rxdatak2        : in     vl_logic_vector(3 downto 0);
        rxdatak3        : in     vl_logic_vector(3 downto 0);
        rxdatak4        : in     vl_logic_vector(3 downto 0);
        rxdatak5        : in     vl_logic_vector(3 downto 0);
        rxdatak6        : in     vl_logic_vector(3 downto 0);
        rxdatak7        : in     vl_logic_vector(3 downto 0);
        rxdataskip0     : in     vl_logic;
        rxdataskip1     : in     vl_logic;
        rxdataskip2     : in     vl_logic;
        rxdataskip3     : in     vl_logic;
        rxdataskip4     : in     vl_logic;
        rxdataskip5     : in     vl_logic;
        rxdataskip6     : in     vl_logic;
        rxdataskip7     : in     vl_logic;
        rxelecidle0     : in     vl_logic;
        rxelecidle1     : in     vl_logic;
        rxelecidle2     : in     vl_logic;
        rxelecidle3     : in     vl_logic;
        rxelecidle4     : in     vl_logic;
        rxelecidle5     : in     vl_logic;
        rxelecidle6     : in     vl_logic;
        rxelecidle7     : in     vl_logic;
        rxfreqlocked0   : in     vl_logic;
        rxfreqlocked1   : in     vl_logic;
        rxfreqlocked2   : in     vl_logic;
        rxfreqlocked3   : in     vl_logic;
        rxfreqlocked4   : in     vl_logic;
        rxfreqlocked5   : in     vl_logic;
        rxfreqlocked6   : in     vl_logic;
        rxfreqlocked7   : in     vl_logic;
        rxstatus0       : in     vl_logic_vector(2 downto 0);
        rxstatus1       : in     vl_logic_vector(2 downto 0);
        rxstatus2       : in     vl_logic_vector(2 downto 0);
        rxstatus3       : in     vl_logic_vector(2 downto 0);
        rxstatus4       : in     vl_logic_vector(2 downto 0);
        rxstatus5       : in     vl_logic_vector(2 downto 0);
        rxstatus6       : in     vl_logic_vector(2 downto 0);
        rxstatus7       : in     vl_logic_vector(2 downto 0);
        rxsynchd0       : in     vl_logic_vector(1 downto 0);
        rxsynchd1       : in     vl_logic_vector(1 downto 0);
        rxsynchd2       : in     vl_logic_vector(1 downto 0);
        rxsynchd3       : in     vl_logic_vector(1 downto 0);
        rxsynchd4       : in     vl_logic_vector(1 downto 0);
        rxsynchd5       : in     vl_logic_vector(1 downto 0);
        rxsynchd6       : in     vl_logic_vector(1 downto 0);
        rxsynchd7       : in     vl_logic_vector(1 downto 0);
        rxvalid0        : in     vl_logic;
        rxvalid1        : in     vl_logic;
        rxvalid2        : in     vl_logic;
        rxvalid3        : in     vl_logic;
        rxvalid4        : in     vl_logic;
        rxvalid5        : in     vl_logic;
        rxvalid6        : in     vl_logic;
        rxvalid7        : in     vl_logic;
        scan_mode_n     : in     vl_logic;
        scan_shift_n    : in     vl_logic;
        sw_ctmod        : in     vl_logic_vector(1 downto 0);
        swdn_in         : in     vl_logic_vector(2 downto 0);
        swup_in         : in     vl_logic_vector(6 downto 0);
        test_in_1_hip   : in     vl_logic_vector(31 downto 0);
        test_in_hip     : in     vl_logic_vector(31 downto 0);
        test_pl_dbg_eqin: in     vl_logic_vector(31 downto 0);
        tx_cred_cons_select: in     vl_logic;
        tx_cred_fc_sel  : in     vl_logic_vector(1 downto 0);
        tx_lcff_pll_lock0: in     vl_logic;
        tx_lcff_pll_lock1: in     vl_logic;
        tx_lcff_pll_lock2: in     vl_logic;
        tx_lcff_pll_lock3: in     vl_logic;
        tx_lcff_pll_lock4: in     vl_logic;
        tx_lcff_pll_lock5: in     vl_logic;
        tx_lcff_pll_lock6: in     vl_logic;
        tx_lcff_pll_lock7: in     vl_logic;
        tx_st_data      : in     vl_logic_vector(255 downto 0);
        tx_st_empty     : in     vl_logic_vector(1 downto 0);
        tx_st_eop       : in     vl_logic_vector(3 downto 0);
        tx_st_err       : in     vl_logic_vector(3 downto 0);
        tx_st_parity    : in     vl_logic_vector(31 downto 0);
        tx_st_sop       : in     vl_logic_vector(3 downto 0);
        tx_st_valid     : in     vl_logic;
        user_mode       : in     vl_logic;
        sta_hd_altpe3_hip_core_top_hd_altpe3_hip_core_u_clkmux_core_clk_cnt_reg_0_0_Q: out    vl_logic;
        sta_hd_altpe3_hip_core_top_hd_altpe3_hip_core_u_clkmux_core_clk_cnt_reg_1_0_Q: out    vl_logic;
        sta_hd_altpe3_hip_core_top_hd_altpe3_hip_core_u_clkmux_core_clk_cnt_reg_2_0_Q: out    vl_logic;
        app_inta_ack    : out    vl_logic;
        app_msi_ack     : out    vl_logic;
        avmm_readdata   : out    vl_logic_vector(15 downto 0);
        cfg_par_err     : out    vl_logic;
        core_clk_out    : out    vl_logic;
        cseb_addr       : out    vl_logic_vector(31 downto 0);
        cseb_addr_parity: out    vl_logic_vector(3 downto 0);
        cseb_be         : out    vl_logic_vector(3 downto 0);
        cseb_is_shadow  : out    vl_logic;
        cseb_rden       : out    vl_logic;
        cseb_wrdata     : out    vl_logic_vector(31 downto 0);
        cseb_wrdata_parity: out    vl_logic_vector(3 downto 0);
        cseb_wren       : out    vl_logic;
        cseb_wrresp_req : out    vl_logic;
        csr_dout        : out    vl_logic;
        csr_out         : out    vl_logic;
        csr_pipe_out    : out    vl_logic;
        current_coeff0  : out    vl_logic_vector(17 downto 0);
        current_coeff1  : out    vl_logic_vector(17 downto 0);
        current_coeff2  : out    vl_logic_vector(17 downto 0);
        current_coeff3  : out    vl_logic_vector(17 downto 0);
        current_coeff4  : out    vl_logic_vector(17 downto 0);
        current_coeff5  : out    vl_logic_vector(17 downto 0);
        current_coeff6  : out    vl_logic_vector(17 downto 0);
        current_coeff7  : out    vl_logic_vector(17 downto 0);
        current_rxpreset0: out    vl_logic_vector(2 downto 0);
        current_rxpreset1: out    vl_logic_vector(2 downto 0);
        current_rxpreset2: out    vl_logic_vector(2 downto 0);
        current_rxpreset3: out    vl_logic_vector(2 downto 0);
        current_rxpreset4: out    vl_logic_vector(2 downto 0);
        current_rxpreset5: out    vl_logic_vector(2 downto 0);
        current_rxpreset6: out    vl_logic_vector(2 downto 0);
        current_rxpreset7: out    vl_logic_vector(2 downto 0);
        current_speed   : out    vl_logic_vector(1 downto 0);
        cvp_clk         : out    vl_logic;
        cvp_config      : out    vl_logic;
        cvp_data        : out    vl_logic_vector(31 downto 0);
        cvp_full_config : out    vl_logic;
        cvp_start_xfer  : out    vl_logic;
        dl_up           : out    vl_logic;
        dlup_exit       : out    vl_logic;
        eidle_infer_sel0: out    vl_logic_vector(2 downto 0);
        eidle_infer_sel1: out    vl_logic_vector(2 downto 0);
        eidle_infer_sel2: out    vl_logic_vector(2 downto 0);
        eidle_infer_sel3: out    vl_logic_vector(2 downto 0);
        eidle_infer_sel4: out    vl_logic_vector(2 downto 0);
        eidle_infer_sel5: out    vl_logic_vector(2 downto 0);
        eidle_infer_sel6: out    vl_logic_vector(2 downto 0);
        eidle_infer_sel7: out    vl_logic_vector(2 downto 0);
        ev_128ns        : out    vl_logic;
        ev_1us          : out    vl_logic;
        flr_sts         : out    vl_logic;
        g3_rx_pcs_rst_n0: out    vl_logic;
        g3_rx_pcs_rst_n1: out    vl_logic;
        g3_rx_pcs_rst_n2: out    vl_logic;
        g3_rx_pcs_rst_n3: out    vl_logic;
        g3_rx_pcs_rst_n4: out    vl_logic;
        g3_rx_pcs_rst_n5: out    vl_logic;
        g3_rx_pcs_rst_n6: out    vl_logic;
        g3_rx_pcs_rst_n7: out    vl_logic;
        g3_tx_pcs_rst_n0: out    vl_logic;
        g3_tx_pcs_rst_n1: out    vl_logic;
        g3_tx_pcs_rst_n2: out    vl_logic;
        g3_tx_pcs_rst_n3: out    vl_logic;
        g3_tx_pcs_rst_n4: out    vl_logic;
        g3_tx_pcs_rst_n5: out    vl_logic;
        g3_tx_pcs_rst_n6: out    vl_logic;
        g3_tx_pcs_rst_n7: out    vl_logic;
        hotrst_exit     : out    vl_logic;
        int_status      : out    vl_logic_vector(3 downto 0);
        k_hip_pcs_chnl_en: out    vl_logic_vector(7 downto 0);
        k_hrc_chnl_en   : out    vl_logic_vector(7 downto 0);
        k_hrc_chnl_txpll_master_cgb_rst_en: out    vl_logic_vector(7 downto 0);
        k_hrc_chnl_txpll_rst_en: out    vl_logic_vector(7 downto 0);
        l2_exit         : out    vl_logic;
        lane_act        : out    vl_logic_vector(3 downto 0);
        lmi_ack         : out    vl_logic;
        lmi_dout        : out    vl_logic_vector(7 downto 0);
        ltssm_state     : out    vl_logic_vector(4 downto 0);
        mem_rscout_rcv_bot: out    vl_logic;
        mem_rscout_rcv_top: out    vl_logic;
        mem_rscout_rtry : out    vl_logic;
        pld_clk_in_use  : out    vl_logic;
        pld_gp_ctrl     : out    vl_logic_vector(7 downto 0);
        pm_exit_d0_req  : out    vl_logic;
        pme_to_sr       : out    vl_logic;
        powerdown0      : out    vl_logic_vector(1 downto 0);
        powerdown1      : out    vl_logic_vector(1 downto 0);
        powerdown2      : out    vl_logic_vector(1 downto 0);
        powerdown3      : out    vl_logic_vector(1 downto 0);
        powerdown4      : out    vl_logic_vector(1 downto 0);
        powerdown5      : out    vl_logic_vector(1 downto 0);
        powerdown6      : out    vl_logic_vector(1 downto 0);
        powerdown7      : out    vl_logic_vector(1 downto 0);
        r2c_unc_ecc     : out    vl_logic;
        rate0           : out    vl_logic_vector(1 downto 0);
        rate1           : out    vl_logic_vector(1 downto 0);
        rate2           : out    vl_logic_vector(1 downto 0);
        rate3           : out    vl_logic_vector(1 downto 0);
        rate4           : out    vl_logic_vector(1 downto 0);
        rate5           : out    vl_logic_vector(1 downto 0);
        rate6           : out    vl_logic_vector(1 downto 0);
        rate7           : out    vl_logic_vector(1 downto 0);
        rate_ctrl       : out    vl_logic_vector(1 downto 0);
        reserved_clk_out: out    vl_logic;
        reserved_out    : out    vl_logic_vector(7 downto 0);
        reset_status    : out    vl_logic;
        retry_corr_ecc  : out    vl_logic;
        retry_unc_ecc   : out    vl_logic;
        rx_corr_ecc     : out    vl_logic;
        rx_cred_status  : out    vl_logic_vector(19 downto 0);
        rx_par_err      : out    vl_logic;
        rx_pcs_rst_n0   : out    vl_logic;
        rx_pcs_rst_n1   : out    vl_logic;
        rx_pcs_rst_n2   : out    vl_logic;
        rx_pcs_rst_n3   : out    vl_logic;
        rx_pcs_rst_n4   : out    vl_logic;
        rx_pcs_rst_n5   : out    vl_logic;
        rx_pcs_rst_n6   : out    vl_logic;
        rx_pcs_rst_n7   : out    vl_logic;
        rx_pma_rstb0    : out    vl_logic;
        rx_pma_rstb1    : out    vl_logic;
        rx_pma_rstb2    : out    vl_logic;
        rx_pma_rstb3    : out    vl_logic;
        rx_pma_rstb4    : out    vl_logic;
        rx_pma_rstb5    : out    vl_logic;
        rx_pma_rstb6    : out    vl_logic;
        rx_pma_rstb7    : out    vl_logic;
        rx_st_bardec1   : out    vl_logic_vector(7 downto 0);
        rx_st_bardec2   : out    vl_logic_vector(7 downto 0);
        rx_st_be        : out    vl_logic_vector(31 downto 0);
        rx_st_data      : out    vl_logic_vector(255 downto 0);
        rx_st_empty     : out    vl_logic_vector(1 downto 0);
        rx_st_eop       : out    vl_logic_vector(3 downto 0);
        rx_st_err       : out    vl_logic_vector(3 downto 0);
        rx_st_parity    : out    vl_logic_vector(31 downto 0);
        rx_st_sop       : out    vl_logic_vector(3 downto 0);
        rx_st_valid     : out    vl_logic_vector(3 downto 0);
        rxfc_cplbuf_ovf : out    vl_logic;
        rxfc_cplovf_tag : out    vl_logic_vector(7 downto 0);
        rxpolarity0     : out    vl_logic;
        rxpolarity1     : out    vl_logic;
        rxpolarity2     : out    vl_logic;
        rxpolarity3     : out    vl_logic;
        rxpolarity4     : out    vl_logic;
        rxpolarity5     : out    vl_logic;
        rxpolarity6     : out    vl_logic;
        rxpolarity7     : out    vl_logic;
        serr_out        : out    vl_logic;
        swdn_out        : out    vl_logic_vector(6 downto 0);
        swup_out        : out    vl_logic_vector(2 downto 0);
        test_fref_clk   : out    vl_logic;
        test_out_1_hip  : out    vl_logic_vector(63 downto 0);
        test_out_hip    : out    vl_logic_vector(255 downto 0);
        tl_cfg_add      : out    vl_logic_vector(3 downto 0);
        tl_cfg_ctl      : out    vl_logic_vector(31 downto 0);
        tl_cfg_sts      : out    vl_logic_vector(52 downto 0);
        tl_cfg_sts_wr   : out    vl_logic;
        tx_cred_data_fc : out    vl_logic_vector(11 downto 0);
        tx_cred_fc_hip_cons: out    vl_logic_vector(5 downto 0);
        tx_cred_fc_infinite: out    vl_logic_vector(5 downto 0);
        tx_cred_hdr_fc  : out    vl_logic_vector(7 downto 0);
        tx_deemph0      : out    vl_logic;
        tx_deemph1      : out    vl_logic;
        tx_deemph2      : out    vl_logic;
        tx_deemph3      : out    vl_logic;
        tx_deemph4      : out    vl_logic;
        tx_deemph5      : out    vl_logic;
        tx_deemph6      : out    vl_logic;
        tx_deemph7      : out    vl_logic;
        tx_lcff_pll_rstb0: out    vl_logic;
        tx_lcff_pll_rstb1: out    vl_logic;
        tx_lcff_pll_rstb2: out    vl_logic;
        tx_lcff_pll_rstb3: out    vl_logic;
        tx_lcff_pll_rstb4: out    vl_logic;
        tx_lcff_pll_rstb5: out    vl_logic;
        tx_lcff_pll_rstb6: out    vl_logic;
        tx_lcff_pll_rstb7: out    vl_logic;
        tx_margin0      : out    vl_logic_vector(2 downto 0);
        tx_margin1      : out    vl_logic_vector(2 downto 0);
        tx_margin2      : out    vl_logic_vector(2 downto 0);
        tx_margin3      : out    vl_logic_vector(2 downto 0);
        tx_margin4      : out    vl_logic_vector(2 downto 0);
        tx_margin5      : out    vl_logic_vector(2 downto 0);
        tx_margin6      : out    vl_logic_vector(2 downto 0);
        tx_margin7      : out    vl_logic_vector(2 downto 0);
        tx_par_err      : out    vl_logic_vector(1 downto 0);
        tx_pcs_rst_n0   : out    vl_logic;
        tx_pcs_rst_n1   : out    vl_logic;
        tx_pcs_rst_n2   : out    vl_logic;
        tx_pcs_rst_n3   : out    vl_logic;
        tx_pcs_rst_n4   : out    vl_logic;
        tx_pcs_rst_n5   : out    vl_logic;
        tx_pcs_rst_n6   : out    vl_logic;
        tx_pcs_rst_n7   : out    vl_logic;
        tx_pma_syncp0   : out    vl_logic;
        tx_pma_syncp1   : out    vl_logic;
        tx_pma_syncp2   : out    vl_logic;
        tx_pma_syncp3   : out    vl_logic;
        tx_pma_syncp4   : out    vl_logic;
        tx_pma_syncp5   : out    vl_logic;
        tx_pma_syncp6   : out    vl_logic;
        tx_pma_syncp7   : out    vl_logic;
        tx_st_ready     : out    vl_logic;
        txblkst0        : out    vl_logic;
        txblkst1        : out    vl_logic;
        txblkst2        : out    vl_logic;
        txblkst3        : out    vl_logic;
        txblkst4        : out    vl_logic;
        txblkst5        : out    vl_logic;
        txblkst6        : out    vl_logic;
        txblkst7        : out    vl_logic;
        txcompl0        : out    vl_logic;
        txcompl1        : out    vl_logic;
        txcompl2        : out    vl_logic;
        txcompl3        : out    vl_logic;
        txcompl4        : out    vl_logic;
        txcompl5        : out    vl_logic;
        txcompl6        : out    vl_logic;
        txcompl7        : out    vl_logic;
        txdata0         : out    vl_logic_vector(31 downto 0);
        txdata1         : out    vl_logic_vector(31 downto 0);
        txdata2         : out    vl_logic_vector(31 downto 0);
        txdata3         : out    vl_logic_vector(31 downto 0);
        txdata4         : out    vl_logic_vector(31 downto 0);
        txdata5         : out    vl_logic_vector(31 downto 0);
        txdata6         : out    vl_logic_vector(31 downto 0);
        txdata7         : out    vl_logic_vector(31 downto 0);
        txdatak0        : out    vl_logic_vector(3 downto 0);
        txdatak1        : out    vl_logic_vector(3 downto 0);
        txdatak2        : out    vl_logic_vector(3 downto 0);
        txdatak3        : out    vl_logic_vector(3 downto 0);
        txdatak4        : out    vl_logic_vector(3 downto 0);
        txdatak5        : out    vl_logic_vector(3 downto 0);
        txdatak6        : out    vl_logic_vector(3 downto 0);
        txdatak7        : out    vl_logic_vector(3 downto 0);
        txdataskip0     : out    vl_logic;
        txdataskip1     : out    vl_logic;
        txdataskip2     : out    vl_logic;
        txdataskip3     : out    vl_logic;
        txdataskip4     : out    vl_logic;
        txdataskip5     : out    vl_logic;
        txdataskip6     : out    vl_logic;
        txdataskip7     : out    vl_logic;
        txdetectrx0     : out    vl_logic;
        txdetectrx1     : out    vl_logic;
        txdetectrx2     : out    vl_logic;
        txdetectrx3     : out    vl_logic;
        txdetectrx4     : out    vl_logic;
        txdetectrx5     : out    vl_logic;
        txdetectrx6     : out    vl_logic;
        txdetectrx7     : out    vl_logic;
        txelecidle0     : out    vl_logic;
        txelecidle1     : out    vl_logic;
        txelecidle2     : out    vl_logic;
        txelecidle3     : out    vl_logic;
        txelecidle4     : out    vl_logic;
        txelecidle5     : out    vl_logic;
        txelecidle6     : out    vl_logic;
        txelecidle7     : out    vl_logic;
        txst_prot_err   : out    vl_logic;
        txswing0        : out    vl_logic;
        txswing1        : out    vl_logic;
        txswing2        : out    vl_logic;
        txswing3        : out    vl_logic;
        txswing4        : out    vl_logic;
        txswing5        : out    vl_logic;
        txswing6        : out    vl_logic;
        txswing7        : out    vl_logic;
        txsynchd0       : out    vl_logic_vector(1 downto 0);
        txsynchd1       : out    vl_logic_vector(1 downto 0);
        txsynchd2       : out    vl_logic_vector(1 downto 0);
        txsynchd3       : out    vl_logic_vector(1 downto 0);
        txsynchd4       : out    vl_logic_vector(1 downto 0);
        txsynchd5       : out    vl_logic_vector(1 downto 0);
        txsynchd6       : out    vl_logic_vector(1 downto 0);
        txsynchd7       : out    vl_logic_vector(1 downto 0);
        wake_oen        : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of enable_debug_info : constant is 1;
    attribute mti_svvh_generic_type of acknack_base : constant is 1;
    attribute mti_svvh_generic_type of acknack_set : constant is 1;
    attribute mti_svvh_generic_type of advance_error_reporting : constant is 1;
    attribute mti_svvh_generic_type of app_interface_width : constant is 1;
    attribute mti_svvh_generic_type of arb_upfc_30us_counter : constant is 1;
    attribute mti_svvh_generic_type of arb_upfc_30us_en : constant is 1;
    attribute mti_svvh_generic_type of aspm_config_management : constant is 1;
    attribute mti_svvh_generic_type of aspm_patch_disable : constant is 1;
    attribute mti_svvh_generic_type of ast_width_rx : constant is 1;
    attribute mti_svvh_generic_type of ast_width_tx : constant is 1;
    attribute mti_svvh_generic_type of atomic_malformed : constant is 1;
    attribute mti_svvh_generic_type of atomic_op_completer_32bit : constant is 1;
    attribute mti_svvh_generic_type of atomic_op_completer_64bit : constant is 1;
    attribute mti_svvh_generic_type of atomic_op_routing : constant is 1;
    attribute mti_svvh_generic_type of auto_msg_drop_enable : constant is 1;
    attribute mti_svvh_generic_type of avmm_cvp_inter_sel_csr_ctrl : constant is 1;
    attribute mti_svvh_generic_type of avmm_dprio_broadcast_en_csr_ctrl : constant is 1;
    attribute mti_svvh_generic_type of avmm_force_inter_sel_csr_ctrl : constant is 1;
    attribute mti_svvh_generic_type of avmm_power_iso_en_csr_ctrl : constant is 1;
    attribute mti_svvh_generic_type of bar0_size_mask : constant is 1;
    attribute mti_svvh_generic_type of bar0_type : constant is 1;
    attribute mti_svvh_generic_type of bar1_size_mask : constant is 1;
    attribute mti_svvh_generic_type of bar1_type : constant is 1;
    attribute mti_svvh_generic_type of bar2_size_mask : constant is 1;
    attribute mti_svvh_generic_type of bar2_type : constant is 1;
    attribute mti_svvh_generic_type of bar3_size_mask : constant is 1;
    attribute mti_svvh_generic_type of bar3_type : constant is 1;
    attribute mti_svvh_generic_type of bar4_size_mask : constant is 1;
    attribute mti_svvh_generic_type of bar4_type : constant is 1;
    attribute mti_svvh_generic_type of bar5_size_mask : constant is 1;
    attribute mti_svvh_generic_type of bar5_type : constant is 1;
    attribute mti_svvh_generic_type of base_counter_sel : constant is 1;
    attribute mti_svvh_generic_type of bist_memory_settings : constant is 1;
    attribute mti_svvh_generic_type of bridge_port_ssid_support : constant is 1;
    attribute mti_svvh_generic_type of bridge_port_vga_enable : constant is 1;
    attribute mti_svvh_generic_type of bypass_cdc : constant is 1;
    attribute mti_svvh_generic_type of bypass_clk_switch : constant is 1;
    attribute mti_svvh_generic_type of bypass_tl : constant is 1;
    attribute mti_svvh_generic_type of capab_rate_rxcfg_en : constant is 1;
    attribute mti_svvh_generic_type of cas_completer_128bit : constant is 1;
    attribute mti_svvh_generic_type of cdc_clk_relation : constant is 1;
    attribute mti_svvh_generic_type of cdc_dummy_insert_limit : constant is 1;
    attribute mti_svvh_generic_type of cfg_parchk_ena : constant is 1;
    attribute mti_svvh_generic_type of cfgbp_req_recov_disable : constant is 1;
    attribute mti_svvh_generic_type of class_code : constant is 1;
    attribute mti_svvh_generic_type of clock_pwr_management : constant is 1;
    attribute mti_svvh_generic_type of completion_timeout : constant is 1;
    attribute mti_svvh_generic_type of core_clk_divider : constant is 1;
    attribute mti_svvh_generic_type of core_clk_freq_mhz : constant is 1;
    attribute mti_svvh_generic_type of core_clk_out_sel : constant is 1;
    attribute mti_svvh_generic_type of core_clk_sel : constant is 1;
    attribute mti_svvh_generic_type of core_clk_source : constant is 1;
    attribute mti_svvh_generic_type of cseb_bar_match_checking : constant is 1;
    attribute mti_svvh_generic_type of cseb_config_bypass : constant is 1;
    attribute mti_svvh_generic_type of cseb_cpl_status_during_cvp : constant is 1;
    attribute mti_svvh_generic_type of cseb_cpl_tag_checking : constant is 1;
    attribute mti_svvh_generic_type of cseb_disable_auto_crs : constant is 1;
    attribute mti_svvh_generic_type of cseb_extend_pci : constant is 1;
    attribute mti_svvh_generic_type of cseb_extend_pcie : constant is 1;
    attribute mti_svvh_generic_type of cseb_min_error_checking : constant is 1;
    attribute mti_svvh_generic_type of cseb_route_to_avl_rx_st : constant is 1;
    attribute mti_svvh_generic_type of cseb_temp_busy_crs : constant is 1;
    attribute mti_svvh_generic_type of cvp_clk_reset : constant is 1;
    attribute mti_svvh_generic_type of cvp_data_compressed : constant is 1;
    attribute mti_svvh_generic_type of cvp_data_encrypted : constant is 1;
    attribute mti_svvh_generic_type of cvp_enable : constant is 1;
    attribute mti_svvh_generic_type of cvp_mode_reset : constant is 1;
    attribute mti_svvh_generic_type of cvp_rate_sel : constant is 1;
    attribute mti_svvh_generic_type of d0_pme : constant is 1;
    attribute mti_svvh_generic_type of d1_pme : constant is 1;
    attribute mti_svvh_generic_type of d1_support : constant is 1;
    attribute mti_svvh_generic_type of d2_pme : constant is 1;
    attribute mti_svvh_generic_type of d2_support : constant is 1;
    attribute mti_svvh_generic_type of d3_cold_pme : constant is 1;
    attribute mti_svvh_generic_type of d3_hot_pme : constant is 1;
    attribute mti_svvh_generic_type of data_pack_rx : constant is 1;
    attribute mti_svvh_generic_type of deemphasis_enable : constant is 1;
    attribute mti_svvh_generic_type of deskew_comma : constant is 1;
    attribute mti_svvh_generic_type of device_id : constant is 1;
    attribute mti_svvh_generic_type of device_number : constant is 1;
    attribute mti_svvh_generic_type of device_specific_init : constant is 1;
    attribute mti_svvh_generic_type of dft_clock_obsrv_en : constant is 1;
    attribute mti_svvh_generic_type of dft_clock_obsrv_sel : constant is 1;
    attribute mti_svvh_generic_type of diffclock_nfts_count : constant is 1;
    attribute mti_svvh_generic_type of dis_cplovf : constant is 1;
    attribute mti_svvh_generic_type of dis_paritychk : constant is 1;
    attribute mti_svvh_generic_type of disable_link_x2_support : constant is 1;
    attribute mti_svvh_generic_type of disable_snoop_packet : constant is 1;
    attribute mti_svvh_generic_type of dl_tx_check_parity_edb : constant is 1;
    attribute mti_svvh_generic_type of dll_active_report_support : constant is 1;
    attribute mti_svvh_generic_type of early_dl_up : constant is 1;
    attribute mti_svvh_generic_type of ecrc_check_capable : constant is 1;
    attribute mti_svvh_generic_type of ecrc_gen_capable : constant is 1;
    attribute mti_svvh_generic_type of egress_block_err_report_ena : constant is 1;
    attribute mti_svvh_generic_type of ei_delay_powerdown_count : constant is 1;
    attribute mti_svvh_generic_type of eie_before_nfts_count : constant is 1;
    attribute mti_svvh_generic_type of electromech_interlock : constant is 1;
    attribute mti_svvh_generic_type of en_ieiupdatefc : constant is 1;
    attribute mti_svvh_generic_type of en_lane_errchk : constant is 1;
    attribute mti_svvh_generic_type of en_phystatus_dly : constant is 1;
    attribute mti_svvh_generic_type of ena_ido_cpl : constant is 1;
    attribute mti_svvh_generic_type of ena_ido_req : constant is 1;
    attribute mti_svvh_generic_type of enable_adapter_half_rate_mode : constant is 1;
    attribute mti_svvh_generic_type of enable_ch01_pclk_out : constant is 1;
    attribute mti_svvh_generic_type of enable_ch0_pclk_out : constant is 1;
    attribute mti_svvh_generic_type of enable_completion_timeout_disable : constant is 1;
    attribute mti_svvh_generic_type of enable_directed_spd_chng : constant is 1;
    attribute mti_svvh_generic_type of enable_function_msix_support : constant is 1;
    attribute mti_svvh_generic_type of enable_l0s_aspm : constant is 1;
    attribute mti_svvh_generic_type of enable_l1_aspm : constant is 1;
    attribute mti_svvh_generic_type of enable_rx_buffer_checking : constant is 1;
    attribute mti_svvh_generic_type of enable_rx_reordering : constant is 1;
    attribute mti_svvh_generic_type of enable_slot_register : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l0_latency : constant is 1;
    attribute mti_svvh_generic_type of endpoint_l1_latency : constant is 1;
    attribute mti_svvh_generic_type of eql_rq_int_en_number : constant is 1;
    attribute mti_svvh_generic_type of errmgt_fcpe_patch_dis : constant is 1;
    attribute mti_svvh_generic_type of errmgt_fep_patch_dis : constant is 1;
    attribute mti_svvh_generic_type of expansion_base_address_register : constant is 1;
    attribute mti_svvh_generic_type of extend_tag_field : constant is 1;
    attribute mti_svvh_generic_type of extended_format_field : constant is 1;
    attribute mti_svvh_generic_type of extended_tag_reset : constant is 1;
    attribute mti_svvh_generic_type of fc_init_timer : constant is 1;
    attribute mti_svvh_generic_type of flow_control_timeout_count : constant is 1;
    attribute mti_svvh_generic_type of flow_control_update_count : constant is 1;
    attribute mti_svvh_generic_type of flr_capability : constant is 1;
    attribute mti_svvh_generic_type of force_dis_to_det : constant is 1;
    attribute mti_svvh_generic_type of force_gen1_dis : constant is 1;
    attribute mti_svvh_generic_type of force_tx_coeff_preset_lpbk : constant is 1;
    attribute mti_svvh_generic_type of frame_err_patch_dis : constant is 1;
    attribute mti_svvh_generic_type of func_mode : constant is 1;
    attribute mti_svvh_generic_type of g3_bypass_equlz : constant is 1;
    attribute mti_svvh_generic_type of g3_coeff_done_tmout : constant is 1;
    attribute mti_svvh_generic_type of g3_deskew_char : constant is 1;
    attribute mti_svvh_generic_type of g3_dis_be_frm_err : constant is 1;
    attribute mti_svvh_generic_type of g3_dn_rx_hint_eqlz_0 : constant is 1;
    attribute mti_svvh_generic_type of g3_dn_rx_hint_eqlz_1 : constant is 1;
    attribute mti_svvh_generic_type of g3_dn_rx_hint_eqlz_2 : constant is 1;
    attribute mti_svvh_generic_type of g3_dn_rx_hint_eqlz_3 : constant is 1;
    attribute mti_svvh_generic_type of g3_dn_rx_hint_eqlz_4 : constant is 1;
    attribute mti_svvh_generic_type of g3_dn_rx_hint_eqlz_5 : constant is 1;
    attribute mti_svvh_generic_type of g3_dn_rx_hint_eqlz_6 : constant is 1;
    attribute mti_svvh_generic_type of g3_dn_rx_hint_eqlz_7 : constant is 1;
    attribute mti_svvh_generic_type of g3_dn_tx_preset_eqlz_0 : constant is 1;
    attribute mti_svvh_generic_type of g3_dn_tx_preset_eqlz_1 : constant is 1;
    attribute mti_svvh_generic_type of g3_dn_tx_preset_eqlz_2 : constant is 1;
    attribute mti_svvh_generic_type of g3_dn_tx_preset_eqlz_3 : constant is 1;
    attribute mti_svvh_generic_type of g3_dn_tx_preset_eqlz_4 : constant is 1;
    attribute mti_svvh_generic_type of g3_dn_tx_preset_eqlz_5 : constant is 1;
    attribute mti_svvh_generic_type of g3_dn_tx_preset_eqlz_6 : constant is 1;
    attribute mti_svvh_generic_type of g3_dn_tx_preset_eqlz_7 : constant is 1;
    attribute mti_svvh_generic_type of g3_force_ber_max : constant is 1;
    attribute mti_svvh_generic_type of g3_force_ber_min : constant is 1;
    attribute mti_svvh_generic_type of g3_lnk_trn_rx_ts : constant is 1;
    attribute mti_svvh_generic_type of g3_ltssm_eq_dbg : constant is 1;
    attribute mti_svvh_generic_type of g3_ltssm_rec_dbg : constant is 1;
    attribute mti_svvh_generic_type of g3_pause_ltssm_rec_en : constant is 1;
    attribute mti_svvh_generic_type of g3_quiesce_guarant : constant is 1;
    attribute mti_svvh_generic_type of g3_redo_equlz_dis : constant is 1;
    attribute mti_svvh_generic_type of g3_redo_equlz_en : constant is 1;
    attribute mti_svvh_generic_type of g3_up_rx_hint_eqlz_0 : constant is 1;
    attribute mti_svvh_generic_type of g3_up_rx_hint_eqlz_1 : constant is 1;
    attribute mti_svvh_generic_type of g3_up_rx_hint_eqlz_2 : constant is 1;
    attribute mti_svvh_generic_type of g3_up_rx_hint_eqlz_3 : constant is 1;
    attribute mti_svvh_generic_type of g3_up_rx_hint_eqlz_4 : constant is 1;
    attribute mti_svvh_generic_type of g3_up_rx_hint_eqlz_5 : constant is 1;
    attribute mti_svvh_generic_type of g3_up_rx_hint_eqlz_6 : constant is 1;
    attribute mti_svvh_generic_type of g3_up_rx_hint_eqlz_7 : constant is 1;
    attribute mti_svvh_generic_type of g3_up_tx_preset_eqlz_0 : constant is 1;
    attribute mti_svvh_generic_type of g3_up_tx_preset_eqlz_1 : constant is 1;
    attribute mti_svvh_generic_type of g3_up_tx_preset_eqlz_2 : constant is 1;
    attribute mti_svvh_generic_type of g3_up_tx_preset_eqlz_3 : constant is 1;
    attribute mti_svvh_generic_type of g3_up_tx_preset_eqlz_4 : constant is 1;
    attribute mti_svvh_generic_type of g3_up_tx_preset_eqlz_5 : constant is 1;
    attribute mti_svvh_generic_type of g3_up_tx_preset_eqlz_6 : constant is 1;
    attribute mti_svvh_generic_type of g3_up_tx_preset_eqlz_7 : constant is 1;
    attribute mti_svvh_generic_type of gen123_lane_rate_mode : constant is 1;
    attribute mti_svvh_generic_type of gen2_diffclock_nfts_count : constant is 1;
    attribute mti_svvh_generic_type of gen2_pma_pll_usage : constant is 1;
    attribute mti_svvh_generic_type of gen2_sameclock_nfts_count : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_1 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_10 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_10_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_10_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_10_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_10_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_10_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_10_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_11 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_11_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_11_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_11_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_11_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_11_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_11_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_12 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_12_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_12_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_12_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_12_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_12_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_12_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_13 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_13_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_13_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_13_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_13_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_13_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_13_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_14 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_14_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_14_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_14_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_14_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_14_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_14_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_15 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_15_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_15_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_15_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_15_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_15_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_15_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_16 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_16_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_16_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_16_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_16_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_16_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_16_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_17 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_17_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_17_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_17_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_17_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_17_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_17_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_18 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_18_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_18_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_18_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_18_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_18_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_18_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_19 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_19_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_19_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_19_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_19_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_19_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_19_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_1_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_1_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_1_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_1_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_1_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_1_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_2 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_20 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_20_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_20_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_20_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_20_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_20_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_20_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_21 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_21_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_21_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_21_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_21_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_21_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_21_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_22 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_22_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_22_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_22_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_22_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_22_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_22_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_23 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_23_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_23_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_23_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_23_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_23_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_23_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_24 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_24_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_24_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_24_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_24_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_24_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_24_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_2_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_2_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_2_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_2_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_2_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_2_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_3 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_3_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_3_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_3_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_3_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_3_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_3_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_4 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_4_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_4_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_4_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_4_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_4_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_4_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_5 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_5_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_5_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_5_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_5_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_5_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_5_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_6 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_6_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_6_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_6_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_6_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_6_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_6_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_7 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_7_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_7_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_7_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_7_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_7_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_7_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_8 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_8_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_8_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_8_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_8_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_8_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_8_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_9 : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_9_ber_meas : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_9_nxtber_less : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_9_nxtber_more : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_9_preset_hint : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_9_reqber : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_9_sel : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_delay_count : constant is 1;
    attribute mti_svvh_generic_type of gen3_coeff_errchk : constant is 1;
    attribute mti_svvh_generic_type of gen3_dcbal_en : constant is 1;
    attribute mti_svvh_generic_type of gen3_diffclock_nfts_count : constant is 1;
    attribute mti_svvh_generic_type of gen3_force_local_coeff : constant is 1;
    attribute mti_svvh_generic_type of gen3_full_swing : constant is 1;
    attribute mti_svvh_generic_type of gen3_half_swing : constant is 1;
    attribute mti_svvh_generic_type of gen3_low_freq : constant is 1;
    attribute mti_svvh_generic_type of gen3_paritychk : constant is 1;
    attribute mti_svvh_generic_type of gen3_pl_framing_err_dis : constant is 1;
    attribute mti_svvh_generic_type of gen3_preset_coeff_1 : constant is 1;
    attribute mti_svvh_generic_type of gen3_preset_coeff_10 : constant is 1;
    attribute mti_svvh_generic_type of gen3_preset_coeff_11 : constant is 1;
    attribute mti_svvh_generic_type of gen3_preset_coeff_2 : constant is 1;
    attribute mti_svvh_generic_type of gen3_preset_coeff_3 : constant is 1;
    attribute mti_svvh_generic_type of gen3_preset_coeff_4 : constant is 1;
    attribute mti_svvh_generic_type of gen3_preset_coeff_5 : constant is 1;
    attribute mti_svvh_generic_type of gen3_preset_coeff_6 : constant is 1;
    attribute mti_svvh_generic_type of gen3_preset_coeff_7 : constant is 1;
    attribute mti_svvh_generic_type of gen3_preset_coeff_8 : constant is 1;
    attribute mti_svvh_generic_type of gen3_preset_coeff_9 : constant is 1;
    attribute mti_svvh_generic_type of gen3_reset_eieos_cnt_bit : constant is 1;
    attribute mti_svvh_generic_type of gen3_rxfreqlock_counter : constant is 1;
    attribute mti_svvh_generic_type of gen3_sameclock_nfts_count : constant is 1;
    attribute mti_svvh_generic_type of gen3_scrdscr_bypass : constant is 1;
    attribute mti_svvh_generic_type of gen3_skip_ph2_ph3 : constant is 1;
    attribute mti_svvh_generic_type of hard_reset_bypass : constant is 1;
    attribute mti_svvh_generic_type of hard_rst_sig_chnl_en : constant is 1;
    attribute mti_svvh_generic_type of hard_rst_tx_pll_rst_chnl_en : constant is 1;
    attribute mti_svvh_generic_type of hip_ac_pwr_clk_freq_in_hz : constant is 1;
    attribute mti_svvh_generic_type of hip_ac_pwr_uw_per_mhz : constant is 1;
    attribute mti_svvh_generic_type of hip_base_address : constant is 1;
    attribute mti_svvh_generic_type of hip_clock_dis : constant is 1;
    attribute mti_svvh_generic_type of hip_hard_reset : constant is 1;
    attribute mti_svvh_generic_type of hip_pcs_sig_chnl_en : constant is 1;
    attribute mti_svvh_generic_type of hot_plug_support : constant is 1;
    attribute mti_svvh_generic_type of hrc_chnl_txpll_master_cgb_rst_select : constant is 1;
    attribute mti_svvh_generic_type of hrdrstctrl_en : constant is 1;
    attribute mti_svvh_generic_type of iei_enable_settings : constant is 1;
    attribute mti_svvh_generic_type of indicator : constant is 1;
    attribute mti_svvh_generic_type of intel_id_access : constant is 1;
    attribute mti_svvh_generic_type of interrupt_pin : constant is 1;
    attribute mti_svvh_generic_type of io_window_addr_width : constant is 1;
    attribute mti_svvh_generic_type of jtag_id : constant is 1;
    attribute mti_svvh_generic_type of ko_compl_data : constant is 1;
    attribute mti_svvh_generic_type of ko_compl_header : constant is 1;
    attribute mti_svvh_generic_type of l01_entry_latency : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_diffclock : constant is 1;
    attribute mti_svvh_generic_type of l0_exit_latency_sameclock : constant is 1;
    attribute mti_svvh_generic_type of l0s_adj_rply_timer_dis : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_diffclock : constant is 1;
    attribute mti_svvh_generic_type of l1_exit_latency_sameclock : constant is 1;
    attribute mti_svvh_generic_type of l2_async_logic : constant is 1;
    attribute mti_svvh_generic_type of lane_mask : constant is 1;
    attribute mti_svvh_generic_type of lane_rate : constant is 1;
    attribute mti_svvh_generic_type of link_width : constant is 1;
    attribute mti_svvh_generic_type of lmi_hold_off_cfg_timer_en : constant is 1;
    attribute mti_svvh_generic_type of low_priority_vc : constant is 1;
    attribute mti_svvh_generic_type of ltr_mechanism : constant is 1;
    attribute mti_svvh_generic_type of ltssm_1ms_timeout : constant is 1;
    attribute mti_svvh_generic_type of ltssm_freqlocked_check : constant is 1;
    attribute mti_svvh_generic_type of malformed_tlp_truncate_en : constant is 1;
    attribute mti_svvh_generic_type of max_link_width : constant is 1;
    attribute mti_svvh_generic_type of max_payload_size : constant is 1;
    attribute mti_svvh_generic_type of maximum_current : constant is 1;
    attribute mti_svvh_generic_type of millisecond_cycle_count : constant is 1;
    attribute mti_svvh_generic_type of msi_64bit_addressing_capable : constant is 1;
    attribute mti_svvh_generic_type of msi_masking_capable : constant is 1;
    attribute mti_svvh_generic_type of msi_multi_message_capable : constant is 1;
    attribute mti_svvh_generic_type of msi_support : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_bir : constant is 1;
    attribute mti_svvh_generic_type of msix_pba_offset : constant is 1;
    attribute mti_svvh_generic_type of msix_table_bir : constant is 1;
    attribute mti_svvh_generic_type of msix_table_offset : constant is 1;
    attribute mti_svvh_generic_type of msix_table_size : constant is 1;
    attribute mti_svvh_generic_type of national_inst_thru_enhance : constant is 1;
    attribute mti_svvh_generic_type of no_command_completed : constant is 1;
    attribute mti_svvh_generic_type of no_soft_reset : constant is 1;
    attribute mti_svvh_generic_type of not_use_k_gbl_bits : constant is 1;
    attribute mti_svvh_generic_type of operating_voltage : constant is 1;
    attribute mti_svvh_generic_type of pcie_base_spec : constant is 1;
    attribute mti_svvh_generic_type of pcie_mode : constant is 1;
    attribute mti_svvh_generic_type of pcie_spec_1p0_compliance : constant is 1;
    attribute mti_svvh_generic_type of pcie_spec_version : constant is 1;
    attribute mti_svvh_generic_type of pclk_out_sel : constant is 1;
    attribute mti_svvh_generic_type of pld_in_use_reg : constant is 1;
    attribute mti_svvh_generic_type of pm_latency_patch_dis : constant is 1;
    attribute mti_svvh_generic_type of pm_txdl_patch_dis : constant is 1;
    attribute mti_svvh_generic_type of pme_clock : constant is 1;
    attribute mti_svvh_generic_type of port_link_number : constant is 1;
    attribute mti_svvh_generic_type of port_type : constant is 1;
    attribute mti_svvh_generic_type of powerdown_mode : constant is 1;
    attribute mti_svvh_generic_type of prefetchable_mem_window_addr_width : constant is 1;
    attribute mti_svvh_generic_type of r2c_mask_easy : constant is 1;
    attribute mti_svvh_generic_type of r2c_mask_enable : constant is 1;
    attribute mti_svvh_generic_type of rec_frqlk_mon_en : constant is 1;
    attribute mti_svvh_generic_type of register_pipe_signals : constant is 1;
    attribute mti_svvh_generic_type of retry_buffer_last_active_address : constant is 1;
    attribute mti_svvh_generic_type of retry_buffer_memory_settings : constant is 1;
    attribute mti_svvh_generic_type of retry_ecc_corr_mask_dis : constant is 1;
    attribute mti_svvh_generic_type of revision_id : constant is 1;
    attribute mti_svvh_generic_type of role_based_error_reporting : constant is 1;
    attribute mti_svvh_generic_type of rp_bug_fix_pri_sec_stat_reg : constant is 1;
    attribute mti_svvh_generic_type of rpltim_base : constant is 1;
    attribute mti_svvh_generic_type of rpltim_set : constant is 1;
    attribute mti_svvh_generic_type of rstctl_ltssm_dis : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_1ms_count_fref_clk : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_1us_count_fref_clk : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_altpe3_crst_n_inv : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_altpe3_rst_n_inv : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_altpe3_srst_n_inv : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_chnl_cal_done_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_debug_en : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_force_inactive_rst : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_fref_clk_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_hard_block_enable : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_hip_ep : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_mask_tx_pll_lock_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_perst_enable : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_perstn_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_pld_clr : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_pll_cal_done_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_rx_pcs_rst_n_inv : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_rx_pcs_rst_n_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_rx_pll_freq_lock_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_rx_pll_lock_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_rx_pma_rstb_inv : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_rx_pma_rstb_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_a : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_a_type : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_b : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_b_type : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_c : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_c_type : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_d : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_d_type : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_e : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_e_type : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_f : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_f_type : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_g : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_g_type : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_h : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_h_type : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_i : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_i_type : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_j : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_timer_j_type : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_tx_lcff_pll_lock_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_tx_lcff_pll_rstb_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_tx_pcs_rst_n_inv : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_tx_pcs_rst_n_select : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_tx_pma_rstb_inv : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_tx_pma_syncp_inv : constant is 1;
    attribute mti_svvh_generic_type of rstctrl_tx_pma_syncp_select : constant is 1;
    attribute mti_svvh_generic_type of rx_ast_parity : constant is 1;
    attribute mti_svvh_generic_type of rx_buffer_credit_alloc : constant is 1;
    attribute mti_svvh_generic_type of rx_buffer_fc_protect : constant is 1;
    attribute mti_svvh_generic_type of rx_buffer_protect : constant is 1;
    attribute mti_svvh_generic_type of rx_cdc_almost_empty : constant is 1;
    attribute mti_svvh_generic_type of rx_cdc_almost_full : constant is 1;
    attribute mti_svvh_generic_type of rx_cred_ctl_param : constant is 1;
    attribute mti_svvh_generic_type of rx_ei_l0s : constant is 1;
    attribute mti_svvh_generic_type of rx_l0s_count_idl : constant is 1;
    attribute mti_svvh_generic_type of rx_ptr0_nonposted_dpram_max : constant is 1;
    attribute mti_svvh_generic_type of rx_ptr0_nonposted_dpram_min : constant is 1;
    attribute mti_svvh_generic_type of rx_ptr0_posted_dpram_max : constant is 1;
    attribute mti_svvh_generic_type of rx_ptr0_posted_dpram_min : constant is 1;
    attribute mti_svvh_generic_type of rx_runt_patch_dis : constant is 1;
    attribute mti_svvh_generic_type of rx_sop_ctrl : constant is 1;
    attribute mti_svvh_generic_type of rx_trunc_patch_dis : constant is 1;
    attribute mti_svvh_generic_type of rx_use_prst : constant is 1;
    attribute mti_svvh_generic_type of rx_use_prst_ep : constant is 1;
    attribute mti_svvh_generic_type of rxbuf_ecc_corr_mask_dis : constant is 1;
    attribute mti_svvh_generic_type of rxdl_bad_sop_eop_filter_dis : constant is 1;
    attribute mti_svvh_generic_type of rxdl_bad_tlp_patch_dis : constant is 1;
    attribute mti_svvh_generic_type of rxdl_lcrc_patch_dis : constant is 1;
    attribute mti_svvh_generic_type of sameclock_nfts_count : constant is 1;
    attribute mti_svvh_generic_type of sel_enable_pcs_rx_fifo_err : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
    attribute mti_svvh_generic_type of sim_mode : constant is 1;
    attribute mti_svvh_generic_type of simple_ro_fifo_control_en : constant is 1;
    attribute mti_svvh_generic_type of single_rx_detect : constant is 1;
    attribute mti_svvh_generic_type of skp_os_gen3_count : constant is 1;
    attribute mti_svvh_generic_type of skp_os_schedule_count : constant is 1;
    attribute mti_svvh_generic_type of slot_number : constant is 1;
    attribute mti_svvh_generic_type of slot_power_limit : constant is 1;
    attribute mti_svvh_generic_type of slot_power_scale : constant is 1;
    attribute mti_svvh_generic_type of slotclk_cfg : constant is 1;
    attribute mti_svvh_generic_type of ssid : constant is 1;
    attribute mti_svvh_generic_type of ssvid : constant is 1;
    attribute mti_svvh_generic_type of subsystem_device_id : constant is 1;
    attribute mti_svvh_generic_type of subsystem_vendor_id : constant is 1;
    attribute mti_svvh_generic_type of sup_mode : constant is 1;
    attribute mti_svvh_generic_type of surprise_down_error_support : constant is 1;
    attribute mti_svvh_generic_type of tl_cfg_div : constant is 1;
    attribute mti_svvh_generic_type of tl_tx_check_parity_msg : constant is 1;
    attribute mti_svvh_generic_type of tph_completer : constant is 1;
    attribute mti_svvh_generic_type of tx_ast_parity : constant is 1;
    attribute mti_svvh_generic_type of tx_cdc_almost_empty : constant is 1;
    attribute mti_svvh_generic_type of tx_cdc_almost_full : constant is 1;
    attribute mti_svvh_generic_type of tx_sop_ctrl : constant is 1;
    attribute mti_svvh_generic_type of tx_swing : constant is 1;
    attribute mti_svvh_generic_type of txdl_fair_arbiter_counter : constant is 1;
    attribute mti_svvh_generic_type of txdl_fair_arbiter_en : constant is 1;
    attribute mti_svvh_generic_type of txrate_adv : constant is 1;
    attribute mti_svvh_generic_type of uc_calibration_en : constant is 1;
    attribute mti_svvh_generic_type of use_aer : constant is 1;
    attribute mti_svvh_generic_type of use_crc_forwarding : constant is 1;
    attribute mti_svvh_generic_type of user_id : constant is 1;
    attribute mti_svvh_generic_type of vc0_clk_enable : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_buffer_memory_settings : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_compl_data : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_compl_header : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_nonposted_data : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_nonposted_header : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_posted_data : constant is 1;
    attribute mti_svvh_generic_type of vc0_rx_flow_ctrl_posted_header : constant is 1;
    attribute mti_svvh_generic_type of vc1_clk_enable : constant is 1;
    attribute mti_svvh_generic_type of vc_arbitration : constant is 1;
    attribute mti_svvh_generic_type of vc_enable : constant is 1;
    attribute mti_svvh_generic_type of vendor_id : constant is 1;
    attribute mti_svvh_generic_type of vsec_cap : constant is 1;
    attribute mti_svvh_generic_type of vsec_id : constant is 1;
    attribute mti_svvh_generic_type of wrong_device_id : constant is 1;
end twentynm_hssi_gen3_x8_pcie_hip;
