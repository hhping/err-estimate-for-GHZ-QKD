`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tXqnX6r65G2XJlzGpEX5zWBG42bFx35+M90XEQtMSqdKwZPxRN0/XOtgBI0us0TS
OBFguq9JgrN8wz2hQem8lHhzLgEVuMHktNnrO7seY39ndhcYAc6IJS8zZNcUmETr
M2aYnPxow5GIegC3xwF8M7mrnYaKABbp9Tyt/quro8YtNJNa1faCfJeAlmZJdbZt
ICvyCTmjS/T8ZiRRI3e5nDBYwhBtCTRzsGsURfCEs4Hcucy6uOdm3PrabEDf7gY1
cpqGX1rWtX9MS3vYZaYyKbIXMqrYr545B7/5k89cB7L7NPLoUkuqNchE7ihFDbPR
ku5X0YEJvE6SFzr4pw2t72rAaWv214vXEVGbCdKyjHDHkCkikQrjWwfRH0osw8kO
LYjvWdjAFptT6CwnyujJQy58aolr9XlaBtdoZroZeFnNx8WM4X1f93z6DorEWJCH
EJV/24zoH+ul368Tq/eoZ+h+SC+eCxFBnfIS5hmdgCVReuLBwqjqQl1PjBF4S0Lq
lSR9eJMeHveX14yyUYzksvSTkUrdh6UOJEwMr5hFlLOXrbWCogJNMRjzRk2vAdVR
dgRMSZvEVIdlPZuCYqkt9hgT01hxCjNW3aS483yP35im7FqL0T2l48xKNt5jRzn4
h+BX3C9vH9dk9/pvhYw+aTf9S0DQMX864zXgd4pV1neltf/3rB4Mj7O2Z8alXe60
tYZpBEEtLKWCaWEG3PYOb3Jyrrr5fxqeB6bJOQdx+gZalDTrfn0iEiCvUZz8fNbC
z7vb1eCm8Sw2qbhj67BrpnX+OmIlyrKu+UJa7wT5QxdhEACNIKXAQW3XkjNLFlKy
o/DpJP+0dQuo16Wbf4scPuhnUoYOI6Ey4UUvYFQi4pzkH1pIJlJvmEf8rlhefuUw
HqI1bgzyvH+Ng9YFGnRAYm9Hti7xHehzZnRgCfJVxSRvNhMd9aRp4oQVxd09aITy
ZSgEqD3kBVmgqyPEY1U64HuEk1rDAeFVckL+u5FdCj4ULi/hVRosblywQO+QLqJ8
E4p50OX+O/avKm3WisB2WqdxvaBPR/cQoRJn4bskvEgaDmseszYp2SJKO5H9bum2
vOLmhqh5dYLT7zPy7K3aQ4tSZLD3+RmiJsz3yDONVWukGEyzDL5BJIA6qb4qKtqy
iji3WdH8zoNTKz0D+Lh+5Icq9rXYxQczawI24YgaH544BiB+JkDunAOFHn427U1u
diBKrW94JTSeAsmqjWckYlP+2tD6qgW9rWUFJ+W7iDDNqQLMRkjhUbzsT6Q62JlH
UweOfYL7RBwOpSAUy0Rq2truQOk3byeXKIxf0W26yO0ESTH1nx+VbJQsmeUlAb9c
OkapfMQNgv0cuoqCUnYvPn1y3z/nNqjz1/YSI+x9A3KYg1Qa45Fm3PyL5YSSfSaq
oCmwCvh/HdKLpL8UHFb3WDzIDVHU0qqnoqXTAYhMs+G38+a1CC1k4ypN9qQSQQJY
ZKcXOQL86lz7uoH6tga+8460RXt0gpU+0JHEjIKDVzmQUGKm+UiMkeDsPWFGO6Kk
oJ2Wk/8sETvIyUQegpsQWlA86Ra9Uf/lnrjWPj7oqykUjBtIMXNwatI81Rq/Drlt
enRy4K+4NDM4Vc5E8sq5LLAJDeFH7gdjYmXkamQYsREUCOqrTRt7CmimT2S2LvAr
O9ChA8Uy+URoRG6hZ3eYcBVAa3IUOD8SmXyoBhhPcsiYU0IvyXS3+rDcesxQnt9e
tt82IQDl+/R74Ds7NqghzVM0tFBCQ30SHoM0G1WFHFq6AHp8STenpuisY4w7hp5L
hs6L94dV5jH+7R7s7fDYslmvGehKBT0aUf6r1y2DijSZuMSXtnOvQW5uPEu8CAXg
TNFvHrVRgfi8N9pbSAaJfwN+huYxM5yxCvTJ/BlpFgxy/tWlpd8W+VHPb21YOQsB
5UZxgOsr+mEXDmlBX2obZoct/pUlTH7tvbohcVw9Kmt6Ora9w2/gzOY9Cpy6EahG
F4XBnmpGW60v3bs+EhJpZXhyD3kO5d9gI4uC8ifWQIlJJdvb0Sp71MANeewRoYW0
ErFCaUh/UBdC8qdbAiv8VUk+q6FAj7o0taRhfoHpkU21x6HSqrKYXDFdJGssDZqr
I448gHc8kM+svaULhJven97OmVjuU20DiUdBXkSvHkfGPo3h5dQMi3TwPBGQrwk6
IbYply4nWfW7bO6xGULpK9foZUafqDMDPh23vRyJgNB7zLtxPrp/WxXIZ3TjHiGg
5gziKny+otsgg1NzwVfw+BeJNSjOrUXLZgdMGvQ6WxYrqxCghjxUvBM1sNVKHbUs
j9Mhcvk66mdqRemgNMswzYTbr22PZ7iQVH9N/72AOq/2hK8/NZgKIrrw8vk8fVhr
r+RcrZfblZPXoNAJmK/F6LR4lW3oJOA1y5/FO75mWGy2UV2qBWbdWeNXdVjg6wRe
y/cu4SkpFM5h6tIUJi9i9uOODweXYa/O+ZG7d0PrIdwHO1LfnW2E+PRRFOjLZY35
UHpeWyj0V3W8r52M5joc+RVt6ckQPbF819JJjDg5SDBipITJb17JOuVhsDUYTbes
Ha9oGBZqFzfUMYLnjhCe/i5kHhGAmperX9nNkKlcpW2c0aBz7YkdRPFpqjbIrhmU
wVAodLS9sYgCR3C6NTcaXRqUOrRpPGcCRHXsqq8URtNBq6NOMtoET3YeYd3GnUZe
PU5dugjyPv2w51Skd1XbpRtIJA8YF8hZuVHxwyUXK8pGgoHqMRyMJXNOoE0jZNUr
VPaw4Wg3lvrxhHBtshjxmcwnj06g9TrFz3W7iFpRfQWzzAzz0bzdk2HZeoq2cHQo
+jy/JvH0A+O+2s4ANXrxGdy/nTcFiWdxcgAMxnpkSdUiZeQfgc3wQs4AhyGuMpSb
6vyhYdQwTFDENsngLWRD4oErDu/1whkofGiRqVIGOKVOg5VqRLKqyOdae7WdTYJ8
LM/SmbD6JcF3Zt/Hg4RrNsdiN+5RBly5yF0x+JliDM2XzkV7rbpF9oXQFTYxhBG8
9kSSyNjCbmhehWUUmIo8s1hF3sWASi+9v9RaMSkuuMNnLwOaWYbzvBbotoRj4agQ
OCXJItjt4j8Xj2Qo2l0hhNdlmCxR4DQJ531SYWV9QEv2biAvgsHT39kslqILxApg
c4/URqNq1CAEF+K9ABnKxSIhLthfK774Cf4my3NQsczrdCkMphFYJG2xj4UP1HZw
5zj0385FjhCFZi2LSZU1NPJaMObvNGPJRHs6V4saEKZ82TZe+RTYc9XxXg5LnINN
dDmNCdOrpIqyFvvt2QGk/hC0zprh8EAPYpY9WJBt7/loCn092UNhp8X7msJGJ/LH
7j1W9c3spBAqi3IkQ5Q+XTvn2e0PiaJAQWQiLykbop6msE85/XbKvaRz8uVaOfJM
R4mPQw8zfI0FP+R+dRladjQeFjdWWbyYcSp7egGzqm1S80zA1oUFLTEOioC1zQZ8
kJS96bVAGOqEe+mr8InBdDsZzc+3AGtb3DPm1wIh6Sf0GGN5TEQSjKWvUxaSOCT6
kIS5ChVwlMT3iP8Vskg9IL80QXb4IPNejrB9+rCyOTCoi+XMFibYm2KAV9UB/kTW
zmmb085xXABPyTaWoTA319vscM5bi/O4ngqM0F6pf/Lqbfr/huMY6eg0EsEg9Mz+
MuGREEXCroXevRKy6+7ANYCGWzWojbbwf1ocBs+RFUYMnwY3ytpihutF8kotJfWt
upcUPgqdYLM4x7//JXFswzqc54kV+ITnQet9Q9QA/y17T3ySetfYMSBOAmos7RwM
Q5IrvkNVGki0b13tArahxiQuUkUvgVPtL7wgX4aqPnaQKSWiOmouyWI0r5coEm6Y
WqshP0FPQ4/ju14T93yapqEYmZbax4agPf8jkMmievCcnn/YPPceIsTKYNBCLf/W
EQVSTPvvAEANVf7lM2RTzxtAaj2aUNG0usYCRbi805cvePtvndsuXggmfeH57+S3
P6+voGpEsez+3aE6pJgrsQs3NqX1hh/3fqoyj4kajRE6RiCwTB1WjCUbZ30mHWJI
MA98FrLqfrbZdO49XjgNEeCpQZsZ/cEtkOAUjiV5uar2HgxArGuGdq08QO4hnhTm
Rx9AFNOb3ZEsn+imMGzvm53CU+GFDTpFVAYp9lzNGcyiU3u32BCObwKOFI8lKP9N
YBMw0N/H81OeGHdAHHT7oWwWPArPxbvckNnhdCxLV9d031nfOTlBYeqaojwzeKii
pXMIhO6T+eSrms5EmXr179L3JTnTriWTt8ffY7BQcXXJYfbikxo4+31MFAmMzrpB
5WTD3FvMPg0A0ZC4vuUlGHiJICw2lvQJHCeoumRIJ2IPCJ3+DsQu8zdIrxyXeP1K
1lV0peFfCjT8YuYsdX10Fyr8GeTrXoN4XcTb9fkdNhijjklIAVG1l9t8qLEK2AHQ
I7MZk8Tc4xBxRYl4+DR4I2sZLOiE1Omu3fOBrAN1VSEHbmL6apSjqe71enDOqFd4
NQJcJMITPhVJ7qEleJ8vx0sTnJI7s8D8J9XdAmwU8AXToqt//J/7/oTIqXaj74BU
99bmLuY3HY6KgPN/JnK8jA3igI/2hCs9nTAkQf9cBi92i4qcS2ve371cLa5xN1o0
+U6Q151NNdpN8BWdQgM8TDt6eW0ZQHwWoXbsY234P4N/qWbrJzy926zpuDnFk6fL
vLPbGFeoAGw8xPgcBvgwe0oIKHnEgcSwgOUWF6rArtIo1QTKvKrIinKz7LOjHhq+
dOAfKjDTA8FOqKzE93hfGMwyvndH4MK2VoCqY0/gfY/iL3i3zZ/LcF3OxXDGocWg
v34bjk+JXxpe52AoK6SkUFCWNrF2KuRk0KOFVlumEakLkNhIvq4k6JWod2wb5oU8
VoNpRX2v2xUmvkVNkCi7zL3cx+mccK/d88NEQXrRSzoCSR6wBinvpPAjcw3hwvt7
Dtzw15m+EfFosFAUKdjXPxpGARFGq6ogIq4tI6WGwK5QD1SA9+pXEQ0PkmYJfTUU
XepKw+FJ++cYxyot474oT5f0FmqT4K/8IR60ItN5RKSIqXMkDfWkAxSMMbzaIEDa
83DDIgA/OoCnSUWWPwZ3r/ztlId3Y7y/BG2U7g8XqZCFvjYIV0At8ssHtf+txcXK
nbNKcSvHMzWtY2TSqzYXlxRkiT1Nw9gpDxBPTJEc40vRH+oiVnyXXTcKPvyZSxc+
SEh6IH2FqBbFIPICQD5ee7TIzc8vE+d0j8Ld4YqkLyS+GXT02WsG+dik/C3xj5GS
jq6xBfufZ0zJkX/+V7AMby4yNE65AFijf3zXiSWE8G8LYSBRyIoWL4sIB5Q+DbEJ
uEqKK+fPJiTS+an3RdpFxkQccnJDbdjzvyDbkAjVdfuwtUBknIafxODVJIfs1AQx
Cndx7iUtvzQGx3RkbmsvZF6My4hdNnnSzhsxH1KNBqVsdbaoknv9ZAqB4tIKo3CL
UeuZHaRdbTg2aUfUBE5aED8d4mGjKcAcCXbNoP3+GoWpZfk82Nfo+eH7W8QNNC8E
QGehB1O0YVRUFeU/+HgA1JlvqKvS6MKTdetvigCzGJnKATPWmZ0BnfSo+htAl/2j
AFKbW/b6bDv2DnuEk+jdaFpXvpSgIfudh1p/yXPEr6VQLb+MBx/70JN0Qmu5HTqT
`protect END_PROTECTED
