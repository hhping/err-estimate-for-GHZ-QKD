`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4rx+yWag3mBsSAdxKCQbBBeq53PzVJ1Gl7aql/K56OnUSfKWnN+5D0wAqqaqt8IR
zpzItu34Yn/xQ/VEgLJnhwMl6K+uVZuew/tVeevas3KrmryU6dYavqpIxEIIdA4H
6LeyjYYzj1T6/T8QFaUBfQof8l0VPEMUJHgg4HjXpi9/MGpUMNj/VvO3rjofZ5gH
qHpgniRp/1cfDX+/fVCftkoZokS+hI+KManu10AaF6PGMf85S4udvG4PiVTExARK
hUJmlGSJhTBkONy7S+brUqZBiMPEtAjZSuS9QkPV4TSqtCtzghC/rj4c3Gf1q4GQ
TxY0h2scAK5zDaWvFL1t9seMO0Wl6PYzVXoO4TitW5gmxlSvhUwniAGx33yrnRBB
pmdnGJiRk97qpIjunBd1zVDkM+JUJ0RQTlgdZA8K1NLmlDnEsebvuIZmeM5lApK4
D+kNY0+gWAnYnbCSdTr9yI4CE79VUncF0lAHaNx9C7kac6wnj7TdKZiX9NYoXtHu
4s0ZyvtLrWlHBd345kDdh3ZyGxX2Are7ES0fDhTC8MU=
`protect END_PROTECTED
