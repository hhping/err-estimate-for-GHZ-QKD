`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kuEU7BIii5Z6TMxG9M/04bDD5xh9UbIDqdPyaWcnTd2Rb/haosQ+/fZlXCtFLQGP
NlWVP07G0yrYsz00aSatD4kjnhAV62JjM4r9l3VdVitHIMATFIFMfaTgA0k++UW+
6rJo/g/rSE1v30dAv8iLNmVbVNx35z8aVcJBdxggQ9wrrb+LJ1bloTNQUl5c0arZ
HQGz8B6fiErzBnDoERRAI1tZV71iJRfSSMJcD/JJlU+LKKMhQSnHgfjGqQUIQ+iS
GLfHlaLXmikCGP2u7aAwsfpcwFWwcGir+ak1vSevMwYFEiozvIepaW7nINZg5sFz
bvUyIJspcirtcg9p//9er7TKVI0uV2duYebJLKSqbzC8kaHVZ1bYikImlr021wSg
YYJk51i3oQYOKl59BfIKwrNKvWTqBmj7kjqRpQUkXqZzq5Tp4Je3qRCPCjUw+Xtz
1XlpBaFlAIhlt3xCDTbL+wIVRfO/GINaEB1cqrXnBKPht4gNTjW6rbDxfN9yUL0i
c8bFdEA0IkZGrBBRYFBAAVShb8jqrse7251ie7581y6U5IG+5br/j5Op0Bf04DXT
jHvcyLpADfwhvQWid96eYaa4WUT5XAR50cXafDNCjKfgoXQz7FD2mlGSzpMIRwM7
joHn/A4oXWIeJtBzwHkMcIs/DSDo9zJUiLtUwZAythbmeD8n80N0YB77twBED/xe
j1FW/pl4ID41sQ/BNb/npmGDCjdeuDbWXFbqORfTsIJe3VWfhDW4VE4eMEziiDA7
3kirIP8/1Yv7Evmq/Vdq3sPN4rOc48jmxYM3jkbEZq2KZXY6zJkINktOM5k/UdnH
dq+VQbLXl81uXD4t+vYtA8llfbnEvpjy1QF4spH30RAaNELxOBYmjd0jtsivSdKS
DX4eAdw3j6JJGde8VwRrBVIV/XD7YUItzD1rtAiVpJ0UYQcJI7L2AM4a/amozFHU
iOU9ZNA+UNVbXW7w8Kg94ViMKbL5fSedtAMC7OaQZbojVcpMbHVF4UpFq/JOj1b2
zQTBefffeQp4zVzl1sOrZBifmQBucnxo/w/DxsSvAXHXNFSD4g7PF0GGsmoVbAH+
HVRSddNxGTX8GdolNcwfT3ncWoGm2xJWTmqwtsH1uaNDvcTKlYfoZ+IG181SK/m1
TMdvBoUQCggfs84vh+N2sD30CcexMfExDF0T+WXlljX3c7WwyLsk1YvIIYpL/fZu
FqUhOUd49/JVFOzLDI6pFML7va1SLQRAchQ25yKIM01hXRPV+wHpFCd/2C9ad37z
zHrn3a/e1FESdf8mEVn7gHAjWt+crOsPln/5iiyA8gF5922K51Sopnfz3nGS0US4
w+7SuU3OjrGv9cD8IosqK8RFu8yjWD8e/K/9UlrZY3f/a7rGfDWtOkLF5I39ATed
Wnf7C4aQ1TiO0f4q2Y+Xq/kDRJRIeNjZrrLLKOq6r4UaKOvz0Z7d58ljLqgRl6T9
gqvu7YVqkjWYGSfG0y/RJGilNtF/Ube6UsMWseHGiZwB8rCOVtnywxOQNgBMwQFC
UUNU9b2k8yWnRWOLyxvEuoLZEOO2XxzSYyIvl1bZoceWeE4F2YxA4Fh0vutS+m+G
ChTnTP4gHPNSyPAWCSOQcel/xySU09TgXgnVZfKFfRYl6EgLkbDSnamW2LsRUfFR
qfmVkZr1q07hCvtzvIvUFmI2OBpdYjtiQFCQnun54WGGWtVK+r0Xz2pz90ktqF0M
aVbcnEQmABPlThkbwMFE6ZrFMymDO6gFq/dQ6vgj+vvrYd6YDHZQWdG8vIX+MiYL
8c0WdgaXnI3V1wNm/J69Nw+bdHjJU4OJ9xocm9wHe9o7l/hqR6tt804tmxPfH4Rm
Bce9lvH1IyVKfDuc9NLSre5qrA6YOIbQgCtBAnw1s9Y=
`protect END_PROTECTED
