`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
StnEFe3+l/drgT5xifY1s5UpqAMW9asm+omtNGVbmwLEjl9QntgWDFD9ScBfvFr6
jb8auo5bJlZsHPWqgXBlcLsUHG0OEucW3nV983mzTFH/oKF2hzXX7hc3igGC+g+/
MrW8cmIZYQHr9WLWiYE83QLc/K3o8QeoHqSB/SHYAiqu/5ceDsUGph/YEidjGIKm
I6hRyIbaCpvyTpmPmxnTeAkBH4/hvTEFZ7RxriFQtSoPObSvUFLepgqhn+bxuWeB
cPhyV5lObsjPddDsi5khzgN7hxYIPm1i+M0MpnnKmt6Ee9zX9rKpW6ix+lrIK+R5
uph9glOgf81aPKnV6mWSgDyf0neeSjSWk/heaslRy297TktTQ4URipyLWovRXooe
dK/U8E1UsD0hERsnWCUQ8K2DtgUb23/xEIEH0DJPmbGQBxaHXqhWqtBxEWHboTbE
JzsgnH6QYV0O8keneYB8kGI9NsO2GIVLQolaFkwHYeG3gK6n1s0ADPPEjp7K3+L2
`protect END_PROTECTED
