`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AW1rDnBLrMiAVKny3XUM9BVbg1Vz88RleGBgPZll4XYr5ceWUu45ygb4Q9M9EN8X
Jh0eU3O1ToBPU9RovLkGESzhfJlF88eWL6DQvUEKbzhGyjtCIOzIVi9E8fO2eyhV
tyLOIP9yPDjHV/oyEPgxTLlZ2OYCivMSUVE4Bv/+B9huaxutkZnrSmom0KY94uuh
2nNUjQW3uNqjKo0Feayg9oWKW9b7r4osB+HhfPa5YzA1jFvCdoNJRS0apCrmPVks
7FAQM4mrrADn5laByiYberuBFLgZnx1St232sjy7H8+6ZNPOiucfxfzco5rQYnKa
Y8k5HOuNO8N8I+4HCZvQdZrzyl3ubxgNE5ZbsJlZ8KLKDmma5AVIeYb/IRutx89e
M+OdNYyn+bsBUj836DL0R7ya00zTY7hRmtCtHxH0h7x4QjHWwBiUxEIXcaT6XqVp
9850oDEA31ufyXd+xrTU8F18v8deH7kF7W368MyWL5u4QLUWdjgbv+8k41w7cSyo
4c6SSa8cl0ZKhuAvKZCArOmXh8JL+m01eDQ2KZe2SjqUmFe1AFlOfYR0ji2zc7BQ
wz+Kl76GmJfD044W0mxsOZdYkvUcjJBH/6feOK+b9g7n5dXBtkg1IHJvdqNv/uL7
ALBZ7tB4YiB0JQra2ERJi62REU6M+xwEPtu5uouRHRq/ywGJtu+OgfUnHoaGISbC
u1yHZ9MijKMFSzoXD2y7AX/27SzmSnGtctwcO+A956tYOI6ImjZNutM7f2ijHIxq
9yUSLUQliha/LOT/eeZyQ5wyQCNhmIZedXK7Jz5xOdho7uoKKlLsQ0YnXhiH6tUI
yF4WIlOdEA9KM5ak7X92951Vmlo7xYN1psCgOK5DY1tToTQPjqDFtwupIAYYspA6
cZmVifJh9VY0j7bdqbsHbsP+CYQGI1LGNW+Wx8UxewAv4ukX/YIYohYMRvl7KtD+
RceCUgq/ZuB/IfRk3Kcf+vkmOfpb8q80azIi1NbAKtCEiDbf8EaAvDfKJDNCbpZB
X6YmxPs7R7PU7/sBTmz986ilIUc6TIGugPCLn0gARbn0s4KCSpWZAop8ya8cNJ7v
teIJrN3/FuC8TmyAmaQYUdS7hG/cnz8ZG8SZa/Gn4xDxgf3SjaZp7iUHfqN9i87J
rcaFnJGzO6JrwzyINwL881ZKrK8QU9YW0QocDP1eXY7nQwlkWLznN+BLx+G1U7Cy
isz4xjpQmfKb1uwUzvuLtRJVgEBdVk7aIHfsUxf6XUVvTfmoQ0FTS0hjTE/TtFu/
2E7A+qTDZbzxUOk3wA4W05IHJi8hquLTCAxKHwkiTJZgJhXgIRwFhcso/Is3BtzD
oArVUtNdOHIxmqNdus1yWFGu2rcMyCpBkEDnyKqwYycQxmIRZcnNUmk3yK1gBoEJ
k4ZjEKjzyG4+cmdyuTauVV63NgZ91izxwg66an/ZSQdakrLq5z4ah92gC6PemA3t
p3c4cMywXkAvSrwR2MF2SM9XpRXlNqM3ooangi0NpFBHloHIENrUGAhTdaJ6tVCc
vWIby5YuRLlIjnmFMy6JL47lDpXv1J5fO4dKjga19qK3dpWVEUf/opdwMm/gL4GZ
j5TKX9JBshjuwvcYm/xm2jWv/Efwb7E1eRyuQbWNmCZ3Ux2HNyZQFqXX7/WfwLbY
rE0vPjcb1WC2H9hP1DDq2PZnGrM2gOQiB6xLVuzFcBRZ2H5xRlPrlRI3LJ95676T
5I31STFtuIPrFl67e6ISp2eM+LSpl2Yo2AfEGJa0TTN3Zyept4fYcTHpEsj9C8O2
jTx1U5VZoGYDOsdlD1NTtYBFQn3Qnl6lfwX8PfCNJF66nb1TpCCe0F+efJurrde6
C5enOBGXTbAUFnQ/s3RcUoL/qUPFodhun/Xf1QCNeVP6Nw2yo+gvHrxnGYM3rSf/
HuV0i16hv5e1WN+zdBw4m2k9wz/sn6G5yv1US6goOYpklDZ6LXPAqVpqHDF4XIBz
C1dP0RVhrIIdeX92Pst/zU8qV0uurcIIFKXm6intKLEttazPakwft5CxnBBH/1HM
8KySf9YvwKS0ZzlMleytNt94tOKRE7FEOUBOxAsrE2v6GQl/U2YT0MfwW2Q1f4k1
HeAxIDb/kaac7vWM4zwvrxqrz7s5mAXY9pZbK5O4NYK4rKchcMSVSzO+4XLNdVcd
k8hayjcYFt28bp4s5JXceIoVoX4wvVFzh66G6HohfW7NJ2RWeKwEIj/RTCi+R6Ar
uU2QSU3fUJUF9ijVE2NSYrOAGrxucAuKM1nQ7BMk48QD/4QfX3l+kUf36aHpKZFH
hoO8HtSnCcJ2PqdYlvagKeUceaL3kGFbyaeqs1gyl/BCUVUpM1D9Ju73daCrh+jX
6QwmTLDtuagy72ZX79Toltt6KmJFWp1NuP6oabfhonF3jdV7gpvo6ParxnI1eEVO
GRsWGYej5YxDU7Z4OtiTNUvsFhY8HE8hJqwHtfJkQqianlxK+7h7t5JKUFZRnGFk
QxFHyYgFvHTMvFBE6yzBk3aAhewnTn//PFxOLijIQYlZZBGvUat7kjJqE+PQ+n+O
HKlin+D754HuwRTszaTvwV7UV7JRdo2Mh5G/85DzfJPsTco9D7F9aHsePWxGxZV1
6bhYNSvS1+FHedo735MaM4NuG4rCtRtnFhIpve/7+lrKy9q7ScZhTRaVGc3YfFYI
yN8E5gHJoPk27QoptydA8zufCkGR90T0KZKGFbMhyzkBf5VjhR/rgRqni1dY/21d
2SW3xSHuM2DhTBGL2qZzUXzq8ah5dqRX5aOn6R0uKzszQAxrZSOMt8mcQulRThDI
ncAgvLM/d5sHP8478bvxx2tbPijsuz0rEBLOeGS/Z06ZhZ1um3z7UVT9sTOXGbuV
OYSxqiqOWgBTjpa1CYfg/1xsuLYMdQpZh6Vir3FGVVy1/02BLQq6DTHVN2wzuMWA
eAp3XDxm/KU6Z/JKP4+QwD7NKna3w5dKlswmW0UECe+guYZEEkmzHgTe3Yju0pi/
9coEwXa7EUabx/lKHJSh3ojBD5C1/mRAMR98+sHQXm4+olcLR3nGLaF9kTkKasLi
4xaZEvw3WK41hiTxxRhUl5Eq0kVoOXIwWhqzx8xSMAnN7WV6FKO36Xw+N9n5Tts/
m1D24+DJvUywOB+3c+PQUHLB7/vKGxsTr8JnTzy7YHAUjluoBD/8ajMZQWihy6iR
`protect END_PROTECTED
