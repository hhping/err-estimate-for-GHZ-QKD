`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dug4woJjguKbmfaezFvq0wf0W65Cy9QMGhCvAaqEDY91aVa92YBp2SpJO7KBQTTj
m8QPvB/vPPJpBq1hRQbtjhAVKEcISYBQN/zr2akaeamgBSpBUYCg4nc0z7CvN0ef
bE8bwXFrSvQp/d1pmxw1L52O7qF8YcYdRTGbm0DSuDbbX+b6PssQVeQvnt80qLVh
VY7e+w5BMj0Z6tInHw8mJDeYk9aS5E18Xm9iFxsvIBa9ab12BOsg4OuFEJ45ZVY9
97g4epQV4jAdAyZ7Pthf8IhcrGCCvgqg9J8Vff7SUYr5Bjs5tTre/34iuneC7HM7
EO9unvsaqQ6n0F0snq3WexBQC64bUyVBIjTqUVO7AQD73W2WTy9wwr0mjHBd/nD2
djiga2POQN5W30+fXm599tZZYIRuPcnW0r0RlABOBtLYQQa8ZNsTIX8AiefanvQe
Uwin9XPjnuGSg9Q/T7AUjBAnjCWk+uNnK5fHTpzeWEtJD5YKC7OY5I1CSQJFbBBt
lgw414uA4KT0ffWNTO2zABnLUNNPDKn9Cux9lctKRLr/kY+4gOqFdMU0SdLE2Gem
vhQ3PuvcXNUYEo4aT4JX6lZkMzob/6eqkr1gS8yKYy8xOVgW2KL6WwSHTKCwMcXC
+z2JldZU3RgsSlFI4G75LGgpO99gj0nioaVjS9D52A5rDF/E4od/G2pl7I1mXagh
R0cxrvtCiSCGdXqalZFRef2BsUgRCxCu/0g21eEmFYgnK8IHEytE6FbhxKomXcC7
X8MDhlFeY8w8pV+wCTeM+4ESuM5BMQyq72AMLU+zExFNSRoF+0wlYWW6UXYmVclC
QEK6qxKQa+kav7aJi/W2IACAfGLWx3soCLmX39TPjiqRvS9zwN/duogmShXOGCm7
gM5A6DTC5YWYjaHOfwtzmqlyWxPSycjoEKQYpDzqmvNWb6Ik0/qsdv023FiMvUbV
/7g4PRGkcmssX6Hnc7UZQYd/SkSSAgcMB2bHUdFeNrXXm2AzMdiEx3X23htSDZF+
q9/12J3VzoL9BdRKEHqkYkMtCiWHjxFSbMx5UgEthk4Y9TGLR66tMmAj/EZqLTVk
O0XydIgSMTlGbhNNw0pOafVEmvMB5L3KZuxZjfD9hauYhenrepPRJyvB5VWDD0sO
/JU5a1Xt9WW5BPwlTXkEhBBHy+9mJbTF3LyTFZ52xZv16GYduqLLAssYm0Tc1SQt
QzovFf771dXUo15WCt0wqi+eV6NbZm63UgDeI4B/Si37bFoyc/2ZKx7a6W30wnuV
+jjpL0H44onS6SjIvJkD648uJ8xBf+xHy/Cgifgaq1v5qZH5FoeBZWrXv9dVmcNZ
bNQwkinF+cgSVgD7WO/DGR7gy1lPb3sa9Hd67xVjE42W+W+bj1nhHv6Nn+AyPYB5
YH6QcN0oFWl93Bo2ouQ/Np5B2BrZRy9X+SOy3+ECJ2vCHGi/j8iN0ARyG80Ca0JY
46y5hNzB9sLiZysiskZv/V2R63UymmHrZIIugHSHIIlt9bZejHiTQizDa8muJzF2
XP9n8WWBEnSz8yjW6eFuaAgyQcpbQ4ja8/07Agir+VLunjkiKFvPK70UREaPI4yk
tJAQhBeo3ipGnepp4fQiBcNmIEqhaWLPlCeaxVKEv/QIrasmwtsHMa0ZaHnbdBec
Erk77ub67KWWkz9CqHDPE6DanyxQQlH4/jOZY2JMWo+8NKgG7lQAEuHG8lpiuk6M
9Rumjtfa2Oo9C5siUHZvxuDeuEasoEKebdtyDIv7ENUP8d5o6mI+jpNide/d0xJk
qyHKcoGGIvvmgnYvKAhBzKpg6nFoT+g34nVls+q1zUZjoBTtuQrAiYkDkuEVVBu6
y7Mqxg4UowpxRQqHk/Ti+feOqc2i/An7uMY+v4hm33tFZwlhtklycSOsTHG01405
WkfdEgFCE5tUlEke955aX7098Dn53E7lOPHHH8MY1KgO8pcEblaBrZt8/ZSsNR3w
VHmoDW6XojYjaPrZiEFp6qOzxWIEb9W30vnQhu5vjGv75kTnc6sg1mTCdR+QtXwW
gU4LVRls85Qd3Vt4MCMQB9eT3bTs5DWSDLOpi9zUFxpKxmYMuJ29EZHZRIqyMZVA
kJBCONUxnkrfRVpDX1FUAY8mHxOza15U5dhtsSmc556Ms8h89G86/v8VKa//3cxS
VP/DLfaqKQvfpkcTfvhXqxSFYgwqTaSTFlsiL67zKvOLo+FwYooGCVBY5PD83hai
JYLxu77boC/z8Z6erQa63yc8rcZOFr+qxP/eBH+AuGxxp7h5KkfLJtbf5Kldta8D
6E9fkJqSagkYdxVYRMEpjP+q74yeNjtDz9/MoZ9DCfKwpl9rftX097eLWnN1UB+I
YHBn3q6xrBzQt0CgQjMpakZHWSIeKdrFlD/XMEp7BBEvfPjal+DoROycCdsHdM9f
UO4tkcn1y4C1f+vb4kVQLk6EKpL7vSEtt/j8idGDmyKFTXJr2kbYZ9ueNsxa83TS
hI4dQnq3zt/Ws4z4X8Uq0yOXqwARgR4Y0VjdKnLZvbGq4Mb0Kkr3BiGHgrDZ6zPy
WrOvYk7wcG8nTTtXsa6tm/03XVnmvkYZbBrVWnWaHPAUrSTFZgJuKeAPENFfBfYt
y1lKF5oAlxwwUSrb2o/uF4D7BRC0thpk7UhoTcdOyisqVptOPZh0SgGKVaxHtnmq
MBVD47jplB9qqcjhdpcc+4qJFquEt+oDFbfVd35/+vqFmfQfAG97fVmq0u+rL6mI
7zGZR8KSt9Qre2hrg5p5WKdIqIUiz+WMUhf9qgwZgsdy1rAjjfrl9EeaULaA+Jby
XQaG35520zu3HldvoY46zydW8Z+wsWlNmNML40FLpTRPhOU9JK0kBTuTYw4WpMfA
1/ufutOeUBXE0eMT/THrwuHKLhL85AvsWKL2Goxm4MuaGmKJnwNAFxORuHQYWmjs
/HK+wi9Q+ZkMgLfQ86VN1gXoLLmr1aF6r6J16nO8Pehw5cyF1VVdMV4XVbHQYBrp
R+32qAT8CEmQhu/dNug3sZK1RnX3BJpkfCy6eiGZR7tWckcmJ1++VCCXbtayLr/U
TuUINHqNID1vLRSZ8MKFZ07T/HHLlhzJkGvRhOPJD8yGtgmddlxrGRdjPjuZNxl8
+2lnSimpnUh/CxnCgXmSoGW6Om5vKXa/wsUygE8jNIfqVz7Y7wdKk8GJitttuWPG
xfjtpAy38QfrXHuBIULMrgpSloCdtfog9RGL30J7eR3tmdZlE+rWGUDLUD+8iHZh
xlJGUQLfEibeRHzEcJovSvktq3cwdOgKVdIY3TUsj0qosAus0HXHRMUYRW8WFIWd
KrQjNnDmggIoHz3bOVWryDVfP4OxzZ+HiTLau8vEjwM7OCZC2qY8v38mqvzsXr22
nvmb5xUJu7Lsc8We/25LVfB+Dbi8sUf0aIayQqt2NbA=
`protect END_PROTECTED
