`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j7IuirV/z4LLOIycpOxzaAHSLei+DFGvROHXQiIUxr/fAHEG/7TvP7E/42rvNDmI
XFE4aHBQFIKKi5VnKbM/8f9ygNQ3c8QBL6UXH55IKLHQkVgP25R/1KKspVv1zAVC
WBmiH4SxQov4NPKdgiTN7kK8YLEgCjJMpXMQpi7j/aBQsm+2jFGRbGF+PI+vasB8
qYbLoUP4wR7yiu/5snQpuGRSvhFeGilRSuRn9cLTKlHlr/pN/PnKjCuSwueLCXPY
EvRFVrlP4HRUYxg++p3Z8zexXQ+3Lu5Wu1BSfvmwNImFDYEfTNXP4RXDhG1DuUfK
sWmZYpCSmJNN48JbJbhTev7djnvat0GlgI+uS27QxyHt93F+utDcIBAo0H6fM4uy
4HJIslYdanjacAoe5NQsh9wuVieVrcmav7wsuGv8f3s0C4GfJjfVN+5OfDcwftL5
0O3No3ipHXtBDkgHl+2J72IvGbkUBQMdlL+idFvFhXlUYQHQsDifngSngfjaFloi
h6zY5v5sTArCiGBficcgpEydC6vEBB67r+OpYxfqRh7nLvIPYqgy2MloMyn+yZS5
SsqixLubm/yrUCFA+MNRqrd86iS57l/ImSm/DKNHE3lJSmWtRMI5m08JqH5DBxkt
9VP0mfTpa0Ea6a56RdCG6QLcr4rAvBFu5W8YewXd/yqAIl+MWJsJgWh9rblj+k50
vF9KfRn6/B9SwB4YQ4QWZ91XZo/xFvo8CZAIQrVk2fISBDL9RTn3QqAJB2cDvOhd
jxd5CVZUmMdajPNcMK8+NrZBkAKi3pzYUaGgd5/4XsOMvGRIbh7YIaCzICquJhye
ee6g6/XOINeP203p3BNmurRB2vO9eXmjO4zfxCuDKGOL2CF8iHkB/4M5+02jUyT5
s6fdy0yJuELiobZpy92baBvanDtom/D1PqxvqPCsNyv9hTp4a1vn67ijHqvHkkKK
Tq79clJWThrS1ieJyD3SyyBaDGwp43A/fDaFRlnly2ijsnU72F7S88OLWho6PDmC
6G1QW8Zng78/DMGx9u6+mkbO0HQFG0MrjMGjGL2N2dgz0yj+Wi0Z5vUGavU78Ink
flb2kVUyxa0S2TGg1N9AYNJDmYLMnX+iZBdEDO9RBq/aZ0UAmMkN8NFDZi0sbQy0
NSh6fijuehaEuke/JhFMyFUrNyQowTm7vFllhbmuHwlpnxvviicjmttyxA5t1APl
70lARrLsCYF6Sy4AvmdW3Kv8AeoFkLYYVUQEoXzsXqLEpPvwU7A0BN9Mg8ybMVxc
cDhwWSmrK908KfftNfyrGHJdl9ftcXhv8F0mW9O0VPc=
`protect END_PROTECTED
