`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+b78bz9L3hZsGqt+STcVT2PD7ra1+Cvl/88l5Pyi9hq+pHaLeqGx38jp41oak35B
jdOLgZSHLuWeh2T1WbU4lLfhTOsZcMeiO6nP5+hLlhIswP7H/BsLdMrxjvz5fIhA
8xci807DfbOKpN2qJ88mXZNwDlu6s/IylGIXVgL2gkFMOtT87+e0McnJex5QKpt7
8xQKA+VLA8p5gi0DhPEWoaBp1IIjRm3au38sw5zEWj6VdYk+HYId8Ek05uWRgtls
evP5WJM3h2njDb7pdYYkDHDKxvoBNS6M/6bKhqVOAssoSQqM831DkHNqjYaziKui
LQpFVt6LC3Egx0hHYPL6QU9AyDDpkqDv49Whhdr+H7omsSutXMsRp4XwoIMp5kYn
K8fwi4zeD6KOadZytcGagDIUVX2Lws6qd0H4I4QoFBkBZta6sv3yU6FCY3GvUQYI
p328WHvlLRnd4lw9ZbrgDYBjLWuJo7R6jd6JhsZGlSkG06vl4l4B61sKeRXEx+5z
lz5YNro8cwMNqBmonc/pTMD8M4DBYcxRfYnMdDDijUXctPT7bMc84zYp3Z2HqCN1
W9lzaD4hbMCzgBZREMGSmUkUzm3ERVh+dR81U3h0g2JLLOjWbLE5rY7ZZCK29EYE
c8fjLVX8ReIBzAHUyOvMq+vitu/fSCi1gKdDCsXGwGfmOu0prK2mCDcBb02PDnM3
RDthRGWhnJyOs4LpGJ5flxIqtcp0PlRxSWs+L0QNUe8RGEJd7eewQIBvKqAAOjuk
GDTt9YHbyNd8y2zEl4G4EZnyiBYwonEExXiP4IzrRWvhd5TQ42xDB7dgVGidFssR
e/YOw7lfEaeRumY7baxShGefomSt+MF+8pV/6C3Gq0DEnNqCT+PJFAVzY0M+G3Ui
bQxrZvSwocGIqvu3xOgTGg==
`protect END_PROTECTED
