`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U7+04rK/XjoS4g3sKZGTQoirJIpLu/2HiotMR9f69qDj6wY5S8nyEz5OLYsAxcAN
cDQJFB9Mzx7rvPV7uXCctEgU4V8giuyH8F9fj18GJhd1em9bbupAlBA2Pa3JIxAz
kFZq8oTikGfyoFTxd3yZLY1gD9D9cb9ZWS2YKZ776jX3zTMch/QeGnnO+Q7rMluS
7g8LQJ/qXSWKV+cInN5pOQ==
`protect END_PROTECTED
