`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y3X4DVrXljGqRw+wU5V/XheghNZw0Cxnk8vT+WPR20IaoP8kqOD6chNgot4jO41Q
yYaCstPQsST3sgyUCODZCBewTpDTvItCG0gaFM3UkVtHxWMpCgpW8yo3BcIJbBor
qYJMGmEC8qEfUewotPB0qwR/KVY5eY6/rY8DnfXMQeT0iJ1l65lrBms9ZD00C5wZ
B/I63wz07rFGnL9FohDd+/gAYRZeq/fqIQ6RYxfhE26hNH71x0CuP7+ZE2+w3I3B
5y31EKGH//FZ2F7HCS3eqwrtuS4TBmEalcmldW9ZrUUylmBR+JGxA/Vp6DMXIEhl
tya9IbmKxF8gfakAueCn/zwhl+gADB9eLdMGtlWPWdHV9b0nVZazSWl7DUTc00wj
NT6rOYj6mEmaPrpz0wiRPh+Q8mFutTMf0x9FdOnv10t6YPLxVSmVr+nAGYvOTA4S
0za/0WGFIx9ziz4IBrWpfZsr4BniadP1Zt5URbG4rEmFyIvf6THzBKSCR1Y+SjhO
vKOKCKsgYYif+JUtNlm1zJ4sEcm9wsnseOf6dROYTkl2sURbAR1HMrmtMUlNfG8e
`protect END_PROTECTED
