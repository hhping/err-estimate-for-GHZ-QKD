`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+0+AeaU/9ooXnADMFlUeKUHDeLEtq1REFP9Yh2dFALNsXX+1fxBsz1ojsa6HtTxh
/qtw44xh+NQ6dv5V/jNljWHJCphwsAGI6weokzvwC8Zz5CAe+KvBd1krJ04GpCfb
WedF4Pn0gLg/khuwFiIjPtEYblXjQMZnZ+4GK29Hd+0=
`protect END_PROTECTED
