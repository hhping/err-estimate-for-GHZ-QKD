`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aQoQYMAK1ERxyj81oorAbV6Cm/wb81PZQPdR74j/8dHZQA2XDl83mEXVeagYMh7h
XXPa7h2EMlIFG6tsYKpTvIEkMcqZW7V3yiH9IUvlWz7ZGNDiXCN1oyY7aLf/FfOy
/PGQmcgUaK9G9ktvPh9lz9U+l/epdxqpl/uITloFIAecvJ6wRo4xtmuGlCkj/ian
7Lh6t0EPO/gGUWCWCe37s5gddia7kC/uQP/ZgNpXT+hJAsqRa4FIueaSV/fUhMO0
veSiDFxh9avQOM2//xUU2tHp8HRLj6knVXbQC/Cd3zUDEsqgGj45AqnrkPLi8wMH
v4fk9z8e2wfGSWLcNoUdISF6LLG7wZA19Myaxrewepm3YxI3T7e8wO75MlN3EHXI
lyo6s9+y5eNfHSXSWC56cJuHKegIDzmEANMu1n7MjdXB22I6toBPPY+CwvP+lbSh
bh4zW/wbwI5xzjL0X/dKnswLEYShFSmbcyrSb6nI6/YxgZ91urf8bzZQKA6W5w93
l8yJcJb+vPA6de+uBXDLDsX5oETtvdVCV9jqqUt007vrtsFJEAqWiH2EV8xfTPzq
yy7Go0POAtT+10PPRl8C4z9hEnIjnEpn4JI5olutK9nMGawVbY4SOi4BCY4y/ejH
D7lyGzI7OKXgGRQJZ0SCTPv64TG307lC1M6SdKK0OpzzQb4btDW/d3hUy7S++0Lt
`protect END_PROTECTED
