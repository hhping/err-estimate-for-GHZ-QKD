`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TXoKDyf1+d0ZdDyDQIQYAVD2UjnNmh0SCgos5COHQyMuirr9HWMZ3Uzydhvk9Y4N
gslpg05Zu4LQaXCrhx9XljBjffhVoK9uk16vjF5QZC8T+VBnvAO5onfGYSFn9JqQ
FcjRZdlLWufxUpYLvypFTTap+N35UiutiZjiHnnYj3/TunTXLWX36JP5xetjDJK7
62QzE/YK4ou2e0+FBOVVpHWzgCbcO+AEggdgHH+GiJrR/exSb3DWbSlRDrg/AydO
w51ulQhNo90bD6fh3L3o1yFoSTlJxrdRWynACfwRK9bmqnLA5XF4V/8j81NOwxfZ
UoMSNCyQ6vBYX2wjtwFfFHtC+UkAvWK3JA8IWV15DRc6Jlm69c22dM0DbmOYGK+6
EBt6yme2+9vL0ZP+fxDi1xvv6BSOXjzdqfSnzGpuLNXe7p0VTPnrocHhtyLxW7aP
h99DAHofvJEYPx5qJ7+g+xE8AjqsL0g/Ih8bI+iebKTpREJcDDRhI0h1FVJl92nu
pi9Z70jcHKDSG126+YW60RTioqznuJtn/etZGQ1rvTqX8+EkW/FKBKb6om/naO8W
vlAIv/Tb0QborRV77ZMq5o7EiWkWJYR06SB+7zzFSe8x4lXX1CNIta3gcegpWXnt
6Kp6t+owei9ZKSwk55ViKvD97Ib3E/NoL4lVALct9NhwmCpDPcF2m2d6O5JNbrFT
9H5b1cRpx7JY6PJ2Q5cW4QtsFaRSn9Mgz+1tyPOStdlh0EHU/t2RXV7yA0bkuIm7
NZnEEGXH0dWvtoJy4/AQ9du9k1yEUTlzTCN952Fi70s=
`protect END_PROTECTED
