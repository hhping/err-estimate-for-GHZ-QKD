`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qm0R6ZY6wNGXWWJDM51McD1YJyEbUdPAeIik7zIRFHtp1d7RiFjos485wbXHHu/K
RCyraMKZkqaV1ElrE5D1o6UvWO6K2R10twuzZjAbjFt9R2Vfwz+GeIn51gEcPiyq
6ptvmjqeTr3zgkc1WsWnHncJxlmGfGwSsactpEQv+fTN4S74OjBv27zR3WwaDfZz
xJTN67nx7hBG8WMSxdvOmBovnPetdLlyx5QtQmvZGel9HuL0i9W+9PVhuKQee0hz
e8tHfC+Zphoqmhcs8+v4unhJxf1OVRKLjel2xj+G5SHhhum11gQZ9AvmRUAMnGeD
WRuEcPRaYSl1eDUnIRfT4JQDFPx6cvV2/C02xNIAECtiKsHOkmuCEz+d06oNRO5a
7cRIx/IarDiBngXmOuDr0z2MUwJp2NkgxxJIZ21btEhLEGt78eSwLBgxhhY5z6zB
TUAc4/j+q6A+3oSYadvtQtJX6UPhzQ4GKbC9fIIoHCL9ponm8VmZGNKztY2xZYVI
ZxrCcxN7vrQtTjJFnssT7Zzj2gAIWchLVkZuuSdMSczXzuFR7TyLealcY+i70Rgh
pO78nz4EyeSmyK1h4DNU/VZstvjaDTkMjWafKTB96J9l5Pj+BrXRzLkysT04WNMa
jLa4GAh4gQ7Q3JLMDWGpfzon+oGoD69Sodf5n5pXd8NS/uJvR8qwps2bGWqOYhQj
OtaDbMWP/xPj+1la5AuOGr4+1AJw5ymVDKCtoOkMyAVoTW8u3wOxrhFzaKCyb4NS
rZ1/cwrN8AnMs3TCFMoJJQE2ztI11Eimf2vEvtZB1SNyWbZorXz4V31OaqtDK1Y5
biCvCTTKd2LAdkMfVfQ8Lo5sFJDArylc8u43Q5K1ZefITeWdgLU37Kkca55PuLXG
JaHm867NJhYqYbsifmZApUT69jjC4MmPXyXycpbe7dHEOF4wZgt5Fkq/S9bH769I
nt7wfFH/+c2ohJ7ws3kAI5JejTQBtebJVE7Ar3Kh4u+9Mut/4fh4f6Yz5fpEPvUD
cNpsBEplDwDR8l9HqrsWzXTlFcIwhx2zWDhPp3wySn92TKvYew1ryvmCQolWwl0f
H7nJNcvQjvxCiF9qajYa4MoQmP6eEyhs11FljcTSV3+XCToGnyChewYd1hdcbNG2
CKeEfF/n0HgDyhp7iPw+IpyofWo4LP/iQPNcPJ9FbHuk7sBMB6plFlTNo2bi92/Y
cFCSYFFA9uUH26CS8sfNUegIqWaOBfXTVL/minfTdJuJ+b3zm5wRlvuIsnCzCRhn
Xc1WPIX/3m/XB7bi7y2ma5PVlcoMLMMvg8y1WQxARVgtyTGEOkIxXbi7rk3fGza9
ItmQSUoezneJVi0p4GQCT7cWbgyp3y0p3V5xgd3384JOT3FKTif75IoTmzMw0pHN
o7GmEM5nI3LFFM30FsjAR/SkVqKqtjDBGDeSwRV5CsFZyj7x/HAbVRhBkhQriMKm
MKmFISNdVvscxwZWMK9Ywfvb2sv7ah2D6ZUsEANx8bGyllHEaCw0xrRMoNFD9Wwm
M/ByHUEcPJznKU+msE6WDmju1yQ7T2nA1D5jKFlIElakiGjmq9sZPaP5ibSZlehi
fGk5ZyoHqK5MDTYl1HFrpM7s3Yzngc6hLu/4mbpw/S2tvxyg6Gy5OikxpRV/rlmN
IzvBLsKzWvPIsRH58imgG6CdU5p1MaLa3/rwxw3LbN1vUIvSylf6bRocDVE3tkpk
MZ8Rv5vMFSumuh6bR9ID+lJJZdMpNr8ZpWlJjwxbYKRqPzptCYzdqPlqUlYDwKFj
SGwcQRxRKyDLEy2PS5LH+UShg3eBwDy7Zs8VRULZ+CaB03yBFAirgcwn4wsIz0e8
FinAe1fh1/YkfQYL9RO+UWlhCpap6MuEJQlx939/MPHOL4ya7JLEx3oHnGw3V7bC
VHbr0GfFHwSiNLsaaQ1jtS1qdjvDHHD/qugMNL8gJGuPYTIBdY8usFz58We5Ga7n
CD7N6LjIG6SXa6++OFZRhXzGuyHYoMBurZgN5YlOByBu3krUXFA4HTY7KcIveP13
enYwkLUbd/MsrOiTqcnNom0bV33heRsntIzQQn1XUpi3jEhsigWtywNv8XxcuOBN
33yJ+P3cJEqqg0por8CwXQssCWXZTioBQ7w8aZUM/N4msFsxO8fcMVsE5b4dEDCF
11BxNulNiOlXVjKvOaFUsBc286b49pLSTnmyCc3gIPIi12m+75qBVCtcB77VhkFa
0fi+p+WpWAvfs42WiR7nK/XLkFdMvTxII9bU3dKbkWo2zn/defvW9QUzmAYjiHQl
rK4uAj2lGRZ/QayEqwYLn61IA63A3YPo52qvauZ/jMWGvFKa4zbX55PRkIHwBSly
vv3sG5R4W2+LnRtiKeJoPAAKPeqj2bPDmnx9wTV2dlhREeu9dlerAzXIFFBoRoaK
1lsilrNaF7fppogv9ML2XK01CEf9mpRjDK1AlvMqVrfaTQ8Lnf9ZeuMPkbUCZC4l
HvJQMix2M6+Tce2IBPqNcNIAyTtwu6Wgj/mA/y6LoNFDBQrBUXVxDkFuEoJrHzjf
VkyADlNWsll6XDb6xO05bwWjfhYX64NhqFQ4f+ZtlvHShBqYmN57Nkoa7ur7vBbO
+K+pg5maYWmNHaYztVGiOqGnIb25Bw23N0ZoEn0E5AY1bdxzKqLSX0aobE/hOBfo
OBYTefICkLhJCPTDtBoW6DItySnryTNSJDVL1qwUf5Tzn5OZSzdQomyhL+w9wowz
gGTRIHTHMSUJuuV92okcrd9bBsGTB8OXGZrlcBJTbXvbjA/GCLmzfOh3ZRYlSDi8
M+Hbdk6ikYgpAojD9mxzbtXf6vfRfwRDMM8jAVHlmotn1vaNX6jjkOq/fOldj5us
BlYq9kd8uv2gJljwKG2m0o/eyWzBdUOVkSZYXl6s2Zp8IYd6L+QhS7bQG0b1hZ/J
GezmC4W5l4KBWDaN4hhJabC/w++fPSBRmXtdwm0gsJE5JRENKjE5qTh5x/mb6hu5
eneYldnTYq9EVHuZMGi2PlQwiTILv5GJMScseSuJh7uLnd8ft1vBMsJc4Czl1xIc
uxdtWfQOtPPZk5eQLxOVdOGUqFX+mwk54l0l1pDE9c8QFEBVeSUXn9X/h9JdK0Za
uAQx8UYHsDE9xO6jmQQOPLqCFx03dyCboAYm5OAcAW1d2HPEJnTj4MVd7Pznq5Bm
Fu59GiMmFtpAVLouo7VzMIt3Y3pIw8Y0wNugPwK2J9BmOOJRepxAdyXuZe72lG6i
jRkJzaMLhiv1ISg8E+veVdRm++eKK+AyaE0qcVsEdlF4nnWl81G/d/hh4fT+w73Q
L6zYFLCQPWT0Mn0XIQDXPtxcPhvd3OEJlz2/gH1lfD/jSylWryWqRPey1frPe1H2
39kEBOK1tnqAt4MNrDZG+rS/Q3itX3sFt8WXyDDqS4scbM0Og2jGDDcjrFlpNoNG
1dEW4R8xHXq0HnvOHn8FBkgbRqWCSLQE0ESwqNHFSE/0a/VymfXUwri3GQtxk7DJ
cdwnxq93MFweBDN0yoh/T6Ct0iPsS92Sjph49NZvsMWRZD8/3wBwvEIXRjKc9jm4
NYjn+FYwYA0xuOQvLrCwXPqOjeulgkEF79wIEZ0HfWrKlxXJSJUmuSs6WiRD8ZoS
vnqKjgB2l2ZG8rZPhLv7lSQEIlQXIrKvPb/lfYyRdIygT8Q4qwuiRZUpYkHM3ePT
lS3AewFpZBz6UEDyCm06ygfObmYmhwWJfzA8DzA1/nSNnIwIBt9DzbSbsK7GuyXP
4wceFkB4MxwmsmkkkkwqXYUbelGJ1QAJzTcTu34Wlu3Dnof8baNUaOHQ4gNrBxTQ
D9BDthB63IbWbldrxI6aUbboIc6zQbTmnCiRMGWab2Mls2IXK0kPfeWuoLsmy3UK
/vtGjCJvTgnUuB7YeI28uGPb/H+CIg6ykGV6n4sZpWiicQ88Yfu8xH0sigp4Tapm
ETagAlBcuwhjlrRG/L2gX8vQV5m8vdf3wJjLzc+JtJWrGSVIuzA0S/b5y8dUSlrH
/D2M3LWlFqZ6DpAb66KYlyx/5+SRhc6nudTzh+OE+inzlv0GpFHAlTblW9CF4gGk
WZtL1La/ZTnK2LQOoFeShE1pRhJ96DyGHhAIf8Q5WLdydD/+TOtLO0zSXhd4fQFs
1hcOwpUHKk3raspofs9UPm+lCLRz61Qda9F5pdGMCm/IAQuQBkxPq12d4vqLIHoB
gg9650VO6H8GogBK6r//78hd7ytvwZurmmziBLZ1EasKTwqKYac9t7mreOOHU/iP
IjkYF/QvFURltHaWk+aknAs6GQBSfgqBXe0g5CZTAaf8XJFGYWPqUnC+HL4tFF9M
sMJyiQAVZA8K5UQnF1pcwmGcMnxDF9E8iwW1C+clOkloPaS4QvffmvJk62x4ob5e
PsEIirLxyn42rim3rw4D/XXKxd00KM1GjRVjthpuDTmH3QASD1cZQf/HJeVE5RMt
63NlZc8UNhPtpk6+m9WEdDd/ekHCNyXIo4sww8lc5xuoX6gS9XhigQO4mwb9dv9G
oge3RDqlpi6Cekx1xU3KBxVs1rWAnp4mXieOqvTDLvIkyxtI84D0+q7t8yUKEVee
+7seieHSrdT5g6UgbzFiyKIHR6v5nWupqZ2q0Quczq4m3tukKDRyyQCgMEFweP5o
vFg/Scs3cODM79BjA/EgM+FsCvm6IqizTTFv1POvWG9iACir80t46NebNb+AyNP4
mjduT+GSGt5WJHie0He8J5yB+nO2JtDKODJp/dEbAbIqPksLmxuYJERImU9MdRJ7
Zqc7SHN/GxpCouXAq3+Z57e0sKGcg1iI+hFdr3dJfCiZq1qvMdKNm6GthGZdoxiZ
+kUqZfvGxoAIbF5qf+mo+JSq/k1nJsfpZ7x2vOqsAQR2rbLk5AnzLetHEEAB00Pk
7PP92rnTJ6hXiO901kIrTYlcUmriU5G0ZIGXQN8dkDeinJ+pJQXo5WB1KB4OLAyb
6LLYDC12GN8NeGeoxVYPj03Pf4NGFFDiwysfRGTHjResr8FeobccA3fpocahysLH
8fnA10h+kHd+y3Sbdf5J0c+k6QPr0E3S86qMmAlBFdKl2Tg4DgcZ0bdfW9P120Qe
vdDzefgCLMhOBxtTwg1PkVJ/6QrjIvrh6cM8M8oWx1JlTlliwwI3grf84BLR5V+e
CLMkYpRTc0CkyedPMtvvnEMUjiieUBZMbnCXOatIqjfpeuPn2bDk+dtmM/VMbtIG
OoJuMcTB+OuzIEp5L4MqVQGcGGKZ2QPoQa31f7aaPlguaZg5k8HxpPAI4CKYkFb2
qXOYF1zIoKzn2w2DboCwVKG0BhwmlVokbX/4gHTWXXBMQlXZGYiOiVXO8aZDr3Nr
gvaN4fGftY+QM7Apal0HfE5ZdiTVofQckuelgLNK3nC0YbSc9B624Z2/DMiOgjqK
rikrvH2sM0UUpDSZoC67oe8qAd8gjh2bQV2Zjz1ZNKkE0BZSh5fxxDTRN6Rrl0lw
OjTiZy0hdLrmNVqUKIciZZxN2IvWG8SkUQ9ytzZM3jEO/rJys5OvKS8CBrFl36qa
nFs+skD4IlmOTB2FDYps66tfWYxCRRo3UabFwarKDRrzvB8iHxlDpSSd9tDt5ZQY
+pMOk5v+1vqGKCswFJwLLZt8m0uQug9l4mBjT3cWf8ucWkRjU7Hgh6sIhS2aVhkE
UnSahnzVemSdFg/5jq5whTrTe2BeC0JGpmli6rl7u7rIrEfC+HxeTqGiy+cWQNTA
OAabjYz1nIAs34ZSY1w9rmmpGLCiDxejudVCwN8smYxJThg5entmustPWx45VqKw
zEItIT4GB6IBinh1ujMkoX7aLFA9cHlgUnjbdmgjeid7L6bWW6JpKb0pPI0cLhn/
rUtr5pT0GAIA8lUoOl9ENqTagnHhj9SuxBNQsPMYeKHGS68PxlaLTMwp89AClQnA
7wjaPHFBrGcBaBoUffEgrRrlNmHparoJ0gA8OwRoUxcoaTLzK2pISceEUQgFz14R
PrBufeeeAoK6CWflebRLi6HaVhr1xc43eCzMPi6Db1vAOyB26qCSXRRj+KDhOqNk
unsJZ+X2hqrrVhNEFQ4xV4ns3rXqSWqv3qMaGRdmIiNKLIiI9G9AtKh7UfdT0/EI
2+nA91VueAoBqZvmUXIONclcMxBt7nxtmJKEwlOt5TLY9jy/LTvvSoBHu0vNaTaF
BtBDttNk/JXkf1cdgBcqAAoDjULOApZ08/qYFr217ijejR1+KjmozMHgY0D9tpj4
t4ltbgow823fjWn+S9faH7Jq2bQ0DZIMKaXlTOr0YJ5LpGIH0h02kJ83K1G+MrP+
9Jr6g0w0xqAnlbUPdrSKPyYKdbTnqR7o33RCyUjzA2AXbAa3V/XxcQ1kcmWni4rm
cfZdefI1b6jiBQw6MDaNK9nVjBGXbUPDve0oeac09monZCaVacWXJUuW/N7FLSaI
hL+21YnL4C8RifXgED70QDfZGvoA8add2uYtKwmSZ1wiNfrF2eHxChV6ZtHCXBFr
7Cc4v9EpNQxDUmUQBPK2ZIvTXxmHjnpFmT0tXYqTHhLnx/kptF6R7LvWMub4vX0O
Rf/IFdSC//M02fDqL8uBFaALjCYReDJ/0vHLMYX7WsJNNzbDjpJ+vEKeufu9sAJr
ZCWydnZsukrEo+VSKp/lH/Rh/e4WyYYxdGKNSPmm1FRglIqkO7VACTitnS/kep1U
CBIj3eRFsIvx/i3tiZRnsHNrqWJIWg8cP/10g23BNB6k2hOVkdBll88M0mugkLmp
yjK432Spd8QTmqyjQT6w/qbNY0yVB47/0weZBIwNqQrZ2rRTK/JjALBTtEzu1Qn4
DXwUm1iX8oVh+eJ8iHoCxur4LO+u+YGr5hUhHLU3JUVnSfnUwpulVZiQVxIo6I4Y
Q91Rw3KQ+bMRwyyFzxPPqi9GZSFNt+BgZiNmE954BrNxlhVatHARaAElkd8TtyDy
RivIhxz73jYK2xkdJwkZrV4VQq0FIIYAXaW9TIDEnsw/s2xtrl3X0axzrKQrcYIP
mqYomWo9a42oF4ntT3pNQctayfX6YoAEZicw/pEb1USKoKvqn+txkPvY8Azgr9ch
InTOSS99xt345clvNXVBKktcyWnpf5bBxRb9A9gortAIaGzK4AkhJlpUYRSbuRaB
9h3oZ+eQcRi21e83J0KBwNJqill2+Six6kso2P7NkByhJto5AVfjdG2vCwC4bAIh
1o8MSxPu1S1wa4ObbIprZC0Ozocf+rGsDxefL3fUjPFB3IhonJjXmPrev2Leumxk
kYjiZbanK6HjbRd9uN7Ufn0o8l5ktYd8ibUVIxVy+v5zGbq21WLCv21Pid70bnJM
qaPABYx85uZebHOg33iWiL8Q5BAmIONeAqNO2j1aLeJhOcoIGCROB9hSGpo7zhwt
awj0TsFRZCLqlP0h/Z2RGDkiCFmoynbaZSHukl8dn9EDLICIUtdS1ofc4SeJnXWJ
zrHg7edkPwzMAtRxo3M09oCg2Jl4xhaomRjhy3dQJG76ay262i9XsusCe2weE0Da
YvHGsLVktWbl2XHDZPlR/tSiap3OgAG0DThO9fyBm3eETs8HPyhI+U6TnGgphbLb
thuN1yWFMAqLPspiIa2Xm4sJs9YkwIJsfvUd5Zkh7v1/+gauRkRpOORkIHdcp6H4
gmjwUq/VrcgkF4RYTGfmveM9uC4whu/GL8XCcgvqqw+vOx+SIZZzjtAbXgUJ7chh
X9pBh2P/8YeFHhw1ED85eOzha8GhAZm1pNhcNsO9fvAEMOWym635HHvQ/qXsEFQP
9W+WP/Ri+334gEyV/hoWwxwUHpk7Oi/nppnLWqjUtu0Nzuq9WRq8FQC1s8uf/tY2
KVn8CEmz5y4IDtXagE4MSX5buoFJayKIbwk5eHEpbM37/IcnHepZdb8LUGUStZOB
Khn5Aa/tcv6kijW9sG81EUN2XS9YCcqVXVrggnKrecbd9u+ZMu6b06g2FhSTQwUz
zBbhzWycDa+WMFBBox5ON9g6l3yhLThm7j83TFMfsIxjvGHQj0wdQ7Fgb+pa5XgW
k5ksb7RsQBiMm3+jrPCojSQ2CwFJZM0HPM0/GJS/oUHvgOjz1VxbBHjD04phjlz5
8TULO0CTnk9dam7Fc78SK8FFCyKpbFN+bEyLX9ezpk/gxdKVYzwRUvYlKc3g2P35
OeJ7VnHv8/7KO3Kgcc7sx98ZluSxSlAkiZ3pKnSOWEeqGzHVpSBjr+fl7T2XhG91
GuLfvDZ+Qd/eNm68K3zRJNSx6jkvurJMjXed+Z6TixF3wpLjAa3CKsBljkmj3g65
IpI99TknJsnfv0S39VPqUHw8+qWVFNrVMqoZMpJxZQs+ux2Q5rfSIpyvemfhV+dF
QJUIp+K/qVe8LI6AdNNqsSoXdM10k+Vwbu0TgubhzfDpXv0VYpnEE4llN3oOkxwE
tzst2mXPE/nN7Kfho7Uteiw3SNcOxHlz2wvHeR//L5T5e4bm1dXE7MH/9DtHxww2
Hr6NxZlprXrzjxzxaSvHXtC7DGjaLgNEjERPYxpp3FWbqKNRYkpMFOYqZBvDeYdm
NvX3rdEBcQoyr+tYb52YZ0cJql4bx5PSO5/qE5hM4J+xCr0ffl6qOpu//CWl0OW1
5dVFocIHDt+bDHpFR8gFUhYJ+FKNJSvSzqhFQ8zo848GwfhdVUqCpxU4RgOf2uqN
X8FsGHsgmgC9NdzA9Z1YHvF/haarAxmW6i4zO7JEYXuf9/5AFQI/mMsNM9URL5Dd
WDLjKi/3rGvOba411WHsXzQ3ot3KAEzeURCNKrUPZ5u2ZdXgYBGv2oaPNrPXlNCD
1vcPMcXW0YJNExaZBY7mFKMyg02sqSBcyTNmXzBrPpfVFqbgv5iP0K/58wM65iKM
Z1lLr3bpqGAfFOJytnVg8JeA/OeRv4g38aTtiQSmli7bRGU6sPSlHC0KXzbYMNp5
AH672t1COCesznJI92aXM4Kswjhj3IkXd4eow4QhWaHhSZCx97YqsECEPGfnrNnl
Ew3cblp7MpHt4KdFrnYDbTNwfZ9upcrOyXQqaREsHsn7Zch1j/vlwcFkJ1Tb9sP+
rYeRno52SKSSTWz5pdGc3BlZZUfEpBUvv3o0g31Y1wIA2QaXDVfQtVd55qbG9Vk7
lJns//JEBYnMldEe9I0zYr9e3iin5+/KQY4ON5lPQvXdy/+RWG1LVnsIDuh6Cbr2
vh65kZtNyCMAbE6h5AP0/pmXR0PZEjZo/CnTTOihkcpAEsOFH7P4GyOL4Vjjnvdt
JsPZbAVcHHPZo2e8pCFpQ774rP6j54zzHEaihtdQKJybyH5VPuevd8D1WAjnPMq4
uLCGWFR1ffPc5yQ6wMsN9k91SgClA2XMgxF/ApDD0D8ToppmKdUI1t/as1TYQV9T
3albx3N0NngDvqQnG6I4goVc/c5iFBEwUPxzcMto2Ev5qxpZmJFg/PVSGWOCeClS
KlFnjHxOCPMZB/tVsuG2Cke1dLmz0uaZ/DWLNvMa0Mhp6+WZ7aEjmPDV6glDnEht
NiHC/CM/MswZ1jyuvV+n9GatKMG9tqzPTRHInzRIBdFWh8TwCPcmoaeWek67/UnR
rIj3kWOiSoAshIKpxFIgRMtJm7heSd2PpK5hhzFVuz8ZSrMIT+zbp9nBrYJONl6S
Olf+ig41HWGEfPBD3lJvO0mYOBK/7ss1bvjXv5iKpvNxBJl8VyjBtaQH35ywqelG
ZhLhPyML3q2X7MHcuQkv2wdnliwGVUYB94QXY5knwMGiiEYUu5uuwPSYlg8Uvcwx
b+vuK0Zbv5IWiObcFZQzjxXDe5YBQW6jHh2CAUWA3cdulv6CLUJCYKc8Lt1PGuBk
PsVBB6Q1TOMuetGQr4ohKpKr7TeoO+cYvEbHuq3C+sRwWthbWYe8eceNK7xOt6CN
DNttx+cVMnnGa08s4Q+20M/EoXh4ZOvPK4t3c0PL3rscfC6sXxK8/GL53gRaCMIX
14x3UALYopMNFeKGmECC72jr0uPOx2VRASFp5olpj34glpxSmKUghKFWbzUoNQaL
XN3HURIYwrhbJKAPSZYC4rHLZjxJMDVKcxj9sNYfCgNLoqBMPQn4MAb5aQcQVf8M
g2QYAKURRyQAexlAOnrhXsTEOiWa8Ots4fMlNzUyntaGrf51gbyBCI12fZ9Cxwss
RxVxXptVJZssqxSucMuyVcIF67UsCub8L7G2Q0gL1eXYw5ssHu0dltARSOUVdqi+
/UJLU4z2/50uNxxp3DYl4nej6sUASGlNHWh4Umjy98MK4sjY6KUl7oKZ+FRnmfE8
8semF8nYP06QHwbiIWSlg5YgrPmw0asToxYXHLhY3+COGRiZl5S3SzXfp8I9c/DX
0o+0dUtkHhkeHmqzl+4Oy+iuiecsVK1Qf/IqOm5uo//3ElGYXlEojSiTl5yBlpr6
ke2a32Zb/qL+qm/C7sRxJPCcPpCOy9dOjVvx9re68Nnp3sjkAGsbdtejSul0a4dB
iJexxCaYAR8tfgzx7KGX+ER7sbWL8CbWOWQHkbB49mXwEIIfhpD3q4Vgw+fNuaJu
wZace/TCUjs7IYT3RPVk5xdTmnwf8vyKxM8tCmjc6QoIixoIhL/9S2EhDuPstEmx
GtK/oU13OMEm1VaZ8k9GhJJmmXtuLFo7za9KD6CDBNFbAWjGay9pQgkEtup5587Q
DqIliolKu8FgjoqCjsbDsCqfsipBF/kwySgDFb57zMIb3iiGBzLM6KyusQ+gsWdy
2sFY+jMkjoACqYjSeGNsp1re4XBl8vBZ0kkvt73Ql7MvTJGl/LMJIluWjImd1KE8
5KOJhN8hK174YFHjAGkoxBmI04WQEMVBahEhj7X8Ngc8b9TOSrrhqetLaYxDa608
gg76VY55rpMAPrSBnwa0SgHMeQCx8fuz7CfgJSYd5lnTQR6Dr2rgFLXaxBdOjXJ8
IfjwIMPjaKvw3uAd0pByv7I0AYIhna7vPkIbYPAKQ7nMsR+GfJih4KfTbgACy9Ik
QLXsqxPvpuJ/oSAFJV54D721ugY9EYSdW71YKP+Ou6V/qyWlm3aJQSt35PRhux5C
SR2ZMg+QGh3UZm340HMSGoCZBYaxH86QPwn8U7OAwAg4aUpdXbvSSkKCv957n5vY
p2cB4fK3VPkODo0HpFOEm8aq21N7j+hRTDjvk+jvVctmXQoDK1r8QxCQs1wpEx0E
+BFk8utDSzxviOVreYXiZJssQphrEDOJHWTL1/XJLaQ9iORSu4JFoT31avuVM+0z
rt3E0v/tHDm4/z1ncjD9Alq1zBbb8WA210uko199XVZo++bNiGPQPHLCVcSLKIIU
kSZ4zMc6RMNXVDtw/HJGyYJPjNLuPn/vPnr76W4uhqyo0Wzx+wbpw53iPsDw6zF4
fX4ZXZ4mn7Os8bLmuJftbyua1Lhek3p7YX2PN0YxwZ3eQ6ThGzmyCn6SH5MRR5rB
rdJH/PIp4lYQUsoiD6DYnyNwAo7xjOwQ5iOCsAo8fjbMzSvECzMhc65UeV9q+YSZ
iH9lh62wRcwFaxrp9041JrAJl87dcjXmBD6+FgwO7L00MvljbyYESurw6/BW0ujM
/yO59UNiLTeZb83zIBG2NYCZ0XMkWt1/eYZS3DkzT48Dwz5/jda3qp4ZVWeNlFUi
KInEyuR2WOs9JhVCEVLWMwavEBrt5Fi31rbRyZSBgrwYGMAwJdLZVmO3jyg/rtS6
sJsriLjwEdoa6b9vujeZhcr2nItk3kHo3CFVoCtcy4cm7yM+egbr2VzTfiQwOWFv
Ki50SmW8UcISRQaYPaN1xb1xhG+cAY79gjxyVE2G0Itn8A1HXK2J8XuMpeXCIo7D
tGuianzF6jwhiL0I24eAtVlRHe71m3S0b2Z3JrZ2nBIGQqTTLJS65ZT17glkx3Xk
YmVvEZxNTD7naj/kxvfrBx+amoo3k9Mi2aNz2dCAZbE9GaKG5y9o+med3of5npPc
LXRKqPozPaC2rxjxHak/ZEX8Etp4b7vsgiqHXxCnuUcge3l+hUQNAVCNRCYiHtIA
Cp/hnBYDipQTJDiwDU0LGsGLXA5qlpMWY4M2dbLOvPUUThwH1c9JUrHlP6JO/pVL
VqCz4NTguT02hd3wW1uZOuGbm2RKE73wspQ+/NmYFB8wRCjiz10TVuw3DoNgDVzx
a6TEjZno/OvUWf9CoPP666Tmh1RuCMlQZeLLzBFhduX7o+ODB/ZEtJ3kw+tNejA2
waZDIw7uw5C91GBwgXsYlN6T1ktQQgtEA5K6Hcw04jQoaUzIijf0Jr11HnumUOZf
luQdE2qO8eT3netNCa/y6E5JBdlMoFQ0+MzeNZrs+8UA4AbvDouW4ieDt68DgHii
5iDBrz88dTt0EDp+GGvYluZLDb3HiyNs+Mj2Lj1OELuliM9aZGIgRqK8f4Kdw/FB
BC8OC/mdrCzcAroF8yvwWy8fNsyYWlGJGzWFWBqoJwxbpAfT7i2kWVWru83fuDK2
brVLkWFTL4gL8pLLZ2Kh8bd/J2Q6U1E/pbMo+4J+2H0fppnfDwKDpAK3bMu+jvSa
usfMS/C4MOCMZcwapsZGbQA6WzLthhriKrjbSXB5gpGM6Ao7kKSNm6i796XIIHZ7
kzDqCqnqTJ5UWKRWRZ7DtxceNAY4mAhbxfYxdXqIyMO/3R47AbPmR0dKV3xXMMvf
zpdAB9uxQoxHQ/1egCNdih+5FJ2/nK6bL+QyPnOvAeybPJgAY7kCnRRt9CucnVlt
NujiZrD/8MynKhHb2DkWZrEryURW8rx/yfeGbcdBxGEmHWvBsHaIJlSsr3s4MdSS
xlrBKbgt9aw7xxFwsWSuyAGHwoHNbZGHZ5pqRmqDxjFEf3FyP5d8QRmuKKmUt9pm
GlNDxhdF4IKN2Bq1fihn0RNPRyNmip6DoQyDDgKvhuDrvjacvu97hkqGfsIipip2
WxiHUotcL9Zs3BGnNVPkveZ+KQESOu1fmoqvtvL7zW9ClKLbufmmPEgPcvVahekz
jer3BYU882gvyAUgu/y9kathQcPVJdv0Cu9VCAMR056G1oxONlv45kmn1bIMuXBP
ZIwKJv9bpXkf48YSa3RAfVxME8SaMsBr1E4teS5Pjx2ZNeKBKa+auKw6zlp1/BWq
ayx4ovuExhyuSr8vV7jQElea/n9HyNO3mjulm5JsrWhM7q5dErNFonsDmuBBXnjE
O2Cm9jrMhOARFLppqjjbjRgWiDYb/wE2XakE5aTUJayIdXDMqxQOx9nsWgua6Tcv
Jd0xpwyCA7wgJRHD2GvDh62AZQyak9I2Axgxu11XLtdShpp3nN0wXG+po7JZ/g18
kP1VaU90ZnQfUGidRvFaPupkZmcOW3xy5qDvm8OOBb8+GngGP61cy3d1oX+LzaaT
wGVpWQJWwWM4pzSVzi5HUSI94gRY+aUoWwITZ6/SaHojOpezQXadqPm8NFf0pRpH
2IiqgIu1DhESTXPyyrPIg5Fp+se+F3azMSz2NWWm1hnOHOtRdumIUzjq68VBssBz
I0ETMmzqwPLuyy18j45oRIpq/ZUJwLErHTkGrVRkCbpfBCr3tzTs72DoGCSG4Dag
OmBNv/YqsuzAfGAluNP1xVja3AigPCFkFOKgyBVMawD2jI/kffbFc5AOpPeYOPIw
txjb6q3OvxEqKXlYBdkooYx7jH9AQo3oPkQT7ZghAUcoH0mbDiR6O9Z53k4mbxus
5c3D0ksQF/hYueuSzwreU4Qbz4IhjmC2t848UusxGpTwCHO4ui+q40Dwi3q14ELY
jwHdZPYqjr4+aaFsN0M9XMqzg/r6TgG5viZyG6xsL5ceyRICpsiaJ0MUYLx8e8MF
O0C0DwHz3N8WTTwWTOC5R674VOiP9yuIAWdrZYodrvg085JvGqj169PJyFgfNC8m
nPxVMOP4tYT6G/YprxjwKh74H+iN3o1f3lv34Ju6A7cz9pppGUl51OHAkjdYvNaG
fHDP61LSr76ol258m8lSWQE2uRoMUMft8aZtQ8mhjy/n7moLgl/szpXzwuV5NCRJ
p9pWau8Gu+tucEK4JxRvfIGKRYjJjEqWRO55we6QVxOO8vOdCTNFxqWV5bXstqd/
rHQqfhnvZggTBVKNCIfwERiRTyyJkKR3dokjW7GKetw14UpH/4y4dbO5gEWbLCes
FYCDSB4ixNu8SFj9E3FpXXdRf2wi5ONQZsGj5BcytQH8CceiB/WsqMPulJHIl5Rd
5N37LTbZJvaOaz83CLYwqOsTXX4Ww4etunq089rl7xzp9YhnMOrkR+MXR+CMSLr7
5QT4HFO9o/6kSWJ8//M/gk+Gx6QSPC0rLi0SIhMz2J91SSv4GOioUKshoq9KOX40
mgttjyfDWSdePEwnJSSdTw637Nrw7Om9RIp8YYRkWs8FAWMT/ebIwT+mRYS5eilB
jWGtspZQQ3uZfghUuCczTMjDFwTjGbmElF8Xf9tmnyLi8Vp0YlLeeYkHr9wA641R
qCvkD14eFryPNBO++u/gJxRpCixeNGoAAwoJVS+RlgCCsB87aobqVVe0CU1V6W6k
Z6h45si9loDSsIEt1FZ2SlXBih9ftfvjYr09IPjvIsIbfoV7sv4u1c8LkG3SyFVm
w5yWNSvGX63dvdScts3eJhepjra6kXpRmKbE+opLiI+BbOFpxl650Z5N8OFKX726
vN6dpfcLWuh9svmaKBTIiQOHrgXy+DEfHpQXhGsNw2YrxqBLQdHLo5aXZVF0AM55
D1xcsn3RuKa8/oGCwWBb3budpD43i5/DtRPuHSsM2G5y66w/2MU/cNBVDuY1+3YT
2Z784rc7Cec6O4X6RPlTcw==
`protect END_PROTECTED
