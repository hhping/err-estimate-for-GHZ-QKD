`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
koGLRRIQezYerXUfIcgzoJcB/K1tE/DvTgYJ/KBVDyLEPRq8vm9HyWwMDNTH9NSW
gNqf2uiIpvXZ8mo5d0A01K9Jft8XEriSfYJBDMh95KD8CbzxlYKbReLEVJ0ZMtj2
2SAdWPLc97P2CXVnxens+r+PpG5w2qkeIVbrDuVgUHZ+VKnzasihnmxlYGTNUy8x
IGiY0+J8YvrbTz3yIuk3TPRDMLHqv3Kj+wAUFNf5FK+aUks3jQcL9CJNDcgyI/GQ
Qa6aSTv0CUmHK1kMzEY/s+GLqq7SvdsNWA9GLNsHxINzE6DgGfoKJ7dml6z1+Smj
asNdyWvLAGGlcT7aXwH6Soe7pwqyjuCvq3DKTT8GrgDP0B5oLjivGu5tyMQsv8I4
eN6gekp8idegV2B30CY7gf0FIruSZulIol0G1R0pge9BUJsPJU3ErQWQ7Z8239+6
KsU3TjBBG99N+Ye1nMCgYayaiVR78pA3Lx0IINeixF7RrvRl5uXq+oQSaIPJqjZ8
eSTheFz3kCNE60WyIPkvVwVlr2gPKfS5P9DfRIaFs+2MlL12ozczFJRXxQdCdYBv
`protect END_PROTECTED
