`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nHJfKoAgovYfsSzI1i70POhHjYycoDM+QkCpmt8Kb0Iqj8cSqPG/mj2vNGtPNTzA
Tv1LH2fYXm1mSxe+SZ19+wRBbldQgUrHR9aSFW62UyAqaSdqEOJPfVFYGkb6GvY2
edNAYVIGeadJpNYtDZW4n/KnEy5rIviZp0GpAEOthwfvoPGu5Ay56Z20TS8emsK3
0iIEkjD7MsjiK7UFeYVYzZY2eaImUi/XT/s0Ro/qYHxDEjjSWzmEs1gIFxnUidtj
QhTpEpQXUIZcgw43wkNMLY1uzAb4Yy8uNiFbEYGLhxHwgodehDQ73Z5WxZ8P8W2S
QFpFASrJVD+dAD+XUpY/BDn8cTSdnm3SP1cEzSibZE+FgIeYKcxwiLtXF9xfgkzz
GT1HYXqBcHGzvlQu+VAxpEdzZ4TBnaSb7+eHOrGzvwQNtZBXwSUZBUMsqbheOASV
hYQS2iz1i50jJwtlgUhjvncOCHls/yPcYrukqtWvazv6oAVLGBJYRHPqlNt084RJ
Jxpk4e68o94QrL5skQq5B9wzWYRU8uFDe9bdQ+48N48bAISmpgWJCWoT2qgy1LFV
GalCJN5uueZm98IalP2MYxNSU0vYBQh7KomSTRK4lSDXJJbKtnTFz7a1Jg0mAFwW
HSQH2wmGtutoKXR6va5j+ZJ+T50OFhlW3roQaafuA5qOn88ZOu7IkJqxVsrLBnDr
Lfw3LJgtdBQLScEHV+2X9oHKjpaKTvmy4NICUrIMLMJOIIK25hOp0w8+47KNA9z6
AjX75e1SKkqKZJoz17oeMqpvbPDl+4nHWgwS/HvXU5GgZjwX/HZrcw/IBlHSiJfL
lrDsaBKas1eP7/LTvBPRxTWQuOAa0SrRwqn+y/0uz7KsMgwQOPyLUgP3OV8Be9Nb
q8md+v+mgXPlXQENkVqeZIoE2+B6NqYD28EUO1hsfbgZvaMh5Px3ZngrIt7j4eT9
HR9maXAu2n1pHyZJhRvly+88E3mZIp8xyG7dLGOmFcb05ZWuUraH+/s67I8W5H2I
oXnD9CzIPxsOuXTkvPxmQhPuZWk4OE9W/yRYZSVUjeaAVr4CuANFnAIGuVcKWrYy
1nWyZbGj7cDWCqAq0XlAdjEFl6FeTGluul1Bd0cOn0kATQ2RcU1IxcVnMoLxVUyw
1uAJQma9zgECmKUSR3L3jKaPIMl6ryikboBAGBLrc1UkFlPs9FwTMncTeGA9hS+1
g9+l6zqWoRfcpzZ+8d7IUpDji+TKFPd7KoyuidYKd+lmlXctSsFmd/DlmuiZOSYf
Ut4kd2pB30HqyZA7KYXL+IV11BoUIXz5BX3cFsxFOHnc3P62MViKO/wnOcUu+2Bv
vo491Vvl6DMEV1pBZ1p6Ko/csa1648pm3DTE4knppPWzTsQUnSnXL3OvsoV2H0gu
oJEDiz6s692gRfsV78RBgh5+FxbhP39I+5zCbzIoy2WqpRjQr0dQfntrIOlza9ao
qSrRoxdsjQkFMFFNPF2uKzjva8kyv46QRmZeRV6GS9KNu29cNJfS9x+MlmQzHxh1
NGt8FND/lpQrDVkgHzgksa/rtGTFSFxaQjN4o8thYB7LzZJDkfDk3u0howQgxzMQ
B7Mw5Nmqfm5TkoopOlQAEwU9NcLpsWvfwtWoghN78T5029EzlpVgvLYYVxwlVHMm
3p5G+C4TwJy/TxwirOwmQfhBBvM17UwWXwiyD7zZ+qSdkziuGaffixIVMPd7JaOE
0VOUZiey5gkxh9jw/M2Qji5ugTG8dCN+M/UBhBAO4Y4=
`protect END_PROTECTED
