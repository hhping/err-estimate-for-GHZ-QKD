`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KF+Rx6OGTQD8/RWPA7y9EEvLG7jqsz3IeadT1TKuDdFUF58K4Xdy6rQLddodaF7m
vNBQQGBDKStEwnp8PCBpVhgdmc1B4YBXOKW3roS2AThalwTUPQBVE/NisCEL9IIa
b08uB1+Yo7niUv+HcfBjwNjwnPVLyqzE8b3Y52tOnVa81Xo9k+lSNglAm4t8ACMG
7TrwPAjO1uKmuTID7zGFe5AtvDm7gdnRQP/axbLd27J9esKjPyPovclVSJxxbVia
tEumjBU5SfYa4OFH0O8AJ8RfZBhECDK9ppKq3Da8/A/6XqiYdbODGcYD0M95WBaG
xOxH7oYLO3PmQA2+rdoePbThLjHj72ooz696wSxR2zo3WGajN0bhdPSJc31RK28e
zdImDkaZV6WWp3yLnzNDibBg1F4kXOj0Z3wxTuwvybJQSBUtzOSPBVbq9wBFwWrf
uhaE/7ol0GreeFIMoHJPQrLkJQUB282WqNW4UTTmWhGnECE43EpFxbvisJ/8D3jz
VH1GUoKVh8DBaF7AvCsWgsBDl5on8Rx6nH9Dg6/d2iT/csDRjk735hcD6sX3ataJ
wyLCyQd/oqHM0CQXEBGHRX6X713TllGQQS3I5Filub0um1Ialz22XbyA1h0PmAmQ
FPjfAQQ70SW00rLYZ3oG2Nh7X75iCCoedOIC/tQrrgCPl9QWIYCO5WgJDLQqxVyD
TAi9DOdgJLbc/Lp2HC1+qj2srf9mCJR8tp7q8yWjo7v3Yr9+21azZq2QeXgGlMTd
PLNOziSXgLF88XKMFuQ23g5ygNf/03Udc482M5174HziiN/o6ln33xjofVk1GJW0
ERL3e68D0PUrTFoOAeII+x3CUrCOyauXNyrOA0F1JnwLg3bXAcRL8uor+jgP+utW
jH//bO/5SWLxzTTVa6ZdyxakMAgYF0JsoAv371lwbs4jAOuFhR1Ai+ePKCV11gmy
qX4/7GSyoX7F8G9us0grnbuRH1IY0fA2sm0hpmzhPwIGtKklAGED7I+j/ErP3jVI
gzMOLTqf8V7YRakeO031NZLu/XLvQaerCzzAd/0fwysT8UmRejQ11xFNPOkS83a5
ghxO1QurcnFNwdze4cNgiRDRvtlDBZlSKSJsmQ5eKbwbJN/mpoR+3fNeZdD3AUxk
+s0JZ6RpE9QdZgu6wSshgIdInjp20idUCgIt2hGM/795R53DjjIwmwIJ5nhhbz8g
voZt/XCxS25q8N67soBUTPn87+5IRFMsVjTUa9WjFXTqVrGmpajjBB5AjahpNIo6
f2DhvFEeDwkFpXG0h35cYIuws0rCtEs5GASFPmG5FeDkrpkGkpRjAvGxp4vpwCwx
ovrxL37Ndp6/kwmUQke5E2cjXPfqGbuxwbYOhDaRoU6Wf4K3XBtKV1x39rqnOVnP
AQRfRPncpGlJFYyVp3Dfb7Cr962UuBX2RX+64jJWtlamcJZZVIWl8JRNNvrfeizR
L2vgjCR3IXNfijny8NlVARqFtxA9ZVIXJtXyxpTdnCD1yPe1OayJQg1/0Y/3Ukti
WoH8GZCBWMy2NP1dgWOTCJDXWhSyOze8J/Q439J3e+Pf+0JveuOcfFYJAvElgukT
rH8XsR3GeB4/5QwCyghmx3T341YzgOCTTLFrUe6MdWlHGDjngbpF39K4wvfgq367
n0KecRHAuV0feiKEUZIl/O2jxEq488Kpf3l3W1aXCnqA2wn0rCOh0z5CfybZgh6a
hH72814n+A4Zb3j8gWTh/yg9r/i8quU1lLKGwrvJ05jb/Dimv+YvvHU6P+6qWFlS
RtUw5E01N0HpibFp8YxlqCubbvv3P5lVX99H0w/KXdn5s7AWkyC+dx+tgfxeMmsT
4Va227+BoF4bG1Tk99jHaa0HgkATwc8QE0fMCs6EplknZyPNE41CggzyejNT3Puo
1OF3fOlektzfEjIof58ffYppNKZd69coHSu3+SsYX+C4loc54l1vlH6eH2Plxd9t
NYQenyb/sLpZjTodRErntkDiDL91zCMCco2W0UCXmgvLJewzqjEH50C9hJETCrdm
rvP1vfK69GtZLR6HhzeXDNAi/E4Gi8J/j6hHJ6g32vqxe6MntHTzQrNZJW0QMZYT
xRVm7pDX9YGMbhx4HI2g7zOtbjvgJM9LRbBHkLWlbddI4wF97d2vvLZsVQ1Dtbbs
xxif7bbQ1ST7WH/SEQEz+NQI6NMEDACBE5fbj8Sn9/5ldj3hL9DPzRq6j4KCr9ar
H8ZFesgKQkUZl90SGRexRTOaMRsSwmZrEYgGVUNgaH1k96f98WdA30Zg2mxRv/h4
nfbfILfWfWP6yXRBQELrBuB975pDLIV6Us+qo0IxNAdj7kbAjHxQwZNn1Ru0BUZm
HQBkqdDmRwCxylnUGvrxm198PHhFsxR9A67yyAebRhJfZo4Q7yaKBahBIU4rXoKA
1ghtlzrTmDGaHwwoZXThuet8tesCFiTbURwRXGmDE3bojrSXPiLNWgwL2z7/2j1O
UAUZHjcYHe619r3U/XYlYnd+ifp9VAHgaqoxUk9BUeXG+Fgq1lzjO5fL2+C3FzNC
QUFMlFCccs5CQs2eXwCuNdG/ooVHpMMZUqbrYtOgVFv52kAxpsppnqrHUuHehHyP
KAByt3+Zb1nIIVxDPd2coNTwMQvgtwNBF5hLWjcpH+BW+zq82/Gtzj9oNHU1jYd0
Md5s/ITR3T9kzrzLVSkmthCoFsq02h/hXTdYgTqtVgXEZ5uvFP2qgB7V502mV9uz
51GfKaxMQeNhD3RnMFig2eBjim5kVOoHPtuLNPy66HJrj77m6IfyYDuHM6XuvwWn
FGiOV6WXmEaU7YBwBXl957WOc5r8HZ15XVAdgs5oRPPM/8VjzZ0VN6ZcX+gDVQ8L
P9T7qpzfu4RlTHWu6dzUzMEYRp6pMAKAEOhDPm+lJSFbA30QWBF0kmPP0Tv5QO9M
KG1v2QEiV/KOTd8szTdXF7BWDxp4WgbHTfcAboJIaqjh4WoQ/Oub4GI2yzQbh7JU
qHzU5p56u3hdnHIUmP3HV43eX1k4wr1VqqNyTF6AoLrlkexXm+MrHn33lqzUL8Vi
NvjkAOOoj4lPpriZNw90BFlG+0PigGDzL1jZTQwsLTtAuHVx76OMS9ZLNnc0FUZ6
2E+nnARxAjx5WHuaLFGFz8DakGx6JRbk9EjCiK2C+buFvPOxmKtnNG8s24kDmccM
2oQIa32Jywq64Dr6U4XUWcQs/2H123KmRBevo1CFb5RZhu5IW2DSDyk4qGP3840h
WN6yX1Voc8jroaCCHJlfACtmSywPv0yNdYS7HwJCJsu4rtPouF7LGTCblFNhcHyg
iYjUMLDOTO9eCjkvv3oz5w1CxrMvST/S0F/ijiX9eeQk/9JbHIg2isJjRA9KPw8E
SdtRKvS+g1J1xZlWfK5Mt9MkDMFbx5qNIae/cZPFlt7T+znAlUzAqB++hRPrcD3J
W0fE5QDmvGp+D9lr03OipF1Pg4RAbM9KuhyzSztoCine3O6HFZBNprcCtA/jlzhw
PadN3cpqEkzhaoGynXiEXvj6UJMpS1MCapvI9GGZWDg3JRF+FXlNM5RVn4wKkGiH
odaxYYKY7IoK4PhIf4xwtRIsWO1vT2H8x9ACzMK/beajYBaVn7NjBYXj2y3BXv6w
qfBZlr+OJgMYFR4uq9st8ts5rnmvTLEmIKNcnhYwXAGtiLO68ndKrFwonypXPWgt
EObQeRVmcor6ov7Alzw+9Us2Rf2NNU7IuAjJjim+p12jtN/lfzw5AxhcNCFQPc6p
3JTgMNBzVesbdmNKQBfxMA3rD/mwWAN4+BF4PMMO5CHxp2P9zHk7YXKTczC74aKT
MpBe/g8R0bobf+uDaGEuajZE1Dlv50D0krgZ75lPWQAZZdW16TXd+D0IoEQpXr3t
3FnEli2aA5xpPZoq0x5eAY1TjS65R5LV58zj9QhnP13AyQilRwmgjOFX1A39hk14
6wJbUU+/2EJfffP828A5glblQO9iems9xIzqU1zcaN3fMp9+WEJFX4iqmbMsyU+s
cVzd9mfcqAygqYgxj6w46Tg55uOwQeIAPiZ3zVckbtCUOPfIyrG1+zFiqxArXXdY
1c8jtnbqkjI+ucHK1/pSeEOLKQwskP1z8TcRkvcQzZhLqeP3lVmmYD6K+OdMoSWc
8v9VFhSijexZqNTFJfv75o3Sz0OJzro5X1sKT+qRgvqzLzSOZy4hHfBDgR5wdShC
4tn0dgbWBBNcG1voiPsrSUcIzvC1AZbNEEq0AWDws2DHZba1xgSbRHPjAjrrGLVu
Gy8x1aW1zqblW4BKA8Zd6fAsVnm/jJPWwFf5tQahu0wwt/BedeDl7KXB/P1lqAgY
PUhWwRtJl//4EkdLrUQyh+FiaVHWFNhtqp7bTW+/uW8HtSLa/QWmPSv73d7KHTP/
T7Gcm+Cp4e6GFkZGAw+diiibEE9zi5jL5mVMhMIafmhBwm5bfu5o2EqJJWXskGPf
sKJRCPQ1AerrmJeVwGoeAQOsctPlKAtUYJt+i4hobsWXv3AQnSGyRgByscdXOl0E
1TrjWf9IoIU7S66A+f6yl4JuGEDJo1nwjh/ZZ0AU2CenS9U2Xn0/0DY9s/Sj0UrK
5snJ+O0IfPUTeYtLt0y2kFtWyF7FB26m4JEicwi4dWds6Kp63tp6D4/wLb9pXL91
9LsA8DHSV9muENdJMHVPQgqNpZDU07Z+NPfvcL+omXVCD7LbHbHeM+C9RfbcbQ6I
8yofU3dZGo7bIFPkoUIMuRLLexBxltgJa3TCJfSJ/tGTZwDvpAGOUUIusvhRnOjU
P8C9es6V7TvmZnxVuKd8Wc1sSq6Cn9Sv5QgsxlbxEADcJueh8Cogc3ZGadQd1Cr+
CIgRRjsbBujuZE9pavbULxZjo9hiH2a6WJP23b6R2sIRgObIvtkWO3Td7UC854G7
67Ux/Qc6vcN9h7P/ApxqBBtMD5ozz3zTmuDH8uz9fbLLUz3l2XVSnzGuhoyHL4EP
GqQ79iQLPgLgIzTtgFtEQJHose2lmxUUD59IIaH9A4OCoC5aa5hSFaR37jf3O0Yh
tJl8xEzAAMuRDmvbXfgrAi9Y527/lzs6+bqH+OSrXWEoe7oo24hifd1kB/sdpCsQ
lKUWgrZrzvcTeJVgEI3uZdg7Lo1y0y6QDZ4nsiN/KegiDqdItcrU7+dyfjOL+Do2
p0RQHe2c1ia7JQALAsZm1bdp8KDQWxNMm0XnfFBJg095WXsk2guP2Sjr+AdrbsND
VOfjUSBQFVgHSgMHt/xOwo6PuLexgIR79eunuUVcytuhRK2p9rIsAznjlE2GaRjT
wCXEngcuLA8kJjPkZTixNYizR+7drWVcNCnqLZE6L4eIzg7EdtBGo/e+74aKOl/n
4T/oMG1tVfNshE5ZGWC3tiCon1H+FV17JH7pJRwwfYvifyZZQ17nHLbWmYPDoZs7
0QokmcMCAX5doSCr99AkIaGzyjyXE3xBgjpjG9T3MIfe33TBUreE1W9RxoHPe5Go
9BVlP8avFnMSvTzdWJQoHvFEUaeWvPJFRW5qVbe8db/4mQcpVjjoWkNoaYEI1Sh6
Iczlc1D+5Ws/CnCZu0GaxQnggg08Oo1QuzRjKBMw5lYukoD9kR4OVs1mNkrxtSWE
YcTaW6F7MTJ5xQVQtpXg5ruZ9OaVjODzD1HQ65SAzbZ7OcA/jvnpJs9dAuehEka+
VOrRILz6SPzi17XovdxJpfQddesVgJZ4NiMR53bnil7fdPPVIWDanQ4qEhfWbiQb
9oPN0kdOJB9INu6jd5u/JWtdNkNu4G1bfhbUVNkEyq0zrjwl2YocaHDt+C806ELP
Q8lTu+/cIfmGaCfWdAO28AOqu9p+7jFCOP14fpD80X9Db8yTkqU/1w+EDtwGJxzX
J1SbTRBVIroul6h8nK+CazP40b41/mSbh4vZzDwIdD7sxmijImsz2fAasJxprZOI
72U2idlsaME4kcqj57yoBGxgMRBhZVR/m8BP1/Ga0mTBc0Oy3r79B8ULY8Cy6XXl
gAtitjdoYEpkv4fbJZyzRCuMm5W0KtdtceXQheDxqAEcs3Wd1JDAM7F1Q7OgWtjl
eRPb6OwWKH34KaFhty8PSlp//oJmnP9TLWTRjBmBkJZmEYriaYacUHHG682IDY84
p5orF9LBB0pso4NSsPK4aOjbCBLYFrquAIIQegNleYdoFVtAYMcskDiuqWSre7cS
JSd6B+VFcuPxUKdnsrVYF/JBmvhfuEmZPcoF6V+9UYNaO1rfglW3eU1i69KtT9fF
xNMP89bTZXEBllBKW3lfLfaLdIuKkS6aUYk7/9NW6OJBmwVMAmP2n/I6ti2ox+xu
Mu3TxfZOGebOPHLBs/iWo8auzrCrXbT7b41rwsk5GgZxKUNta3i6tFYPpMotIoKl
CMW2uj6BpExlzESkl75BNinNwtbDy0pKALKakAAer2vanIlGUT4w1Z7HKQRf77fO
pZgIgW6zlrtkoXzcJ07ACbE54vlooowcDSdsgiVqYJ+zrsWVhCdLl4LUDKzOeA2D
0ibyeLCRtB0mJCMSXja0UozQzjAgW3GREQjRlhDFwagiaJo4djvTk8dWMbIh1fJi
ls5VPMCtAtSKH/LYIGhlrE3a49fB0+p+d6HPw9H4RaiuEqXIbRTXMXyboc/17YQ3
FpqOBrJlKIFaBkcdZTltX5KoeJzkpnklLm3VktPj8J1b6TO550PyE9kKbxOgzBiH
+g6Y9a+rnWtJ0+xhUun9pgOW35paSUji8rA74U05qfxJRvg5nIIV9GF+YPS996BF
P9mgf4dzn0Qn9DJCNgCIk56WZ/vncTbDsoeP42kG4mgMpxGj5jsta5R9OHsw6Kww
bvOcbxdprZcmtdvqBTdO64jCP6NhSjYL8F181bxBlDz2F0T4Tl5X4FaI87a6kZA2
Ntpmt3rKW6CJ3ynsdOlvR7ot297BplmepDz69n3SacnworGIJpdhNRPuznOPt95b
GVJiEud5PXBycIUhDfWrJCzrZUIEf/Un5hhZMq1IhsHxgxNGXXfY/KG8uz+dkpHd
o9SdKi3/dDwkAQjaPH/5jyFde76s+o/Jh5gmGkh8pPC2lZxEcWxqc1xu3egGJuj3
boAqkyCMyjvJ6fEmgfK/09GRHudUM20VnToy7tm8WeCdKt8O6Ci0PIUeve9fIUSb
b5bgvY/FRrpgRjHo8HWkX+6cpmAI5Nn/nRk4XyWpd1embTo6t+xjBt8lh5w5bH40
lgPkK79ZHZHj2+fq1rKuL8j8AErzIIKbuFAqvJljF72ADQI5j2sBdwcSgrh75eLf
f79rOeznMtjqS8WJ4kuTRILUtPVmxzCi1Ws/jT5fElbXOotm9S+RhVUUsfmYDkmZ
Q1llUURBlX2upKw30Y5PpbkRJIxaJT7tIlaxiCHde9R16a+MCsJUog4UZW1R4/uk
ZVkbMuwMFm8lGd9AIZ1YqhVvXAz4orFhmvg9K4CY3CiDsSL8dslME/F2pL+JhUKT
Vn9huP1vjuWxtlILbgy66PhMzgC4ua71dKGEdk1QKBERYsvBZRV6ICABjed1Si7d
RUxLhc5IpwTMj83RK9t0B99rJH5H5DFxGx2x+FW5NXOM89R69gKlYd6jRzy2LDT7
5cv+OhvV3NYC7GYs7vKdM/LdgnGUSFRtI2McDORPTd0VPjuhwWjriaotHvCxP+lR
e5/dOGDyk5H8P2fIIORriJbcMagHtrgLLUB0Eapee0IOu9c9xn+zFZCk8lQ2Nfrr
+DG6j6EcqNvGVcUIvWTY5ysOxR2w548lmOJFECxKDK8yrXG2wTQbGsHid7cJJd1k
BWK9hVGGgF6G0OS30afu81UWnR6enJ1jN/7PgNO+O/rdw+ewzGNgksEzhqCzMgU/
gzIyWm+pjgcEEzFLd+E85Mra4V6TUVqGVKCb4We1YIxZvXHKuN9D5wcomGCw5Px6
cHakIJpsYV6unYiWoehCSJnlrlGDnQ2oleUwuC8zJ9HABwodoN5XE/9dG1gzshId
QNhVjSombnAVQhnBS91ivR0bTzZKTp+bD0CUzHySZwi/wxB2un+WaU2A5zleUU6D
PmO6RsQYFY49jr1PoVH9QGYtblMnj74l3lzhk6/tU7/7m9/PlBZUr23S/T4HjG/z
ewXvoUV5jkfzZOd84JV50nanBR3CBFcEquxQwk628pLZVtdRFQTTRLGoszUwrGX7
wOfreeB5B1zo3Wlfa2xY1uqKYmRXPq4gbt7gKgWOh1n6dPkKNcONSiSA7M5a+HMv
yk7R/w/SSbykNRup0sxoWzAmBJG7vOMpm0ik5K/lGoX0C61cO0I0wr/zmRlfZ0Wo
Qw8HygiyZKQkxDzebWuLG5V9+iguxoDh6FUtFeJkrAhYtvo4uFaLygdDaoPm6M52
r3Y+YQ1xB/Y+XufEs1YzO/AfNjEqUP3ZU3aq8q67Yb94Ntb9Da2EgyouTBePgSv6
Eolw2bCnVOeE6tWfaZUxNf16EDxXVuJvg/w5z3oc8Y4G0HGza2dc00UDeDRAoyd+
2/xvlEMf3YUSsf9V85C+ZnC4Qzdcx4J976JrbUJyCe1GMHt4o0nEdrNlpvyZvCzD
nXgiX1MDqzxPuPXpmp3FKA+kvRV8Zn69S1u+BwO13EPWXs9ach8rHtk1LjtenVKP
YHji/VpDPiYM49KyRdEh8H6u5iCogBffOYpaEfqN8wk4uD06A/wZ4otd0uAulEpd
IH7ALdgYpavSlo6qVPaTS+I2pMoRakhAXXw7rtR5SziwtP3Cj3zk1WKa4gliA0Y1
Q+6xn/j8Fv34sEEvLrQaJ4p6+bS1UZEtP8kIzcPJyHbC8iWCi3dKhL/FQw3x0QoJ
6PQoFLBLYrIOtGHwwo2aVB8KOcVRECjyUKI+XZT5I9dGanZf9yTYlA4SgYXpyud4
H+MSjCHt8uBgh0ZlSx8G4Q7lPrQbBsGI/WQQj8wt/ABUc42qe0Zmo76EUOC81ZvR
68XVS+rG8zB7D1rRCr3hnhFqkeDWYv77/Lo5xTx3ZyKJvjYemHbCUAS+gwdyZDvi
ASTaL660TPJ5xZIyi6WejuFJmrdDTcZ3F5h3e+XYQOrtgiK7tfQ3RiR9Wi0Fd38W
ZSXhxtnrvkmYRzjv4Tb3335drZzTsRfpbTFUGMjZcCOq+sIaWpqLjPGbQOp+WVI1
Ox5Oxqj4pJkHFagiYahBZko28v8b0ALhRC7qiZstZMFaFeU5j7p6n3o91GUaiHIF
kHYccagrVy1kdtkZWPDhCBW9sbQXP+KGHqFBK+Qc5DL2oC+wRegHZIwEuUEVKFQt
qUNZx5h69gg/Rsh8vQoLfsKFI7NrnLZcARpTWDPh5IeusvDNA5OIGCxvLVNwtWqB
HAo1/+pOaw7meqjgiA2mvPKLEsIxurju4bbc79oILhUABNKWUQpJzo3SrOUHBCss
B3duwJpUjoVkbFs8WG/quec6YCMpHMNzhEYyCiJ2LP6IwZJxGEVQ2z5Zp9azi/PA
9PZQ0LZYxtnUbr6dNxThzCr44vaPDBCJdxIy9fQHgW54YdD7PFobLVAPG51kVTOi
tBLpMYF4bSwTusZBewC2aca5+7Tc00MJGSUwjg2adQJY86cNZxWEFbZMwM7cbtaA
9QRrk5fPU0eg0y0Lp48DQJNYq28YlD49rKtBAfAYEIC2en0Kt2hU+ZVZYGJQdc99
deBYG1ja0m3O4YccMLKg5MzhfS+W5xqZNwRUviC66edRJ1QUNBbOPEfPMjktTDgK
QbxCGPoZUDKGAPBP3BBz7RfZH+1o3BEL090LmZE6k627ghQcqpgS/zfh6GBr5Cjl
t/UcemNv+WF7ORb8LA2ZtT/a1bsdkSw2A70pJrbxIZS7C80QgNw2/OkRZXTSLm3N
70YdE4xbPszlCugzM9wbqr+0OePb00eI6kQDECr6ng5/nPHnfkf2jPAe9hBj0nNB
cS0QHCpqEJGOVRJo4UKO/R9JDQi2Bu4y6Q6RD+p4LqXKE+Yc8regTniqrEZpizfi
1RxG1O3LvNvqLKc4IP7uCsIKhl+usK50oz6odu4SXOKuo2h0ZUkj/RacF2v59tnb
a991md8CXJIAqwxfPpBT5w/3ybS3zJ31oxKiHLPrkRtEiLFZcvxc7qpZMMrAd4Tq
GqOtd1b1bAyJzhjU0E/s4/sb7d2IM2X1nBfSN+MJnWw2s0WEcDTWsYHUszIgKDHC
Ii3+U/JgMbK8ZpCHFB0WqAGCkmuwcnWkBULE0/q057RkoGVyKgN2++fz/1jqXgTm
IG6NobTbFWmTke1iftri/J+e4lI8m/qkQ4m8dv5Ma7NzVK+6FwPm2aqWPOydMgM+
W4QQWaGfH/WcdEqiNpr6PWBRAJAHVYsbdETJ9j2BY9IJPLpIgZPh9GEddL2+M20Y
GEAnFaAY7Tg2tnm+IHqe5WMAmhCJtzoO5JrHh4iiQHZ5DO+8ZmIAJr9ZP4w3j4RD
8zqkRsCTvc4T+R7tcQjqFTTy91gZJw1/ieuHuF27U7wdJ+/qAgsIRf/8IkseWrpt
PBdeCk5MjHwUdJYwrlwgU+GwsHinoEZIVO0g4zCfa63/N0FZcVuRDnUVlp7NcjcM
vf/86KiF92USF8sS95XgcaMot7utBX5/KcQftg7N94tlOjNUzftw79aMJ/i+G/3j
L+o0kIs1vNrTC/5fL7/6toFCrbFPIBdV4MNmp9PNUmehOAnRv1CZlWVvMtJysYK7
z5vec4W9tqp0J/o48yzbREU/oV1URsxkSvLzyR3+RCmOQU7Z5nf2WZk+34KLARwW
lV3zm+G/M7GShWvRUMciBkLOB6xENOQMdSAfnV6X+HxvfB2oBf8C/gXeMIbAka5G
UveIX9peG2JKvP49Vsawuw2ArFA6BQA6RdlIUxm36xmUjIxIC934fJIJKW1yzu4Q
wZ2C11CbZfB5ZXEjJADZn1Q2vHwrunoZt9l2weTIhKwSV9vBmxk/ZYxwrXj5XPkn
SpnSGgQx4KsmrPt/T8PK1w3f/BretwfFazjU84mF9GSHghuBJZ5H/c20jAXJcKwY
AIk+V4dxNtwFp2qHWOy7vK3Izbr/an29mV7zUC6Mic+XP6KJyh/ieb3ks0gP8W8E
Ty2X7GmKD5/TgmpeyiPGLvBJtxoxOi65GxbfyADuyk1TGt9hatMycSDiCrwHK/xY
MurcKSjJ6TvrPLuzKrxOrA==
`protect END_PROTECTED
