`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4WCidN31K4BKPPJbVBAGUCZd0kfrIAxm3Z5vTBCPWapOUiDqyI13mIDmJ53DblIj
Rm3LB2KqSCmrWJTrSUHkc7iDl346hFuYK0eOyT+Z03WMJaqRT3AWfLVPr0x5pdC5
HHYSQRRzmi7PdC633gzm2MhySttq4bRHD8XGNez0cb5twX9Pqfr+ISOrGU28FiO/
HfuLwimQFwDCOcWmtiBV/Q1FaCOK/lX7JuyavGrrhTfYda51c8PhhWXrWO2xHTDq
bSCDj/2hNtbcsDbWlXNPP0Vesod/CuT/Iy/rLTWmMdLjopBeFUbzqdOuhzaVT2wR
4ITnND1xatnUYrpCoJZK9A6VrBMzJFAgfXLbKrQwk4Jl/McGVbo+QMMmoNMVAwO0
8w2ZDlypFW2Z3nVtgTw18ItSu/Tm5R7As/GrGxbLLIzdLeqFKVhezcUSyBZX6xXk
NJxvmX7f9B865wxe7jkK/URz3uf03074R0axmeLAiMWrACCiphEMPs213h8RLDSD
paAwNXpsqBj6KUpiu6wT1r/cOcFG91QiW4LaSgkXats/nW3ZMa1b8Cz5+1o17NDD
ySU/mgLkdawxrGCYcJDcb4lCombErA39gO5o03LOJqsSNGn0yZIfkrgkiNLvU0dq
DW8WNWmZPyQJ5Vr2oyc0U9N+RNErfK1j0cz5VqEMhbk3zrprpySO1JZLearLU2Xp
m4IM7JSkhyMpGpqG0eNfkKs99oOR6dzhfb31sMe/QCPXTR4II/1ykwq+MeFQynrL
aMQG9ZTRTSLKQYX/66DeYmFSIDdUhEMHmlOnDYMFBCf8Cc3FdqFiAJN1Ec6bpQH5
5xazAuG+j2S+bOCTB9VjxKLB44b9NwJnCTM2nVK4Y+9CR0mY/JOZMLW9aQbJh3cW
S0uS2hB1OtgHSy0ojMaJh24UOi4JmvbMkaqB7IhExsx2kUqpGcbPTVlIIU2uXXMV
FgWEAMZ9zSKnbBwkVDfaA1dxXg2Wb5CmFezT6emAc95FoyOdLV3TH3rRgv3vnef/
AZv3WU48EPH8zEhemVnCAOi+pkj1hd/dR7sJ6oWGg3RunASBiDhlYp9RfXDO+07O
PvlNqOF9SLKfeRffOtHkUryWyRZ3D8f0oZmLyUxFheFH8CjHBxsqR1PSKZn8Wifn
JtxtoIxmkPgXX9JKnImUHwOVb3xY0QT47wbe2b4bjx5yiJotgpvig5mOULW7P5Jb
kE+fQ+POSsYY32/6HzKR65ERN7bKZwkle+n2roERur8MfDJNZiIoS/yRhnJ8UkKT
RYtlYT65MA+3cz8PyTAEfzg4qIw+u0ChXZN++hm2eG4oSOEHIRXpyizs3/95qPof
GaQBioDBs5LyNxA1jqtk9IJ/c0WbdjB/3WFVDM7G5Ohs9oWmIFG1ugjLv+8casPe
8wNKpglmu+mQcswEkZDg9GWeKtGLFudUBAAgFvGGm1R359/0nEW9M8O0kyCgU0Xx
+egONe+wNzftBEvxCADc+nQj6YZGn+/w4sDDwZ/na9P8D+22qbbYo/2wFhuz+8Vq
DxeAd5WipqxYT5pR2LyXUaaA7mVd12H/DhpLTPKlU1tGdnESSIc+21j7GO6BThED
5amqNfNKu7biLrdXLUoXVYFU//dhSrXBNwGUqlWdVsxDUO2Q8hHXNYUXAezqP7eW
g7RZN1gNqwg08YN27OMnhBv8pUmMcL88EUoOvmKpCayMSueY9bBuVrkpmSBcCE1w
eKhqIKGQzJhs1nNC5IElBPYuNX2FvbjctaIshf+8qxaWxM96FR34O365gkDEpy28
rrCrHGWR4YBnt0VKlAWXNqD3+61QZAz2Oo0OmX1eoyuUsk8vKD7odvqyMJmywaw9
azZDzaizZPOEhygrDx5i5w1XR+c9lmCkRBVZaj13O4zerSM5ygiwQqWSaX6dLxbb
gkvxLHhXlC1HgZYFOp/EKtHucUUzl8XtVaWEqRct8ULH84Bbwjm14lEqaVye3TN7
6ZX+lTFHPgdqorQLjVPwJ9autb1KQ86N0VPKOT3gnAVwbWbnTuDxv1/+U6qgWVbO
nRgvWaquu7CGuIpmg2Z8xc1s2WpYaQJfVIHQUfem2apLSlsFjf1y0KNjqqwyfiqn
kPVRCu9++IJRXcU3C6sMURM9R+BWZTUtiDtXDJOyHkDeucmfumMm0sa8Bc+rMVFp
+BZhmle9ioI10r/wdemgfBT1oh+5HmxGk/gQa3bGRYtPoVSIeDJ9S5yEyRgILyAX
sivleIwWrkg94GM6zuqyh6bmvU/L2qioI/xPwSdT1Gtaal7qIilWc7pvjuGj/7gy
MDvGAiZfyeq4N2dvTwquPbuKzR/g6zhjW+AHFWMBbCNnVWMPvjILzzsDsmoyk5P9
ntv3OUut77edhvSDq4xeNEb3kI79hBoCuJb6jrgX8zm/sLQpn3weMZeTci4oNDiq
wyYNmn+WzFhwtbFFtvsUjk5igCGr3DWPLaQwXANMwpugASkEFL3dRveBonvTa7tr
NsOzUnZ4A+DVJIMtvryY8TGERidFzi8DiiD6L0mkV37ovAt1Yb3WdjNpvtz7BzyB
DpzRRDAOHRwp6qI4TjNi5qWuhon4b+7jPPTgUR/FvCLYLC0nlRb68DoQI/6NqOyR
MM62aEmeI0fRhyF7eOBlk6CxuNrle/2JIsgquPD+hcYsgAshL+cDulCJcffYe8uy
NnFEW1VPOEi/XxnYcjtchjt84LhOgjyD9m+u9D9lu55DPMetEZu4CJefcnSr5i9G
gPisLVhUjvRnt1ykToliZ1/+qh9aYUsQoFr/o9cVJSSKEkMJfj+q5qM7Vzr3tYFX
iEo+uEMa3OtYJ3ubp0CaBxT3LD749fBqj0CxL16seSFsbJehhd9qIzeJymObzamC
WQJkR1XJBoDckIQ2/tm3iboDWptWBLvWuk6sDy7O+yFlLzcMlbpfk8B8Ae21ZuaA
2HSTccPKrzFkxxj32/lZpfZ6YpBXo7aHVqF8QNdqjguvFaGgGNDYvtTskjmWG7gd
LMtnM7V2Z2JiAICsaiYCnGX3zTQxU3/ZNkAYs9AaN6z/yyeLJknnmO1J4x6nmP2w
4i3rvnzX/yI8uOrt3OX+LXrjG7txpSovXJGIelQMIQrLqhgIgTC7q5K45hUoRmsP
ycBczURzgZ0BCdhlq/nRH1Zf596NeErEQ1yI2JSiXKHwDpiC//6U4LCc9d97rPII
SkZWP793MzktYLmUD6rhIaU0x1d/IAjR5kax5oDVedgMZw2jjVIOVztdqyFkUuh1
ZqkzKyG3bxBmGSp71ctjbDbue68UPBAhWoSkRYXN+mEOa516quoUEt9soonH8y7B
er8m2HwHL6tdv878Sv7PqDGtD5+bbxQGtXOW8RXhVICjLxvf7FIpbt6TCPB0Bb5v
zlmpf81PnHsExgYxM177b3KNyslf4hrMFzJYS2d1jvhEIdKo6qXDKaC/MYu1JGYt
+ScgHCpqRxH8fCKk6K1CZcm/ppR9t3brw25b44gdkBsOrmGSQqzg5caxJFOI14x/
BSvNpBWfrLixgAcV2Om8fftnxddCRpgc9IBpMUi2qBAF6PLwmIVJHRhRLwkZSVIj
oud6O+4hHdukWEjcX8yl04ac9nsILfDl8Rzbk1bKzjxb4a8zx5PnQt7adcPi4AsW
RfnJbRmb23//IXEdCEPIWixCCH5WquDt7/xwVyHffWvsmgJHQDTs0R7YAsWx+ArC
8ZhwVS0tytUNz6wwJ/9XxnU/J51/5r2q+HIPwg/iPnNuophodg9texALRT6ZMSdD
3psUDdCHoim6CRsU9PDwFdYOU3q+sCy9baYXbyq35udE/lRUUO2V1jYRwmTTmsaq
skaRrIVRsUSMzz7I3J0JrnJ/BH3ctTvGR8BnCbA3cLARJCy9zXnzBqrGy2lzUtB/
ewxrWwIdTBl96awDfbakceLq6yXzSFvhoq54aW10cWBkenRL2wE4UMMiGtEfRjqS
ohgnzWctMvOG7TkpqgzdhiJJQN5h6Vp6OhfBumGUQMbNE9n1LUh0MXZPOtQr6Edv
Fdk7JCR5eTqpB4Cs9dw9IxCAHWjBwMBCaXlilD86otpb99hswIIAKUmkquhl4yMT
PKNub3DvUIQhYz888c+J0tZ/sKRxC4FH/s7KI7PmM6txsde/70V7dOrfRmUN5LOi
9rCspz1PFslZbeF7yGaw0DGKrCMueM27XWIoO6SEXYrNbQKKYRBHGDGMCw+p8cNk
8X4pa8YFoyxBIuU41UAIU/1sKa+SjMI4zRrLatWGgJ4M46oCXIgKnRyZp7GTaxT8
+Fcw2dj8o2z67qRURvHm0WlPWuNkaICaAktHTK8I8In3oxp+t01WDMbKTwJTRZBs
w/rN13m19t0fzE9NZauUotBWzK8j1aKw31T9czd2sF9IOGEfkspzIx70d+LgoK+d
Ud+IqKFwF9LCMYXr3bd1b3IYAEZvUstCWJNGgsfhgatSFkd9A1gCkUtb9lv2aNe4
08C06vp8+B3S3+MeRPRf3cNhxTAfAGtBq7DZGR+z12AK1jy52gADFArYsQPy2ZTS
aSigc5fVK81gJBQ32so9rh5ZM9MPHrev6kxp4/X8qB6WNBypCtnE5s4xhU0NWI7j
15qUkMN7FKhlT4lXr4GiI+LNcQKYQUbnJ6Qh/PIKsOyGspJLzd1xJWoP6NH9fNIC
BiJgBS9gmJMPHy7R7TSRxbJyZvGMHLRcWkO85/hHgrF1yqaatfjgZNHpDPkm0/rA
/d1TzEVpLdZVAz+ZTgvO34xvCut3NCwkT2W2Xlte9oazv+WKmZOj1nRDXGaGIruz
t1PsfZj7fsWaRDoSv+34dm3H3IU1QgD4Jdm4ePoh1bK74tvMfEGtMyvaGlbeN63N
NH+cMQGlGctoDEIQwu3Kqt9E/gHBGzUNeeoaYo8E0gUNMcDp5A1V8QHNRJGzsIHu
ML63jt6ZR/MnGR6Do2h3/smeGcqiypH1ZLuCohFI0xE9ljVGQZif0WT/T8x2St0V
10ld7wET01AM3viBzwY67DKx0/Ipv22xT5Dvdhjo4S2vKlWQr9UU8mCDz+2CPanL
JnYavAqA79oDwo/A6q5rtJEpeE6WFB43/3P2RcumouGEs55PtrBLjQKsL6jIooIJ
GCuKIjblVmwn+MYz1CCcyhZ4fPslzjdCAvbhs4CXsrPVf0PF4iGI31ufZeuUuABJ
Yc3y12ypipVZy2qgWx9SQqPDs7egKcTfKE8eosDK5oiu7BI8DYQQ1TzG4Joxh+Y0
ALU6gi6Gn1+Em9YGvCWLaUtT1fPZNWa0wDoyX9hkLG5wbufRsu6x2AL+2MZJ3beq
IuqR2q7Dwz97k/pFzngS0g0v74JgmLwGOzlLnNc6kk+wWQ7+q5aTSodV9neRYGuN
7ZWXr/ZfFm0coLBT4SIG2BS4gOc5wQDEhuId76ZeIiz3S6NZmWKfM86GNOibNoZ3
cWLCdTOBkuuXRxUaWVB7Q2Vsn49rj39L9bDNivhw3Ti3C4pB+JwtGwtCMpcnnwHX
AKpt8GMDUW0rfZMTPIubdvVz0mkkTP9Dov9g+GVFHYFXeXERwPG6z4SvXmvcXTmH
SfS5uTNANJr5z7mvab/XR4HZjpMQ6iRXTp1r/6aVeiNMQ6RUsy5X0WA+vGShGyHr
ok2Rxx8g0TqhpLNjc/9d4Q2jJrXFx5Aln7W4QPwX0TLu4UdbgjzExAsiQdF8FzBE
lrVq0DNG6gweUo8bSjZ1MqME6UJjDT7xNrhINNLVjnBjVqdfNn+GLsc9OsNkmawM
EtoWq+BPsTr3+fp5uY56GsK8ts5aG1qVQtWQIBVzGRqWHAiC1MVs7sWr93KPIbPY
cVb94WXEDNVUTIhiRiUwHLhE7OOqy6pu/gqjkKKle0/H7ipS3zvlqDHUvN+lyz3n
l6rqE8OvXaNj2WmODxAepWix5BQlKWwWMSEvTg8X3nP9pAMWGP7UCOzT2UBUnUsR
9XOUEzpXPGGB0tE+DFHfF1a2iTJK71darcfId/EVaJ7N9lViG0RFu8GvJ7gg+vxp
/GqLzTb8znxh3Jk35suw1CI8IQ76c2ywBOC2nobtWc9y1BbLiYQQ+fIJJSzfs1kn
YqTSST1w8dmzwXJLsIDApqXa5r/X/iEgiXe69pfU5YPPZt3rRlVpiSXlTVcLgW4H
aa9NMWZ2o7jky4JCUdogCyQl+GLaXdvksVxpDbZtnV+i5+0Fw2DRuMi3rslOIdNl
tUTXSdsgeIee65YKMxq415bHBL3IY02ud/9S4tOQV0OfPIVRnPa9cY/XaCeYYby9
EufnNmdIbu8LIO5QPcsop1W94hBbBOLaw8QkdRgmft/zcpyz6JL5NjQF3apoLvQe
SlM4c4GbPkwj1btmTp9eQfKos3va0X8XvXYH92ldg6QnxGww3RqSUnMyit4XcM0s
xEVL7VcCxhBfflptc1GrUBQbS0BRy/Nw2B02MVLUq9E+hKMEXIpbeVhMIxv/Ff0m
fRdcv/C2topx8Bv2pAt9V2Xc19YMvqhAWrDSguQQ2+uvykeoHjPplKSoeOl9DMqq
YaVnHehFS2nfiXVXJ9OyB6mNaIAXviB+q7BkoCUPHbd8XsJZ6dXWWbrKF764OKUG
fJCOSySPBEVQtKQo3aAA8V4Uz2lc7ycS374JtPN6lA3WntZYaYGRK1yEIhhV40PY
zl8oo/9myngPalavB0TbvJBo9deOxMotX9YUEa+UiCVqXwpAeRimOJEuUrN0ngnb
J8xwSYvOyOpiRgv1IlCTOz1z6bWVK5Rvgt1ct65VOYrkCV2gLFfMTKCxOCWyRRKF
1RHn46HzH6JIcud7Kytz5YmDZRf8u0isDEmJF9tzbkoyvsSFn+owBhplb7ptBXhC
vkjilY+14/LpSOEOfDWKl/+SndPt+RpF2lr8bTp7wr6cwFmltMv1uZM1hMd/rFit
OWgteMmY57Hh+nlPz+j6i51a+g+S7v3+/eu/OE9NE2A=
`protect END_PROTECTED
