`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n33nzvVNbtoqf4R0RXJkrCUEswhnGD54y8Sn61Fwdj++MigLUq3nEQCdwx2xyUGg
vera0zKU5agL12w9RxvoVIN4oX8z75CgGUoe+2fbSH0vHIg1+tmCREDGBsM8p44a
X4gzjt/gbJcG8GLbM5HYYVno2LTdbL1HNRpNwgTZJJsmqm9EcO9TvwExjBTzsF0A
Yf3BRydHGWd+R5q3psuS8IKlyzuEKH/W5ZJso8DYK8mNZBYwDBb9Z9ZWXtH8miVa
rwEFL10wQfFHqJ6aBvTKblSb74wo0hUSttZHpHWj1P0JACkCadX7cLHYG8n8haWA
qCC6+oayuy+wyKqUxeZ4xZiW3bfWsLapCCzHg+NY43LmwXcFciqRpEbi8ZmCvcX9
SRCVU4CkmUz9NgieGHKL1X6uQXo38JDaPPWRCKg1lAnzzRC+MIs8qaXPjQMV1pGX
HR/7E02B/8tGQGlC4FyoYxcAZoH1v0DyhUHaqeWYwLdvJE68uaEuwdUy6AC+s9tw
nLF6Z+K1Etcg16lBId3aG6e3YGdeRC3/PHv1X1a0H+akLjVD692SUlLPoYqFuitr
ol4PqD574PZKiWFYypCkhJQks/Efa0EvnQHzrLlCrKAj4EGAAp846DVsL5eNhsO9
ufthkqEGAMTaqN3GeTXnxlPpBv308CbtZd5xUQB2O9mP1anZx8wuA/xiy/wEV2DC
xpjuH9DjsM/KkmovQlxN03fqshEXS31Y92m2n7iX0dsaF0kgwN1LriK4LoFiK7ew
LjENOXb+TxubTH+HoWJQ2K9VoD2xgL/wMdWb9hSAarS8uOU23GgbeelNZuLWU8kQ
HSdOxj9C3U7x/s0afifM9Zr0MnvhD1n61/rJf1Pguf37sXawgfrHQhKJ/SMPAlKp
oD18QH8GUjSSs/Ledz/2Y1APEbasvx9I14thRkxhb7S1rj/zInN2nyXxK4Basdx3
PUBbaCo/l+SYQpaGT27S8rc3sOgDUpaSpZI6JvdTL4m28T1MjBBCWzEAjQgpzOoG
bNaBTb1ME4UAl5NS/UOSOn29KN0xq+n/yEHX8TV8oH07T31dQc9cmYyi/R3MYxzb
MF8OGFXQtdKSGobaH5RTb+87sIC1mbl2ecf0bkeZcPZw6CpWjK60MWJo715DqABx
gUfMl4ScO5CHPs0FqaajsxZX5JVssrd975DRkfrPI0mBos5vEOVWHpxz6zH+lmYa
fersezm1DvZS8ZcvP8Uf7kqVkBLXWwtMiQ/v53UIZ9t/72j6jwbR1YshGtWyPPbO
NcPAMhpVkdmnlW9yoCEER67ufG7u5TN3jNHSbdvmtMmZ2EF3Q/YE84JgYrmTPsU7
+6XZNBeaep4HdoxhCP+bx9ZomkR5Yh7MXwqD5xjeAgtF3YAwbBj+RNExKi5g4ONe
oD7YKy1sF6uLKwkFwSruV+RmJL4jv8s4d9M3M3VMp8q5+IeFW8mMRwbcs+nbc/Gj
gQ+1AgSQfn9N73kHABtIGGGhU0y80WCdEK+8F/HgyGRQIPz+UIF0y7M4uwXvQUnf
6V1kwfVDlLS8FOrm7JLY/2a2ZGj7n1WeQMJSvv4ho1R2nBw0xLk1IlLn2AvyWle2
5jP41WQQpXTPtUoIxx6FX2fSMIb5YHgR2eg52/7jcsyH8VxXbjBZxBSQUbFlO93I
hZMBqY4Uqij2rBRVoLS4IZdgulcKR9RrftXFHDOOhimws78ZTaWZ79/jFG/Bqn4R
Y8h4kpiPfBcmx0+WKD/E+HMB1sN4UY4/nMeZqjS+acEBUZ++Q4sVJns3Q0M0MqQk
B4K0Icpc3U418D6Zln5qyoOm4p9gKTzjhzJXBQNl6KMJlBk2TXrmf551/z8UT0tQ
pI8bk6gzLcuVItDR43Loos6Gp0TdsmZzgc7UWhvGBod4vmS5RFh07elZYreM4N6l
qBXrijEcQQtdkJX4sPqLQm9nR8PCCBr7Z/cgpWO2bD5DdGmk3g2znTTMRojdHIRX
qY455dgrA53qXbiSgx8WU1ycY9fa/Sgv/ySVsEDjIp8JM7AA4CMcxG7HFcRacTDZ
veCGVGttSqXybj7yXqL0OPfrVppKAavAELGbdyUrb5vH7qzOlHvUWe8WteZw+a4q
e0m+VYAn3k6Y6oBMvqp6KIyuUyWlruPl+gMqVZ8dJ2qSAJbQonY9wviUsWMbSZZb
U97KJ63LR/hfnbYSV02eLjOXA4gcGkjVdTqhBnEQDVUfau+1Lplkkq9Z9YDIFPIr
f0WG3fYuRXj9A4XqyqOUs7QMdvEV8evWb4LQe6qUWZpf84ED2ESQvVD1lLN2hCxr
iKHB7WrpDPMMkwOV7ZpKwRdTFvBdYlsF9H2CrqK726lXUUs/0LQi2+vdxHfd1Oib
oVA8EJFuuUj0Tl+hZh3TCtvESyCF+Wkxp0z2H9DbdcddxP72PdwSUBelUNUorjD0
qMpBrgDVfswSGI2J7LIG3W6GxvCCN9oaff0qPQrvmd3iuMqYJI3Lu5Rod5C/0TWQ
evTubQ12QHufYl6/JHVLjfzFMKlSi9K4d1tbmRlvGAvo0P5u/bOGVemLYjaTtWOi
wIXA2qrG0em0GRJjYv2nGwHVK1wxsVQT3LZWeT2FfcyR/qXiTbOhl5dhqd+UXvBp
/3FxPNfYf0dEAWcKYPoWmQhS+kehbU4U1YIBtjTKvb+r9d/zgkwQ2/x1CO6JvVvW
gBUuR9oElC/wCwkSMbuhL+TmN2sGZ2r1ks2UuAAR3f1jX5TdXfyzLjsSpqYJ8mDZ
7jQE7m5cQyn4KIJd7qPLPSBv35fuTZxLT03jyeXz+dJFxm8Eh3i3jsBZ8L0vjxme
6xbq7biPRPhdCztRy6bjmcZAzc6CLzgchgl413xbVdtfwupsBBlRc30LKxt/CZ9o
VQzuYra0qZH0PVi5jNZiFYhcRhULkWzfZcU7ETEgUB0AMIZKSMMA6gSU9GcM3Msz
l4NwuGF0ZlkUhxcsLAfef0Vypvu1pibSA2yhrc090uCmXxLr2eODhed22EwdMtHS
Bbio2vF286S3PE7mD2LxTVakI0ILF4y5//OvOMXL8S/EOxpOXaKMutyzuwT7At3c
SgIJCOhh0wt5TyuLf6pvkKkuyRATYX4L0ZmFKn1Dw8cc2diEhjwgb8IkdIozjmpA
zGu5fDITLhAWL/0W9qSOq8vbQiHLanYgVwP8pAMszae+qFxrN5KG3NX5qS9VeqGT
HPUYDe+ipr1W1lxhNmxc9UgGdPITZ2lYeBlz7QaFzAFSA6cASPQAHid4dpwNQ2hA
XLGCAoKZRb9DKnZ/NIE1AL/otm5jomK1RqKQfLytRmh89EmB9nMjHACcheW4mrJv
auurcbQYjl48aTUz+dLWJK2/w9J+CeeJsXGIk7CkdBtKilKGCHMbolkl8SbiXNVB
yEC1H5z7dIDR+evOwWkb6bUR/fejQxK+0yRoZg77JoM4ncIgWEjQY9yrvP747+5U
SHIpKBTm7FkFVqyysQhRgUpQEZHudZpRJAQAA9glDEIAflE5lik0RtmEJXJY39/4
BQ/TtQlgn0rsYBJ8PEaoeXhbqFH2aHdVrBN18Wo70BuHkJnCGF796R2QNjfgxdYw
NsspqImvzN7tH4Dj2yl+ijZn+2z9pkdlvKvC3ZqwPJKghXpb3zAEGasLZIR0a+Z9
m0uwvxHrcSNjsUu3S3Erewk3mYI0idJ9eD1w//pfBXjP14TS3mr1tEF2YpCOHvQl
zJtS6qA+V4WT9OU1IV/+K3zzkFuJtbXcjPIuTFe3/JfgPSI3JIyrkIvmRd6edNRH
7y1SxnzQoaUGBHAzWTr+0y7gZwP342fGXH9C+wOQOPyfIVODk+FNxOH6K3FrLiwV
ltXAyRNBmcw1IasnioDWJsJdR7uMXxmPx8VDxYhfRlFEGVdd67gA+ZIz1Gy94B15
JisZ7tyI0w8eQh9hT7UZ+w5OZ5Mt9grAQ7dNnJEHtK3WUgYlf2vy0L+q+HLJPw+p
Zc6bNRKvvUISMtl/v7AoB7P2pQrl/iJZI1QAR+5n0VnirDMU5FcuTFyfrZQdN9yn
J6IqTk/owWQiAW0xgbPbsAvQ7+CgB+FVdmyChro0LumGj681X+zjp+HV5cgxuNDT
/LYv3ooP+s2JDrTv0/8Dats5/73VZ3DHMWrqLessfbNgoavmvZmBuK8igHavboy6
Gwv8FDmUd5C+nl8bnXTHRCwZmmSu6i/yETadlkjoQgpKKWOv5Q0xw/A1kU2/XbY1
FNa8aZ+3kOB2/3mP8KfczhKz+Hm/Yi/1UQYsAB8NuLifklkl13s0gEGPLlMepX7+
Fo2YI7NKIwA/+/sViOjucz724ftczyppdGbtl7+HXwdliL7CjDCcg9CDpCmfTbcg
pS7YlJXBtjsneNxAmuYNqJdrc1mmm6bB0Q7PETJ/TQcKqWtMR5k8sP6po9OlJxSk
Gl7GAzNOrMozjU6vf26RWGhr8EkKk+bgVSnk/L8pqpfugmlD/xJtRczJA5shnSEJ
junB2BQt5xOB65jRm6PWOkqxnycbVkyN9FsNcxsXwD4s8LQ6uQeibhd5OKXMumGd
`protect END_PROTECTED
