`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JUAe5edkNYZVn8qkJ7aayZDYf22K84nD5iSNoomWlcVhtln83WgEL0rx6kCmyYr5
QYILRAOpo655Zp33+yGaG9fS2cAMNF5DOKf7tWupV72ivnXQ6PiBq5xK3A6WnDo8
x4h9xMhHKniMPohRGWUdbkWA2zqJThDNyZ6CVlO/FSWoIEu+TjgEWT8V07/Zc9DH
4hsDXtOp/0k4APIW8DeGis73nRa5Q0wp1WEo2kPsjnSODE5Lic5T7E6pp8ieMrO8
iWywXEgwzQyxE3zA/ChKlN5HxN3swF8/wUUHBpXO0Su6/HIeyp1N2Ba8PnGVRh/c
VK63HW/XsiWlbvZGajwDEyK9+N7Lyeu6CqoY4mpU71SF6h0MCOGKKURbHqQmZae4
x4IOVsoBRdPVWhWR14Avgx2aLtn+n9Rvp1u2PcSMeGBVPQ2vEOETQWBa1n27Mou6
tqIxboA3kRlQqjbjorkVpFg9XesuW0YhRyrKKci80d58lymUf2Nz3Q+r3nWdar79
0KyunhTHMjJTF36j3Ig8uMuhyhzmVF4olJFfFLszjbt4roMN9W1hHFQYbSUYxaov
o1vQEfYuXFXdfpw1S7ug8g==
`protect END_PROTECTED
