`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RzCKmamVc7wo1A/qRWvCKsXBnuQwzv34myFJkACS3fItiFczWV0DYSmd2RrMRIOt
WtnSnE36NXLX1FuD//0JAP1EKgBtlf7TWJpj5S3UpKQHjvwH8lY9P0n+obm7/MwU
f2KO0TBbPU8EnmGIrdWHtixYDkN242iGAHIzYNuDhe7WU6TdWybXGn9IZE8iRdIB
LDRGT0/OfvywAWSkKvJNT+gwSID8aM4uydxbR/dN2rubaU5ShftZsjvPWrsQAS+c
i1yU5+QTTxlSmk1O6WlO2IBpb0FN37Y8Qdm3otE80QAt0ipN7EU+iqVU+QmrAL7F
SBSN8pCfPXaBlLyRT4fGX+0JVMRaZkHXX93JNq2GJwnmkyWrigMNjXgEu/JSjCTW
Hry6SoDpvxWoiqeJnM+UHd/pTpzs+Dq7wUG14E0M8kHIIxUc6K4+ovfMToAG77Ev
4sOIFdbq8PtGfFNWL7yVcHxQfFBc8M6E6iDc9hmr0Tw=
`protect END_PROTECTED
