`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PqjcqTOXLCOSR2I2g77WrCXXa1HiRwQRtsHJmrRENHOP/DgZt7hIDaCcJEQTWNX5
JfLNOy0Cl2xxTYH0p0/pCgBbrsG3temQF2eNQIA/HEegH4uK2odYClsb7eqQhkov
1MvUjdtmi2+NpzdcrfqLkQKOHlwda2qwqr1WPjIGvLwUZ0w4usw0h8cvHmCtMJ6H
b3AssLiVGi8xWJd4EGhGc/QCBoSFFJ93YeDPcyzQOWU9yy7BGzrlkPSpMdWft3CL
0Z9nEQPj3bWhyqN2LNalb7ItH8m+BlUEYVSDLG2S4LSjuNz1420UklwMALyydG9v
Ivfx8EARZDf35ufSxZj84oKD7u69sARPF36wPWNP9zEvsmJ7qnxK2UizJYV4MMlW
vpIEC/JTxZCogW6FEPWH0oqTXhVZwFrX/peEwf2IpYCracqaBR2UBdga3YicgsGS
U4WXshi0n637S+50b9zQ9oRv5yZxKJlHO7wSRLhUQF42CqP6/Q5zF5JgweIGeZXP
gWWEeEsHyDShs3/I/bM26lJ8e/uE0wdbwf1UiCi1xAoWTt3c8qWc8bhM0sjCDwOh
RbS17GMGNYiwTIyeHAqCVS9wmkqCyyQJGK9+ZE9QlypmbVcwBddBCDQbm5Ai1+lT
5+MohHqFaqLO/eWo9sPRXrHAKz6l8DUUn7cJFarc/hA6TN1OULrS4W5oaxaCLejR
AODISbxnF1xPlIC+pqyAGuYC7x+kgX3Av764+NXlGfrHgmbQTCewduOsBRAuYlkK
QUR7GbxVXosoJ+uwarj/2JN4Q9KQ8wY7h7dtToPqPp7mnfq4ObbJIxplJL+kr4Dz
YTCvwXB3O9FcufJ4bkbmRg==
`protect END_PROTECTED
