`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/jV7RO8Ekd8nHssqqE5C0G+xVFkwlbovZ3kdHzj2bDTBnR41vsdnj5yJaQP1RylP
f1IbrnkEpNFWdbEQdU9dUt2NvCFx2jzZYrEbe38UNyfYi1Ft7FDG3KjvH0/vXM1o
hWE6Jadpk44Dzdc3XwHiyFBdhUDE4EA2AgPTObulLZimXzEqhFc5sBca/BnWWMSh
1OfaV/zNkvCBnKk56an3D+Y/4Y0XlLX10H1vbxf/hMc3MSNch0ddj8mCtj7/0nVl
s8hhfqz+sncuXIOfZc5+y0MYJVqCtR4P0+yPmF1THV+gcQgDgRIYM1gMbcHv0sA4
g9G/9ZwE2Bn55KRyCeBmUanxkRLYvazdUol86CNl3ppypHXWUib3N1bttmaAa79K
tYWiO1N/ws+mxCHnDnMO3Va9zD9XrkeQGUleFEABxN0=
`protect END_PROTECTED
