`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FsrTT8PwgPMDMj/658waH2Pyw/b0z45Le/tISUlVt+e9A0RlFWQYZ6KdYd7eNyDG
7r/yjpsgyqUtZXK5nO9VWW20xs6GQqkFr0FnXdmpNlK8QrsISVz5/YAF9ELD46Z3
yXDyc+Cj8HELUmdAlBOM1aaZ05G84HPp18t1/lAtbWL49xGpTWc1yRzQyA0kcxTy
hNHvV/lp3zlp+eZLMXKDzouv6MdabCygI5v9MdJNrpNC5uuNwebAJjoe732oaK2c
aWQ10lKnNd3jSYNkWKMVTO2xHiiS5HfA15bGEVX6uTi4TfBUbK9gLSLjMkX0xEsw
k3tHvIY/1wxrnmExul/vra8c3yQyDAoysG+LyLQJVTt4MK+rNvybIzmCTqVCjnlF
SrmaXEBIzEZ3b2xbfQpmD3Bc8NlzmAADy7siQL+Rf6/+alrHtiGq6Zqs93fAQNd7
xF/cI3wTdeMRy4975E1sjhfSbb8Pl/dqEtT2kMBTS4s864oHdN5NCPruisQNxM0p
VTZfdCHMMsKOfH3mhJFrhR7e9v/i+/GfX6YI40eQw4jR8BcwC2qGr424vYH+GMwn
x9BgtjcwfKrpamMs6BLN6DRD095V0810xsUmUtfug69+uyccFmV2HnCvDRfZ0Flh
jesyDbQoHauOYI6UG8RwSQ6nE8WcEYU2yhguvbtPDMSSoo4XGAyrEOEs0NQt0ZgV
L5vX+QsMayaC8icZW2xP+IFXx4XG7QgaYHWv7IqkhpIMbuAy+rHD+gp3haswqRsq
lqjWasVOFvqLqGlqbEEd2ZRpmZnF0zFagG4VYv7tPq4TDGa1+zDo3ZwXb+QvamZ9
v/6b3imCIgBu7K0t/PycGb4IibOeeOlXaqAl1LgzDU7c8WIV91TGVgS6gkfV74Za
A7oxDTNxK6qdcvtb7nIyIJf1zIuMtmwMKnzuAddLakNu6OhX79ybhpc2hVYx5sdH
MZZzALVnWjGvl+witIcU6Q==
`protect END_PROTECTED
