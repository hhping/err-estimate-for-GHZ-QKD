`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1N8QV4pyZijrzn4BdezE/rrowg/oD5UPABMzTDH0kEDl8h/QVw7CYM6Qj5RcHKm3
+rWT2LwOnV5TB7ytNcJ2ORJE7iUfg3Q9wItLHGjxj04LJHI7cFwunxfWiInHt1Tk
sxzW1zeJz+H/QgFFVrT1duhlqxjRPusiarNzmZW68qwGLYMu5i/ovu80VOIHYKbI
4T9+CFJX6nn2TXicIUZQ4nK6I8ABzMtlsQc57pBaR5e9VFGtHiEP+3kA4QEaYEdR
fNCDGc4grUkiqDfavhqRmieu11O0qsTzLz7eHy+XLybJMZcyz5SovdlMyRAZBWZI
gYOIvAUp3pZpFiZDOwPOQInwmFu2u8KWAXR7n8/OAP51fW1GkeR6fAOlkjHhkWFh
jCaWeTbAqCRVC4ZrGAJnNCqY1WHFj9+XrGyK1uGAwbHwdz5PAbVICPMW0588ogpX
TeA3uJK/cy8neowBmmi4bzpbgQNCSxyQLDFu+e2cDStBV2RvOR3gnGJAJILBTXDW
iKOdyMcM6huBo/4jL5Bpdn1H2L5FRL9moC/mtzensmj0ZboIj0PERkSWktkoninF
fBDYGBi0wwNK2TUrKMlRvkbUU2Rk1qtHiA8a9+QwwtgQC/Tr/HiTxslBG0zb/XML
FhO84sMp6H0suLdw+RNF8G08LSe0AlOFPH8LUTdronxAqcVQMlUKCSr0s/+bJbE1
0JFy/V7GveRhmVbKbOXkW1aqIUlHDtGqMtbvGWB7LDlcR2qyvj7YqkGythMyQG2o
9y7cm7zZv5LutIfQ8v/e2VHBRWlstAvraj+DR3g2Vl2ErdF0GXybfmf/N6Y11Mno
F9LSWVQbt606s/BN+HB/iNwR+x4aNkqCiwbWZ4fHSf9lG/aErmPprV+G5Ps9juWd
XPWpQtHgOPxLhhy8djTXeiUXHUAS/++WR2MbC4aaiUmD14TGbudVLd7jdA6eoEyc
oFPEa5lkOdPaOy/C4Hx/FM7pCDmZF3C/DXBmDwDSElK7pKNw8Eu+grBIkj7TbW2/
huB9FTMkAHTz47K6nDB1WCKG83NZxrMchCj2UDMHKNShRxwW4TNPWfdis3+PO2hm
HzFZrWzBW1ODWcTArzV0qoE4QAR7vsafEhaJnPz+atMKrRWgQHUnsetSy636pweA
/d7AODxoQ0rhvMqTkoNgVsUGlygtne4isPjd+/dsIB34mV+aFMIPH4bSZQWCa/vi
Pwyx4dp8UISHev+guRFXtVdZBdj1smzRcK62dyQZoiK89CJzDRUODhQpIgcRjcVn
I1Y67O8aF8XhknVp+WcnkxhirS6UKyt9fTTuatwLtsgu5z2mn1cJ7SkZQGc6+4jz
XdOTN+Rn8M0UeGSYvXlXxIH4FnqQ9jnjN0imMTpJ1Hc3lN0XE4Me7E69Z8t+ALCh
w9jPYkN9vEI3modOO5b4t+VYK23nMO/B3uMbvTh0l6pMK7YFeZAF547pxxQ9T12c
sSscZRm5GHawtXvujlPoXyOOTf3RhDVPGZIkz3BWAfImZ28158p5I8MWcttPMPaS
BfONOQm3eTGU9lfLWFosCEUVOJkEEvI5jYQYX/FgEaggYaikMa7cw1tnDqBqCAzp
89AV5HoqLarLHjZgeI/dC2ZSd9sF2NcDjQQnXS3dfHFj+J0PKkngC4DKjwhyFSDW
7xFk+GskAtzzNL+pahIooCM7fmuUNzLbpNh2V1PMgpIqmUMi13JszJP4E7nxnSm0
t2VDQGCarXoXlj+DU3KCHM10l3nXEG7Nv/fm53zNYS/R4cawzaCk4M8qYmr+DAFp
qdBHDGS5SHqlFdVDccxuSa1cf3KG1viWErTr0bBs8z9pegELk0eM5rpjSqDqF1Ks
CmVd+4551xLa+flvRt1mkAbMek1DqFtcPLqll1bTCKb8PtfJfgaV0q+/X3AwvwMg
4Ou0o0kedg63Mj8z/2wOSJ0FysmrFgSF4bkgImVOI2uZycBfzeywyIqPfUvidMHL
su+u4gLQk2tcgV9YX6ehBNLh4EDrnCkKZRZvH+NFJzQd+mLKW4I70hj0thFfyMcy
PtxX84PWmS9fzbBnyCUelIunoLqmchsLcFVmeIg/pF8v6TWyyZtollr3GTBoL/J1
yMld+re5pEc6zq90li1T4Q==
`protect END_PROTECTED
