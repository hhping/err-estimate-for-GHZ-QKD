`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kermIGQywHpVc0G84+zDX+6HZ/sMhj4WlRq64C2QvJWQoYrHolX7a5tNcRGXwYfU
0cn2hNSZPBhv3aDuunUNYiXreiXcEHJf8yyGG1JBXkXlJ7jGoYynnkqsRJ8lC1UU
4pNbcrSZ4jCFNsHAohUP602E/1eVB05mdXb7TLy/9bCRRehS9qVU0YfWd9JRksVc
PAiipkw3ftfXFbt/eL4/NTiujl1Qkykh3/TH6Eucmh964TPU4RuWKCChuODDkM0I
Irm8ojJkMeTM7L9K7RpGDKRKUgnlgn9LN16VOe0CNEftlvnM8kyKcAL24eU0pgWi
1yZMI+q5K9irZnNxahlmhb+q/0EtKfhh5Yj1hekcrAlqZ8BdV5MXTlLoBtWl1Lm9
SAtkZRJBBucQi5oscoCMyTq8fyAhal75k3WriU+NivmYxKdmhukUBKrgxfBc+10p
BZA41T56QunhVjqbVbo7Td73NzDHRKieEbub4snlqkBHHz1BNwDlAqJjIJqK7F90
FXV2SSRJjfFLyOWfNqTCyyfc4cqAsW/yShTqzrrNl9jK2WmYEL+734RBDCRGm8Jv
tJ8ZwF0W5KPXsKBzSuNKpdH0dwF2R/2NYGa2vmRAx1h+sOmNykZlEq8uRdYf7uT8
4zpYRVci02rnIhdPjcKrcquNHRuLzMlAQ8z3wKPdnGTa+DqW2IfvPYQ2tqoFhwNQ
/ANKBrFIHasmtithuOehYLfZCjtuhE+RpIqeotl1HZPBcuWpxLxKF31AM5SMfZVX
oXsoEBz/UNiWDljsCGeNEaWQmjXK5hBXdeBEd6JHRiEk0XMsWb9Te7aQyailDju8
Jnpcc7yVuN5EytTLYw214Ww4UKpuZEMS8AZx+yv/yTflCo8LJrLskea+w2kcxE8T
mf4pBtVRfCbs8wRaWCyC3QXoo3qPIkG45R5S8rwq3VneNj44++h/9GCPBV5wUQX3
J0o7i1mKgLVD/HVg7EAGdw3bQF6ppi9kc32QMaoezACitGmkdNtm7zMowZfeoNVD
TxCx7rtvre+0Uhnm15Xnv5CRESVVgVpkU4YsIm3O851gd/t/j5uHDwNUNqqQA7wF
eq/MhkqwWC9ZJmn/NnapRFgk5G/H/CbpYWUFw9uhXFdXkeiXLP57qoFgz9gBsqdZ
dUOjX4eQuP69mDnrJQAux17QtJsB4Inm8Cp2491Zjx9RFf2pGMWnmHHypvynVjTp
8IKPC0EJBQqIun0YsWoCvyExcQgTeEuI5DMoimGCtAddckWd3gsZysBQfwQ49NQn
4fK9+8495+cKEc6SxpZ3W+mecUi3+IP8oA5FRTeyBWCOjQQz4hIMxVPkq+AE+ui8
ro2wYDVdGBjwVTp5TG2FIrRWU2yoNhdlnThwYjY+Tbp73aKeVvT6HSm9pivIiZ0C
Js31V9bufQI8aFy/YKuZfx+PUexpdiDaVmXAe7OHysa1g7H+MV/7LPZSkN1QOJAm
iDnc5hfrgkrGvl7oEIn5xYO3dWHTcf6HKideB/lCW7yi7oMlPW2Vk2sJuQ/gJqmZ
boh+9qJ9Xb1uglXw3q91SMihTDxkPE9YorntXCo5FpM9XOTWkHyjWHqZgGm7MCGC
VIUov5Rpic9pLDLO2q9Hod2dU1dzdlbg8yBAM9CQQzXQNN6ES48rUBjxu2wyJ4gV
OOpgHvZVZPnMbbrUk84c/bF94eGRIoyxaHW84IXfxHVOkVK6rUpF8TECrwMF0Z8a
BBlL12rYMKNWoki0UZo5fZsKIX8xeQVSVHnliZ1rlYX1uDBC4paXBsTKndSZQ6Iy
MuAMbj7X1GbprUvicPiji0h3/vCbByHQckCjcEvCilZqTfbwzKn22EhKgBZiR5pr
xi2I5n1PEjtNSCOVHAfLkxicnfcTiTzD/gS8QonnODWTaJt13vWHfVhtxHVEg3+U
QutV81QPgjVSASEYN3w6r+4oYcraRSKs+lA6z2zTse4M1BAJMVrAlM57pCACtHja
BoT20qSZr3UAaBUWs4WvF2UKvnEk4yY2UWm2ubJ3TlUKKYw32nCXVp03X3Swe0Iw
1x4QLrgsfERyX8SES52OX02XT95gTBd9iBFkZnKWtgBZJAwkvC6CKquXAC9N1Qqz
EEIjklCJPSMp/VWGUKR5406UpBtY3AVNV3Dpuare9VgVMDbXOIJ088hmf4Wv0cQw
47bCLDzC9nmaM6tI8V6I0s3Mju78clnzd9JuEF9gCn7HvIeRkoywoL7keZqtvfyA
9M6tlS36LjvECxToKnXgmkTUe47pJ3DbdCxf/QWYV5OxOZU3yafHtGvzFonhtIOK
Fw6VR1uHWEsFML+13WXx7Y71qULJGcILHdYZ2xwOMPGZ6bcqEV56CbFvwWh6v4Kx
JxillcqQrsiu8jhSRhCoQFJ33EuuTTqzffPxG2kb6wyIfqloP1dF8C6QmmZJ31Jb
W2t77VL7o/tgk6eHvgyEPA8S8nk9c2/a7SImJU6x9a1QtuFi6vGz3aJQc3JR4XYZ
yyNTOU+9jg220XQxRQH+iuiyzjFphUU1czeV/UxAA6n+yPCUYnPPiIhtwagbPpbq
Z5C90t9OCQ0UWlni62o+kok3dHcgieZaCdQdLaZQn+pGA9mugNXliForpDB+3Ulx
BwZ+nL1arzHcgT5j3KYUG47/Rrf+82cWYrWXMk4xM1mViGq99G30MpwHbS7N5exh
bitWivta8oGjrg/Ifl2S4i/VldG11Fjg9sTlIaldkRtLVNcr8ZP5bnJvyMd5BLbz
omW248KT9D8gP4WhOWwq4XqObGI8FcsEQZy0bn3R8t4Jio0ZmC+Sqp5uQg1aP7W2
4A8DzxKiGFqJrHdekYBI1KymEzRnSSz5H3MGlPR/IXs=
`protect END_PROTECTED
