`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3rUTK5cWTEtIF5gqDfjQJQbrwB0jXQGXvM4vHb4FsIgShhegKFO0+FuEnUtGh+yT
nYX3mQiJybVx5qLaQAhVNQWPi94TB7BbOOWkzfkR7MtYypq8rR0mrBAQ+H7hRBDJ
b46UNKfx5due3jf7DVDNPMU3DpXEaP1W7JChcwD8KOuJ6iCj5ok5AqiF1qCdLAO1
VjBKhld0bEnVhd36t7WyT84lEyshd+e8mZxvAKRVe/KCw15AMBUX3oN/Kkf53pF2
Mns4FnGIXra50Nsbba2H6idQljJns36uHTkkGnErPUYKKUOpGCiF1S09lbQsVXNd
M9Mg2HCmPqF16ELiqgH0evIk4bHd3aYxc/kUix/vtZI=
`protect END_PROTECTED
