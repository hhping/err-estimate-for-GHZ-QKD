`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rJfSaoali3/OoIwRBxuYtrC4oCW+jnmbUVZI3lTV6e7K0gYloFRxgdklCGy+QblE
gcEESO6VQVefr2qFWbF9DV+2xlu+H7WHuaSC5b2NAEM5tpE5Q++46WqvJ8v0KL/k
pNR/Wz2KXFRoO0ov7CRcBilWWdYHfKnnWJN18TiBfExwIkdhkyn4zNL/JhuXJY5R
Qp6L0xrve4zjZQsPv6KQXLVh5UqgPTHVhAaiAx7+9KROT9DdlRO4YouLzvNn+iNH
QxY34Tkw2lKfi1MGPEpwpK5LbhFmiwVZN7zowLM6ak50Eq6wNQXhRP1shO/lmdsX
ZqDJqUXDlYUPo70oLkA4YTlmtcmr5YQDCEyYJhtk/fSI9a10FKhW47uxveBHzwmF
+PjVuuvUzGcI/OY5MyFOvJDmvMIq0fJjg/LTIFm22yZwjdNFo43Au8pmbE25XrIi
aVTwStx8rzxg9+TNfDxVTN9fOxwjVATHV6iyG4bIT+iSTd94BjTd1UfYz0UZer5d
RIiAJPCHu6defqG4PR3Co1U14XHMrsLsTHgEANvCSef/U4ru4XtXUtt5BjoSsCdA
7kWedK6JUUEBmq7f29IwGoi/RNBYf8yNo3Ny4w7ga72RPVq1Oo7ShJak0Dhx58TQ
olD9h1GcV1e1U2MsuQerti+QKzkbJeJ1iTaUKJzq/a+5rpKpxa/dSNXVRuRdaFol
t7EgDkFSvQ8bf8M3BydkL6O1GfM+xz/E2SF4zb14Ii8VFTm+4YDL5fUlKmvJAVBA
dB0Cfy61CHXMc4wzCI4JM4pKKSV2xP503onaJxmarp5nHwj/57wkvNttEGB2vSdf
fKyVSCdvUs+ZkWN5wLl/FMwxQ65VBlIqv/zQw95WcV/xKlQPh07eGmPWVT6pfVSD
BZDJcUm51Lh6I4vvKUN7dElYtnoOZr2DYTtj1OALMcnxOVMbSkKOrBdv4kVttIqM
WmNdl12qmDhHyUWXst+6W9nytfP7P+XeOns5U1M4/EfvtWBvcQ+q7WftVr8sIujq
PPjPQX6DJEEGqCUHRVwnG7crCI2idHqGjJvePaqxf/5EbP5IHnaZ6Qt9XCJAFnFr
9UQM/4wFWBAvXsKduFOgBS20WMVPWYhEzfcsohIRSrivSep42dBXnLjzIOTsVozy
6ncV5jshpf3X5lru+Is1k/8ZGCC6+WplLRNctrRPv/+FQ43tEToYxA2gDkntop0y
N1UsrZXY+qB+Rv1gxiEPdBjtcjTTSp6Y0dxAI6/6d3afb31oxS7cekhdTH96YgCx
cDSX6VzJmOaiC4XBF12OC1iesysNxovywZiwcQ/R4DE7zj39iOOcKBsYGX1ubguO
U60mnEFylqYWlKZTdVPXHO2nzSvHtj9kN7JDVbnLP7Dg14yGDMEo16qqTQpShXo+
xlEObMZVgq1V2+sdPgHOxVMX/PBSqdQSUzQbZdlTkVKVmpf5ZOu4mU8CPbzpYbyR
h5ttNNfPBbtzDAKChyiSLQ==
`protect END_PROTECTED
