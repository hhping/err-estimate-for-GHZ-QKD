`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bgNGEdPbNJMGNb+wH/pRfjyee7bj/DpD28nF0YXvJMXK0y5Q9P9POQ8AFq7LwfVs
Rr/kC1SOaxSFsU9/KGPTsegL3F9ZiTFI+nBPT7kFBYc/73M90N0RTACGBe0eKZoh
1FHhwmX1Va2mT+Nhqo+UU/vsX5oIt6xHMLJoreyQgKpkS4HLpkMEfhsbHX7wHhK6
/m1LQe6jlbPI5HsMOq8PpkjqT586ioa2u884rxDUTfrAa32ywbWkvy9QgykWzZxd
6rEGZw1Z131QeyFfdySEdkshDwosDfTwsNFTqaSKuOzMwX15zHhlnOGG17ees2MZ
rw1x1bYH/061Ave68n39F5OnIQ2QAT7zqKRTLGVCE17Ki443H2nepMhVoQ8DjJbE
/2ftMLX8kbsaqh3Px7TsTcgyk0RLmWpRi0D/8Wd/4STYEgiSmgybv8/ZW9LmCGHd
1VH6av2TVkmHk9+iypv75+Mp7CT8SIOzv1bwRNShFDNiXkB/2oYA0CbJzY49WpXN
3XCctGHTBa154NFG+sFgguF7DrTEd23VhNLGv0hGCCACd7yoGWC1wSX9sWBrU4I3
vAgql0GTLRPfxFEPaVkqmkUtbvMlbDumzqE0dLL9trYVJeGJ+5ibKlP/7ivpGu/4
tJkY1uDJ/6xCFvxBvOWZlwQqG955/YqPpgah3KgDwzhzlE6Q0LEK7jkRBBKAehi2
yOIj5mbM5oJoHSNmqJ9cLz07ylPJQ9zCV3AVq51D137QWMB5unrfQbemGVtW7WJK
T6uO7PfRfh9FW3Sc2LyOfpMdVd+CinrTUCtnKTPjIDphY20ItE2Y8YE44Uyve4rE
9P0E6xyh/L5GATQXsrPHgAceFtqbxmtTs6NwkSX+61X+gFjHQVxHYWOIUAdXjDYS
6ouwLHQSIkfHZXfNIYv2NfW4OP0bDoHCg+eLXAer/z/JmtBnL/rKGnGytqmUhuaN
OzS4Kiw2hd0fDuWg4ckegNGe3rvUtH03ileY4TMQKTEd9RE38mXOkcrBCBwHpVT0
CGT28VNpuGP6xKqnzZAYBj9GSGwe4ME2PFSgIZgcreFYz4Vgq6UX/cGm6Iz6EI+i
kAMkebB8IcvCtESVrIojKDDlWsp0baRXt50HgDiGOQEtP/w2hnHo649ROXjTC4Om
cMRm3M197K2cs0+jv7qX+eSp2sbfzsgd+j+m+ShdiC+ZjmJBYEJk9xK4djF/nMfc
melScRR+nlzCIvygfMuLJrr6uWnPLWom2UH/38HbnqkImDiXdOOLOyLZSklIfqfZ
HYu10dWmb0lbr/pOovYTnw==
`protect END_PROTECTED
