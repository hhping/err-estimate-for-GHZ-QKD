`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2gWpZcRpIZbMgfVGQ9pgfWLiaDx3+kV0lLH/cIpqAtAUEacKt+gHKfVx0eju439/
SKpMYUIwf9D6PHbvwDSuplVAI7GprUKP6fgcd1BDXEfgiMvmYpfX+2D9Z+pq10iL
b7+bptsTRUmgnjPK2YQ+otDkoiTp0eKy4cLSe9mO62856in2FsalcCxDNPImsjM8
o5uuXN4uRi/yK+KA+Ujs8AZKnQeFX3yoTRoXb4E70kkleRj0usXMGLFcFB7C+8TM
CDdJo2JEDL26P1x2QpvzTtRVJIcl+Y+BIjfWOxcZg3A=
`protect END_PROTECTED
