`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fGwsY8PkQXwNUmmUyAh8g/wTMlZUjU04OUJv32IMHlpEeUr6QaOsFXsiHl/NgCRt
GNqjy+HWSptJpLN1iNY0q6Zh3JCPb0LoynwJKqQtzC+Oraas1fhjrIRE1gq5w1cL
l8OmLhGgEhqcbkb5As33nUrEITJfhRlTwT00HUfpzRnvGO3PqtCOgGUBdQ/eIHFI
gHLfF1dZz0RH7jhdzyXPVKWM7qo/nQjYI7bXBMsMuGG5XvYXB4Wazp7iPd+dT5kK
3RNfpGu+LSvh47KQX04jqZIRFDKZsov61EOprx7ZLqROMwJQixwqRK95BzqkWIrx
BUmliu/YI+DuW2qspZrhXEHy0f5io5ZwiCsvwWnwA2EuykEWV2r9CL+vnp8Ww3rU
6QFCRj7xfURSR2olMHNOww==
`protect END_PROTECTED
