`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vdnca+Z5pnE+x9tpk7M2J+upPyvsFjfnRBmLEsNYVJgbm1zG3+36RK5SptlwBOlU
uInJwWUPEIJsSvsblVYZnPEwZcWpKUo3HaYnvpoVel9YXYfAKUTsX1Gsxu7heHNx
OPezMo8l5I3R+ff1VLwEL5ODXIV+DZproJO/+RqeKgZK5PA2iuwCMnbJS0oEqIDW
WVespFLx2QKcc1insK5lE/Tp0OpT+F3HNG+Z28VTuZP5ny1WqWYzKkvPyE88Y+2m
2FCwWphqGnATLz1D5bNRp7tBYsBXy5mpFhnxkgpLbZFePmxnvGCwY/6SqfQr7zz/
gIqNQgzgio0NMS0LE5+PlJgVQHqWOZRO8wR/JZswK5hp7ITjZSjtuZtFwwTvzUVG
XQ/7KalChgNZdwvgdQC1v5CpXKNOkG7d5YoAjNehh6e5qG6YIDfPZGb6VFxlDN1Q
K2sEVCdfYu9fXXIlqQzfqBapGK1LDwntp+9bbtOwd7iq857O1uOh/BPVRCNH6jeo
OyNuHa0yf1o+v1Lb96HyszWSFulZdLkQXDpjxwrv3PrUWiJBzI4+bn7Q48tk646G
IPGgeprx7WmEpeqXdrniTcFsdSdBPHQz/IHrjzmiQoFycA+YlyhLsMpPOCSU+/Iv
0dXllCF8Gwiytuu1QCsdIkAaNepFX4ShA8TFDnWjwBLHQ21ZtQiq24Ydydl9rL/q
0/W5fe8lW6IOwAlCT5fJ5+v0JC7FRM9VAxzMrrgfG7I=
`protect END_PROTECTED
