`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Omd5VQFTpXYgrP0Evc7XoFP+3Hn1wd0qJ//7hwtf9vFUf/PUTJp1viHeOyWyHJbL
VPb+kz8ZEFhaIa1rFibHx5A+Y7uFXWP+kjiycRLYJmiWG2Ty1+2zqRqSn83hFl9L
Dd2UMqC993g2/1hAua9EcH2szmDuVG5UtrzM65ut9IsAQ1KQA2qE27cwcxKg+N2W
hQspT0T927vXhIyr8F47G8gXod2UdEco1DmxVP3oOijebL3dOuMSBtq3Yjqj09/S
AoCBkk5Coqi5g3UzC/h9NN5wvYX6ppXin3qucy0DbzxpOmO/IZK+zFsIYziIY/Va
KXhyEcodE1kmu+g/y6c9gFJ8Kq5hWzvMQLYWLqpq1r11Y0uzTDpdQl5mt1W0fbWm
RaRIHpIT9OpOcVlmTWlf2qHtgSk7JqxGvCDQQka0hUwI0w3FNnPiWndn4PmC03kH
jMTkidJExT0DWLMU3Q5n3RSt5Nm8OG9BhDiuUU3qFmKQ8o5MSosY7Hp7WNS7VKwv
S6dA2A24fvQtrWJrcUE1AhbKoasqXptsHU6BB8L+KaV5OKnm5iE+RIHtURRCTZEf
LxuR6poWmR1bG0Tm5mKa8Rrnia7yqBzu85s3oKd8DOcqHG0bVkeuxAkHHswM9AGr
BwoWYhSKNf4emjY2dP8mSw==
`protect END_PROTECTED
