`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UIVZKJ2tuMXh/ihFmhPmMudYSBRGfTZy7C5usswxW06suEvUaNrDnQ670QvYXovA
GGPfXYtEDJfp1A79H0jEPCdWSlk/lKguIua99bTMH/thLKcWf4G2YiD+XjbNnBCm
3zPHcXonNqIQE3okhl5DyNguDcopox4Em4y9FkwbmMEQlG8rc977PokxeP7t1irw
ZJ25X+r5RKXes295SgXr1nRLWSc3hGkz5dFskOITGgoZRZQvOshUF2h2DnSPHV0B
RTro7w1CyXunM+slouTFGN6LPFNyl1hQJ+q6dLLgjxlLHHb9JYXfktd8M5NuxOLU
bIGaeffBqbtROFWFhiwObSnmCnPALsBPhYnvZNlkZ3/cbsHHcM8j52oRAV+m0L0R
R0HyW+fS8NrEUhz8I1rkGbR9XsnTF5YbIS0rTiOC0VKZgamIRDDtujk/zrosIZm5
wqtP2TVmH4q6JGrwRiHWMBHvLtm4iB+314ZDS4iAwrvG+vpCNfqkrctNx2R2SAB6
XJGxBSaLgFc2LIBhf50+qdQOqp/wTYsvrZBGKAgKVOewLdBEBbRkCAu+YWa+s2/4
kgzb1WXjQqBo5259JCmdJg==
`protect END_PROTECTED
