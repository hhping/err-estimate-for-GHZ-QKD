`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oa3K2A0NHn5PdK7a2T4DZTd8wvHflAuUAiteDTLLRFKE9aYZO7lDpqAFJNQZGcLa
U+Xc3Lm3cZV6yg9M3xvz/m4PZ6WrEf68M7ESJv66sR37XXI93uj7kQET8xldBpLX
2iGlQEfT9O7HyhpCCn+UEcV7Stsiou1/9YjsEWevknOLE6IlcapMqe0pYwAtoFfs
tVDELnauVco0IdyVYCnkZ7ZLMsrEvx3bep9I2FbCw1xwPI6tC47AyiC0DmWuHIij
EHwWgKv6nlA5YkRQVbEewMl7gb0K2UgJSzfAUdckaskUEYSBDCSc8UkB75emSH85
zHCBcabntjHset8UFxeroJWIUlGikqDyHG8qIG0EoIr1ajQwOixQ/LN8FnbbgTiF
vXBFY0nitALW9Mf4OE7gW1D2LbvesBra4EE6ixA6pxA0+BcG4NE5FTINVXWSxUKC
539l3zXmzn7ZGLoHzVhP+UzeaQTW/nE6nFyljtKUGWIa3xfU3uKtwXrabEq9zzdy
SxyardSIRYCd/1k0dWw/zL2uOqMVl5aqZ7b7oPLAolYKP7EkohzFKd/iDzhzO2+U
itlQdWvK5t6JpijSX0GZPqVRwOLZ6Vy6XRV+S4ChO1cI/goimDeGa8JSJuUjINol
hy0HUK1wO48Jiq2rNJX0tojQVEIQW3Njd3K/Jqovk506XpJBptIUTp58IQM0oYCa
zHoYGdB00bIURIvCw77U+6s9K68OOgoV3e5eYjUSff2ZohgC4Lr/jyQfPOfJgTqc
bdlrRg03ip7KoFxiim3EB1d7vhHqiAokrz1uJGw71BUj5cel0YzcBq3GJX+C8/pQ
uBRJVgZZtkjTwGZZ6hyhQa75+7T82pUe8XuJBW5tlIXip0aYUJ4DZgO7l6x26kAP
uHJiJEcYYJW20MP4/5S/dC6yAQdR0sMB7mH+mNw9mAkNx3+4iDVrE65aH6/BRPgm
+gbDuqOE1Ma2rM0iCgv1nm2zNwiwi1OG9dCqyeqXYFnQcH/SB14CpplXl/5uUc/6
osPafftJrCCthINCUGUbwRpeRJIuEwAzaq+YNc6Kpfp3iHwbngK+VbjYBBsCa2bj
Kk7J8Sra+FoGq+NLrZksrIrs/RduB9uuNcSHnt5cM1feIiEeYmeV3TnYfCjl9CZv
JUv5qBcr44ephbewzik0QUfPKolNqSAxit/nLSYUz9dcdjA7vrHvi007vLGwNUmF
`protect END_PROTECTED
