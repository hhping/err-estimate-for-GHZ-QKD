`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i1I1fDnc67H4jcbLGOL1+429aZs2dxdU88ueg+CNsTKOd+KxaHQ19Yy8uAr0i49Q
brApcZhLwA0kwRvh1VqtNmxyAJin0oTBy/HzwswHkBSQAsO/Ph8c4qX+VdBDd+be
Cr5TJiWP+4WdPUeU4cTctMFIQOwTDfOTOTENW+k+w9v66oN9y9tVGfmEj8idyKgi
Kk3Hm8IY+ngpxegTHShT9O9eicUoFEPnk8AYpAoMm0gXeEapEQQ2h745fGkY0VWo
wjE4HB/IfvdKRvO6PpJSr71JyiYHOw3V4Hz4oTqLjFSc7QGpsq69lteAdhELqO4w
2i4233upVB0KzXJsvalWxVqyNjpMWebyyqkh2bxow/UYdYBQpTveYpeAYQDac0l0
qDYDH/QqCPQ8vLcu1vszqBpbG3ZJkudcUCgjXy9E20Ja/rPtYqqOIKJU/9ZTUvBN
ElksNzvh3n/2xWJR7YNM3AA34T721PYGMINuAWkZJ832nrEMEQBTKE90H17Vu2xi
VRcZ8bgRmkKJbWrTsn6FgnkgJkY0YWtpNEafEkbNeuUiL3usqQMYeq3JyW5L/Axj
3ljLPjZS9JQNPlMV9fkkjVRi7XdW91Iku+XWLpWikO8gcj8UZCVeTQkmb4xd2z6J
LytaqdiEORu45fvK/libz7zCNz6QwfIwDGZO8ciJpvjLsASgIi8jPv4NbfxXIPg+
2hqdtx3Kd7yLagyb3Kr+ZAo8phRczYIiSz/lbkoGolhu/LVU2xXM7sfWI9KIdng+
21zoS44jVnpqwStbQtfCL6T5zWXHdM+RV5Zt+h3irKTg1dBx+thl4jxfNgfrh74v
J4w/PgobXBY1um81QWC3AW8PRf9JLwdfMBnjCg8TyOh5DgusGkqvMTEnOvF9+e0F
N+PlTeQY1uhz+mXp5vP8yvjh3KQHnqn4Kg7+v4ZsuIjzxFm7UZ/I9X43hn5tyrLI
vpx+/0JOB/GMqIUupzaO6fgZnVsl55DjUzVkD4pXFD9TNLR4gyZQCDVHTRq6N2an
e8LkxQxfljf5tf9Ox3PtUrwhJ4iql+2qpzHUUJyW+upghLBMp2hdB5FSQlm4Li8k
D0U08rXRBudwbsZ5wRtj7w21iQW4bOTSWLOax2zXH98rbhN1nB2rGzppruN6gadM
7a8jKqbX5mE2WMk9TvjjiQasJ19WCQuDFbrIqM1sM4kHI9ugEsMXQbSewsfGBwAn
ZKieMAgguvhBzYN2Pn/GxyS00T2dwYz2YF9aLaRGKrl8Bbfh1qJrk5RBNZ6a61GN
eQ+Rtl37ZoALWkU0EDWuY9G1AQrNF+dwK+0NvTZbrxcDyzGn5eif1Ss4xJOmUCHy
`protect END_PROTECTED
