`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jzZ8tErNxVYRpuWJwVC68X9sPs6DDIFT1EDQD0Aray08ld7O/fQsS6UGzSEbe0JK
FZ5hVH3QlrmtTHYvC0mZCWo0AJk+N1iSjm83YNSD4m8esvDZ7A4NSx9s1+oGab8D
/XuCaHwnJ4q/lFrTaXKh6ndKu+0K8IKpeac8Begeb51Ed61PhviybD04nxHmMK7P
CZT2wW7arhrFMfyVLsFUkgbnK5KiXaMJIu5LSrDZ9CWJuUj911Zl1pV7pqa+6uIh
qwmmi6MzwjmYWXd/HoLzIs/p5wPeGUE0Cl8isDrFXDrDw8wxMq7ALKGFH/OlCqRj
UAOg9ZJ+4wBW0W1PCIEv128h+ii8CFtkVVJ2QZcx5LY+2kw7Q1lWPul5E5787PkQ
3VOsIpL0CBnxJiZkX+bW18gr8ciL/hUSgDBKu9/68N+z2QxGby1gdNbEYrb5VjdK
A9I9Y8KKkpNVqE1tLkcTM//rvdEz9F39tM0ddt9VEsTTZaOdPojH9+zz9NFI6flX
L0N6mij1mSboGZZqmfnn8OCD/dtoRmSsoL61yMzmdFe9KioZt6U5Ot7bwVDddjC7
UpiuhQPW7j+b3aUR6pc5v5kNcPjMlukK1y4Opin7V/j38C+N8nipjmwRY3lYMinr
hNvc91RfFWr+OrntYujKdDssojnF1+bHPhY4EQsA3oA03XNbWdHJyM61fbJ+I3TD
YCkcrnK7hh2ditUv64DcG9gPJAaWHZBuoA4clG3x09SyHFl/pUx2+awmmrXUnEYS
oP37Fbx99UDwsPNBSoDTdG2b4sWiiu/0APzaPJXirb+mcXiDQ1NpFU376/X53C9Q
RmWVC8qcR6XnyP7zRXaFttTsmCn8EdQDkBWqeK/xXVSVLbLjDRL+rg+LeUHQWb6R
631u2Y1Zyt4VvblbtoCimWEiY0Tm0SVz8Jxd7lzUVLZX4M+ITXC0e24ooJ5zC1Xy
EUktcPKcpPAvrP4kHtpnKL9jInojdrf/hBrzOaFyVsk1dRcDSFRSvJOHIhmZm7AM
5kvQ991TqG8vQwhS5aIDSbUJCntnvBhYEd6jHnAKAkSYexnSvs1HoBVB+DBORBUI
Kwjl5SoibZ3hMB6YVbB7u4skJZW4VvAX1aM20X0Eg/jYY8U62vb0DDTtJhvm5vMl
sQYpDiGJBF7VacxjXlYm93VIqVpEpInFDzoDCBisyR/PCsuuGiIHmZs1KdtId1FV
RJ52uVYlicnkpcHpM982ynG5HiopPvsFd+epp1xvmVng+k7YlPdpI+Lj/xjD9iVJ
Gm0372PyMIwSbvZ9BWwTsnblOpNoLylVPw6HVLuJaIjq7/aNVrrMtmovlUY+9nwT
1a2v+bkJ4enlV7RNaEJhWd43XJVOKThmSrkjWnPQk6VU+2MFaxNzJLGMI7idkMzD
0+sgmSr2008I4hZQqg/d/4ZZXnHOO0SP8wzx49vCft/ScJXcT31TalaROjfAW5Ns
urEuA3PL0LiEi2csjNf4S7BacW6Ge3IOVGOkxTHKmnAfQNG21QStcpB9+2XT2jDj
8R/Nq9Zt/mSmD9k05GtX/gSmKxY90qq0AiFiq7LxoBtN7gbckFRSJl/tjniZAQbS
kwKbbL70nXfd2cw9A3OV+lKelnxl1qTf9xlVOOM1RSXA20GRiFqXU8/xd9VW293P
luHEnw4zHVFBeZ4AqcFapuhZaZe7zUaRQoS9OvP+8JcrVNR7CqVJWO8h0R4pofCc
YcZiHa4w0pXEs76M4x3qu9bCD1kKlhPUEEwTgOw+rzVarTfEqwx454BIIpAlMww1
1O0bvLeIdBrf4GtORsFilr67YkoOudWJ35g5QMaf4BA7N8+8mYdR8VaK8cVwLwFV
QBCYXLRGbinmxsbuJJ+UPSwDs7+Fc1i0oIqXDjRyN18yJZMZKk+3Hnm3blIm975G
1C3E9+FIUkpcWauBwvlzHhagz6a3yQc3zbBGO/u69/fbuoq1fwCV4WfXgqugXNi4
eRRAxpuKUnxuE2Xq7Eq1hBtKDEruYOd1tkWwxP80+HLHhMavCtkJt23rdmDmg8MV
8sxj87uUpfeabZDuaIBDLifvce0h5VyJwYjOp/UynI9jzxEXVGlLdR8uAnParN6z
1RFS/QZpPd+AwjlcTZtA/amlxihNY3O4JAoJCp+6vA2Segnn/mQtrfihplX6jmNH
lN15Pwq4TUB1sZ09fAtu3jjiYbQLVH0sbRmvhjsHccdqHDH5zY8DXG4fM24GPWsi
VnGO81ikJ855GSN46QlfMUxEjo2yjeqvyXPx5xobCHzW5KW3Pb5HZRMAqI+CTD5E
GLz5zN1DuVPYxs9TAGZDeUnwL54fHOa254tiTHCuuYMmwVxS8QUV0uz+pUQG0KDh
`protect END_PROTECTED
