`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jd+ui+eC0/YDcFgAHDQeO7HvdvLGWs/okgll9HnXGa2vld0bdyjWDKR3i84XVqqe
VJTwizX9aC/hp4mOGNppeu3iWu4RTrxGUOGm1+S1tKvlfeGvscW0PHRWpuADltkT
abZ2VaX25hTX+X1npmrvz4hFYXiXpGYd9tQ6fCrVv/yRemMjdYjiL1qN5ddbTsUb
ucvAiOtf22duDX6unt0YNX3oJv/mo6CbKtJwCiVUXeakjoCSP8lHmbwhEDilKCNi
qsBbPnL6m9r/Z1WzXMtzhUNtvwU8tdS4xbOBqPC9RAGSnRa19Gg678vIMEEjxoP0
LneFIj4mco3dwmVlrnKjqYhW5icpkin0IMeBe5WOLKv3XbnftRdlNhYT5Ss0HQ56
txyfE3dIXgy+aHWcY3iSS9qpBjf5EPWchrx9+BVaP4CXfsQymznNkWMzfwPLsIEk
fIEk0tJcIIRUUgqzrG7hB1XTI0TOGd3o8y853PZ5swvT81eCLpHt4pKAzhb5WUiB
Sbi5njEniSUMZPp3SF2nYKEAJtveELB/pKihvsV621muSFxPvg9uc5972BkGYlvM
JDWZBmI2lrsu+qI+tsbgAEr0ANzSJdJ2J2onIgXq8zBvVZE+y9ub4fQdXlbidW5X
JP3QWcbKauXqwY4ygzVQ07XCF3n+7m/G+zEGE1CvV+V91YYzs5ce9EleN/w4MpAG
/X2NwnH0NCzj7x/lyGMPI7l46mjETWbsq0Vuau1hqGE=
`protect END_PROTECTED
