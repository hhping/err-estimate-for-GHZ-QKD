`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3uq/KdlJbIaqf0G8Hz9aD16HNFdfdiNRjUGkYw5Qzns3L+XZa7VsMECJ0U1ZUl0+
EoZpB55sGAadEcBiIEXgdkGr/6J6WKoffSxN92EcrnQDAKYe8xxvKYz5VyEk6Uxp
HQSrkhKgm+tvAUHTSOsEnfrkh3RB/qeerh71q6gzMXoWT+lJStc5nQMLZNTxNECb
gROec84STKop4AcqfmtYVCSWtJw1SjdxSEdZ2hXBQaBVR4+KGywkFkSEeMzW4BMb
hjn8VWREohE/tn/mpruerWMarluEshWuO3YDMFVFXJ7nj3NgnyWzsHXa2AddPhKX
V8+bhXG7mbRBihT2i18IvTkVQ/26ULl6nkM1Ms7W8XBX4WC5OQh6lX+bpx/dsNA7
6wPUsn5A3iwWkhVh/f+mlnMUkbUXnsbtTlUinnOjm2HRLarufPoubfE8a6Nht2GM
KbLhicy/n3tYAp8tapSM7zYlwv3nudS4X0BXsWvtAT6OItduwSgw4ZYV0ufNlMZj
rVjXQQ8jmRuaq1gUv+lEo37yNHn3L6q6kque9jtjl4nBjKgks5nA2mlNPmFrll0D
/cCq4pDTl0DRsmYCTSzPM4wNI3Zx2AF0XNIFYChCDKB7cf7I81n302Ih+DhBaEhR
7CQyYZO7hmHJs8wXxtBWYeomDRVB/CS0fm5u8zOOCCPndDJNbb79G3LTQ054U1vX
Dxbd9rM7v2TE7J3ZGof9cQNgHDQ+PnkziCR2aYoX2BKd7BLxdnu/ogrvVYCrqWsp
mIK+huVMxe/r2xHA81W8y/V+8Db83tdLApmTcNAS0Bbfjmu6wbBrg97I7grZfSZP
maMSzFxa7liyyscev+oq62FGdp9OHfjYyJ1BK6V1NE9ttYMQMi85cKAAFtuPhN7R
1A849Jditeze4OEFHW1SPiHUKYeHU3A+AVE5fHG7Eyk9BAGywzc2xVh5xeUkgCfe
DB1foVpwGdC4foYc/Rlw7xaKVu40MN7cm0g98VSZxSKDqizNa2edFO6AvfP1iyNj
tgLjIBA1bFUTDkWy9H5b/6Wq/DFzbj53Bv3cBHiMbUj1ljOIHZupr2anhjRN4Gs9
vtGXKIn3FuBNXNhnhbouh6ZYt1BtfPPWe4mHll0guT/1h/jQZs9YMqD/08ahB+cK
rz27C447ovNd5U9pIS+q9hwZ00moDlqMsNuOvfKyrB1WibjE9Y7CbretNChIiQEe
j0XAboneQFKfI6eHF5nUc1EEtwo77Dd1rPBRF0PwcFy/lNubEQUfJbBeJzARTreQ
+DDwJaoEQPqooGHVrplBuW8d5A1e2dKZ9/TG+Pp6ESZEvHddyUwEPlLv4fZxrlr2
ARSHOHrYxGnD6iBs9qbl+21fdqT8QwbbuamkURW86x9ZojAAzeLndW8SKW75PJDq
rAqOnNpeIDoRQE4XN7E4NYYoGAo+TQgJCgSVMH2ZJyrs2bz8hw30E/fwCZQkU/Rd
L6akd56Co3YA/ts9Ypqmd+Dp5vIE8DIHbJ9aM5SJyDsPyD1M9A2d3Arw70os6pm7
tZfwoaYLclQYNET2YmLahPGvTjxWWuuBZbhfnPtFExKXp8KqFPjSxGGtVTf6fydh
iVQBc/xYmIvYEUAADvbUSxRIfcMJ3/s+EJm1XN8bsgwoMB/hCdvhUKJwOIrQYJ5W
W1zidcTQYcdDbcQgjK397QJA2NQMUbS1WI16s/6dL8o21PZhYeYEXnl8FUSLivzj
1sAMDVOJoMLgtMO0WxcKqw==
`protect END_PROTECTED
