`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UoZc4sNaebcD13pMyjAtAs6toZWz3r1dZUva7EwMwmWbMf8JyV7naPaypSa/wD5o
CWLf8FvRoQXuy1IpxX6qeI55KVXCa7cQyWpkVt4fRJsw3HePx5GFD3pQNXXO7Qo7
UJVkTqVsw5/3KsUtzrNeqtauKtESBv7jHI/P2ZgWzrgchFGFGk5GY6LCfxX0aEl+
At+Ejsglgx5fUC+fnfNEN4A9kxL9/MWeplYNDD+ahdnwX5I5GXfbyBjtIpzDcv5N
z6m4Tlnwc73a5D1a8UWewCX/5/CBCYMAb2nf6HBy61kk95f97+JQJPfYxfG4JwOa
TrZ9rz6pfzH2toBc7IngqYG9/qnHfcxZyWg28L8ZccMEOQeSG4Y9zIoKBLZEUhWj
KfHR1TeRTZ1ZE2wKJsIBIMUuxGM3FjbbTkE6F1tm6wRUMsoP6JCv6UCY+4m7h2nq
muZQCDsKzlPcEdP4EguDQO2RbWmqzluqD/TKhx4uj8b7d/N4OqQduE8o+3k5DuEy
+hT2GMkp4aiVQI/1bEDMw+3Ccj/BUFrqujNf2FoO29EPX/G9vqF+roXuiidc47xj
Ou8BPihsBFYIlmoS2LKklsAWvtdKw7vZd9GFUVWJ9jihUX8Xul2ZSOOBgpjR6Amd
sNWPIlLaxWgGTUSuOEFD+CR3wNvS4nr5KIwWVAo3/K0DR8S0if66XBAekq9p8cdW
j+oJzlTaCNXjiZC+AvaRNke/n91Y/FYLbU5dyKAi0OtJvf2Kap9Y2AAsz4sDwsCR
CIuLSIiRgFxY+wkx/E+3TgMr4p5aOUsgKISMpiJfWwqsMNni54PGZPnDsCa+UN7k
J+nf5s5QHrnCekwweS9CDdd5jFLwlal70gTTgE0PRYrWm2arCOPPwQhtI/lzI0Fu
H0NYgpzYw0vmhW7HSz4Oyw9U0/QVjnndFbnaZ9DoVh7eQWCqWdwIk6npW2SC8CHw
/IkH9vmPYDkA5b1hw1ZTlHDjc9VQ6QT+2M9s4V2IHpJcW48U/BEyNIwOwMGeiOGP
rU1AA+zVT+eOTD9k8fUManMNm7119grC455tVqjWkjIzCMUJ+4jkdXODv2vCaKXC
X/LFydG7US7sfLWfGe6bRyVPJkvWZ9N9iuLNcUD5v7LxP2Q1WJ5diTW7f2bw6UdC
wI5FQEkhSLmHT4dCA4WgJeQ7kjzykJpsGm9EuIQqvhSkCADqQ3vd88+mweuM30kX
JNNyuXOPSb2dQTNtFO2vPIuKgx8eF7RS6LseVOoB+xzGJcxh7phZ0Rnf647NvwJU
O5ELlpJPirX3fchtn3iYcZRI/Ehl5DMTNSC/VtTyyxKCW7cxQAQ5RcL6Y/x847U1
v16ii1ydktb1bXjgnMxOlcYLtufubgH39yai/T3jm90AmyymlEkOsAYhb+if3SZC
qh1ddFuQn5FlImww8H1cPNLApPT0gFsj6vNK5wuNqy6l32/NGr1Iwr8ETNFSQRe9
aKL/Rua82yqokHbc2EMLW6MN1DQFAe5yImoVjvrDdFcgZwXQMalyG/LwGPPeTtVK
1IQXUS2lIKpWpav6u+7xPVGooySF+3tOsBTWl4wUOKfgja8EavuyV0YShsMmIZr2
yBSTf5Njwmk1V27hFxomdQlTsFvF3ig1KR9dNWSKE5A6l11TPfO95muyCvTtnpuf
i6Umnzv5tWgkAJfcb+Q26FLBZv4WLNcW4tXYw/kjrFDI+NVthYI6TLDbSIoYTjZd
1GVkFt3jlYAbxfpwdr/nB77CouDsQkKb1L3PJmEAJFRYtB3Rhyu20XFsic9r5DIF
WIKW/bafG/otaw1uEbZI/pCyAeAOpijo8IUz+9r16LS21KpYgOiUrwC+gTai15d9
nP/Klhy0H2hF0GXk+wEqdoagyCNS1OaE820AtnSZdmZkyA9uIZ10w+0qg0DuDSYn
y2wsjoagzZsvRN/r7wusJCkZn9YwG0rfujHHXaMd07Fib22LEY6mGKmI4qY6fULY
IXKfLoCF3X1y/s6B3CWs24GsaBKiPzQW2tUTf9ltVgVRPmjSfzrC/xhyuDso01P2
dHtiZiyfcuydecssp9LcXcgUr1TBR/PGf9gdys64K0wCwfZHAYedbtlzXPalm/3x
6DyirjnDmsAncyZwtAOqEE+xyYVMxYfqwtzBiHTdnOL1pL45SsWJ8WZ+NBQHnQh9
s2Rhawwo1LwX6AnvXwWaTJEBhuJgaqG7DHSubo3RzeMzaY4MMyeOgoAfxbFJa3qk
JKETWVvsM6lPfGu50kqkF6LCsPZwRaq7qbdlHL7IWQidisLKDucT5wThN5Qo5z/y
HRYIRfFbMuueVKHUDZvZ6jfdkv5NuXxWGYxo5FXVdNU6x4ZJEZ3RpYPNnttC/aGz
sGKpC6hlWsLIirbdxvui6bP+O9eq7TjMsFe+ntTNVhqkyGMbNYiylbg3nyAIG9Rf
qMzKMJl5gQ2+JwZfRBKGLDikGVXh94EzFXIEx5nuPAv4aBFkGwuEvoy3m6JfICz2
DyXS7jOLqmR+zSXua9/L7QNtOtJAWdWGlT64/f2+nRqWoG+pFYqMOy+UU3Vp417K
9CBiJar0PgXfhFcNWyjC5iGcoT9vdjYhKdVDBqItEg1M9tRcyvI4ymEJ3QfZYrwR
OJ6huykXBRdW5amZ+6zTvx+tQeUSKaDy1XMPwnh7HOnEzQEw7EV+bki9bei4UB/I
I2XmlCYECiQz9hjTyBhddf2NYggZN+ND48+vjCac2YI3a8WroTcK216SXrjDFnc+
DI4h8cpHOV3srTTC7GrFJcECzQWqtMJplDOoT4BaiMYql13wEmFDuP4yW/BCC0Kh
npus9hRLBZxE7S3DtmXo/7VoevB0IakQaHiEaPxJzA++LUtAtkZAFlIybVc75LJJ
HkV5XhfcZyJXmlegu09DY0t8kDlEZF4dwl3F3f1blEBrJTb6kL03+nzv4XQMi92u
XdezfT81aC+ZBcg1BNjHqbrwCppHn6ekUX40OQ/CW0qXk77lE5LGWeeSp9n+u3CY
QYMGV73plzeT6gSxMDd/Fz1AYfddH4zvsEiUeBwOUE6q7KzWJGBKT2fueH7TwVXZ
mfO6/PBXzVc6U7uLC++0q8xO5J6cFfWS7CP6YP6oO9rZBZ9TaqYCag/YLhrxTsbT
ibdNV6zamdrslxiDM+O49zqbwD6nP0ztBZarO5m2bo+s4PXc3zaaLX7SefD3MS+Y
hNGawcUNS280O0Yw4wMLA2zrssGctUAbxyPtXeBcqKWOAlT9XEx6xVqBwISORzy2
YtYqeQjxmmyjI+LAylAxFJnCFcmuUaG+liKRhKrDvWiAUKa6LfyUpIuEwFdjSePB
rcu9WLhhOigfiZxLrNFa7Bs8+b2TCgu8AlQ254ljSWclLOh4DnLaTDXB3w9N3iWt
MKzqo/B95F2iZi2ge6I0UIiMnvmMAnUs2ZwGt6146qICBqwRd3jAS3ISP2bPWzYF
Dt1VHFIEXF7jG0HcWWH7svrafaq7Gegmfj0cAVJ7rsJ63Jeys/7Pqq/8VSQZhzfH
IP0fy4AOFSopll050l3Ng+DJeIyY/+ByQRoSahk3l5sQ9CPzXWQXjnMrwxAVpnmw
b2YFBdBNALJ3u/DvbfrJwU6i/V3w4jbknwQJRzVoq2N0wqn05eLFX6hO9wrX/+hZ
ysnFylhhro+pE2Ff9oPR8mU4GpeOpJeePZ78hUWEgTo4huPLyomlcZW6uqMZLcj/
xaM2SvuLCJybbbiLAhcajRSw+h2SIcJQ/FxgDPr4mTjD0ykRNd0JYhx1XDJK4IaW
ibFdPXZLINqB9MCZtzploBkj2POZi+BWQUckFJEIjUmD2UZdfDbYW7Bu+7MTRwXA
CYxfnGGhWrb4nKi4llnBuIEC/a2fm85pZAPFNtxcWhZRUZjfzpWKLoPuZoqlvVpM
AyvTSQyOA+h9WmF/8UBuTbMLs3QzVN94WWJ1xOrCbEieg2abRx8x+8YOsEJKVwp+
V1pYPwOfgOsqFPn9ZYh70Mw/6WG5egSDm9YM0aYMmeUaDVamxAUmVSHwdY28Azyx
G5JpidJASzl++tYan09as/9qHADJoRXwXl6/FrxLloc1s56BDcsLNIE2QUtZb0/w
WUqo82npNxrM5zzPMWvdhM1qDqY/QrxeapjiNgGoed/pBmGP7ngD7e3saFZ8C3Fd
JQdIBq0DdRAROqmRtrZIBxqEOEDJ5E99xH6r5BhvwXYMoKmbyCN6khbH/3asRJf6
hbMHnSlbTMhScr8LJ5NnCxsKps641ToBoIWA2FMohDN1+6tC8bMe6BP4V0zUofAa
8dsHIVQQRAcpimRHewq+7ro6Hp6h2tHvwU6bDHxCkjU0zb5c5hTEXXW8bpgnEfNg
/dUfcjwNNWLUlsWbJd4cdzH+yaC3yYjAKx4TuPywWvgcNhHoI4fMOwXzBYlfwWdN
ixcNTzN8sbpDyp2q2C7PFpeup9eJXCWJL5FA+rgrfVxHj0Nizgxm2CtTy1YwuMaE
pxqDMC/MF0OaVOH+FRFKcl74xLgQ6mwyvYldAxrRdTytMOPWXRpPa9M3OEaXEFCS
Gjbw/JLW0vMOB4shwXmkME6sXe+PUdirXRLHLcApVQzHArZkak0iWvK/SK5ZsgKq
OF9HEPBXvjnntdo3DlQd+K+h1R8LETfMC1wqs0aUZ9Y=
`protect END_PROTECTED
