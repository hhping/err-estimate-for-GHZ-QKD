`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aTvXbJBbW8xEsAk9sTgn4rAIoGPS50N/PN3Vj/D8jY0RJtjr5bcWvBWqKnVSp5GM
Mx9Rqo5HizJjgQlSgTPEOQFScqk0xIbxSustbV8Q8NNGuGn4FLXU9YeHvpWA2PnP
fNlb8QmSpYaQ+FerIwYsJ4YCigpx5feNawDRfh2kNQ7y9TBr+79SxAojOzELEpLJ
U5nNcsz7MFoXX/5oH2MLknzxLM2SGUOWvXyKhuyJnVb1M3ZtVHAo5h6pnO3eIcCw
WDJR9h4P8VrjXFN8FB8BGxYkNpMi1OA8k5BqPcN9HGY6L3l2QRcG8tn2Wvtm8ahV
50ury7Qum/32zdaDGFRWUf79L6/zl1cU3n1BFeANNCOqviuz9C+DWcAHJXmPGKRf
MLk39HN/izAljDEr/iY39NEfQTeO/lHqWaP8V99jcpKIhxp9aiB6rzkSsBFdzf1i
unvE5vagTqArAiaK2qvWxN/L1TebdBzHsCb+ZIJkgZJ8xfXlTvLR4r2NMaEZ/GvE
`protect END_PROTECTED
