`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
556yKeHd4R0FkO0Tc3knrLmcDw442kgle8jJmsCy0Y8TdeVkCdvvdpbJInaXZ1ag
gwlkQQ6gxfjZSZ+oXRNlCEGF8ji0DmzOW1M9ErkqqiNKye1GhzsE2h1l1o8/NFi4
7A8/20kSiSFMpl2/zsP1H1lJvkqmCsfYW3nf3K9cNUoydO+9akw61FBecyqZkqFN
rSSCaRoKFv7Guuf0qEwj3EwldJPENaSypn2Mq0+of0bWvAJ/OkpOhDr66eUYuW9M
MueEb4FalSQEru9nAmW0YK2yrEA2gIEVZcVfngreV64FGsoPSUbdU78w3E5f3Ukp
nHVDZV1FCil652klVTiHU3vhqfbyK0TsZdR+8hbMBXdrsTmpmIgVyIXTqPn9fnOS
sL1aY7TWpcahZF0xOoHlp2ZS42I5wS1N/lh6X9STufjjqQbNAywqmlrcZCHLnG2U
I2/vHzwU15PGU9nZKro4mdhTSDDKtm5CdnGeTjMLfQHPle8oh33QL93yWy9tzhDA
f3b5EOEcFGG6G6V9RTNl60ENqERgAMYevrnMWtLRYCG7ew8QgwyP5+zmF41XyEC9
lktJcNNvwBrJNnllrYJyss+A1iqXlhdewP8+21h6Z4Mmgn2sB5ftQuDJVO/TgC5T
cQ3tkRAGfE4ohRPrupi0mhzamYia9cgKZwaNHVbxuUEs7nzdJWusw96skV7onC2W
kU/LFPyr+e6/liCt8OItRfuxrMKd7sMJzrGyebqdBiF8Wuiz/Qd72Z9ZKBArq8t0
4nB2zaGdV9VbnTuaBwYEOK9KaOBs2XmU8MbAN4F5EkCMUx78g6iMHMNyma/o0Um6
/19LjHeYrPe3rLK1sg2GUjAd7wUr6imwolSGCgLMl1eKFfuO04c2xJm9+i8gSRpA
+M6KmDFtwccSYddEh7XAQnurYt9w0Rk3EsACy/n3wjWQQs53Q/L4MqaOT14mxE7G
Bznyqqy6lnHzmoNcH71VpMMXbhB7rPFVjqkn2vwdytQ5giii/lo13N3xYtJmeZBs
Wf7/Xto2DwURaWFoC7mBQAw/z1Gj6+0TSYpUIoU+Vv2Z8NIE2j/Yst4aJPVxqIUX
SDw3/sB5Kdv9HY7ofA/LczGYZkqsnlIRwhViyKfnHstHS7CQFChTZ598sEdtRluW
uJwJHpZxhuIG+4fNycR29OBSqdwWaeVr5f7fNvZ6b8fF+NQg5J/OXTQNUNoTELMy
niStqYGHPF47lLcyjUKKNxxucTKPKkbtYdy9Cu0PBl+Bt9kpqC6K/5q9OUZg8tEr
T9782BqaPWeA2yTweUt/vCnR0ioi0MBeszN1cmFzk4aMd8L8o8j4Na77NnY/O+4B
Zy8INnw3FTF6mQv94bPIi3jhITFR0ty40ziWJGvVUuA5+UtnRvd+Pn7F58YJAsZO
A4cnfUCvOTyptYJGjKaoNm2l3X3cXTYhJ7jMdr9u6JiYTU5MdY6yDDvMP/fvzIGk
aSMjAPEWsoesdxTODKep8jV/+z5QzyHNBJMKfTRz97I/fd7VRe/3Sqvs7tYq6lYd
02+2Le6ZLtldyS7HxuESadDbgM0YgoOa6wrbZaO+5zwoxd7srpvq+WAqe2tcztbs
3VZxU955fUptd/zuBT+9zlADwOCky17hRLd4HOd8tL/Uin5cqV6nD78MNyRYRnJI
DL880pQYNXvJ5rBQvEzz3YR+yTc4p3OwOjiBq/sUTEh+7ZsUduMA7vD7xKhzXkAA
YTvajUbeLw8OaVOMmgLLs/Ngf4LMNOewq7FZFL2C/52rrjyUaK7hlmCFnZx8IsFC
ZL++DCd+iuzgmsSP+UIn/A==
`protect END_PROTECTED
