`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
poXvNngZqmfYorWwKj5WVuwzT7/gsgw5Y1g+st5tGxzA1TpBylGNGayaqb3hAgE3
4+XJ/VT7YbAeXTGj+kgNdLjSXUwJXUrr1MELf6KD1Pf5jkHthk20mTt8YRkI259I
gREAnUlbRoURIgHhXoFBr8NEfaaCQ6ryyJK2mCxqG4yZYe8Gn2NJlqpyxatdqLjw
0Z8DgIco8XHnt6WL23JbbX3xf4K15lg43aXNMANuJXu2zDbd5iDTpDn6fSzw7hss
Q1B80GToDy3iSmFq3ogMcsGtHRaawWXC543L5w6BzDIlG8MzPQgKhPUygEU71lKr
lTasA3sUzjYoors9k+UMKJsQHCRSsGAqJYwwTBp8qUIlrXZxKdV7CvZwQ5+sZ6bv
`protect END_PROTECTED
