`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ANFAv2b0SOf3HbvVlnbYX5dBt0LA1vuAQ37FUHmoG/Bx4iLwyFlzpSA2eoNtaDSH
+niPrYm/Zi/BMbnWZb9ff9nLoeE1i/mb4v1DnXo3yTjmj8Fnx/0rm2miJyqMMo9A
9VbCZUzxWd6H3+2lqZgowGveujEcxqatHbcUw8lqiyvoZeNdiqD4cgtpbpzZG30i
p1guWxYNA4jfuWxGK/2Yd0wO4hK4+SICcBqQR6yBOLTeKHd+fmb8bLbRQm688LJO
3zhQycfa27dSQ14+P10EyHDKio8ZS5PfbGtGCfrgLAnxFsGu25Fdhfj7LC5g/LPJ
4l54/5+5Ebyrc87XEzdF3+lMDqPgSDOMfT54DHplWN4PC2YxuvbmlQteK935DH1m
nkqdTOsbMXW1oBS832erhZdXfggvJxbX+SCnhEx/ApHDgZmSDQoDr+KcvDAbqe9v
SCuq8nifz1r3WPAF3n9u3yRHswGQ2IyvCyXi0kfIfVBug0PAbEiQKgjoOO/I1zEk
Q844tVJIq0LEDk0g3wWh2oGuKuRMzHOoCDqiNemv2unwzIXMxEtaU38lYURQYD5F
EvfuKtIP9HyZfpXf3MekhklvN8TbpEh0jcCq9uDnsTGL6xN33jtDEVxsFU84NWAQ
HKBHYR5FOQzjW/skd3fKtvZcDLaTjUVboHTOXck0rgbpj2SX9WQ3tPjSppf6WZ5I
GLkxHiyUeyH/i+vIP8SNVlmTdbNdqO2AmO/3xaZcRcewZcN0+nLjUcGsPJQyzdyS
M+aJmXSigk4VhhTm2qV2++aiogOhO2KP0bJYZKV4XA60i9LOI5JTkb7cAq8fm79G
2yWSclZQatZ7O6w5JNCvHjg2CmdNjJrPVrQoSxw84rZ4dHI0vtJT+a7MSzphPRVP
A7DwLwy+tlhHeDd0beACgpUgRHsXuWx87AYwwQpdXJsH7woTxLB6l2kdL3r/SPGQ
E+Vfm4StD+pstJCiD/PmvhLz/WcbetDtdtYmB9SJVfQ8KUJXwvZYQ96hSzGEr3RS
5yz95ZijBzegI1KvZqeMGGLRVeS8VbBUwuW9mRC65C0iqbKkxkYrLCcVsGwaRORU
`protect END_PROTECTED
