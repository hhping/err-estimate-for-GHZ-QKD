`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q26PsvtTePfXaoAxQJ8xANcJmLRaqKsjM4VX8P8c6PFW7LnwIGubbnFpazlIazN7
+bmpso87DmvIyvW7914lYm4vyjRKVUmz+fDwy7hucWE/dk1gt9PTTnXFrxNVYoy0
ICG9HWmLQ1f4orB66QY7kCDzPQQRWH6Q3MYFDZo0by3CLZUUn9FgDytodXLOqR0K
wEffZqTt95W+JTvOqFOdCUxkGrQbI+qDgoBiE0k3dCFFk2kArT7RLwJ8vMOG1wV1
adArU9FZpksynd6kEl1mrOaUvMZvyT/Ko6OKuaSilZb+1to7Vvwh+4JblCT8WGi5
BQgXVsTTJ64naG+WypFSYChUrPXRXNrdaxXxFbnOWaZm6u6R2KLPjv/g4svGzdov
oQLEA7jwq7mmKIk1mgORfVTKbVw53hZ2RV5+CzJENBSrxK8O/vnmPumsbW6L27zp
G7eE169OxNkSsTRYE6jb3x4hestqJttIM2SLPZ/2zhu7AdSXrCakwumS39QqTZZQ
qGrYvdRJF5TwitBHUpFO6MhupE3h/mQt+wnroBiPtXi5Xs/s2+L31Oo+QqPvywEn
KP1j74Vndj34V+P28WcG+jhXrh1j2q9izHBKyjIfScyyZLqxKGqhJmgfnY3Sbhab
PF0GkbAVikxCt34K2Aewj0A5bIUWEqS48gSe3+jPNY0o0x4vN2wQAvqHX717IZQw
Q2H6GQpMRZvCFD2MrWWyqwyctyFDJg2g9N6E3eV+s+thXC6cRDY+UkFgmMR/ycC7
q99zQ2fvoCXn15VrjzmtLNDeeA7dOWx2OqZYbp449LalQkju99X//svs+7Ba5c3h
oWcejWBo36AG4p65mXdj6961BEqYqt64nOr49DfscWI=
`protect END_PROTECTED
