`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DxkNHMwo5IMsC2dHdKXIAolzs9UgUP+5V1Wc/TqtZq53qieAM6rVbiTK9kg45/MS
TFxm46XWY9v34HWCq1yd6MQ+dT68c2pq/JT7vthsZAOkeO2pCRoo/LhfCGBYYb/8
8vMWss7YevyrbOCqjj9LfQ3UKAtTP6fJtY6c+z+PwPbJYGdJ9+72c/4Dd3/BW6k3
BcCdxN0dBa5YHLIw6epVJeBXEkCpBmCmqi5Qlrp77qU+DgqEvWwurZbAwx9ym7Yy
tBGjVExq0lo2Nwz83gM1chAwLYos0W6Qp9Na2r0AqPRSrXmmKqMC7//qQ9fRNgru
ZFlt6zg0GMWWSOXKsXw/lslEJGE2Hq33mXyhY7dRQp1u0J7SMkrPaSIsaM4pRaZt
/+tJMQ3CWcLBDeWJsOWlIFPT8A9B3f5MqDuAfgWmbxmDT44DFjo45IZfLe/L97SA
Jnh56/SLGNfYMsK+6DjJU77islDdyIPOc5/Ps1xai8+gmsgvYeuLl4Kpo8J7qZR+
YX8Qz3ePuiXzUfDBDy6uYCyOF9sbUom9sFfO6DXu4NxAZZ20umpgrnEY6UCeUMOJ
UgeJB3j+17rkPIbBnPgqQY5TRvfAO6Y1WDSFciw4V7K7Q5OMk83K3JA9qGhjg7Ke
1LWpv3xnW/p5ZnGTPiAwmCq7nZXZqZTEiszGhcDAV1rY/BnFVd6kRMLSygmCRfUg
FmitKS6KGL6cTS0JMJBxtLlHjGajsdHjBURsq+cPu2JXEtFNbcmLMeSkDJ3g+4yc
XlhcqO9dUZlIbbhPRrntFM7VMIWRMwMjWDtm2InzSuOZV00NkP+RBPJfvEvB2o6G
6KsDpxYSZue4R+mLJ6YJr0F6qlztQOYolSfxJflJxdM6UPw/rWgE+jmId6SUa31e
feqBy6QRyJ02+q53NHvExcPhZxe/wG5E1L/Psr/sJMGfCkyKE5rI6koqAqF+RK0r
spVa8OyI1I6KloEA1bIVth54IR4jqT22MP+KroLk7mubBupGiaWe33iBkYxchsuA
NR3Srj0/2L7ZFsKPRF5rWkfJhG4oX4oAqCU+2aHDg1RqUlYU5bs0LOm5ls3c080U
n2yI3oN5Re6ZZNfl2KlJ4/esJr7+t/V2zYvdWbk2/btrzqno+jJ6/JAqUHdwJJM5
3dqUN26Z8VuAjw8/amczzeqPL8VNpj3CQlT2MNXUsddBnRAcBAmOV6GjeYIca9dr
bpUlZ1Rs+1xKyO0kxaGy9gquhorYt7yQmHrL9kIYg3YVWpf8hfhXRqL2zbi2dlzq
we9gaqeatSXSrbADTlhNDEtinWMt+UGr2TqrmfNp1HPjP5jyFisW4Z6FuGMTnAAs
covlIbPUssnksBnJal6UAhtAsx3ZgvQqXILjyJALalA5usUxw1j4R0HIbIvPbrtz
SmdWMVCT3+Miuddhaws9mBqoQ6NzHpdBzylbeV0on/JwxWf9yCvc1OKdjVdzCznd
rbwvI8ODt0k/cK8l83B1D8ziUqL0hIlYiN4962odsfTnCjxSO//9jF2SkDtL+yyU
ZUuExr8XAAcsiO3pcOZ3CUxJRuNkt1SUJbCIVuJkcwzlqHYiBWHW9FDYBCwI3Udj
thF2H5uRJ8XHkE7HBXK4kw8TUyb48iLsaX/LiUg5Cmapu2lB5gqbyfDapEPNeG5V
MtUi3Gg0iFrG4oGveN+Iu26ZT6zW0OKCAe+1nMM5tqF1zGGyB9g5kulEa/ZTGMkL
PeUdsthWkX6t/zs8fS2AGa2NzslUCt5ccYcSNNDooqILevImCOMFKyevbpzl39rk
fHh71leS0874cEUPX5aGrqRhdJZr02GEImHvROs4v8dbnBfnMIJ8l4cwNxoLseya
+Exlt+ESfSzixQ4SV4NFb6/ePMvqO86OgAs+43oMhr5wTIU7ZanhhxolKym06EqJ
P5l5puEwCDSFltRqLfG/AEbZu1U+OlX9+HEqUKsoEy8khauXO1hL+a6HIVhYX3Uw
63RlZZ3o1PafJ2k2AIOcIfLsgSjfGTpadMIEuwr2yIwM7Z28nJXLWY5MqDEB2H2X
XmBQGqIx0ivyFK3PdcD7ZsFgp4MoUoxHhfaH5GMekFDE7bPBNQvHvO5v16/U9UDC
y8IgrDGpbC75cLN/Z3X6ww==
`protect END_PROTECTED
