`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1foHPYIP5q5Est3CkJtFdcnRZZ+B1OQBXKp46LsZrGC85cvM6Hvx08DKLx4AtZ+6
NVF5gCHteR7iwBoZEIsl2pQh29U1jj0ohnoOl0/8o0LEc4fv5kbKuEKbLwJgzwps
V2yWAnn8HjAr9thzWgeKqr2vPobeiKIPBzw1V0ilsbdsFn7Ol+6z4e/3rluIfBzF
jRbrD3ig9gENPKqx3xKTMOPe27Q8SxawsjJNmFUSgxsuQ49fz4vin4dhqVLVUdXU
E3uXwshv2/7XQvFYeM1XJBfLSBEZHdqTIDOwwoiePk/EGKTK1yKUOn2Uqw367CnN
DohsRrXrLioysZcxiJTNTaLlxqNqJR0PTEPKruTPX+J1uX9cSfnKwdCCkbqU/Xki
bvsHiwHXUGSsmXQWyux5EYdMFIGqIWBKwpeVJ3jvAas/Jd6TcDlSVeZPAy0p5k1Q
vBPoAAvR8a4Vun2/MEhtSuoMhXNXOn3RidQuYJnPlk/U4xtxPTfvXToszjE0pPhd
AeMpGbCw5bjVwCx+TNoWz7JOY8aNxn/7U1ZqbQxL3M8/NM66+VtHp0LulY1fHjf0
6zTSpV8/Z6OmhJLM5pAkLSUFfXuxpN4ANc1/REPR8diqIz3LwepfUPRlYcKz9JxE
1+TP3JrrQZ1CexcRnWTwDyLuKbf6N0zP436/JFxgBLu9brX908qNT2TaEETknqZN
wcQ+QhPwKm952aii0yXM0Uqv2ev815BYZbyprxvG4GUNpYcV5GWAuqf0/gKAVbkf
6J+RvSEP7VsQWu1lwD3aPr84MS8mAH/NR6CEaZJ5DCD87k9K8F3/zl4NzJxkKWmb
0m/1RW6JMZVUk2noPwNJpUoF+r0oc3uBbx3hugqR0Luh1smFR5tyyrA/DOTjHnxP
DJUkmfrHLrXaNCjAFZ+h4rES2STjKLOotOCJ7DaeMVE=
`protect END_PROTECTED
