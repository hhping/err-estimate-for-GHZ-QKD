`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z6XyO3LmLzXobDdTFlXyhtrWOWnnFCfS2kcspYlhmj4HrXiVAyX7JbFzIphHUvU7
9w4PZ+w7idi7ekIUPIoNHGydrHVdSUHbSVDiExQSeLacA9gJKIbmkVYeNQLfzlYn
uhvE55vb3ls2F7vBbO1rpHoNdeIRa6VIaKoGSdU0fNji0KxAatNPFZedXTMc46sj
lRsEZ6nhstKNSvGIIrq2Apl8Z9yfKcmvY+wyIrnKj9NOVXxASUmSfBwS/mkkj3/I
cTkLVl2ECaf9JA7FQcWW7Pz5BOhqLF3J+jBXDI5BgXONWKC35WHp6jJChXnnHrcr
HXRM5CLYkDjIHEfdDX4q3xWvCgLZgTsWLwZ5PNXdk78iK2nSWeEQRwk/WoWiY4+Z
skgI/WWOkbY3dIp6amfN7QMPQKWX8Mc9HV14XwS55VWMBwvldYQmC5kihRVTGImb
oP58zAH+XLjbK77EO67pTCfDZUMdcsI5fjN45AgLWnbwh1i8KpeKlmRTyGUQtISw
MMkelNL1RiYZxvpdExsWM1iIzCk03piXyNbCiahEgrBPWGmS/Ks+7xEca9XrlzzE
PxMmb/ilBbakLCjMLWHX15jgMDpDmkgguov3CSRJXi4rIeBz+z1FZqaKjktCJTeN
6Y3/0MFpWsVB8ge/rwSZgXzp+xdX9rghlKJV+v8S0JoZFdKo0vYhIgqH7NcNXqNC
tHYlMPFbWb9j6Qf6H1GB7A==
`protect END_PROTECTED
