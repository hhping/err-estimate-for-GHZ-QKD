`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e/0pLO0MZsGiGmx6i+VgmHmlycIkPyZefca/E7KaIF8Dv0jHOJ/KTApxbv9bcgiy
xhGE3OmUacRUZZJIYA4uKccL44DFIoxd4UICG5KMRXuyarzpvODMC6rBUkde0u3d
WlMAwrVl8YwnAnEjJsLACTnak8fXqP802trH1XNwWYAU5Rt0MJ9QKq940xvN28tk
Yjcvsy3lrsCTyKucX8bvbfYR8PiVF+GLlzelxqWHIRtduOzlerxfllGWyv5Fq2cf
Xi3OCgMQfWyskyvskhPXalJti02ciqRKozaKDD+wNkGEJYj5+XDRUFocjkjwiRYx
6MBaN/wGhCS8bIcrbecNZwI5J37t0kY6PqmVIFbY2caUCXZDACE+SDpDqFZb9njA
`protect END_PROTECTED
