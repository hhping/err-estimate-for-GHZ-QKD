`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gxM5ElRR4H+PZhjn5aDffsQzKxRNKuFLkzWfmYQlm5w46tstrcrLm0c6qNe3N35I
ah9VUOgEVJj/VzCjqB4R54uJJz8+iSOh2l/GA2eggo54AwPAftAFMa6V5GLnCrBz
JonIUtRb4P6+WQcr+AFNWmbSDbOHmvTuVSy+UCgTkkNQgu/ehO9I+g5JJhU3tZd5
YXmbkNXBHcEx7aIHeYrDYnjsYnDDk03yEW1T2aWu0PACcczJact/npsz84zhmacl
IJ0JIGc577JJD2nSOY976n1spQXpkm6HSVJ5LTltyocyzzzpCgIcbu5QX/eaz7ph
nfX+4tuDBWM9iV8LWJuO9Qvn8op98ClGxYNtbWou0qLywDWrk4C74Y6fAd/OhNrR
eNHVHRpjbqAOZl0BXJUG4CngiP86GkYBYg62SslQDfnlams79YmJ7DHMsdXi2ar5
r/lMlFdv8Egba3DXfOEnhvw5bO84j42Q4jKq2qQlq0WAQwe45U5j8A9zDf1pNOD0
tqwa6NyL8BOecaP0lN9auejVMkdpsQ2ZCCzztL/1L2sEB3iLI9HtxOkJVg7xupPG
2NpfhmimgV6prBV8F1FkaUv3auPF6ivqPV6+PpvGltLjjB4Ct7KfwZWKTkfCeKkv
`protect END_PROTECTED
