`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UjmHmv3ethx/lTDN9sNgDYJkcefsUlW60NasyphyYJiUo5Z+XQZF4t0kVAlSc0/A
fEOz1v4dMkJhPwQ8qohz+ME8kMucICHeVli8MAeRc5rMeslAJL1WUXWfjuD5ZUmd
5ctmCILi6FIjXrEUh7/WwZzwi753RdadpUQNfhhJnTwXJKc5qS27vjjzg5+fFuR7
wioKDBSIfAtNGOTsYVpRqbAZVDGP1Oa6mv0iTMIQMEZK0kFGoAX91prZNQOxNGET
ZWKGshS+0EtTVNFQ2oNiGFwHOrf5unJN0W9OSjkCuf3EgX5l1xhfgrLPydDrtEeo
4Hlz19bifP7L9UjdzIzQbJnXRd3KEDLhXTm6PVaVeRgz5rFbwaMIM0iSDd8uxFXn
RR/a2KzCENtdIJuTiRIVK69wNWVtGVqFlZ3pGzpM7iAeIO3WNwT/vBpau6cYbqHZ
AZPPiTVb2UnL90cXqmzZaVWlSPRJ6TH5ci0D5ug0gHaY7ufGk7Vlf26J9YSd+XjA
FG69KNoeMesQV6yQi2i3xcrSQ8SRWoVd1sLcQSHZGuEIfMiFzXhu2MffXLvZNMjT
MeVWaAHlN8uLyM9DLI6Baa4IuQaSrZ86bdgCpGx61QULhd0HBpFpC7rKUZ7UMsC2
dr8twt6rF9Sq7Dl+YVbd1feo9yll3weWm5mXsND4umiQJSWeus5ACtGsMHII0H7V
zvFhULoY+evB0QYzga2gFg==
`protect END_PROTECTED
