`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lCl7A9hAAmZ9YR5ROnZ0GCbZGyXE4IO/e+Nen9lKp44iBu1hm7dUxBd3wCmXokka
bhcW4PBFnSQquIRJBtrjWcE12wYxmElp/oABUGbB1b4YjaLawg7Hx3g66zZYTyCb
4OVT+kw3nhEVgOalq/E/k8lWva4ONVgllg9RqMzmTvSHWyHc6OsvubTo2j1tUdD+
m1lkAKm1lS1X3LXW4zbZQ5pyE36I9DhFXJY8UcrWMflQBI1Tr7q7+37gemdWdnhU
lWiyV88/qJhxAcN2PkFfu9OpitUM4CnDU4rTq6HP9I4LhCtlU/5UukcCL/LqMKXv
HO0y4y/vKc1N2PJEVEl2NY/2JCT+Rep2ySh0BU7/FibWdp1cMK8+UCGuQQhfx4XM
XVUYpixAL8tNNUPE2kBW4ugvkJ/O0XDsWD5+o4QaXEC0d0Fbq0kXCxNnDHfT4R33
o5qQsuPNgBzBlEdajFrxOw==
`protect END_PROTECTED
