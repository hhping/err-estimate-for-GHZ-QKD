`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nHXAkjPz34HdvMyDRZn2nvnMyERfrJPewP8twpIbwFgthaekfjJ87BUidE8t1Awk
cjthhhfF4u1V68onNnh1TQAJB5Q7OTin4+FEb9/0M37xkwxUz6lYiuIS++4vRdsy
Da2qm/ViGpuitIHUeUSVIzQRn/lRPNkfnVNFtLo+/4t85Uq4VtCvjF9HRVFQMrwe
leeuwZ0OT/B/rb2RGr2NhKx7gM9QVmF1vpTW2IB1/HTuZIpebpMWOc77LZizs5vj
VuWuwd1ZCwbLXHr6Tq1XumzOoxzdKtqPhsapTW2ACNxmLxFyWgU4xX30OAJYgaCb
Om2uQuQLBgA4opaA7oXaCOBXvrhBZFWzO2op1Q7xhxrIDXiMIb43BPJB2GAB/uKC
Cnsmx1y07y4rn2ItZKha/a+L0nB2B92/1/R2gdHFxv16qarVltRpQlFyfb1ipRKx
zYqLuTccwMIMUrb/v6J7KU9kLXfDhZZSxeP32vKluF1en+MJPvFsN/q2Ha3SC0/C
W2CbrQRzKArquJX9INcloRbpSqq8fyA4dVFm/+IoPljRvNcsfbjv3WcYHDLL7qhc
UmHz875V5d3lvzpNBEja8FKUb322AKlez3kvt7/qP0YCSdeScRR35MrHTZp48fOe
2KKNx/o4cDKzd0ylvc4UvWVQgSHNEYo61VPoRnQxYucxJAMmgnCSUMTBOCidb1jD
m4FybgjAsGW9oosnIC34bn8w+M3X9ygmJVmlHTahWzyqIuvKt+Sbh0pnx/5ESXe2
968BND0gWSrlRDTm7/BaS4pS5aM6o8UQu7MhLub7cjaC8HtA4d1VQNZAlF8FavqW
5E0FaOt1MxACW7+u95m60pPdOnFSbbIs6VfxDkPQUNCCwIKuQCwZ5+yKjveAsN4l
GcXHU9ES6Nwz+whGgfEFCdlJC7npWxpcUROG5bQ2C2QZNOTML8C8LFJoSFUXPxs2
Bjil6Y8l1DGoLco23PZX7qVL9/78Py0d85FYiQ7xehKHK59BVCeytPksItUHEkZc
lL1H1wy5FZmcd4npeN09qMwuDHWxojApofCQ1SURhfb93bwvbvdrYDMmPNAKxW1Q
9b6OSFoGnrCZLqZ280U5442o0WkjwflcnXWA1j5Ggz0iDYP69cY8t+0TO/1HojBm
Wb7VClF+iGV916hjGfP49i/tIxQGvMhaafE17U3Na7K+M4/DLoS3ILnfbazGY+/9
E8sgnXi1H7s3DUp46wTqbmORa95vd+xjUGsz0e2WSgznHFPpyt8ZevsvcMXpxkaK
akT5FM2SFui/uPXLYqR2H92mObtZAMyB+1j6SZx6oVXvX8w40oUiOZWNrBR+j1lP
uBKWuDeLIH/Xd7ctOG2mOWH3YTQEP06jn539rdJVNgzKJG5WH8hE7kI07cVlNDhs
umOAtD8nkHMAnWWyCfmEaAzDQUt55sTl+as3q2+WvdaAMe91VMNY0diV8VKeTHQW
vpf+7MFw8xlF7g95IkYEhM1gIk4fibvT9TJx91vWIGcnib/L09hBfwcpkcvWFoMP
kbifUKmCzrZd0sq0nDeZQ6/39S8WGUPX7qn6EVwDyBKGjegW0hKHtDRteH7kHVU9
LEOr6wH9WtSIrlUDmA4+/xboygcRvE1ysuvHjqxJGFW8C2oHu+F457nhFOO6mnrw
AMgi1C3wXksmUokT6luU+jl/qW3dLTvHkOPODsPqSf9hyF3pGHvC2cZFoBHsJIZQ
SbceEpIEIO6QmWJDpQPKVbxseZZW1FHWrHydtwCuiuXn0w2O+4SiVBMUEX3eab/B
C+I9uhgOUISXqIrWQnmW7uGwCYcDEC/c9hkQBvVOfyCHrVBrXjGLWIa7HIViTQdy
tUqhrb3NjaUnlYoA+YA51mBsnN4TV2KyAavfTJE++Rp35S/t03qsvgulhA+GeAPD
0gm1suvs5zn6b636RTUKV+r70UcV1/M0nhg8tQ5N+2rxhhSaer+8WK5NV4bunli3
niApDzZ2ULdnZwaQDy+fPc/fz6cHGZO20qgdiP4iKnHNxcm5gNplWpUukSsV1SIw
AaKrBfW9wWpp3rrpLlYB2kJy3xySejImMBgl3AJEC4b8SjZFjCAb/dyP5d92V7p1
Cc8MMi7jaj3tEf0uYU+jM892o6cK8Tz9zi1ZBX2FNYwhmW0Xq8OdhANAaB0xgm+T
V1woqZSfcPNTFN3VMfPuguV+zgppWheCoGYfWWdz+ELR6LI09uYDPVuNQO3ddJb1
d1uW9MCWcBJbb5fpPWSD21NWZ/Gt9arQDTyL+6+p28cphjd41niXJ0Wph1U0yE4L
grzhDl5rqyNoZiKnTtH+MfV1XpEyzpdVTdCF1rm2BjZl069fzeE/Y0/TNg/ptVfM
wqi+cth7nFV4RF8fO05iERTAPA1BjE+IzHSpofJXqW1SZ5iOpf5yJMGagB8TC9S0
VSZExSwBMnusrvGl6iVTN1or2o/o9LzjV8owNeXF88tfm5ecxAUAsbbhp73Fz0v+
Nt8UuaFslrUwGF+7kvRVW5MbA3rL7+08weim8qAZlOpTavx3+xlCw2ZdyHhU/ANH
e9jI8kyqKgORlra9DnVo6LAQmeI2vKUi6rAKxc5L7wIJzfTZ9qT2Ge2rM284kmMt
VIUOIL9n4ceJE8RPNV3TmwdqzOKWtLrNvcrfKshxAHjCVFMzHata8nALELEaf6DU
m5CwTWxOybTEpLnNGdS+tlSqgsKMOno4ozFWnvsK7S5AiR2fuU+oM6N3y5KJyrZ+
Px+SOEjWL9rdDxOp/X1OFss0+ApllZetuxVT5QfhxVEEixpvf44QA56o/rDYNReo
VaLCo99VIFitO+7aL0mSR8WoLW00xjb5d1Rr6DFgUI1fcnFXnWIQr2znmW6HhGyg
gmQo9XCjDlVvTYhU+4Y3d2GGOScRFWQgYDNsd5lzJRAPyNnvZW586rRjoG4RS7gO
Qzpv2V6eRtH/FEs5tK5kb+VRG/kUF+FmtyMKGw6O1LewYksMjoqH23/DggpDzo2p
fUseyCikGf9lVtFtbIYFL3QtdspGFVY+A/ro++5koMLj4qm6lyOR3m2TrO1IKJ8B
9JLe5ZWjoRLPJi35J21D6To6O75ASCdHoGDsMRAixuzHq/+9CZTRMXm1Vc90DEo/
EFP4xFdErdJvxSJaNSvvIGOYhdc/+pvv6gE2UDFfHjnoMfMZMimDvIxgTrfC9ujB
B/L3I6JAVwE88g5L0u+NA5DFRBmiXAPZdi0THq+6WWzzAqbmukdXQD53OGcEUzAU
wtY9a57QS8UKJRQ8GcOHxvTBmcJKAA8EGBIgaYBoyD5XOL1jsgiGTD2/WVXlalhh
acVfjHoNBxhrmaIxJsfbQqpTk0HNBJha2aW5wcKW1bPYj41mGaHOPIkKHRLcnIZ/
a2/HSdYNOjiWx5unJt97o+Eh8wPKPyO59puXcxTbH63ceWAn8IGRuTTxz5z+ynFB
oha430vMHjp/klwKRyQ5sgL/LPluREdd5ajFFwMlX34ce1MVIMVSGKmlpXa86bNh
xrwk9HHdHrbt5OeLFTewS+BLXde/nnwmwFAsEBWIdBVGf+IuxScFma1DIBMr7eRP
qIC6/yB+a5Y8/iPLQULIV4156MFedONsGXuOhtLuXi+TJVyLW2MVEcadNZKmwKJG
1Qgl68ce2wh+lpokyCR+3PIewDMPxGLrthfsQA4NAzYl5dPa+cRYFkgDgt5ZreKU
nGmpT5yjuF8NdyHAQM4XMQfJS1RW+KGJhcCajr2XM1QUL3IzsY0/4dydJqIWdcWZ
IxmXA89mKupzi3wMSLgSZltr8KLx6EE6+Xo12gStkZY++Nbb4EmnpHBA60QqZAGk
oQ7TJeMsKgDapqrAC3VgmK9cIkmdVYl3QI9ELP1YDXLW+WN89zfxFF9UiEdFaVA6
m7IKeyAv8OJYybeaNLNAxgsrP5rQIPRlNYoRO/E0+NyO2xGo6UiNJCxItKEWRMnN
KCAdT+1RvdBUjHqtWWS1E1MTQEI/hmYvadMgl5jP07I=
`protect END_PROTECTED
