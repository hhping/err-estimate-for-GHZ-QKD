`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6YgYL8+DwU6pw6vwQCwzcUtDfpzutTSknXaNi5TmYvAnbW8p4a5aqB5XYmpguPWm
05VxJp0WfBJq8PgyTaQItyK2pH8Mb6fJjphSiKJdWKebbpS5lCe/O/oMacVs0Di8
DZdHwM2wJdpISYnS95EpOAWPZUqq3LV8H5x1WlAY2F0Clh6JyDEx/jVDkNzcQXOY
GonQMP/5WCz/REjtdLuiUH4JxjgOeTnXSxWsMcPUtCBjy3TpMLtcmeS3bBzt6b43
YWfgYzxvXc8QH/pIXOhQMqkV+7noa/3C/7lL7KA+Y3E1xmrvlNpYV+R+jULrWPRj
MhlcXxepw4d8RR016Y1kll0af61SuK8+JwoUwROXhx/uXHrA0C/pP2iFHYmeKrZ1
q11pO9rJzc0TKx07M8IOGBQTvtgC7LurAPPDJ8kFjE8nomKUT1XQxq7ynTdqePPB
jgOpu7Nv0hpCQrbd1HbJur6w7BSt+2bipGCGrLv69A8axajAd+GHq0qBeKzlkkA6
mT6QDibYghSYbRqNjYsIlKZ2kipcC0IJcol/Kk0Mj7Y=
`protect END_PROTECTED
