`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y6dZY4AIBKihSVyGOt5Vx4YlKN5hcfT/+J5dsTBZpSlCxN02nA4bpCAraxB7B1/6
PvzJQemRYCLRT9y8wA0OmNlhWxxsjAbvbigiJovI/1mn8ge6FcSToLJbHXs5aSKI
PvJxgOqMAxx5sNO8Cob/9B43OC9HsL1EybXUMzjTjICC/o5CaqXxSpHiIglRL+5Z
lgHWoiim67Trllqbzq9scR660Ot4DrqPXumdpQOENFhYPos7ansBn3qG6Vkx6NL6
bXOJxTic05/fQ6TgH1rHWrIZTxOPzdG3jw6lfamrrLkO6D2smo1hewf3Fa+0qopM
Tjw7dp5dccDuTStheHyconhswS6nmWsY8GsKTwhgNtTt9yNl7cssCywkqeOgQGO9
Y6OKIBUr82JpvTZlGD/Ce7M9qk76PAlYKeNkPbNFu66VL7DU/v6/ynYzb+6ybBCI
AFox2gm8KyCpj3fZt1df4WT/LTeN5kCFuXZerxkRvPN8tKXA7SBa2zMLmNLYqEKZ
`protect END_PROTECTED
