`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2dU0Q7dM41BxoFIrXv1d7KPZVKNSfe3+qR12yYikrqmpg1f895FKObHzWIszgl2s
A03Hh/ANHjN3bjxDZLhAiCPEi2lXQl8EHVTl3tDJi/gBo6RNX2cmyo3jQNizZLRs
PGB2+l7v/2UJQnT+hC9ny/nt5O5iIsGD21vmB1ZBP8auwu9VfJ0EifpFoXY/z6Uj
lPRXtonJ1R0T7pBsp4+j4MjArTKSe65ekYhjpV3LWU/UkEvJXsa2QGAi2LLW5m2S
BRLX69pyBdL8KaDmfzfBs7j/fr+P9Q2OSNBz4tXj2831paAYhjnQuyyfTTnjXwhP
0n2XpFHpPHfVAOciKtitaMZ7uplo+fBFicxV6DyXaS3wjkOtpsq0sZVSmxlASlN8
vjONJKYrIkbla+pQ++cR2pgtPfSvvF3aUhE3yEPWZtT8g13dtN5zrCrKa3K9UhYN
FQkMZTbkzFZH5F5oQCkzdhc9cVdDMsC/LcPPeQZApsqjb2U+wI0xV+S3C3Vaj4tq
UqiPBhsgT/slpt37ymrWNNdGzJfPSe0Hfv0abGyB7CESvpEtscrXo6wagyzQQbaa
G1Unuzjug81BeB+62/oJn7MOSM6/Em3GZydZSS6RvAf/g0MlPxWIovjLCG4g5p0R
wc+NpOSlvhotLqMi3TqtLUm52ndS2MZShAYS8A/nSHLA6dl3II8pomALpITpqyml
uevBYZiYxZEy5qruRDsLPX9T/liCmVMYgViWyors5N/7LWAp95hlpGhRdNWyWHQK
rV9qKLB49N7Zt/j9EQGuTw7mTIGSvInXFgmtU6kcq8DuMQ6lnxWjKmvKjUk0DI7V
vah4/7squNx/hLQ+up51N1hetTdjTnz/L1Fo51xraMoslSyqBGQe2GEJDR9P8xvb
IvHMrdj3dadhxAKKhcxdeCvzflwMX3jLiLi8khqDcjTt7cAHEoxMNTLwNMhvofUK
PlSbLKBx6vhKIE1lUCcJQy0W3y/oZm8wwQz46tlKXohYNYKv2pqKyRjvNtt4PFCm
sdFSA8Oq91dNJ4RJF6WkdrApwd04NsLRTN69NFkz0u4YQfUPCSAYbTnWmKZPyb97
b98EzbZc73gJPCIUAmbyYsKar7/Q8VjZpFdYgrZ1FU2rGH46adnbX1HxDt3Zv1Dc
CG42STz7lvFeOvFg+Bbkk/syQ2aqcneFEPzv0NKdy0G78pt2u8A58jnBkSHXuSVk
hBcOZzclCT3DSSFY161cZUbdLCp99ck/nuec8j76IQakzZIp7Z3D18otxydhspAf
HD5CbqWZYvhwk8Hq0NAo8lSI0zZGn6EYHTF4ArRiNjgrTowoTmikLYVwv0tsob/K
j8xoVCYo073BMXLRFCuZSxA0TsqBiZcb626vUxEovX0xjP+1+mEEm33PzDKMuly6
yXEFSzWF7p8ZC1LQLJjcUM1gbtYlKm5xc/Q1e8/ZuQAgVY7CTgTOD/hztWL50siQ
Twh83iwHSqUkevcgALk1shVjlsg/hR4tyEqCOHKyN1pjctRMtw30hjPFniT1f93r
lIwCIxuIMc7VrQbSirIXw2N44gFMPmBeyPMkxlFpXzSqYoqWecNKdRWAvcP4ABOz
dnv7b+vv+w5jnSHGv10X1YPcehugz3wvBw/zYtEaFRhn0ZEeLMjC/FwjHJIMHu6G
xBlQE7k+baVCFudfe1ADGUuZQZw91LSXL7u6ZV4R9/TZOe/lcSJlK/yLlzBiAJ9Y
0CO/vl/NhKZblfXIpRdk1O16FQUI+QpsL8+4nSQZtfRk8jwml1QmRc3EI9Z1InDc
JNW1+4j5+INRPlsyYc0J0MuvZ9VVyi0Z0z+Iek6bM2cbI+XSPgd0grxmxvo5jAPs
tK4+wVF277szMZnVfYf1PnacRkCoVvFS3tfZb8AzfDTCyE471bjvjzBVZ6U9Buye
QLDHhtuCN81yZDj4qbT/W9C0StJj1y1+eSNuVfwnDIc=
`protect END_PROTECTED
