`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fVo4nsqEAJtpamzxLfjyYGp1QfaWW6Wx/HHu5jWs6acCQ3uut/zug+muMlnK9OIc
Q5yhwWCgIj/irEhkXJLr+dgIVaI94NIvswIKVmV05tojdOeduR5a+oD9rzRZG3lS
wm5gpzi41iFSMUQHdL9Sjd8BqY6UoHYhORjJrM25x1xS/WdjQS5TAw08wcCgoFh/
NPutLEGPML3qB6Id/As23cK0gNicHhcSvl/SXY75Ml9uAX7bT0sjrtvaU3ubVrak
ChiBx+6g0yd9TTHDNcsqy43tnmethQt2iU7NqaLHotW2xurYFp1NbwYjbr58qTjF
WMUWJEyWlYkWBaAuyraUyfNbPJDvE3O1rUoZnnqXO2yNkc1ldF863xpPUkag3vel
C7TxRMFTEhgttvlNycv8IzehLa6jCytrsbPuafje282OScChhrw4L68VD3hIjaYx
pWRlH38QHSCu3gULtOfDp9/kaH/P8f3wJJeiZCu2q+6qFRX/Ugxz4ZFdJ+iqFTG2
o5JHaWtkDJht6NqNfiht0g/6nTOspOGF6ntCQORlDhzhiHuKU59G5B9WYAuQL2ff
SwMYnsCTQlI8KdtcJf6d2cMAQUcFE/Cw3HsJwos745G+KcQlYDe6g/nSdQxyx2oC
yj5kz2pc8YvL3bA4iolgS2hBYm99+3Sxs1utXloiEV21nkAjdFt8OveQ+96wYGpY
B1c7apAyYmChDgFiOfln835571WjpuWbC69P382Bv++nbGQhgVxLj6ZplssNucIn
TOea0Z1DkTTc7FajlHxRA1qnQpxQjN2gjbr+a3wrS5w2N4yAhc6EAr+XzGxThjbG
N4Y7vV2Dt43wUQ4V5BoOEP30Vi854RByaE76YacN08N0DXbkOv+ntVMrqKPsZw6v
h6kZ05+gG9002gccuorAwDCYoLR5s7PmRUstbM3mFdsKAobHaWJQo5L/TSOcCV2W
KHXYmezIKHmoIiQA6yA5Hm9gyG/Rnh6kV7ELolSrg/650p9/LzBwUbgVakmG+vGO
Tu8a4fFcaBU+5WYs6JzZUxEKTpTepr5lwkVT+dOLrd1CI4eAPoZH+J0KGcxqBg+Y
utpsXMDjubilei7nmx6reeZLj1yXt07MGbQq0fRMRhK6KoSE0rEapU7bADonDa5N
KPTlCGOSM4eW39CzMtAZx7Ej6lVeffQhywk39pPj0xdrvBVRye8wExvOQmSSEJjH
ENkGHqBCEKM5pyZagByk9di8nxGHO6PJvJTTpW9g3KY2sGVsPDthnEzV8c5xHbW6
AHAWLCJhBSV1jVSE41ukfnftcoZfKIt/cwCNkVydyeuo6bMQVVcnuQhqiJrjDDIJ
LB4pCbLGAHScFBIKb/83f6+RU/drGCHGXV2oL84cPA70kNx0GDTCLgPjdpkZRG9j
s75DS2W2MC75dhFlJQDG0Yl+dgOiztHLlYiJCIpdec7dtooPzHmpvkVuibd9OV/n
baxNJzyxDk1nbnngRwcd0q7Is306BgrcB6Oo6H/ZDVcssQl0S1yyYkRCVNDM/sSa
tj12DBnsizwUtD90WG+KIy7uAKUQ6OoDyR1jsAjwuE7g7pbysx3AcX1gHzGw9i4a
nJMLO4sfosnL7sdU5isLj4aTSjNaWLkFOEyildTlRpZldzWFzd12KDBK8m8M9GoN
wTW5yJBstB4LXpqSWNH7g+fcyEwDcbJszTyaHW2qh9bVVzQ1pDxfNP/vgr1hx1KC
CalEYvGSM16Ri6Q1ZfV8mVITsbmXbaXMu8dan2QSp1m9w8b2x90VGda6WnvNK3X4
+On0AYMZ8V9EIDTwHTO/6oi3SX2iKmB2omxB+JkMOqywG1L/axGcfv3FFzdrhF/8
l8gIaB8XFS7Iq3VtK2SJCwA2ykQgsrqLp/6Z+1+xleRJySdJcALEyRBd7fGDf5Qn
2kxJ4PgkjOxOo37cdU8pH8CMTN3fHo01w76UPxdEo6U=
`protect END_PROTECTED
