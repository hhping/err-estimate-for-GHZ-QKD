`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KZyIIxy0sDz/gVSqOjopOSLhVp0olassrag6ijJ4z5DEadN0XZbbUg0BDXMz3SFc
pyvzuTe4oblBwJvR4oL5Bf9+Jw8dp0u7j0FXukj0EyVDrbCN+w91ok/QjZz/gbuG
gDvDFuWoLuJBWJFTYi7t0ELA31sQnf/GN5kgVGtLfzO/QPN02jAziu+TzwvVLZbo
asQ4vFdybbl/VCC/ho3xgntIVyrp5ffMCsR3FICPT47HuIn/WIwf6jCsgwM2n8fU
6W+R5gpBAHWV5JRCxhIOd1LoV0j08RTt0jQqNds87Mt2HyAEoYgm6qmhZ62HPqlV
lZaWTrF5Hetata3S8C70Q4IzaboxQ2XvI75eWRWExGqPwdbC9fxtve5ucWgjB+6l
w3p7JJkfCsfMX/VIavYDKhdJfceo0YJFim5dD3rCJmwpwCgHJghWbV8uzizRSmmt
uEErcLUxiGOA/9LLsoTnxZn61e05B/jTtOzj+iHVSpOLeIadRDEf1WCGlt9KS2wX
o8TJyoHp93LUEtGef3v0BkZvVaTciMbJsMQhDu3YudwW9oUPWXqXbz4owZcog1vZ
DdXBVHS3x14ahbay6FGs4qSVCO4h4+1Qc/31+ZB5Jq1EZpxY0gIh2C8hUPXxC9QC
4ZcmzSpRCuly3pkqmIRtm5w2FoNwAqOU7sYmUNH7A5wlavzC3UZFTJ7OPD/Re8cm
7cXAoV1MIlRj0fOJVjvxmHUvqzBdu6OHNqOXPWcWCllTbFQxxCC4V322vMsCRHoT
iMfmoYLcGAcNiyWzTVpCJPtIrW2j16OL7KvnF8r7a/OzoYHa6gK7QvxJpoRm2GR1
NZj9/AbT0weBWv8733vdbDrMsrM0EouETdhtB7IBqqN3XEmKL1S7KezfWGEZeWcj
QC6soXqfVoFiUvDN0HZuM9/BI6Q/M7F77d295HcqbGOXL85hOTQkaR5UmB9iqYGg
PExA2m2Hjr+rqJ7v+NGB1/oOPCD6TWM7aDvhjabV+KfuWBhUCF5qGlfLSsDxstSy
8iW3Ntnf5OtxeYmp0cH+a9FlaGEwdPEIYl8EfYf3GMWIvCYh0lz4uKxsCTkO3AGD
gdXO7IDLJJWR9G2fUOF+SZkEJ8aN3UojIcHC/xn4ixoxoqpRgveByL0kZSpnSWSw
Esb9RZbXT9VXeu1+eR/2ZAfJDSmHUJhliesC11TBibQnSMIRbD64XDXx92aHMvmK
/JLgVznrOkAHkoS7JpaWJZvUjWPr90hom1o68mAi9SVQFrTJUhOgdkTfUm5rztV7
DcbLx0MktODQx++OZiRfL0aKH5bAPffeEY1EXCzNc/NY/C8XZz5oVFuusH3Ty25t
9nArSrU3HkYvE3izjbs2Cbla1jMYgiRI6dqDOQ5M7fKAnHyX+Zu3XbN5/lSh/W6F
wQHssX38Ybcdk98mAnReX5z66Aook0ti12kgzsQpbfcUQvHF+fiRmEiKtDdriwxB
qzs+LGUnV87mlC2aek1o03HaBmfGpqYPzWR0+T0AhDHycC+/fzs7O8HUSQirTDsG
xY0IXksgI0ItgNH203sou3ne93+N5GY3v2fsZkafz9D/l/mwI8Y3+gcH4Gu3Qn4A
6csYPfidG4MEsDbaVK+B4bq2F2XD+Y/+sRhpyEq9wtpBlcuRJlVBTFAUum52isP4
0gma3q92/srC/osX0DocNvFkWI4bLLjXB6Oq7loeU2KjzVP8IyUPjBdlDEyHuFAn
30ti0UyfnA0HBpozZG3oP5nuEasOzVnT1k23T5dQhQ9IxDosZAAZAFOOxJAcLXa5
MTZV8eV9N7eHU9PxpjDV9fCRQf8VnhTo/Hp+y3DYX396IEH6aoWjm9IwRVXga3wb
zD2hA3JTyDcOF1EAOgblHsdtsbYGIvgsRDyz2LVmLKEJYeY5fP1dXf9QIAL1mdaI
iNlbDRW0HEsoJIIDcJPjCK/v6EwLHMvknv6sAgbwEOjAnmPUqz5zX62XIcgEPYfC
IVPyNiGvbsE2egtqLvB1VdSUdaQ/zrXnIaDZ/L0ty+7OeJZL8ZwDzU/njeg3uM52
b/5H7hHBlsm3HTVTRmh7cVOU8kvFojD1TpxZjBkosDijqM7fw9JoZcgH3aKCsuhO
BGw0jfxTARVObYpQ3ZTTqA==
`protect END_PROTECTED
