`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B70ON0321fwYHjs8egCzT5LdBOfZ2LVQtJfmXyV+9sGrUyzHnUwtklHh9p/pPlMM
2zwdTLWwvfRQZbv7JWgraNElnFyMPhjkdqomgMnpgFmHTV7n7mNXJGHStrsm0Q4p
1WZlalm5Ns0LflzcxePJ9d7qIE8BXVBrY1U/g5SszW1hZ0oG1T+2Y338C3rEURHK
sjVo5yhdc76JZfdEZrLEMpw5tcLlo0VIJwFrq+TdInjv52hpUe+X2R8roCz63SH1
S3a3bINZSsDxiMSVefOCjonu/pZb6DcD+jnJTRcYMyzKO915MR6pCSsuqAt0lPPp
2guZd7QzPtfzbMKM0y0pax1UfPUTrIrErpdnUrlF20sHM4vcwc8HoB7ZaAizOchW
7C6G+PJMJo7OxN6ynxY2/WF/sDzdW0aYldOiY9vQZSYe7AuGiog6kjdvv6LJCIdl
N0uvEgLh+/LVBhj24bHq9YPmcenr3/gIb1jpgZHVY1zWF7ppvqRTXciO+KmnCWkf
qUzGjub5sen6XOwGpWuDL//9VFraMmdhyf4gppxRSvWIENuvg8EeElfBdBcu/24J
8DDXiGApPYKLzemUmrXdIZ+1jyNZ38RwJEtHuWlp9gQkN71b3pcuqOzINdjOnD59
T0lYNMF9cRI+c9n1hHVJj79P6jV9IG10PVJPblJ+ahx6Q2pYPut2RG7PSctlky3A
sF3MR8IXv/TvYm+nIAd1DkA8NZx51i/H/kH6ZFGhtxMY+bPy4Ojk8B9jUzeJ7fel
uDp/kAC/FR9BN7G/m7m+Dh24lH+vwipOH+nFMAg6IkIa7cPpaE8eULp1EVlHLkH5
Z6+1CyHgiJlNSNbAAhFB1LO11YNv/hnef7PMEaGn7yfr7tA6UkGKhkTJjyax2ADv
/ESwr95KrqHEHYi/bYWh0Q==
`protect END_PROTECTED
