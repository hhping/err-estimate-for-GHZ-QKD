`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EtT0ONj0hO3U7ZR1ky5Fw4dsVTn3Fjc9TNl+GVw/YZf5rmO+Y77aPScgHCcLcNuE
mA86TbSD06CaFqYMXn6UzDlZJTDXOnYTRojiMITPK8h8jQyxyl+GKCLbYKrVtAU5
Iu3nY9uBazgkBuKGOOaEubrcar5TxIfwIBvePjjsTqS9mnDeXhk74ktudnlSsBJd
RN0NE09pdMqLQzWSqmIWBMwG0gg8oRvnBTYxognVqavaINBNgrTzyJMSxQFN+oCT
eTi6LiLSCLOAG1mpdZo66kCmCj2Zx5OltS+5oyBZ5ju4WzgAHpX7d2tCBFjIz50W
WnpneKEC6ZwuQ8JK0inJc3URj0BLD7CO5Iv4KqeZesGj37iAe4QepX0uc+tBJs8o
LFTULqLQdpL8nEQl3gsbOtEh/w2ZaZXjsZ7AKc0j54y3yvy0LpxX7jw/WhOZGbS/
28OI4p844d+7tsKXoVI4sN4DSvZp9rQTDjsbFzEgSBjfo9tvSS3dt/w1iquG6V1l
x5opZ79MK0ci00us86lGgYKIj3aWVeHcXdvpvfh1C3qKAILyJYVXpLUpPYGZ6ZWQ
a44IMw0iA20hJKVFskI50T0b9DJSWSgb6rSoDZ5+g/+1gh68lg9AvYucOnmhQkoq
Ptvst1SJ65xQe+rXJmHedwfH4kzm0qPzE26UXRdmJEIW2Kvb0jD8xEui2WCG3ARr
O44HtG4pYLN38nfLBz1htc/pyrU/kLjrOVz5eHuC2Z68mu1cstOOdnVutG4NpqWb
iY67rqRNnE45QAXk5aYMUGxngm/0mcR7X1mwgHdg16M/F40xEnOA9HFX7mHARFWi
bW366TEbEP61Y0x2DROJJJ8YqGrmkLvLV8FjTFmvGJyUcaKD+eu2vacUPg3ninj7
Cz+LgcqioGUM5IfxkgS9HWbiZGgNfMjO8/yuFiJvKNvGBKyvhT62Mut1Ny/vg12L
3acWl86dklO60KXr8gv4mv4JlKLRXSQsVkLX6i9Z9TutixhMx8sK0uMLekMl2wHu
qzdWeA341wnzynKMV/pioQ==
`protect END_PROTECTED
