`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CN1kVv5sVtsq6tehfK+6e8V1VEjkIagLRScZNDZCVS4bu1tSco3MmM32jl2qoW5Q
oLXyElfha9SVIHxgQSMRw2OVXbIlNKJ01fsN5WwQ0f1ae7xb2cg9iJ4Mxwryvdej
pq1AZBn5W8VOE6yLZdmwfdq4G7TwlMlGgHU23IB/bVD66LuRCfYOyNEPHSaMQagM
g8+95zmLmj3Z9oB6emGmztDoR4YuqIzXLaGKvlbGt1tmYoaqOSTR6tv9obTJ45G5
f1j8SQx9qBXonhsGzlFjWcEKmTVrHqEGob2Hc6+B/hYY95vMd3Dd+qj81IZuNcOW
dCuSd5p7MSOQTF83CayBKdpEC3F5QEH7icfWJMXC505m7tCXLxihYmYLNdvpMqKj
Gb3NBnmoLvW1HJT1V3Nb1f9Jh5gBzw+X3/D7RxY2mbGXqsCBhEid3or595GvbRp6
luLms6xoCqPD2ouNy27Vt7z1NweOiQ1TOg7VmGU3JQUroN7HLYxCZSYdIJHnLux2
wos5uhk6iBGLRSLrsGoLLT1x+4F/4Bo8PlwS6Vw5DXRlz9Wd/bcnzsDj926LbWvY
77hoKzI2lsiHagBLiZbk3T4bAFeOWfC0B/lrmSlOxyqt32LCrXZM/0tARImopLQM
yg/2n4XCuVlutcPP4Rk5hAQikLaYLlu/LO6vXFi3Rs/zgjA7kKCJe5xuLYhHndYU
TqIbZ+T/UTBHpFhTCnFlEbG9+NV2dKGhnQyd9wjnHeA2su70obvqQyaTJLy3w/D6
CMI2hiIkTB2AlOi3CNAVJQOo2parAN8zKeZWu1hrZzg/mkClewXsbJJFWZEY13tx
ktDphddyXw7lPozDbj9/hz4+8msHIrfNMZ80TAEogPhHEelzcu9iH4WWQ/VSU/O6
eol6RampbnP0vV86ty/ny5UOS+c1kGDWyYsnreFcJQMLGtiLvKND+U9xVMmnXZLe
GQ7D8pWUhoGisN7eZqBelPi8HMhuogDUx9e4EHSfMBxTrPGZtVQEPZoS3goEta20
jPL3EeeEfDzpf48VnpUkRRUzcNlS+Nk6fJwbPg1azeM=
`protect END_PROTECTED
