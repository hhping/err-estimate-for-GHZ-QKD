`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/waSz56MoXNal5iGS7ESv9lpHN+7FpL4B914IE2aHDINDbCbBTI2fwJKzIufPl02
O3SVSPHoxRP51U0aDGBStdyIiTr/Mdiu/NDzlCIcAgIwZf+D18GnproOvD/FV0/i
Z39aaT2NPcg3nbhnX990LVK+CrHVG6L9TwduPL4I/GZ2kcEPg424dnTSbwTbRT0+
EnF13UUOS3eW43NgmNeLjZ+tUZWqtQBDBg07SkwXq1KMoz+NhRUGSRMCqsA8wUkz
AJy3cwhIYD9SWgkKHVQw4h4tnJleHEYyow0DNId77WqKZOOV4GsLr0zi8uaHj3PL
Zs/ibM/6sJko9NyrJpaw1n4LyaU8wsYp+ezVGIGRm88xm6iRfkIFzirORPLweCAa
sQqcskCmVfq0R51f662QSz1g0ePyIu9rBZ4CoOBceIq1e80ysITTHl7141p5D/4L
1CR+PjtapmWO30dshorezgeVSVrbnfUpmOfo5Ifo9NhRr2DK5r0yJNc0fb+Q6/J/
bZ+vAzVE0fRIk0asQb/PpTnh/4MmyGgoFN+v2Bt44cahSGR3GpmPicOfgvpntEWN
eDqEmL9g+KAkges2Yq8ZoYgjbbagWnCIn6SLVsaj4aC0RXFuy4zxMv/vSVN2Ldtj
XN3JFhWUZULCzJgE7xWf1JzHTQ7ULNNdRaHvvVQwu14=
`protect END_PROTECTED
