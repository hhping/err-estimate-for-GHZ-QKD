`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GdPEsSOa5QROOwTFizkdI3q1Zojrm9xUzX/F0KoqyXOphtTIylNEvSphzaEJslwZ
z+d1FJtuGVAQ7Iap6kxcAVIG8BYjENeVIreH8Vc1suvL7QfAnA5+Su7nWpa98sFJ
qpKMYArrw11p6wyWTBFw0/sb1rnFZrGePwD+5kCm3WWMhdiIIBRq/1EGDus7x3Jv
uP4ueP9CleCsjhLkfpKE8Y/pkCfMvI/H8hcyiloLxO/9ZkAz3mgJocwbG6F/azz4
lQbBfpy/C9yfY+qpMh0B+hJMjeM2uw1tv5sCpKoqroDJ/HevBJS+aFY3ie2wq7wm
ax5g1yEsVwSFcql33nnEnVyT5MQsRWTqp0WzDh7lstAZhJYzY1e4BrTCpt8YgkNA
Cwa5reigdgymF4luDuytJg8JEwYDFdaPgTatQfA7MbMYgcfpzrsPy2lypNDMuYMc
+cgKrbqO99UjOYmqt0xeUWDpXEeW1ywhy4GuAEOxCrbvE8epuY1PfFn/GODkQMta
di+guUzWClbz/+/0yggJVYbgV+RBbwtDdnuOX1YKqTVyHbFuYo+3h5MO1fhILc4V
+whNv4/uViYjBELf3Kd/aa+B2EtsHVgO11YipXJ6ECzWj702Y+hM/0Aav95iW3gH
6+5Qw9bsiwhICdAgX2vYfuUHcQqAnVmXOl9mvUo9c56MjUWlivYpHy4R9Hq0/RKq
jGxIj/kA9LiN3EK29M9mRXs3U7Hc1yTeASj0J+gwWm8n7GYbQiZAajIEubHudWkk
NFYvDLJTASbcGazfdrXv4/eYYHM26/iDnVITxG848Bb3ceH7UemJekJQvtnGVlbV
OLw6k3NWwiLCC7MYTE24Pk+R6FNmybsMWJPg39nJB4EUICFyfmpzMUKKWmoy5aTl
uZyx319XvJR/4de6wWeK2GQo8WdDHUxBsc2qud57szvc1djh+nKo6pV+EYCuaxPo
pcPShhS1wPjg94ysMERTxbMuPR42TC6ciuCL3QKoTDfTt+jsdWeFgpC8/bVmRbbk
t8SwynoqiGwarmCNLuaD8MkEDWTaXd3XHH0jbZlE0w4FMh3Rgc8NsT36V3HGnWHR
oTZI5mre8m2kIVKat5/9hOnc8xzKgMbZwuEw0T1smR6F+pHbE82WrrdYMIQLgPGt
`protect END_PROTECTED
