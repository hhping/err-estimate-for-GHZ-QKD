`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z9cIelMKwkIDmhml3KBYS7+JVDKxSmcueVM2ocYOOUeE2ArD1A7+JHsHZuUZc4Kg
0ofzjI5g7cUQ0kvxdMS5XLRhVWZegS3+KOeTxbSKokXrnEeWPHd3TTGcGRV2MGJx
ZUcG29ZVuXrBcJnItkhkIjy5+o+EV6Nq74FVMLcTxrKzp/srsFs6IlNX1e0ZfcEl
nhGVxJSsLVMAa6ZiDBcVe4xV1zgdVDYDDBh/F2SNAJk5TZAmyj+3MAlsQUpj/myv
72Kwj+Vfu9uSAIhrQbXhCE3QM/7pFcakmiynyX/znjVoYTKKmI6Eots7QnjMH8mT
J42nhIb8eAZDLESFoploqtswl3eBf8Ns2tbSU6w1JooxtfMqFC49JBjhtjF+mA+V
nCnmtosVbYQYQadt8C7olbAYd70oFo3NV4nB8tFGlmrCSoGi8/Udmh1+uu5k9WqV
iJesoSKKrGIFcWLCipJKURntrv/v8ePfTLCazf4AOEN3dkoRMkjoj0pFx2OZrTQ/
DiED73Q3IZodrcHlN7pJf4z2FbuXeAVRcKy3dd6f8zbB7nDkJzSHLVseA5/zhkM1
ZOhTaUvrabGIVASZFU/EIWQs2ts0BEhsrgGpnVGnECdbgkJuJKLWYCaG5PIwO0Zq
+x1wHnwlcFDauvPCGk3G/9TkLO73pkqS44Tlr7keSvtN/VR7UTdHmNPUng0qopfq
wFiq0D34eYaH9R81LmBu4lEEKTai8VsbMT8KVqDRA5bHSC92AhVar4XDcIMBevFb
kTqfrcJzj0nunAX14BTvyeIfILpf7vW5FO21A8Ald5t3I5g3LShxZf6TwHr5FWE9
pwJNOpQlLKCLiXgKciuMoamNRfU/u6MnAj/REEJ+92kA55TcsqFz9WliD7Ge43dR
X/E8Mzwvqd8sUZuEhM4mCwMHuGuHk0GOGDy8/gjKlZY=
`protect END_PROTECTED
