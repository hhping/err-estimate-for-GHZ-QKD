`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7LigpxKdyp/cpvuMLaAnynncM+BK9Lt6KgQWHCssmxybSDJcUA1onUSvPMTdQpdd
9ti9ASOwgV1aV5JovO3XSOD1ZFyixaFRpjxUw2vdd4TNB9ycnfsodCn0aQSGq9Jm
o7zfijYI1rPCUVbd97Ce9zL4tpWQLBBDq4UT0pHSNtdY+WUDNO4PO2wwljhfX52x
2I6NIs3P9WNG/DeYhyr2M3+q8G3QPWhXVuZmW4EAuKNPiuHUy8LjtjKtT4eTDOGb
ACq+uz61XJRm0vKjwek1PSQZy3ylptowg8809vjlmMVwDOu+/jjtMlIKkRWLb1ir
yOuw2nzKtTKIpqWgoQ12C+w3KUrHrYnuttUrTA85lqnPq8Bd10uNvRNH74E2XKlr
35DDiMPaFE07RneJ+wple3kW1B3PuwiACY4gDRPYeG4YoJ7sjNrCz1AhBnPE3aNE
TuYCraVYFP7tv8TSatrR6kPfQ+QV8IxmN+dDPUcPb2EZaDIKsCBrF+oBSVn9vTNM
IEMXesbFPLDk9ng0i4rWXKqneLyqrbl/zduclddyiN3jYT3wlHxJ3WED3JTXa9Xg
uSf40/hY2v31D+UpRdEFHfmFJsl0YJt6gvOKa7tIXzbwuzgzZrAMvxH8qJaTv0Oe
QApbBG01ISQeDIqwzGkvK2SogR9QNzvQtGM71alaWaUb8oGJMIHtgHgegYIfNJoi
k+wguZBGHs0zRfaEcy2NDXWT4x0AgUeY/5G9wYV3AGynJTvlpxY1dQkcLy4Svy3A
6Um5tSqSsZTxxNj1z9MrRE4Z/72Biaq1T22euSRh1YQFjIgm2dCj3CWrCliqHgSJ
xj+GE+Le5wYdGXaB8bh5PX6dEtkHfW0gPHwA/izMzm8nzFt88m3fxHy4kKVEFVaT
03h9aPJBRWVdW9B0qQUvGa5EN5SiiVvmlBInuAvKxLad9zqde68iRkHWq42oZVtY
4xllIrUXk3FUPWHf+Vu068ECY0lezUW6yaLTduEhdzW/bvzS8fO4YwxM0FuMk8ZO
cBPTFNAHGkg6aha5kx0DglmLwxAOjCsqMe9uqXi+PLB6L6qSLrWCxEcZztqZNyYm
NlkCjXbn4XdYeow1GXBX/TtUKedEX0oDyMT80u/UKStQ3H9s+vhrPZNvWiD+IDsm
IECG/Jn2VYxYRUzQV6CoVZbUW2D1mvRLnhQ0w3cZU0Q+/w3MekX+UEuDuzycsj6N
G1hu95M+CKkvYBOg0rkzP0HI5hLkX7UeSzCYgPf9nDtMj330DbJTk74NmIHw0sJR
bmo8+BayUID8MQtbmbwWSZQItzWEsFJg4/2DB9m22GYiWdJFx7N8EU7qgD8qlGeI
TUsN5YI5odkJ04LZn5rzw4HxBTHDjY7+94N932O20/AjcHq0AELSAauf+U+N+cyS
lMpXdDBwCugyGanoQxh7ag==
`protect END_PROTECTED
