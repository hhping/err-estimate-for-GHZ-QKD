`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nxzyx+X1tKsBD3Hlb078gYdKyxhlKP2eYqQJVp5Vh1sRsL81UOOpJfYl9QXnTOcn
LvKrfD0Hkshaedx57xDjdo1WA7ibKeHGvonTwveZela9Xt7ThyGoP0O8+IRh5C85
P9KP3+1QYZhH3fdajqFSkd6j/KpBKKW9xq9fhJlfPB2FZYwvT0HSbpjA99oBT27A
OGR1qKB1952+PrGVo9HQ4XlFarTThxc+ZsOuXy/Na0fnb2C592pO0Hud4+a98W1z
9sFqDQmGUdFgGtBBUEkZYKee5jtARTOx243XDveoymlri/2M5rJuMBLpgxaVkgaL
EppG06jPwuojgy3yq01VfE9JEsccl0fV5D3Qf3r02r+gibAf1VRKcwkqCsoLJ0Jz
TAd6qYoKjablWi1MJRb/ixAzkEi/PZ4yxYRI8Vb8EOH1ZQrLc3wfwYawQQvK32Xx
L0J3rT+2YTXo4CBG0WpsBV18HqouRXNaa0qs9VO27FlQdTVd7TYorOy6DVVSka5b
NM4hPxxNadWbY1c2D5Om3lXffY7KK0V6p3NKRHCPwx4kIAseqjJLIWUcoQ65PFyI
qiT/5rjkvnW2xuGYt7MPJ5QfD6fhOZPN+SLAB1gAugszAVuZS7XZxWrbeD7uADXr
QVuDa0DDKtp9ea0+BcDawzfqpzhsoMlAp2IZu2YvG/Q9O4KBkLCB9DD/EuGekQ7k
vwiIRSEHtJEwn3/A+s/dDD4UwrBnGDWrq1ROG32HbKbvlZ2/3ax5KiU5cmyNxjGX
sjICxZzwZGh0ZLvxmw2gO4BYKfb28H+vDcO39giqe38ayzgUD/KPEQsouAzaVIZc
cgRBaoxUcDB2CuFrtZrJZQu0zbBpHdpOWDTd5HsLdKvjStrpnCJAuNCDr6MnXouC
/xG6s3mir2d2NWM3pHUDiELjDdXGSnAcnBLYH6eySDEGdVCOJ/a0KR0hcCmQzMI6
J+nfH2McZQYPXSRbV5ZbdrbZ1+pNwsxgqURsoq7+2Ss311CRdvoXyOnf1a20wb8G
2kRHdUGdxyads+y241rITy+UlVuvp/BHOr4kSrYvw7ZvW6M2i9yjHyC4vCJ0BGoK
sDIlE1AovgNMI5kWMjO7TQlpO2rL8APUjqIQVvPyqJjSyANrT4J/HRLG8KjQaHQ1
7wRAwOWZ90qVWUJjTrYbNsSB81+B/lPY2zX+smz3XsPvdsUFPtX0U4q882vuJhRO
Ag+NCeQMCyo3DYzhmjY6B9EGZZz7z1achvagXKYJmRlus4/8uTZKOCgTH/mpCp87
sbYXDIosAeYlnUYif8imHTzTwziYO7DOR/WHCpT118DKvbXUPXXiZAQ/5+GTwC4j
sPl8vCSFlJFqHGhxHF8HgJoShl4UqU0S+BInmpBvv81yhi2fjkd1hi2+u8aGDqiz
r+vzvx+6H15b+aaY96FvjrDuDX3xDkmO1X5tqvqr67yocJJ9H88kBtITd59zcGqJ
oFkkFHgpsvLCfFigpFPdGhBza97nhdHjtzewWL1IrlNt7tViXuoHtY+AdUddAlsE
dRKNChqpC0urXLMRwXZWQplF0ZWCBwwpbYUwFngy/cMD5pAbNeCIwlZtuWm54jaQ
RcgA8CvEE4XgkZyTWhkLv1qpHfT5fOJsNRZetPPTbt77O1DIoKfeoj+BrXObRcfg
nHQhuMpW7WqqjI3IIqEl53+PnSL6G5opge3OQufkcB0p20QCEpVuGMScMH8oqOWd
uO7qHgJZhRVxNto67O2Z1llhh5menASBW3TC0heNPFiNXFGgWrhP+Xcj5LemVoUC
xDV8MLtB4J2+kruz8XuKFmv/X9i49CSoKs0bShV3UEMp2+y3l3ANWyjD9+BJ7PD7
fXZi4Iqi8EsdIZm8MHO5wmpjQdHGchPo3L0/oVR8D8PyPTMMRhjJAEba0iUxDRx0
AO0+/X480oKy80ARfPuD7t0yZ7z5R8OVUxzPDB//BUZ0kUrzVv0j7yFKMRk7oz0d
4PSEjcryutTkSdazrDx/jH/LreA9uVOxRRAb2OagmL8SxIt5k+5ujZ20mu1IwveL
BHXVMH1rgZUSzUzNo1Qf9PAEX7JALRpP6BsAjdW7VjW8tbOo0vmgfmGLhxKUG+TH
5xcNAU2sk6AteComt7kYPZlgboOibfpgLHU9OYuDVc7IGXDFiwCCMG53zcyX0p9t
arn3Dt959co7GGqDgUeGlM997p2vXdnHF7/W/X5gTzg=
`protect END_PROTECTED
