`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UmeR7uhTkeQ6YoFD+DZG3MKygdQGQhjFsFrKYv+06ssurLcq0fobctkivSh/z9wO
EiPBr+nnP+bBUxPiIzTPk3gXYpfQAZlUAf68lk9nQGtVD9UyN7FhWXKKL5p9GWLu
m5SE4txXuQTBYJtGDuAhvV4Uj/yXKGc80Wi8RySdFlZz1tpAtC1x48jqL8OX3nqr
UdwIGOkKdajrbdjFYkHKOgPcGuV8RvKMXK6REU+ZddNkmPG7GXQD4f+YKfe5OZVB
LedCKfVZTIx2AI3zqT3ptp1AULWNGmO1OlIyqS8Crp2RMK/wa0EbWLYbCMNR4eMY
9m44ZvrZ8jcAsArS/Dqpe6rmAuO4PhTmJ038BUtAbFaiGHu2aH/Zk6NDtOU2AnhM
0zI4tkmBmLl9TJ6hlzmAcRfyPJg8b4HTOyqPPq18Skjq+EFwcDh2p0ZKjQkz1f9L
xZwZ2l9GqALxrzr0uAwhCGV4D+BnRGvLWVECnUuwuyVidaMjZdX3Zf2MaENQDXil
SLyS9m3OP6iusYhNKKexzuF5G/ZoFhRtDTUDJTHaFBJDRqmzs+68IBwtP4QaX+oQ
t8TOtxM9YzoaETMZbwhM+2VQB/sKSHABCfH3kuQQUSHZaayINTetdu27kS1N9noJ
ZTmXCN0uPW/Ye4LR0IzMz11iRSRiZDpGY/DPbslVajv08w6Z69c2mn2KaPoSi6mL
ooIDjJF0vDZ5eBWW0IOz0GpCgPlceg1RgSByG9MBOmr4DctrEnuReU7Ln3GTDRbM
yy4IFENmZUmCqgVHlwJbPdYfvy7tM5GxXEilsQKaizHJFjkjOLJO3Fbqhge0iJYm
xa59Q5zw81JXi/fgsq0Q/ZrbHjCUbzZ0uatpaIaDugLIsgIG/NaKI5s9ToPPafrh
gRK8PGr3soII6ALZSNk+aZsQkEpo5kIq0gEbvqy8/Jz5m2EhcqddtDydf8pVvLzy
3hh3w9hBtqzxlqPSwLtDaewknQT8nPIvDoGrJRGBjTF5IXUeJFcii0vDL+IpKv0D
zMwChgjXhJ1f7BuLQzEo5/yAVP2Fl12r5PfGx8urs17kMqH+WeDMvWdIFqnDrMD3
velFVuiCgVwULKymQoT/DjpjfmeGQqCsvQYj8iDyee/EbYdUEOIzsVQuz0mygc3T
`protect END_PROTECTED
