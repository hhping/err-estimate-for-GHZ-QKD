`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i4VXgd9Qases/SettWNKzIKUadgA12Cga6TGtE2grb0rsfzdt22Y45BbcrUC+Qqv
s2/8aHR1l99x5EUpaFoYa6Gg9HZiR6uKrBbVOJzb4t4LhISP5HG7zV20KQVpKfQi
6FVMSB24NsnBq104b7RL90Cho+OB0ryFMctGFBt0wdVcd74s+3D0nvmnT3XqW7ig
lCzeVgQhpmd0JgEMfyWzfL2GXCtob6vOzK1cfgnWSU1EhYN7osWxxuGRukxnCz5b
rlvt5iQUWIZZy5eLmlEfdl9jaaZxMeTxZ04S3SMnQXK8NhviEHXZwvUkBCYzyny/
t76n70NH+HW9BKJXv8KROpHAZh+i+jEJGwz0QF5atipWpLaMF1MUpkCB1XSaRkQn
nnUJl2PDdzYQhQ48auM1JeqL6wJ2fsulOWcBSbplx8FlwOiPxdVTGzUUIIgRuLHs
gKK5/xNGvhWR7eFKVrPycrqvo9VQoL4b+QjmEzQupEYUJX1qInbHSMQCWFI7K2QW
UAseILe4tJedeMubqe+RWqhwgJWIbnK2aK/H6ORFbB2T4QeodvDkfScZE0U44+Dl
2u/0iPb58NAX1KwrZNrQpkrJKAzK+TuOEUH31uXffULARNwRh1jTUhY3pwJiGY+q
V+zMErpd5X3xmtzRXRyCZbEuf+KQCFUnOjZik9Vw3IapzMyKzA5FcHTmoegMn0z4
at49p7wrKf4QlvDQ2tW0WKqDmU0MhboSca2MJjk/dKUalRglMzNGbLvnc9QGvfln
SrYEzaZwsHry4L9voiflcMGcIjTJWejCva9ds31ZbYwmjfYd/FK/5WzeL4A9gw+E
sokSv3SsmIIbkkvM0qAUXcCjHqJexFDNLjaIb+wTO+VfE6JiYFr+sDonPFReF7Kn
XCHY1/aaEtK74nc9+K7WvbCWN6h3Cf6xHDarF4VQKPBWKAtbyu3YDgEAwfqLJoVL
0h9XJUSfls0+6xYkMojP2XFjIJIbU3P0Dq1KFBAH23mkzhqspoy8vUWKXgqLP2mr
79lHplK3h01ZPr7QxojSKrFfGF+jG2sZeRHzGvqschT2T4va8nOJOLQZd+E+QOJ4
BkAKM70Q51PJoTLNxwX5Hljg4AYhLe7McGuFS1Khn5FMlWhX56P+pnS77bCnZssK
`protect END_PROTECTED
