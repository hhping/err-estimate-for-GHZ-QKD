`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OxjdfxNf/ADUD0IZ9MO0UgY0SEseAHDj+puvq08zv+Foa1wgNzbI/V8tSaz9foRd
PSXqdbHVxUHdkiAbjKvA/LJDmgZ2YtTtLMAMRhXU0B5sof7ga588dAWHUz5e++T9
hY1dfFXza/k3mAjmVk33oGhl8aXw83EogJxCepAwGSwNsGywOZNbyGfrR5mmzG9j
TRFNxSTqT0lTA4oK83NPwfv3wGmh4cf66dN4ixOb1jEO9T6G+N4Yb2VBdcUbKFxD
I6kIe5yBJqRLB6dLblf2CNxmucfwb/Fkw6pX5FBe93r3SCs+BtasUT9wGI426iRG
rvNU1OOXS8AL5kvXfWqCPXkhEt0Q5aHRkHEhGLrSRnIgi+l7pq7F6DPR1TS4HjGf
p7j4wE6xHrB6hAhXjQnGwKgHmv1rvrOGPb/bti5nf4gTkyTyh6ntz0b18X0DTkFd
iJsEZkEBNLHvNtGBFQQqjqdklcEJLoTi5Rqy6y83nxovgPg4fnbiFMe82YQbHbsQ
haMarhpvZ2JTY4/TQ5aKLw7m9fF7YZV3dTpV2xWr+0oRTrMimsIPH6tSm/F0h5yz
WbQhtqQ78dhxjVJvW6xlsBwBUxFHLx+L9s+TLr6NvUinu1XPr/UAln0WHTMep8kX
uXqaW7P9VJQFsUmKU2XZhhp9gYBfnAnP+BbuZiaBmPNI0s/ov0d0h2d/JmbsHaNg
kSSBpkBWIePjJ8S2nixj5EC5aTEuvnBSU4h1WQNpal5VsGZ9bSfydSrB3NDZzKDd
zHZCnLD1WqDX5YDHtEyfwgoB8rrwt9z6G3I9ObYC70lX+3xnR2ZMtjXMzrm5TW55
VCxFpqeokOCovAZ+2x9IWPVrxAXkrB7bapfGrVLK+D2Y2HjruQzevEdR9bafngXZ
hQbiGSgTtpXRiVQTgp/ongWZlqagzVDV0j1K/jvI0HEtfY0DFqicZmL5nD/WqLFF
3Lo0fCwLHQnTZ5oc0239tw==
`protect END_PROTECTED
