`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DzYjdjLCfeyGQKV9c8R/ttaUPCBv5kLCRqDow1v8qcNWUdrznfnMwa5UoP+oBZei
71jjgVmx4Et3Sa2WUcgiCaKYE6DnqwEkyGH3EARsbEjcUkON1vQWBf6GqyFAiXOA
9SuDQeHVqa7XJsKCPzYnGmGNzRFUoS8dbomH3+VisrRKBfG/wga9t4Ym7EEgCNWp
fQUDD6dY1trCIpMmpJtFoU2myh4sTEQXFmR6GzSTTwF7Pe7Ljk1f1UhLXgFjJ6Y9
75/7HShLNQyz6VM94KTIE9t+VtiHXeZxLdQMVt2ch93PCKRpJAHRZzPWaoTTnpaV
6qstzxwFzDzWjsaxwJdqeog7Ich838ht3buG2hWmV9WqVbKQ4Smf+qTi0VsaxW+g
RBktHs3qcKsRHA5HmkEjC1AI22HBGM6Wd4v2OYSDjfpIsVfI7fjCamm/gmSL5nOS
FJED53J70riJOQ7YQYxt4DmncHmtEB+KJReHFkh0OzkM5D9MgfBKiyJC34wdZoSn
+dOXr3+vgr/jbh1RIxKli9PdEzi0R8RUN2f9wrP4L4cGLUd7OENy61+/02QZ+u1G
9BQkvmFpUXZirw5KO3quj67q49XW8z7y7JytqaOC7qmE7nbdl3cNDWp7PMuZ7UTf
3o1TH9BXicBQYwAXXJ0ooBDw8hhSIyvSQ2Q9546IF1UVK9S8Olt6cPZ5SfyPYB9m
EQovD/9DEuklrJ6/Zuyh5cr6s1gJi4rSbj62D5aytMEuyMWGCc+giJIgn/AP9Z3p
apkCiYVv3r4bJT8lhdCj2kDBv1llCUIgLdhW3TXo3PEbym2Yi6wczpHAUl1iKVVY
UgWiqymXOVaS8nt31UJucLJk7Xr6uHZSGa0Nfw6VPXxnUPsLwbV4uBROoXepXGXn
4V/3x+CvDAOgVHQZoqkQ1GDkqIHJ4VVuTCYWruIfO3cyGmkQvP+N3pkYCtvY30Bk
Bf9tjb2mgwRUjshQvSMz0pXbkIdSKzb3SknwjbFcTn8jbNMUKU4VSrcvOV29mW4H
KUq2MqpaVUpgZFGzTMdbLWsGgMkvDo1l2Jqtffv961cUMqEsEzzWX5WRzc45JCGU
4qzYhdUwuh+Gg4apHeIGeWumxWXkOTWTFN9K359RGlhbB4+HMtMUiF56+8N2miHf
stE2xtkMwSo5OZsifI8wbFfmrj568G3c9I1SFwOZMVDvWQZiayrlEbTU1Yrz6EVD
lnqqVnUFRTXDrm8z6/tVrGeuumDwBO+FVHrEPETlRq/dlMmiHyBJGVAF4TVSocXV
COCrEEc16bGpIUczMUHjBh85F+d6lKBDxYN+4N2kt6U183bzKLXXv/ZemyZxRpoj
fhge5M005tzkrHJzdIGP7mT5AyeCf2XLfmn9ZfTn8cu0RV0HTzyrBVHY2t00EdP7
IMyPKIWU/UoeQl/D2MD6ppwxvJHgCMWto0gSID5UpH3CU9PgtiFxOk/GP5lrbzPC
E2kuKI2gSw4m+GPHloiOYQ==
`protect END_PROTECTED
