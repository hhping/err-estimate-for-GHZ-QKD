`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PI2/DrCZN1lgLkIQ+tn2YCyuHFn9J8yfB9XrVXLQBuQIdGvvXqIQDA8O9fECJQ2m
n+EtZ1B73BAt0JmNRAGJ2vYfKhaangz6I2QWiWyllGTvPWgfZxZEQhAKtd4GuJtB
EAMq5WKfXB4nNBWUCUNteoeRgxbXnDcunS/4oTOfJ523dlysIf9FGAQTp5F2honl
g9uTpFkHiAGmPPmxL4cbd5640ShUGJjWiVZCGnDQPQbGzEvGm2dSmQ0DZbdMAgbH
vJYHvuM32po5r8d4iiKQUOmR45FADxF7X/j8bjJdFY7KcfAEfuxDGY9CGGReblT9
k9Vl/KXHd8FHRC2xARFa/d+F+e5aUADkGTB+LWwICEwEkeLpkpMYloRhj006iNE+
GM2QkdOLU1+JPUmf1jJBLshIy5O8BnlAuWAYnrICcrzV6rsDR/2fqo/jPVzNp9et
XNDwBp7PQ8kSQnBthjYaSH2OCjtyYBFssgXBnujHQbbC9YXsrqHt6lue8VP78B88
86/2vnpKwX4Fn2pBT2Sme0eiVcUW8EHxBon4V1/T56OWwm/IvmkdwVE6hUmxVOHJ
ICcMsgdcxh/jbTfXlfWFScnt0zuMFpmhdWdloz2PU95Q23DOk77ugMKJukPSqj2N
4DK7uH6BiCoKMMt2mOgSFO7kSPYOAYBSQl76ZYYNt50ppPK3YGAvS0hSMKWJNyW+
9ZtGtqIAJ/B5QymEAWsC3o9QBzoWxsb0HjsQq/auyv7kTJe9Xo0FKt27QDgKugGD
H+lbJVKWVOZy3hdpTXOB997Rp5kzpbQOPVqBmqb9w6Uu/3wRhgtS58DDFHR1Y+7I
FMUFpZfaol+/+zttIeFmBP7JI4Gwhm5YtcNoJJIDDw+N+JWU//6ff5Av/qA6weiJ
VOOCG7fpE0+S04wjkeAfsCS82Mecas65rcbNxx+Siej94jJYnlkqLzfGU1sNlhIR
wMziIn+JQYq3CBklEosl/+cSs2ICZz++LydNOSTIblMBZybUH+On/yNqW6j+VSr6
+0BZKaN6bwSbnvY4myqcAY+Jv7AyfEhjGOk1sPBOCLHvDh1J/kVvXLugarCPamep
XN6OUp8CBKJ5/bWDCke3GylAiP7W3JNYa+YHTbSvoq99yZAom/7GgtcOIn2xUSN0
AV21wbXh4b52bUrFX41GqGnm9wtVmKouRavCSwlC/W4Y9hid56H4bxdSA8vpjkH5
LP1XXYT4gbCX3puhknaYzMN4fYat2RzizJEe7lowPiV6I6Va/XWn4/F5QKxVfyjU
kww7wPuj6AaFCuCEGwiRmh2qZZ7Caw3lixdOwaFoFEE=
`protect END_PROTECTED
