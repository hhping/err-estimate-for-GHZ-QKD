`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TBMRRJAB517606UUpHWvt1gvgMmtwVR3Q1fN/pYqweHLY1AWILXWy51l2qAC1rH4
Aq2VKaekizdyKkktYpj/pHwJCpT1CGL6BdVcWgEQAzy6xD2nVp8EOAY+v/xdCXt1
v2LgoG20/F3tLifQ04t7DOCmOBSTRZMeLaucQZ8+RrHxvsxXPWxkSheNEGQ+dB0A
Ev/WLsxuxHBfQP6cxLmoLuFPTysMFZDAVM9h4GenUmZV0Md5VGa+4MKnGNZ0IOPZ
F3pizel/qs4Ei95g2dw9WvatcAZZRzFr3iwblTD7Bv4dVmSCS+6vMuvsi8Nix6QI
/sjMv7XyQlG8B0ShQ1GgxH8PaHMUxbQ3gUQv0gMqgSuH593Rrr3wuklMmFNSiF6s
/h4WYUzCNbaxN/SjQ6Yk434FGTgKg3b3SHoQuPIzcWI=
`protect END_PROTECTED
