`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mHAA22qtxp3dXhQ/zH75BAVi9Ll7XJDACYAmVB3MmXSOq5uTRSo3fnHQNFwGE2Ir
/i/vozAzVU8EWxybfOHdPWDvm+MqYz1V//AFdrYkBae5Y2OZnl/c2Dh4ki5Lhsg2
5EyXQ4w5AnH+htB4EKxoLTtcM722FUBvYtuzClWpKG6nbnmaePTxIQ6ZtLlLEWOs
WpCTnCl/9QfWm8ByYsZ8/6fSDwRQH8IPnKmfP7Py9w/he8S36phxxhuapXmx3CIK
cFdBTj28gVecEVTa323pf2v/LG2ZLcuMYjxaFr6/6Q2iA4O+31AtXWqxyW2PfWpV
4dkF12Ic4Qj0TrOwljj9A3garZFpFuXXP1GkUH04zSVNTQ9IRq0WC52M1uRmgd8Y
YhigAINQreiD0NrJGpC4jEfj7TSUJ00nyl+ij5gBlOufygk7MtXwcLBHwGrzNcIa
Ke34fOvpSCJKPHAdkL8+FsjGdl5YN6AOxDbRzXgztelXgf/GSUcaX6CZOmE3Pvcf
FhyD38XclybvZ9Uw8B/BMql7eBVIL1mPGjbJkfGXwsk6GI0BD2nAExU9dnGK5DBZ
0PCLLOGUGDP/77MmniGcjJ2Me4wYzmnYOE3wLpoL7HfBRWP+d9TpOCGOlNb73Dbv
oSsUxVvG/vDzWwYRZ3Sho9nZhOU2MBt5s9ui8F43wesLqL+SVfnrBXWlBv0VxvIf
+fJ2fvYHAfcj4qV5q6KW47P46KOg+K1PP4uIHperwiamd9N8p00n3+Jf7KUS+4x+
zqrOInNIUUwIhzE7Lck9XLg/BcIQGJiNgIw0Q+hfZMlrjwDCjZAmd1UK6XWivR+F
wZ7gWXyYQRJw2x222voFRbufcIxskufiHF3whwuQDbPtvzLdmsw/HcJzgctXbhzR
4RFF2qrfCTulcR5FLG0KJiBGz5Dn0llhoxz+6bjBd7Ags07uQnpeyzqHZRwkxxSx
1gZecfBvEqp5Cl1mWjaxmx84f1KfIK5tcZhOHCfIQPYK6Qzz4GmrNZp8xWPXdh2s
`protect END_PROTECTED
