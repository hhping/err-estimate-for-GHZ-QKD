`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ww4LogU9fEt9uVgrqvKasXr6llaClAVsVOp4KVXHuk1sdlix9W2k86l5WXVCminG
y2IoG/y5sZdXk4C41qjNeZt4VoHwpC4B3Y4DnV9+r3yA+v+gBNhzkmmgpZ8dp0as
PUOsv2TNNga48ETG0PMhCj9onI/ubRtsAFPxmCqXn5qz04L7WKya2Sh2K6QesFpS
Dl3svNudIvQMaE5kOsX5Tlu3HDQVQpl1JMruLBQMLIgh/MkQ+P9HtDY8BUCKx3eX
GxwvHyMWOQ4wgq8LwmCa9QW1umD6EPnGETBKi1fUm6135iSag4ABkRLa8mfKik77
PfTt7K1sjjRKAd+gsH4IgVhAVlq3BnuF4ss/LarTDvWHr7EBCHlyIQEWmDZ3bOT9
yCBERAj403jOnaCStIxam0SaT6Ly4rXoisugACSrokm2+y6xzlDmLEAbEJ7DrQhY
NWBZGIusvxeYHzQCCKGjRW6kZJMMmIW7trITU7jBZDYPv+XolXq1GUq59Dr5uFlu
NIiDb9g9exxqrIDzN+VVQF7aG/Ku1ga877wvFuQyqcrXYTSNdQySEiJtCnM6oTAX
QdaRcvnYTS2bJ9ihZnyILNQR+iuqGqZsHNwKEcqPAccT73lFSg6l418FLkYH5ylU
8lP/yQD6N1BgyKdC/jTgh0SGcVPlVLh40PiI5JeCD1w77X8OZWTiwvDXp7Ewu5bS
Txck7stOQsRkqjptOBgSxGSOdbgIZRlHsHoIPniRGzkE+QoTC+aZ4f1stcYZiFRi
XkTmbL8trf5Gbja5lDX+9JdMYsApVHzphPXY7hMfHsZbPEU3UW6e08na+qfSt3l7
L+7FnOnYET17eaM2NJq01b5UymMuHeLKSlC3WNSQLebtNeKyHgqDThpYd4JJ9Mk7
xiUUiNZWUE1DQ0SVKLnC1Yk5DR7x1WVy9VFQ3NSs5R52YVrvWp4epso/2FkJr5pP
WPxhTubtF6NU23tI+uEjYYzML25n6dh4dyGhm9jLq61Pi8NfqyzQN1qtB+lEr2Vc
qkqp+OsQdlSIJXHkU7525iI+KkjIvXUUHuLIznFVIzmtWqIuXPd43VPVbhFM04ND
PHIYoTNgfAVbRo4hIsOLoPOTHf42bSHpykzBCj2HUY0fLBIa+FLOkkYoKdfTEUqx
kLgwfFdvGhHbElddBv/t4lBBzVVIGf2XRxrHDQHcjPnRByW26CLge/oz5Vi/FOL+
MiuSxPDkvpcSHi/l+wXIO+k5qK6LsEq7mhJgJ+XpG3rkl0uxUgehPhfn7bYxLMMX
YTCyPX3VLdE5mhdj9UtDxgJyml3lndi5cGqZEgXJy8CWP8CqxzvzW8AwweFadYsU
BzcHyxEXTTPHo40jh93V7oFYtNazKN/VF9mNLqSkp9OxgmKhmX23JC6szIPsE3ew
qins67PYvFoyVBSqZCnVqBRB6Y0OMKsYxs/5jnL5DDcwOorUWGU/twWuOsMazQiL
upyd8jzpz69CJ2YVhAFZDoQpUxidpBUPC9YHkAuImqlHRq93JVF8dRbOJt4Jwrys
xllQpMwblGo5r6VKHeQoGWWXCZdyN6LGNVj/l5T93dwoEbaJJfpQ53yied7QxFHJ
OF3oufDhwkrWkD9heVGsDlK6bZ3xfyxt5XIjT+OMaoxZ0OlR6kKc93QgEaddq4u2
TdRdhxapaIZMnLPQ2TYTrk0uCf5ThpQZeV11j+FTbQ3SAqasfnNg+KQsMP8JwnhJ
6T7NK+Fl47wghYjxbQbOupAV6CcrKhzCLbTx5Uue4CbAZk4nD+syjgN1w3bIRbdm
EackcJ4btd0zZXOS3I1oaUXRPwXz0Ocn+JKxBZuHiqpi/MoU0zZTRFaLsdYu77pD
B7tCzNl53OQaUcYRn1h2IYzv+K8IzTKJVsGQZRcUSTQf6v+/L8DQQ2KDbSCrAteb
RE7/3iNYNPEgMF5pI6o3uOO33y6WHE9nB2/AoL+NAyGUTFXl7exo9eBOrJZC1tvj
Hg9owxmNz6EPJ/23ZcCPo6fKEy3uhaCPJbdUie/ucBVZ6juITar+DyE4wMX5zgD2
1XsEUmQ81Q01TJWaJcENgM7aWVjl8eMCPkuJO+mfa3D3Bq/bE/FqTxISOBFEVA+W
XLRoIWA8EC+PPq7Ng8dVVt6ZQRbZyZ/pM093jA7bXT72dvEFWKck2Psu7djsCSKR
o6+HuLNq5WnkIWunTp4P6jfMKIhGFbfHBrhMXR5KBrXTC0p/66zPRY9N5WiIT4ML
ns9MHRgTxZ6+XwMZne/QhbBbLyDNfWbSdAW1jmjdEa6P4juHKunOhwXh8Y9TJLM0
9YEXb3egCRZHjxEfGY1VSMdmWQV0qenMniqXQZ+OSNSjQw1exMR0MvrpSrTyMyl8
t3JvKLjBT/ggglBNT7JhHpizYAFGFslxeIYBjK279b8gDyAjGYN23/H4esqpHUOT
sqKroem5R6wPVzpl/369XhZKFMao+Qo+OTc0HNUD6K0be5RgZjUeaFI7p2wpho74
`protect END_PROTECTED
