`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hHCDZH+aAuKnPtxuM1St4ms6G/Biuvc54SHYukRBmzNASc56errc9KsdzYd9GxGp
+RhWeejFaFYeh2CYLhtkZvxfE7Am1kQ4vWUlusBB7DAWFWotWhKAGUNU9DkLp2Jh
E8MbtkDPgeg1DESfwrM2iQWNUFE3LosdU7j6gNQFEPnznnZ7rb8VNvxQvrNdSA7I
sSyd9h35WtT17CQbm6GmvJoG0AP6vtYpA8iNXNrFWwAbrzgF/CHr6cFN4kbcHHNc
449rH8ag0afptcGQn623ssgtUSk/SO6BkZ5vrCQP0K6lPzqCpkeKug4qHLj5+V4/
4DUmD3r71R9EKDghOoq/nZ+o/JZI3XoUaC7bqaLiGW2qbfrVgUcofPd7vxehpg76
7WJi8lCF3MCpDmbO+AnE2CZ2iU3KGPe/PJ8xLhLMGsj5+g0q1bJ/M0RkjOuZw8xF
9EU7cAuU15WWatEApbzzvqoFT6zyPiigI06WtkgBmjPp6IMPZt6dSY4R4PeItDjN
DNGMiIkS+jDRmDDMqvHGmwOSSEiPu9OsHHzpAixQxbq2BVmL/RnyeM7EzcLs220O
p7P1MXlAlsP5zzuq4Bg3MAHyFHvWiCDuU+clo4ssqaR7FYHuEj4n5ekxePK8I2aF
oclBIJsI0zbjblZNhD62gSsgDs40VDxBt6cMNvz2JW8=
`protect END_PROTECTED
