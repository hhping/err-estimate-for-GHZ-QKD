`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hJsm9oK++duEq5Fm6n6nrPVYms5VoUBPOjtS3TldPPh99OI3vhsoyQ04j1Yi7LUy
DyUi+iCScpdSnOaUckabG0N3IDPRcaj1mDV43k82TAPC0braoiGjAuMFUzil4omc
BW5RFTiVaoTPAOd0921VUJHN1Y+mp8EV/Nh+xYMTxRN6oob6e+0qUk27coXaMVSZ
n7i7yILnjrDL4UqPl1xzxHhY40rmCFpeCYECqv/GusJXDNx/9O07QS1pt+QWz7r7
br0AGQMjmOIBvg+TTJ33MIG1344RC/7RS2qLBbHbzSVvYFls7MTe7IA72rEYkjSn
Pdwbq+plOSPfu9McJCGKQyuoL4Q+5WCCBBmg+l/tr8oSPegvFspPw8ZvdeE8zeM6
W5TbIcSPYFlUSuWQo8f11BhF3lXY4AnqZ98a5GFl24ghzU1JRNI4v64UpSxY10gV
2EBXSe1DUxkaw8pBR1tuacvV4vxZts4fEp3/5O9OoWvKy0LA5KmvBlkVgnCjbhzF
f+OioXCB7fOTvVtYqAv9uYfarIFXjsfj8CYr2W5QO5XZgDEfvd94xAjRTsLLPX8/
gRar2KGobQin9vbroBCCM4CX62A3gzv6Hk+IXBKWQiCsoRwV1sVNEXU2jkvZLfZE
`protect END_PROTECTED
