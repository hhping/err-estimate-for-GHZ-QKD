`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/7bbarM7VXBFGnJawuo46sIFYu336PIPermk5J8AVM1jFzy5ghK4n+B90wvHjFy4
cXF7wPkq6/8JHbb+NcmmeFiQJogCvLBoHCsGqyXtNjy8PvcdwzdRy9LLKueK2UCi
kA/F4Dkc59Fo2z/Qx7SfC+YBVH/4HTzD3fJ+aCsWtXFl9BHlQmNYAg+4U69QZKmk
gA8XS4e9g4owVV7LeieTj1ok5hdfNas4rCQygN4cRC4RLyyrImZa09qs2OqcuuDj
4R6i+/XMS0OalSzr5z3TeHIDMTwyfQHUUXyeF5RVHBO+STGLbcrM048rNFk1k0dQ
jK1oFPHyATlh6p/84RBigYQfEDF2j0CxwJG3Dk6nzEK+M3HxuxO2mPD9Dbpf3JRR
YOwj0oVpNLSNCLfPAk7TF8NwXztEhVQUI58ued9gQCRWcpve9D4f39M77VwTsOFt
eyBnd6WqV6b+TxfJFuuP64KJ6D7WHo/NiTgcIRXbsqz883haGa5c3XPRUSCucgqT
wLhTEU2b3Cb5yLYgnRpBAkLBMsO4cYylmM4q+GCpl3qOZe94s8j98tR6UaSrZk+f
idJAoBR1P7H5fzYH8pARjFikMxwbfyV5HWt5DqoKPKs2xfh+h2I9ZC2ab18xyI89
uX5by1ZaCfSSJZ23J4WqjS7zl6hpWtgiB7qaTRboMI6MeYaQGy8fCUQAn4rT3DSC
LSBI1s4CGkjAk6WCTF4buKgCXEPM53MFHucAM00OZlOVcy2gbS8RCgobcNhLohuu
`protect END_PROTECTED
