`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ww6V9hDv+f2Zjz7vwIE0PNaCNFWxdxjQWGOHND5BRjNLRl37Nbyh5B+wyrjTqvc4
epNWaZS5yVV5Y7DneqWZdNNCfPTDzh+ohJfj0Akmfur63Rdjjc0ZsB+02oSbY8TF
Q8OnngziQKlZuuO2eAPfHr6BPNvJDJ2gxY/MV+baf4dYQe4df9t6NwmgbctUAabc
YuWLJrXjAJNtmwOmqvTaeJmBPaEae32eIl4rNoEPsif2JP/cUH3eHrHHQbkd2pXl
LSxTU+dXO2wZflbk8nduF9IBPR8qRGtsRMx3/69dBoV6jKovAvlJqPl7isz3FxmH
9tYVrUPGHDuvOpRT7ifEHm/kE/vDbpcWETYbigxn8z7oOX3XLIhDYlZT/qhP9iE1
zM9q8t0QdQdWIK2Nc8Gb1M8sYvJEP+QUWybXMahUoBRMkrGDQaaxJvGh8MzulN35
T3T7uga07pcKLogD9DJ9AIxoXMJ5DZr4PzdMshrs2YXifR2CgDAHhhnrk4jj6VbZ
nPdn0uXsQ++4JCbTKAqtc0NgNX3Jij0reXlZ7tDDLOqn+8ZaMKg3LMavAq6qubCx
`protect END_PROTECTED
