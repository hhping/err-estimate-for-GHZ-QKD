`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nNDHWKTAOJHrJsRHg5UWo3bPIegL1OUFPejrKGlfQbxPF/nPjkm6sp38ds4YL+Td
OWM3hGPSrtSIDNh3eClaFsEFnLTX8TU3Q6RMwoEV5qWXoWTdNcxpthhSCmWbJPdg
mI7dCxei8HCLbXpZRNU5lmzNZyRkeuNtsHFezDU7EFb6IES5miiGU1FP6JS2MXgd
UCaYeXP6BY/1gYBoLUBottSRiIjJaUlV4TBbT/8+FQe3iWrD6u0WJ4jNd5P7Etka
nofRBIOC6QhAseTl8itGz9ubW4MBC+X+DNypm8AlPADfkQYz0pGUd655aezD2sjM
iLKTUdLEaocXJYGZf80utinPmskBx6gAdWO0Xv8DWC+ssTpV4hdDcUjrm2Afs5t/
67+2Jm9BECA6fdiXsNw1qEoZVqI2k6OFOwVtkt9LBh5EjwriNW/tlBzmtdST1k95
c4GXo4k1kzBb1GGc09KI5cMStbJwwDdsZRc384ZHmZ9NaZooivuBvb1Z9UktARZy
NyQQEZO45gvZCRM36jbytH2PKyqz7Z59R8nR+y3Hq4nLRN1+aBAUmWLhlKaRPuDi
bV5Hlh2FjlJEHvJoosplcguLaJXBVqXUPqkIEStoUU10jC3YJHgSAHi/gbeQ8pMc
Yht1fUqOCN90IhEwbHCfNbhWkfQLEvQRBeaNvu0hFp3prMmLXly++D/Qfw8UY3pk
fNWe9nG2v37NPPjo4fZk5n4qeBJ3eyEblcdYJCX2WZGAzryOXgp+qVAW+AbwXgLL
YjXe+7vxN0PCvXEzTLUyuOLRAbXFulQwQmd1HFmQ4o7NkJC7Bymx4tdIYHRRpcfg
cec6cMsUFWivWJi0VjGIsMaRztaqiu0owXBQY+JnCcXp1VNCyo0JVAlqVNPD8miI
P5+dSpr/he5UK8dp07itjHo5k5tOPsWCZvL0hcLmxyf2iSrqQl3TPGhjKQKZlT4W
Wfb4Di/V3XCSIJb5oFUJmnXNXZ+1CJbK0n++yoTAeI40x8O2HvR93e74kBLW16Ee
RbB0ed+QWjtUqMXGZGajU7/ls7OgtzkgVJB7TT2e9z6wDQYGYZnTZGI5GTAlfLMm
9LgPMCpeye9LdI2U7gdMQ60/EJqvS4E8z1jqi/o/yQM+HeM+1BuaaLZRHOymd1jj
PBxwXxZVQ1mzD5YPi0s2YxCoaGM2mXAtDUqIblqZcW+zjhGDetM7QKBsave6Ii5h
jAbLQYBKCnw46wuJR5ROnU3hiQsFtAEf50+DAsHQ3ASugL9m6qZpnyqfQEs0Pm8z
JYvBpxJZeSDY4dR6U3/FbRMaCfkJITjwFYQBiT6EeTUYHFycEi5feY9gENxF4toH
puFnJQ6QxydBllcHnYSvGhmU2VukyqphYeWMKqhyWwSlfHUwKNV4Tr977cHi3G/y
BgnkGMDkVRAOZnWOtTaU9KHwEAbC7hLE8vG7gxEACVkmRW53iRIofAAQa16SNuea
MuCwnEcTqZbNyT6T4TiOoct5sRB6pi/Rd32j6Cys7tLJn66G6B1Lwe4IVvgiszuj
/dN1HuLhIVmi5zSAEV6UPt/MGuzHQzkvqWlcsxss34F5FxaSLncd0NAEyRALn1mQ
oxnRqbzL4A7IO2yXDaXK6tDqBUkCSbVqsq+qp4lOO947+CNTCJrgEsAktYsXlAPT
eGXug573c8U88mYlPjM2RQp/Q9o9fFs2laGT8yF6rDSyAeck641davd9a0yHclsU
NlkvXHUxP3fQtf4wgGfmyN5AMpVJ21sDglZcfdJ7T1/WI4sE3+5bO6OH20Y7OVSJ
Rk46L5+Zk+wUMMNVvrDYBZxn8PCThqWr2ORD7X/8x3mx3dINNHgWkwCsf63EXgMz
dakBNftQv78jXeXc34OEA8+eED+o8LP0vO0/fBqV+C/e4kyqZGsV+0O74e6hW1gn
ZtdHwLWAjn3cPcmcaj16/0dl8TCdWtPN2v/DHFXgh7ssNElK2VewvamarW5WSuAh
Rx5XYMw9/sx4OGjXjbgqLhPVhkbDBTTECM7W4gDIUdc2S9DN///90nhxK272V/b+
ZVzlifWk/DVHBKshWHnH1ILRCrrwFTQnGIpMkbWBnfi0Jve2klCTN88vXtzz8kjH
vJi2SARwspvDyMj2p+NJjycoruS2XjNfVoBTkOB7m+0y/PAppklfkcdRe5xp5vs+
X8RLYsS9tonuVETytgzy4kqfM2tyNMSB7XVA3EY1KtlPvK43l4gSfuGjjqmVPya4
MNZ4qL0gFt1XxWSlrlPm4QGKVw2ofeffS2m2y3EvlDNQclmjoZuX3qa5fSIjIRpj
lqVu9D0CWuvvtzrmBX6STAFkdcxX6pivOSa8kifv64s1PA/0IBSgxFQB/6NCGFfZ
beTRAP6D00JAFFeIM2UqMdVjpg4ZmbsHDnjQt3I5+VAOurNn6QOCzBordZ4PYhcs
hlerzNrwFEbcB3v19FmlkB3lL/4nKXEvWcwKloU7qW8MAuznRtG22lbBmdNKNi/T
gKci3+U6pvqm1QkCM7/fM/1oH/roBRMRRp0thWaJsl8skc3Nl7PpfgCpnj2dW413
uix1mnE9zjInisZ8WkIA1cZWsBP1oDOSrCgK5wPEokrnaDHei5CYk3CuVPhIckJs
UgSBCQjPcG93AO793rV9cR4KdJp00CPoVP751PE+1DdeWTsq93l6NarMc+pHcvi4
kIT3Cmr89DjPQ3FUHA0I+fwCki/3UNoyGyyS/MaN3N4GKDcFwFB7kb2a3FsJEQX6
ATbOYrTJ/fcft40KTHpmQ73X0GX8B2JSvdQPNXJnD4SJwm/Nk9zZK4fqDU6EC4Hz
7nAGmN/+haGSKJM0NHTdjX4B4q8X+VCxDIgBz8M2jdOO9EIKn+3j9H4ECXX175MF
+BnOorJAjwMP5q/qBW/Wrvws/xPSHqbEwGKGGUEbH9R6AYTWCU7yuYTkcOhqv2A9
aHqhRBvhPtfwXFVLJPjuqzKr5PkR1ED8MFmUmgGATJNELUiQJpgNu5K7gr6VWl8a
1V5wSJphidepIUh5Thbw5C4SzQLsM4Kn6F7z7gYbaBaH0FWRDibrFJfvSDboJzg0
lnPl5ohOTOKq3X0mQaCkqFUDpPUBBu2skdkWBOFfCfUCvMu4Hxlsqzm1mkjwkDXi
9lfYJwQljM7q5oJpH0YO8WL+ND3fnfF0axHhJ1Ir5s7XYoYSzZXNFvnkImPDmKLh
DuXeLbWN1UURvsX2ubRegSsrfB7Tx30CoJfPv254QKzyiqTv4M77ESB3cqZGO+4h
mmjf+20YheoiRtty5RTnUgqBQrZKHg7s8IsPqqMM+MClzhg1Hkx0eFB+k404QDEy
ttBT1PtJNCogw9xhCbuV4Ai8w2wY7q0RUxpcHTeKKcGIEm9H87JqNgH318OXBVty
zlW95JFr/spPGAMRa3E/Fi4jePLqxzvShXb5RVMEjuAYdNOuf32s/6qVYQdrx2c6
WjjPEt3+MoOnaOV3fnSsQDqsu+kiA1vJhWUukbEne35pJXwRhlFu1/6y+maLNN2C
DH+Eyph8AuZYCYzf+347/wY3Mn4bQxpmo2BR/USKiiO/qFuN3RLOaoGYJapRi1Jz
EKl1zCm3wMm2q+r4TmsMvSx7/vEFC4J2wLpUnjXUlep5JmJcyHrtHyH7cC8bJUn+
H2zKJSS3/uqfe+eep8jlYYFX2murBMUQDI8accvT71ihx8Y3Z5tl+Dq0XkyZL3ee
EfXeiDRqMft4gAZ8eO8/08xHNrDK0LV4/uFXHVd0PAJ9+vZ9Lhvw+d7dIjTrRaRy
WeUPpArPlXFrpJU0UkcgIMH/gAbg9TuniDEyXrBl8wB06vZvAfFiEQz81U0Q77xn
R277KOu/FTGBv0WpLmJaWHjUqUFXbnmxJqBi5XIFNtJ9xLtCyg/6zlg0CU3M42HI
lP1Q4R4UvJpLsf/aPyKoz63x4tesvydy5ilELqpr+TEmbBtDFadQTD2ji+ZRy9Pj
ar5o3GMIdr6gqgGIR1upN0HyP2K7nsAiC3QpMDDhwLVrFn1P6CYzFLxM8HOfyC7R
D1R3gpjcFBUGBIz9nA3skusLUqK9ZRPUymMtZwaCoXZb1JaNs9p7Qbpm45HugUrZ
fcaxzhkPfvdJW4XT+nlZz7JclVaVGZYCgMnN0N16Cg1HJ2W66zR5s1xsdt4v8Cgb
Me23oDWX5vgqKWgl8Et7bhWw2mja2Y9WBEgKAYIWSGvJz4V0K3ql8QDn9+gV9xrG
bDf9LbZ2bJ1Y1T/BBwTLwpolHP3SrEJtGNMYfw+3ER165Nmwq0cXDN78iJE2PYLf
PYxoMT3AHiwxk7+Mplhjm5/m0xiPhPqUwVVNqDvlwrNKKewQ/9pJ8DFiadc+TvMa
QU0E0hynXg5hETC2i4vlcOhhVrwcrDwCHp0WjbtHuMNkcev5nle+S9U0Bo/6x8YO
8UkeTsxJriAYiXWTyjEv2L0VpY9J4LAHnlI3oQ3zHlkbEYvBFtwj3PVewT6lVjDF
jg84j7egdiMYrngTGi5fHlC85Mm2qGim+/qijJTThh+GUL3Mbe/Ewom340CatLp/
d88simFitKApol11c3qOZeMC4VI5unpnGuRjrhgT1Q9b8ELs2HrBwlyssNjgw85N
vogPl+FXdJU+pRidyGACaFgFvj5YRK1vjUwuE8f0X4IaScaHX13KjJrCw50lRDf9
eyE8rakI0hEa3BhB/MtQMXR0KFkrsXJG1f4CIg9pEXglPmHfO2lzj8UD+UzKyuAa
+8M0Gyvn1ePXRnrpsAueIqV2lU64rU5MRXlh6U2ouwh2Lo0zGA1BNVnB8iSgtaNu
YTi4eKDOQI0PNLTAyljyeSFOXRaW6XB3NgcQaFBpL1Pb5i1444NzgdgDuchRe7oB
InAv9vN/AomSnW4y/VDOlmEI/ak5+Y1Cnvt/b8R8N9BNLOorDu26kis4D7kefF9z
dyTVQG7vRxQPgZGwV3A9zKwm1HirbzFMBSwZu17D20cfXudByMsSYVlMyoMVG+rC
pOcW2RQkSwF6zG3i91jwWKdsLQCFEGShIaxLg3fQNLY9jRGvlVb0gqfbHy2NLfVG
SA2b4BaqZtVo9Xpz7zDNSN8qDFR0xNk2QrwDTUMVID29FcwFJOqFoiC6BA1FstWl
bWTBVFYkPH/UY/ZaQZYOj9j+2JEj+4W7k6308SbsrpW9ub44cVSuKDSFRLEZAO5N
BE/YyneBX9eyizkQyzuq2URb/8VsCvO0RsvF/Re5SW31gqwf6r2QlRNk35dViP3p
00IiR250XjsALokqZPlaO941qWQQc7oE1NKkAgx6E2UzjBogvxS3U0SZi/X+g54P
6CI17+Q+i6qO6zkX4aeF7DnHbzqL5N0te6sh8DLzBHjCLRdxXs0vfRTI9hHCGlO9
z8LiAcmWiv+E669VwNyULAQx94teuGM87d8RVnTED8PEXSdD/KNfqMxkSxV7WDp0
0X4xAbZAgrl3NnVZzVY+mmreFYgESRq0jYNjic/ys8tePdB2cw0WSKHlbLWc7EbJ
ihWkTGO0pqzMIAgKmCoP/7d14pwqRNjR49dPhbg51b0=
`protect END_PROTECTED
