`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N7CASJylkLOUfXzLruBTgDwXnMTyHsSrKm2EyFYaQL0AzaV8ZLX4avOmE7zq1pQN
Sn3+181YCuAKpEH92bcguMRglzWzomNA0H+21FdAYguSOIkprDTMpU01S79jnTSQ
Fs5ocQRREUr3Z0gQtMokRiFFsUXzUZxBwdGI52NRNUfaGgmjAhehgoU5LXswdRVr
RM4RfkT2R4Rd8CqS3x0E0fQAn8G1jBWJZrW2pwStWerz3aUjB+XA7tVL2UmxqWYI
ujnETNJRzFynTzIDSyHmdF9r/W2upgy026SvCNiPcP5L7M26l28gSn4MQ7PdM1AO
kEccCRjPUKgnkqqu7EIhEZh9XokcBbtw/aE6qJ8Hb1WsTRpTYpsKcFRE8l6ujBJ9
cO4lXgMCyH4dOBQ8WNsfeIFsbrMAn69GKYsBjmQKYX5wSvxaneNEVIHqskL49DS/
cgfhS4H49C/UdDzoKIDWtJJWQ+EpeKOS3CTmm4ukb9o0pcvTJaO7LkIs8Tg9xIWH
pJfIHza6aRPMouM6ZJpJN3KJjbPh8x//7dKll9oKZ9Fa+zlJfA5SZv+BJOoUAMXn
n3a/sRNEOCQyOk+a08prLWY7rA10GbWp5I6r6JgvmaEzw0uVfxzxvg0uZSKsqXhf
4+gYjqKn5kEZH+zsGl6bRIHX3fHSNr0BQUBC6hQSyneFQywbIa8QJ0VkSairC1bT
BNbBcaKj2u+LhpPNICvFXB1PQUf4nVOrHFwR+lQJS4E9tDwIcVTfWlMl897imOnV
yEtU6HSw3W/TIgEMbyJoFVup6sfKQGFjMCXaGPc+IP7nTChSk8QAZU/4siayb5k+
xmyjgGFExBQ25iSCklowyzUj6JrVrv4iWUnb4Y8Mz4wwCiAw+InMwIpuGUev4KPo
5h554QYe0ybqWeeqwTUa/AQYpbruQE1h2UpOnCegG05Yclit87IJzthJi3oTQxtx
pPHhV9+I7tDNLVeHqvlSDXRHkyPgtpBNFw0QfAP9kasQeGwA1jL8oxoPI+JX5CuD
mmKhzTgkZYhWtsOVVpFqv7xKytspNBkqDLxfuBxnsUOIThEjJEh331TwV8y0qp6d
mvqHm9N426Od+4UIshfhgOt+0boq1+Tvug5IqbwLeUSxuiHj5gzJ32e1fWrFS+5O
w82UOgC1U/90Uc1d9JyMf7M3ASpb7V53+U+mNQl0hzKgOHCuVBJQAvVxokirrAUL
YMChwwWAh53moCYUXbYIThdSfpD3HZSmnx+Tf0i1CRXKZRhpQDpuU8hZCX3lS21R
9JIhlz2884Mn6D5pfXBW5Mus5KPfLlKmBtXoTgt149uTim7vh2pj2AN1KRXdjHwm
YszDokeQsAMFhqzed4L9Qgj8Rn1HgrZiejJDBJbhbUpWpHZY0IiNjTKc7ssS3MHx
bpV3oGFcSxWTm0d2k9rFu4fpaEDnXEdFfll4UeSmibFBxT3J3pdg1aXOrrSVkIFP
VqHErmdz0XC3/3R3sf1zDMHQvTVEHSPJ8j+Ls31fKu8evP2yo72Pt/ut5Nk/wIjQ
cG28ajCk5j/DnTNucP3nRQzhg215AeJD7W+tKOw618eM9SLxHaiuoh/rYUZwAkpp
w3naUdQ/pkl/FzAxMxRPy86hlOqt6ob4XfFDXJ7SiWqv9lCYh8Zn8PLvGhp2NLBu
u8IHlmUuz6r24MecxyCyJdFaVnVgAFuA+Lt9bkSrDdN/Txb9mwbmuZ7EIIlb3DpK
2wJlqpayK2w76/aEJvE96eJdrkx6Up7Z/tZVH/HOmBbB/mTWVru/C0Kk8YkpKrDR
9WuSwuhcxmhA4DCAfrAmqROUdPcUX8MrvwQKxV4V3hduI7CR1MJBSj6YDVea0No4
Zea2xX6GqNur7hSEkxc8/DH/q4LI+gop2x5MA9ehynzrltXZMQpMyQRCY/CFbOto
Ore1Zr23IfxyaV0TBcQb1lzZyHeDbelrwABcmUAFT0foBRztQn7txQeNNcrBZcUo
31JFEzt3L+QfU4D5Lvl94E5ARk3FS2QCCdn/ffPHMRZ/GCfoOPVPlmLTZOIhd/Md
2vKDMkk2f0lnlBFbtmf87gO8N+DT71ruxFDmFS3i0VUsW71Zwncd5mDVmo9nvLr1
517eeipoZLRq14Yz0LwzCvxIXmb8SJBmCLYAMiic4QtZqsFr1UfsHaoXSLrqF8AA
ZL+z2nEpc8VtNbxG8Fv5GXofoWRRgyXz55B2nZ8taPCV5lm9tqbh8eHFy/YE2U9f
HGmlIwp261b6LWuIMdX9BRnwowy0CtbLIQW+Qj5ddfSxazskL4sobfyLq9gi1txN
kPAN1lX/AYQiL1NrwYrD+XxuAo0afNe2wKFCAJub/CZGHZC704RyrCsD0QglpoPO
LrefFOccdGtCQVPy8rgHZ5kw2OtAEtxGm2XE7S3ZJsGuD5XIcAT/F8Skli2P+bYM
3Qfw3lc9fmcdOuIJEmqWKPme7pEaLh5QdwOA8VHrN+9O5mf/uAa8w4E3WSaUhWXM
MCELdDilkK5VqViB8krvVT9c89DJC48eilCSYeJsnBI+jTalNCB1c79DNYFW58tE
in+JLaHnO8D/BmrHTv1kDcCAJT9Cm92uWcxGo3Gd0S1qs3fsTgQngQMwkAB5gVRG
KFxFkWO303uH5b9wDg6JHYGg3XZ13CDIdWfas1Kpej33roROFitY8panhSh7clTc
TBiDAlgtatQkpmzkZ6vadb8sUjRkJxqJa0BPH42CvYdY9p299AAcZKf2vxoIyTRd
0WlVLPPPBLjAzuee+fDfC8FBt7t5uylS5311Po0R75ZTSg14NLYo2HUchY16QxMC
Dg+BJqH+PKSZ8S9+xhNCrDXFgagknCaDrSFn3+Bi7U9YMLra0y+3mMFKEcClmhoX
79VXhBhscabz3dmdYxokC0oSo0xZjL0twBTWzk1g9d9xvpGPl5Rtka82DFDWkAsh
7Ztcg4P2aBgbyBSfsSUa0wS/JhequTLavzWUqxPDjDOjlduQze8MwwnTno9vWScx
8zm4gv+OFyUaMdiYvVYi2AWg0agn2hmqvIe7kk+6wlF6ShYC8EaoZmMc87PshiYN
k17wm5+UEDHnq8OvLNrAoOEkwFPboBNsIGsY14jpu0R6Siv1R7BSEgei1Isp1KJh
zHVWbOFHK/2LpLKCbtYLbbiEcDoanOQyIZPT169kU1pE2JKcw0dT87JIvah6h/W0
MQzUzCQ2J3HZoBRfRghgPe3NzNj7qYhFBdcMnS5C8Qa2xm4Q2md5rllvf2mmB/z9
0wqoKq5f7i7l8jLynx+CJtdfLx/10gfcKEMUXkiKpmST2mDG/dEuGy3fLYAtX7Wa
dlI94yrgsHeFyp5+si35SgOkE07Tg1ZKW9x4Vc3wVBRjYrwoyHEcm8JUv5C801Q+
g2kOeAQu0oqJAMbAlq8rqIWR6kdZlFfdq9fjRjGshjvYJv27woWZhclR7eD+PqUP
gf6/plULWg1SY/c3VeX7TbKbZagOeyZLtCNu+7yYN7jzoCUCFBJYzlaOeWFvdRXB
ikypQHDiEKBHABXqDQFOPxOgDVcHIrTWUF+Ozm3z+Jc/7kYocry+uqVLM66UK86V
9JmrNMKNpUDquUe4kzoyhYcE0eKnQLZT2xpwbs4m2xi51NN9DmJKwCsW+QAVGvqz
QrqxAG/ceGf96yMTsZqY70AYNdcm6WwrTSbrKFQ4gFP6F4Pa0XweGwalEZGhPHK+
gvJVt5TX4DjPZKlWuYxsts7o94q+j2W+VlIMLi5UxNXLjyTn4q2ssTPzSzqywYm9
wzixnhcfwrALM7jXARh4mpbpubnhEu3kN+b9cf4IFnF/4rqntp8DJaCYAkiVBAQV
1XddLVqvzH8L3iWoDQOYosixlBVjTT58iriq1XUhvYXsQNvNt31NmAcxRGCGCaoK
8qvNzvh7N5iXZ0l0nCFQLT/s8EH7Ld/nHNHWfXghBGhiXb7TFdHEr/fzSbVTZ2zm
rSgnd1Y2bu4EpeLCFs4a0Jv/DrpFl3nNiDdAHRFpiMp7TIJRimZWj7Rj/2FD+psp
NWFtKeAIg18LBoZJMobtnbLDFhLcZFd2+zvuQ2vpkTJRM3Lyb7NzGATdMY/O+tLg
5q6WovPyJZ1G/91evHxl/Qc/lyWx+hHzqoORtVzAYhYXH06jQJ1bIEW9oy9om0fJ
kPens8XAXQtpXgkzR/fkq6zGStYCFbSsFNQ016zRdFtguf+LqhZhUinY2i1zQbD5
GoUmyw3AZMMeObsmsjJIzcbXWNqm5PnyoOsiDH5dESWwEicNxiucThecqwqgeFn8
n4ZPGoqjxphPVbOKv2iW63QAJw4GQxKU+5ux74jStdad0dY7NWpFk8aCjfNIW5W1
PheMZpbGiSwzmeGd+HobeVtFEbBlKPrkgxwEom+t1zZYFwGMuTa0RwbGiGlfVghm
0246ihv6MQfMK6LxxqXUrSL+RE1w7QeEPHr2faR2Nho/+o+i/CBWEbAdAO5elgMg
p2Xv8d04wtoANfjPO7p8Kx6GQx6Qwq1P34tyBaofrsvd2NXvS6RIT8a6CKJu/BUp
bFgNOAcQisbCTrdNUHA/qSCq4NmD5t55LclNmHJUyqL4He2nqJ1v9YABX3IGYC4+
wmW1plOuI3F0swGanNHPi2CVyLvsE5RxdotcDmF2D4RL/jCW2CWOm2idBdPyiG0I
ZDc7uwauyP431IrvFyF3eXPFZdww8OBrsmYLwurU56omtP/NfBo46aS4pHSFMVv4
BUWJU47jTOO9tkivh2rGFbIqy6kcWkTL3RuF4ej2PbkcpY8jgf79v6ZEFM/ltMAP
sTHnqBjpKA5T4xaIDJWMLXND4B3YBYBT39W9bRcdi1Iz6+A6kWgl1M+sMPQoLi3z
ZUfVegHcM0YvPmhPDaJF5T50oOKN3seuN8g86mRfm/Nv8KWbnVBoTvZE2Kd3jRQU
BIvbvzOHKwPS1QHK/7/vek2IyokHtCQJv03jg9yL6xaE3lNe9JmlWD/3zlZcL2HZ
DXKUkfXrhER5L5XpHeAgAyhd3I/wnYA5r14jEg16oJW3KrK+l5fvlwutPjFYEK2m
rGyZnEbKZf8FjoHV7M2LE5v69GaU6zQ1IvVelFYM2tPBvuIrWl2b1IuCu4er9jE/
0VZZNMWR4vcWOvQochswoTYa1/09m9BULLbmqDy9KKIRGvPj6QKSiyErptI5/6C0
AbQ0n/YRTo8yC6J8ZSw8VR+Rt1rhFzH0V5j1zRzr+ps4WpgwA910gQVlcSpbr4uE
b619UbykC6apL18aGLfLXcHXMbyYn0M9q28wD5REm+erIT3JcUJaNl6Zxmvl2pgG
KzfeUFTulvntkuv0UOzH1xm4d+igtf6nafVEkxV5qbfIJMUuBXJc5tS6jn1Ftycj
8+bcKDlfxnPOLvpVb4WvutwBJzuaxUKEzRzcpw+LcU4OzfO6BGMQt/HjL/pMaudb
P7sr/sN+X3tXb8pvl926cxhgn0PtKE3eao9RYm2zHqFoiAoNK0ZaJ3F4tRh7GjLC
bFDJL2SS0V+QP+2Waeh7dMkPD7wmLCbOwQVQXrMMOXmeMyv8UEW32bOluYBJdE/z
oiFK3dvEz6G0MktaLer+8SndFVedJVmBM1AN0cPrQ2FTrwu+y96+zry3xxchWomK
VdjMFOEEERBTEPC2+42oPNCWHvU2AnKjgEknYiz08xW+QEHUte51RjwwAFbygm1E
4XAnB/bU+HayxiR3LpZHGxYu67Kdj8Xd0wz0yximpJJ6I66pYGBpfYpZ5ViMS/RE
K/Z40AcpMNkd4RHssjMR+eNohrh34SClLDpaFryJsc6gnVUPn/Bze2GYIw2/+ikH
fST5Y80b3ejCJwgPEKasoUCncPritXH0wzIPWH+cQb04MxuJ41292YYCpMwb1ke/
siHbIOtO0kML+uuck//nQA==
`protect END_PROTECTED
