`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lnC3VWZjrIoCn/CXX3hqPW4l2Ft4sLy8USezUgav+9NxSWANn0GWUDt1bEWCdfOo
UihnfcAmpUA/f90/daXNWy+Joy3+09zibF/1QMKykVRONqXL9ryexIJDRJf1zjQS
zI/A5WGtfjeL5q4cQ+grj9LPwYVpq70QQMIrod6hi1kYkWk68MAXCff8f873C0gd
koMHNMW7E2q7R0TBruuABF6UQMBt5Ir6fnskPV3SGy3plAyuqmzyvvlvCr5mNT7c
2rTA0YhPhb6zW0Z0SYfBa9NId6LBz7gWtEdqhKe0K/DJcgWfh5epiJ2XU4v4a8s9
jat2JdejJlaBHkxau2ImfJaV0tPRCak3iMHVKvxzJea0AIvdBclgJdZbanyb6xek
qGWxSy1MkfqwoNjdHh/A34p3+J1kXhRg9g9C6BpcanFAVyKHwZeLACb3Izk6UrLW
5pJsMZ83j527C9Qf2C3KEZktzMJeGEou9o2BB8p+w8CIG7a4Ytr6JiznbS8Vr585
tUqei5x1mi4Swi1dnNrMd0WUJWgy8BkEAy3Mz3KKw/YRuzfjq3h5SKPzLhv54Nh7
WTLKqfV6tyIaautN6zD8yWznBaHP+x+ThhJjwM5kV42CX2oplMYqcGhEfbuX8XvY
31MYdH+hcK03gf7NznvJOCXvFdI1d/tM9gTo2Uq+EJbPG1GQ5GbhHPXmn66obwy+
DvjI7VWOiHaVu+eHk6N7hN3H/yXjDnxJH6ahHqUHhxEaVLV9HOpEUWEAW2sGEvQQ
IK57JS9GUcz5K5yL6Bdp95+FQGU9FCfFolgzJDnM6a7A1k2lMxAJufAaMKJmsoi3
pLwgLnoQMGDRFTxyjt3ErR+WtYSKCdyZCDpT8msAipBys2iI3KIJQO/gNE57uTTM
0eUD+qB1UJg6jCeA+86ha+xEieysmDl93HeG/xblQmmSssaNhjGwhenCr7raxEHM
TaeGrHVdUSVzsnSiZhX9p3aMi8td/LpiFkbwL6wyD+qUgwJD+2nlQdjLEp1Vrng5
0yPSIw6a7Ec3HeJqflWWJS14zFVrCeJpIq4swzBWNCYKZ7vHc2s9ZYLCAYZSTI6Z
juWENbv2tEVAIp7MtmtGMiy1Nh59f2wHUL/FjapSzTgMiOGm4zW+cOggLLEx2hR2
ybO882f2iMISFjzoCDCyTZZsYHsQ3VPBW2PJFxwlU5tvmrgXPhXTwZrCdD5sK1AV
XwyrSg05Erf2unNNY/WjPj0uAuzEr+JpSQRxm4u6nNtDEWmdGwUgx/tYSxs30UJe
jSN5CzSiEuudt+K8MuhM92I6EgiZuqJ9dmwkRhlBODtru1UN7r4OgXrum+jhqOgB
mpV7mdJyQbjRhW2HTpypjVskYceMzfUBqSi+Wr8jAWsaZdolV5yCoImTwVTgUW2b
Xh5HLhYZKwODxuQbYaVYCQe3H2wLYvQMF2UojnfHzS9c+oq5/5aZWLrh1R2JvqrC
asw98Nl9PjPynl6jKhwVdSpWMISnbO6YDOMZtg8UJ63fDdFbFXgtouUErQV2INuU
OP0F9M/r+/NVYggWlClLN2gGwjxczh3R21ISeUGbASddpDlB+f9T1Je50Y4qrCMP
axoM2OvpUC/RYht9aJ1agb7YAb/G31niHos69KsrLo1qI+zJdcPJ3iyGj8hfFi/a
HQdZVt9jjlC/4xnBCRB4sFs4dSpp74sJu289i68nEvpt9IcIdnJ22g2MziRtHtii
KHYZmolEknnNIAOUQLXWRbcl2rL+Cd3vY6cUTNeDrtCUdqYl2I2G4yx+kGtxXs1z
y2+MmIt9TaL2uambsWiQuoDi0N6hXAuUEgl3m/AR9EOHqNt/MDB/N8bB2Sf1Gbqt
QdF+ttdt5c7ftq4FXQYorHYdm/zRiZ/NGpkNcVw+f+NURsLVJun1vIjpOBba7EBI
aAekyoaLMgR86X4WfmSlY3GVCdfiHQh9ZkZLiEDsqMSHKbhB0FZfBUVWAXQZs4vA
4aGhC3N2Vroyvw2YXR6t7bSzNcJ9DhsHG/3Gq8gH/+3aEa39AZWl8OIhFnjKO+yJ
RldnAQoKX5SfuX4qJiTwE3Nm1IKR8kqbfTBMysMpIFuZ/0A6rCN/yqYaP/gPAnno
J3fJ0hf0iylS6f/ov0KMilcxJJXGT8DFU7GEw5lBdvZIJNuLfZ+uFO5cbm8qw6+2
1WsGHYgDRboug1KqTDbt4bccBeLpBj+GAoXwaMjMXh0c72A55CWRLzat4vdROZDm
7ZiAK3mt2Za8R4mmgpPU30p4N1w8+mAWHLVaoXuVEKk9hgq1ihIogDscKyWGm2B1
30Gnr5r4CMKfh8RsLt6loYp2wP0e94XoAwx5RA2jU6d6cZH19+PAF9vtVXdCdMXC
vHUTF62efGoy9WKADZtQEP69zk/9Zu8tqyudBTX/zg3Mn6c/x1zFXATdU+H1xCOF
nddxVRclry0SwDX4haVnFL6pqDZubvk73YkezyhbbBXKDYErE8mbq9YMp9PBQj3j
4O/uOPW992kwYmLFMt8Ps0QkkOwxTiFRWes1ULCJlHCTNbIr9X9aoCSTrACxrvu3
97ozdFE/e+OihVF2IHOw7DGUjui24ayd/YNNBnsKemDM1selggqX318Frfu4fG8A
tb+0dptV+DWD3OHnX1wD5UWM1lgF1C1xdkgjtjf5em4iMpKwaAnRAYD9W54RiKOk
TVxAPJa4uOzo1Q8WLTAhAfECdm++OyYGdEvg9Q7+GwFVVJ0PsYBxau6aqzpJxOa6
TdSTeHuHyCm6zpAoaoxtlNnwegwr6HNBhbYhLY+ZidC9c9o2I3xTH1syBVOUJA9h
c7l9dONGt4HyhugugnDeDpnSbaFyc2ZhQm7AD+Jxmw6zG6sGcj08nGzGeDdtwFVM
SJR6s7eqz2xPIdku5fF8nTYr65aF+92qb95vbBoS7NyPRwQI3bxuZoezcNJ2tuU7
ZbXEanvp10yRgfxMgjlZgPHnhvFL3ZofP708wWajppNtwzCjcDvUqP3hGPgnAJ8M
XTdRY8RxP2SgrO95sAI0fmU2fPFOhdPVk+PaJ0PAvaU59HXc8G8IHspWHk2KqQPq
MWPgAYYptSWQER9HwDCp5H6SQxurAiP3CRDTHjZktmXnaXng2wpTFwfvfZu4QB00
hGf6YqYUSKnFX7fuVeL6ri/t0oG8V2DpevF0XuKXgmXol2dO1eQnpUSbROk9Uqku
AgHjN3DK1UzxDfII6j3xroAA6tcQTpjkanEyfCVtfI3GX/jBFWsTipXFGiOPWAyb
vgSWh/fpyBzatsw8S3obXMs2eo496fyPsCnBnI815L8oKXyhjWRImR1hnbzwPrtm
CdQ5ibvy7Gwxw4E6TMVeWeRnosAF49yx6wReMXmqeOP9dwY2ooVEzAEked0sfa1i
h3N4eOzO53j7G29c82TYX7jXaCtUqD8Se9oQh3Yr69Cdijml3oG/NPAu9FPNoU/V
+SJUWiUpnM6H+gXUYILcMjcooM11exBfTE4cJcvAVtuJAKia9Vo38m8I5+JRvNn8
my4DPBxU+LnJYPwk3HfotSY+4VRP+4YAYhclLvWzvjlvkAOaZHwIK4FFc5OhRFOV
6sgBKMj9vTFKZTdjWZ5smhUckxrBi2HcQ8lZFBDCYGQctI240wrMie8NQvjqf3GC
di9H5NSGwHCq/MTabWkzzY936lEHRV3xE7CGWHsjff5UDP8zFDzlRC6TLR46b63y
lQe18W+9c7dcLIqN/ysMkHXPuCL7ynCMTAM62JHHO39YwEQPN3g4Bi1LerBD+Txy
ElAEJ2FUoo9VdxJCdkUZqMe+xmV+y/wPN8grAts5bsKp+2xXPt9jM72v2stu8SD5
Ekh/cYAa+cZpHQtgxPIqY28WOYJ7lGnF4d+dQgR6eJs85i1p9mTHFxwTtnjupDmF
Wi6Q8PaoQaKkw814KVwbXY77EHnsG5PkM8l4AsMnUrm/vGalLDd5wno5ByKx4yRE
pFVDlJrCTnCsOZ5Q7sXt+ZCsUK+zMPImIl7QQq9Y+AHxp49KISVMVfG4NzARx3vI
RpMdy3+PLELwS0C2xYWHdDW1jgkOjeWNzOpVRWx9NEIvS8CMiGE9nnkSh3zECLiy
vZ3TNSkk6rTOfqr+6QS+VKxtvpxrJtne/Q5VAm1rgb7hzbgAfkxdeNLPwYRAaO38
tqmKjSl2ivDd9uVJXabLpNiSedRC3b8AADkEdnk3Zzg9qRuGU/Dctt1/Pq84xmdc
aYZ196FBAqfbuiOB+KBUl33pxy9kkNtCM3buuS0wiUI06SJzgZRblZOxjRkK9Cck
RpFCYVLelHF2dEeq5RmIOC00PcyGnC8yEZl9ET+KCARUCoa+68otF7fcnxkz6gZY
wt2sz+coAdzz29CsYHhtk+eCOzzxuHp2LA3rNQRqe+7boi82J6yR8vA6BqMB3V8m
ib//3B9ISUonXSyNw7ttxTQeVaPkqdHMbUx9jmR6q7Cec/EDPLA/uRKv3tWXM/Q8
nV2ZH9YW+mOPycG2xg8T0j1kOwQe2JtZzM3FuRqkBgCnxV9XFqlKgjJ54BJGSqr0
l6pDeh2dJNuNMhjWeIsCObJetbRjQNipmukrpIIdMGWpjf2bLO0CxmOovpIwr3AJ
dL3S6l687yRRfj3Hg/sWvI+qKYplNBLEcBCfmaOFbAvFxM57zLThOZrLKiiiX3FJ
bvC8VMarklV2DgzA/3KwkdDaoZeb7RIlM1fcbPJOJAd3valPP/CtthRJ4oyGj+O6
W2IeHpk6YlFf9P5Ze9YQEoNJZ3pCRuVbAkT1ISmZlz4EwmPWmW3aEtV/9GQPpfsh
c6gDNQWrqf8V2mm6sgOhf+4XgfKzPAvHugSqODA5rrWB5bOLM9Qs0M5bJVglp5II
u/NtCZaL1piN8Mmgb94rhXw1zlOKbzWQuuYzc72A03TIHhEZIA5vqWRMR6kvHP6y
reAnB6aJerQ3LEj3hKQEy+NasE2SqybHiVuWQA5cvDCvYU1CkhL3WQXeETgEoXRU
taPtfSNLRzLL7kEWDdpaDaY8I4sx7vTlsrpJYl9INK6A4xB/5usKuTreK5SFIvM5
HvYQsEbhjxiy085vDPakWeaIUeEXtWz/hMbayTCTXW1qvja9WU0TwjOqYHuXaia9
wNaw7Mf04TDLdZmoMI1wcY/ShkibOyXw1+9QWmbrQT+OvD6Rh2zuyTJesnKNoitY
Td5e0NERblq2AcvM7CZQ08wCjWYZ3U7mtADknctrRrBpKnNhMkp9vzb/2VtRUaly
clGQUbyXcQKYfaVuZZXD/G+JX5R0nuRARkGtCL6voTrJaSB8XfOq1rvCFykXMNH2
bfwC0DNx1eI5J5u43Gm78UdyMe93qt7Fpd3XEOc1I3lUQt/8tmQ2vIJnBSRciXNy
Qsxy3jx/i/3kFV6QFwG9i2XlpobWvbJicKYhKmY+p+vPYiIdJ3+Tk7lRg1H4JOFa
9pYmWMnn7eYC9b2KQ2VfHmOR7HSpy9zylbX0hhBHfXz4INlzY6mPNpAHWAaH/6WY
S+uWCKfMt8YD/sLTFLbmdhCFkCFzKhhmttREsKcrOVUojaTI03gqXvESF4HFh8Bj
biUNBet3SkbS3xz32NcPNMLmrqAJHIEK4ALTD5lX14qhixjd/eeHyUBIKuf0xarj
6bUdcasjmupEPaQYbibejbVPHkn8ajcKk3LNKRV1Cdr/dUqfY+LE5SQcpeNwTmKB
osNmgjS4bm9TAZmMXcIrqw==
`protect END_PROTECTED
