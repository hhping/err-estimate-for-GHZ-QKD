`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AdQRanLISz7S3ccquWzbtje+Cgs2d9B4k1xdg3PqKMsGnHg5ojd7tDooM010rfEm
CqF2Sq+9hkzYPyZeyGf6eItCWGmJEZR8HDAs8szkhq8H3dYCgIkmskQIb/Mmt9WA
1yuDJ6K0lj8VVY31sKWlNRb/0ZngH8/AOAiBmD2mvmyVW6PdIVByLNLv3lyNYxU3
uFt7Qy1mpUTT6YgsxBxZdFzvXgc0app/ZAzqJ1p675JXlbiIBu9KE9/qtbRcLC+B
L2i/2RO+ONOCjgk0s8M/WxhnlkUfMQbXDeWsFYu4UDEQIOVoi2iUJCi5ei7Y7d1N
G50nZQAP05vSlYMppOyxURGujC0iQ3U/Dt/u6cpBj7wjlloaAaHHdDRWWIxelmLd
8Fzod9Rr6oWFdZlhU+28DpPJ/Y8Fpmnv/NKZhIHL8/FgtexYfNw9WyOoIgMa4LjW
4WE/pzqsgVmSFaNoPdO+dImWKAge/D6swWvJ3sxm4ZBq5qrHLd5vVDN8tq1o77hW
S9wCEqqnX5DcTO2AgwPbJA4CIcEzWG/US1N3HWmwQhxe8uHS6RZm+qlEU4OTz600
3NlizpF3poSKtmMHskGe0H7SWmdsbyfFuwIRM5L/pIOiD1u9Dmur8Yk3UemCTfx0
`protect END_PROTECTED
