`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qsFijnw5iHMYXk4dYZ1cG5NZ0phBhkpTmoEmLfm8GbbFtrs/AYnuqAa5ssHAEdsU
isrNs6J21rZ6wP43V1SIdoEjcslcdC+ysZDPPZd7L0Y24w5ML4dffnkNSLP7ayX1
krNbFUYNC0LytuVF6V1q8cYe4iJNV7UGfalTqvpreByT4KgadVrUxEEBXyH3T/pk
lSgMRig1gogUnIcugF7iVxLWaY3ZjPgM3D8zsN/6W+Bg9Tl89ZsAT8A7JfQOsFnJ
GgNoA/KQ+Qwzmof5L2sbp9wvG2gx7XpRkMdpIt8LnGKXkfs8JCFXNcTxxJGTeknP
66rvaLjWQM5WRW1IpiI7v/wFM7dooMpGU3H6dtXlps/LOO0e5ZYBcbG0f1oA87bB
5vuTyDlgqP/+FBN4HodnTJvL8AzgyBJ+7j4/R46Cc2nQRSbzvIYxmvYLboOlAoWQ
KKnHvAsC5824NaS45chEsIrz8ZmA+nWQ9xru3VFKgR/VjPltUNg7ceHLjrN0wp92
yj3h/4da1yCvlfcGb8B83OQQ2+h/A8ROMHJEKQrqeOG39Si4rTig3HR3fullbrSA
iMT9OKQOZDy/bVyUTOOGgD+EkklUmhxq8fmyvmjzpS6Wdkyaiqd/7W7YOp/beREY
0iNpMQj9b6LdLZyTaDkDYOclItPj4XUDjNqhXKqky0emE7QbZLn//c4QjOutY9Ax
sVDxIKpZioAHDeCiZQyPD9T3nCQySbzwy8kfaxCwOPMF+VCHYu70jhhBHLfSlS59
zSWDGzIgSdXD8pjL5NV9bWFFbtT4+dTYBZjJ99bQ0oFLdDkTVD1uf0ZR1he5L0Pw
yUxKNrryPjpk22lYSNfcFV7gJCB8hS5t4clRpLJTB2JBw8H0zMLdqBSPXwdR1xl5
THCsFcVrVtRq92WsZ61hyX2PZloflRmAkAY0wfLbxFlA6MCUZn68c4uVWTp0a93T
7WSEPGgqTfJuImvNgNZdwJMa8zcbIQ+VxNB88QnDAeaN/brqskE/3lHrp3WTbdNq
ndXBIYL0iCNSJIOH361MTbVUeZ1wrmULyb6Rlt6wLIQ9DN5mJOsWWyz72U2wXAsQ
q/tNgntM5bTkf+2znfp491z6UPlE3PvIVA27VSw2jaYX3tSqqIBId61rD6y9kvwG
U2uTBtt/IOlSNB7rPbPBcy4J9etHUTx/He+a2VpirNe+BfncFo7VSadBtUGXiHFD
mhZGQjuGpC5Ye56YQJNM+RmxoCO84zKuCokIT1IxG3o/WLCLy0xN61d4E5ube/cD
aQ+MKfAAuPJVpApZHn+UdwpFaeDSx5uYM+DanaFbLTlFmsfIngKqwp3Ph1CVydv0
DFgbzzp0lwmUt9F3eemU20pkiTHOY6ifbHd5l+qaFHKHTCl+LNKDv0vSP0aO+7gJ
vny1FKMJyGEtemRssOs/7CRzSecFstzgtdlzuDuio7XVTqJD6in8LZoVmRuLoi1y
zLFqI2eT5kvXSzNO968TVv6GiSUhTIYpy+PxX0X4c4YfQqWvwSdeyJtgTA6jMdvj
WhSpKIMkiSUL1t9jttbAx9DR3QUOHnINJPnrTMJzJAnbQLaFYQLlZ/9Q2Yiiz5Cq
/LYFcSHBNWASxaWMEr0+RCXeVwchi0e8T7KyawJ/BbhyIg9GmCpjZKJwYlrVDXQZ
L5cLguisRCvuPKdcfa8NeAFNgQTAn78jWAm7DDar0mohkQQPHrtyujgu52iI9sAV
/TWvG+hlePuCmkV+xCYUzSQVmpv+xGD0I+d2FazybRfHGGtAUAYQLtJv0201ZF3y
o0OMO8y/bhLUI98Cmy0g6o2fqRs6C18mGTI+8905DDG4Cj8C4gMIttmsjDvxDE3q
/CRkLP+VZAHd9567CYoySH3yPnBEnZGccHfRjL+BraHUmEm5s8mlB7CYNwvbo/2t
G2yl01cbNymE2uhuRrdBKYHIUizlCIFwoD5IajIMWpfmdVaCGzCq8Y0iuma0tyGU
LsTyZTxiQZrmeXwPTvhnBdGy0mnpW0ZMWStpo7c+ovbYalH7oB+EJcnMgbz+lVmR
pzzx60ewg0UndSieCezkXXplJwTkkrLMjO4zQZNBOeWhKHOf6abwevhMFGtJvrWD
6hCkLySmmbXleSqNK1uyxqNLtkZ/KG8cZ/ZIM67/URDqDxxze9vsld1f9U9elUB/
G0efrRGGnY/IPU2YJMtoAlSV6TOZsivmgjI1uPm45iXy1CTvFjhs2WpQlyi6AShK
RFolZWkYCU5vsccBa5FfEqrWKhemnfN3FUz//NzAVC6a2CwzHKnY7YRbL0LbJL/k
QW+vELwVqHyvo5SpFqyuTH4nNuySDzO/xRdGjtH1dHCOnK/5K5QHaJlQ9pqL8Lvt
yy06xw5PHPEiCdbCGv6K7DskgSWogZisKo1OG1jz/VXHhHcTIAPf+xS+Lsy+wUSZ
P77vQgX1ARmi9QAHr92m6EtCe0zIEG0GHKMttqrf0gKEJtMz95EZL/KfOMZXyLJk
dJYrp4o5OwfAdITvxrDIgAnK1/TdYAWyfZtFjFSJtNXTQJK/sIBkrhqlcACr6E/3
LF6gpJJ1ZntCxqvNXop91vcifTQ64MyIyzj5BydCkVXyWoMM8iCW4oe2dPQnskiE
gbKjOOvwcFCy0QsidNYYjFpaim2+vj3fzEwaJnxCI5jWAe/XpH1JI8l76O1tfBis
Mz9CdaumFtd2QpkhdFYELCif27Hw7O899kGhSy2ZemYNgCiMocPI3DDGXQaiM7Op
hd6gbbZyQJ+WQ15bkuA46wN5xEodL2F/4HEr3kpF/gA0xr/lK3BaQjW4A8dBs+Ib
uNdGMGqcf7n10p1aGEuL0Txiuf4lq+25j8BtE2Q1uuGRCzc2oDkI74gt8KDjUALG
Gy4HmM5vD+9C8/r5WKhLD5w8z+M12rgOsY/A9Imxie7jnknJ9YT1iFOYJGAnmbe2
sG4xxhGLCQ2B0DCZiPPUG+W2S6u6cYAxdJC7fug+HGWk+BYmBMiNXsh7wkjxuWyQ
xsc9z0WQe4yCS72MYJf9DHg4p+v65HDsWAWEh3oWKATTfF9uziXn5/WZKnVMHVQZ
pAFcaEExqJJbe3LlIMXwrhqI6WTWu9wyjss9Or4EljRLC1kMRBvFtWRfMERaSCCj
z24IHGxt1mbvh3zfhhg8m56PGT0Yoa1JCnKZ3rENHfjxiXeMWZZQYh/nWuUubkNu
+q3OhRDOSOfKX6fBGwZJxVULDPoNyfgXbMQyzlMoTE42mYh3ZWS3/QL1xCu0OrJJ
fV+UipI9Oi8qMwWPan4tAQBKOPm8l9ax2zMm2gxsw3tRacFxi8iVEKROhKb3OSkb
ErhCTVLVo5s8wQVjMN3m+FtpclJ3uyJMO8vEXyTZ4ZgLjChonfbYO7ylDSB5lweH
okjvDYDQHwomatkk6vTY/CuqMQ6gnL8eLqsH+4rSnAzMl4USs7ayLyo3Qd6DGzqf
UOvZ04VciO9NBYX5P2Yxkhl5uH05Y57MA4tCh1hAYidlKUD3nCA5gzwEc/E6MdVN
ov1qceZDXywoGWEhFvLyQwLnbuOE7Vpfu5cNvCj8aDDnp6RcyLwn3eYCOJjNThEV
RjTYrgFkmkHdXPCt9/YUPJfm53/PNLboqgF7XZYQSPk0k2BQVqHvUH1daQzPtc/6
G7d0clrR/ym3BNrpFRmPVfSQ+UXmjHqcUYlvduyNU9Rzg9ZfF0KR00oN/cv0U0y/
810ABwaKQ1SBuMUifJSHC3sP6KufxIm0iXDemSSyX83DZBCqjlXusVfDz+iaVDRP
q7755en8QPNoF3q2dFYiqvak+KmbPjEbPa8dFM2MqJMNqDfqgqjhpPSNVG+y2mvY
ZAW0hXK0DEHNm9DvDGTdOQ++FNV3Ipru9D6Jd1u03e1/g/325cOn47A7fej08ukV
LDquMU3A1fTmvv6jSwa0uyM1Af7ZFpiqBFC8PCTWbKVg0uIlypCT5xWisOnu1SjM
oFEdBiUzZBCWjfIql25zmksDtuKo9jvAUV8jBank51MtfdTI2o+SL+PJIs7EeOiz
ebQreb4rXp8Wg8hnAOlMZEpUdRLgnlZ1BS3UYFT/JCzHCl5R9aFF4WwHZtHUaCbz
eOePw8QfJKgCp6aABoVk+GZoMIiXxG9gbE1oPZjxqNQrj6IIWO7qfg2Qnbv2xAWt
PDe9GV8zg4wNRH73o9tMJT+5AWf9xMRtvByKfNqVajJ20CV4arhI6ZCnGGE3SL5i
cD28FfC2uTq2VdWNnAbxEh63j6JvEiTftmmsWyQ4Mxeu+5FvcS3/O9RmCGN08bZP
Lob5H8TtJ1o8Es/ompFjQkVpqNrng3JLijN2PINEL5184T+oCb3VGYODp3mYc17Q
mJHVmW7FmMDESbCc9kAV914szsfwtQ2VbMtevIfxtrEzkLPIoVq8bpajPdNsRSr+
Gc4ZwXudwX/cQfxiV0hilJ32tK2f7P52Nud/Yd1NaQT7iOetAWTOaAuNhiLaES4o
3HtXTtMlc9EWWSDfJzG4r6EUTx4KB/ycnFvNMskjqFP3xtVzy/B9HiasExKLORTT
SYBDCH8T7Lw12XrBBJYYax4NH4Yauw0yNzdXH4otjs7vrDA0rSj8lniHSkkxcd+M
7ySBRwX7Dkxvbq2nuKPcGRPQW5+FIAsd1dBVmlXdR2kZjb4N+tjGlvsORkd4KIbg
ZRt+qOJNdlxcW0TYnKtkqibcidobQjOANkoXap0tv7HyHpR3uXg4LIjh1PYRwwrB
g79nN05+BW+a6lddU1c4nd9ZiK/4BMDJFh9hjY47UZQi3SCG/UWqt9uVQdRoja/N
veruENav5H7eDbOFH6JV3ik//rjqQQ2vJN7d7Z3To1zb/JXdWlgbeGNUL9hW9aAg
e7azkWcJMrfXkXclSahl2C5YOaagcV1Uxsj2x1Ei3o4qTc7PjVpY6y6B45c6PYaQ
mqj6bW9Yi3XaX7CjB8rheoMMWuSTgxbIOAgiW/n4+mFzmxZIR7/grS0zhmlc3Cuy
xwuwCI2DF/Fq0w9sKDcKWBlkF/9rrg4lC7X4gl3a/JlejwwxthqVHvV+2cXi9IiI
LRKzquh6Xouc5pLNLbnvXerPLZxItOU5EpBDJ60QTl2efRdyVD96goPiPqYUeLJ+
TJoYRcsZRNPMRB1ojcfEj4Ou/wMdpqwtB0fUorLylRX5W9Dop5ICks9N5Pw78e2K
HJgIVR/PM32y9lrJtMj952Ep9J4YV2Ewazzncg11mQRG8yfqVoTHmFhmTdeUZFVD
pPBRcydkTIH9aXDGFYy9WKCd5OT6X0CPo1mscxHoHk1/UMF18AofWUYACtf9vAw2
2+4iVE77u6q/1PsMSbJ0CqD/ew6UZZvMl9sH5Sz6laHnzni0j041hRLrXqjwku8g
hknDUzc4QLoTQ1MkPuaBVhDQAS8TX83S3gCU5TuN7dl/YIrSOyH2Y5SiaCtWPM7J
w61kvtciYnzJwvac2Dv8HqMdRHTbejQM/42NtIBhm+YzwOlUfH2gBh5hzxWw4IeM
KkEBQHTmz26hfNzKV6wXHMO7WFTGgkuw8SHP+qpz1Knspj2YzbSmQ5P6uaR7Y8nP
y+SsBa9PvRCuma5CNPgAzfCCln7bazYZ9IGLN7PJUwtXKBV43H+9xoxvnq1MoubO
tUJAZwEWKOQcZyO0U0LPlC2OECeQDRYCLEBOt3URykk7ZX93itgzuyVciesUhB48
QqbF9WuPAgGB/k5BbSTjMKruwOdgE+mRa+Y1j4ufnKJUvjTgmJAmN2USGsczbZ9o
iBGTmRyL1Yhmo3lKUh8hCXeBusZwtYDjt4iM08LAbIltnF3JonIrr8+eBnpQufpE
39/jVS63sBFX3VSTRlioUbufqqr1ES2qNhLhOdw7A/QVCMd8nHz+ufz2sW3JwDo6
pmt04bVf9x2sGwZBPUI7CzwXfw4SMCz9QVnw03cmyUx+wQcDLcaHZWaSd9HRQ/Av
pjXGT1O2N27+zPhVs/8cj/n0cc8wKFb1qJ0SDsu1qcSxHYRrQ82GnrCpaDaYzd5b
4GFX63QuTc01oTuR7+u8gZFF2XPAyl5Lk2IpgAPvEK2lTUmnG73EQVvbXqk9tg15
FZ7M1fGlpPFJ7rqYPw4tO0Zchz9MlyJZIEMUMK3uCQajA/me+/w98bhX9SabGhEe
XVRlrQqZRMnF4j3UqzsVsvB2QY0AIAcVwaFI3kop9Q8IIbwFvdQdxG2zQchqq4J5
+ZHwakRW2aX0cMIP3cN7hixAiFBd8Rzd5TMpN+4ojeq+f91VTGZn3XUpvaFHoOTs
df6p2dd2t/7An8RzSKb1IFS2lUDLK+7BsZjUvsjhMHcpCjvtVnoRj3cllJO96FE9
oUQ0VUajTbl1FH+nLnHtGaeuCiZXELHVCk2UX9ekfB+uVY6g8uRO4IyzJUT41Ung
XMye7z0Q+VUZrkpx8KgKUmwtJ42HaAqmTHYhJEvD4saLbt1ALEo2xc1ffHGDac6N
ro2WkHgw8aVahqE4bZWB6AcxfKj8x/r8pClPxeBLTeqnf7ONjqacuzUMwjl+zZ99
HNTT7VRtNcteerPrJiQ0n9IJNy/tNTRFXVTwZdgHyx6gk7fFKgJSH3kznv9TqPsh
PrGt/YSVvTh4bo6tolUayaN/9jJnhaRk3hn09FTbZCqLE9uY7NHiLvc0kjR8mErx
vDf1ZwskdhX0gXEL30k8DrOWqG1Rdu8FwBCkXaSmlQlv4sExirf4NhRmZnU/zzAR
ys1yHt5Iz+4XrFiLib2MKR/jhlEAJfvfDQROYy3BjqvadQ/DJXJm9dQI8vw2opXS
5YMcsaAOpodJJCItoRQrev5XjqOaQLR0d1M/B0kHgJRBgeltHWfkK1j30n2BG1+l
LaZPY896k+XBQvBi+LE4bIEcud6QAOM2t/WxgVpTdRIgNMuYHxUm25DsbYqi+L2j
O4uNwzu09ypc8VXb2rawI3xZwE4YL959wyC7ZcqWFIrlgtyXBf3pv6BOMlfHdCHc
tz8cLOgVfmihH9BVMTiZnS9PvbUYGU7MpAXPDHr5iKn53dQxjTVFF+skzclH1WSY
usk+aIFgo+s+ZIDGGGyRpxllrhdOQwG2ZpmAb28AyaoWqP89G6LRU6BMCPNINs0u
amGmAnHH/CiZ49DROKfhByXwgSJplMNLM8VsUSfjvF6CeDKDCtYlg80qlc2i+A6h
YpJdoby5HCv99DF5Sve5/UCY67sUfavFbgDaNryfi/oMV4U1rl/hLT/rXGDilzU+
zLYr0eupNw3INVf7RMkhOUq4+4Zh0prnEj5yoB/rfwz5pmNTf9PQ10laV+GSVisp
Sl1+oheDccQP9qgmbSwlJfRm6yB20G8Z9rID1Ey//j/DlnyqxazTadsU8XMBL/HM
N3nQkZn+DudpPqIHEuJf9PGMQT6w9NPUfrWlArQeQFC2gc0PDjugaO39PGi4Q04Z
X+8dc4qFyFADtpIa5a8ggnZbllCS4MMOktlBZQ7maJqUpicu9gsaBJqcRk/TfQCR
2ufo+sHrHJuAkV1kcmoCYko5q3X60ZOG1IcS29Owf2FcoxdwlbYoeBTQZZO49gq8
8QLXflukJd6qaGOhajxJ1AAsqNLCiG2WovcaB9EFMAkj/emWA0R3e8oM9+h3kG1M
gn8AlL/LpXflUoCLV4/pwGsYFJIYoTDDxAfTLYtvxYi060gZAXmPVWf2WPar2fAV
Rddg92gIphWz17QCCMd8+uTbmLHsKzNlekiGRM/xtWcppDrOI6rwZ4bCiialmVlK
ZNbp8Zia+ceJxygnoMuO23FZaR5dFDsOyU1Yb+8oll/6G1jc5c45YzEPPRqJfua9
ktGQ6d6mxMvef56w3PwqYELMXJd4PDHyh+cNx4lUogeFBDUlgmA79UMzZvBk3G0W
qDu8vTzFKhn2DCcEAmD1oGq4hfhwYF7vNJm6N2vlE17d5T5RwMwN+qe8nSApocUx
2jbDPZ6w1BjbqZFSKLr7ijQpPC+0a5MyYjB9WmUVQVFzUkb5NZtFoy8fCGJE/xum
G0vTHFBIliOxcddvAFstVfkEtkNc5RQ+sk4b0hwdB9clQ7gRiOJ9NX9zKsVC5MS6
pauxx7LBx1UqniXwq5TVcPMfS4Qe5mg00PTURM9bc10BStsvldl/ETzgs5rrgbr4
MkbS3uAe9VK4iM4SvNyRPkpXUj1SeminHonvHg6jizw4Xxt/Foa4t3KflJEcOvjB
CzkCJmxI5zaGNaTQqrdSdrVd+jPBcZTq80EMF06784/uKtIk194+qs+OFNzdyW7n
kDkaiF4CWa8o3Lk8E0iygO51Kcb9fB9fxukSx3WIdoXRKvNTXcwQ/WPlig6r60FO
TrpoWWsVCxP8ITOu7YvHiIGsJIR5B+PjgfNFMu8dqmMZxnQObCcWhZS3lw28l6hO
rkmTlFqUeNy2G9kmEmQzQ8O+kYrZD3iXWIhpHtgogYIZXfRRbWrTHG/J/9GcbRrc
oWBtfQKOSt+qlt5RcF0i9IBuReYlshbOCChO5DWwZ2o0T2w9JZx7G0FqbesDVHub
uW0lFJsUN/m/rgZEMvULMELanVmAdcewrrRuE1h36aSe9ykBzvD2sizj2bZKCvQM
BcinPrFo/c6WbeuEpQzcRh91F0vOb7TWDWSvi9J4cLSzSE2cYkDI7XK69jKYrmg4
rGjb2buemBD2HtBTYGk8pHuelgUhDIh7st3NYM/EiOH76b4gtzfdoeJXthkf+D5Y
nqv2C6YuKS4Gjg9oH9peIS9yTjnPj2LWiQD4kMBL7NWrpUS0UDyjzak/QtP7ojRI
l3xO6xes0ItXhgVC/atGvxhX8dD4CDKei6q8KPBf/2Lmsjdz3tOmmB9TqquU1lLu
sqwd3NMwFPnUkJFkXilN4vPfe9952XjRV3qi4NcoR1xj2O6ct0Yf0brQogTECUlP
KTJH0Y9ihI6skumCKDE6erbe+6Ewqku5zQ21GJ41xmES5vqczFrKfq7XXoBtrVVR
+cb2gS+eTHUOIFojmh2qZV0w+TAHd3G8P41ocDDAeKwbawXeelJIKhvsolsiDwu9
4wBinrH3eEtlpLEav2VrhuuUB8hXNDrni5cANYQd9JF0Ftl48Nq4jVX6owmZcUqR
1OHEeolrE4+8wBXX8yBnHILH6EdCwEyVbjC20AkridwDQadVTkgqn6gwkUesAYBZ
vfoZQhiE0WUBHqoWkn5xF3Fn8+geA7DQMBQ4hVhAr9OwKSTqGjhybhG08f/yux9f
DC+awPsPbYFjHnj1XvbQsTE+WiSuMfzo6qUjDI7shEisRJi86hQnMrqlqDmAqTMH
kS4zFGUe1LZYPO2FgpR26dq11bYt3av3M6nfY1UQZi9LBgeIzk7n+JB5o5T4dNmP
uRK20iQGSknCh/o+YfwxUn4VDaTyTrD+vh6Q+UtQR3rR4IlG09wW7VlzxEQEkCvB
hN+3DGLEMXNinrMzIq7sfmx35t0TMS47s4/aKPIYwhRbP5IuKl62+tFh23xk/2xN
+TJEBrlOt4VeZqI/u7SqDsOdATFVFc5ssyJQqXCH/7f0PJOy7pKR2m9Kx7bcH9pU
ECVzIIlUibQuBeqAwVSFSH5kFPhwkmGEsznRHiQjLaWsizt+qtdK3dx88TlKtT3Z
6S+kfolial4mYoRtrxNPATofgHAhDQNaIGEnQTMFUrkLiDDFjClHKIb/nn1ViROF
6Yi1fJmcTfIOYM1jv77rvJIzmiRxWHRp2HwqEls+iEbnn6O8WTkI/CcaDA0R9fr7
PgSgy+svicZC50TA+rdGqSgB1aAwNqqV+ouMihlftWLNhTL3Aht6bwWv+J2jjEdV
5PaiqXCETJOwOzVT1f94REfQ3hdSgAY8F2XBil1SmHHp5cSHCMccTwso1ABaxyZS
8efU9laFdGIXbrpnH0gg50/tHxs4Ls7l+92rnFoW5mWuSG69hoIyUdCd27J2ZuqT
dW0nGR6r1H1OQC7KTdjxGNGaoQfiInzNOEgd1/GsLmFK6KhIH65s0NJ8sfJ8307W
Omy3OzA3NwY8TaLb7M5Ut5H9qi4DTeqzcx2gslZX4vM1zBBIlkXRTaAgQ0pLtErp
U3aSWxlVjPpvyTDcWHkz/lhJ/YdzKr2ZF+jyas5Vr8BeKaqTpaKXv4e/iXJLML5B
5HjAP5FJT4AT/eA7iv2lEsDq4sgV4fe66s/4DeOK+ZuI2vQdENT8bQHm12wuyomV
5okea4E5YpYcuNjtgbiUa13wafSYgYg2kinG9sh9hEEEq9NXaqHY+i/L+uTEAb0Q
WP0yzw4p4vThURzxth3KUT3G+kERQl74Buc7USowdj4moaRAeJ2zYpg0+832NUTt
jrMD3M9uPs5PKrGMQ/4t4XH40hMX1mxhco8yHpwTstwCyeDFD/3U5NhMbXJf3P+i
ZXxVIS7qsADpffygZHmwsyMtqLKj9JqIQREPljnXp/M44crMPETWLNkmSzHG8L4R
yrYlS75fWTSv0YIeseulqCEwLDtdouOZ9XFr78tN3FLllkoSlXtEEbVSVQ6nRhix
L1TVPoP3p6/HoAonMMyHyGKXVosHY0x4DF3ilnMH/OWM6jT5L9Q5t63Y28X77Gr9
7nB7qRI0pUxlscoQG6fO8T5A07Q3yo/oaefozVGpMbhYd7Ci7J24K22Pjfz9gQnp
F06kTfWcIVKeVRqa9KVhoRRS56aFtpnRoG4DACQnRFW1BUbb0K4ogpn2vzpCydQv
fqiHUpze5D2OfEt/SVPVtpHkgNDgub4ETNC80dXcPyQNJI7jWw/QIFCMp9NJpDag
1xus8CWNxMY0zJGd4SZ5RiyJ0StXrACf7EmjCs0CHVGcwoxenJZau8oa15kjP2Sj
33F6oWXQCtO8udyWa59uc0dd0s/FNd+dyiPs4oW5n6r8/BjViT7k6ie00lJWcvU+
QtmMN95j6SM4zM4TmlbMVR9u9tnU/97l/E2MYeUhDtMen5twurZ/rzL3Om6iTPbZ
4VdPva3Mb2bUy5H9mSDhsgthlHlOru8cYP7TLFepCFfnLhVPlwnM6iaLKf86aktr
ytW+0wiw0fGwRiNFhOcErtCbbbZUKxHX9EsRopemvqPtHNU8VWxxy7uG5aMC6Ba0
4BEDBPiQPB2u+/kPhjvEwk1uFs1LIkRioY23vQ3eePAN33LN1FNBtDwVKxc+6X3O
hcN0wlKsNuiyQcRXEyx23zdth8wyIF+2HuZ7poc9z+6j7cVWkYZD5F9NRtrXE2kU
qBg6RjYSZJa2RpB+FhDyTXbTJW+TEo3EJ8sSziYM/zLXapmqFqvBUpSPXQO6U7aH
k5HNgn/eLgsbqGJVCk+b/fNH5eF9zYZO4bt0bZiUTMGd7PZDnUbuOPDJAR0GLP4g
kMGk4WOSaFbR7PKL7K4rkkWg1a91VVYOW4CuQtBNfrLIDHircYmvKQAHPOrPfyby
x+yoUtGIUt2+b4nf3Iw7WUsuI9I8RQOO1Twxk16R7iRSJb4OCGgA9zaef5+zlRry
ONPY+1xrywzgzOMibcUHP9RwYz2WMNzjTE5vsG6cvoFmmxQ3jjjMalf98ZO89zdz
7DkwMnlMXuG0tdjHwaq4roOUJE1L/Q8Q+zzDLIvBPvEU3kGM25l6qX4akmbGJx2o
CMDRhISikNwKHcofb8l8o36Z+WPXYark4VN0SvS4QYcSa3wJeZwz/DbQHVMBLqyV
A8sPpvgPVEoFqZ/t7iUAIwJpIx4iic4XPfVQHI4KTpnxL2TAkscIr4OCF41oSxyK
nUXAQzYufdP1sZ7lggvNbVvc155H/Ro5TdeHpJyQVgUm24CblWH3GlKJgBLfX9Km
+UmIa0ckAwczRII2MrbiHQrj+yGlZs7qt5o3QbrbQErK6Zckdxt7JHXTeIec0MWy
nCUNSiVYvC8tGeYD0sXc9nBpbpyTTTDWW7rui32EO+pyS+pzj2O0Ians80tCvleK
I07dYO31UgDpcpBgTZ7u710cX1XwZdmggB2HI/WAwf33WC/rzvhmzYiw0o6fS+JL
Z2WPwE8QLIqrnblfiiH4T1bQyGQ+7MxHzBlKG6XGlYELi6aQDPyBo5zrXwgRCOsW
s5ig1GTU0iEt3hKccspJ0v5ehrP5dtH9YgJ3JJeUPorhfra+F9cujvlZQ19V0+pn
q9cxpZ1uWGBYoZfrPTDbsdcyYVl2sgXySaKzzbUp4Rry5gkES+Q0RyMti7gFFYpk
0ySRVEKCQvHMHR2pRGAcX41uJLCEJx0JBik/o8SlhdImwH+hbFcjkzEvjdvlCh5S
6wMzt+W5jL4WlDScnyGmoDgFDiPFga/CLkjv1q9mihuFVXHEQAifB5Yi28da5dmG
UnX5f5KqvfALbARrR3bth5oXUDgc+RSfqiHqMif+GfmIjAlwVxQ+jeeGRobQTe4f
fKususbpEUOWMx9em7+mp0ZMHShguKTCTbHlXFdOppyiOfgb5I6zOZ6dkYVBCHpU
I38xdBLPMofAqaQt2Ykt+PtIECDGERQ8t5kELsK235iG8ecMEkzA+xIwQDFotWkP
rCmAkEJ/22m0ba9Zj2xQVIWGVLw2sqLYMOGcwXjaNoL70xUkKQZcnwCbsGd58HtI
pdfeCPZyksHdZy80w5D1DNVqoKCJwBXyQO1uYTb/+nKTa/J6f0W6OngCMStX/TdH
yGtN9GJefntP9S6k0pfCLNzMxTHC8kYbIANM98EU3SuzRdF1EuiY7/jY3QnC/s1p
72X6cReoVf802G3txE802HsdKs705ooRnSeo4jcR3xVoiCWaqNwTbTR49h6o8usK
DYJ1dv/26Pw9Ra3XeclNvyRgiCNQ41UQyJ8tJ31hKptRSoT6x/yvrnpGskjaKJir
7FGIN2xwnkJ7LFbUa6DKmZuvPf5naMep1YlZslVgyjEaUre1U88Fx59Xq4wZvcOo
xLT9PXc/nbeX2rL5+MyE42GGk3EzXiSFhjPhHIQe2NyyLWbARe4cNmlLFOJZYybB
aC9IzU+DwsAeVprYIF42k+7JaSdqszeLdMCDsXo8GGDRvcNHZ1agN44MMSWP3xAJ
X+nTGHIxbNuHeMePvB9vtp6zoqMbOEpRUqNXxQaBJKtr2nRr8E9pqK8KwRBIalNZ
mfcpnPlaTiPCuuk9tsQW1KWiHGUVtTIffxf6xGkhlp/pi1q1deYDsuXgGWCuZnw8
VXYfLhbg97NBs98lfRaoy6/I3N6mhNYJlKGAxRO6nbQf8iKOqxeBr8GT8/QMiBLU
YcY3reeN25NSpwmf2dLPuew0q5XxQbAeDlnEtowYwTJ4OjUnmhT6bwk4bpfNAEN2
d1N7HwcWklYnZWkoTOlPBdoFdLysCEv5yI/Gs9EXOsW//12H5K1/E9ouaTLGg2pn
S0SIG0tRPRSogY1oVKo9kOxvavX6Xe567bGvnPls3lhpYpFoGyJMo/oWG08Ud/CW
RjVkljN4EwRHr5Fpb2mQ4dPFn1GW7yI+l+zsq19nU3oJ6rhGBivttRK9nD4df+aO
LVo+8sxMlmJYctCBKuDiVwz3OZfaVRF3oaswIcJQnnnEh4dOlQdMndzV+E5rNYDs
a7+WaJ7WFxJrt5ycTjDVgbzB+oxn3rRmMnK8Dd1Xa6Ws2tyKwIbn1h/VuypZ+2aC
edjPPodjLQPiVUPyyZfXPLKQhVtZ0z86PpOQv4PJhApsGHZFKWsmMvWBzaH2vrfb
92cwDh1DvJSw59j/05Tr2ELxY7ECB+OOUekElS/TGw+4pwJ07zoMt7o7XXFlVhUK
hquL1mwnNEPhidiPY1iquUoAXQDgGJQTEvIw3vuUHwB+73e3kZD4fHYZvPsmUME+
h7f+DiQ3Cfo760qIFtMYOc/YitpPNKUdLdAa2viHsDXGLGIDbYI7JGrr/ds8vhMZ
eILfMF34bJkbBoquqMnZtiIbnaoHdgJ2Sl8zuQtg0usoRO63+8MBlg+cG9cZsB7V
t2Sq237gmqpDFeiWbvV53t5RGeKXAZIjjR04ziwfIOST+DpRrZo/ppCnYQnnvrW7
SwkMC8iy2LmXdZBlU0J2Aq6xJHszAnD/M9IHS+9CwqI2RYNXsw0yh8tuNcoXSJfs
miZeYmzQCQyMPUUneu7nzCa8vFq7tDTkOoWM3KCXrNYm/WpPZWhdsVCVFc2MlcS0
6qh7Pr1G1WQz/CGhwo1qFvOzlv0RXr3RSOnIM8G/JZTC5aDgurGnJfT4VEGpxZf/
sctmT16fVssCZ5Z9G4mZRAd9vswH8czMqnPuXr20Z/zuBwq5VH2EZSxVkhHY8/Tx
BJff6xTVIJyC1tIwX8BRG6oUsLP+U1KSfq4V7UcfcNPmTMNZN9L5qIf/E5JSuMO3
qbsHW/FZ6z3E2t5UlqNLTXNXfvdbrW23hWr5hzryBWguGvTm7AC+oyOqIRBYwk/9
FiHtJ9oEsE3uiIsIKv/BlBxfi2WDsUkgeyZGSNzjnkz4AkP09KEySQkaUNq/xJJ1
KmycJYmZ3MEVsx+3UASu7swr8IsLpqP9rUdj9hOyv4Wt6uYKrdnTSLFzSCcaJ3cC
7DSYcELmXPBlXF2OyBlWIG0fvGOYsfcaVTGnvTgYmsBsOrR70dvqZIswhEXGircJ
H3oQwwyFs+AC4pO3o5gLPq2NVS8LSPPtZc4bX/o/j2mupamqe2MBY5KmQ4/ivgfJ
AnglM+KSeX21wjxL6JA2XXy7xhbQI8oI9Zfn/6kshzu1TcDvItBr/lT89OfENhfg
WHsCnJFw7cCK4J0TtljC8qEs6KBlhA2wOpDx/9KU+pYxCzsFz/fnvltKYhNVoc4Y
VVvt2HeG5Ha0/cuG9iSB/rvg8XaF3QbN5CYnNq4sJ5k2q71UjffcgABmWEyM7R4M
w3vTvsVckAqyXXUhpWIXGX5mwa0TiQmv/nFqAHLn58MkQ+PSXWNoWiaTBlVUOkNS
0Gfk19ZsP1/UVaXB9qbX+C8yo3IcU2RtytMjgpMZ7w1FZuZnJjmHkYM/tRUkNVm1
FpH5xkSplpuoEVS4b9hj/yWm+2VpmeIfjCeg9onqMkhlD5wRay3iZRjY+B6h8RPX
Y07sUJEcSzEZC9AI47p0yRZKQkwgh8oKqsDX2M22dfKdZcDsZ2CGR499VYkTs1O7
892eubOvEv/nzcSJgt3L2OzX72WlBvUaEp2pI89BNdeLW2J6DEMERwcdl8jMhWcr
tA3ov9DmkPE3cNp8I9a8MV8QgSVE0sDZama006QcmC0Omb72W047hvFu4NjEqlsq
zc8LjcX7dNWALePwQOWlPn2wLwgwCC3iMuurGl2MbojWW3h2fWXKx6F2YppP+O5K
9RtyZyDmrvJtHxitAAcqpwfPeBaxA8OivDo4s6GJwrU599nKCoyHqBS0KhiG/mm7
qz+K4YUJY5C85Ifr2hc1jXvV1h+0AHFhDgWaV0l8g/Ne6gg8x4/UpjeI0jxCOZHQ
shGRHeT8Nih8G+cxNGRt+OIrJ60Lrq68XKGP8jynzIdwvrd/QuWbl+4aLvSyLlTZ
OUZfAO9yG8doM+YZEI8TcmVpJVZ33x831nEz5yR1x27GQzo6cMzssb6xEKG0PVGA
btMmk4SQYiT76YgL3+rXB3JtqY+hoBb5VJu7B6UtghjOg28cnbQLPZlTBO5U/JDG
ZEo7g3kXcTA1Pljh7ACu5tVihQEUPb7MjABz9sEMV7a9XmAVOQZdW7VFFL4DpyXq
UVNQV0jM9wnia9kpJNFiebogI6VQcNv8Kh6fQtCFB+DQZQxh1UvMYJHY6ijFc+Hz
ludytipgOlrLLHpM7f9o6D8RfNE0EOhkNmXTPtgPrtHxBwJAkESTQ7vW95bOGPYs
9iodMkBK1pCRwCK7LkXmrwimMCYIiTG/UMFf/f/UemqLTmPDiTqrnqWyO59nLUL0
o/pOr1jTfcDalANc94XvnCRUZSuHfph8+OhB4y9xBtscw56/bruBckK7s7i5B/W7
226IXoLBAgLboWQmLXE846CByxic86veAukHqF8eeTNfG39hFtx/2xAY2p7fvcRk
Qhi0bau2Y3DywunmHCbc2dr3+ZT0P6Kdg2giPSWpVw8HGM7p7ZpoxuD7jMIRh0Pw
+yyfyfG3fIp6Q8qhqavSPwdy+a1mUq+mq67s3ucP28WsjIGROcjJkmHylmfDHfUW
Z+vGJX+89PjGU4Fv5woSMzEMcnq5cQ9lz/eKMe7ZaWkGEqiWIRb23RClc1cNia7F
MjS1neWpjd/Pt9El8a6wD6WcTc8icrUBQk6q30qMOZVwf5O5MgW4EFLuS9Eddfi0
S3Sg/VXi0Ds2dHUf4B4uHGkmLack3vYBmtk0H7mmyjf6wHuso7rloTT1Qqu+mgQu
Vm/TIeLRKt0C9NIUQfkWbf8N4p6+gIbV16TPxWZWxGTz5f09s5VqnlM5RvH7nG4F
OmEVA6v+UfBT8SIz4x2RhM6GiqLaExZs2fBn1GXBNHyZ504qPkPR2QhdcDYFUDbP
RHAhQJ6bfUsXvXFNdI3cUZtVCzpRHhtFdfm0lm/lRn+PHFclUmQOwEMXhahf61Z+
LEQrsXyqMBXM5KUPY1RYs6vDsfGDhBLv7yAwnqjzZ6ap/V0H6ATQznxXiAGLLGcY
5CVGEPGMCtY2Qep0WKVa1SXQAXnMoyVr65mNEAK0TEPl+WQlbjLXRS3HhvyvR6SM
QuuHIyZqSd6C0vgB7vRjIkMKJsqBjFpewtw2MCqnk2flw6l5vw+G7B5Xw2jNscV6
x9HEx7ur9hg/fx1VuAlyi//Gsoq2g7hNmew4FG93r+FYRyqCzVn0zVOY9wZwKBL3
UkZU+AoaOeMBcIgKGnfRrcSwu51cKLTTXS3otEn8sfvOsFb53JLLYdvM2JJAU1Jb
78yaV5jMd0jbMJong5ZJcK22cmEdaP5nD6/SlSCR96qienKvSit9lrKZovniJnEp
eod9N9UBFntzD0fuUyFS6vuEW5x4ulVMOdSYkQnrkW3dx0prGT0mMYSg3aV9PclC
O2AEwPUYqAVwXSNfvzLtxXQs61avEslmHXHDQjOBLGntd1mnyRsJr+tBl78eMzvM
3aK8HlZQdxEeUnocbNbX0F4k4lCVfj2gEGJxUOcoXwkkexyU8UY5io/7Eu9ZKxKI
RgGx3lZbYEIu4aCgZAw/IMsq65TzAoNWD5ik55VwXWPPGcJKlrWS2qmzPRyalrJN
LCC1dgGLScqbKFJL46/qnJL4N8+vKxbdBwdUWd3wJjbBfVpJGO3U5R+2a4pWFp7c
5GStFfGmZEBv1Cl/y65Xdh/iQ1BtppjWe3bmBezYTSfAmfx3cebbslBkxgXFI2Tt
9RHBrS7yYjuO+Svad+PJRawwqgRVmrOq/WH5lZNgZ5pUusBWdxzow2vSsn4Zff/F
Wd7iZS5KrSmOvzDsMuSeXij6XkvHQ0C01ta1BfUDD5kuYm4E0YyFuuobDy4FwFkE
JiTqUzzXi0SwN73/l9xf9QUTeC7ZqEDA28rea4r6DnXfDUWoUjwUs+qBXwqaJa5l
pQMYPxSKo+MBrvo0rbGl4Lrn0zKEyLnqGE020EIx8C7kHsEx+Yr3+mtZTKiuaqlP
JIJN1h1PFZLc+0PD605rKG5NH30CuE5g4cNdpf+BtFhx7E3ElAdbgXKYNbc4Eudv
nVjvvmqi8qRfHSDSHa3rSXsPC1frjZnR8pKPp+80DtDCoq4BYxwPSmX+tTsGByqL
8+n41Cu/pCGq6Jpw30A3Nq0JKwia4Lizd9m7fsnEhXi5exwygW9u8FuDaJKnAtiM
wqiIHBZad9ohSp/UuP3yrqCSG3UVzT9xhwqi7ciKs5aX7hfMuy0UHYmMQm4wiZtH
RI+VSfwIRxrJhqgAUx0iJZLDSOQ71/PKSMu1R32inIkcGFXMoVIj5KmGryz9UsT4
4sHd0IcobG7ru1VmAzhMbaAMjaHUtEWREiRWBGiJZh5eIHkttla1LS0vVbrFQk87
pc2vrZbe/KMboOcxTt8VS9BuBR3Yi9+6DzoQAnKMMRWx7lzp3EJUdn5yNXO6Lh+9
l5yJeIu7F16TgIS5QtVOfqh4E8mwAqxxasWDc1JczACyUYcIg820VajTZuQYRBoW
jsEG3aU8qdeRPwhi5UA/bfYyiWyKJ99Z5Ck7XkbTr38wytGoT0nhcJBEYUzw6c+M
1v2l7vgij4wQnWNYIBTSrHGNWEwJGIFrz2dUhIHqXZ5Nb9Fd8Vqz3oyNAM2ynpSF
kNcd4AGBWpgkuskRjGs8nipJ0fT39fGBhRLJq/5iSSUZdMwOcX3lXcEaqfB5FBUY
nLmIPZGGtGu7sib8otQgGHb6OT6Q0sfhGGosc+lMaOLzudN9z21z1Y4kjp/zG6oL
IRyDRkSjKS4IVs++VtS5A4A1m9lZ/0zbG4fF+uvvprI71aOCUZMQH0Uc//D0GtNO
7F/bg8UEnMlDOwJyTvdHqZgIL9FWYS8GS1vjJ8Q/Vxj6uXy3tS/jpet1m6NY9/H1
FqeC4iFaJCzZ/WvmLWNgo2T635yvYhE50wJO34wYN/YvudWpcmilNwqnoKXJ9Aim
tDYXfoEeDo5XU6zIRDXV0yROREHF+KBk+u0CTLYSTBoqsASyKdslCwVxtjJNluJ7
dSWFkDiqLYMC0iYuh3twmqiw4McE1EO9Y6WvofJlZdBqXgL+gQl5bXsG+JperU7E
8RD799/Q/D6TjU5zTDPvkYjdBHxPdSiYBqHpM1TEcq4QuB4rlzQyT8Qzv63rbyKr
l4eRdYx6QUfp8L8Z7CWQjpu2UqZuFEdvWerQzAhbe6QIj4yaS++QQ0rt9w8Tmtce
LVH5pWYiiTGLF2U95s+AghKJsCoJ5b5I0fy0hvWit0nvJtDC95rePtmvZooOySoB
H/EkEaKkgC5BeDui+5zP3dU6R4gpHbX8ygdrbwnfw/IMqhRpiVf3hzboXFpXPWwN
CrVxJKQ5Wrd1ughmoLhL/0tGu3coRnQfx9JRzIU+C1aRPoiWAPdrMnl3iLrNGytp
69wL3ntrMGIa7M0ng7uK6BSmR0MLstujaBjW/JYjlSeKVvKBEVLvzJSTRgwLrXnR
tGrKXaa1MWafj3TORMNvGqwuSLdOR3szjvNrj0a8b1rLV6Xs0dsiOgdiFvUaCV8o
tLJ2qjCj50hWUP3LEsigf0FTxX+o46wh1aHsqnDrFd8flUoohfkAZQ49oRAP1cLk
FAVcETc8+kLckmARrUWOc8rm7us2CBa83+t+Jf7omHTc5z5nPONvyo1sq2bsszt7
glmDEsftNx0zWjqPLIj0kFnrbzcHA0LLEKxuODsKiSJQy0Sf3ujgXsunjcNmCK7C
4ynsDFr2/A6fAtfqx31apxkbC5iPkxTixnWiP92/juszJSmTOO7v/Ery6o1PjaVy
5My5rjSsRHaYY0RBqKCb1A73PHNqI9oxlZHxdhImBcfsj6C1Mt/MJmeMjkPVYY7G
HzDsh/3/0q+MfyV28x0a83zkMZ39JRKiv0YipSZY2P6r9h6G8C9pEuIO6JLpFrdO
qErHFmNRuXDzTLUxow2etZ61j3UpVY9dO7/wRm0IJmC8FIjRuuxUUdtQq6AkUcL/
Wjn3LYzvT1iXiuSYIpSl6x3vjl96E/mO5zwgO/yGMXSB3uyWL5mI8NjBWkICBUvq
7DQy5rqqJKX4ztqOWPr9vgJcakLtOKHPWcOY4/hQZvJy8/kd9+cb4V/TIboTTbtb
+vJ3FBH72EwPAYXxCISkOTAgV+amx+7Mp2GHCDkUvCsxfzuUJ5GOJYj0r6XsHvwz
2Zk0PYg/S7qm+IMcIRcnKWN/e3l5RLEq9mi8ewo14KdyT6VAIQ+mLvS3/LHSsKP5
4xdpABbFEIcMnAxxOoXELPn6U3lLKl0mnzQJ8J3dDsb9qgVkYScWJlTp30Ai1Smm
FxCcvttP4jrsfZ+wH7lFw+KE6abU84XPw9NPM/tYNRsMlJgn0mHYBgPl+66FBxIV
Y7HqAt2dtQYfnbTPf9ybNbG2zurQ6yJCA368mTPmpxn24NDklDjdjcTAjNBw6hBP
XRzukZ3074iuo7ADmuKp+z2N8JRw1zdBvT1AEWegpFplOyyvyWIRW4opgdLOHhr5
tW+QodWq2s8HMn0oaUsoErBGzNVd8jyd9BGpZ8oauIn9q37xCqP7sjbci5jCUqwE
0efYhilmKp0d2DEHvgJZPpKDhqdGE7VwSue05lETwOAt8QTCWjERahh4wfzQ2ecO
cOlCXmnuBEBBodDP+uRYSG1ZLe+5wpyxkrLEnOOXWSfM4aqsxNnDInhRhKhGIcDZ
xNToxizGVhSwltwpkWBk1473aycbfBYXJwUHx51vXaRrXinLwYLnYdqpUU5Y8SxR
N1YR+1ErIph4/bmkre1caNJB+qnR+9m2L6mLyIYYZVcQgv3zeYFR8+EW8clLH4SN
2fisb1YIjvMmfWEWQL8mutT0mMx6Hatgzyqh75R8UsJZVuAUevA63L+S5w4hNlIW
NVJBk7L5o4ArUCa1Zr7vmkoMNHij1uATYn/aCfL3yIWA5hjgX9SIVDuIHldU5yj3
DDwkF7Bh8KeOqympqQgwPk+89ZrEPt/EIRYQHZZz+2XLhGjXYdynp+04lLVlqUkd
tE/tIGFzh4IhDdjpJOPd4QPTlFLSfIQxDmrGTdlxFKUGs7s/uAVPc95fGvr2y3pD
/NL61vtVGSQK4QJNY0PqX2BWCF3FUqVdRI28EiPRrwbyzkOEMxDgTa1o0g8pkyxT
XSF79LmPgkIkX6c84RJGFhZjUOLDFWvtmqfgMdI0zCUARuAEHSCW7TnnSszQOByx
6nE2VU46cjny063GfH6A4cpS6qQ+iZeUmqHmQa+LK/cuaS0KK7+wHtJ91j+CLPPl
sm8YUqJrq6ZTYlbwX3okR3lOw2tfU3gzG8TClPyEgsJt/MROWbmyF9cDhZcx34lh
HezyIWiR7/bNE6CCk2Lved6ADFGfUEfF3dA/hicrg2gl40iveis78LHoRhLfNqPc
W/DpkgwH1/JW31QEybpHNqBuKIaezoJksKEwcGFgQAwnNfHn4dn2JcAaQ3dULiU7
0KN6nDBpdzJSbUjhNrzrmic5powf+uArbVWtXkoutOsfH0Y/JifoJuQok9gPI09p
31lUqBAtdSdlidNHh4olK6C1oXtDvxnbQRekqAFeurT4G72aiww51shZViMfrIuo
NoRlFc6GO19uoJYqVcAwryXx3GpTWKt0AdXE9eMlg67MMBNYkR7SkSd5xsSym3Te
qXaIXco4Sp4pLbuaP8Dns6HAd787mDcgbACj2VcZmmiH/D8u9V0wnTeI2E4Lm3AY
5hA9aTE+AMs6arh/s8TxVKmahE8GQ5uCb3PiSTaQt+Yr5DVFoBqOqUD/DurHTC/q
qNKjMl0j3LBhCVfvkfVF1OfXLlN6BxoJVetAf2GA0j38tK5vAMBFpFXxPVMEPv2V
tjZruxUmKejkbGnn2CW7YAx7z0YcgrUGD4iPNZpaZ2DHgx4YvXOlblolzFgjNqWN
jMhcEtIrwS3KQgZhZN2SGWpL3VVr9N3e2ewsbvquNSd0L2RyyxaFl0MmRppWgp68
1yajTLthTB/Vhv12YhM+m2Wzl4w+HGhAfQFiwUpjz9siDS1L5tyAj6JV8Tkl4pFr
4oe3FoBs2yyGBmBs9zCvyW3x8p3OkZmvy5bihlwwtXt3SAZDnZ5Ohvx80SrCBnAF
V1vqzIaLdIxl5CpzlBq/po4HmuG7woMt8sFD6qVX0+krK3iT4Z3VSBvyuJBzzwdY
0oxf0Eh6MSQMuoUxn+L194vVVKfHeJal7K5kO+Tvl88Tjhkrh4vBBbCZg39t+3M8
+3hsEmVkGsgtldOmtqQNt5zlQFEKRUMt18CeXdyQFY17fzFbuay8XvaiROLbN1LI
vSoy79GhTUJvWTg6KyRSJyUQvf4w7DmoKhHZdJTdQtt/ZOY2DYrgbrNORhiNAKTX
7Woi09dGRuZK6uHgLkUVIUVgX5E860oiwDm0g0u6/XZfESSpEnDRAbfrm6i5iNBY
nin8pVGA33I0W9mox/yJF24SKu1R/cNsAUA6qA82QuHnrmT1uCGF4lIQO+lA55l6
l2HZAo+UFxcdOsCtGlaPVm7VguqPzyVaNQDqzKZbebtlhGbYFvh2cavOlDY5CAoG
UWFGhHCCFuvJrG60UBRMuS0u57hT/FT8QZNDDDnMFKSsSm6Rzjvm1g3T/Tp64JMr
hri+IjwOtN/b6IeK5XA9xzd4c0EQYdltnhzXYOsQAyAom+vCACAPRqrdzwSPjbvD
RC66lQXNKKcAlSgA+vYDklnwQT51cg8Nc0oSb74qXJFN84CxDrJdnmFoPxKZZHTH
QdtZFlBG3UhIT9cRbP/Ch9C9ml/J76NUI5UImAQ9CTdnwAm0lUUg9XWkS6UUUI7h
5pGfvDG/fU/TmJ8j2UgxtyI8pKogQRrEjwULxIc5Dh1/63h6lYqIm3DB5p0A/ls0
fE0cHz16U+ewuh5AnJHY9ftcJHolMWkwsRu/SXRwd3QKWAqWoFTy1oVmA31d/sX1
ed52KG8tuZg2SRU8misS5MXIcsIaTzu/ukdaXhtxsxNhkUc90Vf4NbKxuak+NwHU
2u2wJTmvaCUW4O9NvDTj3PPy7bWQDhCHstC10hJR5uQ8QcEvIgcaCoQRseRxPzM9
OtGNtU68xP39VrVCpVx7CxsdmVjXWNTAJo7naMIXyHBTixPQEU6rB+famtcvDnvD
I37z3/TDl15ulPrBTYk8jY0ANiy/vuWsB/OC+4CxVRVVIMLwnGhZvKQJBTTgp6hN
K7oLLIjkJszJkA+i4M1FjXZ/CbrALBh5URYeEVfNAgDtgAEyJors0ykj+9el09/1
Nq8RAilAPY5lSzVl+gRaJQWdwJzVSihgIiManDHtkWuQoRqdeg3dtLq/41IM82W6
93S50Z+PWDQ+uSbSBJmqntdOogI8UT0laLBn/xwmGvtb2UhoXXJrl2cTikUUOuNW
RSB8jjBSz6oKfY5eH8K3xyoHVoNoR9xmhJsRZ2/EmFZbnHRyYc7zc5lt8A8FRAmx
zZlW1WHSxYsPmgN/yeSsQipy8R5eAggbyt/Nl0MPwtvz4+ZDbR8pOy54khT8+cfk
lPbl5WDqfCA2vyyqF2FLJwdzczLkuuDA83g12Ha0h1Rz1/QFuAAO96ofGoVjUku4
DQrDxNxaTAagclE9frKAJXkJcIPYRfS0m6gSuhHZIXitL9JnbiqEHZiFpFxANBOA
yhRelPzKXFXE7cU8of0k1q4606vF6SSWrTwgPOjnQ6q+kAseUGwc0De16f7Ikq+7
cRt70NrQ4RLsex1zrESU9u9n0RSvzoWyNUA1KcICbQRV6nKNFsaOMXyjWKQM38vb
mm00jc6oCu9NbVsNFz18o5JC3bU5gLSt8BcC+brxM9ieWRI3OSjq9L2GwJyF6Pex
BdFOPeYQ+8kOahXw1SDu5AkmnKSzJcOWrLmCbkzwUlNTbwO8x3G6xtgMmTmlIWae
a1iU+AZ7oEuo9jbNklEwtxYeeK/hK1zG7ct0qMxYuBb2yvMrNejmebdsECEwIy8Y
k5YA8qLgloWRyG5TIAdqnM5YHF9bkFmIVbki0bI4Cb0IIDR/bPQJIMlq8FbQWe8z
CTlQefIzego3NRHkk0lPLPkwT6jaJ4VxpWMj5g94Lu7ptTZc1xm66ufU9HYwuoqF
vOf3Rub+BsT2qu/O3EPuukXbsa1UYZp3z63+97VGsptpMNxfW8OXyBjbQ9VZhtoC
7hacBYMw5iV0P9jrGIUMSOLiq/QhJvBpbgpv8ZlnnP0kj/zdtNzzv4YVzuB+usF4
LJPFciLmWZyp/JwomaPnuU1sHGtggiK8+/3C5cYJbL1tvJVdhG4FZufcTYCU+7J4
NSMydP/v5zDi1d/u5D7RMaEDF+yztPG7dUbMSSNLcNhghxIbx53fawlZw4ohyUTh
Rc/nDWXyMgftt48+oqGU1brrfhpHajAaxyBs5zJTueDbisXwiyck2Gh+JxCx4Qbp
rY7Q2nB0Slbaza/es7CnXZgK89j7ZyU15c2gOZHLe643RTIvNbRLkSgVpFf8nHS2
0gxEXXKT/5TDy6CXiId8uOxVN4B8/yPbiX4df9Ab4IxbIDFbizILalM2iXBhIPxO
FuWRYzbFwtGzP3X1iiFjbd7JLLhWfFXjIXpPlMPxyjHkFEpCigfbwUb/SA/byixJ
a17v/Wt+p/e2cD/LSgCGevPngrXy0GCnJEMP4KRpdqzOR633fb8av32PND8X6esb
cRI6wOlXt71uk0fZZJ5hDo+wfLB2mgZvEjx2xKIOih7Q/a/WXqStU7vzg0vp586O
rxCbQGdDLLhasG8nRRnq6/JJwV0itmzLD/b7bEz6Ik8Kc9DfhOh2bulfXM++Vaqe
MYcxvgjM+zlkRw2OI8WiUQQgXzW/pO00qQDDUHrfGD4o2q5HZMmjKejMGXFC6iPz
7SzQYqblEo5Sz14KGFFbzwHFaYNpJIBYbyvEGZZ0RgEVvdx3QliBl2Sa+dxrCkbG
4vwYHpL1Wxky0c7r6srTJMDKumzNyWMn3JJWjVpU7i5Mq55EfkR2AWWw5xODAoA1
lMhNowOCMeLFNzUuNGGMLhAtfAkYy9rXz4pYr02BMkWG61DMKQwVLGbg8nij/p+2
6K1UdZ45pS6hidbBigAk5QFzvysvOrfoGUuDa1EkqD9FBg6XXxjV015XZIDknhb8
c9hUeih93WJG8HuBqUV9cC6uCBt7nwNF351/o3OtBUm4dcgPiDz3mbSKi/UA1ahT
DsvGXLr1kawezoATR4sgu+K3Xd/CL1b21VScorJcLZSXaeQYHo6pJW3GoDSlo1rO
ipchNbkn5yyligx/z2VtFNKdNTKX18HbUqj1GBkfeLcP9T41AYUNdaILNU/hMkSs
G6ophIEHjcs13SEqJCle/S8mWBXry6PO2/6irnkDkqBy/pGmN3wp3KYzysHelvTM
1Fj3MQwDYw0slYQOW9Vwo4gX6D9G8FClVHiq5NaWJ5DsMNzlpKPx0/P4kzuHE3rM
M/i/eTciln+W1aRVItCzBbzhXHTXoiwGZn9JC9w7UubZLyYw2BHbJb68LF52kQan
0EBpfQI+f3j+mMnmYWkCHHvs90IkoHmYQfscteCWb8vEGSWDYU+ZHhHD/sZbTP4i
Zi1xP044h/r0qYXinygHtSjDGp14U1TjyShtvNBX+eyw5I26LXR+RFV2TN/U68e0
v6DVEFyEmAQENuIUNoh4gtbuYx8PlDxfKd+7WHXzcKe6nASkxXyPSmX+wE5GnZIr
9VrvLVj49WynjNCkSZvNsEHYCsoraoU4240hYflhVI4CZkV7h6vw7fw5zOUV4lvz
xO+GofWTLsG6qVI+9LZG9SQrnNGxYeLTi57KFkc9V8K4wPGswWwlYFf0t4Zjuo8D
5rx++oZy4aRsQKu+Q7Kc2rhd4jZWBZ4RZHnCYw00x06w39+PsbXWo7UkL63QyaZy
eiQapt8LgQ34P2XE12qUzHyq4dCGCeq3M91zCqL2HMviohR4zZ/HojzH342km6cU
NKAVwIto39Q0Vo+EA3pJlmv9iAZK1UasgqmPEjTO9SOu+Aoo4alZnKJp9v3tFRMO
JaUho/0OLNLPo0WTOU8x3SSHqKMTGkTNbt2ioa4DGsE05xVq5b+2Ln1W0rPXVM0y
BYqUM4qZ5w6hKKAZjV1pRAM7wTMrR7FN8TGYC2mLUvGeOqLN/4i7Lcg8+jLBDSfP
Z+07EFrIUD1L/dCSIzIUivxj1edbeGraDVMNjY8KXS1SxfdUDJZNBBAuwrVEmPIR
+EjogDI+QhOIZGoeU973zgmn9iU11hX/o24m3fPcyZyYW7DV0B6ztUCZuX/aIknW
CdQhawWKXyHaZ48FVwRbS4jnno6aA/ORexstU1QCD7OGXH4OBDgeigKfPthkOMZS
jl6m2HQu0dOI11K7VxkXV1dytOHxe7pGiorrJ0pZ47bezg8Bg+HuDQVg5hh0IFpB
FCq4hil8tkKrzsK+RUUxM8eh0DxKWDmIoUeAukYOwCGXwNCEi8Q1WnqmvsZVK4eu
boZA5ESEg7sQ0ROCO1qzPP6yLK5VlhsNfe+/jVGHoI/fIcxSQoLbb9J8GiwIGw6n
ZR+BE1pSix7TEHoS214fNwABrlpYjxGJ5TAIIsfpPqIhaNpN1ZZ+rDyavq2YIZLR
2l/QHXG1gnWkMBFwa4DHtEgbc6QYiNgtg8fHye9d06RjV6O3/Rewgl+Bxz3L29V8
zt+85fV/F0aIudP5FJyBn4GNzfGAEpQ7y6d+HcxEBPXAGA6kwJttKDS33qJl3hnw
CnkXLDlsf+n9QwkY++xPmFB2VCctdt/fOe59UP8uj2p9xg+oBambXMVwlH8jgYoO
HM38m1c4IwPD1jJUE95HRnt1p/3nu6uEiK1HKhRpQ1pA4NzAogPIMj+N4715mPeT
cNT9xoQiDSvPr3kfMfplgJoOo0djF9K3IYV0Z4FD64p9RN5Qw4RAZIHNX9hLJzaB
MKh+Dv+mzvEElPciLaBlv9EUCVXaRx6+XZenHo6yzrUQVG/rpcRzj+4X9nK5kKwy
JTKGXSGopTsD00r9c+91V6C+C4Rv5mp4OXqHAbm6kZLVHPDHnQzc/ANZtcDCykni
z3B6mJeXXiRILxw6rvIRAUDStth5/q7uKLUN9ug4eFmVJm8YoglNxCyTflGsbt3h
RscR9xAxXANPMM0qWp4xX1gErRx2pD75susEqgpbt9I8Nh+JSthzlt3PSMIXH98S
7x/mTEYG1V0iztVCtW7Sf9G9XxZhSFLX2mtfphfDb9kktRa+/iNhHCT2BGNrq9aU
ZqVWdajYa9tgoO1Hb5kO5cAKJMid1pBFkWXnjjLpfDYwPXPuCQXvTBPRY9hynDL5
P02xKbos5/MYHSzNoqKTTOeRtrSWhLTsyH0Ssg+HGbbB/xZwG8wnSVwTKQon6Jhm
YmzLSSSa/EGHcNFlixdaX2HrO7/nWJH5DtMEMzZeUkakhwtDnmYvPQIatn7P6AG/
NKYYeuwGDSqAB0+vtsU0rqbNUX5ZMzkNeSLXLLHcAWYp+BW6Q9xrCbq72AXODSVV
fNjIIPlliBv0DneeWeP6ZjamlzOWcYemH15rPcn3F5a28/VHTkBJzhLQ8vhdXVi3
1fq4ZwN9XtakZ+LJHW4GPq8D1IgAu5ddXAiT6VZ6OL+A7hNAL4TNYD4Aav7Rpr6H
ZHKvOGxOBXsSCNEYhmprTFY5BNmtuptYOOI8S+sqFJJwYKCVtfCSY4I49RQ1dVz1
H8RRpmciLNpwDb5BLq7kzTDWOwiEoS6mycmSxZ3Lr5kO9xr+chMfrX9DF6S2aB0D
tY55WSWiP1rcJXo3NaCLYTIvlP9uLY/QZJxYGAiWwWzYsmemSHvykYc0m4xHCWxN
g7yMy96TUlLD309al+oVmSBwu6kVhxq2k233AessiQwfWZt1y1YVpRS6uam3MphF
FPoVizep9uropBpTMBMR63eEvT5OhfXBoRTkxmekos7FW+5vfocpX0i3MfD8FFaQ
jHnhs2Gf9ticrZXcgav0z4zOHousUJmrAOj1LKi9Q4L5sT9nbj2StC5DermtuALv
itX/0SwR1KDUiZy606BcT9mNPn7OBecqkxukMMmzpuzAQV6SSB218Fa2HIaNUd2p
Q6dBPSD3Koa64R35Zel8HywKwYueL6/KMnx5wcMFgZrxYoF7hxdhsLAK8dJWuvAh
73bEU4uAud9hkVJQokoCxbYRN8nE7/vctJ1SG4euyTTn6CbXhP+HsYkslKgtuDrT
x7NEL6I+viEaICMxgFwPJ5/n8uuUr9pVlTWtLWwEHYNiOwiggW4NROI9SeFxxuJ6
1KNEKegBXxUCJ9rtGRDm5wY+WH+x8qLQlL5OuOcdBe+8ys4PmJGHkDqA+Lg4p4sn
Ya4hOCP8kzP60khLGs7172Vu/q3CF/dWE0Na8x/UecKet0FJOUuuP9iBlSXdh4wU
D9HpoLQ5wSG5wjI1UA/GsvGYzWPaxCKH4fCHrO/Zu5EuOcnwv932hX5H3Lb+qUi+
pMf53Y7bRBuCQGqUE3g3oi4h0eBghGOb8TLZHSBiMv5a5O6li9MeAXcqmyMm9vVq
3m474nGeZoDeAWHU7DoVMUaZumCxM/yWxjDsEgXmszwYZzY9+7Engh3YujNpnPWn
KqdjifsOUxj885eFnXI5dxOS1jOI7pWo9NTX3SJi644GCGWsXDrHTVYvzMhqmjn8
n94jLRV9pQHsQMsfpW/nklS54rYBFRitcqbx8RrZpQmPjS0/P/Uazc+HWmRJlhDA
jS70gWRPgHM7yLK+5whyvdmvEsbvhUslWc29siy2uxrm+UbOobIljmtaoC7pmNdP
XLMC9SdXAvJ3oWklIO/w8Rre94ksz/wbepPz/v9xFqfgvuzuoZdoiN2CmX4qr8w+
l317/WMprTBbFp/l6omYwfC5TzzhOZQaK5TmtXS89ghmiLPaafP07w1CUiXt5LYb
OE7bQ9WMftQSONQQh6/7yp4+63jbkm6y2l/z7cAAPjbF9+6CTTsxWzzYrdCybSZR
i3H/vYy+M8DmUYMQvx/uIKuUTpdFWLGdN93a37ZHD538hT9klUiQ2QxnkZ4tg2nV
Gumv8sUJdJoElZgPvYbnixsIYpuwG0rR17c+flOgPckNfAt7XXlTAd4dAKjz2oTf
98bUVQ+/BugiR6+rrVuGsp/viRH3PGfjVx44uHeTxqJuS0Zs7dZsfo+NVleW0tIq
+hrhdF2j9v2wKNUVoXKnTNaHERYsMTWi6sOI6VGV07JHf+vMNXqqFoHJ0hKEAP0y
pvdVEM9BCNI+RWAkloxiXYIEVM0LKNQ2kejSBlT/08sJQZJAeXPy515mXC1QLg+U
15ONUWLamJK+A04qPo+h1fSCiSMuWvv4PcXmVlaDYItDwHNbwOYfAIbe/lT6R2b/
1D6p+VFsz+0vvEBVdtrYu5fIoebwbUmNe8NJBJjAdhqub/RY921IXGN4mAifGDLN
F2QLcvfxN1j4v2LghQsToT1uyIiAfDgjbrs1RK1bv/20jMGmtqJ9mvH/AkzQsPN3
R6A8WQFVkmL1I5SMA83vVPRJu0izkMTbaFAErqwVpoNbgL066f7MpYR8gjWkvaoi
QB6uzVMHPUHg24UsgoWzJHm2f8G+eHma4SXmPuoZbjVTIMRgP+qAEi1Pe2Bx7l+b
FdDxvj7nEDn9iTQ7PE5JO2wA1tgIh6JiHv0YwB9A/OCVO0ZZMYRHfzFvfrvrvaLm
qI3SVlp9Vdhh+T6NFZYJgZhHEsyK6bn73BBOeQ+CXK6b2jz6pA2yFxLTMWzIEaBz
QWBLZak/i1udmyDrmLxhl5+RG5kQv8gizkfpjyQQa476zldvMPmOkiNrv3LBKUnV
P0hs5NWtM5h1khDBCjg953RCNC58ox5TbZ8VHjDOJm58dK5lWIg518C8s7Y0qlC7
hMT+G7fcwHMtMYK5jqjGRHzeumtovCQKpIIlo9s3yLkUSkW4vQrn+/9JXPWzrf8T
FEJPjZdq/HkzofcLsIXguXei/JfoN7PR89U6eBOG6a5FSCjXLhsazfOgCsQunq1U
dMOBMNvVexLi7Fl+95j/ObQUsS9o6JEGyTJ/Q0I2DXivzo4X8bFRQlZJrRXA/Umu
O/TagbCDYOcuyTVHxbcTIvqqYYtUrkZ3itoAhzz9bqlx+Dof3kLevQz46CLenc8K
HXCjpadN3RB1phRDI5ftf/MDvUfEjSoHTlcfY71WUjU9j7F+jnQLvxrEv9/78rlx
jfXrm+2PAzqzo5pNebJsPsixyBeF/Ejwk2iKbPno3WvTHoOb61URwQq+OVjT6zP+
2znSdHV3LxHd83hUL0bGS01ekJ1o7umUiumRUaojX0Uo0a6F6bQfCI234BeggPXG
ffs77+IFea5VLppmz2f0IKmS7fsIEiYzdcFu81JbvZJpTHY+Qd5AuV2f1BWA4m6z
Mi8+U6WDaPS9Idw/0DqbwHIFj+VLw4OWR5l15fanD+xBawoy8K2UjLCHcFPI01tB
/ameg8mirmHo/MoZiF47UiP6h1O8OAI0c69RRtdWrO7OHjMF46NSiB8HraY33LM5
ROHjPbNJubMhGT3I6b0bgQqnRm3CY/F+6SyYoY6YvAG6wAsmi3k867vsvzAXpXpE
J32NXfzgOsK4eHULYWIAmbCnSkdWTq8HzZJQOqToHVPB32G7xyO6vBKGobXAqey8
XkTQdxe3N5BhwTmu9/2BMQcYEhXQ1kl9CXu3UbHaLSGYiqCxrudJ/hwEARKVt5oo
HNdTSQwwIAhUAtCVp9CxfDX+Gk8+LShy9SSw8RdZ4FXkhOpyr4LpnYx8hCpVb2Jl
VQzeO5bIRuK6Wt4aUkXcngKCjFd6RUCMS0wD6B8dSML2fofsoYVld9nf2q0gp6lS
DLcTBsPMelZr6n6B80bTezdkt1PGavoyIDLA1NeXdWKUpMaDTv5s5YAVOc2gfXNR
c0ypnIfew3ZbXSA23k39TTsWReSO2X++LjlzV+euuk5G1lGMAF3LovFY18LAUeKk
johpzWCcFOTGthR71W8JtUXFs8hwv1xEzEhigZs5TG65KpzASorr7EnJ5MDwPo5b
VFZNaDeNA9o5zGrmx5/B8/NgG+hUQSH1R/0uq/zXFvjo4hYZxh1ZqpJ8NkFDFXEC
WEh+T3/oSrC1GoZJlxjZa4Wjb4Tm59SNpB/F8djCYnmZGGt4FEu9Jly2dKQMmAqe
+Gwbc+dhDA196Erc9BbmFXFxIsbsNNAZUAKTqP7C3aetvZoqy3t2tQjq9Xwu1+Q3
QKOlEK3YWAp+1GZpnkjZgaZi4zYVH/OztNV3x0Gy8Zq63Y085nua9pogwPZZ7Ya2
BoZCy7a/8OQg4p47thvKLTrFOGd/Z/OPbeKT9cnjjGR7nizCAYSEGrXf7V5D5wDr
xCn1C2RBjOk8dVOZqqPZSuSMyj6qVNzgoZ/LNViVolTXnNd3XYMfIg7y37yxWBHv
XLoc1r8yqUHLVI/woH99eOzsPGHQAwrNnifsr1X7iWqi8MCwfzMeCRvAbS/rJ1Fp
GRH872kFWZ0CPaBMteeBWzziQkymjB/vO3Q0cN1v57gRpB18hP9cZzHdiqKVsKot
9c9syKFqM5V/H0a802xkR+SujdDTJLSw/MRJxDlrgJa5RApJs0e2rjdKwc8BU2d1
+uWRe5ZUQNyPU6mXm80nJ2YUTdnjRoIFwyMm8PYHJJ/bI6hy7n6Uy5denex6UxlM
S6wf1QTcU7k+/U9CsfCozZd2HG9rylcxbI3rF1N7/5/MyXLrwoF0XZKpBhitIJBJ
Sbkhq7AQx3sxI9qp8DaEZlQ6AnTF8Pret/sp8zWFSeHKZ3FV2LgVQSzrIV5dvjhD
DDb4mS/umm0FzWq2otZUKcoGOyrOL0A7gxUkWxr5/bcN4bBbUy9PHvezqKn7H8wU
tqTfHzIPQbwgwJwWg9MXxFNs0+nIxvDJuGjhuSabNm6RzE2FHbAhRUYjA5KpE5ii
GJvj+8KHuE/riC40KcsFJfWiTKsvgUvos39ql+c3VSOEEHEYGMTCFqr1NyKVzEJD
upHzwyU4KywtqOGRVj1kcfWihCPhb1HP9AHZ4JjLps25SqW3QkRDjp2fhQHcTXz2
VhNFgzAb9E+l/1fynnu2uNiCwqOfc3qDdkTVhwhc80FTg24HORR9fOXz69udtq9V
BhCR8j0u5YksRu2hXqwBVhlaJip7hlFT1qSaNe+Z0/8iUQDj0w0+jMVtW1fFzFEO
Q16ncYRrjjWsr0j/sWqW1iNnTvnK1Gl3xy737PhC/WoMtbBtjvpm8gKsyzZGu4Wo
/lMMaE5iWgqKGh4siUPIOxS7CBXoA37Uq0PQeuKgsR4XkLaA8eZ4URiI+culqrxD
BUOXjFVv38OSezs+yaHJ2WJmIlbGQggPDkGtCzEPwMnzFqbkXpTzG/gJl45WB2nJ
k1uNr440+LSh6LuyMdqgG2ue9xSkBHtzqK+vkVhgQpgsizgVjYe6maZe5d93YqLa
UH3WpHblsgwnD89rIRJEkvnPHvulzat3tAq90KBmiRVA7znMjmgGrLQ9i6x0Ho8m
WLzsUaAKmSAM9vk2Pj2DX/UkoZBW5LY6TM3jZO1itkyp0nLyNfUzvb3FAAWCAg4s
2oX5/YGHCHxzi7oQ0M2ij83ZuvySbdJMZSDljwLUC5411wQh0/m4Y0DClkPecSI+
ozAqLbAf4/5OtdzqnqSRLEM+ck8nxoYbeyodqbf/bDC7Nhiarraqho9MW1NEN/0u
i4nWz7tvMWfRchE6S4fGBAyT3ASvv2RznrtcQ4p4H95c5Tbv3NG9gBw6gEDliwji
igi6eKO6bo+oWVYy4Hx7BsU9c93qW0HSoudSPoKAMwQ3yxAdP7kVK+qvEbseBkml
Jxix+nv/v9kehmIWcPb2Gigvq5WIVxbQzytM+ULECaxKDpLS6F1TFVHuQSu42+Fv
gds63wkowUunQdtmOUXQtHBc59rXv2ny0YWaf7u9ytx4cNOn4hcLd8lPqakR3z5/
qCSzeXMANpbTEQvekdTYu/eCgRyinRUjysAlqj2zV3s2TqIVRE9VMc5T7PbwqoxU
JDGBmhTxeJJ7IOv8Mg9DfbZJpqWYK5lFmy25CiwNpWfsUnoPQAv6IWLMIRrOOJzs
hsgtV0LNVKNjFOHyHPwDwBHBGVLftSWxmbHQBL0nK6CyiPG6XSZkYU4Ypbpiqc5z
JKzRv4F/17XWOgAz1MJHrdL3UFM5NNWCa41ZIWnUq/vNElIZ1UJsTHb58iPK0GkA
Jy1I9MVAtBUU+c7U09LJgObNnjfN2s6mgLgabMYGRmo4OpxIHhdzlzPW6UahT0f6
AO7pHSR71z7qG6ZAWMqFB+gRuyP3bzu0oY7mFI89xgxbg7wE811AAHXd5jtdBkRb
gFcztjbX1tectODAnZnHTp4tuQL2PDNL6sWqxebCVd+0/RZ0QSk9RTFzOuioEP0k
2VBq8Qs2mFohkGrNkaauZmLPXxWqDlDZENi/YG5XxRWo08CHQ4XZBO4muslGmhIO
oCPXlRNXY6z2RplMpzj5kgrVSOcYDTUyGvl2AsQL6Ft1yxK2Mjwr3xOD1stuSkc8
z41LHrLzrly1xRegPp1l5NCSxgfjr2Sh8Jx2d33PpPrYcjk1jbCeXG4iyqxsU2O/
J2HazemDkKNSCpVM8KVeNBo37ddv2cBter0waNTiTqpIa+xqvTt5aQeNAZtYn8gS
XM7+KYxdMkQiIcHMAsHpsiu++ZlHXU7NCOcQGW3rp04ZGw05PiL2MGOxiisKSF/D
E/VhikaW9Q7umEs3+Nv2V7t6A32WgDLA/NNA+4jzyKj/boHErXS60/GA8ApAHozy
ojnn4DzXANDxdpomMQYHSN0S3W1tFSx83ytoiWB1mcWiOlqzk86k4wcxtlszb56f
m83SPS4hpa5jekKDQeafFRGZT7KZqH8wnP4Tdh6+pcju9tu9OxHydxOAgs6Qwopl
fvGP9WsfBy0MYalT1njkevqZG7w4U+h0J3VPBQjbMjBiAG65JiK/oEwUZ/a/AvNf
NQem/9xNo/Ce4uxyIDdcVI34CKTSCoRgxo7hF5tFQixBEDGK3WO15cBvJyVtnN0o
AIDjF7ZF837fdcnKDDM+8qVQVUdq6dbFW3TR8XruvPLlUtg1eUBi6i5JjrtxWDFU
uULBML+QHeUFkJmcXVaz7BLk9Qpw8VkPzDxKua/IIx+0OMxi787e2BxBL3oA439h
h7LDqMrJC7q0WemypF4UqKrO7TUWzsPxGA0Suckjn9uZSuiUQBhz/7ihd8LxkTu1
98aqer0nlbRSCa0uLnJhs1cTZ4X8DjSorYPfv09R2ciytqQOB1suybOMZ0HoakCd
VOYEdZXTMYTbuyT6RS+y1xDrCPFvSxG96td6EFEiBjlZgTiScga7L5m2t2t5h5iU
V0J26C8+tjcgzBkhtdNrT7mvN1SnL1DhqaStlmQnnhhSXF2yva5+hZRaCvUPdOvs
hSqp7uUDA+Ls6AuvG3unOFyA8imdUToZ9ovImmidZwbmBwvAWrDbKgf/ym+VdVrI
i3a4QtUv+woyNudn7nHsOcU7F/ViQibBML3YLXqABLIen/a7nLjbfRboUr5wxhQv
hEAmYUPhKpSvRzEFpm67/8VGtTNuRl4aZ7k9IIDmzEnEX8bwUgL2TJOvKJ0d7WIP
Z45Kt5KFzk4EkeccgscdBLKa3A8OVSEiUUyn3PN+G6mVjWYQYziFRd/wMUe47qyq
uyHLkM8lFb4VTgrSxklb4TifPgPd2PwmSeeT9rjnhYKPECieiNQaPMYwKvZT4c+a
zkroHrGV+ARUjCJuxAu+Z/HL0np346UBQ2QIKsi15Yk3+wd1PyWggs5jreKXFCV9
MMPKlYMZdITCWRDFnK37gCCaLDjS0bnFHehhKq9gn/W9/sFP++jP7s2abPmpbid7
hc7t9frDKaRUjtIn51ESC1W96xkb/7X5XeKJY7TlkDESQxMAM6RHB9JBiXEZGk6U
IGk4e1ndKc3DM8PcRI+jlKjfGkl+10sUP1/8z74SLfqXb0L7Vk4Rdl/PAJ8VV+Og
pEph4jH/T3NHXIROQUA1Uy/tJZdJsvvgmhrt7TjkkrYXlyS1BRZY8b0Ee6wF5hdz
zpm3dzvn8CYgLnG+K/KcThTQttHtYplCVClGM34h6CVdkVLVkUVRNMaMGGSpRKcE
BSxtklWsXmVF7+ALtIPxxvnknB62RDOFaSpgP8w+Z1r3bBI9E5bDdx0sUmMnKYzu
gZYJj8dH2jPQzvGbBLo8RegJxVStwyrjTzmTnqmY9XFCPTYmITF1rnTsoHCL92Vx
eHgm4FNWS033Z42akK+fXVrmPGrw1kdMId6Sl43iOMAiGrMt48kLib2e4wMFw0Fq
dBtFscCjT6dwgRKVyDWqqtSuAPS71+hFzxWIocYzJuuAyN2AaTPCqqj6cZW0JeDI
W4WprW9HqC27veNuzSobUid3QfPBLWlkSd+7gGrvVSTuTJf2wIVCeAYfuikW1Thq
MITpoIWZmBxipNIDhrEONDCho1zcFpeZayA4sugR341AWPZ9pT4D17GM0SJYk2nU
3DdNscT3RTZcq8maKJoM1eASAxwocfROLd9tphHw7Hl4Hg4wzer+U1AgMbmqhqFQ
TPQYf4JhrMgPj46rRkk4Q+6Lk5Lyc6F8Ax1eXDZC+l91NpbkXCZmxeOuwjruKsx9
9Ic3biDyfsPPDai1QmaSKoSw/oMSlcrXIsduvUzYn0wDG/lNyr6jH9ZJg2vd5pVf
NL34OA8+9Wl3MR3Bsw3aobt06Bn48jdFG4M3BMp3s3xC9F+qCeSLE+6J9n2dSEzu
nt1ViQbQpVFP8c1G7VdFPwcnDWhuuVyu84MqkTACWSq7vWcNeL5HhL84xmT4iR6P
+kc/3pO01zGdcr5PCk0+d4nqU9ccipQqV/lOMrAEpKzm7x45wEK8WmKr4HlcMHEo
Z04lv+NhbptfOCfP+1GETbf0myHC5YWukbdo7HYf9uTnda6g8kFraqN1LueGet8j
M3mt29XuZ5wsKJ4MX6Kk3S9AVlJvqOuzA56UnyoNvQO+lhkfoRU0o1cYC/DN74gZ
mfFa6TnDY5PhI8AWdWFkJ/g3b1z021ZgZmt2qDDtz9tTLfvVLxBeHUXelHI/un0T
F+v52v0SzjPDagtMjvjnPFVYv0TOQ4qaMT1udK8ZzN08fmlIqbJczRraVHSzm2p+
qIZWNVqFJ2CDZHl6uHzHHLutSsK54nrkQW2Rv2wjF37PmC1dQbF/Y1KfSQdmfiz8
7e6MYz8hH8QLvaUDG5x5hb0p/k09/wN8Oo0Am75Hbk10n/3/yNMbpiw5PgG58oCI
m39BY/Acjpio4VLAburO9X2zLEpK+mUUwybfOC4wEzY5Zr7l+6iGBTZfYoZXHzYW
CEQdQojic4eJH0dUnWdo7Jyl8GLwBxjfuJg4fhyDTbGBY6Iio9eJArzvm95rviua
/UD58FkDdFKiCOMndCXjgcI8wsUxFk7c4Aylf8IxCzL7a90EwHRrOsgbXfgVdS4Y
chLZ+KPMxj4bB9JWF3cx9bKV8HJ/pOVp+B7JPabqt2XT66lTDJ7UR8mWKBhMmInK
COnDg0ohL7MmYQd16bhaQdbNj53HKQurjEKVClZKjonAJLxVUUZsVsiy1oYR1xi1
D4Qtqab6QGkdYMV1GJLhRtsVkKW3oSBKq8r4T4UGHApKZFQGW7ThfAR92XRj0QrB
ewNqfmGdPtE54bcxC7W7xUTRwK8b5/g2y43UoyiZaDHEgolzFeuWoFfMcMT9eNOq
Q34sWonRCmjQJNr7yf1l64W9q6LMZXrHJ7Tj6fFFUdcs5sf4Nb74TM4QkVjBgGxZ
qD8KLY3XMVBK6ph3v022JCVlDs7wXhhBx47SjfzM1A07ETv1AptpWdnT9PolSOna
d4sXzBKcawVq88SkWYTZYaMgOPtttM47w/hXk/6mpCBvDVsIDM6/O4kMPVnJKiT4
SDcvyMFVNY8by9x9p2ZrU/vfm5E73a5Z7W/8FbGVvCB7BB4o5FX20pKugiL60Twr
MCx+TaPKOOQul6+SlSWLwEDbdDrPqRjg2V+LTcMUB4rljf67J+lXxsBXn57Jp/nv
DEuQXPK8hNf2h3mGEiNRglnU/QZi0Uzl8LFIRSixw/F8S/C1/3hmeMaZNT6vVC7b
Rn/V7lympkaNZysb5Sw08y6gMI5heX+1K/FTU3/kLhTn9f69kS6w/2PBMQp01pDh
stIfx8QuXZRapgGb9/WKD8JTt40up4QDeGmliKIYJV8Mub5o9ILgu7wpGWF0+/ED
HCatz7mwCMJPZVAScnVk7ASdoclQxj81jcd9/B4cKTPXPqKZ7PYK5923q5rJxVM4
UlhKLOeZH48qdvrg0MHhOgYAtwYN3OTFbSOowBeps8YVVPfwnf7w9hQrkmXzkTpZ
uChabG+oUStu0b7PWFSzAl0tgeybIlDwEpTsqxKfeggD33usAS7M8CXipyNsnDDw
x/reRu1n7K5mMDmyrnc5s7G5b8EQ56JLQywKKFfQRKaAsWDMilIcxAdqhViUWO2N
NZpL6uah+74bUg3G6e8vHLd7A2GmgT9zPVzE6V5O/Br2TVvjl5rvCqBuHkJVkexg
nG4qw0/lHWFvP2Ym4/1XZ25hthuWTjHNGMFAdBzdRpu1X0odaRdrrKNcO8ePScen
uG9Qkt4X7Da6P7i+hOaWzhdTaCstiY0rXDS2BDHE6C1QeHENHEY1AS1MIuXEwcrT
q//BswG7eUkDYK+XXjKkvD3TS0wQfeJjgU6BVinG+WY7aACHzrcwhoNiL4W0Jkt2
MOeYQICTBQKjXZnPan/fBbTOlD0YtKItwGIhhvzcr+gHLIDuMn+D9L4y6wUFADXw
89YXWGexKfdwH+7zDiWUrGmHMFSqH8d5376DLfbia4YWwqn3qspCGOwKiDWkqvKU
RD+mO9ZAPd0f6/xjOpvpCzu2kP2diwL2d4X6EcJP81BNWVQ3v+GP80nLFN5Nb8oA
ExKAp6ekYh1tkVOdszif+ycTpUE/gKq0+K5B/R5Teucl1zTbCFLEx3CtkCC+EnFY
ZZivdkkeIWNdo9tTAaChT7U8+aXO/JlKHhUkAhfnUmMmj6NF+u4l/q6K+u1zN8aN
l+wBXgBtk/CxinfT4+Zb/U5TxxhzjJCpX2nywNPQF45aZJXOvv3X4FyKElO3QDiy
MCPg0DFyFON1qu61m7O9+M/fl6xe8BWTGlcz2NRiC+e42KiL/Gwt8Ae5D0Zq6j2O
2KPUZwww+UnaVAilUyg44V2MkEelzgmsBUV3eViCTWsNe6dYYIqFvOdA2S+DXIjw
hurAAtcGMJZXhi14uGdXD2ZWS/Sz3Fg+TFjLh7ERGMEwN7gR5H70QvsZRSldnyR8
O2WZ5ylGpK8tTXsRlP2gk/zMugWIFJz3hqg4pl8JYp117MRhS9RRR1IutCJcEtBK
ewVbCGTUOqF5vVF7XY8fH4JfAVlDAPlE7Bv1Ptp+VGjS6sSEHlLkmK7A9j4avSE5
9u/fvQqYc7N0bkqyBx4eZUK23vTFWkDxkJYHTlKDqo6j88qJ8YbSnyFrd8xDs67h
vqdRVyTvXkmKjZvwh/wcV24/pwycNvWs2CrWC/5KlZ7bv1omx9Yfc/Lj66afxMsW
ax9o7mwUqMBJ/tA9Gb0tbebUGxyK+4BUNQ2FOB1EHMYFW9UH0CjXjxH3cYHfBEuT
para57EM93ivR69lvOh9sfGPlAe3coGKTRN87AGztCaI2PTBsJ5PpVMxv4wobWD6
AsjmZestvgqyTrdHECLfdRuw4mrDTnODfXuuxMP6XZFCKtGX/Bh6wabDgnNvKqth
m9L3XcezU2GezbyESsMG534pJ2pB/uKsZMC1md8fnDgNvRhdDyqy18NSw2hIx9WJ
HwX8ivp9DUaI6Wy2LuebZ9UAfU1PGQEE42HJ9SbhyeIZwvXbuhh9bASHxoL1lUPL
2CyBnm845e2cIm5J43ZTGoEwU70GFN5ZBVt8l3e9dxYiMsBML9Tnh+/1TndkO8cL
WM60CbFCmDg6n3b56sa9uwgQOYd53dQxvyIt9SeD9TJ7gy/AiAXNqWWvGvToNPp+
LTmrrdteXoc43G0c6++C29uQjt9fp/3XCND+2t1fGuTv/hjlQLsbyVqaIgeaWTzW
fj/ulhVjkHX9muPKQY2awNDCAhp7B+yH8+i+9FnM/k3Y+MBZcZElkG3J5Mm/fJfu
DZ2orUwrYhUg2Ky+4DGWSNtjTomG9Lwk2YW3putwCH5tZ9tVfkhZkwC7RFoHW8pg
YV5JKIJEbLFNXgQRHxrlC5VnhlhOyXNr8K7HkPojj2rKFJOzurwEvlD4p2o9Z/xJ
eF5lKtDNXnYVuF5btD8cpzEIyGdtDICzVeyODFhkoMOBZ3zs2I0j1U86fGi1Uh7O
KUyb7zSxzArsMPWe5UcALDu7OISrNMc0Gujte2NK6UEviWWkskLzXNad7YigKIN2
zQnGZ9X3mHdHLITdenw5LivrXv6/VeL9aY3PN0YiUK9qr14HxZKMAErH3OT43QE+
XcFa6uqNQRLvlJL4EeulG8NDpm8XN0gdF0BMiLtcmeWbhHnLFAlZtunuqLIZgn/Q
cd7yAqvR4iZB/D0vL7Y1VicwUEilKZ1/A8v4butJqk8EJvovkkJIcurK7myIJ2LT
ysdn0r8AD7cWHs3Bki/GKsTabUE8WlTts4mrlel7MVlLMHJpSKqhiV5EHffw9sv5
bkJX14zlnjAX3JIyxQ8/t/00r5sJBaU9DYF9mieJho2Eq7GgZftbgqq17+fyO5Uw
Ql62rtxbfgdp4BQDUVuaXqwpjfOaj2Mfotot5Vk4EshUhahM+ozo/DhH7/93am0k
ZoCLUTMxJwIXe9FwuzTWjp+jvfWx7zUyk3mj4gpZE99SpUbowiD2yhcrR3w0okSk
Il+9MeL0iuzvlABc976I+qn5aX989jx0Ge87mNCvelOuSF/fDt1uiBXD2UVwrLzW
VkkCqJ6NqRxohTzKh1D7el/G5jy101w20bf2r0YflcZOfOPR5ssRdXadY/z+Ixuw
KeIFPdH+CyWsJa5ad9jWrBiMQ+FZ1U4Hb+79Yt/Tl5gTQIt6FbR+uWbG+lff74CG
Itqa7RdSkyyjBpTJjgx8/jxHOWkRV0qhv61s1vAiNABPuVCCaAn5JH4EVVUVQ+fU
J9ZcZx/QZZ0yMHMnK99ZSd4m0G70Y+z4Ups4xiqMruB0WgJaXrMLI9W3asO09wat
MY077AVDhGFWXGalQe9R0ujdLE7m42MKJwxFgItVS7sX3SkxUnA2Z87gwQNmBVC5
tTJWQ+ZjP/qzU4pYW74NWqC8ffArpRjMEmcv9e4RoI7EezLAFeF/C2weiXaAYHLm
vg7o0NHFRbgIuCX22q4+ISFa7e3KQqk+wQVvuGbbrL3YLhFgFelobqXoOimAK8kQ
NXCB/0UT4LHEDgrbkAwwQnmhBHkvwuCYr8I/iTe5gzaYgtXhN3YFrOe97Bjng+f4
udfB9heCpcdObFhkrmsoj/ZWCVj511LY+UT8NeL5/dvopR0hSgqOpDh4OLp3NTxk
/Te8rua3lFad3F6VuySHHndugQy/IkSXYUqUzmxDqjEGdtU3I/JilPsEPY0x+2WL
a9NZxuESQk8cmu+5ZiHGoqKSFjLVmM69584ZdjtOw1UTd3apThSD4eZvPV4CIkrE
jRqyQ+BvqfdbH1jLgBGUKW7ZPafnvPif0ppxQ+xBduViLGOzqec/Y4Ed+HbWx8yc
k1IZ48YOov1TKRWMnNBQfrmkO473NECc2LqTj76avifuiR5sBd/ffzHlMLROVwnd
6kAxHkKAFO6W7ZkHCvenXGi8kWeQmIhNepgmyjYvfC7neGxmKmTZLsVos2AXuK4U
xK0zV3xeFGJ3EHO+zNvno6NIlVFBl27I5W/yLjLYTs/6sHniD+ib0NpsIH5sgzAe
6CHFLXWaUZ17CQY4/g+xA6Cf0MPFCGy0euq+YftJUAom7gvJvMiK+xspM3lKP+6h
GVtaUh/z98LDvyzoy0V2E1f8cqb+O5/Bo69mTCOxqWE8AkcUJiwOvH8m/O75WnGk
6UH+tCiHbJF+x+nhVgHX31nda8o1pstK9T98reaPB5WMyS/0I+XZ3yvBhK7CJyzC
5Q/jPFOzhE3xh2WXeHPeKQRdtxI2//IWjmvj/S2OIhgJbQNSknJ/nVbZF+DS5T7+
dUO+KLih8g++Tzb6sHlmdO8ika90aBeCWEEjoic0Rz2yF72sHcDuSZmNwMqjXwgh
jnpeKg4BGEACDOz0u+WlufNQz/Cmf+Ui8T4nA+G2DyU7nXb5sll6BK+u/00XXyDK
Zg0ahft+WZZHNKI2uJTWF8su0Tab0dzNOfPXFPBYpWg0nXGaJkF0CgUj3qZ5TSNQ
2VRdPSnQAMVrUIDBAQI0se5GkDYAV5albB6kz3o5hn7pttdvI59aNwZmnkAqvyTk
ZGdmeQn4atDjzRu9JpbZImmSlaAHpSkJ3hJm0UkZocK8lBlOINSEsUrNnf80sKSw
8dz/XUip1OoPbwVeMa8YPQN1/CTwcOsB8StWAWX2gqoRGUkbh7wLmUAGQVg8gNeP
t6FGEBeBEOsLcw58nIVAxCMbJ7aL2TcvVEcHurcfDmmj7In4V0R2tgTPvaKhMAHy
Z+MRLoBevUrii1Zn7ZK3VdycZH2glmqFARnDmMu9YizI1q4ldXHHVY48bi0P+sVo
s7utNTGQImexBc5Dp/nOczWBF1WALGvmtC1b/8rNyepSultTbS/c81joBlpTwSqn
oyF/wQQ7c9ueYGcjDYdLftX2THY3dcDweL8dBNx9K4RPDtR+wvbCl/pmYs6dJXiZ
yA3/gKrNP7UO4RBKkSBjeOksy89f8/ArpP9A1JL4u3ii9mnQn6zufzjHK5TRkW/X
ClJh2JZf9tG2gf6M6n14iVHr+kxX0EFxEoNAgZiZrEiM5cXQhf1hlYcroF+fbNjJ
imdjFkOIlgdH4V4yoAbcUflwjSU3viWmRdBT0hK+LywhB8sUiFFO3p66NK17E1km
CXwgo8IWtJq9pVyeAhb/GTKUFPxRYjdeDNJF7lGlYShGM0cAbq0qiQrwDTVQB3qa
VOzxJXE6kXsocM9wOmStezjhybchVkjMsCO3UuWa4sQMvYBbkTS22Q99QHDTvHLk
WiH1y63++xBwFRwZJv7HCiEgMuN6EMS5Moe8RsDzrK5iVWYbQ4zg0vrLD5R5u1FC
LnxLL/nj8qfCjMQQCLD7DIY+CMI3vHg0ihMy5O6KmUVMyH9hnHxkBarpb2dZVRAS
FuB4lnP7lyULEVNg8/dAzRX6yQfinmtl6ji8/H2Oid2KdKfEb7A9mWfOxfF8EELO
NiibqHkG6th/Q5BxJLAhLQ2OtS0W56PHVt/08O3ShF7wrJOWc+cg/jfKdZC2JZBk
5FwNKfZtpjO3hxfYYVWgoia4fplNrKTeXYhN67OYpjjZqL7TNo8/7zupt7iw/0Yt
6STmSeNfj2K/C3eX8/ujXmBxqvGDZrurz3IcB0LNf34mYQCI76wK2LbL4BvLPhDT
Q5qNrRJRTLZWfNzxlqEq/DXrF9cct+T/QR7LisD4D4EiXBQohpEie9vbzUHU9z7D
xMSKjG3t/QFnkcfKSo6jmIekUqZ6UlSn/f1X8Q5qA6t370PHnl5nSOM8apPfuSg7
3xzNIWUN1TkdFIAs11/PvrDWncdColqxRgR2auKpM0RihCSub29g0vEbjjFLKIXv
oFjoOz7+qT1NN/1/LClKEZpUM3FUk6Jox2xODzewb/XzdEJl/W9s8BJlCR6tQl6f
ZfYMmN6wVax2pMvPGnh9yhZO8oT3SqRhyCV6gTNqBfbbgV+akq+KjwBhhFGHg0IU
xQONORiDbf3mDeRPqqOnt4he8RgCV5fE+BSaHITYdbVDxHoMt51lVVeARM4sTtgf
pwUHU/L/dJgkGzi8gm2fHlRu8G72xpVVnizfKCvN++aMocGbhetKIlu0L1/BN731
Asz6Tcbx9CxzLvypdes3AjCOQqCvng4zrmVF6tgj+P3aSbWKMP/OnfLBG3Rsld1k
WTdVnymFlxbA6U3L336OV4DuyUl45GWJHD4u2qEr9EOnhPXtqjAoWfTkdXNQKw53
YBOz30D/euPlhGjDYSFFuqzgdnKEy/c6qIcOL5CoMgWJ3MftsgrgPO86f2NlkNcB
2TwG1jRYrHH1FhxLXLMXd0rKdOC4t+MeScaCU6Bls4oghoj67Br01N04R0DeF+qR
RtqY0tCcN0rt0LYOJqGinldWvX0BTvSqWtKFVpJ2YcgfibnoiI3Cw/WAh9YUBBuo
seVATKIJwgaweM03Jnm6+VGUs60lx3rlGY4vDCRBriJ9TOzLTWG/9YO0HTXO3h8d
jgbYD6JC/NFm3nE/sbxzWJXmCcI8bGokWlmzdA3KaFWTRII+RXZXfsTdWgzNyCop
InowCJmVbCJ8ToHGmbb8femChMqZ6u6fEaCpwCAMJg+VrYtY8aVo1WbhmaiyLMhr
LcLABZpOfivwBtOoTWMLmgNuAMSzpdeCnT4yN79Gi76d08rdnpsnhOvz/06QXum/
4/GXkA4k6m5SsbdLa2NhmBozqlcPo9KiPs4qc3fKR68/u0IeYQp9hc6ym3bQKPYc
wR8H+1vIDO+cPf73aSFxTThmNSQ1h1KM7XCXbp3RDmPo7jOC3SrVu4I3xFqlW+Er
gVJAOSSdaiaZijAbhxE1k2KfBH//reg1yHxenr8ICLPD3sKqp5pVYxcv1EdEOdMf
qybUOQYe8ebrYh2CoAgyNIVzDaBOtouRTH37J/9Yodw9HRRwfOdYxVTVUsCtDWpw
UVQvIPBeqQFlShJ6bgtCL79rxY/BC02JKdxxqcmJc4l1/m9b1n7VzDbzPeDvWcIu
xNpQt2FvM/chHGFEFewhimVzsOUmmYp/heBeWxge7U8DwRuocFOV2VUW+n/JeCnF
/el6ni+kSJIhsOb2ajMvLRierja1ogN1+OGrZOowAMtpxk4aYKBQYKs9c1es3iSh
P+Q84/AuvoZ77icCZvU2lSYT8k5x1oF2wubtiqhRkn5r620KWTirE+mCVmVzO9aP
8vSR3CrFF/1tngq6sWEe5YabTD4K6d1RTYmWn92U/s9ZFvLaR2FAew2pE9wdvMkj
ozIqO0jgKCdhgMk6+5tERsIIOwZ7AfZZLLRvbJZiEEM3jSefsHt1G0xuxWju8DMh
9w0sqxEn1kooiIXZE1raStBps7iqcKTVZkm0nr4bYCIMOCSRjBPUM5pml44qM07c
RTkAVWxFE+fY+gtZoJOmUJ9+S6F4mdi0SxyxDtspz3znrmbFeZMzVw+jhbe8QGO7
w5W7QzBz2d1bWKbnZ31Z7vwRWQTLYzT8VPreEpko/9xYdxmn2mpnEUiCem4nC3K+
EE5d3/Ukx53ioyDtz+Dpi25XQ4g0Gvfe3JujV0vAUfVXNNx/Wd973Rh+Ww39T9xe
W1tc62KcFfO9bpR5KzBKa6apAc54HdF7/XfJfmSF11D6+aCHORpVS+jwcDawPFpl
mACVS3BuZdOz1I/k/z1UITXUbS3ZzqnpRChLryLgz8zl0p9KbdoRW1bKK0ZS4Uq9
9z3acFkvjbN+S/6xZkUpbQLCosnLEur1Kq62rO0nX8GYusVQ8opW3iOZyR1WkLAQ
1D9+17DiPlRXV3kY+cDGVs+HTcOglKKKBUxwFAVXWZaHmaPKMb8tvQIw/0FhUYVR
hz/NVdolwv7mDMOiycArIbEiNAPn10dx2nOMXhpAMJmRfQo7Mbrl4aX9UR8bCwca
YTmKPvUvmnNgY/H572uIvkLylOaEDmzDPWKonhvf67yIjhtN+rHDy7WhA5q/NvMA
zi2+UYHkKmJKulWAIk93+l+vyIlFJPpXipWhKL/1SE+BeMKi021wfSfoLblJ2a9H
G2GL2qV8w2xcSMDWELEqjGk9gLsO8fT9SQBFYoozys/SuExCVooTLRmY6GotJKYJ
TG+kXN/hCFznTv+IpCSkqjreTIDqTBP+KQx7Lqnp+OrwQ+GZfisWObMoCfLIIrlh
H8cBiJBT6eQBKP2/781n6Q7qJT/Qydc8eDHH89O+v7J4KJuNN341QGDxAsxsq4aG
vXcDOaAX+rcazknkxUiQkGsrSrzTwqKZ+y6KdXvzzcDZC6S6JsIwZd0yF8810yGY
dq2AUOQxlO4bPWLCbzSXumIk/btPeCLYO/p4eSwd5O9AxfcDN7LSoA+dY+ylG1uM
P7xCiwwOMULBovBlXH0SkeGUh7x6YRzrdkm08P97K4CNzk9AGoUHhrQ5H1IOY2Nw
eraS8Z1dfFrh9qkOrDRBOiaZefOj/nY9qsmb/Yn09thxSztV2xOPhmv/TW0Odr8W
dTQbBuw7S1v5OQ+Bp7/61h8erxAYVvk9uwwd7VC1bCnrp56ww/8xirq9K+ckRV66
KVd/4bwnAtirPjZcidhU+4m5RdVZQgiZnoyKPsr+3nz2EtJjGvyQJoB1Vk/Hxx3S
47JHW/elSMcYbrmp1DU4Z956KiTJT9UmUN+DHXyU7R0P8l3vc8IX7THoFX+LrXZy
zklzlcwVW76sdGGmvfc6I5lduJ9CaP6BoMm02CDaAbVpvgXA+XhNas3jp93RND1N
cKtq4u5mAJR0RFMrlKmUknilvcqh9ZqUFzDB2SLvZqXCmaVhzwdaHdr+DsLAQ+4R
0j6c88kcn+weiruOWgzuttHvD9Z5d9KQpxuOg/qEVGIx0wOOxkSftNkt+wf1tSga
wj4VJXaNFf1ESKtpZ3MXNZQVQyscD+OZ3yzU/9pc7l4YP4DFb52Cf4Z8tWS99uUM
7dvWFh/DcYJymxFSEctXn6ZM/3tR1Gb9H5UHWdV74NeDXTh17BSywin2Zoirrxlc
k/f4M8mZb2jJ8+svtpCspuBuy0NZ9s2oD/qarWYtzTQWvwC1SgXs0+L5PVmVXrrY
euJkQFHt1WtLg9UJypvSUEu/gDlSLwb50d5G74LH/SmCauKT/w6QqphMx/JkQJ1w
mS4eCpYD//vv8FZtjl3nxvFmm+Qns+uLWGzZymB0BJM6l4X758eDC7hsfAPtwby4
ZZofKhmBt1kVXfCxopDEj6q/gXbPhLoYxXlno+uoHTnn0GtCfHQix9F8hy7JT1Hy
go7LeuWxLa80jcAMtE6p7cXK+MM2hOBtK8srEQ/MN79qJ6o2WHCTvchPFwstFFo+
nlKRU/kBs4QQ87Cry6i9G5zXMOLXGe5FS0j/oOBA5LQXGa+36FZ95EEkN9qCn6gu
M6wHRzgVoeBgzOb7Al5wsoy7DCCtsqZ3H7usSgY1dEwoWxK+RJC+wBs/H2IzTSc4
Uey2Fuf3kJeOjJtj0VUZmRyYhvSSEL+9NY94bodROkr+DnRnbgDhQ8s/dcWjKQOL
GA+g+xPuuVanPkAG4FO4/rvUr8gioBIygHM4Tdbz37MJohDksBDrpWR08aSnyv7j
3AEBtyKUdTsPXg2Ho34BbY5O3dZTEtQ43755d3LPbeo5bmi7mwIOkXcGJve4nbsn
PzsBXp9ORNDHQgvlpvbApVY4JI/dXEqHUvqsL1DBg+uh05GWsrlH45hc0593lYbn
DMxGWGXmjBv1+mnuoyUZ3OqHq4U9DplN3wNKuQ4dCdHb0BIIAPSb8k8xdVaRiaCI
pXZ/0F8buNKermaLkBNsIgLmYg/3sx0vUo5wZ+RwKqTNEW7po/6xoTh65CUn33OV
Cl4VS6p8VHDD/eiyoPpKJ/9BuO3aooG6ErAfpFpV9gGdIsy06HZS+8IUeXyRmO3A
rvDp8jtwnalykiC+C0whJd8djaWwC1azkNLEX4rM1J7zppfOh0R53ANOeeKxOrHM
D/mrFlsLdu0OBQIka+onU/40eOB8Ucx+vQWzp32FSI6Zq7NyPvtnugxW9cAQxS6W
XoPNCTxgYt1GZITdEbnKIwdUgza2jUZOAn+EOsFj1f/tR0MJ4XE/N+9AHTvO9W+W
qYFt9ZfKGA4ms3egDOBAdr1a9lsTIJeltoq0L1duKGysOtNI97rFL5oBHvt8YZth
F8bwzrL/pPY7HszNPfqU7hcSbLc9lQ+iK7VubonwOeEdsGypDi32c0uHHbwdk27g
5eWDg0ouCneEhBWpqh51sECmtEWhyE30CmFCj9kkA120uT5sbO6t8Btwg5V+Hh9x
/LcSBPSvCaVUW7uNSesSszs5Qkv+9qXqrAhvoYD5sDXcg1DvmEfBLEwf+Q7/CAaV
mfbUVhD1O4hLcU1K2hBcuvh0in4lPJHeM8owIXzi7bUGizAfagp5Sh+CFU2UlIOd
5GGKK0m+FMCCBrjy/3PD7V2YR4DR8OsJY/teC73q+lvfLcorliI70Q2C5X8tQH2D
Sezuu7mLyB/OE0mVth04NAGIal3cPqAJNsAiqB48tzYF20Rb9+hcV97uFlociU9t
bWBH5P/gVIxw0YPJALdKOYGP51K7hF8MFpoVWE1HsW+YY5rhNPWKZmPXoasAT3Ns
1iAl0qjzFyhPEq2IVYwy4Zze+2/vs49wZKOEML4LIgBe0RFYyE41hMLVRSUUou79
D5RicHGb1vwOTPHm5+lAcpfjYHP9wm5OL+ZXfSS15REGf2n6yMFyY3fc62y4DTMd
xcjA4RupFfDpYNxXx+qyQ1dgpg2hwrhVbdcgHS5WgPNXhDCh1dD+LyFg3iswoeu8
DinN9gVx7hS1DpMos6AIS3xoWkIFb3UAqaQ4gjAYUtPKKDEdTKv9doO1+q0x2qxI
BlMl0BPXohzn1p3uhbUHdWJfSQnSY5BTDQcGrmg6ebQg8OUgsO33LY6VqSna0pDn
Vp+7jSHYCqYDEDR92vYA2I64vVDpZxS/nMHF0b/6Y1FwQBHcOmwFtLZ35/zhLLwo
PkfWY8OOCyZOFVb9K1rOLpmTAGTDA8ej3LYqCWnDLGC3R2PisqyjsILlXfOQ0b/g
mbsvecrF1yH1cJ6WOUGjTEr81DprkV+0g6aw8AvyM4CrpKDUa2bWpHWvzpyoBeKI
YNgINalOSEGKyojlMxY5sFLBjoszTtohZA6KTAmhfqgDU42jeAxqpDP1hQmikROO
gsHNHnxsMqWIGMso7sroukdZbtlsY+FpF5a6+7ox+Wn2sxqLMcMGwuKwxyKyCHWO
5j3nhdpA9MF87NOOBdxkWoctooxMPZRNouX4ggSKG7ZbKyibaGUDqiY5hl+sn2Mk
lF9jhjc4iv5Mx8IIO2KG9/wEcte3QxtvmVWqaJxZaZ6qo2+XMSE/q6nfUzuH8F4H
t0G33xgh8wwi3b75IQM1fX6v2KiyN7W2aOssY0PpN36JbMf9imYlNNK940pNF9zx
ezANkVQGwSvKHNwxJtyhCuljJR617y2DZdJ2o5VCKTTFkcQhX0mYGCwx7w28Weyt
9V+tS1MRs/jtm5IZUZOuKirMryLJ42JohyyoM85+7f9Ttmc9kuSDidTJo4bKSco4
nJWO1LPS964dt1ZzgB2iCzPm8q0L8dTsfVVAru9JtTatmSvXZ9BSsZz0LtUBUV3o
oEI/EUsv8/gYm8pMEcx49mFjrTSdbI78KCp5O7OfT96IaRMyIEHPB/Z7l/btDjnw
coS2K1ENTDkAb7bC8n3k6dsCoB+WuBavber5M9BM7ADkAGoCEBfkVXifMyUVkbEF
D986JlL86pC3OUQUfLfKHNG9IUcsLlwihrkZjvXeBoz9QFpMd3FVr11EI0Rb6T4v
KjwdDBWjZHmF794dX3hwexvLUHKlRo4nEyVZd1UX8WbfRMcb2N3S8X/0vSEWqGtX
xGgmpKJlxowAIf6XqPNus+buQshoK47+FU9TPC12usxi/YBOGGu4YlagLdz7Ren+
GkTV/MFgb47vJLV86jalCwvQR/6FIU1BM7hScSp4P53CxkorWMZ58bIQoNATWuMK
DHinCip0Xn7dEKjGPiHqzVs1RAeQsl8+AciYEysh80dh0yZZMLa3Ae/eySAQ6FNM
unoqs6tnXLcQdPhyzrvkVv2TyYzlinXMGzz66TzpBdP9CRUZ79Bh7T6kCbX5UNKK
SwZPBAJPUJBC9RgfGheZteYJsEOPRU+PxLSZyf/RfA6eFa8dQibySEK0IosA5+q0
REd9QyhEVKaDxviRPyEIF8u/zVK4MoBJTDLNZYJoJJaz9a0uHdopE4E7Yfnfa9NR
oEFpVwZHHzXisRH6Jr1k742o8tcwhSR8apykwEMT8eDQClYwQyW69Nc6Y5jp14X8
ybwcdneh8t06QNkP1RMeC1iBMFGJqBhTkD/qOg0puG6XvfabyA2ynVz+jcuSD1FI
4cDDUy0U5DAoBnz59U7+wNIX2UxXk3JAifbHq7dtQCPla0xUQa0CZD0XfBJxaZ4l
QWI4v65/u+zcR4Se6dHx/bGdTfO+F8V9rsa8bIryq5oAvxTVabnWruFzsOugOFsl
N4KarkDMMfusCFpjg0kRP2NNLBSaRXzV7+yI70vro5xLSEP3bSgvwvQbC7oNyl67
CbGcK6AvyWKh6VMPL3Mcm2nQC6joAvbRBc5gge+NOSwF9e8eDPG7ADJhrm3HMHgU
hjbdjFsixkha8ODadvMfJvcfN9nPdKOfzH8PaaUQXysnVRaWN+k3i4e5UYVU1ATZ
iwaefSL/fGsrqA1iB63fKUA4ObEzrHfbo9sXUnRmNth5LzFeYu4cwuvLSibF8cEU
oRDyxevRmqMK2n8+wJPuL19eu41BvTdICL7bl06gKvYHOdXAtz0puAzGGDPhYAuV
5EcB+YoL+lOuxChnfVGSR+DXxWMWzbjWNdxCZc84hdsxmcFE56kMb5jjlah6ux+f
+m6X/lhpmNTVPKpPfo4oKukO5kZYDDdU/4ZUAnPF9TeOira2HkwNY+nZXSn91jLL
rFGPGumXX2RuRR4eJTRh3IRElcK/GNlDVl/8Sip25BI9SlGEtjxHYdxOkyK60boP
rqfbg5qYx0zSmDY/ISSF+q5MDKkoyURJEqGSka1r/xyzia2d6rqygmsDPRs9yymv
P7b7tDNook6A/Xs2gh24qcLH6a8WdSyjvGlbJnKBv+1SDo29G9tgiUwc2sr+veIw
YhOD5npTyiDNHr7LSPJ7JzF9o62Crb6pUf6k00MCdRLou+OdgDVm/sXns2RnXXo4
UL6DduwqTYIVcz5JCmvDRZtzOhsyqBXapc3cGLeUpKdaPcdJJ7bKdXcfAkrQXDsl
4vdfJNYsvZHgDMwO21Uo/3unxJMh0ngu7fC/PUwqUbQGi14I4If4igCNV1wFfEOu
R0QqW74TOUQtNzzC9i56gmoAOh4rRu/Q03cQox8BRzl/OKg6xuSROgGvQQ4fBVuJ
PkqkLj4uigWfZ98qaKMeVmsyuW9e+BkDQz8qWYy4rXPG1B6czGflkbNd0+5BcGNw
rqoKfk/Ob6eOtuEgknfmEHoPynCuEflmNipdpqzJltUrhibkPGZ4CbDCPJTU7k6o
G/lScB/wcHZVEYSd55nGK6tan8i3yaQwHHlYul3UhRY7Oqy6AhS9urbWPcUFQ68i
inIun+pA60H/FHJjFEhEALjPe3BtEhOBjzCDKXwTw25JX1HcAKmnVym+s5hi3Aey
FoLiyBqSZhISgzHVzkGbkW7aGPAy+d9Ipb1d2DAnaHLhwSmB835LatmaKl/qaCYi
LzLLvpaffX2O714mwJwf0VP5zuEIiJOJapAI6wkwMQsbzyEv9s0eJAhSIhece06K
AJOEfQDq4gCRHg+dJETjtUUyDMzCztOLQte1s26dum3wcg4+3/meVZ1WAVKnxwsG
fgdzTFlXEt+/uVNt6W8B/f2Om86xla5+1Tn38X3KPsPR9FakM8rtjrOQicwyzu8P
mGbV8XH0lgzG0dV13RnIXwA45NVfb3ch1J7SVGsOrJLaeTcj5GLEUC+cfgNti6NW
QYumK1CSXqAZeut975kur2Los4w5GMXu6lcGJBomiCMjLNnMxcG7RkdIqL9hSIKx
v1NWZSPMMofgrslmftZkLmZ1kAZFKQ69yUWoS/TFF1u42Wu2cyPmZ3ZOmYuS17y4
g9XdrNn7roPUTlvpurjUguAVMNkPNcDYx80vtRXV4qczeQdtG2s7yUq8olC+za8V
MvKWIYis5rhTkFCEcwupMjRas4pWzRiX2CbJyuvdboxVQee5AMJ6q85lNeY3EkHl
HIyLyQSTLIvfJjKHss39YWDaJfAmp6UwZwDAcwPZIobpdsp3fyNtHUO07Rq30kn0
c4+1kBoTsJ3ZXTx4+G2QVMJc7TUogoGORUE9MGfox5ycI2GjMxUvNS2hdAo1hbwv
Iig7WMf5Nb6mEBMUWOZb0AGaKA+TGyvsjLTgZ2hgfuhUXTQ1CvBg/lX0D97L836K
H533YAUzeyv0DvgIccJ7DsUsfKXaurUWVD29hvmLZdiZd5ByzlbmBTUfRP9FlDtS
qQWw6E1s/4fTvmYxZUfZSDZKHi0TyyTRStO3nWzaFS2Iz1BgRqorzUK8qnRzIUPf
lmQ6Q5TVSgcgwg3ZtIlB6uqmNHmHzUc9L0n+VRARgiUXf5YwEVzNOJfFzCAiLwfG
nsAnmY7Wf82lTLgfkacmm+T4JR25UbYjgHf/T0lftw4j2eQK9Gr3Bk8G3HVsWaTJ
KBSI6K/9enEA685pAuZJjvGiXMzJE+Bcc5rHigDo6mCMGX5XjrzTyMk8588DymuU
jL/v9BuUwqM+ggobZAj1jKcs8+WzTjZ1zsEgMdsiFSE+YW+5dpaytsFVe1uRuZkN
pBCuV6bvak9V4XqtdMKc7Uey9IGazCvyfYQoYVU6gyxdHF6uwy4PY5QoL9zN+ekq
dJyyiwWCwxYQ/tEGOOdBwQcADrydk5NVTCyQjacQLOD4Ngphl4MbfJ2BpdE3eh+Q
wT+fn2wK4KdPxDndQPt+/nfPgfNBL4sT++bKHhgjhZn7GVybalJdceTEgJQFK96M
IiR45w7aJg4LqxGoDYCo8KSmt58CmJnnC5phrB1DeiIZfWOZ0nj1KGLkjAianmK+
YYSnGZmQ1uorLQsogRSSNq91pcbrHbyBsQgoQA5tQ/R1w1EhRMdF/dV5gNQbAzca
vDxbyEaXSdwNSERq9BG06C3wG+m4d29dLtyT7gjspTqiEpaEbMq3ENJnmQNRx3ZN
SywHO0Kv9lcI0U04YcZJeafCHmVYyw0Uc8GPV6f7Gy3dqyVh2ilHG1+XkvPnB5Ew
vyOtEneQei3m7ai7DRQyzjeX8K+Q8NsUl3wOA8lB+lqYkfIDlTZJFCPNDb/QYtNQ
vrbD5THdGk+1GuSiay8vABFWSMXz87bR6H1Dlr/rhDIsKMTLg31EOusO4O0d8TYZ
vKDRcjn8gzKFq6SPKSaJF0bikm9sIrHZMnZ74uRVarVx8Zibvmv1NnZPNLNMslFf
OpgujBcPq55HWHnWWhX3N3Vb1gxG/6DjQkIjfIG2LsaOPf00B3lof0lbx96qWocL
Y0dVn4geJ8oYX7EIvEP3rswHUl1KYaDdRDXywVKBbt+bO0PkajfpHD0pBK7ir809
Fx+uOurYoI+ALRFfhzAsTmw4XfMuImmn294e3XiA/wt2G0KKb2VxWLzp0IBYJa0D
1pWFtQiWF9L5bP6PWXrchBPRb6Uk62AtXmeGvIOfbtGHded8eZSwMHTByww/8frK
zvz510mZ+JD1K1mj7Pot2S3UusT23Zmp8qhfiQRW8kHeUr0A6uh+Eaptpov2nI/g
TyMeVnkCLEDzKZ+kf/POucArdqgJmbPEg50/5+/lHgA9YpBQk3x/nSkbsCS8aY6C
Pw0wsKkXKCoJhdm2hGo6V8CLli0xGmB4WG94cDGHXEljYTGHzODlMZq4lg8LmTvy
6VkQxHlIJPUlk1gJFJ+jDXxKwYdIa+5W6nFTlJI6Jgi1wCHMzNeCd8a7dBeiVs3C
jyJqfHwhLqKPdoUBSWipwPQfgV+trW8YsvE51GAJsmhIdoM1hFafimbiRvJuawly
mI4LKUpwiGj0HCtdtAeX89V6q1TBmMOWEPJqaAUJ6r5RzvjhqTyOqPfyvheef0Ce
Z4sf4SV6rKF0cA7a9NMtb7+wz34VKfhbyT0sPttUpw5TwR1qR36+75SXmnG4h90w
E2J2DrzbFY73iMfalg2GVLP3c/Ri8Qqu20XlcPGa8OlTAXdxa82sysHpEwp73Yz1
c1zpD+j9nf2PhNAsbye60qV9I/R8Xd16lDRjhKoqq3TJ0gO689RnbB/2igVEuE8Q
Jiqsgt40hRZzZplkkGUIW/h2cNPuZNgWo0VkJfXjW+VhcPKaAYCRlIuoKDhYvN80
ZK+FhOLDoVqvLLOYWGJecb00z6ic/7tlxuLPs2r+vSyVelxzF5otm5Q9YJae8tFb
J2hEFPFz+KL8VYSuxkH5QMfT8n3rl5NiJJl1fKn3wMfB+F5dBND5Y3kiboeF+p7t
U5RI2ZedC5GM/KrSXF/IOfPcIGUqpLYPdn6D9GBYrrDdTnGawT6O59ftSBxSEi/w
DkfB5kG+9ZV+Y410fbgRW6z+wcpbl2YTeFU8exwCa4B3+b7inoIP6t3oKe87PHMB
+hVGRNw99+AWeLe3qCgSNFUJxA/N9JbO7mIaqk746v///xiPyPaGhuMbJFfcybLL
iQBTTExBqE44vOm1XpYIySSGZq+OsOyFYbe4616zQfsVbIAL/+YM4oiYYgznhNDX
Zn2vhc7bB0pIRpmlT2DAaNyxZ3SP2XfgW7mpRm9IX8EXnoG21PBOGuaH0Jq0GKE9
lBDGcr+uWkmUWg35yaBWGE6HMPYczfHDurajoKUogx/bcb0RETY9Lzn7BTrtwtaX
S4H2zZzhVZRSxcTP8tP2Pc7Zzr+9r55qZezUBsCkNa7tqwc/SLaxKiRajx9r7LTR
o9NlFvsgmmJFw7ZXDUJpxjmRUqYiAuTiL2qSJxBjPtR4D+YIe1SKj23aOZ8kAN5O
5oVLveTw6bnm+r4tq6Uq9JJJCQW6Eivszf5ac7FZVKh96dpXN6NIFRLRu92SaGO4
r/P422CY3HpX4MEDs6Zyzc9C+WyvcaKhe0BAiil8JzxgLjQEd0Pdv1c1GVbHEc4P
tEG4AwDV+O49cLgUEWMwzeI6JrvWVpDlQMP2fhKhpdt6gWnUX//eCZ7RM07wx/Vk
RWbG/VpD9UcRbyj8zjYOVrSt+4WNEEY1pMeL5gOq9bC1cJL+XJY89Avs8SiHyvWH
/utMGBcgAUv8UlqaKlGqfEKFbl9D9f0GirD7tDRBHxGch+r1VYzF4UtB1H7MtDy4
J29HFTLI6Roy2mcD2zVElmySMr2Um9p3VSLqR8YI/WXXbpoLhPDgjsDGOTu15vzy
+56XWEJyN1btfpjERTWxyOE6vZgr9QWTrlwy3SXp+hLts4KrxTlKne2e36Jye/lV
Y5aavoppzPyzczl3tsGYMd33DjJaWgeZa470s9rcDUr2SSdTiMPELWxUGEk6I9io
tj3/1Ucs2j6BSWnQWfGW0HOp4jANId/VvSnaz+tJy+gZtLC/gU4TZjE7GMMbmM1w
YKxkWIlKFflPEb0R+nemDvknhkM7NH3NrIFnTqSXLFihQ2HXBP1ZFDcD4F6Bfdfl
13D29dsbTB17X0IXO8hBBe8p0Z4LrEJwXkv8wiWPgnHLi0H11schgbzONB9x06lO
Cg0BOJj2itkaGimOCAWTll3qwurU/ehZ+GP0Y3+IWwscOE/rrvqYX408Fz6rFf/v
/aUIWGfclT5fxbtG5ufjpHyxtDzWsJjXG0zz9R29Vryhwkuzy5qIiKQM4GN5TLse
nCxpYJExUXYedZebmrO284ToLPWtSB2ZQDWntxyfZpp0YR9ycnc/+Srh+EuJr6T0
ayRNUVOWM9azu9bP4gEXajYFhWhE4NkVXjmqcezU7mTtsOMYdgpaJfOOFSt9oCgi
Hfd26kRRf6gzMzFceoQ2z2kk7gMTy2z/zzcKPk+pds6ZDagd7OWPh0BSwvha1vCo
0FeDI458yvZa+S0/h0UxJx/xboYzD2WhZNEqcOfyp8LkjKE59cAOd0y9hbiq9+pM
sMOWEijjyK4IEuQYzaYZeqt6eMAbiMhYU1UeIi4hiFztIeMMLSnTIEpBMB+L7e+a
sRzuh6XAm+ZfW8Wlr44SLPIOQh7Uczp0QG5MJXoLI7gW8OPS9BQWuyOtHjkGtLlD
RIP6Dv8eQeseHNO9U2H+EX8Coepu3JhUeY51uCWu4xt5fQbhg3VZYG47Wpf92Z2i
kxTxwsQBqH7+nBgwWahuMQFPaQnSOKOvACkb+XxiDYHtLDZKk6GXqIxENiDgFR3B
2q9UjKcSvP0wBTkchUg9/YtyUUlNfmKsEgXyPizwgb2F8aXkwRg6k5laHufKKVBe
K4MCtbsCkb9wq/sY8OPFfAOjt1BiXHKo823+WCjWt9Szvvt3/6BouImV6NWdkeym
1tc7gTFqeyH2gS6OmfkTmsreFhunErxTmg1YkiZvgsWCY+NLMPvOEHMrl3kQFHuU
1nENsvFktCH04IWZouDH7U5wGJoh2rAuNgU6LeoLnEpnu/TpgYsJL6RGEILhtLAq
oj31gBP9jNC3plAfHz+Nx8vYBHs78DS1hhA9cp02rkoy1nBO8sAuCVmSRokKg+vq
exoBbPtqPOJWdh0CXNNhpk0OtFEYdrd3f6HRz/eyk7D6wQ+LaL72T/sQz4Rctj3S
a6etFLi8s4zzF9/f2y0iCsAhcfoBHnnpsYiDeKKpg2vKGw6dxuWhz/Ja9uIWWviY
8ajuIpBa8GlwoOwOq3zF1QxTDakeGGTtTPoW6lfLXoJ5PA5ftRI8SwNiTkzcH9nn
8FsxYb2G8xHUfEB0gn7pnm6WNn9xS7iN2V8wnvrhKHsEvb5NG4lE71JRDFJzUzK1
zqjTSdInC8sQH4YKU9rBqlLbZLpmqsqskgEp7ziViWOPt+urN9U87jThH12VEMjn
9CHFFi1uFCISXWLXcvCb4CZklZ9IOPT2z2tQYJB05buleKExrWu9mBTeQB67OD/p
OZc4q3N35inBqXPEJ15nvpwwre4kJbiPPSEzCyZ/BX+HVngaLuMueiYB6cDQmcIG
6K0ZkZN1QwT+o+rm8y/cgCXSI1cvk7W/7aiV9JP5wAcguAuwofL4b9OkMDG41rOb
WBFn3IJkQ+F3KP77PVCv3QEFlwnnTsEccCdcb7356xY72sXfWBu3LP2pmkI8umTG
U9+Dp5EpWgiwJ0XXv23UVS3GHl9m1N5dGMUsSpwQOUom7Cc+u2Itj1KJHH5SshTF
ZE7ouVjLQsAV7jm0MiCLonqVFU6Ef8Etqj1OzYhn3WxGPz3wV+66SsJlyNj/uzsq
5WePpfMKtKeCiZKDvpWZOXIKUzc1Uxiwdi8SVi02bC7isVgncDUft//D1HvvgSpt
eP4AipzOhYGovpqC4fDIGSndV27Bb6/YfSG3v+c7R3MQt6UWnE0eeeIsoRTHDwBU
3StCU9s/5OXmLiXENSA0Ex2Hzxo6+2qfathINeJxSt+vRSDLG/XQmdqx0S+bz6/b
yR/MbBozZJChj4bJVfRz7/Zh1THMSNfsqXt1Rs5bsb2mapgBSal319uTxiZdVbG5
RYuQZRxjDQWJRz8/iV9l7DGTvJQpF5YYBTWs4ZTdwBlWFfAZlMMnpCkmRjJk/0dE
IazdK/ptPqyVlfHqFMpEILFESScrhInxD/zwgwMtfnwND9F37Xv8mm7hcUPX5zKg
jwem/PhArr5v80imu+Q5wHGOaOeRVicPCubM4RaQ2dymU9KimzBMZ++EL0fWFNqp
3fZPTkB1RqZD2mVxABoUmBGcvkAbl5SaRszRTrfa4qt66kvuTwcURQbRc3kKYaAZ
hVWDWomh8P/KsGdK1HP7mFmsW+uYZExt6oIkaL52960j1vGZQOVqQuslavfHz6PG
9dipuPPwV3k5HlgGQmhZX8mzn7u5E9X6TgzAZi9lFV3+Y59EO8eZy09dv/45wOcU
fxiXvMEVoekH7y3PWLyS4AeKzIAOR/OzV0VwORML8YFNpXeY85ERSytbykOrc23X
AQhmdW6Mf5815TzOhnRV1GeIOGKlQClmoMjLjVVLXOixtzn4gngfpzHywy6tn2SO
2rgMmFK2XWUAc3Zzfcx/ob4FV7et+Juw5OqepYPkBWqF18vh+zKO1HYxvJsx6D/B
JjrXPHK2vuCbX07jgUiLM9hO4p0w3Ts0CNYYRlDL5av37tlRWobcyHCyXDauEnkG
1hzvP/mN03gV61X+bukcH1J/wPpzepXn/f98WeL/s1ZbaCzRqiT5O8o+883PWwp9
3elhC8HFeGool27fJZkSe1GeApMn4BEiiFVu9q/Qg7xgcm6FTOSwUxwOybd6WW4i
MXG0fIoRkDZYVT9r9ZiyEKbUZn+cRGwn/f5phUR1LNomU9jsFqsSkkjxkQBCqyhh
eqoHSm+n3OP7GJLt3eyHUMCy64rQxJ1bkAyZh54VdmRxDLi4+H7sqJBSP4dYb9iB
GjWloCveYx4mHtJXMDzLEQ7GmO3y+B76FTbULdyv3e8ePYn1fSMStVt/XxCUkD6l
O5udBoCg3syGPNrdKSIRBwZnPhFRaJJbui9ug3QYWDUo+j5A+Udkv2kgvRuzEVp9
SMnI/Qjy4yJNUaihNp/psHW/HoZ57VVLA2pSzXy09jaOuep4OGm84RzBsO7xcOD2
h5VSZZfiKJhRbv/dfpqGymYtjXbASr3mAea5MPWGj4vNGnFdLM0R1tM6RVxtxTVf
SbSTCfvf170wYjXwrpOgqqNVhrooAiuBn4ZKXaOEN3s57r6YicmJ7efu/d4Q+efM
S2oyB27KzvCXzIsWZWCG8ZX4TuJf0RguvVeX4PYEUps9qX7ydiWDiwpXCXx/JE4O
ujmzEHzOfke9CTYw9o8pYNUgxowdWjnWIec9Rn0ig4SfQ9IXZnn+N3/QLEFb2uB2
eXz/t8I83+8CJXoBO09KjQWFaNJIse962AsirgE4FAH0iDX/ejF1dwV5JOpcbhfJ
qvTPs4SOeNpMC2QZmCP0j9fOfjAMRmx4zDhvHlL/I7vdzpsO39LJ17qR46ZZTBVw
scjHTZ04IVqLl+sVastu+mU5HGIc8sGvwmZoWIrqpGlvV+pHci3Wr5dgx2iHoFx2
MtJLc9FLSeiSVadLLOd631usKeNUqwb1qrbCueLAR4A82ph8YRAxUTv+f0LsNPol
CisiJESXlGJFhunc2vnFU7L4ffjoEkTXtuSsePqXyejcmq1knG3mOimc7jLKEGFD
bq39qwYs/TzSorNz1SVwYPnb97mN/LOAGaBQDtpybPK9PRkTi+xK/P7mO3r6dR6a
PIZHH1mSikDJ7fxG+QBW2VaoiAf3tVJ11SSrBipWf+/848GgwO3ASZ1RgBFHvX3c
N41kCIWVipQKvvfWUL5udN6DaZrFZnyUOelk/2gBnIB2e+SkwWL8Ny6sS+Brj/3C
N7oWWWRJRCOKH3FtgXtNRkCCS0W7gzJ5k/UvxKIC82YIJB3MBt6lNZS2ywnjL5/U
aMUsREgBeeHVQ9h4uB3tDcaMLePjwv8PTo3XhXYqf+tstFug8SiFCIsC3nIVc/b5
BeiNrpFze9jzchLYf65wJcdjdk2HEL4d0X6lUy3VaaDComwPWbLgqgiXqSHII4Zs
eEzZQcU75uj8pEg454qrV3AyjtAQbiudvm4xwq6GxgsaZz5mIp3kdRTg6eqctjVs
i+GAOMGdB78SI1IFWUSIccRx2HwFbgttAUc0s7uDue6T7yRvmMr4RXizR8UpWZcZ
byhAKOAVFj5TIYO+Wo1rBtlm6VZzxT/C4A0j9qV52tLGHRSBX3d7/Y/7nYVgVtMR
jNGZJxKG6kie5NvtTZq3afDaoOYES546b4OryNAJ37xDIsbcNaEY1381AIMJ0UVb
/kmMcOwRKch5XQPdFch6fqUtNb7A8x6Pq/bnKL75qyW5gsN7wg+P7H7Ieolxpnkb
hm4b8CJFopAfaeV1UUPInGLt607+aXLERoNASa6e4hk/EoWF36DnExgcd9s4OQCv
ga+G+kipii1neLjqwMBPnA8k9aOEmylQsi0K4N+4EOTbs7JC+J1A/vSg6nawY5zJ
noMLxX7bdhwsOGzy36WTgbK6QWPwWioW0cYzIbYYMMgQ3pC3VaZxEUlsIj2fGN2Q
qDxfAyIamQKgDkRj1MtvQNChWiivLZvmNVKzYsooPVtQ4iSkJPqqSBSA0XqlyHVv
DbxbRKNd2FKzDFxrB0ylQdslGUn96cI5lto185+YoLRFEqI0ipUGpk2KmdVAwRjv
50dkB4RqaNtTraCOoJEQqHBHJvGvNWxl81L/PJ/kcWRmjKOYd1EDWPv9g+jzZ624
t4rHSzVrqfZv3ub4f++Zg8HKL4NveUmnjfECyR3LDbdZaolrbEFRYmbJoWcVV/Ao
omCMcM0hM+2gmIZ2lgwcH8IqxiG9+ePydX0vcQqPKv97xUBppfy4SYZymkv3D6p7
FnvVvhg4/fo4sFCUzv9+t5SuAuPQX7XEEJJ08E+K8g3CE7t5LD8aoGNI88wCNe5D
aPr5Wb9vloh+i7XHPFOq55cMrAAwIU2hi76frvS/8ziDVNpNjGGNLhoJJgYmlFgH
lgkys249JUorbusuT7/o21Ke6gfnzcEeJdTDkWzp5vCedz6WA4yYVjrv8lrQN24f
DiUv97aSzu3SC0Y2n+aJXDpnHF93ZBIdVJA8+HdzBQcXstwce+3mxFQEMwrCl5fq
1g6MMSr6w7RzOAgMcJY7it4+NcSzzZmiEokp6OeZPS7XgTUvRJv46IODCEKjPAKD
UCMAfUi+IISH2oCLrwiqCvXAFZxLa66zfp292D5QTmSFYpn15DeouFjPhyjVcdFy
Ea78isoC+fm00NQPOXmlTKmw3CJLRStK1yHD97hSuEyXrMc+Gu1LF8DVn8Bx7awc
TAe1lGkSQBvAQFRS8czax6X5ry7m7V2qD/f//20j30hC8vQUL+Xbwvre8/DMfqRO
plDQRsNat90JRk2wxKvvuUXjnrxXc90O7ad28wYWPeXZPE1Awtva/gmj3gjkecyT
4i0OGjIWpxKwcA6cTgeP7Zbyx1AyzSPWDP082eozuAP3hECYcTx7vZ0J9jkcPeNL
EMs3+DlfDbl3peQlqszm0RtU8q+R6HmdRUgi5PLjxfUE5tCj4XHcX48ZU9I9K2pm
tmv53Hk8sZv9kvA5XPDK5M/w4Z8v17nyBqEDeQPLxiKFj3utRNluGpLb/gqH/sYm
1jkpJUOa/Tt/NO4SGJrDa5DzTAdsxEC/e0gjlxaEfld+PmwegETaWlmUPJOIQKuz
wm9ux7SziGO+2BY5grQoIjfcM81mbpe0/854OrJJLjGoM+MVEeKOAjRGGwEsIXoR
sa2jBwehOJ644QoLHE0XkSc/X/+zYO0yMmug88YrsZAChbk+c4z2y83Mbf4CVngK
2FlIwjyyNZL/J4URKLtnRLzysGMSmjBl4QO4gZfIF13ovs+BBWudKgwt9LlREpoo
a9s9vEvK47G2dEQ7In2hhTgpqX8hPgFMCIdjCM8nHmbtzUbepkHBJg+35/CZWEM0
9qCQEUZQUagBx2naOeQWspfpPk5jwM7eHbu6yVHvr4/tLF7i0VBuH/rhf+Ka925d
7l+C57tByCSQLYs9ksq2DA/+ui5UufoQ4g4cUl2ksUeXB9HXyFQRu2V/X6+WIqlg
3ju0Sc+GBD94Sg5UtPAitRYnDXjBt3mdmu/amzOGGNX2ztl4Ja+G6TOp6IzkpkBZ
QmOfrM9fbpgVxMKNsxEhF3Z1hFQxAsaUGt3eiTAMz9e3mkQLCpinqunx8XRpLbvj
vNv9viIPKFfV212oMOC7qtHotjsjO7M9U0DCcQp1cWzsxR5VCuxhljojrTYMSjq8
QTFbR98quG1LdBV+ZHspStFSG1WlwTcEVWzt/AvEqHz59TFts/joNz6Wsj+tfe2V
DFDAPn5SOoR//u6qvcsBY9VVKQ4ygkAPMRU64cjXQ+17Z6sQVrpdundAmNE/sLBw
MsODR3TcMxSTG0VwmcmzhKXmcHo0BFO/ziECWZUTsGcuxvmq+IGe7/eVzO93hN9B
GuxeY1lrsuS5/CGMHyn29Or5FkpNIr9zczrN8IiViEpTR7VPe9Ed9DdpOOGW2A3I
cCbRLN4AXBtRaOQgXwcqfA+Y28THdgWsTJQ+t0+gKd+AXk7mWhW7b8HRR4zhpb2H
sSLqbWEsIvdZX+/qGIYxt/3nsqo1kxgPxdfjTMiZ+4IsT18Ogk7ONtO2U0LTo0V+
zj6rAn9ZgLxfNlDIzLJDlJmFxN7l5zRl8s4xoNJDZG6EmNa0I6VZumCU5f/cbDZ6
GwN5r2RAdWe1IgvSU3sKws3IYH3P6jNjmLpBCdi6dfR3IigqvZbBxdI06y7Xneim
3Wcq9mmOOlWDEOfxBOY/OrmPuTItwvIpaQGAWViNFCOhWVSNn2+WheYME1KLwaKu
9D53cgncAtikssr4Ucsy6rab98ttRjzmou1W338YPO/1HwA8VPN2/S4YWe2Juyku
lRhKPWQ0yXYHhtb9doeimx0fKo8MEUxhJaffIBbAogvAhQ+Glht6SVSr5cEGky9+
b72ilDvbZDAZ6sQbTC+jRxm60l1LQ/CS5hHMYJaL8GwDXAwwX1igGz0mrIVBijlg
jjjfJjhyydui5kpEOf0epuM7CVP6TO6ry6mGlDmRzUxQeunn9qqVsHTpPGn6cal/
qtZFrvDB5JijpPmgCaboX2f5xVYZb8A7v7HGSUUsXzYDb/JQ8qgrW70tn98hJnfj
ntj4tzSrfdZDQNC1QV0D//k3XP5gZxhkoKc29PEmLvE9zfMS0T88PzQbiDOHVh8h
dvmYVm2tA9oSiWSPLxx8dlh0ryC6tZNOPI+MZKE9NT+UxAzUWlpTMZsJ/cEKto/Y
3XdeR6E4V9yret9GgYxHbQoP7JCaMSDSt3o7t4/KjeJ5JR4LshNM4S2BFZXasOhs
ViaMEvR7vUjl9G4+phfQ7Pq8ryTvSQjzVfqfHn9dvgQVdohA9o+bLrMXI+zar01S
8zsrgEG2QpJMy/1+FF9j0Na7bADHTVuDT5kcKimlvB8xbHbzwLkouNzE16ysGDx6
I+kfJgb1rjBnthNnq6XVPZ9Rr3gT3yeP5fDtHMmXMzvgKUlRpY26JqPWHiSJephV
sYIm/QIPuDgiHYN3PtDki3q7mhYbPNa48PyxGKbh4q+bKElQojXMC9QooL53eQBU
jAFq39G1613hp8kYlWuGDLV9aFEFxDIztbWtpQG+bOUyAv50vK3U7lK4UuFviP13
U/Kqr5FXvn5orLGB9zYle7SYXbgQWk7qQmPVtrH1V3xkOlVw5Wh2WMNI+9t05ZuN
7EmvwG+QeEHUfKwz8aJcQZ1sZjFiC3YIRoPdnvZ3r63SBxT/kr9j10KLgROYwiNC
QQ7b3I8JVk/EsGnZ4mCpVoJ5BXkZv3KxBUtc/vUywhLR3VoK0IGK7HZe2vyt3cVm
+afh7SQBRpYH47V+mKocsR6J4HDrmg2+2n5E1QhjL48HtPTCl9hKwQAGZ2bOBZPC
fc4l9VrCwqAHUfo1gsQ61NrsVDTeg180dRrkJZI+zRF29Fv2Of+lEizRtV32XNXd
xRoIZEK3nbWpo+SMJSWyCyrHeuBeK8/yoFWHcblVU8KoY8mcWa9h+DbXD1r837++
AnjA/GAa53IIeFKiUQEk8tOWwuXgdBLuzFlI3QO8Zoohw7eKyzKj0g0ZMEeQIoPA
cJGB7FTryw+2yxQu25XY31jhxMy94r9st+KmSEa8/sn8C6JqcKtY/7/cQ4Q1+JXS
mPADxaGIr0tNa1FjOlVo2qfZuuFdJOMkbqbF04jmA8gtNJbluHSn7jxDTWTZDQEU
O5nQlVPi+dWQzZbFNjFliwWg4RL1GbOX9hTbJoX3QbAAyF9idHfcwP1OXh5eK2Ar
9RrN0NCiqfQZ2pdrQnOjoKnYxfwKEnyV/7fFBsUu/Pz3CT1lC7/C7f0/Y9hMoP5O
`protect END_PROTECTED
