`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+zbpvS3fkN09qVdCQqUDhJ6XzlB4DWI6cGNqZDFwtjxSNnuykMLM5KIUbgAJEqFd
TwsD0IvtI6Uw2k5PnyuMpCXIA+vxZFQ7x2XO1fZB2jThcW1cDOQ/3+Wb/v9AfGTj
bWni6g1WvDT13tJKZS/7My33OKMK1xEFRaf2EOwk0bRRfzsPseFkXuoQqPJ4Lr0C
Vd4KgONw5ItJ5IWOzJ5G15Wwxv+LKzUMewHdvg99UKmr+j/VJii1QXGJf0h3GBgJ
nYHvJzUgSjPqGGPg6s3wkye+yjb/lYGOKEq4Ar4TUm4jB3tw/dIEjvHPmuyp9InO
InCYTmOV7aIKd0mIeUN+IDeNWwwCFIYI5bNsovxR9nAleDos1DEh6mJj6Ksba++h
N5fuZgE8pBm6Id/StDJ1ZKzYXxIEon8I7+nVBku82AD+mUidCL+LToJvYFot9KcE
0l5LEC6zJsZuLJFqbzHlToDS5DffePqQ6+6njK6xRdASjuazzf1eKH5OrW6afhry
ty9A8P3Y3gNupraRFCuddaasvniN8zEMq+2UwBQg/1WQtM7WQgcv5rQs/l2oKfqC
btBC5WQoeM9+300sCIIzkzR1U5G4C9zZW6gJZLXmySz4058FAJ0DfB2v8M4Ncc+h
8p8wofLdcVFNEHEwRgUyBZ7CbA/PN2XEJ1BpkPptReZNkIUPKixlKiAC7TpToWbd
zfHqbmDGXT7D2RLLiZqnkQpPQFhvzW4p4aQ5yIOu7/nBmIH3sFzHIDHF41ibt6Xx
bcitNksYDQB5QisTSGhDF8of7pLxCepspcyJVABnayelKN654xLyqU/M6/L5qY+q
22dP9b4bhkQ6Ra+FmOGEc6CoIZ2ZIPXWnTU/aafTldlQkbT65JiqH0fHFzzuG7Ih
hgDx7hKqgDYfqLMtovd8QlNMSSDHVe48dUJ+DjPnq34igCie8bIz9e2nizNJrStG
nTX8JhCjs1HAr6mnX7m/potMIMeejZC5pdtIPp6BCrDO9bQT2pZh+K6eBHDZSmon
QhLYWkHsuEGITD7MrUBZnwsL7vcUSTu0DTAQBv4aJiYRh0R7numLY+6hlEIU72En
14GEDAf6txicfmjSXs5rtsCnM8ay8Cj/QFz5bEhw0V6o4WOMz6oN6GCWgJfGXbU1
RqKhH+x0SsPJnn+/TL9P2CEiOpAU7SiuPoZTB6N85oyGMu41T6Lm3Vc/SKaAuCK0
/b/qj48ghOwRc1E3jvsal+srL1yRVoaWWhTM0shxrc6rCtrpaC56B9aJZnl2kpOj
2S7uOoc7LXpyU04tCRwmICHixMGHc9U20a/9Y8P6lPYCe41s7i8vHIhppDedzETE
JWnSOdF44lpFDCUg2IbhSE/4PKojwxTGEj//dI/oY2L9o3cKtDuEACO+6nYY4w5p
j5zWimx4IJHgLkYnkP3N6xNaJGUDmfwFh0r9b02jcb1h2RkKO6bOBCcL1zqkabq9
IUqYNeHqz3T86w65Pv0OcSWCHOVXoskd4iqKFZdBBWcOp0d7dCG3t3Z+grGGrwvY
pwe253bOnhIAu5bHrLdgBb/4VjOO70bN643EB6g+1nZhUut8ytybJndM4/xWD2qg
84Dp2gXKWEMT6lD5UgdHm6wk15vAX/tgLEEca96tA/X3++wzu9ZfiDDTb58NAUYm
2vhHvQPRgFZrgfvhnECxYNJ/DQUaIPUxL+c+Yzeghk43027rnv4ZVF7RJfigHpPB
HRN8LjCcdcqGg8D04Q6Xwa7pPb+/j88dvj1MVs9pQZ/iMj3VH1U0AXBd1hvo8SBm
vQo6rp5OBFgPStT1Kxmim4WdXEzCIhJVf1Buf4faoKuPLsmcvOkiChsjQdEob1HS
BVh94uZAB6HVt0erlt9sNuT7fRqahJ3iThyZEr79OV6knPko0NnvK3u/0VrHCYca
hEbIZF7YNlWfH4wqNYTuYqA0gpbKSFuP4Ce9lhRPUqL9SjT1OHkPV8IT4cODfaQR
72//6LKrYTJL0Aut5iiGZMHt9FwUArcnVOcfGMfANY9wpNZFzozN8aGKAwJRvK6m
SzeeKqn7A4hEJEgwmy2bA2L6diBeuz9lIgcLAN4UH9CkkphDN2fjSxH/E/vfdaHl
gDs0D4xYXpb9T+HW+ESjlw2sWYUfIaLcnnHgv03RaDSwfKxFBvclwzLwfyTlq3P/
EuMZQWfhl/WWDe1nBvFYa1aFYv2PLa9RWBBH+fqs/9cAG2v5bYw8d53aQcSCLfMp
cjBqq3xCE/D834YvNb5ossgNBcPaWrz6b3+Hao/WL71GAqk7uiqdXtM1tFvwzIEx
gXOGsMUoqQ5SgKVPv7btLHiE6K2PhHoZrjVteznpKSf79K2Cs7kmMu3WIw7gYdX1
0pIoSKandauxQaO6V0U7z29cvjHiErjBaLqMn7AUqF4ymStMAzbHawcJIrwDd90+
yqf+Hl5zO6r87krrmnvKnohMaNc2RBG2bMnwcgIRfA9ccqJDwckfyTez7bnwiLKW
DyhhqjHPfCrRXrT2mhEZiHmdU5xze9JZKqwEwp5hlHJEYRuN6ghB+rTgrmC375TZ
UywNBf6KzAdrJBB/QWaKFikjFcwF2otsaV5wZPeImSkcyaKeOxaajSBez27FZs4g
NsT1PYVosOjHsMldF+sr7+Y9eW2wIYjLlGmc7JbVGIfpJTWDyuh7KYRfikYWau1v
AszkQMMdVJtx6YJiKxaowfq5LovAosmjxIwdTZ/y2EiSaOuw0IFw8vDq+gLTDEHq
b4+gX/8O7/4n4EfOWCMnMRd6OM7T9SPKkMfNEH0q7C+ky+6tWA9tuykVK+m5+tc+
sMAAiV6fDRgeNdAGCgpCk9nG9BNESDkl5ksgsuDcjiPZryjAYiiDmvOym4hFzukz
jf88TAWknR3RvpU+hBvo4w==
`protect END_PROTECTED
