`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kkZNk7/4ndykMF4dWxKg0BFuFCKJKRxclRPELTVrAcHKJNrphiaI+83S3nUPWq/p
XpNa3X9QBABqjmkmxcueQFYb+1G81Spdb3xRbYEjMQRtcseToWi0HiKXMfQkYkUF
sJ64BXJYVg88AgiPdAquprhF9i23/i7zb6h80Hrw1xFHJpeF7s3c2dmEs6uSCV20
hUF0YMADgZ6uyH4qWOla9zjsxmovXXHWmrSb0x6gyf3IvQ/diSCJZcIp3uFvM9Yx
d7t9FmskKstwXjBzGfDOg4MPZ0BFwUgtqLCejiZVidP51V6san8p51byJfteUSQE
kh8zo20tF+niKR7LfEDe/Y33brXnZXSMpd7AXVS6qmPYeqKfFv/dwNa2z/VK+tza
goZQQ3bKiY6IusWrR5QMXYtKwESx91DuTB8uzMTTQhamqM1aiA4naWCFX5s6wPvu
VcQ1U02CE9634ZHO2LyLAjDlHnBJ5y5vQVQq11YxKjA2coXgahpTK4cfE98ZDSW7
xd9eLtLqwkFtUEEZxzuYINZk341q+BtmPY790TXiVK7AMTDBdRKKSRSa7899y6T2
A8N+UsMcyTWBS+RMPWnyLyARYCnu+tdMeVXuCTpZwd51gukF8R2Y8B/4zZYdGz3b
Qsg4INhPCAZS+eactWSFDJQv2XueewZ/xA+fqPH27KHznxrLn5eiHUewdPI37/tu
mMNox0xdepG8HG0ed/9fxIxsyZrfBoNcr6/SCQ0xrHCbaRgpXDG5l36SULO7RBkw
nrwpboRSYUNsq58yOMUhZQaqtNejNpjho6LJu3kvcBu66zz8Cr2OxpIVjONxPYWK
xEDXVAmk3Ic4m3t81E0TMfDw0AhRIbDpNhjuHUzTx+zTU7rrcdTjOgkywGL/jcy7
Uz9UdqD+4Jgivt1vfVorIErV4+zZEeRTbDBPTPnybvWlZQCP2cAzWsvRWlAxRUOn
oCHUwzAebEkqPJYxMc2mdweHonJqKTeh1QRLvdZTmDfTFaDiwKtvUGqncTBoDv16
lX9OTnb+hwpYJ2xp36NzWSIzpeRt2gNZ9qxr5WjGFlstRKG9I0WTuI8kpsmMkLKs
sGn2rcFxoj4pu6JoE8ZZ9YJ4PUBD96OYCFqSqER6+z3/VdDQKNrFE9CJ2uR17INp
SS3baePUnOoKtvQ4y2fbvnS730oGahU7yZD155B4+2J1v3Okwdyc/xJ26hEAz4/Q
x+dSYrtpowzYJKclYq2qplp/+lafeGL38vOqTDXLdwdSgca45Q7MhEsum2Zo2OTJ
R5D4oNNCdgM0DMgivyhPbessohHDy5ayLxvylplfz5j8mlPLtffp2gWXddlT28dO
fzjzFxxKvwcRAfwbmWcnl6aDzA1Xt8VjJiS59S7FAaN2W0uPkvUMt8x/yyXmWfiZ
j3BQuUZnspYM66KO9Cv7B94tTa6cOBKuZX43XXdw9Nz4pTL5Ljf1uDmMGDMdg4VA
9cjMupOVzIM9I4GAK2z2WnI4wgFwwiu1bYRMq5CInbj580KlLbxkdcftovPImu8g
bCAdedcOazdDrn1wZnEE4GDb3rVyOhBNZ0eUGUfQgqERbdmyUIhFSCQipYWHPHsN
Se3qVubA4q6P8HSULjLX1ZM92WBvTLPvgUkqfK+knDzs88RT3kN+pQxTw7m0zlSZ
c41iZ354/IC8yCDNbY7GQ3O/a2ea7baFOneU2euzt1wVFY01d3ycqWSHwW00IfO0
DUPdSs87Xxcy5mjZ6APh5P5RayKylG2jnWbgiXwl+FsAwGiRKA+Q2OV5ThNjl3ed
vZdiUDJWc83My6traMWf8DUJ2wGs9GyP6rReZ7WvwPYLcSbOofUONZdT+LALuK71
C042Zz3WsB6pEt/P5gRpQZxqp0cU78r9k3PSqaH1riWilKD6ugF4xuLwxEklRahJ
xXO/VhdtvDBIVEHt+c5f3/ga4ZmLHxqjpn1RF7ymB+5KkQxcRhbH7wCqEnl7pq0E
a1EhLFOu9TiiMdJ6cij+pGPavRRUbOuLkGY7UuEpQlOY/Ktm0Y0AQ7v8HL+yMvRq
UTyU9xBl0A0iUEpgXjmvtlac9Tf+PwIWUffAL0VNV0w=
`protect END_PROTECTED
