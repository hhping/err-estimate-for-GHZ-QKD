`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VmftBjQ5rcfji7tzC4UbLFyF5ZHVmP45xAyy0ts9xyWqhMotnZ1bxXtwWXrFNNV6
e4WnkwokSmBf9QV2Tj8GBDM4C/a5Ac7pzu7okeUbEpMxLhOP5ATx4MUekszTHbA7
LYrKmOjPQwuC+keyyVwgztkYKQvKQV0DO/NZyMDMr/GBZ0KC16PQyqi9eqiPk+NG
VSeKfSnR3JNGS4zhLm3AueG+SGPEUlsMTLXp+rBJXvIE1B+RGIhK+GnpPQqdKrdC
0i9GWIdhRFbzp0ADJ/RJYN9+Tz0y9eXXLkBYldBSvrSL6Jy/3bNR9OCvwAXZf4AP
zMAyauQ37u/a+Harxg79zWOz7DZuQQfEV3PGBmVqDFdXh9K2p5WIwg/5iDoWjReS
SGL8DZxbLMoXbf0RTdhjVjayRz7vXTG5lCmgmX/Bxuh4rWpWOsWJ6B9auuBWR7xk
+9ho2725RfokdjmJHjm8UldVDRfbSFQbfYWWi9nudGwpc1J1iCw6QUKxccF2i4i8
7UDit7JFZvdO1sZlVNjJT0hLjV46d4QXGKiXbwN5J+OC+ODFr2luBUXWCyJ6GscK
gmMo0DFe2kbxR2U5fRHAQbCgxqYu3BJWpVSXS3xHWrXT+FmgkiEG2/Gt3ic/eEhh
JYWjfOCLrrYJSNFcSpcz21BOOWYq8N+vlCFRz9aKj0/AUtumOJVpYFpptMSbL/LH
vPcHo8mCRJKAE4522Hz03yJpscuBkEjYAkHi/MxsOR0/zlWZuSQ0Mdq4r4/ZLlB5
Ikx3dDw3shhRBfcAZb0d61CK1OnJdKfarLLAMEU3rl9Z6bT5KJtrcRaxK1P/M2kk
RtH3Ys3TGICdzkGc/0DCoXZHFSfO8frjZMYYoPOawMYCFUd31UZ7QkxhgoUlPLX1
hlT4ILQC9HkU1uNAPz6xWzRxX8adm/p7B/NIwcGrFidVx3bRPKUm40sfMHS6GXEg
0HzmwlogqbF5PoE5DxTDtgGKE1i1ZmknC815SrX4FrnEXHvErviKk3chY4f8DLyb
FUSdiUBP+38uSJrASjlimY36iwqsbYn9JI0FwLh/pVauM3d1Jkia9+Fexy9JQ70t
XyYl7CJT6qkf2wnw9auq421vRtU6NLYurlbNUK4/UlRxRVuDMGaj+/5aAgXEYIN4
lbZ5yVaQKx1ut/ATv/Ki6LYBYn1PWexqxMqX6nSpYXviD1Tmt0Seu5d4U82AZFa3
VW+JVsncBxJ6wR6T1mLfAN19M53Rog5+IjVQhOnD8sLDNorVM3aQrwTpTrFGfHOk
yD/+gEUpz4QNBDNXhek15wazeHCIOKZj1vXV45B6inm+utZmKXO5XB5ic1Vk8Gn0
nGaelhWDyJc0cQiQ6RF6Buj7BtakakX/q5KksV6SJ+ploxbO1gY1xsxBN3DcK5X2
Ta+41K92LRWDNHVNIy3SnQ==
`protect END_PROTECTED
