`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KXLPkhGEc5lCzUKxNTXxPvfgYAzWpEFBYW3/9gNsXjXZc0pJiKBzN+oLSFLae1Fq
3CLo4qwmVd1836KJ+2Zzzm6eE/jP/+ACRKVn1vg89ip8UfkyUStOlX7sVdzxoqcO
puEfVNoQuMNqtvGRscKK5w4ZD5IeKEvv1DiPiU+gTP3LBkYXTj2Dqx9LAIjJSutl
ZxqOziXCVmUQNMKFLXdPfYmww8UmtAmy+WzYmSNweM5CTKg+kZikLNZYqS/rDtPT
mHSdeZaGK+n+AA7r+SVQirQZC/hNIlOCK9WbQrAjH9H1hVbCuFbsvyGX/vW62L9P
rQJTgWxVdzbPpp346qgp7l+UYKico86LERyF5sOeqRaIe5ynBGQewISRT4tHRDGO
MOcpEAsT23ty7wCcfcW9CU9rOhJyHmDEQ64S//fIZ+HAmlwhQc8j1DvOaym30/BT
ot5wVqotREuI3cHMug04dX4ta76xTQfh+ydRTQpPeiRswtvbWQqg5N6V/QNZ6g77
FcZ9gsMlA0YqUGgxfVZu3m4tfg6aGFg/ekhv9eX0AxXi9ZffSnA8t7TEUIflj60g
zvgfYn2DpkTtJGAY7p7UCaIP+pp06RtkLUr9sBPH6EMC5HI4jI8VFEz2Z1w6BgLo
0OoHDO0O7/Pivv+lf6Fj5GQA7mvyYyNG4kcZJPEuBqxTlcO5SNxmJtveRhEtvy4X
/5+/1BmFBg08m0o3WnrC//9wDEz4N7hNh3TdqH4tvh4N2U3RTe45RvgGPQZJjCGt
ttetAc2SSpHoUo9gnConupWSTFDU13ogEzf0hOKXh7/lfM41IGlD9fKAVxIHBHHC
SlxKtwXfxZuJx7Pz4Cv0NfdrDbZkUmGuGntMytddpr1RM9zBTFpaMPMalyhTWjY7
rPb+cOjiDtTjw1YyipTHCF7c7x2zoIrC2dVy1m0tapNBiyGPyNl1+UsRW3gIdrQI
gacYrVBRcIK2Zwv2zpbAeZBsMHIRhE8qYdQLqOu+/rZM+WYATEpbIHC2cI6avNFP
RfJFKpwGQxlyTz8P0dpaH3jWnERIe6bv67MCu0QTPyMNgJV1SA5KaDNF1WoMwQsh
P7JeixhQdnlnhv91NpXB4adYfLUYmFbmBCaCG6aWKb2FbF5Pce98vkk8ARe7vSEX
Kb5jmLLhm/4Vk02/iMptjmiwC/ystPQqzSESKXPyJGJuQ3XyB/EdUeNnbsHA+ebF
315MIJZUxw2UhwXkiseXTSmGoYDx08YR4cTQwqcsDOyCu85O/zYT5WCUDlVn+8xk
XZ3sqHf+ox/ipQO5WTwW20R+ZheJCA5YHWMoZrctz/L4cxtv4Scbj+BZFngGfLpV
ZgC0fCwWr8lCUKw3HlHWWypYc/2BkMadZUPl9Atv5QmTEypsU8DtFtOfbxXVk21V
3aj5YBiGljQ+yx+i3+FoKkwEaC6bB8H4zV5idgTxoRAnaOtxgMwiXQ/xtSLsTY/F
hFPLE9uTbmglQvep+wHhsG657wyXOVdWIXqpujGWk5Y5yEhXVNXd2IS0sgJEy+qG
EVleY1TwsldzkX12m3mW1/i2HgppO2DznS/2tJRf898JOzaaixT/o+ulpgEvN0Td
2oSzHYeAqJ6zPU/AkEfcBYMlv53XsUJhw1Aofrbe9fPvZyFKdFdwbmJjmkxIidaB
LZv2WsNPcPOIW/FtHztAnqpiBWNElC45YJLHvwUW0xVjm0tPO+dGsy01Y3k+uyuW
fPeSXmpE2ScWbPuGsso5whgiSGIcXJVQIpPXS+eYi0fbbL8K8fMclRo299gNpd0A
bFg0PtUmYbJcCqakPryrWBNSIQgSDkSWU3ZfSKcTqzhjIWM3RFCCc2asyMyI3udA
zgsZUFf+z9yPRqYpgPAblFY00/5n0RreH26tPYmLPKAnIDWykD5Vrgo3a4YU07hX
wokWPm5b8ttGhbWrJxX0fdDKfC1XyxF9lL+eHHkB5AoOSWcaJ3WPZXXIhkpQLIdU
`protect END_PROTECTED
