`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j8aRgX19ipJi2aHeF3jWVKC2xMRCcxa8+iM9v7Y5SGXO0fL7cnekpKIKk95tFueH
xdwHsqQKIFHthrZnPRtiQ1+IRaL84p8D/3CGfafvoqTndwPJ4dvEnJ4iswbDZwAn
OwvUlxL8kFhW2ftZApQ9j/BhcJSlo/iIkVWLlkcT17YZnXkWMlSJ/tfJGG2yrVoJ
9POHMRv3Pd11ZBcz2f1BneCWhK/ObvDzRVINnWlP/Q8z7Z76ke49L03oZy8dIoOZ
rmWyU5cxIScHxrQ+tYxmS+evUDhs1Ipfur8tTnoQgQMvSKuBqVYnE9OMLcrF3D3c
GuHqYIfTIhmX0dSHtEjuSAqmgbOjBrh+mg37jl38E60XXf/yskX5QUreEB85oTGF
r1dwxFrML1P9MlImlbVfPpGDe7NHGjAWYNopEckT7maOgG4o+7kA1KJQsflNzQgU
4BA2xQU8Vj41ZQJNfkqVK+p3I0EL6aZqnVagv12hOKo=
`protect END_PROTECTED
