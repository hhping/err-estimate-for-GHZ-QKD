`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MuV412ZzCQumwFELVF9Mdnt2BYeT+x974xYi64fdu6vTpPJ2BP9CCmF8nRuHydPk
QqRLjw+PyRlUterxrjtD/ccuRY2+uRE8KPD5X268Wa56IduGTnSvECWqRXy/0qg/
+7xWve8K0USb1g61Db1OBbpxtcJk7KnlUaZVX8WkrjAuSjRbE1C6KkRU2oSs2Bxr
aR2iGiRAEru1b3YimVo1k3bRa48Ks7/ENVj3etPY5Y7GWaefmd5fYLN4GF/Moy+F
Xwr+lFfgSJJjzSWohJ1Z3Kp4dveZKixeNdM59xX0/uyfYNyU95Cm/69CvgL31WDA
Wd2UfdkQQnlOTFZEBYSGQGK46q0rs0f5AokQT+NlPU9CaqQLdT0s2Rd9WiLEkG9Y
VAMtIqdI0rC/VLRga/MtADA1xW+bvTG4XrfPpS8D8TgPdR8/Uao5TUHbBPwZ1nOy
f16K6RG3foXsWGxRFeC7cPIonbZfcgsVIuSXWBYAa/IU4+yD09SpLHDlw2xDVB6v
fuCD4m8QE5Z/4+1S48FiBRJxCB3oNY9HNxYQz+ut+a3z7gEOhzjFKsCrTVBGsA6i
CuL5NaUgu/WxMjzLNQ7TQodwzuITptFn+eNpf3beoaKbatNVqJ8amy6inTFPBVr1
Gljh3s7d0g8QInaUE83MXJEW33aDwWYfS5ZVJNefhcH3OR2Kt80YX/6DaDHwUpIJ
8tYsJrjASHzQDw+dgZGPbAulxz7idB2HTfc7sIKQcoCyLXbyVyGBJFeJD59a0Px2
A+Wfb9riaLwXoH+sX/Gi1+bfZ4/t7M2dbIy+/2Zf1TAZI27s399DN5R3dFJ0znfq
/GxMNWj1sMbT9L9qvOUtFWlf+4f9IZxQ83qWSNPk+8NVMiIe8Ji1PBAVVc7Dz/i5
2ukRkQXLRY2GDYsOHIF0IjEDrQdi7QTYsQJG185UOlZ2Bhxd5o9SwDQOebv4mEmT
u7t6aFZNuDtOBmIpZufICCdE5a3TJrg15YhdePeC4jQCU+Ahc6NFvq3bOKJUP94D
daj6cwREHzEyGkIASbqPEr2dQmcF98ktr2tgQjfBeiIpGxUkH39ZYEBqTcDdg1Gm
lWWVv3iKJ+hbjhgND0hIasEGBrcaMrFHBqlM+dSBGYeOiDc0JdExRvuzATfmOl1E
EFGDq2TIFcnaCyPz/sGXBGb0LUYak57ef0p8FIwr8MehtqaYJrU6elJqNMWmMEU9
BQsTimy+YQ5YyRQxn7hfiuPrY+WIZ5yMTv3HY2WPdZ31QC7vXJKnP7aj+eP8Ru/8
o2Q5afiijtM/fPP+1+frhHXFCmOQpiisS8Da65LKvKm6AddBMhA3RYXUKMS+v5Kr
qiU7kjIhB/L7coxGc3H1utwo/yP6djvwLY25yw7NB/+ELk2gtyejURPauvO/H4XH
B5c+o7Ri0PNweMsvC7/vVhhHLj4GEFuHoZRolyQFJNS7IuTEnsrGZrojdqSk1wux
yzWrwrvVDu6m+9+YbcrRNBqBIpg+awN2lUacB1aBaJUJCvTXXI/vK7fJ0W0ARV9+
I4ZCZ0UtxuN5NtzOTNTeA7hWsOiSJTe/mcA0znnedojmumke6EonRTblL2DdqijJ
jv/Aff4Zv4yN6/aKesz+JkLKxSAEXLq5IxszEO1BYpwC0RxjJN+Tgp0nvs6wmc0e
`protect END_PROTECTED
