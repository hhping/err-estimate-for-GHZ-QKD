`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DEkFauEf5PuA+MaO2EHgcTvMWrwHUpslspJqhd662xECaz4bxQMq26dC6AgMIgAG
lKh84udrIHSeAq1OffivshqX6c0Ibn3uT8SRueVWiDUQKN434n4lzMvqV0UTUnYT
Q2qxankOlwfqYcIfEzgi1fxbFhSzX9jut+vud5jQYMIIKByTzLz3A1y/AxqCF1g3
4ulLsGYGZj53NbXSNYkWIz9hEcZWHrY4OKqPShsN+w5sLbcWz4+hYIbKGHLk9gp7
paaQbxmdIyU7ZTNGRD/LDaG3ceT0BKRe7V6maPf3YoIPzi9TDhhB6gXcijDuy3Uw
OCb40qzX5Mydcouy4B3JmuEnL0cGkBgJzsZNvH3hVhCu4JwzctOaNVvo29hr5yYm
OPSf1VDJdDAEuc6YONTuXnyt2DUREgmGkVlFOBFyJ3iUwkK2hJ+KxrazRMxP4LOL
E8ix5ZTtunP3ms73w9IHAg3CEvhXLLyhz2Cr3Ifn19FvNnCXuw4xCEnCtJFVomzd
qNzg2rihQcHoRaMt8Fv7y0Ft6TTYv6McCLmGEJuI8zqZwm2QupjNyzJQyKr1p3PF
4k2gBINOl6IipLzjqZT+IfbJpmNWXEYlQDk8CiDO4NsIM/kaCZFuUXXlwOUwMhE3
HMoUdtAAx5idhNkuTC+CHPhW5w6D88sNWm613aTv/fQxqd+lZYTgLulXsTMBYO8j
OYifmviyAf3PGtGqBxNg8504PrCyvKhdHX9uTLUDnFDVwd7J/H0GrYp1DIfiyZvt
6ow3K3gqueXV01kNndnT5jbIt4CC5BDtS3wfScHWK1y4mgdTQ7d5hBdT6oFuqetd
t14WjGW6n6jnWPeeDc0SyyTuklf/UHlbSBl0blTMCvwrN+fbbveV/rDKUqVxPekZ
0PENBx0i8j+07Ye8MVkKcAXplZ2mBIgc8EF3HBP8qbf26njzKwbWvetM/VPSgLTP
m9Tm5HB4PgHKGT2WPZZNLHi8SNrMbeoS2b3YViPGgFjIB29Ut2WhAbr4mNdUAWh0
5r0ED1aUs9tUkY9YFs/6sfG2RYkb2YscmNr7iPn8lz19UU143iF/9rmKpzI0RnNd
niJ7vxQIAoMii4IRDIsHkK0lO33Q/SCp7vbOLTd6foQpfrLdIJ1uAChwxM0DPC0D
`protect END_PROTECTED
