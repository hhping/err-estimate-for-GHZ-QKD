`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QtyYFEy9bsFKCnwVH6LnJ1NxhMA3zod0rrPbuwScusHQe3WRYu5sLj87JSfYvp4w
fKwXSkooY/pIUdFItOKv6/qfDE6VCVp/b2SRtdpvaG30/VMy57dMrYtm5fs2frOA
InX4a2w7MITlxo4VDHJoIfFFycovmuxkrZOlG87sagZ96DdASCDa6bYjxlm8z7ln
TRfgfZaaYNay6ULLMfI0eb6vomS3rA2gcGaWYDuSc8OHB/r/zNxVzEWGwiF7RGZU
0nAHOb/hKFx0rLEAR8IAzA+3aFHfSC6WZ41sRF6p2IfripJbj6L2HcgIxUQIE0Zv
9vnommsJJbPMiblEM9BnBiUh/B05548WDECLADIR5JsjO4WVFyRLZv/mpRuaRDMx
reiCLKA3quBKqvQr831Kdwxp9yMQKoSz+maQYRcC0eKAzZX8GzySto9RQoIzmaqE
11eLTLMSCjRdOpEdQ52pqzSkq+YRFnv4bUl745i3VUeihQRWxo9IxD3OlzfYncxf
aGZ/T7DCW/DWRazmWCWnOvm1d2gAmShlYCaVVoGb56O2qiFbbn87FBu67r260YSm
OKDfovTOk1QpkRC4+euxsSoyUrlqd/zEQbZ1PGehGFRYUa5qqSjnhRndtX8imBdU
pYyF7RsIwRURNH0xRmqxKM7J1tUXM92gG+NYJin4v+i5OP5tK4+4H7I7/IYzZOTG
mPe3Da86D91mKcwQiGajYQ13ZfibsEjNb29INIRvC8iSv1G5KGRsWPnZcr8Y3mka
DECsl8x0X6BTiJ0mPJrzl6nd4RCEJUEnHO3st1e+tNSbpeE2rC+hx/G4diK1R9qz
PGnTrt6N6nf+4HAzDSCWWfa6gNniyvws9xBRcW9R9u0GkEJRMn9zp/Y+kbd803Se
7rNyEApf9GFVOcNZlYD1J2ZxuR24JTrIvTjo1HctEBUcHS3BUtgla3gmBkcbs2uS
R1TWYyEmUJ1t8LZmzXgjR1thU+ewI67xYuMw0vvz5fOpUoGw/ychNew0r7YVf0bG
ruiF8XcitdHyzUEloE8Tov7qUEjWSA1MqxkrcQvmbXoFwkpzTdOleCpvhNY1z59v
LhVUs2TTpzX9fz+urCsvNJp7nEdey464RjICal58d/VI0p0lK5pnKoF0kwpBGXlp
SwiTRC8qfxF1eh3/Nf/ckVwhZp347C9aeS4XcrA3smrtZTDQJts41r4ARb80K3q6
izG18tP0z5ZtnLzVuH9AJd0iNMU2a6XY4HD7fykrQXsGItJrOR87Z/prtBJMF6iI
gvfXaQuPFOoExUEAjrQPU0dZ3HG1gYpPp0m8Ez96x2+cECFkRbo6nChZkDs5YwZy
7KG5HoTiuv+6mvc24TmXgIihddUGxtGoFLLDp/VyM/TouNbTm0eEexJpM2k7bggy
5KHr45aMfjP3te2B/ihaNKbQk/mT33Vmm0BwohYaEgXM7KBI2Hcsc6tdVKSMb7ea
8bztSHy1q3WWtBWHRMhZXr5+3gJ/Lm1Bu+DGtOo+djY=
`protect END_PROTECTED
