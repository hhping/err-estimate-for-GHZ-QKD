`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
53UIscU+rLe9Gurysi4sL687c/rWYshCqpO9GaoMDBqLZHN6tvCB8lH9x0fsaxWl
g+U7Jt+Kq3QamunCW3572V2khoQ1yjciNtE1nQydoVZb0yEH7o903tWLALfHv8Xt
LY1LeCMyV3SLCyjPEz6Oczj3kvfwbSbWPI6VV86DRws22/8r3t+yEsuDJ3ZA+GmS
BI0gBgI+nd7qVU9vS57RyONNn1GE3m6ki45oaAOSI1mMozfQrbQb9700ygbMkYyG
JyinxKzfWePlRd1GY6tDaVHj56qwUI+bA2JaRdBBNahKT6JvX0zZLa7D2MSyZ4ve
HL6I6ZNpx3Jv6vjeRn26T5bnBo45RsfoTO5xQuuEkQ1DKpaQMj8+zYx4j9NMsolU
PozqfTOQhY6Q/WjWc6zXVecRQ8LUCn9OAZ6Bx/7WU8SWqC3HcpGLp699QXy4of5n
hNr58gilnulY9QyG4ajfUQxJuCAhTlFLViR8l15qaYXhRygJhOSr3epYzKC3FnFV
BH13CnZIv91kVO7r9LJBxohHMKpsAbFUqgboWeCDk7VVc+IiXsoiwQh3qtlQTImF
7IFsDm7EHQL04LLPKByM1A==
`protect END_PROTECTED
