`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jicYzkPxk4sTmUoGnGkmGuU86ZmHAvXolrBgENA0edIiDrXq1PQznXbvfpt2sJ7Z
CGl/pL0LiNRIVlwj9m3qrknPPoKYYGLgISAuTnmayd8YepUXRJ0vpB2i9bFb+E/0
E7ZD1PW5Z8zEljEhK+BiiBW9MaK69U288wn8358TESzQxiwQagWZpv3/LCafdy+j
JyYI/sJ5hn+YOXVzWc+hOqhFcI/aVE+P5zCyQ0Wki96UB8NtGDeF+sx8xnLbV8R0
ijjKIr68sV+Xg85H+bfXnsqT907oM7UEjlclgcWpKLY5oghbTChzVlEphQSqGihZ
wdtgJzIsFEnZb+NRJIM0RjxoWe0fhqRhweX0sPm4lyAMlzc3tT4S/KdS4qdOPUS8
Ru/rnK/DIKw9GWRr9LH/RsPR4ON4XmTW61fD70Tw5XJ1O7Ikg40sTAlvj432ujMT
zz5TFhO1KkM72l8+yLUnuXbb1Xo+cH2qz5OOzDRMpTIqhDzW6NOQWHMfDmcAnDiN
yktPtqwute4TZGoL+kGfwij3laSVlQUGCbV61aw1KsJjRhwnk16t+enUzi4mq5xv
E4QNvXBw9FR6a1zt1QUjll/UC4dmgizoYOwmFlfu9WgouUWHjLdSRL+Ddgz4f0sZ
lV6CbSRUVistFHptyAkoeU/lrUbK42L6k6f6+JLDuDS+pq9ux3S+oo0qwOmVUbtt
AI9R1iKCfui//z0nhnhNLEKJWMm0G9GeEr8t24tDQiQv8dW5s/E1nN87MLAHdheq
7qb0idI2mZvw7+YPVtM/mrFMOuwDRGFcVzPgt/m28TmshfgIN1Ut5kRR4t/ey2JL
9VTxDPxkfnmHp/FHC9hkbQSl+1XBHrw0AMQavjC/AdeDCigjL7HrVgJh6GUTkoST
`protect END_PROTECTED
