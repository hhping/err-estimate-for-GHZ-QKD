`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uoXAU/EcS1FxYzNGtlwSd2JewxlXHf9yiVYAonvrShyLc7dlAUFeGLqBZdRK77XO
lAwqn5IuUpYteH4+liflLip6z97ToagE8rBTyba9lhKWJI3DpXpSXTaizRhV3jp1
Mpd5kqKYzOBBtwrASokDgWrzM5SYSC/iYziHFRAg32598Js5+un5hOtfBHycvTjC
cdWC+kt8i4EOVzd0Z46eI6aG/WV8O54bRqcxkfoahU+yZjajkte54VIcmUHCHaoF
YwJ/wR/i+iBI1E0PoRdfhVpCwfZN6au+Gz9bUKDSZzIfCg5ok0pMe7xX9r21Bgc9
N6aviRpQxijgRo4VA/iCmfnA+JcXzMWutBGAq/FrDtYI3pCw1emyp4YFv8CFQVDh
j+nyUAYeAnSjl/JHHmLBNgSOW+mtv14ogJzhNVz4DzjQRQNOfHhBdlBrnwILC2xC
zfqr7Ps/oQxjEG2HheNf+me6jaSry+AD9q2FXomGEC1JutTCjKMIo/FtrVt8cHWN
k2MujHA5q+N44Yv0iqO4BNQ8XbN/uhMNxUW/PDwu5oKuot3i0IgYzahwSwNGTWQH
BnkecH1rdQYGogSvsevrYTf9f3dDw7eeeyuwkelVnx4D71x0UvBsBcpVNpa2fRj5
YuFcBH3/tDOAobX0W86pLYViO8083QZ9ssXhq4vOWsPWvHuE95+bJ58jJUR/IRVR
EtSv0OAM43JiUzjLdtAS9tYlsItsAQmb8pQNHgy+/7qf6MfgmR6IWakhVdiurEJL
ml7CTHfU4FQO1hHfK3ROBAgKFFb/vZqpeD5QTYox2BE3IreQYPhzSzQ7ONGe3xI0
OXjk7rBUrxV6xJXfqYklUlZw+jnhM8ixTc0X76A2V4hpNBVgBWDAiV2AT4u9mYWc
yeKzsY7taaEA/8lAODqVC3Pz7utvX48MXCjhdHMknhRjmpmxKnaIe7ON3QviB9eL
44jzI0qOErxih0FPvhno5sCYv2LxJAA0oD8Xl9cG+IU7GKkpziFzrvvjeYRFwcgf
93xER+THIP2By9PmofVrAX+t3LkuNj+6T2wEzdK8pnpgyWnyzWyWzYmpRpxUye/G
LJhSXGPqQeNat2IZ75lSEl1GVmBy2Cq58g4B5arDxoAvJmK8wstG7M1BfHfSeNKA
Fmtcy7jmTO94uQKmsW2aVXRW2CWTlscpkdL5ij7D1a+SpNy1PBifleS2mJ76unsY
uTgUrQEULFsmnxnjIBAPaPIqpLx3ASbxNvcqVAZZWmobvqYWRQAGpnal5tI/QUYp
p8bUaoCPT67LpxazeiU5MRPpxgpzZBB2sODo9lZtfFv0kSzatZI7W1KXcNEIQp8A
x1YDBr9v7+IxIjJ59WCfrGgXStPfwWLGlxTljxZPWwWg6wkNLgBu9aeKUgNB9GUc
iEnHruSjVWeLf712CShdIL7nOMUyvSJmWG0uKwD52uiUlWlNnnJ9rL3jdaFXOkh3
bhsbR+5m0okHkHL8EHLDPhN9ESHCOPW7IS+DSivuppU=
`protect END_PROTECTED
