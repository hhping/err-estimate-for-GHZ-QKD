`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lu7qqVcsjLnUsuSMJlcCAL4qpOXvnvMCxSGaZrt+evdkR/DUseX3W1n4qnjNVdEr
GB1e5w2yR+EWc20ux21beb5hHYmAm9JhyTySw7JKsgAP1i0kj1g0jlzFI+0nLxtt
+pt1hUZg3a8aeKxkNwgYLDP9V9xGvez9PHAH1bPsJES/eT0FdRi4CkpzByKJRiK4
VBfn+ClJKd2ENMa1VIprnC1kncl/VdzPyhY+9FWef1KvhwnfVP4pYwbcMNZTQ6rR
FpjFVA10DQk0wbcKJ/XnfHE5n3vFx2vz7sH4wsGv2vJ8iuSsxGoHce0Fn8MofKbB
+OUVL3KkLQ2JOnt13Dciri9Z6SCeUMpSEvL/0P1xO7DBYLkYmaELcf6FwWRiJWdv
y0p1MsUyY6iG78VnuAK+mwFxFpIO7bncRXnTm37aoALtfcdwjMn+UnhoOmtJsT+N
sH9iePGb3y2eYR6WjFBzjZHm6TmJ7B+GODWa6XuPPEkiE9e+FTamQcw7lRxxAeVg
9EZNXsHw8xbGKXyCZVQBfNHXkFDynlfGRbKoHFDTma6Lxtb0m46P/+ta8V/e0Tjw
41Fe2nR7+6foF9b23UEZHSXEtBnQ0sEmJXNeDA6sUF2lwK7BhdAItyykMzDoay8+
Um7MMaWyrJkAQIVGUdEgxmIxOsleDrZQQGSTbDRGviwDHmnFHFrY9KRCnl/DFYsk
OEMHLs11Z71X7HpP41B4SjCtKzQDXDSsCvkkXs3qb8NKHqpGwb1/YX3pYpruRJRi
821SscSc7A8PuxyDAnskv5F9P7iGCQ/c3HJy5y9RLNH6IaIOpiokAhUawT8q4pFt
TKestf/twL9P7nyEpbrn6D/pzW32WAxOSzAurrcPOuU/evfKfZagNFOWNaC9vGj/
jxezi+qoib4EFFpLNTe91A==
`protect END_PROTECTED
