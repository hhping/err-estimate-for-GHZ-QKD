`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ab0Ahf2KlI7tfE8C1l4zS0KlTFYgyZfwjl9391x5OIZVgGpjO2bz2e68DMYcDbEJ
kC3J1IpVECCgAgV/e+1uCdPwJIfRvI6WM2BEP5LZQsEQz2oO9LcMRnMpXFRGNO4h
Hl0ZTv6HW9TnU0KC4QlHB+XHVzFg/73fGfE4Oeb/apYNTC12CsOqhsf6CqRYI7tf
v5CD5/Bjhz88KMBG8Xfxp2nb2Z7nlS7WaTZvUcKO8uKQysBKcm22GKRFng56L0OY
ZvJOrbQ3+Z1IXyVKf0eAJEXWgDQ4QIR22fhdIws1tbneqMOL745BLftbHy1ThQ3t
73n7HF/OFvqJrO2w8E9W0b9G+yaKd6cSZzfC+K5xDfMGXuAxxYXWRCtDn6njmL/x
dzx8WdgASb7TL/DHyupNIhMWh242Z56Ry/tld0uWYHEG1aDK3/i4RPqFp54TxLBr
QjRQfhkA1Ccg0njO6jSKpb2qI0y6K8Bl9bOffMocISmr/3J7xC7Br2UsC5Y1T8Ky
NhRESes5rZupj3IDU7YNc+/ZrC57r3J1DD75ZSxXAYxV4p/bqgzK8QxOxckMX04i
06Jl5vc/GlEc/g9LUI1f2chgWR450c4jbLK4Q7pTuvR3SoPdnedbZxFB2572aYBv
Ho8JJ25WCRtqr4ysTOzKwVBD7/gC8knhy55UbYj684Ojsu7sPNYdMNpJ1tsySuC7
1CXScwHmCP0TH8+cHi0vapOA5XE1m1cvKTSvZXmRN9nLJWiA3HsKfG0OWQZMN0lU
bk/MggCmIPetOduDijbuM88Goiia2zjTJ1fWJQisIEH/Y5Pbl78QxeKVSnNt0HJl
vz+J1B6y0Eb18lpVCJPOggstmSG6A+AiTTpKh++T77+2vr7Lt/6aB/shQgZ0TFQ3
bmipj5xDPkTeqSgAadGmKiRhjo18X3tLrrJ8RdJc+VTtaGmKDm8feapGE5dHB1rL
ZZEyuIQ2JbFQ7VXKpmIgWf9S2an9kFFLx4k5a1qt4W8LCqSC18bxJACzN6tC1YIG
x2EtMJLzsdP4V+Wmn1e+QdG5lUrzNwSTaLmVE8WAQT86sFoEXgM4c+vGP3+vA/+V
m3N1abV+ueqz+MCAgUAEjyuE2BB+sDT0rRDl0qlYr0zolkpLVan/PwL/nlqWltB0
oY0+V1LQbNT9DFiyi0fHlHulTCBQR0gJvOnNDoO2WI0fJ8FfKZLCguiYgNLGB42F
HrSouiskExz6xLCyy/G7pNwY21EyQdnh3alwffM9NyT0V86faUdHcM5cPsWTHc4u
1ESI4rgwPAI7z/TOYQtqVuLaQ2u1gz1QswYfojdL4YyVnk9QmFUehL/AnKCCPi44
yZWJDhPpGAgU9kh5reuH31/HWWjW0oDU6V/yaGYr+/ONz03Xex4cFtJN/iYpQT42
XDL5FmRkDOUeQc8WUjwM7YJrtt+yxxge+G7/2VNmy3DI3zFWdnGAKzNxtbpPXouo
TpgcIzf/dKMIwuSh1/Fo94/t3jG+zrsHku0s4qGORI+aCt44Fjso+KZPCmCtGDxv
iivMjCtIxyIA1Oyqeoh3+QYExROYRUtIGG4v54uOyX8/yLqFkMpnLe8JqdcOO31d
z8aE7A6K4KSz+PP0roJv/QN4uql1UYP8b72iYzTamSMbPgWvawAv976JpAlwsNtc
XXEoMfXgb8mR9cThH/Bf7rWDiP79VptyQ+l2KKGUGYY1O+wB3zJ2EnYhueZOohI3
1XCn3krcAJOYlinVTz9M0HTvaYIsfoFq+StgrJZQik/m3EQ+srIF1seh/C/T4DJj
k0bMqxwKvP4J7yz5xdiKfgVHbiMCdZ6CKXY40x+PLofemv5OP0cWNSHwG9rT5ubX
jeThRzcZyCnvqNA1Qk9B9CvczqjLFj6zt92/VwXUXBWcPtDleIn/ThAb+bNG3EVT
BCDr2YCysc0QCoH3Y5BIGTNgBV0SE/K3BDtlFA6IOTI=
`protect END_PROTECTED
