`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
46pj+DjA2Gq7564zqQbrXKJprs6fAvqtYzhJuCyAgaSEKALlx1vMnS4xdon2nlz8
oUHKx8QE2BG3ji0WnVdt3BtXwZdDAWBc1TVwlTusKF7m1HdjDcSnwF2Kbj6u9mng
RBIffShfWJv2j88j8afRjPwtr7LsUPDlzrmjt+itKu6mhIOrYJQwrrBlsGkSwyQ5
XCY0dpStc1CUmbJ4AuQVTBw40mxeT9S9yZrJV1+kfrjbAoV7jGxt8Z/c8WPTNoVJ
iYWkqpB0GJZLqeX7V6LwzHXi8mWLOmAE69BI4nsg5fIz92DJkfWwjSjhmqxH2tAu
lN79KUejoie/kjqP62ENiBwkOz5q64vG9aWycQt+8F2SlL30ofv+z0Dxx17V0O+d
ZOtTX9ts/Ykq/sllpSWIbOglhbjsOMKtqRQ1vZqHymWs1Z7jLsLq5/fhkVnjVHBi
z7+Jb2w0ibEk5meOZc7plN82uuDEJSn08buedsE1XQKEIDDotivyNNrhC5txWMN7
YUn1hB+pXhsUPEdKbi7trIXpAja2LOWyH/h3vjHgZZ2JL5hBmPwOYbuHPWZB+jK8
GJTypOau7jipsBkGgSwRfr6v0qUKp7t2PDIvD3OUMXgmYq10S6TBShunkZuj/+ki
gqRT8YHX651Fnugj2D7mSI/Zr7C+/TFxhZDkIXhUVQE4aEFIxs2SbrkKgwgAvx9G
YBpeC16HpR795wrzZiq1ps3r+yQYqvPxuQYIV3Gt9984LRmNnQGS+N6+MBJ1moNZ
pt8wbBssWLcG4HI4QfAabYYvcjofkqHPqNMvg5P+Cko8Gx88F7WcjEJx9FJ7+KUu
LgAS+ynp5WQUIyK+uR1eBiic+JQeKuVtHegi6OsUXnX4n58hPM0qvi0D4lvbxrHJ
mMLrQRIRDvUjSHdhRpmIaFF5/DvemlSGLJ6g6wmIppnduXDYC9A4z8Ede6QdQKBd
LB8q2N692AwiEKA5EZk5rcVE8Vt9W4AZh9pj7Na3ZJVwslgxuf0A1cGxy/XPO0Ho
1HbCL799Skih1/XxyNIhmGarqplqfgWOXRAPucWqoIdUuq+NNwkP+V2x9HSk5wIF
ow4Nqo2rkzUP3sSBnQBumoAN2EkgQB/HcTijhyZklZYwf7ONxCV/rqRm8Aa0yi9t
HLf+Wo1d5A7l0yLcSG7h7LZCrhYbr+1siVmMA7r9lTq8oxao6UI03aYbx28hOt1o
jO0aqL+4XjnFN2zIyfDHhOlwBzWOii50cg5xa5lK4q6MWcOgamB2ksffR4IGb9UE
2tHmVwtlw+J1wHo0caSuzmzqPaEqxjk/9WWEPTpLvdLh1mlI64hws8RYVUU5b97X
yx+aPyu/LtSNt8WFZ1UGAhpKs0oCErFq3HkJWk/mQHr0jjdus7XhHzo/plgFTfNj
GQRQeLdDma6hw5VGTeezB2s2Jm6RcuVqEyCn/gIvOmFaPcs7p9HOpMznH2GxBA6m
Smj5lcsOcHdBap9jujCVijnXtnVSU3EGpnXyNZwZZ57yOCCU6uOiRHF9cYl0UtAL
NXeUjiAXSTTj3eI8HEWp7VViFmz5TN1RAKJsU46MU0ZAdabkpvk/kyjnzjkedfNG
/nUPtusY6jbHtet968FvfX90pv9KR4oZ77q6fmXMwFHqH1ZODbTyyPuUpA3Uhsyf
gWRKzIywFyu2ram015yTH6Gj3lpUYcAZ9GwWjiiDla4bBDZqKzuaYB+NI2TOq9d3
G1wNbIDlqwfXZ96KjPRTI/+If6tH3eL6xZKb8IxazVzNTVTJS+Fr4eeGfsBKQoTk
GuYHen9qeoTtZvxFreQ2MevmYJMsvO92i4WDAfiSFK5RvWO3f5jR9uonTXcDq4pf
8mUcf83EaBpchS6LIGBnTveA61yF2vcPq0CKMr7a5O6ifmIkz0oB8Qn9e7xkHnpy
F2x4mNmxYZVtohzwWNpSZW9Ao2vBXr/LkeGJZfZs8s9l9lgJ0wcyFb6ZcFa2fbfI
bG14eZ8axEeaHBdUePcXRY4v0EKOeqDhjIF3mQOJ/0Sg2ftDcqnHr8xqxzpyDE9y
20nMORZZmCllZQie3+HxG2GdNH77+Xn7WL+sLlhDYQts5dd3d/3hMBK8uIB8a3LR
evlOm1NFjFJFW0Kq7R7rq1+U9XRjCMR4lozm4ou0RLn19nnUTUQ/etTwZnKlJaab
IzJF0cJ986pe4Vziu6SPah5MdVV3wmPi2UnCdMWItH2+rdKTDGYDTbTmQUddGTiZ
2VwrXTrrC+ESlkGWKXP0bhCvjRkeR2S+ikgXYGG0e+Ek3tNQ12no8ck+jrGIjA0L
kD/qFyANiG6XlwM2vFi/8n2Ctbwbpw+8ixm2PW+T8MAifO3fMrmq13YtnQhoyNLn
dVhGZZDxmGePsfdVexGUG4ZUEkqnLkhm1vt+cNo04b5H+S/vLSzwbNKZmGZa9ceD
ovIQJ65VAH/fh8qTY0t6/bQGrQG5BGvad2/RXANydwBWVaFBOc0Uqzl04FjVNVMv
GfOzhUpL+3EtSyUwAOKzwT1VNgyIc3kJT8IqJIjgc6LY/i5TWAvzmvv1xmAuItec
bhhu1Ukwzs8v2uH3vjp9fA7Gmq09e1dnx0q5vz2ZVCaEmRc9J3Ov78N9CLkVm71Q
VkIYKo7dlQjBs0WoyS4WfiStv07Z3Wnd7vr6eBH72B6CczdQXT1v5O5J5tm7NfW9
R78IIakRLsRO/vA8Qy7zZhLIhHPQ9WS3wUf5LWSVWGAawGRbg5eQSKbvBlRH9+WK
zwVAJ4GqzTV8vEi+jbKFMLlDAtVzntJp3perQf/nIlNm/vnJ1BEDCERmV7N3NEeg
RTftNIebazk3zEk6jdhmsfetTivRaWyVlUBsALZ5oJJcNFkW5uEq1TtYifUQidli
M4LtnzVtYw/cW3sRvRkXxhPbqAwqrWQUmHGHJyA1k701K7b81pYtOLrVby+n1jS6
NvcRWUo4fRtlBLPct2tj4Vc0GqyGuESxCJ0VeXAlDNhX0s7NjP8UBRRH08LeXq+p
BGuEaVNZaZBUH7WLMYrUSO4IUoPwG9qWiF2WziPHaqlVVzEsT2f91/QztQMRcns9
1Kcct7HP1H+RgWqDrh/K/Vs0nuhKyRsPk332LWaXIPQxKnBLZbEkOXU5Bz5pY6YR
AS/ca1OFDKFMX6TWA6Oc5f/gbpKydqDNaDlF/RLprNgNmJ/084FKa+pgiuwTFVuP
UwUcpE9ng6ikjjglSvJdNVRQe0QIy2LX70Vcp5a5GifQ8zAjQDLwwn3MR2y0tzy3
s0VHj/U3NlKMwuI2FPl/33QagRePLHqBv1G97SAhznuJqR14czlFvX0wf4OHpKjr
rfM8S9/tSdGdvF5vKE72boD2WTDiu3bFBTlZC/SF4ewM6wCTMkC5Rqu/nHNq1oTj
keD01QDEE0TOTFWD43ObC1XW+puteF+DIFc23mjV8NOvRKRJn9GlEakId92WaHpx
kZEFyAWZe+YNl1+OuC7gDG6hSVdk16KnzxhRITu6/erFQUmBmLkY2gCrr05ePoy9
1GvivyMsIfgyziyqwwMFcSVGUWhyhNY41NAjsuBjnQK6YewAQmvwxlcwYf1J6C55
T1TfblGyscuphSHFRxz3UXDbx770DG+zMYsYN7jpqwe2jm+1kZmo6XHN0JG/M+of
wF47KsOe7TKsISo+D5X/YfQnaR6zrvP6pOL3pFZzHSLnBtmMcyCCq9/2676g9eU0
kfs5VALKLqg9ARt8xGTqjbSYgG64ahBCcS6EWtfCWb3VoTv3s7ZbzIOvDmwyuyKs
ZOAa6n0TC61Hnb3COtEK1PwGiHt59SFJDq5VQXbLX5DVNq9NrGwvp4MDnlOarPx6
i6S7Q/w2ZLcwd5YU6z6XupqAgI34Al/AEBPH8u4KY8vsgx6rw8m+hfp8XP/t5Uyk
NCW2izPWA7on75AUiYdXKlbOWgmkw+uJg7J35srTWlqGCvk6s1tTbeTdzMIu8HLT
dhBiR9GH9DQNPHNICdY8wqIV7JZypLVEJC1jk5oMxq2Uvkj3gsEmCeM4mDPyVQyt
B8JoJR54Ud8nO+3aNoec3wKaA1N+FnsQPHDlKcLRvZWuSVKDiyrM/lBW6K0ZqcN/
60wgX//U/QluSmdRALJRHBFT2K2QEJG68bweGBtiraqVvQuxmUboRwm6jLhmQ929
s1It63i4tgeDd+ah8wmcSU7Oa9WpvDL9VNlxRvMMZtR7B6TEyBM6PExm+WqkXt/v
tmyZLSIjyURf1ZOpWxaVBDKQCx2ZzYZs6lSA3+4c9Nh+OEVEPAGdpIJ7tuSFOa/4
odkuK4SSSkLaXID95g8BINhw0PIVuWENba/IlXH/EgRRHiHXTAXP9N78aHDB+zWS
yuIqK+iqK2CT9JLCtYF0O6VcqDPjI/PNgFRYZedr2HddqqL0or16WhdoxCQfqHhl
uTD4y3WSr4f+L4PY1TCbJwiSM2AF8xboR5F5vwLpHZNWDwNjAwnDdTouTfkEdBrW
xDqKUC9F20JyoPCVYqachBzEukBHSPNhM4O1KUSuJIkYCuw/sXodHFiPF4fUKxuD
hhZPYdvxW59hAVD0l87OD7MZdiTRNafEKkWmB4P/Z4PGf1KK2rbsdWSbx0Yf49ni
4b7JOKig9cR+27PonYqW5bjVkh6UxAmCR5CBjQxLs0yufMPdc+QHGIlRxu7dFhPX
bciPDxf4K2QXL2ihrJ1XVg0FqfTmsnA8d+xeU/sbSGuvsGs2TnEIKV2zv8fP6RHR
L8ytY0dfT0GpWY9d9ZIRAGuIKNeUuhKenVw2g4DNWbz0ffQTC+46GvQRhjrB0M+t
qji+4XDvh4gr0zkAG81EHIoc1IUSEJ/Jx3i3pl5D4w0iBM2CP/gAdTeBTqRq721/
M8OvrZKW21jvn/Xz0T3l44X1aB0tDZ5o+G3d50NB9ZpmDVXoFJCpVaXnOTZ4lxBV
ZFpKjNFwt55p4TFLU26KwMvxuzb1WPD3nXTzxzOk9jk0hAxg7qzmK8d5NnNk4HZ6
y+ZatSuHDtxSse4aJ0C8XhF0Dpyw1CTzvJ8QRH/IPl0HWoP9ujzGYIwG6wvvGcc/
6PGg9FhARUy1MEF/OmjZd5CLw+tQVxML/sLQpGeWuiyaFQXzyGj31ioo7POxN0oz
dPEpLz4TzWnB3LIk7uBU6xwbwufheHf1FSFtNCrgkOiFiNzVhkZp16GfBvRDkXUN
Xq3XGC8s3Gvo0szhV8fuN1jLDk6GiVQVoB/Wgqoeoo7rWkWgDdH7N/nKSADXC/FY
l6DqM3gT5e73IJPitRdeaVCUQFPwrU/hpPsq83spwlR2DvPl6VZ4oCRnPMUULW9G
M9Qq2CWO4vFw2PuEU6oiCK5Y3z374lXP2rnsp4/GOYkYMRmZO6XgszYv0BtaafzA
/tmTL2hYVcar+eRmTgcoMK9r+SXi+OiVVVNbaS7nu5jLVu2Z8i2TI6/ZB7nbbtiE
fGBS/d7BBdlnoblLkla/FrUgeLARYFXX197+CleOwy0AWB7ULmWeJFd0PemMUN2c
o/txdDmKmsk1fAHb9L3ASgDtEVY7MF+NzTJwtIpKyj9Ez7HoK0ej9J6VDK33B81F
tUpDos8BspHBDsNDKiVOfprlpOV2jMNy2cGUKeOqevw8gcfXj/aSn9i6ROz5tjzZ
ktiuVrzp1bC0RCirR51FV7N1DGyYAiwDg/ftX3nh76j19PBZ05A01IJKh1JJ1kbR
Qff769R6F8bYizv+mSheBghl2bS2Q9PubhjeApznWDR27qK2VGxg6StNH/zmZ2U3
En3F+kWx0B1iD1R5kheSTmKzxN3IIPLg7nVdMxjIf4j17rPaHdBdFtsDB3j016U1
T/8CGetNQghsjRXOUMh0DwfKWMcM9yTUH/GXIUJJcHAaPQSLYfY8J443eiKTvg0Z
u1iN1moJfVWHVDgEMdgDeRypKpK5b0eV1mGi4Rb/xnM1XQRAKs1p5MfwDpphy0st
FUtPQFDEG7QlsmoqIv3TpGJjAKpgwejoo0SADUyf4ZgpkPzS3Ja0BQMTLcU0ls9C
eekZ3e1jNPf+AQlVGwSCCBElsOUWsRCekndaKQjtmbAff0ZRwHptGVp0XemaIbk1
KjvBtF9WfAObOr7n7Z4jzfBckZPXI6uzIrI7wl3MURgTArads65Jr+SV1u2VCIx+
yeGVDgtrejBNoQgK2br/akWMIsQVrbbOMxdWfLLlVDxciVK+Hith5iNAMa3Lwl3L
yuJjH2DuNftn1DGvwP2sKvsQV/Pa8UsfW9empvzIWTcrrEXdUuwKcGI1IszCXiU4
LhkMHE/peyUoFb5Epr5pYYFI2Vj/AIk9t5F6daSlKHQSQreQNpITzcvShygHLbqI
hrUbanmyp9iGUMbHoGvy2SK02SRkCDdW8qzf/aW24dUfLPxnGBQiRAlhnvpdXd/v
rTNDY2OUpveROjYGkcpnVcoH1oQ8D8sZ80psbG0hAeCy9TTu/ewHGFmsFHWAsAF2
ns/jQr03JHY4lbjieXS7AJ0MJWnU3iKhWOg3smgZsQYy5h+Rcf2v6XgW34WXKi/z
tuqn7hJgiepp5X407a0o8FqhJc3fZ9m+g5J7h+sz3BOgJanZxVvXrVQJ5K0/OcaB
ddjADPS5ohuBJieq8K3Tbb/wqRMOjwiFX/OhgiplIjHYaYzq3vXBrnAfXbPOiqz3
CFOQXqSx+Zm6Mb3BSyW9Eff9+QSt8xzWKuIMdST/XLXRWcPaZ1pyz2oFKlUuVaZJ
MWXVo1lG8Pqt1KrQoBC8qa/x84hjNpvkLUfnWm6rYLQAMU1NWqcvOTh+WvkfdNjK
HMasGfEtQzMRRUD1aUoLEjAUNWV2EkE6AhDp+lJTn40LEQ0q0oQE/LeiGigcLq3T
Y0Jx5/skgk4JEVCMGrV3RBvcsZe+znD00Cu1aM4qZk0cG1XS9s73bmY4FcmbI1yS
uJf44dLEdFNFFDAoQSZ36/L1bJoXVWonz3Z2zeHh0OSDnHZJbVTjp5F0D7XMy4JF
/+qI3MmIsgq9epBfiGKwfCNa4tuIG1C+kmfYTmDv9ko3OOFE2p16045BwJ1XJwDY
GpPaBU1YT760nPR/rMBlFHOjStdZXzrVrd+KVDVooQpgYIBTKQjwhaExwqZrEfM8
6+e78ou4MjTKMiQyLgoyxHz+ECYD045Jc+v6BYJQdn6mPYMLOwj0PvzWhTqb0Mfe
nv1y0RmuycjaxHgiYqmnZNt19cpq25a38xlzdMJu/m5VAPezYAgAOZ/HT9f9pyYs
TGiCRQb+c6X0Hv0KflgJMhyMs2gizmtfjf0/T7pBD4wq5aPha2S1+jUJM58ycl8L
tC/fri3Te/sUhGOhYcbJyz+mb3lBybhecRNnh/0wYLzNvHK26LhDzNDu68MIMbM8
XBj9QrJnuJevixQ6Lq6DZrr5dbtYlrEzj0nWZqKcx5n/8Kp/scdm+hhLRmvbnx2v
S/aWdY+JPr5kh5ijJh0niepJXCNZ1duNfcAFxYbcaBaTPa9uEnEqGzVQ3mgn30ka
BA73vn91ug3Pix5efLAHjcJOz6EVtAe81Q6rfIlo7oH28Yd+stUvTMBcVqTgTpDH
0ESIUf4vu1/maOu2s/hU6T5ZOVtgjt0/H7PEeqSZ5D0lAIRhbV+WVoboffGgHCiI
4c97FnX225iPVTX+OD5859imk7CVEaUeTenK2q94FNmXl+of0Dbv4q90zX+gRC3B
pfiUK1wYGwphwQVnvEvWrrEubbtv0/Op4haLs1V8Iw/Ow64fZnx55XZLZZl20AgA
XM/2srWe7yOwFraNkUS0frKYrt6EcOqbkhH+X3k87IaezAT71Qn24/Hx1tvMjNu7
sgcr1AeSzDHvedMDlx5lysBW6KVGtJpIhFjxknnTRLsADgGwypP++3CI7dnhSZ2Z
V5QcYeji6Uy+BVjJl8E6n97EoJAe7YNcjxvE/XkibpF+cYhM3G5LtILmVkkXxJkY
hcUd9cBCqPGYdVdXimcnkHS4crnKHI2r6XUe/zIR2siR3L9EQ9GEX8wWaVvRlFN8
stwJNN+gHe0lVAW3hyYdQAabSiurFZgs88uO2ya971kC7/X7Da2Hfxr8VuZgO5y1
omdA4JCdbAAug6kFenMj+aHjP41YxuL3XpnBFR+Mb0bg3tDCs52Zq/GA0/Vcn1lX
l34fvz6OBao2XkwQeTe7YToqeJIf3CL8VkIuvK2uFXHoHDTwEv4pAHOhIaGb4ICI
6wNv/hUqOfAXqir4Sj/PjtbSQbu2ImRZzDSrv5RwLCLhbBFNVcXw1xaTxHKWnkPD
/fhTUx5vpUFrVKVxt2WXwDiwkHusAQQ0/WOYo9beoBarUtHttQXE25bbwvNuLOAk
O7ZMPBemmBCjKEuVf7c8NqkklrBXEo917te8k3i4dL0M2JT/pGCdKtTXt/R/2wpV
x8Yk7aJ7rSFMC475u+IlTdlPaQC/euOkufqpzkA8U1a6h4RUxXQFOpEBLZeJHkzv
45/P9kqSBBIAmF1xkj3IADDhSFjww/PFdOc2k89kvNLw6Fe5OZYIlgMw8AI7wpnU
PGr0Q1VrHTMRC082OdQ9ijaeOc7aezekyBp3H50zE91thQ6vYBDf4M1lDb3NAjzk
T3krvFpG6Wa99ogIYn6aNORKDy/zMpt5syThItzn2T8N4azZppk5hPJKtdG6yc8O
CQRPTQDgwOqVPrWc8dvpBo5BuXTzCEEkHXh0Gc9Do22VwJPqfBstGmjhI1wn0fGI
4p6K1UX3oN8BT1fHmrVPcMjMuPwRidsvIBd1nT9JvsHRjKu/uGjyCWd4/fPVGVQE
k4z6+C7qOjd9F8Q549L9f7ZoLMl/TgU6Hkg3WIEVZisRgS4ozc7CtqV0tkS4A6Qk
Qrr3fL446MMlNHUiSCDvVQ+AElnRt4Y9SJ5iY0FbkP3Bco6dnA51SXSBmPVHgNXT
3xHPjHT36fUQHpPwm4Qu5rlOfJbIDdPl0kbRhlewz8e3nfMxj+oYngUchLpa6Oza
Ghscv0ENZBgcyQoQIgocFpyGVUdnzidx6Qlm4ovzCAbDJ7834xBwGKnnQlVDWQad
CFKHUEXKjqLxSXCJP7rM/OvVpGHAXwaYCnvn5rTmshdmXAv124x7Kg8kKvNQ5kaP
uECWzLJWrp9HaYoTcF34v58EI9aNoo8faPhkRF3L5PSRbdhuxBOxn52QwixwgW9M
MJSLQ4w7aFIPz4/+PoTdxUiSdZSXsW2QXXUC8SqPfKpljoAuwppiHAfJtbJeEjrv
2et6smQ9LL7jH2pyhfP6hgOVeyupImW4B76cWwU1RD1mdgyjxRnkTWEq1/TEQ+kX
nOAsfIAyhaygj8DrSJrcvpBL8i5qM54AHod97DtM1COzHupobwQA1JfrUD+trx8H
hc9889BPvtk1cSMJnTP8PdHBz99P6Q5TmKWwwETK67SIulLT84MUV7C+hdq40J59
9+CA0Qz0WLOwBYmLzX+wvxYOEokrZ9nclARU5XXgxhmkfuvhzMFXxxgss3kay6WX
vmo1ijTolOGo4cXLhjFujA7Cb6p4V3D0vmJ+2PtYZtiN4T7ZBfMbIg6792zlDaiN
AUCwrafRe1FUG2apulWXNz5pmcN0ZUC9kTvhQ4+OWgzmoCPNmEwuOSbw6erKYAH+
1hzzeOBtvltMcNYcB1OghaeNvAWmaNTmgVJTgUO3O4noQVwydsBqYHbClB8f2iaE
uwqTN+XuK7pQs65PD7boMcaDld2kjo8sYPUyjWP5QEFtT/QOweYoSx4JGGc58SAC
LwnloQta0pWMGktiau8aOCz1tKTJKvak7zMej3chEAHxvZ8vaR5CYHiR6hzEr4wl
Wy6tKOY6vzoy43QrjrMY0ePIMYKKet1zqQi7Kdq3AeZ2xTmNxOxsRa9ZLBRLtqCK
bpOnuMegPLCjWJS3NBAzN1TD55g7GXkTfMMo6RFJfbxboWV5dVVSJmOoDIlAZvJh
WYl8PI6TMiJWZbs0AWMHvzJf46Gptv/n1p/oTTlfL9GFbED71QLFzVgy2LQQrots
Uj3mQeQDiJr3dW7qrYi6U/47A9/PyTnPzUbddP5S6OVHOeyQmLykJVtEJjLgRPS9
AUQ1+yM5k3mATbID5tdGNv6tFa8gPiHJ8J8uL2/+G6PpTCcESNRIZx2IJedVHQGq
E3G+uaKETZfiyy/JSsUsJYh29Ak8SYjoE2+n8lopDmDao1Gtem9CADDnl9EjM6uY
HzqVtJ86tZZGqQk/h8Rqa4/x7fqKaJdsCIOWi/iLo4qr1JcU2IQwejsuKNjxdAVg
Pi/q1kAU3oEf2AsYYqkUmLGOhXneoszpRhSadFiyRukmDee7jGFZhK4N2IfpWMZ+
OyEIypBfnP8m8V/V1gpT+U7EoHetc/eUTjxiZ73Ld8ilX/A7kP4A28UZU3qLAoV0
3SBHV1BzGYuyKN/EWLMq7N8r3+qWjGpypM6vr7raDh7iPkd6CiJ2EP8XJdFaPS3j
+ZNdlenJeHUMulJ3NkzL+fmfe1Ioj+c7ezK2wbHjam4NL/ZZA4CQFenWJ+RkHELt
cHq5Bx0FyPpiclhxSp7HzL9ihjkfyeT7OCEU+teuQpLIUdGyOCQN2ypTVBkhA0zg
Q9p2fI347p1L0rj8E25gF8+qV37UGPhP5S9z+UKKynUOFkhN+zMioymvLOoIqlv2
EESBAxtvoksFWQ65QAEZpec2KVSrlZjEMlqGfnMyjCqTZyU6oUlO7xccPc8JlR7W
V4NwEayEBSZNnkyjPTtIA0SPv2iJYgi9mS2nkDabyEWnx0ktD7e3IoB1Bxh+EsKO
5egd8cE5QwPkTGyIDdpwggs7ntmFuI8LJYniTi0IkdjhTB68RiIoaOUHstZb9k8s
gLiGpGX0m7x7U15iXVJUQUq9KcbXZfuD+V4VDD0QfGBWu9dcC+QyFwq1D9eegMyg
Kxpg9CSrj9l/KBL7UVpDj58mOLGlOd+hell0a1S6KDgCi70FA8HEuusTmU2EAbPo
RR2O4+MrRM/NraszF4474XvNrY684spneG3UZ9YbNqPomBtnKa+OG5CYuKmOQ3iD
W/vNMpgz/+Ac1xCkhd2bPTIMhFWLff9UJnR0cJWeljj5C9uM0WhvLExGqkNCZ6KD
RsEOCxCRhMo/98Y2tNggbir2UkO9WdTLD0yQYiAgcu5iq5aKtKdqzt3IZ8fTNGLs
83dtudWfszk74cwt0lETz1NU+K/QPrdPxRn3lnkLdXhX7F5njnTTu2jps0FuO2B/
Y8ArBtFoQXxsTh+oYlJzkvEHzpjKSlSx7va/zWQAVH+RebeItJjyFGw4s4KIh7Z7
m3Tnzsw+UsC/qTnDigoPdlCQqtedDAv9sa7GMftEZXoNtjWfFBitHJUHUKPpZrbZ
66HFsCIL4AQGTDSgGsrTyUXGiqbF6TCwo/vYF2GfIMvY7u9YqXAfsv3CsAcDW5Xy
Wcs/qklDFV69VQl1C++2PtDdbn0ER3EyDeHf+goKss+8tv1NTLrzzjEg5NvfxhBK
fixVrlNJUwOG+RvUFoV1qq6mHuUwZSQB05eV/moiA/0h3Sou8G8kdy3QkXTRKB5t
mKNRLqTuOjqMw8l9k2YMez/ganvnfrdQUsaed49gMJS71/OTlqk2SXTSf1h31kRo
j65cozNWYSOmeihahpFEuICceJYypBmSY2q4IlZDQY6pXmHlTurz3Eqhef0iOcC7
iE+pL8xToZBtlqdwHzfgNqJ1Yw/yNrPSOp5PjY1hX8oDWAuLjpr5z+0qYLLPwvLB
Ysc+JOrhN+1xCTzF/1W8WM67+3ZfRfVedt/gj/SmauR1+TVJFcjLcdS6VzpQiVuJ
T5241LN4yCnu7IozMpdujcNqkPC1GwvsVo9Rx4DqN4VWuMKqlGm7a+0zGwK8eC66
moOMaXu2LSIWB8hiOK5uBbH07I7U5IMMeE2WJC3+1ErV8zVhPuxYVX1QC1fE7kOo
XWcbtH5Qz01YtXg9Jl/88Gp40HNdXtw07qlQOHDZybXkcwVJEESOTKJb06BeRwef
NHyLEzT7a2g/f7+uOvl2IJy/RnQf2Ax/9SNtbhpVL1U7z8k7NOcDnGnn2UYX1rp+
tWag1fD8QhmUpWKbY2wTgTuHqlDqU1SWRbg8oF8vvpZ3xBHDUice72kvwFxbyEEj
a2N4GgYxj832TSjIlUiSouogduJC1HfGtTdacq/xdjrtT/S/zKRlgFye5xo+pBVz
2JZAcQZbFqeIe97ggMclHXlJvfTEu4OU5Xe1oSj44qi1Vc98XYl1lksWyBbcVyXk
iFBNNsV2d/O7aVLQiuDyJGRbaUvAtR+N8mnUkmP9m/hUd36R+pgfcf1y8c8WvPRM
G3pf25Cxk0CootVEK8hAZwVx9adrOWfGJh0xkY8qFKSg+WDVJ//CDXkyv+yXVFkF
ViNplJLfiiu5Sbb48Y93OddiusLGsr2k5ekgIW/yuul391OvBb7tLqyx6oUz/tEc
ooqop8VgsFKYgJ9hpEoC123IUoHWvGrWwHECUhuMly9mlG4A+z7xJ7vIk1I+KIzD
xu5zEt7aOrRDf1P+g05FCZaSttkJG7Ojmr4pv7263l8rstg4AiFUa1sCjAjll7kH
rW/BEaYYmqRQTGB2dstihU1ZlIWMyCQFwRVBoTAg7fmwiz+4rJredAXxrcjpDwkt
bewaRsTO/Msj9MATV9mLPyoKgjz4xqHFbvGzmZBNaIRwJuB/CpB17MP/xDnLNGYx
AvdHZ+mjC70170mTUL7cc9kPG7hATxRwaTBCW9zwYcZEWD4gVLvPqzZavGd8NNQX
WVgHoQ6GxuvteAXC4P9xg+XdVCv2asbDkR5bF53ss6NkT66xZPGgf37mClEtrQzF
KFhaPr+LtWWaOF/f974O1LPpl6WRdwzMhMgfIhqngHO/HF83kh/UD9s3QVw3VpN4
fWULbb81W3PTkQGo67XBUp/wfGi6t+Mz1wBJ7J6yHbwfw+tOiiDDf5z9WnrJWwHB
Ev06l2wdu1Es0OBUFt0E4YN/KKJUnnxLqzJ8ef3w4J9VC4vwTG68w/BryL7HOgnB
rnpTJ+OpR3VpDERu1+/hstpxTREul1HXpfs3+KaHWrFnwlKjjsEa6CLy3Hbyv7rc
y672fTWPf49eavUz6ETFqx5nC2JQc9d/Wv3v/B/wDtw8V6Y6pDhwnPmu41qhvKwa
F9zJsbip1gnyaEuUHZP98rRXwrdrC1NylORd5Yk5c3U2Ipz1pKTfk5/HFDVlJq9B
1K74cVXUjAOBLllH5/AQVRTlXCFWN4v9gy+cVguldmOVgvP3AQBmcI5Ow2ZnvMm5
+I7wLFvOnAd2E5niUpl2E3uTLS7ilUGp5JcDPsXwJB65rrCe5gK/muo8VZwf8UjT
runr9WQ5XuAFj11+dsBpyoTFlujycGdWRwAw+B2+bY0yaQYUsgzpo45OEbPeBnSo
AsBxwfrc8Hc+1rs0UEF3A2PxaLwiIFA+XgGt4lMIEwV+WYR75YGUK2zmN5IUxuUH
dbVe6MF3ObLRs6lQD7tnjGjGyk4+prRp2BgILAi0hH7HMHUsLL22mFB5DF8+e5Ql
0rIYkFqPDd1bjyGk12QwmiHqYXKify9Xjvv00+xhZQnjseprIRE4KYGHIM7a5zrO
LbceBuV4T2Gxv1SHRWl/PIf+m/KYvzfkOW2eEvJ0vFoKhk1Ufq3J40lwm5fHb/lx
qOpgXskm1E5NiG2akVpA8KpHQZTTEQe/LqujtBqyQ21qGaX+6SFqoPR0nMHZmzdC
BGH04+2oHGFhL5BDZFeXm2+XjqhlKXwJbtmcrZ48AAfu4mk15cQYs0MZeU6IzJTy
+BCCYgiDWfWAsTU928QOXUv0SyFtUK545+LmYuIHMYjeOq8EPC3wkxYis6bUlkdl
wE5buva/JO1YlZ8MbRoPW3iFQRlTWiP/+E8S6I3uIVDhVCKSkEvX1s2IimQVwoyC
6riKCmRTlVbIaw1YuODXAa5ylBwA1hlmyAYsTUaxQcxxg0GdnDS6mMVAzq+sFJ1y
4A531uV//dVvOIYJUVzH3e+3NwsYdGzEtQ/xW53NkKF0Z7VRsAIuwHZx3ouMrxFv
AD5pfNIw6dLr+qDvCi+Boil/+gPR8hiCfJ/xSMIIX9z1Rh/dCAAgiPV1f7UE/Hfr
IQCPHhV7fz9mYXiDAHR1LwUfRzzenxnsCIUEvWrk03enITzlRl7w/uPqTmpTPplU
qI4bZ5DWCY4myx1ElJcsKM/5y8jR9H5yo+5v7wl4811x3AV7qT/A76JZ23gfuG0d
0a+H2lKiBOQDZn0Y75CYzwNO9/je6CTQzmhcsdIH8/At8gzcpFeBQXWTBW8wTnK2
UA8zIOV1BiOxR1Sa6p7V1LjpKMm+HUMlPlRNKUCp/CN0M2iiw/2/fevFlunzmAP8
SBe5G8Zid8CcG8QNr0BnnikmwhLlCASNMHD4mU9ZkohZ8/YD99GwGY0U1ZjFWclR
HlPHJSBNu49u5Wz5JSjr8xkOlfNjKkSZBoMRdN48+4i+MggkcgW+zAFIyzIjvoKa
PTAo3wBvCs+f8ggBhaZRlm7nq6sEJNN74HIrwWx+C5YBE5X+8R3c1EC3I8fuBjtO
OtC9gLoJ95kZFbOpcsBKDFRpAzInSH3wfFzk5MXRMsAj3+Zme0S24c2svDx14Tih
o4IID+40UuV6wDEJcU+gEXq0r6sj7th4Z6BjnTvJIsRrelf/OxIQfSaxnjg9yMvi
6Y/+2inaCejS2kb42snO76NAlWIseBjv4KiCc7lVNYKwLeoJy9aLKyHGSR/pPO2B
FjRECvq7EtlEC/inPhj0JjZWVKpAN7l1DoIfBARXYuGByjuv3GJImriH0OXtU3pd
ALCyjKdPmS1bmPwOBC3l28Jr0G/O6/S8plw/SVUXFGRNFOgztGzYUe9z8O0KW5sU
50oZly7b0qAr71nZK9lKfOaI9HMKZGI8qPQdN3ynt0VU33WiJkB+vsgdc6XWd45H
cI83+GBur+YU9pvQLkkvoOr4fYfo/AwNIMtcQ0rxLhtasS9468YL5vQAsRgPhaO+
GCUjAxIgI7lBq1SYMkz2oIRgx6K8GrYAdIKduDyAYKLuMqqEcZgC5xZqAUQBmY0h
Ha7rjq3MLkzJTBOwEjK1KA6ZsUhLQODHGWiyH2LXzygfMNx60lHxNilogAxnw9S3
ERyJuJHZQBO53X6c41q4d/R8YD5pYb+HLb4CHt19ciCmUpqHLw6BG+Ea3VU0DZIL
Mw59NGiPonqGCxC2w1DT8EZF1ercelc8ltUiU6ML+RfHMLAulFEcJh2gKOwF2fjg
vNWpyxaacJ5qE67xCWoagqyEr6vss/8o0qClSC9gjPJ6Tw9InuqiKPj2JggkVZ8O
moflrhOYpWZb8hzndwNOCVLZLTVEEkBaNUic8GT7t+qxyu4If0JiWKRZQqGWFv3E
h2qt96m8N2jiCUsPZ1qX1ydy4VyVrGsY+Q2WjeEH9HuWwxNZfqbNtrUdJuiPcl2I
Iqsh7J0OwwKGSAgD5J7RYBU+PTZMhPyfZWvd4ieg81X0aRDWKwAoUcaLC5lV9TO/
n2BUylcmSQEIAwhEg37fwZ49PYcfT+ZAoZAFp+lnN0nne3/TfVcbdQweYN1BHbeO
VWsOZinIjTLKogDYEDn8ZyU0cL4Kr9FWEhsxgcYDy9prK3AG/sdz8eu3bNV2zWU+
GIO9L7Avl11JgU0lJ4shC3FvwJzrLzuomHFlBmRoJiMVFR++66ox0QxyIn4c76Bo
sKKKuLQNptlWPiWzu8ophUhzvBEqXHu2BjZSrp4ZB9kHnqYATQ0hEnIS+B7t0c7G
HNn6dp9QGcm/tapqHcsZbXN4NGZSVtwoj6Kbk6t9GuRia4/2H/zdOkzCdkzjmmbg
/Y/6r/BV/wgBKsIHZyiIWp0fQ6GNx9ut0Q7SRfmX358t9NCz+hcYb59mSOtG2AoD
IeJjeWzzdVwgjWP9oTCVqdJMnfh/P2fFpmoaH3Q+huJBtKH6P7uBauMyF4jb0L8h
7QgApglXVpX0q3ArDS6sTL6yMl0VPTwEcFkYiRZAv4R3c/VKsJYR14hcMyMSP3pz
EyrJkTQSsyBrYvFyeRoaIMXs7IRecjskqbC16XmlH3HvPtQKfVG5guOace/yhsO1
AtEDjQvU5DZENnMjnniMeC5XMfZdX6kgw2ntUPyDhhNz9nUUBa8PFBuEf4wU0q+I
KLQ5lmX1PaE23mCwRR271+zCvGvNRgiYFvUkPfuwUmUDeoO7eAtL65OWL6MMEdLK
oeyGDHB+uhBjkHxuxVMU19v/ZPjIWh5pzGvLW0NJ/6tPGPIOV+D43NoNGSeExsSO
ri22JDm32Evahek11n59vcbbOynxsHx8eb1U5af3uPieme7YqzJT+dijpJINoL4W
7tZ7kWURKbu68KIgvk3vcztT+y5XKJNmE4KlqLKEWtdy/U+dCvsTCadC5EnQc2lX
c5zAnn3BQw6Zpt8CtJwu1TkgdQo+bx6djRD/7wby5gynN+Lx63EGTqKNRY+9WV+H
oILbc0qczqE3Gg9BmiYIw8NBKUwucoXXY5Nc5UZXz/WObURd4wWJrM7RdLaJ/fLH
bSdJmRcJR9oVEB8RIDOs1L0gXE9zQB1iSagrzzz7KRdojkTez9c6hbHuxglpZlqK
w+oUHafn7aAD3tDt7gWNN6mUtsiJdUsPCQTr8yAUaINa9zw95ggoK2/sbQpQe4kD
xD010FNfYUuFsx5MpQZruzm3K2nA4H2276nMZety3qG8aPlQTXW7Kj/HoOItdkdx
05kmr7rpPTmpDttsn53Yp16yzKhWoKIGXiBP4IgDTEn5avpy7bGBZrwJop3fVgG7
7kPpQzbYX9IJArERbQVPrnmEsiQdMHhXHmheQJquGR0ELiaZY/1qClz4PptAzDXu
lQmp/NKJLbZn17lrT4wnt9gdOKiApjo70UogpAG1QlKc3wmn0dm7b+6lSkrlGbRy
YZ9hGV1Eu4x6Zubvbnx/b11JZ4RJMU1FR9eEf/Gmr8kRIRLwONc3Bz4q4dEtPIBT
J6NLssDHzu/OzCZasJlR0v5II2pBeXtn/uTsOPpzJ30F241FAAf4Xw3Qy3pbqaGN
P3mRIUHgUVYaSOCFMuyskNY2jwb1aDfhGIpsspoRghcUNGrkPY4oKUcZcSFZRtoj
TIx0UJIZEqhkd4Z0eQBeKaRxfq84rdhotUQfN+8wYeT6V2W222lfZ2+fm3WzAnO0
h690dm5fsmgMF7ahTfLgoLDNCH6l80m3u4ioYAggWMp9VlqRQdL5Qa7hw7giychk
6Q518PjEfwHBQ74tcgddyvuJpmlve1l0Ne4/nCpNzdvZN3+Fx19PhA6vE1HZIQNq
Sc8nokcKDZMY5ngPS3FZIsATaKC4M6t+K9dX/Pe8le7WhuUxAR0BreaB/EwZ7Au8
lL65aTP9wPJ+BYeMlGyvl6z1sWVjn7tPnauwheRn/L84eFQiLGBPPab34dNZ8rih
9S/Q6TFtpwxjnNfAruSd6GesLcARz6XnHSs8tCKxr4pzh0dLdaP+taGzRTK/caNx
NTIp14Ssere8U5WTZfXYNi/sFP6seUmfEx1x8M5ooRdaBFUSuSLzbXlJb+9oeXHJ
iZOJsdTeTf9/hxQVqqbaWfacNQaBVTQnVuEKmzo7d3kp2cgQixYNT5MTmBLedeqt
1ON8brZhcDhnmiQFektfHMQkfULQGUassyHRY51YgR00lHWvLyrZki0wPAaceCV5
FFyZmWEtkD+G/OH7ZBgBP/5Q2ZBnPULF0wMZQLVemK4pCIs2ledgp6jMj+DugQ3Z
DxipXXxb8qv2nep6Z5HtvYGh60NjnPhWFgiwdBS314CJylh5cRzPFmMTGd3lciBp
NYaqCcUcsBB9RN1+TS+S/CSDj93mi8YziBIA05IDCLbPKr+XTK/b2tslVvPXsV+x
fSEImXUj1tYurJO5pekuz31KblbF7GyKWBrQ5koN9C9lLFQxprLnsl6aXhADG/tu
rh8OT5QPytmg55kcgKcoUYGKxizg57GQQElK6zp7xfnpBthJLZt6oiGxnNXQ7pn6
IUvwe1QRMefCaspvsGyBXRTi619fv2B0WOFzfzcwW5Xq8yWT6+t0lJY8BbKw4OST
qtMoyu3jrbf6UaAhKukHsVIgvoMo8yKb1we/7q0IyV8o9/UfGy5aw4fGNhqyX3W/
bG6QEa3w1qdD5aKMCqQeThs0TPbU0uKngNxJOxTFCrdLzTAVbw6LLr7nkCgR4dAe
3XpE10KNBJkyTg9ZGLlyemh7IHAlLMAmwvtLJSDttivAvcBkLjpVFmH3JoVhqIAb
pwChZKfr+0ysLbSZDQZunhZQaXcJmM+ST3M9imUjmtAm5kU7zlN9r0aN1LeyDqdP
QW8S9xb2ImC4uHa5b7Cz6Q0I87QBiNpvAuUM70KNS//4ziA2ZA2j5tNfsgSNU92y
aBhuLksmsARh5bYniyo+PBI6yWh/IiKb6PH+t7jEQ0ZmOuLav+HZ4SYHRFGZ3iIl
l6dNELw2zi1VsAlTOg/6I1X/rD96OHJoAncdyDrbHXpulETWfz0iKC70g5vmTLOq
1kkOht2CwoFYFH9XZrphiLhwGzx5vpcHRaze9kkerJzku+U9HPYx4MXeOn+nlxBR
BroMsUS19q9A+uE6Kt99IWguBHfKtRP3E3nRD44JvtwbiZqdMcdZ/XHw1K84j5vB
W2KuySVXvy2Di2Btfw1OuszYhfUBuaRYZt8McYLm5OmN7qLjGuMV/bguedXMhY/G
XL1/+oOlLI/kb/s3h2AskhD0AAkgTmPxPvlTlWgEraMPFKLcD96nLfaALVSo0k7b
hz0t+0kdWAibmC1kavnz0IdWx7Ix15pyKUgPd/b7eYyQrDwPp6lHSq6s5MEslFwe
N/721pTYmuWo4otAuKDAWT7U3/cBvIwCvU65qayh9v1N7BYkCKB44+LLwgFeD50U
N6Fjn7DSCjP7M14H/SgHfazUSyqdfExm5fAkgjT68jOGJtg49B8xqlF+QruEkQNS
qt21l7cRHGDMRzMVM1s6a8PMc909yHDq5YbdFuBnNJbpgAEMmMp5gGI7SCByrkER
DsJF2IpL5gSe0Zeueqh82K6uFH8sKF1IJED487JzSklr7eQhzmVnqVmHONHjzzYZ
zPvH3Pd0n/oVAeAwvvW9KZSK7qXLUn/BJHiHY0n//677jJFYZE3qUVxksrOnaQ1I
ddJOstCO2Xldt1Hed6n6v58tRoA6SAcVRzEe3x4WfOCl9XcgqxxgnqqaGqVtFZ/u
ZjwfD9SWP+0ecvAMAosbnD0FCPji4XUIprji65gefiVLNT694PNpE+DQhW7dT9zv
L3nYOC5khZnLMxS3N8bSdl3KBsAKCfy9aH7YfR+1+SyiH26mJqrKFnZ4NrzVoMmR
5cwpZ8DjeuNLzteD0nuPuqPZlwuv2WlSvC672TuZZ9Qx1ZW9HrqDiCJMrKF8TGHM
3tP5CoboRqh8dFwUwWN8YoFyzJIpqoltCi4XS/McWZA0NfEEbxIVcQxNJQjKaM1P
C03OgN/0+V97w8knqULi43kZ++OJerpH5WRNCNWs1+bl51vQDqzKmad8svqbxGED
E0pU6rkCNS+QLKtoW0Ms2xDQxBJfjNYt04tMi976xG8nXxGeZz5YVtB8xmHA4wui
MMqfwU6jKivgduAXlnaIbgxgjNeEZBFn7VhVYWtcwwTZQH15+i9YnjUqyoIJI8WX
dj8gnJtDlLgtz5GXutniAjjwbUVKwsljLm+zyq1jyE+85RY6IBPUFLbt1W9YEgAc
8XGtDivNALng7czwmQJQjMqnodjcH3FoXs8QUM8AXgs5MqL2yc7EwXyCMOkXk6/v
fmD1qL633TPHlELlqPJPxo4R+4ykEQRHjxZlIsUSQ6RK/BctkXATfJJ88QQhsQCx
QXEcrblD1VnmpC64D9SFjANI0okKGbM5BiVd6J43PNZcpbqx/lrhOGAbb5E53Aen
KwPLExYpgANo50+KBxucJc1CGt6/+ZqqUzGeHOMnp3z2v/inlamSkU+SYoCP3Lu9
KQgGF5arujX6H//VMlt/JTo0AkK3qpvxYk4Noy9JmotERe00NfGI8dnuuxsgTlGr
ZKjRfvWhPiQpXIRLh52SD4Yg/F/pS4Odmw3bWABr1iBU+QMZGTVL7fYObIuEJTxS
qg8mklpZeWZl6+4GC6nK4Fabl38EsZ1cpuV60QpL/j64kzWPWdE0WCPosWuQubEz
n/tsMJtuTA81QQm1OHLu0vyorCXIZEScywd+uaT0v/eRVLAHqprx0pzA/zM9Wxuj
aiheImfbfIdqkFXbgqw9+TvuAFkQqb5g5mzYixn0iJfLh5K5A5FY6NXsyrCNdWm8
Fq2ah6CGC0Oww2Ml2Xbntm+SE6jDBMMRma2tLnC8rXOWFszSVGmpDeG3BW2XPvPh
9dkFv6KAzNTzP3J6VRWIViQVpv/I7j+Xo6j8TROzMDClviqT01QiSlR2n5Zv0dy+
6ElkExzUbEktDvT2xJ/AYz5qlW1pumXG8cuQ0IUt3OQp6CAExiskt6x2iaSj5EHt
KqEfSDoM7nAgtmAByip+Dc8NGYqBvvPxWVTt4i0i3TQJ0FHRz2iffqpZ6DFTw/Ft
7Oqebeubh3GLpiMsmCX4hxZ0P7fAyqSFWvvEEW2xDhE6t+VAD2qcMXhXnyBFAhRu
exS2LfkL8+g/HS+0Gdd71senp7ya2PbFasZ40uEPZBuj8+wB+9Vs3PRrMpDRfKDa
BajUTuD1hur+FQRhTMtxhT6o4PRcnqDhu8BAS2MH2WqoaTS6pMC3zFfbkpnaDnMz
rIZnHbQRvj3HZWlwfxyLHuQXEg/tUc8IBXzRQpAeikSjBU7D5gt/r4H13h5qhTl9
nO4B6NDRp9/3rS0KMvtwIMbwIoj6jYDD+B7LIvSdAsJzgrzqF0eZQ7yatMaFcAxo
jNEnZh0ThzvHq+bjGmO0RZ45rBIew6yMkr+l+7Fun2S1w7tqtddNNAx19BeLVpz+
z+baZA2FwT22ynLyHnmAxRt7aYvj4ObOOghNvhdGBUl4cOBPHtGZ0X1iK/o1CPXG
GZ8SBBmd6wUXlWqnOVRQoYVXzJQ1nClZCndxiyFI5cUV4zsoNTWJBh5SJqdBxfGz
8DOTOxMccgfDkbW6RvxszsPrFW29FSySbwrDD8M4/aWfvJqegpslpTVDWeyCPQ/b
WnbVIkwjwaeNNRwikXnmVnAop2ENUkyADpodBPjuYfevgoikaP36X+Eu+OxdVQKp
qjQbsRKwFN7DmoNwRG3ORyF0NMiifykZuhFBZ8awlt/4uGkH+7T8j3CJ1ZUgqsNX
Sang1FWC6OgAm7Xx1op3/Dh9HUhCHr2SKgBPqfkMF2uKLEY/fIIhRwHBoRZ/uc9Z
MDe3AAxOfVUdkoQ/weNprVrndaPdjU2y1d9R3OQfMbIesIm6alHqPpEluyNembQe
HvG+CxgfswtaG/Fd2tfkdwHXw0FFBJp1InUkce9lIPadRTUkAIkauMQxH4vRatiO
Yq+geU5ePgkqFgwYVpvvomChbPMHOhfB6kj5uejYBPDwMa60NZWeIm1NsEW5H6gB
pphI7ViEIw+sYWbCFA5+h+fAV5XnpjXj3FMen+UiK2SbbkiZ7Se23FaFgwcS/bID
vBlneHoaW4A6yD8gWqJgbUzIMccQd18qfwAjTE2GsgNekkoXybxy23G2CdftUMOX
27ImbyAUmREip0tyKpP2hZg6/oIlbHgUEbcMNtBQa8SODu61fDf4al/3bCyammq7
uppMbpAFMM0p/p9fwIsNAOAsDPEfPAEWTc98LWtR5C4f6J3gtTQ8bBlLPwgcs1v6
9HGq7wep0gv0y+dv3UDtUoSlGLST6t69FfMlId696QQDeDxN1sptvye8cdcG6Xgc
NSqndY6tX2AX+WykGH4SNsXbhGEUGPO58++758lO0iAD/zj/DBExTl2Yfp59zm+n
i5YkDTwQNvpFfgJ+sxQYFcVD9j39jx740H1GoXxV8aG/wnOjXBKeD4FfmQ9rp0JZ
frxI/Rp8ts4hNTNay8jtyXZ4tBv2ZcfR/vl5RmUHQNgLALUeHLdzfx27Skm96JQd
z03Lfly+IQ1EXNlhh0wNmOhfe2o3DEj7XV39SiumHlX2Fa8NatXPmfiG8h8q2QgS
JIM9/1V4Q+hY839o6fOruYUwMxW2ihpOKpUJlv0ONpBoh1lXH6hVlIZ+vKektKtT
sYXYPd2eIKysgRK4ddbcjXpF0/KFKFEsMCr9CnNuhscAsIg7K9Gd1yYEQHuaTOVc
CddVTee8uNOQVXgC+8iLUuKjq/4jrCBXOFcxdNX4baddvlRPyQBnpbHoUqMzGJKU
ByRMfn4aKL7I2CRJHMRcU0nezn61Z1OqLYJEyd+IG3OOgkjquALdtT+JEdwBhU+2
0klfmPA/rrWgnDC+r0kfvVgoYLkjjix3NdMAfukEzkPaxwaIJ5owbvJmySeg5/Xi
gqCmp/RuZrNoIw0T/b5XE6EDGpulQHSaDr8bEF3reS2lncOiz6docUyqpFbXOs5u
YEWHqZqfFkkVqjo2iSA2zwi8RDPnLHfuwpfeQuKQFevJreVCwe7/8QWlxkYCOqVc
ZmEJj99DpLTTuWWYDWQWz5j9auci+1aNusRcCI0K+i21UxeKnO0A98g2AMsMF0C4
y7MNhRJJXjmh6wE5YU8R+gdrwGw2eJvzwTbL04HEu4q9lrO+pROoyIP2qMPBaP24
tWvK8k6guLr6o0racOUO4oa6n6O7VYqJRs8JRq57NiuG1ixHDhVa5iZr0OJ/hegC
SgOJv6SUg9yVGYUkTUt81Yl+ojYYxtEwW1y0gS7FmJjHcP9ax8iR93un28gOAsOd
hBiEGOT3/e8A7aRqHIfscG/3K5BrxkO1R8/vTK5wckVu9ey9HSERluoIi7T8ZLzB
B0bkJUeyoj5xwF9ROL8UQD+RiLmoIt7RNFxoOmJJ3cpWZHqpMbwAJGJN774eoO8N
P2CHcBBkSZb4DzKP5YyfGbmoLvlBbUXlAMQIXoYdbt2/6cmn0Lq5bD0jDURmAot2
Zhs9MT2aBn1hhH1YKEhB/R1WBWfdUDU/vst6f5s5ek2+q1YSUgYpJRqy1CVchM7r
uiZfJtSPmQBwgXcfOt82CsVjPsHPW9XD/1Y064j5jXXdgs8Wv0tZKrRJ9ayqY2o9
UaoXbbb842hMrWUfHt70EssypmJfznX+a2PbA6p7ffPFU0vbJAUeJn+vgALoLVS8
6fj/jc1mwrYHCHNG6n701D2/P3NlAt/zSDmJ39V+gs1RUYZrwiQUb4uW3eQA27Fx
dLwpFI2TC2QflngciJG7WsYdOI2gv0mcPD75tgVep1WQFROZXTxyLMgxNOc7tItt
+QrSjXkNbiffhAH5v1DU2UbHwIMN5ijDJL1uBVqYOE/ZxYR411s+QPLCzh1lCj+9
ZoyxKKDein0P2ydjdZY1qJykTySwt9/hHoxMmboCVKze0g0tkQD8b1C/lg+GyM5s
POHHrdaGOXy4KsgRUhjmcGhBInRDczmxeLsFgZdSZi+MFXWExCpeY6yPRP+VZHT+
xHVSCzA1v8ISbBttZIxMyURqHhfLEJz2MJJ2tI4Mo4TvBBXe6tmatsR2hs5StaXa
zbFqFWUXw9XcMd1uUqNNHi16sMKbxNQej1kSXiIdAAVBldxfg+0ED+VDXjrKcMJh
WEbuSq42ehtBaYx5UoffrRABoB91P8+da/7xnRoQ6AeiW7/XOWOqWkIb6fSR9kqG
3PkYDZnv1AzK/SuNxJtO60jhq5JW9fW6/ZnLpPX4TcIAfnDi0EijFl6qphbJUudH
us9ofkvtB6XAa6Y5ozPnZnREZJHXyf0Du/AsopBAHBYUvazcF6DZOE7fCQ1hOhNr
yqNgn6KBNsbTmClZZrDyV55gfmclTpGijD7Fkasm1LlAMVnzZbf1e1QPOww4Iljg
OUm01hbKuh5lgBW+q344janGt5uHpLJBVlGAP5624dp00wj+v2k/yz99bz27aVsZ
3QEz8OVGdhF+esVdhfX0vsdC3APJajs3E9MRhbrQ1p57gqjWis1y7+CFKIe4sRz1
57G8bsk01GnB/fRwsOySbcHVryZbDXw46Nnn+nbVOmRelIrL00pmrDQjEMkmKHoT
oJQUvK+WmF/lFWbsE1wrwbSuYS1bzNiv7GrLyquTVPvQu9bMYJapJwqwdJMXfS91
av/dRT6EPNFM9Q7dlYKRQ1s5clkBugdu5mmryBo+hE5G667lZL2qacDopXWe2mvY
r1waQjVZk61V9v425jLuQj9t0icJ1hh0K1tRRBfIhGOqKgt1LjIN83qJebjaEt2j
IgYsFP+4+6pF2J4amS6KbMpBMl8i5H8F+YbtkruMDATM9Px4CP6lYR0Jx26TKSwF
IK+iJbSdcDWm8vG+r3SlhYjcfmkayPalLYmqRslCJHpuU0+GlhmlEGIoafqTr5G6
pT39BuyH3ASVEzS7y2b86TULcruh4PZHo5Vd9n/WINh8WcBfKNL1hGCudXfVLgRs
+unnBnyah/isfELRiskfixl1ItwfFsCCOufNsf+ROsiayXr6ArEDxBd66yYpyGUZ
svZ0BoD+JnlrJrkL5ZHcbRUil1ARs0HGicwsEEyuBijZVxMZ87pWRRRgmd7n0Qft
jEaz7AhoPgQ9rPkGlst4ltH3XYvIouvu84vszr3SOw/8IMxah184QnUq5yyZhkTj
qz42B2A4x2BnOwLnr6Rbe3nIB7ayk0Y8vK41wyGzK+FhV9HjUVzkqJYv6ja3iVyK
tpwmyZGBJEySxqXv6ZyVbN0b4BUHiLPQfC9O9nR6L1DGb0xrF8Fs3MyWafP0z6pg
v+QMk3MhSjtUe0swJBznkMKKK8TmGx+S3GWCdc6rs6EYV48Bfz3G2DpIIHHtR3r5
rcfdpPJeRSZ/8d/H8MWDQaCnBEMfySrjmcrSCAkQcEOuGcGFkJpak1f3z+nqU0FY
ZAyOIwJBxvtCZQRHGp4eZAfsVPwAVcsIMuRQLOYC5akEJG6qODy9RqLJZLwNfufV
IujkL3ij0c13Sxf7rJxbn4FAHBFlmPEt1OUpWtnZDV8lfyNHF24ieG3LpIAC8s7r
xsZP/LFWUHZM9FoMS0rkRHfji9bFfOWHwAdwGzRAwChGsQaQxrYPPB20AGrS8V/f
Ruo0RNaNPPGwYDrSPkKAFREPsRlI3NmZ5puiyiZPO/J/+RLvQCgVy4yrt+DIrK1/
v2eYGUHFqWTew5MMN6JHVnFGuy77sud5B8ErwhmjtQGSXk4N167rhboLHvPWeNh3
+r1VGnAwesn/Wu2ypdcCJ4KYhIeQkrYJfpe67X5Ye2qidnlI+eupIsi6EvQC3Wby
A5N8sfXmXekhY1FA7x52mrmHamPjDTVvl+mLdfl0N8d3BeABXv14Hnk/SCkJLlGH
tfGlxZjZdbSxoA1RNtQUOQiltDaz/9A3JQQ8H34iPVm8iNWuTCjreX0ykG8AAF/h
5pqJr250IhZE+CDmQl5o/XpOaKpZhcMRSCRlcMaU1d6eIZRcTNdTCz1OtNJp9oGi
E6NFvpdYi0eN0szERKwWdyOLQqD2mkyYiDakg6JdWA+fpdANx2RsB641NLvb+/lT
nR7cnD4u2pfxkBhGEEM5lWHrVGomnlHdGySrFcCjpJIxqlfSQn12pHC7qMtm9sOq
izIhbFTsHOhpQGF66jroeWj7kdGqXmgluPbwMaBmV+SiGdIYXMivdcVohyVFqinV
wf1Mt/suqLNIpIZPS2xJIB2HXJXsrcWzx0a7ewRuf4aNyB/EEQNkIHHWnW4kzYNt
Z9xAU3t0RgWvYcK/rb0b8C1hyKnF/dIfOgvkcBuevrD9kOMW+/gkzD8/rbuKEBwI
vBH6poAACWJRFiij8hMvWkKtD5rDye3MAYMPiMQhgSE/wwM3w3bGJiyNQ/3pl4MK
awyYvAfaAQu5UezW9P6MQnXsjLBfpDWRkInjOWEVuTd9C6Fa+/UruhdRaKWsfvzw
6ry6sr/siOSTrCDxAG0O3ovEbVtl0vJh7roQrnxXXwtwfCNYX1xVRQSQD0RKjmm6
fbL9VodE9vhtIByIneA1RN1mFOgY2PACQqFDZzZMk+o65kDsPXzz/JVQsUZnuHNp
XBt0Zimxi0MxA9m8Os2kD1LsInnIyh7l2VVDgVgQhEvvw0T6M/YtZSMXzVyoFf4M
NLw4zpQ8yZvvPSFivJuDl6Gg2VYJGNh2WwxLuZoJEKnalMpt/RdRWpFPcUSNOUwO
jhJlUTU2DHjGvbKKihYMu/DKxCohc2DFQGHCBkSYYNRD7gnwmaxnEl7yoibK4KfM
XLNVuajATrVviaio7u5JZUReR1xPYjxkrAKnBTT87SA7nzxOgbZ02OTXpIFYVQR7
msTqdTHCNMlDkqncyxwk0ooEe8lcdAlFwvuYQ0lRjT3LTS1u/IBguCZemnHT8XfM
TNV1qWJxW0jm43CvxImkVH2ZP5c84lVa8P/juoRt4qSlRVcygemKyntX0usUkIMX
RhahOAlH7yaRzH6t2Bp+n8bo6n+yjYk9JtbuYv9ydT+TbkQL/IYkr9Rx+bmWky4B
zgUUzwBzPiES0KLIq4kUpPuTmN9UQTD1kJkcQiJ9+Bj+TNZhzWQ9fRVnEifV0Iwz
ilqHl0Ar1dOB98pDRBbwuYrcXQS9QA+7VDQkJndvXPenyfPXyTC8P5nAa29pokz+
Rpi0bN4r7yL/7pk/M3YE/KX7Z3pd/eWLCHZrRjnU7eYIotMHCb+oK3OlBjgmkLxm
0ncwRJ6OtxJqcKC9u01126QCZi5t5zMKfO2SvK3spgnAI+j1o6NilB1InO0wXjnP
3QvHm302XMgofUBeKQTH8szwwp9bmTRhXR1tR5imSSxHqAMKm3REiLEjHIzAq0CZ
EauM4XgsbVeEEoLKnpZwJsynO8HYgRu2Ba/4BAaKKpFjUWKZfr524GfgcXlKg+TV
7wPvC8yvCkuIund0yj2TD2yk3GD9/nhQyfhHAOuQj+PysgUx7cMi+vFFotLJyfPZ
uzxG9W+cLDm4A/NnlSGhOxrQg+epZSvvQ4iL1MUAvrrDQH3NqGBVe56/uVVA7J6Q
seB47iMHeDnJM5bsRcH81TRAFpWIe7oaB+0OYD0tXMh18RY7QxSicbS/9OAMBeNB
NSMEutcetFPFxVLYObVuH7LfPbzH2g9l3S3AxS050lvHCKcc12l2z5vSUM4GldRM
F7ro1ytjq5DAyd1O/NXlE5BgovvETQUpyUxjbrlUeSTUcM2UMvQ9lW/oQAcVjak3
DQ1uiAtUTM5AktIRCGbPL3m35FCbya39lb42WGSt86MbpTk32NMvenJIE+iMNXT7
bV7PMGIGSlk2ktqJiw8SHD0qksHqR2Apg+az8Lg3MSvnO5XBsjVUU2QR5wu+FrCI
q4Y3Cm4ZGoqCCgLfuzznSf6FNJHG7CnQo67NGfkRr8K+WNLKf9eJdO2za+b0+pkX
FnW1XjSwhVytGgE4GLazQL3Ld0S/TJ444gKrzzYHysAxlTxSec8qRdoJIM8vTDDT
OUvlzvEsp7JVM1hCpWvnNNz6WQV4aQNc9DwXB7NUQxD4MxxyAM5w3EM+YFpciveg
tAKaklvG//+VsDPgglOdyLsSORGQPXTdYN4DdjG0NyuhHngIN8vfMoxO6X0fe9dg
ZEKXDW9f4M1/6Do5ZHHmJkrPRBIY8WowtE6HGXQ7pMendcgJUN8lKyG0DzvCScZP
becYOo/1krVmg0vazZHkyY/6Obq4NbioUbpezXYuHyF43eG6Q04XQ6DG58scPnB2
EE/eHxCZas9tkPuic+zC/DzS9EFBfHnJjJ+6M3av0nDT2fcANQhYYOZSJBzuKuoy
kgUL1MPrHDofDIJ7IOr2L13chgbUfjrNvLmmPR7hbiIRfGm5UJD7AY3Rd8ZlYQ4k
Xw+7UxXZ3QYFSt88FhwTFblUTQW+CWGGyHMB4/yleImKNiOWEs4ZRMpOVYPDaVmV
92L1o/FGjicmsOG2pnf4mB7X+6x67qVLM/yB2shSo9qg6qaDaaFe5UCtdLwR0kS8
fZeTjKnbJXYgU+O4EJzMAgpI+umN4BQtc8MqEDH0LN6gy9AZaJQaQ+oyX83tceMr
XvGytuiZTdSoJypbzXXKXIcvDEc9FCh4mBxYi1hW32xPNXYrbjGWtPTv6U/riHSD
xehlbDMbXE0n2MIkJd6S/Zoozp6LkbSndlvFZ9dMIQMEuSf3GXQOQPCV77xFHhjq
iegKZ7whfdEFY6HnvA1RXBFyVQVWGqrNG2FK8YVSbXc1j/aA/J9+QkWrPUGjww6e
Ssb5d5nwHzkOkKm9N5f9HoT61sy5Rgo0XRYmqNnj9GhpuDDDgiPe6gZeDOz56VON
6ltCQAunBoOFgAUMUeu7SJ/ScrgGfvDPpK3gPHKDRQImA3M7IKD5kVtskyGOtnXx
F0Mh98h/mzOnCnqBKFEbR4L00KQb1urDM69ZLtKcHR4DEiNz/DpXaQdyPk3VzfIi
giYafuzsJUQOkUp0we1hefAXhMLx2D8UdFzkNsqN9ARysZiozia6aNkBsCeleqpC
7Ho6xOt4DB79YEQQ38MkvF8BBzJhtxEa5+AcWuIAVtLKg8kaHDHYxexOSQ8OiFIA
aQF27cN70J/MV38fpLNzHJLS12b7KpJyHVs4PE0rm2tpX6nZLkgJzfouXCEcSYOf
FZwMvyHtL0Az+7xp0hrt4y8Vn+lzL6WRqA2ygjE80tGzDweOj1qOyky2gr6GUw/Y
wciw3VeY7kHglZtk4CIxUeppd/m7AIw+YvdAEHlS3UhBGNkekesJdmk890dkxN05
5nFKrtINiLmmXy/HbWNx7RyU54GRYI+yT5XTwh4BOyEQQHxCeQMDccKAWPjTT33c
8eWonF0JdP0ucSuHqEwl0RJbM3UrdH+OkQMbozM+44yPP/+k2JQbtEPxVmvKFwu1
2CpOJzR3lT4C2OvJ3M4g1vSKXgQj8tH156Y+vOqIt5c/utz4R97+b4G4vtO4pyXZ
tjKGDPIj8TVd3z8M+EbKW6h+QRvjuhYBDDeQsZMb557FzBA/509PwVQHQvmIHvOu
v2k0svuC84Z5v4aqQUJf4x1mcqvy9nagC2E0RhMOxQU1Avmq50KvYMTdNL74RErf
ySXHj+Uckq3rfq7Yk2CDeHizw2ZGXhqgFq+RDGCQQl2E3SCR1GEgroeNkvhnu+/L
Do3W/22JshoonbPVcDBy5bsFo0MJLTCQecihKPEHJ0RWZo2/zZ0D0KZ9k5Fshz6E
AhOasy7dRJ14i+OBIz7OzOaSyI/C4mRkRM8L9vCWew8lS2+HQuKLNXfKEVUv+7ji
mxhPPZGQfvzhcK1oa2uKBljyWKUEy8T713sVdwtWhy06vGJs4WQacmpU/uxeRtjJ
VZ+5wLTpH1bnO40lwTPO9bJyhZs58yetrHd8zqxilO/Hqae5TRZJXJGIJ//2PdAq
LH+Y9gmfLm6PwPzsQTtl3WrG7o61H09OysF5TzyhFayWTSoq1WqOUlag7aQDXPIt
gFK8LQoc9Bmk+phXEQS2tpZxo7Yid7jdwURNnNZFBRCzpkxFiLF7SY60eato4ZoC
9CtVAAanU1UQBR83aQCs8aeOAKcm/kVhS63hc4DeYJsYknrCzLn+gbigisw5S+4v
yluIqT2CTC9YaUtITg/dJi3GqOpe5yNw9ZWqQ4oyC72/Vr1+M7A8zOIqcuJFn3AB
GmHqlt3fwvlefYADWC8ylCRleSllBMQRayRXqX+AQl2+voJhGjzz7ZbqTggccals
GioEsabBK14WNlZXZnNCWJcadreVCCQcWqLgsK2/SnD0UP4U4DzHRunRBpWVqq91
tR8VAyO9joknWSUGKPMzqZ4oAVEpwW1LXyZBFx3Y2RB92uN5U3dDt1LW7OBZO702
cKJHsg/U9gjmg72ySVSc3a6JPF0OH47qt3w4Qn0bxKsxXO22hfzLxsLOTxtqwSYN
7Ujwraxs9Jq0aFIiqHHAJycZPbJ2N23mrN8283BN9uklXrkop8fbeKqeoSqQxcuL
ElCe7fyCjYmt7I+5XaXzr3IBVIF/kTaavyrS9FL1jex5E1LTsdniY0lBPLzcAr3K
TTCookYYNsxIqQsOnb35MykFSy24hWqF1PQhecV6yUPN8S9nfvoFyqtsxPcLJ+IG
HkurvWJq70VYscrydWF2HxlDvdhcg3oLfeojvs9WXCr4pWKyWfId1Xdvrz4/0uRU
85TRhehDX6UJ4a3blljMJ8BmY42AYg6QRFgRMqgvpODLh/+wdP57pmmGcp/22zxG
p+aSX/+E1oJ2U4zKArReUrXgjRd0m9JR+c+Yvf0oUrGW5Ga6/R2WpblPuj1aAIme
QukOTNEJ4Jj/tX+LQ0UU3Ab9sXQSa8M08EZR06RiwOAsQaqA3RzdlS31gakhBHRY
fzuPTddgVhfOKjKP6Tc2TyZqKeSXqwygLNZg8RuhMWV5/7UW+8JXHHtzwgRkBox3
hqsA1w2X58Ltuiqc89OixWfg7demvhzAd7O4mAf6XmPYYhmJrRS5y/etNn6oEEuk
0BgU5cDs1hHfWorD7fIYly062MdC1QdwTZunNLlHTHc8WCdHgogKKIsYU1ZWc/o1
J9CLo8tkX2pabOZb3wzIycenKbq0wibmXOMxj6ZWhW4KcqQsQYYcLDaMY3FT/BV4
HaBkWSZQ3ZaGFiwMxZITsusITI05ykNgGtVfGflJtNDWEW3oAhwj5A/XwyK0duLh
fQOIJTsqCKYcdb1SBErPX9fjcFymuurOVeruT4ORPIRG4FDagvvIAe35ai3EHa12
Cbi/B+fyPjRtzoWlKXloAnujuvNEkIRZjQ4xoTvHSp7hh1l3f3NtCXBxDKqUqlQ9
TRmPL304FQo4omwQXhwDDfYRXmx4Q3qv3CzqzAwQtNJIml/kvqhsqzHaMS0JqrfA
YI/HbEXTOrm2wb+MCIyCFWJ0CL3Fus5Xir7QdkScPrqF3mkD3n887R1qiUVYEM76
kIGz5xE4Em1D5d0XnUU4nXgahxN4BL6X7Q2/qxtBxNOb8ZJin9efJc8IULJDSaO1
K84gsrRe4JAlx5OnyDfkMop6GmoBFm5GW8sM6uIlSTnYPwBkVb5D1Nq+Yh7Ey5SG
eVbysgLcLk3SC2ZaVhDxtblRiIiYxmcDzzfJg71R8C44UF4R9z1FQHFjO4NrD/3D
PlEWSGrWXbZhSdJddkVHiT5hOUcIjtbb12fcxgd6Adg+DOxVxk1PruD/pki2T7qE
g9BZhqhB+fsIv6NQ2UQWeYTAuajMLFqz80qXGSvSdo05hwwZB/enCWDOWyKP1DY/
k42tjBagdaTKMVmYT8YV0hm0JCoTYiE9y2PiVwsTeXC4wzw2dQfM7Opw8OoYrmqk
rvqtXiSrzp2NDXr9CuW9nDqWnD8+jLGqgn1cztsP3IE54/gGr4dfFTIhcRpJlQW6
v5ohsOliwaO/5yewGYKtAurFLu7WnJ5STyJaeh4Y4Es6p6dmXxh4l+YDyt6GWjGs
qK38FJ2/eGVm9gQH4tAeoCAT2zh7zhhbRI/EnIpbtGdyXrHrXsiLxz7Oucp0wVwx
bMOfjkydSU4/QtNwupS402FJuBEczufCYPHMLETiIa2DQIMEQcwOU4Wy+AOvVQYX
qEbxrdBsOHO/bZNLiyH8Nc4qvLkJqxzqv3kdltuuuf7zJGXq3Lg934PZCwQ9lL2i
yiOxzyeI5dR3mUi8ApRCz2EILsK8szLh5oa9/CSgPeAVIkSNOFBSBNvnXAkGElL5
1ntg2vS7cf1D9tOM+g6KzBohhKSg+EVSByg/+X+hiVUIGBse2Gk+CsaDtNjFAjkG
diJ8JFLIIMpPNK3khuQxkW8QuJOxVZqcIaROHR0CkNtqjHUuPkT7mW1+WoYXw6zq
YQzeGVfgS59uKbRcwoVfh0gRyo7eszCEbcuwM3UsGZQRK3nqgxXPus5NUHN6lGVl
3dan2WRvubjwE+k/9zO0rlzyhA5SodvyxDFEnKBulg+2eFOF/ba5dOrBFs3UTQHN
oKrfBuaRg1zW+jzDBiiQvLkHI1v2Xrb99a50fOCAfnezBXf15Kv0jG0HyUDBouQt
5H0mE5LiK7NjhiJFpY8o6UA5F6ihNKkcy91KdSjqb9fH3wrubhuq5qieHEsOv8QK
atjPtJgh/yZn5W8ZIoi/6rkNlfb9+oK9X34rEXJRRwX88RHCD8blZ7tvN+/r8agT
ICYgRZLTgECHPHgoy9WceRnBpuELgqPpwZseqhPYBYflDI4fws7Mqpcsplb4imOh
5E4rP7RPo7SA+UE/9uRam2Y5t4lyiljBxvetZ0vyDCCVEovAb6NpbBEe8esGk+AF
gutBG5R0f/3PKtFK1SRfCYP3T9TRyUrMqB8scn1ptaqZkdlMvSt2gm0dwUAWqqn4
HJlaAemvkwbxwxXm/IsSOwGV6DUUdWMzlME7nbpdCFsQ9ivu7go6izzL53MpuEq+
uebY2UlUCo6OyCFtFKSn9iyx4blbt8i1OV2cSceL0AVC60KB8uL17lt04hhpV4eX
noWK/UceqWKoIBruWYgLhD48lejAniZyypiWUpFpOUomi4uHNJeUiA0nfqOHe+9Y
7+6mMtaNMCMAjQTAihsJL+RJyDJGKf6LPi7HwcTTYvVsb/QaXUUcQodAxSm/cWQ4
+fs7zcumqwSdK16TU1+5Q5DSHSS61WNsNqwBV8kUrw51TmWssFsx5RBU6eGV/5IO
ros8iTLspYrkh+HztwATe3t6Sz62dO1KN8kREg3vIt31JWL6FF65H1BJ3SzWisML
cDPjmF6j++ILXHVCYa0VmHUFI5G+RScDAdQ9GQgUcltBgWW5ukm1EQZnqxVJXcqX
osMwEtxp/G337e+h24vQ4fFaM5+mZmOBBOiggAPiLb1Gq9to61TYwBpNIretQFyH
wi7wbKGA7gZMe8AFJYq6QuMd7WMPBhGDoDc8O2V/snmeoZpCpwIruXlP/yV1HDqp
CTzO56kaVtItwSIxbAQ7h+FMOcWzSaSRhjV2jp++lDKC0YULt2Bcvg7FMA2PsWLU
dcFPOgHKBdVLrKUtC26Dv+6CQQeYgToT7Ti8KGo0F9tSKu9/PqwW0TvdaiJG56QV
v9vA/qoXOOY7ldSwclrWWtgxoQ8L9/qU6iTHxjHEsxp8X/2oyZSsrFMqUbdmpliq
KIBsrsHy7ylViCuU9xzbV7o4qOdKy6ZTo19pF+pHsyd6nUKc5+HJ8TmjvPRZQthT
IkEHiKv1X73qRYhhGMzKdQ8xD3LynVLSzq+s1TZvtvuF/opKay5+cGfQF3I+BNFh
AqD5w17lkeTW9si3ev9p2W2pA+gJl3iX4muD+fj0E0xqIJXUYJ9OYqL7ApaKWvk3
KVww0qXIomw01BAMWywNuh3Aqu0pbd5qOuymdNhmCZJ5lcj2fHdNpS9IHpPDp2i3
/lnALU5jUKYINE//0YGC1Pxu4TilVRQJ7NivxEyIs527mbQE9DU9DuGMgUle3M++
2ekgp4zK3wSlXNQFbs3+maouUVkZPf2rNBLLs1/cGlwK2+nIBmjexsvoqGi9hRse
ERTIgPZo/j/q3AUZIe5qjw0N5XqYl0/D2ywPguKRGZ+8kMO+nUKBuF3wusBdfrT4
bPBOOda59q//f54sR6cVK+eZYDsSD30wB6RzElgK5qB/p458AnRhwicnHjruySDL
NAYS7GjBVcgM8/0jNji1T44e9q+kjfZoTpXLsliEVl9pXFypkte+RsfAArzm5o7T
VOMAx4iZovzkS6jAhess++4sq+ecsHG37QhcYM/X8l3PrOp4xKXTst96s1ABD9Uw
NCsdYFbbkdn1SIiJb+0YfBPPDcggQCu1GPVQwnZIC/BOTASC7KDOhrmKzaI9o4Yp
RncIQYdJ4U4pWNX1sB1sj5TRa4NJYLBBoT6ZVH8cqb6FHUSxA2796UaZ+fzgZORq
bfyNrcBI9iLO3sF2AbY77bEzgXXjrpD4D82FCLgYS0EGfH6ngt5XDrpS1EZogsyr
J6RE45Rope7BwuugISZGk5UV7zxr+cBrYhMkn8xNH85rwDW85REe/Yym9DZBIszZ
Lrbytbt+ZaR9vpO+orwiBCJiUSen3lp5shQYxWQMyRRa2Xj+LLE+FLDMdEiZJe0f
FHKCrYOwhQ6FEPNUaq04op+iSUIamzosNE24jMRypWsBvbJ22YRBxUDR09ysRSAT
kFKHFAEH4GLIusMGG+qRiMWd1f4lyTDaV0YcBxo2Onc8zppY4djOkBXU8E27Z2KJ
vKXGdA/s9fayn8Sc512rRtMFNa0Cy+JJ+QbcQXJutAlRWg5Yu/3InKtiuOdSno7o
MGjAzWU+BcFF8mZSywDN/tU81rCeLCFrupGPQahkpBQI3fJI+953/2ItKCSrcMMg
tODMwiGLeitygaoTZPb6hVms42oU4xvR9vfs9kqUHIeULYPN/8AOJBa9iwW3COXU
Ci+ajbPo9oMAwxc0a4/aymPo3qHTHpMtZs+j4/v+CkLgR6Q4kXj/P6FsSShBxtZc
GArwpQUAN7MDUmt7o7wlGbNPadvS+bp+qw7p5Kt71+6hFUVs8D8ntXCakahF4Nfo
FV81kjLlRqrCLmZuW+Dnfmq6KKgFAjDd9g2jtuYP3AfGCyxONPPWXtmKKh9zJgBM
KwFUl6eOAkXE+mIqO5o4ByrPnBLZ7uglhE2HOi96nT/n7fglO3e8sOvo+NEN15X9
ZOEkGIWD29K1CRqLybpLFylDWIzYVpG3HVl1NIR9DC5b67Ycv093+dTE93zCKzcB
SaaV2LpjuYWxhLILItzvp47iIn8QQ9SUAqcyW+pB7lwIYfccR4KC/Kgo1zUJoJtQ
VV/kVOcIm5L/VIYf5wZsc1Ml5pLU8Vd0yE5BAwXE0Kl7POhsYWzKvWPQLUAO39nT
MrUoLpR/QSG4WhmH3HweWiAMt6ZSEtTp0MV64n1/IqyKjReJCRZXkqwPAZ/47074
7M2v2tIn36X2OV7Bu3y48Zewl5Gv/YNPSQBC5p5iW9NHUCaGQGbnuSlY3C9W4aVC
6NwP5i8J/3TQKhzs8pBLurM/7aHi/oCAQwVh3EkqHQPyQbodTMo0wxcWG9xgnQgP
FXEjZorjerdDZAlObRxsJfDeCVlVUPAq7o0lrruy3X6ryms1P/gNRAysblKIuvk5
o+iv3ZvgDwcSnNDM0f5vKs8eFmneBOLGGFAIOTw76kUa39wIUiVsO+6Ei9HC3Uqf
XS8jd8ABbqjBgQHh/0k8Um4qK6EPSqTD3K2eNvbRoGmiUeeWkWm7uzSYFQxUYoMh
Ktn6T65EMB/xrv9afDt/OFUkrED0o7CVU0QuuhxZ2x0pHRwUlP0/YdpTrpCBK1Gn
a4owH2oSkBu9BttqfcAjLUHeT2drmivK6pJ9oPdE8d2eWZvkuzlC7qmJWfPYuJE2
BoC1Tf7WRXRFRWnzTNoPvqLq3QOEjJ4O7OCbria/Z+UHy0gfFBAoB2V7BFeSE6cc
y7PvmGnV1jfu4K1zJjCaMxMZt8BpQIkWOS7ruLKOFbjYLbfFOG4hul/zjMSMsiH7
b5Bktvtm7iB8ZmxVCp0WpxOV7joEDY1WKjCcIGsmGIzROoCT/jdtt55KVdyviJPj
P8kAICDPRL89+WPQH+qxNNumx9cIuJ6s6GfmlbdQ4b5IwawL7LlWiilxHO2UvwoQ
OPrOxh2RWeXWF4Nr8H2KsCWQa369SpZaY+VOBLlctXT50YpUEOz69O4CKvGy31Hj
hIrM2tZ4c2+5yJPSbZitXK+NDjRf3doQHhLYZsEJ05pmlR0Ucn8VJE6jhDh2BxLx
+Afta+95p9/KvTblZ5cHKlQKfPRSq7MoR/aTM8q/QK9jwRl7Q+mt8dxvKN1C0eRb
CdKhYZZ4DN2C5D2tUgpRvd5RfOU8QXgsXTuYCvYrDbmwZlBZ36apZexL3T9yAfgy
kUNs/aC8bwvYwAv+6uWGcn/7eSQq9dEbgoKjKlLIQp12LTXfmbT1ere2KO8fVbQ8
sXtTMyeW719SIChhrX21l1wXTCvnRTO8Qrp86VVIyM+uCpwXy10E1pm1MW1rTDro
zZpe6Rln7BS6CVv8W2TgT7St7lu9OpJ04rPkzkQjV5jZ0CPFmODgJ4om05Zxndxi
gyVlbaLQlCRhbrvvKydvJf6kB0VJgCLXyiS16ZFULzOeBfSP7VnX8ntqlaO7qtYR
oP0TSAYNwLVcSCHv07mMXbcvD7R7pZorSUBpKmtiFbEKaF4aul3HZZibQWtNWBSW
e56IGU9pAQlhImw7tCKSTn1wYWSE6TTnqFSBVvDzhGjwyWDRMSiBVIzUOP0FWPfH
0Id4wwBt6YfCDSL3MelTzj9DXHwZtK5dVl3SzQVRre6seE+IL/as/di9fXp21OzD
1c55pPV8iTjn+/n68ZAG8I+KHvTmRh40LIjwZsZwiHePtkBuUYBs8BlkMG5p/Udj
SzRb1z1kDxUz+uNk1YVm6AS3WjtASTm1BBjzgU2yBwd2b3hgdLVloq8yGUYTF+JK
rDcmn6PKxt72h8xgrRHUbetiqTNa4r/NsIBmBKi+mN0ekB/zUaj/c8gWOAO6CcdK
8czdms6y8EOGfOnGfAMztKjqv0jMdymZvKUcdT9gAEWQI28rmX8yNBQeHnm590t4
PyRwTkKCqrS4/9Jxae7HoFivoq/iDUGWJ2Q8atqCAO1Yv56QoShogjf9RIe+1jJd
pNfAy2V5n+TVjaTebxAMeczt+FVpWse20PDm0u1pV5zFiRfFVXyP3fvZRv3qYjP1
y/UK0/OL8lCYhuseOc6Cmv1IIwgzc3UUWfW7gepCHML87N+2N07CUmqKcaj8yXpr
vS3bsy6/Z7cHwmD5Sa+51ztraUeQbX1Q3TqXD1mNOWv+4Nsd3oImVkR7fQtQXpFB
qYVNC+PE5l/oX08W8sQIf3eRDCDm/MCIF4D9IX4IH9WHyh3ZVrdJ55GKievCgHjK
3NNRUnmuXb/scijaZ2615Y2RFHabEdm8bvmKchVamok4vLyrWrjy1uKzZBeot5Sk
x5dQLsCC6B5ixt1DcRwTZFpiSVyVF3WPDbgFgYcMTqmT866az4MFkQgDWAZDPy4L
XYGsNpK977e+ZmPg5+sZhQRagZKP0m2EEfFQiO0hrrZ2/h93DgMhNbHRD9CIBT9Y
j9NDqTglzgpusmaS1ZfC8dR01BP/1E11FzahpK4SDON6uSnkKghJrKx2vHoO4UBY
L4aoUU7b9T+LaqWpedSx+k50LMXscXaMDtDC17pK0Dzdv05grzfQbb6iZjNgvCmX
A7BpSzLY85wZuUrucSZhecG3eicDiH1VLMAv+AEQl2e8eORL29eIwct1OH35piL4
ICy8fmf3o8cietqySFJGLU0fHrZraJelCRGjjkD52NZZ8B+l3wDo7Kta+4uhaTcF
1lI962eEQXaRajiDYj7+NYQ+5/Be8tV/p7ZUIbSJKRa0NVERPv+fgxNFx12YsFcc
Ztpy68Drj116bnVlDkGDzw8I25aSb6jqqjE7ZcxaOVDXhL4wm+PyD/K5AQMzr/hD
LzthPmNtKc7NiWWGJh1V1D3V94mED1vgJgi3uxRqwuWVfQFlKEfAvNjVU/lhpr42
/rhF+NrLByHul0vjdWHW/JGjB62zW9UOxmQcpSm6bQL8aa43KbZQpWN1bnoucMBc
y17nR+zsqN/E9AEBY0/ZaFavvxLeghGyiffBdA5/yvhiDkQxquyxgjDv2jWUs9K6
jnjgdIdTUHFGCqPyecWoZltp4+9nLygHDUH78iEMsZua7Nwnvt7ufi6R+swtEwGO
9//nOLGaOcHT8qw6Fjpo7wjIY8+maIhkPuRl92gjjUgdqIfTQsEQzDBhTTuRKAXP
AcmsSkz4+v/1G32AiPUvpqjKwKsLHzPHKbwmGvfvSZN0ua79JZ9VG3a1MFNoyX8T
CZWJj9iTgF4awu3I2JLWqxya+aNsjLMRF9G5bBZvwkCmCv2arn/CnT6vt3FbQ/Ft
o7W33HcJraDPqPljGkFWj4QsGxC1gzET/df0OUJaKKcF4hCuOYMQI6T1azeDGQdh
stbCeFz+U0BZl8pAvu5IwFeuADohKHb+Eutq4agIXxRKno1EO+okFDVGot1rr6Or
k6cktpDrwL3cr3Z+xcnV6TrGMzrDNR5JF6tieQ74TIX3kSM+XmY6+QxKIxHza+xn
b1L6iU53UBMkzpK6xtGXDhoHmbnlj2OFRxco0Ge04kLy/HSBzFd+LP/S+ewaWDYw
ds7AHjVTtvUrYRSVmfO5QDon0RRxZEe8sW8n4ltN0YxdhFxff3livrCXV/+bipz3
TkMMthIynjZXLBBeFZsxTLxk5gP396+XMRnS8yOLuN8WBvuwnyarEy6DyEM4v9Om
lo8uSZ3C4xH3usA1KYn7SO3SE0fvfCWcfEMIBNv27IChwxH8gcfOt+8l7/MwcgfU
U8W4dOXWurvESI/koikjOA42ydC+STawxGevNDLVIGG1EZmCsd600FONEOUCTYMI
WpTSE/wIBHTDK3TAB73JdR1MYEUwJXMXTPQ/gnYh6fwvXbUM1Tqe6vvIAzOuwebz
yYRInJsE0d5WimNQMgCuOoOCwHAAiRJEpx25pR+KAiOtw+Ji81Ff4S/xBQ8lHdys
V4pDD3ZhQgyPEe4PoRQ8Dc8Pfm7nPAEklEyhGwJYkHKUmBsbO2IlDa6f8/Oprnou
xooRkaMQs3mJ5Lb52CPHIcW084eA9RScN7xjOTXoZQbXfcAp/CkUCE+ArJ4CtAI5
ALaJZz8IzYhIlI3ekvW7gnrxhthuMtb01OnLzk2T9AiSMuWGp3cn0VNL34SzgaKC
KDKgIqjk4SfSNVd6Zz7fuDoc8auQYQOP77eZi8YJT4u0P+RIMeP1p7hXiT+iQtut
AbaOBwdHRoHAh15IIBv/bxoG6azBJAbbtq9XP4YcBI51LmjqMX+UTdjX5p5jhpyO
kFT4cR7+KNFzqwdLQWld1tgC1+ZJwO/5apOi//X/ZGdDUu87a/M2tSsp7lYgHN/K
+lZwU8KCCwtgfjebJkRFcIit5Tj0P9tyvJLCejQnt6rY0SGWSbkgChx5vZqejoOR
avgQDNuL6RJdYRZroyYbo2XIZxfLRIxuPW6UbhWD1VDMrySANsLI5+IqIlRT0qdX
2WW0gfAD0Surs4AjiAIKVaOuJW4RUiRs7M/sagtW2GShJLTQDCHwTSatcVGT8p8M
FB8cuXS7LKrpNVRTHcwWCYYhfo/kw3ztUJHzujPrqdX8cdfyuf/O4yyCaquoiLt0
Qrah7pfeIHcVmMPnXrnixCs4P3/g34RbsQYNCO34bkaHGp/XjMUEHf8H71ogHyKV
XKaXD7RGxbkYJS+PypQwNvlkiyYHTcJN9OpaG5XcCZbdju+1J6vQ+gMZViyvuHdY
iuFLXoj/xDQZq8xumAsJbeIExsc9DCyL9kNUzb0JIYFZeBgoDw4TxBgws6waOfut
MXWiU1weBlDO9TyI1MDJe54Tz75zB7Qk4WyK0DpuJVojk0L/DacIdUiCTGJ0paAF
2HObC4DkD4afz+By9F66j+jM6/prC53VujICDdP5iZBHSGzVQWFSa0CiD/NCd8OY
cWIfC3ssoXcMy037iZaXQ9jDlOqAqNsXkFi4gvL+GC4flZUrxJY2A8mmejl8hZ+u
9xMod8pgp1QsPnjBvN2ojqJyqj1V27YaloeB1xNFTYl2kAO6Df1bmj/UhS4ptevD
8gm/4RPiL8XWRnkWqxoy8JhLmNkYdTlGOqt1xnI9xnYFw6MlGTWOgBxGVXhPp504
pKF7PXMb9aOE+jYY5CdYEongy5KpRasvwCZWLX7L6rF0bMXfcaHIXWzAYDAAnLA4
lHQDEkJDN1HMiiN+io+IlAXTCwBHYm57LjtOvqJIdvXUXELzHcsIXTWu3dhMEDjU
L4iSrVpCyju3qJo69xOYrKq9fIfZS68TTOZy/R64pHxZhWP4RKkcj1nMqdr+/vfY
vTIThBmWsE6hEQ2KAR2JnKVKshPTNEFgw50QQgD5kp5MeJajoOg0LCPJoByrp5xM
7nBQSLdaGxbEwpjMqsj6n6eCBtP1Yhz+4nXWZXGeqTYDSsxrIoIcp9yNpzss4sR+
Ht/9YFD4aXuF+xSm0deoC+CFOzHNhCTpzamU4KkM2USFKSqmcnoNcHrpN87xxvu5
kQt7zu6kvFsZZBtVdYuuEVVJqYNDxQfrhBpDaD3OyEP0d/eCOZdcsHv5Y8QTUDf+
7SStTbOgvHRd0VxBR1zZSWRc7TP0+JTGq1HMXt19biIgp74UFcz5NetJs7QZpZi8
xqavYYHhP5SrvTehfhP6lJie8ums7zkZbk2QkuhDPvRFCU1kVPlUilCkgYKfMCay
qZrthUqskLLsxiGC9JUYKBKNmSzjKuAtXV9fK2Ps+LdNZYLCAL97TG7JHFSQKIzo
KSm1pEL8FeCx33cNu/j+dnvRiR+jo09xpPL1mYSYoZGWbfYKLBWpzSqT5TOI1iug
4L3cO55JA3AHAoKqhdNI4tTIKqKEID8gl3SapjCao0kkDhp+EIS9QQFplgs7v4uh
vya8fnEVnBgxSRUbeq1JYfrqJKWa9ZfFjy53nhTDE9Da5uFnm2x81Tb3UYXZM03v
UGtUNYhAebdKr3MRkZlVNadiWuiT4IOTPS2nY1Up8u4jhuHhy6aPRCVrK6bTtw9L
TiDmMqVYdS5REPYfid8IH//sK7jJfVcDiUl0JSjXWqqTdCjc4wSeoEzI1olGavkE
kX1483tTEoRanmei6vSgVqkmlJhUA9uWSt52NDfO374xWfsKseH6v1micXkUGS2D
YLgrT/liAsx6JfOwfyswZkM2cwuPJnhTQzrSbPmCySnp6JPEWe87zjCwZkUmKVyN
FHXIOhctKmyTZEpJomTHLJvRq9C/aPiI0WPzkvDEvFGzAUl9QOxDO+R6CMXRftBt
pxTrE0JedVcBe5qMZIZ/QgouUEQLDbLiR93u5iOqFahUYrO1cqx0DBbTjk1ml67y
PlOVyM1owDYxD+R81cR3dbNm6eB/FPvjr/5nCFh7ubgMcFb6GQcLKHmxi05KU7IB
HjLTyWXShBVldzuP+dEuYYOLgqHKefXiwvh86XuF9eFRbiPBXZJ14fH6VcKRzsC1
KB8NGf7sCvnDJE6RpGcVzfaAunVhsE3FB8425pv0U5Ha2nG3Hw3aKn16b3a0NBc1
pjdRAuKL71V6L1JV0TO3SuEZK8+BwCxmuqYO9vpFdMhn3Luro5zJ4nywbXRsszOU
mWDqOZdmsV0TiSPXJQ6CMePUhARM76sDRVJfyh0XA+Cw7BLYmfYSDkyb4WQszp15
b/TQQoKyTBprOUAOX/VNKvriYqkpIBkXOPkx0QqiC62LQcdQ08PjnTbjgNyzUXsI
csz3Iu5K0pzwT/+OxCN6Y6Q55QwzFMfJvlIldAKZ9cViRewl621CO2Yk/sIxgjs/
8EqQQA+Tu6QKfJH5LMXNdUjEL6q9ugBKBGmuF2DdZ4cNseEOAhDWSmItm9CQ9MIr
icU8EA9ekjBXuyPy4pr5pQdDvdMMCxRkKu4iRYtfE7KbuZGR3ltZGilgSv4RnqlY
aTgdHFa9iccNolbDWKQr2oWWT4kVh9geFYRy9ZFBE7q2Pmd3cI8cqcDfve0LQAa5
2sKjyMNPUmTLnIu/3Gvu1s0exeS/1TG66Y0t5+h1gTT65FAwcIN4w3BRipfv5jqs
C8E5G5+Bp5K33f0id0fdbM48UmoPcqMj6mv7LHnBwbS8w693W37ciqrpzqHejx38
8/cvfRtXITgiX93AqkqWH7IqwO4FdICwATqLJ60r5zGwfZp4wc/MBfcT8P77q2jw
wxeKZ5tPJIt89brSbOBEAgmjT6BpWaMwaybNrvrkM6OARYjPewRBW6uOcJjLqPGx
6XHwy7n64SSgIST4Kt02YX/Qb8XLanKWkSgEMqFw/A9iLTI5xwpxejdk45vz9aQY
rvsYZipnz1TfO9CyWyLo0ZQSvFQHULNbYjYuIbozEBFrNPqwIaIAceCn2VpcsXzp
J4SMXDdJAys+gKbD6imaWPNLLGff/y25y8S2aAx3Zxk0FpUacz7Mv9LAlTCHFnvB
qxZ4eieDvBVMMEtFCxpBPxsYTwPGzZ2Y1s56+5IDpJ9Ioo8pG6fO3QJbpmv11ZOM
Wk7HFjsBmMuUBUOzQv5+RAPCQ2xA+cjEAKHa/K1rg4d3z/d+SFzaQedYykrg5Bt7
DMDaEeCqxIxjzr65AuPZCACluL2msgUAIdxpoTWXw0xmwBlH4P1yAWxO4tfO2Ge/
/xiWyc7U7zPXS19gO9h+VlL+tDK33mAXIURM3anbfEZiCggLczNgV0uabGjBRp+J
rgckBYqJrCkuEHMDK7QElXoze/lmmh51yHsXvlnyCZNgO5gr11GnTHdgBQKCZj7x
yM7rGpHsMluM8tATHY+OwGM3s0+Knj+rFajqMP5kHJsDPuNC0ZdQhAjf9U1auh/K
Xv/POooNKtog8ak9q0LRUDXbL2amwUD3/BPoFL84eQeJHTM2LeJ7kwb9cErqPWaA
LxagoKqOtvpWFCUv7yFZt5UNIK9sVRU1NV9E54mTLwdIv4VRe7d6Av9Ad3GrT3kC
XB+EorRcfBVQ6/EQbft7yJI+XExxb4W6VnV5I4spJ4uLKKAKQJbwWccbtnmLAwFT
wYjyrEM90io6GYDsVYGgW4dKQcmNeYocpASfrFcpzXg5xv3TenWisn7/PxyFp2yo
A4YoCi5algch54Gl0hca/tCwdFMlhufOX017OdRihBJ0fZvJKPtAgFQDDgGerQ4u
27AOKIQRC8+7457cBMTalXKd6smHZ3J+PNRKXDif0WTRSkNoxKzp8CfvgdgnUHDy
NpekjNzTEtpJNq6NQpaQTg4Yq6bsW5RuXYSAvI9p1umVcwsKZ6x9Pf1nzXjtoRIX
8aA01apFeyQHMbdg7Ef+N9T1oqIL6bXzG9XHT162AZmeCSVkv5HfUZ+4iSNlTTJn
Hwui0Zu//HLSosvSe3lxCI1++SBy5P1nXhn+GHMH3PND1XUg83DRNN8NIO7LAXOY
/oWiAycRdatbHJLRvLI3Tpny2+nJWk4sv0UfgRxL2gQuPQKfkGMnLGusLM/Cz6RQ
R3K5u+7NJco0pGHhNjsyA1hzYxrpcr9sGrMs9D1ZysF7CMrorozny8sA7TOA2SRB
ooxryqlqfptjUMe8SNTgEeKhl8YPPqgaEk9aZeXFIVt54KkXjNeCBqYYNnMAl5ER
NfALDI/GoL8ALAqVMH2e6bQDwFjV0FFt4f7eKrZKhw8FjH9TXdI4jvZBqJKh6FuV
oVLuznZm4hdy4lDsW4qflHpKwMy5YkxGmW6lbI/LZZcWaJPZsosZWSBrzvR4mSZF
PAh1Z6WzSQfXX+/2Td7aKnK0cz7QxQCnA9oNFYb2G5noYnzs7jw4tP2zFzevMm9J
U34kMvX1TRp/J4TwC5KK0oYLmcIEAjQck3pfgnqwkIcwjBiJ7sECkuPVQ7gP+as6
TqD82sNRNI9pGpnOUZy0U3Sk+/tGAFQDWs/RG+zxzWNqQshllTuYocGSene5KDcL
zbyTVPvZsyBRGuo1AjKIAZhqhaAS0lYJlKLyDevOBMUe37Gak3XXlWxhLUirNX8I
rdex7979Yh/RRGo6AANJ+U++raaIdI85dnHXCgy3woexkCNgadqXNUpog1HRhpRD
KwZ7mLn+hD6ecp0xOYoY/1O4JhukfGwLlf8qEIUZMrrjYKjxTteyY4/q/vqiGIEu
d+C4vFDfrr+kiinjcN+quw+4q6rNZsITOMTIKTkJVGAnFnrkEAj3dcw8YHT2zqeB
8dW/R6zlA76C36ZkePPsgNxFHJ9Z8DglVsSW29dEF9QYxJNiQZgWcNUwwEWuh6hV
GZ2QYESRz9sipfcmzeYh02EuUTmap6sODxYJUl2UqfyliyCIwhGx+jIJjzWz0t13
8ui8HaTFHf/lX3VIJYOpvcJGOQqlDCmtoIcwXsFEt8/4K7EIj5ax0X6P+LJwMvX9
vD4caAt/AFTiJ9r+fcz8uDitDAXEpvITqeECkRGq3HbUG0LtgFVhVwC4iG1wN+oN
5GuIDVShRvos2YQsyypfeVVBsMtvHLKBf2ySHAxX5Upgk0kLUl4LzyQ2a1COd+1d
6/N9LXFQV1K2w27jVkTYaz+33tb3k4+XArGUKAguLo9R4tcdPSkS5ssaOMOdBZ7f
IfphSFQVm/pI3Oct275QPM8IZFPpHBWbKSNs2HvoCV9l0M3403vdthBPbTxFeBBU
I1sySImp20MIguPXE62eVdYw2TXHywTBmh6iy6Z0x3OmcZv7U/BcKEpPV/Leug5O
q8EcMMKIQRwYezRV9uW9oxOuUgVM7LDvh9pOSmknVPPoqgQV2eVqFte22X1mV4JO
KfgkS9t7Jbhj3Ys3sRd/rC3RwdR/MPQ050Xvzsu/msNJC0YyP9Ypj+lO4WKSacCI
nvaizKd5vCxJLpf9UpV1OPCKnOsoW4Tc6xjoARLwM1+JsmdRqcb9ufqMBSumd+VZ
3Z6xKPK0/2y3kmnmhBV9eJe4zNZXRf+pBZaviUaPAldfct6gEtr4cNH164x3GVsK
n0ksMmB9RbERCW9ETUqpkEmBknjFE3/faqrdFfew7znXdu8yB5V4RaDTmoBrBb21
D3Fjsw/mSZZda54/vcq28+R8ZXg+uenld+08DI3l6FQxIl26WtdmAWqz4nS2Vqww
Nq+ufGteu/cW5AyjaUsJt5KrOO2TfEvePhv0ujw3piE1ygj4NGJDTfd9qpM2Qi+4
9rADNRHClY1pXTCu9UCsUci0XTj8lBBA0j3xirm7w0LZjQGkYkibzaiU76vzPJqd
VlXITXcnchEq8ULKHSpwe4HR/vJFsvw0kCfsgftKJL7Qr244hZSE/CZBvPuQGdlB
RiRIe5KJVytox03rHACiTKlX0Qd7vXS81QoxGVl77cGZnmVUAZ/ZmA5sr+dsRleK
KBsZM95t4Lg5Esr9PrLOHvkP6xVO/8Jq0gexwiljvNclxUeSP6btMUbblvKz8QlQ
XySghr6xbhqgEZmjgymQkPkfpol77qR5Hfx2CXQ/6tqIJSK622Qs0/hxrV9lUPz5
R8MTJA9kzUwJYDDQ/bidijpLdULxehvW5ylZpCbElRaMD5TfPKF7jE6MLs9YMh5r
/nRwgfXDuxtqlgp4o4GQNymEb40ItkRMvBp0PTK8LNfwYuqApFHb7ojQxI15j0ZR
dxM196YjUIgZrHpE0q80PLqB5rHN0xGfIkBAAcaWsCrJn++Q1ujyJVrtwfe21k9v
DkcE5QNg+Smxp8fLGqVvgSr2mFQHzuiFuh0WAeze5mgke32QAAhePC9SEkRrvXv2
/4Q5SlKi1XXRSgWET8lTzvwUPA/WOSp32gfu/x6feXC50mB8hMXCqCKKxbU3U/+x
V91G91a3uS09ww6TBahtfYNTM80iA6LswX59mXuCsGNmAFB/dj6MGU+enFVZ4U0D
dtABf3l/avOFHnwJRTh3rfAaNKVGh8pIh4JkATiL8tN8+Yx8990XcXPy9CKkDR4z
y3EWCoJZ8FNGd5yEyG7aT2jPEymeFVeo/2t1FbKLc7aF/PANzZE/dU2ETpXqe+7T
k/fcMDjb8OQ2K/gOVdbwRDE8KUHEn5+jUTplbN6MSDOOLdAKHkbQ2MIp9Zxe7293
MXVPOZjohMAMUU3loec3yk9Dc4a4gnuImpXMau5Fau90WIHYxf181PvGzAEkGrKt
VbD7TirNXGP0a1/9+9l8O06awxhP4kZEnjlQo2Q42A+IO5BJ/p82pFGmwCsRJ2ik
9TYBCWBq2Ue7lASn34/JnntzKNc8IWpu/pb8k2jvxs54aalI53fWPIyVDeL6YmQ3
sSbn2T7nOSRewHf7e7n8/cBtIrrIyjtIrnXhHMDxSidjC94o2C00fYF480KNzXxM
ASrIeAi7Kr0vB5Fu99ZA0R1fBZlGAlXk3uLsGIHeZXAnGV9yCUQoHSFez0G0ZNYT
GmqoBw7P9n1cVvvi9l4hnUNPUThUzDTkrYc3VTRyLKUPsMw6qlEW6C4IPhE/F9cU
4HzA45FztbnwN/89bLJpaLEJFOVrg3j/JgeNOetNA3Hye8M9xn9PgfZ6sdZ4VM6k
nM+PXU2M7lqHUky+mVLUhS6JyR/6lyFmv5qv6+OFh7sMmbfNfF4Tpt7KFzrdTt4s
6q5A9HAP17gyPCeicnaKpGGO3ROJQoKCdjmFyB/DXiLgYgN1hj1SKBJoIOt+5muj
cIhAqdTuJ4MOXFqmjJ7NcN64skPndJhdUwSS8+qbviVcrTzlMycWuflJz/HwQI0A
trpbtYgskr14ZooMxUuz2x+mtJdT+wjJLas0m/4AkMJuriGyYzC6FRyAQEwjlUZk
i36XlT8+8uVV0wqfqb0Jr384YFiWeDDcI8scslAcVXh70htygg8TGk0JVDgb5tEI
pplJAnUgs3NEOdCsqdt3O7SXKuUIEgVi2OFjAlGbBj9/8pDdoC+YipsNgxHZLnGq
C+ms5BhdLXegSbRZTC8ZpnWAZyHGzs/ev4k9WDv9Bzz7XdPO3tlAqUatUhuYKbbp
Yu9elm9ntLkTh578ZPeL3TNqlzZ/2HiWQQM4oJD1sL4XaWT94sgUtKLAGqRv/Upv
UWnLeYcvJhP2XzXRH00a/8uPgSW4jllQp6FSGUInnYDqA/Z824Kuszm5mTXBl9wm
Rp+hDTZbOlJerrMx2hGQRVfr7eEk1IiZl2+XaBXtJLBr/e52DMc+tscI33qJY3TT
oAfD+hTjwePAJxH7se7zDzofwJxCHiXtzTjQqMWG5Bw+mFXK8jRbkb/b/0936CeH
9+Lh4FCtTckkWgF47CkZi/DKW0bASzKeAo2lPKCJJTsxPTLued1UQJ70GLp/62sN
JoD7NVOiVi3Fjr1S2ZxI/o6zBK2GSvAi8RdJqGSjYCpC0BN2T+Bmb7wt6BtjcweG
8QnDxWDuIff3LLYvpF17cbFh179Deq51q320XH2n7zrOlsF0VTudtZlPokSGgh4+
7v/kCxOvdiuKZMqJ8sbVgbL+wSyr3hl9LjWrXOF1UncQU1sL7FiGFcf7y6VgD8j6
c7kcQZB7sinTbjpuzMgSxxMMRHXbUb9SC9m2upO413iBZiqX3wjspDpCa9+2D9Gf
hyyoYI4z7NHgjj5xEAurDxzRLbtV5TUzPoQOvZasLAyldSeJ/z334ot4Nn3t0ogn
fkxXAzhdXP0QMvHVfIQrFLQDnbTNqLIiBTX2z/xhmjUBWCTAHbDsTpKJGUpy7oeT
rtWKlJ9Ei83oKPHhYd+nhlI9e5b0cf7wTmBYVuI66zYievxTTblBunlAjgkHVSRV
bWgZHGWYiSEwqb4USrsW/ae2VSsNSKtlYd9ktOWBkSQmKnZ30OhCUHbaO8DfFDVF
xRL9dUXmAvNCJGKuF3t3LghjJKU0kPbZmTW91f2arImEACmK8pqVr3fkDXUX1I49
9oVFlF/D/bNc2EuEsH8B6CqTdo5riyk+Ma9HQqP53McYFpOW9+2OKbH8+G85rFOO
aw3+mGCIgg1r/Hmv6PJjyNPk4qBr+78gWAGS/CyQZNIlOP74ljFUz6pPmtBMSpE+
Hi2BKVlQEhiS/V3J7C24pMvWmaq40F9CUP2qhZxN4cEvZHqs3xY8zuMp2aa0U2df
a7ni1HQxIz6b5zV940TnWe6/3gOCghSPgjSAFNM2QvWI9V6Kvebq9sKDgcQScJdU
eLTV4STbi/GqJDm+7rHQ4wKH4uR1CfjNPggQ0ZoXyzLnKoSTw+LIEi5bvMhv9toL
IXbfwD+7X1KvcHu7dytewCo5ZK/MzXoKdeipRdqctJ2fQjKziKU+CD2CM9cfqOL1
H8l8SkVlUyhGM8zHtDFfQ8F/TJ9pcMRcoGwuYa9Ona1jtH6YfuHpmz6rbypVX1P6
R7qhiSikicBP0eJv8BODSIpwubvWETywV7NXhZBkboP+Brj0wIBogbLtvG6vV3md
+IX3yQ76I52+TsYyJrYjeJtgcyiSPY0exjk/dH67Fd4lAvBoQG3cAqnb2B6tyJtZ
Z+by+nbip2hfwtNabNYOvm+9/wmJftCUwuGBkKllvXmKweGMcQc5hLKni5TlLyf+
MrLyeYhvhlhdIOJplK7D7Ub7+HvHKKXXKsAjYS6aTkDvDM+OB8G+TQbmHgyJW8iA
wFzEnVShkT1wdgciT9trLRbcJKRByjWv1Os/MpzQGewTFMHG/fB5dQkvO1IBpIBa
0riQ3HW/KTKbQHJrliNyH0j9ANzAR3VSonNkPkGhxNZted+aIMamvgVIRD8ewUjo
mWgZL6bppISEm2PldkQYWfwpE+Ol9ZefbZtcbOE5UR42p6uDgi5TroP4+miZfbSp
sGl89dhralDcShUT7AlWeKS1TtP6RlWxdHIqV5qnwZLvhEeBQJySHHe9s5oFsZDZ
gUS667tcVadaaqRG/BvCvXmC1LCZvGRXrB9RpIUTjM45jLLggmq19TiZknmT6rwC
wkKcHSR8frlVAiA2CUOOF+oKiz3kpTODkRWTqsldzbFG2ktkX3iU76uaDL2gBvSe
yVxKxIUy4CNoT8q97uZYCGai5Xs5tTssFKDWIq+GJgzdJMrhKQzeS5Hv2u4PmM04
UwYJEEhIS48ZHUGj+6i0DNKaEN1susiUYXPtgYwZ/boognshZZh/T555SfBEI5rL
607CbWvAeCWQiYqf1Pd0aTl7HOc6b8cSOxBdJcTLlM/VQOkqOTSd27PCNtdpEsiC
h/XdnAs7fDUbXYNZtcEltYtT5BK2F7xE+x5mazm22FgR877nk5WAe6X+5UM7S8XH
rXMfFDYBVGhHNw0+56dZilnKHROJIJ+gxC1CH2tIr19j4QYDcH181TVVmKYolJez
2AicE5Eu21zFNBY/sOMTcMhOI3FUHcQH8Y7j18o2h7Bj9bMcypppZBX2OslBHl38
u0OhqKlsPXXw/EPi/S9J6WSyLNkhxEsi4we6gJKq8NjJD3GKt4HC54o8u00RgUVw
gE+mhmqlwtYcow53PrZiWhodgZOH8qXdj7LVh9LDhlnIBQaO3Dq/PBzhsruNA4pG
d+E69g1RqkjVdnsPpg1Ggx1EzzITxaMY0MvU9oAXkAzA+WJ5PmiJsxNw0sEjsdaO
E+pOS5+rRYnjp2vkn5x9uHUxq6iLo7USq7ip6RaAtme+JWz8RDweuJZcgV+xQhJj
Cl63z6McEpl5BqspnjqLcOn/4WhIzkqi7bYY739cxTUKYXmJkzD+THsqB6LLExvr
P1fe25WlVwesK6Xd7QaVKhM0Kl9M7vCgnf3J6fCc8h1MWdhIiv9xCS2uZ5CnHCfp
cZTd1KaxGF04D3tBLH9ylC1pf26JN8M+4Y59oB+vAWt/BvaXJY6OpYoqiXIY2fUG
BmyOCUv66dzL2NkwS7O1iQXoEsB9ryxAgTv8TDED6DqVjqNGruNGM55aKOsJkvx2
k8EBeHYCUMuQI9EV1+28CQLbH4TbkYby8/tLMYlvruv9pXBVUSTcFKuPs971WgtS
ZIsbFQ9Rqho4XT17o0Sb0EIg7O208TPHVpOpFF7pw7RXHwzec0ZPFxGNdVdh0qLQ
xgRSwOMvmJUoaXbEn1pV2cCy2esRx90KGKlaxxulHk77vtt/+sH5p1UvCagSoWLV
3NrEXM9lpDiNB6mpOtePMgIkmLOiI2ega5at6pgXEGVcLU2i00McCYCRAOpmZreu
rBDqYtl3Ok0Ws1GTSn0kq3wifhzbTnOpxQg7kldCmM2fW58RoNIPZZFAdVk+AIlS
h9qoM0/degbhpW0lB5tMeNLgvQMItc+teqjK8ya+Ghvd7gMGeZP3wHs7P+kIxr1a
RAjNxur8YLojWYWCJpBBhHRglAJzmGTmZCoVr6nAa3eBLVGN0xQseqCIu3U5Rj4q
JJtgEx13cbIW0G48+as2QphAJS0qkyZhnT3ItSY1RgItuvGPrXVY3oalMzOYy1s2
DBuuFKuFb/ehrHpCgnrzloKohV8HzIhfAkrM+XPZlsZjm1A84zPK9GdN97bM70Xj
xVfsAlu00DUYSc8ebrluoB6/QITouZTIUq3bJhe6eUtB2z8VWgS4DblqRj9wOmAQ
NO/Cj/zx7MxrSxnOveMavPaAydmnG3shSsgxTc9a5AsdyqVTYV5AV79EffWbPM4Q
XEM5LIL9MNYMeNxwjaMnIAw2CanUi9BbYcWH9wt7avFHYvYugemow6oyfWh/k18s
mT9b1sj/46dPmOyotLHe2/LQjtV4D+id32zmhHcFEyJey1/7Md3OmQIUXxC77Zvn
bxeMki7E4TQGuyOO/epPk5hS5MbsOi5DhS3/q7DWBwYx7R5/aWbdVJWzkRjJkCLT
s3iWYh1/bKPKVdJOBI3NtdaVhGIWkt2291b230P4dnKL7bgyeCtT/zhff+7Vop/L
sUkEFhUHHoVxJwF4Smp7MegYk+RlNjP2/QTODntGf776Xuv4OAmX6dCR167bP3WR
nCvZHKS/lnjT2NTrGfI2NNWhWrfYSBzD/7i9mRz5IU6Q0wKG2Ew4SAeNAW9Cky6W
FScpSGbopN6AbBpCqquANisUNUXLb9PX9wPHNmHfRKUi0HZQpQJGAgGmE22kDxrp
nPEcdgJ1j/xyudyiv6JEiGgGuZ9TN4PFGwiugKjojjWX7rvRLu38KGiBOEm+8K+A
Ijh24RIeRWTXtfDejYpPFkpPluUJOnlYbYYEtxJpBsrq/oOOOWQgSNdly9pxoQaO
YtL8FK/nred8pTGpreDC3+YRHjBjANQEcOICNY6mx5s+4IMvLxt9c/CXHWsYO4Ui
8szc/hGeeCAaBB+xSKXjh5Py4OFVJzq0EcDiJrsni2PCQZvpowhdBOaZJlmdEJWU
K+QIr+AHExAp+BjiFG8IsUQXwJXM+ys2ygptiC8tcSitT9EpzWuHngcsDp13y/WR
zTEvKrzk84eoa2iHaH1wwjAITPQWpK+YSxUSdigsiy6O1nKlYSzjRRxnoI59eHby
b3FPj7CncJBTcwZfO6qLOCTJtvlrO/z33oYc1RmjAl2wvH1vSNAxGZq0XXsKjw3V
c67FbHTYfE/klrlpQjpIvvSlGFSvlgyzxzkFDKiqbzRPWs1dczPWL8eN1wf45YoK
FX0mbpxEeAGDjHhO1c6aRhqK3myI6GYFfP968NZH9V3DRnp86ltiDaTD+QBQlwcm
uG6X+cElidBJNHv/e9+vD+Z5kzGxFlZesr+nPuOdp34GcRcAoiqeyr9XwLf0KcDs
/ZUh/vnP2+lj2wLLS6jPbQrJz1GkhoV5ByJdOtJOjLId5UslhH+MtTlfUSnsASqI
5Aea2C6sX4JT/fbNExPVQuegZJ6E1z7hjwDZ/B4raTNY+HlquuIYmZ7ICjzFuLHN
Z0TFMRofOrSZKoiJWy8R8+Q2IGF6LXT7Wc08coj+jzv9SDIuyQQu6ncF0/Pftne4
y3Zb/hHVAGX88tVW9TYzG0rIrDngvOmYWXTwvHoJbEDIaD6bi8E539WhxuAX0z5Q
/rO3spLHGrr0rXyGF6GMowpx3lMvGDZzXNT7P1Rv3UnWiX/qiRVtE511Utyc65Oz
BHxogxsQb9Xv4tAmM/FPZ5rmdO/xphmwQ48RnP2y9jIMMXn3fFaipBonH0gzkE+e
SwQjvy7ewkOsJ7bDPGFeDKSePvpV/FTeYdnG0c7Mj6UEl1C1Sonj82fI+Q2wteYS
JmjgAcWE17WYXET/hJlhbOvHd+n0xVGwmjcfodWBXHrTKtvEKrkpapi/GbUqE78e
4PZNP6zxu8Y2q+g3b8EWhkc4AvcuhER4P+lBCkgRD8OAVWzs8vB9tw8oADPZuozN
vnlOXvRzkei/OlbHErC0PHNV4mdiIGkcwV8P5UbNk2uFfBTq4WYcoTmTL6g0CEH5
8Ss7C5lnYRpjvVJ6BZkA730/84MSy2frRvw0/hSBfUKHq13RaIwjd8RB4QPNkRK0
Vy0E8VM3oQ8utJQUOLOxJwM7m0gMHBfX7xAsF06TuuM5c+UCC0phnwKx8wCXfmyq
tFSswEL4/nbUZbXcUeqCFlM4spYTCZyI3uRIAnZtbUbaY7hrmI+oS0i1s0aC/kiA
Ivhsh7msohI2GJp6XJ0833j2oyCyJU4di5Z/9xFASk565bak8WPSeEIyUjSY9zhm
clCK3qGW6ecOEUDOWIPfqmtlsKaDCngU2dgnpQ6+2ennidC03nV7Vk/suKrZNx6U
I3oGed1ecxeB1B1FQ6+Wc0UUzpWmK91C2DCJjExfmr+mY7OTteXFNH9SNhJCEfWW
8YaQF59qsf9+s3hqWz1Snj5x8D0t1XcfSFOK8XjqrqQJeVItvxcPjQxGJG3iY6v+
XxA02XBbMWDG0VlC/lv9LWbDCvffcTjPL6M/5ERCBFw+jPzzIYrwa6J6v+NtqPjt
KNREAcP08bUoOIYRpxSEMYkkJxX7Ly2s9xFlsxYR8UBBVJ/u4gB6JD2AIeOm9Zp9
kFJLgurhdWslW9zjrWxcUtDBv4F/DqhNH/ppz28oNG0VOCGLZuyaPRzs8Htkw2XW
YPUXFk3ELVthrv7XYjNwPQfH0FvBf3eP1nO09f/CtNrXS/B2mFXZrTfVm9xtDfEj
nuSszYRHInE2fDv6VennU5fzArmGRg3snrffm+g0IP99+aEaSq7b3vcaHC+5tCCM
JfDBttygzIqWAGgNpW3970lB16YUXj1twjhI6egp+mNOVHM9fpIc74f1pZs9lYZH
UwIkLHI9SFsG7kd/lgBjvgUt9P4VO6ZHJ8/L/Ibg5YcEI8Ev9KL4Xx+ToKNbt9LT
uR6NboakfTvunaVPZavS3zFKPwuuPuUYUbHW71BYP3YF0NGOmnZCqce9MxFFJRkZ
DhFS/PrlxOfTHbftEXggTIZKZZih6VM1Vo5ZfHrnbPJPMq6OUEKnbYf5jAzvHGpm
x79Un27dM+mnT6Da+DmycDgkRSmnFekf3rRd50yxeZ8muptwAtVP7N0aBFdaqvEO
2xolfOt0L1JeuQNCvQEHCRB13NOOaS+tJfVIACJdV182nztHxUQtZMfC8o7ECDlq
lARmuT+zPRh/cgtM2OOIG5Ex9dKwfvMb3iv40Juy0YHTzt+R+ikneRhP4FMpY2Om
MJSJ42lvuFoEj9eCg6M4jol49gV78MzQNwIREGzwKQ1ouVIXe9KumpYA7C5Cd7u4
N+VibXZBGIHbHHj+ZapXeEdKFgKZV0s1xuMooKhlS4AtRsVP4WM4SuupkNXg3JHA
q8+NIPj+hGeZLnl7AKIcnYwf8fveU/Y8I5g8zfmIEblM2qA7uZPq207C/33KEBiZ
WdxFoNv1NDRereThtECU0tXJ4B644RDNneGMqPA9d91JnxAvqgGN0q2nMTqJQzdU
s8Oaae23h5TD/CYwsKtzWu0JUawi9hl0a4zXNX3f4QABV9mxiBbym/QST/6QahJP
C2NMbwH4/Jr6iKx0zc4UUikhYQZB4D1A8wgpQp/gJDzJ+agzklRwoHfyc3RDpNO2
Mby+hjvxTKZ+/pBNB4Jk/nxgrOnun0CDynEYvpi6JxhFEURyil47hgnKyvUMYunz
XWKICgO2MSiFcLWy2LeoplRyaiWBKNGmWWBXLxENhmkHEv/HzUjMvTjyZvMMRAFG
4mjnlyPgMMekcfRIQhoc8z7u4G6pFYf4EjatqaCeeMkIuOSI9TrNuakJqHZ4SM3q
umAusXUpoOGcw9FCuro8hHW4QrZLhwN8YxpXDdetacMbepg9MF1Xp4s1jm5uIKTZ
Ja/HXUW1U8N0FvjZvl3B4rChgzlc5XpzNATOnIO/i4nPUdxAEr0UyaftLt4FW39k
IEnfsR889x6gvBFeifN23+uQ7i3PQUOMgAB8STnwhZP8YFbxc9Ie58KytD6JcXaS
YSu01O/m+YwbCXmvp77ibK6CIo9o//gRrLc4gHoVVOTYcOavIxKtAhVcBdEEb830
wFwpykpGgmP83azHZtHecEfTf6siukRvlKICQm8y/Hu6x17waMcdjwh0LFo3pU50
6xkduVo23KbTbShO9r/9C/Hdvvrl+CyDuVhad4+txVbeayFEQvDNdf3w4tTSgkUV
+gl+VYW0rLUxc+88iXsMHePXki73csW8dq4pu57sRPokcAMDgTcwIIGOXlQC7lYE
FrXs84g0MC1eMTUR43yEYIYe/QJlM7CKUNEEljOHy0sf2EQGekctv1dJ1z/x6Sgu
swa/4t411RSsw/ljjCx61Zx43T4Y7Vb4X0edgyuwW9EwRBsxnLLJ5exGJBTeT2UF
X2+7XoyOFEPF0q+WyzV3sGIDEYws+YF8iCJY6Qrc1GUnNRuy1miYv7bcvRkYH7um
KBMmMx5QX5uH1uhFnfFRuv22tTUJ+9kgmdTT2glNafLAUkvmv/WMgYY11Uk6Aa0v
dhi7ptLsBbd8cJFnZnVnrXuhPwXLsiKaCZpDvNkMKKWdHpxS5iMfpFxKs37I6oWe
VvroBrfhA7I0QXKN4ok495FK1x9ceXrJihdHUZVoe03/tYAoktgnxxvAtK7nEIGO
RZibHGLqdO27wWqUKVyFFr/zDaLmcSR3BvqxDq2wH9SYU9R1N1jOk9d9A5YTIphp
VBAgpwY8dyT2zwmcfjELRTkDMedqZdqGX8NK4lIBalzNLx9lR3S1re5b2XeQz4Ul
4+VfEe9Eu+L86fAcwTNYX3wLTyszCPa4xc12NkElcklkN8EQyz8vcedA5PMTQAQ2
KuVwATupWirD0KISyNZt1hvChPRLL0R8ycGK5AWCo1nBHcdZsz21Bvn2T7wlzckT
LXtGLX2qQ3JBXYOp9TteBC84UeiLN6miDrOeS8AyLGM9sPS65k6DV7G+VMrv4TVm
0D/+meMuHk/XrDNusN5/fF87malWFxEbzB6WmGLyFxM9JPNhYE2wydufxU21WEoZ
jedxfQ88UpKw25YIhCijpyocIYdvtzCAT5lO6s98C+/LmjuMLe02BCnCefP3Q/ai
guYtEJj//l4RUJaFtbzBsQvfazqYno12aroQXzW6yQzBDubDM3GKrrWGeCiX44sb
roLNJ/REXMXdoC+HnlesTym1CWxfDSLV6RipzJTRbPq9FlON8qo4NPoW9QvmUDKx
djNoYN3mzc2p0N4ZI2QBZgHnbgG2qkEPuhFpIQK1kw4A7tOpql7iopQEc3fqHSNG
xp3RtcoR2Ko2z8X8CNkjF+jXEmN8dJB5QnM+KXVvExH/en10DkX59basRiVJjFDz
iivQXggEQ5xllULvmtKv7N+EvS65GewWafIwSzMHVHu1ACdowAF6Xvq2PcM+DdIJ
n/DOfOSqMhRJY2MkxZHTMFjPMfYM+H/dW35dxhQLLw/6RZCk5zLHn7nEnvYHsbCi
Bu3xyc79Hxu3zkMHUoQ0RlJImI/IRYsfxADNztVEWyyu1sd6KIPsZnwAomO+A91k
E+QhNy4u8HWmMXzhb4XEiZCM8g/vzg/SLNNyfxpMXU4pfwQs6fvJ5F0dVNc4F4pW
bWeD92tfw9yGx2OWWUBoWh/fdS5j7Ok+BR1cn23M4UTvLTzCcsuHnAdQFDwzmA95
SVpGjdzC00vZG4p4XwWaiaAFzFbaQE34e9K3O8m1jRJrJfLwE7csBFyxFSQp2mUy
84rC53AarVdvp3JDpUZPTU6xeasSzMluKZP5kZIWDVhNLBjA8mI1DdtTw5vYVyVy
BMmc5aUFiBqmAgxzFvsFwZEdMDmnmigle9ywPKBBvYKweAlOLbYEozos0O1sM4wa
JMIy0r6hxoVqNFniSKIlsT8dQWDPAtYYdpPVxpg1AOVm8zA6fphNHD0mXF4/AxTV
heXv5gWKhNoxBeX2BhozHRm6eXl9NCp4oSQXAMXoehP3Mn9PKllx+BQ9bla6l4tJ
HPXTEG55rRQM6O8/Z54nnFvVJK8DFuDmbugbeSBM5YFKOpw/XxJzzVvcQG3iyr1l
upGzQYtoOm+ApVB74v7KVKh1lyoNItj+n8JcnLtGpMM+YnnBbCd8jNjP9dBjxCQ+
qbGI+5s6WkWc+hUoKIlxENZYWGG3NO9E/x+c9Jufrj+/jmsD0/yOq8irUk/wetQ7
mwNL3M8U7GI7KT6Nx1UZYwpa/eXdOagMKplvBqrC/D9RnUIIXxFFq0fwLSDzR5Ty
FPpiWROQyHCunKL9/s3fvFtD3ev1tsSo1I0WSnnFBMXEvn9ubPpXMKWV5Urk4y1q
YrDoo0CZsZzG4pw3ZeR3zFzBWA516Re9fU1eiCDQuXKtoT6tIq29KxC3RNzy9wuN
PJZpVKQwTNhPs0l17yvAWzeIkShWNR7ShIpTJOzpn5XQHkDCjiV+3JHKNECKkNdB
+5ENC9kvj0uHQqVhqyeoSNgpf2V+dat8FNnHeLlfwL7fdU8PinPIGeXuEiRTaWJk
+1IVzcmlSEZ8vvXAteA+G3/aAkKkIFgXknTHT2JIQoqLFncUmN8eqSth/kyOn0qa
RY1igD3fJcz3+9rJPD9gKdEF0RVJoOjyb3fXwksOmMe0fQvWcV0ntTuMO6iHbnfv
rs0AohjZQmuoLeOdYRkrT8IKIITVoDC89c+RWbm4+wvmn4/xRAUqyV2L4EXP/pEU
ppW5J8Wf+TX3sJdNmcVSkftANezBlgh6v8AfWNfZQuu84f3EjCYMHjCiMx2bTQ1x
5q/3/zCMCo5kGNVJ6UMfEbd4cZoxJ7JfoggUe+FCB6AddoVVJDegxWYzLCeye1cz
hlLbbo4zg2TrwyEgwT0f6a3U9V+XkB6fjQWNhHA1yEX2NTz5UGwnoyQVRxMW+mHD
aOHJY8Nt89ST6YBJERB7i3r5bOAmr9YLFvo+QcKjxB9MxhVl7Vl/1lmWQkvO5MtG
rQIGhafurgLEECSOs45yHUbp7VsfwSelqGkmaQEUchvthAHHNncSPq6MbsaVcxR5
BonLgx9rBYdicUV84Oc51qLSAtbYdGkk8DjgixFIFJ3qw1Lk/zQdTuhtx2W21wt9
GYbgwfVVLkEI9vBdlO/8Q8fdRkKuGNhDxvMGPZXydXRUhAJ2zbMnKbgYIk4e8GAe
NjLZUEtyoqZKTIiL9wZVE0mKpvipZjP4I83lknQRikifvRiooSTjRImDV+0uPNMT
QmboOP0R5alA5UVqWQZnbq/vsxptQubTnxgkkvo76GCdlEf9wopRRgCCYOHj33G0
F3RH0Bsada9T/ArFsQFQvxHOWJfT8+MZ+MYnUSwT3+3RshNbNb+B6ak3/1cu5RPG
YBW4xhwoFTwAoNfmOmenpwUd+svPK2soHyw91wi01l46XZp2nJTVXRqiz9yVU31s
JnzK7ILOSwKrhp9pcKaiM1rchMC2MKBcKOumMP/kPWbJOUghSEEYH2yB35iVgFYy
c5pp7/21mKJsBP34txnN29K6Qidl1pxvtvZDO7vWYtU92Pc3EoAWh+myXWhxlA5e
dqE59PzUI2ySLYWdmVJZQSJEgfcW5+Rg2PIBR/RJcpcuFk2Sn3f5xoja5YdOn6t8
/Sk35NtY4PgZuqQ5mPwVH4Asd1PMTHUa6Z+Rq48xlyes2+vKyBzoBu5RYE/rMy9O
g0ddnY6rN+mc3A2mha+/HdeLhR8s7clsMGQoUUlK7+5n0l3SCjU429deNAXe83YA
wtvI/CTNAbZ48VQYUTrsFmQcvY8dLZEk4+Ft3pocCImz9Znz/qN3I2aZItMnXSfD
DVtZoq9cqxwQ74IAmiq0WtnVolMxI8+wSXt72uerSYL2tEap7R0p6r2R+Mibb7ha
o43FPvx6XM9MlkU5rKuCcL14WYRxYz0je350BO51B2m7UUzcnbZjr1Rcz1sMy3Qm
qwAQ5PGK3jlH79QdhzjvI+iEX5n9+YPc8cci7JrMtcvfx6Ofq2pK8XMYXI7H4ZCs
fxtlB3vYhyk1btF5tTDUqZ59K74EECL+XCDFeR2imab2OaQzS7OQWpnWC3cSQgWs
Xy/qs99GOl0w6M8l2zKbP2ZkvM1KCs+N8ZqD3PZK+jfhsyl+LPA1eDFi1ptt9OLz
WfUGQ9QXkF2ddx2wFi4Y54Ga8FVck3nlJXM1g0iguHiDDHZpbwkUKCA4g/Hw1mMD
vRCTBFWx2/f6dOmkXZ7bvdwdFwRpRJ1YOGAPh46RNpTRoGiVRJV1Kyn3blgluyJd
6v9b0t0A+/acY50oXNFzjKj8hAZK5KJ1tp6ZpVYMrEhFrmvR//SnCBWA0USHQzeT
RdnSzDO9jaeuNN072YBB82028R+TbtGmjDf/u2uXcsKMbs9n5LZYf7zcMpwXmNSl
9RUjfyywC525/lrpjKzUSig3atsowbKlT750D0gDeVFrDZFFK6P1zZOrO0X4E6Zx
KCkjO38p8PwYAtJheNh1CfvpVmw7Ha1y3XZ/0f62p1zBtHQsBUNc/Z2X4D0JTqaV
ZXcag8CeIgqsuI+tgpOXr3hrU2auCNpP7OPyhym9EmNiKwr3CrNrTZI7mVZ1ZMCC
5itrfnTM+H1Nu67rZLakhaEu845fbd6FzPDQDC7rfowpjFWB8cG3kltwzcrdVaxA
6Vsg+oKt7CBOVmMp8eAREKvTLGiNHn55Y25TE5RX6PVWQCB+ui5+25Q+r1ILKAIZ
BZmCaV6T0srfla8AVUdMZHbtJFQTPlZMnAXZoH1VbY4Dlf5JLQIt/016uQoiynSC
ysQIJc06d3OJpy1/mMW1cQG7G4U9O8auSFoBIFw3XA7OnnoHAvT+BqjwXhB86jkc
6o1h3JMhzsUKvmseM5hki3fNVoih3vYk3V+J7iCgDtrJwHrfFVIjxX2N4cySHI8v
yI8nITprwmYGvL9Sd3vqEW9qWcBTshXw5WcI19cC4PccvcLfoEbdnYokc68asUws
GaiMnwQk0wM7uZyVxWJSmMIjI7hnd0JgixSfQnYOSglSA0mf9FMVusdv8mHLPMIX
WgD+p2SfKP83vUhxHgMEUr/vBSYVEMDVYEW4UGte1O7NYq+ID0FzA5sj9NYWESR/
YBJmT/4pNEwB1l0PTF+/a+YUNtxe154Cb12EpuGiv8LQZL9p7vpTGvUm99qsWxK6
9Y/dCDPaHK31hS3XXIatTsH9is4qBImLivZlGyCcBNI0Rg1Mfvv1dEPAIs2PLtMU
kwOSSnxqfWbr9KDar94alsFAJbN/pzzfxOQp6x6wUtQQCBLO7umu1/SNF+lH5XO8
4H54G4HqGOIswWb+1uSZiZ9MhSwlIRC2nJgwuOPC6q5wjFQKjljIA5HHlmcUP2UK
mBybnRxyFjBvO1WjnqPXOo8CPqr/UnATJmlQ4qSMerOhOoSqXHYQAWzccBUWVhQj
P7vaA0I2moRYH9QCbNgh+/X0BfYpH6CycBdMLP2SR1gQLMPXOhEuVlt6Om41sP3x
`protect END_PROTECTED
