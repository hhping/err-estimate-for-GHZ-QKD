`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LkWeRC39hQ7+ePhdes3uqtHvrrtUA+FYk1SmGGP1WU0usaimLGsoS2kJhfCiLobm
K2v+0dQM1zF3cIh74u5X1NTEpNKMoIFq9eiH2thwOcKWenibhY6v5Bj6GK6BFJR2
TgYXQsbCUVGyQ7ihjMSb9HnwLThXwmlJB/y9s9PZuM+7Ld6WEaRU8Q4oBWy4VvfK
78ejNEs3aZC24mH0hmnCNtHsgi5b0MNESSBamhaoiCgfLOCU0ZZkAHMfu1JV8A9E
1a8bDr6ONHyTLZ1MlXQjlwmEOsnzL92NuNrNAARfcLTXOff+mnyfLpu/I55YkMAE
MZilRRSSArbkJ3AAORfkh+lfMF+QAdvL9nPStcu7w8ap9wadWzVfuGS2EaQ+5iQG
hqUoUWCJ5NZ75xux7gJeL92iufsabGShQgnwyfWG7Pn924BWVUxbH3UXIjrq/No4
JK1GGvzkVfm9zoPQBn+ouRBUzZXamC/sO0oBv6AaGCT3dsAjki6kMB6fs7VA20ik
qgSjgo/Bjc+jKwg30X9AFZfSmS2EhdrKI7IaUe5LvhVAZTKmgp5qIKCqUxV0NqR0
1/k8xKPs8h5KhuXhakjFnbiWXWy+C/Jy8QyHEuESaedSTWWluz2LSrgcVQBPJRDY
X7jixacQw0/5mo5IBARZcLqaKSt3AqAt6ZWhijopfqegBvzdluf7tkODiLi9S8Ib
ydaSO7z/GssTCwNH4UJ6DykdK7dGA3jKJxHNA2xxdi9lhxtIvjsxnyxhvvLA+Zq8
4lOcFP83GLt3CixNypn1L7YL+agFaHwZHAYxGYNteEVWm0CiWMmSQqBulrImLBLH
MO1BnTohxo/B5FGYzEXZtrkrShgKGUrYBX1Vl3EmnaucQaw0jZ4mQbeOhcvP1UdX
+ZP+GcFpib7mgv4j+FPUtEdbe6t/Ofrh37HIiMndCXJP37pzE/zkZvym6mWY2fYS
ksHZqoln/tA0E8RQ4d7qa5JJDNcDp9SJuHwNULsXrwDU/XbSwQU7BksPJPAZyfcr
g7RGOZA/5rvXBrrDw+mOD0iedo3Z3PhM2tzzrdK94Eu3yusASqyF/rAvJ2GEBkA5
rvND1KCM0unJrijKfxd59Z5hD9xPQCs0xxPmx2rWqu3VJSqmjToewgUAki9d3fPU
A8n6rP+1mnxz9pg+2kbZ2U9hDuh0DTXltTW4ZjY4h+GWEPGj2ra1DZlqnCxKTBj1
slxhCNs52aLUFtVbqpvXWyyhNxOLn9UZleEcxD4ecv4I7zqwBWG8pEDfL899Haxw
kvQQjWVMovdHeWiG8aJlq5pXgOKDKX+XyjJI5ua0nNjluNa+ODTlLYDAiVUz4SHK
oGOI0LfeoMTx8J1k1prlE1cWBANf3l7XyM9MNzjwMXTp+PON32BFFfA4wdT8mKJd
b15PrlrxWyDinGNh0gTrQdch2+WdHtL7zt/x+O5F70MYUJ+Oog0IWsYrlvMqy4to
aTaXShRaKy9/YO3sEAWQ7tYhKD5l0JrSFijOpQWzLtdDd4IZuP7qA9sATSvn8TXE
dwGVgTC0VnW4lb9cn7bP9jVUVu6AutLq2h8JJCakGj/V453Gnmp4nMPX6KoIc8Cg
20GlWoR7upY+TsldLbzGZtzYPX5Wjf0zEQrI640KIqH/bKb0JxPhk7uLmv8O94f9
pbEgDpejf9HisCN5eO77Ezv36EJ6lLz4ib1wv0qzMEElF9N7etN8sjHah5P+C31O
8fcv2Iccbxg8EGlRdorngtRaVbmGbnezsccWjxw32wNo/c+CT0RJPEKU/Zog6569
xpTSEycfve2nUbWz5I3WopQuva+3MLSIccBbLYxDnL+r9/JbA3lOc29LP9uQptrg
lTymhTmQ1+Mgwb/u4sH+IuwrIiI5tcblYOOP4yeUwsccQOk+QMrvf91TetglvyC/
4wSr/d8BqBQaMzC1EA1rBuhecZQFv31PAhGHoVUGgNYa5LTyVkmhp+6w3vLVojdx
COO33KVkbVxp0VV4H0ITgOgpH/Bx+cTe6FuHrQbVHq61O/5i4GBz2xHzVlRLWoyf
UNdB+QD9FcbaGOUypgrB5dG7zdmByqc9GkjhKr6g/SY8uTCiwHNAo3cirMYGQXLa
uVmHzFSoGMVVPmnFDrk+eX1Pbz572YM84LeizSi232QwypBwW39ZIfw2/UXqzdBq
NAVCT4gTZm1zJwynqsutWEmxZjL7stdidMvwYSqsd2T+J8rf7/3su+PPtLan0CpM
QfpWjiwkKPZqp+rUY6Zb3jbv3APTihqy4jYwVD1T3jGKxXCNci8ib5qjgmCZE/6S
CI6jnTaDxF4yx/dBqOKv0W6nveq1Yqbzt4EjHzegbsYb1aznDzrh2ggZkmBM6BpB
m5C7vSuLGljydTJiekOIj1B5ucSKW23skeHw3MvQdD+ChsSz7QcG6FPYHWvV6CJ+
XWvnPbO04+stmxdHzwBS8Lmn+iMBx+2M59zOdb9Iuj5JDUhyXh6CDQENzwZI5Mkw
qdc/63eTCI7vwe9YU9WJL7+yPCxQxQ+M0EEN+jzIEbyFXTjnaYLohkcTGJyOcHxV
VcDys04+Cx4CxQAFQ4tqX3i9HEJAw8lmmi3CRy5SrYlJJiRGi9P0DkkpwXYHrKPD
d6HxY7HcpDP4jvBDqd1RmfIkiVYHAXSNAaPYnA1AlODr/pLCfk2Qi/c2C6AjhJAy
QpMHUYALGYfPftz/JmKuLY4xjgh9edh5KMaKQ+nEk7WvdeYyKf1DpG3k0a62Lilg
se5aF7/6gDQenwhaFymoyXOv72FjQ3TQhdcervTcX/8M+otvNoQVWQvQ6ZI2uO4i
IMsu5LEWwDIt3EbyofqY8WJcWrdN8iHj9KZsb50DJCWmJFLB76EQN0ZBbjjWRIff
4x0zS6t9OXu7lG2w5v3xjaQ7EBgzQsDPvBHE0qLLOqsbeKURs3Lbinof16sPKmCW
54d2w9u7GZl9hFzYXaOYSQgLltZ4ctcXUFitlxX6zstuzxCZfz1cPlQUDUSUNtAS
n4VDWAIchpzdYSYUQTbzAlZgnmef7Xz38IvTZtEu5ttc22oLqke4JZu2Oc3q6Qwi
Stiu8E/o92Szeym7XhG8aUYXrOTanEY5fm2yeaxcxoxmdWD9Y2FOwVsFJ1+IBFee
fFl3xg+8I63vlsU/lOuktsI42UPTL/nZydHbTkhRht/oZ/696zrbWpP0tP+szLO9
6SAsn0eHSTW3KIQHYwF8TumQ9pXC6+N8j1Oa8Qd+krKLR4O13qbIlWlRa4AyhHr+
H9hHV4x6WP8aTc9OJg0+WdPKMRupzKOAu2sDq1Zmcb7Iq8+s//4LmZtlyihSzVtj
+/ZAcLXXSk+pvKQ4ceml6vDOgzrxjabQcLS4FVWHaIFJ97qjPIKqcxm0Tn4/3apr
vtIXiiHUx+KOVkIW45hmI/5UsFaIVXnCQyOaG9etcg0KrWTZ0QYUUThmiAQQ4mfe
PdpKeEaxzTGlPXWarYrmQ3uXKe4/MkFSvjxtRDcvGpzb1KRs4rxCEJ0lLmQg+ogB
3utEWf8lDxSoPlm1PQoGkOllaAnrYN+xC/+Mt9tW8lfEkjYEAe+bmI/lH5VYg3kR
XAMb9Jmxm4Ap/qIY3NsUaQeAonJI/KDD69+FxCGZFndVPiYTeWqj47XU+ilAmW47
Mhtc55fI+dhwSSpOcfNHXc/alaow4R1AchRSzlyBPmJQcHrQUptdYT3kUoa4jazw
fnIqfzVcV7SIwjK7auNbYYc5hxrTCW2QwREXSSNVWMiw9qIkr1H7LeNl5mYvSKka
SMUf8WWUFhq4fZox8fqsUIB+hMBNA/kex2QJb0i/+K0HkdE4wLOEQVgsOb8/sLB3
vEv77b0hO91dBTIMet8Xe3AumGeCqWdiXJhejRZ2+KnAtKzH13l/hWC+oHYwAJHT
p/ieJfXodJVqLUlr+lhCnrWsxhZHSXGqv6+1Hr4UhHoMNvxARRHVDmsaduVOLTtV
7A+57TXxX5Vcn2MpWjX5l4xHOJxuB/42OlWHzV5cISmhUj3+b1cWJliYni2TDgLc
xeZ+YA8PpdJaCNjZjL+u+vMQrxo2hLJsXMGY0P16PC/ItLZcW83wtOezz47pZ+pl
AvqUT0J3PY0uQGgBEx62t0rjjzR6CwELULXIStNw/FElU/4J2jGwC1m++ofb6ee6
1dDqx2eyPSM0fqgguMs7QLQMut2ZRhbmOo1aEEYCkodgrPcmjW9GRj9KEHlE6C5b
P4ouLvo0SfA/JRgeaalx3Fn5/mQQKgl3h8m9dvFYZ4VOua490bK7OgUdCGYpsGki
39SU1ErUzUDyaNis9dUqfN2G7pp0ZcNBKcacEmzBGiTMQ7lTYO2zTfVopZvpZGgF
R8ZSkVPv02D3hKKjB5ZQWJJJRFXdQvClLqujw6D7Y9brF++KjKnjZtwKR3lbqhJu
uN8Z5AMwpOk+s/hYgbmNoxHnBjFfX1AoRQUHSJRC8YZWgl/1EO/NrG2z818ylK5E
Y6au/e5315VBgtN/hfl0h4l9JbWOTuo7rnGiqBp8WVvDfjMilEVaAjp+t2MmEPxt
12tLaD1lwQ0wLsTgo7FGcR6YudUIMo2vJe7BeTfv6gY=
`protect END_PROTECTED
