`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CXvrfIvF+J4Nf1PytOIYg2UsRcLpR86eLuKd33Va6KxYf2/rwIwP/TwHCvgjndIx
smeKqy74IAQyWE08OkRJIUrruUAXEnfF+cSkz/no1IkgVpzd6vT2lJFEaSjdIr2H
J1GAfYfCWza1TG30gG9H+QJhNU0TEvTPudMl8KhlaOjJuWtPcb6TrqhWYvHtfoPQ
FFIYWTcALhvW1tHYJ0V/OT08TrVxgroFWrYHgKl0oHeCtO1+QfSPVnnPWDjI3iF+
3LiEf0wvQ7V4yM90E0uagPRsuFIX7Sc+/6B+e1JvWkt4/FX5dVXJod3JaYPUjzNg
FjnFhsuDF4hUCQWHLsQGXnJFc/2RRqHHlmBQpLwCTxEl8612224pPgjggLK9cXJ7
uHe1LVbdwirsUyWzBIC1x4JVK1Y0/a0h0hA+s76rcfwo6e/bGZLzvSAkeWV6Ut0u
tt7lpEYTo4JxOuEyoEKE5otNE01ZkBoeWO/rUxZV51Qx/9uhWKN58PMcNznuYf0d
bNdQ5lgRSDXzhorQ7F2z0rRe+gU8ESxphfWgR9ADsHTj+WIS0gR6S2SdNa3kXFkx
OuRZHhtuBL5W2DrCxtQd0ov1So10Q2bO/plCbv5qoQAf/WtSWSuxE4T28ivttzTq
yALxR8migLWQiSDf7A+eRLGM5xzgiqwj0mDzRQY2uUvCA2fJxPO12WKl4OWjYaXW
YP4KyF+af+7e/jD2pUB3TR3DEZUckSeQ3fcUgWrFvxU=
`protect END_PROTECTED
