`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4dq4zm4n4kj6I/xKqkZe9cqMyyJPn6HMKl/dya46AMyvyr7818BR7K4nxpMzWlC2
rvURGkLxC6niDUquikATCzpz3he9oHvNRn74hhx2QknlaYMlNMJ52V8sjgU+a4jp
vSPlww4zzZ/N1lR0AIrYiLTjyS+xKfPuVG4tY4RLO0kj5kjqWsCP33+FVtJq7r0n
0C899NV5JNNCM66OHSAOPi1qXb6fr3l/AWOmMq8YOy1s7Ps/on2T8DTCtunCMqaJ
/UQ0fKTVXd4in+JzlYj82ket+fMivBRglKy6wAjAwhrAwPSKI26sRnE5ZIj+m05h
CoHFbAEgbjdDQhC8gKlIJeFUFjxMr67DSCQQ78vLGZV321EQt0mYB+dkU9y3xuSI
Jwkn6Mp82uAk1Q9mHShkgGrO6gmDVFCFf/SgnfqYWDlvewjO8mAMyRB7rR25vSUs
vlpZdDVo/3cl45mpvWsIf0qAUzonnHQ+thzjejbnFI2RNyYsZbUiDIYiRGF1Y7TO
f6t213N9eP9L/WNYGZmB3ACyxbgle0yjJx+T19pNzWHUSBEQCuTQjECI+/JNueMO
MryWfTWQ3UgkeLAKKSv7NvGxQNDdy7Wk7NKW2hhNpD8sp71OO7cIAw8AVePJc3To
5mbp40ceODCh0kEm6AI4LJMLzA3Zn8zbOhfdsA9qedQ3oLIHapLZpLryFTHcYTHd
7iZRytb5O2lCQBrZoZszK+f49liQrA1o0VHXuZv1d1l/d3+97wTtaqsV4K7ByIqI
dqELtRVOM8iFxLNwosoL/KnqtF67CX4rphELHCiqpz5oFFfujIOq7D23U9HM10V6
KDJD7HvaMO+/qT+KJegzD4i0JJugFJ2CLFkWJ0C5kFcIX+JZ0ALMv30tyKTjHWiS
CZjkNw0+M4AVVDa7DNKwoteBw2qzb2z9cHlm804F0f0rWQLOeQDaa3X6kmHp9XFx
j3XCjOAzSUWNZOPgDLmFk/FdGr7W0u2JAX6ZOhcp4TEqSXt+sZZ9B0bQiurx2cQ7
6aXM4NlhT0VDByWVSRk3Ifn2iUbmZCeQlvicvZtB0oMdC5OOzOm0I/n7v5lWa8xp
XjIG/3snWRSvUUF7P3F7+c9gEQaBAqgr0Ju6MdFIfw+ooGZCp05UzhtHXz2BmNIS
s9fK8sffWd3/D5vWzOpzHGzlZz83VDYuzJ6eiVL5LkVrViH2rzRT0JD4cFCTSUft
esojlYoehrsq1HsDWrqwE2J/uSuXPyunxt/OAGUVGQ5im4OP3tLMiewztsOQCiQA
MVGpotT616Uve+X/aLHjDbGm0ArSLFMF/j9B226aA32RINyX8cZtVAR6z49lF1Ps
By7GIm+8SCm8z+6YBQF30efGZVEFpJob4V7ggVhv+U1qndsb0XDwSxZ89OCTwL1f
aGWTXULKBTroIDafv7u2uEMjrhlsbA91BaIwDREtnrqVDGaRPHysmSZP6/vRjxdH
paORT2tiSMh+EhbKFg/x2Q0wR4HNwp2gW0qHw42LsA8QkHmBKbMxWnAtD7KSQnsu
ptXhpMrNGjFPs7idnRBMVid0IpCXPEHsElsVIrPrY6LUfycXFwW6Ta/b2wzCRxed
pd8ZltequMHZZvHI3FEVWGWvpw5uREH552hkaHUJCwf2YGdbMsgtd1N//8XYptJh
oKzNJSt4Gd0UByU9EHrJWnW19CQOSM6pjCuLce900Hw8D5q6XexId0IdjjT+gKEJ
Dy0NIrUY1poo42ll1EC6rECYLQhWJpszYKvUHeLHcCrRIte9WX0XyWX8zbaHAAbd
b3uiude8/1G2mxyjRmtFR7I8RBQAZ0Un//ALxSR8kcN2xZYqI6gC6MV6pCV7g/rR
BjCPjXSOOiE2qJq65mlT6lXma4vZoUKxBXc1147926tSJzcLgVzONbIh465if2vG
E4DK4oWBk5xCNJTxXUrbANnV4JsODlOeZtpRf4QnD3szrBsNNpGF+ecXNlzQezZL
iU+1QSUaeR/W2nH6FvmQ1pWJ+QqtxxfTKSDdut4v0eBbQ0Hn5ldot6CnXLaobOyY
QjljMPpKrgtYnUZVQYVfzaM5bguYL9y6qELaTkBqj9sR+pt3iS4FBWhyJ4FFdsmp
tkL0X+oca5ER2DRqPXZT39ySoMF0HgkD+ZzCEMVMFk7e4gktijhosX+Q35YWHQ1a
i5sG3dbUGAUwUY/e6amrmnAN6LIJsaoMwgOA8Arj2iAcOYDEiyS+zh0Kk+Pt7zRz
Hh7nAHtYQR7eq0olILUYzcGfm/ago4J747LbtueO3WcfxkQyV7faAmcVdkN852HB
VJ57OmqSrLy5qvuPnzxV6PhknqOvSsmTFbmUNTjtwJHhkxxbchdron3ntPJmsfao
XnETD7SmSaJg7jZzXQC1GtJKVaV8wq/DXaTJ2nLLkWU2d1IQjQJ69wwtMcGdjnsB
Wdh98ZT11L9royMExsG3clfBfixMJeERbR4K+r9DAwXVaWz274UuoWXGN/nuErKu
CHmvbJw4xyWgAOJV/S0VqLw71I4kCHY8fdJA9FgJONwp6eyKQDLPdtIj3UzQy6vH
isgVWeenXewW/DmzpS/S+UKmwTapuDAJ7PWEb4QF1TOrltMV+sEZ6CnNhpt1oDWG
NXS963HwTcv0hYbkJr3xJ2B28rO3i2bTaQ64nR/4fTII0NhzIJJ9dFLawx/zL8HD
eXJD//D4iJZsKWrczZdfpm1Avx9/GmVbAmCQ5IE0h+UB8fN0oReyafI1bacu9ZwG
LzvxA9LYbBKE27VuTfYR083vMggysnAy00NOUBnKPurk3SPzfndWcwXNHEp2Sh5e
ZFG8v76rWLA9mOw1QmEg0EQvZ88UTz9wOjvJCmaoXaQxBdVAiwzVyqgrBoqlOJWO
Z5eWJp0WAU3x8lnQzV0LFA==
`protect END_PROTECTED
