`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sIz8/zxuOAqAF/bldf88YK69Ew22jVVv7khhAO+NZQ02BPPzWqMtYD74InCFfcZ8
kuSwWpZR/9uxJeIf29qSvr0ZSqsG2rYeVYa4a5HvICzJ1fUibm9TDQ66f8NCf5N3
g1eVBpQyJ/BCdlvtZkcm7LfeQtfDBFfufeTARzQoXTcrrhl61MyRkP27e+tl5pZH
J1lbgXMsnybEiTdIvQ1FMF7+gDaWENgWHcx0LUC/LcBJRGnabE4sWEgH7tfYcKIj
kzOVNXnV2tcy1pN73hX/ZRe76xLH0Sm4uAehdYxF4PFtBItPIfcA8+4t5i/Nnp48
bkynn+KoFDqpNGu+xO9WyoLFRkG/ONKpcqUDHXCJAnWwdDqQ9QNeIyHbwtiHLGtE
0ViUQq7RYiX9DijmaxwHHovXZJQ5vI1R47tuJcTzOvNQWWvZGY3IW0BdFbgbpbcH
N7klFxzyqUP2zoJcvniLPwLn0c+4BTH+NfZXq7sZX8b2vuGuDdxGUoXN7tDP16wV
h/ICqB2WV9UAmL3G++jpRx3AkbCXlf7zvO5AYHby2tTT2YdiMTEFDBVIOBu4rBSx
x8iCwFJgX6Ujy4ChyVpnm/S6pn7znvosZ2c8V4YyAPBUpeihJVeoMN9mtlv4Wqaj
QhQYCgx6N1Yxwi4TSUhJsqj8IyvlvIlwYqB8r7fHDC37QCHYSg2Vqa604svY3KxS
9+x5cDM2Atllcnrx7G9nMZaPUpl3FxrYf3xFvJLr9efV3ZSLohf3dEy30znt+J6n
NyuTTBwo/paVZBlcf3Rh1erUxjbluLRTXrm0Vm5WownIITXRmuJQH4SF/Hndj8m2
tQxiqH9CNRIeeZoHSknKgS33wLaDMcI5n5BssWMt01XtTryxBuiaVowU5Cx7CaMN
Z/2itiVdBd5LB3hFyNHxxtcdIX/dRJxGIlRTbc0x3gACzakNcDeum1Da3yEk1Icn
a4lEA5NwHrklE+daNXy2+bnaG3XunrWC46J256w7OQAk5dCdHb7S5cP9KPFPNMTf
Tdsklt/S9LijGR0f02si7hDskMKRIcR+D78v59XrNdljVFGnS/1J/g8sUu8pqY+O
ChgIPVqakKI5kzZnhlkpWxbkhiZU+3PEomcDumDikiiEKPVrXT85ivE4MPSWpCVb
h3/Q4HdE3hQugtFN2LUxsW86yLw1ztnngOguNj4e0I2mOWOTnq9no85H5ILwYNLo
lBb1ZAS7TJfdb2r2kcGdVWVL/0gGdFn9a6D/4fTLD7pNuhBF2ed9eofiVEROZW2E
SaoUqHXzY+vB8US+ACBw1uf6+14PENQ/vsFlPMW6TRRj+O57JvI77DtLCT3uSJW/
tXQXTH4igXQQ/0oczMuq5uNM52rhzcKpz6C+0V1GfgnZUjrhr8iHWtspyNGd5zTs
qyveTB5137Ew7zF+fA6nxjOagMw+jSS5XjxIJzwhjsPc6PRxWKIPAztKprQ7LbzO
gkle7sCnpq6luhUB9ZZl9VnATeUYmq99JZcccCk8DGcx3RN95YS550ahziT+OPk+
8xNE5f21fL9Rrc6x09qu3MCB8giaOE+r9NjVr+RB8gHBlG0UIXgfVzxyZ0ASMA6C
O9ycsmMfENIMJ8GG90IU/PwM4SXwFJcQrzwHxY2UXJFApmA/ZxzmOm/Crorb2Hac
BvvSMIs6PimgrsQSamZvy0Wv63GaOtBiFpis2HyqpJ9w0Sf5N+qYgMtvxWXSyiBV
vM5egItQwS7RP+iPHumbyshJI4wdcdvonRTHRSbsSLICZ1E/QMcR09qNVhmiygvA
oCddcNK+Dwf6gQkkHZ7mwaiBeEn3P/Krl1msWrkgPQDrPJPaoESX54K0+QF8RRc/
VMIV6TUe2imt6cjUoZ5kul4MBae+QIFtYaKf/scx0ADST3/mdBhthBpKbgs0Akty
Pnke5HDpyPCpaKpTlujX4BOopV+MlypjPEx5IOdgjz40Pt5J7gs4+TU4+YgLjRDH
E082+m5LFEYnkBUmTyLP0adkz+aFqi9wKsc30Yy6ev+U/T3zw98tkl1oYyy/RqwV
fZn61dRgQGDkb/1EuaaUlBwpRS31lOo3Ohfvvtf1F9vOrwDi0h3JE+K37RRNDKKQ
E9Z8Hc+yQAmVn1E/KiXI56gjRF73o4mJXN3o0k4sq26SEB3m8yIP6VrChdkIO0AD
jPqVJ6fkK0ibP7NMLxWxAAj7lGM6jspBl6nDf4s2kNJD8UnQXVW86UJZhkXypDm7
I6Bl2MnwRN5SjlnGjqevNqulCVRFLQMsK/Ow2+dDPrNlFpbi+p9WOzB3wCvDHtjG
A1VEYHG/XAJ7WIIlVbgHMgeEsjhThL/Pxlbetwd+h4e7dbIhtOgSfv57ui5OddTc
RQo0ij982U97V8heH8A1x0DvMwthoi/FfCLMHfQvwYbMGM3yD5L/wJSumRkVvD2W
Ym2HDMzOO9Azn2G1x790STtlM5QcXpGXjpBaCNvNbs7mTGjnZoUw2idkhAIlokAP
Mlxo/DpNhnDcUECscZ8JbAYTSeuG99wwLZAPxaTsdT469zr8xbxcxIsYRTDM97VN
UGLvL1cO0MuWmWkJyegdaNhJDEk+9Mlkd3tMXkvezu7iGOV0727vTLAUgv6IRZbN
najrLh2wNRBh2wShCQqwBDSViiu6psST/QafR9GNsUnb8yhusiUYgvB8zI+fujt1
ttZSg7zBcivsgDQOpRrOOmSRK0hTrDVPXPO/1ORJCM2FPL85VVGYL/ZXdRo16cTe
kI812GWyidGlH2tCbWxJuAXAjS8GdD0m5in9A33wqwsFUi0CMa9FkgbTLKTGGFjf
PMCRgztSK1aBB8m/n3HqgShoNI2BDFvyoeS9ERTriOVJJfvPyrTU1GbV+fSKCn1/
bczTGE3uF4lgrLrTT6ACy678sA2PzrDyXLkddJLoQMUt/30WvW72VUajXaFEhQwt
nA2dRg4sqbMPdTrZURdT941ubJuRLn6ai2cNOMJo8JSp/mH/TiCZn3OXyIGwO40e
PvJFw71ikf4O6Rc390s4ntnn1YPMJ50dxse3NO0X+eYY8i2XoA8YbAjyKYNH9LQK
Jm4QEVuZdJkoYnyHYQEu8bardZ8UNv85HykLLI9Fc1ceKvO5iB7TqTnF5FhllMDv
eisOqIakP/YXVyc0gxbuQUvLrW3xUmfV72doEvtxDoV26VAhpztX04IVKyTE2v9z
Ve+2NdwNA27M6BpzbVXMhp8CtB9Qb1QluaOm7NjmSifNVWlCOFX59GGJ12/Lc5gD
4ThteCFj7mUPsBAoo4WRcl8V1X8QFfehnhbqKSuVVHk=
`protect END_PROTECTED
