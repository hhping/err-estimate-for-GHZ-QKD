`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N+HayxoHpXC2p7dq2J/tZOmA7EeetGesMeFzgxD/4VXuLL7+e4KofVYfNA0x2qTB
Sw7vU2gUVO1lNlIdVmCBnv3XWzUgA4xiJr1hz3f50LdD5MmBpuKAGSFUX59nzgN7
onrb0xz0oxpcDOhdYlvObUSLTMdrJZEJnmHepHn8xJkjR9SlTpA8qXL8Vo5fJtNH
ghdZNv/IvIDhxwvL8bTNonta+x1sDhb5erUhqxEVIRvdKJMwbdITVfn0quJwLF7j
kdozqMGCD2q9qb8kI4wvo5ilSwy4JmezefPq//MB5vFSaOIzTetKLGp5pWVgmMe3
jf95YEoFDQFSMbALZsjpi8R9b05xvgc0VBd2Bfsa45W8KRzf+wq5YTEHObneD/s9
u1VVOYOpIAis3Pfddr1xRrWiaJ3yT+VUcqg82XBOMmCzgV8mCTtAOqWdfM/0OdYW
gH8BqUiXeb3hEpl2HapFDHcpz/PXzlC/QrcmQmOVLhDSDxwtiz3KrT6FKYttPysI
eitAtGvouNKNrfp+h7xQoQ==
`protect END_PROTECTED
