`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F3ZvN7LIQn0QXt6sVklop9nUPWNR2yvUkpW6NiTOfgnexQYgw7FFwXxH94UVkV1k
vffYuxerGCWiJx2vwjXOm29HXPMGEy/xaM4oWWzxnMvw4YWOYBJFhCuaT8saO/TS
DJhPsD1gUNHRYZsPNU6IM6OBNcLDfDMxuSUrvMgEZ+wIp89wJtW3u76ZYwlsYb3i
7FTL5wX17Lx1u/+bdECPt4VGNl46Z4KdIH03we17yqt7RQ31Xpa/VgNGLSFZzZcJ
bwh2gCR1OpnCa2ND6sXGI+zkQY4JtECasI9Esejy+Ffe1UM5ENCzPnfP3gahfcnm
ILJz2DzupjNohZWFE9XqLXssfFRNWLhaqgrPrinquAp64GauzbYrxLyVYVIUHEzz
Dq+M1+0j01SL7+OZyiTN3C0AyXCnDyDwawQkVWzqWNG7DH4smRvufOgeTMnXL6nD
e7nYOF/bKXaFe1pN4eHGDZJhiwD5c3hyKGIuHrLcuSjb3BKHReM/52W1fuCoHcs1
K87vRrUJePWnH4ykskpYc5O6FPxwkSwxEGFKUNBmP8XrndHAIaLL26CfwZMNiADj
ikSDO+yuffDdqQrmX4ygeFERDOdVmRqGRYTxJdjdMGWasrnqQtYlN4rh2sxZATEV
At+QbMTKpBEoKto6QfSXSCkK/6z5WzjLa9Ft0R6iHNvyuhcH0F5EwkCADyP9mIMK
VHczQZj83B1ZmqED6C23eOKZ2pXI1pgbLm2yPj0/Eq92vItytH5zWAYSO8EqX2OM
9x04LuxSzF7RJJcYURCUQd+YTotCOx3s60Piv99NFPLF+XHSDop6eX9GbgmBv5dj
qKoiiZDqVSYHmJS6yZV82SzvAHoVD2Ims/PCEjndfTsUvfiMiV/mNm3QevnpZ9gQ
6gsf0zL9kYlq0ZWiM4RksABoSALXPZ+ZjCjMvqJ7GtBswIvYzkjjZhyg7OARLzWa
MNP1b7B3FvxuK62VpTpfQ5DfVpdpYZ1iy11FcaBVAB6VleZRuJXd6n2yinqQrx2Q
hH0FusvLW2x5Ays9vNXhJ5mq/RRT9G3DD+Z+jKfPD1iFOSNo+0iY+ulJ0Bj6vpmf
oRXFQVRuEryMb8u5Khm4B280gbTxaIY65SsPZBQJDlyKubghaLZ6NE63wEzQK90w
SA68fIvVr4rX2Ko1Ot7LoEC/3qPicxA4F5HyjpeK31LvPHlLIQTpTyuNnp3SYucj
s20ixt6t2Dml8MSTn0oHuuapYlQ6IGFujyyEUPDCR063bkIlRET7SQUBzO20jy6L
8IiaFN6bPvWtH3tTVFgQ6TUuptiAAABUBW51Cx7Rbjcqu/EA10EgPIENkYuDug4i
Cy34NAuZtWCVglkGzeduakrvPRxpx8KNsf/UXHB2kQl3tUyXDuTi5wqWMPesDbS1
wOQDRNxpsYAHHz6gx9qu8uYJQoBKS6r1wf3/iFzUub7HGIzYNFOqIbsQkuJZsg8v
Cs95Sp08dTbFxaKb8TW7kctqA8p2FxwHynwvL9uPJ1Ovb9DPGTKgMjjOQQYhf3qH
GTa4pgqNusBY8luC3j6imqSfoxVmt0XWH8yTws0yo2OYpjujep+Pe53lkX+IzBCF
dHBPw6+bxNrgZ2qnqdAqSp5+fUeFJ4F54Y46GTqfzqsz9rOJMJHZ7QClywxeCwYR
SskkA45kiBvtLTo0GVOwHHmh/prQ8htsHrY5na/GW9beocWPQffzxma7wZjtSw0B
g/yGq8VdZrxFlwQNdgtb/mwlTksVoKFdW1TNf6sy3U1u1xINdX7m4+9yvfKrduf4
`protect END_PROTECTED
