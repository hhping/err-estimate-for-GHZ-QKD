`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n6eEIYreOMO0iUpZ3rI3tpPb3Pgz49C+gG0WiLc3OaqRIiDYrv3PRUHbtJTwjkri
sEcmiugjP/XtVb5EARtuNjY+FOvkbMagmgSs2qP3Il1/i47S3aPHtC+D/euu89S0
1hxUetgocc3S/FZwYTwsGEaoP3OWxHuY6DDjx+hIErGqDIBG0UF7GDF4fDBgNCPF
rT/W5ZjAwgy6BIt3l/2khuZ0+HhRKd8Z1VP08RzM8JcxRe8dL9BcS7/gqNg0rWui
zCGxZBlPss6XODDvgB5kAIuazTTx3SVeZ4YIXcOTYpa5Te9es2Fk6pQhQvj+5HrQ
eOkiwz7v6l6S4b3yJVgU+nfbHvVDW1QcvJlziYV0VWks8rsugFAKxjlSvG2QGptJ
HOCZW2raWhisoLXD/aiVc+5lw1lqMrZr4pHJ8hRUHTn2phqh4f3CTzIpq68YyVPr
vNvjEib7HKOZN3+GxdD5rg==
`protect END_PROTECTED
