`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cNe6lnJgEUCI9xItGmmMROnCiIxL9gG/Q31x5CqR7DgWu5XpMW81i9MXh3mY+XS/
rmPc8ANB1CjuWjr9nhfgv04oetgh7s4numZA5rBEma3e3x4E+q9b3IIYMcB7U3iX
CbKzh/kz1P8L0Q7nDiwFSQeHImNiRhNGrW1zQnCW4JRXR2yRzbonZRRON4fDYSgd
Tcs59e4nkB3laLZw8ZUesRSt54FpvPEpR1Am2HlQEELR+ToLUCE3QZu+x5spRQ/o
VP6+Ks8YNWiCpeYETyoYhyNe7JSJ6R6AL6H8XxumMxN74xgOdrU5rGTTCG07javq
VgvHx+tgkxb3IjpAPCEzOGCtPZ4rmGvhwzJqE7uCN4uoiU4FfYfpDijGjcyktiUx
yDcnKh+YhfQyQbZoXKyEFEpgnnm5NrVP+/IP5dRiKcHZ32xiQl++Dk4OT7ujNEUC
vPXpflVzLNLa03hJhBNGU5XcbBu3CHoOTHPh4XDR+ZrPIADvVFfEvrmpwm3oIxHX
NM/v0JJU4GEvyMdKrlBTY6P+Ctq1exNkcogo7vh7/0Q=
`protect END_PROTECTED
