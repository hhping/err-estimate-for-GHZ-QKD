`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yrtWFFKZK3fTjI3/U5QJDgLaoA9MLK8RWZameM9BxQrWwWtg+RRVNRIlQpU++uRO
oZX2c7AzphX/jA+WUDws8KxpN8RylAUt8xXVpBuZfqM/0TKhpkbMcvE81oqbqMPm
5Xk6ayh9l/2KunNWJzDgAx0mRcD+JYb0hMWDhoiHGrkXNGjQI/m47HmfdG9c6HBU
u2+YKF/A0flkYiNjUfi6i0PrNCTNJEjf2mBfFXgZC5HpwYp5dnZYjqXAQvGtEl8n
KN7nwGeIIPzWW0FjQHvhEwTB52OqsrVW2WjmlGHJNnB6iuuNkHkUnULyzeCeFVvL
GZYrd3/cB0sXWVvosW9Yj6NCjjLWJ+ZKS/wc31ueZAITQL4UpvyhorHTiG98JR20
kJEnjgF/YL8RadPPIYAb6H+PQzigY2TxPKVZ/b75J9BkBi4NNpV36tVpiuM92qGI
f38Zdbr2pxWWZ0jpY8io8RsOtqeaH/wQGP/bYnSyLAruVFDtag1LC7iktXg3T4dG
i32AA9CvDmlUg+zZcu+FIeWmHdjmlCdFQJ8/zodzKNyt4FfAXrfBWWgHKKZd1ppP
N4+yGhe0fbXhQzySTKE2gZx4RNYgv+4SPOdB6o1n5Z/sAJ0jir1WV9SuYQ2KtsQt
J9lR8d9oNOU8op85JTWN1SBFYjWAZlw4Oog+wdQN9crZRUKiuoUEnC09sDy9FZGS
jSNl2pG2o4h8qHr81o8JBmj8NUJ9UxcKVhWAf0LUbxZnr3qdEZEalheA0JJcyvAw
d8/OhAFtVRLI0DfP9d1im8Kk9fhnvSXjxwdS6C+Ve4U0SiDq7hLQNyQceACvMbyn
0uPqEff0l69GBXoITeZ4g0QnH/ORT2Cgru1fnbgRfwUk4gfrFirVDkftVMiqRgQz
jY61QuSCS+3BeXk/BpiaxX26vcCyOGt0K1L+T4DaahzzxR7evHqHeawMbkLURrKM
k6ieNn8OxsO/mOHR+efUWLaW5YDs9tg1yYOjEfYULtQK0AnELeuqOkoz1/EVlB1T
B4n49gkWmG3BKZakQNHHqA==
`protect END_PROTECTED
