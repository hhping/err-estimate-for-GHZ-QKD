`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a0ziIfDznjgDtrFccEOR9XjMw5McvPwoiB7x/oMm6+Z5P/yVWKS3AM4XphMbe0Bg
7A9mO/g2LemF/IXUtPg4qTUwbTDeJKyZIWWiDXxt8ykX5NyCf0E76gTXlp3m+9r3
BAzk+nmmGQipSufe54EYD0RVp73jOmEOP6dF9phlOF44k2gNc0zVksat/ywJj4Bd
wG3KMLc5MhPdspB1XU/6dEe9HHAdXrUuit0QNs8Yy4cLzT1THFUaneRPX4gnj9EF
LTcopq66wGUB4i4FZaRDYKsxMPcZZffNLIqWrobQBXJywdhwh44+5ZP+vLun/VWf
CukJFMwn/Xfbw/pzwB/fuCuNRU5kb8ClpuS9Coypq03WL2lg0xor6jG1KobvXHm1
Hit5dZeG0UbtTps3AfelOFRHWjVyYWiSRubIYQFXeRsXjRXfEmXh7wR3barzV6uW
WwtvLoWRk7UWQDBY5P/uIWcY1+VwlacJUoRGpnGrjKCkoll6uhEl7lGA1jWQ/4Ch
BGHRzebGeGb4yxvhrJs1TFfYyYERM04GF8j8rBkrJSqdCODctMdFtIM+ZAiuDN0V
aeg9NXixYyHEcj4pCLjIQOlKV7q+e0NwZkN3aWvvBHogWmPDHcy9SPfkZVl39oIZ
NpgUetKRbcta/Fm6ZwfahEdr5EPbDpCv9SykIy4HYnlsE6hPFlVSI5x5qlCvuNrX
p/JAOTXlxECS+bzWkmBdRvTE98fCWg3287/L9pYHVsFpOKPJv+KZVUCBfX74RfXi
Avev03SZx0/zOqPNh6PHyhQScA4Wn7++x9xFsjP7SFi0+7ppiLot2J8KuLiNhp/t
UiuwAQwk/jbOm3wLk1uK5mXTgIM7krwut5cTchTaSJe0lFPJvg8iYIudSv5gacK8
hC+3GKA18+jWAMcEMcsZPl5sZpqg9cLu5lSJ0MGdrvFgJzg+qg0t1WDJLvHZmrdA
J+TAe8DM0xsPUzUHKTUl6Q==
`protect END_PROTECTED
