`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D8zOdHWxqjyuCatTfv6rQD8wSSempcBcSZU0AH+9ilSDkil+5epiP8wJwbdeZF/c
W7SircctKfwiiJs9IaAF9J0EXfJkaLP28Btl7P+sD9eqEAcFOt4r4gjqAxuCEO/Q
m3mTOYxIqo0UaJ7F+E5KA11eo+ORCzMX3FUPxeuu00rPjHuZt1tFgyfU3kW4aTLc
o8uVJWaB7UwKlVrC07AsVKO/ocpRvPxnhAvbSvQtK+9lq8AQgpEnmmLSvGZQrXxt
YQG6YLY8G86/Yg+ZdW8SKAq2orOnF5DXoJj/qTdIskMewS8ZPwldyf+yKn1b2I3E
YOxx141WO0a7yt5WaogRGrzqmn7KnS+pulQvhdF0LkTSNr+AhKPH/s8IYdUXiNuw
y0x7n1+VBtHVSa0NdT+ZTwjGFxM+XEHhn8CdkhWnJiSAM1FcDnebdjqwjNY1mel6
8oDEKUmwtdrSrncXV+fbNrAy/zUnPRUgoMJYltLekrnynwoqaRsRWxk5U7eoLXiJ
PUWXB1cFBB//ruHQEgMGlw==
`protect END_PROTECTED
