`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Igt9RcCHF/nENkZ1EKFXW61ntPXVh5rDIVcyQaqRpcAL61B32aPTOHLyVid4aMpG
9kqiWX2BjesclolU2lp5GV/o/15EbOYqRx3/VAFP1SieaEqwcL4pcbg4t0FInF5H
/PN1C7CqSvtc+K8N4UuhzKSuYBnIuG57NNP/e6aAuzslgIgdQJ5/3cRJ99pPOyvw
h0lpPWMavNV9SzYYpMl1Xn/cfEd14o8Pll+VTln5EmLgeGXV1ZRzJVMPMOwrRWVz
n6VxphqEg84CPgweHQgKtfTWbNm0N2shT4M3AvPciuX7z1FpogX15L1r+aJ9K3QL
01IhbquEL3H7A0l8BthXFxillyEj5ff5AW8eUM2Wz75yr5YF4ZMveeZAubtZ3LV+
TiWHtGE6f1G7lo3FwEjf8Nojw4LW1qfv2bB7b6LG8edpx0NyPuOI1d4XurNdryPL
H5ezwtwEeFadm2UAnCIWbp3kvoOE7i9U6JgrQ0oqBj5+oOgCdLifLubKfrdokvvn
uqXPYAXoFgrgrwYl4R7J5lzH0X9Dvv4PwXeKUlTdhSRyBEsh9vBG2+CbICj0e4gB
J8gKxJNLbAgQOx3Y9z06ZCW3/YS1iuvVo9eT7qcsoa/T36zu8yZIjStZGZElUYtD
azrSIsZCP7KxEi04TtrBl0dKvUOsC7l4wm+S79taXU6PGZRcOk4Bxx8w4D/kzZlk
Y4pVAiAMDT7bJnkPhiSmYtsXI5oBW/15IINCQ5EkcIBqDvHsFhIFrAJ024mo62d1
y1pN87+6Btx9lFULUOl5l17tGGUK2nHLmj4x+klWk/F5RmcVAuzwdJ57keN0aVUx
1nA0VPZGvgZghdaADUNVeeRA+CBvrMWaFuVYA7IwmssZW5pSYdrkQwXPJD4uF2Zi
YaD8LCDdO14Y/+OqgbE0uldgJLh4Q7VYS1vMV+ESUzWAtexdfwqtyJPR+SrSwyM6
Bm8hVCdFrX+eDpwFZn4Ck1pucChAwiGO9LpVHz8Nwl2asxNZU4rYXoWyYa3UWSxn
tKRzIazDT8/A8hP5jLh805gdnpgpi70uJpAX7iR5rPTZtT/Y9ACHewozmAdSOzc2
29JbofiYrO1ThSoxd1zYD45fNnpuavemMkpzSMC2F3tHd4Uium5uhTUaP894WGN0
DoeqQ+v1OvX87QIB9Zogk+aHNcoVBhKIoLy36AYhvP58Em0PX+7QRU9j0km29bxF
jJiImRqssk8C12Hu3m8v3gKmi/cM7rTtEnuDqLSeo/YgxpO89yAkK4NcxBklwegE
RwDhMwgU9095f6r3AznwKkAdynSjqF6ZNFULv5V74/larYgC91OHuyi3ZDWMvtjo
bB+WrhlbGHT3aCxZwzCYfH/XzmLRUujlMYtidm17gEUkqU6yboJBY6R87rj7IxOT
v/bMGThN380U59BBQDvT5QEfPN4m3KcBY4QTa2Cbsd8cTjg1T+CoAIPPV1tFLiKt
kpOLK7+NhocBUMdGv1CqNTfM0LUUeI01TcOR2xtM6d7ww9acWml5Yqw2p+vTGe5E
nFmNZpmvtuRTfqTnjvOaHTxexCKXmZDT0D0L26ld0ZyHNvwwHkv34xB/Crmna0L0
0sso+nPimxTrQnsDo+ZMqCzRQgC3M7sJqxsf2yI26VKP/P0mAQnOHRQZ+2X4HDf4
AgxPm6wg+aN18a/UAWE7drojNs2guN1j8mCSRRrd+Lti4YOkHanBh5kn/xNWavkl
8e8C5lEdmLlK+hsFv94bUL+nepMGisPqPZ3S+1CJd8x474Ctz0RUrJNdvEp3vYYU
l5T5pwlccJdNzYtzp2kcoNeQFV11chjDcAKs4xMtc3klnGadC9FhSQPak9wYe78e
DBAa1scRbGAsBtnbOb5I5L77fTmRNw3uRCO354msmTLOS/GPiMxuiVSloOkt86Sh
aCWaePi2SVxHhIicLDLAp+TDqVWeQR1C9EICgp4HOUHQtwdGRoCJkcu1bcxs/RC+
8CCAKmUDYLFgEOwZ2Hz4ms7tBnfWEs2o2eMTqIghqwACddCXiW6iMDcYMno3ioAq
Q4RWRO4GDPE31VVMx4gArD+j7tcpQFcH2VE8JDMXffaHedhT33/zmqXNUiOCqGcw
RbxXy2hH1UufnKg2Fm1+t61gow18rg0QNZF7pvM9DZi4B5DM79IVIObz3+daOU5E
CZJTGwHJyvqCgBIMCu4c3IVguNZcsifXx+TDBIq8pyVCae6jhj5vTggQETWnM98j
OwJOPDwGEY0asIjOo1XEB71PqFrbsKzbIT/2NUgT3kNdkNo2hKDDRsEHEcCKJskN
Mi64wDLOdQmeMDg0nPR9dzFG4dGrooMdLcwDuWov7LlzPX+wxzoggoeMB97Jp6ps
LtM6WGYS0qdLshjAT1lAA4MPHqCd5y+MP49X2OEYaQQ1KTCgf29rUwx4nFVarsrB
lwrzIQzfxYjgmsJ55R8pB/2W645wFxIFcQd/ICV0tLgXRQfU+ZoVSRQx9wV/iJVq
L7EbH9LCWW/+pXhj8ROVBYW486anQcCXTXcAqM/fonn+BrgjOOCwxaN7fSMT/oHl
k8j9Bp13TAGlfOHQ5FkJpuKPbYJg/u38TSJcOfYeehtHWYJ8KT7LCb58hN1ByWDO
/4fnlf5zmHjvqGMR9wBqHSy1vRsNYqcqd/RTkXiceeG7ySGetiSJPpi2Jj2FHNx2
SlNEmYClzgAlCHZXOe2Owi1qKctfS6Rjn8RLf74oNrbwa1Aq++cQrHhg3Hw5+J3+
vSRW6P0mpirxgky8GiLFbHAIo2a1nxK5bBTI5OBHuktyExkjdK4BBUPTEVmoBjxc
sU38wbPm/dqu38IzzLKgxdTqtOVJYYlczzZIty1O/3qWjn0lu6FMzQOmmo8e5HGM
1JH0ZEmkENz+YS9YJkn+NbSU3Vd6mRd4t1Y2//TosJZO9LovgglI6Lb17jLtd45O
afzkr7RJu1PXh19O0b33PZXahM+TVthe8JqQz+anIX+rmEbbZ3e2e4NBmKeFuNnc
yCWHc3/jZVFNBXCqIAjew9q+NyqIdOnEONIse14YVTXNXQbjF9uoqJRowEQwK6IN
OLWlvrbqslqIwfcqCxjxrYarxOjxNb/iAu+WmHEvAISL2A8Bt6t+y1b7TYlZ0wfm
tEwYpjF000M4WPSB7vcrXKJ3QMvVkzbmlyryFBIzNzH/HzGEXpG+w6c0MhF5A6BL
WnNAV7Y/8qtlY445Miw7kV4h4DmVLgkIbTzNyphG8uJEbmKKtqn9puLV3z1BvdlA
dVrIP5xucc7qz4e3PVLfAcOm7B9JYedZY/46qjnPBLk0p965vv49Rq08ueil9Dab
wTWQmp6PEjmcwdjjv6MTgkx81FdvCVHFB9qfxy9OeTWyKHNpmvWGd4Tbim9vfk1c
cSbkv25e7lU7/TSLX1QMPlWeiOtETfuqpL5edt5CY+BKBYTvTpUJx4GfmHbXv7Es
8x/4uP3UY7Z10MfFVbnupB/ushUBOOFt8NoxXqnNGsuDgF7ELt1gPVi85ML1pNSW
WNGUta/2PkuqZ+V+QVACo6Dh+30tmQxJdfY5+PZ13mx67uP7O7uiiNk5dbuzG3Su
KGDmvlrs9oWp0/9WW15iDZCE30yfdcrspTwspvLZ9hsrxMBrULqiUc6HXjaZdDng
BgMF19CZF9rt0/lteZAxfZWCyAuAfw6cDxwekXrvIxC0sKScQ69YObzuzeVKjPdW
5E4NnsRR69fto3+NV+y9t2/suvHplDYJ0buIg5XJ3TbRUfmKMyM/4/sZL8jYaGRD
Ibd/EPKS7OgX6/2zrnAtwCu3XD7+kJMYBjd4jc8/PwbV8MtZOHSKqAtWy36x/UL1
Qnmw88sVq8Bl/EByJVMu0iBE8J/WR2P4lfL8ETxrl0Q+are5nSlfXqAFKVKyW3pm
/MmRsMBfNNMndhx/92bvjVj46SErA9Qt/owcQ6ziAgrSxtmR8OHfimDv5V0Dd8UF
C+LpjyuykJwzFCNFGnqK3zA/Y1uO7IDhOYvwECq7zuy1foPi7Sn0BMtHbUTJcCKA
ZoFFCTaPj2WVS+y1dzeAkx/qOCe/lO+dafNQ7Fyrty0kTbVmkzeDjB4B+MnOkx0Z
HG70thYCOCvFatqJpjgiBb4L5PHJw0hJUE9pWkJzY7MHCIAW4x18+MBHAqdNrZqw
s3oFm1PIFPbKQRtJleY0XKcME7OdG2s0as4Zt3KjuFLLj83P/tzAnlh9EHCrGwfF
RFxkdGS32ryl/eTbIZZhoIPgaSw9sU7EBVQPtCSrp4f3wO0SJtqmrzGPMHrgBUeH
JGrbBzDW+1wGDcRbAzdILjPF4npCO+iKe8Eeud+ciAQ4q9hijB7rYR5qiC/W2BO8
1bO17TtaUc9i6/suM3wbDZUq/NhSP/Oo3ot6j0RX77lOV7Gw0O2vJU5kl4h3hm7n
PP3jmC7Tp6uUNd1U0WnQMKYTHNv2Ts7b5v2NxmZhn/4S0yqWAbvcn7F3INa6NRmz
9OcpRxrflHfHbrrnWTz6AkRVlQn3Skvh5xvGEzGsU9XgcoUScQYwLVFQG+TMVxsY
7hGPwxeNIEVd34tjlrImIYav30DpgavCmT0OVRk8uLM+TRA+tubBJtYq75zxZnOu
xhdacjdsYt5S+VrICJizXAxOwoQltLSnIpQVP/biYeLzYmmJuU4vwnKURXAS/HQy
rQKTFg+nqX3HjETDV7WQP9yaoNmnrlpB/VGTml71X5O3QCbNRsUQl6YhCs3/hikX
/i0s3aGCMGrk8jofgE6DSn5tpcHGKB5Z5A60qyZgMfbbDvEKChzcAxa6diS+wBtH
eievU0p///237yKdFDGG5E3dGtzPW+DY5ELJUNfDCJsmTD9zLEPEDOWKG/zhZJfT
562R8HYFgI3ReKHKXJBtnhxXkVHu7bSQdNV8fhkLSrni/ixHNi7YLRUuAWr9jGp9
HKpqlcFgcJpcZTdOuS2gAAdYZq2Cfg1j6uTjQKFoUIIVlznSSWsxZ9rcjG5qkf6i
BaCiUZTW3ww/exlNZz5RVZT0+12Q2cRBsk6yuG4xGu4p2IqMLBsk/CkQAeyPUSgB
bU1aBYfQnOViqM/vujzhmLwpmss3eNyARchagvZM92DoEmu6jCly5Z4prSiU/Vut
J3WuzqZd3Z0dkAlHFk43/TqPvNcSV0wHmLksR3Nd9rxcA44NIRFZIubmUvYf8ryV
hsmvIl3x0IheXFmW9SJoSanuDx9dvISF8poxWWagnaLzZHRGwjBdBulyLiMZ3b0L
72kCITftGtyyYwVCew2YSIupsRGeEY1ArnkHXA1o+Du0elWERlEczoX/ffHXo8Eg
kckXq/z3AnlOW4i0o13fGmcO8kx9G0r1rtmlx7rahcFwrJV36jif7hRZGk46iUK0
TFhuccwUYWJTQ+VKLXLZFQ1V7dkX/46Y5NycVYBBwEo4IxvOehR/rwON2r1WYhuy
EzP9oNq4509B6fONAuU/BOMt4sUng8Uv7ipjQBzR1uSyXgZ84+5NLK7njhkUvxmp
5CVNEZp3jhAbkiDpUa5eyC+mMgn+1QQcB4wBLebnofeS44Ys72+wFW2gfWb6yE3t
orgTK9MM+sMC+H31eWewr/q8zJomAcNH144Fmg4LY3U53dsWxgn6nmN3al9jARzx
txqJ+zzo7Pn1fIfkSDMsqpAEeV7+436A/6neG3M08B8Q88For+dYhQSox/caahgY
G3I9rpnb3PIEiwlWXNU3gUy1byVUFWvLc0Bq6EkwfAAzpuN6zUmKvu4SiqHjtjsV
kuytdzIyyJdCjz2CqcsVkkcVkqoadJSJOxzNnEMjAayp+77XhecYfPJzNnx4xces
re+A/bF0ulZJ67XbZSKgubEImjvX7QN+2cMYleYcUP/to/XRxfAcHJnM7JMAGKH3
1gFztMntJFnDOL18B/8TI+nIu0NqKvJ/HyKRtc/SLVkMmBh5QVwdueCZZawL5IFQ
zH2bKdvn3ZCb4jtjY+58vTY2LONFL8JEVzbGHab8/hbV0gyZ5hWubMGRPNw5Opcl
XZDwcMjdM3DQHwtZQeSwrXuJRWe0uD4WL40RDfq2v6W+jTjLo/uj2h4ucNbLIEp+
z5jvQX2s/B4LNmi9uxEJuZmZ196fbc0iwNWhPCxq4lOvRQ4J6Ta41XffIU4VX2RV
FHDKnKpz7bkkP07G7dVbmJldvQh8xGJWqZ5p6xyavqGsLhL6U5/hKxjVD/guh7PI
wIJPTJIK//zNFDudGV3EyQ4DMBpICq9GywuNsL/KZ0SNrJzlhvugNCaTmk0Impfi
qAjkwz0kV7kKAS1zezkepTNcNFGEa3pX2ePyo07PrrHkfOnyKdT1uH/pifIbRIgS
GYevXtpe8rLAMWMyo6vHNQrEzwXHSzzAODqFwyRApmiAMRHVQBbIRNf8NK7omI3p
dSd6oOMb1CfYr6suaT1+spIZpxUJjkEajq97ocRLdimb6Qz92RE2xVyvrV/QAVRZ
jps8axfupm3OwIvdnfub/1iVekUhAoU50UK9EtWOcpA8oa2YoEyqph9hjUV2D0Aa
1XWX8X23ipBBfEZMFro/L3iPGz3HJYuoRHgTvPaqlqQ7kf8Xt0ROaNgkmQltHxoP
l3HHLxNUHcyehfq/R6J3nKiV+Ln4gstrAgGp50E8J+ibf/09wgdVNqCsTOBsBZAN
oZ8CfICnx8FnCuz8w1mCLx4KWB2s97n3cAmAo+87Y54MMAHdMzen5LZaxfg2mKkV
AGECUfRa0MkCxNjOkV1xP0bKfsfQzGljghN5hiI9ZRBCVR3PP5e4SAx26+DNNh9V
KbLQ+2HSPTft9UMTQmhIHhd+ABDQWV1jxf/GV3skcD+yn1zCGZrvardhKkyZqkkp
6zvfKtOAWO/Bpot7G/SQ4ZuzG9YpFE4vPyO2Vf+k0TogxCPSW0ZieaztxWrY8vEA
fsenHhZvPMZ+gRgmKTLReds7vHYZQyePdwxS7r5oV1pjpwWd1xU1x+JcS37asf7h
rS3ldfDqw8rK+WWvJClcs1zG+HX53hEcJQ+d3Ra9vHDNwhlnDLzQ37/hy5b1K+vF
pHlFf+wfpxEq/8hfAWLpe+D9g6NZbKwrSwQm+8dH6JhU0Dq0RuIMXUQy0uylY6K8
vyW2QZSi6uxyf7dMsYxwf/vj3eUBNvlYPuzzi7xFupEqHX9rD9c0kQLUC+Jk1waV
BCDJDHfi5pplc8B8r64GJc4ahFCJP5fh4j/vZY9ZyqNHWlihM39nADN/2ML+4OmZ
y8DehUwgAjBDEY8fj8Lff6VOkZC49GfYYkw9X6VXSYh7A1eMvG+maDldJE4fj2JO
N3rWH9tNsBcH2h6SoosHKtUb958p4O3rbVPm6IzzliJg7KSuSrZQQadp1otg0Jt0
nF7TaCKNZBWaUbiRtJ9NuJP0V/J+kGCJWuunmV47LuFDg0zyxkH4SryqY+PYMkab
mlKnvQ1tNLlDClDwlovuYBTXM6rtbL8ACp/M09T8NKCkKrCJMjSbCYAtoVZILJQ8
tQu2Wpo/TdMBIZ1rTIWelAYS07t0uFFN364C3re56f7lVyRJin0MiIrESmKeOY+D
zO6YzCxHHZMw+Ej8sOHvP9EbPvVAZ7HyVnjCc1faO59w3eB0BPmYy0wuR/ALjeHb
p5KU/zfP+yqg7d8UOjCXoDWXqr2TT/0eAxeI5DzeV/3/wyKpvC22Vmt6/LXetvgb
5K2x0Ag1uaLXqFUoGqpTeKocysC53qTWKLeNbXJxdqYxCtxumLjkUjpceDFoemc3
yFhBErHVNs4w3oEA/2mZxXe6zsp/CrI0yj/o4oFieBHqYDJkHQSaSUsoH2X7Ow97
B1/dGmi9Mr39nIMEZfg/xbzAUkNOh6FXdJBksevTfsW3WTMLCYAr/bgvpWasSJ6S
Bv9saZofAt5sAolR7zDEa6an19s4J+CByg38Mw6XkKpmkQY5+E+qMb6ipJCXNRfz
CXbllHzfzU32hpOqISmPtbg6dnb/slE5hfchRT7AzuX1kJdT/BuvUL+fczw7eIzn
A/7WPJSRf8wkPwbEiKI//I7HPubCR42dSSllWr0sufG8PG1/bA+G1iPrT/Bh6iez
94mi2uEzQOJzOWS3sXfDTENxdQsWTY4FcEneIP7Px/KlelhGVnpfRZo7qUxf/Fsp
9JPhwHM43kBDewMJyyyyFweR3TqIVc5F+NVgnNR4ztYdfS2c/JQCt+FVW8+aTclV
+w4toa93tSkEq0FeZjv9CBUbG4H688ywN3sHcq0sA/dD2W1UWhmmxVohwLtmGqc4
YAxuySqUcSZgsbBvptX7CyFd1TEgGj1cvUgEvF27FCxFINYgunuvR/UDOalkQRxu
epjjfwuHGPQk2FOTzFKzeJsqy/ZrNpOEneC9+Mh3O47GHoWuMts1yB1ubHuZV1FL
CZspv8G7NVIj+/wxWlqT1RLn9oYu2JbMUKDp7xGVLtjQyiGyVSj3F7SSujPmvYNe
xvvlxsgbaqRV4gpylZ7whbI++Bq7B7bgXdQ9aG1tom0S4CBTmZfEgxLn1W/SvljQ
ZI2Oi20TCCJSE/fNUFBakZ7dPYlUE7/vVVTNcbaFLbl73895+2S2PGEGu2sXpYxn
gHcEsxiE4fWAwktyYFnbjWvPeULpR4jjY/OahJDxODzdOf7Flp9FDg92yO6e5AZo
sjldLuuzYXdGVwDloI/UBr1RShjZto3WVX/8GeXHfz+30WErrLDpjYmM/lKYYh/U
NFd09fUEauZFVaT9onT2bcw1A5Nhzb1px/g1jUb0tzy/kCqUFSCRKG7mPDhxoaLq
Wvm0hsxjbPHQzWEQdaxHBtz14/d99YflCq0svuXETpwaxamTIHXkXHrlsRSLQyU4
g8ZLPKRznUE4Z3laAmMXxwlj6kf8D4bDpktPxAKH9dTAuISbNIi0+HhNswemvDBo
KLhuYrhXNLCA19qNrajAkD9xGwybGHmwzM6vPS55wA0dJon9i1ntBtvao9Lon1U0
b02XSOV+ssXDr9bThOGgckERtg9TCI89bADxkT4iV2Eurat+4+vn4ugv1hvJ1+i3
`protect END_PROTECTED
