`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
30xkY7k48a4Gaeygtk51yRgDTL6MqNlBW0u+OHqBwawDPIqmC6W3ZEAGl5hsQW3p
cYsvJ1jRKUeT24oU6DVDNiJU6atj5vfHzl91LujecB0txWDUzRt35KqsGEDtPmje
xzCiq9kRRLYyoY/PN0aMmydPrd2overMUK3FpAepSEF2vwMCRnF3CoJ9sLf6nKH7
GljV/ElpqzQYYvRmiPvEURpLU08isGLm6iXxS61PxujQy1wORZDzovvu1dojfzBX
Pzdu3GcPHbCM/Gy86XijqvpAEahSxiHv/UO6mTLSrd8OTPdABmFuml+F3thp+bXv
hvbXpp7oCuTbgBz8cZh9OvFGrEC+gZFh82y4sg2ZTOKEi4sr1GH2DVus9HIEfNC7
mWlIcbdRZte4GJ0ohRWKv1w9AeR7YV2nBFvsIfkZ7Eelpt70okc8AkkQ6zGCuEYZ
nrstL1uJGNEElEfnOscSTYHDQXeKLI1QmUTVO7vqZa60MiE3tw/o14LRNcS3ONq3
gwr/2Gl466gF4eTvaJSbGsEfhIDsJ0EP0qj+eOkirclS5UvabVaIFgXrZBwxRKL9
vfcLVtKfATItppufwqf5E0ai04WV9ylQd53B5bm21refdSo8GRVplJ2jnW5mcfAW
8iGHBEtrTAIwd3AC4m0UgJfN+dK4Bw4UzBZ89jICiFWtHbePt/uWQ/dAfTjaNedi
SU4sZKh+SlgV5K8xPE2Jrukl51rZBDAj2H/6DrVGb5p0ESvUAvVD56mYoGoypCTW
KgR5ix9mRtlQpmRttg3wKgm8IZQZO7SH/shCllS0rdtRXUwcSxFriOD6oL/ZaLuT
LwVF+cdcLfotd5PQSFqF0mHIEkQjDPRjp1W7Kx+fJQ1rorwFfGj5DCjS6BMI70/n
osCdKmyg/ax90Gx/EvuOgbiwPMqCpG1PwZjDPFaukHNO5NN/2ZP/h7HO5LDYyc6k
9uINI/CNAibqrjoNZ+tv6Y3O0BQbXMQ6KiDzzZOLTYQGtNSPlSVr5bYT6qMTcyXZ
d/Yt/Xn3HuMYh67EsN/Q7Lzqp3ELkwMFY89OYc96EI/HgWygUsSe7muvDQYuUIjd
zxAKtWnTmNmbCezy+bz+aomW34+K3b3sxqUaa/rBMzhWIx8lI5Iak1OBhE+/4DQd
UgJ1abh0/pkFZ8U8cDMifekEDnEwPAUcti+5LaXI0+cFRFpOPZlUMkwBUmhzWK8G
FZTMiAnbT//+7bUPdbdHODmhRFBOVCcbpNI/MfjUuaz4pIXhec/eprWzwXAlFCma
vMpudP53vnKx5fUpkUxTVouRIj5o6V6w413l5ISj1u900Devz5SXuwhX1KeXZdEZ
2hCC9loMKZ2Z+2JoWWaNi21mfP2FlySSWpCJt9zjyOWigouQlzsVT+qxkSdm42WO
HaR+ITkwqJZHuZlCv5eIImER1LyM5uQKQPvvRNdX3PeV0Di3t65gpL3xUUh/3ZIr
N/p66alW2/YoEUqRzVC7z3PIhtUzcgP3+JgEaP8JCLkF4WhOx4LIKujmT2R1WJy6
cS3b1AWkXpimt9ryfnYIbgbqGyAQmTgkZDlp5oP9Zopp6iRznqieYTs6bg5HJ/RO
R9oKySNaQZe9wz2eDKkMhorzPxwqJ3G9kZlrLAod1qisK5oT2bWWG67SiAbwlNIa
q2wjBB9EpZ2rTDHNydcWHfIYpBZ2wXOukX+mlAoI/PpqJl5qKTtKhR8H0tqdhDVy
YQxXH2ahrl6EAsMctPzVqAyGwV26uCtMBZ3C1LJsriYI4gcCa2y3aUfpUdLveQ73
YaFOX74flbVKyn7XEMDSZDK5nKxVKmhky8i6WLOAz1h4buzOpUimd1bHyIUGnesG
22RybSs73ntLtRHBKSAzg2L7j0H30orp1QclxM69Bv8BfPSXa+2Dbar6dBpwucuJ
pnv/Pu71kE42k2HhfHB6gmwazdsZ44w02ZG1WMQZ0G7QNHTybVCX1a59F6EZeWhD
L5swd0aGeV7kutnL+LcyEFlJ1rLOSAYBxEjw6RtX13g3RO5TDmqaApuZS1iAkqbg
VL+nEb+Hquzb2kW9+eSE61HaAnqUWT9PMbVy8TqRbMlLVi+o1quSod3aD6knxxvx
7SZ5DjG8MpHvym1J+ylQtssZqQMak2xHgKEqrowznio6/4kQvioqnPTamc2S698G
sqFiuFxhviljNoSS+sb/QIIBtPPQViRrIs8qqvDu4CUncOG9LH401VlDqqR0qyoT
cymm1k28kBdf5SBXiR46gV3KsAg3pG3UZhWEl5gfmHtavggql09dTrArCjPTHUMf
G69FXqlN1mxKH5oH45O69wt8SjRJ5iO8DTWrPR0m0Xs5sSAG8m+XIRfWPkzzR8jD
XutAWfT05ABxQaCHMtHLP63j8LL4laAtKwuxaxDfgrAgMQmQ5ukfBO64Fe9xIx3T
27S4bBbQhvLWGPtaTwu0JeJGST0PXbvcweUt3Hfd+Bl1t4d1FihdqiJIEPR+B9Gy
AHmvF9kv8/Z0t+oIk6ps5Runl6o0jUCktfVITjAq3xShs63coUpSWn2PX/RXFtX7
4Ddhi2crsgGxP0h1Vn2uDNw3mgnasBpmVRdBT7Jzx/w4rDr3TnL3smliw5q5kUVD
7G6mFg/hQmscBu+/VGIOxTsxvkyVJgOxb7qxtywwhzh4WGwQ82fSZ5LliCPHc0Dx
+olFLywRSoK1yiAV8BGykkmis030BhGu2MyoDRRyRJ1sUoToDEWH7phqSJ4F3WtW
wPCi2i1XeFwXbIsNe6EDmd8x4sQzxQ1LwHj5cUDRfHAUwCWVwiB5893AThAqrdu5
OLr7KNN562H3ZIcILTnuIT/0iU2XZ31+gCbgKns0ZP++Mb8DtrEVD7546s98hsIj
qjF7l4Hn4tDbHDSsHxj9qkZ3TFcXZUjdv/xzUZQKtLPLBdN0KgqOclNayHCyfLQZ
HAuNyw0QUbwRMjgMAoHuz7SzeDrpUUPwKAMh1OE/jRdbkvx1SkWPu864VfpbfrI9
JaPICe4LQkub3LI4ZFmS8M+ngMQaIZSQXyUoty1FoQxV9eTdywt7uPPSg59BCHBu
ilXQ1wMu59xNE6xEghr3tK17sOChPhYHJrN3W66VSXKUYwer2OLgcC8CVmTNoBrb
jMCg29T5gPQ0hbeBDjpXuA7LiegamyE+z4k8JvIV+xw=
`protect END_PROTECTED
