`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CHSwJGQpcWfvRyWP+OVGpOphPm2//L/RgBOki4cPKlfXPi+XaAltpPZG0dABOXKm
ymEH2PA5ypIxYXmqvKbundfe9Uqz86RTT6n0DOryyYYzuKk/ayFCQ9RprGXqLa2r
PIDIYjKAcXnK8u0KZQmEK68bjqpi6rUmqYcljeS3prvuEk4v6E8h45sXRbv5xqUy
XQTrgoVo4AO78u4WsQ3XKKSW4hnqUwM24Pe7bPrs2QxPHCp49kXQVklX5OTIyl+r
GSruTKSY4gY9gsns/rE7ewe3zoRUw2ApAVv55GKT+7qMJY3416AlWEvp5w4kdhYY
kVHh/5+jzANGe7GmIR05hdQ80VcgJzVxSuP6T65lsE/NAW3TRE5O7wRaBR6hNnRs
BBRqzqy2129hodrNufkGP5fuP0TY78RXE6iPFuvjfgnysVeCSvwMVmLXzb+sYW8R
klxi5PSrh1yWCNeU9hMqujV27OlbnZ6LRL/NaFCQ/YcAPqi7M7ZfoI/iHJfM7NTJ
g5HkCWQv+9u/uV60CoKPHKcQezUOG2C876oRX1JmWEbCIrL1pYdBjZrgx7O5spmn
gJFcMdK3GlSzK3bRD1JrjHjVDXU8MFxOdz0+iOxaD0BWUzEQjfD6sXcQMEpNBWFe
I1WmqKGnIporbvXv6MLaywP90SPI+zoFrgjFyaHnESLnMozmwYpYvGHILCz1ftTg
AY9/kMgr69eCaqKZQXU4n6BZKIDqpTIgBy9S2g79rVtkRn6OAd8iMQu0qWnNB3fl
`protect END_PROTECTED
