`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h/WRPY61UqNeCEnx1lO8bhjZnlj6YdRO1UhCXbfEN0pMSoLzBkx96hm4ChS7JjD9
KYXwz2H475NAs4n8qiiyNL5pgJnviWNg/Q8xXlomUN65/ARz9LSRDrELihD5lMEB
jSKBGl79kPQGl61qM9BAG0fLPD1ApkpQwCAzMSXUVUH+yxdIHk79wp8KPjlSIg17
bLTeUX1xt41quo2dP32G1GUIj3dcODy9ayYh5eEiA14kWwcwaAjvSMNE/IL+S8AW
DuJize7iUKfRah3ti8P2DihCRtxIyxNijbbLeTl9IuEqIQ2RWHqHtbMttfPTT8rT
fNombz14OoVvjJ6rntmfhPg2Ut7hKcCKwyPtMQxhnFmVoMYX/ajuapRBBC1S2j8C
feudJLCoz4yDqLY3cbxGK8jaQSLSj1izv4fmu8rdssQfslWjXYcdXFyWNk3uGm/C
Jv7t1cAdJkv/bj8co5F4VLC4Vr72M5E5RLKSAY9mu+2bUz20xC60FNsCD/Ileu/h
elAPU59ZvqVMBU34ypwybCPZXz0KceBfHMeC8Q50CsOrh+bYSHu2nRx+w7fYHyso
8zz5/cok4RAoIgyztI0SMnIs0fw5dkP+G8LotmTI3pHym1FcbAZ/BnsBdVjjYB1o
d1Eiqu1hmCNKIykD2nG7HkIpuHB8gzauKA+s2J0TRIw5z3se+UwJW0GhCuMorQtT
luHYLMkojmf43d6yYMNtT5xT3p2samfNLgizQbxpSg4yK76U20fo6HjCNq9eMWwr
7GJPUUY+TYJCNwANH95SKWkRqmNorLKjGtQx5JBbFAU=
`protect END_PROTECTED
