`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XGaij3fwcBxnpgckhikLBV1OfSObog5q4mOAKdWlWKY8nuQL8hw8EL6ALWdZqGho
/g0NEp2RNEPXx3ywin+q75Z+SAMGIasuXx+vAzzqUb2pYWHwDGdLpsyqR1ujxCMN
WBUmkrcUixH6m9M/+M6++Ma1KQuIuoSF4/BPiIQ8q8dooI0L6a40o6zoHA7d5QmZ
ZGSIDPC5YXoZSE+itbb0M4BT5+dFUzGxuFUPDDb2CHQg/HMyVGXaVjqW4jfbp7wX
oln0U8CDc4PhkUb80/tz0xoleA8Co6DmHVkk94f8YMZLT2J+rDYU61j/xDspK4w2
3RaFyAbYfIf0rl8CYisGXSy9XhnEyOTclqcRuthIwwpehaMNgDZXYXIFLOSv4xpG
N0q++KinOIwpUs547R+8NRcB3HqqwbWSGLpudpRn5Gy7rOqfkKuX3igvn6CwOGxZ
dlOJWteAD2AsY9iI+rPky9BbvBUaOgqw6x3ruqMs+nsH24fjzkllPpnjcoW+BEpz
dbRN38EEYGqmpdoMHuZIO9/5B1xb0NfYBV9htf3JHBmCTRa5MJQ2PK2TjPvnVuYT
W+0uXptGLU0fVfn1paRPS41HgkvKtrTtXQovd+JI0cj24Fhv6pF5/5b7fZj0SAc7
oV9lUagM7b2oB/gEUgFdAGf6qpni+NepASSxdzYxvkOp57P9vCY/R0AGgozhbWEj
5S4uxHjqdlt8osbEtEMGpsXKWOX+jkBCRvnZpfwIFBMalyGMnOTg91wN+biSENeN
vAhKJM+BWMLk1KcHIk7oGvhAzFrZbqqjLdbxJC0a6/H2JMqwvmGyRQoeCyIQlTPD
rbw/Z6nsORG+q8waRMPmW28tZETWFC1gumS6BYHhWsPEYjIw/Hp+H5mQgwgDZbcV
9dbCbI1DgVm4ecIf2bc+VaRZ76rbubgZZWi6k12rngU9M1x9J+d5CgAng29m7v0h
`protect END_PROTECTED
