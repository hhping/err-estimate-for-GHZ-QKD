`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s0ryoprOxKhZFr6xNzFdYNxrR2WSNOXjt8nQgEsAYtUe1PPpmva7lq8wwfV07Ots
9E6MZ8xc6NxLPj4JMrmSB7YX4zgogtVw5gZhItfhgkHyYyKHjGG078otzdxaLRJP
4A8Kidq32QlyQU+2Qrq+1rWq0zTVF/PxMQr1lP63bpaLxOvlJxXntTJRX6159QMY
0JR1wOkCnH+XmGu24F6hxbXu6wIvYpNzPx1ie6d0QAhwcTOUcRqlMRm2cbJBe1TE
2dBc0I4tgFgQdx5U7rtng/nLsLNOSEX0ookffrZsxphmLikU2uH45C09fpPq/aHm
fQ+ehuozi270XdRrnCXOe772wexFxw1EjCTTHq20b+OPTatyYLJFwUmLgHaaS0e3
kDACB0fh1ArBK2V3/C/xkCsyOjYel97NLfZDveoMrEeAXR5GC/T1D0GHsXPqjLwf
NOEiRtRuXfsjj87dmt5pzxgjnhVkY4wYZS/MTGuPuBFMBXwpjdzsJcklRWkDmyfG
NAXCxpCbtAtEghq5/BcHxdZU7NCjFQvKw5lGN02oaL1dlvIvC0zVg0J78AoTglSO
+uIc+10fG2nCt4KqD25ewpmZhaNV9UtZARorDf8HF61I3rvBNCFN71UGneV/Wtl3
S1N9YrqlE6feG7YEjnBqJSPniJSHtertR7LnfcbSoxRJ9e9mHlmmMMXToY+ALsMh
bZFzklzRyDrblHL+s29MviCnqWxclfMc9TUY0FUORy2US57JuUkI7xkR85L4zauA
ndQXHQaHOuJhHeTeqMUpOZBfjKuyw4/x0vHGXBdrOOo0ALWOp0y3DBbFwFe5mTMQ
fgw+prntVJdFfFA9O5S1+fKYX+0nN9+L3mQDGv4dpqFpkJRdhDiOngwFyMbD86zz
QCfg0ovM/7au5e5TuWn/Nd5+DBfcarA+YPPDpwu/+Ae5Df53W/omCZrJF5LGelWt
mKKjQhYUWgQhyXB98J7QkN+bhFjvH4W9YR+1JTpu/tG5alsBhStSIy0mKRDVQdiX
dZHmfshtIQaXkfhhV9OzwraSR3isKqhJbDlWsmGKoYQxtY2/B6oF2Ru4xlIoU3uo
A6WDWhcQpiWXYMrh8XHmeap8bXkCa6/tqNOh1231+eqkbg7nOLcTH6eN86cMxZhp
1FWWIUaJP6dOaT8NqXv68GY7CnWvjL9FeWOvUIZnilnbz3ZP/oqeXckuLMvgiYsj
sXqrtVZ1CIeU7EYVDs/4HfltzljU/t9d58SCzmM3tJFxQdAOlu2XkVLvPzmKLDcv
Ru1fnacOv+QxAp/eOD7kR+KVslvCsZEHJigtNsS2xy7lcZGJsJbBfRPbTjedF0P6
0rE8GLNEE6iGSEpisEsbssr/aAbKPLA094q8qh8foULlymOTIiN0SK2Z3REp7xAa
lW14IDmm5Kn0b03ONaJsspoO/ZMbO7Qo0u69+FCFTCxHRfRArRTqX10nchaQ5ZwV
Iuudg5rY7XZkk3BGWn/5a5R7ppGtwa6pfKQw1bofvbK7FyepsYgdAiSRfSwGsczK
HQS9Z51jXegQp9NSZEunRyDsrq+VFdAlZB4uBqVZnPuyUl5wTbOLoKGbVsJCkoCg
6lXBV4a4SCM7/c+2sxmQ7Ek9OoAhYdIhzPYDiPa3nhPfoKgnKZBKJNTS3h650XJJ
JM34gl3vFYxSjTlkWauUlQ/LNWePWGNllIymgJqgmhHsqaJzSFgAzI8jpsqFqgdS
1d78lzT8WomT5ogAn5VXNbHUJFsv0cwa9hj+EKRZBv/u9ckcbwtNBZ70K1KZWFxE
sS6i05MfE97HUCHODmTsgpJXBdo5QJcPJjz4f4Ob+1wPo6dsW4A8wi1mKQxoAj0A
Qru6W+czUJT1FI4JCeBcZzpPsHvkmIF3Ky6pDVY9WISUT6unEjlkRkC3YYmBVD1K
XCcbtkuzpso5NrEyG/JrknP0loEIvQxY+2m2SHClAxiEx1Q4sjCqWRXmg7AxIEK6
oQGw4bt5/U06GAuUZ0E7TCmddyAQk1Pg86bnUv1BKUV//RK84cz3iCJDhn7Cm7Oy
8IRdOV4cL5XDr3qWngUJXw1CofVzrwdMQOuzTChiqjmE9ATKYRuBvtBAYuVh0NXK
cAQ0t1Ccm8dMJjbKIMhPLD0yCG5pPLJ6WDXrq1htxFYoGD15CKxGlLjBUOTj8NgV
8nzPy1RWvesMrAxONND0EC+wMOlYwdeYrkj3dpjXb6iKgDf52hJ+eHdQcNxyldMH
Fx5gpXkjSKmtsHuupqSbLFa9KRpGaVpx0YWNyG7mTdUP2Pi4dlCplVSr746Nfp67
DnEbshITqei679kcYxFzOXg2K04k9rVSR+2cO9kD0Js0S8JZTB+Zd2//pycR1E//
BeWvW4kaHjIrMEt6BKSerMJ/OOMocA1k/oXOSReevsKy9BAHLpFR6r2bVs0DKIlh
n5oOglyvBLEcdk5sik0byb1hfzJBqE9mOYy3b3kbel4wRWliMXmiJMgW0xaiR5wU
nvJLQB/eJa6haL5+mvbbVUOjZbfKcpe7BcXAzYsi4Fdi/JhdGcruVkXEy7bPVsqP
s7dEX/7OIKMYJx+tZ8inuU4Bzdop9qAJdSYINsdxzCeRVSTn3ZwKvAXXa1aIwxe5
mqOEheWtB8zdZmSnDpCMqM0Mco07Jj+PP14/6JWHFNFKGij/B9zn8IuJEIbPG20E
Np3J5EcVE77RVu1PzG7bktWksMowBJi8D0bsgEIusQo91RK7kwCyTHywT1/9Pbk6
TjLGHqeSjh7pk1ABblkxklvrahHmgIv8CYW0UCxZYbXpD8sTjSa1senAfWIGlav2
09v5e+mGW+ql6ksfcBTY5hkr4ViahO+PUXfcjjmAr1uO7VsWzspDFOH2dpwGpMnd
UuPQzSuzOdLT7+JOlXfEz6RiCb70TK8p8JEjkITjvisloThP/sqQ1hCseitNFYCU
pefTKgvJKffi2XHzTC4Q7jWt0KnAhQxZoph8xL/ChSjDWZ0ED1rD1xsltNUdBhlA
wytLcnAjkZhGIxeYmF3vTeNr2RFXBVVmC68LHxX7Tqf10WRYcKZFpVqeaL11P3j0
nIt4BG5VAewtdIBoip5WwwUOWuD4cATVAR6T0bJLOYA=
`protect END_PROTECTED
