`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6pnl9S7N+JDq465GcoiUDAZyMzO2iNJLQ6wt3PxA8d+rS0AGMgFaB++rD8eRBMbj
e5BLxCIQ2UHAmdGWJZX8P6CBQRp43XMULgQT9UgalkCrAuMVwN7tNxkeFr/ufcVk
TenZ0T75LrJ0Bh2/1H80n32LQSeKcztkm6WgC8JVHeWzC1MnVVimFCbDOx2UUw5B
LEvTPBg7k+ZwjKq6jw0F9eZO4RgxJj76TXOMs9fzZCg9YU7Kk7cLDpY/t7UnWlJB
dko34+6sr+h9gSsdK56YxrRAhqphQ9GD0jr8CByjk+siAub8i1DMMpB6t+/B6GIP
XSecYaUHEODAVp3MespcWiWzE8+DXpPwgp9cYCgRFNEpK1pbRPN26XqJ2YGdCwox
K1xjsdVb3QzU6W3Jv2vb4R/F/rSFlZ1ownCiHrHTNA811XGO0Ri90dOd0rs07/qK
jO60lASSMy5o9iBt76/IEwY2CiXe32YNvKHitFkxYRv7CdQG+BwTDPDsrDzlAVTa
93SEFf1r3xdcVypfjS/hXDoBp7t2mR8QvxT+Ulnd5hEKhL5Xws26PIv8xtbaY3E6
wKz9ltJI8fcm0cFJgs3VGY728zleqAH78ko2QQ7fWFybOxcw/ZEzT1MtAdZeGHj/
+JYkZR9mxjJAC5A59S872KYcIrT6Y57yx+X28PDQRHY=
`protect END_PROTECTED
