`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w3kUu0VpN7Q0fdx95doJNqHY0Nr/YAggGrs19DBnnz6i0GRV4E3CLIagRrrQ+GlJ
Ajhe2vusJ+HRVXjgzvelQ8ZVK2R0I/9MMSiQ76j4sJcOv7BN0vRxnVlUpvO2oof2
ovLWhIK64WEBDeq40H802DblJbjupm0NnTZlApQrMAnq8aDSleJ8YTRZhzqyDlCN
BCAP1mI5weoR7Q/5GDeV+YmebHWoOD+hYia2Bq3fQJ4Af5hYjc8ud5SP/wIKMS1g
VltLMVlCmbBDn9QMDs+TNenABZspseDUl6yWWhPeNpp45qaRBKIIhiLW+l0B3BjB
4E1LDL/NVTIzmgkia9c3wIKBHwE514KQzwAzTUSFvDXD0zgYbcrCbCxIZMGx0VyM
OmbtbaI3HUreixtJjh/KBN1kO/F17MVB+nkbfJMOQWyS82tDGai+aQVFdANJRKEV
WDIkSzzdOCAs1H6lpKtx6vJJYlBQPH2VgXgNrgaJVjzvUotYuOKpJZHyYN9AByHQ
oXog/Yp/gJEZfkFbhTJwGHpozP1IvMEh2KWwTfKKwLcYCV3hGtDe+hBdTh/wxMiF
QhvhSXTfkCjv3mMxbqdqiMLCBvi2WERZZ8Sm0J2q3teyW8UxJVbj32Ayx8hS1Qc3
+UfGj/KZJFvT69C2AKGB3LDzeXW6a7RGnATZwgn/TZeVPbUq6T6GlsHfJoZReiCY
n4zKnuLP2fIq4sVHEYWDD/lO+sWQEyUPLNOSogZDXjZbok50kOZF6Ra/wyh18w0G
eUB7OBo1ZcTwjFvIY4G3FMPBEOuVQqAFeXNLO9sobeMXIrWGVUAhkyctlavZDJvD
ZJo8J6DeLj1CzCF0KBPNENFhU+W6mK9L7xcaUgc4fgLqT2igsfvFfcnUyfeOEsyd
idWHbLnzSdz7j8P1gxIry23ngs/W9HviEDJNTyXmsMhpNV1ZaR0hFsdNH5y3KWdj
q1z7JTqmVVC0fSzri/4LeLm7cXHUhfDjTyGP5SToPBwsIpKsx51dZiSJOXnYBrRi
+APkEpjyBjrSaE6cViJyCUpnFCv8243LYj5HkcFtcKh5oc2LxpTco4U+mChpa1JS
upohqo9gA0WxCSKFL0lQF+76mXJT8pfP+I0Xqm+hHG6ZFu2xmCxiYpzzQBEX+f/q
Uad/6kkLf5kPr2KIwpPaZRLQHJTyYkNkHfFAvMX47I0VE5UnXv0nxdcW4heFzrdO
Ob9cjIFJUE/AoTYLmBFXGSxVYLA09orQEFMeQAKEOflB9jliqDOHx/u5PgzLGILo
tWqrWKl1+wLqLoBe+WjxW0XBY7HD6dVgRg2NHXkuXqVftS4qCl+ZgOZHOcfbkJef
LbgtK6p1ZeM3LYXkEK2xXPJC3EFBuP1gNc7x8uYWSR8lqpfk6HnHmMpF3QsQw9m5
HZzUEIcJjZnEV4dTdsw7YfGj5y0qb883MmeS+SdqKNjd7xawsjUSNGbQTdak9ytq
IxbOTxKEm6oN/w3AJpbvru0eIXUNt6oe2B039oBRfrhuN//J1mn1EZabF5YYTJtQ
cxpbp2zTMPI+mVBe4ZUFhXpTcgcun5bVBJUIyQiwtZ8hNBQvvr+K9RfAWu7ctogX
bfD7k7nzgxNyL9AppUh13zlm9y5GWiSOXjjpWbJ62JKEAOb2eUD3VR/VUIEbRGHS
DSw+0wdXEc2Zty8uYP99R1A7U1gy7WpsRp9e665zm/16tBYeFbJuZtKoMmsyn6de
OntEGLHc2VRFZILa3NHN9LGWEFQmoUTQRHUF32+Bonjh1uvORU4N6tka2gx/mg6O
43Dwq3PR7NpxcmRWNLW8/2FjKaq6GPUvWFFsKFWBla0ITEnpuFrP0O847g5N3HGj
b/l8st8RxAU7QoIGhCvW3eSJEleDTd9ewCbvsejYNkvwLv4K2Dqx/1e85AHU1Wtr
SqUGPbrD1QNd7wD5yNBV9/B69A7dsCCin0fORbyf4kDxeQEWiZzCxot+SnhMrJCL
yX9huf2ycccdcqlrYRaKfWjBcEty7Vgfa6eBvCP5IKW07e3PiszGLb8yM2HR51z9
/nRVsDTSLv/OB9FzA1e7XYaBnHlkMAWhd/9B0rRkIxo2z2tzm3EKWjJ74mDxl8sO
f9UUMGgn+bbPc96C/ydVVDjF5RoeWvzoaAPSeNNpDMPCA6bpnEO73luQIbik+WJe
fIyPaUshcEkp4aOYI3vnce/41Hsnw7WP87saAr5m8VWF6mIuLtNQywvvYAyEBPUB
Z3eNaIYGsUe484avwgK3ElUUADZFdmctP1jGU6IEybqqUJvCzmCE65yCPOKdS1ir
6k1CXQ0PfK3D8jIyePWE7sbuvtvfa1hRj8blUO1XOCKjBG5skdDLovBN6bAtosgC
Tcwk/ipRYIn+n1SxaqDJnEujCm03PvJsp6BmyWfc2r/4A9dSlUkJEy6QMjlkrEq1
G0vj9J4krWYfwtzFxqYI5EZCYUAt7zecRowsnLNcDHn/4Z+VB4EDwME4Rxywpinz
RinGQYyraCk9IgM/X5xz9yBQBfseHHGwov7LiUwCpMDZGJZt6szm6o5UpDVIs9qv
78CwFViZ9DHneYMl835nC3yLq+YQBNqCpy7yMr/i1yeHD0nxlDIO0gR4fftJj+11
FMj4SQ7hn9rjQnkesm8GBu9Zg4feEvbu+eD43kDXqRyndrPhy7EJvcY7pc2W+BzB
zoZBcKoYAM6k6jPc13oGyJilfLR/xjkX/dQ6rtp7zXT90aav0OSagVYRLDDgUOYi
hxl2rvDdUDMak0V7k/aSz29V95eyCLzaHt2CIHTs0W8Le7J6YuyptT14hSiKgDrp
NAkbqLa7XiYuVZOvLnAuDSaobNsnqFdj459RnBkn6ngTnjCJDM23V0Dn07GC6FaM
DqEgQTkbakVxlozHNiLwAYVGRcGxNmcb+UE4D+3WUkB920AfrKtcUfHOewWvkGFf
mqhh1l6TUDyU1vFME55ifHZ/86mh5/UYcmU78GmcLdG1L+4uh9aKYG+iryieQ7zk
AJpqLKKQvtKZdKudspy+Y7Dv2fCTwHJCcUz0+eLUiFr5RlbjHOGEOskdVYvnx+g/
v6iFP/etBa/d0L0rwy0YOk5oWMMbfwqnpCFVVmqamC50hV3jAfl32GUXCBJ4WE9f
HgYHcl2IQyVQWI5VHYp1fHvi671tlGozGk5wVNuJbZ9FoUAxRkK9DN8G5fjIJaWg
1i+Y4PJHnW6S1SqXyZkZj/+NLujhoc14GEzoMo7uGL3eSnvgBjh9WJtFCAieJSUr
tCje9toC0ChVNOO1Zi0ctb7HfTCrzb7Gb/wjCi1B1e14TYTXPmrRUBbLSypsX5HM
lxc+TXWPXBQgzYvaSD9JuohT3NCVYJuZfQmnMPNKJWM5hWScBgFj4hNzHOCnFL1+
N0eKpkEHX1kJ5dZs9xHxuqqq09Y4uE29/KB32Q6a2sSzr7TWiOvHr9pVNNygZoar
H8pANNTFkRcnUyd13p3WL5GGd9a8/8IsgmSPzvKNtkTak7uLVuZLv7Nmn9LvAt3N
ZUw8h0cdVJf7eR6BY+ErOQ9wKA6+S3C5kaqaDAEkTAPKXwew6ox3yoTg2Vdqnkyd
sxRsOc6TxbxUq1yqzTVm1xeMMjvjxpbBIiMwUZA+OO287m6IDHQUuytfHBv8M1yo
DzJXHy72C10Y8Bb6dyzRBjqiCnrkTJ4vxVmBoVdWW1w918ps0F2fFmVOI/UDtVbY
E3zYGorDT4c1REtE4Nx6H9Z9C0/mHcfjPPyM2qvT00GA95BQQ+idcSENZvbiqmtf
fIGJRuSDtJfCuj5izVyCx1Atf2hXJUkFOiTB0D2Iz0UmnbLzZJRuHay++SlFYOMB
95i6J4FIqchIbvw2pIuSwGyOsY0z7DQtQlLyEV79HXieRZ7TWB788g0zU8hXjJ16
5DCLQBDjHQp9ga6OAwNIqNyrvPLAhutYBqjzZZD7z1P1lEjP/sEbo8te+ghXKPHW
JMjleRkEONXhHZQtODNcPRo/SaQk6AaBaYrJmwZF8LvP6k+norEdV04RXuLGx8oq
tkX7+BEMX9sJlwSgxVXqamMZej5LeFgUmpktTTKvliv6/XMr3waci0/l5VAjYZp+
xShxRLVOYh8bziHxjaZUVHNqp2s3vuu5xreWI8MgP94uIXGQBzjr1ZlZnPsvfanS
mHcrmOMlJnI4hFSipEigxC0TDLl5eDL43vFJ9kRhFLmgtgQhYJeQRhrM3V1lzpPM
o4mPCIFT/yTNz6EgQtv86xtzsfi2Emh4k2ycnmWaTgCXlmmFhFXhkSC63BzultCw
St0RJT9QKF4aivTMR00UY72f4LwlI8pADYvORr11aKUMjEbU1o/wQlBBrsOwLYfQ
Fbtjy3iGbRtiAk1Yf49dbNxfVD3PAvELytNkKB98gbVEfXhiQhlAl/hExLlwNT7f
CtMo0ZYG7zE2oF9GQdH5U6b92MGWWU5XeKruf53ELeZAekJsDMnhGB4LsUW7SEOH
6TltzRKRKR9DCENloNmfr1CFDeGeVDdYak4He6LWtEVb+kgJodGEFWtHNmvyq0SZ
d3Nej7ODPkx4j2Kx8TeqSJA+AqH9mrireFDPu6O9S07cA5rIyjZrkCkeuf+6tobG
JudDxapOyJ770GW2UAUupPC+x23Gl7Atp+5hX53oKC8ITnwOi7cREK4MV/j11ceV
tKWGGIUePWQcrJKY974i51n0XdXGW20JBGMO/y6LCoob3fkRHTU/aWRjltRS8OJe
fjPhF6/DfPjRh22HkxSfjOXFF7bUDgpfsgySWLdmAmhXxm9ZJRlNTgMd3u1NSh56
GlGdSd5uDXetlUo7zFqUWAbbTcWx7udWV0ztgAoeI4EAuFZpE5121y/gdRyZsbaJ
vcZPhb+FlMaBhxxt/g2pYb2qjUs8ceIf+51nVWAK0Z+kF6Z48CcOI+EIR6Kthm0A
PmoSxoD11ezKlZO/KdSuzswd3OlztcdC2NIASZ5eVaxMRX+J/eFoba8+sOWJvLlw
HXzzqPssnpvmBnlI/HMRLDePMtaQm6047vqEPXX9uut+VElZg/XZISpDRJWI55t2
hDSxgitsc6nYDBIiTXY7YbSq4qBuxQQD393J4Bco/X5kyi+VmUPV03e7h80TyGb2
y/jo7BRUFgxUMlHQZd0961FxOaZKesotjiSCpDsnVtmp9k57PWbHTpefqCEoKCkg
1GniogQnN7nPB2cFEWGh4zRTdgfuR9c4FVGqM0GN5fcUU2l3ud2vjS7a4QYcUUPN
xa4Tvmc8ztZq5D6VxFHDgxnPamuICDLm1N/A5b4Bs5q848TvIzaduHbyAAqhHyWe
qHp8XzrP4eCc1FywNiODCjUwwMeF+jK4cAduhwap3b7F8uylRKuSMOt9DIHQCbvf
k5FnmUSfZBNBP0xpLR9Nna+F8YrVNFJZUhtC7iWeKOWSEGl7RpyFAPMY5wdna1mc
5y0OstY4ROyX2k3vix2WumkNOlKq9IqIrzjSVhs5ZB/jFGLS7YE5D3YGVIudpRx8
Ow4d9z9UdjG0vnG0lzHb56IpftU6LYVPN4CQ+3AFjM2W5hc8+SAzT+w05AwCXiDw
KQGA3HXqMkMhCjIFkNmT/C/vfQYqX2Ks7rNwCauF4j6OmbaKdlfcbud0MoZ9k/Gs
7gcc5O0ZS2c4pWE6CcRKQK9Pe8v0RCrdPvVKAXggmgzbICk9ZKEMTSiTFO4dP5Fz
dR2W+G1fmOdiN4Z9scP7esShlehMAA2epFV8zxgOXagOMlvZTx5glRqa250N1vWI
bvcr/vZwrZ36TwG90wYRNFmzuzW0CARsQHOrV9Unp3fNrVJU88FkdbVD1Oi01+II
1A4GwiQzQuq0ItkP+rS7h9gNTBhW7lTS9vAtqmkHV3A/Xn98CHEX+kw7D2Oi6N1F
fcBz4uwcGeCpjyBvGlf8ShcSLT9lyFAzSuDaUNSIUdVlsRO4UWgRNwGtBpYM0A11
PwKER10dgfAPLG84AieL0asMPWhFVO1wWdNY3+2NWtGM8JqgFPvRfCILQEdGJuuK
N8ZBu+5tK0lgarihIa8mtLWZuy4e86EZGiPDu13aQ0a2dgcfLnEarosFAb3u56WO
Pc2FYdUUzNVWmBlZNyftOslFPCny21lUfK6ygLV8qDp2JVQMeAB5QtVYy/6sdcup
Duz2avWzU/4DzatvzH+FzMa1eMVMZAVdsNa5KR2XJdLV8nUtdQwSh+J2vEN9aX2+
xt+NR0AscSZ9Dorv3a2jTaIce2KV0TGa7vq18BSvPBaq1aUlQX6IssYvAh2FJggd
UsKl/qacZNf87zJg4u5O+QiDLmPPxaw3R4Ha37REIaK3Kfoe2/ZVNPWAI58djXpS
JphB+87ZmQFa8NRfnpXgijDUXHKnJFDjzC8FDsxpCtBZGSI49agw1zpk63WPK0y9
lAnlXqQ2P0NSCJvgxmvaTyE0wvKwdhOihCF6WHgizhrTMhZvcko5gEZoWQg+GLcf
frb9Iy+Y6FwimZe9+RUOF4/2Ogmq0C6OKindjCPIf1IXB/7V5cceAAr42iK5q/oB
63jQIhC+pPnZXXOMqfdsjNT7E9BoVmtgeO8Y8EIlTmGJVhO6Tja+bcNQFXe2H2kE
q30MNDYcRRXvUdPcs9Y5wE+lofH1zWWey8jcCBNNuvyboHZUCh/FC3ToWYJki5o2
FjbkdpTezKGDefT004bxaVochAtEMS0na9TT5XapGxQVwTxL+NqmWE375n2TBqNB
lHmuEw+S515s1Ajc9WSN40Yxd5s5O5kL/+lFh1GgdM8DijD1xWVIbL9KppBWEZsS
oT/fkrB08L2JxIIUsHfW5HhHXURYuJ0Cwmga/GIuAqU0TsWqu4KHky4wzFAf5FBn
8yqC9P5QppCvnxg7IOIxqKJnP4MzVlqzfX/jV6mT2g67M2Y0uKhZ7fiTtQzTyCxM
Ej3E/jhBZ5KvI28x+CvpZCDlg7Z21W6CZ9RqPwE2wkkYHAAVglOh3andDTiBF41H
Qi8t+PYfKO+hktIFH96NvblUCH5W54cWNbVqW3Qpg4iMaPvVpET5d0rxgj+zTCFI
YT5msdXlrc0tIMPCnIIZ3pB+fFDg/6W8ynr0hs43KPt6cyiW0YCw5WtzvwLHInli
G7rcDzYYCYfBFvqUgXzf74tgstyv4bdapixSiJCrZZNH/91ukRgKFDwn/PexZJC4
r0Rn6uE14Y64deW50zVO6tVmUpqiRMOh5/zm4izkU3kHKKvNy4IbCBDoS9qy+Laz
g4Wm04RJYHALwh69WL6PdqncaoYws81lELquwH+gZ/iLAFWI2Z98IWqsGnK7+3Xb
Dj+cfeckSghiHXe2VSHbQiuC7qrVHknfVtXHbFerpNe/F5tQqAbkKkGOIO7kHbbH
ZsIjRJLSm4wNVKlGeVYcWBLrLpmjyH5chBRNxyBJ4QMgwCnvuzd8/S2ES7yCpPse
SXYWPNN4KTvZABARYzi3G5w/6oGYyQLruGID5BtoOqL7oLNADmgJVQw6WISryLVm
JY/TemhVC9j3GaydhnXnLrZItvgGUlm/gJAjfB+zoRNrQLln+bNBCjGTMGt4gKHI
4qI4TzJy+sbzmmWmHzSo7317f/Ga+tJKAlN91lPjo4NjX5wAaGw+PId9KR2n1cPR
Kxvdt2/xKI6nGQh0+mvUoCrezlQbFY5QOo9x4I7iLFM9RBPgrG39yvl5EX+xG1AL
Y1lgqNH/cjHKBI4lgOplo3BJN/seJgqTTemBqOBtGkOV767V8Lri6Ek70PlzM1rg
lRh6ZemZQYn7LiHQZMB6zuQjGOjF8MnMjN9m7PcmLjSI+xiJQNvNEbbXsBEzFwH3
NpSX8yaMC+g1dV405ATa9sFAJXQuCxfemvDVUSwQvL8153BJ7bzT/URZ8ixkxOGL
pL8dh+FxRYdZ1HcRnkscCYp0CwShNW2mnE5BfpuCadRaXbnFxAbrBS/ZenkvBsVq
nfgfyItgPCurSermcPkhzMN7p6u6eNl7yv6sFShNGjAkhOt6vHXR5kHDhA76WPM7
uVYs10yx1xwT3r/8uCo+JOPK7GvEFwd4lMlxhK6v7+2xcyIDdHQMsrQ0TYEixbV+
WZhZUk0agdDJGO93iSaf6mohu5hgxUCOGxBhtWdfuxKQaCW/PdLEYm7Omzo0Zb22
rD5TZRLur+8HyqztbM7x1s/APiebhgxchvFfyyJv4HaFqDiBt3uWJ9dwZ04lVfaQ
4Wb8OCOE2084HXn3J9J6AVbuA6X99lLO+Jbm3zGe7mkGRHDIg8CeMdq5jj6BHvhL
CqYvzfMrRp7QMxZZoVt8+p+zcfqrHd64LtotZ7xkJgtBJXvTzohzzwWQCQGgKPKQ
uyohYsVl2EKGLEWDOfk4Y73YqPA+Xm6MhlxsD57eb+6wmgM1HaYDYbyML6nqWdT/
IrRiW2dftwJXRFynh+p1GsKL93uOSvI1KSuAQfGk9ZiYp0HKaqrD4euxnm0dpwij
72TbYwKbqzQYnvH9I56XN2A5PZIzqjNVbWZjjiaKMePxVpwrmf5w0PhyrwbGCim/
cQ3iyUuKTvilPV+XNUJoqDxzGeEP8SvjYtQgsPbF7xzDGzPHdutPNQzET8RLthQY
q7oOjiYX3ipMbXvGkRgLXeaSRBPGjFC2QdMpqLmHSl+bOwAgJIv/AfY8Mda03z5/
HDkEVm8/HkRArnsiDSS6iolel/wLE8eC7D0VUXzeDOCTgAnMXjSWl+EBPcH3TJMb
rOKD3PTnaoeC0Z9ELR4xvch943lw7cxqQTW4V5yWCV5sKIZgEXejffYwqi3BH0RK
h7sA+pwJEhoNbaWwqo2EwNgDnkAoq5wiyEP52xUL3bjYrZ5vmQO+NT60c/aEZXXc
u5+dLaw34Uca/rr4KmGnofpAIc2zFtDnHguH3M3c954GlgG66VLyiDwlq4qhHPTc
riUl3z6R+EP6gkYZ0gAF4nVov/ZxrsU3O6yzw6CHB9GHoR9qoH45jG7I4S4AHN4k
gMCC5txC7qU+E2TAkQVAfMwIzfjOVIM1VzousQh9VSmCnYzYjOHE+P1Kndh/FPzo
mn7RRtl4J+bL0epA6st1/h1hGKgO+VwTCtJsc7ATwUZQdlclfoCkE855NG1Rugbp
61gcrAFz9XLjEJ6ttL9m7LIM/psJAj6+CJBHbFsXve2/PfI6UuHYWbJWdpYea+Wk
C6M9PdUydvYDc3EXbg87lLlDJsupbBe+s/a3uZBMr7HT0qRFNVyq1ZXw5idvkSUY
LNXSnEo2dzXRaY5kAcqqBqCgerZpwObCNSdUl5b7n180IsbXUN6ucWTK22gNQuDn
CSfWp2H5WMa4venmi9pki0pVrBV1xHaz4uJKKvX0+uOWvoF6pAbkFxqW3qxh8p8o
Zuf1yiyZSxxk8yWgw2vmz2TT7Kng3HffuyVRsm+uxucdp8TCOohWP9XRybxvhwHg
jS/Zsm5rnwBFpApLhPBfN0MRHMt0kEQWL72fs5cRUdoRc1MbeFViTBGh8pa1LUNS
fySergBbwqRwC9ApJgaKRPJaFKSpBSG8/PTfH1OOk7DGSK6vsE3YfgwqJt6Q1tdn
2wb+oZJuSvAB+L0lXi9684eT4hyw+aE7DYZuEn1aPbxB7tac87ilRTbRHZV4hk5E
Dz3HDhesUeuSxGeQpPBkPtAv5ONviBQo9weJakHqzGDIZGqv46m1JqycowreYTkm
kDdHZvswQnZxBatCZ2xBy6/AGckj7sUqey0N8sSowpbUkdSAp6hYD2K7SELEVu2q
8umKASPSVd3ujbb/hs6+7iwCexhPSb1JaHdnU2t/24reewS67IFRL7wYDjG2zOSS
qcE1dN6KXnHfU1X9UVtBPMAREW6GdHV2KgtjaSTaI51wtK3A00JshzdGVct399xX
gY7Ha0QrD/vCJx6lmrZCENBhOQ/2Z99EfnVQwK8aCeoNdUtdaT16BsLMdLlmY7O2
NKhAX7NmfnuE+jkpqQefy1MZzb8Tx35Sk3Rc34s+1b5vuYEkJqdLClZVTJuhNKHO
hrBPE66lr44hUBrWMQ5shx+s5Pgcy7xMN+4NOhY9VhoI9bzSeRqAq1uWhoAErx0e
EKq2IyPbGE5HzSmNGW4h8yLaSVhcCzzMqUwjan3L8RZ1+X0x1IHiWN3uAxTMIFQl
VCeaMt61snK3yzLf69nkqQPYJElD7MuMqOIY5Z0Q8pTDH7ncmB6evaBsH/7SdFA2
dsh2YgRPVhiLiH8HqIeXW4T5MAzSDdRIsEkYB9pZ59M1nMWLbjufTk1oGwMkbaz9
21U2t6HgHJfErbcQw0wLQeVT024MB5aOjtQSIeoxNMys1rhKyhT6YxU5sIP+YSmD
wpxFSPmu6uLtGxwgoIHj1EdMCjwtBdh+76cIZMFflmrNFT50KpXw6kk+JmpJZGz7
Z3wjkzvpAPx6xWWmIAtXzvCyQHH0tg+XDf1GrgbAJeXOqwCCMnBCZjzKtFInmqvT
1fGbJylVuFEEGxYmdN+q2iYoF6NEaDCAIyC8bcr8ypcCxvJWpRuOEI3TRFnc4izK
VauUfHPTeZ4JfNbDf5SoF8/yJX7am5bElX4jafmSreDwK3hK8E57Ah5Y4zJDx9VC
xAjTvvaSud+IW6pmTamHpagL4JHUGo54q18NzIwAM0dK+NuYZYqSqNQX/FCMcsQI
k0DM8Dyfzl7bWQZ7Yxip0VTuPafsdHT8chuevia3wH1BLm3DdrkEyZ7YI0ftH/es
aHTDoUa3pHjDi7ccgD/d/wt9hwI7yv+Oy72/IElbIuCy3zvmvmd4lJZ42BFl4tuj
8CZTqfFGETalCf966n86+paIj8USsgCCZei8PCBiQYiAFHwMQQTGDtFhMlWDhvoD
/YGlq73HbnI82OKmfhzACxKwQyK5JfdrH0LBhPFAm3G7mwCbS7pcvpltUbluMZoo
G4CM7HDkGJSH/wpoV+c4nECXJo0Ajo2b/8F2uoYcJpSj8cWIPJxK/2TO4datsVeZ
UH05S9vwyDraEqfgFqmrMjP2Pfj78nWlia39vREsWK4Yy9qtfaD7j9PzqS0BAxUe
88EN7+i1TOgx+LvhXjJXdhga9egxPxlVTuov6jhcrxd93kLkhOz4rwqiMaWMktbr
sev/SE138o9QVuLMPpVFF6mg7Lt3bmFYLbEjVV3qKMnxp6qiWECukiNbFcV3FyxV
FiAb9H8bVn+Y4R6h0FJc/vHqef4QHwOk/cjdijaCB4D2kB2j8DFTn7PUsu0XqbFB
+cG7VZtY0gBUJXEF+W4PgU7LCZMI09tgWblJdveLrCFzoF/WV6XC5rQAO8qIQTrv
mCW62nUS67GdjF+HjHB7UwKqq281zwsqM9Q2F/bhgbEvimGRpjuQ9PNrFMDza3Q9
EbkanE21aLPzXX77WekPyDmDZU2AQc8Qv4HDUvk1mqZLWaE1rKynDauk/X/NUayT
2rZFiO4DTDgGUiJeK0NCwRIIKs1fWCt/PqoV3QZgFKmV2JIvA2dc0WpNaLdbC4w4
wqMCu9Xo7r+9i+jrURIUTmQxl6lcCrEJlXsJmj/rLAqxvU3DKGXZya14NVIwzexf
UPxoKDsZFk/bwnxXwM34rwJnYr9NFJell7pTPJiHikpYfHx5BOXbo8vYq3q992t0
OaN8eBnIoBqvfrT44yWFe/Y6uXvRC5trEGCCcH3eSqQ17qkea4EreeOIUu0Bz+20
iyGA/ZTCDdFDO+PrPH7MynJ+EP+Nl2iHibQFH6Unl64WolLA8ckToQ2fGCe/w7OM
+qCbVkVQtmk3noymJX5sqASX26T/YuEx4fpS52kP65Go5tLqn6K9lQ3qbKIDrIX0
Wth9lCaUBoemyL/6W4WOPAapSscG/L0uyrRrXD3nARLZhii34mA9A1n0ZgreP5+W
AjzoBBnFqnifK6P5tjgihNTcyqTErzTbCioNjX+CDcjwxj7H1cbJMrH1BFcMC00C
sXi1pFp1IhkwoYoxymeFUBNVrEukxueZsBoLXwcmzinOqakkZOWrok/WyDSfuFkV
8x2UjD7Awmif91iAO21dLItH+vVp4221cxtHzAP8F12tnO7aTSN6ZS7m4j6nxmLi
OtBalGqLeO6UxmO1yaeR1wC01z9bMqqC7GNJ91d5IxQRG7NJIN2pU7KnJGXzBkXV
7IeShR7j46Y7i6Yb8iCTiB1wIzbPWSGuTlYGqdVnew4=
`protect END_PROTECTED
