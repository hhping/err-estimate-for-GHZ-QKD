`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
81k2ZEE7bexHS5iEo/7OUWk6np2p0XVo2gSBVjSlDxQglUe+wXydZ+6ENq8B272g
ppwSV/y99Ld7+2VVsdtgm3Om3TjzkPV+crgUKlbSS51cKwBg1CGYwT7EAyD/CbWQ
JGXTM4RQsFqR5isCKXQa5Yo79wSElxo/Yin/QT+DytPgYW/ACeF25/sWTp6JxY3O
VJL2kEBjEMLjkUj8JjOZcjP+TeoJAHv472T1N1q68c9bf++IOjJ/JBxB1qaCqTPo
jw0fWUY6Whg2GQX9S3h3dw9WE9eaVJBj0LCfoL1mopK6n+sBZSTFTqaj7C8kWX8k
1gHP38Oht9MHR7xJRpGzCVZrLhDrAGThpAQzg1yc/9+hrV73IeoVKwgH2QRZE7jB
bZDReXhxH5dJhToxUqihUXZi/NHZ+APlNHqVoGDH9gqedi9lGN1/59k0dXC67u/O
8WWL7+QLdmrTMT0BcRVbR6FKy5zkoHb4oxNtZcxhhwM82hJiBfhsxz0/gPaOPsrN
QF7QQvuq6CXietQ/MMNLgn40Zb6rAlt2lQSJvitqgo9nRoTRRi0LzfNAqM2yBY1R
sqaiwlIliEjFRswL8fBqirROrhgSupH0tsQoIBrFoEeft5zbnQfofxqQW0094f+C
RLUCBsTbj4qfoEXYusfeDFQKyS7DDxG0ygRnjMyJF91xWdMcpxCu9aoyHsnuTy3m
xWXsBxc8xo10oiMzHN+rZdWz87Or96V3/TWPPANWdcy++BO1V4yoM4gIuri47VBv
9bMhrCoW+pdhlLE5o+twU2lRVzwLhG5j8U8rfpp5Qc5Mbw0rysrguhZAQV+2sQrE
ehwN+SuaQXF7ZCg7xtJbpk3q8Ulc5mHsQgYpNCC3PcHQXD5xqPy/wlRWDWPI0OTN
EtHzw5PjVqWHqXN4vjVeJHe0GlR3Wm7kX1yxFkg9ZB2a0Kd1fRYa/svpD/YClsQe
48ckPS/V2mVHF5uBnVTgZ2SMjTbQLJlhQUZTUQa9A2wAtVdxDn5agq9enitCLd1n
RKEl7VcjjxHytFTNbVBXt5Ud/2dYs4nB4t+Tpp6RyEVm45gUHR4KsRgzVV2XhmUW
0PXyhv8gpMMWZmQ7cnmCn/FWmp5d1QnP599G0K7KTYwjJS6BjRF0+i2R542j57rO
jWwBV8yPE3XDm4juyarNTANlwbgX8g9j4+vd+SCowbwgsodQOSGytFok2d9KIsm4
UIZEtYXQTSMS8HNcoowORLeOpHdVzenW9UYNfKyc/Pk=
`protect END_PROTECTED
