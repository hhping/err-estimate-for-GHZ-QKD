`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EjTMHeJVlAj8LRwzNA769DTvAl8sghTa9105zeRngOTHvR2cjuw0aNMMQfJPPVVp
ef36ptceZStPRhcTY4kODKliMbVNbmbZ2/AS1MXhw/wlEwuil11fXaf27tEEZmE+
HPm6QEl3pwOdOuFaJZFhfZZwtkpGrJ8gphAsDXl+XSb+RJ6r54buL0xaU4bnW6ZM
4aRmUs5tIZukWJQMF10EF/aZN/FnGGpGR3/Fggn66sx3HmVPXhuPJJISxi1j3cye
0VcNRqaUcb+amycv3osy+uYahm1Q8+2cIUIzP0F2xIzHUF5kwV3Cc4BSwaTyaV+T
1KKYU/i6pdoTFM13eFqjuQKwCnp+qDo7z6+mWujc0C8io8pLNITDiI+XEk7d+g4d
4V+RlJyJDBvtr9kjgeAxVEDjb7kgQA//+EWWVpKToIr8s2cnRQYUV+92modiqrq7
zMjk++Ino4+er7cHu4NqI7D4Stg9olQI22TofH7Gzt5Q/OhvLoFX0R8AnhMk0EZz
Xo+glLGrdP+oFKxRegkEMZRZXr6sQ+3eq9i/gaNeD/GU5cyXQzFDKTQB2Hh+77Zp
wHVyWgrwTeYiUHCVpI4ccLntIK6qbeAt89nUbQZzqALTkxKpDVLPjipGqgIIBGvH
U2Fa3G/Q1puuK5n+LigbfdZxO/nmubni0GMDAfCXNgQFuSs7AZqOzIXQ7v9T9LpY
X7xclu8qJyGq3UWRXepTOqVOyCWNuK/olubQGvme1dSADkxuR7bvHXUNWpuaOLIY
5qDgUwOqLcXJzCsGbHqNnLJex2IjjsLFOK2ND0W+3zRRbodOFamanQputCpq2Iii
CnenjMV97+8UFUuBGL37NiHaj6GPanPRoDOheDgol6E250wsjTQgZ7VleoUGrTa5
EemBin3kj/5MXFTcRX+4jiYiXXKD7sGl2RHdm6e3GclMMjzmfOgHRfhkHQ41zLXm
aBCAk5goytbgUWNNpEmDqpVvv7iAJhTwe0uXTt0+HvgoxP+9BieaWBBqZmsMJNfl
7sfFfkBa8Q7NMW2IGFnC+l8nX0OtadlH5xvotCCiVGjK6OUquYNoS6ocvvgeVRXj
KI2qkbwd8wE9tJwTIOLp6g33XYNC3PIhaCY+jqR90W9A0wMoOHcMYxetaJHWwJBk
QSDkpUodwHHdam9TrhLV/jbWuJ6MISTLSaRCGhCHwR7wir9hkdDmswDzg3lit6iM
D8rQQvTsy+EML3gyl/UbJXkCqJrhPlfVZBDYf6EkivVAMNNyPYY3rOOT0K9Rm/zU
I/Z8ZqDBnGHJd+6+gCtiQ8Om7X0oBibqcrTGI+pFW0Tb0rNb38xBGbHfoysWgF/a
Iflr3WA/Z8C3FmHcsWzeg8FcgRPJHybCfGZXerZhe0sxMBbm/yc1hMz+LPRCbYVY
5Ey1ft7xpInlr//fN1X3wxdxIGMjNfAjgIO4JzDaad2iUCT39BZsZN28KaW43wtL
FmimOQ+oH78EhkXdZkJAO/4OWRK+TDrr6k2WKDj/9OyPg9mEZN/EzOwDl5oRXUFA
UE6kR0FYlulLPQq1cm4vt+N+GtJRb3A3cOgwpYzpxx51p7H9x3idg/0zEI+33piC
XAHpc0/X3zSsEd67kepKx29rq/GxS/I16PYJuJKMKMALzBmxVJARhHMVgURc5hEV
QTIjVERBhwn7z/wBlIzojWhu3lqyGVP7MFlohU9OawyIxcRAz4QFdebooym6sash
e/k60g8dDySaWNcYNVXdfYqw/Fj824KaFlxJLdnTzjRa02vbd59T1OuuhKZSYMLi
nh5AvwXPxlYoxweATL96rpf04lgs4CdgSHaEvuxyrDEwgxy2Jh4wPJQ4DUIAIqtl
KRZcE3o3OimAf+vuOMDgNmtyUZ94N1GKRYHtDogB6M7+oQEa89zue9todPbOUMev
OEvfFrfxCtKFD+0Ok5kYwIBHCvyi8N+9Ry4XXrp+U2V5uh0CwV2YzZKhZLhSvuzS
RTAIwCF7v193Y54cDxKbj7+dIpBLrBqpzWPxrTWUK6GevPGSPgti/Z51U7K9J6G/
eFgRbgxHr3rVSrQ4TnEMXZqcb2QS8gTk6W/3bQ9rBKcJQ7/Cb4fh8e0AkLct1Gm0
ILpbRsIkYAVPfIBPJ15W0OlGrKBStqCkQoF4W1QchdnyraEFOuw1jZ+Q5T7i8vy+
tSvXWF/piHpoJvHgAZuhPMeFCHY00/s6WfK08bHm5g6ysaPDRPIan1TTf7uyfQjK
2SgPWU6XcL6BxF2BOvwTIiFmby6K3P9yvPym3RNSd/TKF5J0b3Q3sYh0ljTcxqGo
BcJEmGtvZz12GzFF/xQvVZFfOdVuf9tmK/jHsl2LcflrWTh7C0p42m3C5saHfNne
XlC7dX1OVww2Ok366js4a+SGXCa43Y4zkM5pe/rV40kI0+io8AHF4GL8NHHyf0gI
HsM1go/ZNY1wyBgG45BuPLvE5Xt0fp64QHNwYeklHjIW4YTu4BKTehbP3MWHApoy
icne6aUZyGCnflcX7qxT18EIGcE87mWBZ+HV/1r/AO8gYvldQaiUEtCov0AHgxfn
ZNPgkPwNYxXYREN2IvEalqe+5YcfS99SWFbg/yariBFHzncyxDiomYwzUTeI67P/
5cVW0KgOIfeRHd8vkK99qsIs+a5N6vAyqQqoRhCA9yWB8WgSBmFiiC+09GpJjAx6
Ul4sKD2DtFFuDRTc7h7rgEtvBdpJEOUPNvdJinmSFBA0GPGzEgRqV34vDBnebIIE
dGj6GwUKhjZAwVAYnpx1fL9pYLtbZItz+ojnzfCacweRzGXTRPtQpdNDWFpJQ9IY
Lb2FlY+K7aZHGU3eBI3GpG/KmKwCpUavcFSFyV75Ah+G1Hj+9ADTuWcxC9F1dy0X
DfMSOmTzE8O5TZQh7zXZ5kFcUhmxf8C0CaOFZWvAdVVFz0cZ0yGFlKAthOU2oKG6
j2PIAF6lktttXWckoCmP8EH4gxLGjs7xdlLaJ/8BlnGsFZkbfB2P6VnFRomkA8Bz
IF47GicQaCrU4Etlvs748ohd/+53qFCqSOWgNR9IwO1d78G9ZdnNQ319Kz0Q5NbM
U9Se+BkunlS1kgan4OIqKJJA4zwMC2gncx10ZkfeMoVVxUTUuMZxvuq6rFRYZTE/
BAFn4j+Mg1Rf6HkRT3MOUPXsAGvMphK13rWj+G39MadK/8VEgAAaMEPpqgIImoEw
LLNTROmNvveMBSbw0FQwdvj8Qo8oipiHdWJygfUvjlBLgOBDbtlj2sJfRuY2Wa0P
ErkurNdv5aGfiyJ5vrwPHxOLSIaDDF3JcEmSjmnz6BSCUUT+BB5wbGS6ypY2PMhW
3YtFY5W2M6XnxupzIXBes0lU2ktk5tH2Bv5fhyuJwEDq7lllvh8wKzv61EMfzppj
9l+krgb7pejzClreL7FQnDaoswXaJDeYbbWud+whoGY4sGLcUx/I27GdFEe1TBq6
Hayb+RLlnGb3ysucGWzEHYGQfwUNzdbk6mrXboi5E9KyYbdZ5W275bVUtTwZ0C0F
ttLRFGlzftaz94rb08bK5BcAOLiCsnPYm0JeTbXBd/pXE8O3Bttg9Y2Zi+LN/ylx
RY6DXXMDg+DQhqxAH5Z0lVuzDCJsX5za/BBMWxEnjwv4xQX0V5OHGOosVDpir1+I
bW/wppdv1S0Iy5y2keJkd/jEAyBGRij/Qk+ceH/J6OnzkkjUDn24Odzx04vifsL0
azvTEKAWcbSNoFNpSYo2aaQVejtm7Eoa0aE0inbRbuN6je86wbBtUWJxEhNP9qFy
NA+1rQI2ODQImLcdGrQgWAG4QNo/6tnv+yn8FPsd0sdCPt4glzOBMUf0iXFwL0D7
40peMwykIkbaPd2Fr15pgMFbycukdrBAs/ut77rBpLi2o2lPiAeasdLeOZTS/EJq
JU0Op3uHU2ncHCjOMppQak7+jqHI8EM4fZXda5fyJotr4r0pXQVJ+U9LxyA5Yhn5
cFvCtpL1RdGMfOsZ4n/0AX3bF+FHhLqs+qSSA10qbwl13fu+/ohn0QjNzs+CPAMn
TH/2uWu0k1AFO4eVmOTbGNe+UYeOPr8hZsNj45/1+r2WPxe1TId8/+qmC4uh6TYc
msoa3k/+DbFBXEoScpHNdfp8Lo5LvVfQG76G/khGN7+wZzmmfTDjccTfYTipc69Z
oCAX+2Q0XPNyjrcFLHMAWJdwY2LR66mUKHAG12+db67t6ZJUaZgQOTrt9ClLxRzh
9B3wmuWxRIkim51CrSh5e3jjb1Zb4Cz0O2HWmFzMtlwa9EkgPwE2b/5NImyVZFp9
Ua1imqSICJC/L7+X35zYWBJcIHb6J4xsWBTGdXbST1W+VFwVa0A0/wo+r4NJ/i8h
/mvmjIBAy+rhT4TbIZJuMIVrloPowQ+o8eBT6m/VIiq2dHpULkdJpDm11y6/tyXP
jglv0FrkaAJ2GmFAoubFbwB2pocEg8ORgbey0iUZZWUy8dBxpKu+oECi8LDAHvbb
HiWSuFIOcbsUeUAiGYdhD8e6AwqOhJAsGB7tz0wsKS2ZEznkCdfp/p0Kw9SKseNi
48HkYDd19j0aWGtCFh7aBCAmiwpzkLNzFTjWo0E2m3QkkO6jSiw40dASca7eMGuY
DbCiGl418JJhyE/qy5ESGZ1oXsVHKNsDMSfF3UbM0sJSW5fqRMcsw8lLEJCJJ/Tj
MR6ZfMPaTACcq7GeoNoADYCx4PmVpgHEeG67bPYNpDGlqjQori9wfQDFPOB/6Cao
3s6ZmPcQkPi15rjsMd2MIy2S6u1CwJSwK/WO2XIWrRVtwr07oxnHlJXTcQdxra+X
iPn35Xaq545iC/qCjmTnlCsrPlvCrrUq0s4bFygVoU2pobYRx7EE28saukBfpfWB
hpcJbjvRBdfCSk6+hpmXvN7EF/JPKxGOhy5UnjtOB8ufnWjvUM70J0kSBTks3DXU
T094Vip8CQGEIfe5F2IM35XSQ9OksPmIr66WcqT14WJw31btdzNziwoxUVauknDF
nHEo4L/bQPPMm2a0MSanyRj9uPzD2OAcNwlO0f20qxNtKTaFaehrrXrctBmT45Ly
8PWwd3CMNpl1D5eeF/LvSiP7+BhuqdUm+vq8AbbOuoobz1tFcMl0A6vsPtJHN1hB
vFbM9ol99jJnrQW7Zoi4gFbANjU2gPBLGrXBZ82jEuuGZbH7SRZFJjJpqUqhw10t
rAfmbn7tnUvt0uLi25Dx06TA4OG1AVhk+UY0O1sobPsYaKIqji3GegxJBEffwLbF
WhkXGjXPpaP0MU1qddnlLJQBu421qdxegKMbkE6dnnMlqv8kXKy1+7ej4pBojaKi
CWL7lF+YmFOrdYT43qG4EazBnQk9HBNnIO2INXpsxVkSwMim3kZ3l+ve0AJM8oyH
6PEs/0U3QWSf01cmNtuiXEyl1nMKUbx0UAVy30zp0+pTbJwUdmSZtzKdKFaCNl1s
zulqZq/Qyr+avCquOQIqaf/fhpR3zZaKlTa5NXxXS3Lp8Hi4WmcZmrS9Z/3JyVwf
D+0lRE9+w92i0NyYJRGQCqsxqzfeNnHUQYy3eZlk+zFsOfz5ZtkLIZTxpOCJb9S7
hQN1AAVf33niZGVjna+Y8HqsW9m9qdHpsrY25GxOW8KNM7aWmQr0uyaGAopKOYif
tkEjmbTtu1Al4E58ikx03QKeV0qxH9aCyPV+t/2irC4AIf80X9I3+n8H9/qlTyF0
ZOrMbfwRol7zcqX4FrpUl4974RJpHqK86ioJuuXkO/gTJ4RLqYgnqHMbrD5GP0ZL
b1wnyqTF2PLpwDA6f1EV54yz9RebZ/mazVt5ygjAwvWWmHPxEpMrOTnonbc+0GoU
NTWAwwCYaIUXm0dBFRby20k9MTvLBV3i2BHx9rJsqMrBWRm9Ow8krlxxocHTpCPo
V7uXLwduh2pIXg9oQ5sbix7ei74FQpNKw+65G0yjRM4HeHvKfn1/2YqcGDXCR/Df
sAP5j897iXUahN35xx/3GFqbWNWUbmbCnJ+/JDxnCpMYw9JtSJxYdVglg+XjWHhL
vGTgLtUShgIajQmLEGrvAeaWMGsFLblCWNDMjA9eqgwqg5hGppuQH4BKuXyymZai
nT1+NTdgdXWypj7O0ZqQ6jnx1164edL7COjPy/2Uga+7JPA38v+nu0Cdz5qvcbYe
K1KNBIxo7Iih8zE8o0PAFH6fsH4gJBC5vPjffX01B8MB5iUMY+sS5GP7GMWuv6sq
u9Ht1HCpLUev/BdYLT9ABRd6yZfYMWnaeiMk+R0T3U+Dym0jnVAJohbSJGGkOcL6
ZGyIVUu37P2JHfAB5hBQ1lvDRjF28BU5RUY3mzrcw4eKX1WIhAV16AlgtIjIoKrK
WBLM+8h7ZrnHAZgOrFRc37Oo+dtgcU6HQswFmsguccvXXMig/9ZXIpVFZ5rNFY/W
veQbAz1a0DHZOVBq9LxjdMlvzkjpXphBKysnfF01myGIBAL74+lkHJGgHraMCs7Z
/k59JiH2boIGNYJEsaCZ4reWB4oq787YFab3XhiES3W6KcMH0nFsSnakJEihiIZf
vC2EPuR9iYUB4OvL3Bk5eIddXQPwJG4jd5XneYVfkZH2/bitl7y9RQCAgXbI5rfU
y3tBsOFfBx6S2kLDMuN9T1wII08N+2Lbu7o1zP2o1etltck+rJUsQcOu0dlKGpwe
dexQptQqdtR1Bo7KQflzBVHASECeydlM+jHlxgf+E+hnUQTndkhQTSF+lH/oKKwR
3udm8OuOXWc/YjQg7QPhUfm8D3GVKTarjKheq+DolOcy64ngxi0V5N7DG/bYslBg
xnMyjxCPvB+rI0lHfQD7DT1LNAWx5QIC3tvVI/yHDzjM5JEvO/2v+jsnMhCOkyxD
Rgmma9lLnedeLZOrSiNLM/C/rKoe8C32t2nfJWBNajQjhKcKy/eW6qK3fD27dWbW
AGLmfHqo1ij7WdeIy6lCx8ORHO/ZmZE6f0+N20asWfmtsSyD4V3w0QRbsm58is1L
D5pqcEY4+IoEw3TdM1Bo3o4cSF1dh+lCsgt+cNrrzVKTvRQCDmxGF00IzC8kOHs7
3+J9Y9ACLi7sor1t/c3i1qgUjQlSZjGDNGqvnzKdQ2/zI3Wfwcq6a09wpMUodgmZ
F3M+OBdTlyLDjjo2Pn/9QQuqoA3HMUPukC5/xJ1JwZ1pTRw7Q4xMAxGLr/Qb3Dd4
m7JSHeJbQAfG1e9csT5e7djBm0izP2gGIG+snYbjDCId33kswWdjcPh8NL1ZhLkO
mX39hDP/UFgxp6abTPgOSE3LCMUYfhxNIg/8buonRZCwTJfPOccr413Ya8VBHAOg
RejIJl5uy1Rv8ujFtgYmQc9dtZK3VyBHY2RZzZh37rfXX7RWjtROopxk6UWbez3p
MEmwZDZoLpTeXz81zaXkPldQrZ2LM28Y89j7JfmZlK5VF2p+Stkb6kZbFabbSVRo
UaNv3EOn40oEnS15IxXv9/N6ZwhulZPDlVkWT0JuP5ke/0UDKkQcZbl6xusBFPpE
0C8xmqK2jBMftKnYtOI2oJ39nSqZ3csI99zZYTnnDg5YWa+W6Xn6R26bn2s0liIm
BJu8BbsPvdUoT7t/Xj4BBQZWNYM7lF3Xlo9H7nzLFUCCKAffpJSRxMWw8HwvsSAX
gjmFinXtEoZzgyCUTEOhYRc3LpGc4A35bqTm5kDpijLDD+rbRULjTauFiBnFi2GG
DCkNAJ8yXsqZwP3wngWp2lDlt3Ii7EcMKs5xotsqNObeqx1WAQ9lgkk6uNAu4P3A
hBKnas0eu1SkLyKyF+bVoGoRUqso0q+R1ge1hz8P2FTC9AqSrSxoprN7BRMEw8lU
Om+nObDq25hj0pFOSYjidPeUvjuuec9ISpcgT10cL5kYdx3n1OQWD49M4/tCj8Ne
f394PwKAybSQY3P3E8muiPvsWNTDoI/kWjN/4gJbb8Qu1x7iZlnGYbLPAC+bftQj
rqFZy4JtKvVpypYlnkE0rLsVcLwbKSRWvIdNZM2iBp8wlATPk/NlghsSOanaPhaV
JRjMMfC8BuZnVrWfgjUQ4+n8uv7O8dW71+pV0z0ugf7MaaXJwNRHngjtDc9x8ZZc
YRW8QKB0Nhu2Fx96gTvzDhjS/yT7IrPQAFzS8Psj8uvfXlzfR7eylwbr2ENc4h+I
tsA9dEN1ufuLVw80elTh5+rSgGrscp+6VdEp+RI3E3N1w6mmOUBuNq+smKAE8Qsa
NZAPDZIUuVSzbTnSZaxqMb4Dk95LVVJ95AC93tK7uZkOcoUukyc8xX+2u3Gnr7yt
1GQsxL54ky61kC9557aXjEUHfNF+H9a/dWCxwvsDDTWC5tde3OgAl8F5CK19N6Sn
QxtO6IO8LvW4fG0fiTuMAzQv6SU9B5VbGdpA0Dp4gnx6myaqjuzXcjeouo6aACHr
aXVJtRpHxjCcvNigDEOmgSOmOaNQawe+7wT4G7/8yPztVLdIQ9/++pVJZIPizMXl
i5MzASjUDQTOJ9s6jXAlVw41oPa0lcLjoCB5dXBO01xk1BEQPdGzUUU3NrwqmazL
B1i9asJsNtToEn5ufCwtQ/sQqdSH/YPz5YUz37ZBEXqFA7GvPCeby/whedsMv4q2
LTbWRxlRav+P1N9jSQiZyONm1tllJ6EYCpDmwSUxRM2ysOUODkcXE06ScFA5dY+V
aL9zxd78BtMU5jn1w33JOxBlGhi3fQk39qjkMMBSL0O93wW2xEshX5qtDVofldkC
Dk31EyAbHYWjXnfDzUOTSD6qIiUQLCSA69VIkP9Z12urnhymXqSxqJXop6h0E/kM
kaZ6/k8ka5DPLHAZWGJyBw==
`protect END_PROTECTED
