`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sz2nrMn5jPrDZfpVy9DIIQ3Tql0S2BIpm2iRP+MCf2njQQFtjCe90iNg1PSw65+r
KdM2vm6a8okIHGYyHKDbkk+IkDB5pqjW4Yky1WgxeEc0ogGoMvSZeZyUZhhrDG8+
XzWlFjpWUGuTInUjS7mGe36bDLaseojhRI5Pv9S03Xc+fFq/k+4JyIb1yTveQH7a
vKaF/jJYnmBPWs0oMObwUMFfvPUBTFAFxC79gdMZaz2ItZZK+4nZ2UV9IJjEB4hS
1lmLck/CCoGdPA0hTZ5O3Yt9k64SZWPo1tANoF4N3LnNe25f7Di1aA5G04NWqVx8
Tfl24azFCVJQlLGpzgdB+wWpaZ8STcH3KNXvSL1KekQMkxXkmh//So6vGQwIXpjJ
vahJAXORJTN0CbPPkKGMcyWpeUhKLFttk1BT2/JIxGM9PtiwuIwkrm3lO7ubZh/S
bmV3Rx0YzHLr57Fna0/uz8Q0hZEzlmCP7W4juGrsLxnqSw+7mzA+RYPHsCikeVwT
ISxG1qEw+OYq3oqgWkr3w/HaEN5XM8KHRiyCYjAImmh0tRmNq/4s57V67PSA29vo
IzLsL/i4ORXsRyazeD7ykoGcyw490idsUrUQJSdnHvs/W3/MBESwNAZb+c3S1uk+
rkLjRbaGsn4BzIPFT9xQD0hm46cuF5Tw8JvvtoCODY4P5qFBLPX8NWYQ5XdXumHO
+Z7Cx/FgCwhgg8IWPkNSEkgar3RGOYOBLV5jzZ3Bj365T0abOJmlfuNAtB2G8Y3C
`protect END_PROTECTED
