`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f9YsVDdlwNg79v1OE0A34WEE2cJLo7lq44hBLtBzzP2MAZNS+kcyKNejjnF2S9+p
Av3GFQg4JFtvFIUbjJMXMG4tdnYyFAdDMSR76j2SWBLSBR+Tz8p7G9O2PAsTZJsF
wJzT8oB+Pmcod72Ei2XDEChMFi4ev7sAzQNRmd4u6ldckriIevOI7IMwO0e9N0oA
9uy9+OCpLk8WtalcQuNYCe1TLNKI75/i3BGbmuxvegvq+IzLK7t6mvH/Px215/Ga
oGHC2p9eKcGJHW4KPnrGrXlmn5i3IvvrSA1uCGH9Y9PcKitlb9y6cQWrZiJ5YcIb
TUEAWWcnICQmEulVmJ0b2C8XQOwJUZdPaoKry/FXJdORP1C0fx1MWBdxGib7TLW/
y7LhO+fxbaicY9x8m7jxi5IPl/1LhWQKwinBWB0X5VL1npwyK01fD7TVl/xE2iHS
EvJEVmiEWfJvXMgmMEF0U2LRMs5u7S4bF+AKPsV7yEEvyCwVTChSqe6nu6fqQ2eQ
AXanvseSS4tmB5n7QYRK4afJScnp+/0NCWf7qfR2LDA1kbTbkXwx43hi0Qg69MRo
xhJb3tmTeX6alfgNgT/QhoPKA45GW4wnhP/IdhCZvtrX97hz1ZiPimNpn9WXIcUv
dfvyHMJGyFCsmcHLuZ6g/A==
`protect END_PROTECTED
