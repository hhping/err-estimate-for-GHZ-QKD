`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s+0W5i2p7wPUK3M7Z9+N2hb/7nx5L41anZetdzIsRDVO6xsYuhkXiLnkhPCBBser
oW9tmpy6S4J425QTrHrkvQpTPUulPguYLyje2qPZ7FNzKpR/iDkyEH3iUJLKGKGr
y1DRF3NpeVPQKmI/WVvb4npZRZq0iEmx91WWGVkLwB1kdzr5w4JlfaSH9VyQz2e8
0DwhwTERUlEjMJs65Z4YYBzkHpjsxdEQyHKYFrlGBJHwzuznNK7E83qyMnh90eu8
2i7vGT4a5q9dINCA0oRVgeCJ/nWtlVijAIN13WMF0/zjOlk2w3BHfX7nr8+RAT3s
J5ElI3KJXxrtDHR6bcCq09E4Jd1zrzP3KlkSlzeTOs+GPkaZqy91pAYZ6gHGfEhW
h2Q1zwSLLrxOatKextO2+LyVcIp/08TepB4KHV89rnS9ceCUhKt8+jCXHm1fzhl+
4aNFkDSfRrUXmaADq+Z7Lw==
`protect END_PROTECTED
