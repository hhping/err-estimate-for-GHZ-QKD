`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pmgv6rJZYvcIAuPRjC+0cFhtVlcf7APZzSlxtlJsNfIEn7cFFW/VHljYA8bRNdC8
+MjiNPP2Lp5dQf5zhmfx4xbOjmDixvnQJGitCKGY5FS9Zq1rb0DRgqPmEfvk0dmj
uB15g/B3XuDLEN6P4wsj68MhXfmw3/2iWwkE7L6QYC7ZwkZ7FuZ+m2qfbsyVcwI4
usFEm4Zmnf8k1thj4IthWwUXK35C3Q+C3F36elqleVysQ6VstnL2oZd2JLZEa3qQ
vuVeTGAS4G1rAmXkOYyMJYkm61LgkN4kJHUEkIW1Ly7SSkgHLE9H0ZAikQBAc933
pOZpcPQsszqzSIP/8OsIhkcg78Dze1xbmj23XClBDKbihlv/qULdRZu4fxVo+1u+
5qRgONt9eia7ZbFGzE++i4GNizEsSq6ruteEZ7+/Jxa7YiFjBj0pMoHrv2bLs47c
azEu8RFboTo16dCoqZBg3bHvE0BWiH3Rpvgul0/Jm5RjVW2NlX3DigzdGRqi4htC
tnUFBGQwDeJLO3StkbhOumAo90GHhsla7RkdXc4ETArL5jzy3sS7yvuFtu6YJviq
NhdfPaoklQOdEb8IMtkSJzlINuGPb2j9lhdIZ1ZeZtNMWeMNFQIhVUJktExnUwIw
7PeDvcDpvqmAH+RduS93fjemTJWKFp0t2mbrYIfk0Wu9nNH3l/+C1Ka0lWi4phKP
uWXZf4aH3JcMyPW/2Hf+7eT282Da/7dx4jTajmkCEQIh7Qt1Eu0JOWKpBQo1401b
k96zcWd7KNhd1x2GumF/mUNbYFafabVxrXEgwFTW2VX27BAXGP13rfR8uEFjWIb3
6hyAJDl/XhCAG9so/UgEesOf6vT0T6+jBdD0PG5nPr2pyTsU0w+B+inazlRQ4KtC
jEAjTN+LUn8Lymz8enHUHAb2EoaeaRn10aMdKURrOwEp/V5de2J7Ffyml+hK0DnC
NlEj2mlqSq6LV8/e20dfl/c32CDfrSSXIRboD43ZMjn8fD/n2DpFnnalZUGAiGfE
g3VvjG8vcWl+v7tXm7Ph7RTOKsnp8Uz6pLh+itP1mVQRnyk2r8I/1g4vvrJfBGiU
8b8p1uzPOrWzYDTqvC3TNYbi2BeT72B+grAMbOQxdmwLxVBacZiluApX7+tddoP5
VGE6epHZwG5Xta9rwsuypyu82L2uGxSBEvE6AbdJ5iYL2QM9DP4eHEYyCa/rbMBL
ZTVSgmK+3NafyAzm3OJs849+5nYs0me/vJHMHaSkK56G7B93muSS4l1DE2DeF4oG
mzzArO+XUtk0z9T0OBIL9GZv1uEv7OX3pdU7TaiqVkj+rGezZEDi1MDup8cepOMI
EhART2h6/EO8UP+kesbu4i83tmJVyrMbZKwr3TrWuTUT/PfdQjjffCC5KgU2esOX
U3mKTMzRRD3900eX0WUgHOUzw39Au+XixhUSTCuIPnQ1PKnGmf6PQZ50VPDiqoJ4
qjb+2gL6RN+tmHX9S2wlRTp7EO40itncTjW2UBqUjRJ6UGw6LI0fIwhSVkuJKUas
ZfQE6jz8+olaTfzHMKdwPyF+w973hJJavH36hs8fMGYdGEJ22FrTwOapPfCBDzbA
0XQwUqYOpkm8kB4T63XfmRcF5jARtEV7BxE1DavpRpWITk2dknzib3wmjM7Ic1k0
nX0doWr7BVjf7aEnasdclBQhA9k7SwrZueLFfPOxsRtR3nt7FuTIn2JgL17CdxvQ
qPs/0ftDqLZlTwv2AQzGNH4kkc1nMBaw9Sr6zW17O6EJLuiuh8Q3D+lRxxYSEXt7
/mJXRAE6qCqk0t1KMeVAZttskzHsvQVJ2jO1B+luoU+sSy+loTDFv32h0KPJLRzT
t6T9yAOsCw7lDG2YVCrvzRUtnzDGpjT5r1QfKewZG5M9I1fZvaoI7rSVOLVZASLT
D2bKdBA/lfz3LPcBPdjIXyg4LlBz9UpxnJqO8NHpw9cdxwS8ANFtN7U9vI9MSZGG
x/rRSZM3RYDyqqrtYbQgPFW4+GluvMbngPxwsiWGY9XssmykWaKPQcG3a8PFFsdJ
khbFBkDFLgUWYWL6XQhieQH7YwPzMfY4Ts7yEdsrQdjJsb88X0cEPRtgLL15B6dR
CKmitp5JHaH3YcBzzs4R+egkEah3q4ud1BISFYuPRSputQkxw9RX3WooLA4u8HSe
PJYYN2w9cqQn/zhQB0tFD3JKiJyJK1TG0MgSM5fJu+wnpAnj2ZgUlww3ShF778PL
p9UMxIiAAFO/VdQyQ6GAB3YRR39FF3mY9Qk4cV/vcdqDLKPV+JxJk50I/KtGAhF/
9TfFw8HJnBB3UV+6TTpEnCuFHynlrKN9HOxJejBr05wzIw23JFOLeNNXRQX6VWEC
jba6EvbNMaz+ZeqS8MD03Le6/rkd+ESkRIOc4J1YM0z/+h6UHYdKEJnt+kpqhPaG
WC7v5OywU6OUS1aUAjkmDFyoDlwwpVDOXf0NMb9/ZP7LavtFHsd85g7WRL/kFX/J
NEj9fPtcY3hmLQmtSWrBiPN3Dq1rhC8Jrgmskxlu6tKAbDv5aKnJuGyaaJv5I1vf
Dw1h5+CBgUUGeKw67RGJpRU3c4V5r9m3dijZvVjN/yNbC511tHkUpFqQJZiSSEkR
p5lRY2tXYZi63zYKQafR3HdZc6R9BoROkaxCCGoG+kuF+l6jTxboZqBm9CTgWd6T
xPTf5XHE2RGJsquaiteMQW4tN2Wimt+iL9TpZg8yUnw+he3bPPePzRYbVYoepHoM
OmcoDvi/2bMjPzFHDz4G7vYZpszWObVu1v/V4lTCWDToftClVseylOoWP15rI+9j
U+bM3iKJQHnVhcN2j2RK/2KOqDujMVlBuVdsYvIzpziWMchhRCxUwvcqrFytEmyr
Vb8tn0TPLof+mN7JyoAge5piIlzgW/BSPqd5Jr8T95zs3bNIAXQ4H96VjYY+F0KK
M3vCND7DUqMIW1Ii29W2JTkGAFGsqag5Xz/27+LcGIgzaMfh29RGwwVj+1irhPAM
bApBe9HW6pyBSyqkgcTi7Apk/GvBj7tAsXK8yP7Vvb2yJsLR24A5zzuMaKoGuTmi
4Vk9aO0sBUso64eCsLxWyZc1qogT+1y7rADGt4i5u+GoNAsln7bUeEd3Kmhqqde0
dX0diztpkdwHdH8b8oow1bsR5oDtdERnvothhWn917H/LWI6GVMEouV3B9WuSenS
lnf29j50WyiTXUc/ZKCEEaFeojKCbdIP4mA120E+Wm0wgRB54mxnq5nwRYTpfWik
iujrx1O44xG/5gwcHkC56lAwsmEeivPLjEBH4u3P6rnO4aEgYFUgAW+DvYhnef3y
REErNdXIvlnzs/ZA/o7qErqqISbM6rGVGUMxwT0bvl4eZ5p6SjGp25xlAh5FXAfx
RbqXZmPsRhGwf6keH9/o4EiN4EVtt40uvyC8ohZMuLtbhHZVioq9tGWkNFeB1P0p
dRrTt87m9KRWOfOtfJnpo9mmVg3OrPkIPl4FAzhnuV4w5R7HpDCnZot8z3HFfMnr
JBoCTyVU2vlXuF5i62yrrRaRfRXSil4zD5kPAQpv7bShmcvzB8fcAwCQ65v7o4Go
NgCZCCdJC6bwh1U+l4tIBr/Cj5PW57KNuo6y1uy1YW3/W49M5rLp30s1RiTAs5Tk
ygKt9V4yX/EyT7oVRi5zia5Wbm2k+WWsIPrMwzlswIDvIz1imwTJMIWgUg0mwCG7
1ZMXvJdJ5coxoVnPvol1REwVXV/RKzYzqcoey9iOq6vqafPlv4qvnnc5S2uDK0Ao
y52nAS6iJ9zyikQPLwVr2jQYt/AtSALVLI92KOR2hg19jm2p8vdNL1Awyme2WLBq
2YjopEqBdt9bwM3TRRJGWOy4yEkcXuYiwIyVBRCO6JELH4ofpZ1NlNS2UI7mmRFA
086bfz3dvpmgDbUCsDWBeAw0854u7WxO2IhPyc6DoagZX5CwWhwtXAmY69ZwXrFe
mGbh8d+pOc3OZ+ngc11ZBBgUnG7gkXGqDJPUDkIt7F1agmG8fOe5AY9QWx0Qe2EI
hyOFkjbjOl8Mv20GkBrX/TlA/ElTwSrSSLUgWUyd2Xe78kNyk/wwezsGx3GUx8cb
oenqqykA0elhpPi8MXamxqcfbNgl4ZFkMC7BhDJ8HJ9Wjs6Qu3nh25YgeT5KF6oH
id4Td45dnfGW3Nvd06A7r0ViV+UMFpp7RcCkcnmuDKM4B66gyyqyNrB5b3hfpG9u
82bRewoZeSmWgGOtmG2mR/wxm/6gT3Rdiu9hat1e4L38nIGUIZNQKNc8w9AibOv7
zw9/DWI3M6T/gTS13P5UzzIr3F6eCAKXcyOPSwkW7NWDcTliOz2gMOLlElE0NDDZ
0p8FGJwz4h9IJDD63ugeDHUvZla1BZ82nvKJ9Gmq0qFt3zSksvd2Kvkvaf7DbKvT
TA3wQNRpDftBko1NcyS7R8vG9ssHd6xlckHvETYi/V8YQEOOtUlaXkPjpCIL0e7/
Dctbg6wDa9zajWj0RWVk/t5MDRBYCgfAFNdcmxe/Bzr5pJa2dMQiI2ia0q8Kst7E
Gieka5ndu0H+ZGEn0OvRO1NNBzFPKsh/rhP8r39/84LwqD/KjKBpQQpYvIEL+d49
XrpPMgRRf/D2QLVVyT0ZZbKFcmAjOU/y9wh++2nj/S6jWUjWmdbVm6LzuR2M+5bW
gX+LfZ3CvJAyOYy+ljk69ivOilcS6degIwSW4sy4XSaB8AUCPJWKk1lYSZQRwiTI
xbHt/wp7bmddohn76N/WArXLaaBq2cH4Bn8JZocPErOwklW9FHUy5runUI5gTe9t
50p/ZwKYPgMiIWfQ3nSzuyAKM2c71MzGAIhdVmKpR1qSWHHantHE+aqO2ijF4Xg1
Y+h+UTHkik7IPr2ljg7MpcfvVolchu8RTg2kTcGuVhjyn5NRGXuCzc8F/yvxNJK1
N2S3+e+ogSqMaisBx7ZF6E4hUuXG56nmhzC8CqPSvFWQMLI74QmnG4f8s1YWyQg1
WY8C6l7NcCCNAL8jUv4Fvi3nKLAcnJ/icxk/koNX1oXphcrR3X3OoMwbs1wockyN
Zx6MxD9bxr+Th43gPMI5fJONhiGHhD/TJgQIDswcPk1FznAh2qAsDaEJOsXPMVtH
9iup/x56eP6sWU1udXzIHHwcmSsT9YAEPOVTVKPYC+vYPTPdbLr8YATuJUUEwhCk
IIkKtyGsv8/TNJHmQjfq3Kjc9RabpOZVWPLB3vsbnrv+sRizWrNNnOoyYggu229Q
CmoN4emwF2QmvOCSxl0uEMe+gzM04LEIWNBnetItM3Vsk7qZgbHFBt9a1T7HYRiy
I9HkWGXLBh/Sei4OFTSW/7bb5cljTnleqngXewMH4K/B3+qmVU2EMecF88rX3Bvq
nG/1DXh/vYHB4xxgw79dP7TLSgHy28QmNqgjFqdQ61WWERYQFMspxbQ4taGiYYj1
D8JFxSuT8frYtLTvLHaxZNv8vbPJRwpmNRCv0vLIyVIf1ciM3md1NZtFkVIleIRC
kqbbd/Pn6ilJXWeNBvHskBhc/9Y8Meih5FXk4WrKRejdwmdCQVBdSrGx1pOZptwf
Q/C++T/q7+YFdBWXEtzOSm8POrfAvCLyp9nabPOv2uqXuRht1A1OUmp1Ni+nQ770
a7shA45dSrvzQuF7eHJGcOIiDh9hQ2SsX8+ix+TxoDVkcV27mjt5cG762xvoF2V1
PnVDx67G23fjDAUANC6tPVcvhb+JPPBSDYm4+nhyp6x70MkldySZaOKnr1nyxAAH
u8nawtJAYHRktqmAZbtgUjo8/dj5OXNU2TPW7qIG5Gr3e+Ro4P4+LMn12Na7F1d/
qLEVNijcIuTcCT4JsFuncjnTSIf5b3s6WzsNdyzNgJpXnR9fvAGMsfWzOvADSLL0
P6cFa2Adhk/tDZVI2BF+wN5EN/7gQBVrcGiDF/RwZv7zVlPFg55/rkgwQE7v+QFB
tQyM5t6wxnlSDJPMSllNz9YrFAFDDhSMJN1rXAlI4iQgqa54qo6K+5nYLSE7HKJ2
E3IK1FxJ0/Aj8YM2bhupFQoG/AStnzTYbuMYR0MNiR3TGFc+bMwf0pbTF6wT6TYk
N/vgHQeM52vYInC4ZLEm3st8i1hYl4wg0cCrfQIe/IVJG9Fx3ItRNqHv9+Fkc4ul
bzRj1E1DyrDU2+yWIepj8A2FRmVymneDe/OcfqebGMOBv4XmOrb9MNRjswNAQ0Nj
F+jFGcEj74+WvaJiawDFnU2x2NRrgrGYfZPMReuPquWkcpempfTVG6h0EN+YNABx
1CngpyToFDI36na48TINUzEgGezXdO41oLsNmuoqullDQV1Ipi6zJc/k+dbQVQJ/
/bbuWtJrI3bVRGEuhNlAmUpSq76hvH5mzOzc/0zOB2OET8r9nZZtzNLJq57OZnLT
RQBWQyF6JwHOMKB8VMrXK7P+43xKKeb1gGwFUVaLbwPxjJntf0/vegMGtKqi1VhZ
RNTrCu+i6liexnPImN32zSU3WJ12uQHJWDXEriVtSXZxhER0OCZoM7EYFaicsHKO
YexDmo/CWtM+zXKP3i+qRH7rUFK2pTS307ElrfWNx69huqzk36XtD84jrH2Zlo8b
bIqKaAc/YNWT8ClmdStc4g2vK5J1UyCMroAE+Fhd4Jq2s3HFcFPGBX+kc+F+MYSG
kfGjZm5GEbQ+9OOuCysoav6Ydxy64Kbe0bwpxHpKWBR6BmIk8Xv9MnD952KjE8nW
lqXvtOQvcfLWx36av8rqm2t4vcdXCwxTtcFLbuX34c8K4bTQ0PjKyIiSCJsgfOq1
d+OzvV1H2QhkHH4wZUw2+6TNOB6NZgiCjzePWoZ3MMRBQBK63m7vztCV1X6qDZy7
B9/9YhZ3sjvYLgeNea7tzoNDW4dzJjsfXrDOjTKwAZBjoIkyXKmr5zPxQp+NHbMV
1KFicPOhqySQmW9X0V2ACUN3ylPJKkekgAYzOkZQUsj1SkCc8QbjaJja2WzGbwZI
yw4Tqi9Pr5kjIjDQRj7J1BMdb4B2YRC7dRbFGRrM/nU5XcpCvECVoYp/lLtV8cZm
V+KeM6VmNQ5gO6Q4NPfPIXhRQbljO2JuNzvSQbD1CH1tcNev3de6q/MrvO53ilvq
PWUYQ35tOA0wYu9Dod80NqMM03GqxBnTeRJyvGyK+z1KqWWUP4CTlg6i9MGgm78S
K4+tx8+7aRuB5E8cEUOcZlTSeuZfmFf3Ad2Pbcg52kEz/HAfklyyPH2sgzNXuCzs
bDmC2EtFo/0zlHMtVyNcFpDjw/VRHvm6qKwVSIXCSWOnyUoyr3JeCJnQltEGt4FM
SFcRL2NvdidCUX4AAQv9L8Aeyu+cx5o9ezmPpnOu4945dtzinER64hdiKj8jXtGP
Gi9zdGlEW3VS0fnbV+OTGUHXaKeZzUtvsP0gAhO1rQReKq2SBG2mphUOGXt9D2kH
kr/wm8gkAAvIq47yD5S1eE8PVizg9HDboe5n4Gs/zU+KDreNUS5tRIhSj5xwj6+1
iO8zMQ4+VdJbciPYIva6efxblHr4lCMfGqbfgCl5BcvhBAx4s/us1zpPf5A6k7a0
KB55G3oZCyl7C0b5ymkdoriFl9ZkiWofK4qaCyCkoyWW/0iWZvH1OCYxuyYn0247
028GfGJ8P7K/vVVFIMbVYReQ2DI8/Xwj2L/PVDktKkelx+n+5OiT9DCMFBxNYw2d
MwdytJhGvNSfE3YMwcWxDppv6EnWiLWxkOMWyC7y7uDefo79rQDwcWcXjq93K0P/
SyB548IL87xc/dn6XDmx2thG9sW8TZIqHguPn5/VI+Qqwyg7x2E4WNSh42q3750I
hVgHrSXbkgAIg55pRC2ChkKOJKerVUV1qH3CxSNW2EbzjvpFbeX0Uj5TkSCcjAFX
ZMPWpM+2VC24lSF28h+EIbH6SUDDCeFGQW0dfzD/tVmHRxvdp6z3gbqMXVCYHbmw
dFbutW517Kd+c/Gnp+xNyiI/ZLi5WBr/8N64vq8aMiN9H7w38VfcMsydAH+1vaSa
ioC3qw+ugkaoOLLUm2Z24mSafOCGMLt8+YzNxNWqTU4/HWfDnBubGuRMBW2gtUFw
XHW8Of+DiqPbQPPFVDfyIAFZqJOhM2uB7WQw4feKWh7mAstTmHdixNi9/179HUJQ
eLRKz/NoPreVeVeGxNrVWq63W37QOJYesiRTty7EWpn/yEhWkck5HGjvwuhq/SYW
/+2XkMe7RC84ZcX7J9vbZDY+JE9k5o/KhCI8gh4h+gKXbzO2fpndhMqdIU9zO5kY
n39kiWNPrExByonnxMa7lh5UPqY+gyTYfKgs6hUq+eOfSS/scAK58Kh50DT/d9ad
M45weVm2/CCDTTFVgiIrbs4fiUEwIG9oy/O0LTeZv54YW83MyNYGimkxmjRQ/O3p
zmm8Fluu/Qs1qkq2KwgDFPC0vQhvfcZM2oKxmUpzdBp/29Ucd94Rq/45CKY3s2OR
YxhtC9ZEfp7lk+s3llSJBr5JJct3hP92769Ka/55P9nRyFiTGDeQ6ana2pQBI5+d
1Qz/VR2h28zaBtCp4Dy67WP1oZy1tIDFhTl/AtBEbntBTZG8le0Y9fcKfy+YWYjY
jd/JAIH9tggtERsjBcwLWdEowqBokh0RwRYjZEbe82Nql1zorwi7TADmpswPGeSn
k4+exXEl7BZs4f3AKKOU15rD5/9bahJN4o7jGO3RYhde6zH45eesZPgSdV76RwMy
R/fTEp2FT4mRrWp1/vRTSY1OrGhrsuynaBwnxnToUHgcWyLs9vsmiH4h0qEnLbHL
IL8Vir4xxJp7inXjmhGo4oQb4Qb+GEHFY+nWCtQAsgLMImqcKVeDwi9XpjbV/uZD
8tc/Z7H+ITdwyKYjqsE78rS7M7y2qOIOomUfBsAk3KvOA6wVMJpwT8+zGm1AGw7+
mTsS4IOOx3PHsqw9CHGCa55JqwKL5KVT+IoFLTfDxacg3Axjp+yGk7zpyXxnCchl
AbiQ5JcxETErYMFZY0th0pooPIvJIYkyLhrEcmhi3x6oW+brSmLfuSf8/xb5IBM/
QbQBOd/Vi29qxAxQB7D3kSy/tvHoUN7vErYYuWX0sj9tGoWWGBlWqXQjH7jRDX4B
wr3m2uHP4yU2kJ7PIe/Xv+BEUomAl6cJxmmLhvyPY4mNz9rOibiIz1iVjtnQJVce
DuLkm2DFjozw2zAPYMdqa9Mz25CNkGEQUtfOyT6Q7sOUVFAAO175iieRNKpCGS5b
fNIDYbB7vmwcf1aQVu5Pb4rCHYD715I6aWId+BSxcsU22VNhoOyLVvxFGGbBOVJ9
u0hAETMDIkLRNLpdf2grMIwNo0zrTsb9WX4mU3G3OLtB70//LArh7hor4vcHi4S0
kGLVxniRHzxim7uys0M4WvCPxoJgmzgDj745JJSX1JJNeYql/bUZWnaMctaUUay4
3ltzvzZovn1wuqE9XUWC7ixJ1hNlGpt+9bZs5u6PWOnEotQ+/zGlMCBinIhAk+Lj
lyiP/lTEvKrOhDtCtiVrDGxgoR5ShtAZ8ZImOV7pQybO4RLeFAfNZZca5wcQn5ds
zxKpGSBkjiC4PkmWdUx1Iurmm6bQRjTg3pSjT0WVEpitbbjlKriJZ0CjZTTQecHY
AmuoKYvYzs9KyTluHp50F0p+9P/GQtX8xFZFyhdjqV7Ny0E92sM1YwPibENTnS/v
LYPBKrVLUh9AbTHM1QXi6F7pqsgunmhaz9/dyVse/sUZ8H2X8Oi0o0gdlkrS27s/
htR69khXd/B1iZa4UP+UqVFB9bJdR4mSykpCA5di/p8vsiR44yfFICf1Xq/kczdY
Iy0c/QU2HrYfF12BeiYGtoTxvC0iONhuO3zsv2HSEc8Ibw0LACVM+2ki0BqrW/po
j5o0wcgeJ0awfibEHxO02zfe6kw95K2qJNBWtvN8jXAAJmGIFWlxDDegdabxqcQM
vcz6JtAiHdKQ1bdcllyNb6DPEZTMGCj9Hae6dKEiMLXBdbH0jIVr7Sa6tu0YVJ+/
4dgDrN2zaafT7BGSH5PDwr/l0Uws40vpQ1pIOO5V0IPmSXrpdi6julJF/LKUPZTJ
jqyF4pet751tBBc9hPGak4ejZEqWGLYH2/sI5s3aoeHnxPrPONKxylrcG3Yn4BvD
pL9L6u0MQevT2h+fpNFoh4qV9WQBS09SqGWj7FdRrs0ZRXVGmZqlObEkycDZtLzY
emF+meUYmThNQrPJMYEvqSx/n3dFDFLx8g9p4XLWRYueo3X0JBeGqTfhE3MsyraZ
He55nYL/vc46n9p+GHnwMlhJp80LwfKm4cpcCN8Aa8tzWP369bqUhLii/Z3AGjm4
iiSM5HEH+WQaqzojInRNrH/gDd0zdBKFuMb2hZH8+zKadZbE5Ec4eGCJWHycrDN/
LtmMo/yLgph/Y0puGgehxyx3xic2+2cU7WXv09K1LSnvr4M74B2S2F42eBOMreaH
6RJKgvPSBDWUBUIlgfi0MkvgJ3wAwVeL+2baDXIiL/iYjER50aEs0EVet5KuisE2
TZSv24Mu7ncafM10BCBOIac0VHKxXzc6pKd3ArB/uKSCOjy/H5ynqzdagDMVCS1Q
IF8GS4f0GFMYsa1wkhj3TgcTJ9XwfAVOnVQFHkqrqzIQvV7M/veMYiYmNxNTpxBn
0rx/cNMNJ8vrV1jCzQ0I+hkalHRiHOJQgu8vPqxl4ZCd+Z7BwfLpyS2d10EwURXE
GU3nHobX2T8OdcQlXsoi4kAwnEtMdMFWz0ptmexTBOf2h0rXkHbID29xvq1et+Jm
S3sKoe9kEIU4EELQ3jqBPhG3JHzJZCiIdk+QpY5bFQuoItw8XJn0YzxtsCJ/rcht
SEUKRNoRQiKddhi79/mws5dIxTbW/HQyESxofJmhjYwVe7lFdymodU+wCi0bRuYA
1YoSEByO9LAM21rOAYj69S23i534glKR2tinTtRGcywA0idBWG5AMKo6v5yWI6g7
h/4Y6nHGBbtUMuknQQ64GHXAcRHMC//DaevDjHVR/MDjuwKJ4y+KnT6weRwIsH84
vW3EkByb6blThAOxtq3pYzdMBQB6btwWaKy8SEM9UpYmYsG8J1Uvs7bQepVAnyzn
kipIgk5teuE2spc8XApMiQpa/rcF0cpg1TanuhhhH+gCaZGxQpIbm79PIf2CSnqx
HuN6wlHsE++Zd86AtxNzeV/C15gHGn0YoK8fcP5j3Z7jzFcxJBA+AKFZVu5FUREM
glUjFYT8XdmhYEwKddQWXcz6XaBsuzdslxmw2jNwVzuLwgjCeG5g1H6X7WOJFlL5
kKXhw9eSwLmx2yu6MKs9DMtA+VwjJXz84UIBChYj50Fei65UyaF5dD/vLY8Uny6W
P/tjx28pbPFQItuiwMjV6+3F6cyycErwfq9EVUGGh8IHhFUsOvxoFeVNzKPN2A9D
RgntC2uNPyYKnStH4jJWI0YA6s0oo5z9nFcFbfF6gco/xsg7tiOaXQLz6AHamwpF
/FaI2chzk6fSw22y67iF4sGcj64fo/y9qVYw/iT6dVvQpjUvQWtg33/D55IjhsmA
+PmmvaIMLv7ROhbBsNQftZ4sfOyh0Pb1+R/CYa/ijhz1SiWk6G9tkSYizHqzmVrQ
oB5fT5Xk5hX3GutMozmSVPtL1iTZ116iQ8e6+ly3gZ87dNuuTLzGc3HLvmlMCBW2
eKwzCpWs2Y8ooZZj8fGRR4nww5rix7JsMgOIRJAcp+qRAZc/4bgDPzj5IruVHsTD
EuldQbW/Wn7heLi7oZk2DBMVFy7/GZ5eg0KBYiXw66XzLCoaM0SyKL9Nhqk0PnNc
DIWEe7NL8t3A3v55Z7LyycWJKVYQ2lujOVGf72hn/Ydh1cpuDp4KckqXJOm0pqCk
W3BcOPi8H1fBTH3GtkiTbFu9oUVxgAtIxvyJ+l1eD27FmbPJHQhUGuXnEEWurfmw
PerQPJNJlJM10JuaIhSd7nFItxoJKcnZhpPV4Gje44ojBrYMqV1cpIarFfgc3j+p
nBYZBc7uCPgtPLLsxkGDayQHj9DgBH9wxe1e+C7DUm62SJ7C2AqWAfnYrjRvpSrH
OXN3m/TLGz/MxduqcSh1donxtQymxUFb4kHDFqvT/2S6C2G/YAlNMHGxrnACXL2K
WKvJW3THbiVFQy82SorSHmfrRAgrmtLAF3F6sLubGulXQu0m0mmISW043BnvStMF
BGu6swy1vcOc15eNR0NuRwqC6oOy8EI1TLLDfFH8tVusD+ZRvUpJV4L8Sc7PlljJ
dJFv4RV2FAPiSh1xULCk+/y4kZOpOoXr1QDIngiPgqZAgRNHIf6A72SVXcaqUhhD
Rw8EpglR+rPF35Y7NH8JFADOhlyOa2nNsxEN5zArDzeD8/16bnmddRY+8GMK0Ty+
Y3IKLpBYOsAIVNATzlWXcan2vxOgPExHDF4oYSxtP2YZS29vfyedSQvHCL0VzRjc
VFsZr+VUkbBPhDm4EUDIpEeFQSaVhcJwdHVwgkgYYGsgWmxptUExmJpcGMagV+Pn
wFEsCacTsVQWaJQPBwyyL41rShmOJYBkC+MIZyw9CaSw+nnAxmI+IQDoQpe8Z/mC
ZlDdNd/9dUtQn6zOU5mK55VSVLO8LCMi/o21i1giNibikKd9i3lEoIMjXSJyVZ6n
uKHxiFPrIpi/UIXuXdmXVA7Cz97iMpftDLxChKqOIIxOoQgNs37F3WiuUMTJNcXE
fTAbXWAzqML0mlA6nEdnoGcTvjuN5Xqq8wWr3JCfGmqe8UVQaC+ACXPXcofxiyFS
os3+yNZjFX2i66bXfWVKk66P15cnvfQEesrE4VRCjGzmqxYs7JM4tWF1hXWhegev
flH+Ur7VT/ov0sMzdmJ5IM22FhyKKZvCR6EWfq/xTr2Iy0F3uQg7yYq5riZ5hjl7
Ju5gfnd9O6BqFA4UCwsUeCJtC4fjetWuceCZ4L7TFh8WHo7n6v1Fy5h7vzWWfq7i
gaz/RLDnW2b+DziLgfXZYHYD+8vELKEL2gBPPlHar9o/BLFxEEFL7sPIk9uRngU+
U8Xx53eKuxuI8vzoUxJ0uJyb9taG/UDMpP4SnP3TcQ5dvM4573kI4vC1z6i7p/UE
8EQTrOXy5oLE8/G4LpYfMwa0ybKkYaEUJI8Usbfa8ioE6kS5K8nLSftay6EeTjv4
iEFrisSedXaWq5t/lvESFUMd+70AV8FQbsQCLeVBV5BllNLrTBYADgUVJuTwss5m
5J+xgB7qGJhjg8230VZKc/NcJZ2kXy9KUwnEINHVnD+3uZtiob4uRHSs2EHi4flZ
Nvp5crk750Avjn81MMdp7M485ZFNhEqouv4r+x4ewW/BsBoWzpDgQWrImcxEa0wG
gZSsR8dl/IVAOxGmqwC1CQhXYr2yzodER6VFwtxlijItfAsqRHDk8zyLNGxfU/eC
+rXXPS3AN21nUSYS4Wm5CKRdhX7wC1F+bnfwV/hpX9ujkoOa2DwNgRubtrcuh3Je
BB9Cl7+lDOh/AJX4dYaqQtPj75vzvgB3NN/PJEpn/PsOJpMPbCFpcAiYT9stqjAu
IiQ6S2JjDwQflHIxlisRUfm/LAD0bzEVkuyrC4RIXsV1j4IOvrge77E2htuAy9St
1eyOBW0AQCkwI6zrTcvwMzxKe2v6F8A8MzG2viUusEoCE9Sff1Wi2s/pUQhjGM8w
v1kJ9PkunYBVrEMY8vAcdLPJqBqJWr2ttDuEetorRYgDJoCDl9ZHLh3YF5dcy/4s
tJy/0MBzny5pwg1q/1fUrOkLw4iSBU3vszBJjAKEkjTUvUDt74wjgssA3cjc6E6J
/QR0SdWcgg5hTWhItkyelGQH2eHPpoE7rvx5XUgPPZDNJCc1gzT/X3e7IGt4SXWU
mXxu/d2Q/0JkPZZC95z/YM3qMloPzKRDwPYMezKTqf3N36WsSkCDKFlWsVUBNiCM
ZoraptpeRMbclcUvvIdqd0Leq118X+C6SgX2Mvwy7RwyKID2WQox3eU8qmUV5xR3
hsZ8t9rAv8own12sp/kkORlY4WfdMOWasNT4kFe8cEFqJ+i/IrnBYYDPH9BUaovp
wXHu41IHPxthpzWBKoLLW91zTgBwifIy7tMvaFXWVZLnL1dYZkl0FxvBHZ+nh/tI
T6jWKhIext1PgvYz63503pBEE7yK+0eyhygkbA9ijk1DQdZP2YbmPPVnWW1nBZKf
boMlPHc0gS9TLUy+7PZz/omxWAWLrEJdA6RtziJZOzwRT9dv6dO0Wn1x2LxJ7HPC
t97nNIkoR+T9tn3Tu7nsZ64rr3xKpsCkMUobkikzgpsr5F55X9GsJA+/n/vubdT1
Dtw7HhlOeql8LWM+IAX1UElQ3yaza81UE2UdoAHX7lLyYv2r/8obAfEfwRKkwhEs
T8cI2IObjjPScNH+vClbJuho3TwE7oPtc08uTlTgi5J8s803wb48zwn8rr/0MeTQ
c0UYLUktiM4SKd2X0aEDIju0Su+XF2KBaCCMQBsw38nYtPj3DDMRptSq8RpW3skt
Z4wGgS1s1THm2F8ShVuNGbuC1P2JSz5Dprwa+zPWNoZbqKmcsFn2VQhQlLv/xOoM
3jQGjjrmIFeSjL2xfHTdXpqlcm+qQFYEBJvKUpMYijqU+hscUndnA3Ej4EAYGRjZ
P/rbMS4aUAU0z0wUZMwOdjmDpCv81//TOuECzVP1NvPiwg0CzR9JT0jnsbNOm5bi
vmrblQ1mBgh7WT0JBOq1Q1TCLN75lrVHfIF39jG3F8310jdOcQiRoy7Igd4IGZBp
SSslc0xilaObURsnDxqVr+Y+rLiJUDIkSJB0qT10Hp/SuLp2xG9TykrQAgMznaP9
vmfUoW7uXIWLTMD+WMK7XV2NhKehaIdXtatn8w0B6CeeTM9+fZq/xBIs7owyZsZs
bujhPYfba/XmoBy/SmLvizBUU6vwHzL8EPYGIMC0IDJcWp5qXSbkM9+45JdON3J1
R0whNQEuaDcfpg3BWuYWM2HvpQUO5NMLkikGGCSXh2XT2iIdkMDDCAEorQuS08kH
7cfF0LpiCAqjngOfUN/e0W/86dADuQq9P/ULmi9NAFYLrhvNv/Kyb8/69bBN7Jgm
toIeDw7XiuLJ1BuCd3CB8G+O+vWVjhPZGcPEPN997VVrPNhEQ2jteJExCRb1WwDa
wYEww14PxhfiElpXISn1mlKfh3OQ3zQh+x0s3AfsBQhPByY3+z+HT+k2mXwgjtX5
7aKJz34RYWpscF/okvz8jqDvVDIeWfVFo0n8+KB69k1M/jvyhWSMjgPB7esra8h/
EKlfpbOk+OJPBF8C8QCmot28xDZuhBpeEhIcY1wzNYX5hWSg/gIrlcHPuAif62CO
XwNr2W8y1ZxYHYfycDdOZehEXiAiR21e1SVnZgxu1nfnabM4duLC3IpKfm4wcmWe
gYUtpMpyBqGae3Xub4R17FWC8Zkr4XuJgTsGuvBsQMcG2hnPC8ZLgQKLwz7YO29M
BNJrrrY/lksvUolCvct+C2vY/AJoRYQ4rEbfd/V3MPCjtkznV3yYiMlKswiWeqc9
U64cxWr+Q3RZJ6PT2Rj0VmQhtPphz79z0QxR4FYA1W7aOq8/Pi20GQ493f5STlQ4
VOMB+Cn13WuDX4H+nOxpWsmtIMivNSsd9S5v55Wz+W4ozxhRTHuMwgxVwDHx/jev
vbIBKFnQ567oTA5y2PYi5nBcv7k4ROsegFMrXkt7LZ6/Q8qS7B7iBEOkvc6ylbZm
hLOufprwNiaNKOYYrs7X8AK7G1TtnHFDqZ9UaJ0nSW8RhtJQX3ydCGOQYmpfdiQY
pOK1WmDrnrWtDvBdBgiAV0kGZMEfqpRjUe2tReKb1DDZt5xUztca8AXbaRz8E07o
FV3t+rWZWcsVZmXsLMZXyWqRwB1QggOeX8rWOMdX2loD1HHwbM5l5JWZf3gK60dG
Xlfx18XuuHYEpMSnbvHdWOfoIqjVeysVn8WAui7yHFMQ1Ay/nPLrBEnpdndo4w7F
NYQVGSdjFVIaC6Ia7LFL+KNbxE44kVz3b1TSALNuDIKl459tTfW9cw5/roFzJsXa
+RoDy+NUOMiExJGxQOPPqfbGD/f9vJuQ+dLTG2AiCG/MieQ7raZKV43yJLgglt9g
WHQWTEzFxzmlGZ4tiOl/j/eC7NMTdbL2gruj29ln5BmhKPaWR282wC7078uOXVRy
sTjJoz9n3/quXRAt7mlYHnRppEHqDOBEoegkh1MnPdvzaokH6L5636StC4xlv6zF
w8PohaqFkqYM1BO6c4/wDJHdNPsS9ZoJAl5Z1QBJeFFxr1HuVMQr1OvHXA7OCj+b
a4nz58YtxraFnvFLs3/q9AMoWKK638xAGur+78BQ6Uu6aKtCFxI9HHAUffxl+AxG
h8FzYOQRITCK2C1HmBAfZjnMd7V26YO2bHehiA4Q8TNrKu096KLtIkUQoHSbviFE
TawncXyOgRdd+LTWOSKg6kt3UGCizc5LSF3kRegiObCxU9PhuhHjpFe6Mb4lOjY0
dE3UCbWMuekxliq1pGOdU4Slh7aMYt5tAwu0N0F25nRsaPNTDZBtNxYlGZjdduYs
RJZkgWx6GavESHFXnycfsa4sGNso4mcpEheP+/paMOf3bU8/MzpiIPRGwfUCr3pt
vwqLyuCxeFQaY1GOEDirIoziwZ0mMhud2Qkz+1H1vbQyUu/ss3/jaYglqjJHP03A
oLE0u2WtB2OfaDPVXGofFIO2DqR0HhHE/D2jHbRqofbNfQtAgQOmhewZnmIdQo67
E/0Zy/zT94TQrGGAoJ5e4SfdMfM6lpQeXpc+7yly2MGnEJv7/5oLArl77tWGqKYT
wOGIKqpIneSmouCSVQfCMmoXtUrpVYqqtYYPSiK2U6ibCnplkOT24t1IICgBTp3k
i5QZWnp2nzotCKtqg/aiUFN7r+KBfDAQPnuwK0QiKZfr2+/MLz2sBgcNXZzzJBHh
dj6zl6ROPqpLCc/r24btuJ6m7N5cxD+erf36d3eRKiYKi8Yp+SLmUXiNRK8Xjtzy
vUeytQCsuNz99ibZhlLdSE1MK5B8HjPJLRnXXGtVHIU2a26UhqVVoeIX1BiR2pHO
Qw8atMyExitYnxR8s35QkgiEZXikYfl9bEGAqSZLU9A/65Ja45dtz15DtUj9jTsb
wDc8xdZxr2eJ+wUS7EdsljdQImZ95/1Z02/8xPo/mVJb1ooivGZWDRcTczC+vovJ
olP3/JhbvVEDwpuwWxf40EL54ShGB7HNPRtyLZHoB/HvMb/DqKel25gPzTqo/61X
pXy8+D9ngpD9RKeo2p3Tv7nytXG4sjR0kywAop0nCJltwqtn3Vg0O8A0UhdMUmA5
DKQ/Niq+erP3pqmsXGvbQRGCHCQ5lwwV+wNQ0CT5xBA20Mc3BLp7Pwc71bX+ps7W
G5lR8KCSabU/RSScfXNJckn8TeN080sY4ci7AFEUTJN5yHfwczmxgmn5yPmZgd9u
UTEtjl+KtC9eS0rsrohNtzPXB8F612NHkvR3gCYhfuiumymtV8prjKZelZBmPSx/
p2xjDEcfS5afc9mPpqySytQhnZQoE0B8FngZIGxlLvNG9CzmGGVzgdr9TdNaGgXw
6lhEnHAZAUDQW68qymiYdQxS0PD3hr0W5i0eMcuPX7b30OqHP8V4CKZ93JhfvhB8
/0qf0x6tEuoK5WVWKy9BAhbzjA8KEFKc8QqMGMteQx+zVYPSJeO9z7xgNbBJPTE/
UBFwKV+wW1nWk0FqHR8AgzU0gg6f0V2inll+vG8FjRKwuXcifVCZ6IP0rdYJlyip
n3KrVLUI0nQbeVHO+B1aPFxKK5s5Apl+1A9p0oOU/UGN7eUjvjU/itZ4NUgaZIo+
b8uyUvN1S0XmbsBvdMbAhPd/KsBypVRM91t+wrCKXAyxKib2L8NoFznI4Y4h+YIE
vSxGIL/4gtDPtscQDkEO4HYhvTKeeTzYOfIfOzKdyx/0zLkJ0Kjpf7GOdaPidwU+
E/I12ZifSiPZknKl76CxB6bwH3/QIrPTmFrUp3sclp4RXf6FETAiHtXkzkgOZTXl
Ns6YqqgNw884M+vyKXSUDzMIVeSBFmHocMMWC0I72OxSbZlXX63it8vBRNG5ZhDh
MhtgIqzvNPQrUa3m6x24D9O6xFnqCVYYeWXM27sdLaiavxa1mMEEEVjkKtn4qIVT
eiHtaxpcwI4HqBhU+zjDK4Yfeytc+qHQoA9nIDlFbjLjS290eQfpsnp3bJtC+DKa
7oKrgofI4SelsSlLMumZZLUoHQKrmpnhAdluLX7A/jgZ7/tH5nD1xkSfO7/FTcs9
9y9PJBuY/uaHAgvNsHfv5Ts0TW8MrfoAD/F/hncJzTuynO9g2B59Hqdy1SrkStAp
aimhp/U0ut6A94wevnagKilRzDzDbUdJFscvmmedYm+OzgRcGAoMQ73eyO4Sx/hk
9DrCIhEc/mAODEmD0wCWhfEsscbGl8OBN0gRy0HK1va94ij4Owq5l8VHST7SOhXP
NM8gowOZb0yLAUsiGp5pWmRoVGQg2meY6SuL7m/zQcIaym/LVS1B6Sg1x5m3vNKK
prHVJfKy59I0jqOZNLPQ+383b/JcGke5Waa8YdRqinhxNrdJ+ui8Y0v9MjxBCKN1
RWSpFnDyl+pgTkoCvQgzG4DKTOxmrclidV4SjulNmyWtxut/lTnncQf7UPRRyh/a
aI/mmAtekyEsQhv78TMsnxdr8CUvooHsO4QpT0gIuFjNbSA7sUyojqGUd7eXTefS
Tn6ZBKs6V/O99VtfvjH/hdbyWyAlcbA1kGcOK1UEprFBHL7j8wEeCAr0Boyryaqu
DsybM++vMQ1eon2zdxjECk16EbFaoAVJqw0fJIEr8+dzBE0BOqMrHLwBWxOXwBlV
615rE+tDL1JRqrijGUCvtwC2wi7wlfS2r8VKRnnXdDnIEel7aIR+HfBiKBSec3TK
2YHZ5IuLSMadpGen5KrU9eEnVpFsxxK2nawTbVa931bNTVTw2DXfyIP+6WPjZ5iU
2McX11AblZW1ogle/qWVT+ss5oR50ols7B/dN7kouPyWD6LfjPi3efO6bpLnrcsL
n6Y9YJE8TKfoKHzef4l9EcdTbTZLrgIVghupXpjlzREOb1q5zQLK9canmkRQudHH
eU+U2AUdwXkW5O/8xqHYSdhST7AW5HSunzjT5cZ4+05r2FHLBL8lqhWjpHC6akw6
DiZ4NliX7wxypBSUsG5+SN+K26Ks9RDB82ys8QvaNF5ZjUvG+NqTwxBJY9rGQqpG
aBVLHpZ5XwDvGwtQSL7kf8on4RvQ2AZV65Hj2ZPagmfz1yXhQQPqkwbIXvAtgz2S
evD+9+xNOhu0bS7iTzkizqUNzdq9Nh42MCSmwitK1/pfY4HtMGLGUSHZRB/UqG1R
CwwR7z331CoKe4a0s4MMXa4U8KRcjs4n69DFQKvaMsGSBpp4VQjwYNP9/dwq8WFD
VXQiroFRHwFM2K/V69uR5BrU/VYtJ1kbMpYtZrihFc5FIdALncaS8plqtt1tUHNI
r8flLV/8C8wLP5mGdrrcEY+gUgFTC7UXx2TacfiFS/9IhjHsbTL8Mg9nYMVwoqKm
seU3m62TpBpq+Ic4RMHOgKLyELrLXh/UwFo7Fuw9wjD5UwSEkJmfzBBX7XFsWax9
31hgKPt4sKoN+F3IgUz0YD4rfz7oZpBVi92CeTeayvbODtphrbHvKEUWGdpdEdNu
NLvhvD8AsYvt4+Svr4RcBsxcXrr+f99mNEz3P8su8CSMFEmbirX/MCO2l45h5G2r
97xK1IDEXs/wm01TyKCmE7atZ+LPUTKZEbCCTOmVj3WMXdCLv498uJ9OVB+32L5+
vUHyhqv9qYHmywy7agUQu4ZGejD+euebrNAQQJh62v5sBVIbEg1QM3KhQRy63kUd
E9teC8ij/2Ma8Qi5gdIeWWvNG/FOZ8aW+G3lLb69C1ghLh1Pts9cDvBCRAH+nALE
kVhpnUMvP8WsWsL0noHGIpKSbjLj79BE6utDLfTDhtRKOzhWaTPav9t8wgAv4q9P
vZrepAUzbmM3qXTbmsIjGo6gSPA+qOCkl/hkScIcX4EzwNg/HjTFNSlsZ2v98SJz
StIMleOkAS6+P240J8uCRqkUwk3Q/3b/1sz+NSnMti/c/ZW3BHq3APIj3EwdLi6u
BwrJ2s9sBihijmGP85NusIsmTMNKV/66btpMysuoR6n1XuXZI/7akjtuIjveVtpj
+4QAA8ifMIklRbPoinABpfHhaWPK+RImOZKd7nJ23pe4RvHZ6z4tqoCu1pc9PEPR
j89uyPgsnc98mkmzU4eEa9/moI+nQgBgiBIAFi211Y+Xdq6o4zVvSSBmm5p34Tyu
0vllEXZPqNaMuqCOp7/EFGA8N4zrI3KrBlhCNVU1naZB/KlsOyUkTOWGs0ji/FG8
MxLHGlAI5bxclF32FOxzKD18C7yOARlsUVC/QxBXWs6165iKSr/8MCGH4toJXrMR
k/Z89qt5ll+RvG6muiblq7s4QT8UG7kLaWWo4QydqL46eYiXBy0++9y/0Mr62/Ao
yZItN80+U4562zkfdf4YEqORNazxzkB4d3OWiiKYpaXMvjcOHiTLmD3zcIfcVnIi
osW4PF+4MV35N3XrEpCfBlnESnsuq4dUZ9FNHobGcgpIh+Pk1NSQ7dgAUwMYFTQq
OsRlUnqKz5MK1eofMB3KlxvS9gP6jaF40A5O4MqtYAbElISdMy/gb1Lu/cT+xwcB
An+cSOBQnVgZYuFkELeHkIKx6tNsML3Dp5lY6F3VHKrtCW62rdpuU3jjw9lRAsy0
303P62BN22sLIaGi+KCNUpSir8tfNgY6uhKS4nZlg4mNRxM30lQJnoq0FznM1fSv
aMHEVOotEm8HyMfRnL7YVRQiOgcJJF2bJ1Vq9/3IkQCBgsdizwmga/7J1HSd1IqH
3YQYNzheGu2AJf0wROw+wnHeDa89CHSTVeSGt2oBtJoaND4tDGxFEVuHNagmDuV7
lxIXGkoLt+wRSXoRbDy1vQtIkhA78ZyAqsj3M8Zg30UZ9mBdfBPvSJuehuM8KsMs
MNwrhmTPL0ixk26W1SK1bzg25Ce/L80VeYpcvqAbhIRH+8MaaxkoPJDoY2YlV7+J
wtOYs1zNC7Ux3YDA5cL/KneEpu/nyVT+idxo37MoNmWhIo8seY+Z5naHxGY2FfMX
zX1imuW6DjcaFm+BEwTkrs1UnbSxkvPMgLXrBaP4+q2oizZjAtyOOOfBrgGO/y1V
MYGPITQGO24XR/sgfEwzJJUQgO/3OBmrPfkY3VxVr/nAqcUvgBXQWN+dMZotwqe3
3QFiKf8s7Wt4tpYyyPm+gsO5VUybBuwFH1/lL8zaRm3wE2f+Ibf62oQf3s8Nx3Wa
CJiswyczSuNhw/J2x7ZG5pos3SrPCNNqxBaVaVmrqEnDUcLc1Jmbxl4SPOApQig9
fkLxJNc4YSQf79Q2yQclFIYj4w2dk4BEXDm8NsixMFgrtl/4KJkYQZa4n9NweP/I
KH9Id09bKJahsrYtnVTtu3FzElpPF1gB4K+mN6TwUZxxNLffz0Ax11YLYT8mlcZJ
TNoJK3jGbmbPRlipFbeJLNVwGNmkOWP6YRGdYodAWu202PF5iDULr42bPmDwotqy
RPdlq0qBJxZIKQTsVWTo0Wi1+uw9NkkOT/DAPCKVc5H4GplL2vR1H1CS9CO2iP+l
zdp0Nci7PHO4XLH3x6RhJ7evuzjy1G3NmoY7oQpwUfb4yPjxDxPSxLKuS/tW4Ofp
h2j8s3fjPDzvOe3nSMWTgAH9cw9vhR8kNia+gDQ5bvhKFj9wnb6xza9Q2Io/YR31
A1dsbmOB29i9EFq6nR7bsmyqBOpc81G82T9qtk12NRBOMyHftYAs9g6qrYn3CLJ9
FlKKdpDt4TLDeDe56O3p17PccIVGpqxYBX7VTg3GxMKNTdDMOBAGXFQhrnLp/B6G
nKWYtlKOMyVoWV22BjtXO3jCU9tAtTHBS5drspPjNdCp8d+4YOU7Px7IK9V4u+DT
jSmDoSgryEeHJfIs1QUuUvqR64aUcrD5izBeU0AZYVzksMJsds3HEbbSs85qMeoe
AWFPYbAUvs9y1rB7kv27XBB1i/5VjOtrincB/4ok66c0K6ZpAHPr76I2SCpEfoF9
SDrn1oWIWCvUGVqpg5bgZ7/trmiPJKu6MRwbW2C3ybmY/EMV2NGo/53jZ1cTV4NG
3XouDqcxAzK7kC0Ioy4ptiu1Xb67lvv+oVfM+mUwryDkX3CxrWv0Jtr2sLFgTSdH
0ljpCNcx/ug72Yrw87gPhsdTdU53g/8Jzb+nVrAuh9ACUKLCj234AnIqy2cEnyR5
CDt0hWA++LgxrSJuKWtYvedZQIygjyHKzpr13WjANXhaDLK2kG1aSGA+PfzTxSI7
0ugo0hMikvsl/88KdK826eUbYu88DwtDt3w9qXfh92U8HB/0fILhU0hluueEnVe5
vz5a94cqyI/2xBFvMQaPatZc5XfBFfm3IeBvhfBsFYJszucxoMiVmhFqe+vzCqnY
rsQqxyghB0QbksWR1AchoWPcUNNnwTj1e284peuaLTqmDRTEb3LTaHxuwl+hR0FW
o8kms0E6DwHUMxe8sMtTxTMJYUooFJgQ13ghJkZtMhVEX7j7mn+JySLMuC4U5Bmb
/DZNQjKlE24SRIGcorl8U6uEWG9absSlpdP8VKlW0lrSeeZxG3xHdVRwLuz37jLn
Na/+QmCEew+JruIa20ZTCLIvI83gzcBExVqY0jfu5GWh/3quLJo63a0PjQak+uv/
Qt4O6sYol6aGf1m2zAMnqUbsJgnIbWrOPTzBSbOuM//DHZpGkjusY0FUbt0/77hJ
WZ6s1MRJRnmH87GukX2SVxnevfbsVnV3rFxEyOw5QOa8sB4TT5MPvw+VN9w8o354
Md1b+SqBnLsnRMB6quy8u/u+PzsaQT3EzqqK7oSBUoGlOtfYpuBY6wrk8+xu5rke
f/fmFx4vAJt5r6asyw90v9KISPih2mtCeoRdt71pW26LHL94UqBW1LyCQTzO15Ht
HOz4aGobLTx0NHrCRuM3MAziLxWfyJO57ybfOiti5XzKUuzOGJMTeitex3wT6oz2
2+HmPjJ9ovrbejR3lUKnm/Ttdz80eJN40k3ORyR4mb104JIG0frU0GVPqKmyPGZt
uCPw3/ZdR1VwmXfWz3T4e6rQQdsaM6O9x44jWAFFh2h3vOiVSRaJWM6q7IRKxXPz
K8y+cki5Va0kTfoDM6YrNpa+M2xi0GwDRHhEyOBlDikWpik0YsCfWprbH2uKcIrZ
78JrOLzBc8mpPturTgbEjk6HbrQTbZ4Dax5CCTCNiTvs7oM1G6G+UOgAYsOFzdbM
cg1/BhJ6/WmDe6CYvyPi/tFnHJRLzcNTHWSrwNWIVsaYufsv3dvA2zKjh7sSMhAX
J7ZrfcfJonkjZsyZcCyLwyK6NH/zLnPkPtfJaRRJE6LCnk4hWZ5EeU++hkQMRTpZ
Q2Rb9DdxChk2uCmNP+/U7/iAoMcmLpByhCPIsb2P4riMv4u6KOMED6Wy6ngQJp5G
zMD7KfrbhqM/JA0UPh4ecuvB1Dx9tVTnybC5QAtJ1hA4suyZroqN2eKbD1M7dc+S
5w1PKgfvV+V8eNu7gLTgfDwCJHs7G7hgL86tEw1DpiNadsAb2KU7t6sXvATr97zR
TcoDWbraIkYRMJYGNUmaFnckOTui7vNt4cduBGP5ylYRV94DhavDkXU8CT/KVYvd
sbtH44H6OHVl2t9Pp5K231ynhoBL6AD+qiLOkMXah5TGzIcaaBB4WlNhHCHoqCaB
R2cC/mL6R6qOgxrPxE/8uJzwhc7XRBN1FetI/zwxjDzHFgKkMH3d+i7FHR10FUZ1
l9020dBrV1dxBsJAqMRiYMdTqFQ/5sn5YbKclhT043Ihh9QieU6N8UNVLWj9PySm
8ffcUh3Fnam3fywDmHzV3Pi37JjTgms+RTv9v8FDKoD7Yt2qVdn8VRIsLohjHsRs
4QL54OsT+egnYHZqI80XGVotCqlpjQ+nDQpkCLoYadzmuHvMhPwcOzqilQNloEng
6BqWLik/QSj4kzEiT07fNuoz8zYU+XNRg0DirHROop9qjy818c8d91olRKwju9Ws
M0e+ByphdY+Oi3n+fnwGv5P6SCzhLWnM6h6NDFLRJWZ/w8uofYVW76JrxoAYa62t
4BFroxy21zfSTYc2/XrdYprf3IsiotSzXnQL1Bf3pGivrF1mP27Xrsdw/j2WegQD
eR0dn4lnjL/hcnCP0IEI7rQMNqegkJywDkBPweCauMEVIXzvdD7kDQCnx7/8Vt3a
QfUx4SqmN1yw0KN7/RwY5y+lhkwwduh2d1BK1rRtx9yiNAjc1wb3hRlagRn+0MSL
X4yc7yRUiceVdju5JEe5q/qkrh8rZ5ePIZMmrdGrvJynqOokbYpTuJV9RHA6Pntj
HHxF4AW5IUT4wJiuNyHvMRPy6etfWZuWf8shorMaTmLh7kCv80DgIIZQCkEL/cNh
eObne6uZEwxC0OhmBKf+qePHce+nk1DQYA7FBKC6OW/u84Yis1MF0jPjLBnwd95k
4HiGBVJeKWpB0omiVGDmkSdF29kRKrbKiY+P7l6oOOVV0g8Ke2nJ2EyZRkIojwzh
2lN+NCnRkzaboynXp077fjQzxzG8zOJ2UrSoaVdr9mUKv02rmMxmYP/JDuCXeYZY
LQLVHbK51c7lx6q18Qw5sJkb1dZrEwNh4wizXBuDiCJ6Evs2+G/oF6C8P+dBm4Ki
uXZiaeOnXTH2OiPK/HyrzOcxjTepaGYhOdaIYGWcnFgFs5sDKI46f3G7r1XF+jT1
+Uu9CfzLXGcuSt8v9U9u41pmvcFku5CbdGLd0OPmoiVf6zJkDj02oxZxnJVWGN27
cJ7tAwPlbfW1ihfceF9TSX/s7GI1Xnxj6rZx8gSN1WyEP1N1f2JO5+dR/ZipVW4x
n0ylTbdNFO6bwJYaGZA21CbQ7C0gZNWm7WQuOsWbLbX2vLT3mxqdB+6JbN+6YTwe
lD9D9JTiyIWK8AgmsQQYnxa9I7R7MD8ilkeIdeR5VywyVF85rZKwX2s4yaQP3nil
19iFuEVbUQqpBn5HGVSCAI3o3ce6Xqwq4LmSYH3fprOAS85Xr1/4CG5hv0Vlyj9M
RRIU0MVVfUbqALokMVUcgqQZ3cWZM1cyNVcTpqxBQ/mYN99lxbDXEDeMK/QmjyYR
MgUsDnW25KmjENMUV3GirPSy2tTcelSnAGRmNF8PNHSCCREmiH7bIsgo2UimGSXt
dbGAZSe4jValkGWD0quuLkhKdnaRSg5lGWOIFKU1oHY1avWnAT0+ck/uzqohfx+B
1iG0u0fcUxDJaoS7DrI3jm1PfJlCtSQGe76+jUm3SOI2M3BufSOTtChsNdRFOpgM
0O96eiBm+MkoeuWlTqFljeb0hhnjKMQzZkL02UChTCIDKv7QtzX3Mbf6Vb6wT8Gh
B8oiC/XB59kVrTU8gb9YUk7KR9PuvMJD4NdfaPiDn0uy6+8iBwQClb7X7x9tIk0R
LLLuxgyUssmB8xJgzmWDxkpu2oWCvYqVvfVkdZNff9+tJ0M2Mxt5vC3AoGZg9dlc
aCyStWPHONlp3VtpucTEsDubv/BOg5OVvFNUeRompaklBCt7LvBuY0dwlX+KJDcc
pqkreNGN8Rj0CbBEcTkw4IRBY7U4Va4tYzFJIMwBdcJ9Aj6f3Bn+jbCPky52STw2
2ubDFjWsZ+FESlndGmJEpHoRDBOm0pd7E2kSkEHpJDC9lZJS1JavhxLsoAgeeZkX
m4OCQziNqlQ/d4hc0VeLyyyzHmiv/FqRUuRPAPytJTPIwwuxwjLizTiIKiBlYA1/
FYFx9hWOrYpuIPBMS/+oKXPGlLCb4MfBu9UN5sMIV3XWzv5mz1vD3a9HZEkV2ib6
mOasjHhevjgsL4MlEJ1xTOQEQZG00nQnZ0CYmVX2NYub4bw8POanhaNOg7nxt3sa
Ap8VKg9xd1yf1/wq0bJg4l29JShG7X1YDu96EW+grcktq2yYOs1t7Y0ySw6IdTSh
qmxMafAnZ/ThOMHY+WW35Q/oKBOsp1rGtkEO+ZKV9dvfivLs3859k+g45Pi2cg1S
+FH485cOmRCwF8BBhpfhKZ2DZ3uj9zeBfvNu1NzBm9OwfZFddQMgsMtijlLXkkS1
ZbL8lrFck9qt7zkH79LArqwhvk1NpxpE90NJt1V+tHy5xx4cewOqN1t29zkdIMdd
3oP64EVJBia97nEG1TWjeyLm/0k7+JjqFwgpbsdDVqsThodl6/pLBDkqZ6cccElA
EyvGTjw/neQ7iqrHnFTxGuqtqkugN/koqJe8HtujukOmrwBv9nlTkxIG1L4tVbqG
09Hn3m+GRNGb29KR+6SNPbR4Iq/Jxz+pu45oSaHd3XePC9nB5MRC0CV++Ew4uYSk
QuLsrZQ1PmMkWIadqpek16TdKBanH1GoIx4BqOyW03cR72QzfdkPKhOplYCp7H8w
MSpqOw9qcS8AkdrYxsHuGqHAZ3Vh/fCemvS8WaZzX7al6LOOAK0fb3Or7xRxsnUE
kqDHwMYuCWDAYGoOeia1+hgkBZdpK4Qeid1K6davSlU4T7dSPadCbVawNP0YniZ8
klP2QLAmSMa/Moe2ecYJwXqrrrxu2tCba3YflY9CP9Z6GV6LIrDqVqua93WisG3l
2MJ//SPx5q6A5lh2BEeKJLWp+WcJKsCbWwg33s5ylZ++lSSvzsof4tc5z66mFxp5
1Tmf0K+pm0b9ozLKTZSDUjSTI1LTQ5ukSYK+bSXvjYzhiWRQfDajKa3HJIe1Ye6n
5wdtOy5Wml+P5WrXbC5H5qJ9krWTyZgq715usDi5P/56NZG9JKk1Rvc06+G2OKLX
pSU2exr36sUaazGj3Wf0Ic71ZfTGHVWNZ3tMYkhYx1dzU/PShv+QbPVYqPQWEfxZ
HrqBz2eb+lI5NqEzmfgwRKGsYyLOkw/iAG6+gRBxuJlGCC/0oicWDm/lH+eCo+Ty
B1CXt1Ss0scRnp3M+N+Bl9iH+RRYGLtyxhZLu/XBaCoz8aW+5KKRlZsfueO0S9mf
Qu0wYSTNRzmuY1rx3SSsY1uGjRCgv1utIQ6K3cbpn4FUEN0hoAe0L3NJFyqPMepQ
O422liygMwe01RV5NN/5tOyKhzsSIgLLK3Za9jgo6gLxaRPDfHRZdPoOWJSz/eai
uEw4BSuvRijXbczmroi5ob50doMFXrSzprcxXg3Ci3Gb7bHp0SNOUFLHcEW1wP8Z
ZC4f+jS/ImuvOtG87GcpxoNvk0qc1nc9i9tdAonLfMyJTv+LCNx2+o2JTP+aN7ZC
M6nMlpVe3nnbXnX70deN0RXqAPb4iG6mNT/Bw+w3DaV9qYLuSV+DgVEEIy33Pm3W
5cwjlhSVt+boh6ZfpiJgE6m8lrsA0/UXEA+IwV5kiDb2bbSe0ILqFOFVPMjbG7He
vy0KB4+/9psLFD5yJMWZTNsFx/qWnIwwcsajeCSopWzAXt6KLr1TpWZ/loICgKsQ
fPuO5rVw/sa3IggYC+pqtyNUHtJFDz/P3h96GhpTNUTJZyNvR+EcIY4J90Acu+SG
OosN2njH4xVGjAggbTS6OXgmZroFmgOR5uNxEETJ2awdUUrU4XBsNiaDFK7dsf4J
J7uvyb4IoDJcc/DTxgoeCKelAjaLc+/351lPpb9opBGXOKAbitBfBiYQPhlerny2
aPrp1NDEJxF1oF2Q+QfE9W4nIG5FknCSGVPRj9MaboEfsxrqbrzkaydHw/onLiqc
PWcf3Ub/2KPMxlkNKdZlr2R8B85c1VPIABlmLrBLRnSO0LOiM4XvFu/VDs7Y3Saa
Z+J3/iUcoqeaHjNcrHg4nrUTFnt2zdQ8E6fOGw1WxrfQtIuFxPG53AG3c5/ooy/+
8O7w1tj4czPwWe8DwgPJIavIzUoCd5msxBf7He3aTmB/jt3fZwla5Gwq2LJSEhlV
nq5ImM3WBVsbH8VO9ACdzds83TCx7hCRRXvbIiq1GOrzxcFjm8uxyyFylxSaVlzS
JrLI+hybOzW3NhM/fwaGTcOGIJLEL46BmkJQ9toTZ0w6Rlgrh705r9fISlWAbooU
R9oRhSEa21dCgCgqPJWuCONrPFnBwMTzoaW9P/keeqmFK+TyjvosMNcQDLZuNQAS
3Zbe/G3FZHJ3mHGNgnNXs8xvCyVmctKUVfYfybO02eR8Q7eofgpcWlu/eMGHFNd8
RGw6UWIxOTYDRvT0F/C0naDilrqARksXT2DFLenlFMTpYlgGrmKFKOpjiusbW6W8
6+CpcHFifCE8Q89+X7wCA/19niOnU2V0JpSGDMrtrhVpB9VhCZi0Scg+y7igCjag
vAGFMnxccPMgbATEmKjyWfdmflB50fWuhNQiH6qaHcYBQmgLTEf+WruFHfgCwrDr
W6vezzCKX3QRUgEKVw6AYR+zWxG9BjWH6fqkOA0gJgnQEZJDMWuRQi8049v0Pc5K
Iui6P+3iLmu2l6YcpANm2QW37EyGzZ1MGnIgFFXUsJgfbUrzPr+U4RHuCnDw/6pS
wfyLiDw1jXt+jGWcHZ3qGRWaDkSxs/1kmTrmP5WCM54lM/1aVjt0RwTQTY8abKGr
XVJcNwLioM6LiIm32IvhTo37ZxFjLww63HThL2Zd39lzAPoYWGdPq8gRnpvqmfLk
7XgX6Q1DSxabnRQNyfyQrmebIce+KOJsgQw3LY7MLILy0KVFP1dhXYlr+pkq0OuK
zJOQUfMnT2B/XW3djVqeIlDaUyaV6xzldkmT9qelzvuHGc5+ptCrXqRuf0Glk3bV
1NIlE0AmwlOj1nBEDZRlR2xRTvSTk14F5QEW1OupmNkMI2tOcMvJYcv95aL6p1hl
UY8Ow8ns7R0QQElIU1ylIcph967bvHAhIUDZsmUK9IIVT5BYtQAUDk8TUebw57i0
XEQBC9Jayrv0e2JML+xxgdypa4MrENK2Nx8NLgzIbuZ6ZqR/tvs3KYl0Qm5W/vV3
uSfVBuuw+VMe0ge6WibL+/oThhBCgFzjWHiegy0yfddZJ50OKZlVmoqbon1I/TlV
SErQ47xkqBhHWlNA7J3mgqJQbwN1dEQgDByAmvrBpBeYsSVt6rqKvyYytQsvV1Ta
kSYfdMIet2WJOKGixjx7N6Kqe3RkuchPmypflXeX8e5MNb1uGa2qmY4qzplqYZLz
hWhkn+kJG02yuUh0JJTcmurtn6S6E918feit6/UmwQGjUkUN53G2qN4a7AEjZyun
QAAsVhywCFXGXrUzp7qrjGjqKr19q/F9ul9qMtO+2efWmO5Hm8n5ID9QHqqBn2ee
OmaTMqe7it3eivqZmJosxyeC/ZIMy8je0lV7u8iPZJ/Qg4U8RVNuvIXDpdEQaTtW
naLiJiAowJGq1jW4TreIMX+3YLyAIZgc5jJsPyrpria7fHNoSHfMR/aGgQR5wiPz
k4UnHcxEa/FX/AlBQd5ZTKYsGfvV9mQO+b2HQQ07TSw1iEzWNXwX39mxR0VhvpCo
oKCSn257O9+5v7QLt63eNetfaLxrJ31m5h55w8vs0C5V8qBZ0U3T3gnRW4IBJRNm
dtdzdyQptUf3niRRv03f2MrCsPQ6RKar/jXGz2idztjN3wNExgsFx8LKe0VrK5O3
5YreuYFC4LC8J0c3s7n/5xMOAulBlbWydy2Q0Qh7zPJWgoPWrJJtQIngrvSKxN8v
EjOI86RMm1QIOVNKtCJ0AsyU0kdQOPU1LrbNtTpEPykGDxB1wrFnihUFXLOQxvrC
xfaJ5sz3gTXT4aLP8hOJLi8vXWH5iz9/ijxQ40PtWk2JlJ7BeMQ0bqs8nLkanLNM
gLbpmK6tHYNDK02T/Sy58KjhIzJsqAvNcnBdvPCezoZxXn9iGtI8WCAXrZ/ZrMIn
rXgZR2oCVDTXqlQddMyJYu4UjdFhrvIDIiZQrl7Qjm33i2TjhncuUziciokfcOFO
EJr6BX3i4AUpkLE/OYrBEqWGISa5qbQAszmCnjiACszQGsJ+mVPkufcbikFTTZHe
PFJx9jCkP+U+OMp0mHXhKCxTr8oZNgPam3Ct0WpHE7tXTWdwOqoW/cMHC9zi/Vqk
hHeM/sMK+ilNx71xovuPUxFpPfTZJLL8li7BZZ7Hm6ffmq5nJTfuCrlz+zJjtK1l
BV77pR8m/IceshGFQjCKIAIkotprFWev8RKM0xS+r1tse2WS4S9zGb1s/a4yKef2
JlJ9ppBIadtZv/6BxsmgiLxemKzIESrCfvUjCzrjVhKehm0ciakBp6eTDnUqzGe2
otEkGnbgn6IOcIXeOoifQADqhCXWCS85AgIAxo5zHal4PXCYI08eB5q7lUe9MIC9
NqYPBW3BuxvkoWHl4r9UvOBA8+IchW7IYgD+793BXdpWkLN5A0YDbPMUy1Vmb4ja
vgBBC5Q/GYqlYTBlUyYo0o/QpnYtZsapoX8eaLsbVp6GrYO2LnY8+L1E2V7fdxEl
gCMFeKT8N8xBE2pZNGdSUJPm6DnLSC/CzfFzR3RQThqrj/yl/LX7xj5qzJttxBxE
igPoPfVpYOuiIJGoV1tDITHAP5YDbsAdAw50csQZ3cj1bH/Opxz3RVFijxAQJ9R5
4wNJWd6zRdl6/H36eCszuSVFBXMlHwLCTV0G9DOl8nEbcja17oO7a0T+/53pv0NI
aGZ1jr1puYMWdsBULwevno9q4tlFi/A2k/6+cg1ejtlBBeLm8S9bHLx+9ynRfK8C
ahD50UcI4slToOAEXYPgcvolOTBr+AWS6PJqqYGCnyARGb0QDU8tAUQziTrvtCZs
LpjwHNZmSpCJzQ1lmSBpZgyht5kTlwsF6X6rOSio0bi1INdNJEn8p5ohcInB8bQg
c63pHSw7StzJVzeM2Yh1IjQR+3TX+2OQzkulUFwp21EFOgXtWDvwQytun8WDZuxh
PJvUgGLLG7CjN1RK2y1vd7DwK288m0CKuRQBZ5NzyTn7G8ao9Wu8GjVTj+CDCAQm
R+7cyJeSTw8k66ig+5VOszyOOlO66sUErCekD/uhJB2k0cNhVdqHM5Ssoa7G/7P1
xfQtOIirDkPm7JzYH9BEzdlRNslgPl3kp66hhTv5SZk0lj6OOi99nf+sErjtlRWd
hIqgepvPx0+noZAa9z7JazZhdLfwim+Bor7Pzx0Bao+UgDWXMDjEWxlQy3WdvupF
AYm9w6wPy/GuP+npAe2qs+WEZb5FANb5JwZEcCw6j1X5nWC8+ApmLTHky4QffuQp
6wkXEwy5YKddLzzBB5gYGIRcqDp+tmjbxfC0ghTsJCY3ylL4qoPOQZWMCcRDZieh
4jSK4VphQsUEFkJzj/Idu+++7pHOLyLpzuz0Bmk/0cyKQU/btlU2AtK4u0OmlypY
Ifr+uHFRKEqDCiLUN9dewYSFFIx85yVTL9YemYdJe2Ll0wR4j+FRFdZQ2R4heSHb
f6goDAUBEsz8xy/2Fk0ZOPWpQ1T/bekmDJV6gPQ/qcPCROpaREAkE7PdWH0Rg7N1
5c3eHlMP+nLafQTYj2vF6XxhWt+5AZhflt6wUN2HJbKjUcSDXj3CX9FfP+W7CveT
iXA6KlPQbW8EcagaKfCRStltrOrtB65dXwdZI8XD5YhQWN00Guczo7DPn/I4H0jW
DnjVSoJdsgBm4x8i9h2F8EgK3fC6DduyV/QkEgGBo+ELU7l/P1IPL1MP/QqTT2+Z
FFodvgpVjHmUqHEzKBKAHmMQnGBWd6ycsYy61fePU1Cvg0iB92R+YfOz3+YJEZRN
RwtW2boh01hSp10JOv+uKiQIynxOxGKiUecrEw+gqUcaasfsa25Z9yRLGlRd8QVN
U/+VSCQ7lfhpZICB5AUCSl/AMxaERpbhGn1E5Tks2nlMwSlV03Z2DHOD58kNDqnc
fIE5xUQHMZBGdGR2pCnpEnTbmcfGsNAt3uHumEnUmSK8yoBeyMrR8Wyh/iS4gOtJ
hDYM1t86pGMYxbCaoUrJ0CmVLI5E0cOpIQSW8t+QJ+5FZLCrsbt8LZomeW0GZZe5
JyVaeGar77Pq/UdBC+PZNXi9LB6TLHFasXj78mtoNoMff6i1Jcme8k+0AfJm87Al
VCUqd549d14pLAoZ+xURJhdRA/8Od3pzA/RiAyZzTVEv69tsbFEys8fBooToz132
A6uA3iVu2tY9L6hnLgoJIQNVnI9rUFNmFTCBzw7ANhgiL5CkWQsnJXd7F/6bpzTp
nGIKN8sa/9awWWC9zdM0tz1JHLzx5C80p1/5F+kbHskp0ghXQM8HAzrJSvNqH2xw
x9H1DFk/sPn70MM/2y3AjkgCG7O9SpwBS/oUTgHYwn++UBMZC1/OiH4FQ/J+najU
VZW/r/rE10rcNPAXzs/XULFfDY9lJPZUBhBdC20YYqPifSZhrovfkQsQ1IYtMNN6
l7KQJ7NCT6lHaVkxy0Y/GhLvy9gEO6uweg00b1AoB43Z6FDE53ZmWksIR5ArUOtz
gFaV4me6sFnfUVjG+dm9VRIDHShGYI7jnbBlnhX0eGhj4c6i1qDZIOEXcDZWGvCR
WEcO/bA5Xdw1D4wM5FMfsLuzgKRPx0xJzvYbMyCIdr4TBILgpqC2PI9MbUVtyYjc
bF+7TqL8zguU61TpHp8urEMAgcZL9HTh2q88OFljJjKSDVxCqilv0AeB1dOpAWun
RCdS8mumUrkS8LJyqulc6nqmEcjX9dyjxXJgLZp7vPwnzX0QvKInIO0Br2uHPeIC
+t1TGw18RpkLH904sMXk0k4E6VGheO5zEiDSsmkBirFuSIW7ncQL8lxi0B86iLq+
UPWG4NM2eB+FJb9PZPgAHUQrsHIfHy8jjceqLxf21Ip03NbYKrCMhvm2rkTK2DQx
DZjm7+qyR+ZZZN2YX5OmNMlXcG+fTDWnjyJny3jV5oDCqv01/Cu7jow7sQ59mW8B
RSVHa/XVoRLpYB7oBnS4Ib9QZRm2VNDtnT2iS/Q5SO6sFI5lTsuFnREmXKh3BFJV
zgrnXHAO1Omh5oGQmrX1d9ocFanZC8L3U3qadW/6S8HRsaW6wHq0xmWVPgb6dnAb
vuxXKS389dYA+mQfPiiaqsu3gMjED/GVsJlUYLLfuwcoc59AXvRN6J4ghb6vAQgp
tU/3YFO5DULTxCIdelv7iisCUVSa30LOIgIQiV292wcFvc3sudBtl4aHAzVVlgnZ
kmdotSr6P/O1oeTEmKceSY0GwwzEVExGkZ8PJ+QODFW2FE8+Nl9b7QmmO9QntUHa
qozelroPyRoqiooYFX08J1Y31/lOk/h+31oFy3+ME1pIPBZUJQ4zY1U36H4ZeeoG
dQZSKEmeJwvmWpdMQGWubdnPr4yWc5GAlqr7itzCWoAF69c8FM/mIKJMX2ozafzx
eyv02Yf9wjXhbzPZ533NO7Fi1u3PczrSfVkpezzYmZl1IC6t+PE/TL1yBMhTxWN0
QoAAEAdmdLdcwoT87G6cDBkKwKDn0OpB6bszLS9m5ssdfsUzAAuaWEKKQitAESwW
3aqEjDy3OCILqdSQIzkjo4D6zbBkUW5Q8/yrW1t1cQvfVRUEQ++8iwbvo+xiAHoC
D/UP0l3iMB5sDzLRleBshCOsHlMaTq2k09RNk5YEK24V/DJt3O1loOq0zyyFpnWK
1RjTaOgUErucosgDkfk3CaT9AyS/KBL9ddjrdP4xefqzhWBbdBd25b+qgb3IEUxU
/SlKuRg2ATKAbJbmlqSZvxXCFXLdeFOeyptCv09X2KtkA2V4KRcb4XiaOn2dxcNN
iAnbg6nEPaQlCfsV2kRu5xr5skH/rd7WzP3lS/w0UCClNpdvQjuDsfI1YxDzxaQ+
WwC5EVps2wgKNpG3qXI0aG7r2FBPt8+yo7q4McJEWZ5fYJmSM0NSpNglb3FU2OPx
y0jgjLFXfgaQWdaUffRdM2dJh5n+wu594pcSS3lznbiJ+YB/mSsw6v8JFhiv11f5
N8THXA51kfbLcr9h7n034FNIqQSub9kbG6eg9V5GkkYsO4pAeHUgqI1U/k9a2UaS
TIa2haW59Rk9Yy9SMgohLINlFkkdXmQ+hd2Xaz7+vnV6sg9GVwSfwbSu+k0jcQpd
AWgJeTOIYHnM+pbEQ2ZTbu2euiYxup6JUwv0mQF3SW3bn+4wK4GJewAUro3B67xv
v7yV6uSy+nM3qSIvnMMQiNS8XCGb6PIpe6nNKbOZHaY186dsI4s9lmYwRgE6qkrR
AOUWSrEeIxH7Uf0AWU9cirJig0Vo/0MaFM81UY+WPH/YQUvHYH1gYwWHrcTrUxaQ
AYLpy4enrgGvt0CKax7GRCkGyNtLqyzaZdMX5gkmDb5EbZaPEi+hPHlZDg0/CQ2B
/HbVzd1D5mS9SeQEXt+T08lnEPxTWG1Sh6g9/C2MYrImGCE5KcPNN6Dd2uohE0vv
cZBI9WKeYeF4guCBaA+FsTkG+cR2IjacVBL/e6BVyzbY2fh7CKe51I0fFmdK/1jK
Swhr1yTitIkvNLcXtnRSo2x4CPCS0tlLVQVid5u+qsm1kw8AeL10NbQrfHtLF7/s
GS8fKzaL1uEj96TJSMBiV7xVx9HhGyeh94GdNptwatih2wlVtBWgo/T2kPceFf6Y
Zhw1IG7kB5Fkf6GZiaoV8Q6EFExxRmw23gFjjG3qOY/4gVvFOtbrs3gqnKWdmJuw
j5vmWaax3qB9HFw+iGCa7x8M7LWcyikddoZ770N+Bapu2urBe/6rCN2aH986z+wq
VDYp3/+r4uBnXX/8ErlpEylIKux6kD9HLxENnU2UhWRQEcWO2YI1vzUrzZrbeYbA
bn08SEXxJ4RE7pykNOlBEK8LzaHCBIyirPrGx1gKnHqiIjCWqCCWmGICDQ9yzArD
kwmDaLcj5t8GAkhirDjcPcErHIBsY1V1srPKH2ABr4dH3XcbxgdByscF0wk6n2Ls
PLgCXlPcoFKEBqJ4AgLKRGNsbAHZ4rMqqP3FxEwfGETNuQbIiHQDSDGyGgMNgCC3
JWh8GJlrHe0vemRseS5Aw/arB8EQSKLqJo75g6ImHm0LfoVeBtsItDsyPSizMY2p
HtdnQv5c5YiqmMs29Zw6Wxqyo83DN8FfLQrFsL9LLC3XB0+RZ8K9udmLm9utzlU4
rBQhkTaG/BkmlPX7R7IaPDE5ur7kypf06ReX68bVP72kQRCMJjoCCjZ0KIvlm61W
dNydS9ZhpMPMRmlGH/7xmVuZ2LGgYqEZ8lVy/+Qb5EYTZX50jp3VH2STp9EG7It3
Ja6iJkAbaLK5j3KHTxTG9rGTDA5/tApzmep+HILhH7ZpcnXp/sswk4/76xRGtQRK
YlxUvR6b2diDDUMBeB6WtFPuxx7jMt1nHvGm0iNiH03R/MoK8g0L47s/AP5RXgDc
jI2RfYAp1WK+aRHIma75tP1gmwXnWhXpQpXMGbmLE4YEZbPTHden/EUkZvGPdNzZ
Bl1piEj/XHyDS71ynLLVUWtpaxxxdhrIBJ/N10l1kWvXSOyo0+4hFmgks2lK+dTh
N2UZSRVwRS9MvHvpaIRg4x46uQPkUk+ahxtvq9JXQmofAof3Ng9nYD/u5aF/4DCF
zFFFgdIZAyFeScBsQWUriIXL7zhHbKWjiWDP7hkkauSL1itg5LZ00kWHb1omTy/3
0wAcnVFoi1Za6m0KIDYbAfZ9W8kLbjGSEVC6dgiFJqb9bYBx8rtY90o2VZFzMibf
TbNBlWLDD4mh6RhGUTCJo+F1Uvx33kdm5h7RHg4z4STFdO6P0XczmPMz54kLHmRB
xBZpSHSjQH3kZHTt+RfxtrbfFYwOajxjNdwKfla2jY7+IiCzU6kMcxsMqRHKi3qG
vIPkNIWfqNNoT1iZc9HIy5IcF6/g4/JYT8Pl8bP6Dzxvfuf+GNdbO8FeiTx+N/TT
b+F4RvD9O26CTB3bKRolORso6L5NIzi+IgoQTrKDjLZvOyXvl37JG1A1u2k5fzux
8wzNO24nGh9Q81fMV8b4PvwuoSEZ3DzgZhUWq8zmAl+QyOT+E4p7Js+y4rcfaCGI
qRwEZuY6N1ZA40hu/QcfXjf3sI1JuvzXX3i0sy4m0KfLyWLmpcfx9CwrnWgnNlUV
kqA8fsqUDUwlt0Cf3cmPXieE8IfTFdJF9ACz8bWSNgrl/usBVvuCXdQ32KewHHvN
ZDGb0Ufa6ZTWEJSeGW/EqqfiusjgAIsJ9pGx6rgo6YpfgYDgoecYdLZS+CX97UVc
g9CmWb2eeExMoaxgmeccuvjRkSlfibjEe0qCiP+MRrEx65QRoNzocP0tpQCjBl/d
tyhy44JgLvJc5F2iZg59wV4D5R1tYS5O9ucJnIZ0qsF9rlnYXFJZBf7OEPjhJX4l
ctI/Yo/g2aEmac+P0oYsBBXn/uECtDw8FNLddmvLSM3CYjgMfqUDeNKxG0x22DUl
T1qgoCc2N5vmsZMK4E8JSVU3SfIm78hmRgOhb0kPsCImC4aCiAM/Jl3GoppHgwFp
QYvOoa6YAPmSA3H6JjqkImlanTaNeZawzOs0QQmn/qFaCoZhxcT+yQDIglHEVEKW
IThrEl5lbZoCgE09NEQf/ucLnSdSfmfQCcKBsWm7O5Ep/cb4Kpul1SX41YVVMa6d
zW93e86tFzxFhCoPsXxBlKng6EkdDFLGOymkJi1qjxJtzIgt7ymDJFrm5Bl3C3rk
JdfXmQfLF1vTEDbeIfrx5LWx+BUZzUYdZMCcmjZgNzTiugrcgID5NjZhoi2alklg
HgLgL8/vDcrFjp3K7I64SLmhg8Dp3PtIoMH2IRv1JjWahWC54BNyaXx1VHddgF4L
hAB9eWQwFdGgq9SpgoWd6Km4l9FFodDb3Cg3LYmrfb2TMT/nVvc6VNVM8eLRsYIY
VLW8Bj8R4OjWznTAow9ZKO4SfXN/0lJRpTegZK8GpW25feViz0zd4tO7EjaWmSi4
WbayW0JHhUhDd4VuT04YktGqem0LJLj+YgAF0u+2fNIF1t99bk1snFm0DIJXKD1e
Ylkm0KkAxIjZoH1odI4HiriA+ZV21D8gPUnpNAOvOHP/7f/4Ux1kXw6Sxc4vUr4H
GCmYprb/65Ps5IROz0nMY4wZuHUwSq1ndn8rA3FQgwuVQLEIm1NVz+sAZFxl5AwJ
FyACR8az3vHOUCSBtDVfZxJ1o6XbNVxxeiGr5U9+MSbZTOLFfVRxKJUK1flLtoMh
exq2cwll7tH2iHceHoJYHEtj8FhZsPuDPhPaFOo2GQHaa8FeWv9yPaaVRlCSBeXI
ISXp4pRWCapjWy3L3yvFigyYiNOqDX27HIjBTUIkwNPgpfTBkAgcH60qrxfVDvAi
oYsl09FtsvjS0JQgppojRX0ug+SWA/sBXKq6l2yPjErLf4XozStCSh3wwdJAJlC8
KCwM2x0ZUNuCeHarDcSGu2ePk1jP5W2ozlmc39tdnRiDeG+DfwAn8ZcTqvYbHOhZ
4J4ahy1mpSHzi5IJc4xg6zAMwTKHnMIQ5N5oDf/qmYzqY5/0THjyzcBPfWMZ92r3
z8Q2Xck0jUWXnUv3hIyHMj9ej96WJZk1+t49q6gtcJVBu3a1LAXSJurlqU57E0F8
e6swJkFHP0JgND+ymTgciyqsDIZKFoY2mUI9le+CHtlafG3qn/1g0en0qAg4OsWh
ujTgjUmifBLP1KoWIycN9trEKBuNgAt6ifM0quLaG5LxvevFW0uyHRQVlTrAiXPk
IgURHK5JXqSJdTLTmfkCgi7Lm19PlrCNAChRXvCDJI3cO/Z0mFPzydpd7COWdL1A
H+zxWt5F8nLx4F4VhW+oxhP+cQ5D05DkiGiwgu5Ktd0aniC59cB/oUyp4vdQ9HzA
7wWxvRs2h75Ol1bWTqT77i/pomb81TWH7FuyqLUIzKQcw3RNUkeiKunfQ6+saixU
ZqNbUYShn1Z4D5ny5OvvL+oPfCFUcVb3/xMSbRmGDP4DTgkcHfd8tkpW5+SgGabH
5pojWOZSttCof8i8sz2FvFVYThraDAnChLwMigNYIzfaqH0Yv9kpdkQ0THkUV3o6
wrjAk5NdMoRiqD9AW9jjmEfJE3KnoX0+8zu+Pc70i26C8wnHlDTQKvUblLskMTO1
Zn+BWA2AaJ9Qu0SuixYIsMghWn8fNAvB4XuYBeJs0MkSSoskjGgmgufME73ozsCt
plRo9S2fU9fDfzcgHlMRXgMOBYUWbCkoWtzMNUGsfcqRi1S98xYg8nFMZlBi21YN
qSDy1ABuIJQnCP5BraENYd6PbHxqND8J1SEYShPAaXQmM9SP85KiDOvtFMRZQGSV
dQeO3GaVz45O8HaJ5CyyZUT3Zg7b4RksnHjaETojoSYjSmJzz05Wf/P+1GfHePoc
pOp0gpZP4eqKoZ5lF4xvcmrYUEYvkkQlRHC1ebanrYxqPEEVa2cHVIOAGHIchWnr
76YSZE15y3hl3DAbY2NMf0vlXztq7ASHyzdOBDZt31NcDjwppzXHFneu0hcbPbZG
H8jhxlqaIHUqUc3me/uEngISDcAnoi/VmZurP13Cd7Z1kYpz3ExaUmJJXoYaJ0Y/
QuP1LyD209nDGPx5aHusNfMqZFlF2G44KkaqfNfQO5BCL6YahfwgrUs4z0Mq4k+E
s6pbZIgIiLccokx0rmhEHJBZG5rO/8mfBIFM1yuvjAWH0Ooh48Hb+LTSTHcuPblS
uqoDtEdACbzi0znqLLkFGzBnN1JKdjMMQmqOVCLbNpf394FXksejZnnx8n4oDZVX
OA9uE8DcaxZMgYY6q4SZWcEpo28Zz4JYT8809Lz8xkpYik31HVNsPlzPowcaG94y
PigTq/CdbsNQGpXX9O8jbFYzF7y7B95Cai86wHuDozhQ4vdFhiU/3BvYD0MOGTGo
Ua/pSi9ZtoUQyFAqMU+JkDFIdUD/7ecG2Aj3exkEU/sAiw7QlWFdZBdgJVA9ICqz
cQdXhsZQtjHsNfQd5R8RULKcXfFuo1CAwEpP7rnvUulffdcq3Mf6x1Ez7YGVVGwx
oDSnNx68laEraJoT3tU+I0CEdRYNSAC8DZE9JMulwhbB+geSLQHddrakLXr5eDJR
DeKBoKyqYToPAk57L5ef7OxShgZnmeT5vpWjuJMbERYQzESoecGryX7lTqnFyJdF
AIi2Qf3JuFCOtEVX64Pgaz58c9txuBeDmTOvqrZEtlXVo5ZY6UbdWWqMePe2wce1
cTCTRyZz8ayA1C9egn3sAFnaz0TnQqK//aPvfmXH/4+OQ1W6GdQbcvwV7Hdav5Vd
oM2J1FQSyVAIznpgmaHbtBHrnk9onmdtebnuqnJHd4kNGCGKMN5nQmgtQD97s/8E
5GWM9zURRVxNH7mcLTHTw2lvIaT133c4F8HD+K+PDngV0uSilGsgYcZaWwCyScbU
KukDwQFF7mrSqsFrISx/hNuxkcMfMaFxXnTNNfwYvdl8xkgnk9XCtWxGkddwL8uH
qCEyjHpqeTyDUOTM9TjYbFCAMI40UJDTp1neLKIBKxu3P8VQSDLtFXNpAJAWI2a0
Wm8eGZ/QY8FX0YGbyvk/ZPRAgBQlWGN+sIYy8h1h4Hj4mAIpn5esdhKxXhKCIlRh
R+zKExIXuDhiR0H2zRuGiSWt6oUXgwgWcxkMlUaMz6A99I7yjSY5ucVFhXEwjpRe
UuUI253J3FgkFDcsZjaWnEN6Idtry8iJ3HBkBUNZeyp5KvH214f6iDTNAsAerBTG
QzcmmLHTXRdkrr4WV/0zAuvZZXm2B4M9vSw6G1q5zYzSerPqQNr4gOiJty2GyjDh
ctJ/LhC/CZwkKHgpXewmchcLmYIF5PkCcdR9U81ikqnUVwDgPoTyuWLwq9lhSmR1
Zd6fp4t+vzLfIblfa/3K0sJ8YTTqGPQZ3LghwBQ1jyhdSUeHmG5l00EJNvTh70oh
Yku4zBWAkSOsL2puosvfjR45Q9HqvAn3DAzymuIYD+rkfdR0nZC3mEi8JmE87vhU
gvzxafZ0Kdyf+E/cyl6R8bn74xGdGrPZgJuVwYOP54pvBHbBgehLxQmJjzmEeW/z
3sQtqTtIMxhNZX+JuIoiim+KAVlmMYxz+dt6bE8QerxVWqBYhFBX2/f9FDU5e0Fk
/UxCx15b/1DRL0enGZ6TxQxCZgn4zH96xDC0vkWNG9FrSBUERMT/b2NGH7Q3ORC4
B6sjhpv/Nzr+f26gAP0OoZ8TEb1gikZlf0Ya9DflZjzSoLZO29U2+ARNZdl/JLP7
GDvE5rVQi4qWh7jYhifvla50gJzqrPeWgQBjgjysNdIM5QaTYUiWpQqmEN0Vac0I
5yue3RL4mCPicxMHfehF00KxDXTV+maebRksdwK6ymY0Te7p0xXallqNnUR10vSD
hdrmFlPmai8d1Hjj/fm4clPzJgif4fsaLX1SY8HCGdogKKfagzM7JNy32iLZ5lPn
6E5ICbvMlKgCIWEc5KCRbmTXwJyCllAZQDy8eIDFbjaAz8nEYBk3zuZ1QFnfnmYI
RCmo+LhQ7o4+M27pDmkHOqDjnl2LUuMU22A1P7m4aX3lK4MiwqTWvma5OmAC+2c0
re4CxvPagwDggOi1M6RFIjIUOP6iBp6Wo6RSWXVgf17WSHy7XcME2vrDwXhg8ZVi
wmWJ3mRtTJ40UyHRAeNVmlH0rOYkO6cN/y+tNQPTGIRhvQvVt23yTNdO8Aety815
jD//CZh6DO8ifW2d+HNUVbZwJSHpVbMSYfD61ZUtBgIphMn78qDVb7wLUEWqWpzj
6vcAqrsuVX+NSidak2i9oRNu2GkeJxFAI/4jgfcXtqQ9RQpAxZ/GTUQKpx4i0Vmw
3trwIzBQKDDM5xRPNSMyjeSyEQeh1aJYOnCCwiz4ZjOHgxzp8qwXpDsiL6zSYELu
m/it1vQ19TnxnliU8PpfFTFSebTj4bKmRqK04tjjtQsHH20mY0XIt7t5Ty68RgIr
ZRPgR6FwOj1+Q5C5imUY3vv+1HLt4m3/4doUkI2jPuaSUb1IzIcE7Ka5mabR6hq0
AzBeJDvmgCCgkdJOHkoVlJXyXYxyBh/LanCxh4psH6RAqJzhLviJhebdFCbZ++m8
mEOVyUPc11pHWLXsGNYylOy/24ieo4jgVWTq0Io5viAEfr+EBv9p7QuDNMCrL/JV
DC+sVHm50ZQvnn7bx8D7PpV1CpzWqk4oYmZBtv+mtzIKVqPnxIeurMuRdfzonOvs
KRXTXIsHVL3UIx9mWrvVdz84PyUvtfdsRWbbpVCi/JQQL1Sw2sfACkqGZvjiT4iO
hvFDPBJRIkUYCQV69kgufJktk1q3fGgH84msgDyZFhHF+jsQzgrfJI809KwCkoSd
IXOwgsdbbPNfj3hFXHDYRsMrZxwsoVGyxLQzKk+xhq+pUJ98EAfnFHY5TM484/CP
+uuv+6bp0K5d2HnPsHHvbHYvYumKl74MBcsm2BtbiSg4H7Dxi7dLnfKSfnOgYOkx
IEsd3jzrfj1bTAwl4J8sUko97JP4w3uJjSZUV9wQ7QwCRRFrHqGvkNsTYkVaWun5
PjIjq2x2aJ/9Qiktjj7I9ZUT43KHHYd1/dbvYjH7R4hF4I6SxYTvUjCoumrihV6K
EhHAx9MTwwE6CYTS/1cdrFBrQ06QZl0VhrtVgX5T8to3DFXrROxwUCIt0/XB0os5
ORV0SS5juNHXOJZnkh2ogCAFqMQimF2g8Ea1FSF32nE0F2CYqJAJfogJU6+rRYHH
P0V156i4ARkGM8VEoQlMvtPnUylJE1haDkVar5uMMYNDzRdSktyaiADB1D+Abtx0
fXj46EotVoizHvK+Aqi/3c5zDFEbbFrvdDbK3IfbY8d8GtT2aUJENCAH0Jzkz2lU
+8doUtFLmYXOhLdVBbHKy/CCel3XMdxVfRzl+Lty/z0QkVZd2qHVPk/w8H6NyC3Y
AZ2LagkceRLxjV5xCQ8ECdys4OLHzNqGqgRWYu/AcLhHpZJhobYqn+sEGSMJWe7U
cG37WeYp9Xj2E1sDHekKQlyAlxeui8YYuEKa0NlX++qj0PAycYvMiDtM6paE8pSY
CDl+o90H8j06zVsBpNpRJy0AvhD/IMmv1azdvNdM7kViTQrrinKM2fvQGJNP7D8+
9/RkfFSR6D9yWEKpZ8RHw/g1MR/tkV0PE5Vosc8iH6clfWD8WjiY1mXLzxUSjoBO
eiT3Kbmt7vdkcrRZK701Vz6nsGWukgoAeDlRFPDLr2VOpUoPVlKFgBMO6i1lVWPt
vqiOcR91QRutpHv1n+cVbKVwTdiS8FRJ/WK98FObSvoGuCWPH6Dcp1l0i5TwqQAB
VvH8oxrGCP1El+f+2F2qVhuQlDo+LUDYibrKFKg1HqKUTv8QZjsd/FLvvHyFgYOB
OBiV0qHm7xwYhYanrNUo9d9B6FIaQzblrbQOd6st8ok+WAJDvjbAis2JbT7K+nET
+ZiY4SXbEByf3e6QWtJs57vg5Z8gT+Av7nWIDIP7cUmtNPHSqEqvS3reVnPPilSi
gSFHieRWzsOJv2m/gTEcXXVvKgBsXzjSgGYCIrNWYNkmAgFjz/KmTYuwHWGWHwBO
qz1+FE6fEvMNM82l/mP4OtyJN9B3qePe1aZiskjRPE6pvQy74EHgbL8CphJCCb7F
+oYw3EapwCcD3KCE4FOCD5IRiKpWAvR/o3DiHdRHG/nsTdrqA2Xn6vQlSphxkzdd
DIk7XExVQh/gusuHois5kkXwiRv/hgMDEJjekiM3GQ7JpomgQD5mRUOImwY0gIQ1
iWJyamnYc7wYJOIYKSGN8HheQMcKHomn3nenP9jXr7LBr8pOEEnGFVFCYWwxDXVp
APo8FGX6ZFj6WX97COsczyXOsq50A64M1J1eRkxgTDWlbVy0DMy2dzXpY6yId8Lh
XEhGXcARUvr5KVGq+c8kONUFxQBdmF0n5nF6LbGNEPJV4M49SOen10AJuarX6vZG
EqCUBNFUlBKh8Gg0ADMgL48HII9RRQQbaP2VhSKI9w0Y3Ir5qpELvFMqyRM84iJy
Hu6LbEpFaVpBmKrOkykFRjJEdZOItVUXXPp9fOlpjK9XChguraKQ2dWWJo7n8FJR
xWGRk1tGz32yqIMskoGLsOl85Q0C33IL+W/JFcEi7j0sO6NN4d2liVhgpDybgnfw
sxSE3bmdNzAqBI4rDT0LfLvX6A5POWKCHaY544jOROM4szUNxFU3xFFMqklfW0Av
Onvwv/KZI//beu0SPnCqbLlmuAm+vn7mqpIpGP9j4aeisHZRdH+t0ymGTX/rRP6B
3ygdhD7tdjKQ905NgRsKvz6USqurw8ew2u79qWMebLbTacvcXPjAh8rs/gON4X2J
bnJ1gDjqoSq279cUiC/NvWi2W3Ph8HOoARp8ucv0OyLH09oNN3aWbHx23UyH25u7
HWOm/jg2LA5p7rb/KQONv6VRMzW01P+7NjuDX6E5IdgjAWpDtbvhR26qUbM8uOjM
8+YcYJrlupwrZsOPE2QdOFVGEJBzeyUoP+0xIXQ5vB7/KL8f6nttlMy1XvLrrr7I
rw0SccH7JIMvFk7qFfd90thTl+39nSIt31WTuMJIyB0sAwK0nGfEX/NgcT70XXDd
jyIhOp7KQlORPTaC/GH8rKomHPF4XyfoyGeARNCNncWI0CC8NLm+ooyaDcH8T88m
9gau5MyAW6TPgMqbOodO2++e2n4oBrB8zNNeZjyeSIm/B/GaapBVHJpC0YEdUKkc
KTefBTE8LBlBk1c1fiiCX4z66qOIrXfGMEBTUgv4Wr2rI26dUz2QTcgKXWXDgoM3
V+ScChbF/rTIQ/w6CXxxfUa61ywlNmKByZ8I6EWu06m7BOYJvxrmEJ+z6rCg7B+D
e7IhU2tw7eyuFWB/NY0D38IGAu9ezWFjQOaA9hVgkXw03K4dsI9n05Dc1uHCPiRZ
URfOUZyNdBJiF+dc1kC6SM8NW0ZFl9keLXHmSXkeMvs/pfcuoCmq3Wu+puk3KSgo
IIK+KSVLZvl+9mot5N2NIadCVQ10JJS7XSswOGYnYT0+2UHOgZzbO0CFdeTqqPeF
omLn1aUtq+QU3iH2bgXWwfzTsLpzmbxu4Pk3IPCVNb/rGPT0WvUzyQoekQZhq1ae
+chcw2FoJNeE4K3P5bq/uhrQqHCgCUmydJMQOW1vUczTFLmTRb90Xc2dHGqrJRW1
htOWS46GrZf68JQIe90mkHdelA0ezycScTZL1d44uNSYXD6nOo/0+YKoneyHBNrC
Y/Aj5HfvpN0GC9GbvqHCwZ9/W4ormsy4QJQifR4o8hdMpCWa1stXPa02sVR15rLI
G6Fnf7A35cgCJ6HyHFvkkzLH29jMd+aJ6Etsqii4F9edyeeXQFVt40iJHy/tFb4r
zHGuPa3i2sMwcAsycpojQaWp6KolVm2VgeFObXo0N7prXQ2Z1s4Aj7CWnVmJzs6F
uaZWLN+6Phrys90mcUfJz0vQBTs5xie7LTa9Dck3PmTaen/F7ufQKvk+vYOG/8dC
0p1HD78ZkcLaH3QrnEnCc2yy4v1aP8+N/L3E5ds+4XITE6gl06waxlpxC10B8YoK
JQzBoTyjzSqAzLJif6yZFqU4xSZuwDfbqOhKSbvf40NJrco4d98Wng3Wmboe3ags
nxomdymV4XY5wC9UeUJHD6ZSXQcPMa/QRDZkVDFDeNy/0WM0wzGHHYuaSdkM3cV7
orHazawIEm7OYEW9b7gf2zG6beL7z4bBC3R4lq6CPundkFZ8myPyPK7cNz0GGPVd
TJ5xd3pNV3iSv2r/LC2X0ILzJD1IhRZK9pO9myxBAB/gukqCHRKn6Sp0KHnzLEQV
RhcjV9TnC+iB9llvyD6gSSJCQD7SvK9zKR3C9T0KcgQzyls5xX35V2RHICpzApOp
CAVbGbhxfY49LRPYA61264Ruf7F0A3PS7kHtCO2TWRlQj7KBN71W1d0tjJt7rsk9
x9ckH49TUm1KYBHnUd+EjDTKTmFV4pZTtVqrz57roqAeTXE6R2XccGxHaGoF+WCl
CTh9GXFdNUtzAsZxuZKdpDTb//BKtLv8QoY6Iu1QpBLO/3CcoCUk0hREzNZ7Vsqg
3JJvM6JEIve1Cffe7Jr3QtoWRF2HO/W1qHpCcYW13K1XTvrBl5aFm1a1c3FbIz2Q
77LX/1i9ddwWJr5h+1q0Bpz9vZuMZqpgX4CvX6AcHkB8JB5VqnW4fo5wZVD7Bx2R
2j6iqszbPSreTdowaH423hjDizuvGM2KEUd2Eict//0ihEwjhG2adxWS+u7mavmL
bjBITCXtqfVvoYp6D0XWZgyBv5pfOIgajAWBZ4z6XSsItrFXL0Kmik5eFtNilRAQ
g4Nm5tAQ3v8nJMaFTXrJJmFYfZ+HJALMsRjJZxuqhAq/rSxLgIlMOHRov0wRkuAP
ivq2SIyh9QkFN0hu49w6JygfRv7zYKIBe48yiI/OvloThRrZdfPG0GCobl9Wg5tP
krCv8gnHhW+Jiu3KL5FxQDR/EBtGzKfet542gG4zMiiScg/VosJgOt3caKkptz18
vi6MTmtaMmXGxkh/IC6w0XHUGdS86Gm4FUapSfcIYj4k3BGa5Idu9aMvxnjCtmPq
itvUo3JDM1xPJx4rdcyI1GbqU5Gw8o44QM3+CEHPqCOESEYtVTGuzyuQzt98ALSc
50LKN7tRMCzKOHjs5tf55Xnyi9Nj9yNEF1N1RR98AtD57hJxRD/brK8TkpSyleSm
yjCujPxNVdxVgNyNnbZYkT5iCjJnYWfG+ug0NHQaiRtFrHjQyzB1MFhupe7k58dH
CDmH3b3mWcrsDlgZBabATO3ddMc13z7Yj9Y4rd2BK7fjGklCl2qYQ5j1pNzGxKyg
fag5YgVmQTkR2aR38PNGhYclpLcPhChqmvB3YzUNAx+eAp0wns4qGVCC5w075DDQ
TSeWuCvI0M/wQkdALYjnQKmv0UtYp0zE3hHcQP6Nu9698IK/1w3GuFhJwwi6SVGU
nnZXeXnH8lNNsSx2mItEjHdn6m1OvqzT20R8mIQn5PkG7NdIQQaJXdBA4+Gld9K/
t1SP0FnveGIkgobmD1plDKOrh1cB1nVY7Kpou95zC7WyEnn1jxDeqDDFNfYhdVca
xMU8GZfz1Hq2GFrY7wEx4D/3sWkt2jIkZw8SykXQz6HMQZ8UwLIF7lr0J6EtUBwq
hOnU+espG7+FNjoemIM8Vsxe5UMntkc4gfD/+ciGENkbGYRDu2eSqK5tkflknrTG
NH4xDplZ3ohUG0RME5TxiebXYDNVzE+GfnaMEyOrUE/LV7c0MHVvqddMsZTOe3KV
+eugsm5MWZkiV4XDeLMheTpRsj0ZgisDCysdSVmjJJZhKvV00R/NxiJQBTZWp7vB
5SeA1BJ2e0rcXhHzmZ3ypv9J6w+Xyli3agvSmCZTHt5/RWS6if2odYu5V/tktVoU
8/g5leJ2f8BB8xdV7opUpeReP24CngfepNnQvGLyqdAM3UDGlusjdkpTUOKLnx94
5TDP0Xjng3I7CoeIgRj0u/XWHfl9VqJ+iCQDQTpsWXED7tericYaIj8am23TMFXX
QYrUQWP2KqS6Heeojxg47/ZJjnYZeqOkrsvly0Hgd5g1Teen/r+FnsEFxMZrQ9mQ
zF12uKe1vGHNRi8fgukIXdeigukJIKbwXs88uRasUxrDkQg6cxik7giUZAWZ6azr
VHRH/BlxV68yQd/RTRvZmGdtplTYqJu2bV+0tAqC16Luwj4VKCXdDLUnK6M1+SKI
xQ3R3/23O47+GuFfWkhg4+F9mBOBXv7iwy6DAQF2TdCbOZMZRsFtvGZH/7ri89Ct
+CixPn3RluLVXJZDVr11/nXkdw83rCKjhRZVSytDtn7444lFV165xjD62nVwwO0/
YNTHZuIxm82RFr4pagMesVBMprqAYJBiM4CiLFF5dvScyb5SJt2eTQh7DBDacb4s
EEWlVopwi8Rj659gkxnBHbITRmtv3SJjscxTd96iNHuruWzNF+pw0ybmQ+LwPdm5
ctt9w6MQGYN14QtPtaFV3cTf2APagLCIWUAwX1IK/HY6g6nbVxTxwkR1xXfrNNYo
8LsqpuZ9mzuFLdjezm58T994iXfw2FN5GIfTXdBEvGhziWW3SBBixRrZEIj4Awct
TCggewEF+VBO91Z3x0V80YkubMTARCebHXtDqFMcUXknS9MQzh+3B3lLbU+pisgH
RFu8bOk7TGphxJT7TwiBO43+MSxCjRvde2RUK5icTR7sT8EOenKO6QGGKPNT7LXw
G9C3BN7fpfa5u0qxR2g/SBp75B0YBLKatXd6Fo0zYqnXTATrBsrkyv6N2QaPWHqd
9uI0ad5rppt4QTP2nmtWFbRhorWng4U6/2r+2gl16bkM1XcLadJ+JRmeT9ueheiL
90S5vOfNDCRv8BDqdSqlBRFIfIGzVuXsk3N0iPzNDW2+HiRxlS9RnucMS64IzhL7
0U2PM8aGnBjaMpfx/OMGc6Ng78yXpKI2z4B7AYue6RdWjJ56GGS8BK4VlA+h7V/f
AFhkdvVMWI2/X8qsrNRTjHh3iixAgXNTpPLZV7KIpWTYM8XCnm4DUcwjNBO7YlLV
PgELmJVzHUngKgggRvz0PTaDp/6visX3j6kN4a0Q4zE/Vi3XleHRiRhRG3dHcW5F
b60JHyuL5K7GMtOvNayiwVPUDCvzweCCUJ2ny4Et3JKDc3Tt34mu1VM0iIoyyoGG
kQ9nSEW9u1J7Nw8GjmHF/v4XnWIKqcNCt0fuH03QBgqA2yUCYFDPPVtBMj3BhNdd
VIr0gCYr9xqQLUGFtKlyijedzLUbSUnOCAiyTaP3Q6PvAa8xZgSfnGwz+jLrb1Bo
oNv3mnMcqntK+uMPa2nyMZY7mpqaQaaHgDnWxOVfwAxsUu1Oak4O/oqwh2QC4BfG
DG4UzDqcWvArl5DC7rSNG8gTjDnv5T9to0Fxgbimwd+VS/6trJgZ1arfYsCXiNsi
XTxR0AS4dK3sjjcs134bnXjjT8w6xYK3EVancFaRK5Q8v4AuGjrp/vIhFfcl4rup
Rp0z8gEPMyCJ0obh3EuKBzj6ZkQILt2autt8HMq86rOfOQm+9kHdobwIonpj1blW
KAMPx7coq3raLV9aEK9DIinT/0LmsclZ7L7RSm0wBgClGJ+0m0DJCdFCyLWIlAtf
a1yLA5gUQ7PbJ7laztmIr+3jfan8ulw9fmIFbOnrLszzceTcgd0QaFbdNZrYowlj
hZ96iXRFLs/7oeuC88+C1WbRiAo1DxteOc3dOb5OENI0C3EE7sfCoJjEdRVwUkAU
SkgoRCVIyVY7O4uoJ5YGG3mrbmglQ+fhYK5mAFdxdi/R/5XKWwpTc+K0rgYXjqQQ
Dhra5kASwsfORfJH3/3If6M0qaiuyXKoSDLeuban7gUv03N3UnOM7MVWxkOxYDkW
ivL+nyNriOEqb7kZm10cMEtoZg7dXOFm4W2eWAKLf5uDIOn2AdJ0QwWuIjwQ/L67
9QJukSUTMEGyRPpT+ChGk7LYrJdZEvNSHgfs0TsCKNOMx1kNG2UInEh4y6jrIFpi
udZ0Lfl3WQ/sCmnhqb8L6Q5vuSKp+u2aekIIEJtVgeERuM38dBaH2wYDFOe4B7sD
hwJe8mRe1bCOhZD1ldjTd60pjvJHwMiuONLJp9+qyE+N7uqKqUnLHzxJ83t7Har9
Ep6yuSe0TQmdJ3qfVvy1WiklsNkiGO9w1jehhq3fxB0CmbpXqa/ttlDXnzfh9wrv
TQ2/k9Qd+EnSaraC4vp/+uWW2WivYy9ob4v/xQrNg8b0vg3rocPzxwL4zLeQCKIX
DJUP4UQ98Y0vE0A4zKEmOHrN4LasvEyvJTMZe+AWOwSnhmzRqskLvpegk1ZHJtUo
Nfcc3A3mPoUVsMFcZ/bFOyPWhk/J3wBEItImvYIUx1BlqdewGgAT9KZgdi54wNDR
AKgkut9q+A/h4DmVcTP4MjANkSQTT+nQI1/S76jjMtLjz9Fh4bkCmTAm/dspyRNv
vGgldlUqp6okBQEBjzbkt2l/dRrA82iIYXx+Jr6PZZlQ3RjCOK8Rik3rJMBsAVoA
qOpXLUqnK15kHX6KOTgx43o79gND6wco1q8um6Uk8ANVXKxfP7imKtLEILycCxZe
VKEfllzbkBg5/KJRNU10Fgr2xIhwDo6k+N1X4uNe1GYlqMzPVtXrzWYoSIHYVAbT
6qLv/U+h9VwvpQjZUhRUEqxyu902o6c5Mk5TvX9O8BXLvPI0FlZWfgV0JhSqcqqb
aIV1LjzcnZeBnuN6AprfIS1V7+khqXmz9Yhb4VCx/WTlg9qbXKhrWvCAttyT1Jdn
xuVUJoQZeCJ/VrxIr+jbX/v3mqhAjX4o04uXxRwXFGvNWEXktdyro6Txi7kmYj75
pAkleLuxWzQg/gfkOJ1nf4WvDB0j7EcPT8L6adbTWuOkO6T9ThrmQq+u/umCDZa9
16n21g2es7unWwk1MwLh4485+no+p2TrzapXsVnl6e/RDVYTBoc8KEZN+MMLP5yt
gpPvUJ+MI2sZ9dK0OJ9H5jtkwbd+0QoMlTqcs+4omhhaTzP7G9u+BY+UhJWVfCLF
c0S3pWQqiwxs8jC5veeTvPsJeL7LetyA/1I1JcRW/5SeqPazi1m1xG5M0kd50uWx
Mda+CYQ/oS4pF2k+UHcQAEnwrgAkuKw8M50iikMtojjHx7/YBuvEBRFbNm8ri/AN
+tUYYls15lJ6ccumApD2deE33uqAAjYSsTeCrdjkm0ZxR6vN2o7/5XP/Qc8zPIHI
OCLKzKlEtAJ34tBfPD3vLcH14Arv1gjWIrN54MgzhoOqaOX8wpI1/z6X6dYMof5v
ZQWUQ2Vwh5HyEQ/44LB4kUK7UgvWCemUT9iv94ywiUfRYNqObZxeBD77JM91ExW2
QG0M51L8OJ2qr1+ojjZUIDOjgwZJLyH2LlUVj5PZkbyZGXqepXq4/YJiJf5FJ+f/
VL5GwwupgOeL1fScwyn/1LPUdaAPrtIB6USyAPGNGHKrc5/j1IHSHA0KPmjE+JA8
pOFkdNAPfxyOO0AgYB2VXmSWYjTr8G+piuirfwdx0i2s65BuRTsrC8T0OiKvgh0z
C8PxEHQ6c5YECzTQfit08qO5ZOyUjvr/aWCW6OlopoC0fCekEClj1ebwPxLfUFiJ
GfSTeQQVYMGWTVXNvK8cDLot5pxwg6MVpmIQB1P48CnjN5gR3tq/GqQi7DnjJ2vG
rxdPipIPfv4H5I8/agixxEzg+fWlatyNJ/R+EKuvkI3G0/lM3uMNYtrqnc8SmLW9
fckj9zPYgAxrR15jMH6NuSMwh0+Nugtc7UcVsnEMwP0JxcwIDZi4b4O6Q7ZNMK3B
1NSFLGnfOaWxWMxXkZXhmNdvFaIbuE+Rp6L2KguGjemwSmGhnTN/rlwmzP3hH6uH
8QZzwm45ajNeJTXsR4b68uIhssOT2qFUQvZ3GDrYICfcsMzOWm6GmfQSz5cmjFqO
QoCWO74wKAakttgTehWbiavSzhHHkdRPnT4eW4c91sMHR/DcZ4Qg8cuPo7cSZ7Ck
VPF1FLxGXnuuAQZETA6h/LcrM+xd+moCQR5b+cFjc66cT/t/JWI6PUijhmISbWyJ
60v2dOb+QaX94WHBUkGdNhjZoPhvRyjQbW7sbQuVRgdD9wg0kLiwXB4yWNm9hHlf
/9RYossX7dP7eS9U7dhmTZQORnarEDcqd3PvhYvgZDvKLUQMXQQCIgh1hn5075kA
w555ZMzSApnO/x6XvY+aetrG1rh+/bsnl0/fbsRcU3J2YsUa1wfv4d3oOHux0bD+
HrhcVG7cWBp4Dg1ikwdupSI/lYnwL+ES+IJxUdVNn2Oo0oJTiUBVbXJm4HTK9ggs
+ti0BIa0X+E06AaWGOjVnakP/7y2jYDhWloMX8OPeCNSbHIJEV5G/4BP34czPk3L
I0PqDjfth9tIxlzwSTpcrolR85SnzUBOVmtGiDdHuhZXPVQC9iPB0crQN5yHI1rz
yHmKslFaYpx50MXcfThj/wKDw1LWmfAIFd+7+mD2/YHtZ0Y0zv0Rc/qrSir+Bylb
0dsV9/tuocmIF9hRhiXZVCwZqaQtO0bBhXnHBGZRkQ0AVNVC2skN+FjOIpU9CGvd
QEECaD2+gkx9cUfvmOVWF8ErsgNYoy60jizd4GEg7+LUdRXjCPwBAk6D90k8mhjO
gPqqtIke6/SdyR/fIXESbmffxFvoqRk1UvJhh1T2XhqLoF4jWx3zZJg//j0eDLYu
+mKRTaXrcd2MObonHp2LaoYhB93ZByeoYDwdJAGsyPthScDv7+oqF1jWbeasFlb0
81/aeG1br7AnRTcgt5XinAU1PZGNGrlrYceh00GTiMZeZeCRBJl/jLkNxC2iRthd
/bIoqdRBtl0Lk6yRMxKQNwYaaTE3NhMLh5snZA9XWP6+p8yMduNubUhhL/5J6mYa
fhbvD8k/Z/LN1O8WV6MVkoVA3Um9DLmN8jyexb3VTNQ1punwVV+fkkSMHAXRFurW
+8219FVj96YqdGwzYyRMmRs2CX12oO/eQbYLa1Lu6S1D4w1iyBqzlWqkD4OwK03m
Nfa7VW1mumaOAk1V3zBvE45epsJoTUofVQkcoW7Evw8tpzT3FEtO+vc2OVLVcutw
yxi0xdJHZF+5UnqiMSNpYpuNX4GAAejzm07ZvNLdwLUweqbWExJBZt9hLdFR3Ss5
Q24xrQZ2EGCuPIR6B/08+VJxtv8fgzh0UfxoM448gj+5fdybA4SMMmXJ5tfw2Zsi
3WvIph3+Wf6F2UDzQw3nCq5HY7WEL+xe40BLKnU+4r1wvmPQwU43WzQiHI3fDxE1
jfQPBaLqKEEewCAkJeHUP009JZUFYYCy7lL2z7Mi+ShRGwhElzbPQAldfE1Y2R9a
olkJnVEEXrWGd/NnaFULMh8Oa/I3uHglCFWkIzL6oo3sRP/sey7FfofLNXwuBceM
J3U+zi8P1o8toUOhJEjO0Os57f7iomV6+yJ9SSjuub/P5ociBTl52KW1qs2E3DCV
SaE0BmjNBTXAIEy8a6qV8EqzesjDGjKdCokXyfgYxsC07zigtb2C2SHBZHO0JwxF
4PBm/U3A6oHWsKhAdI2cPDbUW9O/PzQJ2YXBxmTOKBEVe+Xhw5VF2Tin+MUUX9Xy
Ud52rrJZa9leSqPgxFwXOYsfI5CdBPdbO48WHMYHVkWryrcqpuyzsQBRVONMGklG
RGwQ80Jsgj3SP0Pfu+QBxmHdlRqLJP7cE/BA6cUWkwqQAFAymu59YhYZNwMkZTom
jWnl0a+LAjiRZBhL8wiN+GjNHzyyIYVyYXGQUQSfPC9zQV2sxdd6PkdP4baBMQtR
7z0MBhkzbNBMRLYwcgWUAf6fv7sEX/xRGZbaq4Mn/gxDAGOwrE444P192EPNDqAo
xP8Fk1MAo9DnaAl/xmf/wM8vBy86BdyMGyaXCWPmp1ZtN2H1EKVv4XrTW1d4DXCS
oKqhVdsNu+3O9tbUD9Q3so/yrYetJs288sYWgplFWB+goLE5/DHZDmKm7yzojORO
CEBZ65ckwmIsMoQ5rOdoDvHYiBJuSyMg0+/h6K/u5hBU/8FTdbMCSlh2lfTxjF5n
kY1ZcgGxJujxhz4+Etwb4no0vg2fOaYe8W0Obb9Lv3NdIAJrra/TgU0XcXgXheJB
vgQlI6483kowyrNyW7MMDsdG8QGYFV4PqhoueNM5FYesW8lM4CT5eHgcQQWYFaVG
9iF/xOnTEvm9C+QeFPiPkJSR84ODIlHO6oNhq6qVGJsS/AET9O//CVjguWCkxowx
tYRG9Ab7LAxMKyqyBXjQHLdgkpdij/5kV8bnUOMlk+z5QOOL+zyRDLVnWK8HPy1F
hFU5w7nL0+2mSpZIvhi567++N3wMnQ/y8WcImByMbwMH1ZrPg0TzF64+CfS9j07a
Be3vU8P2bdXBj700SHmoBeb5Cln+xNV2TxpncIFH651s57b3/cE05yCpzhCfTIBS
23k7FMID0/yhAHxN6QzibholMCRy0Wkq5G0v/lJxdcOUUGjn0hd9w4Vk83sOflo2
oA8xhiPm2OhcRAvP+RvwAqhmhOTEIwjPKNlHin28uYMXhUQlmZrsnkw/LDtPwr1B
09ln9xyvcKQwMoQdxzbMFzDYOSDd9ZIYCihUMr71FkZH1C9fRkMQgh1qisgOrKS4
1C2ftXfbAxLku6ub/dEVWqgY+jA6TeG/1DlonQUSWLpBCtDKCaOBspXVZA5L2WDT
0OruuLtWOIejhrTitg+JPPc/Fo/SKCHTK20rq7IipPM4fpfnRFrCcm5TP7SWYS64
ERrnIMlPLQMQy/rryG1a+iOFddzDQGrNOkmolnH3eLF+7MzcXteiqzHv5YvfvRlm
m7UPkWXnQNiZVX2+q8UXT/km6lEuCJ46u4D2UB22U6biL7FRH0gsCRUC+N383COQ
9hDt8FmVSd73WHnR2Cso/0ocYgwKzsKLfw1J3VpBVuUx9OmNKl4/4YqYhmHtLsGF
R4WxnReg+PlGrGlbqSSfMhCHzz1o53hcYn8T3/DQgSpeDdBNKHs4JElKOXN6ZHUt
8yh9lm8xtizYhP1FDBeZV5YAoExpprvRb7ZyqDsKdefdWg8lF+FOsw9iC3Vao77L
mcQ/TuZttmm/dCgoaPiWv3x7hcrlZSQ/grPhHNxo2OV1kUHD4XfnOVYdfkav2qq8
TpTHhH8Qa6zBL9oU5PPbBkTsAWX9qdOc/iz2GRO5WxMcoSdI90ThgYRwVx6099KJ
a3IZ3NbEfmII5tN1cYMftYPLKsTQM9koRvTIC302Sungv3RpcM3k8AamBpHWk9MU
MDcLaGznyYjjTbXYnaogrqaQy530bW5T4+7gpD2BbDuriJcLHr6DRkn8L5SAp4f8
vs3s4Y/iZskLZOqG20P3Kub/eyX0fZYgTESmSKutWqliAn8HTuVscuToEaQtC9s9
Kac1xq8yu2m8VWyhZ0DRRBA824SxNsZirm8ZsRDQJ3BHMmXVHQTbSZ+pIwpZcuOU
UWrwAxK0Y66Nc8eN06fa5Qu24sm1FW2mi6bdCpDGIgZg1a3tzDx877BCK9ITM13F
yrqf4VPZv1wrmB+0U32W8U1L7njhUaSiRWV+7ybPfOfm9yQ9e9wA566k268KkELL
w5oTMFAKAevWbS7kfQKvuk4jWB+jCM+ZaDA0dJ6xEK0kNPrT2Mx5SMbPKR34cSJZ
9HyH5HHgcSKOdHn0HqZvEG98EeCtN30ffYhuziR2sZdc/slq8bAKPpknKVYyv/nO
0jPIG/HQ8yn8fdMHxOwgsdyCt3b9scRNLgNKE4Tk3GaB4GKpZ3H8SaHqsD1cxcFV
ShUFsmQy2nndvo4mUq4Q0DPGnMiVqO+z5vV25groUzk7hT53XHdRqHpTvWOVX0Q8
g4xYWHraeYHDdj2FSP/sw6kNm6SMptTO4pZSMLfLJ8t6IwXNc2qwad6YmCGPCWrT
QjdOzJQ7dOuhe+OVkdKqFaF+3dxDnorm8br9MmovbfTtvD6RFyI1/V8rA09s34Gz
iUZg/f7rCJMMWwI0QrakoN1x6NMoJ5TdRdSFN9cwia71kMdz2JX6OrOXitL6R3jk
b3SgVi1Z/RpAQazKpfZKHpskrmlykWZjb3v7bcJ9PXMygVuiPOar5PXOagOS0epA
r/0Tw4rRvCAPYgkA3orAAm8owjOuPuAxgE5QL9TnRuKMH/mWUXrvdmnhwyQgboaM
Yw6xo+sGtDpccNjRI9Ma0j9KWFUtAbTFQog00ph56f8/rCPtsNBItlH8ofLESrju
yBtbq5KR0dgJKySNV0B/w2PutuciGdP+r1a4/fx+UfyR56SJiFZINbfqZYKvt0sw
Xs5ni8LW1dRtNzPeja2GGMm9jzPbd8YtIYAXF9y+I4vMISvNX1Uv8rjRr9z4eGND
5HneEoiM711c+OKWqI0Er793aKQ9Hb61SYLpQQXxysFIhuMBJhzSRaOYrr4SXNOS
4cb47r8grgSNLBfMcEEdic8JEsayMgyqaTMV5tjdGCn4XkOh+zqPcns89w67qJaT
jmxPp/Xw/34kXU+kviUS7GT4QwYehtvu5vxa1yq4olY0VKyza5uge7PFYGjpjeat
jetvmKGoY5rQAmw9UbARn+ZI9uyyCqWqsGh85EGc1eeV9TbXDVXUJtl767g/zdcL
YHtcrn7PSZG6/PjUHtEeW1ub1KE9VmzqWLeauxNmACxJ10tcEq1kaarrXQlxy8wf
RZe/tBN7RoZ0f+Ru7Pv+/+EwmYtxgvtxUNZ3tOoUBSyimqqGxhzzrbQDPNaZR9P9
7NRclfkURVGqaU/gfMtz3wF1CpUrI+jrkYbV2XzeMIhUKZlqnpVfuZ6jusk1BXwG
N/h+nr2XPh2SaWS+6eKlGLZho147HHZbh6wn9MsapKqQ2LKYmKoOib/Z1iMqD9va
Vga3nKs+qRoIb12rW1q/TsAvxaqcSVKcuEmvnnppiPDdStzziYJRmJcZab8FJjjK
rGWFIFMgvP8zxm7mxiN8GaiNZ3C7WtSEmt/oMeQBtAvEmuVxD0LBT1nRJ07pBWSz
e5Q69VQYFW84z1KV3Als9LlLbCUCGhM3FQjWOd914uIwefPjGa2LMBI4Nn1+6CTM
HmQDKc2hKVohHOcACVYfmlAHTPPlOXhyOwCWdgfVhJv1lXIciHJyEas814tNPKHf
1h3ZuEUr9TCvA0CzORm3n/mChpNDlClq2HpX3MYa6OogW7ciWcAXVv7DsW1bz+cH
fpWWRSIoqDh68EgpE9AaDBow2/Jd4AvY7tZ2l7IB//PV36aeVPhWuTINVZFrFeuO
PI+kR151CEyKRVkh6kpkxZxE30KqW+1xeNvGBrvl+GvkS/5KSgzf/b8O1qWdv5fv
uglt7I41+rICf9xzCzRUB6aYCGRY6w77lPwzFS0DcE/UhrNI8Ilx9vQVTk+gBgDE
vVzd7Uyf86mDW7OIa8xw/dBhyzopw+ZdkYTl0T1/iO7cZYJkF31mEOIYo2GYtWfQ
fYXxKZrJ/jRPkdRfBfE7UVO6s/elxtmT2Y+UrC1njRGaAI/K4G52AqtAdl+K7tKE
FcJ+vpHvErLomXt6Qtl4dD7kv/EwTNCxOz+AKFpjmdV0bbP2MMzMLBE4UeACTzO0
7Xd2j6+Kz153umZJw1qGDh7trWk5A/VNo4fLZ/JhexPrqSarVz9it1JG8U/OeHq0
AXgK/Z2MNIeNCLVySpyUtVpSWg76LvIKxEBqtOwNfjvaStqttdwqQjCSvl0S95+7
hyL5CvzqbvGsAWzYr3PNcC/RLtnCwHTLgeald8ZgOORHsnHnw6PI7AuYu1nn8Nk5
0ZSFEw76AuTxR3XzfqWYCDWDSebLlTohei2bWlfzy2fWoNi30J7+FOoANq2Ie2o7
cnyvQ54wcRa2Ro8alM1S0aeW5/j2UGhBwNuDmxyeegSdRoGHWXkNLez8IlqJEf79
RY1R/PaGptnfgrqJVAm9XaeD2YS0wK2JZrwz0QPsvJTl+rdYb2bUGwd+P8pET4dG
z4AEjzhv2xK9ASQ3PoRuypzk0iS0uhVoVlMIX9gB/GP+jl9RUKni0boRldV5dCL/
+jCsF2R0lho56YiMzGSKFWP4nCt+MuZMEDJOAeckGcVqR8sk4cY/7fx3claAJGLk
wM7RQdq45OkmJgMRFq5aTcJ1bp3n+SIes2ZVunmmOHjPeu3M9/Umsn5uDr+2EpnZ
d9TqmugE+GDB0L7kl0+OUMA2TiaqkXpcNmTDFZQaxN4B/Lh65kYvTMADL4Qzy4GV
BqM6mBE0WS8Dbm38vg9Zt3unH6dWKt92AubMyk8/eqb90an3ZQQRHOj3lKATO7Yb
obRGaeE/N3RHq5Grc2FLWomdFF4nCfCIPE/wKmqPcVpj+/m9PqhYjcYVukiU+jb1
I1DVHnor9jkeMbie2a6Oi6by3SiU5yK46eqv3YOJW2QSXqk6RbbdB+M075fOsjDq
tzSCLHPSJpzWaQKVcm08yLtyhi3E0bVspwmEY8DB5ebOBcsT0WbUt005V9RKJwgN
tHpL19jeLqMrqKbNtM/Ab7QT4Rh8ZT9efcMOgA3dwG9OewC6FyX8YIj673q/XxDJ
+gBEyTz7GRql4DB8qNsmkcIhJV/vaY6qF9K3yUURFyH7s8P4hpiJcVM/Mtg3rL/Y
cAzKnZDwsFUoh00ihgcV88dlS9xRZDIipj1V5tltUOUx1BnI350XSVWRJqcs7wVy
`protect END_PROTECTED
