`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qD8x3rVtBNWJ5oWGqvy6FrbFIh4YKhxeWr0ihUt1+hu3t/SMn/NtZrb0swnhGJ4e
niTjr+HhMObO0E8kFD7pWecIu6mhjttXANwwZZjKnskhHdqr2yHtjtvdvWAJJO1j
pyNuGK7pL5SE70lqqIUkgKi6H5vYmz/mXQK1XcWduHz0YumpNg2Ela0T/9aLY95T
RZhhdel2xcgAClTfF1pfNw+DcNnxuBCvEdcmpNmo4NE2YT35tCcFIq4xZIMCgR4K
qgxUo+bEHlIn7lYb5YIbBVo9z6PZYecHSkkx2V6sgpVF4lsAVj7aNmfMqdESi4G/
hPame5wWygZYe1VOgiUovlIE1CXkI1t3ZQmySUk/5Ng9Q79CjBiL4YccDiz541wW
gnrVg2AmB3kW10RULQUIVe1wVUkIB3us0qnZfRKLfN/quXAQ66N8v/NKGPVX5vDK
USS6/kpJyldLYnh6DHOQjbqnebwYJkS+TMa0oCX/Nj0/BBSTYofTmb1z9Puy7yLR
zREfeIlU/iTQOK+jakhTkHKOEuYdc9K0a+Ws7vtfDRRwMtTpBdutzleUdQpqkJeS
BKX/YCvxTrLHPIURTKuokcre9wb+wXAsqBAvy7aa/BUGxgfpS1+UCRFYwpowwjaO
8n2X3FxsZg4Sh9fvQKSjvdo19aw1Y5cm3cwe8vTkrRf/2C5oXBD/H78tQOwrgcNl
oYZg1T3ZmZh8Xu1SnPg6CekMGpdUAXrgvSporWXtIbszWkssvzEe8rWm5J5w827E
suqQ9xomLESwHvXWD1PZOXfI6kkbvdZiFqtrjv2iVEUEnA6KgqbgnR3wXli1ueR4
HCDTNXc5D9qkIyA/cPB9XmBFVStXfgr+/4VeS2zBFF/a7Jd3jdf7Sb3hoNqOh/yo
kIbiIhfbNBl7akFeWOXkdP+pNkVFVJluUlhdBm0z67dm8z64Fj6dQizia/jNEJIg
ybVYfNWsRyWFiHs38JqhGtIA/Um78Ivq81yBW2CPYp6x748u/AsHTovgRy4tpNwi
hiw6qIQVNrTvWQ2iTHPu2oau2+64moS0E/JnVwXqCVe4k/Pt5ShllIix+SOBjj+S
hCirxS+N47JGYS8OUi5IniAKdhllZeLzkyhrkkPoQAGJS0ohkWabg0QagQa+Ls21
NO9MxPkiuJPI4ULSAzydxml88QuSjUGSwIi5t1NtRHy6diwJWZ0cibcb6mbXCcGM
pGHG2zxd4rFukTGjuXcUw/1u3V0EBoIBzYqR2Pv/XGV3k0GJ2VV8VD7KG88Hhir4
NOc61ZbI8GhIJgho3JOi+kRLzP/rN/plULlDIuzpvA2S9Mr3oebwuvL88fNLPc2n
NYj5WDw07wybqUrubkVh3Yhy/QNSKCobBvCmzm4djX/dBbDFWgJmWEDJLJDWgk9T
yuXMQNbYcREuBmMQ8YVj4fQYsOD5BmMNy39SmE5jcdIH3IEwMhusiSxGd7hzKpq/
/HLLTr8l6tRSsd517Y6SODGWWd2r7aLYdqWfQD9vRrnGqfTiThFeU0OyKS7QbViI
abgVWLwZnZXOz8kMkDc9DhkoSMvpnUmLoB/8Gqjk9XeFrByfedVL0djzkKR/fyUa
XKcX9MDKVd6kPiCY5qpH5RoGudXAOVv8Oxe7InVOFnxZxgW6w8dmlTmoWcBLYpMu
+pUK2QlHtY3+Dqvy43u3UYqkjQMGc0p7eVX/e7qkBujabBQwJe0xyuj9zquDLbqA
Kv/6fnkglblvyJLJQ00qsJuq1vZZ2MpJlz9xjSQXijSW1f0DLLRvCUV6oPoiHvph
DIPfpG9esJK9AHVHdTU0zEwLg4Xd6eYr1LG8VxE1ExqDWe8ha4iXhTeDWgmg4515
9PXuwFbLRnRmiMjCMMDXgQo0hHyp2FZp3yUOvD/NX5HWPi9UPoyNYGQx5p4kmrT+
ioeomfr2HF0LFVmLBCjOkHrEL1qXNfGJwyAjEplRy5DrRxIzMaQOUKp2Ymm1V57n
VBsmyLiXcZsSoTGTLb3xWH/WfDg9C3qIbZfOa1qO+hFuCvCsHDrNlkHYfqZGEybC
6onZ+EGz1Dhbghj76pC94yEbsT5RZU8/WVPfmgHVV5uKr6cqdmicDbkIrjA1R/PE
ZmyqpCpebJv4hmz3+XfnXng2cvUhYMEEX3mGAuKGc+kPTAmPqw2wxQAGS0xV6/F7
+UxaNaYRtkg7k5a0h1TO0bbqDsZL0llCCaa8CUCFWdjpTUg64bPbF60PkhQ64/Kv
4SHNud4jxKa9lahHSdywARjUGqrzjx5wGYtHjsX+5v4qqLWB3A6mpf/W75kx5oIf
c/ZIZ1xngLOsoU7iOHg2WduHM9L13OzA15wvECK3f8dPERDPCtZAScKDnHk+iO3D
bIpwgEv7tXS4Kk0W6ShSVxD2eSBrK5fjnYTqvlpvt2hWM+iJfg3zC2wIFnN2tLv7
RurZexsV78RoNe0Rrs1O2kunpG/r8VsoAvDF0LqDYhhxdpVcvj9QbTbEPF0hPrZD
K8vFn3T2VHd77zlh3YQFNg65dodJVbW+Dhx8P3YmrwsvCjVWHvs3rF3XtAseVGgO
aT/w5MVMFy90YvW+7FmTwzqaPFOA+a194CHYp6CmnzA7RDv33sfQUqgkdVa5RMVs
MVF5ccY8u81MlIM0rCGu929XxIeB90xZpjbJYKWYiJkde+R3DmAenDi5fokS48vB
TwcsYHYyieDDF5c7X9zFjtdV9rEQc7BIbs61oODQQqvn6t8fQgLo3hSf9DzUBAUr
8IjCLWuuYTU/Tu+Dt3o0nDOa6EjVBgm+hdYpP6g4WfjwDPHzswOjo3URrJRHKhtw
jZ42xKBHyC54kUZP0ZKgPVWgB0eQIiYP2hoRebpDUaEWcELUKKskYtTk0rx0UFAy
eDG2SHUx1w+uP2pcY/dFoaAsI1CpNby4bW9dQi1958ZUwWybHlncp4Zx+hu2rU4f
1DzPBJbR9tl/HdyMLwzvcCpa1rq1MaUIFHcGqbwrh7dVb4KOMn5y9TpQ3arw+aVx
Co+1Hxo0S1AO25n3l7gYI58sykAx5VeeMf6XJxRUpA+CetXHkJeEqspeTFliokSJ
0X7UncrhZX1WkjM4WVsCP3ZDxV/CsrwbDhEAS+Vrg2JDdq4elEcFAjAKb4hza90a
qmBE+33g8AIoeof8Rt0e2zAUwgyHV9C6j6a7tMKZsPPVXBU062kG8qpcuIjRbU9X
DR5oO5rg3oQwRJu8xDvqu6po+zIoYlW12+SB1Mne4v/pHMq5ym1+mZP+3c49GaJV
yPMMmYCCkMKHRZtZruT7FE4wK7d8gJi/GkP7EXcdqE4zBwIrjp/QhIqawb/59SY5
7OhR3E0z2CfetawD3hZQITAW6AtZ9/jMSPMgxfo0eUuGJUFazm60/TIfJ/5EJoW9
E1y3RsVOdv36XXMgdQtKJQzdprsQyHuIJ2DCQF55/kHpr2fVqBKCSNTKjZW6DbPx
3DOzhr5UL5YEN0zV2TahEla/u3zwHYRWSJpFFKC8LFxeGxhO4g94MmucGx4N6s+4
pJI7zWqK60YvFgHuyjol08MLg5kK9v5+XYgqvyAnXvFFmaiTt7jS3kO9yMHgQsV/
ArC4YlZcvNY12aMGFfeNO7KdRIBERtqOPCBhR9m4Ms/MN4s3ap2hbiKsYLGfAl+u
U7K9EBq5L0AKzGw4I+j0hFN0/+dA72Zx/zx50CXhuAtdYZwIferqhgAgHpAh0HLz
xWuWhePe7rk6wTnzFpcoFyhZN4HpT53qBHuzM555Bf1F0on+cCkTL9fuRvsLqX08
3SY4ZdfjwOS1Sl+m59Uxwvny5yFgZ3U9CpF5kipXBG4GpsFgtSGxCczBW8YR/5NJ
jDu95DgDAZtXnyLPnPUgkyhAE+wUQPPHrkR4eUNE3Ufp/i3HdgVFkpIvnVBhHmZg
UJSs8k2GU/C3xr0gzu4gl7DCXryDaA0o2eB3yjaYpqc4rSDQIM0LAUAKKWoPaHn5
tSRytJ7A/v9tMTcdyrkyt7OkX4Lp5ncoQD6i6JEo6FxOrfWDa+/VOlBrG9NjhFOd
1gyaePmNy3ggIVFj6FqY6lOllj9D4pIuCPJgtSAY3+mGZTzau4Ctdj2+SC9ZAJ6I
rSYwCbKJh/uhBO366MdZGzo049Uk2F5qF3EdFH41It1WEV+kgXUjXv0mMneYvvPu
k46MCszUcudx0WTqB6/xQ+rXrd5SWq62V5Hz1MVM3aDQL2wEDxpIAeChb9LR92d4
J8WLBeI1qVRmJavIDv/bA4bfm4hO2pewi7lkQ8hYCFTJJH4HcLQr3hScxJEt3MNz
CJO6QObpXLqEp+ArW6xqVEGJzVrmOy6jwn4VOKMFn/N3/dIkUl+83DEIBYHP4APd
0JJ0/33GLx+JMJ+N2k/AFRbaf45NrvXpa6+5ZC+ulvwWUiWGsEISuMpA2+6VCqfH
p6YtiZ7OoLa3qLTij5mU9zogZ8C8CnlgqPYUL7SGkLWh2rWQjEMHIfCC08JjSVLu
gHxYZ2jALiTZL+woO2/LZzlaaI/Bb3HEXK457LNyTVK70zvsQ3bZNTE2aWcG+DIz
2vUNxXh+F1J1cxj2CJoruPn2X0fg86n5KumahYTwfx+DBpSdLa8pCbqoVEWIyJtu
sv3snB7K8axDsbJLueZvwT54IxmL3eMHXYfOTKOUs8gNk+e9aG3BVwrY4aYQUh2A
ce74E4a1TspylBFB+BA2DFy5vhcm4998hvv6m7vmwPAfCcwLfAhFH5JSk9UU+XiB
bHCMg2t3BzDt8jcwPtZJUPyHqa4We0D6Ib2kgIX1mQzcZ7q2bThLgMxuVo+ZmB+7
//xuo95G5tHDQyMoQJM1UmSOR+uN9OlUk3YTaPEN8xfgTFOAH5z9kVIOaHP6GSzx
a5LG9zbY9oInZpe6VtdXqceQc2y8HpOWRYTAC0Y/xIKwS7pn/iRw9N+drnvmVTDQ
dXuFfm1NSMEkDS1Qk06K5oxil6T80FRqItRhzHYFdFWHFv6pC60Ee9vOcPoUFs7S
ythooeFzM6bmsdjYpkz4wjXt5tQsToVnqzWk2Ay6XNmIFk9Abn0ZxQS8KLIeoKy5
1XS+/HYDzS82LrjUXc3qWWeIjFYM5c/EVl7b19GCr78so6TLjVMm0OqLLeTa8flI
gfmlLUgxXVtN71e5Bj2OXJNFXpgNYVzvPQfvoVHotyOsJwuHB4PVR4dUlSQfRDgc
pbynBHmh4wbE+cGKhDtmJo5ySEugJ7gNiH21yjSr+ReUD9zc3mdsRU6oHW//DUhw
waddTvKNprKbtO+imhyv3QHkEHaHMfW/xBzi7QiVJ2LPxIK2zvlj5WyjCk5hG1+C
L2BmtFvhl7W8kIlorfsjsiACXTdZT8T/NpUMickIbFC1cn/ONuNAWqYQ9I1u9BsG
6RqDSxDgr7Xlr8ZkD8JPNQJV9g2wC+fy8Oqpv74y0kfJW8/eiBfPYkksMybIrxff
`protect END_PROTECTED
