`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k3i50Z7/lz6/jTJFcfjENdFKSG8+iKDmjYwed/DQLQie7pjRZ0J3qLUkcA8rK2Lx
eoPVpwVgtmVbwEdjMzEasxINQIWP+zVz9V+mInzq2aj+JQaUeeZsheoRmtXYK6zE
QNdm02jlfHFPu+igQZW4hf1RUeKCrKgbOpNsZF50DH0Fnr5b7v5QD3yz1s07542I
nFms7uBdjQ8HUNRJj4cSVu/Q17VHuFIBimapOPwAM1AWdB/zu5cJsMRA+bsYracL
ATPTu6nQk19godkTLr2t+CnCju5BrTKvRIUJFqPwFmYLbxeH8k7Miuaddm8ryA0i
ukxt154S4n2KbUhXreeQbTdABBw8DPvBOBWIS7cB4IDur0DCx+anfiir509gFgIG
/rZJJDfeb9M1tI2ZLtzj5Mb2vC1Fz4/UIqF5DnY1m/qVrNxoHHCLWqDwQQ2N4Sx8
arBd4Kg/TR5wzfITtudHxzqhvAepAwyc2lU6u235UINJmT0EEnu33ZT7VFbo9nmu
/C6LgwlGW9Bl8SgsNkK/uGoTIOm6/w166ewcC6yKMf4xtSAuHalSG1lBneWJx4tM
3bFNBLWZ+Sis85IDxfjsQZkdQTip2q3qav5fYu3qmCb8vEs1px+Y/0Mi3D6eWbPq
yD8366cV65HmAT5U3TghY31NpExkcgyFZ7lqkXXPBx53EuHOSCGttDfGO+3ap6tT
jKmdfGSN7Eg0EUQpZOmbraZrTNKQ3il0zuA/9/0svqennjV/GlerZ7By27gjhhVS
O2kDuOrUSZreA2TjaZqm3833pDA3oHzcGtjXKxAyWu9a6YqMQsrzKEqOC4Dn+b0B
XjmX0FWfmXVd+7l9hNXQXRCb9oeYDJEUxFczYv/ELV8IMdTZexa2zLnzuDfBgqKw
6WilgHKLgbvx3t/ibxPET38dWTangAvakPJJewJfQM55uVL16pUlbTdT1P5K8kzg
EjsWyLrhsBAlbHuBA2MDyDpZnPT24djKQO42YPgyiUnDRA2UAbQM1ayQPvEPljKM
v2hKay4QU6w5pnNMB5rBWjBj1UBIu1v/DorMSJbf29zWjJ2SBD/zdR/mvGc1STxM
gjgG9zOKl63PXXMxxzex1YftsVxIfj1739c5xvN1aChUTuDqb1NezyHG1+ld7cyw
Eg0uQ31mWiU60GnYD1gsirGSO49qmexeJPFGiuFZGo/zoHF9kJnp/+svuKewSVwK
+ophWgLJa2ZyfjStWWFnmda4TmRpw+FYWe0lkSht/xznREFOZmP4f3hrO952LEOT
92ne4KW1TTrnXDljLrIreovGsC0n5Dh6C6x1YNJQd5rDrzGJuq+pbBvl27sO/6q5
I4k5mTTH7nHaHy6h1V1CPfDN+A4ncZQWJ3/hyLd6whfCbVEDDgwFmhdlQlCC+2eS
85IQnASVL4eTYwNtX5YjSmBEn/L0P11V2zPOwTfUL7zOkxKeahr2mGDFFV3w4gIi
xaJVqlhWBj/QC2FzrJZknqUrS1jT+vR14km0WOibdf7PNzL/IjpFKC6avoDVXKOD
iWxVJg5pvi40zwWl5AzClJa7gb23F0mqXH3XPGvFHoSo+5rs7NScPTBLE92yRAuz
T/50FUpZGBFZSHjnlUwhlMm9lVaulqMFJTDBZecFE406f+wMua5Z2pcefZolLYnV
qhIsYU2/JyDnYyBwkM9nX7ohZNvFeqqAlKWp4sEvTz+ea3RVRM7cgm8A+5Mgbrg3
ZmU4OJlXsY5pMW+/g0aeMYqdzW2VwDUhpKktfSLkuoxWeJ9yalBlF5v29LHLMOYx
dS73iqXlOv3LhXySJWf75wdhVmZenctzqWy9IUCDBArMa/R8Rh58lZ8bc2p+stUD
a2neRGyLvZ29lVIkX01kSwinssefJut4tRmiOil2oyk01SIcQQSgzA9MT/VJP4i8
qc+ReDnpwpT1qvDFWvIy+AJvORzroEe6nr2sBcKbOYk8ahIs4GLU37lDizJQTezv
ZXfF7RlZx9r2Z9tIcEvtiRM/sNLUM4g6aHkRscBYew5LjILIgQhvzfcrotLdNbTL
q02PCkGkwAzI+G+WExT4Okv8mNMIwDZWlJK/8DUuZCZ/9S5Mi+jq8IHn+KoZkfy2
bC8WRCoiKSF6GL3ODcrsM02q2CtnDGaA1S0Zl4WFWBhmxt3HOUDepWe/1EMjwfRK
2d4x0x+LTaXaatxlBMQQ53xqHp2OGcq6k8xbTQK2xgOjvPta5peSJFApfWsT7KUB
+Qt/g5sDGO55kJmAVmx5NBwTJi3D1dw0LPTPKvty2DMIzZoN3n/0/Zv8pFd6ScWl
MOp233ljpLUT13ScLPsVZ8M480vEQOJWqTWpwEXpUV4G2A3fDxkSq0GTJvPSLT9f
XyvWhiHCk6BxPSV3YQZ+OP/KP5kVVz5uay5mgBy4zGv5ya70v2/GZV59fDi3Kaux
M6bb7JR39+1PmMeB643jm2mA9C7AQ2apulZ+5StMVU9Jep5pgwTsKMu6HUKh4QAJ
aeU4uOjvx782MCIVWThukxFn/i9qAzn9FBEQmrIjB4G6NPThggtlYgiUl6qCdTjw
HH+HEjKvB+bLNSgFQoftbDlZpzByd9aeGZg+k0oABIYQCKw/sAgD5drdeXiAepUv
Oiof9HfFGs0LzCre6YfPgFzjQyLsSa94Q2e9Z5Gynwsgx4Umu2OsNyGshEN4zCIY
KdU5fTv69SVk5zVK/67FOMgMzUjlRJMcrUmwoI12Ta080ivePiLup6Ms9mDMSm/1
6xRGfN4eKAsWhd7ZrQf3dlt8PK8bOgBvOSyaOmF5EAp4+6Gk+FBjeIdefSxyUE0o
HzGSyc+jg5XA4rgUtgnIdfk2ktvbcTzkNuE4xWXgzTDmDBbfqlQHNrKg5/1HvYBj
+cMkt9XXLEofulbFyhjOl0h0GfPOWYYZmZ0pG7ULWQpAUpSvYA0UrLrbAgEK+p5Y
/UdkbHTltauoOrmfp7I8q2KjfyEQXWfZ0/xZRNbebQpTwsnA8svYw0U8dzoo7d9q
UvQC52l0f7+bVf7vGpjGTYpTS2cX8n1tz79qbqfkoQuXxRxn20ILhZt54hLob3E8
98MAnJr+eNZ+6vWf2RixOMz8Lv3+3CDcQpITkImIqHBVBjzrggFb1hxkJlMu8zgX
AthjsqyDJlMyS1I6haGBi1AhvzR+xdFHjZDn9hs0z5+Bop4/OqrPiYR2EhBw2LKq
MBHLGdmx0zDht2ysg+z9xw2OfJQ47w+XjA/79TUYn5XwHoJeIseX+EmrHNFCiJUg
WQO0Wfc+FXaqlwlIIQm7EWDabQ1JEIXbh3c+zPbSURKT+CiOocIm/9L7mMFFh0eQ
ZP4X12aoa9biFBbV03hYZybL6QpyTDIziFuKwWYhnreEHxbCNuAJsNYQoz2vabjs
wyeP/Wxl81Vfnv0cnHgGyxlSbbzMJKCf0+SsrVoC8B8zec3ASR/vxa44Vu4B3NUj
MUkagwyu/uxIcuGHWLZM/JKUlkzbt1C8grYnrlCSEVWeIsoLo2qwvXuVLHzPlqiU
fuATZ+cs9hCwv2ogc9IiMHZiNJYHVRRTPBk1/2guzH+qFTuuzTRnTLwNVFJR06aK
Dp6D9k1dBRX8B2N7sPRCudo4JQoSrEnJxJXmMdE9Y0dA1cwT4ayziBf/c1VPpYiy
1KOaHWclK2eE+ZEcoFjko7RoOF66GSzrJ8UjDa1YpdrdcRFCy1sXPyolexS43xdi
XYjYgdH5Gel9xIPJmbn5NhyEeW0DoHJ1ME/bQr0IjdDiRYlzZxzEOzwNT+bsCEa5
RZFMNuinvUJN33oF1loKmZJhth6LSLFvJ9XmqP6wJiq+pP1foAZwxsVel0LqgmWT
+BJusMBq2kSLfNrx+zv2ndGIJf5IWGiwCCC8rereJ76OdlNzpmO8mS866i7LsZqQ
WsLWEBga+MlaBAVHyW27bPKYiqqOgESRRwM92EzI2cCKunTP76CmT+Qopg+eRtKS
CAEmpaeVuUEhnsEyzup7DIKhiTifucBAer0WGgdjGjthqa4RocKA6NwfznPuEwvJ
MAiiS2Z9SjWTMN7ZHl6OQ1GaC5Kiwme1O+dN6Nh5aSuZ0ozKtqsXBL801UV97kBS
vERs6zZvedLGwnfASzXOCUYRSZr3BKg/il6j7SXldgWGRa6ZLaS/5KSfTO/QKzBx
a59Wd4MLA0MLWNJKjTd6BgKXzrnh6A3xG6VbYGylVCxxxHlCK4mzt9sGtdoZvT0d
71nxpolIx2BnRdHghzaYZ8NXvarBlQuGQhPGSpvYZfpShN9rFzE+PqPwf2aPMpBw
PHg0mbeLlTOo/qTCmIYkbS/j4tEWMXd+GH8sx3BqO27ob6rjq5t+atx1Vz02cfkF
OdsJsuxbW/BM6J1MgRqFWztYYmqEx0zeFw/BPDfKALbGwdWjwG+C+L5DQ6Mjwt/n
Muj+nM/sO7MAT2eZ534weOgFErZ2ZFgktx81W0QcbLn5B/vNXIqYuuiL74mNf3HW
96XfprA10yGzF+eVopRYtm+vATjK83dWYIWFv4YC3ugy1MklTkvs/yRoC7ebJDxo
3nc5HylV+xMnYYW8uegQaUUTqPNJ3uwxX6YBgltLolrvk9IXEdaqS+GQiaOlXThe
xoSkhcGc1FnLwnIjV0AWatvEVUs8vwKpa+DwLcj7Atp9rzlY91LjpxR/CDOGuDKw
XjW9aEYL68sdku64iGu+puGW/URDnA6HSNNcHCSTKjf/nxc/4ntFL6GNnawLxrVY
/j9zDsh33Dkp41RsJxmU56YdWXVCOjPsi5PG3O3FObeGdd6ELICobjaDwIekRqYq
POf+pU9GO3mu1OV5tNEIJz6agVI1gjpb74w+1tL8Hqj4lZNYaa3Rlt2k7kuFqHuZ
PERlJH+ZoiR+NhNHNZC8UmgvcNGbF7FaqGtA7Bte7TDV8INs4r2xZjcznVEH9ZNm
4Yl2PIyLgmkRPjM+1yC4h9HlpZ9iQvjNtf90muzXeffYxHNMLUNPTRhHLrp8QiKC
umj01Y9ODnm3jM2c8JHxGvRtqM2sqbaRGlcQlAWS40g1CkCidk3aTt1AVYR7hSGE
z/BVMgObR8eBoPLmnLcPy/E6P0rRb4Q1ZI9slFQmT2q8s71kpWTdl4REZNRnwbV5
+4jlm6VN1+ekR9XOcltXbQ7D+HPH+FctOdGzs7Hskjm0Oa3xWxHavd+lred0fLgc
rX5f6gJSesSYzHX0RHAcnZ/XZfb6tXX2/l1E1xtzhG3fvPhOLmSFqRB6mxSNmVQt
RIxouD3NQ0fQ5eJsPpi6qY7R+m5KLuqnk6NPynWm5WVPv2+cEcjrVMY/1aO6Q9EH
i2O7zsOn+aMNUlAliubOXLfUGvgSbHGxdRRTfWjI0/75uCqx9xzj5Y/CcMe2UTg6
xbvRjVCDQcw9/WETf918RtZ5dB2S16RJ5RNi4sFljkndCxc/HvzVmq4fru3HFt5k
6hkLvLwGMlMMD1N+bM5OrqsC8wL2lTNqwe92H5Z9aP/Ic+o5Io1uvM5A1W5Eqreb
aX/BszKacFf92mSdlo/j10ahtcxEKD/H5s7Ailcy8eRsNP6xLeMkaRAppap4+9h1
+kuqsgwjEgOuvySDrGjooQLwIZARctqAKg/tujPlVmKZrwdleFQiIa2OBLsAaEPj
74VrmsB8KEcdct3qIUtZlguk7evL/nfdhOAX7QO+i6h4N6VpGkjFEZf6sQKTk3JR
gOuDeNioFrpha8lF7sfSu0eOGcGgv0QJHZyj+zQ8AA3LagyT7iuCxWTcfJlYb00P
zH06V4aE33daS1OcrbRpXVg0XOEwZOnC089NktdacdhECskOvnGMgWk0CWOPKrxV
77rY3b9u6OasQqihm4lFnfnXBme7/zTInQP8GvE8HSgNJ6JjGiBTTX8QJviJJwAn
72Va1NiUO8FT8IyjQkz9NZYGZ7uLEeVQ+dqzzCu8I8HjMzR2+bQYksafauqGTcMM
bNuQO1H1Pw/25lBiQLVdsg048XVDjXzrcJ09wjXNWK9gQBzLExhwBq5Z13TaFiYr
9HomGFHaEyzuV4GpFUsqoHYlencJQOppVNK5SRZsU6qhD27CCWCvPPjg22/UWFbK
I7R28r02b6Dz65XSi6xrFbMNDjFTjevyr+D/gJZfQhzcB/DS4ZgxX1QwsFftm9Zi
RQhAhRoVtnH/8NAKU6e6Ej+9XDxhjlfeLIM9OEFvtfNm9TBG6MybukV2ZhYujSV8
Ezil3ja2K6tXIVMjf+2jC1VltQkrexYL1IA15c2p/5PjnmepGy9hImR9LbKZ0l/g
OCU71gH9tjcehcKRdVp4OILFHQIuwDNBIUj5zdxwKtuWFZoym/eBwsuSgvlt+FGI
0M3u+7tLqcPzMi/3BcUjZjoCkGvKZP2MmZW+mZhwbPoRxz/mezICdalHvBLTIgjU
FaUKo1953q1oD2lPUKRearHGLwY57o/ZV+2IGvSfgr1WE9Ww38QyjDhx15zuWCcZ
TTSBrhVsWZ+Ea8aFFj+nYJsrTalSgIQQDnwTePb+LgpT8t9/+V5Xpgc+nsYVAQzT
f9r8AySSZCdaamT2X2u8EJG3lpK9U7CMkJ5f0Z2scea1SjtUGZFK5rdVU4aFCk2G
TKSaBY9DVcEMJgT6VuST8Xr7WAzn3Hja6T6T2GtlX5neGXIUqTHmDqUsYjnUkuDk
eidgGqaf99nNycN8vdIuN8cH+PBt8cBbLyP7jBBR9xo0sTi6ducY2ekVRDK6NqrD
bjJWhTw5f6WkpJ/D5Uhho36KOQYj6Pl5YPNJmolnNkL7FnXwFdjciapcuscno5yT
eToE2T9+AfIVzDUS1hpOsJkyQ7fjgcAM6quZcilk58YNhijyswuWe9b0Nr4cSh0N
/Eu+vYLK71584B63HISKzpdqCJ5A5FbaqKu+F5C5rmhh06QCV+d1nR1Mo+OIeRDd
s/SsMeZpW9hyDR96t09AsMuwxzxSlJ37wX3LeRGcV8+K/5NjvxCTHiNxaGLvI6nP
NBaumVMj8zwxB2D2Ziq7uXCiASFGJjl91drGm6p/vZQ+k+pwzl+9xsAfsJWjD3b/
7yFowtRCFz/pqo3po8J58kVWVlCoy8+vODWZqji/alCsym2+cratJC2RsSlv/7xS
jDN2Advug+KgJTVBiJiF5ykEW3zMoaodY3sY6VA+CPKCcAbWr4e8iaw6PR/0kG/S
Muve174BpEX86l80toPsHyfIIawcZ0qCefx+7b9X0o4BU/WLPJdjQlGpnZNWE0wf
Fm5RwjgsM6B0tt5zwVWugMWhkgo9Mhn5CSpZUPcQHSKeHtjxQc+IVQDLSgv3XnVN
eG+HvLrImWgkmit1b6gqAVExBmPwox1eb1V4K7Uba2sgFpTkE39Y2pHccjAZ4T93
X4ln4moA7AsF/Coe8IrRf/E0Jqm4OuQBBpPFZzD3/lvSFN1UbkldYnBzdDB2xq9V
Eb7M57yUGA06IUdiiF+GhBmOneD53atHpWtPmnnxXouO/s5azW1DyQLL3qckR36j
kDcadLtP2g4x+/kut/v4I853rS+eU9pgFfy7of0AzUhdVHzwnaGVsFyZCiLLyGEf
VtKwngdHkNqsFJpPe9u1voNIUgRi+CJOywv6JorL8w6+kSUI3JnxOdYqtCQpcOeP
Jzf8m+YipoOMM9ZWa9aZWbG/6GNn28yfc156tR9hP72N8bAjQ4Fc9SX2VS+Y69g1
IFiw+PUq0DLgHmQenKIsuWUfaTvm2vbaI63/IB6zk1QEsAuQMAwTcU7Hgt3sodPz
nFyibygALl4Su9Fft+Y5fBl+0Oax/AhxQYp/dxbTpKal/pPmihXmtG4g9Ig7to/Q
0W2GHzBdP4q1nwv9dUqEmVTOm4baJgngQqm5vfzLcp2iiZ66OCYos53HxEyiThty
KmNsfjP7OgczFygL+Mhodr7nYbUHaN38WKdw1hW7+s7XSnENAR0V65Tey4Q+C/fV
YzKBwxlQLvH6TbluF19516V1zvN7dzMKb74+OVhao8lIJB7+EWUF7eIBSA2Pd8nV
wGDdJv1fzPfhf0+xks7YcnbRTYHW3Zz0ip0U1kRjInSvgsF/Bx1mA4NodXskBxY1
o/ns/ry8lZp0k9IjwstvdDp4MLQSk7TmFxzAKpOluUVZvQhf+vy0yswtAhEO3nNj
tsboyTzT8AV6y9RKVzzh29nLHy/X1r/SfDlHqI80ikCy9z9E4fgLoRUjoCizx8vq
7HH9NnoFsQa/7OsW9qV+IOHS6UCn4+VVgTH6Cs7jkkvONSewW0yf9AKZdamnjzBZ
sQ8zRC+xaQ8DeUdpQVZ1r9i7c5ukqxJZ6CaXr5JkrNRVXh6RDbjVbRuDj8Rg/p2/
a9S82/W/ZTGY4aUAQuMQVIiSGboiv76PcnM1aBXmmTlQksHCy79cH1u52wtUrdlV
ogJONXymI/hraU+s2CvDDn4UExa6/6dIn6GQ74ee4nKhncEF2Y1GVngDYjslb5rx
uf9q1c+Ksaquj0ppiZ7QMsjUUyj+oqfjmKt8Ct8q26O1uoL8fyz7NJhbHPtBmx9X
bYE1YHNIHhE9yVg9mktkkmtNLcTgZfvOzcWlkttHYqqQ3y5zOWCdJXd8QgMXRiGT
LKmoT2+3LeYMT0FVTa2QN8J3lKvpSC7whpDv5beEGOlkc95wDotnHQIAFyLhQZ9u
B0vMFD9LKQVQ82x+boMntODJcRWULcOoTvd21dU81G2KJ/5xx8a6KKKLjI7fgRbE
R49pQv7rwyz6WV1KHon1MUghbiDRi7NfcjbJzI9RY0euOzsPC7ksYutyOOSMnCwE
41BS/mPn4ExcQccKT2aIjSd/qzG24FqhWUfOMJDVVXVbm6l4jx3sjTk2kzCHe6VM
UsxgeiH2NhF3h3KpQ/dU76Rfl8zu1eJaI1Suvr+OzxiKqZKw1m1ZfdRSnU5ClWJy
HSJI0c4T64rcGoQqfSX1cisQIq4gfOta1Bf6XvCfWKClEu+icd1KU4Joc5E7BTWC
etMmp8qQknJUbR/+cABFNR6stELUyl9LiAymISPTpi4ynDyqny9ZhuVZiiPM5zM0
FTHJobfczK1H6e1VjnJvWr/xsOKu8WEZ+4rpmy7IMHJlmbb0keeLozNH+6ImFlYW
AvvVCLa7wL5Ndh/hSMi6zhokmaJwY84aThRnhDfyFcThCa2jEq+hM44qb1FF6807
SET+gelV+nY9Rb/Y22frRvhfT+kcoqtwJ3QNfDCOsoVxd0pk5NfWpiOexnEjnqsK
pniOYQjEZpB9q3t53VUhoHqcyWBN/3ED4BlGM2vg7FmwZauVXgnA28u4jpgiZ6JE
X391sxRGlFF3GLuT/eiR4dc6zdQSSNzwFD7SY4sWyO5IPTvey2dJ0KEdaMqkihG5
KzKWRl0mJlQw+Uwlx6OwnUseKuyWPWgQkctqp/nlQSusEDNklPScNgy+WfNy887N
6AzS3Ndq9a2mYS2pORsMdF8G+Nt+5a+5Jt+GAppw8yw8GnAXCmjNP88hD5VrzQza
2qrkENfYo5VFWu8kkVH0//XijzKQqZDt1+2yiPedCviNnlJ5ZHAlnigJHDXZkX94
1ITG1rKzlFIMf0BWr+v8PA01wfErLMsVzhdoLQrfzOLQN2xj1v8KOpfRkw/oxERW
+PvHL2P0+6GfF8QvgWtRZNK8D7muuASvYivZuI0fxyUKXALKlNGRdNxWJOjHY+NI
9IpoYR2EW4u872vSe2uUySZ4BZv56LBJSjEPCx1cguiV5of74fuzR5BG0rLtW4+4
JTcu/Flxy8Qfxek1Ufb5c9BFyHiw9NAdUDkorRHyrYrHjfC9HrhiEYKWxC/QAgdb
3HARjsG4i4jlfAnymcFVAdGEip1qfoFKXcpok6Q3ZK2iLbtckIfgEPnQUt7I9+iZ
6QlWZWT94wr2jRiHho03vv8i37ijdFGaUiOO3pU8FZq/jPBg+dzXebrooQVkXZ9Q
Fd70xBnE67cJyUfBY76UGRGwgZr/GFhDEKVnFt9RXLTYSNI/gNb6u5r+zEwC8E6r
T8WmuGlnipY5+LsEmK3lwKFwlfD0I6VjEbMlki+zGpEKR19L71BKdzvDbb9jVc6T
FEeqP4T8GTHFsGUlt09YuMk35Wjhmfy1V72Hd+tSe5KT3GSots1+KyYiiqueQU/7
dY2/leJ5MfzN/JeRMigkLCszL+aEvA+yMvYOZggLt0BZpZJ1vsQXqTq6qo9YmKQg
2b8SVg9NqrgeY4ze5HRgkaPNbOm6vZ8TkSrvQ+3Jf/1sx3+HCaqhf+DRnj6X+MKo
GLaCCMV96O3zZvXgidJIGJwhB0+cVgc76SnBr1WKnnf6IwFlFgoVkfVkaf7KWijV
mkwWA18jufEuYYOJWoKjGH3QTTLxfToyoj8NTRjRD3nevtmRRNy/UuM4ZzBNbsXR
KLPHyP1q9K5JLm2NHGnBS+jD2fjaaU5SaJKgsWPwt2tKQtGFzuAfx2v+IVaQYQyd
Zn3bYJ42F2mMVGWzJGfPfJdhNnI6fIDaEkNCdfTVTtcqNXemO/iNWbIDMoD2hhBl
7hgrNn8gBjoE5OkrSjfFgwUsCVgLntfe1vI8qWZQeP6iK9lYrxaHjDrvmKc8n9iE
EzZT5P2zf7rzMXdEhmxbk1Ti6uAC1sbU6jE+UHXuolzW8nbzgmQdbMMcuwE0zK5G
173eNTJXvBwOQHhLFMJHIfQhl7gFnyJIX47yYBjEJp0HCr/IYyKWZe9WzIknh9SE
r9xVGuBCdotP8VBSoKWq9cEFsf+gIlQ3FbsL+jslkHhtjuw84CUuKOeicr80vBBq
5OCS+4eMrQCpx6etwDSqSK6zt8Cz640hPYu7/YIRkYhDOl7fzYWEUIyc+wSmUUUb
PsEipzIE4naQg9ZhyUMJMsvPBqhDzpWafIU+vd626AAwHwawbw30Phkc62J24cf4
+kvpLnelVXGTVCyzwd4ObyVLPQKKoA9UbTtokTrgTURJekX2x2NmmJfCbftOCGx1
PZ0abfyBzuXWfsh8H80PVJpcUPWiENKl0Tjnv0IChsqDrrc72azTgCf5t22DPxRZ
PM/OMUzSXKWEG5Km5/fPbc1rqsIB1UEbha38DPJMp1wO9urrIylKFfwECS7kM4uy
ns9ZZ79JUZ14xQKWrIfDoH7U1I4nHVN1kMQS88af2uQPN44y6LC+wvm8DyDr6fE5
OG8UJmP6RGxQGIYs6/GDQLjG3rcFiYDM/Hv70UCyMLIswaR22CxVQHauaqFKwt4A
`protect END_PROTECTED
