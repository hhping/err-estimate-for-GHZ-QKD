`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8ZtGmSS9nXGOisbXfDzIPXk/rlVNQpr/bvv4eZPLEwQMRgr2vNzYjRfXVjr5Oub1
AjcahQswDsPBPNCs2SoYc3kez2nAbtXoJubXH4mAV1U2uXiynMxhd/o6WOPBmFqT
NJIlnrOqN4oW5L2PoytIRewxywbA4y2jHibwn53CI4pcMFPoLLLL6957g2Ls/mNO
I6ezveLG9AWeEgi/iM9X0up3xr75ZxOenQaduer98UZPCPaRZepnq06U0bqS/p8C
0uPOPHFSFoSEjJGQHQYfAeRHDj9WEq9f5/yg0y8xM4w0kG8z7IlAK69A4edfyeR+
6ZQc9E+slOAJHdKi8qs8to9jToEF139TdCNAb6unxSvKmpHLDbSk6LyOfCNkvql6
RcijkSnOwUTIx8AL3FYJ1NYFo/WtfM4mIIdWDuNyB+lijpkbZ72QjuuF8CrJ6mCw
l3Ym88Xew2O+LdA4WWQ33LaIjqIrPSmYdiZRb09j8ZA2AcyitLEqlG4Ulu8fRF1e
0yS5eYLxdkI8GlEWkY/fY1Iaw71x8gVpuL/AEedigXyvs9H/V8HUIpSEhwvtowwV
HBg4W0b6QPNpESoKYgg2Ka3LnLCNWlCt6K0RATcDe4gvnpYlPO1h/snvuX6OJ743
ULuWhnuEx2JhWVZqEi5odX8/VTQy8BhA8h2d8NJIkqAp0ketRyyYGgMOIX3LkCcr
KE4A+OMlHc6/SXRHdcjb2vIdzh7AzfoA3YxsEapJW5SBprV+t4RBv3tamWh5bmD1
F3ZKA1bPP9aB15cKrMoMh31kCIyCnKtCJt971gGEmggVBf3aR6+3GP8FGEvHFA1Q
wGSlueZuAlGx9DUR0bQCPKFyx6LYklMCojXIegX0Eu7jehBc/DWuCXpCvDLD3ek7
vAwZ3J+e0bihxgp2X3QToasz2uAib5IZlBnTiw/0Tlq5tjz726vGhpE92sKaZb0s
5VNjg3JITkHeXVeTkvd9f0P/j0DAEasJ9XwPxlBKBue5VwAeGFyYmiSuZp0PA05h
8PIh85cgxhLK7Uvn16HSCQ==
`protect END_PROTECTED
