`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d6qg27aCTD/fPSgp0BNwNWjIAxQAYxgmETWWnV0mpezEU7zIfUUyGJ8tMY1neG8a
IgvhwGTbOJtmz30EtIK+STjuR9j0f/Sly/5AaCrF42Wpzy1TiZHEfenDwTu4fCrI
47hCBgI/3DTQLJvTpHaZJQ+9w0D3P2hH9s1wH03NE6qtHyFRoNdHhao7WO6B/mDg
OdhmwVJ2yejDsXCa8H3Yy5z1tCaRuIEXXcz7A7nQX4fbmV0kloBV3Mw9Ij3tRqXo
vxMi6+lLE3cIvEyd0+vQinFN7DazGazwrJYXaMgfrVX+2JsMuF/XSbmA5zziv+IX
TxozphYeVHqz1jrf20Q5o8/p8ThvidFFsjyJhhAKWjJ15cdRehwJP60ucyExtJEY
K7cVZdyHlDVAbptI2s84Kk83Z0GVBnneXA7SlWSBQvRMB8/dpNUikbgHcu7qNBvw
wk6FDpxgoxhmH57/Bxr/0c76jWuKmlAFEZMUmeJlB0B/VC9DbmRjtXCSbl1WpgWq
gBg+Mbq6kkByq8N3IL0SI5bz+cmim1GElMt9vCAyJDv/1aKFEmJroxQp1zMOi1aG
Ah9Tgq0lwyG1kyJEzDrCeIFYw+UGV3PmH6GN24CiwhcCMFMFGwcpbHX7rwTkkAm8
jDJVZwXZDOWs55rH2GuUt6yanaGBMVHhT5sqLfGwvnBO3dHWIbbktIFyeiqVz/4s
NQVReTSIam7DUfceY2DNlWB7LW/d/riwhNn7xSP2R3W6n/DZJ9Q6ZRzTfXXCnaAn
2OZlu6BDTmrJTCPy2i+iNspd1Hrq0w5WKDt+F24OFlYyJatw9lOQ9+1/23ocZkA7
HIW7uBv3/2kzwlxhNZjRBLtDi1fsClC+WUKWuJYziNIH5XHAhP5KiaI799FPS6n2
AIChuKxq/AENNGQuIkUHCU+UI+aUcJba9CAdo18W07Qeq85/8eD8FmPSYkKCUm0S
dYBCrMgUpbwr6x4k/QNEMtOO3f21N+NMxNeT9xTxtRWeq+cbigpG66KRn8mjeR9f
fASa0DCo4+vZ3/lLFDAXgmh1rQRLSBk92OjSQQDWKO6MQ5GkzWcsfrZjEsZs8Vf8
RPePcSc1pW3SnptHcq4fhh/F/vBdkB3xI6IxArBqQKeIJIOjegks/LyQs6IdrDWe
1jc+OvbjcogfivpVP/di/562jAoFqc6HWt0Csa10ogljQiMerY24/z3OhfOGE1Si
xb+dgT3WcsPxsLXq1CmM3A==
`protect END_PROTECTED
