`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TASip4wQgWhk5KgdyLOFh42hwGPPyje7TeSwGFOdCiDO3fdoAeSgU2vasw4ZTqi3
tc0Qu2kjGBy91NwJ0Evx9wJIr0H6JC5WMRfOqyVsVd9SCiuKbR61/QYQ2Pgpr4B/
Zh5zFFou5fTls1NpWTFgYZHY4XYNq0A4hAEiXHJuwhf142KMSvyfxS7gMCG0zTaj
5yVf42+ro76ydx9k+/NWFgUix/8yL3YN4LNRe7mLHaFn6ad2jU1ltJKtAEjzypze
ttCjGNwdZCj+uAjF2ExEapEJmslId4D2FhGgARwXEuvLPExVnrCchDeckhz7yB1F
pf3VXC+MKn4ktVIQqOJx4gYaDkkZSSvwvCKhJzcJj00PkHPqTNirlI74XPDvqwY6
//OJrbzVFqMhznaApDzTHGApT/wb61XGKCaNsamykjjCZOsAYeaHYiiOYUzHUxfb
jWnNj3hr9PExMm0cCBTukjEtxSlmIE8fc1+jRYpeCcsZ41DslOc7XoXQpuuqABoC
gfNMEm4dcyPEDEIcUXTL5NpyEFPCNmw4ylELgw2WC/OspdfjyhuNJTKOTUPBJ9go
syEj5R3+cbhZm6+F/0DYyMEednZPenjeLNfEV5H25O+Z/PvBIf/tOV4WyF8IqMeU
iI3f2Cr83YV544vHWL23sWjb4Jdxq0687PB+G+aeSZn6RBd9djtlsJMQyin10mjU
G0DMwLWX1573H7jdCyeUi+tXoxHWp8djozM06Zn7rqcNohZ18vqIz1pf/x2JTOq4
smi8xKK2HeOOinPUn428kivSZ3SkmN65dF4EI1GthzM=
`protect END_PROTECTED
