`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JYBQ4VQ1dKDanRc3HMkyh+rf882iV1v1qLiAFe9Ooda7gDQyngbTA2benJ/lV5be
LuwSrRkHKw2YKMlu+1DOv1Nk1kyr1hmP2jN2QJnCE2C9PDBdirvzcwkAOxo6oSHN
PeD/Kb6aeoK7EjtBZbpfVJnktJzTUonDY27zVxzzy0Q5l9qf2TMLqWNdBkiGfZjh
CLJJfYlwAOVn4xUzh8s8kEViMUkZSoikOkiYV87moVFHQYC0Ea7zneziOuzmQ6io
lEn9DUrInG7FkTM+LuPOIUBHOXhAi7ZoD5rwo5+xOlYtj0OTq1otItfjvs1lsY5d
2s2hRXMe5Hv80EODZjApfgdS0RXwSQDg3b7vWSPwwXIMRBmpk3kJDCNhl56MEH0S
1oD5+kqTMjweZwGPhhn/Y0Ct6x5cJl94U2/r3DDsI6L4atc/EbE/8nBptDOL6wV0
ZB91JGysTdnEqaocYrktE5mCgUvZuzey0i+tb+1/V5VKK+vviesGhh7hpxoc9KgB
P1WKszsNBLgqPTJfEWD05hsJsT4QkTS26ChnI+uvv0JAjSa/wXQmJmBLQquvsI9M
`protect END_PROTECTED
