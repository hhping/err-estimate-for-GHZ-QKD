`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eO7RdLxNVrHvP+zCEZ89+Eqtq+lcCuz8QiY0KGdiFIokKZfOw+UBW/A624VpqDwL
KwttFldxG27hn7sG1LktFCk1RsBTuZPcfg+7B6PxH/etkc/DbHukqB/PYoXIGhyM
ssvSz79/JjON3QqQC8/ejrjy57t+Pe05ePXqxbDdCL9LWKIO9yzP8+l0dZMtaMR6
fMPSfC4lMoC3GsgIaoBxXWoi6YlZ4DUhZ/WAwVzQzbCGA0xVYnu4OBxySAcKdn+E
BA9ikQxYGJ6qDQ9r6fLmYnMhonjoossWNJILuQkIP3GE+02POnrfkrFVaex5nFuc
PlzQcYNdGavevOb2yP4aZgjA3heRk/5gjaow8u8s6s9eyQXdwWcgbBmMfAAbGJ51
zG2cFSG+tzZhQVjHBjX+IoR1KmJbQxN5u4LBMHrjzQqpP/1UtDE406B5uVf/oItT
FI1K1Exxz171NnSZ/AmumN432gBV0vi2yBbK5O9wN6TRQx/nUOXpitPZNlXJ6ipN
yYus9cH84PWt7wcY+8bTqvAHMnd4omKRRetmHjloJCyjXD9+NG/CUwa4jxcCoUqc
yyah9wWlV3dk43cw8wsdfRyLJSHBGrv3huFf1J1JRBqS1ks4UwUMVtI6ZR4tVd0n
LT0hwLX2dSnDLbFdBtZNgF4SqvsXASq5dNUul3X186ccxD4rOns+REBFAEnnJov9
oJ3sbwcGlgm7MbJ8KC8ZJw+QiUb1CAp91z1qYlwAT9R/ifiOAfNZO8Kj7sHkLBec
fkz5pNgGsvOprFETSjfFRFe71hCCEKgEJ6U/oe+ZY+eO2gTVP08YbKyLTWKPnPtk
0dbF1AnIj+bViQ2hgfYNvFfrcnvRfWADcHMmUBKb7uNZy7mAtPIeRsZo927CSiXD
JMMKaXKylKm2CRyE6206/Fapj9/rlcDLqJ8SuRECtMuFluk95nblWUrIhSEyJL1T
IjTTdV5VeIm2GO9hlmRiAXiUWuzTOQRlTfoUnu8VPgbTNggHYgq57r8EsXCIB1/K
sLDvKGaRi4yEQ3s8BwtMTL0UdI6SiRov3yW0yhuL0z6oc2zKdmo4ql1El2/deoKP
qUpn+2uTyYPbVKD0Si41h37X2+5VQzPK42gKU9+/iW2lB/1Jkv72cxs94TUvy3Aa
ilIDKJBofyd3Nb9TsJvhzmiR2D0D9TtdNwf6roKhb6DvWi3pNwYDkHRn7O1/XdYh
TpSModr0PpVkjSvTBy6xX/uHRlZYtoKkzNMVb50IRBjsMtg2kNQGj2XWkvsMdWSO
NXjx+i2ajwAwYqgjXEvtvTX5PBvKy665lI5+NLNzHIRM/p1xah/7MOPJ3c6prCan
s7etAWn06NG6+9pDubFM2GIXuMBbLErBXkaDcgKj1b054cS9luAn/OeQqsFQVzEk
0L5Znhobi6airKf6BMy8DDOzjUOl+LygE3L82LGs75ONSQ7imx3UZi6bpDqNEIf8
pDBRTCwIo/5eOo50kO6/TjCRncDwwxDxIBuwRD4ea/i/RwSiw0ANmAYXi9Zm+Anl
7FG2py9RXfGLRIOgplLAjA9wbgFa7qIDlNmkOhK5/BkCDfHF7fy9wtfbMjCJuYko
xma/Np+YKk4jzF+qWBJ9/kIvris4R+tz7iOouudeqA0SInXlK9nH4Wgll7xdMm9T
3Aib+mKYcY5v4fw/JbVtUsJY6oCn2xqFoI2RnGIThCsgsLwJiiQ0ZI61NQ3C9o1f
7lcF9Sm5y/CB00vdcBhf36R8ja+KQ+vYLWdVuc8CtXHiauSCjrvgMU0ci3PiyLpq
Q/D0GCAhyhAvID6XWBwbSecmFX+qWbBUtH4Er/tHuvgNK00uSHd4YxyuQxGNblcK
3mr/4NVLxDXDDB9r9CcWgA+VGfHLIq9Yp5zdf0nBSF0CVOPj7zD50ipCQ3tABf0K
hPtBRnBUszZUai8l5ch9mdSvRdGTF0nyNIAqk2MRJ8zoSnTmNOMdw1h9sq6ZpN/s
4ZMCLN2kFCc5GTkuSy8EFLnearbn8v0Xz8dEdNYLlEPkYbM1EcD841U38LinotAL
VyWT1oHKT81Hs6BCWCYaRR09tHTF6oVP6MnRe66mSJ0cHAV1d78+2OvvcAJLbPz4
0T8zHnrqqR8c8L02I8aHLV8wewm/8uAUiCembstcUWXUZog9wcqY9eNej+ma4lmn
yasIpRF3yRfMFG+z29WI7SAVvleAZY8I3EzygGTrm2MgmhgZNcn3tQnfr7jJRrUI
LilUfhnNmrE2Ekf/ThzT2eLdBzg760rfr1XuDgUBBCwO/tIk5pQE+v2ZlzgCX9lk
jnWizcFWmy5UQ/Nk3HJfVxx7AXHYs3Zc44vto5SgLCZpeVmkXVZKODxs9Zo2hEpB
cofrCAVv03iwkHOrqJY6wJwf6We06Hkc8ruGZ50YFAh43oeP54X0zoUO4wTijOV3
lLnsbSpSvBlqJU5qqyIrBvcijNIrHE+pxOZ4xx5Qbnkf58escte/sX10QmAp0pRN
mPIQpNUR9M6eLGTaJaE76ZHHoHFb6bEy8Ku7TRQu57Gz1ROmU3Dqu5sTppMhu3ja
KTK/fyhU/GAgiPMFSEgJHmT02iAON4LiCGg6jXj6PPvOWUb79DCRI2oB6SznazRz
j+fhNHI5lYqskMfhU0s0Fqz6H65OMy73bsPDn9fpKUYxdd+v5U9y28KZBXaBV2Ms
`protect END_PROTECTED
