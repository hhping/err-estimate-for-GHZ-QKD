`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8fEgO7RlzpC5dhUyJEUmOgrtVYNFmR0g7F9pJ2I54Bn7goCAAYFYkk0iiZ8ZXvtO
jHxzWrz0ZG0lhwvBpgteHIn1KDrW5gFzvAqjHi5TJ4KxNMfQMeZoOSD5LrjhSHf/
rqusrwkCxph4PGO26WdKKqnZ5bxkbSRrlaPqmxmmI99PHtIPAK1G3tfdKn9fJQrJ
ClZOylQq5pFx8xoDEqeSJBUxOg5eJ8A5OzcRHoW1WnBmzeSAOQ22KHqCy3eS44J1
5uf1twP1JwI0uxmylWysYD/3P4GTPUd3kPO1wI7R4cY=
`protect END_PROTECTED
