`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mZPGZLhLtwxGPMjPbyim83jeaghdGShUHgeSm7QmlYCMtArHzugKc9lecVXg8oZ9
MYHffNc0mEdn9CuyimqnVB1tsN+NLYiW8uwuIYeK8aeY+M1KGVpOhIm7i/pxEj+W
/Tw8s+2dj7XFd048t/e+/fP37sqLqNkNMjt+ZsHhk5tWHj75xu61tNQ42XmBloJh
2G5xYznyNyzbIP636Eg2x0aNNcVIPRAE7ceM8FP6lCJ2e7vRBA0Co6xZt2q+IWcO
00991MEPSYkAvjlNWz2ssO13wfakwQ2Fak8vQ2PTlyTRMOOPXJ7E1WN4Zu8rxCQk
W+wD56q6AoKOUjZcZe01GXXMWhmsjjWbMQ74sYsib7ImrgYmYP09gUcWetE0mjg+
ldYmubi9xEGf2e6gsNoZwz4uL8uoe7TSLC0IBK0izPn0uFLeUqs7cOYImAAVYwBR
EUzPHe/pK9hT5PjhiCzestCr6g0TW+4MegKRwy3ze1Zus+9C73VhHOOCQhVFOyNP
jXR31bceOmHO6JLOQKBeAfwHkK7WSwJtZjtbHOy8wRobE3OTfbEN7cHXNQ4qi/ta
jIv6KzSsK/ANvJWjb/Mx0x0saMqT7VhmIWgn6Is7Dpl0xM0y/uDdnW7YZg/d950k
pRQkIHONNzE6oOM7WoJ2FWyIIIPDG6hSzguXSWlBFisiy9ZmbrTEPY0RSocXGj50
aM/pLcPjdal9oKIAA0mDYYs2Y/W/KKkMpcdE+3FapjdTG06NLs7F6DMwt5Ie1TOE
K1QwdZcQCWA4ROKOwv+XslXTmVVywNzRJndo7IOvbaUBFUOw+NwQW2OpLW3SZtho
OcufCYkzZo6UHTGyExkktTJRA/GRv3l/2AOlUxUJdweLyM7hwHcfZ88CpzjHDcPn
9hDiOCoQ+08uGE50nhQl8qISt6zvLVluZ+etNjY/6tuqZ9DVDbv/+laYgpBoYPKZ
Zv6QXLDU/eHkkqXTxqONdOsMknXWSe82dRLptD5HVQNoz2uaVedTFfKMH72B+fqT
enNkGkNyZE26lRXepoa/zTruLgFoIZElmyCj+AgKpTrq5s4qduP5GRzlxHp1OiTM
Ey0Efvbi6o+KLN4X2ezw/NkJtXrKTMTwBjofv1aROJgf+njAHCY10mzdI3Lr98LJ
Opx9VIED+sK1CV7AeOHURdsq5nXPnSoNYtFT+azcmRa9G/5mCsPAdhdlBYH+EOdi
2pzO34lYbMw3JCMO06uH6mfHGgHavEGypQL99PSLDdos8xI/l75ZAE7LodGReYMg
5/xTqrJz08AMTkKPSVbNKPD/OUboL9dGYmiZzr30Ui/DfWT+Ud6T7WkVYGvfU4mX
fUEHGh0uzB76kYPjO+xtBDCTmz/5ilDShpqeCSXUw0HH3WMLnpbGcl312O1tDNjn
LdIumvore7ff6CIIzhT8Ia8dZzz7yJmOi7QE12EApFMlXVqK+fndrfoe4sJmw0x0
6fg9ZQo4c/vF1PZOluDdJGVbJ1W2AT5QPRnSfdxKir88nUqCLc4isaeHKVOVWfHF
8QoSFPRhAJqiOZr9FL3C/JbJnhzeIhXTrh83IkVhzb9go4D5n/YH38lgdLZ4uo+b
Qkxg/LF1J0n/6NhXH4YQ6HnoFrTE1PaC8eY+tTXXcxRINMomby0mxjy9BjzuJlpg
VS3GMddPYnEmGg6s0QUj3ObUj1U01fk4gS/D3AYfEoEJJgDaVKrnKPhxT9bM4f4T
ABG3j1pymTkGKUUpL1glgGIitCR1pk6kHrCwzXDVosQAM5Y2ek2VUfI0EI+mYLpz
8CTH/NPiMIiPyDypVqJhtvyKN8B279vtlU9aSVVHdLmutPc6WIkZ+QoRKDEvx1tv
lVS8RJGztf9vfzNFUpKpqR3q8kHyZTfsCtEWh4cG7xuf0oBDJNvWFbu1+F4cT1XR
8xvi5fVMLDFla8cLcCul8MeQn+hrm3WlBClTaqhP8TVVv/Y7g0zUsAMktCU3XX4n
5NhF/i0pcUDwx2j1oxUEgjIy3sek5COFjM2nCATfMNjJoQ11id0j4sRJokyqHYou
lazBsB5xK37B/XyO2SsR/r9VFIg/OSvklxNneiztYNyJqSjkPMBe9Ny/7n/wNRjC
GUIrFK2K+xFg2/ROj9uzeE8FZAB7Hw1QRJ4m0c/KUj0/fxo9l0EtWgdDO7SVoila
vjCmPCJ2dBNmwnQzYNOITjD+LikDju8pVbjsaVS2FNW3ogq5WDQLLGK5nXPT2jnm
QsSnYfmAPeXGpnaq5oqVHUQ1uurAt+H7zjAtikeCdPti3Ene79pInoWmDJgEJog6
oSgbznLSv1SFgSkxvQn9gkHk4PEjDyORRec1HByW8ZlB74+PQNyqWl75hl88J2Zr
1iVQ9TihKwZiMV8LMUsMO4ILWkWLxSPZeuhmyIGUwvLtsAyEpe8HDMBWgJTuyjhy
mik4WuqBFHtH67ngkZQpGIYp4oXtSh2+BjHrCfr113LffBgDU75z0FdD/lqJQo3u
Zv5/BtKoOn5eyWm4Nf/uYPGt20FPV4ybG3qC5zPAu12S4GoIBtQKzIfc4WhFKRiA
sNh8K4jOd5Ilgt8ur8HA5713p1oYGRpqsyf4gQNC32DErI71oP3Ce27lk56HuWKq
2d5KTLcLd8ufCOJWILsEJi03E5nNVUlNSw8Ce5ccv/lhgc4xt83uPDLwFBbhm8cz
f1LgU2qG7BqUZ+HOe5KWEUi8BrJm8/J9EeoARXwBR7+xsVsf2goWpUrNHnHt1anj
xO3ncV2LoB0cSsLHkfRTF8uZE+94Mggl9+Fs0ZWIHe7qzgAC215nYAVOaclFAdKY
DmCnBoaMooJwAcM7Vs0to+Ami6gO6rols89Y14Akik0RidotuINmIehvRYwKYeit
tVUtZh4Nc0V77nPoljtqkivJtqujwkhqrzjAwVoubBmOHZREi/sqBLO4OCBnPBTB
siNe3SwQSo3K7y4K6ukHSa4rutN19v8nnLWMo5yMiXIrDGkV8KeLxmT77i81Iedn
/R/LuutZDYefJ/Q3wJi1f+5yevOAflBOB0mMzaa0ky9PiH1Lo7B4Abzx8nby/ogt
q528E5go8AfZbBm3fRJhH6Y73LhzPSfXvDJb5FuO57UNLq+jCTGq43/v+RJ2UQYd
nAVmcAt+dpThSgPVBh8tv4eAajGbwIbxQ3dsa2FYf5b4dKymuAftGvy0zgegQ03R
pSI8eRGh78+sgqcp5XvWNa9W366ZGiog4x6OPZr0SccGNS4/K6OrrPJkHSk7Lwrq
uPnb9lY6LTWUi3XTlUALsrE1pqRjDpPOlH/al3jUn6edK9p++nLdp8XSQafL/SVG
mGcuQE5Z+ri8cBY35DoPLK98HC6PIDrg0o4l1R4TsHe8/KMt2+7YbGEaRqLzwKa4
4Sur1OHStBonIBhftXPI8jJsHMiq1q2ViYieEZiWGVXI7T573foofhkf4aG2ZJF9
5ehCBjw24OI6j4mPrBlKPM9n+Wx4OorhWSBj5fU/xYvq1UG+UA8p4yV6vFYgRxYs
0czSqp3bEaPZAITZisKDCbjTwbwRZW1hzK7nwM+EJy6pIekvSyWEEneqIyeQLZ7+
WtH9S543KEWcFLiLlTlkz6FO5oVXufYlaEF+Dvhgs1XcPn7V+NQgBxFkveotxdVM
j0qQ8we59GmfqH1lGAOa2MIk4NLfn2MyaRHyXGOHGcHvCPx4NJcQWNLvRWeJ0+Kw
hXBwKHsntEmEeGC8muZiSx6uVFqxBdgGaNG/HqNzPA7PU36gIO8uc1vmZF/hd7/h
BhOaSvqsiDWn9tFSvvWlQzkYm8F6jIICOSokivCf/5Yxm1smp8dLEq6fHpx5p8os
qS4pHWCR/Q50hqy/RZ/A5NKu5+OPoZvkIzJJvgT637rzxYU4RIKqZV7pTP2mJ1PE
7fvCsQm28WAz2Cs0n5gmJIqVqSWNw5OcngO8zT++gb69Pk6AvT1WW1xBgpmUPSxH
lP4XWgpSc+ZJ/SrYIQw5rjK3gyQbHi27huaaZ0nQB0p0dmmti4HsveOkWjn5b5Yo
91P9m8Fk5kg21RtDZ00gIQtJuaaqUDgaSwDtQQbcoz02Tw1tJUiFM8gRYoAwEm8E
Kq1v/1bNvNyNFGh+CCK30mI/sc3JYuPnXjvh7Q4/8FLIyojkL4fIBSVcTqpNxThT
d4aIlSAJf20HygbmtlX+C04yZQDAGF7mMwKMFAqJYKCjMZKyhU9hajR31qakfWbl
0BUrVdpvQ+08aaDyiqQ+J2n1t4+d/jDDHQ3WfUQ8FiECi0jZbV+rgLCfWyXOBPsA
44RM+1DmGMknF+yM3r1OCGgkaFc49Gm0ab3ofON+haHBm4g0xVYQr8nQ3DRTq8/G
UPRSER4OPYqdugbINlA+xcSl/8uBzfODICqcyQ82yzH+xarR4BNZ+3FBIaNfxzkY
LOAe1pJAogzQYT4GQ4gGEonTzHgNPlC/Hj2OeBGNMw68dfRgtwFmv7f6dDRNCmMX
fvWdETXAzxTb8ntpcPOmdMiBK3Jy1e9plyjBVzQFWsWvVzzzmnxjkeEHudo4Vm3O
iNDa1IWGTD7tNofhAP6XONuWqFFLbcjcVTvgNMJPbLQtGK4D9OlhhkK5rn9KScaE
5TFpk5p4IdHm9fAU1iREIQ6IAWjTdUzQn2cweC4hmkkXXmIDS4DwroOHMUVsWE/M
`protect END_PROTECTED
