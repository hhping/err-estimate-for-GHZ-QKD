`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IcFOzTiAM+dN+YNkZuu6GkuX5//CFFKTerh+qtrz7zRkG5z5LHgOIf5nh44T3p2W
6tV2A87V2+Xf9SYrBvm8dXwARtDKrHvfXK5CMwcTXH4F9Zk4swU2Heau9nesdln4
4gxm4Qk+FBGlalo6/tkWkWhc7EYx3gAS5809GnzSQpcCCnS6SGIw7RNEWauoqIWg
dkRctgOqOAl1cBa29WZCcz0sWTOHZp3fU7EUMC3nwu1ybhGLYn2PoYPKb9uNTkWS
w2/S5+wawX5jiTVn2Hhu/ZVX0oix2YUwLI7IMNcwy/QTbBqcbqeQeQqe5+OkT6zv
7/TQvEVqUdnY+pB6/gCGZYtrSBBLGcuxH95Bp1c0sHc1lW9b971pyvB4IWg5YOxS
WlDcR61G24kVXXvZRxXbl5z4hVTyiMsIF2FVuh5wRs6Fp29eovEzPv+xVH9bv5+v
tWm0hp640aeWGAX/Gyuc+O6knRh1gtOnwVKr+NEblnZPKpt8fVJXFv+3Io2Vg004
`protect END_PROTECTED
