`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nj/abVceIdHqvYbLWZa7RZUoY6UiNE0aP1LVTVlfM9VgpCABJnwLImVzgg+TtTN9
z++rbw/5ND13v11K4Gnjt2rddL3sXxA3wDutEAab63fr6ELDg8o+4WyWtEB5Z0bF
wCqHSfiFUD7NiY3+V2ky0dy6quxV9UJ8O+1g1U0XlSfXcQvJulHMi7gPdN70QmF1
W1nIb+NdOEQaUY+0fHx6JgEBpDPoUraHP2Fp6oRHD817dzYP2EnKUJmqdUR4PujE
CrXiCUNCHxbOb3bcPNiKseX546SRwEJHud2DV27rDw1aNTgujR2/Z9aQhAXAn53G
uGVyoT6s75z7peY/Muz0pBHJKZlsmVYsaf2nLoUuSsWeo41KjGTnbHfmLMn3lgo7
TaFdiHS17TJy9uG78qgUVGVwYfLvH7cxUC+VEub8v2iYNRa6N+Hjpd3ArdfegP5V
j9Bmful1i8RtEZ6n1nRQxlFy0Volt6TthbfbuZ6YyKR8EES9/pBDVrLtWFULa6Ya
hQJcAYxbs/+Yy6XbIFjTekbylCsIXpWIGlS/wPFyclxR7+N+T5g/CS0XrOB/D1Cp
Pxl/JEqieNdIXzPaT2UqJ8VHqIgw0gzaXf8Q/PXLsQrVC9tCrM2hn3FMVfFAZcrv
RmBStnBD72cYukMFvPdEzEJg2pbx9Zx4knjpLKDBVO20cu0SmvjcmAZlfd473vR5
tuV0e+jdGnvdnb4+iyV3upwJftBIGkh+uyZTuE2ZYRa4ClyMIoaS67PcbPGj8qUd
wzP3oRvYHuDaZ68YfbfkJ2qF6xIWR4ziW7o3X/puGGTFjbow15IqF0ElA7AgdIPn
z1gEbuink00Et0An7qCeClnB3HyC6CrIJNx28OtOFyDgNwUz+n+5V2pBPKnKkOHh
6gRWfjVwLzkaaWVjWRvXfw==
`protect END_PROTECTED
