`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m2IF8plSSegI4P8RzwO8v6OKZQalNWR9URX6ah55CIVz7MksLUhjuCUuKjXVqgJW
GaqZQh3VjRXVaQU7ocuTXt2y2Vt4VxgBo+PjwAKjLHjrdxw2kpNH6RxuYdHT8TEa
Dq1shuNvxh/Vgp9DHFYjsEYekExgIgQQznJ9iQkOvDj7KxNBNXAWysbzfnh7j6Bh
G7+qt91TuY1D8rdZWKjIOTvs+xHv/30Y0g9Oe6JrIRVjv0eVY9UYNe2PN2tZ7poR
qekqmlRQGjzDneeGnzCA1R+7sEOTRj/rMXO7l+GnOSjbS8I4aNMsMoVWrc6WWpsa
WdgEkOvpKgZbo/TbujOlVXZgH5FX/BbiqJqHCPHDTV67ixZZNY8jDnWgUhIJq+pr
4spOLR1s6h+6cmQDoMt5qpxV9H+X3HC/XZRpkS5q9Ix6y8RPsYaoRXxJWKeh4aIJ
RA5NWPtCZ6OpUlKpgBWREN2zxZD5L6jpT/6DCF+3uEexrveoh+2NC+plCEyE1MlI
X+6gLb5N5E6KZH09T9Hn9cTbB3i1IuMXPlqIPygl6LWk7q7BNNYPp15FYl5DoK47
FURmNmlQASHG/qtkhrTjNxMbUKFztyyW4CeGlXtCD4wPk2n0qnOI/a+MaQw4c48j
+/zdexUmLl8ur5FCStZykM+2hJGntU2fx332Gz4/NvXjRcSybXBufg5jDDAq6AYT
lLH1pB10DfM4EOo0zd6UDb2CwIWQYUSekK3AJwPpP9Av8hdt0RcnZvbuI+Fz7KkY
tvkzioOuY4z4XiAtjz6WOpF9I1qUtAusQ5bMmgyPU7ebOebsQhGPHNbfNQuf0YbV
NO/93VB0fEYAKOSfsKL//D93L52wcIvfN7BuzKjwqtYdZdr/XEHuN8fGiDyerkZf
`protect END_PROTECTED
