`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BATR1Cmmljp3KpacT+uE9S+KPHo8d7Wk0/j4VvXZo7wQbPMcdcoh76n8FOxjjYNc
NzlljAy6Us0oFXzJcTzEH/RjGewraOn0cx4SrvRBKmJr7q7sNDOYXu6JNLXYXkNE
OuoDnIcTmDYRFR9a5yFpGmjjG+aGYZCiDjnKGXAcPY9u7+ZJgJ7R9hoSdA4qqrJ3
gVjX6zyniAKKITH0AxENMiJyicDTRPKAR6fymKOib/On0TJ9c1NV2iEPJnIjTKUY
irGCrtBYKbxDDdGxzwG+3anUHmreqAtzRhd2DI3OfLS5Ci23ryhSLHPSafv/2f29
NJ53QFe+EaHtFgDZnYrwmk3D4Mmr97zoFEqOU/j6ZDD3YBmWn1/M6E+PBC1w2voh
Nw8YG65B+SULD9LmPnCYwJt4rn3MLVwucNFOKVxQjQvIMO0G/lXrvyEkusEtBd8x
sQL5uxxvTurfQkxDM4vd0/OkI9GNZq98k5I6xC8VmeuT5U+1BjOEk1Q5lctz/3Ui
tb9tAUQtll+KS2bmxHwSXMJHBDzI70/zDEWHqoNVwdBz4XVcDYdHrxCpNv21GTgo
ach/BFPsIcHBdALUwRff41nt3LEWZhX2HvT14b4BMbcilQcc4ZWdUsfYlJXaQsVB
oBz2NUbGtmBHoYsnVaRyV9FfcOky19KPSc6CeeYReuVPaf5/zZ4iurgMoaJiOIeM
Dj63Ojr/8TITVOG1EeSVwOs4l9fSAggOEBTkVWE/Jy3XZvzSyLuwYMNAT3RpTy3W
cMvPkT0ccwnp/t/R9x9PeQmlR0mUAq7SVAgVuwZ3LG9lKPeVEzSEYGFtpxanGkWr
`protect END_PROTECTED
