`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q+RzScAdbWcMpRynBStn9NKUZdnUrfs6qkxjKVmorZ1O0ASda+R3Z1v1xh4aegvc
SWSKE2Ys4WbohgGNuKjcc59irBozXJJOurj2+bt1hoP7kk3smtAOfqfeHvE/LK53
23sIQ5AhsPkPkZFmPjGX4W/5v+n+w0nwfSlsEK2+Gxlz0Ywq+TyeZ7F3Euurw5Ce
3kK2jwdHviU3Q5xihb360AG0Dt5/tRq/XP5n76BUUWtYDyQVLt3AWGNytl/f5cOx
Ud8LnIAS+v9l9sBqVAFcsdf7fCyyabfbsw9w/Lb69mPEMNxN5RGxTAs9aqmO84zs
kDotc/KTwtj0hJRQsb3DFo8/oj1mJ6IBT15JYAz3SUvd+B7LK7V0q6aiG+zrziqD
Ck7LSwK+gjH/ClnheaRrfDOauUZBE9h6038PwZtaYvbZj75eqNswkrtqX11iPwex
pZNdJnhHtjQPFk4GgLVcXG+xRwQ89zo6WaRygHlK6y3e6P2HbrQILLwX3zyWvsIZ
LBQEnvvzgm51Fos0URrqmwX4IgH7S1gDGiI9sNRaFsDJx06426NToW8kkBFWX6XP
HFXwAToVMJFTRiJCmpq+x2oq/Gr5MAofLeoyFEp1Gh8XDyQny7o/F+qf+yfptGQM
IhNRBMKbFm6/7XmAeLDmir2ECj3OBLNv6i2D0prGOn7aD1m7I7HFru236yeODx1L
maMzXux+oBx0dIL+WyderfpuXgTT6HHFeHv4dPyjtO0/vXnWjWTIyamtboQ+Suiu
+249Ygi1iCpWYGFVXvxLQHoND9SaXKAbIC2YdWb5y2w=
`protect END_PROTECTED
