`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I2SBvxirvhzAKC3ih9Qde7yvCqSf8Rk+gto4N2/jyjU3Fdc+HR6s47hRbYFkKNrv
z7fey+qpFhY+QId592ZYyKKbZVlDuJnYvBOZJwYU+ttrNQOPv7rZiGRTLpL+SLm8
pxOqvI1Au34LX/9NyA1connn0+YIX+v+auYSE8DIaT1owl8ZMw9RMNCOP9kDUnOK
kkXTrTrl/khyAfFtMy2Iq/drFhobbF8J/ky70WAxHirAnrH8e++0MFeA3f0sIolg
t11MRqcQAYEq1rKhMbgqCBG9JQGb9Rmx6aKJpmVM/fYYwnHv+O3nRAG1zj2qNTu5
Sm1x38VYIussC6yojUGYBUmU3hlDlmVtw/T2Kca+Yp4=
`protect END_PROTECTED
