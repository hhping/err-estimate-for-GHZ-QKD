`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
85AW7X7NVXyYh5Cwyhcj6+1doMIEmnNVthEfK5bPO4bHskv9PIsmfZgXedW7CBan
asL5Ge3s6YTFdxnbrMIGfdHZ3zWiTBtNI3JnuxbWPRMwDetEQRNhodi487VluXqQ
kDnUFipAroRbDZutYDF2x/9mR+yUExPWurpWo9sC89Bsn6ziNULnDoFmqIN67E94
pUNI46zDJgMBGaDeOVxfZjUibs6u5fRbFT5Zl0RO3+ujh3IX1pynMJndyEFpiLwe
FZJ4lVxVWn+WIx+nXURXhRByVs3iq3UHK4IF5aMWTAu67Tu4JwmYZ3db8YxJzlXS
1yTfHV+Gr4XAyb66v6AEg5sM5ATN8B4ooobHPjLVp90OCdGMaYrDA5gne1FDqpKX
VPpreQdl1u0QczEOfUPn9vrBTHjY1svjZjGavfgx45NKiXgeZma0RCuVOnmbcU1J
86shQgsbBIP0i55xabm37RDopzb5fUUAUlrog2KlgrascnwvX01S/7n8L5Aka5Sh
C9HTBr6wWHZ1ERki8+uxOfavDLXJMedEYt89Ko1To+V4DW0Xr5M3uvamYUaBkcMr
JOGNo78EK9SoeEeOLyPZOtor15VQz8p0ltfsLp025cFBhpZZsrnhcZJScfhpXbYX
ofHaJA7MwAPtZkxXJkpue/Fw/GIfwLY3fydS/O0jM7LKKTbMkw+ONpG9Wy/InHu7
`protect END_PROTECTED
