`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q+sSDEzOX5K3aPGaOK0vX185OuhhsvdDS0/OxrnAS/c3Sa3ktDjb7zOqXB39TOKc
vwd/wgK9XsRASrCJYeRNZ5gfxbEkcEHm7xo076quVQyn3PgcndUXLk57jMXb79oo
TOeKT8uronv3X8YU3vVk70k21+SWsHgOLZUs2t6MoAmd8w5LlMeP3M3gY4B5qE4D
zaSp4pI6eNWuhL0RQQo2opd+3QMSMEf6l8InIj/8mtaevD/PnPsqJo8P05vbCmeK
VcqwMVyeNf9kz5qnx1hzBCLWi+J8cT0gqr/sLPf9TEe+B9SU24IBvLOxWMuHF2+O
L0yFIU3K0e2caxKBL6EAxc1bUDYyyS1UQ4+w5lM++18Tw2YNSdKm+OzNti9etYwF
29DgZDGypS59Rk3IwZCfWLt461W14/zSbI5E6YmTF4pQh1qg3HclmKPuM7/6PZ5G
/uCQaqGJmzh1EMQfktvcI6Ew2lFf3d17IORlmGfNb2FljfatU0DGmf4pGvQk0rfV
qFZqUTtOEwaEU7SK5lULOpzZj/ah5myf4bRGHo96H0BhrabQncugXYvxzMUJ4kuK
AamwXh1slXF3r4lw5xvXnTVbOCP+njHrXA1roe9Olhc+rrLIvTKv5Fy3brwE7oef
dgvohDg7Ija2D+huVBYOgbG5ZWbefvW/hBIquRzf77VnZdkjnE0qaoQ+o6itm7hz
x8m5YLY8SdeX6G+sL/WICg+OirZnk+dmjDgrs75G/Xm7GvVP17QWvwTEKOEz/Z4r
o55XAV5BCuds6RYEnaf892vgx9IW6pjUN62dYb+0aRjE8uYaW+uVx81zwnCARGqh
qMqE9VpBjth36vPokhHnP+ITONlAuW6RaCYe1+4dsV5f4xc0TXPDLPrbHRgVKfAJ
tGZI1Zk5pKxMyXbbapqBwYgyZzIHM/TXYYzZpwi7gXDtsiLl9+BJTpvh7nRg84YI
sf338XD7tNAI0Rhk+uTxXDhMTR+SNk4wxZjR8tbD7xVPP67UlbSLz8GyFSgWasXw
Xo+9RrAPXYqS9uBU5QWRXRw5Y2zQJm6FK2WvRbdvTX0HiKm438IAloC+3ulYGxNQ
WtN5X2CkbhLDP92vex8/xsI1I47TlH0pa0neht0ioG4bL/gXp15GDBALVzUTMJFy
AlmpB73ouPAkCcQTx6VhMY1WybHa6r/slqcNovOaakrvNU23TyRr7T7qrXf1g3I0
mzYFBuFa7fCk9nE06+22XTdUv8IqhGYKv2/C7iKGjAKgVu2slPvqqYvcl6hVGxNR
OyNxIdwfTZUpKnD5qXbMyL8I+ZKSnFWNKJ3Y6OFxUj9chcG0u7sFkLAlfgQ+qF1V
i5AdyXGErjb7ggYoWNh9QeAWY1Ijtk5Ha+iE0wBK0mFv9yHZNou8CO9ypZztHhBS
3FxYi7xAQ7uWjmjty+MVIQCERKmq0KG+B9xiLrvn3P0P1aHOJ1MFLSOW1A91U/Am
ox2rx6KQJkuB3aovm5oaYrbh/i6dYQ/+1DCyicHZHU6+Vbr67La1XooyRExPhwjw
mCZxGHc30Js4Ajnic7qydIfbQtboJjF39Rt8bDDUNy5DkpJIqUF8dg5Tk+kFqFhq
7C/+z7NU4Lv9jAm8WAXAn/rMrmQUJC72GaeFA8/VgYV5yoXHwPbMpj1+vq5rMU09
MQi2roJkLt4ormKZoPJ2fubC0mJ2IzChPNFAAmHNuBLtpd1bqRsoPyIrZGLjgU4i
Uh8Sj56EbTkXfFlOKZBZxkR46FM22hwx+pE2mn45N0Gc+5Za4kUzC8bD7kuZdVGA
c1XcpBQ+1q8GDdSITMicnp0kiW9osU5e49X3GnZkYOQHjMd7i/shjVn0KHCaZYVC
+BqRRNxQ/vzL+aBkvJdRjzqH7YyL148IqNF+ugQOUU278VYLIZVswRyvryYhswK9
yIppxJhR0rbePJ6Z5g6Y229H7YrJdqxS+09a0RDkfwRsmZxQyHvwQtj8QeGQy6if
asauNJBkYhGzZ0d+iAhjoAxoshDbhi69GekgA51gKFZIAIPSnAELxuvqunmGMANs
irb/3XBQ+nIho4q0rbwR/WrUyIkQ6apHtwwOEyn24yPMeItCqo2JnjrH4WqjnmQQ
e+IJoVmAumdgSTJWJ7/HW6Ytgt3+DpeQrXeQ9iFEvYJUxWfS8eImv71GNiaip/n/
CbVgliKnGB+csfVxTZ4YlVtc/Gr1oe0UIHskmFHn+mSqjwlrQgsQ5KvO28LID0k6
RA/5ACldswBi9e0pPd+uZp54dLv6+IXI8CXlrFYGR4+C9Vr/KC+Li4NYA+dgBmMk
7tRv4mo2ViBxV7M47z2urfnZ8YZ/As4BjpmHKqh8f2IQ+I3zjgNyvENzECSiDfjY
SXVw1MFDGn7v8ynkBSE/Tt1jKAlBuhPEN8Sqyyo76FBJIfh/a/D3F5q3cjo7zozU
Gk+LyDnGRPqNUOykY5gbcI4CG8cs4hiZ7i/lY9VQdIXz/fcKTuOBoxs2Qg8ryiIy
Cy4jyrFACiwqBlSXra3JG5bbJ+Fd3DP6H1bY91dN+LMFlxeLJYX5tG4OspifPfCZ
v6hdmVecLzwq6+6iSFbVpSp7pJSJYEz8i0/hRiH+A5siBdpvPYPCsbux1li54lhZ
Ug/Gd6n9RpLF8Fqd6BdtQYbNH7LTtchW/EFccaZB/5mOdZatOk+uYWIoQJZxUPf8
VDI3LhCrvxwN+Py8kTl9l4QmyA3G5Q4xHjEDtNrQIXGzGcypBJAbSqFJgvekc7Q5
hTSiRgNAuu47GTOo4IXBEzaxOXJ8woYXeql+v8pmNkm0c4whF/lPNQ1KZBb8vjv8
95//+0rulQ9XE3NXmd6f8DD9NJKC0eRoGEdZVVQZ9VCzDDNwDjzSDSXceagXWLKN
aLfBZcFM2E29P18L58oZe15YGPplHUVn3Uf0Qt8FuFSZOKyhuDmlhaqFNMt8ZEuk
m2AHax/sKHjM/WBB5eikEE2LYwE+Inx+5yzBZyomeeROFjnVC4bC5Gbx2AFSYUlO
zOlVmmC0D/x63q3ysZ7ndZLLbbysOgMLX/DLgCWua2YUOukKudH73+ohWLIX0wxL
21Iw4Cl4Ss+KapAahPiDp3FFrWxFbZ3EPhETkPb4VJ55CrJGfQyXDz8rYg7KnrgO
2HLvNEHfZ9Z0VDCuhF7eFoJQ8b+o2KCJ1V86utqhm85o1Qnw9khFn+Jiiu0ynZ6s
NXtU8gmXiIwLoqgQP0z+vfHLkxtD+ly1fcsttwlwUxnM0XEa/L3yhvrly3Pq0ArV
jhooAo1Ew1yqJ8aB4FYlWlU72gV73degaybN0UbZrZv6Zq05G4smlN8HAbyQEDsc
/83lIpSAk5HsWYCi+d86NxxUu+UjO99V47fg9ELpcIbLaXSZ2xbROuAthoEiSY8Y
V4azwQf3Tgj1oFQBK8LQiYwXsh1zhSDhGrUkFTcPRd7W9NdUB4ICf6XGvLyEQBK3
7/Y5cH5aifXxsW1OtgH9lnwCrDIvs4rTQgxn8jKrM9YltlNf8hwMv3z7Os47HUup
oNw1fKnLBCEjH0sd3URp+lEIaUcLTYcZb8cMnjgdXJNdMk9OlFiyI8I5HO6BYY3M
lQqLP58h2eg5jaZ+kle2qpg7STroSPVFEI92tfDDHjWbdKGLaNnfpi/n4Er2/p28
OWiwwBTg0X/KF+IZTPPkbwsD17QeCnjlFBcKjHqRmEOctm4D8nzzMsK7JsamnLOQ
jAqIA/OqSlv9DuZaVScxQn3qav29PEiijubFnXQLEjdr6P3CkVIQ8sZ4qmzO418M
ZxFyamvJfoFzEZ+3K8hjPAJ5eX8pFJOyYZd1SZzoNGmVoIGaAqk2ttwwA0QGNKdg
r0VM+1e4vZwAJFUwBIRcGWUyvWkoQvf8aRymzF5NExE7K7Pj/qX9q1upQy9/+84d
Dn4ZqSKRl8FIRuldpwrNgNI0P8xH71gwzPxFGnYn3mFF0So3DWr0epK9lS0DLUHF
ZAiSMdz51SthqZCPQrlNATXgo/OAqtYkhQhUXINR+IZLg84ero0KBiCKPvqoDmyc
4y9ZIRomXtUv0Z5cXn1PajvSWiTW3sOgaH/itdvpw3aI4vqBIDt8DHiTbEp0Ytau
gNSzYlTY959vx/EAWjwtwJtozxUEpFmaDsdqn2uy5OeyYbQKXGynqobDeOElrMts
CqbuhNDQaUOdjHKoc0s+Gv61UT4ifb9dwb9qyAZ9R9gOIRruxMDHj+DPSe/foQws
V80Prn+rIr9GSz+n0ML/MbnkzkTsZIrWtMplTlEk8QnlZojGOyMIFyJdqJyAT6LB
wYSAzUQTQdq9v46uZXhozSw+Wiqm4dvt6ehfhpeq1Cu9cj+j6h6Kfba9GDXe7+4r
WH0Jf4MVh5unQNOQQOxr2wKzgtM/dky862tDZ3SINyGCUQYx5TrpVv3zvglIG6ZM
r1gcG0nDHob4zxZR3fXsRMyBavfABV+hKCp7afId9Tw6imiosVxDawgoK0+oYO+Z
WEhgqLZuqYlPYTFhG0QSpDDxBi467G+pKJWItL5sH3lM/BYlGuVH85lY7AVFYjyo
atfdgopx0Q4Qt2nuewsgmNCSmo+1vqDrCAoO174eiYMCMGeiaspEfjfFk2yySLyr
onIOh1teQ8X+e2i1+XRqrCTXmYpehqxd9GlpKF0Zji0oHvxWlVLLDPbUZc0zeNWo
iVWl8Y7gccSC9p+ACS25cHeQ1SpbX0IFH9HzU2+ycLJy4NQAgKJEdiyYI1jNvn17
eTstY30SsvP+iW9LughNYBiFQhQ7xaL/id2oFksXuqPaSt/IFVlgjO4cu1LUWvzJ
P/rMl+RJIiow7b0dskSOTDH+Ay5P/JNgNRxrhvykbKJ329fAgW+X6KwULgeDKhPh
9DK2qwXOMEn9qOycTWBR5xPylf460/oUdOUP99gR8OMUW5QAq5BC/sMDdD27oVUM
jMqnBkCMc2148pBAEeV99SFCXUuEyTNqBWJ7/kIEuhEgFLlkAj9AwX3snXG+a+7N
XhaK2zGQ2oIIsQVLuBO4n16QdrScTPGM+2slZmSoEy++B65tEJLZXNu6dkq4MXGb
HGZoWBCVkbyLcPDMdrqk9OVBGggJMPB0Doj0wjdAsl//bsB6wT/UyG1iL4Y7xogw
PgfU2Iy/QTzphUPNKUUMX5nJ43uBjDerUVx0ds1oPZwTxC/V8Qe7qTI8XhetbY8m
tvXwI7EQtxTLyI4M6ryA4dHi4bmdy7yEeY5DtqYyONf2wngCP0ahzMe+YpUTfjDn
yTjoPUTbtAs0r7QVveIQS0SOlPNjwkSSSJXf691iZHMl2eyuW9ILxIJwMflingSh
xf9oMzJ36etndYpM3Sdke+kUQ7Pz0pte0rivL1TRDBtrp66rOyvFWx2h/jc2I7aj
hX4VZZEpgHN9Lyx+CNDWJpxGRGarZcvdDbFdKbLa1pLEMgQriZlMRZOjfEzmJF/c
o8nLcowxq5dBrNGo+Id02x2Q9GG7csHzsJzmNXcwcV5aVEus0xSqZQtUsMxV8G9S
L7CuKEZTNbWCssRPxTyqV8CVxjIWfu6oogQMNTmE5p2wQaFZpK8sRu3UphLoQC/a
V1+SPcd1PK6nKgZfO/XX8zqzs5NFnZmqrPc+6IQXyiyUOlyDcNmaTyF/wTCW8OSp
`protect END_PROTECTED
