`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TZoBcp693qz3hsn5iCkz+Z+ILSwxyMpgbysEry9UMsZCnxCL6GWheqGZEWJbYL1w
nG3IGadGi0m8PDn+BZMn7vpDTfckuD3iuxTeu98BuQ1hFw3XnuNpWvViurV/WWLI
4Xorz6uQrMcS19OJgjVh/oW3kAARk24X1U4IASr92J0rpbzhNdfTtRaEvto19KXo
do1wQpOh2eo6z9/vvLOb91wa7Or3apVib9BOP/XPncNWuPf9vWmQh7vLLwhdz8Ef
mK2rbYMDl+DQRiOrnNyhiYZMkgzdbJ2hkDi6KX9wKvVnIkD4H37F8+fGTNx+aQab
9bngJYXF/7el6hcqoTOTvmNsGez5wJfLOw05pYqlN1DGLS8QXuaVKPpcz4KCHd+b
y+iOmHmZY2gSuGYMyGK/drZOz+Y971esLfnvQ6nchfr98tZa3L/PyCOben8jMzwt
9qVjZ7nC27AotckgwvDgOC37z4swJNno05+91ansyBXLi0xz8wjHeRfIMZr/z2xX
SGM1v/6bLvzI7/cCAxsVJ4V+l7YmZROek4nbQNfPnepzk7NAw8PJY2OkBLxWaZ1m
D66KwS/uGMMEBDfjVe6+DjJzPiGFsoPNt05bx7KazzgTw9AxxE4BdqOPDorSkmH/
CE5E0oLrpCBHwhm7hlXwNMZdO+HrLhU3QoDQFzFcx77MDjl11w4eJe05QfRPxqEV
bZrBDltyjZehyqRMwRiilflGEic4/sS309il00rKiYe4Fsymw1KeJfK7IAUeK2ld
G5u7AokQsCrwXuAJBgVnhWP6wsTld8pr3xpSa5JGxhM7uKsIpkjOl/Uz58/Gi1an
pbaazz1fiS26+7FXf2rRq6WQl+2qe7cGl2s+ojZWOQJ9sro7S0BEUcAPXIxJfvj3
BNA2M78zmRsnsvMDwjAtIYOyKOKxH3Vo1kOiy0ksIFtA4CHV7C6m1tmyoC67QB3c
Zq5iO4DWhEX9CLxaGpsTcR/C48ZXnxN9R7ho1avoxYPL7qyHjjhAdH478P7GZ4jo
wP04vToFpBjbcWwPYsbBXwss7T/jqyTAJWoxbcFMBS299PVfS43uPr35X2L9ep+N
WvY0iMVGXi3CDLlsfMfQ+NWwgKIgLCxoho+QOKDuGHQXURNa87tkWvQXfCllIsPE
l7ymTS4eiCimLO1e2/bFBT+U2/BfvoIGeptqbsgpl3BBjB/KQ3kH7Z+xhQr8hg4k
RuE3Lx2MoVDoOmzx2mOhVARexXidxqcmZeMPeaI+Aa3p8r94tvOHuwsbzGPo8w3y
K5Cmm3o8/g/LSZPxQ8E7GEMXj0lwIofmzV132g2U3EREs6dYNlP+a2+p8pSC3B+r
8Kyerm4YGEB3g70WCN4JIXnT+9Geql+OAbim7Edw5A8IWGdmvaJked2ma8YiQJ+g
IHwXR3pLen2FHateIpBW+jChbvMA7OCfcdbaUoFaaOezto+JfYFfQ1sRO4vuRUG3
bfyZFqg+Xz0oZbdTnM4g2DESoTTYgcGnwAuF8wHi095XWUcIU8ErtFw4E1QX0zka
CMQ9yV+WnPkggfPYVVGAkbGKDiVP89pmEy4QRXV373ktAxaA0QGAjuyXB9/6ngsO
pZZCtaCYwtyXU/E1fuCAgLw000FcV2UXN4tEnZyEqk9CjcY3DElFncwMYaWdb5Br
gAR9/bgrbka9uOMwy67l4DYZgAnQaDsMPxcBrCX4MiIzjjtTlrSzfXQX83e0h3M7
/Jdw6hEaxDRrJWLm22yxADbXlH5eD+zjNHi+amsBoEZfGirdkB/VnfiznaNegKI6
sqN8mw3mUMn9h7Uc8h25TL7f9gtx4N0w+Fhqk+q5WJKhop9JvfrFY2Y0AZSWHqwt
JYHp8XOKUWIq+Z706Ib9JUeiU15aabeEFxQZVWbTHAJTvo9i0nDs8cdPiI1Mr9Vd
+l0Ma6qq9gwgFW8kH3xH0Q4up2lUwhl0ywobrMF47jdQU1setNxhxfdblqY7lOC7
`protect END_PROTECTED
