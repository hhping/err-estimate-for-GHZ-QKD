`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KyNCVzJqjtWFSTKq6P4+Us+sZCTfcHDTSxQvQwlvDyAYtTsCWtgsoJB6Go6sw+x/
UF4H/6N2H6aojIPwMj08XNoQS5L4DEIirfN4nl5WlP5Kfp+qXqF2iezN4QfXpdIG
SbxnXwkDiA0CCH15wJCgvMxEZhOIffw0hbYfu4f6b0NP5Fgp9W4NzCEmEbUqRvh3
9JivWoeiEx0eiVdvbzP2gioW6KuqidP3aJtEjabe2loR6O/UAIBwE6Ub3SMW+Cje
p8ObrB+CHLYHrCZV4zSjJtz440Lu6n2e/T5ftr7UKPyoKdKHPFZEYwS0FUPKtGQf
+7o3wvyfG/RTWh3KRfWKPVtRAL1+ib8+700dOvqbCyiSZ+3xGG0y0+2+3SzsPdqe
sM4sGrT5WPqECN1ttxdXrQ==
`protect END_PROTECTED
