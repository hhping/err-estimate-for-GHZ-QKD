`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KW3m14mkTLRyZVFQBzbjKG+MrRIn22wLZOeMBrqQ8bQWdC0zmg1NYwmsHlXmcoGq
rrMG6dXHeBlq3OqLZxXuGQ8ufKRB8J7WF/1G3bd5jX8GU2LchLaHycoAzeMfo2N1
RT+XoUhGsoKUv6+WdXy/HWqCUljxONXwHSdJOdmemOLc9HmPSNR/uCEHGsEEL0/7
6eN9DG0qkAgYRofttDQ8fCLfQ9qDwn0ZjOI+1O0EvmwdtT1mu103uN32+a919tKb
xHODuEz6l7mr6PEPDHpNNrE8iJEBWgHplygB1Zl0a/CFBi8TbD270qegjwUtVHwE
80BzyyhG0yz9Suxi6qrjrblgcAYSUMi8YGBlhcYct0bLAfiK9yAAY/wGwWFjzByQ
77keK1XB/C5NlR3xtOeuR3xADz1dEgzmtUxEbKJW2k+q/AGeqcd5clj/q5RY218W
AwWJ+HuQcFHqRFvLVmPqpTzKPATy9Zla4qoq+W5vI6qo/uRyZm5wUzDzdA9FdIBz
py1wBuIufu+46wLTCz9LdpY64IA/THHxAUOHJGK36vLTh6yWxXk9UV7IXkmmDnun
ywoVlZx5URMH3dWrC7D41fFmymzX00/LOXo3JlOBAoMc2ANpxAICtfXhE0pIdI3W
gfbvUnzTM2siUp+ekSCwu82rx5BkjotgkYReIrRFoQA=
`protect END_PROTECTED
