`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z8rsB+Kl3ukgxXS7J5GKrb3QJtl5SdRCZk66PK8bita8oY3T5QCYnaO8cgq5jtyO
kvHhSiR5x6s4Vgez/nxqJncldFezM57gaf0lh3kiB/MmRE737xn4xTRnHrtlNOSf
XmwJMrRWExt8HmGuf3Ib+NfawB0tcu96gEjyM1h1QFKzjkFBXEVHWR9R+GZ0W04Z
VfTPfr3IsGaMVldsuv74nNDODuqR3J0fgggHd2Nfb2lZfOkIf5vaKUuUo8EhkJRh
THR1hNENde70e0++/sC/vkMabncY/90D6KCl8LoZA0YnP1MKR9NM0Ia+OpZHp+D7
V0YZc/D8vPB7awoqSv1tjEmimUsP/0ztxrowr2k8fLQMXlQLgyxkoVmNWqGN5fKT
PYmtZlIEBQXXjzD7HwURBhS7QnolRjXKjW1GH4zO09/a5INaZPi1nR8IHxBWWsRP
AAGRCkLf/ystmXo8px5uTU9pKgAeXccgphLm//vCNHukMAvUd+zlp/KhLLa7Rhu8
Q53jPa33rdVcqg3blaybzSpKdSZdfDzJ4WDYoEHrK4GX0OXUYPNrnnlHuYaxdlxX
07va2sN54buwUDoc7IB7pCbJsjID/v8iFr7WXeY/VAjJxhzhGSkyeWAcUHqlCP/e
wLOo5D2MRfCWtbC1Vv1o9hNJYSu6rXc3PmhPTbBckqV8iZtUE/ECqbvW8kQMCSu9
VTChmb1wGxNHYVykV/Vs+lDCbwM8FofoJdnRrQqvEyzhiTP6/s+1DExejVfMa9wZ
SnBL9KXGW5Y1mGVByFC2O07rZhRLtuuliLBDYtUjveIsvvaPWYFCHsZsP0pm8Wi/
ATuYA6F951K3yo5eD7wR84F970EQIVrXnBi2+/v5n2BXP+LPzf6HVcOABHFz5Xw9
99xp0+XkDE4gOnPg69haLnzXbuNIe/ifhHwKxQL9dbdXBhsoFFIOUwj3NoTBHn3B
08H56ENs7Pbfd1zf3472r6Am2aExg9BbGPc/szIFeNfx1iD3AW9hfATH+bnzaS06
Gl9qCUZXWgPsyD2YzoFn4QvD4tVN4d/XEEnghRLBU2lTUX982QL6nDvLdxgRkf9O
YMGFEoiXHQQNoWNDLHWYHKU8oQXx9NLUWoc+okWkNHll2h/gspokifM8DevtYN0J
1zaeuKMzSH9S+SgYRAWP/4a1pO9KmtRaK0xC6YgblSLdQa4gxclQYeg9N6sydaIK
VbhIUxkK6gNFxGJ0tlXVQgA2mP7nT1l/+GCBQhRkzT0Of0zqbD5/PlbxUOzNkUlV
60KhhxiSUfr0GBwH7Fu+0gfA/6cD4yWMVSdIA5hcdRPlKDEFtuz7idtqV9yQbOSI
/F0QGHEuGCSA2cYDW6Pe8xHu8+Cmalg0kfp3kKeKsdfd6whXfJuGXzCBl1mzs5yD
8EQrzXw5Ws9HBziGtTZL7yt2F/22WgXWbDdHgEwy2tDEXcylsaBCI7o186TIFSb7
pNyBrPY5mzOHJOtkaj7H33aXs9Vz9irz9h2RobxK3xKQmb1Kajj8nYr25uuIMm7N
NgWP9tlccINWPFrsMW7NHzSO5SYslQRDFIEiylA9/3hmDgPbW7VZpZE6YvWj/CZZ
W42LDTUMnO7RnsPDlwQedgDulaRXegQfk/zLZ5brIB0EEJN2uWJhZVOP+aGdV19X
vzdIJH0zm58ObQuEvQOGvE5a388fSFdbUrerreUJVPa041ofplD9vAeCChYuviUg
w8khmcyXXcJCsO5YfvZ8RuzdtmK3L3iCZWAEGX1kAMDpHkDZhFUSKZbQ69S3LAAD
rgtoSS2Jr4/Wt7fCsXXpbkYmtGvujhyEmVk3rJEnizgYvadcrNfvnMrqko/E4Aeh
RjWlfRNpKtl6KXY457AgKG3pWIzqISjhvw4UzRXxXBWPQhkj/ilNrehlNavTEfh5
5tJQCtqAFh1YPhbd4T85hnUX78MG4fR1MJK9QXUh8TRT+gk++ysADf7VM1DdjS8a
ggKqgpxk1i6znxhIRF6aAAzsECowokuVvwj7voc/8pIoHt8vMqDOroe2hBT/dGgM
JetsJadITF+n4cMuv3AdjsQVy+Gk7mQd380ii4j3Q5uL1MkWYYyBqkkccBwxbHiH
5/uVlDFtlOUi37Cx8YDTwoMHwcZdkDFOManaMwQ0f4IWNZYEKs1YGjf3dQbq4C7L
6yul4H6kAAlUuB05hjFkVb5SM/SMoewVmzwUCzKxBm2wiCglcvh4baeL0NuQ4BYK
x/UajCQu3KUSmSlcAQEGwefwvfWf6OJNLFgD0BMthHTZaZy5hogqKPkRV1ZOTAGZ
GGRAi/Nw7UJvMWPXuqkj4Dq6gjicdvjput64f9oWYDdC587zrWDy5fcxdQ0/C1Jm
rDfpHwgKulLhOP8fzwyBKwvs7rK4w1U6OOTOPUzKG9LgHbZMlKnSEuaomh1ULELD
HaCVzj3XIxbKF/lbQLOwZTzZe49oxKyuFYFFGrNfmFwugXY2q6brRIsnwdn3251n
CQ1BzhQxVg6VLz45HgGdJQFTT1Qr9iZyI4/p28PQrYSC7WBENcM/WBxfQTbXguZ8
Kt/EwlTTLISc+zUA/wnvtO5MQK5QF2OXB6jqd2YOth2B7xu8V9XRAsYU4pi3tQ8o
1KdC09poYdigIpt2+GtfdCCuBXXXGvHioPg3Bj0oQRfwEBzCgXD9O1w9rWYgs9hh
D9nASyhZHww8FO54QMdcDMhLueNJcgmaSc0MIcp/81xQ44+doTvuUghSi6ivtVKA
WxXI5eekDMnXdS3s4XB2vsi8X0PS0UvB+lxEd6ACjmA0oTuJAapbGgsysO3HnZaa
AYWmzrh4+beEiD6fiwI2B28d6t7S0lAujtc0xNRLrWu1DAamvcIq3FVAqubSxatq
u9gHKJKRMJH+VZngiI0Z+2mzinL3//1tG7FLerXAt6ggRXlumzJaWAg9mAYgh8j8
RKTSz2k+pmDujzV3J8yIKGBfc5ssLJQLiQo4SIbQy/oNiAGEN6ahrkxHWfS8tvBL
pgBqxksTc5+0EmArgritN7kv796lchFg/lEo7ztqAZiQC4ydfOcZpL3etMkg1yK3
G2b08m/f5RHOWhEhpX7xNfsJad9oWj9/SFbYlRFyqadDO+emVoeqpqEEWejyZj9Q
oFV52OxMRR+hxyVxz49soqQD6LOS7va151ma9NFcFA4bSXOi2yKHaGnPM1fPEbzK
pebBZzJ5Uq11B4gtTd2stb/85p1KAYuZvXPa2sBMyoUJtjFIwy1tKF5n4PlhRfVE
FzRgmiPVAok+hqy/ytJNmj3k5DVdopzFLQ3JkaZCuge6hWPemd8gocRm9aSa4t5a
r+gsAF+t8UoRtMRbCVMGFNMSh4r1ltyyZPyXjRjep+wK5JKfHAS4d60mUthgGMAf
CwWr9Hxzno1AmgY/oqCqC3A7ZySGrBFt2PXfKgb4htnM9R5qm+lgfZRBAmT9ymO4
9FcqG7a4AiOAHkJJ0iEsbeKQKkSWt0jBwchR0ZwtkiutM1UJ4yqqyTpvpYE7xlVw
63HpDRsB5DI8PTFCkarSyiQOYNvRAmShOmrU1HQk/CUp171UuRZFLxAs9fSAkWct
pAfh1cqxB46ow/vEzyZZtK6Uo289d49eA6p9LZAxZo+wiN+KLLYRHTh9zyn/cWMT
6GG8QzKNeFHjRb4L47nBS1+iaqPBRs9K6e+DmwccPfw//GpuGcur3S8q34A5kaYi
qnK0ifXPCMPTx1mcM82nNE5sclrYbo5cZ58+e9LTOUXai6E6bbRZt3txgDL8iRVH
5r0HE/xQ8SHPJjqMJFxYH7NihziQLkFfoBRyoWt7690jt/zJtzj5Pv/hqJ0l3bOw
DM8kJK7X1H/GceOSYGjt3ppSg6Q2YJUdiYDBiaoucWv0A4t7OTniyq3zsoJpXQPc
wX7/ff1skbxfMHZIMNYnW33lkuWa+4kwLnbJktwgbKj5H6hzZ6mewqY0R+aFdgHd
SKebwqAj7s0g2dfvQkqa2IZ4YHZ0ba1UoYb6uWPNKZG+77Yn6/lfhI7eiU3tgayi
ddSPLe5MVcr1nuW4rQFHj274vlD/t1c56KxnhqU+tVYGLwg+6DQ7iudYiuko8uyE
7c/FlsYBLv3aj6hnN0V6K252rVqvF3rVIyzdEj/bhxnvWqIHAeiLavshC9UlnpLj
fb8ReQ+LGr1RYeAjE68EocMi9I4ml5m+snmyaEOBEAww/ruaOdRCPFJXdpW0S04O
92/F5MUko7QyKQ+HZwk3WQ6JQkvDgbYnh83lvU1abUkHd4zeJPdpssJJ0ntQfqKD
4MaoJR2tEhBJh+ZRqTgcwxQ/wS/kIRUohsUkQzEKUB9X9NNuWoaH+hYA7C0QO1LM
l3Q+sam9vpbPzCmHB7tiKfxo0KGngG5aAxkYV157Dc4qZK5JPmp5M+xOlDcCLvr4
RY3fYSMMhvn4JIOKU7LWj4HHw+eOiIwqq4P0q9rNeCk=
`protect END_PROTECTED
