`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pLP+ikX9TS8CBfr0oQnnVms85LIbESpDnqumKlM02kZkL750Kj/9rh34iW1CAT0j
aaf1ESrkoHOUErTAEBaUmHGAixDl191kz5vAX8SZajoBrveqbpkB6orlSOHHXJPq
gfozWhAkllgCf8tfZ/9Rm2HK9FIMuHr27E7SvBlMjc4FII9x0sO6/WEtpZJWvTXy
jfTp16OISsgp7b0yI+ql62rYB9unYmuwF5jGCVNbHA99138uRtRMW1b7Iz3teJ+q
f0ACKrzTHlLTWugrStFFSRuQtEdqS6o1rDenib7lNY9xGTA7J5RFUwGBI6twHLU6
ttFJxuKFBMlAnoA+xL3m0VKWWFRxt6eEB/89hLTVFgGEdG7crSjfEjz5N4Gdt0bS
e2MNXoZ6Stj0eqltct8ulA==
`protect END_PROTECTED
