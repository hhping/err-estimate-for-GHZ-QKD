`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g9UUGcTkFd2FjtHuGS36R9CBuljffVa3u+r92SdMGT3xuivTXQacIXc4FUQLQpVR
kyyocJ/ZGnphpP6VuLE2Jtm4g/UwtDt3yKk11Kw+zrA15CP4lPIx1AcXraybn4aU
HiEsrVxHspjHT6yoSItO7aIDm/9tekN9/Otk8GQPPDaaPbEHTEgg92GBtchEm5LC
dYiwfysRSBtwH4gErLH+/slBu1iqJ35VdC2oMv7Kgres6VagT4ZKSdDC2nMTzVUP
rHZ1m/SubhsPOgBbjVb7ZMOTMAb++FpQjOUBAKTtLJl8nSBexsEC68BGDiqrzg+X
73VCYMon7gG9mkpjwEsjUGLmZ7Z0Pq5KK7gjJvifUQaFeqrwBpPR8c7rePlolFMs
UoZZb+C3nF0UcRI/5fo4aB5fINoSt4NAzm0UN64/GpUR5S58XMWpRUNeKbxQQVJX
dS3jLhk6pnPOzsKbEnoFSQbX55ic0nmqC56uyNKZIA0/X8WK3u9GLVJuzO6UGSC2
wNHlG/ycGN0XCns158xcD14BSQamzQAH+7+F+rp0c+WeVESRQs4dtbk4RDkoDrDo
Bfnrm5ZQMCgUKV1KpLWflibjuGRXv+oNfzeQmL5POzfxyw1u9Y+KDiquHOpKarEK
L+CqmZb6QAJCPQL5WMrTn7VHx2cEx4cwxKkCgyvM20ShlJ/lEY2XBaMsJvMZ0KsM
ZKDXEZNdB2xdqNMqsAmYx3iFpnqje2SyQBLfy8UfhqO7yx5B2Al/olLTytkbE3Sl
Vl9+Oi8tr3JEwl+Y6HanK5+FW/k3vJRz/R90FTpSEoDRiKCwYcTZy8RhnvyYT8r5
9edDhdxmLhckIqVskWBM6gchhWwE/BvioSDcX5r/afDoQaT/RIQVPf7rLTpWPjGl
mLZEn50qhNoHqSRwkmg/l7PMziwaUIwrDGCtnmw3aRxgsD+WUwK6GkhxqIHjUvNx
Q/zpdT+i+omomrg3efbRmQtzLZfXF5qq+5C0KfJTaqz81u9W/lUX4nn2K/x5DUrX
J9rWewZDtx5j61GxOBtAZTdRNE4Zimx1pU5kyIXBBIC9FBGWYBd+uTb2klJyIeuP
Y06R4lo0uTPFdASmDs3bW6VvMz24nh5aJ4PfG0RiuOELK5QC/aAeoFVunfkDPWxU
YXXiVMrIOxAHyvPLB1h9A+ARJl/fs0fCMktlRmCSxbYreol4erUZI+n4hUiKDekL
Ie2VwnBKWeFlU5zzdD9Eup1yuN7mZ18eWh7x/W3NuSl1C7nfdVXVDojzfQVf7V6D
pYak0jv/k2jO/fVEwVHNBxawvSAUzxY7vNSnkfd8anNAXyducn6VdVSyS9DMZ/gg
Vf1Q3kIoclX2lVfw84JjmVrscVRDg8zm4ju2TOd3g7Oes+vQJZ7nYjhhUk3/V3q/
amutkjPPZEYeAKkCd62ZEYIo9i8aOCVnwAZA/4trOH1FaXtPMBW27QhDgGNQ1eax
gEKNyz6IYvfuekcDmfNvgy0M1PLYtB/SvCmiE8cC7zQvgJGNjReA7Ju1ts2SKZKV
+ztcK0JTxkY7EaCuhyhS1/fQ9FhnznkxJHA5oHy3Nkf8tHfGXhQnFAJR7ifO6vKk
D2w4KC/vmN83wmvPLD+8JzzJTPcI4UVRM2FLa3JrtxwNtppM2s7xgxvqREizNT/F
6ufGsYK/uS1xq5CvuJ9ZBre5SiE8vfFCZHCPyK3tBDy1fR9+SHX/JMshCfDG/tIN
Lb+xM8w0Ltb/V5A2D5PMQaH993NtJ5QflbfpoQhKktfDtwPEZWAXV8UyM7j6hb6+
HPIK9YaJZAre/Q0Hoj7g8b5nVM2j+Qczhbo7eAu5mf5Nv5tlUvStYE4FUzuAwlTh
IONN+xiw55SMeVxgCTr/ts3CR1/W/7CXH9mxTjB1yMaE3kLOpzYXNf0YpYVNU7fk
8GejNnQvo/IPtGx4c1VZHGWQbY4S5piM6D6z5R7xMLe0kP/AtlnYhzvAj9+0rT+X
p6TaLq3xIC2GepFsFJFLn0VRG3C3I79ssVcHwbthjPwYjdEwxIqpX7lUOXsXXDQ8
xnK817ulOPD287cGaMLUZVQf1Zqysjbn3dUy9p4TkEBKzx/YYrrxUmlBD/+Ede4S
N5q/LRPKPp249hAU/C4/NRw+3P2yazZcHHJhis0e3wLb9dUC/8pY1WDB593RVHXU
KKfDFv8ng97hjj6DhkZ2fSt7lAmiLaGtPHliWPcyZNFxxrP2SZmv9FoxJWrsqDjL
0QwAYi/Tjn0Fxjpggm88ZCFE+ysnI90ygxMR9m4XanQmIAwZIAKIftaWT6H1Tlcy
4KxgLPpbQMQYwTp32YKr4ksCNb1QBJrY/TdAc7FDCsiq0SQZkFM/XeyxQxYYvSNk
u816vxH5twNGht4kzl83Qf3U0vi4Y4lFBxRNMvfwt1k0oxpMg+Ylc0S5YcmczH/F
UMAG0kSx8gLzQBB0KDAEf+f+J6YcPGwRsSX5ybcbF8m0hjrzUR5csYW36vYMsHHH
MxmBgQ9ywkLW24ZUI5DrmodF6wSIQfEt/Mt4BlZrhauHMpPqrf1LqY2lmHg6W3/V
Pjo4TzxYiv/R9vs7Pxgx5rubqzOxr4s9QLdbZ3LFpcgxGcbJzwRwXrK4T6mp8C1L
HmjHdrQBej8RPVQY3XQDX9ft1nFM9DewJ9u4dzyzbGbi1ThIp70dHwSxjJXJHV09
LvblJai78bHaPslBeBJ4KJ1MFhlm4FBmq8hSM2cuzGyWreuWBsESphcKVQMpOEcS
9pDGgTkcYmfzrU+FGZ1RrOcggBRMVkBn4XmllscllxeD/2y9w7Pd+4AmMAMsz+GD
CG6nk6brhVappwGe1eosUhp1Iu8NKxX6OXAp3Ag/iN29Eol7NQfsiwVygDfzIIau
URVgs9d4mAVgG2JuGjVONBZIfNmp6+30vJuSGxCV7NpurNQKI3jlcdKO5XFYpQz4
m5lPFFEVgw6H8Cb+Lc2DMihp3OW6F/glwf6UIOYqeSR17m/j2LdSJ9GBdfBZYiTe
R6nh9PhFRZr7xKw2MsZZigJCLl2d/cycqQXd3u6XrkUQe8JZuqN91X060+vibhof
ROrznKEjwc11Iihx+5vR8SUnGerPO7Xa5q3IrWn3Zqujh97imEXWu+TLmbfJD/G3
8Y54CTIoDZqoTJZ+JkProCzcuV1utNLQQGyZnfzF0rB4McY3o0+nONjbfX1PvMtt
AQyOSDdjH59BESps6VIqhJcAfh8rGd87WyU9pz2P0cbTz6X5tvV1OAk8hdywW8ff
zTowqZYg/dTbVxTNSqFyNTMgOmhuDYqyEvByth/cN85mKZofEovCqeP7ONXgmVp7
WYzTRMhfijdID16VF/GZW7kd+3fnE/I6G1RT9P6TVQlD0nVqaKASSgUKOVGunSnR
NXlyo05WcKHJsrMd1P9Y4SlWHkIlat/FQX65UPsrP5QXfWmiVOaVAiNwfa8WemAO
R/00aZ/qOG//bj24mIf92lVficUjXbp1tDlOCnHe2+NF0jdrwCTwkJo360tmNzSO
i3VMfP5h5AV/JycfkKoQSNYB6i+IohPZuz27z5ap9VFOyfD5tNxPEjKS5cHF1vEw
m4XgVrHVQdvdfvPSnQpfXb+TNTuCfSAx1wDP1wlzVpkwyaHUpPsOhgJAYNHh5ts1
XVdkWWrLGiG3pLAnSyLe/btHZ2hy8vZlLzZluQsCt4YUCLhK29gTs31qUazhword
Wcrzllt1LSuo2fgsWB4m7WLYs6X14ovICTrVC2+LuKtaTwu18mbY6GTGLSrrKiyS
YuNsbT3K4yAMFhplIjfE2xtJi340R6ApF+hwJgqwzL/xJfHd1/Q98Up0JP4oFUSd
P/FEjp+7GopMXpDkyQXxCxUMPSrqYlmOMM9ASPeXTYvEKP7JnOKoqMdEYga5UeLP
6Uv7jLvblgL6Q8dUSNojDfW0HLkkwNa9zZfszLDMQNwTIEM2h0akXcXgqBJ/BFy4
E7x0eIzRQStHU+qk0ZOXom9WMRfnn2vDGAU/OwA+BxckRa2fz/FNfy4dwIBvG2uW
tWwKz8fglmIOCmWmOopQRnnjh2vuzoIO6OU9i6e+Ih72Yu7YsYdDFntbuAsDV7x9
jo/tPNbE4LMSZ/f5y3MYtCJbtIXGlO3pJburWn9R+NUd4W/y6UT8XJDq3eNEjD2f
HpSj4J6cNxJCqOQ7qr3jOjIUQo37gA/Ys0v98/8K7ZP/o57CbLrWqk3spCHYoHWd
XBTsutGWO09LHevd0HJgR0UOnMOmubEr1gll30nbc9uRJHndTBgvYSb2K9iueO0M
WbBbHI14rTS2VYX2m07LetruwPs2TT0+VKLuhxRJ10umD3DZSJMKup5vKY7jXUqV
m4yQL6re+85Sfb4weMy2fK6GUpo7yrPl+VJW5C3n4QLlcSV9jl2zFCcGmVuCHRRk
NrqqlHvuTZmsuxxofywAkgN18fN1PNYm9D173Xb93h0=
`protect END_PROTECTED
