`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sHzdGhnR87NqzefsltrwGX3+xFtKb857Z0OcAoF/4DIV0sEpDukzVpmQteBQUBj1
V6tqaYsx/GWOsKLu/UmGLLY3x90eCsfZV4VtYidp7GAOQYJaoG/X1kGoYW5nvWTR
TRZk+qlJYY46AYcLgNk0e79BOyY/Rf84hFhtSEIejIZh/KDLgyrYLt9WLG5pUPsW
+FxkonqRMG9qt+/Cxf+UW4qcDlXkOIjvnoPJ6GAfg+hgVTs0xDHssjCzuMKV7E7u
w6BR67dOd5+vG7fYmgEQR0MxyK7ltF2j1odByYSzKq0dNTo1NZA9lPC2IxeJHE0R
ep73GvtXoJ5lalHS2JYG8DqJc/A08Dl93EiB/61zYIpditA0GTEUJbUnaanogNFX
i0T1Us3czWbMC4rsmrDETVrkgaD01ZbgOQidnHIRXaR5LWIFXjI+VoTE3zGkfCsJ
ohVn6Sbesuo6ugQdvXmReRKd+LkHlkhwhiqEsqASe/Leusd7Xk4aUpk0M4hMLSxr
BS+hLli1ur5TSRN1zaracJGxwCA8Ng3jfUmE2lRVCoAYCvrLv6lNvDHYRxBGM2Ex
h5L2iE79Wk3zRbmtmC/M6AJUPIX1UndPptz/NBth5rpVqOfCbVR6MszMyXUTtNk3
MeotMqeEdhGJYI3KeD1EnytymABBzwGDooEdLFW3nHYtTFNWtHVZcW79PpC6lgnV
PigPV+mzioeqsBgWUIVvLKhHiiXyymvTZGUJMm4AUsaTOefAcHNBh66+OxCGOmzQ
959P38+fh8GZFT+LhUS01RDpWtqs6RGkpINeruAWlM14/IpgtPL0JDg/EMqo4hYY
mfQjKYfULCy/hoXpM8e5TQYS+An/LFXtiMB8YCZbxWVyD483mHNzSazcL19nBRXU
tsOBfsngXbFWuBYyATR7FoXBKYyttKyTbupReNRMgtCPKn/9ihWNbeVcPuVNGbLp
ULIBUz99XARi3gOcsQxVXCJltsC3j0YyVfph7UC9WOX2pTb777D3rxHYiSkttgqn
O23PpV8GgHRyvxF+7Og2qFx03T78Le5PbeCVktrEzDGaeK5NUTJLiMpMXHPhJYOQ
DIrIj9/hVbRCQfsSO7Ptu30NfflQJRIc4jDJTvsk/LmrC29UZ+oQhSikiZ9H40xv
pjevRC6i4mOo5yynNrU9rjeoNiSh00amU0CYvSOmGdpUaymriNhjPN/XJOvO1eI+
wCIz47ZtSI21iY4WLq6BMHLDK+G2/wOm8fnkWDm4SnJD+Wgpd9xZR96use0bybRc
AS+JzsQRaR8FWJ7lB1eBxrf78QAMhX48AVHON+606S20Ddj1QkMErpDoAWcXgOwr
DBIaB9+61hHBIeFlmL3NgUTJpkgteqODh2Dw8ESuZyWDnq2U5npTwoRHUILfwkIE
43qC7zBZtg7J6dmZwkf47YPc3yhHsonXmU2dpILWou4ssVSUj83vG8mqyBHQK9Mh
1ptjrSFAC7gFD8YcTTxeWDgKmz8utXEuNCljEks4ZQN2wmljf0MvyEKTIDMrEfhr
7tgVtopOILv+xeGCGDjs//Y6mOHbNa+Ey7RRxA0PKdkbDRzIvumT/vf6pil1Ugl/
GTydwbSXmdXnh+g9zjC3+Hsn0qum4C9ja6ZsJ9KFH5clxNOj7nHOMiznz1Bytiai
2oTk4xopZuKlxkOInkjGGQ==
`protect END_PROTECTED
