`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rzVgG91nfR7kRlYTOWPa+FCy/8YhXnbiN71n5Jx8H5RUqNFIJGhJYKxp4MwJr7eb
OCQKfnllZsqiBL8PUFJj+UcYTj8KTD9tDres7lf3M1DcX3yT97sxS412Vytk7FD4
sbXlr6JpE7GdYdekNIllwSL1RYSjoQeZO71sQpRHdqo/mVjhjkei0AZyRnx3eM2H
biitacBdHx74rhKIFOryuNl8B8PfUTzYH6oRtx+npYNWL3EuDMzrNMh63VYpPws8
c9lhQJY8btfkZqOc0jVD5ZeldQrAnmgNHazT1cNElZ4eec0mha6pcTf9mzU6i9fu
aK63+Wpo1tFmGn7N+mXxg7/ycl1BkerHvjbJaM/tXGEX4LzWBdidsCt6LOXSMtc8
VoMMWCpMSFUO2U2Ht75yjFQIo1Y60TM8rOwV4BDIxxQfooOijfaLDMXNCtULWSTg
PlEjzZQ7HcqqZVHogGgvD6kBZMtFOSByGxxgjdzIBQA735D8tunTqV4LxgpXqwS4
nj+WycVty4HPd1EZpvBcal/CDTMNZd9AArkbummmma+c47kMHiMuTBdT2aUHO6HV
S4pOGWgQjVRR+8QTeJAUwBI/6KMsWIIVRXzF7C+gbSQS8pW5lF3WQ8vzmLXmvpC4
TWqLf+8ZvxoDidd2zoqDDnt14Zzw+rEX/i1fG5gXHdoNlsVchZzciU5H0mqNVH0y
fEu0ozECLSgeqCeU+xxM9DIggUbjTfJur2mqGZ7znh/SALAvZ+zd9FnhWdm0+Axk
+POJMniyNYQU/ZqUwwMrmGOu62CsRXaz8jqop1AdjeOXti5y8nOwZsfwwlxC/tyC
JmHCLGxmN5BsiUFjDG/yq9RlyuUw4QgACkX6+5en5EI+WQ8f2BiqzJXgiUBI/IYj
S/DlN6/KU4a0fDk2WyWwuSvqYOwOqMU/pXsBZPC+nlVWpROaguC7JdmKnBIHlhy8
KzOtVZsfalkZOpjhL21P4yOvlA+XQf6LTe9Zqm4Hu6a2JI2vxJmhA8ZZPZwkNLZs
7/ZZr57Um3mSdCbCDEj2Bg==
`protect END_PROTECTED
