`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B87yJoE6ElZ3zymkbqsMENXmq2QW8ZkH+zUUfz6vmtGsSkYQwEFFqDX4xVFOhBrx
sgM+yNDRoAJD5HuER/6bL8ErNAdqw+LkhXEbm63ZLTaneD+vRXRw/PPipPQBPnSp
l7wCIIqyg+cwFUZ+bKNiqXIztOPRNo43Fxc6Fj8TBYaJWpoXCnhL64DMGjEQ9U7m
s0rVVNhISlR0RC6UF1AnNURDazz1TDySkUFTw0oTJ72/GGLg+/yEsgnA1zVy1yM/
YjD0dLLMmKSpDlXfj8VmKvXgEM8c83LszPwGucbLy1/sfaI5gMZmZ3qFmzw1b6nS
4UxcXoy3juErMdYtduzuqOOy5gi38dsWD4kOSWllRKaPGmWbUb/GPcJfz7L5E65J
lm/fWQHbu7bsTx6VASml5+Sw25il+7GyTLH3xbt9D7ULeqV0c37Av4eO4fFJfEeV
f4SwtrhWk6mYoEc9rlmUNQ==
`protect END_PROTECTED
