`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UZ2I3BEBFmOBWZoEKkBISB6fmZiDezZrJflEtw4AutaV0BoJ32/92o/6NpVWAcNR
JquBeuvO9jx/8A/LVm4RSqizU/g9J/bFcVNCWAQVeIhyVYxO6JDgeCjl5NPLnc3s
ebvILZzftOd64o4X+bPTPnUmCk2B8vnGCEHm6+8iCjSF0P2o/jIOUTsF2u23FlEa
dx8UBlxI6dxSSzI+syTSwu7MqrVwArmZqL7bhzEjRMqnjKpbKzuwJFUdqQAHyW1B
1afUw8EJHAAWQ6rGWvpovHtLfZb0Nw5x0uQYa9HVbUYnd6EJyZ88jAqKEwdI0nJ5
5d5VQt60CqU+DJN8hHlfcJ9NWIYAW08gUQpLYRS6VvwAPN6thCidxuG46RMXbudH
xSe3Vl9IjFloqnM5DaCh1lVj+fY4/+NyY1B28v/eA3+Xx4gvLCqSu4v5iptEKR9C
38RHT7HrXGxUtyrVK4xje8Aut3ZX+g4LW79vxgOuasGfF8JKfovyHbZVXhVC0aNY
ZQuMRuitT03sQho40dGo9rSDnnhL0Sj5i9xOLfGBEYU1jGVhA4khvatbpQdqo/6I
3dAU65Mrzc33p7Ipqxmb0ntVGq3rqkItmhHsLrtEWMx0GsbWZHPvdn8riPgQIm44
7WL+UZRckcZ9mH62nZrdcyLeWcLbpOojK9s+6bIn8GH/dFbA8W1iPuoCYsGFeYEJ
rQERALbPBKNjipurp9OpqWPA/a9o57dOyLgfT+jgLU8nnErZUZ7B+pt1pmswycSd
3hnf3xlEqkUhpJZNaAkJNRxAzXNQiGrEAaMf0EgXf0ab8yOk6a2xVA1ZbpKmpk9a
ZfrEMTfdksRiMvjpD4mFmBDDkKPd7FRMTm+8vqB3E8CKhfFO3TYnMHH9buehhAzB
NPFhLhPrpQdnTTf2iW9m0AX1rydIN1RF/e4UWXMPzrrG6U9JlCigSMx9JmVDdmRC
6pMTQ9y38zrHNcDXK6u9XkicZJqJWI+NV7YL5jFJKfeKD1b96FuXqKuPvLy812W4
a5ila19+8nhZQwjK65Uk9rAWCDDknx9guL/HTjRLc9H5vZV54fWlRy+uPRfq11xS
/yUVy4EXneSanBFsWGyGTwvjeEZ97iknE9kkTCPMddNA+tHptJL8uXpdUdwrJuUt
W2VEXUMqrKBnkNjlopF90FU48YjnLufA1pS1RT8QvfUJ4OFVApFAIiyohcukJlLR
JIvCChseY9g4U5TYPkms8FsMxbvEsxdLoIeQeo3XWmzfk+AtuY4BdYeIe/RVjKqM
KEmm3TZ9ReMPX5TYnzfAJ3EOkRviHGqE8QIAXighOIXY81prHUIh/+31hpOxMUFc
iD2+qmwnt3FLpqTIM0lUZ/xntdKYvay5SbPcIsac17JXICqIY6D9zZ00PCAMz2lH
ps7yR6uQtYoR4N/QLb7hU/8rrFNDtyR1/kkNzA8mjC0hsd8ryh7TdP/o52vsq7LR
0FQgSR4YG01tOrA/NypjhQYIBjFZlmoDb8TcgsiAQWMHS3Oh4zGNY8xkI9dmt/j3
17BfcN1ySGBGYJ5gJY9CUO82toJygYMTX/74epyIVeCiqjGCESgo2nWYsOHa5EiM
R2KWNAsHVKWyrZu6izuw+bI/qvj4vz0EJHSj+0FDgCFBJAceMI2d0M+f4HLkVw6B
bYoH8gm5G7N1+Td91SnKZ/Yn42vD1Qt06TP/CrSpEgYuI9tI0LfEe++lkw9xe2vY
LbMuX7bQ98krdCECH/em0tfPwb3LK3ZOOoIIb1kvEBXBC/uICGQ2K99JPHWo5CWi
dSranIIPtc/90lt/wesB40mRgAMFsLyOgbGH7AqS7DHDIBy1/XM6hc5nuyaNvN+Y
1MTQkegd3r6vj7CZyvKS9dWCnjSOEhKGCoTgcXl9NFBQmMQ71DtLlhEGuHCyWHAt
GitTsHCpPQb+Vl8MxuRg6LioRW8fZRT5n1GDEm3RjCoxQ4icifjsMa4FCFF3Bx9L
u+i6QBePzlr/SnWSiYEHE+XLQD5zBcqiJc9S3igPg7Y2x6LkxLTWuQ86kS6vQ8CD
NUjmKcgI01hlAghH/TIpbFKYnENz/wako8OS3Rm2AUh3FLjye9GQdOuqjoo+O5BV
SRgeRx8AYrEQ9Hhfsj4DZTP6Xmm06cNeSfuMGBLnLE12pjWniWon8yTbjlLkTvfV
KpTdVA3jQcoYa1fWm0I8wergXKJo9ODuLEpRyHJJVM1FbxEdEwETGtRhzj6pGJ8m
tPaCdsak4fXaCyScOyWqTGvWq01240/rdh4l+lVwLGLKmFHtqty5Ow1u33S6rD+t
1vKrzcCTC71e9SMFfoHzoewkFV5wmEofjse/nwCBK5KEKQK1feDoKXQCunz2prtD
xZpTUYqbSmluCAfcyNUSQp1d7VDKy+PYv+rkPiWNz3NWFTOOyCC5x/RHAEMJXXO1
jLyLEYgFhN2Q8StOnaYEG7Hkv3MJ4r0578JH2JJruSmW6jjbzMSOu5tK7j1ddLT/
+ecaaNuvIIDy6W0MrlX+ZSgbUFtPR0Vc8WhxEka2SJPn8is49Jg20lHTYBqtBUI6
GD8+cI9odRFgagNNR8qaow57iW4ZmbeNa+dz1N3pVDlNiYOz/TGBqtfTZrZNfM9n
DOUVtTP4CSxAsYsNIRPf4cLteOEpaiY5urEgjH0VWu/cCnMBLuFzQnIuyzW9bgiG
kJRrterA/TDhY9vFgZYxGfHMZ9nOi8L/vdwWSu/LFTiLG9j7nuOvhT7QWtfK4SUJ
K/W2ZeWUnhUAI0ql8Gs/bx7wrdV9642vUmzeKaSsvY4q4jySQl6Z1f94Y54Glpa3
WwWjREbOolmdhAI+/GqvgSqMyp0f9TS6JzUXEy4HdYRsmY1ArRtgrx0dZF1tIF6q
hQ8OkMQphKuDAo/EbgLzziMEIQixqjf+ZAR2U4xg6RB2/HJ8Qztoxeu3GwXHqzSR
z7/h3CJsWapMLmf7nkpuUAAYb8jWroi9hz+lJ+3SLUhPl21ExPU5fsrXh3Apdg36
vPxmWz4JC6Wq+sHLbNKj1HYPwvb0IiS0AX/kDevAx7cqJVOLr20VQ7Vj/34tUkeo
MEra5X1rsZt/6d6/BLp/QOzETRpceFbXdtla77L5EgFAMwo2pnSxh0CLZIlUS4vN
N/0eJYC+4elv7ILu1BpaQI4O/PTTZ3iDuGNk2v9moFJlUksvIlz/BeVBZki++oj9
l9yXJrqVTXl1vU1vD1Uw80ZgEGRzPnx5IGJbh/x/BKExvadLz2mceyL7EMUoK86p
Gt/3gAoGnGTaKaOkykiuejz8rmzE/zCP77wJIi/R0Fj8iBQHTQsHHgYzzhyl5Bbm
Ry/NJTSlD7bHmq+MKsYOLVz0gFTvxo8pYAl1mFM9RE6YEo52NK8HuTz9zdWy8fMi
waB7sKCuH3rjhGSpUe9kzUyiMi7goBcanhAcRzFRsIhtiey5oKQzuMU5b2+ETAX3
ZN46Pszs6l+xpdQYW3yq9k2L0Czp8glmoINN5T1fxMLqBJs18P9+RkhHQbqu/yba
pKOyDTK/nz7j+u2dUr4B8aMmsUFT9B2wB0I6kbPTc9tcfGl2M/pm+3pQ0L9CcM0p
sykKScKw1sIUn5FmkqdRQCFughd79V/hpmns58FdR3QN9DwPASBBxweSN8eQA11B
k55dyzWRg3NK4L7NhqMKV14CMtnuyKp757lQm3AuUu8axHULPcpUpz97ux/Bc2tn
9K9LSkUDqCcbyZRpVY21HaY56hd3qUENxrSMSSWfGCDokaxRvigvtn6XDmzyt7uh
/Om9E0dVLf6s43cqZdtrbgRAkp5PKc7TQLs+n0OJ9UN42DGRwE9e9n4qyR0E/DH2
AC48+e52IEBwVBu8irQjyxC4R2BjIK6n8vwRBmObNIA8ZAV+Sv0OxXCDmJbZeoqU
zMRIVF8i0E9TorqS8VITrHup+iWOY/gBhnS1WJhp/7lnJitMOrHxbJZwJpNvJh4Y
l++rO2ZB8jMzMnA0b/MUZtgPK4N8Ox/CsIvlGHT0y1VZlwi78bww5qs7AAFqzxRa
JtGLrx3zEhWvSiWBa80vswZkvrCBGxhsZSTleY4I7KzjkgQH2vojO7Ua7MzWmX4J
NBE2PfuJFLRYGVEmXI0SkIyOLqgRmLE6ZM2lakEH1XvinVjmS5aHX13MDzZrT7Fo
//aHOGnw6slh0fo0xL1aKW3n4rNHw6inWafksrvqAMDBtWeqO6jr6cDUNAv7YxBU
fWRX9/DT24RDhSkS4aS8jNACc3YUjemDdqQ/4bfcJdxN8l5Ab+B0Hiqpj9ngA0G9
IQTrf4kJ6qN069YlwMq/3LTEkIqda6P8Mqn0Am3zP6cIUfdqx3tFfeCvZWKOGUBy
e6A6oF3PKmZg/4zD4ghusagFlmOGJ3/ihe0u6f7Xyj/zE2gdS5tdW4ClbT/Zg+bY
XNvsch+dgWSpIQZwwWtVq0I4v4byezOBza66gfr0qMK0q4+ADQDW4IRXTIFDOEXQ
j/LcwBydtr8KM6xEHbq0/JfYFzfk44dIKxJTHFV3bBzwf/uBDpS2o4+79+OOqv9u
zU5U7PirFu7wBD49MQCsQWrDQta7hSe3bOxEJHV06FRrpCtjQbdQ7NGyqdtp4S9K
cCh3uT2mLvCHZoufpLlVxRgkt/dgvkZ61KrBD2FN/jM=
`protect END_PROTECTED
