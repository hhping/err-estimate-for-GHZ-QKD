`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JBJA3zN0olKPlH3eCffcJVsweBhWDOnqoDJtQjHJUVxLs0JxqejraIVY0UHqlCHs
6w5bENAiEj7PrCxt3tT0+s1g94AaPwI8AYPdmSXULqVKunPV3JKgMtC9BL3C8UYC
bq60wI3pfqxQcv7vk66vpapzXqHQswSULVYWOK9crXrWoWSXeEFGscg5426ad6au
6VAIKUpQlKzkE14Pehr4ZE5E/TN0wOAYcn9jO246yN6O4A/9ZIes0V/fQFPAShFg
BEtoBseeZ/pQ6bDuHUDqp3ZJ+R2C24ySLeffE8X/dNaE+jfLTisSPUc8mPYwJUmF
9M+Cfnhfl+CAHvc6cM7bx8X9roNl9OZDISLz77+jrhXyIhScz8dw7sU6MwHdUu5a
HzCC5rhCQ846Mqr/toCgJnZ53pdqJn4aiozHXsfsvzH+pv6fFENdx/sWAugxvndN
sxPKMKVDfWMCO+TCsIb1gvU3BGaeXUxlugRuRlgMX9u+BW43DCiphHvIEy69dRo7
1clgXsx3LD0/shCyFjrzHcmB2a+tASL1SBogBdbqK5by3Tdovt/pQgtyCRHOLd70
SxLu95q3KKJ+QmxdwfhP4yQ7rm4+3JTUvvADgwfM/iKZHCqpljjpjFT5FDjDt8zX
2JvPxp9j60KtPAjUkwuewlW8zZFqxt/TXIZBbmF4s+9OJ2hjKWuZdm2gB0e4JXGY
v/EpyEI3TzGv75xJ/CcsCA==
`protect END_PROTECTED
