`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QWmrPTs2Qc6YnCd9mXYnks7WuIyzr4uSPHvFbtLEjRCzPul6QfTc6/WDSHl4Hf+S
8PEcuZCaauWFW2OsMfx7mho4LVyB05lr94sA5FzRwQr1kUIIIMvB16C5VFTkawXo
7ED62BWQf0728yZkUt3Vj4Uqzez3Bap3HiCHr415tGFW4v9zwmli3sNo1miwDVGW
y+Nco2dd2wzJOTG7ZlANL7Q9US6ON1qwBHS80Qled89lhwIzIw+SJAKKi7T3m+ae
3pgMjMF6v97ZwCEVVwTIqkezIlEE64cSXpPNayUfSrfc2bCYPjO3s3K4JY1ajAKr
pM4xDePJbb6Vh3TXlbT/i4bqAUA4+BfyTXn36DWcEGB4qKt5+ebcpbtIoBRziBT3
Sz7c7MMmNPzDXH8YZOb6Z2iTWebFjk/Z9Njrm2W50VpTLIe7iDC0ZswZpR/+TX6X
uaCbRqTBbcPYAoAmYUh4W2EdAceoOleLLNr+d1m7WJov3kqVvia35CZELf5w91Iv
4ma9cD3jqUWf1hBUj1K3JTNLvRk4BK1ouyML+Aa3uNvRQwbscvaSc1wm2uc1sBw2
igEOGR/jWGi7fQ0FhrFFXjjdpg+3AEnNGSOVBvz5rAQeiSlZNHF5OYc8/iwMeNAV
W8TyaPRgj+oeN4Et1eKHGjFn1mLS22Sm+TzIbWW43FTA9VaKhC4nSarWeaWopTn6
KTxGFNDUFCFVMJwEEUhECdGjE0ffp/FC+hxP+FLaQUP2gkka51H35Nr8/1d/Id9B
BPuKqKmwmKKqkikjAOhD23Sq9K5uwVMk63Qjg1QfZM6eFdMuBF594z5hxV+qwrME
VGqCjbQJtY6FzkOT+OlddED7FWFwWnqGk6+fZhQEpmHlZwVU9Ektqt8ML0lzJf7C
tFE3knk192jP2zfewHmLBySjgRDL9kmDCa2PgATdWnEoDc4MFyfnAF4UrhybxRXi
AACJr8vIhXj6owicfqXKBxbZ+goU96VCdI7/pqk2sKNg1WDPqZYpDJBCfw7gJVsu
9pC80zpRIanszpRL6+MK7AXqildFBGb2NLjvai/O2hyokM/G35k9oGkOVCSN6fxC
3NSzUEGt/CNqolVr+umOidfMu7X/+gQalQ6l8pCQ2Bpfz1sm0eN6IJWmXi1HEpEP
7oYwZYzEYY7SdOXAR/TkAnHlzrjsJGLNU3ml8rgboX9P0kqw4onfnB01gIk+KVHh
l79V3TUrwdeGGcWOCk1lN53JoAWRMZK06id7xZK9WRE=
`protect END_PROTECTED
