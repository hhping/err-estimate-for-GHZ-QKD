`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gjtIk9GYwxYpIsZ4vI0/nYXAiJ4UlN97hX1Ba8KMtnOghNcMCC7f3sqjHek/Ldrt
RD5e4upR5gaaJaWR98uCjwvXLpMs72Ni7N5OljTu34ZNPuQYOaXZLwETncmTfSzc
SCBSAmaz14H/fvjoapGvu2NI8KeTmUNw5vlJigH3VFEFB1PEG2ADD8UhufLy84T8
KX/Sry8/FHPuZ3dDV74VCcJSShw90y5X/TXtNqK9fXHG3tj4i5fw8+dCTHvnH6P5
zU2TgRWB4vxr3XhjW6IPlgHcTf6IV7xZgxOJ+WQZyu3dFxNASOvxiLHgGnj0sM92
iMFQzA4w52lYApvwTPhc3yzuPsZVnTGgifL/VAgaEvwPES6jROxtw3ANd5hNmOwO
NHly/OYKgPzfDXnR901Vux2+xqS0OWJJ2t9+Xh3oxBPFbyAU11C2UgUOnhymiG+7
8V0YylwKLSjkulmRtPexlZuuSiDTkiSfBjqNPJlBZAWAJoMUlOpmsHU6EM9Bt6a2
n5xN07pZuarIs0D4oUp7KWEUo6KFXqparTwaYewGeYNVxtR+PLZt2PcpIHB7JLiS
Uyy6WCTxwadBw8FBp8uviXZ0nJCOOkA56/i1A40VE2x5tTtMxCsDz71MKpUBI3LZ
fT62CvkgDShcTyShYRT0kQDitaZOZiJNpnDLSxje+XFOiUVgLoAw8uBh5SxgUJdZ
Ye1Lx02FbNaa9S//c26HNqvHL2dYxORhIxYCjLtUfUDeUa/ZL9FeTrynfs5doQjA
L8cUPeq0jE92xwsbrvrbLx0nongUkoDvTuGGV8BpA5oVP2ar8exnajwjOckg4Bwz
4/IBoEOkq1urSfurI2FJo2TO00YrHL1cAeXdkM0lmAFggPL3RuuCZwZUPjHdDbuD
1kXjwSTx3XfnJkISRZVJ6WxA6pT90GRI/hiaePfqItJPIoStIaYsDa0ZVPlGC1r0
3H6dpNHL8toVhC60dTGeQElkLtKYQBOVRIAlzDpHDfHBDrfSFDMTbV7++pT3KxGt
SlSUXv22kGvoFDIRLGO+uSzt7Q63iWUJYZUbHIXbRRZ6YZt14gjf/YIoSxdi09z8
mIU8m/oWCSGyN1riliabV8832Ad3QtUASc6our5ZTs3r9FEo+vicqs9c5jijbXur
pHYeKm2zq6Tu3C7xR2lQJiIMVkxfKVrkUt+0XPSde7k8ubUVC56pngGp/7b8/AUu
+rdNvUgjK1BO8OlwQ8VmIZzfv4Zm+6rtvXxfV1InbiTTwTcGaN4FbEvRVPcleir2
9cNuKMR7fsW8Xb81KhG3VPIrzlTdva/VkV+oxAvIjYu80cy0vLrmuszJDAksjDmk
ByCgEegDNLgOsyDdkb6cqOj6TiVizmr+kRe4XXS0I+c356X/GOyCbZ/CTff0ftnQ
Qda+e1efdI5cjpQp4zdn0SttbCH3SMm6dVusdaHMWtK4Iunx8p0rc5SRhuktyR9J
sofl15cY/clcKZFwI8HglVvu2C4V96kwPX21iyOkhl5cxfcHzj7QgkSV9XDkmhZi
H27LaEYSFuQ9BFdaOsBKkmiYgM8hE7apdxwLf+iSbCPF1mry38CJ869WHap6yyV3
BvC8P2+XStJUef25TSz7OhnDdOWnn7XN3knOidMx09BhRdM48SmPwQ+N+jFWUnHx
63Q37+cIfIP7L8Oo2zUHKxj6SGZC/PHpnDxcq2mZnJwAdDsR592ZBm6Xf3jVbarq
r1yIjll510Bm6O5iHYWwCCNRKFESX6l88Yb0ixuE9SVojzt+z9WK6zk6ET9Un+lt
mr4hAjY+Ix18NrcIXoqbA5SzvU2OgBr8nUGEkgpX7RLPIkNDZNYGmPDBVS+XP8sJ
uR3AxTz2ALFdEn+omy4m+/ANFQRDRB6JvCrmGubagkZn98uUgMktcKQXkF0MHKuk
5OPJx7MkvC7ZlrbFJHZH+nMVXPAfBf2tQoUzJNMEMvTuy6gPjtMrsRNBRJgHWOhw
n8DbJMBAx5QQRSwc7RgdgFoY9rnfSA+EEUQqgdWSoQpJ3wLMch/gm7YpiXaBDnz9
BVxFpg88qbDuF7j1WHq9xlSHBPyzlpvG+hB19NI2rb5lJKigXKIFwG7IyQ0snphn
NltJ+T/EFgigUo0yuN23fktnGfd2lKZXxWednmIS+Pa+YXxhSe/I3QVg728S5syb
aZCiHX82pXuyiH+QzyoIWnLZqyotUVhK0143Jjc6Ukz8kJqilJokp6hyICWRm9tv
CdOoWCv3Mg4mZ4JAy0fwHsRvViyDh6oIvo9yoQVF1B/BN650x93bWEW7LQ50Hsa3
bn5Q+aSwOvwLctG2SdJ9HzAFrVxjpKdK4/hlVXYpQHgX7u6E+3YX25IN0fbATTKr
K1EyPO+s2g5gcTn75LHxv5tla2iqL28dl3eZEBsarKlSzbzhEtKTx3lJIu7Bu9Uy
KGCFzDhot3hEraBfESnV7FOQxfsCn0ko6r19rvjVES6203YlhkJq47urjgB1vL0Y
F7bx8W2fvPxEamllmDT9fznzgP6XqAYtZPNwLz90qWn37HxRxnyhF4WmFzK/aLye
teBge6CIRCWJTnKq+LGD8MVcjE//0Qy5FfQUPmjbvh6mIz6t4wYPoIMrg3tTOmy0
Umn7E34TtlL0PmmYGE13UoKykvi7uoH9FHfRfuN/ezLN5v1DJ70XvctLCEB3GBVl
xy3S8iTCR5q8bNJzOFtg8UHKumlhS+BNJCWm8Qgko4o8w1HPohzbo4PpZwyKFQXp
T2pO6Kez3GHHfhI+f95GM0jNH2crpdUH0I5nFOxWNRZ3h2knsRi/Ck8etF1YN/S6
E6qa5ReNVDrk1DgpwkDYpJVgJ1GLEwS2nlpQ8hg0JWzGpHxCZWbmx2Jb1caQ5a1b
sPZgJrJlrlwU2BL57gDxoAXeeuH1nyL+fx9fSk/6AoVosIX+TtM1vDZU6eZ1/Uny
VM1d/CCqoVgZ/GVxy9FvLkJv6rPqW5DHGJ0fgbcL9ZN8JD0mmqZS4jnUzXSpZtmf
TyvdQUxdn1z7W6WUouGYQu2azfZF6H6ftiF6NsHKU8s=
`protect END_PROTECTED
