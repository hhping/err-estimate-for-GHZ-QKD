`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FDpcHVjiSy0DSvKbV4TRsgfn5CzKSiuJtSEF5ZulHCrBeeIVtoTI7INfUDfr3P2z
eR5Y0ZiaPzOHG5g/19F7TJGPPw4KaWnbAa7L5j29g/4Kylli37TlASURjf/7LZ/L
RgSb0qFimcIq8LptOA9mxyTmaGCMtGf9ozF0zZyp7AB1oz0aHnoPq6GgJ0jOpz1b
L3cmBns58VRxhH3yG3+BHciO8Tp2gnFbNwEax+9A0YFO0H8ftXMSy0H5J2/GncYh
vEtH02go3J2AZG/l2AtH4Rj2MQbpaP1s34OVb8RbXTA3sFyVLTZYAhsV1E8cyhw3
Z+HLawVv7iN8QNRD6gE6nu0EWPobkbwiunmn5WRwlZgaRwvgjTQTQH7ORgspnV4v
`protect END_PROTECTED
