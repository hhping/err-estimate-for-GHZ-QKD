`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OdQ1t/cDZG1shH3PWCHer2ROMQ03TbhXI8TijGxxIFg84HIn0aVNh/MABrLtN3Zz
X1K4RwluwuZX6kC5O30/8GNDQxTTkIAlwgkRIEKNnF/3fAgqzu4DYyGvxBcbeB0Y
nZjy+tPVZ4UwKAK//wRYv697ACRu87Dj4GX15POts0T8I2JwBlf/X2fba66KD4xO
N1y+Vse/IbUO5CAycEmcQlwo/zrcN7T3uFGLlArSmLpsfHgt9joCeE+NwSKqeNeK
nLdAafroTqBhNJrYxyEt7CTHfHldgUz6g3Im9thtep3x1xjtMErZwD1GdvLBnKnL
50AbfU6JzZ9lnGD60sAfNT8oxpyvCyqCFiYdaO9+jNnh+MSggyOoAwM+pJpecilp
AXt9tQduanrwOlvWVasd1kC7TYXbHu8q32w5E06JIG3N/3Dpx/jfpbuxfRTkG1OF
kr0IqnG/X5kEsqfXqkRbAIT3qF7vcDYHJtwJmgY//5ZeJ0KsW1IaAmZmzc+RX7IY
pXhJZU55lM6rd2hUvCd+mZt3Kq6Nz1BV7ABetyAGN5c+QmePmGDSovtg5MBG89KA
eG4sX2NcJuZ6ZPSClx8JwHD4B0II61cJLWhx6u4zu23gy8FLkS4sVqDGshce23lo
PyBqKN//wtpb8UBbwkM0Gwg7jhzMBRJ28Tn95E4xRY8pvRJxZ3qXfFUWR8Isl27Z
hCaNEcvAXp7SWMLgGHQeL9eJExXCqqqJc4A+ZQ/3K5l/4ND3iDHOYRMc4fj1p85r
B+rdwkT9QSLs9l2rSjqS41ozQJqcYqzZ09CnFRUVHX3zbOvNY/VpO6wp78AEMi2I
wvrxhDUf4iJW3uRnZEa7e6yZeHol0tF+cOJ+pPYuG3zFkxdDMhVOckWXfAyfDISf
gpxmBaQMD8tU1QoBTNtm822k4GEwGTAiz6bCUrfIOCg7GYD2XqKEZMol+HNT5P/t
Zz/CF5i+d7KYYpRbY3wNZbZSTUOzX/irfza3b847Vy40qiybEZN5cbBZv0Vu7MNX
GBCr42Ajb/gvbzudX6E4DPpwVUWZ+ZcyJZqsu1M/8yqIuMn1zfsxhcAmdrTHlVb0
77wMP2q/98S3hUFWlP9gGStzkXohSnN47zPp1Ds9BjA=
`protect END_PROTECTED
