`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pQAhSUHXrq5FNPGmkACqNFwZ3vlPIG18xvQLI8y0Y89UM7WkLrEi43cPjK7MlXhi
yl2YmyGF/rImucNi+mIPaoJKkghGdN4BJou7zem8Vkk2HWScPpkkKwVmrlQ5Ejv/
kK2qQSzfAk9MC1odEzONZj90Mu6evHK2PSRl30Nfvx3KRtJaT1FayoqjkGlPbwXd
V9IgeGm3TgLCgvbNmrnXbGbhkA6H/mI397BDa6TJ6gXYEVXD2YC1TpblSTULnWut
n+vUAtHBh5qMFRrspsxM0PV/TPVPLug0o9SI6SGM4KhaPuEu0KeUHmm2/rICR/CT
A6b0IHpMp5yohpfX7gJIzMnBz2hlxORqEKG1nGyO82AITSTdqsNIEdw17F4TuTSH
3pguwblHtk/vek9YHlDJ9UHnOCp/srP2CDWbXjod+ZYli8VMYDP+tiFOQ79BUf+S
ELSZ6joKjiS/J1qii41v6Va13cGbZwFOTXfnnPxyjTcoZbs1zJ8mrSaOPTdNdlk7
5pE8u80PhJTY7E/tB60fQWkUeP4sf478D7Cr735Sb+Tt8jYCP5ujk9l43m5tcNQM
tOhnDvpUFDKqL0e4YyeSxcXkA6lmurdrq4/RQPPoEUjMvElTiKnZYEkObdOdRPXO
KZFjIM+2RDUMzGGB+ZBTQOwcPBajav7VzzCVGy6mxOPRXbMhtoyk2/PZViGOd/iL
NrIZN9tuUU9HV/cdgD0q7TqnQeFj4qEFc5kUJdyC9Or5v0TdLSRP/xHbwzMbV/uc
eCGkhqJQy1borchT4tphepPPEPq6DFFV22zgHQNbLAZz1sxdlPgG/ShcAUMmC8Kq
rdFxvTVNSM4J2HyedA0NqtIJFdx4+85qcIsqUK6qylj9bRJ1tPwN9/04FJISC7m4
hkSNo0X8amf10zoWNUJa2PSYw/1A8UPG9xBvyR87w83AVuPk5jlM739rGjLAK533
/ZR+O2tE0PAm7SaCV9bgxwAqjVT86+xSdg4viVqxd/Fl8Ca3o2bOeG7iiO2gyR5Q
KsE3ntYQhHkcMSlIUfTJEg9qkr5UoQgtzayrDBanc03b7goIBgRqtXO5qWlC3EEK
zlDKSCY5D7PhjeTAC15GUOV/erKxbL27652mAPR1O5gXq2pZbvlSMOs4aWZc74Kx
rwElUJEnfbo29awqzo6kmSsE+lNTPtRPLDhZVctIDvj6iqaP4i6yR5YK5bAXNf4L
YmGzMZEJJXDjTIfIITd1akQ1nv5pe7j4vRtZQ9+bLYl+JBWIi6QQd2xm7cz3Ea8v
9QW55TMFpq5uvV89W6EE/WMSc7TNFvo3W/9Hu/atHnM6JuAuE59H6rxjOXQr7Yf6
yjyAs3EitYll5Nn484tXUAvwxqjGf2IUgtOTZiNxkTuroG+7qSJrzIPvjmET8Z2G
mtUP/ywH/Y8YU6t7TP7AZNyZybPjeXcHLM4WPXHp088LHph01UPht7xwSkhtppE8
ln1e8ih0PdAqETCUOxD1/Td3ju06CKI+RC240TfNph+HkEFgg/5iSczTcAe9Pmb6
aa+M/vn7tity4snnJhTBp0YJML0YVYWc1WUSdAORy5mBk+5yW3okKkSAlLYbzV/m
Fz7KxW3JvdrfwrdRO4CLOav3XEhITjHOoOXya3Npi3wAO5IIB+l0NKPvROJmFGpx
PFeePMAEf3x0u+ZQyddF1XFcxQaXHXFvV0BvZD0AD3y/dLEeHDvnU5LLN+fJbocI
xp9SohjUzvkFsCZhCkV3v/0UK8Bo7aeER1/n2uUU1gup5h4rsQSYdNV7uARQKBy2
kCMtFkDOC8HaJudFlTJFsUEXFmyVQ4DVsp5vY+W2lVGPg+csKmpB/Eq/Cb9HggX9
quDDcw/NFz2vFzJxVPQrpiWcOF31ysc3veZl3EfYv1uKOERDIe9LOAtO1sikaDPO
UuWu4+nAbAVfPchp+itubfjiJ0tkVZnsqLZ+1o+rc4F1u2cTKZI5SW9kKtlcefPL
vl2yzgSCklMQUDa8HmpvPe4uYuF15eTHWJ0+5y6m8Ar3VvGRmxqbHmg6rM2PENqO
6tenJrBI2Ir9Wr4QFSj0TuJNo3nvxbj5rtZZa3020Z9W/2O1F7jXtfnuhKAbqChI
HcegBLwMsWUQL8KThyzoUlI1WMv9vtKzG7vaCPiizyrw5fsj9mSbHkmIP8gkTpsV
IHElHdhDL32k+Ywd/7n+dQOX6ROtrU62VMtJIMvzxYXU6vrMeNsSxE63+h1c1Kt4
0rK/9ByR9nI6BxEhXP4LNNFml4TZMR22UJd3QgPc5alAUw41PJm+Q0FsKVdQwB3B
ZG63UhaUVPANKY7LZLa8R/I8eQelZSkR1y5Cj/MBhczmowygmUsrT78km7DIIn6t
UT0F9uXSxnJidhrLMU2Ler0+zf3/NOPhCcmpajE8s1KnF9j7mHxTpNrsM4LAbmW/
PB5ewvBPZJpwW9IkdTYzSn1qJr6ZYBliOWyHTrKUwwB2KLXTqMOuzwfCZsA0zDHo
ipiw++zZjWc+xqo+G22YavT4JxmXYgA813sxjfsGUGQbzUZ/bUTuMdv9hiO1uPTV
rt0R4aCiGId2QicodE88A73QTmu7+Jv/OvsqfgzEhucwC42OSjJkFNOZlnglSDkH
Da9XeQg90ksgEkh7fZNMJl5xABvccf2yPkwi8ylPGGon/HCp09ZJHHloRCrd2W4d
+1g7/LoT94SXNVhZFznPLkMFNyq631LlWTVYXlTMwkVMX48a3fYayGlILEkGKjlO
5/kw3O++K9DU80LHB+lx44gsqGEa6wmZ0kQYH3gTiEyvzuqj8l8N9U0GEe+kQuzT
u/muU51lY7CCuBR5m6GpuRTkWNBIJkLr07yIOgo41pR0WwSoqcpbgHLjktK6IAa+
yQepVWCOU6OD/BUv2tYhJfcidWIksQXIfZeJDE0Ubr3XBNeJ14Qr0HPZkv7wlS6D
EXFGIj9mHXAe4G3RypRhQ9eMfzYx3p/Fak4lNwp7onRddRjkOcd/Crw1KaelLVxH
0wO/cbxc1EEmlHgwDZ/gm5eqFIRkeVnLB5crITimEEaUC4TVNwKEtRlDTO48rYa7
Z9pL/RliQW5T9lD2Y5MftnrBTnm1MZiyNTzVVgLA/gSZPfHEfkzeqwEbl5p3iKuU
2Ca3Zj7KlkXKTW0FoYIDrVye+0KE7uFjh/axeVqsR19d9Z4a+WlaCI5J+E5huMY6
GDVs8CMUFTIQbuefDRs3XDC4iqkBE1tKfLkZ6THaGsXmlkSSaJwR//7tkU4AAmB2
+1tGY/9roufG8lXv2KX0F7EvG/3BRqokMU0OVQtOl4Tz+QiAvxNvx5XSdoYnx2JK
kgXwpnsm6EI5EAcDMzNCqj9xdPbFog8QOWnhEQeoGJ+02TQRPKlneIEa1cXTyMKB
M/GyDbhDixamYGxgYKeRDhmsEna/fKKq1V23uLNrWzPvFeQGwy3SwNF8I+WcLTB+
orf0MyERiQ/ZvZvRzlXt6RtY+TK2l7FRleuUM8K8XUcgVWZVPRZNxuFdFYMgGCcM
bbrmnPzwPW5NQFXACytjtPXX5gMZmApEBZ2a4N+eAiT7MBo6V6+q1waxgKQ5qKK8
s6yQqq88P3ToVMSWFnXmFILm7urOFypTtQyqbUoPOTH0MNi6HJAiuezFF+JfuvbN
u6eU/DkSfTbeLOB6UXqOOjETETFPvn95Qho2aJT/2Yw=
`protect END_PROTECTED
