`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
klSBXSDZZ5dCwXsT8folnJTCy0yF7zAUdmi0m6NyHA1JqoOUZHiUO4rPp8UYPGdG
oJkzkzlH0CHT0Pr9hZDLmb33wWklqZsY1v5r3DJdfl/3zBDeNVsKy6IdwNirdL6U
UyNZ3+of5fB+KG+hVolAmsy10jWHyPzivfCAmVhbOvHG+EBVtWQ5248YtZqZztmb
fXkXFkD7JntIDoI3gyNZuTDu/CIa44/E+YEkut02vKp3OfoUGozFTUVag8wJguKj
aS5LVFbGtrCWeAF5KPZ4orZGPGFgqKMOdkAJPoZ+ni170AVDWfWK6n9yJT97wUmk
RJxs9VKGz9iTRmWeVyUdvOc8c6SzEczj3IAUIrzCQarYAIEJQMIIxer1p8MzbQVb
du5AzGMPZazuev1g6vU4KLyGRrb5E5BgqZtxovhMtqFPAvp952VcD5uCvfOwdspS
segqnwjpXb2XIE6sDozmRWjrSGbkHLuueM7GbxjFpqxXnPiA6avuzQ2XgsDCt2Wt
Bp9knA28yW7zzjwWxBoSV8x0eUfwsf1qKaDa4N7wUEDDGhsTVzg2GcosViG2tR/V
vjDL8cnikEaPmrD5ZRYRy34OZPxeSVlOysQfQ174g2PAipYUybikP/7g8DoNPYD9
HUPIbgU6EXrCdk9LXdfN7YwHSzzLlooZAc4zBKcw3+Qprgyap3wieWRkeW2Y+9KT
JngsZPJ2+Mr8h50ORlDKshafEJ7bvvFT/HXYVGjUd5XXEUWv85mtMPP0sybrlNfK
gyb1CgJ8WF4s+I0/El5r4MFFz7UlVVvqYPvX9vW0FJlRTsaxj4DXPDL8x1lpT6Hv
6he++0nIr96+TrwD7ZygAI2MYNbGkVC25EJQPpMPKwoBvR5MzoKeD3+4GKQDLRjP
CBn79H/KCiU6b6MnvUpTjQQSwYk8RseS8A6f5YL8/MZoa/kY6V0VRry+58tnTp7d
i2hvAS5bBneeULlD1EPxwq8z7FI30HFjo9/LFIflSobNQXWu3ZIHrRfb7w6zgjpK
QCQ3YcogdsDXtUaHLvhkGjV5igbYzOvwV+9Q/t0IIF05YjlNMvvxrsCwi9te+FUG
hLIc8lutCGMUBSecYWppO/FkHhafKbeMsYq0Q4TISGkrWV1vLKGE3aW5m5N9tHxR
6GnXgli64kBYzIHgPeKe2+fUN9hGUkI22HIigyF3GH7BlBRqweOqHFtszm8sleHD
jhpe7hraDos5dySjsCVJ4BBP0ctyWaVEMccq+iDw3b1bKl3gZbxqRn6mdjJwkAVo
VYPNynNKo1MVjnW1DHjIo1H7vM+u/ly0NcMEnkWkEPC+5yCzCGmMJ4xlBtai1e8L
SYoxfrQHkc5+y02xjixyATu910/Ve8u/+1/VixR+oMtm6AlXgXIFsf9xCu7f8kwB
ZTGgnNbq2VtkvffJtrw4ZyHUH2dv7U9EBzqIHDZaOLNAZLl99TBru0Kn5GM9oN4S
bACKlXymxFLPIgr4ORLV9LoXGO5P81LSHFZAAvrOHm3po+vrN+JjNvUryV9LM4P9
F3CJZf5LNGSRrXmbJgGpoRWpuxTaRM0S8XMJvsDPrfUeOpKSJ/luQmR3nKkZ/KXK
lBvolpzwkB3mP0PaxsIT6BwCZULzQs1DpKVE9clg99T4mi94qZkoYJl9qmC8Uqi1
PsxfOX5P52fp/HcrrYTz/oU62zyzll2urKFv0BrEize7x2da9GWdLpWq3g8IBFSm
uApHcU/0Ua9pqCDAkwJSzRcwmDdrih5QRdI5MtYpvpjoxas5/VbCIIqjLrLqp10K
g/ZbP3ee4Pupp5INKbQOUFLcqO1Iwre0tQ7n3rlLzOCr/aunRoh23j29ABgD/PAz
wbbESTATN+FXhYNp6LyxngI+7Mzz5vc5MHi3UJeekITgQL41B6ZA/DHfDN1kWQAY
rg4d00np/dI6/taFDUBT6uxL6HZ7ICj/evwesABC4kv6OgVuo91M/TAdiME1yEDx
Q6VgxtGF+F65M57WUkYTuZvAID68amE7VkfpKp+3xktCsUL50WYikZtW14aI5nSS
Qu7ADf1jJ7/tQRJWFImhW4epTszlbwVl7pp/xlfehwh+ZHcO7BPScG0dbGZpn2i+
eu5VpIamjpj0b4vYanpxG159ygySZca+AkJO75IFaAjADmU4yk5wg0EN3+yykaxU
GEjB1MujN/K6uI5Jui8cXyXyHwLuiCwm2NAks34yzzBtxdnJ1q0pcHpr8wDsXfgn
owqHKWCiQgUQpWIi7ELtM3xC+vi6uIKR64InymcF0NbfoyzzNmkV1+6MCtqP2YlK
2fpX/dVMzNIuQywF/JL28zgcmJsoKEEAYNyV/U6PgCzZAt74PCqOYYMul3rCqc8Y
VmqMa4j9ovigg7ObZcuTmayfSbONl37G6R1rOChwknkO0BCIkkuVb/Akn97NUUJA
rYo8NDsjNsQ/svOAxM5qvpzXd9txVThzjY9r2QwLJVd8PFhu2xw9IBuRR48MLkDS
9/8Q3zZr/z44PsbCmEf8W0hj71+LTPC9mOSj7tCHlOpC2suT2jqMD4EeFE9Dz/sC
JzXvGa1GuSAEsFCNFN5UZA+2e5kJ/jHrNXtzSdMJC96A/24C1GlNe9E5AvLowLVa
Ts7uqjjBoSwZLVqfpAb15C1et6l4fmYVVZ8WTO5cPeQqUBAnDY1jaFJOiUmV1lpG
4hQ1C8Vv5LsTfBztrXhapvANQ+3THh+qMbIQI68oBeKGgJEyY58ZtIWNCmRXhSrk
2lHewQljVhCn6uSjoOmMhchsiP52hOTamkqRmr/UaY7TfWjfi5FXE/UgElHNUuO/
EERjQnn8GZi4fmQsQ+SAuCIoNmi9zH0/15r/de+cPBWoj9NaD/HaMi+Vlh5K4dN7
z++ZPK+Hns2bjKDcG/s68dEqI06HJZbZ1OL5kQQQSTM4FEIa1IMovIHAjLHQTWfn
/kDZe+AdBlxAYIz8VH7lu3pFTU7HnI4X0dBegY8BOEC2Waqt7IpwEZ8dTLkTwAOd
tVZCyXF+YEBlXZsneRuTCWnqnpsjHEbuCkUJIkPJh0WfaTQ08XDDO4qtYJrDpKqy
VKTANeP4n9I4UD+yMXChllXFvmfl3VEbu+x8afshbCOA9QFYKEcChgIpiFtKtuoB
KttI+x/638EYX1Bp6fKmHlJG362FPd6prMYmfYaa+r/l3s1nGr2J7NxTd3/K7468
h/gXpWhAPiTJxbdXobzbaTDHz3jmpdZOMQ03H2Y4NvalpEtbERharrE3W+kUTZ+P
BADiBLhKTFynkMi0O+dKQ3D2pW3Fmbl1TDw+pXRA1h41zS7RYGNtQ1aa15vT1SY3
UM4L4/f/ZXuaz81oUthfqTPXF/ONVIOn0CuAw5yrz6+aXfW71+ZO7zdP9y4TdLLN
q9KRbr5pPT2qMU5nbQ0rjb2beDVu1XbpNB2l34/R9RAhh/N2fu3CCmVQn2w/ytOF
di2eCX/s5gMB6RwNCLbe1JJJHqPy4o7l+B3MtTcMlo2FzgHRrZdV5I+xkpNWrfBn
IDZFSnuRFxBMHxEpO4jglNZrKbXfmVdA/5/zvoKfTqegfa/mrH2M8lF7Z0T7oo/a
/TFhboudNPen9M27KwodF207WDMeYOWxfCTQZgjT2azT8wgeDmQ35vqTbjVgM+pR
Wzjz9VG6go5uSHWrKGnpf8u+X33wKrlg5ggKBCVJT6sbW7Af0+Ax5/JJc8jYtgyt
yvurovUmXOzn+2fcpGWbUicw0O1wvUDuxR5VrtUKje4VkYSkFBgKENgyJzWU1h0k
zFuYa/WMPOX1eOxdk6OWt1xi0wiIG3kVFO67OZnhvQy6j6jSkpUTzbxek9Zsdk6o
+RBg004j8/hsdXQaSab3yqxyIoXSWkwK05ux2liVwTUUTThz4TnE49T/ST54rVEJ
MaIrCFw/lt5g4DLTIdTMtgRgm+RdRgecMOXjVxCxaCE/v104ouvcgLZdELyNZJ6Z
Lmw5vCKdeGww11BTVLKdpTYwODBrVuZCZue10t5oPnJJH6IzOctyaohrcqq2XScl
9haRBBZuuZdzfcOEMB0IJfFKTx3TFmOQu5dvYAJNJgHijo5WAkvSenEgHhUE+36J
W69/NmbM0O3LKwADqsSRQwMUsw1pWyem6mPpAI5XKT1eCdOEMQs14MPXHKRm5yUH
6E0bLG+wK1ZeyYjm1JQoIvf1DVOTmt3JjFPo4ipXoQCDriLBvRrBxirNSQLJWRAP
085Qd6g3pmdHSX+bmr93lCUVq2Fxy7rp32F6lfXYu/0NJIaqv/9bIlCb/tfvQEth
0RXwoQH5fbdRhYcxSMN3Ty2LKYQc+sRA7eZoyfs9eqVgoRk78W5T4SQO9223N2oT
sNy5Dmxeb/iQZwVkgsbTBFCN+Di3G3xjwhGckNMo4ODNUHjoRCfiEpD5i6K2/ZGk
60YtOC4JJL19L1ixOrWFAPzBI9zZEakYWy+w1unstm2qmwA0YzGBuWrNz9Etgg+j
Op7tgSK8K3fZ6f6UEB7Bx30LjAkO6IEyCU5PW6YUHM06pnbreS7crg40udKAD9SX
9AN6gTqWffFWqavNo1CLj9zi+vfWKVo96yTLXbGfkkDyFtWOuvWcCCZ4bIvGXo+O
u06CR0paor3L583kynSqx0CxT43DIkmndcOEBjF4RrVJXlKGhVZk20R3zckz4Vee
9kHRqDmP5IeYI6zRWw3BZf1uS4xJjFJkQKCTxRsPXZzEJg6dU53exKBkJDUyxP7q
0qmj7TrkuYsRnWv8p/UispVSEh6E+PlQStqRPzWA41t3zvZlcMBQpbJu8Mww85IQ
c78ARgti/HIi9szXdrC5dAxreWDvSot/OLe8PkelgNc18GtTPFmou0zkDk3/AWoQ
HUr5rTzypS6P5I0wK5NJN4ajCm2w3XknkdyYZlS7rYCDZj4BB++nJW2PrkEN0Ait
6k5f2SN5KHBZsfL9AvaXx+9r/Zde5+wdSbRrrsDztLELKfs53IFL/uA5/G/815hL
8oShZHTIgacm1abjPgd2pLxf4WfKV3MQGNnyKVqgHLMQuJBE8twGj0SMPQ80NtLL
E5nx/f8G2UrA3pLofskiJjTidUojs4JjiQQX3EMRxlTse8ips/ShdeszRxMjsXFU
zPfbnrrOZkzKi4AuQBoTK+LBKZwGidVnVMKOTSamm9P9MLlcG90NiDb6osOGVUgE
vDvEn7r+XHxTrNVozXmzWy7wWOPs+F8LyJ/fFeLb8ZEE1dVqYdjpLrhmGBRXp8JX
/kP4rrZ8Gr38wiNSuOAj607VCTcMvRFvY4st8Zjq8zE5m5KVWugq22gqhkZLQsNp
3FaXM1UOKrHNT8ew+fzeO65A+X8AMEU3JM1NZlH/ms4J0mFSi76B+/WZKp3azVku
As6EcgpqKlvavYRLD9sSRnNB1hwEdWy/CPiYxHW8pSUXHjVN1g093WayT7Xjxt11
V7/4gfRksN51OWF4YgsCxadrghCemP3USQGWsc/NDheboj11xKQ92ZfGH/PBKLn2
olkgyIZRie0ADma3SoFJ6dG+7qxcr2xA5Ge+7LToZXzNGwsE3i1bA3REWpH1lQP1
lHl5kIif/JF81V+nc0Px77FGmNEjgfgwjrvISAzOs/zETdhjjhWvlM9TS7CNgqu2
Qbzv5NPKJFj5qQ/16icZA2/XBTduu6DRXXR7kxM+Ah/p+GaNotxxNJs/H5KWNoWi
OgcAyk5v/MerrpCQmVFOSuCshZy1BJ0kCNq1+YU5LZNMCZFhES9MZGsUzJoBFV8W
hRIECYxBNvfNPY5NMzdzZ2JoB6Z9iBQholTd5N2G0OqyQrfxstvSLSzEF84JNLfA
ymQZsmgzrzKAn/bou1BVAXmI56nJM+L5AZyqMQQAENb8eDvX8/ms9iFzIVVoeWGP
vSqFKAymR2coWT/EEuH01ctE3X8qQ8wv2ItfCasiPuiRFdKxj8we2HVWGVLXRs2P
0jPnXsJ4LagwTAkbmKzOUT3LckmTqkC//mYp6z1Lop4iFlOXhAl3TNmRPzJiGexQ
hJ+ysid8GwsVHRUK4NsCY/I9zceFqdqzulWzm1DkJvu4bO9bWfghDb37GX/judqJ
B0fIaGwE/bG2hVwu9+NuqKAYAXFwwGIIQRnbsTH0gg9ntzYCeq2YW985nrvbRDQq
Dhrf7Ey6dmzx8clkhk0WwNHW5iXsRZ1ciGfZaHsxb5LFBmzUatCyBX628QzOz6OR
pXxL05F/3omU9h0kNbx/Sjfgw6rvCfKSHlPpsTKFQcuXQz1rvA/7pp01VME//1Qx
K0H9+ACWrkXGsPbDpeV/7j0VMl75Fn+0kjFSnB/RVx6Idia5KoIV2jXHzMLK5ezs
/2VoTFd19XFeXqpK+HyIom2WTGG2ev8hUwX8hgyOEozQjbDaOsyWSXqtsjji0PWm
cZIOO3+qz1lEY2N/rVrfK4x5skZ8pKquhFY7qcd2jo2rzXMlfuxVb37GXfA4WPFm
1UFuyLnj663Efl3u784tBAdxU6WambMXOVVG81cyf0qlKzSAOCn2qDt7HiussEop
qaTpzkW1Dp9NXRGUfCJPGNNMDOTCuDTtFKIgchOCalUXtFH8sd4MTx3iCb0wZZqO
Ox03wOq6pF27R0+NMJa7neM8ytOsQ3XTd6H2DwQoR2dC0ej1td0fVY3baO+1LGUE
588O5zCk5ycQ+aqCrZAFSApCYut1m9yZOF0UeiTXokkmgBp5PjGXieQd0/6PQIYs
NnwIDTr48q45sdKeuuPFRDQHe2BHwmZgRMkGdm1emz+ZIYWXKn7HX4dOnbUFRU8N
W6sO0spYOa8cjhvGLFZUrHkQ3Ok5AcK+Mk9ww96y5IpQe/KuLKKFcycxDGMYP+Gr
70Tf8CugDqayBSQLrcm352pvkI3rmbxc53mEsBqFjYFFjd8/3CMYYnVmx5VGrB2y
q8jk+wZTsWIW/N3Mb0AkN8ZdTmJpkK3X+49yTra3bEeJqYDpBw1x/QgKRse79Mcc
IeiT+LFFcEJrg/hdlFsQ7q7R2R9kmuaEwKfrAS9R2Of0EAt73ycRMzCFPdKinycF
THw/V+zdj9kZ5k7LNzudHU2joEtCIKF38P0/apdqwgnqZxJd4JSLPodZe5SWj9ik
s72c7TwjQ+R6ZELXRd+sw+csrBs9boQ+Bdy3Fya7yoUinnx5y33/I3ZHqsKrHzN9
fiGrogWI7KB74dI8pvQ+/Qwt/NZ5447LUiwICyMxXdW3XpZU+yw7pQ6YtiItuiiV
VTVrPpyEuvdFJEy1sLJJJzUrE1nmh1MHvPOlVaU3Uv0pFTy4ILIyLl2Qw34100pM
P/oJYLcI9ZusVaJmkCImFgf8rhDvfHNNw8LB4Ke7/NKPGOffgfHXw3ZXCPHQox7h
EbPHf9WycZ5cagKSYKlvPcBRP9cRQAYRfnkQT8cO0ASIjUToPpMwRdEtIu9KgMWk
MJEhIgOz84apvUx7wdtoaVFIZ9C4x9ot3SEQXRmD3knaPUA8wywphD/mz25EB8Dw
QtcjmvMLNVy6m/7FDR23kiCVJEAjUBUEDOfcVxr+FKVocfkVVmvWxFhYSdGlRhiX
jKo8PMnBV7mryj6Hc2EiAAIvgIU+K39WbZxe0YhDEoa0uTs4FbiYCQwQFaICb0uk
31Np0fixQD0LfauVtBmK7msn0rc0sgV//JMmuM/4WOQn+PJUd9sV2QNLdQ9yBSuU
5ulJwCQ2yCgrdeuzHhjxJL7wAq+JxGjE/2T4mv3M2tKXEKgMvHNadc29aGx/gOTR
x4VukKq7b1fq/btS3m5Us2NvK7mKIS+J8q23/xej3ZANuFdU/9f3JISFAbcMBXMF
vKFFngD1PHziKEP9eSDM2NVUfNUfibqdmJBrzqjK/yEzn8Ipspy/xfw98+ZYmKCN
earv251uz5DTN1/AwGzIPehjtUxRiRS8vt+7Xq9BQ1mTodAH0EtX4Z/CMgkCkwYW
7FXosJdukoVh+6GCjnUUguJ12qmeBMxpm2yAImf1B5HwWyDjym1XrsE12YFapYIG
RjrvgE5q198gtP9ioYtlWBG10YvuO2HQyNTg/8yFoso1NbfPHFUeQpd0B4I/3ZEN
QWtpdSxKhAZBxd4jqLB2592w2npxTaigCUcf44uE+Jggt/kAQkPTKXfsGfVt5/Cf
P9yufabQuOq0kF5oHGd4dnATRNsvkV4zwOUCSnys3YN5rK4KT5qcYeBCR23Iu1II
HYieR0XMEdOak/T9usR05kWmbDyVAP6tjD0PDwdWtJC96K3jwzr4RUyKF8cmIyf9
oNenIcmHasYCSzGLD+XS0uroh5yJHT7A/fH1whZOJ7ONceXwNy46TzLcmKhwFAd6
MjQ1Al7CBRKf+8Uw+Dh12z0doLhlsnfAGV3kl3kDrRrRXaNKQoLKnEGV1dLBhnhd
/oh2/em7KKa1jksptXnhl10Cg24g9tmLUeHSptMCLcnx9P3DNRS3gricooSmyoFK
YR26ZnTJ7lGM3xSQ7oh8uAGAjAEt/iCda86Up7DtqXvIcnT109qWTQK/C3oJvbTE
era1mjU0shDNkosiz3mCBKaav4rbwWnK1wGuxqfGhV6LJQguEolFlj/LHvDtNiEB
zs2sWOR27oQ41fWc66Nv+TQdoVYPnMK39uPplPmiMi9mwSnCk8QfgLt+xK88KfRD
Ae1EC05X8ZmDXpyeEbLrasYKGIcYa4QBNn+UJG3oWoZu2eiEC/d2DoABqRCrIba6
Bn8oSmxTxEffopBlRVUl329cuMWKwdCoAloHgbyy2Bcyo9FPQDIAQE+oJ6FNWq4u
1WYVTylGz6DcdvwUsTCTJVDrUpr2aZs0jn6k4qz8v+iJYmOpHrQXD4TGP1JRf5AW
RwRRVu2IXqC6+gCjP4/Zr1NCItEzZdbq1g6jHDlsu7qIju19udvE8/SduW5EQYtI
6JZC2Wyhoa4rWHCJN6XYgkM1TWVAbXsqrsG4vuAJyF9a2g5IHLCrMktl6xu0FBSU
SxN5e0qDY1fX2JKDb2KjUClVzLOC9iw4WGI7dbAf/g9DMNC/ga09Ry8WRTUefmzx
FpNiOJTB06voLAj9wBKpqw==
`protect END_PROTECTED
