`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Db4N0zEb5tJpC1MZn6uRC6j1KnXcgTwQmeddRQlepjq1twaDb99Msy6DLaCmhtmi
ueix+28xKPAAFSis+bJg++XLAhnxng+BWPNc0EIZNVCAhshcFg4UpJcOu79VuuAm
jQcoEIKIGt6/zjzVc179iVpgTaJvZsu6qMZESpKDao70/e45rPriA38EepFEhxmO
Aa3NllBsm0yEkcvPtaWsmANjcqBV1iOaPeIyV7f/JifYmV6TEseCzPuPLJhV9qf4
029uNBO3G0oE2CRI+3/xppNHO5QRB+tkWMiT72TCG8BYj4i70KcMZK5MEtD512DG
5WZ3bKoVqIntCfyQGWY/nfprpgGNmFQoU1T4kmawC2kio8DoqjITDUN2gt+OniE5
9HonR26JJrAhwWBByEUe+25cq1cVCpAqh/22cVYstw8BYbbddWX5afKclRPKxFGu
MnmtSqJvLF7+Cv3Xt3/L//UWzkA75Mo4lvOLNaguw4E2O2QdIxPhNOa4L5gtcshx
Y/JGC7Lw642V+KrSI6i2wLrHudmJs2nbY7yNK06/9abEikkgsD6PUwjCuBSOndIO
VLkPLLoLez1wV1O49Np+D977yXO/Fgg6QEwTltyL9eKS4PNr8hJBXRex9YAlOC+S
5O72vcUxzALgenkxFf5jsle66Nf33Khn5FOjOKz7Tio=
`protect END_PROTECTED
