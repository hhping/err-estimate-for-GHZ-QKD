`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qzyhl4J6wtEdnomFR7IzQAaOx+Aj6u5P9k2Xqj081Roa/V/eMVZfcbjLQoqme3Ie
ssMpCJvQ1pK1AgSmRiAQ3dgUtZN3+CRjWt4l3zWJid1PYEf4PxMw7iUtYAf5U/0m
WLZyUiddZ8i81uL9XjnCf6GeDPrnFxqPZkSZkB3cjoXKyLIf5MjVwVPpepfZ+c9H
Dj0oO7tBu1KQ0bEFAsVua39AZ9oiDxrqAlE4mPSOuJ3Ss5PGLaGsy+7OxjnZPdcL
b7smfeBouxZW6LgATah77P3sbjdYhNOkKWlbL7jBz3xv/Q8LPiNOkQN6kI7naUf6
0DljPMoBj+W+72MfsokUNV+/OExi3ttnHbgZyAduAInAwONTriCJFB2+I9RMpcZ/
s6KnoGhtxkX2rFJyRTUQAACNnb2Y2clTSs6oocPKojnCToDHsNzz40BkFWFEPWG1
UrcwJslttPDCrgTSrF7ZcIvocz7G3eJGNVXnnYZMMg8aiMYD80bbtSlBPnEhY2hF
UhtkvnL7NduPSdBfEWI0biAXrwjH58hgp29xF4J62cGfB6kFyn4ONnbfcAuKn7bv
KNmGPArMZn6f/ha29yiaAtv0rnminMKubcj82a6+qjbUku/lqPp/8g75S7RgFt+p
6jPa5D2vorriiOofWhoyjuANOgqxExaMwu7I4+9lrsBbtjhXQmdwImFObdzhDumx
Gtom5VfmfF1JTQ6eUX8BftSVJJEFildG+1QD+CrqVTL57Lu8jmv9VOey+iwjr0w9
qxcfAv2imWmTJpwR/HAQxhn6HvbzEBeCaAkfkMcGK9wKuk9L7rQg1MRz6A8/hNrP
falvcploHHf7QxweZI46LnltQ+vT+eCT4L08odfI7Jw9vzFpMw8467qH6LonzOa3
0LVIZL8G1epE4RtT2R0RDya3PEgnPm17ww+UR6qj/0oea48MZVQthZJiQWvd10xW
fogkoND3LY+Z8LwpZDgvPjOxQsFl8YgZb0ZD39fGAF++lgAF7CRY1J5yOXAHXkU3
lEwcLqk2kA6K7aHRskpVkZ1DtQy2WAYal8awISfX46YkekqfX9rGT0vfVlJxxQ6n
TgZBFsqzHvEJ1nER1IgusOQ2VT2WdqIlY+Tweo6GQ7no6zkzhxPzMK11h/kuxejg
R5dEfZWqRhzggDWmlCe98XYgsKyfeZePZ0kUpGW82y7fnoV7nYfXCwG4Wur1EVm9
RaxfEKTSZRf3p4cLgZL08wD67e6tRYowkd/Gx/asPIlg7NeeyToTM5vQSHEZf/aq
XTFDIs+F6/eIQR+9DF2x+cmU2e1bBdi0kMnZknmitnhQV6Uato2zUwUQc9ciEAUB
LwoOzfLIldS5Kgz7LId11b3wrWpo9YfTZ7JPEKtg0y41aG8L6xry768T1rzEgPiz
4nPOG5Uj8iL4FcXKjhXn9Q==
`protect END_PROTECTED
