`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
asDFWy7/Uylmo4TgwZ6F28QN12FC+wkHSE6rXHnx3c7GISBMte67mGjh549TvjKJ
/STOKv7XqI0wUzUnGiC7pWA3LaiiLCPqsCzLCxieEbvaqB7JzbrqZmn3qo3rrFQR
g3KULBAT7ItxYNJQ4SebmCs6MElG/IIJxwsfVIrLzhhyj7RD3KAAKHwyXL31rQCY
rSE7yXdgBxXExkg9Uv92D/tKWR/wrrAuu4gZccd8n1m7pVUdVUUvhsUf70deaIcf
zdBsKJ5ZtucwlGhFwww7nqTrUqKU3nWSaELIBK11cJ8cYmc+XjNdJH49siDtMPmq
V5BbTH+BmmFLf+V6OtdwYXC03sKuqdhipE9NkbbcOKiQiUwzch0XAhev5TiL2YWG
ozQ+roB1K6WbwHyCcgf+CQo0h3d6DBXEjFHlqNohhe4YgXodRLQiEyqJh26CIkjw
48WUUjGDafVMdTOye1cdCABRrrjE6BheuhEQCL2WsM84CoLuLuwcXdDq+CTyM8aY
daypVilzztbAWHsHXfpbYZD7pvGD3BvH5T59wf0EwTpsFzz6CgWeXC4hzmxCJS3U
wLF4R7t5arQ6GbSQrzuTldKVrLQIS+A2mABNPWoFMf74oQ2jAefgXyyb5kCsCopE
3dsOmkIGd2mD82WJrzeo4E+C4EZ8Ptmw24uoC+3ZwR5EZVW29+wTZw6tMLZiYx84
s7YJqpHDVi0IZiv1fXJhp1WdGsMPIciz38pe29LJJglan+9nCVPyHRH0D8SVNyXD
tQgr3fG+6ByGTWwg12V+lw/Qmmma88e629FjOuPoAdZ3YK2c6qHTrVmHyvvjP4VY
XghJSZj+jBUVA+yj7uOTNVXtsOClds6v9q1qdz/wdkmi1u1TEcfiFXem8UbbMxVr
UkIfmalKX05Bdp9dT0FY4tF3kPyV1bL+F7mxnmxREnXtbEedTX3mh+dJdDNubBNm
zkcbPnE7zyJxPujw9bERM34YVR+gm4iUIKiKlgHFb68AYfhzznkLJawOj2GROJVR
wM/Glk2/y60Y4mTSpWCUmPtD8m2mbnMX5w8ECOoBT6GZB1rkJh84zMqnD8DOiL2u
TAkGJch/c8L6Dvb0BBbLTKI+l0BnPSZ0hz8vEM1RHWgpOx02L800QUVocsh4YDkb
3ym/59KUFkTcy78M85kuCIVsc7JLCK/CvYuGER+wwSI9Na9ICZ5DTzjnO55jZbtC
RR93Y2xRw+vkEXDOo8z3ZIOIrpeBtoAQOiuVmUN59hgWJVq8eTD8bFbFEFvOyQp8
ebc/aqU3a7lIGhBYe5ZBJFnGmYtFpFlgsUQ68aJWezoR0amFA71jp5f6Clvxwu6/
qlaZdIaJbtvh++ICP5bpmTtCccoYBotr+wyr+BGctAYLUQBvTH85+9q2TTWKjysV
2VRyHgiy0XBEHkvBRH7/9I/axF1engcfBk1hdusDXHuOnZ0PSlibVu9Wue/laBWt
KLTmI0A9jiS81dTiv6TndLRAHomKTN7yTTnv+iCBu/9m09kzLGY04jtBcMfx3U9K
8GiO9GZQVSZimpw8avKKVjmsq0MNGck3CrdTeuKmwT1RqpeLmaUOMUtLMsAN8DRN
Rr5MpNugof56GF+BRtq803UOZK4aaC8GG0KPfIr7LmOq3VmIn8/kMca+PGuLzr7n
+7X1TV0zF6nREimvRHXF4wJ8YXD3/yqL4YVXtu1kmvLMaFeBywkxALd8rba7JmCT
uVzRLIHrz34/um5bLWAn9feqwm9V+4K/v13mFkpB4sBg188fA3tXpmIfYT50cth9
Q0veS/kntVAZSdjAfKbNFvqji7LCxH8idEdnGlNDX/6sf+GnIiLaOfI0zzCjwph8
nkjqICNm/1A86BbCIN+GlLI76/qr6mKYDOuk+TRt6AraE1MLQECkklYU3PQFwMCj
0Z5zh+IxkVxUCONCpKFAKFrmgSw8DnwOsItZFc651rt7Ic6EjtQBVVxBzo/XXW0B
6lyXPg7UCUoJlhaITC91/ZY4c1FyBfjUhAsekdTokSlmfVMKNeznhEDlyztV+8XV
q/JnTMbUHYk8NhHckhImrUsU59ALu4tqP8TkB6GH4syAH+AZEeLTYRmpGaMpSnAd
fv2GKSYDu6pMV8PZ7mSLga7Paefgu57FhF9ey/c/eJ3SbLQuf/4D8iRaUaM8kYQ3
IH+6uuPhzgNPvVWbbErX60XI27QjnfFvx0ppG1VxDJpXGZrEgOhSOb1rsZNuYtKv
8mMV9vb0rFd05+aRY3PtHT8ZR/wF4ICzw7hyAQsA/hVFkzTWxAQdGsbirYVmY8VZ
Ic2RP8VmjWWeQP4MjAMR9ZF+9FuOlPQxWunK7VkYWkt5HSoW3Mtaikn/0Yen+J5p
67rGaDLT/0HE5R+MLOx40GsePJcCMqxLVFPe8Sm0/cBeyzRB8/R5jS4X+axCHy8p
F0vDYuELIM62ZrQOk068DhWqe3WTryadz2X43QPRavkAflrE8ndNJAypBq3PHCtJ
KumkAI3C+JWksPYNuSAFdqnajQVxVJHjdhXzJgXt7ZB5DAY4+QX5ud/+bA1EXfqa
Ji42qpVni/Hkhta8S8AWqZqzKQ79iOU18iEOQakwOK0/OGofDeJ2Dy8hJgOgiVYi
zVFvDOo9EJrmz8gFDqs8odqhoiJ7aSoI8QMzP/z0OzriHQE+GfBQwbAgpPF5CZR3
UzWh81VunnRSirJxD3GGVp7vxYg856LztlASShvp13LRRb12HSoOKzq+W10XukdD
dixQSpNagiWVEonrspYwAHNe+cG8o4MQtXgLEWKJsag=
`protect END_PROTECTED
