`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nVQQRX53O1e9vsN5YIp1RVnGogLAz7UefMfiNqNFM1vBB6pv9/DDtRUX6KECcxWy
q82G9efyRVVqBAXXfI5RoiFuTzyMD7VmanRP+IKumRpSRno6COsmjHfpjcWHKKKd
ZBj1rWLLQ60ZNGb1huepXAf3tM9inrqcY4LFVxXtpbq0XIzw/tPx4+BSInYXpIzp
726RlDSjktZV1DlcGRvLn+uOIvWOp41wH5xr9uLQTMlWDIdrj5KlF8XU14snpnOc
e6J/VMxxNJa70+9uNsz3mdC0PNXP7QPo5lyCV1Fh6Sufp8t1bbel7qU6u4W/evDp
OdwxsUMJAnCyCITAgCtoHBiCRzEzWSGHaOw52pQf6mazJ/VAtgbSjrhHSzyTvg1U
CLk7NDKfePHU/v3FbKSbVO3/bbceba9NXs4btPihJZcpXYROQNhe2dun4M84hxuK
mgy1Z8maO5iDHUQkoYtSJQmtbKdNhdHrOPhMx+Tp0Ri7TGtnP+uftzs2t2hQRgB4
Fk6yoKXJ3MCJmLis0Z/W97gJksv5fxaeNii92uxWpBbz33+V7q9+ff82YGLz+qL/
yph+0uNH/Lgc729Z1fnp0u/kkl/aj+ErjIF/b2+0J9B6pmWqyO/vQMdpo+z/Sbxt
rq2SW5rdla6rSZmDr89s6ggyqvkoY1EioCpgneQZRSPIQMeCHVU0V91o6pbOodqr
3QqfyhDLrd/u5N5JyxJRfbxfe9fADAT/yfuvEq0St/w=
`protect END_PROTECTED
