`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1/4fZeLfDB9H14HXX6KQKdjUsAdtRosUBtiU2iJpVvoIZP+bZ+mxxImyFkPSqOm4
HleEotG1dCVg2WDD6fNXUTe3a7ipk4EUTqMhFds+qMY6sYCPBFni7SAEI68LQ6uR
lhkPqqrRfAiLnkcVBUNIkiTFYIcXf7pRoayKO9KKpNLxDJ7+9O0YapxNKAJkLGbO
g4OvjuCq3CJcXk/qRP9lXWZDTCfKerL6fkmwhOsuyZg7YcbgXywlhIZLWs/h11fY
7VXrfJ2Y9y4U58SKqS+NdWNaOI0BljMir84dyqu926JcGyDeFK4WCMhL5+ilJNp+
QIWuXKFm5Nqnj56BeWbnLRhhn62ScL1VlnFFD2cxODIPwXbon/t4rEu36BzatjQ8
LS0bJEkRRxB82rR9nWGQN/6OOQAJMCucIbQWuaTOznuz4oWaDpsu8RFYkolfsBsV
h/SoT8tkjJJOH2av1NJttAlvrzOcXEdC0TD8GW3e4CSj1MnlK40cgDK96xTZz4Vn
Do/C+PlZ8Dz8KIXkNfu+upVFxrLypaKLoeN2Qwuf8vr9h4vXF141JyWjPovT19ye
W2Lc+fo+9Z6XnW1GsP4VCAKUSyYePwko2XeOzEmo6Q3vYmabVRfVFTcIiY7PTno5
QkKx/MTCEjmHqp+DwA9flRkegY6eVhwiKSLHQ9qaiUJM8TGoezc88SDGooWfQE20
QxEmp+UTqb0qm78+NqQvrDW+lmH3zvs2D+XDDFQL/HQTlU5lk3AQHdGMdF+zEnDf
IkZlEAqcArMNsq+5CLGgY0Yd4JbLT/A9oM+7LTeEKWerWo3b9cLYSJkbOICSSJC8
zBVTZnBPwGlytQ7e/xTk975UWqGNUiO/R6FiNNSfkHrpbGdTZ8HYxcCR5c58bQfU
ozq4U4f2SbUzXNt7hNgpGn0EKVnbvPjHM6ApsjPFHJMdlC8Lc7cS9EZD0RvXlwQh
HnjkaD8OSkzbpdlmN3j2bI5+XMVrR/pBL9G4Z/qybNKRvqRBjFCjXS4TPY8835cG
XT3O4FzNM1uh2PaTryvhZpZ2bsLDeJaklF8f5S2ylH9u44PS9qb1YsubSlcjbYr2
fb3zB+h0iDccxELtJQzX7cvP7ZIUuDjfHme3/SMR4OiCBmGIrbY3s30pa1tWt+kz
veTUFtgynRJ2rwiJoH+dz6PwltIjEm5442D3lXucdCaaJG76GoIENVFhDqlec8zo
9fUAekVl0ks4LAb6DqBfrrO5Tw30pXUwUHDDSMO71H6+2f5FqN71vSq5LfOyTezV
hvUeKNFl8ZTXZXCFBfzsAfmorOpHKAPH/pXi7t+rWu8h792XdAfjBUGwm9/esNfc
ZrduE8do/+OC/YdIbCFKpZE20X3nFtdcGaIICpr4NKt9eGDAtkiPOFZ7UyXXL8j7
Mdjuf6z3Lzqcolufk+GUCg==
`protect END_PROTECTED
