`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m1e2Qx6C/62tj/cOtcm4TECbzyU/RSI/+66qAYNJ8NR2mL1Zpn9AjEfqbN7w5Mgx
aBpnhK7wmplaF4KZZgtOXrT/AEAjtt3vg7gP5rckdOd02toCkLLRDj/A0JAwYbaf
ClqZxmj+lu3k46PATrMUOvGTd3cu9DTG4aCXxksRI+gtRBw5xIpz5ZPcNHLXlkei
Bye22e9N/YKJS+h0ciZkwtwPszJC5pj5THokZyynpmHHAnWdNKjS9nPDbJkf/qiU
M8GJql5eysPkWhHx9gsFhjMsVz37spRnrdwjXE40wwQ=
`protect END_PROTECTED
