`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
meoX0gKhCiN5z9Nft/7pIwL3H9Uy/r5CbbReqHakghJdgvYS/OGQ1ix0w3Zr5YDu
oNFDNBYpzxw/QShIMMuFp4Yb6zPEriioF4KuUsCc41594A3BzlU5A1v+fSuifibM
yFva+9eFQg/XgngwQRp+MeV9Nw/e8ZEXyXjNGRG2tIHR9KMUTjCMaiDZCA0iDR9I
K8jzLFi/7GypGnDFXmLPzB0Q28qQA9Ca5DYc+hpx3BX2PxzdZFz1leYtFohBKq9N
Vuy8YuwM41siB510wXarVrDTrX4l5RSXoAp4mwl4jdYK/W/y+gatjiNC7YE+rP7h
gg5AVLzyjkIdv3mBI1CRQJPqmy0huxIRZUIb2sdzjAEkxj2O5X9x1slpDJ9ucb4Y
B59vf8KHgxSScU12avsOZHMcXGkxcktuEEkP/sqP8v5N9Z6nrSrCcGQ6lm04u0Ug
yqTjuJD2K7Rx46d8JBNszd29VoyGGf0BBJrQr4se/9EnReICNAftfutjQavFTJJ1
Qfdx0IUa222J3jHYP4PjCArH1wAdi7ZlD8JFmiG//Jx5vcXE7DD7B9MvlIdjRx93
AM5CyW6ohn0swdwdFvnf/YPnYrh326tb/COpsmWV6Y2MAowooETlf0HQf884/ayp
vXG+Wy29Xu5MOIarQkus9KShE86zJB3djtOdUWXjl7rPnnCMj8uHxS7NYO7I3QFF
76d2zuz1TWjZyfrzn/pi66bQe/iddR9Xlh9a6zycDr5QWHHCmktE1zZhJxSiwoWQ
5Bfvp7IepnRCiFi1rufP57JZZMAKvETFTi9qlehGyZL99EVzm02W1ZSSwXkwrFy5
twBLR/2EBeS+kA0tyurJiaPKEZ8OWhioR3mVxVGxBBncnhYIPt47ZJvqZ/4UinSn
gwHXEPR3/USEQLUeRqSQnKQ3GDBMvWViQXh0yXTKuIVDGYOsTeCU19aNdZYQhvjH
3yqwMHgB9T5ZHyNBEqwrykBQZQw5BUwRGMyrzTyiR2SuQvbsci+PRBq6DfSUcpL/
BSTizCqij1lNPF0NwioHyKbIQeTawdsgOaw5mfWaFWE+a77cXLOOiIJBTol1Su9W
ycVx59kQZiLmjIj69LAG2hzwxLdIF04WDG1raVmFvxyYeeXn01y4afscvxK0LVsC
dzMF4DIAJAyBKcapB3vcz5wIozlmPLZx+P1oSSH0kpNO9/h9fej7NoF20hZSo9ZS
4K7UscQagJ9JJdRXTwyHGMXrl07pIkbOSbtxKIlQydV8JXOeMialbNQQroohR3bV
6eYZ0f2HCQZphorvYKGfiyoDW33iriwDuF0TQEEJtWRaL6YmY/I2Tx01nNcmFcdv
bk3V4971YDWM47j3Pn4ElzyQKzVsea3yvOwWj+CUA9L8ixXsNOG4ltuQfXXRHYyp
TuF+acN+zLt2JwIpxi4U8VjjH9Evx0yz4ZXyO5w2uQ1xjgeLvftlMjJ5g46UsQ4a
EMz5WjUUhA4Mw57O3TNdcA==
`protect END_PROTECTED
