`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bt5aIu3ZV9r7Gi09qbYRUAlHxrLmEdlCIRCeCZHkY3eP09yyAdPZ6eZkgfpgFGbA
zqtYOF+F7FYlKNOa8N/FjF+l3rYN5f2Jqa0id2s5wfhX5Y2b3a+2GUGiWS29Y3RH
CVPjJ7JwIB/CaX+XtGbiJ1w8I8zQq8paAqo5UbHdEuerdLkchckZSadBsPQkL7ah
pdBtkHFVnbpaBVu48Ap0Ue6yPDKbLJ2JIaWZFh+LtZ2fOmNdPs5PD6vYgXS6G2v1
wGiJpdWI7qb9YhpjQy1qnAiIpWSfm8nNBZpoWkSXoP2Slvic9rL8SvDvWc/vkiq1
LIpk2AQeNe84xJXsE0MmBp+bGOmv9sjsrvQlMzGsmhlRVBZAVn/p+Ok+G7cNtQfv
An+lsBUpUoQAUbgKSN+xeDWTkHFFL7fGGrJsWutgqI+Q1y6PDdqYL2MCSLdP/7hB
NuqlhuZjV1LYKyMSFjy+sDjZq31F1wWSfDmTlBaRWv5+7q9rAHM2qas7yQKWGgCu
PNQTiIPBJr3z6PnGs3ekwXwMmP8vOA8Fn/RUZjYOv51X7VRI8MfiU3CAAlipqsAD
5OTx9PLG6h1Gt2xNkClOWIa6xkiL5B8TVHxe6xWSkaXCyUzV9IbN7lRAnK2rWNDs
tglNdRkr97RExJh5TejrvGtrJh4bU4jqF6yU9KJodDxSshVxy6AsxmqooACwiAvi
wOLCwuF9QwIkkhnWmQyy3RJQvgQw0KYkPsAF5nuEK13MUpB2Wfj4bq+O85WN+V19
9qsIeZ6ylgxPxBKrh7pb/KAJY5ReXW5dUg493Wx3CIN87M88jZlnoRVu7AS92kmx
Ob/Nf6JU7Zb+TDEFzje0BFiSqg6VaC25ERD7cOLBVrO/1YWMSQtkDSolKaWBZYj/
L9+++xRvGNIlODA+GthkiqxrSsn4aCfWANAWiqPGqQkG5KeIg1Qji/6n+y38DDBX
qmZ4hKHXDLGn/Nq0q9Svfbw0i8AAA7IahJeK5tbu8eVW+D7bvdY3TySeM1xfk38A
ygYgoOKbK1TV2KuoSxqG/IQQljI6fgF78rQ3DoK0JqjpGsgo5CC303kPfoYrCJo3
WL9GW+rHSrCx6JpumcCa/co7q0xpWl4IxnTAUKkhsLKl5gadFYeE+TPjAczq2Pht
nq8T8yAaNtB0aclkXUoWGQMWtUI75REGgKjRV2aPaHS5FMhjRl0++EIf7lryQ8po
wSuuzXXA+4otZepqSa2fsBUU2f6N6WkfUlTs4aQWIZD60el27cehY2oYJWIvU62g
G9SCcRnY/KyrKX1VP9d1nAZZEYm7EmDhof0YChgngcp7hgMPJKpfWkOC8PJ50sbA
GNsQabADuN7nx1FxsoH1CAXzXmMkBfUn+F7ziFPN2T1yTm/KLrESLgmKh5UAJe3i
rP7Z4mRt2SFFiw7A5IX5Lpe3njaTwu8S2LD7YxUqB708Ej8naFKbXXlDeUxVa1ef
hWAkAThX7JU/4AeyBX/BN4JT9yBkIZJgQZIs1a8gwJhqciJ4FJKpE7XmmQudT3or
qBA2F+xPi4H3f67W8pS+JLLxuLVepBnjaPysGzjivGqGMFm++deK7xZ8YUKF3VNQ
e/dv56RQWsK4rR6TPzPGSS1IbmFCoVPJKUonPfaYbZY=
`protect END_PROTECTED
