`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oHOn4wD9Ccob65FIrPz5YsBWr2JchhdqPbzy8xDEyh8q/tzP6rcJX7mAsBVchweZ
3m1eUNuz+lybxtb55bsEGqDPsrRwiY8iNF3y5aS7L/HpMMbN1sL/zQ/68c7iPRcr
C2gtgnEukpMnO6TIJjOYeuIqU1ou/iPWLRQGUzbTtQpcY4SADl0ROGF7I6azYJpx
XFpGoEF19fCJ+6i9UvFbZWcDJOj1glF06Q45jba7BUuph2Yin0GyoCjgc4/WQd5D
jGin94REgodYSf+6v3KFp7oaBtTciumBTb4MoWsWMbAmlLH4Q3G3AzUPVP5PQvDI
9AekmwObnLcFCijcORLD5DerHXT00tezy5U/wiywqaq2xNUPOCaKfwnM9Nl9pMC6
eiB/ecLhePgboNvmCjine/pnHfNJpBteG29Cq3ZsoAKgHwdDa0dsjDWoBLhfQn1u
t1FIcnu/sxyRoMCEwZPxrc8gCOV5J7HOIjNBz18XwjIOWImVEMNwQNAgEPvkm48Q
CHsaB7b80OfvkBi60q/GaTnVjSdcoO2B5/HhHIcjmRr1fjLdMQzm6iOXQYbHWNNv
vHLnuo4D9T+pCtv2n8i19SLoOAcYVjp4XKSHs3CEXBD5h6VGzswzcP39GC05uft6
FChOzq3S65/tmL/IVYUJnVEXCGKPqD4nVExlYDEoBiHLJ6TLECUaSgM8NS+V8yj9
l4soW+YxnpgYqxxB1g5HRqhqsV/bTVYUnvbNjqcKxy3Pnpk2GuvB2KKFKLFU+Y53
2VI4cUELEyDSS22wWHrzTmUfPZlNfwpmKhP+yCDjr2K3QAVABYO7TpHZmcvO0+/o
1CtnTzRzXde7vkmvDvLqp1X0fptEkIgNFGRwz8VLX1AxijMoomUUYtJNhe5R3Klo
d1f+dlwxG7ziLsabXtD10T3a8vCJVZBTKksKLqeCO3360d18t6nVH4bYfNuynxsJ
nf46bkWJg8orY76wId9odHgXO4nD5/oulGC2RLjtejxMMJNKBzHjoUxl0WtAzV5m
XiZcyX9OTivQSK1p/0AwAAhQKE0SMQGjznTkh+UNp6iDoamXy4nAE5Rhclds3pWV
BnB12+Q53lodj3A664aTorNj5sg5l7A5pgBvn4UFlvRT3qFFGR+vmfm3kBZyn4+2
nM16SHX9kNAHvuIb49ZKpHgXjm1nmHOaWkp6Z+uVQIgJFnPC3uTYnZBPCNQ7TIg3
L2IkW9760mh52Laz+LYBrE18qteiZ7pu57AzpqOxU3bIr92croJCIv5jN7Ms+KrY
FfGbVM9DEP2urR1vwz+n+TFYEoBpeuZGnYuLOclxSRema0BxrqSZ6HrM41Iqk3OD
5zga3xZeim3qC7GStieZFqaxiR+5z44pory5vLIzHWJ5wz5by2186izEZZWvSfmm
c2p+G9sEVE1kBYe/YLBKqy2sud5f4o6s1NemLmcfzduCV+MCCMojT1IOp1D0r2LO
aOt7g5UDp8TBOyWFfvUtkCAD24PZSiQpjbeWRZdamVDlmwycgleWmj4hMW8BSvVk
TxbmUaZOv+vDeCAcfkMJuuhWoW06NU4PRRlN2iig8TAbZ703pIyYHvVkVa4dl3Un
66OXNSj9oFpkWe8RhMVdbzzGbVeaP5v++P3VHKhFiGpTtsJGcsoI8lXsXtRRAIRu
wL1RePdGnRbLJecp6S5BEVqSfq/3vitNX8jzuhC4THcn122NdflYd8rmBW1Rdrfa
hodDslATPylpRRrfuC2IHRgIxLFvlu98GOsgAjrozV3ZguK0+askoO8bKEWDAzhP
WWEsMBeXfHHxLXEOkfzV1wChzhOOeKhH5S1R1cDRPFx8UyC2P/+9NRL9Y3J1MKb7
pPxOfNRLldfd9Up5jOpNfntYOH/V30gJc74Hd93hUNOfHcSQ2KnYyHS4E58h7Hrn
IrYUj8DnhkWBrHJgKNogPIHtNOH5UACgrf/UgjPNbJsN8F1FND4JNfJJIT0tr+PV
XSocUDlUC7AJUGXH/gLE8U/ClpQg5nAra/WUSwDvReidoyGxElGHNIKIgR4i1l4P
EPz/Vj/jCpK9PsOJ11BLkNISzOkA3N2bfVUnoWuMDukrwk/z0DqXZ5lhvxgxjST0
nHMFP1VacQMcfdlEYQSqDytCc2SUay3jPu+ks45FzILocYzTZAouo59YCkcl8Asi
hIgFtJkZQ5J2QU+FuGoSFUqEiXE1sPUh663ETyKMYGpjYGDdFWX1V8lD4lGNqNxz
LxNcFi3Iwb0bvPFGElucAYTDh/WvofeXb1+lugm5CcErHyZQxGgLBlgpWrk/8DAU
D+/qULo3xwOlpbobCuaZJZaAP83eRySmsYoxmB3nROiuQlhYa9gahL0dNCztzd8D
0vppvLShGJMZ9p4rRk1RIEWydM7uO0pt1DIHCJkAmEqkrz/2v32+s0rZpDjInVzC
sq9+kl6PRhQITYtlV9Z864QGDR/2WAW1bPheajison2hOOPKR8MJj/ecnKMMxjmQ
1MybQannFJtwarWtQbZpmUZh1Inwc8LHn1Ilih4K4aYUMPvNXLPhcx6Akmz7qGFe
yOHguxCS8pSjRNfXy4ZJMpfsecLF7crfeU35bjITsYfghXYln+Asawknv09K6Ppy
aUHitjoti1TcqcBusZ+w0hMdPon7vfmXHRLFW2zdWXSa94I/l24mBdHhJyvNBRqS
XxdgPxHyy+p/Hoi7MvceFMI2u0y2pTBIySLc1ro+OSL2OaLvpx+ccTVG0h2itk3Q
95nUXqia1/B25CezL2YyhHDf/3GR5He3Csl5X2QRHAsZNNDwqbX9G7tiau8PatU9
LxfZbd9FkiTjQK60HYOypXeIQoS70uoNoJssmTs/m7YTWdbXDPwb+nefVCbAJjBh
wXagPMubLeE1yZwN0g1e12O/JYZJwOroT4GGZLt8NvIq/if89T755d4tyBrQyoX2
hLx2a5IJZHfp712BidftzmNbqfIfxh7n4O4/a5Gr0YSjrHx/B20JGhWHXpBzLAs+
usS/YwcGPxKYPAFq1EiqHNpuiJP9cFVI5g3veM1fee3DXx/YqFUs57XmVhnIk+Nn
yx4fKTak6aZzi73/uJT0sLmSv1aLXu/xLWRm0pvAseksYXTzlSaOFopbVIikUFAZ
ARBc3awXYlG4D3y7hr15GbuipRiqYpJSwN+3wKAEXgz8LjOEY9S/QoJV/W8CKGbU
56Hb06m9zpcWgyKoi3K7UhJHuLFyMWeYLkPhpI5dPcVKJKT7HYj0dS8nJHmxPG9y
HAhov5qZwqRRICSulmUWrzpbSiqQF74ANd0DonLm9WKc+q7nBcMaVii5giV+wrgt
f9Z2YCBpr+xL1HaCswkqgz+QXM4Z8nOo2uNsDCFAaQ9OtuL8Ll0WE9gEhkFLII0S
m5UAMSd1lxqaTQIL67yRpqJFkOG8gLnfGrFxJSqyo5NU0vAx38CEycd4iBqjVxCw
6OAOkj7ZWfQ5ZbAK03Q1BfExEXqgGYDk2JN2xa//AOcCb9tqt1V4YilisCZaoGHs
vzqxshDL9SZRtOw1a9i6uikCQeQ9UhjdddmCFwOG7DngjaxXQzmxsa7FwDgorVbb
I2KGJL608rrEy7YimdnQ02NTijkkonKuE3Z2aEPYAEZS04ShrbXvL+clhVCe8uIV
Y7SJufwAcn90ENZviMYIF2VEpCvzLu1liZkMoNSyekpEHT+pUwKjC8KtxFw05zI4
YmHuLUX+G98TLimjw1hk+evzUAHCoTuT0t6jkZHBvEOX7LcuV8BY1YQloDVxIOvc
GKETQETXMc44eW37TUvV3vNHiZj66THK+Qszq4MM+/BVBYA9Yvrx/JiZ9e75gYoN
v0FFBE1u2yfsDfzWOtINnvdjEE5AZ9srhl+dr06b8lf/WrhRaIKDX/H26PfTqAFP
VjJzA8B+S4t6JM58W3C6b54EYcLUFt/WbWOFmI4unxg/2hl0RCDFikzY/Lc+QcyR
pROGs4FoKiOG3A80u5y0N80w4fxJcNzBDxLHl1DVis/Msa9VdYjyDfocEsuGVaCm
drs2oERZBCuOJV5YKrHf+o0p7zWr41YzQQjcKQPC+1m2BdXnOC+Ut6HL9vr5cj6T
U6Gbv4p0ebFxwpxsMaf5kJXonu7mJINXy/tIlNx7z+DOV46kndiSt8+bhttqjSt6
AybyVFBemT9AG9Ryn8Q7RX+mTvLPiTpEmPA0kALJBIdrOIt1atOEG0xlvewTwG2Q
K6d8A+zQhyUDoOrUjNPmDBLyYrUtLI1cPOGLymFzxIEg+oBSY7FzRPvd9U6cxCm0
E/gOs9ccHlATXykdiUrMZ4m23YOKKi6d3j/g0myASgTq9Z95UKlI1tdhl1GRKNon
TiRfNaeHGagRIIMw3kGy3+7mc4aNxal9C4kJTl+RwaYpP8xKGFQIpXATpYrRSlCr
KMsH1jmfqpNDP+zOsjRaYuqHRRxJpSgv/Z9MRoZz8k6dBaJ80RZyicA31DXX2KIM
7oDHwbUwTLMnsbtf1hTPHcwuJug6bigiVRCJBjKEptHyP8Lo/xrMeevyWF/g0sqI
DNbERQxNVhyWILZ4MdOx12SE+RrVxMN+/rEShf/+elH2OQswkaKTRauZ7tvxVX9q
KognRLelWLpi52Ug7Z2YLRJGKTTAYRDeabjiJENcUjAhe/n8YIQy5P3uenhrYwq3
8r1t1JbLLQQrd1123sa4b+qc9otz33buVneRtdHVK+yX8HoHfCduVTJMtryP8U6u
eJ1XRBa7E8mHrRMDd9xKyDT+voAxFmN2mHk1j99z89Gh3vwKH5Aa41+1x2K3ofc9
WNBc4DRkEKX66CCfTZsyF3Bbnl1zCHkbb/3F+xkEbA45BTKYYd/0YSu1Hc7gKRm9
QFWM72g5E9xxSiAA3axYUf3UWFW/BFvuzENgCfdpbu0KLpxTrIpjbhhN6nssSYHh
4JVx70jmY2ATRh2dR961sMpKD/q+OT1mdetUu4hf1ieAB29FZiPhIY6ex7EbEg8a
h/qzpTbdudYbE6dMyuZOzNg4q2r7XkmtF6/DMqONwkmqIgBMU6EXtjl/ZrxKiKUj
jfhBc0otdl5h7gJs/d2ZVdia35GC97owspm0D/F12REkf5YZXHcp8YANEbYZGkA4
VeDvmnVYs/TG71g9tjaGceqWtzLC9MqrOmnxf7XC+8LzCcoq5v3M6uYR0LpEP9e/
x/hGsWoDFpnWUleojuWjVjGvmLxa3w/OvOYrF9rhSxTzdF3AstpZ1yMRDf2Gj4Xt
LvDTzpMpn2I8ftOXl5GoH6c5HccJn6Q4siBLUqY+TSIeEPktQJG+hKYhdQ9x+XJi
sRCn18SW/iOrd+3ohX0NsNnuSZ1Kj4W8h0wp6AMeWHvBBSWKL66iywHRUwVDSgba
jOmQef+knPBWs+HsX0BfNa0Np2NlvU2AHPn6HAy3okl1WKBN5y3sSKt0mv+AkWPE
bY5lVYSAtrd6g3dDw64hcOg4IqRCfnkozxx+9iDHO8qJ7ZvcHSpwQUFEg1yoq/mQ
KPiKNGmx0axqvvy92dRrlHnuRFuMxWxHViCe5GzTGzLJLjz88qveHfMKU8uhdUMH
jPt8aLBuNasEbTpiySo1zDwLeOGhrnsHNFlhp56EZG1Uc/3xqrrMjj//rCBPDYWr
TLFbVMEHsySq4MrYwJuuqiMPjdKVuvLSzdFu3qjFeta8dGlQNqZr23snif6YKDD9
g2JVtsd5/+mtVrqrMc6qgi0FfQDmnJYJKoJyvy8fDOHCyaiIEQpxt2z3xtjWsys1
7dIW3MA39W7pIjxRuwNiKlKVWzO3zTkHYxeRCcP3m9gzDOmGo/hRqvKjJxhyu6q+
KD0Nhb6JCo58xsep9B/Al+ACTIjQPwUfnFsP18pQCj4gjj38Y53a5D14o89x3MXP
PowbNqsjnJ2HuHL3/qvWNppKrALeWxdm8/uxET2aZhdLw4Gu8xBu0YKm5OnAx0tG
SLycmwuXts8cEoxt8aNi+oQWqKCByIwhe/HxaOlv9Bfnzmq7MP0J5e5u0hVm72M5
JOGCL3VdB0kSck3DwAxfe2syHDRZiHb9SDzE3OzNHVRvjb2wcebWBdVhSjrW3atM
c2rAyjNCr4BPd2KAk11dMEN6XLPOGiDXe4JFThAkNsmqPsBwOyx5yFC2jQRhmZAd
KdZ7y5b7dHxdezz11RLVtx57KLISYSE7J7vy0MzreEvFW63yvx+/c/cHgnK3O7W4
8CqDPzzOWRFD4S01/Ep+fAXFpCE5mCg0Icfk/AWvbWG1IXcEZJ67sNZ/Ik3RpCkp
wiUts0uadUCUATyGJiouVzz1jdtS2WLFn8lm6EeKSsDwk6g+Z7Lkuj+KXzDHJyEW
qGSiIMwG03jXoXls9+BFT8yrMVhDfFzQzH07/vC3utb4RNUrsMvcv9llasUtB2M3
J1r5kadrZAxWT5njO3xNcDFcq62aIF2Kpm1Yw4fR38GldwfjmEbILQUwCgbT9gbJ
4dX2w/UiWHbbqQ/ypE8B+f5fhaWFSMR92hGbXzcbp8/HGHPdQToWFNiQrGdonpom
EdHsuCoudqcNuXedWwtwH4ZlOUjpAG8hUXaqOoGDLuBU6FBDakTOrwgGvh+KqWD8
D2pFRfDW3IC/ok3ZLXZuQxIcO/XtdjimSgkwxP1cWbHfSvKLVhSA2Spcxkbw+SdF
+awohVj+MjzFUQ+0N15xnHLLfEWClxUZ5BL06qbOC5EV8jsMq5u4pc/Wo4lrTbbU
+e8PJe84XB5NoB7Tod5agsUIIwzrYkBDQsniEtSoXzm8e508qJNnOVIHuKyl4j62
+ke7Sly9vS+0P/WFxVss7tbNFpC07hWF+x1olRB0zh3K4b8JV1VH+WyB3oXZa3Oj
rkZ9dd+QL270shm9GeEjtC6t0A3rN+kH/CZSu4LPr6UdqrPNPGMQ41cpw9zj/Cba
PRHui1ANUlvNuq5XP8MbdFF/ceXap4Hvls+6i9uzRMyTpnOOAefgD1ZZfvzY6PuE
9vzmkRCH3cV85CZzU3U0C2uQuT3z9837YJmowy8hI/yXu05o8PZqYqLSyHKRrmCC
QAb1Rs61IhHrGkAHFVX8f2TUJwUcbLSHbZnXAOp7PuPCjeGdllkxKlHrkHxlpM7G
UoBoM3MPwg8YAfPqtr4eOdZlXNGAjTh+5uu4HyAUJ0X4V0wA+zP1u7oUi5hAPZcq
EBlJxPCKBgwz0JnXf/TtnyIo55tVioBjvxq2tfUw8R1U+bMva2aJNVB7qrx2ehpU
4XDtv9MCMxW+L/QxYhQnAmda8WQ5GmVWV6D/FjH6BfuD3uGjmVhpG6vg2AGE3aRN
0l8xjV3/G5AhJlcht8QJ9Yi5RaHPBIbPRS7QzJZCuMPgxzC68jGvocI8MsK2Rykk
EV3gwcVTh46R6CtaQGJF+Q1EGW9fTqNVEdfNRab+tqTwwTL14ckkKFhjYKXJTttZ
x5UFIeLVaEg7i4BiW+J1aaHjuFiCurxZTZ0KXcjIToYAIQvr09BS4e+NkkOHKliL
B4cni64xyZiFslREJRZ0YDPhs8wdeR0gkEwrxzoRDShvScKyWc9Jn1MPUQp1a0tx
g1nAzoMmZaLA4DpkOaiCZo1Ry9aZIY9p/Yaz56/FHzOCxPwVaIC80uP/6Q/rXgYh
JlOuZenGZ9mGSdfWOmDv5UVJ9GIoeJk6gjWOgpJh6SB/3/vktTR1PSmDrW3uclVK
jvuAm4Qgd3Rnj6d0Hp8hYu93Ed9vlOFe3GUGOD8EVtSEc3UwAIyR1rQYHKA5Yowm
HS3OfkwdxOQ5NXFlpFeIzVKs5HHydpyskVd9Z6gXI/7G+RkAXvUNkBSGZrPaZi1I
750P34umnODH0wwZUxbbF4CqrQL8prfob1RgUhz3UdtoDJRMqtyhAxoTQYemztAN
VZEw8pMkqjSe8Vu/O/LtovUFFkm7AglavN1Fmtxe7GyC4P0P8+hZ3LVyv/2w3bDt
yVlq0tD9r1tyjSw8Dzipo1xPlsunWkc809+3fyEt383u1Q8TKeGfGNtqdOfN5TUk
qQq+E4QkdG2p1dZy/2mauMAhj/Vpys9KwcMDkgGBSnp5JWRLFOUuCDGtbDN9tPGE
dBIdM/xo8TqjGYFfURWm7+dmJRFEZJJIQdlS7xaOh5GA7QzIxfpbk6eqG9wixooP
S8G+4KzKgbm/VPhW8bmyfaeNBdT668Xh4xDvRQexGx3KjA9ckLu2jXiQ7nwFasHv
n1d4Mc1u/SQ8UujBLp4VbDkE7+Lxttg4rPDluCLQpotrmMb6iOJKxIv+BcqNMrBt
ATC9hAHtZKQpeuy+hVyeTCVt+7AFun/lNAfMywcVhhmrtVjlEepQl3hzdFkvioIT
qNZ6/jmD0lsK+Gj9WEQm6AFqozYaNG/1CY5gdI4ZUyKmqYGB4XqS6Ru1IZHeuRW7
bxF9F00/2YqycrklPCU45JQ9qHlIePi5gyU1G0L7t4yTudKDUDRHiTwRRlMvAI0A
1eED8p3+LZshDzxxcvRTcot46Zwk7wNNq1FfbIE3hEX5TH6RcFASuVguIq0YbSgw
l0wVYsX/qeMwi5Y+NawJu188cQe0c2z/A+R45yBo5rNsMkMkeLQEKkKLmr1ou4R4
rUD69LxGAcnk0N+4Fob+32YvVT6EwleQ2rOakQyjKO5MbAIYY9aq5Zn8aT1p90HH
B+xJUr+qNdMvT2X8UEER2lAXTX6wSFEyLkXKuM2QCxtiBQzmEq9mM/tuFwvbBxq9
xUBxnjf0DcMBLUHRWIj4vdM84erPQFu0m69Ikc/tP+DuXeSs9LgqsGX8D3xMw/HG
mp9DRKk2Xl3P88IBnnBDceThxV3w9C8SHTtaXHkrFjqbUZhxd8DaNhZJ7FquiBAQ
5M90vOXT94JhLlDgDYj20wcs+ypeyfMlmvXUsC1iNIX8Q1052R01dqK/6C+w3+s7
gKy8mOaOe4H++SB56PSd04P9iyOdFul/2/DaB3urOoVq5/SV5djEJv4VdYuqpjHN
611DeNRIKkg+7YhtKJDBWt9KVuRKIeoedX3s0/833Kz6HCbqc1LdqkavBqEfHVaZ
`protect END_PROTECTED
