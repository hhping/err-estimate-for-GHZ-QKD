`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mga2G1crXAdNjzfu8ys42PT5/uxE4eb7FvMWfwAhAuno0VkaALRw105VfxIV3qzX
qmM7/Yah2YuaETkKyIbTg7YQYJBuPCqbpTbXAe22yFj0Equ6tntCjlwqtxiXfd+t
j3Cyhv3Xe3JHCBkjZzIu5fv4/HCSvdI3yckyvHj+qf6Btsbi1ub+5sKnEgDP4Qdd
NGqlvrkMx2Yh0WymPQ4wfKsQbSNw/uCSA0mOBKkVaPg3dXO/jv4MriJbq0dYxugw
H8e/+l2EzM/KNRn2AlPfF11SQNsp3FaEJeQm+QCJMpbwAfzsYNp61IPGEbDSueLR
JwJYbn89nyWsYtzVRkzpy/z/jJAYu8QYLIUWq5IKkfbe0tPj9UfNm8AmL5IyFAFY
VljvlCyHYQmUuKQ+cpqTWDMojLzBv601NzQ3L9qzC/DrsDBahPi9GGwn7EDq/U0M
m9qqvsi34TjCDym8zVExzQJ5/BVqvTwrY4LQlb9QES19Nb+kbJoe5bTDsBeVkjky
rrOiDsv3qpZoLGETrk3UwbQmNPO6Vi7W80ZzBS1SqhfO0sNg5rUzfifqlc0EKEHA
H7E49MkUFylKXMogmQWD2WIUC/AxT48mMdjXkclPmnICIaWfYB70kWtjcckiBmNl
nspDNeig74Y1w7W16XlXvkcElIhp9h/u3VC5zxqBxQleDClnNju9CBAuGWAbT23i
p8jyPq5CW3Wg1r48of0/nUKqkv6e93y78RFpAgLwZbtqDxDyPSiIJ5fKeMCXaTmj
NvmwTscRajKz9pdoU8hwysDZLHKmbuPcrjVjvnMd0AU2UPgNaQKaO7KlFZi8Sxwt
WA8JBulpmqq2c/s9PbOJR78z4Q96/rTgVgplaCACGN/yX+nI7r1ZqA9+EUBA0iY2
muT+Q43niEcvUj8cOUrW08YwKIYm2tgvp/bMoXy0gzNkvlt8DJ2dFuixl42Itnng
p/T3Yr6sJE7hC3MSSC1s8hh4vGnjMqtfaxfhbsO0FEMGmBHQj7BzSBR6GkZqJqEk
tzanyPITCTxMBjUl5b2yTOwBFwPtBOWuL5aoB1svWn9xol37bQ4RYYAYaeF/y4jG
SQXHPr0j7MzFwtitWJQzdPEwEi4CUT4qh4ap9w4Ub8ENacYioDBJSqQqJBeqJNIb
McFsYuQG1YOrlc+MH8mxV/RO3A9fywLLZsXbr6N5yY8lghunae/sZq0AgoFBeUzw
jRBlhl6jdg8C4X2RUtsYDGDqK0VPeqmxnPFNRulLbUW/eKynY+0yQeFZzGWqN78Q
WnjgXOfnkbA6ON2kwdDyGkyGrGvIvZQOLgyF4zfprV4WPoZWwTUpMsp9zPOLQtQC
vp9wZYdAKo9G7F8bNZ+gqA6JgJcFS0x5JaoYAJbXB+Ia7E0FwyLteKAw5I26K8pI
HXL+U5d+CGJd8fxfSxayd0ZTihyxNM6vMMlWmUhFq1Y6TYdNSWNLAb/2mT47gyqH
mJIsnJFucUMJt/KKPPECk3swoJk5S5KEzxnukliN/EAvnBZ0uuezsubw7T5Qqn/O
cGQ2UWujtzk4kIdB7YQa/CJFx/WP2f3fzndczPSS289025i3QukJKjqGESJuYmqZ
2trJGS8ZgGd6AQX1v/WkigvAuc0ynOP8KLkoTsZ8k50VHtWZl7M56VsU5Dx5MwEB
jCrj2Oa0ewfFQNz/CpMVHIRlRT9rZf09XlC8xZVxiaoMX3nDznTZFcxAeDZxhEXk
c9NbxLOjwuflYTQKvCAz+8Or9OGogsK9FvkPSoZEPmVpk3XIjDqS0pzafbjYKzg0
zgomwa9NBsxQJ9m0lbgbMzFiNIfh4QGg97M4lq6mFpxZjNHYFN+ePG8dwKyoT5Or
EqKSakNOv8ULu5rhUTg8gIFqXRhPauY7gsOSl+cKFMpYfmmnCzX+kPhVFwpZ7u11
8kzH/EjzO/mAnzti/n7PCFE77c/VuBAcUImgVv5bUNpIRaiG1UDUZ2TNdBs9rvpM
y8cHTPjWrulokQIy9Oe34euPpvpwIjesJYy5602/w3PdLIHhTjDkY//DXKPnDilT
KrR2w12r0jcJNFiakfUhdhrkFV+3zquKZVhLpUhSY3s9girHZdAcd0fuViEeXU86
lTMMHZ4pbro3bXSwpuM4SfAU/ZNS/IiA34bzGMiJq6ug9TCexIOC2SzBCdHncZYH
13+2mOOuk9OZFA/NN7RpKNJqd+sZyM1VySwNcq1eofqZIwJCao3t7cms1J6cZB9y
lYkoGYU/3nk+oiW/wJFfWW0lTQWpgV9wNxuehxz9eGpX3O2R+O/3owY0oBLTtwHi
jYHdzA3HvbrWXpdcLAZhP0wHHzM/GRJ5cd55xGdwX17Xz+10lr7NhTd8K42HQsTA
4MMtUNWZ/2AzSlHwkwEjldf5XNpWFY/9amsv1uHDBkrcg3xs36KbIgJ3eQzWL4eR
AjsyjDjiIw6zUuxCZt5DabDRo+l/X1h2kVB/IHpg8c6Ri/JUXxyp1OFqTu66JOUF
f7xd9YezJXqutB13BW06R8dbO6Cf/HV4h+G4TlO36dvmz94CB3vUKONYhfS+e3i4
80V8iiYAbUl6GnY0PAk3bnpDbdzCyc/nf884RX+JQGJcu9PmL/HTvkwvVgNIKYTv
dXU2r1+3Kj3Z1CrQmsDWkfD7ewerifLKSwA2LpiO3Pl0tHA8eyKjq3gWnsQtOksz
SncbWV3ZeeOKWnZ8wgked4RWDdW3T0ow7PuArIp3ec1ecf+7VTix1W6/h8/iPiJo
KfZhwJ20o0D0YPcG5rmC0EzxBp8fgQAuJ3eT6APLdEhzxkoo0gssXgDRMnTWGcB/
DwoKvhS8HOgnFynTPtyThK9iAChKPH+MpUC5MOawSTEqgchNU76hpex5jk+3iBAU
foEAKJDYrKswsGcL3+NIcKCfw/k7J0PhihKG4bIKPgkx9lriTsyTak7VjbhcMGqG
GvU5R3QLGBoLRNDhnZgS4mRbPJp9ThIN9qwP4qdrvzS3BjRlAKLTxKiyvjz+gcV0
3dIpRCI3siCpoYWBCmJV3Y6tZHhLv5vX7/4laBsJHNqOprCFFr4nnm9USfWl1Xib
bDoRx+6Dei1Qx1SMjLTRxr1Vl+M6kqL/9j8rfxKxX9IkJ7Z152QGJ+5cpsLpKs3k
afwKhs0iojgI7xI+W4lIlQcHBBH+RC4iMq3y2qG1GQx0QxO5UCf+TqDxmQVC/AXF
O7Oi2qT3yNPOgdReUVh6G2vGrCByl5OUVUYEzYBUXsvmZQBAjmP1Q7VGJQoxP0Mw
Eift8KnEbOGEYjqrQeEsJvYXkIsn2ih/akPSYNjoi+oO/WzOtMQlcsyt5zKoG91q
qV1lnatG5whiZVPPXiY3BcWJXfJ9kRPqWyUU2j4KHuGU+NzmTPcT6DQ4DaT2mEGr
El9838aX0yEwXUrT/U9Q6j6d3SVUxWJ/51uhKkJ2nzB8xYVgkMOVpxTArC6odFpW
l0KZFTg2XGZm8nlw/MLAGUdEOWojW1vejQg0NUPKvrfAj8XwcNqpotfQJjDVpS4t
QKfHVQaKySNNh48lKm2JJG2hFkkA1BgAwrDCN4mNd1SSpja1JhKwsKHxmGEP0rK1
04T6olj0nW6VoMgiwg+YcRjpu0qVp3VW8mHyZdRRq21jqqp8HpD/haljIh32+RcC
IkWDPFvxxLhuj6GHKtwcMRK2Am3av/3JVvMUi699zbqqiHpJspGK/9uV0AgRsSPG
/ajILTQ+CnnNudjw1ywhJ23iyUlT59ivld6OTlyqB5ABhq5lTzGGPlQ60PV4xpGC
cBbqTjhxHLJx/z9zS3bzCVquLO2CtRQyywkpwtyf6NuRZ9lHb+8URSXgOCM+MySK
Zdaujri1DrCx84DETZfTfoN/jriuT9obz5u/v1WzTJvyBz1ubqOrz+uEh9NClJpz
/NpDAB8JhvdiIhczxIagczkHoiijeNs2VSuFT51r35cJbf/seneVu6gk+eCxW2X0
phRdYeFO5X0WIPZPdLIQdHRok9ovn0VRqjH3KOPdDF7Fn1bV9NxofUp32iBm5m+d
QAj8pfuLFHOcYRaMAKxRTdnII9Sy+Ae5NCVDFvFakhxjBzXYDhh6J+DT45F+AQBK
kMphJtgT4pRcM+BPCrjjx2pXl7tGTVQAaLGCqTmZhKog4fFy4YKoOFxrWsbeFEaG
0JvI2VaujKKRd/9l9stk5S453wQ5Hws4H/XGjB3mtXMw5p6B1wvJchCbVaYSqEmv
GrxxvMbdGcGCx8jYcZ4OmPQieIgLhak/6CJp4nmFZwc/ALu+50sIEGkZi/T7D0au
ypxiFzdXVdDHkiGqLcoOj8uxSAgUKavK9uFr7E0S2LI=
`protect END_PROTECTED
