`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QMtZr4znlGWLlLFSDUaY5M/esPleL4XCwChKjm72nWmNJBiUmgUlO0edGn/iLsml
SRb4VyD1bACHtnXmSjgYtJ3R6o2xVHH9bjZunKl9oAuaepD9AZnoAsHQYnvG3nfN
+o43WYsOAi00GFVWyIqTDosys9+x5qpRlwY6KWcrY/InMmfDJ1eI3KlEPI8FXA2Y
VKWbVhdjoEB/n3ivhfmVQ6KChvUg8AH2Wvm2/O5F6VU9iqMuReXmnyO8HplymYQe
ZiXYrP0ihGqyJNSMR7Y9SBIONX1Qr8tOFVp6R+kNFVsdtrP+C/prLhOfg7BXxXqg
7IxPQa04rnoeOINk0ipaQB7LfRp9eP05Yzqp7IiRnL3E/brccjv2+IFbP8X+e//c
9S1gas0yJVgvPs+eyse3iLzvKFGmqurFsscISk00WRRuFliwZbqYBD7HNhJXJwuH
qsGlRy6dIWKxkkBgUBqcQgNnpozm/fTwkQN2kIlG+08Vz31Bxvf2KcTKUQgocMum
29KDlzcevyPz4LErBqD8WiGsDNYdruk1knt2wXeZz9TuJHVA9Kzz9kkfsf/Vvsji
G9euLieqXhBK9dhhfGRCtv/EakBFWPZT1nZzPSBfUI7+DP06n3DA+yNbOV4jwJX3
dtmF8NghqYf52nBHJJijQCTjNau48zSRWA5GI/lxFYiQdVsFzEetuopHyLJZlKEK
fSnMYZbuPHev8xJN0kKwNobo58BAJ/MhiiR5/rW39LHySMoUfD9SqYopuQKD3IG7
MADmOzEDsAWzeYEo8noiqlCmBrrGYIWVVEofOyxD2kf4YR382ensvm2P2HAhmfQp
NRUYQl1TCm0dfSK+HSWMYcUtU0NdUVAF5ELwxc9XzHvHCZMq7hJ8SFVh8hy9itco
gFLhIKOeJxSZBQ+zqC11cehv1Zwli44VTJB/fRwTNszxzAgFDJJ8geqljoTJNpp4
G5TOSfgrtienQbnreH11UUj+zSibl0eKxLYngYQ/cLjGYnJa/MjaykKF8rxXqoU+
sIJ6a8YrODb6ilBEy9begAtwCEDJsn9UYBYDnqQETuGSctZ+Ktj322wVnJa+SGBg
4+vFzVf1Bg2feKAZLQSXoFzuYvCPytI9JKPhTPxNQqE2NImBwNMTHQ1+MxI+jCzP
G0xBfOBhZ64w9FNZlDd+9g==
`protect END_PROTECTED
