`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oe0GM0fH0S3AaU42fJCO0vDGBogF3Oa0wXGja1BpQoDo+qcsqmyfKfl850dgTVMq
YIYouMAM+faSOcGDGEfncVL1AdaCmIs3JmzZl8Ku7iI7PnHgPCrFHiE7S2i7LHfW
LdMbkjTAo5EsSoGvdhnKjYKLY9AJHywP1rUkBVF+HIqwRLeeXXvweqajKrCoOnx4
8Vov1fM6q5xDps4bs65lC1HkF9rSTbyut0udJ8ccAjYZUCPSHWV8tmqRSWfFv3aZ
pB4GnQh1DPKN370YuXRD3F0yMkKqMeF4EnF9JlQB/h2HX5NkqQASgcZh6909KlyR
J4WapEGZ/2hnwraHHK27yGhe0pVpAUjSqpbQLMrphONJW9g/pJpJplzXFPCZ3Xbd
Vv3sD0BQDzy+iPTgeUUBaVd8MbAIASN33VilfY9EN54dgBUqdz4tk98oLdb0bzMd
jYxc9AXhB5wBmUIkKF1VslQS1WEqfLI7jRf+4OWEnM5p5/e6vI3aLRw1Gu53Nm3e
GZEJE90f/yAYenMreLPgSDiNYS2KgheVXvYzSS1JIFU9p+Mt8fZ+ZNKcmgM0N7GB
WSRHxEet3e5FmQgMCD2C5Uhm6ebM+tO9ondIeFQ1yMm+xr1m2gFZjPvwl9jVh1Qy
mqr/adKjQ7pO5b6EUAlmIrPyB2dkR2ao4JFognszp6seVXjeejCs2bjoGdYRA0tg
HMU3ZP0xX8/xA7L76/9N2YPHllR2Ay3o26fe/LOu83kmqVuJ4/f9uNqlzwAQUPsA
2aup1h7B4S59bDyrAhxVM5H0pgcJKxUd2aUAFiu5VfSjniQEcx1OUuDCZ1SAIEJd
VHtfpvmVqOhEon/A0AfiizOB3en1YQXfMAEyTc5bszg=
`protect END_PROTECTED
