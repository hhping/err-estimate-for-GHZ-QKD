`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HbY6eoyopcc0IF2f1T0s7bEa8pT2AQkjTL0iRm7CZIg+V0k7a1C9Kw4QAW1ISnTn
qRReB/XKvHmytrTaw+6A9/kkJvDAwe4QPyksvgPeTOs1i5iET7bNCzM84nBrfKkM
JDQqlEY8hp4lnZP1MYSXwWK00W64h8s+Zk6E0kgHnF29sxyqakn5WUff0YkWBlcT
w6xoNyAwHGVms+5qw0AugY9g2ipVXbN3OlSNOQ5o9lbvMJs13YEpBhW4Yq9igB4o
0Qig2kb8kJwXDbKWNY7zdLPqmMTaW/okgq65Hqk2Q0jVAeISXfawV9XR/4QEEQVd
qwYRqHes1CyZXWoFoRRTUQ4f/j3qdyKbo/R6aYL5a7meq1WWY7ExJtv9Ri10f+Bz
2LfXpb56o7lTf/spu44QazpnwHE6WK+Md6jfyvZkXR7ZpZRC73b6LhM7uDbIsATc
2OLt80oZNFK7cQDF8wPCBsM9pfYfutgHWc3fsEmwnfXEJ4UMQa4P74wiYDfrqOtx
MtJq51/bAutyobEIE4k7swm9oIl3Mt5UoHZmQQT4WOgt+AThjhlhk45CeZUmyK29
2MVxZvgMxX3msX0JsZM83gDWUD7RqH3qrvrYlvIrligJb9jWB7NdYW09dnWwvEXW
Uv603e7sj1lpL1EsN24X3N7AEhpfPzx33ORIarS48B0E5vnDNrZB2QHof9lWZKIY
58xvrW06GMVDqZLA8Nxp3JL4dViagvLyR2lG5dEYRqnQwieLGkTe5V0aFUZWQ7g1
Zt6wtgeeyl7eNA3LiqrYfWlX3swY9BP1QYpHaHp2uNP0rDgYelxK3QTJLO3cb85w
15EPMEBOPyp/ZnTwK2SNps9kRWDA2rZxGW+hL1VyYWyMdyXCK/xFFaUFl62IYcJi
ZzrhLq+cVlk8aCT/smVJIB+DUjy8fJiXw11TtMHI6y9ohvAErU+oOZdnMBLXeo4o
MROJs2KsjHQeqwVY5FeMZtKPlkAojWSnvjFW9KFA3qGyBiNw2eLrOJVBBpZI/8VW
7zMMlZaIziOUZdejD5g2NrXIDBiRXm8G95GjSdDE8IUL0MKrWZVgragLYs0eby04
4m7t8iSyFuNwAQHciNWyVf5ekJcPpXsJJ7VerXAm5yQf6Tr8FuE44hJo3gsrwzIm
h//Zcp7TUClbYd4InXCWph0/X2NpJ1XPSDArnVyOPLV5LCRtGC6Kv0Pb8geyBM9p
re1seYiU2bOJJTwR/d3va/KnsxMl1kmOGXSEagdUgEuL/sNzxK7IGKKeJqRrz+wH
U7Uwc9RZJRzg8zs5ajj60U6J2VV2Hxwp8BzedxItz6Y5HRTQEsj9vGwQFzqwvs46
fylXrKfV97MEW4KLy30LdK3xyXpazHNUTVxcWfZa28Zvg+a15CIHLo2i834oYruD
RUrqOOe0YomrF6tp/iUnZgnRrRx6qMhqEn6ug0KjuKL+DgL9YZ1ezijpEl0pm8eA
wWbqp7KklFe9+fY+SePlbeCKTGcbuxvUKgCwWWp+B/h5eabuBDwcFP8bCoWRHyzg
G/vtRb6XbefMhZzw2SwinUKCA7XQ3P8ACva0xN3d0kWMGd4gI83qFMEbL6T6TjAK
MyyumyTvnups94k/IpGCShhsXp7H4E2ODKMes1rdJF4FhhyXyo60wkx7KEiflnAm
UdtSSCCzOOCUPS6aFv5b8NtFWKVD9nEiqz7GxCitnD6g+biNphyeQG7ugnNyO4Xr
cetP71Hz1XtXubuOCizlbaBdMNDxCS8a0Blbv3mgaR64YezXIkXqNEmDFMINpxKN
eBEX7jccQ42RPfF0C4skgpp4SlLn49678o+jJQLkYEp1G2CnEfuyiRTa/kwTvli0
lsVl9IFfNUBTJYLbZlNfKfhKoGRxPUGd3XXzYIwqHjtd/4Wwxpg2EkNreYw04zaP
QK0fgB5ImUTxJC4ucgvGM/tzM/aftcY8eJUW4QiWzozqeRYCaGw3wOX34pU3Yq+N
/5AadG6SifCvANe3G5lqzVHjtTLA/LhOGaUUN/y6p+a8rLbqCeKlN9hZCclb6Ltu
QRuNx9G5/acel/2wT5m+7GNuFL0ksM6FB8TQXpYWD1EFoU5hzN6no7arMIOwLSft
u+w3jRb8wpHQpt3SRq5fEpK0WrPo71HQ+oHf/clea7mT7DfUZE+pICF3TG5xmQ+4
Gd4q35XE1knqtkDQ57V72XC1KvWg5W1sHGUGc3Kl11DiG36/KH2QVi9qymZxcmtV
B/dWQjgpVPZSBhhBzYm/7+xOQtpJouAod/eo7ROjHbFi7p0jgA+mxLGXuiHNqfZj
R3zhiXbrYokUiaemq922Vmr500FXA7O74+z8bNWK2CMGKLiUPg9X28Zna0FGSVdU
61HN2WHNhN5seG2jTOYYxOgWEbPHJ2J1ZHCynLLCiPKkcf2v/uJ/bjGDdU5+VtGn
qeM078csb0iLAw2xtH/S/l0nIsvBwgDl5zYnDVVIpYx5aDGChpc8tZFxm/5/TeVW
0URu9Z88oiTfROVMw38l9xPmgTg1gGH+XwWiOm8+3wtwolKygV0t0dd1Z7KidFfB
3uZCej+3pLF2fk0Bb7KSyjDYRXn76n4hWOfB6nC3ZPLFcz9o2a7UKjsXK25gYSxS
BSxM7iMHT0Eh2CLNiiHYnQAOWHewNLPMgcgwVaRNKsrWqWKyl5M4QtakMKTL29sp
BQJTBDdMV801hCzstTEHE6mEDGM7rkEh4uMkiPJJpm/k8qMFmK+V1ClKHSc1EEIq
YodHLxGuMWeBnQteEoHW7TkJItWk++hTTVRuw8LsaIilj8UpgfTPXSmAcsvspZnD
1qaKCxJh4pjjdBvkh/7dxLA07oDeAaPBFRFyesgFjYY=
`protect END_PROTECTED
