`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SJM55Yn1QntKrb6ADwm/JbDlWZNvbjOwoJq03AjOt0Y9T70+czguRliL+pRjMGy9
S50gctrbkCnk+NfOFCRD+aOc0Ffi0PRT0GMaUlUkKaZHL4oWBWWESrWyz4M5GNaD
js2FlA03+aCKCKUbyfG3z7n+wVIPtvlSMDG07PjU0FHpxgqIOSVCAJLq7wQxa33W
gMh6rzuavHc4NA+cYYYttf0WG2apTODdRiidJj9pjUiD/ejIX5bobKDXhR50DJU6
sEKOtr9Af1x3x12STuZEC2kMR0D7laxRWEhOR+qhfsBFdW7Rnoc435z/2RTvFwbO
1ukzRA2i7SeLZehLESN1IVwqaB2XQIRpjCxhzRZvEwYrt5E/8eFvqdU9YmXzepD6
Qw3F8fPQH9K6Vb75wtdIEYgppjxpFuK62Lk2c2BHTzY73X3lr+GWgyHv4bDS74GL
dvSn9Oo2nhGvP28Z/BMESV04yUm0SBmIBteKJ4X6FRMMrSgtWbQRhXWt1BmNByxj
H3MVG5BgkIe0Rrj1n+sNtRnXAaPMVvQv1TVdVNqqsKgteX+aDhu1NDU1JxCnvN6f
zfk+c1zMAc4tg6qNjcFjrArj9eOP2QSH9mi/aLUg4CEgGsErR2jKk5Fg6mlVc/xZ
fR0BDJO45bZixtWq1nrrH3sl5MjvCRwTKZa7rLZiLaUabYEWHrqqipvt4fPkbWoY
VedCJcpPVn0chs7BcSJEHVJkTdiJpFVkeWshVB5jF5ROcsCYUJ7qKR2dW2WuNsxH
KyUF+SDjn0zSed8+mLMBKGETB+lQl2emhEzdq3QF5TzYODP31vVFaTSvQZNdQLp8
7kJqOOo0pnZm/Ie44wWHGxN/0dPW0kuCq3lcr83pQYlGy+RSuD14HdBdDXSSVvYj
jXUL4R09PJ8ft81vAakNFH0v862rMv1d7VXNmu9FtfnEDxZrvGFyLogaj2kCaVn2
CoXaLpjhD4A8V7OJKHBdk9OH/YWQPArlbthvXY8gSqbvBx/RrGdAz5V6+KF0rkap
4yoQL29WFpIQynYKvmoUej3i3FfFS7vHqC0YO+V6R85LuAru5vYEpBoFdlkCZ2sy
dUKj8j8PMHKHasNEaFvlO1HX+VszI9EeosnwCRdO5j/vrZPQRe7LmZ5zB2GFgmc1
O6VsEde8W0hTaQHxir7wL3JlEHyq1lZyDcPjuEfLSDWvGZvyVc6idq+KnxqL91nw
7OYtzLJlhE62qHM6bLY08eKiAvF5BziQ4fjkG+yW8bx9vjopdpd6egfSFVb65k8j
cVoBUNqXg/kITELivtS5jydGOoyuRUCJ0LajrRbT+05USReLXjt5Bz3fd7IRjHWA
dg/Ux4crNcCsE343Iu2t+o5ie6lUD82mXiQtKnbvdthUHpnSCezvFBLX6IK7wpx4
lTXpDzjD1dweSAWTMn1Ras+yYw1TZ+1EhbuAA1zNRWTDrYIMBcgnsq18sNf3GqvU
KvPUsNjfDDtfoEReYdE2dQ==
`protect END_PROTECTED
