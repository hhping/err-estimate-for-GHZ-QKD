`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TXSy1sLHNAS1N8th5YwX7265cfkhM+myOlHbXiV+gJSN78PX2lw6UsSSqTaN4kgw
GfQGDhSLMxBi5DhFvS2NWXO+xjj22esXHZ/tGOZwBFNykGzdRCW+ErHaVeVpp8wX
t5HO5GiwRTeBl1sUfvH+YrSoSWbGtAd02mjAd43ECC1CXvLS02QvEymEVvc/VEtK
brM4lCddVjlauVPGUOSsNeOOJvr3qjrXW7U8vHPzdEF4K98yb711hMnoCW4i1NX9
vaOmQ8Km399vp2xmnQOb3SwPx0uduY2x/piOncVRGPFqPylMPNVRuvz835Jktemi
6FkW5kZzqUUc2MBr3hW1SwzOTVTTTFIXSKuizx2Gdk/ZH1WbiLSeEi6KgshCKQmF
GdyqXE/NsZ1R8pPSaZ0b3PzzK9O2rG21pUSxJgkMtBDnRle9K/VCOdThFeDlmV2q
xbxz3lFT8KR5A4+AMcTWDIXCmvAZdvAM5TcDq0hidVUdNwYMbgzqd4CxV+tjOhhu
Ruf/blS9+ZplLFfxa4rQ62FCVjwAL7BlbOZgpo/lM8G/jru6S4xo4x//5DyTsNSg
UKZuqlnBv7xiygTJZnGQx5eOoGcKoA/OeYDoGdDAj7VwnaQz5ztYsbw1SupH2sMk
+iyM3LYPBqbJexMv4qP8HlH//5eHNfa1/TzuoQhdAKbHAnfAaMD83llQB4bsdGVf
MTT2oThViISDugPKg6YqR5/ubbTTxoB0Hn/GMQcWoF+HdztD33vgWrLrJNrDwU2R
I9Z069Z3IjyaIW/OT3Bm2DvdcgnuOJt7Zhu2B+ex8C2qYkCF2kq6iTjTKZtCOdjK
3pr3WcqhdENkztTdQNhMLSPhu5T2LS1g/eWFFThGtJ2Gavi6tguQ8Z0K/oIH+vYI
9FYfPe5/knE0n9MayI7KTKkdCFCYkWPRjZSRqpmF+fxFq0ZiPcKqx3IQ8CgqwXak
G870hnTF5hEUAZNfvjLsmv4bWTOSgWsqxGrL32XKeCboUasCrErJuuAeIXf6WGrI
Wrehpno7fym3pZqqkZNAEBU0Mr7guM8sGM8fX0TryvrXNF8b0Kpar/l0fxUOPKnw
UZSTmR4wuxhjaPKarl82UU2Md3ZYktMr21i01X5ySLdzobN+6+RRpc9NBEueScaV
YiG90PMZjP1XUdVzCx2VXxd1zwKESN4ddYEyaT7lMSh38HEyHH0yRKMPlbeJuY6e
fM8waGbZ2wivzD07Iw3AN9kzIwLmK9DV4gQZG3pbPgSm6nsFO8FuU0TnGvEbrSgt
kQTDsyL4ynA11k4ueF06eCR8VDe1AFwThJ2yJ+MhlVDjDwI8033KWgfybylwvMwa
4xVKfFQCD6Uz7XsWz18CvI/s4LbL9Q8LKPu70Zf5Ouv9eD24ZUxh33x6P+M1T8mL
1gn0VSVX1pQJ/pgofZKUqNQ4oJTkTxQ4YSMvqmmSFrxjZN/VQreumxMvEIUZUtaP
cuFn5+c0gGcyESwjDpHpvkaohjzcHaJirebOjYUH5flG3nLXiIU08Y8M+qmENDTK
PLRj+VreIPqoZX92ppkols0C6IGgqYK/S1bFXozH0JyzDlLqWdmTpqCzZK9itPo+
`protect END_PROTECTED
