`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BBLxwJ5/TpyzbJvhCTVmWTw0NQxPFVMcPEaLVuo/D+3sRJmh8ULvaXWGFzSacuu6
E9A4qVB3zqqkATnFwhO56nPqWil9hk/ATo890D6PfIGlpdeMLp2WIoPfS7mtUA+u
qe23s4JL9l5VbIK0fCZqnz1zbHGcsFNbb2c3W9l7twg2iYff4tR7/lbAZkY1EaC3
6gLODLzBZRNQz0uMlOpQ+Qn2hMMUxcbag4K3ZuK0FsxKEc85jctlyToNK9sYtyjk
IX0m7CLilZYi5bz+0FytPrWod+BiU0lUr6IoGYPh7yOKG8OH2rWBGXURe491zi2H
0CiPEniRQGrC2YxY5Kp1ux33AT5+6LvChjhMctfP4tZNaUrexO3339FcUkF34za2
rgVPxg4o4g8gafTcOeX4QA==
`protect END_PROTECTED
