`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0wmCMW3zitSPW+W7Tjfle+SQORaMvGgadwu/+sPzPZGXDwA9P+8ZD23Y4LBrQO7X
5fzYjlrLnKoWm4PJPXs4wf31LnnsooBZACiJj1SzAaNPdnok7DCx95YDnA4YlKpE
5j4TFdJe19IkYoyU7bEOlqpK1huSF/3cg/vnvE0k9nNkM5sxD2xuuVPiWXRuI3NR
QrTG1vToWA9wpWWL/X+zpopthllkjnT4jDd7v7THCAYnW8CqJp0oSbWrl4xGyQpY
dbYln9SWHcLRQc0kgCC62B4/pPj46JeTmz5y1th45QUKolQuacB30KcsBQ7vWOlK
GcHjTbAHHNUvQiQ+4AlFcdXZZGwQ4CRt5iiil1GnBV7AdPQqd7jsqEEhUMXA8Mce
5YDhC73bcW5pS3cgxRYMs0g+89uTA4/Hba54sdpQo48WUAD645dNuKiWbV39H4wr
ujOPf33f34i/acFb7TjjJOpBP/umu+s4sIumuphxFPr3odgxcg+7n85fpIuPXXsg
m9jvRQPWkGaxEVu7wMCGL+IAeOjNXgd+iCGSOqiCLG4a14kdNEkxul1qKBw47WKy
OJvXYpPit7eqXzEmvk+2LALP+AFdEPeb5pzFd58EzE6LLFcFXuTuQFVMzsNCGf4M
J1wTWVYTloDL6G8SbNodFnVf6feXXwJPIGUmTET9rSgeJ7cvLWqUdKfbImr99zw4
YEJ3GvPUbe3mL3mxEqGChNllZMT+uCI3J4nDcoc6BsL6m+DG2BCY76pl20uGrfZa
q7KvkV9AsWROT3ZJuScfwC9f9DJ+3H5xh5BXBMrVIFa1h7M+zOPrgaYtxcoilCZ0
RAPhqgxnp4dUOqnAwP20H94Db5FcgfwkXRqaW7zD3qSDjfNTjZbsbQQMFkV7tujH
Fg1ZbmkbKiK1A+0HKGeRvokVliuOVrAFDNf13Eu7+zl3GQFnzV72VvqiOnuoB/jS
otIGRwwuC9IkuEHYKT2s8Q==
`protect END_PROTECTED
