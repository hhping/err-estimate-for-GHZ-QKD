`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vSFtpHQSlDK2jTnkH00pAQWVq3QtyIxDSHLPsFiBobxXzJZvWBbb4olNgg8LC0z6
ZYyy143i6QgseR7pDDPhGsZIP+a5Xm2dRZzaqJ/2Q8audX1k3d71oc1BgeKA3S8b
i8jezlpUx5R4eJxLNWHs59AuUCqprBGLl8GpLNyruERnXUY62pfAJ6vko3FDWqIU
sMCEouXmf8lEzoTfkx45DUjP844bsZ5yXkMx/d2xZq2lvILTdElopFtX17Bo3SaC
X5ut1sb2Ju6bEXKKYVmJzlyLZICRAPw7YXI5CQeOD7dgbKIggv2a4OXps/zmpL3o
PaC3iRPKJLBmGkzZvUgcqxv9XGOK35HyxMUJJ0HrDhlrgvqf2PjMD2b6CdgHEP0U
fX5In4IZAvATQ5pPyePdwrkvugzRDASzz0/lj7FPHt6Hm2XJoZWllAL5uqzixHjs
W15seeoEWHRN4hmeV2L4+8keGFZ9Fsc7IMCrovX0dtH9BSwDxQ3XRgUrdXbEhgOi
Yb6utD8UfwZCdoDZ8PQS6hjATJQxxAayRkP4EvnJTBo=
`protect END_PROTECTED
