`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UbD87sRh/rCBjQ/CAMzOxcYNyc9kZ3lkJWNoZNrU6iBB+iKLhYU0045/2H3VFAdP
xJw3v+DNVtHuc0/b7/Z3UfdKRUkrieFCfnsiaKKf6bgKcDIGuGbNqhJVNrx1xVXQ
b+iWp/MUaRgk569vOGVOmcm9MO/OQb6V2IEzbHqwCg6KcZu12ETUPeUOCy2AomSE
pJPfNq1MwnXAM6L/HuuIMQUOGDUqDaADc8IOpWhnY/Gdns+JDN4vVxfDDChXAq2b
LVPW5t9Edf6u7mWYs6VrJcHNAdaZ39RjMP7i+74Hw5bZ+gnfy3XSVIlS5oLyUUlY
5zMBB0uHsak1iIHCtQgulgNZyiWwx3VN8CWG3SmdloucpCxn5sQKzvDHeAvz0mYf
4FBbkXh6/lMvusWHthxw5PReWl17VC2prGbFvxe3rQqhgMqGHJJsDUpvtZCHzrYO
WL5Ap2Z8a5unH+AC9oiDBK9ybJzdHs9fA4jYD9sda/SuRMYlutluHgXJ9tlb4JCR
VI1TOMWdUw5QlUTGK4oXYT7zQxs69D68JIplJ4oY20WCCoR4rHnWAWYakt6hZfA0
HMOadXrvBqQTLA/rV4bcE1QyWoycBC4kKGpFUXNiM1vqiLtvDl2iIgcoYvJvSJ0V
n4xwzaiJi+VtSftFSaKgCque79aVLJDbIJ4DXja60lN3v2Z7+6hAfUcDm/WujHhT
YR2Gj4b0T22N6uydLyWiTvd3aW865lOWQGPFjgVjJSgPI6G0bvVQWiG13podMELB
g40vhud9HL3KNME8jdFMFb1CNxJYse4G/3bVrku/sYED0TSBdfuv87H6WN/AmaC5
g9qeZyk4lrFiErb4NyFeX8nJfrHJ32M5pGktVedmFFAsSrFv9P9v7o811Dxk62Nl
SuvGst6/Z+s/iyDJJG4PQBGf3QF99gvRpnqt9Lf56BiM1dp8c8GLDR8THdqqSYU+
pr8omPLjE83WaNkFkqjXalU96Nuoi5lauXpVAK+tVL0pE99VitG8xF6kuLXLYXg1
sFn1Z4oS46usOixcyvHmPwR7TXxOYBXc3NfsgGCVEM5BRcwm+VL2sh0C/IXYZdIX
lA4PGXQFInrnpC2kOsUEs6PLBTAKhIXDVLPJfki+Rmg6Bj2sXcfMzbmxRP5DDd0a
zC7VyventfLvEuV8gLkh/cFwQRImYj1OYSQS/PxLljqOjyBCkXStofvmT7T/By9E
VykQnhVZ7djO/ClTNUuDK9YvPd1ZHeVS/gD8bmeCgwCFPm0pjl340Ct2F09OLH/o
Y44+qxSmdQT6hivg1/VKgUcoWTmCUGtk48Opo4zurtjBBjEM/7tZ5UrC6umgIMkO
FwYhfcForL3j6bczybUqudgKepBsOWnFExZNBxKTBybTExapXqjgffO5SJ9/C10g
gDXp58EPsNXsJIMlssDjltspVr32iSKVQOEvVy1rzsq5V3fuwWMDWvc0iL9as5dv
L89vBt75H+PePa2Zm6mBR+VhsaaV6o1qQXCsTLHVjorb2qTpo6AugEjvGcmcFkpo
ouXfsDhYgBcJuhcJn+2Eqq8fvv93GrR5DSR2QKxhFvmx2HRSYS9wAI1ZYFIuUqxK
2v/T1v/UWp3UGm5o62bVTTYxZVSy3pNY1DjUT/N4jRWOGLe5VHew3bW0oMksuVpr
fEWnteZBvKO08gKeyjmLtPI3AqBtjYDvgp2qWeOw/zatpdQkTfDcrqzsIbZ/mJQr
9KLad0SkOACbGUWS8ZvChQvcP6kIPlbC/auEGPETUfP+dOKmE3NF5kEbPRliWC66
e5BmKnyjQiIFbD799EEm/llehddAowwaglyys+3eapxWFprO2PIhIP/s608/K/3M
cC6C9MSzGV3BX+6rwTv4dP7Zaevn/DF1EuODJEM5uFgCdSBqjMneNrIqoka+IMwC
Z6hxae0ZXTnsyIJbeMVPl+YLMX7QPob2UJpL1EMaCA8S6uKm6g8VW1LaDJ4hLguN
F+lpH8CPawQbB2a87NDY0ForVE7tlRLnVXJOmOEBBPWkvS84ou4Mt925Ld0wlxdz
x3PUfsgB+8Rx0FBFyoMerFjSuc+IEL1jMC8wlU+SBm6t16a+q8FlEFQCVyPmhXqA
korCA77QlWhqg3KK513aurlsnUidpKox7W2kKfQt23aZmjq7B1mMvSVhlVdgJElX
+ByIE/ZaavMXC71vSdMlxdCEQLRpf7nR8qd4gdAe1TaZM2QOpjtmMmkTLbdVppqh
7sU1sB380s+81h9h/T1F41U/8HMt7p+bDFfkNfKDsuC9VgolR83VS/Hnvai2ljcX
8fFHl2fy4I4MGs2Zml7jlPVZlskJ1E8ZerDglHo3f9XR00QtZJ1FrAHEdXfyqoyM
mgMlufJFigvKian3NatY20HFORDoGUO6tdKIwOe7Mpra6OyoDQoQGpY1uCX3xC8w
6wwGdFvWEDuV2P8AsQ5aw53vZE1EBC51X9zjhcygm4uTBYQyDnR0Y3ILijsi2StD
ekDPb5k0u/wbnfEU7g5FbeRynB24fNaWbryQYxH8JZp9LnVwa7fenqPCpLIyG5q8
1IoYZRz5P3hTBkUqQ3kWQYXcxzwCN6ZanVs3wMSN3owOCphEV0RmE7I4N7hkpt7w
oNZA+BHGGqJt9D2bCxXLqmN9HnXBc+SnvRnIsTM1rNfTMeWlDZnyuVFntgYyiIQJ
PXXpPkJtpg5h3wBdERjz9+hfVhxClMRYY9cCod6duCEiVVStIzQ+WfutY70IzZNg
XbW8cNzOrx0JRgZPuSwOmIJ+lOE5GT+HZ1xEm74WH50wyeABg4apX3zckvlviMEO
ARGiScGxD/8pP/3KuOC22JlhFgY4sgKwvBUE09I39oK4UFGd15p4h8ge4/kpnghg
S3WgiOxsW/fnsJE8WsB3XdRbuLjvSt1RaNvK/TalmXMUTBrPr12FPR7nzcwS06mt
zWltpPJ04ykbAoGeJm+Kwz7s7ixZM7PgEZzFLUiE6xSx4hRIOWOATgFMnJ5tsktJ
IuhUatbw85SCVPy3PPUWDzs8ZxJbyMR4xR7RUob5p0GuSrYM1tCOzxeaxjctmgdW
D1/wpjTnJTacguNEWSGEJcaAvPlDuM6FhiSnDukFNNR0VO4HOsCAHn+rcFWEggzn
3wwFGrPcXuuGbcuozSrNVqGLhaFHnH02WcvE+HLaCyd4pBkrijb/5/+y0uhDULxF
NRzGLFi1dgR44rswAlKpgDqwUURYVtp/3klQ2oHt1a2MBgyb8Xy3Wz6s6mp5JzXa
McjcnAieAh8oPFWzNRW7rg3LjGV/6vBiy+CYFetYJ21SizTx+QuQNCotRUM8zQ6Z
PFDq6diTo64ycZ8FMT1qVOJHK8nV1DLQeVognBQ4YV4ppjj7u6KYLl+5qeNdFupT
lanYYmbk1bb0PB6nN7Ulhu7WNUnqKZZWcCI0FxlCT7qcrSCd4X+M0F8E0vzLbyUx
ISv0RkBiP/ttAKN0u24dtFctfPNsW2Xkg1RPNAD+NEEUVn+yXakbqfp0kW3P741D
9v7j96fNmTK6ULchZkc7gCygyKOOgNCrFnKJpWR4rupXB077FZnsmlC6QqrKdpAF
sUPUvHgZ8X6vk6QJmfDtZ73dH/QThDIR81ggi3wTD/16ceo2m7Ky9VBrE3yfju2H
kvfS1ANxuY4woqgNFacM9/FnJIDxppLDqTtgrT2ZKCLwgz8/w0abrnTp+MScjI6W
wLb0uj9+soHEX0ARCSYF6JiEX6vDm8HxZpot2uI/R5qU2e5l9r7yGNAVRjru/9WC
J/2KEONvBDJQjg4zJ0EwpXNgILnmXWC+Hkgzn+A4bMbPXCAKUkL+VfaIg6ZJLdIU
JmOtY8kfr9OeCY8piKZVpBCpJVfqCgQ49T5iSfUn99pLIyLv7gWUdI6p07APeFFS
Lk7Kz0RfV3MzLGtcON/sMZTd9V4zjPS0Yo4vigwlUCqd+WSDWYn1N+az6V4C2nxN
1xqZ0Cfg5d3671PxHTD4gKEjGQl/KtFcHYD4g06Kweo+fAz3Gv4VwXmGR+qjOdtE
Uh74bO0VyM5+Y+mnrTZmNO6laHB9Eaz2PCwYW304zCH4lKb8QKmx5TpHQfaM25Xj
kq8anPbSS0oPcEXiYnRyVnEaenNBoP+T6cFurWNQPiCphqMkjn1wzc3gOt3uxK+1
m9EOoe0psNwGQu2W7RRqVVYyYzAtlsKV/tYC1wsRclRmxPs2acqfBgfbC+rWIq+6
uYJ5dhU0jAfcPKdqpRc/H3fvNmM0Kq+DyE251rcgM+Pdecco0f4WjIwv7C+bTSdI
uotySRzOyTxyvitmRLIfQoFIYGERaIOpACpmc8uFCAp+4oi59l/IBKgAmcLQ7G+P
s7V48IyZ6c9+6v+TnRlJ8JC8qQA6rcCbFUnmUScPj/idZMwqxDPapwLLXT3l6hOt
KLanEoYHdryVp+HIPuqZMo/zsk6LnPa5gH2m7BgYK0MNA2rnQI8nkQTIIpCK4hqw
11jsT/07rzEWSctmnhCUVahjXqvwweW4e7mEX5lDUK4Ezh4+eqX3UFpqmPq943uT
0w6iiGE6zVHDjcwjdAnMdYUgha2t4lLTdbsCtSdpTpJ3CggX3+z665Gl4lhBc1rg
91sgHK0dMSibOBo6zaRAIHnlz0bnrWNftQb7tL5OhsHBW/aU5y4CTMWUu2RwdM04
cYMjBiJHuc6uvqEatSHN2V0EtW4YKnAxfgDvU3ts0DXPOusIwY9VvYG86lvgox5h
ew7Deo02gmzmPZNh1qVWQH2YFAuRz2ZoJ4G6KslZ3S5h4VlsEl8MsiDuHYSdjUmf
LbiG/tNZliTWISiCeOKSH4B7XmbEmeMAh70/89v93u4iuAgKjgirzyMiTO9Y7SNI
HrjfQ8Bvb1f1zRp2mVYnhmvasaG37WycEsgRy4pwkt03kZM8zl0jIxn0zjR+N5YI
BICA5m8psgWkMASE6d7/yFoctdfjeNIc8s3dos4LNF/cSatuZdZGilO4fzYvIYB5
MG4ebjHh/yqsTZTMlzeEvLRR7+AuOeDGke32gBa8q3GqDvnPxAfCfkgoISSJ4hol
jSG9v/uDQ12k2lvVJVxY4R8gwDYIWcLgZCMWbHv5aBV0repmG+B1EWNoZpd5dl+k
DvJo0eCrYYFXzGxSnVM/dnEp4oD+BZDGDKSCNhM7Z3aI/xed7JWEuwUbvgoiNc+B
h+3GppqeQg93s7RYaJzf6Wn3q/e5rmc5jRRB7G+hwsrz1Qq60caMi33S2LVrR5lH
RqoN+eMik4LecIxDW58B4S+dubjuWxeKtxKWyBzuJ8s5gN7vWad80kvdxtPS7NgP
936AmsaHOz2SJ6PJp+AXcmYxwQXc0WCz6F7+w2mQf/2g42iiX4ZYvXcBLQKaJV/9
9dJInxE0kKOGgJnwveGSdbFbBeF2DdqayjfmjoAV3vsWmDYYdQfKaHfN+JygO0IP
7Bq/Gxkq1/efbcbKTOPukmTiP9sr0WfHR33vhtBOoRMAYVF97D98K74iQV0/HXdP
o49cPjpyQYKBc1U+QkqESucPaUAtp8irW82kQI0fVDW2x8ARiWB11jZO4znlhxFD
eNuI+qY+h4SMH4WH2vJkvSJRUtWNHjvEmg+ZSROvE3GGReeTDLeDGGYRDgG78LeJ
HOp40gdDNQFA7NsO6J+EyA==
`protect END_PROTECTED
