`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
au6VUGe+IkObmmpfxV6jWaUS9jjNbOxEEX+/40gAItVOW/oJMUeUnIrnmbLsIh6o
hFi5CdF+W10YjH3uDV0ml/3ta3t1y6DlG0RvhpFB+M0sqBXNIYEF0+dnZXXZIHun
MJWPI+w4mKfwmn7aFInzO8Uywd3lHeVPjFjCDry7NmAl8JZDMAWIg/m9RnkrHJGO
9LsRp5DSbRsXFczzfj53r1bnoGFAMS2t3zR3lbdsN3vWy+NTyOJoBXQind0+pMqu
YAkH6fWu2/suYVUrm1vfVhnv3tvDEnLrHcG0ETwH/aeqsWMFAY4BL9m6egK0tuWR
jpDdAnoIimlBP7Gal8+EJQFn1aG9oNqTIVp0URNQIb2386yk51MlkuqasmLJd/0R
IxBPfDib58/TsJs0m7SuOj314sAaJbgjhpwaUrKwJ0IBbEsOWSRyCqSqsO3ov57O
bav2mppYB00jmF6ZBHNEWwnod0l85GcMAJC+cbmUPRKoH0qtrkrVT1IBAwaM5zFe
sQiU4AuZyaO/MebqMdj5rJF1cDSpJHxA5B8Fq/XK/Tr8ADGKRf/sAOwqISaxwKMX
Tye4NidFYmBrXCmScouqy379XQiZvmul/lEQwBC8ofUKwACdblPlI+vOfF3S9pvL
Pzi4zJG8oISMKTSh258eC0flopXjhiskK62jE/trBR6GAYvpBlqX0BnnO0epgxJO
J4T2zAMFtj8blbfFzB14/AoAJxWJRuQRgmQE6OptIL7QAoyxiQQQiiC/8H7QMjz9
tJElPEksvZT/js6ErxYC59stjI+1pC4SKAet9NhDM31k6UIgUpACuA4q9PCHCSKA
cbLbJbGJ/CoPzVyeMXhvKuU/H92H9IF8nAejRUt3Wr1Gaynu7OWk0XNYTsWlFKR8
Tt3tDjBL/Qr/szTS7PFYZCgsbHz9p8rgUTdqRDu/Bns7M8xOsQxxN60nsMpG7DT5
tx6NPWXjSb4c10mSxPCKgKuNF8Jp5heVZIjTf/6pbHpbqNBsiXvMoCwtPCgfQ3qG
lrP+DbQcWHhQLIihL8jWmipLxJJFYVlc69o7EIObBaFmZ8OQGfvFHH3WgSKJGYSv
I4b2O7eCo9k8OVUY4suFWVlo3YKFAWA1uEIfZ+sQ9J5HArisye5vBof/D7gil2S3
Mvc4aIMe+I1yPt9LYpO/yXFxNQVV9L6/uLFIbEMjH9vIBm/ileMkccock8wVtGzX
4umXXwnFpJvGgQzn6xLklgpmrPCrATuQ7txW7VPSDDXMhUPWVqmkzzElntW2l6Do
6TZHDgo5GmPNYWgob1aUj4oDAQ+Yxl5JejWo5ipYPbSGaGpiZB2S2XD01zGs83FN
sFwwc7K+Kk5WWZjwRhlLOEC38WJOG4JH6GC6oJyzuO+4EadlAHRIGGSAi01m7BmZ
8KaiYUwqu5udolpe3JGxkCuaRuDeWFuC1BbuVM4EqooozZv846Suk28ZWjbwFAS7
4IoAz8WhtMRcyIgSYcbYmveEQTd5GXPuELNWTOyQqsUQjCJOG10MBG8ybxTdY7E7
UCFgpKO0W4Vm3qy/LadZdCc0GDqzpxjUiavxvpKOWPl1yn9JZOcqqucljYV7IzFJ
prc66b9izHzV4cQ0T1TrZMJTbOW3K6BcWYrezR0R0TTx4RcjwsvR/ByBPHb3PZGl
Qhyh6u+yyA80c2ecosS1C8tIgl+yoVFWuOMwQ2XsNL590Po8uNmQ+TUHFk23qjvY
hF4algoXgTw3etDXT6GnlxhfGpLbf9t9aC4v0eQdpYKb1CakZxCmUcPLwJrnUT61
M4P+YEny0nbbvCRPLc5R4eCusM+z6l0Z0HUTq1gCtEruAosBtsvmfe+IdZinU5w0
RfFl2H+0epTvDlWMdbYS49Er58AHmwI2MZuaJisiKkxMGJO+cjJwKN9LQKxG7nkR
JnMT9HP6y9w+xJI6mJ3Es7fHea3B+gN74/ibZ/CyOoq7Nfjcn4NU86kmJel+73w9
9wkIAoxGEsyWKuTieR6/wSm89jCHEqRdZR9XOyiy96punZ4bdHngVgHbeQRUIek8
G359ZurE7tdmsz7T+SNstum0xGr66VKbUiMN1+asDRP4ijhWJLN6rWnor4OjmzQf
gNwkIiPJjsW5/3Rc93+TBk2tRo1EaYJsYGv4JE8mCAlulUA5q5S+5MgCEM/f8P/I
piVLvVRd4gsXjz6W7rUHAOS3X41DS7HffBsPX9ipvPvFIbrSjLpwiGys+oKu60yU
f4TO1uCarjwP9F1zYxCrYsEZhcIuLch14CquSVOjNggkYSsGZnoNKbnQrRVFGSlk
j3DZb3sRWFnSU1G+QOWzhaThDmFALWDUzvKn8um9gV20x18KySPLZREdkpzkIe8G
8EOWzH37j9kGnu/ir+5twUwitx/ENsJGSZdQIQELFJJKkzjkEm1ZPyOL+2eEHifR
yl6mTzAtVK6gkSqpdPt1J1rbd1CGHWLIjKZU/zazUqos31KA2BosgTFhjowMVfes
iIzLZi1Qx+yVp2Mz9qIGMbb0bOBKSXaK4/0o6Zry0+jGqOK8203RhIxo/4QMgn/i
UU7KYhVYtrowrg+b3qAB+H+964nLPTP7aBn/kWE/Z5m84lQNDHJR7MBFixY8G7nf
SawSVLNvVZYcqfNHnOAJhLq+5izpCqlDjzBL3PM9Dc7Ui6e8DjpyaCSGKd0EzEJy
TGr2KE8hlEcbDJbqgxWKV59KiredvkXGOyHVd7foJll+Sdix3l2TBYB15Z3PhK9e
ETfiulytI55PEJMZREVNyodPIOQ22u9Em6jFsohDK0acOqfPVIMynwlUK1WGaV4O
UjbNpBBy109ThjEEhnJgIJ0rup0rNvXnG7wcgxle6G+PCz6gjyZl3ECx4cX/Sp0X
9qqHV4amZet4QWSUsQE9/WNTLAmJCkYPTHQ19SCUWHiKK5bqNd2d+IJeLXUE8YKH
kaC9yCZ2ztN5CLMdALV2QS5dtTYDFCmxBKA8KfGLO31RX6Lx0nwRg6PlCOEdlbt/
XIFGaz5hRiMjyWtnGsVUCZR5uVKBfJdoDJSV21M9KZy2+QQuR/CEACEX0sCIm3cE
E1iCnUuqDuYTuVcQmXUUKf4PO4O1afYCheLlr7WLMbq5L+0PeJaRVKhmpgg7elIr
e/7XD14gxpUVlZ99wQH74liLI+eKUMeXGdNjSuoEwh2p9RLGval25VJETyKWQY9s
5Wtw32r66jE4ZIPVXrKoYiSoMKJatXLdPb8rzROm1ITUK5b+bh6hRTcFJv19PN3Y
nJVN4Pp0Mr5UKIalF2X9AvYBqsbmJpzdH7yaEDNREa5H3jFm3gzLhjl0yKj4uxmJ
10pTEy+2ao0M0ItOkyYYwpKmD22jX1tH9A4tr3G4/zCtTs6gxK4yIoN3GkD5ml+u
Nmz3z1EiASx5L8z3J4QLOvBSWmiukQMtEOMjYw0CcjU1w6gtriaMwIBG8Ba/2gkF
POE9Z4jbdw28ByNHxa3KT1Vr88FpNxMtKH6yGV6NBhxG+CHGKT0Qv9bmLdIwPDQy
RBau5Zqt+XhGRVQJQl0BzwaN3qy/cr+Lp68cdbSyYIS4lOpgN2bFpCkIgAsPT6fJ
8om0xPZC9sdOLHZcy+H/bnc4akICI6mPTOx7VSrNRRzOfvFAGgpOoeqmBBrQTJ5R
KhsOvMYFhYKTcC6xP5/wD7UZCxHDr/5OLmI+RYFmBJbyiD9RzwvNm4nu8zuqMIPc
mc9xOIwR8Cfg92xD2zyRjYFh8gq4aR1aYgkjpayhchp+6dq+852WlEPNKUnmXDKm
payL5JiU5SoCDakyeeoTCV5aLp1goYsl/7QRR3sM7W0s/7ueBAho/Q320ZwHzIUY
Jw8slCQhUeFQnyTWIqs75mdxQIdpXy60I+pdDeIfrnmmBCDaMgAt/wHaR8Py4iB+
c3sj3i05hMs65QRlksHWsShdWtLd3G86+kBgvsCo9STW1P19mv+aYs7kbp7PVNq3
VJFrGpvj3Ix7ptqgEbh9CkpqqIPLfAlK4Nu/SCthGw397sXhSFB3d4k7J7YxQMuV
rjH5eWCoTgLquQBz4mt62W5XKG/XLmuDPR9bMs8TaIEkZpbObPnqLRtWscRY52xT
UTiCJVP3kgC7cVT6c0SNnOyvmmEQSeA7mh/rYbLEMCmmOB9r9Zf6Vr2MFnl2TBEj
rErNOkTlC5UdqcVP/AHpP60VIM0jyUGFNeytKqfUDl75AysAGjb748DZlhGp85LR
eZ/v+U/dYcb1YU1U0QKIJhOh9L9CKjz93dJZcYEk8tnecRC5b8r2n1fBDOAs+JZo
e5tiqGm1LKhys+b1DEJLGE/B2Ho+WoNj/5wZZ9gMfNsK/hV1PaPQch1aMsltknPp
C+2QREJHUde7dFtFaT8zCx0zUIk7PpxoefIbn84HJm6cw/TZGg79mwt7AyYpBlnC
zfb4ninaAG1n3tGXN7m9Iomb79a7gRtilEZ59RwC6R3LfZHSBfCz5TGVO7ti+MBN
MImssMSv5JBeafno9Q8oBTafbNUEjxqZX40nMLFFc+ENhi7TbZ3GAkwexo0KF6Iu
ioC+fN7rS3eABmbRsX3LG60YIH8r34c7VpNC4TON00ZDFIb6NX8a0OpHKnwBs6Vn
4ZjaIN2hQuDkHyQbKLS7gQkcnnzs1XPoCyNGiK5y3pVDE9SxDzI30KaNoyKBE/Pq
A/lLqSgwB24QDZyPJx8c53wndwEg33CPeUhy78xUzWoXOQzbGk9/bz+RMXXmwuCe
e9uf4dse3bm0bwB81bKAVeo7Hpp+qB9Q5UEpn4IBn0IZ3SxT6utXq3zWMuFasTBH
fBFvFecMVVu4iPuniui/W0OFatNvqfBl06f1UMCSgHAplpMb/sRVzR0/5FveIeUE
rGfT2rh37sovAXhZ7rPSZJd+BPDBNpOBJj1wpqS/tKP2nNhldRzaBUaY4TYj0wKu
W10M9zOZwmym+jqIGKIu2Zy0DnRTlns2AKBPugZmXl4DdPQZhRFIAQIFA6JtBh+h
dFHe+hy7niMAPlRGLz6wjnhbc8qCbK7elpSYxO6WYhECKvmnkgmcJsXqw3Fa/tWu
3dfiL6Le3FZmawSMj2+5WABEfsUXAmVmaFy9y12qTTE6TJ04SFO81JMiACijgfCm
pnA4asIeXygKAqiCKL8lybvfiPW2wSbAs1/BfJczNYxPDQMWOOFI+MHsnGSqxcWg
N47hXboxDCVMU3/ckO7ERqR6m+vp5Yu24pT+78gkldCmbLNcTjpWaPG+4D2urkfj
`protect END_PROTECTED
