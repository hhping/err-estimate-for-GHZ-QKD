`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cFJFVQU3F043mz+CMaVj983BwPyp/9a9CGNiYsU5/UKaTEVQI08hDlzSdqSQnXc7
bW2qI7dav3Gu4TqXOCpMamdrGezGSygakvrLCYUcsC4mkmPJ1fyUxpv/gumi0DUb
CKe8k2IQY81h9CJzU/wzkYrlLOveFAQ06qwAtdIbMx3CU3QjvTnpDBHuhuYL1ZuX
zJgaiuYk8BrO6tzzqBMfceVhWM91ysYq0xS0t1PZUCr5aalZSNjdtvy9vkjjwgyA
0fpgBnIw/TcYAyJclDN26o9m0Ufg8DBb4Xk/X2PHoUafT7HOAPE9xfPMy9Ofcxm1
rlaIQcbtyh0E25a/Ec1dQTUSBBcm2SgImi82JWkbT0edpH0OtJ48n8tiXjBlMGxJ
a/blAabRGGzEZck3E6zJRPOMrMQstn/yM2g9DdUjfLSdrmIkKy8vXMj8NWP/bi2i
pEZuuZPh2g1+Nuh6XbYlG09TnV9bxJsSkOZyqeH8WZpWjHJ2ocIOijj+X083bp3F
t2ZWOAaVYJ1F8LhkK5QsIWIaqivihMG4BWkwHm2LOBbsOrqX1rdbcGyax6x4Z3CQ
/UjK3gE4MBf6PSgXUaOcLwKc2S7ihDVwzrPOnlhnIQ0CKczHxrCuJKU8Wqdv1S6h
3KbM7wjtuwTB7b1ZZz2j2OzigBDXc7HWVlCsTct/zTBO5PhuMZt+aXezAivf1EP9
rruMKA3zyiTtQVLVI/3eZ5BkHWNNNl4A/e7cJaen5nr6rYu3HxvG2w69n93iBcTC
CRRSqcAt4XqwQJm6GMiAQJheubJmc6kvPURTxvfent78hvzA06adDRyJ3rdZ2s9C
RlvQIP4C2Nba7veEoKVa0KW/KQ7soHyZ3gHmvDt34xd2grWr1OJXFEu10W//4fmX
RkKyylZzjAwD77L/KC0Ud87lEf/h04rLkownK65w6kSZiKuqHKCBMasbBZAR2Bts
IN+sNAgyapUm1hRwtXpZbwo5z4C/IZppwyiph6IW6ZbL5tbYWGMRkOKLUEnuzAKr
awGZWtVcu8t7x2Wu8k5iqMV9M9X8fgma8NyVZkHbwVfkvhO0OR6VU+wMVdfSKj/A
i8V8+AUHn+TtF6m97A+hTM7xCAOihDd9GGch1uN8s6FSJ+1GmJv3EVsu4ZK2DkVR
YHh3gI/hd9Jop3FaymIVniY20lNvu5alqJP0bFa5zYpnw7Mm0W2nQDBFQyEtwzbH
SFfQJSI4rOXV5xlnNYp6wTcQmHVdX17LghEkHMY1jO7xzJPLYwlPF0Ic9VIrCoZ0
3qC51vFYdALcsURsBTIrSVEe/F2rDffboHRLHSQoiyHpZiNAckwQg9dFZCCEY85L
DFleyO/Yclyvkq1MQo9Kca476wop7cM1DgDCvJgUq+dm2lq6yPfeoUDfLG7/AVCw
wzpa4WOe9bDTSDQUIVB++rQbHAn4Led/9blRkz3mE4ktQ4NDjZ4oo0+23r4XN/S1
86DqaOmylZJ1AY6eSjmD3m1+CEmwzQyE7sM/FnVGENo9+QdOw8wekg8TLNHYV9fp
g+Vml/z0BgZjtIn1ht4BTqt483ncmCwtOGHOipkh2KUj7LqBB8kZXwRMeC3a1YPE
sJN5/q4Nr132docWZgYTFDtQ2u7NzIvsL9cewNVC8y8YeN8Bi5uLKdsdCbjKvrzI
fGIrN9FgsMhcGtDd9dRyWbDtFSwWKfAiFFh1tK22PEk/U9qZXFUEEG+xykpHpCfW
DNe88eZHUuOdablEM6g1FAS8bLU/9GkgYb8Mzynz6yHJYRZcp1Tk3NJHu0GNp6TR
UzDwGOJbZ6qd0JaHt1tDtyKR5Fi4/kmnNOUbFzG3btze7VyOGvyWndxqEJuHo/iR
/XJvT29oUZopxcpQgYm5N5lJQztRqRhW4+zAIOQ+sU//GXQWhTD7FmL40BPrX8Iv
VFns4HPDFkqXj/jT5zRY9MvYtoNuZFMOI6HV10MAOX+ON55rs1Mnc0/+4zyjWtyI
8x8hj7nV+TVFmhR5Q/k8CZ1d2ILtUazJthrfjICkCSouiMBYf2vMQ1tvTdiZPqGt
kqJ/nWOmDbJ8C7wLCu5dmWqAWW+UhR/oCsoI64/g5aIhzsa6KZkvP42X5LtUAdj3
6U79GTdS+qsE7QaCTnvGDZHYqmVJgZUnAYD1DVPn/giWsDTTt4/ao6WCdtnyq87H
6UxGPtxuhOUn1bbBWkXuFaGdO15E81O888n9siEK7QQ3NaI8jELY4xNZjqyDFJej
3BaMp4NS5sYd1VwWPB/lB/6ozFlrhpqXbHYXEDLK/OGo+xB3keg2110VG4D0BR/B
YO7zbuAdc+w3LytZeQiMiMCR2cjKZzyqNY9z53Ohl5tK5MZvpzixUieEhU0TqY3j
SwZbDayHOPKHNkKDk/jvNvVYwuVa+jReGjjvh64tg039ISQNlQxifBiU+3afjy6h
dcLYu9xlJmVulzv5OlMRa0DRVsEm+CSWX5j8ALIVcHhYIDsAMPRfGMN62OJ5kTGd
TzDgVCV84Gil7PzXVNunbbBnaFMharV7kOnhUu6SAa5fCMArZEJ63nBHIZekE5i1
F6AdlyEMdidbRvQJbhKEYpaLm5fIs2Bk7/FUbzSiawUQ73nRy15F1fIv2wuUOg84
hFpMe5OZs7X75zb6zd5xTF6Xf4AdpBoblsb6ZeA2LT3EJNu51NszUAsz3mgvruJI
XmfgsGHO0Eqnxqp8p7gN8W7cpajN2FjepBnjUun3O9arcaiST1h702BobPYQBx0r
rwoYxAsK6jDIZNgSccSDNGOVJqi7oKZcIIt+jsr98X4aGzZubuQ+ZUxjaBDaAcGy
Jrzjr9dOYzwaXT/JAREdczjxkLqo3KnCEbakGzgPzLWjIk+D5bGhnvTskPsDesl3
hAr0QmW8Phf2+CHE6i10NI/P+NWkTrU9PJhB2ZKUDCMQU9cKKZ7MtepFJbDtC/pp
Zjmul58GgdU/+fpGghzw0Jyw5TA0vxMU4sonN36xX4tdIdt5FkUPUZ4SZz7Y2ibJ
6i2YqnrKJ8ZPw/neYJ1d+CZ6mdrcCcTXMjBUYXldp5scLeq7zsiyvlUwdauEZeoJ
gqpfobdmlnRUcCUjCwfehwbpJbt26dkMqwKkVN1DszQfg2CR8ZYE1Gvx/xAWi8My
jBilP9EBuco2/EroAj92L68pQOcpVLwr3s/sN7z0+4LW0QVUYjuQ9xbbgPtjPz38
S8nw0CBz/xu4bGXhyeq0jJtORmARM+Zd/7olJxZ+701OGxCjrokmRw7fRA5rU8KR
PbR8737VYN6Boo6ZVLjs2tukOWvepTnKIXgxrhL6y/WXo4S4ShP0V5MyAf7AJRFD
+9Bd5z3eXECVNQKZTwPojeuDudw/PiMqablxEUe65PhPbMfz/+Eey2w6AvmNzH5t
ozLxBZkVKOawXsEBM8Gzp4OlbvmnRBJzz2Iq6RvAWWAf2XRT8Wqshbsgz7DJrvvk
xcu3b/bgdTHnOPk2N+PwiCWkS7s4KKXDUrxxk1qjlG1eoKn1kB4zdvIT4cRoSCi5
KDMFVG+a2HQ4L2y4iVe7BHq7bTRt5VXe6FBpVhQDsdoVBKl19E1jLUlynVY10UuF
6TVQf8OsfCnmFedLdmE/KXKo9FqWv8LgRAD73rOjPnh6LWy3KOY3U8WQeIpYQ+Cz
qXVfW+3Mn1P64CyAKiRzL3/tWod5unkh3QdKbdoszpR/8c+Q4a/xO450PLCbXCFF
nLhF0TNEOQO8OqmiAmY1sg03hvzaZeWG9GMtMSQ9un9tPbZhoDbsq1T0ZBH/93T7
YfCWAA54YSFaGpwlXDKpi+/BdiBOto+ECmrw0f8FugKq5g5xsXlEKuktzqH+EHN9
h/Zf+ZRlSqWQYiexRa73P768sg/hrqKnBoOq9OGgTOspsRK8Jw0xpOmfVSAR/K8L
pSeMs90wOW0xvJWOmmH+4ImbVk76Uf11HnHPwK9DbiqAMDiCWzONZKT5Ze9ZxJxL
`protect END_PROTECTED
