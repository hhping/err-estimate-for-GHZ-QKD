`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jHHvNvAPOnggzVCX4qpsDpJmZ7QuWfMngTJnp+0bP5lZs6x+tqJIb65KmQeC4uwc
UBrNOHFxzZtNf4EodNMqat7WOgV0rnQ39+6x3FmMh8Q49B7qR5qLdZCLrN2iti2x
6NKznARAL7N3JtXckVB3ZKGqSA92a+3k9thYAxWsp/zm2w7BUBngwpUCgMOzt8v8
RyKZj8qfD+WwLvj1MJ+W1U93HKMVtsp1zXspBrXDiLBpaJ69HEkVsyVAP96+oBsO
tfU1GhgueIjzNF7Aa601pOMYeIvOUxoSngJ7nlcFjTnDAUjDJjQ6xfkH9a4NUWdT
tpfjWOfSSJk1FzyAEkjvpIaRqeQNP84teDwxUtGYLzc=
`protect END_PROTECTED
