`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5eIPKxWoQJofAm/Ta9SDgIEn3M4q2aHqkEDVg9NpaXa05d6lSATtcAx5iYjQuWEX
q/Y1M2k/sbtqVj55HnYPO+WvDEQXUYjnsir5U2bqqVrBVmSidKScUe1kQF1HWOwA
L2O/MNGmKob/BRptmwjdt8HBGpd8lyPgCMlEBakT6CPHVRamQm+tGfiFN8Y59gSA
Xk0Ygb1aIJc9J5oFN+stAWVlIejIKfzpCzhIZxqcCtpONPhOhf+gKY0iIgOZvtcV
sa3Imz1b3qcp1CXO19x0t3hnDGRcxFL5M3AGesTU9UjWChIwzod/PRwUOBuHXms7
SScmi6g8jpm2tv9ddrURzqleL0gfrINrXk0TTPuQlED4mnNwv6D9dArFvphjV7Xs
AtQE7VHYWP2UQNBva7cE7q5QPurEVF2E1JHxe8G61F7lYpsu9oA6isL21UdIuuKj
yqIXHQjxw2SAuEhkjqG/7UiJkAb7cFSP5LvB/F9Jg/RI+qCtnIi7sjnZiWxdu5pB
ddI6igQOiw7w78XWfJrEny3WRQV6CmhmcFCADPqvanAULQ6J+QtQaTGAsdglJ+et
BJpZ16rW7SoG3PfTNf/nbWAn24svoAs396LEZTW1YXbI7ORcHkMzzEMVjYguVmyJ
f1IWGxWYFVf5JQdkB+zhjlx2hpojFpNNY17XSZQ+8x1nOq8g5B8RxTg4QNpX5CCP
WOcqVeHzHOzyiXMWRfoizTmNA4U7L9ijcZDNf18ISwUt/PJn153rOtKo/m+b+DTB
8b6RdbxlSuiG5T2K8BqrEC6LJNPOu4fCqpGE49OknAm+Tw9Vxzw4f6O5SOlw47q4
Af2m76iXiGH7sSr94aktzaJOPlNIYoXOEwtcdmvrLpdgWBSFhpo9x8GVINiv2ufT
Gf4RsdAVEganbijUeSHvGRg6lcrGdOKy+6aky48RyNSxjKFwMDxhMCLaGpiYwMPz
1Fo0vqa5H2KhWY4bvTYeKQYHcHMMmpzZHkcRQfjdFg6rPIcyXfCRZcee6JihFIee
Ils6Z84WQFHpZUNgEXNqBujFqqvMBtvMOf3uI6mA5PY56hUtpFzgHuAs34JcWEmG
yhcTQflgWlg2uOENNoCo04MX89IiVWZyxJ+/LVZEcPEQQdUpycNtMjluOKATL9cw
h0pgccJ6lQyHDeUbLKAaEiW3mtfvU2iHP1lR60vQ0jw=
`protect END_PROTECTED
