`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FP1j3sytZsMinXkvEf/xTcxp3KOoq0OD3K6QK6lJW5zcqhue7onaxrnqvjZEreyi
YSfgn0QyEcwEWXrUN1guvJM3HYiDuLlLVEOggaQEmkfpFPmu/RAEMOAbD/PyK250
xpMjH7XAACi8jRRJxYqDlRS63LB0vGYODjWWu7za9KjcsavPY5tt6ZwS81LDO1Xb
qaXT4jCtgJvB1PpN8c69WMfkrspU5qCRwivBeO8xf90fw9stp8dJGzwvTIS8Q+ol
+uQAy4G8MVkGLhTx9OOCLsc1cOmtKHg+RUdArozXo4nclE+1jaApUFtVt8Glx7gZ
62ZPgAcQRjVQTtEKBf/mtRPrX/FHwavuD59Svmpb+n8feaTfdz3Xz5mLLRjipVkp
UMrqPMZFJC3K7jbxyA3bXK9wp7PNiVJGWO0iMf/IJNa9tZVz6PxzXlQiHcr+v3WZ
Y8vfzB9g+JCMcPrPUC/aUbJ45IuJm4tj867FuktA3OH4wVnU3l0HMSq8R7Rt2oAz
vTA6MN/GzvHw8IIm356AgJIa+0Y3bsrcFFL1QjcyLuDDGKxj0h4qj9Tk9H7OfRBY
CSM31T3iMvzLP3AKBtnel85NSL/gOiLuH33yG/beg7Y9+taGSuGk+oanHc4qeFUo
o3JsKF3Mj2ZrfNn25yuVaM3Uvoks1BHycKi99oKKEMtERtgyDHJqIfonKmEjj0Vx
AtYQmjDf6BPUVQMUOQtDNFd+nGjkUI6CnsrJQku9AY+LbQudB38WiYktt+4JoFFt
zUK3Ss51dTVmQ3Nr90DXx5H7R9Eosp42cnSslOOAAVFxLgbH2QwWCOf0UqxctYfR
LMHhunnif/Y7nAysZoVUPUShW0Bul5/IPSIks2SlAWHqKMxphUNCw07IcqS1QnA/
tLs9Oevwm6xIBbBf/kZupEGwlax7QJ/KsybUqDM0k2nvZCx+ujgNPf7WnYT7Jz8y
pLd82+iaIMnlMAJ/CjjdNS0c8Zmr8YJ1uJioX48WOIczLKKGDpoG55HaNoe7KZf3
JAQK88C+vKrFOSgxSyr27kbkpmpyWRoeWq0U9SGn83eyTqGJhYbyPwrdjipyTp1r
GRzBlyzjzahTM//nzjvA1Df0GdDszhORFsdXm+tDOg3YluLT1f/otTqDrj/CG/E/
RloQ5irJoiNowLgM1xsHLVFbN0bFcol2BDJlTMokt0EKUnA2ZpCriuW6zuW9f9RM
nLgBYjFrycalnvhFpPl3G49PWyRTdNEj0X7ZcEnsogdqmRMDg/Msf1Fdr9o8Evi1
LMem133xsRBUMJ/obu/f1qOLpgFRLdlwSjnGBXUK/EnKj2y/cDpvqrly12FRwDVz
3boBzFH37fv6glLJWsmOxStLphlpVjihXvqJv3t3xaLj6bxn6xt/CD1oje40LUIQ
0IwVix3bRMGaPalYj7xganeKbTqWEhBrmwPuioIQNWYdT/zKzSRZlGiedNaOjg/M
ugCNBAhzjOD/5FqBI7R13A==
`protect END_PROTECTED
