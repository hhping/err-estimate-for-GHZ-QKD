`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
77QSSQZd7B/6HXEB0SF+DF6TNySqzQvQiP+xKAYh1lrhDdCUk/CdHDb2UeMpfQk1
oSmMDmXiIEFbBzlrU4RUxq3SQ+agZxKFdOWAai9oBfyEgup2kDc/64NfzA/WTLy1
Q35MLqDIQaNnUP/f3MgshJMUp/UOLfzl15U35Bq6kn38cTM9JSkJCEQfL3yVyIa8
GQa/4CKjai6cCCX9Vz8eZNjh3eNSKo6C3wm/UK8Y1BB4Nv3WyzA/MQH/qi9cJWV0
+fS/VovQfY4sZ4+P0txuBhDbYsR3YkTOPyOj8JGQ6sIOEQDNJfVHAFto9q/QAMHX
LLYLmNKdAfaGbk5H1yS74H7K6hnyKhecdkv68cnn28SAxjOwhf3bxUuxDFB74FMT
0Jc1hS/w/X4xLMZcphV9oYwSkDjoeKDCHq/wsZ5KhH7BGTbH0YtDEsQl/iAjpyIb
JRyaW6iK/ym58vpaJHTjpDw1ZlujCAu+8d1LhwEn4b0irVRTkC0s+SnIzIHu77g2
8Pa2qnZtmptPamjDauu0s6jD+J8CXIDIw3RJLQww3FuoE2LhYeqgnYX+RVKy9Q74
jBukXWya7Vk39qW94Cu41chK6j2u2xCDKHIKAaV2awdrs/1uYjqI0arXD3k0A0Zv
3x4qmOaYR8qILq3vFJVO92iJqUk+7cvbpREC9by0mmDuowgxtgn6P0pF4Dj2LPIO
M6rzoW0qZZ6YvK+k9M7+J1xga5QlQQykPNd0WQYhQs0UddxW6R0MwbVWk0oCWWSZ
1fukX0w7EnCnld0VnqxdxSoG0DP7ymsEq6xobnJRAQzQ4ecnBs21F5JC2vfzCbKt
zqaoKnZAl27/B8PK7QN9SJRjDn++N4VdkIuIPrjPEIk6OsEd9fXyfI4B7pNoszIe
KmiX8+Ge3LU1sRAX4VF6/rKeQ6DLQ0P3zVAoY0Ugffp5oJZcnZjzMEkRR6nLYtay
X5IGxrWUlptx33JXnNwdovs8Nt0HqkF5DYzdrr9i05RbZaelKa+/3+INZaR0qwWj
WZcaiaU8s8CyaZ2pGTUygl0IRz9iBHjzJpV4NC2pnXQ23plKZNUKxUY7MDsG0bls
+sWtZvsGRNk7P28pMBgS8M0tDfhDUx+7swL+Jj+SEk7KepJrqzl5+T3++lDIHDG5
SP8E+KiF6j2NM1oTZ/a43VsaCOqxXA4I6KiQHqOBNN0hG2yUDENzQvyfzgBNTe/6
XeTz3jOFCokk0GhDzK54OrSA5i3+sirNE7VUddAFxOGZHEIX7MKT9oHl7uI3O23N
6kcyyC6fiNsUhFXTN0rXhjxd4k4/EpeW4KygWeFil3cnVTc12KEpFSXXFpDBNz1+
FVvzNAklZdB6TSnwwZ5VL7D0o3E8v4IwMsJx7aTVeJqkx6OaJ9as0F5OC3hjLiWY
A4j8vngythir8d7JjEVEmrrx7ZT7Wp54ITCQr7nW0xbW0/91/vxC3qQSPF4p6abj
nNPaKlNZj4o/Wyo4HigPnbUirxb++Q9ElFwMHzzXcyUN8QpSaqWaTATSem4cEpva
LWiejpuqxX18ZAGUIam9kt+Ijj+PDYQz4gSCAjg4ByxkzgERrZAKQ2CPvFN3Oxf/
clAvFD56K5bCNizqJ0biTAqI3BKmP4ez8yoHpFe6OtwMwR12GlRcd1ja9UMLe9hP
FA5SwjyvpqSNPdt0x0cHpPoTraU6KQ6C7A6QcNrXqLgCu/FBidZpoY3MDg1zvsTa
7+/oCugUUciojosDR838jCm7nkbWvpLDlIEl7HyVdvUg/xlNarKtRS4tfZEcdTa+
RqBPNIKWh9TldzpIMUEJcHENRI4yi+T5KVUPxkLzmVnP3aEFr/8NAdQdQsht48EK
A8VoCXOCBibN77oiVrjHXPSD2RknHC80b5hCYpDB+HtlSWxv3KlJG2RfSO6K1D8m
PTuOHM6AUX7u0JrEg806v/ndmQWKrtDPvtNlM+6VZk3ukO8gmaq6GEbkAxtaJ4Cj
5gzBt9eMt932DclmzbzHkmmvYT/ZOPNk6R8ZMqEvd47p2mr++DIfesW07npTSAhA
Q8XuqB7X8zo8IQEpQZXJo7yITyDJfKBITj21EA1S+0CTkro+Y306/tvLxfUAEugi
cmM+UsQoBnNSDBw3JLW6dM1267jndSOxSftS4rkmFi5Q5X3X4kKV31ndxLNjSteU
ftlMMxkXU4ilUPKWqpYcvlsJ8ccTB9W8L7BDTqxgKDHDON4H4nwjjoj402ABaUzA
9c2JYYocTBdy72rAgZpCPRZqsONva20toisZH9WU/hxN0PGqivYR4XvGbZhpp9a/
4Y5x2JTUbo1q+sRx7j3Wy6FIIzpUe9eXqLdnWRIkSjkaACRuSKh06Rz9iDQjM51Q
H2f57zNNs5Nc2QpFTezF6AFLeJUs2L3ZGQd2uk9UmuKGO78UY7jG2XYPvvAtGntY
GIcGLtAM07/g3wk2GzKamVei59Dtb8rtHWzJ5u+QTotnVIWJgQrNX37aBwEHWldO
xBEBGT/oK/QpRp0V/c6llmQx5ZjeawoWnaqI26kT2oBje2Y460TXihp23nQSlZ85
vMH5pIUNYjpRmVfD/jWilJo3l1s2s8RCfnnUuGNew0wrt38GzmmefRgYl4I4r/K5
a6CSJLPzbFGlU3D0MKKkV1FStHTGHXQuBnI1pFrbAzB23rRD08AvRKkkVJTF0W2Z
SEhxNp9g6RuOQI/R7xXGyDuQk5CBxzc/ljmudfN88jtiEYN4/e59lnY6m10Tg9gp
YaEz9arg7keWJ8DgT1VFK6WWgl/2c+eGRHI/ymiLYMMvHDytMlbLMqSL6EX8+6HG
L2PuSwtG5a9ri/B37npaXPN6CAImTIoWCXf28Lbp1qisvBXPQKBhqmZ+Tnnuqf3X
iHTdYctlyA5NdUb1DaSlbPBnBXxNsiecf5qQlMUIUfTuJp1YOhyqCKYQ5m5Sc9wB
4373GlLKgwUqv8hgQlNnDYOH79ntCqvJ91CH4uj7fnMwZ5CB/ezva8CTxGPQHWXb
/SXCek7qwwhO7tfg9vJyBFgSRpX4xJcvGuUJwVKDJVn/8SkzrjfrAHac0YDmbGDz
2JTOnrcFXSPljnM0rq+yUFJFA27nSwNpCbEiGWTtlazirattkwUMYjlZ98u346pA
ooSI/UXBME6/RpSTzhZP0zvGWVohQ2D4I3Vmr7Gco3IaTS3QC5JrWeT2HFRq9voe
0YawoqCZWIoKCJBjuN/GcGiOdY9KptPQ7Y20/RLm1cye/xeWww6peg5cE9euA/+D
xjF8hI4xbSdMFmSbksOcEv+3/hiHzLxHpXYmG80T2ujvIkinC+Xg68hhGRxNXlkH
3KedjQtwDRz8PUsMJssI/WgMevmX4SSYZTX2H81HZamqadylWRSF+zJlOoR9nzAr
f4/kmP9MPZk7L2Pu7TPkXjD9nki8Ux9g7bYfRuwSTXcgM56eNHP1YWSWO4RL5w+o
MHjvRcO62wOsgwtzUEQfTWfSRYAmIS7hKZtuvMCykTDpFbnFZkQVcKzr/PY3r6rH
pPmNl/GhvYCAwGtRv7RApDRXKK0iCztSrb8OuxORKjjDwSIrjfHIUC5WBLShjR/n
DZF2ewkVo7aGhm86uKdm28T3odT4bQAlHzziIAKihbqEgD9WAEU2YIEb7fToFvsP
FnB0dofyZeIckMP5gaCep7MWVcTQV6AfP0iQKxMpBmjArXjpDEgtRp60M91gOuKJ
dDGG3qNusSPk8r8oigCDl+6ivEsxSucFC5ci7P0hfDROq5MrXIZ7Bk89p1JWQDLt
tN7obK4yC2XHnB8v/cjTpXQZwlCT75KiGQzgD3FGaPH8heBkblDItDwESxLfYHpm
mY+ISFzWiBjqCzauB84PkmmW8/n8Dg3GlHi5Um469XngDfdMghow0SAO5IMsU7iv
CTDWTXVzzUMAz2+vtI//t5Rri/zYbYnvGCzXDjZt0hRrvVkGTHTHLiCyDgIsNk17
HQTb6Mi/PYsLHlNQ/9hJdb9rE/sdYDil9zeLYQAWC+ZwLBsG4UNjh5J+6VeTDhKk
auakAmyRxZjlexQpg9nRJ3FA45lNXR/qJDIR5YaqjHepIUN9fnltCKrUrfHHdbRW
wuy6LQV4r3kXT+DtQCeCERfUjXF1jT3PLTMhFP/ukL4l4cFSvIpN65HFCF/dZ0yw
brQJnyehynB/5NNbADj8gZDPCNy/p3X51OPXPoK3afQsSsIjyBbRedO0xgXYDcRH
5aIoQT+RC5bAidsY0Vjb1FtrI2C6U25/umWzu1otDaSNa9pzPbS+iBFIwnV+3WVl
CKEgNrDB76i+bLhJ/a9bwJCS8OEQnqpPL38sjKmknVe9ZDJQrqWyEQXbSYbp0fjM
ovsFnIYGDhE3sd2eMJ8/I3T2955cTaN3nf5tE2pdzbZjmrC4bBzlDHPlpdFas0N3
B2HNbpSNOdloXUEvCFIbS6HiAL1FfnL+4Xo/XnZvOrAeaoZTJuwWCQugHnErwHyd
Rzbiwe86+uKp9GJmRTzVC7JD0GRGDKknm0only9RvhXV4LY8OUAi84lw2ZRDHEB0
2Vnxmpu2trgHR7Ghc9wOBFn1nUMrlikclgn7JG5Ut9a4dZ42RqAtkURo5ElF38qt
faWXr/ypgPQfMhgvek+53wkIQEfD2OJpAhDLboprB+dyLlWfR5RTRkeuLG8teilO
5iilBUxldvl4IHNVNVfJGlIxp6kcgGcDCdCWG62n57jI+DaPbbWZ6miOpifUndVL
UBMn5U1/H5zMNucHvQTN7xGvbm0/Qi6tDylMkGgR0mcyN0YKg//XbT88ou2YPC6n
SoJv9mK23qS+VhlYe7PrgYV6IUi9gaCDaBCYW6S5fgYTPpECc70Ur6wiVIB/J+oY
vYKC4gIkK+4BlGtLhoJfjL3UbcXwagSWi52UzULUiLp1fDdhzr64n38398JKj99S
6+CIGSRG5arketSR8mK/eud7kah0ARfMuj8WuygSkYZOwZ0XzaomIiqT8PS7nvwT
UwU+QU+YlYWXHPbcHyvBZ8VXGhxW5h8tKpszH5mgnTQDXhHZUngnYiWI6/xuXy+Z
UF0IrJzmO13JneO3zPr5BVvNfhd4aIrECZNBedCTdeGc289+h+6nrMX+CYxuZdCl
MK1VvIXNOU0QttnLJhyZGdDrMoAnTgyxID0uqbkeN0CtNZHvHh7xIEzJ7T5agQB7
TtxjTnalqEUPK64fjyNu5snvYPLk/qn6KJOxs4iS/fx2JyrwyixYOTpMNQxu+pmU
K8O7UyxT6TsmgnFiqakobGNBDa6HpMS3NrzfXpZvk3Va++22YaSxnJu+7xGBrJr1
Mrmf5+vhNexbRaocOJoyxzH2ictL4fuibY9Z4Oq0gRYO1xP+J3lKadnK0GHCvUp4
kYs6GapYNshKsB31FkfCZtlpTbs9lNzpmMiO1sBsDlW2jv61A+uZv+9708rR88IF
WzoNG//SYx9hVGPsVvIBAQIa5BYzVvaQvGFvXEy6LK/cf5oPw7+uSm/xtcQOk/Z0
ZV0jRnmWktuYjDpL1STr2gknyqNjtkoWKMjuKjLNhZlVL7uixvlYBy/0LB4wT8Kd
+4db3vFibsGbRejEpHAVGDgmKKbhAs+OCwuvxe3hrN8+m+W7ZVK34mF18y+/Djxt
Ws8yjucJLIkcnfay0DoZo02Kre3wEZ/ln5qh2lWJcS3PUfO/Ry/PkZnRVsQsTr+a
jwhCYHgpnDP5Kvp+YjDSjI3gYBGiVKPlSyuluNTH5xH03zM9wT21AXMpYU1mmbxV
cm7vJD8f26iGiax7ii/uTxQwY13gc/egB3R7Vh/eUB+RJK9a11bhtgIW9bV6I60D
rtUT2SclIhnkdcRi+Zqk/tmsRTS6fTPxiEm9Cg2JhiGjNmTAEDOt6zb/5fDJCGGR
Emc2HoLdf4CRctwpDUd/h2oRDANBz8t1jXqAuWig28iWVuNE8HYEBFE4GygIAq6h
JeMqenyylPSFlV8s/XV3qz8MkhAWtg//fmG6sO9+yvK2nUcQ9WbEDJw8jY3SQhSM
IOtwP28fZUWU7Id8vmOb+TzjyjuW7NQxR2ZvtMopEMwIlyYo+xaA1q52Oj8CCWW8
66mytP+YWgO72CeijZlE+K8TklEbQBlXmWH+j02WBXzzuqNwkMdX4bmt2uQMSkZm
/JDIfmyDeVHMKy6k+XOC4E7LkBU+ZysGpPVKSAjhsNwVIPpR+ClXKD+naXIK3ZO7
DAIvH3jJ04Ga1RDWSLeYR59AlGImQ82cPf9iNLAk/wrCsnpXHmIlvfsjAxR7Q2HH
r1yd6PmWVrjZc8W57eZltoL8G8778o0GusxpBu/SUtMrP1i222csyo0jLf8nMUYh
09iTpR6H7ZvPMfiNW73W1PWcgW0RQEgmeVqOPMBVQotPDSN+bebK25baSZG3bVJZ
YE1tms9k9q5V8EgMGALkwzqED4Ofiy3JMWdIoBaHlZ6mB7yqCsucJGlgEWTtCEEX
wiWHnrKOeeEL2deIWW/KcyRZGY7ed7rLoFBsJPi4TbdVL1Z3VcYMY4eACNBjdgYi
mXDeNSXi3iIunUhEb1WsjowrNTKTdBGMapnuXEQU+e/yOA6qgeSNRGodCmH3e5bM
UBiWhoLfsrgfjx/fIZwidHnsZGUdIC2FsXdfIgWDGWUk+6UJ4A6ubmhwI0HVnn5S
q7HsOxhwZRqitnq770vGR4G24eE6fXDdIIbm8eWzWEkYz6WrMHsHIhdCUJwsUph/
UnQN3L4WJugsoRmf/o4TvAA95ekIoB9WC8HlYjEzusb32W62z3yxqJ1+47APMCRc
vBKbrSbwIwSXQ+t8wyGhA0QTI47xPvg8uGAcN+iVQbxKpUehX/JeiW2JsQqU6pKm
iuIkKFspRawwew69gHeFDCZV8RjR0ED371qcgs1puHDpzYh1RRyS0ePA3ityrrvY
jSyBgFC+ni32Y9eAX+YGKHnFahNLdJYEGb+RQZH3Uz8pwUvD6AvhItmLMPpuGZrC
RxH0IuyWClnKI2QeSONcaIoKEv6yoh/h8wD8v39dHKmtnsYcSVfW2w8983ZbvfUy
RBq/yTV+5KkU0PCAWn2qcLTxLtFe6Nlmmaa0xcYTh6KRnZp6qwidEFTtD4hIcrW/
lAYL3kevq61bXTCQh7dUtOKgTKjzbpaUx4RlCEomjO8Eku2QCBAyBjzdneMQTcX0
XHr85ZpVoBEcqIUSRYHY77b5+M+txaTqsGnPVVN9rrhPur7fVGsU1ZgpP10UaUHe
G7+YbGXmjctMyLad2kIDF6lKgNSC1Dr//+A8SCikuLmonUlmABpdARGhG1Y+5p3B
8yurBOYHIwBZIVo+ZDy/CAVAZ9FHpB9Sjs8s9gx+udqORs7S1L+Rca14O2uuAZqn
sHj4P9psfQlyVMVOz6M5mZxpRLUElIrnJUYmwZ3Fi4wDh+T29ZEoPrz45+dY7uYY
Op60To+oKfwX7sA9k5A+z4xZqMv22E5ZdtLc6mvWW0p9mOXL0JU3BwtAxTrTzqO7
EjAzQ3+zDwnrEDY+AI+AHhjHDbiWei6XvqevSXKP2I/MTY4pRono/VKonadWFNFS
vYCFJHpfwODsQLrw0ghvqwjIhKoNOLygjZPxdY3hUy0t1oMluKWt6i7HMxz4JiQb
T+Bt2XIJ0x8C80gzaZY/CwyqRy3L2O26AU7enDRTvmauy5fKJ7JocIHfCGwk7Vw1
R+1onApEcajgHUg/K84a6h6md79S9RmxvlWINEn07TCExSTIsS9x+cqk9cTnhnLo
GfqxOJ6U493HVn4SEm/BVv2A4dcLdaphOfFN7jiNwshzSUsEuZeD7bqx9R4uqT6l
Gxb7DHlIwV9OyOzpYc+BbDg/1MLC1CqiVw5TvGWFnIquOhhpLRyLUIJk6TvNTV6R
NMOFdxLB3oIcu5qaJ47B7c14c0I9dNp2R8zYkf5KuZJIsR+x4OpFohN8JjY1O+Az
b/dbr2j929QoaL8qUjGBkgtQE/HiDD9KVTEu+g0xDBPyx1/SRXdFBPsV6hxMJW2s
ygeDTq/Mqlsb0oOl9lX899oLwL4lzNBseTgnaskyD8Go5DS2L4E97zdpCPGRHJB7
3ex0In/i/mmABCE8ojHBIBXvpQ4kj5gGRaXZRp8KHr3ycOq/WzWunLtvS7HUF4LR
5u6/BKKYunSWJHnNplHP0HUEp1xIWb13toVWfGHuUyd/ZQAUHaJ4ro4Jmq+b/XtN
o41blzlwijv61yHUuopjZnN4oxu6BZTw9BrtvJtlQctpuA09nNtKbrpsz17Xl/VR
KBgEeERyA/XGPY1a1CuEuitXeo2gFKEkjjedBAjy5reZ71pAfq8A9UhozHsRIMMs
7K88PwkptWjXxcOFmxufzvLKxWAE3B5g2N4om3qQxX7CtVcNAU43Lcd/K4HWPXbs
dh4+TjCJbnRx6z/5mY44A8AjA/KSQIorpMaO6hMCESF6DbaOtyGSATMd4kPgK+aO
+xhqwT4cAnR0kJt9uqnxzT3ENAc9OnLCmwb4Mg+dhWFe9xgTeiK+LByYeDMjgvcH
brZ2H9Z7iMM4vKGEH+Eamjyl5AjEz/i5SU++crcH1+zfWddX/e0meUDNK3P15jPh
Iyozd1iPYYbVYX6ZujwrdXxGDTNhULSpzN/gFSRGqJhPlpjt+/4QovV/PfpKG+z2
W1GF+4680G8WKreGxys42OdeV/Cc90DB9YLBHjQXaWUvpvhF2QJ/ohjxj38SEyhY
ElDy8FwvDSsHkPLirj/dF+Ou2xGdJI9Rhxf1inqgY9wszcT0jVgKklyG54PtgarG
uh50dakougEhRV6RVN3mtc8TvZUjqoCO4mfhzpoywjvP138wquWTpvHG8XRBTGtT
yD/872iB2KQddgpADeSFtdj4ReyNs6sSp0wLvUFx4q31WqHJtwfkvyKzvmIqpyFN
Cb0daUciUgfhbv/5zBDvXeMK0n541dPekBRb5niEkc1pK9YIHsG8Dvbxc+khnghK
FCnv5R74XjDJ7cIq7poCwTMRJMKBHVOxpr2ec/YZIwyvSnXu5ByUM1nYMbcTu+O/
d6XPOS/zagAHx2AYCOzmzMZaF6wEuS/AAFPlatp5s+U=
`protect END_PROTECTED
