`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b8YazTQS1+ZJxgesbpnYRCTmDubYjmtH9cLXpkSeo0XZryUktGbX9Wa9Xrq1DQRW
PBDDPOIg550BuD6Y/W2eVTNhD4OwdHDUCmWLUWoPUnT65nLVvUsYzeR652SVomAj
Qiu3nTAdWy6UlJPYDsRyQRwf9dvvlDGObGTtaZZX6tZEGKaPSHYVQ2eTzwzSyqTc
4WllwDY79kMS1fe9GEUGU4BlxZVjGe79QZcCkRL1FFyujd5lZHck0zX4nI67GyVe
BVHZljAlGZiMNV20kgSaEBxHEK0X1JYHN27gahpN1yos0mcNfb3Zn6foTkU5//WJ
KA9Y94q9XDwbNsLo05W+44xqIzM4/CN/+U2UGZk8DvOp0cZ5VDufehciwuvO5wMA
OpInUksjkBolBGTgaJw8qB+YES+VYiIFSInqioZiaDU=
`protect END_PROTECTED
