library verilog;
use verilog.vl_types.all;
entity twentynm_hssi_pma_channel_pll is
    generic(
        enable_debug_info: string  := "true";
        analog_mode     : string  := "user_custom";
        atb_select_control: string  := "atb_off";
        auto_reset_on   : string  := "auto_reset_on";
        bandwidth_range_high: string  := "0 hz";
        bandwidth_range_low: string  := "0 hz";
        bbpd_data_pattern_filter_select: string  := "bbpd_data_pat_off";
        bw_sel          : string  := "low";
        cal_vco_count_length: string  := "sel_8b_count";
        cdr_odi_select  : string  := "sel_cdr";
        cdr_phaselock_mode: string  := "no_ignore_lock";
        cdr_powerdown_mode: string  := "power_down";
        cgb_div         : integer := 1;
        chgpmp_current_dn_pd: string  := "cp_current_pd_dn_setting0";
        chgpmp_current_dn_trim: string  := "cp_current_trimming_dn_setting0";
        chgpmp_current_pd: string  := "cp_current_pd_setting0";
        chgpmp_current_pfd: string  := "cp_current_pfd_setting0";
        chgpmp_current_up_pd: string  := "cp_current_pd_up_setting0";
        chgpmp_current_up_trim: string  := "cp_current_trimming_up_setting0";
        chgpmp_dn_pd_trim_double: string  := "normal_dn_trim_current";
        chgpmp_replicate: string  := "false";
        chgpmp_testmode : string  := "cp_test_disable";
        chgpmp_up_pd_trim_double: string  := "normal_up_trim_current";
        chgpmp_vccreg   : string  := "vreg_fw0";
        clklow_mux_select: string  := "clklow_mux_cdr_fbclk";
        datarate        : string  := "0 bps";
        diag_loopback_enable: string  := "false";
        disable_up_dn   : string  := "true";
        enable_idle_rx_channel_support: string  := "false";
        f_max_cmu_out_freq: vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        f_max_m_counter : vl_logic_vector(0 to 35) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        f_max_pfd       : string  := "0 hz";
        f_max_ref       : string  := "0 hz";
        f_max_vco       : string  := "0 hz";
        f_min_gt_channel: string  := "0 hz";
        f_min_pfd       : string  := "0 hz";
        f_min_ref       : string  := "0 hz";
        f_min_vco       : string  := "0 hz";
        fb_select       : string  := "direct_fb";
        fref_clklow_div : integer := 1;
        fref_mux_select : string  := "fref_mux_cdr_refclk";
        gpon_lck2ref_control: string  := "gpon_lck2ref_off";
        initial_settings: string  := "false";
        iqclk_mux_sel   : string  := "power_down";
        is_cascaded_pll : string  := "false";
        lck2ref_delay_control: string  := "lck2ref_delay_off";
        lf_resistor_pd  : string  := "lf_pd_setting0";
        lf_resistor_pfd : string  := "lf_pfd_setting0";
        lf_ripple_cap   : string  := "lf_no_ripple";
        loop_filter_bias_select: string  := "lpflt_bias_off";
        loopback_mode   : string  := "loopback_disabled";
        lpd_counter     : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi1);
        lpfd_counter    : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi1);
        ltd_ltr_micro_controller_select: string  := "ltd_ltr_pcs";
        m_counter       : integer := 16;
        n_counter       : integer := 1;
        n_counter_scratch: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        optimal         : string  := "true";
        output_clock_frequency: string  := "0 hz";
        pcie_gen        : string  := "non_pcie";
        pd_fastlock_mode: string  := "false";
        pd_l_counter    : integer := 1;
        pfd_l_counter   : integer := 1;
        pm_speed_grade  : string  := "e2";
        pma_width       : integer := 8;
        position        : string  := "position_unknown";
        power_mode      : string  := "low_power";
        primary_use     : string  := "cmu";
        prot_mode       : string  := "unused";
        reference_clock_frequency: string  := "0 hz";
        requires_gt_capable_channel: string  := "false";
        reverse_serial_loopback: string  := "no_loopback";
        set_cdr_input_freq_range: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        set_cdr_v2i_enable: string  := "true";
        set_cdr_vco_reset: string  := "false";
        set_cdr_vco_speed: vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi1);
        set_cdr_vco_speed_fix: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        set_cdr_vco_speed_pciegen3: string  := "cdr_vco_max_speedbin_pciegen3";
        side            : string  := "side_unknown";
        silicon_rev     : string  := "20nm5es";
        sup_mode        : string  := "user_mode";
        top_or_bottom   : string  := "tb_unknown";
        tx_pll_prot_mode: string  := "txpll_unused";
        txpll_hclk_driver_enable: string  := "false";
        uc_cru_rstb     : string  := "cdr_lf_reset_off";
        uc_ro_cal       : string  := "uc_ro_cal_off";
        uc_ro_cal_status: string  := "uc_ro_cal_notdone";
        vco_freq        : string  := "0 hz";
        vco_overrange_voltage: string  := "vco_overrange_off";
        vco_underrange_voltage: string  := "vco_underange_off"
    );
    port(
        avmmaddress     : in     vl_logic_vector(8 downto 0);
        avmmclk         : in     vl_logic;
        avmmread        : in     vl_logic;
        avmmrstn        : in     vl_logic;
        avmmwrite       : in     vl_logic;
        avmmwritedata   : in     vl_logic_vector(7 downto 0);
        adapt_en        : in     vl_logic;
        atbsel          : in     vl_logic_vector(62 downto 0);
        clk0_bbpd       : in     vl_logic;
        clk180_bbpd     : in     vl_logic;
        clk270_bbpd     : in     vl_logic;
        clk90_bbpd      : in     vl_logic;
        deven           : in     vl_logic;
        devenb          : in     vl_logic;
        dfe_test        : in     vl_logic;
        dodd            : in     vl_logic;
        doddb           : in     vl_logic;
        e270            : in     vl_logic;
        e270b           : in     vl_logic;
        e90             : in     vl_logic;
        e90b            : in     vl_logic;
        early_eios      : in     vl_logic;
        error_even      : in     vl_logic;
        error_evenb     : in     vl_logic;
        error_odd       : in     vl_logic;
        error_oddb      : in     vl_logic;
        fpll_test0      : in     vl_logic;
        fpll_test1      : in     vl_logic;
        iqtxrxclk       : in     vl_logic_vector(5 downto 0);
        ltd_b           : in     vl_logic;
        ltr             : in     vl_logic;
        odi_clk         : in     vl_logic;
        odi_clkb        : in     vl_logic;
        pcie_sw_ret     : in     vl_logic_vector(1 downto 0);
        ppm_lock        : in     vl_logic;
        refclk          : in     vl_logic;
        rst_n           : in     vl_logic;
        rx_deser_pclk_test: in     vl_logic;
        rx_lpbkn        : in     vl_logic;
        rx_lpbkp        : in     vl_logic;
        rxp             : in     vl_logic;
        sd              : in     vl_logic;
        tx_ser_pclk_test: in     vl_logic;
        avmmreaddata    : out    vl_logic_vector(7 downto 0);
        blockselect     : out    vl_logic;
        cdr_cnt_done    : out    vl_logic;
        cdr_lpbkdp      : out    vl_logic;
        cdr_lpbkp       : out    vl_logic;
        cdr_refclk_cal_out: out    vl_logic_vector(11 downto 0);
        cdr_vco_cal_out : out    vl_logic_vector(11 downto 0);
        clk0_des        : out    vl_logic;
        clk0_odi        : out    vl_logic;
        clk0_pd         : out    vl_logic;
        clk0_pfd        : out    vl_logic;
        clk180_des      : out    vl_logic;
        clk180_odi      : out    vl_logic;
        clk180_pd       : out    vl_logic;
        clk180_pfd      : out    vl_logic;
        clk270_des      : out    vl_logic;
        clk270_odi      : out    vl_logic;
        clk270_pd       : out    vl_logic;
        clk90_des       : out    vl_logic;
        clk90_odi       : out    vl_logic;
        clk90_pd        : out    vl_logic;
        clklow          : out    vl_logic;
        deven_des       : out    vl_logic;
        devenb_des      : out    vl_logic;
        dodd_des        : out    vl_logic;
        doddb_des       : out    vl_logic;
        error_even_des  : out    vl_logic;
        error_evenb_des : out    vl_logic;
        error_odd_des   : out    vl_logic;
        error_oddb_des  : out    vl_logic;
        fref            : out    vl_logic;
        lock2ref        : out    vl_logic;
        overrange       : out    vl_logic;
        pfdmode_lock    : out    vl_logic;
        rlpbkdn         : out    vl_logic;
        rlpbkdp         : out    vl_logic;
        rlpbkn          : out    vl_logic;
        rlpbkp          : out    vl_logic;
        rx_signal_ok    : out    vl_logic;
        rxpll_lock      : out    vl_logic;
        tx_rlpbk        : out    vl_logic;
        underrange      : out    vl_logic;
        von_lp          : out    vl_logic;
        vop_lp          : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of enable_debug_info : constant is 1;
    attribute mti_svvh_generic_type of analog_mode : constant is 1;
    attribute mti_svvh_generic_type of atb_select_control : constant is 1;
    attribute mti_svvh_generic_type of auto_reset_on : constant is 1;
    attribute mti_svvh_generic_type of bandwidth_range_high : constant is 1;
    attribute mti_svvh_generic_type of bandwidth_range_low : constant is 1;
    attribute mti_svvh_generic_type of bbpd_data_pattern_filter_select : constant is 1;
    attribute mti_svvh_generic_type of bw_sel : constant is 1;
    attribute mti_svvh_generic_type of cal_vco_count_length : constant is 1;
    attribute mti_svvh_generic_type of cdr_odi_select : constant is 1;
    attribute mti_svvh_generic_type of cdr_phaselock_mode : constant is 1;
    attribute mti_svvh_generic_type of cdr_powerdown_mode : constant is 1;
    attribute mti_svvh_generic_type of cgb_div : constant is 1;
    attribute mti_svvh_generic_type of chgpmp_current_dn_pd : constant is 1;
    attribute mti_svvh_generic_type of chgpmp_current_dn_trim : constant is 1;
    attribute mti_svvh_generic_type of chgpmp_current_pd : constant is 1;
    attribute mti_svvh_generic_type of chgpmp_current_pfd : constant is 1;
    attribute mti_svvh_generic_type of chgpmp_current_up_pd : constant is 1;
    attribute mti_svvh_generic_type of chgpmp_current_up_trim : constant is 1;
    attribute mti_svvh_generic_type of chgpmp_dn_pd_trim_double : constant is 1;
    attribute mti_svvh_generic_type of chgpmp_replicate : constant is 1;
    attribute mti_svvh_generic_type of chgpmp_testmode : constant is 1;
    attribute mti_svvh_generic_type of chgpmp_up_pd_trim_double : constant is 1;
    attribute mti_svvh_generic_type of chgpmp_vccreg : constant is 1;
    attribute mti_svvh_generic_type of clklow_mux_select : constant is 1;
    attribute mti_svvh_generic_type of datarate : constant is 1;
    attribute mti_svvh_generic_type of diag_loopback_enable : constant is 1;
    attribute mti_svvh_generic_type of disable_up_dn : constant is 1;
    attribute mti_svvh_generic_type of enable_idle_rx_channel_support : constant is 1;
    attribute mti_svvh_generic_type of f_max_cmu_out_freq : constant is 1;
    attribute mti_svvh_generic_type of f_max_m_counter : constant is 1;
    attribute mti_svvh_generic_type of f_max_pfd : constant is 1;
    attribute mti_svvh_generic_type of f_max_ref : constant is 1;
    attribute mti_svvh_generic_type of f_max_vco : constant is 1;
    attribute mti_svvh_generic_type of f_min_gt_channel : constant is 1;
    attribute mti_svvh_generic_type of f_min_pfd : constant is 1;
    attribute mti_svvh_generic_type of f_min_ref : constant is 1;
    attribute mti_svvh_generic_type of f_min_vco : constant is 1;
    attribute mti_svvh_generic_type of fb_select : constant is 1;
    attribute mti_svvh_generic_type of fref_clklow_div : constant is 1;
    attribute mti_svvh_generic_type of fref_mux_select : constant is 1;
    attribute mti_svvh_generic_type of gpon_lck2ref_control : constant is 1;
    attribute mti_svvh_generic_type of initial_settings : constant is 1;
    attribute mti_svvh_generic_type of iqclk_mux_sel : constant is 1;
    attribute mti_svvh_generic_type of is_cascaded_pll : constant is 1;
    attribute mti_svvh_generic_type of lck2ref_delay_control : constant is 1;
    attribute mti_svvh_generic_type of lf_resistor_pd : constant is 1;
    attribute mti_svvh_generic_type of lf_resistor_pfd : constant is 1;
    attribute mti_svvh_generic_type of lf_ripple_cap : constant is 1;
    attribute mti_svvh_generic_type of loop_filter_bias_select : constant is 1;
    attribute mti_svvh_generic_type of loopback_mode : constant is 1;
    attribute mti_svvh_generic_type of lpd_counter : constant is 1;
    attribute mti_svvh_generic_type of lpfd_counter : constant is 1;
    attribute mti_svvh_generic_type of ltd_ltr_micro_controller_select : constant is 1;
    attribute mti_svvh_generic_type of m_counter : constant is 1;
    attribute mti_svvh_generic_type of n_counter : constant is 1;
    attribute mti_svvh_generic_type of n_counter_scratch : constant is 1;
    attribute mti_svvh_generic_type of optimal : constant is 1;
    attribute mti_svvh_generic_type of output_clock_frequency : constant is 1;
    attribute mti_svvh_generic_type of pcie_gen : constant is 1;
    attribute mti_svvh_generic_type of pd_fastlock_mode : constant is 1;
    attribute mti_svvh_generic_type of pd_l_counter : constant is 1;
    attribute mti_svvh_generic_type of pfd_l_counter : constant is 1;
    attribute mti_svvh_generic_type of pm_speed_grade : constant is 1;
    attribute mti_svvh_generic_type of pma_width : constant is 1;
    attribute mti_svvh_generic_type of position : constant is 1;
    attribute mti_svvh_generic_type of power_mode : constant is 1;
    attribute mti_svvh_generic_type of primary_use : constant is 1;
    attribute mti_svvh_generic_type of prot_mode : constant is 1;
    attribute mti_svvh_generic_type of reference_clock_frequency : constant is 1;
    attribute mti_svvh_generic_type of requires_gt_capable_channel : constant is 1;
    attribute mti_svvh_generic_type of reverse_serial_loopback : constant is 1;
    attribute mti_svvh_generic_type of set_cdr_input_freq_range : constant is 1;
    attribute mti_svvh_generic_type of set_cdr_v2i_enable : constant is 1;
    attribute mti_svvh_generic_type of set_cdr_vco_reset : constant is 1;
    attribute mti_svvh_generic_type of set_cdr_vco_speed : constant is 1;
    attribute mti_svvh_generic_type of set_cdr_vco_speed_fix : constant is 1;
    attribute mti_svvh_generic_type of set_cdr_vco_speed_pciegen3 : constant is 1;
    attribute mti_svvh_generic_type of side : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
    attribute mti_svvh_generic_type of sup_mode : constant is 1;
    attribute mti_svvh_generic_type of top_or_bottom : constant is 1;
    attribute mti_svvh_generic_type of tx_pll_prot_mode : constant is 1;
    attribute mti_svvh_generic_type of txpll_hclk_driver_enable : constant is 1;
    attribute mti_svvh_generic_type of uc_cru_rstb : constant is 1;
    attribute mti_svvh_generic_type of uc_ro_cal : constant is 1;
    attribute mti_svvh_generic_type of uc_ro_cal_status : constant is 1;
    attribute mti_svvh_generic_type of vco_freq : constant is 1;
    attribute mti_svvh_generic_type of vco_overrange_voltage : constant is 1;
    attribute mti_svvh_generic_type of vco_underrange_voltage : constant is 1;
end twentynm_hssi_pma_channel_pll;
