`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8NRCOAEQE7RCMEfucl5gcOgfX+n2BkOhbKBa4Xt81BtKwndWEfb4CoWc7T99xtos
jVTdSmcq9HIkqGrtiAV/7PZOy5+ElOHl51PFVyjiHqZUAMgqgWYk3pJEUXoYbj/w
3CyIL8U8qqKmFDIHAom4+go02wJxZlFKg9ILIgden3cqb/ClOc8LhCFsqrt7M7uT
mmBRUW+Xudf8KVOarRKu1sZYX7t2y8qHu9dNWasfqJDqnSCaWXcgAshbZtNjZ31/
iCcJSMzbuK5kA7WdbfBSRxfa28fwqJL8e7H64udFcVvSa3cJ3nJdfnuL1A2T+vkq
3Oi8A6pbkAZJS+eoVQMmEnIG9dMK8JroMX3ADA4HWVcFw7mULvQ8zN4SbZovzNj4
6KHAhmG8bGpsxwk+Kev7IjKD1qdrhFvfLGbCoFT3UqB+0g5apJelBXRVVLeoNxlD
jTttH4YNipqNKkoZQwZ55jAObJfWERSzYtL9q1ezxG7qVYooIPswChCyFIpP5Txx
JYW5e801NHeeOLX5LDESbQgJS+mqg3MY82XiUuU/WobAwwdJbZgoCEg2lh15klxL
QBCIkw2MaJUn6/kDiwqJj0tYQLC594OiJX9a4AsZm5F65BuXC0yv5PIEftJCd5nB
IjFV+yq8ZnRLXQKDFwkiJSqjwcLQuimcJmfhlj34off5YRaskvv6DWUUnm7sMvuA
9GFclvfwy1fK0akVRLznfz/IQ19uuskb0I8ySH34HPDA/qhHHa/uFvsxpqo3sVsp
g4HWv/bQ56kTI7qx/DUpCU9NxSYMnIJR+E75tWfo2ik4hyPKiwMR+5bpAjn6nbyL
ltC/EKhNffvpmej1lH9YIFgV7s2mL7IihUXDu2J5xqXJjW2FrKp4qxt4a7stUnlK
HorQyP/qOBIvMNjQIONjgrrII+NSCtCHD24T9istNXUDkvmWcqEFQw9cPi8/Ukup
cnKTY5EPuq7BoN/sPOzMzidCHNZ1/JnniI4acSvMGKisbjQD+WCrunatc5KDi2vA
RkzcV8KBf82i2KX87492eNlcIQCY7N6oXCyzHD7MimVdjKujFeNUvajEVA5bpCEP
bUk1fyFPs/YA4sP27AjKHtQsEhmACG0gAn8MFCqpaaUJurp819zwbDD58FfY5B4o
IgDuDdQXYDatlavQpkNoS3f4tjmsQCxTEUw0rkUzVt+lJKn+iSvXF15y23FGwicz
DrhcB83fyqMRWzEbt1gwqpMoMnc5omWX6nyHNpRrdymHP6B6dkaoo4Gp78HvCYUc
FJWGBUS6dsQdVUOdcTgFmA5k2ShH/iL8Pggi2AxKIDKMGrDQ1u3F3iipAVHjpSy0
OcpDmICfRVqZF3lfyxc+XoActlQQKZ71PkRRbSKNF605j1x+iW3arpu8Mdljp7+K
LeYboWdSAej7UGeZ0Rc5hAb7CPlaET/t9I5S/Ms6jU+mYXlmdFjIJmS/OHMd3NTk
ApqsoooQM4Uw1RIXcgvc2RzjkRUAqJj9c/RTh2zU4mXqR4vu1lYxaYNRbFdv4cUq
vBYn9KqW0An7WkVNsnpimveTvUTyswqujQ/vSyF475sDqFdvHO8j+eFKJAYGI7kl
Q8q8LWVNR6gjM4fTcR1Rj8OFIkf8XtY/5jzQX9hqkpZWQCvKPLhx7Hs1gHDbzti2
UwyRznrGIpdBPFRlZYsRmFsnU1dGXhx/wb/J/bqzUjhGPzLQPe21DHeUuVnKqLG1
0dv2HrB+hTrfRrkyX/OQSPitIP3rL4G9HIu+9wEsWWgdQhwKAI/0dAUBqueC6ikX
72T8JGgULCZyany/mp37GbwkicALK72WjTyx15I6XGoenHvEb4nG6UirMmRMyAGq
U3CxBmHeIjBuEGZIyPKE4GelhMHwJXBYY2wjA4/jbBPtqLYaqH7FCyNXysrIkCy4
e2C3cp+JKoQM0EUuqfifFzV+XBmbXYBXwxq+zelCbrgxuJ2Hg3n6Yv7GOgm3Zt/F
rz7mRmclEWoaY9TwGwsSLXu2446RcGnkdS+1M0G5OHkFHSYM/44FEpSk1SJwsFUs
cL1fnvg7F3pXYAInNGybcsCX1f7kakXF5Rn3ay1lmnNI4KIV5zjj2m8+TT5Ih+av
YxpzVdqy7eDfsVBlrfa8F/+hf4LxTub9i0lslp+PyyHNt7bKyK6e9eXjQZv5gszn
wLucV1EKY62XiafTBCHp2N/6Fq9CREimcUw5RwD2TOebP3MvhBv46GiwwhEYFAlC
HuEdwK9gK4FIZzFlMnwFNLo8NzxUCZNDyXQ+h+HTmxagNyRucSf99vWmQz5OpXB6
ZNvuqWaRV5zkoQoMvbE9Zafa3aaJ5YWKb0eSHqvIkkhq5eDIY5ZRyoukA5um16g0
WxHy7WuiTaWbGT5KKmDXKQorSsmXAwovzQIHXBXCd9fZiBEkS9l4MJolLIuyeoa2
/+g2KxVWAy2YdBFdEANpdKX8IvDie+i6DVlCf6KIY25pzLt4szCA9AzlRq07Y6na
dEGU7/SD42K3/eQAHU3nRVvMBJ3zz762qdyJU422hoBnDsQeMdxkIsRuw57xIY8f
8o2KUh5n023a/VMwNWVGfB8rQ+fMmf7EgdtlsmQMcuIhZAkNTXaB0z5Wjbx/Qe5n
iRNqZ4Oo180ZW/F2f9LF0mS+EYmtWiOtIcy9+gMbqp76CZL7nqajrwe7s41J39yn
DRhCoYYxjMv7p3ewFfjT0sXkL1NU9aQv4Es/wlYeHAxLpcPwsD8SP9XPLMtbA+Sv
gCB9LEq8oXWh0HkUQfIF2BCbgADpkD7x27iJGxYdeooTKe99X8Lml1WSK2s9oG8m
o3JuawfazEml3m+dVqqoFq/sEdHYDGn3yDniTAzcdfoMQzK+fHeMWKQLGrCDYnz8
oQRc9eCv7jN8H4Ce5YeTnvcTNdKA5vS90bcZnuyr4AODNNyZokxbLhjVpwwsr4Jm
PK/AQ8+eaYTxoIQIamV6UQJAtb1B8Jd4Muhv+6fdQcRuW83h+j4+bhceghw8GxqK
Rtw3MO+ylEGK8WcBDAc7UJEnqFQdGTw5wh6o8Vz96oqr2HM98/RGbiLA0fl7Rmsl
3UXF4mjoZ1gK2Yd/7fyuTfMTuYpQb9bnHQ+k8dLCuqiAzDeaaWiBZn9c6aP+Sb26
oXRgXdSRP8GDOVu98HSQ0ax5pwLcne4HhTPM6wL76/lsiHB2RSBACmVJFq6aOITo
rkuw+UxUiOsVkvvL+QIFsLs/KvboPN+wnKKPrF5dRk5mce4vW/gops+nBm/JhqaR
fHfl8y8oGfLdm0/ivO1hlW4tOVvL3akxSazdIHpwqvu28SwprOsRDvmE4PBC+tA6
ZVYxkNoKR0uhUxAlF5GVGOJxRUEoufUDae+oH1e0zUa1xrC2jrBH8X57AHrRMTMj
HC8Y/H3CEAi//XEifgE3YG+J9v1a2kAWk5Y/bhBko0LEL+Ec554PvJWY0y80jRh3
sqHoHu64nTxWW7RYEQRhCNraWVCwD7pMOtmQ/tOEtiNMskk1WyTm6VEzb4WOb9SY
sM5BZS++GOuPIb/9doHbjaxLVOzso3QIpbwH9uKdT15VbLqFhXmqXe6A8fROZpxv
TWgVMUvV/egv7csEc53W5Zpdf70rfB7JrBFAX7akHnnLBMUObalRF34wmZdh52XI
gvKhJZX71FdvVgV/E2eJ/1KLjuzKoGoG70UpBf4AKnwOBfLV8tYEElKWHnbm8Zrc
Xldg27qe5YE41Y4/SI74IQozIksUpEn4j82Qn6xqrBNQCbUGq1Vsh240vfTJmHJd
GXR+58upWzXzed+oljH2Da3b0OaqXRwB2LhBBEdkIOmNdXPBfWPh5yuwAsKeFxDh
SsGF8NQ7rwAce9PPS5H32keLN+FtHEURdhteDwpT4qpSO4rItuPKzpVNhUA/GtWb
fBHlo6VNYUYVQ/oerKg02saSrHN3hkrUtfNKt4GUxYdxLmF7vas7rcdjlx8yngCZ
MKggEqQscLzGUSd74Jm06hN6zlGoTgd6Cbn/ooBVhTrpXiZCZLzigrQnC2Y2luvW
A2ZjHBI72mlY9L1rw7GVrr1JNGfHtKIZYNoBLZ48NE5WjzwqjvxHnnFxfIgDnCdY
SSSBhX7MJMdKSHyP7W6oGDLyTFwyNWSj9Ukb9Badc0GrQWdWIFPeISOzQo8TwZ1y
lHML7rqrK6Wucal5QubXG2sbuVGBX3Oxk9ed7slOT1jxG5XLzG5f8746YD5WSb7z
OigfyOgehVPKCpNdvbRey5yFh9524pFyPw1zXHRtL/zXn4pB42twmPiGUo5B0n7p
jNWbESen9Dw0SrXqEpzEPkGWFnijXL2K1QJDuMSfVrn1meYHn8M/+dsqhU2mP3zH
sKGzRxQ+5QBodyCBdE9YApZF+EtT9SXXtdmpmijWJACM6JPAS3OEjnbGsD4xYIHG
+9oJLyheegx1IZ13t0dkRGyAthS1spYNWgwbdEDLtAAjnwAEEplV3/kYX56uzyug
3+dC7KRoB3WGbZHZ4r3sfUiZjHbJ4rErFS7HfHbRdVJjRW2FwfdlAiuPB5w4n6Lc
jekhje4I2LR6ryb4hZNkp5ZXXcXf7Cu+/CySspAK8Ys5j6gaLbaYPaW7v6DVTfqj
g3AovLszPm5U/M+S6J9cmr7Vd/DXCZDf1QATPEY95mDfAysYhmd2jF1iU1BQZVsR
pnALxEn6+5oZxu+eqolOn+1WK5l5C3SzeHpyXOY5m2o8ENlcHTsW5zGLO5SK26nG
6L1r2TlomtTk2ytFiHUsCNJqIDyMyRNdpKG90LXlVUu8Z1Xau76t/PnA5sVv+RCV
ZmWVoKq52BfrN6OTTZVbRmDTS5AeIczPntDNMvSKbnY1VxN2mOvu5BZ4OehS4svx
AlRHChNK1G/SNMWxsBWIpH6e67zsZv7dXd/9cZDSUwEMHWnzLIu1gHWhkYu2DZP5
VlEtl8xNh2FBGhkr1X3faWUcVQA6wo6ri2TCw01CvIAFOwuuNaq3rLjnsrP8jhzl
sfneJa1/Vm9tUv1jhNbDit7K0w1AShcRzH8jiDLcxG4ue0gCuoMsEJvDnfjxe3LP
QfKRP8dPnpHYU8FmFmUOHjBz1JD7ciezJg0Ywg13NfEKGTBiX9jmzEId0yUjh9Rm
UP8kzr3whyXlLD4UmCVvhRPBbnDFBaglgQSBvaAB6eMpMI5okzGf7s9rzhPt+eNl
woPHbWBivhsfsSAat7AWNTR+Ca/omBkI8DMNjzO5WhX4v1FDDRy8jmge7X3Fh0xw
UKY47J5R9eGzMeeeUqqV5ny14zi0cioAv1ILFfSEAwutEjuFT2HUmTpcyIy0aqi1
Fj7CA4Dg06kT6Q7G7H21Yv7/i3r/wOlnRdts+yA2YpgDD7R2stemhorVkIlBKM2Q
vCuSB0nMwCOV+nPpOQCbd+TlI11vCIhyh1mN2WHdtY6KyN8J/Cvjs6aiRaUvGTu0
DebedKGkp0Ngg/18GOXY57tUOM46SH1xWIldArnhpB6oHIalfhpfq3ITi+gYLaI3
wDwQ4mF4ckNXO1tGCZU4Iy4qWIFmQ7kA5ajBEU193YirPb7l+/G/uKAZM0crt4fU
rjkt8bHBDpFThxLAgTKzZRV716/sMv6Ua2fCyQmktXRJRR3JUEjdvc1DE8ZnXtZI
ZGo1LRP35z0WECEAnOn5S0PEUxW2XLh37aXm6cV/+KKE2Tr/tjFPgbM0NXmHn6Cc
3CXeq+LLncdEX5/6H1q2Nlr85fi6/9SK9oW4vkbLB6xCTfuRqQ6iGYOIhbeJYNUT
dpzKK0WU9ezyHtxF18DQw5kqpxUG3AvT0jMNb4jMsxrxuXsvn12+vck3+iX65pB+
MVWS3z51Y/DJQoGP4XgdpwBHOhFctX0y/wuGPBszUO9/gkvJwX2QZt1Mbp4RvWzD
7rDkb6m363FNY6rZsJLS9OKZGbjnbXi4cNngqf2gi8taBBj/3OD89lUNrbot+A53
DLm5TyvbYsbuokkxHrIASETONT9TTrwTsK7M7FC+kppyWxECr548TzbRH6WM68t5
FtUiCsqmblwSTk91ZFZuRY67oC+TD/gRgNLupQpRTjJqTD1EFR2w9HSODAiZ9XkP
eaSUZfOZLTXJJ3Rw6ayN/PJthI3srxhJsMG85Z1TckfThi4jDJ/dbSifUo51AYzb
9EtRm/e1Psk8taPCTd4tj4q/fMnFh0BwPp5PTujsc4WK6fWNIT4UgrddZ7ZCubRE
ajmi9iTF9cuQHvzLzvCALKOGzor1tXw8p4U0ZDB7Us+XzYma60FCqHIN09cKhCB8
b+FR0/M01/6aMGuPfTmeYmsH+y6z27TFRGEPH+9lmdrBvSJngDJHbs3KSqdkc9pe
7MIs0mhuZblHAfpdR0fHVP36Xvnt1WteolIFdHnixjcn3mEGV2qtCbH3wT05CN7R
KLI9FtOe1zp2hNX5kZ4//9HDf/zhCySrylKuE1/Nkj4QPjPRuTlRQwO7JG9uVaSb
eQ63XZH75nMPE37eISYQ1wCNcJANtKqPOx4hrVnPtJKlysw/pUV1dFrIJfl9ADE0
xcFZ0cG/aV7j5zNSBqaS+Hr/0tl8dECmY9fwWIbOamia/+gRuz/6FSCqfB/gGVDC
lijbXmDBbCFRXZy/WIaEYMnfX2qVpOUpruX/HlXKvU+yOZSILi98Dd/8uUUxWkGk
RtqB5YVzERi0b7y+VakuP614BlykRaH1TATSkDFBgxUUq/v2re3oFc2JcGrY+vKN
TKQNoBuoKH1V23DhHiQzgi9gKS2L/jFcHhD6cTIblGkNyOX20UemcZFuPXQyVy3N
o3zA51vg2mQnZ05jmNh9+Q9w1muhoBn3r9MJ4Lt+VHe+ye3Mkphcy4jcBr6bMC/3
yH5xIviSYqc2/ZnKjngRkt1w8d2VBRN6UzK5Cibho03CENphmYtbniLH9dzMa1Af
mVvlysZoDTghCY1HAjoBrbzKzGPNzXrHcM7Z2It79+mOLYOMOtwJ9rjFMWfOps3Y
hBBMfUkEAqp+rq+yYopCQp/dLUNU1YLEXoGcj2BPowhyssUDjUnILLBUlS8fHNco
b133Qf7HUpu4D+GlfTvv/bDntxXdzTOzHA6VHr3u4A1QH9sYDsC5pddf+lRcgSUc
8J+8cWrYDljRpTZ4hQK/PmofY395yYqJPCHHPfeJBZBl/R2BuDuqgkeiy6rKZiir
VBEiY7N40pCAfB0bTB1BCZWHfeldtrK0IuOMSYDivqKtQscahkxkUPdNLlfAx4Vz
5ZnHEZviLPGGVakHM/yYYyfbJU5stdg5xS2L53TX5OvugjzhrwqBL0IoBwOmDPd9
qGFSmyKhaS75zQ6/BqcNoXKBiZ040u50hYXgv8cVuJUhrP007wuOHyQ9tX6A46dV
wgEX+YFjXAbLc5WaGQgDJfiOOFT52sIU+BIqFqwMIBoBZB4dq/H5Ayv3TW7xsCEZ
XsEl/OYTpILgfApw06gWcCTNhWpA42OmfY1Xvwy1IrNexoAHUt/NcRDLpi137Etv
B4WVPZEhCLdn1tJSPlHYkdmDbTdiuN/LMXuT0v/G8ZnIdJDImeAJ1OXm0xC7Xe4C
/Yiq3AqFtSrqMd8/+s3mn4T5sn5B1I1E6jV6bvjxPhX4dWQ4wc7vR0V83doElCdH
zJUzx3J0h9rchviYbdVI9TMmlKDQXhmtFtkMAIcF7OtHSEtsBg+y211hkeYJewLz
WeHaDG5622efGUQwOUFgX5qXnwufwrnfMf+oW8UAK65m2OmJjEiZqN21h1gUEi65
9tttcAbiMZjr6Rk+SrVtoBdjml9HoHqs0SnR14ngdBLPoUrhIJaE3CPuWZ+Tjgf1
JE2AkPyVDADpH5a/IUSwGxKOlN8cVziAjEryC9cvdHvcA0ywZGSLn66yPaCtB6rs
s+dWi1Rqo3hA1nVu/4346UX0buXm/JEdC5fAFP/oJwZUa8ZBittSmlOEdgEkJGjD
69cv2e+ulDeN5gjt/Xx9HRVx1GoL/KEchRgbE4XSBu2TcGFU/41VVxxqZQnQS5uk
gytG7CAXAp29adnso1/H0SUCNdeQUDF6lbvIS+1bb0NOTcEZenKaRX1m3P9vP8dE
4TUU8xGl8Mh5UYoDBzbxPHrjIVkSNRB+gJ/kZuTiZlVaQ5xcMJqj8jkRpNhzcU7l
b1tJfnAmgtthhhll3OpkQhBS6lmspoIZ+PsLRM85rRBq/pp83p1Q1opGapA/OEjU
+gLorKU4S14ALn543J5u5s+EHo7enVtv3fQdcTANNj4U1o6N9ejm77eDTfhqEjZU
SDoJGHHarR2bnA0xAJ3E1T7G+Y6ELi/GhCiploxn9PhtI3WKJXPCFmTemCBnuJcv
tohUfJDY3ALfGd0nkoZwzbUAa8ar4Plz+KUEH0qk/YYnA6J/dqyrhJyoxtfXOiab
bZa1RYSNtYfjP29nlUMfbmhIwPBtonPrHyI+xzZsquywP8xveuH+pxGsvrQ8UYkV
wGlNjXLEtt5EqfvgLGxE727DNJ4gOrRWVOn0k88yRANTKs6OggHRFuPoLK+t+1i7
fDCr16DpUBDnLV/Zom6LfucO0HNbEexYJYWqyZ25zLtf1R5+bCdGH5VqHF1/p0sz
u+RmmbsIDyQEWPiptWyCHHGB/fafN2jNreC+RrdnlCYNKKuzQVUpMdsrYaMeoj27
ppr22xTn+PsG0EZdpEfgewG8yKKjX1mYwvRCQiOy+5qhtVKKAxDNiOPboQA0M3W5
KefYgFpiouBhgD2Y7NCY68vcBz9mJokFywoixeCsHzI4RlxrNdIK3Ye+y1vlT3ie
WbR5V9CM/2Le+LTz855C/cO6GVj9UUYdjDCxHxCn2WRMGpEBtf7a5S58INBEEgTg
HMJbJH6/uQdMTrjhXC8ST6uDKHV6gmeeXs6XtBus/u3heT2dMnmTwGpentko7dv5
bFEt29OwRHfYA5dBYYZjcuhzPjV1b46qfVEmixQEB6e9nAXPaBYo3L+Dgbe8504Y
aQmXOLM2hvXl9rBjl83MMc6tAcGvVVBcUcrPUGok9sekvdF2FbWS396k7NEKrxlo
UBVNV06hwEqCy5OuaFdNE0R95UeGTMe+9JySbFJzjhG+ftBu8I7yeL+iURuFshrF
wVT1+FvBBxDdB/ZzKMfmnJX0JHTRPh9rZSU5TGylKWHi4LuonaGohEWRSr9W/E7w
v3VlaWZf2q15WBr9lij7m3A4gfJ4XIOO/kaFB3+SPotaA8g6LI0LFcvX2OPT2p0t
OtANbfRKwleil+BBaI0cIYZOgS0cmFAruj30/JLp2rDCEm6X+p3sSg1env0bB03N
ePKh1mtzOycGAfOrQfmanueX77RihbcRSPmE7xQHq8Jv7x7PCt1IehleiJcXGWpi
S0wONS85fVwoF25wI9U5XjzVs7VNlxzokeFhAsLRMQ73uLuyPyo2Vp0xyhiAQEb4
ITOq1t/7rwI/+PL5g7sj0fAdiHoTj6HTH3njADA+zjonztL+DrIhCNEvZsiV7NB7
ZPq5FzKw4KUZw7myeSlygxhs5UlL6GkPEGA4vCSh8ansvtYxlNMzwISC46u37Gr1
eDPcoDuEeCUeP1pK88WHZTxHvhT6qeigI2C1dLAGNgKtrTP+7ch9gX4u0sx1plzq
U0FS3Zf0BLxBnKyGhLannDKDtjZxrYXH1XGMHBlY1l3OwIxPs7Lir37mQJUMeGCx
x/O7crwEtMbqxSVPbTr/pVxBnfhqf7hUSgbosGuSMyL9jbvRbIgvbK5IyCsZonPt
h9EuaIbNeaZPXL8+lEPJzj1KFUC2akZsxIk+yWweEiFuCa9zH5nm1fFZsxntvSxG
WBJUYqXrQVYLziS66omTJSWvc0+2STKHrTwufB05BhPZKf3ftgETG+ipcwn5ag1p
eLTFBMPBwI1gmTRNlBETYX6k2BxeNwFnWFqYUMBCfInAn+Ho4kaGgtVeFsDrCiBx
Ux9P17ajbhekg6SFCMRyvsq0+ql3s2c03NFGPqvEGaV79IowmdeQSD4SVnFdY/fs
uwsp8RfHMdlXwbALyImOxHAunE7fQyebHojO1M6MbJn69s7zmzH5J3bCt9gMJ40P
0j3I+NiIIA/GSRYZWhKXcKvqVGthFX5+JXAgDC6cg64+BwnM8+P+cH8kYm+lHfrH
lIDpyIo3JQyQwVzMdnrv914QoeTbcu5bkiCyFhb2ro0gQcfikk4+uof4gv6NlKTX
AyWVpJbHlCr6pCrCSqwRAOLcEcBiPXuI23pWP6FBUIHK2vYkw3fwrAi28cad7WwP
e/goiB8IuBunPVQKkFjyQX37GbHp96TRSTopSzezyJsN4rsKgOU1gv1Ojqc/rpQS
r7IwZewzb/3un5c0JE181AG7xgw0kiQq0EywYkvnggBr03sN/m/SD4gaJEbDPayx
uLjAmgMNaTKu+xZP+Gwr+i/FEXiRprh3zaMOK/mFllswYoJTVlCADZe9xYA2cfLu
bzoorxjOMlK9dySBQnzTge7aavmltTwKnjH2DPN6uBisNooW2oxttVh2q4cKEDnx
RQmnzJqXtuFCfzQiicyk+Fy53iE81khBIvIh2k26hKiADkdwf8atYjidlRBhYZI5
zaXFPAS+wnwAnhb16TMBMNCQp6csIcE97AEGtKTXyF6TPxm41125NuFrnG/ZneD9
T1cVRRO8qEyComSHtLwG7r7JJFP1xJUTlSJsHUu5pXyULU1BjGb5/Y3wBR3Tfg4t
5DoZIFBXNKxG7CUwJafVWNvgJU9lxXi02sRxy6rmqTJLZsqSgG5gmqZetuQPQFqF
+d5o5pYIGSoS1gbNdPv3U0YBSzdKY3QdSRDBLv+Sarrj503xhltkAU5s7nCzDT/+
tGkV1sqqaJT5nx/kpWu0DJt2XjIcENnb9yUZG3bj0Puc4JSfE+30YZczJzB27XhP
wGdxONeZf4LodcY6RsIgD+ireRyrDj9kbRufSpmigeuIZd4MT1avLxJzEu8OH2in
MXFGHORuiJHItWhFs3h67VgbKVytNH0OVwTQi3V4msZYoWStlodNXhGwsvs/ELfl
4/z6CwrpBX48DNCmRqJSw55LE2IVxG2Kod6N7UOqn/tEcVwvJLh8VUspTor6kDxK
yRNJ12k7GIXs6WCAtHDoUCS88GAenoiwB56Kde4Vbp3ZS89YXQPDawh2H77dQ65f
MAK69jT66Ffxl8eR7/nFO5o7HBzrTpXXhulfZ9boshqIWds9q6xuxEsuk2JLSHVF
xwq6upawY0fyO3GKVynVpjYSzeh1aHvP+USDrJ24i175Hg1VYDtx77Ku3ZeuGnKW
+yHmwqEp+g37YVLiprQ63B3qKVd4FBnluIedpVbyZ74ZYdlUMDYCUvGhBEsdLNVJ
zcC6BDaTnoHsTweIVaPxMRpaNUBKRk8Ni14zc85Y/DAry2EJZxqTm79VCoGxcId5
X4njm40LG4OwhGVUMpimhgIYCzaeEXQF7fwkW2VIe8kScO9YbBm5IvtICpyhwUM4
YKbTrLxUsxXA0ll+vbgHoSPwEdAQ5jhmgf96HaAZuhzq4VYhgjUaeyRL31NCofIj
Ys4trct07NFARzZZbBD/ugCic32siFb96czR3BG9cjtfj3ecBqNbnRO/qwUA0Uhe
nrat7Afjcya0zPjGsoR5mlKDtBzHR9OpVQswyMUbW4nHeqpjaGPMCedVV58RaAic
pLDlr+0L8XKg6hwUf/I3udmg3f9RvikriG94pQiCnP1yB0SJVPlQ0t9WNiKOZyqS
VLuawZtFLaQm3MKUG5Xy4Us2a/q2qK7+fl8PcgVcT52liKaXmeuwsSN4mDqtaMC7
CHmdg6sOeTJrVrfHBwibLp8LyATuRMAb+XbtOr0a8L6GGj5TZaDXUIRneXqbSahs
yQFk0k8zc63S/9z4k69AXzz53bHjnKhlOPauLsYC3nEKhZwIdTj2GjmE5IlBrvys
lAutREeCvOH8hXqPOY6fvrdjH/sni8RVi4o0EYsza1hokjp9k2Tv1a0UaXRYWGcO
chI9g9fzGjz4hx0Jkaqyo0Ee/rD0lrSvh6FW1BcvVSYrbBbCkTkey0g6S2aG7Br1
Wx0kzEUqEc0pRDlc3/VrPlbiCysTU/4K1Z9CbZsMH6nHuxpuvfyQ5QFnhGzhTrWw
J/KrU6X8NUaQBlx4Kf0us7ePl88SAB5eM7NSczGUV6ZI+jwH6aK0COkvy+9G3jrY
fqbEREUROy6zfyoBXhivp1PAw3K/AzybaEp7nbwz53zS3WhfA/dmvZtQsS23K2yr
3aef8bN035Uuas+11iT7x7ALVw29e57EB2fdgthg3frQMWZw1A5+qhuGG4qiezvQ
x3NSnnz0MAjEVAOSeJ9b4O0t+MM/5Etsu+LxgDoP4L28aium8/9iyilLzxR+9SPZ
6rap5iL/uk4LVxTMYlX2hcfM5o6qlINmCxj9tX7YDGvfIY8Us8d4s/OYJ3WpUAyS
zmVeVAPZiEuZc8zpTC2SuM3Clkmq38XajAE2+LUGxEBmtE2BJzw6G/qx4xIKre+C
YemMqYN3/PTScz4xHqnf3Ns/uNgDdp4ZlCHVFC4XHYGnEV1iXpwWiAZx52NLJhdo
RFk0DHTEO3uhDYI9ZZIro27k+SMYLXvr8i8ot/O3wy0FAkP4iAlFN127CEED+i75
spNRkfSU2BqEqAGtzl6rHSfkvmvEC3lZYx0quwGg9rK59XimfB63yLxBLZRDbXDJ
9bXra4eEEf7MDLG1MyR51Gytx+73Pf9yq+tu75Jq8EnZmRohIYyUAGinJjDynqge
CXvIf4NfnSeI8bjyro6C8jSohEJnn1fIOmjZSbV2nibUppSiU14SfBEaVz0/Q2DE
EXLlG0QTHWum77zzjstvha3M8S7AeJzZvZjEQKcmb+j+EZUJKNKLVJYM0KlEKPVW
XQvofHiCH5QZQeBwoODMuG12r6juL8VV3w6BO90SxRzqnFUjqAMDg2VNmk0e6L7E
/0KensuM0Fx7KoAM+pNa5xfptasTFfoGNBFKWsTP12o9fMZMYJ1miWOeYQhkMPdj
E7fK5m+VfyJt+7BfJpXzjME9mV6gbMNkx7qOOUY2oPJPSirHSxFKf+A81sbxQg7X
QtZXBYUKLfuUS5mv4FgsTQGJ3iWi8TQ0Ja3Xh7lE03pi9IV3HBd+wxXCB68N8e8z
GLrA3hImmMOLrYvgGAaogfZMR5tVGFEKuDxKWBXSU8FMxbhi7Xs+gVa3+xvZ2tXX
Fmp+UHiAfz/HUU98Z5Yv3e0MeMQyxgJ3MZxb+nl8J2fxFKU2rqrGklO8gR6JHdDv
ajlmqaARFnYAT8ITToUZSjzQJNFh1kwef+/vJ/OWgYtalqfqQrEJWlbhWSepURo4
YpeqbcBgNc4UlQTyExb66V5VCR9LNBz0n5Am8ZstY59UN5/q8v0o57S8K8x/aGk+
CCX2jZdWwG4oWD4VCtlaLELgqWDgDgtl3X9JB7b7YjFr0Ch/E+tBuyCCoFPBBtl9
ZKV+YuKhnZ8juTvw7ztKZrhVbdV5fkT4mgkrxEEN3PkZ5Wapvei9yKJzSfWD+SxC
mUSHgl4iqctDK08dQe2UFhPEz8T1UzC4D0N40L+kBWKSnZYpO3qA33iIg42ZiRMg
zxHurHROpGproklAAoJdVbqLB0a2MyTjqq6aNjP/V5NrOX0yWUi1DdOKd+QAPtPK
OrCjb7qg57bXDR/XR3FLMfeigU6apbB6VOt84oZ5tO+vMDCo3UokA2lPTLIkLx4c
Wq/mgNCAcgxkfk2g4mDvZ5TfF2VPk8UOXGDxjADNesS8FOoOXqQAMDqmeTj3UN9T
HtwITkoGupIwEuNKHB48k1dmLzbpi3TNv7Mcc0yoO/GJZOk8pudTnqAzHw7O9mZY
bo0JUpQHgK24qCZniSJSi96MxXsBW55frj6KT/ChqX7gssusemYg6tm9KMzk/iD9
WqMhXFCc9jtA+pCd1Yxx5MOCFFaW3C0x+hLmV4mahPRQWqFiQLRI1rgyOif9ifRV
UtB6jflPiBAWcdM/pixj/wqRaoEmoPeAIZvI3OYOZ+uKzVvxGazR+HEt+c8ikPd2
ES+Ff4MA/o6RuimlB9Zgy3N9TKXEJ5Jl0TZSihs6uOAHV9iNdlV0A8tB0eDNEJ4+
R4NaGNTCbpEYuoHE008uGkdxMpD67VrwtgYZzPRGXsLekaeP6Gv3QCYw3TVz/bzk
zM+502AIHR/tdMVdKzROlBfTCEWFNdz8YkmVdZmUhsZoJzZUXbqNJVd1Gm/rYpVU
cp4EvRXZIOsys+Z8RLJUPWPS98++WD4+n6kvgD0M3Pzkiv4rW2TLx+XztN0lV2rv
+7Nme/gpPEUM3AsTmaP8WiBleTHPmEg1/5FvMm8ESUJkOdkC4Dmd5LMyeQS86W5i
LuBhxkqHQbrRrMWSzOIGDGUaIKS8g5g2bwnNR5JE4ARM/vWz+UIpURdgtVT5wSvN
xZu4ufEzA1J2vBoZfMQusppcK55gzsxJ1s84+sdj8eEH9Igs7AWJXiWaoOl9AJfL
STYZtla7ju3VdnSvTn4BT3swmt4gH2kriVdk01PN77vhGhClTPDuz3Iw+LPTYfVm
5XExwDHWyyLsnZ4/jZZ5rslRt6pIA7vsE6tijf+Xq6jCwTC964qzyJXAVIra0bio
cImaBNpu1N5yuCIutkNxinZLIT9dKBN6M82RRt+FzSkM050hwXk3nsU3YfnK7Rco
LQsHjwuo61DLeFiVH3CKqcdxtxYgI4ek6QC9YnmMXZuEmCxkkKa9BkpK2pC9GhK4
fSfObgklrKFjK4qF3wjTcBsq/8usODgy5CsnmZLEV6/BPe4VHN5scgnr4tJI4Tyl
vKNpE77ulmeS3UorcEcijKrAN3l1tVlIJ8bILtj6/BK2Msiuf3elbJskgvLom7k9
nA5wbtvKaWbqUrgHEAnnTnA93DtYxM/NAh60jK7GgVLvbIOK+UyMzSkvelkGCh3v
BUPxvrx2cjz22fGJYag0gsArcNT+plJHlPi5LQuQd0OHtT0PDarkjL9YSgXkgaom
hJ5FiqKRh4nYOuf8QKD2/hV4kQJFCiE/iqBvkPGObEmlaeKN5qoMkX0rIIe6A1By
zAoD9q7lN5MlOy5krDiP4YgVdurmsfzCoHesWXBApIudmeJ54xJ1Y9n9kWn/1PZV
ek3bof4FA6jusgqsh/rKqZScAtxSo6E9uQA+3k6a1HU+fy7YCYRKFSuQlyI+tioc
IqleZHQ5D8qaftTY7JCvVgpaXY1xtGeG/c+/qIb/pBAqQxeHYiqUPksPOsOnS+Fn
sdpYJq5SPORh3e8lAh9L0oruyo0zOnwBx5hbTzWFdgtYUdkw//1bI5iGWx4wgIDu
Xgg7Sy9RxDWvv3KQJMifFvq9mtO3fPtSo91+PaqYKJM4Uch7vgP5HVtr8Yq1VQoD
1OHMdqTAv4j2M4XPJxmVdIQSLHaTmpec3m+4If9r2WqYPqqGnGjXlFd5STaOh3ZC
iKb6jLiqHGvxyPVnEEf6ts3fYlM3K3qOOj4jLjpxITTKQC7ue64u0k0e1/c2lyr6
fHuBg+69O1ahvrB+YZ80MS6o2foWBd7eGtOOvRW6SQxdKAjPvn656F3gpM+0UGJS
n63/V81RQZGhTHfnQTMXsfxSo/vmTiHhbR8UWixWUvU9MhyH3MM3AsvonKiWm5sT
CQOdTRA+goHpaK+h730U1mJDcnDQj8yKq+O9XW39A/L+YL/jMEA0y0ZtWnLGHBlC
v2bg0S6DqXpbQxWL9RgQZmR7gHAR7WCPoEpA9qyKkj2FnGbrpvBlPPug28S+EsI4
tCCXhBeZbyOCMJoiT3/ZY5AOWoOnDlhV0S/JHJy6F5HvXbWLNw0M/3pFcXrVaMqs
pU+4/fE/11XwxnrryMSPD7wl3ZsIILmRYUElpBQ14E6Aj4ZUAewBw7WKkar+kO17
RJGNpIw1PivRyfgrKVGgRd+xJmTmgtNpRtqWfOXciHzy7aFTSLP80EtkjQJTCxVM
JrSVgvpTH7Itxep2dnVvaZO9FnL0aPUNGj5iG1mo1LO4n8P1MbIGCjIRf7IqUFMf
tkf5N4x/WZD1AIUTeabaFt0ooo+dHke0nzGCa+VUqqI0EaxtSYKF0ui89wzMTZPB
s4ryOcb53ZNVkZCvrxDT/Y69Y9zfbMPOMz9LAE1SWSna9nROvbtoWVZKhw03Uxhx
LXSi7KExMoj3teajM33lWOmaZmVfHlKxv3thw5hv9w06o71WhzeKB87tbxGX94Og
ETwTiD1kiWdKfPpE2a2FcAhzA2LtcLfMYUVKwS4/gYKPEGvIG6IKBGO4iEAXgbhp
rajXrtwSPq2btPsNMVNYsKimIDd+cdOYFU91AOVY1fvXQ2ysUryudYAUTthwmAd1
EwRb5eNIohlQ9GIRhKpmQ3yGVnh48VmLPVQyR6vOTGDYc+piW/8HTLQNy8XDCRcO
P5J0j4CG0Yb/tp+pMcVTkT664r4UV2RGMV8YVPGXo3p2s33wCUNgvXDr+0ReXoxP
MrFZIBYDp9eDsJyot/kemAOmL7GdbQkdvV29xUFcwOKAmTvQdent/5H7sPjN9L0G
a6xY4deakgG4mykdX8sWCpjpWBaDtqhFfbi1wpz4AP08rjis+oaI6W/ig4Sj9+hR
7sMWhQdMjDLaMKrcqfbBru8iID9wsU11S5LvH49MhLRnd5fGRG9/qfNdQkzLuTuB
h3diF6iEjeNaI/6+N3BI7V+ARgahqro3G2h2dObMq/SBF2YtnND9ux+F1hJ2lq0k
SKkpub/0pIsw7+g46rRGhC8kjYbizfuQDTyOOuAEEWcttyCP1r7Emh1QVkxHU5e5
Tpojh7F6f98aKYWALdj5ArkChqdduyLEp2o3Je7kF08EOHsDpazVKf3sAbxixBEL
DeGHldOzTrA1TGnxEgyxKFMtY8OVgj1TEyrou43+KaBmIMEtDwPL1XZiiVvs6fYO
6uMogfXAtfspf8b750uLVtAgWt3b41XkkYp6OqwgFezkcY3zH+uF11k87WUSh4/E
AdP3SrKtoQEyS9PszT2yQZfjAkGVyIcu1p777L9bEV0M+EDxhv1fdlitky9TSQ34
MPGIaFQ97O3vY23mPfxHKLQ/AkioFKSRJY9drnfZzO8eHg+GT5keJZpSjIxWTHfV
N5A8eK5zkmijKTDs4XUErWnh1EJK5dCE60m2/0+pojtXbCO3wmikqPpKdFUZ0iK/
qLkrWNqmGXCThHc2MXZ6sa3Pp2NJeTMQ/JgucRHn6KaA2dAQAzNOwGqQyNeO5y0W
WlGkx1rzlfg8JwT/SD9J5J18qzgzjuk/OK8Bd+qn1F0P341IRsEDYnhYsmOuHP6J
8zb35go6iXJDxmXmrj3dCz3wqzZjne0f09r3Hug/MxRO/ITWf34lafuspqUsmvyE
OK1LCzZ3W9DVE9OH23lTciV0kR2SFiDgau8K57RCo2JAbKKVP2cVY3DXnqNpPiAP
+sw7JGKgJZqHQnKwDLMDENjj4q/rt0qkOtk6iicDqeb4NsDUpofLwixfAFU4qTNM
WX21at08qFWwCgdl3b1N4c5HpgKzD2ZpZSPiOpuRv+DK5lnH92uIvR/Jg1BlbNbw
fOI0R0pWQtLH4yrBNhQnd3MY6w+dNMGo4qqxfExQMkbc01t0bdytFDSA0hEHh3k0
9IvxRRNDqxv2MQDGT1M/K11e6O5Dezu+lweWHAaSZ0HEn4JhoFR6w5JJ3g8ya4a+
W65Qk8vB7FIus7Fh84c748nEHcIzdIsd1ySIc+0vMikM2uSfuggwQAyHytyT/BMw
Ce+4PXRzcPv4eYLDX98mZ53bFrRNonVcjagQorC0e05w5LXJtVKvw6JPVpdLbbZZ
plONmrFO4899q/EIZMYm6SiRsRL5VXu1jhxfmu4FflIZUIbOqoCdBot1DUefiv3n
/l+/KP1SaQPelAJT9DuLDgTlyGrE/dyA8DTl0N9oqKtsSwDGW7euVbbvpA2TCrMY
//wZLvu+gZfb4+qc9cTS8q8pRSWocJKCLdrGz2q6hdrm6geIfA0yPKDrCfl7pCKI
23x1x4a1rMwM0uPi1rf/tu01LQKW42579BZ4hX+O9MzDDLWbl6DKhMZiyay9etGQ
0opwLnzQJOwhNCUNnq/u5yO21yZEkv9s1d0eC+08gIjY7cE5jp80Biy/yai59+uH
V7SDNyRZ3MHIMlnllUK4zytpwrSt4xZ8Oe3z9wxylHX/rxsTMYuAN4r4IE7FhFN7
rWkJlW/2lQHpT8Rbspzh3vTkvFjG8ON6U4Qzz53VmTNwKRr8qBqJNeSHFGGhskB+
YbFMZuRS9Ty4Dd+glrH0tkDG+Nz3nO5ZYS+iKhSTcYGs/EYUCAq2ZbkiV81qvyLk
ip5VlnjWRXLvpPTf0dA8q0pLrqRWF/2+koOjPHmTd/j5JqnVtUUKqEqjw94QcmC9
iNP7ForV+PBhVqXX6rdIDLL5PwZ8a2UkrThEFGABZcg1Ga+IMjYxfISmZGzRSL0F
LG7NCg0wDPs5UC1ZAWkJ31nOtrIayendxAzZctgWIQVtHMcsm3Ey1xbDUjjbaXjm
httIDnTT62EyTvd7ziYXWT1TpDRHrfeYJ3hBgCQM52hlWatFVdjgFV5PhtZ0B5Dz
sfzqOaQvi4K9OMveS5YQ0q81QGyUFZgI3+Woq/o94nWVPoXi+ExxDMsTmMlxtoWe
PGwzDhWs/QHkPlTJ8Zce2D/cp3UiyyAFFHc9PMbuvQcNDGXgRtYbkwdm/4+FXCHB
vAa4c6H8OgGDYqcqP+2qiQNMnCSblQbeUa8aBjqyjNsS8aPGMbzUGwt1A75gyOzl
ToR8+J8xo6oieUff2LMMAg7ddNyRfB44lxEs4BZEiKYBMmAMwC6abfivHZaG55wY
qYKPt37+nu984ubBxlnE+XDtja6rnzTwuim1XgVKr+25O5DH7N164iZaJ0eKC4eg
znqRYyzeOr9Smox6yu2ads2H49U8AI4Gg8o5oyuL7s7W4VqPXbfGNPppT8iBOY3X
weHG7n6+854zIPOddAJnpFITyG+AhQ8Rrw+8JlGgJNqK52ZtY9d5B54HyLSyEHuN
JrtI7ogLXIeYIQFKtHQGn43YUxImQ1wgXyHjiNXPDlRjlUMf5ir6vHn1Gpc4L9Ci
G+tEhG2rdQk8WS4NeAHfB8bWL1wI5f0NWywv6fcHsxFUH8FuqQA8PPkVpLn2MZlW
FWRx9Sy3k11cGqi3T8rB7s0SCDoFhNpCb/1WxbsTSQkeq+zAcAXPJphy2i6MUXN2
VBOeKrvSbE5SbkqbLmddTHNnz2t1vBSEvco5Feu1XkxHuvhGUOgeMevXDSJsxmIA
W/dtF7dQP5HsTnzAo3vL1kH5RSQ7dN0yvMXIxqLN8AnbjDgGW5lFGykmYdKCFAfF
Cm8wNSW9FSrcLRbta4BKTP8WAJF09I/jCKGcIZmS0J+bPpWC7+5z4S/yaKsWPtbK
+KQA2gWoXSucxShamYXrd+0XNMLoFmbij4ZVqwUU02/nFNY6cA/DyAaU1AxYQx8L
otwm80OE+QNieVic806bmf874z//JUh9v5c5dSSR5rYB46LUpF5n6iyWeYo4FBL5
owVQG6VkFrSD8XEtPKNcJjx3++ol5bOo817NKKEjesLNcuicFOkQJfe19YUVvoI0
PEawrDk7nN4NHsA/zvJvJisObHFmSXpQtUO25SXD7uMBL+Tz994LbEWyyh/Xe0Ne
UGXXuSRp6uC3zOa8jQGS0Di3BP3cTYbtN1qbKAgTyB/H3oF38hgzAgwO509B1VSF
9a7FfOmghcbJN1FUC8OQwp0U1mmu4bJBsmG3CkXsfggd5FjPdkAnKNwTAiGWHMuQ
zJfVjq/5fX4NxIcp3fygCwrw8R0zrIBH6WJkEywtpzqOn+wV+L8fAWPezhr/KlaU
zFZ2n2+ClzJ2sDgnEEHTC841ICTKGglVO474HAXxgLeRM+4eAeJJQfuZDm1kEd/v
0CTbhmTumc3AoupMukrY9G+bGmPIXaCYigIzsQSGh50/rtowDinz+dtvrLOOFTcm
u3WCelJQ2olI+6G+4aIZ/25h6nJYvxs4idGukRh6vzAVALUsy/c4lvz06T7Jj3l2
ii+3Ru595D7tmgWbjgJc2OVwSLmb0Ig5r5swuYNXvKQBZ3pkflUxjSkQwIt2g8YM
eXZ6woNDFOkime+1ZnyEpITFCZjB3b0mmBuhhuz2DbzlquxthGLatfTKOZ5XS7Pq
X7uCKQu8lfuKZ0bVw37t5GiF92/AXTdkC2xGkqUrzvsNJitJEmX8mjXF/6TTrGh/
dAuWPEfBYR348KPslu8FARUVrOn3FnOOV+hsLg3zJrgNLz35LqpqDB+w9fB4qk+6
qdbbwh6fu2qceNbCbvnezBe7uTo4JhiVBmR+MY8MyUJ3hcEcx77JJznyVHmCRJPh
zW0ZGk1UTGVjILh+AVtsnVIV+U0SgFeGzXpB5BOG130cTCRbNHkHOMWntoBk3P8F
Yi9rmQu5IwNbSOnKS/gbih8rCMHBBPlgNWseYdRpLk+dDq2xOQRPLjjGPRuIAtwz
WSzBceU2vLuBN9iqP3cP0UVDyPoHs0s/190TdgvT85euDWhmx+N2SXf1UTnCFZPb
isZe3Lo0GwN2f49VPzgkdKlOvtTfXkfGy0LVa5uXb544yyS5pVWxeNq3R3HX+xwn
LehwcvFl7I8nTW0edKnrivD9uho1mtHvzue7MAopkZw3/ypDwRc63r5Ys0ZSpI/e
8Bwu4opJqGy6vr1+F6f/DW+LjoWmLsE0GaSQEGYXOSfLb1G0KvZKQuqIFNpJO2/x
171GgsBKc9Pd3lSEFXSnIwxeCpLz7UOtIHk0xLQr/MgBM8vFu8GeSVAfJDnpgXfV
Q6VwF4H9ehca0DVQ5pEkmrxorcbMJiBvKrvEIAYcQtq8eLb+zZn3OncRTXlsIt1N
hMtTTLeDdzwvS8S6gu5lJJf3203nMMdiTyQF2/JD99viAEX0ZDAdPT/KyDQRwdTW
yrdf6nYtk9MzB4A92I+nxZY12Bm/9BOmT7zQVvrDBUDmKOkhkUVhL8JbIJ4SdoRb
NsaG1ako1cbvbkNVat2FHoPQb3DcTRkJ4GmzuqZK4y7LZZc1qerFyuzMGUUf/Vk0
d/Wcc+4XMtIaDHU8KoyXHpHfT+6GFangxNEeA+BgOwYJR53yI8dPywx9fVPYdYOB
yCnSzNJ8I98pr8ps7tVxax/mEl2ccpe/+2zu7uv9IfYRlck0UG1SJlgYx0DteKa6
WYlTNjgSTG6yeQkcjJ2s4TfXmu8T/qhvBqciCfISOtTWzh/NeVQBAynnmj2ccTzi
cxPuLVYJJt6OkUELSLnztcHSt59cSgjO8PRUagp/ocGMEcZ4SnWheb4gyVSIbd+i
vVYHgZOLi1De8ZuTFE+DkGrDV6q9K35EIYBEcgr+c4r/vrONmmLNDl6nR1ZPppXR
BY2mXZcNmkR7SKrgerD7RtXmwTD5Y+/qyZqc/azUQcDaUlzelQLPjIgA0uF2Fzl/
+6Ef8grZTQlDozDWJeLLoKjvAVmdt+Ow4cRg9fqpEkDM8Ob/7ldXz6PpM2DywRIu
b2REWwc6gbNWFdK9/m6uKrLjbht0+ZVrxOc2oMy8g3o6AGJ7tzTb1Ose0OR9EY/o
vxA37wMyOffBKp38/EVIMXs3p0jfg8P9aniUF3PQo2gO8lchlr2Ck5rEhjjox9Ak
lNGMgThLvvR21KhhMVDgtSyxYgbuaBK9JoqAiDjKja1wlZWL7F9qg04HVBo98Z9V
K5iFsWHcg8tVTAS7LijzTWz5YwnyhgQyEQzq63WFtroW69oYYWeqpbsoGWrbHC5n
10uf2OSIYOx9AiR4ZAeyRiKLYwNjdezNwaYuaYg2fl2r+e+Xi2xY7hbvk6LbXxir
ceAg5UZlOukAveZaJTd2ow8njqXAgfGbh0gK65J5qDhK25FtQbdK29zZo4wTAA65
7zdOWh4OD6QO0W5Ijgad9E3dkhH7aMvTYvs8FondwMA/9hktw/dVTh9D6GYsBN5e
ngAsMPFwJO0/tisOgF50lDmpa6LrJ5gfKNAcy88zZcwpLqS4pQKy9uGPLxIC2OoH
D/UcHJH43RKFQ4zjzWplGaYXh7DMdeqglqXUZcpgXkW/xVw2LbMZA+f2/8FF1KBF
3Uoe4M5DMq4eoPSrI+KPicOvZzTyNjnDjWo8ZU9Pyez1yZ5sGzT9Ulg8Q5TRW1r+
xSS7lF1EkctWjlEFO4a0G1WV7HhMY4aiaCspH/cZtF6JOweyeotjmewo7cAxC5Yc
+FjjtabGVMLReTy57o6YesVC/hZMNXtVGETavnhUGwQFdXLrBJNFdYDNjZkVrPiK
p7aA1IiV1RifTOAphiBXQn7KFk6AmzjjFGd+zeglFUffW7EZg/e0FHlEawsh8WMj
50oSmt0eEvDTAGLel1cjetBncyfOCYLhwnVOqae3qE0b9pMQMFszMHT9XjTuQDCJ
C6qpY0rJbIfK+rVe28UBDiZT9GbDFCMw7XCftOlzSTGmaFdkrWE0nu6EVcZ2KI55
9WXrLkxn6LBitZwYUqdHhGvGh+tZ4tJbQjooLxWvzIVRZd4zhVpA8UaSjiGcIZIx
GPGIPh/cscKmlhOghT0rvwXb8+o4piVsdSZabZXac2GsuD5ZphLOE1PcJ+l4Bn11
Q59TUFVMyHChvYgH2D4+62J8a6+EXXDsniFip/HdUbMzwyjPrvSfvYGbjtVWC7cQ
m69ctXUunnpdZYvCdzvEHTahiauTJFtV3wkoemTLejWTRHCKFnToDnxbK8wSKMc6
Vixf6Yq8KkhDM88XZJutwkuEQfuvGY8EAO3iMpAFZIksof/y5hr0YMARuAqctR1t
fNtrvX0irUVcEP9/UphKQ1k4nBkcXB5REcTSgPMYbMP6OHKHvoi7YQh7tLPTbqLt
OYixRSID9V87RrC/uYoTehU2smqdNjCEl46Eg+WGF/uxM7B/GqMbljcFk4H8gzLi
bc2zoYGva9JnFfnWvhDFLBHBg9wj30qOL1lnSjbX/T6ITSnJAD56IdaJ9RfYYhrJ
p9xXRVkx7e+SJorb9FeqKg8dfSCok8TwaAC9I+u5MKkO1NF8yqF6AL+W5mdrNLpB
7IwT1RwaYObloS5v46WSjoXJSAyGGFEkiSY2LeQE0UixHECm9DpxlZAyAZM6wTLY
q8TnUXGG80KYfv8LKu7wXEoyKQGothxoshRssE7KQrjVT0uKQz9okA3BiCSBYZrB
n+GCcTtRyumdVqd0ewJPn25U0WB0P76cZO/jsv2PiNNef541nINGLmMLyolUTT7s
dciiiU75ngqPvYpKmQTb7O7C6gXgEvOXpx4TbQvencccsG8qCG5C/0l81a9u9rkF
zO1JPNvwy8lCf4F19GclzW8dJfN4zf++oeJkg/HAis1H+Mf8ufOUUNbtVPELSbwU
TCb8W2+ayKNkTvZDISZmFylhj2xUZesmCDxu+LwSuv6jUe2you9Vnp8i38MzwmJH
twbCkHzqgLJUbQU+CsBzf5iOh3aOosbbv5DnBgHx1oiEUrskOX7RDgMqZOGbzjWh
MSHQDRJlMlImRXhVePUsZAfCkKrTu7MaIB+lQVhRhcwOkzuM1/vKjm+Is7U8mY8o
tL7cwAj6ywr+ywOqj25KjR1fF7RiyjJbP6eg5a0y+HkF93W+aAvunBnkdOEnM617
7338HpyUIJBVJ/McN6QiNY2tygNFAX80aWLGoko9FwjQkuPN1rTuILssMgepNGGF
06qYT9jLOMN4fn10EXfX5PHb+jri+l6hyh2xviiaUKBpNoYVduCAJ1WVwKxQ1Rye
/Y4LaRqPRhv2ZI1szbmMFu9QXWKscE4L9dVztVnGMtw0P1AQSAuau2HFJ3p7o31J
sJ/ujYmhSaq0btSbmY39wiaaMllJSi91RBq2rLIs38j0LRz8XjNZTHKgub+SHqdD
+1X28obOO/2/jw4F8Mvx63q/vCHq/m/xBwvUinCSkItXTGl0n3/VsONMxAJ9Y9Sr
g19j/j9v+BICo69IRSfzckCxCaLe85rUkRLxJFNL8qkFpi/eDXpJRjgJG+/nywGh
0A63JMAZ3Kx6O/7SEVwdM978tq4l5npb/USgISPNIUq+uzc1bzx7OSmMnxZ1sTPT
dNYK5Y7gdyHrAoFoCEiyBg85nrfYtHSIHONIfKDxLytgrmu/Fu2F60BLocrKLJ+a
A2G5qNDcHR1Q9LNZX7vIdMdq3+4v/NU+7Np/Yr2Z5iocixF2YZybF1aDQHS+GPrQ
QKWluxNguSoSMiKyyVi0LXJTL3AD4xOLNZX/38VvTdFeH/U75WsyW+SaKQPG7iZq
n66nNSBlLkeyCHcQg/DPtyX6aWqNHoQqlfXaahXsmZGIW0RzCq/AmtkTmthrSYc0
C8HrpljSzQ0jBlC6uMTSOTnXHKgk6amMzgp1YN0dVI/U6R/x1wxCY7ERVwjXdF2s
97ESgwA/alD+b+XRfyWQOmGsqRiu/SM/IAUZn/8jTnd+hZwajXqb4okKMHBCvZoG
aHqZPvlLYO3GpILG4+1YcmJr/UAzrR2+3/fJRJgiCZKrrWEAM7BkCm/cwGsJfM+S
Z53o6EzMHmSdD+ZRteIEwu+9rkc57A/i9IT7yEyVXl4BMFmY3TQy0+n3BDb5ZdOC
9KEYtjgBwZX+vr9Pup5c69BBGh3Ynto7lO5qaU3UuEaK1Dhhl7CQcYBwAUw4QNRb
uHDzrMw/JyE0Xtxf/rK+JAyJV6ppwe4np/Cd02pTNrt5wAiQvMzZlFli8GrIdG60
ec7wh/UZhDPAnO2+/QCZ/khCZWTPx2X9i1Q7E4PD522sCJLsofjEcl0Xj+TiYTZW
cO4ztDmNSfiF+OfeBJPBHRLp3LsDQUVs48zkM8+W17kopXCvN4jrrF3AyC7Bpnzp
lPTu3431L1xlaS8K8G+AmTJMaxtXAt9Zh3d0eUEcrdYnNlHO3byxMIrLxhpQ4z/v
Dh13mdNmQ/GlGQBJDqeIOMCaEGxQ0hjUxOvNk6si2OQYsC1Lrswafe0MRHdzJAKT
PpAqzOzmGxL5zMtB5YMvECXDdPDgITzIMkw36adzMC7DASo7TzifVaEyY6DYK8j0
iwh2FfCyZk/CJNd5C9IEMxe3GOA7UeSysIvLNQfGuZV91NMlZccf3jH9kZ8EXTzY
/PzBgJyj8IfdzhC/nvGdiR7dEYPGO4prNXypFz3UL/Nma0kQ4Jln3TZdA+RGQZc1
G08qDxbLJ0cJtTOA8lc+huWjntk45VhobDcVK70hcHbuae3FwszBUsYSsyL866Tf
KT1malFj5pYbc8v5OBYWh+ATwbc8ADLmRgG6wUXeebKtasPk2vVxDkL8/oJb9EZ9
eukuYBgUYJlNMP/O3Ij2+nCinEnMMTt9kpUkEWi/OkH7HftJEsJGamYvlh6+Hyaf
pjZ9ewD0lIPHVxR1T2wVFwLHLY8gFzt2HtNZlKeNq1HUVLW7bMwIjw0l88t1ZxoI
l+l/x//cj91niyquUGLFCoPH2lfuVcr+ep1UWT17qsJnFsXMzMpOZCy+Msd+DJog
C+4KtgLQh6D9Vfwdpj3xNLkFGX3K2laiNzZlVSc1vjpSDDG9M9wY7ZUEsaAC9o8r
mxTRUTyLc5L58GM0c2CrGI1iK6kEiOZtl6EQwzDtOFvOCOcJHGr/iL5hHXXhlNFa
tybdm7yPRGkSO/6HNnutz8vXiWzIR7G0IzbvcH/RbaWnMakCw2oDxShuwxlWHI4u
2A6jIcuT+/nhH5tmQCo+Mm1lTeoEwhF6QA2LCnkCmAZK7pGua8/IYFzEF5mmow4P
Ca+wYxrBsikGz/X9Rs/TBDOvvOXwD2ml4osCZjEbsHS5sTsw2fZ7YiWQYZKMsVzs
0uIqvd5IVHgG36mpLpJ4HwILcjXYZqgGQu26D7WwspUBXsJDFhwrDY3QfyAHsobJ
kpXuGh0E9ijvSiVKXDtt/SCWYfMC73pVwkD9mQQC3T4i/kIkb4RC+Fp5iwVMmAao
5hGyuNZ/lzU+hIv1PlSlgweo/ihUxlgT8FIUOGYxOouSjhA4OTBkC8lzdOfb1Kah
Y3swl27SIiZOoOwwV5cRuiPonC0/L8kgaC159TLiYLYhBNHog9y91NU3fmbjlA/0
+1ppPBw7s8ja94kWUURc0GekanobPFh4pRiwgK3kgiwcYw2+CV/2e3yWmXJoeGhx
QokG5LBmpZ5sjtSFOsYjXgetm7Ng7yJMDV51aYl08pxKthuVV46ppFUC9Zu5Gjxm
j3gHyaPrCZPTPCWmgpREj7+kvM8EmdzmiZ2AVclJMgOCgQpKRJcCNZfOiwwIcvWt
eVfjUS8DhMpUec2TZFCx2p35kN/hIDMxU6QwkdlnoWxkmlDLaaPU2cEahGjllh8P
p0gLm/A8d8HSgc9mkRF6ei3tg/tJjxfG2QSKBVbBuBwZ5DZB2w1zGWrkHnfWO3bS
NlGwgoo+8qx/D45iwdjXv6U0GCK3wnNaSXpJysE//hsSijvaMh7qv1jk0vDWIQOp
AYdl4Hee6whPHA6+c9gVDyEJD/8udx55NT6JWaFTy3VBXDJMWxOfenbE3JKyR1nk
GoIy1KFHZcQcZUMBk4iGQQHj9lhb6qilTJ8hLtmLPAf2fiSumkOYXNJUWpUHCbLw
sm3G+a3+0sG31Lby5xc/oYMK1urJ3+eeBFrJ5dva4dBf4KsT/+oVEnRjcpUiWXKa
ELx8r8/igsNPyGId9i/AWo5qwFbk7uuwOvyv4o8T7pQPVs1EizkRZZ/84t/qgnda
5uq7p2R5RoQNV6rHFZKOHRKErDN8gki/BunwhtF0IvEChmwFT725mhOWLsRbhp6d
jeTX04v3YuyunkjrRs8yfL97JbwmK0qsOqPyZ6iobApQDR5X4Hir7aWa1klyvpRY
s7Mk+t/0T1x2kWoCPq4vCxzOwoFZHIAYUHzuLnQstLzRi+bvbDPe2NrCbcMsDW2N
jrbE0+MHHDpdaXRulZpHMSYsdnXlG1/h9/bXszQtJK9IDSBOlfFTWk3K5G/5RaRQ
YYmIyriqDI6RBi0DlAERtW9bTkBCTeja2L96/GtHUdaMWP0njaky3caCwP9uy5ms
+OZi3VwkFea2vFrg5cUSYsyRD1Mu5jVtLDZOa6pTYbY48+g+rUszVUK2ygC5Qq4l
tYM6hPm6w3dLDvaMNtUBqwkeqZcs5qp+7Vov1gB1iXb5zXRN5qqsnkaweqSZrNTe
9TkRUG7t/i2d+J2QOaCpvGfIBCbNs3TidXYTpEe54kpz6FwM3yzlxVk4eUEvOXJo
0F7PqgDxKyoaDyWeHiRvQbA96fYUyhPhxVq3AcGpz3wrXson8u3urqqy43vn9pG6
Eg4QKx84spWcGwduJSXap6k7/eob6t84JKwdWLxV9SfFBganSshR4CwXgjYYTIh1
iJNIKD88kmdgr9rKj8d2yLGJK4i9VvbTyox92ZP3eQzn4y5Sk4E8XziAhSCOXO3/
S4UwI9XzOggzSUOiu+kwIIlSwQ1H5RY6ylu0w7Ugmi18dtaXYvxVSCKL9EhDOjSM
38HF9SkJoK84x+NiRLDRtWHI7T6yFK0SbA0MPsPgdxn7Hmj27GOLV2/lPYAVO+UP
+qkdSRAO6lGl8xiMLsd+9W7zm+TKV72inwODorykqswM7LvSE7NXCc1xqU3mgUM4
lK/1azTtPVClERtEHWOp0FWyTmM6lI10TnlTBlKKr8iqgfuubZ1oIouq2baUnSh+
Rv6gfuGveaHXoldj8HU6AM1G/iJJyMxlGISmh8ZjeoEQodQ5IKsYga4S8jAATbyQ
8mU2SLOsRQotZxWlCjW3ViS4A6vcPGQmT28q1wUr/pPjZxQDgy+JdBaczsAABSUx
d/C3iSBuZgQnOwRuNhJ5GmMvUY712csdpSWbjFN8FvCkY0PnKlInIdOydEMf4352
iaruHni4jmgSDK7MFESCGl5RBG0QYkCJBLfmEphzeWHb8Pf1aiHHmrEk0APHplr7
FBGqXStUH9AhwvEDWYvlynpFOPHWaOvsmYiClYrFyxequHOyhwcpN1PeXKCD+C+z
H6yKMv5coQgt5b2Oea6mcturFyilSn4rUHu3goZ9oJY4WgnJ+7FOI3jYZfyaYhLi
zRn9WKqbK6od645QAMNwDMPK4ycCaTEEWLnhSoULRipkzGPAKOcx4hWUr8BmVycK
EOWx/LS7AssehrwQoT+xFR6uv4uF74CoPdb3JiJD+tdzPSeP9J3XsC6RP1w0ta/m
eHHXLISp6WcrpN7vOmQG5g8Yu0MaKR2BJE33GczTrBD8SR2mkNgnOihVorLSPY+C
oe1Y/REQSa41roJZlxcUv7O0Zgoe1HzRQe2lw7Vz/fvm21GbvumKOEvoOOALnwxX
RhBrZtqTEeuUwMwms+CLKg88/qnfRKFwKkxdJZYs83fWDwYqxz6NJmo14J/Pd6hQ
6Q+bb6yKxypNt9VA8+keOrZKbeX64DI7uWAjZdxuQWEUVTnrgCnXAY0fi19J5gwX
l/aLXhs8OHEpIwlwg3l+JGTSfioeZBCYvRvAjZOBKowUE6LWUAKUT4JbDTulvz1p
cLl+jz4NurkmSTcJJFNt17k99wVPGiy6QjWZc0K4FYWZ0gwgMpQGIunTPKGuNKFO
SJYQXwEOvbxH0ez/c6bx7DyAEuEPmSxyN2zdadsKbhGNIirsVd57+9gkhoQv6K1D
p/pvUqwrB23u4IHRJGxej8rHVho1az+QUY3zvIbdvQTpb08AyqrxX4Non2ZnFvVn
OQr/g8YJY74AGcEHIRjlXOVVH/4seAk6vMf7pqdtSyu2oebrSVkf2UTrJk8SqSQz
Sl2wbOgmc+EKpB8ZqqCCyDaFay6oG/V/sbBpDrNuAa5ikx6nSTUn6OLYR+swhI1S
deyvVAGLTuJRkvJpQRorRWJlA/KpxrbeePAHN+Fn0O3ovwslqb645z/Jigq6G9Mh
eXR5pkVNedjmTItBVE82cYMBjPI/dlOM3GNbp7h6wELbGqeAnvJjPMmIRKQcbuSO
N4SQO74dP1aJktyfizjiaVXyqtmDZkph8XSoIzDqO2i52+RPrTW70Nh3BmsNVJ7W
WzXJ7YVu6PUIOXdjuZIiYLrJAagYnPVWrt79tQWJN6RhraEqYLoFUmEy0PTloK0w
LFdv7HH2U9jvSIP4zzxVcFxNqArqXiRSiXPUsp3wwBfb8J4nKNHJPtIZH17iUn8A
pLVjCZYfm3Lpa8DAQv/72rbYmM4v2OWalqqKNcXES4yuVldgpQis9yamjGodjZQT
3QmKmVnig6dO8bRCfBfVsb9CLOBlPrkp9lFtWnH97J1fE9m5d+bjvu/YlwlhSniS
qz7XiWT8OhMyGeuS6zY2OHefOXD8fMebQYl2+8oHLZvsd57FCBYaTE63A//44Yef
P1/pB6SRALXp7RTQsMR7BmATw3SQUBPSMpbzW2RV3TZvyGgq/2yTERZX3q6LARLJ
yJArNjXQ4LoHBwuaRjXWHOSf8OkShLOhnV7QY6KesjGyMyogivY8yh9fc7Ocm/6Y
z5JWyEUwfYgFktvka/FGBu81toV24jZSu2zmcsuRMstyzd4Mw2gTlX518VVo9t/S
QNZRvv+7VE9qciGkoLaOoPhCx01AeH9PJlXqVMAloszyHYZlMCFRlNKw7lTPahM1
Sg8qEoNCrwztT25K+szG25lrJAiT4VFxJweTG76TLVUKZ9XvXtk09CMNH+BTjt1d
kTIeHDzc0JsbkJwc6ggUVp+0XMqrQvp8J7At3cnJ7AtWVPa1leh4LjoCYwWFV2f0
pViue5t5xLwL5yDBRo+eIn8nuvIa1n54E/EVlhoCLNWKn+5hC/Pz71H0ELMjFfTV
u6wPceEedKaRB1qAHpe4NLsKrJvBYp0IkTB5iVwhkIXuwUFqVfBdOlXl+V7/X9xx
IbH4sv7+4EUL+eha86LCUa99kygvDoRk9c3LnNmerm4Q9WeX98xwFDmzSuJ5CSsl
+u4158xOveyiZovGxQ7ig7HhoVBPJAtJiTR6H6ozCjbY5Zm14Wa3QNPBw39/G+ha
qyYKMy+Tk76JeBML55HPlOEolFnWk6108PMkn1xzmCLHGhzlUVQGwo5V/ZzI6zYt
c3IX6nvJDhpkLdaW+A0QEOxpnLr0m/moT9PnDXIfhzK1HvDuXrhrG4GUHMMocdnl
Wzqq+OkAdi86FuARDn3qDaw2iYZRNXEeO4i40nNDH/mspCyl9qZcSvyebIDCGb2U
8HTZEO//CrmuWCLAYoLqag0ulTz7QmCsho/8mwtZ4VLydzBI7Cbkz7DEEd5T8D32
kxl8eX0lU+BaLsOQ3wZRWGhObA0tunBxM/n0WUbtqg+VLBbmhMTJGSNk4/Xnqxjx
662p03bbCXdTfUgYEewf0NssEOa1UFMaOzbm5YsXWIOEvbQ6iZQVcWC//BKj54XJ
+76F5RzcWHMAcmJJl4TlzgywGg4KK/Iloc/TUS7hRBdTgWzC2qrE8yWkBmDuHP/7
1lV/IaedqirVki+NDRg6fk46FbCKfxmC7rfwt4o89cv1fLbB+M3MEj9mmy0UWgF+
U5KheLTaVr7mbjQgmPlqcHwdzadTrRLSpY+yxmlsz+zclJHVPlWLNlGcN2xY9JRG
s55/ANt3WQsjPX71pRxxGV86CmY+lDio1RGlAAN9EQjEJBoaGhEYbrIRr4PnHaCi
Rtxpe/dy6h6h5RokvC5qPVDaHh7zJa+ZIZ1ELCCyrSXRi4y/yy/Zwm4BBMg21TKl
4XaZF/I84l86nNjoRz4bZAof4FU+YA6eUGmz05tZjMqZjkW96eD7smpEa5Ku1eHr
9Fix0g9Egb8ao84eaaRUF1AMoZc1OrXlANkMlgIR0j5rWp7vSh3PDPik5Ebarbhw
QQU7EliWNPr+KUwf0H4b/iWITJ8lM3RF177jQD1xNMAtypYLIssuaxC1NKFqjyUs
Fw6fDabfsOdITPRZZv+m6s437ErCVzPXlYX2C1/JKT3gVfMk528lmoA97bac/JBm
vcJ0xVdbkT/hsJZHMOel331fV9qK6ornizqsN7KpN4/MnQQFoVUa9MQbVBp2RqOR
hp9Y8Ws7etu7tw0heoyDxw5xpT0QKc7zCgHdhscAV5dH1MAo6hPrSjU7CqRJA7Pq
LemQ3OrqIvEZI7voMvl8N86XEupbSAbP1IaN0B64VoASG9VKHlEii/BDSsUZb20t
b+2AXzfRUDcAyAWSRFHDnscdTyNBbGQLOIV1qMe73trua4e1iDJI4brRjzXn0hIS
d1gvovoGr+tjNZKkCpeQAumsrFOOuMxRLlxNYO/jwZCwr/S+nptOWNtisjRzRVK8
0rDCpyRDnM8YOCR50iFlKTjwLq6cDlVxNxQMV79b3BcGNKPCRznrHiZ3KvMzHrgT
yaKEjak2G8U/wPNhwPQ1qaKnyhy68kYRc0HunR1Jij2IG/BZjdxq/iEnh/2ThDwu
7YkJjiIRgxzT4QPeG/YrPi8MM+aK3zJJI7VEmn11kDhM2cLAkjnv3kRhqQl9C+Fi
fV/tyRB4sMz4XyVxwQ12GMEPBhsY7fNYKgItxq8IuL4dWKiUvxrvQCfC445YjBaK
NnbcS4WCv1UEkQuUcjZJ+XME84NTnT30nRYNsE89VQ67ADntpHas0RglJJqmSPoK
bfwzE6CT4JltjtscFIAmaolOKl66C/qUxPsC7LEZmw9NAquDKipb8qWm6kiFDenV
jgWcjXA2cK2H3FBUE4z/8IHYZWH53ENB2CFR4N45vo8cBTwHjIowIC0pml8XyPtE
GGS5l94RKSQBl5eFC2IZ7RSXlZuMYmFJoxWt0gchB/NUbm6PFq2uFUQ0vaPUW//u
TVDyX104tKvfMbWWEfsBci4DuaUtZ62udIs4tKl3dIKIQtG2TmXQizJK9tdkNLKO
i57REiJL1iIq/oFPKXfquE7OoQAdFdjV/tt/VqvYtgEoz22i56sFwSCtxeA3t/y7
G4uLa7Fdsw7BsOrFFPdKsPVp7LYacA6qSmluXP6brG0oZV8h+q9KtRlyigHA+4Cy
jWKCj4+o/Z1lPsabCgGUuN1e4FGQ5Ja+L2tCBdE/ALMab+3mpguXWqZYhkIIvCXa
cZ+1WCMCKQzv0Loxc0M+fNNoAzk2oSQeGZlNHtMHIgrDIvyE9jqJWVhVAnKXPI81
KQLCxp184ueVZbUHAsk6/+z4xBb7oruK4K8G1nAunxwThi9gGxp+eGK0JUm7cWU9
15xCq0KQ8YSHKADwt0yyUxhlx2YUqvZkRwsN0wIWJZWfGXCaRlxkmcrsDUjCfB28
2BqcdtN29F9W+ePxRaxfhPqwr1PN3MVE6NpTaxZWPePuXWCvQYaiLTMmz+RpQ7yx
OuqA7RdWaaSrHQLYRRI9JBuNf+hA+1f5SUWU8PU6yWYfp8NysqYX9OWPq4rhRpFw
5BXoYVdvfP+NZ16lz0valYWW+Dbwzu/bMVkaqKVxNOV9WcqnF5lUGRzz4YmCDLHq
FgSS8Ne449PMs2MZ5DZ3o0znoP7zYN8gG0jBrFmGGklqJtgGOsbSRVGm9IiEXRIV
MtOjxIn63+eMzf/iNtdEIZYdYy+rtprwr1PX5+LQ4LJ+aeJFunauTsvF6QxRltD+
gvf+6hPxSUERtMMmA8rdyGUFLOOnSbJY7YY+4upa9sWeywNclW0/G4V/yw5MfG1Y
vk5Y3gv4i6Jb1FakgDyGlKq63YGBdv2eE9ZzI55XHKUucXlLeFrOx0E0iGHYMaQV
XiKUeOqQ2qEVh1Ps7rtR47o0/m77cRNNKNKrwUXQfdwsQNQQLXbwdhfgLqYOpBkK
FvCc41iEXlUxinc3ai6GPA4MUg3gI9xZzep4T6DSBItN1D5oWE53M+6ufV7hcjxm
vMTbUDv+4j9hPUsy/jQttDQUDpVPzVYk0hol0SactyvMNtHSZFEG3JAEk7GgdOO8
SzLKaFSfqVuwF7vchxS1VCGNOTCYMt4a3hVklYbEqNkifV05SkRcvEFypXlN7qCR
wOF+TunUGg98DbA+hGJp48OH2Jz5OXc12pYRZ7fZ3Ullhy/zVLdmoppVnMqYc+LS
CjlMwS9IX8+awL3VsVUCd2q/zHu3Y8X3S5TqSYE91KFu5jQXmJw4SyQ+7VlHpLZF
mOiqZ2gvYoIRv0JTBMcQPe8BZyVPdFB2yAShVFiz3tNo8uPfy35jWDmo+vAn3TWZ
y+p2KzgD+Y8qfHEjo/ZNODmp1O6rYrZGel6iJKRE+KkjYBgCpP/szW2+igXdiZXf
Gmpv8ZqG2tfX7jDdSs+NlPoWsYBCUAATwL31AZkSkAI/o/2wH5MRsj/VsDH/Li3t
u3wjSsgMpxBmD6KW4JgIIW4GV56qkQYEY4DknTPFloNK7uYWatmu6eiBi0uU8/g5
2Wbe5Q2O6V6lQycPXqjYGwBm+4Qj5sAPRxIsaK4XRZcgP42p9/ovYm6HBDF3jVlt
guovNDhShE/mOTF4zqAB22py0Zd59jCS+GgG+lnbiE9U7+Qms7vZy0BiyWtKVIG+
A2zm+U4XydKY1z+Eer1cLI7ROojkn/Pf1Pa24g2fL09jm984muxAtseBGqXrPr9V
im0nLqwmOejJjIwhTdwISEhA/dwXWFoX8nCmvF3EZFADA3vBFDTsUe4XFlbL8WKZ
y586AAVBt5ufBo9F7rx3W9Qd/sNauozUkuBdJDcGZhEU48inbMilHlFTm7TefOWh
Lv2cVD004axApmPscd/LAllmR8okD+3fXzgYSptbBg6rv2YsEfYO+hdUDwBVOby6
F0QKl6OUMqLAAPVmyO0qUhiN93g5HCpBc6F2sSFTDEJY46U2p4+g4+EbVBs2WnoT
j1NC3zbyBiz7QQbp7LV/4pMmlVMCxb4ZTSgOxZgIr1K9Idx4AiiSlQ4vuUD7uCc1
QACb/BjgPhbsbe176J8zDZZeVXa/NzUdlkbNIc8v0JM6JTYoU47lzq8K1eALecnC
jl+wnSVl9I3u0g0Re6z3gW00PCkuuAHmdhrWSvAfHxUrTyhQynbPMfqFRo3NqKXM
qb/oGtVszTWhIXaaK5CzrZ0NPlPx/CIoUYCG09IVYBwds1/l4z9c4vfACkJt8CwI
OS2nrhDJrRzR/nLJfFYAi6WBgfkg9debkbKbMSor1gCA7R7GlSoomauGVDhecS/k
hA3whyq493a69t42PdflE1DFM1LnvlEL5cVmU3oq0xg1DyvjlMkaW7NOoP8Ya6+z
Mg3edtH7Q/nJBa07QdCoqD88EOFXPk+ol0ji55/rbvNC+AjzDvzAyMoVrNXGW3ui
Hsuaq0o//ReNk1zkFea27J4MukeijtxA13W3LP9m4ynmkFvt8cCduiuAH3Uzj7JS
arTW/mDM8CMH1vJI7lW1E7eCgkNRtx5+H+U5RPJm6oo4m4DjT4l9ChnvaWhgkbNH
PSySaVYUosbQyMi8grS+4i6mTQcX0lv6e9jvzEXPsuHQQffa3+dnjELEAuL//a+f
aTL+oGxQyODaV/HRu/xckVKYFDUOmRhh6vPjdyWMKkul7FZ/od+lKfKfGOq8j8CS
aC66t+fZ+JhWlLEkfNNP7Hko+U1r4VS7EkSFYGjEuvQPwQhOfvNfuUnZ4rzt0JPP
XWWWAveBP1QN0yMcfr5CgBKjEjfsICjQV6qlXfz2mTqfN7s5jzIJ4bwX/2JnCRrE
LFpLF7RV0dWGbVT+Cds8LMx7L+Uesu9tWHO512+sXFbwxHj1CpSjyCiwR9Xe7IY8
fXaWu0G4gjr5xM7bONWQCxLeNlS7m+XHk14fqpY1JjWEnLnIgX5AgJkvtKmtxxi4
LvFD7lUj74QVoOIy5HdPXQJ6LcN8aP1HRPAQhWwZA/trS2uK7EV7CXTaHHEu4n2r
WLAdigKI31aOq5VRHIZeYwRqr0JkOBzCIVLjWHaT8qTWSJt2IIMrc5U+tpBkWTf5
6ep6vS81qWJYj6YTSjsbKvUdtXKkXkEB0YygyCqwDtfYD2sGqhB29Vs7ARjGoLUc
NSFYm8biXM7QhoBZU6xCTN1L8+4900Im0UP9BT+TUfMkF1TVHvTTBID7oLnAnNBW
xUXqFzgXMgkBr9t3VeqTOnqbNPbrHyKbvJ3z82ErL08VpEYiX9LnEM1wIlqC0JiI
6HXWZNI8tOhFO8E/o+r5JCZVZ7FLrTMnjxwpkrFE5/ZXUgWSCdPjVLPHLJW97aL9
MtVCUuuRQeoI6igRjEZFInuZRVa6y+XahUJNqZLqAV0b1Gaz6OVygdgcynsXg22u
egVSsvtfddWouCaLh7PwqgfeZNLInIqLwv/NGRmAHl3PQAoz3vjG5Yh551Lb3NAL
3LM09YC3Aasn2eKonpjOIf+RGHA7a1IST7sWLd6Luol24uD3aKVPJR9EUzH/Z6UZ
9NMjnpcKotWy+lOayRNOJIiZ+yJeMAvy+wQfSEe6/i1KT77Z5J1ixMGZ726RNMUo
vmC1uV9NHfA1yWxkv1cl1PTJj+pZsEYWyDdHRbDHHN5g1DTLRIpv0QjM3KxgVj76
cc38grRHlGYsb2v+h+YHXQEvIdCVFy7QIBWj3IGFlLSYZ3LBnPdVU5oxWJggmVLB
QtatWEdmgdJ9jZITfejbgUjrsvWkcbXIDomA5c295c4SskeOZsScOAxLmAIfeXUf
v4EZ+S9ZfW8f3aZThd3CmhAPmiodOuMUFVubW90KwEjnyQRhTkFJ+ABrnu3Zsvys
hBxjtjNOB7ijg9bfsXHdDVEF8TNhHwIV2LNcbPJlYkQ1wsN4HJdYNCkWmYOQZLr4
iTcKLdXpSHK+AktQGHHunLTqZ8wh+CyP3/zRQFjIJquLj/uevbft/QQybBv8mDuc
OHPlXlMLYPLztFogCRrvQQsk4zO00P7J/p2vvogMZxDjvWDENpQz/YNmADvSMNBH
gGYX79XLwQGE3mky2jpwxnV+Nhz+Brch+hhSD5U1AvDRHkq+JWhcEQ5Dpx018OmK
bk+OoX8pKBAHPmvQ1enBThiNALLB63W2gK/2nPlq5mgUO9UQcWP8//+k6KDTrQsJ
DpViZyPgiAvD9RwVji5uWBzFL0JFDnCnEWW8WHnRNHyAAcFne9N187rIcvxKsz7P
KSvOzCn1aqbdHUVCZm0+j/PZCECuN9eGJg0LwuEU+HqYn5XIrBfbdwQ3pgQY2/PX
yAZRUQi+3Vur/+6pE30DDK5ejpKT96tAFO4ZbJ096nmjHcrF6d+l6A1T9s8HG/cT
O2MCr+VGZ30iGP6NwcFaE6YPyhWZWj4qkZ7+O4iA/0IeRVW4PxURjVmgFgcnmJjD
EBgOobnt/ufhNEYPZO3rHvaO3fMBA/m/B/H0DTdCwjjLDnh5nhqnj27NHtk/skNr
4V2r9/AiH4571ODKXvnO/r+7+6ZHrKTFvDuBxDR7Y2HDBaarX4+qUw9C3j0Dz84A
7omSrVko3NuVuAm9lWZSynr7g6HBKEX8Nz7V3oK+3B/4AVnrC0n83wFHxgqocXnu
xUGLRMSIKfdvPxImT27dxQJ39d8FXoRT73WnKig96XZZv/JlnMl8ad/QQKZ2eQmR
Tx6qsAqeYsXaukqCu9Wi7/n4EHq/UyGzskPhUoVkkBSFAVNaqUiilelpnN+LML0P
b3rBEPMey0Uh2BVboNvSOWbpGX7aYM+77wQjYnhhXXeNJ2gZtNoHmjlRZn6vgmZy
I1C453Ui4wMT3abEmSIaw8Uy7MgqFYN9M4RUTej4TacI2Nt5Y5xiPjg2/PmGuxVc
twBn8Z9k26gqqb9OMclsguJx4h2th8rL69OK2egqULIRnTguh2G3Itc26O4jdvN9
EPrjTFClQ07vxIe9P9NyzmcQLT11shvMfTA/rOsSK15k5AekCaacQPzZOhNF5HeF
DzIooziCsw8vLqb6Ci53CKxrw/JFftwnC+bSTK3/HBkrqgJ22W3Zd+UdCsM+7B2W
IV/g7eFMCVX/+FVZwOm7HGDB1lNI2Tmk/u/PRsWUeAfANQYEdA43IMByx7srC9p6
Khzt6aL2npsAa5rkV/UK+j+leeR+49mi43JOIZqctknFWH1Vp4IgMSh+b7s8Pqla
fgn2Xs5YAA50Ej8/ic9CDcwihCheMHJeALAaJpMm0f2HLPSuqSqIdcf0ZTL62Hyn
VYpQnz/LJRT6bZm4F1KIfZET4D8+Uv6zFqU4zP9MRHtvPZGB8ZXZosodHPBKNvmp
W7tXVd1aVptCmnQxGO5bB/XqATft4tY/G8qxzHsDuOjndKPbcZaPFbGW/l/01zKF
ACC7BI3bOAwk7xVtXIHtj5KopyG5ETdrn4urO8mgPza38gpcuO/Yb7sYmVd0pIv+
64TVH9jHjzR4WCF+DHemkv7Uex6w4H3MXl0b4Fp5u29bbfsr/e7aGyPADSKPTe1b
WkJEQW8/0XMhXr+8Sm+nqHJJ9oeJGujs4SsZBf3DeNLWwDk16SMCMhHv88DZVoiZ
aWrrWbviXP2f6IwgaACjn0jegvI4SH4R818OGsbsNAisD0wqJyzEgDIeZhkqKutB
x0j9W85A4sig2LF4N8o70N2FU45PQEpsbK/50v+em79yHBaFfUbnoRPulvsCmO0n
+SrPBBkrk/mI2IzmUV3SG0eByijbZ/zyBviv94QtDpMEa2zCfIFqDK6Tt/1hZHne
/D9nRYj2Okx7HgDNVrJkECESPgVH/BkRROohPF4GCbTFL3z09DuRrO0DAuxDaWIF
Sqw+lgYNbNMnnkncY0dRj0OCFS6aQPgQeJq65SeypqR/hI4OWHobHGt7wpbfEj2v
nCwjvNbZ6xbEP4fozL6FWDNGk8fJaH9xY7+H4EoY532WEB3XHdEJA33jErAYP3tm
eU6N52dYZ60kj2cCF8dTIiNQhRmIwBU1VKCWJRMIBx23pSV0/1sVb9xM0TMIvOff
VyGoSFXgfnpgCMdyTSIbnuecjWtsLwS3+OTUA7cwxoHY1ySj8nLnZA/j7jm1VoUl
nAEdS1CsvS+EcwwreMpK3hIENU0cqFMndgXkarNHgWgTJHFlzJvi+LbeVBvCpqqw
mZYSuhoqazzn+YLIblEThTyW1mxfb25ZZu0GDL37mtbAvMXOgS/sEEBmpd8a9U8m
ajhtKmI7pXUH8xHZ/zqIgGz4TdKt1IMc8JpbFhvzlgHj5ggGBMULLSR8As5aX+jN
mw8xl45jlpQEv/hsyrCUrsHVDaIfzEY7FuVhP/P0O3pU+UbpBYkO3Y6f23x1HoDb
QZo3DrmXGYaQmkXgRNxn9CflT3dar2GBzu4oWEJIWkv5U16K88tJCV3X+9gsOCc+
EKfPi8G4WKfiY5tESgtdzqPH1Swwt0oFkqlw9ZFXMl2tBELO2Xnc6CihHt5OIVMI
VYasJLbu4StsTZWR5s1MWsVne2fdMDCok2JlzmjMN1WGzjLT+zyTvGwWWn96VsEy
uWxyboqjZAh/EuRyd36vr/V/EauLDGbwiY3lu5C0uQeqVwfOkY0ZkvGhFOrck/MQ
hR1Wg33UfkkmNcYfkB9ewHMM0toKDNmRqIrnTuuzhAEbajHRjnn1/Zt8pNv6TRXT
HcwuZRPYZK/hE0Daw0y8ILIARpkCP3q572DWo6lJhJQE1ENeZEefsRVghcznuZOt
uX6wh+kajcwOajpHewN8A6ZR9KoSxWeT/aYdXPyTlCGFoJoMmTmSoTfAENn/69DM
Bje0Gc2i+diJKDOgGRN/cNeXDfEylcp8l1MGZBqSHBTwiwRdvB4+q2+EI/SZLMFn
PocwxeApaOQ0CeynH5PaBG5Q5EamRVBQqu9bRRryU9YNX7MCVTUGFEW8Wlo9wlgM
oMsSHBjLBWdWi2z4Camw3qwM26PweC23KgOu8O9geaW7AlJAhOVfiSW31uEgokjE
AJw/ymwaXXUlz0iu/PBe8HRIowZpaLvwnLWA8FSqySxpu69sn9faCOnl8YyXHBfe
ljuu3xW0HgCuZAUrk+tlPG0q96v2rp+mdxzKK7YOrLhzo27h9PgcVAypTff5eFdZ
6emVKFklG0Caq2NY4RG/YJDk2ROdTOJDRE5FQQVUPDkFbJW3tY5+whRBfTrKIO1N
Xpw7BzPkbDacYftgSBPA6p2/B0ZP4xL7N1ti2qlHJmVd2OW8qfDv5Tnr1UiuUFtW
a8VcTPi6ygbbVAjdUoC2BFpomxnQZBdfb21hmaAIrc1q2E4AmIpoAOdLUUtfvqsS
eAZgtAI6LRo0xyioG9HfBTnbREXTXNcYq1ezJc0o1KGayVGawdlZB6gQ1uFK3vNY
DMAt9U/CetD5snU4Gbt8mnNePDAibJLqS8sypNqcEqEW3O8x2gN4CG+PdEEkLGWn
JZyjknAnoOdoc/mIYdgHuAn+k7RQLMYKYu2eQSQfKvlovn/wSNslX/kKo7pIjqlL
TjODzswU+vZfzPlNbXUz2l8CLew5Gzcb7TiCGKWIcb+uwvu8/+W5wsHEaArMpgtv
F2oUvH2b7U1YQG7BT81wbjiT1lk3d6l4qzcJKheSBsijMoQ/8W2hwZMETUFUroOF
JLZ5xkOD8zej1eVwyDH4wkjfqG0psMy3vbPZXvHluP2lsZhzOdtsiarhFCRWgzqP
k9QHY3grsShKycGiKkRlXeFifU852ZoNGzS7yrqj6Xedx+QtfjwfI2UYFoc5Z9ss
jA6NDUIyMmlAJB3oWbQIp9SoT0Mmog444qSFQUGJ58LrEszyerwoqyFFnN/79He3
LP1WIjkMAmZKsr7DHby5vtKF+K99+Qchu0zp/MMxHZ4UvSOxjCrp/LK1DxXfx/F1
eCuFdJlbhdugjmIe2FWCBziW8UE5dOwSY7Dj3MvVcZuqTseU+J86YS7cBQCxVPSW
eG3/bTP84pb8Gztr72Bw/RkAxUyDggV+gB3oAlrHZc6E8sIfI3jFbmMKaP0EQaC/
QGR14gwmTOVlH5pnw478+HdqvUInLEqjAqMYPPfJ/tdeRRZdmGHUNQro61VLSLqm
uQX29vsXzDeR9pFTkNhMPwr/EeY3PUTYf4O/JjQDaT65lfCNn2zk/23ozYOdwVSW
6yj1P9C10N21lBZwGyDNb5G46sa7gwDNgWYphsH1ARqi/btQiTfju+9QJvZSuzrP
/vEjrqfkTHhstZ44uIRnxlrorPod2fJjwCNa6jPjKYSs4eSO5Vu5BbOGtoMKfil6
QxPXfcJNi2/SsSPaEbJc9LwcvvVB7PyhT8bAV39kNSNd6B1xrOjEw5hQa20cKpft
6F27vJw8jiM4l/88liC4zMoCkPnXYtjgtH9akcxO539OG4Corzvm8vNLHt1MaUUc
z/aNzsmpUiSJqf84A6RuxauXNWpcPurJJJzE+t3We+9eYXaGTPVAbl4c6wYZQXxI
4DsjvglPAqrthpWN44eXLeXFhwIWNmAkrWqK6ueaIFiPuBzwwVjztSoKDLDfG9ak
8R6ODMsFAYeRmXcaLF/D9jQ9PWbwNekuACVwleIxCq6EVGykvoXirFrvGfvXI0O1
hgvluK76aPQlWV4kcrTjq79VVI1mhjQV4Be51/7OaYKqrFl5PUAxmwJM2SDdkWlt
uzSlM5IFGFh7ajg54ssILiKo3Byi++yluE4+x0bnBYtbDgPuxyYrO+vdjVjQdhrX
6IGy0KxeKK0f54h5y9PIz2jaJYnXfu73a3PS3a2/Xzcl8WqwRUyQBcWiQSU8PZ7k
aTyk2gHKDb7LTGi7TtI87Ru0HBJv7vwk+NnjeDcfe6FSEHxk7yEUrD0RWEWoEPjZ
sAA3tnBenGvFNiRoCn76+E9bbSfbPeEz+79wGVUcCBHx8MtwbuAEcnm/mNNKLN+K
EEEkBeLwTHrPB/xrWpL+OnwDh3UIVbRf1MDrnFfI9obiVOdI0Ce91DGAcfwxrs1v
N8imgQR37uQdd+gl1FSerGuoAzh2jL2jDW08fZQR7rIz8jNF/gV3TUCWqWwfHuAL
siOu9Y1BBGi3MRtuBZaKKdqsAMPCsoL6YsiYvJaKKmJe/D0Iwdwj3GTjhUeOmA8x
j+GMqn10YRQHX7nHSrGmcyEsONm9GTcTOnce7/BtShz5Vkd0nNGHlRSWgSDQLcMJ
i583mueFbY0XXiB/2qzqN03cn52ZJOslqnkUxaNddYzUDUTCPmA1Qq1FIKRewllc
b2pqyfYIYCc5+IVRU20zwGyMOw+1Y/xbVVEhDiKassEYeDkYojuFjGl9F3ZpL/25
lLwtyAN1B8myaBK2MiJIOBCt07QVYkCdEStJD0S6YhbkhYfT1wHaVrtE7aXpYLJq
wRhA2aR4HDbE88kMR16dn500bZpIyeaJjpXoROhIg0yc2gUTCeiPqN3mu7pxDn1C
NXarfHQVybFAfMkFU7/IDI/FDAHFtYdwVZxUKQNdlV8usyrRtk6tlGmb41zC3Pyu
4xUjBOP/5mcr/RJHlfqEgGWcmigRTFfCYgqmpK6EnGtZF0TFArV3MNz2bsEQLwNz
7kLBzu63z3ABVS7l0pESjsAvmelG1HQEdJ7vNA6mFseKDN+bavceQ0mfHM9qsExB
JHnnfdLBKKoR/uT86sdPTGRnz0IKvv0VrZY+LJ91H6DoXiv9jXHhlfntSSAf5jKP
I5uPfnqPNA1OGSIGNZBGiYcheX0VIc09bymX4jAbMhd/PhqqfAlXYzsWz8ySDXpj
6QKK7Txv1m6DDmkbsaJI9FMfzx+LZRljyvVjA+pC1havq80Pu/HxwJoRxEqSaGT7
1JiBHA1Ack95h+6ICwhWpClNSysUHPYiQTlOvEBza0Mfu0N2xd8I3/bYDqjbZ7wn
ci0L6tUqL2xA0G+9yTUryyEuqfZ/kF4zA9XR5n0blROpXs7XhjQBPNJ3EQdQ7WnE
GNdMs9BSctk76lf4s9DuC4pjITBHsRqH17O3gBFnksZg5W3ge12oRZUY+7z6v7z9
/PhZj+UeymAynEdtuKYv0k9IdylSvYB2iubR0HlPo9ea7UPMaUYcrNO0C7/qY1zJ
EGMRXsybZZnhCJldqZ7vV3fYMTLDr9jWdS+HScEdb4/adRPM2H9XF7GPlXfwal3K
u2pwoP9NunvEoFJ1WD3JGHuZ8YmXUs2/4birfrQaV1DyQgjnmTBxQVi8cvSL/N8W
Uf77rlQcb/+JBU6ZXMhWE3uTQuMtCPRh/SLajHtPew/biZQWn0dUUg3kZpMVf+Wz
nzNYhDqvf+5rx3gKW0YZ27e98A/GDNCZIRTj+Um66IMCrVGESkmZk1xMO9Kk6TcJ
7nEuDdWIQJ6bzvSXvjvf91w6l6GhVcpacUWbaadlHj8UCvaQmGZjFdk5xH1/MCBx
WXS5BSJVU7JO0B4XETD59AXVZ+o6m4gh540qlMIzePCNj6GTJklV1QClITf+Qe9Y
zk+W/+cJXWsGiMKKImd68Rb7lWPJDcAPtashkj4UThncbjVx1hHSVVwicocyO3cp
kzPeMz1bN+W41LdZmerO8fzQjAVSGUD6jf8TkmAPvU9P+MoTRK0nYB4Ks0rLk4tX
eTg9RH4axwUV2Dcjip1JUm6jEMy+aRcLDsMaE9dMZERZvjGV8DbByk4l5tcG/WET
iJiZbARKmGNibQH33aOxBB+xp1byIxO4Zn0Isup7iJ6xnWClmDBYb47jhY20zuM0
LSHIl1Y0ZajKJWnIpjwON1w+QiXil4N9T1uZCaUnawVoU02N977ThAdGTwMvDHsu
6nyFEWpIBdLUw6+UjBoAPFwd/VRP1boJlfr6tIpHVn96Va41yeie8gjqEt3+pJBF
juS26ieAK9QyEuDBvMRd7Q6AFo69PNYdtEhv/A1ZiyxHEMJNHHcrkyXiFy23wslC
0H1ioYmpkTAKoQd3G4RjjtbbmZ6lndriZ3RcpXsbesb4QQZIAlxpHqLoDhwg4stG
2xW/YIriqY6i7MXGrH+Lafpun8yxmqaoaseK8GulTNVQ3+5yTz+ZW5ojSbRyo6p5
GwNxGHWL4DCiTkMftR5P1R+xZFDDPorxjDGoPDcMZTaQMuEdljrdjkj+SSa7dWpK
6nmMg+qbKP0V176qB+D9ZsDevc3JsC/V6A6ZRYAvoW7XMQgzTylmzHnSELFjVF5w
qeWudtCQAe/peZYLEgh6FqbLPD7cxneWIgjUDj/zlYtbRxwXdy1BVebNDC8uLqLt
8aqSx84aoLi8T5b7XG8R6QuCpZlZia15T2F43/AFbTFht4sI9w5NM+gEQRiMf0RG
4zplMtn4rzlPyM9bVROw+ljJL9sKCSX4ft2LVlum8tFiM8so4V127AtsD1WEfIy8
rfUp6ALF8P0jqztdb8FNXrwP4N1wWolpEv02xdqMdRlW+gZjJW+CJckKVqGwPQmw
lN64tczgi2ihDlklDowX4/htKulCoyJss73iMPLO90tpFfHmAz06/5XUIg99wOCA
+tCGnVTNNq7TXt9rOZQtCR0vRZMwfveOa+Xqs+5nIkKVLMtsAf6+reheiZz9yH6M
RIrAtQu4vfokgytlAN/HrweknMHmA1qyI1Gaxq1bekm8uiLSI+ARmaxMOu0QNw3K
TVUDpCgz9Zxg4R6jyaIIvznAGe1Ny5VK4KMocR8em2E/DwUApKfoJtTskXNWDMcV
gByIOUr6GR9S+WnjNXr4HUQqRT+Vx+BMqNK8hTkuaV941h+vvgNlQdHMeYyyLHiW
OJbUDHQvHAZsSWvB68wZ2XIrCzKHSj+q3FyMK7t6eAd0AroqUOwx4jsIDlsa/gxh
XgMRTlZlaqfP8l6I58eHz6vlXt8tPIDqo7fsbmPCXO2tyN9xWX1RRmSMpkVNYBrJ
E2kdPeRVU+oFTt9IPdCwELWRhpKUPxaTIcnLTAApB2N/A0ciA/FajgPtA+h3GrZp
rh+4iiYw9dN1fOBxatSr7YrPDalL0sn7lNIzF1A1nuEGKoOWhEJvYOJmXlbyabqq
QCbObf3IAAI6xe01ys85tn83ZhpT5WLtFVcfeFNqkcy/PndS1bFwp+t5oY0Ukf5N
3lbGh23LyipdvS7sKc7HCKexFVdBrLmqrnNRKZCiImckCilno1wPoOhXEGqVSXKH
bO//xxqTV+jKYMk81FS0AkwarRoV2EP2Tz3yHJxWGQJ5CGwF4268m8NWDAjkctoJ
F/WdEVZa2ZF+uno7XoJ9W6nzq2XNYuBfXTRO23nZoF/iOGB5rWkLsdiO+1w5FV8G
gjkZIq4ooh381h5cvVqawbcY3FA3pUCbVZL9yHmiLJ+LwkIM9yAPzdGMOoV4iAqP
m5xK5eMMF8F5eAsNPOXo0j6dsh6A1CAxXP1MEem5cUfl5W5W8l+Mge2JU9/2GZv5
+6OBrGyiuXMyq3wN+hih0U1mHoNmKIvpG8ujA5697Wz3V1Qdw1/fLpQJeraooWDd
mEtSiK+Rkwmti/NAtJokGxhi/+ycHNAnzAHmiDyIFUE0pabgNyJJuW+Dlntwiekc
+tYOi997ospAeXhnUe5l497o80WrnMUvaw66nP5FNeEMJ1+O5IBjL8nrNxLbqvuf
Mqd6cJ78HUW/CQXlexCmmzRrMGgvq6/M/WM8AHBjT0NYW7DSfGzJUaiXm99FDMpw
JE7MAM2xckoddrUUYmY9mBzixXAlJO1EejS4ZV2XwsY3i88ojakEPHUfqopBrhB7
wGfJJXIIyXzkhlVu70UZwh1tnlo7uuuswQklZ1Ja0qGqy5prcANG/azY1Bimk7Oo
ibUOcICsyRHGg6WiXvZnIsQ0NibUHdGHSHtO9aZH4PbEuu6Rfy3HYvK3cOxohaLy
5ttj30Db2qKURsPk4SyUz5WMWdn7MsCqAFC5ICsfXm/PUU29UbBi7Ipra2JP5OGJ
HQEJOtQ2UH4oSXNGIyw6w6c9bMhdu2l65UwRtH8Lhz0nhcVT/vRXpEzTxruJNQVE
P0GvaezE3nckEDQHshdl4UoiBk8WOYCHsKR7RJyTv8wPIb3YriOSN7gz7/kFaJ8q
8c5qDA/vvSWavjXW8RSuY08srJhtSJb82slHHu2UrRtTZqSMrxU6Jzpi5/EE+c08
UQ+IyyXHchEP7FXC6FWA6aZJymIXgseLaLTAEnsEbTGsAD3hE5rwvjOOqMFS5Lam
wAaEVh+39MeswB7iC1AqaCv4TTRPTwj3sF3TZqC50m5U/r/CwpXSN7EpF45ljp/m
UP2TvelmzTwm5joKs96AMfxG4dUDe2sbXwEXMmVq6CZMmYRf+SiOL7z0He6pYkI0
lL6dahRP3+ZGaKBGMvnCKFb7U7ElqMOR0qBz+9+W72p4v0RQjWtFYag1Zucql61C
1GTW4vDY901gGAIp17LQc5h43s15IjX/2q+X9IdSEhE2T1rsgzwVTgCDHiGVnknw
8Iw77JDmM+QUwA4iD3s71r9v+8FPCEQfNMw9RGnUHze8VkON7eQPuz43psVQSPxU
MVAcVBWajhJvkNPfG9E0xfQpKL4tiMmvJtunX10Xs2PDbEqNs2bF21alyKzO40o8
kq+pSUGbn0uZw70XcrMitrrPTMc1Vhh+GqWHxjlWOH5xm4ZMouB4rux3uLFGkvHM
9M4D9q1suqbjz6XLIvLfazHnIv9iXRQPxrtJdTTbFIhvpK/8cjgYrCJWrpw5b965
YmqR6R8FK/Fd75ZJXloouUIbf+Yk360ubev0UO5adggIRMWipCIpWXcvFYgxDVju
+dGh7Y5aXFtfDyabgFkt8+4xad1pXdjEOJHgViEOSfIA/3oZ2UcZ0rniZ++rtMhA
0r4PZvn7RXGpfe9uzl7TFF1Qzr1g3BLckc1s4ZEL9cDZYKBdTDm+AQtDbHt2pSEk
o4db8GScYtokEjbrl+mS83AUsBGaL+cRYdMHv62SHYO8uLeaoZ8tQ3kRZIJUmXPt
1ffWRUsoO78cr744KzHOHDzFuNYLFLRwhDO/0i5EPAcuHpNkDc3tHRi3gU3MeWVE
pB15geuXfJVFhXsF1bez5QYglqZXzc94q/1qlEl4Yx1Smf8Td5mcjzpFDEIDxW63
C1+FPvXVZUIXFNkleak2jhPG1IMT6Dt0SN60f3rudf4Y3iQYKw8IIW+uIss8y8OE
cAZHRAnfIcMytuNfE4ueOsLwEbkLMyCa9Ti/4CGIqFLG8MmYRb5ONcng2lHBr0jy
N3G0i40hnEvdiXm0QY2vqxdW+OwG0CsbL7VJhIsUJPQVNoJiiowzW6imgi0mHne+
xAj0ocHfQsK0FQwR/5NnykSxwV6lBoJlaHPbhZ6Q5P+nv8pHMHUGKOwYW7e3PBLJ
7xHzvJR22l6BS6BMH3RKQb+YlcdgBJ+4UA6VBolaT3fe7dttuQ2TwNG8JO2uG+Ju
8rLSnrCt4E2PBFG9srNlyLDNQz+Naco7G4LRHWrQECdF90ocEpTMUGhVNStd0IYu
+T2jw9eEOUPb+qV9EyL8lN6SMaUvRDtDuI3jf+GKYd+YLcqF2E6kKBW/YNL7xKMW
24hyJMbK47/+kF92/DqfXy2zhKphUlMAi8d38lV3hF4eWLI6wn7v55TsTu5QhMEp
Pi5aZB5qDztOegHuhB73t3s24j60IthmNA1lZUViwZEExNxzb/GAh/AhuLDGqXpi
UvxIU4Cv9O/p3DltQco0CVOBcBx7pb4G9SQ9zhoqCvuTC6ifFsoONXUdp8Ssa0fo
L6Iette49GEv8CgSPxb/Tu6+c4iWH+pC5pYZzstB55ZtCaxRbz7Hurs2ym88cP2I
TFjs0tPRhIZJuACB9WYefzZXG4jR8c9TISdTHfritoCR4xlsB+iSJFM4JZUQ4jcl
IKiYoYnnck4kK/DkGmUFrHXVvat5uQhOfleXr+DNDeDN06s+NrJrrxq8WEMKW+ke
fP/PRWTcvlBuc9qIXw6f7hWaSjcvFeCH7WjX71G77h4PV2t/QMAurgUebz5d3TrA
Aovu8ktfzYZVUdDyvnGK1mTyug2/vpF08H3Qu/8lAbPYDkvZIXfkyOL0fbN83zvU
hsRlXonzkPRdzR558BAy9FuUXqkwWUzS9rdP4QvgDPl3vqmpZbIobV2RnnxLZq9m
4RJ0n9Hfk6/5VTNqDskYf22U/6RRvdJnCrrc9pRuc30WxZosUYM8HOAL2UglnhXA
88k5hDFVDD2hK3stUu+DW2/w/gN5FGczvhBhfr1lXAZ60EFTH+mHh+aq1zZ+TdhP
1cATE/Q7kxXhsz+SIMRU9mMDAfhCJM5zpQHAkArcO/b85x5OjoSJ1R0ikXQWgjxa
4/L5CSAPLJWFHiZ2n2xFIcgEnQosyFiQi/pAoJYkvQIeoyZwk+fyAkOEjnzwhZW8
vP7mQDM8hdEZVQho7hunGZnroQBspTdjchETELCo6NIm8Sna2RkO6oxgerOBDF9L
Sqc/vglamtj9Eqihrzr/2SYlO7JEJcCbVwVCCv5NdrU1ehZpZNiaJos/c+p7rNhP
9Z1WTLEhwoxkUd7DnNOGLJ1xKb9WH5SKPJ+PbvjcA9iAHFkg6llOKvKhWteVbkLX
CIkewme4YlnnGGPXLbGHLQrvsZsKL6P7jV3jSF0Kf/C9dpKvrtl5J2IF72zBZ/oD
dcvRuAYdHYMle8rtP/DbnrsSsGJklmx++wTDN35bcoaehrMm7ZwpJl5lUblCpMNW
xRsqflSgcdaaxjSzsUDb/hQAFpQRQBWKUm5q/HBlXQTEa8nQBudMjK4H6sAl/5yn
WeeaO41/yFwRBnNhxPTDu5DckXfB3xUw3WvNo0EBwtN6lXWyoS8b1gDB6NsN4Vth
Rwrh6m1o18jWhSnQY8KRvCfkCl3VI15muMIoPe2+glkk5xOrcOfUQHUUpFfoHYUj
oS+4fCtrEVRbyWKVpVbdbYON+O8CKeFwv1qdha5MAUN2t3zyDkFmAhWClWvpZFcC
q/0u697n13U4KvVq5pouAU7q2yCmPBVg5t/poxqDyHWUtMle7JumSYF3J1ADFGJ6
Rdk/yOaHCGlRNsA8s5mqRH6jT0Mwq/3aBacus3I7QfBsQf1wB7SWJwZDqLbaOPKL
fL1g+4ZSoW8/U+nyiiN9LUtOcXId50V9wZBMxiYfhfDwc4DwMjfdJpPDsMYLC8ri
QPMVDfm2JPLwgu1L6mXP2wBl5J5KMz9HV6WgpLmpak7qtQyC7iTJF/i1fRqirao3
GPa4w11r7eIgcVfjMaRP6W8D3NbW44qrtwT5xQBbKkcb+3hjA7PDVOmwuGrYnn2U
whhN4oPbHHaCdn7dAvhbf6FAWltus7KCWueEZAx6R0sS9HPHUHLyspc8Z65Or3tO
YKVMjx1WfneeTQcBeSgDA7uzTGEURntTk5rjVtObXRe+MdsizPG1nv+HCadp19xT
1YJPpjIATIxb+Z/rHS9n8iP2g1yH4HHt26uXBCIaeUZ+bfHHwFS66OJyyQPgo56N
TMz88AO98uScQ23OXNNgWwdSuYBUxfmQ+4HJd36Qr3aXCirq8/2dkaDWjM2WWP8x
UvOhbqYBxLk+sgxM5OhB6zh289whSgHn2KBX1ogxAPkeP3JrT0RQwkGf2X3Juo8z
tic7FYJKpX0hKJNNm8stotSboRWs2HQtOamqH+vahegf9BCo4Az7JrAdvQ8ZY2VT
0qs5YIqo3jXHGmrbM4jsR0cx8iyMMxhZZg6PsDbIoDnKLbOXywtNGkvCPXGjhAHE
fYeiGBnZhhXL7OND6vFTCNo8eVIrWC/8KOoHyGoly42+ReSjQQlv/X05nTSS3EzW
/RxfAt+u6QD9ecdHzXCt4g24LQxwNPbMX91JFZcHoBfirKU6V1f83OxyhQVZQmoP
e9w8GtpsquidWhS7seiQNRNdBjrDESWegdjGkzZ5nkXue14J+5BKHprpp6wsGZ8p
JJBgDWfAfMPoBlXwBsHUUrs6ROSp6tS84ezAWt31Ha6ZqnvSpxxevz26laDyRD+s
h2LQ4bcusmHu5RfdjNs8VISKXDAOJA1WIr2dFYqDTmx881+bNMDD9cpE2WjzzIVL
vGWi5GJh03IKAqeZkoxt5utdNJCq+60rexyl44LBIZO3C8VOWfiOPEBheu5gMEnm
hKCs/12QeswcWqEDTeQUhbTAz2Ba/5DCtbaCmP203B/+3w+6OZgoNZZ5fgisykvE
7C7CelqIiTsK0SyQKdhUy2RL2yGKrZs0VOtQmiXS+rdx9XSTZDArP5KKj+jYgq+/
k+7PAQcpoIdMIvmnk6EXUvwJ3pdxwhHTxsQVD0Y2dvFNV5EDu1lnw3xi0pnurOHG
5WDx4M3t8n8wtMg73955O0xNTbdrulo5aOz1jw4U/mPwVXvcbPseuT/vqFoavOkJ
LHKKsnjnSWieWn1IjyfRBKvBdtm8jqXL3uGEWzJWf//X4LgbYtrFXNcxRxIxT40M
qnxdRMqqc72AW0x6VtxHgPmpf6Q5zutgRDlDFqOebOk3IiMAtliV4CplkFJw4O2F
oHrc3G80XswPhyrXJFiRbnIpi9f8hUkKqO3QXSnL/2PoxqaqO/v9fjB00sCh6EhG
SkTwgWXvsk7sveHsuFpd+DTDid3vV7imReGO6WMMa2lr3ZW3xnfsIFq5xSm3ImAH
V6n5unnCkkfqXj82l8DdN996eHgHAH77HMN8K9cur+eX2DuEaHl9mSX7uw8YVzyc
BtGgB4HnJpuxeyTRxSqXJNIBVG2KVemsPT/SJSv17gCNUjfk1k9cYiw78Fjq2dhp
CF6sVJOdYAkXmzr+llHLAvySjkH0eq9k4P/p+6PdAzbT4gn3HyQ3yD3jp1ClgRXe
sKpvkrV0q9KkwijuFNlPoohPrI7kibJPaGnIT/dwaV2rb6ZOrH5HltJhV/ZMJMsT
ThO3vz6Il8x5Zc/Wr1Nn0WbHwQTObKJbhjjgMWlB88yWrxc1KBOVu/71EIFi4iSR
UYsK6dyrEf/Nxuy8cdAac3Usd5ItFyf+f8pjQis8wn4Vqt14OY4/AFZFJnACjdiq
If5S8zqnLWUeJNT3cWS35lYJWzmBWzZxmtgvLRj9kikIqt91xSouqW83wLl1xIjo
GIOsJGHHq7GfS3UC21zsm+yCg/VB+BR+kLE+Td/Mwt7YtqmtI2dhM4fn9RzU+pSk
zJgdIf5mNeRRjsme8Y2e7gdgSszeyrU5jDlhdczCFo4sw8VMqcQnXd52w074vjlC
Ku1BVrQFLMS8l7dtbNE4/GI56+ssWJOUwh2ZaRInHeAGXFiT2vg9hK+mCPdaZ2uz
zHa5RsgVDxMzol9DDcxWm7mfSJlhk8SszaXRd0SC51rPHi5oDSZBIkbpt+N++V5J
UVUVnyqrJGiinVboP6za9SayxnmDjp1GauXTn99qWxibNWtT1AmUprmg8XB3WUqQ
7hD/DxJuNsHv7A74NfNpkLQz41Xn0JCiXeDWnV5JN8sFPNa9n+5DIA7+TkXNefF4
ZYSrHYHdUDVMFumPbci8Xry3NrgxN2qCNwNz6neB3ACJ7mAxHjuTjo1hb4JiQjjo
WQFVq/JqrghrfsAvLAXQAdW3vG1GerZGPWW3t/4BSW1f9nHy92uNmACDFoYAiJh/
jZgAxIEOOSif4EN8IQY5lRc6wDdFIuH5QuF2EW5sQQy7DjAoHMKpp48UGLLLgh+m
QU1Q5/w5QGngjI/PvJjfLalIRwq2lzZOvTDd4grcM6zNRcXAd7mdUX5uRpqtu+PL
hFHtSyCPpUulT/hEu0h6WNTrLVVzBUNba8GVc1ajQzaFyLV1KOhvIALWjI3/fbqF
UUhbDQ8TrRqCmOvmroA4LKzNpNcuqpmdL11A7gGkmDR+rZOeF4SEJgykuDzXr5mD
/0qCxuUPRhBYU0YCifjOz+kzT6HVf8L2bCUzmUgC1uRegv8swLyHN4f0yBLsFA+9
BOj9xczpByh0JC7ZMcy6GBs2e8yMw7UGmomk3wUIq93wkI/UlELhW5XpRawC4409
Pr5FkelhDOJLeqWn1Bxo/mbFKpUfpau1WH3gcOpXduCnDodhAF0SxVGEMLU5TW8L
/z06wG90sZFq9QussCNoWv3h10f4u9FJaeh19FPrerTvyZzyR4rbe7gDqL4yp8wC
DwjV3i0Oocz11myXJ7mBfFRbziauKgiOSMS70Yr467sE4Prt04yh2O99hDWSefXh
2Q3H+yGRvRCiC6JqIR6W1+g4u9CnFvVjfdw+rdRZC8vjjMV4REcLIlUvuZm2O4dg
tLZ3rDg+0jR2tUff+sWsgRtLFaoOAkX3pe52M/m8FPAw9XFYSh7ELFgp+oS/Ysq2
qjif+koek2uSTdAk9BYJBj6Vb1DyY3Fcr1ahOejse23pVQq59WhVToDUu9pS8rDv
Hf8I3UBbBMh/JqdgP4QEek5Q4A+UaB7Fr/yshe/Jm4Lo+EjYV+G2CE4HClrX701j
lsKnk0XWjQ/3MsSyCXyGQKaBO1xBExZH60yfsaqyJzWRe2Pp6dzRj7FkIfUQvCdp
2D3OUdBZPpFctco9y9OLBlI3/wq/F+Qi5UsurW3wLf23OzSQEiuT5POgfhVtNzqR
cxla3ryX7nfRHajA8hYrqyG1Twq9/fMWOy6nVF+5xPEYViogr74McNiDE8HG0m4j
RXU9nTNe43gX20zb4sqq3f10MNHG6v8WkDoSwG8elRVRcwvAxkpV3eKUaKHq7y7c
xmut9v78FO+wKNIculwnLltMRfgAIB8nL1lv2XpRtSKHlp1BSxsvSRr00BgNX7/n
NqcWkgsbcg/xVT3N0dg5I8E/b7p3GYy0VLDFlsN+7d566sJTjGIg6SoD5bYrysVw
SyUhO+hHRo9oTj0miKlIIG/nMyFzoDkB6uEgqoHl+Po2I9BIQklW7XkOeqF4FPNs
YYMg0hY9BIcDZ0So6YO6lpLFcTWDMgIwByNi/W5diaZjYUUlrduYE6dLsEGFTKGY
qEQE75eIVFrFOs38xqWaLhE7+aA8QDWHhcfOra7A35+WQ++Z/8YBoT6KAE2zzV+r
G/fjPcPuiKrGM2uSA9Rd34ZyxYbfI8cbAWjj3f9DMv9Drgnl862SpL0QiIaG8WWE
FpWROeDbQJ4P/bHk0lbsXSjDdQNucqDKX5sUMRAB0Kjf8g/yAPMeiAt7WblbuUQg
GZLx+peCoaTya45hiJPSCX4P38VPV/sIVaOOV26QVlA7iMlWNN0ScubjScmlDOdT
ZDmcz5VNKBHuXaCNwYRUPbYF9FuzNfuMMbIRsrkf1TaxWL5H3SuCz38CkaGUig7n
uk9DoGhayDjkPi3KnmHc/n7DtkancadabH/TnIzXaam7ZMJhhppqQgmVYGSgEcKd
sFhr+nihx46Cwo2PztQ410REciteKQb41xXvIW5QQHn3ifH7Vznyor+mRXA5gUMH
zwmdN88BuiTyA5zTNELojVSRxsTWYwa89kqsRh2zaNUErzos7w4uikYV44pXrA/K
HMyIrxQNGuD7KRN+OgQVMtuDeVYy9wgM6N2M9mqmGhwgeyBPBnnN9d/zm53Y1lWN
YrabxnPk43M+mTZVqC7Si+1pS8Kiyx5QZ8GTEPkcIoMqjSxYb4jJhFZWyfRBpL0O
2gOibDwBmlWvIMkSl3Vc2K2tjD+OeXJWLz1B5M7YJN3Y2wQ8D4ZIWoKsZ1REmYhH
hyG13ukhSF94a7D5P3gKZh5RaxasCBbAsAc/A9e9YQav38Op60rkX5X2Yul4goAK
0Jm7LpJBLVyExHiSM5rAxiJAuswmdgWNYsXLetmNAJ0OiHJ+bbgXBsI+ahTPe0Dd
lUKR4aMkNz4cYj3uBvdk8O+Rz1TdO4Brp1w6SozD7wm0sLlt6eRDO2AJZ3rsgtUd
gpCE3IdxmBYqi1NI9G/RCprnuN3RHHlA/xszY54+Z86URSvTSTnMP5PaXaNaysMa
tSCd90UcJTczDmtCKlAfgJ5Gj/i2+oARO7Sbijcrp1wYyno/IdvlUSM/4XgPseRo
8uR1ExqHq1E/1w4RTWbW5KDlzyqhbj9l+CFxFdnUYKZl9mhzRkzu29ShRviyq2QA
tF7jes1GVBha/WlW+ze4VxycMGNJLfO+gkjD/mEpXZfXt1hMfHMsGewQXkhABc8Z
HirPQLpHqtqURE9VFJ7MzC4xtmCKVWOCWObanzPty4B01pAPcU0NmAGMU2dq/D+c
460wpWTxlhnsFZwrEFg2xyk+KuORbfPhoTUxow2OJ/dPo3J3EbICn4oNvjTru5U9
d2Y9zWQwnnNHNr5lCtiAd1RlcBh6aTRvApYWuSUTm8j5gjf+YvdprMRCVaYr8JB8
Wp5CLU/poObZwW2+DK2r4jDyk0EBWiv/RI2CSbFiIgRfGpu8G9La4O5LmNdCluB8
MjiwixPEwYzQkicYSlvDVvAoeyouNeDPqH97MadEeswvgvr809rOusT+Yxq1ef1O
saTxu9Lv8CsfxI1249obWasqdIhmDymyeQqC6NJAxpkdGf49YkardiyOhsu+xKxp
7McsgtaC0puL5jikJsHdxQRDRkwlbsYW/M1TedbjMZ5GnIwBpKjis0dkjS6CH2lK
bMq5if27uVWaEYwfBKm2o6WzIMgHIe/DgP9mcJKGFLJbH0x9Qdlm7vaNvFljl+nx
ryHsdXIxkG9DRZtELU/1d8TGviRp8y0ttrRbeB3Th2kKjmOdpMvtKS/9XUvxGizZ
DU+Li5lgLmgCC+2lEI3tfwf9NCIfnLEp/gh2G8wv1j9jUtK45S+1QaVuDdIJUSpZ
d0b6SOAJgQnOcSOV4rRQsrIM4nTSEiYusvlFlg28jSnlByOrBMhRXQvt7tyeW6h6
vypztNTvjpQQANxZwXZTKizBT/0oOXwTcwK8XOI1+eVMpvfs7HK+M8EuSXab8e4A
OCCaYp+kJ/jxJTqpx7fL2D81SBfdgAHDNHqXsrdsYLN6iHs+5/137WhfmsWM+Co1
zcaXNux0PCG51XXErRZU4sEgzD0UBbnw6BaGGcmV6WCB8Lequl1uw4wv919LC848
YNrbKnPpkaId6YBHi546pf7T4PdtKFry8VdKYlJQ8bCvyN3lpOKoc499OgTLhbIc
nlZIeYCWApl9l5hhyemyt5264ZjBHt+vPJw7FvpCs8i2W5jiWpJOc4f+rNCnT7Xr
Qrp4Z/2hay+HbOHdKmLIHzfjcusm9TINZPqdngVHVsWvv8lu91LHupfqJusprrSW
+FpqcKfAKqnL2pWUs+bRzOKPs5GouHIOglTlsIiEfVv73nHEXhqyYeutZ2ZCDLhu
1Mify2+CBHjXxyhqm6e7XoITRiv4utJ5q5828QTK/Cmjl05OQBE+xgPrFOnkAU4e
XcDe28YBt6gvL4/SKT5cRWHKo9lVnlLPTuIxWNoGmiUYqhaVJUfEQIFJ+aAhKur8
Dksim62Tv/KOGQg+VPYn8rm0C9q2Yf3r36Jmf16nDD4oiYy9IM2k4muhc7wR9e+z
2AfhOOlEWfH62t5OZ/usZpbokqPTD9j0aGajfR+9KOJi8pAa5mS20jFX+qpnZd+2
kqTVDrcAIrmsWIpoIA5/iAFuIRfwIUXZXQFnWH613wDrWU4sn9rqcM8mU/KafHkP
CdwD3KZfVsFu25aaZM6G+BPQvXD0GiTp88dLtt7t0popGZquQZjpOKa6Xb0GnY2L
idDutU8xsoQgJoOZwSCJdTO37LYI1QJTjom/HCb8tZTVvLgHiz3xo830XcIU/UaT
ZVnePw/QivOJ8TN/JWkYUDcjWYqh3zEK71BmfknVmh7e2w9z7jgUGNFZc1gWRn1d
Ljuoh/psajHvOe4ZnX8YsJbqt9UDmdTQq84tywMimqAdo+mgLLsID5HRTQrZkKiR
/5hqnxcXHWLvImb5fGLEhIMYw1uy5IeyZjVTN8Z6BH5LGVx26Wkq+83Pe2d/FKaP
0VyvFceLWTa1H0CYr7bl4X5WTK/aI0Lk4uuB1Xu18T+IDPWBzJ8uitbWmJJlAoVa
yszZbyxdyIWkMkQ1t3rK5C3hXIiHcrmOrCaPxZuBhY8XmXHLXzrKXEXyIAss4D+w
3ry1m6iOdNOIvEH58ejzarPV2yhoCeRwlSvcDmHVymKmmsXQ0HYVaF8TU7IzqLOg
FE+/SUWWLqo27ihwmIOX1G8P80AH7mNeHPPwszoda20YyrqhNR6VW1i3kf+PnuVt
/nmWzD4hZAFdXHvIe7EGgMewPIPKE/fggx/wWmV204A+yZcEam5pYUqbUAT/H6Tw
pJq1XUxA0d3ptaE1ri/v/QPWkhW9fzVVOQzwa9yeOgucWsRVfa8USP+ub3PbRd+G
CPYf0T3Cs5tehGBa7xGGHEuvfp6PvmoGjqAL0rHme35d3N66yC4EN7ES4cstM7P0
gk/tUGCzPPchPnd0tsPLHV7X82C4/7DEOntr5NDxB0SGO0DP2BVXR6xtrnKUitkU
HYHoob19iEx6UbJU4bDEyG9BrWdRf5bKg2rxqv1YJyE84W/JGvIZ7c7W3KzOENOi
ozMVAIJuvEel2VUYBUL7eAX6P4YCAUYv6fAfBDV6wYCVnnHj4Z0VgSKAQWoA30/W
1rnLHE+K3MNPx461lYL158XhOOGONZPb2H+s2hQqz68JS7BbE43FHccMZPUWTZ1x
PeqnkRav5/aWAS1Y1uRjc3UIwau27FRlbLuBtX0nC7hEkU1Bha36r/uny/u7NhrH
I8M+Ndwhm2NvwqowO9mjlNEAtETOymBMn3v/z8s8CLYIhVDqIheRTNSjZ34uI08q
0g8aM4uvXNrDlPySVvC7J/iI31kV9IuDDEO+EalIRc7ElnxMnyrmiZbJ36lICP1+
nNWTgh5g0GeqE5nqse7RTPVMqssRBj/UVC2NBz39Bmx1y22yIVPV54LQ7Xby/5RD
MUF8WqgtaHMRgJrQ02eVeJU5puJgzqC0d0A8L/Vy9e3NInbAIFsq5ddtKlr+kiEl
RIeSDJeyDjJcXtqV6HdmcNrB1Djb7odkI72vLJ/VybFwoLStdbnYOn/yqrpHCYSS
Z2xTtuqkA+jmzVLoaf1IRRwH6dooiULyG8y6TFq4WvoW2Cz3chIFDWoBEaZs37Mo
y2tPawiE2G/hESvza7bryrAzD+lR+q1W8d6FYRPQXhQePtO0hsAVnfr+Rs9dhJbU
F7cJwFrkdVBpUy3IMenmKSk/1sllIAIq4hsX+LjKHNW2f5ai/Sued20ja3oK4/o4
nZ5/M2WqI8TmqZZ7sElYSIP5VUWFnwOzvkPQWpK/QJQcCyF04vi3xLzmHjzXn0dG
j+2qwv3jCk5Y7s26sBZhbZyL82izUzWqdyRsXDBFX3KCsPDrG9sdUoOh5T8rOj10
2SzIqpdMXLZdXTHqgYdMY1HAhqIeaL8QGBGZfMocxSvEVvZV+OxU9E6Hfl2L4A7U
Sx2rOKl7VgyVODz8AysxXKMn9Rp3DvCW+bib8prtYDJlR5tf1XmE+Lo2Z9HSHGiK
ncySu0LRwAj5udoZ+/7lUfE3LBY71pVus+t5OrRKo7DLitKlxc7EeIxFnXy0R+42
563pImk9MOLD0j/JQKTxNSySPnUH9+r83AAmOnRNuEH8z4NFvHdx08ERSl4LADl1
qWLHEUHL0RujNKEo6gANoXNVeXkGSci13dKMbsgP/LI7B1HKrE+hApjM8XUsK6tQ
/Z5+3KdhMWQejYpvbELViJmiPzr2OJtHWfLqo8XvwmFXF5gYWaO7mEVcLw1MKLr5
pMWhW5yCoOzOrHB9Wu4cpvb1Au38yY50XHbcxGi0Oc8KyL+EOVaT5rkGk5wKJbbu
8x5HxQLvULiqeVsGacpibOkNfvo8MK1T9PzvPvbObdBm5fDYUsKOEdhAhgRcs0Df
pSCloH6mJG1akL528M0dB8e9nJ7g6RESQItt6yUW+aZJq/uBxnYu0/a5yQbhOmLb
Uq2JJdHZ4xqDN14+vW/GyVi96aW/A8KJMUeHn+qfr97sDheacO/2gBhKofyh9zSn
hZDgZW/cvkFNpTNLeiwTYkr24IutvQTYJjduS2djMXL9c8voBdKRgu33pBBbEoEz
4iFuQiFuGixT4+uP9lqi7CYeySOf9F0HwdLlSdnyl9AE9RBjSfzY+IzbwJK5S56p
hDaw0dYJSeRSTiYuHhTV41pVMs0BZhGcctCgIHooRoatf+VLHXRwb6w65sH97At0
3vnRUpkxpVecGZ80XpGETmLYgLu976FAnl+KWMrhvc330/jr9Kn9pD/qD2YMsuly
2mS0yKjA363an9iOVW2SzK61gVEJLbFg1GUCL5D8c8OOY2XLI6Rl5jz5uemmvrto
DCAPT9WrXJE+LCwF0BGsb18bT06gNorWGKoRLUt/g7S7uIe+HRYwWNUJplJ98V7L
MeUm/ZBxuRGBURqlug89cFf8i8MZglHo+0SbbEvrBiH5yoANL+Q4pJiXlfppPTHb
L6A6IzDRPP7CBc140j+aRIAU31VbYCsSgG9ZOmuYcJGgB4XMG7m/Kdm/090gghU1
juRyG4QMcErntrPxWH5Q2mA4Hjf26S51TMNAbRyMJp9q4XCh28NUVTXl0MpKWPeP
SPTLvcJDC8aHIkvOd4e9X2T3wf+/Uu0UOYsBzYjNrmp7NcK8i7Lyw6zTo7Q2m4wo
/9Ya3JsuvyRngcghaddtsxA44qyisEHrERYtDdCzuD7IGFcWqkHIU1WQ/tpK3d1v
yF3/8DVQmpGzLzg/d1N+pqIUXQti+gMdvaAE8EjViPZ2xBXNcT2ni3NU7KiExenK
DJ9044gmFYsjTF24gwclX0sTC+LycIX4oDAqPBAEY1+2dJTKw5n8JZ2MFcMxu5UP
6TEcZ1idhvamGZnl2eB168571Rqvb+eGu15wqkhhOYGH8LATl5PvN6D2B4lpHBao
e8Y8teijfadAoiaL+5BdA89It34VZV8ifzRVtnZBX5nBgUHoP+OVlVPswoNQQYgs
Y8TI6et62C1Fetv9qsCkBUDJO7mBu5mIFmD3PFX8rUYG8asMpbAW6EXd6d0UQ5JY
gOtvje1BHQ6AY076K4VVrWHUWymBByugiGs1xNpGvLvbC8RBmQzK+tYqoTfhofC8
kJL1uP/rWBDJjUQwtDoswGg38kXUbWsgG09ch8eqm4VBHWPtQv6ewHIOlka30E5G
+0/+JoUZmN8mIKi5eqa306HwDHXHBvhleqduO/Cou7AFpPMzLuvvG63QEx0mnCO6
gPgqfZX9C93FuLVlZjo62BKw+YCu0DHPxQHwiBP52msB/06VbKWoRoFCxQNxLQNV
5oVwkstwpAyuc4D88xezLG1VcxPFImwcs7NsXsmQfz78qS6qSPVTKTuTrjh2Dklo
c4mNo7fUy8bH+jG1PjNEXq9I1qNawjP2TQiTKAgpCuAHlqK9hopO+inc4d+2HNF5
U6jlkTrDQ21vozHmuZArCtZdQhi8+V8cSfrJP2PDJY78Knf5jUoXaUI5ZLBcxP8D
JUNc0jI/riJCbuvXVcsO66aQnuNpQQEKW2rvDRiR0K16MaG7Yt/l3PyAmHPLv/84
rux+ERNdq/bmta0OoGXksHpMQGxN4uNnolKeW2OOma7xlWe1NP+z0a1/D5MQmw10
AS6cVBXSNr5owaDC1ytILTFws3sw7fTmlsDjY12JHYFNYPa4h6ldxN0wnKl7ckg0
IcdVBerioccP96kpi7/jUftNcQYDxHseK+GWWiXZv6zPLgaQEnXFKTaVbXXSa/r+
Heysx8G2f6PPqEwAXNOXdfSmZ42A1uLiWOzle+OdKnADhDvsv7fb932EGOMEgBbb
hpIPZIHbl4Tod773Nyjza8ehs1BSoOh+6/4JJXijMDey+aBSYRwSZp2I9a7zt0M0
0WfxYtQU4YPn5bIEksCmGb4kXuwM62yIzVF30JhmC4GROIYsOT4721tMlrAAhtRG
+TNYo9UTvq5I4rO2WbeOgc/Bz04g0Av5LI0jyJuxapCQdi62PZ4kiD64w8trigNf
4tdAfeKRj9LIJJ/t1df2BD67OYxlU87/pH8U6MAvkjiHXkQhxWr4AtZiefJ5OpLU
y8tel3VfBfsB69RFe8cr47Vmabid1G2KPUpspAIXG12wEEJGbjTrmVLOs7OZyXqQ
qyE2DQCnzDcbHj3Iq7EgUI7130QFMlqnkKD1SwlPyHIc7o4D6wuqp9je4UIWR2Yt
bJFm3135KYGEPWfZrjdUt7sib+ixfQyiq4Y6kfWBhRI9FlS+gjNk7Eztd3vhuw7F
U+2wIxFUUFNwEB9Ckj8JjgZvKJHKST18u7DLN4uSV7D9JS+rNSbSb+z9zZwVBUux
naCwSSTQuG5cTRFwBffg/PsUEkssImGBOaelhJCvg05l76iLgFOyWPnHYCGWmoGC
YWCkIdyVP75WALHuipOMFZ1T5sPtaQ4mbYUnuo5V+cr74l8aP9K2SWM2q+LANPgx
LrzbzW9fvGtfGIVOYS8eXDFAJsHJlel7mhJNLna2iJHOlwdzMc7RIHSQcrzZrqBd
Al+qapnL+nm2UuD0zNfflfddyb68hAltjpBD6mcgBMOwng7QDujxHcGG+qxZ8cRA
6jmOarYIv5j0MNZW3bfDQXiv2qxEKzA3SdDX8vItm3MzawYHypCqtA7vgoCesCZn
A4VHCx9AHH6AyHS3YM6g0LwcmC3LArbZK8GGjDnnYamokWYPTNvMbGZzo/s5xekL
9nR+FCl4757fxgBLrJUk4rnA5V6p0Soz5T8In2M9d6P9LDXTp2fIzYjTAZo1EQ8z
TqBrczcyxPxpe05bMIVYim9VZHdikV9ELj4NxVc8wNOxlwgx6rg2mxklkh253Q8A
1EYhXmgXzmglBxUC0kdiX+wIA4LS/iHoDIOFpSz0lvROFA337+E1c08qGqmNLai3
SfplWQCulydksXDr7TRcsqsgPvl7v5bITUTKVC1Fro3jdeXm8W+f3jQ6DCxyfdYX
pd3aobvj05WBMTHxFqMUHg==
`protect END_PROTECTED
