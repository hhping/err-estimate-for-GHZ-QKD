`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ecaf4YozORKzs3lXYSoPG9CAX38cpaYGmBTpGrGciCQ0pc1Z4Y6e9jokfW12S2Gz
S0uHKEJR9zAHwicLsRSWoKSlSPKRGoIqjNcGZAvKvZxjUhQ40O7ukzagJALDadwS
obaUT4ICRg3hLNo8NmCCMpqItfa9Q9AWzFK7cQFUNFOrOSRJmlhQh0an5RVtiLwZ
NKGnAwpEowQBowDGyZHvWlq6ddB4UtIsxErC9/+rXk++rWzuhwi+z3G0q78Fx3f5
U83hmSxr8WDOQSHacqQKQztd41h0ZDXIB6NSWLkE+BKgDKCL75VQ3Oj0jTCIDe6o
HXO1p4iXN3OBWngPTUjFSW8p0MrkjaCUpvF8BqAxitrbffhy3Eimrw8Tb1ab8Tjb
TSYnHpp+NAN5Wm46HkCtQskpelplDmB5ahjLfz0m3r6xxtEBgBOJbuzN/RzaTcrM
L1Io0jh6IsLzMdYAf2GmEB+SgndMgIsqbB8jHFBoJYcUbCYpeSfNN8aazRaPD8FD
a5AWODi9Y9FobgntYIHcFf9nPTtPfKjHRTq4F8p++BzCAjfUGZWbF4ON28Odigse
/KhK9f4XWMaf2DlsKldAZIjs4u0G9xC2L2neUHl+evF1NNLzeG5jd35Ct1fQdXiw
2k4UFaGa8MsNxgY8EeGK3j2fQibiG2y7SFu8fhCcmbqLiYMr9Zm5P6wPwoSG8zo8
VD7mgok6wdr/HSfhULqm/zGHbES1VQ5fdzwCSPkuv4Hhe/HHM9CY3x6/DKyXesOp
khslJBE2qX8a6hlFWsrUAyLO7wjS3Wxx5x1Ja+bRimlQ+HaxCCTymbQCIj9pbezw
MWLaHEURDtu/njoaryoN8cgaV6rpcHR0CQ1l1c8I1HJMFmOcLXCsG0qI/vM2mgD4
RZlhQWbEeLC4hJIONrTqsxuT6z8kjrd4qMLMojA0QPAW6Zz5RM1f0gim2dkWCn2p
t1E7oBM/0wLZ6z8/T4vIYGGVqh6E76pcjlWsgHdQHFdFN/WbBWywTNBCbWZVG4js
6RG+22yCToMGLSu3pd1BTpOHUGWWQjchj3FugMNJbRLEcZpoDYpcbxpt5Zd4C5Rc
Bia6pnHcc/vqMLv7LLQQf2Di6FNitT+x7nBK4z6tZ8iCyGAUOHXJw31bIj0tSvZw
BtzBD0ntg9NXNFUWbR9VtBMSPlx4GiHWQiQTXM7SBmwKHhkWByFZ+x7oqsT+1m+N
ySp4meIZtlgGEbVgNBpY5DKP1H1Vk614U/jNaXxGV516snNM8NRjxvNqhOkN0th+
sCej1Pi1zOPqlTzlM7wg356cN6wNXUFf9OUd77KyPyJmSt7GKpI9xcJNFSU7Gs7O
KMd4yRIfynf7MpWmy+ZodjbJPjr+DEcdA7D9WvyCPVtBC5dkJgLigBAKv7PdJJVz
Ig7ai/hoGwahtJNzB7qP4Qm2OD40Z49Kcnj8lJAA4rP8wC9aXK++i9VfFK14DXJ1
te51B9VqALlkJBo//xwgQ8AxKDEXv5jCESOxSz3kqOsTZyxCQf0Xj8ZDRftvOukl
PnSwYQrzaFye9hDoCabJBX3S3xYx1gG1D/N3lkLSXibWT7iD3XOeIoxo3/GkcXIh
g6cEEwoUKYyEDsZt77bDu4mFC/OXMhBTIhOI2LqT20X44BSeG8UOpih0Eudy5I9R
E4Boz/cvnJfJndtfmxQe5a5E2alQ4lWdecA064hA7aEQdP+3DaQa1APNOM9MH565
rz/BY9fVUTgHLy56qgq9mygndAdttUTQqQ3vRinwPLAyJTcNyU+AbtWrt3mVzALO
xo8tpjwaP4UvToJxtPStRczISibgi4NHoTdsDdfEkA6soE3Pkz5pQl5Qc1z7ahtF
MikZUPvH/fZaZCIjgxT1NXyWKpYyTavP0Bakty1pyDzSa5QGkzPpy11YToMkojF0
Txp4oPfcHPCdzLBbka3gnaUr/ietLWBYQtiyoUnDoW2n3LbzT6KtPYY6pHCTI/ho
Aj9g/mHTyF7o9MN+OiLukM2nX+grtLh6z+pihQhoAgP6L/JkXXpXzYiUOcw1Kmux
WZmy6dirChtImlUDBi+/Kg++1ToXE2W3jdrgGAO0tFkhRYbyHUgx1CCgCqGS9fGS
JmpAnzQYqgWNWcnCAHzoRRtLHIvWypXfmheMb3bnt/Kel3iM7vT9xOc4sjOhvqm1
sO1+1SS+PWRf36gDYlWFwB8EpOZDio0IKS/VJ3jEtlrsJygVlB25V9Za9i+EfbL0
/z/bYauwodFuyKhJ9KbyXWoZ3wuqxfmo1JzQNfusoIQtcwv1wkqWAZQZKPnkI8dX
C0SjJflgluSDMqcAwZWM0MQ4GxvgtYgeL0sgdchngobUNHaq053RauZn9iitKyoa
0TPANXBUH6/QPUZCwh8IfWF0lNpX+ngt7RWBjwq4n5YlfZby0Xj5s8tqCwc9ieTA
ZC5vs5ofChp2U2FH7ViAeEAomEIGSjlu28m57p040R7LbvakP1FbhUc+PuIhJ4b/
HkGExdH57HUDWp/UODtoTqzLSWsOsGSV3ELy79mbQn4ENML/rxobkwPQjukp3IMi
44cs3/v2oJOBPPt/TiEw8QC6tQi3aGNni+NwhOc0KqoZmwCOMLzIEeTeUWbXxybF
asyWsEwoLo5DN5oiz4ODnEEw7R4iQu1/KkZu3MHyBmFxnBu+ocZC93Xy1CREKxIw
SysDYCI8nWTXCzODhhDuH0VatIT1CGlc1InmEKv4vBH+zrfHlYE82VQXd+dqm1DF
9bsyjGnVCdOuF/E060S4kyOMhxLVMlt4gHq9UsLo3x0=
`protect END_PROTECTED
