`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q+PuVDzr4hkxjEvifAXHlP+t7v/icnHje04hQ5BoT0bX9BtdcRbTEg5okYFg1fch
eh+wU6M3cSVF+x1Nbj81VhOCuEpe/mRrbmiu+8vq1VKWvkZJFWrWWS4IJRP0zdFE
ym4ajD23bmVtzm8SRtyzyi0Vq7L7CjM8JXEd9iP4oTm89rakQra/oTPqRET/w3Ds
mymPOxlLKN1uZshIL1BnQ3pNbgcZYe8SoOfmNBXfLkVJbAFqWEikJb7tWOb2obK4
Oi4Zgt2079Ix9pH3KKhZ932giCzO5T4OA/+ntnzgzAuRXXY15G5ausbDn1PAUWDg
qnkonoqOb+AnwmB/LKohKB4gxAOCJC5owHDZwF3bZzK6ggo1eIMFq7lJXUqaCKqa
4iKhyrOK8gMst2ahne5KHwkWIIZD2HPZ+/1b6yJWDKV3Gex+YopUAIttq0omWyA7
aMaYgM/KqHLejvNhBmipfQicuchUvzDyxQqkl6NK4FmHZW/fpV7uBLfJojknZZWE
HnMMK3XKXRVsYDBbKykLJJjFJ0ABIi5rdzAMXR/eFvEqPzTrazt2CfjNLWcKLpNd
OIg9WLFGhbln6OfTiVNL04anq6i7122q7VnBXoSqfhYSy1pI4GqV4ttAAoUjkHF5
tsjtMofVSsFUF7VI8tBlbkxmgrBxmKTFUsjd6rYPWAi5rHTlzoknSqsnopeTiMyo
Ofns3UxpT8f/9SljtITZTpaB+8a0IXCKRxQqiL4T/9kmy2N8+re6R3ZS/RSW9SA6
qQoRy31y4Wyl1kHHbrdxWy3+XOeD3S49h9jyFE7cmVSV0xA5QhtYwegMIZHw9LTY
`protect END_PROTECTED
