`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dRzVUCgTSskz6YkVyDJvsLqBEv+EGxERlvdLfmOTfytQqiw+SNlpxrRlN0auCkJJ
Nm5K1ZyQr+EaTf+3bqDn0VMtJSDNdLTUIedgGcZuVvpAXR6NgMDTzk0nYaKYykgJ
b58ADT2iSeqjKyEdHc5P3leEAveLArG4DQmk/M1g4WO/swCFCJPNmuhy0DNbH7dR
Am26JGWX1GkDFQJmch0CyiLD6x49RlZLKbSlUJHA+nl16yXyXhwb2zwN2QTs3Zk8
zc846tiTsTOy1KCD9kD5+PuSgp+EUGmJh0cfFn7h81Qr2L4CKym+6jovsSB5ekBF
HVio3TTCXM08xgOODIjRrk5gdvduCKvmB1hAs2PiuwuDowYtab4pMiQIYbPwAZVf
DsobscFbQn8v3QBe8X94MkrduGle7CztQhfS1bJCUInzMaVwCwlRmh80kvJo+55E
D7BHXX96YsapDy/edXtsicgRHzx98PTMTbivcAd4zxkMtpO1wAVPAe9KD/ev1Leq
j5XtkKCqfRrShA/wafMCQVyw1/VLi0Hf2DQY/Gq6QKKN/wVRXX9betxn5oHbAjz2
KCixLAtmtVSMLGoSB/K8fpgDuDdY5lCuWr6h5TvdqIzFifPnutS/FKliKC1OAhXu
8xnfTT50WageBKbpslohZeHMEJuu+so++eKgB7lf8kObN8Prcdnnxl+EKb3dHctF
mUNF6XUIuq4rSMxk7tcJmQ3aBeb+qVA5XxcSdGn6C/P6ByY8i8YRQAgYCVqWKXTI
`protect END_PROTECTED
