`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
42GAwhtgBOGgWHR3ExzKMdSKfmIzB47tHqwmUqDs8fM64aKyXZ5f2BlOeYmRxQsV
niaRov9lrD/5keBRQ62/3ZkkVZajTVX/U1OzkcQp3YMOCX5Ua6lmbqVfsgDkcJMO
5a4UBUFSg101P98JEulC5AlnK+h3M+/969hXFY13VklOu0FJazin/cShCfWlg9Ez
kNAamQpzMEv5hwAXyJdHbbb2VQIXqlgOvhOylpvghHjZJJPSZNusATE8FpM0xhej
SGSIgtzXSUQtpqfSP3d0u0R62jQo6g92oWPkmVz+heL9raCGYwLO0dUtlT4syQ1l
fzPTPZK4fpzK+oB5JxePIzO1ZBouBGxaCkltoXDfU/dFWEWUSzwKV5NIypGNCpVG
J3IzrXb4ih16JCMI1c321YVLNgcz7sWFG0CGtXjAX9Ccf01ZJ2ASeVciO0C7Qn1k
IhLWKlupp0pMU9UMOfDGmF6KugqVL+OfDZtpfi7PChSGxzQq5EczU+1N+ZDMZ30z
5OQJ4G6zZVdmJyp7a9j8M6v8TgfWzTbRxajwtnJWGabupzDRSnzrm++cfJAt/Kg9
nuB32UBlElqVgWn+mueSRFPVePiK2aoQtob88BYslSpthVSGqsGiWfPeBNHCaLYw
1nD34GvGGKpOOBJlgH+OocIaKIpW+kcSP7ff6/IUgnLT3UdXHMgIvtGUe96P3Pq3
iRvqL/tguQkB4tuD1NLQOEdc2Q/tTwN2WY2yh7sCDvaTXsB5bZfjFs0HrYFoJCIc
eoDtBvbNA9dd3p0nH/JwtgHa0A7ZU9qJPLH3rPUlAvpe/+toht8GkHo5nCNwcjNv
NxNd84Zi/wDnNSmb2RsNTVoPfaZHNTrjzzTSvQkRq+T81J7sFAnIAeoc0KcaazHV
HT5J5nFI1I5I4cs+KhC+3P19yZrktQ6Ch4MP+0cTK3glKyVT/3d78F8tSYgDPvId
`protect END_PROTECTED
