`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vi939m6f3PQSHMuFMzg1jjzAuNr/22U3dDxSMTvtGLg5OQKzEABGphNTCB/0LfqC
t7vILxR1BM29xSrNLtbLDxpHgxalEfocpDSfRfGUlpYkECZQOWwQuaYr3GWphukf
z6TapoeLwh1HA8xEglgOXpMaWxWNdXmyScwhVe9uiZfCyZJwfPQRcbi0ifdzTYtL
og3a8CFU+TRTSXWU2O1YnJ2RmzcjL6Fz88VzeGZou7cuRK8YALgPfe0TgkE+C9Lh
VlfQvMia35hI/W40svufbTFSvZR1jUZiHfJhRufWGuSFoFcxwW1DXTEhP/HGDOYz
7Qsn2JNQdVjzbcgfVKIsv4X41PsO60c4Cl2fDeWFTDnmgtMerBZz9qDUZ0D68+p8
mTrcXu3ckbYG4sqXM4c0utUCzbSxC/hCIY0fm2k3XhZdoJqImiV6Px8+Jkg2R8gC
Amwxe1T6M8rnn+2IE9Nw+u1C86ZBPMPYq1EhTuC3bMcBC62aX+SqJ7Rj+EaZMk5b
42GW59OesUFJc3vbiLYT7J16fGd5dwPl7/FKp3bnmAtswCL0gOANUBQFTXWAjdG2
BbzDntiqRSNlLVV59sal5Q==
`protect END_PROTECTED
