`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V60o2sZkKv9LoZ2wJ0tdiXBajen+KdbpVNzkGrDl8Bzu4s+5hXYTJqE9RuL8FMvu
A84oKvdYmssPRaDQ3Bokk1ataz7ZgGLbLcLYzAUJF3te34bIonFMvDhqXP3D8hLB
Y1AM69OR0TpDW59A6aYMJT1ITorLXhlCkT362lH9/m3ZeDH4HNoBaHjWv3fVy2Gy
ZDqzm/YDNOJpxm1i5eBBSYP4Z0uX/P2aoldycbFMpwiWU55yVix3ZGARnLanFsKP
r9N1a1Q2UejNn43R5BoUi4R/ARCd29x4GpJq33Ici95c6uBwvxp1W4jXndMRtG3c
nXmAO43DoQfdNLAPSjhbxuAp8/p9OPiHLp9Bhytnz18NYtEF3Hv97z/EfazW5IRy
ZuMufZirlsQEpN//SQzdcINJKO9hHI1p++FchyWNUx3bw1ge3i+a2M9XiXTHihwi
NTb1KH8iGQ3HJOPov6MvfbusfCAh1xJg+iquM19W6niue5oMX0s6BzBhkbPaSe9W
F1P1p2oT1Bdn5J6YX2sYxOTWMk3TE4UvVTeZSz9xRVR/SkqRLBxKy1JzxSQi1uJ+
`protect END_PROTECTED
