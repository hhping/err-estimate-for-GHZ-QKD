`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LArAbE/C8iMMFe0XVK25pySmSNq/4lj95xmZRk3+TvE0xAXy626Vz3ufK+KZe7pg
RJWHB8fudpv5yOprtiDUIC+eHu1xoacakVsLuHAX4xK0BmQKXkHxM9dXXmyRT4A6
c9xwaHr5ZELLRx09J355iQpnS+gD0J0YMuWdIX8xrmNJmdiQcxHR9zmO+p0754Af
Ioh2IMUrH3PmCAfIzzpVmxd/t0NAz7ICnFpcX8JzZpgTGaqlDNlu7wbfTqQUhBJd
QeFETqZvxJke9AZhEFeEizVy5jNhupGoQbIKZp1BSkOKVM8Q0wo0Fxb8WcPmcB46
NcMaXKLMpSg0BvJC+2LdRRNmfpQS1c/yERvFGiB8zj/vZ+DFBin95DM34VXYeBIA
w0n6vsUFVCr6KmowpqNgW8ourvStsDHwbFr8udGQBF43+dRic+JFReW6L2/xhsud
kToUot7pGLJur7xs6geRlDz9Ou2qa+N006erxh4VeF/979qe+A78KVSTvLcF2jDg
L70ZUVYuo1HIoRQwoilwqRTh5l6lFa/Uso3BZegJrenU/Vz93VUA7fctA/nnt5r4
Iy65BNMFUGsA7/rQK/bVZkIeWwH0SNH3HjbNw2jVtI7gWnyCCsCOxpusawV8jmAS
2/b/CVE0My6HPIparSeq97lIDw06sZNRF2lz/BEynZlsqylXoOFAc+QxUbjrzYKO
Z5IA305SLDb4dHSbyOT5BkvtvwvLnrZYzESdfSKxc69qIxT9n/yrLhHSC5ib+SDL
GmtDGzo4sZHJWv5fVdqW1LvVpgg3Hyfu4txLLSEgO45wL3rPjB59ID8WM0bqWQfr
EVx4NkdBCjBDM7RTIdFobIeTOlOEjdeTTQcS7JYlDuWwiJSFM5dEBDtcF2EiH5wc
VTz5Ti0LARQ3CbnuOJGfdBgLSmG8Fhl6yEO6CjrlHjzHK2TYm4RrGwQWGHonGHqk
jSrq1+VlaPXWf9/DE4zZg6BtvMZgsyZAChcPy47GE0VojKP7RVtB0EQo9bmtYHco
aXrS8EB425P/jqc8BslBIIllotgXS4tpZ1O7+NLHtI6VFo6i/ANPc5kprLIfIdV2
kNJXeqCOn4wER/WcXvH6WL8d2VMtHy161u00/c53F7jXFPdWlirSzSPePHW9CZ4y
jGIDgsCy1XoXG5EIS4lzRx15JpCYwUDWQwuYtbMZaDCqp6VwCj3W6iGT5Fsey22+
+o352XvUYpLMXb6DbczevV0syyAaj3sD5FuDzTJnDBDjszp4GZagd2YZtW/34m++
jttCJa1qysJUXJUBiYokXW0lAHmE6mzYcOXrTAANPomGt7/nuBKtFk/GqOWacyWa
x/w2XqTC90B7K0x7U/JZb8ANURYdRDkaibm4BXJUNMUoDJFfTnsvamS4DZff4zCD
ZJH0h4fSAorIGbdxakHnGGZRCi3s9+cU2T3JH8LUZFTwGW0Hghb7UI8Mq4w+HBXb
86EexrSNaz7a803g+CF6dV4Pvra/51xfN7GSa0klIj3JrtvnbtkVax0RY8x/PN85
40tSD+Efnks9OioFkpTZbN3Nj9ZR9UW5gxh6pc52XzpzRqZ9aHZ112+yU7WoXUvC
nSp4btW7Wod3YNx7aRAITBpB1Qymx8UoqHiptrKspe/CY3dywHplBPgC7jmCGxSB
yS7fTvH3XUQYqQPOLcvW1gc0SWM+gM+3x7TCCeuIzwqZ/a/Hazghrz6xZ8qonhND
yxwrKD0sxSPr/LidsLbVINihhBlhcgC8/rnoM7QUA3VYnmloaaoGJ4QnErtJP3Zi
5reBJqGULibGJzD/VM0hixfCVhCjkpTNs7IKPrY6gvXQwKxamXdyph0u3GH2Fk7T
JK+Zi9HKpaqFyQb57T0x7Xgma+iDgZlFR18Fakw2L6QEy7BWLKL4c+F61UxxPYZW
RZyO/pIj4QDGgRCyVjWAR3DxnyxTXusxDryHpmN4IkbmKmuNgGgz3znT+jm4jRnL
njrpZ3s24iAYOrtD6bP4+ZzRESKGDLYccTs6aprb+W//HcZcnwXIRjgdGw+gXC/Q
zLO88+0x6ta1wCLHUwvj6/cAkgaj63slIB5KYND1MbhV/Tc/FBVzHVg10pbBgqOF
HS/MKXz2q5lDgsnQw+IDFiAn/EwjTyleFvnU4EuvgWFlDVRz5f7oNqRzdh59n5ES
w15d582wWJETCS9H2Kiw9TT0W0mU2oWa3zWTEm06Zarrli3QBTSdcaN1i/6IaelI
Qq6dDTRD/Lrgsg+7+ERtJxLOaNEPkoV9xopv9dqiYC8B1gJFTMPctt8zE2YoyYYs
LVa8mwcM+5nPcR7n5Rd79fCUioql2kCWIusGurbkMxGSsftW1L4FC7DI/iWbSCSm
KrLgYiUEwDj/QmQI6voIEe6qkFC90DQACYMZcz5kmdYkMP97cgOuntBoWLMicQmW
pGpXXNeB8sV1yn0yB1mfZX4JEyUi/HL29Lw4Egwq6NisfDhzo7eQkGAaKFwAAzBF
1d/6yamtlR0qwR7YtzaryvwY4DFVVhCeG0IlZf5ehOu6bHFFfj+DlhKz6sWSOiVB
VVwFmhN7ZiXBjAAteepbauRXdCIBlTbdM++wkzN45Hk3QAsnwSoHVK7i7npSITc0
pej3RyGySrMEQhZ1KhdhA5d2cB44Q938L1iVUhTLPF64wgS9dEWDl9FPwzD/Vl3U
8BeNkzpDuELl7/Q3nZoYE3zKZrTBbXU3G5BfedAKGvGR20QuXifqTWCJd5HuTsxl
6T8oz+9WA849T5xQcWKk2vQQRxpWwaOSD3qD9EbSLvkmGr8ei41eEp8GsR+IVoTs
KwzPINeBKTvghDiVZO+meVCX64spQnymFuBSc0zDCG2nNJpLCbo2BBFkR0U3ypdx
jikdxD/Qh+DlXl/omrQ+ZKP5mFkvZtTVHXFWh60DG0yiaqp3++UeioZmfNZBUmCC
KsFpPrVGty2XA08pLGmSjOUbSbKcBPyAGaMKNnjgCW2+R3XzcRYhSBeTdDDz/lmf
U0n7ZyBob5LkOfEl6dA0Zf2nO9Jv2pfvhji0qme4OssbT+9Xt8ke4aSbKAwGhavF
q/R08SzmCMq9Ife3AJPzdtz3IFqhetIDBdIKL2ugaVWjINswuR9R26ZQ5PwNWNXy
koq/S5Ml/GziRPJnGkzpMkdiYi7ELxgpVtdcLxSF32Y0NLmBBwVdXJ7rFdr7vF1a
mf9TjrOXxXPd3BAH5bPXeTREpuR4w4VrVEY19NmNy4iHGlQNIWMv36x0+n6ZiYdv
hxJtaYtLuAbxd/h8YRPYgpxtxTt5mxS8iDQ+lu8jzIuM4oAgWY08gGVusA7P+a8M
3LgPLuifSImBKkX1ki2tM001kYvvmFn9G6Uvxv7m3ws=
`protect END_PROTECTED
