`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aPGjxNpMP34oB+edvOHD2TQqK5e8xzL5pfTSXgh971Wibukl9Gj0tgfHwoe2KpmC
XQv+H3/9fqsm9Nlj63vxcCOeq7iLujaQpv+I+gt9PdlHzmfiUums+SGijcNxBqCB
TJLB2OBT6lwYQNHES9ksXC/GhvFbU8E26eSM2HwwGjGpBEsL2jeWLS/ONYPPQP59
BLqa2qg/ml+n8Z6JxO+wXOV/ZY+rdY/YwfxUkQk/l8mEleEXIWKpNpLRy6E/TxEd
FQtsXNZVyhs2WrSqpex7NvnNFa/umJ5XbPBXMg/ZOAyB+UagWoUEQKbgKWWcsScK
Hbh/koL6reM9PXIKCQUXXc9FIMUB590BzV91ECQLOHtknEVezWaY2oTvoUMR1pE8
t2WitgCarN+RFFH7WErff/4jN1tMg86lyAZHrR19OkVFSoeQif06GEPwQJTwb3k3
HjxvBfpeqHO4UE96TLbd3rTrfKmGbKkBznr4xHNBnAq2tQq9P2wOYW5RsDM4jOcj
p+3usLsls+H44Ejz6U3vX1ZDf1F/px71C3nmFu2a2cNj+GZbwH0bgbTMDV+74blj
+A404jdZoPvWN3PoPBruDEdSM7MsngytSQh2/vx2zofK5uYxboUotfmokVIdZhxU
aVNNOMv5MpG9Q0IvLlyF18UC/BVeybJaVaScMRceYkUM7ReW/2V4XqRhn2pLvPXV
Rpc50uQU6DH+cps3MyhLjVl/zoFhuxE7HR+f28S6w4oXdy2SmDFevJXeA2bY3uYK
nXa0xFHzj7PLU9wOZEZniO7mDUCvYday6Atyi4sKmeq9ICethvijLdNIrsmsh7Yd
9w+CBHCF/ZrlJ3m8raWJVcwMXu/EftAJhmHWDYKpVoDTy5CEfsk+uhi+GS2VPQh/
rNLeDUTBkug6k+RmwAypLCBH5XwqxLo8Vqto/zIyGRPJB+VArLtlDLApV/zsk5JH
N1jT21xlWfTcGIl5B7B9ZP2iJfh2amYMKT/Wjvdc7r5RwMB8jY+mEoHl0HqthtFU
DGTgWdgd0qhYimFTdiY/Y8ZWQqb051DMVm0OLcJoaaYMmXa9JOHn8haspG8ssW74
fJo8NuzRub07Fu0Pua7bd8/uECOrAPoE5ZZm+WerNM3fXjbqlqLAD9gLBiV/awbz
h2UKMNbghwNfvclifwHdQhWAWjFu47DCS7rqIEIQp2McAYZbLCYNWzpu7UzU51CJ
p7QMb/utqHWe6k+ZvXpVcqvKNzav3ZHb1nQAGN0ES8AS10XwwZUGqqrGN1atJF7U
atmj1xwALaWPAKGDwgmZFVr7dDNJl4/UIGpBdMB/l70NjVAJ2HlsMyQhGSUq9POj
C/NKU+WjnraxP1boSjikRm3Mc8hiL/tPHaMkNGi8Fubf9js93VTmgOi0SpRB4BEo
Y2Yd9XwH/FDYsaZ8/Qc84GifATyx0MTrzPy0UD1HwG5/N60QSa1GqGDhCF35ki/q
AidOgLtzA+8hANYHXHa2XAsLNA5ZSp7lEwHouvqTPu+J0LpAsI/d0lfJvzMnz/pU
uOT/03sT0yLD7G6uGvhMycUOMA5o/nHmBHwpyX7i4xyrp2TOEPsB9cuxn05xqK6N
e43yXIR2p9u79eNWIqEqIKqm27pLBI69DN4vcVTAOIUPVxMv1pCYh/F7m+BPyPHO
NR9KPyseDM5tHe6Hn+1g6qgWs7BkUQxX1dQYLiizT4vdhsuKnmFdFngQ9OkOJtYk
KFVWul/mzZm45QWwEteLAG++EDf3Srxp+rRBvxgEFfxtINHojYEUaU5hEtMvCLsG
Ts1O0uWBZKTnZvo/ldzBcfMizEe0Ufq6YIPwIGFeSR6iZcq7gVfApiFch1XYBoQ1
pYQlp7JTS27e4qhS3Nswaat0NaoIRVX/SQll9+DANPk6xyYHQlUgFJf59Ld+eYT/
A25+bV85CNjgDKUkDHNRMQ==
`protect END_PROTECTED
