`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5F93V9UX+PEkc9BjibMHkKwbw7M24x4QtMEUWjfJy91FIDROxBrDDEu88/m5X5cV
bDJlgVnBbriIWJ8z0tzk9IwgVP/p1MMkyfecOZyzSHzzOYLIDkSaDEe/HWoYaCOv
QDYB0gD0es3uUbTU39jA4c1mEZdWVRiCYy+UUNbeOOgV5RuKJjDtINo01te3x7nx
9CBGqaVRqRCzTAUxK/Ap996q5o1isRbAVafu0p4couKOwhahqk/A7zUUfahmasPR
pTee/sxSweLgk0PDs14+UVyQe1TRWiff4nxqdWXAX9+iqDyqYU6eyRs/haw4wep6
ubdl9WWm9TUcNJUsaots925B4Qv3XiqSIM9lvJie0wlqwBmwVP0kykSkTkCQ/8pM
ZFbIAnREG2euXtX9fHm8g7IuI7rWZQxm27ov7lxh5y7u4KutqMl6u+3FfUtcixNk
rpHSGgs51wy4LmAGVT/NtmXONnM01YsLY5LxTBprd+EXI0UUBmO/2WiRxfnHq1L1
ax640Vh5C+TuLguSpBEZ2b33YOVtEq8MH3SCNo2LwjBpTS5bow4OWrGb7RVq+CCP
2/TpGK1dTQhGi3BQi9Ow3gukhNEcQnz90KdMuqoHDR6yguE2cz0yAmtsJyu35Sg5
3J1T7aMIvAMJvojiOnafgv1OYMrqd8B7gFpQa2osGh6e6tMR/Pdme/elZQPq2kIj
cFQQcisHoaIL6kFUqnKd7+Zvw4eFl9g4lXqiPX9tv1jEOo+TKTb80qOFexRoRk9k
oJrkGmZm7+d4vQ+3DE4P/6T/J8UZA6UiwhXqZQvgFphLj8Ru7l5x73p3OOexC20y
Wj/Y9LlUZmaGCYxnOfPGGRgICM0bDe65ximN7X+jiCOfpTq4pgOSZDjpsjmIkGod
t+GT9/uH+lACRCGE8o8UtkHFMDZK1Gr1uB9IvH2mUQh+GsrtG8f7WUQhmYFB8LRl
fBqMS80/Z8UuXqSxbE0cQFkkYl1Bi+rm3G4a0WxgHqjjhc/NT+AYVF+MEqZVb6Yh
HzM8z5M1XKfZIS++XXxNvXwbth4RCjTC1iL4P74Ett4=
`protect END_PROTECTED
