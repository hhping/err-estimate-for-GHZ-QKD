`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mPP61dDlW9hA3e0utCXb86rRITrTPV0v705Ehq9XHPzfygR9VWJy9SGTiqbxxQiR
OASi0ScbHEn93zSwWngX6aop9ZVqtt1hV+R6rK5eRtxspSAr5mChDsa7+Lp0UNTH
CIZOuBXwlehi/cJTLfYqbSCU1O8amb3NDYw0k+TBOzRXm+RonJREav10xjLnSZ/v
uuXm7uGnatu2g1OadZFl6vX1Ob7aTnWWudphK07w6tlhFFHMnphzEzAOYwxIY/fR
HJ40J3wGla9THfZBxRoiD0IjD3nI+MRdlFKhQd++65JkoBdSrXQ1UJk8t0/fnNcr
nzxUeSoOCz5KsvKcoM1mNbhL/7bQz1emX0EOHf7+VTeCrGaeqIIGIQMyZOJXTAv6
w5To621BLDYFLdYc3LK9Hys44OTlSBwbwiR90kzzIc2WzhoyHfPaSslMByhLeld4
1os3dS5paPCmNL+QSWHBqwSQrbbvuZEYTEcEij0LdyLoXG0bAkPqWoEHCqCWgDOv
RzLkv/V3cUDkrB0NWmBJV60wybZtz4d64HKI6prTV5nsGFD6SkUD5vgDgld3n/r4
mfDhJvodfv8ZsR9JVW6Ebidn6RCJM3erFEg5QtgQlDvqbG/jX8ym9U9vRixe4P7E
6SvBfq6RVYrpLF0fZR8xKvaGPa6+G+ZpLigmra25BHcj06tAxHiN4rzgZeqiZrzu
jDb2ySmfJo17D/E8VsU2wo+kCjekkga1ElnyibqFp0ChfjerAN1eopWPhV6LDFVU
gtNt5FGnM8ZjMoJUWZH2Yv23yWPwKl8Yo/vR3axUBRvpF+7var3qOoKRm3pDIWaU
RRnB6OQQvpse0/EZsjmY74SR9lxu0p+yT9lSoj+IeA5CJpUItpMLhZGUy6dhYQ+O
O0DbiGo6bp+P7mscI9OK2Ak0GURBisqgMisoaui+vbaUQ8rkG+YSU4klKSv81VK1
YhR36pTJF3WiZ2QrAh14rKI9QkZYSh17tTU/6R5YjMPy1KAoKz3NyS+LiH0O+Kry
9vHpw2PA+LTNObh1pC5a7h26Ja4i/mpKKdAaQd7GCil4ZqzuLkBPADXFAgp71ehF
UtTSqFHP0m2dQGY93blH72LUD7N3v9tzbJlHiZnA08dIKGFs+/j9QR5OTPbVATNc
ktBv5uKTlJkbCEhnpMa7pPKjoe4VQjJKUI7h+/59qixJflxe0y3iLrF+pC8R0In/
qV2DDfG7Onl/eVSuUv3outIag/HGmxVev3LRirqelppCTzkycAF9jER6PJxKkGPc
BHfQ/WV8NjkooiDDdfZ0krc1Hiacww1l0VErbmPuLzd+fdw84o0tA6aR0+sqcTyU
ASus7EIYJ41dXiOdAAfZQIJ4SUzRHpUZtNe1phQ8YQOUY9WNIlPOD0Cfy4uzBX1M
ftf+0kiEMZz8Nscge8WIVpY/Lkv7gwfY8lBKNRFI563mrFt6Whyu+8pr0PuTFXVL
Ag7igljDsWbZoLuChE/l7n1sc78kqol0xAsnskX8dhEp2jVnh+N8k03TnnOXpyCC
ggLL43h/JQzULzK7XLa4+vE6oqPznWQXAWMsuOzERlwNjFnz5EPNLKBZncie54Sb
4xrNWXBomTKYR6RTu881YSH/8qjgHVbxahmQXo5OGwIsQLp9dc+k4BceiwRV5Zx/
EsA7AuaBWhOjy8vwoUFAh6pMGOYgKdUz+9muCwu9mJ1Y9cViGdm3Yk4hQKG7NRU6
ROOgDUNfo6Wjha8gmVgQKadbRWRmbXsHcPANmkKLA3p4zAn6yFEs4deqFXDiz94O
JOOV/dt31erjReIlkemjB5SKd3qNKU/KoRWgfI0UM41rVQE6NYOmJmAsC11y81NO
PvpNMEyqe1SOsjFsltSDDmc7pRV1JaijxZ21uZqdjKX2iHIHglc36u0vGliQMSk1
J7AxyCkip5n0/tUiETSiAgpVB5zbQxaU5657sQgMrABsgL8vLXI8ggeKbTOpW4bY
EcOHwQItTXlGn2/iEmo5ZEI2SiVnPQOu3wZFdb3iTalm/oPlmF8fCUGIca8sRTJw
WCWscAKWP7+g2Eu+X+IhMnDPi4f9DEXWMhuGuVRn5+HJ8X3fveAbt8amNgzSMgAu
vRLqT/otGVMjM9DJzMtOLcBGLTIWmARgq8MSlQ4mX+BMuxv1qxvMz8DB7QY39ClJ
4fXdmwfq41qOeMczqlAaHprydJsnMW0t6GjfUruDzZhPk+SBvdEvPYE/rCLWXpTT
mAb+u83KyqYgtMyeFCEs/kQZj8qGt3P6H+5XrG0WDlXqHzDKQVbD4SFcU/6tIX6A
vCRSwR2GMT4yzUmo9XDYv427JzCFALVGOS6hldBDgde0dJXfOLr9CMguOFOE+pQi
WgyvLp8tZnhGQNzC8t91oGtAN+Ama8r5J2rEmLSTeLFtajXnDoDYHD+n3Gn8RwKU
iR4WBtzyOnKTFQIV0JAdL5YAMklWXO5GzUGx6od8cIaexIP1qMqpGKZG2h6of3gP
gP9RuysYqL9vBLGxxFlFSgZtvCZQ9daKaKB6FRr0wCDwmWC/LfDnm0QJK1jinJbp
skSGXGtOEp0q7b93xekzePir8uvvpyqZF61mLiDEfjAB3fVhtTqkXXQpogyCQlXN
WZ7ICrMFQBL6FQxx1kuL3vMQfnVzHKskxjuW7L7tnG+mRSQCPPewOsqsiX7IjbYw
cpnD1tNovB38Jkwt64ViwnQMuDA0UsnTtq1zg8HbQ8i7DiurfKGEwIOLNkms/zZQ
Jy0T+fJ9xohoq41NJq4fAZAE4HmSZaANYNsBaA3YQfctrl1gEnq/LDkLYO4056Z7
bBrvTBcQYlqemlxvqhtPdCQ2e69iN62CIXSRzHOmQUfB1eLR3iIXgHg+wcJxtFLX
LibT/B3QUrIPl+LA0ucr04VDblSLBzZUBpSPQloLdVKIXJC03lpD91ZTTqfVC5+Y
CKJ8DmUjjbgkANcBigzv6hruoV41jZcT73zawfVBSVnj27WSaWWqEbpB/GHYycYh
JfwnhG1cEEfTnCuiOh1vjA/x0MJSQ0U6d3dEVnHK6Bbxm7m4ME0f628vAqIvFFfq
`protect END_PROTECTED
