`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X7P0EQ21JFNd7Mx+WYYfiKuTGw5czNx3ADm1UQIGDjwnMPrpMvQJgbWMoDqgZGda
VRUMONp14OoSD48usNS2t0qyqkJjh7r9wKwfxCIVdnD/sKZqBblfPNJlxEO8FZAe
vT/xI5mSO78qHd2OaXvDtnl9EZUMs5aUqaSwNEdLbiVvV7FGiBnIXTzlYM5QvgeB
ZudZ1R8JPNvx2u/V87JTpWQQAKLutL+SWJLlv6kENRw8IaULCReASWvZnrzFnycS
kK8D93AdRrMoFvdqZtUaKUjSLSSMoW5/bfug95LAcAdTITfOIjMfV/Avbx2Nm+cQ
jwLBcVxL8oUgRir0QlYGqQGdUA12AnYSoFyQI6XWNnqJsnL/8Lectxo70uyMlR1h
L9b2Z1fCbgyI/ctO1rQJLpLIsoIjQFDBYSlNYUvHCEOkkeGO1pJ65Vz+z8iKuhJE
DcedpmEtho5q9hqMHo74WFhHvnTzfsAbfl+ajP/Je5S96Pqf+k/zaRE9EoJnKM25
+++HzdBSj14mmUnA1SpM+U3VWdkopHe+nP9+e3pphpZx/P7quXxar7Akt5G9mwbe
KqFL7+itxBU4NWpwWNzddeLm3HsTuWSVWhBsuYNwDcAXpZGS6AbvHcZGEtPfxKI4
BVOURgeozJP3t1Y1VonipWwSMqUtwqDTuXFlcjDrtplC3IvYN89j2dBl7rI1T2A6
uYwROmsYtB6eUhhWg5pz5Rjs2RBECWFNN48fb4bGvRTa6p32IHTMb5Vj8WFH12q5
OUgyFNj91tTNl05p/pnmy6SxpvXXvk+uKhiBY7eA5I1WLtq80MJEYsLJby6N49yK
AVOqX+5Him2WSsb4jHCdSQAd8ppCYXkfTbhP43MeZDg+rCfAvFywzzK/kUJrk4mk
pJeoCCwdSa81hmGpYMsLJQ4s5UDKtVCfERgtQYpojQgks675lBAswJnALJZhRu46
`protect END_PROTECTED
