`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HAZVL0y5pxXOD8gOoh70oldoFKwSF50JWpOGpBQmtRyzoM9pjGyj8ttSoXM6gmMs
uT6vvVqOXvav1dah74mXFhrHWCKGC1Hury/CfNv16wEH4rzgXCW/lCr4cq7v1G8b
2JOK0AXbTpDehmZMZZ8EfEO43EhBIpgZPi0I3JP6Fc9/sZIn8TkJHSqA3kqBeciQ
65xxg3RhodRTXmp/sM3/4R58+ZgYzMKqvv3M7uiJ9TEmHx5QpswXItGegmkFcUd0
1qFKbgxnCfy53M04+oJCkA9dc+1YgPpHww5Vybiv17RZkD4cuEe2T+2kuRqvOpZz
/vpizPhgkVYVzsbVmGNMdhS55sCiUL6K7VTTeFF83Egb9ZDA6AA16KvI9R5eliAQ
ISGBAKNRiG6j2oJsP/q3DHf92p42bXifs9lBVP/jIYHxcKHRa+pkQ5frWlW6lKjI
b863A1MvejogwIjq/V4WihPv3PwRyBYil0vvgeulbAXHAwW6HRlvEYpQhzizXdUn
03rlOg8TvWK6aSuxxkb/EEWUU1mXr4kFR6yL+dUeA+uSUV1rs7E9pr327AYPepvu
SSu3Lb86/UKqmJs4+ZZAazo6H8Co4hGXCq5mHMUKeI5M0fioVU1ZAUK0pNAPRLzh
jtdK/ifAXGWq/EUdlR8zluH6X02mZIbga19576ia9/L7xgO6oaeQUdLB/jwjXbml
CzPvGYsPN8y524nCeNqDEyivgtxV8JOZm0EqVfghsrGPZtZ6njMX9tsGDi5gi/RN
2jCvvvvk/a9iCngZ3iLeqLEJFto/pLaNCBK+oJQJ2I82y2ORN+xKPg22aseFGoJ0
rMsE6duQM/X6hQHMpKYQkX/C+R5t8yzqN5IByqvA4T/ZZDEePtdmjs2DAUxzbHL9
IH9nlAR4pc3WC1CbxlFk9R1P0P5F9ZU8w2FXbt/XAMB6GAzbZ2zPNKvg5PyA5GzY
sEeWChrnSZJbXoeOVjBjp8M2QpMPkGQsrbCB518XRutB9gQ4QxBleRW9y4qkuy6Z
fyawveFAfPqmhwdQH84QmoxS11XKeM4QEkcipzR+pUTmGb3oJZJpeHUiASBklNd4
cuSDS5vRa5JCPU7pNfx9jle3uzLN/Wx2EUYZe4dUzZBGHnMgnm9EUaPdEZUmsL6b
Kp7hcZL5DNLV0AGpNIxHq7UL2Qn3z8bmt27st/4ATbM8CWf7AHfHVPX16iZgXHE1
Kbgt6PGL28mT2XteDSlEaNUv+69jZtd2filhL6CZwuiAQ9CkSGsmvEma+v6yg1fS
7VygPrqVg7CzENL1SXpEK0iUBvf2J2MCC02RB+FTzyfX1CNSlzJS3o6vDP+PyzLr
iQxDY6X6UcMzofrHhLywPDMGMhHbkoqcM8rNEL+w7BZXgCYR8i3x0HuX+X24UcAy
qFZet878FMrUr4/q9pFEQYBjQp0dNo26A94O03A9G588ranx+ckTmgKl0N7JU34S
TRQI+69AzW4lCgre1ZaD74nTJ2odcS/M1NfsINpQ5gMdN7U3MTeXQhMqom1/fXqf
hTQ/rdW9w5GqnQwsa153+BG92tMDcitAkr1JDQF5SLDlWzrHdhMuooXYy2wmFnza
EH6X1UCD1mEChRr6Jp0TVG3IchxFez+97O/DIqSWiDcsadwIHcyLqll8YnzgQvDC
BFRf0dkTAtT89w91gUd9pOXp5aiAyRvrng1fhg3y23pBsKjJwjVm1/TIjcoIapBH
b0sECrJn3pJ/nD4kxw62X6xQQvj62slk+9Fi08pdXglwOKVcDeHp+0V9T/ZNSFLM
+Z0i0pb3xYC4rXTCUzla0BdTU03F8lFSfTbSe/CSOa/sQ/n5yV+WL8OkHT2v3eTS
SYNBLTrz/l7UINWf5qHAsGDf3xiqIBzvLTDY09LDJy0sId/wOh40n1CX2Sv+UkRd
sEdoLNfDmWuHd8zKrIg+J6zu6i0OBDP+P085HvIvJHo0StD7HiLCNm46g/UepgVZ
On/XX94c+kZI/38pYgf+noAejA0lNRK0IRHSSmNJOv9Rx8k5absJJ7Z8z7Y4qHyk
dCCw+2HwsCA4nJg18xoS5PY4htz9YJsDTHab6t3YMRJGu/muaw60LkgTwMNdhjBT
UFSNUQvzkJvLFlpmK0RyM6SMDlnmMiQiyDLqR0l/nmIjEJ035kUnVhILQKYr7W7m
SiIn7YqQqmt5FFZAZSQS27MwvYO3Xmo8CGWR4DwMxXYwTUYMxFL/w4Pg5fpr+MS7
lHQpLN2c/q3HAn2+kgbFhkn3jAZesO414gnrOocgQHDKSuYlVTHnNsE2DuCG/yrR
SCPRSZmJR/8GUC63NJX2dYLO9z0rutXXmpEfubV5qWxCe01UZjiIg7E/C3ybz8Oj
6nRsZhHSzSdcC1Icn/p0EnAb0DbR8v8X2xfN0daF0MZS8mU6GnDt0MRl41iIceSX
pcTPNwCnC8fk9ohu7CfoUvRUgdeVMyyrAAXOiuTmpvA=
`protect END_PROTECTED
