`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZIaV5bIe4BCHGcvMWm8KP2OJt966cOZop+PL/JCfY7ahv7EkFbfmcY0NEVSGQzE/
5IAtUclSGNwRNOTjyjzvsuyJAFU4Vtv9sqTwNkuTQg0M4msfcjtF8+wT+Fk4CuFo
sy0vsfA26xnoTn1MtSAVp1w3sASZtL8TNoyD9l0KxPU7grjtxF01Av78pqEj6jX4
H3LPKpEfPEdosypQsLAa3tQ+UENLcvr1A9G1f454W+GvVXkcmzPJhXmEc32+1WJ7
PtJ0o02MUvNJFucrWMLoT7GnnObGAuZtlel2JisB4aBBVGDGWc+BASkqaFzP7AzG
erKqQQncigTTaudllmU2BeunUi1v7/2mMZs3oUJHVpm31xaOZib4xUPUUDtZOKke
tJJdjITikvZsoD5HREXrsHWffJLk/ir15XWh3jcXcij7Xbb4VhVLrrg12PzGsEkP
NF2nYgI+l0S0Tzlw3/rpC2NpHu73yDyJkzrchCjbsZ9Cc7hVt7d0c1LjSWmx93+8
F3PDxeYN3fobU0CYgVhPKpqf4s5vV/+CUto18UzctZOkOX+9tQZE8m3NuO7sTKMC
Nol+ggqMsQfatJQVW5G7bgDp0uocJd/jaeud/cJFTaKTbbSsK38gCYLCIdY6uUPE
8WVXm4UTHZUNDR4c5/ymq9INyDr/8B19yf4BFlQ1LTMXUYL66FJjXkGJG9wPthsf
jeSOkUNmMU38aWe8Z02VnjJc+ygjjdXzmf1XaQR0x8MoIMP+xKyTDvcqR91M+zu4
ku0o3TbIMbPyfAIWwQyDW5zwHVz7wtJiInzXpn++LiRuOzPY97VLyqzTl8PTC2KF
ihOQUsT6WOt9Ms4By9wCJtZqIrdefBokiJm6QzJ9OpNz6C3Sw+DSA3j5IuTvFX15
6F2jyK0spaOX3Y5r4l6H1DIUcVTAntTCITb80ecccsXXiZ84AxYWz6XpXnFAri3+
Z4DqBBr2llGjGsuUQwhIz4DSpqlUUL0RLg65vF0xO6H+yil5r/bsdlW5j1IOXsi7
2hPMsAze6Ylaa9MT/kepnpj77TUDn/5VL8u6EE8NdBoBFW3s3Lvptf003n2BeIP9
kHwz7XIc8Apz41WgtIp1+NfYWNBtV8ZhM1R/+AqAf9UMBrE0k1/eGvnWe04YANoK
5BSKYeoQc/gGqvXKG+0gcDq9LZ6OIlTYx1rfOli6qvSVca3X7M4kpiDKbgsLGtBm
aJJRchxWAJ6bPwsDltqhyHRdT4apuRVpVX4aQEsZbbzbfW7+YYwmreGvynXxgLfr
qQAcO70fMKourcRTvDRVUiSfxcMo28YsedX3SYShW7lKm15XkFx4LFnE2YuG4Jwy
KOW1sbCNHJIKvIBrJ/MM8sRmA3CVwXYWpzC7/qjgeiF6IDpcdlEI7TiTpavylZK6
aiwiLD35Xzdwfkf9jYyI2TR/un+Q2JzqY8E6PFHOI1mSpzLgaFX3EfegMO6KeBc2
sI0tWmeddXVXvdche1vHtQ==
`protect END_PROTECTED
