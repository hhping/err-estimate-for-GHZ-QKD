`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2um600rpv8UGtzahmNDutKX+KlUQVRUXgLPONwi2TvA8m/o4294vFaxldgceB5hN
hxWtJxd+6MqBo1innX0+3P6eS6K171VhVwm5rh3DZI3pvMok01uAWksmrQRYps7X
ETWYLe7Kef9kplkvgyAlMwVcxQbymY7+bCW3up/KqIgl684lizk5SK8Dk2FTZlex
1CJSddp9UYpjCQVKjhDHKzlKVE9eMSjty9cr1kwqthRk9l7luDdE2zcFypjuIoOD
I1AUx2FshvmLaP03a2uomj06i3DF90w0M+CXKdsRpOd1EVHbtjt9R2b/zdr/ZS4h
qjk+quH+yVxXvebqedweGKtn1vWvLFmpFZl46vA2UdTQhXVp9V9K39qy8HEePkft
dCUJG7lxE4RSFuzjvJLPaSTIRlVE6Yz2QxIk5r9c4LmFFQ71598+CQw+rogjWL3Y
3FNFxUXR2Zuymf0AS2dUGtcAdDId1EFs+1N2EQtYIm7m2uZasog6o5AGHpeNxx2i
ibC3k7faHnl+2oRrq6FjP1mWOL0VKPEzCKwUwMV+p1okc8mdQDB47Crv0kQJnH0W
KSt+i1vKW4Yd7urczZcWz77f++R8Rdidb8q3B92F89rDma1iYLe61Q17V5dOJeX5
gWpoAoTNwW1XlKcOjP5CTNt8a5XP4T3mX2uDb1ZfhWesCm2kX5nNb8BJbrffvz7N
WChGhdI8UZEZBwJj/4rpDhPF+pNBeeP6xj43ezNMYKnJruC/FT1pSqfU3FTxm0vJ
ebx5v2KRL9sJu1aq5qaipajLMc+5y4FhTAQAyedvAbTPe9ZZKLsE5Js7mxOm+x1M
VRzltmEHG7C90GMsLUcQOm38R8HeESCb2m1eZATTu6qXZMVLerBjwm7MoOyEvSTl
QRV5k/5YVcRtJU3q73GFkUqmkXJKlHTg2YyzubIi/LG2fw7tVERo47kjpboGGpKa
hNEhkVEkINMxgv+NaTGFpEh8Q81Rd7yYmwLhVdD+cmkthNOYKNlvsD5MK93rFBWf
rgpmtTG3riUgfWOVuw/FzXUIb4HmRa78oLiVPeY08R18tscYOTuWW49pduaJUuF0
GrLC8Z07blJiqCiqtSNqbl1R6s5/TsDSwLlhzx9/ktppqY/Om5MI2JQ7iiMyiiWi
RHQqjaeLD3frcGnnGX7hfcgs1dQ2InQHyblRrAFPZMwFVaMje51J7tinKCd7RNyf
6dyQ4KzQuomaMnUc9tBrhaL7PjXA5cYOS1sk1CUHBYkoI8bjev475LyIHv/iLaSL
Rk4dOqidg/FmNze/dJCaC04nSjcEFUBwbrYjPHhGGLg0y1Un6+wOrz4SJs9c32Go
sIOLQe3qJSG4LPqW8jNLGLpFNrnNb11jeMBpZzXDnxTszmaksk9OXBovhxUcK2dV
8QIGvUbF1RHzlA8vybOSLLcm65bjL/HoNSQBsZT6qTgq6NzEzFa4ACJBgahEYaMe
ONVcK/SyLstjK4IiZJfxiZk109erEXvAz0Dv459egPwb8VDwpzZnfDA2kRYRuwNb
HbHlbJ5VxFUPC8j5aMGvM2/2ARYklrqSNyBMaBs3de19EmkiaAunAv8Amje91bWF
a3eDqM7mUqJ5T5oN26RANk5kuSB6aBsz7P7zZtET8ScP8bU7ZZMTy0g9U3iOucxd
PQRXlSnZ73HJ0n/6+1wJNpUaN/wzn/Tn30tzMO+ilUEE/41S09yQvNVfsOxk5AdH
Z1Sze7h1H6Y4jzyI2ufLOcMwQDX23sbYZ9MaZ0y3ed73uOhm7IN9q94X5Dym5vdU
klmFi/3TTuqk4eyOBOSBdIQc686CrAi3spPBNtzC8wS5KZx0xUGNfoWIkLG0N/k+
Hr2CgA7BIC0e8h6IxehpaIeHfaf3rRro1f2HZ/4ajRN3QCCrmHyN/Ua3vxYiCmmL
ZyERFcgKxeKYKuHh/+LrPRwIymmsbJZN6fKQkTgxkMYxMbPE7xe5FqO6tp3sD/FZ
IsvFo14cNqg1LwTUeHdOUtxw/HuvOEVAC5fZ4a1LZl0knlW9xbtg+oEBY/OGwpij
YSUpP05rVrYqV9WW5++Sknj6pqU4bx5QXZU32neaR5c7W2hAI/07DtVCBjjJp9eu
snZBViNx81gpR9udPI0UzcP7RUEPiN0MJYSuX6c9WMixE/t8N7U1QNTR7PWeZfCU
hWp4NQrIeooQJgXUo9t+gtM+NK87V35ZeVX8P8wqMjP10N6jVAgf/3FHu6r203gg
mxeOsSIyFjHy5xxM2BjDxIWKn5FWuJFuJEXM/4qOXaIGl1MeqfRVLwQraaKpVij0
RYDxv/UCZhh6yB48Vvfdiprrxg+YRHwfjPcDcfvuc2IGYYkiYkbrh1OyIDHzkBAI
fJlGNkNgkVhGJ+FsyzGeM2yGlMorB1XiM1hmW7hqgAxFKvO3/K5T5R64rf+OUlW2
9ab4X542JIsx5VKHZu0hKsFJwUgJi1pPCfm8JxXwFE1HhdvQaV5rSZKKcQ8pN1Og
5eEDZikDof9TrgH+VNAr9bMWCe1Vb7ZYLrjWYf3pPrmtlMJmaqsuaDRZTMyPwBsc
CAUqLz3JMuZE3cG7wBQd7gQzwu9fttwTWfY2JDHFSB6cR2zG+P7gYnwjKvdHpQ4q
LJfDyirweM8epKvKBS08q800fNY/bnxbyDsApzb25xm9ludfFimABN6uf5Q5AhKJ
81O005olF6pTE7YLqnlFnZPtNf5VuwTxwItxmUHKLjKN4u2xneqRZ4ckoRzqyxHF
etk+08atcPdATp0k1mlMXvhsr1eTG5V+ObE5/fsZi/mcoFRI+hDm1ilJ0vME7/ea
El+owt1DcGNezONtBq6yxfJgFGA3y31UOnhAMJEoQFI=
`protect END_PROTECTED
