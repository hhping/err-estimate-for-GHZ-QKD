`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gldhhAEEiuMFRdJdzM3eUps4BACcTvCAbnWeycQbDdze2V8YUdMys3iMHdd3E3Hx
dC14OaYw2M2m5QLmxkW2bOtGH9iLrRvX9wOR0SkGj6okvaCEXXx6eE2CwQ08RDqo
MPNfAM50Lu0htvmwRrnqQrjyOp3hGhZMOcGMsHSdWwEq6ZQKLSlkF/wRkk3plq2N
nbEq9o1DOwHfGuYzoW2iC+Ju97GUC+/AOkzdzMW5fYRGvp0kyqifaAxXUQU4jjnu
I7WAbrSX+yOjdokFUqzijSmSaEJdGxokwuVb8yboMEFJaQ+wCxzd+kWKACBZyBnO
fyLcPuNhc3dZY8o9ymYBq7ZYrB6XmgnYeh3nwQvMG8lVHoM/Fl9bM5yH/EOlVjEF
ykoV99TGCD40bnpMnfHZdW3ejM8vj6LIErF/mLDoHGv5Cr/Vki+9fyHbMYSodhTJ
mR42/Mq8J0hD/By+/OwLag==
`protect END_PROTECTED
