`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VmCBVq3PNl8AE7C5q6j6sRajGS1kGu0kFcf5WdDUr4k9Egk2rJVZ1rnmqh3PTNF/
6SMxXG9SszTeSkxfuMcp2pCd7hcUOoj/QkCwX/wgo14AM9ZSFqG4LLm9frsppc26
HItX570td9KT10q/D7Kgpb7gq1zb2pdbTC/98o4xFy26u5U7H8TwWukfwBrOAO3b
sghgGEhmETLfPG5qY/f6UE90xU+uJqlwIDohernt+T6gyOAbFyeTUXA2yBG9GUyu
/9J8wD+gH7LQ166B5IRxwb/Oih6Fh1JQ31rHhTsZbakgRYFHjpQQpGJKgMAka/hz
Sv9wxpu/mtRox59nviXSpOFjPdQ0UBXORBTT1PH+MujYfNoh4Q3kviv4U8N1wx77
22Q/AUVilBDN7KzFRr6RQbsYv48JGYMnSwHxxxOZh262jITNnrB0QF7w7BYPVqPv
7ddY6moN6GlB4vGP42gT+koxG+a6eUhp+OHPU+hPxpKwX1OFznK2RODaK8huoxxD
a69VoZfaHsbRDV5hrHmkggoWzT9Lk+IvNhK60LjLhL9B++A0Dep4G+zioj9VJ4M3
atJUDg1N2qj2sVnoR8X43NkaRWjg7myLeFigISzwDpHLX0huzhjixhxnjegYDJHY
ay0TNONXMLa8h7vmCvR7ds2M9nY79PC11vuq/YFJb3GF6BpslS93MpjTRvlpm1Am
gu8QwGtd51vSiPsSGjsg+g==
`protect END_PROTECTED
