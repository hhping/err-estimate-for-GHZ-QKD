`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2TbyU/JTxxumxNDXJKr5fjBi2RCTdYkMg2+aT+r5GChHLEkt6echWTByog5VeT4d
DOJCXw2q1tALbhO4Vtbu/48lLj7a9ehcPhgflW1TUk9ofaebytc7rwd3lEhQ7s8a
VEW1N9rLfXc8V031+M4q6w/56oR1YQ72YpccNU55+TjU/waW9MpzvQFEflRST0+w
WaABxyy25sfeQ0N/omWxftWXkn4XFK10N+V6C7wliHKhdwLVGdOgi6cWLDjLmQcz
MgAVcaHjP0zpp/rYO7wOBWHK/ze8tXngQErsj2VQq3o0zuezjuKSAKoMp6Q/7oYM
g1w4cgwNmrTXb4nMrEJRSSk9/jgwMcAnCMgIOGIqQqg0dzZH5uqwD7Doxolyuza6
12tgtKfjTJ8nVJpO1WTfdOSUPmfhmTT5DVKfI0/cwVDYc4+MF7hnyPQxepcnQ7D9
I1XVNKJ4WNuOZHPBo3NWzGPEa+1lVf5GdVmyQf00Acp1qZBWXmJJQDkOvkSJbSP2
DCEthh+r1Qgn4jcYyCciYDHiYcpRmea91ICImj15X1KZFIeiMAkzZ7mVFRjIZZxk
lguLHczpni+KIamSVyiA28QDh3N8wSNQ6XsVlygk80v/2Vn8xPj/QLJTEOQTvZQK
9oEVjuJZkPU45tI0Bu4ixbUm5FSjk9l2YNY2nCbsHD5O8TmQ3M5a1w5j78ewk4DA
8oenQaaS5IyVVUhz4MGT9sgEsGN0tIaL8gH7kKFJl2nu93nieM+RTFQwZiq+JNGG
NE44CLcGvUGxGvQKisgm6qEgMseQr00JAuCIp4pHI+tZVr37UtCcgu4U5QJMP73i
GibJuQLzMCalo/qhu5rxIaYVnft/CG1STTbaLHOPGmTQLA3a2SS8BmsJ4bA9ntNj
0Y5ZhLI7pfmKJ3MhUvze81PqBu42FEh2s4OIxvzovKVZwyaQuL0IFeXaXdwDRJcY
dVsaN317j1GXZdUVf0JUBLoR20oSjNvF/42VzT5CIh5ILgrrEjwBoUI+KuCp4iXL
2QGKDp4W3xWYqG26Jh0oWqgcZf1KjHsTrGrydvo6WxZ1JW5scusTpmOufAWvcdnl
AJmCQXf1Qwm5FjugubMzdPFokABKK47Bwn6EC30E1Ja/njJsxwOJ/za17xYpgJrG
eqNNzzhfmFfD5eEGBAs8IrcD9p7v7361ANaTQQsPrxggiOKQerb11TTfjqyMEy6n
C2YGxWubPEBcRKCcnZzq1u625jBsvo4M6GkPKXejOClUc1/XRNrMtg6AO8wZv/vH
w/MsaMW2R7nwct1k9qRvtWJFFHoCdwMy3AddtYg4X2Q=
`protect END_PROTECTED
