`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tM+hPZt58Vmw7uVVRYARxGBq7HWDMNY99r1nHxRjYTHJU2S7RZEYr9oXvzQj7/GA
Kngs8hoztDc1T0smdtoYiexYwq2ROBVRlQTxMBNV6nI2scTGIeI99thlOj+xF4r0
mT7JOsf6NGR8IjQe4gPk990bV6gWguvnPUMcjHgbz1gFpZGJzihEth+Vl5gYR5iN
9k6cZAcwW4/PN32GNpQwNKGvyzMjh+tdr0VzNcL50VlarZue8ry0r/jlEvHe9r0I
2/8GO8d9+M10d2hbHsOvtJd0+GZkScnJqVp2fEddqxdO93eD0OLB6QAh+p1fZdz4
f0w/gzYRdzEua+bjm0RaLMxcxINk6TSBdup0BCaKz9ySGBT6xA8qqywqou/Ks+no
Z4dHCGu8Jvd0OMsZ3cL8LfXGPAQqCaa3rADewlKSP55ShRs6J2GJ0lzfo0EPWEAM
n1GpgOucsGaI+Y0UrQOGJLCfH4h2zjpBdWkbiq3hvIVtm+buJCOCAa9+aLKFQ39o
BxkVzVKVzk1XaGOTpRSt8oASsizoOfXLHXjPuWex9ZajGjvcjiLr98SEwnqBWCGb
xKU9SlwLG/uyzZRYtIrpB5S/EIYGMTNwkk4Q1xKMuSH6I+jkAQU4N8iY1Znn9eF1
Nlmsr3Tk8nNDWVqSiWWA5nK6vCd8gay4p8PJfEIXMh914NyIXdjWYqiKJrbvWPfW
Dp9t9Z5Fwb/X5N+G2P7iIQMaIwJ0gV/ey2hwUw5BnRY2ix+wQ1tKpfUBaZ2SnGPE
q99WB6QKf2z42iCY/szf92DkdH3oyay90VJ8XUfxonev22BYkYIvdH2/jhh4oyaL
wy4Gn8hsVCp0SrMSf7rExqi3oahQlGQuxHUa6kh/Bj2ZWE+kYWflQdDnRFW0PTkS
WEfBHmDYQgPJBEuRV3Qj+9iC79ylH2VxeOVperq3L3e8QCyTiFzWRNJydRZALdYI
kvBgXMiQdmwRMmYBdh8OrS9Xnyjv+2AOBRhaimExIKn+5J+VY0+l7uPjsssSqMzb
M6x1esKmgucQzxpjfkBku6tXSno1Ny1iF611zPlf3+1ilqvmHvrxT5bdYekQgnw0
++2Msch6sWDtuKVzfigczEmHLLICRngiydrPIovMSVh5kXHrgVpzDQDHtyPPRFro
M73VkHPdVrP6ZoOFXph6N2Cuj7GPuIXm7GX90BRrni8EP9cXSV+iqO3VfyKFlwCE
BiUj3UTw7FjZO0RWsJl2gDromvvfiCIKUxVnJwyxoJoE0UTjMrBX2IS4LR7qsegH
QhO7olmfOW0uthFrmqyAEFj9MpALCy83wf61aKS8lBJsK7QYHd7DYabVzg2pzYkr
sRJtwoZSsFMwdha0EvbCyY+J3SL8aku1BnJhonXOjsxy3YznkooJ86iZU+Y2y7Lo
Y9kJm+hEfC4FDY1IwnZcYVtK7NNw+h+oR7VL1eOLBcQVzsDwNHZBYQzV69yM3A0h
JTN14hCs5rT8cyhd3Sk+btR4pQ9c3jzC9ArHNTJ6ab7CAuFxulPTM5aN3YEF2TaY
Wo2LJt+dthG9Pmcbo6quF4f93BaK8EbnZ+Ee7PFh+5At7/idqdZxt/uccMcAaVnK
0gY00wiJd2EsL7Bn5ApfeNnflHBqn1aevC0eN0YKrV1lQ5LE6rk2zSJ312Lnyz+g
Vp7c740NjofFxdIwAoAZ+0nw6YcYLqJpv9QDlN1iGOyocQ/cUM5qOe37m4M11lLP
iQ3dV2eQogXlNd6Wah2iEiOxcdAPOADqzXtun+xSomqbP3Nrk9k1WcqMr7e3S3Kx
bjxmKXU+6hOeHsYHIpRw1Q77aCJ1K8ozui4pSyrDDQwvrpC+aG0qobzeIP7vvTvS
NzaazUShSalOfjojJdewOxg7K8782kqSGtI0BIEGSV3RFq+mXHnbXcKeFkAFrMPq
t/C9P3DajluSZ7Cfdmox7erFS5raNc4zAkbn3w+TOqKdZK+yph0zL6lC7jnw+4wQ
AAhu6vpxr5nvxePFvTmKeZWcWSUB8DToEjqRJuDQIsCBhj83kiObMn3h5NrBhjz0
SRdk8nvKVvhwHgr1uBwY2Wj1c/9FBK65yjvCLEGhfrTGcfMs5Atp9bqDmiXFcJrv
zJE4lhh5dI3TFruNngr8YnfP61lgXaaOXU16yWLU6qWxwmRNeTW8IBF1NdRn2Y35
5/08A0hRjCe5olZVKySFVPZLgeHO75hNUjEiJGH60g6lraRd6Av4/BzflvFC5N1Y
Pt9lDTZfCid9aVO7NADq9JeUn/B3ghOD9eBadk1hEh5AeU4KIW1gkOKX6ui/FOPu
k/HlWRmGOJQiE3Ft6KmZE/JJxX77SVnLuyKVkdwd1YTWANaIbWmXdvkmfAyg9Z50
a+ySDwOW/B09i0p1YApNwWc5rBsgCQEA9Q3vBJuVQrhEchVwjo9ehU9NVVGuLDre
bdWb9fwz0Td44qdgmsDxcUO/b1PscikRibFi+/xAxF7GY+4B1ibliXu7N1Y/5ynh
ySeIyRikd+4sVhy1zD9GOzZVpQDYc25EPDPDrSUDrqCCGhX+tNugg3l6kn5Pqjun
ooFMwQF8eU7vp4C1GRW9MmCQhjcsmzeSodwXZI/zXqsdi3wsr6pJ6Of/m2pmIGaK
OsK1wig0NfH3G1lrbgozt6XUxAmcwBQ97o8QDWhORE98QoseW8Yms2ZqS+qw/jNV
0lx9yoV8VdbaZ5CpaEwujnIl07f6EWdh8yg4KzdvjrdQSjUZiPCz3y6ZPFmQ4lrm
22xAdukGvpcuhQ3LEe57ofInxSetuWoetKsIoq380q3DcmREPLE1wPAvHMetBT2n
8hOrVaeWBglx9bVPWdBFVoCSYQ9DuKcSKqggvIu5vo81ffaOlicYUfGcKH9GUbhB
K5Is7+9qH2TRA8K8PQjd4GP7xhp6zL28i0HjlQvtRpbYUYCIgudDN61TvvnBhEEt
LGjh1w6g2JHrByHwh6zKLLtcX1FEFpiy0DV4GnGgKmWD/2mQEo+RnWOo2qXXXHGx
b+hwIQaBQf3NP7qsN7j6rJX4FzG3UifH9pjczgAwLFLErf2JIBift8NJa+ccSsZk
wpNKYtm6JFsfB2eU8DFlcjkb9iVjlHnSA0Wu88glydPxr7ihuDC4s5snkN4bvkDu
ExzrDHZX4ZgsFbZL01AFQbx2sXHhvcH/2iW1L8wkJ0Z0TeOhspDjh7mpxlp5nm6g
4SYqEd9SZ1QXGNb8O6opmUvBu8iDi+p+xhhsTl8epeTJSHsRUGEp3/jcC93HYE8G
hyinpd4Io8WJffDMbcPjFksU7zhpzjIs5GQEOXmTqoAZ6DB9QNQ8l8TDvvmM9SFf
mY8E4LXM3mnM8k+HFE6aCq+FYARW8CJfHM1B1yqYejFltru4m218xRJAoOfW+vZ8
b7W6+rQwpwPfSdQePvUsv+0CUr7Qir0gNZ0LXL2/yir5eohv/GAry+RYZ9kPgPHv
9WFKHDb3A0ExIN40c6CGKSKmB/hr70f1xLLWrRc8gPAW9iGz8S0Mp7cAiQzUW34b
Q/ErxDAUmMWSjBqyyCEDdTJO2RNmQKzquZNzgfhy5s9XXLWXHMRaesj2SJf2TuH9
zZHubZOSyNEwue4yNFi2Ew==
`protect END_PROTECTED
