`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rIdNv2BZ2z05CPxzykMrtb7HKMMx7gu1sGl0kZ7oja0uP0mKCdLPeEf05cOOp03x
bbn74NJOky73fNA/Au1ky+H9UzYwAe66euYYhUxi+Hb6q7Ckd29Iq6JJOvq3fYQ/
lakBzZDYtqQBePbMcAeRhyercSI+qX+i7uY35IISSQdWkCGLIe2WbiIp8UuxcHH/
HgzPQhOgidCulDVfdJ4YbGbzjHLQ507kagU5A7i2p1OZm/r6iYeXcWb5+kX5jDR2
HDKIhWNM6lW90deaujLDPz3M1sxx95v9jtk9ge6prkgFkJp1qjMTx13ZzEPCZsBA
GW8yJnwRs0g80pae1dGxlFIOiqnVMspNL+3T9PCExpruYE3AF2+yer0WCCm8Xcu3
NdWF76CY680SzeYQLy3UpZcLgwwt9uAbHpqSwcYFxEF5H2f4qZzorxxfBWLgBk2U
u474I/7pe5HZ83hkDDWIfM+0PEZM9ZqETDejjRxZXrw=
`protect END_PROTECTED
