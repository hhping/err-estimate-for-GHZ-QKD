`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8dULJomfWZggMGNJ+DCy/U+FDcW8JBOlasSTOhdnqKWPeEDumZRGPVXvWQH7bloG
hAYbDtfythgw4d/qve4GUPs+Za+zPPxSnW8SE3RS0G3NqzGjKfwf/tNxzOZSrTfs
1YsgHIzSX2NYJKLP8xoDjHXYBHPQqnUYY7LxuTqmeHDU6Mq3XUyKFXr1Qm1vAlVH
5iJ80Q0UQZXy4MCbU5H/Awv+mG7C07srxjzcz2AUMqXeN8KNIjTCUAY7/uyYu1db
2aPY3fEdQAtyyqKx2rSe3RwGNZKHkCCy0czRK7zaZwg1Wd9Hv2ijFnGl2KXi7Fl/
Hr5Tumh2VrEv+GAu99VEi+X/TTNuVp9WZrZ9M4ASH/uQpZ4Apt6B4MUBgV6j+Xzm
AdZfvAIke9EiU3TQQ8ghENREFfl7e3QfInUQnRGbEDFhLLDz06RrxXIhwGGdr+Oi
gGMayIE4m5a4G1jHbYEbhP5FNeLsLyKxtTZyFn7jdKsnhtvuElTTSot7V+ETLGb2
/6nuTyKPuogy6k6jRnTprgrHg1LKd3UCy6wupc9OFJ8K8mtUDqzP6lANk7ZnsAw5
sFaoksF4PCsW3u7mIsaUVhbOgq4DXCBCfhalS1Og8P+3liaxvm2vOXAjBaZnMDlA
YRRJY6BSzDz1mixI4ecdB2kP9iRvAa5j3+pRj/LxXLAvOvCC6T6xgKeliqIEqFMb
tWu41WngjPnfHiLDt5XGNCPE4wasdCUg4jrkDM1+Cuasg/aG4kuA/7xWcOOtlDyC
cmV0Ycj05ViOJn8l9Gm2Ni0iVlRsrNwn2/4HqB2ZsBeOOkLaTCmgLIfHQW89Fr88
cb/CCHrVt5s/GArLkqBocVLmMmGw9G9uAhIR6TwECABS979aZAY82/mPirvB0Ehs
HeToamvUablCXBRU+rC/Ji6sACnu8HQZFwTXm1+v/7TgNXMpFPT2xhf9Ra4Obkcw
87dDevjrEUaxLiN6r8cq3+7uzMkiOJDAg5+UnIwfWZ6+QJwltNU45SzhwW4EUQ8x
f4M2rlFqtR311Myxri68MlYIr7Q155DzKA6w/+VNeErTyljycO9dT7cJPMzFTLRJ
Dza2uZyz/wnlMkd6kAYZV1qVrEZCrQaWZ3rPDwlMa7T3qjSWLPgAwVuouMK1mhNf
/E1MAHF13VK8M/t9bM9BfSAiuj6CnAWORcNdCFZKy7L0YoWhK0qxIITvq3Tff3dc
pV3VUIPO5LSzOVcjcIl9gI/RqdOi3mIe+HbCWwSYuxNVaDNc3KY6T2agxxoWfVRf
OewG1Z2OW2yOFjU75NQ/vfZTwxGofJ6AVtOuj7UzznUWU+rz41nNGVhMJbwGtgnc
UIX7DaeK28E2UYmI1Cr5s5fQoKTuTpEpzZavnCAVwMqTf3raFJq4WesK9CyxHQfd
KCU5AyYhVsVE8RzwKZnIww+kplcni36mHJQon/sX2zcVJuVwP0PXdtS9UoCgEjUr
hxkKV3pZitBDbhGoDdCS+IJe/DDp4CCWG1IejdH3Q6QWIxL2JGGzqzXAG9KLp+Tm
kY7ay3NvMLSKgKF0hys8EzM71s3bXeKUjO2eVn1wGW2fTUI230xeesMLPMyKoMjS
zkDpWuT6CFnIZ3Sr3niepJ3B9gTVaehPyvoz3I3hBBk3x6iZONoduJVOtcw+Utny
9ibs5XjfrRM19Q49Pnl5gZFU9vHZbvISUC07k5OvW4acpIASbiimtLAR1ZTnUW6y
PGpSbXFWn930v9B1VdqNig6ms+VWUMXm5XpTBLfPb9bREPGT2mKEUkPISKi9fvk1
PAc8Lp4GUU7b1W3lbQKDsMCUb8aFBqQ15TLSbFM5zCdzKojgOyHkigtHiB5EPUq/
4433HN3uzQS9I2MI+xuVIxAEUxgs7vDp1Vysd138/iKXu3S/X30RPLNQjscr02HQ
WkHtyF7dU1O+VV3zqxxYKv2NR7qCN/6PCjMhwAVSv+A5kYGHkdLGWtVyja05sJBO
FZW4Hm8NvUBHdd4qkV0uX0zQ2eAZn11+5bTdqDZocDjAHzniYWitxhI/+N5w2u/a
nWENFFSshFJohpPkTzFoKZgihhU6tvPVzEMdieg03BSTwGes8deNCeimyo7i/51k
M8AtLE/yElDAxMNqKFqHkpi986qZiKXOwC2CD1sG+JWvzJDIhYYKYruWjoXcA3cQ
FIoTPlBTDfQZHOoJnIrHy7Rz5iEyjrT4iwH1dgqfkLd0OoI8g0W4JjzTH7xpeNEM
`protect END_PROTECTED
