`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VHYUJNfQPgMy09eK3tfyo5ijVP/8QClV9kUN+0xc2fPK07EWHgpPMF1aIOAlOSmg
JCInF1tswES6hFHUynTmVSNZcm3J+fuTUJIAv6+OexT3NWOXcmrc9Dis/KvOXaXg
3Fm3/MER2ldmYcVCQ7tdJJ/aNP/I5K4wasxsUxchmxOdWkserWSij6WG32gD+0tB
IQs7mvqtefd9JGQJ4LWgu/hTUvtLfqEurcUEHyUjwysFV1CdNzoGYt2l1POsmhqT
r8zxuuQdXCP68J4sqx6Rz9GIQ6kMt8IeAueLLMHd2Zku5Rnb8LMQd4qftbd8/ohc
U8L0u5T4VTJGNX3f4vuRrIOxX6GIpLZQ6HubqTicNq1MppQdOOOZdznQqY6lheAR
YYbnp71xq0F1+3sxnro8mXBALLgl4Wfwwd6fj0XKaciu4FiIDMf45RXjAlwhgbYa
C9SnVA0gqbMzgsOLKYRvHD1Oi/IQsTOiYJxvRUR2d3XmcIYcgtBOlrcwprni+lcF
WUawwhylep0v6YKmaqEVg1UFqSHqtukphawP/RyOWVyYefMChteWwdiIJ/c+sfRW
5T6QZkesCrW9X8XTKILzCPkdVdwEpbBK0i7Nlgl9DSgOcN5Tu3vYK1yyoFpizhKK
zbyG0uPgwEZSJmU0hFbXpKUVFpf/5r+JRQsKCtzvaPUy1U1CiOE/yoruMxL4AkFk
ouZGInYLbnwD6VYyXZPVv9R8emPk59ooVy5bgXX+gP4VZ9qfHv1hcldClS7YUgC/
+qM5s7UnLb4BCz0xnJfB0cme7U0o4uvIDbgJAc0hHdt9KwVqqK+9agPHVqRY600X
sAfrgvngzg0fjA8VfGib0X70fwI155xCn6dTnjHekJfJvabx6jcthUB9xpB2UbbS
LjBw0OHqv3SXtjxVAwYNZtRNMSxfSf6zjTrCMZfHtUso9sRRTxbmJTKkUXh7pntY
huN7T+2UWihfEW57DGPoXc3KNrscxEZdf7ydvNrNvqZEh0mdPlEXVYKu29bdVtRI
MsDuiZKG36rod7CoI/no1/kURCsrBNXeU5JrOOcaE3ECxA6ghNMs3lJN2SJojlt8
Aky1qvWmuiBfODzQ245N6pAz8pD1siS2d02VKC/clSKX6nvLawHkcfaIJNvmUsjs
GJUf63/fRS+fgP6J7FdO4m6t+c3W6Hyw1sR86sasgkyi/yakYfcuQwBtO2Vdm4ST
ZE1RvAx5O8YcmXcSSFoANTMIeplxq8LdcagILLXf56W4opZO3vwaO/KUqHgbW9jt
vEMX/ub7jKR0lSYgXA6vYOxrLZNoP+jAwL1tjtiRD80lFy6kUqjjYWt1zFYec4Gb
skYHp9qk+VJXxSzv5d/LcdviN0OF2LaKPPAcz7SQOCZrNOo0xQqa2cxGOHi1D7Ma
ixGEDLiSdlkFRkqO9gLt6u+QITGAyULHr1QxEk78zmTGYCZBkCkweA4yQ4Fokmbj
k8XNbP+nIIe7sj7uFwdJ8Q==
`protect END_PROTECTED
