`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wosTN6m3J7LpNxeDAiR2zlW4oJQiIdBo+el/0mpJoJ+GQvf72AuVmmlSxHjxlOLU
OrroNocciwkY9sg+efAok4gqQfIhfYdLvgtA7T1KY1asspxmzNYdKf95t8/zM/fJ
CV5BpQfx0vpTFIHWhnjPJZznv0BB04YIl6yQzNPxmlnpXcaKe9jicxFDtph9U+I2
QPJ4bUodw6du8wnFACC34stChqe882B0rvXQWFRuzMSF7NOsw2j14HwmTh47Vaeg
7/Cqkum8sRujjuYjem4ErSIL4yh4TNzkGA1IYg3MgHl17bUegHGIPMhQUy9VQIGH
8iqGY4M/YfUTxvAGPTjxuqshZf5qiKm8c5kSWwvDcFSl2Ngf8nPokk0jZbY2rjkB
JCgUOwO+AYhphCFkyYHjNOdmEdD6jFTl2BhPyFJ/XytW+0zsK7+Cr7NmbI9f+A3y
IWB03By+VKAF0BpUZCJRA/aXWLoyFEiJeInF1gkBzhXBQ5hmiGZrS6DuuzBeYBox
gjsQDwjHnXle9iDdpjbh3CqKMfNDIpn6j4dmzbYD9bEZVxxH5bH9evLcbAld8U98
xO8BdSmpozVMMwY4OimNaXeobkdQudksrY/zzpbr2MFolnOdA7oEGkZRbfH94kqW
pZOO7BW/7psCnbBQHT0el3bJo34Vg6aNzMUQJ9enS5ZgY+Hs4EqlAp1kWtMVC9wM
rUdIMY2rDWdI3F5otDc1BJDp9EzJ3ef4IyRgSLdmFEc=
`protect END_PROTECTED
