`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HV3HBb2Bx0FXEWscYskTqHnSR/1YNjaLmGHMnOqdGCcg7ynCt1nT5imIhMKD5vig
Jr4sdCRmic7o94WaMGH6fh2ji2sSKwzEXY8qH0wLPzkNTWatuDfYD4sG07RYNNOb
frMOXxzy6AfMnTra9HuWDHcyvq6Sny55sQG57NmQ9JKqgUjfOdxaT56zhMyM4El9
8Pn8GeCqoYY8RoYUC9+AgeKAUoZQC4GmtztTRc82L4OEron4cvIWSItIoukRVP9m
2RftfK7IJIksuzWyCu2QD9O+qFHuL+rDkQGjvT4DOAlhaxcinzp7Jjg7Uqv9rPUt
IMTdhHoK7Yg2371Q/0rNvQnRYI/7JS3UrTFKYqwKXB3/kJO4NA+W1MzDuuapWiwq
bbFZS8Wx3DKKVivR4sdekKWjnrd8dm+S7fa/KsTsqo15vxoyE7/Px1Lc7DkrN6s8
OrtiQVQ/5jcJGfhqnP2Ayi2FrRqyihk1cG/dgOImZhowHO14fgImOZ2LwHcS4frx
0Nra87VJPsx619lzZdy5zOeABcejh73fX+CMPWHnEL1ZrrsEO7QPG/ntSgS8OUEo
hKRK8TjSy5b/FVMDnIhGMvCSISvNCQV7CVg1zYKfHxXlPvzP+0+1NsZozvvYcfrp
bbAjUI/w3NQs15IsdmD8pXmvsyTy6kB2SXMEvLGjLY3N9jRAV7U0OSD9EQlIZPwm
AsIcU+7pqR5uLqgxMOXtBIUVfuF8791Q5n4yp9NIdJUwpjrnHOugD+oFAp/mDTxA
vi9NoJPQ4aUJ/yx1/xmtuaNr6dD0lhbxtK/S2qTrFfKD0mdDihLdo/knwv4VeZVP
N0aNr+4cROS1dNdT5Pr3QUxVILd3p5gPc04fKyaeEnINQQj32kYNbJOS8ZC98ILE
AenR1MJ/WhqxUo/jxZesiJeR2+xOon37fA50YPxII5XeZ2syo18Xb4wFJdR8TkPl
PYjb+yMWBCWHVlO0eXOBZJojQ+L2scU6Ma1EUZGNV9rRZMDXBU5yPtYLzEhec2Qx
YDQLnkGvtPaqck/1drBGaphJ5497eKhfflFw5PbXC3IOnkwF7/F3NewGZJC16piv
zZuWYU6UpHSBzAUNWDjV4k0mZTUe6ue8QQ/eszwuBh83tioDqK+vPcVbQPpdrA4Q
G7r9iB+ZJlTx9Vfc+hyegTGOm3pRi0L/ItF/QglODEfEkvJ5878aEFuMTnfrlacQ
iwGcIYEwwk3vWNnfS+6RNaNgZGeZIm0cXHYj4W9sFcm11F8vbDqfYmGuyTjaAiE3
gbo7ymufUTNTzk6bddju6efA0iBrMyoteaxd/zJS4784I5wOSb6Hr0O3MuCuFyPt
EqvmgBQd9Ji2OLfR61QcuIYD//b/ScP/hYxJs2VhvyDaYop8oriHhL0nZi2Lf9aA
mGHC3cFQTn+Iiy2vsPT0DAF72VPNJNXDRRc3hn3Lke2fP49kqn4817J0iaf90btM
eypUFzi8GbNuddER5cPi5W042F5xR1yXSAhHhM/uF9lQ8HBrjj1hrVSp0OkEd9I0
aA4mkzJqId6dZ3pKUTM6+LdEWrLlWLgkCZc9Zs1lBNcx4eGKqTyvkWol3SkBA6Po
78m9XGUXZYCiW55wNEAei2jVKTosB1RdgeiE47Iqc6IInHnyRXYN4hGcE7Qwn8nZ
oSCMFGslKGt+8tcjWIo8nKt8rJF42ICqZwacSBTh9N+XyNcTDr7/OFwgwMS0+q3i
pB40A1gxOpk1e9mgM7t/SNMr81pUqvMbeMMUCQNsRxkqtTv8Rc9HN4gevKl8Nlf9
0GozmxsdWLlB67qG2LpdoY96U7HWJUfbdpu8rAyzqK7mRcpLJukwFI8lUEVFCYaq
yECLdZQrd6uqjWuVhEOMydKWBZ85E60ipBWbNQ9BoETQI8ZzaKBoTi5G/wnhJ1nU
tN7LyVnvZvt8JCtIVLBTt2hOodRc/M/vSnjr4LiwIY7zUNgSmthkG1WJs43ANOrf
pN74IX+2TcJ5LpDYPCc0N/cczUR7AUcZ/VsdIDowkRwqnk9TopJ4GAereDxwgOyC
X0+JEjuO8qV0UiL9GAKQ4sXdnuRRIJBfMB4UEO6XRD1ZYgC2CsvXcaJj4Hf1xYov
FvuSuu1eXLFYBmpPpgqG0ZPuSHpTrjrPpaGF4SVyuHGv0jnEek0BoCLfArY+N7lu
NE35y2ITo/yJAiwF+EH3Otavlljs5+8oYXPCuQ7NsJMwesT++xJIpFEL59cyriYj
KEfg7fkv+4aPsofztkvHifduYbFs1OnHpwdfLQx5U4vc5nq/9vkRlLSUGO1OqYSU
aQGvekgnTtfglGl0zaStaKacynTLeKgClI4v588Ej3Nr+AOy7JXjK7mvKAFBZgcn
UMkB1Hla+jlFd8A1TISRgM8tfz66dS7RTVugoJYx/q62iSTZ06YMPtdji7XwqIJn
qs/opY+VVNnOUYosec/w6lGzaObDwqt8hN4OnFp/lV5rgeKLmFWn09IKS0RaAjVb
aK5JEPxZloroQHyO1axkT6m2HoqP1EqIQgkZ2Duav+/Uj9KzEUrzXj2ly7WWiNm5
b5HWbcZHku5CMFPHwa6FOdEOw9Iw3iprHbj7XceYqA8AofVDR2B3SpBb1CDKeCDg
9R0PJoHqHYKBqxGyMMhfhjrp8MCh0z5Dso00mk7m/REXk1Pg9tfDi/bAPpc6d9Qe
G6vhaQ0JgHLTpXCo6SXolk+jJ1Dywvi3V+DXRyrKqZfoR476dSQ4OjjgAmsWgX71
M8DCnbwPoYaVHX6uHVoMVFdyX/gkP2IF1g0jWgvcxXdVLCzPYr5O1kpuBdQH/9C7
soNv6RKpQG3ZrWeD1SPYU7Ph8GaGurQtOWh0WM//q83SkyzZcEcnS3kr0gEbY+YH
AFPwLsCJsxD0JrnV/bH540k0KRuiesTE9XAYLQ5iou/rZGfdD4YMfoPGP36Hsw5d
M8Xu2gnLo2KfdqH0Agfizz3jqSzTm7evDXDnvKeQFEvwdboygLagS94yDB9+Sqg/
K9NLOv061eEsfc4WCPRcIYq7tbED2sHPcg6XodRSOri0hfVIUhepRa0SZkXsMFj6
Ny2Jl60c7V+0yoDol34J7QtHRElg0M+QbZOBLN1B4/8l28fjIIM4pTwKmkjkFT9d
X77ZJOk8JYMkdCCl2J9tGsmytny5PrQ30k5E4LKBj0JHBzZbqrMt4HoR1ZwyCwoZ
xe6c0dAiYBPW2NMdJvaB0eNyzhrxyqtanwQYeXKTsKQPw4bI6HEvp23MbL5XqIAz
rY82WaLiWBwkt1llAjnkbz9ShozTM69uppW1ZMG/cYZnisvuHoAKAK3Zhic1nNFD
kpI0IjQUh1ynnKDOka/wla7qe2OK5KHu36lL9PoislaJ9TytgNx3zXx1/BhwhOgA
uI48sLye5WxVJAcBJIdSHLNwcfSZshi+QVF4bIJ5IB1Il7hTHk8WVules9DCSAqY
J6tJet2mfX6Q278MwY/Z0Vqz3Q3XBIiPBFKl/GySES+uQv1wHtOl0o2rfAD0KMwR
TEOERxwpItKnUgZviU2Hbp1UAekReqTCLLn+ND9A87Vjwz7Uy3j5bXv2JE5OLY+8
B/dekQFRz/mtw48MrLpDFVYnG2+WQ3YW7Y4haplASZykXyKvKR4z+GSSBi7X8mLg
H+y14Iclkx+JjIKI4dBjuLtEoVmuaq/lkNyO2OLDt3fsxH5uISKFdkgZfvDAwtcq
Mymmuq0PIkhMOH9UXNhYlkEVXeLBh/3Eijr61qNv0ZPBwqdwQwtzQEv4bOHVrTXD
Elm6ApCoY3tKGXMS+K3ato+86iCZUwbpzr0E6MEviWjjcfcVgyTInyglt03iF93k
OkTF/O4vz4WL2NqmJPgAniRn3m4ZgyWguNEsWoDT1dG/Cl2Lj+3jRZArFHYxpIkd
cnQhjwCNSqjbKPvmS45v5NjiU8ubBwwkie6IRD7b5aDvAOJarMnc52oyX1ERKt02
lqDR3ZRkbUGUWTR3zW2u5V28KLvBkIWuMar/jo6k/VTKrTj3UpTULaMRhUqEYP3B
4ZBJgbu4iCMLjQHfY/ydXpTa/VDYP5nfOCd9pp3rzgxekdmbDqkWSL6pkD9Pzw2B
QVEJ58Xoyvy4eQpM8dfrpzgrxHPyLEEkxpCbVd8jdSrl1agxH9KAueCV6pwtkhvH
aDMIE1/fGZVj0ymUYUUQbI2e2TjO/Kgm3T3H4PXkmL1Q/shWLZM8/P9sTLZb8Cx2
aLv2EcqN7C+rDVvyArUFPiJx2g6ztMfIbvlxpxpynC+rTXf6jFPmRL1YK67HoL+E
s2pLSuGEUxc0axin8wpxZcVLrNp5Gfrk8Ym2aEREL2qMkKH33sH2KFR79vS//DRk
enmvTqr3RANpSvMCHrmET1ETZW83cWh33jCuvm790ly5L+RsdgkAjHDYTS3t4Wsj
Ux5uzpycEpMJiiA3w6UjWd9VKzJ8NiYnJHmDHNTAU5vsSzobWWGlJIgc3eY+oKVL
jJ4KFyQx1nG8C9j9VM2rcF3/jfVg8HTwp81ell/P86OUTiSx4FZuaX2zTBatsbvV
HGRpXjhZKQydrLE8uZpxVSnvvXC4SDjD8c1VnrrZ+FO6+e9hV++Ac97g4A4gJ03z
bog1mm/243EKQs1WfUBIg90AiimltTRK2QXEhsM936dL6oNMTSJHjX8ql94GUqhA
HsOD+aGgonF4bN1Slr2Bvx+DLUuGbc0HHfhbfQAyzy+tB6dOflA4hn7A5crGolkY
B+FE/IkszX7oapN+ZupdjGHIskuo0H/QtkUtk6JXnbLPf/eAaXc4Rq9iBbwVcup/
/n247zb5O7HAopewwq8vSa4mPPdcx7jIUvdry/1HhOgGL7nAxh0jImrcwEIdxu1g
FeDbM01rNgGyaVtc6cP0mdO9pmFCw9K9kZha+ThbBR7hAiAKhWKwbUlZAVcBylYX
s7kEpxt81INZjAm4dYA7IxWY3eXYZhBD+/0b9gnqwYj+iG2pDFD22nNM41MgpkgA
FeWOEeSNSrsPk8ea0IUapM558TNJ9X6Ew9DgtWyRjY34jJto78kmUo5/bCNNA7R8
NRzzRD0pF0S+6/V/KTvDlTVa6hRzTFH5n9AM3Z+bVJ2QdhfxKAOZKrk1hUmG5LR5
dIi38Q8iTyXVdAJH3XhsrhHNKTaMigvrSHgurOEaiKVAC4ZzYTsGnyudGTwZpRDg
mZygtUW/93vuQwrcv6rup8cx3bLto+sYqKcoDOSqOxG6mpDgcyhtASQovVSfBxnJ
/HsYB/uBthyqkrVlj1ey209hW3Y88DxsJPsc3erp9qkPBlaVhrkotX4D5ZY85rhe
nwU4T9rSb9YrH4OVRMu/a219CcGbcm7bB+REquKYlMs4cKBLEF7FKrHKl+OmWikz
DbLY5559GlB+CXjMqAQzzRO88E3IEhFhpz/cpisJg+x0xtXX84uVO7vzsaInHKhC
fw8Ie9FPQQW2JAKeK1HVEJICxzfditS6y+/nXrXRhuCXP4XR2zJVyjyrCvvta8/M
3vKRk3gVHhqNjjckVD5FwmmmgmLJIDANxuMBKNbPMVUV5tEDNcCjr6ZYHf58O77d
y0rwES2KvBoJeZgBZ82Gh4cTokmNr7spnfyJn2L4oRuSxI7McgDUJibKVxkft+vu
4ElShoNmjtwfapob2aP+xxCuyqvFV5Y2ZFo0ESCxCXY9dlpoEtEaL2qqeCToL4Z7
E5lHFR/Cn/dQUUk7l6O3EK94QqBwP8TDZyPOygz0jw+VqnAw24VZ+j90BeJlLZKC
rxM7GRS8cy4Mq2OayMETorGbGnYTDP9Egsfp/6k7bP8r8cSyFnFfTt6LwT0eGIiZ
EHV8K3vGl69go3n8esGUVS1ey5qvlLTM0glDR2Fnb3wDzkJM6fk6vjaksTKvyqiL
sqV0kroqXp56wXysHxfxtl1ACfdXRHP8HkB2seRFX8Tthv3Pl7LhwOOXUhjyBmSo
IE9UJsqMIwMfp+s7yoMTMYUcDEZ6Bun/i7UNk6Xxue5QjnjTOr/5WS/C4zxX8hBb
R/v/A0Y2UPOAXCdXIhp+rRfYcT2Dz8KNZZ96MC197+9wbuDvxga3fmpWy1DVXaiq
KkPZ+r5pcfM0hBIKc9wolysE4JMpceCjKPqLaezcqneQo3fCo9vZCCZWyVvyzLsn
SmlpbXbxMwnd3RnMF/YHnoQ+hSevkZqRCD5aIR6DTLTJZKVaQpUMlJ9fXKiAlCYp
lCOIBW026NzxJ94MdCKmklul9agz7GsLAAx1xpNqp/mjksM4IGk2u+bmu1TJ5j7V
SpThMCa9O0PaeMhG2LvAnBWTWBXaHj/hRtq/LFtWq95NYNSymGmNu7azMjshT/F3
BmMiXp1PHJLDLDNbMawI5Rai2104vIe1KZW4QABr6LMzXxj+WIKEtsHihTKEzAbC
aJAdLmUpdrtGssfmPcpK82z670Dp4DhlJkgIuyoQjoENunSsEnUw7ICbZ54w+fk6
ZmcHRBh9ApGvMxY65TI/3P7OFnuoT+Fy5kMj5bM4bDm7SxiykS8ORCsYCouG960Y
cN34tiQrzrLiBQzO2f3DeH83Dip/8w7bOpNznzzQhQcuj1NyITktFjvuu2M6G0vp
c7gDWD5c4IX/NAcSjNRjTWSBEhuVdEaQPwnV8WAoLYGoh0gvNDflG19OlO3TsA/F
CiELqgCo8jnO91e7pd/Ox/t2mUq7sQYDnIh1h/6THYdAiidGzVFD+3dJ/a5rPGPo
CbfC64Q0BE4S4nSquzBmO6o85f+uqWOuC4y1BxdsQr7YiWnV7RCMuonVOAfyOGFM
5E6gL63YjK7zujm4BE/IF5fT6ZXeAIjj5LDLOzwnyvMw954lwfUeLIpFQE4EIlkK
tCPVXVzCInjImyi8882d2srOFQNib9pj12hjVpRww9wM0ZLGAmCfv7/m6RgmFSgm
FNNloiqmo7YIDlWuy+Yh1kU27lh0pcaDKgi9T7PVaS2G7oUusRUMuatOxRG+YiOd
sbTZBWogOGIH7ltAGIiQR+GrHem8OrDAzaozIQGjsMUlXoqKdzdk957+Ge//13rs
QsGWjO4dLm1utc0fd5Gcgv4zoDSNKFnfw20DF+4Voi25ecZ2EUQq+MFQpkIbyHia
1rm/bPF3c7pN2/xFlF9tsI/Ho0K3H5ufQQKaVJtJ+AZQyCoCfEXbB+tShNYZcPTh
El4EPylBHNPG2pr1Bi3rioSBYaX+fSLLvAjuj5OJPBxZWdRU32hWzb5kWt/fP8Ak
iqBNLPXDV29yriNT8mxwO4cHK6FHazr4w16E3ZOjiFogZLV9BbtorCDPxc4mQrYG
0YAOI0q/Zi89AkGNOxddSccytDmaJHVsoEGiRIfTzb9VLl/HJq23NQ2Fd8PU6s/e
XXLWTYVWvPoHp/zxtkpMgn4nhbiCJncja9Lm4L5TpR5bTKPS2CeAA220x2685w6X
yZNkU/AiBRSNhS3u32mz/x5mOrMeYj0AsGcakuaV4IBuOa28wtDwgBKtdGMhqRER
Mm3LD9B4SkAeEFGWfNhgYqyszlAXQz5/KbUymj71nRJ8wQHGhsXy53HHCMubyGbH
1VmmWsogMUPx2YUc+5un6f8uySZxD6zJoPjUR0Q5185ppWcMWOS39CDNUutE70Uu
SWEBgNWkIhmeYk174O9HnbvvwGO7QwCzJGolCOTsWc4C7oCDBE5mPy+TZYVYs19x
cH4PCBTjM9pJQIouMTh3q3hhnplRggJyWsqvCILly/u5wW78ZI+oijEOw5tazkmI
8ZHNiP3GvoYlK2MWaVVxgEBqJIL3NoSrAK9rAqgPb7Y4BNqXOfHwdzIneFlTa4qJ
+KMG9JQw6T0E2mnOArX2OUa1eOwiGUAayd8UUuRnrHg15knGG+G61VVy1m+YNeHu
Gebl4hlvPvPatJJUYaSOvZG5BGQFGsvaT1/2Desm+GA2gsHOOIduQce+aHnJexu2
GIiOnRbT4G46E6k33oUODjEwDnbuWk/v8QluGFbRphmib19gG+MRZ+mf7Ri85eA7
CAo7ljspCjuOxU02Mm++3sNcABRUuCXAV+07m6PksQmY1+BIcj13rLzG5xEXVDmf
Z8Pz8cgabNoBhKabtZVOvXYjh8OlQlDxOwFmRu7Kcp0Kh8WaQkvbkB9FeNJUfRyu
qvWwbRRu4r9oPKtpEJgvKepK4SNO5geWbtZLOKK2sGK50Rd2qR9fDPJpfQcdbKEN
H26ctqbGxYKef+qoc6hkbQDQb7h3dKkKnb17jpK+R/dojLuQHYxE4WEEz4Rv1wmC
7U5PpbK0yXSzpfWfCLfbtYhMuovcCd9q15Gsm3BcOsHNCpX/oLAS5xyXNXbBRVWO
Zwr8aZOrhN6xiCSxKuDO/UR4262S7iCgFCRfkEW9p41punyHUQcRgruIzz3tbmUs
ZOZjQcaStPodGlxlI8Hx2C+uFbB3P+CqoNHNQZtj/2kRh6RwubMsPQW4Rq35fyuR
Yrefxy6JqhXv0j8iEDRU/mfDP0bGREcsR5KCjzFt307cRpEfwBxbqcPP1Cu4kb0Q
m1+EAIf8O7uk3VGkT6KgzyXCGzRHL/GUg9DLUG3eK3xUdntjHzDH59vpojGuUkUA
u8LfFeFlm/mS/EVoACgHCqKm/Byf9FmoA/zjt3DpeuDDsSntyXETyrYE9TK5wZUz
ZoVeLxLlVxnqFyixrTsWmb5ThvSmJY75J6P1QedkEtbm8wsdN64xNlxn54Xp4Z/p
yoZtJs2UAAPnRU37IoTMLJt3EAiTjj08QP3KjNbHCpUOtp9HPXMU5T392CyqjEor
ndBCIFVleV36nSFMg8FL/PNWxZLMOiiv9vVYJVtw3ZVJPbuM2GMEMergALXG+t9C
c9mUOUeXfnkpt96BPVNffWoXR79jAqd6629YTbV5h5SuqxqbADHxJy91EYnQA7Ty
xknD38Ee8EVfdCPAzMsbJOAhbA5v6SW1M+JnQXd4EITRB60sjODVb6Hp5seWiFuP
9DN5GTVvhDJV5OjTMsefECQxdOZohmo/0RVfzx8IMuYMyrcq68VPs/Gvi4NfgOkb
qwOKyAX/ss75rYU/ofqj56D2suV9eApxndQZo+02E594d1cZWLuJIwCyrKY8aTqS
hzg5bCpQbfDPge/DN78EyrRYqX4TFG/IWqjvsCxuLKRFGdWm/asZiJgczxoN0reS
m/UxOgzEweZ05jyXKMC2s4O+psJJyVZpwuajQ60eNnQjKPzQgmuOE8TAzbM1bE3p
1vggFSE4Sy9Zm7H/KzD+GNkdyUg+0gzuJ/Yy3zp7TMGvXgGutSqHOSUpthnX36cq
QIeWJUZs8Mur6UCvok0mg491bUjJ5jwkjeIcHzbwOAYQcZkNhBz7BkpO4uZs+Rde
QhWnGwXzSzjDBn53Gfy9LRwxvYqCMY7tjNPwTyqtDqa32yaZZESYviSq+QL+/OAc
ZgWWuUEre5AIH9YCI0Vg0SCbirqrMqb77bxdNgdWyPYNWz5vnAtsSi9LPrPjmyX9
DhuMI1MaUA5EnFUtl5P4aHCMZZVe6gZ9ZzdtK3oaBXq0QWWUVEpTrH9MUeaOZjP/
FIgSjoNyZ9szxQfC9VdrGFwJCaCOTOeEr+3s5b3QLGw0+w3QbUfuRWcySpoWaR2d
Ps8TCRlkCnXY2ropU9LoEZX12lwBh6T2fsS6xDJnfFEeEXLkXeY/nOVW0OGx41aB
Bi+ECIAmL/RVfO3D/zNCA47y1PJRvdqzwO8temlm8a2oKuSMq7x+mVz1AlJh3BzJ
z4voA1LDEAm4CLXELcPp9gC8zgvzj34gRVHR+7K4zwnBkndXy0nSJ3G2PoVjBMgW
7v77szY0E+BIplcuPP+PuzqEIbU9vp4eID2fRE865NRh5eI59We/+Kxyipeyqh+D
3KpgLYXZbfiqaRlItVpQnfqBVSv4yDREhBjNg4VA0bYiXmBjp1VKeNrMENwTSmdw
l5TawppAQDgU92cmRZCsQIWSaURkkrgD69XSEPPuxIeea/rdj+QMq3voXG9lC6D2
RQ2wGDHgvhynPte5Pz5lMQI7BZ+elg3ueVaD5YlLeWmPu/DIfEVW2zmvvHEbEwXX
uANyj0BymeYLaMMVG8gmSVaEbjeULSZwF+Q7d7RveoJjo25j5JfMfa5peh+DCj+2
pH9XFe5dFeOyBV4V9XXSqGwg6JQJYzwAEivee9/nuyCjsEXomenArqsXVJhEkWsk
ptmkfNJnaYt+BHzlesNfgecLoK1YIvq5YLDEtxmqUNUUltO1BzanGHID8O2xT+LI
AhvYAoaQCj6wdha1BHRDk/OIXsIQa+dPUDndJJoe3owZYiaeP6yDW1mw2j13mbuo
VGhP9AKOqPqzrlcoSLwrJK+hCF+DB89apJxRpCAf7iK1EF0qpaYFoIHXfq7XU7+E
eZ26Hi8LfGZzt+atD87YFXtnHQlSofgQ6AkpocQX3fYvsLd/TV7m1BM6IvD3zxzi
kUAWI7oMnPYnx7rOCgSZplvAsYkfEyAORzY1B3cGzfaxPFwdO5W/rrQgwbuAHzkv
o5jvl0W01Y333itQJErriFtWTCOc1xlNOgMQoF1XgntfGCxukVbYNAEGj9TLIXeb
+M/Idx09MNAR8rDAx0bSH5Bs0czIylisJ7n6vAsfLvbRm5ewKk9+qz78E9oznUHO
AhpIxMJ0HAMKMrDlA1IqUoHVLqNxzW50IlpwhzeOOBzKgDG1XOEaVGba3XkLvgwR
zeSVx0S9pWU+wpMHl8//ri2MoxWiRC/MuPM4xJUYUz2jSPat2JuNWoiawCna4+hE
K6chISPY9/ckygzVHTIjkJAKueGRg8FNrhXdomc385OSZ8xoX6s/s8/U64BNLSSo
79fFQK307yrO+0QuafHUX5/wy8TPJnBRTg40sZoGfJctsCxFMxidVENCu8BpgkOt
6KZ+3shJK1eFpvxqfyAVb3j6QaKCyj8bjPGAPzqI8+y69wJWSuLaBa7JYo6NNC/H
K6KT+Y5/PirvwHH3LNDR20+UwepwKreXptJp+sE+7k8+iVowCC/+LR113Qskq5mL
iqittn2oQzFwb+dcm5BFHDG95U0lL2o5ew2CZC1gznTZftbRh1d6IWmebPOKwTGn
4nlgQXpXeSu862zao0cjbXkj8qxmOzpNqlAkkOWDznfLpEL+KCBGPiD+OD+dnLjT
dt/f5OrRlY1TWLrIazxUyFAfJfhBXZC+Zd/GMgKy9jnRvYVgAlrtBvaXw5h/+Xrm
PqDA2bdYIUit30eH1U9wBXFS+Myr+9KviXKkpH2HYq21FXtDglPTosW/XijRcGXx
mkWL4RIXw0+2VIwSauWEq1QoTAHXQ59OKMtdi7s9PVDZ3fwfxHYdyo1kYkY7sOs2
YILvy15wcT6oenEThcKi3dVhOfNsHwlChH0VvbmWXdkqjOdXBujMsyMVENrYg7mZ
J1ixSeDoXL+i55/UAJob6CUfJv64LgVMqKrOL/8EubaeLnb/CXkwdQ540D16mJ5Q
x3IIhrPU0JmwxwL28zYLBkw/0BjQtstHm4cNuw4J7yPuAk4FNKrwL6Hn65WKUoKR
UpHMHMQPBRX2BzT2/QYxbq70BZWrWrEuowkwm1kFKoOqc56KeaQjilUHsE3DhTL7
yYqRNSxcuyp2QJ0DvHZ3S6iLQUGLqy1ns3swiTuUA92pvwkLM+Uh6HoSFlEshmTb
sLpqEVpAlsxVn+Bx0rwEKjRR4RYB5pTaHXTlo+mjAOeM0w4Vy4hTrKFjUQFRdQHI
O73EBlQ/AZ7tPnuhIEhHhQwCD+whWNiwRyL0qy0iJEzcuiGdIjRRKrfa5syVdO1T
fKXEd7PaI7cAbE2EiC9Wq79cDpOKbl3hfhwcd0mdm+zURgmxE947c8S4N2vrEljJ
ycKqLQ5KWLqiIU1xBwg/GakUnxkUERjP3nmRIL6QvOuKu2byFiM51GmNmUH0q5KV
4Bj+UxiZaj0TRhw7qWdqAS6yph+oME9BnYakhluYnKtzqojBp0dKUjIt10rrj+Yd
prGWqlIw4lyfmlpcwVR+P3bpzus/4+S6S+OKF3b89fr7wCOBMO6RylQggtn8KZ82
QIRCclhHri7nmVugafa4jH3v10cQrBJTp/3nxnNqS7Ac2lLBi3FbtX1PTOiwmtJi
29ukNmGeTnfRQ5hl7fEMQGELh5VANqv3kz9zcrMYI0mcX1x147E7LOWjk3mL3EHt
J4hxvlkOOpME7DTXjpAOgLV4F+lCDcBJzGr+cZ5LcYB9uDTaO0UCiDraC/t8S0RV
LFaRSDBJnOVBUCDBIrwOlmGfukD6tH/yuzHAA9QnVsZU4ZP5x5NLGT0E3761s+Y4
yl+Fu7yQMrd/8O6NES+K8sooe8FgeTwzVzTCevibYHhI7/W/ymEg6oNGzGTYJCQA
xp3O7dXbfmmdJLeOlvjqe+GF+sIwCWEBVIW+wD2T5ueEfXDrxQMeX9OLN6Z1rZPc
oID6cVetqBeAT097j4p3ltPOFyvo2fNIA2zHxtNIbsnxP4DUGcWkJHy40nWi3C9r
Vuk10RvxPsaYZ6Y17SkkzMtQRGxh51fYWhy4jcvS5C2DaSEd9Bt834sGdWBK3tgS
78vrECVkGsugsY5WeYrLkp5wNQJUcqZzV3sN/9sHCoS2qA9i+EbfTHLx5zldD/43
S6atnrQDhuBEdGi1SsHcnSJDxX0F6u31bsSXgKKg+eCeZTTHiNYm01ou+ys/jXb9
nzZQMSF7VKdpfkIMsAZWXLY6YQB0zc8NNgJyhhi07laXkfrGJPRzZZ4p/T4ol5O+
Y1u/5EHXZLX/udh5rLJtmd2gUCjxqXnfVI6K77vY8GdGlM4Xfkx+pQoAN74tEEyN
Hf2g7gcxjpg6aO2K9MId7+Yk2zOloS3Mp+Tg7KUZYN57MmBDJMn6Mk9sqJkfx+/A
cbSf/Fa3Qy6ktRAPaTHQedydZ8+iZmI2coQ1Quu4DTUHlQIEORG2zcp3pRsipwKw
Qnf4GzM+n2VsNESDzHeubsK6LRuByJD87pu/VhF/QkIyxQ9WjJyI6H2YbZLIUCp5
AeHa+sicJiqLMBHi6BWwQllxZS0xkLvXEswrqa3vZ4BMpb1vdYvBkvB3Xfc19FL1
gfew25ZIhDmCSH0W17jt6TQ85Dw40Wy99oJZLcv5W2W1ui/wro4Q3ukIRb91boV7
P+Rg7vw3MCunL0Y1DnlLZo0UqQ1hO0aax/6TSs7eFy8S/yCs38mjQTZbsifgfZuH
SxI3LiNBwjvPGfX0u8PWGhEeWIj3B6+q/ZAMyADOZaF+MDZIBjyQB3Ih0w5FXSJU
PGh50JDY5uW15qlohoka57U585vcR3JUYrCAZwbKGZ9ZXcBj4VWnSb0kJ7p1SCQg
Py8lqI6SW3btRAr10b/x1dDxY/3xoW4Lk5sOeA578VlAmnIGFAhpS7BGdpSLEzet
kHgVpo5dBYUabxOSHxit3vnMs1kHM4HPGlrUw4ATgD6Pe3fRcpEJRtOt5W7p5d/D
PWiMDJrDymzIXe5ZUXkUOFPhXEyfiiSjI6t8ToNTfADs+F1wyYvwg/zJSlx+4yyo
/r5GxDwy9hQ/8IRJCZEah2y7rIB1Z6147ig4HBX1hhlBfmmH24nN3XhZZQRaqA7S
iTb67bmxVaRxonG+aY/938koVF4HMXIamp9BXCzOIjPfh3zrLKCjg2AoB653I3be
qXTMlFa819g0XneJYPP2U2HZWbFb3N5sTL/5YmnYrP//Gkzk+TD2PYyLtX68HH+U
gvtVW0tJ9hKpUT/GL+9OVe07XQsJY+jd/hWtMAe2QaRekaxWaVl/Hlw7Mwr8HoCR
icuaVw6HIt/GyZDVCm6o0eWZf0vIjs349rG4S+rX3jIB22zMEsheIfx6ShQAlzm9
nBC2s6RDCBVU6OlBgeVdpWBNNj6XwEvA/+mbjAwJkuiH+P8z1ccLK6pYA4zbB8DY
xnhctB0pSeyNXFBZC1ogxTB0H91fouLVU69lAZRct6n69w0S5Zklj1dKRnGYZeJE
2mG/WqbFrmzAATkAH5shgDNMCLXDo1mYdM+QGwzLxSejtIB1xRyw9B/oqUu4bxCC
hy+7s4gpu+RXUvLnntC/+dkdylLlAJQcAj8XbppPtRwQ7SsoqcG9yqVVOBvcKCJ/
nn5xF+QmKF062ISlTofpkyyf+lmDVxrjo+xBXkhsscfIb1BaV1GT1NPOdW8EWnbq
3JyjuQfWYkx7fK4QHFLCA968s8h2hBJ59iqWYc7SQNsO+/pQldVHTxuy3ulTbOjZ
Z4M7dDLCMxCz7Y4zjcGaSkptgb3f8diIhnlJBeDGRcFHXURHIGaiDkGjC+YaR6jD
a9zO3lwS8IAk5orUxtaRoX6edVDG7zAOhRVEem82SNLzJDXIzkyLuUbSPoLGj/1U
6BGeOSzktF04Elal9AMqMTR+77L+FbIsGe7DeQJ6uWG2ZKdqGkn+V350h2n4yy+Z
ySb5ByPo/DMar4fmYU+Ok+y5HTO6tAnzhfzc8x3nJ1As158cypGXZmTj4SkRyD0c
Zc6tzktAWMraUiVZ21VPP6SkHnx+2S6ra3YToKyt/3D/PNQc0DzRU7jfaB6kz8rl
bEY2hcLmyQFOUbEh2kZ76Ze+1/5Fx+QIUwGHSX4RbZy2v7eYo25rD9aHEGCKbjnc
XMhTPig/Pr+vtjQ97m908jOPOsptkxGcq6GuoGT92G4eEWk9LzoqQJUauwAtG+SS
ruyWeJWKPUMuMJyFTgxH2O2ALWHsKulxocSX2GVBEJyJ6Y5qpIeyQBCoMlO/Bc+S
SNU76XZ7XsbOwIidCzs+fZ3a1kJ/nkt7WQbWXQx3EMlLo3qnlq3CZs7NLPiiPBcx
ckQErmVfqJ2szR+9JWkICkLvKL5TZc27LXBQag4Pu4i2tdKdXItJKWcImb2btHi+
8OCnD4pCO3rX91t+hlCg06g4Gz2pAaAXHHuMj5fMeWB4Dc9m54QI/j24lMXwnxKK
PCqyfZqwJMgNl2bXQyD75MYgF9k5w7BC05kcblbBdB56mOG/K2y83/G2+yv//J61
ud0opEjIs8DkSVVzs6aQMdZI93qWxWIW/hiZGcQKihakA/jfudiw3G/v62XaNyql
ztTXGcnKUCFnHQWkIhyuhvjjiTB01ywuHakreivX+3lpOJxOoFbhlrjYc/mEkXmV
Pk1i6qUCERafGmkH3qEDLUt6DJappAqehgp1Gu0Ylyqx21X/Dtxnoxbon8Zu1BTg
7qGlfgKGx3LkFyGU7f8NIqj6E9Bn8HL70Gq28N/Ho/diEVMKvXrVged333GD2QFK
aqWTjjIGTHklK/afjGXrROqPyN0vF4Ut5paJB/QztGKJCfnlY8abpUSiYSL2CI/W
OKdizVodWyd95uPW1PjlLF9EFvjTPK+/uBXPn5mJmwVkL0Kzegfg1ievlW/LDq3w
5Vl3wnK7crexK9LV5HngFqvZuOXj4Ez7fwLVevSbM8RDGFRJBwPdGB41JR2Sr+U1
RcJiUeQ62OmXclDVokmwg+sXvNeyM9YKPD/PR2XXzQeMEOEwmqudncaCh1OOJFFH
T7jDRQTU6AeFkL/WRt4mejg5Iq2NSMx3QAnmYswZAjQjSgohzKC8XT38HhqVdQAY
Bji67dgyyEvdjnC5mnLzWJsnRQ/by/uSUvP45Z8FJMcml/uchyB9upf6WDTGcI2N
6Enw+OIMHBzklcHeWPuKeUNLw8wUiXL2/KnfBi1h7A1uLr5FrwufpLOHWimx+WZq
VAcHXuFZX/snqRnS/P42fPADuqdYTKc1T3AvHxtOAyiHs+jF4THMfbkZU2WiWOTj
xxmE9sbWR44A4bS/HgFejRWg0WLxX4tSh9vBSK4n/mSeJMryFACn8sa9yXyh2tQu
QMgRIWbZgd/ZxgV7QPOdejWjwIf0CBz7cRguWYgB5zMBUbTt+7X9nL4fj7bJA4m7
vNbFMR6CVs/TbSWTV/UGZUK892gsZJr+Bib5X6vrEb1WpOdmvZVNVqtyJawQ68Wn
DzqfklEoacGBSRJEEtVbaloFtid+oZYAtIbh023wC/iXmsyBqcyC+9Ml3EJYBNOl
GvrQZ3T8ION3epxV3KxF9S5WIabF5lCTMbJ2QnFMh5r/0AdaBnqQZd1rsxpDK+Y8
6UlLQvcwlW9VB8NLAhoWqPBQcAWEzj9y0C5PK68aKECi48r/4GjQMyEHuS5NZ51S
fQlsOVlcekfn74wQrQM55VD31EUyW+N2e1SmbgtktIrmU5/FQA8sljzlmh0Kucxe
bHphptJ/ZWob5aulzqnx2XI1JdwWFczSDIkhLpTtGKxiT72+MntC2Hjtf44aUuPp
/TxwULth/J/+NAs+ozCKC3V5WaKvaR1XE29BZZIhYexO0RNYafn9lDqR2TJycC8Q
xuL4mZod1iWdGChetKFM8sFKL0Lz3IXlGReBYZK4N/CwWfg8RhlwkwFgnYTLNOer
DlKn6mJTfnmQsyfn8m2CSuNUKNj6NuG+H9ZN7soNT2WstfFpAAcZsTStZxFGpUln
Rgfi96wYjTRDc1f2ps17Jce7ZXiD5PdLPH7fOoVDEaeynZg8+7i5oVS0KypZY1Pk
mAmm69a+bl1oOi7VXqRNHF+99kGxpNw7BB/ISLaChcMUd0Z+I6zjFHTfPrelAhWD
pR61iNxDUhkU277yk7BFGneowZfbRbfz8k2cqoTWOBkA3/UGG/IwfRVSNX2lr8KS
/u8vb5+vWLFxUMIXvYq3Bv5f/HHq0dZL3TubrHoUNhN/F0Djo4LvAJ+WWctaLtTH
dmxssB7bJitRhbKkUYbV3j8G/50L0wSQ7Xgntrb7jCu++hzQ+SepUAGwDTvkj6xR
27bB/Fn97aaWOa5GphzuUVDTTadkhT8igPHR9Q2m7BZrxDz8lx7ABDtqOw+ff2Wt
3lVQVASf4EpNRBNVI0S/OyGYJ/3L/MDsdY9lsndmcw71rIH1qYh0n8dt+r1cI5/s
7Rq9GmteKSsJ3jAjEMnadgjWue35n3+7uFxAuJnjdCQpDIazbQpl8J1Qh9kZR005
CmOfSs7vbrz+WtSjnZt8cgYlqGFx61wLVQzM+cqdYncA9QTllmRszDV/p4dh/zIF
w5yYYv+twQTPPOwTlCW1+wXOvSJ5TmGiDnxQqTLhPdY0lS0LCsUkIfAeqcLce3qN
X/4YCjqjYaOYO54aJD1KGBB+VSwKZ+nU4JhPQGPWSicu72+0xxU6/caWo9pBlkYY
E5YTH5Vtr+bzmdglPzSQ+U7y1Hea3MYIAdzMDWnZanqxNotmcgZhtP1KzluFJEHp
2otfT9Iz8uhuHWgVdo5QRY2w8urv02nlOmUpi6ZYpg0zZAOFo+WDKifM/traMqWV
9/FBs4f2pBzfZ5V0OnDSNL7yMafl2EGAWdx3RJt/5VWie3mCjLm5SaIFF/SvzE81
BozbnC2KJrvG4mL0H7FOAYYTFvQ2XiXCTTbMoi393YBJXhgOrEA4/0CyoOs27/IY
l7mCyeocQmomkqcZluB1qtkUIxovt/1j3tkRfdoYeFgoMkzo4AAzpejxXsMnSnYB
7wL3avU25lt+lL1e8olmuaW7p3ILGN4EL4iTaaQlsJ/lsP4R74gRWBImn2jm8mkZ
HFbJK0D/vhL39KJFdV7oPkZ49BsEWTt1AzVkpViflLvs5VbwBt0ZmF78q2Qd7y+K
RZmrePmsxO+fhQ+WsYQm+hxzehhiz1BiaL0Vh56IzGx372Yf6HQcxeq7dFUQFE9X
kWVF0kIFKr8mfQb7wGknUtWbMUgNi5DtEScdCWZIy2ZZrdSSsPsC6MDD49yw5nsS
5sNPwRZdhPCFDO2rNVW0QNTz5dH3As7QQ59vVZ88vunJSoYOOVtxPfGUBjo6E26t
WCp4eu4o0jLRVUKaylhv4yZ+4/9EHsh+U1aV9Nusric9ODNjXmii/VS9nVa2dZKf
GermzgSo0v0DKQeXacdkqhuJuFtCnYlNmtLqAYj1XTZhnfHPWCktoIZ0mMsj38Un
kgaS/ne95gXNJpPb0HYCDK7SMyJJK80WvQuydTgd7HokXy/dey8rj4+jEeKou2TX
sSiZJmPhrdHw6+anxh7L6bOy6ynFve/aP3wCKGBTQYJT4yRDAP51MonXVQuJP67s
Jmtx0DE3B3ploDVauKLYWeHZD8+y3WUBcahcBnVjKYXkga2wKnPAaT5LpVVR8Td6
5cp4OE8MKQy8HWu5AKgfbD8SUQ//raJs+o/+9RVJvaMa8susbYKY3yLyIy2N452C
qt9dundVEofDVoQOcyRS92OqoGvAH3cO+yelLuuR39F6ky+CYqW6Nwrzg+D+CYMU
MJ8+QN2t1AXvSRyqJGpzl+SW/+8nB+cQA7tgzUGkug/Clc/8HJiPOLtl7fk5oGcj
yPBFLlri7KTaBz6xBOBOpsvb6yFV1z8MAJCZ/CUAqG7Ps4OrtaBQa6LPnGlGZNd1
U/kkz4rVROujvYs16axmZuOaAVmyKeQ4UVN6A+8nWVE+hFS95jAkWCAFtuf3d3QP
OXpRnevDlcdSRsVRGfsoUCY1ePxwRK4F6FzpI8FAs2yMELEAhfK3aR7GudlOh8/F
gLGJ3zc62txcSsMFGOYgKiTKyNWynNeMIRuI9ecufDH+y3m/Z+dtadwcoBhjAyXx
CJ+MmTrOL8KIqHRQARmQuLHAw9aVa/SoTfju27OxITpRX4uMqmvrssTCkycgjjK6
lPswyDNg7mfsS3wvCnwmdNP0LXZFZ7dUfe+jiq1QavL7WNzMr68PWTXzLLQo2qbZ
Ojmfxc8R7BS3l9yuAHXG0yxn+JZBU34uAepEeFtOLUlyTN0Fupe2wEHVpA1BjE4K
yFjzy0TdQdijgp9Hh9N3RlZ4YFKOH/O3eu52FSnkjdFXrZ6n4URa+91b+yhIEo+9
OJXPuOrU8HClGBPbz0ieMQXpCNd6rkN6+iXz0oGQo/rrSzRzPss1puukEQ2xvQpp
TMW2ExRlgR1BJrH0wsxER9626sTRuHSkQSKchG3sR/oVja36JERqgAhIXZgykISv
XxpyadbmwGtzC+Wjm726KJ0yolWj3qlsq+Kc5Qkov0vkaUv4S5Hxpra89knvU8nX
WbHnCVQaMtXAhYXOTy+4E1Vs6uT4HVS3v/7JpjT27mftVi5nf6EGXmwGk/gdzKUX
IcYIuOd+kHSWf1D8ySm+8+Nnzulf8BVIuNd2UlhKyLzQv/ddqpvEemFAfNMzTn37
YWuR9qQZnH0Jet031JPVXM4Tr4O4pUTZPD3v+fzFkNTKeYf6iZ7ywm5gLKaN9wW/
0Sfuoc8fzbNHf4nip5E8/B4nk4rz7mBJkMBbt2rr43rdOdRavL+D+hap6RGuKc6x
+XveORdGIAXVOGf2DJN/8refDUB57t74MSvkOevQ4EYYeVVpr6DWFLN2HtWLLgWS
ByAse5NBjF98ZbGBJLkvq/KAnA49IO6dJBlGjmWxQJat1UY/6LyqJgvawleLmHQ8
qaqTDzpNmbtCn9o8VamI5J2524i0KuwnXJ91NomcujzCxxscExNulgsX5Sn6HeAD
y1zAQ2U/Y7/GWeRgXG8VJXtAPKL9n5+Sg7GelbJaTDn4zNfBIK6TNqDM+QdP/OTe
qOP7VCyMb7ZSSdmJDu2KXHEhRKIqHRgV7O8t73BkrvhVK7CpV/7wdIklSd6OHEGH
l1k+a2fq1jYdil1fUq9wfVg0lh/qmpMRCx3GSb1cyVB0EFO4wGLL6X142sx661FG
AaVKVLd5CbBhBfZSNlzInVxto2ti2rn0Abb8rrnX3mBvTpK7NsCvRS5sWYrDYfSi
ULgZq/lacrIthdQyGtuwOfPgS1eawkcV2RdxcxX80J60Dh2wio0zwTWXLN3sOX8+
fWVLQ4rr/o4DD7H2kQGytCrg2Wt6J67YZxiHF15hu2l/78fAtpumVuZk2GzrQJqR
Hch1fWHyCDNWVScOpfuIYsZ0lsdtDaiMAJ41U2dMclWVjYnDLypkbiFEv70l1YS7
DhjVPatxxpXtnGzAVw2D6uI6Eiljcgcxlq8L0MteTaSum5V1vG3s8gR+phRttrig
imYjG8SfufLIhR7tcKYiH3mwVHxHPTC1Atn1UR9tvkk1GOxgqAQRFQabUg8Cnkg0
eosNYnA8kSPc0+vMvpNGcaUHTILfF2q5HTTqr95hgYPP+Bx1wTTYY3LbpNptfmyU
ehAUmiG4jWGKQIKgbggVxc9FyFKIm8MRHS+Dv9PJcV0aUt/07D+tl43aKCglWcli
3Lk4TKD+3PwXcEKDiW9qCAbjbHfIV/WDUa/VacIjqIrrSZyXUzdtcy0kLZ9TxwDl
pfYbjdmpMZM39D9v27cvVJABICrVn/lhAK4f34mojfHnnRIEYveK946Ma1P4UbuF
/Lwb4ZSA9ybsHOVpRZ5MrT5ojGU8jwTP/yAM47VSs+YppInIaYeUdHvvzcrXww1M
mNCWDW50dRPq6QAWiqC37maPQHGT4wX5K14189KZTxSE3SRC15MD7H5Jbg6yw5JD
ZRK+k9pMt9nOnc93U8p78/nmJkUjzpwfm5AonaTC0N32aEk49VjIYU9tjwXnXbv3
JT4x3zdFLc/KpLL28zJTFFYxyqoyMk1xU0GuAqVpjiG6y9mLf1GVvvwm/4E6rQv/
VBsO7mIKopmaOleYYzn7w1orTQElo/pUkXP0eFidcOJQ0ap7ePPqv8TlFS63ek3q
tr7GNEV7iawbA3wYtgH3DCRS4H1EcS+JmZupKVEMomSQB1R7s2hutmfWPpPXedwV
zC9B0aHbKbboyyp+sxoDnikOJzgWRSgI6J1imvHJQg5vzPeX/c3IULNzaTWIO+gX
/GDh/EV0iLMTNODlS83ccYX87PNaW96MJbdJ5TOv3xS79uihTPBnym8AW/tYhm2a
O0G1/iiDj0PWowxbGNNzkhmZmf0Ujnu+06WklCxLbHr5QSt5d/oEJKvGASIn9TTX
L6quIw09X239RGylgeTWY9BZBwCwcCJsGkC0dblz/Yt0b6sciSdto5MToOpQcX91
9Ii6rbMT+9HNAXpad09VLk6s3ZdStqguqNNo7WGAAufOGR4inXXREG3wM6u7JMUM
Z6Ra/xwNjlc++Brn+tjZpFodf2aidz8T/ynXw283OgDkZStullAoXPtEnppHD+NJ
H9OXw6cjQZyjzvSh9PRFQEspb2OgxpvkQtRGZLwLYjeDCZ1LozGLQlVRLIdDU+vi
tEJfsXEAEWTswjuyBfoT2W8ytBaqmexfrNd267jOWx648LhwhgUYmGYgegUPifJi
6B5FpnoLl29R63woRBdKgappA/W7Rnu2JGQyIAb+pYqcDus0HuzN0Uut9Gz8hB1+
C0H9lTuCZhAwx0m5q+tpVI350B/jHAeakWE8A7Uvm15QAbWMgukY4g068IAx6erc
NIxs/gQf2obutu5FDaQ6lJxiqJMGm4ycjiDU9EV2YRp5Id7/WonBaOS7/MdsdN3P
BV+QUtBgYPVVzxsGFy/nFJ77FLfYc6WADoq5G1R+mLMK+QT+abkHIRLWk2hqhHdl
lrV1tRcYh89IXA8sDuiQcnkBHHwKxyUk6i60SoY4fa8xJQ25qZuI3pGU20xVXrEZ
04Sz6BDdB8VVMkCJYBE6Ma6Jcvh4AgCrf/ptz0WawhYQkl5bP3RYFHTH1AEBAPBF
8aqZE1POObmZyNcCTnKhYYfqJ+dBdR27OJV6nS8M6likR0OeS9QTVsI3xQDxp1vR
opTF6Kk2645xMn47H+Fjm2btZMIqgB4TfBGmEPV9RqDMTbhP5WKil+/V3WWThGmb
M7Gk/eHridwwd5DBbRohEfNzvDL5m25tiS5v8NS8gsvbNkIjIZUvfkeXj4I3j3ar
Ll/kiW9kWGYaKEJqlmZH9TnmbjUavHnN6LEa92bZplDaJD4Q/ikDLcFeo2jC+YHw
IvhW9EoJQI8N1ZcPKFVHkqolIZNjKb4NxU+oonN2/2zpL6S9cbcq9jiCCAI8x1ep
kuKGOaakSKCSL2xkMtCQVH8WI4gzTUURGQ3urOlreUw3xCqRjI8IFIm412rXz7he
ELffxvT/+ZieZ+ivqMdl7crkH4PxMvT95Sjzjctktu7g51V2YiufmZhSu/Guw/vy
5NYdhmIuC+b1KO/jPfF5Z/Twi2Z4DVhVpJsjy1iHbBAcoXo0SRYPDhoGUTNdMdtR
R913rK90pRLwLtJ/vyLtBk/4hItuMMxVfMyAUVrQd5p0JlYVJqabK63a6tAgGR1P
farPd83FoKDXQuenHhYR9rildrNgo8dIjJmqgkyBBkn8Pg5zYqFXuARJjQD5E6vR
u/Iq9B1ZX/ttGo2gHqGkLK9yplg2pL8QXCIsi3HdDSlGXx9K3Vs7GD3UkJP+beH6
CM7qYkaNdBCUZfe5tFr05v3O++JTcj5vgBHY3scVh7V8hTPDRJLvMUVyDFYvdk72
rTYHNiP5ZFA6kKUbD7C6eH0WuP75MbIKMQBsSCPq0+0n3YW4paO4ltEvc34g7FNC
+4cpHhpyn9zkFAuyS9fz6SHYGweDmhrQ/XcByrndwjDJnPM1YqYrjsFepueNqNfD
pGShZoUinBzli2Jn4EDRW6A9UWVUsmolfBVppR6lb0/SiuLGnzXVmeKVsOAu8OjE
YVKr7dXtIeVnQmNmxA6isJWPkoK9dWXtdeUL0rHDy8afcgDYjVcjaeqiJCg2zVlY
jKyYFSvJEhW0c152bK6GWO91cdOuYVvnP0MZN4tUywqCyjfMKRlG4MDILprQNrJr
5iIyK/7Hs2ur7nlHAwRrkv6ck8wjlQdKLX9otpEhelZBsQzXUgjvD7k9WAB9bDjV
/Z73I2beMh2CwCEQOHsQZffoyaMg9BEoZN/Rfuwpi/BX2oRmeniucizs46f8B7DF
9982VIe0Q7tjxNyyX+makYLXV6F7z+YWvH7SpRSYdIpGArh/dp15TJdZTfOLQ+jU
ipg31qSyNncsCsaTaOLOV67xMSYwQ8tH1RfjVBVDo5pLlx7GI1qg0F9mbyyYsn3r
jmPCb8KPEVFFZjSdgkG1amxgh6QNHTvx3BBmGOyc7K3HofQOApVCyaCMNDO+HQYM
a1BsALzx00PCUPvtMH42A3mgdI0RubLXz9gDr2NEsgSX5Opz0/MAau/EX/5sIDei
24LD1CPxk7RoxhSsa4pesp4eMB634o1t4ZcqxQGYF/Zi4M5SAi9c4PXQj2UPdCJo
isGM6lJDvbypKlveZm9ESb0PRZTEaOwFWbB6NvDbAsquuc81qe6L3jXwHP8VSD9c
6yFLDmlRF2PoI8S7Sli0yL1iWyept85iJabu+sbnoguFTZ++2JnAC/kJWw3ISww1
S31ggZm9b0WKZ6MV/anawI6tfztowdi7MwkhZ8LJ87I6Srk48z3COuq9aeQruOkV
MC92FTjov2ryp0S39rpKIu/DUjBZER/hZ3cBaO4aXpmxSpImue6V2eipALAxuUsC
BGhHBwZ4082s6ag06iwUdT2/CqgYUXkKFzfcTZTvACI8uQhXUKItVmXwj+Ti8qqU
R3tetuBeJ3JlcsKbonp5arskuj7i1C+gajD2p7kJAvIBhcKDGzapfGX6sBdtotqV
UXISsbMaDKmvC8KFbo2eBSse2Gs/3b5apGdOJObLCcqs27pGKo4MFt3uYHGyxDw3
L/G1ItqHLJKJAV+xbMeDXvG8PlyarbQCS6uDwQgVa6NiuZoVn7PRycnTiOfGRqO3
glweyB4k2eJ7o8odeSq1VUegal+9b9hvLGP4kil068ijvturLy3GqgevBeAGKs7n
ChNK/b6DfqIu7uWLSIBjVUiqdh+BLy1J8EHTzwbGQxjtZ2A7GTP1knFwmQwfKWB2
G8Cn7gj4RT4MrvYH4yfKP2CD5oxUfU4WC3npCGFOGyYLgOriFlVwhCMupFYZMfpC
I1e8u/lLI4PxVOb3sdPLGQguw1lv7sYgZaHWcTSgWydlX0Hipz31pOUy0+tulIoz
ryDs/5189Cq2VLXQml3lCxtb2sUU9OEBsrLqZl9cdTozinyhSSaf5fHuVgFMEenj
oFY7mu4Hsxir2Oi2XoTkog50i5W3u+r7vBmyNKYepIppnI3Qu306LkCcbB9GsOs4
4SEtg/UKTsVqp4SRULOesjv2ACO2rCTnfsK/4hBYsUSAJcfmkX3pcpH9tLk5ysdJ
LvzWG3OS1SCohkXkicL6dpi568aidPApbZ5FMvbeuJIzUNp9AgPUkQD+O9N2B2oS
QzjdO9fWM44jXR5wfm3fIWvQDsrAKui2xnklJ3lKcn/yQA9VxejmfXxAs2VaBGRN
0rG7sTiiqx7KQ5wWinHmG7GHgtQnSOYN5TAcwrjFEnSfwES7nsk5DsuXIrv7xnMr
xASP8XrB7Gak9Gm2T08IhuwuRYYhqZceYYYJgMs2XTeW4I+ldWCHUzXHn04Y3Z9P
QuVtp/DHaqV7cBHaQ3/aqig/DL+EKdHZoc3ucromTfcx4fjgVhmvkAraXiUMGNIK
Ul++Inyw1F9Ay2DLp1LyK8vin9T8jwb/C9cfWGohQXybxHdQyvUYSc5mD05Kg/4X
URk+qfLyqTsbJo5rmkpKprJCp9j5WnS56a281dD/z5k6yRwMfr3a3jTIwEsxX7Zl
A1qNVZrI6+KWH27R+0cOM83kW4d95A1h4JXBpFdh8JqI4HLB8oU9yeTJOE12oa2Z
RyR5QG+hfCGUCgFkDEYMA1tDa4/9/2+TY91Sq3PDaFJtYUbk1aNVzwaH5qXq0VdV
d7DEFA5LNI3OsidJAnihN60Ky9A6kJzJ/2fWrzSTvW//5R8j+Ubj/Tz7nS+9WmcK
1PnvaEiLKoSGRLng6D8Oy18VOlaaZg8NEDQQdYMLHHDD2dUicfH8uwH9AmGODbeP
UwDF0u4aD4Lp/7lrCbYTLQhWUC0Ja2L+JLC2T39E546QSAUVHGKeK7VxPLHiw8yx
udHYiPMaLMvSMSgaTLUmyVYSdi5+TPCKbF+gsNy7ahnODeb9LaEr4vhZyrTHkEP1
zMV4dl9wunTJNCQ3pQg8Udn6qnripNRXJcTz6vKQc7K2ADQi96xEaFda/Qb+bmJr
KupZ9pAiJ0y/R9nhwWx8DZbkY3d21yOcQbqdDc6cqyxUuvdPsU81jhylLCgN1wtq
77gXXbNPSHrooAp4pN33lULNDlrJlXYpyFD+46efIfBjAHiG2r+AbRMk7sHlW0yc
2bigOmltTmtniaDLO2y+51hpkShySXrCF2KjNcBqWQ0xJFwvUS9gGqd0mEggBe2k
scnv8HBPAxe/FGln3aYifMJGrfFDaBcNbACImGYMDXxMf85GhiIPG1IHTPBTipE3
VM7PoQFjH+P13/ofMzSEMQphSgmb/LmyCic8xXU7BHeIdepboP4128yfX/EGD6iQ
NaiZhTB96kVGSvwsExJXF/eO+Sen48gkduLoIYgzI0173j0Rc+XSHz6u4XSHSOSW
U/CjgaRUPvxvuCe1cLoLjTsQUsWWFL/tL6QCHFbr2q5+26rOeroMeBY3UIIyX6KB
hXFd3iK66a3FYYrli1mJN3ozY5c1U1AG5BoEvJTfR3kLJFFO8J854Y9YltbQfNZ3
fSSQqwlGTCNfVLTH0I5unpydV+SOvXMjpbWz5j1siRgg3f6A3bCOvrqPOf5JCMxI
3Hn8u8IPfCTbxD1zsxM8d6sawUyn/d6NE4YTXpwb67j6mi1kKhoPtgzDpQNfRWTA
1S7H5ACDojrHTXDGAMg8bmTGpoO7wJM2GT+rA2vAibLSfmIeF7d38+A+56F4FZIN
ZUB7CXPrBOVVeiwfnW4h1Xz2iL3XC7+lpfWqETocau3Xkb/pQkKRDa99CFVJjgdS
fGy+Y7/WJJ6UM/pvywGUESpbtXhdA/Mnw1z9Clf4bc5cnvbUmFWfCUbzf+RcHL54
jhjvB9LEZGoNUbKzLjofRbmSk0hqkbYFJjlEBT8Foyurag5KBa/Fm36e/s/v5R8v
TxazYjGmGMpVBj/P3IGen+SQaApJbyu74C07EhhrjoDaA9NJc4F2u5DUmoj12wBH
QRGMevClO9+mL+lb2Xu0IOlSj7iHlE0N/tdIR+120BiZ3LJtvuG14qg6HdZyPsFA
QY2X/kE8RH80Y+Jtfeh7udHvDuoEBTBlIetM79FGbaGdnd9dwtnPFhihTBjkiwhq
WtpMmXyydTD6OD3qgxqIo7BvhfazKaU1StgWmiWN3lYIhTLOhRnmvj8YVHM2lQtw
cqViXFIXKAIehOz5GqMowrMY0HZKzBW/cMdZBoQq82KNLxIfSB4NCrh5UiaXl2gs
/VVzQ0aeQD0TrsBsnJkksFFfbWR7kACLYSC4Iee3wK3qiY3+NxQrmecNGneTfIYh
kcURY3ruiYiIEY/2mb2Sb17ZotYJnse5iE1txxJjvq/F5oLJlbeC58VvkYdTQLev
dvjKuhHcn9tc575idrNCoQjE5JgTn/qyZ8vu6urJQvo3VrkyoW2xCZMF/19qTaUF
Gkz1glYVFCPHnFANshvN96qR2nySrViQdlloCWR4DjsAx5/XyhB8E3Z+Kt6UrL6Q
JnhK0tKCbM/VTaHHVcLvQ7OHr967dK0rLQ6h4W7wpmm/zWka3yAAPfEBzS4mBnpL
nuKnQjnuCK5li7XCP2eLiCqZoFALDepqCuT/SOwD2q6BVIIko+kTyztgPOTpbKi2
3nGJo1NgIxBmbxe/U5V3bqd6ZC7v/SZ5M/Cv90WCoQHNB3g9xynHk+xfkIcQqL9n
PaDVGY7YUtVreYSsZXMQ76c93vkgaLn2YhIQhNNvoSe7QZH3bdPc+jMjt1rI9xsf
BQN/SESOidpTd75tnwDWhCsJQ9LBpl57Gv5fNp9lbgM8geBVHvqMZh74ShD8c1Yb
VTvpBNSOAg7WUcaSdJUcivn08kNoqpy6iU73D69QB2mKdbs+5Vc4pCiUnkgTQkrU
2AoWmUTdsmp7iH2Oxsy641CCMLejPVrVi8Xg4iJixbGM9RIKM5m7rUdTYE+wQUIF
0fJTwdoN7eBBcQKziEyoICOek3zqE7iMyzcnnwNgeuG21JXQ+VU0ffGsmy+CqqNj
s/1HoZCvSNY+uRZwwjclNYbKITmNQSNy8YUUQj7HrpSeSW/9TNuRZ4rCT0ntAfCj
O5X0TdLw9OLy9c8E5eR4mD4dr1ZwUV9xLtaxVT4sfIKDKvLYGkpMkwDBkZGT0+jn
OIumKb9pSIDJgcj1hqaOuSEENIiPiPtB4CQIH/5dGr4qKpc1D2a9Q2gPZFJgZchU
nIHzPxnVv/zHtVdl+9c2FliDIV/zeX+j8iQ9Njpp21cBKyW88SUlY5rx+t98tQM4
ZS9XXuEQvUIWtBNgbQJv0crcpLPOTbGRvHn7y9Qv3LkIlEwJMbF5Y1vDunWIsGNC
jU5r6Y3ySZAWTjtUIIEh7asBseO8pk8N1OQKtO/MzUj0lLGaElWrTDSdkYbhPA3T
6rud/u6NPbPDU9QvkxwYm2FVRklEQha9CLiz9mbOcki3B8GuuQVjQgKefQfh3pd+
rHsOlAgZ4H+jSiVQH8O/AwpSWUMlj9Fx/tR+Br7T6YymfzFgkgF8Y4SHYJM9H07k
sBoOpFjqlDjVhroUmRazXmcV8MlovA5GgZpq85THNR09oTqynj/5geCUWtI+zdsb
d6FsRClQ/xP926sIye4xmvU+6nlnSwLSVhVUIy4brubAyTMyhvNYZ3LaslQ6FhNM
kRx+bgK8CbHnYs966VK1WWgMM/ZJQlGZxCuQTPbtQaFhVZJBNLH8pzYm2brARXg1
DiZQB3V02D4Kvwd6ASwbC6aqaHCmb6SeAX012F3c5iKBY57ehWM8+l/Cd9gyrY3i
OxamlbyETCBsVZBXZxfUDyvJl046U6XBgRs7VVOHKRMUBVle+kj/OBQAuT1BAN1u
jAW9Dk/RIdVudB99h+D9ok7fHdbgIUfX6H14BoWMA+P/jfXu24AyGZ0IO40lfRlO
I7CaKMtgJBiDhCkS0fuVums3LuXz8nN5DQPHP4f6WdWGuWRpbuqKoPqFPMeYkUID
Uv9M758pBtz+i3wQNo0YrMTnel1Z7p0Xb6+8xZ5AKOhl/9qcLQ+eyfoxVJ3HqEQX
jeRStRcnmrXDvpXFzxeLaBaVWwzuGt6BtioKuzbiT/qTzCK0M+lWbGuc3jgl2zHt
EbCDh2Xo5vLmoR8ghF+2S/ypf/jItT9iKEr06cVnRNhp+l75L1NPGBj2vH3F1FN3
tXu8gw/t9peujTwwX2rUuZYAvsOwRLnlWapB3VSUazPR8YcnyNeb4cwUPbwu8nkw
4j1DuyHDplcCDyl9iWe4xetiTFLHBNq06Aolx2LBOz+jJzx1HbPCKcxkXEDu4Q6M
5A7TnfiIO+a2GN/cEV9ERb2TJMHkyWSgtnk+FzYib9eHRRq+TW101AxDL6e6coTT
6B1seBNi8gQUK42o1iqDViprhaBtNR1wLGpschbnQxfTX4Vt8/kKwVAunXsDYmlV
EMpLG5BNorCOgqMvTeXS9nWCOeVq/Hnm/7s8SPyUAZdoRJQNb6FguFS9P7rVrdLA
1/ugB9sKsGOk0LzlxYbDp3uVdWGsqg5sGPozT8Hj/79JPDophXDW+Elon2qSD2LL
CWer4PJ1/teh/eNFFrK4RYpFiFgNNmSLfogTDJvih3AW77GmZztCsjULbPYjn44n
+9UO/nZUH4Ix5tlnigyDiDEV+ZjPCa+1O5NDTcuOPNI6+FbwkdmLzP5oSEfWGB4V
I2yky2h/VPQfiosQCvfpNYDYOlqYcZavWaRBZvV48UqVpm2HPX8S6VHC8JeyfrNB
Y3rLtud6ezc69OcppuECF2sCIc5km1uBgO3QvhjQco1jqhungPixu/cE9vHxCDlM
EEL+QW8V1sS/S8Vbquoc7BITLqZNIN3YS9sj8PaH11Url8nTsK/S5iH3ffHSRAGx
GLCVLV8zOWgVpXU2fHDiR71cL6iYiMdrAai7SllhW/rU7mLHK6VOtmO/URmJWC7W
p7WpKQvMBpch097qNlv9hEkXWC2Q6dU+hmI63VXaCEbcfMdYFAZ5B1yWlH1rFwW6
EsQtq9UYISZ/kxdbejm7i4IuBqVYrJNkQ42Kdq+GYG2oY0InOPGjX57ZcajqJ8Nj
6TIJKacSNHTYVx4TXZG3bqMj9V7zYnFOYP0aQjVhMqx9wu6wVVW83QyRcbZRWgj9
TRdw5oQ5OG7642ANSltKLAM5Ippf1A+6GpKQ0ui6qktNOwbHC8pZ1yN3j2SiIeUJ
F0WwiRoP8eh8e2OFc5RjMY2wPf6BgATp18MJwrUXsS8qlVMtxvoHM0mn6ki/lQd2
lZdKHFGRwxewZi41DM5ReA7xCXz3aQaSxjJ2XYp7LxTNCIg66+/h4Q0Bu4Tn0igN
Jy7QiEOBdAfuri3JLtkQaVAU7JDbHoJlKr0tOuERFYUtKb47aWff8ZwLFrKvjirB
XOmVMorfxHN1pshgS8qFubEHgALIevvljpdCGqwCHQ9Nqq3XFCqeezkDsjc35qLd
pEITDyetVCg9LyFQTGszqEONDX0bY5Rr2hdIMGPLo+Rby5IVucxd7pGh+cLi71p+
r/faP4F2QQh2ReWNiJAqdjcy/RlTy1uZ0g2+zjF1kKLcZOBhfdRuPAwDMYlvG7EN
MO9TKxMRCibY95jfvhehGy1ddDZTqZp6ZB8w0lqhknEerSqAVOl2dpq78NsFsnoy
iLm4GF3+gCzGMhZpTEw+AUtDK7stzle+weVRHCdy2AEatNrBd+etIoNHOCGDOgh8
wGTe4k0+16VK0BaqsGezUcmuXDKw40C1fEMM169ca8A8OCTSFW3FqOSRMQbgGbOd
qSPh8zaB6jAogQw6ijZnzc2IuNHJfJEAwf5UJy8iCFxlSeXCdmAsD5s/PI0YFYf7
PjszJnoWSM3zbI+Rp5avMKQPouJAR3ON/nbBZpH3SzCXszngiCRI5U2JYyZFYTVY
TpC5w2UAH0AFDsoTxcTwsr5RXnx14vDIvLSnM7S2lcShc4zdlUsnPBeISn//KORY
MnNhgp1d7HZoCC9GmWhyJoDgGQX/QrxSm+9Uwg1o2YgJS4o/9MQKTSBqHcXdjsFE
3O8yShZeBCF2RynG7Zog8GloFPJFpuZ84+xcjuaDYtojE03MVMk0eA35QVTTL/G7
mOfSy3i0Uay4pFGs3y8mnegSvhik5PBd956wq54tkTwcoEcSZRogfAYFFWynBXZT
OeirTOpVvceooepji7lCXsawo3yCUJ0dfjdT3TZezYKhXmvJ7jQUyyI9wrnaJ//F
dpp5WlAUQeV7fZvf0eY25E6nEVf6OnKgE6ZholDG1uZpnbh15BIuZ+xJqvoGx8OH
3yJYQ8OhQzt8yvc0kXFEvB65UQdiDm8sVz46vSh7P290f7ygy0r8UB74g8XvMp7q
3493D2dXIDY2TcZSnhwkA8pCuzuadVZafPM9y7+jT1CLFL/xWeyC827Sr6X2fz9q
3QC7Tl/NEx9fZss3MfRvXioXhbfSJmoLj36Nc7R256w/BsSsVXuN6z5e1UtON4BV
ZsA0Hdp/SD1vCKVfcCGNY3Nx2AjtgRGnuOx7vbNUi3wISoy4aMOm5O0CycPWTlf0
7E6gOhUxtc65hc9L1fmXQTAoIZvWeHxjTGkgevS8SeczWDD6BgbQnl6WZhkHfkq+
2UbPOI2pI6RyWbY4JtmgVpXXp7XZ8EiCV8PVzC80gjXa1FhRRnJeAURXhU3howYE
ylRwnFxSqAoi8ImgfFuz6MkGiwzGoNtqI+0EqjiuadP/EEVpzDZRC995yjj3G0wR
8J+3RSkPHyM2HSHTX1/RPt5IUloW4iMUvITAd80hXLDFOkrYRFs+HEWH0kin4Gzp
shJWxeH/M3NyW9EJMv1dFF2yAZth8ffAQVqTSSuWfY8M7fmNBzHSeGGiBii4eX8x
Jio6oqtPwzoHDT2NeXChe9HzV6oUSeLhs+DudpgWJwoBJp+EYQZv/vijdV6braBI
PtY6RO/J1IN0BPFIZic0jzfbjGcR0dW6qpUWSsz6yaBanQDnoWE1Rv48lZ77wklS
63cSXcMDaHmYND99MkkAyWmpnXLQ04j4EdrsdE6/LJ3tBREulfgK/fJbW9ZWnAVF
rwC8pzuNT7x7i6SrfjUbia9MpVcozhxhLzUeZoYubgyyu0FmFu9hPgSnL/nk2bvf
Swgd6V4/Y5g/oHn7OmfGd8bhfwtK/24jNXwnv0AgLlrNbEWqv8xuLwBrenq3brJH
tM5Cc6ys7KeNnftZifYBkSlDycFbweHsBU0nTBNh38Se9q0xPTE5GPwqte/c9Ngq
d39x3p6Q32LxdIq9Mj1lm1uN2l+0CH91FNupCORBAnqIl+IMymR2qfQyqGkIha5E
BSorYUuLhXUT9a0P1x9GemBYe61c5mbFw4b007oiP+eXMKzM9MmiEAWGnlqbl4mx
EgST74Vzz3gIaw6Xr5JvJAZHe0YSpw6dIK34zAVNecz5zyFKgYP/6mnMxqCL2Nk4
88pJ2FcUR7HErzouWhUBtWUTj58arwc9YynrrL/3GPnAOKI0vYkzjQcmuxzHio3U
fayA7g7gWPdBaK68n6flgQHDXW7E88ztI5FO4qKxXzbzCEiYlEZ/zX/cLe9RFYPz
1cZPaDcKzX8WyStRhp6t3iA/usm4gRrQ2JSQ5Hwf/AzZu0b1ziKwH7nLSLHyX5OT
MnLgXsMdiyeVnENOIVhb/XgiDyZnFfDb0WlrCIJ5p7kBGVQiZLCF5BVt5wpE77fv
YyjTvoeRBRw0r9TV1tQY4sNzH1tygqjRga77M9E40Qjg8/1MvaByUITG8AZIAA4W
WTu/M5MB8LTTdriYhuoD4C3iGxuNWE3YhB68tPeTx+ih00HykIdPYnpw7lDp6OyU
TpUGfZhIIxdyCZ5WFPwjFAgqyYgC+/qsr7gQmXtZNF9ll5McNttUVjo+JWRVzkqM
tkfHOSzaSFjZdjxh8ESCJJf5P2d1EXDiMNMKY7gFqGF14j9EOQZn1bp0mF3QXIGZ
GPpxdAG4FT6wTohfOBoqPWnsYbngygvrfFkPgONbGmKBq/Dc7MSzWqn3xuoI++de
AZJ3s2eAyWo4IvKnTwcA0Ip5yfxN8nXnpLXATxZiqKKWDQOny5Ik0SHVqkA3mEbg
JwsJtjYn9We5wPDX3us6DUTzNzmkMDbjdIEF/yDSOpLbOB1cKGBeZHr/TVF5ePI4
K1Za5eYAatTT8IEViwye9qLPXBrUgL4cYzGvO27en2YNyZjW22ZrP4D9LaczEXFt
P4VfS46WI8aRJJxgeTyoIZF3SLIK7nO/j9re/rddyiAvJ72IYKuSejVMehQUirXd
ocL1aOrU/dY4xhWxR97HkKaGmeSqO7WRkcIOWBxy3d877N78U8S92WD61aQYUns1
in1cDJ7+pV6tp2hdy1d51++LzynxVXQU9TJuQgAwacKlWIdwZrW7Yy7UhdCVpQCg
zhg7ABgpEBOSn3WGqSHgfnMyJWG+48juMgzygufO3lMlK9BWe7P9oUIbFD7Wothk
RNjD6D/VMhOYzZZSGXqYhj9tezqjs1GG4726wQzBtDipr5049Fh2H1WAZ9ALP1As
fdzQfOYlxPqJzgfekai54ZAeCYQiPdCnGFBgb7ETk45lgEVCzMnG/z2cUMf26Rij
63za2g51OB6oE2hGtAF0L5nXP4gvc3Dn+5PT0zz8DzqLd6y3XvyCR8T/18ZZAy0j
CdmNMd/6N/8WK+JH+9Zp6syFbSGcx3pXFxiyXXFyUPi7G76omXTJC62mFVQpkx/p
y7zzNLvrDQq/OURXKdPzW1Imm3D0KgCtTXcjGTuqXL2ZAVT9nBeY2BkQPf8zmTgK
vFU6bNYuSSfJwVDaWErj3ANzQW/KlFjC5PUYGwe9+SGIh6sb6ufEPOFsL3Ct5BHg
jnLfTjvpBb40yX9uBKweuj/DTSy6BwyrjE510SpxSJr6apMVtWW6QxKp2ARbKYQw
BXDdIEvZgtghc8ku4Ens9Ww7/Blm8LMQi/NGKp+CbHzK16EWsTOobcF4KPYW37c0
lk9DiL+J854KEjzUW0+IY8HcmA8idIgoZOlkVsJMS7nTJ9HTv0Psz4KyAylxCZWQ
sD8CBmJVcRUM0ConEkF1TEuuP5RGpDtfg8CSFaDoNSpCqvgj1XCJcoaRVTOCZYqV
9gYWMFOnhN2V6oF09SkZyM3UNDivZ7ci+50Odlai5EwlndbXROeeTkaicxmxBLgq
trdN5KBB1EKbQuZv6BxjqzCbOJ8a+ByHDvEahJ2xsRcZjWoj1lxu2x9kQuarM+Xf
COwubsihwUnmskWaB47C1bm574Kg2vhjqNiZ97yI7LbxkjydI8049tDrN92X+BLR
1hNaXZW8GETfBRIPbHHSM9Cw2dROUhTJ8g9lecoUuYH1ehNs1P8Q4hTZJJJkpxkR
5ubOpP0/O04obb77shCpYHMV8Uc5mkh4IZQeAvPxDeK63oph/3bh4MJ3jbfDirL0
Tr4dme3HKt6g3+kCT4y+ZK0YV0uRUuI+Tfk/wrx+7N2W7wVMcckggsygMP9ip9kq
+2HqgaHQVvuJMj5EatCwJri7LM01lRvI7TilpqQhxt7vpRN+YUVFYbp8H8RsR/Iq
GIlIsHZOpha4KbbNWmaSapzKam4ImBCeyAcbzzitml9j6d4wocj1+GDJYX5sMVZ9
fnKXc7Xi0v0NSQcXe4i5wzF2hNYf9TQN3j7LIjRs80fx6d0hlC5yyerCudjmetqP
ngf2MHR4dxC6vNeVjhzZ3rAllFGggPEV1eXtfkmoJjEdPfr0CMIAu7qRRg3OB7w8
srj+DOWw7vBV0FlG0ipWjWuP2yZ70J8r8vBw2+jkZrQaS1FqajM6vxTfRDBZpCli
kFQNri4TYH/3MfdpSvA6Gg3HQr0E2AN85t9t32Qe5YNwEa+1aqQS1+Df3u/Tt07m
5W3T+D7GRRV07x0TLOpmRySZtXFx7HG8ucuXDgotMGPgvhhqCn9hSXJTDkuf4OrZ
0MZfd1/kw59ZeLAQShYSqBmfWcefldOBBr9wWh3lzU+lRMEx9KTUD0miPKaTMcwI
AGs84hVzZtxlTcsNn1i+PM/kXvHlFSWTr1Lk5EO2N+uyNlGWbgHuwCctL5DEiSTI
wdSWklBeDOV9n18yhiUgMgE19kMawTtz9D5YUpoW7eM6fVu+ts0QQMlZxMhBOzv4
P4xECvjwudjjl0koQW1voZlDcKbllVsUzui/Znx5SxbgbZ3Yo+UUDlz7GMcA3Qni
O2nWZWIF61FBSfy09+lYDmog0wS22O2Jm05Hdn4nrbOKhi8a1XQ37Nu+WmQkzoEH
MXuTcJolviT5mIrOcCyD1KHZb08MBloqkkvjqMmK8tJVRfk68PNAIqPJG/9vqyCl
LIzZgX5eOL8jQA1vuAKTFSP9B4DQ8oq4W2sPkpmuhECpW3yHx6DK0ESSOAj1QJ4+
EaIGWIsWxfTj1WSOtK9LCZ8//1f/GXVl35pNCAMYibwJA1yZ8TTiZwok/MD6AJ7X
hYAhh1xIBkok/JOnxG7v9yHw8gUjH1G8o0QwQuHQZ3rBQzrYDm5lZ17uP6YSB9TN
gj+AmgdVe83hImk/2W7sxrBCAUMnUOMZGO+U+vkTedOEU8NBNriDFmcLN7QQPJdG
R9FWABz1UFwfIcfZZvhYhJ8dzSaIZHaNnBqTsa5kvpXOWpuVlSBaQSrIFvL55W0P
3eI1wKRi3Q6XE76mD6gWoEA+EjJlSzWv0p/mUuiyfwCihigcHpZtNSNRlW6Q1f4r
VWg2ascHU3he4QpozH0OtL3YeWFWl816ykYcaQv8SSNEukuUiaVJiW54bvidR1Fz
ssR1s0a8voMoOX7UxhRnlCzAMP5apX2FTIJD2+JNZuBw4yO5mIwa7ooo7THA4Ktx
gR9T8/6JMgz56p5Aw4MJt7W3sUEnSxWYiHv9e81DSmZbrz1rFNjkGX6FbOcVnu99
OX9gJgiJXfBNXVpA9CUq0y4B+0KbONACu9WCquCw5QG9ZOQV2Z3M/k6x2L2nHLjy
LZP1NGlfbBPnsIwpHLFnXSZmUv+ajLCeUSHoeC5wUQieXIr5dzTago2mPzlhwsIJ
/7wJNzOBYmIG+72laBg21LKCf77PniBWJUEuWlcNYh6zgKbZPXaSdPKUxwBxAuM4
tGYMA93bhv0fx+qbp5cwJf50FbNfuxGclNcFI6eP6qXTWudevUAyWw6N8yjyt9DR
oeuh47n/V3SEVCS+R5kVxw/B6l5BozsoQtkH9Mr5ctyYYOMkquCzhSTHghoRrDdp
VlVm+pkz4IpN9DINiXmj7OWm5TYluz7/KPMrhhNuyv9cm/qvGGqNsLkfB+0FjrBH
Fts1jM1dSEXMkujHeu04KY1mVd7zJJa103iQIWYTZQMRQ/P9fTgYsjyNGarfmR/E
shrZ2yhvYM7L/I/XbfC95/FVM7fMDLU74PTuuDPYtSSSH/duhs9zZj5kHUp/hhNn
/zKNR4LdfOZgyVdsbvJCDE7n53bqonrt46WsPM7Z4QO8wZQIL6XO8bZBPBr0VTTy
2cUgXvYnFzLxtCRU4RVdiG0+nmzCzDjuNbsR8aSi6dV6emhRFxdFLC4IVnUvQMZE
IMxBA1ExrAKSCoEkyBkTkul+J7iauos6rhHoVhTP5GhpEDg2qf683rGp4iEkb/Rt
4tNxQ42AAdMFICd+7UL4Yoka/66EuHeAZMtn5uCPNxIbA2RXaEDCyL/HgckIJJDb
ssefrWlpB0K6ggom54MyfZfwP5lBHMTTkHK4w4nYubFzPtHjXcw9Dxy9d29fFQDF
j8VBVtI2BUzTa9BbxGeEE3z1hp9TcPEdMX5yQW2w6gkG4bPQLeGqDVa/rx1ZhyNL
UzH1vDS9RzKcx4Tt2xqudkBxbA07MOMpsMC58cenltrslB9QcvThKBUfhCvhE75C
ZuhgX8NOHs84963j22CpWlANhxd0u40I8I2j0BB9t6l05zHeYVwzfhAsuVgcxajk
iFfe8lmZwlLJtxm5CcGRU1x+MqDBoku9HrXCDJvSH+35R/f1Ykvfaxuu9ibJ+5ag
2WYDlfve3z8WaISk5CEVRHeFXAsdgmya1mgXK9o2T5gdVBUF2FVmRV6IzlLJNMkT
4qQYdddEpLZDi887MyuO1ph+vnYzhYK/O5AQMNm/Thdw3ozpmAUrZRQZuFHSWI71
7s8ysAA06mgbaZp5A4DJA7oLM27yJ/OR8YK4LT6XimTlq1Z/GGhwJiHlszHRi2xg
DSMVIHNiKCwdrI9vcdRShQOq0hzMtYulkUnDcxoTrJD3Z09PVIIQKRDFCEtPZ9Iy
ggjY2VSTIKPYAKyw26opWZ4/VaWKjnQFIAnH3aOsYc3AhGiwbpZwgBNpRZIpYfGA
RjOPShqYAFuKYRnNrRg3jnXxfeuyv5WZfPyRY8XOV4lm0HGDldN9p0F5vwe87Kw2
7SQSK9uGtT8zhoaJNHbMN58O5JjoPjYHE0nLoB5GMfiOhoPy9VOJ48kvXhMVzZZm
ORvZOU6Jy/+rFxCuCDs/yMhEluxFJ0wbjpJHDL95obX9+V7Y1lYOtNcxHjy1uhHs
fcXm6NrLtoEMowuE2epF69Q5ADC9t2Z5NCb8XRFbuCDewLM0wxU5cqsMRYIyctHJ
3Z6lzBSPgRVWH8vmT+ePy4YCKReCa/3pivJ2GcaoBYKX94Z2KX9/zx0GZjaZSqQb
0vYZ4U+vhzoCDeo3J4+AS7rtzNuCx9DygeSPCrBLXRtPJk8TZWZb/vhSpfGfPz2x
eyRW/7NnA4N7Vg2WLl+kYUSFRhXkWUenCn48VAxWgNGFSdkFyN92kuHVWEUz22tA
gwfntbfzj/MParx11oTCqPJzw0LnUQfVjDqNQPB5Ks1Ilqw6URxEGttbNktYl3dD
rZ1blEGENMZSWXFfKHWMBuvaNi4JQKzrQqIKA93N1GtxHEIbpucHrPp4IJjr+AuW
BpGRPDfIDUEQsRzbCGiaQ+XRAjpEPQBxwSa7gSxgVtSgs/hYjcbQcUyaKAU1/FY9
ngr+b//7ud6YYKz2jqG5QfKduimxo2dL3SE6CwQqgQ9Zs1Jo4osxYSJ1OW4zCQTZ
GqSVH3Sd6cWJ3lxuUs6pGBL7c1b6imtyBv/rJlPWkxMd2cF0f4p6lG8mB2Vw+q5p
WFtaTytUp3Vdrh4RkRiOD4o+7m3YvgFgn7CaVyO8Hy+tBAhqRy2JS5VGncN/VUWp
37Cofnsz7QnVZpBcydV3B8Z2r8X9fm3ZbgzS5w6rABt6d9ePaIJnAmGKBqnYIA7M
5g4UUxIClYwgdA9qgOc5KqFSZzJJQGFmvJ/4cue2fIGgvNNvStx8QrABgD9ARems
0oDBEx4N7HO3owzcWqxP3TnZYFV5uCgSTPyGQ+n4q5OtAH92azfb8yGCeGGkktoa
8C/EhiMQI5qKEo58TXjC/KiZyDSfPdHq/6IoXqzyDW+9D+KnqnxQupQtGtz3hCwQ
d4UJLrS+frSb86pb3gfLPje30LPcytxgr9KbmsK11oICUn6lJxdX4FgSbSVoem2L
kDCfj+iItMZtPhFtGh9uRmV7wClCcUkdZ/5PJqE0BWmhflCUi3q9cQwaTRWfjuA2
jvnmJKBmyVrljrip5F5SqXNyP5p+QZyAIx7ZIjH2PUBK14G9g169Kg9K+ZGQPGTS
BPJ2V/lDE0Z5p1SI1fxtZ2kFZ5tDZ43hNT/nVMnOBPRmXPv/a/RbVkfN8NmvRabz
4Im3sDerlwhA0lvyW1JXarfdBRRYClSEph7UUucO4QPTL0nM3M+2d9Fy36EF/7Ij
ugNhbpXkZafIPr361HyRL1Wb4OjYKtHC5hMxQorN3a4xMWK00V6sb9V6n8wohTmA
OGZTBuFEeZmZnRQrClv4YCgaOLCSwVUy50lMHVki9y2m+74FcO1frbSDXHb6ok+8
6QEPytVAclP73ibeioCBL/GWQpACwz0Nu+h8RjtyyMbZCazTlJghUbamXRg8xEU0
JTrYIsqzLzpUcBKgqhDyrl4rwaIJoVuSIlevfgMzTpq7Ttz6ECFIckiFoDMjRubt
FAVgIl2D1OpH4N+vZGEcUg825EM+uXrt/CnIvcLpg6cTuMr7KpwfVY4jgT8EpbVw
JrHSR/x5NU/fuWDwm/B4mmC6RFSDX0tHy2HayeVE+AiUXemn0lvdHBqgbzFTgcso
rpXpmXHgSpVFVsJTx3Fx95k2o1lvlLZvTerl+8NkdhZKj0IXDyhvWpv8dwn9I371
PtNfnNjN/MuI4313cXeUElUllD+YGCNmSgTAoT5ceZUMpssJmvhh5DmayninyxLG
oYx8RCy5FvPT1Rq0DKQtqIq9BbsS5Xhyq8FxXaxtKhWaw7a7GD977jiPOl78JNQO
nxgY15srBmloWhwv/sQ/NMqTlq/qMVE3kq726QmtmM23aDtA36hYyTZCKAwAncIx
iSDanSuIWZMqgx65/xPvbsjpR1b7MDWU2nuhYV7Dx3WwAN7XChqczTcPdXlAXtEQ
pRxJZ69VepnHQX36QX76XrSUBRktEXsU/dch8Ljt/HMxZvT/sNxquQ+8g0+AJ6z6
N5rQEYAHaqW42jcaA/2izXT3HUZQgpTEJCHGmpl1tqSuOsA82YONJ/yFjyIgxMgX
1yMnA+roSkpTJvC8UcJrkNNJzAjcy6O7y27JmVVnM7eKKfNrDQfH/JK/vOHN1PWB
kVYRv1CpvqsWXr/RnT4Gy03TM5S9BGsYEzFOoMwHduLHma5ygP9GoQJYClW/yVhI
c/R81Mty0YhBjPjfG3/YVXxudzQw4Un9TArMTvbGXMKbbBSuPVTA6Gy2w0gHfWSt
xp1jhKmZreirSVfrfNdnv9AsyBNAJdaeJRwDiu+EZY9EWZJ2zAOKP9Dgd00oojj4
8wWMKgP8efeZcJz5OqqbpRDeNjvZBze0P5ZPfwJmrpj8IgpE/SDRVV07bGPExKB6
74cYW+Sn5HknXYBQPIGkQiJuCAU32g5nWTeftP2GOex8xUv4eyiUXxCOPFaflaFV
oV8KapSStZ7sJK8EIREEj8qM+0ycaYSD0EW8awYtjmsfbJwT41LbqLDgYPK0k+g4
YuHUlle2AesLa8oxZ5fZmeejx+njVhz9s50KpMCm18ajWrLR3RZ1aaAjnL+WWGEe
g2HCzk/Z1ImFbtSKK/Tn1bhJabEcebXDIJOX2vrEKTEmAxGtWiq3yUHW2zJEo27I
aF5pICax4ZBSe5O+vYXqeUYotNPktwk3M9Aph292UuLlMrkaTHjAK5/0Xh1fUerD
Sabi8iaux7L/ouMjmzoVmKLf4J9wYzAaBwtPizl+EZM3LSpepk6PpMEa7peMrUAF
+NKPTjzQYkrICPJsZnYqwqxWZN1zX6+kpUKyk/yw7f5bGD9gZWWlWNt0SvdNaKne
FS1f5AfiA03UtiwF8JYGoMlLalU9ExEpHSj14s42orJNYBqJNUvtlrMW9eT1WB7r
1xvHf1wR9VM+CvD9vYyqrB7YGe136Pi6p4kYDyg5FOnriIoh7TFYhGFazc3nAT/U
9CnV/EcVw28FCmAUCEz+ikR1HyeCwJIxs2ggdXN+CZ+xbFR3G3PwYcGGnRsKSpir
FtZsdMNAP1yHeoJCIWBsqQwxDPT5cvhoqNgmMHTM41v0P2SjpzWD4PojZpHKncxO
3r5YDQus3rMKAt6DlBkOT3EIOBtznHOVyG8RFKsswTAbvO4ir8qCeI+Sd/B8ENST
Ofj0P1C1JwZ4oc22viKm7G9xFb6/js8Uoovnn1rWCBm9H+wmlqIB3Nbqbf0mraTN
RQvNQwPFF5dr3N3b9bAQ/cHTC2fjOjLyPIL9bAvlduKAF5fFhu8B7IL4F/x9tm/X
NeYZgi2jXGB0hfyCam2ij5M19U0SxM4ljOyXTczRJKAVmq4ajYOoON3CaUY2OPOx
DrVgtlX7wrLugVdhl7+Z4ecmem0uCcs5QtIvXNJhTWHbGwer45iIwYNC/UDiOASq
QF0CCa9vX2ml2p6lw+68ZyqKZUB7kQsOP1BNpbiwtv9FJ68iewNmksp0mVGaxQzH
ghr07qARH+m818kNKe0ApI8CRLNgBqbJFdVllpZcHRBa66jFPINFUkU/pDm5yN3/
Q+c8syFLkZ8Qduh+/7qIy31YAP2YZumKMoDMEQgm0wI9YOeGwV0B6QYUiMtqhv9h
0IMCR5eWPb471+2VXyyt9OtQIeHOvWAjnwvXlGPTJ3naoVaskakyBr3WjmN7X4NF
KAuZO6LYZYzukMHD845GHsYI2pB8NKLKMEHQTUa0RXyBEwtmbEpQrPAKqfsgcQEe
9Vsq4e39ec/8CQeqcfyw7cerh6LU5hjvCKQgpDILLF5AgSeiD3pNgFi6dveJKA5E
GpOxOda4YWUb2o2Et9G/mngxu1snb3X75zlKK7+La43UAIsTN8+YrCmvTrOwduIE
NL1Fhi1/U0ArdjTSalz0iQua6YKPR3ypG6mw5EzdXjyliPdpFf52xRqMrsZj46sJ
4ZFGXEO7PDlTNm0G5CiUZW7nx0iFkmZSvHyAeF5fpAnrOwqT6uwyudBuuW/mVU8w
HTK5iRYud68g+mfBH02QBbI9qVteRDAtAskx1LCZ4WqsLdlT4rJ51Zn7HFeExlP+
3JaOpAvJWKiQphdRqu6tI8pA4FsaVlY2JUb3qz5qtqtpLkn0diVe3pz6FTQ0qpEg
L2ULn2885aOEo/Trrkdhbsq2imIvnJJTjgovQR7FMR33yEPzIbX6U+Mv5KauKAY5
2xl90o15uOVHPNEHcV/88INOURlEmIinO+pi5LNVVmLZBpM/zxoX7olTjaapBWA+
Wqztwgh0XZzngmnoNA8b07C/ZVYUIS+XvWn0BY7dT97vR73pMWIJxQfTlJHTdeIZ
GViop6N7wDu0jwq+8Iy9PWlTmdakhORejDv5f87RQdES+wvDSPzOPCHMB5w98hNP
LkO6Ub5ofdtGfDvpOG9tx0kEtsmzDuAEDzL1nz3SVLwBT6+y2vMyXM2xItWvySNY
bfmD+wgg/OZHVUSmjwWxUnBwrAanzWlte3S0UZvIjn+grfdWzZHC7rtrdH11rjfN
mvj0BuCfG3DllMCn7ZICb5prQR/f4ZFo+3GMG7hd47ha+jFVzV0jvUzQq2YCyJdY
loNRf8ulJtWvgAc/uAFe6MseVxu3n96RsGpGYFtEFYX5MFERcMiTOL3x3yVzdkG+
1xwGpoN1IH+OHoM1km3uVYI8ej+hWEwSf+fDPmq1U/La8+/UZMAGH70Jqst9nDBn
tJMppN7krFaHT5U8+QCW8B5Rv7KMO7A6SshQFQSVmLb0XsoaIXgUh40xXpYOW2Sw
gpu3gG7CqvsGf5Yb00lbuaHvPd7qhsprmmLP57dbBoSIav9PK87pKFQBNsKdQUZd
FICojCLlVw+XwtkCH7Hqg+VpQ4o+WvM6jG9IB2XM6CwzsljVrAM/A3N7SKnOddf9
Cncw0acY6L/fvq4Sxcn25ILa5M1FA3IC0WCPJ/JRkdckojs5XlYOR1/aMIWnSn4z
f5rCmppbAvEVRyo3qKXZYgrhrQTw9hD828z99MC898xsHECMWCa3yPORUcB6ub2W
plO7LoB0mUBx5Uo9yXIgx7amXiZGg5AH1iObp7I10JNjwMmtJ0c38VyHMysRMeXN
2jqjjXfMoNnjpbr7vJc7egGfIudhkm3YpFojxalXTh1cIuE58MsFKwVCyaJ7WP9W
9eKejmEJQzPFhUoIpIS5xf5zZES5l2hkkBlTDt4M36FNOrnnOFAAQz6I89lljXu1
9VU2WOZ7xJ4eJWgKat5pb5xdIPy/UcjDxFoqd2LAWU9stwvTXQU8jv1NNQ9nLJFx
IvG4L0LQ9uKSaq58BL+57i6Uh1cinug8Ow55KrSJKoiwM4y8DytXiyeP7zy+xyvH
K9tKs6lPJnXNTtKOeeHe6Hp3n1eM6qWtsGyZwraDd9NsqyBP1EEx4U8euys8P+vu
6bbQWuczGQg1KVuZwaxJ22yV5l9w+42l+Wd8Q/u1shN+ngRhDulqXIiCHbKdBUrU
9ZbhD1g/qINUcX20aIdH/F9/+ALLmrbM76LmELIwdml5mWWiOGXuahRgtSro2fz2
kHnyOffVX1RRJ5hhukSREF4hOyHI7BP4QIgJC5qBmcW9vBhRIC8BOSkGjwe4yvEB
Y5yDuzn2h+NhbdzxhMyYIJiQPivGe+x8kg+r9xF/mLOIHPECEiUNJNKB3KZJ7q8/
PUGqUIQXm72VVcbmoAEUOXKI180qU05S8yiB5TZNb3IRjHskDiqiXApqv6zZZ+zY
JVQ/mZED1tldmM+wqnB/xzXtknoJ0YnQ+DBQ/p3U4J9rW1BJukk6fSeZsZOP4wkk
/cRWESj7ZvpnVrxaslLu5pxF0wQIjoQyCL5ZrMV2yhdh6UrAR4cE5/scokXa/OV1
2VRGeZCQYTUn9ScMVXMLpyjTM5RElUB3RqDo5kW3YL+Gn1VO6c9mYE8OR7JquPyH
6lzj6FY702sKaC08wLMBCgpAT11to030jiOPNOz1FdqWfD+s7f4ibkEIp+34H67Q
Z1Hz2wh95hQ6xnMYDy2akjsEzZlQidY+VtTLowodZo1o0wyeen8tKP5/qqjJoVro
7OrcFUBTI3mxP+TgcpTL5W8ZanUnvxao4cs5LTdUwSRp2o0RV9x90LYozsC5sTVn
k+ycDY8FUiwemqkENRPpy6ng0u3bOF6Od03kc/nzMrS/4q9QIO5La93bj34MBs4r
AvlSuEYvWk6h0heTjz/nKuZwmAwbmjziPgOWcFiO58FPK3+qgBqSzZuPhFyXnTPV
6icm/vGviwY66uZBXLsw6hnLKPc3UIkt/FbWYIEF+mAS+aH0gk+nimAlZUWkFzGo
4sCgKOcLrA5Hg1fGvfIiveDdT1aMNq6Zi1BSgfT6szt50EQvumMUEHSAkrzr15+I
kbbHiPbzsYPMZj00ynZpiMFOMDEkriKL/gJkj0lPtw4hxX4S+Pql92Prq3E51nAr
oKP9Qw6UFAbObc3xSacoES+pkmbkyW6dcfTRGVsa6TS+SSf5/MwzfrZMDNsTpLr8
ZN6Fu5OrLShaUzCokGleK9qKlDROo/gex8wqRnjl4xgICqlSBVw+nibvEpIVBs2D
tHR3nU8m8mDMfeCIXQ4a5CzK9VV0tucG7EbQK+EMBwIcxNJhTxHwnp19AHtyTCEc
BlXMSU7RZr2EMYvbjpzO4cdUiyY+s6dUUtlhId75AXyfjt1HQuM3FLSjjEklla6L
sDKev6h6tY0FNeeWulEuMAKjBTCJR4MilNtQavkf08e6BIaOlKyfvyuraxCTYYD2
YEb6yOQg3lSYYf2BJknfVEKt63PF0KiUjSRZwFG1XWxsvo1k+tbZivKWlr/HzCOu
cUbojGuelfEWyWLQxnv1xP76RX168TIV7KTb507CxcvvHepVswDW92Z6TajZokv8
OgQksZbEyjDP/6598vWD2TXcgjsymkFHH10/pYeoG1INianYhTYSLusiI5aO3Cb1
O0JrLwKwNsq0lbH+P1XGFPf3vx6ip9wlcxMgINDcmUuDDNEv3HlvrAOxByvG5Jun
AR9D3MtMlKScRnnF4BbOWteGHL+LjC1xdSSP4zjFlIIm0Np5fEqwkfY22n++eslO
VE7LLwgI/LONc+BSqnQ80x5UsXkd/p2x8gCtwvufLrHlOniR9XnX+rkOgh8HwUuY
MAbItxWs/479VtQL5g2pSvyWsv74OiBhhCYMRGUy50psvgW8SZe34NI9XrFVQVCy
I5oZywHi8Lt8sZbLHCOwi4epDu3BWAWSgWqYuEA5z69Jhl5LmLDysG5hBtUqoXWg
EwtMbKK5GIw+IbqsH1m2vpKciUpUXylvIJgvYiwkqCUhAQzzj3WPyWvcd6+JWJfF
7xtYCJD2O7wIiMyALRaOwQ2tMzMhKrIGKC5wEqjm1X7vf4kTQc/dN0OZsM23shHA
CsTC0AyucrC7UYAMFdTZPIN8rKT+1oVWl9r3tVAN1R8ubrGdGhMNZBG5fY3iPfzn
qWYy08mCHo6H8Rd1mwGEhjQS7r/IyyJD8Lol7YCJZrHDpvND7fC4+6ghLfF7d1Zz
uxu9XBHUFuCrMyacSNBxlOKSj4oFTShQVmq0z69qpOKrwB9XWiPYa3COyFrhMyq3
rzY3Jd82JGmZv/2TRcT1UWLlP04zdwpqVhz+ulKgFhpZ2767bu2u7QigLki5OVfF
vcxXaHdPJCVV3WM89VbWHsUKgbweN/Tob1gHCjdnKtgN+tOOJdrbgVbiKDT97Mo6
E9jASaSgw0RfJh4LKrhuBkrDhGoh00MPKJvnWJ/fHh2aQLy2NZZzt/eRF+/qq0S/
MMR731ltWUXZ7Yd3p139y0V8NwPv53b0WVxOt1Hu9kw2h4Hz65faiecZ0YG9mfQ4
tThWs6holY6owaa69FjnrwHgwdu0CdAqhTj9Lp6KXJSt1Ceuhlax46ax453dFNsv
AirI0umtgVr4RLlYdoTGvbq4HzQcyXN3JB8v6X/GKzbJZmjkcP03izY+MnhxcJqc
bL/HKokW2aAmU9j+e7C9oaiYGfGeP25+GeDx7RDyMF4BXRXdWIXMQAtCShx13gXA
gjvaaz9GlJnNJVCyc9JTJHg6NVlhb9bvztVQQX9Z1N3ZNktXfJ/tTvAQzwuAowib
2mEq4uRwxi/UP4OqCIaWDPfuk6RiUDt2vT7CLqhpfqDkOLPkWGQIRQo+YTODkXcy
nkSDXsKq38Nrx8mubGWD4+76GeNE25sB3k5SDjyMlENLXs+NEXRyn3LOjOjol79J
X84Xr20TohwKWhzL+5hnQxIpf3ydIVIyRTh44p3a06we+tahNqMSwCSExeK1+NMZ
donNxvyTd+qm7eRrQfv/U9GbXSeOHu8i4o+fi65stSspfle0D9CmdUVfgpWx+LiS
4EOAPJUp9qah+sf/r+I8ZqUMKrhdWwRsO1jln3Svx3Pt7lNexzk3L7x6ckP6sop7
XxTh59enHWFTxKcOFkXv+YH5SV83ktsLZO8NZnbJURHj6ha2DK4W7uzl/xHQHF3c
BAg/IlNT/szIg9/g3vayAkq5wMiZ9h7jmfOJ23H2uXkywBxw6lqRWKSRksIstlVK
PU3Z0N7C1PtO+12Vi7keqbWWdD5PebW4FjkCZOJIPMxIDeYSPrl1wQ+1P55usZXJ
hoZuUyjhMitnObKMI5JjxtGEH9k9x5xu/hPmDwstu9OYpdGPTlL5MXxmvJC5/p4y
x4KzHZ47DWhSf4r4MovYVVo7D3sv5a+zCEmwPDNOMs3L4ZjPrC0d5ylMExrFa/nK
Yx53ijDfQdv6oY8fOofc8h5dUpzjkob83cHzfeNgmowtAsKMdX/PvUyrZfgzjz/w
aoTRycGqqsDYeyB546WRINSRFd3uWIw6az53LnxaJQgYLcSp5w9tT7j+SB576WyJ
m/B8w93GFzkMc0BSbsGKeo5yyAqdXP5lNDQCtBerVZwyRw9fvPP8PGuGsXzovXMg
yuWoQ4evNp9CIV+ams5K4rgyZiLFNO/BG4JTlPlM1aAK8Hh4MjoLEDzPQRWx7Vw9
L6KLS5i6YwUXG9Da6lHFZrIef3c8NGi93xOyaBF6QCHJpny9anNLnj9EjwT0KcGh
5bP2nIQWsOuHg+VVA5jj6ZIbSOMOzRj1B5xXUvqO/01QrcgK3dE7bTfTwLJzVXBy
Sn59y1Z55omz1cyBrfmOVV5CM/RVcPGZQeVDsRWyumXq0hwvqHDsxvaRH+QPNDix
B4O8ON3ISxWJYFsWyh45uUO5PjNtzOq5Ypqig+za7Q8F6AWoxsKd7cwTDd2rnsjw
NIynCP5W312+sQ9YguAjTj9K4xoROSmjd/9xAjRRfUTDHXUSJ/xDEd+R4YwsvJZ1
TJSc86y/ZnnYhGI8KHxYT1ExuHOgaG6lGEWXMGmBMBVnowcip7W2TkrufG38d9I9
WRKEdnPkXksKGzBCOmusEPAF+7gcX8rwMbfLztUMKd5i84SIl2z+o9nspmJcZLQw
/dqcMytF2DekNJfkcM5oQdEHBPjR+9/v03vlDBWIqLtLYAOorulomfp9Y/BU1E55
bud8s4EN7KHUkoVun3ztUUSJ295h90u1vuWYq9CaWGOgKCF/H7cfz77mAsa7VCjq
9e6HG/C8GOufOdsnl+06Yu/tJcxNoB7cb8g26/mepILxjNsOXzPfZ8dUJ5LDAsFo
NwQTVr5g7T9g64MpaAyFW+izUrJ/ferjsfrV9rfrdvyqwLxczBwtmobHNT54y9tI
H35U+91TBGlsPZLQg4rS3z1D6Pph3/O4DBA/Xb2hfsnlKkrmI/LKEi2y5DnTdkbG
krgUvQ/RkDjs8P/K4AofQdxTpSQHK/75/nJs1g0s29ws/gc+058kBGxhmENOTBpZ
eY84Pki/aPhygK8/hm0rHDupETdNP0n6RMv4eoz++UMmVULMvs1mPkAt4gBLH0cn
5L9DpoJGdgC+xBCFvQvntl3M2Mz9XYiDg5HRm2ijESqsjxQqwfuTrPSrQJntnrb2
AFhEXLNXRn/C2UZmt3op1URsNaYUZMzaYw6Zvm/Kvz1sEu5la7/ZnWb4eCiZFMHl
gEESWe3d7NeN7fymrNk+uTxhgH7lpHjO24dsqCIwAbeT/5rwLFKNw819EkpPzy/b
MW5HqE2thj3SvmCGAEBIcARmqY78vgwPXlgeSFClYiGgJM7aQaMQxHOtxrfPU0qO
fFvNb09rzc/zHwi7+ul5d3hXxwwSyfZuVUfL6/Ps9pjT1JCvuZ+y0g8/c6y7wNoG
iLT4bMY095/Hr/vyivvB91/airIFy3ttvbNiFsEnUs7nxMgq/NwiPvlWPx0WtgLr
MfY8sWIvvjGPjfuC/Se1I2ZGFwz2zVRfc8zLN7Z34Y2YP/YtYC/r3LoTMSAgWqUw
RyG9jY3esWxUCYX8tvK2pqxOrYyUqwlY5zP+yYsyqU1GUDf20aklAyTeE/H47Gha
WmRwH87cjOD3Ef9A6RdPWZWIDdse25IVbqLOX3U6TPTXD1+5FCW8dTOixpffLy93
WjgGu+VXZApG3jTxNzwqNC2JzaPfBmkW3PDJB7Bv+J3n6+S5R8ootntbZ8Ykb+wB
Vb4GoWMyQxyM87bwb3SQt1VdRXpSIXVoktDFoOtcK2aZxM7fPelb/yiWKuGrae6J
+GJ+k+8ibSuDPzmIKmPyXzAHSknblk5E3WRw2Yk+UWBxxVLNJ/cFNqS1AikGp+Je
ZMbLJq4K5E2fE2ano9GSwDMsb9cmo16aufcVlf/rJ3PeJ2BbD4GLYBiP5+taiwgi
6JxvRP5iq/8hCMG64jJBGXB6vEQCV6Y5DTi0yeiI4geI2jLQ0U2ElqodsbicfnG9
Yh00xZtE0SrrtxKY7hpY21LkQpxHGRVW7iu646CYy0usYXZ2G1YwbidiMzJX+L/l
fXwEBIJQxVYGhn/XCz1yJbNb0I6hO2MtJJ3CSpTLCBS6rebbVlnKAtjS0H5//QsD
VSGfmw4QDkDJmjYtkSpAKLKclkfpaiO6fLOiCJeCQ8T0GeorJtNKO8hpXTQQrN3g
m4QxYmnPuvQSpjrBOgqCC9813GiLTfZTTT48tOII7YCDCuMG9W+2NKKSsctCJ/gC
vS9LyfOdFVakYAnkAVCQ/bFUAvPmABC2m4AT2molcvt5/tLwXr8EJcGXdSqVa5SV
AM1Lzu45jhSY1KEbbJh+14P2+CdX04bFw7g4SGY1AIBra72hpIv0xEMAexb83lIL
gxZEMXxRDRm4HxUnWnkVuJ2jNL7tOeVh/6g+pZR/630Zd2WONzNO64d3kN2jBvg6
N/UJuwIG8G+lIjGthcL7YJLlT3w3kV2tXxuRYgFWrkqR23/3x69qAuJRQAZPkvU3
gVOcTU48B2YOjc5XHGgLWgJQmL/w5MUrPhWKEdM1WRHEku5hpk9R5OaXy/RtnCmh
Fk0fADC5pMwcnW7bM00stEI0sD3obeWaUrRLRbJEodEXlIAB80Y/ltwCks3zoJOz
wdNusHaELHfJ/nn/L8SGdnMeD3jsqqXLDldrkdnhSKEyQKxGc8/XeyhlyLHZbdnD
VmSee9ct6yOVnIbh+1zV3ww82mlEZgqLVp2BmhRY/mOtg+I5I7AjfPBot8JWTB4Z
BBOo/rJSqjWTNF2hEnNh1qqELN1U+pXbiygOuCcfDhgzQC7ELRlhZKk86Pb0VQMW
0NpQMogwce6kSmZ2bXifCSSwRaQTHx32Nk5LKTWMfds3DsS2rd9RVUnafnFqjng8
CHOTQJjYn13lf16C004Huu1+/hRaep8YnUyrAZcD27FWKmNxb3rytCgvAjR6pdht
x7km3xpiAiDN5mnVLcH3RYaP0kHqIHjmbAuj81l2HfPZXqFokSWyN+FGTKNR2jEy
yi6i+bcWw/WKkoPfDz6MeOkhsj6kbAq7/bxj1X3wBHZHGHSuRDA4w3WqsHJwVrcj
SoqjLYZTkDKHQVVSv8xXZYl74w/vf+mj4DfyJldVWFOPujKz7841Qe62LCZhN45x
CB/Tq1a+rFDP4RqPI8vfaMHWMmlEbVfMefY0vwAZhd/DiuzId3+Cd0VUtfnxKsQz
I7IWtRZUTy8bML+ev8xZ45wWA6rxU58V8x+yxiVmBVxP26O1mYUchqtROb7Y6Xod
fTAQhASxTf55AEE7gWYDAi7Dr8baPXfYAB9yelpl8+BacCSp3EEy5UhRvvfSxl5w
Q1QMFzzmCv5ePM7tkjInoJdzOkq+wgC2Xy+BrcKceUK6HshtdaIOjxkyxJt0Pk/E
2/p30xEYwithRyLNntHlR3kYkFV8U4urA1ylSbwcB08pvSfPZj6kcrAgVTCsEd6J
QhAMe8nr49aUc85kEj3qo+Q1c23m4A5NQWsyyeeOju3TBrkwpOjyXk89PpoNdHBl
L249rh/q4NQ34UmZfe8fakLR/RO2RzHHmgjJvqFJNYhkHPIhBQOofMhxwsmlO+3w
sVO1UpY5jifapnCxgMuJD4CMEo/J+TQBtPPKW4dEjha8tqLODEjwGfiqXIDYqk3B
DTAweXJNOKBLyefJGQSkzOKOPavyCaEAR4+63KN2NRNXyx4SN5hOB52bukKNY/FW
gqwUpXWPkYQUHE68w5b47xKEzX2hCivGFS/d4KBSBNwKGnVK7HKSMbbhaxI0bjul
7BcnZVGncGu3gdg8J/uTV05vfudMomnpyyEL6OuyZgW+adkqArmyIye/2wM7gsk7
Dm2KFRZskQRjwyXrvbxV3AkuSi9f5IRMoxFq5fqlTJzqZBMnVf5W7kKXKgeujDAU
YytnfOFgAFt50/Q2BD/Fqw/KfEE4/akJEOEugM5Nkm+p61uaDsbLrpdw4U9wZFbl
Xp7yDlnLacMfEXSUkzX0zp5baQzXOQ81fcAjZBqGB//8KKOCfOh9/lef24zl2c7O
usaU3rhRWGAscC4Grf/mw2IF+FIyXIpCJYu6GtyGHVEMj83Pb5EofOVXCEZ5DHSH
Fp5qfKkEYjL8oXav8EQQFsc0CTKfKWV6t/hw2Y5PldxDlQ2RX89ryrJtdGi+QnOT
8lmlrccr/Zn5SNOC7b7iHn8Kpsylq6nSaZvjysNy2vbeDZ9u57hyVllOCSTfdUU1
HEp/RWNUJKlNclfpD2zkoWHn7Dj3iOudHLhuswyFrs9M3X8h4QyM28g/c5dQRhuP
tK7stj26x8HYzwSBrQNy1akpeW8roJAud+lnYxgiRVOlvZkgaaZeKQpHChqegtXD
zVLtkmqe6kHGgqmK/SUO2h9E6PPF5kWv0de29tqAs/Vyo6NDgKGxX4fEYMuFCFtK
NeI5Wx4G+5S9ECQ2CztfPnFpiABP4KtKVXTknNG2sbHvdQt467cQU6uMcx9phkFy
8KQt65Gh0ImZmEejMM1L2oK0cSDM0RBJ47mGKjBECvGoifGJrqNTXLMs3G0L45CP
g5qKShULPYaA/+yLnzJxl9i8Rct7C6TObq8BGaaDhVKtN/CP9kyUhCfQ2oXSqUVi
cLTe8if/ms7/TAEZMkc1v9QHuy9adjy9JaRPy4eiSp8gFlpd2gH0TIR7W2hKS3Oz
csEg0GPeSk17t9V3I4FGI6rPbWcZCZ0pQLzl/SG7BZEUAgZmfnXxLfafPxO6VHu1
VaGH62CSrcvJPzb+9CLs30w9WrX70ti3v1/l+n5l6DNfkD5fTruYsGtDmQoccPQW
dklrcWeH6ug/1wkLs/RhoJrg06CGXgXotO85HUGz8+WoXlhm7Nm7YWdtgLKbKeRN
Sh8Topa7SB/4UWmO75EEFuk2K0cx/DWNd5nUF8MPD4vBqgMFr9sxY+lSVQNaosMJ
9sPpELttKvkTCzBOmBYKHlhZwxtFiNJuHWTQPapWgWmVlKMOUoFQvdBCMl5pyBU3
yaGyssu0BXISQmOGXA2QEpFhcF6TKBokwcm3ryr/RUdbtoFMeZciLBvHsTqxCId1
T9AHoGmo6tFzZllCPxbTiMlt9koc2Pv/vVXL7xawv4cZo+6Sha26/dkhzc9NRpTe
FAD6/0ICH7KAXgAJEa+zptRD/M/LRe8CxEAVD6VueQy95p1theTRb2IDhrLeJaFo
n6iaYc8WTxhUVLHc2PGbMsmNeKEcTyHD50BUStt9FdxJD5WTAQPf0u5/SoyYVese
lqO8W0JsQicE85qzEbSagimfeP3rlwrrkxOnOOVUwSueH55twgpKSthvbqvu8zEF
3dJWInuL8oMpYPPKctpR5rA5BSbWwIbICt76Jqk4rDZRR7qQ4DA/y5vhDSPEzml7
c9TfeFDpx5/MI1E9r/FF9OB0P99GjSPNxbPy02xbYFNpQvcS1r1ilSmETmStqxBU
LSL9qA5QtHXg6YcnBt55lf1oX4MBttmvgKL1G6u0YuRtQGgPS/H5R/Zjsdv5oUgL
KzDOz0kVjsK/VwCGZVrWrIDvv8CWJYjkv75QqGwq6o50n9FSTsyDG6LcoSz5qnaD
OR/htQFDqC40qVp4eFZkTwjsk9YmGA0udkPFuyvnXE4uaqv51MYXzTIg/yzSPdoB
OzWeOOCgRHCgjJ1WlOkq1eK4QGfAUJCkit5+6TYjuanRoOKSzPV3LcRKLpCG/mDn
f1UhP5Do++Hs8PsNQ0s2MaZqPIvhBJ1j1XJANu+kdmrX4rrHbmt5Ek9xVk7Ty1mw
9lU54IPxacRnMm79E7dd7Aqcwb+yvYGr/Xk/kFVD9AYjAXIwhKHKhhAVbJ4we/r5
joKbFAVKW32on8qwb6SSSh80SK6VTmKJiwhfxYC9rf+LA3eBj40d1QImr5gBH+1a
QkeNrP470kq0TnhJfQ1jg9gCIL4Fy9+zoRiBfBEGzLAFYHsKJA4Qq05ZgNa+YtJe
T7WajSOk6mpj7SfbgIuk2JQVMk7bEhM5/8BvzylEVPX3N5VC5T5BuTxhBGGlKuKF
c8JbxF8dNq8oSTHlR/kMPTx5tZJMPWusKkzyxYHSduy79a68lOPGNUf5ANOJSktf
HC0zkSwL4BQ0LOdo/2Wu1d6FfnYyS14PuGe7xznfwMx9MgBv70T5wApSHHyPRwbI
qRQGDmCCH0+7t2ez90vFQemc3iNJ9kqTsqCqvEBLMtEO3jTMcWHWZIwtc52QHB3j
blOhDiIjjLysgDqU9p2cNb4WYuRZ41dYu76jjDTOlZ5N2+EQv9uFzmKkGHfu8QFM
0sQzzIi977r3J2i3JSmN9TOnooHcVGvWY/dW0pifxH+1qRAI8A5Yz1LZDp4clFRV
kdISpYWjHwkuZD9RWN6Jva56T7AGfEYqRlv8y3K8gJCl0Gt7gtV2E1/uAqcRqLbw
0peXz+HNLFjUzR87XPuvykfBy3+YynjJThWbhdrNyYBNZ3ONrOnAPBjJ29ImNc+S
+HDwIFZOGKS94QHDDfOUFZR85C4BClsHNbYoiEEwUm3BbgQRvcvrnWuVSkG4ai5y
SKf66AcwpzYEn8YbTz3OqM207VLcWgCnqy77mUMjXjkJGDdUF3Hlk8XHh9kM8gDX
JkdUAFb8Qyu/3acpd55e/JAMkExsaZHZrx0qfGj/yjj6nBJnowa/Vcf3WXGsYFuc
uzkex6W4NwI6sVFyK3e1VBRHsc7wNffHQUovygDkR0cVmySr6Kf1R2+mPASlDtT4
YPlSIyvo60dkjKY/e5viZr71CXu4qsh2YzhpzV/EoDprVVaJzeAfavVzTtrTWm0z
1CF7SY1Z2OsOVswRzxxwMmp/Ro2LzPV+P2iAtQd/CFFjT7UXbRtQoIb8d6RUmInQ
+i0wKwsBUbJI8gaHXFl9FP5x+mieOqHhrCJnvzqWIuI0nzbnChPa8imRISxK6WxD
WfOb9O7TraYBXwmrUqnLNxsA/ACMV7JtL54kG1/428MhDxWwLgrw7x+tZB3oVLzS
GU4ih9gnDsv5FJQ8wHfRZ2oY1JhdYqhsf0jd+rhxxCoyoINRiE15VGRF8nk1Q3tf
k8eV0xOrJGUl4vl9Z7McXfF5jknzM9w5E04tjS4sJQB7YEUVetAB7eWd5urAX1j1
QDF1dhpQCIQh5NGbKEOzTwvS/DX06ZoD5L5hdZEYgJ5+HUiD5CnGuolSOVFAqFd3
vNr53xKih4byDPizo0DvmhtGDwGp33CmbL82CNj1uVCKkSjsQ7PImGo6E7MHrL8N
jr2s2KLMUKvOa+jpDnDiXyl6AvM/49hCO9xKA8jmHRIR9X5B3cNUEmFzRm9j15zM
STaNpBznNFrko4oxu+vuw9l9Q3IqU+zYUlGXS8jJTFfHmK5B1zaGuoh6+oqjiwCL
n5EqIGlttGZXvWNwhtVVNaLaRwPUQ46TtZcCB4JbLWIpXAmXtzUan5cNzD1sWqcr
1YlFNOOVkgt4MUokwoIy5kJbfHfDlcrQ0LmCdYV2mCEUWc3EemW6izhqyBF0/mWl
FGLy5sphJsHj5karjsiYTvXjVWB3DnSzHuoKHCGLEQCkwxt1efYK85GxpSy8gJ8c
D6oYQ2QWqagGzecPk2w5bN+820CxMd+htOy/TZGzx+yISVpsfQSh7Z2eoTMX5wI2
mvrWHFzhJo/EDhC0MPi27Np2dsu8gRcDlE58Uj13OVCpENFCBEysdo9Dq8qUgw7e
u7xNELyR2HmQSPn3PnfWFhhtdeF3mMrLiClQ9X+kh5jBlmjfesORr/QgQEQ2L0vm
Q/yiA7BrObqiqjNqH+BhfPb3nCkZfpVyGQH7Nx9B6uw+J1QnDPOcrWmPiLpai4iR
T2kLCKWDsRzAexSt1AY70jmTRoDs0bJya9T1nNq1PN1VYEAgRKwIvV8OjQfVzzUX
dWMUWDBhlarGPJs3dHMAJ73MXO+fjeKr0Jaf0SLgn98xMhgIS8xohGHHg4PDnNu7
7icqud4VEA9ZAfReampfpuNkHdr3Gt7+2UGe3j5UlziXGkATc+IEXOBmi90BSvff
76NpvLRdXlKdyE/+krVIwSusAeukFBlCFgxEkjQvIs5/VEblMqbRxdTr+8PQp1mu
bu403jhdoZeP4fq0206C9V8ZSuflRqT2di1aHmV3Y6PZHYLRkm8XhpTNJS6rNTsD
bvN7A37yQm42plbRFiajhjABwVqEgA/DWGdUB0pAs8o55MFDrto3wYS8vH+VavL+
ugaNew/K8/S8OvdH7IED6yDBRSLB7bAQHffGpJtaayt72u02Wmix2+tgtOM+6MVS
93EeZWGbDwq0FSvi13nnxsXMIMbWXD6/CueNYUuGbE728LCgOUlMD3eKVDr3Tke7
hlTL5f+kDKnJOL6/DF+nbSKdC5NRRP45sdO1BfxvOtm7ZC3cZ34qG8OXvQyFXpXw
iNeoklcFTATLW45k1NNHdElApA+e/xLcJz9LsH3FMv3A9R0dBv9Vos5bTpZk7pBF
G2EVp2LPKdSG80mf+rBaZYZw4Ncuev+vFfRyhQT6ua12/vqLP5hF6YgfmAKJJ6Vg
xa593RiVHHlYK4FYit8V22YolxtLrVK31ism78gH5h+JV7AvtA83flgm3u4jAwf2
S48jAM8My40OzqslCdofJWd2xqHDVIlvabAeyaBSZ7Cynp0Jod3buUAF5ySZsnHI
xGbX0OomXOnPzsKLydvjQHWA/ePubGCL2lhPlYd7LuzdtmGA7ca+teHDapl6TDci
lWuDWPySakDW/qVFTnpuHvhcg3T6cwoAHoZwoX034RVO8jcX/NHuJSj1mK76oh7x
bLxDuVy4OepX1gbZjsScpGyQ1XvY8+XHaSiO2/bLsADB30qmiuMwuAqeLNwVYYsW
g5CMGnYXhKgQXORWQh8Fa5iig1KRpmj45unCbEZIclsD/tcTNTdBrKrou38uhoOw
RXA8IxI4C3T6i18DkFBZd5OA680UjR8VOa8YPF7n2JUjennDHEYVLq0kGFdRS+3G
xWEw9L6E7ESfczdecqmVIE0Kyeo/UyDvkS9bg28Z7BMlonvYGpOJAtzVqIkok3rD
qkfDSOliyCRwbZVvExUsbRc1iMhEDddZSig2UYCcn/kri0pjKP1+EREKmVCOJg8S
Xukqyg8oh3amFV4Y817ehYk8mi3AwWGl1JkSgy1YC289cZda+GI0pr7i2FjPC850
yUiA32f6TmU5X1Nne2MvDpISGKwcwDttQdC0N9lJ51Wb5aNt70x7FtG10TNoAybM
HKAAJbvG4DyaaWZPeWNaBoLNeHhdYmadkV2i0/IPlA4Ha4CXH/pcB1S+BVx27slI
kJXvMkdReJBFOOKR9aNkrjwr4f8UQbq0UaH+bPkcT8ioVivlXEPKSca83t/AvUvk
kOiA4t4ewKwIDvGTxKm+xQkpc3Rz6+g1XiIuLG1HBCNvoYnPAp0ZheTKKSLxjy+y
YIA1H5fY/jcahAtHD22ba4HdWoKfA79w0lQ6nFzxuQXcSi4Y8+wt3UumRX/GbCVx
CRVrMdeg7mlK6UVRq5Fkjwd8C3hsVN09iJaLKNR4raITXZFbZhdhMFb1vN8FPHFY
EWqY8G2VzwIDb5d71C4YodITxsKpkyrxN8ZsotyOaJxfj3y2EIuXA0e1iiLdjI1J
9qqusGexBFTT36jimL4UGEptQJd9XC6oRbULmuTLM/1a+iEp3IZMqk7g1ZHfGdlT
1zPcbpuIG16FqfDdSKUJU02d9/2CaZW/O987M7m/a5EgiH8TVV7OtyTS5JzAu3m1
AtORc0bjY154aecfeU3yUrE3bNWK78vSPkw7QLNVwEokzOL1Dmb/PRXPaIJFG8wa
PhgyVZoKR/jt0nLSUmEa1p4kKu8yqrIblZ6Th+G8m9XbWgGPN0LNIL2KQCQLOuKy
130eZloBQcpcGWr3fBZ/99YCDObaQw4jpkspNO7nluRiwdd7xV9XJjZ969Z1vd5E
Qq7QATprD85yJrVEqpiBertYeaCDE/9/fp1eqb6lAXo9DV03OrBFsfnXuTuEXQu8
2xo9H/1eD7yrD5HL9WX1Sdz60mRIeDlTNnV3NRE45Z3kKD7VlqnmswMIXyV1cflZ
n1LAJQyxe7LzM8TP7aiT7as+dzzaKOrmxAn2aws5Asci2505vF7ZQa0nrMjnqS3d
DZyEWbv01sX+oeoTEVHtAyoVi6EHOlBHgLLqD8CgyriFyAQAQ+umNo/o1o6CRMDP
FMk14YP47sHNpFjF7CWsMYIuHuiASIArVPS7tP+WHdJxhRP+xOpYDsGFpG4kHLei
lFW21Q3zpbiJKQ4sJOIcKPMdkoWgbSHyqeTTwqJspQAUSePatiLFDD5UuXO/A9Om
Wh/7ce9/2I9limlRg0/h0yg1ezu3dnI3+K2gY+RBcFs2nm8nlAUcbxAhcqN8mzFL
IkoAGchLf6EM0CDCbviNw0BOnqEL6tb0pL5yt8WbQ1JhDc0JcTGYK2F/gcxiqfXT
p3ECWUPPortJLoWXMLLZ40ONNa0ubuzxQgL/lTA9B2wIaFsd0mCAvy0nVE6lXAkp
yioTNO6Bglbx0sWcmChRpWFg3zJ4TVhmSxEgpB2E/SudiD/UvGr2ucXT67dAIVWs
tpJTNyOeBTWVExrX6fF9eY0t7JoUDnxwBO1RYIaEm8zbPciUeZa6c/HWRPkmkQAE
RG/cwbLCHJRUKxxBBo8SEORhtFDYleCBLxXJoka0kCfw4ir7iJM4PPcmjHUwiNJk
RJBOGYbWc/En3tXlr6vXUEu1NThu1+rWEzmajQZ0IHCsA+2GRrvrnP0ESbCCLRye
Sd9shyeKaML+Qb4C2ZcILwpQSarGUuPSPSm117ms5qd/kAWxeVBtcECL1a4E6OI8
KFO7qXIYHCwRtiICzmk07ZOUrLVcxNs+F7FThXOzrnuLVyPXUOU8efFea9glko9Z
uSoREfOZCLjpZ8rilezoKdeXJTXYiI6PZ333Oxf8yPkhVsCvv31DL/ofZC9rkwoD
GtXcTjWrZlfvnNPh/vl2J3zEYPTR8MiAVtTwIX1xfL/kFNtSZ3Nh0043Lg4PkukA
/ark/N/DXzp2F0z879pGhGRVUWJR1gArNhWttDA6w9CNYSzoG05WNGi2kikUQ5i9
zmwo71JO7PUav67huZCp1bFvYd4QwavUY+qZR3yut6S/5WEb7VTkUBfzimj6yiDc
YGQox5ysPXD1WWELBzrgcrsRks62h0/Rn/1DLmNQG/Od41YJ+cKF47QL2/H/rYG0
ANBKzGgk6mY6pg9eJ8ZBDYKUcEwQYVy7cYNVltFdu+YRYmLUDOiulzhjigoxha1z
uq4GlJ4rkgVfpn/XBO8i1l7ADfYGoAAv4TtXlR7HIGZttSvvcdHF6OHldgz1xFO2
Xffm8YscPlecxk1FqROcMj2RH5XweCq5GJWKdqsLk/QG6CTcuNoVB0ah8HN7S1Y9
vRBKFUXb0PVJrOlKdX3/RU9ew6zNbZQgp8dxVXqvyt0+Z51/lOhj7D9iG3WNwXQ/
OHxZ56x+UdAhHWJkHwcx+qda1u5yPOKe9Pauf9u1KhHfRla8P6bWJ5IRlTaVC7is
CUnrwDl/BphRlIBimuVgOeh8z+aysqOMQ/gEr2JHrT3AoJqUIffFpLOq6SX3zkBs
76gEpNfxBjNy4D9H8SE8uAkoqvGhIyLeGNphFxq2j8ghiS6rn4qv9ID9UeUMb/bS
4vRRRQ0Iytn8TG+fun2ENUx8b82OGTIPI5czfnPJ9RAnP4wna8kqBXSQmtepwcmT
zKCtv3lzONvYES2btagyB8Q0lbKdHwLa1mA67T2+3EIb9S64qvh4djZOS0NQf5wH
TS5fGzNF1j9Io31mC6GEwJhnPu6Z9B/FOWh+yzmhSxO5bZRoBzvaVpDUg4G77ey+
+n3S6aRTDPyHi3F8JQ2rV4jmNdB/PQ8fuXVslt2lAEf6s/+iH3G+y/KDnUqAneP7
/nDAKcJR2WAXyLZdJ9tBcw2lu+8tjIdW03F9s7reHb+CAQAtBP4kUf6ormA0NKOV
Jzn5M3uAw7aXHy7UcQ655Nz/UY50k9vFjR6PoO28esP/kKkRdig5IMxiJCpZmO4I
EllX3BMIi/dOV+j5Nky7EoyCukXclhswAB2EsEF6EJpUYBYskseRZR1mShyK9w+2
Ewlw4lsDs4jKuiGTnzsw1vNPEFc8/T4/Opd0N5dDyzT4PSobzFUSSP9MqYpiMijn
a3llhqd19qdWRtTwhi3I+R7TGHlo16Nl+rFM15dGQDw+oy8eEulyXeeAmjrZCDn+
ZndrWYWR/w2wH9MpYOgeQXmOoQUouj2aRWCaG4Yd1RqTeedv/U0BwgIP3A1mHs4m
YpaF5N3CBafdAwCqIKjRAPgKAWJKy4SynZOR13jRJYRVGwn41n52/LvJx+qmhodc
IBdDQSPW8peLyEN6DanoDoB/EpfaJo4yODS310Ys8hsKbVfYtSr6Q2OMrUWb3kZ/
F5ZRikUJ3TavZH2QfwYDbJQ48ti+vTNwJTz2zmx72T8uLvBFp6DdouMC9IRDu9lS
1KhDL3+eJU4Jq9zKNnx+rU6rGY1/cq9yJomWol/wqGUeJROcEKXOSfaOd3h6wh3v
9iLVq9suyLt7Uzub4uoRfaPcTnKwCBo+onuYGFdgk42Tg3qFTX5NOJF2JOMsl5Us
rnbE/Wyt6NlFVV9yV/XTg22TwJyZVOBugpceR0dTweeEli53iqqO3iImgWCaxDZl
aHXwQWo393cSS6du3wbxS6norcehhcr0zANDZTnD6voQFxE0FkownmSl70Uw1fdF
dXO8KzwRAHXGSd1qoH9Fo5lynQDZKs+fyFQRKAENNAdLjDivM5ImsM5rZiDelOCv
iiRrKeNIfnHDEXmozGD43JEW5TL2qjrEKloHQp4MR27egYiwFc5k2Qx4VubaV3Kp
LZCmgisgys/XKQxVyBZKAXmdKpBkGlbFw+MlbknR70eW2JIgdWF+OJd+QIm7L9y/
BU0ty7sKGxGeqApFGpOhahUp/fi+R7/gi11GUIBRV+mYkQqfao1Osjh2BzZX3gYX
RNjyEfEA41GeJ4ixujSu4xZRgQ/HWdgRrEkVs5I1XIX0tCzqadWC7erNovYJZCv3
1OoVXr6RixNEc76ztGcmi6Cj3ScqPZQ3PhhylfaCkv5YxHoUTornJ3ctalYloRY7
tyGPORrtjqfnErlts7axJHcxDL3gX/W0c5SchhBMMI7BHz1KwFvrQNnWIkHiXHgl
yofAxN2HK4bdNQGlB+u7Kuk2nl8LZMV+AojCrnf5WFppGXoV/TwVbf1NMgi+TWfT
xS1uLR9CO5BxOA9FgbxXXCu867Wz4VX+X3aVkOJ3mdiLanLR5r7bCa7ftKm2Gog2
6oNrBi3GNRG0YrHh0dD4J4DYMACG7ouc3chy0chzhCeMIRLTX7pitu0waO/s1taq
IoTdG0Wmt8e9PIIHVQMkdYXF6KT1WvfRSZzfRFFq5woAx4ctGvNVU/frgIr5YY8R
E1KoH+b2Hb/4vn9j8EkuqRxkLXNzrUZwYS3Etps/xnIk9Hwb9Elt5lVg9Y6o8NVS
0UTFbSNWJQls9ugrzsrZQff4mpoP02L9pYFhs7xwgiSf4ZaEBJyLJ0swJMYdFDFN
rfxUvmZDlGajDqXKaolBL0xit7gdCaKy1HbGaAwm28qhUBeTm81oKfH7BRz4QG1k
CYNQvlK0gDG/0dPX46IUSsJYozdjBr4xIcOYEv14eQyWN7+OLgzgF64osnIrj1tZ
BfJcoN+8dy8Ep88xqHVNrAgv6MSEyFCMFlCGXwcgxf0nK6RmRxX3nCC3gwRQa8cq
r5s7gUTFMNjqAi08OGRt/hA4nRWyZ7EGZtrqz2Ta5K6L2XlON1yYPAFdHxG91em4
KaxOah+nZgmjEiniyQVvCanjHKbz2fOF1ztYtPV5k3w/CS54PMmUxNEuk2k5vY3x
1NOtflD7myTv/rnPpkES+ZlOqiPjwsqXsnjBACHZiPOE+IxaGudKAqBwXOd2Zrd2
ti5xFeTz8W8bRMj/YdgU4i7nhPnCOsQQ4EaSH5U3cmikRuAFLqRoUXZ08HqvEnx+
`protect END_PROTECTED
