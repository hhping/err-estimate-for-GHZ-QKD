`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/bQV+PhOtXy0gbB7HGPaa01K1ZmKrVrG61NEmL6a+GcmiZYCSDWDrNf4mmB/MD/T
/GJjaZ1t23wMJaZI+8xT1upgUJx2zy+KNrAm/sMN66+Me1grmRw0aW0OwRXw/OfV
fEqNQCkckGtd9iZwCWVkWkhqmOdBmHoqzABtPaXvmg07CPosBmXbJgtch5wSwEzg
z6jax9kYKmZ6dufYxHBKE1bHYjbdxqZF17bOKVyjs6/jn688s9+HzLVFhLYDNp+h
I3wtsTqyJ0c+IWm1/9YI0xwDcUJ/LhXnnD3YgVtI0vm/yT2XQFCD6JyQ7cg6JNkc
HDjMyz2mYR1FhH2FZ/CHOzI1XqUchc9T+PJTtanS9qpNUu5BrmTAHdtVpFXMJuF0
ob2vWOFObeUdeG40UJvGOHN9LrAHl4IW/lCH4WmW6fMpe7X9U6F4tPYyRX3Qcdb8
FTuFI7a6Wr+lMog2ASjHWHfOxOiRvkc4k8FyGpZNq9Xv3ZaeNsxs9GPeh8QqTT8I
BExEk1t5M3O8k5YPIyD21vupbCqiOyjUCQ5buoRVvq88nmrNPhKgOjq849q16DRD
gUirfStcQswDEMzjPtyvj9RY++o9mteEf1q9JOwNsXrsbc3WMV12dfr7uhnnHtXK
8HjBMznH2Kuv6ToEgmeExK67T7iF3vZ+Et348NE7jJc=
`protect END_PROTECTED
