`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a2yGlX5RpR8a5KFewbzzmMAbOadhYywEzQaut3E9tzdxUq38mNIKlNs3zYTZemZk
qG2Hm8aIieUdfoJr4y9XO2K+q+kztXg7U9DSbSilSU37uxnAII79apAB+byUHg2Z
b+dHWU//DseqG+7meME1NFo7ClfhJ0q5VeF8oEiJBXqZ3+PW4MRlzpvFG48BbisW
Cj7icj9t3G6EjbmnEUePcXty2FY3yAajMSwlGo530hivmzf5bde8ckGHc6yHVk1k
tvNvglYFXcwkKSbmPy0a7Kejf7WS5csI0Fql0E65VUDiy6nIgsR9h9wftLp4o+j8
q4SvLXOo7DEQhOUPxSRLMCipJUu2mXabEPgsbmYUYi2ipGAMvzcOvp6eUReig9lo
+JBvYyOH1FT15CQJEjsINvjZy+fJYH+KEtyVG74PzE9UlwPci34G0LpL7u6eGs3E
BH2Lgzup9xu/Oe0Cku3wCQy6EAueyXIscwHj4xK32Cl7zDXd29sGBO5zPNp/tKd9
NzSTp5aVbI5CAdHtyxZhjzidak3XVSyQiiwYX8G8qJ4+vC2hscSt2WehNQ7gAEC9
oQ7wNZw9sPwYR24dhZKmrkxfpfVZlSWczByrAw+EGv6Og1sCNRVaqu8fuYMueKME
HmbwiKusHN07XpitQvzzRSjHCTYpl8LgXVEYALaxhsQbjtOB96ZGqRAUr5mRdUSD
AYqfdCYN13aO2OdkvD5QzqjXyvSNkTa+6ZSZc9WUnXzzCun/wkqMk8CO2cr2+WXc
2Y0xn7gKdE19SnurefbAo2tUTZh2zPyK+8oCOkhsOM21Id6BzJzY1fgDqx7YQ3QQ
9b7iUQaQeFB3lZDPFpAoHlobr64jN6H0S/6+yh0oqzdNFTdZmWj+aKzNeqM6pp36
v397v9R2bFoRYJ1+FDZ2GQ==
`protect END_PROTECTED
