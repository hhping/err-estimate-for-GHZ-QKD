`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P32GEGH2XAeHynTdkY6Q8EID482e+xLXL5CTC1cvmaSXjcmFHnkf5RTsOktaq4x/
1sqx9bknnsKMPR/SXEUF91HoixLJsOc0YbpwP9fdIcF0DDz9lR/oGTTQg2Lp3Q0J
8zqtG1IhroFZwqiTtpG0rGkDvZH31OCbRJIBRPzLvera273wHfd8L18+oAmb9hbn
S+BvKgRS+Oz0pXL+FQPnG5ClorECqj/lRpb8vUykT4DCbXNGeDh0ZM+Q6xf/1hEY
CCGd9A9+9uofkglgOQkUog4SUYhS8hRZcK/JISC1u8Iqc6UJhVXByPkYupskvUls
vCHs8pFBW898Z4G8Z/LP+ekux1Mx5nNdv2rEhB4eCY4PLles/SI+gi0qna1pBSAM
Ad/P+dgU3Em8gooi14Et4pD+oAIhEUBENJmk9OWHS7A2xd6g6MQy2UqlXGGYBrbI
Ph4WIB+bi7r843RDTkikv3klgVZPAUcKBeCjDHprJETJggdDfGVxdkcTqAYJkWjD
cQ6c0wINJ9WCjTA1k9CTQprhqvyRSCv2mY8uVPvsu/RiPbxW3AWZ7YnMPTQLiOay
z6zWxNsQhc9iZVnq/o5Va3OYxMEANjscYio9uPL8ytSSfy1jp9fHF0jJyv72j/5e
ymVvyQ2/PHNIChwWCi0LPfDUU/xHOlkaocrLq6bvU5GYYaU+6giynuiqY52kC04y
3YkvSJvYLEgaC9ZRFNASL/1/NZOY5+P+m01Fgn08m3eTBBob8yyJEemMrYieUuWS
vhc/5K694/KgltwaVD6SLcaqKUy/rKrco7DElrqLF05LY7da47upYt/srl5K9aso
nBWmVQcWnwgKJ0/9Lvs8NYY7H6htAgPj+r6z4qsqRdocuUU5qgqEs/BWJGAwfF1P
kZnRknWp0oTHPzpUmFhY5Pea5upOcCzlbU9Dr4hOvDySaMQf4ykzHyj0jD2qhqcV
ZsQhGX3BJ7m9zCICa0l/eZ8KYWD9l9j7RPJy9eeehjPlhKfy61GaTmG04tD1HKob
H2enB6X8LX3lYFmKKiXi8nAIKsBME2WmA7Iul4dvHL87AoFI2Gy04CgvTCWumeVO
gUsn7Sqb3xlSrkDCKkNjDjjNy1SPFtwzn09Oq30yPFdjuOEC2jc8Mta8wDpPpjuL
tdHUDkdr00Gk62RR3tMd83A55VMWYcIb1Da8wRPtOkZtIVwSpwAYkc989EB7tIsO
nx+x/ZER2azzEogdvpP+08ErZpy+t26x/3UNrseOHKiw6yck/j8Ms2+FeiMLV2Bb
`protect END_PROTECTED
