`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nrn7Qa1Tk14ViwtAy6Rx/Yg2CfIX4OYf6R75GQo2HNu3ADkosu0Bp4gPH+oKarnb
aBXYnHsjW329uj8HvQ4DBkWYZ0Epuy8d1T2fYJXYEWhNDon8JPDcHyYd+JCloCNY
oLK9KLOywEscR1Do5/c8Ho9L9v+txjpNwuInav8dNFD0gm7yFY6ng6HOMQuqMTL2
c2deNdNRRcqzni56+8h3mrLCPjb1aM2w6ecpAq2jDV03fNnBubi+PNK68NgNjtP1
qLcsS6dQQ77rMzqaWoAsFSUUIEeu9HqVdpyuCYrBR5Z8bcAM1wnQu9+t1apQ3asZ
0O+StZ7HqeiYDIrvxHceHWsjwy8bfYQoTNpoi480k+F6dUvnvcZR/xTOg+RngwbN
+XJEY5AmRjq0GLr3qnMf2Q==
`protect END_PROTECTED
