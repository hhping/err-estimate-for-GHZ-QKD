`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iWA80NlB423n8/foKjVWoYSKbKto7zfP20/jcNXQz5vSqBOzEzOL8a2uR6yYl9pS
X76AiBvcNbNy1FKhpPr4cjmn4mMNLpUvif/XUsRfHYypXu+8VTvaAlRvGZlU3kJt
cD3xHSRIJ07+IR94tMIWVVkO7tpUQiyXqEocTQka77VfkiCJtBmIKXsRyMcUO4A+
zFKZdKiXzWW0dsOokPJSfrEb04Z+YFwPtLM/4rrzkJFAtAPgvEHfNpLYF73TdNqa
n9oaouG4ph5tIjfo9b/eoIMLSnRaasGSrGW0NBXl275wFwQfTJBEUjNR97IrasGh
FiW+aN6pDvM9PeJFmvDjpaKUMkKT3mqbZOi7T3U9XuGysWhEwmYymh1+IxmcTZUR
oAIpS/fvtxb0RX8OibdgYgO3a6SCUZaos7/82J3YrnljkCKepO4c7f+ruT9TaeWm
xmXqjvCDWBQf3/tXmzBeO5YCMBPY5+ll/vDlRV8ItsH9jZF7yOdUkSNc8Hvjnkxh
rIY31jS5cNfNJNGHPDowaWjaXK5ivdEAzmIurg3oirZ0Oq1w0WEXI2KYnbqYolYj
qqXjIgxulgCERWqctQU5LfWcv9P2xl622Gj9mreKsZOuwd2IIENK5vG7XXj+oLCa
K9vVtWCz8ydTF3LbRYYVFqdal6vnH1iiqvHzFcV9ULIElYHCi2LfCDHbaAZ5PdoZ
kROLOQnp67Y5zc+bRyIkImpn2zQuxD/MIkfgO+upAbxTiEek4Cv/fD4lB0MXaeKT
gUoqquuVMMg8n426L0c/kPGJEUSZVaTsVFe4u2SiCZ3EG8p1N1KPSA/zdqRQdvO8
URE0NSrNBjE3VU5BLBHaUfwJ1URKTgaXd0ZplXtcbPFqL5O9x+G+4EyM55hfmjTO
Jnn+Z6INTHxFl7HsFt1afFqDOcgmrh0iJbmdlaIyz52epLjy8mZNiCkfmw39O8WK
FoAkrj2l78n9FaTJM95rX7ipkl8ahiWG/bDz0DnNffq6HG4Tp2+6jvJI3pUJW/e4
+3n1sDmpsmTjoZorBwrR+jaP8R1vdGQ0O6pYz3O7w+8=
`protect END_PROTECTED
