`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OxDUYUF6jrnJz9DVtXrBAUDqV+yUCmAC7HQUhKtd/ZUP3NfpNqAB1+VqTviFnAPF
bpFYRvt52zM7o6hmYn5oZjTYwadNzv2wd10xFWqtH/aPXK2/wbsT5OClKqFbQVXx
qj2skmrPx16umiloY2zQK7FxEZbl8Xp8uysqplzD2Vup/ipI3apMmLIN6VucCTe9
jpi7wwo724rQt6AXBvd4yjOa1IYTGlqUuz5Yt6vopHskqWiRknibGDigWdGv4Pkv
O3MdDbH+esu7n7s7PLCxwlFKIMinhpkZGuExHXHxZZEu3gjnTsj0H/TIFF0K94UR
3YChxwkhaeMfNDYJ/rLiNl926xaQ+h49UJVSVuXQk2wT+/ZEkWimmmIoxwEBJy8G
pwlNW6B1dop7SfPUVFjaKpQjIKRbGY5RObXdw2jLrgihOj+7q6GbxTnuxJm9wRKB
LsYvGCDgLO4QkyZabCyXleLDVaRsIMWF0qwS1UXqCns9BTSSCb7UrIatuCyg1Xdl
BV7ZA9p5ijsEbRWuFr1a22psASBh0lVlC/yfKKvn45EKNFm0yUJjFptdQ4R1OK9Q
tq1UqJblGsW52ub9y4fpYfdEVRhG7kIJpkSUPtSJlMezLUNuTeeLotyWikAdAPk/
4kbonWMWzeRx8mZb1Y+jU3zCO57ttYuEttXaNbwU9cScd9wFwLV8eNtO8LE6Owj0
/t0N47WIsBYMy+rmvdB/MmaixbIT3Leqt3qydwa26m3O+aLWtInO5F6XSXjYo4Dl
t6mhh/z0Az8QffiUPM2vUeaoeORv6ZaZH0+H0gE66gr3Ic6EhY0adhs6FWiY/lTj
vjyq+tzGnH+PJqdXFzfrHkTfAnQa5H7MMaUPplv57h18ocD5owB4lj8BT2m1GqOV
VlF6qaYFgSrd+1Lczytio0ZF1PrUfYXnM/YGO9llVU4/8p8J/ODiqb3dfEhR9zqw
enmbH7B2PI4uu0TRok6MJ0VADfdfmT6Kwxuo9AWvM+y2T95Vc5xFhK16XU/3nkjR
hDgrpHQl7DgLfRE45lUXUZ+YLyIo5m4pRlsO+NLIsJb4w3UsbD6WN56/+XIi5qHm
opmxAiL+vHpw5fniNOuVBlVq/xq7RZh4vT0QBY8t4LAnNfaEpvOdjhPZNvqEmS74
DaypUIIT0WsLTMfwnViy77QPT3qKrZMNtxLHrKhQJMtXt6JV+DRKrYGVm7tdhENX
DNNsKFXL6MIlpkgDnyvsbUaGkHP/8Xrp0O/IJR4UC6mqUj1QQbDOXIVXo0feycEv
EgYeayghQrJg8gCQE30sToZ9+aywe+mpQ61f6w06ay6i68l1asv3l5NciJSzyIf7
RKPJRA3TSZXXdlfzE69bjLE/YQpDQ+Xry/fORjYt5Pe/jKHY5grqlTsbggdIK26w
X/xgGYI38qli4fuRRYeUWaJZwwBiFUX/SgfcWjafoWc4cyfBeHXivLODp/If1eSe
HHaYie/eVtPwdWplkqTujWWMlcT6mlOTF+JNrBiYxbe+jAKOTyCeXUBJHwlAuQsa
qsGxLSDCo+D15AWFtxFe9Mytwtj3gcq9WKl3FLkm4TQ=
`protect END_PROTECTED
