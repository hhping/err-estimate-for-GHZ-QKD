`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hoGnUIeNWc/FBJnoEsy+fQrflFPTAHGmgslI8P3+CsQ2vlT9KlNTQW/B8xT99sr7
eQ/ezO9KXExI6sfkqOECfRQPW5TONh8aG7vGs5KkD1sQf4n+kgAHNTLbr4JiB/2/
D0frB+rnBxgV9rbH49x+h29PB0GLJNpX2HpDNh+xgfKb3a9UMU6cuIux94EV0RuT
Ai5X5mtryuf8FfXXmqcncLn6q7RoZ2Yx/y1Oy+uIM2oK6sJoukiT6KW1af55AUAy
c+eWnIQaBv9z7idoNDkpp+n6rSgYV/nB8xsnHdC2hvWzwDoPfii6LxrHZydkSZEV
Voy4Umsvnm6Iy103vHx1n6Sd8MN028dE08TnB1e7My4zAfwYn2X/DDbGjwQ1ivJK
Xic3+U3hPQmdiwkFZyPl26ALn0hdZMcfDRPoViIT70t260OyELRaPwV32Rn66s89
tB7kGz+4RKBiyl2PpOM1/jOuunUpzHGukSaMBP0dn41NiG0jNMuYr/mICBFhSfxx
gHnSU9Zbp1vSFFX3evY2DSvWNXVb4o0mMrIOl2iRwunxnGUuoVfEiEJ6TzJsdMpp
e7j4L2yiCwip6PA1JBHRDevM6Soethmx0NfS8iK7d1PbtyxTnnJ7In8CVbbeBLZu
4jy8Ngw1MQwUAr/+cwgPGOAd19gwrJLT3iV27cV4Gxw6QHuc7EZduW2XehuyH0gd
RsHaszce8ZvSzDi6v+5ljC4H1pQmKThlPDp/l8PzRm79PeGuBgnoHkhDQo3c9OhN
D3+2FIbpKV8hMw9YHxYhJN1/2h0eHpM9SLGHlEX9EjFqVA87dsyvAPrlpStwqt6R
gea6ZvdNTV/jTiETm+sa+cE70yJIcrF1O+FUET0wkC0Q3TdkkVXVjgTEyufAkeZq
qKutlvOqnM5N5/0flhiOCGg5k0QDPkka9fh+wBJDIds0cd6br8xiJ2Y/fIxOWi0f
UbzdQerP7Z1ToCpS8rPulhS3/c7RMn+3YWD/t3BWmgD4lhlgDw8ilqZH5Vhs/FLy
vWEnTtlm7yBPnIX2S/W0dN6RwLR5yIuMcHZvF3hJ5CwPj3b39ZkTXv88/r0eDWN6
hcv+UrNcTqUQrfVwz0gBIlOq81VcoRJUfTPAYSK6GUO+pIXUNh2cmTv7UBj0cUaI
YhBoCC2yE62noVixqtx+SwNbwPY3hPcqQM1WG7sfS9dzt1xpHQiS8N69q7HuAz2B
nl6zPMKcEkNrqwXtzPfCYzISge4HTSJuY1H8cfRd0G3JzMQ1RlHUjUFlYMwZP+sx
U/GDh2pJeJhxTHO21B6Lz+pr3GLXkCtaESPDBwQIMeEpq7uP3Mu8rxHH/pq/ih3x
8oKFbWZF8w0TeMCSZqNLMNZPCXA1w65pADRPiYqEi1Oq70tFFDqHzV2zBjmtx3D0
eidWtuaVH8C+XrrzH5Wsj6fdoIwkWelVp59mwGTNHYc0nBbkpaMdrCHcHiS33tWc
+ZHGKkM6JoUtKgBYkc1uVsGCX5W0EV1eCiA2FRuoi4mSlcdLvitMrudaqC+wJY4A
FQy9USR7R6McXRjEnj50dODO4p2HpBpzZUg8L7o+s8rI9FxCbrgrqFDhEb9SNcQw
e2ov3+NiwvDe/ClSbOO+rkN9NRKfX/WgY3p9KyrNaOaN4uZ+hCI8P8bs4JsCcFwd
exAubcv4PSNbAeEJOg0al4ybrZc6vAva854SYoIvxlSJRx0G/G45qlh6akHTVf7N
nJC4it7GqtaN+X6g/49oPEa/0kLfYncejUMZuwCzBtI/QSygLLXeqgTSvhJnPTo7
b61qXIzAEgAjYq5wP8bJztk6nd/G4wnNAL0Sdtn/i9gyrCc6+P/YjsfLLueYalLq
PZFMKvPILqHBt0/mKt6HD4/AFJ/TuxTppG1UbDNyrBAuP92RFpjXijyaIb033tFD
KbYsz9is7LxaqJDvWqpBBKO4lSGD6IPgVsjiLPjEkeu6X5xpvXkTB8vWJt3QBPas
kLdHCKTeRn4Ozw2p2hoQagM1qQ9QZ6xqLY9g8RKVWM7/EMGecmA+92XBVSYDpZf+
t7guN3QxBZ2WhWfsWOiZGm5Av1uDhZyzWqBA+A5t5HDSZmnUKMTJ+SFq2osiBBZ6
bcWdNGoD59PxtsPH5gS9M+uT63d2q7V3z+FGs5gTnKsv/b8W/H/Rig1CYsyTGwij
YCsnK+1mP5HLgpyFrpGoQTMfnLYo4LWS9Czx2R217E1wII8OBLoYlntdtAcT0k9A
e6hN1/D2Obi4MGV39QgcnJYmWeV5Cp1JNmSV14CWwJVCX4tYszdNtw///WOA0Z+V
s04VK3lEbheDGkcVfntNUFhGq/gGCMHOf0sxwlae0h/3gVVsnFcVYCiVmBnebMlf
CjZp9CDCeBsWS1z+dit0/dqDYXtgOekvQts06cE5LJ8tsrCYMw2uU++LxW3+6iD5
0w4NI5o9aSrcINZXIZ8xq3NjMYpGadiMyWF5uygLuHDVHrAXVoTkenMv2pqegmsm
i1ypHSlrDhihKaaVx7ckAC9yWGt3hb73gg4Wiifjrgca1v3M6dvFWsqUozOa6MeO
64SFxi7QTRayc7NnP2Qv8TPkTizNaaPXCwWaOBErt5tO4Qt5rwPg/94lJcpNWxSE
lDMvmDKp4Avm2xYzByp0iu4+knvg6406tJucZn82l5W67NxEgKb8PLeHes4hd3kU
nzeWMP69zxSJidtqtk1ji+CF2ln4JVZbp4kUdLOlGPP5gY+A3La/GYcNimF3YD6A
IKSp1EQ90NN2ohWCqPJmSWgE5suf7/iDibC9btXn9oR/giKXtQIpL5d7nnV+Nvf6
NmfroWqvMFJSd/lttaI3WmPlWmv3XXhfBukSQoSQnTeBR7nZbH1RQ3ivGdkkkg4R
wgD5vrGl0wSg0hwakfE8juFYaLOzhg6Hlv9b1zdRVKGHn2Jk1jk3nQrc6VnYyJl+
QZM+i1Gigec6KrGL0qC2yyyiXej8gzsq0hQVf9UYXTRHuCq/sIT5AZX7jhLZZ6Tm
ftEhZbYRW+uTnKfQArLP3kiRRIlau9YFGhO2LwlbkgJ+p9yw6hvRetCitsNPhYWM
X30VrGNJxP2YH6lFJ5kR/gRqF10gtKPWUYY8vF2Wg9C9NJjOU9TZjQeebt2nmMR5
`protect END_PROTECTED
