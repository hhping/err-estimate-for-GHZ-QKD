`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pWVseuV9vVJS6/tfVY3+aXLPWTGwl6yF8h5ydNvcKboEARirOT6eVeDiDoR1t3k5
ag7NIyogn3XHz65xDSdJH43kessjPvROCAnvS2l0nZ8Wog7q5jLAWEkJ5daeaO2C
kvJ/vGY/CxWQo1p6P1AuZju5ROuRLCZeM7+OAyRhUtPSDa6qfaRAV8tmUSwUYQFz
MMWAwZ2DNeBwyDqCsaMnuBd+ZD/31txowYlFDukmRu7Uk3hPiTS1oXVDaPJ8TF9l
0WY4MUvCUo1cUF5IUbiWOjtAZaqM8muGaaKCUK0+hPrVBMrW/VUf+DvqD8IOo+W6
mTARwuPeLYm8Yc02AbI0ms0oU4k6QIfIAlCWNc3Jxc6bR9JU2u2Fb5mPIFVLZCfh
IW9i+W7VOsHNYO5bTi/FuEfl8cIF36o+azygqID9PUExQ3i1TmkdZR6J3Ef5lXm3
PUJ+RcWV6kB24LcvPhUXRLCE4LJ4g1jWdoLur8ZH6Vtv64WC6Hn0jWUopcvmcDfC
kIN9qG/g8Qco/bA7rWHAPDir+shXTE14rxJy6e8+zzYNqxim6ELiqvwr6j/Uw92V
htesQ76izJibdFUhdST3htm+Ppe3joBn9H58L/R+w4gnsZZDjE829WoNEs9y/g5n
o2yWmQEP0UNT7pXPzGDrOycQ38fE/BP/HNPrCq2+J5cfXFGhaKNMH9wxcyExWG+Y
soigII9jA8zJX+ssdiWBeFveutI3BF6tpi3woY/yRtbUgLprXTvshKTGyETkE3vY
TN7Q/ZIIGBHOyKL0mr/tLfeIf2TxJcX1dKgoXRyYbJwj/LgwkXPdNr6S6uU6jsHI
ZC0sWd/2PzBPUrCBnU/UHN398JYnIWizKW2Oa/K8mUobkI4eiXAwEosif08Xfmc4
cJvORKmIF+c2w+x6BITb4ViI2dPkrwN25uUkTqCEQEy8cZ8XlyutkpkClQeIrzep
hi0XFXeMqmM9YDkNpV1lgWxl0QP/fkmsH5Hkpd4AYKxxl5zMOqJHjwkvkd4yQJae
UpWeiqsJKwSlzEyCdCVhIhBo+PE3fhXf0lfr11MlwisvygX7sdXTgsDsKr0tzfq3
gM6vWHPDUnk9DXA2WCJMJRPrmBghD/UAF7fPMpLtGRK6+r0rp+wkI/XAKJo9ew2+
DY/KNmBb6nqgKlF4159WmG3LH2xKvN+9lKteerZX9hMmJkJKleuVEFhzrxgIzWN6
f27nl7r8YyNRmajvIPLKs2MyAVbuScfr1vj+AKwnJllsXcDAOILInZiqAY9CUNMK
+iK9wQ6CEWR29MnlrolyRcQ3b4uFwVuxG88yiZYuPqSdXtrTI42Q7589yC31D5oN
6IbssLtL6xGDCOhJJNt0DFGtfzQvhbQNCyZN4apk+CcqtJBqsDfdcTg7eM0ScYoF
bWi6RHK6AQfsgrqDDG8HBNTOo8CDfrJasqQbd7HsFI4ceuqgB/wRyErEWbDGa32w
Y/R668wQk4TeVouhiOp7vNIAzMnCcVP1HdJYBZ8G+l5DLgncTC9JDONKiM2Bu2C3
rTmuYb7XoYA4FXleLYKmt6FVRzTZgdYv0JMxc26JeZ+ZXTNuLCTy0Zk29B7NvY+N
WfCYM2mmrDPuB30mTm8L5ihYx9ynkhgvWX8Y8NKK/fXpAJ2cl4FqAHfnvtEcIsZz
05Q/OgWkiX7m1gwTOeVxdYVix5EgBbCbK57ajwavYLOaM46kjqB+aTH9kX4RGfXm
NmGU7f+jX6G+5W7vU7UMvZY4VEYhvIcqzTvZe8hGM6H1cD64I8lvrdrFk5sr57rF
4uLyk6KOT+YI3GqLHrxVSkFYbizo8X5VmitL+FotVbYUA/a2K9kxI5yiKrzZL9Hz
RmXYuOLwrmQri6S16K+wXeYczGbadW7HHU+I69klAlCURY5HVXf88t6Cp0o7ed6m
fHaZjf5dSFnT0XIIPXkPyYkfXxvlO9pLhz1WOUFTdGjnujL3LtKgEN7k+fEJ457c
Iv7aszQMFV3AvNDPlr/Q+mGeyFdGJZREUAyT4apBBSE3yFSHJFhWuBlpRNCGVhru
naYzgF9+Ho/y8uSyNpgoJkeMHaGHZWQw+5+wzh8/1DkpXHRxA18ecJeGVfWIf3sr
ezwI+qxFLjEOBJPWBZ4UqusYgAeMy6wm3dLZX3+HlKIJNIRBsr33cRv7yl0US46K
GVl7Xn1a1dOH4a4fb0TqJ8lM/7Ns6C4JuerwrPC3nHsP1aGVsoHcpnUp35VgydmT
1CyLb8GtHiA0N7knrFtPlygor7bQtfAx02AYw9E00MwXT7lL7LIeuqFNZfxSszyG
D6jOx46bZMNrt8gi8oJ/lJR+Bqh4jqclKkHyvyQMSTYex6F0VmKrtWL6EobCKkHZ
BLy3vsIGc5PFeguX7oZGqJ9oQe/LQ5gtU7g3IoJx+lQrxIkwKXNLywBjI8f8wRme
Gy4XLtHALQ8ykuaS5fQaVh7aVD0pvLmwCMglBkpgwG1yawgIctiLupjOeoA9lnSH
MNUMP5dpkSZJbFsRE6b5iMn0loFN0d1Ic+ybygo91Es=
`protect END_PROTECTED
