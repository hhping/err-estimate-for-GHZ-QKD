`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R6YNgNHLmN70J6pzLjdy6aoj/Vi2jAjWhOiSkxjERtyzOwulM6LY65gxwRvW0h2G
4QnDkT0+UXz32Osm+Kp1pxgGsnSM4Wu74lrg/1ID2JMRNlKtxP7th71PEAvHBuDm
Vx6vO5hhxykEtVC2khrXD6fNIgog/1sCCK8ueQl1E6l5iOM5Sv4TC2g6UGzCvLpu
oFZ31b8UVe9x8HCYGVXMIK/CnEgY3mfGI1XTZg1ok3osSaWhsiYyTTS0sCrJMdfn
dBlfniq1htNsVagkMdIleDRxJyB3O2xFKKciFXBxaYja7uHaV4lhphwcQe2FxXw1
HTry3uIT1L7N4cFXoOajmj+/L/nmrxblL3mRQhGXADiPKUVPK066hSPbJLFR3DZo
yHOB4uSXAKos22KsPKlideexUI+6xZykZFi6OqyrbWrLL7nTxxDJs6HhnkQKMn6l
piBPVxOfJnXrK3quz/TDfMKOSeM0kJyXgam/vYFO39IlTnJfpXnqbYKfdtTevNO0
yelkh1gxQDR35VqO4Kp34SSs5k0YGptiRzv+UbIFQaK+K82UHx2ASFe2yIl2GPpz
BvqQR4KunJ0ObmD4Uw9OoZeeaFu3i1JCTSw2dEZOgbLChKmiOc2A2UFe1hCE4JIs
uccStyAP1TZjJJMCC/X/eB4/jm8PzKuEnVs/82xYvPbzJe/qhKTIKMJRH4VFAqGR
xCHc8ziGMCfNsfrzX4U4grCR3HL/2t9o1y4/HayQO1TIxrmzE0WhkveILBMwKl7b
scDyC7t0q7ZRWBaYgqfSKBequDqZ0QOvCzz8mH3JVZlIDXBO0B+oQjZ6KQtWrV7a
3z4dQMlOIzjoVzzj3nbmjMskwln0eBEGsLlr1TJ/GFWxNy2G7W5NyN/tXA1dqEty
fhXQfLimYGFaGusfpBpF8JA46/5a8WGEWg1Z3rvFGKEwhwn7a8wxDLxD+ooJut7a
Mh4J6SEzaNBuI+ztIliPGS/F6CcnJtuHrw/TqO8eFIZh0ok/9URhp+LsnEt88ot1
Z5Y8evPT+crqNIpZjTg8WnKTzaiv4vKW2I/3z2VFTpdL2WqR7t0ZqXXyor3hBBf1
3GduiR2LuODstlNyo+nWRW++rkAqOeCJVacj6lFZrXRy4HQGVbRmH7quoLZwPpfW
kaMCqNewV400EeiX7g1DhkAWcHzT5cJ8tptx9F6EYj1LmlrxK1ZRfzI72X2drQcg
Cg8aNp4ani9WK/+vl8EZlG/ESDNexOMlXKiuE7lwzkMD08558z3xeAqekECdHlS1
g9oOXNxKlZ9m/mwVIItU8tuZECFEKanq3W9VbHgQCJ27WLlDdDrjAI36jf0v1gIW
iZDmVOizNVXd2pDjaoNuy/PF6SPHqXQFL19Q5YGU90/wc/EP95pLpvzJxKF8O5Mu
NdtE1yruoTt7o5BStPnxIF+wFVNKInA7q8ElBN9zEow9+0Ec0dXHxIPldhWz5daD
m6xBm9y5ZoQez2PlXQyjH3KNSdyfHGiJWOx1rVQ+RL+OyTg5tFXaadwfIle9HEFR
IXS+62TK8sXM7nax0wxzSEHO1R4Xt2A55+hSAm7fRC0=
`protect END_PROTECTED
