`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/smSB0s1PYBsfUv9VuFoUaUOpvzS4sPjRvvtnGW2wI4T8t4Lj9vsw1JBYjayNpFS
S72wz0Man/mGsIOWWtdc9jKSa/4x4qifLwjAcbS9t1Wi0Ca0nSzM3MLgFuC7ULM5
PLczsK6D+cwHmwYouEgkxnVIj5xMV0Aff2x4T4FjnbG7yDfjZDyJN8p1U0Ozt9bJ
STEVCuCw7x+X9/gpCRRlMpf4tYFFp4Ja/J2NGZ26YsWQkZcl7thAYeggWOqw2wUw
9bxvCyhXqGna3k47yAqLQJRtFbDyrUEi3CibO1cSHHqgDrFvYPWbw0z2C0Et8fD8
EtOQnLfYLv1i4LcajmO42HeqDKzOc60QPHhlidFloQkjkELuKte131igze1Ao/1I
m+vR/5m9MPXuwXTSo9MrrOY6Bvd9qmQMm8/Z3LgHDXFzR8Z0XX4OM1/LZYg8Rba7
E8f0zBOr0u5UR5/6gbCM9+z7+dRktCj2tjMwecNjVQ5zCZCMpeLuUJD/54C+9VWM
H9fTdzndGJtAkFpq4IGlYCzhQaAZxA6zeDN6qjc+Rw9hnEezQzLoxcSJEFVEXGLG
bRyapuSxMWLVnKMeWdbB2g==
`protect END_PROTECTED
