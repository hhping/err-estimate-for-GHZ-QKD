`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Eya4UXIvr0hVsCqGvi/ajNlejm+kWjunAS5+ecUMrGCo5cO/id4ohuPcFoWqEoYM
OevXzMPWOPtdGh7ucdXs43pWl4Y6gQJVr5SCKt7+wkFXu+Pnff7XxeEMGdQZyIdn
Czkq5XOxg+DPbrH3j8/NPOLQ2nWvIOd5KdgkBxB8IRO2cdpJkcn7HAHGB3wk09+n
NAohnYDGOqKsHuMrDgZVaMmAhyrkYzsr1NMCCwh5UNGKQCR3lqpdwD7rKSeKRoK7
P3L63chlMy/qNsNisnySjxcmxmIRRPtD2J+cBppnQcTgQQYvPJ4gX9eSC/GLkmeR
9eNIU/4td/ie5kHD1kUBH2WQdlcJxBtDbRSR+w96OvqZmi7E4jicYxWSp78/rLwI
LFLLtIrIWX8zr1WBwowkgZWnYtda45jxW9Ivq7bs0HYr1O317hX+o7/OISaQEQX2
k8b8Wn52beDJa1GztSNbvUiTmeFK81puc0Biv6bBYC7ATWCardPLY+oViudMsikh
yg5s/GzuVY41fTole+IDOi2jyWbYpyIXOgZmnQpl1OryIZFwUj09OPFMx1UsSef0
j1H3KVOoRNXG1TLrS6dF0xW3k/QMrzYgjuwzHJv3HeDOzJh0/oudBJmThZLJ5Xqx
aGOrn5uHRNhUdMQnexme7a7Hv76PDQd+qXWKa0coKVUwHkJ3Zk1WtW4TW6X/mwC9
`protect END_PROTECTED
