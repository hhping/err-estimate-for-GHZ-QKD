`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HuK1LoX9qRlnGYhcu/BN/qOpuQoJS0ZFiym/Wn0VI45CQfp+v71FYfrKFrB3dL3/
LzGGzpe/NyWA+hzaMGiilR8//cGeUdSPOJbq6yRy92sevo4N6Y6mVP0OWDkOitsx
SOaGw+x9bf45fFq7k17fZTWOXwdMYGyKXQsAiMIc0os90SIwo1N0M5NTP1n5EAbU
s5Tr3unnYN7yTaZrQEYd6VjVetocmwy5G/c2+bng4+q7DGqn15ceSvvkCrN13aKF
1OzVcLnhn5k5JdOHR5Qm0cPy10yORGMscg8sa4V7zlZIG0G5j4yGokdrpbaRep1z
tDHSObBtxBvpFDSlnCg5dX0iyP6BB2puJid9NGLYUtP0aNSlqMaZOMOvdNUgvRe5
B9ueOwaLt4+8kfCkmCogUvE6HhdQRoqPXLfqv6WPlQqoSMJn+7hsRMtYvDmQBQOU
VabFRbErXb0N/Dcb9Whs2Wx2mnd+ubMCh0c/WWFJn1kXbttaaeDNKcFPHceC0MAl
ujH517tUIdHXosQWW7oPapcsZRPKoqyABPn738yBnAPZpG8mowceJCmv0DvJ9YfG
J45AUK1h+8mP1lTqrCBYiul+P9bEGjHsLrT6AfvVjWa6s5rApEM2wN7/yIk9c13e
w/9IUk+5pvj0yGxF1MfNIdjrPzFdaF1LT+Fy/0p97VUKHllOmJ9EqEPgx7JNNv9o
5mNaYa1T8CXOIfrO/0NNhYARBFcYyhYZ384IY64xzDh8SF6NYtBi7spWP9WzmpxZ
arpDuzA25oLvolDrpJxg8qY4QfgyItliMiUupu9kKrw1bfa9stE53/Vd4oHD13EA
IjxU66q+57V7axC3ZysZAOzKA5mfYUIwPsyerH4AMFM6WQMylMa37fz/YaVqyxOj
PdrMHS591mEnq5znW17hh9VI7xtbxlm/GKCh7ULrRWVSHLfjbzgDQTtc9IK/Py1/
1vK7Qh2uoEtP+E0UeFTy+g==
`protect END_PROTECTED
