`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EHS0jvSTJQYwa8ye9bgT8CTdB8tFTR1e1DEC+oN9Kq/ueX84N7VQATa3MCue/0Mw
/N0mHp1UxKFKQ/4+gAmIu/B+Pt9+QAM/HSay6smSBnhhZAY5o6NMp2AznoFa1fud
OuLWN58Kz7rh1YRf0J0GGiuh5cGvwBpT0yiTwLpGudGNrQmPErhPgAXE3LfUWg2q
o/Fc014qbFi7Xrvrbh8tTLoiYCWcGDbNZVEOCW0GiRLGgeqK3yH3KhS1Emh8UUqo
/Rc6TJPfDQagKwlYYRKru2f4nmbLXp5+J/4OsCwuklp4CyDj/QToKWC5MR533XpN
Z57GOY9CtzIK5XXkgm4nfd+yhMdVbou6VEouECIyPgO0msBWhVOJeiO0p84n89Wa
6ufL5QFoyXZ4cWXGsltTDHLG1sYKebSij1L0fUxwhzc44BhEexVZYgysYLUkCGte
CvAjpg/qEOhdy4dRu3Uv+knmyeqRwfCV38+L4CaGlP0++geURDkpb0U2O4yp2PlV
vMIg94fBDcdb/AHy2JTfWAfRkEqqKYwUxsEtN8TjKYSvVbsfyQuiPsf8bbfiCX2W
/tYO9fP8pe2Wva7y2JgzmNKtuobSphhNpZM2M/ckwi09obK+/pQozN0o5lIabBXq
iXJxC9wcQur4zF1p/DhSOQ==
`protect END_PROTECTED
