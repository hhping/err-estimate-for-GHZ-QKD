`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V9oe5MxsA+1IVuGXY0jd6ysIqLvvMRHdoJ2fKi0KL5DGRJMYZjY8Y89EywQFFv+d
UsEdnfp7DkoEZDJWWRHxdNv29rOsWsIBVlLN2pYL+wBcSJRWtJpkXMAo1sDcTDuR
4/Px+LGUf+2bH+upQsateIjhdba1SZf3Cl9lPTCYUteQuEOHtgdL0B5OFeJyChMS
QeMxQOvMeI+F/kep6s87CKcodZa8DCmzkwastt2y3yx/ws3c5JBvka5s/tIW5W5Q
/rBDaTiND1cic/HrWPfA6Lsz0bXO6yRskXcqJVgPcsz0MvClYhW3AssKpC8zGyz6
Shmi9nNB4oqOSsFnC7/S4gIXvvXtNIodWfL9kXEPZHul21RQcDIj7VTUCabRcdVw
Pdi8XaNi6FjGEcG65PY8v6ypCLa2mMK7N6Hu08VNzRe8fzSkX+T1/MpKVwkvldMm
+UEDsYsaL2+r4qdeDDJfqw==
`protect END_PROTECTED
