`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aEX4bHH4mnWfU5TvZgT4dKtpwB78R43mKFIs7ub76SRDz8K0lJu5BqaWK6maHAsl
eGOzv9R8RD1roGwbrRhNg+gszGUD9U9MDi6Gzp6owxG3fB5DoUxn3YfBGHC+Fcb6
T75xVr5kGvNfWUVFQmDq8p+9iIpnBEB3YSl2hfzmy7DAZCAd9W4QuD9mWEldG7XT
5TGukPv4nXOVHAnybBYdKxbQNk5F2hy3OxUBxUsmkb7CxVzr/ec6CN9JK7X+wo2L
DizA1GfgSzS7kX05+KG4YGwhUgr/yUMy7EpFaThbj9IrKu1FQQi/4hBX4kUv4iCy
KWQP5LAr7RLaYf2uPcdHnvHHDKpI7sSqg7lTzK4J1KB2/5ZFUeMt1hqckYSEJixf
ccHJ7LeAd+TRJFbIwM6FC3M2ID0nf07NcVFYJeHzDQ5HQ+UrOo76jCaAcIWzaOZv
a33lzJQSsDXl3GHao3uXalnTD6g9/kUjHSmlwwXSVJzbpPi2K3iCsm4m33e2kv1R
GYksQyuBMfxX1GkASmFB36uLtl+jogPtMeTpQ7CGlnqkCnPL/2PSjj2OEhAMTQAz
+aKJDMsrqxn6E8NCvsruNSN5tia3L2vtKEEMXIYR8gN7Sxqnx26wAc2ixyBlhwO6
zxmFczaY0JOFgss3cQ/Y27MHLjAUCZZZC1kzcJ+V6fVLHiHo/AFyJIlv6ejs3eAg
weNMQcCuEHwud0xrD8m8hm02ok5lrl2RY6epuv25wSQ7hRMe2jGLhtZF0+2DooJh
T/eWnpoKygmSFLzdiJW/BvJxAs2lbRBD/8H8fkd9VmcZ4zvZNpEk+df+gPPHAsNj
j8GHpZna4ou4Pr2elLLipTAOgal8sVHHPDMobgH4diquxx4YsZaonECVnu/uZbGH
7FT+I1nQhhY8xT+TH0PHRHTPcAg0goCLtWSTMHBywzi/+jFfCkBgQXEa3ruGu3DJ
DKiXzeGtru4tOVaDNypwUni+TVz6C0QdprBO1qMDoKKHyIqkbSHoLnU7e0zzPcNS
a0TXvhsG6EXMIdphOJ7qDsjBiYP3oose+qBiZid/ln0jbEsqgcbg9nUXV1qodAhk
cW1WAexqUfIcEP9wNuJ3OapPv7Psg3Z9rgZjA+Yv1HF0WCSH3eXXKjI9x5TM/kTm
772NsTQ+cGQB7IAQB/Pd9dmHiVeUZhA/oIsHLSxhN/vtaRWCGSYDkD9M2+w3hzSC
0s+h1bxbLWztxI8YQTb33tvlEkg9pMg79VJ5T6dmNuYFkcnhz7Z06Z3SXD4w5/PX
DeIRfGibkp6QvX0ck8OK7saf+XKr+RU4X6TCYEGttqqPhAZ/x4918M+TGv7SgJw7
lLgBmc+MFIkErQEncPgcCq17jdP79cyR6lXKwzp7UD3A/040gmox+ILXNIZR/mlE
96WMoDFQ7URUXSERn6GHCTl1l6HAiD9/lsubyDwopMbGig4d0BeiktxHVSPOs+nv
Vrfg3za/XhfrEmF9OcarqeSELXeH0kMHO4fG8U2/IG3CR5m0JRckJAKVwtqvjx5K
m1Qr+AlPPr/g1Aqewe4yDy9d3y9lwflK1nkUuKPcAdMBKsG+5+jH5m3HbB2AHEmk
GRabEC5judzzc76rNw93HCigytJsge/tj2Ty3gKGk8Hg08RV+BJ/c1dPOIIyK4bB
D3zjZiRn6miMnEePlvU/tjYvcs1bHWfdDo/ybfiWI51/NxGJOndnu+u81LhCdf+L
xFsIqaS/P3tw4er/1X64a88jWnNHy9EIf7d2Q7Uhp1CgrA01X9/A5o5DSShql41D
UGjlkMQKUl8bEP10pt5aNbBJLj/FKirnddbsejxVoEEJIulcb7KWGpj/DoBNV7va
0C/E4dE74tM2kIO2f/j24G9uiSSsMFgWSLDvxHQxiP5fqT2rY6MGJjySR8hVln/I
4kU1pmzRvX/4GTRzrxtSCTmfF81At1TfGI+9/UD1EMSiG7/Z0PN9eA3DEBf7uRHh
wVzQob5++AHGGsMvDL2ljIAONxDg20uPISbxjokRPMrc1sqn2oOdHQ8+fZmAQSUq
kqqtsb9gq/wQhhBd7uyDD2Ts+tFzwSDBuoA0nYQ4AUPNT5k48gkiP3UElgK2UBPG
mlWcw1M27u6TT8dY4slt+PNoRldpSQM+zbtuE/XHB9m7fcmu0lgLcTscsku8h1NY
eviu1GRQT+nBvPhpnJEHFxuFawBApGlJOsdJewc6nuOcXwCZ5YIpbv4lyeUbLDpz
7We7Z7ockZ6xv9hEobfTWYlyzcH46JX2qkIhl77LqzfbZ4Y6Iy8UOi9bo88dct9F
G98uPDIvZ6DisSsARJ1bHXOTHFObeWYpA5gpegFLavokWLheAKQx9/ZIIRlru3aY
kUOaO5VkilkUJkDDDDTFEqs1TU5FdlanR5h4BAM6DdrcaPiwIyAX2XhM6+DbENUS
SBNfxlItZ2sP62C20Ht4Blvfpc5CCoaZdsE7yyqB/KeONAbl5WWlnGJwkmwFeV+k
W12ajbWdbt5WfiWNGbaDvw==
`protect END_PROTECTED
