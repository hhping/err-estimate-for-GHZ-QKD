`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dz83umiT3eekTCI6brIZbtfu/OomeT5CM+/DLyiRtpIbrK4MimfTYuG/oLTRrjBh
VHcXeICbkY/dQhJSkYtR3yV9Lcajncbn3zMKRUt62HLyU4EOOI5yK9E6TQrTLkeQ
5mNNW6faCeq4XGhKzkjdj5L4Pkj50MwpVCPT84HdZ7H3ZLrA1lxeTj8ETwNIlrO2
ZS0HXMco56acykXyACNZaBrVSSDFY36FAd65v9g3TD3zntiVTbwdqaZhTHq9EKyv
AThWrr/LU+tFPgB89x83ONfGbhzvUnrKmAupQngILqPQXH8PnswTvY8NkTekTRJ3
LKf/U39hjskir58BfXZ92a1F46R5pNEPB8kBibIo1FtAGwpTpK0F/8PBGV6bZmwQ
8T0XGpDV0BWvU83unzQx/HQ00ueYgntFtJDImtuHLjVt++zX8TRpmRhlEIOLReXi
9/+hIyBuPWW8ji+KtqI05Bfhc6zOnb0ku3ONo8yRp5keMYZyZ0LfO+ZCNCdPK4lm
j3ihXATWgcG7c5Y8uBY1U+90ij/WLwnFmseNaqu4QCeijO5X7Zg2kWxuv+2z9Owj
vdJDRwkwpi5z4+YwIzYinvnpPqZBPRWNaA4inowVrzEspXKEEbGd3zQjpFKoUHZm
7QZ8xRAXO7WAdvB8n2gEk8C8GdDS1wZEOc8IUMJaB2DHBQlXLTlqSCXK7vEH2aUi
WgZK6I2dMvuNVZvaEDsvr7bo01Y7fYQ2VtSfbEmtON9+Fx6DRDwIJZt4nX9LvM2U
cDgTiHO9hwdliqZcb/DJ270zi8RsnIWxJo23E/VB0t0JmKLjANrlQB1WiWymcGgT
QOA839RR4pPh8eQJi8MB+zIQ3Cpf0Sf2w+7LF6nRS25k3xNeXU3DXAEIffOBGNre
K4s7vMS0EKC/5SCu8AY2bMS7nkqGomHf5EUej2hc2hnutlVoSObCL4zY/UW0jc/K
0urxn/9xIBOEYpAiffjdtxjApnbcNh7I3xiOeAyt3mEJvR0BB4o6+q3hGNdxPUsl
WJR9gNMXBJbARbbEgtRPM3Sicv+y769WihuR3R9D4lngtY7/y/ZuEL9YceE5fChy
Hm4M0nNwenD1vocFUEquBQa7pVsiCP3qa3zQkMYONFjRuRRX4hcaDHduX0Fz4GTf
anfewUSOhYH+8yFs0E/aG7+whDnryuYbLkMY0KDyK048Jas0v8D6GHCSABGElfd6
SudTOODmB/2bbnclWubxpYPjmmOKVEKj12OxWd0s2IDN2/l2gpG5fwu4Y0H48nIZ
0LLjH4PaXX8pM8vY9cc4j3fpKwJ2GM4Ks/8IGA9GNua99YOUV5t/sNkFchWxCbOF
Y99Mx3in7CJGQwKkcchFoX9c8PAH6TIrzPdeWvcbq1QkIWRfBbMyQDUwQPr35RU/
VsqOrsvhWNdeAY4JFJzFK8b3jGTxfncSX0rGfDvRf+6R6uayLroKTBlrt/QcV0Pz
+JrwIlPzcxy0eUN339rJpd3amQDbuUDs9BV3WWKHVFpucR0n34tmNzgfPHg0jo2p
03XbroHPFCDZvEVu//4vFOLWL17yy3gTTR9rQFwHMbfa470MAPcCLxQXdpCWjjC4
ObhIw/Jn3KV6Jg3FV2hLvIZo0UkrKuX4LRGAsuiefCXjEtMc9J7gdbLnTOqsJ0kd
azOEuzVg2UeDM8uWR2CgE6KYyikElt85X3qioqXAH95S4Cl6sZHLmktOAZq9obRT
mox2v3/driWy0lZCcu9o6z3+2jooZqANs2jRXDUWRUjWJ3l9C0cxB15wOS2vNB79
`protect END_PROTECTED
