`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZjDkzaM8PPtLTrEp/DamWAOkz2KH1z8bG0erkuFPDsRTntlt55z8jZKdSMp7Fc3O
T1uc1Y1z1Ta1fRGPs5JflpiKFFlnCEq/T7LRJ0txuTuld1QLiQuNpKoLvp5Hyfqs
ALEPjiHBjtP2ywA6o3fBLSvsNqd3ONyzhe6eMnuYLXmtntpuhjsgugxgTRo90oQf
pIreQQi/NT4qnW8cDlbtK8HfTWnaDIYSkiGiJ1OQD042DqDQ+HI/WxMOTocTPyFt
I0XNz2OPHWFq4G3fd9sPW9Qh2GCGHtf8j83fUzhZgFZl9Y+XnUvj0E5zsugOOurb
EadqR1M6vu5dlGEAhczv9IxqRQiKe0Bj5NnSiZKokhErls9pHbPy7KasJo5Ook+d
se9IdzS9f3vIR3XcQe29ekpfCmDgD1Ot2l9guziC/gPMlbJwhK+6aSyqZSZWdixZ
TWzZbfRRos6UPnoaYtUwwee6rLH199OMHxhwGhvJJIIBOwPKzsWJdIBWTGtEt+El
ak1LozUJfFZBX6/YGjaGoxX7e+vDV7tngNgHudjWKX7UK9cqUWSmH4HaQ0RIykx5
ZNtDxZVCQiaLLGqPMqhXfNucYtTxvP+FuYsQLu8JkDvjjvdBSvBnA+uldWm3RfrJ
ehE6K3Cq8KKxqz60x1sZgDMtPFaZu6zHk0GB1kmDNVJPImA/BxHBq57fEvpOISB2
KsQCtS8Jt256M6Nazzuysj9i8W2FB9uV72MsEYLACmSp/k4m5qJKiqwvSJ4F0Yaw
EHWO97Cj0t8DkC66H+UdaUtVzqu9yJIdkbZG7I+JQErU0jK4cwlyd2iwBzYSr4Rw
sfZv5Ea8hyV67/jh0INlJnGqbsicJzREUpxWAYbJ0ps92AEDiCBKtadtw6LdtrrB
2TiyYAR1XhpbBoippyhA2k279Oxzzna2kQaNnlTeWFssxYEzU0Qh7/rLYYk7tk1x
T65aOnInJFoXBqVFsJwFD8Tfs1laHDSwXOuz65+0b/yqB68AFK8g4WGaHLpRfquy
VH0sg0mKRcNV3a9badiss7CUZYd9OVqx+DxwwNda+xNIFly9xnnrMXAOPyyi3ZSs
d4tTN6YhHWRbz8lwqayjpkVkrpql4ljN7lMkcgftthLyvdQA7wlz4moW9P7vXM54
lZQie2ufCNrVRyejyoD+xOZbkSZrNgZERsX3USD2MThmJ06QVXx4KaS7OONygl42
eXbFIEqe8d1B2LkBaFu0rMiO6DHNUocqwWlj9e6aU5zfrtyqj0Mj8CgcM+xPjmFY
3PYVwl+9ibBkLgTb2fmHYaz7dniKe4rZWRMPmCP6zT5Ge12BVdR7i+3JsAEJSIcm
IekrUDqU9e7YydChGgOoqzbiBk6pflI2D5nGoMTnRwpvXMd/dHYqTaZ3ogk7m2Qm
SPDAEF7oaviIRIwTSk0nr07s3cNplx2h4V/vGsVBjRayXZkN2OtpS2u0YKS/f+Hs
NmN7WKBezKgO9EcMQurbN5uhrF8IiwhQOiAbZrSwyJ/tpOS47NKIeLosRNpsq0pd
iL7OtKJIY67l6kWeFpoN6Nkej4D+5lYYxL7yr5DtEZ6Oj8nwS+DDiM7b4z7xCQAO
fg+3ekC4WpzePIVGM4EhXLTo+bdDa7WwlgUcKhYVV4oEYqo0DBrJYPEXg1CdkvSr
bskdRWibD1TKVCn4Ji3m/rex9paM1Rc8FnJK4rAiBwR0flKSDJOL36sZFrzKoxLA
Cx6t03IvjzClniPTK/XxOBNuEgJ77PtWCEFvvttvyLBirPHc4Dy6JriaU8SifC54
ujndQ5sCW1qiyDAdGJ9N+b9wpDbjFQfP3YDY+TIofm6IFaVxV+/ttOJ8VDkWZGFV
IHJsd+3QFLtNtPMKNEXritKsoeP6lDgPkbkKJcPki7E9JjknToe6O+2wUGiDrJBY
nUWitxU9crpMcRQyIrHvaTdzLisovHHfA0jqAraZ3b7ITeFCueeTd0yprJ2XnWMH
7Gmt9Nsqp1wOIe5qaJ04DFu+9XBwOj3QsnObFvcVQdcPdTp6gtz/gileqQEaLhDK
j5whV7QdD8WS3l2j7S0cm9EH8x4IJa9tOqLLR2OOC40GMgZLT7jVXxSnfHsqdeBG
+Dlu/ehawFD9+jr4TQ3e8dsESq59xR/EOkShnr9COoJKSFUPL6AooClkaJSulAn3
MQBDYBB86k39XBx4adG0/yAp6leUorGUSauGvaRTlfRK+jqwMGtl0wQtNjmWuvJ4
y30KidX4QYnfpWRf8etpf739YyFtrJmSNsAdV96u7902TkFKvRkoXoGy8ZdKnEMi
9snN7tl9q5FVkeXgFzId0cSNKCVeVZqeTwknbShU3HxWu3hM5qVzVyx8zU9LRYH3
7SfkftJNNaOAPV13UoJchVj9X1BVBjjABDVUYwXImih3akW5b99B9I5mmyT9QJcZ
tnNWJYUygpDCmhV2vd7933s8JqXTOoF8rPM3hyEOvOI34m7BQ7TzHU2zmkXNu9mf
5iDMfMfIWshOeFV8afF0NU/efGq/r0O/ky4VUyXnsqMeljD9jt9Uj+ENVASqIBEQ
9whVeARIXqHGKSoGXZOZHlFoUAwiilDeXArl0WYg6/vhOMrM33QBtNXbML4bM2lJ
Hf6p19Y4aFthjKtqcwQX5oBoFuIfpPC8jB+IuZOohr9V3JkbALd8bAsRauyQ70z3
V/sOTqtKLoiEZjp4D27B3ZeL79Vii0G+kvp2QhaPS8tSuKk2XR67rlcW/3ZLul+T
QLd/pxnzkHcoyWaGxDVhyuAppj/+n5GL4ZIHaHDWqEUSchLD3W0TlG3GisQLgrrm
M7+ErQBcmilOyiEhTnjP3Ut3v5z/d/N0KyWayLIqDJxBo56MAkIBLueFWx/5xKZY
C/h1sKwGOrUjiRajcJBhJo/WKwkUo4BZqK1vTspuCijod5dDRzZJ1+91ssv27MYW
+j2Evf6NtYH43Jg0WM8I9r0kz0U9QEehgDUt1l0G8zGrXpwOdgKb6+a9AQjAQFrf
O8AMfH/AXpVybnZ8Qr1aKMSEmr2zkMTwh0mXO0hKNTsvjzd9OxtNbKJ7UPBlgb2h
In5oWqHtBsYMruD4syaqA5kDH/ntvPcoYZtMcyyCIsHWun5MRnGztec5KkviQwj0
iAdOhzYN5WsBWziccJLio3Q0Qom0TdtoG9q1/EQCaaMxXMNj3+BENYR1oSp3L3uk
oWMub2IuL7I89BtRgpJtle1W7RWyFfriZ9c+oB8+Zy1mIQd8tqS/e//X1ZdGOvqX
TBJoN0UwA+J2+Y47pXqR4AY48xV6M/FFYKNBlNbVGMrl1XRe79v3uHod5/Hj11/g
u6zhria7rjZAdZqUQGUiaocYBadrR1MHWZX/Wd3SfmArjHVE8Tj99P/gaewHny5d
LV4hPGwdEto+/LWAE7PlxTxmAVlJTBNEdlg+EbI+L+3+6Cnm4J0uW8RwsU+v9nrt
JvM5UFHFYRMlIIGi0hS08YxDTDRLyQ1ic+jNGDH7ZGGso35fYdWcUHRRksVSkfGH
Ypaceq/8/AG9yIYePV+O6RI4X/ybuTaVmtqungo/eFkGVrlnzcGfGheZ8a+hlHwJ
IwUz8ZeBww6pPTIeOMp7/JS5OLdMdNPY065De5foy9CuU6/6WK+Q0VkF78KpQp01
mkevgDzFoiMD0+A+uO6HjihFWlii9quAeDnUj7KRMUEviFb28mr5B1qsvFX7mLAF
+/wMocrxZnn5x6+RBj+hj71NUzKRflleKJGh50j9IfqU/VcDkJOKtYX94vgL2TUa
74BAsW9bbp8Paq2Hwep7GIk1vyfxnMidtp13tI5egBSqRMAadMtHeBcE+XrHnC2T
KQ4Vb0IES2KLUY8VcfUqwjIWqHyPEEvEQnw83TXnS4fOUYsaM9PBasZ1wKVUIxX6
c3ybjP1gu3wWjOoSvsN9kCTTESomtZvo03SoNeAnAdWMn32n5tmyyt5wAF/tZwa/
`protect END_PROTECTED
