`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6+YAXXc/VpZiKDvs8XFH6+b4Rft5ka0rtLmhEYXN7dVRMy599s0+KgzAS/QC8lW3
2W5E+sr43Cad/vlPoV2a6jnXbCR4Ir2/rxzakIAWajE8+QI9u+KTNghPG8z4xBp5
3UffK0WZBPuueXzI+avBgYiaIYGg8VEkBLUg8I7OpRSZLHVA5tCq/zcyq8tL97Ul
/iLXdlMAnTw88cdmoG35XrpkKUOwP6FHc28EpqpXswAgLEPCSeeOeUo4iPQ+Y3Mi
kktWSCNDJcByp3bMeELyuzlweBbjpdgD/r3xafSKMhXb4l0NOrrlK02EJivOT2YW
F0lFExjWQDZcO+bhYc1lMUEHz6/gi7HjKGqk8EuVdEoPUxKrnA8lqc81+rTREtxH
qQETym0x7YOelkEktOqmKkS5Sx6KAvtXqhVc3l8kU94KZB+IK2vSaBuiufshi6Fr
0T0TePXufi0MZhjMoJ+dJvUQoYuHPYrl/ha8ouwDOGW/s8v3Rz8JZckYzyLOyqL1
A89z4EOqs3c6t9Nb5WtTpk8pAStBPaHN/lkeUk2J3ZamT9d+OhSjGsqrtqwLSalk
4eG5/xOyNUi4Wg+3qQAoT6/AUHv527aFBrBS0hl+8/UxScAS2myQ/QvKJaGSsQM0
fenf+uU3syRiuoh6Ud5/mBXE+8DcupobWg3lEf9mdkSsf3qKyl0tPm/sQD6lep5j
h0qE7MOytFkjINmslDtuMOYVXQGOhTVJI3E4gZ3u4zD2RPQEunHTnhCVARHscoKF
6XzaOLwID7fFvaLtRaw4JKqozI1OhySeEYfda4vaAlamfNSs6lwW4PM7LbT7sVWg
byVWgFewKk50T7bc5ZlObIa7ggzNZS0EUa9eFvO9gE3XONo9KoSVibHJY8gbc/5G
CrjDred+BKHgfZR7pdmB2ZbxjgTUgllH13u+Fc3FEgclfVRP7ysMchdwyQSeQJoW
`protect END_PROTECTED
