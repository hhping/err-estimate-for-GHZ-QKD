`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XlnBeGA1nEbXTXz/R5bg60203ZJJGCMoJilkbLEz+OgUgbrUGS6Vv8bFk6KKjump
UCGIfk+4YS1HY2+vjjwu9vDqBoD7pCaHKvzzy38NmFFu8H3QPqtDWCWk69dKnwvk
7aE4fDIxqxTFMSlDdrD1qIJECgBBcjKYcj32xV/zhBHHAxjOPui5EiKktiOYFQXn
BJx3+lWWbBL4LzN7aLLecjAsWS2GdKwvDZfCyfKNkpdfrWIN8y8hKNWRgBqnZEY6
i7sNe/exuWRlGU14yabUEONl9iFxTY6HWJX+axY4jlhVXyuIOz+EPZ9XZeFvIj95
57/aJGH3mAfq/kr8mPVk+0OfIIWvcN1V0pwpzRkjOTry+yMVb4hjp/Vftj/Turp4
t9S+WlqSe9sD/YO99lTfsi5EI53IdPmmL1/CLTPfDCiDjRRQdPC83WXhF5Y8voLs
/8RxKZJ8T67QiNyauhHTKxZfMa9kJfjyNysxuqSSShfMpCWtGetex88ZXZLMG7Ss
q1iA8Zz2rOPr47Z7p848IqetMhf0EPInLJ4ST85azmSVUkjXawAWxx8zcZyR9UJA
`protect END_PROTECTED
