`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+m3yN+e/aRwYHaTIDdkgr5bgFQ3GAKmMHezWhkXeDGBXEBaMdg4UcJbOVKKSGKmX
wKyVMeWUibbE9QOXLmktkWRtFOpvdOXC5haLS41kqHheIp8It9F4dGRHO7jxRRf1
vGJh1KSpSM2lNNf+3cLzFQlFOz6swLIf+eVeDm+V5JyrRBzPMoHb/SJuvUgbGgUh
elCMytj/2fnT/x4KCbcdxB2g0dQ58yfV4aHhQz5L9Mpj5/YZ9VWBmnnrqc3hDC7p
idKcfJWWwXarYKYBsNjCRP6fLJC9JlvgqiEcoD6KO2bXOMP8BrJZg09PqZAHHz8g
HQTIqPg8Ix3HAvK7YhgPRTtmjWLCW09dUw5YTv7Y+0J6PWCN8XPqtGpa6wD6VtXj
ElIPYsJOMu2TqZZfttbI1lECH+K93M3URJZI5YPQVk/O2wRELFuMC1UapVzcOHlO
LScJboWwCvJet42MTRPvSQqs6lr74IxPuubkhvHybA+60WZPtrY8Beefg7HwRojl
NOJAWCnbmojotmOADV80XL6U5ku2GCouKV8cnmUJbeFBSQFhFTTwkwfa1YAVMLxk
KBxXiiZIaNbpqsFwoRxfdfrpI1WkS1kDMN3GaH/hq7VNiE/zyEEU5ftJxSAAZgj+
p08GnGyxAO330+sLt72+22DEivjueAL+DDjaggWcGdQ9V8BxNfKUqDEXlzZib0AP
kjb6hnzyl8IYKrZwSUiO6C/xExE7mMXENB6isWqKsRlL2Pr5PXbq4NCGQvtJejnc
BLnFF6pfQGcChGMLU6lKS1VRHIBD4ljDT1HHK+glS7NxGiB7/Qa0Ptv75w+dHXwv
Q20wZEiYSBFlnt5bT0oVnWxNGSDRG04QLrcEaN9R2/+7mQxe/UCJbQGBmjAnZWcz
/qAizHKoO4Wwzy3GEWPoeyVMH9qIsnnAhxf7LNNV9CgfvP3Tz/UG1BxVC+keUWNX
XDf4crCzKUJvBkk5PjLsNFG+IFiTxL2zwksJXTgK/JvdPmlxOjNEKkdvvFbrxlyZ
BrcP7zvNNxgmSHyrwXVksVnTydF8F554eOFnG1H+vxg=
`protect END_PROTECTED
