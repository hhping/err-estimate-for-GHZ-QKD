`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lnz0dWSpBgtpIwnSLFq8cBUYPi15CJxEC5Le7N5qUPDNirq1mBa2zKalH+kydX0V
Gf7UBU4WsAcQGnKrSRZ1c43fEeeURhF7YgjJ4WBFy646NdyrAxbcTKM/o3PRCK74
WxHlgopxo0SX3htAzaPPv9EEdhFkasSvB1SNA+0znycnH4MBAKoSPTfd+QaONCXo
ZIf/4194H74w4SMfOhC1ZnjZmram1hAEwdaEMyuxdK87h8YFrFvK5VTsRN/AVVCh
Fx/NkdCbcxfeJ970+qEcTTHTkpIKwxe8CFZMofPlNohLA2rJ5cm86+z6gMPGQDb5
dWo960EaYlR6aTLIs5zUB5MDaBNTNkiOOqHk6BnwCxJBJcl+6DxbkWDIJI5bd+T6
QCtuSOhxuEIm0sl+HojNMuV61SpqgWwrWarXGWeSFyKDoI4YM7M9kx8LtajxmKWr
JXguhwczdGHXOF5A2nBnYMxceKLFRBqePJUZwmyAdyo=
`protect END_PROTECTED
