`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XMZ4ie4tq7G2z3Avm41y0lITowk9hhY1W9gnRAJki8MVwiWoYx2rF7AMBy98cag1
1nmj/Mux8sxVrvx7fALVU4z9Q1S5qB0uaV2zoWaLqoMmMU48cVOVoW1PafH945TL
9cpOf4w98c767gOluFSuYrv14nq7ZC3Z/2aPSjWbr4WUFyI5VCO5gAfLEK2bmo8L
mOIqq8H+8TBrBnx0yKDfYlD+A+X1/v695pgbVSYXrErHxG0FC+Pq5svCYE/DrMB7
zrII0HwhZUNGjVS9M1qwU02hE7oJvqx9R/WtBUwZfAJeLXBH3+oxv9Ga1U0LS8b8
78M//qFQNlV6sU2bEzz49wmFwKKI6+23asfF2ENYV6yIohnjQ3xkmC1GTwbt3WNi
/ZhseYqsYUukHsO2VekpPFuAKIgn6rmLLyGMaEIxK85Qk8UJ1trF/WPCLJM8QiKG
`protect END_PROTECTED
