`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pc99IT1JyLvtvvb0CUt5YFMMprLLoCLhWzX+lgq8/RQOeA65oMJlpAsw+ZjOyvjQ
o3WLKg/oSjWOBqMAsw8QckJyhiTJvieSJfULtvJclM2f7w8uAuI0mPIaoByOzWw5
72r4rWmh6WZixThsV4J3liR8Ra+otRBRn9UZnb/CkZuPMqrxD0BfDPfDJNFZt2qK
PZYzQ+fvHGkiZrDcfgJdnybmfJj7NE84jg+DD5Md27FgIvMVt+zl+nJWn7p7Vhhi
NziGlikU7ennam4IDw2HhgBtm9WusZVPPWfKZJS7mxKFsXh0YAYTt6iF14hsqJth
QbaihVLOhRrb7JlBkA5veNpHxnhQUbrqBFbjU0xi/uUmS2KQYJKnyxW2yCHC1Q5I
5Yn6Rl7IzdRCzr9MLRUSkQESG5R8+JqXSSs/8auYy+/6QfnhGlx2fx1HTjcGMfU5
+nJiZR6aUpglNt1HG5fEUmfxkgWIHk0asOFkd1Yar3n3dZ6IZMO+tJ+MGCl93EuC
a4Ix1jKnDMehVuBH1mMhOocQhYC7c15ArjLuqtcDNomx807KeLxKDJtwON+wqyhn
o1irSX+lU6ZiFb+Gbhab647PI5YxDMYPTL0Dduc2rjKUQ8XmxpPgl60oiMNrftDD
yUme2aakgFyAZ+ZJMaiAwXd1gBvnb4kvJPFtNYh0rFDkNJOb67UYFMmsSI1XSWKE
yCr9NJ2Kwpndgu6/NiNoSXG5HWIT2YYBGIaBK2WF3ynO6NNpWFeVrvVE9p5eXD25
EKU+eT58qGL/f5Pjk4M5DTPAJQME78ukNHlbiX/8sLaa8/3hhsqMDdCw9clBngKX
dfoGZzDdk5aXJHcHUOFNGLNXeb41ObfU25Il2lSg+KdJpAM4/k91o6+ptXRyMDrP
apK8lIdL2nSAcY11Ouy4nsx0svx9HkSUeYAHN2VQW8UbmkCZf5bSWcnZhlpzW36s
k9OKvFD+uFeogHhrmE48w8VT3h6US2OdjcX8niUV0ik5biZ31vct5aPsBjPvf/Ey
lLff9aWhBvf5Boy20mDTXDOQJlH7BTBCrvMMwZ2hJuwZCu6B9p9bRGJN+ltvZEBf
Wju016Ktc+GmC+ylmSm04ULqYn4yPcLK9OdL0qHDm2s=
`protect END_PROTECTED
