`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ayyl2KYTZJLdy6UwOmU6qb7oQIl+v3bGDRR0wCBRxGp5nWyZyVTygBSKuu2xeGNt
1mxhLDJSOVlxq9225r7+sMNe+X2XoGj22OmIGLomDJCpBP7hP8W6/tdsls444YhF
A1hcTR8F8ohjHSBKU4FiD11MaNJCdxoBFxvvh7QqModhPGdXpAHQSPirW8Eii5+q
IVLjCfsUtz5rziP6Lf1rr+MWt7HS6eY/jXdH5j7YEhupnTTxFJtHpNDXTkGCtX/T
AIs82Di6SWxIV8zBwLwNPwnPzXVYgmowVtOuGktWcaCkH9rPKzZfI7JI+5cX06n2
7i8Ao5tD3MQsbo17GDGSRFpkEA96cEu76bVzpDp+Ea1escs6XX8WSfnJobntmeKK
QqHa6LeqqRsFBLNSfBvr+aok1LC5FrfZHqde5QPlI4ZQwiYC5R8WDrHicsBjuHVo
JUgsY3eS643qr0QmDqVVLpW/n2r5OX9Rfg94Ut0GOLWwtADmNGF4YYhQEmP+Ow2O
t3a7wKvT/QpJd+Cg74m7pA==
`protect END_PROTECTED
