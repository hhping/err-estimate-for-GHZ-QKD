`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KMtu7Lcc3kOcF4mjb9IUzcnlcuoUsrY56oqrfK8zvxSF56lDEHcRM2SUrwjmHTQM
4xDZzIuFgqYFmlDO/92620gEuJUKJ23ss4nNhcq3tH1knQeI8OPJvQAnP6T3i4Ae
UlyCEZ9tteBnJwFxSbSRdFOv6NkdKCFZhl+3kTgL9XqBZJnqT2NE7NRoPdE70kC0
69luTfnS6coRo1ggJ7USms3+tZQ4E6KOe3if07ZAacuVLQkT7Ru4l7BqpUBH1VLE
d1uWo4SY7JTq3aM2tq2xWdXSNc0LfHGDuNw862yyMDewvclnl2UIqghWnzbDVlIP
IenLJRC9cpPpJ/QFYK+KRpGm2BlNGy/Gff/IK0AH6Vk8s/8WIbkzVBJEVB2/Mngz
5YskfqEAhBaY6Mg3dn9FMRjyXsU/9XVViCb9ttXH1IWHo6Lbw/Gl0YrelTV2GAiI
eoStnGDU6yJYf2sJFwkAENf8nWiqAQzj0SEjsNQ5WrFJMR7GKmNF0duLovcvpsnr
uwA3rP0BJIcs5yF3/7vcJPDORgTIhFgPU1Fns0FYho7EJBUAh/aX17YV7LiqUcWm
LCRgEmmkDgma08c3Esxt2gWEOPOYrsN1biFJTJlCpXeKnC9WdZFm9PzvjylPN1VM
5xKIasjETHqlQcwJoVJGKWJmZXufHxQqtb16YBLYHbWmsjtn10pHELZLMeQe0syv
+ezHQz4Xy13k78gC6PaV/RhmY3nXp3CVxiiJd4rs2b7Ocvw54A3FcGaN5lGJ+m+4
htbhMIxHYcrkxA1YMGdYuQ5dfrq2RNfgOFCDwk/+Wr/A7JVuVOr3AHEPwJ+sVD1/
`protect END_PROTECTED
