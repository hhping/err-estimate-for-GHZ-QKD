`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jIJJp/ousAe3Y+9Hj91L8O2P1fqwFc4MWevsaQOqgGL30HY9bC2qQgTkeOE4mUOz
lm8O00XlTNG6nEgFq+rcaP/acda2fZWUSWM29HIlsKr6+YRyCRyy12vELHtCzLbv
y8LuZEH/EFgNWksI6x3iVCviiSk3kcrRiE4LQXB4LWa5nylrUDo+Avm3TPWgEF7P
ji8MyCfWWRJhnac2tSdxMZ9IavGVs8kpstAZ0wk9njsmRqM6xBf3M0Gy+BTI3tbZ
OYg2SJTjkN5IvfDChcNHNfin/VtfaaBDnvdZWGzBdqIpVPqOHXJNHvjRW02nXHid
TG82F2OC18K7xYhq9JkBttKpLCvveKgtNTi87AdBZNSxq1lt/ogBqHbiwemWQ07E
u5IdZz2tsrmeyXzs9suplovDPyzwDGHGpH9iEY/976xKqU2otIKKXCpu8nU6Rp+m
sYbqDFyyWqTv90+dRVA7+HNZD+ERm8AptAkjlXYrJuRSIKZuwneoR/cVM8JxJeQ+
/VyY5tLD1qadjogU5RBeuXkssWMqTqbauYRy4rbj1yMMGgp4QznydjkOR4AL3Pwl
h7T3Iai8LOFZ1TQM+hUIFr+6LQIrJixh2vsd78kBTN8TbnQbk1FwWOW685icokNZ
ocH3Z+vQZZnc/w0oZ3iEMeU7pjlEWggBMTSOb+NzoHnLujIHH4i9Y3BXc85wSK/Z
Ks3+TOrtPRsvMg57yPX09QLTCuBTjuoASn6vWe7lK32gwF5HwyKFfnLxv/Wbpfgg
d14+4dssIeGJDO3vo5xQaKoDyBT7eZl9MHp6oZZMe3WbLrAFBlpdwGpmXWj077Mx
EoqehND4HYS6NVngPs1ye1nyKKCyfLVHtNrTeRyJAD6BMQcNvvH0WcfxlCn9q7Z8
`protect END_PROTECTED
