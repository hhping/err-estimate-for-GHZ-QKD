`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c3jAI/+HlaPbpv41/dS1bPiU58xdyqc1M4SECGp6O5z0oRTw3gUO1mIpeApBT/la
OVUuteBrxq8xh+f/v+3ngq/0BzgEPH93pW619T4+jso3wK60m33cqJ1tVb7ThM0C
Eu/PNeDWa8YAL1LtaTTv+Jq2R4mbT8PE3pVD5qYgq2bTbtUSV4rmotXTCk2zXOLx
UEw919nLPjAN86SZPIvqclSC8yIL/ga6hluWO7nH2m96qzDTNISVrzLpsnf69/ZS
1T3ISRkf7ibmt1E3dcuF9hQlPxIk+uzfB/0yLEJmw7h8tchiqPIPrReavjdOJIHL
Z4E4W301M3Nsh94zQS86maUNjZjiRWzf8ov6HhaSJBiVxmPttcl/ZLAhWViVrd+o
3oEuaDQVCrn5L7KD6NkA5rgQmcreYLgmsEre1dp0EfdbVeO5Zr8EN+QaPL4kXDLH
TcsbN6eOL0Wj6nD87EcIyXyllC81TpDEjb5gUFBcCVZqhxCYNKKcqdoGkhV/xxRs
rbA49AdAh4uzOTS22C9vO1+JNavxy/i9TwFqCAnk2rH3GeDecU8QHB5DK264vxzN
yUMCW+hMGqaQc9T4vOGrVHYvaXCL9QlaHu6KOi2/M55FyA2T86ivJRWE5sA1hjr+
EbQakHIprXYKSlgNf3U/mQJl9+oYABUpfd0exgj3MfhMuibrZt9yKLOA4TOJYGay
MGu5FxfJvTGdCRuITxoqxohViUACKX9MtjLXHlXmaH3hLnoqMjYGcvQF+HMR0Hov
ya4v32V5uTFuOhMM7gmBqwCmD0+w7qyFLKO7LanErtHpc76ESDg4FRhFBnAU/yqx
NzO5y6lYtWTMcJw9PXqXot/PvVUskECAjMQuH26HqvddyQqW5C6wKy6b0SaiR4P0
0WubX6oCTOdH21hXmOc0KgKgMgN5ZFSE6Y3qXr7fFjGFNDDW0h0q1TY5DwUb3EjT
DeyPjiImZk943dTtys23g2zBcYqWhJ8TIjigjm31ndI=
`protect END_PROTECTED
