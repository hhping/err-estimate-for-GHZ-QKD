`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K+eu6odEsxEqsN0uwibJfdm7EGlVhXlr6LWBvJzHL49M1EvDoALyZn9FeYZ7dhms
FjML7av5AF1BczCntwtGTd9fTz7q2WNWKbDzmgEHRD8kUuqhFiTzRGGTkBRjYtEK
TdW8dIkHzNzsglGIDp39hfEudcYoQXMY82/Z5qj7mEunH/c0i79K3fE25vSbTpZC
taawYYmGeLrk6SP5NC+eBOETICc++Q7fLB1nD8G23r2HNm7Yq5JrhVusg86JVkYq
v4of6BlzJg2ed7P48rh1hFqyfvDC5fQSyhQnXV9tzBnT17Y29vlBQmQ8eGxd/63K
OeD8G+3xIQfgYqtXuCFWTTeVeRmRY+SuptCa5I6dZi2XgyXiukoqHh3fyNTwcoho
K1e5d2yaS7bzhIyP4Xx3c0r/Uwux2oaOWzhF6GkTrqPP9S7RSoLWY2jieaSRdAvR
yj1jp7JKFzkWGbyzhVbBmhRqahaEx9Cp+AQhCN9AhoCEUW+M+YMQs8Bi0JikvOiL
3KI++7+Y5DiibaeR48P/HZWxJ2cnXXQIm9nUwIbtOu7s/yNhGFUd6qvvahs0c566
0/3Bipi7DhNl7Gp4x7uNCpG/VnMruGWX53kmJ3y8kTnF4HlSXVx+1o+CtkBDW0oF
AgenWATLUuiZNzFfwhvLlUfSiLGK1r+4dnkL169gp2Ou0H4zGDBS6yGgvW6eIUcP
xX0qAB9eh9ZRAAkcIJuHuSOsE6Ky3ncG8f0Ettmqw3VvxFSV3klsEaexrUr1sJy9
+nenf9mOGFOW3q5UTZVovujb2tDgyQc13RE+ziaiIuPG8a2lOGV23t0yRCLQ7/AR
phzrfmIxfX6TsKGHw01oGlSvXTkfs5rKR3meeSd6psjxy8gZkeGBu1z8+JKPO2NW
fOymW437aE9+oybga6RY3hhbioA71Jijx2IfdHkbtJ15LlXR7XEyQ6g7cLIugbGJ
wqikga+F/FqEdoWkgkmnLjrS6mujvPQQb7lBaYsYP/mNiaPPIC4MjLJgudGIssVq
UfqI3u0jG3c+IXChSTXoiH6gCrEsGmSE4Scc+5fWBGHumPo5+3KaKwpZc6tDqvo9
745WEGRRAUD0WpBn2Rrypg3BLoww+NiKBgB1kHOZWpwDbvjfh2l6j7U6GdxJsWOq
/KLX1tIAsPxmyQcGFVG00Wy9BLeBZ+7Vt/ekSssyO45mxesQKNB70Dant8o+pOBD
3An7CqrqNDNeqa+8OpNRlLczNaNLfhLqnPIyD+qr2HOuewc4aSIV1Kct4fiFEzjY
yc25ifD5iJah+x0kn43AIdf/wgX0GuxyG7d9Au3bKNwCMzCByAwJVtcYkHpLpu6k
t0yWqD8rys4d2AVQOEAzPi1/J1py9bmPEu5qhM4EuCYg+BSNTT2ug6IDkGCC7ZqI
/v4IRTIpP9O3CSK/O7unLudSYdBTjSq2YXEAszWXwrQZO2c8PU4LSy6f3LPSn8+3
Pp0j4Ayr5YZxZdYI0yzCmQiO+jt2acbvU/8Ab67zR+MqNIp95Eh9Z2koxtW5z+Ej
TUPyuV3o1J9fP49WHsmT4BgeLug12n5p3E2KXcBTEfbfCniUfIhoQABjXOLmS3Nv
Dc46/9oORzS8AvrLUMQ9N0UjLHVDu0QQwU1PADqze/8zWEA0Cz7/UVOuVZ4MEp5V
pBS6LH157MQ+ouK/xnvPiLEusToPRVfNfKcTJUec8WFC2cqcGnD3S+T3nrwG5APF
kKQJGli3MInfBpLKQWFfMGptx5uy+ZyTRfcAT4PP3B725aEcpt869sfO1mGgLUMW
UJK9zdW0d/w4P5HQ/oamihCYKTlnO0SRB9S+p8l0l/lS+LavZvgfIbm9vxXDHPsP
yT7JzyHY4wcrPln2aqeqvCTVvvR+E1RNoR1JPHwVGJv+Lj+t8yqVJ10f+7V7Kyyt
gdHM+NvMO3bgVLbTYL7ngoZiScWqbY7KCIayOEWWyCK/AJPXcRPZzwN0DBVdvVsG
+dS9Ex/RVtnFlYZ2c1OWiecaYaU5PwRAQoSi3V+1yW65/MUZb62grkgQiXTDUhVa
ixnZowzOn3iV68OerRwRQgEfDu4LN5tjeOhKad/6AhGO4Z+Tj47x/b/R+3M0g+NR
JYSgliF2FHsq6vkU1TqfIExXQHOvHuDWz9nqDK8nxmgCXohz/VlG2XjEy2lnkr5O
hYpS0yodRszxTkOUgj5xPk/Mb2rynAPx2J2qDDYPFpsBDjc6FOfiQh6mKWhkNGtJ
6ZSf2PPJNPO7UWqtEDcRsdiDnVB0MkIIBa1O0BFQlY0df/H7tWJxSSEgO16bpsKN
KB61fjdI2GprhEFhIrhGtlRSOK1rscIa6VmZYLmsM74u6rrwPw4eeRfowiN05XBY
HmznYcYi2HcAvQkc7fI5uXKeGj1G9SbyN7LQY7TYAhTITJIZWWJWw2gQhtodzGf9
KbOdZwBcBfyM6X+HYA5jsBvEbfWmfRhopNNncA9syQ+m1gWXrIUglaZaucyN7kB0
utPZi+xSys9UpBiggc1735yl7aoySlTKYuGnLUEtnVZ6kvhsv4uSxUsoMraamhtM
dCOQmVKKAHADVXV6h3oJ1LpN4ciJ13YD3JvzSa1wIzbe0CN59clRGoqaB2dn1csY
jzRrrZOo3gjp9eUNo+Iik2fnxQ5uwp6VriY8BXTi4IqPzcWT0RbAABoQmSRBPw4b
BEdLdgzg/8Khp7RnDuTGM6WbC8O8o2cTOJ8ZVqPUjODZ9AQIhn/8em9URsPQfC5E
kcUD0yQ8gvXHo9ygYIaNUEnRXZkSPbKY8Lm+nYJH6EcKdir+eERfBcSge4JYxiIv
wgOl6ohBBs+LsVuBgyCKghUvKNDDZ7qVbqeAGp24zhFsIJ3rRlgt7hIjMDl3HSdr
A6np51zIN5zsysVaME7KnyW0vLgOuGOV3h9/XRTjb0F47Nf8+6lJOCOHxhQet/39
Lq0IU6/+WkDaFLDJFMuG5SgGUvBUn/4x6Bd7Wn7uCJ6C599ty3gUYe+KNtxx/pfP
t829/dU3dtIDs92F8Uk3lxAgHbf3cArtNIFhpjgZnJ95AuhwdkvCCMGk5HmeZeVw
1u3MryMNbknSoYh7dkzmT4AfZa9Q5h1WEX4XOpMeo9nYH7j92WsSwPm3IM7ioFko
3rDDMf3lcxskJvi1xCMKmA8qq9zOBNkuTJ7KA8r4TtWbadbShVAbEPNe/Z0FguQt
Z5byS8sQUOjYmygrX1hzZ//TZ9Jj2pJCbkDwC2qs23yf+WaM93gaq/PH/8IxZOVn
uNIMd1YP55Pbv0Sl6p3BpI2WtjONdoAj77Z1YiaONBceCJdXav47mtoZyUfKrnll
8l7J8VWIrYKHHkwvKhs2AyLlOYACkkTfLZt/yU1AeuVuWJdAg8HV5tQuua3G/UbP
6e027p9SmHQoj0rrH7+wk79BL9VrsH5XBlcB7hIma37Lj0r6JrlARsj4IonyFllf
6nxrAr7NMzSA0y43GRu8P25daua3QMS1J/ZeRX6SQnuqhkZFIZNbuj9+nnMMxCWd
SSWSHwBfLz7NWIJn9GWwgYiNH5272baITmzbOndnW5pzTqQMEb+HXBF5DXwDVEao
eYzpo5CuSBLGxrM95934pOM54rUBqKqTJ13Xi1F97V2gm2Tix26+ybq4nAQN6fcP
bIsV00isBlqOJWItS/i9RLGvNN3l4/H4AugCTjIoN8k=
`protect END_PROTECTED
