`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8mOq+0T2uitbKIVa2x9GQVyRRrAYbhRox2eYncmzWR9yZdk2faK8dE8X1BlL03pX
MGigzawXD3En7wBT2nGmzO+pZCD4fO9yYKaMGKv/zvJeVOAmQQi5j4gOrE74kFEC
SOICm58TsUL4BE2k2XPnvi245XrLdp96vKuQsN0Z1ywbnJ8/lspBK0qfYcADY2d/
hqf4GkQqZaL9fw2dOduNVR2mJu/wO9LjqWFHVyqaFW44MkrY4O2+dpmdtUVlPLKk
VkBOUg+AHJbHr8OnnBHOKY9nDZv36wfA9G4QryzfWwj/Y2aOnXtSnpB9x9xGYvQ+
8FVzE2CAH/7ulGxeE8myyVLXFttzuSL/wLsPybiQBvzqQL5/iXe64zav3v7wU2+7
t5Gg8DV/4Rz64SrjQYUg7MBYTvWPVqLEQ3hlF+TmFsJiPWlAPXQqbnGsqKTJ4spV
8h0Dbj+6+uZ3W9Qr83UzVeFOBf/Gq8hvJV65xXaL4dYqrrvmU0NxL68fF/bB7/yy
cU3eUwFkod8+k8lbqkLKHpwEeYzxezGF/Y6od/6iyAccK8LU44jNOTgga6AmTcID
elVdaFGRhaxCo0X7Ui6XSOGqYN35eAb57pNY2Gd9xmHHd1hnTZI8H3qRmuHMG9t5
syHOgtYs7VHf+/4BBRBGpHgVbMVFYZyTrMOnmuMvpE0778bmHzvBU4S4CXZc8/H/
DWQ1JLBgEEPDSDzmOggBNHYepVv0O/aHWqbpoWuBm5ztjuUKRBLw24qVrJSoJPqk
xthBD2i/x4wkGRaKDTrcfUTodybaA3uGtOi8HRBREs+O3yx3UWS2lJGFb7pv7zjs
Gj973AV17q11vtNhcrFrGGIDldix/ZdNOpnvqw1p7owosKT6G4t/ZOJEvt/5CiN1
KxID0i8N4MMWIJ1ZFkNIWlt2MTu38Q8cL3pwbUDoVgdU2D7e6Yg49OXpT/4HBgj6
Hc6xfjzbAUedftbEqXJhfARs+E0/6iTDcwPuki8yco+sGmQPLh5JltVsnLRIobYy
iO3bZ4TuYlmANHEAMoA6uhZ4VahLWHtBo/+0gRTrolk4mJBLjzu2ZZk8OayneNio
XTV2X4Hh+PeQfao3GLlfSAeg3MKJIk7liTfxTDUyzP6lb6StQffMcQnPvPB55dPq
a5aCsCY8WbgjFi/xrhFGBE7nynGtzH5DjO/o3vD+yj/mM1gXEgb+9bxRG8nBWT6W
uIIYFJ9a06K1qEnWKQhwzJsiZegfYI5UQzeqls7I0puXrg3q6bPuK2bqQymey14i
3EXuI3aouAd9RB0nnIUbCONbpixjUxurSvtqI+mUZNygrzyzdoFeByNxcT2GcL6/
8ui7iCZ19ncXIT+BmMXW9nGcn2npAeD32nMcfh7wwEjE5JaMBPlbWm6gcHfmFtMZ
3NVT/UhzvgkCmT/9AY5al0xlpo/7KFzmHyBDJV2MOhqbOmTFGNkFxQNZGEFIoNQ+
sLwryKPsAxEO8Q19J1tmwuGIwd18yLRD7p5y3N7SaDGrFZcowLqMVJfONH69Ct3G
gZw8W28ruO2z0OlLPeIiykM+f8dJy3eowLZM2YwDZMocu9l5Gbp6RTKMGFpUKMos
UDAjiFRR0RrAoUbCgcIimb3oS52NVPIktWuklLGMyTJct5gs+ZGQGAkQM82cB1JH
o2dyyyyFFhtUA5HBF8olpbBVQE5kXeWkSJBmJOnEbImMmFN0TF3s4my8xhzRUVni
fDQ6NuRdbVEsELCI86Kkpfa3s7WJCsjq6mi9og89Z5dkpcP9QijMmu9Mt8KZord0
KZELmTnzltkhgxIfb4iQQibNDGhvjuKhtqc4L2fKguY7fbZc1rLMNaELKbLQL9vr
6ethZLBrgKWuvOijQq50Q0UV0PSjxdr1aFbpnISSS9e6xZ9+rSsDrfuldMhP7cLA
qgCvK29sZ1LXWtuibf9GWhS01hBgVAQLUqOjTipOqEg=
`protect END_PROTECTED
