`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qrRKLc8dN3gnIGWocP3ekw09eyp35cq3ii5ifRzAITDi0/H865CCl9eSjU/OBWnO
KSLTv27F7JLWuyN9ElHRVsstmzeGAEZPbaC1tvoi3x5Fu5sz+FFzyLq9lxotPFIl
OrmU+mB9GqcG7psGidCRYOnMeCnINLxY0flyGb6ALqP+8P192thctkrWkNv78bUc
84oStQ2DIeZ9piypNEaqvA1dGDf9zJE9hHmGcIl4WaFvU/oRDjd/yY4b8jvK2e+8
j2fw6BVsh9m7ItSixHfNyAgDZFM35sMP3O8ALkKcAQ3bqDSx8LOAFNiQz94yyph9
Zq1yK2RyyPb8EsAO4koFU6xPik29ykHIP/At26wpw1RkUWOEn7cQ6MwXWTgC3xb0
pknB89r+YifG3Ywxq7qiikRs511q/arWcT6lgCD+zDtcNygnLSsl+K9trUbD2eh0
0omuDnY5SonLNH/ojlYAxkJPrqXx89O4fjE9GLsi82d+Py1+Fu1T2yxrwSDkpCkL
2kkVGDBVcVscpVhCLHoyIIqHe5caxfcODwoXsywp8KlPd/efmAvI6q9TZDNF/R5l
UruU2I3U2yXFLdlSuI+raOPYcoebcqDf0tehNGV6B89mcaNmZnxeesx0onYVc1aI
Iz8tTXZCr6wByJqOCYq4HUmF2Z46MgWVkVt0rPLo5xGbZoNZ+hpZwKmWibFuw8N7
YGhZUiMrpE8SmhZCPoKft5O713d86rmCRLM5niHA00wbVhHUkFq4seIYL0PPtX1d
CTCjSYd32SYQBXwryHXBkPwQuEt1jAv646QNPKb1Ta9IkQEfMvOUUglO/5ONFYq+
HHd8NqBvlggHlm5WQa0Ws8JN5avAIAEh+04om89GGpZhlYEwJQzDOA6hwWH4pJfh
cnHLJZMHWnDFEKRLf4XYu4d93fTCqQF1J9Gyia+/RbaV9XuXtS6zyFqvX28L2ODm
VzpZ2wJ4bLK9LRMfxcABjLIddrfrYqomoeW1DG4HPEQdXAADHET46YnGJs/S0BtC
buCDPcwxsswPz+tO0z54wWb+NjSmob4LYquPoam9Psn5rG6Nn1X+DGp3gtWFZhXn
AbZcu/GXqz/n3jyWSPtjbdp8O38lH7hA0ESul3sGa5ULsXAsom9aBoejbrvcGneq
IqWnNKiverOQiKOf1hG00nYPHZae3feWu821Mwqd6Ktg/Jdp8m2p95wNx+tKjpZ9
PGRpgtx4EAh9VQyAcVpvndc2PkYI+r1g73zNFQOFMYo69jT6iEkfjrRWQx25pKud
KNXRIT7w88GE7ymnujMS+TUOvzR+Uhq39O4fMI1Dw/txtcKAvXK+sx6F76wOf4MM
0RB++hzzs+PMIK/JmwVmYMsHIlskySmpTYn9gOjl5KR6QbGKw0jboOnF/laKK6B3
dhFzYhbL6XuKPZiO1ozXFV4uqc/aGgLoV4cxpQSKkjETQax6xHlSvI/dWr35Manm
buFujNlAvXePHT+hgHe1mwvmrNPLWfbrb6aAj8peaIpY46IV9HkJ3xWmXhK3O4fw
N67iSFklzXxInIhEyA5TNkj5qngubRls4GJSaaqH3rdZ4YvDIk/QrE/V+5BQ00QZ
3LonNrf2tpDgahZ8wqSoTlVnmOL5z+2mEyBVAo42hxXjgd8qlUDCnekTYy4IF7z5
tnotiSA0Bbt3qo9m6PKl1b52QnFShifpH/cbpbm9IjZ53jhWLq27/6NCwlLiJ8P1
SU0cPlJS3U6/Qu72R5J4B7y0ew0X2M7N6OTW+YyIcimFgkybBWxje5B/OE1pNVZ2
GU8tB2g0pQP4nyMS846SPqE+R86rzYbHFzI6GtyiLelR21La5aIkc/uqhnZErd4q
IgW3BWR1z6AIcQMHDAvUQQMkmrQ7K2+qFlw0MfD3TDdCQI5Ha2D9WB7vxQGorxVH
E4N5sr6k0Omi95G86j4NucOsdJfEog+dT0uEkc9Aruzg+P4qNXAceVZR+1uEoNCU
owHr9e+xhx2DMUQNOOArBzw83BAFM40N6jsvN7riefda1SqBVdXAsv74atUCfww4
pkrGX8x716rOnyz+EnpNcEanpDs4W1pJB/OxraSDYgFPR4JwjyUAhXrNUlw8ym5j
RRNYuDhM6G+mfrJHDL5V94RhmdTYzFktVxOn+gDfUvl2gvNdJbEobRYeBt4mVwQk
Rw8elrbhwbIxI+mAnu7oc/vGoM62lVIG7wVlJ/oO2wkMMEU6yxc847JSLEdoByw/
fYH5xiKGhigWPXEnhEc0/H5GBnwvMdurGQCTyHYYZrSqGG46UCWB9bRMzBPBeYEW
7uX1v21iQJjC5OA8c3pCOGzTOR3IsZ91XzWpY5QZedL285INsm4QHfs7loL7Kb+O
walM0vArizTZR5reDK7/lyLKZIikqoekrb3WkgZ1xR5MLkWqyXMYpBg2WfDqn2cL
vuAaajnNr5vybtlNrG0Yvyj1BSaY9Z4W6gJN6KBixF3hsAFvk47eop4UZWWBt19G
lqYExg40cKNL2nCp+6AF9+8PHVzn2K0a7MzBaWh7DGmBhYq1S2it1yHLBnZeKqEB
wqAUcZ5hjaq5gQm8Ok8vMT6P2YqYuSPU7xbfB6r4s28n7Nqgv10mpYCll3StXcUD
ElFMP67qSHrVL7Yvo0SHCTmO3k6i5q3MVJ1Zqu67eazt/f9yT54t8F4MTOfij+GE
qBJqu2ZzjxegphxA5RfCMHp+sFzNpz1PkAmQQmEeY+a12NkxM2ATKXcg8guhs01P
N80TeQz0wlmIfDhF1T4kLzS5Qcy+qLzXLbCfN1CapB15wpMOrEsFkbQ1/q4DVerY
RmsUM2p6Xqi3oiPSaDofWc1JcxwdpewNmRorrEXvmjDxShGQrHYhgYl5ZTnPiqrP
Oclmo8R9B6XjWmpHZPMlaXhyoQlle7Hii52VYbL6dlkk/Eli4LPO1i4RXgFeXX3/
u+zAfyI00raZ02sHpf2wquW7Sb7XKdb+VHgubJu+MUvQAKYeI9aIvxFAC9VZ6LPJ
ESFdnh5w0eUl8jBviQ+ZwmZ3diLvNbUunjghCDsfjeCnPIUyKOVG267U5i/PcMce
rxdNh/EfgWiglbyNaEUwLZKpssihbKFFAY4Zt8Zf2xIGDtE8E0FJByyFAHcC3McX
Rr16OCE/5LOqEg6DBvQFbaMXo6cODb6iT06XME8TH3fp010FCwwgahFonGxs04+/
rkcqIcEv6uy5YUgj6vJ3OVqp+ktlVmrhl/kMVY62y4rLAV2jbT/NwoTOTjoP2Erk
3w03bi994QQPY8/9qsD3vFsjMMWhqPP6im1cIgdNKFVD13vHxEAfQ87+iyqhC6pw
1KxcUrhLtw87DParF0m2hicaIlvRWEGarA6mn9GNmetDVs+lkt3b7L4W5M/W4gTQ
SMiU8ayv+Pw6W1rqYbx227Pv4/4r93sHB+8OQ6G275UooxUKl1cw8hrs2ZsSlks/
9JHFkBGo54PbnziKyDneXZ+CUuULNATJQJGKg8rt0+Ke/e33K+Ka/DbbCSQzPVhM
zuR3zERm9XCA9ryiLsB7yZRuIrsOdgZz1zLBa2VE6AeIXy2qRj9II6wAdnsm9gp/
TKyHZWVXRJgW1i5k+OZRKsVpDxFPnjoP3gfbbisZmge18O/50M1/KrwRTrLbO4xB
XL4UFqXqBXb0bKQkdP4tH1ArN/iwq0gAkLlhg9a1t072h6FZEZP1fd1u93yBJp2q
BR8969D1GokAAXfC/8hmixKrDOD0B+1n93OIwM+Q9bk88EnPKOCP9wEk+QarwwIP
0+7z4Wz7j73DCsUAyK2ZhN3Tm6F7g5kKNc0m2ahXAKfm0M6lAKSlCPtZz1VyhDa6
2H6ZVwWIqZIEF9qSE9gUvt5d+94pxPrsQLME5o9aRAitHvrUr4RY2UXblxGKteHY
h/ylJksk0MMgoa6HrB+rHCDX9daq5Uq1I2xyd2ozZsKN5wT7/H0UypNa3MuuTb//
I8ZsrYH3ZFNs4SxmvmCCIry6ivobPHq4F3a+OkhpyihLbNxnXOxWb5eXU1JGVj3Z
7/kmaWUMpthCqR4jMDh+L52WxSHb8RP4unED4ztsyEwRxLXp5vV1vWj56WKNW+1f
W2d0BehA/7l3DT/53TrAus8GFreBTuYRfwEXvZ6e7BxaR1UDiiehP6Orw72o+/Do
aUqxy1WZDGKvFoCq4WXnlRvfK5B3lnnkLhX37NMP/d2oJh2GjvAaI20/SA8DRBl8
VqDm7C+MmLZNjbSb8cE/4krnMGjaqOpyEapvLQfU9GV/2xH8/EUOZ0+Qin4gTeKh
9+LqI/RjkCf2uixAUlH+kMTIkUJB1jssvThG2SaW8olIvPXR8kjF4n46xN6c3uXF
zj89mee5YpI0In0COtd4kiaX8JJiCmIyj/PUPFQQyGDrKih+28wIbiQl//HZ2z2K
L8wYCoB/Zh/rnYNJQgzNxFln9od02NjHtWteB7SJsSsCqcewVy7aYmM30DWfwaE3
s3UUHdM1OYfespIjaui1hK/Tegq2qGiH1ztKkFc+EOWuUyIo6fqkpQsgZ1rMBCVJ
ZuokZyjw3n87m2oW0xP2KPu8qV213ikEK4z2iNia4x3Q3qbCuftR4fjjWkNOVkew
04AitNFj3JeaQFXS9LgGbL6D2c/EdnWm7B7KbCXdlpJzEqudL3qGs3JmVMurkj1R
VgzLbPZDm0SB24OC+SroETANLW3WtO2jswkBbKUE/GqTnUBSYN26bpZ9+fa7LGnG
Spl4UgIYnQgrTWdNX4z+H604TubbZsqCo3QkCi2eQhPz/en4zKHEL9NR0PTy4VEr
NMNFduxEwauR+PGKz+Z1RwbGKvnc6G8T60/OauYr9mdXio3t4cwLYlTeV6ObinlB
KG0TCz5QEJT26MhqdsrdmMGStTFNeeLxgu7ql3RFo2bSw+B3fIagDf/a9QuCYdWI
cJYgwUaSQ7nEDAMd4ucNqhwR1Vq6WK5pz/BizrK1fookAhNyH39qJcdRUcJ45BiK
mWkhRysmrNEUSpDyh0Xe2PJRPfU0D4d3eRcdcjq15RCGFpOe2VrfridGwnt01SCG
KHhNuF0yOQJOrYqDPDiJZFNjfGRxANeAOa2rH5XoEviLhSkrTpLb0TBT1LEmjKkS
/bMIf6nn5o3sc7c7sfsjyAxfHHA1M6oyqS3+k6DLAioDJ1MEocpUnlIcv5u8gOQS
nQv3fvQCvnTO3eGCBtKckpN2I5IcidllOYGlMYZ3g+YaI2PP9knE13ZCe875mxbQ
Zmk64QlctOZxgpK9+w6gILRZa2zEPbsm6a60kFfHuhPCLwxlsOeSd9jTg6QnzbFT
5hnpw3z9ofl/EkfGkUcOL3cG8R1Lpbzhsgs84ZN/xVC7M0UhN8cOciX1wCwUok51
h3GDkHyLrQLTwxfMXaJ5jY4eYsJkc6R2RQ/ya9vb+2Weu0oFSqhTTy/dU0T4/ENh
0/BtJUBkFhTf56lRZtoWZX7pqpgVGYn5feQRUrsxIxcUm/FJpJ9T6hKeIy7mjasp
kNjEzmhYPIS3F5Knr7CnWEPJcM/tYOwbS9qclLJi6LgrDqzy9cm9I9fXfupjy7lz
ZSLL3iPMmUfH2B1C/cGh0W0wdYPNSOMzvY2N8oPcVRO+jB4xTCgoH1M/aISe/s4/
w3S/C5dPDxbhtytUEtBllxV99QRU8nk8g/m1iCL7Irj3J8rlQKRfhf3l6tRmeD7Z
y92JZrU2xPM0nde6g/S/oxgJCj+pvagOIKu4BZvZweSxT77Zyx8yg2U+c6UwSmFM
N0CsfhZSMyFdrSNR/7LopDpwGwZTL10xIY367Bj7gvo5ozSpg1DrDcLw+EiuMElI
cyiYRB/HbXgXusW/ehWRtWA3U0eu3AThY7JFrevI6C+klHw1p728FXrBBr6/nNBd
iL1TgUzMQxT3xmq7x8SG6FslOxXKwwcJ7DyqIh/SGgneZzP2PyapW4PwPmihRV6x
K1/AqBID4DLJbGzbnp1QENbkPHizGxMyf6dIhF5CIVUmIMzbV7sbKKBQpjkwHv04
qyPeZHsVavzjCcFTFLy6SqtSkpsqn/qGSwPI8ZJ/G90N8b6r6/OuhAeopGMVf9pa
CCg+tFNbD+zLEQVHo0LEP3BgSnbpg4M5tW3jWaxd74HuTfZt6IEHx2S1gfUSW3HT
tSbLR6LMr54H8MamG5Na9Yb93qBRVtOjl7dmQppAJ0Z22KTzMbhubZ3VcMd5mgK6
aPDhPquTLmXjeu+h+KbhX5hATRHZil1iunn2ll7Ta0H5OLHixsvKCyPhvTxZf0Cs
TPSAE28/XtXrcTKl3rj2Cq/BXmlK+SqZZgsJT5T6/uV0seUsbe7wZIXwZtKHyTQW
9XEhExmGj/8VwjzvCDJszN4384pD0PVqu31Xb25PKKvunWyQkjhwLpjM4r8oDXVz
LcnATnmEqMY2UMXma35T3E0XAgeRZTW0U4fKpqbm4BJO/YCtKMH23rLOlbCS4TeO
zuk04dQlP10nnFhTKRxMgHipmGuWAD/+/gbK374J8TCmlft0I7n+Mbf+8aAIOZmF
0RxFG7UrDc4I3pCbJp1niClFP8ZSkEm08T2F8xgnkNbxKS/sJkiSmlUKn9qug9sz
pAwVoFx6U8W7mT2LAvmLZJg6gZt0e49tpbsa4wBKtWegmplYaOkL4IZZZeKy5/PA
oxqKufQpwsmFyM0dcxZaQsG07ktYan1no/hp92hi197YbgdxnRom1s0T3GQGMucZ
E9ncuuRecyvtBQWog/SvW8vRJy3/nVDA9aaNzgPN33E2ZZxt1kzt6tPl0fHQsq1m
gOvIZ3Nu7tXORpnlUpYOz6lm7eGjFPzlGHg2Lx6aae5Qp7QiRZhPK+EnCSekCt9K
BRWUVs5S+ns9cX7JVZDKmwRbBHNdLiwwT4w8n/d0QK8EdgGNO2sSzGinDnVUtrMm
CsuwHc7dPeOWFgg7Qb1Z90+ZUzukXHx2+HVZ+Epq9JrgJAjKuC1r+BnVzg7LTffo
QDRk1ePQ9O0TjHdk+jGZlOmqkrcOPFlUOQMu2tn4WQEQlmqbwKXLv9XnlZq52oe7
pmnrA24epqw6U/HicDJUU0X9M/sZXfCpjQX3+KIMWz1w9Mn/BNxb44yVit+yOMhL
+TP+YnODA2ttQ1QTlolSdf4drkbXOADvMuPnBpLptppPrlvJXTxJiLZXvP+/hNuD
G2ZtnkNG+SU25bn5ubDvrlBA8hMBZkZhYrNixCUCV3BHo67kuBCmDyBjh1K9k9k9
bdHRnp0D4D05dMscugxpKYOeX5hK3e2xAn7fxorHSxs7v7nMJ33nmJsgnoIhXMFn
YzRgVNUYy2SeZSZ2Z51qbXqgh9el4aU3Th2EDqsS0iXmgE7lxeBbv59qmWsUQknV
yTwa1Hdf0I7TglUU+mGH5jAJTMFlFAjGrz+45ikr340+6w9YVxVcfDNvRqsYe0v8
kRPny/yf/n06fcXQsmAGpVxrv0c0T95f+ib+dBK2mVN62/AjlsmfxVEWt/Uief56
To9+oUZhXEmcfMT/5DWPrOE37jchFSSLvvzeKaJAHGpyq8mD0zWqgFO9MyKSCZhy
5IdK/z52BcHVC5udI6S45Ya9Hxa0RVexcIjM8KyAxUiCQh76xZvAkDVNmNeBTRq8
SAg8LNz2lyTG4LwaG14cp31Aqh3E8Xo5qe/4rQWAO33+mq3r47N+R1AegqjbD++u
XwZjk5554dEVhr0T6Ry4qfDryq7U/UKm6hXknJVBSuEpRF78EUNg0FVxYKZjLZRo
/YMdqzapuGFxag8jT2GH0J3t4itZKJaGpMPchTvgh5+q8gTXF4l0AvMnLQE4EOjg
rU6J/NPBLZAmVWzkhfYwzx7tXrNza2ZEAEfAq0vYS9EqlkzjXrG+1Octei6kiSqF
SXQ/Q+8QdyLt2zwh892h7aDPTs0VRflyFgnWiQujEDu42JH6cfo2V/blHyuj1iVI
IvpQmD1Djnvm5MXYOnqIH9/U3IL2UZHVGtFCOz/pU2wH27yupsuiLXKSmMusv7fd
XdmRjRguPN3ue5b4vcpk1HeRPrdJSES36P/1IVcQ4f6SCdDumXAS8nnRwV3VSiJo
bYivOk1Vn0yu10lqoN27KSTQfz0oYIUTCacLU8G0wjVv3rWR4yglpoxqcJxzWpFG
djwJnC315C+W8ecYr8vEEKQP6+g233hYLjrJlImYeKVMDqr8V2PeRZqJ3vxU+kOG
yyzzErzb+APEXLMra9bz/neiEQawMXQ9DjnyBA8Uv6PPxQFBxbkGPVfSFhPKelsG
gHHUDI9hDF+y4a00y9yLUYsKrXtzTzZ5bh/VLQPkERMqLpQGtenB7Sgb4CXYpraK
h2IBpQoPd69sD1Ldb7uuoqedOBd1hkxEusb9yibFNcXtHx7hpUgNCUFkZQPUC5gT
ywd4Ho+9qAuHZ/WD/hzm99qn+S+/DZekAbyoH9mBCGb6+aK19Vii6hbn29OP6sTr
79QODSmwkNtLZoRlRq9CfEz8g4nTo+RL/Cfi7SO8rlZReIRGE8x+yDwI27PAXoJj
aIkOr8GmK11YvBIGe9Mx6zRuYGyCIo+bTysS/PQ4Xb4ko9v2/7qKAhJj6pbv7iSn
qY0SOWur8F2Vzt6D4KYES+t32IZWFEok3Vzu8DOzDotGx4T4lcviVwCxwNbJdGvR
4FNS83/bgEFHenHwmbJiTJGlWJY0O6vVU6ws825878k4eZGo0Hb65vqKlQiyVziR
WvXCBpBiTS8HGdAAdh2mOMpUqxgdQuo7qh5m8D2GdB/cmx2mgv9nzwcfgRwM+VkL
Wp7hVzOmqhAzx+AkB0N53KygPJoTlp8TaQgqFdJEjwnV005MkUR4Ylp/FW0Hv9pp
efKgryfa8OnBeK7IENiCyQlIcOGa0TAPV3vB+i3vFDuo3/zWpIitn0V1jDU6B6zD
mC6hgD4tZC4zjeeW2mPDFa0xwQNbjte2VN1xITOqZSiIdZxG48wSSS0MAHXEmXcD
kFDXCzEfxNOd1zH9QOd+hjUnvhkfgiO/1a2wxkVP47mp8ueGqR/UD+ZIQM6ISu46
nnTJG5tQ/8lu9SnKwH0mUXpDcRv5yFROws5U7exnNTgxIxLuJB1g2eklNNo/bZWC
Iueku7uqin9J3j5lwNQaZLzu58bNM+GSSiviIZEKCoJ+XgW0rS+K8qkBLYSVhV64
6/oZYQuqMa5O86L7S2E3XSj+y6jtvfWyLi64j+bZBR9L7Lmq91ouvsMdDXcFoH+/
RZ+wJNdQlp/Nr+xfV46B5CJZa2BPRx+Sd7FEJRllwfRTv4dPrs+atVas/glgZ2/N
DAjYSHM82KrNAFqohPY+D+6xcCBOHV9PlX7nqfBvttrQ8qKcqg5Qg/fCepAqwRm2
rHGjYac0SrEK+bpEotiwRmMTbRyBIJsKNlJ5+oGdpuBn+qzgBgwU5cSk7NoqW+gb
qkhbiV7K7sB8+Awb0jrghAqHYv2HCOG66ftfft0y8VHgMDS1GtE0OoDSGjtim7sE
LTGi1lft3uWY0doCbx+QWtjTTJQnob1CvDE1YXPZ6c5OhzE0zF7KS5FVSWFFNTov
hb+I4VS84wkKwPhODFtwuvoI8dtIRoCfxmymIbFssph00RFddwG7TBdeR81V193o
VrF69zDKf7m9/RVzgmfthIhgREjGG2Pr+YhKBwirKlAn/RadGydkXIlCt0s7+V3c
ThJy/CcTv7me/87FswOoitpUe1P2n1QlxLmZhgsDlImol8lLR/f1HdqPRPI8ZLUD
ne2Mh4zJPBMD8hCDVs0h/7k/hNWSpg31mDHSAqcxILiJC3b8V5fp03dOZ/Rv91pg
Sj6Qpk4FbwYtomvM8bkt2bBEOeho+gcxhNFjib6SeodQm8dPAfd5zWEwt6SbUsY7
1O+EOTTxE5uoeUPSvbNGyMSAd8iPL8Rrwbuk0ol004pndoFB/3Qbq+pXUHXGDoLt
VhyDorfmgFpBcTgsecyJE2cXnZjDqKe3h8h95trlPLDeD1PFJtKORYSo4d+0auSQ
DlXTqxyQQeCpPRZ/lC6tzY49drAnKgvr6j2Hu0I6VjTMx281YqstTzpg4GrS+L55
fVtfnzmLq/6cJZ57iQXsg/rYY8WPLtxDB48NM8iinPreBCshQkh5WU1RsRptGbeB
6CpDFmspiZJONWLKdMd0I3nWAApGccjfNDVS3RsQ85drMfQiNC59/IH5jY0X+17R
MmNRc9UQ/No1ubMkWxk8ChvTcRUIHfM9lR2lhzeQVei05MLzjZX3EPJzJqNyQ061
4mhCFLDa8/55E2ETB0qZfeNl2fi8mQBo6i5zd5pYtGDpmoJYY1m5OYxQ6MfD1NxJ
HKO7Dw8waFueMNo/V4KcUMcwmaeVRJmv7G6whhD7w1y5QMzKsB0r9x6RBUdKlwhr
dvfx5LL40MwZBLgK4v/8gaRPaeqDy/PmX0ERiuE6IqbpD6u3gDUn0YgcbefahkHv
XnTQ/qRa7a8AQ4/sxuFUFI6tXgH+URX90tRJIwO+ZtnESx9m3d7BBYRNL4Pig52q
riA61wvKBqaVhmFACI5UfcDL+V1k6QCXvx/wiEdLRgFTZ1CsCVAI2Sa6AAVRXu3f
6ZlHiykQZx1Z+HiOx3kQqBsN7/OBwDvOdnrfBjbAB5MPRhTv8gzf+t1WvJvZu78S
0b8TpKrPB5qU9V94yN3/cLJmlVl6w/SNc4woczsiWGK4tLJlnOojhiZMozmOjmSU
a5qk9TLovNfgmTCzAB30GwAey7y/aQqozB3tCE+yua9ZVFUqazLg7Mze+E+x3B9i
7qHIX/Ik9BoOh7+N8VfGbmCRn0OCDWXHjb7iMtI3SZMy7rHxfNvx8MxP6TS5U/ts
zXtoCa+wqGP9k1BtEKbT775X2gqIlfPDvcf0ZMeLc/W3x8sQ3qeDeGacaTnUJiMB
TJB5OQmQBktaPwkBw3blJfyhzAhTNuyTb/sTfNNBQ1N2lP9i5NyNPArB6KJlHRjG
la5hlsC38JN6YGVE8NDTpe3c3o/mrtWokymFlxYMKi4lDgWeuCirJMxTf05izwLu
ndOKiVAk8fYriiPFC0eZsAzv69BnzpXiYp5mMVMKrxyg47spixfI0VFUukh+w1QH
Xhj5HziS6V1VRxQIWmfsx1gAV3lFIqVd/RJ7Nn4MwJGs2nQ6Tx2o6x0wt+rpM+KG
7b0nF7+MNNhtQ3vgvO9fXTfsO8rPtj/0Go/Oi5Hhks+SKPUl4O24fSL3PKxTlNXK
vdOK6S+QApTIl+kjSpxJk35xqv2y9ZAaFa9m3m1cWUcMka2jSbRoIHy9BWT/feph
Mnf7YOF3L87pPF4rS9AceMQc4OuIQ8EvewiB0bCIGqVGwKdkuB06NAoUuY6kEjoF
yrXttMahNIm0Kq82Tg2aL+7XStDfxk0kApiVilNPTL3IfVGCulOXNyT3qTlP/uuE
/eXyB0CpQWOUPnIfuzdODk7EeFaJmoZv3QNat7Zb3kyquLfmFyR7dZQhw14Yiexh
g8f43Qt2Kv3nKeeTVxuTKu1CWVEk12WX3DwK/FjUkJAXWUpGWSN2Zlxc6t186eYr
0Bdgvx+zt+QlKgtP2F5kJMoxoRqCJhk+EjlgmtMF4WOw8L2trTyn2rUR2ajSanj0
X10X9mE7NnmYqpxDVNvhSlcMTXHWmy3VMgUioXzx0S8QPcoQbSJFLHqjNki/CKj4
xpcbJRLJQ2qT87cslKVjy2jH0fRP/dte8/7kYyq/3YYHKXFeARqBBOXiKYmuOhlt
/4P8iquyofoPKaIRxmEa66KgtCf52o8Ynke4ncxKF5fNFRuFuAV21McYTJXCBkDC
OwqxQKuo2WXbpIdjaxHlh4XjDzn9grCqwoxC0FGEhZdulAUuDCft7EXzC7KyRm4W
A+fSWMaRFLYZMbg35xJPZC6X3VmbhaBaHhVD3Ezy4kp7RQDgearzz307RXA+hhss
GZjOgsZFqy4gCf8kVUJUn22slh1+NVH38ebEwl4McuD4LShroG9uqaccbumTJu0b
U7SR7ayDRzhPeJ2vLwEHHGHDXTGuix/FR5JNhpPyOaXWNGvDLIjyc+Wc43lBfrd8
ChLCdR6bRsPaeH3JZEq5QC8LyCl5GvOgYOTAK8lx1LI6NDdQNy/1CPO2qve3SCNy
Qoacx0BLVdXHrwgdmG+md0B/EJfvofmBz60UvltEU5q3krr4gDT1wVYt6QFO1jwN
a7HKTXtun5nqJCpU+E4sVXWCLUDM0dDZZ11zs2UV1ky8ybXPkxAdDJk3LJcey0u5
iKQPxM/OLFnahKigXbM/INZlQAIbvXwMp1u30vELJU2XjXKGMIxX8i9A1iq2EdTL
fP8cWZlxudI3kKmxm/ohhgoCe2X/ycTcvmKpwP3oYuHct3961AndAY7n9A5c2xK6
YBISy/HJ+kF2xomPpz2Z5NCJFYDZGJdRHkrcR9nopyoarHgNFoOPtw9MF1WLZJ8C
8LLakb5XmwceJepbGZfK2+yO+swVprrPQmv+vQA1fgmQ/zgbjXY8IzC6LAK8Z+VV
mv0pA4/bOs8hoswtVBuM2j7HYqc14h1m7yBeZ97jKX2l+UxcbnbLwCBgKQfq1Tvg
gwBI8wqhJkdXRhHif5UwdbxlX3HBWWSuEmVBTQLP0XaOC6SpsDtyQRMlisUv9AZh
2OpBIyr5GUvY8IcvJEINYhEU72zQx1wtTXkXPSBJpGjMMaY4/UbHkx5hnNw4YAi5
uFgDnyV2n2adjcOF2NR8i7mGWe2FEQDGr3SfpVasrB7D5K5Jazkdm5kKgKPHgZyr
llq2evV3WWroQIvB/JOv1FH3Ud2Sbz4DfjRZ/6AZfXc9cNmRyIM37VFOcKzwhcT4
iOUrjZ0B9d7B5Mt8ncicWfzvpWL+LKtMmQK0raNBFfSjDilA93UQrgxSdHIsS933
gZY+qcqMhlHF6PW6/xLzXq+cUSgXVDUy8CY0by8nwU6t2OgaMV8qrVl07uMjHwuS
FTHCYQ9d0bmdiFhYmAg+YrBBxlv911vB8wPJtWMnDSZpb45Sp4oEY0IUXtuUC7/s
23crUm8M670Mj1pxFkfAl3PaBaapPkH8NuiwscDMUutXpQ9ArUgRleCuxxDuWSVV
bvMIx7m8WRja9qKEKyODXOyXzw6XwUVCVNn8vatnePox9txPy5SE5EEVt8ju8xM1
lmbaggN9bBwJJayFbp1ftryaY1HlMZ4lXOmpZi5oGMIE6iR53g4B0+znwTvqhAbE
cyAwNphaOFtCfR8esftIoM1PoD200iMWj3p53j5Pm7fmCCL6SPpsrdtzlXYDOjsb
/zg1gauv+6+Uz+07GNW2jYCI6CaN5DpJ4H+OatVRXLokTVeIlP1pwSIKOhwu8mWz
FcvUzCHihEtxtmY9A/Pg7HCUNfml0OKYVU8VjPY9DItlGSgZPxIJCHPaqBnNekqU
8ElVD+BaUp8ChxGT7U9zv5VUiZ5r3FAZP1pUdOcDpRaYsxEq1b0XoQGgEB250uk6
Xdk7D+bYL5ehIAWyU7YBucS5kjkIcWR5OXIEaED2G0rNG8GJk/J6AejzS/E97yep
xMc28W4Spwf+GcDHwupbWk9QvDh1++2tAHA5oYStSDqWQ8Gz0Pe5zuMttzOnoFbl
H4BpurJcQm/WYGC8y9Q816QRm0dHBcPMk8rCpjZKYtODd+x+YsYAjfv21vQflvh0
yCxpo/JhzONCGDLnYiqyOfHo+WNWnVei+8L4oGHEmL4v81g8wmM//ZArHjN6+Nuf
ms2wj1s8+Bca7QtFogNgP+rTxtBYC6NrWfyaNVGgUm1w4z6GQubtQhAGEgJAHjoG
0M3ECk8mKY0qu7Z60XDrlmJi/z6sPa6Zdq+GMM8F4xHBWX2b0k7bWQW/My6T3m1E
6CZ5YlW+MEOGHN1mEc65lKPp0KeuYaF9mHXoPSUDHc+UJg8DuvQRdcP5b+VhAr6C
l0ZFh2ugaE2icNp/foxOGKW4/Cv9emWbUGE8hDRzHL88YncmWvIo1pr3cZErqq4m
Xeo4Yt0HHq5B7vUilUzp+jBygbaXoaRsm26ylIak3SKe6BhMwWooASPcpbyextVD
AGE1JMVdbAubIfGGqsMpm1zbC+moFtbfE7SZ0UMAX7Ijym/JPf0kJye8AtMvg0Hq
Sgd/JrteZaO3oRYap14bEbVL6Q1YiZzblxpFFDkDfjtPL8dvuoQC0bZdFZlaMKvN
EUq4nLpyx7q9h5SsSwkEG1bjFhUxD4ogtSuaxjiD2QVkzro8/mScFrnN8GcNB8Qm
wV9mSufGXajVfY74iqnXAt0yMMzI6+EfDCmHfTb1Nof2UhocrAWxIW7J2Ep2qO7l
4HbD3o6qnHItOa7g9dzrKKAkUxAySqUBmi5HTXcnpZZ/Ak3jaycZshTc1gLgplbq
IF/YXhOjAPbvFZ2fQSP7ac3cllgWqY6aH4w5uGUN85EcJX/GvGeVePBNH3V1qG1f
l+k3sq77MbGp95uJtOuNjb1qiqDTaABFyxUZ+G5EH4T8unojuHC04pURO4Z4T2Kd
JRIRodNvs2fREKKXmWEVR94u65r2NPDcGrV3L7LcypPGqJU+MJjkB8Lsd7GG8Jvo
7U5esLskDQg27hLNy4kKR4r9xl+TiR9aWfSmvZP+f8qz18SZ7bvGUGoVqYvBBYCW
Qa/bRj1MalcsODf2+m1aTYjIT+HqNitGqgglwsVnuqgC0BCqs2sAZodQ4Ou/zLUw
7CXbKC7SJdwXMBUfIVwPdDLP4qaj8GLJZ3CGGfBJ7/rEMClDgGoGJf/W4PrfgnwG
RFHPaBZV81UeVKA/QnYq0tQVapVFlMAr0JeN+v82QENML2mRWka0+ikhZhbRTxPC
iP4PA4EXTpcoii9FHfeMX/3GoAC5kVcFUxzUepqdujmUEU/sBEx1GodeCO7tR/mE
BVDWChH8ZxE5zpCX34T1Aw3Eq1lQ2XjQOBIf80Nk7WdUhKpY+OSkMf8hrFiOHs9C
8YKdf8T4/1zKXP7U94yfmvI7UfHBBTDXxcllk788gp/dsePtsRC1EGU3RjH6CwC4
tzxJIhWxa7hhlBAbxCCa2yLPU7V43eakT6wcvgzHNmVkXuhEipARDvwvIJeS4ZIb
psvE9GbY5RWxI6wlKaPgqoS19v3/h0W4wWVPJTMm5hu3nio2aUmds8/2MO3K3OGE
ipqlvF2NShjNmX08BWrmC4Z69P3SkM4SnyZSF5aq+4CmLZA/e4zO9PwGc3elw2JI
Ipt4CXScVMH/DgBAivmWYD8lHc/q4gUlIm8hPwFU/9I4TIQNpG893gxWcAG8s7Cs
1T0OtPDmnhsETHnIPZLtCj0vWS0a7OQOGZqMqUY/EOpwfrag/8NCBPImsNzH/eKP
Lh8w2Op/XYD4wpCRRff2Vkp0uH2SD+8BMi+rEqcNwR6eXthq4kCJs+N8GHWjMlmG
SGqjuqAxH3f+dDr1D+z6BRMNDBHNSOycJmkgKx+2AO1UGNOG5ehsYZe5+uhgeQBK
UnK3Kiz4lYt6yJho0HnjQx1uB+8rMoigr4Hzh6Sdh/l/gXbW4lVDLqsY9KgOGwNy
dENTjQtfcctU+paOGU78DAR8yqKatgP2w9jYrFQ/gql7yyRj7ovZ4v6/r+OGg1T0
0lNI6qCSJSePcRg/2CQCDIo4ObsEbaDrR1zudiQlJKmErwqTHlfeSJZ2k74GiWAo
WDxrg0961oA10D2jTn8ANbJJfDgVKylq/RGGwroajxIAv2kMXk40VVmNV6RpnXkS
Xb9vIcR3kXHsW07cVlTTDA5G2+SRee0NQ0d/j7UHtS6bamBR3Gcx3FYCHob079Nq
EHg+QOZofxdNMFSMo3pePX4II1OxEt2e/7RsWqG1yXmg/Zytgns3GjD1TJitfYEx
HQpKW1XVtok87wURkHDa1Xar2dddATiImMbZrY5ulnob3rAuQb0Go4BulnMwJUOV
KdIVP50l+KdOQeR9k2UcevhPXJjv7d91N5VR8QfFWskFCDuQ/eF8asR7aLzEzbPy
t8+lelUbg7IyXAbcJtvniu08GE866sC59ZrvOgUnyGeWcv13x/sjr76426VAmRuv
2cDPyUba8fvzY6LzmrzVtYxE3ea79SHYEvL7XvMEFk2BIaF6L5byknPDfblGoQ7r
a5jmlM+qudoH7x8prhC+tUNcilGNFuLhYbi/KJiD7iXZW724gFK1RQvFFXtnOxRo
YdkyhK0R0+cMgiScf2/Y2lvEHbexX6Z9ZAR7zmbJvm4veCr67a88otzMgCVFD/Xk
I0jbY3Lcmka0Y5+fWOksYH9gRhk7IDOJHzZKBlArZOXwE5+rtc/n+0hNReHhLil9
0y1/yuTbFHro6Z+iqliQLL+P0OibKlWCPr0pSJ8+hZvYqpbt4mvpER2Toht4sMdC
+mS7OtcLrvN/R4FD9lodldDlJS1KSkuHS1SV5TZJQST6+CmMj3umhoIvRUz4/BFZ
kxw/oabXFotWlVWmFdSENobK0urSoyBk+lmndr5+Q10tVFYuv9TcVqZrw61LsSS7
YXMEHed7FjVIKm+PMdXo4MiMmcZgPySHBCkiB9adr+hmHUJcWqnwxXA2dWd8GPQj
ls0twXSb8sGtIUBwTAqQUjIz8BW+bnE5/JEyaQ5RqtjG4FxbIrEs3ItMLDBSMEQL
DcdkTWcPdDdra2tfoXPLUaI7xDJeioEONgROX+I8Z3jOsF1GU9GP1joNxa7lgkDq
WRkAuI7EwlDjnWtLQ9IrSqb842tjwlJBYf6WI1BNk3WLnpESODVbyGMFebnon2mm
+VtQoSUBeC2xeteHiTz+zhejMvjGAsAza9jpMEXkX7YTNMViYI2iXlo7KaLkQbjk
Eb9iEzYzmtTZrhZ6Ij9/Eg+3J2X8bYCHZqv87yBkhKSOHNoLhL5rHOtFvxJaOir8
39ZKLVo09kVu+EC4AfBJMRP2GhKNHE1UeY6TsylvOHwQrBgvOJxtuPzV04MzcCU1
I6BVC/Zo1VQ0uhmQVzegCy3+i100bAWq+ljVd3SD4Pb49V29RkJ2o50l8ffRnSJL
QMSandp6QS8j/1ArK/62zKqPhgxPNNLy7wZgd/38475VeGXl8YqAI13R5fwcxbpi
8htFyFBkbei/6oOmoYKbNxYBtxETqfqYFVbutpeFBl97EtN8pXcyZ41z0u8lIGIJ
pOTFoKNUOXLDGNfSCF+J69bhUqCtNq8o13LnBonvPvrhBWsmYriBH8/uUvXnX1cg
xwoMKpUJ7qqYsOIuT6/e8XTIYnRhYhzXFNFm1sZF9omK7JtwhFJmcH+HuSfatM6l
Nsb/zUnXMX2J5bBZPirs4o090fp1SzrNRUn1cgXSeNBy39MQbjcc/Sy3bvtuLGHN
qmVq0jzgoHn9sctlUn6zqIUCtP98vL5caWhxvj+Qagp6L92NemxrKDxtB2vf1YZd
DnkESiNZS2vEA7CqxKi8P/lNUceqVN2wbYcms5gsgbQ7blM3y01VmPLlSR2z9hi4
MdGhUwgeUByuxSXsvV8LUkg2nJVT3o8U9jUUqhvNem4PzxM61eHgwfO0NYnMDZ8+
L/QXhidpVlO4umCBiunfF6fPd9jg5XAL4TcZE9KxTtXw8gx2zSSIzUGV1yVAJ1Ly
a9w6OBG1QGgpB3kuXHMV0TaIvJDD+B2xldNMo8GhV5cALMraE/9p41ItqIQnF7jd
FZF5VS6Wigu5EmmRh0/aNrx9SpVKcPh1YhCf3sKsmFjuUaYY4/UwZqpw1G9edmWp
dG9Z3nRADngSPjUn1W1YgW5uiNv90Mafmvx3XdrbP3gmLsw2fT07rxRwv4SzwEtu
5pXYJnebIdfVJBKJtZVOwRdi3fLw0cteP1FqwDuUuNpbliUByzGsgLIqlzwvkjiv
ok7ko7SthuJXUBXhrx0u/oMzZldv4ksoSFf5m1f6nnWLSf3tyiLj6daaQscMGrrr
5p64HnJGbK1AAi1F8XmcR7n8xzlSjlaanXj3H5fNSmthjsrYJUNRYt0RQ0B80S8p
zeCvffH038NnX2hjZ3YVeeD9LGRL+1oKPKhO+0D5rYyavevpTtGoFVP/irJFvZoV
aCpmzuB1GIWqOy8o5BoEG0pvYFnIMAdpOIM4l+Qazs8=
`protect END_PROTECTED
