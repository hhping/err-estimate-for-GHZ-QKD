`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9knYu/yqJTIyJrvMw6vJl9MLZslBnJnfoBMmWF8SQTtAtFdVF4GV+9keEflCVdI2
SQD6B/raDnd3BnbZBNPwcHGX+RelV5SDVcOBPJHe4fwLh8fXuElk1iYggjBcoFXm
E9Mu9N2/I6Mz3iCPZLZogu8CKmaXp0ncVwVRH6W3zXNFwsMm2SH8APi9GwawF4D2
WPNfj7Cwdmo3DarqlsTOCVFQT17ZbXgXueN1jyA946QkuEyevyfupT448vr6YB4E
taeRiZ+EFe19ppdDni/BjTZdv3DA8lNBYPTLtqXfMFNmG+i7OPfWBLoXlUSafSCq
da7wTXMADTGbe8nfUQKLnKFxcwKKwjpggEcS0iBiS7uFZ4Dw27onOYPpEIl2f8WG
qvQBh2S2++So1BfQtXFNUzvBqVPYVv4ipWj6sZtR+m8=
`protect END_PROTECTED
