`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SBUp8ntj0NcjpuRBvQ0XvYSStwgelb4QxXN+Y9i4xxc/gQRx1sufhbWAbsWE8BWf
dn/9x1vCQWbXLDpOUd+SxMSG/b5Q3l7pMG7LYGd9sMo1Ykl8BWyZVI6OapggCcn4
laxjdBu495rbX4K31+CwiYkvqg498HhBzrPf1rqJ4BNQTWZhPX3udWZBOTcdyfEb
6s/dAksTsBEz4dqESg4e565Xd4uuBBR16E7ZCibrhNRhsWhlF5bASJ2qFT/Tqn1R
H35OwKE5PFhpQQZptzj5s4t3Z4BtiiqEYm7K+F9cF1U9PEHwHIpx1k2jAKUxUdRq
IYuViOgAisk4/NYf0X+bddy2hOflByxF4rWYPL8yUF22D5LHIgSqeHAEzoua+O5a
ZeUEClrSuplhmHOOwgp5RTM+WJIZIebsbz2TASLiN9nEtcTJCcfiNeh1iy8u9IbV
51rn9Y5HnAYgRnDAiBmjkj06wVU3psnW9T8IwfTA8Ivjupp2nY3jfYxg8xSYYyvh
l4P+SgaO1gMjNETomD2l0INT28EaWBrKV1NMO6Y21MZCEPP3EFFXmkAtwtoIaX+/
DiBsiTxbip5CnGm3qHAdd4zxwYRuSdys8O8C1IGf7j9/shgYkf+EGG3g1/eYndU0
LBipf2BDU9l1aMnWnxysRZcLZBeFc3/2OiTMQeMooeJ5ObdQaa3P8rdEX/NPI024
5/6prhCg/o0EBoQst4nepxfOrfAl2oRciB0JQk3Lly/8e3F9Nx4GU5nfgk8aYkOh
qJ/NXSGLv1LMNZDqJRPN+0+WDnniEp++K6P4RmEHztMfgz+xKjJ663g9G9b7F9NH
F5SGZotF+o2F5j8NBIaLRZnu4VvKw2zD6nLcpWV11ikGOvBBCXUC1A1k3CAFT11t
UPS0/752daqabl/CPZp4qLNF6q6aOGrqFqilF3iCpHpx3c6eDUudbzduX3TOtQ33
RP+Y7TIuq7gAm2Uc5cP+8xxuBbWoLJDwhp8vP53Pud0nA6psQw1EDw0tV/O6RxSY
nCfIRze3fQxCSel1upkQjmReCLvNkQkpY7IyA9V0TckgGj6hFaHugN+BJOK71XLU
AscFJERU/ueqUnh4Cw1jsa/9uLNUO2Z9V/So1DavOZspta+mqAitvLjLvPxdH7sv
0HuWQ2Yi7llOgQ+T2crQEvHbveisgZMaJZSYZfjTaIlTFLZgdmgs3NmX6UOKUded
XLof7s8gCNRVASZk36CTS8rNc1XvCRv86eVPRI7op4Fv000kU9lv8D4DWxR+ar2J
bqxVD+JyTmv5nSRV3ldIK9A8cVCNJNYzmQczShNwG3lqHe4hgTWTwSWemuDesbW8
sjMJZmrkdB/38tHLD65h+Q==
`protect END_PROTECTED
