`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zBrDx2EWT6nj91yzQK39XNWzT3+ECxpDbiiY1Kj8RM9h3p6sHYIH+PfMcEY0aLTB
qNPxqIKYo9oVi1K+rit2xyBVWjNr1Q153vjh75OWwlN/5MrlmLz+BOInC3Q8r8rI
5afDdrILVhqmEATfe898IndMagIZWaiT5BfoTJdrh39wwQwu5ID+xOI/rveYu40T
K/SVevlPT1BdlrPmFfdJqJKilfqN4v5EqTNWKNwRO5pWd4UpJoTyZc21E/6bweu2
r+JwrxrnC/ID39mqYlz3t6fQ8un5ZcIEkhAj+W4GqpcXhIL2yp8rst6YO0WIxr+g
6Yk5cDbzZ8Ob+jTOmivI4CFOTLukJKPU8uIlnQXyw3rUmQpLZhe2b3B+/hWADm9e
Z3lAodsPyz4EcsIOs0s6BsT+aW7t/VIACtdCSkKSzBLgms6uvj3GzPC1t2kKvl7q
LP13usOFbJLGCQdq2BxmlZNMXbC7nJP3paead3ivnsVSWNi/KIF6oUoJBtu2XTSO
ZLyyeNBHByxE6HzwrZCh0OyoD+W0uppiMokLI7HEII1ELHo0lv3mTQVJIK9pV0OQ
HwtKYtv8LZP+YoyYq7d3nllOyR8e/QTdKj1LXlV1XbXS47aIFHWsQwo76WMMtrRc
cZylApUxUKq65qogmriEMJEooZw0DdwFPsTfm+DrpvhbEHWDQbBCqwUMgO+ji4/2
tdsBvt/fqqzWZRUl74sCOVNmqACJsrzkTAas1PVViGo2NWw1UTAJYLmwXwimT97d
1Ap0q0FzvSVbygm7lySxwwQ7xzYllwGbkWtKPFi2tF8x5hI1avTKl6ju17CSP3qm
7lJMHkrwOb24idZAMdJR0At/1URvnBxe6P0xtZY9DOAyNlTwRGGQDBwJli1eRzRV
ywaDgqeAFB0QzRvSON+pagFKYIQrdW/niVS1Vg1simLpSVwDSxscWGkpTKZE3sFc
eClN332SQXwV9HD7z4XCdJEPl5/jPLCBG6bDSoJH4ROKWpueWoTD0svnMwbyG5yA
1SQjGvxbBJAhRokRWmeT5fEqLZWrcgN1JJC9KpjOCzhB++XDqgZ2l1jkFROSqh5d
pz1ttf/E/oIrIyjxx6x1Ck9yHxMqA3vxr7bQPCms+vJ75xXsrMEMo/N7nRDtX6xs
WfpW7Z4K6wo9NlskzYbtQDaJ8AVLyYR321uYzrPM927+fCscHZPXphTMVfP2XVZo
ALoAZcEAUbcY/Wzg99cQB5zD5LNvmMQ40lo2TzlxmI+11aqc6lBi52qgPJ+daZkk
cLF6rsI3N30wO+MYwF922A==
`protect END_PROTECTED
