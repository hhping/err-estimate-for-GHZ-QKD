`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tJET1dHkogM5hIrbGAICaSWTod75kJ/gRW20XIEtDHhPeu5VrbXeitx1OJKVNZ5m
sq7ImTi3WjiT3zlM1XqblixwERG/8G7YB/QXI1iS0xtSelkAnfB1hSy8+8XeZXUO
50vYzuDib2UbmJjGN8MUZfysTjDAWO5YXEOk54dZ5FlxE0xFtOrXnzpUOy0D4iiY
Y3CpPo+nyfeQV4uF2eG9tB12+RgB5epdzCUStW3jZcJNQfnXZMsRQ9KAa/Q0XoMo
xqqCeB9uBVUe6QsBQA9zOKUxYfl4j3je6UImQTpA7XxcusL9vmMnt5VKInhTSkHr
0x83U8KWnqubg5yTLmEP5xE0F8ZFxjuWgZbsVDGob8roUnBEIxFC2+E3/ZgnSrdX
+YCq1fRhi209Jneu25Vai5/sWIWmQi3Qw8lqAecdVOnYZ8CKC6luk098NCO1/9Ct
iwIWarl01DEctpAN3HJkbmMUi2b8es77D7/jyTsTqUp/bpO3XPeWq+8bvRf7CJ7w
suHGcN6rWuJ6KZUcwjB2tzS0QckvPa0YKANvq/Lr0FLNjNlL3zpQ9kWmAnVd+m73
L4oNQhpWI8Mkrqpt3LK+FxrjfHSADcc+hQD6VsJ8Zr46fazaL5cbi7qZ6PR2rVAd
Ju1XTm2h9EUixV5cyYu4Vkw3CzYLbxjTvxboK+jN43x02V8G8wQGMOclNmB5A7aj
UE1NVwk184LT0b9unSTQ+aQ9NGvpoXsIihEAKdL85yOR9Vg9PL/8O3Xbq2d7QUPT
fCtLqYpCk6WkcqAV60N9OcIYRvM7qopKrNjsvHbF+UFGZ0jwSmFkm8C7fG/MO8XP
5HE6olrXTV3lmUrRS1m9EohH3bkwNuSauTbT8v2jpn18nGtPM7UIt2ecGbhijROF
QrD08VKgW017yadLAGfBlwnnC6PQ2+6o+xqi7drWqaTU53mY34K1+RqFpPHlylt9
kqOqUtU/L1Ta97NFnbcUm8wiyJJwHbh8JAXydxbX0uuU4MQP9p52OM0I4d4Q1s3a
kYdAO+LTaBEFwZG6LrfGJ1CHpz/AgC0LNXHUcwlaL2dh3zgh8tpYwtVSZp2K7llq
ifpLGpRjJuljKg6CPzBccn8E/Zy6JnCE48WqPh8AoE/yRgE2ydIdHnabeGH0FkNk
zhIBlvNUiwiBVxkxVS5bXyl/XpN1R8S2wdaeFOBiQuupZFGaRXBNyNWh8n3nJlsF
aVcRCW7XHn4ULHkK2MUy38TU2JmtimGBZ/d1VlQEgpZgA/A+G9aao99UsmeDIjAC
HP7EFmfEYhHgilb0EQr844gMTUsdtb61SMRTMzGHrmmmNe76ooTsbfh7ArJS5E34
aXDrG6kFfOqfiYVAPmmcbOtMJHkKyGhnBpBLq8rL3YsfUnGZOyziG9oTfqY7ua3F
Mr5DQn52SV9VM0r62k8Gmg80Vct0oqAnKF0H9zHyM3cwz6zij919zjumjpzi94Mz
vG2ShOiQF/gJ6cNr+x658MvU/f0XMCugiQ3ujEktCWx4Bgs6pQYRWBYf82NmHB2c
eBA2UPmEDGZvYea6HhjDlfstSqTqqsoNFhC4giJNGfUw3TrWMZLbJtd4svKYsFY2
/qZrdGMCl0tnu8uoJ0wLGQ2w3HTb3zfZOzgsmr72ipKCsUWKA3/CdkYUljD3XUOQ
IomAL8YzrIY1QSC/YUEBvhhARjkpNWDdYMpBilgDclQXfIJbj+EesV15ZiFXYokt
QEZV1l/7sG3LO2Ep6yrfFbKtISIQCAhckWVj3vhCX1uYw9LKdPpCKQwI7Gfe3RIx
X+RWsu0eiS2t76f0lflRYr4z6BNGQ9sSIzVtSuB3Rz6SHKREL3IrKLjRVqGIDMe+
FTonD3MsZKr73KeoA/RgvJ4WEDjjkSiBNQ6gY+yXL/frNX2i3bi1VREVwzeeV76d
2hmeAimX2mQNM9VsDVDFifR1IvvIFJCcmuqhPyrjRRntgHTxRp8XBU5DYW4SqsNs
3NI7ETQ3R88DaI2hYiiHtur9U1mL1x1cBHilCKGylWFLu+iLPbGVhWLs+WQp5o8i
5/pP8jRy4VyO5lVA/c6Vu43uuLtXDXUdv3rPmW/YjyzonPEeOXU7kpFLEWjyTk0Q
okxL83qhwDQLDE6Uvbg1f+QxL1XVJRfc7hP2nRLSKnIvYWxgzxGf1CuftzLLHz5U
eKTbPa3J1ORDN//sekTWvTb4zQTkAVmA8t5UoPDBdZtEMih5QVsISLaeUcYlhSfs
GvCy7UlsuT3DRnXdvdGu+58jzivijFMgLt5KhnJ7RJ03NHUOu+Ldwr9crSA804tA
oxaob7y20HLCr36HOm3YMTYr/+G1uE99en75MkHbNT+e+VQEh2RLDe7ioX8e59ga
4M3PNphnnQ4H1IzGts9IBaCgnznblK5/LLBP+PTl24Lo3p597dmZm+fpdkFmko+/
5VxRMMrMRnCQ9dJ0/6q9IOP1kad0OgNf6h9wD/1s8TwstuELmZxvBwHkTKca4/J5
UfVsoiSTSMOtn3eXOSmhqANI7fH8H/dlsYWMUGqMSPgX5Htn0k9ZKtvBIoSDF6D5
A1oVN5LFlmzXNPQmwWHyC/WxBLjYs0FqMbLNRBcSW23YbKRuBfkDizioati7dR9a
wSrz3+KVx3KBRKGTBHlYyng5rh+vDCIyoIFavxqEgJA67IdANvy2YXZY1m2e0Ped
qkU/2FMI45HPQnUYCp+p7MmO+u7KJxdTxAi8mSL1+DOWLpbN0l//98dCKXwm2yUU
VeWiZQtSBhC3CS6uMKAehFp0uKNyKYIM/zr22SOiQwtd4ylXgPD2dj7brYIRI2ay
IyyPP/H453MAPJyq+hk39uyszFWeK1mHrKe1Ff1oBeeftgZMypKRLvMd5Aoz5SoG
pufB8UOhc/s9BlrqgNFs/v+fF7FYXWNa18MbzZxoFD6dh8GIuvJr3KvcRqsaT2cz
7YqhSeRRcSwmq+ns3felcWdNWNwt5YqwGaaHj2Et3Z4ijkYqAUzCB/Nhu65dIxxa
W/O1ZFCvJrDqytibt5EqgaH9O0SUanJP4OAMeSb2D26lYI+53b90NJ/j/CP7ttwD
X+ZZO6GSIMrSTzv/7nFY4qcP7x+7klww04JCjAndIog2lNhwG15NCC39rj7OhY/E
kOcE9veJeJlgCV0T70Z2JO6vagfFxiB1whzwh+hNtU4=
`protect END_PROTECTED
