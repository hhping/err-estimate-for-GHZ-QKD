`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ThqWFYSlPWgixfbYhF8VlOPBVOvfHXIabn/Xhkl/gOBvvepQCez4CmojllRNvPxY
4jHZ6BQ2oyisQjgpOHmfzl6VmgZ1h53UZC7UKrz/DHwAXmbCZKLNenxsPuT87K4I
ZGtv4TmTl2MXUoXIoi9AAV5/9HcTkbJIuHSBEBGrAt8sGpZUPerK3R9lEoTTrIY2
xqfAo+v7LoLAl3CY5m+EwkU+zr5msszrrHMB6Av8eX+VPkJko+soCmqiskI/xC9h
ETcZ89JfLNRQs0jQlETF/nepLm+U6zx3uHNRoAQ28JoBhV7YtvDavE2MUv6/V0I5
wqWN78SKSFulBh+MbGOynnaITWljUy1Ci9uqYuL8hl/WWno5I+dwpDCtNenQEQDi
G5ks7uv9E3ZKuUnOWwxvalHN9WjAmnIlLN7Y0M/SzRrRSJWNe6AaDE7B46FS1DiB
30vYsLHhjrhdUfBPM4FHowMDW30sWBOCXPa7qv3tgEAENjfW6F3ewCztTCJUuq4/
GOeQXG7EX6qzsPSAtmB/ogzuGpHIf+ngbkC3Zk/7yc/rRNuL4phgyy3AVTrggIu3
`protect END_PROTECTED
