`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TdLX6PjFo+HR8Wo/6ykphfymE/1ZdF77xEIso03cm73MOn3+tTnPnUbW5/vO8PkJ
C7QtPPDYMennAnUqioUkBx/rI/CY2mAmXSle3YMcZJJtgOexBxpvbMgNlRYsupi/
SLsKZeRSsfUcW1aDnzmpwfB3P1ZC9UeC0SH/q7lz8avERSpdVOfcLhctXRIZlkSm
zualsnVO8OTbXBhqVgkTpp1JmYd5bbchCoO9tIdELN5v4l1Y6zf/y2Lv8V0CnfAj
mbxlV0jyiy/YYYwaMoFWg98qdTQKGOJf/T8LFVmzfqt7RAhrRhq2sVg0Kq8/0XGA
jP4Z4AzH1f1q2dQCVep5jWFDO2Yf21juI/SGUA0Q/Up4iCkl29cTmfSu5bzE7Bw5
VS3n/33hWS0UskSCuko37GCOF15z5U83rHaIu2wDhuTAbqk9LZQLIt1auNZmB4wO
rg3SqRiDetN8wfJyo5C6TDnhbPsxhdKknfM4QMNHiC43Nghv0aVWRUwE83K7sEN9
HXrN2Ynat+2e1UxO67O+OFA5VU2U90MqfR6mT4WhOeQOIj4v4dUeSA/kH0av4RhT
h26QRnZW7jnE3K6xSTuJDrVRoFSdhEVttBgXi8d/a/32igUboIUkX11f9s3UzU85
78IHng6Rc8tang67+vEvr9CnVH2U09CNpGup8RWboUjWd7Nr8ct05D47JI8HUZzh
TcsZpUCngjuTH9CAXS9LghZYojt+cVpbzcAUjdzulR7n5V8EL+HHCixQyy8itlFs
BYBPVArma09dpOqV03H+sYRYNsiuosP3CIm1pYt9C3t/o+P5vFBIkH86g9SPe0XI
dTpgG7ivOgMLXunM+dZWSjujM2EO5k0lPwsJL7mmnAjBr1rNQf5FY5HL67a7b+ul
1LZ159FJwXvftBNP8us+SVDggAPK0BKX42jpRaEDWe3J/rKOMFmdu8ElP3JATydI
53FZ6PGErncPxyD0afQM/LsElZ0/T90KR4Wx1W1sjrTkmgSE0JJwwgULdOhrYjUk
++Awf+7WOJKvEpzv5C3a+nnX3HJsWgFYp30r+GUjKjQWWIoyavLJn4CEhd6lAd24
/lGj7DYpghrqD2h2NFi5NcuPH7sul7XOHCp9lG24P5FE97JEbmrC8hu2VWZI/nRP
YjsTgdZrjqDhFr1YD+vpenXGsovds9Qpng7+X1YCNxPKwQKvgo8bJxHejdnknP6C
n8aLOAi3s63QeM5uR5/A4JaYTuDMO4bSLHzrKqcbk3pJUb+oqsIxaNUH2YdC86JK
S6LDj+hX9EAPc1f0R+EfYQtoqGmCxF/6cPaj56EDUXT4FzkcqBNoE6MAxZj08YKq
pioIkhl8NHQ2uQS9/39z8t1gyRnTnOu0C2P4+YvoLxFKbNR21BC2KspM6+F4jOXQ
qHc6K7UGI9V/xI+09WjCgl1nWq3W0trJuVN1uLVut3sVIvJZO0phHN5XUeIsi9Y/
SiArta1mtbZvRtSPnlznUxrYg2TRONvLyQFoFfmCIFgqjcFpemFN+ipFutglCfoF
Ve1Y7FXN7tJL3CikXWObqlbiZp5y5IYwcjcfEeCBlpnaxI6H9TmfURS5KYHeg9LU
3At1bAEgsFszQEEcSi+S+2Zmp2HysttZRYIASB5Tk/sZp7dlmECRKQyg7JtJ/LeM
Q2YiXj9sUhaHsS2kAGxfDilS0nCRq+GsL/g2b5xY8DvV+ZCpx4At8e2zRzrc3cVX
52fxLTz1MDATiAZfxPuZ8UGBJdw1zKP1YtgQKPpnPevHgovToK2V75vjt8LIO6TN
66Qpujg0EeX8dH+nqs7JRLNrv6pE7gvwgICG1MrgAE9DHBa6omVV5CfXM+Ly2Rgs
JchncfRMdodpuCpNPVUXqdwLHo/mQWi8dGvyAXl/Fb4HB9uBjkM+Xp7XVPIbNg1r
+M1CdpWfbk/WB5GDBFWklWdj/WeRFE6x5kMVoI/OUWl5NqceoABKERgBXIA+B0aL
zVB2dc1eqv4nrylScLKpsxauQVM7+i0tEw1ZiEo6pZxK5baond4LnI7cnEtqqUQ1
9B22oKvMDbo6F0rh4yLq+2Wlo+sJN9XrxZ8PYHTyJsERApQZkbMB5fJYvoUGkx2a
kFM/K0Rz4lafNOevCZZlyZMBJTr3WL6RqOOPx6IhAYtE9kDHP56Pjz6npcWGpT+P
MmPu0qZyrflyCgr41jfymF0s6GtR49RLpM7DgQm73uZhXII2QKvhR1NwHH1rShDD
TJDm8PGUG9w4dSLK0cvMFM/7ZNhFRzYsEmGXhp2cBswTOgYUx6ba+3xRkqhp3sXe
K8HXnTqoj0RYjEE5wHdZCesHJxcLNEvSrTFEW8/nTdqc/YzLLUohlUDY3nSNr5nx
E4VxwKfhoz+uLQ03wUquQxyvXUvknN9mOuLxDm1ZIp951SUtnS/K6D4e1F9xjKpz
2AHQm3ocCQY81c+1erg3bLVYDd1qR3ISKWz/5bBKtLywvQPGuZmmayOQHP/usi2i
bJWTI4UVuZvAhwEZZR46yP0akrFPd+21tC0Fg9k57qeHJZorKmjHxswgsUiR+7qi
ZGDO2A7qnVdRKcNPr7Ez0cgw/OqS78xKj19zOOvnj8Pqz7SOpsGZIbhrkAkDSPCa
88blYHoh04ORFvS3YOCudp0nIoOQgzEOr3cxclhB1kMuVyDhnPHIfK5L/f6IhmWG
yqFXdSW0Kkf7JolrzgmYEwD3gWsNIaLYIV3mjUUw2Mgd4OLCEObgzIRNvb5+c9q3
jsdfwAjx1/aso/zNPAqxE0USS/iuKHVhnAaLriRvEEm0CpQlmY9pHB4vvQ5jUUUX
ThuZo9GaTmQMKpKfjUK5/aBMn4PmQvhfuSpFJ0TkgFFTSkssUmeOXEO1FRrr76+U
dH5WIO475gkF6/sXUD3vnkz+pMmtXPLWWNN4B2sFK66OGzS9RCyhTIZUzP/fC5Zt
EFOZaUOFor+nuOs8xr44AlFXXJvZ9GtrnMCUi1g/ryZzuqJ7eONJCGxAPF72VErq
rxcZsKQ4fqhUuHMwWTvfpNGFrEdHaNzhB3QGr/mE0W9R4x4LI3+fqeEMi+ESdqCD
7l0o7ccBulDu5+L4AYlPXKGwTB4qLSmP3SXRpNMYFPK49qPKd/HKehO/K82wQ1F+
C2BQSwMwZGZ7K3UIO4X/c3OoU9ipj4CbdmVEdKlPv5umqD56sYACEGrPVu76epUp
onAbQWBSaxNgMmuPXrnTzf06hOKDzCUo74Er287FBk9Qsw62TiZ9l7xtHuS++hko
G0v/zez5Z/Chpws8D/kqwH5J15ooSBxEjQeJBmPP84qcW5dHPtq+/+tBAzH9T2iW
OZB/OGyfmb/KssWCXwIPoaXJSc3oARpVerdleh281HO/eOmOBAfJ2TFuMwBORSva
cHlL2jhBF3niNbDRSKE3GrqsnvZkPts/ElilBEOdJdcm9EfOvI0sJ+HjZ8MtqpX7
eqsc3hsVpSCylb0kacx2WlG/PpUnbB6EuzObtUAqqbuy1TSdtIDgdbevlVxRaIqv
20nk/iVAQJgQ4HOdIuK/DXiVQtJ6TlujsDDYcMb1nkbFSmrXy1jALCbmLk75joBb
RQKaiNcnMCrjHDi2sBUZigfnEBqkpcMZPAiE7RqeXBvbYVs5G4r3WkL6xrT3unNy
KjCBe5U9v0UwnGmQr+jk8y4ZTLGLcib7HGodRnzFXaUX0U9+xfr38XJADc5cxq6G
XAIKr2+SXqp7DHy6F1YP6aAeuy+lf8MNGfWatXvD3vW4vqXx1wDlzBS76sWkU24z
XlhdVtLaFtdXFjltzrDbISKHN1FSjVO3FoOTAOm6JHzyaOPhOGG6/78TBF+3yIXV
V7+LT9TW6WXSZaYmTIavse+RHnG7YU69sEWGBMMau2iXCxT6skOvFyfuzWYBfGE7
hDLkwO9xwPlKkentuCceWP9/odRnpsSqtEE3VRFGCyUcKvSRiCBZhl45Xr9V+2Qq
vxTHOkTqpexWE/EOjZrIVcgHc4ZdY6oqXQ3DhHAjhYG7drY7qvCjo5/Krgod41jJ
Qkz4CThhNrLrAzMcS7s+eU5Ndddt31WSnZs8ciRYS3rmnY/MptOSxftLeaG8sIJL
J3JIfpPGp7LU84jRmaLv+1RUMwdvUEnzEyUt4ZdnC+PRBe/Z34LA6x9jLjgfNpVJ
e3cWHvBKXQ++s3MosXlU7Fh+x79zu10EkgjtwrulHaxDA0Xb/DHDyqDZL5SYogow
IA/PqGVAPF+wvjSn6WjaRCOt0n9buy0wlYFPe+CQiEJ3NTnq1rr5ukhug0dT5/vz
tpMUtM4B2KRFg/Gd11LmS92qyarlJ7PcKbXtYIbRLlWKndpZZvE9pd3r95VjW2TC
HXlgdOpfgrpEelWs6Ht4EXOD1+kju9RzntxD8yIBcweFHFFqIWbpU1thfhb49Xg0
ZqeykuXvYyClJFOs+kVYxbC1I/rlZX3VyJ6MHczu4BviqBZ7pk90jbiKOexyhPQd
GeYZ9hYikvLfHXIfB0Sks9N430aw/Vujkrk3F0PlELyLFe0yxlLoq+7PbRqxuU9K
eiko3s4LsD3tJ386sxmV3K2jhY+6mt+J00DVamEam2kXZDlAO0GUne3bEjv3RhmA
NcD9sT21HMo+0lmpg6B8v1DMA+g4srnHnoswv0ikP0pu9MMb64ujYuViDSZa4mXV
spw/+qRKLT6+Cz0r/18Sk8yZly+eyCvT36lRnffy3+agg25Nqm6Xb5PTuPGcYQVT
mNbh+o+wJcduRRcx7GBOcOx6tRkX3agRk9w3TukhecG8PliLSgfjxWOVBrU+RI/k
H9zJTu5sOUQrqKhaB51cIydvyq7FjyNZMF+mPoTrHngUhLUwg4gNf7UAyJbfD/+y
gx1IktGDrdoHLZ4uTtguLQSg+WRSbvJQIXEEq4c1H8Zf1+QlRj5xyCbueg0cGJ+S
KaQZjmd1yzB/GdrXArSSZ/mcXkOBcXyAs4eYQhQN+RaWhpZKUTD+vZEi3dPFuVkn
OyA3kMXVS8+F0fjo2Ka7EKwtT1vypfHnJjIslUwJ8NxNL/nECqE+cuqY8YMqSTe5
EvszJSfF2uaCQoa5KFhDDvkgvGcb69Awbf58KDCQVJCI9dGpXEn6Iwhz6zkFfAZq
GvZTcE/luPHwSaDqNs1WZigDMzlZ/0aX29RRGZOeRAoeffWrgBe4RRK0GTkIYl06
3GsX5HwWY8vZEE416rS9/kbjw2vbSlIHNEgKl7HGunHmgLpHdRHnuj+3kZFAD9l8
ozv6KD+I/zTeuxN8B0ffA3fbBETUkustNNK/RdjP8x3kTKEH9BPD2ACv5EUvl1ZT
kcJAERkidzes2ryDl+WNWcrjyTsieTN4ti3ZEljKtjxFKQ49W7CJYWlC1vVIB+H3
2J/xOn8yZMEB+IpD9qTc3JHAoZxFeP11LWDQqQHAXWxqJiLRaICkIEY9G090PppR
qjUXcce6AhXWreycrwXxnkPuzVKFmPKTBPJmLsDic3NgOh5Rj44nkrC71FCCaIgZ
7Wd6bmJkZ906RdpoObB/rjOzTJIPCx7o3QuqOBRaUvO8UclSLPrGKeiGiuGpKaCY
2l+YjmkFdraPYX+yix/jw8ayHMyB7x5IOeLE4IJQLsnRfSiAhljAdmemAR6zshWc
3xuJT1vGKM6cr+LQex8itY5tI5NpMpsRwRO8zT7fiBKXuk0FJmB83IIGUYDAmeZx
YVNiX+yt2TCOPJR1LWrN5FpUHpOZ8jEC0705RP/waZQ/V0spmYJXjf661aNhLqHv
LmuhwP8VBAm4tHXRNzr2g/cnO/RZ1nm/ImgRGiwZehfRs0IGZV5y9BiQNQCCbxSI
iIkGEPrfvSGYYUJ440uXJXraLX6nOXFh5Q20VSq2QeLBuBI/4AIORmxTgsUnyLww
7FhNX443WGZY4FhilJ6Y+Im3flEzahsemvGFJa+ci+URdEtBnhoEf8mgpSURI16r
JhUYjFcgksctwsIMe7orSNKKB4+f/Pd7PXZo50N8fHsiI9bGZwYmh8bHoAJTj70A
oKzK3ytFimK4mgeg44/PCftjTQe15uzkHxLPMWlJo+Mrw4fZ+hZ9gXodJyXyTS7Q
Sqy5FgMHijpjP+UWdKbLGNBn1PIzqytGVKsind2zGOkuu4CIaQAZ/CdioObWUiE3
I0ZLcdC0/mds/oAuKlgGJ3WSXCt+SsvByGS1Zfk08928LbkbaeYJIDns9hOCKorf
GrGTL1+VBbe93qyI6/mU9iPQk8bLlxWkGd/D1X61Liv+JmyWFPw+rxEMO94/FptV
6ZmlO7I4YLzBL7lATEsECHrgwO/oSkhAVS6fPkD8R3nqv3mxhbkpAxtSMm/zRuKf
gN6ddy04klg71AXCgDyTAjkxTxn9eb4lSzRdsiCxKD5HUCGZHAaYrG1ExRTVY+fC
2V4OSKXWfa8APUQhulfbZg+i9bQeafQNiM0Ey678Yd+3wkVJwbbn/YCv9O9CESsY
iVe/9wBWkuXTTdxxt97c8A/cZGu0QrlrI6yIuRhrlV0Kq3/mjUU8jihCnKbpxkPh
mKOhyF2jXFhmpJsm/pRXs+6qAigT29YEDQTvUdXKgpvc4baOLIsva2Ta64BFtli6
K7SwXABdFIewLN8nH8bg3BHh8XXKRp0PBA89JKW//9WIGMcPTk1WtX7AqtJT94nX
QgvZPwNJBwKFEyqXXwXO1E/EAk+ZfvUqIzmZBCMacPtKrKX23qbIebU68aDkI0eS
jzlfH4jpZsGuSqc5nSxTjH1rdQ1FCdTHaSnWaRJvMw+PmRbu3gx8Lh7MWj2ECz5Z
6POKkrM34tXl35Nyt1xP64BHLFLdni+t/OHUo1j4mQE4nMEh0uAu215JqXoFSJ+b
APeYCpZ7HRdq3aBIQv+LifuoyG1mxScMXa+m+1ea7Q89K45Gk0s+uV94NEYyhmh2
BBGIWYg5ndY6yUvGhuluJCyPhGIw0FcljhdioCJcW+ByoU8mfzjFUd1mtAFCJTZ5
exL/kNtbDhwkU+/6UmZh6PfQ0D4+stqZZ8kZusnmMSCimOsW9Dci4mRNpUXStJOf
d5QBU+2/SA0p4iPsm3VUjFXVVdfdpmeu7QWpEMgxlMGo4dBYBCd9vwwjLLTf7qOq
M599pTiUCeHB303iA6NRoTtJVsEHgmboz+GOJPrTmVFXFS7Xb2LvHNR4R+KeGGBk
1zLlNALZ9hkVnsk4oqsjzeu0dr8nArcRSkkDKJ34lWKYiEGll87RTuqTqGfaW0kC
4vrofGIwPRR9AoSyCtTQ9y9bhg2OlhzGWwK07W9pOgczOzNuOLY74vnLXFGFKw+J
Vyu3p7NGAJ0Ia/2lS/rzvvmLRwKf97brHRvItZzyFbJlQ4B55ab5KkSKOd6zE14N
xm7MAmOuivRgSR71ldaUvoYK71HpdTmLiFBDHPttcAVpeViaZS4pEqEzyd+dSPjF
MkzUFDYS8bSb6WG1oHzxaD94K3dmZCxJ3AQb7B95s+p42QJYf1pno/2i6rfP6ger
M7cgPLE55HY3iDgy3Nungw2ybAtO+eK+H+yxv/TwdKQiUgLoRBmL8ubd/FpUSrop
aIH7MqRm4of3+p7pNX/MM5qiwLQVbt5plV4ZJO5ztIk3N3e5ZYeCGHMBfg9lOFjZ
jp/F9Nmh8YcKF2nNtGEpjClk32S/vQruiPMjqWg8jsS0uvQq+8NQVQffWAnZ7END
BmgUF6JqJll5U+KOgjw37OXBrBl373S7NzkO5D19tnVFSfHLAW7q7xchRNj1RnCH
dhIXkfwh/ZTq+NBqWXQPQ6egWFAPA5qqZq3n5dR+Ytexyp/J1ztnXqBy2QM5q23x
ppCuXmkiQ7WEeYR5S63bGF2ZJ3qAxOfZzchkKP/R2l5BM3rLa3PCsa//0EaHMpvc
TdDps4hsNBgacU0T+wUXoO4SAFC8r3B5P3EB+0Jct65o1KZBTwaMuzCLkHsPg9V9
ZBl2yCmOgH6pdqo3Nnqo/Ihqd5IMLnKXgsJHfjiPeiUNPI2T+nbjQkqkRCX7Bbq7
Am7C8Mh1vniibhRtcA1utxE+WRaI3BTYxcIXnKTaTYal5mg+tH/bvIOGRkQYjGOA
5YikbkcTdmXSSZtAIaDxePj+0y9k7oUgyPVkpuZajKnkbRmujCWXmgAcOEDoI4U9
puGdpnEWXifgUTQOoFrw7KV0ZK27Bcb9lyYEI+r5K+hleX7aW+6gPWeIdoYMdveL
4AEhlwUt1aDKtf9IJTWR/FC2gzzhHMq8rhVZkc63gtixQSkpQBnzAWqukkWIThoM
C7JaAOq9UVvQMwu6xx5ELwPx979ni3TTJHiHcQooOLRfuZP5v/PtA0CuDkcSrPYC
5vyNZv5C/kve4FR+vx+H7NRPFCUDIVCvuahmT/aMpqofjPkBCpwvSP7K/GlszPGP
au2A7N7degfbbJKVC1qr3w34d8GEbkiLuntWovRWtP/i8ROsk3i5LdqW70Laluqw
bOFIdMcnv8eJpwxPXsx0YAjRkJJj4EXg+ZkKHx5BwzXXavz4D+QQIzhmekeTkVrO
P8Y6/tUoe96FWmzUzr0EwIe+1nwI+IOnmxqXkPs5AitKmv1pxmWFBHnZPWSKMQqJ
kaL2ndBwWP4TDPelupuSGfJRU+chdFOPhivEFSw30HH3qp+VZNys/Dk4hfNrMwjZ
0VLVpGUOhRxRlRgzxB9RwrkL0Ez3Ixnhez9q4u5BJusq2OO7kupZTe0z4ucPUVmJ
d8TKEtyhebgojBXgd+uQz8014VZflj5BtdfdjRRvFmWFvazhj4ebg67RjMtK6GyN
TL7s6QFwxttODvw3yqb3VNddqfOyL1QD4TLwbvYyS0eavSj+kzgJHEsgKqliRXAp
0ke/VHFYA9RKzBwlC22ER80/YPQqpXuC5MOIQ30DjsiLFO+vfXVZjHP0ylVPV3Wi
U6Zi23URYY/S0naGm5fDj0fiBPX7wn0KnMZ9ulzyDbVa8CoHVkeFaO7pfrtjENyZ
2Lx49b0X92EsgO99WJ+ccyxqjxc9fTO0FvjmiBEG9dj7q/J7i3QwLpRXJlS+TvvR
H8BX3+4BI8SOMg15dNw/tSyHam6nYs5e8fwAKf7kfQF5cSM9ofUmCCq55Bi9vaB1
mx2vsEmzaqEtgEf9avX2oy7hEyIL3lOosHlHBbaWUEFnsf/SixxMF7lzL23pJYPq
7AvavBmZClW9JfmrZWzA2MfQgG2P1HLwIkp8W2fMx0M4a17xNT/i+CZxJSfeDXMu
dCDTHtfx5RdvpRedyyAWA2gIIqUOeLtKffvNxgsaGULN3i+qaqhpBgtL4haTfQrF
aK9Fp8rmxA+P84kYKT3TAy0kczKxyrxYnPr9f7rCOh6fR4JhKDW047e6VV7agdVI
JDQcDhJPCLDJe50F7mMw0gKwTtSz+NFo+bLD/8sgR45ZNOX7KXTRkZHXsn127arn
SdpX9WQMlsDn/7/6Xic1mmphLPaFZo92STjKyeiCvt55q2hI8jEQgVqvo6VNOuHL
LLxScbQDadedQef4BU6eMaQK3BCAnuVqdpobFo43229A/YYnU2ST0nFQ2pA7TzMm
IjR0xxvNMXMgQ5vNcJAdvD0nVmXrWdXy3iKQdEhKhmJTX1Et9kfet91Xk0dFtHIi
04zx5DMdJ1tKVK29Hf+WGybapPtYU8e69FDT2l8rCSlOpyaPPrDXTZio7TrXtCvz
QVWc12/u2+5hS/uVGHBAcWfSffgfz4/B2VmfRAYJ4uwqKaErP+bPApKr5DlUQ0F2
ymK1MBrXMhdz31SZ56qeg91vwT9pXjliGssYyYQ5i59ND+f8cqyhpeU6H2ZFAPdm
zy1y3quMtVPNVqRkW9tb+pchFaxaqkf5jlFXWx+R0sdcinU0aZiJAOOmsg8R/cRp
/TcXEhLDEuA6NCITP5eQZvMsQZZ7ZgwpB4Sf0UGB5YxA9eB4yC42AGWG/8IMnOD/
5GugCb+iailG3VL8ZmNeZU7pI/hcx3Y+TBTuSOGWP4Kho4Pfojv6nXXqRQj0195G
RuITjgGpn4Wt/JIaXfU0rGvoZ0JTuFsh2j3Ur3/D5IICMJJSgMB+tJSBXxvmwo0S
sXPG0yDyIIwyQ15uA+7uFdiBay288+mNjy7OK28cWpj7CnB1iFbN9CwUB/EvImkx
T+rc5uHLQ44iTrSh+OUm56bIx9WVmT4Xs1YZ4wO6m5dXgX9deWyHQEclU9lPe69w
NH8m8uMWQc0vJmUI7JIi1qRYCVteEl05Dqsq3tbcgSXmqE96Ytacuf4Y0jdGSMEa
GWVXH4JOBUaJLRq9y6YMYkNr+ubEQs1wonyLn87j1bee6Hq9I6TOb2fQkMHCLVmg
+x8hBOwu2xer9At/RONPTtLMoWbB9RGgsI0fHyTNieDWujx6wpVfkdvRGePeC8Sj
61Dhqk28Q1gFnkniiGTygRLx7zz958Bv1qyBlSSakv0oEMgfBAm5dGRJ+ep6s6An
jwvdT2+kv6hYqwyvXv2kZA+AlVxA3OzqV28TOz4mvoiXKOGHUB/yz7tyAsbSxsJL
sP1W1Af33T/U00FSoVXAuJbRZ42mcuCl+OMduvMIFxhjZqdMFhQLf0yr394m5hya
pDuqlxSIoq/awidGYrzZJB/sB6Ugn2jW7Ch8QXiqbSeyX+aYGdQDCLciUYHqzGAy
pDa+7DXa2yxNiBVqZAuNHDuG53E9PZdSKw/n/mfVENU2eW1pWbQdXpy0uwHEyxST
pOSZYzLc3KwnevhbvNu4u2pPo2VYvMom+ORrw626gXUIZkEI4SWDjxaym8LKrUMa
IMF4+iHBj/+l3nhyxSsksfLOBpEMSCYCpcGXX/hRt/GXT8Z+eb7N5vCyph7gyFQ7
6qUM76i5LD/5IMfsfhQgUxzO1Zddz2cJOtfy8iRn2/9tmghIVUk2h1Ii2v4qAN4W
F+d5sNH/mGut2U9mM0AotWY1sQqo5UNSh2tNg574R0KKuz/ILRfMpkQEgBOwtmiy
mtsetvrnK1HuMPVPBQ2G0kNfQxRrM5EXA3aw9vo3j9BmfWbvJvEbAzn6CLLYodFy
9LAgesGagYpgR1B/eooHRdbUscrLyj3RZZf0d37bV9BMjuW8obfvGVltx/C7Yefp
BSlN8mMqU3Pd5s5bRPqbdv1ctalOa6gG7iqEnuMas12tjUqGQPNLxljbe9kGlzDV
uAF0XQgRFUXhXGUDQ6mf9DqWdzmdnNyl4Y9WUat5YjUwY/d0EcPHTY6ihX3/Bie+
tJHzS1XIsCdrjX2HmHco78El/Kq+RLabq1t3SkeawoJUanMm6V0PqfD5IocxK9rH
OBTIK7Da2GIKCfiFQZ2T6N3B9FSqSsWLVIwK4RWaVle8CrpZr9D6Zv4BMQ8IR2OU
PGM0YP3q9CccMvZ0r/HhA1nL2ek614InvSv9fUbkzFsRDEQobbojIZqH/blx29tr
kQ2gtZeqIldweTBd5rjNkBypMEuuOdIQhDTkN1bHfKhrahI4Kq/UFV56652+vO3u
AIWLBqqbJL4ppzc+37Z2VQw+ZmiHd2w9tvAdn/laG/nXwhWtAh+b3X2888JUt7bh
JAX2m+0iq8nlbeEmEzYiiBdXUwZhfMZR4bwhdAc4VZuiZmPcM3/8PdQWajBqh97x
/NYg6IdjyeksC65ZwPBpYoZ9IxeVkukhIRA9yzplfGoRDWDOWjpslskdDifS7A/Q
/LBNow8d0lRc6vvfYRGCS3GNnfNc7ibgmRwzCEiG9TPoJ3u4zz8Z3ayBYaLgfTrR
re7iS4Lb4EKGn94uL2g6vfWqUgg4N2/Qh1TTkWalSfMTQUppyAFIJ9bkqza+KVZt
j1B/k/tMsWiHcdYHnglYeMDc43gsLzXf0HERS2nsFOxlgiZmUA3n9XGA8fN2vfGS
RUJfRAnVuIdG3cK4YqRalZiFU4u2noGGdgwlZiAgFMApgl3VwV1VGfHdXFCB5ncn
ERX/gI5TWHKq4gtR7g/sUnUKG+SGqHZm0pkpZEXTx/LCWIeCjupFHEOhc0g9r6KB
Po0+IcOuFDsH/UCyR9ZhPchuc36twKE/ImAhf2T6WvKaYekEOA63q1f8aBxaiI9U
GIKJKCXcWNmpNm4QOIHA7YBta4EcVsbMiCdetg6+vgV0NW5p4mawvjhgOx9lldIi
uG6ni6Bxl66TDGE50aQGYcgEm4w4xGYsDLGlGBXwrphW2JZg7DRcYr802WlWltgD
xkVgLREhFFRDY+NBO71NJvByAONETlzcU702oUlA2Mll9OwCLpmHyztJg/zvlZr5
jvAL6Z3dMwP/VueGL83kXBhl2YviZp/f1u7BpQlI//qPpsK5ZiAeI5Cq+7Wn4ctt
br4WfyBKXv/++ylGybxb/6NbEOxcdZB5f6zEVSj2506w9f6BBp833kNzPSByA23e
LkRtrmTpe1sIkArcXMUSTx1r9iZwdeE1cY07EoOY779/PD8+ezthP3nzFAerGWJ8
4bPwC2AJKsfwtacjwqbVIuvMPteUuXZw9QUvYJAeEsf8la53s0NKsogwp6Kl1wqH
/IcHXp36o+BOaNEh62zaNbcU4km0NZ3YS4YvfTgNj3R/YBZ/jEg3lWDh9RK07E6G
VMtnwngcIyTvraKPC+96wHV8trZ5lTuCRNwMtIHA3lOkam0E3MO+N09VgUtQMOC6
y016ol7VaT9JYNhvBfpViHik28bywmxhYzbBaz7un9P0kcRC+LsaP1sANa/EpKgG
s3zlmUJV1MKUDOrbQYV4YmaH9N8TGJwyQutDx4wNMFQIkbWXhFF4qA+Jgwq1dZmn
vM5u/yfJ9GZ4MgjfGI34apQgDYp4WURctwSS2tZPXbQO5OpciH9rkvaBvhhpwWTZ
xN3hq/k8n3JAMBdtGpVbTn6xvIbNrisqRiz930G0QqntQtTsS9jwXeV6THOO6UBV
UWRj8nszil76P2auYAY7A2r3UqvEn4SXsjTiWDq6N9Pau2S/cKMwJq1ooFClpZ0h
aGD7fN/qrKbiC1j1mIVEOfG4WO87asLgBbzNskzKWtf83qynLqHhACTPRsKwf+dn
Q55BAkbj/XeUrEvYAMNFOt+Ob869FRBx1AGS5TlMe9elnKs90B0RVFPbb6/wDDC0
vy9i5ogT3GlN9xtTJNyw2ClcUUxBx65q4LCsjxvk/oOHsbg0m1/AR2kHJmKW12gG
e0IeoIm3K5GUqJvKy8KShiCC42Jq/YorZ/pGUePep5mc3shpXcLKnV8Es9aW2GIM
6ZMAr0MP2nffCF6hQc2x1xgjqmvj3bouamuKCHmsP+5QdfrBK9/DTOyi251nDom8
YWKL5/zeQGCL5As+ffv6HWq01e1lxHKK7847IWsrxoqPmNP2ZrvAT68hU5YorQyD
yfyRkSyFsLRTBG0/faKKFBatrma8623iqSL1KtLvrAP8My9ouy5eyyV0cU/ETyVj
2eSdLtEcW5CMCKDeigAj3gciML0eyLctsbkjGLXeW58cBpZbbqs87pUcj3vgsVg2
YT9GNqGKNR7LgMU7wldVUmnb3GBfE3mhRVaSp+de1WzVzAl5l+JYMqoZJRzrxWZz
7YHsSmjjMEvvLwzcm2Du5DEhko3BV7uUz1i2hLWGPIGFUwBixo08QiXP9/ncIYCR
TquK9rVO8CSnRvDxuxo/RFZhnWZkcVa7D6uJfrurm9T/lbSEa9msqMgd4dC7RY6A
ELn9i3oyptrV6K1vJcXNgWbGQMOYnQVxLi5CvVJAjJEog68OgyJGcr6WgBBafKQV
x1incbJVcX1MOeLn2Mwb6vlZY26LLRL73ZOU1qfp3mnPvoqNIr32UPt81B7aGwH9
/8ZuaLPRiCOwRgDCDSrvFrLqq1OkQ1lnsG2gvFFjBQfXa3umcs0yUpzjbDymEuZS
Q1A+m30NwemAV3F84N7grTT/8mcfhc+NysSOkMsaTdYpqmAdV2ShRpH0KQqqo2NS
f48C2uqA/Ucn66X/JZC3F/fsGA17FSH0+KSeJKpW7cRfLMbkF0AKGytAmbHRSMkW
ew2T/tcYTqhDX4MxxryU60HKdcYJ/jcTms+y/Ul6iMRrDpcGFwqz9aKQJ8AYdCz/
uRqmlDu1gZR9Wf27N1OtLKkgpjJXXo0l4ikZ/5fRd4bwVD/jCCmqQ2h4ywueGuXw
6AAWaGznSjJZ/CAf/nknuvdLfhA6jsr3l938CBQei0onFYa1Z37RSWDW832wfyEI
aLPiUa7utkT1ALI/Vdy0ltkvWRRtFagMdlvL0mQHfRVElw+RzrxmXJfojgn2pe9m
YFEAdV7dEHPdK8bS3Xz8KOSZUw0qFLxeUxKbxGkFOKvymE8jZXd3lWyY0Zsdq6au
xJ29jfoaf2bAk7CIHRFeG032NELl5dbgV2E3NrM1ausShpdJtbgmjgJvSbC25oIR
iziGmFaza0NDKsTU8iZ9rHmKmqb4r5SU8syayB4G//6569VF8Z67Ps7xCIw3zRNU
PYoRv/vk+IUnlUQjXQLb0x0Bqxt/Gwo9JOGRGK95wkRhgOqQxMhNHImY9K9lKRoB
1wQMtAGF6K4Cb7p6HangBMVrw2zeWHOKvyvzua4Z551osiIvBvJZHosj6P858asF
Q6I8exog0pY2DwfaDp5DIMDYzoJVezeJ/HOMDoQK4cImU0qj9UooUq+feYb3ovl5
//o3zYSJykqYtnh80FYpANJXRTAMHVGffC+McWCLq352pA6rj+CBVA2uyOM+zSYm
m2LqiKwzNYSsGBr4uY4lOTSg/UNbzMk0lSv7uJVvWz8dcm1h6VWX8sPZX6aCM3vb
fLZnPecZev5uy4CpKlgye82oNfh/w5d09tBvF/M/34zWKChLn5VrIreKPDxMxsnL
HlbIRCoCxinPMR6KDEFRpib4bhoVr/vc7HZ57Ohfu25TXtZQLBtAKuSYJbAaRZwT
gbefLWFZRPZXTUYtC3ZvLBVO22UmmYD75/pZbBYsH8MvfYYenTTB/+OV/LKdfTzi
cOzto2KOS4V9ozxq+22Ww9LCwjkqBGS0mlpIg+OKT9Y7Xr95ojrzROs0dtOv4QuJ
3HuM776KPXRT8Z8KKyLgO97mdRCg3QwIjq6y23HLf1mLOjOUcSiR2EMrSZ5QH3hh
VtTcC/TOqydCNaZLbp2XfryY/D6WsgIb1zKofGWAfdaRMZLfno9Vivj4Si4lZyZ1
CKwLRhDXg3BRpOYxh26zD63FRhrP6YaqF0wLm0p2V1qZvRe04V5MCkyO9/BJ0Ahh
59+pvzuanL9kGpdNwlrIPcTLFAbCjpW1Toq0tZeP3AlwfuKSCAEseYCsKS+cCvfL
NuMl6xEjT8ILwt8fbj2DR3z0TNXnh3g2CotJQ0OpKZiJDK1i5+stCLs+rOqlaBUe
Znv1eymUjmxTrebHbgsgzUO/AU/Bt9yV1tf979O4UmqNW5n0kiRSpVC0IMi48Rh7
27aySwoor5Ia1+42CI5eRR4BjzJj6LJPsB82JrXvEWXPhKKAZ8MmUyM+YXvKCMle
zkgmCz5wbE6nDmeZPNmBNqCyedqb+63D+4RTsQa0jCTjwCobQ68hBbgCMOK56m03
F8OkRj0V1hAgcVBx/h1qZQhHOsKtf0/fyf5eJtGsytmGsacstXtRmEZtO/OjYEbn
s+kumpr+AzAyQ4yjS0RYr/M5Mr5kw9fHC2Y2s8VIU+4zBvXMTm6uI9hR9g0ZobnM
s5EIbdWq0zwcOsTOrk4+/IA8C1KAtfN8z/mH1R3s+Hy8XjLxVgugImWWv5PSQ8s7
uCNUwBsrvXNAXvisd4gWWjcqbhgn9M4SGisJPJsU9S3AqUeP6PEKCv/FxcV46OOa
PMUTpePpwcETj1cNSbZuzxMKu4PtwZ1GriNC4wkSbAHgBB37JzDNOkzmV4Cfyoi3
V/X3foJ1CtMwfsUka67ipYa/E1XlarA9WrIFKxqViHbTC2kLRMR93VZ9/EmV4a/U
vM/fFNc41+3vEhBTUFh9YS5cx8XLCFWTqNqZjCZcAP9+8vjNJau8S/AilZFbPcqO
UUmeafPvAc9iDJERghbcb4oXgZjEBzbZmEhs+VIs0Edos9pxHAt7y0qqsoj/rcT9
w21yz14bumCVCKM++t9+uOwrOYohjzzE2NEZrByAHn87YvDtQp25Rm/6nVr8Tv1G
TQ7DxALPC+426TNhAj14W3bO2Br9rAc4kB1Q7fo8ns3JZBrF8DlRKiB2/LoHKLw+
VGxkhMR0kQZJLA22CeijZ6Q1z6rwi9Vt8T5O+5NYyAVWcmsSXDD7xOk/3jtKhPMs
SH7FYH202BqB9s9AD6eVq5nENOFu9WP9XYhQmwidie+1ku/DjltQCyGpPl8ip/7E
P963J51ZZ+p2ygBRgEKpFhYufuja/yH3xwaNnGMdkP6Bd61M4lEyr3+pM80quIUP
t7yAzNDZk/kzbLj/XtpdjByjWkEXU8movpcrWUqzevOpnnl4M8pjjBXAw16tPDEC
0FS8xP8OUbgJ2pEe9rqVmfnyKaK5Q4y0pJSUrylPPM6bUDjOlc3QIuYbo/J//mF+
iz7bcLi5zeDpAetymXVkvzAwIKVlOptQbX3aHVAK5ojnVccEcERwLg7mBxGbnhc4
2BL3JcOa88eLGbH/QfMmRivluLm6xHUhBtHBHSLaVwBVaas8QtYdTIgZ+twvYdC2
2mMeXJlNdlCk1sx7l1KFVaoKQqhtRtO1IGtCFpDPlr2Ci2FmV8iEf8UlheZVpAoH
uq8bxzD8vAnL2yA1tFaddbCHSo8+P1mphjKbhZLRgnSor+dULQCYEg0+WeJ3Jf3c
i7UVaAePTen5Ogg7SIihqpN6Sb6mkatiiGK1R1vNxjnIxzYjAzNMtYQnJMi8EJ65
PkCsmXzMILWVHXIfE3TVYr9ccnYd3uBMpKpMpbx+hvLfDJvMIqFphDMhZ0XmRfW1
WIbxU5A2RxlKqu64BeGLBne/OKJR8S5hQeyAqkBpeuzYTa1MvkZ4yemPF9DP2jgz
d7zRlcNywBo5zpjvz171sq0ZALOp9Dg6nTga+PMLG8k7v0cKO46wqThIYnae7iWn
kLaS3WrWG55J+kcXLOlaULLvakCkKNKEXOPYp+oJwzuVcQI0vMJ3ftMJpcunCPfc
pDkzs9153Sykg7WuPk+QQBQr16TyaqQJ9dlQLNGQIDyqMEAAS7AukK4uwh57JM1D
pMcP0Po+x517DFCNWQ/MAT9KvD4XOB69+Ds4wNIFpQ75EzNYD1JpVbiBRieRo9CH
aEe4XLkjj0Xd7qSLzmGZ8BKroULX2CLeryom6WzaFY4r8Bl6jt07W8Z0RvDm9azw
/8zYJZ81n7T1HEO0GqNO0bG0kbFwT3EixQtzdmagOKus5OG/ihToBojCvWhil0LP
rJb1fmBfQHlZ6RTWOzlU5nTLbIFV+ZguM15BNLNAY9nV0XmuMauOiW+L/Yf/TSYg
6BnxHqa+pRYaghz0iSXBIgGAsczkmrGRAMLxE4C413+Re1tPK+9nDtR3neXLCShc
kNT1/2Rltiog+7aiB0Ci5CajBUCeEhqZFnQvvQk2GTEJb9hankoEAPLhjcaVxNui
Q/qHnQ+sQvNvqUWx4jLy1LqubqoJcRV+Uhqq0/a4T8nA4S6v0AbqAjeYzP+YMK7H
ZeR+XGSPkWxyaSrCvwxfY6NWb08VAXbg0UvpzS7sBknjvKXYDVYwjuWa2WgPJCSQ
agAvj7h1lS+2k4Qd3GjfBrsgydxLYBoI/vN1NVrA6jDEzsyl2l4LTVm9GfccYi0P
sUiIHE2Tupp1vHtzH33BatdYCkaxZYH4ukh/fPF2R1DRcl+MIyWa3r8H8cg8szel
RsRtK0Jb5vyZzls48Bp7gBqZqE0u/cUZO3R0cRC1vXYh5XYwD3VT+0ujaZ2T3TbM
sRq2WNwrIvKlt+MofcpKivpOuD+76iU15B4z2xVpWIPQgLFD3AWVvXUZBXcj7ItY
crDrHnStq7hOXgY49M3MZ5xw9I5A+l6D1sQeGV0F1iy1G6oShryBcU5KRmL79JFv
TTaq44YXegfIjWw0/2q0wR72VU+4AbOk296YIuNjArbqbMYld+PfhdcVD0bJ+2+h
rP7MBkapQZ/Jyz3OTWusvkhNAOe84I2IBrUYTTetXzwg71oyrHqC+3/rtToFDdmp
v5KDDmx7sfKSGN+Y95WgaP0sytAXA4mQ+FdEqthlYp5y1xAd8/TFtui7takem2Gh
wIomUP80NCKNBYiFgyoarE+m+URqCqdEjn0EKR1vT8EMBnDe2JFnQB6uDCc0AYme
hn7jtDad4ym7BfK6wi6Vof27i0/t+EE4BmQ3ZTEnHfruBzZU2hMEmnzF1Iex1P8P
wY6f99LpY0DXPamQx9Npuqp6qId1wZR8WjHhUYmgs6AZVVDI9IhxqrfykZ6N609l
ZsZRJihLY/Ma6+286BL8UvXrGXakGOGqqHca/yvqSKiZlo5cROywTBPju+yaXqeF
eVKlx8YFnQ75NiOEqEYrKjOvXG2KBzIcewJTAtYemaYN+mTi6XZeF+CXRGshBGF/
Qvm4xSqjLFnmvK2eMleCLiWaUWhX9EZxNAwNwQlsHLcSHEdqbRiENUYxfvdQOXf8
mtZZeqHb29cWmttgSOlsfHvGaBB1u628xQKV4HaRhzDe8VyVynZULXPJhdFvqwOw
aAoeKu85SYya28pkAhibfNic/uiGiRzNmozjeeMHvLq5eGcZ2/WT+YY5MYyvMB8B
J8V1FeNMqxhwQq7GhZmFMKN5phfmqMKKNKhUhY0Y/Y1T5zn+nfEhfhAB9MW/Bt62
qNgDxWlYk6pTHVlLY3sevSmrtj8Jw3qiPlnBVNYVvEs4PyWZFOcHqaf9j8iRhTbG
a4P9H6g645RMNx2dix+9+SKiNU2pfEHgYtjxr14w+OiOcVcxZ6ZkYCaomnNMJNPl
y4fY+1Nw/+0323tb2FuA46WX7TyCHt8RzcOEpz3ALMeO96gCumLCeDGNVtzuTD/N
7t51FXBbPx2YuYuOY0tCXiAS7xSjqk1tnJe7/LfJ7/QVhGaUhYxwhTKqzOkftAor
JSojN3rBtoG8FP76wLU297ZPhvDAZh/OlGnI1CBN+GVsEeQsx/PpDYyeniPqGBUZ
gEpjm8794TE8cbupHc9urxzpZOY2raWVFSIvdFQURdhNbRQTCWRbMGzCekqnCndb
n6p7Oirj/1hXINCqLxTLD9v/EaPMgmsiiWvqzDEHiqYe6ugzXASoru/XcebgJZAu
yzsNpWxDKFh+gv283iYniTmnoJY+KTxtWO2YuRxNrYMw2V/UwvAQPo1IkYzAH9k8
0DVBABYsBZMrJVjhsTfeyaD70HJBW6Ub42e59rBKdTwk8hdTPd95cdIh5V73cYTa
c9aN2/ppmmNXKP/UlWOcS4dgUTR4E5aA1toTJ4ibtkN+uTc4BuHE11cp8ZCzo+Tr
1YoMmlMbuHC3vSvSUUndW74Y/FDQmDSEJH85zQJK8MqCA4o/wR0oP5pxeMYwG76r
Rg4mkfa5V39Z8r2ZJjnegGv9Qkv2CVUFknBNTSSHcXQZ5DC9NRbXU5J6RllZ3j2B
zn6bP7C5dfcRXWBzhJUgpTScLn1oslXAhMcs7B3GGhxfFjAc+XYb25Zr+4VIZg05
GuCUfnJWqf3x7asOqR/Q7r7SP2e6tZjq5uvf/PzEGjkug0cMGoMCYXg0jXKml05X
Oy0chjE2NZIInCObJX4dr56s8W4HZKjrc/rQ42otK7dJdy8K1g5xqiEbMXfClR1T
B3LMDeLOhY54tojDUbauIk4QrZj9AtJjfPEUn/A2+/AwGnv3Rc1gPrBy/VUUicHs
bMfeTsVO5SAzCs9sGD1+Mkan6bEvVRrkd2sCxbva2e5r/o17dG7pBWFxCE1L2D4p
JaqtzxaG7Ym5FJRSdiOPjMc/FvEDFwL7+SSl0qutTSSRuKqJ7L6GTfHrgklKhD8P
nYCgbJo5Io4AUeNuaE//w0Wu1PblEBUhMIUz1B9oJHwk87njTq25LtMppfhSutxi
fMCZN+h79d+UYtgKP8b+wpLXmoIW4Ddx27/D0OK9cJoFOUmN+Yxb4/H2IxaYHlHi
sh86GdUG2scRiCh1mVMqQ1ba68Bshs6v4xjpm6429fQdup50i3GrkoBZivhX1S2i
3khbRJNdob26/F4MgaKmVW32UF9tP7ZlccXlkdGuQnWT2XCMEw11V3dP5bT9nFEZ
l8nEZ7ZfZE3YP56Rzfgi2x/gxbB93gNiUWtL09XQWr6BggImFNfubWKi34UHaR3x
HcwhBildUjX5Vvx7pbonPkGfCQ4DRGpAcjlagduPauxu7xAKDhpmsqcGRp9HtIQJ
MycA1vEIpbGjA/ba2T6hqVlkkbP5Hx85E/kjIx8MbqGNS6EJ0tl4zU4xeKYhEVlw
phNyN1Amv8cRaQcC4tGmhy7VGNz0Cnoa69lRQEYkprTQvLmUZCKHDXNsl1aDKYO4
zYbQ2HAdUGSytBsycQpA+tA4J1hjXDbWeGb4wGFITes5r/M8qC9fc2nP3UPmjR3h
OBs9FkPKktsxUD308Wrq8SZE4QuT+rtPCbtqMdqFJxkuZKaAisPMLBMOyoZ5C/4P
95UNeVysAh4/t0BAOakRluelZBI7NchSxlSl41w6XUdeRpa2D7P8Dxay5aBVZVhe
akfsyzNrzAR8iP/nAvltlysmrkONuS7TujA+rHwpiUEhLZSgkZFBS8+qT66g38T0
GFQQUN9pOnQTFYPynQguN5AczDHrL0AwBKjcvrTyjnGjGxqdF1vpJGNyOatOCj34
EQa1xBQoqQZ5XMti76irvfftAA0aYgPxW0g5GgUYPDET9M8ApD+QVzZlGkYapVFL
ameHDQ6kSXhxZBn90O/wlhAW/9ZPFEEJTI2LX5WHr86ZV1zsJtj+zWn0N/qEOyzt
FLXCY6lctVzC6x3Jsbf/aOyXvcSBig5bzbyTuNedJHaaNptBPYdj2goMtHRM2dYk
7vg9eGkquWGJE9PkRO/G3WTypSi+VKM/xccJn2Cx4130m/C/V0dnA9uFWS3Dg9RK
HoCoJ4z4AhMwV9fVccCysELeLhy7OP0N4eYT7hYNmRaX77Ibv5L44/zk/YDj2UCZ
uNoYpw/kUFuIU+DW/i2toK8I0aF04d4jR308L1FqB1d+8rMVebwARwxMP3WvDzjb
anlaQPa2ZbEZFjkLWNC0OsNqmN6Lmv8StUYAx29jsdlRXfb4yreZ0muyb0Qi2I7B
ergJssT1QmS88gIE5yILbbM5BB6sOeIxuP9FZ30s3Q7XAICsjk8SuOgekS3RD6GV
CiCTjHWeH5MZUJJC3jmxDYAgfBAMC6Bqmx6oXXTQXZ4H6e1FtSxA+6uZ/ABMJa1K
SSZWEqGtkSqYC/PTLjd0NrHsMVA/I75VYlZtvzDfDJdihVSAn7aD6Dd0h/ftDDHt
WstmJmUuYPYRv5cFhxJerPJ+3VJAtITMrldj6QVff4V/ZzLPQVX4fHvqFtH8I2tB
laq1Qb4Obp44KegwKY9Ofo4R1joe9hyLY5YDsJkEqV6Rt6hZy3vc3xF/qJlKf5gM
rBS+pYxaHfT4BdZOI9wKrOFbCz0ilCgBU+uIg8mKrbqbWWYtI50o7DHt/J4IRVns
FrmXoh85EoQcU8RKQjnWWqm6rd0Z/AC+qTnTUyGOfWdJG7n5cbRDqnvomyyf6Yeq
09+Glm6RI7BBDkbIOFRGncCCUnCam0hhKy22g+mnsyrWTvd3LqPW4gfUdQ1MvLR3
AGKczQT7qUHepZxWftUrwbkj/+Z3T8o5SroOlOqAklQPalsrdbaRejSLMlCGVVVa
6xrCzWt4HKDa0chILdeSH5WXCVd5wCRwc448fyzQBPgjJkqcDcpHzvlzR2jngEq7
vb6Xe1l7phrwtbgeikhLDYpVvJgTbcVrgZMXxFTj4/V9I7Hw4aOy+pHk1xNugoOW
tdvIo83KU044/Fu6iutbIhILNYsNubMFTaCiilX3zgP7sz7dplWlQKJ96TEJL4Jc
RVhN87DsrgZ24Y+BPtzDatXqV9Eh5m1kPSm+1/c8UGMKjFl43BOcfN/DPCY4Q9Ye
tDSLnvV1ptlLZT/YEzJPwZ0iSiiAWv0HVwYgQLyKw8axKXVXRVNpDvk2VE1DGqF2
a3/aLRvLnULy2wizmkXDNDv4PjkwdyFlZx02ibG/KuG0IaORaroAHlReuzUoATD/
XtMOIelD4ZOz+XN6ZcH0wD6ykSgB8kQSM3mLGCZAMl+Mx9qi4oJub5R2/5nINbDT
1eistRNLnMqpfthXyS1f7hQFwFmk33MvyZOfdp4WhYfHIO7fzAvkeZjpLGQOMIVx
/YIN9PEa7QkaYRNNvCOVPyyoTVwETe942HNXtyfauJCD/Cd4YenkqKMcaJXprFL4
bVx2cYq/Oz687hSikNqQJzV6S/n9kqgstq0l06FmMCVAus10uSaG+fKgR2DzYDHP
fjfdgbxt9KvI6gDqAOKcROteoePux6KKpDddy0MHOrbNo/rpaaEopskBh6ADSJJx
sV+iawXa0WsjXWRX96PxHML8CsbDZxCPnmj7B3KWJt+effvM7QtDo0UJxyp7F0iV
zFXjcxUh4jqHM1FfSF7uJKTwlQJlIMncHHslv9CNP37X8jIVxfh0rTF4n24HRULN
XSi02LGMTFfTonIHSo2x2+V39UF16jKJeXQcRMwfi1Z6JgWUJxUhKE7PhU5fSwKf
sAgjEemPDarus7XOBle4WI+4V03YwW8N3jOdyZvP4TORJUm9PU2fmCrTResKxRra
EDD0bSWnbIUKJ9fm+HE1KLZGWRnN+lk9775LAUJ/ccYq7s/QsFRREKthQHVCM437
jJzE5V+yg0CyGkoBkYYkPeUe8B7Y1EbBe2nIw7qCY9CIDXqOp3JAjplsYUcYEsqW
7nvVXTiCIJqDiDXFoWx0Ysu5lZKmOanCd53SezQ/kq2untqbxUO0uhEGuPHRvfsS
DbK8ZkFrFuQ8HqIJuw6yxeLMBKPIEkbTDAECBKStlseW7nE3SFOfGWfmisahPybn
IcN2+zIjZbEqEgTN8RgCv18n5nECRRoEQ2rdsyjpHsxXK1in0aeZQEuQ83gioHas
ySK7igu8hvdptI6kl823t5nxHpXp/m7KNFNUS5pcbJgJ1lYrjAEEp336xz6LW7UU
dlUuP+81tjRsr+fChlJRDF1jxNZOKN8wsiecfeUICkpJ48WzcxcGI11UElxhYTjD
O7/uiH9pxJwgTJQV+xa9OTXqSH1qlzJExQTRCoXtEr5//7/gEJTUE/eVd66rAt5T
v4ANlg6GZFVt8zBVkuwzRz/OHJ5bvZ0tiaLgDoVenr2TgQzAi94B/d/zLu+Zl+rp
tNWH4V3zfJ85zHIHT+2jI71j3lfRUbzkdMaFlct6Hmp5vA0F3U3ojes1H7HKiIug
pBuPG2uTqOtZsaxyrMKO3KAVOrMWOobeV8qEI7sHk9aaM+rgCqwXsPi8aEGNZvqm
oyZgPnqiDIJdwgYXcaL1BlEuJGUU/xqg9c6Phn3someZpqCChHKMTBnfEsMOIAYe
XYJu+t7rcMBi/eEkm4D4sjpUCY4nGpYlF6v4hk9DA9BiS2BZp5WKYtPPLykk6rT2
yw7F8Y2s7myQhZavODJB9T9zMnHToNyNf7RpU5la1tF1Vma3ZyO54sCkpWfbleme
MK23r57zhMQEhy1Fdbaai+mtV/AMpxU1Levy9b/IEJa14FVPd5IonNO0Ay8SbjZG
jvW73RBirMB6gpIBq8cRDpjutROzSHphp/lD4FojbkBBO44/AUVby8mGbwwD6e+H
a0ujcssqtwW9qJbdLkMYAyY1ECqAcEVy3mbIo0uaeAE3FDLLEPYeQjKEE+Ulha1I
qFUBkB/Ebdh9iT61u2vWg3E/pCmstZxBLo58Nd0B/Z9VasyVIoEbTuRoiAG6XdQi
6WtG48lGoAnPoR87240ZCBt9wHJI+DXAZRlpOdl+6XJr8Oj8HA4CY9gKh3AfDQYN
MYUHrotUc6c6+xwr+FjD3QPw/T7nq6RvgqYMte/HGU7IH3v9PCUoWNzQMIJtY62m
R56HPk6vCqFtjwPBLZth2A7lRno1Er/5Oqtivi+MgJ8SpI/b7vhUXh6iVoHqzF5+
FuulUkXNHbnWVo3/DJZNCn9ChEcyqrdTCAQUIqMOeCH0keaIvh6gtX5RLKjNxMGG
EDndcj+koiaTKTvHtn5l28qD7poSfZCiPncAejAjVx28U+BDE6deqPE8xSCZgTtk
n7KRab9/6RF8OBSQfnOYClsvgIRp94TFO3stpG/2fYjjMZgZJquIiH55eWvppUyZ
TNpfUxG/jwuAbhgd85125bdCdEaqm9QsNaBOU8yXoOshL+s3YjnBRRAjR6HUDARC
MkYXN37cQEAH8hjADHO5QjVVjEAVX3orc7VWemc6Z3VOo1UTmYWyhno5gyWKiwai
HLiKrPsnRjWW5iOXmN/Coigy4D6b1gjSJ0q+1Fj/SOCjWnA1ZitI2DWTvNUI6WMS
yBox60n4FQVe4nGjhSvePvEVFI4RxbKNNw4ZMV7IXjVWUVq6Q7v7E2BkszsXEW3n
k62U6XbVxQ9p3cSk/a4vdU/RvyHFmP1rVN0AkiJGFcJqejN1zRYMAwCxcd8vviIL
PqULxmw2ZxT/Mr6xt5kpzAutfBrpsTcW4H0aFOdzw+GNQdzrqOxih3QzeG2j7Vjg
+Zek3zUbM2XRr9FwZZtfP5KMAoq2MjclCKYX+Ca/77wt+oTU8Foq75UebVQqKve9
a8IvWpJ2XmaYMe5MFBMvZ8jkMwNLBmKHU6y5ICvX/cdwOsPt2157Abe9PP1qV4MJ
cUwCjXpYvQuBC4v0W4sb/j/GzwHc7wX/bSoooaODSn6mdtNNqeGKrDoORAKBzBNw
TVoauWSTtERu+I4T9FDm47NhUC7/Wgh3EvJN++9UVbLJ3eMLXsyOGHA5XZ5ou4Vh
IhJE688C9OK58AbCIEnYCb6MaRLHJyEY30n92PUpOId7yDzsC1VWWmrg4vz00gEe
Yls5KGnpyP1SP9qaKpZM/+d7ZpqnRojhh8okZ2vD9wDETNa0WCoB8Ow4sEImZ1E3
TKLUEukQ0YjYc6qdt9+tmdxXKTs8TpScSQ3G4Zz0tViKc4JuQnKyeTREsbyOQXps
sXfU/zmbWOoKzadVyDZP6S+L7ycQdEpZ8T62FR07EbshUD/heDAblUYLZVApltLI
SmyIPYET3bHvk9hkxAtDVA87iNz4RC+q01QdjVSlc6SfImMNvpFuAgYGqzHz6YhQ
F680sVjM7yXXoQr4d6q55nnbK3ryI6fwwMq45bpZQugAvNYMa3DwMNGB51Q8fR56
rMfEOcWEvxsrUJ7Dz5Qe8NTLfIpVWNFnTtOe8zDWVAGJTsyWcz1Q4jN9jwtOfCrr
i8VrxXo5IVtJP0br97j91QNY+C7fiHpmCktHCt4BP182vBGq/qu1FdZ7iwZ2H1UN
EocWhnQAk7OaSLqq0d9fe20OCjNsdBqp9+69oiqrlMxv+wRWwBASonZY7/uNQecu
MWbb6OrJr6Cz2m2Rbj54anXHuWd3mWlcK5mRhwNOwYZ1B/LoIubAZtuzx7sQXa3t
knZbRbiIr/f/+cBIDJptQ6Oy+0FHYts033ACUxB+uqdYDth50Ibv7n01eJEwvcqJ
kHJbK1I7C5I5/be9FaNcavLfZCKPHqsNY/623gcnZgkPoGcwlQre9XNIgwFG8ZN8
Gce7YK0puTLU78VHOggdmuR+awKz/ntZkegWGi15k/FGahmXu2nwCjmu7XgE1Lza
Ay018Y/S8lWFaAVWx4yEiaiW5Yf57TsigWrG+VKMMGzUmuke4uAQlHystSsLwTSU
S8wojAXyY5T60w1CdQpQ/UPstZc6qlQg+/DBPbE+gUGTRYlwiSBbi7ZJ+K5ZSK/W
rFU0Pl8+/36xB85ct+Ev3/NsisTZpV40H+N6sGCi6MfDxzos3T3jQm2srTZCx0nv
6Onr0CDgawJERPnh/f3KAt6t2Bd15N263/qLvJtMIA6XIC+HEfJAUctcwb/TvhZk
CuyY1fn5Z8zkiqmwuMFFntXrcYTQo94QlzoJxyix3cYJHzsgB05v5K5v1qElcIFL
+VWl31js6uWhRRZDwKOLhhjJHRt1u1gh8cNbEupcJV4JGoNdfEZcECm022PbuNxR
BynfQV2O3ryv2jPmpRm3YPo5klE8oCuN7hcePerY6Kx+s6Zd+yH05C358i0DFWy3
1z0lfrmE/R7Ohysbz/14ox9eAU+wCg8LWGoECudpxx06LF/4zu+gXCpVpC6bnvKf
ghhZfXJbU5Ojiu+OAxjymt8I/yduOGpLtx8jbfc3r4IX7qwLY9aQGWFfipsYLrXJ
Uy3s4dWVpX0qQ0pUmg2QdJs0VQhz50FR7mxWOMXXzRO8V109WwP/UCQCaamol8QX
zgbPE4az/Tm8det+zLqM0u/2Zdl3P3UZvGat5/6WkJX/5v4EgI+NoI3SdigbqqJI
aW0mAwmRO5s5wFYYT0/bACoKbVIaKy4oWpgf9Yl68b/0VYyGiABJZhDVCKt3ubXO
J8fa9m7IMnaSJXWy3jX9qi+Q6BXJJ+JFQpebSI7ledTfPYX23TSNIlk+NNK6HNuK
/YhoSqUYaeXGU5zylHtXykvc2KgUfjKoTEpO2zBquG/Z5jAFirM3dNQ755C4GAy+
ajPW1+XsDKqaIk+X8II1airrbaq70E9jqpucuTJ9UNqmeMs2iGwJDo1twOmeCrCk
wb44g7I1X9RKAE8nqqs1VdOGzUBBFRI+M0ZnjfTDsF2ADodeRSfONBj0v0+c4G6h
CeE0PzdawO75XXupcHTbrDSn3d8Fdbtvqhy9t7i4v66/61OeFUt9iFIdj57oYftr
k99Dhp1H/Fgv6sraIMdIfe3DLkqvifIIw0k/p4Quz/6xHu5GpAxH4k0hsU4EB95O
/dOMksyf3bFzf54YTwfTFVrJvTwh5CDiWMxo/QKt4ySbQDzTRpFyVM7Uv5zPkXnd
Kflzw2KYXhgdb34RAynGDazwMWr/eSL+Ug4DRXLE9pRn6AaYohRBiyrLLZlkzp4C
DoNocQY2nuqkJ48U/CR1jsxMzoQg/Gn1d+2v4nlY2/RmLERMhvGQbud5SDpwLUoF
8jE3BNay1H63uTli25BpJa2/Weq3xp2/lY+pWfjp0YG1RJi8ZUd+DWi/M+38bnLY
EaEr/BDDZU3AzZBEwKbEve7sbJT5SjuRDurm9QpPOenS1MEg69bOQHtd8H6vAmIZ
b7rwRoqREaLFTtAQYANuxZGCzRXlxuLY3pEK2gae9A+f/iE3V2gyRN3vcvJKoGEA
D8eBcVQU3QJJ/6HWtDP9jXwKO2wGgfCul81VhwmSuLRqPaWGnyuwYVTEZQbg3p2D
u4QW8e9G+hNHd7Skp7ODgs6AxeLUSsTrQlKJ2R3ezl6cYb+2J9xGq2q3oomh5uGV
6wusJekHaBmO24i8U+RAIq5vhDHgH1KdC0Ni4KARQOHjX20hdH59zSZjEOlX3nFZ
eXPv2UuIQ9eGS1NivNN5KHOJcEgE50TuKomYctazixPH1lfHGSYAMJGYDKP04pVm
UvDxBxOTPq4pueCfhyoZydNmvo1ma85zv0x46ieHEhV5TC7xk4b33c2RiC0k3iHA
AcrhexDND2eqg5Z9emCZErgxkRvtlbwpyTXbQK+8KjcmztAt49Cd52YjawYoD47P
BxyWnrL/MOoV+SH2z+VoVSDBHM7dQh9MSPrwsuDJTDMP07/178HDy3msrybO1ERd
mH3PK6S0qeuAwgDVIBebNX0998dMzWfAtGNeVQHl52dHUdHbc7gVSdaoNeFKKqOP
sOEOqGGzs27Yoo3ZxFeTYmLRATtBURUzy0wxtJS4bXhUbeBuJkC07BTAMKJJiPhQ
V/M9CVSkd8Tt2kxDaQ4Kg3L76lwSY+jGJavXI87UQm8Y+DvnQQu2mq8d5wrJLJLh
RX5qt26CiEllyHD0lr8iPsRgx++P78XMH9vqwe2mQB9F9PHIT9/c8kfu73JqNSFv
xcR4QM/G9eAjGiV2ENSk6QoaAVbyaX7kcHy4Oq9hF0bCZ395FE6SWQPT9vdsk2Xi
FTC0pHeiZ5f16RXHOEzKcAylEPFmgRJXKeNHJL6dpCUPhiRXAm2CKuA0BN9yd+PW
EQ8sRju5t1NVZD26qH7/ZA/0Gh94B4Ck66Gem9WlKPkXZoAnRgRBlBzG7gxYpx33
f9Usr3BYANTdyyVgYdvbHlIRpPf0Jneke2K5e/sq2iGqkqhshnHz0101Af1TVn+K
kFCYdukgA+1Sj447WVMVskTcz0BCYBklJY7PUrbijFV7r0wmJchDPSi3uqCzexQg
AoJFi1GvQNrs4kZJC7xyh14LmhyGwI8DwcIyQLzK9M0lzLNhhEeekSXHYvqMLQgJ
tWtuSxMdCRcghyhhEPERbX62bBfwosuBOl7hHHgJIW/ZM5weH72y0bB0MSSA/+c6
Vjg0HS7owF871A8lbajlpmFgra/f6f9Qz3ptGPXrHvj9HfLBilcrOfXQ4d5ehx7t
upVUNnxKJ3C65wNug9O7LSlqsH1Aes4BD1DWfOr9JvwESJfJBtfxB6qkzUE+xIZA
JnoPAUS/rVxIBtinyw2WE9uC1QmYkHl9jcT3m/lsNnM5pF44OjffRPC2nxyyXzr8
vyjblGAT0j5poQrKu7xWEobXyKb5Zl/n8/nzSFcZMsHYuyYxSteP/JvIavDLZ3b/
zFNwvr3ljx2k8EwrT0J32C6aAbjmOIKP+8rKUfzSVmKprv1Ue+H6npp0COcVa78E
y706PWpwPxyy8G0hh2J3l/PBzDplhwMv6mITsh8TCRkIvSAhLQf77oB6IySlHS2j
Nj5wrAnFeCpEXIy5YJdBq8Fsb4oZJVFUlj0otcU/lBvjztTktKPS+J1dSFliQPlM
koebPGFr67GE6wJi8dv3NPu5UuIe45dtgnwAbaG59q2l/CgrBEBLDTM40cAAeKAU
3hqw/YtnE6JxHUhwSmZ0ydqTYMth98Jr8omiqhC6QbHOv8RX2ONfJCBiKbDJexwb
DWKLd5lirodffEk/Zz2gU+nWvYZNkNoIyv+roEuF4L8Rq17aXtjka6zJ1DuuWov9
1myPs4brYopHZrgOfGH1UYbu1MIccFDNHZeDMUiLN0bPwqWg9Wbl++Tx5FxeXsRh
/gYO2zPmjFZcQQ2ESBylLY1f8XnSG8/BFk+7iBilIwOYhp4xL7Hh0MPvE/INdWac
Jy2o0UgZVyk73KtRZofWW20y2xMmLQJ3dAOpum2G9chYX11gvMI2xO9W2PgSRrZX
NetDwulDuJUZcCBX1NKlyzFeLvgRk/SXL65MKGEJivkecs+WvzM9JEq7Y7PkqV0w
+XyZ3pXQxuomn+o9uknaz+ArAV+8QiCnk4Whi5ajeHCPJdPXvHw8epX64QVLr2JF
hqvqpckxoXlyPqScNCOnwnuOPN1/fqm7g+M0xneya144mcFZjD8IgjOevZs45eLW
yA2xiDr3l+FD2x+7liaiGR4TOw6E2LNuDnZc+17PumczgKTmRHn0LMIW09AMJJsv
PPLD9PPEO6ZGDrPdgYd2Hi244/ZY7s8ZSx5tcYOKYGg+ZvibTs/GmcVY09v5dKbe
mzkwsYNKs3BYHVSuRHWtwE8qGUmgyDVI6IEnJjJz6pmzQPW+CUnzLjDwgKh2ZkK6
kiAheIUVZgKsUUqU6hQnJ6dmmwD0C1cASTtkhUozN9aXwnvqaewjFN4k/hkZsibX
V2k6rHZoe6zoIw3PiE4rOyqJ82Wd+u4k/jvqw99QISpzygA4CMVhcDw1BBuQ5HkU
9kijfAreQrUxPDyL/DHnY4+RPx+GSLQCgLNb+yMZFyjAoqDssrx+NW4f7eqNdpDY
70zpnqVCa+gQi7I4S+R0Jcu+1OU5iPhC8Qe3J/v5Jargf7UWH4fxf8mzk/i1F/1J
xJlFltDuDjF83H2/lLUyNQtk+7F56CuhREuyc+02pOke2uZVMoe50VWD1uN7fqpO
7oCfnfYrBEv3qcoLWKsHgncRS8CFppyRQ5Fr+yRQFpcwoFZopRKi4eF6tUnYmzPo
llhCcUcanm3nYrCqFKDvMEibJoW+ubISIZTPs/3G/9D+Q9Ag9rqPsyJJqWX5ohH3
1EF9jDmO2bKh6YDGFJKv9/V+wvMISBwx+SwlgU2GUMGl0J8q5pjWX6oKbl/3fq5z
Z/w8G3Uz5FQm5YjxVfjexGxcvHU6ekwkxePItvjR+qr/FQIW51vNYUHxq+lxIDZz
1C1TU/CMwegNQcOSxzRR1C2+0mq7VOv8rGsjZpEy1JqSRWpND4qSfFjcLjZgBM+r
k5mZNQM4XjDaGMa09ZLrDuiDmGc/e6OUAdx1dggQfXUV9TLWrgl2CZmh7g8wa32b
zGqqdRNnRsvFnlcSaajtq23J7gMT+/LIVgzT67svNAsWoHVuXWcTvjsqc0eoigPE
fwq4Ylf0iGgBfeczOK7/MvF9uJOMGhFY6uM1q8N7Nqs20sf6IkahVb1k45sJEKnV
5/nbYesg+FCxb0qOudwvnRXhOG8aWIyahrOvd+mJ7f59zEuc7/aAcFUYQNhMACcB
kdTvx4AnKzJHEFkAV52VvGG5shUGUCc2X8X4je3nVbQlLEDIZmA92yuGDxjSe3+E
2Wt53GHvTw9Bi5cEKLZAcejOktvQS8PWJSQh790amcSwUG3DULYQGkjDS2GXK4vF
Pygw30JpUYiy5KmwbUu8pKChVaZyOv2jKw5fKpmunqrdKNk7yBJh9fL9Vgg84tbA
cIuNI4a2HSFICnElr4pSA6XxDvyF13qzumKmpGWITq+iyOFfGoeAeiS0CSSiRJru
uMNHpymgpO+p2V4/V57YptCZrTWDDjj8FAEZis4wxszdbrxLtD/+5OuLq6OHpltm
RmiwlUjatsxHsHbyaFCE20V1z7rJCbw+wDEHaNDwRPXzXZxAuEBAtR7YYjGjBnfM
XXPTUKUiZVGvfOeZyN3SRjqy5Hxw4yPptTX7kFfJUKTf1MZYhonW3x6/9sT2ExT+
UQjwwGnb6fFuoTWchbQxg3L509XNrvxSccg8C2UUKCNl3mVDANEUlpxMfkC+8PfH
3SmDTIs1/0ghBVVCitsHW+llAvSu/xT6ERBxSnDirQwDvsbacYHmO855Fyb9ckHD
LIUgrwd+/tfnG2HCO98gxlr2K0KqZLRu6YtMwDv38vgTZOXySGNy/cp8DU97AS73
aC7dQlw41EdFOXRc/NnfnVdVDCVh8j18sYGDXtBvmc8mywen1WKkr4UuAHDHhR6g
xXKAuHu00atop790koEG84vXuhSjXNyiJWFDQq7R0uVFXaoUqMdpVk4sUTz3mZ6q
jop0VL84JxHhOoKZgWoHCmVs5gob1W1O3I+wRoApu0lZAFnsmvN4lWL65p1wjVxK
0cxK3ZXLJzGZg3QwvRnlOuGxqq5tfQV8VXpmYk+DaNhd5KGoP+V8T3DmL0mQWM8G
0LqYZXCRB8hAhNFm+qzphc/A8X5rquhD13LvXNpu8TFNUtelYHbvFthnAk5xOXXB
A1xZ1zQzlw5BGUnsMoOZrcXtfwAHOPn6nb35uw+bl//LIn8cqG9BS94b5af03lPz
meZ+P9m5uOgOCgj38GJ6RYj01WsG/jVYaLuvOGNpPUrgKK41p/f/2VZ/giAXMT4K
4ZnKDEeqLj3aO2OD/8lcUui4/pwqESXXp3o/ez9XJ2VEGnGpLZrSnZWU9ZkYNBTs
ZzEO/tzcqXhyiAEe6t8U67L8Gi0d3amnz1kqiMqRnGWlswVQ8QH4DRF5c8+If/jc
PLtdE+cgFR+fUVI87cFL0UQU9+GTybg4H3aaR5IGKIhemiGCB0HZ3rVyrNpI+gZG
CN6fHv5WjnxRp5Tp84YPXKv9FxG3VJDJLdDeew3/VV3xPJedUyujj3MCUK2Z2hL8
gWTrb5j0VLOySZX8oVT5yLrKmx+tUxOqgvpgu0HW4JTxpGBY7Cv6UKhsaN2eNgrI
VFzaXhf79yAStaR9T2Q5BT6qazn9LB+LHSl1VL/9zJlMo8/o+7QwIihVwXOYb38B
B3AH0HefnOd4CGyaG94LKvPN/cyfG/BSfDT5770D7bRy73bkZ3juaG7H9E25RR3+
twOrQ8rWzHkyzBqXMb84o+TSkr61Jn8hiyoWf/uDbLYSJ7YWAx56IX/z2sgttaY/
ERk4s1CVzqd8KkW/KpKFPDo+pYclS1xBT5BPWfKZj3qtL05NXyn//5IRCRW7qujj
jvmpj5NAH+bHslV+5zmaM1DEgqunVuZ6ZhJJrhUVTEg1QYfV70SB1cxqRuX/v+uw
4E9XU0R7yRCPVni30UdSbPpL8v3B37fYjHiHNReQSv7JOzp/XoW6UL3c4Owenjrk
b38uyGNMA01+OE/cNN21DQGsbiiXNDEk6Ff/D0wT38RBpQERGyUjNR/rH00JsqjZ
hXRl05pmgqvacV0Kve5wMEqfyXZMyNzrjVPMmdN/oy7TtRC/F83yIG+sNaNHqSP3
vRtYf0NI550Jkv/K9/ceRsAFfeRCfDbE0IEvcWjxL5V2Aml7d5Mx7B3z1q9umuQE
qpcPiVyEOrLWZaAS2DxWH3zUrxbOSf1BMNYSbPKGwe+RZ2wJcdCwfIRBwt1Qmhrt
K0qrqcTPAaJJDQcDnCEUg2WoSpIfzZROG5rTDGBBb6kUs3f3XOkx6ITpn61fdGTT
EA9BZQJFsEgXEmW8bEEsqe39DfsWBTqHUh6gL3if1D+ACTPTROdkRipzfFWMWzC9
gNZbtIzsL/t/FKH1DOjSTLY7c7SRX4pwc5YX4aJ8+Ay7Re2sptDKJV1OQGJ7EDww
oFzMb51qHsmSbjhDCm26el46Aqv+BsR7BiexxhedFHvSBFlhXoMpONn4GeXYK703
xzJShsegZ+ueao0GOxBnMPvh0UcftptN8ecdoWpNiBV8gQdq+N10BxZ1X9F6WQjN
WlNrkS5Erc6VL5cuVQ3jdPu7yTmxUlDAs2CpWnklZXl/xZPM+qqzVW37rYBH6dXr
BxdSYdL+2uSMncMhESiw9f6ubVHqsc8tELzmnINPRoF0jZzzQavU+JNqm01Alpx0
q95nYPFQXSxYIXiZ8H6fG0A9I7nVp+uIWe4UXbzRdtNpAyY4zPOloSnvQy4ha97F
3T/LiyTULQSgeHYhV0BDGUy87H6WHAtL4VYKbY0vnfSHxIPA41ZeJCM9AhjcW+G7
/vtGrM3of00Tv3iyDgaQz5bu3lzGVYzSKQfhDHu5ijj93D2t/Kw2n1KBFrJ/HAJN
dQFaoAhxNhlX/jsUg8lRTvCONbuQDQae4kolrY/P6zqD+AnmuJCmc9QLCjdAAYuY
wckKPjGhg6+eFDvUOIVEwBkNl1ZrvgJ5Edlht4f4dGNUAangA7ssTXmT3WGiC2J+
QgfgSjrgnIp0LODXreyUW7hSMAYy/TYi/hVNSbKRkcLvA/jbkf++wW+gpViFEJKk
4x5QQ50c1Du2WdeQKmV0xgn+2Th2NEfF9cXyyZ3D1agbtGolYCZeiwwfDPMorrr8
uCl4ENJH/3e30t2nCj+jd2IMhMxD0HhywOtAwaASYPO48atzf0D4z1/qhwJkT5/1
esfC7e1Cek5R1dN525tfSJKpBaHuRVcE6ButhGesRnWWdEcPb6F0JQQrTXriHXiK
VWEIx//L5jUH7e2rJyKBVqwO/JJA952zSL3pyhOEwGnjxjLjY/P1cXk2gB3/stD5
wUhdI7JyeIWf+887cDXkzswUKpNL4gYBUB0MM8RltRKmB+5RFYdl16gtA8UMg5so
R9qdsvwYgAw8SfjVG4pnRpZagUOJsl2rwRXsFYwr0dN7Qm8bMT2AQBq9Yy1woesN
OyPigCVx86qqgHKBTvnmBLjCzq4dh43YITFMQsAr9RhPboQrGdAQQhNQQrv+4Rqm
eBe44V1HnzLEM+bi5aiIoYzpL/8MqGD3pWZjsW9azrK/pMDUP5JrCn0Ma3uyzvzj
A9a8ACL5ciE+r5YOY+Qj7HQq9wnS8U9n3v6zov+QbAKnNh/eDptFo/TU/I/aQP6h
b0PElmjhIGWngcnIrOYLP/xfqoKAbxqzLiVxa/kKjwt4QI59rdCYZbcYB1NYm0uM
vmpGzgWEwTPh96In9o8NYciqWVybzf+156K2uvVsi1NB3bpZcwdYEV+6mia2U9Ik
JbPME7hCf5vhzwCKIcBuJVo594P+k+ab2xNiJySVF5Cx9cll7+TqhzCkeIPJTc9R
Gqf7sMSsfjr/CJ4TJGxOE8Iln4Ia3xaHdr4h7oFNGXAYZQkGhbVB3YBBQ29pS4cq
BGMkcMSipiv92NNFjPgmeItKx8VFejjsrJrsYs7e8avCiEdUdyEwrkntBb6kQHri
moWEW6wa5PtKimsSZW2fQMADmdc6AE79B5tMjNY6kDYpxuXBv6MrzwcNKaRYJAZo
XFTIbxBds+b4zOr2w6Xgq90ZXVT3SAfvst/pHJ3NHgLvRv3he2HkOchFw5ZR1oic
XrppQPYZYllwOjnShyGouZzhgnBhOSlQXLQFkad/nF5HF/M8atV2ADbJJie8lyia
7r6r3AawsXHRDS8cP/gCpXUWTKfq52EfUFe0AoXmJ9tdrl0qHlUR13IxA2Qetviq
6NTTZGcaMXHWdEfTeMoxUfCxk4tAyYaB9Mvwhe7bhT+18SwKHIXL5VfXkgO+a9l0
FXMNAf6tTYe+Vb6TetKOSTNzqxwFi+fJy1F794sCtcEr1iqO79/0oBuMvVyyDYhf
m73o7dN9wj2R9x4swqEU2jl/ZuITRXLA9p0TTDLJLHjxr0JODLzdd0KjHe5DmL13
s369IWMuBlALWP9gyrMU2pRRuorMr1OF+yQsQyUsVyzS0RKtWJV4LdVAsO87dGeG
Ovj/SGbXDY41nD3iVuCNEjY+QtdZ2eySkoSXtxNJBI3V4kGHy1TuKNZkxp9964eA
EkdAKT+etE3Esi3461h3KvHMA/w9OX18jqbGCE4wuHVt+aXDDdoM2kKvaHJPE57e
s1oEcSwBa5UaM01PvZL6cq6P5d+rT7/ifrwJEqGflR8EpMalSQiwr+tYfykEzpcg
7XtiOrsAPWe7k1V3EIjrp6f5e/+U4/ZyFX1k4qoLBQyduHb6Ce9Fu8Aoo0pJaRw+
Olm6Td6UoR6XKdo6ABihB9ngdn3p6+J3y2PYUJVmtNeBVV6cwvJFQ9nrmF8MyI/I
dU8zqhTgnwRUq7X8vf5uMI/jFjRnD0wHZq2UvfIAvsaSSSDLPzZHP61CnEnq2Evv
KJBlHu77ZFLvGHl6mXbBUysQCyiJ1uh0eVu1T/j750TObCZRWF/vxupG43VihK7e
58+Xj0QKSt4m7wojqzEvbUJMaalw5O5xeUN2/REU5qIXSb7OBFmUzxsEKbQREIMr
SuBwp6tHV351e936WdlcTxUSWwRmLsX7jYE1OciPym0Qt3Bv3Bj8fg1RsdGejbl6
ftwhOSnCeeYb3RsyZn+10YlpbQe4K6eXZWNVMBQ8BMjwgSwkeCj2BX6h+aw6/BjF
sTxhdodRoHQciZjooq56ss9c9Vas5WY4Iq7C3n855vtqzASv2EC1aY2P3SdlMpnA
GQ6PeknV4KUHPW9h52xgGFPpgqIq+iG7h9uMf53VI90p71nCtWLNxypIrB0ToHS8
iUt3ntkJmwLpkH64QoJIwBllZYrH28ibXHB5J5ssCvSkRl8gye+cwemdpqzUqiOd
/yrp3FlVg+HHFi0zRVt+2SXGggV4x73gBs9Drkic2QyM0bwbMcCWidUN5pcMiYqA
XVz6qNmrxDwbiqhJxle9i24MVFoD41jxDwrvJmciZqE2YwWtOWYj3uTT5JKJmWUo
GzmPpmsyEfZP5WEdXs1qGQVSLmjUSmk3PDcrcwXondxBFgq/3taSudRKTAmNf90I
l622QFs5tHLdK+5e/12aCdqeqWZIK8Cvost5r3xx6PPhk3Lptw4+H15UtS63HhJg
CDvSp5W4YR4mx/hisISbOeIN6tldoo/Anx9D7tmHMbVfpaCGSBAGdJ+SFJHTN/MG
aan7kxa5qVMb3eBjqzMzF+Wfy89gKoZJv2X2PbMzeWKzGcM0IIKFC1dWuoWWk+GZ
d085AVsGm/J2mKXg4yj1kO4HRUFOq04QTcgLiNGGy1IE7IhnCXExdWB5ZpoVDu1d
MyfBPuDxRSaq8tW2iLhMKSkgjrvIvzD6ilwOrs7iAbMMcq72Blowlr2E2QkVj5C6
BOqh4EvmWpSK8gLvDIpWxksFMwac+pinutQo8UdIrzndw2D5ddHn2GmxoCVF0lhX
kRURV0ItIKqkUWMbhP9AqRPznri7KT8+aEOc253dfupadlX8MdqN2NR1xUg0TjBm
ALMj5MfRQpRgU9ET0odVDU3AFGqeq7MZ4cQ4htNDAft9LPG+ffh7olk3AeeLX69Q
M8TQpfN3yjSTSzM/3kNPpMoQq+moba5O8+KbGWu+zycAct+QFCZzgTUmFg8wB1hm
oMp+b8wtzVNybzIdqC9oQe5f4g2NXF5h+eXFBduiwjP0bgyy7I+6MXiNKRCvgOpa
yIvaVnCVPpI5re8FeyJNEaT7a5btcpffso9XiaCzB8dvPsKmsiCMEhFhZrgSFMwh
+qPKmmYW46+uZ0kfkK+uqht58BtfeGDAvCfRW0aXfK5L7YyjpMEZbsGJAxbauP4f
0ocouCTLlT9jqzKO5jj9BXAfSDeGBnF5swRQmyXJvK28n7af4a/oGN+nLJwA0IQx
FAAymJK5W6SwzlM3vohlaCNfv3UxuNCKasWa7+NkHdfc6oZUX9kk/NvPtpm4ThZ4
9DQTg8B3Vvdt7261jmTx/Mfhj8COSF+odcjr20/S7LqDNz3fKP8cU6bt0BCXfNz+
mKUAFj9f3bAM6nRTcnKL8UmfTOIJMz8bQnuQ1tpTSQwMVeMsLfPPFeggV9wrcyc4
PQUj9kmOuAIv1tO1TKJ+RPzwN2nvTgsIi3NfxJqHyo42IWSr3iR/4HWHPFmCBYH2
wjjLG1qQq7ia7lbggRB9DOhIwi4XugYFbHZMAKB6ov87RlPoPqY9BNduDm1L9fdV
S6IjdHNtZEMSML9/84HVfzLhunDndaBjqPCeNwnWh3yhhaYjSVLsKf6nU7owSOQx
EcVCbIvhNeH8dOM4pkVg/jqjROwUyxIMLBewt+DonhbjZx2IS6mpQbyAcAYWV2yp
JqX5iBTWGkIywNeTawtJ1cUsgkrOv9Rdyn3KyW3w7qeK7NgBLqLGRwEEA73vLcCa
jd+xFVXTNgjmmdSJ/x1oopDJqKJCIWVaYNAQfn3piIRWgH2/4jZbXQVbIRNI+D0i
nO+H7TMiomGovWLQITAO6W3ADZbpOMJJugb63L6hMRjKhhBXE7tFCFZvOLLz1HOo
9aQ6ctCdkLHf88/Oj4QkqJewZZ3gZ4hfO9cJWR+gjv6zGfqfelHYcRBj40AjM8MJ
jBooqIb4ZFaNmQ0L/EId66iJO/McXpAQPobivXGyLr8+kz514xiGw9Nd5Gz1hqVr
z1xvXgnlc6EvXaG5dUP/RY3p2RWBsYOCs62PqahJr/M3RsFUZZ4GIxpTwMHjvxG8
HySyccCRbfBooib6s7hMXdrvtMCPgHkgpKX8KHZJ0Z3PoKSlsD43HppJWwwHBEZb
qI5762mj/9qAepVipx6Jnv8JoSBeNRUV77aQurcUmxyegcNhQ5T70AlvSjgxXqtW
gYBXiLyJEgCHYictd/RkBHb0oG9wgCPhAIE/oj2bko4NREaQBH+ycMxXdeq3OAhm
1rXAQpr5daHGlyIJE7ih3I9m21nDOvkuA6FbUmmx6nCFxsarX+RyY2zVdBrkNumx
oOroeDl/a4+GoObeSMlD9LxHgo7vO8bQB9MqaJCH5RYTvMBD5gJqhMtQmLIml1KE
XEfqoAcsMX3yBmaOBMMqlDLCEAwEQet3KqX93uYL+u3sLtVfD3OImdYuwWCAuj7c
8X5KHLnTcXIS7+Hoqnxx35j0XtpioJNuhZCAVJWqN36oJ+l30Cst6HmSor3rFpNj
60oi+TdUClXSwkcE6qWsnpZKz4hEqGrS6i6rrgCtmfv+hrTzRhQDUr0y1HhkKPqc
V9+WDpL7gYiQ3UC0f89bUAldiHBrcxjRgO9rGgvLllLnzstLyhWkRKsBbe7PookR
xYs8XA8CHKNSyaLjgCa1v8uqJezZX0oA0LGi52QR+hW/XP2y4XD6pf1pBrClLg8N
0lAAYFjR0RHX4x/raq/fwbB7qtzbNqrd4rTXjJ3b3XOi1y7BLWaPeBF6loUwhx1m
PqYIxlvuA4TtFbE11ZQBf3YviHK68bM1Vr0qIOu3S+lfCdoehbo9rnt6NgBy4tdb
H02LxdZGEM7tUzlFSQlSpHEIi68gbgKuam7rrmbmYhUZIrTIuGO3UEOBHUOd+o+/
EQip0R+9WuLs5KEKqBGy4QVZTECOirU0wbVb2p19Me4aBUWG+I6hoOL2yJNDubOi
eH813Tox4cJ2sTkVNbqU7UiT5z0f9qgk6e3NfxeTGaU1+nI/+bQ5oUjOG/wPqIBm
3xNRSb0OP7JFoup4EvnBltnnWi4szknH3qRaZDEiwy8cqyVC34DUZSWMV20MLMQ1
Pj9ocHpyi3PoeySCXpzM/3oOIEQ9Upn16w0JGH5HJoSRpw0gmX9TBDIAIT6kGZdD
oi4vJfzcAeon87nqBJYYeNy5cKgXGNPFJVYcHkdN95Kmy3YtKoqWFaWaOkjJMu6T
h4POMdJ1BNb1HNGlAol6DcJ4jGmZhAP3kSS7lT2GmAnlG+X3hVmA0gyYW7p/0BrN
VGq53ALdemBUMEtxfbiTmp5AOr94WDO0Cubnm5zz0l0Dp1Wj8vP8QQFo9dtA40tZ
3T1HfOHacZIIgl4RNTnoCNko4tZn7KHYXewkFuKZbbuIb4LarLCaag4qf2Y4GK+d
zNob1SCFaoLNm+ZM9C/z5q3f76iiYO0A3bAf4yPb73c9AmpITIjtCYYP7k7Io9p6
lKYcwMZIwmcEnlxbddW9VjsYotOPTniJo4NF0Jjht4U6ZcVZeJGM7ywq9pon2xjj
v13Dp1h/yRQJK8UYJXHtUs1pyZY3kRYca2rVLOWlbNQjto3P1gWxg8Q/QJ0nYSMO
vCvDr/GqfBQcM5OwYcipfTJnv/3Slt71zAiLCNpKipbEL/EoN0IMQg3E3rjMugGx
qA76sGezvbxB4Ty4l7kb7gyeVNj0OVWk7c88HKLwYDvGbam9oQtrdwRsobVjF1n1
rHf4BAvgOH/XFKEjse+vfsqbFQ1tuZ8s12d11ECG4eGpp5jLtp6xq9uXE79zMPYe
AjrkvJStQQI7Fm49mrrZMCiAaIgVQxe95vmNQzd7Wuo8qwLjdlKrSUdtQym27J0Z
jm3jGED5LHRo/Ay2N3ugJP966LIFCmvOCN2ZU0I5uskuXPNmFLWh5b0R+ObUsR+2
WUTzmwXJdoYP8MejKfYeTvrGWSh7c7FQU+WRhGDPzT2Y0ohkh3Du16+McJU2cP7T
+00foi1ELidxeXP0FmaZk0RMDRixGKs5oOZwnzg6M58ru3+hMoS7rENa79J8Q0Hg
Ib3KD6telhT1UB/xz8Fi07vIGo8vBJKOTe34aeO+sFKz9PC5U6VZ4JIIERmHWc3i
+DLAfXLfPiAlB6jxVEbkoYsC7YUZBi4HvFUJtSCmaKei/r4798y0MKleXFUXi5pI
b+Zleu1G5qx4hriRxq9Fb+CBdHkyD8ggivXN1Rf9ArcWwBtw+ov8hoFPLp4DajYV
4ye5lwWJw0YKkDE9Ptufa77lunN7x7OpOyUpWCFWP/gSdslm7MkB8lu0EGuI5U7/
y3oyCxvBYasdQygcADggA7e/BDkxovKXoOIBvh7/AXzsYmmtURjzfHvJAJDbnMZD
TCCKbcrkYw4Ww1OCnv07218K2zQzHdA6FF/hWwWmA75QXS09ArBzIJgZ+QHZnn8Y
B1qn3FgYcDnb+lsKFbkdrm8ZQK8BbEi6Wou1VHNRjc0xrgYJyqExY3s4dSEk+IFw
58lroVsRXwP5NHM0QcuBFeB2Vdu24XzDcR3L4uYEgS5L7HB98Z+zaPzHS2T1EH1p
pz1cceKH8gPTlwSva7MfXGK+NAZzWkJ5LJAZKtOQilm8eUaOB0U3x4j/5Xfqecr7
U1cQWWPa8H4s6Wamb8kUhSa3rz18TR1wsFJy/3FPP41PmBjOyynhsYKFFPdctzCN
aSu1U55fu9VFsVJ2vvHq2S7yQEaHeVyaXQvixGgM3n7aJc4WiJ/ICqqUsE6b4bTg
0wXaBaoIvUNv4BqoKkAWnZmQehY5PP/XQ+K6wwnBlKV1MS6jaukpMfl5n6W3kqKJ
ppl6HFTR9W94pqj9a/ADiABshiEWegg+p1eN4R5xf464xBSQKLDbb08y6xr8GoTf
oclWXSQPz+9FD5vQWmn25kQa1Wmkkv10lBuSe25i+U7kw0YajrHXi1lD3juerv88
7ARujc7+ld0I05yRQgC1pEzrWYn6EEPgHoWjHD7rDhdZqgv1XvQ3gQfP/hHGXXfL
PuPzP7jJiiIF2k70jukMQex8+2bWFGNfnf6sldaBEINQIArIN1inRLku2RInXI2z
6CVIcT+bpbYDsGRCWxVBjpF5a6mRRCsyRvWhfRqdYNTWCtA28DEybgCjnOgKYQdp
sZUYykkcrIbJyYEW49uhTHEa08leGXLXMYidWqpFkg4lVdSNGiH1VL7eArCqRibM
KEY2PH4fZ7G3K4VSLGZG4xbQEt08jlCv+5l2lsI7Hmwh6rmzlNpadZsAbwn4xS05
3I+Rz+vrjHlz/vAeatxOeP32T3EINPyNrd7O0LAnTVKj5mPLW5WMscy3ABXAzqZ6
LX6bE+rRbUi/+QMdz56gFzTQMLWh5kaW8m0bL8C3DsiVDn73PrEpDhx2C2RlTDx+
UZJlVP0rutEuKkZBcG/Yo2lvWjZmTi4kcfC63xyVXXLtDVZ0JRjj9BPxQO8uF9a4
GkFUpWOQG6WlQvpfY498WG6DYpWcOUCUaPokBKbpE6wFWbPV8OrAC5RhsMLa/mGg
dItz3j0MSIbPKiS+ed/0n2MKflJM6Bb/IBxLEwrqrHO80OV6TCHAMxy3+drfZJwT
VApKskd6BeeXwp9nl0dk+dNfvjh32OY7F+RZVGV1k20QKvz8tvf1TRW0PGBUjaSj
KTbxd4IBVAgJYG3TEu6WeoXSR3ZxLw6J3D71F2+b3rBFGPhESMzmP03vq35dxA3K
Vvvk4Kfvp3NurpgG7gc5+CL4+7lZFWljeDZdghEukrRjbQTshO0J8SNvtaqK1aT4
ajznVsYDlAYvstz4J9GciM4pvIJ3h/TrVli4a2zQzD5EFXk/RFxITYBMnp2QOYJA
Uq57HN6689jfROi8CDUZfviR7MkKC25KneGy1qVO+Zn/Ev3fxEihfhF2ynhFkZ+s
BtUR6LOwNETbxufnXeuWlVvKFmAV9d0GXSTzj9CDn0mFeJV0aKfM1SsrvfyXcHDi
jdgPKlFL7Wfz8lEYfXdDtiJYYvMWC+yFnXYKAYwy6lxbE/mttkXtihobFQgC1Skb
s+pMjqdDDY6sOaBYicqAQS1y4eJrFT882y/CtJ0WeY1M7PPguuYU+Q0d4BJHTg27
hlpIeeki2iszVtyl8nP75QhzHCW4k1DmRhsriefCI32Bz7B8mTQYdklAQ1j/5k4j
7bHsIe9a8yGLh9RyEMXJIoPfz0TMsranvWk5idrOVEreWXp1puUzSO+tOhx7MSoo
gGdfi3vXrckVtbjx7752zjLuK+M2zn92x5Xi6DK2pyW/HJ2Bd4tGI+ACDCPnoFcR
j6OG8CusfoirA3WtGTW+/+10DjbvVwqE7W4qh6NcYYljAR0Mui/T1o89r8rhvZ6o
WO5u8tdP81gfkYIcL5oAjgedcyYjfBSsGUVrtWjcSqGUPM65A2Sud7RSoEw/0sNd
sgFIEBeb7BkR+vM2hTzSGyyv87C9CO0yPjjjk5ERaGFL9j/gqoAMDjOd/uVdKAvb
Rmz3BKUirN7AZy/8Q6ZS/NHws3k8oVk4ETDc+HOmd59/6ItXr3i+QN2mrHrRSKBf
br3JfrgnEQaQuxcOeS6eIIueYQSUXvQyy9BZyqc9otDvBck99gi28qAfPv4oaU99
IX0Pyq7qSYDNt1jYfsmtaD5I2b0arZfbGXC/oKzs2cWhOqnXO4kRm1VXlQMhiYk0
3PYo6sx5jFSExW6nmvpeMhioBGZeQIDXoU+KgiqSgKyBfTFIIegHhs1Uwf/mOz1f
bLLX0FJU5zSaqUx6GAGhkIOB/gr/3HgizQ/p3eUUS4ItZM2xBPbUlHlPAJHp51f8
Xv5j/RIGHPq1jksNy4009hllC5/cbaOKLDKQcnaZeocnWZwjPkOCPTF1WdNbmRe1
vzxArs4IR7sRuPFlmQysQO53nD/JMzbasJvI0WaXWL7iwVQd57LmPQ45RX6aOXVR
IIU2f9RORxKAmJ/DIdD1g4OMIooYCRDG6KPmmjbCRBcOXsaU7hRL6cADH7oLkOya
TCK0U05lokcqtFrvraa94ENWEmjHKv6RFoWx2FHLILROEXdfvSy3OIpAT9EQlwIe
C6Gi0RGa+6T2Ru5r3udxsDGdyP7VTcSyebjEv55mACz8PWVJLRQzNKPVuzEncuQs
UgBpmA8x0a66UwZVytikdpFY2N8j0zUioDUoDUqTovVGK2+KPzuQk2TY3or10Z9d
E37Q2mckfioTQEGGyrXhgpPHEMxC2hrQ2MtfHyWUrIM6QMqJi6XQwk/f75roflaV
tF2MwruwL9fjfM8O6N9DUOEgu/hghPEIYA8IyQgn6/zumD5ddOyq/5ImqUhzh9V5
o4ojsMTVkfMNxeXrYWygSXlaSMjj2F+Yd/hK4+pHJTke74BAB4hvtv4Pk3aJ5wXy
1ueTbb9cYCRiscrbD5Qpon2JY0HkRW3bWqRZJTF8zwFRazbd5cuDYYIFi7xnPktS
KKn7/Sz7G3LBxFLa3k3Aeu5v1plSwqIgjuoO3w5ssXiUQ6gY5jn3D/b8NKR2SbM9
heBO0kvcRXmTgHNshFCG6LAl2tX1eKE6E2cfTp3RLz7q3HdSwrBuoWaPXGLOD3Zf
3kMHtjUnfDAd0A/rdvI6vhjbxkJySoz2WjsFAmGPdtMQk/HTLHdZXTciaetB9gdG
S6S8m5NlItts2J/Ii8+3HJMv4Bvh30r+WUdAx3uJB3iQ8OxULddVqAw63d2XjNed
F7BEekWLb6E/lLN8qstwC1Pn2MKgXYXV7KsPLzCE8m5+JV1EYWFsRRJQdTrPZ16I
dYtsfj1kaQhZU0fKYe6hWtagFqRsrHtnVxL34c+4fCgOrPual+6FsiGelYZkj7cY
BrLTvmV2waAJj1MdzDaLsOqZHWkGERwVs2wvIyFvVCIeaqsf5YjPnyY0DUdrgnRq
3sI0HQqaXut05T97TSATredy5jcBM4/lpxHDzr6OiQkkUWDf6ZDmcT1bnjmklzoU
RduWmzMhzyXIk5aSF7JfUVfDcKZkouh1iCATF52Yv4mc10MxarYCnS9+wG+tq+bw
KINJq2E7489HBt5qz7Khp47Ek7UmULOAFyRVBP7o2ym/G4yUDiy+5eiQZsKIWghr
D5H6cWAP6Ks01u+TLhgXJrN1ZOKxQRxYfwfBKiBoNFh50eEmtshPXQF7WmEUoLAY
IGncrtPKmjTOhu4xTZE8Rhy5+gPjFhI0Pht6lRrS+oRslL5ypB+ZnB4su23T5vDC
zf+yQVPP5qJgevZARnMOgZp3tAoSOTgaVFeBO3vQRG3nKKPW/uk94hYsqcJ9h08b
Du9e2e+OaeuQn0DmkNlBROWGEhxqYbZhM12dYAetb9YikIp8XPI5XTh/3sfO5fjN
CYyP9OoDAh3pHkKfI6PqB902C0I5C7xaERQtCMFFyiadLVxIE00h4OaIjR5JZp0K
VFHcAACglnnpzR92qxB+DZ4/k61lYBIMdesK8O0lzGeVVqoZQge8np9KGZiWF/Ks
BLTzKKYzZI6/5dnIVImWT3yyXjZZCBilZ8ieaAd/yslQewwfJI+bpZqeXxRcF2e0
g6Vf8vCiItiSWro8l2xmZmmBhFZxlK62tpFFeP3/F5AS0nYEWRGdzbNeGgRew3Mc
undSFk6UH9ZdoDBbA5RXfJVsU0ZmeDLpf13l5BmOAz3QcQILVRthtFSvPGJk4Zsj
ZKDLKtYqnyM0VOcjCG5JnVOjrRWL+62esOJNDKSCkxvRo5SvmzXXrONWevu51m5u
iYQTQeLh2+YhOT6nCA4fGrNazP+tBgWdxMM2B2jTKJ/kpE/jjuENMfuWz3Bx1yMh
3jnuWNFlEO+FXjl3nD+5UbIROTYXrCAzl73a22y460ZiomJRCv3MsdeZwQ0quRig
2AG3ujv01hAbc7rQvL9kigcCSihcX5jiZJAzqdeDcXLS5pA3/UPZoLnYYKR5cHSG
6e4NfZI+AM3pZLq2vZX7sM9zzmArh4h8zQw2Cs6PPCm4jzXnp0LH9IRKoQdNqkDl
KYRJTRxqp2aeuV3zallk7UuCb6ZqO43SWjtpLsr2U6UAbJ8Sq+JXF8GyU2Tufc7n
7whSJKhcnNgc+9KZ2wxEkdlhlG320FuFZ12jMPpD7hd46FBH1b4JTMh9FUSRkCcF
NC2XQy/kbEkpAc8y2boda6h4n+JSagAFPNODUNypQuhYx4Vfp3D/ve9Z7BIhwLBZ
EUtXSw7xaz83lMaYLweXhZ8sLPkDZhJurO63Ccv031TyVXEwRtRZ5fd0UUbgXFJ0
7dXZnufjtptzhHMvqGq9D6xoBE1VN/w0jP7tcwquaz5G2uUCMy1LOGaZivtjGyLr
q1ZkkVClCcTvYPC1a40NzgPm18IXi9qZmrtYwLJvbVOzEKP2f3gF05xPbxUDcqT1
kN/8UcQaVXTtxnxMpb/2L6Iqarp2eLuwWT5YxxWZQJHb38VnD/yNfau2IyotP52Q
k8n1HvX/BHe76TemxkYIsxTu4BY6RuPG420VzaBu1zzQ8NG8jwi4FUs+iPWtEUHn
pv+KJJjeoVOEUCLEuwH+ND5q6vGbZOpJHmbhGsQBbzyHYwMjbxzlCoz89pDEyeM2
3KHWTyncjsuQDkWKigtAuTe7pIis9CUU3LDkB9mJfkcmOI5Hbjq22dT81Eq6n8lb
ZCp5rsV8z/fLfupexh8EHOKL2RqHHEw6/+wl3jQU11meOQ4geP9L5fPyxi7zfDyL
4m1/AI0ERC7cqln7n46f8oZK90ewWflZaKeL71i1BvH9AYirN46/07mB4MzZeCoO
UN9vMNnGcOjLKcxFQG6K8LCIOFSmz9LtARaU+ucj2Ctryu60jTx+wEGhBpWIszrO
/6pf5dt3JwWiVZahYXCD2Y/i3imOergXjp367fTHtNjIcLmzJFiVvlHpvvrA0PS1
Gi/JaWtkmiQvW5uIequIwjJBx0n+5iAgtYYEyl3ICoSrFgIhXcVu60sAyhqQh9wm
8rgOzc+Fe2UtPs6IPAUb1dSGXEkTRI08nSYGz5SncKMRfmbkCOwmqi9v2vP8PNOc
CANFiDZrXZBmDqqyGDCUSjs+sI8d0rwB3GMnSZUC86XBgiOZEzgzVix8jXLsXOTN
HPHQVUrK19nC4m5ZL5rybSKbrOsZA0orBDT3WklnDSDOQgDuA4gLamBAJM55iBGH
+jKWMSIht323ZOJJJyyp9zk+edikVYBR/mTjCgbtTfzCc6DmUmsZzfZR0o4/wP92
ixYLoEuEiTb0zAcp7aNX4xcCzeC9hUsZu8XRGoj80QP8fpCn8da5b8UiAP5TR98M
TpRBInfRRKyoxzA80WvraNwEi1Ylt04z7Te8WhOQy5vPZjKWNhQvSHuFvKGF8h0B
i1yLGcTBA0AJziUwmtVOpNzHD63cra9PtTRHBkbttcHk5vHhnGE6+E6HznFqZRqn
t0FvcdogDIWQUaWd2zoXXxoElqYBeooGtAaTJG8vaCilKgxJPPXy9tK9Ffh6vku0
Pi06NUIhvugnuB1UsPgpUqFMfBRVffPyV6pzGTfShzIi/bf7wI31VHgZN5LeK7Q+
EechbZ1FPdllZbRbv44P3sjQ5+7DCjN/HdKm6yYtPCZLEhxO5m+HaK09B+s3I9r0
bfN5YMMdQWx3DN1xqYXeuC2id89qJN/dpjZVECrmWAorRdm6OIrgGh4n4J/z8BJU
Y2K1NtYZmxKBJ4Kiii9D8aLFmB9hgCKGRxgrZ7aXzQBE+oJMHBWaLO46vRt3PQm2
5QJmVIdgeeBF3g6iosCDNHk+kUef2kQ8aMKuwuiWQ1YbNyOcO06DXpQIaav+5Old
SaUyLzxLo4MM+uv4s/ZA9+yFaHAb15+z9pwHQI5hpUEy8j/5YV2OH/h9y/LcYAMj
/IM/HGUDniXsxgspjxt+pDDkHEcSIBB/p4ja11Ab1bcpJT/h8dDd5oPPOe+ioOO0
zIVmEBcP9foPn2/OJ3jQ2mtsc20n9lLCkcQz6JwQO1s0u9nMiIfd6BZjKX4Somuc
JJbs9e9qcCLMN3C14nfPv/tcyhH+HQKGYwrTQ7rLeyTeEynmvJQ7uKj/ch/+IYSj
9NM9kY1v5rEjjWtgQGAczzZWCNU7j2U2eLMU8viq3wzoiFkdfG27wRs4y2EzOMsN
OuCZ1gRYf+e5W48GvJD9zO5wjCgUDzKGnx4NiFecfmX0dhms7Mkfitk40kFkg1F8
Vd+mGctD6AYLVz9MPRoqR4g6ilNxZbRpVtk4iGL15I6PrD/e/Mzc2qYh6nbrwOL3
CFw/hhCEh0uTAbp/x7A8hBWjyUKnT7fgThI4/XDPC+7qEgZ1b3vy8BAb3taG/VVy
ZZxwnZciilplHVk8iwdaQL7HSoKuuBvFCf5caqeCpZ+d3GkI8bjenl3JJyLJSS+I
15DSBRkOo+GeO56mfAqvURdgJleBwbdSkL3BxZqU9aU38NTMc30g5Ihjh1pdkIP7
bPnEAQWTg6uiKHlpmB8i3bWF+aJBaygIQjy0Djb2tBYR0llmp/bZ1AplB0Rw6sH1
i7eZusjkxXwGpYsMCI+Y+ymmIdcNxQ5FSJrTQItlBWT23KoPoIa8t4pKdCEBSHnt
Gn/Oj9bQrm+SaLcWtP52KfS2Nmwbibhf4VVl1PPvZsQSDZa0UAu0Gsqh+uXrDbKW
T+kue3sXqpcT64n5pnTbUr75jxAEW5f+UjHa50ER2arCwIaJ0Xxu39acPjukhzEJ
Ucu8JUxN2I2dtycTOh/nBy1Je9PJYJxOBxDnG85N97SUXJEIoqQEc2IhrhsHSPNj
NwdRkGjojEEaoFA5p5efyrNwaUNPipgYtyugx5LjUrhnywos+GT3yLOBNS9m0il6
FPnnctdw8ah2MIlFEB3h8wURKa2gPkaqT6mJyoomrMQrlpDdVArWV75uTgUm0KUh
x4Bru1IYl4KIif64lywD0l3OLceNvwKz85WbFTwySIdDGF6c8F+IEEE/5ahN2CVI
FXepHYDBY/EFF8Wg0L59c2JqBecWNokOKg5CNk7Rb/fD9g+MnE/Wj8+1He+bDC+F
ahNHEIR4X737rREFCSUroRIUj6p7p1ZLA7dGoBHBYs8fF0tgo2wmuWzdEPkEGiFK
2e64Az4UpxvVBa+N3oIL92crUd9y6xYlxr1r7xrKCTH0kYQ9+Uv5qomflSzY+lxk
Bk9ggcrwfNm3+hU0JRPIKwubx4ywq5Zook9Z5guoSHXVo8OX2vXO/f9W4e8NDnsJ
66J3w/xJWKqAwBd2CNdCAhpZL3VN9N01m3f9Kzbp/FAUVNAQ1Ag87C85XCAAMNQ3
6LobA2SQ+UTxEQEzf+mocEQshuXRY93gjuCWIPQaRinjOdIn+oY1Yv7pHbBeO0Wr
VF0p+CtajCmzfe7rmWDViebrbgY0Oa6KKj1I9c+WRFi8LofTiKiq61JMqowzmA0u
eBn0LAMvHfdX0IWkleqmieULPmRysVK9hSDf/KMJjMrwhYF3fby40lQMMyop++OW
zrJrQN3clbZZH/K3ECotT/ptqLuZyh6SA9nAChluNBwB9an+cZa2uW56g8DiXfnf
zoGrZB/goY6wRfDslZC/Gx98kG2v+OEYcUHy2kFX15UMtSjWBM9IFFPgu0JgoDmw
YO/UnvKxrKBJmZPlJBAKlrMXza5e91+Mt1WCpQaFLq96DBqn7DXHaegtgZBtFmOR
sRHxNZqOOYg2Mqrvp8DjSTUYbv6bqI+fV7kkeooROb2vBcBpHtSx62oWUejCFG5S
AuFaulds1hP/BoOiKvNl4DHBiFQEHoq1AAoPlX1uzI6RFDLsKCrANkj+FQuqGNHO
hYTVueMVtgAnvzwDIE25qaDJhEQC/0VY82s9wv7Z0IhlNvWvvGDbl7knZlLFxz41
tzWSSRv2yr/9c5RsVlxnCIE2MWfVPmWzqUzD/EcmyvlguX9pz1vq4Rc6DXGgH1iw
3Jz82AFQod8Rg80XkMMYgf2PJeKjI5qm9M2netqOxFHmzXMqop5hkIxwX25qNwV/
6TJJEpQ7EMgumtubOsVjUc7CAaWqM5PxtpDAiTdkd6x9KIHh7GEiALV2Hbr4OChY
sc/e+izzmjkDLGRRI/1gurFYVdCnbQ/Vy2rNmZIBYzGir2Ohb5Oj49j91PJ78bUL
uPe5+mI0SOpkWuJ+Qr/LbuJUd69RGT94SsEA/4wp7IP++F1bbic4S5HCquAtMawP
ChUiWmu0DHAWhX1xkaMosz7e6mhyEEbh7CVSagRqONLH+lYr4V/Q6kqab8nYXO0i
nmnATyUJM/Hn2ogLckEkc/GgJLsRxWT5KQuD0JOY4iQQFbLCuNLaZujwKoPMm0PL
qlWUQs5rEwMfD/MPAzH4X66EN8KczeKUKGcRIlSYyd3Sqk0wnnuFecEBgtRTfrDn
hbEP6o+0XAcQQ1TBFgtCAPFpYOIapZpYLfVqYszaOtweG1ycdCEDxO1HBMV9qhJA
MVbEkKFrj92IV8pMgx9bHaROBzR3bZlDiySvlGMp06Nn2t/LBbzUaGZw+ejTAcbK
Y6JG0l9woGqCVknxMBxY8V4HhQmS7O9U4L3zJmuiq7ebItYuHbndPY1vBjNdhzYx
+NEu0ibIp2c1F4gr8bqu7MX/kdBPfcu9bUNRs980ZyJnzWD2mHI936SfD1c2yfV6
OI0j3iFispSaTJt8aBACyuV5k1FGp9s42mCklWVwIDGxUP+YFT5DQfza/smyak1a
pOhugiYXTgYqJZ3MzqR2mv7qOgFo2eiXOs2Ma+jlSDLTxtKE+KOc1yY9LBHO2AvZ
/ULs00M5f6kvxFu3Og0lrga7nz3NNRk9wVIY+/xksrNigh3BQm+8G2NaLCqNGmV/
p5fzbZyOusDY8WmoXa83gYY7GyZ2xqV/jDpiuOdo/uYAyC9jAQklf0XDbzR8m6LH
ulOGqRfSogMq0vFYYaPPJ7Ziy4omyvhOuIbC92JEUbBLFPvlpoCB4TFMDJ3EIv8n
Kp6xVR3U65mLGUjnN2C4tcETmKH5MyzOe+kwoNlLQTLRF2j7Yxwl+uibhBenHGLW
bjw6mDZP/LT89RasALcy1aVtfKZWk4SMEoeAA8QNl5PBZe52DELv/XhKBAcRuwfS
V+ftHPNI5vqPtV1zXyezZtOJ1T1iJPTs+yL3tiPyQ6zSuAuZnb87wMlCId5ccfOv
qyAUJ9RMYaQuE8/35momdd1gfxmQAx8WuBBejhb8GEfMri21V7f5y3aiCUKfqEBA
WFfMWA47llxkoktyICAeygLfk9YTsclQT8DY1E8u2ji+9KHdQeegAMDJzEix21ch
+qs8+8Awv0vL1bUqMaZfO0HBvrGYELajLr8exgfTsK9PPjmXYwkz2BZUoGjr6EC3
FoFCRusIVpaaRq//t2FhBGUb98K9WnesRnIdx25Pj4HZC9M1t3MAhdQ70J76kbrM
LeGUYtofKMqXg5h5+yA3IZyCTxu/K65DTOW2kaD79wv4bhk7t/naF/z9FBpcFG63
m71ifZHndcf1JbMVhuiVETA6CkxsIXZbx2WzEmQ3CQB69nVtEwydGLqFkvcCWiTT
D13Czh0cTAIbOw6peNUCZ9BQLX73mxkWbRdnQlOjK3qh/yx/tHtXUxbCiFI4tJV7
sz/jafeEKZL7xDieTB/ecMJ+XQxULJ1ERYv3PXTmJighzDP9JOZ1BfssmOxcJa4s
+BzP1z2DuTGsKUaEQQXeeOzfPLuEEJ+YMFcvCQFhxVF+2L8rrcb3DHnX9Jz6ey16
JuL8IRDboLIiCK8ddfgw/EKHaUI48WPfUJWMKqj9K8gOEjLr8hMv/eLn3ehdNVhf
qOU0b2UonT97Da4GQvFk74iZGx+gJL+/SKMfe/dWxL4Rb6tLg17IpJHA4AoLsr60
RMuoPwvQdVHoZE6bwDczfC/3cOZsHNk20tHGjwShe3TL+LgWxuMc4/EKX7RKIQjK
FRT33kRu4d8idWYCbVdPPllgsZvbsxbHDp/z2h8VFK8LdOreua6+RVmc92tCBnOf
Q3X695ABf7S27abXqqgZDzJHYbhpfzC0Ey79ARA/v8QOS7wpc4ekiunbbwWekqsK
Y4JWg6+ygRHGXJD5q3+H9Zo0Koszh6R1VqFSMRAjdiEamBiBqA9UrL+HjA96tkEY
1kmMRThfQX8Lah6Wf4ifQV7HAuG+F4jb6KPz/wji3eHCHIu7r4x55HeNikkQJoQ7
AmrAy5RWqNlxaHBUaBFdh7PMwUuVqmzEgjLtCcJlAtlYQI4TzfMLkLw6KHTJy+si
h06diWhlIqjY5aOO42FwrKs9funpgq8z3TEWjvftHASEj0EK5f49O2zOXMqLD5Ms
BRmwYphwOCGo9CItuih7mxV59S9vEp6gXRroIudZi9EAZeDgvI3iWoC9PMVNbKaM
01pU+JcPqp2uGWb6O6J2roo9zwAZKZyAGru61JuwUOF0WbhPGgrU9pwD7gMlafzc
QhTHfbTYyh1aQWtPp27DIs8g/WJlMPH6SZPxJyCVKbzlHsUO6dSNhQJfmyfhSaeC
rDNXkWDl9d+QQpaHQexHAiIbmeC2nW1xJ0VdyHVWW0lpD2Cq1dDNdleJAZwAJvmW
9NqXGYyqnrhs7EGv17cbIukiDJwYgruo2+TXmmwsfZEadP4IC5YW6yrU7dWnVhIv
SN2XO+HmU6BAQvhRIMChzfFde4zeuh8qxujazTAX/9AOnbq+g10N01bxKPrqe4QZ
P7eXI6ldAb0IyGJkxWXNGCPX58/GDHEybeXvU9fUP4c854esCGJVx/huqGSlpmmY
w0A/dHNqDfLPN9NJXN+zjvNnYHs4JgoXo3xuaTet95Fc89qKKeFjMiffPLyyVXEJ
TVNtwV14LH2paTHuql4oz39R3Hcul1soRnWeblH5W5p4CRvuCxA9DIadUccqvnms
GEviAmVV7XBL5OzpoMbtdYjc1bwrt7G/4ybpbf9GtGfChd2sMjQF4i6YaXKShWZc
gdKHuiY5zTo/46SckluTAx6frug6KV+DrJGEVKcJYTlHaxtaRk9LylPVOSjclWR6
cylpQ2TUmLUtOi4ymPUrRUhHRZd5AjIAYomsfxPVLbUwD5QktXnul09O40y5bOnu
qhUfCNWZw9WqI4i8zhqe44t4XuuKCvtAhvq+v3MX92TlcACc3heAxoXuIja69JlD
IL1hM/jNNp8hfI9JDgmwWrOq9WBFLPnW5Xi8tSuJCTbchlXQVQa2u7wrAzsklBXg
DqxGERzPLikYq9d0Uh/WxHdrXHH8Fu90LHdJzreNM+ASRx1u4q7TiitZO/EP+TH9
I7ji840yrKbN7D+Lay/IOwX/bUWx0lgy20Yz+Fk8RSNyorVjhBAnEMBe8D40EvKV
PzNybYSwXO3L3SBlfj5BbZ3TQonf9zw8dE+SR/Ks5ACayaHa7OQS/trZ88EJ5MF3
dBZNtdxlukkPYCWJ8DiWGNQXOpxiAlEDFG72oNL9ESXlcz/Q+pDt7dkqizi46pHJ
GKE25sNz++AcBKDrYgSgVJyoCwYIoQDydv7RSQhUXrYVRrGwA134BFHP4n2StkEx
GK3sd1ThGxX16yQpLgQ4nv/lnVIaR3H17vSIZFpOrc3F8ks+H0edMd1SWSlV2+9V
j6NrwwcWrhM1dtZAQgO+HFN/afE3NQJKNfo/+GOQrMsHxSZc+qwIRhMGGLRA6lUZ
I1uxrhkg1WctEccmBhbUTmlQGtglot/equQHloVnCOyHBHc9S/0eujm9nuibxxbt
iqGGWJFkLDc1vsGeBLZdOvBpkOAnrulSiUtcxZda1FwqV40+3OcoE4eMSZQOP3La
jx69Yqo5AwqR7vKOrRDM17mlcqADBd/XO7eNNvABda91ETaZ3Do4okH4jDfNjDsa
/41pDW4lyUtDck5IY1PfihcWsfSuFraJdZ8EmX5QDxGJZ8mOLRHXlM9L37jkAo8O
3+HM10vdaqkQJoY3nRbFW5daQollNU/M10hR4ufYqbUWJffj5lZoqTjanHfdbvBO
uEPU0esMXyTejTHefYH2msKXSFQ0WacTK1mSX3jnOJskoajpl6/IP2Eclo+QlZi1
03VjCUW4yCWgj95pEE3SPQGJ9hHWAHZE7SZYZr5aVAifCyV1MXqSMb/jQrjL3FyC
33FOeo3Z/2PrrEj2QDxDCceFpdkAm0hvGfn0wz6r537ROsdBXwJp5nPAHQCODMZT
ApaA6q4/8N4DlmkomjmzW+aj22Bvf9iIlRjSHxPkloG5nnbhoJ1UaoDMrKzbr2s2
UOdISjZelxdgk8+Xt8BauSALtsr3vrHPsoo3w8wUc4CXG69oC9P3xPREsCuiMDH1
S6klCIFJNEFvYVuZqSeIdczmCtG66JXWJrUG7OqrQQ053HzpAA8laK/PtN0b4rMj
bjHWeKk5JIhDTyqe4dbH2pO76aUp2/xJkXY/mhFxbWJJJiezVzQg1ACoSXY3M3Iq
7K4HEP+t6PTEQDHzUHLVtKvIYlHn2QOJIJkpN+Z4tkLhc3IB63542/1LPLcxuYOt
6k8dryEMdlk1JCf5YeVrVKDoCc65g+vvVlbkzgtqmeHxwZjjPoK8/ITP+/NR8QDf
DzA1TkQBVxqeruRi2NPyumnqPJegBPO2ghyahnjRB6H6MYk6jRvxpUdC5PuCMeyM
jFenEp+J/GRvbMlm7HaGgNcI9TU5BNkmwfH+mz0B/r98UQi3ckfejB5ejYejvHOB
KNIUltjPcwiTUgIhfD7U+KwdBn2Ogiy3ivunhsfQVXOyWH8OdxcYKrP0iiL8F/o0
fv/sN/oVoB47CvrPJ2/Xm0CdlP26ngnyWmVOiDDGRgV9jbt2TFduvdROXz5itX64
XAgAoJAxqaW14gA7c1RAm/6q85oHskNizkbCI0pbTn7lSrJHbXCyT22B46Fk4CVj
ltK04wtYioH9+gFnDFl60cR6KpOdl9WH1jW3VqX3wVR+iqm3r3+9P5tgGjjqQfnD
OqESadfthjF8bF2AqsA9JKTomWaU5n5vFiMS16yCW6mqT+O3EaTNSXrubNLX0y3m
e1VHVrq6QPNcV602wLpp6VuZCLuDh4tjLg9GDc4A5xh5odq3M9XImXiD5n/IS6Vr
zsxuKCBPanTrnM1CM/LxZn22DtAhx5wtUxjAIILThddoVr8gHJ6IU4diK9bXRJpb
ShGiqYfOFe5ofQxgVKY+de3X60AEdS8wrT5PpE3XgSRYqfWJXBOeSmTsrlfP7A7v
vUAs4oXU7vK7v2ff6V9dZPfiV4SpIQbeZNo/bk7YaK3u46XtvXNA9+7QjSJxk6X3
2IU0bIvkNZt7kzuQbuF+E3Ag3dCzhGVgjs3j5kctGu7SabZO4ubyJ2nvSHYFsruU
mEL4JmQ990SZNwkeh3/QXNO21WNGxlMZFZO/Y9g7VCHN35eH+B1nuUS+uPDT0lFw
LW5N4lv7N/QBxgMycP5yDiQfsCyYzVf2b1WX6FCSybNzOY1H2gbHqiefJH2S/aO6
2FKW1w9R33tD/omouYKEUVEWxQZ+gKif17q6zhukk4NJZo2gbcob2zLO0Xk+hFk0
pdnF3HTPdKt2uVMhNPxHTe1kBgG3Phuib03quxmyGXjFX5lazpYadb7yGu+qGWWQ
2t+M2bUJSVYQWQZO1VyY0BzxHqZTne1C4ZFgp8uFucOOgXXbf6ZhJqxDM1mR+Z+I
GCmeAcpu4q8TT87791EIIDlxiFAofvMnD+qfs2wcC5qwa0IywC9pQQnBTTA+qjb4
URQpx1Xt4lzCrSmbZDop9TJIgyJRkcpYqBa82+xVDI5OUS+sndMbSXyy/iqLJR4p
CYTlYA5Tvd11tTshrxfMda5fz6sKjy6S+vDHEOUNxtdvVt2I0LChkoMNoYl7avM7
Dwm79R/X/6mMX15EcwW/WPqbZTfOTe287s8+56cxbEacQbF89vzn2SW0GTNJ+STI
FIdIZvfJzddF/syDCsmDgLnfHTSW9Xs4A6x2ap5vVrl8lOB3xZWOZkd0m9yyXVLl
HSfYDCFGxLRa9TAVq8ixKx1xKwep1M5n3wvFrpRLIp0Qa0sNM44AahEIYKJTkcIp
s4g3l0cZo6mc4zUel0xBSp6qPBF8Fz4w4E7YI3i8YcAZtcKXYA+1t6c1ut8KoTDB
jjH6ZsI8KdPYfB+y90CHmAj9Z/vvtJM7fmX5803EDRkxyvSfli0b+XfP5k5hHp86
hME1YHVgI3IzqwmhfpbSQiC8ALftgTicE7MO2qQvIGcSAYeIf/Q7A/jyOSyPfFlf
6HnCiaAdLOL9BezNnWTS179w5tucUnKSGmKnbJ2hIEMRxssWhxLkgXhpVsRN8WTj
a4mcgHCgi3J0BvWfY5LlPjwWcVXJVXEgsPK28FpipKq8OjSAhtfYYP2Zy3F+jQQa
vPdjeBXn7qUgrYYOC2cXLwoSX3T70IKA8UfgvV8l7PiTtDuGXl1AISTO89ur2XWk
9sMc67YGCehW3roL56ME2TO4y2wgfk1lzOyd+V5tuR2t+9MjYdovlkMgXHsKeeXH
Jh4OkaEFCH5DqHI3+ofcweRw+Z7NoBaL9USxS6OEmOpgCd9B/HJ4o5PiQ6PP0RY6
qQHgoL7OcIry8oC7XEnkB8vx1Y4hzmZ1Y9sTcOX/had5/cPmBBiaGh2sA9njYch4
0bPhUPcnDB/mJ6UaQXmV2989Ll9ByBL3iDy6a31tCmmsv0roljhTMs0HTLJIutNB
IC8RaKI3vBmCS0xvP+S79S/dc5JkYgjbGbsKkiSTVeyqnLeV2simDdBBQlKkIEJV
yrDrIh9lI8xE5mNfNyuzwBE+ECFlb7LFlgcLLBPXQS9LeDsxC5rrBU11bNFmDezC
j1WX5Go1mkbWLUg+Okj1mBFUOlkhnujbfBxX0OET/TwJH85vgSQ5ib0oCmKIhjxf
O849NfzWfNkT9ADtJPa+9dSFQ+N1h+u0qmNlLOC6ted89kcDr6wjenzlrRiQQQ5L
5QbZe7fZ8b+iz/4OyNO21GR2tcms2gjjFUa/4ro+TcEh3CJsLE3FpiliKUMctl+l
8kLxNUFhk4KgZE+OZt2XmdSbRq5z6U22CgHnp1CaK6Kn6jezpG/MO3COkuYTRRFd
b4S/01bfgrxc79A/fpoK2YJ47/t8sp71JXBkPdErnz6LvtyuBxIHz62qudqd1Mt+
TnDMK6lCuNRP2tiaQpc5PnaNya279JrdQB/AJKJiruiJXIe7+9bvgiQSlC3m9oI2
XWK8q1eDq1EDAY99fATLVQomSQhFycDCMesdjNePzIA/6iWKMq2nGoB5HxLqGsPm
3L8/PW0xPZsgbNQdx1mGWOrHw8jySsHkiIZekp2DV3U2cJ0hECVG5YKEUSqGO/Eg
PgAWlC3q3JywRFg9oNKYkCLMB/e1/nfSgnnIiI753VtFZ74jXjzvPAGaTtVgAU4U
D8Vg1i1Z8Zk+ZzWZlG4YjJzZ8KxoXrrPMH9X1/hnUAUXNe8D9gLoTbrNAwG5bQMY
TEugcYVmBbToklSxnrCWHc+0Ly7PQ4PwjGQ6yE/Ekxro++Ai/S7fR71uKnW/sTPN
STAut5FTC/Hy5MtUNvvPPUD/hum1VIGmEEKzQiEGDx1GZq0vfRCYS7HfYt08T1p7
MUgHFUej2AuMP/Kel+11R8lRljuxk160dlifPWk/J1B1EKcJou8ajLS81kbEPQaH
0sgu5T4o9t4Ab1tKCi21g4oUzpvnq5Gagh/6/sqEi+ZJlw/WiUmXuJ2TnRIO9XKA
YDcJUNrM/iuj3tcjlmo+0c7qTq5WbdPukIGz8gakAK9+19StNFN9lUx3JSlZTkZZ
rGHptwOtUrqcRUOnYpuWC1daP22ZGdrdcpUAQDK/U4lkNByHlOk9swzza2Y/AL9z
HKb7FpmfELvtP/DEtNqpnx5/oN5ICJrTmxN5TM3SKBbFRLvk715G5eAMMTRtwEiX
DRXdQ+FQwpY9gWmsmDrpJT5npyaAvLvYAcLB/L+mi35TTjHNsvbWAes21JsfjrlQ
KmHw5NZDIjyzUaFrJv6GmSufq1nRMTvhOoWiNGPoE7fQFrVxsa48ZZ6BNfmimPia
giBrm/zuYGxRH3tu58Y7tWD2yaWDZaM9Uoyt9vu4kWAuJAqkiocgBanX5vOOpPF9
mplEkCUqH/QVjKapvLHxXbB8atdsUqFl611aPOCWn/eh/rqFWdScxV9OwQdegdo/
/voDZMAST/+TSQ7kj3s39ysi7oN+ScIkMhHuEmxPyhSisJFgaQmE59s5BoIIVwfX
9qM1WYisp48W94j7VBeKa9AxDIhuH4G2nS2tLJ6nRSiR0q6PkxMNiC4uQTtYhkAZ
8wwm/x8tkJpMFg0VoxuVL3RfGctMoanSBxGis+KII1zDUwm/5UUcVvpy6F7//s5w
+kdxFnsEaz2aG8hJ16aH3bSg0Jsc9kD9N3RfErHTyCfZ9uGnKRxYh+f+wBDN5hoX
PkYZApbfddAHm05kDxk5vrK1fCrG/xM/Das+qeVddqRL4UjG6UyuCtNjUB37j5AZ
eAPp+6TlR3g3Kyz1OidRqSjiTnHeGModBV9kCfkWPVSzXODxgh4+hGCqPME02Rgx
bR6CMNL9xbkfeb+J2KFWdOdSmRELYd6/a6BVcBD/rmrXj8KgtlIRBOLgmUe6qryp
5o7YvU/DiG1wUxJ4T9oArv1wAz4K0jhv4CUifrE1PqwfaH5MiOL7BvQ++C81qWbO
sj+bJwHfStwRvip1Rzye2H18yNnnPSUcAB++Zf8NvJRyTDw8Fc7g6Gkrg2qNFxSL
I4BA4ytoZA1PVz8qrFG3YX2/vQrR0Sl5lNk8WJ9++ZYuYQOonChm8DWcf7/M+1IX
xMTcTyUgo46O1heQ0+puJA1tBTp0nxZv2CYuxfDKal3Gka9DlPsC59tLBfJ2gMZc
tch5JiKof9eTbBv5Ni7Q/bcNysaecFqTN1SeOh1e8lS3uCMJNBskwlY2XjJHImUp
D5EKWj85mJdNcrV6G5/b7EfceGqqZavkVbk+SEil6qnpQQHR4gWQl49Q4ButKijf
2aWeK017uOq13cU3J9bw3j2xlsi6uFgezZItWyfRLbTneZogzys16RDMSmjkHgG5
xj5EvJCyWxew4sJz8uJEBW9iM+DCS/kVrN935jV9CeKKpF3X22n+ToiWdNGpoulK
zCbGGSmYESDlVcuUQdrPus9vSoH422dmfFnXofLstALwsaD+i9w75AAu6WB6Liyd
YYwlQUzZdRJ49S5G6dDZOLmHxsEhbMx5KLb8pZMe0Zf8et1sljOzvrKdrFwk+lOh
6puInV/ZS+JCuBQjLiN3MYKlzYqVcTBI1N0gLtRoh8Lt1WxvW1Nbi02IUA+9V6ST
Q29/yFFdMo1A2iX1/5E+eiEhag8aztEgRsneI2hFFGuQ2Pu+UCNPSMdDFxZJaeqr
Kfe/1HYACCrtvAuptvZ183Sv9989Rw0x0PDrTyzRXdcachA5+9zrTAT9H9OMFWje
R0AsUL81X8oBiehn9l+xW4wJrviOttapd9QX8W+PJqCh5xFreju828dValjCWI/x
DHVMfMkHv0GwudTopAR48IAJBuOY9dIj1agyVVBnrKvn1CN5WGOGEqoaKq4ysF9t
1bzPnQvXpVWmbzXM81pJ1XeLhrp8V/VpL5HxOOyP3Zlpu20s16fYeBu2KahccDXl
wdCyEuIUmUnfkkBhWE747Ek2XkO324dkazxQxbSMRiZqCgq9LAmhAC1AJhIiFvNF
quvuEcAHU53JLevwKKMlf9EN3TUYDUfBv62qnl/ZV73SBVOz3gDwF/uWZy595jJ+
P3AUdeKEStKAP135z8vSwFVj11Y1dq5d+2M5vzYp3JBDrGaC27cgPleVlQaxPoL3
hJR+9evdiGI9ugG2WWFQ7FhJL1/rxRNowCYbwc0JXg4OgRe9PqkXAnnEuWMFB7fv
CazuAxNDFwIytaXWJjUFAXFZB0x8uDew8kek1SZZu2bKAc3RI4YizLXfZ8Kk70Xt
prMRD9V1ltalEjGv/rwh8lqY04cuT9zlB6BSHS5r+A9snubYu4dBN036bLdSpLzq
EiU5FM85DZVT7ZeZ7fG00MLkqGWxJyS0DrGM1L4zfj0XpURvYfeRTMltXKGxu1aQ
NWEQfe6cDi7HHIT0RzZmf5DOBO/bIOhS+K6CePThMVxSUNNaCruRSjDmxcEhaksg
2wahttVY0/TgSQEohzPCticah2p82UhdwDyQDEiRPe+RNyEm/bvL7to68v5/Peau
BInxKKc+QJwYwVGuGPIXgjnYfMk3ep6YfaCWfx+Z9Ow815+652RAG+1uQ7rHS4kz
x9FEagnv/9oJlDAyuPnkOfcJte/JbgLCnZPMEZrZPQEwfnoiX0v9CnD12241Th9a
Acd+VFhRrFcf4fnKebfvOCFQRSzM/SVawYV8Xi989AaXF9FxzNXkriJMDWt3D2AK
mjLXsBgepYZvcUVU4NqoQiwOKFvaveXku0thKVIX4uKZZ9WtyrrxXkIYL/fg1y/m
YQuOfCD27fUxmq9wDy9bKyHjkvqjUkgFyaqlVZLG50omkmttjTlIQKMVwM60kYs3
xZJntwOS3UvVnNVWHDgneDlU5qOl4JkUTT6I714DQcoCVALUG+MFGUdw9qhQAMGt
PA6vKe/NmQJOmOWaJh5Szrft2qY1QuY6bLAWtCeJ0KOxEBkEmEkcPjCz+14EdMpa
uLU+qhDxJe5GxpBjMBJauP3olIQsuOZ8M8qB66hmHACszoGWLagX023QyfTocTCp
5pZfCcu8+Pcu4GQeYsNBu+fuNbjVFVwJoT2Bt4PhjR0=
`protect END_PROTECTED
