`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8wgsw6S0bB1bvVCZln0oicS7iCLnhedj1+4gebdVX1pGtIPlCqicOe+sx2bmZ1dw
7Xq4a8jow9+zkSqQfopC8OqY/4IkMrd7HsdqdUyVcYbVqh0cbGk8YhT1wJut00Ti
E0y+feg4PpfKO0RfwAV5bknc7RLVFfkDtafoAt4H1UcDjUv5kNLvn70qq+c0xLof
jTgygD3fr9EJUJchqm7stbVdfW6kLeKFUOmGO75VI5EtVy6v0lnQcg+C0TD/21tH
hLP6lboSMfEZLDTLRR9amy9fAB+JMzruaA3nDhJ7Vf5m0orGSIMRHz4MTRBMWd9y
/OcECAOUztOyaJ+1cXX9G664nptN6y7TxAzMcsNpjkkq2g2FBYl6UXer8uuq+3ir
ADF/pK5HMupqFc4tQROu7qE7BE7DBkNCYUHUeF+XI/7CCk514cALHTi14GMN7XaM
pnPRk14ExeLMxy1UD/XZw16/eZf0AazniQl05XDfnrGfZ1/JUHn33OLl7MCdxLWD
LcIA4RcnairlX+AulwKIf/qFzL+tnKCSu/xY3v68eAQpx56vtOe3llV7ZqdBjhF8
ZNORhXYszf1zgvGbihR1Tar608O5Eqa2LCxQNZcMpwbuaqYA/lhfb0XT+oPFv/HI
OD2jqE3CAQhrtQfxBNne7AXstZWx9mtdpUTEy8wYHKE4ashh2ATrEnGF1xdE9pJ1
KImsdRrArJeDGpeeP8vRHFsul/bFq+G10A6qHLYt/Z9kVaMva9Zr5zuiJqeeCBpN
r9PcDo3q6lD7ucw0X2E/DJrJsXjUpm3Fe+XI8uopThM2dg9vaAg99qlGdrloktwf
gTEqU3Yz/nI/ZekgyN06jA==
`protect END_PROTECTED
