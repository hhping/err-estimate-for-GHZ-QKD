`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4zp4Z4yQkyWyzVJsha4sBCKzw73FeWn7wp4Gvzd8SbFxihv+/sGKAAmT4/7Y3VAz
F45k4Yyjq2naTcMBSngYT63iTIUkNhLyC+/7SaC2yS4WGW/BJloAxyd9ViTWJ3s7
LMEOBysEZbp2at3btCFWDfiseCcKnpgd7vwW9vnNSpeJd5w+PpB7rVAe3BPwGpzz
qhJOtrGUQf2C+oO3KMxqoEC+cnMnlJTCiztDmZLRgI9Rappi59IjkyNyEtezCLqs
H/xpLIs+9zUP5Q0vfiy9ni+yXDBikmmjn/Bvmy/Pp2ILB5ikkVHo6TNnogSHkycD
11hvsfSnFzG2QLw1WGgbUxAhWCWuRuAIxQiSC+cCiZ8+rknR69gnLu9tQqkt94OU
WfOwK3wWlTmJXFVF9gJiRcxefSnmfxX4K73cSYTfKxUoGfqc4TxGCTWngGSQ15Dv
0RA0cUrCn2mKPRbKTWFi6u5sRbrMyrw0GdaXHJWU4pqw+SFtPaAY0LF9YsPWq7+l
nydZLg6N+CeGcIQt8Qpgn7XsaJ/gE06qVfXdvOvI7XK6xCxjppKZyPLMULHB3hj4
XUcup2iZv7j+eOagIfEmryt3fwJQuDazViFrdVz/vA4dkuiLg1ohbHbFiBiMkIJx
RaKgxn2mG8BD5om3NS4ziOyJOUS1qLCNZPiPiyEOiJak5FjsS+/bcZ+uX5wHqP3O
rfVeIjZatxg4qMA2Q06BJDR/1dK1VFSW4YT14T9zgATPlcEuBFpmeA+Z6pUOxuo9
4s2shMsaBId4ogyixgTQQDG0kEl5JINyXsDWZoe8QHaVnIVhk+LPjfi4O5mh0NcV
3oyAGrpQVkGN27NqEicOLHYNPAUHJdV8K+5WUvygBsXGNc6U/VQL8AO/aNEdBIW5
QF8OzCGdHf8U0OqkwLPddV6Yaa4prusskGgTDNTcYpqEI8TWDiPXICY0YRKiMmHF
aK2vrvevN2zNsfPZND3fjn6Rd1o0v44+1IKW99I0TA9lWNRrUcQROCGZwO3gDC/P
3cm72kEcEPbLvYLTNTdnntrjU7+TR4XLr7iW4PAGJ2lje/R+9qFPj7em7vEqbII6
9QpLb2dVhJl3L/hXHP5sIFt8k3b+meFdIx0aqVlpSnEMA2DOMLS7nMm0U0kkvMFZ
4FiOtTIkfkQj/T+PWjHfYGX1a4N6+Ml1nYSZXMEgpsLyCYAvqxHABjX8xWrDXPRk
8mmsB3PU9NFhSNfs695gKgdKZYRG81BTSFvv+ayEbNDjv4KuWTl/OPlXwhhstTA7
Q4QY1KHFhjzfBGG7DRdilCygUQnSqPu+OqW1+kt4PYfs1yamn942gCU+YwbGwwkD
nXJlq2xRMn+QSD5tQ7uf3btyKSW5YyXvJI0AjepXhN5nvO4TL/QD045Dg9L6EkDC
D4sHGoX1zDrKoXMugQNyQWNPyR7AgfGRigtlTTpOH22nLyVpXO6I28+KKUT6XR7W
+g7yyqQ5TTOkiPUtXNok/jrKsD8iPcjVWpUNpiCZgbplG54EqVodt7SfxEUGBIpo
1luFFhyl48B15TzdEAqVXSmsZjskeBIUM9YdR4hSZdqTXZBq9CEq+RkNofevjNbw
2T0l8CnHpILVPs/rlLgHgbZidIA+gc6BZT6vsy1h95tsUf7LsuJRfb/sV6BFTD1m
RB//U0yhIBX46YZO9QdAehuczOkE62Bzqp5T0kcNxGh1POk9tBYylncFFVisxERM
ifDBS7ljYPpzyl1e8OgIEee6l3Ej+Seahpv9g6fTiwFD+11R6hVDLfU4WNixp4G4
pucr4LdRitSEwJCGLUCuZj9TRMm9ldwjUWd0wOyj9by92P/DPHjSPKgtqgi8AOyC
3FQ47PT2kTO0B6U9ih4ioUamiZm42DsBalGMHUi+PFTjaYh3s4GArPNsA5Dp7fiC
j+S5hCtEhdbtwPml6DJHzXjdF6heY6e+kzR9jO0H1WOjdaQsFR/2b7A6opD/YzRg
GFLhttsaLgW4n3vDALS4zk4Qp0PrQE7B7Bs7UMymyS0RshmDI1lwYCqKYX3uaSK4
nj5ZZsEAn+GJhWsV8vecixXzxS4K/GbX5jVwT4xjbu94fw5qmg7Dh6krtqsXHryd
JsX15cgHCRBoKixP19MwZcTHXiZE17ztxEN0MaxjLqpLhntnkLRXOEZ/ruDLzZEo
AcLffHyCyUgdGKPZbUK7ms9ZYYAHyRLEh2Xki6eimv8yOtEEtB/e2T0D4Sd8prf4
bVFikghTSyRcFVPOfEsIfkdC8OK7yx7wjHPs2s36dusrJHi/9cVwAb/0BYCjFz1u
x5OgVpraXmAqZ18HKw/+/Ea3cXHyC7/5nYZ/5qGnQzIgVrA92zBeFyUN3RViG3QT
HARfUSeK1yGFaIjFFrXyPrnwWGj7mPk+BSDikqN5z29fLTWxy7WTkA6ww9wMuykP
RXak2MeZjFXrySDfzyhq5h1qdrMI9a1CXeQTkJ8xf/5/rx6VByWkXFN4Ts6J+T6s
LUSKU7pWDJnYym013iyuv9QtoqjfBd3txx0pP7KllXKpTYcyQBiwCAgFTw3mhlhk
xRXMrG/YNzt8mfEQtSGYdYwqsY+Y9dgiNrAC9RKFNbrvRjZcNKILNN1oRMEjHhhk
ifkg49Ju36O6++i3skUSg/F0c3yv2pJv54tUlPznsc2srqSLR1HkqYGxuhgOQTfr
WFJFDrzhHCJ5mSCvvQvVVrmbsdTMP+OL4xNrKIsM8jh1zGZc5U2If144Z47Rpsi/
5IlAHCV0yg9nr/j+8SJ9ld9SBx3KRK4zzorRnST76ei2OMXKE6Nkj0WkWH8FtOmi
oT347EVhJb56mK1c26CrRzonJvPmOWURBWOVKR1fFD6Hdp8dsUcvdneMMDlIM9XF
JlmlOKBjRnJUmYkCBs7NnKazF4jxfx++HA/K0MUL1pXorTd+k3xwUzz9A/OZbOa0
V6AW9aepewSmUTvUTKJjJuijNh98jQJtr3rdzHBWTowtAawtDVd+1YbTT+uCj+/t
+mCkVQxyKRgSgdGyz3xEBJwZOFsZmzyJV/yCqsRDKIWPDFiqMrmRHzU1J6b2hQGz
vE5OSvktkosabZPqrSPdy/1vuH2d1gGWVPu1T/mTgWOj008TqUMyaucI5Yxx1tWD
Dg1srX/zwS9RYoE7E8tLRdY23W6L0tchtZ6PRDiuMG0YLetJ55qprDVUpAfEkixq
WvxxRcx2sS1v4Voqe7WAo1nt6QION/kDVl4QdTUaYKRhXMyTeSlyzwfKHlNQeTrN
JzRlhqTP9tP5K2LJE3BYrGRa+sKuluIf4ZO55JJ8mPt+dX66PErhpj4GFQjPMPrX
1K0t5pKX88sd+3Mvi9rmDgrpiP+Bb/i9+W/6Bt9Qi2zJrDQXJhTGar2q/slT60X0
L7honp6XcLJQbOY7Nrkd9EX0YQxvLcR0qmKLutAN9SO/mATZBdu02qD9RhAu6LL5
yi1hgt0LkggwXcOTldxcR+/be7dYy3xFrC4lu4uA44XJn61gzslUhFbZQgrGNMgY
A5x7TCpWoPthIfqItQPTSxqwsrhNj7c/MHR/usL6pT6C8Sed7eVGqBN/envMIlAn
zRG/rX1RG81lpS4AfChfiUhKdw0dFNMO/vFXEqgMEu82CIHpObbrB0erlSzCNKea
BexC7Ic6loFhXsRINrcAkCKTGhNaa9jth51o6evVPgGMb0mDEdZzhQPIbDOhkqHl
ko0C/Zma3x0BgyPMuVJIDXk55ZBmuxuiEtdyleD3JKKBOnLj5Nn46vIhjUZgnsXB
iDoqPbIt2fnnYphZuboisrpnry6ugbPcyXVOFXRj+fN1VARuWA/dBUjcNKnI/3og
aXdxXhWxcu2bCE8lBWdppHcmip9FK1t4qyg1K0IQBzAZiNbxGnwM8o5wFIIxUf9z
CicTOhLJxLIBqM78oaAWpyLVKwBQ1gNqNR3k330bFABbk+RMu+ywZZgJMmOD2owS
2wCCl4zJz2Lyo5I6hf9LAKdh2wR0JNZn2WrLpc/LeNV4bZzYtpG6Kl8YtFgpS8FF
aniFZLGxbme/w+Q/sAmRCOfCAFvz1mWA+Z2lCDuUCurG9PR9EyluR8akyKmqJv0Q
wO8+zNTvqBn0IYQXXNtsdsqXtEfU8aftHmP6nqPxv07SKNnvCftwvpF6hJoIv5Fs
HJYDM/PnawD5Ts0YcxGqT+OlhCNy7rWHwWsDWnAV/ve4u9/tyyYzp9KYOFvezVMy
L8XnRds5XwPJz8Enyz2wD+CUfl3mcAT/buZ/jLulYwYOcMp0nL7JIsnkcBPZNWI3
5iWcKuMc++kVYywMbnOTB2SHlLxr3F+WJp3YgVfZ6TayXeRchh9+HHNdW6yLfiyY
VzxIOye0z+mWFfPfGCoLN+sGJl9352jZLm9QjsQvzg/4VymVQ03WiDMGdB4eLLfT
KCjg+SY7Riw9sUxLzJsvaepVGnXg6LBXyruNXgbKiw1mpESpjAlBkEN2JJz04717
U++xQ5tlRJsSmDi//4PpBCiT31t/zdRCopeWrUICwLO6cPYiKU5Ur8RiUXRCK+3q
zX04hYCqe/DNmjvU5KzRxqAOEqPPhuQ/xbJwgFoQnyO8z08QK2b/8rZnZ18okhBm
Q/W4N5ADf6QYcrGTXdAGgfl4RODSW1QCnkevc0+9e/yiCjH7mrypW+P1cpZp3ngY
eQVTNosogQEVX/tCFAT8ykzvF5qkWb/QudNAxf1BuGmVIdrU8Iq86V2Bd6Kx/4l2
cTBmtJZTqeNB5aUyKgh6zZTj9H+ZXpA7wQQcaC5WLhvcKcQdkvgmLw89YHMze7i3
Os7zcBZWqFblK8TCUIdfE6U2qgQnZsrMmDK96l8xqwOBxGGPktVfectoh8H0kn7f
F3Z8LcqcblzmxbH2I0Ejw+2yuYF7YJ8uBf9HA8md6Aj4HphJj6sCemt70wvFO2RU
c7YlKXCByHTXI9D/p9UeGuKizAj6g2QHLOZo3rLpecItX+czrEsQDwngBy1HeT0y
OSKOAbyMYtRCP20WIV3Psjz1CAlN5xK7fVz2gkRDnxf+MkilXhklsChQJd8TRt9J
5pyzY8rSvjayroGCTCjF9VPh5D/9IxOVKzP3O4RdUqoWx35f57iU6P+JF6d5VMTz
w9C/zyUlcucOz70FXlJCNvcKXi60kun7B0nzD/CT4RrjNEwtLRbO9chii10yNwWz
g+y+0KtTtHQIFjSLpshwflIejZ8Sb4gD3ePS/XdK0OskVFhlKWXVfKsslh/MiBqq
T1Aw4qIsOMZydbCXiTVRkUiqpSrnp8Cyn2pzfMBfnojq5uc3rrMMQv/UtIVHcVv+
0CTOXvtTz9BFlJbGncaMzl/+37s/iu8nDTfcmRelgE4JUWOi6lwBG/o8yJ0NdSGX
wd+xMYlNOQ6matnkwjCHlrrWMOEM65WcLsbLWWIdVRZEFsr9iFiWJogBaHMs/KOb
t5wolX/damhuvTzQwc3ElBeGYiWA2EQnGyNlx7HYE5cUCJzA3ft2+Trpt5cuDr+s
c2pY86K71dT6AoQWE13r+GIXPgmpLxUnNN9/yxDOWKhpJWm0fslpUvhBS7/wE60Q
pDn4jREfBV8pUj4T5o67NXT940yVUVv06hGhjwu0Gve+96tSthIu0jnCF52nTAGK
BcF6ut+1kJUj3pbk/oDVRztGHAITFmJi/UArbHX1fivZynEJ2+BtvagibNsHgYhy
S9F77pZRS5297qGYQrKKYx9uT8lFstmTNOAazGOHSZWuoHs9XxOG9di9BcPHlT11
YcUmDL4uD4CkFCOP453MR7fNtvJFe06xDPHgK3Wm8bgA839hJ6dK2TQuS8IpkcXJ
3uKugtrnUOfx42O0JRrwYUpS7tclJYgJuUkh+1nFE0CJJfJNTpmAXCfPegVKMdl9
ldZwJ0mmpdZdvbMa9TOx84lznx5KYxk3a9cDLx+9h0DfGTVXnBUGx22z7Kgw3sIE
DaQkt5O0Fn4rFeo43pHLhoYDZjW/yAPv+O0xReZGn+Nm+zJXYbjlRR6GBHcNO17P
0Hm/pHVXDzSzHw0Vgcqg8uryjLnscE2coMy8/mOZeQn3UJhfA5vAlor6W/8DxVrQ
ABwJN+DA2FKGGdho0c2Jlv32loYUFqHQew0Mefc8qDR97pA/Fr8iDdCzvK0EsViG
fCuYrXksYUl8AKz+nbuSJSw6GIArAzXUWaDAYvzUVoqjNLU8XIy5VKUO0E9KvyIH
9gHNPrt4So8y7bSstiqfmB23PFB4vr6k4TU8gMOgorh1u2gJT6A32/oVGQ9oqqUn
B/4TSALX2NpE82HoclD4E9nwP/dhDEy0dhSY8ylE9YCkLR5u9oAtdxPTV0OPIsSe
MQccZKm+aS0COmJR3AQP0Fj1TnTedR+ORfHGWjJP/BV7o44L5ArwFcDcEhiJlbg+
gZmx5cw0oBQBzxuEBGI2rQLSy5372VvpCxnR67drNv+kSuYdKdhswR81okJVS00e
vwHQ6dEg/pd0nGSZzNaD+0jVu/MoMQ+s8tueDqTtwLyXKaCcpuk/ppQPAxKP0q/O
QgGCx6eGJsAfFAjg/jGvzh2DmXLzAJrhEeDJSuuLPQm7yXClLYwu9A+ISM9UyS6J
mb6Oze43UUR8PnWdZJyOQS0Vjr7IbbFV8bDm69tEJoZLl6VBf8xU9nZM211IzGcV
JahNck+zSahYajCANKJYcrpf/IxRYzEyWbqhkkTFGS/BOezWE2iSdwWCohJsR0XE
4hv78lv/QWeKYd/OUjHexVX5121WhG6NwVocgQFsoW+EeVUYXhCjtolyxCrwzQhr
M0g1VbJ3ih5Bw/VF/IhN2V9FLLadVDAX7EtbUvRc/SGfoGfq+3BmSWV+ZFSVGegr
mFL7Dm9ev3gqAJOXvoVRcKlrGQKpZbaVVbeLalqbPy/44v8HvZhbd9PQ/vR2EL52
PDf68IF+zid7mzZR0cAQsjJUfuHPzrr4tIdZ14VNhJxnSxQvJN5GIV0VyrjET0P6
ZeQpsa6OgfkGmYLJxq3Hrj4Srb62wCfp40s69ttZoOWNGqfplCkysRlQxSQ4kBXq
43fVuKPC9pknPPCJf7Dx5cYpDdPiEY4UVTa0D/W17OuXHNv1GI5+LilsfyuwX9r1
/j259hfNKunVlHEoxmHIVgGwsLfb72NDIORMVfQgIMxFA9RWLS4Jlyw8wEXB2vaE
PuewWLRGmgIZWN5n3ydKxYPcFSJLC80RevNdiB64jgtfwPrQ4RvNolstq0ILKkOE
V9AsoCKxJJxflN03N+bUOifx5GIzGFA041oWrdX9VQttIOhlzh2y+Hkh22ZC/Tws
mEI9RP5unirJP6EGb0sCpQL3PnUstA8KigKcPrPUD62F7DMaP7Zoel9qT9i32aQa
NlnzOujoEbcty5s/i/k0usISvZpSAMFu/DRidyt4Go6PgDD7lfR5hWD//nPYplLq
Y5nmjt1ITHenfDJxHChKJp2Swva/6nk3aszGAmbkYG/Bbh+9KConKX9JxAdgWjiW
AXr19HkLWk5my0h+TrRS8enHvTXLKX46OI7FBiAMFT7+qXaam9QxjT4eeW+tOh28
/mKWKHiYAIsM0F9idgZKCzlyD1IiCDsGOMUVbj1XuHr1A9NskvlfpWSLuzgJFEM8
0YOlOdptjnGEdu7F5Hr6s/cAtIgrMdq1ww3JlmYuwmEWtshL+ZOci0tgDQvEA6Di
IGuaITORbwXJytg7fiRvP8d9jnq76CJvyEjQBHlNC9AWCMQAeb5gx4pBDQBrwLti
pJ7lRaWtbanxvAhT+bfBbiv5/JRJsUH9nSbi78zcCiUpFC+OTeovHJ71j/psyW5g
697nmQOlmeDTTbqg5nN1NSXSGhJaeohFIfUbzUmQ99+S1pmUwi8f2LhIY1kdAWsf
OlHSimPnsWlEECwOz8nkuxsIqbstlp7gx7xakhoavWScu5CI/kHc7PuY7vWk2tJr
Ut8uzhXm+shCYjIO/A7VlMvlC4y8/Scr5wD3wiVd4pP9+aHSYMwEIQoefKttYHGX
f//En+cGdrjnQaLyRC1B0MBCsItfbh9y47/51f9fIJq2Pb04W3hBgY5V8LcoscuZ
xXWMi+fa/Sw0cSGriZ+wKlUTboxPU1VXTqlxV4Jgrwo2wnWHfZkNrMWl90dj96p2
3e+1WXYJbrW8xiHfjamhptUuLkJBaavf7gSzTjZtIWM1vYloJt2g/L9SCEPZHw06
rqDCZJWaymHx0BFAl12qWMz6ZTzzjkwN8au2ThW4IW5hARZElyxTAckLxn4jDFVM
Mw3CfeYfvXT6eXOYkhNY8iloxOklK8Gi+O+NDcrUXgDdsbejLtvx/HO3Kla0Ikgz
OS6dL+F272s9U4T+DhQcbf+vLD7Yofb3a+iSZFmGm2En5xdkqVYZA9gvdgLF+Vqb
iix/r8krJmFf+VPnpcw4K6FQuzkOKhq9Vz2q+xykYYPhXWaKgT19+EPIxyEdzZVu
bWvKLGKvlWeMs1UVqbtRYGmrHrOfV8gTlg2C8ka+3W7JzBU+Ldm66lVnpuFqqttU
ArPfzNjAlAwSojeDwVuV5zk/O7NYzFXtibIiLyE92vw43I86aiteLiZoq0t/v2jW
+wshy77V8cHY47Df/BSSveXshSY7eLuX2xA9psREcOwzqL9QaQZSoB7WYVkhwFhv
nrg0XTShcLI0af1kKSu1FyR9eRDcFq4z1evAufULY+Y80GPibaqmixrz4foRCjKy
w+l6yjyAGAEEEDOXI3DNqI6vlDaTEcbv7CY0yymDqWdF+nAFi90rYR6lX8VBpoNd
WfA7LEWoAKAMzAmNSwo8yrTpeg6qMBK5/GkiqFOPuPXlZpZp2I4wJs/T2jzfdODZ
BDyeisBhkNIOyP0TyEpYGw4BCQThbWQ41b076MAcNyDmPlan/F3gUb9smJwIxpdj
MjQAlBBhGhV/C7Dx7v7aKMwGyFeRiqsYDoCMUARs+G1PM5xlsgzMS6nQ1wTIJHEl
NqluRrxu6dWishOayOb81OFVY+6hrUXNyEHXD7LLQ8o9qudIs6rLJJmUNIViNoG0
UWy2bes8Z+nX4s8ZoFgUuwkIdwl8GOZsHfz7ye1r89gNsi6j0eshldFmIboDyhLb
O9fVqSQaT8DgRhU3+qISqvet6Hh4wSOfvUwayvmfkPhoeubGBZ9cD1LJ/T/wtXSb
yu0LbdeRJr+wQYfQUxif+fvtiJwN5BsJXHb2Ia0RLXa4FEp28bqfLixlQLLyGDRm
I0ITzLcib9WiCZJqbiMTZwXo/DZ1nydyLN/h9Yvw0EF/ds4mCfDE8Uj43u/402zi
IFtzZJibVBNCJhN+8pIvStSmDfBTSgGSkNrKLSYwgTSu2OQxAIQu47LUWIBAntIh
D+V+/h/R97aDa8dmf64WB184ij2PAGCC5B0IA89agn0tyhYKJAVIEEmkQs8GGhcs
3kH3TFM+v7DOSHS+SWlDwSsYb18FSdRqznmcWVAvV94RX4Ob1UkduJqZjPEhVScv
stgG0axe5AwVAKeomb2Lfz+J4o1WQEhseuOd5q1RBQ6caXdCStls1FiP4y6QDi3P
R4YPr91x2G7WdU5HjrxifRfymc2mtQgOWSszxP4Tri7KWABEDmCETilzce28aMUh
Idx2nrwe2/nAs85L+ePITIiWcmrJmcIvMf941f3H1WQNTH+lJamwShXG7/S72NjZ
hhD1DkzGd3Tvh6DR/9B5qWgCWGS6vxFkpX+R9Q+mDC2+iwEtJJ82Mnc6WHez91T1
p46cvhhujZoh1ZiX6KTM7co5AYPtjM9/MU+WX+OZ+t08xYlORNYdAIfy5EGE6m1d
eA0t404CKWz7pXXlXfjkBpi9OHDcwuUBNPNVWMz2Yp/6D+2TlsreITVXK8mZj/aR
DDzFs6St4hYOvmDr1ABTmb6vDNcakF0H/uUN7CiSELzK60UVLmAKzIryi1GCf7Z4
RFofxIOXBpw7cskX6LVycRPkhYMBtQuLYQLQ34YAjSD2LlgmPtWWy+Wr7dBaZtO6
PJiRnuLJrA5JcWcdw3Lv6fUNR9VTUWQ8SEx/zwKFsbM20qtSYiqo/z4denPS8cB8
q4qmB+uRPP7rDRjAp6svq6lOCZCL8mlGgHScpCI9ZIfxX2GzfPgxymbY78Kz6/yF
1UhOVZV+xsuB74VVq5RtdcGTnI4iKwJzfNiU/8wmu1I23HAnEGdRqYseXNw5aQ+P
FA/W+cCubhZe3XWZHCzatpOCLMmiLhjdtBXF9UDB8KYN5sTtQOJM6MW7I7cKc8HI
B2dPj/HgeXNG9f6yFl1/0qxr0Fcx86YIzzHbJyv4wCrTsgG+E7B1k2lU5R52pJ0U
RtE7EXAlpF9aH/MVbRwAay4qkot3Lh20gTz3SDyenZpErlQnAmfXrkz8NRFqrVk8
X0oV0iL4Ux4po3PxLHflkZpjDy2zmN2RoKRXqJtM9bxQn2o/Tx7MLAecH6Hj6LLZ
k7NmEHPTMb4mzQX9oRU4y62HF8UVJrEVXt56ZoluOFpEbeH1lXXzXld7kOix8AMa
R7VgBv4MUlFX6K718uSxDDLHUq22BuUelbU6FrAblVabBDdTkg8xLFtxL8B9Z7yN
79QsuF+MMbBGMk8TH0QRC+fjZ9I55iaTkS3T1K/8UR2goQcRYlHhlNyUzhSLgTd+
fhXse7BvKJyYjiHmZw/WW8pcdFox23CKm98A5UHK8reM4tTMi/eohKfW6+U0OHjx
O522BEnCDi6oQFKOpjNFcNlALhLktlqkg0qQezGiPy0owIku5SBBXiTXiSG6G2lX
K2yJoPyjyLcYrGWiyV3hnCouvdvaUufDCrWyt1Ut0GHh/bnejzaNtzRB3UHoWZPV
MfIaSdf49/YaPfBCpresbQxByDYWjrZ+Z8EMrW5B9fvZ6FZyyOaVYOsAG+Wiygk3
5CO6wKGSPvqmnNZO3Fn1NDtD8UNMCJ2Fmpx4y7rGI8JNSa3o0yel9B1aSaUxU2Dz
ZB9mLj+GLYOlSe0C/Y8jTxUxwyqTHi2N7d0Oeb9s89dOFN3a/fquiN1yeUso5960
8K+DaBAN93hUMJk0puUooBI3yJyv9wAbM+a0LhfjR580m8gmoLWHXyDoVgxDt7Me
K0e9soyipajTol44eiQML4dUL1DHKzaL7LHRpEudBzPbNvIbPFFiBTeqI2223mv0
qbvX3bXlnazsUDvN5As61AAfo1DBOWXeiTqHkKjb8bVdKdGDBI9gyzI1pAglYt8E
2msIw9canqhjqCAIhazBrywxl3CV8TnOqQLXygEep4M/V4KjtLmEjl+tcTe9+UW6
i+cjXBGrvhFnLxLQKfNxDWQwygL8Vo7V0mIUcZopTMmIfLlQgKGyV9n9eGAWki70
0eCfy+5xmG9W15rAcnaUEXHtp+yZxgrc2Be7sNpyVyL3uHwTNMVGrmS91nCeSnkv
4N6ddR+3eJ4CyN2RP4tITxiWkgWeHluBUGW/pDx7aeIo3k5j0w1snfB8jB+Fp+an
LPQ7pqMRPkZ8NHRurbZgWy93VsuQ/TVHsAnkeh0MZ0vuIiGPvmE6IP6KHQDcYX0o
mzqX8I+9GUW9DSNl4NDO81M2Wr/C3Ggq63y+0jGMb2QIK5ep0vvLswGiTtmRT/DZ
QQT3SzDtdHXmeQnao+hiUx7SmudqPTvG0JCeVxBe/oqt4p8sMwrk0GUxYdq/1MzH
2lqUzeBX34MLad116zWrmS0lmDlP05z6MEW8dIzdm4F8Sg8AII9N4f9E1oGisE4e
+obqJe+VSAAil0aazJ/u+mo/BYR0/m/58JqZkQychsBjksAFF0o4bEFY7zVeqFaM
rD9uKskjNyZtQVfmdPZupIPEx/NrGYnnK7QW9spxf2OTmM2/H0l43tKzv2mXy9YM
SELLfeV3Nealki7gvIASbv52Q4GYEB4NMSdQfF2gpE8mlsY29U92xWlqCIlEAkvH
tAaCHsU3eEBckFnnrXo9XgsfEZ+NVwHqQt9WT/Wcwv11VJN4BFod87qdDhyXCgEQ
oczOjcp16agX9G+jGfRzt7Fy+QMJ7c0ATSOqpQ3DCP5QSRh39IuoxKq5txH8Pn/D
LqJmpsivmWKOaGSP0MccIt2/gpritv+TZ+w0qYQqLpe83uZ5li0yaKloaquiEUfw
i9tfxPdPgVBppWNsOev3tHTGZE1m8O4JFWIZK96b9Xoe8r5tJcEpf/uKVmtF6Hcy
L/YLxP3TI+UyJl0LVqFJJtWZj6w4TvQ1frrt2m0y1bADebMDB/Q8hcBm7VqHOYIM
08ijuAfn81+x2MYmra48fHDFL7gs2d+H4xMMQxcu79pL7A9VPamqo6ZuyAmYWa9s
Mzg1lXPEbhZyRj+4kQ4n2uciIUOK9nf6hGjrNTrWj+P2tV44DBu11TJYs2MXUsUw
CZJAeZ6zucd7FGQKDWFcBjUOlgrYfd6GeOimj9OioUMDs2B5J3iIcw6qGoMmDP/p
KqRoBdunDwjowUs7GfvLMxLoqQrY1fVyhj4NMFUnTTsRT0ozz5286kaj8lMnE177
MXh6qCtlwvD3Zcz1Vvna6Qrexh0Hp/8Aj83jExhsQ0HjE0IccVgmK6AFdzlPGOzX
6AIInzUvJHcjw66s/wx0RRVqB7wEHXeYtgH38MFyxh/0YFYFO2UKSC4r7V2Z+x9t
GtUWfJSbSVlquru1jGy+KhPYbW6PJ0z22+NswNb9HtbO2Ezwv2F0VpK8DgNBfMXG
BIuIqr8aS4iSY+8NrXT6BuAsbSNaLxjsNWwkaMv6WIIUGngtG08hiEuMfWPZ+nBS
egK+msp485S6k8jJPR5ryezqE6bzNa/tdFFGe8fpIQ00FzQCw7wt+OyZp1lrK0od
glkSKJAXMlbRTunKDcNaYQOtA4b0/26gAu2GltRCWVUfJWw8EqZjE4sP+Z0GRznq
99rtWCTGd8EEpOlZiN0AXeykDm3bdaENCApRhnhn5XnLzr8gSg3nsjcpu/Duo8aO
yltKxcY6diJ9aBpGZYJPIAn4Q1AriKs34qEs62W18A8Yo22aZDUCUaz6dpkbtwPN
0+aw71X5fd8OCFTdkztQpgLPnUwvdg8R+TgKRRU2R22Gg6CoSXNsdW5lbrvaznxz
8fGU0rPE+ZymjWRV18GDXX4JXukE4Nonpqj4ifZZ25IGlPTrFy4DHPIOBaM/uW4W
bEinrSlNaP/5mVruQWYX+LFFaYdwZBLI1pGqueE/ewv/7lm7oEWck58lxkan2C8b
7I2KbhY/ZTELd/sBPt0eeUbpKO1WHuKZaQT2EfQTg93dZiKg8rauRkCBYwtVlGhO
qBYMINj1nzJ8lF5jl1vQuVjbH47fRfpn4YCMBYceVUWgXq6bmMK65X1HigSn5mKh
gvm1RweTDtARaQYyFdjGOQln3o6GHJmjjPMFEVLV8g9cWdSwQYve5t0ce2293TCA
YN5oxzXW8KahRmsjitgJluVbTj6Sy8tzYpKcW2k6iuzhHmjnNkNsn6S88MsNK84d
8IuGQEAp4bzPRuew0XMlTFkcUn1Ynr91uCIppwG5ZH5i23dMt0SmeQBtVo9ZzArW
FfvA7XVcbMH6Fz/hQyqj3LJoRO2J/DnvbhIXEnqxQaEBmFD5NWPJi85/3kW/J2iK
Ky61WF7DMLp/dfh6vuIf1aFsBY4wutuJy6JZ5T08/wjMfwCbjWe3nW2a07JVGxKb
dphqY4/GNLcnbEl8v+nhgUFJE104KRHHu0xHxgzvsfJajNxM5Wmlinr6t8RVEwBD
56P0pgDRaYQrk3PCOVPv9G2ekPZ4h7LxIS6UaY2QCLvVjZ9NQa/nKO+WEt1VOL89
+J6eZwALzTJAWSoJu2fhRX3TzExugT89fz32RPEbU5quZZX2C/OuOXO3w7J5EZ06
lX6YybLdpSu1etdBEz9dBD+LM+fLRoxB8cSFc2zw+nsA2W3FHYBSLNxMYnRdAwzr
bI59FOFqncQHVh7Dbq7wkRIY3fwFgCB42yPQwpNqUUxWGjxN4QCzMClnXH3GLFDJ
lU7QbtbuRAIYyFV/BBORc0XxGWnsnJq2+oxY/TwuB60+deobz1H5WBOoEJ94l+Vk
KZbBOL5IwXti+ur2Yj9ENPS1kqULqtWqzeTyvCk7A5cYn4HZW9N3mPCEkBt5jcmz
/sqXNPLS59mBeGIsEFNKa/dtD4DVT2UczhUy43a6kiONzKOGiyFGB19b2lOO/A6D
G8gA4UJrRzq17eULt4pZqr569P7dEloQzy+9k6APQI8095fm77D2pvKuScnCoXU4
05fK+nv2dKxQ20oh7T+GUgsvViMUvjZBpYRs0XqVbjGLq7+pEMJheXfTCaw7XJZW
HSxcGvX6uJMKHDAwJkmGBV5+HSDZpscUSrZ06wiJJjmow96clUoyvdyaQvGsdJlC
AbxOHr0nhCan16QsG6Iw84hFRY2n0DwBjuVg6KCF+fGkwco7Swu6VvbNc2XHyt1Y
kRJ7vU5ZqlLarIbfeLXODavhboHAn7H6NODuVt2HWZPi03ACNiizddmN0WNCstRI
R4L8IAeh42JVZmhuy+gm7ZJVoVhbpQ739HcmMrzu5xra9NNIfszTAvG4sgdof5zU
iUphu3UJhsi9jcebR3FV9vx3eJo6DdW2feRCiaOKrzHSlvzCNCVcOOPhcqGcyhPl
9sLbWV+jzZzwR9zuK+nE6YQOnAl8uexhisvwzOnBUC7aPfmezkL8Sqv0WrnY52ns
KoFQOnEgDbs8tjKmh9exP4SCJj8ZiNPHJakBELZil9lpg6dTSVRcUIoNW3chw9OJ
7dVGxMwHwfGjmMZIEaf3cNSamtrCM1NNJj+hhT8BsCaCH5YlzM2nRrChnSv9p534
nyTrLJOP4M0Hgvw4RamwLJ5uBZubUnNzaNzPaRnyy83ZVkeyFMqW40q4GhSkZJeB
7Y2pUKzsckHLINIX+OZYaPW/+AI/wvRuXxnqGhz3qjXmAe0GZajr1M75qRzoCIwh
HMI4ahroFdrhibCgeY1w9C7SSz0ET+5sGspaL12tasHX6qO307/cUmVbQvJ6HnZX
Xn1Kgcd9o/Yn/engS7eCnPypGaXa9BQ2JRrHKht+QJlmApRsw0iu26nqxQNYg6Sn
/ZtW7/hjMdrzuQYted6QUBjHSE4oqg/EpdfzrVaHrkbbIuCqMEhAbqXO3bvZYkJY
MsIAANnrxpU2pulM4y2prpFxE3+H3wfudsZXoECmr7b3k+SY96YckSfEA+PS1srO
j1icOISmWUKg+k4UYXgJeD5AknnJRLPkmbdQMqc14L2UjEI/cjDfICGfEfIrzaj5
e5ilI4rVcf5kr/PFo0BZ+ReZywRHxbQ9D0wME4iWaw0/AubkqxUAk8qblDaqcO1l
5FeayIZWQPkPyXEhy5wq9PCjIOO0N0guwWBYimJ/jlg+7ZNQg/VxIXAi9jo5AFF6
E/eDMhxm6cWFuCAaWQF4xxdv7J+IkgxplYvWY58HkIbMlSD5TtRosEUhZzMhqFpU
WAkSncPmXzRj6Ddz8+h6YwvrM3z0Hsk0Dqx20wfotYQ+l0VjXBFeW64g8OYSrnCO
bbF3mV4PPsof3k9o9ZBjvgb1DjTb3bTWyq3WZmAPn06P/1FMYzecC1LcxSBpuj3M
63C+pGUWrqyxkHT11j9N/bWJVaEqxSPXtkBa0HBgxDtjWUVxT12Z2z4aSQJ+WMuu
GIGAAco4fI3A44u3ZfqIH0pSihstADfLEO2mvZVPJnbhiKZuYsRfUoIBs/KmkIzA
H18kusZ9LfYEQeRZjp32EI1enKBP/pxB4ZMkXEFILEWMWfBG4nb48BIxq8cZ9DZi
U+X8snWR07EQ1S7Azr0kuSoYBI+ksJXDjJRR2oQLKQCQDezxDJtmKkYq6PtMd2Bd
zj3beQMeHVvHNUNkW8Bfo4voho7Q+V8SWaAmkBko0tVLtGcxYqEuRcCM9maHunOt
GOVB679zJ8rRRBPCuAW2vXciUjIO3P6IOVv+SRKzfF/8ayKmqaWPHw8VVo6713kx
VTb3xP9nfcXZVC4kuBMK+AZH2cWmLuhRVxRNdUUceR6RQKLQl+TxznACilTzHffv
dpFIzlJ7hYoJQ2fbcv/LBDttzFlYcTkZhVl0Fn8BdEguihP4NKeH4eCAx0YDUwZl
jxEeFqBgKzOyLh5l802TPlQu/WGmrAckt4gjHY2Rxa+zFBQVZ1BBhkWjAhuCPt+7
o6q3wp8rjPU44cx9/AfOWb2Fog2p95U8vX6E+9p0qrcIv4tTIeEJobWRWdNtRtLR
RgHDjpgaj1tHPhph1CnWhY432Niyjg/gy/T7YeBjfCnNttKx4fKyMR98ldNPivNb
X+dWBTIr24Qcc0BBaZDBYL7+atyhsxaPaAx/hp+bHPOA04wF25YCYHPe49/u2MZj
gDRYuBXmNn4VGWib3KMM0WarXeE2Bp37fNSy7QcHo4F2EHIS1rvvUHlQlHX3/6k3
sPe5B5lXfWVer4nw2E8HvKf3/wA9wzs7Qk2IzR4HZdjWzfPOaHQC4I/RzqIIlDG/
3YF8SZO13K2aelOBHGFozgtuAPwezwa3UPVqXtl4/LlMg3yz7+txE94GUdtsKapv
lnimO81uhzt4wJ4V9gQaLLUpUqQKaYdcvOYXgqNqjhluqYqxcHtsZHjPpmS1ODM5
PONPV3xYD3TXug6U01mf8Fk2fSD/edix//NwHk5itL3MYeIC5/w3X9q+dTMkqeTS
+GpNXYKYdR0su0QHZpldYEVKW6uNNpPLqzfI96gH1cEWMyMDXOVQFPrUj4lkOs4c
OL/gUUee+judEHIaicuxEXzxpLyg1eI46+ylS6Y8j2vg2oknuxaQ7ioLaoKc+dWB
n/bFUNqSb9gUEO15ZK08qRJaKgqVsqwG5HFojzGlIVn2hP9/bcrGoZ20j1dmxLhQ
zE2NU5iftsNmGHdLhlUNxzw06PymbpRG8spWC3vNhqC8WWqpE8ktCfNWL9ensTyt
Saa8+yXpGBP1eQSqwTNZ3i1qILrplw/3gAuZGF7U0O/n0ypxOpdG2C+k3VijBaMJ
R5rF/mh1v3NvTpM229pleKf0oqLR2uTp35W7KwzO8mmp1SbFE5OzGxKy8AuUmJfC
J2cjIEDle45CBCmlVjfuoeMWodYoxysFmScSaSgY8O8ZADm7LyTPyEeuiSrvpxLr
ohidl4MgHHRt0CaPm9zP9ryiBYcCsvw+7Ax96riqnsN3EJyVW7OiqxYWga53e4Pm
AJy2OQGvGhF6yXple8Yfwv6dkuFGVL6IIP16Uvfuk/8wsqaY0RJVgurJGdeF8w6i
vM1GXTmjoMqcynqemK66DtiMnVl2m2dGbL9F2hgjthBvXoVMn8TIieFMCB6y9lYD
tO/lYu53qktB82CO3SV8Mw0ig92zylCTwZLrG/tL0kRUJq2zYA8ESoOrynzLPe41
Cd5Jo5wxYA9C5EHF7pRjS/V4poxcLm4GOsX5x4FtIMRgXZIOq+IZKr3KWH2M5UWq
+1cKu09gNnL44Xp5dVbjyLcd8rHaUk3mAuZ9npAeDLBX7/DiRy9AvwKGgR2fogZi
T/VfqOOv28UPpxfHFJB3lddfhFpSs01jlttzR7XKRpvogTX25c3c5fkIlFBLyzJF
AJgG/PFLnEU0i6m4D8UrY/YLnimRzQP2DaRdPzBYkGhdp+46mPbH2g6GiXwtw6Hb
Vbg29ERC3PPS/1LFJ0uKLKqfsWoNa5YI/JwQc/6xhkEdOFo4R++Uqqvg5mK2Ll++
Ix+KtLt3zvp4+QXf/BT7yQ+Pw4l+qoP+W1gTGTldypY439H+c+SiTNbV65+sZdAz
wZAmHut8AeLV9GtxP7EVdLpu2jo4QdVmbFZDiUscqwPKdzFxOoa/QZdzVxe+4gDA
AcXMqB+vbOGQGMWzsod0wNFcy1c6qAnbv3ZKC5o5PGDv1Y54jlChkN/bQt1FR41h
vIFYBB7CB1RvFF+fqDicaMaShPKWKehuKGv5lgmNlzvbWFlwhgeVAbyn7xF5wWaw
p9/YHsrK2XWpw/N/Ah4zyLPz3cJYxefYUUswDb3FcS4+eiHg88KpU1VfJV6UWBvc
CpKo4atBXMcpuKJQeJmgKr8yE/fdzQohZuNlGH69KHwTWEVQgN0wbYm2XeRg7V7F
sQhnfSs4gP7hxQ4lim9shbFbeP6sR7wp40o2vlyPOHuJgCt2RCg456u5oouUyvcs
lmRNQNnZdXqzMbH1QepyvI/kIxMw3X/nbkfsMVeoGDzQHmhq2uiBXjQUeIeW/Zte
1QgCjcbJUBa8s85ebymxvhAHml+U8cEfzqYn8GDGidZgnxOKG5lKFdPIM2FYnepb
fdzRVFms70T8+erVTs/nfxces1Q4MQY2i0aEPKMuYGN5GL31HEXYGYX/QbLAuGF/
vRHIT9KPvchtvLmwYwMBoWyl6UJkqtElnFwF6eHno+iM466REohacuvauNaw3OoT
hVGrr5hu56vednTMelYu95usMSjqgmN0MguBG8NnzlKyKoS8WJ/Or+yBq+Vtnwlj
+lc7vvSxkDxrO/YU4FpIsXBab1uawAnaV4I6KsfGz8L5aBb3ccOFuOnJFSepEQDr
3PcPWRWEjepBphcuKqt05F341NjvfGpaUE7wlC2LXXAuu5tL845SkocsD9HLM0ck
xK6vKJsQCW8WIH2kAHzNGpt8AUysWXPPPOU6vIDDTcXNgGGtnr3AFdqXjjSdhIXa
7OUAyuQ6Obhsni/OiqYoE//3ep9E0uNf1x3c5C2QVQEVViRQVIhT9iwKmrdKFBrh
e7gKLimJQG6EyyfYYUaBmFb/2CNHv1a1c5CCB+MLbd7sJBwqvoOxu4lLhYC00iAL
bWdHh9rNBsPt0lkE1pj4NCqdI5d0i1g9UDVAYjNrcW7UooaAjLp1bnVIGp0dRuXd
+nqZSbh7gg74iFQpjOvshZajs6f/emIf65bGWmNw2KREzgGFaBV+uUgKVrJKgCVS
fN1VL6hMnoRDOA5UNFUv/aRBKvmJbZZRj0462aDxf7LugHJZkhs/p01hvlAH2GaJ
TllwMOKFQGhDlxAfx5rIkJz3HbZVbwL3oaLdYq9EijHcDVujx7dcc7iOmOu0BqmV
abk/mUniV++Y/+PPEWM33d/6SBAvBr2TDDrYq4vKP/vMOg+cJTx368wOe9zI3qBn
co4gSBwR3nBUWRt92hreVvgSHQNtfygq7HIQ0SCSiOdHiSVF30Ht9sVMlce/f3vL
qHLKMD9HAnOxkIXntikOWBcHd7z2B+GoiGll+RO0ORhbWwT0uRv+rNPi+gTUIWNV
TmgX3IeowD46i78aiEEH0FT7NhreXwOouDjDJ8/sETAO5BEsOB6zEqeSyUH/UUQR
ZkEy+lE2Ab4ytXOckuACFeUo6FVGJDfHs1mOSzdlcy145WtnB7Zps85BvGtJXuRu
bSbjT7IDeLBYjJa2J8SXhqwbEqrluyFzBNOZJ70fhoH7keDtFVRS5wR2wAjU568H
2e45FzdBeoeUoGaX+u2Ie5DeeQmJ2KTJ5CL5gjhrbul5M+uxmuOQ30aeHVnzE8yr
AGCZHtLwHelacpmkVabrj/iOo9+s7Arm3U56a9lBodJP0uCMYLt7Vl6txxzKy5wg
cIVnLHBx7Z+3IeEDnxS3jOGoqJ+kWV8BGFf6tsw8uAT37xuvhi6NcS3XT/UE7NsH
g/1rOx3vfJAQc29gZayp1noMviXXxCw7Pnpda6zlGq4GfZEIc92DTmnjgRikU1+V
akj+9gWVkmZJq+fi07wOLyGQO5YNgjH0+ia2S+YOpTfLC+vhW/WgPEJr9vTDbIbi
9Qpcps2G5K8XIk9JtxnIAXhGQRtdrljG/w2oa5ztcs7gJrSpq2Rba2aZeq9BEB1H
4FA2PAZ5/wJ249kPzsO/gC+Lu94nT2adClQQitH29irJHH7uu85pPGGQpNDp1ITn
7Zhr5FJw+b4g7or4unC4FJA1PUUnaOrs7ePCHNXaWH0Qw86djrTW20HgJ5r6yzVz
J0aUe+VYd7kHzYQ3Pek3DxPl/iTAihxXvBeJPcCtx/3JDj1xN0EdP62v2C8v1JIM
t5fc1fLJlhMyp/AVqHWqClBWddcuT6dLh8BBkYWo/3EvOjYp42Azh5ZHKDAz8/6k
WeTpOgEH7B4oNpYaojpwAFl1fINEKQJdgwzKgZanD+G0xlay4vXsSp/7lvOL2en6
ywvy9ED8iNQJWt4ZO2GA8FtmfBqF7w9VksAkTVtQTq58XwgEfi+GSFDVuBIqfyEv
MzX/V0aDktIaRsYcUyirEUBpX3marGd0wC+pmbBFYjNJjjZAo4LNdfWAh0Kd59gS
hd8SrXFC+BO9raaD9Qs0UF3CSl9vKMoqjeadwcne63XBaULCNxjIlwtt3hl4nzf9
TT4R+M1lWZN0HqUJYjsEZX0L3d6f4/1qjRqDs1ELPsD64bw3xxxtIOO7QitJQ7ck
L9G0KlZwsUrGJOfI4uKGhx15wBnyqPXdrxbUwU9okLEzcJ9IPtEKe2Y+NIBJf7Ss
b/tqR8HdDGjSAAsssdcWGqAVS34YULc/lIzWpT3dcDQvvOpecpJnxXNRhjXTTNkx
Zx0vu3XMLsSrbkpyzH7tjZEBAb8VNmCn40vl5H45VttowJ5OPWeFi3XuOIPOBBxp
apAxL0R5LeQKu+B1ucvqHqT1zjoi3wjCNaTar6JkNuHjpQ4Eu1lrzHuk3zLlXnI5
GA6PcZNDp40O9nw8SfFk7ZLHa3CL2bknv1fXbr5VDHdTv9Cm5EgRJ9ilxYDPsImV
4NR8JOq4TT6H+Oqd8gygmWEjaXS6p86OGDY/zmE4lHzDWVR3cnMRzCuhsiu3yN3R
M4KzvU4MatVIL01HnxwFakZbjNuD491yaPmWomSjWu4EM/Z0Z1edd3IEtTJC6MOD
WOfSTpl+ZfPPSkmLxOXHgBJN38ARsYZ6Bduee9wZ15YwjFusod4ra4C5WuV6aWeX
n8UgYvgfu1bbTtzE3qY5nifINVcabxgkZjny6nO/vl4ceVcgqK7fNrnFRQr01BBm
436dYQelsKHtO5ZGdy0BKlxXzGIu9SW2vOsMhicWIVQrOkgRl0RoZ29D0E4FCtJq
WOvZ0hBUZ2eh6nxNnka+ihqsDK03Jv6Ji70Z4Aw/nK+Gk5ugkXJ4IoegMM3uF0O4
UdwWUz5WJsxw3gdNl+JzpJQccsfxEKICpVlR1xLgc37+OO2LGZAQOgS1pmx/NSEx
h1BV0XYEJEmH9I+Wb1s4pcJDlKtPk+fnFCWbBTQAgiUTd4zytLl/ntUemAXg2tku
dnXMMTwqOuHv4pZrKMxmL1F1JFeE4aNcOhIRGmX6k4/JuPHDpa/BhqPE43D9C6fL
0W8U7N3eEMfVOkG0kZSZAcY0EcXpQNdqmIZdl5Fygn4m3Pqx45799l/qhS89IMfO
EP4qQUMLOUiGqMIPxxKrEh4OAIorBHSpUbO9JWLSMZ93bYa367kozcbQgOEQjYGy
rHh5OI+Hx0yo3qJVm1bxMeONp1PKPVbyOxf85IfX2PGWKJOTei8Oc1G7xTHRHcrS
U8mcTPO7UHMAg7Rg70g4DkUBeDBpkYmj0VoDvvQbjvtQjskizAif+TVJKqIj/VpU
Zg0axGoUUMgpl0vKLgxlvGPunpCY/AzCxavFnRcDVUVz9PYXImLNVp7L1n7h3EW3
HkEYrKKKjc3x2OPMEhpgnqBB+NYwwdf5uuDH83tXaSfn4f74OgbQXD+eY283UKeV
g2U+UsrGQ9u1Wqm+mzp3IXFS/eVDIMBfGBX4AmLsDzKsVBth6MsDDieHHTtpEoSy
/3yXhdePfuu+NkpUYQ3eSfTm5y6fMsvnaBFUmrd5K9uGSd+hZ2L3xjAZlVuT+bEg
B0v3bMztAZtghXbz3yTwQnuUIWk6FhJMZLJEpdUPATR3iu0iRcccgLJCd8/Q1eI+
eHKFmOJyklOYQK1ogrz2LI8wl5ySOjVinChULXt3DNg81s3hWKuYT5M3MRGuFjj2
qihGmXcxBy6lF+ibl0eM34woColIk/3n7AqNtFwVGEJ9QpOLZH768Dlte+9i+6hk
2WSh9FufnEL1UU12c2gyH6lVKSq+GTmjg7YvXLqbdmSAh7ms4DU8FDkLDCVN0vyI
ENkK1k3q+j9ouhp3TD1uvDfro7lxkvbVkzeApCE6UFcvE0yuSaakkf/zwOkEo2ob
fVtN0NS7S8HROCQ+mCucgHvZ+6pF3Hy4pWvVNKrjyz/dBktOQdEyVii7H3kyCF9b
nbGfCInkEcoGDDLlDqumMvM/Wr4tzIo6fHWOZSorbeeTfachVc+LUeWaxjfkZTLI
xcBtkR72gi5PH3oS/VTL+DWCaSYcJacLM+Eoh/Egur414x0fA+kwyDLTHeHQPE3U
kfmnCDK+Xsw/dJglHVlxP2TxrbMeDPP7yiFdiVAbhdxr/23vywok5uX+zpt6PsjQ
iFwVYTcowipg4P4nKcFqMLeu2WwKhi62cFUzafsspaQDZZn9IhZ3xfzOf2isq2+0
9RaZQECTPNEw+CtFqwAj35NJXCNTGDrB0xKzuKGqry7FjHlYkKiw//3S1Ou1XGht
KmOTzFGKqAmqIUUgnvRjKun70NcT+w/IsIu29eA0uL09vsIYZ6pjxur/DjgMhefs
srkljHCyoxk/UCHOKZnJ5UfsireXqDBOaioWx9HWuNekHkQvC5k3lDQwG3aIMR6Y
gXQa7cCL62L3DDMQU216906NX54kgFtjzfIR64Dc2JWWGfpwNUGBrz/vTVNHb3+T
5k5cJM6MNVnO6TUlHnXFaJoRlWqCYzLrQmu4t/0Fv6iAVVMTlkWiyR93t74YVZps
e+BfFqP7u1P9cY3HilWN1l/uxtlpuLyyadopAPgfPpIVhAo8SidPyCqcJXr8MtYC
eG9Mp+OXq+7Fo2iU1A7tWnoEdyqeILnWle9D1Cwxab1lyzlWYI23zX/7QZGrorNW
Bsb7dqv/3WKGwL3Ze3jCFywvFLNGKNSLbxYctlF9cpUKd1IaOq7fSCBAGcK5ftD0
Z2ibexl+UnAxOGfshcVx8Ekkt5mBQiZtwGPI3iiu8OT9kyVPQhdx/cbMgP9L0fnx
o8XUe+3Ek2onoTP3r2KNHS4J7OzdrToF4ikk4Sg5d0ZjiUSR6KH/C2/gA7BcMIRN
x3BdxGaRzQs2KqfaCWOwMKGSN6aebdltPgvtUyJKxVZ0pZumXFyOn1ppo8ixzXg5
BlDhGPRn2r4xFXFeRDy3IDaJBG/GEGyAgKrpCZJl6jcZ8sIl8brE2bmDjcegj4go
HO+aHJsEPW9uR6Lnprv25x+aIRD6/7V6fo9b2H9+PRZ7PPkElUk7/Sbyv45XqDk1
vSHMqQyzowtQZESr+x9TqsCOac+xYfCX1a8z/RvH74Zk1W5xn3AAetyl2fU1d1AE
ygR5juqFCrBytnDLoDic+JgLuDHtIXnvuk4cba75nx+UPSvwBI6DM7FNDluS5ZRG
oJDGfnhyccT+mhjrbmTkni1f8pQHosOFJtyVProx/K7UWPrbB3dJ2HwIaMM+H4zl
5zD4yMkWLGMIMzvSg9DFebf/m659BHbMdgHsjsZYZBTrbU53cQZzmsjKtcLpXSla
BCytLQ7bwnuvtOT9yQ0cxuNlL9dZOdIsl0sFvvr3WR14BT3imczmqDRZ19nLTS5a
5apc4V0NQ5vpN56skwbg9EeEUf2Ya9NYZtXLQxPqS4ef1cusxvG2d4X9Fr0mTN5z
n9cr4yIyKCFLFe/3fEBu+utWZ05oVE8lSBnm4d1fmTCvpeNNUB/RvaAoQ1aF7Rjr
Qqj1QgxZKUOXVLYa54uvb/yQA8Q9TRFYVgqGS4mc41WIfHqHw46g1fGWS8T+wOSD
ih6siHHGcA6lgfAw0OamhaqIaw7ABN7uYDCdBmX0Iy6eMgv+wN1mGNO+b57mlDg+
gIkEqo8Uml1s/d+u4UQqdOa7GmrSrkJW/q6PH71ToqoCVIuCenSBCAt+bJAtgH3S
P2W6bFOSszAn2xShMN7ZEbfwvTzVZb2P8B+gFacCTw47Flv5wuKaDicXCXXlSwXx
xK4HTs+/kLY8bqy2yyTUooiM0+LainNem55iFQy/E+98WdAIepHLWkqT9zYhi67n
f21Sm90xcAomH3FpdZEdx+w0xbW+Pw8fK8/fohWAouO7kuXgazoOf0Ssv4l5B19z
xGqSCjlU3hwvHkRcArK2uwaB0R9XiNoKYZXd6e9sAm4TqCKNLoEm9Wv9rC1eDnjo
gDrvZ742MijXsevME9dSgFoMA5glgPUdKuZ8HIxvyS2mVBCHZuSghqIYia36nqiJ
qQIxaGayk2+mVG7qdid+MJVClRftrVVQXkK5bxWAthlkW9aWxGmb0eSyOiDOeAwL
dTE52vfhi34sY7LveX5mUO0xUk3uKjnWnAv+wvuBpzDdmOd4FoUoaGvZqVxgUMrS
zRvmSO4kvFDLX5a6eSgnmIRuc7Bd/ddA3CvSy781lV5RYDk4k6f2uk9SrWURnv2d
WRQ9dK7HRLSTrHI03pjlPTvwWkBs8+CIDL1iBEYL6P8pq+bwpRDj4XwrIVUrDOMT
W/TJJCYAmBJvIBn5pFUMhEFbSjUVrW4yjSF6ttlGuoWZ1sSUFsiZpivhMhv3JkYw
ZieH1d15PWqjIVY4dinCmiNwTkJSTAq6Ie0/foJ8KFfg8v40tyDfyHPcbTziTzyU
sQDPcEs10Iw0jMqE2uajB1FXWqTDk3KCcpuP94Bq/Deu0OXgBzxWN0vhwoKrDXzv
c/5zlTR6lG8ESaTFtALPZw86ZOSLBlu9ruIikCQbRwZO5r+wp7TARF2XrDHODdW4
QweAkU34Pr7wIGQdVqPtghogqOVaZkhU5R9XjLLyJy7YDPtWaXnNfXfIpDUVs/vn
xsD9yNcj1eHSifpG8wQ+Jua7vSPqqAHxeTCWcC1e0QqSxmYPWieBKUWOvefSwGEn
GT5/Jt4dloICFabSkYo1RCmVuabc0ADmM26DvZM814XB6M54OFOeQhuFCjkHwcR0
6m8A+a7r9zOMHcskWs9TEMwjOFeWWY7Dy4GkuBxJY6ewpx8pXzKme85uCvxYfzsq
KxDWwHSNmiXsK4/DUKIEFamQUflPgarWBXhIVvhphTQr4k+UycijhXGEjtmpkAK/
NLx2rTDP/fqZ4nv1tldfI6eyaksUpfj9UhPQZmTgPqEQoN/3MWY0AXx6TzaxzAVP
gPFBF2E1aOMAJZMWyA3xufd70OJtEV8O6YiQFLJSXM2r721ejFgYNNRohDmNiMIM
Cy8zU/X3Mz9aGe+tqTJLZKVPMxYmX5Iwzk9NrJl7opJ5bO6MX/ogVLo/KsW3huYa
asHwPcxc+hFUeTGs4GhslsUsO7KUQM1wUMqG6DNfbufLFokkoR2VtA8VMXdtQ1WM
QzqZr5sQI2xiTOptYchSEBA8V4cxWILTO6kS9/qALQLBERCc0n/nmCFkUS8x0JtJ
by3pSf+t0r998hwTINvAOrGQv3QeMuyimeIJg86N6Gwafe4irBit9W2MNI/UttXI
DMogpkU0M5qZ/0rXStG3GGfMTCe/6O/ox5vAX9KQOi8kmKgUIR9a763kXmkQfuhv
e1M57UMLpO8lw3nREXanfj/vWNPn+Zw6TIbYyqa4UiZFjat/Oy0iG7JmC4/2wCCm
CvtVKr3kTYrDAfEwIqJgD5e+7BvXZT2HFpl60mLz1Gme5/5hXfgdu0CmjEBrAyuO
U4mA0WkAjJvsiOHMosBuNVsmmwVgc1DE7uqvG1kcYKY2fcR6dkxpwf1EV8V106LJ
Dn1w20h6+YVEGwMOqyLT9rN7xQXq3j4PzrRbU2d+oZr/XFVwgPAOmS1v3j5ltvGa
kkWkNKMKtiRe7EuD3f0hFMQExddinUxrojTk7PHSH6HgLKqpJq5l8DhOJU7l3379
pwVrLgePJ0grYCJptdJmVrSHRCYvNu7jvQIUpU5u/2jmoR6rheaQ3S6hwdJbTjve
ToU1Wosud1k4y7e6Amp3wjrBziE2Efmr68Og6XlNL0bN7MfC4sUr49EMBftmMzvr
E+va4vFilKSmhshfJr85mL+UO+q071Z6lYd/wTLLb+AHx2lZTIZJh1ft+2YZ3KWu
XbIZyzP1n0yjGjlcBAtRcpZA+wiczkUcCvimW1kCcxBNxv2XBu0BU6Q6zWEPt1XN
WOFkWwtUYGYAxmFb5+TkKWiqQg/20fCAxb8B0iVURmiPhDVEEImRlZFvXHoxIeSK
KNW7noDvGbsp1yFRtszssvg1QLLg16GCnzyZEzfG4j/j8H1OgY6ED1xQ8T3UthSo
FEjubUw/H6ZfaCR3DN61mb8Mihb1t6KLYhZjPJDpdGh5hdKj9ovAv602NC4EhDUV
nzoJDuGK+8S6gg/7mgF56F/HtkD3IAhsIBm+ROGzd2/eAyDkPiaGEbh0urSDH/5X
7UNj++KxeC215WXULXpKhWq5pAdTOUjYkKX6LxIj0rE+HACHmH2Vs8UwZTDj0qdr
fHocM8NeYIhS0PJ1WZjtSNVrJu3BB78zOu9u3ZUyAhHqkXat1O92nI/wXXHgvPWZ
zBSK/5ITOsGJMhfeeYNviPba5L/QstdbzPWGOBj9y6a0gXYPinykSNLGm3ZYFVjc
wRsJ5jD67/4XgZzM1EGsOxdPbuRLGsdJiLC4LL1JJKv4dM/D+uC2T5SlyDlcA8hl
8nVFaQuRPnroW/1oq548Uf+dwQmtvJUVFnLAHNh5uPp5/mx1p/UzRm9EobGC+bq3
dbvXxqWGGSqOVBr18mtx7jBs+T/2rNF8o780q59Hg0NqIjruaFiEfdtRqlwrdmwi
vGEhuj24SZAxVXQm4hjLoR+mDMa8AgCF7mgIxniw2n1T+2bqmmUea5wGjztAPKhx
V+BBV8vpB2bv2/9AnuAg5dpMGsvp8CvAZFv159aNfRlWlu5w3lKrsTEUuDXKEdRX
MMO8pc/zsN/XHdCymoF0F4uuO75p4HdKkfdq13cd0+YYbFdZMqC/KmfWG3jPNHrq
cXcZBfA1UJ19PnwBHIhqj+PO2knaekyE9x/n5Krf+50cNlLY7nljA5LWXnaLCM6Z
lAaRd0qxOiU2sg4IDckKDuxuYYmu68z9eJFBXjaG4HCvcu+y5EBjrnInJxFTYwFf
0+swXmCqnGFhqHHFxqWDy4z11ttO1zF5wxXnX8l2qs+zfTlSuzMrhPT45AwxEqIS
5ws/WoasXMx+zoL7VtWLBmI0jbFG6zTwZiq+HOueQT6R+0BrgcQgXlmdyKb7hHXJ
52oxY22Xnl7bbUizKfJaurWAbZ+LvYom14hZy3J5EZMHscJ5CNo70NtHgF1LRD3i
AQs09eb+GGh5idOYp8fri6Pt+u6rVza003z9k96yAghTBEsA3CuyIySEkOanBMbe
oFTxjEwx9So7HJYCJfU6xAmTXl8/0VeL6iy+HeY7tjzeIjyUpTsQkxVXkWnLdlGH
IoJZig5yB55ocUvw3G3o9jalPFFYMgdd2cray1Tc58qoRVaeRRBMPKAqp/0sBrVb
O2qcdSd4QHABRwZ/6XbhnMepAQnZDEd++fIA/AoL/ll3owoqwVSkyH1uVTClxz/q
5pTqJ8DkFXA4XqEdq5U4pVIKMeMgOinWDU0thhHbzCk1B0YVx1Uhpcb/L4kRMGAX
KWnJ3miLvsYX5sHlkCYdVdS/kNG9//SvGi3rREhWaBCJ6bodsFv1O9gsFhgCKSby
UPnhxjXtMKG23AB0YIqkdNmYr0oCKjBAWqbbrBCN79Np5KhmLluDPEW2e0FDnMKX
nNeL9Cff7scoOs2IHLoKtuMJCezBVqAzcrGh7M0v12s4AU1p3+iu/Mkj0AFjl82a
3W1zcj5KV3utFfx9q9jnFfdCalpA3CzYCiUFR6q34dGjrjO0rhYCgCZ8Loail0ZI
h37NY7AkhR81puKQOr4XVPGEBNj8YF3vjU+A/DeadRwfu5AGUU1NjEKfBcCD4YPz
YJ2nCBQlauh7qDEFJNXjD+nO4TyDPCC3Jtx5BsYX8zMeRoSNDPWDaSi5oZcKS90n
eA2XMvtSVGU9C69ZJQYnZ1nsLSi5iPFn1vfbelhQzLqRuzT++9G2k+9legwGwBXI
bsCucSH22MXqQTvhccaVFW5TDQT5lsKEDYEwQQxOEEACRRFCMudNHpQlh688fmBb
szXkE3ZQtR7y7CzAQP6VMOKhEODDD+rHPLrB607QvUUimXLe90kPrd6r90qvtBaj
+hrBy8pj+7I1JllREj28QxKyOUyI3OAEoKI1mMYBTZvFpL2wpWg/SDQR1MtWhk2a
j2RONaAM/stvarG2Myk1B+AUOUPCVqbt1ylHm1XSbitlvvo71vxFId/7L+5vQUKG
t/h8l2lIuoD0Am/b2i+B/RhoK6SRTTraLQskAunPuUME+2IKfQVLPeoMXOX7f5ri
YINu6XwMxB2NhiqXvpQY0dGN94R6cWoYW/v7eVyQkD6WD0/y6tbgtgFZTGcqjcJ1
VKqKX0ZrkeLaR/DKZRnftLae+1yQA2yh+1A0ZgUaeLWhLeDQUF9c/8pMaRNhKN9G
QBXZWdnr8pyZ5vBu1Qe4R5/iv/8qgQZ+YMsn05a4Z4+cNcGjuq2qWkCdiFYcQUmK
FVwKeXYZjAPrG0iDolCH9GY93oxdkCr65XPzJIERhqvkv9idmJIA9MKoFcE/7AOX
BRhD8AmL3dTkWmvh2Z94yYMEgOyJzPR2AQY9TxqcehBNHyuV9gITQ1rgNM9dBLHW
OaEcn7gY46V76bbbCVzSIEp8OpDakbfYo9NHdjP5pO+Gy2TbjuoQy5c6X3vPbHqM
jseARg9mbBBJi7fwLzqG/WPnjltoJ9i8PLh3HskNMLJIAXuLhge5agTc6ib6yjWI
19PQ6lKW5f36QxYQXr4qj90cFcop4TXvwC3k3HqK/V5ctqmRZ3A77Il11jmGMKh/
qklOigkMElU0JngvzuYOwTL0JM4aYfQ/tFJ29FKa2rUQfZ99T3wun6z8qRUx6qYC
dDm6HEFS+RWlSQGR3uSXfVDuHXmmyjTynNA7IK5AJZGGcnJBd3wEPjhIjr8nVbSb
N3rn6q/uiNCfnnG6R/SvEpmicQDCAZ0KUA6F739hvJiL3Yd0Mwweoo+fIKZ38Ax6
KpvNjuzazkjT/nYdi05rHqY34Ag0Qwe7jGZTu7j9ze/PAWJ8ttlEr9zo9DL171to
aZ3DvyISBfp6dwjmgeLdAVF/hJoP7sbApHrY+KJWGOU2o4Mpeik92kHoD7EeGEmu
NhnH0n1fnUpmG34jxKAnbLYo1kQ1RsNoWPYFsjH3LvgA3xQKNeoIO8elOjSLppIi
H1TWGuoOjmUPbYBp2D0+oir5vOsUCRJ5lYHYgKn2ao0oO68kijeEdqUZdUssIAfw
T6yy64Pq3gdJq9tP4SXQsQp/aPK6occYE5WPXjZDkbNCIfdnorUoPNNgQF4YOjJh
d/6VEPo5+1AMDood+hTCvI5ziBYaZMh+iA6sWAvzBqVrzjIP/u70e/2W02qWQjYB
MGuYXmAsWWaGSE4K/Cyg0HLH/FlZs9H+QuKBxLKeEiS53VsEXeC5B2hfq/1qIJ1N
PsroGo/fAuMYjGff6nfIm/GmfHMp7ODLJEdd19CO9IfRxzdL7opGvGbZWpADBJzj
nfHQpm9hiIbQIhoV/sgTvhl/RxBerzYQvTDesaSUq4Z/0xIh/o04N+JAEoHnB0G4
LlLUWzejmAhFeVTKOmZqrK/vK0DnYErYjoAwbkrnEqMjDNBOLeTMkjbExmg+h0Id
724fio4cWDobgetRJA0umRN51ZoeZKQ6+gkzZoShfGdUcQDVpmGrLDalwLzDeufb
ITnokNJJHGNk5dHHm8VTEuTaNNz6Y6Ocu0VB4f9KPVzQK1mVDNvX/KSK7rX5rbBn
mID0Hz+2mnmzspGjrn4tjbNmnxtP8psI0cCPBSjok1YCPi0p/0lZJJRjjM1jxlvO
YYfScm5QxoF2tptgrODXNLdp4QnKsYYukmeH7OpNM4yFxXPy1rbyWpG9ft4JfUtJ
Yt/l/OeIwuuFbm6COR6PBn1v83qhLf+y5lNtSDJwxTOx3Cu/0nFRDncuO+h/u9ER
FtJEVgowxFn3L4pJHyXG+PzNWmlqGNvhEak0dUGaw5c6pqDuDSjHtKTUHksLsFZ9
VcukU2cwVa/J9vSAXGsGXuTLk11V9AeMLry/R25FQ8nczajRWKuf+MqFaWytPwpU
f5apGLtmKZC4yPjaWW2e7urY1UAXbBoSbqpWtc6YtMqZPRWQAK2ReuqWbiVBS5MR
Hltqe3+IRY/HRaDusc1HQixLED14C4daapl8AP4/ZqHJnv+5wqWKqKZG2Dfrbp3C
ZK1Og/n6D64q3LmzYNdKCUwr0+cSajJipIuwrPZyJU7GaqsY92IrPmcfX1jCGZY5
g/WCEHFm1ZfTeseN4A+B7FeqlB5ncu9yB67FrA6xKHqDI6Ls4sTqZikyA2EYIT11
jueDdUgF6qvdvCVOw/1vBlww263u8xvGxMIjeFBiZdispxZBo6gbBWkARR1oQlZf
dKWwiz7pJ/VwgyUQR2Zw803pI+RQGVzVBXGiydw3C6AjFqHZ5M/HFmB3NekQ/FKY
fh87d89DdpTRcmqXAWDTh71V1PeHeX5XI9KVJYBUqWGv+01CMIDIhGPKj7JejoM+
pRxO06TVtjlqA2FhkkOS/TiCZgm9aJ2T1MJDpI2VZ189RQEoTVbcFVV5f//rI0z2
yPI7sd0tf4MAgywotsmhLyB64N6o853/1C4CD8DCAtbqur1jtCYSI34FI7pIMtuZ
AGBIIyifLJfWaOCCH1jMQM2tFyKNPndqi5uxCskoMjuyXMiueJ4hQQFaAsL+edGL
SmPqpYsr6PsedqnaBRwhUblRNmjck8Il6eNcegwVNYTlRWnn07MqnQF6Q13MMjtH
P/Z1hwyiz8d49m2ZQ+k1wiioxpOE2357fxgWx9rbTs0FaUoqJILqtuqyiXdlPLuk
WTUC12wzhvwaA+eDcQM+vp4nD3EDlOAb3w5ip4DUR8isIyYwg4gpjqYD+sz5Dl+J
6lCruocWbVCbIATdvxCqaLi2f3YZ4FWuBKe8Qb9a5YbVpFL8PO4AKFr8+R3jBXMt
CERRyUKbiv86Lp3XsKD6JBiJ6W9d52j8Ck7uSF5hn/tOTU04KIE7L3hgZtbvwopS
NLM/EWJMBdVPRwr8tYc23QCHJ5tTpe2/VA1CZV7QWvWNxGGB8AVcyoEqKPFybv9l
8LQnvanYwUrhzGHvo/Z7mTIlb82hQSFpFSBb3TRcu0tc3tdXc8xUeJfCmNbCAtz9
HYQ2J7qrwLPBx9zWgCo9U0hB1/epYP6o0RXTVvYRfqi2aAUQ4el9UyGkR+JRPL0D
ctB6jPG6FuUjaTLcyZQd6BwU1AhYUNDcBbL5m3r6IFgh1wZWOb4wfRZFOEOAxUO6
vgS11y/vA7ZY99g2fJHJTGkdRPQM0J6l72mZ8CMvAixvtX/YV0QzleGmmivpbdff
yirO4wHFqPS7b+SyAht8S23Z9Fab6NoGgpautqA3pRHRROhDHI2RmaaYOvLOc4U7
F+cdiJymnKYFtSXxhrswTf54CGyokhr3ZiVar6Fqsqg/aEQKOiS9WguE2DxN9v0x
/OCfxiTtHCnUZw4+dswPC2KKXtYxvqD4f8L8n9rsr5CXZ34PftpDlo9kfu5ZT+ui
DbysGdlY9ywH1TTBZVOCLx/UWbran5OuvqYK+Q+lsFgATOWTCfv+WmmNjz8MV8Qn
ux2ByIGphM66VJYuy2mkOcoPQ3kGf2nA8v+yKgXfSzboVHrXh2HCthN252qJL+sb
SyfUvcHsw2ApCLLnTZgwMw/TB4mD2Qa4HtyHN18/iyzScJdGMZci7z4FJTn/gBlY
lV217sxMyc++9UwKG3rMsUHMGg23RqD0QuXPc/EvjelRmqRqm1jcIjKMbfvr7rEd
IwPN5p0RmuQl49B2GTllzkcGO5Oz1hVfnKBFAfkKyu5Xz+Ph1bfS9jlK/WrC0BT6
TrJSmelDGH36GRIWqu/08SLs2YF+uyy3Vb7z3ACRoiau9N4OCj/7neeFYFyZp9dy
DIYnKjrm0IyHcEnGUr/ycWgph5OBeKH/ZIrcMpzDhSNKExbijIECo9fqDEo+aJGy
u+1QSzRMAXhcpJ54MAR1Co7jJTptKDWwQez2E/Z1j6k8SdUlbUxOj1Ff705jg44q
34u/tMsm/2wQ0vIay6H3fn7KpDr1mx7kAcYf2ObIVdc3h+Ez8rTxaFTJYnZYFCW9
apDFpLDlqxDV2N8IcV8oeX/cBmntcKmVXSgM53SkAkdkbiF6u8c9HWZXQIX1aLEB
zYl/Mx2Ov2Y5ndDWpA7IsQw+bQ+MFYfrDpfuDqOAimB5NqVaXdnYnueW6lsOL9mj
D03dI5IbCqkJGUpikY8aW+KKHFYqpU7pvC6l8Xf7Y/t6W3FrmR3L1s96HGuCq59K
HeYtfNcOG+fWlI7GP99441vzn2ryN8yMEIGkaF6rqS+IV6rBM6+QKSdDgSceMHiE
AZdlmCT/Kf3svN/H+NMe143nzH9F7Jqx8uCwUA3tLs4Egd7YL7gb/mpZ4aV0UIVz
sSiUEiHTjLnNnKwXAZNZqGJHVTVamYMOK/cXrgoisoMeycPjG3KKa8uA9kRw4ZFq
xbiRHP0wmqvyzspQHzGwynNCi5sudEpObmP4/0qn3hMLiM02fqKmRtYsTYR3GbsR
KyouFj8vw56MSEQtvIQLEqb5ZfXxRKRwJ5FRaB7beIG09DV3sy5+kbavsYtE+mf2
fzgL8L2TncWJhMmXNqyQLGgfjwON9+QjwRbj940ZWRAz/83zdwJpMIjfoude+Olj
+xyCb1fKjpCZ+AkD5k4XwjUWh2FWc3RNJ5suJS5hTlInRE5tYnH9QJGojMDBairY
mp2M2/+YrQb7WKiW5sq8zDDUPf6To8mUdmXivYunSA2XJ5s3Im8ElkwJ57S0lLTT
/hqncddRXPmDPAaaIVsgDWoax0bBN9T+p2aWFPyv5Xm9c5gpGmkZJj56ZRdrmmKS
MIQwbp8vNPfADsavawKpHDt47TKU1Ryn4xoYXCJoCo6xxxOG/y2KyT8gFuL325/8
cFyIG61pA/EdL3brndMEexhYIFEWR9fSl3KyLw9lgbfB1A1C2BWu2Bzp9k4REoGN
TJDmNAvjk+Dn4lFhBS1cVEUOI4dygxF8glrSsg1lT31dKr+FafKeggWsP8Non5qO
PYpefgJrIMUy9OQkk06twurmcv8me5YKkVD00nYtp20+Es9OAPbwSdCvrzq0g+KL
e1U4jvksD76oFkU/W7x0hjP4lNcCDI/HWnXjq2C+maxuH+FtOQgCbSxyFclVfGhN
g/2wHJum3GVmdYUpg+nxptFq8ZR6ckbNKW+nBHVmx02kw7W42o4oqp/KfAEOhAwa
V2i6L5MoOz4KVyxDsbCsYE34Ht+vodgLUYZaZICyEJColEs7f8gn+SdrfkPmJJE2
WRhBi06en/TyHKci4mKobIdqxKcV7etTak09njw+AfzH8jYoRQKbowyTh6wJC0nZ
8h1MZhJEz5CRBKvaBgUKtF+7xuqmAAlIViYxjYPSIMSe0kC+UksPxTJGvMHMzGHG
bCY92qMUByA+XbmogY+cX0ZX6Sejm5ARBgeCKP5gDRo5rpqBOFUrSajO8AUzc9SM
RjVsl0s8x1fgxadIAIJL3fA+lz/LDo0JYH2Ts0nwCH+70htKrtyi19amtvgIotU+
bYJx1eaBTKojnQfslrJ3MGyHAEDUeU+QVQF0m/ccwGT1GqiFbl4bpoGxER76CQdy
NfXVGa1hPn5q6wAPFE9tca+RIUlLP1Z5YJxw0xYYXxBckkH+jthp92gA5oUuKvM6
/xtsgwqZb7Q+WRacYlksqnfFZ29HtWLYiDBZPY/cpqrUe0hSkCesnsA+gHQXwH5w
f9+OisQVXOJ5CYJdBYOJV6jne9vNTdnFuBaDaSppeeG5eCjnupcowBTf8QS+whdU
6DrI8RdqnYjIfaoFpm2zWXHkyIw0MHEW8f7VDMAG5Q0rsJxJfHHyCN20a2CwBTft
UsFUucz3cSiCkprfDK6LqfD2qDRr4fadA5Ecr4y9XQxQ7kfwKc8to2kDeGwziK6v
nYfPcoPVWHu8Pno8DgPTvjXm8Tdrgm6Tu5BjOcptFXORPF+TDFWmT0GKAkGdvN0F
MD/gfEy9Z51BxC8p2tteEXzEGVZIzHwgU5IgxdFNg3fK8jjVCXh+7FysGdbw2eBc
CSKgpTQei/Pd2lc0OWeBo520lWAwulvp055o5HhCkp8JCB/oyY/ziGa1ErS8ZvKM
olIM8WAC8p7R0JcS49+Zmm7Jid+98ELeGk0iRQ/Qu+Vl7f2sqKFhgPTeN5DjjYhq
tmFAKlw1Eis6VSvFOKuRv8hnORlJZCjolpZaO3hBqtl26gZ8n8t8NRihCGxaB/S1
vqTMgVogU+zwwdyxJYlqTq95cRa/hszJEB7kboxcc3BoCXKZcXNdMkVAGXXhowaz
saV8c0dWdHegmRbAZeMVYZO1bl/AratGfBrYPpQU2YnTPi7W5Jl8iehzX1u1ZOFH
OOPSipObAfZvcBtuJbHttUaiG8F8/X8bjqjnLDHQjKXj0i4iv1lldsvntFBEE+br
pcdKlMcqhPLBp54xpvlEtgW14dbz8yYqRKakzihiMem/8ftNBC8WqJjXCgSKPv30
CNTkafgbo+6pC5GWEd/XiU8jelLrDOfcHn3E1VDuCz4yKJq8L5c8w3QFZhDi2DPQ
ZQLBhfNFBfdVNPvEtV17m4BIX3o5jUyQhLiohDGwEs2mjtAiV6/a6+hPRWSo+YxB
DzD9vVQnOsOkNWCkByHZUGASvBzSfnJFSglZCBSt9X8TtscgdYPUf1uluosFI5Yl
8VdQM13/gqLxKWWBkT9gBg0qKsADd3WbII0SBfZVDYa5KXVFNVJjdMMD9RsxT1lD
CU/RpQYqnca+Zn20zH45lQuKXzbx40bJpns214BbiEdZfwnd8NOral37Zw8dB+6k
EVqHkx+XMSBwo3LcZh05argrk5W7+2ooajO+qzcHUbK/cT1/kk2W41hloR7GV/I3
rk98F21Gu2VWCELV/iQZDji2aEOLuADW1x3ZsRyUDV/O6T6odCe4hh+gZsg1Z5gS
Gb2Uy9vvgrfNTwP+QWcwptJ0DiiLrHYjXWsK3DmdLVS+tipmp8tymxbkEDiVEdKi
+hq7S2H1gPlTQEtCDbaQlGLprhmD00hUQmkQsBSxievXnFkh0LM6bvxj8ldR2RCh
qBFPT+QHJm4sq55T+WcG/g7kgqEINKNWaFdl3twe+QkOOXMa0YqQDG8aMtjA+rhV
z4JrfUgr9pQ33VN5KblMmGEXqFhKEq+I53vc2V7Kbh6/+ueMFMAwzr1boGezcDNC
hw0q++qgdPBtcUfgC4q8yHpRXVOGBehw1pLGz2T4WRRGq3J/Iut4KscbCe8UqA86
O1TUn+UliOQAenUhhjDkUB5J2AwJoKdNSn7SQT6BhoBGgK7bQTZR/11F3n6j422G
1pl2hMJDzD8/eMXOEKPw/ETuqlT3n93ZmT+bJ4ylYiRTA6PteGMb4Mxf26NuF8cu
VTYPXmBR2VDFkLjOmHUUkRPcPjazBc6XximloHS9xYq8XIAG52LVtlLF6GaXEwcv
pEtoaTJTQEgIqQ4Y5QfMX6I8tHZLmazwMIsT6iNpUZy6pL66OHWnvMTz96WFn8b7
ffct4zKOfuBw3Nkq/G90P2olXWwr2mSgxfirMj3WCes2DhHjSysACrhHCmLaRnH4
ka2gbrNmXHbtdU9CSBhh2swZ9RSZzg4l83NM201/AGpL+5kVvf/8dHylscJUET9R
/NtFe1n1PsgVX752gSBw6s2flNI7u24tO1JrrJcgz8gEasR8olUOUchRrpbJUyte
y7wGEnFk5d24uCGCOIvLuA2BlNFSvS9pjFOwunXZ8BADaIzPKG4gKgNpuKE3ioZm
SXEzpSQQdn09ec+Quj1ZmelBJVZ+QnoRy2/SsK/hRMdkycFp4EIe0QWTjsLSfmIn
RFJMlBku93bGRf82apz2b9TeSUTcWhSO3KYyw+0jMiSuUNbQnE0WaG2i92qfGV2S
ez839tbaWcqoW6F1vBCupDKIKIlYr/cHW0WyMg2Z6eeGoFA7B9CNAtAaM+qj3dZi
0/FvkLpYsIy1b+0+P8jrsttGvVQfIFs04yPxbQ4+XXq5dVF8NusYWmjk2wHX2Rtc
baB6e6qbHj1jLxxFflSgT11GC7kZd/tVQbFBQuvX+QSDCpIb5GQaXuHTptbZi7pE
Xmvvc31d5kiHXcNK9JnAV+S2keCRQBBXAWQ2yEAtG85pDNHmuNmiHxjcuUhgBISe
aonJIWIwTQKfTPsl1LkL8KpyjyNI6kNbUmt4OZZaEkv4ag+nQu2lQsu9q1lyONfw
hSH6EHxDpWpU2TzF0h5KAzW4NMBh4FgL0yLaAFAwj2qKZmuUE7xWA/BV0Be8rVl4
vIIsBi5xSNtDz1E4CO20v1AeCyV/F2+XJa6VWUXxp7u9Bar4zJH2eAn0qfwCgaRP
vrixnBRGlY0SVFnIQ5Se1PJlhSR1jM/mnrSuLzmTXkY3Aj6nHNLifsxQ76ddFllI
bzgY3D4RqsNNDFhlywu2Gtrzj2jBDBBkSVN+7nGVYjnbUyxmHlA0LDyquvRZAlGG
MhCz839tv7M3sWCZVrPhvzDDWC0Y3R7iqKUVfg4dEpvrUX4F8yiVNBQo7zcrvpmd
3WUNSFQpRQaLeouTce65SSP7CdlU2v7G6fjKzwYMzwMgnC+VeXsS2gEFEX3pw1EB
GzBFw14b3RZzPGzzErIIWdw6HOcXGR7LI8P8cZvydoFgHYrWpgzhDPkmUcyWK4AX
tB+vyIZhtX5JknTjATCf4LdNjrwJ8Ww/Ssf8Rd6ScMVTUxCPYNuskP4q+EDEfHXK
dFJZJoTtOxUeF2r0V8/44aPsDT5yQYQ0AONadB+fdCegOo38Sm2axpcBro6Pn43v
1amJdXFPdrOIOVdiTLyhzD3RQEULcX1OgJ2EYW+qKCQ07ymp0xpy7Ij5xJ6l+49a
MkiSFtSm3eZPnC7Rph+Kvk6aNzwY4LfrEpwKPOUlxPh/UrFA9ERtHDPHIohVXvU3
7OYmXgv9FrDZloF9i+c9UdIHYfRiSqOdZa/0MXq4fBEVY87VkSIj7Qt7shVU+oCj
igu5ujVzvhmhv1pqK8YqaVZYvFKlZCTlZN34KFpQXfp/KlVIxeBTF0K5e/GA/RZh
ARRPBckfBNs0EaKqXixOT3uLT9SH3eXEApzis4Ha9dkPEqc1wWrMUrszfKq35mK9
Vi0skjSL7ku7VRhFK1Vd52ZtJg1uY16XgN5lZcjIyxuEDAdgBbO9yQWDy9AZpp5D
qHlLBJ1qt6j7Cg569HLNgQQSeYzIpHUucrIZiAoW0zFxCyaTqUEQ/OOnZlTt1u9K
kWkdaGq4YhB4fQYiHpWWet+XwJIi0OcvewckvuduoT+UXx8QcWyZ6LuyqWbd7r+H
WQaxSh0jjyXYuqtRe01Y5IjEw5vEan2pZzpWonoX8swVwQ5+9qlR7IQ63W3AYWh9
U8np70cRjtEkt/RR83cbxjMmwFHkk8B3OIihdPWRpP/Tuy9RwnynM/TZhyH31Mzi
rv750AKKi0XiRFClCQPw7lF4X+lVyE45O5JjseHb0TnakSZe3/pguHZXB7YdoByM
6xpqG/atXt8amJ7vjCnkSbXO6k8B8SoEf7Us6vNYq7XASH5TQetxBFjC/v3xkN3Q
C6sai+3qj+dPZxLz3SSQBrp0mA4Uy7NCTjVvfKhQ1kushLm4O+AfV9N9alsx7idd
17l0skfzuwhEl5GekFn6HbmN4QcuoXbfflAyZMA0Fs0TlY9dsRVbx5ojdBA3dvCd
iCE/En1Pjg9Lq7S2864LQCSwyZDP0bvKvXQxd3Rw8FBMw9J1UsxHs5Oxbkk5/8cA
gc6Frm5E/Eb6VaOi2GjBeXiOAkfL6zlYiBcRNpUtZBQlwaewrfijPX2A1TkqWg7v
q8N5T1Y4qK5e8mK+tByCGaZ76Pd1QsbwGbqR/uOrjVjbKdOvpjACiDhJSwlYP2wy
1P7JHVLNzpCPY7JD37MQDQdcfY6KdieX5UCL4jE3bh+SISyJYWZt8Jnwp89lS7gn
vg5KbKv5kZiiumDMMFYk2ob7CUVw7UcFYZf9mkCLMlr5tLhItaNOeCpluPudrzY3
LW3T6FQGfC8vff2dmBGx41pH4jAEP7VFimB45O04hh2JrFLI7Wck5kuQ8YqtPRkF
dIUefAsBrjf1shxuin5S7siZqkJYzRDSGqE8l4olvg8I7r7nHIU7olFUQkt39o3s
jTQgt+sxISnx6IuXtaa1dxm31EcVnHp58mSuthaMQY/Ki5PpgibJkKDktJroTMek
i003KKsY8+anMm1DV/BzIK6oVehtzPLSa1G744KzipR+5AfyciaM79GGbvJAyO7r
VxGWYsr0kxQouINvv/KuKC8wbzzUMSSaSMza+R5WpjErEZ3um6KQItfgb5tGdvLY
rJJfbp7xACLpxlGCVsx8lWxA23t0v10dJo+jzqb1KNLYedyoIIhArCqCbqCttYOT
5WiZgunfpmhsEAK55iTdbYgH9GALr6m3ZvxcssELpydO1fk9nAOEztoJ113qvfys
gCYlEHro6EEG4730c1ANkseVk4kHsOTNC8g74uYMrPwexHdc0rIdrh+s6tQPIvxm
rbtHjgtM7rC69x2Kpp0uP5IQgLzRC31HxRJ637wI259vGfclqGmAHoFO8r5hy6Md
RQrdxwvTgYEmJ9wpIKC1Co+uynAv+2ZvM+DTSlhGK6AQtm6UuJIgaMEw75newJMO
a9hOPpucGY4XAWyOzGjc/QZxQJz7pyRXKZ2N/6j8lxMPRVhtg/elPWGGFKw7AcK4
F65jUhLl0ItTUeuRlIVju9JJ3jOT5S3ZtuB74RmXxBmuF4QhrfFbQ+gkwqC8ejSN
3MEqqGP64ofD79dGwB8gqwfJSeSb+fFIvhK3K1BH/AE5xFERoKF6sY9AcH2oo8Hy
74IaDyyrwPAOhH+QP5uc1tQS7qOP+/HR+SxJn41CeUdJGqOwoU4QLfwLcYAwpxWV
+H0em09UHPhLMd2PwPljtEcucK0jsk0WzQ58SLyk5rRUwce7qQHQ+/tyfAq8+9Ez
L+XWj/7+DxOPfcSPyjFBVs0L2BYi5Wp67DDEDun8LvT0CVBvcgl8eS/fMG32qgIp
5U38hv7WwX0bYyt7sT5qWbOfVe4feH2yIudL/2wpiCoYA32dlSBxXMBARd4sLuTg
T7S888yns+5i8BbN8WdIBXWkuW7+msX+Oh6m8R/lweEesUPky9IPcqDgTRRXvMT9
z6QILGWbstDNkyVRWxUFsEO+UpLB48cdnIt8oJX10OWCflQ+sYUowq2Hg+iXfyxN
K1gDNcZFoBYrqTEygzYVlKf6tU2GMXDOdZo/DmH9W3pePEuwECzwrudTs1xTne+5
AxGbkxNd25el1GDKHLmXl1xVoPRLHUG85MlYueXyYBqpsSZKvrTwx3Cq7yJVxkAo
JekRl6kbbVbIk5ojNGX3LH0XczGZQb2THbxIx4FeVe3YNxDxm9fvG6sKIhA8kIeC
NTptIWh5m8mU3wxP/2T3Nqg4/kj/JUxM3uy9hkuVmWmx+QlRmxFzyQOozkszwVAu
aBaoyqbmNLSI7S2KNIA2+thARfndNzxxt938NWwbZHh2xoj63yoCjlm+gldKGQ8K
hHw0gEfXWPYrfTY9qko+XIRXcp7XrH/iS0G8GpFb8xzs8CL63zBPLSgob0V8/7is
VVa18oiay+ILFTQAfTQfIOY3ZQZa1oPAsCDg7bzVJsRazKxlI710Nk523qoDuWJy
XA4A4xsN23i7Dd60dQlxnT7lkIL3i9E8hPHC7spmA7e+fVRZDcXkZow56UifZjul
N2lAnWIo5ojrnmm6eYmC+actWMD5wpzQmky8ZNmQ3prIE1DWbQjV6XI+UKBCytCL
97kvGfGCkJa+0ndmWnHDKriV1XAsAiPZTOplJJqaNhhBk0+TUrkrIMI3uw14r1MM
3cpBs5Ft68qan+3MpBmJsBf1trDDFBOQcEBHutrhGEd43Zxhu7hIKXMPh3eVZtSJ
7MdNSY5vDedYZ5hBUE2X61TCA9xvsB+yv6c5zLRfLO210LacXKm113gVwHbBHzsF
5/WvcTTrUicVl3Yjlmof/Cbg/G6BhTSc0uC0ExEmyJxzZys4mWTaVn3g2bsiVXXR
Z/pbw+X0LgrZ/9I2GCj6chjBfJIyz1oVdWw6lIsD+vil19j4y+fLJJO9Q+MMvl34
Cjt5vkgcjTu/6f3RNBBaSrxkUD6uy7d7V868/f7JKVIJJKbQ8jOjPeO1YGAtf472
V5m18ZGAeQvVu+q6I6JMYbv1xkwC+j9UdSP6B7ssZgnaRt94EUj1MLnDCN43TTxE
0/BXOXk7XxyZ98+qjTw2eqQRhVKabxe+Lf49JZFYILQFsKfKHPR1Sqobn9uREqei
AsDhHxceWOj/RHd1txReZcwdU6dIK0nPf8IdPXbsL/IJckzrAfhsM2f8nBIVFhEq
w353oHwS+hyzM4gPTHQmwTzloMowTBFJK6b+esAdfW2IjmLMFj+qARDZtYEbBzdB
1mVbLcflmZ62IK54hXmrleHGt9bwYDysw810LVHVVYDhlKER3Tkdw1RV8YsACHkf
QrumnMfjU4iMZoAMdAtZ8ITzfncvmS1EDPcCIIgGB+8UOg4QNi+8xqKIrdr1pJYz
fjsOXjS5rAzRepoWNZAqn+iFDML0SJ7G9eTEyofM2p46A+NPdNPCyvuuNr8zMX26
YVySwZBHh3oENRlaFy5urzz6ReMN9G94kqLoXgVd+pO2bHQ7eKPmuA85BtKgMdFH
m/euQq2Z68kfS0I9jotAtcfiorNZK30iLM2qkqXzpwSUy8WUyeEiiEaxxrzNZJy+
qjBUCyM+SUZ0qXo4/Nt8l6Igt8A9CbMlggFS9ICHmgHSqHfQ9je/+bW7czzSz0Az
YnoA96HQJFIN/KO5uEoIizJRCPKutVuZzeX7yShVxa+nn80Q08FKKLjrvVzb4JNl
1Vt6xdbaRa6ufxcrWB1yRBrChufO0V1VJubrEe0cjJxdFWPECQOEAs3YdzPx1Atf
aQqq3VdDi8e4+zuPMaxSZhuidODwZXNsniRIZneLCU4rYeMQD2ygsKF2sTWxZIJi
JSAC/5M9R/tzDRb3FWMcG9YGDParin03tHqX8HqQR2d3Zf3XinXKUOmJUufOQYN5
Zta9Dybua3VP68wTjLqfbIxMxgYUfm64/KA9Xtewdy3rVSz1IpqHYpEF1hzQWlC0
zpfsFJE/sgsvz5lJ+CYPSWvwLdo6/qQvYMq8ZoFTBjiemLp9NfuX9I0QqUA/QbNq
gsMHmQGWkSzj6YgVQhCl/pXNY/KvGkxm1sR2F0DMWx/HaYW24VYhpLIjTEJW57zR
a+Wc7xCWIfvKwYr/dDUANA3PMXYoVe7KNP2lSEGcwhdDqHKCoOuc214JIN/sHzdt
Im/if0zx424OrqZ5RVjHy0e5KZUCjzb7ewD5gMnOKUGDiufYMk3o0UflNUngWbtO
TohcU0nl47v+I2w7npsHcaq7z9CMyE9fEchzlYyiwVep8yBuldjUybeTA2q/wIYe
uGlmJS1XioatxpWnWQlglks/VxnCPRLAF/kIdNZU4JOKu+09S2VrQLT0DCYr2peR
czsZalMrL3QjP2XcR4j2SGvNhCTk/cUaspTrlGn8R9s3iPiZWuGXvJdkP9E1LOzv
764CJn2bQlBrRNfVzEg9/x4jxtgHs26YJoIEEGE9NA89tQmkyiHIDFNbPQetWjPh
RnCHtYC2Ls4qOZo22TMd3QIje2Bs+1EvtnbYOFZU4cEo4LVwPyjwivm0YXWcEcdl
hO5bgaH8ifN6RyWmCEfv4uLnbxMpFiAbiSsLn6EV38mTEpKPyXX+v//p/8Tf7yrn
Lc2538E1m3XIJSrCSwjQvJrej3THE/o7n2pE+rUM1OyXdh0aEiH2Auw66VAp8MMH
N9tCLrGDYo6EASMu7Fz4l40jPkGZmGyQP2FvIQjC4szcqfWOMqvDa1ImGT/lYpj6
02rds7moecbiKfkXPt7zNC+gq3aKOw4veZHcx2xo4/gbcL+vxesdVn3Be1kTcKDW
LoUa3yubWYvE0zpBcAljs7XCvKu3cXfp3+3H90q/DgfIgL9nETVhHFJVmAC+0hD0
62rR+FV5TB6X7BXdfinDCzRk7NQ93hIbLXZeFVW4K4Te34W2Aj56wlMxahBgONgs
ObJB/9y1S17ByDeUTli9Nae7xpfZxHHdMN576QXVxV1qXL+29V7zrBcVvYR0uUV1
Ct2oALN91T4MSConvMHJZlfycyIMNVypApV7UFKYJ+NVnQaEEXCc6IJk9ykGa9Wa
jxID6b/uHFcVV62UN7Awea9QF59AjbsZ2Oji8a9JHtUHpMP1eh7CT1R1BhkdW48U
aXqW40g4ShInorLqA1oOq3QZr2rAewccO14QBu5A5xbIFJyVYKiavfAWCIoDvZcN
qrEfNOD0LVl7UhRjlnJpx8F1XJMlzYQw3WP+1mSlfMKZxA1rLZKWeFwvEpKHAOod
JSs4OqGOsCxH6h1pswoh92WNOh2f60vR4L2QlJqoZhHwtonhQi0H1tB6LcB8sBHj
kP6WW3DJbvGfi5NnUU5sc+/hYzN97wTM/tmTGpnXjYh3PGyUR9fbfRL432Op5POD
TFjWtVT3msQZnVeUEfDjvm8smiZfejoCI6TanenpFgFT75J9VLuD+vtjP1sGYG9a
xQipuqP99Nivs3FMhlFLB0obfJ+ko2daqkqtIODhRyg+dkTGKgl5nUe0OScA9w4+
0EzXy4Fc56CQ+AsYXLWLmb/CkZIMS3PC9h18PcXLM5p4jZclNAQ/NegfqJ6dmi9A
NvZMrZRwldyLcR2xW4flht7by4xkFW7Gw8j2ixnRJ33elYIFY6wf1vEmvaAPWvXw
93YgdBlm8OxwVvhRBJEwvd/YclycC3cRj/GBKqo2FHRYq9DqAVuHBdhDiPO8JQ3E
GiwRTn32lifKsJ0pQIqErpcEd5XiqPyWGHeOCZgExH5XESA18bX1w+tg9sLrTWRu
DBqzMJCqiLkHtI/mjd4pBLHvUD2dSTFkoaPRE+Lh/Bg5/sHoT6fxmDoLJuXdbXWB
5VhAVPmBo86ssAIMl9sZzEkAXFS/GuQGa7xx/PE5JapF7rEE+6/1qkfOQyNQSuTC
K9XhBlmse3NkIeTHnh4ombOhuL9nW2iFqdM//QNDKjJMx3YXgJxt8WvrITRAwxgJ
5jQer6/xj6fLn0cWrEWQ1H4OVqgE443CW+52xxo7r1Co/7VohnbJRJGOT1Ncq+d3
Zp3NX8PoKfpDecxeSoWXiDW45TynyunMHqqBDNl4YKRbXqy9v5i3f72zNbkKKwA6
pVtrQizjEgEACjHFrtUP3MpKhGiIesA0QeM+U6iYsiD7ufFG6TSMiuPIsuE/knJO
Ug04wmnbeXHA6/iNcNY7uEiA7DzxMYsnh125DKSXEtnRM2PjAkkOuN0gX9U6VY1U
SkBxTS6VTEmbixEbnamc9P4fXMC0IDsMWZCDhEuXkuJn+I7ltyxeQ4t8AmYl8OCe
5vtC5jt4b2UH1cmJm0xLQvviJEIfYtVxRQ/vfXNcyUCzJRuYedfdFqT6ui2yIISk
lrNm8JJFL8TIykV9DySOqYrZGhSbBE1FPXl16lFpfugjAVcQlqw/je9B+LOicOL4
n1kAUPOWy5ggg5qiryD3JRpbIObKyI2vyOqpSDEmqDL0Vra984/BPQLJmsGVRR+P
FvwVCOvytZYACYBsW+LKdT97LgxzntrtRcX0NwBiyqWFU8y+jTL24Q1BZQ4nqav6
xvuytggbuqH2Hg0bVCxkJcbrrX0HpwXRRhi5lLDYTJyJPJL6MMdjtjzrzr9Iswo4
06Sa4+ZSlzkeXn7YORwWtL3NfTwSuXxkTMIgytZH9SZo1KXutfg5TZDDIMd8JDzA
m0jAAxVDumAvZas7RHXd4PW3OG1mZE+Vw3h+qJalcjwBgLuxdk9m6uO9a/REvE0e
lEyHsuBOrUsNfcBijutX9BVkeaayxZJeaO63owMM+eQPSo2h1unCn7S9dVULb7hZ
VGvRU6GXF4OmfFBIywCq3Qkopm3uvY9ApFy8eagfh5ESor5EeYbheEAT7xzvlHmT
J+S0ZP13mtaq5PMpkwMfIDbTidOG5siMkyt/pCJjSpGjr4fYzsfWKLcp8y/3p+PT
yLkK/O0Qd3Y7XXRllXi/pSlYgdhGKXJ/9nGHqAqTkZxyTZGw4FeATkTK0I8EmQk/
5Bytqi7QT7Gu6kcPtlvDlbcuYSE0nq3ig4daKOQBk67fSbE9ntlIUnbT2XhKAez1
HmvL8XLZAKDNSI7pcj8t2wKOM2w/lujDBeFo4WYqXSNTRXnbC1kS1tF32Fg2oGlY
1Tm6gspq3VYYPDhX0qRACWzo0nzzozCJDPqaXzgYlhFTFt3whf6rJG4XRn1wrKlM
fqfqVxZ5hddu5WXE0eoQ60wl3fRuG36RQHRAupPq6i6N84HliatGKTRA3ETA2RzI
fbpOTPrPhY/YiCKmM9J+I9lK7qBx9CPz1DzKZht0cHDGtyJPEtJcx9UXZqDNcj3M
/RfOfoyAwTphuEaJ1UPCjI53PaP7EFMhNaU5j3n4a/yOxFF+NUG77KxZ/ixSrN6W
/LcobgM/gutZlZAWOnR5X8YWmbJmcOVLnr4kuhXoFI/jZo6Ue7B2vgzWr2mztEro
wwN2aJeMmbFyu1Qi4lfK9FBi/WkSfJLfsV0RjHZKbl6hWOmzXyW+bC84zhnQt1sM
aIKF/O12K+c2lD7dqSU5z2TXVms4ykiTvh5chK1sQgngIe2uQqdb47nIb4A4C2vK
cYa8Wf13MrH7fPSYbkvXpxV093scHH3q/ZpVe7sbfDRNCXlE9bBvsTUVSwbBwJiQ
lPeB5i9aD2y5qbSJJPShRWSKO2JHCDoO3TlMCqcu6FLIH/qDU6QX57nEGVphvxg5
02iZ9xlyXYXSMdoStQCN3AthBjvENRTpGVOVTjPfXZMd5vUhS3B9iZHYOJs5MSy1
dMG7kq7fkIGDRdSjsTiGrqjHCl32hBKbUmfsxwulLxNpsyUrAYjrzaxVEFXJCjxY
825QWCiaptTDcyRPkcV0+6J2OH55lFFCYFQmdywvhYbZxQzKXAUVRhRsYv2ERwwg
/KfTFkj+0pMFfDB5eNwyjw3kbuouDmQauB7vFfi9w2KxmXLjeIf1yHRwe01LUynE
w6YAXz+fgaXFVE06i+lwiLMsVOOHuHGnG4BAVFvCtzOC0lWfUx+QqGXrAgdurCWY
yHVinniNciOW1JKVCzu/DA1a+JQ5p0Fq9EgOMp0A0Z0epa8b6Cmd0OAt4XJSZFhV
37VIbjRbefsFVLbU/x4oBJ6VwWciEThY1JONzl2I9WWkItZFwlLLDz8WCT/VPuhR
pMwEJgnrzvq9GvseWcoVBiAWXtgx/pfmkjKMOS3CicqSuSAeSfbT/pFFnz2H4t0U
mBA2IgR78Y9fC0dGzaLzvmCh9yHis1cZ+PDBgwRJDnW/3Au38JXE4Di6Tnsn+RRE
StDggqVJYIRMxvY8T6ZnX9KuRbSR87FhfGB5QBUhuvhO4YVdzCJqc70KIjA87Nl8
pF3qdlePpYZDSHp0g8RgyeFbV8huQu6AxNFntH4Kv2uETzNhIu4OWm3MMyOqaUvP
1wi60k7yh1MVpDZmAtWuTKgPUO5onEhc66/o72iAMblEnVcxSMi3HxC1X6/mDojI
5jr2DSDTuqTLjEPdS7UZJcjI1YtzrSkE7SwQAik0GeDcBK0QYzE+cs+Toa40o76O
oRksTC5YPVbqcoQWnf132Of+Nx2w/C+QvZQykvWMOvYkQVoP2uPWd+JForje4JXv
yuwvA5eEIEu5G94uD5J1aDvtcNUqVTl5NCTOU+vrcblqq+wBA6R0A000jG5KS8qQ
UOLQ/zRmXrsDw/XuYPDuPeYivpta6bNkkkJ++pyD/KedDRu3fx0J3msJIiTtwV98
l0Ivr4i77o4Mw6klAamQ+4WSCBaHQpcVP/6lipYmJe02ODjtmOtlCEtb+u8+QkbU
+T3DRd1WtY2Bz1aYDvulLWe35IGs+aMdVTWlzOpDVp6/+yRW+anLBpNcfAeaR4Ou
94byosnxGqTaoCeYlf1bz/AhQWTVWUa+T1wmPGUDDK9ntX/gTvVGnN0kzZRk6aOy
oe9B3jVjaSzN4OBOADQvVeobReRl7BLWV40b5AEWJv3ViEbZGuv1PyO5e0mk4yxm
RA8ksrgezWvqESpsDHD2GUGoz1dYwdHkb9W/K9dUgVWrb+iXj3wqcjgzxiME2Q7e
DioFyR3RljKccHFAFRHnyJ2f7VC7jjYTUURWpCxQOMQUo9ZBh2H/Rj918vQ429zv
wHfBEj0f2ZSiErjmGcGJ912EaJ+Ni8RZAcTn+z9/9LYDx34532bDgI+aifrwlwyQ
t1xToetL1mzSBhOgFEkdLXkVeXJvnZ2FarSSYUPd7PRIgoIgQrQdqq0Gyz97B1DO
vBjOF8gJ/I/a9rMf7ghGuBsc8DYX8xaCCRKkWpRBiZqbsQKVOIZvXMrGpIZtF1Qs
XlXwztviba0/d2KEQgQAKDvY6fPcFsNr7xHMhTF00umdX6gRlkwWNLdIzA/CfJID
QZpLHLq9fFo56r9s9LE7l3rLszl3tEBsLlDXRb3LviOEqkwcX79gginuOZCbRCOY
0WXOHvUAPrWXUm+H1i6TgeRO0UWbmZ7lZ9oDyZgcwsaSEnd9VbH5U0WkzGpFzXbl
HfQ0ctY+NhqkT46XthE/2OKSsU2wNmzT2nBAdnkhyyrPIzwo9qv9649BB8oxPB/v
TL1KeVngo0bz11bITi5KkKnHWFDz4ti0QX4hp2fhXDHh6UL5FFH9EejdFalWwppA
PQ/wHblwS8AWUqP7WyyihWUd+OUmKZpncWUzI4o15r5IQNzGAphI1V8QNJqfg+/C
glzeSu6XGF3QCfY7J1AT8OqbkEsx2fSYmA3Y1PztAPp1ASdwfXY4fpd7P2M0cVaN
ohETWsgo0gKoEBMaECYtOs+PLNRIOUEnxCeScl5bC3ZWULpLjxuHGGDrUVWvfPJ4
EoSgwq0/YkcrCWM/av1RD2p6e4BpOthE+OnnPx9MNGsPTh0NGHUV76j00eJArZD0
YJeKxThyU6Vgm4KjeFTTxURG7YtnPCZ8qfRIiR80NCRhDA5ykjdkE0CL+0flLX+l
WolkdSOOYvUylxvJvewF+absDa8fqPK0LEcOJH37egV+/A6jrhPhCaooD50O4ns4
BtYO1fdBhCN0wItHHiEWNgEwVcG9Fsr1eaqrLW+mk2UnhFtlhKO3vRf+iQtOdWH+
fReqAXTWMHDTZLMuGyt/nFV4W4gwQKMUG9+2EAi2lZCWnotnVL/H2a1LTl7RxtGm
6n7Z8bsvvpnX9BC4BAjQ7l75BHWg+Glchue5xal9RGtFvuaQVGy+WcBWDokVBnm+
vXBwmL6b4xZishoHJIiZck4kvQaV71mGOAKvrjWrrIiYk7vixeuZr2z/PAN7yWhU
/9Ie6qWkEHUksNSLG+eSyXmA+6Na+QNHVBRFsSpNO6azx0IHQKS/aS5f0S52IIEs
/iEg60TF2eU5hJgNg9PgzfHVmTfmR3+vTin0rtvUGiN4oWopjEgfDmmHH7XCnvdY
Q0zbOGSOHldq7rFNtmF675U3MjxP6/3Wj6WmLxOz70Up22+fVrNUMEWLtFgSXcq0
vK6xSvQhMW78g0kIOcHvsx5yR1KicSOIZXWdWllx+jnUDKKT/taplQe+divJkedg
yftYQ6e/kDC1u77IFHyEw42zl1cGeROo+2b4stYpao5w4i1pSaWXqHTap9lxj9mR
3Q6BO1B+WpwPqUsQ37dvPTTqqMIpQbb9PdiWCnd/r+gI0eiFD1lSC7pgXJD+MnP3
K3NMdvYKJHhzSETKSnpvYL19zH5BbQpLw6s1WHllPFE0y9XX9EfCnoMKl2/I3Znj
j1HUl4c+k0F7h+HR8tpasCpHQiQOJvo+yOrY/FImxEIXxna2CQ+GqnIyjnZQJNRx
YA9OJQqACkN6B0jM/1hW8q2M0s6FNHMQniy9g3wNU2KMR1Q9dFIt5YCg2fvWGpj3
5XlIEjrPkoY8ix4Sdnpg3Z7xUbDTlK9wRJmQy7fhb/0E5VEzPGR7/SXufmwDFMMr
0AQdXsglF2qk9EjJhQbSFKt3L6HOHAXnEus2mvKjOvWiaK6k4MCq4DmAhE08E9rK
AzCqR3g/IePMw+sI312V5KpyLkcal+e2j74gJZ8X3JvWGkX+INwKejaN2KaMa5wR
RMbMLCuuN+gXjA5GeYaMhCJlkQiJA/lXu5Z/TjW4n/L76YjFF0W3RCaDT8SeGi7C
pDNLmyDu5W0dS+RoWDImyadiIACbVeciqLtoM+6k1A4Q29AwI3ha5hgAg+pMfA/x
AB9KFJP6i5F+4o19gsjTEg/OV25YtqrE9wSekDvEw1IvcS/cMrKItVJwAm7rwb80
9B6tbMs+RGdVkNyQDwlTLntds/71HQoJuAiY9yxFVm9vSObD6a6FgSHGXRMooZhD
94HoYfoqDMfGUrrees40A/TCQD4W2FHrCyMdvwI4pbv4vUJM0FJvv+JRTJBTVTu1
iVMugMp8hxQxXprfFSi8AHgh2PuWaCbRKC1qjAIFpNfRJ+dc+C7CzhwGdrSStfBg
w/vhihZMejjoI5GVsO9h3dsFfOvy5FnqJrBVkxowBC+vMAdLq4BjDAdIOSYC6gZT
9LVs5pC/eHs37qGrhGuR70bAUdGKs46/zOCGaklbbau0WAHvK7xXKRt1UK0DExLa
Xw2ltwPEXV52Ui4CW8GDoKOoc6Zj09ul1ZkSnVjaLpD4728/2z4k9FNeP74UqRRx
q5hjFyTnbJlm8Qa3/LS8QB45nY2khepRsS0FWqQ2kHgBrRjELcYITCgRgq0TqqN3
co1Ud+5TysbtRIBYknpcR8LOCnlpM3V2OFAv9EL/3gxfeDklXy0cQgpYTZsMv1M/
zzH0kFf/Ci5vI2k6KZI0mQ3uickQtlDe5vBVBB+z0GyRj7Ncs/lDVxBUZpZHg+75
x5wxzZNfvmkUiEiuvi4luWkxudYHKa5ARFZY9MHm3BZyypR61oh+iTgVw7DalTHT
bcY8TW3BbVESXDGE5C47uEM47FKdrma5JuGb80FxWXUJX7gMa5Nm6i8TnbQ4iTqe
2TOHhUapx3v8OH8AqtfKcOr7qNSHMGPJhn49K2LhZSaRLrdzO52ZyN2X0PkfA8Dt
G35BWhRSPEzxIGQUv3A6xWIKAHXfrPfmpZ0I1chyR1IBRN50UQ2Fe2eVzlbjDmOs
yKZDRkrnwvYFhoh1CIHtxDJ2pDohkrs1dnri8ZVx6+r7KjKk/EvH3t+8g8uGr5uO
7fXdVGSlg8A+NTtGD4zfBRJusVql/ZKcHgE+ffSSAMRDDFFs2f41mUtI9Ul+57t/
J7F3/YhStUCe6f28jJ3PUavogEzOsjevwgH68XH1Jc4i1yYmNiYDI+oSMAw0Ku/o
kyWnfYS/PDjqtQdmkvQszUH6UddudWhn7mK1SUxd1UAKiwE6nyeCzsXRL3E3P7eY
hNT5NR9V31aUNZC3FV2SBLBmE6jTTr4D1266cfkInsl6t+SPCgqIZUcT8EoW3pz5
Bv/4xKiQrifwCBbK8Tt3PXlysWVFNb9r+22Ioh0b5JRaXqWeVGbaJWvNyyYx8+c3
gO02N6EwFZwLtSigdYdyP0S5jY2g7ubovPnO5/MXVlnQDX5OCFyCeyJ0yw4m/tO8
1YGXhKIxNntMl+INDX216ISdPmtLbn7wJyFRSfT6XQQRgWgwAzsVFUFhVugph2lG
ZifF+lS/7WpUzpEbAKuTobo2O8Ohwr2HwOJw8UdqkNZRwDUVVt5o35Jc3+YRaIyv
spY/zn4McbJyhlQ/6GCIFcbHgdDW8aAeylYFCZtnu5TrTpC4gB7uG1mk4xl3TxkT
vk4g/hQyqaivLVzTQ/6YEa+QCiecEITUWwfmr0g/qecrrLJOMcxl3/yj+N0nm/WD
Jy6HQ4mXgkjKMsIerLQtgt0yIiiD1Jvj1v5cFXTpawfy5PaM4zcx2dJx5NRzY/Vy
0cJFvHDo7ZlTY9ErUSuEqdTkdLWKjlMT8hLxAfhv69FUJoVw7eIrPJIGrGj5wl64
SEoI1EfIFtb1V/46P1QowILeBg/PZM9ptbp/Z82AqPx1HR1iSnIJVC5x7cL8ddNA
Or9NnPIErnywTDdvWl+8YdQXIeZawWdDShUgtwNf33Nt+TmsXCfTGX/tRz7q9KsN
LeC8hBZQLuitHH1qPd5PWyA0erUGvtmPhlB7vf5MwqJkdHUmX7TfFr5U8st5DH3Y
eHgwL7OGoX7q1AQ8+UtickLsaK8J59hddIJq5ornnqc9dEW6uzlQb6t072f4x9KW
dPW8oX0kNFo0XL8TrBUPNzRlBSMmzBNKTk95ZoNJoaRZiQDtggtGWJK/gLSGRuYE
3ZCIBLFDbWJE6HYRkw7KEgL43dP9z88jHVrPGkc21ZmIYtULqOMbidypIi5NWzQh
Z4JREW6keMuQYkKNydF6Jip1B07sTUB+EgC/fsuvMSUILKRwp7/kT5bv86OUKmK/
1fo9DwomWHagrIUgxQISti0DVMpmSJojBpLf9gzuFMIjTjw8bWajWwEyuewZJRDv
+LFcde11H+cvnF+RGQo3ctrEMqWj9hXMjLpop3k4F0rmbcqaLO7BBJbPv1zCV/Dt
trb/v37hwU6h2S5D8/9KP6C1El5tgqNMZp18tbKx2t2MrtLZ+60/eidpFrmYRAC7
KSxiW/yroKfwVxMp80GrbAKCCKnSpCzeKOKNjUfFsD0Y6DRW/5O7eW42I14agaN3
CwDcHc182Wd6SNq+0DBElpJltR8O4Sb30uCaOjcOGltquW3ku1Qmdo+UdEKLmu+/
BYU8z4+X8nh8EkW4SBc7PXOEpNt9oDBc1h0D/52r197Se4hrwE4MR7Lb++/vddUR
7Kqar9FITMO1Ro0IE+K4O3Lkm4jg2G7eIA2WFrAw/Rco+Ma1nvWxgEYAaw2SVS7l
Yo3d5IdJrLb8oNpNieU9Gd4ZRAqPPXAqSH6kSYg6ICqbLVqXlKB7q81zwVSUNzTY
LojDYPGi1kj/AmS16mbtUZOx9Z8JKFGIkl4Pxq/PUzINn4nNcp5F5dMc5hoOsJDQ
tjf1WuEft6vAbSZtwc0uzf99AIDdhV6bJCcftWKjpEB2VszrDLoF7uXQhrxZEpPE
FEdANqtC9v0p2WdPxMLYI5B9A5QCaDQ3BDknbhNP59f0o27ZkNZnJGtPOssxK1cU
gzsXJSUq0i+u3/yr2KpTrWG87u501REuUDM3zPe7AG2hKCuLoOrRIRrM3n6PYrzD
DALDG84EBAGhbgx2lVE4UvtVEyi3NRyiDrhTCMZ+No9znvJ7qsgIzpDs48IOWF8L
5QnJLN5AU62omDQ4sLvsBKXGxaLQhrq866dzpC0TNNT5EInjk8xF7LhJM8wRTd6W
J1KboAqMMBxAY+Vff10fklZdcEv5HeuxhYGH9lxi6Zo+HI5ZhFTr5SjUdFFypoSR
8prJTRDqLP9L2bH4Gf2nCvKPtuA3LBfo0DvoLLJLzKXJ7tV7ZaH3YX6HYDfCH5a9
Zeo1GFcZDC/PEeaNxaTbtBBEf9C+PUDgpgTq2lK9isk1o8yfIJdABZHJK8gmPXq5
IIGMWbJPZbA0qNllhxRJvE4AyqW8ijn1mzkp3hAqo/AuQhaP6mUXMA3n105d036g
lcZ5TQbgFdjHy8WQhgTiTmyY7Tws6ryqblIBXs7OrBviHVWCJLfTuWRafKh24rN1
Ug3oDkwohSbdjJs6ayhGewgk0u1NMFXJK2qBtMQQxQH4TVZDlqU5WHWxDPRJRa/X
rRiFL5shMzZpw7YCQ3TsxKIo+2wEG80LPTA3vnrVoz1/wBZLeLECz86j1mZGzERi
lM4p0HqdGuB3Y9mMwSrtcwp20ndSO86XczBpALe6B51hvpnMQUGDqOhqLNq9qBpo
zZI6M2r3R0rgMhaPlGdeq3fokarF3spZEJjfs4UaSYaTHIQ/AO2FVhxIr0VcqA+U
/jLGU7umYORvz63RASRynN75USp6JFe8dZppBzIbwtjq90xCgrk0GIAXN7U14hv7
QxFi4Fut3s6A6wqeGfMm71rbIXAH0D6/cUqVzYM3OPm5vT4hlOQ1ke3acrr4eNmn
BIe0W15BIwfi1gN5xDg9xnMD+3IPYHXnmDDWo6NDJz8/4mkSD7nerTs9Z6+KVaBN
Z7eWjY2Aj7zdZ1MPFgbLwaqxjjo1Izwj7eKeBtQC/OxDDqDfkcgDtdXPiAzXsvrw
bJVuijCkeqavOfQEKhxd2v/TOb/Y56GrpjKYbWYlOJg9oNif9mofflXktWywz51p
SRUl8bnJmbLSIzKPNlOOLQHhDWJb+b4f0CWivMTF0uydJnN108mtrK1XxUzOBl4R
VxvI1A5LhnYi/8RnkPzZi9LaGscoLQeynPPzCkB2saJS2Ug4WrHPAQDhry17ai/d
w8M1z/oaI1UywxIueY7R4+Wm1r7ur1Tq4iRsHuLUV3CN9PlXb4rltIVB/Iff7ooG
MrfexK8cYBT6pnLzLZ7x0UZRgpcJU9AHjSdn4Krf0P+JITVjMcgwBbi8Kjc4Szgu
YQsGzwClkA5xDdY4pJ+IDTA7zkAHgFXD9yS7uEM0HD4gWpy4/vV+m6IKQeXyDfXJ
kpygwhaf6ZvrVS28TbZZDgWDuS3tgaevDbORdHkbHuKL+s6WhFC+RsK5SDYP00K2
183Br5kOBxH3ZaJDXAT+7wrO+oRa80NKyUW2L+XO+cWKgNwhgCcN3XvxyD996ygg
kkgeXD/W43iuRb2vVOUDRO0aXGfHFrqfyeAfo3gplXlWgtJDQnuhGLQeHDRf7gY0
F0g6SHWvG11tkxBTYomKV5yPrgMIKDdQgdshzeyYnDrdjt4RFRMho4kfP4YSPs7j
SBzTYAMjUd1u7kufmeKurc/gZ1hWaXq5TqB4lLLwG9N/ospwtdXSBhW9pP64F7Uu
uc+oEvRRzCJI9RRW4UGlHEJril8bbfsZ4JlorCSDjf603XMmPCjg7/WvcUJW3j+Q
fdCHoqLPyyn9FluOuNxktvRtIiCiTXaopbjz95z7oIexzNjnelx7gVwS+XCkVyW8
1JpnV9zHZ0XblLXED3Rdd/ks3cjRy+9o/30e/YnCi2FuLelHAG8IfRNs/C9KKY3v
vcsxY+JIS+1W15y04jDdMgg+fXGar5pUWufB2sR9ejHT0AmmfTTiAK3Z89bqYhtB
mTQie7JLLCRTA2jtDA9jlD32tbx8VIGYLB3HlAdBV/dUFIm/CQpvGUGDZhtpPTmB
OfECKmcdMZTBolt4J2A/hDU9OUeRZTBTQuUlHXLnNylTLMy9Xz0spvyqzEJDSrxG
PxSGrDKA7L0o1PguNLXJoA8KY8nKsL1jYMYnYCtm0LsnpDJ3SvOoEKK8qRAnJk/n
Y7+8X6sV7NsPHMG17yaIFjD7Pzz0M9Dtu1+tVF/OT1U1hIbLWnpK7oS3OHMAUoal
gyOdSv+oYapoUVsrV0O9Xc0ap+25QJELYPYB7o/C0ni99OYWwS+Zf9dSyfTeSG7V
LxhK4DNNmtI37L4xP0cl+Q28dmsZuuf0JMF0l4ddFz08aVTid9xABQ36IaI7KuJr
QQag5OjNTpjrZYa3ISWQAkAMJMPwaEo8bXCJO9m3grHLtAML15SGOX2ihQRXctgy
FgZLS/ZYC5goinS6uhP9uAmdhZbYQYmO6TxLRU0Xm3C//jWo9gpOh2Z3v6MxsAby
79At1L2ZAHYJ57lbycqLAN0oIU7Uu7l+gqse1mzOXZesjLZwhOqWNjGLZ0lfod7E
pw6D+f2Xf/ixOaWy8nmkGp5X9DTcy1aLvfc433fYvTaUiu/hJepDK4v9F+4KdCOy
v+1S7Q+HdUDI2TCNsjo+tsMCSMQS13IeoQ/nVDq5IxztXsQlUrvCDJUlHvt5lOLK
ocigYEEvc43w0YwHeHa8zKSCHM3xB8MuB3la3yX0lKUL14wpeQQw+ct19543rocD
TMP20R3xKPjQqM2fULPgyS1ihuqvnmpJm7GbbpQrQqTzJXrGu5EBP2FzGQz/YbMg
Kh0DeuPrfn02pdWUVi/+6jr79rodLBNiYkW7qwOcB/EoDuNIW1oZVFgole2E04Jc
1964MbN+Cnkl/zAxXQn6c+E0m5t9LLiq+tD5tZXqleA65yKnKp1QlpiXSjhMnvg2
GnEuFeyENLdwHkvoKIHBI4QroNmD4a5m0CTjrw6MT8NVnjh7tAtV2viyORe1SQfq
o5vdmBXZb7jgZVII455dcNl215vv1DZWK9GZRl2b9AelCL35oihCaUjpV1boomSu
5CDRu9MosmxGDkLrFnvg4IiQt2KXe4KIA+ab8QQ7guf9QS2zXzpNDTuzxOdUyYUZ
Paba1yuRbKSP0NOHrGvsfnGWoaC/04IZetzaWBDQe9gNlN1Bf4IqyGXvblaPpVNb
Qudb/CO66jyJcC+avKuDA3v1d3Jt0UXVeVjMMFVK1VH8acdvsE6Ar21rt67tjJGi
tYizLnzQKu7z/0nlS5cyhFx4/+PCWywUewuV9fCx5uUSCwJ/ttOmGDHpc/MX8btF
elqZCT12aZriGVb/vKTBEHrMMwYz0XlrFe0Bkk/WQezNpuN0NU2BpZNZtMKzBysN
kPadKnBYeTZi7Yef8RgwBapMA80NqCj7nd+D0eMt0OrPWXh8ZsKguSdOprYJn7cE
v1AKFRZZ2TzV89PLknfeDW3JtFyPpip8fY+gdi5dGzAmp27zi9pmewDWtvjITkb8
GEqc8waBS71/4Tyb77nU1IObEy/3h9ZQH6HKEEtfx55g2R+ELtV/Dx9tLZBDnAVg
3JxckIoRXxZW2O0FdVaXNY4s6dIpzGST0/tASBMz5fpp9yyORvyLwtQsl/h05HXx
wwwYtWY90rH+nmct6HjTL3w/G8WI6rKhN5fUkQgI1Ord0UafHqO7q0m4Jl7Pi6qR
MvBCQEi6R2AMXSQPqkeG/opUv3RknF+j+KQIoEeIpnCVdXTcUfiAzmPPNRSW3Z/l
FE/zIUT2DIJbVWW4GWxOofy0dmY0TOkSVejeDuPAxVgbgLiwQ0kbWAH93TXRv1Zw
6O2gIKCr+J9SXi4slu0hkTPRBNhngMmsDPm1TuKt3cFGhD8vGCpST3ZrcePf/yZW
nv7HuRXgG3Dc7oOrde4Z3m4KeZL6nXoHBXMsOrWPPq8lsybj86rKmsHFfTir9I1R
vkJM6Iwq9fkS5QQxfQhRAYGHv+R/gbZzTTuZM+nQAjvAu/0kh8zDKqi9B6POv9z9
o2Ynk2hH0snxyQbPovzA8ePw95YMKb6YjJ6nh+yVFRJjMkgxjMe40XYjjGrDDwvG
wC1UAX5q+rLStdDc8fFkNRk3FD84kduzOwZteQaeCcLOaoDLWKKe+nNpjjuBL34r
GPjFLw/iNfLzaKuYhzJcXF5Z7YzbYMR0Dw8GEcmVVBisii2hGDY6Reph8IWXSbot
WOzd6VeBb4G/lHc4Z/i6Ms87F6X/s/utOjVUKBQb13oCE/KdHc8dwd9x1CL6hYwQ
sLZc7rT6vBvM/4trc4qHM3/AsHmTU4CDX+QkdOIUFO12WrPSbqorGf6QVEOYeaYn
HaBiw3pYHDKGWfYZgPcRrbfaPWO1/XMAQMZlReY8g2QuHfFAT5mXkg3tsBsFoI6q
xrnTtLhzE/4CiOi4+eRZsp0yN1eqOPJqYgSRiuDBxkeBJmx33zCxhe2Xgvl/EYLf
5uCRgijQiN2BuEbbTupu3rjzJeXP87YxFGEh8+Xcm01ELYOAyaaAVTF40w01SFxf
nIJMiSIpi+mFsqXnkRlIm3WMzyt7dCv7B+EFn5OLPfeLKLBiXpFwtGAJQ9yEg0AV
XTyOyke2nUUbe+P8Bm3wsY/zMv2e6weSzU6B0b9F+1O1oVJq5Bf9DwzamyzBvUQz
kurd/2dkz6mVP3AYGfhZU5hSGV84tv2/YQ+xE6BJnAzj0a5e9A1ednPphgTQ2cUs
TnA9MV9mHJTK72XhSgm/dKURT8dqm3wSWBUswDJd/I8LJY7llrFynj6K3E2smWrA
LRvlxACmDtkWE+FcEario4wSTvDxBx1V4AfD9adj469PZjiGGNGp25KnyiH86Orb
TleYvH6+hSW2psO0PKr3Pd9h7tzNEMjevNFbfFK/ZV9NULy/l0fw7U/g0q0QCI/V
SERQOkE3PIDIwmQ5BWkJua5ck7IWpxkHuD747wMwrzNxrqT+idyp+HabsMMBt+lV
GuHQ3oV++auMop52+9mONKmIp0/u+v40tOAkOc5kiGC74GaGZ0yOjIRQZijB3iKx
2CFUIxBg1YNx1BxpiHKSdJmZxiKTKwieOqhy5dBOqERQZFByIDmnXjGXWiLryH6g
OwRHo8wvMWjNIPoolmhEov92iAqF2qNCyIEZaguKlB5afKj3tkPAZl/hTdDtAY47
UC5QBCDWbbPzrjEX6ZXG//OnEnreXYqidTmUYh8Qwb0a3fK+0nXeL4I6AspR9f7a
f9kszBQaletFVzlKSj1swmRbtaQhzbJCjponlF+IlQ9kmzhXsTEm3WSLw4MH0AHH
bAHUWdw5ST8pV/3N/3B3PSseyMaumuc4Fyg+k8X/hbHCyL5HECAk20teNhSM6zIf
DetmrBMHFLr2cd5GH2JkSZ5KApkRfCwRsm5ndIKOdN+g5LMz/thUK0SZftNeBbrZ
JWYC8fJOSad2BoyfbOsP+5bJhCdH180/Ad05Wiywmr9O+5znSShYBiSnlreL4yw1
Tf/I0Bg1ZYzgR22II0BQhsY9hkHP4Kpc1XUIRu0d7wY/9IGl2BwKbK8+/JzXMwmX
BNQARfsYk5OLd2vkyzSXxxPCFROq3Db5O9ZA50svC4Cf55o/zrOHajYdxUaYJxI6
1GdfjvjmS/MAika7m5Bt0OF6gPtXyw0kvv08HHMfclR74ljBEcioq7URS3j1aNrO
/Gfa0kekCnFB25B7AP7k1R2hqUJFZvsAKGmY5+lS6QwLvPlVoL91qbq5eDbDUqia
H5jM9L3m1YAyxiv2qvU8SQKqFbnYZxfPY6fP6FlS+w/N/DvD0tO7tjSCO+7ul9uk
p2CPpyZzTr47ozIavL9ua6fPWaEkBhwJfOdEulApQcuKm9z7zakpoyLArW1TRepi
lm8lEb0uR/YKNp31ttaozrJ34Ku2kLXhAcuHgzIQPwV073ayFeWzBd05c+ETtt2A
ProOcg2auaUiwfcVkeNKvb87WvUcg3j546WbvdpMg5fCGrtQyF/10/+7K5owKZkh
T4z5cN9+bz7UW0SRS8JVrLV73AQuJOW395+/gOAbkBxNAzbJGK2n/A8pZkPcBvaT
/V9Nz/5vkJmb3Yi4JwD8gJKrmW69jXKLGc034skgjntjasOTaNx9JEgA4+87suHP
JBgBWBAZyjnn9hcyoTOVl+Akzhh+waThWrXGyfkPaH2CuWOTgaE8R5GaT8P8snDB
BerLx2+a8Qk9dMXUrwc4d7xIknRpdAO0p2NeT7Cf7zbv9UyDJpeNaPZbh2vuUAW6
QQVnWV7ORTvd2MKspXx8B525mMFHqKiTzT/d2bfmLEZlYFa9T/+YBkGHatdyVkEX
N3Nv5/YxxuHjl8OPGFZ8041W9h+zK2hvgQoRO3K9KzR4w8+UpVwtt4U41Q/3J00o
C15BItgQbJ5UruMgTIriQzYpsc3qEdpvyiJnCXWsMRWrQgE4yo0h6rYsdtVkiHA6
166Fc9mi8NWoZ3aeE88eM+PdP4LNsCn8IEAIkGhWHtnp334hAf6fTK1M7GCaYzrN
eDQ6kI8xmh8UUIiSuEAFwX6RraaHcKKQCsNdJ+am66/H8yvZ8eyDn2SXgiVj8/yj
IoEP9Zp9PHNhPEybSYh8NnJWXRcqghy3TabpEqZHj4Rxdcd2Yjxc/1e3XbHpRphT
rxh277GySaKNU35MciBz9WGulS6u4PyaOyoEqVgAQmyDT461tEszXC6x6t0U3Jj6
PwJyM/cdVtKCdOHFNTTpORjt0LtTKzd3ayGVyQpSKG+CcngfG5DiQNiqDkBPlE73
XysMh8ixvObEgZInIqh0mekP3wcds6XcGAjmrm52v+Vgq/qN3JQKNmPNW3CsuFir
/h5WCo/sDgg+k+LfVTzw+4Pegr9srkkkjBMhEi4tOAQwNyLgomfubo7qd2L6Zfmv
hh5Pq4YGhTF1OO+FuS+Z2I9Gg1nJfjChobkfzgV8wqEMMdq+x7Uw0FmbwReG+mU9
OV87vspMLUa8PMFvMt2++COmFOhpPfOJMy61sTxbhdzjlQ2ssFasvPPh4ZjmPoMo
1+aZ9OQjAl6rGz3gMYpP2/0JL9NZPf/dsGMG02dpRw0o9wY9uG+/uhS3lOKhKwzH
bhlhf2WlJ2Tz289HYZgIFNATU54mmYYKDRUGQqytdZZPN7/+RG9xK92p/MMt2j8D
phasIwbfVe/14gexdcIKe26NgwAvLnZ2Bkok7+SLdVSIdvF5NjqwBwpu/RON72HE
uelqfQj+kRWq1L/9yDCRJCMlbpkXC5jUFZfqH4bes5EOE+619rbPmYE8kiqUESnA
XB6BsKzvIAwtTet/HM3sHuSr1PUZ4PZ2bOCeLBYehO6P4pdjCNRSv53xaFEMEdXk
OE6R5Hf/8SInG2TAeAKT+niMFAifi7Iz4icS50o9lWs0hnfjvdOHLnCljkfybbA/
sHelWS8Ty6qSUMrhu5wwjel2g/VvnWEQ89h4g5YN7aS8kc9Wt1eYGnsyS7TLb14N
ctiwgk/bGCBUjpmce6MfGxl8U0NffXE7asy5S/7x95uejxELX4ZEoQd6u98vsbeb
7p2RYPdbkoYCRy6q7E/cFOP73H0rW4sFfM+P8JuS2ltzvJpD1YHFokl3T12P4lzM
MTKt0zL4BF0R9/+JwMcUrUX6YjSl7guOvEz4ugmrRSZhLICfwuiTSM2I09L3Bcud
jsr1e6mtBc846Yp/16vWBBvSvZfeNuWV1YdT8eXi3IRq579c15qFA+nOKLKRFry8
aFeTS/5Ag8lZEi2bCLGMRku6FClKgOW23D4w8jQPc9soZfDIiRf3yEUH/OYr+SEn
kZjD1mwsCFQiRjhDMza8uCK8sReej7SamXSw/dS9K/gAWrQjl7Ivq6tGee9ii1cm
ehifQm5oQRy/AQ2jqQlDpHKZdXYRtQ/A8NL2WZIWxE+DF5ccgWWELXJZ/AWesShk
3JkW+wmhs/HPb+G1E6NI7OuI7OieUW5CUOJ2QfzA3faKxWd5vZSGgTbK6/C8duNt
ePWq5tX80O0tCYbeG+x3goV/f6t3h4GSLORtb3roBy+XXfti+5lld9qzR5KwwpQ4
lSEJWaK2SnElu6JjvJ5ZcCs/sxv7/roS/M19fQtXieCcDpJGqdvMTo7um7ks6yPk
DhNNeu7mIAL9UwwgjOEfOOhSc3JkfnNYlDCfacAdM1JvNnmvgmVNse10GnY6DGSb
W/tSp36apFpsk2qF1BtOobHM7nYMUM+XpAogOSLhmaf8dTXP9Ff+zQrpUQa87A8l
K+HaWihY26Ixw5rio1s6n+kifvxCh+hlhsmcvmzYOSo2hfynH4iy4SLDdcusBGkv
GO6A4ic4tZb/01ojAmkPAWowLWO0i8/2PqFdCdNr31vihmGcsdK8UwasRYKJ3ebX
eOZf0ltDi0LyiUhGRp91N9OQUFk9eTDf4sBgon59hJbxpkwjvWTryLaG6A9Eac+U
5dTO5+MTeNI494BqxOX6fOyXRKfGB3KJy+yF/EILvzsSbReF+mBXCZKCv+dvi7hR
HwpvP/cE9JOv4s477PN08AUwdC/4C7EZOdyJtq8JbQLhDK3VBhz7g6+Ei2n5GuEI
V95soJX0NwaaELwD3OOBC2TqXlVP6SqXqEEtHz3I+InXkCn+a9Dl+2a/YQQhnvCz
ZozWbIL5fBxtc7UsAkU4R8xUPTa4qXmKP+jzNKE/CtlONRFZuu/bkkoxWmb65MwQ
434/vFzhF9ouSy9Dk4LjUnM1UoYNixaAOg8Ity82JBqMmzR2zP4aXcwhFqdkGQu1
fY+YPniJj3RK86VRfMTtHJlRikvCzccyOrlshUoZCpUFGdEUekIlV6HDlYmtop2q
1POYuBXZbnDplyFBxtiEjMGaWcp7ZLjOYgJNmLHeXEsdMVXi0pzgo8k27KiJvDZ6
5VlyexlDx9Bul0NwbrJbUw2E696ylIJK+u4n6C/ajiIZKQvT9w0GHae2N6C7w2zD
3r6TmOzyPJLOqhTluCdxZXJYAFRq9f8Q6sd4OujlHuXkVI/QB43Xe1o77/3Dx9uX
q0Fqb43LnkX6LU1YKVSE+Lfj7ga6pKuuC8fWqK8pvGXE1PLie/GK8mnLaWt0YaDL
dpiisIYEHytbHmFSK/aaKdT146u+/u0AzXdfIsBLYyQYuXSSv826/pbQgrsoM0vw
TI1q5DLwFQw3x6OKDqkS+id5ZZjzGuPsyEZnVWZTQ94NCFw7zHM3YQThe4eyemW6
+skm/03o0uINrEwwh3ruSUDfCl+jyd2qT7vAaYVgkUfXCuBHTgtmfVQD06z5dUvG
c3dweaLI926cDBhg6i8/f2lFO+OHB5PqGrp77pqJjF8Q+/WX8bYkL0ubWEGR7A9p
6W5Frpj0EhwI0fUgv9eL0HQNsK+niuOskB2XB3/4uPlx930v49XGjddB/BCs43Eh
HCLaPfENbQfoKPKztftVz0bSR6kGjv2RY64VcLa7CeduHKS5L3ldmsXjKubsS3X9
sqIiB4KYEbHFgMcnJC0WNJsAEknHKzFVFWDGjOk0gf+C51tHggBCyU7fs7MnQltY
U594Mdhh4VHkk4Z0f/+FMtcY66uM4qA/nldCJQmKR2onZuaxRWhPxR2FSXvo8LYO
jdkQaKujS8xdFor0Ik+y3ZxJ5rYeD4JiRuFOLdFqDcYwZtX2+EYHyiKkxiRgZ3GB
NJ53a//0yJrC1cf7OJkQe5/uPgRxXkm5y+dbacjpHLnDlk/e7KgbsfJSgg725t7M
50B5xFK8IVD/BhTMJR52Akle42hw9Xze4iZeklCha+pmjoikxHUjtlODz5aCjmr6
WoXTxYOehKC/FKAluot/ePvDKWNTCZAnhR2+dRXyUCds35T3ByjTkqnGAsVzEK2Z
i+Er6R8dj48qo3ILvZODapbhuHVdXptm6/Rpx39jRMPXiNTfujUKZ/DYLXcen308
JzpL2/Q5iYj0/dKi2dLocF+YTrfCClss8nEe2npWogfzXG1spgdUC3qF0VmYPaBM
tQD4YXH3K/TxUseeO64qWgJgiSPIUBQchy6B32OS14vwtYR70fR3Q99PO5EYn/9G
27Wfi0jCFbTCHzFbLavQJVbcTWbfFnusGnXFd4SlhritjMVDJjCBeA/fqyrG0zjp
JXimkfnn4l+EjRmA9GddbKo/dUkt90B8YUkBvv2vgTNSWo6OL9Ns9ORKJNrB2dfO
8n0VdbGuUuea2RgEYu7ePmbFnRoVlMZ3GfqQzLdPPQH8NUkncnjG8CCjEh+Z2G/7
Zs09+i2JrIUiIfdjlvoouBTP9wVGB2fvfNaZYIfIHX23CZhUNhjeCHSrpQeOch7u
dihCaSlMdtLcC2SvmVOAb01x3BBzVEVAIt8geJZBBaX9O1oLlbGPg2hu4B5Jts2y
EwwdDgZGMqM2PHiY53UYFW8d5MCdlOjlr81aN9JH7K5wHj1SkTeUYEtSGFSuAr3O
M58NU7rhR9KOZ5StTyqrvu/YZ59CdyjKv1yuspvJPbD57uotM59qAEcpofqn0wct
oGGSGA54az9NGM8XlD2xyiR2/y8RXnop8vknxXztIAB0OdboN/6J4tIy0DB4nelP
5w/JXtL2eOqt+yQOJ0Ire1IVBXTx/XbWB1TpJxe82IRro3eGg5bqCJtvs3YIMVy+
s5Twbp/FKpNLYDKpJRn2CX8OPqHbsmiT4wvNInFU1HPVWavRmNqT4JvSDbTZcNq7
TIGaueujH3j0HVkvqWIt4pjHle/cmIQh5jWEsZK5cuRAoZPG7lW6OYHsze0I/dve
fgJWMAr67MxNJipB0nsWExRfztwQSd5CsyMmDkPkvDa7Q9jIMrfUu+6T7ZNtx8F5
I4oSM/H/34o+wGuAt8DXWREBLJif5Xam9eBIWvjIugLGjs1LvGcNHWRfmcPcHyNG
CxVZrMqmoKnSeS6FuN0FQ4H6f2LAoSy5ylVjJ6bQ3hyTT+MrWCd358DMXt4V4qfB
0PRJTWUiqShPp+u6EEP+9/7arVYLAnrhaXogxINGD/f+Jy4ntUBFHgj1vpTY5IpE
ikmjKgNNtHldW4JV0QvmA/xGJP84iPmYQrJjWYy/kQKKYRRRBFoZXKnpM+xLoWIu
xYTgaFq8JXR1TJURPF3H+uetS7Gcfyk3RtPvuCb0IW1/OoDrOhXxOIlMENtdGyK0
vyRsK+y+dVD1rZLWL17234psu5+mMNYSIyJLPACfew9lNqgtNd5TBO8GJkUWRj52
2GjPGAG4XgLp/msjp/+qzfmSjmopxaKNA+jfAhDons0+8YlmoTLEEMjrOFUaHLy4
dFrWPnUiSKdqlJ93luepqJQWVPLKH824EpiS/IunrfNjUcoi2aZ9JgmRSqAolxIP
pze+QDUFHdzpmJMxLijjGDgdptGqNN5L8+SAYOXvhO3/fT4b1eHvHQskiB51TbhP
NrFjEc4cXH2LTqoxDXTvQWE6Hat+aiqm2uclDTRK1KOmUVrGZuoPTvJycP0udRAt
RADVpaFn0K/pqTDBVfZHC/oJLG3L5rkxOSwFCWIuYbxKFqc6dGO0pBW3HpDFDFDd
SPv4OfU0yRE3FTuc+55kdrhcO2PT+7/V3G7Gh8QrRz7MmdmMkibMuNjrpEJPir/b
lnF1RG+303Fo8+UL7LvP7y87NVfilgdlA2wkWbFIAwRHFTdQg/GzRnzmIulTeNZQ
BVBEuL6Dia86FuMsgzt9OYO31aTi5H6aeCbH8+g/M4w8Gt1Vi7DSAV96itDtvuf8
9k+Enw7hTsnvwVT1DfROVHRCTVqiCrxZAx+ia9moZbAhfERsLKfuk29T7J2+T850
/JmkP+1/7keZ9biBc50QWoNSYZGdpRLpu0GGKD9omwHYefE8r608dUMkhKMU4xB5
3X9L9fD6XvllxIW4ADutzaVPq4uDydeRSm8pmkuL1PKTwsUzcwMdALwurddN0DEQ
LqQjrDTJwk8zXg/zjLBxjJP0q8lHXnve+8ix3PKm3rfALcqgr2526rekd/XbNUSU
WP1kYQfT4GXdZj0RqO9SJpDZzOYbKY7+CnWeO6Eqb0p4lVgEyljF7cLoR+6L4Vv2
+cOuy9N1aM88XGkq2iRTpi8vpV96YQfBg98OW4KotA3mqJOuFTZLaLWCESX0td3D
hh49OiK4tRtcOzjJ8iuEhHLjKKEh4MMRL+KZqxa2xQUpgp/ERp8q/YEKg+hPHjf0
IV6a2m3yv6oNSqA1hbzhLW68Qh1cF777a5Vq5toj9JvZvb7rOSJW6pdddQwS5E73
5t6LUc2UBU6oqcqx+YgWJ1KA2ysVUbWCugA6eN4K6lCvKbvJKrG8QEIA1fX/g4aA
tomsWSaMMmzl68wbWXuvPcmHnirbwe3ahnND/pmjsE+FGI7SP7UQBPNKPXMbD4Tt
WCuKiADpKc0FASJPRV3qu4Eq1F42MBP34QfUWCGrdW7drXkVoyO10jVyExGCoEBb
hPiSpb3GMbMX0G/N0YmoEnw+/a6V2LlUWVzlMLAKG5NV3hfqc6zC28NhsaKVeHTg
+lrEtF+vVdWOvBgElW8OeKNJlfzmiuMWDj9Ct+cdbG71+pSc0wOqJrJQzjzpBQ61
RieVA12teueSbAhG8nVqHESjLPgCWUO77iu0NUCMXMS8xM/rrsbXtK2avE93vBb+
UhKZZoJ3SLQMlPF8nCqD5EKYLZtMXzrDnQ6A3ztbCUA+el9tzjlJJIaaMCGMXvIc
HiPkvCv6UyTk7b/WT2SaGeFN2uW1B+JOmpkx+x/llBmcCyb1jVTUeCeobBVw80Fg
xddz51JN7OpV4Tn18MXIFnKbQ5ANyQey5NzJZ1pCkaNzPLI/kgV/NCVru0eNW8jd
xc4nQb8E8mPuau/ZSlCXY8qnvk2/kQm0JjSlZ9ozveVr8PePxm/I5HTw4lBle1of
0qOo0sATd1C+UnvhIXSH+55w8FO4v8RtGmeAZdAZ9nIUi/zeioM+Nn5PIgRIJTOY
eQWGojHobVQQENL3sDRYoHSTfh2ee/JLbEGW3W6RnimFtenZbwPoWlF7ybCt17zC
ks0ujhJ6MuxOPFjQB4+Ng9gmE02Qro0CVpzDJmWknmzwpo4qDFy6L0A1uFsUk1kr
OGX5Xjf2nH3WNPWzf47uW4P2stqHvlPxRe68GTEsjRPlSw7VcDjVLXJp9GoAVpbI
e1R7IQcP0QAfdVH4YKVoqtDJGnVg+JCFFGt5U2eww6JDHzxqtvg8AEVn5lngADej
x54gO8NuauZZNJ1dl/L6vtKS5jKpPNTjDi3i8Dr7sx9CaC932w2sZARrYJtUD5gi
lEkdMrc+ewcpe3QUk8qs3neyFsfFEiixOrTRqIfoT4bpIrox2v3HS43d4C8VpNm/
dBAzqe4KJlxjLK1hPP4kTlQEo5nDS6jAFRDJqUn+q9JiZ7eHVVV+jynZJpjigSrR
F2Fjxcty/00NFldcNgvbEtPthl4Rt5QOj0iqlMrSqxAzMUmrUSbmNtHQ3eDJhxkL
d72vzEZPedCCb/bXiljNcvAgnLv69z0yi4V3UHMVcmIyV//y6HWP9GEkfqkJPRiW
1qV5c95QhJ5JE3aA8a8xsYOiT8dVFcYAu0/B/zJF1ppMzx++bKfCZMAPmv5ClAAE
lssIhopIK7L+EbgkmTTffUXL15kygdJ1Toy+X1IbT9G4xGTq1SNeLVsG9nj2nqVj
Sd3k+U6/NtmIlOWSBHRvrSBjtpmjvH0cNdWyenIwrit0tuejwxGHLAl5NgKyrD/d
aYjcsTmbBbqlfV1zzUkX1CR5JWzU+5G11LfLsqUTDbg+HAQRykNtk9HAORLqahPq
TnDkCls2WICVLZ9HrysMtCoO3ldQWK3/vFZU+7//nWao5L9Lz7yB2tH2VGd9ymsT
/bLvAS6Q/zzhvznp047e0ZeIBUJe6kUdV76Ao84Xd0jl6EwPQYQ8YG2te7eDyISj
kp1Ez1Sv6XHLYabMJ7M6LazG63XWEloaU6noXL9fRDpkVHZ/nmv5tMvJADhjQnjm
wXguv2X+P2QBUmFXN4Fuj4MmHv7isVkUDHLDFcP2mzRTAMcwrPGT5Bogrh8xIeML
5xlxc/4O4+RHvimCSYCnHs+kYbILDFkcSqNmS4qIWzTFT5jF2NvHbzF7y7SrzjCy
8ltIO/QNyuTtSE0SqAgfm2ze6q3SaYd9uVnn5fM/AJGKPrIcwyLAFJblK3tH2ENQ
mvs7+ZxtNuwKGe6ZjTKCY7WXoQKAQDWOXk5kIaCEMMy6I4eG87xVzO10w8LXkjcE
yJjC8QC8NEdZ4LJWsYuY+sxgShhZqdXmXeB8Qv1/VpRtqUCgKgucx1ISo9CAZzXf
qR5xNaYI6vnrPRyGmAKj332mSugDCYUfp51+QWUSoVOArBG+wuCtcnKQdtPwPCuR
EQcAm18VgRp6rqo2Io/qSXxT/h7uu5Xqu1trXFrB11i97uUzi93Yq3eRkGbeq/tu
kjie7nhLaHpgaPazYU4bvQeInX/xchut54m5SBFRrpmVkGiBot9L6UUKfGxEpmIY
UvpJCHfYd7cVK5RmlpjhI02sk1rT4D3hAN8oAlNu5dK7DdoeJN+QAGa2rawf/8/n
6m79UFDXPrP17VQfhWelBDT8/lizP/jx2ebl/sPaW9akmzqlQH5oTyV0o4Sgy9OC
/1Ma5kEimngVUuTUzNBT1YSHij+/X3S7ZWCBtKoItjtGHIe3v2toEIj/guxH14a7
qvPLjanxHqx76jF/SclxkrmUjo/yuE+gFFdKVjOdi/qZlTbXcQfpJUYLCZJAba7p
yazQ0JMph3oXmdH10FdK6FfaDMxCuKlRQ4OeYkFvO+ewMlba3P03iSZgnwTvmY1b
JLWRo746H5JmMrrkQeAeRKCxhQ0mOz9O/k5SCmZ1OqSt2JruZE7QuTGXsgcQUteG
AnL7H/kifevsbXnbluLyTK/yxf7hLpxCu1kd8lls8aUTsEKIYGV1a7tf6h+vEE2Z
ucs1uUNsQIHw/74LoTLbqe2+F/ARBE/Ilqod/MuQbFnEKc/MG0cAAFnAV0P/IIn1
xaJJpSVyDe/95MyuKh8EE5VhCSShHaP7ZX/RU6xhs2ItOCMuBAcOmodTrCpL6nyW
2YI992mFq590gI5FPw2IpoMkCSQqFoSy48krAcCa/i/KNsmSXHQk9HENDdhk2Myw
SjynE6aozFQKpvxrF9Dr3ZR1sgK1i//9viRjJJU7/v5TXqeY9Jsxn5pmdB9Z0qrm
3hLA/s4r9k2Uxf+IwoEEpmuq+gxtY96h1fiDsdFXP1RzZXk93oh+0i2CvOixXUpz
EsjGQoimD+qmfBYalxqmccD6V4TsokEMmq4fEU6LiJZQ6uGOb6TFPdrXHvE+hi4f
b/ejczkmZ9xPAioi/DwhQIImfjGywClEV9pKYAh3G5HrUIolTNoMtt9BZ7gBAaY+
6M6Io+j+1b1qSF6Fs07JbUll9elODGU1Az870uHue+j8fMqpOa6blsNyYGelV9Gh
+VTizVPU9YOlm7N+8rKxEiUB8xKmCVpIJ8UyFzCvkdbCl+YVFrgM9RZ5KdchEe+Q
0UtVz1mdgEX6KKRsYbj6IU9cqur54pIfhX/YSyDS+spFTZgqQMAPMKqw+kthR6X/
scOAApJzeiT6/9UuUyfh6WlOHVs90SYfoww7ss9zBGUVcOC1wRtdMqu7PMpTnJCl
s/ENGgvwJljwOrh319FN1IksvsPc0tI5I3JPKXetTCmMSnijiEf+JEBFX8KaZUMu
IjA2D6a0q52YNvcKeWmnqC5euAGdqL5Eh/iYErsfWmUZxWPsFhWWxPawpgv2yYqm
W4S71dGv0qUaWBg7M1ppyhRIg4SG+D4LoBL7bV96brHZsaKBRo+SdKrGQcRKU4tZ
nSBr+jfqRIhA8j6h/Ya2RrfFEnWegISF4QlBkh53QYPQQdiP/VILxAv9ti0mOuuP
x/mtsrZGo2TYBeVLIjhvLKMzfEeTXb/HcMxh7F+YLzpNr+WYC0CNh79Nogto6Vhy
+2VWrW6hzIq5Ur3yC3eaAccxffzpqm2O8ztMvkbJV+UNHB7VpcAMK/lJwcIzlD9g
O+MWlbvStEyMAqXyC3I2LUWaDyc/UnVmfvFQW8CDmKXqwum0ce4n8hO7ZuO9Dez7
TvvaYs9cMYsx8sO1qokoesqn8WKmpfeXhn598GMgSTbvfAJGfBH8wakBa+r+6Yav
84PngLvYyrmR+otMHPX3427dSER0EYyEpH/88WYQiw7k3O6kjebWPB6Opsc0uTT7
ot2Vu35fiEuNFuym/RvYp/YLVVyZLs+8LJUE91gY34L3Ojen61mC92nj1O/7pzD8
W8yaZfu2PK73c1HvjWflUydK+brTgIQ+eNcBCqVWBcDOMpmh77rNda0hoCeHXTLM
qsZbdEMvTG4EMJAlX4tFUr7WBfmok+mqb/gKo0PV5Evs2aad+9rrKN5nrdUJjla+
FuozDh7L01Tm6SwCAmQ1k/ZcEE92NNwCVH6QLmJHUUz5sy4hjDJJ91CC3eGdY0lB
a0TaNaUkYkco5H4TIExbR9ZRhHNUJt4m3M7Srbu5NMrOmX2DHJJeNmRxfxk9/JWM
B4/5KIkrcUBL8zfl1VUMhZgfAznnQ6IjMaKg1LynLmB2vyYFlUVMRU0jT4Gj+due
IF2Bjb+efdUuaAw45qL5XsT3B0egghgW0rAe0yfurBQannbabU/iPzY4kgSqHEqI
5mgIgqzK1JVUwd7t9/80d+3JDaGOoVVeZPcgvPnqe2NRMyOU8m7qHEuVomZpOvjc
M6mstfyTw0NP+C2Y+8PrFcDdFE9glJJLEP2bfO+KFQfkXQ0LPzugXNT2kNILDs/B
mw4DF+jwR9ploKABNE3iwVZLYe9LqLlzxrfXvBTrxRIT8zvRxLvR4mKjIr2WJeZT
FRDt3LS8doTd1tkOcKhno/kyF1ijMvcxhNVQvp9yJvZk7sAHSwqUned24mVkAt7A
+A2MYFBO3TLpoQgysuJF74TZ+rr4ZyZ79RYm9PoK/MkeOEbdaf9pU+GRH1PG2k6Y
zUiFva2vzCHtjLCrF5j+AuI6CeaUUYgmkbNe9Qo1eETYIsqsh4zVM88fn1/dcQ9r
sLDLMTwxVffZNQTiQCZ2KPvGeV2ktlWPxpgX5k6+0vNiqy4FA1joAzKgE4LT8mV7
BJApHwfJpPicIGvysuqWmb2ri0Wlcmgy7ByOT3pJKWkeJw46qxkYG1nzIKFlDUnH
0kiL52ZtVYNv/165cLimiWg+RYNmfF3mY4+D9q2GD0drHhdCAKtwZJ/gsJ9lqU1M
snCjBXGtgo2FfM8n7t2bNJhzd5KxrY4KXLPaHYMLqIyNeGOqFF84Nfc8iFhuPpSG
VSuxB/tRfxuqG3hh0d7f3bMAmPGagVI2ZrPMUyoixgX1SOxTLjF/4a9Hm9er2B6a
l2xJoIH6mnmHoslKLqsMnf+hgocjWBxwff3DhJUe2Eg8M5/2GjtF/HPVRACkg3Zg
htLMybrByG2qSSYnr9G3hO47nzPVwIGygFaB5pf9gclnsniR7DKEx40ord3XbtiN
JilUoXbr4Oqib8+s0qXpZwIJBswZkLPwLq+j8ct7iVGfK/8JIpevx6PLjCuqpHdJ
mcXOnQxn2hpXH7it8tWIwCBp2x/qkQlJTkEYLeltjwQfV+a+RFIk65GqvcQIlf68
aCru5JxsBehD8Hnt+InsSSuuP6GOxf17034nyLmCym/WdcW6mhPZGQ58tjp2x3P/
axBVHYz/nJ1VPx/WKHXiyffrMheW3DtTOYBKMkEJE/dPWONtekppn1zUeRE2pD11
POjR+Oqr1si6KmVWElB90yJEcH6y6UWoqM3QGJ8NLLCg9NzuvIWuuaDSh/nmadDm
7CoJ/Ct5L/HOMuyUB4Rr8+1ERDw5JHWp9+/NHSFspT968TfLkXowgbJhlPsWvOAb
636binkCLh4AfAXPbSuKuaMZcHJ/CBp46JDOTtKZtwPiAm7CGUK1yxLWQrC6nC68
ojRzei6m/Hfy56gsr7zYPFyAY4Qd1evCTHPLlKm8CXsVWGHHFVL4fmu8L2uuxOEo
jEA3C2EUIiVHuPAnxzKMU0dWosqqziCXUmcRO6Bcv70aoxXoONFsOZz+5Ux3ZKwb
w3MDs6rbjO5X7srD8TQgpfiGhDWvCSVTrxgFDS/xTumXWeRoHNb1835kVQDCA46T
0oQWkySacyi4rzsR9YFfcho4vBzM+Frma+EOc/IVzoUc5/cpwhkJeVBcggAdHcpN
nU4pHgBIiyv7m1MvtAQWPrwfZkTnUDkjlyyRxrqzDSUXACcd7Gz2ws6pVKNoVWFJ
u4qKHUcdk2xrQT7qPFRq+XvdM5byo5tn3iIzYuHtKubUN0HK4t/R/2e9S0oLMVyz
PN1l4167A2vjcfeeLJbr5zfX5ElnfD7QkxHJyVIyKQyW5pHWnEjQD/waXFvrPp37
d3w1ndPsA8VMntLarFrEriqjPpy4Rak7QChtifNLMKinDyXLx+chBSCpD4VQyVqJ
Vg8XqOwh8wI2jaR73oLpgvxySMNu8/grSEP+nNcwSpZkQCQCEAo6FNE7lq4QzxBT
OyuCXlPQz6rBbr+okXdE3l1hKDchQjZIWZ4HdhM52tFIGOYp5OfuKhUzweCDH2M7
2NziGodDaYzSnAVMiZNczxV3QL9EdNYnaaapRtBY//H+hao1g+0tu+Kf+NIIwoDI
WPkRpUu4AzM7+xKoLTiKwWvu9JuX6FFORnEhpcneCo6J9kmYdxYayfoNpiwtVteh
ycBpDYBrlbfUfNsW59UU6wNONiOrNdPbDyr8sGrqjMLcFEBFiwxlSSdEOwnEkuL3
/+2fswRbfLsfvLyQDBWOv/uOQYyHTC60eA8aPgIQDxXgxS2teWccTjiJBx9L/0ix
sSSglCgU/Ipt5QKmsWJM71+qPwTKJ6S+1lTecZ3GcZVQXUhM1oXJ5UepfHyE6ZwR
qLdD/GiUj6Kqm6ifI5+g6mVttKBQFVewTieVr8u/w0MvTOydWmWod5iZ49Cwj97v
SdDz9E9n/GVWoKtLgdnzlymkr162JXbwRlKu6pxCqZHkHmleAKo50Y0R2ulpFSWs
UzsYMbob3Rb+ypZNUOXiNubp9bjZZv82xb0/dWxEZtLhjGp4li5cBKxXyWfaxDGN
Xzs5pL6eaEWfqDJ0jKDYs5z3flKLzzq1NsucO36g3iEmYd6ncoqrT7I5RB3UmTAP
h3Ybxz8iz9lOH+pb5sgNNWIPF6pjF37dUKQuGtWS1RubRFZXGmFNuWo7x4owBqSd
ktn4k6yJ9SXyORqmgwsQ0ZNPWGu2lGFcW9YHdnMuK8v/cRP6EHOf0BvV6GD3p5wr
S4R8qq/GAnZhh9N6CL8OA6TMVmA24HjnhD/GKqTuMR5aKsei4sDL3+sGkEgr4r9j
/Qjen+/joH9xM2QGjhG2Xufw62hubbrwMs+sSMlIFqQ3LkdSlqp4G/OseYGeqNNR
QxVaMtVpYD3fCoBSjQ1Mc8rOt8NVv4yZPtj3N8grMcNVVft7bA8rfAeDB7BEMlI3
z6Jf6y3JR/Ipq3+1eBf86Of+ka9VRC9ObNd0LnEPJz/6vHqCPWjRBnLAE4K6keyz
EiHG9wRxVYjioY5DQSrp/r77nA2O62iZSkH9x4jMrwykP0nx8yMt/T93sNw3UxDs
05t9JcBHHjHfm7n/kaiZPU+y9BaQKOCA7Krux0/WptNrtyno3h/d9Gf5I+vAMlQX
hJe9oeCyfB0+b9FuHVuwFiBlRn7GY68iu/M1iPlHl3ZOoFInh9hdYAXxLP6/cQS2
4BLvCyFjZ3vRDvo0sNfM7TnIOEG5jeWOrbmH3kn7apolg1Fa2jRJbqQawwxU19PN
nVlMwm92j0FKIgsagCRRBhrF4ofJl+PykTKof0g99DWrWFoVf3UWUqABpkcSG2qN
NsZedDcOKdKwKanzqXMVoFK/d6MW6pD6gsgydA0mE3JkTis5T1PJwxjyiwDz+6pv
z8Y45pp/ctTTVyblf0kloaJZodsp2s2U9MKVbcO1MS8GA6Kx+TxTWdrnjry1u2+4
ZO61h5jOXJd4mcyuHIMpkkW+bOb78gNa1X/T34TOMBv3MiC8HI2B7zg7fjzN2D0k
7ymgT1g/pFbqsLn8u/voyLHUCiry81g2VcYV/U+IMvCLPnLpSrTtAHzrJY7FdwMn
j/xrzm/pd6Jcs3ex5e5ZaUxoK/t7ujWwWP91hy1nBYX/nxS+CsyjegYET5HEkJUr
jWri7giJoYUUm9078J+X4f6P6f8nrHFAqKSo3IPnTVAiB9VqavVW2Toach3OzdTw
odPyUBhmc97iFgbd2wrOGcWOBHdURK39/ZJAdlx6r44Bu22/MS55EEPNPJ+CNue5
jVMI319AiubjQ9lESk7oEz257DsJ+n5gzHnlSDRJB048S6r/96f7mfPakxs+ynBX
xkzyDjHDnqPHn4DXAX3/uRvlIrBw1VShBPqb0jeS5T4X64Lcsq9oFSbOTBLs5MiG
I4pfg4y7W1c+zTEpIvw0cLuWRWvKGEIqQLynM/qqyuXtZQQTnVdv4GMkxUFciY3z
82a1KMojnjcVTpkwn5UhnBE+c3prPz3wa8QlZB57D8yFE+FyHwQmmR6AJ2QGaHMv
0ljy3no+ohbIR+A+yDOqFd7lydOmgc84wHJ/FqRE/IOQij00ioJtrh7/s6tHEHBD
LjXoECRjB3Nt6BKZ2QjckYBBXgGGDS66ryUFXL4SMf+JZJVgJa25OoIjN7fwHaTn
3Tfdw4OxScqPE+V77ozj5IQfCV5JJLZolyW2I+rsDh02cP8RbgCOFiBhqUNcct+h
36Pay4ihfm7eVoFFi7UhCkQNcqS9KSnlYRADdExDDwRV3ocm1753AtGJrqMuFNTS
i02VB5f/XpUHModketToTX9DhCEdzadThgGB9njsgJ9WY44J/wEmKvPp+/RQE5+p
tBlg7sbFcnQT9N1bct/aBM9QfBPYUABCW78XXJXfL/yozRJp/shvR48YMwySOov6
1snvpJdDToa9gXVQNwZqR3syWUvCa/6vXo2sIieHMDO8PG6oWeMyZ9CFKhQrCJFC
U8J9uv8tBOXzWQ/hzj3zY0z01EsczVIMySDPpe4dB/6fviedS8Bfpo0X5ewQZe36
41NEEb9JLIJoCaO4UGYxcsLkQkMtMgb4N2GIo+aUqROTG988neVG85vMhyrpwEzW
sdB/D9myEhb0bv5Qv/5JbiJ/AW/SnpH7CXWPDSr05X7QU66orV+earjprswcrUUi
g8zod9LCF/X+UuoHaITLjzbyd6zVJbZDP24P9QdLeqoDJVJv3Zx62mcPqozcDPH5
LU3QulCfmoqNWdDzCyri/KlY2kJUhk6zDBGTbc2YVyqXNGHo7saGzxXLjsCLpQuI
KvRORocjVp7wch8NipNgb0qNyaQvAlBoLCw2m2hgi01g6KR/7nHJtpsj3LDj4rRh
dk2PmvyWr1ZCoOECUXuRcVSak/+67v9BbgsSLPG5OMArRlWATv2IhZXNK7tXRAKv
fqhytHc8OTJazyQ4y+X2ZgggBK8xed44IIiXKxy1NSpuK7tB6Q8C5B6rsQhmaNc8
1EmcaI3ZwbjzrA2OmOtxX9l4yNx3BgjuhJ131zOwpIiKwKmf4Mm5ptuG4bo+k3WN
VVE1YvDqQF9i9oC/7poJ3FtkZ+GqWHTO1ZjBCyoNV7GVHOCajl/0gO7NPAU/CpU5
J6zdnn1KkFPCQo9GtvusEhThxUZ85uEYA9xu7b3fQ9lyiSieabyYV3l9PkzjqEhL
9GiwjCWf0gKxPWRG9IMn03PHCWQ7Oty+tuTyPEW1OmBhA9LWM+z7x3k0DTUQgyrx
s6bVVU7AVI8cZYX72vZ0+nBFBxXwrO5T9wwt2F3i5pHVY1awI4nowS8heKOTY54P
GQFbldyxRd17gr5rpr412uOhIcNhvPwqkyn0POtO9qIViYxj2CPNfEf3479ORcg2
XpzPC+alKZRqsJg9JpnHd18Xba4tCf6N9C2EG+locefZVagn6z7T0f7hGTpsX34A
lyxnteZsSG3Yu3yqHpQbF+epWXdaIkC3h7vL+v+aZCK6yJ7l9O+ha3LgwF+L1kKy
l1b57PZWo9r6+QgNH2gDwWEtwa1AOtcARYrDowWSmzVkWoi1N6jUkPACDdtRqcPf
R+DZbM/wz1qFGzdxrPMypbsuG0hwwRcCDLWvgHfZye1Hg1H0CXCcvzghudEtw7Mu
qB/j7PGwTMLA8LePvp6qoW+0vkkUl4nqvBXIwRNzf/GedjTnaCuld4tqZTov2+St
Kqh3rU0J3haPSzTDcDlCLXnrNsI7YSP02Rg0CARMbTvtJX3ABCRDsg5gWxDRkQsq
otWNniwRMl5N/5C7PUT+aP4XtQ9weVBl/EjMqrvg/xMzzfDIdM0cZYayZ5/c+L17
LmRpuEgt7/qUGOzR2/srI9vSPiqXNi7C1tgBhuqWJdXBbNbfQrdW+ZGuMnyTxxnZ
5HWp2Z1ETThxpknwMPaBIyFoBUYjGpZs4s/kK39e49mJB/9KwnGSES97NNyp7BP6
pu6EfnRNIh/3xvczEFORN+qSQ24WKoYwFstZ2yQUevIdqpQuE83mtl8d2P7ZOdDh
VFyxVR7WL09Oqv6C/gh/qtgnXwBrtRmDpgQnM1CMWKRFWYrDYgawAqzfiGopWANc
2N7lEhTdSF1Oqf5Y+uRqydO9/xBikNjLZcjMGEbi0sUB2F2snRRKnIz6hcHVQF/O
tqnUlflx/UUW0sdRxx1ciHdZe/WFXU2ryHnR9QGRI63MfN3HTMiFQ/9laCB4C9G8
BwEKHmsVzmMdcFXXIO4RGMnvUjlOmISjMsRoxzCRNNYEOrou1Zhvehm682l45RNK
6mmKNVNU8RXfPvgezs5ADl0CW6iQFuUCdzsnHyiIK/9rDvDSHwJ9+BnuCJ2OkCUN
/g8rC5/XEpQ04BwkWd8ZFz09CvA9fwrC50EpbDyuXmIo2slXwZvBImKhF9FQ5C6a
G8rlQ6JUs9ZVPLKLTzk7HYQap0JK2JAb4YO5XETDa2oRlNoGwPtRMG139cvIMmOG
4HVF7/zVxF8+cN2MWOLLvKC0bLal9mssQFhx/jMDNSCDk7jP2lzhmYSde6CG5Abu
pWx3y+7G0au7JBb7nAjRj5GnzYOI/IfGJk+9hV4nuLpPI2WWbVlsF6ye+nhjBS/C
ULnm07/hnGcNoSchv6pz0s4dSMHIfjvcWlOBAE3Kmdw5puAQ6yI2N3ZSsm3ineCH
eG/Cez7bnUbHfrLWLja+elNkPsLVpjZLBe7mPw0kuTlntsrzY0yCPVEuJJGHj6fB
oQDXs3Y4ab7q1mMI22hTJglbAdxwYJEVVvCkGAzx96T5eELInfiGyWp0lnGWXU+V
qr2XXqgD7Or7g7QfTYdrQQwoNOIPA/lbCq/JEOaDfoqi8LUNGwLzBCbEeYS5++da
NON7eMlqRA2GDw+PDblGokby3x0mumQQFAHlQrhNGTjhHdYl0+CsMQHpd5YqdSc8
lCqoZ2uRpKBLmUiI/AHgoX4ve0IeVntKRasZu2XM9xOJFr14znWslArdm1T3cxJS
I2y/BOR5rYaTrWwFv5c7cZ+J+VZn1TQ5PnSuf2NGa2f5rIfcRTvDuyugwf64hLZ3
brcwg5buZFAWEbmmu4PosL7wqQHH2UQlZ9GMHT94FQ2VZA+6zhCYcDNI1zkCJ/oV
ZuS/IeavIV5+tRvy96EUCStJq9p/0waweNdTQrtdGlO71FvBRFQYfV8zcXSIOtlf
erpuB7O3l3ARgm9zyS1k2PwenJmXa/a9jSWvUBueR3SAbTyMyVVD2MwnAh7v/t6B
CSU8hY5IrVv8AlTUYCaRMJQ4gP7CyoMex0V8RGs04yoH8sOCu/aMXqQMhz0uq0C5
Q2rEwno6MwRnQtS87awmmhUTQHQR6XqtT7CAZwG+GdRFvo9MvcucC6voCpDLdpnV
HoG3QC795lXKmjfRKystx4+mPuTmK2L29vyil/dKS1guckbYZW4DAOy1lD31aMJJ
2LBhqiyIKIWssPD1F8fH9qgPiEq+pFjOUdlpNhmIV3jnpnCB4G2zYu2edtq9U+Bo
80JqPDqnYBNtNEYuScLou9VzlSNiMSlTuIiVwqniWUFzBtIyAkJQm9RVmO9oGgsq
nyw/3XGvTLNWti35Pb3XKRRmgwyEz4MQk7xXwyUMCiWnlkU6p51muqn1kvX8mdJD
cTT3CdTGJ2WMuQy8TFNkzhYIBkKQ5l2bQHbyMQVBgnl3Rijbmdaquy3cwDS/atC4
wWkQEb3CnfQXfvZgnc4TpMzKa3U8yNqFbEloLUnGF4NXt/b2DGzCL1/oqSCaYqlO
I00RcUpZKDcgtjJZ2/aQTkyHKo3XZciYWGJllTsHIOfJk3DYjNUqU9Zx6RT923Be
DmPxoHDRj0Q0vxWSwCqdA61oIDe0EgRWG6rj2b3WSLysZgGK8ZQDUHwqqzUFVhhC
zudjY1c40mFIr1ifCbkKXD334KtqUDPZP1CerYYTu2a5Mh40hEco+4hlgp3GnPy8
YO9eui4BuJIJH+xgfZJ7Tx27+qbn3Gpyi95prGwxrxHvBX09Jx9ytAnjK6HWwfo4
k9DiO34r6If4bN/QjlSSwZyGHdzCk99EH2XIIdeysniUBZWNHaKPPBZN4J4CwNRA
DkQIoJdZczyHCE2NKvZHivcYbhnugs7JQxba3WCeqkuK/hTW2htgPLeCIrvBantw
XYVi/i9T95hbqEyWfFwXxZ9BoSv9K6gGaoLfHL0TGeBZimYHYMAt5S/y7qO9c91F
mQNZ8v3eNzB0o8QxHAI2w7EyvIQP8uWqrt6UWNvu4QnIsK7E+V9sA+6w19GoWjpV
AmK/ODwjRGzfIZHmLkVHPd4+1GIDfkPdkUaUH0spgZo0gf8nbum/EiWSmJ5NlhjL
yMAu9EclG6tMsknOGlswLtFxVu/BLLk7TwTQpDdDTFqKzV11OflZMF9eE8I5k7ie
NLuOJu7SzQhPrR1/w3RnczG02+x+zNGpo2YWUZyo8lE9dmM8ZjuyZcj+Lwisacrr
H3VGRobOoh5FjjD3yCi9i9HtgFY+pzeGnO0p994SJvKygzs5kNud4DZPU14zNVOX
MRudriILl+GQE+Dl0SsdhqDBNITy8mu95j/mMYvDQ+HQaKMaKWl6xc0wet5Af0BN
+XdI1HJQrc0WE3/xuRhKydXpKVbVBv5hmFQNBzHbn9cHsimqJ/Pwq2cuM1OXFGju
grz5aMGxbIZ6i33aF73CSZWhjFEo/JSjMNTyPit6Nhmxk/WLwM+abAy2v0uDfeVg
ZegUIEEo6cUgOvLXNGZAq2fQMl8LDwvy5ovGAZoBaQAJLcsF1jFNoNc+J3k7x7sZ
RnSQ5Dbl1vqYFIOK9gI3qcs2CnoiH2IQSsaZ2DyalJXWG+oX95EtRkneeNpmDPzd
WQZZJIbYSAyfTlUclWIO8DlBgC7sUbHtl0Ji5jCZcJzGsbTXYMqGICuHbfaHXcSM
Abmh5OBzjHm5SudGutOJFhcb4isiMA/BAkaNVmw3VKAATu6Hq1/orn7qjCu+SUdP
YPl4yHkoy/OPGuy1cUVjK7X7EkkQYTASf8h51IUzbuU13PaYvw2IkDXsL66H96En
VSl5ZJQgy9MxFujZYMqapaxH2Q9QK1MXbJYr2QLwQudgQInvPF0f9oqw3tf0Abf7
FQDUcPfkZX6rAhYtBtm/uzgwBfLQutp+VNG9J5cr/1+NIUgQYK7tJ4eIb8cdTENK
g4npfL7NQtgztl1x9dSQ8mPBtd9wweAsMoLJ409oTuvAa9UHEpeCkvZ9dzfROQpf
M3kWxjVEjqXty3bPggnyE2MHPXFhGPcmaB500NhAUcpzUrWwqONuP/brzn6RI2Bn
+8wzdG6iiEA8YdLlLR6OprF5xkmPvnpq3JQygchsCUpMGmbT1vS0BE60CL69cVr9
oqd0/ho8yqDCG5XIsEWKQzyYoEu/WCrEmExWbaPZQAUuysw2HhtZzoyP+wcD4XZg
KW0kEgNQQRG0+GIXNx8PrFdJbkprbjEjXq02idJx5LZOTbTI2Ob8Rq6M+tOzADgK
d6UPiu4B9H7LRgQIqGi9cYvL4mOuCZp7p+XBENa9lP7Sy44P8B+hLVw+cdyKtkVT
uSwntGSnzSZZDU31x1SbgFBUIzkEyCsoHTgimTmJ+wxHP6pYYm31B3MF1//hwaec
CXdjwqvzlEVTJKuTlcgmKtGxJn4hH4p8F2jGYG2pzI2yahMZU+VYgMS0JUeWvbuY
H8pLFczk4AhiUUvButSpyGT9iS4gZ5Brf3ZaX5MwY/WFPa+DqzRGv8JiaD3jNukl
tzZq9hmMP8l3qLdt4dRFbcD0bjWQ992eTfxYVfnIA816GcbDT2MlT/zhhl4bX8tb
crAZKHK+QyX9lK4lVUS6MzCe6Xxrod2AvyAsA6+7EORWQ4iBr+TKrjh8/rg1XIzb
gencJ+4UPZiBqcB0qws1PJD6gN1XFu2JA/k/kKzQJoYsc0LwtYV+fnn7K30cv38F
9rp4pxU9MVLQg9YMO+MUkbXlp4/67whDdxdMI2ovhcLOrIDMjuuSLgjdlxRz8T67
ioJdm29ZtthzgGvBBY8FlSCqpSO1Nrl0j3qTVmajb+uWaKIbEPvjRdoGh9cFxnIv
/GImuZyd8gBXZPhADXmu0tc3cg7YiNW8NpHlQy2ti2yEEkwGtoOl7RqXkBMykgH9
e9ot0b5DRgoGm4eo5mfS03of3v5hA1W3swqGgXjISioDjoiZW1plUGB20dqBd6co
3aWBnKm4W1XCTtdAFpYgM4jQU4oI0O9EUC+dWmYQNH8JGQ1UHSCwTs7XkaXFNuy4
jnJ0MCr5fJ9on4pMojTtol0PN7ZiyM8rs4GdLpfWW+Q7CJiFsWVgnMV1gwqZ/p1P
kWu8Wil2QXuJ+jdabXkVMeEETEiT8a2LfE95JLnL0B1ZhUJB1Bh0yuwhZ/30vGOq
VoEpsb66TKIFdWBo25zFs05/3tLys7eZpebZKnyt81i55mnyj+ARK4H5H3a9ZYfR
Etgd6ugrw2BupvmwPZNRvElko2qWM9IT8r154zcMFoMlWKFfmMMH4D+YbqszjkUp
yh4JaHz7XOdPsZ0o4lmU6LOyN2vvNsmTyp3Ea6PlJrM8PWh3H7dqPAD6ytptV6DS
kr2b9ykh+3jwpR/wSX3HTlMHZhc9ofHDvgES596KwyLQAqSfQoHLVWhEM3IileIf
ttBxa5mAa0EpVs01QzIx5DxV3Knf1+qPgr2vKw1tEBEO0u6SczhkM25sAwahaExd
/YneXZv/nHY8dpImstTBpIOgz9mHDBjBPx+dS8uV1ZVsBN2QXEm5fvMYU9lX/2NT
+6TeOorvawpd+K3h8Gf3xSm9s2mbcQfGaHBYZxcPqcHVjijC20ULYbg0bWxaVU2A
1AesCYPpMgyQ6wt1nTMGX4dyF/kvO5vkUO9mpo80oL5NcmSksVPNMIHSjkg6aJoO
lJtwEoCDyLuWcQrI9eEvelVxSnzq2o3XQMU33dSpBe5pDl1pPk4MjOQZkj036ndW
hWkA9Crf5oZuTKCWF+KiCkRqVQ0lBLKE4x7OeqQrAY9Xe5aWeTR5Q6seEmD7DBuV
RKdlnhWFWx9iCGEE3piPfDX5cNwwQDqkxoTW0Xi1RyESO/ln975icRoS/rmOt8Lg
+3jYZH5RVUPOCiHVHaS0+mVI3l4WluOmOKZiRXmhnWSQK5/zFu/z9VSnrpHHYVra
AlSrw5A+Rxzt2jsAhQgv0pPD38l5XZPN43oS0a1d4wvdsBwJeJw0Hwi0pWGfUEqS
maVLIeqABOWd8kXBk48fVlVq8D7LMCoSIekL8KZWFzWhEA1Wj3U/NN0QPKu2fl2K
t9vnsWM8142KeAT7q8WdDD+F9jwP7tXOUIPhEYCnIRVHA4z4fsBxWsykVSI8kWP9
rTk4KPi0ofhaNEvL/sdnwTczrLUHbp7cLN6/lDgXJRxx0i3ik4dHXQZcj/GXMdbc
1HNpIIYY/kVo9P816iKv6KkCB36l5MoKScO45OQlxb6lT5o8cWp7xDDWdzhX6wKj
h3AL0EhgvCKwJkVVeaYB3aMjLiizSAYUc+wj8ftWjcr2z1iUqVNSLiJJw3ryGXnZ
lvkn4zoAS+BZlvMtAXOridzJkMSfFhzUV2YpOWbxmi4GRL0uXDgawIxFekL3cUQB
ohQPV6+jJUTrM+tuZB2xjwS2fCNjUAHjLffBnsOwlfkp2Y15aQMTHUpBYhM+6Oo5
oxYaiW9/E3e9YyEGhQ/4BNagj9+UVzG+GC3ySYBnkdNJfhw0fMaRuqEx1Ibbi8iV
CGXTpioxV5fTWsrFZqy4Nm0ltLb4Yym8AXJ82mcwfbIJ6l730uC6syWPxViAAwPw
F7XuXwrA6+EgzW+p6DfoZuS224uNeZdWpIpX0cD6i6+LlyCX4KmnXgQlGTmV4lz6
vJIUdUuSFeGdqmgajBoA9w+mcSXl2h2XnaYdF67l0EgJuGPyQ4GE1VSDYk9xUFQD
BOJzA4m9mraRSuE3vCVkSU4NaQQHhBz8C4TKjFrwUK0SfXfe3rHb2DfDB7F0Dg2U
oV74PLi6iPu57/x1xF7dOqScykbtfe8WWMl64EKk2Xgxarv01/Dk9+rp62fz0ANm
3S1SD3V1P2OpXMdi36tY6Z29EvUoVRX01vvfOb7RMUh2iwPvWG3X7StGHOLjbCgE
YV9VZOQzZbPQCWogRxCXnMOQ+EZG1pIwDz6bAC0G1pIWlIAsWF4wgm/GL8+G8ncb
5YNK2aSv19NSwwA3AtX5buuUeQX8NKtg40LNRW6+k6/SFHtUm4Qv7k2ZNjqeia9r
we8TpFloL3fZ3HSA3m9BXqkiGPhZtSDlwqbK8JuNnbZvRMIXaAD8EscRWBJ/Swxh
SwhxvjddipWmPyjTyMPgaB0wPX8xfh29QZDDY0R9aeU1CnbTUrJmP8Zo/Rld/dgz
hZpIagXszKwUSx7yW5VmN2oLqqe7r7w+ZGSWZpfw07XrD6Kn0B9z8oYp1q15McJ9
EGu97tZOlKRiVWMDW8LTmpxSkDNDq8SLDrsUMz4R/62cV5ycx9w0LYB/M6glfEKj
QhT7EMJ2Q83OaIs6S77vYpMRC7r4Rk4bP6fRJRu90/8F+TYZtGuGEW2FRl8ErUq2
o2xVY8WAVBSHse6DU2hGRvo/k+Oe13DJ9txLw1dmnNg55qN8gmqG0+zKBNVpUtbZ
uBVZlVWDum17nJ10y4jPZvtgcGasPDAXW65UxR2oVJ21BdaZoICUMYaFdUehPBxs
LqXoNCjIbmYiZWs70oJtyPJUxT35OGMaO3BmrPKcaxXKDT/GPwf6panrCKN69nXN
eeS282YPTPtDNK8JWWLGvB6aWpR27Z6MUepKS5m8/DxrACdXmlA1j5eQ48qDNSfx
IoVhUc2d+tFNat3Qyb/H9cd0cH84xYn5G/PtQvTtmSYCbp1NOOamXHhApgJKQUkP
WvbwXXKXKgPdnDx5gIKhk5XWiK5otAWByLar2Y6615TNORyinCWegao/mWFU65+0
qNa9M6lKm9+f7Bhq34iJqbMU6suQTutFuhdGULsrFChgEG+vPWFM4Q2U9oDgFhs5
eLoyJ0GAwyvnU1gNvv6CVSeQpI2eAUmj9x4zau7V1XeOr2Oo8kKaRftoAFFs97JJ
QsAsPhW3+1nbd84stN2xN/pKWmB7u2AWq9HpItaZM2tyx6i5pj0JAMBPTlnDMW+H
Om1pMVyFAzDTXIWOlGDFLNKkDbk1BbZJM11jYtRaYn6YRVW82gn/TeiM2WgWQpU7
xFmNU+mg8C/2pxfsyXdu8AuIxmkSIoEUGCUnnRqQk3CmXl2Z0DCAdOCsStMi2Ntk
GvLKOb/2MwfgnM+xPDTihAUdYafss/+8h4UhBjTJMplUGZoskYqcNv3YFO80J6CX
cB0PG+xm2Vn0xy7FoPiD/HYAgcyPNYbMfvaWPz+d/R1iAsW6hdg2DvjFe8l/MsRS
pyGdDY6Ds9AsWsYR4x8SDZB7s38oX/2bDcIqxF+2K2wLbmkf8QBnxsP5KChKGPfK
wkHyrxnT0A1SDCm6k9bp+bJEezzYU9+aT+4/X1VGJXm26gKW23j7vXA4nE3Cn//M
c9QjzGfVbGwC1Zb0MqKwHM0mrAO6hi+E3ho+PyEwJIqdjfel5DXqRqFNAm+DUq7/
ZAb7P6lL60VQ63zNJ3pCsFYTZ3oDskl2A1VV6fot5SdYCYKtFRZJtD9UMi59tMKr
3yzFoDpAwkUkYxwn0Zg0SnHdJiCWL7DZNJkshAQGUsYXVREv85iXJZuRG0fuxF0J
LbfnWnsS7gOQ7n8n1ooVbSdVRvDShbnVm/q8SYzbXZdUnz1F4uExMxfRejgTiB/J
NH8n7PnwiyAhCj2toBqIiG+ePapJEcpdWgegriUGrAHUN2qz9TS5BQBuXhVatcTp
gRtgamPcdAeyDF1uclWIEIRNYMhp5DAoV6v09gkwn8XT/CUW0zBVrlaEOs+6nStF
CGt96fqkdveUBaIAj/54QVf8LMW1DKHFe5KTZxBJ96+FDxZ8+s1qJk5QHdi3oXE7
CE63avkqPqxsGpT3PoBvTiVGGsToknVBxwA7vafRjIvtc5mnnBpYu6fAoXyHUmk5
RBVEqFFQrodjAOe5ZGhgR+h8Rubgh1gEkNKnAF2HgUiqrdcpRpbJnktA4wevcrbk
e55q7T/V3++XrFtdOCU4xuAmjH2Fg9b1qhBiivCxhYY1VgCJuITL3Bnn0yoIgBsz
AL4xD60AZrgF595MznX1wARL/hvyzNB6bsviuuV8t98gBmipUmVSZZJD2G9Y2V2L
DrqtYt1YvJywY0WRB+WJmXoiaiLjlZxsN2DNnYr3m6/BAYclewS5DCz6T7IN3cnA
ypexeRQi7cA6wVwTjon2D0GOO2SkA8Dj8Kqxle6xhn6LqNaJDHI7bTkD/vDVAA3x
EacI1xMO2LKkYICQc9IQ2ybFg4tesoI79yAacGkhu/ArW7kpUEVxoZBk6yNRWjyt
FJVuOmBBblizmI6uPjkj2bfxY9tpSs5FinMDytXoVHzh/7j8xA9DizTCTcwoQ68u
88kVlQW/Hegb4gYric8ke47rPbid/HEXGZlhH86eW/BSY3IKZjXvDXZZcogr4CUd
tJx+6Jh+mqyYxNNuZbrJOM5VHZFjCbDfhPBSdUfJw23ksRDLnxhnx300Qe3abHJ/
nl6e0+75pakY2t2DvGuvl0GxhEYnv3PjyZ2YJWb5zjGGK0nE0TPgwOjzhXH7A/3s
+P8pnlioM9D6q3i+VHs7SZf3h0tGiV/ByU2LjWv5Uq+/Oy5YYN97lpPVUqY10H/h
DLGBvNjxjvN8bLXwjG/5FgNTOjFvunQAwe/Zx21Ai0xeEhltpe715OcX5GArPTHE
z64zmdBCsKhbIa7/r2GkDP2D/GVEV4VoVL8BtQYKvEd6Qf0z9saVIGCespdIffIW
qOtpHRp4arz66e7pj6WqNceZ+hVmcw+dw+I4ssnfHDdqVmX9IuqCb8kkqLaGjpMi
A166s65l8fhsZxF+wEgTij2BT37PpTi1JQFmxYY4dAbsP489cb6oHDJgWNdthvK5
jtpuoYfUgdECuwlAdqf9ahUmCVXiBipQJPuDT/v150CCsdzgc7SwtlioA4DulYcY
EOEQAxNAFayFam6j1+iUmbXQW1WknRzN9ulQzXsigPy51qj1DIOx17+DEYGrVnf6
QSlKVB9lgAnelRjmzV4g0LCwDNIHEc52XAwBr/K1qSM2YDgDewTzVgpXMNmFfVqL
ECJU9KIIMn/RYlwATZcBgp3S8ZN8aJNoBZFzNKrU2DWB1JgLiNnY39dxI6P7/GjN
OYSCAl1/D872dHh99C+beyxg5SJ0SHTC9f2nTGg+dajX6gPhwX9IGopJd/RU4WSE
Q2cDuVPoUtOt8tP9UOcqhh3j7ygq7sd6jwjNZrZnTNS0ekva/6yAuEzNurHJN/cB
jATLzPKJZvaUzYTmA1o1sY9+7XZ6XYVdB/1hYQzQoMjc4qh+eWL7cVBfgnaDkaHG
Ojn2tYLiHCbXUN7ioyGO7PsY8SBvVVQNUeSprg8AqN2vVLmz0WqUWHqOOm9Pp1oN
j72a2nZSmrk6qMKrcDdJKPl0115KWuwg6qDD739hFY/8UhTls3n7YhrgZz/GRm9j
Hui8DBfqeHMaNxO1IGlbuM65w/UruVSeLnKvjDCyDMgWzYKOIJsae7eYwyjlIeG8
JTHjAW2OQH+51ecDNiw92xfK9oP+Af0rk7ct0N5PJAj4wpVUFUEMc05xj8R78YUC
UrQAFK74eeLYoy4rHdt6EoXtY1SgwnIuzXTyDdGWBWJYU0VNiZBX5xYxy7locgpC
bGNrlZdpSBx9zgDDcA077KYbdYJ++mY9LieLcbRknv9ncGtqCWvFBXiGxBgqCLcq
SZLPtFXUFvqdQDmYPegJYeMyANGu4QJQRiVz840TR4din4nuEVs6yWJXRhqOqZZt
bXqdXPR5qL3lC2FELgRCabEiJuOqtqrAD7GEV5E9jWoyDfJqAhq6KwB3kzeK4+3j
b/I+sDDU9jnodtoh2INbb5zE1yazwmVbld5SXtrc4iqgjI4vjR1mQydA0fXcKNna
+n+2uYEiFFbLCWr6E/7A2Q5JlxXdNpLiZtQCeixXDNvEqU16TvMAc0wxLWv0ZIRl
cEKxVO+gYP/qU8R26c9AeGPqiE7klMXPXKx12bOirn8RFkg5L6WcPdi9ZCIBZWKX
Q0VCCKWyYpY9mhDzYR21jqHw00Xpusui1Jcrypy/Hf2ab7hRMv/xpDgCDzOMcTfA
DKHffCmqq8qm3IuH5cd+WxYwoCtsneNh6cp+y83ae0dnewW1Yp4i9CK7RGaRbsr/
VTsDL985o4CEovTGWEhjwns4kVozplz4UzvfQgv2Ey58CGZ8TlXiLZVmZPGpS1E3
SeY5W1Qvpcji8fQfbnWxxH/wwV3/Kt6SkqGLdloU/v04thNrMTaampt9lltsweY9
No90u+acCAodnpcwK1ogQDybJcmmA/4UbCjSIuHcccR/vIj/alAC8Hz4v3wksv5E
LW51E+sE+4cIm7gii3uaZ/O8nStFO7jUzocAjvXj2n7DuffwKuFKjrKfxueU333/
/o9MHqVI5v0tzaUA25Qwaeee48wZj+E1UEaz0DkdS9gLwLIBLcImdYWwc3Xjaq5R
mRDDsPA64O1Z2+65To3u+ZucCAHHJQVopHwn2evqYAYwHRjy9X9vjr73xHc7MMVu
4f02049PBL3rWXc3k4YS9M6eONGylhsDzjlzLfz5eyZSExaD8pQDO3A1uj6cC2HK
MHI8XT7fhDmrNdMXI0bMRRiHTxPe08x0Z/fKXS3TZVO4rBNysuCM0esJA3ytHBY2
5UJjOxVs3+BDkoo/5ujC7IxcZLXborBuxMZTR5O9vKic65qT2MeRu5B05IjNA58q
vA9bvPrKhnX1BRnIVex9/qEPOYI633AKvMQnjOGrXoDiKLvt6QOt3Xz+lTiWlZP2
O+P8XzPDuv3DD1Idfdsr6/5P7wuOY/ZRjWYY5ynHZw5X9QVfkEqQl6U2892JW30e
G3jGM+1I9wZQN5UITfUq9E8wbyn9I5bAdoUYw4ygfNr6et4BIU701QGNFkQDAwBh
EKiWTvVXOKzep4pqj1Yox2xFUMJXLgWW96f/d2V0GvZBSHX/iZY3ZsBUZUB7cdkc
28/hnjaypZkDAzl8Zzhqr6lwer3W6JsJOycdAInOaAQONq0eGcJJkehKwc8UeGPa
k7IhzoLsiljb/rEMj2qSZx9tng/ky5MnbXRHhT8JGkPDssw1UZDFYwAhgSTYRPZS
a3l3+gm5XTn+Gvz+kXm4d4Tdlzzosazt48IOCopCP3IUeKG1e6uoMFy3XN23rVIb
Pdz2kAUJL9wByB+9/TV5XsRUFLYavKMIm5J8UDrYRzF0aUz/i9pwOjWX9BZ+ryUP
bDKPKMtYvULqLKdhDkxqXPTkyrKPiUpVErwupvQ55QusryZYyfO0y4kzHRjZBrId
MTHckLr5VzHwldQbA4R4XjrvBGIZ+ZYtvtNBjxtPygIbGjCiVKY5jOmN5Nw+fOuW
hOBaPNpQxoNR5KgF/FsU6303t5inh+N8V5flUFR+ZtpRrC/XWQK2mqqhMqc1NdPp
5sIJKwwCbLwOzZZjsd+E+leYKvExINWvzAMgvd7TeQqXBk/XhwjTfBBKAC8WpBFz
6WKvXiwabSApRM5KVCanmhjlyIOUAGkk7yQnugyR6/lra/0P8aIjW5/1oUgC+erK
fLJRYMH2z1L/87TS5/sA7yJQ5aXaBqNp6eHtO2oU/dtJ1jXuiaL8ojCMsAppglnO
6kwJA0s1WWS91aqy+ZowMQX2uv+wv08LfYlJQmQ8QA2AsRR50cWns6afH1n1b7dH
RMz4Z3CmBAEhqjGJx6NM8pevewUbx2h18OVsJVd1B+zeQ0V9sQFmvoMRsNZfikT3
VbMffdEeZ/4QxHKuQmFWAHReuwhQQPohb7Z8XPgmJXN+EahiHkIc8sEkYPWIAXiO
V5YBfT28OQ761/EfaIS6IW6tMxqBtzULN89GeD5vanC9H7X0SS31LhzKPAurrWe2
W8DCwsk5tGAVqCIomHdAQvUDzfeOgWVTjFtqHSgOP7ByKem92g8hgBj43c31oinM
BTZdMF7P9e4O89Xr3ljLrkNzcAXQfRgT/ywBGhAY1QoEzcugejfZxbnApyzVWlaw
8WRccyY1WFoB1v1EPOlxNo3RvFlTjCcBLI6cZMEgba/Z2zSBR6mQB4MkyLotdamK
fnhliQEBoy2lKb+pha1jb/TMoL+lwY0DdzhOlHaWKRwS6Kph1x7k9dGlrtFVB3rr
2P1tpn9aFTEJcSMTacl6ZXbOHx5thUnliLpcTpuuOHeF4LR6wz8PTIMnubyrvPsj
8cs9D2zOtbxTFE/RXaSJ/f2eA50LSH88lRc47sVZiMIAdRoqPhgXVxuv3Wy2AXDI
LDQS/dweHGSF3ta7v66hYm+YzlPqCsbiCy2ncfJctZ+laPAB59vufmO/QQSLTx/r
IkGmMa1Ft8MJMGBimu5agBjbBPIVnxGUPXAHFF+MN9mmsOWg3+W+HXim+TX/Bt+v
vf1vGCGJ8og7VOBKLij4i6m/PSCEhk3FyoO+T2LyYdu5QEVtQhQYwtk2NCFrYDri
5ZX1bu0p01llCKakqcmgBsK+BVIdeadM/IftNJuTYRnl/bn3+cEMPOUgRuuwyIRJ
Ao9NFclea+C2hDD6xfaqs6da3KbZwxHlpGd9M1ZudxzGhla1fcMAsqaL86CgNCK9
cHnxOhrKbEbz//0q+wbq9j1tPonjfNz1excYCQYXe8H3nHDAC9zE1uQFu6pcO5nH
nr7gvsAXxcOzBiwY7H6fKx8AHJfbMqbOqLbTGs5chl8MX0n+Y92GlgE/lSe0K4+k
juzhT/5K7wI1XheND69ZwjEHLJRmFddMyyHXgkXJI6QL7QKCs+j9ul2mtHb5UMb7
5uUrJb0L5vELKB8i6Fw+oxXrx/gj5pL0ysCwQ8j8aeucsY7oRopI1Akwj1Y6zgUC
7tPMPUvbR2crCylOdXnwgFNFvvPWnOF74VNBBEqRfdXNKNGByJ57tTSHAvHItq/a
71YI3Njy6rtT6z3mr3v7RkLDzMN44u2Lr156iPjEYJSxsQ+p3TYZG07EuaPMtR+g
SeQJkaDfs5PA+Y6rSA4JZLowIIIal89FBpXBiRbGbEmTUrX7Qn62NzXqJy/EZtXm
wNwHKI9Gt8k0nKoUIQn1atb92qXNtgwtLciFrAskgq3h0Fdy3y1zQ6P39ADleiqp
6DV/BFfjKJ1445MB+bqIIAb3lSQbMglDxdvXh9YcYdrURldanyGfxjP3XFlrUHfD
AhXVyf4Q4CRYEWd7H4MY2hmIjs8MfwWqwEtgXChTK+yNK9TYreJceub9Fose/U97
c9BWQwMgLNWazmqRczRKQWyGF9eoGUTCA4ZJ9Nfc1AiW155siKjKMnZFgcoN3b3E
cKMeV/1vmV1sR39U1G2wPPSQinGMQSRIfNxBHt3SqDjRr8Bn4sJqKGl/jzk0HXJX
sBflumjWL4HSjH+sfiwA6pP0KqV3Wfr+O/aOWiQaTWMr01oj6RTU2Dy9GOtML4sI
emdvOQ9tuI/hvlNKCzyjRapzc0voHmlYJ/ydpgcHxDKgGA/CUfj5sifnqC2e0bHl
u58TnI9N8nz04cM/Ws5YWgkUPp3+1gq4G/sHWXkl2cEy8TZQTWVZWWgifPwL39UN
ovCBy0F5gDrh9cemePONk+z6j+AeiNYZ+zSIWv3OVdSpvXGkO4Q6qYBqN/wZE9uz
kh9gDhyeqpXhksYUian8a2Wucn8bMov495aygFquinX8ZbZYM70RBEzcNRC142EH
Nf21n5814YSIzH0z0KXlWG1mNt/Idcl2f8tms++/fJNMPT/GD8IsN3maa4Z31D6F
Px8ylTh5R1J7AvBJ4boEnX7+dyRz6Odw5eYzswfiEyS1CieVCLDwHmctRxeLXzgs
AmKVpKFNTZ8jcg7hERBqNi4m6DPEyjidVoWFlhud2QDHIVcaaH5gG+Yk72WvM5IK
O75USEFS9PKyORwLibT+VQ8PRYHM2TyjVxxAYU8pfD27WlFu4wVNy2srZO3qXUaX
2lp8XeufyvQT6+EqM46MHERGHGTv35UHVr72ATjUuFvAVzHM+3TnoLEMstdKroa1
NfsHLfqD89sjn3IxhLd7+JcKFNVphMXXYrDctg/WOBRnwcSrDX7yHfAYKCnjSQRl
UiFIpJ/cI/+WCL0hQbqLoD2g44JHD6+v4MrV6eU39omMGEaaArJgdwsDgI9shtq3
9+SyJ5VdRSj3fYXotPN1kQVS2Ou6ACLLhQYrqvcQ0WXV6xD11pbR160mG8LMTk3l
1r0Cdpn4aPtf622dUB6ySyo6VwN/1ynuRy0xu8n+CuLNPTsry72qsWacbXliI3C/
GHdm2Cz4h+wpy0BocWWZJJhqFHAuZ+gOeszLdGEJz0+9cf5xNLoOaRuUFNND/nNL
nnFWmHy0RhePYriugYl85SlZgRKIJ9G5RNJEwqyHxuI8HgzINnIsLS0+euNpEUZC
9TRmSX51/jv2SuhBC8P8Kq9P55dMgDRi8X08zb9sPkoBStKv8uYw3+sg6yMcn6Gf
qAac1G1+uV73LgPvmJcs1DfBgwx/q1gMkOh7A+YQ31oPGQ/VGbCzP41eFmE+afL4
vg5XWq+Lgyv6Dh3wIuFtA0/JI+HUivuIErTp8I5Gxla3pIw5s7TgPHx59KDBvqDq
GJC+igz1/BGoiL8Ug0oRB4iNv4Os4Taew47cghc9OiXEUKRsgvBQj2Ahy/HoRR/U
9iYoihRKvZze59HkaljaDcDsCY7t9jibH+CHYrh2WK2ZhFj612xzyA/behDKsCCm
7XtYPPiKEtZDu699jjX9ydzqqpoIbmFyjy3/PPa1Y0WyK0jJIC0MVnmXzhImtvFh
bxzRUFkwNY/Nx4Wc3hphclxD9Rs6wlwe/FbhCWS81ULaKAUv6ccI1AkUXB8MnpCh
NmAmCi4/Ngq8uAxF0Aba6IwPVIt9Ows89GFh0GoONGLLDLByWswZ7aTLqhQNgLKl
7+eEJHa7yjV5RXvWd26nSUtRyiA6E8FC+McGarLYLoJ+I9QzDDwzz9wo0znMGvcb
4xxcjf9tO7OYNrTBTBf8YrRmFldYGdy3Oh1Oa08EEdXCu0tNrS2AcdPljxgvPbXG
6s5EnnNfWupQhqLRtIfSVIt32zx1q3sdr5hPQrRYe1E3XRSrMXrbP8iRT3QuNaPE
GGwDNxxzZRVBK76Th4hdF8U4U1m5D6WFmoNmPOmLWFFbQJG37a7lICQ7SC1e86kt
Rnodenv7quCAiScIRDAr5kg8pQZLbhNoEo8DeW+5anpj+eruvLJUrP0dy91qZZ1L
cTN0dSt99Ltlyxac+4Mt4ejPJNxgEvME2YOUauFatZHBJJ0DCups3FrYIUs+L2H4
FmFhjmIRglutfXYRNfcNMB7UXjEfhnLNZ4LcjxE9rJLUrlSUnrwaYKA4jIgS8P+l
MH/RHiqxU9WUH+3QRayt6QrU6XUeNkEJfkqemEuuWl6jHMajFSDUz0WHAvsjWx2j
hiY4wu52oDEyY1/12wALGyqGsWVG918gH12jN5IvtsfJ76qWowhKw+zUE+rFsrzZ
U/gWbyjFxK86PX+TWvVK88VmWM7MjFb0fnWAKLx5ssrGPwyXHW8b7r8rS2PQeO0E
zX06va6v3wqEuGXaRoSJyUpqFb8zp4BmfVztDOq3riqBLbwjTrIF9GoJdeuI3wPt
WfsQUpBEuASg0qbk3/0CCJ/XLSoCt0+C04yG4WbtlBTQTwtjmGP2R0EcUjS98hcp
hBN6mje0SzfuzYOECY+QpK0M4a0I5XYq4q6qhRPZDIvphSDiNSGqB2KE5TcmPjEA
CRP94APJOmqCNZnelKVSJs6HVObBvLFpY3pGmbTlyuawHV46jiqQXPFMKjx0/YLa
I3++PdGzWhJigERQRoJl3dYMToSkMoRFR5JrdP3mVFuMHQYCry3dm4KO++Q6SJtr
UcHe+qWJXDyQTPXfNwTeNACB6qNeSkiBompKqyEdVUEttbjvK0l2NOglLOEG2Gtr
v1GLTSpeqi4KzbDccxnBFVpYnyrhYu/WVKBOabzUcdk35xMFMJDD4YxOEJClAzDK
SaCJT6kpCkBJpi5ns0iOTEtKFPU3Q+0IdVoq/CTKY+bLAjYiz3Rnq4jlpSxyEFSp
t2QYF4PKgAqMhTFhjoAYokolu/Hj/AI3RXEaCTNhmA6UEZM9qqX14NPOezAlR5K0
Ey4yQaiOIC0VleDvEhwvRO0+j0GOvxp7DEErQayWmNVdai7Hr99ULkE5aXMrFzw1
02WP6I+vvCP4X4z81MLc1PmVLlPyuF+oXQeA7yjC3oKD5Aq4d7ARfU8KdELdWSPG
Ly5UEqVomnBZpIQILfxbATpuo0NR1BJRsx7O2AA6G21zUuTBmKqlCe9hlmzEFcUJ
d9mAk9evGqHTzphxpGKwJsJUHgvEnisSy946AwGXUD70k9sqkxFU8rzWZcDpGs+D
/Q3ALr0+nQT/5X+paHf3ht+xxT4JsVFNDYLyp8Ru7r+Q4YN4K3y4TN96QuaY5rBn
+Tbebgu8dO9GVfh8FGLFuqSPevvSBlx0cjduBn/byhHm35l2d38KfTW0wVlS/j9r
/+zCme3MoNeknuKcvOlCs27Tmeewwe76zZZyXzry1kDCRR95hNZZNWwhO3MIbDUe
36s5toh0Ew7rgYBsJihw+iq2ONhnkw3Mqbqh1uoE5mMmGcO1wa4ebES6XIbU70fU
ReahmC6QeniC40RPcMEcQe9nkO8ZptUj68/dpkwwSefR0DVjL3ToeKNKtTE1PhFn
4xATaqGQPLQHjM/EQd11qaqoU+RdQG3R4t+P+S1FxMcTaxBFfOSj9Qr//t+0fny+
FWuX/qKK02LIHIQSjaGUuB1ykLIWQ+uTDxAGYI4DZUL/zEFjm71KSi7TlHoTFLI8
Xxb6hmHTdpkAp+uNNkeHywXIZGKhnHqb0+LcRbtI1Nc8wExsCcFpbjT5HMZJyIA0
uLuKG411wInSV8xTCbzJ5Km92AQu1rqm6sXp0FvnsZ372zbO8pAgeyYLyoN9+sc5
HvAilb97HQCJe+E8tz+ZY0CPG4700fhCCibvuXgUO7quc80VPuB0ySI5b2bJrxgG
am7tK6HZxcI1+gDNE00G+P80IOnpTynilA4kLyMtoKmvWo35ifDvANefVQpv22rl
2d3Ao/bKiHyISZBGvncKibHwq8Woi+ZnITqEqaflc3gv6AzutDPDVGXDC+Ew2FVt
OAigmKwtYDqG46ykaof1qo/C79W4PRpZXuG962yC4fWo0+LBDyf4CtVASIi4Osfi
409wscVK4fMGvihocVbeRIHV3P9VqqyXXlbrw+c+Ql8sWbgKO+bj72fuuNmk3sCA
S8qbhYG06eiGNZeQP+QlSYX17m0QgxeICxw8kHTMtIq+jMplPOuDcrEMn5Si/PR5
HRiiAtGIXiuN0QVM9VqBZgN8HT5VbMuhhhikDCNC5WThfYQAJ8ExibHZBxmUp+e+
xgug6CZquSwEIk6TDJt5W9Cq5D+GWrenXo/n6zaFpzWiK+5Kiyl63Id3HLArRolO
5T8gH0DChj2y7/3+SRsHoJjdfz9Rl5doE2xKuZwIZ3OCF8CLT4z1R+yD9zTi7D7a
U7n7pzww4SS9/v3c4URh+eaIv40ZqA9tjxAJ2ZTCTPQy/3/5dk15T2hL7jVRjUc2
qYJQUUFNe4InQG7uSPdAXMJuYrFD558dD1ab0/Df9EvQKtyjUX1z6V7cQJ+AI0PK
+KEW2/6g6YEtGjfYTsa84wbtaqzOHRDJnlqMD/6jIm8vgSsxOLmA7lM7cCw8nII0
AVEETE53qebDk6mpquWHFDhJQpDebQuIoJMtS5T9VO+R+mOzm2e+NTYFMC/2GFj8
4u2qaGoov4RnIFViY6hO8z2EWHrbSdJLcu0RZgWrOz9O3msPcS/Xlfw4FOgyHLSP
B6clzF3SCFK2m63qiDeWKiCoPFpU6rZlV7c03n79DvjPLamhCoJcHlBvIIVTDcib
GD+a8Um8x7Wb11ro27CkADfy5wNIGjGvghimM0j6XNE2sqTze8F8mnCAWpXeZfsV
8/gE31FjvUpLFOhQR3BiLyu0sSQG+SmLx0vDL/yvjLnXA9UHK3SxjEYsLojG4YuT
kSaZrj/oKkw6Rp5/Q5D1l97liDAyrDfDnjUnibEyWcSZ9SX93/s/pmW8CG6NJX8G
uFjmA5lf+ZSipwaPJsar419bYra+lm2UJJvaeJGoXFwl2UU8Q/RQQkXMlEsPKKtc
D5sd0bQAR6r1E43SmHvz+gY9P4Vp4k00IMqCia/JqVAN26CvPKJzMSUULhtgis62
hJqi9S3rF6/1WNSwOOoTFon3aldKpzdIm4+3wK3qZGeDBFBNTn9WFvAFXohtcFeU
zbp4Ou742NjHoWihVRhwtQSJVzQF/QD06kGSwjo7my3kOSfvoP0TPvoJ+XjwP+Bp
OCmNYK1nltJMzkE3YC0AIEzfA2Efgr3lkQxt0fwhufXb5T9yCniDxJbNhXUWZuAQ
0Z9yfFEphy+khho4Y4cv6fEIej0TvlMNhE0lfGoEgDp4NtTjhkCbDCDc1w0gRKaZ
WWafSQMdHWJktA41Jr4EbePzqMJ4/egINjKjB562EEi08MoKY/Pb3J8NkTZvpdvq
pyuT9INoGbUEOMrbomudUXK8EKUxVwVxjXWvcdsobvWmEd5iAAtuvciuscOPy24D
EnYjhfNS+uIMDuzKeZmABp5Oy8e5pnhtDMrSkfrLOcTGtrbDENFnByGhArcIll9W
jXvKRoHjniLvHUxdLYXIgkt9ER1DW6dw9lfh6UrQPmVP3qXLARf2SfTz99oo+V6i
myI77cXHMCY+LTnE7dG0ApALa1fE0je8YVnDuE5c30l6Uwv/weBCBP1WXkbpIPjQ
guRjZziZjemVPjt1bfv4p5fmrGLlrRV2qW2xhjrM+L6iI4GYB4YzU0EP2oeDs9ac
+vBk2EA/+W1PV4XuxkVOL/MIe6XxLzYMxnNaQwW6aXHV8lcjeHHLBAeh9gu3zCbI
R1zSxMrF3nVaz6uflosDtDatzzDjtrqDz59MegW28QYfIjff0E2iy8RmehWz45yk
j/aQ3AVrhqc4nlq6PrClo+zQyMSayXkqy8ujKZJA+FNpenx/VOu/Tpv5wxtGucEY
Cp7h4Lq96iLhpjzvwtAoWr0/v++6hV4RSuj7ieHvc5Xslbux8hexQg4IDwVw8yxi
sAcey3H6DSV5ye7wIe9anZWSKKoIB01lQRZk3dGKS0oolnMJu/KeBayoZEVZy7bR
Z9FHklLgmTM1SxjwgqmtIJgojjCsnCUgrIsWAza8NIZPZB4JeMhcXri+13guM69D
ZajifYGONmpoaLrcZu0Kh95zQjVmfsGa4YRPOuwCmZbBCKuprvOmcU2AeTPHqEJx
YA+wLX9UM2MgTAZKIqrcM9bInqXN8LvGZwuj15hcbpfCw6BRje0Jalsyvlj7HG/z
GGP6EovpleSsYcx6Jl6fTyhAWnhFChGBMhl7RUuDGzYYhnuLHUXWSNyYkcr2Iiyt
6usgGMCmSSSQ2WZzsomwqFrfIbANEX8UYvMfqgl0k26zy8t4IeDfx3U2k6ALpveJ
UDsCRmml+wqZmBBVun09Jh3f9uelIak3LjzWbFUOy16W/o9B1TKOpBY+BsC2Lp88
e78QRVVMVnLsUQxwGhWEBG0Es3sM2W9jUwISFyPSekievryNAzNg0UKCLM8qTAdy
Js7X5bFJtngkURZKEfhHxEf22VzcO92s0AymT+5qOpVagRKRZw91WBLnEpAyAXws
7JmOekEyuOdDYm+1liPVYR1qPkrBEH8pOuoMmfpaToooZKnPl9XUdk3J6SmNt6OE
Zy3gCTCrm4VFVPPiU0bITswNEqSLICos9vnHVOogA0e8VKyeE+nVG209PsRhsn8a
YagRAI6MEthCfw6xiIr3xfv2cvmY9ISYONQKkcpzbxIM9ReN5slwQieyVwIiBr9q
r6wG44y3sGz5qzou3lJ9OEBzYqwIQpAslVNlezEFN6XI2pkI9CNxHf44TltDcc9/
yMMYlgQkf8JdqnPiqY5UoR436AuBstf66wVL5KCtn3dtfVQHxoGWZt853w0EGQ4Q
aPp5XVizzLG3TTMSdkisoJVcVochFH1E+VAkQGdqemZKg2ulhSlWi9Ga9D9NXe7G
RdJy4+/aqNwg6XvNFRp/5SO06OKKPLlsPQVRupkHUKwztYmOHN7BXxsEokQlBf6F
Nb3Wf86plaItgh+Won7GoGEO7x8XB5FroEdV5kRZTRv9L8IGF9zqxfXZUudgcqr0
gjTM+sm3K0qKSBh6YPSGlA/K50BP9iIk8YBndlFM4o6JAKBO6Wlf4CyGyPCFSPEM
WvbtMLUhOe/g61N1JL+km7RHXtLkyTAAYIPdgHpqbGusEsi2PiiqeK5L9w53ROyN
zjOMZmKSKubMvD7CDKNuN0KZ3aCWGanx1rRURYVK27kQXWLH8In7xEuaWG5vsKCH
gk0qkwbcYzvNFLOf3IM0xlB7cMjyKtr/8HSEgt2hHbmcI5U6Berd1J4u3+WNhfEo
hBMkskfRoF3yqQRdbOt63L/2frRRLid6X7BhCgcT41POQO0w1nvwUX/9ycMEO4tB
TkqbpirJ5+Ce8rz9gVfAnOIRJxX+s9FOaeO9GQiztCKLLRkPxyX4EH6h/A0nL6Sm
lJyc/vQa+YYPDo7LlScrOPA7/2qxP3m/fdjkeSSGOLFU4AYvR2jGcp1AzEFsVuE1
wW09gjE2tnsNnR+DkFVFwuddRyC0DHV48aqDRdXhSWqdcIJ2PKlLzmF9r8P6Rzly
GJ2/qy0SzlMjgUr6piRfrZ0yccgTfujVSNgEuyeax8Vi1nixAWvWczipjAzuH3VE
SLC2qZM/tBPLL0IPLLR8CDccAtCme9mMdyVAphrLgL2/0xvedfoSYI3/WF9rwaC2
9xeLX1icRDiTYrXcJwRRgVdk/flA5F/z9gIHiaSl/9ShrQ0QaJRzdokb5UGujrzs
oohputkxqz1dY6RBXWRTQPRZ5Pm+srSF1tnhJSN+ovWi6L5l/N8jMFY+4X3uL2xG
Is2TsWx5Skdsh1M25yRiYxYQaHEhsacsaSsIY2HWI+BSwzkKIrJQ0nzvOZRIzEO3
lohAIWfBmI8iHQtn9b9RQhmBvgcYWe5a8CT3KNDoB6pHaMN5WxoGhRNaQ0RdJ8tP
vEwqPZ9vJ3tSlirFhFj+lu43FEVK8raAmJFWFZPIAErMekje1IxM6hccut2DSkwf
q4irN2x1tNX24+arfs7P7aCe0r6Tc/A0+gDZ2MUCjkOmyykdGbx6n06RP37Tsqms
IpiH1OmvEaXUIDUTtvOe/OiBErjZPAqSztOpfkzTTyj1baHdT3w0UxD4CgiyD1Nr
6zwBvQgyut4N+BLuBAu6ln50NY0M0eOoIqIioX1UFcB9YYzA4Y0RBd1klB8VM4Sx
HHRjRZOv4q2dkQjVHQGv9NHsxot90fK8U2Pd3TiDjqpALkDJv8Tc+PetRuXuePIx
vCT2S9V+qZNDibBHSFdlJodvC81wOVQ/gKypKQWDwVgQxXScBjUS5zc0IlnrafW3
H/ZV7KIQ5rsLFpDrxg/xYgQqLbiLFbJlIs7njc0y3tew5KV5aDO2L9ijxqrX9DWv
FwmpBDpRt3kXCiEZP5tK82i+buMlKWd8TNIdLOiYuGdeMODlsJS+R/UZSEfKwZIE
HBoM9AnD8bFddpPxla9lcZteIMT2BVa4FHUyzzRnkYpdH8JA7Eu5y+Kapbpo37Et
QnsxhMEtLGwfu3kaZR0wKfSI8U78TM5F6AqPl4d991RVaXcflIAowdtvY7Al59K1
MGTakDJg/cj+pQG7eJKnzkTaBZZq9P/0gZ7wDFfHU7VdoO2OhoD3GTV8UaFfK0a8
uCE1t0GJavluPDL29DtmOEE6SrKiQ2XU5VpDT/BLmBta+b/H3c/Lp21/sq1utZWF
hYj3KpamS6Wj2T3JlfkqUeCsH6imthDcHhmpHJw8HpXuNajUQHyKMu9npi2aEpxx
PxI7tK0I08xwJ0gsE4x9BpyeEtEFQ/+u3VHDcdYZBXKoBnmxhrhy2rS+mMk6dWyo
P4MYLjRD4/lwqJ0di9f32ewDRVspTsrL9qGM8hVn9x61zlCWzNViC5PaAh0uZKus
NIrNtI+2gTNOkaCMfTj7Qp7KDD2RtsknxUX0wnml56Z2j0w+qHMs6ORq0bfyPyDs
wHMb/O8HYapVKKEDdeF673xgaRA402cU1P/7yc+ObYZ/WTwBxSKXKNJUxShvmRTr
35MNmVCaJGoOQVbBQJ2JGJ3aC44xXRc9758f4vTcMwDCEiMCUPlkEEo1GryizkuC
RjKDLQL3fLwa4ZirS5EW4P4rNKtHl9u/W6p+/6xh9kZ7cuCg5HAQ8TCW7AaSnhqD
y5yDhgT/kdDZFxkvd2H5xa3MMMS9wR4ix8RN5wC6u5SwMp0qSI2FlZYs/HPbesLZ
OUDTcura7mcTMAuArsxoB58o+ZZD0ZIjeiGAOsss1FhHTtXsjmDucdC0Js/S3E+W
zGgNCkStY6mC8Ulr9w4MZoXQjIciLh/j5kNVpKSLxY5aNAA0/2a1HuVCD7C80LGa
QohjoRpWABUw+G/tIh//6aNtvm6N82nDru2XBkEQY8fQr/82Tln/vYozQzndaVHy
WdvpHeaUjawAdxF3dh0ZHDJkkFDJvAO1/cDhzDzg4I11nXlTf/EG4xZ0UxAC3PRv
AIWFoI+oIRdh1UdAXcpyEOBTYrItC43NEXlgj3+/BSPJvu4Z8ha5aurkbkjxskZg
etVA70HefudMZxBMhJ+necUTp4op1R5kT1S4cYpXxszpxqqw2TeiF2cNtDZ3ymbv
CUQxTyVgU9H+B7bnwudfPvqPEJlXve2QWvODpcEyb/DJhDIbFA77qjplpo8HiiHJ
2kJn550qtrjAsE+tAh24jTbkORFXAO1+nvzAyJQ86+fZGSEMCPnr1QzfCSTeGV7u
IXDDSbvBbct/GslHrLZIag6Yde1nfpGpDs2VsOk/bh3Ugy8nO3kAqTBUvlBrq+Fx
k6Ni30rzLgApUp7e7C5E7U2E/7Q1Foy8l35R1L2VYaLeV3gZuWnI/munRsHwBvcs
oc92UJYpr2fvfUfRKOaLCXS38LJU/9Y1AvypiggMIBTNK5eii0ASYcR6lZKFjiUH
DfqpjRRwEoMjJpE7AUxsmgrF+3n/37VCxiYHyDSzeKd+mJ+s37HSGEoV06l4Q/xn
bLsB8e7vFjAee3LowlhDneoPpwUM0m4giBM16gHaT0iqA1RFwB1dr3noUxogugyy
XyV9xpWakLS89UBP4YFv8whBW9cMo5rIo2CRhLwDMBazAPqYZoq9hA3tzQIRL/7C
pDZQBfpVY751SXiQ3wvktUTGB2YPuDU/Htk4ySGiRU/ddAEzhu+u4Kk4Q0UBoyOF
W7aqtqYc2UpkHnT9Bc335xeJi1/2hdfc7WbcZ4a1HJXLJLlk/4ej5J+YbrJ3j1E/
2M2vFYQkdL/MAcW329ZJSVll8cmjmcZ86wVK7W71AlbZhqIY46UZPjT1Rz9pphm5
aPTcVV0pE8TMN4fN/cbzWPVAjoTkH/cm3JVJIxw7MDE62A9N8Q75FwpLa/aZjC03
EVA8aSPgGi3XNFZQ5BhIj2QuV1WkiG4o8e338Iz1h2vw/d3Pk4sjeixQElXjC8iz
CjxgvrUHSTBchU0BQnL10KuHaja6dqdg9zW8eOV209slb7hwM01KLpaQ2SzfbcI6
tAk8cqTRRMaONVvDiM2dpvYUIqA2njQo2mEuDkNXNLYYCstyZ73G9Uq1wjVc7AsM
SqBkuJ5p4hMW73EAfnZIiYoVdYZYL6iVe92wwYsLTiCZTu+nZkGP5BbLX0sEw3Wv
oAzVcelY/PsqoZ271kXLl2nnecPQ3WLX96g2AcYQOAXM0WbruwEAXYbcOw8u3Ez8
QHDs0UNPR9eoV/VlWJHU7a9cbgxBxCOPvLHnkI0SiwJhvg9W8dsErcl7vuvJslLZ
ISGuFwaMXLNmXMm5bpTy9Wk6AXK3JUUbnpC7P5HzyZnTiYDAcMARgeZCsOiFznqk
I1I/lQQqZyNmrmL9eMjuc1xdUmYUgDBE6S3t/oydLdFJrIJnutcPKuEWAF/r4j2N
YiYt7WZatr29IYyQmf9RGisHopnKZt5aBI6b2nNEwlHZuc47H1VF6WkaJYa8fHb9
IBMNkbplbFSXnQrO+sCuBkSuc7GV2fASukXmlWOdMxKZgqv0zNF6d6SrVM+j3Sl5
4a0d1zkClNUzKjUOHHJf9hPfy7eEwVVyKkaP4zBLru5vYsIqxzOzmOVnuqSvM4qK
aayEsu3EMSiyPOVDATW5kkknbVyg3SgdVEGrr/7gFOvNbJc7PFBPh+APU2YH9vho
g/EPbLFlvNQ2nPg5lgY1Q4wGA/D92Z4z/Ic1Zd/TUbl26IbnQ58t5wXu5B2j26Ri
2ki0zaTYtEPZlxSqbfdZuuydWuaeigAeUEILK+tFxNApBHlAzjLKlhYdmYtdIxpD
Hteu7pvK7zaPUSKL68RIHK+kspRIw8VAeOKsaYgemKAuPlpaXDKXK+0ny0RrwFor
R8w+BJxq0PSPLq6jyFnCENoeI/IR7Wjz723O/ZjQeXpX6U6UaUXh2XYBBtXoTSCF
Orye41UIszsKgbZ7zwUFHyeDiMo29phAxlJl2voIhrQ2rhFc+sLKHdmNeGbA3tWs
u7SN3oRrTgNG8R+NT7sCYB5EyxhjSqKmv9+NXUPZhheIAAVG9KIfUn9SRiVwNFb+
zqpJgQmQbCWZ3tu/kotBjvrw+Jd0JJOMFeOIdRVDMWkerbRAUd1dzOptWrkxf8Yz
2tu+kopvZ1+ubejVKzTyvp4N84QVIfCPieFXi29VgZIXApxSEgxvoxqWA0KiT+qG
i+Rj+1aMwSH9lmkedPgF0SSu/Wiq+3Se75qaLwcAgeySUqbbK6NIWNVG4Ga+YBc3
ZiNi4y3LP76/McRvYxCQM7mII0MxVXUx1Gup03CLc4pJwd/EaCFWfhZ2wvv/hnyc
ylLfq9fyyIzIMrIOn+Kh/pD84qfvHin+dssfMHWPBsmk6AY15wwB1Be42EbgDjz3
jF12BD81Biw1gBnmQx5Gncap8Jz3BDOZoJzCpMoqV/CmvmRWxWl4jFa8aqMnR1Oe
6g39zz09+d+fUM9MlA67pEN85pz9dwEOhtlsdL/0KEm84BqFmsJLSFQzsnh+WF+b
dWPa7a409YmcJ7Q6gu1ZNNoCO6AioB92HyZ6UsH6wpAUerjnjGvdHD/Le/By7HHE
EW1wqOfO/T61piVATZMtySCMBd1hrNOZqcuUXA1fptcu6eTizGXDcP4uh9ZnR2s/
tu4DVv8OtY00hpMx0/hu7N/PzkXk/NCrgmzQZ9WEbvI5t4IfHFSe6wMdHgV0i8bh
dT+KL/BUFpX6DVD4qbmcBTdrTOdti/RfoF55zNb7Mg3fQs3OXdFNB6PVUKnHTwg+
VQPpbhxrXHMyvHmuovPxeKkprzeawVXskjx+mceveFrh/KrsyiC1gIw4vEf9b2Wf
3DX/De7t9DlcxR0NT0AOcpsd6hOcczPCeK0UyRhqH0GlQMmCj6FopbiG5QY6eam5
SkuE302Pj99rLrmFp9eua8+LMBFTRknxHO+1G5XBqjN4GFVZ3C1fnbqvtISJrwAP
QE1n7kaLLhxzddhRU4oyrSsH6QfBSng9AmwSGgbHJiYo/q4bnQt7C1P2rSpWUfE/
7RDS83Hh+4oeEbWZUiTIRL97poSsd29HyLW4Wv7+SNdavwII82KUsx+4U3DuZyel
geSmOtdR2bZYEYOu+PMcuPczriCKAnwJv2+4U/05E6ZFZBk8oMX+k1t666WJuRkr
GIC3QvcmW6maZq6LKcWzBUGjBcOqFV8gfX+F7bvcLr2UUbOxFfIKlpPm3APo098V
pYyOtQVzFuB61zsQnPXfqxM0Ptuf/ehs1Rg7yK1g/7l63oAwg9UrSocJKpdEuQAO
VpGKGo616dQFwpikSZ/EcyhqOHh9yw8Xl4T0i17bh/9R68sZIdVZ3Wzl6+GJ69r9
+IiFIUGISJae/g/HIu2/wwB2qAZv/bph7p34iSD+WjK1I9mIIRZ0g5UKlP3IzXIP
djHnbPqo97Bmk4rgE/YC8SYrzYFqyaZYFT2EopxKoWuDoOoY4E/c9yQI5wvRWEap
0XJHDx8vJT6EBjecLdUr5QUNDnFomwDzaVyB0X6HYHrUCATXcmTJm32FIPRB+mOR
gM5Bi3QWgGyR5l/xKeKxAsODjzSz8X0HTSTmfJEqA+Xdd0hjn+IqlWKZRYT6/Z5m
QO6eDtMPWWTfjkIuvDHtcROYzidvUhcnJX5cbsvY9OohfUdAiBNeJ4dxeX66PSDa
6rOQ7zKv7nND7J76dHBp7VTwoPrdYpQ0PeBpzEIUW5hV6qflozeLqThdPAO9TqOP
isK+YXFgrRUg2rK4vTbmGn3k8qDbGnaKbDwC3Df2nSWxq/3qJzkutabHELhCwMxE
Y+eNk0MQUy8uIDSr7ZV1n8Sv4DYYi4bFK64KO10VVUEHzoPZ/l++kIf12+7j1NBC
704rdKVw++Uq4rR7yBLDMG60/KL1rn4lAeKfBUnepd9dxMk1rQJWBop9U4uRYa+j
KFjeD8Q9cOx7bvYd7uUrgt+QfPE3wgo+LV58xOGo/IUMePMDAgYcvXW2cfgnM13x
WkRaUPB1iVC0+icE3bR/jVBI/UuexmvgPHBoGcIcTtcJBQ+WDyo3Ssi9WGViwMZK
OppDjw4jM1GT5P653rwyVa/Vv+xEexMZoqeaB2JMLYpHHbJr/Tsnja0wWPAWvLwm
rgmzGj8b2F8awsavXrbljRkcUMKjasKjE6+ulb9C5GPpGqyiAPVl9ZWVvkjcFa7J
bc9xq/YO4yT7k18PU6mq2kRYV7RO21A7Pjz+Oa/vfFkWsEmHAoc1N45/+Fve8zm2
wom9mu/4LB53k/5MpKjnuaJ1J85V+wuCo4aZaKZ6K4RmUdW5X/2SJSKzHUY+0dQi
e7BGUXLgCr2Q69/1DoEG0B3L1oI2armzG2NpuAYkMWBKqZuQnLKMXaPlyLhJaojL
SB4H3XCUIFX4MzIVGStDXCtCf4nvtjKhLfl+O/i3F+UWWNqwLO+L9UA1/XAJShgs
KO5aJhum4M1Yje7KsafqvKPPOBHPdGa78tC2hTMKNMZCQlZZbb/LNJPWewWayzBc
s9IOSdMzdXo4C0fQnFIPqmXYiUMLrZ/LH/7je5lDfpqg0aPMOcSTePRl+ohQan9z
F0J4xMXT03bxxBLfBNXVivU+744eKvB6I4cyOCa/tVc5dTjC4fQvTy00ELXK81/k
Gv/fkES2FIuh2JP3m5KNPV5/wQj4/GMl/jcsI0XnYPdqAUTg68o9FyWJfxHuluD5
BWCZBIXckmQTNk8A22hNHVBGVm4gMx5x9ZuCQmCt5DQIm+oi5SzwpaRX70pL4ISD
0aon6UtIb8ReLnSWC53tN3Gj++dNFpyViIgoiubSEQ4TrdLC0r7F1XCxJv9FDNUk
lBjSTNoUQf5dAe57Gkv2q2/D9qj1+sXFpUgLd9rMYMbuknA8L6R1ePsJpZkYRfM5
Iy/tcia11Od8kXXOVZnOyQ+kX11+lJw9i3PCpub/zoH7aXK/SzcHDGYsc6bpgjsm
57xD7s/VeSYjeZgEJ7q7g/meDIN+OWV6FdELEf/2ehFtAX70bkJJECWof5wxOWU2
yIzqdk6zKS4kVkMha5xBCNJNxkYdM1lhzV111B/yf+GJ7jesx79SIRJwhQnq5JYe
Wtlwa6aMZUuuqReCpuUFt16PtXRK8ukgHWgNbwtj60wgjbs7TMyopjKTUEcOWY+C
f6xtPtyKkcX3Alz9VSwkbhs+AXmfoUEQ0Q5fF1/WRl0Hla48Qm5+nlg0et4HfQet
JIhj7sZu7Lq1dTZYViI+rJ1c/+yHTGRzJOqCZvRJ6RPKTU582AO8jn7WW8NcpbMo
Sy4M1kNxulr2ny2BsgdG1j8p6Q0Qi4SYIBiH9NSXWK9cbXdQc0rdzzBP2EzRHkis
6gCr540h7xdNmRwYdTLrZ4cNG4PZCt6MbRZ0wNtkIKPpqf/d+aW4DXiKnIInZCO5
tPpCsoCNysOgdC19juxSUqqUwxABP4Fw3z11cxnYnT4xhLCo3QLCs4RgkisGrZ7H
mSZcqjFkbMMrolQ4cLnD2gz82NIDc89hbwP2+GljSlTo0wb/tjH6F03j7Mk10Iz8
tPjWXuM47RHPiIEMFyRZi059P9yPeuYZcYxMzlBSMaBY9Y3gDh7949XD0ZIWuLRM
MEAOApEMdhnt6+z+YrMHtrCpCCTgZ/tz1tmm/TAZ/DF16SbP/IT2AhvK0vu/PRan
K7Q2TgNaWvc82PwbkpJ/uJR8K3YIPyDI+rpL3HWpYHyhWXt9CwmzRtrbOI+bw94R
XuNe9K+ckY6w9yzp+W7XSHP2EX0xrp0A9Smu2Bh+T2mr3QgNINBYoyfsMbeGpqW5
zGHgB90+GFlDJWPUBlgBGNVUG8vfp0XE8lGEr1ty9ZOfzlLwAZRQXg4LTb07xpS8
zyQq4wqOw3wjdj0OWfW80OUxjI+JXtz+KzC5lY6VdPm/2iS2qhV+C7jixTLMGxjD
dJw4pznNuDf7h12aycTpU4ZC/t4SpyWV3X3Disqs3dNA00E1AY/AxDDqyQWy0lmM
SzP11/nQ5ek4O+n7RDk+sz3c+aYsuGQrYubKzFcTO7Ni5BmXsriz6H3lVFb+Uqio
MxBDEEDicDvdfOUo/eqvUO7oZt9nmtOHtpAVEl+wIypA3Z+fXsg+Dw2z2yMBjRUo
nKy3DVO171ZE+R9x36UKf19G4gMXXSWj+fpsm4dr2YBKuK8UURYyv/+xs8S5dIBm
bWPd+HlaZ9GgIjj1eNliXgYP7q+dteEf+Z3NDi2awFzwg0ojmgDK4fnFG0IIZYc3
rI5+65SeJWqFGA2ehi7rkeVDcfDk4FHWXMUBYYRjmsHbWCFBPOK9yakTtX3EQcy/
BVyQFD8bFUJRTDpzNXOmV5tvyycAMb6bLqHG+vZyCdaxoKIUaxliqQN/4wy6HGvK
mOKoAEvw/9/f1vkv6cnggeXEH4kKHxjA7esxxKskKd9VfscbilYZXLrTrSfQpJxH
JBJ/WCoc0DN+YLqT4wDrc8/qK+Zy6QlPygY8T58OrtlUZ0Pbqy+VyKwa0Te1gc+q
s9tj3Fl+YxY6Z/tuboRXb6XEdaKolt1ep9dDvMMmHHrhwgCrZxsVUxWPKvp0R76f
LjtVXNi3eKPg+Vzl+lBhZJhpNkxLgabapW4s9R6h2S9HEArIlPf5knw6EorUgyoz
UB+3++LG430Wr3UycN7PV9NhmP++OHpMbbpBgQ6096YFbqFGq/Qm7UBfl4Cs7+2y
+dGpk3FEwRyJwhx0tip9eJm1YPxV3ZVQm9uEhRFnUWlWDMjSWiYBgGd61/Rdwdso
ff8NcZR/VbQ/xpqH69eiyvFMQ/IjT1Xnu/JgjzzzrHyu7fqVkXn5Ki0QO6pCd1QT
intQLtRZpPS/KzEb4p6b+aXpq3ZhuMnWYU5cRh4dU2pJ8B22ZaOlALFAtj768INC
rFy9feEearjfeu9b1Y8zJj0qUrrhO7WoOHIFJgK9yWGcUj8cNwgLHRSEBSBqBCNe
UwPSqnwjiAIsrqgoqAeo6GjPDXntq/dWNZAQV1JreioAtZHvB1Fjjg6GbwXQ47Le
FkRmoO3J5YtVSFDIhCwI9iL9NZLIJjvqC4LrqSACAwYruOStF8UuV7D728F8CXaf
GIhwknIpa9I2txNc3DVOmVHJM3SOZrc8FKa+Eo8xJicXZEFNuAB/tjwxevn04v8d
x6Uq6HKgWeuMd7wt2W+ye7HPvU0gSoosHTZZc/tO/NcFR3XvXK8M/sscealmeZRz
FPX6gbiXP2Dy1wGTWr7WtKx8isQ18NlEhEKWepfh6eUr4cnaJWeMfeEus4tCGz09
cGZGqoSsQjIuNet9VQ8NdY+7p3jY5SDiQkj61k2K8RF0nR1ohwEsctNLjKSxupmp
c1WDQOSg/hJszEStAxhHiITbimuHaeiazysfFRSYwLfPNadyRI+U08j3hBzhSIJS
h+r9LyxJwWPAz9duBfUNDkOWxKZ/GiSyP0v+ZBuwpzB/mfzjROxfdVVp3Z72+Ewh
lvSGgEkHKjiwQYH1J+q4tHpNboDMzH029zVu63TFESCO1ANb1mAjQsVPdQlpD/H+
gseF0wBwPKlv5S79Y4/8jiQRiBrK9aomthwYztnxupOVEPj8BXUFFb/M4Gn0J1+T
fukth+zfsWEFGN+HQnNNjm5M0bYBx01AABNlzwMX8PCmDSG520IW0vJcf5v/Fyuj
1gq6hVX2bX8iA/YAIwMNMG1OdJGzzhV45ejn7aXeNXUS9k5GZB3ZseF25MGRDkvY
287d6li6cXJoHdWPuAR4k751fYfBD2aBk1COTRGRcI62ghZqIap/jKg135D06RBL
hRPVbPuH06wN7+QDmMW4xDsX0wqZ4y5KX6I6QT4lKhn1LcL6sgNtHd42YlfuFUmW
F+MVfU/Zk07mTOtztQp1wFI4v2poawVKKCie1tDQWxkf8lrS7itNENHviZpaXRv7
3twO+zXdzVsD5l+tioSkE4aOFbvhXys76c7rOh7CwwD5zfVgpr7IAAOYAEozowWQ
oRCyPzAS4emNzOPvQUGET8F6xisn2mDobyooTMCf1FGzA83oL53CIYK3rIeYwOhu
haI8JyajkTyC0Zjda9GhWuE2tcBir1+x5DM6LvkLLCBwLE40z5x6Q/t/V9T3H6q5
cjRRn3nS60gkQYOtTh6dQIkUULg4MkOXie94CpXnDC2aQbsP932EroeH4TsL1X04
MRxIaR5YVeCtQYdQXpjXrRv9pdh4zHwREPgHS0deABAqq0+x8GRXL8EWPCNzN19V
LWW8qWinvFT1UNdnkm/MCcVKZ6GRBstelRwNRsQUZmpGTC6BUdYlhAzWgM6QHkg7
X/qLCWcAFJNsSS8Rl6Bv5Jwj6sTzETy95O+lPTuEb1hQs85ywYnlwezkjPZ+Ycin
abZOJh7wrKWWyiOlr5DSZVqNdvvTn0pobA/J2eAz6yOwiT5I63Icc1O549FIuWQ7
5N2zR1bgr1ATg+fvJz/gkrZkralDV67fmynS4a020w5ReKnw/Ux8nJE+ubL1uFt6
6xgVMOQK5dL4eXVvdkLj/6PXKcu/zoDRGmoGxcT3oolH/tPpOSJvdmAYpYAW59r4
cWgaQ2xClXFPp1OBde/+ln2M53WpjzBVUJwlsI19cAcC55lT5LnVPJPnfiAukH+a
JDOHy8P+n/OBF6no763xUyvo62I2qQhnqYutk2j+2zb6v2dQ9zCmN4eNpWZ1nmmP
wLnS+Jo4tId2QhwY1Hu+JASwR4iU2do978wILAzr5JpfofCRcPiVtnENTSpVNsuT
w4TQ4ZYZCsNCENZ5w2cRw347ffJbS7h1Ik8KJYu5H5HlNNRubMgZstV74LDLjAIN
rzxMRkayfSzPRblkQbo5oj6p1jKSSj6aNTkf2rd3Q3XodWkjLcSrrx5QXr5f590Y
w33yCnqFmM641h+unj4MfeB1eItjjSXkazVLxKY9N+p8/whgk20YJA3pYXZ/HwL/
AgdbLtfd++3IxCOq7ieQL+H+B8ZmjgsDJY1JjJE2+qFH5BOnnUBgNcCtfytxWeAN
4ccUO2+XQLD6S5KYXB1uh6Gh43XUX/h9LmrYJohQZTvBmcZMrvFv9UfP6Ycinwzj
2HdiDcC0xO4SFyGZY046+oJvqAfehCM8Tm4U5oNJDgB3RcMbuNuAhXO4MYOZn14j
41ZvDXe39If7A2FrEi1q8txJsxFEH0Hwcq1jDmc2xcQA8bO4e7pIMRB9W7wj+apj
/1b5wHN++BCGHwxpSpGqh9nyC+0anZzYeuMDykS7XAVxl1tiKBSkvveMbNLbYvNS
HwusTEKfACB3rKh4NkySxPutfstcywyJoip9FeDW37VrwyrmQk4chhYYmtB9l7j9
hYyAOjafKAJnxQcZGK4qBgewrDxiLmBl6slnBz4i4l2bJ6xsigBMgFqvhqp2Bzn6
mu5EnMtisqwosEfbrZHfIhsk3zP1z1FsrsK+rfVGtKOOnL6xsR9BKpNmSR8pPTGk
aPzE8JIDwQR9yKa2sA1hqG+9NxKlXeeE53ncFBIQRXeLsep8/NmTTweQRngLiquk
SRRZvFX3SdPbeC1/XiyQUO191A4gO/vsCKADMm4VAOvCawcNBuoCFweFrHk2ddex
gJ38iZ/Yqp9fPlpU2y7jnB+CFYsP1vtMHYHcKzyVV1xFxGJOH9IEs0cnUL6Ivyzq
RHac76U9YCWih380s0KPd8hzjQ9nSsG0KGU21R8iCIwV2f2+MD8nJk6krwpQp/EQ
Ld8Myk1Sjc9di5vaOXL+EqJJUjK3ncc6bILAyKwH8E4hjCYShEnb8ZYzlTw4QqCf
vTJQINdkhiVkTRzV6mB/PwArHz0+OLxKVftvhIY3F5w0d1EVSqZXr0G1jYjBSpHC
15zWIK+fQd5DgdBFZH9UHgqDkortMALESKUqvfAlXadNWPr7+qTVPI7NwcYYlkIP
fwPD8EYnbPpQ+3ha7KQZ2fxnTdFQ0fVR6xWpjqZXsq8Et3mjFdnpyidaI6cr9Ikg
q3AsP6TOfTJrLcI7BA3FstqS4tcrR4zkz3Gv9ZxdTQMtpFgLPjAKvlw3CDwthz3V
Ulu8RyyxgjgrPvp/0QT62scoah+MVaLCsj2We8b6zfi9u4e+vS8tmuYIX+hc0qeR
+vuVAoK2DBh73qw8W6OngV/ziDX8PFx4sa/t38vUfj/QJfsFqqINBH7ix6Z+I2qC
5hD52nU7cw2IKIAIb8IrysURpiqbzllGmI6EshwWhc3+6yxD5ACeDZ2mgX5wEcR0
z0aVPM237YatiNjNeqbreA3+LQ81agFeJD8J9mDoS5POv9RKO/QQTAiaZctqZ6gz
AMGlXP6wN39iyZrUfGfqo+MUrMCwxc3nXVy1C+hBuocuHtYeFo07+J/+04ZaLINf
uCSY5gvV19b1tsc3O/N0nWATpXUgyDzixaSwuQI6DZ+Iahx5j58SuaWoLVhUzawM
pJuEUNvcu/9K1WF68Z4ughHnPtzHp/7/3ougZal1E+oENg1DuJ+yG2e6fL6BRe31
eMFmyXAU16m9ewJB7Kc1H+TcLBYdQntueHpJ6fHetVlIm1Kk9ekiqHzn+v4aysWY
XOAJjtSYDyMcyFECDqWY0aD2tMrcnWKoyW59pKK1tCXGjS31TXYoBkcVYz/wYzNl
TpVAh8A7ZzNN59ROl739fb8ZT5Pe7Og5usBepBS8KEvZyiCLM3oh/q7q/YIY+Azj
UpA7RB0D5DPIRTq4RNkQd5vRmTuSjcqne/8wqCTBjspT72xlLx0lEjXJbU3oiASz
/8oD7c9ChJdrdY0h7F0zir8a/mMZ9gsMCzUntQDXZFnaFgME+268Fokhrj+c/D4E
gMMtivq28Gvpj73LgoHMGpSeMZYeoRQ2dg9ly9jvyD3sDZquMKtHdBIg0EegJ3uY
b3zAqwk5Jea6AdmcPx3Dk9tBH8KWL7pEnsiOQNn/7Y5RuJRjsA7YQsmvWQ5t4pUH
NmEtVumKhHBMTXK1h+nEFT+kr3qVHmbIJrDTCbEEGe+TjCSTzpugz9dJh0bb3Q9D
uNDV7oGeA4XuQoeC3QoobnMKSsAxDGG1NitqVZ9jVA5ufs17wNINd0UPt9shKR9O
XQOLgZ0nrcl+lYt9qWRIJ7wSETywtNaIbAdHrreCYfesszrWmQkGxOzwjyqDYVbo
l+OxelPWbIBOx09ULrdI3RJJHwdDroAh94JMExIOPmivdsXkMjFgBOixnNzHZEqa
XNKkD01bPNEHqo7B4cH5vrK0eY2NgNVqcHYT2U5Mc2kh8oio19qx4aIKY+oRQHyR
pUteR/o7v1QiDyRSgh9wrMpOl8aWcfl38y7vMb3kFPQP7FcqTZsD2p9HH3WmouWG
RUr8Ur8O03qU+c2CI75yGv7CW6K8lXZ2lBSSSk36Zbq7ANeFauAtn3dzNRIqL5Gm
AcFdQkRayhHcECrvKL8v+t9xCaOUZKBvhe4RbVUkpHyB5rAG1+dC7VGOmQOtr5yu
5UoHCj5PlIONo9DsRv23jDq/pYm5lgMAPpu5hqEic24i0NUISViaX/eIDiRSn2wS
ZwA7x2S6a88XHj0fA3RcO5dIQs/5alNME1HUnvFvui6xZhMkxX+Fez5+jukvmyX1
YnPRkgHluoOD87H3JJjFg/84fnGK4tMFscufSqNdkOlBlW81o+Ps4vSbbiPbJB4T
hA9302POzetTAYcajOBvDu29szEKglxY4WLk7j+9vgIc6WIm0hUodDOHuv9IasiT
VSKrBnDQWNR5G1Njmau3KTT3nOREYl+VIgsNcK6xkfD7i+FLpuedoo95pIsRSys4
y6kjLuS5YecDE8Df6PN9GcvJnBCCpsmwpPxkOaBuqMOVhKCp+JuHg5EXRv50aNET
MCkTPQojFlIQgN0sKmNBlCPhn9dxVppdncb3/eMhirD1YxGzmbPQ74IpHubREDnA
kWK3k7IduBlFh0apJtsR8JFnTEtJhygLUFRx2ERCjKA3Jz+BGANHJkq5abl1LAFm
8v3kl5NgxAFZY0zS5hFcvb+gP24e/4dFKggIihN204MW2oemVDafs+3afZAOG17H
ZbzDYXRnjt1FRjFqMO2C+qoEk/PeBDPVAtXZ7MCAPqoCNXumq5T5WHYDD+VasFqo
Votk2cWNUGFyXgS0aQ+i+a+NAFdOqET3FWWb4PYwNG4G8OAZOcGIT9FHYmH/MTKq
Ab5pYuK3YUg/EjRq5FX6uD6xvZ7Fiyx/ZMVra9SeZ5RzWdWY4vra0AF0bV30vEbJ
zDPCa6xQd9Qu5lk4p4z42WtvwKEkwfUD4tv563aCxm7eGMlVO47ziNQkW9d4vUPd
oZO2GU7EJBZj5+Y8dXavjwMQNxeFW9If2/cWnjv5Wk67cJGWjw5HhzraCAs+/D9k
/4d8oqLygEfjG3UYB0wDJaklb4b8s2M7E4g6Ds906mM3HgY8Yxrj+Ihn47HhP3pd
ugT/modLd+8gx+EHfxFTAh72kApXAwddob7WxbzoBMp8Tw+VWyRvFp2s24M/Tn2q
oQ92OoTbNqwwmomchHEuCHTnxxYh74JzVs2Zi9ZjvTMzzq2ahUPhAF9pGGtDMUrQ
3ey3XU2NqE4Vc7FfWNPthQShAZ1PO0hq774p5aeULGavtkttZHouNWg3K6Zb2QBd
jN/HepSn+Nmxy0qN8ENIie2oVQlgyZYwj8SxVCfKwwZD9RD6HNLgy5AP0Xd2JFSK
IQwJoNXbIIoS65lPmqQwXVek56O/neEHyBkDiL1LERSHw1geZLGJmE6fRg0V9/iq
qSGHDKgov4iJQlP8TsEp+IRrD2NGzM0ZctRRFXZxQvxOCIWrxVxAfTUqzqCeGbEK
YvGGT9b74l2YHU3MaSMdUrK0gbUlabzmHHeL1z0dFdeq71VAgmRZy+kIJXvUA5jj
uOMMSRVWfs97QTJ3QHnIcgLKSFfC6PdMD1QttogTGxuZvM18U/ekNUANh+NCKEaw
ooQXg8S//0T/SRU4e0GRcvYXOTzk6k7EZKb92jvJZlzZf8aBHaWfM4F9xc6bmFHg
HuFsUG9CUy8WPEkjIim1cZttFzn7olvE3nJIPDM/AdbD80x3XAJXEiKEGutzJuOh
8lIF3cKCQBNSF/X7WeEnB0Zcn1ojd4ZA75ImrMd74cBlxRQuhOGWhV+Hj+vIh8Pw
5YCH0x42r6pLS9qv2A+q+YPBl0UrUiw8is6b87fUP9XPDw1YmE3CuS/PQzXZVbL0
donDrgwaaWZbtCuDL++Zr/JLyPzv5XOAKJtVK99+3ySJ/QT9ovBvF6OLKcPk7wnG
wLM5beXkYv+EKdEzRDTMLZUmGyTOBOK9iToINVxg9a0cmDR65xRP0Lm9+ITyyWS5
dlDbFGUZj47lj4PGg8pExSNSECqOEsTYnEk6NpfzvGAFP4mjl+NgpgTkb0kL+QRO
YqjVMlikVTYYDkiKKjcDPYcurO1jy6gEXYZdKbQXiZtkv6897zN+rVlPrb40LvFo
s5ZtJx9qDl0Aix6Mz72l3zcNlSmdhWi5V40WEoFP1vySGk8BfPoY0ZoBTVkXXf1+
tSSCKrauJaYtPr5p/oVRDpmGU6nYMw/fjzsU7ejEeR7y4iJSnlAAZHliUtTNZ8zY
T9ZAU26XXwQ2qXvqLZQz2j7P82bwZm2Xf+eyScNAT5XmCXyXr16WWrSn2tafmiuB
TcpYiDQCok79fx8lWu3cQPNgDod5MCfyH8DSsw0MY3Q3T/aPjES3rBaBGybG47/S
viNlQa12u8yZ7exhpwBewBA2SPm9QYtT8Jp0N1PDsepP5t7jkpXyjqIjz8ZEE3Mx
H/d5sXaZTxwKyq9+OBHBcc4FIfaIyiBICB8ZnQz2Z1KlYl2AqUXXaRnskGrcWw8w
u0LtwY1CmzpT5egiHiQDuYk2J51lfPU0h1vILcOQ3sx1UPTc1i+aSq8dqNXyOsvb
2WKtGfkxdBFsd0U3leWszmP+t9XNB3tiXin+ojh36nvHEdeA+vpM7jVw194Mqq1v
vf74VMd9Kkl0g/OuxJsqsdqkoKIgs9vLFLV37b40tDUU6aS7SGqTXtC+EyAoGXzj
faaaSG9wZh6MwDKIFM4IXqEtr3YEspz245XtqkaY9vSHTnhpK/kgZD0zFMag6pJQ
z7SOJ1qxU+QCEKlNJMWY7CTiocDKrgDONZqsw9spwNJHuqYyKRDd+mMRea6sB21/
jKGbngD8YXA1ztC12UxnZg6dYBpnZ61vsX345kkBMkxXV7XHhYd/dseuSatDVC7N
JSYkxPFPKGVlWFc3pZ3U2vrUU9UbxhzcQN6i29Nysn3LHy5BWwyAyih1tMENMN7G
WQav3CXBk9UTA+1IxdpxPTaI1oddD7y016JSi4xBEJwhyp8UjB3yJJwH7Hp9Itqq
Xb//HjuezfG9FsyjquwAl8LHMagMda9PtLyTXwWUgTCrfgWHh+7XWTFyPJnInoPx
IK0caNbz/hfl4APC4lM+dkmt8YJ6JGPcwsOahW94dzlfvZxag+NGlqBkTWyhsifD
5vYwj19iwok/ejSX8+k8T0fwcaVCu6K9x8WUp8qL19/rSyOsRKCPvZG+ZS5FasGv
E0C9zBOXMHzFiC/qWNPmj4fMfDF/7nIPv06AzZ3D2ygkh88xMqYZ99ZpIEXQU2f5
dP/mOy77QHQS3bW1Y8IEKFlHqwac3cKK8zmZTcWrLkMFwt0P0AV0bfT9pivxyds0
XPFv5t+L8nr+Jkho8L5catmqNidDCILhzR/7TK38kZSqb+aSAtcGFBPBnSZ9R52M
zM5Mf75PBJ5wDYyuRcE430fGUh2iYBwN5CLUB4khiknZ+3bbfWolINzrvs7Opb99
vnjr9wgpV31PNBIU4ZJxTMhy+BrGJ+fbYpelG+O8/jemHwoBEoz1X642j/DolVj6
iGzbu4B12NYttIazmvDMhY6/3RZv/n8Ko7uxgCRHVGpu8UJeT7zYguIpDymGH8m3
AEBASEtqBZQk8qQMtcErdlfTNgrYDCqqSl4fUViJs3qAxKt7NOjNceAaMVbDnHAH
h4XVknDvSGlH67iEhQdPKKoey5WxNBckD8HcA7fSuFiuH2O0zwH5k17SfxmYRRH4
tOydNs332ue/LI4mNyEjtOHjg00sOvThtNmqvfdon1qhojbO9S3I4WFXgmQNPP1f
E4YqlxSzH4zskpFmJMuOf33cxqEa4303DaLybUIUQjoyXLTWtHBVs5i5jkbD6cjd
Ul7Vg4Wb5OqblGS7PtHuTO+YOsB1pIY3YMXCC7p/LndKR9dUiXSasxosGWpAK+Mi
EXz0m6rjwEMgGLcJ1aPa+xWn/DgLpaMoCDjf4L2XVOhPtOQmCYx7pQpiBz6s4AGa
rDKRJD8VZV0ryvMjgPZ4Pg4fu9Htf6h0yVcbe6yDNN0cVEfwiU+8eMDv+F42wbOr
5cug4+Tu42EiOrKkNS1l6KxnmM/K0WC+Bp0Ntt576F6USA40PYwGFZXynxWdb+TN
itKTPC58xte4b+19EkV1DmMSSXOuB45kfQqFWZGjg73MFBkSyTfrE0x7th/IkipE
U6avzeylBkkysCpGUH3OiFsY9lz5wOLQO3s9bLO2EO/qAldWyYfMFvAJvEUwMAtU
yMR1Bet3uZiRelkdBPHxhRfDS8bhX9FUEm9Ibe+qBWfLWKXXlO1vkXzF0qw6dxCN
O+tpJiEPzBh90T0TU3exM26LCBmvW+lXA+jc2J+chY20FBrQEuMBpB3yfUxcLNGm
+Dh9L3DRp7F50Wb6yb4d9/YjU8Lmm5q7w4wjTWNCD2XD2c59Vl2ni0PLD8GV1LKx
uWyO+JHBwMQTwjI55hYHRVwr53aEmyGu797NZYN3I7iyW7ypLuWdhf8o4M50mW1L
bASnYm8c815chNXFsaX+GKDfpBXiUyBYdzAZkkeh1KJAIt92vD5EjU5VIDGbZfHz
3s+vwr9YpQjky4VbOMEFGjqZoiv+pnDvUXSXhR4+PDrJ3zrq5gMRww5dpdOdIfBz
s3gcA8JlXhcTvaVWndVq0PTGzRvGGywNDTLtthsKDFwWdEQoevX7JGqFuwh7MyRp
Iv2LTvLApZRUciEUO7LHAy9iD9FfOXkIUR6metlUvyKW8RdZksXWmrXuJzqL2O96
AEL6HXnNJHKmkNJvOJSIxbi3an3Ox0gtYzPtzT9Xzl9j2gf3jYugoydDWBIJbWGh
Jpi8oKV5aLuGGpMRY1reucAO006PBZ+YnBG0ziGJSIGVM05o6WyP4MhOlZcz3vfA
2aBr1hWthWr9shWgctYSFaGYIxACGLBWB5PqcX17qBEE8gXGjmL5NDAsMnXBXOtU
jqFZeSVdHnI357U4XthSAFoIH0pwxTvU/qxJZ+y5jj+e3uvpzBYU9mciUx4cUxbu
b1PjJy/enWEPfZYPo4daTb2DVJiERgwDPHZyYQ7Y3K2KHTpO5wMlkMuPcXAE1Lf+
ITbYqKspsSkRsIkL3fS0LwfztrTTHXC+kzrNde2nZdPum7Kl7BxWzvQLXGEPfUUx
Ygu4W0QNG1CXjRsHiJnu2zS4mMwPQUiFhtT+pAvtltJ/OJ178ZSUX+6seUFmjhFO
2lAacS6MD+SkDeXOP/3Xt9z71GBjjrLZ/aNLTOpS8kpU4YNZLdtu7r2fVaxKiDGo
3s6Pnm5Jgowe0N7HSP9ophaHkNebulu4a3NGUotf+JTIemJCsoJp9GbVXwce+MQc
6z98QespvUsX9Wm7FGRcmlSzv0+wqDkrK+T0OsJYygWJo+TlV13NoysemQx6ME/h
nq5oXmNWcNKyZUx8Yy8Wkk6rSOSObhlF2A3FmKxYC4ERcM5kmykzmuMkbnlMKY9l
eGbZfVZyt8XA9CAwbY5bEI53gQ/2hLDuh3AnBC54dpNtEwc/WBoXN+74lA0twjof
1N8oouOsuAgSDv/VnIs5aqiHip3L6dlWw4ovUXDvsbBrS0+8YHKI2fLwPhb8eKDV
293bUqtajZn44SK6gWPKuwmhvkVpsCc6UJ8z0HKgWbo6TaK/WwbTCAfQx2/Mt7Q+
/RT2z6F1c5b5bhhMmwug9RZU4x3lpZ4MU/goUF+0ozBVcnsVR9SrWK4Cb7CK983t
0Y2TjFaP3xDypKZ+g2GJ5NVIl6m9Ss5vEbWrihgTUlcLWzvHd6zWamYauN+BJcBh
Httco0onxPMDDBNhrSOiu4B9txX/34kZnLStvPsYgZyWm+BqicXXz0RC5WJ1XaN0
8m/lYxccZKWWrGcB4RCQRyU9IEsSNGLt4AMiuOCViNeDxWbCVDvofjmnADHDXvIN
5YPkMRu/Arr15RC5Fq4omXSKX/XiyLZA5sdrwddszodQ/ZBcpcP+rIvNKQ+y0fVZ
jERNrKGHlea6puzKTrsDvbURk0bp971jCMZcAhTL81JafQzfaSaj9t6jXlkG6Kq6
LJztdIAUbFZroPH6+D+hzbUPZWBC4dmDzPcTBJCPFZTFjkrsiV5w0zB+cPq7fIaw
Py96+rPUHsOFodN1czVCsTegZtjQhu9JsXL6WMUOGhmNb/wz0G+Z1OiXOq66+V4R
/00b9Cf+Tljm4etFGA6eRpUMFFMnsA8j52BVp1qQYWHDeAz0lsysCbxCU8FgfyXY
MzY2N4XAYoAl5TwZpd7irwtA/BWoWVS4iulLPjEYUX43O6qBytrwk8PP40V6pxbU
oz64hKJb6+VPBAJUKDYmhjUZP9OBxUSvEWfjXMYlDt3KZQx9wAf6AZEPS68xXjqS
2wzF3NYVR/t5+aR479to/gDYXH8qWhOC78K2WMVjyM4cpxzp6hG3vmt4/ESnhgOG
JXRnV3xpiLL9SxoPxf3b1VkIGFgRL78MTEZRwUGRYQ5QKs4Frc3jI2mCchQ52mDb
w6Uw3asNhv0f2vd2eNPTtVESQIZZowtqe/ItoFtYksmxg7jVAeFfsdS6g6tOXTfz
Nehuy1T27XFFHDiXppo3PI/+VawndPTW9+HIv6AWkBV4MnIeRsOtBOr5w1++sg1V
kJd2YuqB2UkxVI32gOzAsFtvTos00KyeemO8/4AIa6tZ3fPQ0HNaBN9O9ePSCpV2
2jaGqHwwg40RBR8YonxW9TXPqAPix/K3aAOBhgqGk0pn9A4bvSZKKFWx4x2trQcb
iVzRBOWDTx1188gfurK5LAD1fWdBzPg9qwKa2CKwiQgZMvVjrDAa59wgGheQ7msV
NAaeWza3we+HA43gSTHuTaWj1VeHzWmnL53YtFnvJog3UGbHiJIUQXTLdKtaJtJq
c+m09sdrsxxM0rOwLtxgonqGArTIRQ2Zc43u58FRJ4zLiNK6vEy60iEQr1iZMn7f
gPIhtRE3luVxYo5DPts7PLiLdr4/mtifCa1WZorya4ZlgQ8PwgYIz98k+dquifFV
HePr7Zt0ZBKzrALsous1Q/+Xs5GCONxJhMd91Rdu11IP427Vbyq30pOArwgCoo+z
WND7Ad/xllBopUNUvH6bBFuCO5idum2FqP//ZoTcUxcUgBwoOj9cDSM/rdjfX889
2ZwYF68gNh47mJip4fO5//w3odO+vn3igl0m7/BfPx/lnits47TZbk9Oh2mvuoVV
WtyDpOo0pVrwsPITuehQko5ALd0M0NHfIlWz62iTpMrHk01LCUf02yE3n/BhPzSO
VFUplFELfiGlmodUgilq0fPvk2pYO9d1U34bWGHUKq7PpOcxhZbnJUTmhpyPeD6x
SkT8PrW6rY1cRsekYdzV/DLzK7pQHftDxhuzw6+3vIZ8xqO4Dn7wwbvr/vV1W6lF
Qtj3Dj2CXYWQFNlpzNqoiP82ELPnz5g0z5L26OCeV5ncXunQnH0Js7FBReKrxPu5
5A/7m9sZ+H4fNhYsptQzjd42Qh/Q3HZrYBH7pptl1dyU/KrjxkwarhbH+ygU4Smh
9fsc14+8k07MmpSWQwGvonTPuVHeaEewmUL77/CW3qJC+OzyIg3P9wB6+cjiNTBL
aLZyE0Fj4nhti17RliY5BldVbXSE0AVB9x3i/toWK91tEe1HRU4pP4ablyDl0nD+
+mFMXqRLsoe1FMsBh6J/dXyM+MfKGAsb/AsN9cEHCq0XjodDbWk+ZH+xx4cyWM6n
IY5nIFcIMb5sbeXzdJyFLluFVL33k68GqbUytFWESKcl04OSTQD7KDw2zImoSFkP
RT08PR0Grsa8GBpedJQM+XP+wBXN4KdRSn47+2W9MRtz4PFi5b2q5/NgssoeEOTa
2N1NICc66BDD9Qy+6ngOFwMX3Zji9pbdbhlul32KZOn2ZzFK7CDDix+mWbQihQbO
swbgqH/2WChn6W6+3Z97bXHYKEkoIPR+gO6mn2J1P26pOEu1iiyQMl2zq3kOsVkx
M35WYhiNJDrxg3Tjx6Lu2cgiXEDuoKlqApX/GnFUEqajbSh37OZ6u7xLEDj4FAvz
7nuWM9DAfqpXETRIq2sszR5Pa4g+w99OE4HLaFO+JDvIvZS0jCl6r6jppis6o2f8
vjVKUDR3gIeGztAwf5pNjJD6P0YQtPYAgWNZcMzsAkXv1ET/rJFyx/+p37zHsLS+
uZxQV7kTPun7Rl2XVr82Z9TVAZOH9H9WpdIXjAnQBPWmBeNCt/7K6zBBKIGQu6qa
Mpopig1aIpNNqnJLVWAAZOJPB2tu463/7JjnEI0Dlg2fwBS0v28C9vwU/7wKpEJZ
Fdt12x02EjEVJ/wWHeRfeQyonVkbcqVCZyOAAtgLjwX+NvWrivNkyzXkk9JIESRy
ReVxAkDtFGxl3H6iq8DFR5QykrMHrxLZHSIYWRF3gKBVrUsCLNqqzonXrP4eRoxk
HMqPkuQqfMeABLzJWJRRtWZcnDUibifQO1B9IFK6WwqdzIpAZgrL9mocckGC26m4
qJa2qhSwxh+LUxVZbTyPTEOKflLbd7TGhKCaBGTGnL+e2U1BXQ+QjsngJZy4XxWF
e7jauXmuaAmG59vknCbKebduqynHg7hlOqCSboKvxbEuqeB/AGt8NQ1hmG+mos3f
CW5U/5gFh5ZYdrcmhL9z5sjdQLXf4BFdNxw2Wh++vNeWYLOiRFSazgV9MlDqb+Gk
w7jQUpNFTnU1ZltoQeZVc9rxhmrhtsBG8HsqMWokkgrBvNsEv2L8+vdGJ7HBsNOG
dmvefOIBAXugN+Dv5jFhvEMR0L7VaE+1D0sM4oBEmM0Wq4biCLztBgC+Q3NNJmgh
pCwyOJoKK6Lya3lTVoaM1dPHPS2Se50I9R2FIhfaaBWloOdXxebOd7/ad3mwb4yW
v86eZgkQEwA5KPsvxvwvEpQbu57xD1IFZvedtBM45Gc2iHtRXjYhrs6XWd49jhwB
MGlE3dCk0FOcQTRsnncjTHC4Jcl8llJaAAK9Cy+0qFqB6gdJAz5CzDpVJlJT6L4e
qQQ5wfAZbvdpLahyq5qYsMoV4sikZF6OYxf5f+KIqFpTodUpOwrGeovxxluvx/MV
4mgVZN2Ho7nwEhKYJtsiCR4DRmMGckjfMBWpLHcpBhHtI4LBVCqfr/Ubukbgr49L
u5r/tSUlpALaauN5OM1L94462QNSPsw+qeKwNdTr8fx0a64a8YP/s9to5JyHY+/l
O2ErUtT03sM5vxfEnj3Wz41RqRfnP61zbgOnuSGyo9Mz2z78IfS9ibs7pqQ8QwDz
czBrznuPjt75/Sz3UcIiQnAciWxXqvEwLeotisnCJfnA7pWRo6Jko/i0QFHpoEhh
OAsWcNHVy47XPuANdZwH4Yvn48iXzsw44epAoLcZ91gK4EfhtSV1lIZWOLXGhuQ6
o/k6J5F6DcGslsncxkzYR2fFuig8B8+A576bivDI5MNd83xaqj2TGjKgd1mv8wDI
YB8UB9gcwQYQ+y1ZW6edqyppX5ESoFNOdkI+PQnNVOkmWd2Pym0fyu0y5+JALGPL
QlJMrttascjS5lb3/Gr/vLquHwXGztBCzUOOm986uhR4rfIG8EuHZAXtICNbpKvl
6ZzT8AFUK5cLo2QGNlUmT3QhFvG2tkuQSSSUML7abNF4oFiNQo9Px6q2CAPQtNSZ
jZj3TaFeU6SHqSmUX3PIkmcrJHEcNSPQnV2oTHBE9r8j4Pk3MPtCO7VTG43C1o/b
hKM9aJY6CyJNqzY2jVdgIqpLgOiHJQrpbWrme9upPEiewZuwtrHdqPS+WtP4gBqw
AZ9r0sPCBHTfaRjfsiWVc7/GuBqAsRpTBLah/0SuFyuihbF1KgR2A2e3xUkGbqu6
FPcOQeOcstKGVmx5DX0I+bf59rWG/yzw2ikijNk4pvRzvmHs/4waVoISeayayJEP
FreH9TIfH9pAwa9Z5ErG8+1PNHDNMKZCH5ZqLmM2vRuWzPCwtp4GcS56zqLTGDcX
QcD74CHlr4gsJVuZIt4aBQXgCmgbLvEAOL7X7evQXY/Wex4sYSNFhdbKgjtkxE6q
s4Ux49KYouyuGsgEboElUqjsZ7vxbYSs7sBtf/m9NovLX6FtH08DLkZj/bsh7ASZ
LOHDFJQQFpbtHobQC+UV5RyjrCZwRfnq5aHvJ+UkDGZpHqeKZfydoIIRhKOhdRHM
bZnFp+T/qJen6QXJyW9/TmPCKIaXXmlDh3R1PlTxq8EwvO2oKhOAKinLWbtn5Odn
9xXWs2gKafMZjkW/BS4p0aZLdi1X4d5zHAghskz5leA=
`protect END_PROTECTED
