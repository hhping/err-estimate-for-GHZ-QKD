`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ehTyKv71JHkBdDPak7IHTFGttRca2r2GFr3VUKh29ephb2wujC/HAvPy/xpq6LJI
FaAGBD6qQFEuLr39P9ifyKB6+kwPEDbULiI55NIjXG3jA5QFHQti8aKUeHbd3Lot
ClQyKTodToe7WMkiL+0AMPf8aIxwVqrQvj+feNo7/G0G5WbSVs8oPTgFW927qlR1
bjpqootiUyMaIq91TB7wn5wURZ5B9j4On8Eu8osMoyMnRNFqTGQ8MXMNr/2fgOsP
o5VNmPDrW1fZDiK2O0Fb46gzEqDrHlhRatfs0+tPOxYtqmPJFrm9XiCtnJN0qI3r
9ejJ762R//e2/mHbJKaput4GqGTlbqsqLx5lhUG/rd9nNw+dBRhcUNUHWVSVQUFa
wkvo+hzKDqAW+1LylObJ5ZddEflgIfia5O7KO1HbKIEG/G/y6pFbtHtUNHRnqgYy
iF3CMC3JKMu4BxaBiwEVQ0mm7feRoYIDVD64nKiPMhDa2HZYnWAti8vxZ6eiZtlz
OllxM9NtY+QA/zrzxin3KVYVAo+4RWW7n8eSEfct5GlIMqn+uFPNZQAB5HxqS9de
5IaeqIjAfbR+0tAJC+2z8DYdjCXw/bsLq6HTQgalpjgGc3KVJhcfPtzPCqfc4njJ
KVV4BOfFFNKnqYKGV4I68buk6zaYvJykbcHhSgZfAQ6kT/zJjJfrBtMAjU6cx13z
AZ4jH1Pl+DtEnUp0zRQEMRkaQ8U5U6gsOTuxmx3XGrp8vYQMZK7WtqDGAzLsW5Pt
yhdv2pdUsJQWiOiyW/sRaOYoSqdSS+AyVPUadHcy2JttNCZtirQTcmJrd6Rz/5iO
`protect END_PROTECTED
