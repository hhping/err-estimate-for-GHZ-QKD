`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qg7vWx/a7K2GXqKzzJiesXaBVpvyY5pllu/QPPjN+czqJyevaGL9CHuJAMB1EWTO
xlM4bS+Yn8AIwMcZriFdIhn6V5OGVdqoW9C86x+uP25HRA25adoBf3pSuT6JNLPz
gaarJhpwylkbVcekWWcu4lRMWfx8a8LP04HDbP7gWfLKuXe0gzVl6jB4ndc1js9x
x5/B+ZLlhzp3ohlb2OAPb0SObFcYtoloviaXr5CXF4bqT3mIeYwhTMQ4mkRQK+Vo
qYeX2JJBHSmcO68s+SIqTofZosCtO5UkHlsUSVctgoulh44+cF+WkLEtOlRxvEBR
sHH4lC9UN/zqDo5vCUXZ2L9r5Zy6Jo2lWHId46PsJzndkSvT4rb+zO+d1Fe+hnZG
4SoRkkr1yrvCSFzXGDfZ91dURWTZRUsWnpZx6R10GOSswTvLTWGMhTnuWQ9cbvsq
pJJP/+z3gs1pkFdg79+j36htFksJtkP8EyfKTc/S3f9jMgkEjV9IIzfTbk5hR7ae
OP+DYsbFIzZUCd19KdTsUIke50TfpEsF6b8eZGG/kZYj7oCsEWp0PuEUCqZcKmq2
77pQ91XpmgH5OGIoADklrxQ6noGHdvqLAIQZlf6pmOGfUf7XmcUKqs5vOb2m8nfr
oHDmf/IYZpq+mrcWm0iFBcKG+mtFKTmsfT4BZ2o0CI8=
`protect END_PROTECTED
