`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RwPbxXNqLSKoDAonJVoKF3Aj/UcqRsbd43Rml0WMVbz04Muyd6auHLsquwKVLlTQ
6xyDMTYbkkogFYdtUgYy/uOLwF2xTBRC2o6OEbsVBjCHaLBAsZjsBsV2nf7I1x6k
aOObfHUe0dUMy1DpmNtPsW4thCa6TN/7Jqvhf6/mFTwY4DpUeXRE3qa42PsPzQbC
RKJ1HJ4nlZgztAy5XyAc5GdybByms3/uvyrGAb1/Xwp9owEOwzMfvuWdvEcDS6DT
glQbkJbY6Vnrzh6XzQuBhuMc/uIkpL6/zjgcVl+Vm5fuhJQsJLLqD8qEVu6Pk/21
CSvksC/9NsLWrj4cfbboxKZYt4dCkDIpZyyBz61VuZV0kvBVWuL+nb/P2IyuU1Hu
1b33/4dHu6MNF4teHcUBQxZfLqXuoOEDrhaybJyHtPHFN5cEhnPK+MoNaTjUnDJk
qq+fwOA0bJE6jwVZWUbQWRLp+qyZenVlWMEwSu6ICw5de6Dakp5b68WrEy3jfZhv
c0xj10SjA+ARtTbWM9k4JCArxEgPjAwJ7gwMz1i1/A4lrSk0AjgJG9aqH+nnMrgu
DZ3qQ3A/+JQmkjJGawNFxmKgXeOz75WsnYFK/VhKdEqmvOddsGBZA/Fo1wg1Tkl3
pCNHaaYm5b5qBCjL74DFWQqsW6lnWf1KxbgizjJXFMsAEjAnaO11misjjfpKYukb
lJ8Wxy0+uJhF6cryAWfGDTm6TLTVmyRV9Ev0s52eWYMZIHSF+svH2K/fx2rhlVvy
Y5pNWeNbpuT4uQBRtPDmoUZJgLMtZsJ2wT6R2uWsaAY=
`protect END_PROTECTED
