`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y8+6UbEhsVha8GiIiW3cK6iDzpL8UH1tmwaKAT5zqk33D/vLe+I28JvOH1r9lGVv
ZOz6Px5MPWtbiv3o6oOFgapKclotW6jLTx9tZcPQrqEhQ5ISl/9zM4NPDpFzOTnq
8VmSZewevIcu+gVNPo+G92bCTZJOAV9ifITPhsC6vTnTEGui2Xlcob1vFjyhGFi+
bDcID58EbSr/ck2eeIrIvSGPIN+u02q04viEbrxauccr4Tg2TCg3gGUkdJOb1fiq
EZfwXWMxV2HrlqOBFmejxJVyMDsiB088Pe4n7MEuUJy1F5AlWsZubMhRO7L5SY1c
9KdVwDAjWstVe04Uw06KvB2g/cokSm3UIFTCXIfa13nnBv3HdINBAuUcIRRhxdH2
TdvYQ/K/ci+2OS1AsLx/xAfBI/li2XV22hHJAk0CjTiyOLLqDIHs9zePcTRhPoHm
0BCnVh96WFRw7RNB8CHHUCgmFfA7xTpLBa967146+dFnYIc+stgrohShzfGGTLW9
AfVV309B2zPsBAHfKYnbhxXeC3u+oi1nexc+jTYL1bKWBpokpQUkplRHCRO1U313
8Htqol5dZ/R2oL+y/2lUWdSqXdb75a2qdCCg05tQHOYmrWx+yWSl8OUxBwmNVvgY
o1UMVGC0I/a0sDRv1uYGGWy5U2CqBA/MDob7iQePQ2qTrhjzGuTQiBebeCMgprq8
GDH0rdTFKG07pHd76XkGfGH/8UYTslBiiBBvlpINzTLL8Nb552eUxHAoInT3BfBA
EHbMnHcptqwp+LpQ6kp469k43juTBgrY7zWpDVd639WjDa633orA2VDAz4Jo2MHy
6XpaHsUQWUEe6rOo5HVK+WJa2MgVSrsCroFFMW22BPT8i9yD3hlm07AB7VKHcZnm
wBFSHLe9xS1A4H0/qg8ihB/ngzp1cbK64kURumqLa8WJ9KAoxCKURQAnKAZ3D69Q
uHCeoFQe3FZtHUY1x6qUN6LTfwWVJ+BoxaPagltRTbz9PqeBpwi/ebNFNgOpDx8A
YsTyb2NSmFdxkXne6zqi9xcwTP5kMbPTcCdeKV9Lai6IiA6WMPZdhF5VX/erGw6f
/64DGkuGK5uSBagGmW7cAXucABUdjD7mqptb/tpa7v9+sBnyFWlY8aEab3c71spQ
6L9H92tEJjPrL6B+YJNpVxeeQ/zigPA8cJb+2p17u036bu8qkYW7yx+QbWLefeAG
Q2iAinWYyrxyl5pQPfCyE86tL0r5OzitjhFKS8YtEBFfmn0kof6buoILG/jm9nm8
L9N9YT50F4/tcm+0Ll/hSjSKIOCTsEri5ddt+NOg+C/M4mz5ig9bBqyE+IW1+A4m
n5k5vmJuJgSGNTIjCFgUZdloQ00t1lfhcULGsqgfXzG5IKmhTLGI2UhYqamM8ESp
oT6vWLNn66I9gl92nq/0losndQEo+nRkxN68Qcd393dTalKJyzHfsy2k7U5EqPoq
01lQyWyueRpHthhzu3s6ixTsLE8OaklQCJOCst7fpno=
`protect END_PROTECTED
