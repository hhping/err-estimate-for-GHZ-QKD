// log2_fun.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module log2_fun (
		input  wire [25:0] a,      //      a.a
		input  wire        areset, // areset.reset
		input  wire        clk,    //    clk.clk
		input  wire [0:0]  en,     //     en.en
		output wire [25:0] q       //      q.q
	);

	log2_fun_altera_fp_functions_161_f7x7wfy fp_functions_0 (
		.clk    (clk),    //    clk.clk
		.areset (areset), // areset.reset
		.en     (en),     //     en.en
		.a      (a),      //      a.a
		.q      (q)       //      q.q
	);

endmodule
