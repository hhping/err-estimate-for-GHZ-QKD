`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r8kNrOqPCvJYp8v1oMnILZ4a7HhzWI7ABmc6LKvPU7L2FmEdLNwgtkWU+1Jcmgbg
NfTYizmMDaEKNTLcxwEzJCkMcTDsAWTGWXoJyIzdNyH2P50QYcTSwiFULclv8UWP
4kBmubSOayLoszsM0t6jqA0758luzota6fJZdPkT92XaDei7C3yy4NYxcDDoyWwG
Ta1hQcwR+ufZ8jI+sLZUozpkT2g27vbj4srV7nPhEWBLTH1Ux/H9AFBY/4yE/lT8
QqMjF2m7Q11Rb/DgtQNY7t/46/41V7HdXN3weS1HSXApRNwPNser6SRxO0xGDdE7
8/q9G6rfKkZQfqXyt4I9fLUnnhLkKhmSL6eMc9a12UZW5sg4jkb9c9J5zbIw9eXz
MEtgoFTQaOdLbXTevWmNV9+MO2CCSwwsOtuaNhcRsxIuFZRpeb8xm+kmX3X4VZFH
Ldf0qmTjl9MZ2k39Eht3/CZRSuFJBnCIcxAayMvD7xL8YMKtwXIZbDSfV+owaaPp
9Dc12ltVpX5PWyPvfGaNn/g9Lbe2nBn4L+tEVeVviXwKKgdpCZ3l04l5YdV76tg1
0Cen2IbVfg+kjewqlgJ6NcoAtVyTr6EePfCXhZw1JYcI5RSRGCmUoYvzSjlQTtOB
pCO7E7b40gOa/k+vxEcU5kcIw5qu9++dUgAO02sv77xVDajF9EsyQYhV2FWiyFnn
+YJd1Z6AChCvWsHUlC+Dy5t4ukkqUwSMSHpzcfoedzn9q3n7uK9hTBiXp7A0IpmG
ewXAcUXi5IoEkCkiGOLGkodLhcw5FA2QfOxSej7mXFEwATuFRgASPNY71q5duC7+
vmsMsyfQIUMxiECWcxRSOVGgVdnnFZ1LiFOMWjj6a7JJ8F8fYNjZoZ5wX733gMHb
ScXhom51D96uja1+h4b2ElPFocPwORID+opacOnHD4GyDFVhctVmz0Y8l0ksy60X
8hlVNVaPAddIzCfUmn33O+2NIJ5NeoTiR2fi0SKVGTs=
`protect END_PROTECTED
