`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CIMN82mu0uCQB9XrRK/b4YU3lduM2wLCtWP8zipfB0YGAKgWrTZFL7KOR8rSReOr
TJSkzXS5PEWSkeQYr6z5Hes0i/cliNnBeZg1Oa88mNidLhQw9YDC+5K3Pc0qI1Va
gGSuLFRGtm3p3iXGNdspAQM8aJwgMWqm6zbzUnLxpMKQmQI90JHgIJmkUp80le2z
EiyMUfwkj1b7C1NF9yxFtcYmcr3IKdtfF67hY8Jdj3mGj9GSvMFrWVh3DX3whXfw
9998TYZZINh57bXFN7YviQhyjk6eKF+e3dBbr3TrMyK2TJyKEp1rN8975T3VOJ6e
fqoRd1E0U5h3P4zfy/gYAfsyv5MH37kIiqynDI/CKiGS10C20nTMN9BlT78Aaqby
edbX3ZSoxlq+1x0m6rJLxUTf1JxLj4etomMzkQW1P8ET0VGAeqm0VU4sdyO4Bjio
BO1s5MHekXmDu11x8OgtHRToPxVnrBWdWq24nPvE9vVXM3U3e4YPi+f4y9DyYVZe
l/MiJyHl6wBcMeQ2rRUBUbnJ4AXpcpc/1aVau4NWC7IWn16SaTaKV9kz+rYYAUxv
MK40gj2ZV+GubMMH8A5hsMrqbjLWmiz/1E+htKmWrMQE20vmk9N+Ap/juCuURSg7
zadMpuZnREni5cDNO9nZxTUjYsKsqDALssVznFqpEQxR3nt91CN/sTTASGmEwi5i
hvmyt7DW/pIbR1IoGRmdn1ioGmXofgQ+EaOeNGrbFOesUlSDUxP4wBfwHIv2oEdC
hFIto/quKfHDHJhtn9Vafrs8j4wE3KzALIxf9O6rgFbM5jTyKzT7y/6Z7SuOe+1S
l4uBuJVaeVMNzdB3HuW+QHgyE2FScsGw/pn7M879WmYZPLvZFItt0lnUMI6qyVxc
0k5p3CdDdzD421g8yHITq6M4DykrJY3MzzRQeZYNYb5ftXalvZABZDgEodNDuEkt
pegYi3ovK4yuq+dJW+mIerLh3AOx4BZkfy8qjY6Bs7Jfoz2HPdSWtpywEaxeljzt
TQP32XicubLPNcbANejudHN+YC/lwIqCKmGrFND7xyBdlIcJAYMx2o5CeyjUyKDA
Myc7N/JgWCCCVQU1ty1kcJOAZDvLGN6Y2PJjXCJrIU04ybFX1wZOeoM+4HiZhH1W
dzXH3ePSvON7W9/f0Nmkl7dopk7gKH8lRRaY9rlcx67+hGtj5dfE2ToOznEEbmwG
8R4pL++Q1KKO9rJcQlZkV/TViUhAMyOUqkFHdFkoZ58puHxjOYCTCcDOUlvH4z8D
2U1gKqzn+cKeGed4zKYOgypK3AmKUnq0YIx0ipJUj+kdnS5tk7h7Ps0AwBhDRuUm
f/EiqvPLimUiYFooFWsdvhxog/TfIhr/q1KtUrz8mYhBZ5gdWceUIOMkHO9hLUi1
YwxzgdocOiqZEJhS6+v+89JIX9mRyA4ymRhudL/cS+fg45DMjkUY+bJTF7FMH/e3
1EK/vZrvGxDJxxoySB35gyPXyd1BqeKHdHt+SYAqsyyRAljT5Y9xSHR3JJG2iwzP
hyxN6UxdrLDhPkwvVyesRLAeI3gGeKSKmcMctVmsWM13cSbrg5qzuIjvux20SICd
ZcnKJJ8BZz6oj14zL9lIlwW50hXAMMJ0GK8NedNVPgw=
`protect END_PROTECTED
