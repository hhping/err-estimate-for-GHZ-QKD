`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PjQJoGGnEfOeu6iog6l/uMKWPiws0uNlno6dej1fU9B1Y85E//uv202o8dvtuIoN
jvTtw2vr/LcY8233UO1MMN+xXa+/3Kle8xHK3zRmYAkBDvlyXcO91j+T92qvbp8k
1vM8xq3RR7zDjhkNDArQ1UY2KN/iM3tUH3ouFBiS8W692xI1Npah72OQp1x4NpEK
IOx7G2oY3VLRKS4V7Nh5ZjYsPlOTjUtAFZBfrIVQs4f7cI9nIxOrTRFJsDpUaVKD
U9KbBlpaNIEs+xUJVeyv8kCRVV7Hcqr3msTcAQqsTnrIg8f7X246M39UECgaSpBo
AaIkiAGD/VWuxfe5I+G/NNLXefbJgas6LdiWbMOBXXlugltaQ4kSXsLWwHVtR7a7
T9AVQMN6vw0RIB+4OmRyQn2f61vSieVMBocqi5kEZwOhj3VKQ2vASCxcxsVdjYBe
6SjGokuL7cQPCZDvcdp3psCn9s/uxq+JFTvG9AZ28GRqKnfFsIiyjKZXTBm8SK+s
zbpIgh8EXEwRbiTRbuyTVjub2aKFPjsKwjCxEQ44LBl4bM170y6YsQ/pTDMlWIgQ
eHk67vUFCMSIyz+tfEVtkaEM/aQiprJJQj0mBmRBm80XL1RvwhJSrf+crgwaSyqh
DM8r5heEK6pxsmXJksN7RmzS6rr7oHmubXvNaxkc+aRIes5TtFW0poxXlwxZK1pk
aoGQYPu8DhoBdIFkiYzu97myJRofW0NLrwjvEez5aG96YzB5k2QvOzfo4gXtBpyB
wwOnI2Bm5cG+FniovgL571UiYuP5Q+uEq9QHLifDApYaJOcAH8YfDIf/OauxOO30
e9EWsOjGpO0CKpdZMDihItPlk8FP8+OIFTo71UEBdQU22AyKpd4K8QOIOIx0Baaj
O3Qv4ilB6XhfmJeg87iet4GlrLePjOKUwkjeERjr07ismX59pY4NRQJyKV4Ps4Q7
k6w630BrN8iwhsDi1A+VZRUVVctT9WXR3rnJ2vuPYL/HX4GHBHr5yGtjz4PqJnuE
JnE0RNPRqgW+j5fYOWraVSQz70ickbF0cvHphEpU8QVqeIY12amGB6GSg07uW8u3
2Z16D6NrFxzpc6Pzx3jTDHjFAf4yOsiM9IZwbozs0m4pYDB1ayfZYg6FAAkKpwau
lUMHBK83nZhKIekFNb9VWzjbpD1pTPKVwSlnPEcFyLDf6ZW+ooRS8W39JBvBl01P
L0qYey5f//86r2QZ8zMe1+27wtN9x61F5tTejqGatdJ1GJGEk4ShB9i5xBUl9PWG
4ptozr8pc3XZgJgMmGBLnw51pKdKuizVtYjjXATsNAiFdEjUUSG0/uMesLILy0+L
e+d9nwxPayca7/PI76NMqATgwgdFWW9sGggf0igXWotweCBtaFyz6DDMW0StyYyJ
`protect END_PROTECTED
