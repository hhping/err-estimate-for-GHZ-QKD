`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EU752zifJM5/Rr1lnFJCbuJNNrWj5DlOJHgaKXWQSnoLPPCPn9SvJnqCCTTvXFSv
bjLBUlSMvhKcfGY1apNZCmOj6Orm0mkYg9bYJ0IgSJ1peT5k2S3Bx3YXlP0YGeOn
YFsTcmljiKKDW/4y0YCb8fUC95WdZ/A63MMPkemBplWAcx5spsgqo6yHTBCPa/Lo
GH0bCUrKJ5nnyUA6HUtVMEjr0rGWyWPVikFTYaQJHGa6dkQq5xvb8ZfmGA4X3PTa
zhpiXX27HFSFHycVzgbjpbT7RtMyD56mN2r48+nBDztvCTKDbiLbSXHwzSZ9/JTB
N13OSXcE3eEpol6iGDvdjuVK3kj5/zaFbpb2hJconJN0mFQWYUwWkA8r6zbW/waN
YvTu0dnIrqXijFIz/6CF+W7/eLPFd0VC0d49x0O6UisBHYXl7cSPkPOcm5HC3gbQ
ks+NE2rmSZSj/cBoX+3/qpVS4PAb6ZOIFF45BtRUwpeGphQCoiYT9sbT2aXV1NoL
TelaP5TtTSww3tJrBcWxdnW1ZqhDVrVEMAKMZr7pPdqFAMyEZS6tNXwma4G/KRKK
1hiW+29Hd2Jkv4eo1uWBj6MhZvHTgDmqkgTAW0l9tbhmav3pd6q0q4/6hfZMWCOw
O2phT2iJNfcf6Jq0m2nCsr39br20ROh5hWkmyIbG7qviYgjzyBX56NjLbrQ71SK5
ItywREfshDqoYoQJbs8mJa2M59bMm+PcwhVjIokEvrPPTJzbFBDQKPbtKejL8Roq
8YntNjkJeu+2HLVndZtSfgx0oDh/aBOntu0ifomwTAi1pweQXsyQH5avmaa070rY
SAvb9jXr1sFJVkvTLH0TS8DVGfAvc7yXJXV5h4jdtrtgeB5XqGPMWyfQeoWylh/v
merM90XHK5YuVZtmX7wD+EbBZ36+CZ8gX0lnd9Gk3kqqITelKo/GahFwAs6TdzbC
05T9cWCKjP3sq73pWHY1hRIVxo5UKx/xazJcUlDQZ5zYu7iinyvR61K/2DBkJq6m
67hSiaV0KVD/r+zaZD6J/VSaD9r4HI9WLayBWLNO58CmM2jrjQbYf1/M6QA3ZFvm
bG1I9YDTXzGpbLMDxo0cWlHaVr23ippJ76CIY0EJMLM0FurWVLrGTMlvBNac5VOP
+WEmDARBQcwr1OLHPkS2qGruOdBKru9HJ3vryKRZOxN4PFVvd9nG8q23/4UsKQmp
HYoybb4sILdd0vVPOrE03LuvX/+jWpJiKTvzRv3aVwr2HpDnvAvvyPGW8kn+ImZr
ehdhpT9zmEC/5xaP7Cz7DuEXLiHHO+ojLXzBY50ltmK9vaXpVCNz3kwSbfZzHG+n
br32Q5IuEONZbEM+UBpH9Dp1EcXFM4SeQDua9zahmdxwc0BE1wJK+CELBGgcrMaW
vgBOwDlvKEvEbnKcZdEodfYmWx7QrTZfgOhNspCrF8eGc77GxflXtvzhkC8iK6xl
a1t92OSDZXe1AMD12ubrcFyCsmnQlm9vcGFHw4inob1I5Elr2s7qmzZlEC5eHUJA
AEP/EGM57HlPuBKKWTyDDaKyFQysWO3QjRD7kuC8psSASehfW9zT5/6nleYF0Dx0
weR+VHiKTsgnxxQn0NC/1VufalUrPa6GWHP9E8nxX4qGKskuWXt3ct0+wm8yarjH
S37FyNV6OAxxWT1HaSCHAg==
`protect END_PROTECTED
