`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zDSXTsQi5oEskIXzo900m+z8ME9QhoBUweZW6c4/WvBl3QnQc5fLA98Uj4Eb2UT1
Str24fTY5tjuojGkmzeNN61FZ8Bof/xKXJlBB84sp9V38hTZX9zIM6Q5+Al7fxfs
9zrZaAsfT1ssddVNeBmhVwCBG9mWTISFahbQ1Z5OoHfAJw1B79Bplu+UOT8h0ORS
93/PwoNnUvD+utt0fNXDMPCDZoGInngJuxWFoNrk2CCoJH1Nyrq3eNK80Lr53/G9
LrSpgGr+ho/cuOyie7vJyfiKe8Xxtwk+qcbCoqLxXmU6pw8wTxveIHh/+hItCDIC
qSjUW1UryKCFvgVU02MEXChS4rhebGekl/UtKRe1Ak744JzzYi4XU3TZ/3iJM5dP
d+7rkU331S3gE7P0PPnOxJ0SnJ4/fPvgeinC04ZNNoXNRb2D9QbnPeqqm90V1Dgo
tcf99Q7VLw2VUaM6BbBShcEfENYJOjcLYNzhHoAkCH1wCJHj9prY9HWOaQyZmdVQ
SAeWeCYmgBXN0R6aqZOcalQD7CuCDGdjyU4H75Z7ePtMkfOje/OzwbzAAY25aOID
V1K6BYXySFIq8UySeH6ZzWSZ0OYLIT/1Au22M1UkBVE5DbXxOjbFxlFNddVw6pwG
1N7PS5TmkDc1KDMT63hZGyDJtYbo7xqsfZwM48bds2UaZuZFdlQEP+oqH1K7mMVu
TNUn7dfe1L00frgYmx/6xEX21YhgNlJYkNLFdjKVJecrZflGyNbx7H8afsIQbqR0
OcLTlxbSgnhjLAeteOjKKoRKFpCtoN/MdZReZxMGECW7Uo+UOxsMB7LyRFyeFPqN
NdR9Q1ECZrHgk90Z8yP+H0pY5cNlvMfYSZJdSdZrtsCRL+a2C5JeNL6z25zjmDNN
o9YfG4UTqNMqslwoVJB8tw2UDV/Q3M+u/E/J0hKYlXs+3qr5paOGeoZKkm6mE4Ro
b3xqK1fAWuH2Mn4lA10mmS9ieA7Tvaor2DOVeorERJg65uhA9NEs6lRaOxICyCv1
drkJjQaO7eyppC012DaJeyrQnQNn6yZj7Z6ujpJLfAz2FNAXdwhlOfCi9NtEirot
lUrIbK9zE8/UkbJQK0jGXgO5pDPl3Xb3sOHOg8gh+B7IH8hqrd0q5W+VANPQ9MfX
WcmK+87QVid8zZW0fOuQFJzpLIz71aUOzC0as3cAvVyyPaBWY3zIBw0hnUui096U
64WHOhyZY4oProtms8IG5cfchtHP+qKaYJiz34ItKhVUr7Xzc+5VL01e9DFoADE6
jvZffqLfEkBcQdPUZmb1i8Cl5rWuAGAKx7DvkaGQj3ywcfBPoa/pPqBqRwz8NmaN
H5KSW4P33itNNDYUZVvT2MNAuQPTgGnyjwF/UgExN1MCxI6RlZkc5NKWE1FKZQWJ
DaPwFi5L+1NFtNZsxb7T0H4S+T9Z2/RxzvPmFHN19ZFEgRjqI/RDKl9QRkUnQSMN
3BiSecGv8CkN0uDgMsTHv9xj+P2Laas3bdLgXyOmzWFt8gaTMVnii8H/CFZQkEuJ
uHQ/jy7Hmrg9ed79vr+FB/347tjH9w2a+neAdWXTVLdP+LXg+u/q8GRvy+kRAmey
KC1WQdKn/yMsiGTH8FDV2n7ndP53W1M6D1iakPRNd7lbyP4FrYTGoZkSVt+Mcwip
vc+v2K6NRuvWTj4ONH63jw+QQ76+C/edMbUAVLB5k6bnIOM+8kJ5WwzfHf6t+1aa
`protect END_PROTECTED
