`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aMfgCrnYI6hzUPrOcvytBG1tmM+x3NDNM//nmtu2iKc9m4SZc804gQRtPspaFkSg
Qoam23BkhEK0HEQVlLLULmTloL6LD4dOdnKCTN3KyCknZ7/nE6hNWWI/T5kkmtDV
mhhV8Avc5/MJEQj7On9x7RnU6dsko7yraV9hLDq3SKR7rS+Kev+d9h1qh6MvhqiS
Hr3gUzzXuuTu1qcpaO1krOaHrvr4vptfWNnn6Vu7Zp2pWb3bPQNoIQJesJ4NFMhQ
lEO3uRcWo4kYgE060gLzVvqmxcuiAaRotRbr8K1rd3V7UWZfSj1Rlm4jB+cLgg7K
vpcCjnKI9ktCyN89oCkJAHKWzwpI1g7lSU8EkqOQlAEYlzIHCbpM9gqvouTevw81
PrXLp7Dm0lFM2CpxlFXwAaMguzZZ4scwPIMblI+opCF4O0gNO+VeXSg8aTJXafpB
tbUYx7TUYp2aeHOIRkO6mp92ozQWpGqLAdCi9t6nwG7Fx4c8ZY6ECokqkpp9g/jx
zGyLbJWVoLDkZ/9SnT/Y9yELd6B8Eg9SznB5ky7VzdTkNZaE0H9zIwirU1000Weo
gSw6u/tI5D9gl32XR7yPOuCiI0H7BiPshlFhozdQP2riNfzD7TJVbeclrX6l2ZyJ
rlBh93nS+ktBeseivPBLcQx4ShpkRfzbIgog2K6D7DCGyv/cH31fTB010NbVlHmn
d5GMFFBrZBuO0NZft7VG9SGq6z84xn//lvfI8gI0MlWyMHa4f6Ns5Zew31RUiH6F
9zd6bAfexMbz0BDvYuLdnocqaJTcLhQ3xU9F351BAzWdGzVIKyyz0J+3v2bqJjEX
o0JT8cBJFrTjdotti4gPUStaOposW0Y52hVZE8U/122lXq0SKM1yu/6gLfDyfRrb
TtrpmkDm4rPTsK+0+Aa4+Gz77l+oOXBMr6XP8Fa1AGViyv9S6CmSSv7CEjIpDe5g
T1V/8x4w9rHrdobgnxDMqRGN9eZrDyVN1zDdtw+N3mdZLDflhGY4hXY+XYRbUxRE
E08Wakc+v0RyGRNJ8v69DV2pZgceeXMcgyv6OjAVNMLtMIQPbr34Ppv1UC5uiqw3
lQCI9bTNtWESqt12E3VKvnm7QFpFIfG24lyCYo0ak+UBabbLmC92/WmCUMPeDmQm
uRoYa0qftECjzBkwijgCEc0QWDNqSNXSFIWJ3Q7H1BMjg3y6QmIGYKeV/rF88A6/
tPfvAdXsGmTNbJRxPViaaQlLT70AOKCFaHbTXFm0w8CfjINkPJCIBAAC83Ujstit
0UzWgnLz+KF4IttiNhqOzY55f07cMNZEwUp5SXo0jgQFLmqpQAqpbm+e1S74n6vM
qIrJ74fUFuMIh626GSsCR/QBTZksBN34/KNgKS0/yw1sF9xoImBviTq014L9kWUE
/O5QPFnWuHlBI5OSGdRGdijNyH4lqLh7HBVcNqqfHPT1rPkXdAUbp5wo5FpcCHA/
+MYHMZ3barrIgZkh2fWX9lXgvw2AYLTWlmmpUZR8MG+wAancuWDmMquKsb8fJHpc
CRmWgWhpc+lOmYqdX+Kq9484ww91zqAzBovH653o6o8=
`protect END_PROTECTED
