`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v1UVj2jORo5tlvb5G6N9ZDrh/2QpR0kpRNYwBi4obwquA4sAGmKq05dQfurQD5yo
MTgwCgyJAkku/H5mD37NhVEh7fuRRPCjR7LSmvgl/goGbD4+czDw4r42f+OQqMsO
V2l1cxIA1HJI1EwzDXfhmJx++ATebavsnqITzwDafWqvwWqeHZCQrBdFBidEGfw9
E0KFCpJoC2DML824YiTlN5N6Eex6pyxo0kfHD+h7opJys00OBrv3yP3I/+csDxqt
+SFoLuyOeQRE1kcon62qa6U6cVaLpWc6qHBCHF/ryejZ8Q0o4AHvEXqD+Pbh9eIf
i+LqNBYM3EADSdKng8GOdPVlSNqalNaenDivYE95JsnhJVcCHEMbJZCariJSgx78
/Qj2NJhKLoKs/aiFQUjQPedOfo0PqMyI0SY1Aw8Y05g1IxUIR2mCxl/3SVihxnop
gSduFqOdicL+E5Bm216MIhtIjlXq+IkJl7UX/tBDTNvOJVKUiSuW2z8RfAdJg/er
u3IYNr+7N6I905nv4mhjBzN3AEoDMBc71ALi0mr/jzNWidRr6wEU5hQRZEfMveXl
b8ccgpO4OmRCrnc/Nk7rg+bljgjFV2bvYK4hU5dtlVmXfA1PTHsTtQ9I4cNMojQt
0trwu8LbBI8eIKJI6E2/wxxjajm8GRdAj8Uy/ayaowImylozu6DNX89f0mDaNDdl
3p+ZvuJ/wbraZHEqbE9y4RwSrBj/JUTjARPuH6nF1UQCUaV6JbmYYO83s8T0pn9Y
yDmc/W2qqsultZRPZscNeijDFeTvnrD2VY2G8sj3sfmLZzwflhFubEu+v+fN3n8U
`protect END_PROTECTED
