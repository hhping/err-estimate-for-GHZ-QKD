`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4QJ5820gY7EvdG/8+9ZOLj+dxyJuRa9yDeoLlcukqGnyWDeginIiIeiJAG6VvgHF
F6mw0IXO2NVN1B8X5MruIG4WHIiu6w7sFOcn6xSzsN8GSP+1FAJMeeDVeXKYLlom
J4LZvgHFtaLx54LXgiB0zlRUlaFMd2jri+sk9PfOubHJwnyXUQPSA4xl11dxBZ9m
46Yyi5aF4mt0ijN0H9Bd12qHtH6Qf8FSfAdi/YRM99wMi2n/mJEVFgRx1JUOabov
5/QWDEaD8ln7l8AOQ3arECYC8jZZfy+2KiIbaMZkpSf0wTfx+eWMHhcBjBJQo2l4
xyy/g61K1V2n+4aD0L/+zisuf6qDIBPxLlNR5/ffwPHeuyr8oMLrjTUlHWI28Jhf
akAfQRD1vuubQeAEI4zLg57BlA+GnVl2Q2dikhkJQwFwmKSoWxepVY81mazJKlIX
3d5PuacssZrlwtXipo744SQV/+7GxR0Vmo77QR8KcSW+sroMmxuPGcHqWQpgWoia
MGoXJu1PdcL78zcw3En6OYp6zEF2DPoQnl7g2HYtbfIpy4wizktjAL9y47XY/3rZ
kx3bG5lT5W1DCdKexW8Fdcf84PKTjHFJDnwoTLQwuvTHoLG13Y5o9E1Tm7rPUfXR
l8DPqudojWUqm/+fzw3v1fS1RaDzVqFqferbnp3pCG108YQlqPTwEIVj/I54Ob8S
zJHAKxCFRSLyiPDU3Odf6MrZ73NLr/Q8IkI05HYbbmw5c5xFRa3n3iSqvzi6L6Rg
XhmL42Ly8q6lOtkudLLu06QCNZgwTeBYUUx8milA1eqx1fHWq/poc+DMFxnTdqjA
ru7THmzBSU0Ru0l/T+yAcM7ZUZ7XVuMvcl6JakRveHx+yuKHrCyTkn23ghI4zvs6
S969VVzG3PPIjuXViVZN48KqAc6Fhn9IqTwlXCtK0HDxzWABb3Dng/gB2SLx9IgF
gNuCsJhFU73xh1BqCkwP4R60I5m10wHZUHXP5QsRojlZprN890LcaNsFq4MyL1hW
IWV/OQSw0/DngwCZpNe8LuoCFBC6gH0Tz2NIn2WudjU2asXnDUrhr4M0FuAAEW3V
Apr8EIJ9N6f0/hAg9jO9ZdW48RzH9tqgMQBSORLktkNAG55plvSl13NCfxcZcq8C
YnR+f0sT88+4ssUdmTOZBzEIqP6owm0pIUvRDgtjUSkxLHIL3Rfp/oSdKTGb999b
jaO6dN8M/uarnYpRUhBUSfPs31Bbi5JnXR0eEQd6t1jpwpwQ2Yv/o77wYVCNOIZ7
GragbkGUrAl3l0k8FC44kJY39QgJUSd4RgQgPm8iY+f6Rx0sw+xpJrbU/+VfJMrn
RKCwrq0eoOpffqajNyZWBIW6M11uG+LRD5oPWF/Ge+BDXedTTP21uTVOqr990J4x
IGiC5UlnlLVdT0eTe9mi1BMMZNsoGv1uvSRaTuU0A1Fg5+aXtLuaEEcQy0jLBey6
GY+XyRB9yPjPkWvlznVsJDIKaGfv06P281a28ZAjjX7vgMshGZRhbv0GWzvtKsh2
nxV00h1jQfYxpT5oqOF/pJUQO0n0DPSEv0ZuM5eHbFckTR/3fbMyYyWLimnGUTO1
gVlwjjJuZbs4s0kGuGFi81rcQ6jlY40xzQmtUdA1mTsjJhOOpGuX33ypUa+QJ9yO
ZURc9vcQhhrRHESMbsdnsHlQymJddQwXv31PT6W5HMfXuzccghzTldV+O6pOS2lJ
tjgeA0PmNAs45sZBKrBJZKq3wDO4oSW7X2c69ZYqH6hRkzg1v0/YqJfvdlATz/F9
rZGsbHLkij9fN0yT9btXgEKaagSxQdxCoWq716U4a9iJj9/mP4ajsva93aI3YH+w
DvqHJBnpxaXNc8JcKRBdMBb8yZYVfb2qJl4GB1i1pVKu2/wz/4oXWJTUa+xVmL2h
0eB1B0luajxC2MLSQs6J2w9p1ogWnIBBfJCqeVn+EzEXk+tsq4YHt5vgJ/tdd+LR
Ok5ghm6ZV8E57rzukCx820STSTOCnsoMYo9RywpUPyJh28SDWpP7c4IpuBKZS7+6
Mk+dJ1xBJemXqeu/ksruqRFLQQASfmNEoNQsO3Dq2EMsecmQKwU0rl3KdZseBUse
WWdvwvYrzrg4LZBVtZLatLCVJrRO/bmkOMRS/RvIUsnNrDFvysGtbsf5yBoNBw2X
DZcxpq4uXcpteK0kGvMsx+eSz/Rd2xFaz3So6qp8cnCl6gnypRBjhUzRej1CsCt8
zTos6kq/P1n3ZVKHOTbiZqGchhVgSH9/IQsSvWRvo4BnCuTE6VW63m20aH737hCI
yHxVoiyiCmLlHLsgPAp8FxPIWCIpm46EDqShrKavgVkQ/ch7nNHLEVIy0zxC7Iyn
2OY5KhUziFvPCbxJhvEWWRGlm32TN6JLEJGDgoIE1KtnSO7QsQ6jybU5T3mwxQce
8xcOcXbk80JJuVxImXY7oezJUsKa3seJ4eQ2Gl2t0TwFqhgGhlhzEO90hTiBzVxN
+emK7DBIicGCIY0nVKJCLbsAVN7gWGAoZ1N9OndjsZYeNC2MaZfld8y11P+I4CCS
0UYJ+l51cNZbo0HAO7lLIt7NXBovWzyBs1Nzvw3zce/L+1utJZYQC+ahPSEXHpRy
HKBPk8Aq4T/1SKsPKXkGEBMrrPZfnWTaH7e8am0kxOxmftAXGlBjk3i3oAsv7Oc0
ZUox0r/hxSLoA/XyKnKH8LOd1SU0LFniSxE8YC/dDt8wwJmyMlsSMWNgy5wTeDTq
3f+hKwZ0B6Q+bTz3H/u7UJUxSr/bVOkqvHurR8iHHpdZ7SprOdJKCsec1Uls2yzM
boAk3AieXv0xGCqP48yY9Yu443QbJqh0j/Db5smTZhPb2eJ0Zvdwaqt3LF+J6O9D
PdrFqPZdQ3OUtmzbuj1Fk/n6dkwMnCYbgfQz5xjSlV4bA08gZpT0IVDufTrmPslI
qhjTf/pHZV5TaVeV8cvJ7qULaPCmMsTxuUYzz8Be7PH4BIcezi1bNtfDyr7pwE4P
5xe1+JB47UwwStmuP3IyUouOuGelstejikpgR7N2qb0e5xaZYJd7ODgzFM5Un+Gh
8IKrjQhQAsRUbB8uUoFElPWmO1G4LqG9FmRcR4Vl/pcGYf15dsKnBfyMBPgjSkJ8
F/ZszAp4G77KMO5qLxmqiBG6HUvPZ/Sf4rWaylOrQ4U=
`protect END_PROTECTED
