`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
COH//SUCrec4/bH8kvAUCqW7fHJTPEqYY4D9XbDHirlBf5GvNnah9yAl9O8BYHDS
UTvi8A51ZMFGJaogDcvN6tjGNtYbuS0XS2M7VbA04F/YSXNbU8uDKiDZrb8jv/5s
Ou3i8n5mlvkzUiBY2LdToVy2nLcLyA3Smm3vor3EQ1iMHhp0/THFAojfHCORERS8
sAbXuAJFWTW1eG+dvDR3cSpbOr9QOiqYbz4ppT9VF2sIfZI17H4wt7ybR8G3IvuL
LtJlGxNPMJbs6ae2GT8qtkfiBEDK5bZprrbRXVjF1xHwHOGFeHhDEPbKqT11lYbJ
Wn8oj7Yn7l5SlRNjT0yrnyNh82YHdQWaBrmUB5TS+D2OIWDsKB2/+p7eNSBAdhjy
j6HC4jA6LVk4f07Pu6Qrq0TQOfnRncG3k0484KdhhrccunR7jT+nDjHABrOVqtLo
50UBzq8Hn0dvitpvXtk4FdBIr9Zk59kJKq2FrcsXltBWxE7pzAYiRylFpxeJGCIo
ivCKYdmX3ytLFHBnvkoR5nOVE50Exg2jp59uuHiFA0QYGlGGJjT0NEbw5Cdonxb7
6tO8dvVqEPCY4hTWNy/ZNwFV1gdxmXzg4zFp0u+sECVI68xHDsDfDLWjwEG8+gLM
2KJUTwjE0xcIIg/22Jx0LfbnxeVngnAq6eEEZzUpNx+os3RdenHCOrEO0VS2eCba
DXi2bnmUNsZSi24PqNNSmRaNwcvp/msiNfAfGUlZiq6JrOY4epwGM3XEB92+JM+x
PeRpmvG6PpOFG9lnj5QDWvAGlJ0VqAj0KjZrluOkhHbE8Qt2JBFZLXlJF3at14i4
qKsXgMsZBLMwOOZfnUXQ7hA+cwZiyHfeGMlqvMk0KNinyAL4c0L88y9fBDp8rHFy
efuWSo/oM4eN2eZ88lgui1UeNYcKCl8pdETdQLZYlzQYzXy28rPQBpoPLKqCbmHK
AlY/Kv08ZFMfAp6mdqjGBYQQDl4rZhvY2EAZCSZi//GZCNv+n52gaQbkqfARHUol
4Jz6COJw7y79T+Bs+8Z13Ubv0rILi3ZVVDzhG2ZAlpSUcmRgzuq1wVO//4kkSy1X
anToijfI6oyVfQoUydCxMuW4/OCjFkxRL/T+SdppFHKKp8p9OLV2r0Tlwa+OPhn7
HfP8uuF5qIFeiVXPdAyxPwaWwh/PA6lpSmbBP3qYcvZCxAiAR8kVITD4DRaCogTm
JA0thyKeKVI2LVtFCwptjuP6IDhwQ1NvM5fmc9CZWlGlCQkBxGnsEiVqkgtUCAeh
ITHGucSgcz/dmPYaTvAwO+JPvYEYaRQGQ5+FfN5hHFdVHm8nyfwrFVdR9+Lu9qFx
s5Ut/g4NKigcWhWD4sfIydsYph44sUgu+crnKy5xxJY99u0mJ794YW/8zw3Da+Zm
Ep3AAbZ3dOgzGsEWGjl4b69yADSijH+DFWbhWa9bbRYATpV5M7ZlpY4p/VbMwOLZ
rMylR6j0N36ChYnVqRZAOuGu2yeq4WzEviPlG+HL6Hk6qfAnuck7r9OreF3r5dPp
KLoSa9DfA3RDJi5wwfeizWC9PQUho+4ew6Op8l0hj6F3JUQI1+uiCcnSs9iV5+wz
9p3/QAu1MfKcDeU9GBhf/OLR5zhQIm/AhnEVOnuTI5BZxJ3WD6+F3X1e36DLg6o2
dhZ61l/EoKDavtmknhwJH/+OYMhVB2tUG2WG74YYAArAufFOHnPzsvFh3GzCrgyg
d4JQOi6kdV/sm0KegUeSIRUXV2l/Dng7eEIhsFFmw48jUYOvNVhtYA0SlV3frNd1
j3b4BR/r6mOprNfxEf9KRGRndt0VthRkrAmPjrkUPKgBlny2Ett1cv7qPe+0OSVG
HXY2ympCqd6gBGer3AROOJnKqWx3KadObikrnIC88aN1uBLY2JnuXrYLBcSqMph2
8SL6fLv1cJI2fo52FuMUi9152ZoT5sfMJhXCVidJHlRvcGeka4GtLqIyIt1TSFNU
Rkpo1Hv8cbXcn7vN3cMsU0V7wSNZs7gxLBXpZvck4+wpEXzxTV83tTyj3PN8YPOj
Pg4puI9zXEhRoTnc38CZaiXDICDjrj8gsfdLasIPQgvMskcpN4XY9BmCEIgst8NG
WQjGdZKQzK0MPrna3AxQ4bZmA1xUCiM5BbsMRwJxiw/pSY3w67XJX+UgAYDiY3f/
ZrOjNmfPUG2ip8OhRU0B9ewQCw4p3UACJ22xIFkULzfJmRVQIRr2w5A0W/HTUhrI
/VW9RW3Vy/F6IOLng0IywkxE/uCqauT7PRWwwHhdJ5wS3bG8KuK+qW9f/rDpkRUS
/EF4aq60GOA8cY5FvXTmgZmhCF5ThPBD6PtBbvU/ve5tsYRt0//+/veqdUxyxw+w
cXghv0IYQ71miUQtMKsXP79l4ylniCmGTf1KsdwBVMNmAxFrYeiiszLB17pwCjkl
nogP1tf/3Ye9kXUm8Jx5HGHokLUO+iMWyC/hM0s73eZCa9NCL/Myx6F39ifJzxqI
1izdLQyiScVytdPcRBHjtqHd0pU1Clonp/xYfT/R66JS+ZYsFctmMs7a2bpIfqzM
1d1M+kjMRKqXisUAJ/wQKQuiva+fDUCk8ppgrggn+S27hWfrvxrIT86T300cut3m
RhjbY8h/VWByy1aK8MK3YM6sYrCxmmCqAcS73pj1qD0BxL3S/KP0hHRDr9lMWXDj
h7allkUfxHR/ItMy9AR8ih/PZCYx7GGhe2mO/LkDli1Z0NQwlovxFAzQgoUdAyAI
maSEiV/yGweH21coclLmqMTpoY+EIYH6Qtxv7KblhmFUCLpMPYBJ9Rl887FoPyMh
M2mfrYA0t3blmLxYNvBQg/2BIjMK5skPC//gC2uIMK9/dm8VJlft6/abb6H+du5i
5uRSD0fbf8WbId8BHwdEGd++9HJhgxFgRNok1v+UyiEu/hwdh6M8ZjUyZAUuUTxT
P2QmHrV3Q/VQimy43EUSdm+yUw+FvXxn1arvdC50xnEEZC9bIoza13YOclThpC6g
8UQ7KVZUGrcMPixjRjBRuG7HFnw7zDx0jyyAXObqZGyHG9LB37LiPcavbsCWJ9FA
EgY6I3V+LfA9CLsANpprRe6cXsxhdKMrGbmxxy8Lx9l7ZUVnVcP8s9bx0uw7FwUT
qOKXXVCiOzLbZbyeR0auxmc81Dco0P9ro3vcKnflWiKJGfMBoNlqCRrIQ+p4aTHj
3F/iIq5RYXpdZI7CTr4EQKbEIczzsh2ClSyzu8a5iC+0h2tK9tK3xC1sQWGHropP
MkH+8od3Ivi6+cu3x5ZmzT2F/iSg3mUMho02BVL5pVbtdzoRM9ikFUHFnle/I0Ds
S6TxrG1Qx0xGrwbMe29Va5VflndajVwFtukiwcucafPaMuu62xJp5bJuj9BotAUi
WGFpM1OUkzwQCLb9h+vLRhlo7Q8tkoihtDG7GwkCi9V/itNHnmrEvbM2D4wxYn+i
wXRj9ggkkYVT3tDcXC+tUq3LZ+cGltiAQ4tcRkodPWid78uRSv+PeIbQuYGV3LdO
d+jcTgHK0/D8S0kVEAXPNycCfwuzERcN9tp+7fwBsOAT6nRCfihrz7SCNVxcN6Bi
hMe/JBkh9+l9/UqQbk9jILy/a/jgK8SNapwQPMrz7Joq1YhF5MJq8zzn8dRDaAAX
T1YYJ37aoiLIyLqFlRxkCOHKUjoS+K6q8xmqdltL2NwQn+RGSONE9SmN3KlMZIRz
7vQT2fmY6M92kSN2ZlgcMRETAn+gqgXSAzdFtf+DosnO6bK+N99Dhvi7afcEhCxv
o3OucVp83nAB8LpJFAwFIJ+03YHjzFkHDCv8v/iOfdZ4pln/31KBePm7uaLF10m2
A0sJa/78jQHv9s113On41mqwgoNA2p0N5QP9rNhHRNbYwfkBghIKRBJyopB2lOjB
VBdDCGPB8vFGenLnFvclIOV9hUPCU/OrbZw5NnOjbXv+4ukVvtbkYtJ8LOqbYXGN
iiylhB6ln/1RwfQUu4Q/zKWIrYNy3eOd1NlpAt5IVxO+3i0npZ2dINyIMtcX2euY
N7tIe1VKjl4FQ9bJnPLjCxeda4VraYWOiOfh0l12TK75otcekBR4rGFTjshfoC6T
D5tp21zC8asVSDHJffB01azSRmEhw6eLlumDlm6p4ETG0BHVD90tdol7pZJpJB3S
bZQXt1z5UY83emP110KMawiImgK+zqWx0Tak1qCbhp6oWITcNu8bpMKAG20SmVOO
DjChVtwWFq4sbeSP72jvOV+6qdh2e7BLwpZdPSjp1Afm2geFWVOB+igPE2ZEwsQG
tTf4quF45Zsj8qHyoeZd9AR7Nv1aV0s8HwiL/qZRkKm0a8KMcIVYJFFsmpXQo9wG
A1uh+oijSjLa2GqFPu82iZcCRzC02IsT5AQslKmBtwyASRo770Fh0C3rC7vhGzS/
h7NEQpGntlo66VGCcV0413MjI9co1P3Hi7kU2DRzZxrU7ocEJYvzw78Y26R0R7wN
pRXHM/9F9D8pzMC1M/hlwHZNghsWjKrm4m3F5jjuveFB1vmX3IFMwOaXLBSRc2hZ
MhQmycOP2DVyWEsHjj/euMX9TG2S5I6mj0uu6iuWMLYSr9ME3IgEuHIo6/IEhvfb
EZ0DBVUCyLI1TVhpDRjKNaxunfhJwKv0crxfkZLfrBWDxYXv8zARSwz+ouD5urFf
JEeI5xaXLhtywpmoyYRBOJvEpWY4PoJkGk88csVkZLKRkBHSFObiHo0BKgvpEOjI
e0lXVjhQTw5f+7PmilB7Y7B2AyLw04rdF1UVXaUFkwegSDy3tU8MQsVoH6vC5jKr
V8o1coxJ0RWyzSB9YuvpOCyicU405Eq8WmrNHyr/Sf89Ca4b1atGoga4OfVkji/P
kans/TdwIwbsVAqdPTV9b+U5ieeyrW19w+GQBz81Ekzmw+wpYAqbxv5LKl+lck4I
CD/vJH/LNoc/fQPoSSwCU+ByW5a3iB63XqJm2EHMmp3qzCZonZRAv697keaKL/1z
ivnjEI36pq3uCbirGb5xWQhfmzYjfizHt3haz8OQ2NVo/GqFjGKWdvX3P+Wu7wSe
zYxOqBMhck8ghXXszkFF7qRIs7LQfMMeZKp0Gu2tzeEL/tQLoBA18J54ymP2ImO4
ItqQP8JpKaouElv1nI0sa2y/TJLyLLBqUw+dtxdH/qFHpiztCL7p50hK4l/MneL4
DGmpBA7N59Jg0vI7t/CoWFOdJY9cvABYpPADcj8iqIr7U8fQj90b97hGtr4VbJCr
KctqrEJ7qmn5//l/G6S1TiP08eDhpk8d4UGkjwDIxgHP7kCcWTbFPX9HKqnm+1mn
ktLCMyVzJ8sha9OzHToMQRslPACROrQ7TmgbfXvKcSGlzAcFDw4VSgvfU04kJVGb
dOYWxR2ixkPlopOlmyCQLYupyy+NV/yJrGJgXuj8W/GpUepgRUz3n3jD5Kem+UZi
dg2g1lC0Oc7Q8zYBs1Y989miWjNwr3fg4Jb5EVoxNrr6+ywka7AX9yB20UnGIFcY
Pqa4vlDo361ioXXXoWtWoUYBgptfnxYBZX1qzpd9O84ZTkWWvYv4o2Yf2DEv1yKs
DdMjoAVBabJnnGYpvdwuG+XR4MYLGJNCV8BBZqEwhYY0tkv+rhUxIBW2OfOTgiNo
Fl2dYIqAag2y5EeXcNm9mtR5uYN2bOB9BTZx9a68C92mx6fy9L3Pp1xdnGiO4C4j
Wzm1/Nu9vG+eovyVkBxxFq8viKnHzfQ4DsB7Iir0EAvTlgZnteC0iPz1PoHf208Y
V+JhgdKZHjxSR1gI6w70gWmGIWGZBgs5F0wTjo7MtjPbP4GQG3EHz89Y9rlhDpbH
ltRg/NC4DRWlGgnuf3DPby4l6GN5swy6kNlBAyVF90QgoQgv3D/s0gWhvUxmhSnj
owwZa3ZsEmUOGPPOAHzLXHpqu/fimDRhDybLhJVSClCuSW64aInG/8/dN3ofbF1G
myYzv4fN7El6L8W2BDSv+yERuThaaOp/0sFejaLN9UbV1Gc3cracOKCwQ3zZjUjF
RbbzsBrndOYB5lFkD7YxsKDEc6BJVRCDrGBgHiHUuP/o5dqIEBCPGyTiG+WdS+Th
OcCm2TCaSmBKxpIBZzeYYa6Snl9yuf5OsjYPiFQGgDGeiXH4ykzSpaazauKzCRtO
UWOhMMeIlhXn2sbhVHzYxOaDeMNNORq7pJjOIGRAhfQ7fXziTEfQfRNdtS3NkTIx
pGf2BJ5pJCbkxu+FvUuGJKNZVX0Hr6iVDgy2WPSc/HKkBVvtgDduBSlFVrheRL85
xQ+MEEC5SUG61LAOQh9WWIDsvLcixE2KYRf8+eHuQdIfK/m4JxcWmOKWvS5N05vz
1P3+Z1W4gUGiJ+4iP6fdsTmLzgVFGTtzLkOvSEhbdEtm6yhxOjaUPZilIQ7MunGX
OsDBtDK7GSkci4lUEnLRaUOIJgYQqRGRtiKjHyPhzK1qrzyx5I1IACKyzpPDP122
0+ZVzUZfJia8yz+IO4UvRIKzIFIK0aUUxMGNuRKC8ikHGzWxft2zUF9xMmuWmUsa
7hJD3wj0FhLMJFJgxhEcwcfl6hCp0/5kMemTibc7ZnmC8sng5fArOPGBfXyH0uvm
DK/UemsueMj9oQVZnulE5ytOMpCM1EVhJwNBmBkvDjRXG20MbvfXTOpN2pORCTaN
ApPBON9z3JaEfBquRjg48+YGJFvLs+GX4tQikM9xzZcuaoSVZCc5jrh8z5JCy6qo
q/beTEH60XKVBfIaMLQn5D/oMdtBZV20elMJDNIMW0N3CD4FIdio6O83Sdhk5+iT
3G/denQ93A1Oh3xYZD6EWSQZFPuWruQ6+9y7sJf7/N7PECJi2qj/pWtsp9qnCWHL
3kAIAw/BAL4USBsiwdwW1mTix1J36HVXmecT30g03fbq6VntNUVkL7VE3undIdRy
JHUbEeR22wszxNJKk7TjfOT9x2QBNDikyS8zJQRxgAD6pBFsMrcQUTdDQW98OVMx
riqkZMcq5Sl+PAkjdgE4U5luRiR10q1i9rBShFqfQQbwBHOef+C9CDGIgxcG4dgG
/F0TuY1X0okMKnXOqO/pYEORFOw35ewjEWOh6vQIgyMjaOiq5+Srcx/jDg67U6d/
frtxWB4AqA8FLGPVG7Mz62nwwOqIz9ci3BcnvfvVoKp6LJqUDE2zTmBv5pntjU1K
le4BeLUxziPTtYPh+VgROrkO9TIZHB42E7JUGfoUMhjcnsu8Kzw2ZaQ9EnuctYUm
6d3Nmsbyj3nvsiSKyacsyHaEtfwKhK/sroWNE/CxTCYGTYLMXqaNtrif12CCeO1i
Ht6J1tbpOwcvXBr2DhbimMo+O5yYBo0muI509tYPQlj2txSUKycPdntvUGue4Qn+
Enrp0HJGOjn4WhEcQc+KLqaCJXwInGrvNSpdAd4LGmbbqqbIc58sUwRW3I10TToI
hAQrYm5SZX3gEN7fDu8xir7jbxtjoQJNfYCk88MEp0BGniUMqBct7Ja5oESS2HRa
gIUQUKewQLmbW1sCCFsWsvTyTI21eqjzuCIo7DFkjo7WF7lUe4ZXTkKb/qRGUPh5
Wn1prBMPXYfSKseOfZV6g4KIlSy88SIBiDqlFmB+q7aIASJUjAlI++VTBTikU6uc
9hkf9fdHd6vcXKlHvE6Q62Llzx0Nk6mAQbR8FsHrIm7d54AmxXe7IstStS+DZnp3
4//n7Ny9u5pyiqo0ni6jau1XQQo+qHAIB3HmCP/VxH5Aiv86v5cOWYq8Hmybx4eq
exj5XSyoWVFr4PgS/P0MK0xW8m2jYPW1GGo+zbIwUmC3xotxWHSCOaa4H89LW6Xh
7NTHjo7c+2pnydBJFDezh+RrIjc4V0GTlAWm16Icaz/GjEB7ukeqRZogS3Efhy5C
uZvoAKcsD1IoHwiU3VMy/OGz4G5DhJoUyEA74NJeljZmTENfpQZiKsKb+lXPhQkb
H9atLTR6xQf3EXi1+wbpFE7rUrOAER5gxQ00lUXpd6cWFomUJiMJ6o5sVwPkLaow
fQ98JqCePWhHSnMRkRmPTzVOdDUEKbiyW03vIYrXPfzETXhq4IuDtma7kk+K1UYa
oKuSTV3E6EO2h5HUE6j1/sshF1o0B+m63nRWEseCUXxx5BQDU9O7XM2PwNJ0Vt0t
tzqgmiOqcOFPY6pY6M+jG4uRj0AGR7s7AvFUStRIA6L9NK4IN7MF9zOim4J5zUBL
Wp6wakljuyRVFziVnfjs2VEcQueS0GcxMXais8A+cHXNWGu/+qjTkM0MHYzNT0jG
L/qkKlTvvR4SGqhQ5HShZx4Lm3cUkVMdH1HRX0WS8gQEVmwm/MYQhxJ6v8KBWBkQ
HIsyReUXz+o7JD/PqnJ7JWX4Z1nst3HvK5VkoriyOjbnsQoFWeKa2gIQS8Fgft/H
dLsE5gpVkvOVdXF7gSL9J+PbozoTaHGzydt5/IV1k6FI0zUeA7xhInS5viPV85DF
wRPZbDPa4nC+psRf5Ocw8+t+QAzWN7ee8B1LCfsRF98F/g9PaV5NLw3p31o1aIVQ
uJxHyvTtdK3iaTBVnCJJIQmyVEHTKhgStfHNaUCCliU1xIiWTxCDxGcg0NRwVEOB
ubltQ3YrEZPkTBbxQtGg81PhGyfUIZP09UCqDdxaweM3doBeB6ijw8ixGzwEYvUE
qbRYj5sgOokapVyUW4rz8uH45cOdnFJegcgDqIu0SWS75Yy2TYFawfv6Bu8IuLd7
VkdynV5R7IAqFPs6wda/DvpPyOlPc4MVwQ2J8FkC6SYTJC6R15kCeWsbYvbSD3Fh
15A/PBA2o6wBaOdR81AKaAPvuEtWm5oC7hTdD5zX2AWjN05Vxg+3Re4xOzDRoFdR
KOfLqk1vRKaeMNAKGiBRhA7RcCT/nyCzMJlf4uxyqQ44GY11zyUMewdQhWvxIse0
eJVgx98oJKeQsq+F+Uq4EadtU4lJePrEuvONF5YR3HO7py5NqI/tqgJrzcYpSllQ
EYnNQvodJnEaxMrDFWUzUVzk7CnBVrZzduwkbqFrxoR+EfC7ajhHn290oY+umgZa
HPv5lME6UYsUB6pDAeZydP5SsgE+T+o/16a/H8TXIxLN+TCh/GNLpjg2KjxVF5Nq
h5v8WLByyBLqsec0k45X+QIofT3k/PC1xH5CmTDlzaUw+Cjq3WzcsccSbgtzuagR
IQSFWn7/BqdIUJFGdonxTmwb6jnKcHDsumgyuECfg002svdLNjioMVvx1sXbtMq5
46HKnMqD28dPri+oZvzvC5Kt1cOgdWoQl0BKRk2utNRUtNIz57SbZjKF8sfFOJ+9
7bSSynHvdXM1d6YHQpPI91z4TNs4oWKAQ7ul609BQfaw8bTGXPJF0+rXXpGaPmzQ
KHMFxavPVzLIYRtm9HMo26LN9Q+sl4FPKHa5KHEhtzaziwagwjFy7EFaHHQMgs+I
SoPrAwY35u9C0y27dhith+QbHKPQWi5fXmBPugMtmlNvH5qkDZpPdnWbdGZV2jGQ
0fV8T9D4yijAKETVrtNWemDxztFhP3ssVhgkVkgVVejGewzYJ6MZlcZuB0pLkaGI
xQlikZ/qmJPahojow7xJRO/ad6GgzaxxPHIglwxptNL8CTJjiKmLm4vXPsDLHb4f
Bv9zKyjxuDcigViYGEynw2h7l6D0oCRx8/jAu3mxoO9fl0S2ZvLYqYSh36oGrcpL
OvaMJhdRI88HNu6OLsGxT1nwOKS2sO5yh8xFOHvKYjOYNulXQ4/IU2m7oXoQwC/S
CtC3UvxpgEDYEsbDy+3n5AAjvRgKESxUpF1z02yVKgxDPU1ZBjlX4j9qyVii206z
yrusUrHZD7DNCzMlcKNnw/RKmMTMgbRdjda2bJA+qu+6VlU06hgoPW9rneqmzA9c
a5vOM8zBc1C3nJ7C9/5Oqb7c1xD9jJ1ehIf95c7B+nknPAJAIHpgRu4tujGfnMfZ
LZ2Ezqw6aCdX99CdDuBe3jn+rXOQfEQf4g9snP6pdAkfPIiWNzXDdfqX5VsHvjPm
CIPivWYdSz7M01tXPQRevmAIvKuKc+qkxLLCTb4h4/r2PNOsg4clKbDfwHg6GEvW
pz/9krN1Urc43VnjF6Gx7Mc9R//13siCFE7Iagvra5GJSzoZ+PBwPrjSmgYyTyiC
vjvBgXz/gwJYPD+P3ryJrxtpwqFpP9JoRu4LoeA1zB21hxj2G52IWsaDqqv73KF0
iCDkwqcd93qiN3HkbdxBU31dXsm65pbi0J7+JzL1xFjsnd4fuFYURy53v2vDuKl2
m07+mmCFdIp1NwMhvZMK8mn+f1QDRwtbQ998aDJtkpIjtD+XPmDcbTy7QRe8wFCl
Yygu66+h56M88Z6RcrNoALXS3+sOH+RtxfbkIBUtwrWnknJnIEMoITlINKvUFISP
/oS7v8Dh1q2QrGbvpWzVxEFWaOudjzX5SQXEh4bgrG898xKdD+cS1LtpY3ZEvRqG
BLLjU8lwZCmeTSf8XoFpx2n8d1Wkt6WKIsoulV/P1pkC8W4XNQLOASmSUCoRutm7
sxfHO/K/s8jVxA9s2dSZvkEHdRwub1RVCzmFxnxhWGW6GoGxP8ttZgV8x8jXAbi5
ar8z0WqBtRMFG3jJCzKFxEUwzUMrqaOkINgOfmuC1SStOtunbyUWoCWANu2M+YZK
2DzmC85Xaoypoxcs9z2Irestjyc6hGQTsCPdApYvt5PhJE90CGFq9pC9y3DotPOv
vHugzQNcTXVI68AEr5waDQ5p0KohiVq3g+X2XCCFrliocXK49A0LzCO5nco+I0XD
t/Jw5Mc6PZJbvVZaTk5Dn4HqIkIyCKNL3kRZfkrMDYEXvza40pr4tbbhre6Cl1Bs
tOjh+UTYCuHqbHZvt5XfdaDe3pa3UGyzzndqVtlCMw5fPiBoHX8ZSkUyW5i/Omr2
3KwyIOHkl7Tp0nALO/+YrRv5RmNAfYTB8GDvjzqD6hvoDie4Vwp/gOlsgczUYc1O
rFUJR6vPmSI29rx8xANyWv9oZpL7/NMo7sfIYEAhr3awxTTpOiKnNiQrsiAWbsBP
+e7e57qPKbzyBKT5XRzd0n/iLZHMB0we9M7jr5jDV9XbdLPOVXbCXdo9wQGI176Q
N7P7wDDfv0yQa7TAKF/wj2n82D+Wr1hHTrQq0bFXi68pLTkYVCpVRJ2cFWH2b6Hx
3O5LLcWvIfLwTYxeQPhBPsjYb5NKjlJCoTbDmYDFl1wyVKePzM1gKp0uczqnSdOD
D9xd2iyDwJ5e12Rjpv4JObyyMVhmlwW8bf2W1AHJm3AIsz6s94PWIgDVTGRC+Hzu
3uM1SpLVxbnKG2nk5bRDb/jVVtohS7OSheJZ6AsdgwT41QfUbXUgkf9RPEa5wXQ5
pDjkUzG0YAzmbz6Dtb0WfwWQuVOBhgPS3TQqLlv+JpzPi7Yz6cWw7LsxdM0qWHxh
u64VJoIH1vWHkkxY9KpZDW/yZlC8Nck8/xL/XnpZqCG3RnWpHYFbXBBHFd4JEuGI
K5hJqddWBK0z58qVaX+wzUwlviqaUUev3L7IwTTSRGTRbs8gJAk1Swy7D1sqY2Uy
oFYSDvm//gYxEfzunUofgTGgz36wiwifVTtsPqTx+GGUpbv2ow+8/eeR9XYKiL4a
fvvkYTipdlX0KNEpE5GjcZPLaUyXknJTBTRQzMaEdCwT2k465WLUDaDWJxWnAhGw
noj3wO2DqwpLMhi6HbQOHFM4OH1tcVS7QRIAvcYcI0F+CSYpwruQZ9DULiPOoTG5
EB7akzke2ODnj16PKjCnBrRWq9nO1bqFofObcKZjiTnTVO1SLP9K4FzXGHz5Mx8H
FO6M1FGu/cLw7mwp8DdJMiKHN1RJ2tCzQoed0aX1rIUgo9PqfqgvUc+XVSqAYlXL
PAU+Ysu8+GfjsxWSb6WOUFfNS4HTEwDyhOxqKPJaOfce5WvLYCS06LyOg08p7bNb
Up0+TNZpJt15VPr71yo7GX9do61TvIxkvZ1CQ11Ivpr1Knhw1M3MP1EMgp1WiV4Z
w+JeeXt7h0VfP6XlmQ3jobmdOp7Bl3AvKF3OJlI/9QupLU14bVb+2BOYtpdXfyAT
EX2f6c4j5tjrouQUVfmcIIUr9QEB/nNyLT/jaDiiv0DJDMCI17adzA+cNq3ppC0s
pmdfCHLA5/zd9vLFCY5WbP191lgLdNYPXXAmfTWrD//3jC5DkBCxGBpd8kXzu4Ky
+QkTlv8HU4k9l0uHmH6fknzPHJr8TCG2LS6OFpeWe9QwNlPWaLgloRcQmAkx9pr+
7uMqJhfURPKY1e2CNlJnSU/amhwFAmIB86iDf8tXirZVpfHU+4YOoTrB783Df9a6
MtruLV++Bb9mgvxsoLIuZ2ak5r61n/Uqw5ncvbtBOcz8KBZdk7rYh17EAk1yvKhg
uBWeTUSb9XgdH3b0lOdcmvu+A1paClaxBW90KO6QVxufyBjcFjAmj3CQ61NyZvne
MhrAPOIJ/qbrnVpNvv/zbzAkIUHOqIYoiudtdDUSaapj3vQCjSkUh//cP0eUU+RJ
Idz8nzXNe1nqucr+UTYWGMUuZ+iy9dlO+rv3EDYrfzx2v0qRPTphM/gQyWvupDOf
9mpnW9B59DfEUc6EGXTcPVfD/6IBvpy6jOHnSqlSGBMDb3LYufodIvJWIZvHMoQK
BqAQ/gDl528Bk9JKsnpmE1gBm06z6ZQvqSDs2YWeSA52qJ3if0U1v6ifREzztSjz
fEwuLrlWv3H7TobqlyfUjUDQQpU4IEWgPnFJLo11/iXUiYwhz2c6mZ3vGGnaYGCU
wchG5pFrQbQJZibzs0Qs3zmubKGoKO6y0dHj99Rr7llqSf/gKD6/akKHUsN0SQyW
3LrFTr7WFXP7pYgqQMfDSQUYlM8ay3yaQqtmxaaQ2IQHtYgHrvgtTLUG6/jw3xV0
qcH2BYIUBwUeBlMgaF+buK6LnnsOeEsf4SzB54NnK5is7/+V+RdGRKde6WhFHmgJ
WfqnJFccp0Vx7oBKv01+TN198uTxdMjHTuKUb0bNAWhpIcTe7Ht9W03XLxCf/ZDI
39PWSlN6FAZMLbii7hqJfqUBBkfdOHgiat9j0GHEJ2OII3nDfUZEvJiUSWB0xQNY
FwMeDjHeEciyHfYPe4enCZB/wvlsP5O44ZkL+ry9ncLD7p+BfyGXUIuJCWsmJhEz
brqFTfDyjM5ZQgQlkkbZjS1brB8wBgK7jPA5GH31WaFMO/LMNZVJQpbOJ3VNpK/1
UVIe1Ky/rGZEwHbs5l2gpwG8g7cXV7iYwWm8i9Cvd3DjsHh0fVcECwr+FrE1LmnZ
i97Ra0/ICbwNq6JybN8r0iGxg4jQAYKggPOo1j3mvxJamXkDt/yunnEqsqvvPIIO
FXu/5/OrlJYj8BAI/fq9tGtD5b3r+vWvwHoDfW7YNSATsSDoAg228s7pCLO8CeAD
hdtMIxmMjEIMFZCO6LhLRTQwiWyj4lhwWQpFgYeQUIEinPShVRwMMBaDWbdCVfFp
QHbVQz5MbyybxYKBmKIot39yiuk9laxwVYzpnE/q+bq67PP6cDKbu82Oq12FgL4m
UlPH9OGrgsMbx3p0cmokgimeezy+ClitXJO8ZLwC5glb1AFoizOdantCn8CRTiSh
5QzzJua5Lkf7iUA+T78LR5bXb0huz4zGLBs3UANJhQEqpMn6Z6X4KTxV/jZoy7dA
zWw21OSFO3g/B6xkMwFb1eBfjC950kyhzCjJ+uL3HbNdQwrbHoJ8fEgxZLBG2/Xb
Mo4/+IY9dMnaX4tj5NE0oPEmYZe9Q9AsE1RO73ymBdvBuzB2mZq8twQNgZqOvsii
LCaCB9tgcU44FkaLHsFPby+HFLwNkVenBfmXJTWIKEheF/qLd+mLEzIeSZLUWp9n
En31klCM7Tld+rialQNY18z9KuCD5CgJ6XZVui205+ysyJ+MBAybFvTj9fk6WNUE
epus5jPKJLzjdqlVbqYICTZXdsoKhH2EdSqu6Bwp9XsSw1h8eguYhv/bP8bgMEP5
ckzmiZrwrr9JddZmUN2mhiKkhrY0QRjhLXCpBXbppczvMIu9oFWQZr21gsOLBe79
kegbCFsIOnegefINs6nx3Qsun4K2rh1uhns5TWh9EHBB3RDcfwppEpWGVOl6p2XJ
Vs18KFI9oaHiyZC0AiNuHL/DnuXYI7BnW1dxPpsQSZcrNUvznZG8negZBjsL4v3A
M6w7Sa2YRkqod2iv5rAgjonMPEAqaGvn7j8NF51q4d04WsOZakaLPmjVBqTBdZ2t
u5peIbsjmc6EhLy/1dryurAT3gM/3CTUOzh/sunsoc+IxZdeFUDnsA/fWiio4wEs
q1eoZeiO8xiJoq0Fs2dsJ50/PrP7iEgLpJJxKsHPMHlDTvKN1CFs2PBid2VZ6bWS
K/tS0sZOB637S8BSCqFQQlvRdO7LZrzs+4WdCtOinwB6ZxLHbZ+buv8vh8/Qc7to
WNILU3jOQW1Bb4SRMkj06whgFWxTEINamX4TGt4z6IgR1l7IjoU7bgs+U/veOj3c
KWAKkMfXx8WcJ6S9bQmAE2F5Ke6MZ1PH1soAjZhvq4H4tEOceWl+q+gIeO1u2R9/
mVDumLs7X7JGTfSv8nboSPTAsXR5mxfiSBck3lhOIeEi5mT6rIXcSxj2crzvj9FE
80aiposOMNDiCRMvL3FYFTPGFaExF4latA1qBrxBYNCqyHIlB4VWavVRZrhA7ylR
00hr8NPbSuXaui/aBWJVzraSyngo+UudsSNOEHq2W/0jS5BBwwpHf4SwiYWOotK0
NG94EzVFl/a/aVT4zhO37JRZ2HjjYotGzLZIDO8eMmnRqv4JjUenIzG8eWyYWTze
kzNCzW/QiuldmV6RmNJSPNfsV0AfMshOjFkxdkdNlE+B4ZhQF4npPIpVLIjwBh7u
rj27uCDITLP9vsqb8gwFje1msqBneGOaGeIwPOiDWdpt6O3I6o5rL3CQyaERouvL
uBWbL1YAiMATcvKmfk3DY80q4r05QbleJKbtMsZ8pjd/iIsUwrxFBpUH+17S4Ghe
PjPybxIwgjc/5V5etTjnclTuKAUEDl3mhe8H+Y/9n6UdG6Gt4KghgueMGkfhC3PB
a+9wvhsvKwCnq5xuDXmxKFY+tRjoBFYs46Yma4xjxyIWIyHkZo47WnxiCgijscQz
Bd+q2S/rfH2+13K3AZiPvQlXDL+GRmSgLNZk6bUmvvogPdgJTixSRDhgn8JpkjMd
tZowwX7jJJhWoevrB9cFNSbdVQURkaHTNvKTZB0mOpFeVcYWcwtuFusq6/z3Yfg2
ypBKicfmEg2Bf/g2GQqBjPAqMCEHw5b2CFwdoO2vyxq8syj5kp0f/a0muGddimBV
q8tk2aMqBeyhpmOFbiAdocQkfbrtn420UYlQZ0A3ErlIWfG01DsUdeozK92aNfRN
p0WBi9UOzIEXJ9O4s8i55qWJxTEeOhFlgP68Z1yHfp6U1h/7Wy9bCOCkY6UFWSt7
F3flQwB00REOjrKY8+tiejgpn0f9Vo7vfm3Up+ak3wRcn8Ffg+DXvFybFzxDxfe3
F5cZ2cxphrfdfRhIoxDQC8VN+57oEeKRse1lu9TxjpX5nVYKDS1O2rMP67vDLW2Q
Azvzaz+1rp6y/vCbhrHZ1QwOjYeeTcuhtKksGw4RRcDJusACuMYNw0aAY5DQhdNs
dHCFEDwE4SpAWBj0uhuy82zf6TFq3QdxXjz9MA5/ccZetwX374ZY+PNYdv4K0AVG
Yj/iZAy0cfUzhhcRfhdh7LyqfhLPjhHl/elg839i4qv8i8J61rZM++LhPOzGOWuF
vK20xUZQKE+tUsLDmPz6+StgHCi7OCwl+npR39QyABnRRnhHCfWmzPuOzTxCvszT
jMG6tSJrKg7+g6nLHlczO8YeZPc6qsZhZvYuN2m7P5jO6wMBxKACitge2zC8b0J2
q0HWeUE4KrTdCqwuJHG8fqyn6IxRsfMEn1iPeXqujPeTGONjq8GE1WHuOZHs+bU/
jwMaLs1Yho4GEnKSivuopMRQm/KCz0uZBt/jQrDVjoX7jAq3pU5pFRgRmrPLI6ws
jkzOrFE9v0eTXfXk4daDOQKP072CTffy1NjOKjgGcHw7tsYvDSbHFT4iDnjeZDN+
YedwExhriA4thm4WX5HXfwWS7nRqK25MCBNTDYShSorwMbwz1oWmeSlr0yS1MB3g
0hB0x4g8c8O7KCyRIwzAnQnJlOdlym4FDEeoeKxNBv90YvzgZYV80RxfKXnau0dO
JQR9/iSeyCq5x+JHJtA19oWeiG58TsOYYvLHSAbUqV3i5hGDEde2NRCxDaYEYPm9
ZFBgA6x2TinRnZdezSy6ChJjkVD/jbU17xQ1qXcEmtV7F/sDuE2Xe+9Wz3GK68p6
/UBKhKcIA9BuJKwi4PI9Kaua4SyVuKHEVSQO+GngMkWdxS3EufaUMF53etKT+qDk
qfZzGi+ka9B7tdpiMjG8EbkZ5PgadSs+MlKk98Go5/01XLJT/bS56ZlBH/RjPqLl
TdCbgi6UAp4G6LjCzxL2lJxssXQg1WpSW+enAe8eKKJzaf3g8IlwyJli/HBvZBbf
i9ZwRiou9skjI0njjeCe3tVGFVGGtre3sh7rXv2+PG4tP/JFDJjcO67lhnhbIhYd
4iVX3H4W2PzayINZs3RE/OXcGoKzI92aBIuwoP52xsQ+2Xf1IoUGPwGrKqLA9+tM
4dWqK24XiwmLKsCsrrQxRG/8fhJq6ZT0qg3AqmnB7BJ6E+oG3nwsV0zz17DwGwAw
h4DCIymNj0NIK0Oiq5zhPFCUZ0ZbfnhIu6WDFyVl9cxsO8iusWb1JgQ0Vjtv5BFD
pVEvNIeYefrukwvB5ZQ45Nnc2faVpdXoUtyWlQewxFEemUxZP+FUkhlktuCjexw6
QtYfV/bTHOFkoCIAur0JsiQ9YQRrXfJStIEGsyeT+QUQiJ106JWK4zLMD0Z1B0XB
Js/ExjyecLFDiSapyD/ouWZAAcN6I4DcuLoquSzM0OvFqXoZVgNg33tR7FTcKWTF
agRveHw6GNnLmPr+Vx5SEDox4IaPZ3rIJUDtBB4g9lAdY3FsVDFOAAOl9F0B9QvD
kyZtdw14e5SNp6gfYvmTTiUkn8DYxMZ3pAarv7b6ebE/ThCMEtcMnxI0WIwHHRAo
yOthL19LKc5ATRmVafcSgx3uy9XyvGDNx1S5AxLADopdcgj4XES+ZB0+zQgXG8wB
Vp6UYWtla5ZMkuJ19dd8g8F7KEQsqkSprCLs24MDp7RLvOL6UAJDsx1m0HzgVVDk
x9SPD7kAQi28XP333RD+kFmu1c6Kvf/oaodiRjG4Oi92WuUYyG5bPKkFEOhSQL1O
Z4Vsb0m7od7tLllPYwU+KZ3nKej1zXIJYQDHgWvsTqFlcBnT8BE7ZPZdNkTEB0Ik
avDpmbT5VC4Cuuvw/hOvKcb0S2jjfU1h+BfwgjbzY981IqJRwSeQ/3oh8BXUCb5j
s54LX1/u/+stYMf/bwqz/+KeTNZSeSDK/pKF7seSREF6XVj61K0VT1PsPG00qcU0
R1AHYsm08csTfA5O45SaesncbtRZ3yTQc4putN2rI0l6C7+TwU7L+jeuDeF40fZL
2xcYLCDqeXhwH+Lr1nJ+jAIH5CJA3csc10ki5t9oawsSsFv7+iIBWDPyjFZaNQqN
+y3/C4eaGKuaIDSso4k30ad5YkmJ0KKQrRmEqvyRNBSDYNkacjMa2oTJ1UWrh3G+
CSvB6M0PZ9RntruVEoLyXIGmC8fbqiJJ80OfxjU8E4FzkEpqU/UKUeYEJe0l1Awa
3ps4834HlqaJOAHTGkA3pMTqdmCi2V+bZ+cSpYoXOXHCiez+Is72iQ2h73Pcqf6K
T+L0sHcm5clFRY9Ce3SfOFOPyOPDkWAlrzhBzQ2yt01ymYh1SziP9xTk1DYp2GpL
s5oL4n7tlfig6/btUT8zov/tIndj0d2/0sT+X03+m/JRw0YPlOQs+/4DJLmtaZf4
nAS2Mz0xEWkuiAOZNVGbYpQf6uguP+qF0cHnErqmQoQQe3X/kWQwmLZgrSnKaHf1
W3AREUvzMw1vw/PyUADmlNrHs8D08c8ewT40VI53qndOX/RXgdd3HXeO8drr1cms
B3l0uJHH5Vc6AkB2SvpHkxHrYedeJ0h8PyUCWwow83YBkw4MiQDPestPlq4UUN26
1O9Qze4sXTT/u7tVg4/LkiBYua0Nx/+LCb64mDCq9zskAZgre4Um7Gd6JB1L8OW0
fBQfJbIRNyFRiUkYkDClZgXNdNoNY/GfuULdvEPomlerZrzZujBlVszeZFby3p0e
RYPgzlMXtpZ35sGuLcDXyVHPAcx+K0NgUZN1Z/PuIrHfimDI1oUcklm6bPBNRZMz
JPkBr0z1wLyYn59Vclhxq4uKryV6PaBi04sIUrdnDE46nCDRv+UWbu75OzWwJwAU
w7kgs9ca0Ru/OqbPrfLqpWFx6+sLNJMPzxUTSIJOhDVWAHS3XWP79upJjk0OA0QV
uIJBlopp/WNaKB6F0DFlmMPyA+7/81ennbClw9relvVSBIczJVZweFhJCW9tNY9D
InfZejf3RmtUEEuOf6Rr9GxPRZUFye6LmV3xUDtDD3SAhfWo0OGO3XndRqfkwM6w
Hur5q5+CUvVJLRMwSM8CaINK3nZZuFalL4q4d+D5sbncaupzDHUxBeBhYZpwcwz2
e8Ltvm4s5j3IWiMIqkVEGHKBDP4nn8lFoXANcGACSfTCGFFd6EavUoaWq/7XrGFx
0VlZhIWMEQ4vkZHey5w2kKvIcgK34mvvlAY6F9WfdJwuvps1AgDAoeeszHimAbVQ
B+nZAl24rOxdlraCXFk505ZTyB0q+eScc77SNyiewYzmcFT75I18qvU7h2+x/JRa
d0/b1QgkogbJiAmcyJaECTVKybAWTBe+mrlQI7rz+TTgYjkqqcufgU8+L6+MLvli
8qJL/nUJAmFFgOz8KegGEMWpCg9q6UzTbuLmlwzDfRhzKH1tZbC03Fh+JxaB6Vt5
Lrtht7SB7Py784HjcbBwZooMU831eIdPIMeqLJpfgHnNYoc6tjGXfi9GUI7xCY/e
/Zl5cAe8zbDDobRoGNwmoE4DgYvwfEA6WZhvb6BLk7eJSqGAZjXABj4bUAOlXBI/
iFYSR0vG7VjO4gh6ty52Cm9vlNt4KVaDy7HkiY9ZTLo9YGkL0ZIjvjfND8nlYGJU
bHxWDff/cCyiTXL9W4hfQ4VvoPAHi1buPr3ZoLvnArP4/zVHMSrAEp0wW9fkX6bb
I+3PmnCDRAImRF6heIiGrkKSdrXj5punspVKVVjnRjrOpE87uj1+PfS2qA173j/P
7o/cLibVhy1rxJoU/Tk2aSPzRoohkJ2HnqwY+EYe7GYTaic5GqWgP2WhIFPxt0S1
ko7pfR7uc7w3ju+FGzhCJgkcd11QDy4le3tZmtMrT6D9B4ttYZ/oojbKX7OenITm
kO4PoPOi+2DNvVLoJNDbXJzl270qLY6ITCTolgYs70MQGOiK6J1IyQSEFFZEb3kH
U6f764sZGYCGrJN6nDAqIqGXTVlbEqU99discT9NIBnuvn7EIa7WzlXh+MjP9dp2
WM2S8csm1ixj7TttIhct4IhHpSLKv6aQYVSJdPMJyoYYhgxzCvrEuKGx1wJi6rmI
vKXEWSSCID/WboVeIH6NFj82i15flY7AXMemfEJ08FJL0JEG6d9FqU8dVL+kQoMP
N76t3eRrRPBpneWomqDXsaBzT7105t1vo9623z3g0oV+gIVoBhFrrEvqTnUXBgFb
dByYC/u0qg1L/FJOjexUKZw1ZpT1Mub/Letb63U21wdo2yYF7vSHouX7lDOT2M9A
v7gL16sS6nCdDBbc4I/+ZGdE+Vl/lZOJlTlsQBP4PSdlpUC2yNGFFHHoOnc3v1XL
8DmgeGjiTwIuybIjNz3ohla7AwUZJSSQOgDkIM0NOxQ5YYaCkQUWdJXrE20Lh8j9
zQk5VbT7ysMl9BEvoCUXGzonjots7ee6YrVZGph8sf0QGoI5yEel+ufWmiepVmVa
QGq0JEemm3i7u0v9Y5G55UzUuTnNEPoCYYgk6BeZJqIwYdOeJnhrPJR5UJP6ujuI
p36y+FtluklfBUWMx/l3Q368GKeMiTK0AvV69TiF1CumeiAQewyEyHm8TaMSA92f
EqwO65c5H8tNX80mQHAtv2VqncVQ9VRo/9lE5H+d2z/CFzIVGgGFhQ6z9Igs0HEd
VNCL9hlSQXnpFwzq0rznsjtAj3EKznP7JtOSQwZdX60fSGPJGWt2KCRPBtvsDaGz
+V46Lmf8Wt+GmmBgrhAElpmIdzKaD8gMVaijg9z1s9lfdgQT2YTSBnoBt+z1bGRk
wTX52vhYZRcifyfUAY08yZgwGTdisU4crzKfqY3XgZKan93OmJZ2DumN7zYFDbbr
LO4N//8Jx3JyncjK6xsIuDalD60dVEcPBTC8wrZrGglDgTtqK1V9zZ8drR+E/N0X
SUzZDPze+nX429uDBVND9BKWrY5R1nVIwxplSmonXiZ4Ez3YjQEunq79POGfoqDz
cRQOogd2TG/Y4iMRedsO+/JItNYg9QmiKVw1qfvaHT0tew/90c6TX/9Uy4+HH1er
PQaTvE0gOW07/Xv+87fUOgVkEqt17MVuRXCNYC/kpI8MvtP1BoYWvShKgnV1U7jA
CkFKMwvXyTMQAztW7rafYg9MFzq1NRxxt91zuexVWD3ADN6jJS2r0SeMU7HZbOk9
zhzYPA6ygrzilyk+cpVb1QpN7p1yDiA5YtRjChhOticpKUFjB22A4JIM+P768HlI
pT2JBKHlik9EGiio8GfsppVCUWOinOUgkUYob95r+n5Cge7/PsetPyyxVvWCIYGx
dCJ/DsNyItX31CB5ySBjl/ZwRZnfFqClToLxN61uz0b6arJKTZHbseUh5xohWmHi
c0dMCNmM3oKZXhBQw8kgNBI+oPTWZW29EUeVLn//Fj1K5uuIYzx3/UfnNqpQJu6c
a4pj+ZTJl4C/vERhwMwkbyirhK8EfIpx70ctmVTuhSCeWV7T/Nov6pSxrDfcLhNF
raIgL0EYo4QM4l/SW3FlytEKlKPmU1WeAZabpak0ctMnHYTEh8iZfXMx9ZHoVvW9
sgXKNCtog7bijX5mC6jhvm7243bCVUhG4Rh9iMCoxgs=
`protect END_PROTECTED
