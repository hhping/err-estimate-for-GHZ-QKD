`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6n+PqmjqbaQXBDfzrB6cZn/dU6qoOcOisflOZepWQffR9j1wTMEcN4ucW8m5/WrO
qdc4JbHwHX1QspZhHN6GA9+7DwfNB+cZgUnJyc9MqGQyup2UoakYB5amuQQzbgJ9
/hihJ/zpyPZjywp9YK5a0cwl+knvNuEQE2Z4UGvFo4jacnI0wnm0SahoS4DGmYH6
VP7ee5HscyP8RhX7xygeX7P63jFuKo/+5VqRF9lBGdyVQgTWR11qpfZJVycy5NSh
YOymk0UFxKsz1HEFHhjxFEe0WIW0LckeqFff7T531RyHV+qZXzJWqZicpMYZ/Dlb
FxCr/v/J1YsBYsHhcc0OJSKaqW27uOGdkx6pCjZZBRRNw8doaTsN1juk8QOGZ4xh
TGgrbQlJVqkUv1kRYCHDIryxbEbubIpN40iUc9n/e8eRW2erzxMy+8LFtTEsXEAV
hRPNo555+0bZDZT/9Dv8geSFoaTxaV3qCVp0NL/GGD0MbC8R0MbahA+aQYh12wZR
ploXmgZ5ht+vLWOyUAAgl9Xv1BRu1fqzOLrbzGug4peucpVAl7oyrXUq17c16CB3
IJEK76N4ACq8qqkxogoPTqxdSITPkwJUxinZolI6stqDeBN+Xze1c0/CEhuFi0Gl
cR7g3XCEVcPDYwTI9BVYJK7Ux/3cYU0oyxwvhkrof+vlMUH9E79sbpEjfXwbheSI
NEtKFyrqZJdNSmCMmJ7N5MVg8SBOz2B522z1Qs4UoN9KfXYWTnCNCgixKN1nhMTC
4N2a8Boi57hYvyadyXnvA60YFPHOVJD0cYoQt3mOb5I9K+a29Xyn6U0ZR0l+aww4
CgUE9foMA11yK4AhoNQgzrxe5RWFBpdTgpPnqfvjzk9AWmfWszrosJ9KdXOe0SZr
Ni5cenDZOt5XroBSAbXJiWk72R6uxJ3Y4ZPsAlBaGERyxt+bTGa1w5U5uV43plek
P4QHaP56auf4qDVYPsIthvCtU1O3UOhs2cLsvKFO0PlC7RSSrqDNM7tXqNWdxk69
N6XKwzq0DpiljNMdbTNUHug01xh7L2YL7np74sr3fPCDSZNB3dCDpG4JBJFyx71c
v4cihtCgTEvythgJzVTwYq7k4A5a4DA6HeekeIQc8Cvq0OZH1Mr2cGk5uCQJLeNX
KJRGHXzyw20ZqNuS3SRczZ4aNvXtTmkG5vXBIKVI3bSpsuv0qPJc9EnpJ0p+GtjI
pPeLD8AlJu6PGvrv2UUvJFpN1i9jbnymZwZXeT/BP68kYq+UVZy7zqahYt+MaJ+K
cYp0kGNqAalu+8l9KDZ1/gPZvivIXx1tnaKH4X5KQxJdVawqjRVc9daZip7U309L
TZqBt/zz89rtps4EWge/puh1Ea0vg1VKzjC1CMIwR1TFnQmRFH2W4n2PFcI6DAEh
ozahAe1mYJqKfns9axXEpjIVAUGRJd1Kklln9W4mburlMNbuld7+ECgkpzoJMPyI
X8wsfgk9ToxlTmgQk54H9yxzDF5zW7egD+/ZuO004o+n1c3IGANPMvFgiB7vJEJ5
5hDGmP0e/3eSM/F74uTV68cUoA981JqTp+ka1BQZVRsg2zAhAMrXVpNvoxPdWD3m
15RoP5gIjoPvb9Sx5acYdNC48U3cYpIx2ssriYyR2Pxvg9ZjfY53cHfcDiwl3NNY
gx6nKOT67NUyyr8tSs8fnIVq8ah6WtpUE7w4bKAid41J1oweHST7kua15NuRbAoh
J3WSsTaSpKDeb/mpekWWY30ZRMdqmIg8XXB8ePH4/ge5oi8zWdGNNWYAdhBBQfoC
VphCaD1XKe6ACcr2qxWFb4aDbMsukuE06Ge/AfpYY9UjTvysdY4Zvs7IEp0CJ70B
SxS9UMPTqW6lre2B3vNxyRL8/NM6yEkthopjecYoLsYn/kABxwfgePBY7mEox5CM
iMxRuh5w8WOcj/mfZh9J2A==
`protect END_PROTECTED
