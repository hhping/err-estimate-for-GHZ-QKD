`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M4Z3ivT3OExef8Za/bIcmFP6nkQDXwyFgxYJrwkMQiJE7apAUyjrGsuDMCBoDwqN
H5Z5I+RFBDXugcx/rPHbY8/CY0JaVmMsLnvtNW+iQILeIK7REBVf+6byAmvUMdMn
hetmDP/rg/wEw446Vip5NgyzbmfpPfpHDswrg8mQHwfZz99+mWJK02qiNwgxE4kd
tFLNByimpMWekYdZZ7SBWPYM2lDYKtW1pshWjstAilI1+oTY3CyHwM6mcLgA5ubc
2Rd90t2E78lQSlzp3eJ0JPeqhoS5g5JwrqM3ZJl3gR6aytqywQOnI7vyxB3yVU1M
MCO3itsvqntyDhxsOUuvJ2EKwo8+GTUYNCFb9DjhwetcwguYrZjjCdRmFSDwuxIc
4sSYqhCswNvm/PX1yf1CDSmjgfHoQ+LbNG/a/tMWym3Ti1XDE1aIg8zDdetk9enB
yfkfxUDaYiURxpuKm492PUJyNuhLyzY+ET8FhTk+GDhH2KqQy5cLZ8LbIca7nyPZ
KvZGt4wP5ieGVQCG2Ydzk8ITgSnRTWYIBXEpmUyg8Z+j61j8tqHdCmmB8MmZdpkp
DAzuvVsvJLhWOY/J7jqnmShwKZdUYGbDIrD8OfwdUYVyPJbWQNOMjsC46AzzagM4
3CjohNSy0WWYYmprMZGyMaeTRAocwkUXpMqwkTnPVOoQD41uEOr4gw55Dt6YG80e
EQ5zGc1LM1VCjwb+JGhkdOEBVWP8dokosJkKwD30L8cAu4RYt1qVGlk2eojDZ2+8
kgob5ZSn/K26RwROEbN720CAFT9BvWrCb5CygpDlD5BnI4I4Uv2aGQ11Mi/8zsdC
fiYGz3iTJsUef9DJ3TPOJ6tD/KpZyy3fDgHBmIEcy2pHeu5S9l256GMTpXciA4l1
+c5rx+Z2InOZ6zXRnV08+jlss3A0DelNFBtw4sncJgA=
`protect END_PROTECTED
