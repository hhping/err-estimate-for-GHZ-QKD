`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
haimAfmXoKTK22OD2x29WPuzA+1Yrpyh+x13kijFbCOdtw8NU4lw9mF8gZfTKOGN
KP/tUjoM5Bc9DCNzlsKyMnQBrklVyUebSAqh/69LOqLegsvTLu81x8wUj6vAFzZI
cO3I/F5cBjBrCS7yOCZy8eafBz8nMIi0kSV28qEU4Re50owBXitghiXBjd7O7xu6
b/FMO7Dr/fsQetJ+pVOSC7HBYRSWnFGo++9f5p5uUd0QBxbEs7WcU1YrDX/nnSzL
vPpXyVXTi6nVIn1je5Tn2Jocu6R2f7/T+pYNBsthkSEMShRhAOCUnQGkDRwn6puo
+IpBuqBBP1EFIAf6uPPpf0eRRfCkM5+UqKOyQHR6WL3uFMUieULCdN6N2QuAukOp
XTm0Syux6wmyFFCINcv4tC6H+ejCxD7Okl0nVIByZYUXeqzDMx/u4i9YlclXAGMd
3hFMsfy/ycEVlOwwqcPONO0pvu3CJQYwCqZgNSMTgI31DspaW/N7YZyLZoIBR5sR
7++The8a5E/XG5dQs3Emeio88KrxlXVF6lZjAFjG98ckeEabsLZf0y1md5NzrBvA
HsLdBWZMYrdi73jDV/2QaRpNJtisugqKbyz6Ps8zXc0Bxsbvnh/4kAX2H0l1Kb1I
6fLevKXUP+Rp6Zm8YpjIPTBddbo0WKv6afc4Fe1YqAx9Wo52jZxU3lo4pKVRmWbT
Rx1hkneiGTaMvlO1va6m/OVueqxtmcGk2Eib9hg1LJNrFJh86JNBKLGLuXNvNUO2
qu+ILHEIA9Ef+Zt2KhUAoFAjra0d4FUv53igE9O6PRlSD4FjYdB4aJPFajn/d3dk
fob5tpzWPVdsvqztqjjHJnCbEYa3hx7LosMTdoYRc/CSBqV2X44okmxu5I+nXyDQ
eE3SkGl85R8yEiW51D6S6xPq3TB5UTt82DAUGYZYxLO9gn4DjmJRppl7JGDk/7t2
gc1kFWIDAVfs1DeQ8h1qbBFCx7+rZgS//yB/ZEAtafPfqLEYAbTEL6R0qZoMNZ7Z
ZWZdMxnfKaci5662KyVPdmWpbe4dyj1+5TQ5Nxf/oTR6tev3E88bpIQw3cMDDQBj
qPnCRpWBVNzvndFN78OaWB/oPH9DtC1TMH7eIO3oHL80ZrGha7otVn5BrDQKB+77
hDuLEMnDmvyGTPGxPTlLy+SRHmvwMFDbLJK5ehZStRYDdE96QBA0lM51Y4psRJpt
VpB6jUtfF+HlgNjdRnSyfbrG+AID7ebfPinddyFLh2ao+iXzOePySnmR1BbiFewU
d5F9n/KKnrpJ6rObhEGdogvs2vt3XIEc+1PCtOTNJr5I6hIBBhrx42JjT07PMpeD
Uju/bckl2ye5HcZKVuATh4cUMk3qSBApq6Vud0ajdRcBww3tlduzV1i/zUY+gub4
05qfzREZy6jlE9UXvmNmCIwnFZfbupcinlryV0lPE70EA7WV3vjF+h7+zEAOwNz6
0GcUP5WyV4O35GLAsSTzJxB7C72NCQpPWAyW+s9gjdJ1jVowZERIVFlOmv0kOYky
akBNwYh7B9E/fA6MUppIlGLTa2buH4P17JZtt3flD8IHiRFKgx5g8eHunTk4PYB/
ld/MAu3+3ZB+ZMQ1ZJioqyEav4F4RD/TAxtzeJx8wN5dCEDgwNmkvmJdhhw3/95u
wELjrh5dp8+NuAQWSE24/+ObQmY5OLHPByA/k2hjUVGxl9/cfSvuCLlqnX8HWsOX
7VDJ259+ypAaRkWlaJAqmItb4dNBTSz5ojSlE5Q3bR/jFK02TAvBASgT9watiHtl
m0cdLyloCZeubu6cl1DRW6nG0CnH98BKjoT7XsqPSWLK+FiOrBrUdUzhLGXJiwSQ
BSCSzAmYpL8ojTTxIs1G2mUKt3KlCcTaecfYOwyDIZ5U0sVX7MfQT8Syd6j0z2h+
DBnRyag5OthqJ3WAwmqpRtzeof8wafRQG0EcZDbcpRNLpD/yMXR2xrItIopn0Z9A
29eY65aSuizXJcvaNb9cxotJQqTs92sligXz+PYICcUpjsLn7ZgwGMgy0a2Blni8
eCtnW4/hFEYeRpX4JhJbksBdUBdp9nU3w1oi4aGDX6W+QkCvjeuQ/joj/HQm1ZS0
WX5EmOleMADfFAiVIZ+98PvjB8qMfncEmU1l5cgy3zx8LeAxw06FUiuYBVIaUKi5
rBCI26t4hnGn7H34xuqIsEl6r7e8lkmYwGdn7OMDRnMzkqHBl+tDnjtGBucSwIwk
w4vOeW0Mm2oyw/WIc0K3qrZkJjkjZNCT/ys5OqayLUJP9BKCHR25dh+S0/Q/HXQv
JLHGp1yGiDq+4yL3M7tqzS1NXTXMa0IMSyrJWBSJmQUt43/K/NHnIwzt9+kFVp/c
AP2Tua7lwXP7k9K5fgLIWwc9XTlDUHUKph0BlCfo3/qqUpuJ0lxL51r4Rij1aoEd
KHAycZwT8TgjPQDHzbnTg5tZrkgLYb46Y0z6CU532Ztvqk8GgcTMWStrz511q+VK
RCrVkLst18kvXD/fKFV5mlgyaonSiWHnuxwGHFhH1nkByFvOYLwNNJAilRkaHxWU
VU3PYH1zWZcSIIJmAbATg0gy5xXaOvaZBuimE6uOdec7ZhEZ6Fj1LE3CXtn69/67
9/ijo6olwVCdA2D+IthbleYU1bNOtaT6fOmSaAEoUAHt5pk9F85q/e7tX5cSxLgg
2EM4gmHUIudrtnjbUtrPA+Rr+OPVv2qmIIG7322v+jdind/Eb23UpuleFf+opr1L
FWmrJUeCcgHHhEqZImIx7OoSlDUt7KP8tWnie2Z5SRvB3VIT09Hd7kOv9E4a0U0R
Gn48nu8EmrFMDaBAXMI1m43b9BtVmSQGrTc79wZZQP2kGHOyWMIQPdRHyFE6ospZ
OzCpnrWB5aCIk8QnlRK2ZmGPgTdoy0SFNBUtWc/XB95MD6crcTf28fGHnvrYpwI7
C95CJ49NiwTurhdAUhcL6X7CWRvJN3y96uweuvaG8z2CHpeMKLTLewsnfOWa0pN+
eHHte2T0VvTrixNXZkC9g2jhIHEaD5OYUonXEJY1nXWVvfHMjd2n17YzirkSqQVX
IT18eoYPQ8sy2blZ6griU09ugXJGjj4bfNTYTe6QnfEDqOqS+YYfwl5q7UgvexnN
SrE8Okenc1dDBUD8hLNJXkDB8YmyMHbtM8tNmgaAhg81pkVcUP7aYSelYLJu9CvH
HsBIhA14nfyCu3+DKhlY35hUJrrNhnDiCUOXD4NI9p7y87pi/R/q581mwh600Pyi
30XNWDvyQx1rw/u16px4AjZE6wHj07x5ot3GmAIG3FPLUiTYyrsjGC4VOdc9fHYC
8qPMTXqHCL/ilwJuCW4T/TI+CNsRTHzm7/zYo4XM9UXGVbY3klbFH76rpYsi7IoX
X0L3eAsViIBS0GhadszbruLWXMlWRdq3jnGXHzNbJZJp2RTbEB60IKGtK/CMSPue
JP1hsbkpdlxJeG024eBO4mRvPoY2F3mhSbX70DxXds6hAmGYu3lTjKlz9DmNJPov
7JGgQCib/2IeYBy0Wn4bjlnAqqUITpn9TCZbHfoemKG/qwt9CebtYEI4POQ/IKCY
io7BUjLRI7wn1m7umnIdIXg6T76wNSg8QdszN7mVyqzd+fP8aE41v2Nc6BxGkZNg
dWLM/JcbskkIaSgmPcPUQ3MxMTFkKx+zDUPPE13oyvfJgeELb9nhQQIAHfdToVhI
WkguMe4OKguKsECRI380VcM1OvC+/UFnUzLcDK7z0OnX+AdrtNZM9ic9mdamYy1x
aekFzqtd+ywH6coQCwSRwNh5mzcv8ab636rwG2jsK6TDpLXi6CSmC5p0wz7bIdeP
jPQ9Jo5Ny48lkmTG817OpSHCXRwz0QlpmauOFdejrPAWHmWnWFNM2IvGO1YkPCvF
jA39nbAjyMZdm9Iohmo8XdP7QImqLu4EPMSuv4CiOweop1JBr1mGAdutNgLP07Gz
ihQbCuzTnPJZqjbcR8JUjuIr37hhgc9V8ImZcu43LEjVxmDvP6T1HtNuPkyQbSPo
ZHrn23R1RdAYdo5j4n00XRod6ekunyv/qXFSDjOvAcv0j0iaCWkE4bNZoIRbCqZo
X284McmMzUg4ghdVnOiO94QumusSYgcOQ3DIG3ePT59Lf/FgFzyxhXZVepnWXAAn
J4qqeFt/sPAME8LEhPLQrbh/NM/1C2IhBRDZNUYiP11Kt6lVX/AwPKiRLDNg44yz
YNpwcJGUYBzgFUX9ulhHX1En6qyv8WfXlQk2pkO8Wb8U2MlEdOeCQ5VAaTw22+/p
HacdfW59MHa+fqg1RVdt1F6snN+17OKT1meLEKzMc0cqXfV+d6/ycp4DK7/3rw9C
DftZABilii6vp0iWmr5J5PwICw2aRgc6xpOcFZrBIuBeOArlX2BizjJeSM2yoDWo
Xxq/1ebyqX3xQmuRF/yH2FjgQ3GsMbi2U5y7JXqy6YTd5jm4FPaBvFgxLFLWJiZ5
BetEBAmXnqEidb6gWZVmq8R+BJRX4W3zthF7Db4jz5XTr11OJsVm/BUplSF3cxH3
hlwGpmUB33lYwslsbwtdnSOSQY/gxE+XepdFmz5Po9JLUPJnAeJmPZ1zoCDhKhhA
HQowPPTfE8cfL/QCAGE/oPKBiqr7IMqPZBIwVgpNwlDsWMxEGSoHK9LJVpBCJ61i
XRMjPtbgsJYRNMY+qmDlA0PW8jeaPJ19wqJV3ryZ9ICcPXerseFD3f1t1xfQvoBN
rS2DjihIY/Vbbubmu0MR6euz5fQ1og2t9jIVtC04LBtxI4tGb0V2RYpRfYX8PLup
mDbOXFhrl7VeGr4JwpzG6mh3gSf5hWcmGGu41Uch1+/MNPi2wY2A/69rBfV9eRPj
WFK2JrLHZTmzrzMOxRSzbFcLUOKwg4tNLYxUR7oo15U7rXr80f0H2T2A/X98S5Z2
aUxftOe5kx5pAEfmKyogw/ObjUCaAHY22Bj8ayfxzEaAd4o016HpwjSGbxqTFOQg
pulQWaDNggrs5KX5KcAu8q9K9um89QBMijfTb/HZA+DmTH2ENmT/Tx1KP4DhSu3K
ul8FAuSbTScoGiUIy+YYkpGlLSgUaJVeEsV5eAeHO/h9lcUajL/neXmtsA6mncVv
cVPG7OtvA8PV9OVRIC1EZQwmHz7YcGmIFmIZebagjetyKFBt17psB9B0iu30A6Be
uOQe3gwh+6THgX8l7Ath/pPWp82fDX2Bh4NP7ZQAgvU0slyOz3dw0TpwNTONmQOQ
wePjE4Ghnm8uq5rEtcXkgO/oRmTmmA7G/33hnKIkLDF+ihUysdClgLj6gpSvMBy7
5lT1kiI6t+1NpdokdUjkQSSTtu5oR8T+HpXfnjVsbayShY2du4b55EFb1X5uUoRo
PY/317ZDEfjzZiwBu73G6YEoWMB1FdQ91rJNu+547xh+myecgwFB3O+An7lL+0sU
Bs/7uPI1+2f9hoy9rxjyy/j0mB2XgLRQVd+zc/vlGlC+1DLLLEND+nX5IqsAvfok
RFY4zjZ1pbqSvUbhE/spPffdR8jqk+xDK7M5KRlLVfATYktTAPXoVd8ejsDeZjYm
t/tkux7f+SPludefzvelJSxy6D81ER2kZqTw0u1+2gSIA9Gr8E77DI+cEvOHoPKB
8W3DTj49AEACV60yanXNWrkHaNslmyM9ou/5nZs1CKXtvxJlTuPg6tPxCqtTu5cS
s6ZLaEwReI3sQcS9vVvB70dJf5XpgCGVIyujgCQDg/OSaZFCeYN8GMNHqsUidF2w
9bBHT3xUV4ZtLE7Q53aXDRQfUKJHSnQMWTSh4nhCvjJ/WQ1cONzVwcDTgOw+06xo
xwH9rFkiNJlZVvLnTfAMZ8coNSI4SVldpiBrtd/mNIX46xE3nOJjkUZ/DRUNS+sq
bqT16EE4eNfL/4kYoEuT7BW3UDC6dUlltOv4gVdF9OqhehCM0e3dAvDhZVKOuxEL
wodjJ1N64fjIVpNBXbON6rPlTxz1Tzv+dz0+eDiLH4gsdaq+tShPDPcz7VMnYdIw
zUokVh+YlwfxNeFeJfapq7uxENf6FzpNEyTOg7dOC7Gi1W3dR1aLnT0GBeOwvn9i
Dh2O9fPUml1ibXVU0PX3gJtkJpAr94aADY7zVv5o6NrkLsEyejtzgX0Zn28RpvlJ
fkb7dzIF7PEBLVKoDhhaXw2uPZ0hhChbgnxtpZajC/m8usbBglRuas/8wRZmfrcl
NrJRzAI/Mr467Uc4QeBysR/F2lc1kmnVjRK1wgAVL08TKxRU0Mx5MvfkT0dFTvtT
qBvbcwparMxVLmlf5+RSecos93olB7mxUeACJzLwE/7tyb69vUC2M/1/htiNb/kp
skOmTUEZAHARvgvdwpRHLX7D2c90YUOdX9dn4+uv2V+QNzi55BH9ExtA1jQB5y94
1Im03vg/AbiabSy2lDhAbwIdK6SeA6BKIa9wa8WmxriOBazSQBGO2kK4VPX65Fve
FhnLRlgmcnb2M5A2wahD46MDGhHBASqwYzPw+/794lPWhd1xBuKARg1sp/mCrFSs
i9xKZYxRZlnjrqAycfmpbxy2HmvobmMEQ8nakicuOT7t1y3WheicrVQarhl2rfdC
xC+Uu7MVZcNPvZzgNSpcmkirD+lyjgA+ylaz4Z37y0hJP9gjs0bNsIyWa7DtojNw
rt7eguq3U/B0sls/yeNNKiOk+RtRsj7+hzHPUlrVLoezNqGRDyF+PIe1ZMN5jS6y
uOBQJZypLrqaO6+IKuhEDPCsSwf7Hz3lau36uZMlIfMAW8CYKl3KIlRtpJ/esJ8p
d8692+cHlnqlWoTKoyQVylP2mmw4HguSadJPeijoQ3w+W0UUBlTlTsAYRBGS31Si
+HQ1QgJrgfe+TD77/4Ipjqx60BtWN9DBUrskbBF73U+BACW5ECum1qDBUwn3iD2t
fBpQW2uZizxiMOrFpf7DLFi9iIhJenhvyZRKDcnhLzGVi7ntLtIADGDSj7tbhXRB
CdmIiiEQHVWUdCMM3Sw+WWpmhuGsGwwwwNBYCkpepu3hwuTatG6fou2wzIJKA8XW
lfdG5CMqZ2+jl3zbcnB6JE4x9Omzaqho8mG6+1JIcXijL5sc99/Z99BdMPCCOua0
`protect END_PROTECTED
