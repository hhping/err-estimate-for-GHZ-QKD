`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jFwu2IOZDtYT6Phl9/2vsN2mt+lshFGuSHtem9RdCCehsoINxWGb0vbT56n6sq8z
8dY9qNY8G6EV60czFx43GG7XXH3yF1KmEsh9kzQKT3fZVk+gh7hzuemdr5Tu4mvA
ObxN5dDQHQ6+bs7fNRnuJYtpG5S+XuHZcgRsJGKamOL3mjSnsa4Mfy7yLHgI8pjO
g5vw0h9g5ts7s4U6PFlRzWN7x4mmoduaJpi+drvoNBGpC+yAKqtjnthCuSotYJxu
MlHKJ67jQSlqUplLD305phJ9z0sk9vz909TRfz5qV6vtTXPweIiYbrE3NxcArbme
DvL0vPMFpwqWKeEEFFUvffy5kQCpM98PCy9AlTm4f7V9MaOftn6uSQ2FnpdJjZAW
Z28CYa95ArAORtksnEUPjyzep2y9Sj7P9uDohLYDlz7u4wVQL4xbpaXD6szwbsH7
6JZruURSOyxpyEvBjjQX3iKUw7HCPTluQ045CjNGcZUg21+Bbp5OEJIs6XtWi2aN
J2C3YmzJ8NoPGirPctgCpRFuY30wk2bbl5zxg0P9Z0nu7+WJWv1JjCPBCICdk0hr
PhnYeYU5nmKgcnyhVm57duUIps/h6F7b+2wvRXPn2cI=
`protect END_PROTECTED
