`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ytm8/WlSvn2MN65X6d798ttDNdpAK+6vqoSNQhTmmElBbOhjm7Gq1EJ1RCKXtvW9
Mh8jIoY7C65+3o9u55QkAUzRlUJ+9AifZ7oesEC9Kay0rGwzliotels1Ka4OsCFc
QRfrJf2dRoNV5l/6pAEf0zinBvLUNlHBzHqEIwe7i29apeJH1IGAhbngR8P5bhph
GTxn714D3JTtD0QxZCToaT9y9VvMxg3iFr7u3aWxpcNd68FSQZJmC5Z1k8IVGO6+
/HwuF8l55ujdQbP1NYo6NeWqbAE0YJdEA00vGpelpm5gRqgQbznCxZtaLVCPxBF8
R4Jwbc8OfQAQeDgO0DxyQ5/RzJi48D4V1hyCykuIaFPwobI3V2551Xb8uvN+5zC7
amKZPuocUjIW1UqDFVt90Nbr9X5Am/aYhCYLDDvvX5Nkv2KJ6HAPAsVdwelK4JIm
shMQPnR2sC2L0HVbCEaV8qv/N+YnBAnn1CTn6LRw079UCAJfa/swyAqSiSlBz+55
ipCYxA35pUGSQD1YEx2fh4sxraUthbAdQzxcnhqX8BvU2LqTMiVtYEkubCAaG51q
cNA+R3Ejp8/wdZbvdOdCLZhDCkVzAkdwGpzMemnFl+fIO208JHtnVWbCNqPTNgEB
w5MAOX+gt84e1bWmJX4dgBBti1SEGeOTm0rKPx0B9mUSEXsCpcXH0CpeLWwoDp3o
`protect END_PROTECTED
