`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/X4S7AR0MpI1kBG9/iYRvOBJ89pud9nE5GfPPo/DPEdfTLXtt5EvxlsIJMAvXQj8
NlSQXcHz+rqB0G7sIhvnL/5Kl7YjsmdReLxt8qI5jSnpmrHKzbxU/9xz/wYgJtFy
h2ewgiXjrE74T4HdZeqHCz2Zm1Wr3vVKnq+ddRWg8speq4tAIQ69mADuzCNX/wNY
9zJD8DjPgYtg87xIrwXSLwxBeVfR7k7m36ZcFAq8N9K1d3zytdzTDcmsBMRByivd
MpGw6n73QHedaxkoB5HLggPKE6STToDlVZi52PdylEFmo+c+3CLYtVf5Yh2XLczU
2DEOcCjCE2/hlV2mAl/a2PhYib4sPhnoHIu7a0cEJ23DPrq2a3QLosCQN7MvVlFG
ByCLVCCRpDH1F7+W5HOzzpmRmwbppdmWRNOh5kbgQPuVNHQjQtiZ6O0eaPj7neN2
DrYIKM/6bhI6ZOJ95wGyorN6jvze8Jizl/XWj5lf6JAYfLyu04Ce7XxAkNuhaWu6
r1+nOCywIRqr0N4gkJTgClEs9Eo7hJxEgVeH7so1Af3JLX/1QSIJEVWayikFRvAU
DXIRcwcrQ4yOEvO28qTAasGTyRo7uwcJTIWXHFhJ5OndMip42MpsT+uQvNthSlT2
rzLK9iMdQJL/HW9zroKYsbrC2nEZj+izxdW+uj8WaCzANIrI1TzlzLYoRojRJKEo
kcs0amaak7ZQm9nIFvigyq630ExWwD104D0ngoGZeiz1qJ/BJhkjUvzaT6ZguaVO
c7uNMiuKDZ1rE3pl/ee0CzlWZ8TQB7KXiYhb6de3Qy/uflvo+KCj/mO1PAffbPE2
tXMi2QFjtVsqzTtSv/6Oumi/UwQScpZvasRnD521CZvinC30yoRkJyCjFA7Rgdu/
/BLQuNd4iLUOy47PhBAFXmzIGdEhFqDG1TTq2LVfV2djg7+Yg3NE8sQRQ9tzfegu
AeeaOOE56zel1q1/hXRygDlJYasMPmB5CQJyfZU65hSkn0sRcLeHU2vrJyGAKnow
w0Vq2zZUFBcRTWbeJql+2MFb4+5C6VvL8rPHDXkr1YbUmn4R/wj8VX/EAJZAFG0l
x0ZojKB9NQG0PUyPDVKtxoAHVQ4iLmLdNjkF5sH++2Fb3WT0zgZQf+RLOw0lLytD
6t0Qhun5hUYV3IEsP/KjNimHPKlY1S4S3uaDcIlae2B8b7RziQLitTXsrhKKdul6
s9HSsjCEORFQvOgVZ7d7q0Msb1nAppQfeqcF4L34wpNx+XcFSmMiu1SiXAcufX6q
rfA4avsFr8/ZOWawJQblu+kuX0/jBrtpesD7K3ImkZKU5jXUhxvtR1SEJniCjnum
vh36WyhBbHwICWEzztC37yUk0hwwGbdmYXMNJtX/RM9fwe5VkyDuk4exKgPzOrSq
XDczpoFyK7uZ5OYF39MQgG0k4OFxwgBzFILlSbgkDPEioMAL5gqCGPU8juNeSxJV
NK8br+oDvnZYbdmOqCXZwJZPmSkIOVgInZShdtL3zhfhcK1NzGnpTN1HGhrTZizD
WbKUJLC6DY4EBPS7oyhOdMTYfMk5nmenG3lPmjpiPgCdnDGGXCGbFypcZnLAJqkw
abv713QaJqaLtp14bEhCypw14peRGXC46qtrt8kEhXUY8i4u1Sqwm87QM4donMEb
nMzqKL1qpNKLFUI/98qLBtclLmZU1jcyZLekJga3FDZAUFe2VG3gWdhd+L4YSDOo
UM01XgX7FG0CyPMB5TA6llHh/m9MswbqPUbp9HnLDt1+ySSVEP2bsw9ySWsByAH2
QNlO37ALQQcSnJ5x8lB0sdlmJohSW7QbUA2fHlTzloElFhcNV0sfjeOHtJLQtNkT
Kk+zYzDUfm/Dx1ZojXlBObqtkrpqSMMtg9hEPy5KpJ0Qp7qRBzwq5yP2nYI6kAq0
TgX3XYScAljNuvs2k2qGV/HJG9QRZBQk6s90bup10C5fFtA47CbKH/fK1hGHyBHy
s2lxYrDfriMxO5mG2UX8CzGfElZaD05noEIdmujf8gUJn3H+wwAgYMmnA9E5w9NL
++P8HGobxF85uMm4/ye0e4aRAWHFZ72eq3B8b1H1IGEBISVfNNTyxhP6mYm27lay
T1Eoa7eAdX94qzNy+baSiHCmsxPqmaf59KQqOf44kyvRMrUpQlPkUH1TbGPssPRi
GQuzf38MSeVaVygMV1iQEmH/mHsnNnvMrU/+4HH3/uOn821Q36YKULcn/3qTV6jL
Yy+x2/wcgT6FEaxGkjFHGb07v0ZJMfIWEpQtAKi+J/CUvKv9ptN4LxmPGnFbG3NB
aGW+3ziK3C6rYgeP8hpdwcw8QfeiiMCGRh5rwUxqRPu2+Wq0tC4FgJfvAuvzoS0R
jy+RV8fu4bNFve/l8ZmkgmsuPzC253zP4CJKbHkFVHD6VXP3QxwRQysDv7Tg7F4v
kiJxXENJB0FvziiOTFuKWtV0Ck1y7xlJhTzXerK3PV0/L8jw7OCvUEdF3lznXqM4
/x+2O8HBWpOrPyorsSPhd8xY8fdZnFrGa5IJtU9vbaX0Xkl5vwKc8AZ+CyV9T6c3
6C3u6H6zVFrit2U9M9Eu7KOR1/FSzgzjYdulDYqkamRqITEXdpHyicA/qNilkCKe
v3kIsadOc4SurSPwc6fgPqyASIF1il0jJyWvDKlgp0+PjQTOQB/TiLy+ejyeJV5A
R94K5chPyDrJNVBFejIoB68qnbVo3/dVFiZlT0v5qpop1oVjZ0o2fq3waUqv6QeE
ncZpdzT/FdlkJCQ8kRDmX5PAVu9jvAcGzaDcuLMgrt0weIzO7QcJiUzhg/PrMytU
9uSbirbKBUP3CV/cSrTS7eIJu+dkANCYizw3A45OHOmQeb5/ZT3/aKwEYNWXn+Wy
S2xNY4eNT3hg5U0oWzlUnHdI4ZjyZccIhK0/EgjRJEuuQBjuZlIdt6A26rCTdx8k
7RcZl6gPc3Malw07/TOmqUSo4sFArzEghlCVlE9CJOPiD4LA0SC57n1nfD7PrcOh
ZRmliFH7Njf28NjEvwa9MhWz/Y7R4NgeVEv68FdTx8wdkYuoyutX2r99VwEM+9ca
4fEIk+6Nu4UNYNaiC7aAOPP6ynTaoAmzlqEnJcl4huKSXUR3YfCMRWphKsJL49ry
yWhBz9x0wSttlWsIEi+zE+ExwqkNweFsVYCiilg3WyUbnufeOF/bVvspvb1VYW9W
gYzyXpMyk6X+s0Gh9Py2SuxEGj8Ex6JKlE+7HgiTkBa/uDjuupzyEjb9Oz29hHxT
UBBcdsAQbE8DIol+CuXPBSOGqTUL92RoCRLsbq7zokxPAp0o4Lg+en/CYGrMKu8x
8F1SLGLrTB4AzyBcAci4vmbSxEzLnbcw+MvSNojuzX0ae75fVkMXRrIsgjSH0vKk
`protect END_PROTECTED
