`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kAwv+CKphh0cxRxDcuP5GNZSEAEiLtg5Kgj46kDitFZcbLV4xPQ6eYbt0cmUEuOj
i41oG6O3VqEi96sv9kK41yUxYcv1js1ro3KkI+plfd72p5WvbVKHh2+XntKLSWwQ
arXzWUGHsIMw11mSIOqp0+JsBbiYUX0tlUEYLUEchhjZ0wwx6rCbfhe4YL2fmyeh
+RYtx0suonqI33uRSSvYemuCkEU6YQjXoOE20b9gGXJL682HmuS2pjCbLO9tCZg7
v/zELFGzva7KlojbBhqr+Uh5h5Evbk55UE9oS8+UiHoHJcIwsDnZmhHXwlm1X8dF
tW5OzQ2RWRquGM+b7IQalRwyivMJcbvVRVS+1wFhnzfrBaXY6UqbPoTdZn2lgOAr
NFwNEftFSGrYQx+aGQ0K8mQy2pjCS1SjoXi7y+1vp42/9hVUuwecZJu+9dSSwBUY
aMeyKruXxZ48gPlyISpa2OxL+kvFhErIEI+ZBFgKV/r9IAkaoK3H71KajLUbW66Q
ihGVslyIO9OR16CgHhS5yJoACqhIPJv8CgRqLNgySA9YtHXxRPy76DcnKA95HlbK
Grt9XWRH3UgIjUulCR6vbarRn39LjHUlYTEt1g0KMiTw6SrEg2iG8bOGPH1F33+A
L2LUY0rUTcYgBQsEArEzszoAnRkWzkO5GhZCXDUx3t2yBDY7qScswaDEMiPcqz+k
zrsDYBxEZNTu62tvlHDpWa6bn/cw/lz1HUoSwDX6tKtJ0dMKF6yomYSlPnFmHYtY
APKnyeXPsCLfVwA4bN0coKZjNUutocQMgxbfAerjKWe5+Fp244KAVir8tXA7L341
Fjjc7uAu3lbQhsUeZYlLf1PpMrvCgaaEhD5AsSAelve75wCKNhAk4YZHGY7ljPZY
7O9VtXtjtZin9UJ2k3Veyw==
`protect END_PROTECTED
