`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3rphfAjBaR3Pl0rvvZ1chwgjkfSDinXWUwzkgp1bgJCCQBuDQcNYpmBzS1Nhpi5J
SAqlWVhNavDdk7rzXZeGl4NCmjhEsZxppKBG9c/ERYA1aLnOv7pBw/gw/B8qSTQj
RJ0aPZrZccumTV1mKpPwx/uJya8hreiWSdx94Uevfk5HzECmy6zkzxsCd2WNA7z/
1MNTyAeNFPelibvCCJvbCMATTcMIXfAj9qb6MK8smRi0lNaT870oPIQItVTDrdmB
wk++8bRhPTuULw24bMusLw6h1rCky3d470qpCygUoSBauSLl6x3gGeipi5hZP8pd
NkwXm8NOvYhOq40vXwpDIwOVtjhXtUmCoZFsnCiwUpOBKxrCJ0/0CRhFjXEboS7E
ULOYl0VlbnqIdB99Q2DTI3UupgeEkZjfvJ1iSn4rTgPudR5pjDy6JtTL/bZwf8QI
+N26uRMIo+s9fQs6/foadg==
`protect END_PROTECTED
