`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IYmYMxI5n2q4AsLjBGOad0CdN8tj4PWF+bsfZPn4Gx+yyZOqh65GicCERjC9RcMx
17XfFjK9cxdfYjvDhOcQ5O+7XBRyBGV58RnbP3NnWS0DYh2GFocl1wPvoSAojcBb
8F9N7cMU0TacqtwNquRdia/s0SyxojzMrGX5iyAswayUiQrAq7uh4qUdxkKkEuWh
FyZEiCqOU1K1LS5CnXQMWb3FterXAOOqvb/SBuQMExhnPBdX0UE9m/bnJaH76JOK
3b+e6S5oGCVgWjAAD98eOV1qd1gUrM6YOieGK70XS0o0VptGeKpIuyD9rYo4pLt1
NKfFjDu44d2LWByB1GOeAMM0nRiGn42BD5qS8BfpOM5Swvsr/3oDwkSS/Opi4iVi
qQ8LTnAj0jk6vInCEAnxAub2qlx60LG3IrttR/tzNgwiJV2G5/GtU7FMgxs5NVw8
kfXveBOCjkyq0sXxUlIdhmIuUFGUieoyo2Yna2dSduYDZxD6x2vTAImFsyvVxYcU
A4JILZgFKhqELwrx3Qp80TTQCTOGpi0P4VikH3RiS9ux3iEwpdAHhk6VjbC7gO6G
hINHTrgoEbbVXLCEp+JazmvvMgeCu/Ge/ggJMzF6J8wbk0AYK4VjpPMiD+7yRRm2
kfgzrn7+OKdlREZVOxSpuzgtfavAH5z3oSCsTmI6vgXlyG9tbKWpL+4o8S2ml+Te
WDGcX7HHdFugkV5DfWt61H9lsCbmSvm5a1cAXiyzr6kF0ONlTd++XKJrz7AGMkpB
VqWlG8YWTSpL5/CmVYCngBtdKm6tXuOnJo4mAf5OG7vtMsNlJiExBaQ2sPpuZsj6
Tpv3lX558w84tHMJ0eQlVC2YauSYElrnE+Q95XpUADf9W6ymo1duTpmCn2zk+Rft
1qs8Bp6LdUJz7r31mWSx15WPPHcOekW7of1dQQvusMJBrtCZmLvbpeGxF6rYUBmn
JYJHo6mDz1kPmFhAQrjJ+h0ZvxBKBs1RReZk3OgpU0upMRddzE+mU9lB6IAquuMK
qZ2oAx+FvKNBEzjIJgXaPdirh+b5/FH4MNQVovdD0Mb4jExjok2cNRXsKzpY+8rX
8d57zB66xhJBNJNDHeuv+VRhDd1Ugl7kkwVK70JPwZ0vsseSnW2WomAlxmNfIAWP
xNfbko2JF2OGmFRypZ9HGiMJJvNPZueHrbpFMeoYiR7IJR1B6MFEgb+svoHZOgGC
s9QsGwrr1KsQPTMLpHXnsK97ygmrBKO+hXhuMPAZ4J2subjb7GWm4QWddGL2x3FH
z8hi69rxtpmwM4TBFiqaL0+TptAIdJ26FzsWYiz+TXeMqGn+mxnmJFwmffERKty6
bNHxzXJdCA0cEXMz+orsy0hZ0/0UPhjnLiyDEBxDY9h16zRzNlqvYB3f+kyRvA9f
5W1I9BnOWdQejEeBkdQWrdLGQKiCH8wJMP1TeqLhZyaTpJ/GYt8D+NYuEkWl7HZY
t9sdYbTeOH2K+2RN/wwELAYNbj6nDZ+ZZsOoyDq9V4YYBnjj0FMg8Xstx6mVixkk
Kgc2OcFYU6Zw2EzVfsnFMDsmVMjYaV0NKLQRfe/wWodolK2wezZUTrDZWNrAOBw/
i6edu4FBcSKGb1I5Xc8f7A==
`protect END_PROTECTED
