`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RJmxU7wUnTqjO0lW2B8qHAm2siNbvAWIXBYZrzReIpDLONDeiA7BqSeh30rDz7RO
LwpTKDJVmK0zTnjD8/Pf3mfLe/MH9+oUKyKo02m7PVxyAeyFt7+Dhio8g8qBQVeF
vyNz9y3vYKBOArctLYt6XRWmexeCUO4JHRZYPowkmtwujGoJhBtm8W1sgYXPXWR+
tnh+CDqZYq8UjMXxQCqUwne1lCneI0I2rht4+0jEjOC0nof/SD/fmm8blb/Rgo9U
EavWms0ZEQM/jD6OXCay45kjePgx5z5RyMEAtFcHsnZSnu9WatI96BMhjcHU2U7I
kFwXDjdw4dPCL0DFn7zo+tatVgy0JX97U0whxXxI/6k81gGGFRpV/5kwMpVRLIua
peRRl0hK6J7FBJT0ND/LkqMiuFZQtotlBRkpeZI7LbHCYg/yit+GaDlRNljctMua
/PSlEivPDqLaR/6pxtr5cTQJseeMjWWzxrm/z4fV5vk68nlFmbJt+FMGY2fAc6mx
dD+znR7UEJXfbAGZMQ3ysGfN002mWLVhdym4Md+YrT0mycJRJick4+dRdFk5ZTcM
aKXdiUSefs0CUGRXvxDusUk/vt9rjlx56OOyQXanozT5TeRa6wmuhma/t2BaTdXa
2tZmlKDpxfxQDPSC/VHGGEWt+tQUyXyPP0saGIChL9/6az9X9fm20TIQ0clydmfm
ENLkWX0+UQlEyIBGCi8OCzUxBaguqUMtB0/X3u48AfQMPZ9ZShR0sCM/8lDh4xP5
sDNz4SdaY7kU/z1/Epmazg==
`protect END_PROTECTED
