`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d29GU0tQMqa+N4rtKM9/hVcl7j7zKOG68VqPTk/Lr1ycsskID/gTldGfYK9WZqPJ
ZSuob0zPKIxp0N/4oeOgHzcrLYMGH5elck3kKrldmuqr0EbvuekXyVjF+6Xpd5CG
dDMbKPjcUW90P+nRjBUIUiFCFKwUavMgVVkbK9LbJKlGyynY0HQUK8OgPa2Ki6bf
c0L8zIdQyW76s3tSbO7F7TYdwVh0NB3WGe+PI/qK5pWcAkBGyRozaq0YEdMqdt+U
JgIpe3I2R27zUu+vmTCen/Oen7Vx4Vh0Tj2dVBD4qdnoPlSuV1et7NeY6jBqfwTv
Z8AAp+s5JsEbDTzAj5E3gEOo+eDRauAIzi/iDxobehLGxFesqgWfmompuzWoWMPA
CKOvjQdD6J6mxbvnEj6cuq2g268/uezy5527RNqC3eIU2Pjzgb/yeOdDpsrTOH1U
5FNT9IT4k2Ez3wZtkE+g64bHLHt6OVZq9laDrGGV+vOGcXvrpvrgCyEnHvUgNJ2i
CGUf7LsN/sILpakr5v+bVBeDnH/vRJpKneFMakQj/wgtZ6hAAZPCPhCAGz9wKYlZ
nFN5FHUbT4ZTdaWlPGhbEY4kmM4Z0W2Z87V3CXNX9dVFvgqc5vfZvffhurvsGJKj
cn6mEWFr76Kv5/dUIwacK8nWrocgC+RN/ZrB8AsLAisTINfDdUnLIpSCvt058CRm
3O/JoQ+jsd7eUqr1ZghCXhSgKncj/ONKaMRqKrF4+Sndgqdfx6ts8RVYOy/LbLTG
iz7gW5QMYn7aWEf8VvzYKRUvMpnGpoFqQm30I5DPssDng+DZ0OlH/2oXnOaJ6n/R
G1Bo5QqxpPWXoV5Sx5T2BBX0wzNKEViZ7taqJzaZoTdh8CfUYnfuqt4RMnqbp8OJ
/TwpBYCEYRD84qQ+oRB9Nty+IMBP+GoD5QhM68IxIuxsYsqL/y4tbCg3RPk6euc7
X+Vm7gTaFFxMp7LV+GTaJGS4/L22cU1tVo6JwBvr+zsvtdhX/jhFIq28/MA8NVzC
BFsHtsMwTe4eYiB9+szS3WfZiXqHIJ8fIsfSvGZ83WN7zpiAHcW7A60OQ74ENIRw
lu2s9blEje5Rvw+feIpcesJOpSsIFq+oMHeIqTVOHDYZwfyqo4unwRXk8AjtL2lD
Pcb/dbMEAk6lmEKGnL7uym55r1iWzYe1RD/Yq4f1K2UxMbCPjHhlnEKLg69x6DfS
WBRYQzklJUMR4oqk5gL2H1yycxzpyPHCRoqfaUX6oU7EIeY0+oAakLdD8RyjTU3I
rpjVWAQhG13dMS78Yw41gl4qkoNBsTN5cv/Ff67iUz6NeZ6yM79rcvVYZM1LuK2f
fn9Vpuajhdupj995BhsKw4YwbbLfOhC5ogHVtOopNn4=
`protect END_PROTECTED
