`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hgFy/dkxfYclV0TDP7SvyxYWNejqD9uZPqfzNYXdhf3y8wiwHvzEVn5FcdjO1GiG
3qbSr0HW4J7ba8Q2w1jp3gL7Y64Q+rXzH2loj9NTZc79i9u8brn2sVQf90YQu61C
aHPK9iwJq9Eahk69FBkocMB/mruZM2broAtDjwrMpd1JSNiVM6LpVgi3aucZ/OX0
`protect END_PROTECTED
