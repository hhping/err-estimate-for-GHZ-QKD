`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sC382Ea1FxBZwT6RH8cq76NvpA/4TICMeAaI9cSRbjyYt94Y7sTrnJTtdresIZsx
12hk4NK4e2MXA1LKd9Ga3drBWFVcmbkvTpX3u1mCGJA9pkngm2VshKB+iKDCalZY
j5vPdbzFTRxKcQ/kO+Hz3vU8Bcotrw7rC7Ekcxk6uizk8+36YHg6hMOeQe2V08Vq
wvmRiM11t+8O+ZgxYKhYgo330bWicngx7TrT7Dde5n7xhd1QUId8WVGPtPBfK0KD
VSACIoohkESup2h7ZfWBB3W9SdnYXKslfBMSRpNvy7r2c56FS5xjwDJ6XdzLMA2K
vEn3umebEsZWV6k1StpzGZeE0oKvNFCx5wW/XQKc7ECttYyfA1gblT87I0IIz3Vg
ULJjpdg79+a2GT3zh+/J1EHqd3+mQfCYTqIptTOu27oe6IUY/5IhPvnR2hunix9n
`protect END_PROTECTED
