`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qmp9CXlSEt+5RkRKX8bKiLVh3mu91qQxP7IjFOGpdNPFtUmIeLcXEuyWf5gKx2sq
Gni3G1nrueoSbf++EweeNNjDFDQ2R7Ly3hMUShLgoRAMIRxDGKksGFvZ1WhebK4E
kf6h2ZhbHZHdEcMGI6OSbgkYhR8Li4hNbU06Vxf7lj2qrpx3+BqQF7P6vhzwaZ+O
VhseIj/raYKkdGvFVmnb/V6vhH6xms9Iz8fjFDZoEGEKNV13wiC+NLqusXVedqP1
HxvUj693RgelOKUMIUPkGqABojExJhDlyGnL5FxPDpsrwf5uuVWjn/Y7xJf9eyt6
vzxpCgbYdR+X4QsCwCJ1XoMQf5bgYlp1SBoInc/bvEJsyX49RLuKbmUc8RADPDku
zOkADDI9vbtN3mOtwofBouPGBuGCC7E29shQtHOEPobk7KMa8md/u4jDaedrojHV
6vPFmeKhkZvIrY2NQVAYx1dHgXuTVX+UkRBm16qjaxgB0muGpTLnzSS4Km5Gbgvt
Nc5F4xKmOZuVBii/ROg3Cx5UKcoGxaaOF1+WUMI47exquewJIQlCyCbGRrJC+jm7
ZFZ/zqc8Qhu5nhly/7G2yxPNahn+se6KBZqJ+QRZh8QKf/Xt9HLqsxcF81nbY9zT
NjDrYAA0VSGaSeaJ4TaC07pphIthWopSmJQC609relFRnXaZlfBKip349Ds32kKd
wmEBZiOd3CW0uj1IXi9ikgDNij+1HGRaKhVhr0KVzTaEPa63HdRRB6BzRktBYFMt
H5+WFeeMLkJtWOvC0DDUQ9EOUrrjMCtBu0muPHc0mep9qIz4nxEX7EJ37UKDr/yg
g7hQPiKgJskJXTm8qNNeX2ApxjUZhFF7PxQlrMsoAvdyp9ZKomy4psJ0WIpyPFGn
bIl3kcdeQQeKGuTTIoOUNWGpAj8g8Yz+m1BOCndwbuCb3EMWN4LbPUL75EojrkDm
dY9TrXEXYW+voIxwdcPgZzpTFDWNGv8pM49gSH8RX9w=
`protect END_PROTECTED
