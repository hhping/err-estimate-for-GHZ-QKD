`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OYizvymxwuLThv0b6p+UrX8+4L+DvVgJ6kGUdybQh292REdsEw3FakVUE4yZe950
WnuDhwOcGiYqdFN+2OaHJwXi65iYcixb9Vwy9USa0+5bDtNw6jCd3JyBZEAvoS6S
9msUdUMkq+ZZfQvXfxoYec2+c8B1V9OPZaF/ZoR7B/IOQDdNzpesT/X+LcCfjiUX
ReUik/CeOBAO042USqhQnLelb7TBMBcYGOyBMCvMOYlBML7ruzIs03LoUlwZ8MGi
Dy5k6YhK6s+tR3cW1cBjQxjQYBkoY5zzeyek4cdC1Xu0rA4pBm+E2M75cpAxVfqz
Di3OksVhczMNw1OYalD2+2NlpovejYHSJdbSTSPvt4uGPB5kx7Q8e9bbgzq5mOFk
i2JCDBl7uWPF5JMUPaS7h2C9jwdfKoSJqwahV+mZaUc4I47iKVPxdjgBRATfD9k5
kmW+fCbbA4I3/K82hoGdhCwsdozTjV6vdnR7U60wSyrF0PuIwxZcoi4mXGKGz0Ej
iBTf/e4gO+F6jdg42X/L1eDjBB63XH+W768EGW9NtOC9IwgDwydkET7QWsQBp3i4
9un+XxpGFM1qVNivnpJJq2JQVc0YV6vH41NAa3Bq2YbM1LbfP53k/l4z6HRwNqbn
iWdu0Cars8XOIkSzQDBB5Vqs/Qqai9aeZ2Lho51SoS0=
`protect END_PROTECTED
