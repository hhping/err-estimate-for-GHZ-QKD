`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Fh4jw6xcl6+hPWc0c/jjTBji53w+N9koVjvFf47EWR6lV24ch1aiDOajnB1z6l4
aYpMovpNWGcuiefEAPkGYXbCzMCruF5EKomgd9+37TznfSQFNr3QmKE0U0rIHOjX
TdAzrYGWSVnzBU5aCdQDdYPi+qAQmH76IlYm0VjtP50KYmGevAPHGMxDSqAzzoLG
2ficyzzNVgwb3QIzuKeMi8O+Js1jsRGE7HDeyHh/j0yblQekO5Prmkc/RhVXPqlG
ieSKsv/8FSsB/6YsGbYEg5kxNEGdUOD67FgUBTMRRHyVWOM+1FyWDDgZqLQm1xtc
XwZu0SPhOAWbrLZ8b4EoAJI5hPY4lM+Kcz2uVlLGcZVr2qnRPnEBzBY6Xi2njLgP
s11Y3cuhQ0KQG9eVT1sUuTRxRMwF+K6dY8L5CbmTafF4qVbDZ+veGeyJFlQPOEwE
P/7pee2TqlSq1F1PH40LrejUYcaZT9BQ7T9WEyFjcRvVX3Z7bcx+gi6Wd29mXmJu
RnNamj2JBjtJyDDV7u3hQMY6WqR67dDToFy4CUvFUj7fpW9eVQADezPX0Hlwzlnv
8wDBm5URn/SAdFq4O6tU6mI9CiqlBZlhgm+1lzDxNruxzspcqjeX+1/m+zJTm99l
VX7pF74L97b/Rg/aS3Mof3S0L273h2Rn+hhpIs49oqCKmH9rXWh3hp35GDRXzG1H
dDxj1I+O/u23rNo121Um6zPxI+wO8FXMAcpJGcXJMdbhmWKXyre1evu2TZg569q1
`protect END_PROTECTED
