`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AOEYotckLZLS44DBRJEIGidK8s4TpqgSqsEphl2PlvJly5eNZArjz6Q+wux0e3SK
5hr2yKCy1QlT+NV8vCoB4I7WVEnqqMEH3TOueK/BuX4V7tqGdwCxjmi0pJmFduEI
H6nVA+VegchbGCwXNXV9gG4KyXTEg0SzA4yRuJ3vJoWpPrv+M7lz4yr2cBnIj3wx
UZ2kXR/IOlypIbEn4bREqlA9dCr5G8CpA/PZ8n+4bEMwBujf9c+L4+eV20T8Y/5k
/5uW5DdPrjvwgV45ngEC9KUIQb1O8KmNmBr907HK9QmNs5vM3PAh8RnBMkd6sSDK
QkNSY81hvz50B3em61bfHVs6bVFCjdADVpaJcyynZF49zKJxEwIvqOoTF2K3B0p7
kfOkrHjD+Riag4C4nsis5AXTdLagThCPkRiTaLfNrkqKsc9rVexSE+2PfINvYhK+
wlUEhw37KJ+Gui9d+d2GjxWUHGLfs3Ha1D6+q4rylBM8cI4sD+FESmlQiQikGd21
hzWFY5X6+ETmbdSZEkDv+FigqUgW3pmwPF4XgtBsmmDopPVptPdX+Y2ERI8LHRaF
klcEsPjZHcEP8Yjqi/Z0EFiSl4oTM9IoyN1bWK4WR4OybDKSYjojM9tI+HXmS8dG
tmIvS+uzpGhjrVNmfcYgWxvdC8whf3x9lUxE5kEln3qNA5T81PKm7lFlVuq7moxI
8ElAjM+NiKFfUgZZDh9VGFaf1494uEqgdw/fF1Q5Mr8b+gZNyEW4+8fFDl4Sd+uX
Ja3CK+OdVbJ8HXApgnYA1UMVUehKCw4zHd+sYM4U3DFePw6JJGQPQD2/nwOUoton
Fo+gWBwSgB64vfOSq1j+WGdWT8BpcboV8Fv2B2ermJqk1tfUXJAop4BL9K8AJOfl
Ku1u1EfkS3t0ttiyDMPReP8Pi5jwGNWQxJ5CMLwATu1oph/paXHSlhm024gpBSlH
bfrkYzL0D8zC2epLgBY5+iH6tQAWtZR0n4yg9ULhHIQ=
`protect END_PROTECTED
