`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vfeMIfs33N8/Ekbc4ZnOoEOkC5Er9TjqjSortpNnEwmXCAL7488ASapLLGNnT7SF
Sessj3Drs5jgUDPrlKrlcnaUpMfaYwoLNbG8yuy6HGomef4amZ//erXa8s87N8My
q9l4ZS66faERkVMnt7gilyFCM4ZnsBRm5YOuXmAQf3LaSCHCERLYSDUaFtrFwXpv
GWxGPEhEAREPJnBDMYKA0fpzsAVfP5JJBIS9exAdeIj/cy6C1YoYxFnV1Cv1hsf+
YogbIKNk9yf5J/RziJLpIYFTQdfenVo4rqkccP6h9VRZQnkhTn9flZO1KvwsLRDW
8VVrNEA167csC1oAVR0s1ihTP6cGkHE98SRqglBgGse/elxyyx8Sn5wob+mYH84s
SUWR5j9vHdRmTi9Ivpg4M25U/YCJahxSXpE9TRRPqDZ7hPuxqpL3jpmb1uEK43t9
eyvZHMfuAqjg5JaCa8v1hsNmWB21+LDpYC39nMNWNxM6JYd+a472zc4Scy90s4Le
rkhT0nY0cJn4qSxq1Pg6zqFSxin4vwabb/PF3bagzmKULw5R+eouUI7GWoZNufQj
9z33U1HlH/7++fR88RI4phTcrVNfzh/td34LaBN+BF4EHr8JSVSx2bemIcQlCPfr
5LL1CUHB7nc2dDE3dLmDWnguJO+0jE3hqcP7xylQ/ATPbquUTMde8v3KaadGjz1B
HHIjDj0GamIY7G5zXLrRtt3kCX9TOfqN7T4CrUODeQbCCZLqRs0cCxTguwvzYDQj
tku+hTusBL4fEuS/PpdnC/E9j/3STC5W1BxMcHwVfHWkKYAVNwgfF70PbSLxyf+w
ZgSS6OSlahSvn4aLXFXpeMXXlaUjwQ2Y9/HaNvuCOVB9vzKzxPAKl75jFf6ZVkQr
ZE/fBgLxd1iohHA5JYLO5NUF+h6e39xRnMCMLalgjAYJLO3MYFc+WVCDXx2Mh83L
kxaNsdud6wWiuyS7X+VzZeKL8zv1V/F0JouoWyAtzYP+0mYSl7H/lNuLmYWln4Dd
AC9BqYFTG94eDeMHkXvjn5Kfrz4fx6Hi0+GhoG2iJLwyzsj09Y+v6gfzvQLsXUm4
6zerRAPU2cWMPCqnkA/CWFba85S56+ChohtVWM4aB1Sp8zhuZylFPLt/FdVObJbk
pkYSSxA5ysO56Wsr+2g2PGrLb5w3sVF59YU46MN39XcRAj+4fzo/BpSYoept950d
rRCNjeyv5DjGtPl5lWfRjCce4Hg0hi+xnNzpLlc4+uurIg9Hg1+rLY4JGNKKFttT
+KXBY/rPbROPYJiQA73wn78/KF48qtt7I78Eg2ac5j3ppBomh9Hs0AAWeQ8VMBOU
ay3wutBIMLzXeC9EelefZ1Re/olPE67B+N9TJtzs6Ir2uGBZibPi/FKfKdDn5tsP
nQWNXQ4vi3luBVoRBGwueCVurQHqpa4xnUZtJkVFTxb4XQb0REFC06CYkW7nIWS2
xSJU1taWRZv9SFeTsaY18UWs7UpbB+B2gtAxLN0jb/zRILybNdT6iRCiy7iGzWke
5wHax06qIeKBEQs1Vn3C7zH0Cozrq6pBXJIxSvfJ5zsf/8zEY8Kaf3KPVMTqgLVZ
epHxrJf5Y+uHkZaQgNMC/wuQ96WkLEJ/09oIhZu7VSsyS8+dlG1Bagw8cY7wz+m3
mLfuphADaOIyaZ2dVZ/LBQ==
`protect END_PROTECTED
