`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4/TX/GbgGdKtsCota+EKuVeDBzhEDteftB8Vr00wpow/It8g8a1C0ddmxWQfvMBx
wemNRAU5LeJKbY2ZSQWDBIAu33kAPMKTHo0oIcIsY7bkLh1R8gYKEp+JLfpTuSC5
FzXtPGL/Yrfs2e3PKi6JtiqcvMdBfKMqsFjfSWUzbmnx2Uu6IsEqMx6c6c2oStMa
GcYSd+dktsE8ecEsiB+MtN9cPMniVh4Asi92TQPBrzu1yyQsHQInc8/lSFRq8XFd
2P/AGnUJZrpqD/tvxUdzBiP80GeG6J4sTeaiRqCGUDsMZ/MZt7gVeXZDmhL+RsEM
XWPMx1SeFM9c4XFTzbixUMUvGvtGcNFh3yCDci5eDrfEI5cDYiFJA1LjvnB2PCRf
/w/bscVypw28lPm7IfQxHefGWmn+c5/ZrrBzGgE08/qE8t+Zf0rwk6sE4bIcsqog
nGVv2X0nC9EqWLaRHN+h94B0Un9jfBzzRHBMXE08nirmrfckGlUOX5CMpJpY+tih
Ax+pAHUdqglqqAjtFGE0sqYEGeZxi8KG3hH2hSXYFLwvst0v+NnmNLCLAOOChQY7
6Z5s75DV3daUV5IPvw3puPE1ml6HQx5qu5qyeJUEHLlFmj/OMIRBz/uqE1K9P4KJ
54bdoCmw6JeZ7cAyr95dgLppexG1AQu9Nvb/gJQhxPergZFwMCW90FI6ifZYJ3Nv
O/2LrMnspwq2UGU5qeBgGAMJj5U7OeX8I5aZZQ+MTaKmjNV3DYtGfjFmMSMhGWg8
7PmXbeWUBfPAaTkrhZVlhk/GzqPIYns0oFtY2WlXtWzGkNzQ7c22nO/9PQK2eNFD
wCAYFTOGrxDaCHztAV+vZxTD9YlChmsojXDzrCbPmUqrSvRndpLGFV8RFKbY/Fnx
WRAQbD+p/3aPFNkc2wryCH6HQXs3FvGPGCb5MHVUAegYYW4mgFoXbThgaehFwwp5
P6/RM95JfeodrNUbFj6XW6M0OJlBpDFuxVm2MBKfISbKdrcRduPWA5RoWg9DA86D
deyCb7Gzl2VgK3qwrw9LTgbsBg47L/jEYo38sjHEX2JOZiWWNTCHU37tU7kPanAL
D6vfnr0o7hKJSKwPF5eWZ7kxTO//VrsQzuJZYP4C+Re0RfcfDVF6DUIMcgPfaU1W
0xR5rVbneNQSB9wXn5Qyab5SAKnRfhy7GMZ7oPboO4F9LtP3YBGagY083DBpaqor
8RMiN/b33qq7DqiZZ5lIoeFX2emKS1gHByehP5CmwLlLyucF//ND7IQLA4RC2nWI
FirPm3aByzwG6c1F5h+PRJAfSnKLs2s6QxUgo8vcXE53O2xDU3Oeiy5uIhYBReto
lh/At8fExxL4m4wbb8j9X9fV+3KUm2wAmwg8UGrc2wN2GZQ5ZCHgLqMTjrzyY8P5
9jkmVb1IipvVNO7FWVvUGmGBrSPgmudRO4RVuNnf86T+BXV+eJMAPpa4ZyZBQtRK
/uBXu//PFJfpC226bn6V3tMy8ZBzfcRpJdBvJxwVreTG8fOq0Q2n3YSCkC4wG32a
C0TfCNnuTCq0D/l91uY+3/LF6fZO39Tg0uOf2Xyq8NfZxFDJIYwZQLU+19fXMzfA
K8XryMIaRrRGNpdWrMAkWgThz55F+6KaCyMnNgzasPq6xQL6CrQkYVcCHLoBZf25
PQi0BsaUBp9neVtCtUk8iBScKE2wu4QUQoKSNhcfjSvkGgKPou0zlGzKtZCy5J9u
ifAz9ptS8zFWmasJkDOAXx2lCBisTDX8U/d7L1ANGk+CVEsdwFIoAoHXvllc29Bi
RznbC/s6k66sdfGzrJdVJsCmYYWCnJV7QEQjeerJi+jjYW9g56JDIIx6n1TGdsVK
17gGdeXk73ew6doFYAc82JHK91YwgMeKb7g8sAsyXnmEZ6tcHXufit1OAPTUiUrS
dHEDfBXPCPjg7IUYdWQSSOrQvPVJhEgcPx5DkkgL7tJHzKiqY3tjM/1u1Bpsx1Q2
oT+mLpQ33MJJDcVBYCa/yn6VBeZvOCZU7w5ihQLXT3lGG3T+tIyRHXLR7793rDov
yqEKMSWux+uqaAg9GC73KjaPJbAMk2xj0lEmmSH7ykRjfMuKUhes7LLz2GAj4L7i
xakkR7VLBS+bPgiuZbunLMGN/Aki5/Vj03FdYhgKg2znmQU7935DqbGpw2tBBOa9
T1r4fNt6WTJNNbH01ZJ0qR/Ak+NB7WiTdUhRF5fiKaHwjEFHNFS2MSh55A5zrpWT
Q56QAhPdAd0mrc1rRVQkBGCGfziSJ49Y8QXuSbvysTuLRis9/eGJ4L1FyXHyJ24L
MwDOPi51rUkYaUqYQrUheInMBApSYBQ/WFGv1gw7qWH3hvP7n6yZKSdP1jG2xFUv
TxS0bDDU8ewIn67Qej1BdQ2YbWyAAItWtzRDQQLelinafd3FbUh3tEMu5tUYCMUN
07ZowGn7SW9mcu8jHUZIQEh8NLfUOrFahRLs8m8+HfpGeQDYTYTsMQsQ7yPs4w3K
jp3ErjX4qsVwdr6ooCmOjDr6hNLCSvS0DczxwMVkWDn3Hx/hkWLm5aAJ+rnjXaFP
2MTyumkS8xTxGImCva2puxcsZPwrGwsF8iRdhhM57XeGA7Ft9E+y40kASFGn1R19
si+DHkL/BOLc/ctKPn9WA/jzAcEaQvdfNzt9BEaay4qxandOp1OcpuOzkvXj6PHC
wW8NlJDSzPtwbLIcrCISe3lO9Lt07I6sjZ125X4kvNDbk18/XlEmwtzzCpqsvyMz
JwYev1DrrjhAz+/LsLR7sDf+pIjMYJGarxY5hep/E3uFxGRzVHCvW/6mwvn76JgK
caPLOWzuHzeNb2g2lQ1vSMCJMzdqhyvUWRpCNb1uThKESwqH6W7sUtnFRXJF4gtO
`protect END_PROTECTED
