`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mh8huMteo4bikLWJXX8oV5x/4Bb/U+f+4GGpPIphmV3w2ZsLxcA8E4gMHGluVzor
DCyO/JpVLYkUqwjz9MGdOS+op57VM2t1j5vJDLzzOkP8LeSNeEUEDOzwyxCyKCuB
pmnaLXDRmMg2Q+VnW+SzAngnNlY8LoLs4or2kCseRE+KZWKBmmT2dTJPlL6PhDCH
Gmy0b33MvtI5Va40WD94pR2vwsxQlyIdKWLe8NsWhp4XNepz4FnqBK5KEt2kOYLj
wjS+rifK2tHabq8bff9fIqDK12Ee6OD3luFNlJoaQjHqlApUjo4MN69KIIgzEOnz
osn0yFjKC3M1AyF5l0pY412YGhpemaxlk8pEhF7fP17awoH6uFx4deuE53j6BA6T
499VPi3PhXkiYB7pc2Id2oMDmRi/gnv4XL7yjPi1uth7Iedn6ZHoCSnfuqf2Xde1
MBAkGuaTvBNwoBHdB+ND0p72qR7Cy0+31s7XycUGDCTfVykdynHiHJnVOqTNKpZi
igyhiI01U0J5r6Oi6i+MflEyv3Xe6uMz0ZM3j/aUgZvqfZO3sdEinHnPPHjAR52V
2f2yxBU+6XmC2LIBR5iu5sR9fq7+HVgwERiyMoQsWR0906xnpmHNDsBVFCjQyLaZ
SYYMs0cU5QtxRWqdUkJFk64GWak7js+2nLfqwpVL+tFKKOqFQ1AjG9udkOu8g5Xj
jjjjnsBLWayQMUoHm5W/9goMdhOO+06FMptMOYABE1ANRzPQVQWsOQGiwsoyrmEk
PK7aBZMPhqyASrmEcJFAa4DDeOeH6DSI8xYbFxHxIikfXiS51I6+Zr0oX8rOEFQO
ablWnpA45RLVZrhEyWE7570cfMfgNOUMJUghYAjlrG9VsaW0I2O+kOusiLc0z5Eq
ac4jxN/j2B8l90qjM35cRpJNFMi28Gv/+LlOrKdOGuGsEribf5GRgqgh3yc4tHdS
S31dAT5N2OfI1ZogxdkGm6395wcE99oVTH9nEJ6DRKSv6+hU1PqD81ls8ITGuTE+
MGC5UpESseoNDdHNUonXUuYDFdYlI4wevByiy4cz1a/TnWDKhUXVTB096BHj/8B7
neO89XwdFNcsuTGE2WBjr1FOe6pstNjPLo5D1iXLMvNvCgQNT3xJtfU2wnMMEpiU
wq/W6QXoS+B00knGA9XjHoMo1zs7lBNAt6p7xT5lPJA1KTuNXzNi9cyfCHFTJ6jH
b4SmcI7gfBNrwuaEiX0nGAOBJrVvG7jQ0nCFBcDhMwSnjTt9+dUsd9Ca1ehvYelc
w4SdrAjkr3Z2EVni2Y//vAz2XPkBMSC2ySc63EW1QKF+I/pZyPqlApmXcYA1o5jd
EgkuLAJojJDkH7GUz9kWznFek+25rNvlJhNXHfYb/GFfatbPDgtryS6MUnZ+9tf8
kKEVqcgJcvZNxxnTs/flqemJaIdbNMIycQN2kM+jf+d5NC1qFvd1T62X89fxPX/e
bgvE5Jysod5VwcKF1nE31URf5YYgOBtQErPxftBxYUvUyoxecD8ThTPhDk3LGO8C
xI8Mi/A2d6VsGruGey4vQVDdrauVAvfxlBXxEf6HTv+fyY3i+qCJUl+8SszrueHi
nyaCX/PC6vRb6k7eQjIn3E6AAdO6NmCzL+bCJjAl0RkyZV9x+zuk41qUhgYgzD2U
WwTF9DiN7W0eJyerWdo2fM2yNBqiDi19OaReZrc4s3VicTPqw7V7RQ3cBN1+IVpm
ZFr1ngamR2NmaCWTslpMEl1tqog5lKPamegmb5xHsDXNMz3287ZUlCmTJW5wOrBi
rwrbwasCO1PUHiKhIie935vIEY9bHKbUbqJ7nbmhZuCRjRHplZmEl0pNLXB8BwPz
4ZrG0jIRbxO28mEnc6qHgbR9kOxblPtzr4CUUBJlik30ipVaVRH0hnzQvbHlWgEu
/fVnDhQ13N9+3Mz1Ae972h42q6IfIpLdkQHfRa4YjSCFn+bflORqTUuzocsojCi0
l1yta1kyF09FymLS8mFb0NxLFkN6uo0Ib2Pmip1dG4nRFoLeqTSXJpeQ+UoD+xZE
Hsk9T+bpTh0wOu0z9ODCV0sxcaE81sYb5SwrAPiNDa3IHTkmH6/OyNm0zjOaepEj
Vgw20Q67ydRfrSOWIFsNPrxGqI0VBLQp9tDvndWQ9Kg5TjcGJasHwxOAHyIvbtmN
fvyjx6kYv+ZKMUdcOirqfDjL/LH/f31BHDRT0ayonv6xwzo6IwMhEczhTvn21Ffx
2scydBBJ+g/Y0YuiIqIwwR2NFDsq+bEXMeTukXjja/B2CjXd2aRbC4DI64BTuXzo
KxJDcYo+JReh9J/yhH+3qzeCEYIPlaiwnO7Jv4CqTdTSYCkgIAPqiVZTScnn+ryJ
5oOfGFEEUODvYdj3+9KJkh4IMeAydTtt/kQhYeVVUB6ZFvFkalqtg8p4K+i62iIp
4AbNiSlGTiWZTTWV5RlZsG36RNp+NTaaWXD3PsijoKh9W4jMQ6I7C0I+PL+hJsco
pxAzR/D7T0OneR3HybK83J7RRgatul94uO0JLgnqB+ev4WxotDvVgxqfmwySWhvs
6OHEHVIAI3lVmlgBUPoytng08WHAZUJViAtJecI+SyiW01MRW3rsyf+E0De66uvZ
UZfesrtZcMwjc0q6mO/coY2LXW3DFzgwjKk6eUTGrGiVR81XooQBnUBKuMBJsLXo
P5iiojbnuVVNaYyaQngoQHHOa7PSlS4ZxahsqpgukGhIhrDLeZ+YWh8BuO2d/+6k
KDNiDQ6XUfuOg/CeKKZTqpoYZMh8wS9A+pEk2Jgdfxa9lcSJr5Sw1PwQozunrzrW
V7ekbHNaHX8CNGDjJO8WdXR3d7K9ipY82kZpFhta/l5vVFwGUVg+h7lKCVrL3NlE
Ruyfx3G2YsBkxwaOthgNG6jJk/usP3bRUQ3n7iFWZzk551xDV6FAebCOtSfVNgDm
J/3xlAlAdtP0KBNWZaY5DQSpSlSPFzwSK4rWbzJkwmURdxcHqXPREoY6HB8/X9lW
Ra02GaTI5Dd3tQmVUMFZNxtmeXY+4dOd9yRnxOjHP5jTfwUPTQeITOtVVLwvhyaU
5vDczaZZkfwnj7wgTgXy0ir0eDe+4KqRjjyS3BdQOS/a/QXDFLSj/+1UoL6THsxR
How50HHhZurgJvU1XMvhHCNiSgv+/3zM3Zauf4W1Kv5qoscy+Q/RjH8SKfTftDxT
h2/MQRNIZesos1HH5YZ7kvgyMobopXGJdxgPXDTwYqrb9ipZI0y1teqnwh2sf13R
cbNSYREUvxQEYejOIpNa1vpjtdNyTr44PYdHe5k6KehnjREUI67hEsZveGnlQdmw
Br1manXaq70WwZM1A0BFC2wsytTBbeqmehcDd5LxEPh3vSBKYfTZMUBtkyT66hei
vtd7z+WnX1pXj5ZfWuMvNxX6GWved34uVls9jgA+50EPSVHoVLX3JseTAwb4KDCR
tnhUVTQrdohaAcvZicsNz4Pe0JOwmDc2Y1tkynxpaoDJBFeKVwyUz1zJ8dpTTrdL
s8UnMw+G4MLkH5qJYcjJeO70n+uuq9YmAeqg2U3OlnYCJ/JxoKJ6LbS85BD7onp2
0OnP1yt6/JcV9U/dXXY8I80kyVRfIw1ClZbeUU/bc+i6oEwqJc8BWCXdSwSygzs3
RyFj7jAj38CisCfeklWee6qoNx0yn2LZltheiSJi++DiV3kJjGFw4XP2bmHqGlWE
xGBkra14++CFYKn2nCzEBItFTnSh3C0FEKOofsztIO3fQqOGVFAV44ufdMCaqaDP
jei7e/3Z3V3xO8F3H4Iz3o/NxX6iDNxIByM+ccCppSb5pLajnbXJyTz18/WV5u63
szyzEBS2HG9SuMtyonlmuhIghO0PHwDysQSFzyjzmZX7Kssmm5ZVJr9OatlVH2oL
ua5npuHpRyAE8GHYZwNvTA2hvnmxNl5T+U791BnR72nbg/QkH5Xv7N5bwbx7+wfg
20VQM0udnz9P7asc65F+GVtul/CpeJ4tx3G4uPTCNu+yF7S40lP6wU4uAz8jSfGG
x6ZKi4M3bReBVzzuis6X+i0xWHRvKUsfOaWvqvTkoMncH8hFi2AMjWE5iIiaZ/0H
+l0CWLb0Qmcp3Vp/1ALKXjON//LFMbbr2rZKDtTnAn4ayPodJekRvjkSxPku8ZJz
zkuC+fi2ANSxj0mHdj4KBd7yq985t/gnG5nBhMmHVFwhrU1CGH4pGP1c6jUObqqO
0Qmis6AxNnxDB0EfJWNBud/FBtmPQj7Vm43FJiYsZ90+ON12KmgJnvOIJuDN5fbR
DiD1jXL4h389FFLSr7G43MvU+Shh+qfEXzyv5jfeccAt6ysJ553CoKE9HO3wjFXB
rBs082fhJ+QC7nYx/G/ryqVO2x/Mpcw0j6FNSr/oYCjg1gT4FPKUbsbDucWMa5Cm
PpXut/yjwzjhp2P2YNiXTOLouCthIE0lwKanYC/dxf0IeFDq+gcaoLuqk/goI0rJ
EG+eNRgEEJPBTkOwtHiDJdcI8VhQazzPhb3Up0qCGACtzwZze6fQjj+49eKMnv/d
iT1reeDJOTHEQB3L9u3b2oSO/L/pGZRfsbYob4VGLMR8Dlb1RbWuQ4vFSi6QN7GK
7DRqzT4qPBaGpF/73Fl27+j3TyAv4YfJBxVy5Pfv1wezm+fO/gq3gCuXX8FEZ78+
4PV9z7v5QCD/dDzL2cB4Be3A6Se95LufJGewpjw8YvFXgn6BMRLTRvNaMfJNiXy3
5GR42dNKUgU51DfC9SjAHpgMVuh1ESZle+7HiUOgf4F68mA1I9R1CVYlQUAxjSc5
9q7+PZR3Y4ztIS8Ui1+fA+baDU0bM8320j7enWhAVG0YtcSDJvU0ooY17gN44wq5
hpZgN9RaJiTIk7k8S3BM5Nc3Ck5WKiSzRMZPQNVM6DkXfPWhGW4ThhUUHEUH0/UP
S47S9mLNq1DUiJFp02oyfA3F2v0vvRM59Xbju4Zi0OItS5GKXbhmLypDYVPQP9ZS
E16RSZPEj1UZN5V6mAKWKoJ9JNAfBpbWH0v/8orKuOoP25pSOyigXR+olOltXwlp
ns2+ZBJrwUSZfddIZyC6i9zFuPj51yZiC/a/Wz2+Tfbh/ggWQ3a4Unpd/5T3gekI
wbrUurNNvd/DYdGqYXnoqN9Z90Ncxf3T4B1Dt/TXb7ixTqKJwxqtZRM0rEDg3TxC
x6NyuEh3JVAcaFBiOyETVYdzS2QoOdVHSzNCGcnC/HeZ/q+SS6FG/A/4yybGB7me
42GNLgrCN7A5gfyTP//sMvE3kgfrYdqgTBW9xBeay2eJCTXx2sj2pKfNUI+vLvFN
jGgx1sMTa3IuU1h0dDZvk9FEZh3F7rfE48VayYhcUUWSDNghzeCttgmb3ZyDRl71
ICDyG9AGgPfyzZy5ZJvkUy7Vl8meY4vebSnN20gBaovXdSEUUtDhRV6q2ILImddE
nx8TlQvYxPaQW4gryBv8VC3VB1NLih2cj2pb5rS7v8tsBp0BlpNnbvoHQ2HCocsI
aAQoIGYIrB0ceFHJHZ81ncytKH52gEiPnZz4vqCzfQhiOZ1X9fqcygM28NpP7bP6
FBO1NOz+SM1cKs7H4dOVEYBIZGVR9P56U8WS1IsZqNC5NLZ2lOIVLoiLEmpymuGC
dt4h81LfRlf1O5fhxk6wcwzhR4a7Hr5mnv5p9OtXI8LFk/nxKHn7okitskeU+qu+
/rDbEw4FR7wlE8Q+iaFsYfaHQcYyX8SHRsyTwuTL4Issn1Isw0jx/7yPgp8nQHa3
lYW64gKBzqVuUxIpq0KDnZansIkX/V4GOq1EtdZfhLsU1EBJ4QWaBRCtf96fxOP2
EZfeHevpqt9p4Q3NVDZOqKk3l72S8+L3helZCMe7/mky/frL6xvGMJqSK3z0Uz/r
mUpSrtPAcVOZX0ShWeIL8Sz5RzN6Sqw0AbtE4Ht8+FFxrPUq+asGjRyQpZjddi9F
nTvXjbq7udJukVrb//XYmDdGwMl9WxU2CV+SfarRSMus7kPo75wEOs1HIAnJk+Ut
MEi3zsN0JM/emE+5sgpr37oUGMb9SWOZpHpbPlQvMp2jn47vdZ9OfW3Bo/c/ruFc
PmUXbK7mki8Z4OV75KJMeMEqOW69r3KvPFsUclnM0Gk799jL1FZQyoiKBEsOWH0v
rPWI4I37U/H1dsc43M9O55SVdoG+nzyDt1fEuafgsI1sVEOk2krLQRA0c5OnGAj9
HRRw/ofH1jAPyr5qyOJ1H5b0Z3jwTgx1qEjVfI87cP3DJ2VH8VWAZHWKSbK68avM
Pw6vkDj7m2e/luFTdwD4SIvflwOyz3HV9jlm6tObhSID2r/2SBZOx6E8dGJ37LsF
mKapdigauLmt26OFKAbDhjZ8ZvFILa3iiEvMmkHauoZYl/8za7rak9A22uzdZ54a
8jVqpitH8VTwTLVvjIgw+ryooeVeUw+w3nAMsr+Z9EEio017cS36BaNY5/2DyJ26
CXJiXF/BudxXYdw57vbrYNxaltD5ZU+yUXDzM6eD6JPiUpVXENR3MCoc2j/7m5uY
kSq+LgeXt3zSrCW0MqsA9Vee0siytvKN8IPeZBSAZviY54Gued01IGhIubD9rHkU
r5KAoY2MRGr5fhM2I89kKEbi/dZUNlos9NnKeVbdvVyLMLdb00/Vvbs2kWaRG90x
3kfmSj8LxrEev0lV6PUC4+XvcNKAwgfLa5drygLGp5IREAnZWWD90kQ69BwYMIA+
3eSiztdAJXSP9UIR3H7IfXM6Tc0ZKRGDa+4cFtbbi0K2AJyfLpkOeB1m7z5AwJMj
R48S+pCm8Ji2PmKuXRa4ejerI+FsYbwq7P7ske7Quttst3SMJnArLnpgUlyeHuXd
Hsi5+Md/nCdLH3QugJHjMuJgVMVibeTSzHOcdsxalFd2TaCy7E6m7NnbzGwPUYek
IYnMF1h8ew58Pe+A93LwJKKpqFMkkw3cLqhIvOX1L+dDxuSrcBNXWzVtbKPM5Rr9
igIAb+fnbRpGxFb1Cc4pjJXxivXKGQlyXnO40A1skgblsYYnMNpHxU8xmwsRmB4f
kIj/FRofxNTv6Ewtfprn4uQaf9pBetzGGFMDwO5g/IflhRB1DSjAU6NFnHegm+NZ
6Avs76Th2+ytUpDkfqULhvkOAm1aTbfoJWU9uZvfbe6Ruag2XEHUKJNbNjuu2g2H
n/Ti+0013/1h40mk0MoMCjK/3m/EB+rYcR1HLKJpS8rzOSYriSABIG9WO12ywqXg
Xxv7D6pcF7j3m1NPZpNimp7JRoXdzosehcvUC0kDfUa7ZQlV4J59Ov2tVdVODi+J
TCSqwOcADxfiwtOvIWQiz9E/wTdvc+Fz0x8H1DJx0G/zeQsJdzjaeT5oGQkqqZBK
+2ejVR1lIYAXk17QnMtHWz5ZDkw7/b9BNgoxxgifRCfemRSivWJSupbJ28RJG2YC
05F9jfI8DhMcfVjN7buzmHJRTEeXrhgaSrLC5pSBSnK6J+IdaUeq9B0+UKsV5ULb
FZ5/5iIUUw0beRd32UmoGHX9hoPbDm3l3rLI8zpD05mauVTyq2ww0sVDvWSaZ0vj
siRRi3V7om1oclEQ7ay7S9gVHaEZh6yg289q3nLQ2uQ3PFqtoMiDJpKKRqWsvXRM
tUtOeiRyPf8KWS0Ij0z4GST0EDOoBD6OF2HQApL5Syy6mRyjKiNFoLSR1F5oCHzD
dM12PYlF1CqEfL9fLEWuxW0+ZSvJwwixI1jDiMkRqr2bp6S+9L9KZhtkXUVWmM0H
jgqJzGruOPnMyCtaS4BY9WbVOIdyZE8TY9fHQOHlUTpCUZmPZgS/8bZsM27CWUP7
xDgLFYXKm96nGy1aF682/HVNCT15o/s4/1VFZq3bupKYD74ooaqvsqsdmjN+8cqm
fvstycvHkFOlZdUrG8DncJ/BK2/LfsBDZ06XmpufTJB2XqgqXAvJ3FR6jykp0IwR
k1IIVfxYA/wRSUooPbJBpacMkQLlQ0zGpb73ghMSHM2U45rrOYPpXP6Ehg6SLWAC
HEWI6TRCcsy+r0Xs6WGTk4sNrHKE3N1upiXL9WYtq7mBdXKGsCgnX4sqlbdaZS/u
thiV4l/uiolYO1nBs3HZ7l/vNuNYI0oL/fnCZoNvE4djnYfkbTHEuBamGGFFZ1zB
LHbXLOK2lYeNwUdMzid8Zgy2aIkfAhZe7wiWsYtfcJKDug3NW3qUHrmH2/bVEVou
xqDGRBa91X4mliL3ENY1hs5FjiJfBEdPGBojvB4DaTa6Fu4onk5t3LR6GYTd9HP7
GBa486RKE2HFB02bWe6VzmacsXi/9wqkuMwq26Pdjn+FTur5CnAyVe/VUtdmyDth
O69eHl2qPAETXZWHPd9gSRSM2v7EptKpl/rmUmCg9IS2Ra9/zAYMpCX/b1YK6BPo
Vj09GvZaOrdGvQa5bfzMHWwfmfHeEaBd2dhYCvNdHR1B4e6dLAgI82eJXcnn3YsD
QossM6X/Ve8aqwjRrrfDEJkCKf5X89E/fY0dmmy+tQzo8cZqdaPfXZXDfvmmwFU+
kxchCAXtIzqeRH+xFmFF34s71erTAwImD9GDI0933QGHcA/hJGVC8VHtDOEqEaPn
Sj5tYzhSB1mU2DigDg3wfJ5ONOrWTDLjfMtYhSNQJ5SrwR65/Xo9ieN7hnjXbE42
WPEX8LViy/PlKfvsoJdrrltoqrHKV0iLCeMuz2DuQbTIVNp2gvsZykc57kb2RSuZ
DRxe6zSlYGs+WPraSwmKAjhPHYHDmxiEc/EY6QjCXsBi7Dj15yFpX/tdJ4GHoIDV
32Obm91xkRPoYVUPEkLGHAi1TdB3NX/vnT9H18TYPnb+PJm0n1yn5vTfqnbznu8z
ZSoXAAtI0eHxqjvcqBSGZTEEZIBDR54UnOKbgAehFnDj5IfzmwKXUnjwL8QHdy/5
TFjEo8fZMwZ6omVqvt1qVbejL7/Hlwqa9y5Nyd52kU2Ll0kdUaA8/AMQJqNQ3AfG
zssBKrKYeERkvbb+GtOa1QgNeV1zgbPtTll+2nJhpdUQT8YU0yVSKgfN8X+4VgXR
UriQ1cqHB68OZmrcMbY4cHuYCW76R5GqX5GyP8Mq/+EoEw7HwlG68RA7bJuFiBFQ
o8zKh/JYGajkwyHAlLSXH/xXMQsB0MiWONLPBAOE+rP7oGgu8BNVjXIxsbWYIzJZ
UvWJAaKcuH9PI41FZcuNTjTVcRQx9u90jbuCjBqWJETQEGQmBGLo8P2Rvfxu4VKb
s8pGSQvvlnShB5/LYGJCReG94Js7VCX5r280oaiv7BhgrHNEc5oE91gIDxNnfs8l
rTJkvOGvduYD2wfhudE0zU0rOz2WKYyCyXVPeUMwTqp1mwFGOq063IQ89W+wFhPv
XTV+vObyxv75648LHCfaVepY/WBpEhUcJut3xbokt4Dpw8Hp8m02OC7OfSNDuQ7c
ttQ35ugoqCLRSrLy5uLmqFUg8EX0Hf0pBrzvBSZfUMkQOXEG6Razj0tEblrLh1sF
ePNGJYWzsGPBJlf6WxdbNOERqyiwuqYXCf1iCgtX8+vFM+ZuTAmVxKLJswHUr1eZ
BS5NizffTY3wUu1UaQrmpZRBXQa4BQEzVt9TPf4TusZTNEh5D2kI05SZlUlC7L9n
kfUGhnU3quCe5lbImFNNqT9jLytiBvH+vUD9bEJBtGqePsuqCJ7jtKnr+Q+GZD6L
iWkCYK8cvKhoKyS54kLDC74Q5VF1jh/T5cTR3WKi1jMPwWafjEmhOkG7TlYYaWac
CwKy5AaagCydPZzPYOHPYCAP78bQblJ7B3LSsfxcjHWUcAtCBC//YcttkFUYGwmw
CSlMF8gYIAJ9DgRk1+DrOk2xlfDhgfFB1bhxYdY+kd1JqrkU+LDwaRtm9tMCYtRy
0UaL2vg8EahwnDUo4Y+WE4rm+RcUshN2WHfVAPZcX8WFLj5n6JAYIy5zzKBOOfME
RBcHOOYESjOI3XgnhwiBV5BsKM4iPr9Y/ktOq/uC6nKqrMZROuglfvYvQaaH1R5q
ZsA5XibfmKX1eGkxZsATOojrT+4WU4I+YwqEVpx0vIcBGxE+GUqFiPdxcuGI8imZ
zhj1yhpCfMDNAa/E221pM+xAfYWHTnbDw3FNHKRZBfx6bBtHJH60r+4DPus5G9RI
DQ+YY7FANmBagX234aOnaP3ak/zn3dPStL11l7mR/R+Sag+ChvXleWLykJvswte0
3ZkpmHwDXex3UJfuBmq1NqFUNF1FBynQywntcGeHte2WXeYtSAJvxgPe9Ink/BHF
P/YsN5dfP59jbe1NllfEASLjHElhnW+9f7g5iqbZd7lRoZ8gfRj4e0QsUUEctmGP
V65Kt6fA8vi5ybF6AmjoGoPTIf4CkXUrvtnEpu8H2hslwkv3OftJZf2fHRpym8DZ
vx6WTHR+YiK2YfBZcK10lyQXNxRtny5CeKN3OFbYCFwaju4oEOPslgaXG/F9JZAr
/9XdJZmlOOL7xKHFM9rafFBFkbTnX5D7CLXXPzHrbz1jX+hgRbgMR9cxX2j3uP4c
KN6f++1uwoQJp7V3yAF3veYAvNrg9Nqsm09rkkAtGbLl3fWxKHHnSBLCN4VhEU4o
i432Q/zMDIb+OaZQpLeu2oiAL++xh+Jpc2sVt1rK5K0u5vtoYh6ckb9yg5kCkDse
m/hwrO40ghOmdgmG794Ogb1/RSyx5zi3+B5SyKfO9j2AyBl35+qY0t7ek3iV1w20
TNp+3+u9NJ0SWoDU46EFk3iacpll+eQbb3VxhSc9/RB6/0c11GBhdJjkkyEnCMtz
swilYMeT4gPL0jGk8QtKze1a5JLeJ92XshsBmHAWFaqeFAn3G1fNHMCSnJkhaeB3
HJ4ddDwTwObzV8QpGJt0niP7Uh8xE3XP/zajrXn6Ff5R5d5Re2Pf95r/RY4Wu5XO
Z+f/hcatOR5eQtZo0ckFhRLqri0jQrRLIJjQTsLkAGBkjOkpO71RXLvng7B7aNVW
npbgytAU+twmRW8l7FpOlx2/RMz5pGmXXvL4WIWeXcGm5aH+u4DhDwFXxTn7pezF
qvgH5bukCjuprAfNWSxSjZ3EktxBhwqAjRhbNjUbAsd6fGLJ8JNwunUoqlZ87hxb
PhkXjbJHnUbmR6j4ESwSbLkxznzAriDMC7/lv1QvCqo3PB7BNEvxh/7K+7AgMICs
PbK6c9YJp0Sgg1/fb4NTULjNB4jdEo1JeMLh0eSBtqQQLkc+0EX5WaLamLxuGd2h
Yt55Fa2iiKCznnKE8jkMHbMVgQKjkBS1cf4HWleV/E3HTWikIpXzZB/Z3d4iRQC7
e9M0Url8rrQZHe3v64IuAsd2LPT7Q0ro3mcLwtNLnN8wj3/s4VowkCW5JqrVeOps
b3j+J7e47CKFJNbYyDJD+13jiDbAMMAkKE878SU3cYvkbdXSm/xLWZmKbSVv0sk8
8+Pf4b0Iik7kihEF0y2fDaV5T+yp4U1L2oRUy2NCX2nW8+zM9hChSJuoGGCG1+Tn
e0vqLR1wv3mDUixhhp+vqt/VW1/d9N1AnUkHPIOTWgKWdfZqTZ4B5d/R8rBKMbcy
vZzZtwTKB1n1WjEw53/pTmj5kWdL5KyVZGuj4Pj1fioP06rfb2jDlkbKaxymQ6HX
snFZYeD1ndXVmyGL9AOG1hrsh+E2s0PttCuaih9r4oJ/lqVJJrint2xdml6ODAKZ
ccaAteTDQVMM9RheUCaW9Ywzu6qKNXExFWVnQ3wELs8V5uWzHhNMVU8BdfNZZZGP
w9BIpjakKDk41m4efdycRFN7qEvLeuKp4d71FPRVoSuLEGd6VyPzWiDUQHRCe/Rz
G1WjZONpdpCLc1EJ07dovRk6ep8LPNCmfsD70qrqs8N/IYB7+lECMJkxuevhCft5
O7T/CFRo/wqTKi9O4jjJUK99eJJj730KDukkkoCDoyHAI1djpyAy6AykhAOoimDa
xDM0oR3S8fOmOJ/JbK3xQ0efLPk5bMsJAJbQTzWk0goQe9ndpS0JHEvRrGciWBPO
GmzUBunZS7NxXpSdxyQiUJ3J4dlp2G0nailEbaP4GWoIwkNUhk3ZVsBfhAnh2LkH
5VJw74PJamp7edBJE5LQqfpjXhnasAYiVlFMKQyNJl/6+CVTO7JIETF9KmOqRiVa
nHytPHy+UOuJ/1IuhsBxRrP4i/OK4csAjNrhEMJvgQmwHuD59xdVl2Ysgsc8UGky
hYzz8pl3ONZKTdh0Qc9itQxhEpPUyGcGxbOcy3QxPS+4t+iq7dAK78p1AnlgDZpt
tBA+E3zQW4HUf/01Z4jrulbxJtJJClixiC1/gO5dUfBw/xHhnsRWSOV/mJa6ZVoI
Qus3ylZAqYal/8pseikbHMk5LSh39DzHUntduvv5PtaYo8pz5aIW7DwrLoWaNRGC
EWzfoRKKh0+Ye7M1NFx6rVZXq4xgeL6X7hUHVkA9g1bODu33YNzIStZeTqveteg/
B4XPANw2C7gv0KzuUd7FxWRFypO2DAdG6f1Z/Sk7ZwaS184WWe20HvxqaYU/ROLQ
LPUtYeAmsdotpguoa01XLJ8byr/oX8YoOYpgnPj/9lmHtPLFko/DMGJ4lDlPEBJA
rhvBML1ayNkGNSGJQ0MjmNDzeJuc9U1HQqRD0X5bZ/EnG+OxrnTbkLRpO0YwugBv
5n/KLZnBFLcasKk8O7H32DqGqLa3Y/Oj4MnNlJWu+oJQU2SyP+SaHq+NKHu2o5DG
fmECKUndSgZhhpoXnFs9Syx2HmO3A9lxRmItVdm4blKH9yeTxuTcPNyxkLpj9RjB
/QDxb10JnobJzVhhU1vmklWy1MDlsJBSTaMbafuaxZFvwFN2WW0vNvhmN6HLARTD
zNQhuIs9EqfLcGRe6F/B+VuYFqKcH4VZzQPVOVTTXWNJtQPSKn5GbM+kWcY6QNDa
2v74WGPQUoAzUoXvpy8t2PFQmOhimX8RfaSqLG2/M9FdOMKg3Gx1lEIFQ92IFAvZ
k6YtivJHiCQDcTocwv7g7bkbjl+mTgQVOQw7aRZDEgz5N9GuQdnefcDSror1qGux
DB8/E08TVAKO6awhQ0xMPCthZVJWu150se09xf6njKr+mOAEXowJ1wGRvGibcnZC
E+rEub4cWIiaeod7CbCaj9yucY4UTLhT5OnlClnfH/CTLtEoBS6HMKATgwrAWIz/
JrA05nX/m9SqN3xPYatLyCsFQnjsN7O56VR1xn4XcbQgpF9G7J+GVJPd2eA1kHFe
bOLQARyfqVFqQQbA3gwFxE1tatz3I3frwVTFs/nTZo98x1F8rl2Sq8eoEqpzIF+t
c6wNfvpxeYwtH+mlZNs+WdjgOtAR0VU/1znUcLpJ1nYE2sX3Qc3GTEQ/xJpHRqkn
cg7WOJunDo+E7FC8Yth8UP6XRpzGGykCaK2ZMTE2s6JY8wB9M/IrJZjQjTjp1mtw
Gw43Fs0LthElRlSIL7M80KcrVYdwPK35Oues8pAvcDI2SC+dVN2CkpbZgYcpKmxU
3+EROuMjuG103EcFpxrjJqdEekTD6h5+1Bjza+5ZLOVGC0kkvmnoXE2ntUgC8zQh
OhIlj5ebswLVRJapVkKcovt+lra8ywlkWWd6EJ9m04gO2RawIE0qi/PU2ESD1tRt
6aX45+aX3ItwXe1MpYPizz35VD6lBVjjSFL2GQGyB9RMwCXwD6Ds/Af4626U1iOT
/H9N9Tqqva5OCSodTfQSkU2ZmkkdVHL4EgFV9Se74KX+8OiFhgXqLA/O1c3bpPAD
85U57CDktyaPquwNYe5v2huUIVn0xEy7jIYjkNzryE15p3xYb+jDVOeHscwP2DvC
f6dCJycxWJg2XLKtO8fvxUZ0S2GTIsN6wnWxp9CB5bvUnPc3DUsPGEN5yRlFpeCP
xw6NH7rJ5TfWUK1ATvIEOOOJ3Wtgrd8Llx932ZDK4Erwd0UUJNJ3BWX0E3F88pqK
Rxd50rOCSBJ/DADfxVs0zcrcnnoB5n7iztghrBM1u8Fxe7c814fcsOlcaIJ8TvCO
7NoaYza23RHb3BXVNzll1aeRg6Y+hsra9VDVzkyzTVG8J9ilBtNbb+4EAKeyQ28W
w16htixry6x0SsTtTJdsSiEvSgR85AL/SbbSm2LR5DrQHT+dPLpYdn0FRTrAcaHO
7kOOcp31qQUYUlxM3w2GKty3mkRWx+w7t8HsdiXuwLZyxxPxkVCXWBmdlPB81ZE5
tqfR7fM0EUp3fiYFNPvjaDb6HaRAfiL3KlD1NP4CaE9D9WACPtYAf4t0anM+FSM1
LepnbWVxOupmROEqxNDhsBPQFzQLR3GYJZmrcQzubniIue/iegMWpcHrZYo1uICz
aOcmEi+fg0XHHjBZyLMM8dejRi5NEJmvLT7r7giCSYQuhb9GMH30/J1QJSXUz5cj
thAstm8Q1sHhJkZMaUCDM2CBUiHpUwSjkNNJy9S3qIHHjxvF3a7rcXM3sYtDp957
UXT5VTH0iUWgbKG5nq/Y5q50xazjqFlRwzvMioIDOEYIknIBt6gTgx5k4OyPwnFO
IocCIMkPrxQBkEHIy76cbIDnvg18zddZwGL9ACOg/78zefjlTwL8IZ6C/s/FWBWR
v+eKclAWGo36b6085qivsyCegbATE5MuqIkqoVEz9Vgalp3Bf+rq4MqSXNopAKm3
6DMxvB65l6ubjD4NN+n7DrUri+drctx3AkNJEhshQpW5RWlHUrziIc6EMhEGYoHa
7HXRZmEnwyTuX/S44QxmjJdIxxzStWsHc3wMD8FTeKZcELtAWTkj9RS6c0/NdiiC
xr8/JcSk3V4WOF85ZUFFBwct6pSG7XtyLgCSUUgX3UX5L8tUPps1EZMe/eZQI+Ag
RvQhTRdrsVTDyTH38G7Wb3GLLI9bChChb+WLC+Gy8p8Xr93QMOVE/594+LbWkKLi
6aK90qxR2zwiZWjVhWgPPB3uzYUGYbpP/CpZn0VR1MTwyfYu4mJGpOBFxALFVMYP
PRkcuZv+kco4q8Q7d5uOed60w5NVQ2kifle2BjVthuO1HAchXoSutw/Tcpl847xe
rbblCsel8w0RtpILRmEyPM7FYPOjZe3RSiPQx4fHh7mthOKkKsQw4d6kbpeuZUZQ
60GJzL8XLaq6BDKRjEK6CywM0+nCemr0kJA9MwUq9l+qr19YARAg/PIlP/eQSSLE
5ihK1c5XGVQxrSJPEBWChhqTaXwebj11EWk2xsMhxMbV/w6OLD+GSYBce0vz2Sa3
Zf0Q5GqgGszkQQvBhbDgIkrQtBXOcU4m6xHRNcZEzWmT0pwTUp+URqM0tY7gacnP
fd1Be4IWJJZ6sQdh4/cyRrcR4wF2GnsYRvtHdve9SKTp1YOQvZi07GMg3tTRP34/
xi5ge/nK6biS7bts2LzzzJ7pot1kbKEOKHQo7bTYAqMPfGNQn5BAZIybQ5INLz6w
a6tZH/NG/6GqhmzRmajDv7pYwy1/ceFDEkHbTGyknH44B+m+/WsrB9oopTJC5mI3
SmtOnZETS335+nWKRJHk8a8SAtV1JMC+cPnEqIzTWQDQBl2QuhvfT+k9oVUcW4gK
13TOPevkru76OD89JA35Czfdg81mq5PvFP7HXEqSw4zEZKjly0EVyAVA6qQLNcvn
5dIPJiuyepdSiMqagApYtJHJMYnLguP6kSNB/ShpxS3B60ICNybzmqNGQCRvMcty
v0mQ9zAj7v50aPZRxlocGop7+fRlW/B/B1SaaQorJfVz9RML8ceAvcibiDk6mhxb
KrFAj5bVSdjiJhK4UfRTX3YSJTmIgyhHZzJg4M1WPCK0ap7jssiPRZWvl/lsVfOa
1GYKQTw4xT6jKH5bkHEHWR9taeUZZhxf9CFXjMTL6MFOt5xGOSYIww1UOu9Xyx/I
0bOyRy7KdQY3/n5x+RiDFU9rJZnO8+Ayx3MyWi4x7cCMw/4QldZoPF7tfmJ0yMYu
QtTm3EadFWKTO50tLHTazWP9QSLxydTRrrLarwSSn/or1eoBwb5ILIKNdbwTwX7F
6TVmgXxvtVfyWbINW2dNHDshE9stTfmZqFe11PWDIOwYnFwi+NbkTNmJFNzk4UNS
dRa+mQhIGe9X0E2K2tIx3C7MD2bYUMV+xjr6NriO9yIFSQbGwrB7jdPiafWJbemr
nKwnOlgPFWTHFuAYso93OONztPHYGcDfn5GLQ0IUTt3wP9ictCd6EgTVCfgYJYUb
Jt9PQbVKRoLmAoP9yOFUNRFc3RN8yBcR6jMA1Y/C+foXFBjuyVErhEC6BfapVn7b
pfJv1o8AUiCe2+5e/ROFNs1XX7hv7qAPMMs3bEqoM/pZ6JqZasXZ+EGV20jJHvw4
L/DGSJLijQx2+u/yPDeLMa9ppG4CwfETb+f4nAj1OZgnvg+6cf5pVOfvDgXs5F+N
UW/Q3RfHSfiq6wfSRn2oXrfD+2W0JQ6GdA52lQU7V+FtFLxfxVZvTNjVNVIvHyir
fKR/ycWOVipfvx0c1ySSIeGV17/1DZG7N4xP8LhHnW1I60v5YXYJOg80Z3aVGT59
4pECY4wpkoI/qsPOlEaf2sPeszUcML4G5DG6NBGaQ6BVDT2b8Nc/gJTyDMYGgK94
a9RPsb/XEbXfkLqjDKcbJSmm+Y2MdFS+zSJlPU6oK9n5la7hWN6nWtWn7mShQvNd
yvNuOnqEhSIf7UpSvkjolC3W4jPLij5yQe19cpj8Hw56aR0Ct8Vl8mPMmyNSiFwY
5nF88e8+As1hBkpkxHAfscNvMohdAVvEqeSVYIqzKRuQrJeEgO/4F42BfOgLq8bi
osgzLIGa99BPpIUcpDjvat7Im8wEcjUl3Ua56c2Gt1jShICsxueu+3TktqcJejcL
FjiuC0BAwq4jPrq42VQNyg3Su/pts4h9o4q+UR10iuQ8zBqT5z8n+q2wmmeBqjeH
pCVhZN+tjW2pFgr1oEHsI9UOPzPR1kA38PAFnJsg5KaRuRi0LG2QFzu+iMQhvPKa
WcquESTybBh2XfKCkPeAHcKABbjJ42r8utyc8SLFeI/LZVMebyr7qBaq2S5bmkFN
OvN479LN9qMpybkg398szol8H1JjQz675KmVXnzOrkww24If3orTNNPzTxLqk7T+
kyLxP3fmudAxlWVG0bWS6ut0Qur0lpw4sYyO/rzk25/FFAZFXq3ip4HU9W9OAIrQ
gNM7J1mM5KrSUSGz8aDDX02FcA4+NPxkXUgmpocgNlSGZvtP8TYyM1P9wwthSE1H
Hk9b363Mp8WRtstB726R4Yni7GIkevEqEhhH96GTQrKg6TUy3j+ZQhQtYEB+iATo
mpRHLtqW7x7xqPXcDy2KhdKaDw6MbsEgp56VQoRKuEcTAscUIsGHQR5D90LqDC43
VVXW1kAIlHd6M+ptGM2uolGp4SgMdpFyS022OaXN8cHeWfa5zAaldEpYdgMm+5Tt
Sa65nonWINMIw+ZEkwDviN7VfbA1Z9Jf0Xrc7HHI/INMukijratYoKQoXB97+9wF
irSwPqfpa6IW2gIRtqWRf/sG74zIbj6713XviGL9kS6O7IX0f95DDMke5Hr5nwtr
zD2AtQOldLINoulniLOFtGe5S1GE9feT8U4Zj8bp2GNrVLpESoEEpnwzadD76qDs
r43XVdsiZB4bl7SUqND+dmOvRhDQHhZ7tIj1/+NOpUBErWzo2b4cKe0k4gxOXGEh
IMDWjVX/uTrJavreZYZ7OcPGN5fRYlfpA8XJobCVvuwidz70kghuIwVS8R1zX8MG
sYOeobB81qqqQnbDo8DrgdlDVda9PrZIcMuFPlmNkxEvzQzXleyZy4+u1GCPJGWh
UoZRHVJJUEWrkgjFoVCvMJOwAxI/8BOg4GmLrjDm0QfOwNGh632uMGvG92YO3AXV
5ksdQp4OsAJtchPpCasvPO/7mXJ2h7PMpyUhm5GMLdcy8Kq+++O+PAMF7C8SxIz5
+NfwYQXybksx1qZCqiaOOiFqYJiFLUdiNYmuuEjccrDsCOCtF8jfcXHJhkBypSOW
nhj09yI9DwBElEbD1J5Hs2KJIcfRqzeI68ivGkXpw0E36M2Vorhuo8W9kRAnWOmb
j5t2yHeURXSMonSxLpOLYM+41gEN/uQQJXyrdM/7H+ALp7BT/typdOcf4lTHEtIv
ejucEGqPTDzbtKVI2bLmNFnqXYzw7lwDDkUukcJbEYS5kIfINQFONf8rJxOYUV9d
pUpgLY8NyHUQcvPqEe/pJSdNPgXI1Y2gq8oSXBq+o3PRRBxylM8ht6VNdwPIAFFN
ACE6dRG81YXiU9piXuiji4gGN3MJ+78UiFdLWnTgr+ZzTg09yHIuhSg9KqvSyJXP
3XlWW5MHoXSw4hchs4+pjJ5VRHZ8lUQUhhVrAUdsGE5H3SdpbYnxzfiZuF3r+xQY
asNUpt+5+5dSeJqiDCRmc+Qh0kUdArIqUgxHKivc3VZ/fj5R6REulnLS/jJ8kxA4
pT9/lj5OiSRK/p18wZb0Mebw+PNzKr18NLdHzny0JINrsE2qu28cUbms2qrC0wQf
RVhb9Xkq6aiwqcY0m/enVULzieEgYNGajez+yDJ1EpdoWQw5u9SocqNzwWNbIhbv
sioAjMgJV5LxNMkWYjek2MLwys00JdZt0OSB+LimXhDGUMIThK/PRZtFki2aLs/x
kT5hk5IhV7Hyv+2pWllCmbW2M1ryEYSPrJiVGRvdX331IkH+J9ag346HbXUS1m5a
0u6JiIJl++zEKLgtlxIXlIA4O84QRv55nDTZlRZYArh788gcKxCBYzo18ehA8efv
vD4affSbec0vvzciloAhePFvcka8z80YMd0OaPyz/cGgBfksutpMU/PGheA0V2aO
zH0SHo4lIU4Ca/4SlGcIOg5FGacqsYQr0fopEpXmIWXcUlBkSSuM2etcL3JOqHPx
cQ83bLEC1ksIUnHH8MoWSJDemLD+uZ/epTLvyxk1isPBy6PJOBT95CFyjMimMeQ2
06CJAvHsWfWu/AShbrAQAxUj2KzOfm6ezZ4vy5j/JTXZkA7w3E5fwnCC+txuSj8c
8Rqp6RLWImmtvUxTm0n8AQennRFlUPX5gv0+kBoypNqxvCyG6xf+Cc6zhVuHImvJ
5tHsebrFj2dp5HgPsk8wGzImvaK01d8E8KTkKHfZ6H/N1aagBhgJ+2AxuZ7hcvuf
IU/U4NfmEleN2f6GyTbCt7/I9SD4yijty5cC9f0uiZiySXqKpp3haUfeiiyqEold
DC4U5cCKBbWctFbjsDs617O5E5s38c7vOgIZeSxFF1mMY8ugh6K/xydVwkKUqvho
ISa4WYCd7FZdRJce8KU8MdELTVV7VeJeW9PjX9hbPx2JWGJjNwLQtTYBPtPpXiuu
irmvicJy6ikcHXuLd2Sc09RE3ri0M+yjqOEnMuMsU8UhvbnF0e+396RW9Pq+OJSN
vpCqJ0tistCiYNscVygIrLgIr6r0X76s2Ldzh/H7YiVzOtyxeeTAklsC8zo3PKoC
hUKzre3FGJPUb2MvhTxoNuYsFfHD8Wrh8Pd2eUI/TBVysLEeio7AbAnprbL8n/lB
qA8PsWIbP9VJiBhkcH4rZPR1VEo1uTvMgMkQq2Fv3M+qI0M7RTLz15dsmCoKseQw
zRDKGLhg2HcR7eWMgbL+HnX1JXeEF8gqrOjWU6BQvWPpwnTDbk9zxXBNT14C+SqU
KcIv0KspEL2CxwgASLbITet3baiZawBh5WseofY2nWNpILPStQNZ5MSXAXHR8+GX
Slttg+3gRGyD1rLFX4P/VksuyxS3pYFxEuy0HFBuL3Pk1JC26YP7Yq7jqkXizTi9
gWj/R0WQv0MSvipEeRXJ5NJbOuXURe17Lbch0FxnjW8W03gjvKaeo/OIkpY3FkBU
g6ptzTuYpylWRTbr/w7jPW+OUZTQYgJw7fpCfcyInyDsUilUPBd6G57YZid+D9wi
3UEyn76VHMQn59Eiop3CSbj7aVctTnptn2YJR8l7cbg1c5gEY74ztimm3K/5I6vW
S02tJH5dvoMOoSn7z6WFb8lNfWMjk/WVDYdeBBVlnFXkSt7llHZ60FlERN5gnqMD
Zi9OoHiiWUpiU/+DpecSxuVzcNy6pglzWLEZ0sSTFNAB+oEXnkHX2KnbEVpsACHO
3bucCjUS3+C/kTC2CUdYfHVY9T25uCJ9kCfnJd5fHnOZSEu8XMWRpBYFQpxBuNx7
PQwa8vWnHdf5yaFhIu48J4q3++BNc7j5OgcBQ3BBEjGZiuROP5GpfdLDCTgaHCHb
yrrH82i9lwfXdJs0V930EAJNOrbQz5FkEQFtPQOGSm87OKch9JmmIssTd9zxL/w2
fg4lXV/23wrnkWbMMZ4ZjaF460yTuN4OzPmst79kw6wKcjr2qGJEwpVxJaEvC/nS
LmHkmU3JYGh/NI9udG9/qA6bLznb5VzVF8v+H1mBrZrVGZSSlLwvRZZztpZ5oUbQ
fpzAYmYWTi3VPkv/H4B8xLe576IQddR7xRuUD/F7Y8lAauW4lFlecf80wi9zTw1o
5WUfizkacNfBPPIkLCBoViOrrX1d3IbgNnrKrhvP2Ds3ISyPehXsU3kRzc9pwtyf
eWMsUzuJ9pMvUWHl0S7nzGE+dIqRYK3MWuz7HmM0IsT8FT8rMACMxz4qD3riGjfd
c6tDk5evhHvY5aCaUuN8sPBh0yXO3o2ZUkoEyxGvgy2Jw3jWFgXoSWVM1ImXceI5
j/61FG/WEox8j4a9y+p69f61RHm6DCGc0LCl//b68lgCbmLHsgO06dJuTgJDLZoP
nLQecjwzln/n4yCnnkYtBUdBx2qmWS2QXvXL+JpYh2zFBOy2kgsQccOPHlfsRYW2
i2MYz/y9dNe5LvglIWDkFqzSjtmqd+NWWEftMwsdWZA2YArXU8Alb65JPxnvkY/a
9etM6IMJVTQBIp6daG4Jbp+8FeLsLyAKPbPYBIyj/sQv9zXWg97HUw8PXpJl0sm2
pOrSMQ+dII2n+fO321quL2kdH3YrxYrZI3nUeJHblQcutJw1qSHEqdIIxK0Qew6n
4Ma46Epp5JsCSbKdTwrDZu/U8u4EGa7EA30SB91tG7DYsYEQXNxu5wGU6wlOaGWK
IHy2bOFwCnzCDHJ0ON1wrfwG/nUS95ZsDdYa1MWV5QUSisvZWfTbyOsfi6t6KzaV
0HAQ+GOqx23oN14nV/nR2se7GvEp5HbB/RTctqkMBL35Qi8JT30r34Cye3wIjJX1
NDBxqQbpD72IVSgtWtce03FuICihCN211wgqoiO6XbkJMgC9awx+MlyFjgYyDILQ
k1i5tBtiKecgCWILKhchDJIjJ0cC5o4VKaFmcJltrp0rummn6htv/GIMDCzOpFJU
zTsfakluC9CEah14yAD5h507ml8jXyQ/W1hZ1H7mtggYYPe+EyUKu/viSsgJegmL
tHIBBrb3agZmk1PKfeYr7iVry/yq2tBAQACjwerZ1QAO4Uv9yiTLMJGYgCEJikCL
BYllSLLlqoQAjVgI8vlbS7G3YHXNhBtGu7uV9Nl0qlha/ISz3CbDTi3Saq1bAj7G
+27TkVmdXDWGHRtqqlvrSgDxyMYRB2i7A1Demo7n3GqSkSbBHTP9lJPhmeIHhhjm
By4u1HG746HJ8W1KLBEZpxdFpoVzcPRA1YIeEmLEwoyJXs33vEpnHUqlULJA8NVB
qXHq7MB8zemr2x7iCU96HNF/KVLKZr7qm7D8LJVyUVrngPtopsffcLw7gFHV1MAA
GvPcDfN7nZebEcB5cvZmC6Tq7hbBJg9wErjBIWQMZKGAaD4IOuoEZJ0K7iF297G5
WN3WmvizesZmXS8FaoRrwMkiW9P+P2v6r5kilHYpI3HdDJb40c6awZA0qANYfT40
bTmDb1Og98lkkcLriIBROPBW9ZgywDQ63pceOGhOBOL0AbCtc7BRgeEKzQPwcI6a
3EGOQ0jKRDpAzrobS334OQ0DFqcyOm9G5yJXeVgS8okB2a8DA02fHBMSWcZ1cTej
HfLOvWeC5Dsvt48qrTMFGtU+jacQI6m7RGjle4FReuWduEv66cOB77ZXsAJ7pSXE
1SLFVnNU7ib1tkQ5q4y03eIejoDlQXssPtJxJy5As/dvFXTPSPMI0Z0uKUp+ecLC
OGGjI0T4pfPvTA/fFkRvLKGi8Bz9+liPmm+MMl1EcmFyd5xDPCi67PWezTNgB494
smdnUa3MGqfF/RK8FHIaKkaWFxRJ254D9ZdR5V1Xgx2Nlx5GLOhiy7eWvyM7b0BM
CNspFMHtHqQ3XNd1YJFA1P8biNqqGLtPO6wTmvznpC7S8S5csYMiYf5EB8a39pT9
etZu2USEFGnGqo1KcwA8stLH1a640zUXwW1YqVZqfPPufLmj35OETF5OHkYATlqr
OmbYOBwlA0gHkp52UXHCfXURnpMm3XFBW18LoZ7Qg6Z9hBzOkoGH3nxpniYGttfX
ujZuTx9K7/tSOA0O17JxCvbzJ+A98F4n1Q7gQFWAhwJ2kJVNxL/ApOFP597q5iRl
xNQKUIrAq8D0jK1M1mNfQtWdlgKMaDfos4jeJLu1gYvyAf4MW0PH6RgE3t4tTbyP
cf4VpNLpZmGPxvi9v5PUDZbrOSYzisV9dki6ACN/MpBj/KD+/Ws3IqUyYxUvU0yv
K4pKAU5zBb9xMtw9c8CtybKVKPkOqPMHkPDHQgSdJiwt1ZpyDGLLZaxkYU8t8BeJ
evWzA1G7X14OOfKrwdfhExP3e/cv8P4Y1ZS0ysVNke+52Bg8PEop4JYlnrhDg97p
tsnFgn2nx+FO4bUcA5kqhd0lUYdStCA7os+06OOkTrr/kcILVshc0u0eOOn2uzwo
TVT2lxFG53A1sTDDgUuEuggxYHDP1bLZa2SlTnqmdb11ZQ63NXeMtQOrmIE72F1u
Bz6am50l8+o01wADzmXFtoT22tdgF9dP5S/gbr9kbNim2wBh06XIy46D9tq6cegs
6vPsGGroeLyl98NLMjOHHFD+ZFaGZ638Nx5otjkJzPN2+UmwsC6XYg0hh+ZB4w1q
uRBP+PS4sf8b1ZLqWsaQSoG1EMYEa0jPnThcIdDP1xQP1o8sPdQoBz0H58ISLix5
SNCAkCpJf4iR1oPWMaIqdT3ria671Y9wSZzWrxii4p+RsrWWNxnWZfPNKi+s9+yS
BcLiZmGdPToIMnQ8RN8xB5GEiyTXROao4z1BQyBcE+uf48wlPp0tYH53unyEL/sF
Hw4lgsRTp5mAz0OLpFNvhs7cq+o/Q75nnOVZWFF6hJNG6U9rnq+jIIHhwNgDPSR8
yjZ17oN5nqUkx4rtZNeKmsw8qPWTwcr2iqaDcVZYQa1G7bDzieWD9P5rTVH/N/Mq
zaWu55wRfOqU05ij4IKfu/ichlhpfIWv/Qq3BURB0Hv+tZ27qSwZIgf2rONLU/xw
Du6HKTc1VYTTsj/Qe/fMpGzuIVsh6DGxPO/DZtTomt1r6zCzxbt644RVzhUZZdbL
HiLlhxbIcZ/Bcg9S4FZ0l+JABZVSSTWuy+wj+6X2fXsU9IHvZeG1b0vnxnn9qDgr
9sqse73D7n/qsCRc/ezUkgRhDYVXB0gYXhI9o+d3fiYyNQhS2iLxopiFIQDS0WHj
ZuwyTUTUtOGi9+ArrvNxFnRVeao4GtvL6RtsGta0kXSo434W2quVaPKMcP/60whL
4vy4CuAdxDXClugsZYU1WBULQ5MGThmqx6yD/6Egu7P+xnmq1+QFNmsJEXhLhHne
Vr5bDbSGRbbq64lAMly2qY/pILKQAMbhBI23RlACg8vndYY4hRDaaUJVxeHBXbpN
/jvKYXmGHCTd8kxqD01z2nWrRamkJ+EFXr5P9zKgE1Bpr9m4mwoPpwo7M+L+6GC/
lcv+56Qts39WGnwL16oC4btcmz2HYVBxS3AfzVUPmJlpXPw9fZQLwRxBbJteJF0y
lrKtcKaHvM2SJt7rzh2LsSCe6k4/PvWJ/Tt75IzYI2UJPsDoK5hEeXoLGvQbqafm
BaYD+rvm11HVKu8F5HXIxLfPfOOsh6vjHCsv4SeNLQOAtrlZZuntIMZxAVlevOIL
SNw28fo2ICYj9WS1cUcgiOmWWlYiYQ2z9ChOON/EIjqR4Bkjn4yRdFk52wN8h8gD
CQ+xj8NXHcwHvs8Y87pcPfNMnV7l/CttVgq4d2duxF+tnzdHT6uxcg0nsKreIL04
3NTdMqtr7FyTPBIlivKtC1lun1Trfgyt63NMe3veyrEJLCyWfLuDQOhWCba6nqfZ
27iUtOpJAnAwobPbnKFl0NArihmM6NvYaFfNxl5lCvXnOsjnC9sMAWEc8T51H0qK
XknOsLYWwS/fup+Js79G6CW1bH1Wx2u6WezK62qG9AqQRM7MVxvjNKx0bQp4clVN
aN/D1ffHAYsL5dVBbm3kwngT3Hh65DVPAyRv7qYeezo+DX/H47iVr9+i2j2wpS8W
6bfmK06zDNmrSJdJSt2Lb5BnT0tHDJiRBl6Jg1iCB9yolYcO+X1AyKKwyuDjrKRF
iAzZN+oB4wKrY+mHiGHkn8cP6n0FKqes9AAWmwi8eQ009WYAbY3CMgrHNiK1TkZx
/CxUSFGMCPSHCSr1rLqV8oW75lhGzfLvEzYEWFZVUTVmLpI2QERFftvIAMd4WIrA
/3vOnFpf1kqsaLcOkWHgBRsUdw/1Luu6ji9ET8ZxGM6RduKNNC513QJ/04ZFDZqv
eB3FoiaQWAg+b9Sko8hgXMnRC3V0qm63pcKh65NTb7XdHTk/AmBrGNqHNAHX4/1g
/XX3FVhwB2ox79U9WU8MtNe9bF39w3UaBzzWwohobqfbfJp02fnqcRKNWvZNu+Ps
6tpkXRaJWUvFKohyd9HM6R1NXWX+1sQ1zkqNZ6M+n7d/wwYDjYjeOtLLKG1Qe4Ot
iwdaflEbXpxxRmIQ75dP0f1fdiMWldXJk4ZiX0FmiHd2Mk8HiI61LJ3YxLbcPTuM
N5PsSLu85MF91KzCwON6ZSBXYd+b3ZfGs9WUkfsv+OHnE9HCXkVLlupWmXkeKUvb
avUdEbQkwvfFTOVIBfGbGxSr6dr89z4m9lFj15N+5ESjsl97Jw9R80ukDOmuoOkq
CVeO5McMXuA5r2mdMRJEgm2PI5/gjC77BIeYCOHhdoP4aq1A1nWZugPNOim2qjZ+
8U6hun29s+67WkOP/W0vXkQ925sz5q/6MXS7OK4G5Wk0XfdpkgbSnWVIXD3kzUhg
dsgFLXXI87IdkRo42Ak8QOQxo0LQLtNk6TJFbgYwO5pIzRbyRtiEkin7h+w8w/eG
E6roXj1CFEMKkzBMcoMzT1X2DT6kN2aQsCROzds1XN9HZQiuYCXu4Gf6EKQ9aYVl
ACSdzvqayNEDzerrOZCR+IzYhWmE93m+a8LiO+faUROktSQomctgbzxc/i6sSoda
k9Ubt1mSE6mZg1KPegEGceGn1e46HEujmS2WPSg4HiNx0tWbpOYJhJ/NKjClyFg5
JJcF9NWAO1CAjUMjpCv0/uLyxX2FbP8BvBG1ZYvNRdZFkbrOpPyrRniro7nfN0N0
xHIP5eEwBKPwnJZf3A+Lm1vby1LztJpq8eUYN13H+0OBdTnKcM9zzOPGobhkC6Cf
16vwt8BNt67KD5DBPUMwmYeQIpadmF5HCfsAQwXcBV68trcOXGtNW0b5ZNxuW6eY
SsW3gCKwWEmPvfBChkDAIulJNGYbvwpoaarK7B4N7tZOL5oSuG4f+rU5smDPds89
MRBZjEgeYtZckgbip1CUIHD+WrkeH9SPUXmukkbCxtYMImy+aSN8xz5BQxAu5M0O
wfCydXl9B1y2BAIl79W34F1nBUg98AKZWmvSzEWemsm9t43vbl53NQNhtBBanNIg
L4DkhFZuImZcc9GmSwHMOo0rE3/nAeG49V7k3Sttq/P5lc3ehTin3Gb6f4g0ucTU
dnkCYjNr2BVib6JxU4OhSoKEZaGmmU4tMl0eDFVg4RHdaxRTLFUDDChQLtl+Vv9Y
z8kV/aunbYiQg3GhYFrj1tzZhxeUDHpVYoOROnEoCUFpK0unRDtnoQONMTNR2FbR
0uM0eHynzutnRxSnps5+6qwNGBRdUMkfIQWBJnIj0huPEGqZh4oIfYyLgBFuwSd1
QVKdiLJ8DPUAGypcs/bSc2VcrTWXFt2NPPhAeUeLHf2Zh6Y6++HAV8P0Pdglyre0
3zSaE0XzozKTiZr7v2WCmwajvQQ8+Sr7moYuOgB47vp75PJyu4+hTAPrZjs9zP2A
T/qJshZ1EiCS2pymvT62NAJU3XcLYGzNA3mXYtDxCRax3wGu8aZ6oT9X9ly2U52/
ki6WbSORrSnDABVDOpAoJaiDazKJWfE7hICJQT2o0CnIeWgxenHJZmAs1XMaSrdL
193hWI3oT3QleAmpsDbde/BoRN0uAHYSjZcbjFfeWE8/aw87tcQb9LXpzaqcftzO
npbTuGQL+80gkglIE7Rw0YAGAZcligojLMC6IRYESZv5aPhmeYp1Cg3khtzProGG
7j+bSI33d7EAfiSKkTANFu8S+eoPAI9kaE2E1gayePZ/lCecVIZ+bDPeMMHYSx8U
Y4hkSXhE2s6xpPAms9A603VaqP8FpoVkOEychrKrLn8NWZowatwr43fGbHHE0V9W
W1P4NVwB1U0JU/A+h4eKlb3t42ZTuvCZEs+aCQ6VDGx9nEwENzG2sbNZSIAi3Wwx
B7FYfQ28OIEILikkyqthgFdCajuRy3iznWh/1DJyWDyRmskrUokQo+Mv5uIhA2de
Nv2bFjiaWlenaw9zuMViIoBvnPK5JDoMfATr5qZVjam31gPzoo1Ia4GIIazEqBeZ
5jjjdrY4f5dp5wXYC755unl7g2EOdBYzaNy61kMnDBSmrTtzC8+wX0qY5nPtyZXS
ciod+ecDbBLK4xLeH9mBEt/Z0vydRKujhKQrJ3nX1FrWi9Z0Hax0eFjRTyM88cvO
8rNI0tjAKigG852726kY/PSlL/kJFn3uYIT5KLkZr+6O8RyogPG13Huy9f/rOeLb
DfTt0rJscDGYitGsSXusCWVieEfhz+cD/x5Bkde1IWZ71n7kFHnVC+rPMqwqw8yj
7y6RJo5uNVmN7e60hRefhnS9VFARE7J+MZrcnLU6KILhr79mQX54x/3tiT3GfTwl
mYysd1dFybHOw5hMKgUT9r6TF9Xr09peE2X728TNGCOodzbCSqALgALQZpAG7ZQC
6lqCmh1GagBKePzTNFuXsMnp88AS/mWY/KpTIvttJPBtZOj279bWm78+WMcgr8be
9vNAwhM80C3+6oIp4iBteBGe7K9hx8pR3i1lpsa7SISbCQjwVNXhvUr4ioOaHd9m
21xR82/Zly+JLbkkyItI6OqaBeYojQAwBq5hvvPOl6n2dPeuxPHriQ5cmiUV3a1F
MR0JUFMPcpX1mwOUDMIZGCb+BcEzwD74YT8xfq8VeWAWPsbw1iDMsQlFqGR1hIE1
krP9BGOeXO1ttACBQOOX6GMsyhJh6X0mU2poo9qXiwk/o5t2tdDCVBHJkZmL9XqX
c3y6QXyigzZNvfgRWrKZriElRMhpNArDUCL/0qFRwHOTbwdR4Iu9kauPVRJhsMDk
BFP1Lrc1CtfMPxJ6fCzeg/KF0EU+dJDeT74JFkfaIpnluSRhr5PcudjJfrZ6NbM7
WoaA/WzXscgTAqgIc2OIbqRFsJEz1u7PaO3y+vlImSVyvkvN52xpjaFjcyUDTgJ7
iDrW8oyT80xY9efSrtnfKgK70WZOJM5riGuZm27WxfN329v2X4rz9YVlo3r8Iqkz
FdfPkl4GnwfbJ/iH2CC6ed9Vw9SozRM+Lt0pReOAJjXrB+Vb8jnWaFrSLJ5OJn3t
kO+UJzITRzUvXc0MfHDEarmIIVVx/LR/7jl1LOxNDeLE7k6vVJngSivDHqIuzTQt
ygoQpc76CGVQg2xEwAVU/T87W1mM161z2EEfvpyb5WLOSLzcoY5df8Q8V8SJy0YP
MulY36gR0uPAfvHNGyTZTZ1MaQk96qSTcc1fkc9lM4uqXvru0cYN8ezkvt6JEXkD
RH5Z7tv6SoY4i4NifT1sQzqbHsJ08Se4kwKvURF3aqp1Bqxc/K0IOmw0rNCDIQJq
vuKGQ2uaLD6zTja5lNDJpWixxb6kTm1KQt1yBoTVowasqxMxVn1TJRTPR1fMI2tD
zEwRK6DnTIsXpclIXVDc1tqrZWU5g1oSW0EF4uQ1bNdLUlM4Dg+vYbn598EKsvYO
CX1u6dFPcexKXe2K11PcXdY+zFA9Jw44Eg0AZOcjaosq+lr4+w3abRLtlLqWbmTa
36HsPvf0dvgXwMmfpowsoaNNjECDmh5uYRCSd7lFOz84um6lgXnaP4ozVwxbmfPA
b66s0f4txuoYL3gFW0pctUHuF3OewCVlZMHTEWHTeMzIHd2r6z53ax8Y2vwxbltG
A9rTNNTLjJZcMiz0ROXtdE8GuDiOcLw1ueZbC0LOH5Fn/YBbpx+Y5lF4e3gE19YQ
eGBp/gyWjOu930YaN3/rm0+OX05ea0bsk3zocCERxo5YxMAY4YRdDtL0aIIic8HL
aVXSTPVloUryBcSagA8BGxQaKzo9rEB3KDAC9yHNsQ2RDaFWRSz5H2X1d2u7v6cV
qrgbE90mksxzBDhBoHnOScL6Orr2g/Rb4AV8mLTYeTepkg+b+5j7f1IllZrD6+uL
lYiagkpt/gpzXSGe3raJYoRzqv5PdZftJshqAxgY2vVaYFe7dmv65beD23qKuOr1
E0AnFkdzCRAPOWmIu0N8Qo5fHBSAHlbhXQ+MFrqgE+EP5frJsxB5vySRvbiAiXof
yLggXj8bvDT8wc0CQAmkJclr+kE8B6Ojb5ftpzcG1jMBk/RRq5pH20Wtl+Z6r6Q9
5RcLmrtTb/3RLyvIo2aTptPQMM652qHK3TQ973hDTWgjWxZ4uhvEXmJKqU7Jh34Z
li7a7bbXYAtGEKvpSNCxsiAPBIe06hGijv2Vj95MlTV79zHrHSO5Y3efaF2u9A2f
iFgclePbLySTbrY9IutBEa+eXCIKNT2vHNwJNgxzTUcNuMaeXEGryddT08D5Xgm1
+kut+sEjilCnL/3l2l0PvdbWgp/d0lOs/7VOaCuGSUqQv7zEe46GoDzAZDUkur3e
K/VrDE6d8IVQPgA4uEZgMqY47od0TDNa4K66JMm5TjqLZR7nu0cnexQSAPCu0Cye
GHdTLb6TRXlOqCEZtN6HBm1R9UkQ+W13MVxNAqNIIlFdax39Wp23xBkSL3VaH3qz
HJ6YxkM9pUnnlIs1De3dYoF48p7hPcjnGL0YQ6S8LEWSNZI2bxUH6z+NwGgAqv9Q
nGkhcoVvneAdukXDB5Y2UWJNdVOV/ef6T1RIOEV81MYTViBhex2UCnsr8RlGhPiW
c1Vp2J2IK+YQ9p+f0NJHkq89/b4aeLL1hWpONSwZ3X/8u6SRINgmRypZOtovwv3S
PMAWNARBTrJaVBxvmyu+qMLoZLw71jZ6YfGyxv3So5t3WtR3whyAcfWaIUw08oOz
2tjkUE5zg/7pad5k1dPemELLa6o79buYEVFMctJ2rB7b/hQmof2HJ/AZINPd1teZ
lGiDewNEqsFecGqU5VW914De9AMAmtuAdCam+MNxL4+tnNI+48PV63W32b5e8bJb
m+0ntjta+yjo5xMzdKSk9QukPerBpA0AuNGun/QDeUea/3+EBJkZwvN2NLlSvWE3
XqLNbKjhms35Xu+9DTtXPOJEuy01fnLsgUfNfDnvZA17D+3AZI74fD67x09+AC+K
VRq5WMqBrwhGDINKU2zVuXYy/BmwT31lrRuILVGJQuoFVVvTzKjTaXobO50xH0ca
fJN5ujlZXFa6rAPq5Xi35N2Uv8REzVB/QyFX7vljM13jsE5Hc6oBK1ikSRqlrz+M
H0+bfpHGcqk/jFBvkldDm/Vtkzd0eZti0gC5ScDpOmEEAU7bc+0DK07tf/GNXLDO
YDimEekiFlL4hVQvQRY/Jqe36y6at0AnkCxSYMDGMlVkiGgklJyBKEH0XnxYYD5Y
yqypalvdWioSn2Bx1WwNwhfNExTuu7p8u+/geA2NrtVHn2RiiOy/duWwP/5udjGD
IaJ7+mBAl5GIb1U8vW/cMbOGLeFmDu/alqT7H6AJI5QRWVsA+B582P6SMFxhHMWp
f0pCGe2lpPiIK86zNuJPNnEwe4QDNwPjbiyVFGwCJgVCbeRGhJTwnwkGCqGgOD8R
zZXD0h754+22bBz2d9m0rzOvCDjylBdUQVf1mxqkBMSZXouQv824E4/heu4y/Hhj
tRLX1f2TelrKOsoUx3RUjwn61LyDsOkIksQuJ5kr1eqTwcVQzqHn/uhbb1FpbpNx
zbwpjHL0OGashEhYWQJS6VVBsklxrGBS9LAvhnMSZYCJBf4CP6O4yr9NCEO4U2h2
j+XBMEgQQMbiZt2BW8uVb9rEJa2SKE6wEcWjLOdLP1iTctX8/TyPIGkVH28C7CXk
+Y91t2VhL2Hcwy7ri+BjHFMAn6K4wmZslzKv/VaThclk4qg6Whr1E+ZLgEkhsCo0
0jIbl9SVxcORO+e+zd2kYUv0dBA/VUZMnQ/E6d3hBBl50r/RF8l33JaRNWOKxzL4
NpLgdos/2zh+8zO6KYcJ0rL28VOvZ9r+JZc4TBrAf5VynBXl9qcgx5lxFQJrg3sL
3FGyMu9DWQ+l4WQn1jtKjCogHNVDSfD5quT2aYRTVyC2HX+uBJZGIuKGsATfi91Y
DkKJWCiMXCu82cteEI5Tcuwa3uY5RgmYmmqXLwyrpU8LZk+1LtfDf3d7QMBuBrGV
9ddyv9rw2vnReLMdRrQF3HjAAepMoSQzphz+3d83nXGIhwrrgH3HKr5AavysE8CU
yNqTLEZGtpq2/6nzkXF0Qq0ZT9n/3tFdamRNFYXk80CpvKasbj5ImYjL1871lcPb
tXx5coGFrBTniB671xc/Ppi1MCnj16IDEJXY3UYEzr70qxjYExkywDHz3jq1CcST
92keK6S88fKCAC27sO4GWDgEnwTPwWmBruKr/wh1U5UyoqhCThiEYzWwINXYhkfy
D2NkMwkZX1VeCoFHWIz81X4+TBSlaM5riPHf9xiGG9DvvBxqXs9xhuz9XdIHC0Bm
YHOvhATVY6RXRURmvNBy0N7kT+sQTxWHgFh/A/zjA84GbSLV/t2z7UK4u54td8cV
u01nwJEVs1OtWFWzOUScBzGlCBa8OCe/2Wcfm9UvuvIFNgM9nxN4jHz/l5L3mc10
FGJVLZiBQT7k5k1Gf1htgBMpcmDKFhZsh4bpz/FudgRMNhgWNsWt4JZJl1eq735b
AyEpDrSj+BNrpjwVdBx2f4WjhvgWCrIMcxmPy4MvG5fV7j1/9FMNwwQUxoc62EZY
gFW+aQDycLIXfIKPkcnTRVkOb7zcYEui4k1np0llrjFb2D6qFRirX4TVvI6bfHtB
0mZAAApn9lFvQ4vOVdU8NoRsoMECUXVxljUbIY7R0kUAErFgu4hORibM5u/Nnjr6
70QhGr93roeAJkkA4lVfBBCvKI0l0FdrOztanDxxqh7TFtP0QcXzQIXKDramEuH9
SSWWtD5fpTZXTI0peG3KMsbuDhQG8GwpW4fya24Ijx4N9dBf1jlFV8EO743+CI0z
NO31u5HBEDwvbfZcdE4w8BtGshFmGM6uUyY/mFa3bBEJOuEvIAartyz9rGlGSfj/
KfvttKadnPKKJuZx5Bk+OClVOQisYrUtWItyt82fyKVdmiGWSkiHFluC6noI+Pra
udMl0poihZYbtJK0EYz2TjrgJOhcK/Tiy7no8LHyOgXRK2zbodwv6JI/XHNKmzE1
EsDNEhcS67oO1Jh/9VrT0tPIhAVLSDgdxtEpvvOBTnEWSv3xr/7wOLMZi50JLv+4
mtWSRSrSlcFnrUvwl4u38R5T0Aau4gxTBp7BNfzshqyrWVIoGTPEuAoLs0IvyW2D
jceM0DKQrDZOjIRx+aLEqOg8iecE0YhYSHRLY7/83xyYw20wnWamPcVay/wSE+VN
5ERIiKEUTLwe1NzZ8O4T1Fl3vR+ULWkOYOrvSMrvVLNFbgrh8x/HOjD8NXy0CkyG
eppCLqGJY1YsY/aKH3Q3KZZsQWXbXQuXLqLidPDgJWzZBQH3ctEoJIVP5d5p7SRp
zcZ1BJv3I3F6mrz1NEqwgN2yZ7yArs/+AnIBwl1/q5Vo4I4m7kcMOLa6QeBBkRi9
L2oSYwOCq/lW3y/USuXbaqph6i43tPSbgRBnmnIAuJ4240PEs0yC4/OBtXUA2o2p
qGlBJKG0TsjjTdaE75tpVeBleB+I2j2MYH0QmAKrZN2MP/33SbLp9D6ia5+/afMk
59GGGaTZaJyVKz5kk2G0hZeJhzDTG7xxNJd4A0wl3xnLtE3w3xfp9AUUJwtBL8yQ
g8BVVlcabeetvtKfBbtOfvO0RkCSS7kvKMuhaztiyjW4SkUWgphZ9Gz3sgDlETjQ
tpPjeIOYeP8gv6FSixn6poClw+k7mBlwjEu3GPhXnGkHwfoISEbRAYy7XtNrpFxm
aBhvMzLpAd18v6hW5yYrkZlCQl2XEa3+Du/vFB8I5A5jVwaBxfntsG/PEz6jElMZ
x9kUgn87DtWKGrxqFVI8Ay8A26fN++Qz7w4bxOikBzYfIAAeciKpX+tPKM2CuNkj
CbpF4bVy/ZABUjRoMoZscbwi02fWk887kRylzh3RobOkS1hsTYwnjL0ilgUXQTpu
T4QDYHf4DlJP+IWd8WCDUHjCC9cAnRAAmWq3JgS6uQkzVKyrPtEaC2otUW2zSOz1
85NOwMoejB2x1Rg7x+OYbZMB+Jy39ukHMwXaNpTwbY7rrh56sEnVRA90cqv1J3ls
ULUD1WMdgpHBupJy4hWZq6Eg6sEdYSJJ3iQtWhwDhBzAQrNELa/HbskVHC7eBQr8
j2EMuEeKBXl0MQAR+vhiSaxvMXHhV/dkK1HIDswo2+49cz8RfAPDTfk0gBhM9OMB
rhmE7zYEsPf2IIpOq/uUcfIcYznnIIlhXGZ5deuLPkHjAjrEfZTApUwpPe10S3Ws
ehA5+vLD8zxuE1CP79JJCfCKyy4wVM9Ga19UnSZzM+pplYrTyb5LXu4AydWskjxO
z2w8BUDfTwd4hhLfs3NDoR913evLYkzuqg+bR3KXn3FhAs+kWxC41Jy6zbM8OYT3
IUQMTQFyT5H/yB+8PSv206Yx6dVYERk8ABUTUr9vLqXHioBX3cKUakYK1CfdKDpp
Hq43LQ9eWrXom6S1jfUAAKRPgnBUjaxFd0HqzOnQ6NdxWSQ9as0k9ryZWhoa67LI
QDc7cenVv7ejV++DUYZJyn6BgvKRUG7iBiQaNMNhmUGaL6TO0YAomgXJmLMiO518
4uNB05vkRVLFqf4zRkrX6z42hP4ZjyELvSWXd8IZFGx7SY0nD/6mFD/oeayNdDPL
oMI1s2zcl7wpQqHalllbavcPLVhBFqn+8/VcdC2fUENAe3X1aodepchs2vynCib+
jzAxsrZ0pad0eZPwgmqmL8TpdD6sOAvLv2uurGMNWCAByxUdnmSNQ8M3/ohmglE8
Bt76URcA4qv/MspsemSB9al50pLvvDG54ejxJ/eBBDIkoDC9XRv3Ud2vna6qf5Xk
IQp8oZzR0VON9Gx4Gwetb3B4BaA2Imb9Jok2GPQf0g6upzHDJKXYs6STr5X71XsE
Ak7vkWVgl8yUcgxdlKGHGFSDSwgrDMKJjESxnko8zjS7FrtzFCbE+8+Tubom9kT7
1GijhEszMDRiad2c5fHyke2L1QOGQsNVSXADdhUKUnH+krWdlEYhWymEwejQiClv
Bi6vswA0iFpRsatiMHhoomHUMfPDbB+qP3ToVxKkKFvYczIIxwS6MYx7hcVjD/U9
QYuyleqW1ftrhyjNsW5QH5bPXK4I2goYPpm5W+VFo0XOsqK4LN8PUy77KJ/1PKMm
vgwI8mtAr7DkmoKs8uEME1hFUh0fPwJrm1Y9ldhCXtzRTn6H3OP1r9tzKvUUuHHr
BQL3kgbvKQJ0mgSBjpuhGV2MS19+uhalCvgNhSJ7/hpLx3s1hcnjl1eBUBt4+swA
UMH2WqIcRSgrMJuLLhGUiFdCHdqZ3m4PDpzfqRuJbyEQAgJHhOlXFH6nlz8ZJkZa
ZpRAhqhEh25ZL0G+QHd5AeP+tppmF0LYo8DpD8ZTk5vyiIEQkwUCGnfxpA2sHCEd
tZfaPyfK3VgyD88xDakXL83+lJuZDofV0vyxU10bMQ4xDr7RE19T0KuCtaE/rDnO
U4WlmVnIZprIOs3f8b2uvG13om4DDEJWKC+1fAqpLP3iUwwVUQ6dlGrnzGBXKg69
rQMn33D40ZdlQKFCKvlCYeVSxisXUdTxHohUfgehx4lyqbPfi8yJKk6nGZA3oSTG
CMfIQVrW47BArfrp6Bp8cGqEQvfByf1zkObEBSzr0x6NpxW9L/o/gKIowzTARZw8
7tRbD0ox+66xSugh+MLumKKw+zLgyWbQ1Y4gCOVJ9xJMyNZEzjVui9VGBaPBtbax
P8/iQN/9lTjSFhZ4wp5rmDuPOF255N+Ui2AJFSs4cn+uY3FHlzj5qLTKCXX+bsvR
8kGK9N7/ucSfxXgSbDcQBm4lG5kEZ0xSledRk/4DIdJKxWzX5o3K6lfAKv4QccQh
Ch4VMKbfXrKhVQ0G+Aga68MpUT0tsbvEzFIIb2Ns4FtuB2tB45E7C6t9KRh5ONTq
4yNYYC71giGFDAKL6ZTS4BXvlzh3WMYiel7nj5plS+8LW3xinHMab4aqRZ0PwtFq
yvDEWUOdwRkPr4NO8TtQKW9SAjxi/W3ffHFVoICLBxf6AbcUx1DALcmfQVfcK0Ob
bXbdWk63edEGQZXA67yR2JyjsMW+UmKutWUFXNTHqi9inMPh6fUa29YxfmMojvCI
8NWJfFbwfaw3cNeWUe576gl23p1C9UWLFUk47OGQbiNGgZ4vtfrPVGaQ4NXaCaOT
41xdb8Fzvx/RuD0j1bfxgzxQ4T1YrxP8GZBaHCdUnfY/OpZy2HWcEgbutRZGuOsj
6LUK8PCEsXZHjUZPDECt1vMBL9ua593O3tPhbEItURYYsX/Nkx2QErnBRXboImVc
Xg/bdeqL6/3ySEdjIhENayobp9/xjfKrcbWQoNM1mIBC0XhyBiOX0AtJ89nz9JRJ
rMRGrpDg9OZWlQVbkS6x3IlZrV6ifMPxNGaRh1lmtqov2723voLPKfwBRZSN0+5N
mIP6bUx8n4vGR1zAA/y4FdtlPVKhfCvQ1gJOVC+XcLcmOYFKIYaM4s0YMX+4+kxr
+ZVBfg6z0c5KDMAU6MOOTxE+TTgI70FwwvKBsU70bjKgMRnuIQCuFejIoVXlAoST
01xCDVCduOz5tsdGu5t+/n26f/EKk31R36+0p3GT6RSwmEzHkpu1ZcP4Yd8VThpU
k9UVA/B9pM3y75MnkuQPGyYHUK/l6Vz0QdvRpe9ujz//VDIxUgrXyRW+YFRSFi+H
3R1LLZ4f0RokyjyC+oWqH3eTljuljWpF5lw2KXh2cAL+Ctlda1t4GvZlD8bvagxZ
ss1XiAsIR1mQDpPYAXjri5cAggzl+spBEI8dBRWS9U3wCYERfPm/NG4syqiWj7Th
PukeU54mub03VJxd7p/O573fwlQOHSNtLwByot3AU03Nz8szaxtv0TPsoLu6FgwU
KX9c9KYfWPF/LeLzS5qg0Srj0cwu1f5vtwwexWv41y1s4QeuvXCN0NcNa8zFDKPy
IhoCS+qwUKy9Y59ueceAFHLNXn30fEzCNhReMh5hfHzQ2d3H4+qSCW8Z2VEkV9X5
CmNTY+WiYkkbRiQR5TJ/of2qwSPiG+G0m+qVaR3VP+ysOsAA2ho9YcPeXz7/uNym
9nXmSDnub4b1ienIKaC8tEz24yTJ3+NHWzzRr0D0aiu2jWxYdAkaSz6vKjsWAIrg
rniMIuAbIuuXovIyXkD9XdMV1p3QF9lf0DfRt3goq6x3pIGUdAGF1bsWVcy/Yj41
O1pXGZ1Q9eJ1UfqlHazR5k/euxKy8QnElqbTcdj0WuLP8VlStGgcwMD940qSXEf/
7syNSTcz+//d2J7RKn5j6RquVP3Sx5vVu7wYbvrob1qGe66qTS8nCt/pDijkrjHl
3AbOLGy78JY716lA2rlBN1RJZB2F3dTntAMypTpyDIZbrhoQKJ/0njEzx2FcTOcB
iWdRe8rb39O/bV9oQIgJHHvsAFHuVK8LDzlYzXjRq3PoH2OkvI/YNhXuOnNsuhLc
kkoW8Q33q+rBUgARTB7eKevBbKa5Z2O7DRDj2TKEhCiH6BitifX/4Qp/JcvNifMc
1kLMh5SEHIW0Uvlq5adsZ294VSyUjVkf+PMOXl2T+kwQ3chLwht9U2nNX5DqEJWO
XmJuyzAOw0KmoZy5mW9dNogwjlL0Kqjf730ca1y0h8z/6jOOH9mCsfuJOtMmqqxb
lHFK/HaF5dXhmX/ANuVm1pMDzqllqhMhEICHFKZcsjeQw07jU2HtmUH3EEmKHVO9
gl6AQZOOXLy27W6YVjGbT6BCBxRhx8BTJBrgCN8p+XcVgfk9A9p8yAQ8y7bQ189g
8WoH+fnnAMcXSbBBOKAu3tTfceWZF6YXe3fYfGIftSLvIC/q+0Aa7gMl+kDkLSjI
e4uH3jdFj6gO0m5f5NYmlzcbawdnlWYMxuWqECb8z/5QQ0z942iVWUPdUuBBCkwq
2OKwuY3mh8DY8EHBYQjX+LPDyIIl4FpqW+jTauD4jHcvBNx4B7ID2mP3evVDPWYM
d43oDgS/PS59E20tGRzBPNi26+AyVDCuzk3vlC5cvZjlOLpJgOGFlEs83px951Jb
5NucYljrvJRSG3EpOPf5mWbzzQ2qqk7SXAokAcLLSl+YDL77o2bG9M0Oh0jAcmgv
Y60D+E40I0/ieZmkGwc4lELZmfceG+wrDzArdEhfuvkGHlUL1HsZXTjYwq1BMQZW
kK5diVnNjB8hDwlU0GDUYeripjtj3KMXPEgkv6WGGkcG58IC3h9Sa89fg97R9KT/
AY4+PXG+EukaveaPMcWGzN+l6b4vrQ2bQ1RC/MEAbIxM7l2uUcCK2tAHwC0gTivi
brjkkOkoXsMnv4M6qac3Q/4eK6ATFLnygaqkbdScw9B2x6ecZ3Iy8F9tgTDRcKwM
T4MIgEAv+v1WJhth+L55eYYohxj1tYZ7SSQzwd4ADdZ1tkUec7cN7MRiIAn8r0WU
ViMPsGaRi2NlerYgDnCjVOFpeUIpHW9Y95J7IluT78GNGjFxzGXHGXmZQ8RruHpk
/AAtsU+4NmyLgeMi3pzLFHssyb5YN15iizJqPOrvQ9xBR0FTRTQiykaBleT3YyT+
gzYKyzTN8PTWt2dlkLeqHMVqvVLFeE0AWBFuhz2fxGudCwpfM0nzIYg5DNA3xdWP
ZAaGCTEn2QQ6G+Y0j30yaP4cODni5vkoMJO44TGWHhBSyatrtFNO/UjA0lGe99Q9
0SWVhgbSgMfw5HGwRY5N8Nh09ZgvkZQnxLIoi0RCeWDBfjCCc6Lftqr0lChj48fg
EAMSd3Cec8eDzfpHXVKgJcLwXK0RkA/3Kb7EXWjr8F/oaRJiceYN5A83kCIp0bVC
ZwMOQkaGzSJg5FA7l40k6gB1j09gCLm5RJzvKQ95zJ2tesZ/6JesTZ/fDJzAdogH
cHdWfeSw5iJqZG3xfgZXil7jBQ4SiS/beUHjdNogvshOoaAgGFrk5ML/wnXqIgdn
4yNqr/TJBl/RsuCI8PXaUoyuHZcN93Jk8WDadFNf3fXPV0PE9x6QXqAa3iHch+w3
UhPjWeJi9TK7XZoN2cz60h2PQkHfiC3VjEG0/YWKECPSpJdNV5WVOZyWtUNkCHuM
6VZBwlDZ9XUZR4vness+/M7b/vZscW3pi9LFVPZ2h55qNN2G43mtQwhJt36N6s64
ItlxMGE2jUbscphgHvrcoltn1ktknWmN/eC0a/n2OHVMP5+5PT7hyCK+BYc3xR3+
Zy96FW0dTSV62ETi9j5sZp0acYU4yj8VtnJetubBLQPUNE2azG0QOP59brldd+R8
xektDHkW4IMNz6xA2roHC7V3r1meIUHC5uMV/jUhrgABA+XUSHHvEOCpSAFwTAgQ
vj0S+P4716kqVSw2ec4CJi3MA62iDbIQ7vqmsY09biht33tk8+alLghmRvOBRTRk
VbdkgFR6a4SE2zXlVriYTrg3DJiH/koIdmdkV8APQOVKEccT86hh5CsLY3x8iRQm
GhFPptwMVXGPNOyrmpXQRXxj4S5E3CH448wsUgUYBCC62bIfriieyfL+H7kvRXZL
bdMlBEj2zP3sCDp9V/ta8pYkujr9+07xIrt0UkCUIKH7EBHzKADQkrSjBNDdNfmT
ItYJhFy/Civm4Wu35tXewq7M5nmPmSwgzRUcGDxE1xDNGH20QAWcPmFZPiMf4Ii4
T0ILUKh3DGV+Xej1C+3E0vwqi80cBblhzMRqTgBdNXlvaFpnxw5Cl+RT+m8g9phE
an/Xx8BY5kSMvdbEc8+1dwOr0wL1MK7hY9ZUcKwzRvRLuE9dEhn+hFumBmQDxLsY
jY5EiXd5623PGjvGjXDaxZmkmuFl1ZQpdNpH6yH/V2fpf89crsK8irHK/6hOPYXu
wAzGBwddq+ZI3yw/jN1XfW/PeMAC1dawefqEokEyvWzV4AwdHH6HvXpIUK7uYmyd
Qii4PoK0vhZExEcwMaI/B1syq2SUjvuwA+CEXSR48OfyOQfyy8N/sPYNhSQz9/Bg
cCdYFqzsb6MejzH9L9pOCTNmnMLFmYHMVkg3hsbEbAgYoTpQFOehczvEfBKqRqQI
LnoLcQT3c1FgbyodLTaC8MWVcRCzaUYdRZsjQAn972cXCHzMrzFLBGk9F3egfiV0
/QKk/l02UfHMujJRk0NZ4TIs+PTGcVhmDziWW9AALa3lbx7MlcI/1M0TP68yn2SK
mDNQzXwKnNmt1FGXPpU8S/Idz2jNI61nBpdwAB+T/3rHxu3ZwpESkItRuxkieD96
ya0mku3aFvGNIhQifw28Al7HK1iwnWZ+ig5ZxnYDZD7dNhGRC82sCWOV3UZg9HoC
0SM9pt3UhXTmlDKOBXtZZNbKupYCS8e/E3nYAumQ6vp4ho0ht6ptFSZD79IQwqsj
gck7Hy4a71M1j6CnLjxGsjBesz6vF04n7GPmkiR0S5QZjMT7mFKoJRtQNEcydb7c
+92vFbvrCgPd7ONOU6ZuWzuiG5o/l/iMH0RiLPiSbmUWUFt/ZV5gIpOP5Y8PY45q
5WQ0HcLiisriQJ6MrOfbUMaRq5kH9saWiqctBJaxFO0RBX5EI4fJ/xYC12yoOZex
mYH+hFIeHz0gYV1SdcvrJ9tGrYLy+7xiLOl3YJuVv6eeBrZkMu2+qA5Ob1HtbTI1
v/iXZFYYJ53YlbDYzMaeByyHRxBdv0dUuM63RrVLA0/zhrFX2EU87LA1ZEz6Xvro
L7cKAYJ9z8YxTs17BwhGOVS4jsu5YU0m/j6KB0+pCN/5RRGjZeTNIsdRnSbCWaTZ
jRs+5yoeR6HVtWovpTcoZcXl6pXWDcM/OvxprHeQInhJlL4J8y6B/ZsNLViJo7ep
PHt9jgNXmmfLd3t/GxHLg0nYNhhCZrcxxRM3O9UyzgTShH6gbwg5gvUCxXU191sh
Ua6xwYXRJAf0nisj0z6b+1wyBDQw/QJjuZt/xkDddvz30Kt9pnbsLk+EMEgPzlrf
bRSQvRaxzRb20te/JtVXw1lS/4yL+aA0VgeX6EynAC1ntrlbk5D9ieyHB9ZbAxAN
deLH4IBzMU4ulZRmLUyF7WLuZVN7SwJGFSt3gbizYsIAkDveAtRKQyOKBbFgHhR5
MbRMqPwe63pdGle2MaYChwHRsfeE7+sB07FWrWrjyGXaCGIwW53zs6gbLad3MeSZ
a2GM2eR9Up0lhy6ouexlHi4JfZvFQnEXgJsQatxs7mQOB3lgtPjSsfwEAD7jfWXT
8Q/y1IMu2F5crlmUJAnXgaeusc8G1HhevkXOUOlFj9ziRUsFzkiSGgvWl85FJNcv
Ok1G4WALcNTRIKUUAwEh49qppxHfsfafl0uPZ3XRBd0+xhlVaH0TKD/tK4++ptHq
VhkFFPABjHm4dvhUef2s8jS4afN60gq17Xr6/q0+s/aUjmecG11HHbfCyI85J3ia
HD2XxARXFM3VFPEMBjAnKfMfz2peG1QJzFzzkjwls6UPHbHBIXFMqqB+EUdfvKMU
z8s1xg2QyNEYCb3BoOjzo/41eg861GJBUMW25tZ8H8u6YmUqbvmrCaya3i/vE/Qw
1DP7nXY+ewvO+os66l1m7YRurswBA4hMloS27HPpxHICoKLWgbZ6J5+26Emgukfz
MQUGn5QH875YJg7ZbmeuDNvZMLpJsvSlVCbXu0hf+z6pl+woSUjlj/gURMW95EiQ
JFKxWLllt/lLe12kk+mYLA+2AzRL3lwM26ruC7LsAgO7zvdC65sHZ/gviEs/+wiB
WoQ5+cvb2OdwXCecp+Gs8lM3uuBoHCxUtwIFarhiRQ3JI4RuYd4ZxiHlTkSWxlN/
sptCMXk5dVRAq4G2sFwpJdrTYko4EUghWerg3MazW9tkSGJ79TQLl/lo66zwn2K6
OREHkiMOcKrMIIiSQC81nwbeCZFSK1t/k6o0PEi9TfaJ+YJ9r6cTlNxoX09BdwKf
IRAB7B6wN6q2Ff5HE38Pptwe6yMpSzEALeEbvNxW4c3yRR9xsQKa8P2unJ6F4PfD
Y2o/kOG7UhYkZuNnJBiBY98Z1p636gdDyr056Ug47jciFmww1L10sHY15G1suf0h
238NmF8rUdGIVYR1BgKFYx9r2fTD2MLIPwEb+h2WScNcnOh9ubhYUCufChTj8qdQ
hVfJuTMr+L/YI/pAJkLyUcu7SRIUjBcDBJMD6qVCg1JOP1yoTXZoEhleeld1qLxZ
GnzavDCUlGONTDrhJEbZ9kz1uyn4Rz38Mo76bgrLpJZZW2rm6EVJNf6/RheKYsh5
LiqtnNb6M9UdJIc89aL9Ld/l9xAUlGZkwMSIWINvd+t0XKzZR8EHryX9T27CVk62
2rzXA0xhx91prxz8WguRtwYmUfTVZ0ajXdrXgBCT79VJPi+xyQo9B9BWK2YyX/2h
SakDI7hl1lz8GTHM2CQSbzXAQxsGb0i4LIIy0aTHxY1rzbyMl4GWpWpq1kjlrH9c
vQ7Wnh+ribPTjoQNV7h+fcJBE+u2mg7jXwI3S2wov9DbLG9UxBTrKIiYNwSyto1h
akB1npC6+AW9cJvF5hEIbWiVXzjO6vY/lAzdLzJQ2F4sogn6jiHNC6YlJqdFcUlc
QsCDQKZ4WwSntCRDnWpB6i9YchWV5dJkyvZCsj9Dtyje5nQZNgaPhhF+X65BN7sI
HjNiWP8QcmJEguWd/W7tKVatz6rYv2+jcepLXmlALz22smxm4bpSJPFjbcZKPyvL
RabqAGwKmBjkp3FDGWtoXxCUeCWJD+lzqpksS14TtJnhsWgRwerEL2KYcEMPQrBO
2QOxyfvOjTQHIB/l2GTBAI4SiBNKsvwdiOpKBI0v5RiYiNLwLKBiTO+lNw9ms6ma
+ODxprbwM73v7siUVCyff6G8TfutJDyPYv11Q+PtQscE+sCZbPWC6e/RZXSfYGiA
tafh+yqZwpaKfflO3TCSaS+EYUJvLqtjcLSw7aviT0BUuZXMbVDghnAKwNO9wG2D
NAn7S0bf9TIdrQ+4xJOOIxzphDsdj/2OPzX7KUa0nAsLBW7H6EXFh117sSLhBOUD
tSCT/qDUMX47onVX8nHAHs27UYNrFEVb7bayCL13NmBXYbcJMt9BZ/RqBTctK50k
ZYnQ65/ju25/j8OyinhRNnOTT4cNdqJ/VHAF/j6m/Yt/3EZG0mkWl5BMBiDnE2p6
hl3K8/mxUPqpdBnx2tVEtqpKOA0kSWMXv4aCAxWszqwoBohF5athZ7b3mhbNQDvy
g9+YYmRonPVABsv3JaI8dOokP74zMUjFJxeB/uYmSq94qavkxP6wm8JBSwWRxpNc
46Ou2INF2BbjUzVsBc9Kb7atSocDYjBc0KBofP42ukqZr7N3UMIKqbnQBdwqY2iL
BY3LIOvkwIHk5l8ulybZYNQqQYStw5F7Db+Rlt2g+4LkWRv3S+lNGftN4Ot8IVIc
2vslwFIAoAXSoX+DmIEEXb+5PSIn7vbngetWsgVxSSh/TU3dWeSzbH8O57YA2LBB
lWtAcpcoBDObDLwtIxSIlr0dSaTUgXi/jeFm8DVrO3Dxyu/fxuwxVA+MaEM3Q/of
5PwZmQm3Xu9cq96o6EO/5OP5jJi5YuCjmiWhM4fiKb5pWNyxTbSxJZgeZn1M8f2g
2SkNX7xkflLZUC+d8PaIE3DsyEDB0tyME2nHRx0jzZb98J4pdzl6UEydd7UEbrZp
i78zNav5RqW5xmrKKjrN4tr5qyMY8Ev+T/tbCGp+aKgMmw067Cp6mjWr9MAAQAxQ
PEMLZxIzLsHX7gjyPWNALbbnTpF729espLSHzFBcLCI0lmNry/8CGMPdGw/+GQjM
mPs9HLZ3GxCbILB1dp/vD6PJNa9O0hwaP7jYV7Y0HUvCBp84CX5ltW0KE1awWcM7
9Kxu6j3bArwuxqNhTd29NmqvOLICaieOE5xBc3b8y3TGLlHiewCVqMhfuV8Epbhz
z1rVYqJiwcfSqIho8m+y+zDB5/e/4onltiYkPZZzM9rQciMqKajJnmIQjyM8egOF
JW8LwoF4zV2uCxDXNn9tXbGQvSoFScjavN2vuSUl60G413z7+cYfEKcODxpQeEML
pAHYER3JSOys/2ZaPRirYYKu0+pJXtEcVSYmHnEfXqHFgd59517nn5tx6R5PAgDi
Aa6DENZXuuUI594Ic28RECa42eUDqRUOPU72kYpDZxFhkHWrsKe/EExNFl+oPi+w
DJ4vilqFt3/XpynYs3X7PsJ122i2OjwVSltGVQ8DqLDymTmGoMKF6zr+dquJahkq
K6REbHclPIkCvznTRyho1UGBjrS8IxbHJ8lATUTFU6bH2P6f/92q60oceQEs/J5n
sl+bVXrInqgsecEoHUGyekuJrqx9RI3r0NQLt039vQa98FVc40NQmWOnxqmeVoqE
CTplS9wvttfgr5lI46d2gNPUSrXTq9mKui6UP3/Y19pmm8bc2sEgon5UnBaMTCzI
ZeZ1evsAxB8H+hYLvSL0/xrXGYwsgxQmO0DII66aqpmouKSuoC+1LvYEtoPDJEP4
osnQe6Lt36f7W/SyzAw/9KBnZ8aRbakwhRTv7r1NXuQskbFhKrnBg9jMY8zT+WEX
YpDpJesp/I6p1DujGJwP34Tjemf4+vNaczmbXE0BiYcUgVIt15dsYShdc4pJVOy9
MJlDDOj7+g6+eKchB7NMcJLwRTBg77TscFg4uNSUa1K0wci3XLwlfF+XYIZLzElh
IfT9ZcrWp7rVkwvaBuQi6cV5GPwSi0EQMU1S/2iBf2K8xOx3cKbmtM1+p0vjHFrN
4wB4hWuT7ekwWS/CRC+zsaRhF+l88UfJBqPECJAjfzr8EJLFzC3yO0Oa4CXLtP4D
Gd72rbQy//ZnEQ9XGncmGlHrL94l6Mat8VBXtgbI8WKr7EoBJnG/+wdQJu0E9Er8
8dQbebcoUgEkmg1UcSAO7s0QqIn6GAXtAwZ5RQuZIoUacKtm9xEKyUec+bZ+vEx4
al1nBJ1xX4WeZCuWV9J1XfP8L8oz5WvMSPp3tPeg/ffUiEMfjXOzhDHMZ8mLdgh1
tfwz0x+IlG67XX0cNhdTk57x5kW0RhQh1aKJzJOYnOoQP7ntuMi/Iklpni0sNC3J
7u2LopY6CbH9gZbCzBvlSpulM/FVEbGU3DdJVki9bJkjw4tQCtNeJ63z/770Ih9l
1EXp3fpogLbcGGwbRjxT67DKOnbo8yjBrdg3IBuVlhoc9FleEJvF64aQMyfA6T15
hiGfESbF+a3TTO2Kp3TTCu04Bv8c0jz09/iKqsYAAsYnz/nl3WTsHT7F8NrRjSoV
tlK0B4NgokfHilgQq+YjhOEttUbcY14ZCzgK2RaXlkxDeIHSCK355kMWZDUYV0Yo
JylyfGBieIbX+Mt8q7Z9p47TF7bkkH5UQMh4TWZDwKARm54x35vWz5WSfJqFYWPg
CyIsWIvopN1eB0UZLGe7DZKQ7jd5aTwh+luSvPqYLJezel9CHSxr6xmuW4b3wtDJ
j5UG13hV8fDTjSOIU/dyGzbSCgQJEKZfsixyHel+KY4DAszqzHy/zxIJ8BMVP+2h
TdMSxtphYQSWo0ajNrA4Zg6q+DgMtAhYQT1FXPAfOtjGXfehIPGxydq7noFngbYB
OjQXwN/coX5GNY3w2cgwFckjuVMTsFCnC1I7T1XU74+D5KBDeSnnjNtZkvI3CiKE
BgB6ZIC0YKPPVrW46M6UsEaTsAALxBT7Q37yLTPcQs0J6IsVai5ep4UH7EvZyNYa
JD2l1DeDIEGVKPuyqKal1E6CslL+O9WbQm0EecrRndGAtWubalBrMWd6lt8d5WaS
XiUYRSd8fZeSrQRC7cdngC9fsP/dNugM/BySdRAavvDE/xE21kCT+TOQg8TpbP1f
FFSyp6Han0iLwFGKf5lmXRoVQqo6fObGl9nO9wnpUEZ9WS/u9BFf9Ad/RtAz8s6e
LkY5mLr/DlTraHVhOf9+8hNSJQt/OMOWxziuYYeMj/owxY77SnTmJIuxkH728/Lz
GjJojSW6UgA1HgwpK9mVV8X2E53izrfo3pQ9pF+H2zUNy1SM2spUcRKSTVl4/jZh
H4CumxxGSnLGQ2yAknhHyOaksiiJ3W4BXcsGectR5fGtMK0u80iPPIhWi5KRE+0q
xsAkWtBCnbeg8aHBqH+BKqOjazudkOxsH/iFAmYhk2HQTQY4cB4BEBahmOGT1VL7
//OsloX1/EyC1zBeLCAYix/mfKn4MyZ/xMdqGiDLLObYDGwM4/p+00Qj5wtn7HhN
RHfJXNW8BCkVQnnNn4fmsTgnUDXRXecsTwFy+Xcjg2gzpycbknhyM/r9OJ+ecUcA
HmBFas0QQeRCe0yTLoSjQO0wJ1878ZjgbrnJYureWSLaNcS63SuN8jI+Vm44cQ6i
aTV5kinV+yhXL54ieekQUYBspvanhhQtydXxZ5bUJruP207zYvP9/3NSzNTVlqRD
I2b8ib0qGY53k436GIurJlpL+KQDnSYHP/daVH5Wl1ui4GV1EaH/Zzn8KpzMsDyb
SBdp6soJs5dfpluvCz7c7adTxl58qb8IVd5lI7TSbixCi5n5g+imM2VzbYGjCCQt
WObWelJ6rMaXWWIpSo1L/CFl167yUOD+kjPvru2XCQzLY8HJgbONiqtZCKb+i+ul
q2vXlyoWWU1ewBlGquchUEMesr1dp/o6YjasYjiC7ny9W3k/t+5yO2H8XDuqhBkA
tuvgFnde2hCfqlI12z5axfFlvnQZb5835d/uDhDGRSGs5BrOF6OhvuvGmOyHHQXm
i2+WKt7XUYdVsiDBr1ZqXSqX3TQmD3A6ledeu+UdSvbJVBOAOTID2GJk1icKZkPS
i4rqSl8gZJWTs+7I66yvH2hEFAINO7HHz/BZbhnzM4jrQjbv3/vsQoS6S5XMtxbh
+qpFOgz+RqIaQKBYlZAIqctyp9OYf4r/MXeYhk6XglvQwCtbE78C/R9cOnLFqxkB
FZwzZMyqugfBDlsiSOSY35G1BpkAcX18jZVIbCKTC6ZN3zy7/+GTpQQCFAKyFyuM
xD2TXiZr8T53lFoKendcAcmtlHe69cds1Nfko5b19ZmaJBk25baYqKVIliivrES3
5sjOcyg0DjCmMRxWEFlrmSuusX9oO0vF7CR8fz+52RcZ3Cqq4atLPbaeJYVImjYj
Yz1TIscH8HUfyE3YpaR7vcGFAL7Ju/VOsv/x/yf3IZSsg2lyGr0MJL79X08T/XIg
fvPSgCYjoaliLKHJu7qL4tnzpoUW4QY4TzzrK+Vfo4WD1+envcJ4TP0i0+yEekx/
C0kk4l+Q/bR0dq2bEp94Rwy7tPPbi6Hh83jNl7+GVy7CnnLimrziWoFL+VslT/+f
8ID4UweLKVynLimVqtu9UkhWajHvsnVuGaA/WS+BokrX3FmdBqBcJflyg3+15Ffg
ytMsrDTNROkt5RmFIw4T68EVuDyX0D41zFl787iv9JD0YXjHtkFbIqvmAihWwy7L
DkyoGr9c7EB+qCCnWOiI0th+nnnpcxSW9dZxJsN/s7CcrDSmxYxZUJAa0FBQPtvU
prIOqBZptbgzX/DMP6ZIeP84SL3jufFnVFNWF323T/UN3aSgkEIRFKJgz3JuJ9bN
fCvJ8CKZOR1TSnoToFjadOcXV5FQXO0U4Jahlg+WR9MQYXgFrYMu8CkY+UZ7BOnP
JjQ/KKKZlJ54mrdfyhSwYsPsPoq0/OSgpRubdwI72cBUccaetyskPgRKXGWe88Ln
oXVZT/L30i+8U7XG7MiBtmoWPF8Z6AF0PZJvLwTzuJAl/r8wJ3chp9VNCp59AiXT
lYKugdJnxjrFjA/gTxKSTkQK3ThgNfwl6Tn+1piEj6OYKrUmTTLcBSjstr/URsJc
ZnymyAvi9ny8QtXmrDMjNVx7y7yNiaAroM6ChlgN2bHLcln0DpzOLMzgLVfEZgv5
r9m2XzMAo27yKG3Vz0lLV/aizt715Vp9kbkOyrHXl179D0FRH4iI8hJAq8Dh/2fo
QcWhUU/2/c5sgktion8OqeYq8v8hLoNwQqPUKMW0yH4D9YDdtBmadm9xUxS+AAGL
YAopMlK/07IkQQOg8Qh3xwP5uJirqewy0iqy5SHaUPo+E+AmCQVCJ2QRUwwlRSoz
2QHiA0U0yHpbu9kB6kW/+Jz7fqmGtaYPM5MAQ2m7YB7ENdWZxX8NL4afAgYUhFVh
G70Aq5DjJ1nXJ6BHi6ZTtfzIBwJrwKe8Uez4Y87uCs/bxlN1C6me3yW2I42dkfTk
YW9teEq3xtcUtRgppfHKq7J2T7EMANdfYxWyV/cgUJz+Y9EyQ454ZqCzCBVV3/TZ
/fKgyIi4t9ZvObJQSIbLU3ZzGecoeo+eVS+95iGOwVaWPTxzHx1DQRKiBDCYizVr
w7ytGwfvk7lT6ryY+PKmsg6ZqeawO5zkcfA9XEFKRaA6LjmTQK8V5DALtH2bsFA4
YHCMZhx8OekaKSNGssUQZM5Ojqjvgdgp807Mgo+x/jTq9kriJ2t42cQGcab35NOo
noQd9llb/u6oD1Pbg5+310orxYtqLkogNQKZIdgZoJR/NUn6lnbqHK+0ChyL5oIO
oGaQuHXmvScrDvb0EqG0k+fvrvOYo+9eSzjNPh+GDwIxRdRWmYY+PB57JHoAR3YQ
6C0CwpWuKT075Mi0yHnFH492WqN949GcCAMnFytEE3qwxkOboQ5Qz96Ieq1Seppz
XhR6b5/PeoKa07nO2bQO9rohX1RwkkiSm3e00L2cHDHYjyxPXa0yGXCeI0nSU272
3mJ1THO/1BAzLX//zEEYaoNyYB/aO7nrb0pbAuXa5RKiheVLaunxv+lNGacoCWRG
QWfxS6T0XCqHsB01RUrZNLvP0AiFmkk7jdPgzGjYEW88DLWK+kmrH+3aHYIU+E9E
Tv/CWDoCiiARzYkR5NEQB4x16wX6hUnkJw1siJYtpkT55N5XRSMAfUcue29jRMqr
n/WzYi9RLgjzFVROAx+gU8/wt2MNGLVfpntGwLpzR1HpucTSyPK91gqPoBfi+Hgb
sK29gT0CVi47SUsHI1hYEoNGtrJuYZ8A/7r7QgQe3yyd/XIvSTrR/ZIro1avAlL0
O8wvsAlMkx/KzKRtL0YGqt+30OnfCEsv9LpU5HjHse9SUvDYGaGKAmwJRsRQyr7B
nDZueFnw82bdzHPVMHmvmq6MA/pv3uGPYwAuYedLnzvdFccbXMuMGAy7fIbw1FjQ
/PGXt8I3G8dphlcfw/AgPAFl3KJHAp8Il3qhB2fvYJFFwhBNKSLEsnEB2toxwlyB
Ys0oBZNmf4ohCrVJKFnmOi/c8vMqtYh85RgwuvvlVL+P2yo8adhBw/Upl6HsxN/S
DNka/G7FoGbCDmVX1njCTCP/S/8dPrNp/spKtuNYw9WLRs5OgZvby8jK1qhp5MeK
D6cDp/DEMXMLoIZC373ErcZm1iR7+hQYJc9MQyeQXWqnID4A6k6nn7Zx1eymkl0P
7U+cryCXy0vEbw7lA2A41t+HskI0W0iIlsFxFjSgDArt/S0z621YKiFiH26PgzIY
Tn3Abm1T7VgASIrtICeF+7hxN5eMX7/3xtp9ffMsQiarVRjyrlMSqG0n4d+H+EQO
RRDAeHmjm4n0+feKM03eAAy523K2P7NSiKGOcBUxFUVolra+sFylyFbknbEVdU2c
HwiHH7cTz8PsnoHhcK+/EnFLbCDPCr1FQnVvsZdnd1BiFp0IQCef8L4gS4frPQwy
UzXQImfinA0vU4MuXdoWwVYCmCCsvPfAMazx7p90fs3Vdq5AJiNN/4Mzsm4d1gSY
cH2HLiebOrWdQpKKm1vOh9rPO4KI7E8wrczHnc1KRNTq1QxD3I/ItUxkUf2ZSiYl
7Uyd01WkaBabMrIkjRWRkpuGm9OOZTifs48fDX4K+Tokl2EQXE+vcXij9uHgUyaR
qq+/WOE/UkGZW6WXF/vfClqqVfRB8MDg3YL03t2RSiCht1AeOV3P2K9fTc0kT9WF
302Zqsa/CD0M2dVUZE5+lKu3SsfbbUwRDnR6M6TZaEN7ZPs58OBCSuvR5z0YcKwc
3l7KLTQDVYGy4hD9+jTEnjqFv23uAM47+V1IvFz/a8Qyj5wqO1aZZ+jMIN8qGJXu
nwECaOcJ6g6xcYm0q/FPmt5ltnX07VlwQck8VmWdUvWYhYGxteFDUbanx5iRve/F
saWmdsxTGP3cH2rqO9jPeN495+HairYmyUc0CiAJVKMRupG3VOSisGmg4/eVgD7t
OmkUwsuIqBv91KwC4bNbesZ7vBKhYEWU/SmlCLRxMgry8rJ4N7Msvdh7zqqqBBhT
pAYobjbdbLGmq4sxCgvq0TqBjmcOe26w+rNqpVVFWLon/xxq62c0jz9XJi/O0Yf6
QmSzlmgdRsN1gLTjWvXpqpZX4u9hKm8gtUof6drp82LxHRRy24m7tSZneMTgStNb
mTRh8opcL245ta/Wm84ELgu0yRRXW38siTSjDwlHBFFvqU4Y5W7Znh11VE7URl6b
WJ5BXnjVH5jN1/noPRNT975n3I/mbdkjjPGuaKS8m1eWih7ym85CiemDmp3sbHfk
3JAd12NgNrnjB14DuSEQRKf5Qz+zl/NujjYiFEXAD0Kj6kZyqP782T67OSv+4dON
OPqAG1rj5E8J/H1ScieovF3BxXNV1u+/kftXDsLCp/liXaPih940qkFw6P5hsPr7
ilPJQzwPBXXCwrPNn5fImsEv8P9E+zBST01Ca0hM8GfNb86kSX4O9XVAQZVoyMXI
UlwKaL2HwiUAydbwTtYXn2GG1UEg/0tmbNTcKsZAPSiBSGZmqcYUnd3CyINfpFwk
C1Qa4o3T3T/yuuQqgTdxfonGkr9ZcAFv3lNXTur/1+NGNrtXD5+m3+A2dgW/N4Gn
XaWicu6B1A7CmdcM9AUCXpVxYgmE4W5iKevD2NOm7uqzerTh8ALoMtqutAo5RBie
ij8yBQEIhVrhYm1Jvt7QEZoNSy4EZQYpQ5R3fguiwVxtB/Md2ToXHKweY6tiN/bQ
L2U8cQiEta71K3CpoP0ZcQ5kjLNt/kxfOZUu3QUNmzVa0L65ud+PAkClxJ3/ZrJp
gga3YXupkeA4bnd1PmxXucDERoldeaHhlthAl+jxD22ymNdg+DXYndcx+EsvrCTK
ZTqAkD+Zz0qlm/JZ9195q0IoPorsrPPlx0x+GJC09t/IM7oZR+1b7LztFbM0qlMc
uVbi0nqxS61elZ7ZSqDcT9lRAyeoC46Cd8PfLn8fchiypqdI8y68WGlx1cE5HEru
90j53EnDyMmQzps8RJfVitOYF+9KFknb4cH7+9+DkVca+vkvsocRfyMRWewC9gHw
cMR85eVUr5233DiBOYYbiEG3gVkM8TIBYaAlT8/ssnpaetxM3JRFE8qRrot5fFd1
cBgadIw0hKGhT2alQmqlRKe41eyyWsD08Y6HNTY3YLfcFBjdHMswMsA87f+gX+wt
QsMMiSw2a685UKTHHgc/rzE1Feu31EMbUbgHn2ekbV9INBS6bBBiQ1RETH9OAYeW
wuB/1kqZWDgd+F+WOnbV0akOr08j0cddrz+4/nLuqujFxT2eqhjCzyKayAZ6aJxr
F8sKB7FPZtaGAWYNhlo4T8b0dwdC5TiSi/qzEe487HSXQb5X5xN1WOxwxUrudixP
olb+LPX5zyIYycKR6PGIf0Y3GuM43L1eSWNn2/y6EApp3K1lrEWwFrwZt8J2/qnG
lUnDfaSDAK5MEeWFvAvFjLginj5TV3rk1A9f2nzD92wugwOqbi83dsr9u4wupodc
Ml14LGQKFqfl5zmcg44KVYqiBxtuHEvp5aiwwZ4mzh8SuTUl9Jo/ZzyQXTQPCPqF
PdZxEf3qPY5Xn3aQdeVfP6/eN81eVkkD2onLm9zCuCqEpJSr89bAFw0SLuAC/Rfl
TkcB5SnlO0YV4RaD27E3aaAU1cm4Z9gbU7Nhfc0aTm2gDR+cuYZ1lH0RP4ZnG95f
D1zqCBJozozJa9IsZwFRwExHFBMP45UCKEMMeknbpUBwxdvbqj5Sy94/y9BO6rT0
MhOzK/wzRIbYLx9CU58FaU4zq7+uEz5nl3kW7n+gWhUonVs9iSY/JKYMNPasdlzV
U3N565j2fKfhrRMOmtRsoSqye2UgRa/BbaQ6fD09JA/D34Jp2bdCNb7X+QJaAn5W
tBsKRsZ5WVfWhQsqa+RIjj+q65S5qV5WFNoT3XVivDKRHv/DdqV/Wj3XYl9Fn//e
qoPnfaUMVUHYVwy6BoOKAD37UfiGyo9ug3pnR2XDb8ZVbb4rWP00jPEDshyxPJQ5
JViZ89BaabMEv2IAORQKyiwwVcfoWftDSNmZHClzhRBPPHTgaPW9wDjvfgmdmSgQ
VuybNc94ofIZT316Q0m2qW3Szwh3lAQYjCDsu+gbfFTi2k4ZxzYjRTYsL5n8I+1J
Re2Nx9LtKiXMEt2rkcq+5cYaew5OLkzrdkLfMKE7tqB0wUkPKdMYJCjN/YT3C0HM
hH3yb9LfwThDtwcqGUth1tv4Svj4Q3c19N3lj/ji5O/OJpbl8GIqKWSP+aH+aizX
c+vkdW3BL9giFQf/c3xFK0HfWaGkRMqifeEEqdvpqNmRfGMoozbcO75wP8Y/cSDC
XitSt6kqkfoNJtWncLJXpS/kXgUTbALch0WffhEMLPqSZLWpTRSpmHe5pxBY3AG3
P+d3gTXU9eo3YfZlsGbbs7GLZ4za9mRNSqecaBRWpQNjvoU8m9Q5xMMiudoTQK9o
otuOTnbCB1QQFzbqoIPiiI+p444X7LCKtmtflKnGODfY6qem97UFAqpSr9Xn4RzU
cWZR7o3ojnjQgZh9yEt4muHgpSrorP6Oy3VSemleU0OUJC6vVy7k0NCrQQll6XA/
MYNqgxaSwyHL/5wXJar4fcihDz+K1pEB0g/gP118g7TIU6Dme0L5PpqXveHnrMqI
be0LNL6OfCD4+9sLZTsOOgwyoDI5wgTVJjJVbwZEfTSsApKA2RUL+8R6mJlCwsxq
k8pav8UTIMHerB6f76jjf4g1lz50NObQV+Gsqp8Vo78Aw/TJOm5uKAQmeXh+VmtA
nitxNTquWElGvKCCDN48zKwEozFv0mDZ3DA9msAUWIzx12mYtKiMXRp5Fskyy4iY
E6HiwVrob22FEvNU+nKRF6factqvTdnrtGb28R03CcZ/PWQFwydnUJ+byQvzYKeH
7Op6zVY/VM6+XAwL0ld1h1jV/73YpLvi7jH+iuKCUDsQ6owzd06O/EBoctPze9BN
fWFLtO894K87Jlm94eHeng6KspD6QRAHvL9z8DbTN31lOSSWQqCqZNIO8DZyeuoE
rHY99+2pzid1WbkAwIBrHnhdsQjIaa6j5GbdPlIOG6+ZcRUWHrAHSHaK87riGY+/
o+2I1B7TGxC54/IdvtyEmkcVeS6AuDoBwIfdx3nvjrnbnK/u+gHeD0wTRaN5MmqX
gOtk47N5WBJqc1zR/r+mvYQD82DZpG2Pe9cTj+oQC/M9GYfIj50zxvZ3P0O6/PVY
V40ZIt6wlWlnplhfrsgM+rmYggjsVgCaUyYcM4bt5SRqtIfAzGMqnaG3x/hts687
n3vsQkpD/UaeDXzRkzxdptQHdINpP7pczd0lxRfynGi7dxv8yQqmmrcJL80neYM5
4+sj+Gs+WbgwIkM/6zsY07f/m8s0aFCg1h0ikHtspSWeaEGLhRNBDSpXEp0OEQpc
ir0TW8WBzz2G5RfO87R+JnPioxBYpoym88oTBDnole01PvSGAyg1yZJds0tWPUqZ
YO7MhZhfYb6viVZXJy+oVVL1XezVeH0RJJXCZ4q4mbKSBpmZnqPJKueuZGW934pA
Hokq/5XaKX+quYHXX23wEsDFDVC04rcmVWpmQ8g5IaaZ7Kk92fdhV4tXsOJD1bBy
A/P4Mey9F1M8pDXqCIm6mmXLQ8+5NIqpkZU9ZX2p2KAYjLzUpwZ/qSLW2Yx07uUs
uIEXz++516gAyzCIxDVIS4iv3SJDPxVdtxsLIswv1pH7PyltAwdqoPPUgExLPsDN
GseX1CcAEMzTKd9wzKHZShGNOEl64xhTB7n6cVBBfp/ItOfUFTd0BTFpo4lgw9VQ
yRnFp80m0NgCwKdQjn9TFlh09TY+B1AVeRyqT9CUVE7o3Emxzj4XQTdwuqmIou4X
qGvCC8481hZz5jyuszOQbeR6KZxgY8gvWFbax8o9rDkRqCo4zTrD3k55P4uRurVw
U+8+1v4mhOYs1hHdDTHTdCGJFAlPjLIIA5nJkHgCmcRs/wCN4ftg/gM1oMMdI6wU
CgIaNO1KJyKv4Q5mmTqr9BTnrRrXOubhvhf0HmmVagpCOSXwVEpqGjI4DzZVOa2Z
h4+2ksNgYwx68OOKFcsJ/HCnGBOPS9+T6JHxymPSBHTqW0Hqgwxoj4fIoxdyG6Ct
FboLhL3AgKl3DUbc9Cs9Bo/bhvpnBIRwWrJlSYrW1iVp34iRiJrQH8PrVKSYRhWw
NO44oNzQWpJmTKtf5PB43LxaZb8zFmwJr6Zug0LHO4Zf266rFWyzS+ILSAYIt+oe
ukxDhSYOL+yNBJmCZLaibh/+aDbPYxeeAVfF/hTNW75iRELm0v/f70v9f6K3NMcQ
7r5qkRXmOYXpr2fi4mRwCwQFkCgjyOfCs8M2CegYo5hD5M2GdDn3F4RcywMdUKJf
+Ya2oDQGkGtLE0IvSfFvtVsRUH6NoVJnMWDatBmyOJdY5nPyFcDEsZnIrZu7I7Ho
Nb2+X+5+Im/ADyDVHZKxGd5WsyiXmS7QasfP7b/EoxzkqU+BFBfKEOkXKaXJj4FL
RV7wMxg1xJqLGYbzWKmPKsiMxecYtXlYGgOv5ziDYHQ2jBWqZ9Cr4daHlqnRSmLe
M+JI14MYht0hhuSa1yl05yeveBInLsxJdasEPE8EErzqwSQXrSlHxvZDinsnOsNL
2PCozpSPg3s2v1QPZz7WVRtZO3CXwpCQYyGfv3Ofc0OtyjUEnmlsgpG3i+tiEFAj
F51CyljRXz9GZTcTQOx4oT/3wiHBY5mP3seTGPa74Q+Zd03Yx/CSG+mmGhm030k8
x6DxI3S3DAbUxnMqoiVMKCP+2FFV+2WDrNKMdygb8INtPBe40S87WE3f/8nPgkuw
gF21RIcSWEJlIJOliVJwJKmf19wT7NQslaPP+adyjVcOLYmFZExsDcByh0INJ1un
Zmzpq2Drg6fmsKbWimgN511g881smhK0LmQF9OM7X6mpQ1Zbz3UwceWlus4iQNA4
AtGAfsEqU4GNDlSCyAhzn1lYcj2vQJUzfid9A1hK2yZBF17HTXdsXjKZS9vi9DJJ
e49p25yD78ohcAuzGl84n8+ErdnIteVcN78uZ2T7g/0h5o0rsM0WftWRPUZ059LV
L9l2D9nEB8chz1Ob/nHla8PCF9uDmEMdnDCvDTXaViqRZQI7L4QMkJZT5+PYVXU5
EC6aMB/xHGD8UBG4YaLqqwA4DdIiZc0mk1bqLbLFRbo8z/fvgQVOo1eSjuScPMoY
b9rBFIo5uTyIWFLekcskEr3uJ4tFv6Eh3gEJ9tu6S+JMrmluluvFWO0ADDYRpo7T
JTka78pwA54NHA4Zymf0B6BNPblQkepWliuSqW4nx+0obXoEFaSa1fWGSflehn+F
ZnJMr3N/7g6TkS3Y6J6Xn5oDNwHm67uiXIWLzwtWrXiAc62SB0t8f2AvxAJm9ijf
9Nk2LUVva5825OUphaIAiI3N9j4wn103glTm923O1pq118hWpJ+B102PVKl6trsb
+EMVt1gNl2/Z3SQ3lWmpgzI2AixkwQmiOXEt8zjh2ySwSsZOUp4PWVvwisgcDI9X
+uWGlK/wBtZzQB6RZ9J+UD4pFMyAUIUwHPRTYpzzHby+QvYWtdInXHxYabP7h0AX
ulitG3Eexp4GVevgNAJBmepXlbWl4XZ+MLzS2ZPsSBTxoZoeT49la2ybtH7/eKGP
3iCjADDU5CqWHCYjPUAXO1qryH6Y6dBgFp4gQvFC1jMEJu1Dx/kus4Krd9mcWJI5
qqws45AiVM3awbFL5b6IoYboiDPOyGBXJv+aQExveIgcqzrgYsxmzAFH6Oo/9Ja4
FIZkVUuFei/+K2Hod7ntRGEa8ok22o+86HUG4YO6wO6fpZe4lRE5BITxN+x4o3VJ
FRpMeiGvFhVr6n6reB9RgAhA/rLPtbDB4Ng1FEUvWtPfRBL0NyRpSjZJdT7o6CSt
9thZcrlfyNTfE5WRFZ9fuKVmp5gSj4Ak35IB9GueF7XYH0GPKbyUhkf9cfNXGOn6
pVnNSs3pykgZ6pnxuV6YH5Zl9/2+OoT2zxvHs985FupCnLw8Nufi14QFzF3vW4lb
Dk9QTP/APbwowXNXd1VKqiHf21ax3yYxKQ1rNW6JrAiupoI8P/xh8bgu28TqR9Xx
tZmQ8/dn+PA7JJAOE2/y++VqZe0S+6h7+jN9j+lH0aY8+TNGyRiYvIV5KcQ8Dwra
hMVPx94/bc3lnyN+v3PAFduHI2CuovvZGLCzGhemXMqSwoSdjX/OaY2WvQeRqlZU
tzP/kyoq2SihFW9A9fOMQX53G1umnKPAxsLDDmHCo+qkahzc1ZcC8w+HoYTA0c5f
Y0eykmInvATw4LQjrCGORKBUO9oz6R3TDxzCoQl/KbGGMHnzrtMab4sh6sp8Idal
THr2Wx/1q9qoPk3fk35Ikw515El1sFqAXHgk4D3s+dNhdjdy1CTyMufL914HGeOz
wG5ynyTGlc9jq3os+QjV4qxrdGowR6/0zs2jk1cvug/aZm097y2e2vux1644KBxL
HAUx9Zezl1oNOxVROilYqV/X8Wkq0JrLufrJ51W6I/4XzCpR5XXKSAy9GdXmN9/y
EgGropdlAlG8ermTrYVkXGa4db2nKmQNmEEd9eLzh9K87GfeNB6rfVSw/K4+jeA+
pct/WVjMwLkL+tcMb6O8yRTX2KQ9XthO63KUlX/hKefFO6ewdrl8pfSKTc3k1fK1
sH4PeCTgGD2h0fqkh9atGVRWF4vxv668Im5DWoovO6Dzlzsjvrr5CxTly+bVrvQe
sxTs3Oyb/uT6YpGsCnDi1UGYoh9NKeVJqVxouLyOsCEQLlrIC8DP+I4U9U5RGA3r
pnDxHIdmyj9OTCP/xoSOMevYYXjirTlReKxk3eBto1r1PO3waY3ikaHCnfIK2zq1
HrvlVNApQ+kFbowUY1zC4GtoKCaLnrFuVygyY8mLyGY4Q/84ChlJ2oYye8BNco7F
4bVocKbODacof1iW0y28sLuPYV0LY8HBlDvf9efXPys4y/QnuWE2wAjnLzlWyXvw
01uGKyB9q9Vfl8GWKJgs0lpne7nBQ5YXAo70NW/WzTkUr6krUft3GFW2GCa/FuSa
0pp/TrAIfUh6Rg0fB1rtr+jCZvVaJ6LVmVo92iFNwq/DQIyV6/F6RjkV8rYawBjV
V8xeSUy6Ll+QGfnVVh3ykqazQ4orbNr/zYw0+8n+uKWeU/pmY8WnIfEtj50wd5sO
BU1mkqdIj/dYIzRVmgbnKVlaZKnznWDy6QDBoJ+nQGwmGi0pC+Kh4V3ItW7kG+kT
VcvYr36t2GSkvPqRjTk4UchIPGwOqlcJZzEjVBcFn9zEEB5RU+H8eavCVcu2F2A2
zIWrC95mHwqUASWM4h1xoDp2M0BsFu4uj2qZS48DNt6JPgTZDG0q2LuuggTlDNDz
3cOuG2ByrSXz/it2ANWsla1wHIzhOxRSheYPdkxawa70uWCcLeGH07RytvRzmbP+
dAKkeD5KMWJPicXCTk53gNpA8BY6g/wjpO2pzYTnX4mb5NmP72Iy+buB7cuo6d9t
ruZcIMJL5cpu5v+M/BAIvJuAJY6iUALRKNdj3P8G6eB3OV90JjT4KD99+6QPivNx
inkhe5pP5sTEzQD8UQk4htNzR/a7qqlXYJR+qrJyEW9zrOTWnYy+HwE+G9rykeIf
h6UyhrkkhazljtSu7nn1yJrgLmmcvf7Jpbv2BRwxX53xTIxmwPv5laz0pXl1FS2w
wUQZGdTflfurvmkLN2zR33YY+Qan6OJ4C48+dCuzaqoz1sQZ1lr/sts5JghC4l8Y
7yEChkB6aAcEiBnEnma0Mp+rLthA+nx3OrlDjhUafKln9vHaxuVZoTsXvUMZefLv
bBCA15j+dTCkd1jlf4j8p3m6Iq3r+5PiTLkF0dKxhxGltpL3QCVVmBAMAKZILpwM
zpDcfqriW9UCiavkDNY9mAaFeB7vdwLuuFiqJ+dHIZaaezKNn7ScCGZf/knXbcHJ
R68kShyT3or0N1mkkO6OGLyce0fJy3/ZfB5Coor1QaukrKFU5HbfZI9VvJ2m/gwd
5uCYKdIHl7bj8YWvg+IrOrTeUEU1HBgvHGlbE8bR++X0bj1kcRNdk9plen8kdYRB
RJGK6n25YtfgfyZK+fhKYMYEkMeFCTPCaw9f/5+mXBAyardPxWSgGbfRY+7+IvTy
HRJ8yQq4ZpU7e/bNXjWeFS1jANis73PQ4a+usRcw20ezHe/CjWDUf1RyrA2ThuJJ
HkrtKqTmpAneJk4Mft0U4b83ZYicqdBFK7rTxhHoSmw1+pvLNlpM4wuoCupMQwU/
MMYl1GxYWt9M7UegRXkjcWAuCR6ifn5eviBLyYPm+e437209TAfI5Djg1MZyg7Be
mp55ZgXGGw6prtxt+SuKqv67SycbLPluK99B9X5P6lYfz3Kd1er8jKaa7F9L/WC5
p0XpZseVogTnRI5rApXrg6igwomU/o2fPEDrggt0kWnlmP9wZ84sWIEiFH0VObjG
wwtNUiRBRghTaU4JkGXf42m3dlpZx77K/yTkkonHpPP9GjFFsI3LyRCmAfr4E66i
JfEEgWBIEtt6ld4KgLgxpKA5/SW5AkdLarKJ3Bq9f0bjCwVltUMGFL8ZFvbhlhd+
8KxSsBPBzWpil8wq1Qeme069CZXbRjE7EFUSW/8UZr4XrM3c9Qrzhe0wV5DbJg9r
uaZEaQb5gxdDoFzE2xxJlsvGKfiDiEqxnKLDfQWv4Ra7Z6aeMwZRFB4Ey+l69vT4
r9G3RGZiwz6MMVRtZPW5XrmBj/RLAagS4xJbNLAz812IjmQ5WwngUz2+YrCamWEg
sRju3QupBzr0KvjHCD4gD9WqnhnQnNTxIiKf4ab7R+wYTw9GLNOKEYMb5XfTTuTj
3szjeoOZdvqXz0qHL3yq8yyLwUtZqNPTBo3cALoYVP97ByGQVTZluhsU3bZzpSxJ
dfTqdxNOelCySNfeaNHBuIVi7E0YDxgH99YB9EXp4Z30YPHG71PlD06mzzToqb3U
3tDwI4X1SsyExmNv8a6KKR/Idi/YcAQE48feDBAZWYgXxPv9E4EsbSEgpsIgBPdH
8bbWA+a+f3qs9aJPBSvJHjix6iN/tO4vIH6QnN+nOtXdXdko7hT7aedeWBwAjoFI
TwHXwJJ51WgwYhvVAXQ4KKY8TFrcoGVk8nNfZu/bZh93qoHYDjXCfslCymFNYUKh
gG4muXF91IaY7TEz4H2X8hByL6qQt2S46fLVe/qNyoPJbc/LtIy4rGdsac7Przu7
yAZqQegKNun4AMJ5/liN/yq0JTeVzkKF9SHmX6pQbKgIPU4jY8bRwkn/svkhgYXv
YaKHjQ9Sk2+tPYQYpO2yrYTp6X5DrubmUk5IGaADEubVVU5o71bDVIxum3CjXsyR
8aORpI+3zlaGIpkvFoNLpVn3771STsoXzmaFTpDaqGRQE6V8vwLhfmWiIgYIO1Gd
RpPLY071YSG+o6uqJdchhXMZ+0BeguZ+6PwKIQ0fxdDkqvgiHnkrw41B98HDj2Wy
AmqG5CchWR8e7rs/FWjkXaXSOaC8frdLgYnDxqkKS9W036yFH5TiNf6OerrvGkBM
5bJ7K3LZPeeaHOJvG9OiN6u/tYEX5v/t71sceYnkKioxg5OrPJt21UZVAH0vjYMd
ZLlz7p7+HCp2jk42kJ86gnz7ROuzEzPAc4QIJAJJgp14Cf4TmZDhaW9HhPM3NJ/B
1e1dStdWRYeQLqnMNLQi087kAQoJGIlnGrWCcbU98zFE5YzUd1n5e/H2x2z01dVe
gLcF8x0+9KFv6pCQEYc55wflmiB7GZYpbuHVolFTiiUGPc9d0Y1dJr6/PZ4dwKuH
LO9K5ReC0uygL4cFqXJvXx0FgdNlq4Sz7ZmN6R55LQlqHvvD1K8IumDzedNWkQnd
y3udCgRzkeUIrdGzkG2eUmva1PMKutYNYGqLMcjDzbCn+SqpFr3IRmSPkAsw5sE2
i6S1MK8YkIXgMxMnt/DP0yrd7WQDkraAFTQCULiKPaBl3OM4XzX0iW0ZSGK9dU9O
LgVjt2magJ/4fX7NrecxQiIULHOjKJoYxVxknYIMBUKpMl56zEOMvqJNt6OK3ToA
fpyRlx6afEd3rPV25qr3bRl7lsz3KC6uDfelAQEcgJHWFR3YkHRz//uUdwl9VESO
9BIxhEnA8BBOva2Kc65Hc0NStzBq/YdAu80FFhKOrdiGVzhcQkd3evY02KvPbKXz
JCSLgu5K0IIk0+tE4yoC7NetUXWF2m2/NMI/8CGtmDMsWi3tHAbJeXbyY4mYnRul
m9vYVFGyecdwTQY3BpuHHnCbj+yKG+ULCoDqpohFxJyNqAqzseBnb6mdHeIlpggz
HKqiBnxEsZ9KL1UghHHVXUa9wFmR6IBOtZ2dNqR/FIjXWfBGGRQptCXNKiezrdJB
lrKsES8pagbbsxwUEsYIW3/mQB/HdlHhQcZYJNM2iPIQG5thNidJ3mJQOlfUsM6T
p/5ycP3uuR6bYBRIUvMemaUTP/WM1l3tDIxY498CXTOXkoypS4M8Rg2qnrThbYU3
Wq00nChVg4l6IN2kngPyTm/vcNIoNu9LwwUmoqi6QhQP4VQi7XE6q5eaJIWYWqV9
XTk9D7FRqS57DSgId5NPOiAlEH8pyUSyKDnrlQp066n7LnztsMsIa9D4h5Li2gfK
l51RbTOKMVazP7xVHRYdPBr2Vg1nVLBFkrGr5pwXm3UnaRwBacicUI0w9ajF6sdd
XP3o/M16mUZjwm19G+wLqw==
`protect END_PROTECTED
