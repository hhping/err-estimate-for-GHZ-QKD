`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rew1j4e8Ug+wpGaQjiZevgzr6tZV9xm2m02qoaZmQoJilv46xIgnDzd6ZCiz0+6c
swR0tTz0lSOrDWlK//JQtFzG05HR2l5LyLd+Z18yNkLMOy+7Wij7j8Jf/wJhG32Y
vkxog+xcIT0b+M5PoupX6HMp/HNIOvG+h6RayEWLzIG7YqtBuOvf7+QaNOpp2J6z
/EoweBEc0VEnAG7sUXsapxJeZwgXzYblH0GvIB10YjsOrLm33Pq4MCQ5NAv7khhH
xBzMo991gtCabQD7753L+VSKmas9iVq/VbB0K9M5aGatzHZPDUZPZ7EyiTA5y66R
Iu0ydJLaDIIs34prW9x+qyPEcHZ4EJ3SxeS/kkzCWF3T5eLrvutbUL+6s7e3JLR2
2fjzShY3neLwCHqYFz+I0TYZUxAAZgzy5L1k2McqgEL5xxgGE0gPosIP7ReEGHK/
AuC+qeHYQD2JWzRqtzk8btaO5u11pC9eqC2PTemi8SU9i0F2FgwqPZDMCpNtNBZu
IpMNEdBBlvIhnvt0xwaKkU8LRTrScBywBTYq1JIyvSQaPJRfRCzEjcpqrIIlPewk
tKipNgaMGs46+WUF+VVRUOkk3/oQq4PP9P9YXVcXNvN/JZLy8DWiFNQNn0OtruqI
HwL4ghWP/91IrkFPemh+2jud5m+qXFDIH/PnMpFK/e+5Ao6Vhrxk7cPtfwO4+HJC
4U4NmJb8+ZmKFwpbXKoNgaZQNPZPCx7z2ys1EzFv6uPExYLDdgSfOmb+daAtQP0z
+01WRf8DGl2HaefWf1TXdEzr0vwMVTo91/KO0uptbKPoWYm3Srm2C9u9aYIZE6nD
V43rWpQEHj0WF0GlhPXCB3O3U6XnPToWki4hqox+CxQdkRilnhQ6rYgDmfHLL5Cu
OZQmhy7mJ+5HAzFlP2VHhpB+y9ZJ1dBVe9G42ngKzOykYVDB03ePZwccIND133Bj
z82nTzlHDmcBtfeXtXWBvAtJHovyZMJZuo+9bUC0mdF6O+5VkrvFmSwNEI2UlklW
dEmCeTGIUi+R/JfuGNVOcx47inlkgc4ZKhnWSVDvMCLXxl/x81UkIZMXbK44Vs1h
EnPSWsRY5EkKE1iheCm81BowNxQzpINt/I7m+xm0wVK8B4q14yGv0HVhxRAtGxnT
dNX2Ecu2HDboS3ok/f+azJKRKQNL2sbI+/bXlzL+N5tyfBKXNVCaQxTdZ4cwXhpj
++k5ohV6WYxBPQ2389d9//J+2gYoN0Q2HpMry89KzgZgx0ZAxocnuMkbh3FO02tI
h/yyDbzgnoa9nr/KnLPM1DTmILIaBYJYxWNtjg/eJr8=
`protect END_PROTECTED
