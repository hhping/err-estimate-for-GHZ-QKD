`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FVl26niIrSMPI8Z81aixyPK8jBEn9oJyNkhuwQWYgeVT1OJXoa+9BQjLPsYZ3T+Y
1zTRCU3NN5GGR4JqU0DwFyDBvuJ2xqSzstx6UacpyhIHT/9Ww6YSz3FM3QW1NSgo
5jvXKkcZFznuHR7xU16mUlMszB//dfF/y6jHj6wVxy8EPu4rB4q9mSkYmTYG+Spu
kt51tQAy/LpA/VV8OEVzaMoMzapduKm+iuB410BpAckbQypz5CBmrLitLN/sxtwC
m8eQF2g+zTguTNm7nwXmotYEm72hhq0Ln0ArbVO7sf9IA4wn4S2ADtrtTgmVgeLC
ZWUhnusWL6Nr4PQGvhdpxBr0zhOJQiu9mhmiIp0XgcmLIKsLO1Ipgo5QxisFhUj+
9jpW6z2cTp5SnD7ducNikhKTPyBTtQppaMLxEsCCNVXDFcNJstCyptuqeey1Q4Bb
AoNwpb8xFe9D4ovAHe5A8cU4hFz6xYQU0QYz5OHQ/39oSfnhXZ8ToGSFtmBEa1rN
MHXDjmypTxcxoZAHGxgkZ7oQO0iyl66LeC98gZKInOHZBynyZ3EPpMBJFwSZGkxt
/aAK2/q31O2pk5K3scr/ij68l5NmOvlUbRjS63RZpgR6XMvuS2glWuje2sx/0l6Y
cnN6OaHruNHi6nEnWAtaH2cD0j53XPTZSna3AVkId8AVme8pAaEXh2GDgKM0k4vV
Kaux4Hwl0saI5sYcAAxAPwJtoB66yBGVGMxld9PZ16inb07FHacbfuUyyesscoV/
mH6+3J2SJcZrx9T1jnDPbyKM9/jphjV47bqJUVLLupj5aFR5VDhUq85L9LocttMK
NX9LMrLtGsSs9R+jSzfV82zhV0LVp551MJpXQSNZAzK2B4/cous3MoPMcbA0vBho
1pFdZSjZ0Min0Ru3qxceiE9gh6hLWw6yZmaJ95L5IRXTU9UR3XsxI1QQzZiwIMQ5
2CG1wyhj40XN02zdPrO3GLLvLPQqFtI+tCp6p9KFsTuzoUJsXaDc9s5drgdp3RuV
+7+RdQzFUZ8UbyR42XyjtSXbME7PLO9zNZqwtBprgV18N6OiZ/xmRPH4MfGmf7k6
rXi1FPXCLJsuq0z8w2QnjXMpfHW31qyJ1nGPZJ+v+HYh+qToGeS6/Xg2oejmJCva
oMgqeZcLjjJLtgMgulRYpfmv4Zaas1qIthF0/2qSPO2sqaf0JuQWnQb0fw7yf77y
VTvz0zgGqN2MFo9L5BDMOXCL63jueAvZ13yTz9bgNmf9TdcPdRhqsGU31nwDEN4j
fvQU38OkLWMXElUAxDxOkdpM8uF6dgIdCFw8Xy2Q4jhR0fa8s3oPIdpsKDFP/x3I
oX+xvU7f2SWT+P+bGdA/pCuFaIDBhinkeWbwlSz0RlX8JKUtC+hkoudlrqtQ6XW1
qQpan7btIGo65IDN60+UiTPcmSeEhS76XiLO4imlyIykaVTpD0viZ7yWt/vMEOZv
Xu/ONonIivdHiUoYISEkp9gQlutfQ5z7UlTi2kUJ1SWtbb2S6LFRY+f9eY9rDGXK
LR81NtRK2lWP4zxxHTIX5K99ZUynFw6C9pn9+9Q4QoqDo6e8j2gLT4KYSdxSzYVx
X0EpMYv7sFfAgpASUbO+vPMmfedSiQhVjPYUfrzLv7EvWzdlZbG6xHT/O2MiFY80
3Dalhcj/5oFLe4fyrhKoTQlngqLwa5BnUy8m4hpTBHSVzNLuSUGyAn4r70SlRB5U
yVaYdR1GN6pmu+OJI6UajS1DyNqDdrxPWEkCVR1TgX+KfDCFfimD+HU7vnZbLLka
rZ4NThcqjx5Y61BmLnpB2rPtH8nLEs5prLgD7ADCJ98ohpjfqWnJtUE6gkd2Aype
j7MYIhhhjiR8TI/butcha/8tt57BtXGaAKi8or3I6wBBOpiqaLtNXcqiuWQ2H3KF
cuZIjZwp2K5zarcYzjx2NzzXTZjqj40ooHb5/hlacnpsZzeFlZatAS1HFL6u3Tfb
8C93Hz1aFjVjTajw6r3w8yf0thoFB6wBXXhWgMgBqyo4Alvbq9Td47N+MKFfJZdD
T+rcSJoJ9V5REzc/RbD6mERk1XqUU101klI5wDLa80GzOWvKQeu1uJmWOA7qCZRQ
ZgLIsYm99DM9Z7m3UsGKKCQWMZf602FeVWYlbhB8ljBTmCjg8Q1KFhfXnujrtjxg
YICyfcRFPf48eZ8bqnP7QwXJMKr7BQ2P2ifJlK4QSNjoVliD8nqe1V4UvZQGoyVH
fUSF2aX9tHPyn0BQzFoBGb/9ERfy8CMsm8I6SFWIA0jNG9YJY0u8euZQOYDKPXiY
0Mo+I72jyGJ8O7l4IKLheqIhwEMZJExtqTUziCqmaYLFiU5M1NRuGnl7NUAa7CAq
Hi8Ix17JwGOk7PIOOFSB8uOeMWHi6gXZzJwfKDcRRfxKHINVupo3Ryw7q2mZuJU2
lX18kHHh/DdNfYjZQyPo1XBGV8LSqRE1y2Thv0IL/pUeIediUTk34MWMa6wv2dE3
r5jF/t7rBE1QkGkCgjKJj4H6970b7PnCNqIXHJvss47bKrWNxsNT+liNXm1aAYqq
0ywTsQ6cSthNGvdKt1dcg5Hev4osOP6Sksp84HO6cBamFHptJDJnr4XDaSaU2Cuz
NinmVtwRqWZ4qi7b6tFI2CRw5lnuMHkH4swwxHI36atewCGZsQ9s//ZhNl3Nx2vQ
qFar3uFFbjYgVJfLnh9IHyvDmSx8SrZt/pDZWOWsYjdNSt/SAGbvUVUngx3+dsqk
qNhgnqRARJwhhK9hBDBQxOkB08ZMpMtMQBesYXgjV+G/oCSK4Ikgebf0YPEKoZ/1
qtKtJ7w0nsv0SFx+VPTdHa8CUFRHEX35xPHLO5/nzEaoAYXjyENuVZkgvj+pEKhi
aru1PytLY8f4Afb/cGEcr9o11RDQkia0RoUYPbMk2FYHIr/7Zu7vm2Rp6jg+KIeZ
tWLXcU5fJDp+Nvt4BWehJXj1hHGy/zWnReYMMIsA28rhUrEJHdEZwL4YP3nksUAq
UTFIJR/mKivvhMv8+f4OlfHdXvRVPtLSZVQNMRVXRd3pii5VNyasG6DJAhh+eKPQ
WVKbZftAvoMhsXzIn956L22DLrAMAba1PF2UOqNk1qM=
`protect END_PROTECTED
