`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5gw5e2c0f4UZu0+JkELZYCvv44wvXscct/r9T6eJKzG95p0UcuABqtEOtaFO4wUi
MaWo7lyJ+ELYfOME3+tNs+4fl8IgFjrFTEE65/l7Apj9ibp2TGa0w9SUQGomBAH5
KHm1NL+HFlD/Jbdp0kj8qwdAYXOWo6BFOqhooYK2mpHi6FOoBzx5n63mjXuIAOgY
MNgBmobAG8B1U/fWzvhOdXp6mktwEoYEdFWKUugQtpam+2yqOHrRDlJEgkCyuYtM
n6rCpFHpXsaGg1OT0biY4ZUBbKjsUshmjfl2LbucOxfCG13MMCmYCWbd5TDiCViO
ufVUoecxsTbTmBGI9WPZgRSD+aP1BzHXpfHRQ6tuSnsTjwZ1wSSesXWsw0ZXHYEc
uQ9LJ+/4r3eMY4a4gvqNYrzll4q9+5Aoy5MZpZq9/pfA0eCJ9tiPzxyJYEncIQwz
3nWEfQ5BGDVpu6kacDri5xK70ozShfukeMsdpfMsb0F53xJVN5/uNIOJLi3y+KNi
7Bldr5kLZtSKzUkkuiDkGa33zxTCeRN4uG3lUXIxQZL3yZDR4zsu21zosJkGLtJa
kq7efvrZIDgbgq0j7Xfj7nyIsxiaGJysSEsdOQ9k4P7uICCsyASDp7rT/6D7wcFE
sbtcXReZdCvoqnmmq/8e0XLn5RxwJThJoGMJRJEirk8bHatEdXRW80IzCydwny7N
FQbK790x5UZflkaikbznohwOC2xWT4nZrfOhUmZGowRWq6n6nUzm3U+PilEjLxsQ
DjArMujA0gf8tqWdro6Nzw==
`protect END_PROTECTED
