`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ykGDTFEtyUIgFWythUtOgaOVQ48gWNj4WBEM1V7vfPSazr8V9Vi73HMOeRBwMdDQ
6RA4xR3HTaxfgJNEUUlvpcUNRVjaOTv7aDsRTjShE8s4/DRmdUgjV1hpIt6YWEAT
/WGrvKntxlMmF1gal6wax/Oy6MCNGH1XvTg/3vsYUwOSeY/KIcUBhX9UBB47nY8G
l9cnxMQ5WIrkiAkml51MW6LVksLI53KwZGs0ACd1Q45+7hObVXT031ZHc8+Va1Az
HIUUB9CEaSmEg4iNVsL9dzQ06ac3j4t9A71lWC1nU9JgSeWdDenYOCuxj45rlAN5
bRy35+a0uuZtYkJ+2nEx+CTG6iMj8QGIUyZa7snRmnOYyA0VszgtQZ173krGYwAv
zT30d7RFTPzUsCbIvARudakuNljgRa+Pz3la7kBC3qLa/TL5KbO48r0sYbwOKmn2
FfOxoyHi2KXC+CJPLrxrHCPBuXWIZLqILzHqwBDyTfVv9Co+1Rxohy6VHSZr0cHy
H9Mo4vTpR8l+gZmnuUqYPrbCaJUB1pjAVUtUeGXqbXeKGVOg6tl+o7+Avuaf434x
xzzVvTOZupf1peK/VJHKnTgAAMd69GwVtsnPHWXris1kttvDUzSivzi3vC0N4lyY
t0t4c79P5uY4caQsNSrsrfPl6a9gRBTGXEqHANYZC1E5iXNJqKfd2Tt+Q4iSMBdW
DOK7jyYjyc8+O1DE2MBqr22KeI5ObX5qowq1mSc/bVajK5rsRjDPLWo4O0ekArHe
ao7KER/Yb97FI2pLfN3vtY5K3PmiWUOEGWJwG0CO0/4ce800nQ2q2aBhk+nlA9mK
mjT4wg2psjpDGODeY35iC+krqBoxb8zoFfW/KBHnELZ2s5ue6cjk7THroVVJ0vlA
+mDZPtETmqlyrdQG3pI+kqPDx2HwDCcrTi4wsA0UDyJ8bHl1TEzTUJZXsy9aLg1T
G7vIjgx/fp+79wuAlBfwl4t81rr+kRyzj7WdBUOZ8G9r+sBqJszOmbWkU+l8QZ8W
h3EFoR6MisGeKM/mfL2dZwdd2bI2k3jjfURU8aL30YqCGfjlM4VuURO2EP9KkGzu
P35mplze8iAaR4QxNY17Le3KODjQ1fFefXbHXG8IcQoijJBqnwNfIBfwFMUH+b3c
HAMv0ABiApe5IQCx6QJOwPSBCvOODJChUIZ/Vckj64HDrSyecRPzKo4bPkthGXOH
L6l3XYdCoJZ+XUUMFyYqc6U+S2PRKQB3bvWFk293aeRp7P5RlpaLnS1TCrDuRyWA
DI3hLFesNs3oZTkzGq+za7Gpf+Ml4+dmF++tJifA/ovjUlCkfSjYYJklqJH/KEZI
FTgkrseE+iB02v0kWEGhLFtEpFAcFRmCNQV5Zv1aW5OHJlHB/rTBaXlQP52yBklR
g+RbqJcDTaW8qHiHs5sgO4tI62kK+1t2XeCEuiKYjWtoyKIyxiPSPa6LEBaziamC
gI7C++59OdPBGfrZaMwN7rkJqb1UCVlR1uSyqhlRgRruKr1nbApYqDDqtdO8Jy5R
Va6ezgaFqwbBJXltYgqARCbFKRBD+XYAn8e5TkE9BZUljK254hVMmlObHfbZx3IK
42EOmUcrpsn6pkGbA14KcL4IeaZ8h2LJMOhj0UYIW2H+RWBUVQx/ZW3bLxq7PtpB
6iVSVe1+8OyDgnnROpLDE2lew+Qy/qWKqXFUTR1ZYMI=
`protect END_PROTECTED
