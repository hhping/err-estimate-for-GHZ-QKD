`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JmWbfQilJplryeV1v4otaoie615m7yeLDSO0VSPF1hCJL7ZZqNNwA4f4pNlvpoWr
eSRstuMqN5UHPmJ4kmMTjIVvkAeWnlBq2LRZpgLYurfeZ+pfujInS3YG2Uu9mWtk
t37zLyT8PsCQRsstQxZfNW/SyOL+6ufWaqwmysZ7Mvu1YryoaLnZVCnLgKH65g06
M21xjrYFydRDQy3XfG4GDShDKcVhu1aD75mYICUi4G7jwp9c5ZmqI9IOVynM92NL
y/SMV1Ai6MNAT4kSTAbSt8t2k7tu3GPVUEpliTQcFuYv4j+G5/MCgDgDM0ZypERd
7ZR+QIDJahbCPOKkcUMotalsG9f9mbA9g0brn46/mu5DbnQTDZVakfzOfs2VedFP
hc9ZLn6fMnu/2BDP6CmwbJaq2CNKgqW8/6mnRcMSfpvGhiv8JLtikrTEyIasUjVe
vkBwesOC2NA/BulomRMy3rUap9VIYUHRSLJgQVymx/dPnZtA7bm6WXddP2yyIciR
YaoysPyXlS74kcmGeowYEwBpvJP/8jOaudn9OLj2wJHJ0jrdXNMqmOFRfauRA33b
pUhaiJF0S/B5TWCjhz70r4wx10fN5ujHnObql5LfNV21awI3NbdiiRxrugzFlmIp
Zre6JQ1gK5dwWjsfe7Enb8O//Hzin7fmtA/EUuBZL9VlVo/clujUJQ1zwrv2sy0V
NpNuucX/bq+kovzLititTqi4rW74j7Q5ZLzL+MLo9vK7JFaE5RgywGpatLAuabjK
a9dmr43T54ubLqaDcik9yn2rG6/Y/FTdRdpikwcWIAG4wWamUSwmAO8MyJ8BRRfz
nLXloSYGxGNXYA15RZ1vm2heCqCELvOQopvWvGUaIAnX6zSSekkvVonseu7xcrr1
pSmUGN9QbPFjiBo/ifkLhj8g051pn0kBXVLsYfpPjhrz1gYJFPZ8yFMnSno6x+Ag
1stX/c2xcmD/Kyw7m4Q4qd2+Up4Ddxqh0sbPIcu6I5PoQKtrkyqR3/gmN98yQjxi
9zW8KaL0aiZ+BONFB+kiJ/EzFha+x0+pcgh9lMReB5Ek2mTpwv2WtDIXxJi18uTz
DUMzUvN+TiF0tYIXLySZFa1zL3Rrm+5VE/Jr7BvDo/VzElubQ4Q4yhTCgCUdtdB0
QbMs4FaUDxuxHHw6qCqtTTBAZc5BP//YWQ5kTiJs2COwWDL+3HOKuAuvWbig+UhX
i0UT+7sO9UoTttkmacNupwfeOw9DoYOayIl5uUli+TuyG33mxR4fT2Md6Hx+zwCI
BgNMMeI9lKeyTDUzmYyQD8Q8d2LEtCYamiWzEik+4O0sP9w6r3jaJnJTiE/8Q3+t
dOb6vyYVR5Yvcvd7PW7cE3XgwRGUrEL0b2zhnYAATMNkbYClxMvDAn/MRnI+AVrw
Gr6HhjnTQY8RXGGyvgas1cZ505iC84XShucD21hTPVPz2vy99pJPYOvktFK0zAnY
cc14EpXxqTAzwIsaLzWvtsHHEzK/N+a6fTQhvUB/MvDIGQbwF8FsiqPhM6iyCfFY
9UFrRH6CIhoSKw07NrLYXB+LCjkPrKPZnoun0KTjeQygaKJlKRzX/CXvKxhhOIN2
I3q1h3R7fjkbL/ttogZR+6WJHwnqPT9lg3MUc/UeMahKgSUAqXrmmlJh+H+kNxN8
bS1a++6TzjTKCohhW0tOA8UiwdGZiShIRU5stQLaIT14snaWxx5TBpRa4VgNR2+V
f6csTpA16NoZGDuerywHup+yP0243FSF7jNKNT7xrrCfVJCGQlsS8kLQfm33XGPb
LDwbZ4NtoNkPr9uF+FcByKmE0gRMHRQd7NB+TmYtwpEcbdWcJdcQVFYcjsiAECNg
d4svfpRZ0Zf5ze5jbme0dODDxcR6j2HW5L4B6eXf11JaMa622dBHqES5Njq8XQng
H/Ll4h3jG9kyVTpy36111cttEW3aAD+CSgRLenuucde0P7yTHSb+HGd8+ARjSAsz
yMA1ZAPmY335QGH10jFLtTzs4iASD/TsWqJ+yUPv2AypqWATuOPhLd8FNg2RMkIp
fLiFhqjFlKdmA++P7v7VvpqStdUtu9PnfA26tzs9Z6xl6T3hKtrIuSi3t2NsU9+n
XWWbPk5ATfj8yXbOHtputUNzzBpW4MW2BSiQy8XRV4OKUpkYd2Y6Y5gAz0l+cfm3
zvD/K81UGn898T+R6nzfj4q8l4K1A21Q/AGFD8Ba0tNFa6Z6tgyAXUQhhf+bSBn9
MWJoy8atkhBf+g44Nmm72ybRaOLyHFsJ495UX9tOayufKI80ZMkJlJoOtJlxw2gs
OgMvKulEf1ZZj1oyJmiYHX3Z23XnK41ZVoEe8A5XJ+pglTSycTsVHFv66V0jeHAm
j+IBPVU8yGpqJKGnrk8ZP2Ofp5w0n7aeFUAkCXV8c9nXyA9K3WPWHlCOGJ60BD7e
me9EU7JANH1SzQSV5q1zke1U5Cl7Tllag3LCFfSd+57/yudq3d/4zbDn+h1PKkPs
c6fuu4SKAMNA8jF03EFIk4F1mg2PY6jH8MTLzjBEjtTKcNbDRA5xpx4y8p0HON2Q
I9nLx6ZNkVrOZHnYpEnVqTxp6LarFYNH/7syL6lNpYNZdIDTjEnAtP8duO3g+u16
h1Wlfo1c3zCi9C3c1NmfCMwuRadvcydFiOWMdlWv9N+ztCkpM9VKTFd7y78GqVQZ
ttRfYNRXijCUI+rE40J9RA==
`protect END_PROTECTED
