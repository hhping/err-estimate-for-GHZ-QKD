`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lrAp7USCmKOAa9R3b8zksGd4EuJvNHvOe7Zb2F9A/ECMiuEl3Zvxu9RqL0SFF87I
EBmXCev4OM3yRJceBWGrkg13GqF9D0KzQ4NHpUee28BLtdvbPszOC0sipPTFhhvP
ozInVfObZJmTlScxD5Kb8QRVmX+VX4sKWrBYDn3MOdc1+TsA4D0FILS3L3bRwuk+
kHqFwVqtSwEFFg9ZUbOByVOyHx1kQWgZoWmAA6PFUGfe6y0rvCFdK3DgdYdXPp86
CHuETshL3d0sg9EU6mFDXBokcrK9xeUdBg36vw6BcQajx1RL5UOXmmgh58efa/Q0
yfdZedowNGkrxvnnDhnGfKAxMR58Dzua607mhUcRlNa0DGxNNE06Dzr29FGZKoFK
hOGkce+RNumxdpU6mI1a/rWayiLIdoeYj0BdL0i18LUm4Yoo32yITRxQ+blfjZzX
trnm9KQ8hnOIHhTMoW6uWCyy//EgMObmpc7tU0YrxIP+PN5IJHYVr0aQp3Nrr88t
R0MwZVcyRTTO/fGyxHR4YvkyAxQeqU3vy3v3hhoeuSTWDvqR4bGV6u1Ec3UBbmdt
ELwNjvHkdlICtZwo+Js3wD3lJdas1S1kqAqiQ7YfvEAb0l579yI9xh+miX32FIbC
ZyaBi6t0hOzNaEidJkkuJgGldDNGXDlRHP04cAJNYR33xqVV0Rp632YqBf+Pmju+
uAU/OF8sI63yc+Tx+9qZ310kddoX6Hby/3nnZJB7k442mztC0TpQTNrfQDc8YjNF
hYSBuTF3dw0ntYwkR8E8ekwSVjAb4fVxkhHbc4IaUmsiCNwU5iu+Ryf0j7OnljWV
t/NMz9XXuGFAnBIVywtabYF92mPwc19IA1Y5VxAvT8hLZXz2zAsEp5PwkSXzzBl8
GXYH/WlqGtmWup5x/TZln+ALfn1xlRmh9B5xtoh7XcNbig0brFbLMZ5aDtXmRzrP
zMFL84AhetG4hkxb8nYmqFhAQ8hZ293LsPEXykVrgn06NAydeBMgrPingddnNOXZ
Y+GBoS/GP2aGfw3A4oSGc/zge86+xWaN+zZ/zlWEtUtufB52+oI5G0kD4XXO0K16
mErBhy/nCO1fEhcI9Wdk4ElCr5mOc0GFdvkL5v/b69tGpZRt4VeHvdOp6xADipYh
e4SExKOzY/4dBOBXlhpT/Hau2P9cXhKH2LYWvxUpmi+GO0Z6AYcUp2s4DWpD4TE7
2lVJwz5BBuNXja+Oi9rnp5a+W2Bm0zXNEj5nKUhbmZquz5yLXO4/Gf7MGcLKmEpB
sj1/d9uDCCDfdjXUkWjI85yTp08oj9gaajt9LdhgWfApB+E7iSq032SgRHS0Aa6d
pbbJNJAzmTi/ikEdVgI6Z5ex3ewQYq0aBk6QnBD2ReinxiEXt/nwYGzjZQiqsseD
e+gJtZJRraOknEE7dPOFk4Z39qSLc7TZyOBMPCo6PwMoPxVpk4p3jWVZI0+IjFT+
Xqp8cY1oh10Vt4YTeWvUaub1sy1Bg+Yr30t0Mlh6nR0ZjdM8kTr1DgQ08ejjEH3n
7lEErygC2rn0PiPKK6gD9/aEUzoxRDdeuHdQGZTl+xLkl8+4FZEtHDnQ42Wlb15+
SN1TMgrMmM1lO050OxtETOTTXwtDGxX9p4OZFc5n8EaHFmn2RJBlKDh+4akfNua7
UUsIuUdWLlbma3DdcNRK0Q2XupDD+FiOO4kLsKECJMprjmdrTTF9+RLq39SvzH3X
2FiaKVJ8rZ/1diJ+aX1OCDHIJg8bzKCMG5C+ii/vxbpey5+pMdfyxKKEvd+5WUaq
oQ7/lMPhoGRz3Zndlo7EbhiB5HT6Ysp/xFheTlazPmJqpuRPUANqIAShTZC2cidl
1p+qbXmkZl7XIUfRwfvrgPMHGHk4A1x6UWYlo6KLNQkDXn8jOsbgoE+Kj3dInMjB
4ru7KXZMDw6GKZ7jhZq/erdYRa9XuT4yvGfXRnYIUgXvfoy6Y7cLv0u2yUk7pIMP
u/UhghkeUSpm608cp3UEIVlULF3ANv2KZCoQ9kUd9X9e9MEjvONtOi3KnVlls7oM
01Us68Yx1BqRZg2H/hYjwkz+7dKkUbLOErO2+IqqHM2KZO2UCWvFYlMpRRsES0Ws
xsoUdVXy5BkwkyQD7/PBvHpUaqMH9ffrpIuIJEd3fZiU3/6DtWESlTeuCtkC3B7H
AcKHj2LVJ9RvQhUET+Ec51Xtt9+L1u7IyNiT3cD7sAUu35GeOijmd0ixzrAWtNt2
1+GIDM3cjhdaFWdrG5O1vlDBUvQX/At4jaWIAtdFuKioflUL39RHhoKjkxnrrpiM
kCDz+9YSmMvqM+1yRYWDdc2L0iPD4gI6ssSjprSvu5BhcXZOrpuEq4GLnmKjYNZL
otkFsp11pGcccAOaqzvwfVhu6zPTjL9wXqTzpN21scBRxWKJjuCilEVnYd7annMV
36vmX2XNCAmUgInB5JDX+fzuhfr2nTcwPMGkHvoz8+FbRP1cS4uoEVypmJHkUhND
QN+I7h6XOpyYKuHzL0RNzGSsbucbxufNQnbSHau1Z99lmRM6OD6wNuy8Tqk8ACev
iTFsfHTnqTBdo5LJ27dWsY4loi42Uie4tzMoosLqjAqPwQ9H26SAOoopCniiig9m
3kLtQrFIcJrxfdB3EL9c1VtRkbppe1A+JX5qyTbGpuK+10ZZ5L5HD+Ea+rsgk4t0
reZlXI/qU6LaAIZHHBiSkwDaw1ruoUUTjqM6CqjJOcjj92PLso7UIbobekLD7Hrj
Y1Wn/R8YG5ftiQB0ZPiamPZTX0DkJqidUESokuRhJ22BqRmEeoYzQ2bVMDj8Ew5n
5/HQbM47dK1ym2XORIHy6a+J4Pl2DWxNihsprvw0nKQDlBqtfE6mdNtixS4cpZX3
w4dTC9CmBLRcLKb/hTOjY0G/Cvwkqw44oVIf9SdhoTwNQZtUYW6Kj4d401RXd52t
kjK6Y4J8DyGjWkBpE9Sy2otrioeAwL0VL0FKyw+qnKCjKG1lgL+ToonOdJpn4wiS
0meZg0c/yeueAPuOsZzlKmFe1wiR+vDnHWC85x8b58LhnC9a++Gp2i/7XeXg4lal
baH4EdO6xYRJ0kKoCAjtkcRhO8X2eUfJmQC/FCxZ8MADBCgYK6kHH3D7dogM2sas
BvgnGZa9z0q9n8fmcJ9fXb+UEf2ykG/Ife8yx9n2ncTeQ4qbdN42y+fT/A3AN+lY
3sFBJ3ojREEcJjFglaWGKYqtcFRDArpvuGBSZGHyRngE4en+uzqXiTbut0WB1Tx+
QKC56wrnc8kIQyrefzbnKpQSixj1r9wdLn+tDRGcIbn6BvKtG/HrRANA0W0ngcry
tzGQhRwVgcwAHJcrejj8xzQyOZYJx138iOEvga/P1ZHbGaBfp0N5VDAfrQXG8S9m
7jb/pYiMmQWNx/C+DvGVZ7b8xU7jXTplOC5P9uIUMOHhwL8N4iM5BMoA5v1DUGQ9
ZsYbg75gZ1O5Mm4O/iUhPbUfYaDIHoMWSRSYKN4F/KABKCEOGA4+McKVnQCXOh+x
D+E7QxWZFYXij8a/Xh2IV0Te6zzfY14JqI8oWQdAiMPlvJfvqJlCifN1cwrAmESc
BCSg9K0Kw6NtmXJMv0WT3CnK+z/fFAMvcy6xv2SK+TW2u8QsoHwv5NMu48pJBiz7
nXHaffPBlEEzDAgtCVXoXXb25/uCSYAX06s27Nrr3GbPqePIxbyRFWch+1q8XEkh
My/BKZursGGX8VY9nZyElH8fgZZhKGb+nITtX+0AW9abFDjPaGQ9uKXAQJHLkNd5
rJKo+ZMsqlJXdf+3Of97NE/H4wknlBhRq/mJFHzNjtMT3NIP+e2qs7Lnv5bzRHnR
8Zs0mPgujw4VFf8U2iMsfELZ2SjVM42LT6lmvCu9P1+PlgoG8gvIiR2ytmWPiX91
RxB719LvVk9JBQ/iLm+lttpdeMMOO6mltAMmrrhY6C5OUsSvC07Rf0+7C6F0NH3g
fC5pUJWC3L7t0SR5Ick2QunviW8ZjAN8HqPUVzByJq1p7NdG2xvNiWlF4PoE6y3W
Qy2AWL7EeiRglvhpgeACIL98Dk5VOMXc1y6yTxBkbdy0lwUs/Rit0D96ZX2oQhXx
YadsAfLxozbx1S0khJWlVE4GEu1iZTWDA4eByYcnmDVH6Vwo7zAcXz0Y1Iy9Qp2y
H+uHAoMLfksYLcYFW1zWIBw0/AGfkG8U+uwncBT1Iqf7XetAg7bhemuf8Q/Vahm6
SDORQsQHPTHwxFVseflAoc2XGyhHbo88V3lycqK2Dhvbp7uzaX9ON/YqGV6n5fDn
f8hwMLr2JEzSrtzIosSQl4YaueYbK9+t6JvgvFkXO0776820YcM+2FFfL89L7UUR
H8MshkmbD4uZBfsdGAvWQAxyasvnWzr2bU+PPDcPZCUQXDCzQi0n1c8DmW3HKW9C
ygx62SSNaHt3e0tjfB1mREhWkmhunFao3GZA2+U++povQMiEZJcn6WpybdNDBHkK
A9+L5k+YCuE11rsCZ63W9aSEKBtlMChnDLKoNNu3K9+xQ3ioKN6AT4wZfQz2OAlB
zEd6ZhCDvm2b3SpJj2wNNJZNvfWeHCLM2gtr+6vz/pWGBAWBNH6PsgTxsZQd+jTQ
0Binf3J9ioGjMu5l8IFus2jzYGENFRdPqKGhReMLqq94qHImP2KVWBIZPnIiIp3s
FufZCQ7gEqvo0zQ/7XCJiWxs9oI2WKE2ScjVKY+tjQHSO7QgjW4C3QiBox7ieF/y
H2/4GNbC6hrii7ZhnhPUQb28kbqk5qPS49kYzJqP46LKvH2+CS6VrvF7z/mndHPE
WrV8Y2Rp6JIKXwNgANlyqLjSUhq54pnGQ6BvTSYkUgS8chsdUEgAXyUZTqVgdoOx
+CtMfToYrq48efZU/33HnHC+ymZ2gA63aS7wwhWCfJyXJ2+nqNKboD2mx7iIWg8p
oZM8vrso+hvF7zNhKIW3bH8beN0OTUI5yb6a1CNgOVncvjLcobQTo0W4gl+wfxGj
hj5d0lZpHDG+AQ+FfzUDxLyFGiaixZxJU1XzOQ7PHHeKW6zcSAeKEMXQmBRbyvR0
fsODenW+oYKIgdhkvL/7PbbKronYjJEJ/eHPQN5x6+/xuxf6dCa+yyUxNb78gktD
ya9H7K8oaJcnZukJZ0wECp7b+nG/sR+uihDXMWPHHsVJJZe36Gchmdu0urvOMmgB
5HuWaEILdvsFWsMCeXCHVqhhxDP3/iO/V5P1zL/sbdWCOEeASNjTm3doMgus7SjW
NgHaIUSpuLb3XXewi9CMrWjQcaXoqgqgzIFdH8FF+0Oj0klycFRl0YyU78Sa1EhF
gj3lJI1wWXxIQOz1b4MyNxVI+TugDU2KikRgf9vUsZ6KEs6r6KC6gJPousE3kESv
BZLrQQd++0Pa1tcy/S4lvxyiuXqXKYMDQxf9jcaTKLuUYzrwbLz9HgCCnSTg7/1r
frm11uEPtslN0gpNqQCWvjcfqODcQ3bDltWEv5wL5nzFgir8el6p5adwTs8L09Lf
lyLQPLtYwH0CIpyJWuvXz4Hw/Rp9R2VwHznNflckmI07fgyTxS9lUQMIbELLm5T+
dJq1tXh6+CODC50B3COhihFTgdIWrRibaT3WOvw7JmikKq4GFej1QupjA2mO6qVP
C3U4/Rk0g0MqdVmSoAQAX0ptf8tCrAuZs04fxUhKYN3DFmGmqmB86o9Dkt6cjoAE
gKoyhG+IgX5t98oi9Do+p4kKWwwqb0EAwio5Kzi3Jh+9/N6GGgLdJtPiVNW667nL
2TzoUP+oadVtNF8Cdvbfn236DSg7V6UW7AtCiS5/cALiscu+cCpbN96wW/eN1rp/
FqKsvgZ/4R3GgOXcWG3h4fKouyfcFsdSkjSsU6mtF2KS5GdtQ73mRMrWmiLkh78x
hMEnDavtc/09aKN697pHj08p+KcVGT+L5thWHVfRQMkq4rhRNKc01dV+w4mMEtnj
l75XJl0GPsjTqUZO0NMynYVlNZK4WlMzNhYOiMkf6T5VDznm9ggQMiTFeyWVoiQ8
TymjCcLy258d9CY35xCSHSOU7yj5M7zekKo5QNFV0O+4f57ibGslYS3W6i32RnX9
YHzQLv9tXKEHCDELAhEtncx7qMI0jZFn+ujwJTMhy4jta0ddU/uf9ll9MeCDv08u
rAHMQI3FuwmEKUIr3FTrBrmXbJ7B0LrZzpDmkhnRa78BG8D3jhbJ8S8uePNuPe4N
8XEhRDWz4qppuOV7sqLXyWnZtyc0AyUD6JQMvwy0gNbix9J+nGbiHs6Nzn+RAErR
O2vRfe4dGsv8UBM8rj7Uh3oET+kwEaCWFPiW7LdMXUBP712F9XdWKnTcgZ54qR8L
qHuAW8mcmNcqjH4ub90dFRk8AmvAW+w9LTwYYTjq4QhQ5zPuMNCd+8jmf6R2NV39
1qbzsQPBxtSCmtNcfp3YP+E2LSjhE+S2IN4qFKoSxKx87E2QYH1hB4fsmwjZFqYU
raoizdmUAl0/x6JluSUBunky/55BvL5Vrz/8dAj2lKQkpwj+vARH7V401Ix/wPkW
z+2etraslpCCTpLMdRHduJKuVttiZxF5G17kq7/8qcT3h7tP7IKebeygb/PH+Y43
roEhKai26r2igDAe/if+Owg1T9jsOwCha2aWebMqGwpyicE9lVWPjeXSdWXTEg26
p3X6DJPz4F1sFaSnEe5C2S24Fszix1L0F6wIKS4Qee2cNylnHOnY+wsxb0mNVmoa
v078+IeQDHvDE+64DdXY6MLkwVev4RLSr3MXeH73iK9OaYsKvQqCpnylhUvBQDbf
l7xb0ugXEfNvgXwA+Aj8L+Pa6vNbCIl1liunuizVWcbD7E391HzHDKnvDRV8++Yj
3tN+Vx060Iw3mjFDDdQ4Bowm/KZN6WhoFluSCXoc7ksXveMgqeJdw5rWIAzt0nNa
oH+lHR+fNHlwQgdS7NGB7ICy9Qq6k/uU+3HATtJt62wAnLjIHuNG0qsza0CTMT/o
VYloUh45YXf/vwknuhmbmpGeYtGWwk54//SYc6NtyvNsJ6Qv4CA/ypvj1NTZxRFa
Y2RdgFGW7sCydQJ43+2xR6MnFFbW4OzbZcH0XYAnRlhT9A/kJD+pFFCkOGa9JyHy
OHdCQ6YyBr0LxaYFvFaQ3tW9DgEOOPyd21h3W/7wI6hVLTC15fsWCQh41tORIbDq
Fl7zbQqJlBLFKSGnvotxzoh1zDj+rh8iqkuQ76KWPbSRfzoGYuo7+axjpQ2CAWtL
SMhDUXwwA286kQO6eaTwlmbD0UpwBfKowSrpN1oYbNZ6L/2t7OqaWs7sL1sa6LGI
sDr1PWL1EdgBp0WDOdFIuuXpQLTdnKTMkACeux50BS8dRLPtPLFmekueec4sf00V
qJjeZM74UFr0famNch4NayO4KZZ33dJp6K94hFPoXtjqz+6qZcusxDMuyr/bFPDF
GlME7EthKTIvsVNJ3dSicoqivNy+axmnEVh81Nw5oFNyTCBKC7pSsPDOXYO/z80R
qjcuRsi587i70Pk5KQ/o6eGsCYqOVHKGXPJ/Rh9dqVvfVXLq9JOUWRQCb248mQGc
/BKAJYpuSZdbmMLphd7vt8plO4QuwRRAqK8WoANrunWfM8kpxuDfdKhaUcS85QeT
15hrzwXWq27ZenmGifJb/0kkrEQjtPJd4QhxQicSrsZhC3xd74C3vfTQ6oB14ZVI
y1vuIHgGGOa5n7PXNBGiwHf6hM1HQkHYTs/9rRvD0Qq+NHYkqWhlVKrk8IZ7p5ch
yki4MvNWXThbm7pXttLQ/tvxE4vKLcIbJ8/6wpn0BH6zcvHCansw5dpgWKlyzjMC
N6wnJ8H8TV0EYq3q/fqbV6RnXhqpq+s1lhDev8ycO6aeIb7Vw4hhYPii2rIYXPsE
fqynRLWfN2G99ohPY5FGZjsbkk3wza1Dt/RqxGGN6JozQ96eQ/dJ1uZ7Lzw5OiM3
DMVXr7xnQ3Y/mqH6+xUYz9RSoRWyvZSOeQqp5OGsvcyX3o+vDqI4uptJISF4rzr9
ZKRq5TbMvFu/ZxrcDVuvXTl4Go34NbteIQl/oCOhYRBXU2k938QMjRQ72KdN7S3P
RhvJMnN6AsfFs/fSJ+WuYjr85a0mFiqgPrebaD0n+l2CE8BvXCG7kG9v4bgUrZtU
jY4ODu2FiKiFOdgkPiZ1w5MD5fxmNARq3++n8w5+a5HgIY5NXiBQ9Y2JGLIlYTbz
o7OjtzBqZ83o7doyg35+7Hja6yg7A7jWKjWqHP/mweBT3MZ9o1RSL/rI7kuTTVUt
gjXlYT5FzoiZqJX+9aYPsybldyrPFaev0GWzlhrn55g5WIHC0Y3UpuV1pCiZrZ9a
wphzGG9bJQRHPlfiEvkc04sxYdmcQPT0zijVlGkWPUcV4oT8nDcQ2kX3H0O4AM2U
AaGHRMx0KaMTGfqKjgt8L0Qe0cA3VQoG7kBsCq7XU/efrnDtBKXwlSbjh7u4Sm9Q
DCszQscjgDB13LAUJyTOcRQ0lB8PK16eTDA0zIM5F/Y7DM7cNv03RbDhnnW1ov9s
ROU3uJcEo9+q7OCZfCQaHeURUeAqfc1bXAf3wbvXOz34SV4AxZ3CwFppumkYzhEl
/ZeyJP9yeww9ZPsbc3axnOTvlpLuvwk0UzVngs8hfl1Ao01pG048ub2SFiyna3Oh
CfrqJZa7YokoIuf5pWStEePfYZ08OM2syOVVqjkmyNN702GiktlwrDlmc4ZbM2wR
eGLVd7ufCbRXhArDUFUnyc9I+8uaFp82xcQvfH3ODVHjGg9+pG4DnJqYttWvIknP
mjw8wESfRTE1WUm3NNlPiN4eOPBUrB3dDtakd01mXAnt/1+Me0dW0j/AxASYtoMi
b5G6FSU65vQvSjO7M+HD6ALY3pLhphlizVICn7pGdTA+SWxtHW1FPQ7uANcr/bDU
/GMw+sul1Lo/TLt811rSRCOMTK/Do9z0qTg/AGVu55pmDHxZwOGqyMxy7nyukHz+
lB31g6t15/y/51prCsRIFLIhLsAFOtL+Ned22JcOZkErlsyckJ5p8X8T6dO/Z4wi
ErkfXBrd2Q5xME7njN4HO/mXXXskkm5KC1J8ib5ObzkOvt37vlJFLFAtrT4SDyLr
teNto9HtVD2QoBE2jR/w4ZX9aE61+9pkKjNyfFsVppd/yyZ6EFsIN45qqCL1ZdHo
q9RbJ2Qf51mauKcYLHa/RBg/58ylbuXWJVBGNJVnjeMES0TyGiyr9q7kWAPSqhF3
pv9C8KSY4CkdPK+Ujrt3L9RmOJAWm6UH7HgwFCOejDquYtHd7vSAxN2I7DFGtIvG
fSXRXKsUd4B57wzFLAwdtIcyjUmnt9lbUIU692zljxjBOGG0lZATc1fuHd5XoqG9
1g/FJOLAcr5sbhurNXwnYtx/5DBnlo0SmUR+fAIM2Hh4wAGQZmRsjVq3xzrBvq4j
owB8DfMPv+0PJC97QODjn7gHTUuJD8N0RtkGWLvQK8pi79wZIZKLdk+RipRegXLc
oDPBrIAHybpieMvqH0X6VaQmejc5WiWj4aoJnMULVuEOsMnRYttQHOy6A6Az71qV
S9IjlcjFcY/Z00HbLF7O+uFYsRfQFVt/fkJy/NQVyFuK7WgbjcL48Dg5wNUGHbw2
EaDW/CjuOVEIhg9LNUqZ7b/CIOBFtUdb04tR5DxAoqM9i6Pjr1t76xPGwneY3WsN
p7p4B3BN5VVc6umpdUm6zWV3HkaZxYyT6CXbp/oIGKtNJxST1gn+bRcyGNlNCdD1
Piuwn7BA2bIBFBBhnSOPW19jUQPet9pbDK6LBTkH2Ew3Iip7zlXMXICzMfKG8cLy
kbZ0YLKfiRAdLm1vHHcwiSeASt7vqRh6KdfBVZl6XPKvB0QQKq30bqwasqQMlm+b
0mV20/8xnAhb06Xh4FELi5CubWTgSlA6XFV+e7jP1GeJPCHYSTYBHxjN2C1eXglz
X2wj6Swd+Tn5ZdH1d0coazD2fJCku2WElnPosXQ7ccY5xY4ZmgqiHc2uI3rX6E9B
eqx5xfmUtD0Mq9+ZIEn+oEXyZwm+Mz4+ZT4GiSQ4PGvuPBfA92mmg5/xvtoyZQxb
A1h8QgeECMY4d+fgP83FAG6sGHMPyPmZkRhXfd91EdpPt65IOdpB00XLU+eRr42X
kZOwpuhQ880zMpAmWA7KkPcIknlbkomjFOSwPNbb9Nq4bTETLd4UXeemBB+Q+g2G
gbLKymlo4zA3ccTVrEZiLox+lgvrHuSXpUJ90Jv2yYf6v8+vnpqOhbNmd4WiKMl4
FXChF1EFxB63LNK9APcxtkj6H9Ay14497tvZJgJJll334f8pHbjTzNNJrk2KBnYO
qh6bWjzRkLewtmuqJ49wZyILAI+UhsDujh3/Y0f3xxKha5BFpey/2ur7uC40dPwo
QkLzsOisq2kg+R18OgKljdM54zc5U/NH5RgHAQUQ03m2ewtEcNwK3tRF3qQssDwo
DlJdVroB3vRm6LXh5Yr+nL6t5WGWELhTPhC9D8NNZssWAk/5yD0FxlCGNc2oQ9vf
DKniyUAlYff4/sWQvoJKZ7C/u4vwbEsl9fcVErA+lT8jMlfhI7s9w4mi4uMZ16uq
kE/1Mio3gotAwMhzkD/AAhdAcMmbx+x0xKWBy69JX4hc6SMjIlqog2RXbEZ4ocxI
BLOaQhrysyEY7JSWws8owwTh80rdLxQYrUoOzttNJ7yPwR7csoQ7edxx3qmXb9xr
8agPxCyRQ6YYXz9TSPr/A6g1+Y7qM3661WAToXgstNqEmV9qFI2dN0Y9v5uKiuM2
73ud6shfi3sSfJgAmOa9d4x3YxMJDo59lNArK+4Bt9hlfUwlJxv12lPlYpoRrq1y
F4b//TMRJ6VM5JqFMR0cG+5+UTwLgA1oDYgzXhjwbErz1SCxQpxqB+5SMbu1FGat
VnCJwDUgnPAq/FhGQO7amWfNVWFJpYrTOQXfd7XobWqNZG3JG5d3fwPDFCTBb9/Q
3qsprhH9mRN1nofpu/fKLssg9ZT53Jvwf2P9KyKUcviOvkM44YL13zjFgvU7F8t2
KCEz3tz/nNY5us9z3X9Q5K0C1p5NeZXY05np0sigWaJFLWqc5CXvU7+K/9Km3WXE
Jwb2I2nc12r5wJXcFQ8G1a7fghpqSmG53tyUCnLatcGh3S0buJKAQBZ+vbr2PEtR
H8PIU+k9HkR2btulVOOFa22yiwmQsekU6p0wWTSLsUrRv1Nym3KH6qXsazU3ser9
Jn4fuXlXNEIuhHQx5/Xxrto7ks4S23YmY/VaixQyFbeI2uyC6L4TZj2OSqbSwTj4
yYehLOjvr3optMimO05FIuxjOxlr1CdFmgBiyAP9n/SoF5KdWnKTMm4S9iN65peW
FLOYvRpwuMqxbqefcBBwgvTiPaoVIgpWWYHEhZgvwlkcpY5kw6zaXDBSkzwZ0pMS
B0828XQmpHaHwTyz8nw3X98puMrroY75RBKkng/MlTpbPiWo5Eyuvtw5tjCE/MJM
kr0EL94LQHWHgH4CQ7CYxlQBI6KYZ42m/NFabeF3ZmMRRbPy9mLupoV1Ffxn+eT3
Udxpj4yOkjWwhWPa/3dDl2yctBTjOHzi6ofvdC6kvoPuezw962NHdUSptDFtdLMw
V0R71wg1Hl8pzKEgF6blgQ77oMbS8s+O2KO5xEo/gllXUcbFLH4GoOCJkv/R3vP5
LpwVIkOUqQmS3lNMrliapmTLjngrA6ZDBOA3pg/5mojXhqWVkW52w/AFplZyDhgr
M9vdwHyKX+xVuOzPXHm81Kc7lTLXGmYCbRdwuiQNxSNGv6+w7/gKMPDAbhFAfX6x
hjGhZ6lpZ/Zf06vcGsdlDcYrXTiZ91dEtTEb5I7sFH9IvJ6qrjOuWHQzyyj7SjPP
Vc+94pQNT5a0A4UBT9IOJslK1M4wPOEytpFTwacoyDiFAOdNXNxIFQCmsnXv6XCQ
6qLmTsfdm5Qng3vA72wKwJgid9oLUifsXNW/I7IpDae/+9u0+2SElVXTfv63LVRz
qM6eQLQL9htniFCE65eS/NH1amy6WJv+9etyZ/2NHWe4xiJFVZMs7bWogP7WpRWH
o97y+FS1nnxj1Q92buUu2pLvCjs36W6MPodTDtNL6HnO+JLjJKP0txHoZaY5I58b
rct+ui6TknOW1Dzq9j5bQZwrjey2rPoGdF2SOpeawk/LkGR4JBcAVI+haTQs9IAA
REAbgpKeZ7i2HnyvpnS+7ldYPdLc0E1o3ZaktbY4IYa4OSDdf+qNjT/OCBaLYDIJ
OD8I3YVEmmk58mHJUYNidFBnThMlwasCVNl4A8ugnRHRjvcQw/g1BnlJg/nXurdG
tROyiZyhFArs3c+8n4Y8Vg/7rrCTIK4GF/PeDRPzBCdFARoTwAYgBqJj6fsTIqr2
HnQFrJ+qZuCvOaiCwox29fR3s2tP33+FoScqQFR8kt7Yc1aT1LGIC4igGDj3l+A8
FgOmE4tPfXBmIQrxe42UvYFSpUhxLW4l7QNWrL60wTOHI7uR10zNV0L6GigwmaCR
zfinZLDnIbplet307uv9GrXXYa/ytWiNZXO8PJngq+E7m11p+wkKgbcdeA6D69TX
PrdSLHql2SgGc+xR6Huq12cvckWAJzDuofVJW4cHP6va5RRb3+jfYFramluMp+i8
zx4lgpEJ9Nv8Apgh8301sQb6Shd/z8t7fTfptcTKFYPy+UvQNkV49bkFj72WAIFE
KgRpyc2deIGElUINRbEJYvUD/DjHd8atJlBbUM0oRz5zA1TLHaU1W6ie+c/klXMh
MTDz3nBk97UrQmXh6RWJiac029RQmwNVc0wRNapok4Bu1iMifPTsE8/fSmeBIIjw
ekEEa2/jyccy5nFeuInz24woj1l8x5Wc3hTjE7dWQNGg9A6hJS7cyAa6ix6Ss+9r
XRB/XEHEo5plRUW6UGCEqTB96a5KyUy/dSpQtp2+7aRgm2HfbMntSLBN6OFOZyl6
fd/hRuH35xZr+Gcagk6Op3wmKiwa7KxNeANsLLoZAIAU0pdK4Ta77NBVopwyok/u
A1faZj848WDnFHnzHNHNAqMA4U5iX5o5/k0sytdUUN+O5LViRuAlZUAzkKHAdWd9
FGQtqOCMgNUXSh9mcZoa3kK5p2Oc6Bu/Uk/cAOMQhAs8JKg46RV5X4PG61ilC32V
uKxpez6vr0mIhE8s6xLzP1Kmiq9KKNJdFIAge62UGaoS1K7lQXstOaxKMb+1QXJS
QMWwrpL9kXe+HMf6d2NLXOimuZdjr7jKLCD25LClkSsdflauX7eyj9W9DGS2k0pQ
kaZGhdxLQr8E+c492zOo5WDRmeoxqmiRuppNqgJEP6Ygl36Y0aLnQUyR+G+jhZe6
Hm2KEFXoH7BqPCkZrI+KGm799kpqw/bjD2kiGir6dp7WzgTbiWVJJXxnqUSwhGxA
iC1svS7XGM0sLSYzBHJ+vtAOyj0gsAgM6+PjVh4/1ck2sLD2dQV00LBmcwEek1Q3
1QJjQr2oqtgEvojy4yZWS61LbdFZ7tTtyzzFdPPZ7OjyatTSAqmFfdneZUTmF0yi
tK9Hk0/GNx31eZ9sIIE/iuLiqbIGXUWJlkJPsgwWw333TMiSTHeqBwOXi1h4DBwL
AHodVZ+etdo2dVcs1ipFr7w5PqIgZasPMcl+2K7vnuuhL6cn2Myz9qnSNaf8iDG9
tYZX1UkWJzZH4UpRC9kOF/loShBfa4DecWkMxnubacTQZwv84fhQfYgeY9ubQfQ+
MkWAjDa5JgNYqxodRionpn2dnAg9CT6acgfMAPs2SMvFxjcOMkjCABobax5aCzKR
fmU2YKWeMebkp0+yknrzb8sVEPKXnqLeaZfFS89ANc+X95jyynE3Ijw0FpG37iBn
6k+IDUQ/HDd9ySIGzPUArUiCUSSXkK8UqBTVqUciv7hGLx3QruvVpB+0KWdkjnKk
pG0d2+lA7o27nU5Yp+cyUVNeNNsWQKLGLWE1jF8ZjAjOk1MjCDXQZN/AXiSC1r52
b1QYEWlDCQyPtwsvwuqyNiWfBtSi/CRbGr3zqhVAPHKSet6/E9U1+ghrWa9R1CNR
8X6Potg+6pK9Ve6d3dMkctpSBnYXSL43Ex5jrRS8z9CoIZMUVCYNhnmzY4jSphVy
Rmq+sCr4pYLrKFiOBVaCuVNeRF/nB7/2zWGzPlY8ibJTI7OKSLV6Xm/Ee+eSyKr1
oYhBJ2BRMrguuSo4tN1BxH4ZkDA4FVj1n33z8h2qULh0sD77Df0Z8oXnu6l6RYJ8
XcsMK2mXyk2EZsusHGwxwo+zseybgX1Wt53CYCz/1SenP9QD8ROXiu9I8T+Gmz8o
YvhFcCiW8yevORDklIuvQtcCaL0GX/2K2kmUK3GhrdahCcTzKWimIMpWOD+t7KnL
sM//WnPyxEYCyAZMbrmMY33aTdTuIy7SjoO8bbO/z3KVFpkvdnQ7EQX6QHJSmhlu
GEdm+onqyD9ElB2A+iMzCP2NaPpxnxLP6odyFubZz5/4bnro+clBdLL1KDdVDf00
fNoaFLqa0vh15x3xi1MF4quyEcFVfiRCG5a4Nb2b7QXtOv4KQHAFs7yARbMKMFIG
pq2mw1uw03wjYhy2rMXt08HQP/b0YZMPW/+dvQ2etItnvqCq51QH24KFLmTcAt61
2aKUO2DBlq7ta0k4P4NHVLnLO3BwPJFPPAlyuBgFSM5IYqZkAXmrJD9q50lFXFKU
kH1sjP/R95msRFS6V+iKZXHGHKWwT2ahQsRP4qeJNq3qw4oXemxXKkDRTcCoQNq/
Ou8ls77wnH9PTJWGJeOIsb7FQfvCs3s5yY+e6M13nGN6zQxtYktF9c8g+zHjp1eJ
bujPXUFo401yetsMMi9tOLxSTRJDwmAeW+ha0rzccaaqfTGK8OF3GzyEGPdkQH9P
KuFri3+PhGBF7Txaj6SmvFeq/HlVk4XrjNi5F4lxM3MgaTV5lYHyErwDVzXb8R7H
8OoVelrVd5h9zhJWb9BXNny7CFliD9Kc2Rq1RzWQzKacSN8SHOp8TfRTk2PyTc+N
vrld5/KH1salHUDECPEyniBT2Wqo+QYGWwSzt4nUY5PzzcEPbVDzafnP6AGON0zO
QrGY1M4bsHUcezu7TVHuJuI7luPo8t8zG1qw+PUcBD9YvflGzq7li74sJ5m2gQPo
FjDmMjUK0kqH/L+lFu2cL0dvtItn2dFLnQw0vzI7gMYs1NTesYC42RAA9lDiukaY
pAbE7x8lpHQzj1tFmhXL2wHFeif9oo7koEGcllzy4RGNbxhm6Wx9NhXPn9fK2UD7
MAne2YK7BVTIcZxD8rk1lyzpsxbB3e0XX7rtFh+P6FfgNo4hbq+3TsMQWHT8Td19
eAxMQWo0Tozj+jn/xxMHOedOu3ZY6ngmuL9nuMv6cmAJ7AeH2/Muq45rQicjLy6c
Il1xpbbTkY8V25wxEo0HVPNWyKwWfTkU+9O1wsbvEz+OarWavpfaZTDGO4mjEiSC
a5JhBZOs0MP4QuVL7Z6MZp4U+wtPuLfW6j0x2BOUH3CHG/XpjK2UpEUgudqpjnmK
sOUKjxjj+cd+J5Bx3O8sBWO91jQ9Khlf01c8jmGzASbP7MuqibFg1u/03R+fIVdP
oW/fw6Ed5moqa0g2MVS6eeocCUZkt6X3X5MJTSa8AwTOqTsD/s1mP92m9pEAQn4K
IWx/kSjotLTBk8vrHgNkUnF0L5sEkBjFQE9cJSx15NF843j9sUyvqcfXwMWA0i81
mXj1bo6gI2sve89YjjcB9aEpVuCYTvRWbspu8xJbUxQ8AYyaYS5jzIjQ85zWkP5j
Nsn0/RdmcN47QBbUR82fbZwb7uQcxly7c32e9rHJOm1oR5iKqVxPcs/ozH6lmzze
nxcFiLrvAk8R7DHd8FM5NI04vPHNtvhi8pFaRfEHNNvOvhvT2V00tZVonJtfw3wK
Sx/M8QpfT7KIZj00gqsyGi248FzllLxEItd+YI5z+EZA3kS5nf98opaSvzZwf1wT
TRJ0TeC3GoOfvdZOKe6YHASG0ybx03cza9Vgn27RTMbYLtbWWsvEI99+3NuTz8Y3
DV/bP0gZnWr47SWnbUr3WVT57NgnwtA1uyCH55wpWFI/gT7yL59Os3IeNzbIzFWF
7OB9LshsZR4wg79WwRpVvgqe6goJDbbcJjvwhCymQdLFLjZ5oNY34a0j7+M5DQgy
9ZK6TbfOnWYUg9E0SD4VYYzmKATlvc9epw5B98pCDDYjtJmqeLcO/oGU5V0a/vhg
d0Or68ZbSzjJg1RhW49LYwTdeQp7BePvDd+F7IRwNXVaAOlgLCLTDCy/TyiD2RjQ
MsnhEhkMcnc3hgidnQLgQd41IFyC+ZLLt5RVCGSBS8vgTEkhi01VNgFJ84FhehKy
+/aygshOOjfhtkmA5NmEdLY13YjzIcddXPJaaWwo4QavcCK/hxYilvQHayn8N40E
xLVUAu9oDgu52grsU0ime79uqwBB2T7uFRGmHjQKcdLsC9vrDXKbYzL6KmsO423V
BZ3/+fHtyVozKS7lWM2YV/vVQBxq+ll5va3C3FF+ezkIN2Zz9zoNYQAIK9zvTiGc
lCflVG04JUMvjTg3lVOfGT9DY0d2e3TFXs8T6696SJBW0++gbsG6WEWyRHOsHAcB
lGnwlgGOX1KA6o10ic9yOhZBjrntldmgw0A0VhGoCU0JWyFZ6Wr0pt6YAPx0G+qc
Xaa/FVfBLtT3TcmLwUDCiyJeyxnUSoIlEBG1PwUv6ZEyakxY0rqD32YGfk/yz1VB
8j5a/fDKbsQ44oy3fkVtrkcPy0Qi1Id20yI0T0vvWaOG72zJ5y5qTy+c1aSDIRzp
R/DXEeT/fQDsu27CfBOFXCRWi+MWer20bdhJeo1RJ1gFyHvEA0aIcm0IHf9dAtEd
+85Yh/T2cNHlq/Xd6c3pHJ29j7jUWq46tPwOn1GhOg9eCHQ7XFMY0gO9YyRt3UBg
vMwO1Vw2DmzcbamdL2KyEbn6JK2uC/byqkMMNhJUU6QnZ5Qd7j8BPFJP+IU92A2M
G/xgPG39Z9+ZPLhVsJCSM+0Mq8Q+HoIboQ0ONJyPB2t38cCPeAXUK7hne55hZTdE
RYoLHTWPwIzcz5u77H3pwpQaOGOGuBX/RQzyRpdiEN8GqcWOwygS3XwpeLB/MXpc
hI7v9HwE3gL7ECgicWnnXdmr99btQSgvCmucGvQ30+DxhVaCLcqtBSMj7eXRMkI1
Esi5h2giJ3n6UTj3RtQ3cfcgHoLYfwkDheTo0XdnUTuzoq7kTxPdbYxgenskLtoJ
cvmv5o8psDgeIzc606yNKFsdfe7hsZwI+j5QdxudQso3JL6APnd64GdOSH4mJYNh
0drcJATt03A7cj40NMB2WZsEUHQRFRotr5dVCIWtCZdTrQ4HSaDb+f6/d3V7GelM
i9Gzrup964l1uhQXY2PCutMVRUTIbAZxOQg+5beWae2GAzxOI1FY3IbAb1L1NtSK
uPymBKN/aKEUVe0RTjciGCRswFOmPyCRvfwQlH7NJJFkMz/Covftb6Vlo3Zkhg1S
epGdMOILH9kJhkpFgCdpRfqyIIhPdEHGo59g37fwK6LRVZ+ILZMJp2OTkyrX7Ykf
2YOiaPRwu2eoL50sxtOPscMddxDxTw59qlHO9y3h1TIAinCaF0zSG1aSv7lxEYpN
ORil1F8fTCAThJTrjODfwtku00cBr8VlAd9iHKbOLae2ck/MmRPXhNn8qHs9LCZp
XzB8P5iS2fS0Fe+vJVUYKDr5ysLWTbre5pgYsCI5eqNGiS+89HqDlt4WVTlEARG4
silV57EfhKTDQA/ZqOHhWKuL967Ar09j+TVhLGYlDBHVyW96ISGBL7j1UtD4beXI
uoDiFRoZ4OM0H1zCAnY2qpi/d3iUtCmaE0P1X/QUdJsljIfcQFpfOA1qo0cmiJVh
V9rfTFusadChsuqWqmFSCEgAtlF73CZzyk54/O/ot5BG0MaLw2huxo3gK4OUqG6W
Hf7NcBXZxkYxzuZq7SpPT2Nc5/pl4yuTAee1sbuSDvqjqGFij0r2shv04fCF+wtq
P2MW3urLM1PQR7LGNjfRLFYOeaZ7jJRInZXnpVVg2J2wGMjYiQgO3y/O/s1yiRtD
CNqmVR2SGk5ldpTl8sE1X/2J9qpYGh0Q2bjw/crEREn1ewRWxZyYYiaHrHjqnT6q
htXPdHmU8oWU93l/D3UFmY9AzuMNaI92fTpi8Ui7tENW4J8MWpz+LtzVhejjXGJh
zTeSd9x3widDf15ZC7QPFDoa3xw3CPlIo6h4XQRECG45U0nZ69VBksHtuioaz7iI
Etrkjdxnutzcqb2xJf7CHCoZL6ty51YYJz9eupZU6CqpipUBlpyfeZLlwsRi5rw0
9oDm5uQKAYZzkzrAm/RPK3xqVrM+sHYbzT3OrWQuxso+2zsXfwrWDSj8vAH3VLtA
/9qY81f3cx2gZUwMuH/O5hhYMzJkOtI8im6XF647UfMbRSM5Q24WB6I7D6TJOu9x
fhglD5BZd+NvMgJFNATB2I0XG3MxSn8GWSse1G/ySZDgJY+zDhNVVJaNlAYd0ytU
21xNR8apS8aJJEmF+mCtDLOpezze4Gd6LwRV0/+xynyFlI3NHqH/irRnsaTSmzVW
o6gKHyJ52/DL9RJRGOEewjjuipAm7VfNBB4/1bj0B+aie4uIBpvatg+D5oDzCb8C
RslRARoe7HVjwxqaZ9v7+WT1ZKwloUNmmkMr7zp/5xngdRFVnO68kdwychAlb9qK
Ido2jlULDGepmCxwPlgRBYAREukXI/t7KR4REU+qu0wrr6gFL1PZ280OpFFMruL3
uGQvGcaM5vrYSXAW9A6/ZlKTacCc7NkRmxD2paDgYBMpe9zWPgPdQHrdmVuZ0qeV
Y6gF1LNO+pXvXrm/6Vkok92ez4+1r0Q7Gl+e9dzTbJJ6SkZ4M50oixHfZdljgte9
jPXTUDTaUGReKv9pBB8J/Xe/mM1J3pyncabOgsegxUdePMJ6ozgDXuwHiejQVHNA
l4NsoFaetMeDH6e4OYB/vVY6tqIKuCnWrNZNQW+WQOXYbkgjRMWKeFWWj398FJNz
4s0wjPci8zcTf2U1hvvDH3/MwIzn78C/ylpPnNhhkN5IvuLTIAGtu3GvXStgOKII
pBtS4DCqIS3LpRVMFbsbRJg41Iy2w+/o38eI41t1fGYEMAto8ruX0q3lTx2TnqOr
qJTFZpAQLpwXuuFKMZWUdrNm9MoT8kBuDO5VH0T5EZLtsZ4izROnWB67wwMjQ2g3
3+A2P7t6UYzbTBjesBYSlmTjzF8dwwsBra6uAavBO4ayOldkuz6oioRRu0RJiht5
nOG5ev2zT2D0VjGsdZFBh9HLJqBjM7kwykFJtjkg58x04BxyAa7gDIe64lnSFKHp
1Erx/jpx/oRxyZKV6IxZbnZmy9ERAi6iFHAhS9VKf/PGJa8TM3g79yqNMkESR0iF
MXOmR2BDlV8g2ShAmGmfp8iFae6Rv9FvJosfQnZKTHSRNeFgAHhnuaBDdV/h+kZq
iyq7iOuZTszrBJsp4BzAl8n29ZnukB/QmIBN7RuMs568m5q8T68MUIWWV790lh3I
zZJlQb+e1Ty1SS0+vXBSjNFXfdlqbp9LXS2lg+zF4PNSItodFzy4GgR9CZgIz/P4
udUP069HT4T7oIqCqoZQgB+SID93H1rnH/8kXBocVcQchCOxJ5e1vulPog5t0J9u
W+gVtPVmQr4ytHgPAl6ZLGHt/K9vhbY8+/M6ZFDPzsp439lLcn4sxRU9LjtbzUUv
G8Ys6jIh3fB0p+f335ouCp9Y4IplO+zbe+27Tpre3Xa1JkVPSa5rscPplLQ7xT5I
nnpGFYX73+AYiR5rqjFWmhlgTtwkIoBaM7Oul1ZbeHVZfHr6PjmtnU/jxKYRddxs
QxO5acGT4lFvkYKk5xpsYoWiFcPxjMjgDYd54sEPoyRnJlhZPahmR/UCbwrfBxoy
mUM95z/iYcHMFJSdJmWFsDQgSWeK+VczS2Js+m/4bApz5fJnIm08re3PrX216VbH
mUexqZN5YHA/uIte83OQfmKcRV9JkX0Om8Z/8rKFH6wvuodK9VWHfyPiqWgYPypl
kBnaPMdfRneruyI32sq+cMdqjHf0aNoPzk2d0rDcgrXEQ/hTndnCYuJdV1t0LiH3
SS8Sp9T2LNV0jeB6rznbP+qX5+RPnRWJfsb1unt1gARmY1lX1tDfKPGUMrqNTDjQ
wUo7ApgrWgK9j0Qj5HpMoD+IYDGxm2v+vtHZRwrgoRYZHQB8efXDQGvYx3OiBfGo
JjhR9ACzoe8GSgVxzr4k+VzqrfzxBdP0kbX23SytfIYq7ZvZAezlL+Fr04I68Wu0
YWPQo69FUijT/BaQb6+bDY3S9sJK5yfVkVnvs8xP3IRMYZ4anJCO27+4FjFIohlD
pP5KZkNWPbXdeDDk2unsG5GcnKN3/bCT6uhYBshgbdSoJtnAPBP74fwfflfWRkou
Z8VNYZT/g3pKW/M1g6qYWCQxjeUUGVn5KxFr8+UypjaL4RageFDDABTYQErY+FLz
JrzvhJVx1b/gC7BP1rpV9/65yrsWlD5qJsiAgqjPHGST1hXp0nP+ZfAojy/VapZI
QX0N/BvEBrg/sPAkS8QQg64Rc0WRpBLhMBn7fc92VcQixvAW9sqbesfflC2ambWP
FwHAMS0S5P3cCY6qieQvC1XYEO7Pj/A1z9Gjkdi2+E92d5hwuNTKcGuOzl+vBy1X
9Xvk27VXLfG1SbcFwsp0xkAzbBigEvZq0e82SOjUhS0oZ0p0Q5njtcxNcY/xEIYU
Awh/9gA2NfjxN6mpCnXzXFIfLcpABERURjR8NjmNc7XaFlAZ3PV1cTY4n99Qq1A/
3I5UibFnkCE/EY3xCrAgEerbnKDGg+TuQ/NfbBkINz35bNOoBh/y6J1+RvTxf3O/
1eu2Yq2D1mPOAgNGYL5FjADAp/KKlUCi0C77Yq/z2lOW/D2rb3NUdBUBXn4Vcffg
kKmVCPDPi91IGwhQ73VJ9ElIZ2skBxH131yT/7iDYEdJjyNHlBXSeYuWYm/eXqV5
ikzDPDZiM26HaSWKI8zQIsYcbJ1T5DyPCiNeN25X55K/AJ/AZ13Z0Yb34/7gNCAt
4QEf4cD37/KWPDVO9YFyVU4ULdAWx/sBZe0YCvZ4runPba7U4OS97SEJdTdUYhBi
ZlGwIvl/8r8Cos0UFXMpl9PeYeUReZHWzr6MNRWWLgjOKfCg5B7cMWABSAjs2jZe
3vvAXJmn5ZwByY0KXjBNJU9wePkonpO3Kl9YJ6qSvCoOWSOD8oEswBNFoo2hngS0
UJgrGyA8zWUB0AzvmR0ZZ8GwQ9eo0mLeWAf+r+2MuCk5EYhDBQD6gEzwWqs+1xbW
sAW0v2zXu0YEaEud7gch6oXk7wbeEEim+CKBHTUX9H5jcPRKA7nNI6fTxUlLwFfm
cmXkO3uek6vSG2UxP9nhGAOP0Z8OiJFvPk3bWxBXtrSugkaTTrMiwTzpz3uUKG9Z
uuMY/dyt963ka8wpXTKtAZpBN8MctkDpCTTymsw4MpnBCGjx2Y6onOzTOP4Q5Kea
1n9pGSQrXtleeUqnzoGP7iCL+nScDblPcCxHm+FfyM5X/wBu5nY3vR6m0Jimt50M
q1zJcjrLC1HVnaNR+wVic7lFYHgUbU2cKO4RcqA882V0ZVe3MHwYTp16hUGCGBl5
FTueHgeiPx6QCYkgMkjVYZmg5QaaaklsaD4Ma4d1guQ9UV2nuZo12IEefa9L5VNv
cbRVwzuApCJyZ8cPAes3yirKnyPqfcNwiJiArTp4667cOSzHSFAHPSi9P5wIVDr1
uLWKGljAQCYLytL4VrQlcrDc28n52uV+dSmqq7pI5I+1bMsxZcrPoSBDKvLDa5QZ
zGyiuax+3rjaDkwBuSmhsEWyXihDIus8Dey1aUNG/RCsl+qEtKV3ub9HJjqNF4pK
Y4mwafq+yyF5pLahoR9zpXe44J8FwIk2q6RoFMbUqkvmYV40Pnh/9iXeNS9ScU2m
q6QKFAQ/qKVY8F7iKnfhkWq9SClqCaggVPdGW4yDtv95lyG/syQQT+IVQRDdwPxP
dKOuYX0q5TfIOIIkmENoi2FFGT0BvNG/CwOi623GiJkk15d3eydwJuu8rvOpu2Be
NNK87wz471jmESFkN6ifESS2bncfmARK+eTBw58D8h+1ZBnmitqkW0HMVzAwcLI2
mN08cXZTxU7hOT+A9i8XeRFeUYgXpghWjN3kg05XMd5XcWvTsufgH4afzaTNJmvV
Sw9VHQfErtKojh2kcr+6k6va0E6WwYgyIbPRx17zspmarrauif5aaI0xQhuDBH1J
BqTWawzEq4E34D5tQqviDYVrRpHrfeCjYJYpcorL4aQH7etA5oNr2wyTilkFRLjc
I+feeG8sx+dQ/iOKYRF1t93BVVUP1cS5DviajnYOL7dxYFUWej3A+nFjgaIaz5V9
NptTDBpH4A/p66ooQlzHuNJMT3DcasAK1EeCqnOBmIoyDoN/SnGxP/MNBtdkSUnt
UT6e3nkXbPTnxftpFkHA8Sd6wVdffBKPYEOOF2wFWHPZ8ou+jwXPdZguX9kU7Udi
4dVrNxMsxoJleSN3KpR0VmK3wARTEXoCdyjinmHB9PDgY17kwOF5gpwgNblp+jXh
sQUh7Tbv3A5Gd6MfyXWj/8WZePNv0M0G7JKyQrvKMQEXtS24w7AZv7H3nVHLgihw
B/IsChNnPfYdFrnrA/jyQgKGFke3tvWPCw/wDy+cjliVptCpKQGkIhkyIY+HaYjX
oyVK3qL803XL8eYVGSYYXdUS6E3Y0WolVG0ov7DvQWTiTZ7nVJAR11L+V08Gr04N
a8C8Sk4afHgNcrbNOXu1rD8/bTh4UkNrIDd0SMy1lQVhwa7EtkNNIp8DvDtas6Zp
NaT84AdETiuTiSmJSoPUR78s6A2BRhxzTAQJgvaaBbBKIB6auRK9mI+Jyxezz3NV
+71/XtxEQttJ1gcvLy/serzP5n42BgKq0gfNMtfXNcnESmCVTrXNftNQvb1U+YLd
BEh+WcooWITHHYKSBqDChYE/rwpLhxoKtoFvZOkMnUQsIf9q7B6ZOn/aexdPlO/m
Ly5xGa9w5SqrtyYY6KtyN227k2oGyb+1/Yko8HuzX/9Jv8st97GVGtoCy7n4zpgs
b+MqqZ/QrYahQK2hwAwTiMPj58OdEWqoPKkj8XcKlKc=
`protect END_PROTECTED
