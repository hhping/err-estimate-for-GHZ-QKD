`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dg97mksk+xnhHv5XLue85r+LgA1VVL9sJk7vnOobRMQdOHECua9OveFkHpADEQsH
n9P0RopQWFzbidO7UEZIgOmKUg3QtcqPWnEE64NRwBUtf2fP9s1xk9czHFH8cCj4
TCnfFLCBHXrmfAO3wLMRyMyUrNYvVzEJJ2nCv3TBRaQR2O3D/KcQCoQwGl8TRDbb
jbwupXguP5D3Y7HPWMVzpda1r/zdwRSLAmunAOPdNEmsYUGRiwWPTDulkdFiG+xT
vX/4M5XbCxXadkbfKcxEfeVix8z1DVtBuSmt5K+qubcFdnn0QzNov6O362WWgCr7
Kx3bKUGAraVsgqj3wAivbGixCGQ8yGjMkjCRDpbiboZJQ8kW8Nz1u6jThnPNS6u3
i8I/+5zo8SoJs0ns/S5sDpqrP0Ec/Xt1K+usOb4ks93UBYnphZpgvQ4ezh+Gg2TB
EJrlAdsxqIFKy1TCDjBoJAhwFUH58ffaqXRc38zvJUzHiRejetLpJMtWp5sf733V
NJ2Z/qDUhiR/qOWH1OjjcKgvIJ+iXV8jHLNNgKJhHarJ8dgxOibMWu0/BOduH4DF
5RyDdqr12tA25o/v6Tqiww==
`protect END_PROTECTED
