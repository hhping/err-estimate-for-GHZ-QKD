`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k+OAda3W7/UbG7OxH5LcN0uxhvN1gJ1VZdAXnwduW4PgUbrIByms/IxPDwLXfI4q
eE555bG39qUSUur68o5L4xYoLipQG6Xd82EctuV9B48RdS3bXgvmtarS5+SAAwSK
sONbHYTxFrMPy9u8FQvg6t386IxBPCacfAG/TXNwYIJcJAV2cHEzC8q+bm3J/+hU
+M5aXnjH/5h/+y/bBUcWbUZzz50dftrbQr5LjpkTX0nYzAe9TJEC4yQ42o46u0Dg
Z3lY9DVTS2vkhjXYv/lJ4wkyYqesENtOJVHoHjCp006DJEiTCYSvupBYDLi2Jzq0
xtY5HUxLre6wFZpf7xHs7WPZpPmdsOjmSNfmFCGhzq2XoY+kria7CUjABIhidhUK
7TOEvfrL23syl3XVUmVtKmZTyCwosMu0WRcG5OO3/KDS2S49J49xaaZWYJS78Mf4
Tp4x8jT8BomRzZXtXL6E8amKT8GeP/CAVRESSF1PBR+5385wOtV8RuQ6X5ow78Z6
O/gEISyXKU6g4chjeKgVhsjk5EoZ/EEZQhhMrYIU172SfkZBfUJOascDtSBL0sIu
T0eW/nIly+A3wVfh5VljqZJn8fcrVO1KF5wzAHtLI79iS3hNGrDj+/6cjOR58sYV
zIHPdmIbfqb4A6PZ6oCtWSTwifdeMz5+vw2jVqO7T5KwOm+qX86WhqN2aNCTeeUM
vBZp2SCq5Tvh4qp7dTrvluWDnAJu0vtcYO8G6dBUbAKrlCCF4poZztekA5iK/bu4
jw/pnzkosB5pMXROJh/xulr2QUQpHBEdPMnwo6bIuZnoJgeAKzE556ezoYnLWMCc
dMYFrB8J2lBdQFkSl4iUS15W7UfHG9Xi1UfGmAk2qnTiqn7OzoHFlDrq7MRKlkqZ
YDz17OxBlr4LFImM534Lo6bSaODxPw50twsbQeTeOfA=
`protect END_PROTECTED
