`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fjs0KbdT8SlJkjwLq1pIrZazynFDeILU0xb6FLc8IDhvrXQbh7w+bw8K7eoCy9E4
CGKXMbAbQwmrcruvdWO7MzaypfpcfZxIZ+IFpYJUrlKwiT1FgAz2qpum8ynLc5Qw
lDxeVrGT8xxcO8tUdkWhIHJSjzUT1sxIfvArqVvNksCOqQ7kIwKguuaM3UVvLaga
RRQ3ySldhKpvvbcRxxNSHl/Tk1VeLuroEN3kciTiNfO2U1K5veaOZDdS+tpMly93
PioEJAM8MYMNshWcxRGr8HtjBJutDy0uLGJd5OQgtJZmURZWRRkmLVAkzPAtQ4Mh
SyHKy0AfMEtP6bAO6BjJbQsU6QHxzopR68TTkt2IHpQ3XSoWHwqe8MeeKwV7WAAm
a5XutR5RVKRMFfzu/duYCdM5DUOiBepKNml5nOxicM+ws0mx6wzfOq/Cn3J1wuGS
Keu9DJKcN2SwfXIWh/WDYsIH0XVC5se4qSD+qtRYxWbQit/f8eHo2tDkgzlrUxDZ
3r59gTM3UORiBlVys2y58VRjhOqCxlNvcVFqhDSd4uIM5BTkbgJyPr6ROSmPzDrn
RHBSU7ua6CkOoBgqMatnKlok1OQs1x1ysLsdMPKbEKs+ynqCjvDGxIULvrSHPWBr
c8iirMD8CgfyFnqwP2BqRJwjjMepqkGlW0WfElGhRhcmkjYbfLkGqcW1wWN/gozZ
h/8B2I6QEUb0oVJqyV510eFOTLcXoYvrVx+RNyYcmTCTvFIb9JLe6/EeUOc5uXbp
7tqArI4a+TeBs0vozRHtQdxwRLUPEXLItcKhuT5wZ2lsBwcNQTpcYA7TjRll+rRa
8QdIf5zH+R5r71Jh/v3Mgiu2TewvYK+8Pgk9wdzx/v2URECbJmD2Ix79wiBbYEIN
kUpwBu+AtH9SzHRGtqVGHRtelnzd7zoCPwZLfp8HiAIbdTC5iwJZ+IpD1bajpIDH
PjL/5a6q/hVcA6KVBqW/yT6z5cPDrW8B12hhrTiQXFTbsdvoKPNC1JZUuhcFWlvl
fNwTggFrAwAQamBbm3ynCk8IG0LVI/9KT+uchap7yFkfWk6OyZLXwydmOjJCPvvT
ZC2zf9NI7LHYblFh4R16VWfFQD99phWRZCe0EWDBnqIviKDppg6Kef/yvcYTjZ6s
P0wwtJt9RfD80Ir6sCO/OxC5kyOkZphv8nuhALlAgmuMflholNITzJj4zTjWvWKu
NjQh/HW3P2sne9j+ySpA8QGi5syPK+ktmqK6HEkzvFN9MbIBYF6o3PYv+/GV0aIZ
D21zhHgrfCLR5N+TNhjUS3TPV3h2aSGjkfn8da5IIF7/Ws634mfG4pvaWURr32vN
1j9qGTXzi7VJcdHp50nXeShfzU9aPr3dnCWV3b/gLaAQ7Wje96rzpPMlMwml/m8O
PM/YpicwefyP9I3ldqak8inNCb5f/m32J3W39eO2lYb7uhraA87xn1IOGcI2QrZa
r63wfRZCYWjzP+M41xMFxHRV9UPYg711L0e4YrjykhcJ19WdFR1hl87E1tLwrJ6v
fH/1k1mK8Vs2UEg3QChke/DzjRGJDSTJ9cUltyD33aaM8ZvOqoJXeco5W0J1fLzO
dWLcwHnUpsrUQWPRBTSP/hM0/jD/2Nag089RV0HkWx1QQi13xv5mm8B9mxgqfIVh
/xixVnOXglK+fVXKOAB4xxLPRihGYsyDm3ft/jeygKHjv9mMAEDuDvanGQPeJ09m
9A+XXEvEr8uqbSUOMaUoHuz2H4/FKFI8vles3RuPLjq4QQ62GzrSN2MxQ2/dIyMS
EFba7tBgxmg9NRlpgnjNVZZmEWPWGI+wCLganeGrbm3EQEl7oCS4cATry5DDywo6
0lIwNlq/XTY4/OMasc4YeC+j2lCU7afnoFC/VmiPM70qW/7yp9C9dVBQmIn/1lCh
X8VwZi0cnUEkK/0sTmjgRxWZeMBxblMbme+JLsggce+xgn79PchFavnzyyBcUAAL
8erUeEewLXCIX36PrNkj28jHIUJ/160rCfGZchqFMWrJjTwHSZnPNgGSlGGYEAU/
5ucWa3kZpwm6pLr0YkzskqToyvkvnq2XhxPSioaFWRK1EM98Go/G4MFbJz6SU1ET
ZuRftFVdj+nFa7rJUgV3IyKkgOSEzLqDNYE3N+JB9IMBamC2+Qkp2AZy6Sr4JgCq
yFPW+xAK+JslKE12Ps0kczsYfv4ukscJPEn0zl7I+d/CQdLZdHIiOOeIFE9SCRd0
+X4xHWLJ9ktmoHbxvZR7y+4f6DzO9wNz4QzM2rr2Xjdm7asnYUKAZL2eVqqFhJec
MTjfngYS6rizoPQkwtpXujaobg+W2rkQFTW7R4F3AnAPt4OK7fCDiaeCQMHWL0nB
Ii9qp2iTlmJKb1a9ehnGkwntQoQt00pL6EDI9K52tTXxozlpdEg0FcIbnd1QeOB1
2UguOu6VVcY5M9r8R5o+0x2D3DndfBPv9mjBQWP3g2O6cXo6oWtEANLPX1HjO382
xr1LAHcoQWpCNV5y1Vz1+KD/IbROHf0KlE5KnhDtkMQUj+EeMEmF5QRvw1uMhA1c
kvFD7JiqbIu8Wf2Hwh/m6kg6rboBjkKnjikvGvXYeBfHY0eAG2FeraPq98BUr8OP
0KsGXG+lis00rIsJ582ougp0omkYM7b0cHCg21L1w0pDjYofHngz+TZtm3puyCSE
iwppCgjs8rMcLZ8EhUEal8LqJExoGFBLq/5tAK0ywfxxhaC/mIM//PP9UF0yZY/g
/10y8WC6p3rTbqfHgr7LLbA1KdcT85oyySHlH1JKqXJGUd7MDrVjDwbLUVW2JibK
vgqW5zwCf8k3NoggUSlv4JItwZkqVQcMDD25DhYarMPrZLvjdF1J4hLKl5F8K5sC
ZvkRqGNbjCbwqRwDB2KvimOnkl9LchoLbXpOBqt0S3s4uTsiqUjXc7ap48bWECVa
yKuDEa1QVAJN+jlNSmg58C39fKCV+EnGsemQir0Xwn4sesbd8o3a9CgIjt6bJapp
6a0ShZYuPkthe9FBTOoaRSFTn5pVDf0Xqa+iBb1PXgoLyP/9GgJsZsIyc6M9/CtU
L2XueJW13fyYH09i19M5vt+e3igiAzClxi7shLXGrKs=
`protect END_PROTECTED
