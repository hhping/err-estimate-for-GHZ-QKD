`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yurlRyhIqFLZx5PSAM7+Ho41Hbi8dffY77O4Lf4ZOIWhCBWTkxCmA/wdkGhmLYqF
KrF0y02Lcuhxi1KRk/GND4UX1QQ+xdPipetAjCfSc8+6ytAzBl9+slv1G7iwCDY2
FIN/es0XHqaah2gjJO/NCr9F6cQBbKLeBoICVVlZjhx/jWxRcSv8SsQWFszlrIG+
nVY2OldpoeG/7qlPMKFflcC64iLWc2fO2vaFFafTLYCPGU6tAvJOOrDhJhJ21ouA
hd311vqFwwT5deh+NKN5LlqEPnvLkLf3aECtQ9CYBbpUh7Z3FeFBWUjmYbG0wX6i
8td1mOjC7dZNa445NTbeTS2N/I1gpZQY1WWIspZUFhK2YeY5pf+Omx0JG6Pj361l
FqwQ9cEt3ww/BnwPZ5YOpMa3KFIqmEMwqWuoBdcNI/RR+WhKnL6AJlqafjinBcBw
`protect END_PROTECTED
