`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ArmcuRSPx6Dt217Uvoh0OIwutZgGjBh6MjCtm3aWxsqu7vLoFYSDN3X2HBU+o+Bn
DiQVNIdKk1K57d2YinjF2lPBZy0giCKj86zhpDQIOErSxCGD4udc04NSyLK9Zbs9
qcIuMG2i8u0yj31NtYl6Y+5A1XaAKzPvrf1oykkNV2Dfcgvu+kr1AGiLESW0GxG6
pB/U9XNuK4gUFYBmS5GIWk5JrmoZUHYyo4z1Ci9kfq8UU5u/vPLZotNkM/5vpoZf
ucqOnn9lkb0CppYFuUfkE5FebNvAEvPrJScoKG/hVUnIzkx5nt9bUTVIv9ZMLYwi
Ak+jPQmrwuz5VLFDrNACqHe5Ki/uWCitVp2vg+6d60/edp2d1Uu1ohPfK+5x00v6
CdkaDSQ+YWt46aFkGMlAh1oqEwcMNlvGqsUiiYvFgecpcLHQLsj12GpxF2CgjRlc
pIJOKh3Q2xJAtKJ4CPXaAiZVMd/ZHVaXwcFi6SGna1B0eA1h1foX8D4kmEc9y33Z
cRVJPGUyu/zHpudDTlJaZUwwqLQMbUxrzQAJG9GLJkJ3Xm7hD0QwDU1reF/TDMUc
+HX9WQAr1/hDmlLdM3bpGOKIlitnFPcL1KSdM5qLfk3Hf+h7uLCwSDE7m/WF1Ryn
/mg+kgNlPN4yuIdHY9AWoiL3v66q9kQjiZf0HwVGfamj8Q/H645Rbz0siM4RBkjE
apC1oJ+7O7T6BWYWJN3H2cFaRsKXI2x60g3l/wjuXVNVdJCdFcBKhxQvNKDhAW0G
veSWmlE6gry6WcJzzqKc0PPpYhwwIP/HaZXn1ekXbMbR4nvrjpwFX/TX4JtTFpqb
4anaA+n46Tl6eV2qcbvnkQ1qxJVCx6+gcGot4bNimadFy+jc1p1EYGQCnJztT1K+
5cIxz5w0dtDDlRVIw/x9a+arp5Jsw6aItFOmj9ezszD+Bq06PpzJ37lnPmGcWSAE
+D1ezCbLS8bfKikEvOp1J9zRWrz2wE2aAaPJMpHA32zarFzJ9zRdzM4pRQyJxvot
dP9fvxblQiKuEGj4FX+pEFnZVPjC2hGcnGIYEqrzZbVip1ocEmfh8Q0UNfOaojSs
RiTrNsriGtr06Mx5RGS7OgoILLQJZY8GSZIC4G8iQ35iRCxXDeia4jwfM0lAWWU4
MRj2xW82x0VCmK48nBpl7Pd0jFBfQG8xRU4Z+QWMniiGnZcA55oxAm+ahwqaGkkA
VupbEt3PppuTu069tXwPjQlaZWIE/2S2ibsF9DJrPCA=
`protect END_PROTECTED
