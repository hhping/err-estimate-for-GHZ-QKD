`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U3BN9qn7NG7jUOo0hRuqEDtUdXWnaYZfPSVuRcIZdz+EJ8a0tVcJSnefkv/ddRia
B2wX/quT96QFEX01p53l0shFeB6KcbH6wsTiivOdFm2FhERrtF/OKa7d4JaFDoU2
mG3V9+W+SvRv5vMfJiDGe2Zf8btRFYKov8nEgjzx+c2wxUYETS9ag1gvACBs1puG
jS+jcbHv5BlQKloVHE74Kf1YMF3GF9/PEy8bgQ+gK7Y1+363lT/sEiNV+ApAkCTc
R1NzjKO+gIC/2I3dbyHlliwnOvTtfP3LD+ssnffp80rDSqW2/B7q+BU3K5TRTwH/
kTwRSG9HQ7WllFwSutnNXq6E33eSNzX48ZT1rzQ1FbxwKbnkLJfXyYnZPYkh/uce
khPuHg3EV2/jbxNXl/wPYaP4XYhF8wYt4i2gymeEPMxxteriEz9z37u5qOHteHVh
+7z1QM+vAuIdLeLQm6ZadyVOMEpyFN8MIku9XuzGi3Rcs28IaDt/hSyHvScbfFjH
msE2bpBVAID3b/bMeL/ApBBmKOGyUQOXOF9Dmg9/js7Gcx57UR1tYj2f9UwIv/r+
jQKbFPjpY5E5dEMsmUU0O1CXm3G6O4p+kwoNK97n08/CL0urLRG7GXvUGtilA8mT
8fNsXPj+OEK3MvEQqjzRBnDbbNOGUbdGxFm6CJmIaBrIRPzMgLwoOmcAbhQguXbI
AynZ8R+wraurM2yVnJdJzs84TMEckCj+DUPfJ8pFebgraGYC7E8Jh2mDOi00Vgv/
KjXSke6mVjXtVJELVGcKa8qpeRBM2zjgM5EWZpfLTN4Axca5tFcLGHaHAK2U28OL
KFuRwRRIFITvIc/6ogWl3dhxvgojNWlZne/0AdZDi0D+D31H3oP00+u9DnaNbGS9
elWyq4ZqPuxNC6Ypj1bCwVszb9gmqj9pSXuX/fWaSEoOj1CQRhfU82PU0/7bG/GL
uePtgChsoZSV4wfMu0MeiD90/h/ueyldew4e+JVfqvdMWljJIOi/edKZs8MDuyGz
JfCQqyQDc9KNqDwOuHwBZIxUz57Xusp18VxKaktH5EU=
`protect END_PROTECTED
