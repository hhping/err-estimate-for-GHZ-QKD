`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KBUnBQQFBa6w/VCQkqVcCFjCSbNfk0BRZtF0bmNHJAC+mqf0SgUocec3BEaeYSqW
n9t7ybNaCl/p3R9A39AqAP6XyWCnGB862MofjWZb5Jv/rzB5b3N7g/1rNBXSY46m
0dovtsU4CG6nxeD9UlBRPx7FQdoh4+6auJ6ds4WaEH1Yi8/pm3XWtg5eHH5k9egO
v+7ZQZdnFq6t6lohUwj4L7Rm+GCX3WklWuwZkCR5kYIL2wtRGFZxOG+GQKpTj/0J
Yv7h7k0VLQvs4I44HREbKAh4q2VuoMqUO2liXs/BVC/Ki7kwkfh3o+fKzXBcN0I5
6Z9ikJNdBIdf12HHYPdKKt//wNz0qfJ+FQB9HZOTXoNMvZg0yMq15wIJsjerVeQI
ChQuk0/eNa+EbyB+Bzj4XpGVKkDdiLQMfZf6W+iVR8QX922z55+fCrpbvjJqWnYf
CbsObFYLCaAvTZa7djZ67QKj8tN2NYBXXxt6N/SuJZBWQ7BHlCCDFrgdAmWe/QY8
4FVNo08kOLxI5emag95r3YnPkrHi18QZzrPJd6psn0pTk89MdGbFQd2EsEQXaDLm
AAS9bUguB7Ki6psTJ4XmIEFjyDNQjl+wR5YBEvydKKTtsm2rVFvIG2HGpnCwoQxg
e5HUl8I9A+kOawQN/LkSzsmMc5UMAwQFa0AsdONca7GehzoXsbpAWbV1CCjFViax
Ic9rxeXyzQRAmoi8Bs7ScU1Pg1tcPmMVLsLPlI1Y8FevxE0Sftwsc3uZZ6hUvsnU
6T7+reb1/nZVVpgE45xxaCwrq7Fzp4h+EcC8JC8q/sK5O2N7pjRKpMziR3cB5apd
TRDf/DV86zHPn7KORc13+DPXHHGp2rv79BdcrU/mehR2a4i4K9fOjEszCfBqV2CS
ry/ygiJg48ekIcAcAxjdxP6MeWJk2TxwCcif8VXLeO7AjjuoQn/EJzM6qKYWqLYi
juq4cglstud6C2cQTqPI8JT7v11KtI+63QHeljHdqyiCkx2d4E7pRB7cKm3qNkri
nd6wYpSLLtVZmsmySlMy1v6sFGtT8yA2DGvIWj6rWshvb84d3vE/5h/VX5QWw1yu
bJy2sqYc66fpCARz3GLlPZ2QaXaF2JcE+MlqX2Bsbd1BBKMFJWCSuMF3eeQSBRMc
gasHhppU1RqaJf6rzd9lkkLlF/LqCbwT1Onx8m8tO1gLAOuW0mXgJLXmsoLSj+U3
6lVvx/Dn/6cWP7qhy62NqWqFDj3dhSp3nVPsXoNkP53yQLN2xNi15JmN4/mEpm/F
lch99U36X5nR9lhYNiWFEYXQD0aTdJb8ab+wJhY9t0smIkbCfB+ev9c5Ho3uVybV
3K5K3dGovS4MIfTcIXDz3VjCOaU7vZGYK+yS8Wv3wBoIosgc+q7ekZcc708swkcV
ylizDkcC4uT6X8qFKNjuh47DqOjZzrqbw4izg+93DKwSeKAnrVQokWv32PZFB9Ve
782juky+J0QuzNimZhbkFcmtp1ulzjAHzkQlb7Hy4QcTmKvzH2IA8kASSNFdOUtN
x1nBTPllFqpxYuMmxLNyHOgalh9+0npNzXnHUqgNLqQtCwFPj+3w+lito2JvheWH
5it7ToERZYuij+S0q46fOEkFA2cqKniESIkKD3Hvk4+tWdJLia39WNaLczU3I1JB
S8VV0t/FJNTp0TrhU2DSca2Ka8iWWBj8W7yUoCUd51wOeMzyAdJF0W5GCB7Y5EiV
t53U1AxyV3eonrb0mB52hGtsfhltCYa3vwv7jwx2ydmyKzyUGSBcjye4nzkOGI+k
eYcdO4j+SaJ9q4djF9G9Fpx+6S48HZtvrmInKrzcb2Rk0k+uvMXUfaKMmq95mq8U
f/6w/JEBhK/HIfo+p8UXTCQUiD6ATdZFG37iE7l7UpVzR7wNYBh1BFBnw1cXX6ds
gA7B4FEQl9MXOyDwzZywfduJEBO7pFQbLZUxMeI3Bxgu7KBKmkDJ8iwuSVtM6i2N
sU6o0K3TG13Oy5qKnHjKQzkYRXcaUD1n8hLIydTX65cCnr+HA1LBvdoDqXOXNvhM
RK4JXMryaDCefW6DFPUEHZj1+rSwAK1lK+c3E9lQwq5mZkcIdBZMoz2aj1lq0rzu
N1YgtDkU6t9QTk3Lr70QdV0Mf4ZVolWPGRIiRP4l0+p8u7TqM0WaNhjFwr9y/nqw
N3cCGYwAPHaNjZfIKszhuJpTPk50BDUqLRT0Lz84dGqkyL53J8V4hiLaB5wjbcHv
6cYRJ7hGFNe+OoGyqd7ZfnsuN6EySDM8vQIJP3PTGCIB7jcc9UAJBg1Q/Qne7OQh
X60NE1zPjf5Na/VLPr4Ex18vqNd0gOXR8cPccrQtiyak7U4Fw2hc9NAFhaw6Kz5N
bGxBvg1fiAV6pvxwp4a4WreUQ5tGxYxe0u7JSbZZrhjscsuNkeHafPRpxDhjTqW5
BwTWwMdo9mhpn7+Sh6vrBe6pwd69U8zD5hGN7SceVYtpqKm+z5vjnh9mSFvtYhgP
Yr0TNfJmb7ZFl49R7qMlrg4E+gyaI1SBzUMaYYEW15DbxO2HSpkvvezXhD3cl9LF
6tpxvI+toKE1zQVYuq3uO0UHo/rk37TxIa9OUn40McPWy14T4h1JydPqGpTMGfOP
s8/ijowvocDDtBT9nO5xWP0FjIWRbcYkYCkh/VD25HQBNaHsxvf+ZSgFwzKDrEGq
75gO1L7ed6Nt4o3/79eXFaOvKoSae6//AtuUea5VpSuFUes3A9ilYXh9K5guK3vV
tJLoh8xmLmEs1IKkUfNllomnCCCYerjuV6oGr78TcVwZfQx/SeNrr+ePmSkrBNI1
eHRAX4kQtiIo4f1TiCXqnxZAZWtUzh4it1pnp8u+bLUr+vi6AkesSb57tnhwT0+8
ELazU0FnP2mqY/qzdornuX1KNw2cSZQkl96HmYiys/JIfHdQQC5nvwCYojxAz+fc
obHEDl9tfmFSG/wEY6lZ/1H2hgpWgjw40WXpaNPmFkxWXnKuYlrX9MLvlvhaeJzs
VIa/i1XfMMOB+QKAX6rh9Z4RYeC5GSd9V9WtI8A8JHkz646EXjQFtxNYDh7tbHpv
NWI/DbkRF7wk2KHmjJI0xktAORwaVt63xhxcVcxYR110ecINBitbnzmS4oZD9Cv+
SxjQ9kembU0W15V3J0OmBINhcu41kZ1Gy7Zq+ESj/P9AV3XGJ8IpwrzeFXTNzHPu
LxzU5+7gfJPmCapKDxo61RqEZ3bgVCtXRfrL364OXuNfWvrG/5tXZNSbaUIlQ+qr
XTBXejYp0WvyFCuqRcP4zfGmBAQXlt+wGlOHozcTfo1pUR695/7kQ/v7f9IYUQrM
Wzwn/4Ylt7KJdRu2OSZ5PiyKf2YrK6swF1z4xKmWBBpzuleav0D8TZ+24jIx0bhI
/17udv0Z2VTyc9ukhwgl+D1wsWfeTappzYHtV6gOP2H2qScU1DlBBcCeI2OYArtw
/yiiaM79GNG4q9fsJOjAj6AIWvZBbt4bTws7yoxgMg8yEACWq2or0AiByfq4X4eT
zMCr/+CbHGvvlsIlBkBS2538k680I4YGTePJnmhwUtJUhCTclu5HqQNdN0yA5vJy
8UF6qBtljcI8Z3WJBmwZZGdN1vlSy7hxeWfba+IgaQK2h8AlZNn8bBMhTqd1G4/X
IXudQwfKay85Vnmi1YowtjwOknUdZhDuR4voOQGs1D5BBGAeQGLHEVsp3cF/dabP
/y0OLu9bYZ+wRQwIAAeSdpHcWalQLLDbVH6rDphxct27g3k6p6gtIY8zLmJP5Y1z
TOaSLgcEndyxFzUOhBzTHsI10k6p7qzm/ydRqTPUHRuJXXjIGVtv9ochW0yJsB4r
3g3pPadeawr5VcC8d00UFMSOXNIELQNdXmudLxcI4j9qEzQgw2RDCv6BWLjtAyqd
6ltrgREM1R8i5XE4UlIqXZwT0IaisdvFsq1c2nKSWYpqgAlaShR9Iv/DqtP6pbiD
1yImgIdSpivLRzgIhc30QKUS45rxBhRvXuDvNH24XK6uuTa6lIH9BTzp6ye64LsG
Y14juw4557cWqBW/B7IwBPlanaGZLIPnU/LI7GqAkRBNIkdXPcDx6lVXy3uUCFp7
PBAQUFGXt35pTF6bmV5UvwzJzHqWIt/1NYPX7JtYDHTFaxlqp35kKRxBMQr+4fvh
tKXorXuWSTzotNOWVB5le+t1L0X9sE3kWszDkN0jeYpVv35xVRKYvPqkYLvj6bfQ
kMIQG2u/jrF7Plb5sz5eBCmXG4aySciutPZCw+VBdQvx/zGMfmPi9GQHh9YLQmQn
Z6rUb7GItUlcr2OHkO6et40nbkl9Omyz6kcaj8JlTgseJzuSnILjdgBqFl6T3NPB
Rjy0XapDVuFiBu6kf/DD3k5Rn6tRixuAPjLH6ilXL8E4mOv9mpnh5ihQmuyQZNoV
FNq+eTRVFQ3bQPU2Ss3MIh/zmqkqxXQyhH+yYVAomk/M0+IutM6vP7b3AUU4Z8+6
FCHz6DHciL4tlXtk7UTCYc82hO4uOowGqPA+cJqkdSNNRJ6i8lcYzkNi0CfSrLKr
UPWGybNXNoiKgyLQ2XgNk4ZL4vMF2FQLc8v+rtY27a+RaxVHGc93OFiy2EeiEJwd
R9Og+3jC4Y8UpSsHgXK8v171c6NzxUvvKUlwibvx2/y+W43bq3YouSSadB0W7XXB
8wgaMFxBVCiyqrEFccCY02HHTCnocY4Maoqef/gpBb5UNU+vNoRSku72OheySfpP
7EUtzM3sd3c/BxPRSMZiYMjZUub7AcEbNI/RkgIljgo+vm4BibjJ0/fo6DuIXqyk
F+fLPESJnpfOVg2VdvGs0cqAHj107KBALPQUTUj3tTWTosHM/+yNYWpHqRU1AreF
Zan1EUy+wb94V5Jlf2qUl4ljDGzZDZ8WgMHJC1di/Rs3BWcrDPZXAtcHPC5i3r+O
NczdtaZnFRPaVdEJ77XnBc/RM/VtV0JGjJhVrjp9c1naYugIdA1Ha01KyloTzesN
uvi3jVlEMmUOa/JFFa6HkXpvF/G631M7tDbnP2hjOE7P74n9jheM6mreY3aenyba
zviETb3L43PG5FukiXzqkYd/8Cl6erUp67sTHBuojZKOU7F+rry7zzG7jVS7VZyj
4Ax+JJrDC/DecnYYeEuVxA==
`protect END_PROTECTED
