`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ohP75D/hqe2z8vheYCW/4WmPYoB8RcallgtNudWN/RlsSdSrJWF++TG39HM4pVBD
xvwi8uXJT3tZnUkoyAqpli22OIkUNh1VltXBgmDJo7sOYTx9L37MSTq9yhxI6Ua3
bd4we67NSDgxVJCJ+Do5YqubLEXAS3L3/gw1zUWrrHJ62LxOTgo9DLnUw6I5wVVe
d26tfSOzow93Sr+jPWpYwQRoxtBZ1PRXatyRQuaL+YAn+HWilyEiDVv9kr4jAdHU
3sLNWPLrANLVgjEGAMXlc0FRjJ5C5QcYTd5xCtlwisCxQ5mfy7RHGDfiW4vdn3oo
wG8o9/q0WIdFoAFLiqbDbvjBRS2hxZlWHOfVFqikvrcWCuCqUG5Cxzn9vWBtZHl3
cncD+hub3opYqCFMjhOWLxtjCcROEFtmNNTBRd2CwkDJIahqx2s1DxNrcmmNbGEi
gWV6Wn3ignOWsfxM6DqOXT1C0DtzrADAJ+iyJuFGJA9PYXnrV+z/CnOaWalTArWs
SjPUVx37VGfPTtRS25y9eU4fV4YfTnBavpq1002KnfzmaMf1q4e4h4EVFVw1OIXk
HkzaOjEOuVjYQwhF7uptbqM6ym0rk07Q66VYCGvu8CsuXMWtcXqbFb+7wrGxnROb
nKMZjZc+JPyMuqqqur2JMl5LEkZl7CRWWP/Fofwn4gXn3VSna9JMkSxfKhuRxtpd
ZWrwYWZyfrLKHFIs6rMSQRPk4xgxLn2nVLWTau+XtfoiSS+t4iC2HtW8zIM2pXno
xwlkKpPPPbFfb6sdJcrPYKK6Pw9/Ep6zpfZ1FPoWWvj5LaP7ItfIT08QNEhfOHO+
KVl5Z5ye+meGk4bR3E7gr7c6/WknWlj01sVFxaJhWmKFDSSVt0sC6sewXQ7u9HHR
eAha3nDKX2tzVRjet1g6Sg==
`protect END_PROTECTED
