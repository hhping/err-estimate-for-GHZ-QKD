`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vuUjtDqofqhIDj67jDKB3MbA+faKqqyh0b8Wl66UsSXR9QFf7j0IxeHvSBRFKeUr
SWVMf1v7k+fX3GdgPC4lH2riLMB72oFyuIhWbyOjDNicCLMeiSaUybQUkcaTaNiU
GRQOBjuYsyTuSuFuq76nR87XcLexyMWgW5rOXW0LMTR/dajlieV11aCOcUOtD8FP
Lx/5owiS4mjNo39k3Qets/sQ+45puA4Ak7PSvCZsJ91H69CQK0TpUfV7pDGWf0/M
P+y+mcxaaH9dAxu5hjyzjfCMwx2e5t7Go4F6E9AkBWQ9r1VBg5i1Pi1lCA0I61Qx
FoQ7fJQtZluQMlvfnvFEIyw0zD+xeDOxHeyu4a7IwsvD5LczUiOwIlqZ5ZMGOwcZ
a8awUvxQA5Lbnk5zcLeZWwRjqlUtaqsJMYZAh/VmDRoVw9MCu5Xj9NTXxCl+EnCJ
WaMgad3KuCaPFFFXGK7a1RXlSzRk2a6mB1X/uG0psqk3qoDTSeuZ4mn5sJAKyy9+
X1mpgmPEtNYbEuVsq6wKx35gB36S5jnURgI87H3lq8SCcp5D5MLVr8+/BNBbkMID
AUfYC3yI388FxYmFeDVy300nrhN9sday9AhjoZp4oiOdPL0DF26mPoJnZM5L5Est
RzXcJ6n3dhBRFC8XMQpYkK22ewzFNagiv0zELo+R+FEz/1qLnaFJUDOj8u8tO+Zd
7nUhO9GsnbFIjy41AgQyZF1YrXF5Zt1JfUeCpnehlLG0yD6wKsNS4QgfPuaIrnHj
LOhXZGLLicJl6QGcxrAgBxOWdC+zxTHikCmHgOiwYyQIws+NqTy4S+NNt/LR81Mq
qGgfnMKtsEaBWA7m/TWWDu3spmP+wfS+QDivmEZr0J7TiJNpdCCUyTYvTyh73lk8
m46x5UFhREcl3DrIiktWYb2I+4ditYSZkUYBt8K5S8rlt8u0ysxn/1Lewk4V4qir
wGN9VemfrgXiC6V6qGqnF5y2FTwvPkvO5qC+V+EmISO4ZelVf+nw150FJMPkW3SI
`protect END_PROTECTED
