`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3WIYXre91DKdCVD8RQsrJ9K4AzogsmiBwsZETOxC1T3pzx+1zu+P+tW3DRtlvfBJ
WdassNUhuk6fc/HBfq3UhxthAvmtoNeLs9VJJmW0QaNEA4+z8EMYGny53x+YLctQ
VrA9eCxwjEavLQF/YjoMmLiJKLHK4Qutx7fsieJuRigxxHMYrE2ROb/MRpmKxhL6
vYyRbBPi2WCV6ITfeFQKd4ZPqN+BEstmV034qOyqvi7/BV6UHXgUWpYfkCvtsAU+
xEmDV1geABibFtcI8rJCLLmmQ9qVSZY8a0H6l2qN1XE28meXMTJ1DBXMfomYsg2x
9q7txMl6iVlMWgPPTJ/HI8Q/L2OtkQuphY05ndKSJowmcxp6wVmxrFHoS99NrBFP
ST8UxK9hY+LzxQZ36P7E4mV4i+ZyIj6SOvrRi7lsM8E=
`protect END_PROTECTED
