`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jZ4k3tolH+LftAMWbloxmgey31biHy/nyrn1EvlGkP32eNMETEWJtYNjFNSElfEf
ttn1fd7Q/QgsarKQQUbV33MM1rUXJ9FbMt0Jon21L4bOt+GGGqzqNuS7qw4JAnGH
J6pUmFU0Hx0c1OKmKCYz/Wf13PzJNKvI3qqpG8ok1t5jJYBQwfLCeDRh33vXPXAZ
++52WFuWkdhD4RUaj9RjXPHjWPVjbeLALPMsYNrfycZK6gOf0Qg6/c8Ih3Zwz6X+
f4tbCtihnoo2HRCOgY985HCB9cGgJkoQoOBMB6bY0yPnGajFc2836+KQ4yZHn7IR
kgY8jXGGLihDtM+k69zOCGK3LFkr2/OGyudV7FSnVAhyimp9ufA4VJjwaB1ZFfEt
fU0rovEmYMC2ZEMftUsBYfLSGPm32YUY5La59+e2IboRtmVKwmmgTkwJUxLWspq4
tynmtW6FvYU2JL8wGZAG3IMPlksT2PIhiNrmIiAbqnYDAnp+usecIRdhcR0ukHg7
IlBQq4kb79zCkP5uG3JfBACjjYqPsMjm6UYFThl/VMzhPqeHus4B/0X6J09KiOre
GcIVLfHotw2LHxp1gUU/JrFxZGTvR4u4l9dATHT1fW3cdbI7jRkgAgfdDU+w8d8h
r68vJO1oG/GUaTAzSiWQiPtxZ2UCWzO0giWk3o0auao/BtduV09E5w6lAPvgZR+N
N/C1Wltug/QgqWJTPrL773f9WnJ6mtLBMShnKlfj0oP/f8G+F4bNULINhI95mVka
J/7catPEMFGGApNywnJkUJ9FhLHdqTqYeUUKs7Huyu9vQIClb+Swj2YgU86tLx69
y+6JDmt4vAd+pvA25uzMASm9JIirNxj5RoWEjbQgHbpYbXCLt35Um0pIv7wdpPPe
u3DhM0cYdGUCLQOJbr/T9pGxRZe3cqx0dCOLFjWoY0vXi79lyHgeC7DVU9yWynBU
o+nQICVpv2ofC+JNuUqXygByxDDAKTbOdu+bDyJKhLp3CJ09MOiuD6HUpsqgvtbp
JhmoYGJm140ZXQnOTzaz51a8mhTEN71iYQtj2WWgaG1PW/l4AmUxNJzmSDDCW60k
TgrP7cJaPxadRCKLuzE0+jhnxyz6OknMHzmdvw1g6QVZ5ryJ2ihyUPwRtmJ9E7vt
Q+eN/Kyo12dWh/Ie0umBT5xRDtTH3gRYuJeDlWuJP9cwEgO88TaS7N2L0L6lt8qG
RaZmx+fggSHDZphDHVaihXvJHYPWjXJkcK3bjoP8rkHn0XM1HhQA6gy6r09exnS4
s6iTlwjNby4QfnEPW8TUjsnI/thMxEDBdbHdvhsOhwO8x5mMTypl0qYR970SKgbB
`protect END_PROTECTED
