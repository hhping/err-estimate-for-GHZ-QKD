`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JGi9hbxU9TFYyDhx+l8ErSDnGwAmrDpZoIQGtaL9AP5Bp02/ewEchQU9ZghfdNN+
4BMaZDUL7zyrxSmyFYoR6urVuPVLWWsnfi6/dvEoU/0YKAYsxTYm6qSLyCYfankz
eLY/+k6AEzAgfofJPZTtDn/Ouq3w7dxDZgULu8gU53yqKq53GT7tAf3t9JiBkRTC
9oWpgadvpUh4QgpucoVMig/HGNpn3w7zh6ks/gOfGqb+Mr1BWEoKuNvMeScCIeAh
rvvpMChPKziVOi2uknw7MdsYsVGiSCwBFnEAl3bol/QagDq29uadEZRMo2jyiPaM
aG1r8wHC/bXlTjWomlQAreV+jztrn/jDe6FASISlzrCH8KJxQD4JrYUJvvLFw7sR
OCuDtS/HzSr5g2VlXqNqxOXJw+86NVcUE+Iuoj0Ib1U3Z1TExgMKNGMHOkpk02jG
ssEknUeYiW4dmTaFplEvuT1gJmScdP8ji3XM0gubavVRft4eA+UmNVB+Hl1zwf+u
tXxuSz5vxmLK+LXPCRCQmz9Ehbh6ky2dHk7EKzPBNfTznqWB9H3JHnRobQUc2Os+
mVHxuxqUjPGZoczWOJsUonIo/yaaDNaL6edVi5lg5ZI=
`protect END_PROTECTED
