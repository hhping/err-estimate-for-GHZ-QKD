`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NErvdEo/yiyYZdDirPjBuoxqfEb6vZPFhh/w5dcozT2iWHfVDuTdW0WnXrHF/11v
II7cC/6hikkVRczqu0Y1y73aZnVpPEQOKJsSZ618CHlh4XPvzCV1A3lyEMGqb89b
pmOh/5awD3Z8yz3zILTadW5RRY6J42CAFNdLaeDbSx2ZvJrJtw/j/VqNomKljBsd
XU2BfKOMbNjtqHi2Rv6GPKSBvBKbCzBs56iH5tMZ4qJLTFAYr3G3J2aQTAJVDLLh
O/zMoGjb1jD39RRcFNn/dzw9OSYC/LZ4n0b9IB2RS7cmQ8GuHVgZMrYR9Zd8Sltq
gZPtaHU+IL1fHA8/PkywUhkhndEVI7r/0LGeNwVkugWJQmfwQbjYLizKmq+wCOKa
/6RytjRh7SP+dZQFJA208MtXVuH0BoE5Av/dK/jFy6LZWbz3lUIycoaLhbuuhis1
TDBkebCUQL5YVyotBaNLXmOSz7NwhD0xfeSVT5qKfsBkOk5jbGHwdc/8b/oUq+KE
VjbWhMOuZVfydID/y9KQD2OrG1D4gYNTZC3+T/0mpvCtE//ra72vXmwbSzW6xY51
zw2ldEtyKi+w9TiX1RFpiLJfgNpxJfEVdBqEMc9oJqAx92kzPGJBL5mrUg2qLXlJ
8iDyOQbH/soSa9Vxjp4yjNY3YDSQjbMU8oEQJCFRr0qcDaRKiWIqqdKPwbL9uItR
paRzEXfljYzDe/TYpV/apPDoRzrzZt8AjzkvamGuuwBdENjr3wBENWti/MnJkL4S
Uk8hMFCeh5tDroE0TGGRMjTiAUN0wuqqeGGFPXDYeqslWQE2CQVloyVeVFpApM7F
PvOCOnFshvNt2L5Ylw0IZCpc6B+cpRMkRcgDRcQ6YU9S3IDyq+qy27IY7P+WSbOI
VnOnL881GBUvkdzzRPEXFcFyFvYGpGqNF5KCrLGG0OdtljPcrSBRt/o22epCLYK5
xoo+jOLWUkGC/FwxG8E105TuwTU+s5sLC2VjbqNfzsWLl32/QQLqA9EbFY2hKF1N
3Ih2EC+N6Z9f6/woDBTf2Mmbf+LVwksOt/oNOKv9uhI=
`protect END_PROTECTED
