`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QLxfiia4nNYZ3nmXg+5gx8NZ7gyYcixzS30/gd3MJSDmU9EKeqVWfuOC95SKj8Ip
Ah8XyAEETHE0xK3oPoZApcM8GQaiWSFmtdzaUNBGrv9qRnxn9Jlnd5Q6q2iAZYR/
cHrshnRVcbHMZ1JoG/+G/ei5djQ973wMEQIXLOoON0ULa2PKXvOBWv+rEd4Q+aSr
Q3YFmt9PLSKudBamLGcPHeAepExZETSIK34HlZcXhWwHw9vobgoNSFy9mvRgxS7k
ZTeWrw/Y0fFFE5HgaZC7xf2PfNjkIY7HyiZncmLE5ixuKye0ozoe4E1/Zq+wphBt
ZikQBFfD38RpI7lX0iYpptDnS5sAY0Ar3b0hFEGR3c1HWOixR3eqjcNaMEqjNGGT
XQFKaz3xRr4Tfua1MRdIaiG0mQxLIZvJgvHoa57mGLJJnY2mFYKdBnOoh2IbKi0W
EZmaWqPaxkCW3Pc4bb61Ag4b0E88jrdC6+5heI57HVFPyX/u0of6wte4nYHF/T3X
5qj+EWHnBXop0l3HyD0uBceEYOvgh6mNfAtvEyaUdVF4ICfyluCAJh24JGVnfql9
psJuRB35ursgNh/NKUDs0nlkPB5sX6sXCN+8wymfelK4xlEMx2Ad5Nr6tju6+AeM
5CCrjle9/Hrqp/h3nK//tMGHxXzcr+tWP13yT/2EaLqqxnV9A390rdAkMP3+/V6R
vQ67Cn8b7uz/t4YINJdrZo9ZrEBBEpF0a8sF59eu9PkOw3PD5smCdccRbyb7L1uK
/Y5nlsrHSLVel0yMpFbDhquywwke5DylnK7nd6PwoKoiRsXtXZ4wMis4XC2fOx1U
mkYt5p8rC/uKGKfYK6FmGexizpS9gSoFaC5jqoK/dyQ=
`protect END_PROTECTED
