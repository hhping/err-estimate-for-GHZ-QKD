`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DjQ5M/wRdEpR2F2OJQSoIkM1GMxVHbgHlkMsB0P/9YwAMBOSZiUK7htNZKAz92po
JNiN+QeBdzHzgPGZr1RCQ+eiz8IyIBBGkf1Gc+Qetukgh4J6ln3HyKEVF4FTNZ+F
mbx2edTZ0E4c+CiYMR0x6P+GImTJpYkpoWcin0u6kXN6EEG3eMJVhU91G04fDc+Z
jm7jQY7kmMlPx7dd6NA7bTsUE/5Hodr4wMz2ZQ7B4dKxKmmz+dUIhlIrTFjdYbhA
ENqtt2FOel89vsJivL9CQMkU4zFySn/148UVefnyShqqXpw9rt3F2o5Svg9Qw5Xu
ia7DkvOGzCHx6Vgp8sJSGAeBNYbjCI5BT/w2dSclKJuNTp4axrjJkdhu47/fVrfK
e27opOWwucuK50n67/tB/tOYm0Pe/Uvn/lygHf+sxMjjT52nhSC/kk/fc+uJBRGA
6VJfkboQ9oaM8Z+x7sAksruWFYxjNeP+rvHLTlMBBz478Tfk2CxbAlV4yj1+HV2B
5yUmFGycsh8uBS1mW0YVsuRDEVaWven4EwRpoOGYt+HOpUK/gevZaaJOr1ZsJfNP
Bj7kb1ZlPjX6ObyLVX+HHsvuk8Q4i4KwJ3deC24aVT5BB9oKS7ZWmhnRgo/4xVj+
P/T4KpqU8oUsat7TVv7inyLDmO0SsD3Hb4h6Bw/4xYc/y7yV+W/UwmgA1LnF/OwW
G4yzejgKudBsUSQGcFK87/avPlrv54S3KGUI9ZlHXWuG83I56pcp16zdcXrkQFvD
aB/1KYxH+sS9NcbDF9VMJGR5m9nP8I9p02gm8L62lFrIN+nyIxOu5IfpVqh/pDrj
0gX+r4S2WLZ5Mgn/yTFmZuX2f+ZtUV5W1RYGmvcbW16h17U5GQP2EQ1PUw6vXBDd
oaXFTB48vZLSzy8PuZOfsEycw+R82d9aEx1LtklKxUEiuLLoRAG1kci3/wQ6SSvb
zhUJzg//cLITqz8FCGdPvKCyy1DQHi8cfS4Ug0A7SVR807TPL28i1TiOe6zQ3zVu
0S1nUa2HKrtO2PAUGDG+4vRdOqQW7AMAJ1neL7pWKLBzUc2HOrwMFnKEDUvf1y0W
E70LmPhg1EAio3YrrGZ3z5+65rUdhn23G9Yh9dt4oa0hmXvjbv1GCoZoS1o98840
xzDLAwwyIRfNwlNGJLpMea4tOVM3aqn8fjMWzLPTozWFYOTdxrR4PedfJZKNAbAx
KZyGl+/oknmBWRE5gidsOe5FyL9aL7MfWEC2UyJR8XeIYAT4ECw4R6+I8VhWiPxc
mX3zlnDrk58ML1XoB+H6ZTROsPYmULSXGdWxjn7uTR4vxc6eVo5G29Y1VTUXFB21
cytApUX0Wrfy/YnAU4wKGHP3NuSLUvoEofWOKhyf0g0sPeGLBGgAA/sL+06gXPhX
8O8O0JNE7oRJ+/06iiUUEjhMzR1NLWvVVWrWPW61J2YrnVfOUQtcp8zT0xw4KcWe
+8bz/eEB/Eul0wc0b7O4t1Gn+nOoes2kFweW3lLvP8u3YbviU+0h6KPDoAJcw7eU
KrZI2Rqqg8HMECT4aWtdHBKDcyeCDmssggqzVrH1bYuFF2ffZl0qC7lhs5Nhzkhq
fmrxkzEqPVk5op5oMU1Ie8jXzTUHqo5etx+OmGjlT9ayHmmTlTBjWGdPgLJIWT7Q
4QWVPqr5/B/pFmf/OLSUy84Kln5cqW7MA9fhrws9dP+1QEuiVrg6r0l3oJugZNzk
wbn4H2FsmApt5nUlLhfC79tLXdWi98eD1a8QoFrJMsizHaa7aXK6f2SehjWOlxtH
Ets71V2JbaY1/whSVuSJdyV4j/RBpC11+PuoGeJvGbSxJLP07ID5QM4ZNFFz51zS
S/O27xJSOcY7ovDRP6sLTmcHMLt9nAJduXk8XXYlIOW/NGcXhEeSoboDReGr0qk9
ksKouUoX3ya+WmIjCOfVwptSAVeLgt/0eDr30Ao2u+rr3OuMv12L0gykjnEz0LMq
17EVTWNaccpNANmXAAha43HnGa11mV8gR8xIaTSkr7g61j2SGbnVTUclkc8+Kek/
rj7GbbM5uLx3ZF0A30rtvxodHpXsJyBviNn3AvHwBPQhtHFDZd0fnIf5i9a4Rb4e
IfLsuj6WTrcp6UCuc84nugb2lU/eJKx0Sf8ECAWwNUd8aU5qkIdW+UOOueXmUtxs
8TLGAMl4F9K0pPCBEgdHlA2KVYCnmPTa1fLcbWGqb0Wzcuca5Ez/noA2giMz8CAb
tvYu/UZ/pqofXs8nEBLqV9v5qHPYIGp/c1rykDp7eafQe8uxxn1kO1NbtvBPgJ/A
w+o6WDCErA5c20Cr72vzEmvq0UrImOiZGF3cwIWp39cUIs9IbeliyBmyPD0TvHRA
EDC3F1PlEOdHZqd2dVRFiabsVaYgPDxjbtzb8ckxz7y/mj76Q4Vnm2orJSupxImD
Tfsqe0eB5mQ37ZmFmi3mKTK4cDVJO3Q7Ha439y73piqhoOtUj2RwRS2GNiYA/vVS
I7pOSbcfLBqQKS0WbUvuQCnnI97XMD5R4XeSwUQw5h4F2ud7j41xxkpL8ELOhDyX
uTOQCzgv13zOMVo02Gb8Oe46mXxWDyLhw1N8SOjAJZrARMUG3xRfyIKwCi7nZspG
ulAQQT256PfKpODz4sKfiIROHZdQWDv1UDZjmEZJVyOjw/3Qavs2/wKGbciFV9ae
zF5yjjx4zjGWtWHpdGqInKlPPK/VGUSlFXEIVgPo1cju8gblkHk5CfbWgm8pNytQ
jzmYYD4oHmDySFC64dlTLH1Qh+2buhrwwcKYorLDimKBS8KS4zRFguV4v8yHawX5
S4pfQcQ/61THsA04TsfxWWGxO5pd3CxG+32c850V9b8/okXab3tZ5VrkrM0u/YmX
LngkFpbilbUG87xji/APUAZdzCWSbe6M16oUT/CbCprO9xTtq1wslocAwLHKOVGr
nHDAzPLs7w73ko8rBGR7WVwBUlhg99SuA+DP8+tkhW/A4T02+aD/rte63hHlEQB0
LUWeMzp1JOV0fL1YNDGArbnNxmAW/lK3n+MP5g1LSinUh64AeWSGNxerBgvCkcAE
noaPzUapvjU7eRk5MNPOfYm6qZ62Sk7VneG8gYu/QRykBttJpUue1/noT8JGjsSd
uqY3yETqo2CdEjU3+lK4iDG19MzGejjvCEZ9yCweR0GVpYf2dD4VBUChgQDdUKvB
AAmDCga80gHrihwmfp7R7iKyAtXB1lmsbqUwOwGiavOE9nGgw++Q4fsMC9e/KKMy
CINUddDDkfBHwWVgFmpehwCKxc/d5UPHPdRoxTuN1Iw3NNGBBn44qosATM0qjWIA
k5PesFTd7J+hfU1SfS9NWBG4g+Q3x9ajk+Sx8n2+91I0AgucBjzpLGtY5hoskCSc
gE5zIsJV8vIC//R7EoPUjo96K/CTkQvU336qLOc1cU0W90iY6vzE0Ub5SSGfX8K5
ir7iev/R0r5lefGgekGCJkYrNndA44qYw9n8OFm3sxOmgBBHT09fufGqwUn4Cs5k
dLCfyDBnMC5ExVnbBmJalirANNknrRAO1mYHTr8MwUfSCX/qERKiZh1d9ZXbUb33
WaI8vyYBugZEUHj1CLALqNTlisXC9gqZeyrScUEOe/TNHaTXud9Af8JxVZSCk4Dp
NN2kAgHz0xcSKsAO6OJ3TZ8zFDu8LDEcsPMcI1TYdJdpfbJIUmRrzofxiOY+lCpo
YgqKUim7EbXb3vlqhEIYfxpZnPhkE2ah5j60JOUCH8hUe7raFEv2hBt7jcZPsoYl
JVryByUgi5mtKsgXh+WK6GAYEf61LPV6/KeGkKob6bbBxyOTD/gGTOZcYBQkJszb
+2BUugv3IKEOIBSQN/Z7Mqykka70xB+sqgUDTVHCKvE1XpboTqiDPm77eqc1G3VP
dJtrnBmuril0/PIVnA4svnuJtv3weQcpofu2ekKRsMWMMk7qeqmCnqSY0hzPxTFD
tI3zHVdukICIw4ANEDdYcXHnyB6l50vkdVT83upAOzi5wAwI+/72a/YfhdgBgIAU
yz2SStAUxQBLwruc4scEZE8LvTDCgvjRG9QIfmW2WuIPHGwiXNXn2a6SJx/28TZs
dbiSYGrVSeB8BQbAM8P6OJ8QuEwyFhNqHyUrL1cnzN4UFErZKLc/5FHCNOvvS4D6
w15+6nAa2skh1cjb5hYVhWWUGgs4jJlK0xVt3AfdUuMWhqGB2K8qSYpRE/b4sVvY
85DO6alxmL/oKCOP/xWoqTfkKeaUrLiE9csS2lwUDNHEzi4veDz2t8QdJDDQvOeB
8z3g9BsXFQXCEEeKN8Dbe/zuXtWvN2EfJHuy1ORDcUjNEPLmnXca3XKXJiuF04iq
XAHVB42OInrAEVyIypoA6BeM0/KGS3Ba6tMaIutSp21+g8aLUHJXnEWzZa24GxBd
5MkCleIQmguJ3/9nWiG1BHDVFD4BKXEU0RH6JRHMlRzAizaJhsQa4Wdh8NXBcGV4
HQRtWXNI0cbwsYDVNLGR9CAn8R0zhnDsXaj19Bnb0hRZcgCqz19HBOJQvnV37dpS
0Rc+4fl3YqYdh8vgclr4zsncFoVBxspQHs+pRLPgpVBmcxLsafKM6l75cPY/ycSO
A8a/fS8lKHbU2u2+7KociKJJh01SOD9A4bNSit8Cupa7Nr5aPzwhmD74EsVJskJx
ELWbD4ABgSZoUe0eHLaZpI9abtaPMHGwr2iMFCwvD0qZt1AvHBAfE5b0qnUkjIoD
qD/fv2kqzGHf/lYgPVsm1TrZKeaiEUKNiIfEKzO4DLFFp6055YQC/8Bb88NxklCq
JuLOhQVObznv1AHwxylS87BCs0+EMgozeIDEhCvnE1xSCMW2uPJWijasNeymVx2U
ynLbqyrMJtMkDK0KrCBKFM6sWyX8gkFaYkBPlPg9sIAgSBElUDvtr9Y86L8juimF
3DprMq7puZ/nb1eidP7OzvVIk4o06pk4LPAxqbdV24U359rPJ3jPXRcOSIJcNF4L
6zDsS5kNtVwzWel3YzzTe02vyOJS9laDD7CtL5DeTXlKywLeG73DSxjUhimKoBXY
zoJ97m+9lT/7yXy+DMUioNfInuX9/QYkAIN/uI5SmhPd6yW47nSiFrvL2MAET4CP
DUsTXiy3kOHj43asM8fUH4olNf3Ktmt09tFNmsHepg1DN4913wwexuP+FapVPlUe
i7WM1HF1xp9FVgO5e3p0ZsJ42uN/40mB9RiRewjG6Ns410juDH3kWSjOJJMOyXDe
scpz5BnqqZb7aZkC7vS2bMcPP3hFzGfsUSpek9hrc/jJwOwen3GR6aQ+jRrJ6qU6
vxV9rk0nMz8iKrU5QvQk0ulKRC0XwB63FR0Mjy60lwNRaCcSlT+YDN+CdciSZMA/
9I1Z/7WiLMJpW+jpaXdjyf2ELfFJ5POhFAhIRLqMDv+v/Gk3fgQHVl46DIaWGc7U
EoCx0FbnGtCcw8dxY9bvEBFJCwcNRTxZ/Ogoc5gDNbOOG6KrQtxURkc8QrrzsmeP
9XrJE61hh8CvOBZlbpv/DLNZU+ShEF1ivq2xGY/aQmBRHAK/izrZyYQYqjcNZgc/
jqPVDW+U+Nr+iEEbFJetUWeuzqMh8k2WALohxB+GLYITKKzFdgYVQuR9WKUmLP9k
CTgHPFKLEU/gMBlcJ5NLo2Y09dzWL9WlYHdMKBtiGXFMy1oUEGxuBVy5SEObR1MS
kuXvjBU6MVtxQXeJSxxdW4lqSjeGoRzk8BriM6fxpBqXdQe6ysQpa8/+NeoEiKZH
1AJcGkuOtd/3VucCPJh0OwBG+42PBfTHhLtxeJ+Ofm8LfOt4Ce8NwJ2C2VoIfwmH
WjCAb5Q3BLC9IDz/vA/wJxyBotw7rYvbvUNISfcmLZBC9m/MTphf9bbcO3UY3sE2
naSTBhJS691KVRfsj/f+jZsRieE8FHqHXIzD77ObOkf+tJHXC7v16tnB46HBu9Vl
DCTI2CJyfFM6ArXxRkwqAAsudkHVrJlCmsvCXPHCMN34eLoTt5WD+GYxAkLTmbje
U50MfgOjBvM+5Gj0H2k91aGtJTtByB5dl5V1jwGgLezSITTX7524fU37RfG2iT76
tTHKswH7pgJue/PN4Ul9fxtNQ2QAAZS1q52lR4D4fL1S/VBc6YMAHqaz95KQvzeC
HkThG0oG8kT51nbI+LLKTokm+JHlEOI5PZ+BHZYuKxhdsDXaAMYJ4jWwaor/u7QJ
9NEGo0aRxxi9TcSZjhGb70PQYTb1pfBMyh91k9BH6a9gRh+zwCiCdWIklpT8lp7D
lqYnKSBg2DNAcLdyz4MLPek1/8LZ+DX6l6HSN0MRsmJgu4/kVsV7TOrYxgYxzKpk
eVlxzOepQO54S1/5NcnkEKpF0/C/ViXuZW9uCZeWILLDfr1EqbrNPMbhqImXyzaS
zNvy4PowujD1rQzmvfXbzQ==
`protect END_PROTECTED
