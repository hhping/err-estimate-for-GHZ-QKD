`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
emyus8hC/0BdAqGA0tluH5JYN80CJn7P+fOdBCWBTGXA9v9F9yM9nvTmnVna9tdH
G62rPeUO8NJk80bVa6MwKwxezFk/i1CRx3sWviVcgGOqYVsTYxnGHeyi681EPbjW
KHwrgAB9enH5c/TRaoizCrOPdCV887YPZx2ZoUKl/5zpnU2gFnSCTeVqktJIEcu8
GIVAmb4ztoJVNLZ1hHaPYYCwIGUpnek0f+HHDxpJ+VQ=
`protect END_PROTECTED
