`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kbEt6EknDRkWVhgb++nAxZpPyXMh4V7CZNh7fPzK/2Hd6mzzeNN8BHorja6rjAdn
pQXn+ppptjs5mqjX7hh+jJPwoPDm4GYmXYPN/T8TvoTixiyDWYbV11WwNnTsdFfd
5RC0inE3Im0ri4zxqhxmqJrrnInKV/CqoHMLFQn/vJ/cLuHaWU5k5oU2yLV+NuL9
YQqajzvW8vXf0ihhcXwckIdk/GEDLhjuF8tqAoxcTvSvMzxq8ebH0kiAIHWGzfO8
p67MUfICyLubECS3AHP/5tEd7BFdqEmenBljMKWJb0UD2TxgRXxZWf54Ch7nN8t5
WMFtlxjghX0KuKrB++u9dzcxnFpmKGrAJc3zsftk9uaXk/gMduZa2OYyn6igwIVK
CwiKFzDmYtYw+r6X+KtaRE34VjnCbTGQnwxdOoPtoMuaU9p78y/TOV5atYgJDoiS
Eu64+xfwES8h3J9i30E3XfMGmteCd0hhi/eUZ42Q/yOuY3dp/zrDiXt0MJPlOJX8
wCmarHgehp0/lsdeGFC42/x7dWoZNJq1J4bnwy/uegDDqsecHssBoXj6ItILk1tS
0Jigykr/ku4lkFZilWeCeVItVxH38zcCbXaVE0+8+Q/Nivg522gmeV1Q+gzimOdJ
ZsT+Pre+gG9sIv9jXqynFRNjQ+yMSbp2NTyYymRR8+oyVfbGXiY8BBby23OWPM2/
g48eG2z4zoSLarvGrdgezKdqN3pl5sC2eb6xRNAMKVT1Vz4Rp1WRrulth7yHzJ0z
J0+G0j0+fcIF+fmyVfDPtmJUD67Hi34H3jItLiPtQm0xaozDQ6NeUOtxpqPk/TfN
4CjhudY1pk2GAdlLe7b2lxvc0dpnyAbge9wvrs1NZJ1Xf0inEpDnAY16VGFHsxpR
HEekkdXDuj9FOlfAfDrH340X6QR8HU7BARcAIGVr0QlIsa1bjbl+Iz43QdSNxY7+
NfW3D2LdZsYF+LVrKcE1YabDMcnLL/p1zfm7aGEtK/q497JR78dTOMJ3i1jnA2SE
442rYfDJ0D7OIHF5reMH7jdJPmvudaUik5sjv43DQx2HbKBE3KuFFO7Lx5JWXfHp
zsYwCvMjUfo4gimEaVLz4XYn7FFJEoT52u4k8y/sRG8WmrkLqM9zZTr74S0MJP//
54FiIc/2zWN4iOgWbsJdfDp1kVmKhyMU5koSEGA4p8JIhvn+xeGhJtYykiW3WdMd
sAif7i1uDR6oBnwnObx4DD8/s67ylA6mlyOvlSWGPZpbXxaJrAn0c7OfNCf/xURe
vyLr8jBIKtthGHG0omNjgx11VYyJtKHfEv4bKOX+GFvfpP2/x5Q3hWzVpN/7Gvi+
/lW/MFCPXYx5ER7zbDsgo+VOg8QNH3A3PNQiPawIt3fWaleLGhGH8dWuQ2eKRTnp
29A30IletE81mkhinX//OEzn9NIJpVsOTLhTUbl98ahF+C0W/BzpLtvgwsTxF0Kg
Ndb6dAmuSUUgwJUd6wmyTjvy4LWl6FzBuPf/xlV2iEAWv6zasTTkVbNueRYtypee
FAieUlsWsjc85/mtKRhrJv6hC4onrhVEJ/XS0hVuuTuXmH/4UirO/vwQ1Vya8cey
ksymkm40n2lIMMf8ENTv7ewxTzhNtFsO/FHK2z3bdWYh7GqZsD0DJjjFKaGHGOWH
eGnXRlp3l3lmT7+hAJ9LJRQBVsTF3Am5uRjAeoJv0zLq7CxtpNcW8zdmu1RkStuB
C+kkqiz9ZEfaoerIK4jRH6lOJMnJZrjEy2LKVIAaqZWVjJhUC08Z2h0yaGlvBwPp
GcVUKkiDrkXWHng3xw+ZxxUDcFtATRxYp0CkxmHHMLmBv0HwHruqtYzESAxlqPZ3
aUW7S/FnAe2opYHzxmW4giIa1NDkD0HfFHmT9iX6pZ9afRdHJq7ESE83QK9qu/U/
y0WthfS6kkMZQyqSlZzIpQpcKiY2v5iQ7jnVZfkzgALQKfl9gboJN3CeonbEFwnH
8aANIQOMRpLxottiOch6qUD6igfrCVs5Uxh06IGeCfAcjtomxHpJDh4+NnrYvZT2
eGfnS4G0JIRoA+BdJCdVjN8NmmomVkHzjrEADwsuTUYIZHvrq6X9abFHOXY/RS+s
`protect END_PROTECTED
