`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wt9Q/nbcI3XPxC5rFQbl+nmum20HjedZzQactWkMI9FBoZu1ew1lQ08+d09+Z8IQ
qZQxlgwgY4rNNaJvBXseuLecTIPWTIcm8lsFPAB1jKGJAo2/L//RUudGYP5N8lDJ
Bw1KQFfweuhhDThPrQCm68j6prldQmQaEqXH5sXqNdtF5WF+sIhuziUgpTzzQzaf
RZGfunZ1npmFK3TAh3Ht+XOfXYBmGIcXWUZadg8ZrPbmmoTk70kqXoGnTztS2YPL
/PCEPIBexhZ/SzO4DnD7ur+9APyT2nJLWg/AYvqoKrusu5NkyKnjMK1JJ55iZJZK
2w+hipN1ppOtLNejD/+ktL8NNARZHbiawuPS0gSCybliJTOJ/UnZ0DKYtJAE0eIv
et7GpTbEXDFke1lyhtupmbdG4APta292BcRV4gJENab1tRG4n6nFOlXEZq8DxC/P
qTB+ZXeieGptZfsc00Rqa1z2Z+eBA1OFnaSXKwrB91+PccD61LV/fjkuGLBWFPFK
SMis3HfwC2tszTFlwLlDMPPs6JfvXtRwQS0x329veXGFFoMTax9jOdK/8FT34byS
UY1LPF0i2SoCzC5oIzHR6wAe/xQCcJMnKHgn/Cz/AQI+U5nxUv9nIb3gBL/N+iz4
+8N7LaEHl65q4q0lf8PcLwQ2+Fje3KyilPpsKvO3bZkKSipgWa2BpGWYdqIV5VqF
S2WrsZuULu8JHLdRxNjvxs6X6jGGKLsrxUAJgsn9sU24qQpVawCFeKppw8U2XHTi
wPpAu17eXLZz+Nz/yjFjQOzD/uuwJEkGax3gmw35qWNtcpLaIxcOkCJwpUtXIoe6
fAtolkBG3pWyd3Ld7KgJY/mtQ/f9MCr9h+/CigXVAxtBv8pcVjHPkJZFOrGqJEXb
rT0eNS6qSyUKB/MlvK1a01VQXYs3bPkKpVnKDlF52MD0EyW39ffYF1gIYq7lu9kn
D5svLzJ7/BQLf6ZQ49hKTaLExxOgs18L1Kb67JvLc6kAS4cu7h39VgWVArb0TUNR
vjIOGe51sO8Dx5O+2T9hwj2JpT3O/N2Ti0tZqEtXNqbtkcfEySW1Pd7JK3rZljW9
Zsz1RzmmV6+TDZYbUysE6+wHLRzQEtHtI0nFJCwTguR/1HYe1heyAUJl1SzSUf2n
JQIq2fLcVAsgjYtbX++PwO9BxYI2wDnSM5LeSzXPUXFrPWq+q6U/5sFnuObXHP4A
EKhp+vzYQmkFLZ7+LJnvPzRPzXPwgOhwHjybkS0wuTniwvUYQ+GEqv5ou/twYw2o
KPJG5YBKTmshgY7DTiCElZoMchBU5JWvZnfUJh6tpTQn1F36FF5+oHG58Vf9kbcW
duZbv6qsxIlSbNFYl44M0Pl7vT62jmW1OdExYtB6jrYTLuXjfx/CdSw07T4BwB7V
bOnjlcTbHT9vHX+7J3So46IjPp7fnuJLAHIvx1bD7OIRKKVQxWjomZIGJWsTXuls
8a7gpL5AtfB/2xC+PGaf5W0EK5bYRZ2vWzJx5j8f3X7Z6FZTyALqY4S49O//qs1H
My0iKcCyj0YkhmpjtM8n6H0wpzEpJXZ6iKnMiD0SZllTgQyzxjDVf922+Siio63k
jZ+OE14WVSJ/mCc8Xt5gIopu3fljauQyJjoU54VqfQoQ7h+fZJDcduEZ7mbjnX/Y
Bnp31SiW/3z66XUiO9727Pc5rETDwx9t5k6YhfQFCqu5+U2qEwyZ2PK9mPPY8pxW
zF5++t9gK9YFnbSECq3I6r0zb3aXAU9GR/Ls2PQ0cun9HpLxyqCLcWDPEHpkP52b
IRFBDp/9gnJV0tSWbaAbsnD5K/GR/TebnStyidSj54ZkiFREtOlmpgBdf2t0ItmL
RkTO028xOtVEgMr7cECM2syU2oo9AWtMPySb83lhvlByLqNzG9UtywgSTuay5NKO
Kz++/MxgWwiLC+UTUolflTHg7WmLtbujd7c4HFms+8Z1qs5vttmNRfgi8Irv+ZW2
CcWTaAN4CLiokWHMVupSKzu0TLSgNsx7MN1p1hSnz4aLkUi3f8Tx7FYBdxyY0M8S
lloYZYDUjrepyjF249nYZwEJzHk44DlBWNnkkY3GFTyhk6+guoRnMrUb+TBTtVt3
aZL/RlcpkY0xZgj553Vt/VzdG/jUfGO5eMT7++p/4jxLOo/+EkVlSOqa0LgQY+tp
eB3UIOe1AXB/szmHb2ZiW2WJnf6IHDvCcIesspJB3dmsOZgn3zAV0G33LYVzz045
mu/YzADL3+J+Hs084rmLs358DGfNedptyHpgjECZPOkXlNDGCA4HiT72L6oM+eAH
Rg1Yk6BenzPWabUmZu5p4IxHkebDrtPfpfL3xs9hwPf3fC+TxFwb5iC/RUz8PX9T
iScKap5igbgF2Csg5biaGfGUq3am+vPI4ah5/UvEN0KY+idwPJ+ZvIj8IbG/GASP
AniqIdsNLopnD8NWgHIVWlCQlKBgHJ9CK30zxnadQiLA5AOqZIE18dJzZSfzCtSf
ZNca0RqYLXO0AUyOWdk7BYk5ZzcLcAVwnOknV+lk05sc8eYly6stwDM5v1W7zczb
xYhtm4j/KZCTiUIjzrl1mY8yQcjiV7ekQCrLyIXsvJRbV/BgXFJWoCqGqiTepbcP
jgePe2G1wLjllUdtgHobs1GNEqQ1d9h1E/TKE+rB4zgNzI10c6xcLxqmNv0zPWBj
WTDXCbsHpHCb7Cqr6alRVpO7xeNAPZjRnhpAmYivyZ7BSoiVmiE8yCMgSO2e9W0Q
MEy284D9+/vdbnywhFUa2JPUdlnKcCN0TJMDfhWQqlpn6VodBqclvcWfKK5iRB6b
vOi0sEvoBjxFKZOvhyysfE7/yNbQfksJsihoXJ0R8zwtIqS5YUGkCvA+orE7cvw2
K2UU+sa32l7k/E/WvNAUaYmnSUNY26z5w5akgfjLV1byA3dIHvf5PDVaxVubwxeA
IBug2101YHa5ZG02swhSItYDQXhy2Y+xA5E9rdgBdSQThoDnJez7gbgSrbX4VUIU
pwbroOxbycmqYq3JWcv2OzcgDRxez/QYQksiR9icDz+WDWdtPxPxQhyuz1rkiqyO
0iFF1ZG/cEFl5KFCwXggyDXx+I2+roCvIR74j0mhvQVUohiThcGP0HK+2aUB3cUa
vRKutqpqdejeTUhx8bfi1+EoNLloVD5g1VKqz2L6dK+NiwCCeGkb2zqnq7JCwoNq
MZUNiv+Ur8L1eOUkgxBi4PPC9qhq9wTnccgt3YlrD7wHmhGHK+c+K+GcbhSVpJXO
JCBPl8iFM85sQG2Z4MgrtFXxGBQtZzqWnqc+JT3jrM359REs60z+tcNTpcxkC2qO
I2EO0T3mT2YIKmto7aZrUBsJAegwHsjWahiuBGbgYuRUpTa54jKSuzyWI4d1+V68
QP+pmr41jKI52I6AH6K9uTiTnANHKiAFZQCCJWUItOwoJIyeqm7y1yoBF7AytBB/
0TGfwOZBj7Ah25hNy3rXajrx463KlDXxo1O2jxTc+spbWP9y+EJFOKQkkGSH26Nc
PFTu+PjAIZrUF2mXXYAgnJFyZ6fVtFgBAvR3/SeU/64qThyf2kIdWJU0cDCYBuRM
m6oItLylhcCOgja9onJQHHhHP3aKc9NCMYjroB8Jl3b1sOy3mKHeE9sU9IvK4A6q
jgbUisr/Y2EbroYLF5qnERqqhZr7YWzTJ96FaUrVEcUCgo83gh5+/HVdP8VZGlio
JjyayZY5Y8xJBp0v1O6RSZLSPL/Z/Gvw5JHLBX4BOF5jOnGbTAjruEHzisIdbN0h
buJnV8UlveasRMIUKCSXPhsH6XvdXe4XjTI+q6LK9+HYKnRiFTbOQutLilKua6Sz
7aWD9hdsuMHYvYxP1S/FYzUjhEbSmP2cCr4ilJL03cdVugAA0whoXl32BIk0K+BV
gW+r9g7JB1PeHcJFweT55MjvkiloBiqh+MSwahgJrTobthDou2BsyeL3c6OQuVSg
GcDQeFOp+ajOVxj32wkpYevEb9msdLfmn4a2P4SYGLYGJKVocX/cTqGcyhitawOn
cQc9xL10Lcox4lC+f9Y0UooldDIgjD5uZxHAZzdAXmsmVlAJ7iMu/Y7p6CCrNuI1
/SnizsyIPgRB1OCpUnO7BOIMqRSgKd8844zBA6p9TUMF18q+YbwRS/D7nHzHTtYl
oQ3c20MXFYN3ppLp9o1y5mIlcDp4ohD+l4IvZh9edZM=
`protect END_PROTECTED
