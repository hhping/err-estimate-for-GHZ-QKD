`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uMRIYp6fBJJ6vQZoiM+0UhO4lof9iu56KtaKfgaTX7d6GN6+OD/Xp0bYGhNu25eR
tMEjAIrK1fSWCn36VyG63P1es5oYjazRyhiJ6AXCSj83fIBBG99YxjyT8nN2zTK/
Upn/6ozVBIPZG5VP/Ffr5N1uWBfn2+WjPBiiEY1rsJp16z7Q4W6RC54PlwGmS0Ls
zr7hQwFQT+/Vg5CbPyps1NOikiSkCfLbOIVDiISnckXl1moiPhQLz2A5lUL2QBml
PMMqghtPMKg50IcBaYCNAvN1Bj5pcecyEGHLYvi4xxXUvOCcTWuyT8awvz1ZMjRw
cAkwG/lPvylHWJGPvwVy00QMmjK/276UtPnSYlo/op6ZFEgnzpE0o0Sz+1SIljHC
irEsWLVhOwjR+9da129mExBbOF9FNynlFSPzjPT95dQ=
`protect END_PROTECTED
