`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QuwIR/Vy0/s2wLqTaIl526Z+mea3s8kEiyxQJ9klcHHhqCNkvmu/RZ5UjMq7J7Im
Mv7Fht8qBk8vpBuZCx96x+QKHWI/E2T966A899GCTT5QR7C1qMv3AWOtBG00OfeN
3fV17Im6G3cp/7J3SON+/4MUMuOWbmt1L0PT8rwSctER4kgwgyvZP/jcV0T527aM
5LWP4TAhKWlCEzc7l0YMeAHY+05rjmVtEnH6sVKs9ztaU5JiNFaIrQZrb4F4eTWF
SeJ4waFL/fmuFYB2qfIIVlzY90sfI7Snopbn4X4wzBn7RpY/uypo9RGx5r268ojb
n1a4BWBSsHcJXGAgF9VJAk8ZyLXF6iNw6kBh4avFU5Bvn+i8+kU3F29Vm7x3/XTD
LIBlhwbUeZTemyUzQ3mw9YD/X2KyxYtTmAmLt32HrHRriFRTWxVMJwfr70Hqzn90
m95FdfeZOC8fvsEBhFboEGOwYCoRN1WXH5Btgh1JUGlxizMiOge5UD+U40Noz+i+
4MYtNTqmUOs5h7duj/NCtXfYI8QfKk5W6WoDUZMDuIRsuU67MNckTqysNNm/c/Zs
B68gVuO1B10+TzslJKWNHiubAnlwXJ21jCki1UQxO+4NDMUGr5BEiJGqFWn5oCXk
Oe39JDRJ1jrSf8J1/OEFHKAV7ua0BmYftMYVwrBX16QKar6GS328QrE6JfAmx5oR
6aspg0mNfHD++XniqsM0dOOmwSG6PMYOCWFOzuA2LFiCdPuAmLOjACwFmEZXqnQi
W9Xs2MLpW95XZVyVnZwLzs4GaTC+WmR74CctpKGC5dU8Z9gD29hasU8ZxIR+ujjG
VWMvMk1IET2C9s1lO3hlesF7wuIAWbKkEphV8qmBg886CWuDC3oesV0avDbq9qHo
mEmyK6IwExvf+42uRWF8DUaMJ7zMUqMMsYMvOZQsHAnLlBvu/burpbTNrbFN1uOh
q1ahvN7e9Kn8ciweo55l32Iyt600IM8ubGC8n9U9Av0ONQNGvqcaJjPkkAqfu4YD
H2EsWzXfjYJrebdo0veGpKTZtW/iZl5ojH3u+TMPcAPq0386OwCkCAvR3/0X2DIz
a8umOqWbv7jnxJZVkHz8K1BFVpK5jIaTYpOV54/y/rFtGU+VdKocgP703Aew4j5Y
272EOcioCEIZXD8l5h3LUmi77HUIQ/xYCnIK274+BnOVEyoO5qKLxoaU/+v86ErG
Ulmbn9h7vtrea5W/PubdfIHLnY14Z7AlFfv3+ecW36XKaabXLpg4VTtN7Qcd40cl
y9urlR9u3DKpqk2gFJitSy2dnyuLf4yjMTaGAiXC4+0s2ViqelFt7l4LNEB0N5ec
RCgGKVst1g5xpIngqGvLO/gZmPuLhtPrV4/ajXN6yMAVZdPoVbyl6J0tNIi7PaXl
oHAgVBDVGk+PEA4XISdqH5QEEz88NVaRe2H7hNFDZNlthTfY2JofxJG6LTg69BCi
KnkaX0/4hh4k1kGnNBkGn406WDMMGCW0zMfFwuWkiT2rsFrob5NI8uOqzwrZrU/P
C/ROIJSsyITZyFHhGZuicIS3afa6yNgm8kzjJYfIsWTtwqclDEfdHeUo3vnhgekg
yVRc/e9fxfNjbK7+0ifLbDS4tx+fpauseXdfBOfmDBju4G6Q4A94IIpd19/FWPLl
VaCu2qiU9cTr6qsGyckKRS9POC9K7LyGutJuq0z/o+YnxcZx8bYhCYBkyLeoAq+I
p8QM7aOfzyoa2eesx/lTkZle3/TMhoThnBZvCk8Gr+YocaYIkSEewUw7J39fa3Jp
IbKUObvMXoeANZnE3JtHmHHcfUVgc6gDDNuVvpCprpR597sqGq/bp+By71Xhdlap
t8uDSirNH/gJIbevoP9e7jMBrqHko6YTTPDO8FLiyjg+V2K79mLFklcwpGv0TN7v
zhlxKXQK0HQBF5ZXts81HfjBenAxdE8GpNLPN4Dd24V28nCjHHLwAyLr/TpsxKqx
tZsgbaFOfkgpSLycoosQpKd4YEhO/osOvU2yFehCm7+e1TAFH32spnCKv2AN+4NW
/n1gQGI5BkfK+fzdHrEBldEAMhr5jVCBFd2g8MBmJjvtguxO7wC5mJRAcIH8poPu
N9OgyagX2njp5y/BaPpXJv9Bwwwi1uyuV0xMVYusFk77s6fUiZCQ7+/qPh3mQYZj
0DDqIWMAiGJgdY3sVfFgoh9UGuo5yev+jjSiHJkA/OzU7Bej9unLPocG54CoN9im
VTJMP+S/u5iiIWo/SNFuWF2L4KMgZ3Sy1XlsP7a0yM2MVAJnaFcWFEyyRYGyeWjC
4z+5HlzL3iHEytByrxo5q0t1ApkH22XY57NvTrrPanvMdbG2RIJVQpnZIbuMk/Z1
8B159X5BrKpCQB3QYSyyYcpDBOr84CYr2XeTExjDf3ZFO2WasGzYyNAnU5I/gj3v
7SKztc6uEpXNzz4zIpJ4jOvWgyoZXsqCwxYom/1Gdxf2uWpo4E1UWIYeMfk91b9k
vje0z6lgbkIKTJJ8WhqY32kdiQc3YjB619aCftbSGHweTcCdUsDnst+pqcHtr/TY
OkCW1TyzlUgKk4++xtUybt7UH4MrrxyeIo8hqdpEfAaCd29zd4tmXyqkI91dQjC4
xA0wvsXvoTNSfTjoUoE5vCECCyIQld6TsrfZ8dcG6nLkzc/U4nXWQi2xwguj635m
YiXduGPiY1jSFiklH8bvreUMQThp5C+I6BjeZJdyP3pRQbYQ+s5PciL8CON0MPl9
2x+W5hOXHPZJ14P0eUahb6m7h9x5kylTBxqH2sk628kY7knEIHCuEaOmxWsJtFss
NJEd3wlJuVVu1m4BhX+yzAGqe0aqwOO7b4SuTq0o9L2tMqEgySyxk7ACNPeEHzye
H+q6rtbrrWjjsw/o1OpvowKkFN9a4aKfB4WCK49dSwSi0MAI2sZ1pid/xTx0+BrH
i8GX+E4wL/yyV9W9yr+BCghE+JHtc0xS2STPHY7W+unSmf5QfmyRYCWs8di9+sZY
z1uWODMDiPLoK8ODelaKYTxWFXjNexGba6em6J7c08GSfZuIXzjVXwnm9MwsMmpu
J3j1Jjj9Ho7n6Gm/056/ITu4MVASihmvGe07KvuxfcyqU3Rqw91DbN0lBdfLGijN
irmmsBo44Qr/EyGkRDMq6NptXhjNKk4+iLe0bWxh9DRRxAPbz1a0kK18p6kXnLGC
zsDEkA/pcbMfDBESBoDY6uzNW1ukkv8cU2bU7JmxcKlcwrZih+aLys43dWjaXflL
qrpvCkLa+VS020i4ivn+GC9cMGd0DzfZ3pT1eKbVT2iCFhRG0k2bqLxNEgfpUKOC
3d6ls5N4T5v9ggW+E8Ds5b+P8tmUhDb9XIBRIqGLWNpbRT3KpvWvwEQ+Ha9h/Y10
QIbgcGg2zsDBl85GMeeUw0ejG8Xq8RNzEQq7y/kQ2F0YnIQYE7YO0eZ7KuPz4/uU
P5SVHTI1Iw2aXLKA5Xbc5IDfRnblIFW22vZNY06aO/VqkslG2EugmyA0EUuRyiV2
HFDRT41+9bv74HL1c50ey8IPI+vq1wwQ/4PkPAQlBB6qhEvg5WUdCL3H0QBXAYXb
tsWVPy4Q5n1FJb6zm5ubdcnp74vPo3ALZzw0JdAL1Ww61woSQz3Wv8CYJGtzMJ+2
S/prDmrc3quSEYEuw1cbCAdIL8f5l/xiy86X4hJXTd9fI6VsNpnCN41dtFOFOq8i
Ot68qi8aSpBchrA2UhfHlAjl7XPXuX4VjyXCFlspz3Tza9ODO78lJHg4owFYGHe0
oJuavT+qWLjPBVVHfRDozahiKqhVPjGzbCtosM0oy/BgYqy3s7DWPlpCAQRKpgZw
QZXcAARmHFUTJDfUYEhX09fT2DsAc949HxBM/G5FJXsJL6m7oZFmWKWqIsLdhx79
ozcvZ6WHhNghA7mXlqeacyvAuByhRJHw+PcQfhP/hGJii8i8VY+ptA+uA2EP48Lh
DYYKpjNPm1spWoU/roq2DNvYrUoWNTRRbzGCl6os6lVM1EirE0Ebo9cO1PUHQNRt
iPSzgRqL0WdgmrRRDgyNLUhkPCsGjAVy7dHT8/v3lH1cfI6k5Lo5JObBYKujfo6C
tvNlXGltdsbHc71hNcEgQNpj/nA8ePDu74UxTtMZxc+dh22K8Ph2sEQIeRJ84py3
Ut1I4jYAGleTh+4om0sq/tAPHKQqnskqtSAm5NbWC7iTIz9+Y/WUc7weuHp0dxog
gMCKTxt67uqeL1pud/RuJL2kIlXgaa4RZUtZAws2rBSUXx9J1SXndxqrs7oyJkWa
/DLOHa9MVNacS8/w4mCWngD4IflETYfyidoXsrqMc4lXT/CYDBiTsU6NmKuHc2ZF
Rp2iMzd/V8NqRY+5oALajwtAv246YmAxx1S/JbDiEVof/+lfvyW5SQ1zW7fuX/JA
Bh4CQ4wItQcC0jeRYEgUgleOK5Fru8XP462vq8kqjJPgl5jQvAY3LXK1jTfCxaEJ
24da3IzapVnmj4FLadyzw12A2qMt9nMBgyVr2Z7Zpbm1xSdyUc5qmqhf0vjQDUyV
gTtNIBFof/cJ69bp1/yx8PwK3j6YMWcS9vT2FWFTFpVv1xfuelfNQCOaC8kat83E
rZs53TFCY1QgjYFryOfVqaWDvb7KR0hBFmSpsVtLyw7IMoSrbnemecotytDTqwXL
5uTzhpHK6uNPYMDaQxySKOuOwXbi8nFNhRY3PQgHwCQk6GvMcq+tbGBy34zDaHtG
x2DUobrptNg+K3h0nbCqlA79JZZYyja5uylnTPohNUiSXMrE5vteAC3RmwKz/7PT
Q/VJxDAYLrkKZWJ0gkbr4gKwhRYl20QppjSt33sytXHeEyBLcvJ+I6EpBwisQcfA
36vhHhfwuAFfx1vgb0h+1xOxSIeOfaHu/WFBdavxQWjCX5OhyFLDKkOcBfS1o6pB
wJkLHUc2Awygvsrripe9Len89rBPWZ3Mwx106B7euGXLVkgWW5zG1uaJ0e1T8XxP
YGiIrjkF0a6WUWao1AJBuiVKK4sOL2jZQdsiO6uZ4vgYncjxTV3cLy/lcBuv/QJt
xGkSDTRB7gprmxVOJzfnNdLK2OV/dhTLyZ3PEmCXRTP2c/mYT/IIT3RigMyBawgQ
hAXLca3ksHO+asdaH2zSKy6+3kSTSUUxV0pOZccL4F9FtHyUVym/0wVGCWXSilDL
/HTUZZEM22ejmUOWmBqw6HYH1gIxsoEY/L/beB/7LlSw4e4b+er9LxKWrbcmxV61
Vp2CgrvF/UhVZ2kC0FvsWXF0TOeewMrV1/02Wv5OIeUZihIDqclgkbkpxu3DqczD
6YeQOrG+3i/rxQgseHMQUFDa38rMVo5IamK6U6b5ftwROSsP7YFogbarXBvpaTGw
JjUnfyGGwQaIhvTDNqDd0MOO2ATrK+SAmdF3UkOYc3aGqUC1qohOSV+Sk2US/CL5
HXpT7Ud0xHsMyEmeiD/n9cYB6LWqmqUAHea/lDBn0VfRfG6rsgO82vT4mBUNq98n
kIJkxGUEzgDBAIJMO0UM3vILHpWqEmHkWLRjgulrx49QL2GJfz8REQJsFv0Q57FP
yF/ya+ul9wybgSFLFJ6UFiWy1/EamEipIO1faEq7k4ULm9XjhAOPxOZeoRvAMHSw
4OWmvkTBXbPhXkt8qBFay9YYISjcLCOuIgHEETgln1SvRRbbjwwjVXBVSuAK3F+I
9s9+AelRvFcQbqFXJOO1lzsMuE4tI7mp+KeR/ywcNuw3rMYsU/zD6rR0Q5LuujlX
tz6oqd1R33E6GDpDVtomQnKmInJk2PZA0jzapeFohXWOwpDanUAV/ewHWSMz6ATE
HXPOXvyD90FhmrV5J0OedVC531x/jHgE2rtPShWXWkI90kO5fccg/dS3xABajd2h
6GVXm1w9j98/8B7tNs3YzOfG9fU4otmHFeLlrTvEEnwJtpiaDvQZnZk4eKrAAny+
uBrmxkscoESQhZC71z6mJHq5F+dTp02QmmDrVfwUSlKgpW2kg4OVcK/hwcnobmmM
Wp/f6Q5nXgUPn4CrdS3hkFZds+a3ZZ5KshOa4VBkhGKGbR8z7fLoCZ/C4yydiQOO
ALpiB1++HEYblzSguu20uIyBAUqCvFzny4BZ30hDWORlh55iTN7i51hDhzakD57y
dqoNV9vMroTQjDupSamj4rWx4VUjeiyw7O3jLGbea1/kW1PH1pdlgMyp3IW7FIQ4
95Dd1tUe7OKMGZv3QZ2vF2PAL7nvraKhIG+C8XnQt+U4SriJdDI/uf8zPBw8Ftoa
8+h9Wgn+a3uAysUVXGmmrosrdS7rrMyGK9pI6iyworhv+eTGiw/1CeUh8/C7Eh3v
OWfuYvMGVYUYu54zhPQHKJsmgZV9cobL922a1rPSx1U51K7oKDuk8jZomJviLpD8
9NnEjAAjpHcFn51V26eatsCL0A47aOUmruSZ7kaVaszwviPCm52UWxrTraiNNpfZ
93f1/sTH2jNYDOr+OrDjaZLVRmGFU5aJDG7VSTBRB2SdMSkItiiRsrmhYmPn9173
jHam2R9RTgH0zDT3euvEnFtAmIcJgmCo0wrjTyLwoTenxTpFyoZKjvTYNiiNC5dJ
thFw4e30gbU8Jcv/5hIca2fLBno1/8Xf9HiG4ZHhubASUTYVxrmAtFRoNk1Kf7X+
su7sJADhFzVc3o3RMvKnEpyrDluiNA9x7i9RkwTSj2AGw3LUPTb9ynDc6yj95jNn
pqL9o/cNDIKBEbtJ05HvGDSakQTokheZ8RKc0wXmrWBEe0JqJNhdYx/l5kBr9Z16
PFmf0ZovrflrWqHCjs/UkPsdbs2m6Q1VZ2vAxftNIH9m7zsnClfzgLQZZVvIOs05
xaDPy6oU0P5S7sa+0YbxcPhlEWaLlwKYSsYZP1Z7RnQKRZe8vXxQosXA37cGWMVe
WOobgvxq2ZFWLrUckKzcf+WF6inXZctU1p9pMSl46VjWdiAfN+EoufM7Zo6eAIuJ
dxCIzLPytDfw7rvBtTZ4KbblK5TlRSaRTFUeR1E/pnLFJNUlYSJPx3e8Z55Gqr7m
ZNZUdR9C1ECsxj2KK47NuKgFDHFhtfZBG0WwKRUqP2ZqsnGAJpHllI25gcqroQPw
Vpq54l8waoQvNz7U+Jx/yloCOMOxWjl3A051jDbRvl2KH9SERJoYu3USJQGg88YO
od5XqTlEBgsQqSYSfQhf+de3NNWNPIjlQoYPpNLKrcGCmRh2oPqpQ3uphDWbFF5M
07FNlVaG5KbICVTkHTEzrzTs/CSH4TB7ClDDbDdUWCrus4RJZoVuBIHwv/wxfzbY
Qq726n2dZOmzsEGgUiq6Qjx/dm9hDCQ9PEeEFU7ZDoTZ2DIfN1OpOZvUxP4SZ4dJ
M9qaBlQt1H1jsXjaO+kBnuy+Ganj5DKUAavnpinLUs3S+TwIJqNnbSGegKnF1h9i
2RLZ7DOcZZ2i+KpwwXlKyZm1Izom1yullWwInSyglg/6darnbxQcmPye3XTDmo6B
8KXhG8HGt3z/Pwsz9N0nuefWQM/GTQDnWe3hM8luNlsKqwimPlbfz5hUoJ7a+79l
4KbRel0ffix2GFwfXhGCTY9XhmugE6ltzI7kb88k2+lge/6goSTlP9SgEyw1nDY6
w4ZCKpw80EN60Gkap9VSjEcy4eHtRQ5pG6WieVvfuYPAouu8ItUuCJ+zegsa+Iye
Wccj68YanVVSgmqjIJI/SZVA7gpKI8fv/Bm8pnvHvL61N7myHWoF4tCc/0foYL1Q
u291qgrtHLJccOZFukBc4xoDRlwyFjGTOqXV6YQ6EYcIm+n8eYwu31LaAQ7raGjs
cBInl9J/du82WjhlWv3NQKeUC64z8tUkMRqpib164oBWndAnqNIaoIa1UsOj57yM
DuIbgAb54+AGTi8CJnhcH2aNkLpTQrwd1NgUhub0RqA9iIpHRVfR9UddSrAFE9By
hy2R9cnrMqrpPCSEuXVZipyL/Pc97CFcejngZwadGLt7kLonBGnCOos8uhxUraOS
ARtuWJg2Z1jtuSgzkOQIr/MxfYPCbU8/iBe/HB9SV+xaeWesgGFOBnbTTSxEelCY
pqhvcx9aQZxQnG1Fe49T327xB6VkySiqZ2ecztuhgazPOkTS+7IgOdc8zooKEDWS
BTP7ZoRVmLuSM625s286TB8PN5+JnCiUwTVfm2Lt4d/qfgkbam4kCYquSJ6fpVbH
xmW5kbP8lUJ5NgBWJ+XhX3jR+49QD279ja0RHZopy4BERzmHFl8XqJhoLoOUhbXi
Q8Yr6XZjqZHKMO5XAA9KB/K4Ucb3hivcjMF2OPUEZfX3mDTkrjMXFpzx6eu2yLBJ
rhyEalwz3/d/kG3te+2B4nso+pC2T4VbgQRJ7nPcArX/Hj3h+qmTkC8w7gAIKB1o
8GH23nnubMQ5Dxm9B2x3+Uc74XE0520oLEAv08vzyAjKR/OxjQvXEBGWAYleM9Na
cDlABwvhmStHRBaugLUlKrKRw6zcfn8jctgG1ndmkhFwsZrxg+y42IEG8jNF6qa7
E9UI6TpxsHJ8mYb/toohhcjfYMVRtpvrGlBlHjA0eQjZpGgsxbLfqlLLzGeFm7i9
UqabiHy7Ooei+0fPlu5ziKaA7O+jZV8V3mDmah4x8n159JCgi/Z4iALbD+6QbEV3
QABpWioqzUGcVp5WE+A1Kw37flBgAsHIXImgrBdMrrmY2CC9Y9Hse+dNi6W0GUrU
Th0eQ021c5mQ2kCeyt5yO5NX4geo2GT+YnzOlLIunDUexw9AwnPMjtLWIe0+1gc2
ZsIv1dtn89zEEowsM/llxB6KbFU5/Qsr2qXvYAWp5zHVWLqeKfqyOoPetVdb0/3q
HbZYIF8nLzjS+w/3ts7Baqwmky7K05brKt+udFffvhFg1pEibpf50Y1Cnkn/dme2
h4u4ZP/SV5KlRGI+MfNhRRismVGAIWwYjnDlkJIQljN8imtD8G3Bf6FP60qWDBrz
murBNqlABbqvq9y03Mtg0sOIrx9wEWFIRDREKTu/kgP4JU6QlbGRdVpzjUBw6fNa
n2Kt52ymf2dYiC13zNjzrpgo5xJDceEoVDevsQnNJbdiGJnphmE7KNHqJXylvwTH
JV8dC3YLUiGMyZT8/kBZmkpE1vS1hKiMzE6ts9atn/nnfvlQ7sP4gWFx787Vxu5h
n0LQLtQy/7ydGAxHvGaj4UANAS5TkkkxBPQZMPrpR/ywT+7bteH+NT3dilya1mME
NuK+8/OLy/mUxy5KruwtAEUK/NRAW452yz8qmIB7lFlLU/U04ap5A2atmNvCs7KJ
hq5d6VlUi//i7Wub/bPTCY/BkCFYmbqsAGuYGnH9tyuMuAJZXj8lUBbBdfMeF7JU
1cxfOKbjPcOHe5P6B/vpMeETvBrUWvqbDtRvO0N3nSTIc2vxh0LYCgvQkuLrr3qa
IUwjyg7IQtEtwJDYHAsW1w6CQQ4uUckVdmMHIyUoY8dVuAwposH0SDihci5LmqSN
Ll8jA2/8wrXB/N5N3iHHPNTgCilIea4nJp5mpWKXKwfeLRiFnplOoOOkL6qmcZuo
yhROiu/RxHKH6qWgwVaQrnWUE7qnR3Xj0LdQWtt2EUmjnyE9OwB443uvAomeH7Pe
3iEcmhbyY8/oNit6NwvXDdFwthHe3J95sgXDkRo4e0CfJ7LMYXvMkzXgrein+fG8
pc5i9oN5qpQ5uYfMvNAj29/B/ZuNsORr+3HY4ds/i6fz31dz7Md+bmZ+qxXHia+8
wbjHNnPjLJwSGEh75BPOxrWnNyGLy+A43LplpBXC/vs5rPG+ifxEC6OvovU4fwEQ
byIGbf2fzQRn09mjZkjdYelSZiD3KIAyrWjEalZYxaOULRG1qYBivEYUnYZ9bduJ
dN36tSjFpRphr95lvTmSTknB8ZoN+qseMikdT6tGQeRryIZo6bAkKZAZtBF0XvIs
EO7IYduPlFBF7v6PtrtKqL+9GbCh7Xv/DA790g2DC7vDahb6o/aA2OXNNxLorcuJ
WL5qAwDYefgG/gTubUCjaDVMV+gYYu8o4/6myE7ZUqckXHFlQ7EFkmTqOmteq5eY
6r5PxQwAa7u2sIBAgSSEQE6R7OujzGeA4mUuRy2toHvWaTcKNLanJrncF7ptopxu
2VHzcs4FHr+i4+lx9hVZ1/xYUfJNNFHVDyn9JDQXIzZDoTwDmYbIyvbzvLZe2HQV
ErkRHn+EDSiVOaCmIQYiJzgRqSjvAeYzH+JaYNb1WWxGstNEpwyPfKhcb8Lwg9VD
dTpkbDWzgxHwOgkWCUefTgSJhhsQfwpmlbbRRviWgcYgBlhRSgMTAxsTnKGAyEyW
kz5bKuoWjgv8LIK8cYBIUdIBURhEJMNT8RwLynnx6ddNAGkCESBsol7o7hudAGox
llYP0HOdY5KJDD0Nv2oYsv9WWj8e/mptJD+9jwxkU1z96IRfRbignUrd+7sLO7mN
75TqHXYcHZK5xVib6WiC7NR8aAY4ZSU5sOcXQ+uNDnc2kRc/l3HhBOrriKjShzd4
Jg0dI4LfBzKfbAZEjNw+yP+4oYfFqSFPs+nDmKLuhyFIAy5U51gO2wFgL1Q9MS/5
ycsTa8lce3ZqgJig+Vf8wg==
`protect END_PROTECTED
