`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OiIm6fXGQf3H6CdjLRLmK5r+1I79EsQzbbJchZfUNWpgU/zYnUY4acSCDr8KNWIO
n+iAR3BkG7JlPuxtEwkVwiXjgoAe1EdnNHWsI6dNpihNAxeH1ukVLeaII0YlSBst
Pym1wx/rwJxiAU0/eVI7gBXQL0WI1HPubLt86YLmI8ffZLXE0Suz96bAMR6ZjSw7
ZnLECdGfXk42CI/Q6NWCbnERuT6WwSUfUzh0FDN0C9owFiDLGhO7fR84Oe0hDDMV
0W9OEp2cJdHkqbk9JeI0HtdqFiBGCLl4BRHA8VVoChW+NrQ9Y70v/DRrzADGam8j
RFHrhJRm4SrGTDdKwWHgN+25GUnprJEXcGCKJdSb0b+Dxg/mTKuEYzc9JVYEMZOF
uLycer5OY5vhsm1N4DDgR6AtUcU55jLIWAAj0aduGCXNtEJBLMPK+dZD2cVMp4dT
x99EpfJ1TbEOZ7B41/NB8nY8+LiGrPC/zLkXmKQTUi9RTyJOhD3g/S3GpxHq1Tvs
noVQ1tzgJcuz3gBvm5fGzVbraUzYZ1C7dnYVEisTLFDRs9V/Cf6HI7y378FPprpu
ovq6zn4ld2dBuuFpTbQ/ePPCjCceeyr/3ryuJ4cwz08jv0lZBjCIPUaC1FmeVNJL
hWD/fdR2FAaijRgT7R5UkScYE4sJQprrScxS3Dim+dyie9Eim4KQm5Omjv6IF1TL
O8wzErORjymwB7JHS7tS7Jc47rlg9ojKN4L86YJNxF3fzOx9LTGgezJmyV9xmJBQ
C2XUBJw9bU3DTiodh7876ZRyDm9poVsufHmQy/o18z3T3P/F0al4+8piuDaRwz8X
zwScgT1EfR+fcS+4YUyQKoekbNv48iiigdgQosssEvzW+nJmHzOaaDGo2oaEXv0k
ZSKx3P/VPhFWLy5Z8VPUeG9t3tUDG73CrN371gGtq/J1pDc1+wugKamyaEJxx4KR
`protect END_PROTECTED
