`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gNt0zb3E+MlnBahvuQgAawRkE8BYMYB5t44V1ZjWBWaPZA0vX09VdrtCQjUBC97r
7CGyzFYluHv4w/EBLPLZlzFJ6iftNtu4Yg4b5ginFR6PhthPDRvVWNB9lYcZ7PAa
LptRS42d/eK6PzgPXnn+7m+sa21EopnwgwhX4KSztBwnT1v16hfbNn64kC9AuW7r
B1r+wyJtnY9CrcxN4DkXlqHC4NdnWjA1kzRDMNvawglwyLdiT+UKj7m8Ruv9n4rZ
o23J0bo4A+msvTAT9fIv94pISlKoIX3lTLck7td/gyadKizq2tjaUujjBmSpx00l
kaA90DIdklarMJ9vtkzAMtr5lwFx26IXXwNx0JQMQQyeBEBrfQLyuom2LAB5b7uk
viUNx7gYR1rMXABXn8YvJNFf7wwUK3R2vCXwXgaedGrQLqXaqioi8NDrz6ahyV92
p+otCk2WGksQcDTPqZPgDFKNzSYNwFgYPy4xYZ+gom/9fPBw6cPeAHyfa1U1G4qB
B7AC1QzvvgIHpjWv2hIrmuzE1pG37dY6dRZtPJNhN1/yeokjTsyeqmqjArVr5dVJ
AKloMm6i4Pma6FyaGiLZCNOdKaDYimSGb/2sCKh+xGF2jKZ3kMAAgXUWIUsn91WR
cgAlIjKHVlesW8pFIhN6Mz+QrIle/jevnulSaDWCgVb154dXxEeGXLNYNHd15wCc
agfd+Te350e0VA7qXbycIImSGIbShUyYWEio0iyHUkuJtIq+nz39+Ufu+mS/6gc+
YfE2KL98v8HqiBmZH+GMvExors5+0Utt1pEwTtvE6x5qUaqlxyMZtGvqx3aHa0AV
dYXxb19Jni8p3mZKzyzWpiRU3/zHFK++MXJ13U5fYs8=
`protect END_PROTECTED
