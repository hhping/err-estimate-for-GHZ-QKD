`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T0QtyQOxTvGK3gMeG1Nn8DLDgi0EofPQk+GpgeTDeSWcTQCZN5snTL2qZyG069B5
3Tjb41KYDt7UA396uAGsE/rt0sp/Q5QbWu1vUrGQdRLgweK14z7wjBI+ucb/6CsZ
oMZ89sFTVDsfPpoA1VKGYKQOjFy4jwYMzmBvZ624hCJ9NKo9zUT99aLOHyLMkxS8
Ab5QPrmu5XRxxiRqHelx99L5mqPfOQtisB7f/in1ifhDCzBIT69iz7FnfUmihE7I
DGtKuX3YaIjATjyJ+XJ5SM7T1e6mqMPV1YObjZJ+8/rXdmS3Mppr0JW1GdE3iV1K
M3nPYAe2891/d63j2RxU76C1WliayyV3MSGpbzSFkfj1/SQN3SGMA36M+9lW/9J4
+4RrLO2De5bPy3epB+p2BVHTl2FbVZIwV2QNbagYNQifOWu5bHy9pK9jnLg6rxlB
J14uxJttEO/yUeokgHnSyE/Dy6vHCduBIV/B6hOL4XJqQZPMPIf+JeMBq+hhYXlm
gDi6j6KG9p/aUxrdaxafNrkhR/QhR/0Yg+FNJ0AVif66+r0mMUlM4uy5siuaZc9v
Oe/AgGxLrTUCs5SzkI4lVDHd92NBi442D88HQHUSiGbXeTrMo9XL3Kbvm8fnouPK
h7sO0E7Z0k7BiLH6gYFGvALOA46biSeihLPB39gbeT3K9Q/8D5DWxUSNFddS6O88
RCsAo4yQZXzvy4nwpGJzB8pXCYDQcUdy9E9v9PmbuhdGe0KfRkjTJ3Y2kfcANA+E
fY06Ii0Mz1ytpQw2KNqIUZC/B1q+Lsp+npWBQZfwFwDrrL0fg5s2lTqCmPViBNI+
TtRiMc10wsfovisi8zD0sgKoVUFvusmAxmYs7ifMaXkjjD4Ndl3SWNvNRSkj7ocy
in3rD5EYRnLvsVHCSsfAv7iUA+8P26V1klL+bAgQD33ttPA8kedXwDkFRMuA94AX
P6dLTXvwn0aIXi6+cmtzZnAgqcNGNHH2L4kpcKq8lT7XbABzv1tuyZTPc5I/7v49
DeF/ALeACh2eH4mFV1iJegTgKCofvKqNoIv97lCLkGhoqbndpBNmZVkZSnTAZEDl
Es1Kxrmco5MOMOsrmsInY0HzsWDYIaqFE9IblfL2wpBCGE836KoHRcuB64uq6pB1
v/M1cL/HmU69V/tJdSWV7Pz8mB7qIhJ0mPrHOaGw8yfT1iCbXwu3ew4IeuTr3HRR
uwRwuph5se4CVGbs6/jwFYWH9M8SY5tXoA+6npVu3nB6ud5Sf3nmvaODm4YpaFvd
PEdS0A9OjmAC/m1MNjbQtM30hLyW0uYMXzPwiutBxai5lhR8bsFAIHz8p+jNb+QT
z7RBKEwyCbSqNs273SXl/jdPxm/Qdwri/5mx9aFkzEHQTxStIfJAlOmlwbh/c/E3
drC53TAlh4anLnlS/CmQghxbRpx03uOswtzgWkz9BIIX3p6rZ+ES5IqOK9SSIaeY
6BJ7sk48Ei/mNJh6IaK5iP9+XPM/iP5TnNOMJne0HZ6H6P3nSYGC4H+lTFnkBowd
4Nr1Wfxonf+2i8VPD0C28a1DpHY+wLfqyjGEJ+pwnTUuqJJPSmYd2CPlk/i7rLKc
aPu4rXGsovKj5cdCKWtXXYU1GHj2kwZ2RI00K57OBPAkpnXvkmMAD82Djfjt1YPQ
i5a7X/vPsFr2cszcP2Udd7vEBZVkivecZV/71S7DX+NjVV0I58ifpgZaCDd5T2q1
pnSV1ibmPKz9i2lsoWTWBGY3PpJpQYx70oksARgL0eecfjBA8TzdeSqvoH+k5H6X
JK3SXSglWWN68KL+uId5z+oNOWxVhclxQRX1u8D+jNqZu5I3b2PBwTncKnqtnv9v
wiheBVzUiy9uNqWhtXRknjAi8S3PGYaWCRtbHUEfgtLu2y2qBNvYawL88r65vroD
noLkqMfuUFPVZLO3K88eC//TmN0bWGGaAdDrxje70P41ZjhEP7BISOUYywRxwsB/
8t4yq3w+LtENK/d/d9avGc3kXY5Jtg+0tYovxZUndVzlRyZ+5zH2wOGx3ciMCRYe
6DK7ah7WuuPFahrESr+TyI9VVS848UB/GD50tEuQbI5lkGOtGMsHJovNJCDd5FRx
duEKY78j4cXXLIZqwzFIQV2uG0Ca/6hbCZHd/D8nVwxERgY4fAqRAKOy7Tueg2pm
QSoda1dd2ldF5mXY+3XZ9dkpEBAYu6HxDXvNIQ+6nNs1bACdK7oFF6Dfza86VXc0
mNznMauyE7UP+wKZVnBIeGa9dCXUc/x9KHayAma/Ox7BsN1CDMHwL7yNXqjr+o/R
SFP8+Wpm1RVXB4oYEr13vmZyV2CtoZsgYKLQPOXKztA+dGzGY4HYjjDDfD26lIar
Bw3hzpa4UiBBqKn2Y/GbpAQ+APJ8jZkCALWUfgY8zND47B8Ms4p6dD/tJ7zf8eqo
Yr2TWVDm3jBqNuzMilcPNGpGtKS960IXpCGS2wwUd6M67JOSYZqbvYdMfJExtzhj
9dnM2cLIkWDaW2FwlvdOSsYU/tC7Nt4szmnRfo/b8k211SdMGf++Relavt6zwULh
3v6g5rPl5O7eIkBkaiRg0Hfln+0DwU6zXSGGs/gLvEd4CSVbVuQUzM8u9SwaK5xg
5m8PHg2qkmt6i98AqhwCeTQUYwOFra1zYowL+EmxeJBEei61DYbzoRupg9V5I+wZ
XD96fBWTtHeN2XjzQoBXJe5ymanJayUbonpS1aPpvzRzyycvKnOqbUkUHuXWbDAT
sMlgEJjx4a5Ckt6ykF+B7lCJZ8W/QAKKxccsCq7A+Vn4FQAEBPPWwK0EuHhPa25h
`protect END_PROTECTED
