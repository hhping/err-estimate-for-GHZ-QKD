`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2+nIw/sya3Qpz/Kt5YbinECijBPryW2oJd6xqzhLpsbVQVWsfZSuYHyZzZAIu7gQ
gOhDm/oxq1/7cP4WeucSsFBmScM6dQfes2purH25bUSpsbgZ9k8YGiMHlqZSfShB
YUNSMZtjj1Nqdpuv/NVc2eZqVqrkOvNorttacyo1fsneoqSOWdMdbRpXd/2qFovU
9ajz/AXUxvU/DEzJxulEhF2FTCLv7gScfaAl2oRdlVQpxbgNJXA1nGQekGWLzAHV
kbdYHG5gDs9y+5jx9PFGN4hZcLSK4mYw9vV53Lsm/5w=
`protect END_PROTECTED
