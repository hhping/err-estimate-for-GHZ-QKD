`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s40+awTv/HnG9zdyu6t39FnUvPve90uOq1yZzYvvxb5gQQeXqaXEHL12JpMX/MFV
CyZogGd0DSkrBPFOpG1u7LgSv6U2kjO6+PXuIcKfbumBlmZ0+EmgNsshbqeLOw9+
QKFrwp+rrk1ZhWhwdpNw1CzZXPclXlcKQ20nIRRVGEDwiFBvZfRVR3sZrlFI0KrI
j9astmrTYidAxLKzdIDGdMlT9uMXaMUIA1WYEzuCp1wSzQCjRj7yrc5daqabABT+
MROHVkr0N+lm6KQ4Sb01MqwBTL2r1srDCiNQMJf8yrB93AWgytOsQtmyvQpji6T4
Gh7S+S6c/UDDTDba/qyl96nVr2DAfMi9fttA0zPgbZ1080zKHKm0pIBr8Et4fdtN
YIuWnBcbkgNu1xGESJon02ATmsxCYAWkjdENxUGveAHctxij22Ri5qywFi7C3JhB
+UXm6gJIZolvy1STyf4LJi951jd/w2n+TwfMPXIzOYyYxLxCcLfBhApP+J8ltPX3
BV8aK0on1YRwCWA1w3UqdYUU+ue1lc9TQuC09JSWCWEU8WndVakcUQXgjN5UTrez
5Yu1I+NRKR54Ej4GoAwC/ARUVgdx8Ig7tuxCKpe45ztjkMZqMCs2v7NIP1BQQdD7
x8qO+QRi0OL+NBCokv35ZBHRoioLICCLCEpf5QDQTAcHw8rPRC9c92CE8wHrSlI8
LUrEcNWgYwYyt54HpwL9MR4THEytNJQG3MEHcY1brEneQsL7KPxufg3PVOb5NQVt
4kyY1roTla9xY6uPVa2x6k+e2iSBplC6vaFLdMON/ftmQjveW6KdO2NyCfur4YVa
XADUAbbGMjAbNHJM+yyWzaFjyEAeB76xzwVgsDEGJzGH//P/38/GGYpQ3h6FD4sM
qiwOdWEVI17oK/dZ6cFUhz2IxqHcJBYL/18Wvm8HDd2SovJ8AxAWfS/m1K+v8wIF
JDX1msW7GdO477pHIExkUly69AkEDy4anE2AbDEP6oUsDvL6UEwrEfAupJ1E7Jw8
p7ADcLQ6Wztu4F8Y9k6ExDI68i8RpWC4SyhuxNzZu9JT2qwcG0ALL+BdH2tMhVa5
egcdwnWT/9/7K1g6Lw2xndAgIeFAJS3fZslI3/4tDXuWCnQ/03BCQFwvf3jQ2444
H9qJWCfyMlS+HB1KKykraKRMcZXAmNQMNLPY6KkinjtvRlODiT2jL2RcbcdG+wit
c45ZH6k9tguSYCZeAlZcx/ThRY64ytRuE4QHQ/vORY9SjP4c22IRHcRqb5akRyIP
FZ0Hapmb7c954PISw+JvWEj9uco6hd+a6X0RC8eOrIUjAG/XGq3dQl8wL7On0UwL
OwMhPGtrcY57h1k/7fOhsaejf8um5N4H/yv7bmh03YrCfcsutawVXF9HaeCm2QOd
lpcs6e/8R0JteMh2wHdzMc2N/b11ExyGUW2nEB8c5Jvu+T8jw9dyUSZ/mnNremYU
nLMHYozyqtbZ04a0WW08EHW68ApBNEoqEHvieHGIw/gvoh2+lYDzylENiVb8wzHO
GbQmZGs3/QyRgZ9wgd7OVt9Mb4QW3GJh1OaQ06L7sDPvcoUBjcm5nJ1ee0xHt80w
MXExm43dZrXBf6l8IRyR+1FR2/U7CqHgBLUIum5jDBR1TtAvLEbNK2u1VJ5gqh5p
oEhR4FXdx1HeDorhHRb9KMk/Iqiwktj5UWTVix5/YBjrjUyHgxm3j7mQljPS/dLc
jOubJ6MIAWPhdX59yA59TDT6BYZ19h6Gpl5IdaDqLolCSulOAQ9MMVJbqraglrve
JUJAjjrkuDZd9vV1kRUO0OnIgEBhf93nOw+ukxcaQAk4eQhzgCCLIyonkmqI2er3
oK6+hcCPlNJ2QIXx+I2KXK9jhPxGvDMNtUU/4qn2AXwgCkdcqSaw35/iGfyj4Qkh
j1FJzBdr+09i3ENaZ9ccdJwLU3uBU8Ed128WxzmvnQYrCXQDy+RRUQJTLVSvU9IA
yfh1tZRG1niOJIpD2djYtDJKgATrXY1nAWjF1NIJXYl/h1Sif1zi+HUAguiZSVFc
kDEzffwcCa6cb7eykAmAVNTaDb9fKKzVQniEY2tU6so9CeAa60EKAy0l1jrwbSIJ
G/xeRz3Ht73QYUjkG6AJ4TumEi5uEmN243p257mzp08fzHD9hb+5ors5KWuLUZsw
4scSVFz/W42nE6S2DIdd7IHGsVQx3RRiDfrygQEC4werl0rJNgnkQI0V6/fRce6f
le0RMwMb9xfDUtWV4OHJhc6LGG6THw3S+OowZ9ef8z0EfKHNuumQ2DPcywBC/JKj
rGUJhFRuXJ79C5RtLHB0RJVQpdh5aieklSIWd286t8WWeg5Bu6etihdRWG5cNCme
GpN5bhhteqAmZAcltd/t6ZWVBs7BUOKKOrJDQUoUrfup9SdJhOW14uL5Wn7+kUkA
5iS6Tgb4hF0QkMlWyEwhAYy/FYjZgOjzGo0SUTB/4mGfS+ApT/O3BCPUyAxmow7c
xZhJjd7GSt9BT8PefOFK8Vvb3clFh1EkF5GICYLua3XbpNoZaSkxD7tAgpwUy0Az
TwZfFl+Qb+9sVXRIZn3lMoZ97cirOsQithkew8k3A+4=
`protect END_PROTECTED
