`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Trs5sjhDPx1gHGd1oSs5QqUf/LktS1esiEMZD4eElXDUcrz4WUm1Sdm91E9G/EJF
01nhFFkPkHBr2+s4uQcAM+j5U8wuRFERAL0sEdnsWTwBgnvTQjRCVfCBntGA5OQd
nWzS4FM2XW7QfnVeLcvcoTGPAAZs+1CuqbD/Mi/gmQra0vX6nRc7EVILiBxVJTKU
JfzqW4Uf4XaK6YY6ZqkjrgDeyM7tli07lry8MHYXddXc4MaCvA8+b8ROKzyurrtP
+HByLd/d9xGbEz9HqozcdMHDGGGrt0M0H+4w4up8udWfh1e59g8IUf2cg2TEQvH1
FXBkxYFVFGPTULLq7uznBc+UrXXtAXGmuZjJULlBuLwxhe8uDtJbZG/NvscCFuTY
/XinhxXsFTgINVqFYvFqcXHrECGug+hhS05jPKf5yWYPly3G6VJNSvP0MbFFxbdJ
3Kqsz62VIQwg0In+vtleWwAxMQQ414C6bklMPih4avk2yIK92h89dLy7culXCpi5
ilLY2PRiQ+F69xrO7Gu88SwsqsyYPRMKBDJLMdofyIc/8d8/ds+bkPKSE6GBnrwy
ar/uS/pmvXFdsxXr+iOr+NykPy6OaraW87a2Rjk1oNh6g72wUJgvo8s1zdtUrACa
gXkd9b5HdK0TJj6rIBYV6qKT+x3jSUGYVmcPjXQtoVNOpQblukAmfqsEIMk8mp9A
l3cZrUWD4zsL5zEiG55xDvjN7W+ETw3rjlQ14W+rnIGSP+CtvUO5yCmfwENk643u
MobVjum3DfjW9nwTKwfAZUVrGSaZ9d80M7JDJ7YQpP/0uArCcRm8EpZHCavW0P6W
j/fmZX2S1sP7Sceix/3kL8jV2vLCW7FCHIAfI/IDdnxrWdhkFhw2Kt4suwhzKESr
mu5FDY/W8tYyH945vOKVz5fl5v7gRpcSf5clXLC9cmNyz26Us2TitdFkC9MP+aUf
x3up+5QngECRB3yPtIN4Vgu7psubwMs4XP8lx6fP5fgZ8qqOm1aXAdtxzcilid82
wO3ahS0L8lODqvjQKx3UDCITspj6kBevOG0VTBkTbHbNxiiaEDgxWoczrsD3Elo4
oKSckF0zvJ2toPqT0i75vHXqew+06s7WpMy5cdpui5gZAhrDSpFJiW22iVCcD7rw
6+c2FZ0w/GsgA/rnqe7ocR9XgiE47Y+C3WluFbxWn7Qz3FOoBEYMTNyA94fzW5TP
qwX6NcAQSCm/gb/Pju+CHm6mrwUtHJrV3MaAYCR0kcDHduR6/B9rkAu6eXGO/XJ0
rdS9MaaZXo7HTPffrdp6TP3pJ0W272COi85guG1JFTqBujwWtj0arQGPfLFw2aTs
H5pGthOEQ2yDGW/JxFPlSavvgL7tkddMNq7qUUXJ9mo2GNt9vwtkyW+9F66wwDPG
WLli8igvDtYF+qoSLNIRuLaZJl8xghApSy6Ysi6f1qtPhCdkj4roaY7hcvhijmQd
5IMVSvhCA3ja6a0eiHD1i/7waaZ61124Xl0p3PkGaPvC8y1datlZLIhlCGJe92rl
xZrDyhPh/Sm18Ul54idMlcEYA8+rf9VRYz6uOWVdZ6wdYL+76ta8XNFtwxo4Ta0B
tDTrHSIAl0CLlobQK2kSIButHFUT/COh73/JmJ4es28DnHZ1qAlfR8QHKewzJ2Hn
XpwEE1v5gABsYlZT+NsndXT7C4n2IM3b7C07GdniHww1pKoquBEzNNXBv1kYbEh3
BZu1kmI8uHBEdCDohdgIrs14K0LoXo+7abo1yXIt86TbgbWWOhLPQjeZHCKb+9Eb
XrwrOmOkYqnhRlip36yARDwopY74MjaDMOK4VdH5uv/JZuNiNe4JPE+QM3IzJcpZ
Tb6DMd/eGwgluPSRblHwiRvk2odbWo1y7RFd6Os/Go+OqG+bvj/NXxM+geIPdj8e
otsZ3/Pg7rCZ2PNGOlG5oJ3iG4ay249zQ1XBUMCMFnDyk2cVycyfGd3DtjLnGyzu
lhOliCw0mXWCJRi0yWKv32IVcEVK3wMt7K0Xd1kVO7tJSinlipTQHzeOH4expyX0
YlxHkXNZj9sfMi9n/bQXQGFdfziwyODOOIzkhu86L2OwLqhfEk2BzCQu3kuIQHQB
JI42Gqc+77t1n4ihfXBe149+85ItZvL0vDp/JoLEM8Z3I2UJXDSzlg0dI4IHTd1p
zPFFKRlHaJQeukcWsOB8i7QZBGjYQTuJQqzAE22CJyEbo/Q/Tq3UTceYugDy3LHn
0Gldj3Dcu8tm+2djBB0eKqiMfoI8lmYtTs1e7xqjsMoWcaajd6Nm4iFCry9xB00o
08bIs0MZvetAv1Z59j9RLDjoZohueZG45nhHWUhurGJv850tZ9yMBlv9G/Hl3iy8
PpnGnH02h9hCfuI/RyDChuVWzd84Kz7BvYh+U+1VXfMbcKKjdR0gpDp2BWllqDOW
6VV014juoEb+C3Swr6tyiVwNDOeEa9YLw3vpEDGMZPgzQjlF+Qc4aAxmtKyFDl2a
BtS4MrSf51OpXngLWbbpuO6U8HtVcWGRoYMYyGZzwBjBlp+eUZpvyqNNZ85ebEp/
XRKqycY8gUyGJyu78jJW/zMISCvByui/h/VV+UuRwAur9z2jYGOLQ/ErFUyPTJvF
1bQS6cJp50/umoGjv9CvK2s1mKjULZSDzH/jW9rqXviOP1JgWBPDIJBDhfdkVgP7
KSY/q0ajv1xJ4HYF3FG3isCqW1BjcZ5+gIGaYuVPsnIlTWLznrsL1MwypRB6Caws
XZhBfi4sKq3GXbF/auXYdtefUIMwHxaxRRlTrPq+uxcxeYcfN9w38Nqac8CeHmx4
jmMIggPdodkM/Cx5xz2mzuQNPGZDcnvL0EJDG1EwonLj3XGe58Bbt+chMs/0tU+b
9BNKRY3stOQbgp10VOQ+aVI+5U6NnW85Wb7ZiQQRaNEBe0qpAYIjXui+F9xhBtp6
zBUASkb5lw02KB7PEtidyC9T2WuUK5DBcOnXjkbdDA97AIgSi2VNw7foPERQHquT
lA3k1l3GangdciTFW/vE62AMor1fOHputtq9qUL+46F1jMP7QnxYIrK2k6cFwePo
3tr1QxfHa6vl3k0wDkmozJ74D/xlxPGEcerMIgomG2FtMZ8Vb2I5aNh7W+5KLIgd
4joW8v3kMTbD0Elytg973ng43lRYFpr3Zq1uPVZbshMA4Gghw0VJ8jul8lx5kBKO
HZBZ6hJ0493ZLKyBL8MDfaQE2UNNGDpEskuxglc6I7h+VrfOBWgkSkH00U0mQM4A
Xitw3mjXlXSe1A4Gj+QAynecvdaIWLR33JMbABVBjCymiEqK9QiPyjRiR3QcWBhy
dUUEzdOOHDLHiG401TUvUkkKdCXyAteiDK1oaBoxICD85wi7CzgwN6mbz4YuIYIe
aKe+4FC8Bs+E0BgpnhE8IqVFpfSyQoQRyl/s/MeEb/9RE5Cb8alVWyr77BwTwCEQ
w7H7I65v6sgrvMURkiqOeXlo8PTr98yJrPy1XAlxMmTa4GaVXOWqhxqkJJYQbWUp
tMsLj4N1fhpM4go+dnlrxvBX5Or9A/NqLnvTm5rv9OA=
`protect END_PROTECTED
