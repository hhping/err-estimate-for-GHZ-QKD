`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oM+ph9gTjbZWkTOLCnJTAsLkBHrEskOpF1iJANzpcU09KNUHaWXc4e+Ce/jWAJ4T
94mU9qnbg8UYfpeWpsJ+FCLRVIuqfU179FuHUB/WAhdqhuwXFoIWKR0imhsH6xkC
rWTT1fg94LXsf9TKF29zi+haq5jUxRO+hu7B7whDjtCs/JFHOFY/i3iQ1KurNl74
ujX4vEM9B+Wu/WgpfFPcgCLr1Z+gWGB+D/KiPElfmvO0LauZVam5y57kxXmyQjLL
fKnzCIXKqT3HvqoipTJ6b7BCvwz6jerUIqgbDz0LuVCUuUad/wK5Tc52tl/tO7gg
d5OQCc/GAxlF9YEV2Fcj2sHbVItrPU6Wug/ralducuABKCtXwDOI7Mc0LX/1T+8W
8TxJjF+pIYffs1ylXW9TuQwGcA+SVEVfSwb4/r+ah4JSkBmGK6wX/PtTwA6FTs4m
gLq55MigVaJm53lx3J3sAea3V+7r+JVCgppUklt5n2ncV5Zqk6SsWTNeie428C5d
bDSedzZfJRDf85EKbiZzpl6sBXwAzvDLk6JFLHAmXZ2YNjWL9FI2H5pHQRiS3q3j
N8nUWOF4k7SmHBL7id9cfM3Iw3ZFL3JhmDYR5koZO6spAp/FHXHhSo9EsnDCLMmY
XiI99bGyIZZQTKk1cajipGlQ7rOPvUiR2S08B+EybXo0Hm6+UMF5jnQQuusKle0g
Fq7Hb4cBYLpWL/OfzbRbypSIRO3y+r22aUJoHHufTqDrl5Ov5FAP/ebN8PKRzQGQ
jQ9KOsxQa/VCfrCSnWzyYR5WGe0/eJY8S0FqpAGS/n0WsE4JYafJ9ZyXcAnxmGXL
s+xpun4NT/R53NsFh8VnabdbiQmj6KHbm/hg5tFYy26SSu14F7SzY1vdYmJRPfab
zf1w2ioPrFBLin/vWbg2bPle0VeVaAfst59DujYzW5/824OVi97DNbR07/X3PoLH
aRLk+iU1f/A4Ble3BPU6atOzYwmUIClrSM1rv1YHzczvBdfzD8fefdnlfRR51YAF
MT5ezsvoVQZ9YEFUbidUtLWvN0bwa/oG69z/nRjVygU7aLXCJNqADmsg8alJ18mx
rFkQqEsZPjHlFQmrHCVcqFUp0+PlP/ty1HLyXE+BYnFnOb6Sz4C638fPRBDuAROP
j3WxcE74dPOh2hoZ4t7Y5I9NgM6JNXbvrTfcn6kIBMerdos7v+Cl3W3SzeRIso42
Umz/ARDLLGazuiWF0FgJovb9CFf/vefBRyID8QS+6c/Xa2cU4DjuuoBuS7QHN0tj
tW+xlEdJUufRnew3eKDT2kKHuMT6NZfmzRRKgGZQSQNnyrnQR6RBjyWR6jqd3vrL
1bHbhdYKPPRErTW8DKBJDV+xuBynO1gVUemV5Vr3jJ7iPIw5t/CUicN80wuzQrHx
9SagYevIqUpfqcTCNN5XKvF2QxBtV+04a8NxU+LaDI53keIdV5XGr/ASqVZiHHCz
4JqrUmWpnHP7qOvlIEKFwBF3BTJSpx8Av3ax0NcQQ4qiHoowQbHKlaraKczADPMK
ynnE1lVA+Oodon8uUBYdmbxgLfigMadSJDJ+WPo/1OJcApUp4laQ56ye6BMlo4Ot
w/jDmwDAvcWV1HY1iXxSnjNNxQ7qkHjbVQAJRLI1c7YTq3knAIu4dwzXdmXR6CPm
qZmjnvwfKOCaOWrVH1LQU931tGWOwD6ScF7X6UKzvUZ5iZ+xFCMEw/6NZJxGB+xd
fBoKkdE4dRbSZHzoX5QL0NxxwxXKcPWuJQD3GmJ8V484OatNVuP9sN/qyWVJyxxD
/WeFheHiHokp1jXNSIFKjg==
`protect END_PROTECTED
