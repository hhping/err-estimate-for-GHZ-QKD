`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DWKMsb0F+/WT3Y3hdXmP9wYnOkfh4yh8W81ZVjs1LGxm9kWBcKc7iX837jBU+/+g
UVVEqdBn47cr5124zC6IpZ8hQTbYs+og73LW2IoWgmBNc7yUkxSP+hVdpFr639gA
BTPuvzuTuHYKBwLEhrE2mZIDUdq7jVmQfYxrIU9XZ2EX9kTLxmXNBmqP9ZHLlzVJ
maz0/Ngxx6tJTKkcItUz8meVk7K+Z/nJIgawrkpwXVxTV8fCCCCV//UN3eEpWxvY
J76X2NzuFoOqBmYszhB3aJFwI/8E5qHW7nC4cVKZ50EWAn7XrRZZKLDkAUT9CIcR
QXVY1ODkvBlBf1yd+hlJFHmaoF0ZWxAnnEOiQiVJ2QcH/JrheMZaRjCmJIBGdm/5
8yF5pwLqQlzh3z11LgokQBL2ggxhSwqrfS+D7FJk1PsQDJE6KbSnwai8LxKuQYhz
UnSyuUHrhzWEVNylBwWBeeCcLX1RZ0pU0cdw4U4ivcl3hGOTQ3Y2D4BUdLIy8uL5
2vmEYY9s8n4lEHtN7obb+3YCvu2kv9JkgpoXxI4yrbByFaCT9CDzgkSbK0xle91T
JqtGFyZtqeLsBn9gjksgQBKlewQLizMZwv1DYt3qrQsQh/8OglYrHpoo9ECuUeRj
`protect END_PROTECTED
