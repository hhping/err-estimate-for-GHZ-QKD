`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FJLTE+0MgQt21map8DNP71t2K7k4nY2YLdTUSUhMTbyciRMjPHIC2bGatnrWDb8R
OCIRSissXe89tO0M7noclipKd+MtzdWvZ+A0fIuEyt/QbKq5aYM1HVLTKDD8mU4z
vUiErmdtzP9UEgwaSdhOnv5zWHzRJ7WzDOck02prQf9YMZ9BRiN/b9XROlVIGlhP
vRgcJPYJJHcOOZnuSvuwGAYLzeVUIXIH3H9uObAPuizYGYQleFiuQGS70qcZlvZs
8eUUar4Zko0TrNfJpXPRwop4WEcUd3mT7P8zbcvuMtLQ5ClucV2TX9P6t+0rH9sd
MxdUoTzSLorhIOekxCqdk8SbvZB8emnJbbghuQRZWHJ8uQ97j2Sh/tXjO965UDuz
oaUZ0TtQUa+lp9Gyl9AC2pqLYff+mpj5wYDRc1z9saTTtZQXTi5r6FFZmlkybpRd
kF1G7EPWvaUMG/LKVnFSRxcYnZXYXPH9PZtb59ZhW/SedZNLN1nDI5kq1BGFULkI
L6EHp39bKX9nWqoBr/NyH428xPYvt3mdK4qHmtqV7U1tK95FOYhcDNQaSeudReQ6
qDroZvXInrcLo8zE0oSJ3/qzJq/MOJi9d6xRZAIAzcZMyR+gxCAW3XlwN6WPv58Z
Z+cPMSmWtUSobn6r58hYe3RDuxu2D67tcDfY6iy8ernQYDiLYY8AI3Cegsu2V1CD
U2GU7/M38pZMxmA2IdjAVZXHO3jI8WoIGDPSsX2T1/29NB6K6a8kG7h82Uk/SEuK
nDAO1K4s1S1Jip9/6uGrcJiCCpW6aOcWyG+SyTvonVK57YQbCPq0zS5vuK1tmic9
lUzi9eqvyyCrY+OdQD1zhe9lD/E/sFOR1+ejiGqs2qLPEam3VxHW6LlMvfr13f2f
5fdVFmmV7l2wUN6XDfN3lOCv64F31ZJh/pjJ2fGrxgeoA7zXfmPo79uKcHaPVWbO
irMVrMA72bzSOCxFW7OW1hKc3x7SeqqoGKvFPuXeL29seg6u2FeRqEvAAj1rm9Y5
BTn/C/NiGVZXkJfkUDa0HB911R2BAXCRrCSf6pTtN6v+i8yCWyQTBxPcOH5d4pu7
MyxGT+8+NnyP/LfShCTPfg3B0uOycIU/rQqZfvEYRh4mNwE2bx/l6bT2gfObGVij
VzbtWPj0UzDSNXyo+HfP93XQi29ZxQQCCT9IuL6LqbPBhOKQSarCFNfRxKTLDBUM
elbuM+EnNGfKTICrjwUF7nNts6eXXkV1UQ65wKZUKfPN0RtudV+gE5UroesqX0wS
/f/T2v2eiHfoJzpIcnfYlEVIyOtTMX0L9c/fI+4UXIzOP0YYWCCHqllfhytPyeKO
JCNRnBor3BvdogNpVdbI6/hnjqaO5BmVQ0Lb5DienTExtfGxDqRv8YzokQfzDVCY
mvEXYQVlzfsagnhNRxRwoplMifydcE9rPT9cYEktJNg/sPlUXSm3omjG7rUqjT3T
H78GRPWJyrkhBNe9ZIDmMnlf39m/bfJTHCR/11Tn4J8K/mtzA3CcHJ7ObRr4vgAO
WivemezhO6r+Jv28m6NWzdLUgeL4rhbLE4hm6Mqb1UyWzzQL2Y2I5ZXDFfEjg7aZ
+zrhG8DPXnh5rXUGsrRkiO1GxHjSkWt+b84FEF50hmDYXTS7h4piYGSSVbHtGBwV
G2spub+RP3w6/n9GWDdKIKw1SmzygwWwrLl3gD1kOHr/hoyasRpI0sw86NJOAGW1
vEIZs7w9d+vtw/TmtiIl8huFsMW19yr3xnqQqEMVzGL5CYg78V8cZ7g9w+hq2JW8
Ih9B+aNe71khrhnM/9+1ZuDO4BOMh0k9X7uW3X91W+3wLa+XCTRHM8wmt86eR96S
i7SwpiYhyuedkbUAfvZPaqdwV6GXqltOilhjvlHGaS2EQ1RbQpW4NWYo73QKZZM8
fokkCs//m7omMVSYbWemsOkP4t7KbcsXYCnBZ8UdC7TWRnFn4NrhBMHS4n0op5dt
085ZMCXxuSwZbKSdsmtl2EBv5OVzbx31uiuI5auGpiki5bRMo0xYHAT8oDbvuRMY
oFEr+MFEkg41S9gopTr7QLmswvHpIvPhZ+GpbAfOOCpuNV9pieqjoMZTduS0dIkl
3wPjpP7C7enD0+ChII1UPeo6Ly5zyxLX/9dt1I9bNR/ieeud6jwgxQ5gFwv/uJza
3wqJnkc+B53OZBZepk2x4w5h81LV2HnaiFHn7HyDWeEStxOn9SthfvrFRKmwMD1p
gyOZJ1iLBukcAYywXKWRvw56fOBHga+RETPKyIe/murWhi+ToH2vPyHsFjWWmYUN
1aicG8+ywZJ5GYQJ+uXO3jbIeWjG0IhIKLNW7HmCzHyonvzPZ3+fJZwafrCjczBQ
BwluhT2kFujB/O4VCRp/rtGoGNCWMObzgsbeorAqzkjhPXa1ICYtriB0P1qw088/
MqmSFs6Jq8prwMMoDfH3yZNixdkrANjOCuG+1WIlUvI++oleUva+s5yv8uwcOob+
XEbTfbOGfKLDTPNhqE8JS3uS9RWw5g3m/Kn4ex4+LwuRcjRgvlyJtW47cB92wDcs
yiy9BQI0Qahy7HcQAE+F90vVK8CFKcHx4V7c1vcSxQ557u0HcI/CyKdCPVMzmpsK
TvINtGYIon3V8D3OU82EnGfpprau/i7q99OZqVES77DjiAOaH02xzeLs+6SoXCkz
uw/aDZeB//G5QFkmlTYpTZJHfgL0NNSuBkotqgpGIubcN6MBjqhXeGzv+UROHCZc
T8aFLbexhPYj/27f8ei+q55eY0VHg06p8Isn7A2fJXD6nprqbHq05hO4wF3mbQwn
W55Z1vdSeEArGUMz9o7Uv3oTvrFTVgH2ZG4GfFhZnRhCzdFPzPQIpXD9uwpmx6+4
7/PFbl1lXkY/rrWgBaPSEIBUD4ybncOKjIWbGI1G3qVGTPgLF9+vyuXV4Ki7GxNE
tMCUYrmlM3OEUIM2Om4aRfONA00Hj6UZx65kx3Izflw+uhz8pa22DaWDFza9kEPW
vnwzxksAqgUYn5pGpudHtjjWs/QCACLx0Q4QbY8yPASZNZgl+T+itsulFxaRaaYp
x1fFhI2FSl05RbOK9/wB0S1rpcchp93acyYDGx3SQ/JYbaFoYL51+E1hPFT0Bs5V
uiV2TvtiF0N3raD+XnwuIMVFLG6vM53ULEs0/ZoAvlku5ySCQifdIJlHhguPsAsu
tPPIdTPz1u0RAQNSmsmipmhGkGr2/+RmXN4SMQxEV6UNvHu9f7eQOvMUYHy/dIsP
M5hIcEOUDpN+LlZhw1iaWzh8roVz4XStdLtAmWJB6roW3BDK2ogFrQQkB8Hptz9i
XTE4Yk2t5KfOglqZ0sU5pesXSu+htuCcPjwO6ofGH8cknOtooWdnyv5RYphh42Ax
lLMaTNnsU68kfzhf8knS0yZ42p8fpa7mASdE5had+v3TPzfOeUz83sUzN/qjsUdx
e7983aUJGoQRKsYAV3NAnm9+4OcI3shKszDXIjs/W2dyEzGeKtOH9fU/Jx+qRJVT
yPnvn51f7EWojAhE6I97n57/R21fqmHUt8d4FYrQa6g5XSYo/S4z/yyt1L+hG3lp
93uQRdkypHq6QhJif9OIUqFeez4Zu7LHYcWnb5HvGqpv+Ep89o+B/nxyI8Tr0fHB
bU/267kk/+WFID9NQiEn+snAgwfrQ8GNQQfvLRPk63fQRNT/9GvouiVd3yR1W8RH
bN8Wocotvd1m+fvN78ECiFfZsKTsRYgKLaWWjfmd9RRZXBeifWmkgCEREBT5xaK6
gGB1LNMFka8raqjyGKE+Ij0YS3I1GVRgyTDVcu56NB2l/pNUY550SiEGb8J8oTyy
Znu3UhqM16rlB6vurtQyc9cPKSavKku32/lCJCq2EYUxsZ1Yib0sn155Po3SHkvI
SxTLDPC3wR4LyS1bSr86jzci86xjdlt7jAffqbT/FDFKuxEqO/g7ZrCdRNGcrVAs
I/ZqYksT/Iare790vZAzMqeLe3NU7+F4zKX8X3afbMre+jGqrUtaF/I2QQXy2Yye
nzdvFfmNX8Xi5qxm3Uy+bIQKeuJXKQqyNcmsZOmFp7g01UugjIcQM6MeIcW70rlt
XmulDivDymW5oBYzFgHbOkm3jSien+b3vFApOGnbJjXoQm30/dtcT78GEka11Tpl
+rEvHuTPcJGEUR22DP1wOd3fCN45gR57ZN3rDs00WrmyLwiR1mL07mZ5eby65Mv+
yMZWkS7ZJkNHlfHsFscPDTshIYyJCBPnLpkSb0nlxOD+b/NJfcXBMyvuk3KTSfCm
+GIe83kF3LVTyBincR7k1eW9kUBKGE08P+njWOfhC5hCQGT2nKYUhR9QKOzp+9/H
La84ZVHI9gxEjMAxiH1I1QiWfDVexPOkftFVEbvo+CsMgJY1YkmfKfUsH7NNLePR
UFZkPcGM1L2wmVvalJ3drATG5pSqsFMlFqeXvwJ678PVLeDFPaO5rrwpqphgNtmP
Woz8eFbyGhnwxGXaVEIhHsCKbzDjnvVxR337C6maYqHdZDuAS9rUZrZlyXZDxJ3q
f8DXrhkLnryVE3GkqWhOaVVCrF6x2XkjOD9MzhFJJ6V6QOf89OsaBZzGO1c7/Db0
PpDCYLvp5/qkBY3Maszlhfs4zfTyCFPtrPwEfg8TLmiYlSZrLmqyGXYey/1mZtLt
qdMZ4e8nFZD4hJJnrFon5u22CgDWb5kOe0Ew66uecrBJAbZKpVa1YObCMDQIDPoO
kadSCSQbbbzsXah6XP8kStbBwVnsMp/K5akd6f8mDoS0EPYI5EnZZ5N9aNJzR6Pz
e7OK9VWPjYT1aslVuKTq6dvA24KU3AeRaE9R9z7bu+N8EcQlfk15x+vVOzQqyGuB
9iS83HKa4q9Wzd4UA34oPhNTkbXk9Gli8Y5TYJkDnkoLUEvPRG72gEpj0OWdw+X2
Bgj1PDmV1zVs/DUScm71rri/hGDYhlEj80lJh84yjloNgitNmym3y9UtFKdNzqZu
v0BQLtepEEfvvLjJmQGVTQ5iyj7GXymOyvU6CWkslNfhCcONr6MWFhZVzjFLfc50
JfapJMrYbfq5dygWmsHDiJVIXPg+SYZmPHVJUoQwPFYNrjr/5qfvkmdcNrvQ8qF3
lrq+vosW0xFHZFIXAhpw4BIvwz8m0puk657dhIdVR2ahSOevGdFVvxxfprdjRDyK
EV2tAiV1BMIudYvLp7rHIdASkMqnUzs6lkaqyFAFsJvqSpvWQhpYzNn9YMgZMiGO
eUXv4twCmReOZix9EhijS/Izm+1YaDN/zTfJC3KOtXLSJgG9ykt3iY7ZCo3PjPiu
9LiahcoOCvIUY0qU3B5y+4baSD8gLFpc8XoKyWloOsYCN23mb0iSjkUXoE7g53Wf
tVS3VsUbn7t/0eBlLdJUpNs6k37hsHgcr57KKZnHNmqMcIYz2wTytNK5Cf1qj83W
M08gKzwVKbNudljrh/CvThVACdDHXBXrIXcjGkGMek21cl/UuggpSGf2jjIQozMV
HRY3ZvCsC8oxJsScgPP3/bnXQq7FqGt3kPe32vV2CwvbMd+Q0AeuY4P1QCFz8gRq
VBlUSWzZX+Wfmihjamey659Qe8Wp1P6830HyE8Fjadw15UEdnl+L/7wdt9fqY9+f
oa9Inm9dJjDVbe/NCmNLwER9dAi7Aw5TagkqPZpoMy3swcW0EUGsICMwMAcaIt01
2VnUD0pa/TCeeRZ/kvTzmox/qFXLtNpcxHeMq0svMRNntA1kF+f972l+LISNA8Mc
1IV/PH2QDGxuuhJCgaX5xpLKxGopVJjLsTHewlLApNw1mCROKvgym852Gdy2xUSj
LgAaMLZt5BqySmCENm306SeAfFLKHFhPOzwepGJepdhNwsVS4Y46C7nPZ1xJu4Nc
GfCvTmio7X9i9bHhxrAcsbP8CgpLZo7O5E9HdWawYetUSsjZRCyQ8NzdlOmWPpLi
JcW00EIAbKwOYcYUlC3RD3FD8b4ptHRMCt76MAjwChHsHCKf1w2vfeZVHcey/o5F
aq0ekjaBgBHpv8TeYcjR71oz9GixROTxZghhudqYQxESVYDQyKjmtnAuAd26ctKq
+Z5mEC4B+iiQwbgAdfBUhWnxKE0iGPP6qs52UsSdduu+ietYORrIcZ+CxidQ/3Kc
lIhuecQjLjAsHDn6fsIZEmbYcXTkcWOzqc0IwxzFzrEBAS1FuVYCVwCqwqVF4ZrZ
vxkWA77jpO0yDoImXTm7uJdcVoXs4Onxm25Sjf4uPeGclhzun7+iBZZViK6bZWDI
bA83Yzxtk5v+ZbBM+jC3IOSZZWDBZFBmvYOuaDsT7/fccvNMmIgzODtgoBmFr8zl
2nIkW6I0fVKSBSjqB4hiONT48rltWpQt9NEzyfHXuNqAOXcp7WHMsiASLHPW47P3
Bzf6A6J4J3SblrdGvKbSlgoSY4OirNNpQPlRZuKQzX2kzPpEwubdl7LEZH5lJDEh
Ka/Fkusj+4XFbW02k7qDHFD6o+dSwzc45cvDRmzJh6nuDUr728bmyIKkj07CrWIj
9qT/eTHPgjP87kY9xrsmZCk5KR7MGC/kCaxj+baD22EcXs4/XqjpxAV3imhCbejk
5nHxi2An+phoKjdLGOMt9ddLogZ+JC7ijvMXjYZx7RgJT2nt/dG5jEJY8XG8iOsT
eGURv16uNl04KE6V88tixJIviP5Fb1LBE8NjjgsI2Nj7W3joSBuKgGxep8qIFheA
Lp3uft/fLPMvRBanFvJE3qd2ljBWAkbJouaJFFSF0SoW/QIJ0MoZoHiknGkhsc8C
F56FQN6947ywbgXCkdhgiB+kp5rlbpAy0pGxhbBWLYTrgvBDOUQwEeXoU5/LsBTK
sa5xtsbdfsF1GYkGpVV05yxv6QTt4vUAtym/3UE4Boe9yzVSWY89oD8ZEp8fbHrD
FF57x5gLfkNPRrlVaIoS9hCtYIe41X+lpUqfdm0KkgyAwYllMeVSn+Kz0ac4TLlW
J59yBhpjVm2hZJdl2Yriq+0wI5GGrX/fsQ6pRfXRiqmOb9HPEl6gdbeEaKz29Zwe
2U9bihMbHGaBMM65wQpv6QKe1NmNk5sijzg9VK/HsD2Tw8kdYDjjoZfmqE9vLb8x
ITGdY/yZLAFExddDC2AU9juWE9v/f/FxRtdf6j81ohXRu3ng8xThw4Y4dVf1A8ps
A/szLnBsZHpmTEWBFXadd0h7vYYymJIvCF58UdsZNAsdBwgMNI9f7HfWIsWgHWwh
toemiedM21eXcwcFK4xOA1gVIuVunMfPYCJrWfsFYStm7FRxpNKTrFQpk66XfdbG
hpT5FHYSL4QSV6eTE+IePfHG+g+DyDnqJu98jjcHKtW0gPNmjotEOLuUDB6RQkij
fO1FANd2wNvdcMDAGBE69yr2gpdWlXPzCEupDj9n8Aa7nW24s1usDyVsP5UxWwD1
GOtqPmwnPtUdeOrI2HG1SYSdHzxPhF5bmedmRuKMlAQ9ZAzfdK2QFCJ8AMHA65pX
SFaR+guYfrKiFI77jkjPrcfPxZ1cTSq1DWe43uQWKM1vmvrwgmLEN24xbjmsO9fX
XZyF6KKoga9nu315RaQExU9eGbTLUO8uVV6WYng5wRMLuemV6HwbUFQzs7XXXUbc
EEgjTRhaRcIe/6vXPfXDeILRgjhm5NDBpornAXagzv8Lhcv/oE6YGTahxfWKwLwp
vgPfG/wykXQ+5sfzyH5H/E8E6AGuaprAYR5fXIeon92uKRwrvG3aqQu/LY0lnpeI
LV5T9hQ2J8W53e5oazQBlqE6zA6sc4EGU4YRVEEhyy9eLutXELxPpsuMVSGv6+CW
9dtajAKpN057WDeB96cNVlTl4QvagM1h3KkG1Hg4nTlshTsU/zhBskFR0dYZ3isF
zig9s+d0UkgRgVc8+hapmJSK5qbFy7X7Db9gp3gv87NO3gxE0xw8fGYseURHk/zo
eszuuPFAn6CoLJhqG3VZ7fL1eoczmveoQh7fQKvFmsNC3XvgJ5fG2r+i0/eKvv2F
49ULk9SHNWNl+7gr/ESfng==
`protect END_PROTECTED
