`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JT6LJhpoc/HVTVq+svNQSmNUdDDra7bs073+nMHeoHLMynWyB/dAiQz62xVY5USq
SgZ7eY4jGCtXdIUU2mMwrtuNLFIqOtLCRVA8JwxsabtA3D4ZwQmb5E0OG6ci3KMJ
FY+WvN7Fhy5zR3uSFcnAxK29BqsTpS9PQ+/mthASrDTitbqrVQJZ8pFjTvCG9b4m
t4mHBvkm10wFC0B1yCsdtByabxDVad9ylUNTRmotzK9PeE+Hd3r39Z6s8y8UXI3Q
T/NVahSqBGL0rZ+9kFmxqs4gUBixzTYyO3x0xjSvbiXTiRcTOvnKsfnDYtDD7Nu6
m4L4zkp2mG/SEi4HzwMWaxECPhVZyAeVebz4d+PzjjZHJw+sCxyKdtQepKBTR8yO
GAVJBFvvbKC15Lo7JoWeqi7a4CpBq3Y8KITYHZcsDzSDWVagDc41pqUgDxnHnyli
B4GWCkUzd223kf0wiVYDNQfS7wqisWoY82csI4zkBQmiwsRx7fMQVf9Xar9N47Au
3cixQc16NzNmDa1c89WWeqgaoX3mllvzLmcYJvfnAPmMEai0xnYlGkiU/Cu7dLLX
MaM4cLDS7qtNu/YXIsXX1vfZrF9BGiWw+kCRtAasiXAMRn/eiYIEXghbgjC537Dw
LwmhsklfvIvzzl7W3PS/v1ZczYHHr19lletkesRvajuIBL6MMMhc6w/EXfQ+XDqn
EKYXECB3Fk37OgsFKkrgWgF+5AledH1grvFwEjY8ylgtcBN/JF1Y/PbC4G0nzlIe
ddTeF+sKDP6iAYYDMuCHvFyDvvLyPWGYoaZfMYzruBN2gNZy5eBVVHfGQT0P3Y/Y
LLqLuKs7L/UoDSDwU7859q4N+qJZACd6tO2u/e6IBJM/7JtoDaQfWatDCQxorrHa
xEm4YvBWS4k3jxMUQ2Z+yr4bwcCSJesF/1Rqa/dim6JS7CsaO0s/2/p6tcMnXQal
WC/0y8sgCRjBiQgFHmEuiPl69kXE3/UOnXdeamlbBeQ7NeefF2yPcBh2y3A+eC6v
suAFeO5P5+j6ANcALditoYhcPzCSJ0VW5e5X8ZVNymIGYL0YdOWDJh+7HLfl1QT/
sU+5Yz9nxjRfuJI9dVxjPXeTEVUem7uP+1bPYWYOd1aG4VM91uaCx0S54iIfan7A
`protect END_PROTECTED
