`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8OfYD60yapuEabEruiHdLDf1Dnrehyz/XFHVaknttxoqRDQorwXfM8l3g5sLWcoU
rRje5kJ1TNScgh5wmNe5WHmfqL41aUpOvdOD+LQXKUvPR5RPZ2yZFH/wvCUIuiRC
XEkxcZvq89978WqmY5rvN/NXoiYxzFmD6shMG/bq3+1qGnH9HzSXW90r4NfYYHI0
3dDDElIWIrecZMDSy42gm3lQCQ/rhvLW+3lzp1yS9yJNGUijXz8hNxatfa78n6xE
C8mRhKq/DlxJyik00ilJRcBzBd83oELEVEWOrbFwgGimMnQ6YYOACmkNYd0BdyFT
SBNsiaFoWUilt1qTOXot+ZV2lOQgZP735zivBQT7UFw5x6baLUE1VPORTO+8eCZ0
8kap3OJkYuuH/sCiD/m3PHuUjkJUNfGEM7KiwEwYyZrlGas+TouUuSDfJP3XEC+W
rXMrJ8EyuRIqgFabGNF/RbPpfQPuhMrPkpoGkSyPv1vgsswP9MomM68FYMbhZ/ve
Vq5PbFpHnDktgu+O7aXZyLfSZ5s15RTfv1UIi1woUkmu6XNP/UXOsldGzqcAeVN3
Xl7uQT+TOrMEA7pBN54NQFzE2gCQdIoh41RvWT111/qS2KsC7r31JtGL3mWC2F6n
1CGZt0NM8L4jhNJo6nhmt3BBGKQkdkxhNgbX9tdfIcLmMiVZ8XZJcXDDVd8n+FyM
64OF7BqtO3pf0fc0xxRJJ9BWnjaXSwIm4N5dZxUvClk/l+GMb3rmDgYxjhgoSAe8
QbBE40CaOVGhtsSR8JqZ0D3pp3TloxdSnQF8oDpejmD8zhyO5ei4bC3jrHkkDFEv
9ZySCWvKkxDLoEDW2mQUoX0YRjv7bItpZ5hidoLPPA+AI56txL7gsB1eiplHGW3Z
dqn/CFcFhxC67UApKI/tY7MS7qJjBxfDESzoQM316Zs=
`protect END_PROTECTED
