`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9zCKWqtpyjTX0pX7heyOimNV6K6lc9gA6o58qS2LhkdpeoBCY8ODjCZBHNPbtu6w
iijPZhfe64+Jm3HvZ6updZKkB6m1bGNrYhjyF7bP8yfWIedIPXc9GCxY6hCGyoDL
FZFwaZlsEbjEz0WygVjPi+ysevGKO1EenCt4GV8ZsIGZrNh7DzJnnD/F7s+/pfyJ
dn+R9IcDGWWd8hxi2sJRNecci2TVppIEg3iFimyjfnWEvBivSmD1w0T+q+bQH2de
XYi+3zKjUJdiy479PfJaAJrxt9p/f1DXHiVo17iLiZmLgvXdVJAyXelcwPNohyJi
adX6Zt/RRjUJ/2QKzHIoOdN16Ou7G72rcB7qeyMEsdkUxbcTtpeFveXflz/hBV5c
ZVi5V+/A9PzjbShu8gsuBsjYGsElF6Q40dIjZx5BckvcMZR2iHDrm1uh1rkNQ5yv
hBUYeAZFSQM9x4ELulhFvsWmvlTXebUMag5KsjZjlCXt8sZewfpqVf2p4b3M0+Ht
KVCO8WmlNA6xbj1a8u60VCHsLuiin1ftSkhpdubiVwPyWWmQcbY5Niw71erWqan4
G7b/ym4jAntOyG7XJw7IdHGlsSkXU9Ox3y0Oly9ZpD+lqyOTAfbOJUdmZTuOeEQH
ND4QAa8UU9nroTvDe3VrUw==
`protect END_PROTECTED
