`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LcoL7kf3z2SeV6C3/lHrzOqWm0CO3WeW9//bQbQWPLZKHrrceGpeIZvEs/gqzwww
6wCYscv/oftM9ZHWdbuROcYJELzja7GOisCZzR8LEX4OXk7jdedwLoz3EmmGU3YG
AO4j3NlnNKY8kDjZyN7BrAmCeTJ63duH8vB/wVrZofn0cDYZKi0bIy3kfAGGuW2R
Ys38/eJZk2ukHvo+eM5PL34SX5Uh08gJ/3Uw48cM8HSzZi4gpKVlTlXXX8i+6JEe
/J2h434jDUgz71C4VzOy5BS20tou3t8yw9HrE+2RM+q6tAe78KuJLOv87Ty0fSkv
zi6nkZEa3BNmPLxBAZk8SYfyZaqJ1WjSTjuxakfDUNYDVsyCljAe/EaRojgF9Bye
6NIuOT8gxLW+4bbtrXDgfnEit20yz4+7Njbvm3Awm5bVGQONOaJv4N/XcHhptgdO
PW5rY/GYxIuuTyUqFu873jzV8Fmf9jsXFkrKsd7BC5x/9NGIMZLxjXw6LAJGBpvv
ugskjAJemH0/GSPqhZ0uJO5lP+nXLxhJ5tWQw2VEuOo8iQc6FAfkFtjwT7AjVd59
7Q9A8hd8IjmYxbfMMMNfPx6di3y3je6BRgrx+xqUwbZd1XL6F/L2CROgdRylSM21
KhTjiKng6T1CMZ1j+TQdz68R5AQk2/qhwXzSNatJWAmY4KVxXO6iNBChX4NS4gHC
bQEdrOIAzVTh9jnInIc6YxQdxTHPP/Wrjta8CYFF+6Mxr+VXeY4N5zzKPi5rUPgZ
WxQFoVE2ZxPfIcDzennwqHPcwSMKW9eODRwK/+GxTH/IvzjlGi2rKRh0/KMY54ff
riwgw08UACT3jXp6mA7wZur/eZxHNnqTHeMczidh04+H/kMCs4QXUGnaosFWBsMo
LF7ZH8+0v3WGJUn4UxsveOoF75safcW6uCxqy/YVfqQ/kqbeJcg1O3WeDqdtcJBq
GwXEPAWJ0/7h95jqNaqtAFYWEyNUFlUvJLGsW94IntHEDAw4Nl+nQJWhrc/1CdxY
MMnmJxGz6gX/c8gQ1a0NBUtmlNdeu/4FtzDyOnTGvVMvib63VHJE/BBZIYSEX5Ca
1921qEHYrGXGkojbTSUapl51Ze7gYyVg0/fJAg1n4S3yokciTZXrtQZQzCEybSC0
7wIjw9P7QC5bfO1rlNjKzSo7h5SPpjUSJhDAu3+3HFPJb82wkf2OyG57LGjFjoTe
yiQvmKocV9uCYGF8EUv3lPUrqmzVHCrG0YL5tMXRUkEt2pktJKqVN88+ggi4gKAi
G+cGp5wH7sEhg2HUfhoIRvUCOT2kA5Aru2i5jYoB5IC3iqPR6Cl7kESbm6EUpMfi
RSC9h62uSAo5B5hQ0NZn343DRGleK5Lv51SXsRooi154rnwTtH8BYe/rypYdQRvk
PiVmgkFH9oMJaWqYB7SLJ0V9u0Sc46GehsBvvIMu51e19lERCjeDXSCrAdei/wiv
4HnU4NtbY3aFF7dhFVWIlBIRHaf58CVJQSGZJOANouGX+2eNZlsi+kKx64WtwfUG
MikGj2XD6ywYeDH6tGuFbPRZK5PXsEvPYMz3xz48l5krKvxSs5pBvEWZRWUdnY7a
DEMBOm9WupCfc9cZa9Z2Ww==
`protect END_PROTECTED
