`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eR2zoCnqQuI8S+B7rHP1W7rcalpl7xn5GHIkqIlmDfl8j77XdyWrHQKMPb4RcyG9
C3/K27GTkamI6orURvqD59ATptTP6ARJIo13ufkpmxpR8U9UJhTdzsYbp/2jQ1dX
pCfwijwWpCzpTaodNWKA5NWTV6VmqUdvgImvaNdOnWQeVk4pZ31pphWh68/EYLkp
iEoMnewHXuMQCRc4WXoC7iume13gigFXGsBVpRCPKNk2aG8/nv7ltKuu9cndRLQL
EMW2ioCVVimGdw/Bn55JxVLRupofyM0+dQtB4oLG4FCenLAYZ1YCpzVg2u9Wr46r
4NJ+m6DCXRLxrhpFDfpBWdtxYg5xViKz0Y9XL2ANcyxHlpFA+ZYOR9UzVAoPsx1T
ROiqglYad08NuCIc7O93HYdMeCPl2ZzsGITAdB/YFZ8TwCwLo+INcTJV2oi9EAz6
Vzv48UfCLIn86KJEF/4F13Jk82Pb4LDifpIpY9BOn0w4qOctzcDotQzqZjmST8SM
TuoyuCRsq7I+MKGrOWTTT0igzlrG/ySTcP0h3xzlMsDEXW3a+rQMVz75N6DUGkxL
cvwZG2pS3U4YoQk+gNxtYTTOU72DeJIhR0xWz9GLCub9GcDv8yylZ0Fg0PpC3d9K
RyylJKm4HS/T9Sz4EclrlVKqOGIdnfPysSKMNTvz1kgTDKrAKg39Vckt9v8SYcE9
oxqxK7gFI/ECpoPkwiaJXEf3664kq4h7WJow1MiGluBOoyXFGeol0NsocjN0uEM2
Q04TAtFcSO8WdgEqneFr6nH5y7CZ6p9tbd4+IiNeFMMR3JhvuEHC7e9OZmRqOd7E
3Ahckp5KqG38+T70mbotZvFCg+fQ5DIeMmGcZBbGABcjPc5GvpGWlLwy2dWiJ2pT
8OI9onMLfWdJWW+zIJCRO5jrHUX11k+8o/w8M/5FgJg2YYFHibed8NN00aUzeJAY
e7DEdUlhq1psSxwFmLN8APyZN1XrLxEyw/ZAZohsdVN3/T08/3fEgkW4zknYit+o
fwdhly4NTem6DsAcAo1lIkEDOTSJolfKXzZnqMhPTwMD+hjrVLm/9+LmZdFuTSP6
l2hk0i1VpRyPTWTA2mw4IVICh+sW539ywjANtsKyQ8OsUNDkkKp0tpnJZxGCcQuh
up+9TWqgn1ECWPFYNZR2LxamQVci2ATOA5/90pAkS9IzrjYrysvTi04IvDnqbadr
6QWUZvCGlG5RpRpI5RT7JqoSeG8c4ZZRpy+HTdEv3VX6nnpHgPHxuxn2ZlE2jRyu
bsK3PyKVeVl2Izd51gEATRxFJnGKZUAIUxV+9+Dev5TnZlPZdY7YMGGhdvj0duac
qN2roAj4YlPY2KIZvvjAAWj1cSKBBCTKul8Jv5xmWStyPmO0qgo34bTmIKDCJ33p
L/9BXGrl2H9SwVLwM5biORYVUGIBe2R2B5IzQOapTgxQQwHvET5HJHBZ8eS1VL4U
9HYa2qc5KvlFYvy7inl+3UxxkYncvKF1iX8uWwyzEVyzVuDXch0o8HZLWsvo2aad
kVtlweLNQFLW6/Goehj7oobLipE4I7TmeOLw7cLex1+XdDynwvz16bjk0zCITdPt
LZ3JjXYXCmjYfDZcSfoPF2YnfpkBN9RRozvYYPkB/zWbn52WGdTfPKrSO9KRnOYN
R4zPGChvdCyqzPmUQJ9iTbqslNdvMo+a7rEGV7oeUMEZ3RC1hbG0JGrI8dXEXA6I
42Gd4YXgtXwEHYfNRX3acqpaqsv3U/vE2iFWk/X7g0K/jhIUO6cMnCWvBWmXqrpe
RZoUn1o/EXfbbdkUlIztl6Oi/EMZ4FamY8gDnc4XquFO3HEIc3HNDbm/bgw2fxWZ
rTNgvijzU7jtw2SYeFX2z0zlWmDWafws2V3jmCDIHiyN2F7EanLGRs7kzuCa1jBb
8fc99OSPGUVgGaFcz5hH+nE/fTu1G6+ftR+Lv2Adm793nAFsK5PCouamAqerpJyg
0ZIXzN7zEzvHkDJN6vVCbh4BnTI+ezuN/OQnsEXepig+t+VXG5RsI2xUr7u+lLvh
POsCI/8hsJP5mgLLog9A2OI6N8eGAQJqCxZG/JhlDPwxKKyclVMjWW9xMNS+WOQb
VrN8p7+pe8ZdN5hLP9UMGf/5ljzQqa43UGBI2Jd0nB7YYBHEA7pmPf/PhcXbkqiU
Ksmmzf5yEPnf/lFMpTGc3HWhUnwOWAbLvcOd/2FZQ+4Tg8ypRoYZ3Qj+7l0Sb+8Q
f4OJ9mmHHYgV0lKRlBl6cwP5zbna1fQx5K9VuI0oF1qKldLamFHBtkgH7K+q+5hk
N+YvejYPGzBtpGMCD/QsAuZXz26lbvQqA0pNPcRfuR1girEHC3+gzpbJ0s9MMM3h
ZZjTGySFan4IUGz8oAjqZw7N1wjQURQMv0ZRyzgUHguXyX1NPiijDxJNu6F5mggO
PACrDJjixB72PqqUcZN1d5P9oVlo82XMcsGRzAvt93/9HEJM9NqASvflPhUtexXO
IlUPnL58jB2plz5VMDnRAWpVhl7WYTioUF6BgV7yY/dUmsIImRd1eSG2bT+TE6OU
aR5Vk1ib3zH28gq0SrkbvREcLLVBoc1oXI7ruNBo707lT0kAasbXmJbQ6+T3WB0w
hwXknJOILgTVucaTrK1kpfB+3ZesPbDVKT/LBD3FLFfEfYBEuZN4+PgvrI3QXVdI
xekrarqdGiyAkYSj32DQ2cGVgFbg5iw+yzJi5m0XPIAb7X0cR/zsg4NNBHHymd60
lE/iRpNsnvM39T81Qye6MTDS4bu3unlgII3nT5eAR+T/Q4wgo8Ej4vYH/gBHQhZo
8Yfxjufo8OMQa544pruUO8HZ2GgBV4qOBAkawH5hqRiIV0H573Tj9mmwG9gPtooG
o1riEsu9Ch1yHWbjop6IvPAqoekgI8i7Iy2NV/WdK1ulK947qqppenuy+nCbwA5X
SM095ZXQaNhe4sCaoY66JRnn7mII7O9a8UwreTM5YWEDg6Nix9TI0akNoWRDTJfR
cIiUqSD0U3HFOMwjeXL5X6/AkOcjVkZ3TABliGpYVS1DF3QHTA4KV/sGn+2Es4ez
FnJxBSWVCPP7TL1BOvHv+p2ruMwHJg1uhMV5cjKUVryUrJEZ+kJUu1PoybUfDHdn
ksc3VTmuTHaaEydRCMaXi4QcA+3lXlmeWqTplKK5h901YFy8+pR0chhtnIOHkhtV
PSJ7z1Zh5hO24x8VpROwre/zssne/8UWHj9h9UBGygGrwOLDhhgUrJmRIx1rREE5
6Uh1ADFU7Jm9o//XVbArnK7l1S+RxqrArgJeZtFEO/2wQD04NerfWRePboaLBLrC
SDgsg2biepwO/g77+8ARmA==
`protect END_PROTECTED
