`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZKBiiDMR6V+CFKOfhh8vUGs6WaOuhIScsvygPnl+/DV45kBI3BEMC8dzENAp/d4H
uUWTQfTfyQIKaUHxHQd3lVyQT4KBVm5RqkbiK17RrdsgAbC97hSgYK4DVL2/J3JK
ydKw8HW1m2dYWrNi6d3x+ZDqTwoOrMp1wB55d7LOyvpZjsFC+SrX7hobt+HjThl7
bHGV+NP4cCwKU3pJTh/K27BLG+tLuhYDBUd7RizZwIu1a9InQEM035iHRC4+Gd0v
MAgKU7rcSmcJl4FiS3zqOeiW15BgKCWaqy3VAaPQ7fPsh6PQz5+e1plAmhl5WQkc
whs7nBLfx49O2FULObA8FhDl0pDSlYr7iC71REhDP/MWd8a9Gkwvxcl+o2lbFRgU
o/6oAkgC1xae8hcwtTdON67DhXmAgxlMhjHt8y3LaYVuOmdmJt6QAz7ctgICQK+X
HNorkwWDpjNEnkHn4X3kzOJspYG1tUYb9bmsYxG5/CyNzMEQYM3OsZ80a1w7tI4h
ogMp6TUnAQ9STgeaDMquV1iz0Q4GS2WRrXeodygpK4tjFiVFiVJ9tho7bloE0kAZ
/z4vk959tOvpbY5+wTCK5D+yvMTJweF2p6JItdujh9faNMyzmnIiME7iz+O4/DDl
lQh7SJj9/dBohnsVJWWOXPipUITlSgmK9MBvXyXUDKsVPHKpHut+sIQf2GxdKej8
FOnTSKpj6n3eVUgzi1eE8IjfznbO8rmcAQz72nze6jUnqE+MUUM0b1Yc8eFkryUA
KHYHjNf0S5F1sqZWi3147vjSPIsQs/On6TCgJaohYNwp4s7wKsyGN9Z6tprPTpkO
wNMo/epipK56wgWc4BflmU+TcvB30T8L5tTFz1yTcP0=
`protect END_PROTECTED
