`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f9tbYr3K+suanvj2FGmbRMdkVXIbOAEYzJowx02QYi+mguxLVLOuffeMb28GnvCN
6f400Yvhwxg8Bm6hpFjFr7WxmTChRh44uATUlXDN60vN3ocYXtu6hR6CwG7KMrA+
x5RN2E15y8WDr0gfIkJkts6KXVZLI6qOGMV+2nvP4715IsCiiLITcIrst/OtgLpn
8UfWrGc5LI7baPYWwAoY0zZZNaPc1ttVfYWF+1tCnfDpI88rpNKZEZxT1VA7WFpD
HbkcqH05roPus61Me83VezG7ZVxAXKxz7elDofASB4v9jqCgXLVodcAslamHTyMK
OSivwGKxvwHWQTUQuQVHZa8Jp31Euy8btbNtoCfun++4VzaCnol/9j0zDB0UMCZ9
70KjYx160Amrkd1YXilINKVAFDq/az91CdAO5MKziUlCI5CVxweULnooI+rAylEE
Z6I9tKuKUjFrM//QMELpiO+vLuz2HwY9XOZrb51WBdfI6zJGbEOefnfL/Dpui7BV
2juqnaE+utLiJOdtnHNvqTwjHbOxLzqdsTvi7LKJIgNgSheZGv+E2Mv0EMKR0q9s
ge4Jr7tkTmh33/BK59KwDMtdqage9hTMXe0QpgaU/xpgGFakmNIsuKhuPBCQsZV3
TasxTWNTN8gDOTRAup3UiogYWvfDcqkmd5dIhR4r2jsw2tSgfVSyAy0ws9lgamnf
/S53E54cDOfIlpBsp7Syj8EVIwBiP//E1eP+32Az1Jzc/5P8gz/MXmntBt4L7+W4
3hmcgKgHhPGQoVx0bGn39qYfTpSMZo/sO/CmnEQ9p2FRvWGlgDv+z2T2IN2SgFPr
LzD2SxQZdp5uFg+qBUcfj7EY9lB5V+GOSVmZdXBfG/od90Unm5va/uHHET+2wet4
lt/+W8JKGTnUKr1mzrwfD+ms5qJOijx+3JbEa8lRvv727/sRHCoMIsGpQuUh4dNg
eilNcnmN+k3RjtT8YkoCL9CHvDTx/GXztkAmrDmT66l8vaHayhJLGdOhWAEUeGJH
4rQx0TQJmPc6Fz/nJjfsPd3gx05lPexym3NqXU1tvToRqj9Uvkklpln61utUSjVa
lsKASpwOPXfcTAi7F0vTr7B4g61h1RR5QMtX2QpYb4643Z/hzudYoYqgDaKFddqU
qiKChZJaGEGFYBcSkU1U5LPwmPlEje9HG3ny3Y8WkZRbWUjXiBps+DvP59lUEEuN
CS6aH+l7SvubVC5ROJP5FwhBPaadbIM8liddf273/aohKoND219Jxsz8AOppSkjQ
Is0CxP8S4lucp+DpzsXfqb3c00YjlwjLRP4vHy3PDwzLzvmYsOVvtTkA46MQBvhx
kTuBTyNl96Y83/kR8WvL91Kbu0PMSnPiNBrmq4si4emHTZVYbbmvH71NOKhuIpdB
urtRzyiUeiaKN/aRtcsZby1tlcDgyH5wBJZWdmLSk26ZoLcT6EWZ+RsToWB2L6rv
zdN0GTkkrUbnkAsTXExE79uMzSnFz+KFL8Vk3BTIrKOf7aYm59Q5yVsXV5DIAPQQ
B3BxTRlFsxMWN1WO035wA7SkFog6gKtbj/b8r8L8oYbRX20NTej9RTLkgl1VonhK
nWYBtT4IJvd0He9UYrk67MYonIO2n7u5o90h+/A9SJgZ0ztf3eTxEKJHGeT8y5qj
+mNHuXju3ZALEQSBNU3wkjZO7ZVH6uOO0Sp1DqCSr1MkkqvqnUEjkt38sywB3RNf
3Cma49i7LVLTB2SdAQ5Y7tNf/ldy6Fqip9hVP759SgdPyu+lNC+rmsIgI50ggaxo
Tl+qucJxPYOSZqiJLa39IJEVL71OmHYQGb3FVY0MW3dTJmAIqWk0yy27d0BOT8mZ
qNjpEH3DNeCH+cmfUphQRYm6kY1VpPnDvCk1EPNZKWQdQb4Db38g8kwIkqNuhvc6
QLUuKm0kWm9myh1O+tyecTNVpEHtD9dhjKNw5Z6LUJrWTJI2S2p1C+QiZIaz1R5B
N8jcIvnxa5lJJCabwV/bCImkG42hkezRyu5qMbWyQJYoO5sd1YF9QIGdbUb/Je6q
KlsLawASrwLXQtj6Y/9slFCRcNRuNXGq0e4E1tptm3NEK3SWsAnvC6/uB0wtDWmB
cMBvkelRbravQxcgqUvJ7Fe8x7A5bcsg7L1V8g4qlwMPQcqBcGLEKMvtMUZlcNAK
0TPtMk1/oWTvaS1XSS/ntA0HOIWKSLt91cSjrkKtHZTVnW728p+C1/4RQ2MqwCu9
rnv8JSsZPj0CL6dt3tPtoTQEqAgvu4A3i2Uy3fJOMAcOXwiGarnSYujNhiCv0v3k
DRan1Yx6eC+iqnE2m0d+1Whm3tONn3ddSDuqb/n+do+wZOUQ77tyRT7AQlQUsy1D
+VVQ90kEyrzaRs+aIHjCr8bU5tnsDQI664CEyXirm1IMVSaQdHH94/fliqBRXr+e
eeJWH1G3ZT65NA92ph0MWZn60QQNMTAtLLA45zqmdCtAYsRzyO753uD9tk2HKA/g
wlXr4KGbXuC3TXtEsT/3NwKEWgUauOOyyqoYoCrf74kKUwzE3wTyH7N/QTK7XNhQ
wwB5hYLc4cvVvmovhrWJxZ+m5VPxI4N5yr/acqkQMZMO3iQ4SN8uyR8frrQQmkQp
Y+g+w4m920Vk9EozKo0uBrUH/Y3meR7NPprn1ZTH3aJT8bheD4a8UrCRmhErft4v
k/Um6rOewiYxTrB2M+p4uxUR/XJtpnKwrBKzZHKPAjV1KaYJSuaY7wxZUTxWsJK7
wU+eJ2wSpP5prs86mE7OQiZHe6iEoOJyBzcZqnzA3pfKwhWk+nGfFpBnFz4M7byk
KXWsh0PfVLKSbCIicK2GV/tvyMn/iPXIWCOiIOmqXgDIafV9Ho7QsOpqdQMAfnI+
qtStZYkssldCdIWKjD/37Puqk+qToQdx3q3lh0PtvuuogbdgFlNQTOEfmWCPHkZN
5KH9F48UvEGgWiD58oiC9nvuEJAC0OupBYJlxkNgqDI4avp8RHsPXS14roIG8ds9
0W1ENI+SNxbDIp8FRUNHteUgXoEIlnxkglNDR2QL3WKZUGFR1qag9xFvbbE+Dvq8
IhKsS5cCY0XERdsLsK4VACe5zaASBt8civ9V5h7cUdY+YPwWSkbZR+N93YvCgTK9
Z2dj3UrYUZ+ieekIqLQWtLsX0mARCc7REATqceJdU7ZC5rfmuYXUTeNAUU/mC4/x
yKn+U/Puck8z3XKsCvdOuYE6hu5E8ZbcUa1rKOSNe7L1Z+ky1Ao8Iza6mqUTda1k
woIbcZveEvK505SDmwPziSv2rpSjZ8SrqwPljXxHhAbMz0L1jW1+MqCZnPQJO5er
6n4Kxr8X1hQq7a8DC6NVsFeS1lY/Ox96qRloIFExj1c+RBsOQvbVkna5JDSLFaUP
huk5ZGD2K3Z6nWdbYSS0j/iXf/kxSN/TwZHDi+SuH/JRS+TeOHO3TgCvcb4hYCZc
AOizzdNuk9I1uEmt5ZQY3UApiRCMS3RfQUZ7pguz6e2HRuLHdgz6k5lXNjrRWNp9
I7bve49qES2hTCA4aXrc4Xha+eUW/1b+p7oTmi4EEAGz0RPPoOnk0bZw/gkJBs1s
GzxUE0krR6+4ZKVvQXPFzPX/WfOtSb8eE692qoN+pWGy2qZ/kpJBY3zjHbA4vxc0
FpV90hVoC92JTwIECZxxD9RAj4VNQJely5a4DVmucymSbFnWjmzb1dbxBCzubaKn
xw1JVJbadojBIcPBJHh7CjiLh8dJOykX9EfrpRSwhiJGic22Z0C8wi41sO5T+nmw
MQwoX70hz4uf85SqZzpAu/DLI5gpqV+5EfwYfkDuFqg+Jh8y5wCP9rCM5Ves0NXX
tDyu2lr1bWq/l+CQ3bDHW/Na89A7mjgWP+hbICb0E/m120wxZ0iLwz4hCKENyC8p
m0KC2IY3F3+T/dctsV/Co3X/mrnB6OF4uJ6BMqIsPuGSnykaxvuGYTjY3gAAEGKz
U3jDyI4Erqwv9/zbd664FiBND4PEHjKraqwxal3K/GEqopdw2GZodcvffOJ5mDXu
mzRPiwJ29aGaFTghSQr8cU+rdtfKcC6DbpMFbfMglhUWFGg907hGuA1PJwBseCde
dC2mPUxewW45l924TF9OzmF4MC42bm/wzCQuDVGcDMhgNi1WMUuWNFtqWwHCFOV9
uqO0IMPLDEiy+E9OkLfmhAlUFf8duyB8GzbvjLKjs0PhhqCWvfnebuW8cZ69tPn/
TpT+RjYkdpJ1yyNjxqG6TPiZTvZOrW0kacvFUMsmPKUqlKnSvlCD/iwGpLvcuFDO
4VzVcezaGHgORqQAAqv+Pj1XBwEYV/X+Dd7+jwYGyQytJFJ0FcgU2GNlCrzGi/AR
6+v7lgMkUoMKB4YOBTdeN37D/1sVvHQQcsz2iX8a5vG8ZNz3ub2Tt02PLWdiqcKF
SeDwgFQfz7ge0PmEv5D2PUkB+zzLP5RtOgHVcI4c8pXoWKwvoDfJqjMWeqkS14eZ
C5sqDqZh3DCqiFXFY+NpuibM0WEygnaAWI08NrmAvq6tgrpnRVj897/6X7rI8XHj
a6wHR3x/+7SmacKGPVSaJTuiORdYa+Tesi/Xrv0cmrqmsS7fL1DL9oy0rThkndmD
FVgqwbFkwSXFe7t3/mAVE8mKNH+AazX48hq4AbEpeDKVRmg8I99Mw/5OKgZUeTSN
vIgg+Hzx28tu3+tpwI8v7/S4yia76JWYGH7iVscazRiZ8volzrsNftw8p8KGX+HF
1pJ16OAtgT42r/7H2TDwBLzjk1fwaED+i3PBL7AhCb6hmM4PS6S8cq5MdfrcWtkG
r/zxNlic5Mr1gg8U2Y6fxL5mjqtzBx0GIn0ZSci/dXz7yqXIqsJspEB5mMZqvqTP
+N5TjzmMALTz0kU9TNtcGI8vDEw3fkHXWCLD3GZgWXiT9BW+CbRNNSfPGQ4sovWV
6ywX8TAb80GeoWOqsYs2400tjk3rG8SkSQoIDzrxUA3hNWGt9uw2dmhTIYPQEBbS
c/9yutuKG96qLLfMs3uxMrLlLW4zaLH4tHPnBFVeVGxaplJLAM0QI2OpRE90j/al
ZGAL/Jv4u710WM8qF+npC2aS4VqImD3qJsevYEibaNyofIo9OvoIOXOiAAAxR9OG
fy/dhd2HWE3SKiQT+FnQhMUz+npuLp93BnhXyiJPr8TEQlG4Xh/hlUa0a+i8rFlI
V7x464ZS4jpdql1SrUubifULRkRkxcWmQ9nJC4hUdQmtEcTbsa7wn5JXJff5qXDL
I3a7eGhNylWuECvJOe4YemK51i2R8dcguhMFIMq2S9jCrVsRxGsi/12nUnnwyB5R
Ep2AvVf99Xjtrtk0uPmTX8Ph+6WTdzZ10IMdFxhLPG0AwwobPcB4Ouc8w5RSoMeV
/oa4PMiNFj2CbrcYOzIpPpmCK5YQS8qcBy1YF6LNRQGqY5iz0SAqAZPAHBg7xZsg
jmdz1xTZ3WlrqSGfWu4Lf98eT48vAId0K+Kz/WtvTNXAwQniUhQ2p9n5dKozy+OV
JPN4dk/X/NK/7Mu0xciFEQ==
`protect END_PROTECTED
