`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OeJTWR0ofu5bLDb+piRhOyIWIwygKu7RS+Aw5YksFJYGVwbvTc/apGViiAyc1EfI
1sO0kDgR42ZuUsUebwNyuZKUkSezPKord6Vq3OQhD7+4dhWOdI67hPj7h66kUPzn
9f4aTgWMmJ8qojmEhbKEZE1Z3L/gQnbR1b0omybZxLfhyzeqhmvVesCsWam6C2LB
CorzUk4ne35IYGo/n+eBKWoa+OJLMxCABmTP+YQqjYUjT/Bn5Dr2gDmu6fSuFWVJ
9qf6Ek8reoI7q32sfOxHu6jJEx5sN6iK2cTRlKXvInfDl+315LegEnbCbLZC0qiC
Dl1HuCe0MzylHKrqAniDDh/z7kWghICsikljOxf0FEW+4YlLvcmCGVKR1sVIOCr4
nQTpSXcE2AemCrwIQ4IO/ZxJ2ZSMKTEHmnPVK1IskWH8epe8OsD2+OTlYNpetSmU
fmoJS0EC5pfTqz8u79m/aNcaEWCFHZUzpwudYWv5vbP2L4LhEyfbgwughYJOOBV7
SgoZxizz5gkN1vbBJZBWE9YZ2Fw1WC//EsPoGqx0qYS9EX+HZe+gTlCZY/WItc4V
Kr1Y+z2uX0MvsCnDkwLx9aWNGkOnKms9sMqXVzzbz3N+CxT3UKCGgBWtRTDBGF9P
YQmmhxmKFDZm/NaWP3CGceD5LZitAO796EylNoMQUDoJRx0uWBFSGu3pOApVYv7w
O5sFBgzZHyAdRrFZBUm71pM1C0Cqsqofi45kmBD3x+hpGr8Y29mjMlGyDNIPhJ5V
j2lKQfwfS6o4RyfBbsa27ozi1N23iWEA9sBIyxet7spRqVbmgDn7Ah15/8vMBKIn
E6ICWr9yQAPMn4i6tOvdDQZwWl21kPpmUpJa4/EtTH8n3O8YkQqEq8ryvVrvjHCU
TYaqw9/y3lTXnbUfrNWp2pYcmCJGA17cXJ9hcCMi5FhZYsBO1C/C4wiCv0Zi4Nck
FxDWH62v9pGPP34cg8f7yHmUDZQ+UPV/4B/TOtTIQiXqAEQxMNHURfvH8WMeXyt8
km6V7FF+etvInm1O4JPkzlgROBqr3pgRzHvlJlfmr1w=
`protect END_PROTECTED
