`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HbzwKdlBmw0dqWX25UTgEoMyuJLbi1bNj5pWHl8hTUaAIBPVzAz4nqAtluVRecx/
zPmrTvXycScMKwHdFv6H+rBmKcCYqYXyUJNVHLMKWx6EZwd7Rj1AVJvmKDArHlHW
SNUGrlyZYkO15RehGLoiOkeWkUW4MEAtf+QBFbZ6jzkkddOvHxuSy+yq/8JdcDkh
/87eYyQrIuBsmMizjGvpE40qPFCso0mLvBYSt35M3bOTw4dYIN7P83ml2Svv8jdV
mleEjmTMgMAqJ06F/Zr/2KYE+TihR0BGjhQhKfLIOX1YXdREtQ/E57zN5sqZ8Zpw
lMBgcqP3ktOJqnh9aWn/ukqi92WibJr6c5OhPNblAPgGbd4kTZm2DxmqcaMdkSOd
KhmCclHYeNyvW3lhWxWOYNWi3w8xg7oWD2gN5ZQGVhCmw4ebIuyjMwjM+EkINzLq
e8lo9Yc/RJ3DvQ+Jpk3YoOCTx8opWjO7ty1qRGxqKqN8yGlQvEgaQJTFnDjzTc2W
j8ks9t7Vpgi0xGSDOBHOkvxaO/pjkBbJlR+APIc0r9r3STx9P4P0jqVfZPabzt1/
1QTJFNW/2s0nYl86wZxxB4Ka4htpIcbT/T028e6r1djtW/1Ps+0iwFKzwLtFkRip
9nrYJdTzB7AKFmqg42YkdHiuVNIZRMXw4oBVqsq0fN6UthLWI2g9ZOpLODjqu3tX
xqAzFtFDnXyK7/37j3zIsFoCurQJg1w0sPjtzHgRwkUiqUthfR6TY9bfFzne+bmO
TiYZJrNwrw27eobJAdpxN6WpQeiaG9kRX2F7u56Oarl4ACrZ7q44yf/kCiX3DaS0
xV1etSJofYSd6I7GaNHhQW+QfFVU8oG+tTGNoFhX4s8GKu6h62ujN749lVi+Ouda
jNj4tHq99z9kkOqN4NLfS5AwajR6aH7sRqWSN3R+CRHtSlRrh2o2CwWceQ1U1b69
NTvbjIyJLq04yCsS5tK3GJIJnJh2VtP1RJ7ViweCdjar/h6UJT7u/IJ7I925jRi6
5nnobNreUkIMlgMH9N/tAGT8Wn3uoX7+BXNfQDU+36IqfG/YOHWIgnK29U4WTNz0
pByBvXAUdER2tbhNd1vNI++Bj1wSt5P4EHfwdC6V6pklHwlKhhxO8WiKhbmXnK0b
Q8CBZtxp64Df26qvo/ztTE1bCMeCxPTkWIztrxJDKsPzOhrwddD+umwQXRaOJ1/m
LPlV3mVlWmVquNwnys1S6UY4H6Gt/12UfES+PDOjOYBZhe552kzTLgRoW3sZ12K/
1LE60QD3vQjZZuuiTAtDpQPyMkjifzcJgtC07w4c/PZtghkzMBHINKzuO6a3dxvO
B6IylDAprPX9/WpjARQh1OP2u+ZpFQO2QnGJT+ry1uc+1NhNOajuYFKU1Vh2kV31
7QhUwU4KLDUjV4V5SowuhviBXH9f9vQREIOaNnfo9DPhmbEW4VFE+A8fnIFjiLiy
l5DVKyO/nma/8FUakgg0lwow++coJL2QVLB5hdl/jcTrZEuDKL2jDEEShL+oIkNQ
w7l99zugeEk2CyKe5yGm8j3n0xsfWIR4ElbnDUyBnP+D1maPNX7yOXsblKYJ6dUr
p312TbcgwSzklKs3MWChVwBtYZyUImieVqUlK5t3gv5MRni4N+rimXUwj4WsP9xL
pAb0HEDXDS3e8nth9L5MpPG/x1KFvhBqkxLgAH41YvvdOxjXVzllT0QBX6CmJf9Y
ekDk1zWydgf2O5XqosmLr9QBkwWkta2LVhCLNpoajKaZUFMLx4puBreXNTcfamzD
fiUBUDHcKVUSn0HTJDJBWLhDt3YKIZi/QRSzhEY+f9VwcjiJy4G9OiwfWV2ELER+
xvadHADOx3gpwVeC191Ye08y1juSRAbcvdbUHiFu5algZBZ4e2UhnbcK3GHQhHhn
8+W5jOHEHXzK+3cKmsMqYnhcSON1Gssi2RG/jT2W1Z32jR8FC4MHRjVt8+jSn0wg
FuMRyqQu+dDj6KMdE/SwX3lkTzYlPzwEhLKzDFLGHuc4QA2Fh11G13Jsfs9sso0u
sD840i8iUSDAU8PSR/uSliBWXajCWmBDZ9fDg1XA1Hpn+SsLsce4snDWpjX9EN89
2h6z8xP8nyoMxAGMdbd+4dOmwO/5ZQXijXrZx0svSaImKdXsS/+CwOPKsZXbH2ef
Xo3Kl/NtT0FrENR4/A2ZfqwcYtPbZUed8QEZ6MS+q+nHtJxX0JxUD1BdnbO9MjKl
M8/XQwO8s1NYXVCFA8f8bAcdEcnbj8xAoo0voYLSLqKMawo/F2CChP056c7dlUXL
4GfgMQVThBTJBQrz2daIp4FETQrWTzKa16oEUpL/xCXb6UmQ9PQv61R5xOhlh5bU
uPse9QkE9x+uvlBfnErq3yi2ApdFIJClzQctTR4Q1cGXV4mPJPHR4KbER6wC42AV
182GR0vDEQWtMTDcbT8D0aEa64jMLbptGHZpL4jCvdPLizJqYNe42baG00Bq2O53
6wWWO3YSYgRuEccu+49lZouDx1b2x7E2EIoCj6mcS2KNDMw/Rrzdai8DCW5EZuHN
nAluDhxIMtCGyrwE9Vn3U3m9q9WpIiBCOF9ZdLTXDmVTpGpJfaqsdQO8fDLgLVon
LiFdIz2P5HzS3t90Iv361ERN3vjnfZR+4gUhnYkjAQMhPCiW9WxFa0apKFR/SiPu
nfI7+eJvJ5U2toEuLqpNLDwUo7mfiSRYP4aLQpCbtV/ju6JqBy2ElPzWfpeOqimW
pSFiBbQuLUXfE5IlI+AB3Ym1JfvOUd4iEel13mRaiq739yuWmfvScdhLmyW7WTxo
tWOKywwgHkwN29YqE9rVlqcjRSzflFhS7YBugtKDtbaxjq/zJ8kbHJ3jWjLfJHcc
cAGNGq+p8lcZxOXtneJHUxiopFcwKRK1ttCPjWwyrKtUBczmT6Z6VFURzxZLxkJS
zqD5dGkou9Ghhwx76JenkkFdSiAJw9xVVYMmPja9cDA2J+nvMy86sMpDsjoGHWJA
YDJsNkXSGeExnZIHsBooYbXB5hF9oy2Y355JdjkwPwTzkC9pzOD72VHPBiDZALMZ
hP8T7ypBsmRWHzsLhiKz7pMboRYo9Q4IhSGcG/IMUYw6w7dBP7yZAxTDWohrXzV9
pq8BZx9b1IU+le6GSTBf+huVykQlP4v9GZ5ZuAHSSaYzgd2/npqZVLHp1SKNFmPK
A1Lcvr4s9/XRIAFKPwzsq8Trfj4NXGNymBUxtSlgHYBDuaGXz8XJNvl/usoOzXlr
WLBnS/xvFJXT9FkwRSAm5xjAHNeLvKbaF8rVm9sMtlx7RC1U3jx2Z90l7Dqt5nVa
yizb9J4UiiWGzgS9tHqTjyHZpouOFD3Cjz/ZnOLG6zDmCeVqHQ+j7wcQzYvCjYDs
+QqdyxTgOoNQs6E3FclMIgo94WQpXFklmKBwOK/MftfwF8BgaBMcZ0Cty4tPYEZB
yJK38aQjSjy+jCrusUmCTatwrl7pMvJ80vuLyzYf7KTHHKyKGfR0OtD9G8jYzIWe
Lxdz3EccrqUhY5CwPFZrBAdzPqfZMU0uPxYdFDIfKqafOn8umjbf9TVFCZlRe9f5
xepL/4Geiy5mNCV76cPEq1p/gDNv9v2s/spybnqZ4iF5orCdowqWclZV25btaubi
oHD3OqNtZFJGP7IAZn+BIT1jdA2W8/PzoQLDNLgWmr0KPGVau96uAwtWESkOwmmw
6pnYpvPYkJ96QYPwBIBhYJ+dcxr91NNY8w7AGdyINKzCGbloPGTy3J+lQt9Ux04i
DDBsBsZtxFFZ86GDw8MQ04OdvkEhL0xXStmNaUsuWNx2028YuyCPtO1NAINLmzUJ
55Jpyb1vaSWr+z9ziQdrGmiwAvhlGR/UY16+GzayjrSZFu3wz51jqtSJguLN41tO
PBIp0XdWLz260i0MA4KGW5pEuRaJQnftUmCtUfLncvtTBhbmu59cd+YinXV1RBE0
+Tl+O7q8VarBfEvWdjRYK2QderccjbteS/l+4LIdXZOMWHKLyYRKG2V7tvoM3Vr2
fHNE09Bz3q3twguky+4aSSZffo3drh+s8eaZt7BZMy8rglEq+yTpI/7hmp+WwGw5
2vzF5FW0oEeQ9nTp1htmu6g9VTfkCw7INCD7Fb89OHg7u9toeTzBRF0L2os6xJJe
Fz8ZQhNQifOzC83v6VL8QoCJBRTjWGGFCY19qJKcpnvPyhHMKjByqGBEACAMxPxk
1dwZCufBylRKh1wxmM8pW7Kyq+UzO3bIyzGV6v89JpT6Rbo0tGNcowutFv0xePsW
Aozm9/PXFGzNnxCg8MjEV/lQiYmzjrWRhoPSkFj83JyJtWH1iZ2+e1P/1Jtsoyik
16pZQnlM1KSnPW3Ulyjjkz/jNHzdm9nvWqHEbQsAtDx3J2/AZ6UAq/l4PuVcAfm7
PStWQnySj4A8aRthFrN5NWAwXB9aIbax1rEsVNqN+YH+cPq3Gy3aC1ppV9GN4W/Q
aT0SE9HBcIZ4D72AQbHIs1Z5pP0yf++g5h0BKzcJMTi5KWw9e20ZgRpp/LW9jlp1
4SWFrCAmHeBuM9bS1XJohjGl8K8IkihBTELhd8NWvNypUxjcZLV5oi4rqcRkaaCC
xdpbRnYihU+6vDLuwG555NdIqDGVVzaIaZXzjc2rikdZnZvzY2sFBDUNGC8LwVKn
dqPnaGAdJdUWNdeHDpF6XWOZibpWxaBSD0waV7WYWrkZOuHMjP9xpfMGlBzWyvqR
DMfuzFQGEncqWEDkR4Iri9H7wm6sCirk7/Iy+29Vzi2hQq+gofnA3f9uTSSASlr2
OSnaR5pIcAESYo/v3aoBM5er3vY9ovnNqQX0/byp70rjoIRkjDpfJNYAn89oAMy7
sE7CIEJ+djTejG7xntGI1vSTUbX2/L61I71D3T52USRhOoAa4alTsKhYR9+ZoThd
k3a8R5VY0J3teFURncnbY/O5Q1kgPtygHk5n+wlslMlD/3oz47BWH4+xt7TDnxHK
PQMt9KiLVv+ARh9sa1G0beWgcYtClxKogtsAIz7v7DrZpvbjmsm80JIEgCOvcWjq
HgsbvC0Gpvf/YWmDobUa9TKsm3nm+1MAI68ZIYfVkHdTygly5BlbzSU3GrXzlmh/
XaiDZowxsi1K2RgkIxmhH8EUlQFXKD9ejuBIuI6pVwi0KiZmTjd8vdzQ5G6HuQle
3uHIvnLK3cswFSAWY5bsYpr0Tikw8TLIuP/ASAtgAh/SzmjarXmWYK4fZnsKioCu
P9WJUO7PCHKM9W9HPlMt7NvqArKVlVO/ULFtLM+BR10UyhIXmtnUFQ6HDN7UdKKu
6qMTO1v7lcFaPcWuNNYXTySec+0sXAdDqgiQyemaWBqw/rn65f7UiW3/11MByPto
pt4G376Mjl+7EAefs11GpkWjrFk3ktED94ETkQdlWAEg9y+CR+7F5BESXquw6nZu
vMTOnzHr7M2ynpzFZAxFoLm0eVW3kBJIdAbIba/QE4ySSbaan3vIYWcN1jo6/h4C
D3fCAQPD/wM4LffaL42IScP3+wt70Behi8/OILMYKUd0d5lB0UPky3noYujmEUl1
PV8KP5XGYfISs5tZ9n4cmGnQOpkpZ+MIirbdYLV3f65Hzqb0kwamp9I8gwUe+awy
JyqAgT27pOCoUzQq29lZljKCNbu2QV7ME9W4W+calCAfZJTetVpAASgckBZYYvYj
1xtbSHkpqcTTLTFxy70jQXId5T2kcy5OvEaQ4RuyvL7jeFFVBfvlqOZsxKxinjoo
2Tpg3sj1KVqwlwzUApBveLwC4BG0yGYy/lG96EdsZzpl3wPf/3+Pn/W2VIw1t75d
w9Bzq6FH2IIB13mF/Xw7/y0xnaMqeZzXQoQQz4jc1spNF4yCof/3aUvFvax9/Bqp
MGbKwQcfbhX0ix7FQT5bnchdU5zgEzgh1A4K0E6IoePYsK3i+Iw6CsTR8RhlwnMk
U1K0E4FX/dJaBJUOWvGTUGNl9wYc7Xb8SyfFvv3S7JnnQMJkAa+xCN31HC1vIiRY
55qQVlYDhcDi6HJqMOwWtEdpfKQRGxt3MJE4dpTba2/qnRTL3o4ZSKPvFHbkuyXa
pcBp2VdM6CFb4tB0c6tgn0LIWDs1+sM1Oh7k3GrmvghN3Mn61+ChuWKCoxxdiqev
jfAyiE9Ve2V9HlaUc64gyknrMMzoBn/1I/IigCV/fQ1FERZIsdOLgd/nHKoXecqe
FRu/UtxUk3Z+u5YFqLO0HOEzsw4S1Nk4wPX5mQrfBiHHSpUaC437KzsdnkVbClE6
2bmXQL5D0QImFZGr1RZBHCePJYCbO6EGLNHkCgHZaHB+WqxsSXqd4hsdaqKXckY8
gkzIXX3qKJuXcYjBRPN5Hn100UXuqEChVAvzeJLD+D4VY5fw0G6PwQcS/HrrfFgX
Ze3KmlKUJbh+LC664gsbIKN8pg9jjAxJhl/QNvBUKOcgkXjJolHeVyu+4MlnRkfl
+4t67zqG9q7/6z2muyTd/eAaCqzVr59+Cz/lNPLVodA2GcXEg3HXksEFKolbPcEr
rU0gSPabqyF5ViQVVMW+C6UdTDCk8HhcdFjj4haI3KOryH4T37HiI9+/01izPXMm
rLH4MUqs4vcJ/SfJj5i5XZcjGUJzupiMc/tNQMVi6jpPqu24cjnio7dfHJceTz6E
OCMYHEZvSYcircDsHxYEu5VVn2uHW88IqsuiiOjJR1D7lwwidKsBmMqp0BdjxaX8
bI1a+Oxj3M3tO9Bhqs4cptuiarxf1xQHNpwccU9ZbR+eR8+oxmC6cJMXA9TBXEjg
kXdCYganldjtGbgXrv4Ab0/RYt3+cCyQO+nIN/GV6GwhBv0OuoC8wopwzCFh0DLg
J4cUCXbix70ylReYSyI/gdLbSmYyPxxWff1HUjWZuzuQjz7v8nXfmdlOLiNcDiN4
jSIdDWGpINIrCD74ZYQLGOqT76hM84ggQzVhoN+XS04O434rbzFtKioJO6ctLIOU
/kgH0aQbCJ+vKkpe/KSLSy+/Hi4LtRCeNfgeVF0SK+bYMlIhCeg7N3+j+ibHwX74
CUUPj8lRgQgn+yqrqtZ5AHBEIfKX94mxdiNfGulTpNN+Jy1ySp1/yn+tnsdoHXRN
CLhUAzTQkcKvClDt/ILE+mTyuLOteAdPVExcfLGh/TX4Zh8UiDAHWbp+sWZ0Csde
gECKSVyt9wlT5ExBs6PDDAbvV19MEhi6QF3KlDSRumIP0Z6dxsFzMnl11oWJX57M
eLOAgi394yHvhoqeJFNuXQZERb/Tc03PvIjx7x8i3TGbkRrGAp7zftx8x1Fr3+Kr
FJqmoa67JJXgnwdKU7/JkeqpgA8J3hPThxI/ddKAdeMy90wo9WsOFLOV1jmZH/bu
znmKZ6v6g1DAJeoDwLRvuqJz2aW6ss83k7DUipgD33VAykn+lel/DSRiE6f6E/iZ
AjXbkFVJDVa9QAPEY4bcOcrOSbONolZGG3UNEw2H7wfJZmUnB6qHp7unitVSA61l
KYpgRhjX8huxKhfdD5GMZub1vyB2RWSzGK2Dw+GPPmU7r4VWG+pHDzo2hOwkxokY
A/IZG4Cew6c0P84LGfuh1zdkyNNfkkUi3NXwq31V2zRKgQSzsh9DEDOfaxCkaqBJ
RU2E6TBNAoP2wVG00v+x4VaFsUidytkacAmhE+q7J3HoAIuWVnOTSEkAOP698ZYI
5EjkhX25JrO6tWEseJrtsvOjTSYt75e8VuIgyES4GW7G2ve39uPblQg4NNEQCjzU
XjDCkILhRp8a7WxLKQTZ0S9x0AsBZ9We/xCI3QPM4CuIpnNYii4RCjqYPTEeO4sI
DcYlzfd+zaVoocMdth+QodOo6Vfn+dbiSj4HviFrc1kUJjTr3BAJN/nko6SM62TT
s945L89GhySfZHaYRV0xSSVIJv087j+muZ6M5syGkl+9LHAvA2JxjnJBnhPCWpcp
SezLffH4EfFh8dw9UcHyAHV5uhs1vFJjHcimoneLx24c5quJ2DdNNlPNr1vkhiBQ
PcX+s5dyy8OA0H8vyqnq3nyTw3I5YO0pwlyn8WtIS9BYQtWncFkEebg7mnqfDdxk
FaVUOA6nMfXP1NLmURGk5fyvmj9IczMnOC+3tEHH8lPQElMqiLNBlhyqoNm4m+Hh
njb9KnPwmrEKbPIrX4Sn5H3/DSBqljRgzFCfqGlhl1fCkc1zCkwQgmGOfeV5zU4h
8LqgUq2tGTcb3AeOMwGnz5bzSA8vOz6GWyoMcpdmdZEOIDBew+qMufbyA7MwtvDg
cLIh6NCr43qBEwhkpJrBhnHWb2OMpPrL/RU2Shuy4arnMygam+zmeTePufyU0JyQ
2Ad/UoFBcwIzsCg1xAGl57kHcofBl53j+A+2WUr7ETF59Sn/dn5h5fyNcVvT0vhC
xsg/tQYvu9u5Uj9psgnrbYUQJouOX8I8ljF6DDko+c7FsY7siCkpGdaci3S7F3+F
ki/52UX90Rl+DPyAhJYgtiebijEPECiW1XwV6S9K/Zb+a0FPIYrlfGIgAO9X/uaA
tTeV8KxvEXhaVc6qhNUoxN2Ky3BzrspglOvWjhjTia62D6vLc03tx9msgvucudsU
3XfYpHocqyJczeXAU1PITFON32+a4P21G0UFkm8iC1SE4RX7fRG/1+QY4xySh/Tw
OkIqxeJC7ttUklqO19r/owjX2Usz4RDJpPR+KDBl7CuTZ/nrpwAKQ3nBdt/kWS/m
Du/mIg0Fq8uJETPAjqWyfMQolTMCSRNZKTofVez/Bk9Q+FwtHQ1ZWfwElAYZxlbS
8MqaPoxCamo/x5GMy14NalA+aFMw3L8l82EaXgTDQB28zESaGcLctL76BAbJ9uXy
OwDQDvqq3dPfBd9QO41TW5IliYaujyLnC64rUjKrN+SzeNHDlu/mM/W7E56vI4Qo
MgJpYbPVE6dCGE76C2V2CN83Sn09srn7PilWovaVyFmAFVx2RN/kK3JPGUYuobOC
6zlWoemWQdLIJ3V9E53CHAqtOXR5pmT01i3cvB71qEeeCRfiymggT9+GvJjbZ0sI
30UQd/Uytp66ZAZwJGBTsfyvlXkpkqIbiEglnMeXjhLrDLzpLZgaIYApu44vSqQ6
cnLtiwQnbVug/8DVWXH9YXgk4ywjBTdvWCK1ucFn94pFQ0hZ5uXt7eJYTPXpqz9O
r0ZWoQfbKB10xZ6ijfV9yq9+xi115byJWh4+4B5S/TmciMiHReKdhgVMHtiPXJPL
9ZYcjIaR/sf8rRGFsO5HGbvAeDtejTIeARnN3wRSWwXKl+qS3D/xfYfyHv2rP8Xe
Yh7XRTzbCd/I0TcS2qBfcw0NkqVOYcbkr37t52tWfJHi5SRlhokqgQ3jXRG2eCvY
8qUXcivwiJOeB37OyG3QXM9ssy4lfJMbx5I6+5aXZnUBZuK0rqJCfi/L505d9qhj
W5ltWHD/K+GPrhubRS0AuC5LqtnWiNLg9Uibtzv2rvuFO9vpNTFTkXZU7skoz6aE
Aqv4jBmUmtB0ZbFDO60M4W5TuH0hXBHzS5SqVmj5kILU83Ge395lDlMhg5hFM3j4
GFeD3ThyylOJmTVf9OZTag9xkVLFp375MZ87wv7PieX7nmKH+d9F3eFbBfdwRlQI
8S7Az5CljQ8bn1/gZQBsQ9kDf4UcEUkKk7G4mN+cae7pZqZ7IYVVtyHig4O1dOYE
HJrb9jE7gYsM0IagqEQ9e2mehviEVegIhQ6IDAAcjCp99kP9v5+I7DfLWDLYKDn2
Z0ZCg75B4H9X/ZyyTTDcaYDUBG9sHNonmrFLNer0gx7MbA0tyHlrCMLwUengW3/r
XzXU7p69k/Ctxtqf+C2GbnPLp9w+98o7te7cSImzx+wuCnjtvBM4pPILzodJlWh+
dyWly6M9dtkxSdvDxgR9dQ8V9vq98msBHK/gQlBb0LILfSXn9dJhhYMLcUgIRpCh
lteCuIn8ShlxCS/oXcEC9JfW9tN5QZF8FRizuNshAZLoH7rTxPF1chkNYYvHxDXA
tDz+cSEz6rIxU3wJN9uMfJ/UwTN6QKNOOxc5MQb9W3dfWMlFw62BRUa9Cd3ZCIyL
fXjH9r7HTCANYnD5EuBaOCj1QkpEDwTGaztnWecKOcaydaQPRbHpPZDDWDxjBM/2
AxFW2dsGESo7tW2XVI1HjJIlKsaPlU2Y71e+GusP9jM9Boh6Vf3UgIlH8LsCHF/k
2dJ8fO9e9nBDN0crGvcLA8WZaslhCPFThFepivw+s9dkdswnLN2Ubzosud+0mTtI
Y8FRpH3Cia2IpZgMdEQABWGpvAK0jc61BXxi2dgxdmYmoRSiUf/TLPc/oefLhc7Z
UNivk4aOdk4ay5tMQQjNos/dQAxK4D240OkKHe62zaDOnCeHciCgWNMh9G+fpeB/
m7Et8jb25GGi1eeogrSAyS/mzO+rzu7hni5raTO/RwIzCY6wPCqHAVr0b2vKsYrN
tGD5Rv3mK5t388cWDePB3ZrVthFB8ZeVl/qMRNjbVK8noYeC/QjNkPahYQy4TsBf
0EZo6Mi9J8Ycvte1c3Ie+pW5GqdLaNrRkl/muzFZuTq1fy7lev/SbZcU7ikwJGSn
Cc0UuwwcTTPhsEDGU7L6uJ6+5co+JZvfAftCuMFvmA1OjFLxv7UGlPlzUaTLETbj
3lYUn4QVGJm4quHDQZal/Gmd7Jm9gu580xcWjcKRXFl0uRijQoPSE/C+kAiTVPfP
/0oIbutGIyXo0NRVo08PbHETGqjoWMW6Q3M2sltQvYIfGaMt1HAXeTw2Gz84ipHF
XBy9y4q+vOZ1apqFSWgslfMYIa17ybvszHnCpavdshbkyBdMtLebZb5lyEWEVI7W
p0i4dgKUPkWVAsLMiiVnPp6yVBUQZWMHAAeSLhh3YP5xMQS/UUyBgRMPV4WRas8x
HdV3SSoswweAdl/Px4/M39mm9+JZoEm6sOdzUvld5ZbMbYEPvEiukucd2TcLMTA7
b1ri+e4mRu04RIMPA/WTWtheZJ9x4fgQV9tOzCV2P2BjKM32FGhJJI6ZmPt3C0uh
1Fjoqidulcn8lCUPFxU+Q3RU7gSrghVksgtQLuhgzAoGmB26n7EJ5+yiRdkkFXlA
7IYSFYwgUgmFZ5BDuriWALWLwDoFOaqlvjENI2iaBFJb8lbOQ3T/339zFDu19oXt
/UKVybfypvbhdRJNzfTbul2G+lu5NQJaZK85PF/Nkf30rXdTblcNB5wvoXeV0hyl
ban4Ekd/GAaoEht9UEgqaHqW4KbFQrnaJwpcr3tyrDuJ1Nv2UnCeSTb5FCJXj3bU
/0hPAvoxjk0i/FUcvpsg/uXsI+KplLYksRfHj4WEg3P2kZNa/TA7THcGkDqEoV+w
ojaqKtpHdu1wJxQfdQZY54fCmFvgj/hNEdD156vmlZTts/wq9oW6IEc2cfvPBdsi
Rt/ie5fmHgJW2UCwUZDKeabp38iXZSzkJkfyl/M5tnTnQsOw/Fq47RwCJLXE6ugo
QBVxyyP5jmWRXZy5S+QJc8YRKpklYZs7J0OFxdqo87leYCz3De4oIG0TIXm0Ni2P
RR3qgbdOp23afnIZI7ncVGHAqi0jhS6maoW82C9+FrrTGzaxqm5t6M88C791zk0s
L5C9fV14bOdZLqRnD/BCwTYBlKSR6UO81GmMTF2bi4h8ZF6FJxbUSW/DtvoLzeFZ
zwb6x4fV5XD398Y9gDDgMLMrnUzncHGPxwLz8t9win36TtWxdt1uedMdEmpjcHq4
mM3Mj79i9EMMWBZXHvGg1EN/vTG9RbY0t3aAAeLxZNDooa3C7gwqLT05ZssJRuvY
1zkwxKDyRA3prsuK+K9CUWrTFDz8+6BZ8hwXOYmvxU0adljCfktt3sHEjfa2K6zy
4YtXCqyMQ5BgSpeTXTi8wJxjmWfsw86mqW07mMKE+kGlJDoWkdj/NfKri/RjHe/K
cpVzPfyQjX62dQI8/XwKv3gjuAgyAT/nW6qALTmXTJ2XYWtuwaFURVRPlCQzqX0S
kWXziC4eN8t7s5jMJFfD5f0eLWZ+16XfMP/VB0W6U05zDf2dyUrmqN2CUOQCfLGU
vWw+3qBfl/dxxTlmXE/5LYzk4c2J7UGLeVOHOUVJRAJExjMBgHmSapjkNgKYmV/j
d/p7NkNwHdqWtv8BWfmfJSJ/CfKF8SzDXpgY3eHTH9tfyvNprV5315H/scrcscFT
XA79Iv+xA8xMjrhyUs60JwIeriNX0YpylezMNNC1h47zZy+kbJCoAMB94iGML928
VwE1Hs+NpzkeqlCIvpNgXcNG+oChnbIeab501/G1J6ttDAWlWWnkBCyQSpEIHb19
j6BTiu0UcaDVV29Lv9nzxeI7reDYPc4OgdoQyfjV18id6MVcAXPUWHsEQ6mmMZ6G
9FLiWz99ZKfGkV+9TwVW5UKYPofP86zZrIy1OnJmN2ZfK+ClOAT2riVkdSjD+u11
8214G/VB93uX7M4TveOlt6bfbQ9qNw2MJmbRhyT2EygyTI0V/C6afyXw2/MxCaSO
N1uPLww5KoV4U5ynxe6SKSWasVn0XktkClr4snGiuH7jDxJ9SnPx5Dh/3FMnnx9/
CUYNi4nJ6ksZlckTkq2zqiRnSj3Xnv8mkM5iNnF79bSa3gmU2t4IvvvOsSYkQEz6
wADtYbMgmkZ9SpO3RY0Q/35xokuc9uWVHYp0kO7hGWT1Tx86uXfx/drptXGAQsGd
55yvuDwdk4wO+LpLLMr+ehnb+DWu2KhJlPm2Ca2h654K8mAgXYVHrqS5075wISQf
C9SfTyvk47PHr8tnwncbBUZbms355Om2SpKSNt+Z+3VZtA/PknrfNgCgZtnIR5YG
rulJfiAuE5AiZDId2vQUx4J4K9uOVUdxrYlZGVg+FLOdL5CjAkKv2gOBQvCJQT+L
fKNL+oSZpqcCkTjUeE1YQpPZH1sqC2DP8gJyHoYG3O+td42P9MLvG/G0704h/dhj
JsIXanxPJV7uIU/wk/3VjvOTj4o6m4LmwnBltTHV/zGtRyc/fvG4vRyjD7TQ9VeG
RitShFnrIW9/IUHQiPr+YPwJ0I8hl4pbF/OjhFosfpYwT4RoAawSblJqqzJoQghb
oXpuhmB5V8IkswNd/19eomTEiWYlN7RPSSh0ByE7um3PgqjvWLxiTrbJbL0YA0sD
Emrz8NfP2nI4nhQ1xCXGSYXqJcOHfJQ/5zwUiqBRN4DV1rQ0mACmsbh+1QFNKvlP
O/mTKTt0iCYMSw2bm3OXvQAle4SOWl62LvBCcGn5NoRpITH1VY5I6et/Y7+a6LhG
n066tyQZPDUobHJlnUyAM/5V0XyIXyrehnktj38Vp+Rh3NhsSM1mmjvRT5EHUhPM
4YeEXHAZH/u5eqYJiy/3na91DSM5dhXbWrWJh885CkPVfEOYK81O2SMchj03e8Yc
pnJwAgZwquZBlbuQg3ES2srCiTt1CXwS8YfK5tCZ12JUxZfvc9TVo3+NxxqQy7aJ
MIHmTqLBbbnsgZA5iTm5RkVxjRGBhjzh/t8IKz2JmDObSu5habQTXOyFtA7Eoj5e
9VWeuMdWluFBcESSbEJfXGlBbVAci9EaQvbvWV3L01SBI/pZuIBi6F79x1eXmStk
DUjE6I2w6uECj2lZ50ECKX7uJz9eIZOyn1MdZuAwQy9OH6CsrpA0VMUW+k9dlMZt
5QpXrpz+nrn6XP+KPxzQGIS9j6hewly1SF8rI+w8yXyxmx13SZILNnwV4Lh8NrQR
a/Z6i+hp5ebUgUvTC2rCmrCMfcnN/vve+2MFFOj5rDXqkSsnt/s9/qOOwHQXA4T/
mzn4AALdg2+ByDyAQkwEmtiJHWJQJXc2obFt9MnDZmpLBbVHyUrBneObjKXy39EJ
ujvtm4Ye1Ozj3wAPD42RmfPgtK7QVdFfkUxzpTDV3Pl3aKAcTxC8R4m+LOpSiSUx
TacPG11lT7SP5JlfCCVeQsOk7vbzGtXdOL1/N6MWoVqDSqkOiituKcymjyz2Ejdb
EgCLY09Br7+OAQmXoPNQQeVZMzANR8wAYwCQZDZTPuxJZC+cgPliHgw2i/f1SYo6
38BAF1RvXQSNXEH8IiAugswK0ca0q2c0WZaQ2C71z/AufGU3lmo1FB7i/KIDwLhS
bjjuWdTsg4+vZcNwyF6KdaNtx+kezV1x6wrMETsVyqi+LP//NtLYZ90VZNB/ihIk
OQSwz5kqM/9pXJzs6oNFdF/mbOMngbgCxDSnDh9kkZ2dT/y6qr20qJ0mL+cZxSLw
enHgvQeuqU7cdd1o0pJdvKFu5lZoN5aAVDfM/rJjdHIRVtYljtm5PMno7BzLrUgO
uAcwZSR91aF0wxs38Urcl57+vFSvefygfOAdImRdNHkSci5vUeewn1RGA9NL+/Mc
R4Qax6IeCNXU2ZRPBBF/x5/HrV3VXA+7Z1adst+Ow1X2g2MgGHuVwqkCYwXzTkgA
NwjnNJPjLj9H6Spp7G/zrEpU/FM5bMqGvzYlFBjhDNiw0LR7k0nKfisArzSXQxVr
o9Hsg/e5gauJ3xR0iX3AfLDnHcVnNWhBjIQmp5aIDBXHaE6BoMWxVisVSf2W0Wus
Ch1lgcHSkhSBZTrV7+sM6HvUomsOVJpZJyR61xgubKujq8eW8LhSFI8noT38rOsD
wn651TDak3mIN9z+2jruwb1Lx+tpY10NAsh5JOG+BABJGLSTDi5zKd/O3zHR3v0O
dPTaMmqnSyf3gi9U6lDXmyylhusN9UPLC4JwvmglymP0oPzn2JU7ayR77ctYsTvb
oIfppj3KaWnqF81bAK2/6fjRyMMUjrZnED7cEgB3lFirW/xDZnxtGB0RqclMmC5S
7OrcibzJ+10j1oXHEXCGisGtK0MJqIZVVdl64yEgJ2RkgUf7nTMrNgx/9o9Nw8jJ
Cru9uHH5cJFnFGpNtE76goZfYZY5kJVlPQwb227IZ2c2zyoOlTjQNzvOzBNf/ljI
adClsjUxpWaX3QHbL+AXMhZuEJRacAgq9VjacQMgrS/Fm4X+yL/zf8lnXH3cmMew
pqIdElP0Ri4axT1rbve0sIiGBS8iodJhvUQzYFDLNwPoCRVwvgUqQHk5qeWe5bFe
1/8nf2tuZWRVuko86s7AR/6BVJp3LApJWb9Gy2Qizm6VvI7ZZUu37vhktEnGi/4Y
2WshNWbDJAwuOyiLCJvEkTAoVwJr5Co8Ja2C1xPqM/K8C3lGnWQz/QoHYAaK3nbW
TpyBEf8Yx4WXPOQU7J9HQbU7gZbh1KWiob99FHY5pi0SrmUWcPFaUjISUkkiOyM9
yoiqVRyaX+D/FMHQRZTgx0QWO4f9TOhcdLX5hQH1KJ6MHUD/CzmU0UbeLKZ5jte2
wpVy3T033rvNcDQnXtup9+5qE1eL8lURuZhqeMHfZS0w55pP9jfu0qTjT4BYvBrP
jwe8BLgoSYuW4s365c43wXwaKGDtNf0boxNLXOQqqdzmPtHvJQvPPE2GjPW/+8Qi
KBRaQEScNyzOEfpHfmbP9G5yDew1s29ny8JGeFqbTn0a/Z5uPAvl+/fNiJXLP5J7
igtPUvgk/1EqTrApC5ybM2HCOCyat5AyWkuROLEAyO+DwpPTsom7j8ydW/mZe5lh
6ejTa6T9FY0pW/ipUMdPF04gRCiFu2g+v7OnaXA76mcHtOTXih6tVP45Z5PRJM6q
ZtUc8bX7jgp8Paeb8s79+Xb6glNUFr6P44DDEDVkoBaBCyRlVIXlw/E3i7OX31mG
+AkEtZe00avs5sP37G8nUFN9X0tByGTdjR4xHUfp2n6a++xWZ7cCKenQB3DAAZgt
acJO4lcWvN6ZyRxqaSju2ppB+dkszYvC5YMy94JZhwFFaLo41Gtu6VmqrPaOyQAd
W4imvQjQq8CX8+PMAKTR0h+rrP1VrUQQ0Qqt1tw/+KIVTSP9scklnuIRveYDEO1z
vPZJjX4UFcVF+/5T+8EdVma4l23QGlUTLLJh4shgjVQO0n7iNUsChyj4eZb2Fqg+
AzxDkZ2jmL9CCxbH2Z8nOYRHfjyia7MGe7dWGdMy+TFa51BnymJTCbnKPBXrszF+
BqazGHukuyIsOGJg4YWOU9buQuGQSuf1iRCmy87Lnz4nH4pKUCtUBVVK8gUimyTc
yEGDesefFcu3vI/6GXf6aZlj3BPsTTFF/7wRDsGPoHID5ihvWyJQCDE+3FBjJGuD
NoM5/hR0TF7aQkEJf7roGBzfZCOrlYiGq0WuNqZ+NXyR7O8nMjxxeQTBrBKWFx0K
ltSvx3ql9G3EC02SgnE+O0+Oz9FP1Dlpq4CvZB21Ow5m4IlWKX+HmyykJD9U7/J0
BfY2wmLHWkmZIApAiyW6ewd6VBoAmHyDzJMFDDjAVtmJfHfzPETn6b+rMtcMFOt9
+n79RuCKMuwRkzCIqrpkofocCySkfMe/YdusnOGiMMtOeMfkVYruGEcgxDupw4Er
9cuxaGU6Hr+jBkZKD1XWCbcMNlU4nzYaPGD0PIPWd9vfIxhZ7JSXk22xj7BAVCWq
+KxTxtqFAx+ghYtGuqSIXCLiYJ5np4htNeF0pBMDPTNWFx/WJTxbmLsmTZeoJHKO
fkjHXlxDOauV6Bbldst0wmUsHxEaAOhknsC2dH5PuO2EfaRMxlwmQxpOmtqnY18c
egdEUBDq9U+5hd2GMe0tPJDzZJnqpKEzTeFzKFEmPyrjrPBkCd7l+hNO+LSDhjut
r8IDQl8pemLHaGC0PVAVbMWaW3qRZG3SaGG+DVcTCq9VSaDNmdbYoFQ8egVlJs8p
bP367l/TRfou30K8fICzl843tyjXUMXYuQ+2qVHMXN74/MIgn8wUYe0Fa6vYbRKX
L8UzKVjt61bDc+Lcyc3ecQSAL8qkFmOUT04puEqi+rsALwLXu1ZM4sEc6wfkkvIu
GSx755Zxdq8viUUYMFySWDvfbe50xYjtbd9LG0+dDeXka0j4AlWPFCkwBLfyVxYD
70Jj8id1y8fAkLXlVhfolDZANUAPtqlQXSUr/qMCH9hCX2TVdVducaUFLtdzF0a4
dNBhs9tMr44QpMUekd1RXM6VdeudQ5wGB6ugoOb/kCipVZmFygCdn2RirdrQUqW6
3H5/ODgVN43RIfToye5Liv6udw7zp892DutKpfAMCsSRsG11ljSJ8wa8qCKmNIPx
lN7LyK1sJ9OUXPdrGV9s1ITwVk7Cy6rFNYJUdxpWVLjiBtTntqKXg9jqs0y4czkj
kmAjFbI9rsVUMSapojcxZtCaDizDKpGC806ecizdjdNO9tTuONAmSCGnIEzSLLvn
hVZx/rcvNs6hHF5nedRGMHtkQ9150gO0eGk0mpN7E+hLPmpAldYqjbqiwUtODOZF
TDwB38FDUKXhBXjPU3xN9BybK04NBaf8qZoE8NOqT5x1VSnUNjuzIXD7KniNKfiU
abWy5DSDGIOVOBG948qzdv4tyBamV5QgP/m7gZwje3Dry6JaTZBEQheUAPz2FSYA
X3ATvFfQ8tW4h/Os6K6578ATzdSH480UQLmebYjzQKjSrH4qAY3JF4ySvqqrXEDc
+QCaDjGvgNrdXcBzr1vTB7YzNfG4b31NcwHjGaxiqJUSrR0OsSkzoYSID4xNVO9A
SLaTX3OXTFsKveNbclbZ7PKRlLqeZFGk3S0hsOrzbIaDfOxghW8XWeO7730ILHya
NCEQaSROmeZo/P4YDOlfxBtyimk1lCwik+D5oLgnEtlQpAjktnryR3vZ9hK7CikK
pKiKFiA2GMVmW8rIqTFuIb+kE0KnYzfGM1uY+meib0tA2RLNrKE+VKJ7h0p1K5V5
WK8VdJSdAJ7MEMc2KQ6M0wLPFNAEjWoFKMOlGSRvTxzEMVJwzjZ9FCPf+qKncewx
76gGodNVvyJG2jw4a/wp8aidgkwrzeW4uJq93Is7GekOk46uIn5PBpcB6c/mv5zo
u1H3/oqK5hgz0IN/2qt4GkMjo/lglmlpqa6U1lSAB7Iowemv4T3N4uZHt4iLe1Vs
itASUBeS3ynqyVOL5XfW8Oxm/1tl8ohj63PK6Yn8eWbidsvMIlJJqQFsG6OykArv
rGL1EpgYf9RTD5L0Nl8yy34XhzT8/2z7C7/9U8LAdsOoBtvkVB3WWFtKMdEhWEDk
OzhAz+uGk7izYuG0GUBKsd21amv4ShbQEz1zcJL44o6SElK89W4hx/azNTamFZ1f
sdF7LOBmugUFRqGGiCU4SbIEm15qILQdgLm+Kvv1Ap3FCSxGL2XHTNh/eaU4hmwR
1VnXiM/68HCDUaxtM35JC+jmhYveXGOv/Hy6QDPewpMmApYDUbR4pw/wRYveoN4Z
F20uBUBvK662FlqiVISVmn1zIXOUO8mdzVRwQU5+WJ80oiTV9nOJH3Dc9pc61pq5
qJMN89mWx7u65UosBrGfkfMREGyVIY1uFS12EZR4xrZXXWP+80twL+nUufrDVjHF
ediEC4SJFjcVa2mooWYIYg==
`protect END_PROTECTED
