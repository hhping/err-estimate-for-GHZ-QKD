`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CC4THEAsFtEoPSJos0IU4kC8LtGoKpumNz5+IDVHheuRZjkCab2h7bDWEBcTFh3V
sH0AAlN4ao/+H5dgaMVZ/7rdkyrivk5wAus0Zj1vWy/k6vBJdDTGK/cABwo6iaPL
H9f/BIymPX/3DXxY5dAFkoh7ATvw/+QxpBQiX6ZZEn4T7SnyjOx8bflT/xziEcj9
liLWnEKeAxZKV7w7nBzuE71HLQK56HivCMIOTsKr4GofZOQtfgXGa/wPs+CEKEx8
gRRC7DPYEiiPBLfsToL8ttjncpWWLH06x9+oqHH5BrG69gcbSfYUEre84A2Wzch8
cYki6qFj+UCc5VruhGXW3dxsgIvNG7BoEZRT11zzYMICR/ZO10RWTK9NzaHh5b8L
`protect END_PROTECTED
