`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oQzviZ2oG/FPSN3rVm4hAi/dnRB+spL6ioub4xIWIc+fzc2YZb279Ng/6A1TRIx6
Le1IK2KizY7R+hXwye0dlL0Juv0eSoHEZFM8xmXt0T0/ITRK08vX5lSck0s0MC6U
h+UQm/1VNS4s9LOr290nb9Cx5NrKJmdIOo4y6HghrUG6PBXUHazlBOq/vM/AmSrD
fEZODV0K9uPYs12n30dIpd6rTJB449nvpAxL5NaI4OOBlrHCpp/mrfhuSJ3VBIGh
am53Y0UCa/eOxg+n+u5v2O0VrKklgDpJ1oFJ0cEbWNHptq9PofGYNOUtwoMxjGYn
RcQpKLBLjwKi1cDfqGkrXUuFZ3oafm7AjguZNK/ph2G3kYAtT9v+4B5NbR22FvGo
xk8DbO9Jm9t6o6/853iq+GnxsYrKpN18aDIesOUg1XWH2nfKmgMDPXFmLIuath/p
p4BAlNQJGjy5q2qWvAMuEY7O/8gdEDiSD+evOg50N9HX6r1Xi2uA53ZYPxeaXeAa
jV9fIz40UL9QNXC6VnQH1l/OrkhmEGGSHt6XEkHqiDz84hA9mlzNH/n9+pwO4q7f
LoS10PopEDlg6+BofWtwRG5Ad/9WTOk/FzvVTxcKd8XRQYQB+uQhNgNjLe81174c
og65VmHYAhGdP3N22uaBAO9FTPDSn1ujggYAfjYZ7byfGuT/zJJ+a4I8Sh1zMy4D
16P1GOpw4ZyyKhNTZzJERlcJisXkFV3LBRMqE5CtmkUqeG0AIaEEmF3D07K7uYvM
hWHSusqOIHS4kyG1YsS2ufkU7pk0PK666KJvvihzLITTXwoamrK4cheFwjy3m2Gw
KHoOFc6RHyJ5izjZ/XNl0KUFEi6MlwsGjmHzGbuT70XT8FjlkFA1Jgo02oWN2sf6
EGKO//OXfP6gO/8nOgRa3XjE/NKf7XesV5/bPKWFYfam8jFjdZ2VRHZetZYmi+BP
O4/1d4ndluezpATlK1sUNRxjkE3bg1uvlt3nB8u1vqnDWn9hps0YL3aDDbe6YlLk
sbCx80niGrvjDBmTg5rjLkzsL1UlN+ZkLi1O3+4J1Hln6vpw+6uiQQkuhHo9SrjQ
RGZLEHywsQ0jUnQZ+cGk8knKS/7ZGClTiQhoRAuwcQojRF7KrfPPr4a3zhfCkXbL
xPnjdZxhKkE0I8G/oz/BGtT1tHQh/lUKZ29CN5nfci3dRBC9nhWKRlXZCMixnv2h
0F55VCHoVSBNnHQ98x74E4Dgpuw9r+V5hpY9AyzTadDdaXdkR8Zge/iy5yZW7V19
OWgERbPjhpZXOF7Qn5OWB9n4QQw9lGbQ/C/ZEAcpgoSn/DXVzkcegwbGO5ZIBvMC
LVGlqR+fetOrydz1hQUkdBB3LuhBMp6G0tzxOqbtJrbSHx/mxMUqH598CrUDlMXp
hfZWjP/JzsgKNGxXE2JEOcnQ2B3VccOYgOa4/d+ljktPdypT38YfXZN+7QU06uYo
FppbNIYkpTMPB/AnENNMG2cPzhbOs1dyeDcNRNupSBrCwkmJ5fiDy5s843chltFW
n3nLlQ02S5nLxXoVdKwcTQl47MMKM1cDv8peAymxenbOGdDI2jgZxCAJrRxhzGRF
1nNK72TQPb/wrz25mogLf+SVTK1zGLsMOliWL3Z+BqCt0Cpc+kXmxEYUEcp7+70j
uOk0EJT7LHgsQT3vlXKo96LdJbneG9JLRkXtV/we9IbxwKbkpjPF7pUU6u9HiDaT
Y+AugigwvSZ9CKxdlubPrH9tgwB1ATQtUMTlk+HA7DnporufkuHWcgkdwSczi63+
plVt6msVlHrDA25t6R3+jQmKKIf/9K7SGCAMFl57EW1hALvYonQkIg4D4dUwDfgt
eel2keS9btfJka+z8iqsZcwbhuH/mI0UiEzlFzKRR7GB733IpMi/27vw/Ozu7fbG
A3yryeaWK1uXPdZdN8subZ+xHqvQHFY8qDV7AaujkYFLjIAk5Ndu7rWr5bs2rduK
ySJi2Pgr7uTDwErM/KuTZc5atB3CmlNUFJTDnThRY9jTLuc95jyGka+waFdJcl5i
9slmayqNN3+tkoXZM7jEj33QqvnwLVwpboUVJbP7hPh8dmW/Xw/ReyYFfKk45KMO
tj8deOfiSI1EnS7tKrGqdu512Qnwc6aDhSML3uQssfcq5D0K4ufjA4qy5mIb23jL
`protect END_PROTECTED
