`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7ZICBtkeRvWbKQEq9gi63ezcghFViQSA9j4gCLPjgpqQAJUY83Boci6NiElblWfk
vWkrFcmdMBN1NAtvDPLZkoIHSfSq0O+2rUPcp7yO6ndgn7LoIe2K6eRuxw2lCmNW
ypLgyzh8FmmBXxIoo+37c30cIMaWnCBC/BX0xjhp+UtfDUdcXHTdAwmazwph3H8A
K7AdVuZy8FLbDwtRkleVs/zZ1E/JtgyIH6PySZJwb/9ki2TA9Z9z6CQ3ZtGgGhBL
6QTUFQwX5Rv8NGc6mU/eHHIfPTk4hbuWw8Veb9dyl/7n3W1+rg7kAu/2lTtlkdtz
a5CtQXUIxKmQdJHLCcXiFg==
`protect END_PROTECTED
