`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Gq1bXm1mE2w/Q5qaY7q6HXFzUyDrSD811WCQfP/e/kgJiVGXbNk0B+rzIP/r+6f
tqOKB0+yDwmyNvDGEaeh3q0DLBkrFfkKq7yc6aeW7n+00imXDnsw4SRncaq/9rCm
MCVGs6C8N7t9w1Hid4ptNNrSE97lmnnm363o6kPus37Xr9OoNQK6lJakTQGukhw0
bYxAdLtnXx3Il1By7U6qdE7idjPeEGcTw/bbSt5TfmeFhGm5kV2o6XZwjDfCcn7L
DuOv22ZI6rKJCmxaKGEIIWnnfZNcc2xEiG/H87hIUHAVptm6uVrYKkgytYa9Hgj9
rtTTZq7yyl6/z8AIAf216aaV/865Vrex7r97CpFoQoVMoWIpH5ka9q6j3im9JeeG
IPCg/cmR2p8e8Sqvzt6iowBex/peTq2ne4yKTCuno+koIULBurM7aP0dW4yUzHDW
33E73hoanvnKDvy0vA9kqcuSOC8Ltwc9mjrYRDVyvaMQrmHjqfFKvEAPHvcW0E43
ET2AM8UXE93PGjlc6yO4oLJ37rHBEimotyvGbgr8FWKv6aLuLSQh26Q71aDHaeJV
Nfxe+Yl2RJkhHU7AorLcJ0LVxBDQeEGk226/qg+HG9NruQXN3iLNIJkoIfJuoHa5
tIaCcnn0sH9jblX0eH+U1y42jVbmIea4zGkY0ypzGLOFqrdxGfeG0HX+vRojon4P
WjFpH/Fj+ZEWY2JcFRzgId8Rt4ebZCx3izsj7C42Kbtp2la2uS9Lxc7mFS+zY0Na
pE4dvCh8JQfXIK+sfdf/s1V9G1Edb2lXRQzyKawto1ciDCr7zlzyCRI85mFN3LdD
5SMmA8sPE01LA4LAXrdXnCExhjbftoJ/aMLnLHix1Su0TT+1aEmuWCJDsq9TAsro
Bd+CJLLDxcczG5KKoFWigAHE1IDoUFwIqWiIcY+Wg7q8cu5nCcJ7egWi7YTDOAyc
u7quaBcora/1QthBYwZyOhLKmeRuSuPMXkKbyAM3t5Y7/aCW18i++5QWpOJZUu/q
H6IoqLhmBZZCJspH63RLbA4FzQRwa4ctOB/Yxl26T/WjLeGEJh8nmRpII6frtGlr
r+051hFoAO9Wgy9dlpAFPI1H4R6gWKuuF7AVC8fk/npaw0kaP/M0kL7B1+3qtdAN
0oa96xtFuUixLFRb8pWfXO+SrFAvuxlVQ2kA7f3cM4ozVk5zuzZTWsWlBSJMOu+d
LHszPwmnZE/gw1O4B+1soDWJgb6a2Tmf84wQkXS+9+Q=
`protect END_PROTECTED
