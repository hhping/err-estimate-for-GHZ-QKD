`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fig0+zQbGtEcg3zBKmb4QP9z2ZqI/YtEOI3G70/bem7kaAc69YCfCr7uEEOuDbWb
lQbLIFSFJoeXYMt1HLFq85f2XqIjWBIAAs5SbfCUnxPNAJ2S2IyE3bCPMpX5JRjw
Dh1OY4UTC7owJHEXbI0lYhyLK79kECL0NvPplP0z0HzXQKA8HIAjFyJxyzwlGXPk
1z28j/lh81KCaZuM9Ou1AZkmma8n1T+4YARmhr77Yrnb0Ad3/SH1d5CgC367xrqj
xYTkEgV6Ww1vdADDhWZ/BFX2oo/YLN+lnq2Y2JUJshLboF/B23hvJaavzFJDc9YS
zsykwdHAU1u0Zm9UTWD9Wo2KK5WhucTMSbODnJcugDbWCC0Ayi1+fx8w9Js6vLWD
SBvV74wyxsiJm8UVYX2HyJnS6PsZPnI4EwpSR8DrPASyHdIlLyjooFDtVQqTjmoW
Xk80V6RsmhbHB7Ck00nePIU5IErcj04XXdvDlejoLE1U1HRAo9pgqHrJ3zPLbgwq
1pmV9dSRVxdaY0Fzo8NMsqR6y/sDk7VQ6wkLH84UJOeTQFeP0464fNdMF3j6ZZRV
v6i4UdcW4AELs0QMfmM91gDPy9V4h5K/2NqYpnhvU04iIIbs6H1noQ24D7TEpo3I
Bo2JDM+Ioo+bIPNPnIKn2DrUVPkya3LeRXDzquHtOWpVYlgumDUF4NOWhOVkVnDA
Te0doBvbWySoZyflFajunwW9zs+gnLzYjMWyJAczkUcr2RHND8n56Y+P4KII5kTu
uytg0xuaN7mPCpCjAmOdOGD5VcBylmE3nf3toLMfFZqTDKs/4nR3zza5nnAooWUD
T6kdX9iaer50Z3/ccAag2s068RgtfbPeIrATvV/xEgt0GT7a2qRAU8guK/ZCxuXg
qDotjn+pYryxEIhWj6vd2OWgHgl7BMMHj/cqDANdgfCSuX5Ogv2d2IedIFkrxn9F
x6iRWfo3ECIsExlioqbzFuArm0nGO803bk39arHO6tnqMhq1oLGrv9CsNgoXuj6F
idqsJhb2YLi030IN5Lvup8xBpWmVQngOlAUTfiWf513x+mvnps2109zpp3QKhL4w
StTelouSjWkxnvy2HF0Txmqimx/I9rYbAbjqoN+4E3cI61BPNI1SAsYHMeOkdTmQ
pgdl/Jn6EH9FRectzjph5w==
`protect END_PROTECTED
