library verilog;
use verilog.vl_types.all;
entity twentynm_hssi_pma_rx_odi is
    generic(
        enable_debug_info: string  := "true";
        clk_dcd_bypass  : string  := "no_bypass";
        datarate        : string  := "0 bps";
        enable_odi      : string  := "power_down_eye";
        initial_settings: string  := "false";
        invert_dfe_vref : string  := "no_inversion";
        monitor_bw_sel  : string  := "bw_1";
        oc_sa_c0        : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        oc_sa_c180      : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        optimal         : string  := "true";
        phase_steps_64_vs_128: string  := "phase_steps_64";
        phase_steps_sel : string  := "step40";
        power_mode      : string  := "low_power";
        prot_mode       : string  := "basic_rx";
        sel_oc_en       : string  := "off_canc_disable";
        silicon_rev     : string  := "20nm5es";
        step_ctrl_sel   : string  := "feedback_mode";
        sup_mode        : string  := "user_mode";
        v_vert_sel      : string  := "plus";
        v_vert_threshold_scaling: string  := "scale_3";
        vert_threshold  : string  := "vert_0"
    );
    port(
        avmmaddress     : in     vl_logic_vector(8 downto 0);
        avmmclk         : in     vl_logic;
        avmmread        : in     vl_logic;
        avmmrstn        : in     vl_logic;
        avmmwrite       : in     vl_logic;
        avmmwritedata   : in     vl_logic_vector(7 downto 0);
        clk0            : in     vl_logic;
        clk180          : in     vl_logic;
        clk270          : in     vl_logic;
        clk90           : in     vl_logic;
        it50u           : in     vl_logic;
        it50u2          : in     vl_logic;
        it50u4          : in     vl_logic;
        odi_atb_sel     : in     vl_logic_vector(2 downto 0);
        odi_dft_clr     : in     vl_logic;
        odi_latch_clk   : in     vl_logic;
        odi_shift_clk   : in     vl_logic;
        odi_shift_in    : in     vl_logic;
        rx_n            : in     vl_logic;
        rx_p            : in     vl_logic;
        rxn_sum         : in     vl_logic;
        rxp_sum         : in     vl_logic;
        spec_vrefh      : in     vl_logic;
        spec_vrefl      : in     vl_logic;
        vcm_vref        : in     vl_logic;
        vertical_fb     : in     vl_logic_vector(4 downto 0);
        avmmreaddata    : out    vl_logic_vector(7 downto 0);
        blockselect     : out    vl_logic;
        atb0            : out    vl_logic;
        atb1            : out    vl_logic;
        clk0_eye        : out    vl_logic;
        clk0_eye_lb     : out    vl_logic;
        clk180_eye      : out    vl_logic;
        clk180_eye_lb   : out    vl_logic;
        de_eye          : out    vl_logic;
        deb_eye         : out    vl_logic;
        do_eye          : out    vl_logic;
        dob_eye         : out    vl_logic;
        odi_en          : out    vl_logic;
        odi_oc_tstmx    : out    vl_logic_vector(1 downto 0);
        tdr_en          : out    vl_logic;
        vref_sel_out    : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of enable_debug_info : constant is 1;
    attribute mti_svvh_generic_type of clk_dcd_bypass : constant is 1;
    attribute mti_svvh_generic_type of datarate : constant is 1;
    attribute mti_svvh_generic_type of enable_odi : constant is 1;
    attribute mti_svvh_generic_type of initial_settings : constant is 1;
    attribute mti_svvh_generic_type of invert_dfe_vref : constant is 1;
    attribute mti_svvh_generic_type of monitor_bw_sel : constant is 1;
    attribute mti_svvh_generic_type of oc_sa_c0 : constant is 1;
    attribute mti_svvh_generic_type of oc_sa_c180 : constant is 1;
    attribute mti_svvh_generic_type of optimal : constant is 1;
    attribute mti_svvh_generic_type of phase_steps_64_vs_128 : constant is 1;
    attribute mti_svvh_generic_type of phase_steps_sel : constant is 1;
    attribute mti_svvh_generic_type of power_mode : constant is 1;
    attribute mti_svvh_generic_type of prot_mode : constant is 1;
    attribute mti_svvh_generic_type of sel_oc_en : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
    attribute mti_svvh_generic_type of step_ctrl_sel : constant is 1;
    attribute mti_svvh_generic_type of sup_mode : constant is 1;
    attribute mti_svvh_generic_type of v_vert_sel : constant is 1;
    attribute mti_svvh_generic_type of v_vert_threshold_scaling : constant is 1;
    attribute mti_svvh_generic_type of vert_threshold : constant is 1;
end twentynm_hssi_pma_rx_odi;
