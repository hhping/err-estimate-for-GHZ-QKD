`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
osA0rD7Gbed6iOzwEEsl9zwzJsayHdUDj8ob7Hs/e3iRT7CyW0BTFt7X4qZU9JFw
nNU67QuNU5O3TZJtbBKNFGtUdSRmHT6pO5Z/xZCHtXneBJnOn6ptc1EOcTVWascN
uknCD+BVhSLy+y+2SkE2X2MT/A7Tj+8SQtz5pz+PoeSSb0A+auQb9IGm0OAsPmFF
MkAODl5i3b2K+dmWLZG66FwFBMMvX9TyK5TMSVfKiHdor5b4AkwKRsBwwnDFA1vQ
oq0WQh+wrRIXLjjLAey44sMK85+c2M8+EhwyNqABwD2TtnRUxpDXCkEln4tMzHbc
FmMmxl1hKCH3zA5TP+NFXPN+mgRUQINZSuDE5h2SkOxw/cQ2hp/tLobMuhC78nWG
jySWEWodjl12ajr7yxrZnC19yNufazcbmKkXMEfLEHKO1BqkSaKnFMbTCc2MlRJW
9ZAc/fX4P16OjtWFNNB/jKcA3fcDgX8NNP9XtDPOdIbZ8f37uKvKhpgMjHof2YsR
PSqOW5Rvp9wngTVRpGqCMn02popcK0AM8sL/GkHl9W3G1w4xfUqIYZ//4hlv3oT5
WCtXd7pFBv9OMpUbyabj1YOmHrLOzICh112r+4ngy9xPKI7JKXft65xuvBpSRvfQ
sRfzKW3Z2/o9+1nFiATI60skHFJ2Gdxkj4Tv8iBKvOS8bvWqoO/gVEkfVoVrogIJ
XQaUjHWkvye8m1I483HVhvEhXXvIr4L1nv11+G4zD8aVPK7BwtA/3hdbJywXSyy8
dmxYDVDE9RoYaYQ00QY4stLFnDnIp6103jGGwhdLDeuoMtUEsPI+Sz7rrN9mKpcj
LMjfbfCNITu8TMxINe/miQ0YXQ/YqolntZKiIUxSXlJ5TqaLtQIOQL6Nh3j6NryZ
nADEwThID481KtOpY51ISOIFZszKp7KuZEro4Z4EFc19rMkss7DI/uPx+01pPKBF
N9kNOS4+nY52MHCphgLrvg6blbM5Dlpyx5pkNAG9z/0ss62rA9w10SGGyxhAYLle
M/HcVQtZRLLX+vOBEFllMEOSAf/opFvurVO5U0mP0jmYTuXGpiQEoe2eZ/0thujw
H5Dp6db2Rn7Frpbg3w25nmJxIILsAmyT6LZj45fCxutOHddKbIO3JdawuGlHYt0F
3yQpW3BToEkHesKtN4+JBRFHvwoJwPzS+fCHPigWqfWETxE7C/tngGZDKIiQU6bj
`protect END_PROTECTED
