`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fEKGgHwxkfmtda1rjLb2S6+WU1IMc0ro1Q/6KF2ZVsb07/ntBMrW7u+JbVmSGaDB
/83LZwBYP0nZC7Mt5/M4dc1J60VOFpTtmVVdP809XbWgYfkjl/xANYgorjHccg4p
juF2fXKa7zXZheUmQCm1yppnL6YjBoXnkqTVrnnS4ozBzBy1wLXvPLX2K4ORfED8
4/ZvfDBvRnK0F+BIKw0g1lxjfZUeMNvD/MhZNuNy9lDAOl49UGiWI2yL3rFGPJTd
idnXTI5NBN8Iwa9Oxc21tYqPV+MNANRrDbI3Aj+8fPOfa74aQywSw8nDidBugX6a
sJq/CXly6wOtZhjpFf+8bcmqicNE7DpEVIN0e2ba2YXPyB/E/JWP0bPwAsUiOqqu
MAFk5LsYUfjdyiyaVZmIiAr5pA83TYOvaKRe5tHycX4ZEpm2K7CwHZibWaNgO6Od
UFIpcM/e6QaBLxfQflg9tfN1M6D2cU8g9XN2e1lQJ7793ShpyO347eePObHnRTnH
nZSojtl+Gq/r9H/roGeiMm7vWVaKoW4C0sPKlkn+5LsahFarXSPxo1Neks29s3ri
cQM6nzNTMcKCHaEnRA0Iw7S1kx8BmIpi/uhnNlRNhHVkxB33Hvp/bSA2zLdcvR+/
b3eUrOGs1DV7o9hCTlHxoEOrUpvV2+SD8DokQ+NOu/EdbY6PQXVpksoFGJUimn+A
Uxx66Tmk1jifvZCFzGgRDFbWKozn5dCEw+qTfWAEbvuN3iTCsJ/YzIWNRRrTW25P
`protect END_PROTECTED
