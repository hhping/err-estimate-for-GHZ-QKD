`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B21CGoWxqqFT68yv70V8+o8KxNo97Y6ZJZ2EfdElK9tvSpd/co5gcAiV1A37Z+u7
jz8k+RpKVwzylv6Rr6eDJg6d2qQs16xvhMRYUv/vsrbuHOj5s79dYWrFlIYyDuff
xJDxgEYQBOwnVAX/MRFtDS0+qPpQ64TQOsvew5x/knqFtXxd9F1fctNpEOdz+D+E
+bRS3NcDZDXzuVlt/CwLbJ3ovYsYka9EJYvwA+SLO9pAq4MqLxAooDO7URjx3id6
luiIWZtdp1HX51VyaWYjrmCN0psgNTo72wPTWsEBW3QLHRfpHIIbapfn4queH2y4
njMA++ChPgwJ22YwyUn3YRHKuCjd8MV7Bdoe1KHXMHOAKFxNWMO5dAK7WxvwgBuD
ZikZ14OJGPHjTgt1QfMF4i8vKA4HiqgnKwU9k65nmkOkx3SXMNaL4rHXcRYQC9yv
k2DKTb6cWC1UkfqoBy5q6Og7gwg/Igc85+kJpnq2t7X6ljxR3iqx8Kc5nGNwIK3b
3uRXuYlAsaNn29FG+0uaH2+VnYoCxrE7DtZMvWW1X1kxkQ9hyhhdn08mobCk3VvP
eAgjhuEBoH64KKSoyGwaRqYlam5u3txMhPacoGnjtX87WWDG2Ni9KLokDpSCOw5+
`protect END_PROTECTED
