`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b+hlfQSaYg+2Dj/ACV2pht0XtSF4J0ZqCBtxMis+gOmdFtb7FwaUV0PwaBoR39eS
oO8C3K9LGdGeqvZY7iLiNe41RGEFBUO10loNUo4bguymXnoGfa3SWp8raZZxAyTu
I+lG0T5aB2vupZDkl9ahHRVxV7qfMeh/UUOfr3NhswDb1OZU7FfmLvuVFyiHNFy+
iOA/2fIZ9LUMoNh/kkVInqK7FCzPNAm6Dnm8IArCqdn+OoK4aytSJmCK1ZAiDrC6
tKH8S3iCLPtnY4ax/PPGH/f0xpn7N870FX4wvjVtY/Mr1JGQOF/n8OIe2t4eebVh
n7KyM6W4HGC2cEiq948VQk9Vk74KL4lSqxluLmi/Z85JVuGt4FqlGr/Y3fRczGLD
78MWzKx7UJKu+IWGnS7XwosLGb/y8+QBnACdbTktiMNlVu+OXfFmV/IzAb7+JB5C
khjGz9SJP/sS35VWMpOE6VogehhDeWWw19y02q91EXzD93vVv0nhyHT2Z+XEZASA
qW6bfF6V6HEc+Yk2a43gBJabA5tEfOw0sz3wdw3DvB9B5ppD4U2z7/PpAcC/BmAx
TKs8CyTdbah+0IKOp6RR6w==
`protect END_PROTECTED
