`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wESACgVP+B5hkRsaTvFyEo00quBPlNbwqhxRWTy+f0LpsjxM6Aej9ZdoTzRXfDvI
quPpgIuQ96dIe+cSo7wTY7xpsGVtkFtwsWfxdjoQFXKGY39foJdZrTq/Q/HbeaJw
kaJeaASqQEErZsHLUN5EDblSMDOGahF0xwXDqGWnNjXA0Ik3p1QoqHayyP34mcML
mHVfqruX/CKxiO/orrpBs6jSOhD6Lni74OKRw3eW+xU+bJkp5uDRls17vwoEEuMx
34kr1wZa5F3czKaXjDDNaSZQ+/53HTYY2A1oLacNYVtXXUSynHAP+4q9yBW5HMp6
7E8ddCRemrJ7csOZA8jKF4XSy5pOQ3OJQFjgOF4oX+vtzVi8Xnrn8Ur4FEzLRKbq
hSb5csw03c3eDl0C/3nRF41EB5XjNTJap0O3qDAUVzRKRxLL6P0iSAyZyWBUrhYL
`protect END_PROTECTED
