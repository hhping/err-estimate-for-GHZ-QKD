`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GOEe0tGjD0LOn6kRb1CMvlzHsvHbV+q/XeSdglkxmnI+8kBzKhZYkZNgBRnmI4r+
ivYRJGdklm+cbUlWFuLXawEQJzJTmPLbmXc+Tfutwzvqk0tfg/jBMzzl58LQlDeu
qAaUbpMYb12t0rWm8MIXBzGI9Jq6j8zap+xGxtJ6D2eNSAeyK2MDSlBoRqgbyyFT
cWmsVBjFZ1QbroZnyatiJQxi3XNK0XIZJM6hmVTuQG/1gKCvYj6gmwLWMkVYS5La
Oq/Rucu4zwMJEhfYCPVZpag7zipWtdxSfHopXGEqqLROJ37UH82MMy2NQ/AOFBBC
KoOAKUEWIpn9PQEZCCAjH62c3oMSOlA089LC8Q/vv4WalThR9AtMeQObSm/ny1Qk
fls9n3xZ0fnLcJxU0XGe3fRmsHs1obGidUKcHrY4jtH15V+iadyizv85ozKXcWMI
tetcIo043/yJVsWkrg5T7kzknYLb4tRtOWz7ofiNxwvRSzzIHaEJPZqPVdqrnggA
FhbvJ6ILYauKV3UBVJASK2q/V6NwnDurt6pgXE+EglU/8CrlCpudnPls96/lCW45
g+MdZjoff2FcsX9jWPnFSpEWP6RWnuTmccdZpxQMViZkgFuS6spYN0GXi4ehaX6s
nDqHp9nDvK0rooXEsN+u2i1Fr7V1GAk7xz2zvquiDj92gsxJcnF/jFJ0RPyctqNd
9XOFjK3Vq8P+fjUiSNPavYqpCrfbM3w/YkTkMEMoyPz0Ks7fppyvbRCkHwy//rUz
npzSduN2FJExAE4cbWmJ4K++EEEtG3UHM/d+hK198xNln0V7ojeuWwavYQZJknPY
MM67CCptIvDrb79gRwL13bXZNVCjbb0oMtv8JbhrcePNttcFUpKnrQo+VZrZbwnE
DGOM3x4IVhQe8UOQThDjfbngy/686zz+7veDZ3xLntXnFDgGtcnQI8MHi7d9EcBw
ZkR6NTUomLCCeXj5vfWm5FRQ72Xf4oICjTdmZdj0/VC6jCj+2IGYKUaOgVBi7zS8
HEN70AaeebP+1eGN3rDOJQXo4Vnb3sswMbxp105hZO9eB7aqfpFm7fn7Ur7aOxZP
UOJSafH77pIsyj7rFzZAuk2lupDLYZOa9N8gk0TOksdqVHVP9EmU/H+qO3XT7+/v
lAl14/6KxTts2DGpBr1er8LC5oMbQCUgOk+Yrd+486jA1P5RAXBRQxQWZgJ3xxbv
BOkS9nFZVX/gK6CTwUBKMVhGfwv/6Osnx89udt1Avewv9b/M/NoWqVic0oT+Z0Kv
mE7pNrZ4jImm6d3ob1eE+hxWy/jDF4/65bTSncWGfVsWFS5Kw/yRV3lk307+XslU
N0ZQBcAM5y8j4EYZ7lD+q/OEyJLy2oNC7tLq6dvK8w95Q28OAQuswbQ5lKGpWx1c
AfSsSb2sF0ybEziV88ZGll1jH7aHZVkie31wyYso+07EvBelBhZ2zy+cPuzboYL8
ilil+epRfEHlAYNuE7BtOpQbUqRnt93bt4+7bNSmOMaUqIZlX4Pdcp4LgGM4HvWy
HFdsUeTbbXbkOFR5WkB+RSvUSN6GXtoI+STa183nDJhR+xQkbM6m7NHieW/2PULN
dJ9njGapi2yJphaWCaHy5dsfuwLttpOj57mkfrqu9eHoT7MOn3u3MJrRiZ+CxhLg
EG+LQDnIpu0a22ZDpLacMVxOKXpjpPfTt0fR8uI9V/l5vLM6V0ZuaGQqO7NUI+Xn
W77a/hXgb96hErWTOxNqhbO9LFtgEFr9STvok46AxWXCEguHbHnl+gw12XdTEMGf
sgDxs/5JJZx16/hjAs5AO8E/f9wXBsWdLzw6HBzHtGPUXw/yirUFRLFnwQswxeuK
Z7LnHKmMl7rKOhNwDS14tAYPy6sd91CDO3KeWclmmFyDkoyyyb5lDcwZNrgvu5xH
a/qK0SE0duS0WjAvCERmjbnlrBPWEmns9ZAhpUJITpGElbP87VZXv+K4/94OQRVT
PzTTmx3fR9ilS0zYD0Ha7QUHbEjjQIG92BjlUKeV5mzeAyVb7aZSr8zOGwxNbLbF
ggWkXIZ+GFhJfyGbbVEnSfo2ArR+RY7iJVmBCGAUMU3IE6nh786Md07E7kF2fayt
7u3IFJfaqb5EiaxT37XEN9o7yUGlQpzMwGBg25mpCHDq2n0ABorPqZ6HoMWhKoRF
Fc8vP+ClQNZAIyolNlnsI5xpGBnYwzbA95JMggAiVOuu80BTMEbxXqoYV2ULIs6A
aMCyGCHYKKnkMXqOM8fSaL4mwPWK4aU9CNQkQIVRl5bYaojo3wG3BlJZ41Nd1yEt
GNevKybIIypI1qjRimz+d5v9Od5CMOQoZjtY4aWC0kCUqgyFtgybm/rrFs4nYgST
sLFyRbLafKaoSM4kRlEDe7u/iQZ7HZkLM5K2PGVar1/GmGX+BMDhQ8R1eaDaJHG7
LGWSkpIJhgyzqJ5qr0h2EAc9FFqfJmLTnWiYgME0sdDuboAe6tlhUk8xK4zhkGIb
aaK18K1WsvAF1wcAG8qEHw==
`protect END_PROTECTED
