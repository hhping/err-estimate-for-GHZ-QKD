`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yHQ8mV1Q1pByIX0cKBK9vrv52uJfFpgH+pd4w0+3dQ3FHvUisOLFqe2OFjKXF6cT
KgLOzso30B/IiDkmRbm2qnPr1sMD82g6XmuQDBWCGTbVSNllQS4a+b0Uarpi4w6M
oPOaLsHBC8AFOfO8BkG8UxQrM1zckRcOAfjl3EsK+2xothrVhzzcv8H8zw91C8zR
W8wYHDjWTYUR7lYFraN4RODq3iFUw0a6/t1lyZOmcI6Fj3EwZY0GHCIFWspFWpVd
eWLqWCw5r8SZcwdpZMOGrGpZf/FM7ra6Hw3AmFzCHxVufV5P+zNdB3NyNUlX+gkt
j0ueC9i2oqgwxsT9d/m08542CrOZHzHAvoAR8YBhsnPDN4+LT7CYFfODZZJm8oOF
xnDtYHfZpFibxYzqZUvGf8etEzXky9dfd86HlOGD1aCwueJm4bbvcl4eb5nui/eS
aL+ccUIKnXYBgJoezVTViQ2UfcVEhOIIAXq51S7wZjMMmP58s/GHGxmyADZDXSQf
uaSR7NI1bgKvs5itV4VaXwAVkP024yx/rbR6tQOuCZdkqXz54W5l2zOpgTzQ/juh
25ZWVlj4W0ySZVQqtXrChnwI6LiBS3usmBv2RZWrpqzQcOtrZ2cXTU5MAqVh4YzI
IxH4T/ZWuDjZTJf+RM555NuQJCAgG3tkUYhNuvXqP9WM/WdK4aFHDw64sTYgwQv+
aGKtQYAXte6xoh48fW6WSybO6qJMWU5IAPln5lEi8z1tCjbynHZGkaiZe1YwlXhq
4k78+eAeQBtkAdPAk0FGRpSTtm/sPI68BcHeo5eNjqAEWWYrnNndB7GZ/6E/L0r9
TJM+T45xc9gvW9PkO5mhm7AGrOfRwSfE6/j5B24Fc0oXA/U+n1dIbFRNbmPNDFfe
Oimm+GaCnGAult5UcMRhD4Ddr0pib/LF5JWc30+7bSukW76lXP4uKO/vif2rqNX8
/bAVCeH3UNbDq0sAtClntzGQZvNHfndPuoREh9a/L+7jPEsHeQrbAbMlzGM+QbgA
RIf5N534J9zXuG7GKnzlmVydK0KwgEMBF1VQ2iGmc4gOKpOh5YqNAeNr3CfLDvhz
xW8lTxeVfEKvxO0hnanuAfOnCfTusmZadcUax634z+SS2yT2gDRZdK4M0uaSym0s
qxUj+RxmbaHZFvnYGBpwcIj+Jlfblds/5KkhEBBcNAiovaO3rNrFhE/x2vxD9ChD
xYH1QJbJ8HrCi32BVwcwSGDFnpYuhAvGp5GciXiUwIKguLML3uQQGthuJjQxDusZ
/OgAbnhMN8X+EYYZUfUwUh/+xjfNlevLqlTjI1L8UhI4P8Ye+Nupuh+C+Kw/Vni2
Z4PvEFsRCSwPpvPQIyE49Jw5nbOFYWTNBpMoWUXdqVUQ1fFEr79z2LV+pYDHZIMw
w4ooI/tMMDtxsppA7JBeUyfKWCHEQuKVESP8y/IJYqW7BK1Rl9lFlxRVCRg+BFQr
sEJp595QTmvsImhokJ7urS132jgFEU+y28feBSL9uqM+YRrpd9GabcaMipHo2HU1
GfqgOgI7mXnBRI4VnSv7UfIL4++1N9rom/xDaFT36ThL5J9Ko04yFMHypQYgS+8J
5pb7/jcZr3S8V4hUk5GtgH6mpP1Yb+TO6NT0rRCp8IxEUo0DgMQZnE+gbEBIF+5B
SAToWhM22cJPNZvnNOdz9VlCUmI/l5ba+cfAC9ibOFMhmCaK/hYnrOeBpWBXuZJc
9kTqihGwvlT9wO5dxD7v9XkurlEp+fmffS3w93lKqLtRBnPnhqA36ip+k9FawbDl
zVZuieTJ5Yop2Fl8VRY8aAlnJRBZkBauXr0y5KGYdaHgin9KlwZLMbqJ4O5D20Dd
KR6XXPj3xtNEVdtz7ZyLPq81AoLUXAX7MHxPv482dMWlUvEi6JNFy/eyuop7nOQK
DP3AkJBjbk1Ke0Jf1JdHMyeLR4xgRDXOW3yO99eziB06oKsnUkhLgFegbKZA3VBX
XKZSnMMZaSB3XfS1UwOCCebG03jiwisWwclM0TohSZPUEfRH9qY9n7rAfHD6h0Lc
ImMfbyMQKFC8tTJhtu4ACTJN9XGXjoYJy+NGnfJgrAp1wPZdsEAt9y36CRvpgZQs
`protect END_PROTECTED
