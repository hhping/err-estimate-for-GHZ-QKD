`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8KETOCbNmFL0XL+As3WBMX+HwyjHygQKUM43X0Mpd5nuJ5SIwTR6nzrv3OJAR2sE
fse24xMHWPHh96E2p5rW1nTg9gwThmVw527EiVCzzPkL5AC25fgF2uMtFy20bQ7I
V6pX+ycyIg5DzItjzdXywWhfGEoWgkhpsV+PohiwzawMJCY2Y94jgQHnurGj2OGj
1eV3Jeq9pXLNDrp62y5hW2ko9wi6Bi/S7plcuUPJeNHtn7KkrWkVRyKNFpcUlFgk
MQ7Wu8RR65l/0r5oLarRO9KWJXfMeY/so0cy3wvYDQ4q85czR8u1XTD7xCE4iPmE
Pfe80d2XV+OvRDEc8dfQST/fqvvdJa9J2OuZkN3OILEQzUm3rRwWr/Cb7yyXmzoG
BJtKwdCciJ3OpVCTzcX3BMzl38+u0KWDVOpeFJhUh3eFIXX7NHFHVJys5iD0otfm
yrweZUPmvrxz/frXo+Sly839IdDwlHtDgdXJCrsuB2Y7i245rY+w1J3HpDUBscH0
6Xoi3eLF38acM6GDEU4KnUETSLuEJAirIILV8Ccn/aXOVr4xI5ioJMvZBr53z2lE
4EGxM36XjkE0eNyzmbqhP0nlhqPkQSdIWmVLUCHLsr8Eya4z0HTSbEREcN56wUAc
y7C8q5GtADENp5JC3cLW9RTfhQnyKpBkjgEhdTXEqpnx6L9Fqd9Z4AykUu9KUoUA
VsNAmPMlIJwui+x6oXLz29P0GjbxBquX5aM/gpeYemK5wbaB3xAwB9kLej3RTHt9
ESa4gUKPo8652G9eWXCT1TCGJXSyAF56KlXakyBeSpNgTxBHDkmUR3hrS7vgVaAj
aJCb0Swn7ZazxSFRn/064piTrh2/40KQrAP3eI09U4sKF1e0g7ZHWFPIFRjHYDJu
+it0ZeK8+SD+tk9QW3IDu8SgMb+cLjO9gLvrlC9Zt63KkMfad62trb9UXhAfOmY2
HhN6aGMCPZirTlOG9mY/gAO9MyL6w2O/0EbkE6M9cSel3eVBq3XWKEiWNwTC8Kpo
tyZqHbNgytQKZcBGeXty8wzcvKOH8gjM2hUrONQJ43dRhMgpRVpGv1TtK/C5j0rA
DucWq/p7CVLrx6oLA6TeEeugQI5oI6DstzmL9RAj+Ap+JAJ6tlBEk6IkMKOqDsKO
Wm1sB3uzPrUdV2p0qJEllXQRiVJHjPcu4cS/uqwWPpvS5EOEZEUvGn/LFqIKhkoJ
kx/M1n7BMMeWcZYysnZHu728Mo4/4eZ77HNTBNM/QKmkxY+FxP6nblZUF2eCSu/y
Au9gSIMUqIvtO6vwkq8gOg1bqzN+MXar+am99pyzvQTCLzpEk0WxuIr5uv94nW8q
Bu4zHsqFDccUWM51XwuD//4yrwYNyxhVomGkbzyn6fxiZjzRor10wHylQqQ73cl4
gGhWV4nvdrfKZO9xdIjzz59NfQ2m+vLuJxdjxa3Fpar0r/ntM2+FkzQdB0WflEyj
qMpCNU22AD3cPKm1oizfgLAsgA17A+PJdjo7+3p1/LGDXSm/hijYeKHEILq1ivIO
qixFHrvcF9ZKo6lv0BI48bXTarzbQMBm41Gb4hDrY0KjvyDOSGY4/UyHsGXD6gNI
yDYByqBHzcy/IxdA/WjiHQQDl7NhftESVw3UY8hfYXTkl+xbecBsM+8Xkbo0vDbf
xNdzNbaYOPJ9spf19mOwdBkR2gwbMFEc5+xDbuK/anDkAI3gie+WmQQAtD/Y0wk5
gJ8m+QYzgOngUKIS5GMozOnq9jfqXRQA/YryVy6L8lzUMbnwWsnAycXQLPwGAzwM
qn8LXNsQBwR/1qDhE4hzaVeCId9DC8pe2qLIJTQyiVBOR413aHgTTZKMxDyoyeiB
cN/AA2ezHnZCqRSf8o+s2Rg0QGxIyWPcJnm88LC93W7njmP5UYNqV5c1+sH+CGVa
oL4cmnJPVW0mx/G5kiKkMeYWzrR0rpE/fhXMcIFGO+s8Z4ZIQ/OYGPmco1+7sXL3
wHGMGsMj1BHeWBK41emKH/c6BdDuFCQJUCVnh2FwUULtSyVk4ZO9wNfZk5/Kn19A
9k6Pob//lzK/VdVT2AWVABnx02tMwOZNz+B5O4p2oT8ct3kRWDDIx+N+Gywjcilw
rNQWLywkq/cNdI3rXQ4BnXEVF/rc/+WU0Tsq79O7lbE8CsAjvRNLcq9T2wK3BkS6
g1138EdWF3TIS3szd/KjyUqqUoFpuDt/Nl1jMFrihEv0Idt/h03CG3QE2CM4dx1v
SKWYctduwhwRbROj/0zYnLv8Spe3qZK2zAij7s64oQ9/s7gThjtmVqBlNZiCsd6F
Ov8m32EzN5Q37tIlTP342jChrW6GLJJ56zyy1rDWQBJH5EBPzJ1TAZugwlu/RLiJ
NZnsl2p/kxtCv9+5blfzxaNtmD8vjbePuis0vGsTFBazEPnyEmePCQlIZTPtvxF/
l//S8AdlBYb3MOW0jeLx1PE08mVxyQpICKJClHLM0T2Oz1YcuMreOFP9I7NHopA+
JHpAhNO8qebmk9ESOZU9hYULi5LyL9iO+ImySzdUnNkA68npsYXoMzk6qT0TRJQ8
C0M40bo1kEKDqhoJYeQqJ7lkzy4sPO9AHgm7RELse0gpVZvmiQ9yBVxCtsH4KcEs
vE+W6t5NlEVl59oJaoEhKM/SARPWV0G1M3zwIIeHNZO+8m3yiMC+boYG581F+8W1
oNfCUVnQD44KrYxZeGgPdXP3p+g0mcBWRxO45Z8zm3CSjb1j7SvybUT4FcbHvpcL
K/CDpeXtCG2gJDUwmx8h3r7oiqNh5+EgHwsVjBL/U6MREIj90An3snB4y5aPwjEl
YbpdAgUH3oklHBpsLAG1OQ26s9pzJP1WgHGSTm45jGWZHpI8t/2t4xnAUlRaaHn1
q6zyKo4R67UlHQughQJeJTew6Wi0XyhGTsT7QXoGlUOWIjImwHpNnEEpvIAgMNs1
GP3bmrdZPVX+ZUz++FfgCK+JFS1bPHPOGaicBsly167W/XvqMgyEBqbhp26F0UNx
BfTHq3Wfu9WJvwjt7g9GoAm7oCB/PcyyUJ+rEL1OqfyyEgCWl3mcp0W/qn+v7ZGq
ZHINyApR34fGRcwbHC89aaCayKzAP0+Ih1T+C0yvrgLWCx7EaV5fyTPRS/bPbm61
Ex3TI38nJSfhyOnAFW6YlvugA2mNm6XTYt0E4WdI7aRJB9HOm4EyQn59gYyngjcm
zNYARgJNbR3semO5Mox5vTAvl+mdD7JaI4I/QVMDUpOmB1w8TaEUJ8498QRAcowN
8qPJuFu+fgjA7QbLm/Ma0hPecLts+andlQaROGWwbXntHwdkMfeDcBrc6hBQ2Xow
XnexZL6nJhmu8DeXlnqk2sc2eWF8FHdgRNDPCDcEfmRsnpLM24vUlvKqiwxuNEgL
hVLVIfozgIPldETwvEdsvUEtkOFyBIDG151SjUHZ6UJyMXCymVKEinmrsBdWmc6n
XrlswyVtJMvccGUAeE6PaunRIUggYbq8h/2bXYDJImZEQuwWN8r6PlZ4ioyUrnM9
l6izbS8tKv1aW5tS1xtZMNAPJgOU0bidXBg6Lg6Svdqcf/Q7lFQl0HhwsmZpfmMJ
FQhA3H7u3PYWneS31AmSIKRoggX4LTdgWSCKh/hpOG+IDHEmGaR2nkGYTv3Jqb9x
8+4VW5BBab+TQJRE5bXGAGQxW7MRctOpb5F7/+UzWd7uI4HRmwwOLDxcwBFDtYf3
eyEPKU/dEdiz1xDYuJWH4BGAe7Pu0S7hp927Wv2Q0UPWmxwTeuxvA23CbL9YvIE8
F4JiOpXT1jPRbCLZQ2wvgYIE8X6Eh3O4TQKchupuz0uqlvUWnjIoBbRMSXJCQM5X
MpAx7VzqWp4MFVPAxBJAHuHxywkgK69dgyWV3zjYsc9IbAiiaUINbIVzssLOAU+d
mtdbKEyqSlRAhceqJADmd07a7hK7AfLAzHfeAPT2oHV6zYs4GxFE5Rs0EROi8taB
k9rWRgKIvCe8d/ymFrGoMHbanDXLZIQDhvkK2TIGYTgYCy3ddmv833F2ll+CHpI4
vRnnmYQAuYFGpxTFEZ0u6tmoiDv0ieK+XECPu7Nqxn3PLnff4vRArUZDIMiwpNYz
jl8rrt9PsQg66cnuaP6zDVj4GHwpjGGHg3Fhx39OJylx+TxRADjYSQLOJIUKoSX6
2nntsdCMuwCiG80pzb3aAQuBkx1l49SMrT/2cpKQtRQZuIVAbWRuyjR3RynPYRIr
TAWHGdEchaZSLlRrye3g6zp4KDFeg+oZydhIk7IeiCJLSqyarivpFVWLph2pPtvQ
uWH5GnlSK8xlhca+Ia0Racxg8LmBB8xPT1vsR5pK2OWRuQMFEF2TbaJX+Ab//A+f
+SHqCCIMRpuatfdlxnugC+4aoiHM50dTFdCAx9r/82UcvvNkLfpaBuweH4uV+plS
SQ7I4czXDNh/1Sd5qkkWXlD/QePOaa7aHX3qwE12vJSBBnDp9RnoGJscNYrbntRa
JkJD3DtDtf5UNdOWzr/6LdYYn5+BuNoe4nbPcEFC3gwZtpT3E5w26ijfz4lTJPbT
PLrwuaKzX9IG52WJy5VUotCZHNNNVwu5u5Oi1sRLHARB2DiJ8qhU/BShf2jGAuHM
25xFWm6qudl3ZhlJvqnNVHnfO/I/6FPLCErOgG5iijxhZaINpIvpW0Ov870Q5DuW
fGPIJrC00oEG41NiShwIvon0ecwjsuzuwoirQhWaXunQfNAvlq6JGt1CpcK6zpdE
wTfE35CEIO4wGKWXBT+nnSWxRzKUdrmzL4pmOer9oNC4Pd+XUIAuuPcczoHLDbXm
v5E8KHj4xBYoZpQZY8S/d7eg3ucKHthgaTMWY9vBBlnTxYjIKd2zYx3FGDzoCSoR
2pjjufD6RujPoaGrrfuU9S1mhf2Wowby8m99l6cs1VxM+jAGIzgkVcK0AWjUYH4U
2hmkf3aSNEhzZEGrPo2REWucxbaGMLgP6GygijBKRdZRx3C7heXVSYpNk5BO9shF
0YXVCFvBiFqTxrbSa0LEriE2zJLf8toRztsXtknrUGwq9Y5yfkf0veOKXK8TPnZ7
qkSJkZ07Fa5qtDMqaN48fN6g4wafmW5ywTvBnDnFUdqxmWOcYCpDPLFrj0LG0dcF
WvX5aCYSwwE8UdLRAB+8CiWPwRDNDe6T2b4CIslRDPoyEzPxTZFvccISuRoY4C/B
keKK6xI++xNwFehRBcs+pbaimXRomynono39OOtRHUdqg6Gh6Z5yLj+gFTeTrTjK
GaauC8GmLINc8/8U8TmWDUMtynWDepTdxeCNN8XjqtS8J2o8yLmBFA/ADhJ1tRBO
ofW75nvXyeSf57SpJvyqYNuilC5uHiXjIp7MWnjGO9MrucChgRPFisHMnanmRnD6
APpnfYQSLGEp+u/qxEqIfcw2znXmxWqPUFKtLelu7+ZcfT8WqkngJQoUBxuD4Z+q
30NpsXS8QlyirEMZGKrZ+rgFm3GXXd85vI/Z/5jJ3et2nIgOGlnUVR1E/PmHkX+u
4d9oq63asihptoQy6wr34vB0PySfW+KaJBNpvhZzfmXWf1/SNu70xCKLYQfBI2pQ
Txfzv0YprU/rqhL8nOcJWT/G3RfBVnMdsPKYpwAq+T5CX7Z2Rsm9IlJuU4805z53
QVNSeyvXCjogeQw1Ms9SZkI6h9JB4FxBRg4ufeOwzuZnXH8o2sHQtCo3krnZxgFX
ttWPuu2o8q3p7PQxTOR3yTrA+IC00iIYpJVSMPlC3UM29bfY3nL/0cnuERA+BY3N
6W/MLCTUp6wT5F8qh7ELYreUbkr1AUHsLMXywm4BK7T577vw3I6quPAASGhChNsl
KuYEdFzRguwh7qNnOf7jK5+4Ls9PF1LHFSTFFaLkBTg2Sc3wkld5bn43kaKUKezj
24kbqEnRp3N2f0e9chMzra77nhUgDpfOorc51it/uQr3n08wCibZFQX23uGkgONo
Sq0qsVvy4laHRq81c85mTLCuo8/I0x8Sh0Ski6X4txh2fFCiSo/k0WTHzsFv560B
rWyfn3J/Kf9PlVwzjegNSbB92tzMAIODHZwGQNMUS85QxFUQT5q5/vtPiqANYW2u
EQJeuQOM+Mpaii6L7fqac0Lu1MmaAfhaVK0Ya5HuVh9COALehdhSMZb+zjiXyXvm
+i6s/JuTFczbjv2JuVu/MLYervlU58O7ej/o/EGQOQCiLr8KZRok8XtWkzq9szw7
+dC2enbKNBqyAifP7igPeb/PQYH836zZ1Xo2h6ccGs3QQ0YFnlWYYPxl8GW7xkqs
Tmc7kj5dQM/Yq9wVkeNeBDxp4LiwkZwz/1htJDo+nvpqCrVkMuNe0tb6ug62uG1Z
7ude+ovoAcmxc/5FWMomF6FoIUdZsZBdor7gFD88SxYm4wtbR/tVRepP0QIRnZMG
G+Q0YjeOmOc6nzst7P7/0tVnYuHJCG6/0QYhuIvO0IL74hFf/MGjriQzamvFxsnM
6yOJTrK0PVP+xeqZG9YWqZHi5NUnAu4SJwEALJgWr0ns+pXx65CWxJQhY1sVPZB9
mO4V5RBGwSuHX9ni1SwhmSuaoj3d/6lGsJtpfWtbv81avlE/NXbbD5HLL2YYFd7t
4njaYzZgt/jhukPOCaHadmoAhFzS0X+C1mB0H6M/WFve+jZ2qVIcwleok7X48Zd+
BOw+3qPn5D/thqcRQOgSNCFMh35Sh9roFk40+2cCiTflTA8bnhNqZ9aMoeLvyZh/
D3FhFeggwqPoS2w6V3QkZH9ouFiC5vYaVnxa6IO0vxoDSzFbkb6EOH7A3t7Zns4u
RKtzt1NdfSuhPlhgbdLWAXPYvcBz0FyvfpV/xIqYDHchfYmdG4jECyTtMx28AzuN
gPvuu/4Jms86DgC6DWF4vB+4r0i+t76R2hj1YYJStosBGACZ055kpbBimtrevh6d
NaZZ9UPXFe2D+bbXd0Sp8nFzgSQ0BwCJafUMFrm/Un/eMtA2a2zSJek3F1nul8ry
q8sIuJLKBoxY/Mj+KEFeKTKttGRAsq9Ooc09V27h/n+vcq8oq2SfVsFWM/fyowaH
LmKm757f7GA9TcgNdssilFO+1Fu3dG97jzHaZNnPXJ1u5XajsvWjyWwBGTLh9Sc2
y6kHuM6gte4YG/vVB8VQLE7hL9hY8n7FrceFIQM2USQuQNztxHFvIUlqA8NoCpC2
mfkbtisZWpUXK1htpmEf1piHc7+oKuyb78/yhEJufU9YOKiLeCPMBtzy186Rr5UM
8M712oESwbw8R4ipheL1SvYoirEDYvviOFBd+bCudHzndqPSSiXUUddmNki4Yoy0
Ve1x7uTRNiAVJ6KFsIpsFlU66oUn+zKNTx+Ee3bXsBuPLeyRsrX1xgOBgi0u0PEA
NMj9vr3q3MmT9MNyd+uf3NjPhOA2bMejQpItf1J6FYdBnEIsohrqni3MiR3Q4n6n
Xvk27HmJlY4h1eg0y0DjnIQN8UcfUsjGwNanzfe2D5ULExodt1gdvvWYZJdmYFfy
rN8cxS1jNQafvXfbtIpDSvXg2w+a4koI60FV+dfdbdyfKbEroqHs2I3eeWhXoCvB
gEGVJfNZTqecuXyAf4z/L7qZhTd0Lg/aoUYr+PNTVI7fd9T5dod+h/l+hSqtYUrD
q/SMQbRCqvti5kZ8aL+15OSPq+lXoirJMA+qte/qEz7TimseucCrY0uQPPQkf+fi
pSTJi8cEhZHCLF/iBjtx7sd2KYnlXIuxZWIoRRun4y4SOGVxePazKKPtbIM/cdaK
dxLp+ZnRCO2e1AERi2/xl4rcCkv+umf8vwS+G2lySULwTYm/VrMA/pzelYuaym8e
jXPlP+MEavUI6qXfeTJAzMX/8MBmXKD/5pmNCxhQvbXaz6TL4nSU0qRyzytvhQ/Z
UuHNeiBSSCvOi7C62Tpj/ldlRVR/CWEN/ZKJcNymEXbru0bXMmUTWzoS/cqfee2q
7bHpN70N44lImzTn84anxoGHBb+7mudZkmdxfVceCQxBpP1+/KB7d0GwJVwsac4Z
G6F7qy3bGtZCchRi06EafFHc60YDJ7pZPWzNvqZC5Dqz9k9ZwZpcy7R1EkliTqHR
0O6QpivWuopAaC2NrWNrVF8ShC8MCKWdV+o7kMbPLrCV4A/SqmmIlx3yYgF4cEaJ
2GiKE+gP1WKF1s4qB+S4oq5sKtNrawysviKALqF6KZYLpfGjvZFmFXR40El5S5eT
kYwbF54VQ0sKtFPxwrF4eM1oNCl4N+8frOOoAvgeuv6znhv6cIijhA0Ystqa9k6h
gxRpC+4eYjZSrWDmgwrFYj2ADXDXFAfiWqwpXHNz2iN+8kaZ99ZhgrwFC7Bi0ylT
uWO3Q8k26FhV3u9ln8hY20AbaxqqBhLvdkGBWtRcRpbkuT+bItQufhg9MtRWYCJa
seAkQi0szNutdeCG4uPngECw82fbYaUKBkWyiyH0XWJ3z8td3JSBrY4bDJg0BkMo
0njc++OUlZYUKi7jbq+doQE+oeI4sJmLFOKpZiSgbOzNHBQslP6D7ivwy+9ugbbb
FeIWR2TAJjqFRL84u2u9Z1dN8Fsk9zNyBGZrhvA+FDvX3KN7qw5h4w6bTNQUhtNg
umwS2GEcG5GIGr6ubPPxnarmfIwH60VIotzKvHWi/eNoEQeRPG7k72dTjxiEv7q7
QQplJKoAQJJQ2tZ6NkvjozSpyaaMPE9A5JHytPLSaDGM0gzf9hyKmNNLhBl3Ns4C
2WldpBCEvf7CHTly8DnvO9EmTcDfcMU64wyKTAfoRdy3Qw+2LGxWA14FAkqKLXfS
Mo95E3Q27niXk99m615LZcEUznmpGN6XZNln4fI40t8lGWSTKzXWIsnEWQZLRXA9
pCbR6CPsrleqXPI9qmKQSpsPZ1MUbhjgQAeOAxhTI4mo9PL+yY26n+kXlksg79A9
chxJNm3HCOmFoFqWzE0AcKnD4ljddcTYLlbbYt3eKD0nlPHdtHepFcvYtAQ6RXMV
vYjHrZqOf8/mnBiwuWhNoNY5zHwqlGBHgk5hB/h0fDsbPQIetRKfASZVZRHeRa1J
xG1i4BzKf+eRmt9/0XneksPdh7wEHdJrvBSjO3oA8JNokgOHZ9x6qvUWUE/DrTzA
mOJgMLOtlnhSHjWLEXI/It+ks1cPC46cNpjr45StNKbGDzDeIgooQbhLT9wy2g4j
owibenGPc5Al00xup1fPRO0Vw9EaH1Rpx3ZK2AWUKsEvOUmeoVMJdHsFFCmmDbfh
jf5VrjcvJXLjHG9zgITu3WqwkYt+l8UVm1NfjkHErF1swMHnCZDZ3zaCQ8YPP28y
l7tZtq16ut2Ck6/H/WWpYLtkjB/KWTOCScfM+9wgFH6igXKUuREwQbiRRC1+3HiY
c+7JtfCD1fTMdp2heT2DyIfsUs0miJAtAAMWq9UU6IC2ZzuI0OM2hCntEBeiH0HM
SiIcSVjy29h9/OXA6LIDsw+w4iQHi8I66lpA3q1G8tBVo10P0WG8CAzl0YlCedlX
De3pv3juOUjpcPC/C+mouQ17aYLEvqip6Ontj+DhtcITPr+CNG7TfmNrKPMUMDfb
1VAE22jeszEaMbDvzsODTJ468d+alUhyTkpBgJLRnDRj3pqA2/Ez2LXU5VLcWqyO
Y+AVYyfvdZpjVEJIZEyzzkeVRly37zYjAWnSRfOo6WbudM1t7+xQyZD0g1JD3izn
L2XgZJBJlwEKWwi+ZK8f2mHoSmO87penrFqMa8s4ZLWGcoR8DN9ISUyltPNyYbmN
0WB9rlpnW006/FmuPGFTiffXX3gwAoBmU9VvLKZ/w6bdDs5t+3dMTTS87rJGzkM8
uY9pCUR5UaCMqxjAcG1Lk208sF89WvO12yS83GPUnmB5BOOQyXABtnl4yCbco6cp
MAAj9PmpZBLnlsYv7OaklDXr0kV9clgflwpuZ2B7IVvi8S+3GrzXc3BairaxOe1a
jva7A2mitbiAWloGk5GT2q66dvMt+bDzHx2TStGc4l2irNxiFmUTMbAxBZPbYFgD
xoqq9O9mQoZ7wDPMfzjtfc2tIDQ37p6xZz/VYnROKLS9WsrSLrzcd7AjP1ovdSjt
mqrWdkHRg53X/lQ0BWXv9t/IwRaoAR5kuMtfNujGir+XPGvl5avGF/lPrv1xKxJy
FZSNrL9omIiQEtU1f/NL+VWaKPZZxCyYNuflZUGsI6NES5etUpPTu4LKe5lCXjmR
PWXgxgmNpHOU2Lem4ishBOZ/EJ0haPif2Andp5M2IsT5JQ2tcpXT9ofrbpkCM/iF
ZE+gSKGCOHZkHKnOLdwfzpeiM7P/1alyagnuoRz7GBqf7GnwMjHFyHPC5QGrHJo9
VWH81riaAlku3knzMfKuqKM40YWFg64R7IoB3jlW4kVEJxEBHfcxbTxx2GQ0zmqY
F4NJd+aNDZNEvZdwQcH/keiJe8YhKdviEiOUcamCOk1DcWnZvqQbrdYzEMmdlmnv
aIN/ifR2EGRIJ3xKaAZDs67/zimjFPjOjQQ1I+MxpqmsB0Hrvt2bXl7C5EhBDHnx
zJmvBAPNxJVGam0spemF6fTkCKTo3sJOVywpS1MgEPv7ycIt226E8zdPL1YOzfXf
JwsTiyiOfm0C0YUdM3H8QRzSYSZ4KO2fpstvBj4/kw8Pq6GvNHyIxpqhKwR/VbJI
/d4W0rQ9O4Zb/7nCYfVYhIukycFTrwqODl70cQIAowWIOVhruxMk4+obnk5Q5p3A
X2bSYlgA9AfnwbdyipxeZd9CuQbGzSptZqSI0anBApIiC7y4fLqoBzyEGAnFUr/J
OfaOsbC/sGH3Nwlx3C76LiGCuIARYeJsH79OLY5IZXiUOeTim8CVNuIRA0qUYh5O
ezq1iNS3ZfoI2VIUCFdaAgl6TXTwkipPzi96/Ed8rsrxRppSFYZ3cZyRbR/p4Jga
QETPhSnQxw6xB0EDDsj+njmva2e+pzupG/iHcexVdhPnjm5HMJYdhOXeYVqYkEXO
Y1CroHxutOdm6QrpSm5DDh4+zl7erkzDuQJGV9tsQmDPdKpcD3CsppRP1FfR7Tg5
8bmzun1YLw6sBkhn86ALrz9aSqpS38ZGmKSVCkdqBcARdjeimWzEpx80ZSEmRiXl
0IP9pJ0JKSWp9MZVAVUko0o2Ti27g0jXjxGjf6sOlF6IrjzcsXUT3Mr1pDwhZ1/5
fRQa8aesETyHApxuscC48p0BJNcdptTMjLeGDl6xcMjuOXzInNt79VGW6n6s+9KF
AZkwMv/BZLZacK1tt/fx1OguXSOQMJd7p095cLpA9Be/m9jVQn44bttS1uFWaW3n
O3UH9QI98TZ0yElwgES+3rfBqHvzIu//smNKZj33T1rmQZY932wg+7KS7t/onwcY
hPrCq9Fp2SRFjjYwvKItwvS7so9Y+N9ZroMnDGhVJJwbVhH22IRwg9c1C9//ni7z
q1w4upICZ4jOJWTP0qhH+yKG3qoMM8KIZQPVK964CxZR/7t5iNr+JUR/IQi3L92z
Pdu/68oTyYAAhFUMh+cmtqSCuQtOhJi8DjfX9npu5oruIoucQjFL38jjIruA+UXP
MelnnC0k5o2D86AbZ3etkr2hWmQ952chDGvm2W72mSMQvrZWSf13WQ96/DnIPPAK
jZspeQKbPuA3GEwTB2AIRDQI2jVuU1Y+ep1qp9EVCjFSby0/p2B9nuJpcGV5SC5k
vaK6lHG5Dp1WbSjUztzQsxa/ZH82BrRk3Zu0Mnd2oW4iL56qZLNwxWvLFDYiRT7N
Gj5D1JBojJP3BJ5QrTPzrGlAAFI+b5WPjys3zFa4pNlnoXjAEBEj9dClFdeFSicY
mDrBmxhVllpiQ1S9tc5QwP7oLrxXBOxZ32bUw1Oggb29nNQqoV8eVsOlaJhbz1y5
SrTaVCgSQVdTWM1mbQFbP8rlYjQ6lBYTgVdBTcVeB/hZCX2zAP94aC8PC3HDMumL
CDju0whzCuQubl65Xb7/w6LnjxULh7oP/7+ikgMJxRJYvy8my5GhM8sYpnskO5ln
oG2GolaSB864SdU61uxvzMualDNjCrPWCp83qbsefNbBQ4SQn0b7o6cIV9K4+seY
LvhBoeUKR8DBIBx1JcFMDapImRHof8QQIRxfihySoDH2X5y60NwCla2ip8q7fFbk
04/UjTMti7RyWJNwYVvuHlkL5MPXabW2Ny6bW+2DCWxB80Si4umYrjR84I0fnBCe
Rv59xhfKl1L+UOeW4/jDXjSfcouFONxu3iw9UyEa0aZrHOPcnSLxX83H4Pl8B2x7
/WUDxSKUQPPSdP3E0A4nCLP6kZqvs7gAQMkWdw7Vfbs8g0C+0lT1BiG63DUk38H+
KmJzjNDSLqWyQvhZyTELIyYI0CIOcIYplQWVbsKfvdRzH9lA1b2ojpjI4fOtqGy9
zjPKwghiOS7A5niXAok20aZTPH523oK7ooZsZ/8uTlnNUgNlROOkul1cTPEW601V
ols4E+FDoejWURhuQBTg0JWh5pbOO7MlCDjMe63aL+eCqfWCfchmhWcFAhv8uCnI
HGx9qfttMLpntX9em7NPZJHDtVgcRqSvZMD+Gf3aVmdCvxOrLtemx9v09tg+1Doy
y2RrMmSgxibGRt9rHS2KcQH6ImL+rV0iN7wZDE1FHEWemGLP0eW0IeZ9GS4hJzpK
XD87T0MNHhFNTDHq+9Bo3F925iQhS5rNlPdELB1XhDXfAqQntGYqeUxrTG/xpqpv
blkfpAjKw9p5JbRNh4Zn8gkZBlqs7uyEudJXB3Hh8r/kDMZaneSp84XvQwOZckGI
r9bJQxOndO2i/sqKCIcjnpBENRFJta37pTXA9foGU8eZNTsgNe9Ln77hk55UQIiI
m0aQEYvED3OjCQ1KfqeLEHDHr+GZpDPQrsKwoOel8hhiYJYCSigWNDuOTziYv5it
uyk13X3M7SZ7Y7UW7UriM5O8s1MtiqCXx0dnNsfnnU/5nTSQ755BpIWzZfKkyEop
UknLkZUxcHbZLqsyAZlwKef3ji1xRRPyWzRFUvrJ+i+2j1deOinPGds+k2FOoZ40
Ilvf+C2EGzZNyxGDgbxCBlc6UOHKn+E37DZj75CgYZE2Km1gg20tUpVoEGw+Vk/P
IjF3FHenFvqnV4hnARdvs59g13BarEkmNvRcuYuCLRGmjC/RrEejC+q2EgctMVj9
FYIC2NDHoXCHHYnWGLm763I8FN/igl+ZZ+F93ZDaXl2psa4Idx64KGkTQ+xJIakX
F7jyCR2z10IHmVa6ShNo+JidZJFFlWzw7w99eFiFx0/SoyQ+Gj/Imd44HldV1QXY
GKT2P6cE6l+KEpAKq9mNSie63Jevy3LGZufwyRIzfE1KBsORrVjfKy12TPcXo7GV
bL2COwQX/SjjUNxmrKZHOeYAOVuljN2A3dx9zdd83knTID67rxs/Lra87egiYXQX
u71/wP3rFVLni7AcW7QZIloFXG0SR8VdvZ8AVgf0mjyVPylo6zPdYmaFADJCi+UW
+efMezrboaeTyrJAc7vI15HX6jJ7rAd1tbnhx6QDICr+vH7mzfNY6KMINcE0j0zO
Xg4B8UqFLydLA6lblMeECapnlqTB8D+9Xl8SQW212eaW5Zre1GxnRoJlsqxt6Hsq
bqtynmTm0m47JvO068fc422LzPrlmD5rV006x+kTxtJyL94LHXRaIfx5H5g4PZzr
/ebaixTiHJrIvKmn53KH13cJbdnML/l07aLnyTB1W4m8ZvjGuKvAl0iECbdDoEoA
vflS3rxG9CP0o5Y7gTo2ENTPUYeaSjqq4Ag3ctAMGyzjY+VbMMcoKWy6KJv0v0p0
5JEz0WDJVVviNspHwCDNs/i8Xo8VxVE+LUmDOGanFZjzGGzFMYap6Il0Nfy8zCnj
F95at9s3VD5e5bKS5eJnYJDAX9a02PjVXMTWM/LSWkYgxGbYW7OJjTumnUHfrPn8
NsmY1cn5GC+KIxFfd9aPbTeWMtn9GT64jn46/GecHrP4sybOpdgKREpTwr8YjA+p
E4SHXu8EjLNTNvid51B3CmI4DwslCiCM3wjFCyXPKjdYAt+KuE0uDipGqGYbTTJN
v2i3JN0EfhHGHLaQEOkqQvv1xDZmRUiXqweY9kTR9ywLp1QOIxhYN2xW4TNFEB2+
oa7R2UgmN5BKPc+4I31XGPUKbd9c6KYPZiXwJe1bL2mtU4GqFAKGKZ8HGFEB4Pj4
HJo/8MqiR67z+OQMfES1sXHrti5/8qkxzCqSMR81PTOzxSriBMOFHvtgwW9dp5Ph
hW9FN1CjPAODVDpRXmbs5xgzSfdD+c01eede24bbOhQhYw/5AW7ygX7s0V/1bDMK
XNiPFAyNQrdcZjwB5M1LmZfxf5soL1cQXWRKq2CIq037r2MYroV8uuL23UlDdgId
CiPjlbMbLbQ+YQ0jDwfXzl32SrDcj6Lauux4FmF8fax/3sFrwZ6p5cl1Gu7OcS1v
WjD3gCeh3J8RjNXkBWaSra078IgEE2tcRpoBPAIXedyzHXBtRbX5ilS6xGNHX1Mz
gFRUBus+Gk+4buDEuD3CesAzrhbVn9sZmoFdh89GZzKj7Y5mroJWMat+dXf6Y56u
q/yg9o3HITyJRzOGnyaFct+v4ynr0CzRY6MGMzEpnZyz3e7r7DU2+uzxzaKJm+Kw
91uhvOb379+b6zrqSIc4ZwH7DzJeccHJyupV564EjGOHP52o4MrhIKS1oX9VU8/c
v9wX8luoDk00vY4mBstGfffHWOR1EoYsZOxkFfyC5+V4/FXndi9/kqcrmJXWyNF0
2R47sx6fOQ4Laqp9aVzQsKsL6ro9WKNPA0VjDB8XaEp5H3Ylt2YYYcVD9RM6DlTp
m0O1dnVO6PxlEA8M0r2+QMdSTr+MyMJ/AR0rZ1e/mMeHW2hCwjHiT0gXK4uND3i+
C+J63ZcjFDl2b0VsCyKMeczIz7tP8tNWsGDZ3DTaMnIPu1yeOxPxgKxXLvOHJRib
P6fcAxGqr9NTPJ1KTIy6n4EnckVLkli7B13UTlmuzokksQdLUvCxBaXQx5YLVaU5
uJBqqC5dTqqH9g4my2h4d3Hp+0pPSJUK6vnIIKWE8XhKLsEp6g2r5BkNb3PzuzE5
c0CNLvJAuReJrhZgIvRKsMHsDuY49frVEor77RxNK/jJODpBBhFdi9HipCnJaqs6
dUaqJS9/rNM/g6r7KBLVgVAI0dS7yMmTvobEVopzpoav6sOWFrkmmy6Ug8x6vyNc
7Pd6JCYIekLG7TK9i5AadG64ibTRm0DDch1aN0ObkMowxz9NNp2LQnZu2C8m4lUA
9CObAzpha/sdBK4uBAkDs2QyEr+VqrAlSdySyCKV8F4fU/9ZOQE/PUNV8u8zIWa9
0wzEsscot3NerU+tpCw3FvZJ73wmGy6oVWCoGnWAQVUewWOI+/cs0TCNLprrOT/M
xOzSODjpQ0JnLOFPuyTLlAWhzarVSWRPe2hnbPa4JNeFF/f+YOTr55ccllzIw6Ir
nceSpnEN+Appj/uAVlMZpWA+Wu/GYJYEgGMtinsCR704X3EBQBo7LSx9FeF7gyaH
L8RC/4HhdMDlxZz7qhiO9B5h3SbL4XcohquZqQCt4G/rEt8+y1TocRXTy6Ax+fCu
ZyPHgViQmTcPIPcICynkjkiLlynAS7rrJ7dlW/+REhn5Qf1xA7loq6WdLKMC4QZe
6o8ylvRYCaaR+Sya/6orIKeCwqmgyfuLDn3kYSj5CbwH3QaKdkbYZUzdBSZMsD/5
x3opB0o9inQEOulhU1alw/4BTIAG1rIR3viMWeGFrmsi7gBne5SlJ5ZaybHt3Aum
SKH5OWxfjZyJhL5QiQojE4BxXSZ892mugLFnLLHmwZLPKpxqWEMdwo7gI6Ldm/N+
ARrhcq7o4FaG2vd9UbO1J4/h25+83jOUV9wi7RcwbWLLrZAoq4f/5CWGptXDAKmt
3URbHUE50S1vy+XgV66eX+/5Q87MwsME1WAQo9K1+uiCBObLFZKC0UsmgPf3FzUi
8ObW5zEV5qA19FdC2O8PX2qdEQMsJ4nMAy8f/lCPrLySws1R7fgjI3DuVNUSOtb2
gxH1rHy1xM3I6vCjvtkDn9mO7lo1ZeIjDXAP/SBhCBPJa3gvhGVdOn9VyhH/+oCo
5aIRmlBJHUweQvaZsKOofJHoOgUJypNV1//CEuwKYux3WUoZNcaDY70ZdU0BoDFr
d1woPrfZZRfNE9qYQzBRQPrwZrAKGcriKKMvOuKQaTBt/P+S3G812y6ksdcWAsZS
SAN2NP6jmrgXoPbESkStLUhgthnOmiEO7f0xtELXv1VAqw21cs7hAWkBmeTNqCgQ
nj4J4gnflCjvVWy49fW3xg2djUyH3FFsLCDVGLK6afH0D89I4eK5a9zq8AOOUtLP
vqYGroIAf1hvVnl3hW7gJiip6LZe74QGiOESPKytwpafp18a4nIiJ3XeZg1MlVQo
2yYQJfT6tYCrJWbhkEJEboNSR31ZzfXTlzeSJZNQB687m0IhtclrwPVwFVUzs3sv
Wwreuwjhvpcx+AbLs8XzRJj2VQkc6K2lm0SQS+z+E8jutfkeU0094mIuc/9tXUDC
hn3R03LBCZPlE1IX+sW93AaHpAeG9uuw21bRnRQJDecRMDBRnNX6TRkcGgsNmoQq
lZRLfuuMNI+Oinv1XWx32445gd1eQyEgfc0/202wvfPQ6tHuQwDG14N1+B05V1vo
QdhPsbx4Bm8BqF/Gj9zbAg7xBtr15OGSL0/IXa8dU0+qcNboZMU1XrOkE87h2Yme
1ya+RoAg9W4oDztREK8SahpIVlnMuoII2TAG68aeMMDialQNVPQZjjy+pp51Z0mQ
ydRNtWL3QHFxYcxsd6bKBnskv77TkuE+GQqRz86G41sEv0vwBSqx/I6JppjBcmND
PELf0nX3dAkT4kYXEpjwkLFdCcXGHyuNcxmb7HNhNChLNRdqnH/FrZFWdc+We9ta
OXMS2C5w73ySKI4j/szFWZpkT3qezVkUjTjxJCzQ2PK/tZjktIo5j0uCuIJ/hxLE
mjW1x/M6Pd2Buyiu+ILba2ExjTWDR0LrPcHXzVIxabhGgDpy138A8xMzvhXw3wyi
dvkPcr4htbtgHBvlWriDKIJRIO/AXT+u0sbPhArElr7WbLPJoQDzJ1ICv1V6dXKv
jL3wyAcsFF35e3bMQdnbDSYpM7GcFxj1KcT3Z9Oy8AgsU1nuSWkTSc3sMNkDo5VS
GS58Zu9/fU6kchqnQlTD5wTnaHPyLZb/+Jp6j0rGTYnwF1BgtMnjhAz+uKJCN44O
5OqEGqLZy8h5l04t+lgUjQAC4avyDXI7cEWmF7I8o4zLymgFAt9ZCTP4DieqO324
4WxKa30W+XuRPPcbH4A7ATzWf54E7Nduq0T2sPfmr72C3gUYSF/Ug6xK5BRUA2zm
UzX0JsgmA4XmLt08lQ9UW0rH/fxBmxsvEKAKhHdP5qSPNgH/yuAU/V2NDWxQPcuZ
cwkwB2FW5bt+r/VEufwKiv5vUDzGlFZ2tDjXXCiD5Qq3RRGQud0p6u7wGOMfNYO1
hE/dfwA4xagtURTUunDCz6490QIMo0g9nyjdZ4UCl3BmEMI4NHPiccIT9uwOREOk
Wp30VK5DcZ5tX4On3vdWRAKKTjRAHNjehweJZTTWHp0dNQiEJH21kafmxS1vbA1a
+61aybHDGLmvQc90GN1u4XNZhQj5uKZfkDHK5qlWAPlTPdAW6J+RDoY6JJUW+n6T
PzrLro567pv1QNllmj9SJVKvWuz3hNAhIIdkzxO7te/kZp7Os5nxaJIedhdl0RlX
sPY2Z5xdCP8bAKDySLAC7N86Q8ty5/xTetEWHHKfCcWVTyYLqVDiU9u3QqmnITxl
qr8VP66Ec0j6CzNVXeqxKdPwqFvrTH09KqYJpTjEhhjcIx/0d72vUKuCF5izCJS+
+aeBaeWyWRH5kJ8jl5kFp2QWSynTigMuNlgv987k9TH9ARzJ0BDRM/whaRULH5df
XmSfc9BMxdph327BNuCBu5siH74ionU+otqXvRxNRSMWMOXHtBoSPP3TXv1QkoVL
6UXsBfZFUfCbvQnHYkJhvxJpkh6GAyTlP8SYA7BlfoQ62KJdVhtMuq8oqIeXWQc1
3UWuEyeKojfuIAWNKXB+QZxumknVFBrrbAR1jSB9zZy17zjmiWs04p2l3yIMThAt
xrL44OMSR2LqVy2xtUbm+Z5pqCzKLpJWihtg6kdkiv1+h4FlY8SCNUNZstUvxdwy
GJ3A4pSh5nZrq9MjHyPNBERbReOXtWTWVffFScRKhagpHG3JZ7keP6x5WfjP9w+1
DCS9y0MAh1R11jBbHQi347cg1evozj7nlLqyqByZzD/ij4Pj7zTaLxqy+7dJKxtN
D8q4nq9VUNVtCERl52m6Z770J9NUZNIZzln0I/NbNnaHIqmfChpfywfAmJNoshuI
5snGtziyjdZrKSPFN1l7ma0I3vCyaC8qDAzW/DLEPqFZRQ98KaQ0xfo8JZTfKG5L
clJyo105AeBnT4kbILOmf9sQUEU9iymEUziu9YYDrYk5JZBgXMtnKBHppAIatUAK
158mvlDDDEEVMfcTXaS8iC4XPTFdEqQ3nnXdJTqP/Wq72AdBhNQVkeeN1QbTefzb
72rhubZEaOjrepfbZqFoTvkTeHj0h4IcQuasrRGlRRgd3G+4XE6kXpmE/DqEM8yt
t9DWLX5XYdi9hNfIy8A7OyjqQoAM+4/zxskgTnTExqOUukxoqY7S9phvcQnLdJf1
pVvAbgFHSHW30kK+H3fJWqCh14i7XX7ii5eOpaXM7wensuUm5Yq1R4qdp7zkAoMo
D4MywUGH1qdIE7a4wWsU8cfEgeTLiGaLPzuxpFsMzif4JWit14G7jbQ82Ar2rZqU
72C8Zx1x3ui8NiCU+rKNxYtRzgUVCETNKynZ3BvWT1Qr7iz3bvrygTDITmQK7+B7
JOd1x1jOt6FCbhgZ19cXjdXoo4laEoiuEYA6afH/UIPdSBmRXRNcGG9P5RIQ4+am
7/u1bIbdFUwNFFAQ0Mf/4XUWcLjsv4BkXu2uk1/5Ob53AtrrajTZF4V1WKX5x7i3
+2k3H/Tg1tHL92QnpKwx38Ly7JE6l9BvFsnYMftUJj7x3sSIONlZfKGzqgsCsYKh
+4NGd/lauBB0TbNd22Cy3jpVKfvEpuC6/m3ppeOuLcS17g1wAR5Hja4Zix4Jla57
JttTsibDfKtOUNSLID6Bz9KH3+7wGXlDIyOPPpK94SaPMPq8D9rwxhhqD71TowxN
tKAHlUaiPn13Q2c+UEXfqWghed/Xv6JvZ3AV4FdVKkqHLA/RhvVSaa5noxGFKMAT
CppinWUgqwWIfz8jyVZKuVGPFCDOcvw3cgKAuqGIW8OBfjbhOKB0ZiBQ2JJVgLL+
aMEeNX3wv6c8chp5fyV/cQDaBXHTAAGqA09Aw+/TtjvTgIhANc/rhF62xtorGlqt
u8AVDu+oTVNpoGfpiOrVEzj0UD8P4o11XbdQuLbE+/9cOQkYrArAP6aYwM/spvFY
UY7VN3nIT5VDpd+EwPcjYscoB0yhrZ27I2A0RnvjmCLLWA0CeKy0bDKq5IALbMSZ
R5N3s5Wnd45tk5OSEQVXrQGRpiafVNuekvZgI6wR+if0WV3gV56pwkreluNTq8LX
B1xWt/dZJ3cUTFjNFFRfDtHF0+/mgYkMKoFhXtXCb0ca/77IxNDhoaVawcmFzepO
Jzn78jrPouc+X/LKGrghXmGGAHfKCdjQqoS8TVf+FU1q5BbXHkT1oN2cSH+WKXTW
S9WeiOjA3UBHU76L2Hu4suOEdDcpM7/QgAuiW14dV7ZcZN8zdPn9Fpkjin3kcjRl
bmGd6nBCvuMJhgA7JH0G7czqcjzoG5cA1rjkBgxFwHKO/6xArXhbAerFKzaDD6Tj
ZQDKydm3+AuF/j8xn8L+pWrwBWe93Ezzwy7dfNVrxepgkLezCH7vrW6QvrrjcPQN
+n+Fiigjmjpx76YTHwZgCIHGWLpMCBHvNYClr7tx6rps+S1VZaT0U5m5NK5e6ipe
raP4OJ+SFHdNJXW/s++hCLWdPCNgM2D0amCBlZvZm1QSdMxlQi4T+Dtv6NlW2cOx
ieG2V+WEI8LFMQm9kPnGJn+lxAkuTRMFAhacyFqbSxcWHHQfYghYn95nJrg/0zhm
6ho/nB10+Y6bkkxbz8lkfoMFeNAzAhqMURI6uYcx8gQWQhdLrsnp75j5Jfg0lWN3
x34o0rmzQWzGdTsBHMCAVznbz3nCUMt45Ab1JuPRVsZyE8FT7NOL02mIByICDKTl
X/BJrLd0Cf3fBEw2R9btPpaNkkoi6S020ofbcX2sdLeC7+LF8zKz4TJrLcNi2H2R
W7/aylqfUc7ocExIOR5p0xjkiew6Nh4Wj/vlDLENS5EwGwu6DAESAkw4SM3cC/ZC
hJ64vvOcZumvNKax11MFTXAXIRFlCn8Xs1GEp9K5wPPpnETfMhQHVbG3quVHWtUK
8LL+lSRk30XCk3vQqrFhYO2tPsCcr0TVCwP9rMOd0pCuwU8vm34EqbXK0lC7s02t
R2Cm2G0vPxRlNn60Z4hAmCu6Y0txGSU2QFY36kAIWGPifv2CV9k56Cpucq8o9gda
V++pIQClNDPwyu1qzp5tcjII+mcsphFQW5cJjQUIsERXouKjHbtATHMKit0VD/kY
ZX2lSoTffwbSL876hlD+cMojmRIY6WEwhyK7gYUc4Ka7fItbRXro1d8m6Qzkxz+4
/RL3ta1LJJ6/kh2fKCtjA5HTVaLrObDh9KEzD7aQU/1LlKyN7pUmHEjynN/jEViU
xwSZIEJizORuRqucB6L/Hk2csaB3duye+4sj+4WtOMljHNcGPpo6a604kjDb1uB6
D04xjibm4I9DBPpGAL0Y686N35RB1i1z6icApxhv1m6XeGZx3BzOBd0weZYX9HaL
c6Xwj6USUsBngeYk6YD4pcjiMkJuxvGqVeNc1l5xMRYyjtqwC+EG/gyMAhyEYyYT
PTtsGoTmkxKWz6JCriOzRTyLo7n8kB3AzBO0tF1iUig/QMSoMrdCjRVr71ahPNzh
0WyTMgCMiTBnX0Us3mbTkHTpwgakn+SzDScwKqlfcBDtsAkaikLtnVfpOsGIY8t6
oPJq+lEm5D9vGsM6IFKSWwtzwc89kj86nO5cHN5+Uedp9CghVCYCwY8YPV67WeBR
OHGvFwGoIhDOOWPwZdELx0CCaIvix9eofpnnKizDH4zm0JlWhFGy/UA3vXFpLPb0
hmQa5mi8UHvahSg6wRbT2Bya4+E73BYZfwDJ/3Z0uJubXeZ4xvGL21BV+gt3sUqV
MtZzM3zZJgh4K5YUuWgnJM4fSO4oqN6U3amgzD5fGePIScamlCv12EhzSuJ/HUq3
mI5NWQLjcMR9ZwP+WdPDMTSz3HGJbfqDNoHZXXDKJjXkYttVJ/KUbDpp50/jIedt
RgKc4CgEOAMYTYzJ/qDDrutiz1ls2M4ZYBJZ2VGqsi0YjxNZOGw8B8S7v/sO8820
Kusx37ndQ2D/x+MhIYNNYvrxSlZKo2RBPuulF74JWng9hMwyYfyJ0ssl1SAuqQfP
sJdqbpfghC/eLIKfkoWbiNPGlytHqef2IdfZJ5jh8fFCmDUrHbKQrRRhEuWH6jbT
obxLY5jy+Bc+pFKPpZQvHFJRFIwXTg6/YH5kbYxhNyMovmAdiOt3ggyVxg5v9Xb7
n7pU9GJuBYOTgWZWOw86zx9SpU68lGOMhEQoCSr3zyQEE2HMxiQh/01nX3MBw+Nt
+A3lg4NxYPAAfWv/NU36o3hMDR0lajBX+w/tQGZ30JEPMCh+ewEhnH/4NCMvSRG5
pBendbhTnVieQoWgTxyBX0O63n3N4zy0Cx1FDBqjiM72Os1WP0Gz2DkAYWyWjCdi
bpEYeR5uKv8KOzWf4lnFDoMwcU6eFax+TrtdhCLyxarOkDgcZ2gsDL7w1J3knaQk
Zh4pafdjH343XS/HCF+Jr/BCENJMBVydLlTiIFsWvFqPJ4xxgTrigdrWobO+grU5
8NpThNYCFRcB9+KUQzN66v9Zn50KKSFjtoLBVbfjzsgSZrFIhqskMssci+oIQF9E
A3KcajUmyYoAMwrmbhqnxbhhs0Kp777PbgnjFRjqjpoM72gGbII5tkQVhEtugfW2
ewQg2LP/0vsFvHNJR4COTk8btIzaprCIH8znLcpIjH1FYqBN8HVhX4lhLxBTCJGH
6M0uZsURl5QCIJ26F0QoYuybJ9yw9nhoBkU0ALdTvGLlG73xIrEvTDxj93njjLLG
fJhSjHVweSKikfNtBfNz+nYvWpgorxusLJ5/Jsq/pT/ixpU5z7BodJL94+6J8dRT
UIYq+i50rwzayt8dzXp2CHVlCWWu7sSDIuHjb5fJPH37iD3IX/am5KuLh146aXte
CjHKJ2aZGlZK5v8UpkTmYAnP5nGAvoaeCt8LBXEcCaEN4g36ObZWC8MxIQnv++2Z
NxCOgjW6ger/LcN7sdTBHLj4FpABNqAQi4iOakJbZZFgtx/+kusCxnn59P02/2G+
UO4y7V/cTOSDdu/9/RZATR5zvIZQwiq4dTsaZJiCf9Mj3tjVVEwN5TVd8EvMxsiq
0D6n9l0ZytFOqhMDWyIG+2/LXUsWxrJaoiA+2NgZEOn/JMyrKU4xTuztUZiilAAW
UrrpnyQwFzclkoULgUwHLp5erX99vXJGYVHgz0FOQS1HxV7QOQGR2f1+OSHy3nW3
S2jDfpYOlTuROL30ansC5sZ6bJwZEOTZiGhBcD7mZWqrM8Drjd7OnVe156EACgnw
dYodD1JCRzYNH8961YIHjNjARcJWb9N8vG6MpkXbqXc6TiP9JSyNTbdHHF+Hj5aP
f16lynsK2q570kRAcWruy2VeTwjeb/8r2KsZI+NgAJsAplpR+vhEJsj9Svcp7A3K
s+x4p0hbVtLES0hTobPrXDo0me26M2KF2z67Zh3jhJJaa6caAkwym5I2CWILMqhc
8RaCHptPIz+e9fs1KYKOzzMDT1LOoYXyqsCkiuYPPU/E4xszAWE4CdxSJolCQKcW
oZfmu1EGgb8TWKJHLXqk5iAjVpnmTTA5+WYbevbuckX1I+H9YJ6ut8TdXC298H2p
4O6y/yRgUMr3Q0tFpnAA2kPUD/x0KL1eLvp2d1OUZZT/2TCsLK1BESTaU+HhiuNl
SESh5Ezi+tPjuzsAb6PS7db8GZ29GXaLMW8tVJpxs7Gn+vTbTkxE5E2gfwzvbKjL
zj0jg+J5rHHVJTNLFg5e4FEMRxNDNmMLkd83Q1aTHnP4MOhuMx3i7Zreq6S8YS8T
o5d6bQ2ht65GVuh4CupFo+9kyovGjvIo6yud+7JNpDkDwcRva+jVKKbN6Ief0NBH
GZ9m2uGzdGwflxX7YfM6o8WfJUpOGqIatzoPPA4QdPDwIVVItmiezml+Ss5BtmKr
TXQP9J6TdzR8UJuZdTtJUwARdmrijfkdEvcxhCoJxlopJxT/+JVdeIZSV2hz6np7
d88Pvmxbq0E1UPwTSfO0CH+qAP8ClVLiNhNgS145ncibORaLiQlbVZJLvUzCkPkQ
1hzWkCHk3+XsHYFrl478pr7VukRb736UVB4djOgx8khEj4AYN17vZ7g02gnyMA3W
snmlrJEeIuWO3P4mKXaRcnPyGnZKfAtJ300GMjL8XRnvAx0z59onvVvQHn9fqpgX
NBJxHGTCuDxDHXQkX6z2IuMW4SyLMOOkuYKum0PYgrg3b+063fKp7Vjjx+EYGQce
VzU39ivSaLnZd6Abpu2olouyNCJJcaokFP3AgIASqKyasgOzgwgZuCZGROro9GW/
i12avkAZaEWKL/SnvTKyvHr3fvpfl2C67bowBeNm8qy2XaE1CTSETzghnAb3C1jQ
tuFc1q7MrWUyw5pomD4iO0iCDjp57xItHQHRAcfP4uUPzPYRna1d8UQOX2XE5LrY
HyahRWOsywX6etmKbFvXL7HbQ3YcUg/x+mgZfkDBDm9WDw6HLJWodptRJPleyvU5
0OxCo1/+A4Wn3d7sn+SoOELv8xNpXu2ai+5BOMQnjKUo6FJywsnsUvbo6hs77Ahu
3rZpWc74CZFkOY1mtDdTRosXlh63FHxrTx0PjAaKPM9Pum0HAEy6YkdsrewF4/cP
OiaLNQs5R5Zv8ewYBxz7JBjMR88Gc58OVLEbGGfmEAww5o8TiCmtCNRhnBkXDonr
g7C9ag223xvRqeH8Ob6/jEsR47j++5wqlzAtRwcI5rwK7oHYLue+cFoimt76fgAe
8zKBJK3CFtXAVx0V5BM/XEFl7XVT5c86UmHucVsYqn2cWCltvOIXVBs88wMfaLWt
S5HvwTTXESe1FK9Yecj5H8oldmDqj/B5kEBsdgy5OGZ2b4cQ4kEHH/Zn5S1mXw7D
KcOfJdSvyTIojvDWiHr9DyrQVPjGtNkxGtfyvhM2o4q/4guLcD4oZkTb043mWLJf
o3+iNMOdCkIvZyc6WIGlIHpOipJWGYK/MsvqmvzZOBb/0YtMq5g3Hd6i7BWJkOm2
8YMG4Pwv3X/KwQQb3WcksvGbJTPlc1M2bDjUhoPaOC8mR1YWIaBICAEFG8n97iIv
A+LkDb/2wF8sguS3Lu8HiZ0ioCt1sOz7aOZCCoJwvzBWoy5Gc5Fi/mNGPkevonOL
xmFj5RpMBqimGBY7tui2BldkiOFzWmt1m3TJ6PgMpQdnbcTnxvYdYQKbkcI7OeY3
sjCXfhUEQVfIPfjhFcWUZd0x9A5AMaNiu9xlv+EBgfD7uceHTJafj7bcOHUi/ZRP
nsk49A1urkiJUtYh0jcH2Pff+zxUQg2/egfZawHPzzlrwEMZhexmMxBLTKuAUuFb
PD4GGENj0Z+rWZ9dUhyAoIawdnZ/QA1ghQIne5BtJfwh+2hGsn12AhOr1GOwBeLA
gkVxB9qQ41Wr22jQgedrQh9z6oGHVICoQ4OX/5OoMhn+8PH02QFiNZhsngVWJY92
NUHsOGelWO7jev2/30KoK7UiY1+jGpvjD9jmIk3833dGxwh9AuO2ran8x4OB413x
L3+S2jmNwkz0e6jjOsvMrqGKwmI82V4wf5L8QAut+Lcv4x8ecbfvbWB8o2t4oltI
nWYTy+s8xOj3ic/77o7HLqI9lYZ83feoOBkDfj9oiE5GxdlfIkQSek50XfR5PAnE
E2RVyYWDyUKEY+qRqBnHEZJLoGvyVU+cvI7e4ZTHulr/4GpaxSQrHvuMI/azyhI5
ZB3EsRSDcy1Q/EPHCdwf3xthZKDyJkXfBJFKat3WAPLOsJ7wn7KLZQJHx8KDISL+
1Wx4AOmIbNwoeCTwxBXjhR8XXa5L7gNO02hBVFqchiTqAfNuEoAMScdqMXLfQ/Nt
SDevEC0Aargns54sbYwxdK9tsxDwxsZ10DmCaPQrH8nbfZI630p+A9MiOTtokrKR
XENhN6d/D9ce37rcdhR9xLKr3agUW/qedQQ749ZjxfpUGDouChA8/EfeECLrMI1S
A2tO5OGHWd0mBrTY7JtCkt6L74AhlMYlNpCeiqEmNNpV5h/mBCJUvEz8IPxN0BmJ
j1ai8jjBL6JRsYp5mrAnvyVv2TtDAZi+tbLBCPNQm7+W79VR2+B9/f6r1CqSC/pz
8YM5ULDxMATHPkHv9pAqWpqtz3VN1LdflTVajCixnfPPDLZVWHUZnBQhXRTg6RUg
EzhX/u8x4L79Azoke1E+2zo5Ea6oiyBnl1nwd4rESB63KYDMo9ux+2+IIJxJS25C
q7XiOof6NgXnQfbpuY4Ao3vSD4d6sog77ZEljkqWzulHFhQf7A+z2xvbdEeSftXn
YVDOEbBA1rvvfK9vUYI62qKcvKVhR2sTtcjRDICQvkYLKdYFHUkhtVYoDtXV2F6Q
eif57VCEnplh7mxPZcoeGZeJgf3vSieLbo4fFSpXXoWvvqEESoRehEWMIIi6Wyk8
Enm6HeOm7hRGewgkL9hm8PhAEy2tNpyp+0YGJr8yo/D1UUfbtvfXMJot92LQoBAv
kDMykg8qT7dMVFHxiXjeefbKo/C1v9O9q7th8meegtkT0sYuxN9/FgQKLmwiCiRa
oDg+bZqTE6y9jegUATXMOCJma75NkqYiCszT9hKEGzll45SFASY4zijcPcI+RSdX
qHh5Y7jwbiShC1xZ33QYw098VG3WmVmyB+6uk7Jr7NYKphh41P9mkt62YjZLG3Wt
WhLuI4VzIB/Lgh7NeOxfs3q5deiFNiLQk6+6cAWKFgiELWTvSHD8TV48Mb3sgrif
MIX9xsSEEbuAq8ZH/0P1KSRqoDOMtmFiDl6EAMpH99rO7SieBxBrQtIeMylK7uN2
9oC8keIYH/w49Wnht5fWr1o/4EBOzyHmCnH10R63i6A6m1gWVm/eOb1MGIlY96V3
vjrXr2o/YYfhIWl7NjZfKZGZEGGjAgSwbWNY5547+MK/dtTlqLhG9B2h1RFHMAXH
/M+iNKbwyo+em5XJ8D3IkIVYOzRzwiuDS8vd+jwEZA5P9bGdsYrCw5ZfrBn8huWA
mZAq+PxJsCloa7hk/eme7TnN5o5owUiS8TjXMvRpwwc5+3xULHUTCZ0XthD6AoKJ
rBAuRkw9CQkxGpWl6ah8UqJV3PqryGcn61uWrR3k4/xFC7yjLfzDtjaQHJ7D0Ae4
bLH1nZcRWLpWfzUa9Y9c/Brljr02JWEhfCJIZdyD7TCV/iFTnfPVBVR/CvS+IXeD
L9OQYnls2GnaiXV9ukZ/V5xblH8z/wNLrj1CcV742my11NGfBMSEKChuj3Okami3
aIl4ub3lzIDrJuwIw44UqjwpcBuHEAvBg8BEF9XfoBQi2CbIXNo/5tIMnnGJea5q
P7iBhLHe/thCxYiF2Sr7Kakd1rWIbsblCn/uzsZdIU8yorNMXjzcfmDbDX6kjGk8
zaLjWIaJZOenVLdWM1etmeKKf3xukC27UiERUpuI92HAjr6+6mZPoD6zDk/1RHrE
2WnQ7ZGHJqAQAB+HQPerIk1c9/pvd2/1paWJbpHGwp7SUQhQ4z3AO6Oq4X6YUdCY
6apxLnsXDeRz5WQPYggGQVVFjKTSC2xi+7HUL1FwNjUPjO4FhMYCfHFkoqraP+xW
XLM7od4UAGuzwJVCodOPvNZCukHTn7JUS6FsJPWRUWR2b68aZjZAAlrweCMJB94C
Ab1gFrlkzPfyeFSkags4cav+Wig8x0hVARa0SyhSbeZHly5Piz6zbG2q4WD4aC+y
HS/RZbCvwGoRcRhd9KCsApcaps8tE53x9/Mx8rwjZK/XMHbrQC0GRMU4RmBiXCSc
IgnI8uqcV/nr+S6UhnASHS5TKRWTgzBByptyu1TkOdyre1wzirzjpnob0s7TanzJ
WAwgiAS2BD9nkZ8xWZEgOkGcrkbrVFEhIafEiWDWosGdUbPmkuk8XeMDJidb0hsN
TkXQZMmRLlUyFfNV8Eogb5eCZLl/Ri4ftEsgnBUMuSfLYJQG/pkuT82DuPZRHG7Q
SmplMx/Rv7z5STAK+W4GoPa4t+v5+CYdi22oKl8/ViWAjBpvwugttBGhqW18g7ea
juN4EQ6nurJIQ+eDhVdQ9ZxJM5p0m83AZK5LCK5K1IqR/mD3xUdVQpiiA3+RjLd2
ptUno6klGn2l17O19GwlCfvy81gZ91Il3FGcSYfCyfG6wLBEZEQSQ26NdxKFulQb
LPK3NuANQkVW/um10Dlax9MGVl6nd2aFPPSjFocgDMt/ksiXaKBtiMLTaFkSvxS3
lWR+iifx9w2K+D0NDeB4wdUrBXcBhaZum9hfCYAM7PrsbzeRHtktTKATW62DPYPy
WwJ73YNNkfZa2dGD9uLC6w+emJm7/YJiwW8LQRCaqd70egRl5UGdpMNzp1Moc/hb
pGoxA70TAeaQxi7up2iH1JDNC+Rma5gcsH+ijWMT6+98DBRyxgXGmkZBAVZMkUWP
drJ8glVNud7HsV5uCM5LUHRMpdQAl41HiOl32/ZelR1vE4yNjg63rV5k9nVBJIs0
BrbidxXtD87fUO7MSxUkUHreA4xKVzdmzBhkAGD0yDHDB1C8SXXJDpt9Reqi/HUn
zKSKX/y30dVqg/WgriPovZEhYw1jjXBHBGw9PnkJKgB7IQdjv2NLWlYSk+Oae7Ow
RFIdpTakoIZrhX0COIuy8YWAygO8Dylir/zie/Wfkq5Y1uT3WOC6JgDL9jmbHH2H
7Nu9ax3SdHOIm++9KIpamTGwnFUPw0BeJLL6GpS9O/YgURFLB/MMy1hsLlDkuUAu
Ri+bcwt2l+2phmtlzGEhjKsNbG0ljMD7urw5PV9B6VAFTqV4SG8NUFCjPkHL1wU7
Pv8iGodz0aS6Xt4LyAhHFC2dcIOYuWGpLqH9eNNxIYfjr5NtiE+PT0tuokuEF9rC
Lt8jLWoLBjw5pQEwtpcWDaxcdoFZqFstzJto1F/CtnMioX+gQvoyCXnVPfk4r38X
0dc0+LkFMvEcAuQdZsdzylFTgMB5J/1HW0jnd8AyZYNnFqZIjmJYa/PMAtarp8Xv
GH+Y9/s5aj6WoEQDeQGlJex/QDvaTw/QVkyA20FSgX1DXIx6Tc2VZ+YP/vLdLrxO
o+kLhTjPp6J0XyM/3XQ9L05O3xtb+M/LegznNaImHuRYVAEIyLpKgeYzVYkjSWeA
QbS4tbGH2bypyYxvBRkZJg2087zwiLDGT2p5SFh6Rsq1+iQXWSUtSyIBzkLkrtN1
72BIxG6Lr4vJcCdo1KlnyGNFeXFWSfP6jUbvSicM60P2aWQXHP+ekAxFFqrIl80s
nhdEhd6VX+znUWuRsWbkXXRGfk+UK4CjxuVkYxC6EmgW3yURlB9qZMpQvntWJ+ON
Vx1MbzcbD2ggFCYa4+Xq6kbbgNlbfOpk8tkoV4me6NbGje3WyWg3em2/3SvOJhQO
J8MnQtCmkqcu+WQCt/+18u2WMQjSVZsFzj3H+r4gPOVVTWh4Gy2ahPNeU3N1Avcz
jxRV0DCjCL/pr3IJ+1aVmdCMMRcIsa0ERnmDxxz4awRfH1WVxjKXJu+lhZYEcDI9
Qm11PVMC8pzGB4YA2vhZJzVIhQMItlI97pv8YCluYeKjd6eNafVezVAbqxx8An6H
YfFnZvzeT3o3LjX6KbeuBm6PIGYUTuOuPvVsn6r8xjHjtaaLQ0kocNCsdY1mcR5o
i5oE3TCaVUI7msLwED1U02919KQ/f4eQcD5utDZpPV8MaTrAFByNiMC3KOCnph56
4Ro1OSthUhf3zQ3EnWN4qxHUfMEwWbBADfwdDbH11ZgYDEXayF6C82hIQKWCiqRU
+3j1NTJwK7ntsoStq1fnaTTX43grWzSKrX7n9h/s/6AzJjWvFIwnki9Pt83YUDns
c5NnoeGbREYtXb7jQ+xvd2N0qf3uoD3cI/Iqla1RDsOu9eaAj8sFHdGIHg8VjPGk
b5w7nzGdaIPbrYcTA6NTtko++51Xc8a1rSSOxcKthBVliZwa1eoniKcc9Asewb1q
GeWJbnsZ6TUi1nqm4SftLsb0NRhLsaJ1O0O/a6UgcR6foBeVmtKOmIFFWCW9SSou
GxaSFwQuqrcs8YfRUKWNnyfvlPEjGUwmRCA71XyBlQht1LFFn8bfNrGCwuuuakcT
h8cS1hKJ9bmVDFyycCrOWUCv5MnUEXn8kNvRGKSBkCzUG4msqghcJAKyuUdvTzQR
Wlzb1yYB/dvuen86epEh/eRL4lTe3CXyBZn888DREUiX06nH8nyaU5njrtRvB2F6
idoetoxsN9Fv6G//wyFEoWCG7pbnm2PwPmA9GVDP540VXUKdZyNTHMvA4RJtxS9Q
a+0QN/Dx1ue/mymJIcs0efp4t1ZbnDpALi6ckqb5VqQ2GOTjfNRXrE/QltsOMHb4
xNLPQXr5zaJLnLT4PRDH0ELCf9ppL2fY4fLQHdLP3DvnVpvj7E4gsv6m/Mgja7SL
5AGWxpGbEveyNVIBgjadD0YqWEHcLh1MxFtq3X2598KBd8QXosDMr1oQU8R/myTH
eVU18HKsTPZoFPtXZgW69BCO5rBxuDv/Qq0IYkehilZfmMfn/QP/85EDwINJDhXn
RGubYmLQ/gOEGfy4xhJscDP061q5+thYNtdSkrA61wrGxdmZcd+dbS7PSxYi22UG
SifI1zX20Ss6m6rKEn/W9OFwFAdPbUhcTzg+xYf0kXuFa8vVAJRjbHoaWelTFxUa
rw7lRYsimnpcMCuqhiRo32Xywepz5Hh1XyOxpeLPfq1VGmaFE7Z4pE9bxJTi6abt
F9lAdqcI9HBf7aSIzlmBiYbkJigte6Mw1xmXSxdkCizH4EXtNKyxy2bJZXDlThwP
Vr7RArq7XiSaoOCObdeG8H/dXQWPpq7x73554ggiMH8xP+t2KqkmrNTRWevNepTq
rWbdd31YYN759IGsXECmCKaa+Jx0EPYQNxW3X3DHGZDMgg7J7f0FTaPlaL7CUsC8
0mIjCnIYfNCQ0KXo0DgVITFJB+oSx8Z0E33829K6/73NfEE4xo1wMDuZqJEfaoZ3
XdN5biyu/70zriouMqUaP7S4XggkjD4lJTLOEHHgOA2gmJ56Es6NLo94q4qbcA59
FAHn8PUBI9smrNppoxjr248Q3jI9lNWilWyNtBhHDb78jiPYeO36lXbgAJPrF5cq
Ee0pAkuNlY+6BNGdWajZZ24f/XKTC4WyjmxhNhP0o3VUfYXSSj3F9FUfwC26gaZ6
k08zc+JcYC/CbvosyM8GRpVXr8REpV6MJ3OV9joNK317fxL/jF2Qd0Yp+gdfPAve
f+w73nzoBkNxjQ8uouWOmb0gJUWCtmFC5hKbsfWhhriNC7Iy3q5PJ8+RSJyKADMi
z+tv7tfk/pEMhq0/8SUeo/SnMa3yyakM4MT9AWCfIVpLAZuYwBZaezo+OOz6XVtg
NsPZk7VdWJ+XA1boxNDdXuiay1kIu5IqQbqso4yxGMyRtco2k7oSWF55UkxwLkU2
DNSsWnetCEeSqPA1qA33I9cn4+FKNtBje+EELonKsqu/bVXQU+7SerM7MarUov75
P87Zf4n4nrL3NGlGy7MrDr9qpGcgSPGLGRn5w4AxxlBgZF0H7NdTgQ6uxeael/kG
9jVTqxhBs75nzmTARg7luCrYQa5SN0fYlbHhIKGiUEaXgGtDwClk3QnvZ5dnYHi2
ircFQ1lIs2vNBUsK2nzPX/6PoMe4RE76VgaAIn6/JgUcKeVg6Of7jjDUQEFxyfF8
/RSCU17chJ9kijovfrhCTIrsROQ3Sc2xAkvbDQebEbbGnx/fhvphSueaQTtwfkls
Uezceb5++dHQzJY3zl8WrNljn1GpSwwEyPU/61qIBYLn4nxNGpA1so5dLCT+EGxS
MpXGgpYYowJ3KWQwTPFQs+EsdE8fdFoQ9I9/nNwrqd3wsLKj4Ew77PNZ5ZSwgNsn
EsKuzCAEuKTI8MG0c8de/SZqcLPiXB5tPM2M1xLOfeoXJ9DM8CincCjRf4o+jBgK
pb9/sOsvgfEivyq0EiMLh9qukJElnpLZfb/0/w7Y9rqmf0gEXAEd6Luis4SQI83r
M3kWgC0Jye7uvLr4b91es9enR2vHAy0fpJB+dgXv8kNDpaLzLU3lXnmYFjTUEGWd
FVv/ziIiJRTsvjFFIP4XkeLiK/NWH8w7em/DsiJkBN0Jjw8q/Hm6k54ExyG7GCgu
Ss9Ixui2h1AU8k4gL84oEZYCivm1wTTt3N+HYglF5/G6tBWu6+i8bep5KSG0QnqY
3fuRkbCW9lnmSxiq8WaRLNhIg1XFXF8vadpMp58KRALMCii8/WvTEGVsa5Ud4z9N
0nWHqWxGx22uD+qoEw6vuT8YEhOAhbbjPZQ0LoVfhFSOWugHDcZvYPZe6FCme3lC
MzeDvnQmI4iEhO5Fq71j7Gyhu2Is/H7yP2hRJBZaJMAsdI6R5F0DOhe9RykgdN5t
2cmI6c2b5KmB/J6s81n5/5gVqWfFxGTwXZxEYig75uU+T1xw/JvSmpnVKvb1M0h0
BbVdb7wXrTUT5vHi+jGUEht/c+hn00S4G4PnOs6x0sallMSMUK1X8qGBOLsFzQ4K
o26HEaLTkCkvKLALnOYR2EW+Q8Xyk3icd41pkGxI1wFxvxxApLgabHfDt39oSP5j
ELRXQALlJufsCCN7U07Fb6hunkOyNKZoPtnWMvd2mVG0F6kHsg51P7tmFrgeRAJL
WjjMq8hRMarmwQGnXHBkv0gLtJXGslp5pPxJVNP7Yr8cYV3CWPJpNEKgs0oiJsz0
vD/NQAzoqRh/GHwgaIKC1eRp6IiPpTHwXbcVyB3Vo4fXC2tFDjCk7BUekDI3VMff
InSlgJ5A2NPMSkl7wXPTrcjUX1oiW8GpH37Pwx1yHWFezwMYTZbDFEBG/KVl7C3o
BZ2G0Ew1UnKAj4HNbpFgZxi5Ce0jrLFI57KTawQ9289CGhzvmg+RVLHLfCF3AKiz
yM4lI36BDnYIEL2wKyqc5QjLrZ89/qM9DRJDYQXizMJsiSVnQ/y281Go30qCqCb0
QenWxnqBUrUeEBjUpbNopgXQgFdjh0Z4PNCuAInTepnEMNNQPFWXArlVAgIs9HJ7
b3YyluIJzjdfpaers/kalfzQJXIW0v0ZborvNuzyp+QYKDBK23/Ri6V6+ptJj+wf
2PhfnvA1Q0roRag8vKRboMLnDiFUDxa9KDSpLbETH/u3FHKFEWCBayrQSeWM8sq/
lH6zNZulamZxp6hCL38XRl24VWiq2En0rCH74AwYV6hGMDlRMhaBij1QecOL9jXI
QB2UICBKquZRJRfz1Lu/rSo3OxBh+MS7KMS3Cbhh/AQ4AD/4hftAY3R2ONqPkMAE
JlQqU7fGr2V39cRKYJoMKpdx3xa6ZoNaogSJAXA2DNVLe7Ed1+4lVAxTI9Z9ODsL
6VyxJLfSd6E5wHDOUmydcGelXTQvoL9ZJtNn5cw0qb0ZErpv38kp+IurOXSNxQD0
7zryjZxIOIVvNQtuh8Xcd5psQkkAR/k7b3c8IUDQ0oOdtviQn8P801R8kWBmQAjT
OF4bADuGJA9i7b5rzaBLePr0+QzSOx84kGsJ2Cw07fffjRLAEczG6FbXuhbhY+HO
QPjvZKBn7pbVensuQ9V0NpgArrkWNiW53+Yv5cgdScmnZSRBJxnpHFY6RTLdQuhU
6cEleIeNJJJzANMe+VWHY4GJD6FWp7oe3gMzniBlWx3RaxHcuo1kiYY6ntKTSVWg
or2E8QKhz1ddtlF/HQi49AH5/6p51imbiMVrHebvUpBujYTr6JUmZ53wGmx4Z8ET
bOycvi2XGMkYaWoiGEb1M0WG1N34taGcERxvevyWJklIJvwR4EQqNCjqIiElZmgi
zIxvCUvNQ9vTeFw3r/xwnApUtgqp4E2w0xuqqPUAFzSc+N9UXXlP13Gwr0XpKUfh
D/bBNxXs5JEv0TCjXv7gFq7MA7PWdQPAHoUmil1r1U2ZupFqBSEBGbWOHe+qhz9m
oRSg5MiECUfp03N7xlqPBmUNk/T9fUmau7FYeHTfTOqH7jMkuNnvogiA53/uW8Jf
XqKDbQOxw4DUwN2VC2lIG/bq0NC9gLG4KkCgz9beXJYNMYmIhWUxutfR/6jeLisR
hSm0lPxAPYwlhIIAVXOe1txh98ik6KZjQOURPUdvS7UtqWEBPfbDhFYFO1161bxy
eC2mi4A8zN5ScLLN0pMRAu9tVUMD8wmHtryQFhJWZUezzcP/AWHvRIXbaTJKW13n
7x1iA2IYVjg0ZLjtDZuceTrKguezLyb3fXBA3FuK/dtPU6g3cVdmQ/vD3VQAX+JS
x900NfZmeZX7E5hAEgv1uC3UGB+jExW5Hh61R3jEJTNN5QRiM3w9hj5t87cFCHIN
0j5PjoX6/xwyh2cXK0D0KO+M+pa5sZzJmvxX1ogVOU8m0oz6wsMHjA+jLwJzzbbS
yaOECucV02Ce60nJCkZjqoHDrm/gyFdY1KCerTodjt/nd0Vq3bmTN/RjYpbZ+Qam
CgC7rFRUXZQHVWC0kc0tM6himfpMs2v+kTtKAyXOOUt7XcNFdvyVbSRCTLhg6moD
x9I+nzJ/+gzxdwCysZx3+Ko6RNEvOKPa6SDbzhDlUk8/LM8/l6izTSLu48zG5eDD
dJ1I8a8Yj+Wnzym+95NOQRGu3aTzcY+uW0HoNBUlT78GJ4Tj6o5o7yd0To603KIM
Gl+3DIstMOPvZe1cgvCQI1QcqomZzyxGDaUZ7ynC1QzNjAG5QXC7u8RbGaK8GeqH
Zh5YLEFrKuVE+TvelF6/9QQYfnYcyfoowlL4l0m5ON/HjM5C4roxufrXobJ7P4+1
wgM7LRx2Wef9eH+o36d08c4U62qnJvwLrhQqP/dOfD7acIprTFHrsj68TxNpkE5X
8wUcvBPzghl15hRK9TkWta9+mKY4cL6kI/rf+jQE/lm2svOdUSpEyTt4kGNsMXBM
ETLguYK8NYF35efYf5gsRNizOVk8N4L88tdm6FQFE9kyZyHdfmYlclvJKU6elLTx
xiS/hsuL6Go0oogvCl6/Ym5KHmlTJVqUcPHUYH4IB7pcGB8BqtI/KCa+5zbktGj5
RUZwnazIAGzJYnv+HJ6TH6QYpWgZt6Z/r/r4d5xP5s2rDV3xDGdmt5WaYm9Oe5cy
8jl3EEOTLslHhXkfvjjDrhABvUnwdiT6xsjgzxJbj2GmiR7STPBSj1LTFHP/RIA+
NhEyoCqMp1LXxgLETI7mhv9lP4kIe0dkHre/TgyRkBGc1PEwpbwjjUFFyJ1p+doC
6jwfhcxAMDAK7S8+QO88lgO5YBCVHG3O+TOWC3CjJo8Y6O9E/GIK4qj0yrg38guD
qbBy13C5U1hn4YDlLSImDUZQee1gO1aalp7oAEiYcmyIaW+RF8ylF0ZaFKFRsbr/
lTi7Busqvnrj+jhbb1VRd39SuJuO1tKj0XmG4Ko2wWXwhIpntVixYscBZYRTibJ0
Ws6YQwrKwWP18fnC4ag1Bq68bIk3jnrm5/ZXj3EdiAqHLGzngsX0nteAI42udbjZ
qvCM6MbWKsFYzO0Do6ZQqDYShU0tkAtQ9eDnjPf64//3y5zB0GlliCwHz9j+MmPJ
+gn4NtfgTjaq6nk7vPv0veK0V2HAQ05JQcQtSe+t3bRGUtiDETRNZf2SxSlNO8zR
7HZmZI4MXWngPxS/ioUbf+ZERJqAax/A4b1uvGpuIGOz42wSBFZHc6YMJYdQ0pT6
QNvoqMpT++3ZzshJcRtNi0Ew22KwNg9alOR7EfleQzDl1Sa+Bujil+Kp7hjgKyWQ
o86gVfzns+CE30TGK10eGBALqmcm7z0HjW8GEdZUbkMjTDd2heyLlV0a0lupqoTh
8J09zeq5Cs4+t8YLh8SkFMyVtIkCw/APBX0cAm5Caa7j9pXTzcbv5Vj9QB9HErPo
38Fcul9u+hxwRspdyyy3AI9guMMmcRAp/zSqb2Y0ngwt+DB0sNCUJzND2/5Agove
t5zH5uUgbItOzTFcY19wwvcu4hkWh2NiPFffbUprLUE402uPP8iK4/eL3FQjhIHf
hsqCKgufdTgMD6lPo1u46gGmJNTc7322H8YkEDp7i2twgaAOP6zIgdt6pCSJO1IH
6tFwr/VwLsM/1eKvcp0xvcTiszCc05p9/W2+QhY3ZdPt1kAUmol0x0YiiUxOWSHY
iQG4+sfr/aYneFNjLaKbJS3lYARQppjK1GVBMJAizBGoXxTi4ItDHDXaCUBgmg2b
2qKtxoFsgowj2mpSYB1Kbkx3Ildog8vml5vUOLtx1BxbnLAphcymAe2uXCPTfC2i
tlSncZbcBeqTrLFjiAn4lw05qN61kHKUZaPPx2PWfUr27Md/kKWXJS0WYfsxM3Il
tsjIWd/1iUlA3uYgrUyewYHEW+GWgiOG/b+sV6xVJEIPWH27F7bsG6r28zD3U029
RqBnQ7R4oF2PVeLtaAeKbxh4InfE83BJofERdMiiUylu99kEQfgeZMjrQRwjLbMK
qrxRwOxg9UgT4h/S/nAp0U2mqhtgJHJkyGvu1RMPr01sf+F6ac/GI2Qc5cqfgO8h
ngJiM5eTuhIu20uXNiZLCFEm5UIgc4BZB24In3sVVnxGaH57epeQDf4b8otdSluN
dIDvq8QN8oKwvusZl8+Z13KccT6gsjbFl6HuVYC2oKSk4XvguCyC4Ox7wOtGh3ZN
GfmMJX4qEsvGRkcDyXf/llmXn6Vib7FfCP0TjWTo7gwVEOIKujvA9ke8n8p45qRI
kQIXXRCjicZrffog57lFzj3fdnphsBTHxsyyP7bTiazBjCjtDNPtwuQviiV+VM9h
HyUwBjR1sCPcy5fwTUiUGuT5fnk01QbT0AkmWTWUeVn+i0A7yqDGpYqsFPNRTiSw
ZdFL/rWvvC48oz+4zT1Mg4slLrJy0EbMymL3wqAbrnpFMUtFuik4rMVJEUkkY//d
Ewm6y98UCtpVqYuf2Qu94GBC/wP/hgkRi2mCTQHZOSsDc93PIV7aPlKlYKYifdst
GMkReHNE6oNo1cgq9IeC+SFyRXjKmPWkxeSK66sC2TMWKc/jSCVxIytAZ6VKzMjP
fsL8/ai1ziXwBcrIgInQEqAQkoQf3wNaIfr49rcuU5bFYPhPMVdXxlVqgB3qXu8P
kHzeGV7ieEJDOE1176k7IGgjcdwz1g+5x1JoS+wkivV0bofqQNVDxoDm02P1pZxB
DAV3B+BlaFAWM6jB+waBXiW+5Eh4KUmO9yUu5y9CSffGBsQndXw3Dq9kff0UPWw1
a1wpxM1dbPPtY4HmY0lI4TY4NCxLwKWDGmaJJHWJc0ERq4aMlCUU0wYVsdnt63qA
J4yDtG9ZAGcL7DCwIZqNgfkfVwFB310E2FJIJE596OX//uSNtwSh494HK43rCV+g
t3NbGBUy8tFIaJDu3q1Zo+KAzwlDgo3Izi4iBdA6Y4blPNdx4lWwOEpqH3vgUrAq
wG9vdT95t7u41KzsALMcQWawIQl54UPUGPJ0XqDXDG37QkIq4vQU5ji8+nM1BPBi
2C+eE3wgec82I59IYnh1C1Y0JXIyo2J86Qw9kkMp2G6ryXCLlihgsx2KbGP8kmZ/
OOSzF0qkLySKg1mAcp5RnG8lWcSSGXQEZllkn2WftESQMYbucjtqOPR2Y+Njd0PU
9dAQ0O8QPKK3tyxDlV0hJC7gVyrz8T8NWyaiHsrabCZdw28co4nVf5zJdv/qCrqM
MR9vxJlkipi/CuHneo+yPwas/MvxjxbbmI/3SSd1n9/gxQz+lr9HmftsBCb7Jicg
aPpvPK7f8mOgCr5OOQ+SS56rC838mQCbEYCD9M3wRCGmOnRV683CMEh2SzAqTgGc
iUNB8UcCIoVLEpCw/S+ZQEJ/WkuXlT7PW/qA7qMzz0J0OvxBrrIK6d9w6arsfej7
bliqiejh1eYRwaVfSBRo4bFjL8RlysJO2KXxrWmJf3rBgmgWk75c60w5ff8sogdG
9LHJM8j8agXCwoq4+prFrm8GQCPQrNWu7NfIEEcCIS9GBt73kfQDOHonWZYa32fr
B33rwYurYvHWYvyNersd7X8gleg2KkLKaRATrSr/+CEOgjWhpgeZxGbTAan4Qt5K
5zw+7ut6ZbS2UfNkR4ZVGL3g15Q63CF7/9cR6mbu/yo+JpquGa6qBJ77Ml+8OPJl
mTwHPPvFZtzm1cV5P+Y3X4p5PcRoa0z0JOiR3c3vlmCRrvubsQfafZBq+kfxT0F/
WxxKaNzFCNyjRSQ05z/NDXxMUx6xtHWGKAVpjd3E6j9Q19OPWgnpNvmmpTyVlPDN
fuDmcQdf1P7HtUhAzLEzMDyOdRR9UUkXjzj6g4PL29QI43Eii3YyW3pNX7zLRLTd
ZjYZwQDnUN8RNVuJbOy1vo9iwha4wdQVZCJ+hnJYtz3juZDmzAs/XV3BWXtFjWLM
DjZt6SnWOhK64rDnx5+iqsBS5I7Pax1ADoIjM6ihW1yF8dkdgfVj3iF1pHTzQWQS
ElRIdIyiPsBs8nOf5MA3lxUqI7KrD7AIzxLj46RnAi0QjXKcI2PFKS1I8m+P3uW3
9YxxvC4jgiNZeic5Z/S5CKOuWniwlo9WYryXoHMVHAaw6QD+xfdrmr7f0zHE5Iwz
r2sBbOwAiuGrkM/Zp3x0J1MIBi8J5+Hyss2TkPw/D8ShuwS5wQpYk6PkbpouxIcH
CwRGocvuEu5x/5tMA7vz2GA1iyMwInDCdka3mbLFQCwod9pdOID4ungHQ4qGJq/U
E49r05PoIvN98bu7M/n/26SvBgyVHfkFLEr8vvZY2uyEHUNLjyqd6goUcvODiswu
2WhUdkMJTIoy1IwQswb/yjzjlQaHOcTaRJx705qgsYEOEvRQhR3eCaQaxTKzm/bY
1xRqMnlHu0WKIineDfnTK5W53ATe2l3TK3VBbh84Ox01S0X0oBjYzkEV7NGW1OD7
Cf7lf0AYUHuw0h0vL5ON9/zR+gAaJNVOEWdujUCjmmmk307I14qWLyiu+Wa9K4vB
4QM7Pb7+BeXr+ANkxN9Dus3UJroA+Pk9asv8PXepB5REdFrPVKS/OAIcMMS7YykJ
Ie9TI7kblDo4KfzXhRS6aqV959pRlRQ0W7eE798kZZ2Qx+YBlt9ns62fAzvs3Bl4
o+Qo/eDdfiahMp7N9zFv1d72QL8x8fOVsKRlXMhVpufLZj14OAQIHgvezmeV4BdD
yuVG4uh1gGZbPRDFedKGbFAesyyckJrQNS54LiflbRweMfroZJMNcVcYsXc63KeY
vocac8zL/pFJ/OBTL+iXyO/baIVnyy+zI4d2liza0niGScRLuI8xwki9wUNCZ78A
Jad72NP9XYKLTrUxl9ykrF0HGNS25oWF+wn4fzziZwA0heMGRmxBv4ga2C6OUKes
WUFsH4QvQz+lCQORpVZKN0WNUd5j1L1aHCIvwk6tULfbLcc5ykD/flQ1QI/rRZj+
w6EaEIK8wXkMhkNhS2ENu8e5zVrkqXoa7CayfkH+q2gkSJLZTByc44iIOJKPODm1
xeqAgsXnVAJUGdC/y/VzXi4Y31Y+YmWsi9wzYxIFmNGyT82l9lw5dpom2dnvPxHo
ELYukMKBoJeNRHPiwSEazQGw7Vqz8uXMtY+pk6YFKSft5vn4IvXJ1KWSAC5bRX1J
QaC0s++4+G8kKefD8MhI0O9Wqh4H73zVh6AL8wfbTUiGR7GhdTqu5y+lx3xniGVV
tA8r8qADREjn8fTxahDXym6TbFsbJy6xWTp4r2Imp2+W1rjCEQCfBF5sPu8h9dY1
swmHb8zEpjuWZEIiaKfrg8HtqwOACNlWWsT1+d7bgpbCw/+cJQ7jwmPyaOZQODDG
O2e6CvJLhMKt6jZCU1JQCvTN+HkGTtbGVdbGg8b7kGlTrc7+QPRTWxQC1FD5X2bC
6dcZZ3WPevEP7LKpJ4s16uwHRjGgr0+5jlnw7+GBFwqaicicCUs9QUv9CFibwdao
PMvLdR98yNYkRzCmY33d6ZMHTu2mPKblU2n0yHOf01jqvBpbjBN0zSai8+W0gqTE
ef+QpGChj9MidpGhBCyOwIC1SbW0NMLDf4AozdRHXUVRSTw52+9y1vc+LAzoqIp0
vkUcyD48bWPKWAF4wrpTC3QiDpFygEKhWGazXGwxMysHqtKfmbMv3UcQx4KA0I9u
s+h1EEaGJPw8qMk6fQFJBJWWeYi4drQdOY0PAs25TXufoL4KIl+M5NotqBPB6GDh
pwcN0z09UhiId0ccN9cebwbXkEUXSjQe8Qwxhe7YFi7e6iYcSpa0nqpH8bIIwQpj
zVqR2xwh0yBMxcEha46HhTtBbRWW8wm9YiqhIJpeN44zkhgEuD9i6IciX5jXyjCl
AdUAO70P2l9ePXYbiinvev8bTJbz7hmah5W98u4HtfqdgKDdA1nbpk6vTS6wj4wl
vE7ZPbWIrpN5hX2lVrvKoIkUwDQjBtLd32dNDZyKUhYsfZpF1Cb3xRFtfkN6C2Vg
C1Z6id0cPbolopVqB581U2L9zbm38kjwE0PN5yvVlr/GuQ47OGhaR3xlB4LgZ7oL
oNG4Mg7swfr6NOEt/M3AGfharqGQZDDKUX5BQwWRFMMxfvQ9oB6VCQbZGVZjZgFT
IL7OMCsrBnrTc64F1nPNLIV47+uWYf5UF5f/9hflDB9egePXbVMMLkeDpy2642Tn
zpFN8YgC30ngXSG3oVaJ8BcQbP0MRC5v0WblheSHZZgHW9HBsbAJ35KLCRSmsbbn
y8zCmSOTv+aNrwBJrdibdvGK3EqoNFQRaOv0n6GYK8eVHaVajDtJsZBT2eajxjiw
KuKsJHIfmsvK1alxk+tt/k8MfuIyvnUqMeMqogQaKhdlgsNRfxHr8pDURWbr5HFw
5bg/Ddtt+TGXq0jUXSoWBY9kIc7bmtjDwxedzVqfHxp4plCurfMFNFPJ86TMg6W7
HKNjG7wg9y5WD+xJeABQU4pKJwlbnJC/tkeDnG3ReHqqGJj1p1z9gcl1pd7IMRv1
+RaqgDoVU6/IDiyFBUQs5ZU9OnWGRmBAPaLUHt4ykB2rkJYWJTUMq+JwSowcefab
LcWXzqcYUAA3mMsE+4BowDvgBLVZqjfIcHjqAt+nCezASZ6JNMZvkA3BvGn0Bho4
UmtGISSR9Oc6wmSzA/OPk3Uqpm5GokWUlmFGxg7CNc28aKO+1PO/1SGJyvtrguaT
d8EVBCad6eo6hlSm81EfAYr3vMIXCv6IJHSLb7eXon3FykLDxDOojO8+phmFZDh6
g9xnwse88jFiSrY1/VH22DJ5igpOvUQ6JDO4wvJ1C5BrF4wH3ZvbjnN+28aJKcTI
Vrr+ar2SAoQ3yznMNwMvCZo9n77sSeblr31uqnPCv1JD7HNG//YiXMmQ+X5WY9tY
0/duCyy2B/7/fRVYntuNYpQ9KGs+bTxLKSXup3ZZE5WJw9MHwiff4OfV/Tf60qLd
VTrrUHypo2gYWdtFX8lTu/Ovms2j9EI+EQ1D0f4cJF9Prv21R/7vW2TvAko1F3ub
OGVcewvqGMZ2BUS6XrEB6jF98gcrkIgvaze3fDmihPf+XG5XifgdmrSM/pxNUGmp
bYL7tw1vsg7bXbZj8775pClik25YFn63VVc2RbyX1YzyVff8W0ZpDM2AaUk5yoEa
A8w7YYz4HdRKPOGwMaw07XECqqmdJ2HpbKILSu5MV0K/laO5PrTDF897Bew3URWs
S55In51R0p/tPCob4BFXB+AXaksOeHCEyJne4Ar7VUp7MVh9BkB1NPphSdq7ESlO
b/h8xIrRpXSNbvPANipZv8FX8wHGrGvuRGnMIPJPMSbP4NO8G0GcJXpEP7zIXyA1
gg8ozSIgLVR288g4Xdad+SpgpEMCDH+Ui7W0JG7oavmtXvoMhVI2CMQ7qKcIJOKR
Q1yVPFbf+JRh1AJf1zeDkGNQpMHMC4gsWMYcuee/MVH7zWv5ctC3Cne/KOZgJy9I
gN5G5BrhXTuzJS7x/qmVCon6XjIwryWIlkPDQNdUyS4bsRO9Xef5MggHmr8HWkFM
EWmSFnUCwwpLFnkOU5EVk/8VwpPqWp5094ponaPOmrpOi2R2ze+Agi32f6kuUFJh
slBdGZiWQkVfeQclPLtVi+Fsamv/JC3dYawrXwkROczBfiuKL/OENRyNTWei3TpY
boFLaA4VhLRSxO5ycjuxyu2Sh+9FCJsSVBN0f0jgV2UKyyUuI3q9vOo+WGRQxkbG
IZNIXPDvxF6tWGCRoW1hU1uocmpOxxE/j9uRAy7puUjyg6W2+KwomP7c81bKSjuu
SjH0PQRBxY29aEAiVdxv2ui4DVRZeOHNQf67OIQJbU1VV+zZBUp2jLRKU+etp+Cw
WaEfimW1F+M8YMFIV+4cheQ3RM/eBVMVerE10JsGIkDCo91K+lCHbmBZ/nBhQB7A
HuK8thR1ZP579xl1+xZfHn4kDL2/Gbcyfl5lGEYna+d1OQrZlyeQyV7h2eHDBf2M
k12pDilbzYQdjAiBwtCKpOFQbNuq0ZTo14rTNfMgNJ1u9R8m/nVZ6zfukKL/ySpO
8l77JNSjDOQ/+1GWojNYGgZZn1obxEkx/DxPTmV7rcizLA450X3gDAzEQ2WAPoB9
Ud5A8YyT48+nHmQU9DuY/q087mtfwezGyHp4pG7WwWKKTxiMBME6A7A6wtsgmJtE
ejJ5OtjKMVbIsJ0mn9gMeHU/bAKihx2ci7TRpUHkZyem5zp+fOI7On2Ge5W4KDHE
kz7VVP5swg74ecE/Y8rTSgsELICQFBMPr/lFrwfD7vDfVZr9USgb+z5mQ0J0XNDd
XNTeYIiUrVqYGToAZoYVVKeJVnXqQpfcDadrdGlYlUmyfrYLyS7tKqAieGKggbzL
RdyvXICZLJE1pq9rGR7ASgPCJeg59TWH/5a59YjBaUEY4iPOBOw6G8wrSykJBfIv
9xrRPX4TRV5v+nDlu/hgsbZAHFO4fqrpeIQH2U0OK5pZHjkrPLrVjwnXJFYNt24O
x9P/hSVolxiJNJVTHdTXtnP1lUOgkGjhVBhxmKaj12e9fg8Kl7MzGCiAsRGNma67
Yb80QI5z9jLoAroI6ATFgnCJP50coNCfIdIrog07gvPDi+tl6xj8wSkyKVybuDOv
1P1WrlJilbMKt2GRUCoEWQEGC4Or6xp0tmTitEc14BPtU7o1P8Kl8NIjDsvhA+IL
yZ6yb7jiHBDNE+jDxe/wdNlWwaXXqlYUzQcUNPaIIlxmRFrsGQ60TF/mNT+TiqVb
OMnV5aa1xZOuEfznX0caEZy4+1YhXmjD350astzOUR5i3VO56C3iniWl9UzS8MXB
5rBTg4LjFyhJDLxRdQ4Z4XKenxXsnK/p8zCkS/OrgzLJWHPhz0rY2bNMwS8CxLtf
HCC7xoGHqO+cLVgyAty/hgAFaciBYo7jWXg7+MDo4ekoMYmvOQc3pds089J8xeiI
Vr9byHrgxzaCtd5NJboIOwn1vDv3WnBp407ZxELYjqpqAbUPhqBGyl4kWs5IJwuy
IwuD4lfmypAlPvATK9/Wq5wtSfxQdXqAh9Exe+90gAUfKHa2vrLLr2kvCkJfYvPJ
Iv6t/22BGRlJ8HEKJFg9vPrgXZfgF6mXGhjuJ3RnOBe7H/p1j2BPFiewKUIYTpIV
KJVSRwGvsFnqDJSZKzPan5wQ7wu0lAOeq84TyKGmICCXYbWSUFmclEHzpAfVhnQT
Dki9NwAx78ScytkfG0EDCtZWuYknCUQjSqC21SPjgnx2ZDaPkXTghYBC7gNXfvGM
n6Nasd5hjBXldfMtKTK+QBVbSA/ymoGyfmGS+qng9zJZ/EyhvOuku7OaKbxfs0XE
Jk4dPd88FaSA81ELPKdFGJ+ZoCAB3SlAUqoLa6ujRcEiNmq0N3Xn0kYQJDy52buM
hZ5pZm62HmD8PXaYsdhjzYJ3qmueSt5G3LPTJK9m0g8EE6Dyq4CDGkb9Un+OySMb
yk906/qHFSjEQbrvl2rFjf6Z2aRFLjZf3Zrx61obd1DIaDTO7CQ+ClcSE6ZceSqf
138E1iI94TXaj01O4YQhESS9gS+Xgw/Po+lOjYQ0kVDCWEXzxReSnBIoBjJHaXVZ
sUW96yJUM2in1TBH7pmXMZnXpglKkHIYHx/AAFUIUuppwZup3W0RvmHH+4nRpQB7
ulRKmeGK+gLGTJyDSaWlHHP+MfLkPY4+UgbiEBbevhjm5O8F2mML2c+e7Wm0AHVI
rMXFjZzd0SbajilL6ih6XsLgAbUcF0yfKtGwpexcFO1urTMOM1eYmUrBrWfyzxQQ
62X2mZMtCZ5Wl74mBI4BM3QeH2F4Hf0w6BkISYMy1cPcNfGoDKtbhilbdi6kqta0
Uzu1+eKNafGfF7+w0ZjK67h9k79UfwlVmvAH1MxHys+PKFl1lcdw9Vne9+4yiQIH
AEom5U/22SHiXNCnemr4WiOLKIAigkCaz6m/0EwdROyZLULm7VXT8KXuvHr9u+hC
QT16DCoFsJSIL327g4XwwpyYMSEbG1PPppCczKYvnhUTGAnOT0+VmZR20Dg58NXg
mB4D7YKy0SQY7D7X43vNb/NBByu38y4I/NmFlhKVEorN5CUJ3u5rWDYZU5jykHav
3ZptNUsPVHTRtHxfTN577WinDoBXNk7pLQQ107Vx+dXTC+4zt/iVVjhDile/K7an
O0J6IbI4llMapS9nufG5/MasFsWe1Bkxhacrd/w1sM17uGaP8x/SWM6Z3tby/R/4
ejR+1AtKPdUdoXB1DbTYqQ0+S79H83h7h7B0Ws3FjdyIbJBecC6PzDkB50FHUOwm
10NgyNoPdtD/CVn4clBINt0KeM3KD4rmbl4VWaOEyv30/6GLHY4QrpD6tQx09xvN
m0Ttbdp4xxG/XUc2YFkHAKpqjlq+TeIgdVS0lSaZeYKAm9iZZXPnxxD6NuyTwjsu
uIDPMvfGG2yve4JDKIJMmztjCW2YcdhxK0uLi8ZW2OYCJLKeLu7CRhz1qq8Sv++Y
m2nWF+YaMaPCon6K0JbHaLgLSAT2iId6Y4UuUtTRCpVzknfm5BayhYUGYKTfA9Cz
I9Ih6IEZFla386B3gGDIzk43dbY6okQFF9AUG+2GTUHx1zjfUhQuBPglJELnCruv
+h42oQnLdBjJJpS5VabnW5GJmrXIKn6vtCroGbMSQ0ule9TJYD9HWaD4yO2/zNOX
jEaG0Y43QgzUXobai2zthIFGY0kLPBAT0H1YtvoQ48DmOpY2dQSSlQbHmwM33bI0
qRhZrv9c9rS/4szzVcWs7sZbqxRcc/OF+smHSFmMCUxuB/DOreIKgaNbG0pD8RH8
ibhG1QoVf9URBLVK1ZNSAuckANtMRTF0NNTtAvgdHrIMG5URLhJ/p0ZmSv8hr/Gw
FYMhxNnrfwGuABSWYu31IKGWzlYd2gZoCP1AS35RqHWU1laCXsdqBq8S/d5Mv1Lk
39bxxDcDnFKStS9kMpYqB/VzoJNZNLgDRz9Rq0LcCLzj3ZyCJFmICTNPrHrk5Nz6
OI9XORqz8hy8ijnxICiMYhsz7Gd1kDwL3vNgrrRcesh1s/zZobZ5QkyFEb6hX6KL
jeJwaJNuwfrSkjblEYRk7s1c0QEsoVdL2tPCHIjWvM0c+PG9oED8TNF/v5Pt6DUg
/7MmpHei84LAcpGMxx4JqRpILPo6E8tRSUs765KwqXscz+MfoY6GM80JQRDIKocU
9CTQg84hh1PUbrEGZjRfoJs1gI6Dn/1FZXoaMke2LuxHd8S8osQJmufUzdJJbWZV
gjlziHYNhR+ZPgiDYC/XrC/uMRcZCaemjWfBQHbqMMqppy7xasZYXRB2Spgs3k2s
jMmQA/FiKEDQf2S5WGR7CgGCp7bbT+hfD+d434tHuhbP7/5b/TifEQRh7BtuQQ4T
LPc52nWYCw/4diGX9t8THNSMcYFuxfS2JiNVMdL3XNGB2R6cRrUUKzi3oXFD3sIt
ME4BF/MMOYOyr8SfWY6JGuzmap+0kOgKdzjxrFPD1NHUDbxbEh5v7bjIzE3lEjcb
n8u2QFmL8Acr9mGdMgLMtuFI35rUSDHmLkrpEVh/HgTHnV/SHM6f5TyNy98KDP/P
GKoG4mbyh187sgwI9hHL5kX7IdhoUyTMZIoZJcz8zA6zrQOgg76JltFMfttS/a3n
EBFfU0WpptNwXic1IKk2DtQbu7lMEYqHvKPdyg0W+aQG1qpAebP8b27CFBCHf8yD
VIp2lGX+RBjvqHS5wvdMXgbgXUF9WN/7u6cH8eKusAHy4wxV+8n1lSM5n6VFjt2S
dRMcqSvsgPG0lAkdIseyDQLrmC+TDxoxHyVHZnJexorWFlE13fsRbJQIoaIjA6wd
nze2OeveaajQIH7JHaRCuD8LC3HvVM/bEnj4JW5jXExtebOjleQontIhTTbyeWTi
fVpPp0bQWHpXW8YOlPurPMk/6l2bld/vK32PWKkSint+BRvtGr3/Kvi/gaa9UhhE
tV/iKUqJBksp2/psre+poX32Cwq9gLoQHZ20Piurl3RVtYhYS5CmZdhjv2ugufN7
lkVgYSVHo0B1EQSQEad4EwdQ0sX9Fg7F9oa/LO4vApI6H88yDxIQwesNogX3d3MK
MIaHViVZjo4lHf/XBFOtcgAf/ZxvueV7JCo/GMI5sYsFwwP31E8hdWUjruk7zu6S
EE5dS0dM1iVSe9NWVpqYFXz1/ocflmhCwyfObHTLbP6BHvWKYUXNauYhPRJPO+DP
LXPSSLaJew8GC0YFa55akUisvMxcAletdNEAStxqUHagBso7XivU4mUAzq4GnznW
+/Mxy93iiSB0LlA5BtxTSqxkPCbOTnXYeAWiJqo48A30o4X8ymwWGVkfB/i13oxc
y4owLgv0wFKcQYvRwyg6ZnBdQ3L/VqVwq82hBD6HmAqaqc4mvLgZSMA89ilXQ73g
1dYW+tPZvF/0mgBBo12ftfpXyqK+UZ/Tvv2jjzT6VDwDT4SdyuoQY9NNv711R5Tp
yQfddSR9bo01/fnKZ80v167z09CnNwmDyiS9A3NFxjQAW8E7q32owRhFrGII7tk1
fpvwi0GidOt4TmOEDeSUmd6EiRxdG2XkSkKc982UlacMMQfxlrQ9OuvitR8MU3G/
bJc2F2j2TZJvfm6BwjAoqMadT3lyimoUU0kfQbElIgDVh9oEewqP0quzp9aN55HI
yrwMCGCtvE1+KQzqB6239cRQvpJOn1rtzCRu+hpGsrQHMKalw4JpmXeZS1r8y2HH
CgoKwyUlRRqTbsgidSPP+iJ6+djtYJ2bv48YWe4WiC29QRMtnJ8v3Tiaq0wdUoSX
KPyj5I789ce+cSjDvE9bJVC5Ufak0de4ePFrLgbGIAkEk8YDwngNTLei9TuLEtrb
e7s3Iq1rCFEticnfg3CmnQY4dzNv4koovObf/eHnBP0bTWN+/XxV85pBnhYEXTVo
5iSOgOO4QcHEv77S4mI4JN07NSF5B+f9d2H38by436oVz/7+VphzLQqT3UfDZLqd
Fol3nYO4CaHIcIYrMeXX5BfPhiAytley/50yjRw8sRRi6mc18tnHSCWstMzNlrao
rb0nLeHuLJ8KXNZ0zrKn8b1fWxt/GPAas/CvIZsZqg0apQ4IIkyeDYW5RH9L6zzW
eL7WXtrsEJBN5zR2AmaaofRuon8HNoxT0JHJVipLlS1tSohlux0uNelsJMGfR7QB
qYEvjawxXNLbpqiResQREKdznROJUxtHpYfNad61/Kvpno8EbljFf2tALV/boJeo
/h17+j8W2jSFVlpXEa3bBVKloTj8c2os3Yk3bstPZ7XKYHIbE29WR7yImxVOPGJ/
WJvkO5aKHPo/gMMv6kigqT3DuDvux+J0mqHc3Lg6ChqK51wX1isC/R9mDDl4ztn4
ihiO4Hb/f9Ze1FiKkW+11zTgDDx9duxrEj4TIO5THvPZjIqVJtoomffV4aR/M7zS
HG+16Mrkvs28QersOm2Qm2hhH+BXDiwV8XQ6vsvOINftudR1zy59QgT3DaMqStlL
AHkeYGVGf8uxCZ/DjaXyg34taYJ+WHhusRfayZvO0BdmwIJknJFvxP2gfuUhwyIp
sSJBydkoSHBnKPu5g17jIgEr0A2hwA+Cd0Mtv2ogEZJDIIbJ0hAnChVYjzRsIHhO
r6UGPOw7TY9+XbZxscoIQ063ftHS7H4Cc5Rky97aXzhSluIeSKWm8tVc0i9S+VZ+
wW1ndI2tdCBOpeUXfgPYjR2G+f4Dpr5aJ2ngws6A3O+DGmZkQnXEr0fWz4ik1aDA
tslyjdrddZ0iK7AnuGP27990Fu5W2QRGS4XtMnZ8O8iBgX/MqQrIpwp6AHUFJ/rd
5/l5qJrtlVIFngsBVEBEAuzEclto0+WjCM7i8zFCrVH8ON3bhURB4fsudG4BgWTg
27BjEzhpllZs6L1oDxdwZWM51H8MoFCZR+u0iAEKIEZhZSvfpaj5rg/D1G0p2rNO
gEM3VHeciCy42CA+PeJt3+yBnqALmB4AuU7jUcWmvfBzzIkSKD5C5cpiyUs8WJSQ
lwpWvn0bbaExVCdESue2YJbZALC7lPS4/QbqrTxtVomalo4d/0pJ3p0wd3PT89Mh
zHOuo7yOxzWc/7GMTY5Ft3duCxtop5FBHAo8lOuvCgSVfnZIRG2A7a7FifDqZByh
Rwcpol4yc1xK2GGx6HEwf0YqDMpkGwVm1/M4m/0dX7FivSF5+7W4ck7aeQoFUmJk
gbltfxAnE1GW38JjF7/RCNpEKPePVrZLmY8DteCuvq/qWW4oNSAgRWj1GVy9F64T
noj2uEWeahjwzSHyPDqOaCXc6SDywXcLR1QdUXXS/RWZjv78Il/vHTmlB5da4idF
Y33X+4MSBoT8x2ROduqmStl0ufRRtMPoLhIBht4sJl32uRS1Fol388Uvs/9wqcWi
qXyWRZzQljjEEzxwtFkY6bQLmDAKcwPlIr8QtaUEVFWDF0s9xAp7UYh5Wp30fYH9
eXdnpjbygy37Jqzv25MPMAIQK0VKsibE8rLQwGhxBNBzKEmmOaPIWGJQdnJS+bns
/cU93lmTs7o9hb9TY+JlpHOLbi0MFkfN3EBU7YOyWjN4+jwvRQFzWYe1Z4zwESCl
IAua5FdGVcKLW2gPlVKCJSx/QJRNn8k69yMUO7gIxJGXFp8rrFlZzauNxWO2xOyY
dr3WSDnaliVj0+ZdxJW8Z+6uJcBmYoejA7cylzkIqV22zbRGdY5u47paShKoTzSF
ii5AXIXZCLMPafscMX4OTxaYYFJaUzSIcmM3ZOUTCy3Y1R9tOcirmOWf+SPIPQxz
au4nBoLsRs+/RbntKkPXq+3EfwG8j8gYxqGYZz1sdLfAHndKoSUREGTHjW0mqx2H
ikLy04FbrqJ3DKgz23mMDukApr+n2AOS9aOHk/3qcikZYfrJ/4mWRXo8qFpFDacn
wwEFbF6aPf22QDEbQ7qKtwd/VCKd/eXhMu6pOwN42QNKAE0ddK9HkQ0AxwZrAapr
XzOBHWxamp2SdJq6gN9nCYDNW9MSd85O7iC/LL0TydsunwGEIg2VFexmPuAfrJEM
7hcjm1U7hyaRf8H4nNM0MROwf4xd8oVTZrnSAK8/iM08RTQ+fYxhZilgKs8bwf+O
5MOfjzLPy83d6JeltBu8xNk3VV3gmctDBQrD/o6RwS6eyNJC5CDZ9+UKYvPFMFr3
zXJdJA7WluPNNwA/uWFxgnsQrU4lSp53q901qKfg9HswKhH1CMCCe8YZ3t8NP5KP
saqyP7czxyDFo94EHIl3VchQZVgZUDjQ1tVIxHDsDr8y+qtWK1n7DFE6nMcznEcn
Ldv3ZEhOhktJuXONer7S4YziYKj//ghAYdJ9JTgsfDVriiMBz0O/hF4+sxPHO5im
Bb0Q+qBq8Cy/fMKKLUGeyShbgxRKZlFeoeYiNZkcu+JHpvrRJVkzAzwi7r79kxYR
5nBunzQQfDfE8srFcljaQCqVLB4S5jHHRN/HEdgr/O2DQsA1GD42eyl4I09Dr/6M
jSlebzrPuwu512ZcRmWmpwZH7CXfA4UV4Hv0bmSos/cUU5wE3xUf2LTsk9hsQAzO
Zx3iinCL1XNvhrtIMVcIfqMzs5xBaRGWwrK089y6/Jyk6uvKfW/9xsLft1rr3OVX
sfRmQgjJHwkMG4hLWr0GYUsQWYCcF9jipeBx8IYodUEp2g+rVzn0CO+Cdv64jolT
9cWnzsR076qICzsQoAZm0YBXNsLefGLMJM68MArlctbvEPTZf+k6G/3uiEIqNUcO
gHI1UNAK6y8rtu1rfjhjIgHB4nKFC2tiAZ3K5TOK9WHWYCYAIWNuN5AvWCHvSTm/
b2hirulFwsW3vosFLXiV2s36wgDhbdnSJzhdi7Fw8C7YZ+gCD0gO7nLs/bnY/3QR
sM5lKNPxkBY9mNbZA6ddDHsLXmTz4tPeHLQwpQpywiJrx5oNtd/iTWU/d1m53jEm
PO0NJLiUbDx5SFn+yDRuN82kVvW/mEqW5VgSuw1pzpCXKf+qLsDnuLLGRk0D82UP
bmtGGWWGfWH9Ru7tvrGD3Lj/rMBnCqFIC8zKgiIEk6QG9EwHLxM0DZIJOuDzGLFe
3nlnN4Zhq027APK/pTm1NJc0KcbIMsY8lr0dvZ3mIuDqurSQ8jeYBrAyiHeYm/kB
wF3RdhGYVN/8M5Z31dw4cviawUYrlBRsc1jU/uFiE6MA9/MsBriZLs1TFub5uImT
Z4jc/g3jUSC8JRR6qDCP3P8q4w+AImT/p8x2YdHjePdht9a/EwfpWLDbMNCGneD2
fDaBeO6+lJEuuWWnW5ulqT3xAiCif5whEgmeIhy5E3Qj0mfsEwNuu3Yp5gWPMeD5
b6GCkefcXn5mRXpl2XZHHEGDamwF27pzGJxVYc4r+g+GM+4QEVt5JP5An2bIGSOa
l0wGa4hiKdBX9ueB1o1Rzll5YBVbS6rb8oqoDqSfImYxze5v9DyiZfuXjuYfvrQ0
G5BUCqMYjg7Ml/9JewpAllySdJforsKjk3fJnHnoTT/GMJ0SH7ygb3cQZUClQttV
F2A919Ua5eB48xeqPlgNSVaelbIZ1Nv73gs+7DZMn8x9GkYXzWsteeGYt+vuokgM
tcQedCXe3oRGLHdnmTv0NnsiH7sm+BC2sVa3PALuuashE/I9PeddzWQt4kJ0xCGi
lfW37o3qwQiKWio1Zdu7jyhArUU0jMmguOnJRykeL/oTn67rOlfaTX0NF6iZNMAH
8QMArXkF83S3xsFJeDwgmNEM5JkY/JVUj3yoN3xsbTpR2iFly+ndrYEMS/G9Nygn
Rquv3/IpHKfPIE7K5xRu1LUKdwYsdJjLFdeFQXubCbtDtkdNvBagKZ0ByD3n3ccZ
/l3+qRJIIAtE5WXAUqfthkxadRuvbx9fdpY+HxL1Ws4AfZyoStcqRfk6zA00y9Ed
k9ONFpWcFVCowQVQ2CiW9I9zZomZxP9PVLbyRUwpkf7lPOCYBUmxCDczCpWl1tmE
bZ90rkqreeK9vsC0rf/JNxL95kVGtLqGRoX+1Y+jxhB2T37yPccKkBwZkzFOWiJa
V4XcqUXhKCzyo4U+MKWqW/4+7qxxSRtdPGAiiFt5gcRecP4sQEkQPsC7Edd5HCHp
nZ+IhBxyUJaNGRHWHhTy1wcxCnYxUCKS3LuJGkDZTPa2jatSFw8gLLCZwkWV17EA
205Vr4rupHoO0pXs6vQQiMCs6686YrGAITWKqvNPyic6kdpjaYHowAODdho/yZ7a
+40JoaryHQm+cDds6mnYSOSeyoCRn5ONjJLylNrvFXUxlM+567A5b3JvS3e5EfUj
6g9G9bwbbAFAPa5sz+MmeJIjvZIDTZFAw3uPxGjn0odf1+UznvlMilW/bplXlQGb
dYK+QUfG0alnsYSfCS0LL+4TbBw01FM3kW4Dh7mfwY+BmdXTxeCD+9rI0hH4aDQQ
STe627EPYv+aWG8NA8Nji+VeWz3Q8YY5LU98P1x12VER7Gb2dwROQ2U8JSg3WNBM
HRROiuFSvx7m4AXBQqPP4SO0LvD8HVFA55mpGGI5z4K47JFaM5MpXnDoeM0005md
LtEAZKOKG2pjZXI8yKoulOqfK7Pa4gdHk/iYBsXcS5nzCqkP94WyUAQtL/bg6CRH
3onKqkZCznd7URAozRxyfY9Mb4F2P5d1DSWQXYBk13XerKC6+Nn+ViOw/YwGn2CH
XoI9MvDI8puTYChMHixixScteXQtFHIiQ8EIUOI3uXS9O+G3R9yijbS7v59ZXQCA
2FdIe3Ai1eLEfKCXVLtslitSZEBS2w49AIwVIAlBCjhMgX3HjWBmg1Rf5BvNgLxc
8x001i/RXsw1wgYqdHFFhkjJL935vxU/QjtYrlv+hzQC1BJUHQ+/HM6UiNIiV5E3
+eRgyUAUhLFv5cZYShZxfBR2+dfkC8hG5hctLa7WkuDJZkmuUkUysmQBPTET1AEi
PZlMncQjvZC+/9BlDw89QrNXAvNn4dQ/x56oWeVZSR/LxRH2RHYY2bOX/RCFZOuH
bOpofiyBdKpqqOJw9E7kKjkiyy9c/YD+u6fmf+K/A6WTMj5QA28+RPb5m6zDZW1t
pN5E/QlDiOSn6hlO3mqpuirDY2lBA3uMuGqTJt7j3Wgpb4gMPw1IMOLjnBAy0rwq
Tre1hAfi4pegqSIASf5Wjw3Ap9KmNrNIpOTAvqWRiMVm62kOMkRPU/e5ebe8bjTG
OOzGdUyDvLywxHpzM3GtWR34fadcgLZ32/8cOPoazpZKAx+PSjBo69hlKwaJr4o+
HxV/qSo4vCfH3n8QHyxseSAXHXIUSCbhEXyJz/HlYD/6GhcBXItDqkxnXLhJtRp8
kwpyimpKXd2S+MViGZ/qqlAAZmgRc1RftOWiyjAomR+h+3Oow+9yKFIzxgfmrrHx
blQF5X1viy+0upo85c4xiYV2QYVU2zQIkXKARYeu6hxIR5UJ5Am5EHHAZrRVDRDY
2gMhAhE/OlIXT3efUh1iHAfa6m8hab5XELRV5IYK8rT+YbiqvGYa+L0ehFCOsPo2
MbR0VUQPU5LagQ4Klr33NIUaSaff+X9U158fWvMcQvBxAND6MMPBY6K3/XrI67xh
C7j8ziz7bhF8692A/AJydLzfiAnexTLarA2Y9iXVaOIhcH63QO40EgHaVadI3x/g
yc3hqCZadJlK1tHyLRDGuUvZ+0Nq/H2R847pimz5R3kpo8HZWQhlJAnAzvl9G12T
d4niAiVSLQ8QpP4jpt1pNDTvk8NyVRGDG569DChIecuA1Ux/yEpGGQTapnICi6u2
g43iZzv/YFpLb2xV+zry7e7zwQQHbmgQ76rdlfp0Hhx329qQDRNV/yw9UgPWhLYb
ZT2h7SqqMID+SWtEhAfEdyek0SkgPXRxr2se05yeP6LOtc6pVHdShG7fhdlHYGvL
kLlC61YgeO8xsn85muYMJ+7gE77AUgWuoNyHXWH16+eH8Clxu/+D726rDHZxO8vX
RVDC/c8RENiXzNWIt2HVoETEKhvRnXCWVgdok1/b/Qk1VwGQF6lgnHp2qE2OkOFn
kDpbW23L2MCyXajX+nwPZSjt7FiaNm9BiSGr56BQTI8RCcC5ikzKwBDFoBx13/qy
SyYN9HsLCynm7ChTkwYRyhkbj/wGwh/OLOqivpB/DmBcVRvZwHJWLDMKP5AHiQFN
kw+l8HMsDAQF+mt7wjy2JvnORfrNLTPz9+059X/L7sHbK1Q5eTlr8LypPDfgU5pB
tjIZwtjs4g/nnfc84T8OtEHQx1IUroYuhkNbNZ7h3BRsQG2rVWBRWBl1DXUKrc/K
13N2YtmL/gyDpGipEHcpmuAJb/AlxFHM/NPODPBP4ovO7ke7e214EcjUZT5j9nSR
SET3Og3ncMIco14WCYJYwSZTcjuTAtJOjdrXa58iy3R6lBHmSX89Yubnf8LSYet+
19ioPe5SnaIB6uXan2pOAuEVu4ba+1GhJnk3eL2nZBg3Gt+XS1YJvqpHx7wCdSXZ
Hu0g04QHm9vknhxuLh7c8pOfPQXn8MDSJhOpVJdmxMtxtVZSKGqZNtJtG3OmWYb4
a0RH5jgDDbk54eK6XlUdqljiporlA2Kr++IBwLqIzk5ePWdSKHFEpTwCjb91bNdS
sLHsalaX8naSD1u61g4yPeDSPCX/r3Qf+/ZYHlruy7QCeoq+WO1/cQJeVZThZ5U6
Cvjo+t7OacmHTag2PBYxdfGjCadz9ZWaNTqyXBLRpFqEECzTufs2C1vHJoYarXBd
ouYU+qdSHraOfhjHU3WNES8MuZ2xOjIAoYMKPA4nO4kFz1V3arv1VHTdZoSJ/ZF/
+Fw4G3J/IUx4s5dMoXKamKpXre1gNtxrvhCIu9WQxrwAgd1WCz61qOenYUbwyVD/
wMAq3vMDFKcxiyRng4Bo0xgScVpHH5A1Vhb+3qlWRA5gVBBNirid0W/bMI4jLuvh
jIy7fUAkYSWEFfaYLD/WXQmTzqJO6Qsu1FAkS7C0iklJA5d6lnQWs1kEH55jLyUQ
oUJQqNcgLvDQVwWDEDHwXS4N7LKOhNwFxw+All7adSTzKwoSxnghPfS0keJ+/AxL
K+ZPDAFZf9NTWLXJLkBmZVVOE3hrcmHDYbh0q6gsq2rvcQ2Wl0cDyNuFcyAZZHJQ
BCV/5DGF2hJ6o4DhUicD8jMBBzZwXUEbFKRfrGUpxw2bMxblegZvfDBkr4qjkyj+
Z+HddUh7Be2ytWtSYuMDMCfyoEa/cfqyuzEgu0lPxblS70ixBtug4DSOsHCAk3ge
YBR3CsFBm6wGE616nZRWkh9qmoiD8+XzlnWg1RUpqrzgSw5xpN8ynh+9hKF7DwrP
2SLzyT8esvn76CjGo5jOhxABKCPr52fo4weXgJpNx1SOJu22YztSqVngglsLRy7x
ZQWkXfR4fNPUVcPWp7nOi16M4XrfhENkg7vTu3e8XfpCTLl3N7Vj4rSmSfI0eNMl
9xXxBVa/QEBLtyV0ICU+3vWP+PahuHhVh9yb/qu0x9MYJ9oDTcjrMYfT+x69efFe
4fn+weQ8JfRG1mO8Esc9mFqdPtRjW4xknFIpnHWTZ5YhL94Ro1/kXW8DCHfFc6+1
3/w4fLcvXPSzyVYn/JKnrXX86Tk2wsjUPbLcO9VPuI/WH30IC0W8JuXtv+aMcElP
0rU1LHdeBLvvQ/eNmyrJ8nBTTDqFgEWNWsKmLwB/31BcjoSWONZnZDQNqyMgj2S4
XVt93a+DHH5wJ/Wk9kdXZXGH27hgd4392hy15zDl+rBN3+6TI1CEuSYEfzUNmAg4
OZvuN1yx7z5qys+DKOS7oKr/h2v/RCMko3TK2C8rZIxY6xouEL4koDis/nIkn53N
12y4Qm20c7Kpdl2jjvYFhdXJGurYOUb3UX3QznrKVGAdi59P9w8g0e34fvDOHGwz
cTUUVt2hZSEEv1OXBBtVdOMRTbrIXmFHthqXalH3l5Kz7D/kJ75fGzpMBfgIUwDM
yl9rd3e57nDT4/GxLYqYVNAswF8PssxtxwqDk/mkSdxGzjzSyPqpAgpJMvceaFLi
f5LqVCi27p03YxPfBGNoWl8bPto5w0nafQ2nINe+VHokxFC4Ksvl7MGEJMYGkA9/
cnNDu7Wpkkj9gGlDoZ2L35D7Zrv5Bx+zraZ6zpsxYnLHR9ERrexQdKPKtGJF12XT
+j0lhBienTJN3s0jh7HqpYEeNHvETC4qFSE0ZxuVr8V/r8Z4tXM22c6IXAmwP5nw
wFl0vLgrXT1Y7CRfIeduKEfBUwJE/qEVoSfrWq0KoIuCFcwaNlqMFhqFToCYpZzy
V4cxkcQ9SS9cCVTwfDGYAQNYdn5Yz4wdoG/B1tMU1xQmTPg6X5/xv3UZEIgLczB9
4wOew5pu2zN1HL/lokhbJeHi/dV1lYiP3wC8NOryMCiIZbhf8Y/vui932lf3Y1xg
0gEobWYEbkRSLkKXxYc73USJcAXtgYJhtIZkmk2HNyGuJZkNdXL6NdwIvuT26TGT
UjKkqtfAe+fB7dESgwecLgbsL93yaf5qePOKT2700Jdstsvnnx3cnoOB/ULFQdp0
OA1b8OG5BknXY1wHgY23DZdThheX+FM5wnzGn7IvxxUfqzDbdA6l1wRLpFG53xBK
XdyTIHljf1ZNkFayhhz1EHZviVob34220+D/PUulJaOhO/1o4oUazvhm2dpJLVZQ
WQG0LJZEpFGPhvdZ50SNfmg4oI7MajJJlEQaoOaxlD8lPPXcRoPqKo8jeYz+zrOP
4503Vpgoe0pkTmpIb55EDlhyV0UH565H5bck4TKadQpKTG55hV6GzoIVaV5NtkWJ
civNXbejQPrYgaY8cfcPUVZjVBRwYq7vZS9dMe1ywnasMkpQqVWzM6ZG0Ttr00PD
G4A5EyM9SbGTCcAcrLe9kWhF1bEkGElxcv2PQEGIv4+dw94IQyoaEkX3iU+VRcmI
mgoLGfy4dsWAR/uUklPBIj6vvnIkFebLa0yRPL66O+KrmkWGW57FAXzgvXgHtK0f
3J7W4A8Sm6SP5lP8dXsETC7QWZ6TrngGhoIGT4jPO6exlOtxdc7hzLKSxZf0g9sV
y3lYrBD/RELm6/picLFCKgmDDRyra5H+9E9EpY2+H9uHjV9wJHFJkfZhrtG3lnqT
gpG/GlrYeueyJuEh4ZOmcC9rUur10GHfRJm2DGc5LKZS/Z546ZZ/Wi+KOkepVvLw
8BYcLuVtKdWRl2CI3AiCKjLJbmupeiybm5ACwYdKgez3TkFGfxFnr0AZnq3rVgeT
OhlnJub0bqx346qoBpiROFi6qlWi22by2kJ3pAXqhfz71fZgv5ZMyJvv+xtehJ4O
Kjc5zs6BpUlWBoXvZFJoXqJgvfNXMTDNsnX8xfV9Fq+EIdmsHLEnWTphYkRFQmvl
j13zMaELN3+Swt3HmUQBCUkdIuGvvIJkufooj0oJW44NKMJl5u9M3G73nLNCkEwO
uRydJ9uIBduiF1wpGDOmOpKnxfo6H+tAk9fSH8YV6oXjesbnTFZGBrrOg/GShEyJ
W7UtizYTMC1LHwZc8NOZVck3Tu/7b/mA9m/gtofVamVAaFSNMp38Keup6ehpV6x0
PPNLCk3dC/dOLIFa4JrUFPYapbt7ScOCj68XVArL81ABfsnqI0zD+HOgmhnZqkLr
/mrtlKB/Mbkmfv+UYDyYoP1OYoflaYVCqgVMOoUzsCIQjZWyTd+FN+MnJo54SHHW
8MgtlKnSpjhvegEEmqqnJXpdqDNrTdoOKtdnqESDTeYGkX2AduZwZWJPnuiKXWKt
Un20lsSoCvr+tdKLPu5dN2mvbupBpXPU4aylAq4JVVfzykKON9RouIy78Q9cbA/E
b4NQICfMjbLdnZ222VG1aUNwUNHMpAitA59f/Rf+tAFm2nt+9Uh3aCNnNgLmqGJF
VhRvl9DZjNVOOz4anCTPM52YQ7xlKM73O6WMGSIEfPnpcHri5DHiLEH8mlp/B3Co
bBdapXZfNT+prE+W2SDGH06mfDbz687GSzBMDJmwkOJy9mHLThWEtgFr8mUbWs4G
RtDVho3+vw4U9E1dq5JXd4awWvPWAggUBDdd4/FVM/mrP+po21nQaCvH898Jz328
4/HIR7p1cl0+WKr4ijmVNMSBF517+AkA6N/BCWiq+sLUQdVEiwj+YWgKXGKjQlDn
Wi0Qo2lW1kMu43Lo3KOqbGj1ORFk+L4ac1XGGNC3MF5i1Jx2ulq4fGXEcXZMnwcZ
I0fHQqWzn/il4ztQrQKz4/IJn2hOONEFNGzxuH6Lnxu5CUs8LYBE6q8S1i9ZgZ7M
/KJEIHqouxwJPfV7uGhNq0oLjgmF+QHsudyh/zQ1B8hHah6PjFSB+DNrQOFp06sZ
XEGWyzi+FU2jGgJbNN12+x/uRFmeLnWSv7k7awZ1hKZUSD+xLvep9WEi6gRNdBdi
TsmWR93MEVX2b6MtuzhvE1QzyXLquv3QkG7HtjFjS/o/zxTPMVezCRjp0bqFUc/Q
p4jnxlpxC4aeaaySn8jGHQZVFjJJ+vB8yPFGU1LmJdbO1fq7X20noQZ/fMY3ZAHM
nOXpIi3VM9AgGocrfavHAn/EzBVL0ntwLeB9iPOgmOUAFjPnK6sEP5LCHeWWFCzJ
VSpMYo9PJELUAYCk0FtIGMPZibz9tCeUGT7Ezlu3cLluWL/wMsEyyMSl2iEH9s4z
Eot3FjUVBHK7cn8d5XnN/SHRH06dr3Vs5Sw2a2w2TF/q/2FRtn4iofQtbmeZ7V0R
CftBcEWbPauY4X4p23q5VkyKfkAm1XjFJfq2bmoyOd4FU2CW0cUdhfK8LHmk6XMW
ClstotWwCjgBHqeHZeUJJ/16XwbZYWT/bKyUCVLknWTOjmrz/IMaM5SBt98uNkcO
Wx7wNy7quoMDueLcJfShXBSqc8EyjD4v+/M+jN9CvQKMJHSGlwuUSJxbfpy4PFbC
VQbQ26W1V+L6Z8rlKVzG/AK++Gn7SjCp+h9wr/NGrr0a2KerOXoFopPuaKmDYjqy
8PZ7R/TpbguPWxXotCv5rmgdedBgcgUATBlx8DFhm245J8NvO8+jv/l/XD7f7rIY
aHGxRuWXXZcMoWPVmxLGsSNVW7L4OFL2M8214p2Z9ROc95PNX1s6o/qIhD3wsssv
YAs10TmsHqYw5Y6gSyG+kuv9HEVP/v8j7hKWp2fk22bVHbnlqLyHdM/DqiVRZ4Ld
bNVFeznWL2J7iEVyQ9OTGIqZTvvjuzSTXAb3waUnKPk6Q8Z7ptLYRo5/v9kDh/R4
TM8zv3IrhOd30jqq5b3Arudd0/d8Cm8l7fnaBStGPlj26L6h78QyG4gqUqy7efcV
QJuFhnFNNoN60O4qTcx+i8zSr1h5bp63z524kc4Z1aSqtuGqEjUTBNcwGcjusmLM
JIwPxjdzFvroBZKYze25Us+I/e45Jb/1N+JSwqlolkRWeRuwvT+aDARZZcPTcdjA
GStcC/8LpjqdHb6RymCrXfQRYM8Eq5PI8dSsyKseuVaQC5hdJwdw8l6W+1brzovf
EBCNHMW1QXBWL1QRsfz1Gs7pYbH4o29eK9HIBvLWhAtKmLcR9xlxNMDC+uMo8GEb
bbyaP6xuL2I42pTtbh9ert3omMQeW/IjMGoLxwFA192XEp42diajPq/Umcv+2gGl
R7Flsk4CbJ28ZP8QDdQc8ShFVO6G5ax+RBm31FmY9A1TV/Mgbp5jEz5VjorMQJFd
Vxr4X1LFsGtBiuVAWClnLfWhTdlSat9t6rZOPWl3T+BqBNaeTR7r4tDIHeKSil2r
u5QlohSz6MOYSCcnXMmnxopkb0eDQOiiww84GasVXIAbpT5kyLGp24yGE5Sc31s7
86lEfuQRetczfNh1PmE7hBS/c31rn8IeUy5S3D/+MetOSLdkf45n+a1hVZL2hj5w
18iSmEUw/W3PKCCPpFd5I8QEE9iIU/JQBXabFfoAQY2UXSOj5y3kFhyt38Hgsp+V
zNOob2BI7LK/WAQdgkGb/rSSSAjQY63vjIjwYfUzaYjd6s9eU8C8n5yHqP9Y+4tT
PtAhzE87iW0jfy8XhtoAG+Mfos2ce9MVDNsME/rwYlYZv7X8SpIwPX8tCEMtqnEw
1Nuzy0QFiVEMJq1QdPzamb+tw2lSp5Vn8F9XhpaKqXWEL0pGHSrdM/bLetYDF5n3
sFVzp6ZmfpSZNQXtwgJPaDea3ak1HtsJiAQUAP6p7FUH7HG4KTJn+A9TkPj5t0hz
EChRw/YeBUIDAYQVm4t9ntfoEvyIMkLpI4hw4daZaHT4YCo3XB2edMpMaqUbDh6M
hkU9ovXvF8rLUvw5+/tBhfJXMZNjR8+PaEo8nqnrRuyCTl3hQ6o1yXk616TqtxwM
S0A8vf3o2q77UDHZ5i8uPUzT0BKUFhAij4QUmuPK4tGjgegqbOhHgcBJAhyqzc+7
BN2uO/yiUEqJ9gSNMae+KEoF+zBuuzwtFZ9Y9m8NgID0o+6CsfEjxgK+9G0f5EJM
Vvj5nYHRYpwGpAn7F0ZSIPcx951MtTVsN+INXdeUrDr/7giP5lXD/tb5+Iv8+msv
63Q6pjjurs30UxYm1dT4F3KhO324XEqkdc8ZWvCyY4UCu4FkkKyQcRZHSME/nRTP
7++8QODm2MZ91nKDkmsX43O+KtImWEw8g4o3xgPz+mtIDayfPfX6u8DEi0J2X00j
iGYyICXOQACJMjAHcRhT/JwR5Y2U5VE+qDhwm0LtxUF5GOIzR5Aes8cjp3Bcjytg
7fGzsSVnEEw1JUt1khkQaO2M+7Zb6lOxxdQon7a493/cqRl0gGIAYYaTLplav4BR
dsp17IA59xmM4kGVcscajl18bOR9LOz1anwsSZGkC4aHNHL19vW3SDFCU7ZGyWuY
OyiUanxzQqKBHARkGPkpxvSqM7CKODdh6Xtb8fFt1hXDZ4LEFF4RjEsehvbZhiHQ
XzRRHtnTMr1OMkZiE4xtTB7ntCGGPs+NdLwi3DfZw8joCEG+3u15c/I8Io/MpyJF
0t/5CF1MtkwQ4OX0deXsHp/ouTo+NTlmpxg3nWiH/OMAWJKnMDbqG535RUjDtzEX
3wpmHXY+1xXYspTHZHSrqXRIJmM4ZvZn7ZZtar7/7EQZeNs7w8WB16RWToap6+0Y
x84Xl1Kv7GR62xX3LrL4usgMmwmfBVY2xnpyOC8W1V5RJ1tK2/Hyt7J6WxTiy+sr
jOYT5nCdxqXmd+MNWB6c/ZT2CoRaiw0lyUfPxQO8+/FaBCgINeMkHmWGqF5/+mdQ
O8aDt9AyAKqDQrlOpgoOZ7zp8L9rEPtgUJiOuAjMpGR4XLBP8zNC6Z7FJyWE0dyJ
ZiyULhoXD2Zc8hF3gGmLwGtRs4XYzBOHt1K6VnK2ezYfdu/GeaKMPqOqbFlMz+mh
EmzDXo41eJjMhEi1eAqdxkl6l1iM/OxxyntReuFsYk0/MiXKlKcGJ2uurNftEHoy
W74cmAEoL/oVdeyPgHBscpDe/NRzKwgXGmqokifVmJVeGs8kUncaX89Z21GXcP3M
IBAtDZbET4fTsljjVZQB/rEbXFIkaTUd0LCkDl6rQT3WIG/PjoG5p42HzZohpGDn
5Ddro6p264/XGzAAyZ82pz4OS7lAcoMGGgns5J3JTMo3RELasPNcS37orLPLGc4g
WytoDOlwLGKJGdq6uMC4R8jzvctkYpLDMqzFCiXesfX33rq1BXWtpWqTaVIVcZVp
8dmycVkI3mpQn2ytIUEeEGRXOg9CKwgGIp/WH43Bip9+N7A86AeD92MTAblmSoE6
1s36J5otQzQO0cAx06oXrB5ThMLE+XdXwmbsE1pyxnDj8f2KC8KglYk3pAxclIyo
NZ6BtQuuKv3QSK+24wgp+G3AhsqwIr8OSc2Jo3Ji3PFkc06FgxN5dWz2CvwIJ7xg
keN3skEedc405DdqdY1UHcbeu96Z73JeJYJodUBNhnvgKw5Y79fNRcql7NeMQ1fu
lBb6s7rXu7bkXDsJTgGTY/BBlcSlaw5cakzJybnEufRjqDlHJpGO6879FOnt4OcD
VbMDMDEwYgeBacOW/q+JMJTrQyHhmK82VUNpFDAPYMgr8pbqN9te/LfGJ3IVdiY8
ysxerad+7bx6pUBKIqoFEpnq7KJsVzHHRukh6dysri4hF3z1Z1C4lPsJud4W62ME
Je5vEZd09gFiXC7CGEtJPusy68ON20/qmKyFaz+MwQJPftD7smERUwiVDFDdINsx
TrpUGOR9ckYm+lDI+WLYoupyYFldwc0SPHQzqvIz+/gRbeL3SNC0sHH8Zx6vz4ny
b2qApw7+yRLzU911RDdc8xBMpBTfgHqp4ltXjXMP/kGD69AvR31Ms/NddekrBfDD
BXLFGjkbuu6r6NI28g+7Hj+8aE/0cLJRKZe65gete1qKlTix9qHyjy816ANVHQF0
I1mRrqVelhv7V4vnc08ADg==
`protect END_PROTECTED
