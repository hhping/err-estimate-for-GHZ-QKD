`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sjpbFKIuf8cpOHONVTVql+nhMESJ305tjj2MnacsX2WHFNbIEPaqvjuQyzdZvsYB
ovI74f7ozFO4xJ3Q+nRucsici3+04Rtj4SMOTUZ0YVuHxh+/B+Vlvjef3ZFI1bbU
XhmB7Lc42tXSpN9DxWAR4lkopziqE1W/GDCiJXEjNszS3k7IQ8ZO61xpgYMf5HCv
MdopQp/MNW/QshaBAfJhX2t0acWjjjhtpqDerbUGAmF2kQik+VoLsGZCmT4K/AOI
sNdC27rKoovWNnXiYmSdcLiHu5JkNKc11t0utnjbsdfgwf5kX9M4F5EfMustUD6z
BGcf6DQow6ZoGz4C3ilsS961hNtj/EZNZ8vrF8xpBV+Acad0BhxcAfhh0ESqqv4f
s0pLumDOhB01kTqPuS5WJMBLyOHO2FV5ISxzeGi0umGl8JYG2i4AqlIxu5i/OVfN
dKeKwkhNQs2Zc4XFHJExWN/EzY0WxuzOsPuKNsLlMK0=
`protect END_PROTECTED
