`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fj3s/tX+e8EBL4x4Z8mNDvDvV4yhLOAQ3MuDxHb6BL0BR9X9oJaFlwDz8CIiVDe9
sQfOC5iiLycXEiXIRnLA7kOPlKIetvlXC890kXoPwnPq7va7UuKM6OToC6TYtNz5
F3TIF9Z4kISN6BvJlj4PhiUZQL7MmJp05YPFs3SpNlYW0YRa3LnFqt8+pT9gKBU+
PKaK1Hz6Sb9Fbi8fOqf7QK0y2bI4umeLdI2LEbuVknYpLBm4alTpEuYqMmIfLHiN
0OZHLTv/tOq8AlPqgA88FqjHCObqpR5GYDvfF1Lmf4eHxf3wQyvZIlEuFBtAtfn8
M04yhn4GOKIb8Vier7lmI8yuecefxggfnkAYvZHo2WzMhIywB7N9s+21y2PYLOJt
D0SxSLux88Jx1birXkleKHkCQlP8UQNJhRYjl8gJAyNlty/CiuwSSUxOWkuWm1yX
Hk7Z4uSOC4FM6f74sPx6fFUDPvKoxLT52u3UwuUacXaeNcbul2Wxl9O/QEwUImgZ
5251xzW0fzZyHdjtVJniamsrqPfCUuj4vk0YxrmiHC22Be8H6ERkvDeslOak1zrk
+hKsZUhCUzGry5QKprxXtHViPvxhUprLn4TxdJopUoso1eradzwP9fRL+IZ3dE78
9wEDZVW9bbe5XlHaRFrUUXafbRPoMhw2yp6zjNiJGTN/3Hfex3nfJJd/pIemLBRU
OEpQ7IrYLztbaKoohZv7SMUfEGIRwSiUGVKvrcJJGef/BhEB13E9dDkodFuOjY1t
q47KiYpU0H0cEXMOJty0QgaVbg6CB9uL8yScP4IhwBjgu0do4D1YV4cP8hil+kx9
ES0xOoKG+gJpBTd4I91pZwMYf/ZNss2ume1hXcqVF4YueNWG4ELeVvo0tfSm41af
JM9drwNTQ5Kttas0bZ8UIh8geXKS0wexk2W56iFy8FQGsCleOVSuPPAFPOTswRtR
WBO/4hVQycuF8Znmc+yqTSsdkn4S8WP55pJukKyymP27+SmwrkPWxtnIFaD+rVbt
CNQ4pDOVHSQ68btlWvgs6AJu+TJAIvAaWGXoL8eqF9zz161qbU9rI1RUFlUTguOC
xYwGmJJ5G/HKQY1SuhgMBE/eApsAyGNqyKxMdIbueTaxJT8BEirdVpJ/du7uOGuK
ja46ckqRDz8AUebgwjbv9qMHxPif700Gv0K3hFgmMwodysEDFiwvMJFeFDE/ovsh
`protect END_PROTECTED
