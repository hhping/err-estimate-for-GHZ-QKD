`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yr/rZa6mU9WX3EHNuQA4Sj0D+mCYxQED2P1GIYvHw6kIk5Qsd391nA0gA8f8OIn5
4abAWLoUWd5ZjgnfM0DH/8WoCgcloF1neBJQQqchXTV+A727217o+zvAmN5PQd1l
2Quc1vSNQyQ39JZo9Z7TXai3zZpsnHwlPzc0SByqpPsBtYKWUDhUaJnVhRoqoTFG
9ficC3gEhEKhrArGQpQsht6wMR3uUykatQWOyDXhv3lC3SxrGoWSS6qDC4mnbZ2n
8eSVRzO1hLR8iwyZ/gdDYG+wZ6XoJgeyxIp9zQS6Rywlu7qwvx6ba8MHfAF3xD4T
2rluQVXG0Hd1FFSixkO63YCpI+C+lk/rIMzXVojzoQqofwbJjOvmiEsl/CZugz8S
8oeCn7Z8tLRUqXhiYVYAZxAd2tjTEA7ms12l5bnVwHIDj4IM45M4L+ddinNGdfr0
7uiFEkvOKeAqN52ba8o9cDArGbA/aYoUHX+lzhbyLZgwWkDp4TCij7F7Lgyjei7Z
Fh4mKuM3zkmxRGyHUzPgDxgPZXGgAE8M6xfPCOFM1zAGUB2/iJtyswuo27HqXyKT
L2Xtw7ZFq1EuC8WR5Y2Nh2rXpTIHY39l0YY1ab826fJ2qU39VgjkqnnwX+pFjpIz
HXo5mwJ7JAGaNPtYo24VNMIJkqPL6XW2uEmYzeG2B1egH32VN23T8X1+51anj76A
KBmsRCgToNZKcwzlTtpDjxiaGlpejlcc7mNT//tsdTtdhfA47Lou4XbQz9JcoLEG
AdgbQDX4rqBZlM94+nt8NaRNpkZkUsqzvffN/9m/zX6Hg+EyELxB04Pea7RlG7UH
dWhGnWqUTFL3eKjJUtrxHQsnwZzD2kmuyHAlTFetQvaHXzYcIQdtj0MczC+03AKO
`protect END_PROTECTED
