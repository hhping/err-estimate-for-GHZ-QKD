`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MThhZuEAUCDv2Y29JMKp9qapyt7Qu0ysSQnJynZPckZ2r9PZr8FCe4F4xo1u03Av
apkU5l3UJeDP1SmJm1JzfwpONaHj2hvHPBmuu4NZBAan0DhNIZ8E72YN67uysTQm
PqEoJ41iKyTLcRozIsyR1EgB/gRlBsXVBHDnNX2PoEIkglcMtcu79l0yYsq4UaGi
zrKCpdILNoyt0/99ue9P0UlE+QVIlIFHZ1meflQrP7IKZeRBjBojBMm3woEgls+N
P9fMDUUcCOZhwC9siEWs6q+8hIOANt2jIQFpTOntcDkq4MjrOBk3I8HhesQQOyQ9
Q8EsW/u9OkpuSpFoXLBNqdATuuShSpVCP28vitBFznI28iOU1L+qOl4w2uQdec4f
fLQLorVigEo3bwVjp1gMs524VVBSO7JxbOVch0CJEkZ1fwyHsj/CxkWGB5MC/Dl4
0qnuGvQIHSFG4EXx17sw92Da4oanObhBfPoXiwPvjfWyeyOo0+SwmBF32cxss2By
6q65qTJs6/zT1hN4v+C86dScPIvpe7Cbya7YIwTujmLqJuIY9FwdO+72svCKE7L1
6e102/cSo8wyS185P9QiJFDm8LcDvu6lenWF7K9DYwkZ5wuHwjmkdOqJ2GykFi7M
AV7pAKyH9fQpy+kLi1ehECYXbg1CiovaOg23POIbcNZGeWnI8rz+ykX2J9+PLWBI
4aiKjdBDFK5HT51RwXaw1uqKHDJXqyFIplxTyFj4EWycdr2jqI97XWZGKaxR8jOS
K67PXgglY9KiNbiyfpXMxXT/ty3HNB8gwIvG7VT6PXM2GiPVYl3rRY/+KTIhTwOC
KRc64aDHUSPRYuSP0F/SAO3qVWiwWlJ1siXy3ZGDz2aSPS9gfpE2cgRpdqDyv+NU
PEfLeQJmDq3rsj4SMifX1AQg2Tlht+0GilPEiZMXww3N6Frj9W1Ulqc7RGwtk4AZ
Sz/OE/NxvV8HxnmjBi15OjWMVNRG4phn9peRmqokbyYRop8S6wBWx3BMpjmveI6x
E8dP1J75gkNXJhHBJxckIhOyLomcNgMU/Hvag+cN7aRhTG2CDnlbnNl/PAk9Oucx
gePJeca6YlbfOLH/ydVf/XzElav0kL+uPwc1RT07wFF4ZShkNckC9k82C4ljJTc1
XnIJWToPjMwM939mDp2fSt/DySxmrr/tqjEOr8GWuep4BQteN9MGCvOsL3a9nktw
M92OsFXjbw3MhXNS4MH1U1BG8eCJnYUsWVI+eskLBFNnZBmiFGGaKBu6nYu5Ol3q
U/ZIYIZAxnbDarRCzETUvSMfllA4u2yy60dOTUOhtmAGKJEiJHGfXijGikvJCAUh
C8AU3asrIQDwr+sZCOji3ndqt5S1J3WwNx3qtLdcw6felbfq64VtKFvOzx1XKvT5
S9kZMOpBCMseKXQD2W2849Vu8J/jkNSr7/lIsuBJSAEQYNdTBLB5ebszj5rJhJo0
YonbGnq5hLE6SfC/PhXenhUL9oBkLtWIXwIh7n713boFVD98SVwQd02vLNLUf66b
eF55G0qUd5LIwat+w/gV/UerauM99ybiDFk9doqXv5QqP2X1/wD4gldJ/kjVoylH
PJbRoDFFp/xXkaPDWScqIDRp7Ab2oeCRaWcCQSHIpxG2TP084USr2q/hlOXi2kt6
zGIFMaaO+NjPEU3o5GWou/mOHOU/ah2RIqleFYnSxrq23CWL504Sms4Z6q44GdAB
oTNB+hWdvdBsVqIFKH34F6IzhUwhfcCN2GbX6muVT8bMcqNRa4KM3uE8rkO0+q9X
vCXoFq0WhMMeKITpGK/FFTkmS7lgVFu40h22LMc75jmkoAjr4XbBAUrBUg5WUUXT
eTEjl8RmPPtWDUfiXil6lBlQu3SCmr3YzR1neWJi76e/fkM3rELDnLbrXLtPh8Nv
UmyjqiRCtoDGMLn06GNnaUhNXbB4GH+d8wXZbHGA6hxFOi/VcZiEeyEYPInPp/X5
hNZhpIendw1gd/fZ7IAU8sQuPkOF/qzCifjH4B/SjmDuS3g6jMsBqfh1DyR61D+w
I2ZobsQIQSaD2TzRVuD2sLGqTQNUEj7jhppCwgLuwhcXVIXMHp8U0hgqJv/P11Zs
rGfLCwrSwUSCQvglzbeDr5gYDfZsZONoF0CdxSgRytutvSKa1NeEyaORcEEZ8O1s
tHlgNUuRN39cYO7rbLRlJ1SnyBgiKrCvBn4iFZndYBc1c+GHOEQaKWDuEJFGd0II
VhH47DqC7hEFR8/5+88NlY4kqOsQ5yevcwyM3CIDQ2J3MMR2s6NixlrTD3AFxnZh
44nIFsbTd+a3PXmorHnTXk4/CXInrEceyxADwMpTsYJpZTzWjPCrdXx2SytEWK/k
yWQsQJPa/+ah/XuCD+ob0apXY8edE33LhyQAca6/NkbcThrHWKNgX4kldjHVUCBd
2UwWuZMgwN5FyiSZ9Dt9jm/0tXyTv7aey+KEoAbG3zA/gy8358mdU6BUcHP3GHlt
va6yjAT0V0VGzCDQPjTPCAM4jJejlUTHkUaZg4zZNpx2nD8y22Cjjy6KfPefaJ85
MwrhWXCwMkwavlLW5b4W1N1FjeFAkGkuTrZfDoJAKWmttOSp6S1j8vN3LO1xOgBb
FvgRWPQq3Aq7LMCWdAh2FzUkqfLM+dkxlDpqq0J5wO/uCXrdar4U+V5gHouwkZX0
tvvQD6Z0oDN+WIikDgb+YUf3btZkqx1EjhkHD9p+Dfqg6+Vv/V4QtNNntZQ3DblR
iqMjB+ZybQO/hEq0GHZ3nx9Rjtd7ktMnaalr3buz+AV8O1WL6xmshlGhmd/X0fBV
+mCPvCvuSqwcPSM+m/PB1Nf2h0Z1UQtio8eJt3OZzaYi3E+NJcF15JWUk7c+N1vU
JaJEVLMvrdF4t+nosg4GhCaB95bO9X8XiVGC3pLFH5u2wiulCfp+lHC3Ho1j+tlk
3n0DV24zsc70bJH5nzLifVYrWls2FU3mElnxeZ5QSWSsRFvRgbql8X6WLJ75Qk8s
r2qRDeiZHyVnExulJ5V47xMABLLUvO4F88TGLOhvPfEhSadYVbTf7MBQuKU8p+pP
nCKch1Du/KUIZtEQqOFixfvdRBaX09q0JAmiuCbW2DAWwiNnQ0nz0EPrTFxY4MCF
EbtqYLRi77z6IOaNup5h4HyOOsGG7GRgt2Yf5AK11vGUEdcxKc4DdyQ3cXRPOQba
nj5gywW2cYAI5H8IYhIKzZ5GA+HjaQyew3E1lNyoB6xmqiaW8zhwdW/OUpTDjD8c
HIo5hFY4Wdu7ibHB2kQWFVv9lvKt+L6vu5k1yAIuDRDhmUY6goBswKL/jTBUr6zI
RzxIFrpEfJltoiE/beEw2rpr0IXOq3fBxHUBI/MgdiRDvKJsMKUT2sZ08NFwJMwY
pIrNlfUDervX+imVqfFYMDTwpYaJyGBzrsbz90HxgwApG/AiHE6K961Y4M4CSuSQ
ZpF7r44QSJWDOO6NJZS0E3RhEbTot1QTAYN/w7s/KIFDnzdjYhkSqvK3APbxSvo5
Bilg2GF1HS6ABr/iwvZkEHb/6umBGtrcEi5ZhNJP9eTV6M4P+xrDxdX7YT4lk5qv
pnjwQXNNts0xFAcgWfWBDuk84RtE1JdH2hCKVBdCaVzCZW2ROsnxyyKjuYfjPghS
12YQS35FmCmXscwFT8vgmwtuTWl7ffA+aBXDNvfMEppjEbgGfQbEg/rvCfLiE+Ih
EsV2Dhp+vzMM4gA0rFTa2xjFSF6RlqdZKrwyWjZvoqYfyVQ8UT4eUCndCB091iR4
/fO1DIHdYu9xZceDPF0Eq7BSZHeCZV0Mk6OeWvScfoWjyz3jzSsSx5R69aV3FoHZ
`protect END_PROTECTED
