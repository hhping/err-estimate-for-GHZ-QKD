`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Z1Z5dLzS3W8LSdTC8acuIBdyo+oDUj0ad9Q020dJy29j2hOB6qKZbeoc5d6y3ai
qeBrOX4ZdHFkRLH5HEV9qY5Y7CkIZ16VpsAfJA5SZiR3pJDPAvZaXjS2XshS2D68
wz21zdLxtb82h+xKotbPegbDzytfi+5m3rUvvlU52KbNqopv8lK4eO8xH1ax2Awx
odGJ8wn9824Mf1y8i6jjt1hD2Zlc956KTqgqm954kplY0ApHSSd67SyCcpZgarPb
Jczk4rFi5VBv3NIzOgy6awrb7Ill6aYepGzlSFHgn2IqMZjAPIg05Ih9sXxqF7C8
QIPn3d8xtyW9ZXL2lFCpkNQV/zaU7l0xugY+BrRdaIlz5s9Vfd6Z66ruQ5wVTAK0
NAcyGj8Cs8P5UoA9TGuQn3Yb9U8Qdt9yzGq2OyhD5okoy8TY3fdlQ4V4/aMgJ7Xi
p0TZuYjIMfvZ51/PxMjQJstcZ95X2/mhRH0oUWL2OGSZRZnKik3y/LsnywXmKHy5
Kg4CtKKu1y5FUtwsn1Tj1HsMn/6i24IcLPCILOC/XWuYylFPYhbLTKDaBfe0kS9v
H2juL+7jEWrP4rPeqqLnx7jPFA4W/kJ3ir364nuUq82O6q+LBHIazPKuhTrTxCeQ
Wexw92o1ww+x2TwdR04xbjm6CStIQW/o5YK+E1i2yXS/nkwe9k96O/dFWxDQlypq
vooCZQrcjxsN270AtiRuLRF554tlA0+Na237BuJH/wgCfXvFD5C8qbFsDaSWh97G
2dFueWV5Rf0atx6+UExMMZPxNo+KQg6+EAv9gnnhhp4KKlqqM3z0k3IjqLKPekZO
Y+lWMwpBTTch3h+bKwUZA3EW6pSp0f2Bm/B8icrcoMM=
`protect END_PROTECTED
