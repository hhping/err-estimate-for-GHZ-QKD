`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cal5saFujbM6Jv/rEdhAm5jLTSwjF+sgpOK4HLJCIUbIu0sw9BpyxEZMwKslCrtc
+020ub7LUNiRd1yFllaAKiRan9F7gmjLwrhMSBF8HkNdmvNJnXzO9ySRm1bQ2MF9
GUzfqyspDRwiytmFsnxnocaQkVDTHjtawzlNVkbE2ftRANVbpttf/5yfIJy/vloR
FrV4uuDhj3ozSlciwsdnANcETp8DS90ydeWYfMEtQ1l1iQTgLe9xxCzzZJBsTKMH
5OVHxBIIj6fGNcvu2Hca2G344b+Rq6gB6kcF0+GB15uXDn6WO5NdmRt7ZTtylajB
jGqtAXUf0wYDzYg1nt+Y7LpY/MHj+5mDkm5+yFTtuX8UHm0USKB4JcFzr/KQ84cI
/1oIFv0jz8yCBVfCub6mP9o0+EIVZfBivIFp8SYM9vrNTPnCrD4H24qL3ZIyB5/l
DQHmAWfaCte5bI/whtc9j953Zqib6OBihe0QSjfZ230hqMvYzGprKxC8jqiB5rQd
4d80h/g22GS9b/DvudrLuji7lwxo3VYINverw/ByvetUHAE+k6pqGT1a0PY00nMg
t2ncfwvGwIFb88IZLXslgmHj9B8tqzmVxNFxv+uZTaLmm3uuk03qX5f3Xi2QdAss
DF5OMEkrS/Vlpe5XJxDl8uR0k2QBwcZjNiXu+IXiejJtywxcWcrJ8wzKK+mTzuQZ
8YnHzBq+6laRmFEE+/TiysFDmS7Lntqm3GFQSsTa3LjF5oFrTM+ciHUoctVB5R6N
GaSJNm/1LN17vw01AKvoUw==
`protect END_PROTECTED
