`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2daIeVE68cDg0gGxJbhi2H0sAlUuruo9oywkO/cYE2oOOteSnDzLKmskNx0NiZ5L
QxXncmttWvoOziCEiZyqYb4PUMgu4zfIAnKFWZSO1T+1mPsF9HxHekOqL9v7m77M
9hDwl1JIQSLGDnMpzdoypB6OR+n9pk4nw64AJ5Oi9mGoh+4c+ORtSjQMPq5TXdjT
8+r8+uLtbfO92SQaPHMVlKd+tpxP4KmL50jmDBf1mUBWEtalL/SM6oDi8RE5lG9h
lloNwem58QfCh4UQU4b4MgmBj4hul1LPJvsywyFNXpJnw00givKtZs5S7VMRVme9
S+MJgiNmxafpEUOCMygITneg8a1/kXH5Y5DH62BEDUVXIBAFj+CNsmkD6dcYWhQB
Fu1sDyEObYzwFm4gtgYgmlhc4Cr7YABoT2iiKiD+tmq/IuqO6A9O2hZYVeE1dLSj
qTG3TznJzDyyGh0NVsQKgJ61mhw0e9KCYGYzm2YZBXwXprVN/3X8mCWHycBU26yN
olO+hO9Hq/i4kXDGt2nOFSf68qHCESUaHIa+Nlw4KifYbTvQrvant6ByWtuQafrz
ALzjjwKDSCPFYH1Pbxx8JhtC9ncu53bA4XtEIGxetOV3K58tiiCO1PubgLNSOGrU
nV7Bv0Xyk2xYfRZcBWI4wDU1+LQFq9Jjxww5qgu+CM66S5ziHQx1m3sRWjtqlRNB
rL1zZeg2UbIXdZg45xzEHHj8OAR22T5J+3OG3IzFOY1vq2reRTcoqeMX7mplXoRa
zyW+aJHC/hNoyc7busL3r7pE4N/SwqsHpVXdtE2Y/y+RzJrC9r+8NqwFGCjkaw5h
hPl0o3BbFbWlXgh7perP63BZAnQsOyEWB4cnb5KAHXkRf17EwlvO1ZPbBdb2XxF3
/1UgUEB0oKeNtv+EsNAyvg7Ciz+5YJxDPzvSJ4URZvbW6ab/M9GNb17uwX9iP1QT
lh2mhgsUElNBsnQxW9pEK+DSShh1E6eK4nMhVw9mRw5UybDG1oXqlz08wSzAz8Km
1bBB3kN6+DR/yVlMixwxjB7KVF9W5T3GGebAigCpR4kBuZKZYQijXY3j2WacEMId
I25/Mn1ZdsZNbvTWBKl24X5N17UQxsO2UzLMUgjR9d/wLPpFzcUzuMXU3WDWu2oA
vBsLuG4TtFh3x3wDwMDaGi2HJdzDO8Vp0Nfx4VOiLTN+nnbva+o8zWS7j1MaGMZk
uWtdrg2h2VRP4ZZfQbjr+itIp9q+0lZ2JOp3AGwXz5TPJOJUWXKodpzGmiP0fLfG
ZwuaXtJKjNVsRvldAYl0Qs6SnIZTiNpff1JAry5++yyODqUwE25Pk3u/JVrWqA7O
CRBibBdRnJ0l0fm1YyPi6DaOhV0vPLZKGAyqUjtqn5GG2DIRls8FFKuzsj4r85vA
0cwc+ueqxtpTT0xrHm5xxr2XY2vQUIA1WnvAhsoxNVenqGMbp12CvTSl0kFVPZkr
SRDhH88caSrlPAVZJXOzKipNSSKhw/iceSZ5XBpjuPcoCviG3WEvGjb/lD2Kc8Yo
EMDTXafQfRraTp0UGoJchxsic0X6dGR1xMg5MT5LsR0Gg5N60+qmKeaG6vFnquBU
JjfaVVWaPI9H/vwDG4obLuV1dJgsaWj+xTyiLgkbpL4djuCS30IQVK/l56u/M7AX
pL5IqCIuWpUp8020tf60+vXE5IVaX7h5iYRR+j03jlaLraFK6lEVhUny7FFeKKe/
4jMA1TnUSQXyZwvTDHpScyMKmrwqThiba25HtwzVsc+TsL5KemrXrCw3wOVYA4+2
TMqB/sS0zmoybGl+Rvyxv/n4cVvVo+vU4qumtNZpIVBcbtmt7fH+r4plqEINQuxD
ah6cTvvN1iZ7W9zrOTyzzl7YXIeP/59Qf+KJ8JPvb0R9ivmPYW3cIpnTJGFBb+I4
qy2NInbBgykBOgNe6Gp1A6E4ySK2wPWy6UrQmFEfY2hC+OzrSXdzizA/YydehtA+
1sehPsuwzEkGOH76lHwHBDpd29XtwGAsjPYSAYC4f6r/VF+ZwOswBvTXuiGQp24l
rcJ9Gr3tGvYDtDK36Y/ukNYCJdMHNclvGR3uQFY/dYK0EKVIZPpcxFqcpuTsw2rU
6L3NzwJL57ZjbjvFvqrOGRAphXHES358BdULHSeUh0r33wUhe1spSWDwqd3Fs/kY
+CrOvtIsVCdJji7zYY4wbl6rT993OyaM2lW91JxisWcQrXahjM5VqGAY+Nz8Jv37
Sn+ZX0lA1W8csbn68SFRj33XHzrHWwO8YMy/oFv+pb4=
`protect END_PROTECTED
