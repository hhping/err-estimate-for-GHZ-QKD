`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3UwBwpcTQk9JYprYqzsuld9+Ml7thVPGo3sowTLdJboA1QiMZt+gIbyrJikqDF9N
54AKfcbujOfzZw75HE8/ZqBM86BOl5TQrK5IagoIPj+cJ9dhdDZTq3Wydcv5oScg
slBjx/+YkFnATw1YEPxw1x1pnx6vL/kg+OR2TXQIahjkO37ROkV+o8IsjwpRlHVU
gLKQZR0KvVDzPdiUV2wse2B1OiTIVBLrQw6EKwuSK/dnbWTDl7Ph0BjmjwXEYUEA
G1TTakj1TLDLNH0pwOQsMe2uqYlymMe/4TrExF5cjL0DbiAzjt5KRDoJvjGJQ28R
YGAtvQrJlQ9ZfJQkGD0Ip2tbGG8u8MDhKRyCWI5R+dwshDCB4Medi8IGobSQtPoB
uFvLzVQuooB8tpefoJx803gpmqVB1tEBT8bSfsvFPpiQE7VS/f+bC5Joyk6mD0Bq
u/s6e+9cHrA4FePOwb/G6jTt1JhVaQTgLpT3my3Ta5M3OcBugxsAgmfM/r01GcAK
Zk4R+MlZoc3BcF6DGal5EJClFkUy7g97Qt8rrt1whh6h4Qqa3nuJk7l94N/rAH35
lIgtb64RITY4TUPnekprvmWoQLjh8f5AmYes6zLxGmfkbGoiUbXMx6y1yjedHQvq
ejtLdWMTinWFOt60zIGpxONtLQEN5jtWUhc94WZ1ok52W/so4xA/Mh/kgTyb8C4t
ncI8B5p5d9oM0l58wPBb3rBtLKGuZNmHkp4p13B/sBEnHIYSBfV14sjA/k5m02P+
y8V/gUlTV4WJXbjs3GzDoO4PmsHORAhfKQUCngq0U1TByBvfdpjh34sw8ORxKnKT
kjVA4biqMuKGSE6Urp7JStsbp6LVWC0F8/Uv2bbFdg+j7/Hpo67ac8g6VHo1rK3l
O06j470jmdjvw/3ZsLP3XdBk3RzcPVH+0rB2Veqoi5Rtbe37BPpnaeORJmZ+6VFd
p7FcgEAw9KVg40dY/NheFkv7mG5vEAGqyD2DxJldSoJpRd5FmZXiN18bzOu6k7+h
5FgWRyKnOZMxWVmlk4J4LWYogFr5ITl0nQ+GYHbatOBVMVG2XzjqhA/poCAWAx0u
6EMZSU84lgja4LF0ILFlYcCp6hVlsEpvVConz7Drw0aOQ64oSRAB8vQ0RnRU4D1H
n2TNsJX8NXi8EqPQMrf8Qc/+Ka5aIOyDmHdBkmi2yR2SkDQdEYMFK7Cali4voDQp
6BihX6L+St55tvud4iRV3x2Cpgq8UNVX+TEHi5xzzwfdmcT9AJpfDfuZMgq5akxp
KNjQHzMqc85A3/LvL5HvzWdkf2rTxssvCQGklxDiVKToWS5QPFxkwCZXi6v3PcVh
RSSRhdDpI+uuehhHro/2EKFsBWDD8bEBDY9RvL/XVOTZZiGwr2JzpbvEQDKOWmHJ
dgEDvKKT09T7gb7bTVBXlDsfPXgDxbp8a8taiV8RC4kmpT7moc4/xuzRkrMxD/0P
t+kh4VTsg2kzt8nTgUcDGuueHW+MCARWr/zk9QpVpMmANZosq4colodwkvvVzHRY
k/aTNtz7noPFmEdpOgzT2OtQAgSz3xxhRWL4f/7vyMtj6jyooe34dTZTSw5nBlb/
E9cSCrvkP8aqBuBiBVQrRslXo9K5FiVhA7jbzf93c6C4BpsHjmIm7LdwUjNlXaPo
O89svabRcRasc3bo8G4BUS+0B0X3PkTCnR1zeXBcfHgOzNZeO3vqtbI41kAHwCn0
BElNwHL1olqgoOz5gPQu6Z5I9MPM3pdJJ1mEHxaDIsuFfQGZgVCBXQja09ND+dR+
3z8En+xAdwXXkDWcF2PFtm+2TmAB4825AZmm5Ns0oNyXBj4NhkQc5flmsQEFcV7k
qamta+sugAVHB0PagVgO2wz+T6euxlJFdUp91WG26L/CBmSKu7CJJXN5hbXQz8eZ
WxB6VQhPDnY6WCTzkr/iL8LL18d9QXIcsR6uNpYzW6yGpHvH1JqsQGJvrQeFWGgM
zAS2Sknb/sEhtPlmlGb1dzDifH1dC0tgpD1szp16f8TZbcYEx4LqL5IKV+5XzXYz
+EjMnfB72E84jmqnS8WtDZEJ3QqwP0nQT9xbn2+LgDrJor8hrkrXO7wnJ62wzunZ
NHqc+LfD61zHmKx44y2MdraUYYQutbYmoUljkrVQyqPVzwfo7aVqKVt+ZmTsSMDW
crTjiN92wsSJK2c6UQvB5q02tu+LYvh62EvjUjEDM4a/3v6M3L+haueOWPsKb32a
uWBwo7sXpRBdXlYGvAaxXCda6k3HJSO4kojiWbqssR2+GLkYfwu1RaQvWmCJiWOO
cKDr/HaRaixFgYEG29PCJ2xk9w+FQeMJbIlA8SQGWqyDtt8FwyWrMn9Gw2X1gXXg
Xu0DRkKu5yasJVXXOQPUTvvGUqiYM68F0YoWBFAo6X6zT7MYMIZqimcMNduq7ZaJ
d/6fqAGEoHxfDjgMlpPJxXSWyMSXfuw0mrZUPeCHDdGzp/audZrVyaZoqyLtr9Jc
plW6qDw8dbEgidy/YUQENYR5x2l0QQ+8RZeBESxarOP4Inoj+x3+Zy5AMwxXP196
uEcvj+5odxyd4BS6hq/qvIU4Z7aNgJY+RqOvNdXhIX+l5V1ruCpF59XXSP4+AdVJ
nQvAHWhUOYMth/A0W/I0qOdH6IMKaVjRyzB59wkgRVj8dRkcH6uErHH+Kwb2bmuy
7x/NwHCgbO7ezkZmnUFfbLwlwFd+y6Hqi7Pl28TjTakER2lTNnyufnITmp21cIXA
YvPYBtcrF5ZvKImd7Csl5EksR/oCe7eY4AgmfHg8qspCHvwuWiguIW7tbm7vWqCX
Zz4xVcptsb3aIFQLXyxRo+N5P/zLn7zo8qy3L+/b7DsBJ8uQRBjUSXCCVLfvT9Bz
+9cEdD/wlLXPPkwyN05vaDi0sCYz2i6BNNYxISP3AaKK+oi/Hc/PI+QYnYh7qf3Q
YqkA0wpZKpwwfBrWyWmaUm4xoPS9T+OWYZpdt3WFzqbfF4lJOUnF0RXd6ZnK/AR+
nkP+oQYg4NxaJ6EtU+eX1JsB0HCic8UdTmhJRd+3GK9qGJKpRP6Ev60ebx7BeBmV
+8Wrkl0oaFb0VtV89WEKPFkn/0CK2X4Dy5aBIKlva8qkNG5QetPzimm1vsTSVZIb
E3RojBCW8psSw3oY5jrw87gTh4JkxRqgT9IYUiC+0G6EoiyFBWrP5qNW1dyTFVBk
4f0Y4qCRYspv38nVn8Iyhlkx192UgnIBEkYN/Fbg1qoooDekcQcSqrCSn2CXcVza
hfkcaV6LNRZRGjCxWlyKEfeH3kk2VRqG2YwIp7uQSpOkBxYkcJWCuZa006LbFlgN
IdaSNDyQ5kg+ZRlj/DiPy5P9W0RYkPX4Azws3sG17TWEfegYMQqJ80GsYRtt7Tr5
+62kVY3kb/LwLwE/G27lXpBXXwK1JLAQYNwMgHQ98mt/iV83TWLK8L85bLu9zVjU
l9dfRuQwwGuIf9am1A1dZfGSZVW8aTDOB+gmPGJd36vkwbHF8zb9f44jVkntO/e2
5QU/PSMEjjvPvnKBwOwA+D5bM3U5ldWSj/ZKiPx96aSmq4ikMJIU46EW/SVvn10i
qUk+rd8O5C9/fk0ITGGNgSpinemZ9jpM75nYPSk5sVdekBVQTm8+UR8O7vCDfZME
mZFB/I1Z/VSuBwU5l17jFUskugL0HD1zsiQb1gbYXXx0t2a2mC1kUO6yd64jU638
jQpZ+5aCoSVpIaWI/eyeS/OSQaK33avLu0ILEVnp7N2N57tHCaDFz70jfT6LpdfR
8j/XuSYonGInw6EgwuSHNtnCdGoMM9sMHj05wTqzXzrQwWEbbCoaLrvhBWk7ZHAV
00PyYARHNOK9NU1f+57K/sC3GWG6iSNi2szEt5NFKlv6RdEjx+JpytUn8L23tQPA
f0cl7UB7AWchGPJwUYK8eElzHAlyoRQLvMRat7kuXQAIAKxgDHO3nxotIEHHFSfU
5dXN4DbV9Wc0o3rmDHXQDlX7hrmXh0Q3OmapIslveCZ+1dJhQCBxVbXgGE+LEcQN
5a0EucApa74R91wN0zxkJ02JE85W9q77OB23WXtsDFozbHori2phhMojT8jWDaf+
`protect END_PROTECTED
