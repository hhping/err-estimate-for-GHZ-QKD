`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
puKKV5o5knTijIOqyECVNFZcHrmYHHXeRozb14j37e0FmEZa4sOy0vHBFegRSnVh
SJHVR46nWmxWKOjphPbdFLJNKSOywpOu4x75/FOesYUyKcjbGRwdHS0rz+wsBWIT
HPrUP7sqUdTIc5k0ey3Z+vQCfqCiVlWDvF92PQMSeRZ44ad60xYw1zGHRsYLIde5
Ksf8+YpH9dEynBwmAV6+GARbppxj76cwAlCWj6UNpZCW5H1r3AUNMlf1wy0Fg6qk
bNgB18mLGaqGrFaZ1XNJv0PXMe+elx+De67r8ASt2OXT+9VudoWjyAdayv2/bt/r
1W8JlgB4MoAjiZsF6W4uv8E31XIBkGbKNkoqA1Vogn5nd/mm+vH+ej1VJKdP/7EI
fGOqZOXCIkmrPPJegmXFtEGIp1hxnVjOx+lUBp4nB25wPNFAae+j+PCP+RPrY4pE
EBfDqqL8u/2wsh6qall42QYWU4ZT3XRCpUySPLhvOeo+GJ2RydpG+4HA9grDBF7s
mihrCql7Q2B29eQvxPwChbJ1Urm6T09NGgvO0sZWHZAAXMpIbLHdJ1f2m06G6iVx
SbNLVsAjUz9M1XM9l1gFAzXoiKYfB7i6rT3CcvFdqGzVXD4efxbxof1qDHwCpK4v
cvp6OR/DnENcavcbw218YnEOHadFGOIBgpA6RHxMF4YNFtk67M8VLWuVLomTE+RF
5aac2ODDbVPdNlKFNMJ6NU1D/Ld61fa9Z/cS/QQzh3Axa+0VeWo+QwOCKoAan/6u
hvI1bgyqr3/W1dDKj+DDfrdhWS0cqX55G1HrWoSLXXkzKAibCFbq/UBvHZk197ff
/1SJhwfoCVB0Zisne75nZ75C6rX9aNh4pBrSJ9kgoZitNk18ts49SiLOVSzoUIJH
Tr8KQozbWcQGRtoqzPUmjqVwdAf+sixZAQRsjyBXbpzD7ZGKP6Ah8q4wOzIC8pH0
GUfQpEXJ6N6fMCpQidZRTpDIjx4gAZbuy+qoTFc9AivumdbVdU6UNYxts0+waR7H
F+0s3b+FYApSFUbh7hy9mVkuDQNg4KhIyvhErdgWfvc+QDgjSGhuHc6yukdVGyHv
BiWiEmdYl7yDMbT+eyoKruOlTlGpvEutqHv5rVX5vTGAbQNJ/0Y7Hsg1WEHElA+y
z4jbdLthyUZiR4dBGCDeZThhNpu9RwhryfQqK7e00lIxVQRMG75fdPmV2oUhtj60
lWYEf2GZvB7EVtkoN+TPtdmmpzze8l/midl33NCc961LKgr+zr2z6uWVj3LF4u0y
szfkFobJ7V2Zj/reh66Fe7IFTNqujsMy2z9pzA/iMY6j2DOwC9a0vTknCzjrHgq7
WQQpZkVg3my3YNMa8vF/I+1463SecpCW0A7VHpZvYJ9nnnxA1kCQ8/U0TfmbeE0D
rYtXx+Q6iOr6d5u1t+R0YANWGyOjdmCXEjpJ2CkyljaZeguT8gOQMkRDt1bOHIlP
3yXt6GAoIo2K2w36aBDmmcbezKw/A8WgmSRCNX9wTNUJIg3EBK+ki3qdoiFRpfto
gQT0XJnMHF+P0yjKUR1ZvoHRQCUFtyz08r8A1NSj8WIiVBdNmFzwGmN5zLPdRIy8
h/RSUCUtISrBV+teU9jfTIXrk/cQUXYLaseIndl4mJUv8jihpQD+iZJ3EzOuqb51
YIB0jYcLcbpOO8aWJ4RvZFu4/H0d1HI15VS/6XcDxQmjyTiUu31vSmuA/Ya+pPdQ
VwaWPe0OmN0Xsw6TeXwlpqIgSr++hJ1JsTSbVRIKlmURoA5JxVwJ4R8bJOUQXjqn
e+q1NqYM56yJOIE99nwXaCKHfk1KgJd4oUrhSIw/H9ksjsWn8hlhyR+Dd5keGyvk
FC/9wEUQaHXlEJr3+O0FjioJcag79bjd56eiX4fQxA6WSWlr7FpgDzJKUT9z5zV2
RPdKsL57jAru2/7b34Sxd91m0yeVeD/Nldfl6+svMGzgK2mFnCPtmpkj5gLr0JNe
9e9Rha3cL6XpD/HH92ZIQExb/+3RdmLSjsvl2xPTAsIybCJje6MOT7UwbS+6+8Oe
NFv5pp2kUJZiDTMAvB5cdCnY/gSbi6lLR7twMnOY1UFCBh2I44DOEdDDimoH9Tj7
StXQJr/H+skVbwmeGulQx6RCJq1o1y/rpoE1bI5FDhbnHV/4EhyIoeZ3y1SiKXsw
o/+k+/sThVPmwne81I8HfdYSzR9lJFCcEfIyLoalWk0MhNjc3k+IFl3bvy/AnQlm
6HuHltDlRT6nv2TKzPB29SwdAgomAyR3GSwQp+w1DVGp9W8dqU/qKuAXpvQJvpPb
RPMeLlAN2GghXSmRUdXGcyYKiKGO4XZT0SPoYIkNixccBnwGQhf1vohG5xZ8qdgE
CrJh2bMxNkQiZEpqAAFrUoTV7GTL5YbXiNyuKTYqI5y5HHtcCYgPTVaXu+d64iGJ
mG40VimxnU6DUiZfB4KtQE9/btBxq/w6K4CWjkDPaAPPzI1fOsKttMtsuSPbtTC+
2wRquoVxOmn7pwcnbLkTfzjX52cNd8W2aF+tvL5/b5Fc3ZKioU7//r4Re7bSBOLv
vmZf3MTnOXRidlihnTnYPO9QYZGgiNp+w/5sMji2ydqvL0xxTqBC8gpo2y/PO0lH
V4DPI+lZAuvnEMt2Bw9F3R2+kv23kaXt35/77BqUeBWCM4Dkklcz8dD5H+IWwkof
aGRojtDLco0zFw7tKCwtEm+fw5VU5PbEtQ/nRxHYVhY6n6bfyNIdy7eIyUO41eUZ
0/ADvedo0OEyIqSTMK+9a6g5os/iw0KnA/AXWYuSp/O8q3nU0RhY7WCsI4iG+nXF
EwsV1z98YDh+7GATx16hntjtFibnI7T+n6xnknb0KoPgR5oSEK43vdjvFCzk8AUw
jRL6yyBTL6n9/xSfCvEQdzcSd67c/3XApfsuXSRP94pGUuJn0Dw3qN2g+mjU7Rqi
ExF8y7NeN9NCCGlPk6GmQXmm1Prx0rBazh611We9aIyghJz64+Cby4Ui0B+tu+KA
YT/4t7vIZrbkUW+LzA/WwDsNOlQmzLN45Sq8b3aDNZeZcxdWws3Py4xhAbxVOzzG
6OF/xY1eheg4wWOGc3uW5JhdKCGJMyQiWZ/okOddmFuPRaOXfu4FRvkbYTGNdeZc
c46BlysthYpYyNwWwG4n9X/shiWAqStmy69I1ljbqTx2ofTIRearxy6uKneJoGdL
6Ibxj/4HXRM5Hn90lfK00IFZ+jV3DHUtT3h3cV+P/6GUCfueD4KYNuYyGPYs7vjt
P5PsIoUet2quz1WyRyt7/Q==
`protect END_PROTECTED
