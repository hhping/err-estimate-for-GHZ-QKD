`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YsyJeqd5huj3bySobZJ5wkTk6v63DKiMaCqezviDT5xVrZcQe81Aqdcqh22dRlpr
LrnNf9O3r++nAb2V+9kQ1Be+penXNSpVaYflK4cTf1UPG7artbLPenUYunlBXEzw
TjeZ+cg3WdnBOLdtmsZ1gtQtBXf/1RbDZ5HlZYnSAf2FjYiYUIwqiNXZ2kC1QhNN
aVXp80znyWLmwhIZhriKT0HZYQ/SXT6CJCdTyXKP/yYbyoPIjmyTorREV+9v4h4y
88yDw0OKKQEKkur9R0iDZzSrE/uNs9K0qrQHiCDfPzEdksbkIVFgig8N+41NLxQy
+srtIXCycE83IZ4aCNfGgAqOpR3vbBSFI/guO6qXAd35m+BJlemN8pSMbOLuCwpn
q9LRb5fXiJmy046yMy2bugeAvimXmfHcraRzhoc5fUcbvvGYVTFxNVB5N6hKFACc
YGZqNmTURTkMdbVN7HaaGuSci7krTGyNA9AEmPySM/c1tcGpfJFyhoe2r9WxntdK
rt4qhd3hnuf8RVfgpQG1n5kiMQQTrgWMdnJitQ8wm6x8TydJFSTGeArwjP9fwMmJ
RwN22lsYxMdkcC+7F8ZWIguBTZ8/gL9pzzYlQRYTs3qaISQ3dn37MfsEkgUM6+vj
yfe2RLHNWd+VKrO+CB+pjUy1fsrps8oUVOCbRTdbPIhlGmaEk0O2ymQx1/74tdCY
uR9zilaaBIrJv18OWb7RRPWE2PGnCARBsfY0o3ju6mmeDM9bebCEFXEAB+FEL25S
TPciCg70wsWzvuZPLU2mq41K4hDsdsVauD4x02r6Lz42QTXrhqH8M71ZsGr54VMK
BIaRsT/m+iEBdvCbk0AGaYTCuKaJ+UyflcbtAw89yHD6icYeY4pbA2Wdg93rOVtn
YMrPaQ6nGfQlLaWxrt0f23WP+7qo86ayw/IHlY4xA9GpHROezxRYJErU+lGryEyW
QAXFsC+LubV2A2sq5d3mCOb3aGce2BZmF6mzPI+z2IJ+q6f7q/lXV88SMw3YsB7n
Bf5NaB/NNDkB5T7NAQwhj1bdY/Jv9yqz1nQl8qgy7QeTZ4plz+wZQcx9MkBX6Pzq
VFApZFJl8ENn3CSiAyJ+ElBwVHalmRAAkC0eFDJhOmXoUT5W0OquZKG3B7xnXEst
BapSvDNKvMmCU52P0GwRgD25vgYdwBPTWX/IGdFhDEB72vMM+4IPQphi2MSHx1e3
3O19GE6cStzb12cji7eZwqlcTnstDFhmAsiOQkqNIh3Yk3bFBWFmRKgUDsBAtnW5
stMUUATvTopD4bHtL1ZON1/a1KScApBBz2trIfZ59O709U5KkRevMHrzoPlitA2Y
C0LuooJQbe8hIsYRohCD3A/s4SfFltdNrOrErDFy7Oky27j+i8Ya3i+UwuHzWBDA
hV+dkK55BXoOdaWzZKEoUSkEJPJwPEOXF4onMgSh6N2VIInphzInuZ1EIxOjLfME
p/tqguEijHTUWGhHBtvh6l077A1g3tDLWpz/nObnsGbaU8yDxL5ZsTLYEnKLeohN
Mi1fFq0kMNkz2mHANCTGU7q0DnAJF2VdnqOHVtkacSygCznsc3zvkb9wPAg7RiiV
qoZRqYEBYNn4y5PzWE/BUbskyv5iCgz+A7IUphN2slVg6KUKAjF7kQ+UGBHDU81/
nuPqNpsHwETQ1R8TRfZMOpIjbxdIBJQV7BuZQQ5TATptEoVRNvkW86OI7/GNlqeF
0F7gXjeQe7smT72PNPVXRuJVOLjXjvJ5VXQFbsdMa6TLRAT/ADYDzQhtxpMeXGAH
A7LeH7Ye399LPR5XyFq76xQfOIH9rniuApLr0+gRwcV3P8yZm3jYYYKKE4Flf+76
pHXtIX/7KCVEL7Myq9VUn35AceyP6dgSU3/iMKDAXYWcCiVxm5zHyNs4e06LdRhC
9E5vLUXyuCcvCJD8gw6/P38/FSpLd31mvJ06Dcw2p3zBD6oDLl4hnIv4m81tiQNU
uyZTIqEW7RGpCFrjBDpbYgaovORnmUHVyNBxtR8g7eucMsYAnB8QNbmse5AF24P7
m69QzdkHLz8G+IB+w99Pb7SKt/BWkLhEUmOtAzKPwJSX5AmJDjPAhHOYApa8nq0N
ElZN5lT8TRiJiZZyMa+QbFs58rbqImHoihHRGYW/NjTD587TFbav/NEVUVjFWqiA
sID5oVlZyFjT6sWbWzDVI0oikuyBQnm0Nd2zFQp+84JYQK1yuN3yUTbNWGcxn87w
LNLKiTDCwwzhHwNx2cyU76EqeF24+aj+iuZlAluAedTwjdJ8DNhvTsPviLN5DVmp
5W+u/1SKRNnvs7gEY9LqbogmlK9VgPVxYKCZ5EYUJ+yeCAtp47jkMWAwr+bw0Gx0
nsCZRAC9V6P8dYCDomdGbeLqNkmnwh0yg17u9zsNtdubfgMMyIjWw7+biZqLWRHj
L134NgHDa+zxFwDPaSRe3cwNmTOSRdZ9HJvaqtywWKkJim7nV8ptMpmAvoFPfqb3
6FDJfQRxpiwELn6dXZn7M8RaGKblLpUmy7AHeClep5tK4HrdT0Q+Yw4oxvwxalFw
7oxxm4DdU2A86NIBojXFMutVNni5EbVaYTBDOjJidCKwPICaJoiXHelq9vHkY3GU
qhRtm5bBJ+OwTYUSBgXRGouP78R6sppTt72SGAmRfDxAxQnqfi9nFxj/qjVHvp2u
xLNhOy317OeCwGITummm0mwl6hju/0O6QmODpNL+I5+FkMgjhbPT6DxirpwDfZhR
TTRwJTsBfGo9LEM+/CwCmJZl2JYjJqvP9eUWtj8wKhjWSMWTPG+FyOKToD9b6WWB
JaTbXYgdHpAbjoX0BjSoOlAnz39nwe7SPMQiHWOvEtYCZO1SVvvldAcgd+Iabq5q
JOCO2c1LcF2ra2n5+ZFYFiiIZYlcMzkKCiPkqDw2v4HQ+dIYLR1ODz/dK27jSBMI
S6peMLXOy19PIa/DZ7ECl/PXEB+ver+pi2D4hPZm4EOKq9wJHMkWRpPzG8cKpbzg
ieOiXB60W91f5CvCTDLoNmypyVkCa7likDcxwA1Tl9DrIERNsFy3kFRShLZd69xb
DJr/pJsmNvjFlDqC12S3uDu2tO8q1JYAwtxM0/c2foePpCyg7jB6vYpwYQk53b9o
uXWXb0buvonsoLbcwUF1LURzzJiPxE0J6VTJlfzPsFs=
`protect END_PROTECTED
