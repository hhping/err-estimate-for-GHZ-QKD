`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uva3iwnXAGhJCS9opHostKlSHfHUvu5cxznwNtV61cb79raFa11+J6kKZCWe38Ek
TslBnlCwYTYfIvXvdqDAQ83Z+VOAqxt9odOwLjGKU2r/+FVdI0JcyUPdFN/k6y16
cxUxOy56xW7Vj6B/m+mlJVvMbhah1XcCUe+D2qcUN7JIzMKPQf08/drbUU8/XC+r
OcoMoIGR4T1y19SFKzt+rQVaOCCz22R7v8VOX0zkKezVYt+wMaIheu4Ms4vWiUch
QG86QkvHfK8lpUVnOOhb6eByT4D0t47JX4dAfp+u8KtIDlHvfGPZfVwbLWXiTNRZ
3VUjLEYNxS1uJ+vePuFUKBkEdNbY54WfWUi/e1LZQvxgJ0NBDpqN4f35QbFAZJ9y
P/gN75sx0HY1i1JP1jxBvOqE7nuj9lcGlUN4jDIAx5DohWe4Vk2UbuzjJDiGjdxs
B/UVrpIYVJUunobNZS75dxxWqHglxRxHrvaUjVyC+9OadrvK5izkgmt0gHTx9Fya
3Pq51KA5u+eYNoC6psOTvhBIUVyZyzF2PcwRJqbK+USRaQ+DwyVWEEYHF+qVdGul
rP2OGYr9u2BpgvUPoiWMepeLHkovt02aDlFKFRcxZ34NlZBMNATv2AVBqHgxaL0p
eO/Fqz9ALNX97g2B03UB+acmGS00sQmZUMLjmy2uVlw=
`protect END_PROTECTED
