`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
10lAH4iO79dHeTJDQcta4huteMDkNlQ2uC8fv6Kb4MmJ81hcI3ZspfsNc7Y00ciJ
jW7oUEbJz7p6Y2TQYWeQio7czYgun2rgUhrboDCnvcb8cFq5r+GJC8CVf0Dghg0H
t0114DdQ76nzY/w/YB461+FUWn5yisjcL8oASIfRb7TSqFqmGOuZUyjpEOdrxazq
yFGfImmueQK9flpG/h9QpXxcwaaHVNhgYKnmD+gOD3dcX8yrUxJnhhf6L4ozktTA
Z+fampyhEFL6kzLNGB+sXOLyq64VlhA/pK3zDd3qaDZjVJqjf6Zf794fjTDnWq1Y
OfUuNNUfj6Oe+gk4BQ5VcRYMGQulridS2IhCAyOFXcbfAtQSh6w6Y2KmQz/4IZRY
/he6+EKFHlulvkYKUCLP0WQbHaXyBphDt7mQtg90De9mpvYJ6RWL2pXpfnZ6GGgo
ZWWgRsDMnjX0GsTj3FodckO1tN04EpfM1G7qaIGSX+sNXCz4pAGVFfQxC/WXdpR9
`protect END_PROTECTED
