`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AoxY2Fq/XxA79Agug81xVfnFb7LyJPRZf/S5UJTwdkiBcwYqJzrRZm/eLtwjbArP
Wnfo5hHk1XaIekJa5aDjh2MW2HvxqK6d08ZFS6LoPa6K2U72pWaFD0Hh+E2jdA1K
BKMptlUzxGEVBp8ExTO5q+KtTZvS1A1wRvCZg3WCh+t0RXHxtIDqLZrTwXDxumQD
f9d4FuaR1S9MM66Czh3yuH02mEQaTdZPPndcY8NOn68NK5EuVxxZyS/nF0kzhipo
W1g1fz0QHFXzgmG4r4nN3GSencyypOTClFdv1xFd8acOGFluJiqnb1mmKaFGQJ+9
BxunP+nBelybSiT1geyZpxHMmpGe0VmMqzLPDyqMOWTyPrsyBYSrz1DCemHaGAz5
BrdcxM1F/t+1Qz1NEKZ9BzqSJYd7IDM/rFbwQBqj2qER7FHIvJ3ErFyVu2fzD0D/
FryhrNXRDpuvhmJP4rmmwEZ9mYshdpmUSApp9JDa1iMKA5Q8C6mZ8b3plTuEOW8l
J4qhYqK1txc4eIr+yg5N116y9UWn/Uy+/N6fLWgN8G1yVE4Q4YwYZJfDC6pyN38c
TZQdBTEPnd4q9zPMwmkhZA==
`protect END_PROTECTED
