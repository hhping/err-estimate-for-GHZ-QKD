`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q48g4kqhdPnfjSYPhzJb7Ad2URs+ct+j9lvI1wpCiHLfeXg98DGKBgE+5VcyDonK
7Q5njSiZIENllnOV3WaEvybBPvklvXED9iN4UoVgRUCfE7BZ7CfiT1o4UK+EYkgm
tRX2dHl/4+Q8wdimpbpQJ0aC5cwcZNLB1jCW5LOVypkXjlMVIbIgdlKm+yxQ/m1y
LxLm6ojP9zYr7dHIypxD/fbyOJKKsJCiUx1jm6kwD9BY5TNKEJoRrH44gvgkyUO/
8PgbQpf7QSDhmxq++oAvrSUH1KWHZJVOhiD9i/4RhxmtW/3zj3oCOMtGxbLZYW8D
Q4qn9l1tfQixi5rS1uzDg6khKAknkVnUN2n4WVL4uYbIRuLFf1jDV3dvRRiNfMgk
1WoqvkVHZhSGq91kh2aJLqyAlZzCv/rg12IefzN1ncrnX5jqR5/FGpIHCdqd9qZW
PKaQrFhHdY7PWYox2R7NtTqNPmi5d2dlbRNoTSAlB0tuV+n3UNkmd3yr6PL/xIVn
`protect END_PROTECTED
