`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QmPba9ZnEcuuxb03tJrC17TSAf8Zvt+gw/ljQkvqunqdwe4FqrTxu/55Pfp7HlHX
cQoYyVnrXz2so027ry0u7BGw7J9CJpjVobVtBHPy0wx2T6+DHva7mVYrXcbPKqEt
o+Vvqmxbni6F8A1t9mnEUW+MNM2WzK5GZZVwwu87InRrIeyqfeCM7uzz5K68szdK
XNkhf+/IndHAF6F62sppi+vs6qRRfN06CP128cvZzG8tZn8ce91sV81rjOvy/2V2
z3RGLfxoQVvr9rvKmqX3ym4Hun+3PMj2c9nsZE8oJBxM2CO+QNwRMKsDtUGxpOKL
1Pn9zcSaF75/9wRA6dbNU2XU+4qYvXQdbvstXQVB79cqtoVuGexDmY05FmYIk/Bk
QwDfS5nOvtuXXgcVR24H7OhRX9K+GBQtuABYg3+wZz+MuvCY7qHDuYad+NsFPjYP
79Y4L/Yp2+otUjZ/e1u/SwBvJ2WMGxKdFd/xrFmj2mQ=
`protect END_PROTECTED
