`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+taihgOjE94sKm35YiEKZ1m0RCHcVex22v5FJ6+7dwn2F9MRhB+xZaUYDezMd8DV
noPVNonW5r9i01tolouYySBcJQ6fLxDWrU9uFdltqMk1va9VFSSR3brAbDyV8ogh
J4zunHBSdidPBpNHt3dMczUwxiLXmWbaeFbinS7WTk3AmK1mhFWEdwqSREhhD8By
eYjt9zPk1jmhhcqbimAdsLvk4D+zxGJxu7x0uzWdDMuvEc0OEEPuXFB/Aqdld9gY
7Ohhy3gnrEtzSAPUzH4CH0KBtOQtOf2ZCkY3kUHb1OB/XGd6yrRnG0BHnnPg/Xni
CxN9PA3Vu9WPdGQ72IpBb6BzyOZXjVHX9NcubjNxXAGmxWkudlqdN8eMQY7MLqkE
QjKlTqmVzdid1UnNF6f6jYjy+tvocwNVx7sfarZ3KeLkJEkoLWNsivFcyXEqPe53
Dgq2TfQWdWPkYFNuX+LjGfU9BfSaHJFEKNNbFY569p7MLi85O+ZUCaYj7HNjmWFI
JqR/FL0PGBpbVzdmYr7PsDDg02i69z6eOkFi91k702gTv13dnj56EFvZt/sZ6qyG
ikS9ya5Qqrivzpy01RrWct7/m2kiXk2OL7bG/1ndg3jZT7D75UIRW8H5ZjcfMPEj
nF81HNzsl/MmKdc2WhlDlY3MRLybcH7H8kcv7V7uRjSbGq1rbSQB5zdueKXy/29q
fq3Ib67MA8yAG3VjvJ2UqSmzIT+jOjeetCmIul2aXiTNYtlybezEeHZq1ejVWRGv
5dVep/TTr5HGZh+Qyv/s0zUmEI8nO3WrJfjW5JZPllBFxVeN68hd3db4/EwkE/Uo
++tE+TrikPIyKpbIZ0SQ0/POGcV7XKJKPSFG8KOpXH5koUwJf+uKROefM44vwXFt
/qLBxHrw7yxhgg2KTfAb/NTL+gBND3AFojXDDOCZLiVmzrUdndixp8W/9VJz8ogX
3OD7dZXKsMMvELBcy9FK3mjnd5rfKXjYv5I/SGmW0kMi9h4Vrsaox2O1UGOckssN
y5on123yFpurN/y4ai+SD4pnhkheIdGEYnY32DTt93BVK2g7q6xDyh90r4q/RVLW
qoe23460T1p1Fp2qgbURpi8UvQoqVoJaSvY2mRvOFKKJvNzNqAI61MZVWxrynREW
nYGGLzPNuyItnYkvaDwG4gstpm+J38Ly8tWRgDATA3EwLVqNER8U725oXrCEKPgx
C5t8H9qhiIG7BWAkBKjrmNDNZ0YBiX9EyxfiiESVc/ljYY8NDPZQblvx+qvRIraa
ipcB4bdMglos3cEAfJOW3/4Dq46ci7pGqT9PK+PhMVX06wgSL0zYz89ZRGkCikip
6RqOvNF9Q3cDmbYucn0/6CpJH8sv3KEUOK2bTgcIskzYsfcCXW9lU/PlKk03KEMd
qIUNfRgv0DLvAM6oI4HQO+E0szDgCnGThQLLDKlr6a0qc9qzWG5LAwStoYNiSymu
2w5yqOWfxw+kM7wPDQsXhz2ZmuSGJxdu8QmsJhqnrwT9FGYlOsyrH4tRDzrNAgtD
2D+pjMTjnNKoNYqjDYhkUhJb+61SRtSbYf4k9GOJsIcHfHMP30/sPMz14oyi/8B+
9jOC8sC0iX9vW0Yc5HzDIp9eJr2524JvEgmInxfvNlJI1j+CROb/M2N3i4cCl+lV
wLNDwktWMivmbTYzFoOTWq++GAY1CX9hqsEzxBPclzuLm4Z42s7P9bHn6Uaq1yhx
rRAx6+pyEFPUbx+vHZbPO9Hae/0DKkCtWwOkrJGTmHAU1vBINKqYkSzUUOYtRxI7
afghsJSvWfZXIR6/aNRZIa0+pQxnMbtQkcWxDuj2cReMgX6LXWw6J9gkN+Hqlq2k
f7t49Lt88OQ2+R1qh8GaCGmP/nesHVsRYMf9kTY+c3fraI8oY0vNZfqYoTspr2KE
zzmqtkR8qowT26F5xbd1NJUQynP1GFqg5hUT9JqK4zU9lFwCQoe2dqu6jHDqWB8X
C1rYdrKxsZw/koxFzTqVv+TGdopC2FjttDtxCmMpmaVvhVtoDHIJ4Qq0Q6cHhZJm
UVA3tIxnM3LSyP4DQnXH4Q==
`protect END_PROTECTED
