`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7VN0KK1HDjpYlngoPOc2HCsW4t5PslfQd/CsDP+HHHXUujK3KcneeiYgypQrZTuN
n2pFmbaUGfZdGjoa/J1+FAayci4wCfKEl9jFXPyhxOmHhLA/c/WRZXTOVbRH1iOG
kRRWKJjFUDKUcwc8XonvmghQ5rVGGy075WrVqBDvvjYPYB7I6QB9f3iMBBDgSx/k
JqFtigvp0/i/zqJFRxAB6nQcua9061SVO5yvPhR62G/Z9Cxq634sP4YIX1f/Rjfc
VDpdyAA3dvIPpDjWkp7EXbRTIDieJ/IvcxjGN5dYvRvDaBXsVAL6tppQEcXVMaL1
o0tMk4g6LqBYQct2EFkpTUYaPP/bedATB1CNzxz7faetKRBwEu4+amhSaxQKL2/B
mzhZeOY1vHiXlU3CMHcP2QE3yC1qmSmz0asAAbOCbUlZJLDhuVjN/U/qW0RLfdOi
1Q7LwlHB2fjGdaDGg5hrQPZfMw3ViUrhIZzmQBSFbZR+pNDp0/2gcV8d//4nT86b
AjUFmMEHbgLvH9ONR/Hsyf+LveeE8IFf+LiFpRmgE43ZSweMWEmU+6eoXWyRV0BX
Zihg5TNB05loEqaC9OIu2KBJeguBQKAQTb12HnNov9NFWRYX3T0qDQXIOpPySvgv
UtqStq2xWll5q7Pi3jtGsWuFifM2gibX32RPfH5fSONhz6cynbXrWnmRsl34MXJB
4tLO2u4F3kchY9aBiwWk24I5UJ68QhYm61e4quf+MM0fmZY6+BOy1NpiIoWyUhkh
xsipSNnmvOjiaF/jii2sQmn4zdJbX8pnlUBjiZRzokIKs7riegea9tld/PQXOCnk
7/F26AHEgAm2KC1Z3ADmeJW0jYUuuOSErwgRbiHNqJYknljUOdAmBCR0TQLRExmb
E2Tcxu2zS5yQtFf3ICyCjMgp/n3VFZBFffgBEfttcchb+68XkiUiZFgdYZWgFmNy
Ypot2SJ28womwbgzSKTvNwrM30pglqhX4ZdeiIDRcuw0OR1XYcnoS2hO7Yvsbdfz
QHQV1TgQHPs5gDkM0scb9lSy1AJnsDq0cYO/gQg6yAk/J33D8kPy/cdoVdI4PH34
8kbzYUCgqhpvImHcUBklwL/c33SwdO+eXAZ0xwDdEFUglJMrfvE7upi2NMGyqMKU
yzl6r/YaZmQezUxXS+W/4qSwmP7mVFE5LI04/bLT5hjzkDcus6+emt4r1WZhGS2g
axmxJfbbZ5Cgkb/7rwHdZW0YyoWtz2uq3Y55AOSAW9M+Jax/o9WNP35VCFwkRDgK
Q19Ii6JA7RwZu3qOTrxX3HF254yAUhcnVRYBa6s8t2ct/RWl5LzxiY1TxehYQQTI
DEqb+le+QHBpAf/usQrRPnJJJwe8Qb2nAZmv4Pk8Cszj+Daiqn9ub0QYd99iUbeY
XSMcwQQKp3Kcv4bnb4KOuZKqLWsTdApepuOrUn4WtPeZiCI60gBTLzQ53YwrI1Yo
DdwF4y9H0Dw5XGaTfCLRkbZG1/mgHFOz6uRdYpTd2MO2qAanyo7dkn0n0XOAq6L/
XLkCNttxwO2Q5yyAgaAkrROCgjtRL+Lx90Iwq0D/L7wqPmWZsu7WQwNUrRJTp8eH
2M5kxLVURccXYxJrWLwGSoy2JP0HV5ygSo78ltnHnCS/xf8NkG1bcCFMHYxfHia/
TQDC2V3clXrvrJqvFdWTNeb/6UGMbnZaw8m+moPiAEV9lzGu6C3oAthSLS30Ou1j
ysXn6Y316/C2lPRsGmerMh542qS26Bi7NS3TLrRGQoWBGIscZIS6YKNtbPfeTEIe
`protect END_PROTECTED
