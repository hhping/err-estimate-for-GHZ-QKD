`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
67nXzJx6R23HWqBOkPQYLVWC5ybVMarFAmpG1puFUOpxLONfbm3x42tbkDQR2C2m
XnArPSrOYwADu86PXfvSXmb2+zTX23baS+3XvOTpejHHdYNcfxGSf4U4ahf/YbPM
bOFTVhITty/KhrIZnpwmxvwrHHP1B7UsVIJaV2Xt7521JveL/czjcCGYd/Cgu7/5
4HL4oA173cV0QsT8AP967h55CnX969WZYckmG1C8xR4x7u0ONjF329yvIHx7PsY+
JWDWI5psUOoccIWYrmZ66vwI77DGGNFF84Wq/+bwMh3L16jNaOS6qCCzzKybPdgz
cibvrcB0wZFcn53DUVfFGJ8H9jvn0nSchtC4diqiDginPVTPJkaUSJxwrS6gxXhA
kdNbUzlQ8sods0TML7Xg3fnQgjayut6RSZ1Skki5EnH5iX+TFDWMugnug43BvK6H
LZDgWTXfh8me/mowMnOni0rkKDTU7oCYDsqPJpmpW0IBd31Y2WDEVFvSZoeoaD2I
ImTYhE75/eitG3O9c5ix7lSqVcyG7pQYVq6Wnz6kaHLPw6BTsSAnh27w9BtUiSIl
rV0UzwkqYN+YvQbyx0Uh3eHPNvyhiEAsYMbOoQjeDLwneIczPqtoihXIkbbAZ5A2
29nYpsj28Pt80F4cWN6N3PjvXGBWlOPls9jj+u0xYDWaXqwWPYZFH1I1h/womrsl
eN5ADQa5LlUlpEq+iSHgOQhZIbhZGwj54QFI5m+IjSiEiHz/10c/0YciJ4hB7xJ5
ak5Q3hzOx2qxCNsNp3OioL9WiZ2MT0TLlPFIDAikAO5qGH6KguLvW999AFu/Ara6
T6S1GbV0PqzMESLD8PsoyT5FNqubyNE+Ti7ETQ5NzZv5Dd17hZRXf9Ag5isYCKWR
86xhhv1t3uohp8a5CXIzFHU7ZP74vJOM9vMe5HKuTLUwjU8rLaKB5m8WzM6Pzevy
X449u4+1wef/xbwuSVM0oV+HNs405F7OA53YH6nSzCDEJgAOC4VdZCm5V4TJFGvg
ash47ikSfXPdrEayUyj9tqJ+vON7WKSuBVAVsUTGd/r8JOvBrS9r8MHfmv932LEs
wvYfNSuJYWGPOWMMUdfmqpa5DfsRPQ4Q4cSX9pM7lMmFU2DdZWyC7wMZ0WC87Zi6
XuWmvxgOm5XIk5glo3JLNAuCMI5L12Z9utRU4ppk/4Suhajm0BMJGGzXlHAOMGzm
YoAHndK8KO2tU6GHIi0hnWDTjNBg1vTnjkyoDilvUON7UR/0yHBZQnKF2xRYNeFg
55Hn635uZSORJplR8SDmjixnwOtHTd+IWtGls6/bOVE7Yf+QlveiqMXxbxOoXLgO
ccyucrz0nLdR42gfS8sa0UQ12jazjh8scxQQY4ufFbzwNeGVoJeHPQraSOg7M6YM
cf4DJsNOS/zeGdV7aB3QWA8/O303CUYH1IP2zyoRD8t1D1HFOSUKrKxa95aXRJnf
xHMu///EHsjJguGOVnEoWnBgZhBBtEarLp8MttNcL8zsLrMxwcpjpEpx+50JkrL6
cbV23iCvILpkMJisYLwvLgv2K/x3PcpS1211oCh/zBUHWkrbQipHbfD2+8NeJu2d
AJnDMF06ZUeHpCQufzPtjRMngukqyAY4qB6Vt/D8kAolnGp5Jh12b8iB11B9lZen
SSsd0V8jWSzVxGuTptvO8tB0lhuU4IAT9HXxd3jx0onM1UmqGrj+9WF74xDD+/N7
2/xN4PNVjZhajs7w3Q//y93qUZgH0xgipI7u8x3izXaY1aXnBhtMJd1XhcPh+JkU
B3ekKSEyzhgm0yJAg9eNMPSqi2ooYsHU3xqiLwclo4M+cfiDSJgcve9d5FZQhA7W
RT4mmmVKIabzsJ7ZSLK7++NA/z6hZkmZW2RziUXKGOraBxKES9h4cX1L9vEFV+px
sxl+Ckizu009p4oDMTFWM33TG1XjHQKpDNvDClbB1YnsCydtI7AdWiUc2STIG7th
7y8xzfVNOhAcuf37Y9q5VvZMhFueRB7ypDeL9uvhdMVS4SL9kE2WAD32ehELp/+k
byMiLZvtrSFkGSTxCG0yoknFvTsG3e6ETWPlXpcLkh34XuMUkfWRZ+OKqy9zdA93
S7YNJovuql31KLXXUx+G3jZBvhAaNGKV/7BKnHq9apenVu/1cLuWhqYkHJYi6ewJ
w7g/pi2Wa2tnw6WT5PoIlaFWDsY+QndSkNNfjeQArGdF0/sHxjstthuoMHiw2ady
Lh2/RZhbWklQL5bxaE1D07fbO8oHyRtaX/7RFLYrNE5anMRwPnaGZ9EW2Lt+fCkc
rfwBpHxYMc0PlIA9N5jKEnTMkfHq0qnQiJZjhWQi2nTHxr2J+KbNafW00MJICTaJ
kyRHQPrDPlOrdThDGLc705d+ncmXFGJrrcXgQiicOPfw8Ic48ZOzcquIaNmaJGh1
lq+f5J5R2LZCu7chz9Kif+ERZp4CMFp5s2nVv8y5ch1/skOEArijufvFExwghEhf
yZCeiMtbtzs6LatJWIhVubA5J8jN4Fdt3mwALVElmpGncj3YIS/aCSj4RTFjfiAP
dcL6T7Z+kGLJsjvDWyFrku7mJIWGdwzhgBBS62e+BI6AMhPT2I2rm1DwhgIj3pvc
C2KzvZII6Vkc4xjVCQf7AxCu2D5ZFsIM2Vsi2CJI47RuOOxR/jWeZokKQfUymn89
6YwlrOpbM8KbMSVolkRYI8W7/Ek4KJSasUXtPtsfXJIkrBvI2wN3Q52z7Ob7lTk7
3CxPbMr5SQmJmD/WrX8PFY0ejuYTDaKVhSK2HpgkiFHBso8wbZWJ3tatZSLRu2Sz
4yqO1FzKOmLI6W5ZZX4WRWNhd/AYW5ezwHqn5SQUxdqgbYIEFV9engixn156O+9V
TN6Le6D+rCYaV+SpfrWYxjTTAqgx9S4z9S2zbZDtHfU0E+s5S+bTyatgMvY6knM0
ns8V9nR2l2smJQfaZRZT73ZVj8cKhM04jnle60g4fbuYkNKr44dHIDvfDoX1MjvU
Lhn6RWW7LLIvm2e3S2bZI2LTfTtz0TqpDqhUcBhfuzRSb+Lf133NU7R2lopiWi6f
7lzMc3Clyvvud8ud5H+fa33Q764Lvg+o0ri9mK3UaJ0dOdHjqxFCHkO3sah4EL6P
eLV5WaI5CML4RfP5kKiKZ9pGPldOTcDgH0yJ977+24Bf9zA1tOLLModbsLouIgzS
dSMlxScoJvGuKRtCGqo0uF3PhmFO/OgvwIESwxagF2KbalMZ+4XE19CbpAdtNFvw
ddO2W9hx9hiiiNA5GDZKV6kvBU+2DeFcRAX9AQXmxieIA8ijLN5MREQRW4AhrI2b
dRX8Ns3t7TxvBnq1MUwJ0sHH0T/5+wTNdcreBeCaTEbf2tuB5TV6aR+nIm3+W/y7
jJMohseTnMf0g3bLrreTPra6JcxpE/DIE8gJ+bEkza8ti3C/e7ZUEMnQIBTbwFA2
Er4S34fnKfF9zbwLm6Hd9jm7syiKrYUSTLoTHi1RMv25khb+GomF5UuZhDSzC0ws
cYZkbhv9ehsaRtI7sNzspnoGImbPD4PK0FGOrL9HmED9Iz6vvbv2qhCWsWR7vw/g
VtL1OWch2NKuD1i0e6U77D9GKDS3Vt3BtC4RGi7aU6RvTtPQSV44KRV7Z1bpzku0
8dw/v5K1gm62+CxsSUTiH/9OYS0Ntpf6m2tT/0qAp4fnD7WjVxKpdMTexytL4ckl
Eqa2ajmbYtJAUtUcCDvuSSWUsXU07vUxjZ1X8gO6H3HS7EkoMOiQ+1LvXQVbLBmr
ZI20bBAxI3zx5PaTwpULFus3roq7eFmCxQllW3coyUp9YYL+PnWf1cWxZaOXGSWo
76tJ8XEu1CVgTWy2l5ekDrUQWKuFPkDlelQGNL2hh3ZfJXz8LgHPcHs71pjvFeh/
AIQhwfeyZbTwDvWvxVI6m0kUozX7JM8Y6nz3I7pyMnXiQTaVmOxfRVUFzESdtqza
QXp9MuLoOpk+wA5tLJqp7XVkhG9wlpUrX9IS3n7sRb1+1YQgAXfJP3j6ycr2DhRg
/DqlnJwaFnocU/f5bjkcwW6LpY9ieuqjlOv0pnJOCda7vbK3CutP4yvGHwCqmlwa
g6vJIIoKlqSyrssl9hlUn+PArACN66UrtvO5lnWCy3cAS+xucBp3cbWUlVZJubkZ
emCAKkYkKuHPPlEL5bJV8bjP6R5aQLR0nMUee0W/ANmxvEhbpK9pSdPcB+1oVvCY
woRxMSIkcEmyaQV2dAav66wX5fk2o/rpgY34BbSDZ4CVxc+tIKs9aDqLsJkK+N4Z
3GODkn0paM8LWfQ7wz5FFu7aKpsr3jGuyLdPgtzLtY6hZsfW/MiuzOsmvVzdo+V9
lSHdH3fvuIRnqZVSpKEdsxoe7JpuSNEwwNC+Sh+E1OKl5p01FUSpN67t/KsTExDa
Ts/+BjrFvC7yjvvJNX+55IKcnJ282I+g9cl1Yq9D1Ghch0kQ67OdHMzbcwtxZ0mb
ZjGN79Glo5q8mt0+GgcoEY/GsRYFyhW2qu/RIije0UkD2W93LEJnyBf7nhQ7npxC
tQJ2r9T47dddp3PM0EGWDS+1c4VdQtb1euhQL5QQYYr3dy+5EwZz8Ej6MlR7Ht2R
mOaTrTLGuACxW18J4WFHjOpW5c1YvEue10xdoaEwwMbEO3baFC3HxJ0JmBsUd49r
5wAR66Q7LdRpfk9Yq3tii5jInu4TxHbU80NAOY65sF2po/kpeSFUk9uy91bHCdEB
ykbO8eDCqx3huYXAeUm5qx/Wr7eTl1FqojO58GNjsEGCDHY5Urv2/nZQDAI+E5TY
3orNj1CFX6dq6BY4hAUUqf0j4av0F8Y3gcHodCbUohXUprXnOKx5GOByDWNYX1MT
VR91Inqsc921Kj0vEhqB9BjRxHDthI5QnwzE5i8A4F3vZJJXPU6yKupKhPV+g2Bw
2BUNb/OQCngRGx8Fmf3iwCPcU+A+4qQP+W42V1rc2oqNDTPjW7ZtEyCpgXeLrmIM
yzmBKgLLUA1plx1QHxFi0VCRdO/Fc8ItMsVbYdydN0iW4iisIMFTpMX05ogszAPF
/dI4pqw/COjV1zShuw0xQ5PvIQa38I+dG+Ax6oHFjTi9Tw1BpZhxj9UXJbZmWaRF
+SV7tog40YIG/P3YEHzN4ZtKdMoowLrXy6FlCseA41ODRD4pGkBT1PmSZvXZYvdE
el5fvsFcCqOsQaedCZeI20xaBnYRwl4ZTPNxw9R4oF/mKvz6AEAqptf4M+S8hte6
MIHdBQVw6MkTJxBsEyMItxzaaVd2QcTHr/8nf90vCnZmK1Uqyv/3SdFB2V1IcUk8
vTJMgToc/s/NaYAqvLsuYPlrVoseHmahIV2NikBO2chbmZvzaB8OcNd1J8U7sR9u
nZsoflnLEa2gAkw5hDGEWC96B3wa77mAf6hrjfkOXTPmirqVIqjw0aJDCv9Mt+rA
9hzk1QwA19RWXRN8jJkTPftss7w86534xGELZmkB1qYpa4I2gzbJRTQQIU4EHZh5
l/ASFwZ75H7wrnGD7U/n7s2EAnFpcbxgQl/hrA6Brr1/iEglThjF4KDgCOCycuSc
Yk9hUh4kvnh7wATXpZ7ZynCItlJ2b6255QMx7LqhFM8HnZG3uzTk1rhXeLlzMZAV
rHevQ8QM8DmGErLfFQGKW/ghDszinzaa7w87Q7nR2GPypH6C/Y0SDD0k1XvEFJfs
ODjwGOaLjebTqAuKZW/KNfiWZVhzmPlYIirF6GqXaSRP6i4Z39O82pW3XLps1Kti
yfUu7icGQltJDjTLlZy0mNjwAAtOdtrbaLX3CUiw7lApgtUGFNJTQgBRijJ0o863
0YqMch+bX4SFECm5a/+AtJlZ+aeZBUcEIcFH3KY6iY8abZquAsvfodF/qLLBny20
IN2+kaoB0vSd2TXBGPksia0rOtmZBsLlGaVUHEyBEtUcqs9xfvJRLulqn7EwBWlf
GOELGGznVdF3Hs9P0aNMuVaKIsdvUeSTEuEvoOJRw+5OHw2oZIYI5FXTiOp04IrV
efWoI6e4dIAipdKGeIpQ6vxj0BtyCJuCD7kA7l6xHb1aoPi8G1An3rzE/veM+zhO
J42oH/Mm3TBKPWotXH7S/cL7xnQsvCO1RLXcnCzGEbzthcOmMvzdNnMPQUBAgV6H
aJeLDh0FzIfCKmzchU72YV+d3D6r3YQVdemRHuFm41nPaMl8mpU8azlytRG1QOBl
i27W1xIv0XOPfRATEvOG4Z/8eIIyNBUf7S60PUttWKOxPqCCTuo6bZsZSZd4ZHBH
NBxhS+XkxBtGWjqa/O28gSEPDS7M6uD5w1tVgPJRW2xFmj1iOtizZdfniJiIL+ZV
fP32NH4Ov2iyjiGE3W9iW5/LdbfzHa102FYPXViEu41GrD6QDzApXzirMvRWQaMG
wJF/C/e+9VE2E4VLDzyQs8UGdZ83ENCJwVrXvdILwGWhkprNy3/2CuvUMB/tazNV
wPAy10o3uWVbsEO6/9e8Hc4oqF+Px/n7qomNOWRAy95MT8P+Bu03p1isp1l9BT36
/3ats+2yQfFpckPI3BA3G9KLyuezicnsDtz5FyAGXP4hEVwcVIyYE31Z2+giU1I3
R3gYcZykH5kv4jLmcxh5qp4ex6PfDpwwXw0Wo7E6YCV5NJqNHzPCUHLQGt6V2gKA
TJpU/SFbaR0Irn6Bj737+ACmCnVg1daZjwkJgWzYaI2tShw9ofTwo3nqwTNPiQXs
ohTjb5IFdmzPwXfldUdBwFq+dlIwPZR7jstgQUZPvf3/dXoE2mrS9nd3DBAII+MI
0njewwDuN084XZ32LEEQtZLcqOaXYCXsHh5QrrNKnFVEmsNHGR5TYk3WQCnqG0Ow
eK/hlIo7kkh6vaeU1ir0KhCJ8JAjxqedFS9v5Gpfvz1c3ksBtVS8frT+4SrNT30s
5auNmN0MEY0KkYEJoGsdUwM1Kg0MhOgMfpRfYjnbYoHNlazYZYmMLTmRPPu8jZ1P
7wvkA5lS1i+ItJySufICBB2FFv8rnVSJB7QG6giGNLiMMqBCnlOH02iOj4DGxSXV
fbI1cJMx3zl+tiRkGuhVmpvF4UByVKxGXrMI+3Ms+naPl+QQTOxnFl25jeEWjZkW
QOz+vC5f9YlRMSKaeOh9pLzF2WjMTiZVcmA5eJv7ujAjhOxVoDghBQOHC5hU4Z5u
DNl4N8DCqqwja+XcjtneBetIUIwB1UVn/3IX4antWXjdjD4QQL2PV+LHCx5UHBiu
g6d+/eub+x3XKKuNA5EelFpzGzNx6b6S4/8PP4zVZ4D2EMEMtvbTCF0WPAQpfvAA
4h2ResaWsCfJEgPPbEnh8WOYL8a9qr2OINJ9JkH7YXXkVl14p1UnjW2NIuyurgw7
A9b9rGVnBDKwXnd1tr1V2v8SKLpfVbW0MvlSlZYl1DxAv7Rg8Z2KYHxaF+nF/J1U
2b50z7LvPlOll5zja2f4vQ6HDeNLzkhEQe7hD8r9pZyGXlUn0N6gUGEaPctFw2mr
lnESYskvw9992g19cU2gIVQtItEdzrM1nZ/ox30+eg6/ggZRHQ13MIhm7HuKePFB
qkf1ujtq7RAZvdmRWFheE6S5SGcCk9VqtptDE6D05nggCaIGHfoM4huCwviWAkPB
eKdeKA8GF3rI4Q1YNu1XSsWe08nPl/j9GCrcbJBk9CQ6ConJF7A8EA+sTt3DbSyg
eAWVRbIh2JB7Zr70MuTuh9TpF7lAVnipZ5y8dORZyJBGga5toaN1/L+KQKV7PJez
WCQaaXySVGaP0mew4gGT0Q/wqeiC6+zscXC5HicN+pV/Rc9ez3dZnIYdTfXXFYi0
dykTvv1DbH24cX613uTZiJdAv7YqQd+ZFN1L99oiZ8xBDEQeIOUvtom99vX6wt8m
+Kj6he+O1Rw0UyfxrUeXRPvfgPVRV0OTfUUW3gMDo7vHk8KKH7ZfbVOXfnSm4PGi
DllBh1apr+AndY1IDKMBcH3wi+NRfoU2rF3IbTjA2fFM2Hdg8Skcz0jnHFSzi9ln
VhmsyO/OftdZxrqZ7qgjkc8QyMSVal5tnnZvcl6ZwHiuSlmt8oH63Xu/BhTfcuGE
OnH7xEuGuJRt0DXGh+0fMQ8x6QyxZZlntg4nEXg2XCC1c3Q7MbqidARiX8Vq/FJg
WqHlStyBo5vltdu/VPNDYByNtqsjFYiTGkC5xX7ruDSo3QVy6LknyZHyja5lN6Cv
29/3idtLXEw5bElCU3FR4wPxukVAwEfiEsU7/XtCXX40idA2healSnHS2EvnrCFe
5DA1HKTp1DGhe5F7EgACIFhQz25IHKZMVCWNCtDQrF6F4UQJ7Q158ARhyBZe+FmS
CyTMer9Zs2j39gjmPxdebctN5gnsmDNBPDKNwta6fnb7h8jQOvbQt/B0K91MSgmC
ojwX6cjsxpvf5xjDBirFgA5lpeoHwlYCwZ3Yc0YU3KYqww99hzP9ey06T2zcmAs7
UvAbZxOYNgz5+JDa1c+k5FxZnXAewcjlfrLaloVNs/Hf+IVscnX87wUnK8wI+6xH
AT8CBcsNTOHKNtPfpt0YzrNwyOUrYLhUfFItCy78Bxwdo9aSu7dijtr6XQAm45as
QWsN/7yLt7E07yGU3vCVLHoyubOokWEwLvyoGF2MZFYkOlsvcvvljyvo098oliKN
te9tQpIHa46R6yuntQToOD3/z3p9AX92wALy7uFg2epIxohvygsUUNgcj93T6Sa4
PrCqGq89wK2PXOXWRgjbiqZyf+l+0klM8nPYxwr7Ljc9OMkcfnvYtCldg3brxOfB
Y+GY+O3y5ijnKtFdvmg4Lzn9ZqmuADklZYbnVPeVWNHhEzJh+K8Ti9vmaVRwMk/T
pCy7XlGdBAVT0c5VVIR5X7SeOs4VOzkTiLvCid4aLEKE9S7DORaMkopLjs3Ccu8F
+bonQOZFoLoXYBTgXGChkKARY2FneemPCzWzCmR2ZD85YmKTt2OrwAMMIaFreDPu
BYUVlPWjxU6n1ZOJLDTg6IKhWUWQ6kPlMHEecd2htf5eaUV20yJlSCeepPs+to15
0nDyWwS535OkknQXWkBaYH4ccjWD70+5yFzpeLSOuCpVIcBdHwKi+JTEvxkYOXjX
tlABai8YvajOHewSOeB5mI4XvyIW1tF+UC28vgXwFioMJI8x1JWAvBqEePXZqs5m
SEry2hkrmS1waqgAbXIGz5JWZ/Y7jH5vNMVg36qcmTtAFq008+lzsdYuK4lqz360
wYktnD5oBkBoUPdyMXckUyUurQcaULmzGHTqkbJ3Zx3iNFjEGHzCO2WuOxmjkADg
9ulIiRoZrlzFfw/m4fLicNCgTOodEmmIT5tJkPDHCxVJOUfVmhHhKIn9UNYPZFd5
AlzymrWAbMi2G22T0/SNaneqjTRlfas1zg3tVvSWxu32lSyzs3Ei00ZWOy3cET+z
1urdpi/vW82DyBBqkhqjuN4v9Si0jovOK79TAGARpkJmKVT5t9GZqQ1HyEecM+CX
8rDc6bCGsnN0b6ho4Al3ifPwIvn2q3zKprT7hD5GzoYc2Whfa16N/7W2X3tywHkA
+4APEG8xW7hp7TWR3aFSqyTPAcezCGVApP2yMiegGBGKtOT3MplVH2ce/O+ZsnHU
UV6CnteQjZl5QkKm+8ciAXUbujcH/W7P4g4WPG9+XwYf6xJjLOW55QR+OawBhoeJ
aOqnfvTvE6WdVwNVXovlmtju4RUlFbUdXasHdJx+MI/Q1vUE1xHw+pJV8Ie8NSR8
H+bs/zEaIQlpvtgiqlB/dxyMPB85sZArWk7UrsmyI0oHSk2brhsdpvNq9AzYnuzq
Eyc362Qr06zykXcFMTpygluAsbp1ymz6NULPT35ZY3DBcN5IR9a9jrNqq2HVgx0B
ktEU9X7x5ocjv1/61OIdqPBNH4TpD3rU8xX5PWF5Hgka6PFUKsXKAU4sj6m9Mv9q
1R5GzzXgPyUKkouVWLJZMTAdDg8BkFx5eHWYaXfyEKbyOiBB1uSzs4Daf8d3szkH
eEO7NtgxUrhAifY4DOIJAYUGNzvHGH1fgp06q2r5imaboLJi9UsawMCxK0rEgD5I
xzSopBmcmv2wO/4ttUjiRqR6KcNPLrR2wcbTFgScK52Rn1smT2EBO0takw8FyvnU
A1ad2aQZTc97julnYWZ8FodDgHE6G10oPnJvtBd2QfYtLpQL7gFEvSJinpt8Z8tA
K4/v38qTgcf/BUIfE6ogN0EhBsn85Y3gis8DpYlhG0HaVj5wJ2DY3DqYLJYsznUo
cMu7fqLDUrfOYlYB0TV74kPfLi2X7Q9s3O9SLrNbJ+q6ZucO1TkZr4b3zPS8tTmO
M6kMaXzPNoz/ekrN6OSVumReBh7wrcWwjbWdeEBOHqRIYOFR+MJMaKhwMzqoawWe
wqFpuZCxgK+bd7fzIn8aH0RvpJPZB1pn55Ob69JWk9UNjAXQwge+m4K6vxvCiqLg
Q9rChYebMDvuBdBQuOj2vcbjzPyF8Y88lDuHUu53RoOAAhSOE8SUIuY0MMoIa2mw
DKukVyW+dWKa+myQrRbwTOnIazq9PjXCSGLA2PReZCbRJwgEOXp+lBh3ny1yEo9U
phKHpCS9dg7CK99naXfRsaragAV9eslZ/IScHiWu8pbeI22mP6kwBD7HFBpB8IF5
5Y+Tea/n0421nQefgAAUmmtBFFVPg9X+NuDcAlPspbq8Y1A3+e6EOVkAtT5rZEkM
1/1NUDcYqQrpzNVioLMAc++ftwx4sgliNPY08uKVGaiE0EO+FB4Mnb16KxVgDyBw
lybeAVYB119CqgDipJuBFVm3a4B/kwlQq0t9rAi3iddOAsLfBaI/2s7oz46o2Err
jKBQicAD9mFLCftEvjcLecmUyk8rOgsJ3O2Ay1DXAabfNNA9rMphN76kNYpboKPQ
lEORieKvQvEa+yHQYmvoFaJPQV7BJRUbHJBCswXIz2jw5JguU/bqU/NfdjRKCTDu
7XsFC0QsaLTRjnzJENMp6i79CUHXA7G7wrfaFjYBCVDzfCQo9HgcCUKqkxR98HZz
XT2ZCTTZp1x9dTq+0fjfXyfRob4jpjZqV6I8JN9UAy5AHqx51R3NMVZayZh5I0mi
Q0sp2b71ZWGvd9Q9627PYJoTU4/wwCcE4fgwxgvbUb2vL7/ZrwHbVBTbN+vBmX2G
uCs1RTIs+gYK118UFKAOKcjS/+9uS9fzr7QCJ/74sUDd/mZJXrfcsRZnyz2epGwb
SdVSGSnbqTWa8CSUukcN42+u8u38K5wQYOD6UhZvXg7jKLnJM4z3GL45eUryI7Kv
fUwtWFTRhp40fMDCSDXywLY+ZQLBEufOAYjCMPUha04aPJB0QGFfEV6qD75KgAQy
ajKeAt86r1g72FSQLpXFkNp8fwU0t0E/sUpf8/FDckr0m/N1JEFZQqxEQCuGCIZd
klB4wXTbWSWnZs+dT5LBMUeXTCJJfTpi3MTMOvMaUl8Vomt1GVoyU6fOK6OTCOtw
wmJP8kb11RxVq1IRSM3WCrV+kbHe/sWB1Su+4xIjYid/LcMjrkvlTmaoYvQqAbKS
`protect END_PROTECTED
