`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Ce7stuAj5LBmyo5iKiVa3n4pKANsO4tsC+7BrZgJ0uHngRbUZmBN3G72WVm+l+J
LTlCprTmBPfxKt6DOj0cOzHPYufAFqgnGwItmSB+3mIeRHfwBvQS3TwKN8OBoWTf
dc2yybqi7s4Tz+LnJqBuKGbhDueE11NOpfj4FSJPniUZkBqGAH/PEwC07fJkidQh
/xzkBFQ1rRW/fhJIkt5ZIw==
`protect END_PROTECTED
