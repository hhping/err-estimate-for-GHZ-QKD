`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
afYr1L0w9HjQZ2H4R6vOiJxsXSx99ne+B5CC+ic+KbqllBTd/bpi+f8zbVEEKldE
Vh2EZXLySFrpCbOqJ9KOJsd1+5mIQJQAS/kR1Dx2RCeawUhqx9OmkWxW4aW+K+Ql
plSXCTwKEvdAQlhXoOuB5dVc4cAh6SHt1jzETcWSAgHEnM0gZIevxN1bwm8SRZ3P
VmkjXW3Vm3UebiMkHD/3E0D8w3mMcbxaM0aaiH0kqSOVwdyHv8dYa7gg4FYME47Z
6+S4+af/i40dzL2Xg5wYohpV7Ys/O3bWVSSojo37cBMXfjJkh/8TonTS/xe0WF74
Q65Bhz0ZkNS/hP67Wtys8fXIuC5WbvqYVswfNhNU3/QNDhyjabrAYZ5XXuMXIaOd
2RUkjDqZY8ryVc3UvdCDw8ur4/eud2UkpESKw6ducyfuLosVvg+7hn7DNVHJZaOZ
BuMVkJPnD+14pkg4xzCNiYuvd4jO4CA5tDm0JGNdkwopcr7lneErYBr5INFfxWSj
bCb8Vo3UptzVqvC8bzWvcjDG+W5o1ZPbJ8fRYo32ubG4mWCVp6GYkmPxLff6ntsD
`protect END_PROTECTED
