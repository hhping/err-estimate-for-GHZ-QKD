`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/2pFPrP1GsVHXCuPTAcfZ/lxSyHRUO3rQb/8MYOL5GL8RWSWrV5q1r5YBS846Ol8
cohQs9l+rp4m3bXldKTnZAkXUYfcb9upLoQc173LGb8RJmqELOzhTQjQTaVVJ60c
HhcscAP3YxYilHLRsFj2T1cok8fu/lhQw4/kZD5rRNRFfJFd6HEFrXEHcmWdeT+T
2xOi/l7xLvLYtiGoyPAeSt3AXOMSe61pqgEXcuLEJ+LcA1g7ppUf2DErsPSfI8gD
pSVJfs9v4Zs5X3l5g21zUGpwun4D3z9Mmv7ygqMqVMLqXGT92tJcks9kH5PXvXmB
QN73h3F289qviFVFRqK1+JBiNGsvlGbHr7PYNVtaTTnbNd6yW2Gp5o9alz15eLTL
JJIG0sk93QpNXFWgDRYpQ1an/ZAR3VibzhdAWl+OlL+yKPpSYavvWJE30TcDfitS
gaL2cZOm23G9+Qxk+BGpdexCWARWMj7adlxdtGAYQG81JutmIIfi+oqRGkuVE++h
LuANQ1bJ5yRizKY//0DlGmsAD1uCcmG8Sw81oP2yOi00ZKad1OhJ2jayJRzML9I1
JM51U0Xjpo4nW8uwE4REJ1slU1azyq15d6TZTnxD2hUsk5SVfBgfQkgB66gjxGeG
uddejUgM5wu2bhSKwskbzwzJuUjTmqcPdIQ0vEORLRg8k4r7zU9C/XI/l4imzj3l
Rtop7gb8sBa0aIJQP0E4qmcrMe1YpqdYNiMTbac4RhI7gjt6dUnBZJTwPhx/2y5c
kQsdeIDd03wyWM4ZTWrzAtUBJNWRGNMcLbJuvWiezc4Jb1SCHi6RTmM+n0wekog9
kA904R+lHmRd9B3i8ZFQBjT7/Xwyfb3mBewhNYYKJ8fsWL+6uzFFy/5kqtMjPJLb
AGvBTZ6f4qP5s+wQVA/sDlMZ4XfXAbF1lAeGcgmSqE4wu4ddKwZ/WJqDbCkPmk3w
eemXicKA/jCpDJ/O71HwZ09nXZohCWbJRi7zYB6nkRK0kePZ+02iW0xE9nnDdPRR
hQVsBmTUGEQmV6Bwb+lEmuwQWEC9Lnp2tdgCw2cmdYT7rG6HFasKOgC8C+wpcl33
XqAhsYr0B5/ag5EWrnAukcZhI/LROc7WrI1szUSGJp5UNRS/2bvYCI/VL8nJ/dmp
E4W5p4Ozmz/GBCApba6ISd2S14PZdnZg8a0ZN5PJpuz9B3lNupMSe+S+VzqBludu
ZSqUoxY9saUUcIkpwhCVJNe604ZodVFSMWLa2IMYQ6P9AzzFXRLr2PMbMKEJ83mP
wLrw1/MB2GZq0DexZsOc2C6UbVbIcBVUB8aRjwutW3xRFOMN7nIO1w/9mJY+C6ZS
VWsPF4uIOy7bM468TxOnapGU2KnKNjTE+LqK/XLulijq16UpTM5MzMHtDP1OxB0Y
TtMB96pH9rlbGJrH40905JJwmHIjx/Xw+6cwxwq5NyBvFLUgpNND4AImt2+AVhxK
y3BASdnCtuHaUwUIP1qsK0ovUe/FRY0FVOIEXsoelaTQ6Ho4muauihc+Cq9QqFm7
sr7EZswi6d0Y+XDRyLcH/D7lAejIhwtUs7Nf7oQbrvB6nKx3k8MXZJoTgrdOHzJ6
4gpqlqDRLnfr6FmPrP7IW4/RcuSa+6DGl9MZ1lLy/TZGII+Xa8AzvBiz7Gk+OO1m
BQ6w4MpQFHTtbOn+5xKbjguooDW3JMHR1J9ywLjWlT2Kt2NXohz+tQcSnuBVTNeI
TTlit7XESRYfFVyEciEyBC3nB7PBPWZe1erY0Ff1MHvl95oZYPK0qkHTiIqF7i95
8rkUr8vEnYDUQBd3Zp0+W9B9MyLgvWLY9GKoplaAS2jrBTLI0GajYkSgL1QESSo/
ZD8f4Me8myjn79k/dXqepA/JKMkW2Tgl+byo5GW78VihuSM+4A+VGg9gnbDCuOoC
YW55iwTKD8bLAp3iSbNwRtM83EW5PMTfXpNRJffZck6/2QJwwYjZH344lKxx2lj1
msaBNcC2/PlkOrrn4xr24wdV9XnoO2A4DMj2sRgwRBCUjhPvyNAE1KAskgoflHW3
fzFQRdy5ff+juo/q7zFM8gJzY73+GD25rHs1bvO2wpIEhL24Jt57ezcgbt12q5I6
NR4XCRBKSO0oHl/VDcV7qg4W5Fc02SUVJLIfyEiDtcSZ5tFt6AUhFqye6dcLxUfT
k1ZuFkzftK7iRYdkGZEPmVXRS4pkJI7zYGPyes0KtJspKSYU0XIyvdPFhohGuCw+
9+K0R9NjE7N4Av01b9fqzcDG9lWkMIHf9jYLEG9dmhcFbMBh3IaXoJhqkw2CnBgO
qhpMTEdyxBLmEULh8Eum2kpVWpvZrWskUolo5rQOmX1r6qIA9fKzu6a7FrbDSnnu
uBCYKfj3Kjh3Xcx1ynMDviKOVzwTOyQcWQSKGl20ghtsqY2QsHggLphJDr/MeaI1
8wlq0PWF77jjN2l0SyVBk2uAyeDmmJYAhADToYHQ9vkaFFpM4FUhPl5kCYcfvR4v
JVPUdKqqHjnRe/Mx0akydkCcSKv6OtbcYrEWp83QTIlNcqS/slPfj6YB2A+zmhmp
cwKEw0c6NmQFHKtO5JgyZ9Wr39IcjeFQZTtpZQ7iv69c2v4QUgJguJj4YaJslTxx
Bvy6kSLBHNSwiqcziuuR6rSLAJLfbr41h2MQpmyi4EMFalgvYwd7h0qJAoVXMdjU
5CaYiSAfJxK2b0VetFIrdxg3BalSRtyVi/9Bzgh4rsj3txIoMicGLrtFdHdLCKcS
hweX3Jzu5wtJNQH1Fd+RPMht8MJP8t1I5SOJjEc6eUGlxDDiW6rrekmBBidN/hGH
Ox+6vU3Q0O0zFYg8w4DlmyPphL32P4+hs4pbCDetUCAt/pF6Mqw4qRWoPbvPMkpB
mZhhMmcxeqNrctGZXDpKMfaMAZtEbhkx1zcSemMeCZbWHTfME4PsVAh7TfP5qlvJ
qdIeCmfc/HMYHxBSd1Gjd4G4FtUlDxC5q8s/8Nz/Z+Vqtw/j2X3Q0+BzeiKlM83y
1fRevcvkVjXvXx43n6tDjiLfFsnYbHg3FowroOKH/sU62FdUOTc4Rulz7hvhMYxZ
perv/ETfsbgtq65EgXWaYDjIj2R5BY9Ff+5wKrJK5a6sE+7ECcncBmlKYuHuUryt
DJ5xOm7QD3aKiadCMyIGeVhm45V5vjASYXMYfS8L7z5+QtYvv43FKCaybgtp0YpG
zOnZTdjKPWaGWVmp8AItHP4RqAKzIcw/R/njKHIHoAEBnKGm9VDCITlCodP8jhYm
l+SR/z8ZJYG7jIZOkmF1L7m1mu7zBNUhtWmzO1biUH8od+O0mc0qrefWQ3Bq0AZE
iOt5QWo4Rqs37PLyISyjPQzOq7UFldtCT5IXG8yF438qVMEZvrbvAH3/c4+lCUVh
1kdFqrtsGSUXAwVJuBY3aAKO1oV9Nfj65HUF2X3uKwJhWXJmcVFpuwlnBtGk3sDs
JxgV34NmGahmCGaR2OfWT5xog27udehQB019UcyJHxgkwKRfg/03RPrKrlywNPuX
qawA4vKkTN32mfmdYP5depxxG2yTJbZazFWjpG/+ZmiNwjAv8BR4UpW/Ujtc3XhM
6i+OTwcdAe5g/UEYTl+IFH5sm7ZLJFHyiKP9tFTRer5VZI03GCHpZA2fiJLNj8OE
Vm8GyYWIoQy5k0Hi/PAih50PVJ62l19WOC3CLRDYApYt2Wawl+2+Pp5OArG3UvzZ
zx7KMuxbNpzQouxJahDoAGu7IB43ueV4zQxRztF6Jwmg/gGHzu/nEyl65d+tXnND
aN97VfyAv+FysWjAoMg1Ordqde4QMH/p6umMHyAX6namz6jE40xyF1JWxUT4wk6B
OCRFtmgqUPXDUPuFiX5PcRIvDzCtu22TwMnF8zxbXHumWp0Yr9/VRH708J8q3I/w
LDSSzywxwl34VioCjQBJJD3H0YLHsE6eFHJyACqo18JWKCZ0IeU5UzuDpe1bB/Nb
4noSDiRjakmqS0q+r08EhH7fF48cOm3+IiN4DPBS6zDJ2+3f8fuTemVOhbazoj7i
ZnKtXA0VfWjyqeeboujUFBFn3StfyAiNXhusGUWR1ps+1MTf5rxPJsY9DExkG1uy
rkX147tddkmGzCnb864sow9XmJpyzvQhQEyme8bNDc3GmvoW0eccusJbPMxtw+Vt
DJFVytuj6cEQnaqwymtpOztFGMLqykKFTpEiPe63PN/LSgCik4P5YYHs6wIrZCui
KtQekMUnhkHnuEyk7K3pzxrkQQ0qrYzFyh1yX71kVQSHhY+o6DnTF7r9bOjxyAnX
Jy/43LiYQNCJC3mP5qWyWuLxfhBfCyWe8hx0nYajQwMagxCNYnZJpP35QOX2T3Mm
rk/gMb5tsPipaiPWycjSqUMfQVYzzAQ2tUMcnVP+9ZXav/0kzGW5dHtuJJ51CYky
EzSvbWB9kwle8vcm5HTsDdcjahunCDp9NjLHCHYGFvXNVP0/liTL6ikPM2BS+euk
Dg5RN4CDvipPmnxuNpr6iwjMcsREcqq+HcEoJmCj6HgbBeF/i7stTXAq59svDc+z
pgwNKm7HaPC3fqm4wR9eOmplPdJqTCwyMU/g9uNn2TMYL256EXD114nrgGJxmzN/
oZIj4vGNOCb+6Jsy6mzPoNIGBp3W5es8Iee2bJ8q21V5vjrLtlFgw5MnygNSsZ9Y
A9sBI7HhwYICFEm2HROwJmHxsi6dyXsKfg2Q45BjWJYu8d1FXGzEaQQAuLVDH+nh
uKHRXgWJHCOJ1NQSzNC3poiTqYBFZucFavN3kHAWnPDXHmheg4aE2WVrva2cv55G
+SnxJxhb2YPHPmenxMBXxo4IQUu6en6DHmiAXypwKXaX9AEaGNxSdQxW4dylFMSg
6Eff3hJxKdD4n1J5I2QVnyJEHQSOM3IPK31oaO+qkP+/vITOArLA+5N7QkAkhHX+
WJpWUdp9UldZYhByMVRkB12JiIrsqgcljeXwlTsHsXZ52PPbddqzu9O/nmRzBMr3
kAHIh3VHYumzPrDdR6ywitsygT1C7fnhbdmFAybs8RLmDFI/y9EQ45J1pns2X/p5
JiBdT1tzW2LO+J0pNpJKn3+7e3ky4smSmUPx3+Yoi//zRDx6nmFIXiC3YqXUEmm1
uzOit0KsSNShJKcOFMoTFAbbNuPutwbqSLxLZhwoL6gVc/Dtz/9M/oQuSmRkagIF
g5a1IvVMIRQ5N5UBtSOip8lL6QXac3+r4EFILcWZRRJD/bTJe1pmUY/1osSYUYTh
zDNC9Q3t1fZjjtxdEQ9+6qMN+tp7oIcnSI1IlovbILNogpUsSSXEfwNJ02mEtBVR
LQlDXrgSyEkPckMCPCVuJyO9FIGmoKw2JdqpMSDnSOmVwpGryVk7qT2PL6ExJRv/
y6+jwsVMw1vAK7rlKk0B2rUmGlbnROO3l1lKHR6+hjxLsoBP6X+Zaa/eRTmFbH2E
PRsPbEWIx8Fdkq6TkHWDdjfiKZd/wzsXdP/GXel5TogZW7umcU9dc7z1yiIr7mgU
VkbU04hclhZHGFr9In2tpMkqIMvCHOFe5cks4b/a8BZ0BZor6tQmCpu2rCcfe/PT
MqLdQwXI5/LjSOxoJBUOkriXIOyWbz7CU8CYrZTHnDItvdklkTEOMu/fWh6+vDD3
4RyWeSh/COhuWjsjTJMvk44uulVp0qx9qYKo5WcRaoptuXrL81PL+QrK+ZivSWjv
YdMoNXEMA9c1MvmpVxeKAZO8TZ9hV3CKvI8eYtQWt3bS95ylpkoNy+X7zgnhOM8N
GBpsuCnp1VkFowr+lvk25N59mF+ymRWr/BTBvey36NoVmj/5bl4ehZhBoYPQRv85
wjjd9iaqGqLNHC4zsHOH78JAktoqqcrJmWRwzzsGnDTV9ynQQIrkEv1HAu2TgITv
vZ2HWrWMdD5lU8ZK9P8dhzu793tSTWJepjSc5WargSNxHCNRU9nUHl1DEkr5cBrX
ru4Dt6C3K+8oKQkz8oXHa7VBAYARTgPnIE6qbzVFQFC0h6r+QgR52hPB+pFCSm2C
SZYi+0dZPZtDYJxuzVAMiTxkbiiJJmXk+WhHwgSMvaP9wNyCwfVd77dYi8o4/ouZ
CFa+OSnrqBmCmXX6kiRxwh7qO52vPwa1xdYrBQjfJbLCwqMR0Yi2DPa8Lh6Lp5zx
ETZ3Knq/KfTrNM/WmgIpHbkyQNmTCUtHe2zx1rtXmRC9PenFd/FprJdwJft9sG5v
3lXP1wuCwHYdNmrSmqbOtTQEll2Tk7mYEXboxxPSq7XDKP/81iNqrzme0Z2lkl5T
41xesH32CXr2rnSar387foa16K4sd5OXKv3FwhIDr+Vr3RkJpfT8dYN9CD5X0stM
okthVDTL8YSHgbziiFHE30PTVl5xB2vMJrVDHEr2/9SMdeqz6/BdZy+4/oNyoeIc
rJ+ZDSLszp3Y9/6dmVc+YIc67/sO3jMNgrNB2FLQM3nN4EW2YiRpt7lH+Hv+fe5j
F2osu9FtgSrbVi+CAPHKNqsm9hVxoM55SA+Vso9Di5cUxZgVY0WvEVF8ON8d1tFo
DXfmG0xvxy5QLFDeEf4wsZ4u/mkfEHBkcCvj4Qt3I1N43sgZINwioQQ0EKm/HM2m
H3QGysRy8DV2Bdki5YJjyzSPaahxaM1Tid8RXtLkfgPMS+9YnNyI+ihIibXWowUB
sS34KnWypyx2TpFY2r+sd3F7cVk+AJFspRR+DIKI/k/3v2WSnUSU+eQA/i9uodaP
+Ltlao7LyzvI/prI5lmPOXWgd446kXKCqPfG/VOCsIIp/4NvM67b8E8qo8gAJ00m
1GnqIBR0t12c/8+dXbqA2f3Rfks8po/0D0WWV1NogkRPRMdCsOzRj9J1Y8QPze7m
Tvztj1KkYJUMqjFGiEIBeX7Bzj0xls7uRhCbPbh8dIrnl7UANtSxZGnOx7ldPUId
M2X1UJntH0CzTZCTbrMsqE8V2H28EnJVl+Xbupsw9+slpZnvBFlD48yF7YEQYOq1
wM39ZeWo8UUODLAK/CKv7bIdF+aBifbf++IwvHL6yJhUplLk7f5pCT4L69+YWeyS
gBTYrT9GL0dsvJ4w0JZCTvRon6+ff8ciFdwzW1VJ/1znRek5uMIxycT7HDHvczYw
Qt1qkWVR5WcKja3LOfOg2IS3bv6Q8pZ9aDDUICwIhPLmqJYilIRVR1Zig51CYzFV
u6E6LxEr4My1EnPv3rWIIK+VzekSNryrm+7gevzh+T0O8D8fN0lo7s0+YColmalR
cKxbu7t0sLBCX07+/qznrqLLRWXEBAsmGioeacOrfgzpFPZRaY96AOtT1ifMijKI
E6Vf1H0RbrDah0Nup2B1BjyTp8/2dVi5vavkyFptNfk2AV8JIhfI2zPCaYNjIk0B
COlixSB86SRV4ODMkygvH1F7xZT7BNgJj8Z4uTwqOd/AAhyTnccEs9zAWB3d30JT
kymrNEw5dnf22Ykzj8D22rD3u9WES+2/sFpHv2sJsmMz9jOzdSIZRiOGpafJSFzi
bZkm6lD8+3VTDdpQuQrcEwicpza0yMXC9nXUZyux1NLvjDVP5O6TqOajGyfSvuel
4xLIQi8M+rbGSmJfCqNj+XzQweZKH1axHIfBMtlyUE2FoMSAY+6csZDGI4w/T0Hn
zVoXv3L2h05URzUh7EnQwrPR7kOY/hQyGESk/DFxU2Ap8wdDugGHRe3zKa6M8D0E
g/rAO/rOQ/QHmQ71RNJkJ41Av00JaJnaZVh8VOTnHmJwzU7tsHmU6ri8fRzdJf+8
8/qNWDp8qQqpsgGB2cu8pGHz9gsslbkqcFWI+MYE6TLda7zbrxTv3VGvH9GNy9ck
Km1d1JUvOgGxL25rtof2rR+GRrmGWQASrY6B07KaiY6VZEtdyxGxl8s0GDOEj014
Goh3NJ5WmJ0sKy92WwCx2FB/Y7Zm3jz6UL32+gBWL9D0cOz6yLQcVlsKM8m5mesB
WC46/3EtM58eMdEe2Q5b10EHmu+ODg8vK3gss8CseIAtP/UTQUaMUMd6p6BRWPwS
wQ7G0VHTqPKe4i6QwNhbFEk/HBZCKcpObJ+JD7ai7Zh3kddp5f86OITFjIe/EANc
EEgah1/GrePBmZlImjhaJOh2/zUlRaGmYTiyLsrvTrnq9VETfHMr4bip26mpRnVi
Z5OT5Nym0EQvyMCHNJ8BI8+sNrsuGcCCsvDbh2eEYrsaL3PaXgRijyNRZ27P14Xq
qDub3husfCABg14RIrhfl1hE3QpG9dcST1qUDloVSOzPDEG+zyTXhMdf45F1Rsh5
LvTJgSRkTpDxc3GhWf5JTfyU126DYIl94rOOmBjeEfIABKK37RF0I5Os9v7GUXPZ
kspPNZNDaU+WMmRiHqNGmpdXA6WJ1JwNa4SznlV/87rkESNRdSOpehND2SrqJOxV
viSquVgvhdyfsRUWD9mX1pTOxIDkuLZuCNqDYzrvSosZaySZgefj6xC0N3nWz0Tt
ahVOgXm4H1gy7v/x8iUOqXu0IQJr6jzN1Y8pRfMx25RZ0lMPS9yI7zC3L2sFcL4X
o4urBRxjB5ofPYig+rayU9Upgsqx8RjrwXQ5tuaJvyfSqWM+y/ESvAGpKUCNkI8+
3HlTgPMen5P/afF0D/Me6iqqEe3UTuaKYXpkaeUdw7EpYuMDfAJiJ/eSDQIhNENH
wW/JvognSeR16QaMXpW+QIcAZnssiJM4M4TY9WGGznhE53c/nVTqNQpec9GI8Fo5
33iNoVWKgQrjhyEP1nSKzuymvXill+zKgkkdRDDaERnY2u1fAPvtlSP+9CJboBSu
zVPkYUuv0WiGPE8vxR1RHMK+1BDLapdE5NAYGdJTuBpBq5Jq+5YlQvUm2HSn7+EV
TQHC7MLzHMQYnTOZwOkpzGuyKEgNaEg66y8TWHAUasCoR7P6PlrvPkkLMpQnkgUU
4w00VlFwf97zvI4roqnZNcf70vKwca/tmL5TFSB1Ofbnys2mWZyjlPh07LK5G8NH
mdXP7PUY5LdCjyE3aZHKckoFygTJBAo+yr9qHGMflNxm1Weea/cluN0oeuOQ1cDp
zuzeH2xVY/EedisPfrbjEegHOZIvxXeatXVItYvBxYpe8o40h2OGSseyGsz+uNGj
Pm4m0nLOHSP/TsGlesK5Y1Vhddd/NLDtDLoXAz+iTiPxkn+duq3WKvK0/BGXUJPs
j7wqZLgKH+K9zKLSceAc8+AedkYt7Jg35co3IO2OSJOiUWVuosePLmBvXB4MHkNK
SnfcmstFeJmXxfKIlNzB/Eh9phPS0G7WJ3xTujARRXJBGUggETEF9P00abmlZKDq
Su+QNxqXvgoJTkAvp3wZqAvmGL32yXdv95EBkcvWzd2nfmGCNrg+blSBEuQw59A9
q6z6+6m8a63y++wqyySRNABxCw4fh8WZID00ENO4JO0Mbl/O87Rh+tt4KnWSDiLO
WkjAjRN4/T/0WKXvSY+Boq+r8GVr8UjeAAyJKnLOLLC8ktLl3COd1LPbqHkZMXZj
RCZQDHP8Y1z96DH5UAR4pNpz0FWltyFM6bREJ8S1CE1qUyYWjfz90cAIFwV2zWPv
H+9J2JLZoM1zPYgrhqzUjP0GlpFf0Je0RAW+9IyL0lojnrJQcVgKwLhsWaHAJFwY
Hd+g0rkaA3306cOTt7147OQF916qIQAYdPSg+3ltJoR8M0eLqDKiPqfVDK+UrB7w
TmCRMdNZl+Glk0FKvHdsCJ90gKcgUBVDjJ8YBsoR+QrRMKKPpOkYwgcWnyUBUcZA
1faof9jSZCzE3X+sW5C5T+uZnjB3vV7nDCtBE+ldpF1RMCBhUOEF1P3FguPBRvmA
2kFnyatGIBEMAfj4zsTxn7/SKJhaAdiMVI9z6p8+WwaqOlcDXHbCebVUksuvmuWY
Qqa8SFYSgvwMnXV5CZI5y5yKcdQ7GUf32hW8FtR0uMXcKfUnVLDP2tmg6acmyZWL
ZpB2ucgcomzbz37YnOw7KwRKGm9w/wtuey6Ep9qaja0F27I8isYm369dR7dGf+X9
8IsdzcPlY4bADrzT7etW1I9HzQ0q7DUyNa2s0iG11p1H8ovPbGG04kiNxhpuW6Y+
s7ikJDtKcI72jxzblAMXGohIapnsUr9pAIA/4RtpYRYYhNHRB5kf+zumIsOIKl2V
H9L7ZpX1DHXWyDm6QnnMG+mtl3IWSLDUmeisp3/MFOKEm4UItxmVY2JcpPHQZlUp
2GefqnosjPJV5fnX3r3FcRJNfb+TfEFMCINND7H/imL99fpP2f/yTJuY7C6e+wC8
LHxWflSOcJzgkGLkPzo68rowAzGINDh+34hKWZeJPiidsJj2sCk1I+PXEDeY73fw
a8iKY73TA4t6R+ZEOc7eemblo67tp0nRpJH74m7FytsuSp6r1FXZi/41YDu13Oeo
e1GocPORQaheTZxe1ayjImxiZVGPL9X0GWuBPqQM2eF4pt0bjXt5jVs9HzTnbSJf
0RT/D1yWIvbssDWAwUH3UFzPGVar57DmoohjaJIHso/5yzSMrAM+pGgRnUnvNQgp
ZDUOyltXDuyZqsxRB/5ydPwVUtO9q44ZuwJmbn8qHiOdyQa6sgHmuBY2rhEFRn27
tT+bBXYegGDk2WKWAYZPPWcBFlLVYYY4MUqvL2PYftVN3rlkrr1j14QPPtFdY3T3
pTBsIgC7koW5uDdo0iLkV/+nAsq9LxzoUzQxtvir/HKC2EOlG7FjfbiFKNPVuRuT
GEPWUCRj+0auxllgxPSwMYRLdiMTyW+f32apl4xxZUZNdl5Y17pLQw3jCEXQ/6w/
Uas4HPQmeHkTHe0jMIXirfIaGK0cqpkUBusM3e2k+X8/AtEl89ci8cyaRnSbKOpM
U7SYWMmNmw5+crLT3E+yA7f9ynmgjCsSKQvh9hvSghOo7FgyOAIgEQEoD6iXE9B9
rishb1poSItTCt6ClZbKbSFySNiMt1mBulOljYuHHhDoSSTbM2OtgZNH+WAxDPbH
C6ZiDeDdaM+fRFVfZo0U8JLccBoOn6lwpZV1n8qWY8gtVoFffX2r5YDYUaCg/qSP
cTL3t6ufIL3ncypkBdfAl2oiTF8QGHfTCjQAhX/UOwTR2c6aAdiTB8nZqfcsNQHN
vPlBSWA7snubrMWN2xNhOPel+g8Y3QfNiPGrIGf//fm67TgFSYDJvxdrx+XuAAWJ
y9AeqBNVzckfMD18VTaq8TCWd4Wr10XsHxQZhqv3hT0vVR21hm/p7ByA+ZsOH+xc
0qQYAh0LbQxB6vPxMlxMVGyiNskGkr3H5nKfvoDq0hAJ08qeN/on3dJ55tUgHfud
laBJjkT2W7Riflidm8bnki1Jb+vEoSOPD3tgDnNrB5kfDOd9XNdWtHqMV6RpDDoP
j+qdGLSkbvlFkR2Wb+X/83XzR/nqjRlb5hYFGXY8ZMVQE825rwz/ag+8OQiJLNjC
ZEOlVW0q+HFWsSgLUEd/k4siJ27eEugZbA/JW4Jm6CG6qq3dyJvA5Y8tUaikoeJq
3YnnUX9EwRKe5voeuN1uBeBoDuys0mQAlXO7ri1XIZHhevwseUdFHWOtRsC9baVB
dD0Ldc7VWA38X9/EfNMfWiO4QbD5RY9rW6IcUVX6GWbDQmLcARAyafwCQUprDDlc
3NoklOty2I/3cnB+WUaNKHGdBiSJQfEFIjdg2byVrKaC/5fg5jA+A4XIJ8jDQ3RA
tXcA8wojgMfN49Vx3UIx0hBKEt1CFn6eHhogOwX0NGDa/iGMVvdKaftI+GITPbf6
2h/6bo4oEAjYWWfAEs/FEaANBzH8OFhC8TNR/ArWcHC47/2nyTf/6WD4Js7oV0O9
l2hfuBmhGhLXOr6IDSiDowscOlL8JjOWv9CIVnx+1K+RTLfGDUy8cCUQmPiUwVr/
KU9jBW0Dd7gHMcE2W+rzDYBqu7C0xuKD3EoDq/IHkWT3+vwIEl01Nlf+/UnWJT3k
4/EpJ6UFZRFfR0Ifp7AJtd8fwgB4KNk10beJAw7u4cK50L6IuKd8P+Pz78h17o2E
WN7m+i63Y6CVbDza91qvhY6iy96bL81ISFtxtvy5F0UoIK99izioRaBiqm+66rek
HLXj53El7G5tpQer6EgJr/1uG6TKOcuoFzeb0x1GVKvxPCrtBFfO9nM++zXHvoB0
pf2ocNAuWT4b5aJk4iFU9QXi47sCulelFnI8V7Nv74pUo3P80GGb9YMsZGO8WI/M
y8PVLxwxByTG/gzup2g1ssvzvwvEuet6Lkz1m5uAijLUZ2ngrSfeuMKL3S/QFuHZ
tUz9Nc/GVGBl/gBjn9j/5q608JS0nkZjjAyipnh2lUcr90yxa5M3MZiu6a7oXXG1
iOJtj9aR8iBmrLMA8GYpX1PlsSoHvHkPO6wx4qSJOqBXG6V5AbDB97HJeO2WomBK
k5bhLlukQepudfZ7eU+o13g/ZBlAyyQlxMJ3zADbwH7K0XrJepE9yLvUJxj+/w/a
rN8wDYebSV842o1RqEBLw0VRTxPtXbwz8Av0S2WSgOKUUudTULh3TgS+r9c9IYmQ
n6AHOEijSZ+x16asT+3URSLimG1DyMLSBbdU0lTHIPBaWtk5MEbo+yLyYCT/oCGl
gMHwBwU4AjJvMXEkPzVr9hB/N6CbEB5AiKTQT5hqP/Qaq+4hc6oL4CLWFMOuW3WY
za3UMP9N9Jd/OIiqP+5xJed32HF3pQsKRjCGK+9uCO8etOWYTNGh7IQ0twuyG6WD
LgJM+cAEZki4D8BGSYgC5nkSBwClI7RBj3qYYAaMAfptPCdLH3YXafr+voujNm2p
YNGr7vITc2zSY3ZkYp+JK/DSDBfxQVDnlmrXj1klVGRqgyKJwnuwIl58U1JpNgom
5l2unxtK7z7XkUGXnjzj84srEairzL+uQos3nXi5RvLzzbfTJ6qUcQpy+IQXq9tY
OusPVCqfOk/0xW2aODZxCa2Z+d3xKkivV5LeuanHuXuIbVciRkka1ZI6GjrjL6No
fSIanAYWx62mt390eflL9gdhyt9NcWjwgRQoIFxc1n+KEFlq0JFd7SkeO23HG0S/
EpeKptYEGM8kvKCi8KOdXi12xqvnpvEFn5hZ/in5jde6rUHnLY9lDIkAlWK3HGM+
bCmUioj8Ov4C6aoTiydOQoxM+MmawMqGSPQTCiDksiwfKf0nzxi6s4iLxTtb7cqI
2FHMKjegzFbBtnkYVRVygAqoepFelG1uf6+jMkmafhZ13dbWCLbWn1w8rt/Q0BlG
EqmiMy85T2H/H6TzUMCtn2aXA/Gfpah5HX+9M5cHUCTE9SSgutscWxw3kx12MnPf
Hr5UvUjAcTwzTdeihbcKEIWr4rwevb0uDRZAw5+YFYuBS+8/r0u5bMNHzBCfRl4Y
14pWL/b/Gu0iA1OCG1X4THHCnYg7+9OIFPqEyybNX3vyecTyBS31UMJ9t5EAYgT/
kIELDhVAHmtYpQYDEjcr5+5cVADa9AkKh0dfbcQGL0dWrrofxDsmagjv3ZzYrg/T
5mnwDo/ENkuhbtvutY5OAb+Q16j76xhmDTGoMuUUOnW7yhCH9/JB7ewjurxDaN66
TCj0FHe3g55ME2ESwxuyA0EeCLq+7614tUBWQ9Tvp6AI9w4NMFHP/ucuj0pCYePz
6uBZgclKsx556sWgbJ58/nW7NyEs+LG70psoaEU6DHLoSStvN+tmSV2Q4tyEmX+E
r95VpYjBc8191WIBsS6d+DolBkZlqo9kTuWFG+cnpbyDzeGP1NbH4Ke6y97AT9Jt
r92HapRUflahHBKgint7N2fJD0YqH/ISRWimUi6TGoAmuV1GYYdliGasvLVlHSF2
LMfxHmLTSDBl1rFGwHvxmZ2nZCtZUcN86p0beYuST8XTpa/r9iL47ZzsfHAjgnGl
9r8MNXozQ63tE+uLGVCmvgxdWiqEkMK9nMkAJPxya81cCUA0E5Lajs9dyzydFIB7
xVVI2fFo+g9JH8kVWBzInuzZyyFu9VXn+GHNrRyIOX++P+5i9ohXxMBodyV/cYI1
3aej/pg+spjWlddYrCNT4tAOBK6cG6uliTVPGxct1fW1vriyv5fjGN7Kuw5Kia64
hoMfoNYuBk8q4BXcKbluix+9K6g0IGdBAHj5lHlUS3y3dVRGxQkc4y0OIM/Ay9JC
sjZGlXOLhWC79qhE7Vk89bZk11KdVmXHwMQFuLJIgQJw4WPW10/+9weQ7a4eFL1G
ytzEEgTjw8RIF2ykD5Tl2cuKgzWFwSIQh63X3TvxunnVFlO9ZtZPQpxbx/fiAH75
3tUnXQY9nYMXBLm4lbvXp7t9HAB+/7FjmQ0/+Fvq31jpcbPVthpc5zkB2Fq4xLaD
93ESjaqcL1f6s3s47XxyhKAEDJN3MSUAgx8mehemi4FDjZDZGdxGzG/8wZb3JfEk
cirzaZ9fLWFQ/+qXX0r/KXBmLENcbP1scIyJVKrybxNJsu3ciGuJT539Xrstbc7z
El7Z4GnRgPn+aBZWPsTYYInpXADcoeB4T7OkFb8K0lNi6rp5hjfZTU9qrIXHWgF0
v6gYfKC/GoCGhqzNGxvHTTgadxvc/xfW9EuEJWcGi3jmhY1j2bzWdFvR5ruYqpXU
58gdhVs4xtXvDOpWbv0aivEywziWNhys2159kujjrVYTMphk7enQU+7L3qx/jLqV
N7AAlD/IJrqJg4qJLA3jgslWoWc/xIz/A8Z+rjrpKzT+3S8MzP6gIVmuxyat02oP
QqqXhOm4QbzEBTM3RiL06MhgCLe8N1RCUSnukLOAdEBEzNnG9i/3EEg+tgPhHscm
QkBO8XJgD63FAovMCrvF+kKd0LlpGs2eDCM7cJO8rJ6jjMCqWq3yW1BnFylLew8c
zqFBL0HrFlrZDUhRkEbD2M0wQpb/HEhmQbf/hm07bMKKi2UPJ9m4lcRVWiIZmXDd
ju7+KHU6ZYDOMN2BtdmQI9LhAflQnKSYDDDc9knupu2VTYXYZEXyePtcn3PLxdgJ
0KWONN2eD/UxaSSBiE0Ux5mEO0J9LR9IMEbbP9X4l9D4EhyMJfL9DnJeEpUp/ZoA
er+V+PLwvpem1rCEsiUHmjmz4jzSPqaZXZdPOI2iA+CnjbpcvJgFeJJFhnP9JA/E
/bdIfLLFTbBzRtCeOStcyb8hpym8bVSbuOL8fwemnlLqWKPXNydsKQ8TNzESfvK1
Rh1iZ07g47Y8tRMe6ZejAOm9Ko3wGyS7Y8GhxhuM8Pyx8tb04nbJ26pU6k4yH+q4
upDNuJOeL2qSf5ElzxpuPCPiQtn5Z9xE00Ab5UIybcIrkBNkchfVHa0HnN+YqXCa
yY3GQwDXVqpFFJtfkKd+4Ey7scPSnPWO8idcRy9C6/hP65+7hsfzzBBEYEX3yR34
GyI+dAvoQFerJXEHWs794SOzMM8h2+ZPPZQ5Uy8IxzuSAM4vt0rKLAWWIsiBGSiP
3CYkEHRH3p60Z69PNJXO8VulScwnP31Ry024OW9qLY1k5S7WWev5Qdsccx7brddV
Wcc6tEq3V0pAyCSUIgyNP6fZXMSlmVNFIaTUYarRsjEZ2zTE0oLW159QT2DEqXUB
l0U5cs9v2yH7s4hFQSANOBOHmtoJ2y6ehtWsmFqVeBnT8aZQ3mKnLFddbgrq55kl
l43AtwfnC9GN9Omi0QC7vmCN04fAau/aOHeB/bIzm69hwozQRQhdOVPb0p9PQbly
yEMZV3ooBVftz6KC0yYvGPcM2f9tz7qlhSi7RdV2E1o1UK2TNr/7YsZ6yQ6eK5Mb
UHEQXzX5imdRD3j/GTZRsjKjmXasxSeY+HI5WFP9RuKK1mL4jIFDGhA4ZVybDyaX
r4uIT9566EuXXoQ1u8ZMfX6gwtiuSY+TEYKsasgHn7q2QpzoJW3fmw1CXbfofue0
ayvnJC742lfW4zJfEngCzyPIXMV86Qamd6kxLrf2dih4OkxiWrO5tYpgigoyvzqT
rKU3FvNUbJ5gD8yOV90pdlGwL8H552UjpvgUQ7lQmQ4pLkokosvKGLfK+S3iBhok
y5/1tHWCakktX4XN0sLLUTdK4IcAbDkgXAGtTM2sxKZ4du1OVgsVWiLhTpdchnRG
zITknllnwyb7bOA2Gp/UovbldAj4f/VUkoAQv2+ek+yyVb87ajdT4aUgQ6WX0uJo
+j8V93CPl6EUZxWDQ31XwLPiC7m2SRJgME5oc8kYCQVxyPNophbyZQHWz7kq9OR0
Iu8eCOGYG2vSs7yPX0wBuZCSdUMSejwPe8yR+T+XYJfECdG5Fsc1kJnv7liqvsCx
OeXtIiCBqDiqQwYfGgFhPb66JCe6APdwI3uwsQ7GQgiLbxMq7f9leVPt4N5vY+ZV
lB8SETLEa60/VjT7sOjtpDvHJjchiL4M9cPvyojvJSQsy1spjdtnI02qc0VGFAnC
F1/Y0J0XiPVzG7g+bv++7zxC4bwMC8VkiWrqLLLpBFul9zyQ2wT9zy7ppam3YDR+
SZ9kftjk8XHGmXIe5c9yrJkL5wQwB6EMVAjv2s8XlPxz+CNKyxSbi9bMbmuZXh2b
7zwrTKZ54OF9+gr8YnRZB+s3BEEEhKzSVw4QR4iTfhd/dJmTC2Qua6YA8G8RTqtX
EHpQ+/z7E12SiuiKFk2gRkKD5+e29n9LIr4iMPi6isWeMEye5vgzZbiYvvWxSNTT
RQLqfXV+lNrXYxKP3vHAj3aLZt1epUQIhp9iszOzlrFs5fDtktU+okwKYMJqPfxu
5dAGuRwtwz9zPzEut8F+ztL/o6GDjYf/09kJtZAYswsZv3Uoy8usjgKPz/ZHLbFW
PrbRvBorEK8vzd12nqDz9TwSTLkgvfxZGF7tL6G+TV6abIvzmV2aJNOjrqKNB/m1
AatDJhzr9/F7pVO5gRrmgr/sHk7YvMNJgSrY/AIebHa3XoIIx7Rwd0QB1s3lWMw5
iFlwKR2G4AfN2DNZvWWxW+U9mZXpgHD41lQ4GxdPXGvTgC0XyYPmSqwyI4A10KUK
8YcmT03OGs6gGtD+io6DZcQOSfWWCXebnrieEzDjqyZvkemPsK0+glGuMBlz/SJ5
qdSAXFzuegrsonZyevOA/5ADZzrJH9sorezgfMU9Clfg7n3fMZRi/cIWL7/wtG/H
StpZvEXRUlG2VsRCI3MKJdACZ83LSN6RGq1MxwOgKkHFInaoZPcwOCR0X1C3IAnm
Rs28T8mHQl3ZIrKWmV3068FZiO1/dnfNOo4VQPrImno+OfdMJ8R8PVa1kwQEt5vI
ZyYAyZIIVo40DNuOvE4K+iUYhde5C4An0cYt2qRZeaekNJXrEo1Rn8Ujw/6uw9wm
U7Q30XA7S3JF+wLCqWlDPCZBEfgkdchX6pXeNQQBDID68rcqCc0Adp+XjPqUoqX7
iHPG//CPAU1QzyfNSPHs+O6de4qH6pJ/LNmhRHbUlsOKn781tXpE50qKoJeWT5YI
JM9vYLjJxI9sDsD00iHGPUQbVxZaAzyTqk6BgtxUsaBLgB0OgtoeeQmtPwbR1Aah
fztgVonkfA5YBCa9qZyJhL/xvCQeJwtmF0V/q4+C+stl2uAF/Yi6EFSoiceTMw2r
+fZfw8oNF9d7+zwjGviLADXIQRQkfPrnqbiMR0tX8yQQoeKKya1wr5McFYeE+68c
DRgiot2PVL2zrcMVeFc9zhCNx24s/BQLKlPnS6NHDkwMo6cwPeAtM6hKjod8BbLG
HFBicq+KhfTSz5P0N86f92UIe0eHNZa6CJUHkUn28w2EGJwn13SxqyZT6BL4kNSg
97Lp+pviz9B/f6zH6yfrZgnKwt0iF0GQrmahMC3xhtj0rXCL7RaU/dO+hO8A/ajv
fHqXwItk75Yn7RFmHliI6vb5qkqBBGELyHGyMe5GllQ+vQYhkse/1xxqoLDAgI8z
UnB4xvl9YMtM73JMijjLyUqBUoY9jlv8A5L8OBm64laopQmd3JsmFC4RF4OGE0rg
lwbh7v5NFsZrG22K656XpmkoFeTXAJakH00miitvKbRrRDn6++SBH0m7QVXSlwe+
HKvmJDw32ZixsdzBNlaZvT69NkAHeS3NPmR7Jz9n/LVXZiF2ufVMKun5rkOQApeO
IqKesnydk8uGOJVRlO7bk85ol1lise2Ppc65Rz48SAPCzlCjXir9seMWjjxsRQ09
TqA9mLHpe+GNDZddy1CDPZw1eRMpEXNXlTEUpCZTXml774nTvx/JpFpeFWAXLgMU
wElGyeCae9juxtTcV7R+dqHoEzqxnNxPcsJhfpzfb1NCoGOVUuzvQ61E+jwAZ5EM
4Ufo8P5Q42RfbpkMUzo5LcLg0igucbGx0mHK3oXdKmDCB/6lqaH4Jf6uP0LroZfs
kuDfmof4FKzDur8QKo/PNeZmpgsYV9yPfOsjkrxg82iAeYwJxJZoSYK+YgULFhJr
Q67d1CgyrBikTSFCBy5b5lkdYB4Rv1Nro+Ybr96Ni8X3YRYVK+aBskUiG2JcWC0+
BBazhAphUWsCAIIrmAjU6aTodwo9+vA1IUuLaEdIkmT9j8Gjclj9amhNW1FUg+bA
UhDLsmnur84ZxkK8F9ki7k2ui0eJysN4aF6VAcSij03rnY9xoS74nRJL7oRw8N4N
mqlEwheg9ssqQ+MGPbpW97OAYfH6iGPYx9T8v6kkhg1IhxikV5KVdpQWPU4S+A5W
DsqO/2P9RJDll9yxXMAD3VDgeXz7D1cvM9bCuJB4kmAuRdCu/SdDG1kAIohXbfIt
EAVlTbstPKasKN16VvU8KO9Z41r+LF4eKl2ATmjop9T/Ys+HZDLndjLgD9UErh6d
TbYoNDBxt2fswl4L6nvjelAzij5eJ+7cDACqHFvRQrlu3cYBB6+vYSY49JRN3Hje
h69rFv2FGu/IP2Juq8nitKsvXHyi+8fD6Oeo3H3NnD13VU/rrztE4Z7gpQ+0n46a
2D11DMmMWCTqV6MTEXwHllB6fHuTv3Yyqgn034wylz4ned3speHSAk2HZXTZTR4y
p5NKjwkx7Eylbo0Y6FUon3R0bBUMYEyWw7KmDqcwAqVLHMLBTsrxPyrZkskCqsJQ
lYfbP1BiOwlQ2KXPzZsdXsg13DeSJbfYDObnaxLbqRMZoEGnihDNCODDvc2YkLdS
QJnhnvQIpmk6w+h7VMcHLdaVVku945Bctw021RJfMBAFzCFjGV+bkB8vGuMzVU05
UuRWxBCLPJdjKA1NvWQHdYJZcBWdWSdqbfeKYSv4lYZYe4VEWFCfoN6+cM/tCmDV
CK+GgidkTwIThogOKGk/jt3pROIeAuXQVwcXTsgA8u8hZhnQs273L/I2QxgcjH0g
UN5DQ8dpXpDEaXDCGkwpXHyGkHmitRLIUP+7o5F9MR81CB/MKsUbPi7bk7wWaKzM
E/qdL1XQ2ULvEGV/ilVExWGitRh2+J+GZQfCcepg3mowAEC3RiudwppcSJt+2R2g
bEVJXELPOa9RSSGfeJk80eT+M7UQshTkj8FhRyGGIurHKaKVNziOAB4ySsUUVxsC
aEkE4jsZKL9LNLvTG2BmAaIbVOfl0cHr3YC8gew/xW2nRenPnvm5DVeDzwoCcu9j
kRQuoZEfBj2GGxtsG03xBzlrbK2kCsv4VB/w5MyQqrVFHCgWQhF1MpoISZvDQv8L
TDdnPk68aagO60FxeBH4cYpcim10M5JtyOu/ZbotvkWpE/1JGN1ycE39CDGsZdhQ
GrixGmlTr31UngrvyxgMPEK1vbYb20kQhZzCbi5f5KxHa6Tl4gvQSzr43auPO3Fg
AGM5srt7Hwzz+CijeW82QKAr6R5BPPJc4x4HRtksC6BT+f4GB/XiDGWKPNJYV4li
rpxIRbeilfLDgVWf0g2CYy8Bbh9KCxrSKq4bArcn1TJrKS5hncbL0tXPU0fBemuK
P45muRbN50zCYykgQkT7OXod8ncQe5Gqo8Tm2Q7hxuPcyma4dogtdf8MOMJk46x+
MiXNNpNsg/NPhVwcRHNlV7FeXtB6g64LNnSS811LQaUB6c1AJzDyS9O5x3iwjzVW
lzELt84DeWlnvSwz3ZESNImoLqtyZzevIUfrWp8Tum+g2Ka5W33dp0+HUZBaAWwj
fAfXg0Dt/QxGuUQ02FSWplp39SN7zothRI+10mGHcfnv1sUxJ3GYtm/tLlvjqGG7
OaAJ/JgYYFlVn+zbKMCmn8bPDE13+Wg9oecOw1hLfgZlQNRb3exntwfTMSyg7aLQ
E2GmxLRr247UlMeGPn9hJ3S/lGetWm1f1lqFEZmqD+PJ3+s7KKvUPuz9B+T6ADqp
szC2FPp5W3ezGRSZYHLC0DEV5kkCXJb7gIcWpECPpqKrrQwf54VJKIAzA2TYkUvy
ZdaQqk3pC8rl8U94m5jEiG/e7+yFbbQ0wIGKohH5TGC8uIdUHIZNAbmL01sXEeJ1
ZatqIJTbRc3PurQAtpCtobWxq7CxYl2t7ISWM+BAG3+nQC3CjPkYMmoa2Mc+yGFP
5l2k0lHzTPKxSSakyxuD/7vJYfvwPwddmoKScec8zpmHnPyZfc3rv0bVRyspPovj
QFAwCXjVv3JqiGqOK5yvvLrFj9yWY2WRsLL5Rvor1uABDNFHtE13LmfOGNn/qumL
MCwpSy5tyiQUBOFIIRM7RLwxSO64uVzgRLbOe+S9V++cHqMsOvK8xq+9SMrhRNF4
KRjm1xEIx6zyyx1sD5ZryRDcqpVdjKAhdSBVqaJqgcQzqQ21g/WFT/7QgwmceYWl
BaCr1MYEx74NmdemcD1KXKL1bRVrJu43fwoNCrWGW0iaCjgLruDZLA0+1vgyxPTW
`protect END_PROTECTED
