`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3+JMQOcgqw9P4dNfWhEjtNSOtHRH6ebxcih8JgexWkJo6A0iu2yQN4tb6FaTgYQ9
yjp/X9HvQY6oFa96yJCJAfJ3lelRNzZONwxZnakO49Npvpr76cFSdICWI6FI/lQs
wuWBlOpe9R4SqCg86UBtQuKbIDZoXiBK5wBAyne836Y+IfOdqU/NOGs9U3JYv2Xg
JLvASwOuP6uDZiszpBiVHT52zpMM3+H3oTxKgYKFq6hXmqVruv25tYa9ssuRG8H6
NhifgBfyHLrcZwtGorZiLRoTuCT6k7HL0ZT0g3SwLIKCuCjXW9PTMAweMqLYZaeU
HEsvYSfX5SuBsoPRceeH1GN1mvqKLRzOa2fLOqyKWIWalSgrGoh207hYaN8e51la
1HL6OuHfAttm/pr0bHQjc72t6YTRK3NCn0SH28+fXTnLylpZCMzuvziLiRMp7FfO
eKBPnJwirmLhrGf87YA4eHTtINJzFQ7BqXpzeIzmwEnXcZrYjnzA6ArrW+RZcf7v
liuo20AmmLfCJwPybnzHR00Sv5+aQBKAcvZxE4hPX/A9bW2i1EHNZITtp3up7XJY
BqPOA5BWdCLuzpR/zJRLOpLLuvwJQW90rRJ7JdBqVbMJXDOfMukCtxzYz9DXfvnG
bXvw4aS5MTMxrNglbXaFvMyTwag038LD5akBorrR0zYSWkU8Xvs9K5b3MgfmPHPm
OJtJqlJGigkRdyiala96p8kPK6AwCEiB9E+akMDWf1pNumtS5ZO3wMgI2f6mFJ8m
lylko5Ammr44Ug8S+Yghy7MFG6R4VF8bFqn0aE0RzRlg677euR87qoJL/k/phFpW
JLbQuzVQ4dVmHGTlJrSIpNuvWfgY2mwe9QjksetxDTu1UL9L9BQqOJP1wQAmqYTR
y6EsngmekAls7EI6FabX0R3qLGsacDcn850It4jlSQlNG5L+8r93KWr8P8Ky1gsy
/pU2/gVtKa278fo67DelPWy8+7CTe5Tr6Ez7bY6b1yPu4W0SJkJtCMQzapNOfgJc
inBN/bz+SYLlt9kOT/a033pdesX+04giF9oHPUXYCUbRZwrG5yBDjZ0/2hHTbnz3
y9zZLduDVzhdi+k5WKgD+tVqsmAVd9h7etIf0o4Wp+iiz9snt1L8VORbU6viqOYC
oK6KrtINK2vTNLz923heIKW31Adj9ujN5gbLJUXq/6d2nZ6Ng/G6vW+FIHIg7QOh
K5onxSAIK5F++aSw0mHRQW3RRLQNNgLvu1yTxqO9Oq7SthlvVs0rMSzfZgjkbALZ
1A6ZMJFhU/GTpRNBNtxQIOgQGLQObJCtSNXDHrlx19uW3ZUBf91XpJEI8sEYeu4P
aJ5IFtq8txQxMQwjRLyRVAn7SMFf/7txVvR/EbSJk+2L+eRKeCw+4IfkAMgPr9S5
A4C8SkKG2ZTeHfD2mk7+8xJdCHaLW3JoQ5v9Y3YuFN8w5LugScdyphCKxbz2+z3f
7C+KoarYNQaOuonaYIWjODUoz2XV1sLwkLgxF6hpZnFHTx+CqSx6vEz2oHm2C0eM
1XzpOFAfVEgXNFpEEPi+XexsIZYpZ6BN4ku0V1Ra/5c=
`protect END_PROTECTED
