`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3OTQaDxqmzYRfBIycNBmZdBQNXlysjZmZesawUPY8kHhMlmZ8vLOc7SWTEBRW/Ct
U/tIvE3RJAnmjWSJvjk6tgbbdyb/e7zhqLynS9zqJQ2PyytHvJ8VtaMCIDxN3zIa
nd2mH1nOfR7Fb9p5bs720H3JhglxWPGYx73D2ZJzK1CwFBBYaY9syeb/QO+gehPX
iUkhCV6JhQoRXnQqQdNLn3Nc/iEvs6NUd6CFTsU41fUGakruzXjryYVxeBXW0uRX
0s4/q4HsALE4+aYzoh+1h9I8LrlZneT92SNDNuy7v56LPj6hT7Nv9qDl2v8G/LgN
rg3MIP5TtyxWMoXNMSkE800Undw67skvTTd/uU4OHvvoNl2pA2pI/217x9mGtcg2
XBuD8OvBUhTH2u+YUXhJu1tT0vTZYYkO9KBUZr2KIGriekhz7N/6E6Ids9jTV79g
0hQfcigT2BiVW9rEPR/ZcRktj74fK6GAXX1d86qBsZy5hb8bZ7OgNIPDA2bFWncv
vJXFZBN/pAqx/Gsy6s3yG9inVXXRvnXe5MBc+TDSjU/DfSJY+lV+5C1rxZ3KlGh4
HT48KFi87WJXUPbpApY2lRDVNKn+ld1JCIrBX7oBQ/krOgG59itpyPLhBTsd9hr/
QhOpfq1YbGGrfnTyKtAlJ7qJ7iakOsoqt8YdkqMp+j98tUEvShIe88itgVcehyuR
u4kXnqL31D/CaWIFxkbdWzdQChf9rOLxtNj9GYslUuutifKR514AEQYi+EDDIKtw
9ChXxW4Wy2WEdFSIK6kMBVeArEFYzQtRkELrnNulQ828UsZt5/t3CKRS6Qo37Fmz
+VMo4dcPAcYcAULYxSWmi/4Gk+wfTar/GquVlaa/s/WvVeyXU76JqCPOMFMb5NKr
msB+T6ZDCj43FLZ8KTBFIpbiBX0t4oXdyfQTeTdMb1wTIyFs2zt2SnQfLGowbez3
z032DkxQfJ6LkVDQdPt+fb0n0Yai92/KwoBJftnJodhEfvBqFnU/4tsWz1Q8QIGJ
p6fRp7xd7vZqK7gBUenrS/BA849tDvGrV3h8AsNeo4auHvOLCN4ogn3WLcqlloV0
vFVDjT4igqCaQDvOIvDe/XBNad0dWj3TZy4F7NYDUv+TgW8GEc6sjQcPYxGi8L82
RL3pOPwHyYxwq3odSOS4ceMfLDrgXrD9HD8mgzW3ysgWkyKXSSPWa373I8uPJPCz
qiSWjTYbsgGhSF9dFoR5yEQxzFw/NFuem40ppao9oiYLZ4bxjRA9EiS171MdmVk4
L0b6C0784bS830ewPrF9Wi+JU28eMutUmCtxvWvz9bI71o6dRgeyYs1MWCbO7i5W
r+/rxl7Bf+lJIXjp59iI3zmsX+x5/TK9qv3GvNbcqnFDu6Jo+CqOwjnR5EAlJoyo
jbewHRIBn4n89k96lu5GBRoYJwRk9r9addsXJij0A5EVl2QRPLR2B1XIfVISmbHl
2EHCGwkJiqXbaPSV/KA182S+ypEg/8GACVfKSGIKNv5BWQU2E+GpXNYpNqQ33+zm
9GaoNiDvfMDFrBKHSJbJsR3lgPCRlg9Y3WPMFY/ocSbqZj4ze4f13F7JLbToPQeR
jY9UDZFNUD/oNFMeGp23i9g7sY9JiuSZ1ei9ukxF438lSYE6jaokzGHSZz4AMS0X
OjsCELnsz3T2ZQeaY9GmDdqNdTvS+RsCoVqC/k31iQtFSJwBs119qL08Bm6fLKu4
aHB99aBp8JNTkfb+UToSNLeqsd7Iv3aQ/f3VW6HCcuc=
`protect END_PROTECTED
