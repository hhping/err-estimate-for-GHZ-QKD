`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z8qEUBgas+7h3+07Q86xD5nDZtS8B3x0jlhf5dETmdw7paV2qDmRqj8tVC+UXovE
hq30LAbdJwV0/TiDLru8OyZ/PuT8Zi5bMNAMR4C+Sg2yuyvY/SC0E6T5bQdMbA5E
+nWW8SSb9vgvy9ddpWC6XhU5D0OY4edPYmH35Sf+eW5IqL+TdsEMeZPtx2u8nHj9
Lo2EfmlNu3JunIc/0Ok87sRZMSVZgoZWC3vcZdkfiRWEhdUkdrDd9AhIIB/kq6jo
Np1JrHkn/Lp71TN8PUPnXNHFuOI3uEmIqI1pKMnj2EYFgcq+5D9mPZw29GobPwbC
ZYU002A7XOLAVOfp9mqHeOgVj0tpkJvrSu02MQXrsWMupgffZBNxkqyClOEJAB3q
IfSB8b4D+EWsF0XckzIIyWnMzZu3rznrpR5sez3v4mCo8WXKWrFZImD9bbkaNfFf
T0MDodU05rSK96F10aOMM+V2dhtwuVwQXkEYOYaD4o9gbnfZ6SQvjuNngd0+0L1z
azNLZGWVv9/0+jVV72cNk+cGkJzapKjmBS7AUQD1LowZQODGyJuwckiLAaJ3GG4B
Rf2wDol4V3gz+ShabChqs2EcIdQmwtEDNsOG4Kcq+ciFYdNlP6MW41aLNLJ+Tyzt
`protect END_PROTECTED
