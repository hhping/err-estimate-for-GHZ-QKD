`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2/RGvWR7w34mU1estkudr50sV90xQTSq2auHEHk/LOb7x1DAJ8ybP7XiXT+GRfrg
ap9xzeb4Ys4N3PVcOeJ2sGLHtnLlnHO5bdA+K9112umaLuTsp7zq/2a+vgv/Cyy+
KkT+9V5XCeQhnEUtiWBkSEOKrFho2tF2hnP3QZyF2tynDYEkQ3TRjQwMFqJl9o4b
engT75tPdIDngSVqIjonF5p1ghs6fecOpa4NolyNpBrrCwRKUflCfugR5r9sIS++
uWwWbJSGFSZwJ2Px0BuClJZIXkGzW6dvxYKQhl2sfEbzMTqOZx/pkxJtLfTCkbNu
d6bt+Fy+3k9uxVnx+6Hgix93pljMDstrFI7AMnjg+f7jGOInyXgQ9hPU+47E2doJ
OMi6CpAMasH4mFhcF72DgyPb2bdiGGVdO/PGiouPfTDMhqvQAIK748toGQbUuf7T
SdrLeHfKoz/rlyWzM/5CFYzJBx/aqCOBzpywR9mgaCOSEPA2lO2FxyzxFHZgpbs/
DuwCKuTronVNL076cV233GZN5xtLnd/kwN8yPvEkgkyv7YrlUDyuMjsJO1Ten+3x
Ce7CY4B62G4HH2/pVyzo+Gf4GdMCn3yLkpuq3K2G4wVwZELn4YmlS7svYXjrzSO/
h/H8VPdawaOUlsB5xTnK1VdAFhTmzKQHg4Ton0JBci/y2s6iJ8CcnaVYHIETrak6
sRnWzve8nCgiBPjGjlMFri+5btCMLmB/2g2QxqkKO+kGA+gXzBQ+grrirBVCxif8
CmnWmkIaV2s5K9fSSIa3oTsm8AjQLlkhPqoQkEDXjgJhapFsQS9tHMdciY4DoIL0
XnmivsxZDcWiMfne9YTZ4Bu5R3Y1BXzKU1AaDSdKsazvjEJ4V3+8MTv0NF4zs6q9
MEawtxerspSoegXlGlb9qItu57xS1fPNeRaijSpQlpWKRwa10o9N2DWOM5zQHlA1
eMKYEj6IOI5cVDvi1ayGmV1IwPN0Ijc2xXkU0ge+eM2sSBVgPMZB75BL9rYbHWbs
lgEutzyEDI+SAKIbOKKmtDoPFOtYwfCN9M339mTfGj4gQ79gKkZgbEK0mV8qrKSe
iXfRMi2+iVio2v95P9Y6UMRKIOWXyqNhaXOnM9NoMiBLiva+poCZWs9e/1uQXX1+
KksafsuUAWxQCwtrIUACt4DPIhFBEM51qBez1jkCSwQEtavMSrz+4PsSwT3FQN6p
cPHfFPxntHSFKdAL0oApx7m6Mb2Ddb/31A8rQMvgGh4jIZMWh32eEBhmjr2UIP5t
cBENqQuRglRw/K+qnokd+BqzMEPzYHLvmzI9WOH9rQYaHpZ0TlwQ9XvUDTADvqdJ
`protect END_PROTECTED
