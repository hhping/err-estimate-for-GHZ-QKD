`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
41JwVY9uG20Ny9bNGMiD1sbfRBEsbi4MPWUIpy9qk7wpFRF8Kx1moMmOUcu2m5w0
8aB5tXj6Fnu+g+dJVKK96VaOOuxzn3t1I/JQDLaR97q3n08O2BXWuHFZxGLGZRNU
EP2ex/8f6uVqsX3POQ/VB/mJ/71DQI//+akQX+iNJX2E4uSHc9vH3v6i9BPRmuVB
NvV9CfCNQFZRz2EgoKvXemJRu1KaGl415KrddxxOugobjBUUR7TBMqNhbPV9pRmY
rEr1N1ZhmVSmxoBM3GhPGWtJ/VYZCycu6CpvtxCweoOHDO8Trp0q1BoLdWcvxgIA
TkXw/yncBrB+6NVBQxJr8rFW3xaLU4z3Wseizj+1QpGsx5hNMGGG5mDvMkUj8dlF
Xmc7wOMpaAQdNhLWwe6rqVnYe81wEzESXFdlNmDC5/pRaF4niMoj7IDh3kxf4lxm
dPYQCRfQT7Japk/sm6pAc2Ry7Bv+wApJDMfUbYQNOZxnsWEhX7fC231USkN0noow
63RCMCbbAhcGKB7W7nw0FP7gWNOU9ATwNv++RiUhS2yVL+mwopAcyMr50buDXiYG
63Yim3hSHOzR/rB4M8hQa5yf1KcvoHHng8o8QrBITNqybzVSkFE4Wwk9tPkFlhao
UcXE9Rix84C+/ReHH64/SzFxIAQyIqn4tbT/yK2ALIsBKjpoV2Fl4y0wdaLqrd1a
gFR6YNLcAnNnsiG8XndpvDZDGAk0s6myAJ/SKNZVLthh2VjnnQFlgYCnVyJbbIpd
BAuMg4/O+yZcHo1hEjFjCh7T11xTrF3D6oSoyVI1Kg378dCyJahHMHkhaV5Lg5RD
2OObEUJm36/owXv5jFejZvC5bbzn4pBQELZQ1NEB2PohJQhm3rf0ruv9GQvgGsun
tf+2vigO+wIUZ+i/owRp2y74MFQMGd6wWywSAi+SoK5Ym+TQ49LFO6lB0l+yv1Ta
fNouTUM6Zgc1ISsWbgQ4XGF624wNPG43Vzlxgodg8mtuy5OFbDrmT45d+qfUml6/
Sgox4/1bOsarM0pEPFZZxtqv3Wz2mEnZS4HGnaqfiSrlx35u/1+BV/M4fAFNQ8gE
Oxglwsy+RqCEjxUXCdpYd3RFiZuacoyyM5W1kxyOU5UYaRVyfNjKYlE1yF3l+48v
9IXYiISOsXYVp2FpCLNooxhj3MUTL0dtlDr7u919SMz7kA1dGWlWyntwYRgA/CN0
RE+U8FbOCLKSdRX+ziHNW9AqtXmNI6TQgpeUUnp7txZNVZXeltLigPdZOB2KstYx
x/Wev+ymaN2t9pYLV8KMHG7ssD8h37lNPIpouMd5rPkpGN/CQEG19uEpWlhRObUX
n8eIlJpQaXQu45ZIHO9EU2PPyy1/R88R1KVoEQC+CqN3qkkYztad0mXdDnzB3Ku3
bLGnxJY5G76z0AgxWK5Rk6JVXElQmUxvzSuPrODFBI2Y+JHrworhPq3fDA8cgfgu
CSQf9+uUypZUe2TmWTQzGNu9K+flYwBMlKB9xsZJsVOKLu6yZsyFMObwOk8PvAyY
TfGZ4A9kLf/TCyGFNQKh97UGQ5GfXLdN0tRS5JydBFTmdE671af3HlAC3PJeeyWs
mgruBpLxHNRhTChSvbttacB+x0VZ8I7y7tkqbCyHfv3ybVe0fRRteMtCSbghkpjN
mz5diseGQUFqcu5QO94eHY2nIiLXgDTIGHsu3C4p11NJeTwyE+iydegumwEesnmX
AT8O29pTPsnnY9WlpGJCo5uwg0+xR1vft+rQ08dPcKDmhH3fjMqIYvZdkHwHt1OY
g29bS/icXC6ejIwqruc9MEHv6pdULdTrkE4Qpf79m1InD5Ksb+wRV1LgNLMQTojH
sns8khiQJgZKNka686i78pClENIJh4cvp0MUWeOiHSjd5916vUp5RguQo7fRhZIi
LXPpHg2zxEzXSSDhiCVCdC/SIPLvH0CnYsvJjDaujqHatynW2s+Y6J6Q7mtVA3Eg
xBBxhMCM/ey8z2zD6pOMyBQJyyYMyJfoIhr1dv8263bO410lbwdq2X0satc+CKo5
RuEiVOX5I9GdF3YGMPdysi0dVfJdmCNJ066mXbLxokyhncPDod80Cr3i/i+jXW6r
DEfY+dujc3kfS8576Nq4KI7zKWdsCu0jXgA4g6xhBBewZ42QbTazdjuwv8z+KC7T
98ySMXrO/7tyWThErfLNkU9hLOVj1oBajeEbuSEb1v5wuK3wj5Qr/A3p/Fxk+rX9
tz9k0Db9m76Mb1XNeqWI4VF6cG4OqFATYlmRy709sw1KOO83VUmsT1XR1P+ANxcE
hpYS4DsmNvIw31ti1vcs3v8bOcNCi60Cn9hl5ULGVVC55tZQoOtuKGBpdt9R8XkF
5PS2o4j+RtTr9EJuWYIt/ooVlJtZwHiO0qeTLpVxpnFmy//+ULXJoGEsMTLYwUMt
z0wyt4Dk1iERLd251tpryJrizueOPqk/qUZbiy9x29R1wC8PHLYSZlvtm3Jp0sPi
rPmw6VmW0ErWhgzjBAKGceyb9/kIvtObK+3P4mPUxrf+x4qhSCxttTPlm1IDVvLi
ouNRzzcxeImMyDITISb7nNiwcXIFAuiGprYJw3Z3j5tRVhMmGbEODBq8O8uBkUXz
juX/irB2VoxGoKO+rjq3P1ehjV0vV3WWR917+6yRIwj3kcWMs4WvlAhVn9sAvf8C
1H4boWSiPthrcf6F+gnbBYKjJtJiQEexWRqUdQf7GMxGpBYjG1qFac1DWisYmJxT
Y0M4sjHRSTngohs1IsBY/vtNKSdfiBGP51GBI9cdCuuwwgCtf1tj/lQY1q8RpArt
gWHRrIWqsoui4u8JsLNiSdNraaOTMOLDewwHxkOEp5EPYrNLB/TfxVNTj2b4tXIe
g3Dpnyynoq88iVkcDwZH3c7SFHjBAaMKvHeJrZ2zdU5aGo7Mu13NBtbk2BdWuzuW
7qDuOjAILhlytSh45zLiwHjjl6sZuCtzoP9IWR4xWB3FQ+B5rTFY4sdIJSET11gD
I2Ps1NBFcoxRrsxq4n7jGOYuOtXGuvyndlLsH7pijoHxLK0V27oIisTsFDn74A09
7vNBPCyWNL1G2IXAE3MVn3vOdqjRfkWJpYzJlVWuiM+9nnDEUsRS7AxGzpxhTNM5
1dmFL1Mk8TWT9xnMeR6WuXLjUMV2dRRYu3pKh0mChyW6bGSJnJKVgG2UOzPpw/cq
qEZ4b7PcABU2QuIeEq47tRxv4kidOuZmVzuBb97ltwEdZSb33xJ3TLJOkl3XAP/R
`protect END_PROTECTED
