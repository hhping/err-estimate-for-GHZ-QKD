`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ylNDIR/UKks0UVFNjVmB308LwJedQ3Bt5hVZqm1DLfkbBRWCYKANonnymE9CjRNb
4zPPghE7huzqrGlN0gNev7ShJHNSEk0Mg+8CXxXZc9+BbC/EA4sdZiCxe+2pZ47D
Y7VRAqPgvLRlEGwsnKDC1JSUor9y88gtPqcQkNBdMXG9pylLEz+1+08VL0sCXCyK
PNy0lm1ZurE3Pj3Y1MEMWOV7u5uVTMURQYlZoTvb2qUMCOcTykOMdN/X19VkeytK
J3/BRRYGQruc+OobasYVtP3tPDhm4pmVF+ZBQhQkpTjmJz1Oew8afbjOyP2NZ1wV
iYuH0iWbE60Fmc03HjXXjqBVX88j8ux0tLX3trpT2PBajZP9d9PRLQsOxL73TEl8
tk7uavm/k6Iv8vVR4LPUmcF5BxpPCX/W4RiCKDEDLMaPflKIcW9EETGU66MU1IjP
2g327IExh4s5H1zod+ZipgD0X/+mBffKQleBvW8nbtXJqScZshPKckLZ3FHrgyHj
O/g89BHdJTxQrOYz5jLGu64CJ1vn0xGErPQpOv+fjAE=
`protect END_PROTECTED
