`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2ESmD5bNT8KxprS87LaP7XQfwy1cLf+8O60ldj+9HXGZZGxBwVBqIKiWUfwxNSg+
EFCxFl1k+kK/iwBlkzv1TRFtkwFJCFhDnY0X8b2fIopC1ZPzAXY/oh5O/Qo4qL8s
fgJg92GnB2gyQmmW0CtnYmUv12qqL+pR4fyeiqLJXPuSPF33xjjUduSu/EkPy+kY
oivLQv7Qlw0PyLU1pdAD4ZT7JjbW2+SZMcVjx9Tl035m9Qduu+ih99jK90k9p/XC
MVRDCw+zWLAcV329vFdZLwH4tVETIyFmqw31eQTGR+FFzGlrOJd0N67eBM+2N5a3
w+NB+6jY6bhGQBvnoY90Fpn0DKKh6s/98BrEkzvt5BMz9Snh9BEgjaWFEPXsICY+
JUbbdLoN7WQsXOTx4UoOOGcyGrDSnpgAlGgf9v79QqmMdDsehWRfrYpqTV14P43F
nRwcHsMi41VqTpXKPfVAuPOZ20M63uWFbcvbyQ42MIEP8bZKm68V048+WMTLsO/M
4dEQ8rdIa5z506rIPzJhPCnomOkWoJuUH5PREoZkgr/NJHR+Af02FwTOB4jcJBIv
`protect END_PROTECTED
