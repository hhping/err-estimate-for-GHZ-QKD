`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mzAaDpw5X5cJfEtWnAKeZqBcplcFKspdR9ELk65/lPcDt81Fk1+E2K9qonMU7mIT
QhOlZvbUOWVGAEv4ZYrj4oUpvaLf56abkAySMTWZZLnp1KZb6idbtUMmqEqBliQX
f6izYkxJgUPEH71CijBuXnzcL5uR09LOARfOhYKB8KUK5cz4Lj+HOpwrn6H48Sfu
wtg60qMw33v1ovMR2QK11nkn/4EHB59fGPDhbbdET/R1U/v/GeqquS65rCgquNum
YBVhqmr41VWV/SDpdl2iA0eD/hLQ4xJnVpLzYgf29tSfD1saXg0mMFClMYFsKDH8
yTkExKjQWvS/uDM82LIXlSIFhWIRBMN9hYWMMNCKjl0ZG/UPLHOvMrKCETSEQ8Jw
zjgtBwX7hCal4L+ZlmIj6YkzzX+/uCsGlNITF5NQvJ6sLSJvxvNJiIS5qx2koAkE
SC93f3sLgR3kOTG3hEea5ZV4d28pr/zbt0BlzzbRmVA=
`protect END_PROTECTED
