`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RKEqkLVAeEihsfjjCEec/pgg47AcofXiy6loScmpjd+ubnDRZOm1zm3Rq2Y8SeE5
fZuMGzythJSirSc/7A4rrrzpTDmZCd6sNPuQwS4p0gyrOlR878ZLpVmKukgxqcMy
1NdRqi6Ijt0FmGewo6P7HQszQLqh4J9pLwotJhvZ9Lg1vF71e8tpCKKbagbhcbE9
eZvHOkQ3FXel8c6puAncKgL0nJ9nVSVCOj86SuxAXWZRgtun1HQfKj+8qANz61Zb
NZ54Kl2c9sp57/GweFEHJc+WSiBWI07Auty21lTJI7XrlJM+D/uEmAVqiNaqxaYH
+UObW3OK/ApsmtITFHpyqcnZkFNF0B+A7UkgL95YelKVJNGeuVYr8FQeBE7e88WU
6dPxkX9qljg3w75pEysmubcxdVTE71u4M4SIf9M/A3gk1XSP5Tc4uOhVd5Yuc6C3
m77wplU34hAMYmvD3Q9CgENeg8NU8qjSQv4MHLNhW+p+08HCH1QXcGptBrX7v8B6
WkxWJ6u/j4Wfcj17ArGQMRRt+X2Y1bp+MO2XpZ/JAPe4+JjYuBjNBidDOReko63K
bRyePSoIIk2QS5uoGZ8+yFDe66UqKHt9drY3bTg40pdpdXFkRuW6/XB703NuKICX
rqwdhaZYWHCmtmMtikoxFBBaHk50D5mZaRzeqNkJCqYR+yhUi8vmpV+RwEEaSbPQ
Pu7rpEB9CsV9hwhwl6uQkSbHlg6Kuo/USEYUoZ3Fo3SAvTmcN0w9H8eeAoZRKsDY
0ZqyzrzdEB4yiURmHX/TXspvkSQEh2qqjzsSk4azt/Vsl5Jgie7BlC7Fl7AvFhTK
bnG8klC2oSC2qJ6HSP6DvixL7hVR71HUxY9IvfRyPSOR9Ki+REDMbZC1wf/2KPg/
ITDAZiKSP/77GXpj5Azu2+QiynYDdEYw9zLRvBSrIpcW8aXne6dqCPJjKvs373og
+FuqgzSGdveXfpPQh7uJIASJEIfM0YYSl36hd58J7YqgVSqmRjOi2anYVIhjlqdj
aJBJDD5ubrNE3B+quQbuaE6ZSSKRDA1HeTXwdTgE9ZNr7+yb+VIcZQ1qICVRbikj
LlkajvSfToq+MwX1db3yCL0qYiu7aeeVrQhHxdtV5RtanJR+zY0TRCx806m4AUTX
ez5LBbSyt3YHAFHQusenn8QB/+dPXEU4REuJEky+Fo71d8IYp2Iu2z5ak1sUhUOm
T/6HfjGyR7SEzbP+NjQ4VgzOgrpQxuuNYUxLVCpuT2r1qFVbeHxgVnm7mX3cLEHw
j1+hMKp61MAk+DSRb/R6gZY/xd7OkYe5Hmhw7ZGft5mBxtpEZ51n3sHYMfrCNmMc
2jE2D6dPmrbo00MB8AGqkdiR0aY4YTQZanctApe6/iwWgMjmkhjsBy4OGZdYRMgJ
XxCq6IKwxWfZjqMeejnlk/kzTJ/UIxH1BdIYd6jL5Jxxvh9OSqbKIcFnT+cCIn/y
eyFHitz953EuL2ktrLZHh2reqdpJWWIus+EV3/VdyOCpS2l4pcMI0Q0BEADcGVLP
jJFXKalHLO9FRZyeuMpe6fOdiksX+Mpx7coXmm1vuHAdpbC/3a7r8aB7B3/vWpCt
3JObeL8uKvLy06gCIHD/PgLugG2zkmY6YG6RAXAg4PamG8mHT/sp+i6e/KKSP72A
1mssjogCubVJfDabpf/WyX+oz9INemTP3j3NJsDauGHC5TCSDEMNM/soDqwHxBSl
Frb87kDkjM4Hff23iAvpjRKDLmVPap5CC+FqgLnb9w65qKaYjr/6Ty/jl/X/y9+J
hdXukPE04gsSYkbFfMQv6JuflX2oxXr/7n2UzArswNsaHpgk2yEj/zhixeiAYCgW
hi37emg2DpEf7lJbxHzsH1qXaz2bGpUiOUrrpIqw8xLwYtI0Kqkgtn07ha6OmokN
EetVxL0dHdhiQoPa23M9aaBt++Bhqu6+TTT84ziOfVvqDjM8lL8Axr5I+oak0Ded
rxpPFmXoCFK4JWQOgdu9359RDmgXhmVX7a9JS7gwiE9X0r6SKDmS1es5P8lM4Ff/
+v2vvN0etJ7hxIbr8IMA9OOPPcFTOjxQisQyXnaR+BmsGfTz/MuBSj59e1QWxyPQ
oF64GVDh+HzD69ucutNV5pMmi1lfwrJjQbqIS5R30lDfv0qRR27LbOCdyin5Y5kT
iR3IxLaB6KxbPJBsut5X/nCgygjXwQ58kJoV3DglVCppbW1fPkOTO2ZuA3ny9ImM
DHgwj7Ahuxv9wvwGE4svdoqYaPGowIDtYZXnvRj7SM9raBTKakTCYwE1xskX5ujV
+kyaALL3qwHHmhFBEyb48W3qVZDmvPN/f6f2dP3lziY4pX+ajRg8t86HlC3Lc40D
83EzaMT7nW0m4kv/KvkP8/b8Kt35Wy3DUBRejMznph7nmpoQStfGtqT5KhT5ITs8
GBI75WMANrI85k/UgyhrM148qunlQKVy+RNdsv5p9gGTiqf+WvJ6LSbYdqd8vFFl
xoxsFKlVN6oWBxUhT11TDEFjxKT6ratqFyuXvUeWO8i6DeJ2mLWlY78i0SRTQU2b
iAgLIYf4EeVLSFYKPHzEcx+jGl+QqqaY5vCcIZdyroVigSEAaFssVmxSkfx8ay1h
/JhaAUDvUtZSzFYk0L+hSF8m78EExnAhq/t2yUPjBXH6+EGKN2vWECJZuhEJtWm+
`protect END_PROTECTED
