`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MmQeQKmgw2s45voQkQqi0cC500Imgm4iSOcOKeiGRgfDxOoc2NiOPgJbyVCUvd6u
VrQ/EvNrYfV1M1NcVxK/UZqyHb/5hVifxKyFT6Em9VEH9qmTQyB/Db2HhPialMom
HnDgfaIB7BDBr8p9caCOuyoRxiHLtvjQGaVt/+4wXU/dQ9NAWk+x8tytw6IqkkGp
9AHSwLbJL+/4N19UdmxJrMIJWN49+AzD2EcAu03mmWIXRFeIE5yyNH/uvMvwFiMH
EYjvlmDS9GLuD9Ton/zz9q3XKcQOKpN5V0u5WI0XHCYAKCaiZxJPlCl99216O/9r
ENDP1wV91DIVMrjAXhfZwLsiXl1tt/qqtVA8+allV+J7HabVhe2n+akudWmnLPoa
uX4WOXiRaBQGo/NGe4gvWt89DhAD8Bigg4fok0uNDdOr/UQGWyZjUF7eh2I53D2b
buoyz7Dv3CU9PssU7N66eMa7EJkVhHc6Yjpn+TkJfksc/hn5olGOVQntHTs4d0RI
dAlxtmnDjOROSQWLx5CxQRBxryccXoRXBnOWml37zuIRtxgWPMz0JY+g/4aDeOnN
j9/txJ5i7fAwfVGgDi9es2LeQE6oTTlNZJikAtXBn7JjPO3RcPXjdTypt3qU6OuH
ysEWGuMw0iKRhlTwzz2BQeic014GOPT75RmDXnTp19UPf97BQ2Ifxd6nnr+333Nd
I5SJ8qnjHBHvH7uzYnRK2FVRHOftiFfZeFtOf200Pnm2unDqBmJbKvpCDJTRrfUE
OgyogGieEjDfrf/JT6hZBDMayjTQYkPI6yBBQNA9CGOODLX/NMFdYSVfex9SowJF
vgY1tcUAC7KqstPTYUJPQSDo1xGrUrYbf9IrBrNYcOb0n5vIRYyyVUe+CFOBJ4SE
ISYRUySQW9pOQ+J+11FeL1qc/TNJgGGlcWNP39C3l29s5UrEVyqsdqv1SABaAvTz
zzmbzuzrq2sHmbPqUwcILlu7VakokbXmYqD//lYobDjhU7AyNuljgPRx+EQW3dlo
1jVxbNti4321M0g3cJezpYDYqIXESmyazO9gNFlIKIZ/ZlaF3Z3mRj9ZxMNDsejn
ypJaeS6nnDOtlnimVv+WGs71mhDUrBLfG62tzZRPWPn2ilwl5kfvQaAuOhQNK76P
ZkG3xW4P9gL/QOgSR8q71+StnRQHVJPW6InZj7WEb0fNjMQEIBjFMtorcMKmplS0
ofrbE0D6YvaSU31BBQObWQ==
`protect END_PROTECTED
