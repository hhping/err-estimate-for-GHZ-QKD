`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hi1BgVzg/1OaJeX1z9zFDvb+S3MeWXqAw0I5Om/VHhlGbUnxf/4z3Xli+9wfcYo2
mogMLbqPUuLkeJMeNiGHQFkfg9fOe4/aAOFV6+pWs5npgqCX3bRnvSi0wMlcOmJI
xpDYdnvx409SBx7W43rZzWs4T1fACFpaiEGe4qUFAZJ4FFkV+nPc1XQIpvgJD4ym
U+fKF+rm+UwRfZDNfzO52mYEYDqnvW82xpd5X+eubUJTl8L4nECa56ueXBZ7pWWl
H7T2e0CktsHFB99HoKdpDgtbsXU60uItjjFVLWk41+8wxO9jr0XfnJ1VDluC4Mqg
gvktpq4vmevlnmaoHrH/MArEOCzhgMCt5iX+4hiLkMAEeftePjVdzRpnJ7JFO8sD
X/4nN/6HyqgL+3/bKA82VXAzyn65+L4IZULTY9qbo9bANmU7p3kfev+JnXWnW9OA
pu0yAf67/SX8385tg7/UserEtT+3qEN+RffIo809JrwZ0W8C4FT3xl1SXtR89R+H
`protect END_PROTECTED
