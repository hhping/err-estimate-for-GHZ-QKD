`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5pzaqs/fc8iwtHov/tE7JjqtsZrbAo2hx8uR5tYWn2B+UPekUZMsQay7ZyqM24NE
qF6yBaPOcPx4iG5ApOXSeD8csfHmcF62n/kSBvqaVESV510TEObkVrxsZARG2AsV
7+ueMoC8erR5LZVL3bEMNmLJ13gnbE9L9AuqEpfkQRqlAVl89lLflBCIVi4dEmAe
nQc4UFGBcsXqj/0ptODXvQ+ipzixoZWWC48xz1fBSaKFQDdyNKGRwYmBjDO1ozyG
rVo0sdbxh8Q2SE+SWHqinkLy+iUjkF8NdH2nWA0sALmfEhcxSCcVMY8wZpZoPxD7
xGbcGZgv0xPLwqX3XwmtGG0eDjFNbfcL9fNP97DyUgdDjF4gAxrLDpqfabDI5i43
amn8jXTXwgbfzYSG3upPRaLOp+CqDjcm9w72eHQ8rMEi00+bb0reakOLxY8Xdr0E
essBc0hpzj3w9qwJKp4D1kTnn9bDLg/DWvR/SHC2NujPK+Kbw0kgGOqIZ+BKVHCF
pHYzVlDCJ7dvFYq0wSzxWn+r/KLCyHHXiD0C2/1+euaOWkgT3R47loZhc9/R+95r
MBDbgZruSe2sIZab7a4vn5vRY9aFbdQGdb+pyCexf3lQRK5WqMHJIpl84mb47S7P
qOJm/6JfojWg+fNq/NPGRqJWomQReLwlLh0JLJMYvneO/K1bX1NwRLBNlGelYOy2
NU4mkKt+Jieugom5jxxjsbO2kSKD3Ptpd9i+/pkO8Xn3gnxX8xQFJYj0Wm+rz5f0
zfVP4+UJ0uFLc8ya+TCvu1csZnDJ6erGyCNNtMHmEwCVTXe59JFl4xPp3rHAGGpN
62vkxCcMSzEQrUtxcuQ8071NGBppXmRBkEHmXjz2k691SFDC7fIPJDBpTF9WbuTi
uB1lnRvzE4uPjr28/n5BaoTcwzSsNkJ7gC39yVdiEEThDqZkdK1M2pfpVKPMmrO3
vbZCEFaR3WtDOWc8BDWE8gibKM7PeIMQca4xWINN7QSVNjsg0B53NwDMpPTGrvXp
md8YKzm0ris+334c5c0M4I/rQIZbP+SZOPdwrHRXmA9WObMmT7SHZ59aAS2jo7Uo
oNPRlmp1y67TY0PjWxA6a9F1ALx1kvHXql6vayUBBv0ZND7p8+Fb7FsHoW3aYphh
l4u84aosXCrLimpedTam0sivHqQJ4KXOo2WiRgTI7mLIYCg1TfVdCAUqQ6JUodMJ
e8Zw6+VwooZyrJ8KXCSAN7J6Et5q2r/R0cpbH0uE6V3gQh2webdLrE4kdfpFcMYA
dIqLj3EyV7ZWcXHUIvd9UKCXWf9XYGivB6tB04VuY/UMHdOr8nUQRJ5SZ7b+XRzn
4+Vf5U5VmW6NRV9+94fKA5EFVe8nAyGLsoGlGeaRHxRShJo7qP33d4lQW30mFUsL
imWYbp/jRH1kCazSz1+JZ+oikx2KezLW9ygUP56ip1QAQ8AtZ/rlukL5Ti1uLBF5
QVT2ynMZYy8EQqa76WqcpQ==
`protect END_PROTECTED
