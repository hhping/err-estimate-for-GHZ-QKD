`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5sQmCmmfQf2YY5P6t5tZGcfrobTwikZwJ9STGuKbbP8EUMDUXeyqknqkci0JGxML
QnO4nKJ5c7t6NKBttp2NnIml6/vg260GAKuMcffLu1Tju11IlsHdgXTLDR9IWVbD
pwAhdR9wCWuHVxhV2JKvS/sbyGuIQKnI78GIp3HCJHG1+QC69cyjFb+/qQG7evAV
3OlFPzqQnrYwNw4RiRHiup9v8/JHA4hONnLSINcwgn3MGzFGYRq7zzMIsaWsXMIf
QiIjjL0TezVtQy1Z3NsZF+qHRSObnvvNuZkp3Am2GaStwoyvjlSY02d7F/XfIeg7
CjNkp7wMqr6E98kNoQr5aHVKx5djsJ+P+bk5IB7dSxTkWfhsaI8wnry+KE6pLGEN
Q+bC9ENxZBYrJ9sTiG9FduKHuD1g0aKLG7ZBdNPu7JpHRw/ZKfKT7qZxgHOxl3Qj
ieZtF0TPZocuW9YWCZrsOrC9/NZR1WYxtHVoIN1DYx7yAvttj7ne9p2O5cC8B4UT
LPnbMx7uoEDiRqcKVzhDnPMkTmE4qYS8CQJxfESHbl2lcS+9X8igPfI34yZ1DLy4
8Icq7ou5jiD7g7OR9q7CBbVB2Fa73p47fTCeO7yxIsGXnjIaF2yf+4b/mZ4aA7br
dAN/wM0WIj7RiEHc/oWT4qK/Oq2tVX8780EdsYLhN5/tV67hg7UHGsCeBAbO4lM9
+3Hp320ZwHCSlPepItwabg==
`protect END_PROTECTED
