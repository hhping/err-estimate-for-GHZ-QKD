`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SAzCwFFFbI4U4KjlPOacEoZWGBs1QR6P4zNTzgRKmi6nU238Tp4BJJft5E2Jyp+q
31eYpGVS8gJHU0e7IcjSUaX1iPOSha+xXbOqhXiA263+AIo84MUaqoyuDnbVA8oS
tjSOttsoZVF8WEcyTcxnnBrAP605t/mFPTG+lwfaSjmygkwEl41QSCPvKX/8msGt
/eaRNo0utTVt88pSRQ0d/HQdx+uUBh1p4fSQriN7uvjFYMecQSBtPQnXZfAbZ/4o
yy1aIO+8/Gaybtda2rCGBnGRbUm4gfF5FTUe+MX8uIBpAZEBj8msIbJbuVmNNYH3
REZGvRi4SzYESfRAlOkns7hmmxIkoCyUwx4yYMbp3I9WhX3EFfLtJAEOg4dLD22q
S/HJdWWc+STWYYftyCFx9F14UgglHfirlxwcqbjVWC0WS6BDdNzbHvB215FY40Wa
GxRbILoPAWO8BqfGsNavIMt7Xiq4AOjVgzkwn9E6ZpNot1A5FMqJMx8AoX3HMJ7b
NfQ9CKX8hoINIxYHjHhcffPJH+jvl5VCv2GLzKbHj5LNls+zNCKTgGRlcEPmAJ4i
hRODpZlq5/NXZfMj0V2R34KsT6PruD+dy9cKooL9wPCO+bC9psFAIGl/IrW0mQlk
SnR/cF3B6rgu4pmC1xH+J2l0wi4FcLqLOJccbkaY+/Gzus5eayKNSeM2lP0QTAtY
Ci+vBIHXz2KbzGuMwO6XGagEOWgMW4AEXRY2vE+rTDewGS0zHt/zxrkyby3+udPe
/JkSKcNLdWlVW6NKDSpN/N2ByvCUzqtlpOR8KR3KzZRDbTWbD2kUYEoU5R3vuWRc
/JZy1bfFbyOi6WzZwahOefOity9rgnpcbEIhdB6T/irhvLXM68hzUMhyRkBwnXg7
kOfDhfsu6+LoqlVsB7ALXaUSrWgAt1ocsbmn3fDX6HoJYDLH1SEXYOqRCRb8xa6s
WfV78Pr25bVbhaBeGHIeQG+RB+vXF9NpTTmlVBREl8j7aHElzwbPmbojpSQT32KY
x8WwwRGOpYyP6TmCJ0o2ZvClOCl7ztADUD3mIpBMhPH1Kgp265F7zp3neAH3OnM6
M/DxG/zvh57AO9/MV/qNOiRXB+vDuLrxc3pYMi1I7adW2zFhbZRKiw9emB6DKXp3
A1JAUM9miyxOGbdJdyGrCiOeXgx3WfClJdScIFOUnNV8nJ+AGyZLfEAw5hKr43Jq
dqUg7b/bDQSl43g1BWEu/3wd5m3IZsuuSH7lTn3H5dh3aJksPVz0kZfHc4zKCKez
i5Wsz1h0/NI2/MBujAIk9WUruA00Vxj7flxmxWO8RSX9hLSocTvURN4+Rh7xXh+W
cFFyu5OtwA0dxriAU8gtnKyJAnE499G/0G25YRgAKD5vP9bz2XzeLrA/u+9cP9s4
xhS4AEPbcsa6FV8kAa4mNpzTfQ1okJbkROuufUw/7pgOmf+uyjeDPBDDYLuPDuO3
KV0fGD/1ndCnGqQ+CgUbeeNjBSwMum6jF5ue5ewKbrrtyLW56ZSfkEa0aa5YbzrZ
lHoy8RtdQob6HSKgUIiDG8hbs4qErOgbKy+e2BiMfnx64y5xkerQo0z/JsoQO9W8
TahC+XsQq32DIJL/D5FZqoo0tgKfacP9VWgKPQakshPdDC7RhQSj4IZP9gB7KtEr
YULmhdX3Jf7e/iVzlmYrGJy/kC1BYe4BS1mEOSUS/Iae4QlRpSE8lgHz2Q/J7xMH
2boz6rU5z4DFvxa1gFw5j4byKmQ0lkI++tFDzSxMkq9wwZ8xRkLJVREl5h6I2EDO
IrahyU9oRadPKynlBtVGFrb62SQHJREi57tAN4reFZKuFtO0/6jAU9EhBwysBvl8
leydmhrZ7LtY/CUvUopp/KFJNTtFO150GZGirMW/t1Axn7xpttSdNh3Na8hYK+fH
0gcHkGUc45HeHu0Nv0L5BMXd2tnGapIU8EJpczE2wfhFYNec4cNxuyLENZh/rqh5
zxyZM5Zepg8khUBx0LMiIzXvznX35ndiRoOLWL2tDQWqUCil6VLXZDCpd482NKEr
JMoqI4gCZ4jk3WqVmrLJA3gJXKcYs+SsrVHuIF1eAWJQ8L8OQdHqY4YKAfAGaAxz
ZglVjg0kHvHrEnPAQknjxQ2wIJBk9jyaO0FIFTp4qC9iCW8qKICSiqokAz2TJ4zR
LItTUITUrqi0D9d+Jr118x8kPdFCj5TODfStVHXJpgOv/ed7ZI0H/NFKZM1lOqp+
e8j7DeKT6f2jEzRqmQZ7Z8i+ro6/zhMpLT4uGPrEj1UjnCjYH4m6Hh9YGmIMessS
XMAcKbPKf8ofxqppIOwP+HOaQQ5QmAafVtTy2oWSqgORJnFU97CK/guiRrFCRfAF
tip4iYSDK/Tl40D4jZjfIaovpM7MOC0IPH+qwbjUiHCwUQ08vXLkGUNwVblO/4EG
Eg+xA9KYg0SnI03BOd3L/k2ajgTREZFHA15G601xq0eWpw9Mi1+xKRDKH3i1bc5r
R53Xh4nAPJ7XvsphZSc0lcHram0fJD/D/1juCRnhhVXVmtLjmkc+/F2mXLGG05+E
mpbSWj1t4FOcqIwlYOsrSfLxDZlqlXORjqXb9BU2c8tJH0tD2gN3scXdzlD6rW4s
MdXhNSLJYSyx44Gv33zH9TJhb1FKT4K+frxH1BaSwCGRAqLoOAmp7uEJuvuspW4z
eI6HX/h/kjTwA1D6hAy2apooVoB7Dj18L007Tqr9nFoqyjCGACw5jGUtT1xc6iGL
xeAM4SvxFKS9hN3EwzQpFClgL6ZhdreLBw/ezy/EHwUvKd2g+1aQpN95/csEmM+e
WOCDWh/CSsYizzc6+GlL7yafkxjpc7EDWZckehGp/xi9hz2QFKkwCwjU3yO5Yvds
qN7NTXf5BiqEyRVKlpmf4+evuthYNsm0BC6Pfgqt1Omiy4ww/uTNW0omkQgy1oBD
yEJ//mkYWi9Dv8dWBQAKkbdhq2Nq3Q/QHhWa0VKPWIOyrOPEIL5bnJLXWVczllv4
nMhP5Sd67iNBkt7qux/wLakk1hUo9fejx0KSPhqV2QbNseq2XMDzaAjnOq2F7FrI
wErkRCkzh/rFS/CymGU5zzxBZst4zn5KEfMKLiNKXY2HvixqmHgVzxFGmgcNA3fO
R2Wqs84toCECywgoeaCMRh7ziyuSloUmKJWeonRupEew518gVrW9NcTT6FZ30Isc
+yklcMh9G2rYlmJw1m3zoo5LfY68d2CoAxtJ7DHomE4UNqTvDpl0U5aZIAQ1TJ8n
Y1tt74Hi7su1sIZIImSx3lHAAiCzq6a7G/9oQCt3ZNukqT9EAIV2Keh1GpYewFP8
uAa2mpdmWpg1eUITz3tsM8MCTOr4Kwuip9Nen2/VuHRQQVGjuellgVJ3OVKMCnAr
4nOjmDOIrTtO47quO7fr+Q3ZyapU7pFMmwAVi3oiVTKl8s7YLc46osOn/vRid0wO
OzKM3vFMy2e0rBXSZcufyzhggaGpaPaseUjiMWQrzJj6j6a3UYCVFBSa3F5+RUUX
44Jfx8drKdAckTmqW3XJzf06s91m6TO4nQUzcvUgCPAYuOzq20gq8bQXUeIAqCL4
3eIfVRVpawEY6jvXXN5mHw==
`protect END_PROTECTED
