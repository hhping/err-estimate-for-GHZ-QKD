`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wycEgckabGmH51h6velAi83GWzCuHjZFVmAv+mgPtlRK40U2gzUGef00CjL5EStA
CqpoCenG7mGCOAIeSF5oFjxwf5EtHDAD1YFDNIM8xsi0+zvEk8bmv8nkC/M/oqlt
pHBcZ2d8RQwvxP0ZQN+TMnn9IU9QcjSI1xiqAQLOORuPNz4tzWQ5BVUeiFrQlpcd
+plWkozofjg2la2iAE207nrwShspqgnejpkvWpj/JTueHl4Le79hNbAaHXR8kbnd
8Yo08ZUlkFA0kEXbgBejvF2jGYaJqOQ1c8b2+GCr9p4wH8zPW0tLnc0+Pkn/LHMc
9hn4/DYrY8bx4vXwRJKP7gVnnYZZ4xTimHQRll6y9cvkaSASQ7lCacOg7Nn38a4s
ZMay0czWB/oaP3sJVp3adzujZODXS9LDUoMz8ZqTDki+15qXX7Zmm56F2kn4QcLE
R5jsTLeuHzunOiR8/mvzUZWzT1kHlRMHBzDhzJywJxdG9cUtBv2Mi4PHXjTcDXO+
sKXVi5WGlefexfLBRNH4YCod++lKz++y5CKi0YQLwMMVA1OXrXjoohsqwlaK6cs1
vjXV8f0ITdi7pT6807Z/4u9auo6co8ooEvN2jDJanli3Ul0DSwZNdUX5jCP6Aaja
Is5hZjX776T9jbTORpyWUNGFsbS2Kz9tgmGLJ3lt1FqpruLz4P8qClJFPtQx6ZPk
zWEHVV4M6evXz4VNjqtA4uR35r+Uj2h1yvPk826PFpLDWGRe4GfVEmOT4Iap7TUa
UZMUy8k7PAvATKVqbPEVBeObabsJAbqq9rLZZQ7DlI3yNInps+pCVGRel9UpqbKG
gyRbiBL0SFpZAOhWq/awqTW6mb+833UL2N/bRSh2Ytb8rtj2u0gaOO/ldS1auV8F
775F88hII6+DLxtLlvR0/zuV+nPFdrIoEjRpKZQFfVbdzRMuAPBVSGcklcz4Cv1D
M3rs7pfqYlTFITF5GtOuKdQSvNP1eyXKNwX14XxHQxWg7jRzleYtzFYWaAHfEgDJ
lljx9dB0MhMGESnnxFTW2bic9R8TR/mhZ21N13pJ0YbjQdrTyFnq5ch31nEuTfx8
CuWY7BhGeQrC+dyU2uM7MPEO2aVJHsNxyC64h/jcn27p5ccROxrZ88FcK6v/Toh8
JPLBJUU+K3tdITzYfEoTcva+2F4usE2O/frV/AwQ5rtl8Z+EiCss46un1vVwb2p4
UXiTRvRvuSzsblscypCTjBanFh/gSYfaemp82KBDeddAFTFiQRmrnGqSxLhy7ajV
l4NHvIYVYy6UkQNkfK4BoFfjqH+VWvgZBgN32bzSCC5vdShaGJpUR5n0qVQMc3CW
1FJozgaIPr4kXyLD78sejcerOU/KrxrX/zjtlhm91Zkft0tCztMxM9leXvidEjHB
07n+JQjSD0txEWNRIR3IIZyJL19ldJVO/OzUse+LWd9EjT3cryIUOvI8JqEsZJSc
H9f8L47C52g+o5xvWiSp/wLhxtV8uvbyhtzGfmOzUwbc3P9UJT7lsDIMLqnTr0pY
P1h0ck1riwvEJ7oPtBSr67UsvQQcy9JncNxfZ+I2TwEoftEeIfK/ej04XzsgMxeF
z/uvNQaCo+t6dYVqFBsb8vlCQ19J02ADwMP+2xAg1REs8j0dLvtajC+CDMk2bPsV
MvY+0aZO7gFJldz/Qv3JhqZRspGFhjqM6C6FD7Tq3xtZwzqwMAIDM0qJcRZi8rum
hGX+Wz0hzRZ2Mv4c/47ytEUKsFuM0h47tl8pcfAMspgJu5dggixFTohrRXRa1e7v
oC24WP4ra06CsmgXHnTTPqkEa6hbPvxunzjBfwRfuYF/JzvBFDTMh2Ug07Xo719k
5RvVlsqP3a5rBH7BWbr1hfadUfbuHBXuSKNFa/S0CNYdDnHAkn7ptYQ3Tvdk4cY6
E0kK4b5DD9PhGYm05AKiSBIgpNo10qLL0dEyXbHDa+70Jdrq4KCW5gCCZ/aoiud6
LHTThLuWHryYX+Xn23rkZPnrd2uO4GDm821596DH9iwkHZj+U29lsHdo2R1Ed1p3
xpqBgtoPiQMPaVUHXN05M8L+hZ0baNN2+EtRfEzZ3yLCAlLzinM52cN1/noNJ6TN
sQlpwdKZygQ9Q71jj+Z6fNt8/wjqMyBnSE+Tks6C0mGJjHoNMudTzBhKpk8dT3v7
zc2MifzezSIObwniP/WoxvMw0XNWrLUzrsZD8KtcXckhUm1MCqy4fgEvyKmNHsZ4
sGr6q1r1GEuavscSKWPzsgDzmSYzGXHzodHzDUCjFIEalmPiUs+JxyTDrzdgwxWg
bhXyV0PvsXVakpQWPs8SnmdrYnfrrVOcBk+Ou6vlbkruRnODFHqMIeO0jYq81K6T
6x/YkizR09m9wiHGv8DTl+2L38m6gMusFB9ZM/F4ghsf6rZxIVaIoV4MFtwqZLUd
1C5Sn18V4/1HNNlNcoS+8t6e67mZUfo1KxJuAM9CiooKWklmGBDl3I+375aGbYDW
3F/+hpvXF0C1hWTNanhWEkKCp5sF1a7BJJoMRzVsISrlUkvLHO7N4BHZ+xQ10Wad
DreA38gwyep1nphVctkOqYOsgozyMLtsqSm1RgYwd/QnKrJxRF1nx6f1X6kRK3L8
cZOGTJtZ478wpNgEvJGfTW0MInMZ1g4ht6Ln/k2X5OwaLq/Y3YDlZ3JyVSAwz12k
13un1X97SsBe7dfoX7Wr9VVS4V0hH9P5O1NAK49/Mj3BKfriahB9MVC8tav3+J07
WWNVr79tv/WsDmLd7gjRyBOhA/Rwu/VnHquCnBkvWiaJrppkGB3VwvW17iBmaWtF
7Msx4gIAONuI34XuGJ4WYWcMvh+MA6UCwypUW5nMJjlAw5oBswzhDVqygEcJ5bCA
a84VCKDbZo81F25Wp5ePEtDKZle85SkSzYlcC1TCXdxc5djsYybsnguAucGtH9Gs
wI2X9mxc8GSvvgNqONvIOTaxGwoAEAgf8uTzsjhaEgDWq1APL/gWWVAVr1A4RiY6
NFVDK/9AasbDvZEe+sGfUIn1s65Nw2WET7P0r6TKuCjtbbY1WttzhvkXWmu11LuL
+kHEPtby8ENSIxI/47bWymiTYnk6tLZd2XEQN2zqHP5WLmJMiaziWIpOrIRHfuX+
/T5rkfVRZT9wBmgCE8O06rsgE3tLFMEd1wRQZcuAqD7iiDK3BxSpXVCFKPxeOR16
nzWJtz1W2Cy34J7Hc6gUAYLaBfpN2d3SMKWOur2Bbp+fuBvT9FZ/uFvCFmp1sh0z
5+g0NqBW12uPDGQDuG0d9dc3y4L6SaydhYt2pSisS1s9e7MnYe/r7jykEZGunfoB
m8Ci1hD/liblm4p3ChRQbYzY+LSuq+mKqDpRH2PD1xlqamkqvjTNOXmdgruoXFgW
OyoDd6IwN3i6Rl6PQFbWNYyzfo4TnfAyVZ8TtH7SQStt6UUGvhUsi1uNXVpJPOz+
wTwWRmlD5Hk1maR3pZUeEZTBwxcAP+wx39rPqX/QhRJwdfRXNDJQ0fi+7c5IhIp1
WlX/JvJvPgKahcIH45jJEsMZPpBP5osZ/BJYoM/rF6Fbb9Rj2bTGOmyV++4u2XEb
ob0soAiynxP9IRdaAvsabiq1aoKDTi69xeHe78XmunCGFIwa67mLkgahLaVa1YSU
VnXc9dzN6++zF0EFuDN+8SdluAOVjkuVC+aF3Kza/TDrYzy77183OFHmjhmj3Awd
b4IeOElzWMHnOZsQv78t2pFT0oa2FVij5ony48IsD3V/flMSyii5JJolWAQwrvu0
17QB6jeH/7fWEgWbmVdChnve6MdSPxUM0psz0kF0F+QjGx/sqCqkvUjGH4PVIyUl
mYmFRX0onODmU4RZkNKTnBp/aZs7xadF7OVwqydnIuBIoJrYN98SavpLsZqZCwtp
9PI4uGo8/gEXOvtSI/y9FBlpPlz82LRrtjwFR2FHeBEkCW0jlWe4CgWoVKVv+Is6
tritztem4EgwVHfGx+LRghvWKmXozLHoIgtq50irDtQVMA41lXrzG8WjGk2Ng3bu
265iXDbcestvh8GiBYH4FcyZpBG2qajjAk/tPAnUC3mgi14iRXRkkglTfnESlBNW
WCUmcbVPPAj/u/160QQFKdBwbmaQq9kzphW0HZc0/pdURULxQcw9WiNYQQEUQ//k
NsxcxXoKG1gJa1Pkyar4HXsPIZZOPJ3AVGpMQ2XpJ06Qv6Z2BofA+K7Kcicbyft9
UDxgDgusHMm1EQ6YSWZhkaKmrJVzNC2v/IxalTVc0zjuYVypYlPZ2as2PtFrVwU8
ZoD+w7eQx5ti+8J5cy1tQnVOagXWfI4xWIDCGX0hUHa5i6Cv7xWjdd2ukmOGolEl
R1T+Pu9IGSAzJF8LRp5caMlYLcpGQ40ap6jPBBuwhKo=
`protect END_PROTECTED
