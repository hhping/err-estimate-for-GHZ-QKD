`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+DYe8i6hkTFHl9Qpoia9LlAr+3Jvg7dUxOKMOIQln7+6Wyr9QLUzOcFA4N58dghh
LQ4FFguebkv2f7VgYcLgLojbQu+a/Xm2pTjK7zqH3OuU/lAPxRhNwGKE71Zv1tQ0
RyXWXcCLT9KZboSk23i+GB0j1RpDKW7Khuctfgj/pMuGUzFr/x2fVCZMmPhejppo
j5rrsrNVJFbIREAoBTTjK3YPjQuhYeS1ght+t1gBNGPwMSwlqAnXgkiLnGCElBry
9TRvZWRWpZbfenGLY+QZibGfrsxKCJU+w5dUW/6MR91h9MZqNYCJTveOgL1glgyI
4/ToJgjV3Bc/VudfhEKrO33HpYBUozWzgRSb4kAAv2RV9BbXyYT/nbdMF25uzWEf
59FGAARugWB1WJQgAfoGAH/5zQx9INTnoG8Yh0BJk/h0QZrnNV2jXLscOBPDAuLb
pW0RS28KcsFRI7f47AwCkmxndDgqnj8IzdKYCLRf3c60t4+FUmId8YcSDLWBrYj9
3GiqwqVza9u7BZlJyQF/of+DDNLs1LE7NaMynljoLxEDRw4BmXXn6g15kpk1LSxk
ag3w1HoNDFcsCIKELEafNqtPb3repodR2PxkagnbViF9595124GTXp/mY6ODGiJE
W8wq2zoNKBAno8dIMvx52VPn8uR5wG6tyD4OHKSl81i7AXpMqKUnhCdMRMAOxyVc
aNcgFpWXktzC0kSlMW0wXxWOdFlXGOVqqnRoYywMStLbJoZ3SWcR006R4gidGLNO
jpxUJ5B+nqSJ0gVXyzzpdtra4nd415FvxxVnxGbPneI6Ge11hT3LUryw2aFkrhVS
4xb0QF/V50TDQu6jt8L93HF+VJmP4xpN3DcoMsq5kPfLCIlABsHTtv37m57tDId5
Q0hcQpDzbVnfpuy5F378PMJEE/WkGsgd4cktHzqsqYEtmb3GV1e7dGGu5HxMUeMA
ZDEgb27eNqgJw2kOhqPhJrRKM4OpOYfMYNrSyLqBJ3H27OCv6chlAJ/6DekFDtzC
//Qly621qRUQvteTrRm5hwqxuZuV35moLJE5vc0g7NlSsLq6rtMUKE5GF++osTe8
dL0UsVec0F+vKIV03rgu3gn3NjxBQ5Tia0YiWSdcWx3pfO0Si8pFlrt+G5qnG6rD
tonVRrVwy8CxZUi5oOnkEnanwUDmh6ImlIdP/TENhITchYXBMA0RbuLAPaFn7zc3
f+b3cBi+s96+tL93Db7riFYyWoSfqFoGx4515V3+DSMNZTC/ybAeq7E/Nm91Pc4X
BBB16Rr+dF3ws1IUha4Ikgr/6E2TisVxmDpEPXzv6RTEw3XpXjOhHUHBgK+rJHUQ
Ol3U7uG6aobYI03/gv0bmvvXn1ndSm5+w0bRXN4xCeg/Iv8UqT/8EB0kgNJW8rtl
epIqVX78JPqvDT511WJLpEk+BWKroyFXMq1Knw5iWEQ0jJPyNugGmPLRcCGZtebc
zsxpXWlFgbGO7Be1cVW9Am0bZmegE2mkGR9PmCZG2+R5Rb4zUm88arJ7wTt60fKy
veBlNBmTQwZE2TGlPw8DqLRlvYmtlTzEuuKMou0IhOxNIJzNRCho0y2/FaT/jkdo
0cviIhbHbsML17YMzHfFtLvvRC9wyTLgI8zAFr++8pIxNEJsDmq042BInSRawgP/
QlwORFQjgDF+b4Y5OxGN9/c82vN0uG3L73UySmfegLZFzgpSpsn9uGXYyEQ4YE4b
k6u88esNdSx3Si84F0w6qfsk1or9qaJzMdu6Hr0hPHCqWwSbZ7K9AQhPJI2IJURd
UEw6kSxlzZjwwi7Fu38Lho5ThGmwyPCFBKXXovlhTjPJVX96POzREcMwUrSaLIKm
G/eosmqaHNud23hxpl9cWpO0GmxaB5avVpLiej8Au4nLmqeBvP2fJ+F+MWuLXuE7
ManbRE28fy50CD1vTCcTR9UZ7ArTwyWjlAqPH5HeJzIslsm7LM8x2vOkbzZsRd4F
NZLYTAghX2RMNVkeh9PT54t7vK7hHnAhVfE1iecepA3aMRh84LvB4myFnek0nD80
/c+aDWq4MSZ9JavtKzWUEx3pRbZfrTakIOhEFeUmJhn1dbXTpMXtrC2ZH9XYlHXL
zw8FvlXgTQ/1hjCgnt1S2P/uorTQp0yhb72UMTo+Tsz3FiRKnAih5gohjAr04wxj
e6Ru5678zGtlYJ86+2Hz4nAkGG0ICEtgPt0pPmcnmJBPWwHr9Np6Aah96T0ouyQJ
hO0ZmLvVrCZtSvKq3sCCgNj05DBVNuDQILgiBjjbRiAuUxOhw8ADcPttDEMbfeis
l9sWhA1vafR4HWorw2uODkmLxdTXw+KI97YbBJwWY0Jfia0kuybs29FQ8IiBqL4c
uP+A6ZkMPmqs9D3okzwYy15zIVTKM6K4hVGnX0vWyoaXJzW8JYbzS0wiuh78PB0e
TtoPJWn0u2PP7UVqm0EqzJYyT8YLsGHoGtNq6wL7MHY/yASv6QzrhTYJpxkfYkxt
gYwPh0H1YGk90/SxPzXnOQ==
`protect END_PROTECTED
