`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/AMYlamjRspkJKW2DYvc8BztpkUezwdQyx+UvPi9IZ/oMh7jy58wDRj7ocsQHOkJ
ASeME3vucodaKHc0TVljsBWSi3drORwDW7JupvsqHAv/On2DSOg/TBBp/pGbZ95A
0c9J8D5kcfRP62JnBVfKOiggTik+p33lNYy3eO03dejof+dC9EaiVG6CUsGv3NZo
Dd7waCBYtpyheaMN9+vzjdOVQSo9a6Gn4M4B7r5k112RIIXnK9j3GZpVxmz3pvpo
YuGcZA3OCEz0ZRQuEe5IaFKVQwqoAIrQGmWY6hkyT0ao8hcGiUcGVBuY3R1SPkb8
jqYdpUSphKBL3FnMuz5mM5FE28wSnvNg0g/gQJZIWnNIrUHn7fFU6VCurgRJBs1b
+55e7/5tEUzVM/5BYtgsajqxLnimxbPNSTfxohPpc31ak0csgjoaso3WvHUY99Zq
KyygBRdg3e1j7s27WZ/OsXFBvR63tAiNfZzuTnXBauuJLoUXP2PEp0xoz/r2HqRp
OX+Nt8M158ZnM1mQ0JKq01mm5ID89V+6VgZhk4xg/ZbswJUhgQKv1BGBa3A4Rq/W
9pLG0fkmnNeW8GSTfgyno8hHaFO/lyznDnkob5Gk8DtKDp3GzHadq6PvQ1TIDT7m
hxZFW2mGFMhQJzN7kG3N0DKZmCLhqhE9y6COJgkpe8697vk+RVcEUQWgQFSscyzu
TX4Wjib8EFG58YccFD6jdsHmcAElFcZoIiDoRmilE5zTWdfvulgEqKEmcuSxFCP+
mfs2NMj7PrEkUEtrQsRlomNKd1T8mbWqB5wOSpN9dDU=
`protect END_PROTECTED
