`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ipTuhneBD08vT0Zdnf/V0yvYtBP6Wk0lRv+Wu2p3u05jaWYW+ECQGoQxrOkbmj1Y
hUBsluuSh/h0/N65mTqnIL7zqfZtzOhj6L6cbbAuGzO6VneAKW4v4muS8Ce1Y6Zf
Hl/Pb1shhRviYSZzdMWwxAR3eYv15Ayz/NMOgixflMPBJGBxRnvnrjBeQzwie79S
Z4ETBiUs1LR1S3LHTWGP2jf2wts01eRERcTdlxmAREn2y6dV896Ky+WmYx6xIB2P
IttFothO1acKOkE0oLzwoqIq1sHGoGABygEQKmQ7Ja2h2dMHi0cGzsLTzQUF3pjH
Sq50KzfztUYvVYUZS58BUIbpODHdf7eFdB9u14KVSEj4Ne7TCEw+DLl8vaYpizav
D6hrUVmevflR3MnXckSnCVUhbrgHjFM+V70AgriIdqjgFI/v/pT7RLjYTyr4jQnm
7alYDkvHLFML56MoP3EDX8sc4GQjohfm+k3xKSUzAm1vBbE3ajbXZoWighlE5pVY
mO2sVNS4+dMSLvxHjKh8wu55P/ZrkIjD/uyGzCpNHTf84Mgqz3O+OgSAzslxgsYh
MkBvuWAaB16VOnnkzqMNztD+LLaSTVLkrLOIJtStAZJ3frkTCDXs00tezUfZ4aYD
Ivr5EA0avU95Mk5bV0W+HTq273G73eYgsop3GBgOzjWmneWQPS//E4kkZCdw+N/I
syjQpAOjyUedoSeeNqFuqVRGr5ftYHC4JnTpgOXqGg8xCCXTaqccrQJZXgzohHX5
gR7B+G7CHKGA7v4VPeevVcx/BSTKwkQlynx+krjVdoQHz5vLJP0rNiA1PVZmJT4p
3gIZaLwoERBWtZIM4lDD3xmZ3K9nTuL3LClqa2puQtNRu5UhGLXDWZUiFSvS7iAw
liqBdhnrlBkO4jbNLLxGbwXtHxifyzX7Bi7e7CZrHAdOkN4zg+sY3ttapVXfyrwy
MQcQZPQiOBW0xNGzDMfQmyGU7EtJ3RjxdKgaWfKq4wpMu/2yPGekAMsvT2N/z8MP
SkrO8r2NCnRWGhx2PozV3gLt7cLBvjJQjZjfbjurLHOx7ofVt9XQ131IinDV/yq2
wfvlbTW+ZgIaj3mwXpCc8AvlJ7DP79VVKrXItvSaJGs9fWt0sZZUzALty6cKEJfs
fTO7qhgvXYKFusuvmmdTZ8DeVQaoxfBQ7obdDgpEQBnbEQy1kL5l8zig3kggaOkC
yJ8EXrXKdnlz5gTrs9xAHV1cE2zkPe0+2pG4Pdj+N1ypDES/dVItfl3DcwXDDvTV
UsJ8djWGpZd4QiPV11MZmekJBffB5r99wKwhlomgPp+fIJhL4J9+2x7cAXNvDukO
njY9FiMeXChNsrmvZ5ZBh8NXvtYGu9d9vvSE4Cc45azxtEt+V+kzFf6q3qqhFp2V
tE+va3m56sUIJWMZ7vvl0vvv64j82vtTved23jdZuMfqGv9c0K5eI41sMVLJ0nwx
Kle+8B/iC7IvTlY7VMd4Wxoz/MuRBfVOEyp8djGJqi449vGwWcmsfmmjZna1P+Vq
o+jaCtTlb5IVgiH3hs+mZyUH6pUdnvhQXD7GvzQNWu0fuz8Xhfy66tuTPZculoNT
ipWzciMXWhSniTyjv1ZJ1xG78badQMibCcOUEsohqx1jMi/GZqEhHrWw14+HWjjv
+Kd8ePlGISAHPerN2SThWqKWHbwqXbMZfxp4NJ0RkWP5SN2fixGevq1z4IbuYNVP
nJasYaWTUiJoz8nsRKtqiWKfX+QPNjeUtwJ9i4WYOM2yAlsPPyp8hHUDzRQc5aPw
cXH2vMMWHVxfuUSMctv/8tXTFp9vh7cDFdpEIGLA6wAYhL1+UB5R0VR4WdcvZXtz
plJZIZtWjQCNoV1PfPwNc8WRpbxvOHASXYGcrQ8X1gz2FUShMipI8Obf3kDxulf/
OAHaE5oiPk806vUQQtxNllbfAsK+fqinHzaZnFxD8KyVNJ71+RfZMTwiYP98CZZL
mDXobORF00N1/T0sXd5+lwq4anrU996Qez1vIvGjbGoKdsrf2hdeOlgC1cVeEjsB
PxJIMydZHMlyqD1rr4bfadjhgau3Bq6Ld1mbQdFbt28lo5jVpkjK9KxdxparOccZ
FOp+n3E9vHeO7EINrZUm+a7rDR+YstyQ78mYNz2a9N73LnX6T8SS2GR+1QeV8ZPd
+SkuMJzyTojRL9sJ2/XKsrKl+tt1ISEXBdjxdU/uGoO99V3oPRu+Saom6imPXBJO
qRuIhIyQNo+0vLKT2mtJpjod1xHiQN4kxul/Q99j0YfyLhRPVhQrGt9+XonZs9xU
185PrujYzd37ZttsvCfJDGyM6zvTqe2dZedeH6mnUJhKKbDoQTV5/Rs66QWUtBYP
6BeeQPI9EvN4KPcnonOU9/5ZWvexjqeqt38UYNwM7zeQRycnvvUwx6BPnJ0kXggv
lx0J99dbhYaNrp+7r3WC19dgzplQWJRJQymosaOFzN54KQiQ5ozbezde4bseCakZ
GB4BoiqkUtYTjK0V6yBLa5RrGD+hXAf9KC8PNKGJBtw1M54CUqHkFY7JWFHJuivu
2ZWZoBftH1dUOc8rI/ofZBCvPuI7yiFgHVXKiHu4S6Cf24ES/CPHPw5McC5blmH1
rsdqd1WDH7PRP2seHl01y+HYedRG+W3Fu48dSS1O7ZW71RKpqlk1qwwQu/IrOIQ+
VeUurWQDbj65Gx9CUtwV3LCoFA92Hz4Vnd9TCPpqhmbcpvmbxQs4NhlmjW4Xp9XG
3FsEQhc1uwk3ZCko/fijeAPl++76wvoEGEwHiSoL8zgb02DFyV7jd9aTiOvRJPkE
wiajtWZeuwUdfGFry42GRGvUzMU9fd2jZJRz4pv/j3diN8UonGaFEpqqvxLVfxN2
R8lUTvdhKvSDd7UZynBeKJi49gAQM13Ywh1npv0TkEygBWRhwEVJIvTEZeLP3K3u
Hq1GAbIKcKdNGRZ2GkBKZByUnmasEUEkrMGrb+/pGO4ceSx9aA8frDELiXhpUr3w
geUEuj7K2VsJ7XJH/H0Rk5pD6s67T3Q9qta0R+Aj1qA1chSL28BebisR+IC10Gm4
AExm3JnZPDwa3Nn09pHNKQgs/Fg/efwTbQNm+SZQlgrQxMnnpKQuEmbaYD+P2KYE
RiyeGx1Es+cfmX40sRiBaESiiArWIkhmPZs9E1y40zC7dXQOmNVTeDC7Gh6wz4Oc
lBIBITkLeDtIZaK5kF/kQ3TgzAejPGw3MXTF7WzuXWT5olbNBY8zoNJjinxH+JYQ
lcO98nhSNbnFkuIqaMbK/HHQTmArNSpQ8b0RvEq94yxcygeP7bWgDhCFrWZ5reb+
EMqvpmw6te4oIgwc2bDeaWJdeCNEs78mhVQcMjlZCmEloTKao6gif19/MgwW8sN6
BfZfQVxxLXdUGI9fVciOMvdfml+9MNhUWsBPGK+7TOPzeUrAu1GJrO5SLpnn4Oax
X4kQs0aESPoN1xKffWKzEPHSukrkpnu2JhR4spNOnzd0lSMIbMFvfpknR7fYo5kD
jXxvMO/4Z+E9+6bSmn0uDGoSgetLXCQaPr0cPJ1/rHQ=
`protect END_PROTECTED
