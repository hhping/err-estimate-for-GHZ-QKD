`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dWq6OFDF5NDtvu5fHjPa8GygICvteUzVAQXt9AhhMfGUGP9Iri/xFsjWtiBsrNHG
ekDhE8eW1htyOYYN34aO/bCzgwJ4kr0LHaQ8qwnk+ttICK+gzEi7XvJfqQiRMzne
GayT+d/ycEoAp5JYo5Fp0S14CjnaBhmyo0sjs27IkoLgywK5l7ERYxU87vHnsHol
DrFEAfPNrza1sXv4oZ5vQCqsv0gdFg6NknbJjUYqJjEDlWwO3r0RwahPHMMT3kk5
lzEaQ0qUeYsBjPLRDtjB3sV7JiEvqvtAoJRNlRHnt5woISnZNC0ht0dB1MhKq3Eh
gC3fKcuvHbAFuW833O+GFVlQ1+MpJHUw+aOagylAlZQgWW/neEp9HinbCORFlG4T
DElRNUEGD6mnLLCRxleDB0haiVsX0zRuwhQq1FTEu+ZitBsv38MygUjQL6NMzpFe
UZ5fryYW1TUNX432qwX+hfyUIWiLmG/zUGZdWwE8CYOv+eD/tqFb0XmtPqsNJccs
ADzvZnZrw0vmpTKHsvcWvoHGn1FkIrs4J7HFoJqy7a1A3OjdRx4yaHmzM9+frp2O
qW70+76sDalpRHaMuNEDOPlxebkuzbwKLnt/B6AX+Gd3mga1uSDG+XR8GePNHVXF
a3JD+N6jj4rdBOHamjSf50gtu0dkBi/EyoQGeyfncoJx09gtk3pCtr5xBXcVZATx
meJTY2KHtJ8DUm76t28DarQELEr00gbMYNRSpbqr9eETf8V7TFE9+d2QGZj8qczW
r31MJLsh2Lq6gSGT0zZP7ZFzoryomtB80UkfyX7fk5mLHiCBSC8J+8wkvbGMon+t
OKYEUzFoD8Zrh1wFW/8cGaYRMqqk5gncN6I0FLTjGxp+lxYk1gXiJCq5GGJdL+vk
pru84itcXVR3OWuyRMXYJgwidSByM5Rug6Jjsv77qDZXFzUDD+5z3oE2/9H8oODc
oce2ROXVD+8GDODtbofMsyzmtQh1g6fgKhYdEO/lQzdl4upX0BZqpKqYude8UWZk
wZBJeByTcxjTv4sRzIhf5mU66So6ZzNbVAqgEXaTmq1QUN/hDWj2VIlzpuZ/VJGS
gVAZssI8YGRPERFtRUWkG/OOtc4GOMc+Eiy15dNCsF+BmNrTcFiaviTt2bTGpC8q
RPdsukpo9+cDh56LbH0kBhijpECl9QKnkaxRB88Nqizu8SPJXxG053h/CneazrrL
O0Pa4U2ZIEBdQOYEkLIuzlYUOW3sM7LuSFcpS8U1b6VtlZi0uuqn1CNU5SR/zXIV
d2/HZfVhEjHNnu8GAvB7Uj3YqthdZmXoDHZiH30NHac3Hqiy2vsie1Td8+x41yIy
XY/rH84yPCSuJcNgRZzB1RsD7xRMAA0UKE8u3bjKb6GVQOaOSs62SiqQTe5FtUpd
hT5mReSz2jc431qN7GvTJWceo1Kc6XegXgNBclpf105FtS5KW8r7MDigHOXZStnL
2AVKUf6tk39/g9ZQyjdWe3ZOmK/tePQEm+XtqsEQcV9Zgu1HQCtTJmsh4d+S8kpr
uy+Yf9S3rxprfc9QdjmJ43gYHLFUVatZ9CaWzHYmv/wthz9vSSuybrYclQbR1TfW
EL4vDXrl57eCHOXxAxLi3GeJKcYa9vHj4MAheabALRmw1ltYyLXpL2BUl0u3w9i7
x1mtKfGLaUPFTuVKtAH8tUBV48zGl5Jp9KP3i+N6aVtVCKzYiTiahys8kv/kUukh
CbmnS4rwQTTl0BHx0g6ChBAK2V2Luq6ML1/U516ZCCFWPtutjXeuprWNBfMbADf/
y8q+47DTSUwkebkfMJT8Qgi+eRDWOx+bd5avgvRYmtqyr5yGWtDu1qHsbvjEDfaK
KOU4JOtqkz1W/MR9PzzxKB/u627ppsZnwn8G5AuIBGpQgdvm1+dOCfl+C8MJN1Yj
UlrzECCaLe+b/faEPj8kfcTb8GfVYrgdvqc+lbhqUdFCcY+XT5pLFsSM3VsachGC
1jYcXILYnIEY0apAzPeyTq+c2laWXz0PBLu3CQiAOmzFxJxJ+i4AibeYtKtM3aXI
yz82HY8CL39k96loc9QTTFguuxBhV+IorGdn4pBCNfMpOeK9dQeLSgyUBCLzdter
vtpf+9HlgLP1jXKX7YrhkpQFDDIh08mygN6rLl87Y4+Vl2ZHur5Ckj7Hx2nDK7ql
Ed+MtpaSmV/uH43E8PbRSOupE1GZF59aRKwwrSVekUWLdl9UbLRLed1iUHkssVur
WajnlyeDJIxWSeR63oaDgLP78V0+SspLvpB+YKVxqup+d0ys4/twczAUYhLBaBOK
eCw1uF2XZ08VdA85kS60PHa0DW02fG32KcRLmNdafyklc0IDRfxekwr8yE7ZfjQN
WmDsNJDKs2zdrmBHoAmvRzthuUnXkiFis47miwx1K6JBPD6n6wheaeHkIU7Iwb45
8lXTjSwLGT1PmBNIEf9Uo2CmvzkxpSpb34w0KPTyLaEH5s3Ns3/Uiu+0MJKRVAzr
39mpKQhiak8hqB6xH4xuXi+sh309hyg5Gz5UN0xEip0RsgnBwWuqGQDrM//a8WBo
/tbZzllLF9KbZ0IZTv2bTOwYglUXtRBeSH7eD8or15gc0J4axoLTKfGD7YF/EqPA
yXXoksg6z9HpOs3gMe+DNv3rpG2+C977zI3fsOgtCIRaT/wDnKq5bWXF6fPtsest
t/soeNmRKrVGJKD1asebnUi7dimhzIL1mhb+sQHiF10vq0JZl+BMsJXYPfLEBOTH
OTgfStJx/RICUkcmi3nhr6qS+IuDPXWfzuQXorkBKRhhyVSONS4wos6aDut8g5D8
8rVPd0orLIB52DoyQ5K9u0j0+x8UTnf9xY2rqppGUPUqXXW41o3zD0r6kESedRqh
cB5VbSPlsA9XnQoZIGx7DoxPYcGxl9ujpo+BSzN+CwTKQ2nw215YE63KId/m8pMu
s5xewPSZfr0CY7zKvEDR5gfyFJNprumQP9f6ml98G7OMlqXgCYh93mHSWt4kUs9d
to6mv2e1nLOm4ZImVlAGj6Mch2oSktgcpI26pbq7DaQ8iNDEdkHumwfXIDxhx4ef
1ccordnXDCmnzKOPrgPBIqQxwgUXwUHbELWs86u+GST+A0CGVz5kV6eFAym87K1w
t5aymwdQXta26Cy/8kS1iH4MpZXvT+RmM/L2/HgdbDBXOPNyUKLGzt7TV85l86bI
iOOhnGo5u7IR3OC088YR+qVxBmHk4mJuaGctFfw8PrKTyTLcWBl0fOEz+SuJl6nW
p3fElMljuHoy+ZiFqDRnoybKdyMnvV4kgrZ7szLkPgknEuBgR31MYv7T4/xa27Sk
jcrClEkJLg9bKJZz5SbCo/dRJvosA9eE+cKW5kLfGuio6wS8c8ntkRP9SnRWDcS4
nduY271gZ5Qa8KcDfmzHWF6y6IqOJrOktJ34k1B/19EMrXnvHtW1+b7qDH15QwXX
FmrOP978jpcnbD8ItY1q6sAp4sKxOpcPTvx1z6tI8H8QSvwvgR8qjAf9xPj9r+aL
LZf7YK/262W1bzi2IiXCQOp/fnhXxbRIz3Mng70W4ejNsuBlzFC1IiKie1IiNyfo
A0FKK+VdWch++GV485nJCFWkvn+lZ5IWHp1+jzPuLRU0SOpqlFs/eqJwmT8ydiEs
uMIzpys+H2Ijf2PFbQ+LjKnvxFI13q63jxRHTpqoZrq0FjoeZZUb0fbK3D7NFgOW
VtznK/qu4nsT18KyssunX0eQUS+RsnLLFk4E3OZQ4AxydxzapC3MXIuCwjiaDnI+
qgLYxQ4kfYY9K8XjuhKBnurhFjMxu2yfWDVYXIrjfMXHMYYjxjZeOpa2gjUlLYXM
3BWgUdCq045H3y28MLtZodGg+bPStEg8xoaGN6PMCRqZYd8DkfQS5pgxe+ox5zlL
nT4bbuToWeQCIwGRtVyuQ2yHTqEnsUbuCeirDhmC509HcBbJ1gD4tKVF0xkQhUpA
Mcgq2ileqmmC2u4cIyNb+amttHDRnMRFVeZ0L1t2w/rhhczI0qY1MUcodn3pzMwv
PndFg6q4TH0m0e8GpWirwKz5t4U90sipjj+h4VWTVPloa4sidJrz1cUHfP9TUIqj
XAS97ff8va6bocDzeLaFeHgyCceSW8e/Ps3bm3G0BzeZ1DAiqnVhmbge+mR/T1Zv
keprGAEhX/qL35iCZpk5ohuxO2ihpT+RNKsrpMX+SofH2tDi5Ih2yG5mG2gfW4oL
1UAmj8wBm0ZY41J8EZ0V5XeHP/a1aePsSaDnvaKjBmism7JwqKV3kaepALwZd2LX
/JJihlH2H/Vd/oDxZc1xSc4n82VD67HdtgmHA1pa1FjmZZNk7+/aB1MccKXD+HXz
VV0vukwARxyJyxxncvSX2FXvNX2f+VXTFGH09bmPxWgpHUkBq0fp9VqYnPlPBs8N
uxJY1QOqb9a6f3aHPeIDGTQttbRwb+JdjRB+taEUCUdSaelZ/NPqDr8XIcFd0AGh
uEARvHH0IvHdFMezoaBkGI4V/90NCkIFrLMBQPTsMmaEZBtDn2R6fEAB+nDOF7Wz
cNXxWjJOap6xt2jU5FNERElRpt6Frnz/Ybs0flmjek09MQHB8ywwtNKgK1YEqJE6
FXrQFsC3Xzt7Z9h7l9gqSIwmxiralyxg3bi0lDVpX+PA4IATLzWfZfto4m/odurt
0/ZGK0mQntBt75vpH1NmCscl6TXZdTTh6QEAenkC/OMQ7MLIKBaoDvWZATcuGp6w
kGFhRZxrvoCdtAVemW2umtN/HkZ8MgR/ZELmobPdsb2Rtf3M4w0O/s1zZAL66Tln
eHkh7w5A+Xi+VMeyjtQs8ONiRaKqjnAGFaDf3a3Z7B5H8nYWOlJhgM56E8eriQwb
W1FljrbmLyQBCKemty5iL8DJfKSStrez+D6z+2e0rr6ASCE4BxpL3PdoDKAN+hTH
2iu/l4jnCavTsxtlThSd9eoLvnW8yJjUWMexz5g1554qeDcmNTVvzR/u7SlmsuJy
aw51qmInmQz1rpX6cpI+Qzl2yyb7ibOWx7aJI4TGmA04vM8VUchKmwyE5r4iXL++
SA0MvR01Ac5Zj7weeJluD57RqQfdo4jQ5I6QqiAw1kAxEV1q4v+dDYqi86ADqTBu
IMYZ3Q3zqZP8Yv64r5bzL6EFczg3TFD71DaFCXKuu2dya5AIbTxXWmPqj1En26qt
zVWj9Bl6/F1EA5P1CCHb3fwFovLjTRaUVIAmtn0FuZnv5Xqwndk6bJmTVBs6JdIY
rP2yled7zXX1BCT15RN8ptEhosRvU0p8FAv0KmZuRchlVHSjtgovng3/Rf+NWLRA
4904Z1goJ+ExzUa6hqvmgAiHogcpBGOI5HQgtwyF6/Po1MHikEotM5q7G6xrly8u
xzEvxJeLMuYEWPCgFyxcYxkBFWYcTvN2pb8giF3exzPkh/FCHYsuAd4eap4YvOiy
Os72ro/39hRb/nU0UkE2mbQnSSn3ITFpLJYGpUko4dTjWLJaCrjAHzuzIZRfx4bo
OTw57ThyRP7lSV00YAYmDNwfwbMVqwh03l9EIL7RTSqJ5vVcHJ07XY0dSG+qiNve
M6KKY9r/1TlKjRMd4uJNutw98Iu02F04BqRuYUfYawjZcT51Aw5tMwaGCDhjCMQL
NerTOI5oqiofvU99jf+kBxn5ETRJkPz+mfQL4t3Zg+M6m96oiEOytEAwblTYnqQo
xnSBxJvqyZpO8ige2p7+HRJRbfN2w1GTBkiYX95K4cijIkFZwFosdbA6NiX6UeuH
Kh5ygNPh0kTUmAXOhZB6UhbfKvezSxyfQPJASYm9ixxqg1hk+LkZdUfI8HUGh93+
PAZJdh6/owrjOWdEtElx9k8aOhUCbUPHkZsGL7bwUDnap/UGd0lEwVMZ6EL6r4hE
p9EhtDiRXz7Bm98FABu71iRGWsRH6Rv4jT38pB4rMDE1Pz+nLk3xPZ74lfDYe8xn
n0LOBSBm6M6DEfP0xdMD+zFhSOP/nDWf6iuiap1g6cDP96D+oocO1H0O5Aqr3SmL
200gbnEFKShzhekTRQ4kH6VyvSfvVdtIn9CX806ZyByU35PB//68/BEvRaqzuYYP
RCJ7/LNS15sd+i0bN+t5STTRCfJjXlseRpI+qy4o23WCAZ8kEusTtEs5VpfqhenT
LkB+8nt79kwD9ZBs0DxwlQF758A+qaeEaJ/pBw9ZcKuVF8FhLKZtoOG29P6ARWVu
QlxQ/KMNFVGnDN9Wn7i7WLXNblroipNC4AQ7pAQw0lwc4l6XBru76z7D+KvxHMvL
Hl01B6as+9rWdSHWXppYVD6JZHpTUuW6ERSZNGhXk0Opsxxr72QPcNWfUlhU09Pa
wn6QTAUBjyOGOLW82XAfjT8B4QVGaKk3ebvf/2Sc4wn+ZSmk9PzMyTgI/cKCMh/4
ZO+d77p9Fhj+OUXfs8zvrtetsABqbXF2NdhiPQ3hVHvDYwoZeRgcDf+J5LRy0/vM
+9d88bOhhz6IdXbD+lueg67QPZrPPNuG9y24wfVruqcmTMXVFlBhocJIrL7WUif1
OBfEK04ENjoMOaCBa9SzwbzEvOdQsWnmFrWDRFQaW/MZAEqpW1jIRci8/k8rnn+O
Q57ztRGGnrfzPNCwoWUgOl1laPCuFTxn9U+Ecacj1Z2GuGQNaqHMBOEuD8xADvoA
ovLiw7eWbAVJMshAxGxhDDN4PBU8WQUlOYYLCVWtS5FaDM3tfFhvo0OSITKOJ+Bq
UYhMXpZFGSe2ljKUVaX7LDuU8vmk9/4gsl7ACLzwyKw63JHgQAGtIKJEMQO/psVP
/m95SVHTJSpIFLd4TbZzK0fZDqwREl8S0x2fXWHf3YtlzRbKjI81neWXhpdhQGBP
MJa6rP+JqguH29LIEpS/FLZo7V9uH1D7e96ytlrasDom/ZLD2bYdbvE3NUxo11+E
VdUntgnCSEMRe2iOx6OdUNuFZAVY0Jc6Xkimz3qeVwqAq5Qhh54WKikwWexR3Lcy
HbBNZVUENiZJjhEfflKPvkb667G1fsBIkZC1iNnvNQQzyCgcVQeIzc9Z7agNwnHG
M2MYVmoghc91kbKVkG/MFX8A34tYCgDBYHmlZQTCzagyeCTMTyOFWyhcLwPWfBT9
ZMnfU0cEh8+KZ2GID21QrJBSu/Pxe9T8ogP9tAFJeDTdb8qU75YEZC+TgdQEVMeb
7/41G9/bqQK4ZkO0RyrfmAkydnB3pXfdkQvaAN35o8zHra+ycTDBr/euboxJ8xUA
uRWzM170UpTi6MbIBCCCSZJRJz838i5JPFITD4uVKNDBRcTkTm0J0BVABcOxUxSH
HPvqNJUTtP4Y90WP/n/70Xc3OvikbMhPu0JHzLQ/JV/fMckIYeUgRbPU0b4qoaQE
RaVXLF8JMHwYQFAIXgvcrBvTc2wAGkArWvKubNh1BAQq/J/2n97vC5k0rbjCmYL4
tuD8FPObHwN5YxgnAzFOXDGKL4gDP6bRftO96HVe3NcWBUVFz3Va8s9FSzcf0WfK
uwaOYKWKepipbym+G5FvTPMb3+FAYHlprwhuPjFgQ76jrtP8NkgzmKUOWRsH1lKE
rmMIFGePmKxAEb/2BQwgJURhsjl+SGDsK4ZQ0/rkKCs8On+TTg5SeCnZ1qMubMjF
1pNg7B4JFSA5a4vp43DTXsCrpbo1pzRkMRjhlUAdFbbhiJedVj0v7CnU5SOLrIuF
8L0jCoTkt6iW5P4Xj0eMe8REd30ywD5pNHUDcEkHPWXi2KqnsoehC0IcaSPwm9Te
LB8T0CJSnEQOzHiExSVUClIoI3OzXK3CkSFGxToan8/lslioIfGQ6YsCEIsWrHR/
F9vvanH9MpyGLC/N0Fs4Pz53p/ks9kY3EEKSQhdRoIJHp4rNXQ1NNEIISDKFAhNp
o+6X24aUPK7w86ggxpoAD64VN6bJZoPotsJ4gU437n1UFwMsRYsvNjr77J2e33dS
3hzGHTZ+oBBv6pg/IvENhvchnTwyqeYAOIsHr7SEk2gVEjmf5th3ttfLzrY3aX4u
LqmtNc6Rr/aiHm5JvjsXi9qCRQhLaB6QxChT92uXtvqd8SnExvfBMXSJrKvGFCtW
5mCwrcaUGPi4+OpACmC2x1OAos/5idYjuBZpBFnFPBia4iQEWR6ARaw9lEGQcU+Z
4ts7PhAONeWhGfh74NFD/c8KKPWZSfaD1ZmA2MlAydBHckUyS6vxFJjw2G3MY2Sw
mNuyjym59jQQ5rc1erFJB8zJoOnPXJfMxmJ7dXMfArFciwnl05l/YYLPrGO8rWEF
VDiGZM7rJ5UmQMGIM2DArS/BbEPehWTW1jaf0DLk7Hu3LWm6CYuXurysaF/JHREM
VE8Hcgb3PRKEWj3YphWR5jLcRiZcnx+SC1d6prKVIgOT1X8j27ZMv3XyW5ilrvOh
tOqaoA8Z0U82eTFq7aOibsTy5WXkL9GhHjPxauIEdlWnWW+GZITsKvOVMBSnSZlL
DORD6LJEBIbPKQkQu6G37kqa6ILDQ1J+N/Caefw1QMzkmBsQwaGKI0k928UfSc5H
farR/Hq8vp1+5ZSrr3ny5F8gONss/8+Tk5AVLD73/U9yXTWfBUuQiSIHFgVe9oOj
o6JznCvO4BwCLL8vxQcFTH3wwvNl7vD/Uguv4XQ7OxtgrCjbbhao+vksAOgmo57y
exRk3DoIumbmpsaZ8tKv9YJkO3gQJgpvSFrZU/40grA=
`protect END_PROTECTED
