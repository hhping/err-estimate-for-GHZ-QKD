`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/VJ6aBl14qV97g8TC4nAzTFDBltIs0sw3kod62x1JJxoN9siOCxFiTiBKz3sQJUv
y6a9RlS88sZyaSca8lVVSy2HnLb9FIRXHPtlj601q7lbg2pbVbgJK+1VloSFfWle
tnA/0E/eTSCJ+zriAxqLFOHZGQQfZLQ/R3mgB67ExifebedS/olz+hSx5nI265Zx
RncUdGooE681gGMhqYQBavlzMPq6cNUzSnrsfQz01N+3P7ZSZOogpAMw7mcxESKU
hWF1knq+NzPdeNabpQjMrwizMtalvSh3EcztE0ss/dvwDqQZNvAWqlDASJjSXeeR
CCnXos/+DIIeLS8llmKzYRbkT6aOYN46U2N/jzcRreFC5Bl7m4Erx89kz3enPOai
8RBKHl4B0QeR+1qA7csUmM8roazzYSa8KpWxereKs+1+gjRVViDpkQuG6e6YVYSo
ARtTf6eNzha5Y9kvlytWEL+JpyjokzNwSHDnpAS0HPcRfXb1AqOkGzz+GuEBXoJ3
XaYUdj74vN+z/qCUBTbGooco1KrAwzbkC7WrpxJyd7FVZAZMGYJ3BmpPpNv9Rfxv
2xz+8IujgOXD4KkoMQ7h61T02aTmdG4YLiz+CWn1o1+2I5DM8UqfPm0TTix78xkF
9RnX65mJQHUbtT4XSGGO0Q==
`protect END_PROTECTED
