`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WWsHFwv+8zkS9Y23q7R4sAYGxZJsnJqa0MbEEsvjkzM803N6n8Kznw9EiamyDNPg
srMYkwv8a1s8hB5Z/YNNnzKOJevvIVOhe/X1EME4US4mrFa/0puCoi1S9g278chw
ZYm7ml2egb18OapA5rRn5UWSAZfReoEo4VQokPgHbUqpFqIaCTE4id9lnukOIsjq
LBSJ7MyhVrzGtPnSemNoA1Bmvak4VjM5501WIzkEVZ6vsqDIy7vf3M2cIQzTMzAD
QMnSAEFQNZpdJL9+4X7e0z/z3exxX6kxebkp7fj3Njvlq12XmjFOZzP/JPA1aCdq
OzfjvyhbInx2HaFCFmRaDoZ+fS3BPZgBb3CmsDZUwQMse4s3veYFqzynKrh5v2yz
3TKeVybLWie3KDMfCmLEVN8YF6F8L85GDyL4eR7jU1GYZqmXaMh9pgC8HmDwkz18
9Li83mK29jOe6UyWty/PYRsYzZ4sbA05PMjdTChDh+W0ifnC9yykQOEGJeonwK82
BCrD8zjyl7VQt/RqTSUulSt8eDdMhCgKSRNPTdDdJ7vyenIzt9ESpi+cGPki0AAA
/ftqmC7aN4K5bOt3YI/rHGeuAxKbAdpYFxsUhrCCt/pnWhdOWS1KgZtYSv2i9INP
NZ1AWaBh1xJWPj5a0BC0xwpRoe/bZNdX1hHAce2jpWcchVhQt4VLU1qrLaNCOe/3
iPt60HOSBdQmlsNT73mOZLaCAf3Gqr235BWXsB1Inh/MpWeXjmrKRGBPgwjip2ZE
A9WUdayxzIJtrql2i5r55Agq0AZObe1MvTRPMYxTSBfCJzQZ5k1SXUrjIbO4yRWg
gs4pxvBhtiNnwwfOtQzq+MsWQcTT43iWHabCHUGkxUooylOJcoNFILW25VafRVYW
UzFc8WNZ6A1lXAIshR+lzh0A+yrjt1m3dxyl2RCBBx1i6pqKLQDyN+LQz2sTxOZO
HSSrO2cV6rjezlBrjyortN0Po/0EuZS3Yxl8XahhoID9x68hP0uM21GfRH2P08iM
zkbEXNXjO0JE9Ph/Q9zRql/v8ifYLVNefckrOk3vlq0AEqP1REQMpxhFHlCHRkfq
Mf+vnnLRdZvug/5rMaeKRAxAc2ZtcsveaPDCoZ8R5MDQ/nNCcX+wQaJL8k6MWX2y
IcM9E0Kf7gTmT/l5I/SBeC4OZuqrFhgAEyQMPwcsYh85B7YabqB0eQKLiAuLqSca
Uj/x9RrEFtNOTi5LGjAkhoZ8ii34VIq63VDkPg6fYWCDPCPUpkvDxUSCdIwBOZ7W
zeblSg8YJl5d+ZwTmls69Zj6nMp2L4KZwTGzohoWD2Z8uBr5P1hBpTYIMAp6YZik
kMo+7PPW1MIXB/g5gurANQva4m5sMm+XIt7W2guiXB8GSjr18au4NDBgJk9TDmnR
LbwIqxd2+VdczdLQj+PKojR39dRQ0H6PNKqYgy9fjpr0T+ux/KV062Nmc/0LDh1F
kqFqStJ1R8JOkZtGmHKb2RJSFlIQFN1gi4jaKqHeG191AXwUtxLrVTjZRu4sA732
S32qkaBu2iZspcBL5TpKALzApQi4ILw/o/p+Q4ijs5CnpxIt5NOSR8wDgRL0yXhZ
l+WLsQrLuDJQ3MyEtTnyOBpPiqqeOVjk1RSq7YRrMZVOej+3JrwKhb3vwZ7th5yg
8Ne/lG06yuAirk5YanH7kGc2gqubwQAK6N+OsBjMJbaElbBhS2cOlasF1ntcNnI7
37x4fxl9X8pyKwo5g8A2cQ==
`protect END_PROTECTED
