`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/LUmLxObnmwL37GzoZ4fJ56VkuncGBngFrzxRLrobPIPRwRgs41p9w/NPr4y9ZpT
VEx7idYJYZ8wAxWj9MdgvhDdcy6MHVb+HjpUdKugK53gIUFPc3t5/QG6LFTW6vZ+
VXySg7sBHSQEjdKwVBRFoRWUC1pCbGWZ0tCeaZYklDdDyIRv+v/V6vsOcXcEyGjy
jW3mir63x8eT8ifGRduK+Pbq/oZFoCnocm7/m/RJ6mO67twxxb3d0dRY70l6dKNY
sPJadZF09SsINNmkigCtJR6SISbUBXD/UQ0jHmlVxMqyQSBnKymWKUNXIVq5VG69
9Sqlm3KdlJyokmGscuenUuAZaS+tL6SM/qL46IPxBskLGjlt9yPhioCiUqHGJDzD
cIuRJoL0k4MXccu4IXiAkrNmZdMsjgJuXquvlYJ4ZV2rGRp0E1rY3o1c0cCLQQ2l
xzIVxuS0gI94johvHyOODHS0FwA5NtpcwVdqbsXMe8GC03JxttEgD4TvGcw78woB
aBYaUJP0JfWSPS/tIjVwo/NTzXFBis04/GGHQouOWtjL2DPRkXuviJ3X03FMqkyd
PMV1b7YXplunNEpxMgjYLYChqb7lynsqsTGEpY5ldCGxsFfgQ99YlALqKQe96bxu
X6XdqR9rGXEpBTExDoFVL0VhspmUrPpYj10MFVBezZRIFFooqqcrRBxS6cIxwf+q
oP+406n0dBZvWXJ7qTPKgVU23NuMsEoTlaZjTs32pnkoCnbnDT+B2ybGTIIX1YNX
QKGqu39RHbdVcOT1iL1XRkaTz90UZNhlcnLybvyeWCI+6azOg5LFUmMBfnjgLD76
ilEsZiFk0sTpc4uiYe29livNEeyo5l2ciWpjYVwupSQFoNj+v084KR+3SrXeES/G
TMwRURgVlmDtiRI96OLwQvxO+SUatjKJp4tNR6GtWtRbxbPpPPIXYgHjUzr4GG6p
66Tk4f+A7puiwwPiYGM8w3BvmVw46GwCueqjv8QGeo2dD79R+9xLIpnenwJXqwvB
m8vKMEK8mhwRe5sX6jd6X05MdEoPYTuq0X3Lr7eXUjM=
`protect END_PROTECTED
