`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nLj2YvnK2ydG0NmS+FO+4PIPkM1IoqJRfhbhYNymiShwbv9A4Aa7Ui498yoq5DaS
UkiCMnFl6HD3j3khL+gAZIvNKf1c8e4p7f76O4P3o3xsRWeT87iNSqQvJ15M6EKa
JZS6ySyx1DQpnGt035DU6/Te9nMwCQb446WandP2CBnClrbUTIFcE1QfyAyBd1As
6NXQWNCW6YdQUKCLcsLXBmYoJB9uYJ281co3hSP7Uk4HmeLWK2c3XIvqgutMclEb
VM8rOHkTKnN0fofeEJmsFvWzNZm1tjvZ1WUDCSyuIuRovWG8SQUJHHlRn/+pD7xJ
5zgzkScqTMy4Xj5T2CWD0ww6kmHx8cAHdZqWVM6K6XNiRviIrfPIeekNIAcq8Vk5
5+jBYW+fzA3GPINbIJynYEsOLSUqBQfdo+Vp7PmsX9GxUthDVuwgR3NWxI3QmJPN
5VxJzjlOkPzbst+05zuOlSfLhV3o7hsworTK1XXskVg/IyhEfwd4B4nF16G+ejQ+
ddTL6nevlLYoGDsro5O258nvLk9K8QDBn6oV8w0CkoFab2Sd+dSai1iyfh8hNoy8
l46r7J96S5SsTne+syJcwo0LzZVw19zLr14bnQLL5EmIeXU+xafcB/Rzrj8dcwQJ
cnIwq05APt94Lek94kdt2wf25IW9NX1e58Mzuo3TqUz2vfr9RWfXrgqGiTZSrXSm
dX7HR3u1fqalVpTt3rwgvliNsZmL2vOEBvPOhiPQ4dY66gYYTruQu1gC7XMxovjo
e99PE6g3H02mJfnzp17vjB1qBluPrc3u8lXmCPlXNmRVovW7hnCOuUnU8Ll6FUIq
YmeXpTQBOGvqEai0kyV5HVpu148eTCkqyfBtZBIUHweJKVGyoakb/8GICn6JsKRr
sz8aa9zqXi8u2HiVAi+JV55PhBpAVYaDShbuYzNFe4U+tDhDGxYVTRQ1Xy2Wc58z
4O8HqA2XSl61qz/aAIEDh6y1jpDRibSRd+CUlX9SwegmbOsk5me6vE7f/Ru2BrEN
Ad1Hq2nF22645grMyg56wveHNaaWnRZgYkPQWlkdsKc7LmSm+T7lZPaGGm03fT0C
rcWiiPOUhwMwASvG/jcT/d+Wm3QNPw3zJt15D3dPat6Nx6kNtL30TkEWGHEoGVfI
L3SJqmGXtQUtvZuiyRE0Fo2hEqfjrauYafOi78qOaGk2mWjCwcDAsg4lIi1H28Np
3KvQHdSaF1k/O6IfQhW2ExoZnlueQ6owgUj8u7qkTjzMxGdKnTaF4d886mWU/py1
ysQG+2Ykd7EHJxZgvIVZp20CfEVKCqKTfA/PGaTgRHA=
`protect END_PROTECTED
