`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sd09uyQMzkAlGJ1N11csYwqzQtEN/NXRYY4NiFj78UB3/SxgJ815nyDz0BzslY0j
aZ6XRfSlzpsWkIi9GpCCUNZ/VR3Y8KeiNouX93dQ34IagipBdzhOwlLkJ/ddkXd5
fB3/C1TulpmroQlIJqk+ae9AW6Bo1cXTsmOj2vTKOex4/7msgiOXEMqJg6rOI9BA
JfWJ8y3OYD0cscIkkZ9QnH4zSiMRX5YTO+w8EftpRtK1gkfdnr2oXrogVsxvhiMY
xTvffsmvShl0kJ1u+M5gFNRJEqctATPqlL+FFmbywTcVTWCJZ4pvixE6S1D6yMop
ZGm5nZFfefScSxatOUPPCYQV2ZtM6vn76XGbldu+POGFEn9wD5cuwM4YS16gV5Uc
IXgecyXb81GILprFhkzW1GVkdgm6JQNF3g4qFBgHZyeDXmiFYsxjYOggHnDCdf5g
dq8EFyjUYyis5JK58sRkqNZ5/m6QTskSzPmogAjdVph1dstUN2Ny5u7cr1FZqNcR
msk6oJqCWO+MmsUQkCRYxAbrKDJhnAQxDZ+yIpnie4qdmrk9fKsvaV522zLSSMQE
BU0MEl5GKrSssPVGEGJbJp3bZBr9XtX+cLBzQHY1NJ1CKB8zO3HOx3ehHaIj52Hq
ELDEnFyLhj/vLaFqapaDpcy6ARwTSzf8uMlWeQbqHWDOdrSEDobET5gmsUxicboV
+kkjxEClN97vQQVdDxkAYrf75ocAkhxFqnRqwByqV7byxlQROt0/J8RBJhIui/Td
`protect END_PROTECTED
