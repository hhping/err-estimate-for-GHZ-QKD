`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L41nDk9zPPG4ZG+4d+gxqPY1xAtKW5np6TRxprYgtz2SJGvvaCl/85qaDBXSYLjt
5L8Xf6I3XwZQi1xsWVcmhSZY0Fhi0EMN8fknJUu7qMHVBBrqV0tx7GBlxSWmmwJ9
sEJX1Vtr+0zbj1zbDV7SY9p+q075NrVR9qaO0jZoADPdhQP/Oo3/ovGQXwpzyqSc
nzQSnBYX96XgUncTSNRwlvTcVGcV23oHQr4WrZSPG3NTdLC+TYDJVpVzUbrDn5nl
M0DDeVwDa1J6yxfapeGC0MbTK0PVUoubtWK44mW+Zg2/+ygZRonFN3s6gL8uhMAD
At3SaZZFw1c24YIifz/9V4/Gy1Gi/OGNT7Lq0hC5q216+q5YfrD3zepijpDFkArU
36oKuSnFE6pNZ7s7/mhf3ZTqowdMiydbHE7jzPkPB1cYe+90SZFbI+3/7c0hxesh
YyfTnPB3NN8a8AyQTiabqIL2KQ65BibUWotWh1pW+yJzHkKatFQhM43VsGBMoZ9Z
LMU+X5gaAxUAhHsMR8AfXS4HYwWZZc4Rtve2fv5/4ymzUHI78+Oqj8SZjOnzmecr
ftfXIfhAxdWkSD5k90W5GJjpQ+R/d6O+tXLdcZiWFTu4KJdMoBgs8tF+086RCxc+
efKIMPU+cv3sONNyN+Vx2uuvPT78xm/lKfjKDDeHUAjx2QSkp8i41T8S38POXVbd
rwLIxaCA3vjL8VugAVFpm8jJ73NPACdjSiK1wZbG6mRdToWO3KhfbPMx/0UyE0fa
A7yVXX6Yln6+dX3+ZGzDPQ==
`protect END_PROTECTED
