`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TxH8LlcwKAk2522nisT6g2jzGKsVn5bIMaZ8e3FtaRyc8i8pn4uZJjRp3K9tLCPc
ukZgowelfPn/fDTZm1uYrEfeRIF0Vmw3uNzMGIPKV4CnjTYds4K1CG7jPILDj+KQ
rOIB4R1+yzgNDhGo9mAUwucKR46b0A9tFyWbvGOXYqN9Lz2dXpWnXhZNLhZFaJTH
pUIk0nDKYnDrmOrY4PLmD1iWK5U+NLJ4TaV6+dOA7aEYxIlEkinD8Ni/iMsDO+Et
CR+eswiWnzW4F9I2P+VJU9w3X8FW7ebp3sIawXVK9b0zdl2LrlvJwRQKlzNWLRDE
DcyPjg/INJKYE0rp79Ki9PwzMg2ZPGw0lkrAiY7NYYX2RvP/x+oZmnZBSzYkGCFT
dvCr/di4kkQXuFriNEF9Lf1QpVItvqgl9t7pxfSRH3frD11w56ZOXC05T8KDIIX5
zMNlY1+4ItoTrYuDBI6rHzuCUNQD2Yozl6vnOfd9N0KYO46yWey5y7vqL1qEb5Ir
AJXDuyQMmZg9kdYPXumb8JeqQ18QCOcIz/qjwbO0/Dtp2vEHhXwwCHREKkkehX5w
yLDJy4aavuSDU6BHzhi0n5Chtrh+xuJFM8Z789hp0BooCaHaoCJbtzqGJn8OaHKb
vk9rDJlYhvnauqXcWKh2H3uU4ds0PmMnr68qRmPNWNCzxyOKs3aaM+8hGs9zYG0w
x6FLCmT7KIzmeMfOjBwqYE7JlAgRwrvcLsmMoY/hAVcd31PiLhQHRtDTFYb8uiMc
5wJRGeZfItjytpxh02gZL36sOX1FAqz9C5yWPny6fL49a6hd9LxYkULEWU80am7j
QpJU/cicJBo3+5GFtYdvVC99N3bjrINRM03+LTDoUdE7Uwc3FGtl5tPuYNvG51Zf
RrIxdZJjzuHNMDqyvMIaqGwprfkszhu1aQIAxJsEmwbQ7sADAIkWjrn3Qo+Myjq6
eURA9il0mbTGy3kDogjbqBzRccwTbJ+Xjdk8xCqV8ipYy2PlkGHA4qUKd4pmWl8b
Av1bwU5sF5lRRcbk2DmgjhAbAhUmzKyMVLXEHcx+hZYos/eNus+6MBcwsO4Ebgg+
Ec8e8Yq3nbvD1ki9VAEFoimicqMFlpmQViSol6y3eBhxgmChPSpKxywK+M5Qx3OP
44SGgrZ5aHDownvxLY5c9xsmBJ9/Jhiax4kUwvjT387RUg6xan1AR1v/3ztCUkxK
CS5/j83QnUY7CnSr5VvnMBiyfGRP7DdtHJbVJaeLhPwT9bQASJPFj1qBn3RLYVHn
xvVm7E/AZEWRxw2cLjFr7IcE+nxIsaRfSkH7dtzO38k=
`protect END_PROTECTED
