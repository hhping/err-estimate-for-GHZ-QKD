`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J18rIT1rVw5BEEHFCXAvZnGnyo+wdsSsboW6jmuKX862dLwMDF4kXHLBeQqGbwcH
vsm2wlSeAixUhnsJ9JfB2n4MTWadwSbGVbadmoPuQSHpv2eFkso7xyWa4NWNrsCz
2V4dA/R3GmhCAaRuots7GH65dSOCPjtoA8Bd2bCkQv1DTVi0MEnIfGKeMJJ4B92R
ZlFuwSVP0zuLv49dGwVoSQCP1/Haf57f7imRpRXfURt/QmSC0DxFk/jEGv/7RnFE
1bxHFSd5Ve4aokmWn61sdGCPp1izX8dAud+32+0cw/YkAXY8Z0fq93XmJ+5hlyik
Uk8OqAFfUQCURaS7qfqwlfkgkZjMTZr0abxiycRoA92fsKrsP1adJH2e4noKPhRW
iKY3OLiW8+eh/1/UmVCOaP7IP2epJvCkViPv/7Kd7v6EKRlXj0mV73129XqlxcZB
wniDkBLxC15peHHR8lGjUVz+01dkb38p/UCT8fyI6OR87h2yWSpyuBooXLd6JbHd
`protect END_PROTECTED
