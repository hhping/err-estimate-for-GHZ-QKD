`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D7tUjCRSwWr35BM4wgTQo71A1bXKtx4fHMpPHoCkmJ1D6dcX0iHG3qnERTy0sX9S
9NwKijtJ2aBCcLISPqx4jLAfK13Qxhiubs0do51jRSWlDzLNwmUjBtc5V9s3efp3
x3/TGgLwjUpTAmCEu7Hi8P9OOC6orQNUoxWisJS1qN2qEc+PhWsbRMObaKMZakVI
h3OhO4AV5Sz39rkDXScyPKgjAtQ6pGGmGYEFt8wvFMP91Mddag8N7ehRGCEZanSZ
szTi5EAbujLncZZ1RDKGoDdhcigeF7aWQg/4NayDNwG7YNY+lLLaPYQkTPSy2kpu
FZNXT4jXoVXjnjSu+WT49OM3sV1EuAdaLA5sVhNArw+2xBk+zul6HJmvd0nvMSg7
YaeiEUvxiFvTOtpSE9TTb+1uXgCTDRdencMIHaNx/MeX1tC8pQhmglF7/R9Iivc4
JrSzzLk0jvuMCOlclpEjkTbDn4OzQXnF33cAkmHDWEEw6baUriXMkOpQIlkomSTP
x0xWbhJZQ3tRNaIF2T0E/lbq2amHN7tKsV6wPSSEJrvgU2Rxbt1iQ8nonqLgZ+rB
GqNRg9WCwPSqfysAHfpEXEBOlqDbQs1MjUa/1TW5J9ii1iNN5tIhgs3mqKHw5UqT
je43zsQa7ND/FPDIhz6idMAFzoGW04EVl/1QcHB4BFZs4QYkxy1zVtT5lCGx7MuS
EQwK2kL+MsWSRtrUiRj21xVykkaXNJ0hnBHeVz4lg4XhIQA9But5Po4Lmdj5oj2s
8dgeixBwOUpcN9c1IHA3ak7hPMvO1cqrx9zNWrW5LS+3M8ubjWrhWqDjf4EYHGCg
V0tp406V2DkjquKUvs6mz0W5D/pYWtr4Kj63kSlpzttz487wJ1/jgeH93B783SV+
aiyt9askW06TVkwkC8/m+eDV3QIlz55D/CESuxS/rXtpVUcW9Ouu+zk2FYyazlwX
h5s9c42RYWgM6fs3XVeVvEFsDHRSwq+fTdJf/+Ps+Au6EZSpH3b2rSgLCb1wCtm6
blLIedno5egyFJDqcOHtISdOxBdZ39Z0d4ZOwFRnv4oGbvWdrXFdIeb3lhAyb6vH
P/78SAgBwjG6c8NMvQvm3+JJda1xf/vfZfmfRnAEjXe2jbu0/TxbUtd5Tv+Ho/jz
8jMeFpH8Ry51mj4S++gKhriGIcuyLNSBbfXaNI8kcuS1X1sln+khZU35R+rOhUUF
/04+EEmojW30eV30Ay5tgRlK5joN8ovScSMCGSEB/YUk2Cl2xeMoGw6XTvuiX3Xo
fYz/uWm7aWGtSLgYaN7a3Nt6+BefeTOTl+auxAFeTmdE75cO4TW7r0VNP9zCnP9/
uIvE0OJzrhqyiYYvV1QsAhdbY4uvyKNYVrKrIt1pP0Ned/y9/AYcCJZBW/c5PYko
0o6QlaSjOX7WmfnDjXfAzeSSW3Exem54Ywqp4WCLn52dpo5prVy+LE8PmMcQv06+
`protect END_PROTECTED
