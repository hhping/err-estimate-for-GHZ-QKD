`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tQX6hxQRg+Do7LQgsymwjzPb6xUuKUmFdRJbFLry/laENQr1wUbkxv432Ph0EpiF
0CDw0f2v3o2PwWW+/LH/1PuEMllZ3T9xx6qLI06erGeynqlzJ1LAiWjpFpP0AcGJ
JQI2TEl1EeaiYq3E8dwPu3nyGci2AYzIxGrb7MLuosAO6S+eUxqy0ZkCug6WERfl
9qt1YKkMQQ3Z1bhgt030EkC1xNpNtnyNooUuv/ca2I96WpdfLokWdN8q/Q9agRao
7gKxbJbDpHvdObKGPpBh8Py6tpuHstq5V6KyT69GlqJC3AYQzkdeDwHISuc1M6Pc
T/Sifwy3/omri56im5GLO23WPVW/PXjZ+Q1l0W68SXuG3wabXNUMRFWMyEz48twD
WOhWlL30FKYJ6RjpM0JLZZCts2WyJnlijav+j3KsVEHkhq9Qx8cMVcg72NzIqhW8
JwxjogbPoBqgWBQ8o/DbI8qQu3/2mA/W9Kp9BJOpikMAZLVBqa8Qo6HNtSxGbadX
bS0xgjizmkb+TQJSYbMsqMOFrtm8cowidXoq/5xzyyc2g+CR4FJmrNrRVzEQ8E+V
LSYQDudbwetBjcGeQvtZifCXYmtyf+becoyez3pihDu4gLgZamPia3eamvLTuUAx
bzCzIC+M6JqhB/scRjS26od6TuRmQKafkfQAWlgn0MNSAK9aW3nIjSR8uj0kFQns
euILVVBQw6R3hogWFIUO53kbwAv3YUceKWwP7rU0I0r1Pb8LY04yn2DkKwj5M/Uu
2FQGlvOH5/c05mrKofDO0GGL/42GRNlFprbq+BS89cSbT9hpjvK9D5uZBGVQ8cXA
vtR0gc+TR7fMKHbECgs+BhMARHxpBiFAD7lRzPm7fG9tXmFArrkqwofliWRa7pn2
meNbgMZkMdRj9rpTWYvlqHnGhMNmqPa/IkDGssT0LtQ=
`protect END_PROTECTED
