`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BK5+qyuFHWRZGhaYSZdl9acu3Bj+tigptytN3I0KIFeEc/GbUOVE6jYZR/eyxa9c
QKXZYlusX/grj0jdPYw52cY/SRKQs+qvAGRrQbfVx2jSJdhYTClfoEchUaMMKcZ5
nawMLJ8e3rSezeUkhxDur2dEcflU/29+eFMd8iSdWkbmsOLfdgqznRfRUk6DsRcG
C0JEfiwd0pLwYuUXHi5bJow/aJOw1aIkvWqgD1lc474UU/DecF2/7OGdpY00QOiS
V7xBa+v24flFF6vVyABTUAPnKbsktXCmJrti14BDW1LOGKqSkom+XWOtu+FEt7iv
10xsy3ZfcieYddnIKgHXyzz6dCZ+9+SGeOuyOFlzRLnweUGnOI2PXAnFkbFo8hzC
DVamVb1MA3gyhXgv+JSY+2q4Bhv42/VSTToVsOTJNE0rSRbsNhkwfU+G+Gr/fEx3
c44OolkL8FVl1/AFLInF5D/yyk0W0c446nOe0Uzuh5Ya8fJoSMqQ80Iy794iA49P
Fw34xSBeMWnsvDAKcrzMLqH5TOO1S7e/SIYCCY7MBzn8jO7ZOrcIUG65DshL1mtD
ML7WKNd1aAq2TAaf6NAgCEJiKQg95bj+wKiwdgOuQaw9HOM8ZHjywSdpJ6i2d4ff
hi4VZ8s0ORXWN4D2oVZ/Ggoy0EYjsKWCLdqQ6vkOYNS0IgoBCrweEbRJ8ADgso+X
dJjzH8pjXMOdLmQBzFk9CdYL9Ftish5IwVZ2l2gTzPDP+Ze/2zPfzmAbeBqxZG1z
IqeDZtwXxVywoigPj8ApxAmLzvVpsK3fTJSg8NHqWuPPN2Fwn8mRvR9L7UQgcjV7
PCYAk/RXecl8homkHASdpLWim9rueB0+AzHbZQa/UCU45re9d9R1NwQXgQCBMbXT
XqEWLWFetnwBARe4KRivwwHWm8Ab8G4cE7WQE/PnUcyKsJxHX8ViEm14fN0SekD+
uVJ8mUzm5xXhnj2BBshTSU3aJeuE3OFX0pvMZNK3EbZIarnZQ3Z301WFUyohH6pn
QG80WLDSvtHgFMGINnaF3lJuoZbumsITbvRvQrh9Fp18kvnYGTSFDtP9Bx/Uvf9c
P/JrP9UxUZF+Jmw5WIeEUsTFxXDvfUvXxmswPogmEwueqBfxqNzC2wRnAlB4oDM7
q1osCOvguehD/rxEtplHWRtFMAyk5FgA6OYamfgOoBeU+qNKkM+z3bzsRe8CHKU2
ZQ3d9qnZGHZPQnDT8ThbI7b+uqpzACLvYKv++gVZlQ5K4za5vPuhMZPsG9lKcuI1
39NEYgIxPACh2SBP6UQBUctCsR8mxLnAHzhC1WiGHdJcEqIIEYkeoLDw4bGBFuaq
Ls6fgnYuvHfb87RrY3468pAIyNuYRXN/lINqMcYS1sRUNYHPP3m4NxuBs2folxG4
4m4LrVIsx6bOki0mqXpxJo8c6taTpeKgmVIObo5R/00licmcfSxUx5OsTsAGIz8m
p2eyuxTpIlQTGA2JalXvSNHNdHv4KtJQigyzaKMsyOttYspbKHjEV0Nb0xvmGoWY
F+rKhWTAYoq5QfNIlkbmOaRWWvog4LzZfY51gQVxkI5icQxuBCCp4ga5M08Ahdas
xvO5e5TBxWzbZ3fLtRVDpK9Fbvw8B+FaYLEIsxRkUppeVqGXrCDJFzixR7BrDAuR
g6XPIYh9fuCaAQmoYalhuj7vKkdO/efljIld5Bzyxi3ftRX4nsJPlCnoWDZxd3zF
d9BE5tJ0pcr1mzl0Ndc/dmVEgtSxGjVB1rzoOk9t6y/mJn3FEp77D7P+wlo/gOWu
cH1JeQEETPOCAwLqIi1cUh8suub6bmLDslCf9CZfXqWxLv0MJcpkFPP1DTMT1nC4
ML2KNpV1O+YEIWZQQyXUjD/bzaaZuw4S2cyUPNJoFCznk3CK8JdwdWr9Wo+vILfd
WRwt/vauqKmZnzT1QgCfaXRzyULh/W7NtiL3WnWe6YWyc2ag5NgYKXW0g0iDaNsR
YRZZR4MuLmJUQEzHrCkhh3SRZe7/pHe4buNCTctYzfyJTqZQMFEE1h5PQOUBbEyj
7PTicSPTeUByaEmmwesOla9G1Ficf6+xY2ZtYHh8goX8f5wa9tyvbQKiNq+ZgWk0
yKDJuhAu8nhv491vpAlpQ2j7wp5c+ckbrgbTq4jC5p2wmQGFQ8ka2lWHxjw978WI
XTU6RnSTCaq+Cih+Shmu5EbEQLQsGtBM56hkWbglocAZbwDGBmfff1DMVqcID3RN
MqYl9ayoH22ilYk2lFhy6zshjtUJ2QEx4hV9S7dLOsCTdiRrcSzud4zKtYOR8RDa
OTPnZIDdXdrUn9xxwBGn0LrjMkqcbPM3qQ/EaFcK3jm2vHREFaVF4AAJt9vCgO4A
KzujhnNtQ0EY9/iETn0D5Gzwfbff1BmOcPpJxEHWDTZM6QXo3hNrwUlsuZTRwWYg
fWCA37o5jeEBl3OJGEk/c8kdIh7UXD5vwlFFQ8rr7RsiRTeFOzjlXp+HWVtVwOSR
NPLZAv8OLMhwuY+Wt0Lz2geHQQ3IjGW9gVJdhLbKKpnuGrYzgMg14iFgZPg+JY/a
NMMSXK1EUiv35h3GETNUNDtjOAE5FbuB/xfugOs48/ij0ZEV0kJn8y/tNTI7HF74
QlMS35Pp/CX+jAmBuC6upp21hihp3TdDR7fnw4LQDH+WtskdUornT7Bt3B7z8UAS
mW+PMQvxMmDpBw9rNjV1iPPLTufaH4BCEWIhNz3t8Cm8KPzTtZGh+gcKFtdMGdRt
qQ9tXRXQQdaZrNqIECfDuLRFoR3CnjXJrTVhnAe54TAgF1CpxyBTNOQ7e4yF+Bn2
ELeoYEFpvJKNmNzqPS7H6Z/kTL4s5YRc6O/iFnUqtYuPcwt8fDKWukRAlIJz6JTo
a4/IJQRscbhX3U8CIe+6OkbtwgK+FQcfmWGuAZZLBSbvhjbYZ2FAyAq/RULaNBgL
L7xvBOwTqGqhzwyJvSSe1UFk4QhHIJ1GJguc8SLRQnjnLEvOWFLbsM3Fa9YHjwZI
ThgJau8TSV/YeqXXkCo5TFbUb7Esh7sGq4BrTNbeiUPOwJIFG6ZSFKh92rHwwcbq
neVS0znZMV0bO9CN8dkRWHWvutc51QbigoipIGwhxLmEUJN+cDqIOy+KMQYhoaOt
dDEzOBcaoEQTnM+P92INjouZtD7iMJBcWS9ZoenjXK4ie/5lj6Oa+G7tYK7oIJLh
w+j8oGmZoCe44LL2AgKsUi6kwvxsLp6deiTFNfZSm8Lf9E3FFaGxOAVb28dXeOSh
5bsvfgf210QFfKRfkBQNG86v2FoFvlaBpbm31tLuga+77Q8ZRyHMXI11r1mNpVlj
XkLRFW+tYq3dsQ7aBU5fQwr9aSdXNol5DP48AboAyDWpQ3mwIvggAMA71Zi8dqpc
4lTnXQqTk0CmmbIbfky/xck9oBv9/jGoOJA3CMbFuo4pQrb83ScnXkafqem62i6u
rL3c25Kju/gda2y0PznssiSvP9EOzxojjqHsLAEq4E3uECdDw6Gq8vC3HyhaMDnv
7XIqdOJUQrvu8ChZS2HokTZOyQEkOYtEwAXP6Piu5G29tvhx3ID1Ugv71qnAzRfD
0YarA0YZU69KPmUtu3Dejg5hhl1Bs6lXJ45svRJngDdsJGxug4O8UoiskgEwJXtt
OhpUdOtxeYpyaUaNzkOSme2BFuEFbakTj88JpaF3jBfjI8WV4FTWuAtXr351DdvW
nTp8gmBeCeP04xwKlllFT4p8c3j8xuijZV6h8KgudY7r4hsV2SDwlL7ZQ3QR9dBo
xfWP2Sf74jiYXMhOBVlHym8aLM5T7D+eVhPwqubSuC9vDrQYBPfpnolEi8JG1GWU
M5XhBJh+bt6rCJk4cBhTGyzHGIzy2s2S1ptPa5yEvMX6c3ge6rPZUcqmqF6jE7At
bTcx988aeG1WfkjUwDkh0JPAiEmTDlmNdkW/Bd2zqALqE4ffTU24t2zeEKKjJB2N
0HqNXZX37mglvdMHaGwYlr38O5JCqYyTcFOdgbGZgWTRmEylLnlXU1NwTXIm/zhV
vKtf3rlVXsXDCMZ60xTwoObP/CYprDe8MhTp99mg7EFn/Q/mgQDvUFIUDy6KGkMa
KLhhyVMvNJ/TGBNVBnZVZEP85XUe+tvGDwN4X0lwlWozQFb+oBa7WU9MfI0R+8QZ
a5e2JioddyrT4nm+XuyoTvmBu9ILPh4r/BgtqqHEZIp2zR+b9ekYWQobzLgOSL7V
P8LtKmsVbDkRO4GPEkuxqIFhAvsEzervx2r0CfsRW4tlXqVRUeQO0XkLBkDwPCmP
eeF65or1qxilwalLaNnZpFKiEgm9R5i8I3L3we5y03LWnmbEbWgHMDMSgoZsyw/d
Cz8IvibMVB2TR5NjhuMeV46JbYYRAS5MVrEO4//eY2CMf0SwLrlP4cdLnJfFudE/
Rv3ZopWgxlVTdmawjpUmFovYsbPjtvEPouwqbtDaxGqK501Z2xcxdfGCtTyavCB0
`protect END_PROTECTED
