`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jaGCpZp+kALE9Cb9oAkyNey8WDMefT2wNOI/tPYLibX3fQBZhRRp7GpX67Znhc7W
Tvc9MkTt8zKjsEHEqRbMM6kpbZfYAIQyk0ehzGAJnpZGLdkfO7A/mJQHkLCw0t1w
1QUOuz2z2JONuibFZAI3pkOLVBKB7N6mW+wSCQ2JMe8Akf2NMf/FV+5rT3YypAAM
vREGbS5YNEfiT/dR9I3Z8k/MLdFTF1gOx++P9u+yIPZG79OARFUoZgg6OzXDQoRd
3Tqx7CB0HPoEBa68UGSrFadWzYD0CFxJejLzRhjZMWJR388KoPi6oUDhmh/FN3V0
2kx9VtaOCu7bLVvWiBaP54tmm5hjcLNsH00vcqZhXROkhzvzzo0klBvktUjF9eP0
SfL8O4e6tOvCPT9IqJKqzqtFFDzgALNIF03XuUUh3b9aWeNY1LiLucLQYw9etfd9
hysz5l2IyB8C+N4AfAWMP59LzhNJoqsfcIozUIQD+02Tmom6Fzth7o8ReoBC7gUI
OmRXMZMNEPGSsrprjvDR8e0dtYvFPfXPYuXa9lNXrfH1/2v8pSiojhhYZN8MWu1l
l0+vRKhGU6JIqBIqXVanmeEqm8CbWOXfOVuZ2BjYTQIpwoqb9ae2KKCGA3+yj2ou
HpxpqsWeK3i2su/KZwY/cD99J+jI3n4pBplWIiT0rN4xuRNQoApketinAloqF15g
KCIwRB6NCtZamow1oGWNC+rVguRtnfcsTbXoN+OLV6uudvY/JPOem4cTmv6gzauJ
3Iy8qtwMk8xIgY1Z4D89XOFXJcN0LSRhiFjAshRyJVcL21PWQbW9v0bFhC4edLNx
jgQkwejDIDuBwxdDZC5CHY/j+y6XIP4mVrLPpUjzogYQgT4uLiarAPMAqPfnhsMf
hbd5ulIdbUsU9iAHeds9ADkqOvu5KQ1CyNvBT0fhx6wwq/b8KwThNxH6slNbT2hO
/AYOvgpHCUMzVkhf2i/AD2vyZ+SvPHbCRcaUqdv5Y8PUBdHEb4CNa6M5qQudzXiu
X91OFvPeojtxcbjtmYuDU+84p0BcSOLddILnXZqnRNJJXO/j0AT8UNJBgl977tKG
cKP0H35Us2dITbvM6stQh2NlYu7Sval3r4d1kOL1PsfU1jAltvyt5ebp8stON2Xy
5wf3ihF4ORn3sql8VhFZs9kCXLKQvneP5uxFL1t1GyrRtrN5VpuIFrba3i+wU6bT
u3txnrQ5MvDa3uHT8HZGQ9U4dyXdil/Hl1UFPujqEK7DRHMTRVWCpymS1yul5vFB
jNsqbLjEr27WNlsOwbCcX3AmGLhpoCinQ5WUxNR+U39JLLAUDZtE2sz27uqUXVOb
jxXZZvTfC3/lDy+Kpx0oSFCG6ZLskb2hpIT5p9f8bFipYTKvQ9mYjJYj0u9Ck6k9
D6DBf0zCWSjRcN+vgqBY61V5goirLaGaLjNtAL8K2S+mX85u66viI0MXhMSLFSre
PkUp0ZbU3kt2eGPf1lgpy7/IWc+z4UrTUIfgqWP1jRksNPYdksvJwWQltd5laJ39
V1lFx2wyq5O0rNbtnklV/3J2/OL+KYM10pjZJkuoQ5ebLRydpbxfU15CxJVunMSS
QOpDYC+G7mNQmANhVr9nsbgBuuG3Xxy6qcCx7yPvlteivLZYXfdFz6/DH3J8oLjO
nknG+/JWSlbtXNhOMfVKRnrWiBkknqDkdHCDOIbIZe1dknRrr3izVCg5r5meF+rt
kptLxHLj2I87oGSm5EnvKcENoA+Uf+IV6Wgg16fseNY5DoQexFGyGgehYYQP+gQD
ZQ+u9zJhTLl0dzhrJRjpK6Kzy1tHw1kjxsLuxPfHCQD7I4hkMVeGZDiIZgDs5j7g
m254lw3Yw0p9hY4cHm2swYqyuvB9S6LoJ/vkHa1/gmS4XHEJFqJeBybJlOrHIUQv
ygPMZabaqNeO1Z6QRovHSxqAYbgBDEm81lhZ2C/bYrjrAMQT065pyg7opeiX9mAu
gUvqkqyP8cSd1N3kYXMRCQvOmHIjj2Q8T8nzfjFj0MZ3obP+aDOhO1ekAOPhwBPu
kntHgW7G0O7e7nxEC8iyCe9ILXDRhesRDkdv2hsSrZpq68kR7JIEX1kc0QbREXJa
2O2703+DbjqgYn8/qlvZtj9oLFQovCl+BrrSAnLclWOWu8vxjRXY9pc6SjTZDlw3
wGuHiF8wLUF1ra9KrotyomsqSnZnPfups5YL8jy69HpqtiGsMbKTTIxgZC9rPjWh
4URNZilOsShstwOC1+nErIWiRMPeF4akRaplNJWTAK1FWTLY/op9jGP3SJChPWKZ
oe4ZeKcEmTJF1r6YIX2iiUhtH3lGJn3DAYAJgNTUy4u43luDS5ZLtYpp/FWmF5fe
zhsp4sSunWlJUwvK35VVOE9Po2q6VOrcTVjtu2VLTtSsolO/CdOGHLyuEusyzmRo
LUA1Lk4prm6Os9ngVvVZJuM2lSX8UiDWEvGGizhjyfyKKB/aQ0YYtni9/ik4nuND
0/ma8HO33fa/i4KRKeUpWlKasJ8xXXmqTj966zyvMAPW5TIj6UF9lQwNYWj1mn56
+QDY+atIxltFBu6CgaDtaiGkjj1gdj1ntd1Z0X48f/xGE+rWGYjrg/4OIfauYjqj
ufYelNPj4r+KizaaP3b2A5CSp1QwwHVq2wG+DzuJbceoFeDT0iV7VvC4nlBPabTM
qvCe3/feKtJ9t8drmAhrsKHBKQkKYAy2HEWjp3kn2sAWQTdBhOL+ywdm72ShTEsl
J7pdKu6VrxqT5q1NRM+nTTRQpL9BVK+e2/mgffzggbK91gZ87EXM3hmOWaLI+D3s
xgaWsV+9IJFrVaD17EaZ02D7tCkSVvW/coE2+ZGnm2bUdRKvcTzJC8ORTJ627hS4
EH+MbLf1Av+LzpQIyPOkmJsUkFT/Ux+l8hk++0wQQvykGJ1ltHu393K3EMc7Gdfc
FBJxJIf8iyUs/Rfas/WHJ8AK2832bEYMVFekMuppYRYqeEAnHbvGhxrpg/spYWXL
ySFdsBs1VHn+exy4iC7aJhM8xKCLfnbKkCt6Mh36KUFIu1lCDJw7TzUTAS9/lkOv
Zs5Wtw4Uj0IhrTCSVTSSB6EzXYmRi9vzlBeprQ0mhyE1d4kb864IZkel6FuRcKT5
wgMeL4vN2oT5eBch7ht8Px8dQ6AOkX73zmiJ7+Z6XDFoZdkW6HMC/HO/HeICfACw
GZdlhpT2XmIG3lRJJH95N6Vx+G2gVhoomtT7Wev8NabOohCpaiD7GgI/DxkAHVMS
G4Ny2fKf0MxTQx6sUQRqKxLFUNiWYZ0rD5SvS485tCoqx/onxp1nBZFjgTQhPBwY
y5FMwkfYSH1IZ58iGLOLNB75dn/HPqwoZKHDPBw4KOohmwkaQ0kmUVJVTSaPGSJO
evowTaAgMvcfMHtOm9kM3G7DEPTN4QRYRjWUeic65vgotTtxuTvDayaQ5TgGyFwk
3CmcPZPB/mRlfw+fmEXy2NMi2XvWHv2cBofYR74IHblQe339f3lPgxJ4htgyCosv
UQobr92RsWDnCiMIZgxo9Hy6FknfAqBSc0o0B0hbbW9UijOUKaszk4npdxH7qo9I
EZIxw11ujMyibAIzvYmkZDSTKEyR7ZAwDoqDinaZthweseSHHfhNyFykDjZOn1Tx
puuDzWrCT22gSTaMUNDnTx4noC9hzGxS5kKjpnpH5AJz0mXbGiYF4uBkVwR+4XpH
fPQh2zni2NGqeqTSdqFAJNYhNpXLGs2AJ7v7mqez+eG8HqppDNker/pQv/hPxg4x
D3CcPgNmWQgDlL2PPE/pVhbgalTgZUTE479fSD+2TSEvOnPfJ9ExNnizf4rVvA5m
75hW9VdK7ImudqQAhH2rP8ixQ1MfpY18urzLY2hOmB6yhNfj74ZrnvxEHaGMa+8a
b4tIsz78uMhLdr/E2o2flAelEFS1c3BssGZNQK3mbRcg/Phrh82bi6AnSoJn1Atm
BA2c7+pbzDzPGqeGUEA6A7qNmVpEnV97ddGmi8Cf3E4VlnNEVO+1PoL0ct9KsWAk
MjUg1UCeIHXYk+Q/YOncaLx0Er61U6QgPnaLijpvR9uI86spwyRRzCB4NgPwl0YL
1Yj0nARxE9VD4eVQpBzehtPG8n8G1Ho/jDssXeTfu3Lzc+gjGPwq8MsbCWBDCGSt
7Kz6V3B6vf/lr4rLlVtFoHV3ppESAXE3E+Oa+S1kCF2HsHkgq0w1Y0CAKT7YEgXi
4L6ZdtKCbjXMQfJvCeqpDCt9zwuh8PLQvq/sexP7jVuCeTfpsGs6lwKhGtzMC1ir
SQyH78HZPXinypwcCQN1yUOhusUN+GxYYlvZ7a+k/o0lSrfQPW1oLrW1g+6HqPmM
vcXZrdEUjOIxp6pzwyEO3bnLf0y/Wdp0JkpkZ6KJ0f48atPfXkjHX3+F1WbTUaMq
3d7jawfDZKhmtj6sUUV6qRXUE4GF3gzL2wP+BAel3MYsXVGfjzmq7ClchqxUDRDE
CqA/RE1stKvrHVWitQD0JOs7dm0jp0XObaqiZhQWWFLYOpkT3Dj6Gx3AQQeE9KRf
thMsUMySroUppJL/hOLV8dIzMqcV81LyiyT4xvWmX38LeeIbCeo+kZ28R2LfSpQt
/a90i7yiejPZWsA3PxPjhdo67A5EycUI+RmK3/qs2tVz1oiTG08B+l5tov8vRi9E
51cx3DiMxoVgl08xGW9MS4r+h+I9ENwwbQDLbC957P83gupNgkEkCUepjfFrGUae
ZIT4rBHK5DOqlr2lYadLPlbGIx1JWcNXCXWk7Y6cM9oc6pvtljLmtj7rHdl/yj+W
mPS6BibqAspTuIXy2o+PFhrwqL+dY7FKIuRKICr+/ug4Umg5O2JdKwPtT5lBKzUE
an+1CsFaCebYk8SGLw8J2zWDmhG0TQgYb2Po8QY7iZlGlYbnegy97/0iXlDiduwC
iU5hbHAVNP6OWidW3fgdVo3VRxURhALONrTFIfoA77NtZ+p/l0DsFikV0No9fMcQ
FC+bxgtiyknK0xVhVR3mDwyKi4+KYf15+JW6jt7Y481UQmxDMQrrrHz9AlZ9fmV1
2VtfeVmus9ml2aBp2dKoA7LkQ2G4XejUeW2Bgqq6qwH2QmpSfSP6xh2Xd6oZIcmF
5y5cuFjgH7B9sRhEXGzaAFvpMhQ9XVo/RR7jWURO0CnlBH4/30e+0BcfEoDGKsF3
2TIOtx2vyF5xIsBx0qbrsvArnIxS/Vz6LhTAxYZdZemA1cyeTcVxHf2fIpS+wRdA
cP0imedsKg01qjMaINxxLzN/uzFkdS4AWxLcvMLFZJpafsTyseAXCrY9fimDWNPK
M6Qew85XztVF4rrML600zryoI5+pHk8KbFJpHwU/j6ZFnJjmeq22z9D3gamHsi1v
LNEq7trqE6iMk/hGzmYUbMEGjBAYrWQKMzUiN1H1ZNtFrVvuGKvKXmIGPe9HG/Om
6ndI8Sx6wpFvP2t8vCUpwcbb6o9o2AQoKe6fegv8ZIb8bJOuvJYdi/MmhBupbkCt
SQ8kEqtq5RJL3nxJtwor5smq6JJxXw0MHFhqOSK3JkbkgZHOPFFcFqPL+KpwR3FL
ZCTQnDN4DkGVosVd4v7B37+D325tXicel05MMyTZUgzVvzrbzRGWxS2kqNNU5EZp
0uMxaAky38/TLHwm9Hw0yZqWd5K6tUBLl1aODM7D1lCONOpbaSMGOzpDNX+vHFkS
833ncd56+qes5KSkZH1OFzwwNzUalH8KxbIjMXkG9duSrVbJCckTLnRgC8lg/QB/
V1F4uFXrPxXV5x9QYwgw7IkShwmPxlnbAYU8QTenD8imRQL72Xl/r+b5uh7OnZzx
t02fdcwmtnVlPgSPcYhUHLsgwARpJupWl+4aIrPyetq/VIQND6ukqI4lMHf696Xj
0Ke6YmjsfE1clI3vtaat4AuNGd+XFHR5o8GwuEbAaokULQuVDfP0C8IB4TG3YOec
zTCPzYcUJ4Xq1DKffoAjZbooaVZCKMXZy/lDTmWvUNyZ/2I/cxouVzfOprAQIPys
/mmuu+jV6XZgmLDRk1BLOvuT8XP0rcubF+n7yMbcP3xC6+j8T6t+1qmmgj+7rwQd
QVTlN+ImHddzDoNNTYNw2rAPSPBBeX0aQXQxeToAyVtRgOmSiXyQWbyly+OcQta1
zUhALbUFcxXdQB3O9D3FMoWDM2Hv8QfqvhQCcfZp9lSHtUcV75Xi8EwktbaL0zSD
FOcVwqrL+CVIQLEcriIb5HmoaY9DkbwCqjuOi0/czg4QJgxCe4j5k7TwlelRJPvi
bGwffo9tKydRMneyhD0R3Q==
`protect END_PROTECTED
