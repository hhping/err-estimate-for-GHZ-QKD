`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tK8ZAUh+LrrvNF6xMqrg0UFi3+X/38bzpH5PPXk4UO1oxEvdizC7CVa8LVVeOo13
TMdmnOqs523oP125ArfCX6VZKmTMOIWr3REnFfaX7JJhME9KYv0KS1Ec6/3KbzjK
a5Sk/lKQ8BflYV9EAWwo7fslazZFS305EV4e1/AJ2zb9yQOjJhBdSDjTJK49Y1Qa
pu99liychqHLDpK9tbTKVBnPuB/TQuwalNSH0bCKFDHi/KQtbprSMMlkEx9uaBib
qKCqunAhdFFwym2obYdQS5BSS2TUpEj7LHD4fVypMsmTJYILhq5yz4Gys+7o79lJ
lXl5Ogg+XhSyS4WOmX+oDJVjMr6OdqQZjfDDqTr/fayXML9OMPToIwCRQw1pFo4Q
OailGLXutG8gKnxiIFSiOGJWiqCOs3rwYTJZzX+ZE0o7Wf1NfTr/wkNg/g01tiih
Bvdi07qa42CAkqjUuDN6149k1tgc+BEa/tVANUy+qsLMg9HVQapb1lNmy6JUUpc5
4qLPxWugK2RqAwDAMKcq5uqRwOwPP24Ab+ZY76Gr2vYwpNUeZf/WluDVpnADsXU9
Ce49wFcpylZQ1oT6KrgjTw32UUNBbIWrQK9IRXPzqmw/vL1uH5MHLfyrqWOb566D
9HnF5hLf4RS36ZLhqzbG+pHmckM1xGQ+7HUdPu2c26FALo5Xujeb3EoYxxEYqV4e
Ie73jkrIi2QjlYsIUbgjSb8nz41kB8MKzMtlb2bKpWa6qCSqWRjnQR/CDWQHD9pz
jsfHDqWfo3YHqcwAnt71w49+STCV5IITNVcm7yz0rD8fLK+9Vkc8pF+WPOt6/EPo
PvcFVcMQbUpwRWBJF6tKWpUBCWt1GujTr1wbBw9Dh1wXY9wxo+1LnpW+OWDl16LF
L5MRy8LLZorg5+D9Kg921DwxBrUR213SajAqqzR+6eq2d5uTS6RI/1NEjx52t3OF
aFiege/zBZ1YBFUFWs2xBQKEQ54mFIYkM22jK/E7G7lr427Wli1laAy5ke+0q0px
wbE7X3XcTjiG9JhD+8FxA4IoSYCh2gaLNMgxsG//3XrJsyD1H2yxY5Z38wY3cziE
k8bSWvgd3pQ9QOKNbOzXbsH4datjmeKxamcwRUVh4gEbn7ZrGYHZY7FC72tfwujy
eVoNt8xx5UMF1SO/H3tl/eYOnnkBQBUT+TipqeahbHc4TofWpIlMDMbMdavDa+jq
iuI3dqCKQpFirpMeYBus7l4c/538aZAd3oqtcOkqFSlUSi4PHvb4Tz9l2RMt4Pa5
c7ZhuVqOeXW5GlIWGBmyGq+TkfoQ10dcAto3t/WFUUIkWaO6RU2G+58oXwCPNiDa
bYiv+gCYPu+MZCu1KtO5GXndaPwY5Gp8ysdxXmQx/Q6BvFv68Vw7K7Nxz5sMX7jm
bhIe30t64/iO0M/WQPjwp7Vo4HBY2ppp+YyBsP5E1dqdBxoElwx6NfQDSw8LiIu+
SY1FBSLcYMnxt7Z7S0RmixK7RDkyVCTOLSMlfJF62Du2h2i/V9j3GUTMRFwCnH4e
r5qrxvH93ymxVWPWcWbmPJn2ucltDrUJftIdix0cfsv+eBOV9A35S0m0eqf3uVtr
jc/4Ei6udwp4KI9hyaxrqP0Pw7p20PlqjELa1U7oMAohd+kLnF1TBwcSJ7IWgJpO
gRyYxwrKc27TaMHv4o6v7Lt9csmZBOc5GHrz6uVJwsGjEMdvuNnFIc4IU7oSzYS9
Pmc9K64sB8rCyQ0Ywr+UnEYo9+uw0n/qkVMvrrN2GckCvCmpMpJnXVA8ncAAcNUk
pp90AWKVKHT96X9Gj0C9+DisVXZonmDarIGdX0AP59fXcbCIJo7mD47p08pUkDmx
PlobYELsZ1aPDpMUfv3XyW12HyKN+yLOnz9NzI/6BzxssObFhyzXA8pwwR070Rvy
/a02lIyr2sO5BX+xd7qJ7E7GBP2rqqREnRjR4tQ8yyvG65u6lUr2eo0xyTyJAG3N
RQdAmOitFGVPn+qVMQVjaUWBruS1jJVQTPT3eFKRTuHd8XOQYZFR3kfzlxV/FVVg
YHwireMVniLXt00VZ3X75FXUMHIVrOSr7IvDEPlpDvM50I+e/baKc5hfEvhZYir4
i2NrYkgIj8K7lbSe3inCE/kC7CwdnI1UlyAD7p9xq8XS1R74pCZgTTy6SI62DM3C
fKmMab/7DJSwUsNFa5IsQ9p7l7ti0qnYWY3LGod9/TVK/6FyxR+dep9vdTmlcrBL
Iw4c1eE0J416G4UqzaqT/SVYlkXw+AjpkIy9G/W3SRf/U6Usk+CZWqVu9lK/Jgcc
145UJZhXbUPd51hXNkVkh9I7YLlHlyQuEqi/dOCx5YAuyOyLFhebf40LbPqKwrTq
fMM2bP3ieDkUJbeIwI55I2QRAzf+Z/aG+gXqECHqTpZNIRtrcq1uyqG4iUTbUoIC
RhUVg9LNLSHAIwFIji0gyKn+FmM0469esplUU7BEyCpYEYPXXuXwIJozCe2vB65c
tX+PeWLqMK1IlzdyeoHZePSISqTVaHNzA08cJcwAlwBzVyPSpYnLvRniU1PIkCXI
4LeLZ4kYIymOGKDzI95ymS/nhB6/bR2dVn83ZWHqhVFm/3Yy2WuA1L1u5jfpbyts
kX8N90+zwMt05ISwhTIbOYSZzoOHZDuGmkpv8k2x4o3LFfvRv4vgN/P3+ZE93IFI
jw50pfNPDuj6bXDujFwT121zVybSWt5mnEftIQztFlI9U2/rd5IorjiUHvwzGHOC
D91J1fj9CcFB5I9IwM7TuRKyAQGo+LsyAcUYOsADZUyDa3S/KIy+DqqOOEQ6q7YS
fnumA2bVgJDinwjqZMWi2R9fX/MEykMDUPEjUvdXzrVEkWLhdbbi9jdO5VMJ0Ib1
VZsgquE1ooWnW8snlBT/Ux9pe3cDONMDh3rHFfTVfI448fxrKTR6Yb+Va4lhzLfJ
LLc02ZxXcGXsQQPyqTfIIrRdxAV6Z8oc+Tb3fzhJkrM1LpV/qt2ipc89yF7QYsrW
fKuM48tBBVkqdwLSIweGWyVErcC8Rdk4ZlLOtUbz4mb8PPn+QLCakpUPAkUFjvbe
izzqXBLUBg4W2gF7007l9aYJOrHB3nCnSVF+IP+LEnRbZpWE69jtYlmL06diV8/r
QAMr4PQ/JZesyFXissi2JYJHcmzeR/YcoFRX0yqmUBodShpMJy/QrgfezMUmsiBA
5caOJxZqO/ndlZW9VtHZT7hY35N6A3bckJ8oL2nXQdyOAimyO+5OfCbrhSogCont
U8kB2nsFlU1I+udR9enMAA0/xmk0ZMeAQ8neZALsFUzHNcxEIj2ONuC+oDHGEcLF
RPqY/rnYJQa68YQxiFuOq4H6OFKMlvbX0fqLBc+fMQGsF11ZSYcTA47M6esw/BTw
WPjCbek6ECHt0vTMNRVRP29+G7BL8fFthbKcVU8dsvaFd2H38w2QUiFvDXQXGMfg
DZyRU2Ew57t1SFNq9SPEIy6Jvrr3YapZ2CiA+JABnkPADzKhkFO7rbxFuYDNb9jT
+AeEajWCpLzKMGV8LNaiz4UJvqDnKcjMh3fJQMKLOQfyxIFJd6DLs9EkgOmxpMAR
FhoKbf6xEbcd/zury9WogtINohw2NF3+Z+7drLE191fU+QvLcF4IUGhpDTS39pcE
yESqnAjNAwFhHT7dUuBh2B6DXjAHDr4lHGBCogbYaOgIm40I1bcL01Bi3gk2LxKl
Rg9PmK0V00pw5GrnduL6kuyQtCnf5z0MVToc+TrqGveIgWcMV0L5bDFXRNz+lVvq
5Eabj82Ej5KZF8Opr9ohWWeO8VZnX040iqlGKbdb3Qb4odoNM4v58xImwJyu++4g
gCXGeYYP/xE6nOW9VP6o5WkfREq6yeYNZQLc7Oeoy8/toWcYY9RGAQZ2Z+TnShiT
pQzF0G/aWchfgzqbPZ4ja8ZkZTupA5XxwrIgthgXtG6SD7piMtuTi+jeeGQGTBUd
umQfCSQAfw473JRb8nc5ebOia8XsVGlBLA3ljy6nxKwa7YL91eoTA0y8zBKMyTL6
GH/tXnbBgq2CpN0+HQvUkth08XtfKnoeSNJMlqw2fceEjYzqD+dQUmN5fsXPt6TY
3bKWWgWCey4t2okpDICMbi2aYyk5UWY6jxvqbypCRznR/LUfkmOTmfKGTB7pyyhP
hOXFcdycvGS2f4jlCrXO0583VtQHADbaiDQR05TCXWzlw7OaQXWbQPhB8/ix4lcV
`protect END_PROTECTED
