`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0nW+LoT1gdwz4tLRo13z0ui4XVp2zWYPEQ730rF/h5T0oreDnP4H1pEeVKyJG2W2
hoRhuYP3gPv0iS5uu6kuXqF5/iQJoaL+iroSV5+JFxHeCh/Dc0IJEF5aOKXaNwj7
qCUumSV4X8OJ2RnjYJEpReTXcFJYGMsmX8oJuh+RBP/iCn6N36vQFPo9z/16fii4
i72rzF62OEZXQUgVY1ueuHl8Wlg4FddTGLZ1RwjrYXLILvNrEO9VnE/ojKyaWq3h
6UXBUtQQpcM36p8ybzb/C/fwTaQEAqNkAyYwPzYUVHp9sy7T4ICFle3kYvdMdNl1
yxNXh4CbPSXN8mbrIlB/LYKQ8QDNJ6J7LzAUryS6Mcu3NyLzSCJaO7ngwzcsF9Dc
SIC6uXYptP6ExYmjNkGEJCKxKFOPRFSva+oQRKlUQsW19r6RYU1+9zmRoSuDl86P
JZHDuCTDy/COPxAuOI1PhjWYASYFBQ6IhC3MoZ778E0I7xETB9RlkX2XqyPi4RUo
NgWzwO4pMwjX1FucEc0JrAIbQ4uxmpGpFInOz9UwmX0QzpHg15q+37XPH3mhIx2m
ukLECD5/i0FhB5p9gtXzBhmz40JZ3XbYzFmSaQbW1eBQETnqlo+Cz/wESTxbvMJM
sXZkcM0cnY2Zwnq6GJ+zM4NrSUYmiQHj51trMiGkBJHVBpheKlhJK7otD9EsQ38i
IgQGTq+dW686yElt04u7KMeYSm0ddJujzsUTYM+Fw533X+00gePRtNj2XiWsfDvx
NiDNx/I2hLJr2YAJeMrw8YaurQlVi1SFgcZAA1LBdcymvz/I7EBmIFiRnLA2b9qI
oEIRUTjRI9hgVvsJy2T8G66ZHGUZk42aJ1sAH8zZT3KlEn2qHzT8qK5+mEh6ip45
llj/rsOIihRud79565/VnyyCzcqFBj986+Xn2E+TzqQ+5vGQXdGYurkQA2RmkAa5
HYSZbijDSuL+6TTANX6dz5wVqx8Mfbl0jp2GBn7+CYAsy0TVHvMS3UNZThe5KD5p
3Az02S4+ibm265Ye0Dq3Ly7Hc1mV1Qe+Ot5v5nc+uRvQPCgmajCB+GZntTaDSXh1
bGFozQ/gTUHIUdPKCmaFbRubXU6GjvR8V+xnXpE8wKjTEGZMyVrlzIszU1ebNQdv
s1LXhui5608x/94mvw9QTO+QD6eHEfdGheTEM98lt5wfYp//my/QXoOZ8T+g2epD
rTz3VFcWy8AlSyUYKt5Kw33qLKI3BLw1Ou2ggaBAz3YFrDUCHVpzUqCrR5k7a9XN
MDAbkzlNNYdm8YYKkKOIYHU4OukUJuxqAnKmr+xEhAcSWEuxaooFpzbsFVUWAEyg
ARVqwRRoEinHQfZeT7e5bm6Ug1C3M3NZFydPUM0dtuv4bpNkgzndp3du2KfP8KI6
SqWd23njd3fzE9zpgmF60vPRRLHvXhstZhkEjPU15aBNh0LgdhmzNUJDLxwSqrcR
0l94AYdlQAT2VHqSacnX1P4NaQW6yaSqYuqohA1Td/fZ1TKMyig7Pzd3pL8v38PN
DJdx0I7rsBhB3A3Uw1wGGiAkyQZT7WCc44JyKzLRKDNnFE5PWcYErTu1sADqXTmv
3I/eacsLsFYPpaloZWw7mG/ssZ6FWYCAOKObIn6pz4Fo1bEcKigd9AlpdnQnU3jZ
DvBnoAEiLlcfbgpZrtZ1T7Rx2NxrYxDyDRJVT1XmHkNyq8jnvS35mMX3qvRPBECK
J1mTg3ejhRxLGd54pacWnj97X43/OWkGtdvYAJboJpGikWnGE4zROpblVvwr1BSB
sVB1bwORgTH/xhpFNKRW/3G1urwzCetLkX0dVSfhqryvJGPj/vxDmram19gdtwur
w8jcyJpJIq5yKRO/4/bj2J5PNSaZM1b3mPlZtN3tNPX4qe6aB4450uTIAhvfapf0
EKN2cesBicehtngBUsQjbNyVGrJVVYbVN5txCp5fYZGcsVgJh2jkSqFr1l23cUrX
mzLtcH4MOj+gAtNUGzUowm9NcktKt2Y0nv9WGKvJcw7f5BCmKNsj4lheRRAJG0iS
GKfH+8lFpzZb+H9huEgMjcqjYfG2rWAr9o6izAAR8WF/sZSENnwM0ei2IC8hiC2x
buwTaZCDKLDGqitg5ssTNumn1yaoke2ivbxPlWE+No8h9RqC2vQbRTZ1BeT40L+b
o5jAs81YH4pDUAYQam4vyFW6lZM/z9Kg/S6GczcwXLQdHacJ/ztxpUb6RrqnECof
kleS/OZCRR23+rFajv7sVfEBz5Zf99E/r5Juuuo1s3P3R3GWi86TMWYAZ/bRsNOi
vFWIpQPFJzNM86QXt1AcDSro9RTdVSgFUF8DChlILCD+QvSeeMS7mxSHYws1+Kqn
1A9H34JmjB35x9Is2XvUwtuYxpCHPfLy0G8J85FlPFrv2j/mozbn1GW+dtVr3YRo
F1Iw3VJ1E/6r0Vj2pInhvpN//uX/rwlY0635u1O5noONQ10KmUdhcxzBU7BEoUMt
yo7CEqCXXdUEuuuCBuRVlQoKEZpKhUMo0egeFkBpr2TApJFqmzuwkeKZiV1ysFcF
9vMhlDQmXMNbufjSQLAMXOk1ckJEGHWXFnSnEv5JAhbKqLnixn6nu99JXH4yZPNY
W9sNfDx/HdLnBFCDo/UnDEnorTEc5Rg9HssTK4JSl6xVttDiYJ3P1xUIWS4WH7wf
U4UsrvAMnL4aZJBbbjl0S8eo55Ug/A/RID1QySBS49SswHG/FEapZSJck41R+xRR
+vGkaKSehb7gegx2llsHjkGeRUmiuZIV39Jk/978EVcnFDL0K4PzahKGyGezJHES
imNm7UClLW+7CzCDrI/4+NJgPp0iTPqa7FVgVONOSZF8M1bRB5Esb3GounneFTsW
jHWQYmxjMx7NDgZc+G41tMYi5MbkAPETp17h26zUWo/7a2lqw0HojlXpfnojeP5e
WU5yP7PSH1G3ovN3TnUnIO1UWm234+0I32W1fguewjq4lGbXODgMJQay7fsvGbUl
JxXneZcVUsOJ9klM2DsSzhtpAG22EhRz4cuk33NCP00qaKAAjKmWFhTbpadQbs/L
5e+Vw7CxjN1KsmfSmbNgznWoGvsQYmX0bQcbVLCOzSQwmd7nnxmNCjGhRfsFAqow
Kp9DgwXc+SOGzNJEPvnFft//ziebOND7Wb8wJ9OSNsl6qKTHZs5E4hq2XiONDfbX
HFlZn8UVB7LgIpKSWty6t9aFL3PTO8q2iZQBjljw1FKswUorEN+Qz4q3tDnI50qN
lIvBbBqXc3c2tG0fRT+DQumNPa0xBwCrJ7FqkE67uLGCBroWaZ8Wd9cMifNnzCkq
CwyTj/6bD6M+ekipi4nJA0gfnIK0ocaJDXSAqaBnbzmF38Gth+1AZVyE7yqozKvf
YFR7vdQ+3c+MK+RyXePl6Jo+dm/ja9AzWjrlsOkQGT1Ma7UPCOV4R4MHPx6O/7Ns
YqD1FErFMTbTAexs6eqrtN5I4f2Q72dEffp31xqM1D3aGiruqAPJSI8oYoj3UC9S
uh00M8ndaLAJGf+JxolFr//N/9Nwlf4CgHF6/kxCMUHsg85ef8jHmjStkLylYh5j
Z7806QnOfBy4kaBJBoCiEziSJUUA9fI5oa2EovXVkkG7fwX14d0cUV1olrvQmYnI
dy/310quiQD+jsKw02NBYEab6jQbN8pNwhbSAYhkHJJA1S1lQZND2kVtYBKhR8dn
ihIH+SEUwOluiAcF0k/V86Cf+8OkSRHccBfr3KoYv44HyFIdLTs/27fdc/rX00GV
tityg4X31J7gbhOGiiGsSiqj7MLDnPNwWqIbN3LcFphZL+sD5AzizEWTRev6OrVJ
M7pcgIGAcke7KfWylq4yUNvuKNXFxGMPngc4G1/r5cegPnhFoxX89d3blPvXjYRq
7grnBV9aKXTUFxHtFWyRflSIFfkB/rQ6kzX60nLqqRygJ4UVxCo4CAHN3XXiIUfE
ARg5RYV+kVxIXcdpyqvXRpymHM1/9kpoWxtSFPABo00fkiN2LLxKT7VjQHjMIRsu
EKiRWKrewhls7ZjQOUNxHvprvt0lvozIOvVEQYLfpk2Ez5e98ogvV63ad0u61IpS
2d9ARfAT/SrCJ7WWnjTnG5sp3FyXB+pz9uz/6OnQQGjToWFEL1fuL3dOBJwvyQqm
Rp30tBtKXgsU7qJo0gv7Kk5sfqhPMG+nKruzSyIXUd8Q6swGTnJrtYY2vNJAAIJV
yNdSwCPArbgJubfk6+82NIIM27RBnd2yeOeh1iHB69i7MAM6tvXcfJwdSbTf0D/G
vHJCcYYP4adqnUI8Qs8UyUPeHvql3Y9mt2KK6v1F0zO27U1U5p14T4PRI5rkiu+H
z4a4YwRlOqxDpgvE8oho20A91EH+2zGlp75busVNbF5LCFzLBJIDYLogOEYYIStz
KtoeTNOuvirxPgw50LXmguKopmuqFZP3he3qriYmUAMUO7956Wh1LtTKYC/9BDqD
dJegX9QknwZC5YTs//dIVjD/CZ09p8+iv6/jhldOiZLIVZpgnHA393u6WkRuHPsG
wI8/NK9RgZUNh3Zb9/c/+grCBwOZ8I/5pKKeys7Skeh3gRxxDQ1Mf1iarScMJXIc
zzUSSYHEYexE8Foi1Zm4MdnBwwPRDw2gTMnv2g6NyLf2XjFIE6Hc6Ll6peS3/usD
5QT1mfWQQ5a3eV/ZoHHCPZoR2D7/8s3BdsXzDOvO35zOQFkSkotgjMEOuPnksVUz
WWMtSRzuGqDryTYdER1VMxvvEwlYcfwu+NgkdTQa6trItb3VUqjpXyDeYY4j+t6s
iP1fKejrMRJzcPrS4ES3ko+4jjQNjiereZOuBCllhTyH2iP/giF3JGC4nStBQC3Z
dwirIYhgMutAS8mWlW66FOdc/RuPtGU4ivBJBZYgZfFoJrSZcL2TlE3n/sJ2+GAC
PrkL0UampvWipzjK+hhgMQdmJGv0szdPqdj7tf/ox5sPbmnDg6X/FEAV6iDdHlzs
Tmii+ePEgE3ctDMbu3RslDNe2mq68b9zGnz15pArK1Yhp7sz7+QkLiee8MHU09Rv
hBUFeSG9qqJqp+lGS8+HC4j9atS6SRo5vSuaGeF840tlUQmlO+JxfLHjmdfsDg41
3gzGtF7sZ3xtqJ/PZ263LG5kRzQMya59MI4djlJdn3RevgGKKMykVn2hSSfihjjQ
0O+aVuG4rLWSW9C+T1Em3wRi9n2T9baApsOuz/fHGRBgemC3iSpmZvVjgy4s3Rea
hq/ZCe/ns7telznyFlVf6/TPQf/6yCKZjwOfLNNvPiItW1Rfys+RMTYhHsjStaai
bSiFl6/OJJD+JW9mQb2cnA0t+kp0eLFxv9PJtcNhVFkFK86tVyn082TgTDVS5tVF
W6iGOEfILKlBCgMMUMe4xWA+DvNQBqdr/k2OEKCehj3y1UA8k5qrbPj3quCXpTEf
WN0etygnKmlaQkMDSIdpc0Jf1ycqLpQ+vc/z1t9NpMcrKcYuWFMrOf+Di43/qm9x
cQR9zBPHwymiBOk2g+97fETytJIVK9hMWRwqy1aw28wV4qTH7syJdjlXqxoImxMJ
bsFeWcOZXaQVcYOnimrhxRY4sFgOZjluYz6j+NtcBl7Fs2L9VlLWNsfjQoaeJhsZ
TC11mJaQLfulbMz1FP7IIGapjX1I98yCvHS3k0Ap5qZMhIl9EiELBoLUUXjqJiS4
HnGUtPqvOc+x3N7ibxaqBJbNTcdbERia5npR0weNDrNj7yaxVjK/rHtiXbg7kHGz
E0O3VO6IjqPhgRnO3tUzJZ9fBjcMXCiuKHlsLhKf5aukC8BrkOihqR3adQ0MHAwQ
WAGQUhSft4qkzfGatTTHtMVTG57HY6rUNE6aQQZcVGU0jcpO4Mxih0lVIRpnAHed
mATYH25XcU/dn3yDWVf4kon6yJ8DlnlWbg4FWRFnryG/FSCZVyopXcFG3M3rrN+i
ZT4ZHgik9gx5WJg7cDhZyFOJJAKWE1y+tXTZ1hgVBPPZpxsA1vl4LZ6wqSARjVdx
3CCleQg4hU13mcC7kKeSZusL1l2sAHXTgKtlJGJXYQs+Du5Vx1Cs9zI3Gn8krK+9
AjMNw5pzAOCCK5oKL/M2aRywfRJsmX7HmGgCMiQELbW6HzS9jPZH8WBjzZamNfj/
sJ8MR9y778q04n6+3EcHiBnQ4qAyjpBodd2HOmPzzG0j9T4BqXCKyGII6YL+dZxi
cLs1Oms8yq6oN6VfE/kwXDKu5F5ZsLhhlEDNqn/X47rmhGMkNBfst0hXErS9gz3m
kl4CNga8/VPG2VOynDm7COLSRp7yZ5bCsyfJpL9S26mAW5Z5rtL7e3XiBBcT1Own
1PTzHcf1tVM9m3QX19ZrWVIA5bL/PbYtChtKpnyYca1ZmYGhSbpWvmAKBj+KFJ8m
EgXaVa+JciitSmE8VWLykAnFo2y/lBGhPvGeBs0JAwjxkoYcbfS8T3Yt0bkeu5H8
/DncdXq7R6eDUVW449RrGi0kTiJcqw4e1kScFr2TcZdUDabnoLUUwbZ29jEfrzO+
llPHW0VQSmn8I/+hVFs+qTDezjY/mDniRcUS3gDRIQKZ6TL44aazwhmDrmPZyOFM
m9dRTC9Jm6TA1A+3iWPKiJEjjaPF6phQ6CqJenQwDGALangfaUsXYqdY6h197By6
JVuicdrS9xV8LLt4178Q5b4lkIXmA7QpgqqWowhoQQfwJJ24NH328rsbqje6764J
vs7y1RJ8n5wlZLii/VcwiRJv0ito9rqASjrXx4ClUobK9uQTSwtxj+F0BrU96oiD
1HyHQMzMOHJk6P7gVpeAC3BzzIU/EO53mBzH+x79sFqPxrSw8hz08mT7TZP/m59C
S7ZUEHJv6+yBupR6RKCdJKIDwgWa0saZIg4/hsJFIsOJ01eyCEifk8/9Ldfd/u03
ojYjfxhxdfPjdWeepeVIQjdfwvr1M+oQsPE2pOq3xJxvcPQHPMHzDkLm6WfAbGxd
i3+UpQkIWKiwroNbOfBjN/icZ+c7L9HtLm30O7Km332g0Vk+X+GW1hHFSWK4sP71
wjcs07JN7RmbEOfMkVOKMO2HO9dgiyTN3SJZPfUqVj/FUkxW2Z1V7VSMPIn8DMVe
n6YQiKU4WhkH7xYNRwklu6O9H1sXGbn//nDra/u8wOtY3/wqZlxoN72OpLf0hSl7
negj93sRd7rSljzBDH+v2XXGG8SyqVjUh72khLyufiMJMDt9U189NeM0AH4wFbJD
kONzXHuPKUYsVsVh9PvYv9IcoLvJWQwhpDXYnkiqxtuesZ/TVNJfjdbxr6RqyNWg
x9XcjKii7UmxeZEm35ocfOqjjbNFXwSuOJ3IahwoZdnBDA0Vu/ddYi7HnaKBKbQV
6rKqqv9fjgVKkUGqw2RbOZzoDEcwWJWGoiVPxz3G6XrwbxA0B0c1TeJxGY49Rtao
Ivxc+DinbQFM5QuZP5vvuEJjvErTTP9sEV1bgu3ZbEe9w9v5BBd09RTpda8gndao
uitdlcTEy0XbkVUxiIXKNqd+ej5407QdFuEsk+5K3lktvIceTrniSAu8HIRBH1gI
BjCq1NGYdmguQ0Xe9F9AxzwOKQEzS9HCQvUJQr/R1XGdN0Hd8S5cnf7se8pwRhjg
Bh20h4kuSiib27LPgsacxdrldVk6k1wSoEgs+55bzPlPV3m9yKneMFTXcYwnniAh
myRHJnFZDU1+FKWa41PqNMFFn909WEe8zBBDABWW4TtqcK47qoozuNm96SQHihPU
I31kuBPCLR2xrRce9GXRdNZVtVyvI4QoufgGxWUZ9FwLbE7JgjhjQiUAIfUDo8ya
zSuul9dlmUSK+vNCZ1eyVA4K6sKLFMOhVRbNiGWOlvKvVzIcWXczGXME6/hNF3E1
72SNWBUDDPzhMA83lZsuLn/Fde+kxG/0jdgLx2MAFg0PMbXyfJ8luRAuph1y6u68
W8EClAiz2YdDOTh7Qw+2M4i65v7KBNTp4vykoAnap11L7CmNoMVeWIntjxAObWte
y00u2wMWg+1CJqr6lKcjdG7jPZLqpX8BJcrilcD1w7WJjwc8l01w/JQtOh9nvMHb
wNcrs9OfHUj4XO31HyJFbv4MUJNYhR+bmTSD6a7bwZEhZb1o9nDFS0yQQJFwmvHv
7AGXluA3sdbw/s+rBOmp0lsbflnO6ehI8blsfOCloheQEYC2r44dlntwro+y9YGp
COyls+On7boA42DCs7Mn3CjFrWDfyH5eWGQvy59pTGZKOEM6UXYm2ofQDme/jbnk
vXws/W1lOmdZ1Je1vQC1nsQJ3xEEEBIRe7/qCfUDKHzBAQ7xmulj92mnLdL6YLGY
h6xzHXCBXRaXhepgjDeW5b9oUjXuVcuqAys8aBjNVJmwTFI/fwitCGETwcSBhqMr
Kkkwh0zG9ewj5fWUVVeBEfrsfqPXUcwXmqBk1YDCGxDmLgHekoqlWNHnar4QyN8i
bJcxhDgP7pIZ9Ur06ja/McqWzu/HITX2e5xL2ycoXank0S6Yrc+lxzE0/soU+4vi
u4gMxTOsd5JIxV1BbKkqN3j8sbbPpWGDIanO9kv6vegDgHwPU7UaEmCAfGLwd05P
El0u6P/gJxMpIf7sCss9FYxKuBB12uFD4iyp5aOP2ROYFId9pjv9kiqScBaGlIM5
7tJKO7Y28/lz3zd8MEEE3V1mmE2NMVEGNYsqyJQ1OSjKs2ZChVj4Q4PIWi6MdiNW
fIWo7pocL+gHmY+s/e22o9y6jyL9opCg5VI6ovPiEYy3oBd00Aiel1GdsenzJPmf
Qqfl9rE/UUywsgsiZyU9VWLKY5ZUdTa6i7LmsQHSefgrJiYVScRg+ywaqrBcvX+1
hMUE0N4wjWf2rIyxahPOgsfI49yU8RObezPQQ1W0UxTegRPYE9CUUFBtLXHXWiQ8
Ouc+208fg5kB7GksblArdj8+K+Cb8blrI8jCdmjk4mNHWjEdY5PNcFn/Zi2t8JNO
g0Fd7yP359i5HvZSWE44lg==
`protect END_PROTECTED
