`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FrkI5nmkxoghqGVaoQfKAR59M1LuR6ilAt8MuyZJCQe9EDUFPk5Zex4vNG+hHVHN
tEAlVnP8xGASe81TMK7vEsNQNMO5ZjWCQFq1lYSkg0LavaxKNvksV4AXmxi2CPSn
QIc72lHgMlsJwvHgvQYJb5IaBmuJwHBV5w7dsb1ACdGboOxD+6lRjYvm3vVE/53H
a4o5NUGcTjW2BjuJfxho7BY0ZPArrbwk/kzNHjL06qezFNRyL52Q6zC9PUMX4ZJT
Ivd4KOlXGAiJrr9xsMMik8bSD2/LXGfDSF2bQp86HtEmlEYH4t5QbYJ3JksHEoIN
5/5Gm5AkuvTx224RmZYW4ju+K1pgrmb6R+Gbj2dqZuL1AohIT6LeP3Sc+34oZghC
yfqsSawAL/UtK4nrqIOh/XMI7B/0orqP5MWIXMq3D/VPtLUGwNzJLHHhufO969x5
hiAnNkx0o4NQzGIwuxCa6i77E76LkHJmybvdb30gj8PIN4XW3vHKZqwXHlN0nVXz
QdnrQZDk/jMTqnQAlevr4NeLbe606Ip7MHmEPPjBTv9KSU7dIQevQsda9v+nXyx9
S5Lrac4ZKqpxZLggiGyeRodpsh5crCm+Af804151uL+fns3oqXqCP2ovtwwiRh7N
1EWmGVEQsiYesxBvMafvNhPwT6NpT4WFdluMby65VNluIUlPYuIEpOzotGPSIg/B
T3birblvzLiZdgRfFPDFHAh37SCSSQ/OTKx6GyfZGrM/oKtBN8oWr9d4iLGG3nmP
4y+TGALFnh3uduvg0KfMxj0MHH7qBM2zMKt5Wy+ybXYn9HNQJImhW8a+tbBqOP5v
acYcCMAvihhLcmzl7GM0jqpaBaKP2ZIggV4rwoYPuCKgb26LW3oujF3jUwWpuctk
+fFi6E6BtbEElMjV8TZztMTZ8BbNiBqGrjc+Z7k9ZFqk2F+OtR8pi2C6LT1hNUcF
u6aAjAns9tmtwhsUadgIiynpQ+AjB3KdeE7Crj/nKOK9+xuFkSnfE4DDQaAhnt0S
gaPKRyH7hTLaJ4D4u0rkaFs+x1JAW4++AaYjZNvIKBbV1TaOsUamCh713s7+J/gT
Q3HyVk5CJVcqkDk7LgyvqsZ3AKFqUst11e9c3mXblwE5190MijcDd10qUrtH9/wy
2VN+NO4qCiQamTAjLZjUXLKcGn+k/WJWXtdGR/ku27dgEF/OwnhlyRbWahxejVdy
yEQFUX+v1kRnLL3VhXq0ULvpsvV4A+7CnndykjyPYNB5HBTpkoimlllZLyM3HWVt
d3wOi8uIxmQwVTuJ9MTuxBGEjPPvlXKO5VO7BqX6Mvrln8UUtcybtOslplswReyN
YgJXBLziUA3WnIDNmGfbt0Xq9lEPj0/Fs93SwLjKlmjHUjhvu/vJfOdY/zFYFSBY
nSsXvF+BL/58UnvJdqN/5qmp0vADUPZPQdao9Z8V9VoLiEeUvZ3+TPttVJ+bs2Zn
MT8yNYwdB9OR0weunBn8N/70MgMkJq0nl4xhNjZTiRO+IrCIYpkVzUr4ojp/FoW7
npaM0yBKMRDZx20zFirlmRQHGBeEN7wBaI4Fy2W21AEXQZgV7EryofAPieiH9VTG
viI47emPz4lqSxJ91xNn0wLMkt1dxxCFx3k/BAZViWuLxOs2FZvKgDi6N0580SjX
If/CvjaSI1Fz/EI1MpOCy/pgh3s/h4GSiajCbM9/I22yWo123aVZhMKL+wUHDjIO
`protect END_PROTECTED
