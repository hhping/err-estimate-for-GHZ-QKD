`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9BFf9WkdlhNNjerpeolEZlLMH0iaDFSfgPTPEnrI5LZgOf6Z50EBTQLcFDUtDYfG
YJrOpTCCbzd6wl1pLqgtvKb0oazDIksqaQm4bS9TDtVLjuG02uvbndw8FabnnNpa
vzACWn4WVYa7wEjNnC6J/y/OsVKLRRqQnFMcVSCEDK5zJORgGMmstXytj0hhvzzN
ti/z6HmJvYAvuleU8s5uASLd0i5cjid+UrCIe3LrWsZwjHG1G+C0OTeUP8ZpeiOQ
FNDXh1/LNHOfeduCINU00EcyonSRY1mgAAsbrVbLpMgqUlcUWRt7d8CTSq3VishF
h490uokTW68mx1QmSeRptn1WBLp+Q7CsenrcmYYXO54pd3L2yHWpl/gidnvPE7hL
IV/jGM+H9FfnfFpZpr52ZmzkgptfB7oHZvMVfoSGOf0pGi1PiP4CFT8DMk567Mnb
WBI10rkBl43qac02PFJSoqAHvHpxgEQ/Ik/cRtLqwHXNKgfc3Ygpu+jd01rtPPdY
sneZFlUzSp3KgAt7+ebJpJJ9XbdWw4g2onYD0tvOQw75G/OlRh0jZIy/y7V0pXAW
Im2lyt1BjTicpJzwUWmhzbXPLzgwk5/yVH94Ifx9bXHcznV0+D8EEBJyCsGOiBQ8
SNRue9mlmL9Bxzz0cBnXrXTQinvBNb8qTBraAIchMO0wqhNV9GlRc0dztygdOjwR
Cyt7e/64rbdYSaTMfw7URLIf6MlqMHq8LwLoV6t8uwTvvASQAWWBaEQKJXWZfhN8
dSCbho3bkeKOaccYOn+q7xz+diGyY4TizyhORFyvUqg=
`protect END_PROTECTED
