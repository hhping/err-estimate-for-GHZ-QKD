`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PO+NyGfxUifAmNMQmWeQfp9IcxBhRZIDr0OyZGlDMvYhOMej3kF7TMyi+njUWHOo
jWeBAxZCxN0+36fJ31pk8mPA8OJcvYOcaCm2GLV5GaA12hAFwgg1sYBanYeSpNQp
5GBUCVx99G7KC+u4BwhBt+7gbrlPfQe3mY8khR0cKrYmmL57/14ZYZ67E21ADbpa
0n/e9aT+3lXzf3aaR+nv6RpggGwAR0k1CDALbHiSAKq7Ghf0uUm3ifrkaH3oMvRE
NTb0c+PFbuE2iSn79Gx/8Kh5Y/+R+hagWA/4Qq1bsdR2PNZR8k54tNshmqeSHL3u
A3ZAKlLAA00iuat4ygZgZhiqHyjivVF2LH8ZJBoRtrbyU+ywEYjL7DaHTfBpefot
KlPU6cbBUbQ732WoLzBChvnPDGP0udBM8g94vmx1isuiDm7+rZvlsX4bpCXyq1OF
DcFShsLNv6q2215UjgLfC0BQt4NaUIJODW8ZApZraIM6YExzaNAdmVXsNsHizkKa
yM5bSHUQQL027mMRUVuJ3s27aGqb80cRZ0JL8jDi4m1UV78wMmmBOO9lnVzrDsl7
yvbi4hNgBfMJNjkE5XwqG66oAxKta5AEIKeYTj3mJUabqJrg+AGoxFvZhVLAtaGx
SvdP9km7uZUxiwWIyqOe+j4XV3wWt9DMRXbQSwDVr6pnTL5K3LbDEiNHq4b0XbnX
vqq9sflkrZLtejCk2gLNBSOMi5/a/6QN1FkCaEiWNNeGSGZq9ZaEGjaZFNuOs7Km
2JwuApxPcy9+qdgFS50xXbx617ukXhrfucIKlbaI8e5Hw6FUzSqEk9ZVZwzeXTw/
nair6IBxgVkbMoV6eIAWRqKPM3IeRcQfqTEPMqNtnTHi5oebr3WTXYkbm7pvMzVB
yDl8BeG2OXs3ThvXaJHM9pjdkykwWDLhSIFyrBnaGBtNciC7WawxfxVIgEXGCrW+
/+3joJ6BSkIIzn03r2Yb97WNOqbkSNbPJPazqPnY1G9I+MDra3dVz+S0+dKZUVEr
yHhwx0bgqAMijLN+k+aQyh/OdhJBeoqjMV+OmO68BsitkULtgegqtgtqdweV++Zv
s1Chb+FBhkARt3HPQWQDMCX7wy7EWvLhfGL5LKQYpz5pPuLAxtMx/1WLl0gO3t4t
yYSsCFm3Xho73rm1oAC9N9/QTXdCW5Jr/WcOCxnISht0ngKGng2KtDBEmAD4a1Hb
CIYeCONbJNOumeTyEtIORnyecGC/t/hCh93W2vb0Q2P4v9nmVMKNOAp0kLM+nfyM
JuoReOY6ZLNFFG7l5UsA9+2014i8nxQNm6Sy6fEYSyqjaPC6S5api57X09JpnVIJ
2MZibDq4ewSKJeY8Bb19SRSJMdjsPeGqcGFUfMPLH+h2S3nunHxnvScBV2qanGSX
/oscTPLwuLBwa71gpoSZ71IE+CdPlsa88Oj0puC+r3c2OQKHKDJj3LYgEEuSo8Ry
BL4xO7ks0DOoCwZ7SJ7iQKE4d1DJT1ojCAOn5uRabrAtsgyqcOBvZcn7b66kdRTX
zgivbplsV/XZpT2ll4flrCsj2+21wGIKjZBpnFa5p2BmbbaSmFaJ3zFOFtYBJ7TA
uEV6vovPVI+svpyUI+PHolZnhrbD8sK21/2eiRzuzH5mZnoZszyi1SnxvcP3wveT
vwKMTEkh/OYLtkxOp2nYr1JPypNSj0gjBm3IUcmLbA/S8pp8cSAoZJn3Kr3P6SZ7
cNzygJckCzebwUMKr1QThntq4DXXROtYazD4O6YxM8zPjU5/+2RXAEDYKWfzDFIB
32UFdjfun82ZILQKjYEQtPM6OGfdykv6AUv4RsxoInkqksZ/6fwfyDiXjVJ3DHz9
APSDDmWn3o2TVBLZUhSqtZUqv+fj7kC1BLvFkfi9mWhNgHRwqSjTmVquLCI6D8En
wzbhA6RiYa8nhmYy9dFLy4c3AonpHnVLJ0EXWpFfd3l0/Z4lKNYROksYfi3Yzw5p
oza7JRf6AmHiAh/zUvL959Nzw/wDsN7c/f6ejwI73dP3ZLHbM0iNmwsThvcmi/hP
fs46+t4j8wJBK29+Rog8XVGb8jjg9lnZgY3kGC67N+LzFITE2Ei65IPH2mL+PzQY
RpWJ8QosTXtvc3on5K2U+Fwi6T7sXHITWpdTOc89Ff/1mFdP+sci3ajYKimyX3FU
VqwC76h60gs9Gg/24A7yUea3PsrZBWjLeVYnf7ODzfro9Tmj3t2h58d6QTknOEw/
MOwL2gTE3Ozmo9s04GpJcdEiqFyLE9KtY3tCMoayextueo95JCtPtxAouOhMMzQw
62U2B/WoUcNFApiv+75ITVhtcjlJJkxy2Ikg5tsypeWF9rdCs3pEq1s12Wf9W5rz
CDYMrMos++KSOo4ZJ0GZ8agd5Ifq5lWzvedYhhDtHZyZLYia8Z+t+oNQylLD1KSN
jsTOQOI+iGColxGNpcuCuKy+JtpssXjPA4aQYpJK2lCMpqPvGbgX7fx7abNUMdL5
5+Vq3nkydp2G+KM1kozMnwwfEXtXpbM8TeyI5d7buk1l1Fv7BfYltKeKtwY0yC/o
W3YX0JIzPc6ztXTcVY3/GHINsxsJMM9ZEADVIaX6kYQm1lT/evJiTysU2Z82+Ace
kEQ9tIOqSAfkBfzaPKTZvsc4D+1yjsXKY7R1a4H1CCVim/TaaXWDlml9zc0plq9s
4kDNp0bZq/wUekZso8ZhLvJbrx4gsyd3rJx4dtX/aG3TurOo1zo7OK7TF173osA1
aKGu+TDkKijWW4rmdkga+HOMBxE7UGBhitF+yA+UEl9Da8egJ98Vcs4uSlb+Ymrz
0cddfjYVfb6Ordm1LhtXoErT4LUsmPMtvZrQgxW1fklfHgKtD1Zt/F4d3qlE+qqp
TPWvCOHLadxyT39wwr2JTbBBzetf88dC2ovvfY9j4CAoLhDV1GgjHVJfm5KVMo84
iLngOs91QjjfZSFE6B4VKTEb7MRz87C1dQ4+z6FFVYhKB4/+F3kcpxlc2RhmcT7J
BqAChGlrvTdZWjnGjzrh1UeCq4dXuzEy+pcYEfD5jQbADYfwfYQ8e85/plMuEm4o
xcOrPkYVLQgo2IrmoRsP4Kaf1SSBQLX+JN4bGGYgI2KHW5UfmPSsCRcdIicQZZe6
a+JkWP0IAHMHI2ZhiSz8S1fGxImPXCEcE6wSqZp8qKxm9mZ72AA7oxiVXMkqSvyb
zl4QKPypRRGaWkJTFRpGHZBC+OfQ8Y8Tu8ylCr6uWHY5ARR4dENlgWY4pSAGmila
E7wSNKoBiURGasx0MykfwrYK56XIDFKsU98oGFinDXsez8xDV5uyVDwE2lCAQ7HL
QxsnEuVPVhlUQDoVt7i1ErA5eJvI5aPyueeBjkhou1RkscWZC69F5gf6DcVaes4x
brrOsjUkK+pQGnc9wtcc5fypmM7/d8hgKq82fEnEBcNzRbJv3yzdIRT7s7RR+ZTH
ID2QDqZXcXcIJMPjtgZeYIBRRfrRKWKQkgR0MzSNIxuAa001TJ0cBPxCys0aiUDc
BUqgLZ/JuG5WfdxPfjMpDUTZ8kstkJVS1/xuLLaZ/4Ljrr20QVBc4t7cbPXNMlqb
mFH9Ld3qL/P/vMZkFusPjD2R7bMkGMy4TjW0QiXPOqZ0h65kpdV4zsq9mxbAdaaz
MjTktkg7jko2MeaK2+oJh0O2ljBkZ2HNPWiyl3U/YrsxaKAHb31RFab4pKqv1cSz
vzvQHL6P0AtjIoS+1ma84qmMSd+vqRxnxpbPDVVSQYbscSAMjWgY5TUSIsMdDl/y
gunrgux0k3PyUdT+D1fkHf6e1UO8l7Bql7CXohPliqJ7aE6jR4a414N2mqVcaCFn
O3Xz3lxUErOnYui5hFfgnbWo50zfW0wN+Evi6jEA+L0JzMk272CSfjFbpsiDYYk/
+1H8K40207hgIMmqmJjjViwYLJe9PDF8WHI9KROPbD2Y5IE0FHRSz/vHXCiqcnAv
rI6c9xbnUClbovKHai7BjZ7AgHTsPjTLiGkJ+lNDgT7sAzSdY3Xfloxx5SnJMfvC
yTS7r7CDzwSDQ3SJHO61zEbs9Fj4mZkj5OyC+U/cZQbVJWyUlPSxhST51Af9uIft
agjjEiFFEWW1MUjRZKwiWqdaoxjFFIjiO7T9yEFBrcRLzp08yXi8rwGybPt3BUrz
fz7BSK4PB1QqztmuFh65E6BWOVS94eOyQqjOiVlAMe4g7zEHx9yrrDBtG0NrzIYB
z+eyxEsqhuVTAjz4lsiBP1BRLdoZ/MZOj0xTz9wsTfGnIhuVyyDrKm45Fp9O89e1
9BeOMQFLSdMn6wTmIr0cQqAiYVnCWC23Ts+yo8b8JFSqKCJMOLzFP84gde5JfDm9
pPTs+95s3WTQE/RNoKvFdl1zeauAAhPl7v52NK96aw3C1/hZbbkDC/n4FjcZ7Dmn
KQHByxdVye7GQgmEV3eJvqhPZg+Lybadu1zA/ADqAT9i8bxrI9EyY17m+bcuc0im
Q80qd/MxnDMJOhpHFj9O4n49j/RulmO/RIIXbAs3CF0uGdJoJkDR2G5fthgHUFz3
fH2nCK0DsZZza05oo1llbd4kZm1UucRQ0ErR87QH2Lgj9GAO1t9oXvooFuy8e3vK
gC5hyfEwfQnFTX8dCw8xtWexVsoKjY1AEUNZqS5B2oUrL2LTAJNb4+zTsymR3kMW
KltbPg2EtyZ/arc7KsLyr23dbK9oxLJVMZpLbwZLgWw6zDQj+HnZEI26vTVQj/vF
sZEWYPxFZLAoW4JZV+7Dd22ELiYxla5Nfbv0tlRoPfhTQLOwUvTpDZhWYsUC7iKj
2VExJY1BsqYTphOELJDEMaxuITD310Z9mVb9/2NwFxFCYFPH9urvSXxa617P3BR8
aVG9YH5uSNrGly9Ezk9Eh2Aeb+7VpTiF6hOVfX56A15LkAa42ZPwjQ2Lh3hifQ+q
7P97Ymv843/yBNeaEle5f+4h7D8ieLv+FwLgWk0pd9S+YXkk5Y8hnhiYmyQ3AJDT
v8XW3Uh5PxEW1YVNK1M3APwJBXoyksCpUC99wgrGd1P1WxRmzpQW2MpFfqqJ/elW
NB8ul7Q3daDEXffmMkWugsYGesxxVB6ai465/p2dH130/x0n8KzNwX8k1SB0zJMW
djRU1yp3NV7jYnSPmD8pfS4qqeneJ3iBZYhS7C7qFLQP8L/Nr4uC62DiNOcM71xV
qlmPMUYLWErkCKN1EYXYRx7kexihNi7z8FnWnkCxKmC2HwS+7yPqf3P2N9pv90Fp
WlT7D6MKkIzYAhe9WquMqUe0V0MULumlp1SYOXC8YoblPUOK6bwO4zzfWYQwyJrd
lZ9hBLpJ1pGQLe2NAO8aiTz39fFpagRv0cK7wnjmtbp9CUnXBA6XrAFDF5TH1IE7
U2uqMik9Zmfjb/ci46VQLdfq7KZqzBsLSQ/+NfwITSblwGGPva0hEQPDbAmKZfI9
LgUg4/8QfdejwNqoafaDMWeUtZDqEgoGo2RKCtWJoToGJmWa7EpzGZ6NSjhTQlsm
iDlNyoC5XVDJyGK2cKKWGHPIdJP5M38Q1QogqVD4+PIT6WpMaPcifed0PcTwNDxr
sakFFEw4JvKt+Ajwpq3XQj+83wxvQY8AXii0sVkayqyp8WmXRH4acA6QkLrtDTHD
mZY++BS3CsOIhCRnZirRTsEvtsHxAfcBgNJLwce9yxoKuqR44CF0sm42zw90qt46
auz6igXhFlqtTNpQkccE+RGHkBADvVteMtmkQBKXYZvJ7BeDklDrkvEFGSwcqSvE
g1WvjUUBA0kg4tT76hKEFn8hvrumED1sRCSEkEyEO/ZWJAOd7vR3vVNpb0qe5quo
uX5XphUzrHgzgLPOhiDHPOriqGH8TJzxrtuYUTK/49Qk7yf6+PeERdNx5RsQh5DR
8fJXxB1Md7vep4YXCixd2JxeHIRR5P7B013DwSiRAftZ3qDiQFmXI9SxWJneDTav
vHtgYC3byWr5PsVy7yXFsoHOYQDWBy2uWTLMDKUihYSqspcvmM1byy+kM6GaYPhH
`protect END_PROTECTED
