`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8SINpJukKfhjQgQNMmvXrf1iA6PNF3UKxsh2ePq85J6YWUV/U2Luqj+QIrYLaywV
QEmXRXvfOaAH7B4bGmWL6GwMPDpoaIVC/CKUh83ElbA40h4IgyJWun3MBm8VP82G
x4WMLiIpH9Rm8eosUUWGqUeZSFjc/HXt476w5KNcQwwvLgxWmIelLAcLk7RBhsmH
DQnStFQA3JaS1GCV2x1QpLW2sgMKTFyfJjqi1t3PNtyFPt/awYcn6vdcAHt9iODz
5NoExILORwaKl4Z/6bMOy5I1wkkLsAkmlWtoiZELSmReN0JsOfEsYCowdxeEgDjR
3Z0GxkzGQXHYVJWezOoZnwi+L1ZfUZyN/1ppboYg2Amf+WqLMMMxfyO6JIoqr1Bq
hWK0MtzveVOstTV4OxhkoRf2Vi73FHbCtWaVMS1DvQtyGJu3VsKQ/ULW4z8Rhylt
RtG4FqRT0DzF6y5vPXY7sA==
`protect END_PROTECTED
