`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pvycKdumO+Rixpe8+QZEBrhli62ivEXokm48t8ybcojuz0RYI/YgZvF7FNihUBAC
DFtAVVWGJWiNgyLohfsXNVTSkbdJ449P/NoZP3vsLEccfey/1XPXBv+9RHZsE5bU
mvjC9YW1ItCYG1/n84VJT/dWyD6wlYZEU1gmHRZXuARQFTnBe2zVd6u/DW93AJCv
xH4btZcSihy1lujtkfG4l/QCnCNRxXUiai62UX4KpdPTDvZQOZBPDoj6tNZxltpy
FcOLFVMX2pRYCfgUVHlxp6zXUDBR3Bsqzq5WQ8bBqAn4mEHgSloImCPR2U7aYjUM
MLZl/tlkctXQyQxmOaXad/yn2PydXICzczbo6+wp8fD5V8jRKeFLPYMYabrDphSI
KTD0h+Ix8ecEecDEQQbCQddDNR2UbPjFhAfeK9bjZO0dP8LvsjGndEb/p7hCzGS2
SQsQ2j5BWVIKpZQBMBkdK6TD4C2a9QBUiEK0p0oUBQ5GeaaNynWP2UDnbch1w7/a
2aD3WCOSxxKu0I6qNryaHZfsokG89E64yALIepY2CGdcs6aEscqi5xzm18gZ58s/
OG9ZrmdxKOUVGcW07I5bcpyNnaniJr/gyQ7z1XGmc1hqEvdLtBVLEI/qVtKLN2sc
WF4AJ3PxR69mAwEFdZhq07mtdj2bTre9udjpxMn+MXwIyd4zOQXHp+cRQDa9l6lR
ih76Qj9msSf4upp0RWyt5SHK09v/BrpRDoFDkquLoJ6+g0C3m7Avq1GCBOxIJUnf
AUUbq7LQKjx4WCyOokNLhVtD//TKkHY/u45Ps3tiZM23Dz40adLVQ/R77csZ8PVP
vXQPbIpVFjylFvxfox/hrFNxrsJ9SJmL1g59M0Q/u0/jbP7zqTJQ0pBzLRB/8PWr
StzXQAzBV1OXFCGksBmrKocz9kSje/kxd/4jwnJKjfQHGOYMrEB7ZnLudlotJTGF
TVxP9+YTPc+owiorK5vm5dmlzgObwXLQV5vck0OEHSFUKXHyzn3kaq4+p2NrZpfI
Kd0e3Fa0cUBvkYHHkihkHaflQ8vtgnWiQqpNehs9idQvCTxsOCEg389WiUexbB5k
FsdBNhUJgEz9vXewN10ZGE5jyNrR9J6lsXQ1zOJOhbHadIQcU8SKE9pvQk4GpfSP
47Af1Q0KV3R0TPqjCgsdKjO7c5HuvMVOVvWzOb4x1lE4VEYFiKLIUU5oMQwkSDHf
hbJZkuSTqZHPunj8LA/uZ+DKBl2RScQo4j/BmKRpNMD0LKG62is6+roIMZGo5J/1
hSwbD/BvRyxiYS/mOaLjzx1MkQS1LAfH87mCzxoj/kjcIhOMPr/XLzzB6jn+pSBk
894MOpZEf3WoakpnvnNeO8zDCV53pu8K3UkdHXMJydhbPD7gwABLRXLhj/zrkUFe
dHA9dwuj+Uh3cPYDOBZZCWfNMdUNRcyam6RNTjHx+B+icCx6pBFwY4Gn5ZAhGTLa
VeRsf0uOlNBtR8clwP5DATjm9f5vHbtCZV865QaSsRCcNQ0QBiLnCCETfOJx/ZWW
`protect END_PROTECTED
