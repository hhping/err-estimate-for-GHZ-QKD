`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4sLbwiy8ngdVkSPkLgmF0+sJ14CL9n2UQnaCcbhrFZzU1Yti7HBHHNiZBuAdy4A5
tGzUCzyKlqFScfVEeoU3SffoKotw6ey7tKyfbrtF5eBPA/+/dxhcmHvkFDHsTOMx
m3fXK1iX0koQ/5b94PwKXfX5Dmwvb1bwTvuIzrVz3LQyc9y41vBcEdYYuLqrNyH0
a0cOPiMkqYAmMF6BWrM8woVnozC4L3r1QqzUfQ+qaUgc/wW3FgiveyBLubTX8Pwo
huPr0t3d+zqKV4/M3I1CCJ16jtzgGs840zBPIAS/fZqAn/JsVc6mCSapo5U/Sf9n
munKsDfz5UR0ZaIgma48vUWeYFt0yR4/TDpgqu0XXqfNrFxKbbs8KafA27Y64UQa
itN2fsSvX5/xPSPRq83wnF5fAXvOlZ0i3vFPA3cCxeYO6xfsNSSG6zfL62PMWhYt
1LYx3mWX2iY2YoigDJOtAtOsfx/kPPTVs2sjuWqbpbmRwxVnsY2Fr9SkwlS3WIjw
96u6fsQeZMWlfT6TlxsxZQNSFRAww6wxP19/jWrYzuukt76mGN6Q73OV577N/1wc
hSmWTTFu0oQXKLdQW7D7LiKmxT2D/IUvhrQfTEzO0bfyLZvyiwmmU2oGwnkHkEzB
x7eS60kMgKNj5I4nRXX1UqV2+0AaVON+eBJYn3IngkcEPnvzinJT3Zb7bPUmU6Dn
bINLQVKISusfWmKVFJvYxOOkXDC3VC/Ym39Wbalz8i1hNxOWnTCnpClec9ilKzbk
`protect END_PROTECTED
