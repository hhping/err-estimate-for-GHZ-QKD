`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M942EZGT/ffgO2oyxZxQRaLJCClTiJg4jVYRUNZ6M4Hmq2UqxgL3sKlnMAxhof2z
LcCNYuBvBfa1FkT+WbrQM5c//lvzmRqGh8P4ejAs0m8N90QkR4ppns0ve8qpskz7
qHVr6n/+4aDa4i9qBIVu4KkV6n/jxcHoegRlJ3IMEzDPLWfhEkz8nKg9pWVBxub9
DzR2HcyU6pC84b6RA7Uv8VAj1C2tJIt94lz64EzSyVS92dyeOQzNAxcxGaKH4jLv
sbNMne3eIJWetbdRjffOvoUU2WsOgsz+0h9FJpI3JFZP4QwvBq4w9tZFAjagVCBN
dh4FtNGPu5L5YeK+pCiVwA+1STASzE0Pj3oaNH/9cld0w8ucV9h/uSwOixaiZ+4T
DvWbc3NcTNjpJtkreQFC06Bf1+rPW/jTTjyXwRn6R/Nwq4YkkoDlAeJlVMRxQo/P
iL7sFjVKdv9mblkhOeWUHOXU5vKhkx9ybTQOpyQv1xfzsYoafScoTZu468hbfKIs
oG869pT4u3We2/RCValue8vbP7YQMddCOr5JIsYVagJY3RX6Rbw5BlHP3tTGVDHJ
CCMlqZorX6M5aC9w3Q6bNZegxEuQ0tCMg7iNfapNDl+N601Y0wBcz9bF+H+stzw8
+ICwFGvFR565D2amcxJhOshFLsEjFeWGOU3Jxqq6olw=
`protect END_PROTECTED
