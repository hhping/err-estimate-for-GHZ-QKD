`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d6dHsfPMUvdpAkUpkbQiEiIDF6wuBl+WAYuH/pNKRAVbx6n4o7p6j6IrOmyF5AVn
ofVV97oQJU1pFo6kclchD02+0Ij+yJoXybO6VNnnkgzHFsCYqZmJz0AonTwbYGmT
TTb2hQnnScBzxcCztt/lmLUYIUmBEzGlTSyqIDQVP0ZTmPTTdMHZGXttNBWVir3i
SmPs5nfeEWJMRqYnddkTTKUwty6+Pfy/lAqlasnZBVwp0G6vuvoc2egwfOKzkHie
xDcLb3nDMmatgAQNt9Bm35pzNth/5GCwlVDsntupnPo/PYEeV2KfCaqn/pHdluFF
yrAgPrORdfgN2ksv37QjZlz4v+ZEBE3+EmlyYiezOmw+Ap3Ap8abIEZ9DnfcjeL1
Xq3GtzG6HVzcemxS1Y1WkavkINj5xZ6QbyUxnNi7Qs/3z4itgiRWVPfAGhiP0M5p
mJvUn+1ZQHJjT0w58F056h2GgfBUf6r2YnjmNvy+HFlRfQ9OSPXqESc4qtiz7Db5
jHfQ41tKgLoiYced/kzziryB0eMKuRDVCaDLDPuxn+hAIMnOaJ0jNgKUoXZJfEr7
VjpG/so5YBOr6gp0/OiOWDyKV3YqBOWJgUG5ADIJZduKVvaut0eQvnDhSDC2DNh1
PqS4SaBBNoE6MyLXYPc/XT3UOIsFWE0iT0JFxgzKrSe8o2M+1oxyyoNtt1USniqP
RsHGoPu1a6WMChGaf58MN4ek5hDOZ+aRS0v0/zDcDrnynI4pReKIwKfdnZ0/KWpf
euGXlGhZgYeWiIOAt6iueDZgca1NJ5VaGMOPQuEmzNcmwFvIhIupqYAqVJ9DC1eH
Jve7p6MkxZlZAqUVwSPzqBADGC4byAAIq7nizvqETNCK03sJb329zUv77NPQUBnu
oslKmSLk9JIjAPGdfuzIFhA7pJPplszcdWJblGLbGRJc4ZpXxe32701o64etxIkq
wWpWrsDNbhmzEzp8Wk3fI1yvFqUpBpdwFtYNIeReIt0oZNWt1cXnGmAAAx4sQjoV
8gmNFB7f96Z4cqa5BUksCQcVrsefBs/Z/DL4lYezMYICn1o4Ba7SecVZnozT9G7y
Sqo/pO5o8zbJMCMKXP8a9UctcyqdiAoiWgFcao4RFvn6XH0DSJtfX+3keCwwS6sn
yQqZbfUi84tyWhmbwWfFn/zmEijhe0BS9HP1oiyc9KVy4phTjmFGAp1XXFfK3Hn4
5uy8dJL+TJkoWnRoNt4Yo9kVsv7HS/LZDPU5lo2eh1XkDng8D8lgJgHljte2KRth
UPZ8DHUGzXSAw89SG6/Veryng/olIPc3wWcYc9PRvpzjyVeIEZX+21GI/xoWLfsM
tx1d2Z/GN5JP9fjbNGEKIs8a+sS2zotDG2l8PaOZedEfP9bYauSks4AuJprtb8KR
GiP7l6a+GcPJqnnd/HC9/rMMxMz6YG3UwLEnwQ1pMpBgiTGXJ3c7sSJWKu93In+0
izoO0z6Sut5KMdgLHtO81fqUXdoxb1j0okb2UWa5g8mwS4Ie/XBoG1bufitszu3l
CwqE7b/TJv0JiILbNVSMJfxx1d5tnt2RJGrdNbDxLUMsrLS2+h/eRCg0nBPCwDZI
`protect END_PROTECTED
