`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZjQ6uKZURSHheuvZn4Y0m+MpvGE62RMyzME5lbowFluufZaMx58q6OcZHUQY62Zr
RgqOCN6VEFWRZqTtDqM2LfmPCMiMsLCgqchoAPlN09onrzcj61V2KfbvqJhGUoln
NKcs6UqxSZuLeEa89axaqzwtgETjQa1ERtHyIussfmC2679WQROwdJaUjMGv6MMU
/ZA57FAdPLrgBBIfN0zlOai+ReozFcw32VbxQDTr/lmM2nyKemZG5nlFZC6w7Gqk
JXSiE3DpMHflrrd08MrjXKiRDqvrBm4mTWNlrSwKlR+ZbwZtsVNd3DRyfiY8b4CK
7RaHXfPBO47NgedbVCk9Vvj5qO90XQtUoqNcq5xKXmsMK2w/n+ahVh8h5uK01wal
1MSHKY1BwA67A3J9lJtMcbtKaJAm0/5O6ql6n+ryNZlbpo8Smnor+qTHMb4gDRQ0
P8xy9/8MnQ3akHyWHZPJ31FJ4fPPRqGVuUlQH5gyvyMhFGxNM43xkoHY9ZBxU1eZ
Aqx208loq7plrmdINRtUOOd8riUPuYTmKwI95nhLcmx3DSERSsbfhjFU46CZia8a
HXuF6RwYyzkFUzsfZD9gS2FFftgOAp3albApbSHWlTLmIWvHyraTRGCsiuljsJ8M
OyKvNFlBAzOaKpgjExyjG6cj7jTT4gvzx6cXma8nWTRsa3vGlsPm4rZnudx1ZqeT
zl6b1HNFh2zm3FgFjYBify2ec6IQGRKzcv7ehQ9eXMVulpz483+uUWJcXRTobqxf
aNUOCft7QEyzCtcqV8BGEE3SLjIMxdXdJ2y8xp1NLH2HbbcCkGr7kTaBhJe9Sppo
6ROGVlIP92L1YOe1PV+GixCEMYSmNlORPJryVZz5fe3kYEkjLHZOowQqn40c7Fib
z4swQBWWMw9e3n7YZ+NDu5dNjNiKa9Ak9KPQlVRO4ptXmXRxcdVp3HHpXsOFvY/j
KV0DSsGgcMOZiu0ASdfk2znq/UtQrSz8F2dcOhomOGHbTcGJg8xfI5iPM2yKVRiw
jJyoJEzDMbCyGhM7FDJU3vc7cr/FD4AAxH0uh0dN7s33ZpklPw+HSiNfRR7dNob2
oJ5f9wPGdJwYcF/o6tPPoNevV+2aLHguF+cRpjGl+fza/JsFLcLZZmjyHHyOWxWL
aaT4aXPyJn66TuAGMRfcADLckRiMROrsv+yDlWZqSEbi4WwYV9NQax+ovxMIKesC
SUH7DHNFee5+TCuesvW480FMaCrET7ZN3C4ZZtRBCzB8SDNq2c2+hXEx4jdSPNoc
GdFomy+5pPPAeKgoj2W/H8bMkzI3KAdKIpGWuiYv4HmO97GLCMYeC5lkizqjvIUu
MLp+nEcmurWFLH/yntnEys1B0y6cgNBFgxFblLxr0DKRnMzUoNibDnjgF7wROegl
3L1LFW+M0IXOz+u8Ufr+cwKRO6WbcICjNg7kqsUO2Z2yL9+SnST1dzSu79CDoXEn
Wu/cfdPhOVkGeCmSMfaphl9KZEdSLH6C13Xh5mQycUA4SEJYOJe26PMYSPoIspQa
Beo+e03Sg0SfE0kdHRQpCweZGxe5IDtpezpZxIck3LFiHReFWPeFwMZfcxv9BGlg
eyv/oS6T650aFfv3SteWrr402su9QIGnqa6LS8ELfRdiHyjMdQqEMw9qESNbtOBU
`protect END_PROTECTED
