`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
le5ZfAddCGOFrqYGs2fh8CUQGIpLG5W1rsc/Yqo3RHYn/QqSxP3SGHydJy/BNedK
wdCV/FJL/nLVmvCkAHIUTgW2DW9qeZyTDyNOkOr7GkeuM0P5mQyIcdVipcBQJ35f
cTJnPQo7vDEC+MpVl5xOYp/yr495UhhLM0QiaRE6+0P6jnxjxm8MUCsbOJDQWI0T
3GnD5YbxZP6DHGrPyiltPJAVzCH3+xpYNlx68KIXjKC8MSOcUWiGdFOHo7s+KXrM
Lgc5cR4onEDjOSlZTFicx3ttK2aQGSd/j/iwV92bWOJkf7+8EGQA8WYSvQ0ThDSB
sF9xvNY0QRpTGPypPF89MxavZreQEOlE+kuQxQobqyU6SG0Fw38C7VzlZ6x8iS72
6IMME9hu/tTUS3VNNsP1SbgrvWVfkpofme1R7etGT3gNoh9NOz32/DBIgr2WvK3a
fOL/KE+C/bIeXE1UuJvkJdZsaF/LK+7+rHyxNrhCRL9bFux4zazVrqMZzLtx+BgT
GZ34vLWkmlV8AV3gsJdPYSWEjn59Jhlu5Fh5pk9okYo5J55wRYNKtMrADgRUmBn3
nVKFK2CVxdCQt5R3rYTm8IkJvrb/x7IppSilmNwnd929aNFubxxxNeBR9kQHk2UX
VcVybDJcer0wNmGRvLzZCn8Iwgj7ZP5fAK0BSlloV2Yd5f+XVBbU8NcMLWdCB/4M
GNxgaNL/OxtjMF5ttoVQutPBFYmQUQCAMwBkHVO5ixoBT5MYgDCx6svTqhfSxZFk
kp+TFfjOJwGwLK3xfMJHhuY/QjF3JLhF/IMdiDaM/4lEraPljcP/cT4pgEWol/JR
G09QTmI1Jj7z156hASDYaolNUB3Eg5pcshYnCKRexBfRiw2t2tPRuZuQGBa/O9Bg
myjGsdjGh502Gc05vLrrP63CrlnIb2z0NbTr190e2l9kWJjUpYS6mm/zKH/PKjWJ
E6Wt/AgVDmrnqlVZcCMKt1OmKOSFkrXLKYwZJ0PSoQeHUUPVvCfmd4XwqxFZA2YU
5AJXrUxcgB7sWcIdQIIHI7xnYmTMKjO3WYJXP+DiHwqrO90eZA0OYOa8ZHyYq47+
rSIQIk5aEwXAPLviKAKx1FZ9//WRlOBXwN9VfM8kATD+rd8V7BF/37SCSIu4I9KM
V0rLo/d89VVDkXk+Y+q7hVvCJV6pkujTX/fpFz1iDsNlDAeOb11+ZD1e2ZAMUYiw
TzpznQP52VeWFXxbJmF1lspKOch3jRZhCEttbfuWGEcNTAcLwSF+TaYeqQt8KiMb
+quwtNyJKF2xJPoyxGuXskcOiShuXAHxDnrUEPYO0u7jrxOrGkL+UJLVRBhrDbAG
loSMRM1/Ep8yFpcSq517ho1PVFgKG8hjryh1oxAK/TAADuXMG1Jzo9B6AwZh/Brp
jEmjqsbASZCxvpTvvMxQa2AzS5dYFGYXqJVvTo5d2ri7j6JP+MHtVj5bhoEKgyhf
T1y2pHJcTqZM6Tp+Lax+2wdwVeBhbae2UBXCXyEaHVao95V7RnFCm6xfJtDeN7t/
8RgwnBGPSwENRFQtCDyFy0zmo7DZsAAXCPyeA1Bo3VlGqwA14CDwgH5zQc7sacsd
PPkKVCzmgnQDjtfE1IAfSg3jwiEfkepzSXuft9S/SEg3cViZNfnqq1JnRuM2MFwB
nWvOs1f+qS0jmzrcC/HlqE1QGIcxX2V3rbCq/DvTItVcK/5CN3WoLI+x1q0ybSfn
1yv8zScqaZOQo7Ya7zHyErNmH9mCAzQDMVOOmU6tigp2F9PCPsogtaBmVWGqqliV
DLVbY1m1NKAXupEhqhojwJzQ9lNu6s2UkENMWkAP2w/aa7id6ruF+Rk0Phg/zfSi
PV8Ru+aYwHI0D0RLh9WjJuZm4HlukHI3KbwN3wOtqMq/xGQaAOihEsSkP7/jTTfR
Irj5LbxVtccd6kJjmsNb6bdyfUoUrP/UPmmrszdE6tGIkcMtVNkPe1Im0uBHSKyR
sVaIIJWAC4MVwJ7ABk2Z9sf1xHLC1iqxepoRI3LEe8onw1FjCEadpgQrCbdsgQls
crrXbNvHaU2WbleGn02JWiHoPcuXiGrwACJKulPwQZWiP69P9DmXXNBIQnkzoemQ
FUh8OdPlzrKYgJsBmZ3HDszvqCH2BRjGy2ojRRq1fCkVo8Cz5c/feAIazYEj74Lg
4Y7iIA1mzH7u3xPHY/LKk25z1PwUQ35XO1QFdpmpoujHYYLVdHcc2HLz89u47mcr
JCBY9F09dtXJoq/MnWPrBQfBsbHIAAFgIi802zUjsOw2nijeZ3FL1XWQ8LUer5Vu
EweMWAI/6P0EZC8gGOY3QJK3SUQC5Qb//kcfkpSGlJg/GJmqBXFmoLv6y0yo1sAF
Ur0FwlciUZlSBAYLEdzy2Dw3hrDvYT/2Shn+Ea2OiV9vaE9QPMobqhekOw8Uj2aE
hbwukBZEkCzsd9cbm7izOueaG8yRhsTKQ8Q1DAGtg0WJ2QiubAGiKWhiYzjLTrTN
IriDCD2QtTLYX9+SNDACzHcT7p0fcmyhOdxKzmwFWE1yQ9r2SDS9vsK+az5pRKcB
Ow+HzHABfqtH6uXCBJnuuC/pj5gTG9+30CwaOetHi7LF5mQEGajY/piOpJ8Oq667
14IV1q2fleBKTzr6C16yZbwnlcVkXY7LSPMMf05b2NVXBLkt0QkVe38stuB/eI/I
Plb7oothyKbri3AV1uHVlzTvddrHWifsmSsZjE3KdXazvxfpzrDXcaMzNEWt979J
FXa2BmrJ62U7n5+S5kEI+6zfG6UhGqz9GuiRyHhMS0sFUtFl1ViY1uxJ6p+S0Ta5
iCyIskyVBFsZDzXDJuN7+SpCH73xJSkEo8oJijVjbDB6lxXtMw9jLFMc6Nj3zWKU
1MTbcDeiiy63SS65cVPzeg8AgH64Za7qbR4pxYUjb/4/aRNLEubVFnyf5xef5X6o
glCS5Cs4BWEYutlIJKToxGrkf7f9FmCADCzlw5viIdA3FPVTP1mWnZWO1tSokcbL
qdtqELTSn9BT2DOOTFE1goZEBtFfVNdjo76HfvVw4ZWEL1ZIBrlNAAlHEni6DJR2
awLrh+IBnh21DH1WgQ7KFcTYGIGUYIq5HFL9182Cv/ilFUKKEkQzlocxN+XkFGau
VKbdLocffYq3bZjjLNYbYJrAcrGS/pgFcd1KEa/4IGzLX010MVJgLvIAHHNvTEWF
Z8GmpNAlauKYbVkm3uUsHjmw2F1xEM0QBg8XNQUUdFMkQODD0Sr1CGxjwyuwl6oX
gXS+lhpoVFjnE9A2UqozCA1MMqZSsu0ZAQLO46Wj9738iB6acMo00JDQbttzalG0
Fdy9oqCjx8TTQzOkYO2wAdltryAIqFSQKZKP2D1tlQwKkAZUGtfgrGtlGL161k1q
mZAE7P30k6C+j3RVMYWDSJjwawB7EFh+6qxwycWrApiHzOuFz60U5hfsDvAKVxsZ
Uk8ePcV3W1inZUWK+wbD6Gc6WamPWatwF9M9y5TSWHCCGkzfa3y7ZwhtRCmpIZRO
aqZXFtWRXUQdIdp74fFmbC7W9P30HjxBr3mCcy5oaUWMNfw/H3ZmLpF799cign3a
msVM/1T+v+Cx/ZMzVyTdAGJBMBFeu11AGQ8qacISXJBHQAZPdfn/BLN2RLVw1nXc
ZKUoX1y1NtUXXs+ZuDqxD3fq9lzoeU9MYBJ/v72IYcqw0uPqdPJTPqREB8+NHlZ7
Tle+joqequI5ERfsU+bDBN1CVTbjRMkEwbXrt5GwFKXNNAk87h8A3X1eUaCm4EAf
9j4iHXi6D2pQCGX2AelzeR7bopIwRZN2VuvfaVcyOhd/21o12E3Qt+/tIgfwzbMI
K9oAlY7SPwkxqQmueNYFDSu9VMSqf9+0Ch5F81pMc2DmGtF5sJOiRZsFC53Zda7B
vOBFwP2B2ADxDu5ATbUUA4QqBZjiY+p5qp6ihgU8iYy9R58bxq8wlbrGE4kUvbGM
VG/kMQocLlsYhtFKZQpqQwdZhcwL2DQkbd9ZH9OYzaEtxN6Lir46bctj6XDUXLeb
kD0KjuXmvFPzIfK//aTtZG4UjhA81PMfF68HBPIzgwLgcnpDxkaYEfUHDSTWLtTc
CTg1fGa/evVhRivt5jcX6sBWWNONbrz+LqGexOdDjHvQamRB8fu3OhvjDQsGOVSX
8iEdNAWkifpxdbQicOHBC2shAQMDeEWLsPIWushHB51WEgDpnJkReagUlm2VlPRE
OIrmcZDjHD8bWiGrIWaE7BYQuEFABZ7GDX9dP6arBhc6o5YRZ8L3O7sTYAMxl7bw
jM8Vej7SJVCC9cAbjnKXnjvN99Cbq1KkQWohyK/A8rpjHtiKDGI5o6QAmSVwekA4
pHKN0r35E3U82YjY3nJ5oqQN3cEPlq9mFyoPZ4LufgIMD99Ap8xvElkGfTExhqje
Z8tgX4Pi7wolENGZupQ1owdMVf3Ud6tq4Nuy7sHF7D5xQ4LQfjs2RjeIV1QTfWqo
2MCWQ9Xz1IncYBiGgQFqPqWLckUDtzHU1KOQigh5Xs16Gvv+U0TtrXCiHfQmmfWd
BlBNSMLGw9X8HuVLlGycTy1a9pAGsMrPx0I7Pyt3ZPXGiXK2GAyTt41RTpzKEA1q
xZ5kdlA+M6SujoDsw1CCKJ9cIMyRRI5YQZr0eEn1R/wcSkDp5nSPXvgM306dXLSC
09eStVgFMRB2OIp5fdNrIV9n7qi42DCls55KScmEd/ENaWI0Ur8bhuTmGPpKTe1C
42Jlu/2u9k64mhFxsDUCwtoHKr1+ZJO1W8oUh2MDhr80VWZ748Eio2dJw1evlPrc
y2wMHJt2layDiO9UqViZkq/YLhdN8tVoBAw+roDsrBMPemwNW6CVOnbSGFAiHuHI
KxPaSYQtFn+Q9zKabe0XIZHqcKlDuxSUu4iN7ZL9sXM3fnDYv2A+IZSRu1KELXeJ
5Ie1ARXnwcXrsQrqlF2KCs1iR29DPhpIShlGDbtCUvXAdzECXoXBKl53gu6/puKJ
hFSWEeNKEGGBbuaW32M8mqlG+aGhndJFlbklpdwooADYcN9nVyAf+qw6Rw/hob02
ipbafKfjB21hF0a6GVZMX6oRXwHk8grY2dZWW1R7SObUymTwHKs3lNAv4v0DwHg1
Uy7yqIo8tinZSnhkOhfnt0aQ02nWXIU968cZd1YWoeWZ6gDlXVnG4SGZ/g46cclo
HiHxnfuAbXzDdEWHXpj1GJWgsEOiKxXvEd15zG5YJpNDcGUqRyaTMK88apBgwXZg
eqPDwlkpS1a+SY5kxjV1RlorVt2t7E6XK0RE4MUIM9i8EifjQc98ui+LKxzkS21k
X2XA7KfR/WJ54ur2a+TKvb0QjbZ0smDwFbyvNbrkEqc1OXRdkHYGLoOfLa2y0dXN
wvRmYhmjPmlSopIR1lOM6bastFfugin9wBtrs0cDW27RkLY9kVESzCVj0+27m0Ln
4UH7I5iAXmDisYUawdv0/8ZLrZgCeRZJmiPBsuT5fID2THzMh5kgtOPxl5KGzXQ8
G4ts330OF9tJ9/08cj5IAEroIBDXmgqbi0FXHWRYc0ba7RcIpf9Ajb0+/PyVqKxG
AEvGL0KiqD0nlYJTYmyb5D99jkdXQFhA078hv0BZW0eqxb5mLY2eK0yTikxvtZxO
NGaKBPwxTR4R5tzL0J0C59E1oonktD7BzLWTXC48PucyM9l/g1wt0+J4YoYwkkwr
0y4lW4YOmeUYs1CFlr01ZJGYQ1nVoy5xN2PtZekUOjwYixRTgmb+se9mnRgfme9X
fO6DvFJXouMov9/68Pu+INg8yfCxOVdE05PIyPHvcoDhYuDGpdEC8QFxKHIZrIn2
BXFA91bNHGPdmVsi+Jsv9/U23t9e4rd3KFurhp+3qK9SdwSjznc0EwbXvn77xtfi
NpuaDuCiFvubpRzoF1w/ipset6s9iXk1idP6EPup8OgXzSFTqpiqq7o4vB6KW4vv
EzGWHAeOWWWB1ZUQGZv9PA==
`protect END_PROTECTED
