`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5DHd6utbiBhbQn1fJ+BSdTWlKh6dGF8sMcf/BKaT87r31xZWBDjR9gWr/phSGVty
ahjIulJHyJ8oyAN4ZlOEhEaL2BwTv2hIoFzcbFDZa1ritddbkRvwoDOnjxeWglZ0
+y+Kv72+Zp/DtJj+yRX/QI0TOvE1qg5LMPZdTrlfUnp6yUI35tKaw8OmWsyZYqtZ
BjRYaUYh+dt4HERMpKRhD6JFbWTHVu47NthJ2btENKqtQHKfgw9upucNAvokDurJ
2TrZI1d+1JZXBMnLnJUP9X+C/tym5JTofMVsKXOqV/ceHDKWZIjxTkhN6dDbHF5e
E3NbMxGO7kjpoJyPBYdUw9tNQx8pCk8aTBtrJ/VGB+mzvicA5l4ulKKQBumz6AS6
ljJ8oXyx1zYeDsyHNPqZirOFXp5HvI+eYLFEKeJ342xCguIOY4Fsxspmh9EQ1Y4p
/Tryv/H+1w9UAzoTTLNdf5GiHx4Zpik36BV4wSH61YkDBz/5L4+2ItvSTlDqPfoH
qtf3BjudVJ95wy2YDe/wf+o2QWaoxBZ5WONEuFMQ+sKNM5P4LAkvjcWLt3oTc3Go
gW3hWAwndN3oaLET1h0WWnfHSoy2NUvf0tG2VyDA0J4CobnBaC9kmEJRoWD0Y4n5
YYHCUcBs3K2UG1GZFhZguWkWwBp1DpO/vkjvGZeRGG2plX0lTsCGNrcn591+iufM
Zyin1JqtPcbkgGwZOW11+Ih0voMYIzPDIZ4YPnRDtNUuaHWV5PIm9KyINAooTgWa
OVaLJn6qlg8gKDrW81Nl8WwXPmP32NSvaC+r7TND2aiYr9fX/P1CLkblamtlfrhE
4vSVW1J6mMiogeuMnuui8Xy3I1ladQ1jz8Ct66OnI+rMNL+qFjn9XC6w+JV00XSp
gCXZCpaJkw9GSSGz+rlFr02cf2yNic+idkwBbNbz0TY2pAgJjQRgrJ3WXMjoxFu7
J3cJ4/WkBZncKU1jfapLpA0Ilywi+5OgwabC3gU2vcLxwpSUI2wONiSf6TDspcvL
8HKsaUyGUaI/Tby84nzcbwBOSD/WSpuBI5bCymDaeQ9/eeysd6Ebc+hnHTDOSoeA
bsMU9Jkbg064s6S30V7WWi2HHokK1q56YxIBVvkuy3cr0WlVJXrjlL2z/HMZJ6JU
aBh6SCNg6nn+CmWsdUbNEea+wtCp2E9DmCRnmCxKmJbP5rnyEiZZc6XWOQoPEeUq
9NN0Ra22lUeQpjjUUZRFfpC/EzDCrWbU+DyG1ArDnGvHesQrjAbrNGjM+89HR2Hv
CT7JU3nIj1Rn9aSkA3NEq1SdgIbmX/K3n0ByjnPZ4WXVAaZefyJxBBr+UUItgIZQ
wRXpiGNvakKuoAGk1j8AkiNqoQc4WtGJCLBlM2ZbJpzQEOv52U50+WA9SZ57g6Y5
BofDUmZ9nATIiqRYUOnhT4MF+TwQ/GZIljBuDwLD4pUL7k0tx9cThYpabE9l+Cuc
1SrMPHXXhuRbB4cH1SmTXAzQl5lBcjlnJcxA3VrTc6hf0a4PAaz2nwNJ7pwPaxo2
eGeYaqt9YuSwzyLBylt9dMyJ+xQFfnI2I4C+bCmbzfe+EMREEQrMBT5L52s0mKBl
cT9RomY74wCHJL3DZkt/wCSTFjar/Mk3ER/LKpd7bKIwSuxSstvr/AB7d1YPnYVE
LNLBaBqD4H5qKhKbYvrUJwoT+gfLnY+8BO4IT+3s/x+eAbKaOqkA7ZZVgSDnq2Or
6A10VQyb59aC1fnJvb1Ql81ls2OdpLu/V2/piba+m1f/P5651UlGNUir6Ffq/kNi
e73tzdMmCUvPHlPJmxgee1WWURz10B+edZIFPeRIaazFziHeYsl4isw/zqfp0TPl
YhoARXJyjWuKEF8AcMmR2bSbY/pvavLrX7MXZX7xGNFUDqrcZa7dhwxv2yhWrKTr
rxrqkGCKxeywsSVKv5wxXWQbtqUibrcwTwpKV0EMcErLYNDAu/uBbVBXSyNTKb0j
zdn+NIG6THyf2G7V6TTEPMW6NTJ4cAJK0aCPEYzxtLfrgJoHr9ko69y/vGJd6Vnu
4H0IPhu5UDMHCjkg4/8POdkbl0mmtELLB1sLV38K3LaKsMivtTA/ulJ8iobZv0d0
LESqU5KjORNm8nk11LJur/ehIFZrsJyGSBNAmkaJ+fRC4CvX7faYmnHk45yNFiY6
Lu/EJs51sZWjCqa0NE13HotmBQ5qOMnXPqUrVGC4jmgmRR9+i0jHuEPTmwh8cPeZ
9CfwXdhRTVEyAIL3j7gxf3aL0d97O0kZjAv6Tqe56gERg94ugXRAUjortTyZ7JvJ
P6wwW9+PKkx2CnP0GY4OB1Wv8wSA8+OY/GTxVUXWHVrSjbtspJffmoEhfHqaIkkL
+XvtKQatXafWX8ye4kYibV6lIO/ZBAAlWiz2A5ZwcG0vK/4OCmmFbJXfFIEGUOjV
b8pQHXkBnV44EWod6SHPKdrUEr2uoirRukYLYPbC+wu3Iv7oS/+z/ZHp+4PUilTN
Q7JKnUGe0EP0VdofX8b6IPtcf/3Jjg4Bw92thFTnZyo5tkF5bFOzERvQMPVLfKVe
Ot+qC/f98UAsv8CMqXhMqW9OEqVlL82B/i/7T4gxilxXLL2X5wSa13LHLwAeclmP
I2/GzU6wUJEvaFx42Wvve60ANhk8xbxbAa+wWYUmO97xrWCm5Kxh42yBW7T7tH9N
F+yPbWIM6KFyvPJBa74p/v+zoBhVMq8P0FfQUPxzJgKz7U0EwrU8f5wU6yBYQpBt
Pcs3uxqN7kxqHHzffsIKsp252uUpy8ZMJCHocz3SSGbbvGjifxHqrh1h0gPBg7m5
xyezcbMl9e2Wcrua9jv0iKruyQq55IKAESB9b4Q0znIS2oO+CZNe/RUxtGaAJaZ9
cMkbYkjA/Kxr1Y4V8323Bkt55bGcSSyl8Bxba5teuv4=
`protect END_PROTECTED
