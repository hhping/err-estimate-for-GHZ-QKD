`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0OI5Mv6fwgMfhMTKzGsuz7sP2JGgKUF1sVwTK8KLxFDoulKTWu5YR40y3QBslSj+
mK41Oou2HkMhmZtBwjfsgERWAQhMZ3gy6crFcIace067KHfUW1Y/y8EniZhS7xnP
miqtaAapFxeTtNK/pNFV0QBPpMy4PfE8If98ZJOFXZQVPVYNKkvqdBmJD4TgHL2r
MLlTa286XipcyvF69SD/BD3ze53bmZezC20ZzJN10enKPezvCnCOrQjTWqWXPgUt
qGuteh0X/ByhMjvWKcDjMTdj1IwxHATTCqW7lDLJ9A6BEPGtlO+zPy0MAAbfiW1V
DasSwimplGZVC4OCTh/uswqZavdqmDcZ7wtF7cIQjqskke/fUB+gHPX0/7PYTjoL
uTZOYxJD0dzdEx24UJJbbW+OMeUtsGN366UyXZBUn78ar6TSAXrp/1ZCr+M7xD/O
JWXDLDI62/0M+f1MF/Y6oTaYVwHeH7rQRbGCfyFGk7Jv/AWRsDqlxq/6ew2ENETH
M/WoZ/iGxGd0FX4dwHlKXSpheiTMg3BcSveu86RdcmRDWT/yjKNQwDvdMiwz3Ulr
qmUDCXVvHSpeEuSo8/hz/Sle6gtpju6ieDllN1QRZd1PviBlYFwk5hDzd0mB0/t/
HeF9SmroCzyOpO+qzW7QeYL+/rX9X1DxYQQwerH3CeY0r3YplEeuN9/++1Y5FC3G
KIpSGH9SvMZhiak4tVm/D+ahW0c60b3ilqe2hUstCwZypbvS0fiueN1WNGAz5G/E
QRWNitUUmkyW9UUuucnxcn0B+PQ96x3aErBG1whLPS79UeLFmYf8bF1v5f9UWRgw
uwnO5+3pgC2tj9KmmvJXld/FVDzGLPF1VVJUEu7aZ1tPWdYwccqc+9turagK6qSX
LYR4GQv+b8qyf3DOpxSqMJBDm10g7Kd4C9JjqlLf3LYD3rqPUPo0JDeLXNvW70u4
vfpvQ+6oxyDLGTV6QHKFgktV9YNDInC+wborYinOUo9GRVNnPb8jmmVLQqgzwrJP
NB6ytLmjdDZU0oeqWbWNoILqkFUF1n8Lmmyngm+TjTwXceXb8vaRBL5E5TdUj+FD
G+oxCeX8/Y4iXy1QKqrG1IBojAR5g/qebodvNDt/t1duy26BWoOj1aqpvEtWCGC6
b+NOVV0QD3ziuBRMnt5uJQOhjXl98L6avGEBrtXuy+bmapVCMs+EYb9BKmSbYk/w
RaC20/LywEKWFJiZkZgFD7i9zftT5N95Ndl9QIQkZGBhsdKY64QBO2/BRdLGLPPY
sN7VkeHGdJCvM4GFGswfhxAS26s6gtEJUCfLQm9ykPvdvACNXeQg/nFBMORnxVxl
PypM+xpqi1K/MYENUDY4Aoep05pQyaP0yP/PTIh7weqcfdb6t9RJNsBaz0vPrV6i
PJQAoia//e5DV+9/8YGZGNtuvPk3HYZqPOPkn8k8j3PhRNczjdeNsU5W4z38hajd
lj68+FJt8XaXC5STJjaPhdny6ZLlZTHjOoNC4FWvzA6Q1UpYfHqL5UWYGExXMmpY
cAybEaaGA5pAc7OW9Ez1b+rogcSxASrvLcFrfrb+0tQAsZVjKpPOQOS7H4wsIxKD
ryRFSvKZs8TiqecI21hDLuWzHPtisB1fYfIdqYR7lvAnbjg2dTuB58d6FauNCnUE
EgwRXK1LOF2Cy66K6cwxTAa1OPUaG5sm10dQucYrkJgc6VutELGzAmOJUD2+pCqt
+mwrXBhPH7Ue/LHZmwRAWuDPcIEsyLYcqAEY6g57izyW7Cj0hlhEIWo2uDTIw7fs
yIcnwGKAld8sMC4VbbTNrDNlPWCAae6cc21odxIrn7OnRRXTytcGCNSjAPCag3YZ
JOAkr6FOx8iLI/LUhdDLBo0IiKt1IGPSYAD3d+jfCxF7XVGMGtygGPFDUZmTStqn
4kwkk+Rpxdaf9iAC7lRAUU8SXpmekOcsF/PvXFhpRr5Z2gz3n+RpAiYmXh+oy1Ve
aMeZwwPXZTHxPzRn6SPxvC71S5hDqaxU+CkwQ/lyodTVP0sGhKb6mnKFg6PceukC
kYiuhc90xKigNSU2BfE9ZUx52Bp8skRZkgfIohVynm+h4UUuokvt+Cfl5+2IPxiG
3mR7HZur6xGl2Ru7/rqEUop3M0A+VX6/2Vr2j/VMKQPtYCgqGbHpzKskCv9Rt8my
cvF/aeWrOdtWhq55RfYykeGJN54wLF+Vjv0S9HedZmc2QaADwOPu0OjvxWmwTUYn
SHAcTyhbR6RbFgh1GM0vqrIPhjFCByT9sKKH/FsuOqGJcd/vFBm+Hhes6PbvpXEv
qTSgtos7lFJedX7xxUJAIsEANMCyDFRpdsZInJZcj7RuiOAebTDjyuJxrwgHpIq+
DwVl2xNWM2aJ1ZYswjKZWMEVbIYanNdN6YCL6Jb5HMGIihMz0CbVReCJE3XTCSyN
YehdRegcSE9ZrR6I9LSDyO5IcVhS9BoHBDit+TEl2uB+af6hiWexKjQnvZQ6XPeh
2xHaEmGgz/SuWsO2HE+1yYPJ8LH4bMz4hkTgGpIH7MEU9Zl6opiutabcJJQMkeLk
Osrc9PTv56giy8q5OBq/oKS4YkzEIYRLlolmdivtmMPba0LWkDtit0opsA9kclfH
lg7pj00d7+yyfxMVU4/Hil7wtfaIWiZHB39w5AV2WkW+LilgiR+FDCBIx+GbeiWL
WISwdKbOviRRgkQqPhcS7lKiyrmoeusDXOjq83x8CFJ/T9U9nr7rjY67RU7zfcrF
eZWwJTWOXu2vIKZY3Ax2vL51WdfITL7rqpKX4eBOeXmcPTW9swBPi3K6DohPAii6
oYzI6pObbpTnDQUpoP5X7hL43DvmS2lQmQx9PIXqwj+0gfN6DzAj5ERSSQCwq8Pq
oDGnitfO0kq3k+O7BzLCJbsdb9tWFrsU7cNLc7oSue72NHo+YyD4UL8oA9vAJ8/5
Mb+kioH1S3I74IsO0TnBih3FV0ZAVOMtjkcBhV/nhRxkiIVRZdlm3YMpVJ1Q+zJp
4TLPjIkbN1q6wmbI6reKds4Z8Cp44OaSWRz821GfR49ev8mdk0kc37j53o7LqXl8
UykpnWcWBZfdFenTsFPfW+7Cyq6EqPxferbQYIIH40lBvD61+RP+07aRMjYBdP80
JKhnvC8OEHoEkCLUqrKo2Pw+PmSVI5TPvVa0K5Xe2+rMUR/AknvHjepDmwbVY3ip
K3iYS3TALEVJT9YAhCebbWWepHiocMiRQrwD9UuZRffljibd0si8S46LRkhDFiT5
uSb4m5OWNKbgY9CFkAkb0eiEqDjm9EK5RamgCfDYpfhZhnI5EaxmwI2RbxAzPWf+
Jb4ATe15UC7Bj+kXNxY7JNtN5h0MrhrMgGhzSnTJDMiH1UN7WR+1HCY4WX6Mp6+d
fGsLwwSY7mcyA7XZ2TJLV6FhbFDALgnaRmEREJt7GYtewD6MfgKYPdV8dVnhuhk9
5HhMgmTC2WoMdEwi0lDp+dthDCzyrz3ZzZw3bvvOKEEVeTptuMMtXapMMtXnSgGm
R/zaJJuuXHW4+g9yRcOg6QPdHM7xn6HqbTUbZatwXxowLdBFbJcMUguXgeA7BML4
1YHVFk+0+Yx/QJ3OrnMLrxMf6Pxgz3/xcJh+NudPJGKCqdBGFiBP+DJJncCwRGLX
yuJs2BsI7aIqiV/ZDT4+ogilnMYEc5kIHoH/FFvezGxWO2sG0M3x0mS70td5Dwvf
CgDmC0SaVa0OXtgBfZiAguCAs8GXPIQlmVFNXK0p8ubHfuzUtHq/UL/NlYKVW4Kq
zCCfKsyfdl3FbWDEPat5sDYolsufU7WwMGRTNp/gR4xhf1xNrUPDzkZjg7cRxx8m
C0Vn3+OAwyoG2FjkCzakHpJZcuKXvnIFZPh1OnCO7UIKCoWW9TeqpxrO7fpZ1qwQ
JGMA/eB0ssjKigsu6NrwiNOBxpR01zaAB4/dAjm0uJLMTaAx+qRDACph8dxO9xQX
OLO30brpyRnQKdnt9DomX8WJvVMqxKJUl/487zQU9zJOV6TLPoO6AcFgCzBeKANX
dsQVFfTMEHGQh3kmY1vb07LJ7/NGV3vW2VbQFRB2N9+wRgcXxqTGdWPxMKx2e9VQ
92AC1IDx8KwPUPRfTNYaGztcFRTZb8nxzOXEIUX/KUTOBOFlBKttqlgcHReS+e1t
0drJddGFSuGZLTvUrEURNf7PwS3OBofBkX9+VJmy2ybkhim9v3gyl1J5eu4TAaXG
ZOV08D0QoZK0N8hXKjW6ubXr9RmNqPA3LaG7ZVKuy57x9im6yqnHlOkhQIAvPHvV
ynTMqFALpxKKQEIGnY22lPw+z5+bwi9kI62tbgiq9BI/KsnFCaIZC4fP9e7wr+xW
60WlakCxUJgOmNhf/w3JkPGa4I3eIa62H07uv5gToXAbBMc0gfHQEp/Vn3Q3TKhS
otWS1DHQAs7Iq5eZp1zmzobJduAT3OOlGxGcTuBrD9k9H35g2tUHuP5Pgu49REBd
M6rNXuXunZNI0d43wu7GX1bcYwC3BgrXvDGqHQFsccaYLqiACCbfqOD6eAnjRP8u
iaTnMZhPbFcaff+7PtM/oYjexAlBTE5RAWQ5RnU3RiIQ/PW2AacVRYQUjpc9S4mK
/qz+7tZsyiClYl1DGwBjXNfXdXRyj85OoM0f5TVWZFwWi880JELli5WJFdOgw2e0
kuqTHbLpUzZFROz2fkd9iJMLDvMESO2mDko514m+G/u3ZU6hD7cJ3wmiOJcBJPXw
n5TAiXYvgZKXTesSPsX9kU6F+n2pbGsiyEvyi7Sj2udpvh8fSANR9U60Jmx8jtdS
EGs0/laoNa0ga2dsTAO0CcO8zkdWj2pCTFskpImaUBC/9aa+J1pRkjyFGU/QpHAu
nT0RjNbW77K5skacUwo//EVOFDngDU5bKEo3QB5pqN8elcVa4OTyGrQyYaALk0lH
sKffsfq3RphaoSLCQIyjRqJAGd7Vpx6S263lPbWQGOLmEjs7FjXuYjQbR9a7C6SH
yscN3VfJEqLfq78K/65HnQvsnQGtKucQzC2uTA5uvx5dL9T7/qlJON0KtGrts1IE
Dr1zy2oF1cOc+GdWCL3OtmcRYBtjAWTRevcj0wnwN4YyDTAeliLue8iCACPoqO/F
YUEAZhJJWU8aHbkgbpI8Wxl/wlfRjY4c3C1KfFdp1p/RNPZNalbFAQbe0feeVQpp
CO4nJAromnvEQK6+PCO8QSVwjhEC02IN+KvGQknJ5k8pvOGfW4c598SmIxSvdJ0L
xPLhCbLcRCXLmJofFkE+Sg/pclIqxkFIa46MkzV8VDFXUwH9oxed3sraKPXqQx1B
ZWDjAWlO/CtYpzmvlvq7NQ4QkfXIzHJOQM5zhdtk4ky9gVaGgT2+y/TUPhFxvXHC
JcQrCxf6W923pIXVFF3ZTsO2hcgk5fSszc9It7SrD/Gjj5FSqtnFPRZOfcvsCVfV
xLSu5UjMNcMoYMEutS8DDbyBnTAt1SbY6YUDUdXR34G88+bQ7idX6ZZhL2UmZ+fG
bzwtxalpX3LGVjO+QeBa3ki1syjHa013rhxBCux1Y63efw8SL1piMunqLT0T85sJ
UukC3Dh7fcSL9VIu02O9Yiuvwelx970o1ZVJ/l9EyouJMtm7cdAJAgm71PWj171i
94X6znZCCy+ifa1Ik6DKhePRGur+z3JEZ0n6xd6JpTmHaTkbtYQxjPffE2h/+uZp
YfcxWsjaimk63pLwP1OjUK3y2SnceyitgMTHjKR1XWy1TAT4RekcOoOB+FznKt0i
2boBXUDnROBE9CQwYGg1LfNkbKYybdcCVblJN3ZnTRn3YcVh4CI1NylPz7XTaMz2
xvSk9TB2rsh+JrzIh0ybgx6JpccOQwBrGfxZCWIy6Jh3Frdw9q5gvZql1ZAcEFzy
N0HW2JGmdfEJ3yiunB3+QowlP7gtmnXkARd0rL6qlHPr76IJMmJp4CmfmrBA/aqU
eZHPMuA8CT6gtgijmy4QjILMFZy1kUpSCRkL7AUvPUbGBBDAYM2v8/IF0NehKDwr
yVk/vu6AzX/BB0VQa/TGB6KZfT1HElrWP9n8bL+c3mNuSE5ZuOmqfonzmTFll/LQ
5rkXgrdMr7kavZK+CcyhTRDIRUJnwJZZFjC/SoHQP+0B31Xq0LQrvjjNlZuFqeDV
xSM35CrpgR/9SrniP6g9CsDNe9s1dQW/qYlYlJ4WdTjZsNlNfhNZ00HGTfvDE8Rq
kGpzLInC0xOP16BBQFlKF8m26He4jNf1EKVrUQqRh8Hud9f8cIjR+V6REo4ccR78
TJetrrYv5YoJOXzrcXBIrZcFR8r+kT8cot0fcuNaC+rrGv4B094u4JacmpRuXfjr
lFkAyWW4QGdNFKmjYyARMhpW7Zcd2comkhd0GVwDUQo7f/8Drw1Mva0iEPOw0a9m
X/YC/CWXfeZlsn4tGO6CcBxNh0THsUHq9WR4X6vAat1fxR9u/OvWKExxktgyXXa5
81OHkii+/Bjpu85oiqs+/yTYJcfbhTjDqPyGUHxAedb1PPkjlpS4FrhcX3a6jlii
0Dbt0ha17pA+VRZHy346tw775OY9Li+sGuR3DNaNQLBwg+6lnyrwPTR3wzs02bsZ
4vr/cxgul60FbU00SrVkvWvVlHx3UaUkucvXrVsfXY0hgOm2HVeLuE6eSPl3+/MX
AF9xfFuR20DeyWDrcYE9aKZrmnubojysydOV+2SxH2HZaMmhCS/MgkTRVX5vXCQt
2DDpeZdAa2cW71/kwOaSuNGStNx6YZPHRFWJmZIRh4kL97qpoYB2TfWBa2ds+h17
1fmlkB9rOobJgc6v2bKCE1jsHVukFc9bS4afCDpgdaLR2IRkiUu8nmP8f8GaAq94
zHp8i97u08bqakBEq4A1rvOeJ/CR4wGUP+akKW5LiTgDEOAm/q6UbhK00xinwLbF
PyTj4+93Lbe+9vMHe5ZoSOSznb9LTm7FIzb+0LLUhFU/csP8b/fu/9eoTQGX+7Pv
0gNFd2G5Mkeyc/YCu0rapw00otS5NMIP+/6Zym/n38/Qt1Qrn5Zt7z4oEU12Zkec
IQ0Qg1mX94eOiLtPp4D5PAytmyb1Z3WjpBF3Y+23RPUuzpgaCN1+YaJApGTgkGoU
0SS2+ySdOmcUaPPU3h47YQ==
`protect END_PROTECTED
