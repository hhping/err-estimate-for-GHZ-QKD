`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TsKuE4Vi3WO6au0dX4KTcDCOB9NPghBufc4P10nyu1XoWHoQkme4h+lPM40e76Gv
C79yTRYOTj+Omc8dWGco8huvJV7XXPd9woHzwOM079U1rFsuIlRDIG665q9HzMFt
KjrpW+GHYi0XLKq1ugIwMYXYDlECpoKPbV/JADPgYFoIKICG5of2FuTZico88oYc
zh6yBeEHi1XLIcLaAgouiQOLmglDDfDZXjBCXjqBG+w/bcBgY5lL6LXxWRpohnwx
2afvlkGoM0WTUKZgFbiB79+yzBD+68rTegdLSj/jKNQzBoGDzBLdM8abAu6Y6Ppy
S4L6c/oVWuKM4nHk0pf0Zokdj3OY+Rln/uteA5SLQvbTxrDkfxD0/UexxKkM4OY5
QAPs1S11MQ0ttK0UrGXym/nzkxixjXdLeCE/1nHF9Vi5rC+Bmm+f8FV/cbhXLHJO
eoREWm4AowfHPIqiuuelCVbb+KUVCa+tFYpeKUq0IALOCc18o+OafkXnNyRmiRqd
UA0HFKJ4/1YrYz7cwCWzR8icNHsKSz9j0qOz/B91Vctk2hBTDxe17prt9WUH5BYc
yzYStFaUsqFzCtX52qZ8T8TBJI2DG4Kg6bOWqfC7qUazVC0+w7uHvtqInZR1Dz8B
aRjqmSFRGqfFmLcXRXZ8bQEuzTjY43SCadvlv9Et+Z0sWgY2e3mS1X3/M15Q5O/+
xxoyf6FjPhhOT4+MtCby0WvQo+Rgy5ZQCAcOQ1VDcb8pvways/iOBMWDD2UUPS5a
lgqJ2u9kkx9ogt55VF4pN8NcEaAn46FyUTMmDbULRb/ruupik702S4xPl1MXnQJU
aUtBhH2xf2R5IEAdRiT0Yf3FGGl68rEY6RPHdj5ct6epE+8+a1DDg7Bk0HnEqNss
YW8VOk38T0hZCoP2I+dM3jSXvYHCNIh8Qeeybqn0midmqgJbWjaWDadtC8jrYJ//
YHj2EsclaVJdzr5JPBB3ituJhFfX8pysHPY+B1vpz+nU5q06mbMnnH7WuIm7U3rG
wIzBPjI3PZoz3bUxTRDfLHgVKMDdvmJmtosofrXApO5tqZnP60jf2/P5wEwftztm
iLGWqyg+m3VV5sfCLyRmbWUaCRyowmtmVl5+F3j87E4UoZGQQqlWNzxvtNT/1SWn
+Ca/0xvKs+ak4+c3oqPDa/BeLOnk0QV89WiEntQxsnPjoRsEXn3Fq7do89xW39/H
ydZnCxNCyuDQMECS43g+WMLYGFuY6ifBsBQ0eOd45rh4S+Cpg7z0eBjtMNHFwRcY
lZCCmg4Yhns3D9pzVHTsKkAa1rrlFINvtCYTxg+/gVJyOa98K1+REEF672CpaVP+
ffs8AoGG8FnKJn/Ersg0KeZkLx9y35jc4T8HHNKY9MT33xkxcb/GZQSa6ANV8Z0q
Baa3oWh4Y0MwUayHI5Zz3w+v2ZItK8ogWEiYFuVhB9zbnmF8HEWoFxlL6z06Du40
Dv3SYRQ9ASW4sKmPTUH/qewgzIv/75pVXvbUVtgz5q7gI9OsfLkIMjs6B9nslL/u
VDFS+5BTRyVWgpiX3qUMWtf3jnt8NLyNRUV4JCrzMvgONmwcxcIwlEUy6MGXc+uS
Dy6IJ79T1DJgmqbY8e7xkoTWeIJiJBkg5v+CCBltDdGcgvz5gWsUeXcfBwMhBx+M
QkdOTlxInoKbXy0TFY/J5J8xLN6HF2mr2+SBYtzWutCQlcj29zqwYysIqKRFHYCc
WCGhI7wGzz+CERJKVnV//Bm8x9a0SoYkrTnq51RNE2uzPPjIcWYpKudssjung7G3
PIZ3cwFiRh7St2e6+28eN0nhvEhfYWsB3MPMUvQsPSZbBZKk5+7FNOoZPLvCiNJT
Z30/+dmcfZhs8vPFM3xSNUXLRuib2DxfiMhMjxrUhXgmfYtvnGVl7Dkv9K+uGBJ6
aoxWCjGfFDENmHYWrpEMelW9c8m3zVGNmAuuap7yZKpbf4Yias42Mbf3EI/gmNWX
sC/lrWptU5Y1gOjVNzbUXLUHc9a1V9qj1aMuk1PoENxYLPTOKTbqI/4ZEcbsCpdo
mDTjcaK6JHUP91J54OFHfFZW11o8tk5kVwRpta3c/BDGgbespBpDMLe38pU9OqnJ
pHXqQU0DxbRp1pW+382zLg==
`protect END_PROTECTED
