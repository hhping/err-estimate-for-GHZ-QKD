`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xtF8CNc5lJ5w5Am+GRbZ4vtUSBRaMIQmGP2+dS6JliGof2pDb4ST9GuqTYPrzYb1
0VlxG611dZqYq5jQM7GJW/FyRPW2ZrRbNoMLZfWZ8rRG3H09gj0F8oHrEQlzlNuk
kuKtSyGscIAGKSHcaWfG9kCkBWE9VrwEcmb1YePB7l1/jmh+cGKSGxRzKCfey1WZ
//mGVSDANDeFxRjrJa5CwsmEMI+i4FsGp4200hE/gEwIH9LF/eYuxn1rh3MTZfZy
E8mokc+fVIBhFyS58u76Styktol4K01T4nwqBbbaj7RD1tdfXXbVshv40ODc7cjD
XjTROUP31ltR96czlRagR1U3NKRPTkA524PmTu/685NcoLxUFfCTRcSHkubZGzVV
j0KYewca3LvZKhGf1T4g31Cfe7tZV7SfG5GJLWSeozfVfOe7EeNwyPg3aRF/4MVI
Ar8oTRRgagboxRvhxy6IYZX31GiZ0VGxMTXLVn3UnKLCLU7IEHxgrrneqNtyS+Ig
zUlTRkOizRt77tQEZqy5Knb/55FfZwnxzPQi0mal+BysQjlSOHWaOoSnt2LLMhC0
GIo4eJyAxsFC5Z8Mwo/EuYNy0vxP/jgM6PXam3J8WNmrOtI3N0Uf/cFI/HtcSA23
AzojZTEFUIp440nPrmW9AY9Nc/iQ/jQIxW/YudNBxryS58PCm9E8U4cJeLoxXz9f
tW3xvX1kcFMk/7iXSFGokM2Z2Pyb8j+FvnQHIxVoV9wta639pInOQMCzTvFKC1/s
45VByH8stcyVzrYY29xR1KSk/+h9g4uG9PpzdS7T37m+4yvswyMEMc348P8G2Gfh
4Gv0LjIRD0hZtmNB9GQaXLbX1wWR0hy3+hRxxXmkX1lC+ozm63w93A3bqblI4o3k
sN31AAO5kNilgaT6h2ipQJdqJ63UD403+1KOx3WUnQT0/KlrwzvWbvrc6v3f1+GA
Pwmt/RDg4V2Sg34vJOtZfq7fpcrwLjwQf+IiSCTL3Z08WbRKSlHFGXBnn+GU/6JW
NPJjWG0OKbK0NRun6kphGDfe+eSq6CFYq8YUpbXjFrYzTSImnseb1PBRQSI5GROX
/B8QZdvCbaiT/VFKeM+VNZzJq/CwlgQKOIAHRz+IaaGs0lqmp8i1W2wCowGDki9p
rNawu9xnB4sLlhwAmQwviK3TDOSLXlFaxSF+h/MbykeSXTlythwDAAF/6Wk7YrGV
IieBLRu3eq9E9YlDzk+XEErXfSMehSBHFTwzjaQSdk/oz7Wor4lhT6H44Sy1I1rO
BfhBUajQUnzqJBdSvsq2keEH42GOT+ux4VtRDbOeOiJskhe+rc1jA/z7FqOJLAWg
NUH1tFcWvmmGnjEQa3em0I4eVTU5WTFNCdnkULPwg+/OYUnyN+/VEWX/DNY6Uxn3
jxTOnwSxIEipjwCIWFguNhsHHXbuqm125iwtftu2GYms5knmG5rPanM3v08WGK88
lFymiO1jn+KO2vVHhqG2ktc5CpxvoCMgVcqeOvuu07K7GMNHLG/vqQkny3r1rAfY
DXjTmAbPidN1vHayUkbdxYRuar+3Kt3/Wf0Ay/4XAG5EPKlxAbhEOK2z6GGVbWOr
F/rpIsH76A5oOiTzjpi+soMb8TpT2cYrA+8xxjKvsq3wQnDy7ozYmTx1QK2dDAbl
ZIV+ST28DrsvfZRFdUEwqPT6/GLIMmVMFOvqc69XlbsXWJMmT0lwOsjbK0hCnDBF
KZlDbJqY0xZ9Nf35Tl18zFk2OirjaGr5uyZ+xdEPK23dZ1t/fwBXiNr3VooL06hL
JRpXmZBLS02if2TxE5+Fp3rWEdMaOT/zkMgTXdPCLoAzZ3UcPM3gJTS90qiAGE3g
OGlzh/PrAXmAUEG5xHthK6QIJo+fS1o7AuAicok1JDAHI7gkUNFTg/7xlgkrPGCy
i3T1yy32aAzPXKySDhx49i1p9JMql5fCRnXYHmgR70k=
`protect END_PROTECTED
