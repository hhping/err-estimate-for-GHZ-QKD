`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rwxV9/bIjgaB4VHd2gTY3f9R+jVDdOKGidSDZInmDBE6RqakZ5fd/A7swyaQQB6L
JQfnE7YUpadT9LwYGxS+dqfrAiqq/3Ae32yZOTLWWxbz3kX4gguYOvko5KLhW7zR
L5vvCeOhNZMvUQvVppZ871nWHNam8Tp9TH5eY3Hfq15tTRUjYAHvvCCZyVn4Hn86
izymXIaSP3kDqUSA9piYP5P9UFxfdCQECjMSbJjxry2Z7b6jBoiHdneZSs2akOrw
LEl2VbenFEBTuSxKpN2RtjBEToqDGBKH3RoiYaHXFbt1EYlMQZB6SK2Hv405WSnb
L4r7g3XcR4Mhm2CT2XHHuoq7ZCgZVbNW1qpuq88nxoTW0KlkxKfMMseIZI4DIe5Y
ZJU09/2CrTpu25X3qTfWgl/hp0V6Cre7ASSQ+Didd19jvmXn1zQ3TqCndyCQnZnn
fau7uIR3NLLWggzFADFaV3TZrO0bZxHm1X1lna6JYkGgw7wXuUdrjlD91MZodRFx
zf68+gGhTFcZF+mBAPmb79/xHW1x+tz52xZ6f43z331aAAJmlBZL1z3vitZmCXZg
ZLDPASHaajYaop22/+XkBxW9rI0IJy/T8IE+eXVnX93QdLs99odXhxIg+q+iB7G4
`protect END_PROTECTED
