`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m8akHxbNNCzN1ICa0DM3Jrdt9RbQY9zsCyvTbzCHpI/VHjiUTrqz9uFlCq72XxBX
wdOCXgRdQBKHAI1Bg21wE1NqQ2PvBm1egmA/FfEdLyIzWzoHy3R084rESX/ftw55
0tuJoC5Gbwq8y6lke7TaVzpIVaUa+Vp4EN3sckoVuRM4TdpfIjjhgues2wFuDqRa
/qLZfw52YpBRvByjh7bCKmVoMCzbkW5dE+xfR/aGFz0MLuzkudF9ZQtSu8HOLRwS
OsCUDExRtGKfp9To4eKhZ4Nee1cDszkeWxxy52eLBRE/FEv/m0MvTizwImkIRuAd
n0x696f2sjXmfTRtrLxi1C14sEI4jjOgAxYsO9WKAvgQv5T6o8xC1R/oXKZYi8B4
DhzCMwgtM1DnQytd6MZ2wDOTKjj3xIOaCE7yBm2PmjxA7otPazmhUKf3o95nog62
oRIc67B5mh2vlZCPCUIXz9Vc106ugo5l+kZwf0hrf+znQ+edYBetovr+lOwUchH8
W4Yub50D83v0nrVRzFYlgPDcJRe9KNHnSGcoo1v9HRcaNSZmjZ5axaEvTOrGqESW
t4gx+qaFGIwpsj0XsUl+pqcVf4DuDzZwRG1f0bvTXn2HcSBOSWZEybIFPTpRolH0
K9TIZJGht3HQs3RgGNd5FVLPhCh+XcqMujJQ8HSJSGTTyJW9jgozJBPQdILa+S5v
ydXtrnmWoaGIR1Qt5EVCDFXdV9nQcCHHmL7jETXGn7p8enTk3Z1uliB0oUoki/F1
PBI8eFNAiyCmvjY15UfDYBTWvskQF3Rq7xEdYkmoSQYgMjMc95HSAyJM2UpXXZ+n
Wrzh0zYLmmh0R4DkDDrfUVlShdoMC88fMdQiyC2xS2eFKCnpv2Fy13bLN8cy0cKo
dNGPkoOOshsiC88qvT9ZUsPZ1vY14Xp+5Fw8W8Mn2jkF97bJxua1b5lxTyOSbQK+
4iCfkCXLnsGalAJUFsLdcmU4DJzvQRPAGh9lS3JnuorSmLIbi9AnnTCGsGkWcsiE
k+mU0KxR055owFCcj6Syst7uF39995SnAO4RnISKD3seiPL0z0GA1gOi2JAwBKIE
7qSCgLmB+hJap2mUtddavYxGeTClp4yGUQ3CzPWhnkoi9LKC7YJHlpIOqlA2LL5W
pdtBofLokrGHJ2s+A8BoivFwe9pDO6w76OLuio43zMq2dxuq/obvc2dVFIvaQnU+
7RKghmoMtA4iTPPUbTPCfDKgWArojdF+szzlyiFAlcelBalID768igzt5pQFYFXH
DvOR8bsAqi3qn0SLhOTltq1YRptAkgZssukwhXoisHs=
`protect END_PROTECTED
