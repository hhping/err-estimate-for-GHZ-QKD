`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O8jAiD2shNUGHVH/jBs2FqpaqRVIuOij/orFV3uQ3kp8uKYuHD1kjxCqRyr2voPB
wEUiDW6khjQwCGTeVWZkK3NSIhjkzTjVb3nM6jbmSd0wMRwJ4nn0lq+JC/oUfXr1
d8Xv102Ix4gxmon4SLum02drFU1kzx5qY+EeOj42rZ3h3a77P7T5iOB/2fECGthW
O5JVnlcHwNagA5+tVh4OSvmjtwbx7GzBR1UYBmhCdHimTMRahLZOONaTkKPn9We/
+Ntrto1AA38gIdte2RMKd0a64RCLVF9umPWW3dhufo6P9fH7I/lPdqAf+X0L6B/0
zDeyoQDqC+BzGvmBoNxRUk9KhhxytuSPLA7yskw1ww0s6jJDvHMwPS+fJRcDlMS3
oZ3rXdsJDMupcyYSLfl0lFs/EN6ouXwHRPLmANGQv2xjyDeMP+dLRkSSNVqgPa+Q
MyazoMujwV1xmwXvEk9PQ0gL9wmagGxu3YsSI3kqkXSvwGTera5galr6z1t/96lv
t0P4uUP9smiQcbi8Wy+XSMCz9vdh4dGyWadzUMsurov5348qOcUcj885PyAzJd6K
25WqnS0O7Xw/gIVWWGS3AAz1IeEjN0A+XrlEowjhTgBYKX0YTT7CBKZajvLoy0eZ
69b06Y8RhH0Iy2teZTtgnzrMv/W/teIoRrf9IFKDqZlBxiGkWyklrRuWx3mT/ee9
wkujl/tMjds73N/rUaZiKeqFQkVb4qpI6VA6NwCikdYytGjXqy1k/dS35KNLc8FK
7lu0GR1nO39rMpiTd8BxqqI8LaEv4+6uN739TEq/eOP56FXWfnEFnuMy8nuVL6w3
5eTMEW3iPZIvCYK5V3HNdUMIdRiWWV9aq2rQG8K2CLdWis6NGa2ZPVBSE2O1WuHK
L8Wac3F74oaslPZ9shW9EJ/gnLouG8ah3XP8XSRDVS0fetrDHiCLK+kWcREY1fbT
3MSkEHD5J2XqJfkcKdZHtxnG72/QfMyJ75JSGK24qgz5GrHFBhcFBQPkzcytrrP/
L+vQvoawgUxZtIaZ5IVtTDk11KJpusib5SbLiZwLiafRjIjlpeHjRAwRSlUKhWKP
ZnamfG1KfmZB8VVJYYr1DsFnwaZw2DMoIU1GRsy48hPvx965iHHtm5U83MoN6EpA
`protect END_PROTECTED
