`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kucdjs1OMyt4JcSQJLvCp9Be9b4oleBaNmzJFpmW/S94/8h/LzhggPp0d6WBqXZL
tJZctdf0Ua45pynH2m2jQR9SEBJme5YJyiZ4mRKk8rJ4UmqBcyWVDgW1RKyrTJXQ
yFdh8CtyKGpFgGkNzZEDAiP9A/mHiwt/8XFEQ7mowjDhaS2w+9F31Gs7eGcP/q80
uHbjE+1w3hEw2SS5IjtDhURd/taL+IseQGi4kAEHHLF36Ds7Cv2Ke2/JB35qmD9H
7ooyyOie0BHutQTPElyVGnpSrZOV0aF++ZnwATsHRDdsQ965ini7Oc03z9LhE4qB
dZy0lfXKi2Q/KQ2F5/ZvV1Y6RCIeQ1Muv9fJLR/fMgpkqkESXCSvCbnjPSCe5c6F
3lIlEoC4LFp1sffg6xGIVyi6U36uTN1PyDmSDcd6Ueciwrzd0d582d1cC7Z7qwt7
+01EJdyKSu7/6wCQRvEtLFXcy2JIFsXEVtku2cpjMd8sctGhhnQVCEXrJxjOnGD9
zvgRkKpA0RL5839KPudxvnaN79yvqVybpsP2zZCmyZ88Tc0LhTX+V6MUeD4+HXDc
h/zNcKVSu94hLhSajYZd5Y+PoTnPRFdjmd/CV2MgG+KIR8wEF7YK6rSMC3t43Bnh
UB6ns8mI4CiOLcvnlBEgxChdXRh5oLmJ95wiwxbNM4VGTP5PtwbUbRZ4z3g3iSVh
pLguQu3AWHwjGzRu425+LDM2stQYlTw99UtYW9BoOB7MPbdM/ji9dNvAsKthNnD3
Yfd/2nmQALodY8fMR72vzWs6BTHZNxEOaQJbdtnpQrH8AcZNDeF0hnoCRWk1k09P
x+dwR8MkLu7KtVZXYRrAG+r9itqKHyJffP8HVRM/byhnTq2sSRIxTAgnKZAVsLNK
EsUK5PLMl3zuS8Ti5dQW7yEPBjsjfXAAS7kEbBGkrT1xG34/WQ+SgAdZxMW3Fy8q
b3ka0LJFfIEI+pbVo0HTEpDEX5oboChif1imxXTajHIyCVrgG+QmUw8Hx09P8gfY
NTm/T4JQxktauHRU5TPp7JdAAZWY+wSmdg9O/BKzoPPElqxoq1xi2jP0h4/mi1wv
gpDfcrgbEBzmkFXiqt/kMe1fqJiRGX2jKvmABv2+bxi+spERp5WrxTqMjfpcBHFQ
gnLXEiGaTzykrs3J21aA8B0Pp7urAO+JOEyb4B3FyTe1M8bA1vd7F529XZylvpX3
XifrvaI4d1Pi5gBmmzLPGkr3kKY9fmncihKwLLO1T7S5bxY/HiKi6XEEjbDr7cN8
MXZIEqcrA9rVvF3++sK7P/z7rzhJqjsyX0b0ZdngzzVagAtzgqCDwkKkzoOAk3Aj
zMH5lzAd2StjVyhQv+PIEP82Gk3q95HUM4ECiOOtxAoMmz/mmR33qrjqQRAWGusr
dH77hFoDWZ3YNPLTHGujm73uTnsoshhD8RZwRiwr/Rtf6bf4NfCXZOcDWsnlLDuR
RhjFmDdj/X6yp/JTC5JDNM86ihQWfYQWdq63Kumr5hJyTaePMmDT8RjNL8n6wf63
7uQ3uHHViGei0Dg8SMB3UzjrXbdXaIRONjRcNq88bpqToFAFSopBvKBtZK2+6Vhi
ivPQzax8rk6ASmtV7VBYYb3Kg4LpGZ9kiZg1aOXsS+i6ZHm7GSAac1GofVgaOZ6T
0f/1636tomdI/JxuR55qNy9ONdzz5ka/1WX1Qh9jNBMtHiCZpmB4yW0q/EURGvcC
dedaaWCpiVl+0wIWd2NayHVHgi+csyCRtFx4bYpewyLcGfBUB1EhY7NC0b3HlcU/
82Q5XgQaBGvu4bdyH/EEiHOD2mvb6ibY3/5/WifV15/SfRVt2Bk61m5+OuCxL1xa
hfobav3YI/m8loqYDy/cTenvjNotqowRkktPToKGDa9LH0LhGwRyXwRbOSfIuHCj
Oeyrf3XPFq5TR5OSgx1/45vkOHbpsIipNxdv5kd8OxUa0q4013Eh5sdJ01GbLfF7
eCqSQu9mg5FGtp+rcqLYKxNeaYmaKlLcwYN7sjKzc7KtciobreHbRRF39vnIxW51
5DqI2INgTQVLp3l2Nl4OixjedCULxQKPOAMbnXKQlryOkKh7PRAi1hAGWins4D7J
t5WoNnYefM3I/J9nvflLH5TghTTjoBLPBBb/8mToY5ktAmsEwWRGe7zZ727YRemx
GbmgA1rSzDfjQKCD0nz6dmvL+s/RFZhhp9L07++SrML/92IcGZ1Kt3hWgqi/7cEO
QHOwPKZccgTxkp42/DmEWZRxoYLDrqme/jnflQ9vlvdpn+fyZue7FPichvtRHEBS
F6iu9h4iRIhwGJoqqK+sQ8kCIsUQnxDgstqjnrUpPTHwV65n0MEETGFuKdPU08fc
F1/az9ImvIxhSEYkmQKTmO9EE5onTKQppUaJ1IyTyYAv5uAh/+K4WQmHCBboj5Tg
AVYO4xUuDpPgLpaqR/VUSd74oxkaIl7zRVUr9SXgZewGlUIbQ+9Y3CSnJenKlDR6
nF86/mmTsyolUVM4Vnc2mK1yqj+Y1tFWJDq07uf5Z2XUKiePc4ZdvMo48/0v47mZ
JvrRz1pg7QSQGTTe1QtMzTSg7fl31p31HgiQ7/qkgT6Cuud4e9HwjLYgnvGGwoQ/
r84PUzOyRP1tRPrbTvTajFn0Gw2b1pTm5kCPKiHynLq2Wv1qlIOkImVOcBgb2HhQ
0ki/094w72AgwNL5f23KVmYeZpDYFcqIRY9q3/TSnFfNjHyvXEbayjha4G01ePo3
FZ9VYM4ho+5VyzqThljMOHQ+s5Aa+oM6xF2bcZNTxbAenJCgrPoglrAeNApJCz2X
voi/u2zHFtVCSHjgmT2RIqYv2RnzVXi+jhykE7fKpWyCwEB1huthdAvLYOI9gQj8
YsIcgcGBB5hpjTzlq1Pd7qbALCkbZ0DV98DrrpG9L0kqIwWOdng33h/gW91YOgId
u2jd56gXQlZfVLMCzmjqhkknsbkWWjsG0CrW0CDre6fF8hj5GfrIw7Mi/acd6oGw
Fk72CMc1mraj4bKi5oAvSzqGv1FtTCGs41yFd33FqsUC11EDr1+5fji0hID/FApU
k2DQN/mnVT1IuVwbrQIr9pGBlx1NBMBcH5w6I3/ajL11zuJCVhj9dF2m23m35sQU
XKtAKq5rNuSThtwAQvflgmp0JtPhW10kiO+6DtNT+GXZU9D3SZKNJvmLcyI9TNbu
seXD11/Zl+wAQAbIWcKV7MFY+Jb3bIoBNajSetU5aN9/WYvZWCFktgIHOyZDXbET
zgXTWjqtr1Kf3i+8fSOlvwKdUXYPjEnGvmgdlN15n1qj1SJgc458LPMrgx+itBpl
hBp4R34Phvf8jKSDHl2No19pU4K6mm1RXDF/H0fw/tiXT2tZgUIWURVc8T0MB+nv
zYWxsli48blU6EUkmS1MMJHMqHJ0zm7+L9QNod8wK8Fv0bcqCKhN48ngUFU/Y3//
EXJh4nucCFpiEhvY5R3wFHDsMlTl3wi/C4DhRPZw3i19g5KT6tJbqI/XKUUw/0Dp
sxajXTkfcAoME8J3wuZYGu+fMC5FOf/TvEmMEZRZ1yoSruiNLlx9jDj5b3cvVUvu
dN1fkBqGl2SlPWhfOClTgsHsi77mmstyacDZlV+u2nfhguvx/KnDIBsTLcsmS6Uy
I1fnLn9qpFE1da3LhVVPNWC9TVdKq470lQ6bYLW6WlsId6iLRNAvqJP1XYeyi+/3
0Rtmw1x7dtLmRG2VbIGhXGkYMVWIsYwtQk7dyhC9Kqs0IpblmMnGVNrDNJdsxTAg
CgAmvlMa8CDdsFMwzDMkIgTD875WpFfKuRhH9CJjQMj5roUUOuMCqjGMTR/jrSa8
HvmDCNTQaDPn/cmmelFsVvXJaZKUS0QPqLOPwIIlhwMB7huiqYndyyxywjhovD2U
76YWAdJBCjsioBn/hR5uNuvAVimC9ezN6Z/5iJPd3LQnGGjgqn4hkefsKfCuhE7s
urrHcEclGyozvNh4mU/HTA4cvd20AMsi6ZZExiCnH5/1TKZh3FkxGDrv7kc/Y8bE
3iQ49AfJwbXdoyoFLlf16XPhABYk7NkW9XAl2PiU9fB+MlCbytgOGRZ4WkfG1ZPc
9vRztnrP3Q+qMHbzfu31Mp+pT611zyabQu2kOzNvQvQUZFW3spjTAbnSW5QtZZn2
WAfffh5Bnn8/qGIXOk+ZspYc1cd9P/IL9le0+UgXkJF8nR3LM1qSDm4yIJYf5rhQ
lYeWs3eE79wghkk0A/US+PIff8fXGcbt1jxT2cwHJtAHsl8TdLAPZkEws6is4tcY
bvQfhrpREwGPIxN9BBnbjjM81ETXHwncb1/CwUYhdwr8VfNv3HdPLTmnDqCWmE2F
70B0SvMK4vz1/uFPeKwN0//2yQsbD1r+uslT1z5At/+9DDN7T7HsEL49kADJb2Ap
eUsJ1JJJO0NcI52GK0VvDSdrIDLO5wSfXTqV0bqnPT7AVNRZmXAUwHhD9sIwNZLW
IWf7XMsx/0DjbqfRONBZZ85WPJu4gNJPXxNgdWby+WQk/SAw4kpcUeJHH0OSyfee
lFJ3b7MjD67YA6j9QC8MbH0g5RE2qYJQXAK3Scj9xVp3Wol/3vlLtcby+01Geeur
VlqghpDBi55fwht9SArrABTlNM0r+6S5gPifArPx4Ntq1Lr2dJ3pqChtSflmvfJh
gu7e28EFC6MVcNuAJGcjDiFCvjH6hq8LxXfB0gHZo4s7yrpVsXBGyzR8wzDhLsSo
ULO//l+ZIB3EzwxlBtJlupP45WiDh4SHwodmRlnYQ6cPtKo78+9XdG1ONEHDr9aO
shm2jxk22Lodqdr1XUVqLqYBfXPSFJDyZnVtvv7AfAuzB1Pv3Blaenyb5XG7yedV
ly0g7SLcAhdkXM35rK/9C4I+fjGJ5oyBwsaF0TpXBbnwT76N8SkKQUIoxCP2cT0f
RTfhw/rrtyMqpw5jigyKFU44Gb37VN3JR5mM1RAxh15Bg9qJZzj59ttWzMX0tqnm
RCLArevM7Ki7BwkQof6/hwdzBA+ocF2sftFLE6yw0wQAbRH0Fbb6blPidqxlt3PF
TsxoFQ0wlbOxCJe79FHbiossvJXA0NF/r43cJz1ggLySwX5GlUU3/xWeVMj3fbNH
SM3s+ljhujHEhrf68qmakLfV7MfUMhNZC3qRj48rK+JtrY+JmWukw/crQrBn74o5
fTUIWUVSocyEeAHFqp26NGIS28hziybedBsphd3lkHIalk+fmEcXDlfs1RbHQhLM
hnCsOvkVNrG5jbAj8ShG5EWVxmR2Z8g69PBmTIN7uhP7PFwcauycdZZJEC6bdLsP
kk8qHfYjR104XvnEngusxVl7313L9Z8miruE5SAQMEZt5Rl0wpdc2UtBw522qIjL
ByA2UcxXS95+qNFDST/xdT0jHwAyVseBToWVcbXsuRF92fGwU9fGOZcxH1jhusxE
Ud2/iCX2fFFq9TTMZWb0JFqdn8oFzkShvkP1GQ1m6AxKzTjV1KBMbNqwp/c5cXfS
YGP3P551G7nzw2Yn/pfddtHHbG8ye2lwM9+zA0XRz2gKb6yd9g8uyepNGhto+tso
Xjsc80sRc1H/CbevBhFM2Xxa7xEKARWrIlqvVMLIGLrcChs7Kgap1ia5xllI30P/
VIGgay2xfDP6I+qOrVYJ73V6F6VNCB144hMXu19NzWqaxbWIf7B7/z35h640L10h
jJisyMaKt6onk4baWY9saO33ZZ8pUjWepXFBo6SYohsx0uPRSK8fYyGPXQjKESdg
KLBjuJkZEjb4vC7hPWeoj59aFCzaEYyULD3ROF/5p88pXs40DHOq+wuKrzNXL+8M
L9ByZnNCl0kg9Cio5J2kLhNyT2bOZUB0xTJ+hWCptHcaAryjM/SfWz0JGUQGgXBC
MZWnwShOMkwjamdgZKzdvPzPmBHYILtYOtankdMsi78dWOFGcvz/+laXegmq5zpp
o0u26W8uGGG4NSdtzUJuk1W5KVB5Xk1OWKeVsXeNWdb90JGXIr/EypuxLSNjKztt
okGvWxFxsgnm+R7zPKOHDz8sziBBu0v6DePtPCFiSj7qW9qEQ/W+vUCwtKa7DvQv
yqYb8aae5F9j5PDi6duyj0U07OaJ4u2+j1q42B7t1a0uEmCz86G4xDzAlklgSH/7
iZdzW6ODd8lzbakU95foxuVhg3k2n/s96amd+ZHB+/Q4T9kSDxmXSG+E0rubQTk1
wnqOZFT5kiDblsdN6Vd3MGz9+W5CLl22koc75Z9xX/w84Y7BkbGlo3rAWOhJ6+VJ
DfLIQLQiPzo2sN0GSwOUdFdCCti6c2FgWfJvoEbNACvSKOcy13At8wW9PAjTcskQ
aSAN+YJYTHRlSagFfeBWYUBqdzdKkxvcy0lKyg5cQ0pwg4IoIUGYyFbILx6Yax+U
eT1WJFZxMff8nrCI6A7LZogkB4IzJoT0BH2m7RDJ7gmrHCROSD/3Y0usfJxwH/c6
yKNM7AaG3gL2C90jT94drv9Nryh1Jb52Qg8t0N14WfrJcsO5WgEURA5RRN3T9T4M
WV+f0Pu12s8DUIpql0hAaxfWlMCXlZFFK1aRSHm99M7LposbfjglrYnJf9+++Xvp
Z4Cgn+YEx3HRbdQBToaGBxz7lN0mv9aDnvBGskGViyJAXKehHoxUpD+m74ZyQaJN
wbS5GZ/yh/0cBQe7LBghdIJKwkITcEevWYuTKifyRxzuOPnPVlOONYgOwAw45sG0
cJr/gK7cRKIPRPLkm5C0ZR/WXfZrQP5NNqjZhFlekR/cMceSlH2QQczYLFeJmCmv
f3NvmWn/LIDtZp82Mg4kxvoZlBH3wyNn6TwabVCnnv1zCaSi3TXb3tL/tFUZiJ1U
PeAkF8WnJ9Fw5tG27SSWBu5b0o8atgdcxbxemE8I/SF0kTE0iWQSGGFkdCXL8uoW
5nHAxKXA9AJZdH6SvyYraIYmvczu7cpC7J7HEUVtw8uHbrplF2j2Y3sLx7mZOxNP
nnCB5KUnhvvSLf43IRqTkkr1DnYcx2SnXcw/7rQkwwucVwsPQjQUBL99fPYEg1Sx
k5qSXrlJ0Cjn3UT9BRK6IdjAzaWMQbpbj+2G5I8PIyDdiA7ZMG+1UcBw/NbGrWum
ET2NrZvA/SPy3kWYeZfemrvbOA36bUjPaNBqxr8qV+vOnkbJXjrdwVXaheL5Sy6O
zF73Jh+egJQjUp3ly4LvcmJ40M1AFdA+UdzSXwXNfxFuSn/+FhrjZf6/Fmx0eVu0
CuBDKy39E65yig5rGTcPQynS42kqQHtkokUu4Nc3YdwDoDZSr0d18kWwUam/L82F
N0eTXOtGZkQXGdkLJb2IlGhjFpDT84qd6MuJWYnp8muK7M1dJit5nxMOX/jC5xgs
ZPdC4HHbLw/69lkaO+wO65qDO3JC7lJltWo4O6xhHU+aqlDQBzlPx/fKg8g4on4K
BLhSenmClDSq8kQlr2LgVmrYWX2v4EFqNco3l80jgoeq/dENjnBu8xH2Vl0Tscej
IS4I/iDsqxXMdqAHKAmnyDoZiqQ2LMvGRW3AhSPJHSHWlETFe3ASJZhGhbOfmKQv
zuQqZWy8FDcUPSMLkIiKMRFOW2R5tNUV2n8wmkC6TrRDYxSGz6XSPfO1DA3FNidv
6wu1uPTns+HqWrusWHb7pweQ/UH+k1xDZX5+0jMjiGfd4U01yuHpUGzanadBWpik
tKZWxHcuAhukg1yvxm/C2JK+i7tOnif28JcUqK7foMj7B3ESVHtXax81czJ4WgNW
EYs/F6X1rLnYh0tRJn7CyCvbwUls8NAqk7iXemVi8zN8lGPJxkmTevYb8ith6rdC
0ljMSb/rVxAOX1Y5abs5tC6lv4PF0VPrmPnq498lhkm/Pkhkkd66CVK26K1mC9bA
cPNjQuZWiQvIAz4oFjo2BmmPurLxKYcIx2CqMAlJTIW1dCH9E/UGtqaF9w2uMKUZ
7U8rYxaww6ffBvTYrTL3BFkslOvFmLkgddeEQYuZhkE68cFq5qtJfm10YgeCsQK0
juIynFSNn/ttvGTKdc6vQZ4YJbJ/96bgdGlCXaAv7vhysauvtoZXTkECPxkk0m7A
T54nhdq59jYMpWGSEFHIDkq4NLCfYlQf2XlWvnGc0KbX0480qodvL1WdMQDrbkBK
+FlnkHLp8Ttaqdo4ZsYZ8Yg6/I/l0X01pOP6bajonCxzzLoNBI71vlmwA0xKZpVm
kzuk9kMPkaYzBoPmcd2DXTubkj1ihJ3qzgfc+lFbKtVdmfu51rkx2HdSEQI+/uT5
LyCqmSFJhNm0IrWA7S6JHO7qZnoJ/+aP0TrtzxL5hm0VlpRNiHQEMfchT/ZFxMYN
m8sgcawcou13Vil4U+pTz1YpGb0/2RCPhXDreB6TO+8Fd2LTim2QZY2E8EFzJCGD
StMpqZD/8QmKqBsXAQqkgfmd/A892Yrr0MrgC0Z99MHp1RnlYafl2bbbDDYuRmvc
waaLIizIe+ikT11gqlDrlcVVsC+Qp/Al5cZ5+5589EM5mJ+W9/tvzZTP+pLaeNe/
qRn2wtSCL1uh0S6Pfzy6LTQWqqL01nIrpGUzIJYTRdk8rr3ItTnI4EML7FVnZSG8
JPnqX0vsI0gnl8nKWfvDn1TNcHnOclYe8QVFKlwd5vYUW4/lu+oQgBn5keFj6nCS
Zyr1weaadkGikp2gp3NEc0eCE1BYckVD/CZq4SzXVMM84VS961kkXWqHBoO4P7E9
xaQQ6d33DgEvjBq9qQPBkstbr/+5XIxzwIVOKzW1VAh2ltAxuspDFFH2H80WFU5+
ug5JWGE/oQ0/oftnv6wgxBEL2gl3ecUJFa38IzN9XFIruNIbLL34HDZJiBEyvLEO
TJ87L2AkbkTun5mvI9i4agOZym/tdJBx6nw+OwO3sLrXrJ1tGICHaKUSVoEyVe5s
1lkZgV95SQsVAsIGMUu1KXDOolUd3IJQTOK7VtDpngYsZ0vVfRGCNbNhFQ4ceJNo
uvLyBgkm62B9CZjASJ1TBme19e0pZgnJB7yZfGHtI5YKlCl4IIXRl3ofSn+ptduj
wm9z3LxAl9zyeHHARlErnJ4fEYO4+KPApo5ylfBwnCDNYUklnP3ZW35sxYv+BUO+
nrNNn1b95fvzSeOzGU1Q5T76H3smKVF+V5SiwuRTG33sjnFr4u1p3zkCRKtwKKHs
6BZaPixL8T+Yt9CxihDBal/eGL+Oh7/2JFAfDhh5O2wcxYPeNT+V1c7RHV45AuMW
4d6Vstkm0xIwMSkV4kWYpnBLHu86pFZrxIDhoMxz7lpNBzqtGpV8jbcJCu0I+Ezz
C15H07BRokQLSgi9faZgGbdv5xUtf4yYp5pUkQjuxJtgW51yXkWwYLkoUVbihLj0
dgiT76ifGl6CoFFG4uwYHFH+ipnNxPryKRiSDk6p0wsFtej2WvqE4y2yO4Rkud4c
SCGetDHcBn9/lgmd3UJOsByDN+hOUvMmbZymoxNm+Wb+3q3rT0CQzg2chU++CHZ0
+tA+zfU+A2PLXTEZv1wxjZxUjeAHFMbYxR0oizQuKDuMb02iyiUDaqskQYQWiKb+
p3VT4qzaYfL08wlQhSBtiuQoBqhnFmYhEO3A8j8dJo4pmL+S5Hs1k06XqsNikV/j
Z18KZyWv/Koi9hGlkIXIvuFm80S+/+5ECHFWPu7VFjtRKdamkIE+1cG/Duu1BLlt
XAajZFSd3kOiu/91hnT1/zEV+/+KANCYdvZ6d4Ezr2zfnAJ9NDZnN7UUGePR89Hh
3vdDgnIZbLVYNk3OwIiAeEhPwUQRkubuF1jPKTtrQj1rJc/NIpB3ZUaXLXKmS7bx
GYJxv0LsBkr2DZTZXr4vo28cFYB+VYa0tHQGsXCsI77sZV1/HIpm5rYIZrSHYJca
S2i8ioadvbIW06kczSyWAtmejaNqbKGleIm06SIHSOzW/53fwxG4Ze4sZ8RPJOBg
qktjB3zNU8NBwuhKF+P1gX3Z1IUzJkoDn0+1J6ybc6zAcFXwiRdlgI4WE6nf3b3Q
jOQ6TRe/J2yE/Ex+styLBMAORZqMA/MZz169p+Vfp/J3JTThWf0NL4ZjvxOnRGP+
yhtP9WJi03RN+UrM1RNB4AMxaqDoT8F/mzYw9GPGUFf1PGq5k57kTa6Oof+2REyx
+dseN4lMtfycxcn5ZuMlfBmmJiA/5sBWj11eqshwLOLhUYUoHtoUGKMuLtnf9krD
GwQHyq6KYlZLHb+DrtB/HWbFnqkr5gAfGJB7moCdb0SegZ20DjHcYrrR7hDqt5PE
OZVWTrLFMiHsZKliXWsX0R0a1vtutBERyvfR4HckqfE=
`protect END_PROTECTED
