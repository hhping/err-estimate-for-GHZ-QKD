`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ANjx7mP8+tiTTQlW/w3zyOt4fGoq0/0r1WoEyDkO7x5sGfGMiMDUE/nSZ5rc1Cai
XDNI+ZFpW4ScBOJ5yEiaWXnytuLSCxl/g9s9z8Z8oNfRFRiI3mGxWDQU4J5MLCXW
T2hSfgROxcY89CG4u2bkSyRcY4yO3eWy0CtVwPLilLEL0BEbowhvm9iIQulYEwr8
16E4Eg96Hgvl1uI9RpWHm4QNC69OelecVhNhrAMWLsHtOHqMzOl2NlXz5LrtM5Zi
dKY2iYUbk2bSk9S5J3pQE+85AKdEXEz95SNxCvrfSjFFIYiyInOuhHn7gpxkVsAJ
/b9nmhwmQ2Dg0jg8kYwc9vWE3/Q5F07AoahBZjX8MeG+P4EmKj31knEx6NewfZFf
7NODOK8HXC886NU9QVHR9PR5SvXTSHlv+MskvXd+LPSsRIKwI4BCNcIBki2v6Pbf
JqEJNxACcudYxSdcA14jmH4NxmH5nJfCS+BXYBakVMBmwJvMNAAvyueA3uS0Fb0V
d9zB4Wkk7zLzNFRVk+eqWsZvpxucG4hZ443bIvlisTnz2jMIaHaB720eR6cU5by4
`protect END_PROTECTED
