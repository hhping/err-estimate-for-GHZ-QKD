`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u9RlSBr/CDjboIhP/j1fUsX8KqqJlfX3X5zCKO1aQUoujHXuDnQp5YUwuQpTcKRU
PdI0tYju1zec2aJGldRz7/mb6EhBrDl81H9egza+UVcPRgypyXL3+BtzGCNXtLYI
VXRTL79niOylvLrAiQBV5j0dzXyMvcP+QlWpa2qP6jpJgnG4U86vCU22bR1h9M3d
0Zs/01hFuKkjiSMy3c20HuawiQ4y7Kr/JEnco5uklZU7ruPgFLZQIDV15sbKXxYT
Io0mycbWHhNPOLq4o6WZnnfAzZCxzuXCWSg/sP8jzoIIFsZzkxLvouJH9kFQ2J7p
O1lNlP6cGg1furfPe2cyMRrWgL6bRKfvdHd5D/REoHgKYGnG1/yx7d0tavC5UK9F
ez204IB3j9KMyDxHZW1FynEGmMjNzsFNe6FMXqZ55Xutok3Xt1EFqaYS8hB2/D+z
NMIZmg148gNRwm4u9E/G1Iy16SLP+fW3EwOVh8RwQ/kRhAQP8ENNViQf/dQQSaIG
6LloSHUDOjSIdycAFE8te1TKmZn4F1SHMBexNJKNyZNfvJ4TgI+CbILvASUH6ANN
4lAkOXsSoK9paqxmWe2dNQYfhJwQvpoTGOCNoboNFH64hhdcC3fZYp7HE1TriFKR
BbPsZUUSh6Dn/paWLO3+tNL+FtHB/yqTk+2gseSMvkal2sQILEmhkdRKeH0f2My7
`protect END_PROTECTED
