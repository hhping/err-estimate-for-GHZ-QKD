`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vrqO7LgleebcSG44VKZJZn8SpVT8oSXkiC75w6BfN00usbyp49lrZQHO/vOKwO+R
qsvtGs40Rra33KlAk+wIE0GgwAeXwOJV7p9KKAqjakY6D58oyha2bSbLIvOUdaEc
vG/WiHG/ktzJ10L0h1+Tes6Du6m87HfRvlrKuuKRFjGcoXjlXJZoes1RVJwlfqig
Ee/j+tENrDQn1j9oWVHsHlb69whFe3OfeDLj6ACPiAnBoYj6K3QRDJG07vRpLod1
GgogzIUP7lo+kU1AR4IYsqR6LzBCvl6da6tp/A7aCiuv3vX50tlOEWliB+KeCaFm
zNtC14SF4ri4bJuXOTssN6zT9cpS8+XB71IYMlnuIkK7nt4uhBj5OAGZrw8U3VH9
9naz9m6YiXPg6ScdxphaufHKxOGeO2b9ta4ZyRCX+fn5/DkLO59MZ7Z/3USCyiie
UsH2ghFT7GiB4gM6lNS4RSdIQqkQf3iyLy5UcpbaEbhEyxLk70z/nlIihwvpPHw7
N8WceRgehfce4FeGicaMZoIy0bDuFCceKEHrQ383+Xv7DzSFwXEPhQ6VJjpv+2pW
aOBTZEDdnZbkXX+Ri5Tp/ltqsD6Q1OxO9PXf8mUIxLd5PFD/MXJZps1yYl2GPJ+N
G+udJD7XkLMMfBx130ogSkWIYqF1sNKlzUjbRsXqXEPju6LlFwmdViZLIQfdAQCf
BfKBXmnpNuLz2LPhsC9hZBHVpKdlwEBtFXuePjMWsIMmo2iJcJF0CnXB0TLwv675
u0qt6EdShiHW45ULUpkcVgtcaAbHmggJ3BPh9jkx4Z+7J2NXv9bJBnHgEU4bUSry
hfDTcr6XrcnoYZ/ceUGCczf6ZzPfb5Am/0ydA+ngD8CV8dbGAZnhRY+55iHE81uy
gkk1DWKBzTbduHucMzM3T35dFVCDvZut/ftj7LUIBFZfwIpFHkuQNb8/hGSJ2my7
jp+oR26lD4/RL71Dk1aXASzwGE/xjnv6WJr5k9dVWVqNhEgEjlsz6fMnmIhOMJkZ
OK+4HBPxYTseQh3vZuybR0TKXzHnq11ImGGZDilxhP+3d06W47CsOVc/N2ocn4kw
cJHE/rWniazU20zVPBfnnU/SIQpd35hJtPFpPYIe+yBrDSa0KUMBhOCxKwLO4YY3
Si3tXMmFtAR5PAYntRuu1Z2j27MQsVi7Og1DJJUII7vm/uvLRZOwSQH3aDLHwfDZ
VMtZ+9PUkAuKMsN8jKXLMVvcVp5FNnqM9MT6gtv+wl5WfMo9+W41Em+YjncqUIPi
oez++unSurTrXFHbvWAU/1BOvC28nmZ00fHH8vjx/In8mUaochpPETQLHPGvSlmu
S2rq32lVk0MkZDhwBuNJs26fAWv5JjKP4Iys8LQKk+v5T8hbGaI6Edli8/Dyth+9
OkJa4ZHc177nfpdziYSblt4XdIgbIkDudY/HDoGfHdG7bpSh6i753meDbX2OqtAv
gE7OqhK4RgdDrPeDq7noiBWhsa6Df6cLLdeoqJSnZHskavZNogd1J0RaHtL1nIEY
pvTTh5cRaLCjb0a0dmuYAfgDB8ltAv+1jFj5lipg7iEHCWwruaql+CvkYoRyNkNw
/bxDsDqWGxOyqp7uspQEbgXZo6TVU8ht8nA0bZcJJfZqWgXfoF2KvBT8dL//YVdl
VHheAw321nmDQu91eXtPJvEqSZCe3AbtmPW/UEGC39Pobb6GQiOEUSvUs22sR80W
AVL5W8zfdLV1n1jroCQa6jYfBZrbBOthJ2HVZ5Kh5e0yG3wj0gwEnDVP9qJKjD8n
eT9MpLxezZjgB+8bZkruvHBK53k9j9FXu5Vx9wG6BvJQGgiNN1JO6Vfhp9WO/KLO
FRXlLgftGc28dQ4BRk/ZfCv3SXak/jL4yHaoMJ4xxhXSmRVmLrF/F8GXUapu6qey
Zg+JfVbqbfm6S0QO0/1XuyDANo7IFsDptW2wiNibJ8uuOGA7c+njVahH4OF9ELJ6
JQiFkX3dLZ5FgTdQOUVhZsMZRKm+BM7omGtlI1AMowcnYe1HDXLXcv2udnBLW8gR
I3j5ERHsiCuWaqvUJl5PwTWuttPyZ0VsWNwnhWmLvtns8G1tRQNiYtU1BJ8Uh58e
QxeTtfT+T4NEQaQVXLOGBwBURVLbIWaEuOlXxMfXDsr/5vk2xLnZYAxZaqquBZYn
gTSjP0b8wYwbSr3e6dvZwZ6mkZdSyicVjfmZrGfSHNlppOhGrH3oBDmg7bPE8emC
WoXUpakc+C3BTqGL/ZFlWgZWMeqfcGkqSWfOVfG27B63aBGCv6UNBBtgbCZw8S8n
kw4Y68/wO8yj4gcBeDISOBpm1ZdHn7KgMh3ZUPYc3OoZ9G2jYuA8ztmDc28T+nQk
LQ9jsUt2fHvV/aFzbGrADmuHwo1XfD4Ew7l4VVhhjr0c4GD0NjxjMVdChIHW+lP9
poOLXRN7fChwGc/hTMw4o1hcJSoNEdeQEhG6FFlCrTistm5i82rZMTcUr7FeThxu
y/hMPceprCYKq6Z2VaiWCBMvTbbFckErQW6o3A6nXJy0Muu1eme7dALj/B1i07JH
LzKMtZ37QagRhIPTim+WCmPZN1GfM3jPPBy9gopFIc0nOOwuqSzoN5GhLZ6ZK1J8
L/Mill9qxZUFPlg7V/vLji0s49Vewc3Uc71I9Kbi+rjhQPDMclQSRvzvtSGJ1RpL
M+K7KZqOyv1viZ5At0/YIw==
`protect END_PROTECTED
