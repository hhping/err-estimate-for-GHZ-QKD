`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JV3QxhntAUsISzaEN/8c115yeUdr7jy6OLuI4WXSpn8KyOuWOqCO0zXm34/CK9r3
kz3gohdKW/fkNDxcSW8hqUtdp9RMqAINlEE3+0el04eK+ZWS+ctQORHljXX3cbms
vmrgXijR28HkLO7/d3pI4vitf8F4npGO+hzaY7JEKuzYQPRQkFEKaU1Ty5mqhnIb
gyp7Tk3mgYHgQMz4uquz7qMK+yQ3MeTQCioWNkaS2/d+eD+JhpSi/PVmX2fP7FNd
PJ8AL7kiOGSBaYdoSNuqaau6mFY6yMmz8/Zh01oAQInZ0+wTdbjRY/swjE1lICNU
FrTTdPbV9hzlToyYLRnfHNemDTeq77f3TUdwVkme/oweYL8zGjTAyX1V7Werda/Q
q3D5cOPsd/ZPcx7pyRCOxFfvH3SUCd6v3Fq3L6jvY1IyTWq8JOtGaTKOLt5bNl6t
ab/zqY+cfsBQZQhN7PRI7SoxjxZ92LGKwY3U5jRVfflRSHSifuo20RXGKrwCfWt4
xmOvgXmX9uAmwfAKIFBYpNLDR8ReY9Wk4ZxD/KjTw6R1Tj0jvjWUMLWf2FImbyWU
ZKhHuaCyy2+X75fk7PJvppWriBK+12dE/bahmoAYpn1SR94x8GPVDESefLxDfv4M
UTfen86H7IhwIMZ0qmF2tuXMixXtwdOy6iFyTUN1+Fb62itO5K8o14LPuBQxTMZ4
+vwdbiTDUnGHMFqvUwVfFMw4UA7YtMjsnB+jTpo8044vqpcGt7oMWGQaK9eiSbuV
L29TRgVrwlJXmIgbmrpTV9NUwezwtLP46Y7b18SsFSy5EWZFcWUl5NCRjRT9mVaS
ahAuLvVOfmh+EQedeC3oJQ6O0642Zcqz47kDXv2+9+4SKZBfssYSg4o7C+SGsA1G
oYFg+A9QHOCUa9/kJQBsmKOu+0pH2lUfRXCOY6Rgnwx/Rw0R3KDNgOXWaOnzQjs/
p2RiysoCoLbqwrvrNdGy+M75jr2zYXUZIHwfQm4HOs2Gmyyf4oKsJr+/RFyhEZoO
`protect END_PROTECTED
