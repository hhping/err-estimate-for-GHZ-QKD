`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KhHdf6aqs/gQ3Zag5tdCk13OrdU+Ak+oe4SdNYsmacB/81tkQoZmVotV16nrCW5h
Qh/cXU6AP4eNsGLzdKCLHh3oXOjsIvW8rHyO0M3M9zlPafdvsN4z7PiEkRzONzW9
YrnZKq/9BT5GYhAh7+Qmz7x0vqip33C7/QugVnYvPYXnv152jyexwDC8zRdIE9qp
6P+0TR9N+kYHjuLjj70vllL6SLgPfFf4/CAf7SU/nPY5MZ1PCxBah6SOzlildXJX
QkxkHlxe9IasLfmLlRbnQzF/JEErbs0UmgFdf1yXG/pWTOMpr8KHv/WGJqcEblkE
e+cYZ6lvgPkKObS+kBqAzG/QpUBiu5+lqH/Hwzqp7O9eW6D9a2Ft3U04dWtYrTuB
P94jQCMm+Zzqp4aV0gya4vgGOkuqXy8RR/Tq+HhnUOq8ye7A/anBRl1HSCUccddH
qo4pc2ChrFxzLAb48iFfP56zvS0AmPDHUZ/DdwJiFcIf/Kkupwr6CelpFppGyozf
t/8UJQWdLurEdmMEUD9hOP4dejLXK+XCeRdNd9svdAZfHOABzOOQXE+lTscOltbt
YE3dDSGDpvv3xjvaR2UL6bL1qx1XEMIbva0HI+DGbYYfYstUS7poh8FE0OUvtwO+
9Iwmhr6pDLomShcnULYgY6La1wfu3GZ8mAXlJU9sAduAyyxu0cmNhQ/sDOn3E2Ah
RofWVjVUafxUluuH2ekpISd1aGb7pjZu+gZNL1/c4QGYi7duJefRAchS6/mdG5Ql
wgDvmaSTCBiN6rDQiNosrPY71eCyNDh9oNxGNManGzQaYSwh87PSU/Wd4+EHayBm
AW69raCvdln7chfmhTsEl67kWokY+jYGSsTwdhzMttT2OESZHTP796BWuWysnsv7
88ZHYmrk0eEM0aOzGd2U7ZwPF4aG8TqYuX2WQLT7EPoA8+NO9MJDMtwP2oqRPIUw
bju7Iyu4XeUQpF4KYUsqOQ+VQUYFuI47B0ZvqtrpvrxYG7Nbl7451RrcUt+cfFzW
r83/JHRL0fBeVwLdpTWG5g==
`protect END_PROTECTED
