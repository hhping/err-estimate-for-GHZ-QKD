`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2EQQ9eQTV+V4KFE4oeFWbOeni1NFpLISiKUAs18scwH9MrDthecCJbf4L+UIQjgm
8TWd/+k6YJcpfquDazZBBMoXQ+7bB1Uw5mKjvOPoPu79Rn91nsPdn/wreeNM0eZ0
Dd6MyxRXxdspRBTXaJpmBSlbzH1at0nxKQg6NSgUAftZInA888+o4gv5dzSn8MTE
bXxcoNQ/rEtuizb1oRwpAjuTCpqJJ7fIWP+cGu0wdZDipgawYPJ0XG6pb/OMas9C
cuTlGyjVoPBae1jTOzLfuqnt55+ery3RA+5T7lzWSZN/ZshQv71ma0lIA1LuGloT
VDLr5lWy6SRVpyNnkJXcVlgDzunjV5Yf+SnocQCH8uPpOymRuGxoXVQZwtJd79fA
hJUq9Xsq6n3MmrJeZxvIF8VLDrxtuay45+iebizR5l9jIHuw4eKTVB3luBGci9H8
MFTEB8la3FoBaF4ue1a7gsMv/ck1OETqq9nsPRh31xUkwbg/Y6Hy+lVzUw2SdF/1
RRUh2UFYiznLbB0bxjTHHA==
`protect END_PROTECTED
