`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CgNqKHxrBi+L86ifKkMH8mnSTlcVtq3n3tEmTBE7HpgEMdkMNpvf3qdtdAzieQr+
We3huCZ1pfNEzi16dUdCKN+YYNL+VX98CVir6xfoeYd+omD3Hqgngygns3NjBLR3
5UUMbEgilHCCp3wNC0pBXwHo8tAohVlt60TScn6jtiirb2MgW+P72Fk9ZJVmaAw3
atEpddFGdcSJCBgXo50CcoMjjM08sM/R69x3RGX8VnIwAZ73ahdOloBY6wJB87rN
fxh9xi8y4NNrUx3ejhCgGtRe+9r/f95oz8kKDRGKEAtEfLITVChSqdVeWOpyOR9e
U0epDdan0QTBM4XyzRUUfBsEaMqeZI18es7b9vlWL2uVINcZ/ZjvotXq1Npyc2p1
nNg47XfAroAcfITLWahQjSmjp02JeaUotzgdBgbwDVBZ81euyAya48wl9a9Pjppl
akR+/wBd7yTfuj27BpVp1RgfMgV5w9R7YKOjLeR+F8eAGGu6HOiLO1kz+UTp572+
guNylEf7p4+9xOwhH7P2iPfGofS4VRXNns+fA0tLF58FSOChB/qPihGswWVORMTy
s20xobjCtrFjNjSByz8JuW3G4JACQiKpvUZl7yK4o0na9yb/JmyB3VzzedaSefTP
SASr8tqMVaoZTzjEYHOTVfMlzNCKoM9XvNE9HLc8JhKt+cruoQdwFXVkstz0YMgn
1/LTQ92kiJcR4AdUsoSgmH2llWWaZ/HjnGvnYX3mUfEoGBITqDhyXGn0Dk+7oTNh
52AiLWOgsIFre/Jed1Bc6MOLJgPIuN0ynymNn161lIHGGCgFllArYszG2IzIKidc
OR6uQ6lclbzImmX9PmXniA==
`protect END_PROTECTED
