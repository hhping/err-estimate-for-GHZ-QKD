`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mNPn6xlRfch/GJZtUB3phPZp4enFpHvCx3vKE/IX8KIDkcAkIkCz++8qw3jOAfKh
6lztDYHmBn505YA0CuqPDXjidreVE/bHta2BXycqw/JExiP4Q8p1uy+otD4D4GoS
oedF/sUoWpHC6Bt/RGbMswkYDOkhEjb1r5sKtwaTR96I3Af6j0yesr7+nXWpNkY1
0iJwi0F7jljXvo1ggtEvh6BOkZ8EPbId9vuY9Jtev7jNJSG5HmWCxKPmWZvqjFAi
JlZC4i1JNV+QAWQ5/o7VJS1A80XiNnlVJ6znVib82BhXQZktS4LgS2A0Sv7Xsecv
idG3e/QDggIxdBUTWtSx4E4r/ZV+JkEBwNp1NutQrb7tuYum5SxH/t+D151B0z0u
KnCND71n6WvL37spmQ2qgvEwlAP/tELssUzudBjPLJE9kQ/KZn2htl5z9OqPRF4w
UvFhMeCu4FLaS/ADXISvqLOD7m+XHzQuqzsqRnoqEQeNOKliwGS01yoTf3AObuS6
7wGN9E0qLAppemmhx4SjTscBMTzXpMqEVV/xoBgKfVAZW5I9i4HAEmPa5mSx0ZIH
8T8m4m0WAkRvif1ixVy3bShaN5m3+R3ljGJY5nNhailI4tKLzuKt9v9zDHuk4CmI
lxBvi/ZSLSNwglhDbQ7ljCxDy3y7UJWaPXsA7gdrApDC5XkDRhTVP1S78riG3u99
Wg25STjOE/1lzo45Ut/mqRGpyLHkXaE0YeDzaWLmIF0kHxSnjdIc8a5iBBhiqmEL
uD78BvmoV+2zNjDp8TR1o++O0N7QixSpZ4McSoBtUG1bGZzyR5JAM3E9Qj2214uT
f+4jDlH9oeKvFDMAGvndS7DsKaMO9dJTj2C5Ct+Ip//p0A9qxD8gWkRT52/QuC3A
Vv55a4hBUJlqjelSh6oysaMCW9OPXEJV5usaTAroyX7qLvyF4vj5YBwll3N1o1kB
5GGNga7fFiRmZiCtoOk7ZLj2ScJ4MrYz7VEUdw0DttJfyf73M2n1edIgbrahUuel
edZ1OU2XrOkYWENsQzizE2WOPKpEtHR1KSFyemjgOZFuTR4oNAG9WZI+WPlbQTdA
6D+kZhuGMhmLxIkoUHnSLKmD5qoxTclOiwTjusaT4agNbGz/0koytW0WKkt7AmoR
xUpKyaRR61RwZMvcF29m7eRv7AbvJgAgcCyJkDGkKNOQj/eHeI78/ITccVy/RlN8
3zOZGPqRcnRfkL2y69HbOIItW1A4NEJEAM6CRLRCk7FPL6lQ0OhoDWZu79GHI8fM
O7hYevXWf3jIOaDIROc/CQrO3ipCykvFt7Mi6utW129vguXgpzj+CXdqBHA2zN0n
zLniIejZ4PibYBrJLlUv/BZlDe2P2em8PbBrgNmcY6cQETl36ps7BISRcuXkRq3p
zALDkHNBDUDDPxNPHn2VXUgNCiOrY0HhNg5a/1MZ66+zZ1CvLjL91sPvfMvbmcRh
XhydKoCaEQo6jEVnRhte17qkyryq9suQ+HhK5Jv8sM4hqt+iDJgFziB5hi6yBFI8
cMdw3vJM5290iQFyfmN5GThOBnwDu+dwdLZDYvDNNU85BP7IxtcN4yrKyX2BaFej
aBdz5G9nUfEEFXwgg5o5RSxQAFNkSFRLXnUHsJgxo8wOeKU1ztThI7/5+PQZDZa8
EjyzQrr1Tq464SHPWzUHmEseaTAJN1DGRI+/HwxYMJMUYGiuiXRCJmy+KdggRdwa
/cxZblOjPymzsAtN3m4xVUVh8OMKYI0AmXvgaOejlnXKBIxcKoUBUnzYPopMIdfN
u5yC+PMr98yzt/E33bXOB6cdUZF9LW7uyXDUKdECUQbW3oqj0cTOfZ3TJbq0SEeE
grqxSs3FWR9zb8Orw9JIeKqllY6TrPqM3RaKpPG0Vh+X85HlSxqYprlrAiWyfFIz
RaNOFD5EzwBr49nI2ZNjm7R43ZCSrZlUrCdAMBcM7f8WLLGYg8NTpeDCLwyptTyG
7DImWCPu13pqTwvK1GK+3N8Y30ytOqolzWjsIGtI+YC3/UWT1Ifv849WULMNzjQr
NkENErLMSOnyVL8gyNPV+i+q3oya4uUA6/fj77LvSFAocavToyLo7k+1gZspydiy
66TuCCENuNqoYsURDN/cTp/7Y4oRu/ZOcKMdcqHXFQj5nDzrIZ8eoMclNhpIt4Gk
pn9XPKr2xIF8wJNHcZ/WzOhRMMFerYYuWFltf8L8VMzwrQXNhzb7v/2Z9KF0Q6/s
aXdX4GWM6pA4rYAZq5oJtD5pjDB+Y7AdgEMbczMRAomhKmCf/1BCz84t/dFwTxSj
JOHyu6alnHEtHqIxNquQ/4O4twRb9NMblRkIYzToMdFwoG2g6PpB02+imnxIA43a
+khMC4P+lwj7UYnD5bjh0gdgLpL6ZZDZItL1kW4HFS4+LW+jKI3/4kbXAsJNiF3c
kpssG+efQxq7e2GpDTsSGAXXpHOZIQqbeNZxAtpnz0XzvOFwX/nX2rD/I5ImFmhH
bQIekyko5xrWHPHKUqy0kBdka/9UApG+NTsdvWn/4iGLkXWv084J9bqhDsaoL/Sn
due8YaKIZYWlg4er2n9BCW0IwyMk/CuOp2syeUAs/CWvAeKtZySsf8IbvTar6aS8
XofVu3ZQOccCDlh5XFr+pj44M6tj+/0IV1MO8DvbL2X/VbF4C7TVcyeFxhpXZLKf
Iw4kVcPw5HhIVvxTjACJHZFZco8oVv8sO3pZKI+c63iRPH/CK/Nf7NbEdIqiILtw
k9zuAAU3vqrnQudKxn6JuteAO0SXGSfU4gmUm5JBqPOoTijhyBo/l2GSBLa3x+K8
Hqci3mGotrdRZc00KwrRo1S4v5iq94/O+M+ZdSElSs9ysuGQ212uSmYOkBHcGmDI
VQ2mdB89/AB2izbRS/EwGV0BPxSX2XnU0l1j+4Bj2qRBQG5RN2htRyBszNMl9iAb
TgUSR6afn6bA4iDMK6S56IoeeaVuLSLNNlAYN/1CdC5RUKBXrrWlB5IhOkeqWi+3
iy05Gsa9SNgHU08ZgXKRyReDIK40W9qi+kMF3ghOp3nnfB5zgJ2GYRWjMmPcjb+u
gqh9yHj2GmjOEO6W3bB/8xrNYE5A0v3vSoRu9ccq0UHoMvCLGGS7w7kbxmxS0wVC
mxbBouwCVQNpcMWssck470pZUZ/prjDjms7bQlnED5n9XcR7S4M1KVbS+gGbAa25
XtI4bVHPr+9iShM76OYfaQ90lP86LC5xZ1ps0PNqG/NWMWog9HMEHoId75UVxylm
cez+NQInNKBMHiupNJ82hdTHcj5QKodiHF3v0PFxWl2Y1Lt31Jcld56JSMSTvZEm
mCdrRddiP2evieU1JhzAmEowXh7WOoWl+R5RHKQ3bl/dpQbwFsc4y/XpJw4fb0IV
XqfyM351STE0t1UfoDFemeXbsl3JCnspcd8vK6HkU/uSy6xSV37Q6BrUEZbIhSh8
CDKQlMUWtwKLckHKP4QP+eBtyIUcbdDJMySDI6ft2vpOlMAZwFDM3CPkXFNlO9B7
7cf2XnUVHj6/cr0Q+IluvUu076T4uHbpTVJnvFs67mU0YvTBRxvSNs/VDpznsQiR
1hyYT05sWJxTSz5W8wWOxXTWB0f0dRlwaTDbJyH6/yLoqvITyexD00rTJUTGRjuh
RBWtaPvMDLUECWAiH0ZWVtXnZrpNKTWWj9or1+EJgFL2XhzCmyquyPrhh2ZVh4OZ
NvMvCaMPINPsqaznLrTB/TIzNc8Grla0iA1PI2Pgn3HpdDVeOAjCVR7tHIWuLAiF
I2uywVIVwV5C6MfQh8AdteOvh+K0pgMcnlru0ZajONU31B6cJR9QOhn7zbgz8za4
s6TQheU0ZTVHTAqG8GgyMf1l81Py01VxXd85x89J2P16TvweFavWaPntzElQhe3p
ZZ3xVSinS9AiB16jMJ9uGqQ3O6JAEgI9HacJPNM0J9hf96hEIrAQmqVO89ZV6mTF
nx6dK0/oe0ah5CnhLVhoJD6sxIcXS1RoFwf4JsOjm4t+83vB9+3pf+Zii3YPG6Bb
fDweclxArXqmpOrLJSvlbqS1PlJlV+3P0VnntYH0nI5j/aRFS7lD+BGs73gmBbwm
Ui5xtHzPsowvghpJUnPHK9HA6CWJFMOztNFEd+6GF3sbkc1fMoILMbpMbbEHOmzi
jPkDS8HU7OtxOi78C6+1mGmbiz4C1E5ezMUwRc6eaiGaJ1DFEvv5WR828KsKJVah
ujUsuJ1KMwv79qZ+NscXaMkB780vgRDZu+JeRGiruSc9zwSNaOKhJV2ytspWvvZp
FHYxywXEJFXTTTv007HUNvWwX5ucDnbaI2w3lDqlYOR+SAEL+JE7LMdUgfJTOWYH
yTTwjH2cXWR5uo79vkVagSm8MlUlC2UhNkD3QLDY9mXDOzywhnyWWJ7fCWG+6w13
xdTZ2yb/pzrbBvvEpaYa77WJLVZaEfKrQBRPSuDI1LkGVwIKnLXwFGU/UX53rTBy
hWvCixLZzoL0h6ytoUhUdKgzhCHv/NjLEpmLlfATcXFp8fjLgsRKumPouy95EXpm
3lFuYSu2L4bH8khEt6cvlT8mkoeDHSQgpQo4OA8r8pacJ6Ehd92u4nxGfOuzdz4S
3iVLig6wMY2hNt6xNk7PIeO7L/BgQXh0BJxhQKDNpyGtrIIEOvWoH6t+JUxFdTvs
aCXHMYHDmFJA5fJ6AcdCJsRwtDgRvR8hPL6iiXXsRl42wgqzDiWPwixW0gzRV3hv
VT4G379doI2bKOGTx6dzWnaIdNjUzpg8lSwGiEAw5Wjag20WHfH6qaTMoZd9tiiL
P5j4hoJO5qSk6JmzBGOYKjztRo0MK8neQ3O5pHp6OIYZSzP/kEV8CFnRTB+s/UKz
+bo/rJmU/m6QZN5eJc9mqTdg1xe5+CrJJg08qaLr8dOUm1rBZqLQPICsfQ1LcSr2
f/AhIUCdLdZfCKW5WPC8wZ2zQWm199TWxrAfplW+hUZGloTkIc47eI4z/swFWEkO
n7PdAbyoAvNNthIq/Xngx7YlWRhPg1N8f03VhcCPVBwS/mxdO+HCw9A9KBO9Ynox
2Z3mogI+Xhqc75V5WVSg8mappJY+Kfxwcc3iPhOcCy7+gq00ZC6zrkzJ4cyPL9VM
u6Sga3CzmXdMLrNdUOK56JAKoOT1h9gHsY1slVJOnQNZJ6BhCiQHElpE0+B/k81h
0NsNxai208KaEINl2cezRTiPoDojyRd7O5dcgUQftZd3FMnqAxUN9Jt3y7OuxW2x
KaaHrj7riFg5z+L4AKK5JhsjYZJvjgXsAfQSUhpGmwuaZ/DDYgAI1VA7D8pNmGtQ
0dCTLVVtrIH71ZvikSLB4U8Ec8/wHDlm7FICBLu0RfmIZBI62IMgKQwwVIFC5Dpz
TkkYWqvbHnRwfKsFwCl7vfXkScNMJwveG9vDVN5OiIL9mf2lhepnV3fTUs6VqseT
xDSV4ncVrmbpbB5x/T5ts95GyLTemNpTr8Z/DwQty7aMmF0udAlWPVNaIWEx2rb7
vlsmjs9Exl3KdJSMZPmClHgTvsowg176Z2clYzK7r8JP+sJMPqnWWzt0UDmFqH1x
8omtHMEILr4zmMwhfHESgpMLgSKpFQ1jh5iZWzVHesA=
`protect END_PROTECTED
