`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l15F+xzjWD4T4B7l8TkJSIk/1L3MmXJa7QrIKy9Q6O7lFCxtAejJnz3WUbJGUJ4/
+j0xdGg1nw0FWByQV8oeqKcYLsnfWwu7nMIA78NwGaDC6QsfE1VVtA2otCgtlRDk
Vg/yc6NslG4UTlMjfpL5FduYoc/47diEzJtnyQLrtfpkaUvJqhIH6U3WdWqVfAfT
rxfqxdR9np7R1iCoF4yUTmCoA2hKonReG+ebpns/Inv810CfsPwwbF6nX+6YKmJM
Ac148o0whx4LCdfa3u5fzY4ZFkTQnOLUKkU2pplvr6R01WHylpx3jFD84kN8QILh
71x+AczK2v9cPQFneUjzesjzYgBNroSPQ4fOGLmaz78MX9UcCFcVC2x3FiBC74tZ
lfZBwk+oao3kCLYr907HcT19WLOSenGJCv+RhXXRnNz7SnEPSCaH8JfD5/wXhM3R
2E+etngK4R+XGJ2lRWGwAs+tnbxu0iODct1+iuDq/uZPdX7U3WGT61HmIPLThTgV
rGkwz7ymhUqir2sFQlHPnPGnl81foRwN3FtzBXWXPtKbU7D2WWg9xZBGSZuY2BgQ
2uT9pyThuKRPSm8w0BVMqMeQfKjU7Gxs0KKgxIFvRu5R0BnbVsADVw44QofUIOzD
kusOBujsJDPdsyooXOBbWEZS0XXKAKDd81DkLZXCQXFr1vZXlNzll6fKmzF+uGH4
Wg0cjI5dEdHHKFiY45nC8E9N6qLdVqPOzQiIZ198irf3snpMdMJ5gFieVsSirKYZ
0f9cQRrIQ4yV2VrltGIvrqM2RjMOtUV23UO22V2Doke2+ofI9KnOr7q5dbUn5gTh
1VcQn+Rq/1TrC/t6P4MqXB3VSCAhO5pEKQAi8FqBX2nYwNShu74h9DQAMJow3djZ
IdbmMHsAiAd0rVMR+70oO7nFTzLTpFAtS7EsK8fHNJEJ1ZfhMcuyAUZkJhpp2X7X
BTOpKo4WtVZhZvXQhvTpdzq/sA03RoITCCskFHbotcL5xJtXK0jYkjAZ0PKElEfK
U/+CaLDGKduUqf/hqRLD5qLHTUWoiCS4GAYsIzet9/pKNCyZ3qhfZ0EHghZakDX0
znBSq5pYmoq2EtJyPT9zZyQHWhQVLtlV4YFjr29qIuGhwobJfrR+eRbTuXc6stQh
gjwfJjvzHVJMfAGT7FQY0bpMGU3zq8nuXRbgge6ojOnsZ1NX6wmeJZ7OJ/ULOym4
TKzrIqiV4XhK66bJzkGKcZJVB2AyMS8WrFItph4UldsPb3weyrYGBqvJiqaYntcD
L2mA7r4mQXip5DVtHKdsNQ==
`protect END_PROTECTED
