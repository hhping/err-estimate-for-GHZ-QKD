`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M38yd6I36LQPS4TIBd0WfMFKY+Ry7ekgodMDe2ZPXsibZfRhu6Mf4/ZcrDudODYY
tcW+3DG9Ygb3+rLm57o5gTCtFZ1jJcW4yTmM4HUFZZhuCzeG/5wQ/USJKKlVA5wY
P2YfH+IBewau2ulaS0ix8O7XIybHW8IEMt0UdXvZjCwmqIgAnO/FDBDZeJmf5SDy
VzUhluNzW3avFs5/vl8XZhQZ3byc/nwEMx3BxCKlIcpAqY2XOErQhUBwHrvXAJYV
5ZQNdua/DDAsRAZLsEa+cPRKMv2Ky3sxegJKzc5GSyx+KPNhx2sUWtE0nrvNs+mT
vzkZ7SIvEGnE5lDwAHYqu5ip/iuM5IidZsOFY8lX+P4=
`protect END_PROTECTED
