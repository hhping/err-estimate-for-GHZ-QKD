`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mkuwWhEJeQARbn4T9QhTnV3R0kmYvtcVOYCIwp5D6ZrOWda2E7ad+3lXEdU27XG8
LjM6vLosH8upJ3gg1RbvMCJ8mtE4KCEqyZpdzX4pFYqsVMjTy/c8IPmLgJvfchte
ot19F+3zpgccLE5i/FqNfC1Nce5g/QNeIttRNhglS9bg8D0U7nMkxef1mnFsUuuZ
RfdfLIXOd/PdtqppgcL9Do61DiBl3+ehVkT0zT1Ql1vM0Mryef5bs+zNFVUfnuFa
Jrxyx8exK40WuGkmDvTCeVlUH5NYGlS9rdcotYeHhnKnUoiNEnNUv2NHZuxPH2m/
YSocr7tTDEisPSMeDHRCMu1HOR1EGhqK5QEm2xRi+y7zcDKxRy3OuOH2tx2eXrRo
Rr4MpqazzSMrhi4maHeLuUOFZyjJDIR3kcuGHYrsr4d7eE/5SQF6HZl6PqVIi6oY
4ZFohl7N4MZle5zSsFBzpdkvWq/Sx6kcUe5HTRMPuc+u3/sVWu09W+6qQgeSfAuz
PiOiD2ARV7YtELhEu3gcLnS8s9AUJbXVRdm/lSTLsVpTaiNm3Gcl2k9dM/+to4RF
L3DG59YJ1Fkn00sFk+UpTCifmoFZfLQlmt8ppsEu46/eS3omtsqFsUzXmZisTuDU
opyPnuKQptWmwnv2X3oa+t/xtxdtWFYFXGU1FDZtCNhx/e9K3tT4C1urySsqGPzo
UVd3y5ji6AyWQyrYF3eo0TU7Z4Rhxfn5UFf4Cc7/accF467CcY9osHNYo4FaoRAW
RynC1yYOTgvPvZSrdV37PcjlfHyljTyYcMbBS/Ofak75WockCZnwIqDGLvRCz9xm
C44vEDbyd7L2zWOylEdHxtaiRD1iNdjrKkPGFKNwDbseWOVXp2+yrLanBtbMiqiP
FLrqHuSeICJChhgaunP//UkY1zIGEpzed4xExVbKCS2bSDZSkDE0a58UsFvUi6+p
gaExeOPnd0Go/PLfXZlr7jb9J1WuTlpytHDHRwGKb7G/W6FjahRHMRQravrGNrlI
vrBy+ykNwvFMyyOKbj5H+b77uRcG3hEhfPMVnIgesLt/SRd3D310iYlf41CSNsUE
sW1l03ROZWLSwGx0WiTJlzD5pDaCdGKEYcC68iyEWB3Azl/XjCM9bUxHZ5h/mWKg
TXNeIgPX1RrXX2kozZKTUYN7DMZAxe+034L7d5zBVbo2lORrFs7bwGs/XlESdnTJ
LVCrmbuhBa8MRIlLOHLz5ObRz7O4HkBeA+ilQzlxLqME+XnZJWfhhxX9oOlwbPwZ
qWV1hUAGk2QG67E6wOoEKpC4cthYLVzTEJz7z9jm44U0/9Tty75v4rCJEjoV+jNK
l6WYMUNwsMNgXcnREZH0kP1F1aCkKwWlH/xYy9fFC/wnuNxUfRQk3mNhJIbWt89h
7tEb025Zfl9HoRGgI8lo4kxL8/LyCGQR2ER48fnhP6We9dmg4hJnz0t1n/pN392e
URfXgISMqx0IdYu+L3VAdgiTsVTwwir9YPEbOZulNSynKTk7FgBKpntpyHAsKcuP
VnSiEA88WWvw6B3Utt3eJymPA9m1dqUqQ6ArN+1ZA+CzteZRbUuHIUH63FYmCNY9
X2YGIsuPBYskRS3wgwCmcoG5F6Eb3DdjnAFWFUx1nxr2TB9F7QNlLbMZ0Wxg31eX
3tSI3wHIy/dtfchVnC2pr2TeuJy6m80+HXC8k4QXjgCkWIYHySvAaDMSlMKrinPx
/3Q0i2fdFK4MBn/m8dGOp7w14p1l34w86ej3Yk68S164w9E03v4ooODpmuCOSTDa
ALgBLOwUo4lY4PdZO6KXovRqoWc1bKDBm2dPNz3vMVfSLY3JHyZ84a8pc9g+M4ik
z0nscEKo8jWTfdgtVXbZS/Swxxd8omPNARDe2PgGqhXgL8KikRbSYImKS9vG7Qn8
e12Jl8j4JSZVEOGT46o0aZGuvl82xSj9YmeAy+++c0M+47o9olIf59dVKRH+I7aw
3NiBXfhrWzflV+yKT0q7X9wX1rmYsSavO8YipV/EmTcboybvT6v95v9mOwuY/6TH
K2ECT1ZR8GlCSHHjUhqWeen3NHEIPcZh1h+A00DW3puX3GWv82l3//oP732mcgqT
Ovf5BoUWqgQQBeoRWq4Nvb0vlmII4QYBFfgHeLcKzovSJs8teOMGKH8vQtAq2lRw
ol3zMSD/wO5cWVNwahKsbIWUVETLdREgBZP+AUrezT0O4bVxHumZKIu0zW66Cfd+
NnlQju6KfGFKCbQQ5CCBmwj1jl9cZVBBKgQy5ZCxQx6plQclXywrw/Pfo5L0vvzs
9aYYsCXRSTzXQ6HXYeMqWBVGD89q6Y66FnFSSMEX+TdLtg7UNxaLQ61p43MalzgL
bzWvaamhOst/YJqBIkp8o/tpgel54OuIzVWk188pwhD/+mXiNCdtgCCamuoydnS6
yt0pViDMaBcjbpxBDaRrfOQFxxZNMlRFKa6jTLbWMVUqcalrYt9XV/+HLy+qUjQp
8A1bzgIdz/qcvpwkZkKQAmG1/TO5ffV0nEiH5rWhgrwIIQTkgAUuU3Ax6MRAV38a
RYLHnMi7s72RFXf4FsNVgYecmhH34BjRmOQvAW5nui55YOanrwAihm8pDnEN3NZ9
KE/66Ix0l9JIXtvHWQKHLil3PzrnlUp+cx8txfYbXD1ZOxMqxLROhb/F+qE22AyR
RF+lj3xfYhQX36CO1GB94MguDxBaJy+9z8nGt/aC9FEig2cc7GGFNkJkONgHBM7I
SR9xnCYblCCgcgvPdedEQKA7DaaqR4+c4pFVLS0GczE9pKu6b52nfVoVOhQ408we
WukzawciXMvj6uExGQnHrBpkF7pQ8XTdK6+nyTgsXmuj8EQMzZQIvZA1T0IFiTGp
G0oj338TbcC5ZL0URgvIXnw/hfGA+3dodlIdm4pd/RAfQa39X4tDF9mrqVHO35Us
yd86ZJ7sBxAwteZYkwrTgsvoIcuy48+3GbZEoTySn5UheGn3kKfxkwxab77e7AJR
d2qSjUxuEV6tZLEGHPpodNodXsEsrI5GYUzU26kDIIQjfro5LfTDu+SHcUjyP+6C
Sa708iseipAQ7CsHFNzUBA3CpSit9ygq0PD8eEJf+8xYQi7JNcRBDdDPslzqVoeZ
UU7zA+jVqIv1xTHw9CcmZfxeQpN/VQPm7OeLoNp1nUIqJbIK062CoGJJJWWB24g4
RB+gwF9Y+qywxZX6HmU06BfFEaDOLq05fdLbVDDwjm7GU8IwPA6MKNTG74V5qhzs
h5s8omfBJnTx5Xt7q1vVB0DrWVZw247rNHApTZis2rCSkFMIjw0+mIiDCgZFhSjL
rT0INS727eIT5FUH3X/dj0H8ICo4lLI90Aa9noMsYH6aQCZ+9OOh1Xzeey9/lsLS
JK84Vlg2jcrpzquCDSWUaHYXQi4at8hkzBeUEE6pjWw3EZ3qSueUX0ZNQJr6uOVm
KNvI/my+D2mbUlPthHMs8UKm/+SF7D7VO7LU7FdMEC+astychY6ZS0S4PgaiMzhH
qqxJiMhdGCvJarRPQXHVu9rb7O+YHY9gfInL7MVpgDY+H9pKX5FZSnCcHxmXAdlL
rBhY5gB2PBCCW+58ro1SeLUgLNDNutywKn2+YPO5ySszqNhkykGGidzCGZldVVYM
shiH6SZOFMaZ9mCgH5b7ekZagR9LnZCpJWtCxpDQuFOGpK+MIi2IE9AxNSqi+pM3
3hvhi/jj7EjRyCdoB8UbUxBJdRFo29KkONQ7Dto5bx7zP5qzG40oP7rxBE8AAygG
oVDvp1O6Oo74p+H8zEd6gDolwWZUFjJy6TMAeQeLsK1YdLl2qDLair7smt5+y9hU
weoVM/1l0rCsen8fJL+S1QAgR0pMoDbT9JsIKpRWeCbvtuRNkyXjbnAnICJyLQZS
3eL7vbdM/UEHLXiNp1U3qAARoxcad3kbSCDVQHMR0n0Bt8pDn3p+1pnufxaWpiQ9
LBPeWYEbXno1EKn/QcJemsH+clYMNq5xNSwyFyGWq3PH5+65CrNrd2zV/OlQus8k
8U15fisbrhHDeydM7CU4VSxM1UqnkMGBqWmTJyxjgTf3Dt7G8Qo5N4vGaVoSJFBB
Fmraj1R2k/OQ4OsUNzEFQRJ4r5fSRTZPV4IpsSbHSVsnnXcZc+6q3MQG1zERWUsu
fMfQ+Dx3xMRmVw0QHvVINWw5sEcuYdXqkFao0PSw7B6BU/HVCPt96dtsfSYLvpqO
BegYu2NzJ2pqafcE5qE0vLR+KGUtsdkuE/cEO2NGYUVFXZRZG8LHBT57EIRY8K5B
9dU0Nxj5b7xJbS/hyMJYw+Y/MndqdxFyGASbO4qjbxcLhQ2wQOKr8FSkfIuAwTTn
t5f6n/zwRfa+hWp6ddzKfTAKCVMrAc0O6ewV2xV5WjzDWb1xU1htv4F2w5cbuYuw
/v64dbHnpKh0WzbWGs5SvG8w8g72iT7oa5lnhZ9mG7UEDFOoayssmBLmREEBrSmu
IRm/6JE+S989T74cWxSIBBbATprYNkZB77tU72RX4eXieqnB9uEQZuQ/wnHCVMfJ
IrM9UJMCwoxaV3D6G4EGQGtmqCurfinyR2kS0CQdAOAjutq96u5Bi3lJoCZ7mfr2
yMuDrlIfCM3pa5o/J7QAmvmI45eHrnJ8S9qGTwpWbUThE35PdTivnzY7m16u0SWp
SOEhAHjYruq96ARsKkbIkuzZ1+URADRYKg0a3+/BzPz1Jsxn5HmiyCkBYfr/Axom
dzP9lgT6v/TyBY10DXRAyyjNTHZwEvjc+jYaUC33dyTZn7zZiksL82Bouvdygnal
lMVrxyxBxVtc7lg7CU+VZ1W0ac7FFi0AxHz8n/C4lMTgNdVXAo54PgJETeLw12rm
wQWJi4bKaMl5WJKwf4EOUUYYM8RWfZ2q/edweVXwLwRaqGub8efugp8fVOxToJFK
5a9Z7Mq5s29DGJbDY785tzAbXNY8mbpy4soRQB8vPp08Iydj6ioWU8YZccXQIGfc
hkRQmeFkrqu2JINkrg9Z7KiTekQfPulpiXeZKrevs69TWjWfFldqpSU4G1nEWcDP
6KQD2JWMyAhTmHLENDU7iLwcXtJUIz/u1uK+XTlETU698x+DhgB6uWhxGrqWVhsL
pMZ8cYbr3w15vIjDQu8Ns6NZgYWv7hXsZrxJavHlXNU6X3EadXax1D+38YoQf/Kv
bxDcw0DFj/TaZ+ZTFkgPxvJxzPHOAGIFZJlos02XY7aIHCNgw4bc4zbPsIjl2ZDq
dwYpO4CWC8D28UF7VpmzfoiZDf/0XvFI+rN7mk2sN1taf2zEs9IP8ilFKk0iOMEa
XDuTC25+1M31RqMECtx9RM1wpw3FAIrl5Y7LPGQwVdSt8PnhzEUITdwxvijhwK/6
4MLQJpNNooXPmT9KSl1uow2nPob4yVo5rQECmCoo4xuPAnljK4tek8Ochm7DbdI2
`protect END_PROTECTED
