`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gCi5jytOp1l1uiOSFbQA+yl9fQo8l56IyPVuxGxhnJI8BOXAD5riv6Re/XZ2Mc5s
FgU4PJFGyEA+Y7xemq+ycoAQM/+FjTd3vcRilIin3LhEHQZcUL8WmzouHhnoHoq7
ZX1Y6tqM+23CI8hueo2+TkxStyDDmeEA8Jv7MC3SI0BXEAnuN95ZdHoVNZePpwb8
2Gml9aP2FyTOHt/AGVIj+ZBkL+KzlQG54vAjYtGnONO0sskV+ieQck58Ns+0DD2C
v+Mk50t55zMV6PpnrRYAWTvNoec5Hg2QMhr8leZhHJjv6Fg3sxnZdbBz/gybkJPh
ebsxWMq7NOCg6Ly1eYYdn4lpYvwrEl4Q6u9sqymosplSIORiSrfxC9znI7UBXArc
jwr7HyH7T14fUVLFP/8OMhP8biowGk8tXVXoPSArK1/wQQ6OgvRBL2NShZsIC8ZO
E0YIsDa9uzrIq1O40oAryrJK8X114YMXkb375khadkGApZgZfRuUe59gA4YBCAcQ
TDGLWyhG5+pdfkSq9joeSquMhE4XRxmJTQb9e2vtcEZscVfEMgxlcgJ8FlIu9yAq
184OGRRbzABoGRSD/UMQ+oiiMRntkVG0snpbpz7cDJcMmB1EbhDOmR5YwxsmdYyB
MhOsivOuk/zb3HUpNYFBMa30JOfm8+crd8HMdlgp6N2LEE/tWrF3dFLvI+4pAI1+
PtClanRuYsoPBuQNU0RZ7AriglZO97z0BF7C5a+2oxsJUY4bz6kf6faPdTmf1Kw8
XhKNS5iLOkPDVsukqzc+6k6h50ren38jvvyQw0bmKC22+HzAxMtpxQVcsYgQJfmH
cc03Duro7zsgN3eUPWjtOjMjG7OIlxZfY2dM7oh/A/3yMV9NR/1Uak2l6KiebO0o
3ZH5Wi9dNeEHTlK7j8mfpVuC9LKsbobaUkWFUorL+REVkrU+TWskXRySl+2DiX0M
+DQEVfCAfaHx6UW1ebt9/xAxhVWhCTtyVrG5LGeNk0v2o8SWcpZ82ZcNynu4nsyr
dat+zH5JkRGcpP2frpv61QdRD7SEMCLkhNcktotujJh1jJhl3su4fgurEAOaAaoT
lj3xiDqukyFyam4EbotsYe74nFwf63WS1t2GeaHlOrxgZcv3MfqziVhcnnbWK+B+
UGL5MvQvCgsZpHImwHNUMWXoZAcPrFlwMBFfeItgcnxLHG7wYvXKDVXj/z7hWjoz
tOlzhIWfNHcY8ZftaIxiNwIC5trWOE/JuAKDKlV7hFKbGD6XcMlmFXmlCDR1tSOu
E+n5iKf9u1rSXqGLIoGOSGiTu5h22DfFD1zHPEQ6sh3pd63rp1swA3OtqkcvhSaA
I/yJq4heev0VNdaE5U+r/JVqdfzCry+8TzAIfQgvXeiY2/bBAsQBEq7a1N8W51ez
swUCP3weURMiARmo45+N+NAcAR2CeBliDXfRzUc83QkmSyBHsmc8vJgmwz7dPMKg
RaEMiJ5/ZnFFrSSti9+uMmWUo5ryE9TDoTNmqWZ0F/NCnaO4FA0DFN6q+1Iq8l70
0HXRp0Jdg9b4m39bEDUklo3wIlWfFUpwxqlDbQwpKOrV0VBu0I/fZRXXmt8uS/uT
2a0jTurBCaNOHULxW1H38cyovp6Q3ekFIBvTbKNtJpyL96e1FCZp7vVplxuCAUhu
dmZg2JgKu55PG3MSQqmjGhej4vu0m7AZgGeJsU5EhHslTw52j8zolUCno1gHoDXQ
2CA/5xDU9t9bxM3VZGsnDzks8pweRYBkhskougMmu2FU0Gi4UYFa/bRua7Pzo69r
gNdw0c7hhPyU7mzMO7Ts/bQKZu0Zv5bTipqthdv+Vhhvv4c06wNi7g7JNAQbk5we
DvaApaXjHQKubzDrWIjnoKnuENhz0eWJ11NQpLahacouG1eSc5c2DXdcYjMi1/Hd
dVgGLHDuGdiLRwTu7qqvlDINpv+IPGIr8sYLj2EKna2Qpid8gVw+1cI8x1fhMXd4
KV8D1kVXwPMQMeLfnYEyJvRDPQ6e2ZXMo7Ost6DNHEu/ZvfWJolZBat+XMeo+uYz
9h2j0yAgsDXAI6ZSK6XhBXgXpO4+NRkFWO0dK5dHZKUrujSchGaNjBgKgHZy4MUu
HdEIbqoLfXqFnKJ2RW08g5RkHvDzMIYvh2AqMeVzMprEVkjlwBUgYzAmZf4aaOtO
WEsCN0IBWtF7bkDJ4BwdP6wdNM4UdvgDUpDx55ofqJqkasj9XSgLdBDSIS39268f
jlNMdhFGViRG2WpHO6nGa9zlBuBMXC40j8Cc7M18TPPHdLSmiJxfTwkhK5S6cZqQ
hnIk1zBivVZWyZwLksg1d17tHrY8Uovkc5PivA10C7XFqtgoxd40prjYsjSP2/mx
XCLBLSHI9apyG4KVhm0LOokShAKmslGZ9XGZpVjbS/Ncyvd9cQxbvh2bU72YPHCZ
EcOmizRzZApRWfwCSpPpZVBvxfU0AYua+/TWDgKDMZVI0Bqn8EAeVuzH0GORwbV3
lKHUgS6JWIvTSpzffsaRyc9f2LyhEUolJTSHCqptnXaRNVkVBW6mARXi1LtdK0Am
ePMYQHUfnGSAi+67Aba/G/4c+RUmC0TLZqXoisClU1c6I8wbDgKW2t19OGTe9Ynr
u+1iPU6gc7G+j/EhT2CBVXowsWT7+Y/GFv4cFzfYxvCFTlc3J+lGsr/8/9VXvXH+
N09E/ewyJK6XCfMY4KHZSYUx19W5z3IOBMR1DRp5q3OjXibT9HxyNjVfySEDbvU5
Z0z+3mftddjxyQ8g+z/tUWDMkZMVqe3IEVpAvvQgJ45oCn34BT+FJDXpUMvVc/6+
3+uGLd2izRdhMxEWa4pRy/jlrozrymdftDGxijon+AJNYFJctAWqWlTvvumxepSn
csQ58Hk/oZRGrKdE58HqsGrI6Lv72r58ADN+dC3FTf51daLaHUAc5QsZDqkk0lkh
gDoFsA2LJAsmje78hJuXQqFm287xp5Cdh0CPqDmqCXAmBIoyB4/tfVE4Jb+8GziV
jOaSQshSMtTTfMRQPkSjWkmWNwPdSwDTOMOq63C5K6H9tWs6d2x4DcXeSSq1hbUh
04WDQAKEBFpyl/r6pVODnI5X8RPUUBbs383dWY+dAQhGai5alSPtqhglJTOMqMWi
BDsYW1eHgqAAtViT/W2L1BSCgZRJJ93LguPAHNFGOqzV8Z1ZqtFP3h+ImsMZ6K82
4pTbnRvbtoObJTKRV6P2aIJFH936MxNKY270pL2D1uCgb7wIhKGy6rENLMIeGHGr
UvoT5Xdjp3beGH1BUFXvYbaPyLjNg98D8sfFmw/POQX2TdxlVEgOJYebpSUFMkmE
AOzle8O8AcmlDDXDsfTiIzZb1mV4BHP4XJOloryNKHTMKLZ1VMY1hFFSIi6C+Yx0
MuYlQgSTl/eaawSUjH57okHN4siaTJNCC1TRP8qJmVoF+v/af8sa2uRBciiS3bww
DU2Ftrq2Dfz92Di5MM5RJHX6XHKKK4c8Wl+TaePcEn+e/QI7exfLnH/hlsLsvzn2
d0IH0lrQ94Xe2PEvZfXnbhvJxl67XdQgWMJuIwDVmeuLrBT8t2MIolNB2cYeLnRc
svelcYmw+8OVJD9z5ImQWDX5MBYHdBTuSCfgrRbN8jHJ1/w3vVNvN21PZawIO3Dm
IzDmk/BbJ7XVRz5qkWL3DS3dAHk4C/xJ+CYMpRSym8wvnUb2HcFz9NEeoWe4e3mo
7rVR3nm8vvmJGw4cyjevPlTtxRx1OH9aBltgDb/KMkwEQfYYzXBdCCOUkm0mJGMp
cDFCWoeqTxyHWQ8uUBvtuJw8ebLcbPR5idt170RlKcFEjBTOyt6+mMH45ZzxzpsP
5XQnanw/kKFDOhCHTvNIDHRJQyk8yI1rQqGfwBGWEt4OjSWLVz/RgqsPqoOGyNN8
Rx/nauZx7GZv4pgVRtQUZOwp1zzf8CkCfvsd4EFCgUH3KdOJjDiH6rj7l9CDHYgh
1L2t+EzSd0de2dKD1wxHQEf/b+OkQjCHLhMRq9jZSVMHyz6ITmPZfCKDS+O3Mrpd
hGMvhWJ/OTwn9j4QK5BsRtWiXTO5zyMjKX7Reu9Lw2RdTirFTXf9qVGivDidaJhS
kYHu5TwbtEKfm04Rg0L8kYX2QSdPbNxtrgsL6h/pwOP0QcodwGre+FDj3iXsWZOR
sPl0STW3ibSbogehdbmFzhBHmImXxFkzYgVVrT87eKdnDiKUp4TKgA6r3xM23uNX
/Jk21P8V+9RQKLOyj+13zVSLnc5cEiJd7B/pd/BIg0xPI6lDM41ga+VKUmaWoitu
ui2xx2659xnCrq/tt7DX6XZT75PSBoeGn0T7oyAmaxNX8x99ogK6bwU59AaBeN7k
6rLT9qX70/xnEvjoFqTWzTKD2FCW71sHzAOogcG5EFTDzHGBiJJLn7Eoam09pnh0
vjUGTUPVARLmM9Wn2pujKLJMJaycmKBnObJvPYA/a5fzj1mazz5GjdlaQ302DIf+
UNLbECQ00Dsmlm+MZPGHEfRPnGpP7xEOTaTclMyHgJdGqzVYxk6vuw2lg3tp57Me
5N6qRzMe0e33tffnx2Bu/loV7VqjZN5shpzzT3OcgO8TaNehtS8OR4pkxFEPzxn9
psWiayik74/VOcEKOPk/B3pTiT4qQ6fnaH5meuXy41A8Qg7+eAQL3AQMF7j7GN0H
CUDp5kRPtQeEhZ35wa3OKQ81BZ58xeztY9QMAX+MCe+Utp5HwpzrrH9E9R8my09B
rjiBG5G+gZqw/TowBER54OQmmIl8tBXp2N+7pknVLKMdVjvmnDy79469dj6YlMpE
4rYPhoEo4ANPE7z7YfGk9qkdvOa8P/2Z3DG4NvKkjPvVLjoMXpCr6TTBQaNRxjCV
Nwk0geXmsgusdgpidwddh2JheScXrzvxQ9yyI1S0BjAw18Fp9Z7rp3GPifCrM+ql
epyw/V4jS0TjvuDWFK9NVUjeQ43sCfPXRjk+gIfI06N44KWghPG4zC5Q5o/fSGc3
4QcJwNqQWvUM52A+1q8QefpjLOPrGIPvN9YNGnhpa2ipPUigpOLGuMTeoo+o07K8
NtFM+DKJ9FkMI5bOvfH0gmm1bn0mYRajBUj05PoPYDHccB0CYxEbblKQz1KA8x+H
jFktUJK3OR7/d9aKM8jH//EfFTbJe2Mxh28pRVbw2KwlMeayh07h9qQvrGsMUwYS
8OEhBrhOqwehLCDxMWozlQvCkUHbgMh3QPPowSshkQeEgzamSBeDe+eM3lXNMQ3G
JlzMTq5DASwP5yKBwfa2eBfhNkGFQlhf/OjFBH8gq+j32w1yVjadSgSk7NrYFiHU
gDAWG+WttaxsDLbJD8mb0Ey1Ym+bOFrhueyMcRscvPM9NuiFfhwXOhCMfOGT7siz
YCUWS2xGH330Q6i2jyH+wbAVpondHe3vzW5JqVypQPJrAuyXMJRVZwD1niwpFvr6
uKfIVnxf2OhyB+KLAvcbxlIRZcjzhMDrXlZilayI5q9+RKSutvtFAxU844O4ffc2
tEnTEytPrnIYPtJkAI8gWXEWSUhEkjOfnFl+UiOnChgvsMrtVnrnU+CZvIpsH+9S
7t4xpb8AyJQ6dptQbxIAzic37jjPBj3kB+/EiZRAJ8CazfdNxLtIBoQBp4CltLUZ
RvmsbyDFjnt3w8muODg6ojt9jW44GVSd4ayhfeX56d5zJ65josHOvBpwCbJGjaFM
0SrRh5Dc/vy7DP0GuCO7fnzsq0TNGDfbtG7fj2k9B60FURPa5WBcq/xHl5xo10JZ
Zk+6FPA0d7Q8lhpECWtF0OvpclN0Js7+T8aXoaBWirrtj5RrjTQO/yuJpY0RhBnm
GjHzPS1EQxv/xCqiV3/Btgimz1RtJO5gZD7r2+0UWzUZK4yraYip3R2aQfasU7R2
RIc1tvefHfJAmYsrGLYQufVpmnVydL2vdrjKnJ2/MVWPpeO412wGHnx53ko0bN5v
8gMO2lVrMdXAExzDmhCH0k0y/DoAx3wC8CJ0ekbTCsMEzGhkQ5qc9w646e2wrMDV
IEij9X4H6Et/rgXVvoTlqjvgSR9MmRWcGT4kkAJ/vglzyJtM44bAk1/safO3UfRx
TMqFzPEWtRLPBjCBiwfOjMWWXFK3i3YvVi4lFsUKzb6a7oW5cfDWiG/4ZZvCpPij
4OB4xo9fRedc1Ua8LnIUx+JmkBhEiBY6WaVZy1dBCi/jp6u06tttigrF8mrQkyDI
f/wb69fyoIM5Ma54iOhTbwf3rnuY20I023LsvG+avqE4pOFPlf9L+H2CUiSPhnKf
plHFX4X0VGhy5/JHhx4ShF7/wWugCfIa0J3ydQ8otXkYGuLbAfGmyQByVX4W5m89
Wfy/6EFMujek+JK3aCBoFu2duR4SHfQaDwCJf05/LByEYkfUOo7rRoIrLBaeBwGe
F5QbO1IpeD8w3Rs609KEXbceLcPFlgzXogQ3DtRX8H1z/1s0Jg17csXdzKotaiGk
KsUkueskBPQpP3BOpeed6w38k0GrUmOggY8Z29+lXSEy6DhnS4k2ICqMfDl2WXAA
oUQugPQdrXKTNo3txC8g2f1o+rr9oyUvslnd1qhraZ4YfCwmo1iOt1S1AbVEdIq7
QwTIQnhoTWGRD1LkelHBdg/ce/HFyk2qgTWLTN50KA0HdDcZ+d6ko7b4URbE/jz3
9KvS2xNxwqyQggemyFGpDLT8+6YnUiq4EHRMYm6HAadnK+5F/ks/RZM4e6gDGLwO
Z8UW/puQZsP5qd381pU0UAQ29Wmer5XyTmptm0Ma/LgVpbpMRC/7y6SZQ3J9f69J
fEUlISyvpy2TUbnImT6FE7aMFSxxRKyYuGRo6OMATib9zuVMWTLpZeRb3be2AIN6
875OHZG7O8Pt48H0azLjtjtmY++NY2TksruH9hU469fHIc0kpV8uVUc3hWKSVqeS
LtOTgaFLleqMZAT2Rj0+s90VgjeomNRHNZENt5Cd81+OGzam2Nx9w8SkOgZVh3ld
Ding9u5rdVAp3nuMglxLL4ABN4UMRO6UXOd8AGHCPQc2O5Ap5WsV8ATy+SztphWt
MV2F95yQJV9QJBglqZ2MEQbIA0wAtzKmHZOTQDjRuhjLZHPq0dY0xN+HPihk/XsA
JFdQrMOljAR8SB2r7rQUOr2FL0oxZ1pMGdaUHrmyLs7oF6QctK1037Ndnjea2GH3
HTam/dNnkNB6QNmI1p7pulWMOsDm4uOBchZguX+tsQfDPJGIHviv4yfnJ/aRvto3
Wu+QcvaypTQFVh3p8jvzNtAXVs7VZCdn3TQVT6cOu6/Ly1o9OF3NxHslvy3xzfXy
h+T8JTmKXjbQ5CyV7CQ7BZ21oz6fm4yUjmdfjaMWqbrDD8vEET15qw2UnKYMtC9e
Zh2Zek/1pr03YCQjLVx1XAJ4G/XbPQkbcCj6biDbAeR7Xcvl3rOzuUGnOS7ROHua
SLtUxa4Pr4UFyxnw8IqNLmUY7GBGt0sO0sQu+mS5u1eS/tx+djAUftZxgjhTuV/8
yc4ksPdBWNhL18Nags6kjFKz+l4maKhcCrW78JhH93E7FbTAUXgxcYP2YsfEK54o
EUT/pTU8b3PutN03woTuYWG1jTeH1FxcarZy/9VcswmkCxAtzYlt/i21DARIwmWv
zv1eb2kY4xGkA6Ykfe31uE1oesn2hOK+uFhe+8n5BsO6nznk16L9NTg9RhYQYOYm
PamsKbrzMRD+ZxdmIy9Ks19yXpuMsPuXV2an8p9JeI7HGybRRAtcdt08/i+41aCB
uWMVg2UtV4TN7gOWzOiV2/HlEa/YskQMggBAOToWUBGytfKAAOnf73DbMRpTGwIB
e6S68Ws/xavfAaf/vbUgolg+thjmk9UVMKHVFtWyqTbk7tFh4SLEO5FaDl8QIu7R
cttUUc7ggim0hk+C7oVfVKoePqqyn3JUZc/sRqUhaW/UlnSi5m2YxsEue8PhdeN+
rnbgI6vxTlwd5JC6TzPTd2EkhrTR3tQk6d8AaAzo5w3XS+YRUcThsNxaUOdhdseo
y+jNhw9u7YcJPpDz4g9IEluaSqhPXqgZvWMzB2TxUfHlA4LzixbtDpLV4Tk0MqXr
64w9zZLl9yWWWz3V/bltbzAHAqG6SPC5WLbs8tBfODVVsdOiowZo6P1r6mWdgf9T
NVNm1Yj78vSSjIwaCUS7FYhwvD+Zov56hZ95erYX0FA2bEx4AHV7Snhzf7wq4M8t
Qxhq+OpnTVJzTF9oTRB4y8aarrJ2dO2p2Pb8S6OY3DxjgsppxrQiPhhun25E/Izi
a/XiophfMs5L6aF+t4Vzcu7uo7WacU/EICahKYyk4rrK/X9Axgf+eShbAAPcB0N5
sJ55ETfNXHJZvokhkVIW5Vb5IlpHVy7CJZ6bc/9ryQ1m835LWnspB5ZDP5JFNmcx
o3tm8Kw/bQTXjF0XIPJCBkGGLBlliQZ+9FakCUHp9o05XwsTX6OqcIwL3GG3gcE6
oUGM6/Bc0xRFG0wBcT2vSkMmxL4Pc6C2R6ktqgx/I8grASy8jfJQBUITno2o3ABW
b1liMnG13jXyjJAm2h/flhUvrSr+HvDDjUQPhlaoxAnqkqgmk0DQrUNINs8HPn5G
BjIFiC7fs/DXTu1hXNgD0znwXOE3uE/h1nbQIX4p3ePPF8EUF0lSicgNabnA+mPf
CV40dBotB6/Wdh9Sa+GyjQAiaPPjCz7Iqyax1nt6TUL8CGJTDwWzdHw+crd+eyZC
smsmdBcgOzrN8lCkF4l67lVdLlZtYE7E6n+gcKzdZmC3n9mhsKLDY5tyPTBsx9Y9
swEufR7G2GCDt1BcbUpzBTFHRGwRtcjdP4sQDLm9VDM9GdljNLT1h9ocyBBzoC8b
6/MDQoyTk3G2wQQ7F5M4GSHy27yh/gMtG5JHr14O1J+iSXhRG5F9L2AVziJZuVgC
TPKf6AEY4aSSJQcpcwRwO8EVqyTp9Bmlkq1bdUM0IJvDJiXfhDs/eG3w7X+DaZo/
GEunYFomPFqPkhfpAL+S5F4jr5w4shRcz6qYzlLtGg6FIj6MFmxGX4+xRUG0SKPu
MYHuYriWxSpET23clGL9X2JrYDWJQmyPOCJQKTV0kzxjWaIjp6D/Kjrjx+czyHkL
DZT89jVuovK/bcE48xDnUGZdq3rJ3vQG+t0YrdZZUxuhrPqPPHt8VraRHGu8LM4O
sjRqbHFwsa1oWfi19rXvvUeUFVMiRxn3CenlAHvxPC7hNfR4Kl3Vt3yfwzfRV18F
Qwyj/85153AnFkkoet+/THKTwVYI63SHMnKA8YQWqng=
`protect END_PROTECTED
