`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6ZFxUtJg2UxRuzKzySooLon7WC6mN/PDWssmxhC7EVnRC8y2PEZ/HDgKgYpT501x
n2i4hDQY6RAMvBjhbZ7JOLmokWomBle9ftVMd6t/R43yLG25j9zIv6XQD3LKkU6f
bWs5vluRqjs4BO0rg+Z1HGVHTgi0rRaMvMM4yGPdWtkfcj7FiG2AqUvuTTpAX8S1
55cFKkHlq7WEx/HkSpZLx+hcFKlATUkaVw4kbBoVn0BW4e1JKy6bnD32smGyh72F
hL8uwOwkSRVy5AAIeDAWzbgrmUo75cvR/cAFnbZNSzUIxbzadyBfL0vYYnJPc7Oh
lKFYinFwqlFO/H1U985KX16iSsiQPyRn/Wqf91NQ8mjlOQR5Hh22OMVYjXo8sUO5
gqKXKHp3Csu5KMHcqfTbl/+ifk5cdcst1s9a3Vmf1AtUJs+fhaxk14CT5/bL+Jx1
bIHuqcOi54PMAcGptkYoI3P1RCHG+zRQdNxjaAFGOfjh8t91A3T9sMC3NolHAl36
31b1h2Xq2y7EkW9M9pvEUp9AhUkcvTJ5dHzcgFIBiMcpr5rFAFLPXDZTAwh3bmZC
f0HdcPI4PNj4k5VospmDYFWKZgptZIrH7JnfcKTDi6FwWkIkkJ0FJkcW4un45qic
Zcap/iRxArEXikeQssJ2IBvgWQRYqVNWyo68LcxymB6GLTGr3WTQJ3oRaEBsqBCZ
`protect END_PROTECTED
