`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EDWPcVoRw+xlQAxR38tJV9Io8QNQF4WsB/c3vd9Vnsva5PmRhvLcxH1V31SU3dVf
XWEOOCpzM02/MIm9W3L2ZprRnc72SCIOj6i3AovE/hpmDn+6npNUH+wVqmPsfMDh
PVpZx2QWJ56B4WWreUo9YbIGZFXtFfUhekNaZLVrclQS5q0UN6vZkaV9t558TnaE
9b0hmU4DYt3UmVHkoWomMDlqJw8EG3xpe8r8Iu3HeARv5rRzGPMIaqSZtMPsb4ez
1f9gU32wWKuUU5hzVjMCuPqDcN2/xhp9NEZsgeGCrSWKXWOpFPjJW4W21+PRIvze
qXuV5VfUkV0jN3RN1yD708X2hMpdL170/w0oydk2SfNBxahGBhGoajIUOYT3bHLU
XtfcqrpA4XeogdkNDXPhS8HMOvLotfTxdwS30beP/lUPGEDPiNNNDcZA12cGnNHI
sA2VhO5GG5ysFP40f+FzmsvWNJFiT3jfEJI36QNJP80bzvbkoSDwYvz1uioAxxbV
TQ7/dbcC+xXianQ9JH4t/5f3f+6MSQugwzWPDGbqcFgbELfeZBy2WAhgVMCnox/q
FfmE3lf+If0qulREz9QTK5UlJV5z9rVlYj9bJ9QGck7JZDAOndS7amT6N4EoftQQ
2fGbDmtCZNw83/ZpmGOpA/eg6Z13kC7ALDWaY0WOGZbkm97LRW/zK7gxtIIc9blU
7lrkxxSTi/d0Ua33C4zWc9Jocs0uhRHK5wicAbMf+1RwNxLViSHeA4DTnqLEN7k1
GikPlRjXiFdW9+fnWvtJ8xR7stC6rO7I8KI7Ya5v7z83bgGjncV3AhoiZww1DrYF
wfQFQYQEFY75nOQQb1GzJYYguqda6bPBMjFCnTwkv09o24D1k0XubYB5ixhIGl0y
wHLApYSs1UA9eJjGhFQfbcTdzwLbsYyjGwtkESvD+UoEN8FS0xtsecmwmOOgtvzR
oWYLwJMv9/ZF1xdWxRkIWuQGqX/uICDLOEQINe0Evxx4rZJfIlrlh1LspK3QqL1W
wEDuz9jB0xPZtVj/9kfPRLsuB2xRy+0jIkw3SThmey1Z/DcnTOqRP756EoKSBYNj
W91Dvy61jYT8cDaTN2d2/aOZjzw8SHhoAG9t+lAcR5OfqrnDMX/7WSOjAJKftVnY
Wl7nAlxYjsGR8THAUM2c+3vH5E8B40jjEFskrcxAMOPSQSWaiFW6lUXqUAof8P+M
Kb4Rd/MXMsjb/KuWaghzqkk/qlvk5Fwo/K/Pe+YsD1YlSLaDwyCUY73YXwm/QEXE
5G2iA3+PLDN4+8iSwdHB+zQ95b5k90pFpwdVk9c7Sgs=
`protect END_PROTECTED
