`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
byVFUcGeHPQrryXIzN7K3d1OxNdR+1U+/pkAf5BAH++/BPuDnfl3jXg2aAId5N1T
SLPodteo/pbFhZGoKAt7rzxGEXOIGY6ou2BdjlSHLD0v5tLg7ForkKCfBUWA+IcZ
pp3lw04/8BZiNJ/BlFxe/tV/D2d+mJ2R82EzcLBVZSW/Exi5TEemTFRIgsb+3pqR
ZVsPDRIZftz33KmrnFdw8Fa43PmkdoR/9KWxR7tSXYP0/05pwcnrQPTSTchSJbL+
+jU0tvO4uqzsPRl1C7klmhAjYfEnoHe6iRXBqDNHkKNaVB1IfBLFxydEjtHRCSA/
XBq+phHlipGl+nz+9TGKqCn3VPVI7J0Vif2h50XEEmI0xrFwzB1fREut+3T2ddZk
mVZGUZQT+IUo5Mu5balIKxegbFLdwo8wRkyp9bh8Cb6d/5odqGeVCKucjLX1hhl8
a3FuADNarfKdIbV3LdSvhCQOrFX+wz6IYZMWIrBukNPY7lawtDMRLrslbfR2w+bj
2za5F2gO5rn4Pf2R4mi9mCOAdz5CE/0KFLcptHWjjEBxe12PuhHfO7cuF9m+AVsi
ow/60pOwoKpUD3rVt2Q/Iu5U9KCXwqaZVIfIQCN0MhkSEgOia5HHBU7+axgodR0v
8SaI/WDkbFl2f09x2WVU28BdFeDOTErU+uxJymR06Ek10+DezDVQWIEhZx294tI7
`protect END_PROTECTED
