`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6hO57HJUIAdBYAGbpZiaDjXWgMH/z3oylBhKIsWLxcq7DA2TRbLfEGVEfFh+UuWM
Jkze2sQCRJynENX1EImfe3hKqC30j/N8d33CubzPV6ww4JDEL3wmYnPO+XSJGyjx
XOKiCey4np4Nr6kz8KPV3AI9HAYDtXXbiHmuFaLuP7N/FwJZbf3BAa9oIEqiI6hV
Pp++Jt9Ct0LLHmwzfXlbWaFKGQ1kBwMWgkEHf41PdN6KtNa1BGowpIJRoz1+bRtb
bVeTbNX8/MqXxWcV4AbfCgsjGZosgBuB6HrzJqUcrXxacJabnQxFWwdYFsM/4zna
6peHIEMyW+WMgrcJoBtII6yLCFK5/LQOAsOnODRBtTQax9AF96s74xiP+/eSBifH
xyOJ72gSiPQyp92innGx6maCUyNDjQJpleEzVUn9aYRUtbO4fVv6nuEg4lWVmTpy
dklaZutQ9XE9qhuAwFrSRu4BHm2BaeIxA04WM4PLBYHH1Su/GkY5o+TPOxtk/1M2
XaUDx/PkTN0raZlT2Pagw6NS1f94Z9U18oDTwDaOSktssqW17xwiNiXXBPXfJNbC
v3W7qRvMMZgPy47hpC9gJjIuZ1WVMo+tvlCutLIP7IU6xYqjWBU0fSYEutGA4WH3
HAwppIl2A0QiDjVl+LT4X++m0RJNAX9rvWWxV0at71OGYDgM4zKMo3Fyk0OQtKnr
sHWGqAT0DJjDqp1jhho+lwwtBq/trhHHp9gWw9s0PDbJkjHVxEgFlrZ+98C4V/Rw
lWa508BHt5LMwVoaGza5TdBs/OGw1PeSQ74gWbr7OUm0benm8dg1bqnbN8scpMIx
Vfn6KpJ962Ea/Ra9cEjZsn4f5jTNUmrcFzJVoVajb/C9q10UGFSn5FoSBWEEN+h2
uXLspEWWsckJJcJEqxBSLpHDuVWrn4IzYsi0RJH6mHsLcimmuMN+2H4Yf6jsE8ip
CzJsoQK2nkBXcoyDZIR1YkQnsohPvyi1vxnYWWJKWeeKs7gGkwv39mp9kenkK9wF
BlMwYkh4lxIWsO+eKTGAxcO/fTom3wJmBNsRcq0IFo/4izp2tHTb3baI7Cs4f3C2
k+P2ebmArosrVfLToVP9V2pK99d+LrIPWnGDOK/O1PDjM7R2vxDY6kA3IV7Sb6qt
gtMH623drLU7LVujULzyi09ckQShB2nYaaZCBZcYK7l0t04yK7okNb6QJBiw+XLq
`protect END_PROTECTED
