`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XN/MX6gTp84HTqf08IDXQFkCMG9DF8vPb7L7CJYugga3hywcvNHmAfbHXYoy1fpv
xI0ULavYaeQ6q/ClzLhd2egDFENrwe72XnG50gZaFkMSk6eOUalmpsXSait596jj
oROYcwtOp++9YajzaOc5RdjpQ+RJrOjKkHTbl5WNyOOXNgkFVHUl3wJhr9SVeabH
hcApiFlZyAzfrIvRMA9vY26T+KNesDq3eAOwrjmY2pldpRD5Cb6WPWNFzM9k+Hba
P5Ce947s1RPEgLry83W7GQ9LdYmpfmXDQL23B2h04K5QYv/9OI/2D0P1cQQvKh+z
ETGZyMjSQg49s8vmj70ZJHYo/y3y58Cw3vc5xCi1k/q+deTwHt1XW37kbVU7o+MM
CmcpCrB/lcMbB6ioOoXjVzhYmUQK+wob0hVNa9O0K0gqafHj1tu/Oi7RwNqeNTP4
T3y+KfBbjvQlVHcwHrSKiOkst1PbH6qjP7sY2z9jkg+cv1kwcqUoCD/nMLnDgnrq
jkUgA38LZXfOyPfSDV/QlRbYJcn9KJz1xsSiVVc3gmHyQnJJz4eoIen3FUYYz99s
0wBFJSxN6Z5sFy786Ax3wBT8QgNuOg5FxJ1f2zLJT+QcnA/iimOdboRHXfWFhw+H
sQ5lr2hxjxUKhI1wZFs+6mslDnuk0n7wbUJE72zzTKE=
`protect END_PROTECTED
