`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cbyWvNzhNBhN33HlyQm4YvrsYnHpd1VNjYSq86V58HYMbHJZ/f/yE9eMyOYp3y+a
fPukknONWwSOI3fIR/nsIpBPH/j3NoA+aktQl710IQfKlZBEv5TdCEDTUkhZe2uh
JKmh6w0mpoOWO2fDJwsbjCl28mUg4i9GsTCU8a9Oth8ON5vqyAS68syBNljYYPyC
ItauFC6CmgB73Sgzos9oYDnl0AVy8Ip+GfjOGp83YXBTvaTmjRSrI/zwbghwEW7O
G+7V46GBFBp/sbGahr/Lg9pDBB0KLrpC8d10VJTu5k4QgLqVMResjnYbEl02ox1Z
RpgXcOZqepypk+I5hRb+fJKKjYDY9Gpsi7CgGWbt2MPOkWKDXQiKg6O0Akv20mel
P1FnhTZ5g0/gZUe3WaQawvZELUnDBfg5u35dsQ3MuZQGdQUMODLyY/3P5/mnqNUx
Pxr3vwtHKuDsC5ucKA3MsqCt9JF/gOL8GCC2Zc6PuTV/zp8zyCvktaUdzcuJG5q9
BhZmgdxAleUVB83lRZWpp2Aqwv2WSR+mlDUFOPqNbwTUzBSWNn3pkQURVBh5prvv
81Db2zMwmFhilR5/Ep3EWEav4DV+jguuqNCn45XkbcRcjWap5TL283aqqKHq3K4o
17y3qn6/fynxn8VvK5xH2r45tj1icnwCAHJAl1xAeqCLB9/Sglmlkf/VP22vlUDO
fY44QH+NIX3ZCr970B2ryr3bADVtR5ZA5nqUBbpKF48eQApG1pjMk4knHsv76lyk
xqisVs8M2cIRAIn0XCFXRSORb8SvuKgq/bvZ0yh2jz4P26FZIfxQFQJxH2GqQTYw
A26AqZVdfZaM62PNFJ6+h2H1ocWxj4Ekt3uBrIlqKmK7ouQ1OMuENfV1IPd6GVH0
QsyzZ0RF2eLLQ00cu+rZTDqbgOEHyV0DHjQfTtHzHSwGWd/MRXDXUZU7RbyiH7B5
f9wyGSlty/kHR9eC1TyryraUvbxgaQkw5WCD1qLN6e5xSl74NrTn5hs9PyLEgR1P
foIGYkBiVSIp1FPAuc38Hj1WNzA2EdBF4vac03vv4A6RtL+DmMIOq+yjIbICqrNI
W4wmEMZTS+2ZP+qfCK7JQZIjZNfgfcgO2s7oPyF4Z6Eq0jyoEyTzl7+qkdHb+zco
7rt/ZlJLN7vO8+EkqiLb1Mqe7WgP/ri1cyBzBxyO0pfuxrsjeS5Y7E9yg0DJNUSo
9msN7ThNX4AUmu1euHftejLdtEIYljRFdrg+Y8RtUfWCwuEgbWd45Lz+YWWsPzv3
cy9pcygUznHRvb2ZdN2tdL9Y59us4EWsD6c8R1192us=
`protect END_PROTECTED
