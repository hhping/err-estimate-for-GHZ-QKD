`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m6Nc8ceBE9THCqPEJquGKLBIwA8w+TKw5hWAD+czB0CF8963Ewa00PvOquBYbC0R
JLRbpwOVJMJjesPHi4x0AstBW50GfN0lewKkttPET12eAQ5g7hH1x19U6ifjyZVm
Jiggt7qu3H8HqhzQ3Zq4XnkTWiscicihXoWXhuETW54gX6D597Xym+J5J5UI1itC
HXuUDXor/bB44j2lwIhmYN7wcvFOYOU0TLIheCFchx9kqz6kxcycLrS3kWVTBWkU
zk9DiYo0pXYFFGownYv6YirTdHBrQTlHgMHkySXin8fNrN39wgdqSYgjPyJfRmwX
N06y6tZj1Bnhm/4nvdgnVPkaxvv/GoBBkj/PBuj70h7yt72a+ctkUp+a5hmeU0RQ
+3gebQynrcGQaGOmExqekgt7fd/+vcaRLvbsrtUg1AVHCFpuZht3TJMopK4zJctD
/Rdy6GxHz5fVLQETx+dYkD5XtY7dIsfC93Pgk6S+0GmX+0seGgB7hHn7YFKd7scQ
AX5gOIVsAVrQ+6Pl0yVXwQTRkdBbcXztDTtsjxdBqrtdH5mDZcdd+CbTryBxzcsj
rVDegBaVBIqZGYHcfffV/dZOuUqMGf6DAP19FR5HjmYwbQt1DfAjCUQthTg5LhbC
/57wTU/mUNBtic3ZmebDveL6S2LS9Qdrh8Exa1CEQG6xTLHJVcVXpq7+PkZc25IR
C0tTJ0YY4ZIWdJHZTAEbww==
`protect END_PROTECTED
