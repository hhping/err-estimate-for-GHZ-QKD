`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pfj0r6GFAE1RbcGgC8X/8iRG1VTmp6KLes/HisIgBC2QgQX1HZkiAGaxtdGkW1+5
sl85z1o9jtlKLlEvb6rzNQ01VBaZ/VRQGOcvKmS86DQb59wTd/wduUo0vqcjVkCR
//B0SQOiQ8SOwnYfiz0hZTsT1PHsy0oO3UVduw4yw0D6fEGAG8SFyhNCuNy+ZJJT
nw88VortxtHS0wQGvIT/c+8zj2cMr/mv/0Lv8xlBF1UXmiS/Vq8v2uKNqWpMXfhV
ISh6wFlJJDDDy6oW0+orTIBts0BbLUryJbBHWo0AYrYad8OcDLQSYq2p4UpnumUN
spz+SANsDL2BxoibhJTkixNGYub4BtpBZDW3XZd/LzeEykOOvG3NW6OvZnF8CRYO
HyrvU4M/0Jpfth4ICopH88ZWuThmLo0hln/iSJcVDYNb0e2R5/7WjluFtM9fBHhX
KL5f7Fxytvn0o1Q8+wKjoxN+8mtEF3hY38RcnPxTTPgoB0dRCCWn/tMR8iiLq+Q2
Kx2EELZvY1pbeyn75FheBEgg3JSSchqvhQuW3tSdsQz6bthiPff40cdVRRriS1eE
0xJZtLANBdxN1BnAcyqymmytj5OtIFwjKfOQeqW6evfWGqQgNSHJKgITbwJ/vgXo
K6vzAHxptjoJivi5GdvMoydAWMFKughJmaDn6FXzAm/8AW9YIi8sBfh2yXDGmQ79
BD1NNXOpBXyM/KHw6M1dwh3acuoZdYmqHh9t476Gd2xQj8zdzjzyIlX749CZ3aHb
6Zd0L0oXFPaQ4uH/ih1SQo4F7FPOzxW7qnGjAJmqFabUq/q+2gady8/MlPVBI9CM
eQEa81dcMTp/COUidVxtrkmvqB55K2RQRljQlHje5cutTnS5NY+Uh/MJgsehz8/C
NBFpuKW/sf8hU+d5YJ/QarxBr4Dzuwz3pNVfhLKeGD5jtyJP31JziUpLp4uqXWGg
iDdCADD2BTQcCRAEV/45Q0NgC09SduQdcAf/AtJozKcsB7RYBYTpmUAL61U4zfMw
tlCzNitTNL+VLYA+VuwfUCNWmwTDnD8p7HOscWlsF69xUT3+tK/QfSWcLizoswN+
d8z1YjMtpNdq2++haPnf4pcu4rtZAq0TVOqxfvCn79UL08U40crk17fHmhm/9dIm
QNBtvjdChl+3PhNiGzvLilov69L9pzYKFMY3EvBgm7uqGsPbqtI8ELg7pUdIUCzR
TwcP4tiRUR3U5vYCLoli7Uohgpi9mgEwNRXKE4e/FVtO6PXQ+9+xJQ7R/oiswsJZ
CJJfRD3OBxGC/Ye3SOdqj1OCdoIBugwB6loZSM4LPtjufirF61mZ9fZ7yrV43IUx
`protect END_PROTECTED
