`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C6Dhs1FhLA7mnee6jth2SQU4St7n2SivWAf1ABogxUkSyVbL2q5vcmRcriAVrEzV
AsX8mlno5zwIYaGmWXWZUsCtVAeASzJLLh5JPqP49KNLp5FaPw5joio7q/90rxA4
53QCUfXNj1qXHKOzHSC/FV3rXpTrJvoL05g9kgGHVgxJ1uqSSIERWOHg+zljektB
phVDEkflLsOFiPrpX5czuzkNbqOSphL1vtx+6oGA/lq21QYO439tA4JF1VruuaJp
8Q0NKN1JN+CubvV11iC4rro/PQkqye/N6s+VA/VUhY+la0SDO21y/T6LcPWh5wqJ
ec5GQbFacYH5gSmlG44VZWp6TxY8l1r4anAr67yXQQBqWc7vkfBF3lp9c1M6Vr1Q
yBRvc58+EdqM+07YQG3gvrqTPlMv57EpY2NtHktsYr1cG6whEMnoQtsI71n1pLVQ
rix82Kt77QNSPKbP3B+yxOn+pZ7nwpcygTYdB7deFifZX6seQYbLebALsIo20IAq
eVB96PKUtweNP992319YdQM+HaHxfSTKJp3KZS86PwDH1rQKkJnTbMkt4fBGLB5g
efFc0gMcViSxu7TYfAwYDefLmkDdSgO4rcChnlZkZyn14Db2PvWuS768Wnqok0LG
9dh4Ic0GuxNEcU+l+Z5axXup3wcw8hWlopuMlsAMhu8CY6p+H5dC5+/Xt8uZXi09
EP7CRoWQCfs8ftFxeUZ7LgbsRnqRxyBLsVMURDQJ3iw6IqQ6BTFbmaoIF/1DYFA7
wMKFes8WDWahkqNLDBWi2dCv69SfXVPZxv98LabgEfLF4qX5pyHJS0dp74qioL1j
a/ihRoHo1Ljz0vc2JcnigvwV5gYGTasereR3QPgeonpYmdywzWfslHcqq0ZIW1Vs
hpjXgKr/f0epGxGOL6y+QTsgI4A1ef0tZFEQsDzf8Tm0p7O+WsKdfZAuLhQbvUQ9
D/d8uAIP2mHYyBi86L8jQGUhkPZQjq/k0sStiWBPXKde6X4Yc8lx3vZ4oZE6HAdM
rZ8pzSLV+32NUrtdPvO9stmiYJ8VpR4/txAWE0E2xPKpvn89Hf/Ql1WBPEcSBA6S
eBYnvT2bQ53VO6K7eLQcy2tnlIDY2/frQwAw9hKx9+LTxG7ElPzbz9ytiaarc8Nt
sBddwnHinv7LtUVBmABhObauvofdBbY0OrR9x9SC8BRt4eCTxELEhyuGsLN4BrHZ
eP7M6ovXZE+VUVAT8H+SZcUNJjZuVgMLlEPQVFNY30rvmrHAtAIhadZKLQrd7pXP
4QWGoQhFFyskYF3Nda4tYgCzZtEh+RTFO3HPt6MMTNO+U1nksAfLFTdarLUl58P9
U+ejfvipe3XtpdShFj62ZA==
`protect END_PROTECTED
