`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PwrM+l3K5OBpAYvbp+jf64iL3GGDOGFHKcZyMez1g8/b1yKDcuPaEGrI3QrUIRQr
g5rrmgUBUxxBzRb9LKppdhzrbDK2TqLHZUyRnqphH/rFgIZYxiSxlh+bgeK4cuIX
KkGDUzs89I/M5K2bCiug//lWk6+ityeKCrGeP+HYvpIsVw8w1PyNXSD1zSW+Vk23
Y3y+2GXnHrcmiHyDI240zXT3CnI8dy9A+Bnzj6TVMb1LLjOrjjB/XCSg9ScZT+R+
DCLOka8+liHThkcz2TUX5Fxn3EWmdY9DzVRW+o6ZUqCbgU1wdYmYDamCcjXZaBf6
jVOiVF+0cfhrHsiSN/lyG5j11jm6b3E6lS2kjC4fNQxTrzXmViNJ/qNxpX02ZTji
1QSY90SZIOqozqPsy7X7CVf6p8LpfUb9Qp9zLWPKFhOZB1DCcwY0HMdVx+hFk5Qn
yZCvmvztyTdY1Q6ZEbtNQL7USDOx8upFI3wO6293qnPZk0AWPQxuFngMN29smOSK
P4y2mg1SE2eSMm4TJgPAF4TYSPK839YYlZLLUa/vTmM=
`protect END_PROTECTED
