`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JCbAQ2zEaE7LosPHlqHruJiGKyGqqR4BcT2hx0aGjsAqPD7TFtTHfuQFVWjv1Crk
w5gJFjGfELxP2kqifyfG1KexwLFZk1oYp5tteB66NoyfcYuZapkY2Xg9tN3Jd7fr
1LbXN1f4pzL2R/KHqdC8K1+xGOixgq/hbt1chOqB9tiHzCMRuiPmw9JMX7gCXGcl
nRUVxezlY1iKjEKW7ZET5Ftr4qSlEOm/hjFGo7VmUIUBCnNN8w5fbdPlbewIZfEY
eTIDrzLDv0UjOqlzz0OEvTEHCgoZ+f6ZS8CivzYCxrxgr381waAlACWOiatPAB2/
GxLH4hxli8zQpn8o2QafacjLoBbED/Yan8WstEk39tonHU2DkSnSV63pKnTORm9V
A/+9JTOv1EvyRAdGa9bqpPf2aRVqX6CDUWHcb4z36Tnpj8EzxOLaeQT9NfReLlnJ
TWYcUDXo+PohBoWKHuTo/Frm8pKh3xTf3joowZkuZhm800HmdTeLt44vX1NcK3th
k4ZTTEuf2OOE+Fwl37mixQQF8nlc/V11vB51OAYSmLRqcdFeIbjc1DbLfQeuf1lX
GoJfxY9aMV7cx5Pwk2R1rGabRT1e/urjOtY5k7smN8GoR96RyJQPPxMRcO6XSXDw
UxuhvMXzs1nZ1SLqSeNjtfKO0ObmRbD1cOQyH1Mf6MbSMfeQbExNeRBdNlVXrgyP
Xew9jyPpl2nk/LuD97HMkdCjPzfFviPqRDudOsxfUlBBBdYHDX4WI6x/heuqwKHc
4A+JKhImiq2hV1quJrE3DGOjqjYfouIzRxEI1Dhcjk6jzy/4/BBA80QCIl7GYiBD
`protect END_PROTECTED
