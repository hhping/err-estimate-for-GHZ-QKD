`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7nNpuIQs3sD0+hnuanrG+90aaAk55ThHinAm3m1HmXLDGnDnAl4mPbYYZIMAYU+J
Mi11Ga9RTfHzsv/VlgmSLShBtSpFdD0aO3okPeUIBcgLcOSEVy3UoxnIqnQYZFmQ
RUrZlOEYpzqcgtXuYSMkV6e77BBKIoZCa32eV1XIOP4RaT7cmpV+ghqKGzB6ToeB
ty0w8Xiaic5yrMq/KXhZ0vFSDn5LsYRiyEWHvkN7H3FZMAPw7HJdsVH1iU3udB2E
kAFdd74ZbOkD97kKW3pZ4U78lL9utEVt5INVOE3w8ggHpuYCGe8J68trRaFANruc
4yTVrBObySBW4gzdifJEPmWjkIw9w5gWPpzPZKggTkycXBWSY22+Rh6tYc8pzpcu
AoxfKjbVdchGmBaa8QqW1ORivtQ+/UHNlMHX1l/iV9AME6cHE/8wQvBj+0D1WFg7
iGVIsxx1dKuwzatEtqpZXu1BuAlvkCV9HMmJ6AgA164kfcT9tAH1HVjgMkPIVfqZ
Jzx6a/IiXIsiR2h/0fWrDtdI6F2pwccPbuIBTHTFKl4lrEUF2kHG4ENXiXnMRT5I
igL3f3EvwC59rCaqXeuBbFMT8pgUqGgZwxHTYpmE//zg94SHkswUOWHaOGiZNZ1L
hEtH4ZitKlatZSYdddp7ZhoPQImMYwg3R2wtjB8UxmDyGXMiLRwAHU8CU5xBzEvp
vuXEHdgdCll5haK7oo913no3d2KJ6SHXdyPYcLTXoLclWc55T1qCMVGh4UHEKnw5
Dk6XCCK8y3QmWgbvw60HXGX6IqE5vXlgIFfB3buBmybrFhQl0lA9q35dSdURhNzG
a6iPYq/P2OuToyJrViA7t9T2JribDHrGE0SpA/WjyEKMSFpx2Lndi/Y1eSp/lp+4
nysqFI5uctEdIBaaFoQ6PQLy9YdKKn++NeqwtmkO5Wl+faQ7643poLG5BZ0Qm+Jc
5vQlqLanmFCkY5DrEHj45Hz3klqwEyUO5vnIzWoXJRCmdYRPcHKFXzitDgUrQyIh
XMUY35M2JVq8ezE24fPdXdImJ2YhPosTb9WeCLVVnW4bxLvDjnsnHbrM1jEtkXzA
sRwwNnqcW7LqD9wp03RVd+QJsFCfZ2M/3qJkno73yWM=
`protect END_PROTECTED
