`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TUbpAFPpxORGBeDCmhGN8nkEIqfnIR7Lr2tHgkDwXWu7TQzGXNlMMqnWLojhjH/j
Bp0cdXyTshESBK/cF8J9b4mGI7GVCFjGzmjrvkHGSdUCTjhyb65L3rs6y2irGd9b
HVkAhULdWpKpi5SW6LxDNHiIWNbRBad2MqEGj+fdGB9d73nLKuMZQHa5w/sDqITl
S7rjilIrDkYPNSj6fiPrq9R7sFIqWggu5PciLVHQB2Gbb7xen2KLGuwCXaYUVzZa
G4w3elyKgETncxLa+C7zXG/MTSSmiGPM1j6qHgJqP9NZresgYTvPA6Q6Ac2vGhaD
hlUhp40zZ/RuqcSsJdC0wB8/Y6TfgY4E/VKcCdjqoeUwt9Yq7kWiwiLRKCRVzmDr
0oDc2wRkS/rTnYMaW5FFKnxmzkTP8aOP2ejTEX4l23hy/wRgH1oEXPcSctw6VMfC
xvZ27BlRQ1NkV97bji0QGQBq6VXKwQleKxYdu3cxh1EnJrFvgPOUf+XrL0OCoZnp
fxKuWTTRRvbtDL8/6fI/F/lOToeD9ei6A9wv+luXIzhPBLeQ9r/xOYc/hScQsDv9
QccpQ5/XXdb2xIoMe1fj7P7xhLpip6kwLw+mZXDNqvRUS/M8di0JOlphkyGdFs2y
DhOE69sljE3ffHoyL0TBbtZzSdQ5xoVo0Xw1bdo71kRyVeoolLMv/FpqtrsxFeg2
78oR19m7/0ZNdkX2JUB+1XGXvvI/pxdjxvRNmkfzoGWvQS5GNn6MVsXIoYTLsW+X
XgPcxtmLQ4KSZNqQ1BZRevwgt+pYwmxCalZ0NYpF87ZpYQ7b1wbEmcB+3gi9B2b2
IXh7W0fmsk1D0JVqr/Qi4v6xhF/Vx1mP6K8PfUNGBNkp0TSxLSAXGnSTkZV4x+c4
ADW6fkahLAishE82nL/2yhDQNbTZ31s0RYlKgBrgqqjNway4QltGYEA3UvLfmvh4
N01drVffIjVpuzMg/90DqBpl/VFp1nJQGo7+dvw1v4PROWvb68zfouiOsfL4jg9x
d3MEhDZNVjHcLa2A+uafKhRRulQkP6eRxL/lJgBSBNurAmsfpeec2VXud6W49ix8
sxLwSuTKW8ZpcaosV84FbXTyNLpjW37OkfOwzibXSxhkoWGb7p5Nk4izdBVCmFkV
qCNSqKdT6LMl5U4ZyZjSJNR7U3Sk56aCT5yXiqfKJCxpcPgbh2WhUIhxdTRjohL+
vdNy8RKVGNBQhzsbSgxoyWEvHY9Arq0g6TRHYd9z7tfpWcN9Iccl7vZy9vBnkcha
m7axYVYZFk0yNkmmPRU3Dwof2cQbiph/mlNqIKqArNgAW7M7DLMP5G6/lXq3QEl0
cszMB3dQnjyyQFISAVD4uPBGpENXoRXSFYIVfiC3Ko/Cm98h9sabpzt2YXkwcpQ2
dxC0IeOo9KKz8NKY8Wz2W1u+yzChIWTgu0dphHykfmKYz4tsHKMnId1i4jtaSIoJ
iYZByCO8vCt9AWec5H9h4g==
`protect END_PROTECTED
