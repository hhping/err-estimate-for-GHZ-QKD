`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lxIgLS13eIPaWA554uoi3vYHduhf6WPOtQ/paNG8a5QrqmbETEh60x509und2odW
JkYYBLkuNp1sI8fAscp7TTky62VctxyPmPOz8SZ6fGXI4XFA9IrnjBpNeX47x9ul
sAdCb1vbmwRZ6qeKGdhTGWKdJZbJO0cuJX37qSC/kG8nG02sQoAlqEq1A2Pez/ZI
VrZ74noHQpCHjNl12qlyx28A9dvnNdSRIuWzEE2fFYubDGpZzAgPGTAa8fWlhaW/
05TlUO0K9662HVi58TmFc9Fok2PO795t4e4Wcd1wrK3oYgOcjr0KkRo1tM/1Wmr/
xFJXHA587mftv2EyGLGoBGQc6sVm9+mdhhULvdU4naYxb39nGHsuoNyttPGmUhNi
o1toz3AA5xXoN2MhP1/6nyiM8Ap2GpssRPohgqWmlQNahj0M5MC2GDNELRP1EyJR
J2R7k5nzdOqBOt6GCdizQlQ2eM4aRxAM9Q8RzjL1IsU4V+Jnckj+cRmU7pMvXeaO
L3BA/oA6ARJHakpcrkGKXrgTPM0tO9cUf3MbltPBRbHc7LKBz+ikB1lRQ0p88Ob7
ypasjrJmHybgagXwAf8A7o1TyzfBIrNiSGi54sY/I3DcBtpaMqw6KwEylWwOZflX
GjpbtNoowpIl+A6lgPQq/H6zy6KQe7ORTTIme+TzbJuPlam/XTItnU6Fb2GBK+y3
WS07rg5WIeZsj1xg79GulZWfWVM3d2WNzTQ/hj85fRrXwlUFHtr2otPuczCqNs3U
zKlF3eenFKpb4r0bygkw4Fk7tTlcCkma1yaBhzNC5ykmGcGESTlmHh9fnBpAeYVC
ESFHuHd3qQIkb6ez3XXWGCarzxaFi2nJ3Z0INtA0Tj0LpwAs5tnRzTrm/Jnrtvef
b8TSGKXO5U7chrWSjCpEx8+UfWypuhxnwKvVLNcj5+Ukd7UAnnd7E0+5VIcXS6uw
knwttON2kbIqWXANa+FlOzDAS0BSmDLt/QCA0FgZLT9RkeQkg9Xc+6/nExUfB76h
CIUSp9ScUFgvQUMFKiFqVHHGCnVMVtk0CK4WyJ7KCbEQTE1l2d2pFxNNtqp77COx
f9fiWmT7ZBzNcFDWh4nnZAVgcTTKc+FiaPNs8wYC1s5xzVCjTarepezPXM0YAJf8
PI8QjWeQBbCTcN/Re6nnEyUmE+gyr3uwcymSQqaXyXWomoKDlA3KiMVwrEY0wtnB
RDhH9qFIGoB0NHEXU/7FTeg93/IllnAHBMhWq7PqDaNAOXSLsFvlLMSNIBBQRhQ2
sBj+vsQS9KTfJOy4QxsT00Vp7d70bCvvxG3h2o3sjdIKSIWDl7kTveASeQ/FQnfS
QlgQccSjypGdY7ROgw7wTrib5rmYcMTKC6XXe/1XChp2xUV7D0mNoep61faCkg54
0yWbYXV/yIlf20a1VrcCBhi/qigDmDO/lesQmo0uxbF7Vx6RyjxNdK3fZyxLOaq2
04aOtv5C0aDZIVL74X3/4sIHLF4Tb0hyvJNrKPuYsHwWOx2UlHbF32xamm1ICCRY
ZLlHS03IAfNy4acs5xL6scGAcaQwwDD4/4sSCi+NZvIaMgqN2nghfgRTZMvPI8tF
dVrnE9ASjSAQ0MxSfRkVX/qn7jOZ25m9oKi4FTgUN8wBmmBJFdlNsW+TS19drXkw
pid1lIR0jqK2uqczcz9y0d22NUtCAq/Nc8X0GfwPP2H2S/LMnQ03CVwn9GE0yvYk
dEdoT9JvNH5cAsC28nObCGC5oSqMPBJOTeblx3GQJTXU7sXMRkVdyoY2sSzongmq
OaJSyXvOa6vNo+6VNqw2HrDq83LOTmnE9sXQ6WmYEI4My3ycB/+X5NMNIm1HgR8r
3P4iOVf2HoLdEsLuaJnFuXC8THdDTsJGYlhOHF+OB1d9jF0CPJv4j5ApDYXKIlhn
sQ/LjyQ0KDuqOT8qb/Xb3aor7KHiYz1fhwzJyyMks07bNH9WfUH9kpjZ7Z4FVXM3
Nwkgru42sUlIXbN8cHMtRRojuBjNRnwKfkmDQg625NMYDXgsKIP8jXMSXgNGWBiT
1WDHcBZWE2juvOEe7YNfttt8UD7WLbTW3W2fulGhNd0IU17lVvuTWJtbDUItINi6
4xdCnxF2wgm7q1GMel+Ac6hC6/D0UZVjkxaFpTx3Ark3GkNkSHqdVsExpx+p7+eO
0IZ9gUQ/DlimQmQIkVdxSuURtzdLFzxNvyud7T11TvRFkyyOeSU0bDgGkWC0JJc6
wrsvVmm2S4ULyjuNBo8tT2XW8hUTZiaMW+P1Hf29OgR70nQybZJUFBQ5ULCNzAPH
YSIlXGrI/uZ5zl0F6yEyCp6v9nUXXMRedLVOCE9/xdztKzLE8xCkSI6uVa2amNqR
DRfxP/gxBfICCckzaN6B0Hovvn9TgUYy1SSCH5z5Cuhj/4T4kP1KLFOUoBUJc0k0
ozDF7+UbPOILGW+CRMNlKvSuCMm2NWQxru4PwYMP7wRIyYx3nmd20YmTkvZDNfwp
+0foLJRn//yirON9xfR8XRSVSp/mw7kPdDdUXcOW2Lztn77uf5SmMvbcgGAj92dW
bcff87/Bix/qOq+aSD/JKfLukxpwXt8KKgCsN4HwHKU4X0Qr2taEgjV/9K9xOogb
moL2nwAba/3QpfkcKFE6MuVbGEAmfsQkT6rdSbSS1JS8TtHCu38hiJsODq5g11nM
CFyDlaVVC1mVTZs/cvpOAUGaH3z1L7cah9gcQYSZ+RHrvKsdoTFqsH3vbFA2TZQ/
vJX/RzJXkcmFx8gaUW2fvuc/GTRM65KqeloHB7iZY3hQ8pWvbTOqooWDURaEeLau
zhQvFErVNhWOcsIvii56mvufZujzV+Y0nDE9RJUHY2qWNB8OAAFJoQH8tHKIyQpR
J1ISBVM3uHT4ZdODKKJlmT3bMQbgiNZFT3tODKzW51jndu7eL+oWqmLyo9qD73tT
Yl9wbzt0M22I/jh2s+b5nc//i3pQnhhYJR08navykvMLZZP7y1sAOvw6nck3CWfb
MF4/HixVN+LTffG/0H8azirEzGRw41bxp3CG7jceK0zDpbBkdOgNkIVhtPwJxgP6
ylMbm79Cgkus73lsE8vadhp5Yi5jYlOReKiUCVnF+nhp5w0xgkC9P7USsX0PfpjH
FxZ5Mk8Ix+uJnKRbycazTWS4ZFK1aidGtSfwugvAMLl8EfxF5TBxop6XDrToCn4F
UzDCKY8yPJDgacJTWjNUqiD6Si3PIZSMQUriivtpCEPbGIBm8TVk+9+Z1ZOOhg7R
SvM6/OiM4Y1vuErX1/uODqmcpi/SAtpSiXGwno6WQDDGVUK4/QXhSa+Qs5dfN59k
WwW3MRGnuoiPqD4s72Rhch5h0nqfYH+gsqFZMGVP3qVbRAHZbGDSC/xwuchloq47
mcbZg/jQ7oD4jFIk3DhGgfNWFaVQxdjx1Su1pP8+W8jDx3xNFEudPiy8kCf1yjiL
mny2GOW0n2MVWHw1BOZ4a0dk/j2oa9GHeg4tU8ESxiMeH+gw8Sv5f6WoMZXYcWaF
gaAzREtVVuKleOP1Uw6jmhLBQmoHAvl7H+weRNzT+kwgioKTgBr5mwuhHED5JrmB
HnTi5zFW9a07e1cywvQ6KdqAUFGlBVPs31J2b38CR2cuv+p24wJAamihLU9taXNJ
Ho98GDZEIzDnMRaLY0TwB7UqsImP/R2LdKesFJQjb0PMgonebY4moVTlD5c3y2gb
UGNjGlpHRJZgvWKxg5N/vQ3s4HVKpGj//baMF0c99/zt67N6VwVlkJu0X6fOh3cT
W7MALy9q32smiEbH37G6WG+pb4Yajid8v5svqUB9uu4L6UE3vSt3LaC/IdDsW1au
R901F7XE8gsStCHZJbaVLBQwO/nC6SaMlNDV6w1bgKGd1wZUYWQ5tYS4m0AYOfKO
eAIt2FSH8G2qWN5fXyf0CBku72VbX6d2GPqJkPZv5N+1TVc0Ceb5JCRXiNI5oWm5
zwtW1P5SkZ0yFzCtX3wwJp0Uj54lxiHwkq67Lf51Ci8gvmMvVnfxMaFAYPKqc+fK
jUUz+J0Ga1DO7hZhRRSWmY/A8mbwR2WQj8nj/8CY53aZsUHHILPUILKQud2k/YcI
Avk2iAp0GrCXWGwgcpzYek/d3abgC6Cdc4LiHDvgkdn/mklb7PxNbo50rZd6BJGw
DFYxUx900KQAgEep1cwAf857LQlCtNkcm/Neml1o2KfV4EIsJlRrYw/us5gYkKu+
VoXEpqIpFnDeMFfooRFo83FEkqFDWcj7NUqW+FLbra8c16F40YvWVbTcQqJSDmvB
WESmRPWBidquWaxpMmvnXAkas60O331YeW/LZYSLZepGOl87dUioRSsno44yt6Wo
hVZXnjBBrfCK/OBUXfNX6p8dBHs4r/eJsaJbKM3qRQImP5H1rbJmFDX6HbIQ2GYX
f3fmKN9bUmpmr6Z64O6aMBzlbECerqmj7NAMiFi0wxt5k0mubaILZOyUtr+b1q+u
3qMW3vosyC2kK0J0WcUudZOT+PFisqOAuHQau6wiwbf8wFITxOeNMQPyjW10j+vn
kX3LIQWNegwLMBb3I/1OG+qingo6/M8fWw2SyfFxqki32a0rbAIffEmJnWzySlE8
AjUni1ymHnV75QrMPtwnJAdOuAe5ljQF9oIzYlLXnIxwMndOiy+AQWXzwZctfBxx
FJ0qrO2nwL92c+I9oAJSh6BEQ1u2B80wG9FaroYBP1p/Xs5f4+Esbt5qynVW4uiW
vTZDgguO7LkapfPIs6xE0E4VYeQ0rdDhw+qGUJKrhGmo/MUdIeNmnVpUjyz4O6dm
laMJ31JAQKC7Q8hI6Z40XO3aDVJ7lyNg46GV6eV41roGWWBvFQW6DcWgelyxntrc
PqnVwwcGcUlMcihu8U7jZ2WkVNWEaVqbWruEKQexWHibcCwn+L3IetimzlC9bm21
3zxH1pB3N85nnoFWSciWEbRPpxlQxP1eGp1ca2fiCbB3xD9B1Us5qcGD9vG003SX
K5RIgQzZlkilU7oBPk33RBVKgo57u3xwPm15/pTDl6m1PuLCd5thpwFtwhyp+uhU
w3TRav6EbZeYMnsgEPK5nRD6csKafIloNDz2MEsqpzietbOHPdNwxn6FCJd9E3aj
XH/b0dgCQHoKk1VoDiDiALDnvMe2UfcOmhoUS/YAgTzpdC5kjy7J/elLEOzWW7J+
U+MMUT9VuWZYhrhm0MFE4WZTHDZ3ayw3zd+M63Gtm8han4hQuHpZMq+lqWvqrNB+
FdhaafIrUkGNWSv8Yv4oDPO+qyzPF3Zl/ia/vp51rYaAvUu6VGsOfboKtJ8iIA3i
/PIEoLx5/okcLLlyZdOeYExJT+EVsugdhdlFFr1E2aJyzjmkmhGrpOuUi76EqYwR
m+OeorYMGlNzTw49RXhraS11Mx6ajnNbb3qy4KmEx5heED4ez8uuSTN0GDTHQwNY
RCjzzbPqoSnrQew3MqjolQg1a9BeERGZZNZdeUs3/mfgsCVFeU3qeR/tN91BwTgb
Cvm6EPSIDYjosbXP5DgEBr17qQ1+ffmgBVfjIoaTOqMoVQlV44+gbVxLHutUggFq
kIZQS2mi2m/7a46pr03TOibSCDoapBompKwFdOwkUZ8IJyg9RADRgKe63Mm7ZCQ/
sz+EXsccWG9d4I+u3WReO9ABE/xanCEJ7Ub3p2Y6A5Y4+5l2uTlP9dMWfJWDSWjX
zqP2tEmXl8yqsCJsRSV/eya/GH1I3Sy7rS6kI/4u9nsTkiPh5n6vsAij7yaoXXN4
r4C5IngCvi3LKXFuI1LzkCKCmCYnKTZHHEYOO7HsFpexDhiVlZ3wnSuVpujTwWvR
nfq1//5zaJM4DfCJMZlhRfN5M4o+yM6BOX+JWLulFK28VXFT8PlWsr200lMRI+VG
QvxKMdlDnuX5QIdhB2qtkbpptfctSZG2l3PwZ/QqtnkPA58GScJq/YVQhcqTgZi+
OOiIroxulSeiwMwRNvBTxuak/ZfEpfjkC7ubig2m3U6SPwxA/BCRLsa5lmQhRgH+
qLg8vE6vFSG0XZcJ9D9kdUq91CTs3WHRUjEEz8uNALmLhZ19m/gn1k/vwsLSsne6
FvxSN+SsnurQx23ih7kyUGM3afp+7vX5EfgaAH9SoNHTKsAB7JotUGxiIqvaaLYK
CpLy2de26PsPLPeVGhjuB/yTxEprI2l+apQRVP8u+fD9qDcpTrLa2LOzQB/kwN9q
IFOTIT/4buiP7EgrtFy/ZH5ibLTWuw2J+BZdAnpXCRGpP0KAarP8t/pl4WJ85qb4
BnlZuRy7eejfgtW2WNP+G0UsuRrBvEadVUAVAc1mwL3SwaWeUvQ5WD5HzeENcAyU
CBzZRTwbbd3cpEK8h1yk8w6xOyThB4/LIfGqyGlRv/MhIxcmQHSUVwOtkQz5NKEJ
zn9bRXNt4aKcm9RAtFk0prg3vPxiNQf2omyCE4IzsMIZPjRvK+JktkZjxm3rUPSf
RoikEMF2Z94nBtRkft5zzhH12qC5iJRROgNDqjDvxYvljNE2hblbouEu6nDcHu9S
pQZZAw5kHuFD7DlCKyH67lEJ51r2P/A3+C2IZf/bUGcpn77gWEKhKhP67tiIOvtA
4RC8xLaPUyNGu4BhA4YGr6EP9YBfmJt5gs+7qxZFo8B1IKS+n+RzSXKLGkL8N524
PnHeL9pDdXunMma0jzGP9BRYT79lCLBEzuuz6p9fzt8tC/9DN5863czf28uy34eE
YIRd19noAL8w9L4V9cgWNMWIMEBv2nC1a1HtDkSdf4v52SrJtg+TYK5r49J/vbHr
YlkopVHmIhGPtbatezsjLx7AfIzvaTDWiBR1CgksyeZn17NRanOefmi7jLmsJCxQ
lHEpb2jzyTSAj2xKp3/6ZBVNS4xI7J7V2Vh7/EWWgTgxejVf6GCGi4l5+WYXVe85
SibLo4NMSBZO6KUneI0IFQC+4Q5KZ1H6YTe2BQLpHw3CgqwnH1ZppxzlIqvKxzXk
Sf0nb++5EqD+zna29TsJWKTREE+EgULDaVHwxA0YBgeOkM2KhsVU9WKt/Pt9e2Ps
v4q4m/1Bit6y+3QRZncZa6jqvU9s3EFF0WFY/dnEMtfOidOYN/6CGNNVW1sX7+9C
RAtcag/fL977hRfqNWbcus9qq2Dm/JfI0nhuCeZlRhUacV+YRmscFEJfOzrlk2c2
O9BR6uGd+91rvkSDEc/QhjdGfWepDJz3jSTJ6atwZPrgq3xDTdfI4TJ+zVgs4aDy
7Fc/y7EhSwT4ZqA+xI9pigYY5DJR4HbWTgDPFpaz0U8SUI1qWv/vSACMAbg48cx9
SQpuVJiBWx3dB4jxvOWMM6raGadRMDxKO3EI8FZMBU7atcttQ1s04Ft9rtZxF7rN
01dOjjiJibT9VpyJFLBJ5MpSgpP/tL3vsiMwO27Tz/urrLvrmpN54PcVprg5OSS8
DAlEJQOpne2ZM00BDzWTTi1a0Y/1T2qO1PBsZe77MWL/PCnWmup82yNGAmTbe7Zw
5CVWD0U38F//wfqyqfWkOXeuOmlsa6qItt8+0YqHWLVrTeuSsa3zFJO3iDxYqvrK
bGBJpBZ+qUmLlVzqHGce2EtwRbQEJ02AJLawDONJo+vQiSfmEP4DAGLXG9l30QWn
9YWTKO6zF0m42f7E4+SlyZ5/lj/PXxakTjU93bhwUVE/PTFV7oNZT/csL2xVu/aV
P1e+YXAWq09ZgMoBCDMGqXkdMGu8T8Yb8u1hI6yu/dEUqhiuY8df/VmToa5IiApj
xWSeWYQ+daBbAuTk0PdPdbuyLjt9X2rehQf/x3tzJaYtk9CA7QDQYl7Iiuinb5AH
+PtmGS08Qqo/LWmfO7tepr3gbj91KGqcdunklbcKf1/IItgKlkeAPgT9WVMDzLQW
QJmEv2kM5KLIa/4QM3jymaWe61OQtxaSBs2BVtT1ogCOMwu4tGQTN76sejWgSUcO
7i9e35Y9IkMYsVHRjRhlHbkCt6cid/l8FQTyQ9rpgnD4DtKRuAmJ+1O5yJd7BbDA
h8WZjhKJSNN+Kr0vJGQ2yT43JsZ3wh6FRGM3puppz7CiYs42S4Xh0Y9LIHHhmyum
rtt0ubx19UkIxjLAAaCCa56cWukzWLyKAI2aLvyKLpetwa8WNOdu5yJwj6E3ULtS
pL5M3+r5V5lhl8LfRoAbOLApMr/T+ffnseab4RC7AtnnypvznQcdiY3WvQlUCzav
phJukLD/vZCZJIOAmUkeEG9QsbQkINDvlJ+azci20hvM4nEZm5ejHf+TmMmdSHiq
SBeWfNmFN/sYS76AOTTrdib7QfYQt0mdzaWHlQAL+RuvoImFJ+jsGhDZ2K5v3SHo
Ac0gND6fv8vlbXXe1sGi9eKXZwhv5KhUUHsj5+vM/Hfxpo4x03xvaKERhKlmMfcM
shhrAy7KftXq8jOP1PRXqdCDA97JFp6zLvAKl2KH1u5z40+ntILsSDdwjVetIuST
+VzdbCKm1QLVyl8HYcjNbc7ZiIqCYbLb2xxmzwTLNwN95QzCltwYiti7x9By+W3p
e/XTTaW44AZuycrBguRQvkpHoFVvxHEQ5nyIqLSXYP0M0vS1/HZYF/APzdyQP2mv
+ngE+uhkLpQj7vxCRMI0f6e49t0gKB+aWAlCcvk2GurgyMY9CO3GUuZEIFcCE5xN
nmt9GpUQuTrJV3pikAFLm6eKT04UnOH8v5gmE1LV+f5Z2VT0Lupq/xVESLeUbvCd
3wSTMSXMZxFWOLvc9md8zoLSd/8zcXo1r3qS4fHuEcAFjJGCJzuwnlqi6PJZ3P4J
HPMV68Fs9rzjfexcBQ2GPT1AgemDA1EuLPuhR7txJjwA1kodeT2tHTwrq4Ymsrzw
8+6+6osb8Vuf7TpGSkeEFGR9H/G28UUeLhnCuMIncFh6HI3B1kZiZsrUqfQZQdGv
yG8wC7PdWxcMchal4TwFDZC317O0ogWp2PxnLdfq0/zO6bkdfxo8fPywPgFpT2rQ
I0fqC4PiJgOeQ77QjpgC6DVIgQmdvSivE/trobC35gBSKs0E71GA4l59oze3G4f4
Y/RwpPfjSkeZMME6YC5OKBwRcn5/7mX6ENb+uoHCBrzyp6WmX+/euiqfeTyz4M9h
yjfzpuPSMMvTgFgtic97C8GlxrqPya4XuGudbe3jtwsn3WTa5HHyhslNBVlVG2Ef
swQBQ2pT/j7xOYTAzB3Qtnq0Ojd2FqoNQBW1W8zOy6WOR4VGFQseHyyML2dWY9lW
EFgqfBok1KmNHDTSJcycmD068MwY/g9NvxwtWVVtUy/gr5Tqd0XMpta15qJB8TFM
+FYrvaN5/v5kHAjXXXdhcVghl3yMUvDZj7+eFWV6mKnXGH4qJCQvLvQJCYhjM2Ow
OMw5xx+/srPQ4PBNP4VA7ZVxAyX4GJVnvCXFhTvyi8n6rJGxJyi1H7ktk9Wpv8QW
qpXRLLn5byH0w0shqh3gQ1pR3we3bdldOmsk9qdZsaKyeIyG8pq1IzR1Indfpiib
HS+4/Dllvhm9IQUtWt1YpCVZ51RjenYQMjdphL+N+EvOGv0shtyWr0ghGbdzoF4W
xkHwN4F/Q5LRckFXSAd68cL7MBIFGRMoh9E4rAeQGzxr2MxV0avH6AjbrMD97TL3
DTFvEPawVX0wGznH0TD/icusYFB1MbP66rs+5gZpsvdJtSIi3HY/bYAv5YOWkowr
8wc65vJ5SmwSEGsweqlZhezeM0OnLwmayLfLZIUFyRiIF2/d5DdOxphmg8xr+KN0
Tq0AYbAmiDtMgbvD2DlbwRH2gp7rV/VtH/KSUlxxj1FVDMO4sssOOzeOELGvHgP0
IQbajft1LP4ehA9WJL+r5LNa/csPQ2hK/6BBfD9xP+iG073X+GCy15um47/TLDOu
pMPljS5fMXdws7djrZvQtglESDYz3DpDmGSTBHGxVRdfkVxNErHPzB3QwV+pjBrc
cAT15iXLakDM6+HRdWATwHs4CSMg2JBLaK38k+ICpf8g3tnrwt15wcQd/8EUhtQv
/zDiZ9FS75AOeGULYlkoWU6szbbzh2GzkVXAyX9jWaxdU4j5zN18WrIxscXZlrIB
nvqV94pJkyjJYNruaCanUcN6qNAQW+Qf9dZ7tURYYnXfZpJzoi6yjqto3qEP3N4+
YX0J3SN3B/vl3IZRPcc2M7JFau7Pp+O1auwMQGYnzkw5/1yEok9y4mNR8GBPqMbD
xaPNxPuRHEkTH0PRJwlVAZD5Es4MIOM1YIFYU2o9XOZbGiLEzncJPUZGmXynQqcP
dWh4uwoSaKUlsQIUNo/8XJwiVpQoO9KDf33mh5+bjYp3OPaxdjJw/5OkzriJT4mt
FXYOZP42j0SEhuMtoOEvdkDPDS4W8KU0/nAM+8F0ByZzsuIuqEBpH4Y3XSpYHjfl
6XcWbdNuaeTRHCnjdow8oh5NA5FWLBWPsItiOcsh/FJ/NA6WhP59A5gBH8j8RyXG
0a6pV5SRQr0R4Y37lcW+mkeTxT6PPjRBx/owbZ2KX2wlqQ4xtw35wb75656lGntA
62sPcAHaURr0bb3zSR2nI5hnuECh8lW5XYa3PnVPZoHIWcCdzj3lpVn+15vvh6t/
gIekpgjQix93JGZS7a//9K+hHIdKNJ20GD8VWQJ6t5+bZ29GjyorELv4s6Xqchx8
KYtYAIVH3p5WaWj5CgTt1cJ/ZnOxWaoUD55o00wLC2qDLCvLSuDvHfgsFJ2v3OZs
zQtdb4OCmT+NhieruFYhHSvatTrgVTZe2yvAHWsEPDpsP5L4O9ETAQJuu5VPO46W
dVtuuEa1hNgkQkgHqhLp6IT/FFwVR91bUGIBWxIoit5DkmVIE3rsrrLgO9j/ZSNp
2EYe+4LnaGVwAQQz8ZSv23l59hKyJRdGBBDf/7ry3WyQQwXZ4anoGGQFJkuow/Hi
tZffkWWMGnj70P7hni6KcuJLXDdnJEpf6JDdaYxjsKPp1lYtaVy/oAb5+kH+FPP+
XxYN68wtB88jqGzMkBXj6ibzrDQNubFiwV9iNHqqC8eYZVGjpNOYcnN8c/2suKzo
pSpPMoR5XggjZdzZWPsdfh1GvELzolXlbKgtG8YjtKBgshqodCr2JljApEXfQ7ya
2F1hMhZqLAKU0go1+vOVKhCunSXYi053CwjpZjYlx8sJfEBNqwjfviNXmZpGbZba
T+72DE48gOVBj8QM3Ygf2Oh7abH+lZWHCex9uiZKoLFu6G1+1ZsqqQLhEV38LIcM
TSRYwn20pk+3feFE8NjVLNWrKnU1k9NLn+dONKWcehxehs2CGPmK4MNUWM66cT+8
2Va3bOZIqAdYjc3zvc6gTgCQ/uwXP1uWx0jc/+HwSr1kbKOVbp/bEXf26Bk6RtQv
X2d6LCgtwNlEANLFGvGSZeJroz/9+xLVfJCXYEPcRYGORKBLSQh2u7mVZ5Wf9wk9
DzPH+Ayv9F/k0CqjI/nhBATrTC3ZNoFflNx1r5QXZrAET/cMfKjBg7gvGOgIK8CR
WisNEr69qfcy2AY82SfNvGhZhpZizPilrEXOAgpgwWFBOxvfCFjLqbyIrT1WJju2
4yX8JPJqyanHAXG80JfSUVgQLP/OzJEho5yJHYtpUHgrKfPPMuYtL2re4V6CA7zi
AID5BhPwnuMUZ8oK8KxwUZXIFWVEKMfTuPQhsj25nuf4EZW7FFCypoS6dqviE26L
EwAp3kDB6FgOP5/yuYFfjri7YjG1I4j2us9g08GYSlig4Y8y/DQ6R7bhz2i8nCwI
BBNTs4ey/fSRE512j+afcdpTr0VKozDbMVZTQytvoO/FYPTidFkmZ8IWVf+AYdME
jd9ZeeGNUuSoc9TBTw1SIK8u/e6Z79bS4SDWTQi3mOSZL1Faq897S81VScQe/W9j
C4CVq0BXFs0vrIP6oYw+DUV3+4mwMsF9pMc3oKzPyLVliskdZplWe1v/9+SXKqD8
I3grEH8ZznoTlsKvRq24u/aXl4e0XWu3CHTmiQNYo7QRyqqydNn7aFLFGMIjiNX8
UtZbvJYTJk1+S7d8lud+cRbI/S3roSwqDYE0XeeL41DMF0fjep+p16UJF+/UF3MN
azmzalk1Kl/zmJNuVrXSMBQnSHDe0wAN4wf/Z+ajYY+UREFkElcicj5U9ly5mAUR
gu7KAdoJFERb3kr3rCqQIw7aSDRXXjo1umM2IK2bJ59G8e+ERwuGGY7YL7JmYTWc
EqJ7qw8NHYlVSBeVZc4bHaTwLCDIs6ytaFsivFL/FGy9nLCfV+o6tpaz1lN0rNw3
qnXvrmBY2cjXFjzYmATgzqDxVLqMraAhhBiE7TzO/3+XO0BMGPZjP2AAzHMsJYu1
i6Cpw0CrHBESdurEsya8QCCvWkYCRn6m5SHhupIM4tuvsSl20Kq29MU009YiLo/s
Nu/2r9cAcH9afuVVAB61dy1p29dByjSXZGWFvB9Ozl/ko6VMwFKq6wrJNeFOjdcH
to5GQtD3JsEnBlwr/ZC94AhGREHrw9t5huT44p8Z+Er9CHJzdSAveKRubz6HI3Lw
Y/yNkwZ3++OpvFAJkq5JgXKGVH6b1b+hCvZFgKOAcXWzIEHC+XqNYY3r0PEtSuhP
fKVBkv2cySKZSLbuc1PVv6OwfMlcjk/FKD39kj3lh3J27bwdxtMNFa2U83LVQY9L
Sl6NfB+HocXAsY54UkIPRTL3m+e1XAu/Rljqrpy2jgIeAuN3QmxHQs4NfbgjUli/
nde/RDZEAwJFEm1PlsQ9GxYLda3K7VXFIY13eN8CJTmV5DkG0NXle+fgrO1X0tJV
554q9XuBAAEponnasVhxlh0rGcZ879WGLQHt6nh4ZOyqTz8HULHO+3TikzUM7t3c
NfgMiwdEPYRkLeUhAeANZJ3JrMIwDinaqGAp7+gKwjESf/9VES2AFHOx33hfdAEu
5ee+KkA7fc7jkkJ5AlhRAynuKIdaOO7XAJ+qn8+eC+tF8FUmFocnhL80fpobvkD+
c0WA5J0xxkxvkDwPmL+rh2xST8zX4bGFRLROsVV0xQ85hjxdYstmq6NCpKvnJvoB
ixx4qepl+nxdX4vcvDvWLi6mcgfhdqS2gYjyH9B/Wtkrwn4TTwBSmEkyToc3suxr
+1yjUwbqZqGPNqEOF/qTvCyDSkohVC/qBsfdi64UpwrlWHQA8+/IXxBuV2SMmsRR
ysHYvZgcqDMgxcAXM+JcaFzzG/YM844CdduvYTJqJdbxA80ryodSaTqlKUhh2e7q
5jg11Xduj4O4Z5Rc4J8On3QOf7plWgSPDvq7TvKp3C61mqcwGPUCOfF3RcU3sjj4
d5+4jWrl7AbMXJ23HMAVmgktjjlUX/ORHkPTijS46KhRbJczHGNWiz7S6sxUsi20
kF32VzFWwmFXe4L0aRNMUnbPw2ZpjUiDunAf3J9zAsGFFY2OK6rGJdIQfcx1MxsQ
aQI0XC9QgH+R0+RD+3Vfj3u0E+24iimxqMt6fHrb9nae2jvEhv3tk+hpm/5cQYev
HGmfpuDphAket75DUknNbU8CbFbUu5cFSeSqVie/Jsg0G2/F4jJUAxWmVNy3F2FX
Ne1diNpSH7BRNbWyHG+r1w7jdWoS40EFxwkHN31SKYu73B1/rmsIpRHRak53Vxit
Rvdk0yATEhvKOlZsHmAiQ5+7S5ACPb26ce+L/YWzQhpqiiJc14Ow6wzlOy7V0Sgd
UVp38vXfHEWXHVa2OAO0UnRLUwzenCg2L9jzWbhPb6bfoYq+Xtkjaidq3nIVYyaU
nIHE3BWQFP82h2MtpB49CQD5y+TvxmsCw3JWATy0XPxYwYlrrZ/w7D1dEZnY+gqn
zW85kfDjUs2Nm431I0N6C9on6yxGBxuLaZUH93HtU6hmxfa+2sgxaECtG4tQVJxn
Dn3jSpZdSZGso+T6Ord8pkX40sWUOr7YLpncCKYGST6QtwCcn/JFt6hagcHpBz09
eW86CsdYePISonghHZtkka3tS0/NfA3wX1m7+BlIq5XTIUmyiwUvtfBau5MIyL5X
W11RrLDUHBpYSuajC6gsqq/YoRCZoX87iknFVKQP38KuLdJU2mjODwBXa5Ph+t1y
jDotCNg5hFX8LJvUqemT3OQj0iPE1D7Bx4EDM3D4mgk/p42I4E8Lo1/C6EF1WY/Y
Z9PI5fHD5kLLazD+K4eB8/3ndmoC4wmV38FKnhvg/QgMz6x2hSpe3R1wAtV6xKo4
E5L+cwmRRSH5dB5Bj0PBZEQ/F5nT7v06nqnEYkjQFjUuo4XmBttIvY6bA4zhcSsk
TDUC7tFjhqWyCQx1GPcQh00LRUGI9FUXY+PP6Tch86PK446f8YTQylU4Q2GdHSQn
svtKz5Y4VztZ+SfmOamw3MNvq2ZATgqN8kl5Jg9aJGcaQvRkVWm0CtuTO6A2CDXC
HtPGv+VCB05zyNXkctrvkQQrR6WYAxuheqTvk0L2G3Cw4vSA309YKVIg2gW6Idjd
E9wUfrANPXSXUgB1JLwjKMdVAvnD9nNrJ9L+5INkTYJntPbIAc59KUByVrCryaFi
JN2jdypMX+1e/w8zzqDfPWISYX6iaGDSPTSTrmYPqtq3LTe/qU/gUo/rrcm+ga37
X5r7MMeSLEt7gwRGTtoqjJ/NayA2mmw1lxdX6BNedtKEbLuThQ/Nuj4qSp3wt9UN
WZk3jO+RE3gZ63I0+DJ9/go1lw0SNZ3Y4tUnTXSSJQmfayaWzQGLXPDlaOwJIpKz
f8uaCnL6PKKT8+gJ02JHnmOLcs2B2Zs9ZbxmaZ6XU7iHvk2jianVgCrHN+7jGCVL
eQvvU/a5xDCc9kQNgsHpaq98gw24KGHFhQ3IhaKTH6c/aAR+wZCemSeUJFJjWRcs
lHCGgLVAzxfyPZ2HlM/qokBuxGymwPVYZaeGRRya+D5TS8Y9duDqGTNXYgZbPnAr
74VotzWRehVq0BL2uey4nBU9H9Dz3P/z0i8gUf3aZjKXEdlZwA6kLhTlo80NzwJL
J6VMqbmBjFSB/NHeSs0g4p1UGhKEaTuTktInwiIF0NRgYy98Vh4tXeUQlC/PAmum
Uu87ns3vaPRFFvDXBF/b1yrrdPscdVznn0PdiM1m0ZyqnrYet5XbD46Pm9gH5+nH
THTmCTZI31FVstbRUwChfs3h4t3c+NTX0WjIF93jOhU0etHhNX4iIuPyOMfP/LeG
0uYtqhs9y3/2Kjsxsyo5vPL/7zyF5skb9qcVZxiFSnSxoj/08+zPtDNFqu1aebxl
4L32Nh1rm6uVOHW459RDkks7KxEljIN1taj+86I1COUQJDL2VXs/2Woa+SvPzKPc
RM6U3byh4tvWQfkCzccD5iSQd3vqtOX9BLHcGC+fgHGihDqi5/Bpg3WVlDBdTIL8
x0xr+ftAYWmMxzi0pEGMsOEnjwP1lJUd8e3KVIH/DHOwrFcQNh1w7ZIkeqXIowhV
JFRgzT4uuFp1iToerCzMd6wHyo50iqpkl1BPztwOyLPrFZEdmDjBwPYV6kmDBNm6
sDWuChN9xax//oPYWv36ZI8WZwLZRsCxu3nqqSPAwOlPzp5i82n66oZ9I3OaMxGE
VJIGVktKAj2MzpbL7Yi34vXtEyEyhVVDpMXvtKiWo6KIo5NalyaeVKYNJv819TCh
5wfcY3KN+KI1LySmiPAJxOv+pFanD5TmIJXi29WzIe10RI+MmpzyBuYREsrSSwtH
5CLpL9gJmf0AiX/cZI2BrsuDymo1XmWkze/Qw2HPk4HGA8Dp6kIertHTBL68NTYF
/hZPinUTTlFd3NGb+hA+0BG1NB7cp4JInfF55wQrJsMw8h3bFX1JbglqaD/BHGT4
lySGJmEfFz5OYddvTJsPYDASx0frSqm6cSBvfpxptn9VESraG08DPe4VL7yB2Rgg
ZTwCuy2bRnP1u7UAVVvpn88aNslGeu+l1szTzE/CGdri7chTkqKtdYIspt7a/EBB
HREPgyohpxr2Qz9oKXKcuK88KxBJaYGp2L7/RmYwOEt1d93gHu23poeFX54MtV39
Uzaj84XE5VH+kUDzbeZ2ELN0V6pCYrRYUN7y5WPMNvSj6iU+QKX9licT3yZ9/nNS
ChJDIYFx/Pzz2+0kNxM3NmI6AZit4vTO4xN0agyrnvfbevH0Ub5fvCoBCnEqPX1E
pKkeriAUAGn+IsRF6dXq5FkZqUjHpIGqPWfyOaDOLSpooCVjcLa22p8tCqkIvzRa
ay29uRrD+PnegX6RmgtuQ9u2JeFsfw83o6RCJzA3mRubgm6K6R1DXl3v/AYh4KsR
otCIhJtdEPiRzrPeOli6ZuKR0MvPOb7igs4HKF7V8aFSDFymsjGEGbBCGEu2dQUm
c71jMC8tZfAiGdhce7r0Lwb0AbhH26iW+aUBuqpo3AUXM+NKSgl3qsdRqZYxKWxf
4how4/ub9tGY6DYwrkkucjlNdu+OFcOLWp3ObEYEfNJfhoIYRi96s6/SzswxsedX
f2b7V0IlnELWJW7K7wecj4FXJkYPDjV4qNO95zNS22t6po1fnAu6bnNg7NQKqFSI
BUehAtlJfPUD8trArOWP1yEaPRDi5Gnvlj3WFMA2dqIsO5cbfND+N/Ug4TY4HW/d
XjvVc8PO/qdlWFRV327M1nUhGxmFo8c4/0J4rYqMP7Q6YBj5MT3aXf71MlukLJiZ
gKjj60UMpNDB2dkTN3p40pRNVSr7uRW5MVI58N/y6EgMcD6aSUb+FcM8KN8LWr0j
kmC92wMPdaB2O83TLKMBXJQ4lTqVl3P0X/xOxqXuSTdVorXyyGjALT/RgEuCvHmd
yy/ZfxTOaeZcwgT5wM7/5z/GTYfs8DA7eXJRKeHwNqhirqVb3sw4hyDZL/j22oVr
QpI14lzlIk8SBGX5XR9bqL3JS3V4ra8QtCPYt+53u5Kp1HZkxkEXFQrPLw7Va6R/
StdQ+VlYp+FGWVaczJIE49s8JfdjHx9X0bRAXLIOrvi2li2mLGjliviDAe2svTlR
OWFnWjuZmXfC5zDyo7CZEIPofN6UcI2Jc6gmWPtN+/MU4+o4Sotia/k5DE5xUmYu
RyOCC6+7c5UvPevgiTnL8Vnu3uYxNsGB559PunxcPQfC6BzhpDwib+KhyR0hoz5L
hSLZWvh6IzoJRJZPP9nvg3OMUntQcZiQu7Zz04dBbV/EcRtjbp8KOqW3nFI4wTdA
JhCjahPUj9nGl+jeG9gtzDvo/R630HVa1s4Rgcv+5eiSkblKOhozVAsjF/GUhGrW
PdZk5LJEMsNf+NsYXorl0EuXo6QScXK678QeDgI7y8q4mZ0XP8OhV/SaMStg7MLg
6/lgl7gIkMDYdlQIxWNCTcD73tWKu52wcZOm/TdIzbRK4d3jE5rRW+yDJRQwGkrM
jaLYXAAJJN+ry5okOMEhTv05IzrnIyrByQ5Dp3DsowDoV7vF3XzLKxOmfqJu1v04
CgwVSJ4bbAWO5QxbhI/IeKcWLic/UMuVrwS/E9B+kREMTIbTEFXoY74FvAjOJOrw
j3isayHGfkw4WtF4tfiN4+gHWV6JiRBydbHj0vGxHccF5s4XWRnUe+49gL3EPaTo
hiLaGpMOKSvS8E6RPko/D+qYksD5PS56T7SyomLvEMWQOuRzUXj0c0Vhg9o2+bBh
oED5mhd3ZGR/iYBW0ITOKJo481POxb6kMgblMGuDTQ9+0HPZz+jpIYWf0lrH5zIX
48t5HkY3ZBPbsyYNmtlvxoxFcKtUaGCau+1J1Vf8xHIS9+VlMZ746zUYqLlCt8Iz
OJ4EjscYcjYsmbVBea2aCkM/vyvr1FWRs84oEfCLsiIL4Oh7j4TENKYCu+4EN/0B
DrBAAwhtcWlhuj14s7DW3xzppDOgnhIoUH6j6Nn2DJdGQgU2j+BWAXyV5BJzy5sW
Rc1nHn56vTWPWYN7dHokOs6g8J3QJwkLIKhTUBAAPj3ORXOlNhUSato4SWT5sQfb
fp6eP8HXE4h761xUVEPtP6Kc7m6WpJwmQjaivuOOTWo54f2nEVJF0EA57dHdimQ/
0ncQc1SEbYGwkOpVYyl8ynvAEhsuuFIJVsxfVMuruRL+rQhNk5xyWMENp9/5VVmV
/OfhpLqwrzWUKwsh7GgPjS0Yk3IHgX9sXAIZyYzgHoffjHgs35DRZoGNjifj3GRe
eMnIa3DrH576RjxAYGY0InxLVndZoYeWAhxyef8G5QYrEv9y+I9omZjcIexqZnYF
5/5fQpf/Eu6zuRpjySn/hQiEVCUPkH5+zjh4Lktox/6SoGWKR0QLoDCrlt2rwUcc
VURSG6GXVm3H4W+7MZAhwyqixdoNwxFPuSkVv0iAYCxwIYsLPKlEhXh0Ke3nPaeI
+73fNeoMKtbiyf8hp+AjN6xkM8jjB2nwbg6SVrq1Icrb16pSwv8lBCW8aOOLPs/a
/Oo0M29Pq+QXDsFbxAkmd9P28jETPoGMYdGf4Q8Eaw+UR9EaRYPyNKC1Bdd9Mhd+
85n9UWfij6K9alcKcTakMl7OrvdlFuGg3JNUCCroEIuNjtxgAD9Nn+OhB9lciCQs
T9gy6Zsk7Ow0txLaF3htMTTcQY78RhRYnnGCGbxXDrmCBKnYynzMYeDwYpe8fV7C
nYKOhdlBeZwJauV1lF82s+qEcRiuAO+318bxHQqbLtFH/8Q8K4nkfoKTpawUCz63
OA60b3h4HxFhXCBJKYfPyz9Sgd84A/+R9rJqKlHcnJ2fBu+GppnCBziitiY6B//6
a4Oh8+70fqZfImaSVVCN1Bbq2Y2JOVDpe5hd5CN2FBhFDGAFuJQIIgHrbNrUDnah
exOtcsG079obS3dTgS21Onp7o1SiZ48CvXbY4a65U9Q3W8+knH2l8FxJewMILMQO
INeOxDd88mrRiST8Pa7vmK4e3Z5Ql9GUB+3JyHt5YQ5RBHw0qHCQ91BbDnsKhxbe
wCBhZaXdJCcLOTjSdyAkep044MReBMppHsIZ8XVVBTCPpC5MlCYcy2GLpkXgHeNW
4UmhaijKqy+fgxQ1vlKeG67dac/Dw64l9IDBqRqGQtKB2ugKMEnLRBI5wIFxG8n3
vXU8CQ1euDZUpMIvH5ujZJwYrlctXkm/CaGDw+7WHhXHLeXQkphRULpfMJgZOVXb
/dCG8gWh7kx0B1rmU0PHmTmssuU83M55aQKa6x9TP4TfCD6c7SygfpsgSMbuuexW
nwAjLw1ANyYnE+j/7fiZfQHmR10HCcQqt0sH6HF3fW3JlfdsNGI2VjwwGQqZNXxd
lJ0LA4Xq8OwrFPElJwCM23lDE3XKQvcdO+Wxps7olSaHd7to5GMUYGTWdT+aquoe
+dow1/wmNkaPdhWLikgu0Kgw+8imjSokNLVcPEMEM0doQ5r8Hv0T267B8MDYdSGX
0PGGULHPLZLn0VK8Nw7TtufmeyGt6Yv7b9NsA75nJgR7QFL8j9tvzRTjI2XaZ7NS
UCt/Y7ymGDi2X+e0OKSlVnxGdHBs+4EN6q3/aDmwQ55i9jk3as9l3Z5U8vQqyoB4
BC9dkqTNUzJHbTkP28nspfG3Sj0AKTZYTmk+ASDPnopKe3uP+rVFqi2KDXEyR+DL
f4qQsd8wQrDYYttgny7nhDnz8Z7OKGaIN/aWPktRNZ04eE7HsBNVWTaO5SNTt1Cl
1AkBZC3mbUwPDnEP89cFkP3Y1gY9Bwc6Cs3Fju5jKVdAJbiWW7AaMwl5sc4r0gla
ig9dMlYTjOGjq/eaoMDOkCsdYoOIIqklbJVF28zGg+HPkKPt9YvcXxb3VGv+Oo1f
oW/QoO3kF5zsk7lknzabbxK/h1hK7FxJVwpQl94HZnSjmjzxdXG8fdh34CkEy3O6
lA/VNIJLQXtH52LiD/0qRIUtGY/zICWxOXI69ivACeg6o606U1Bzz4A4QZPT8afN
Xhu1VSjtXBBh4duk4XjPla/H1vIHgDuLDU4bZDBHAA3MrL4i95rPBd8DR5iB+XKr
jRjk8kirqCWP3geVfz+GVjf3tuPQ6B1lmTiQMT7Ed7446NjbWOO1dSk7/I0VlI+Q
YGhwLXVTmVshKjQkGvUrkYz8aLmhzL5hSxsMGezy1sXgo6cLYt/sbNzt/rw+TDq8
2U3V8bXRNiB6cAz7+/jKS5ZeN5Dra9vL86yfzcERN3/EQgRme2yCxxVrZsWh117U
/BKzPgbwviHp8QKTKtFiqpSjydatID33dcCzdgvHP6HxfT5HdUblb18gfYT2m04K
GnMbdWkOKzjKz1nWi5PsZm7Y08catVoXAbgEa1ENIQsDlFdl7SyUIhNB288T3sIU
MU8cn1+7WVRhL6ML3NRXUr9Z7bVeWKTpPbRLkHLyEhq/X+onCHyy+gUfWCOkjMr6
vXsgD64KTgPlqecKNVW8Z4RrYN6gSGIIasAOE+YX0PkSV6XQkwlkZqGPmstd6Y6A
MjSZyZbCNTqOwwttyz36DlMRjUqqFAiP0/uJ6C4GZER6Ltq25PM60f9prrAij4MM
c1KOeAHQIY5Lkzquet11Wt8Oe71viHvV/mLhd5/xIXVbgteFvw7k5Jo2tP3J9KE/
Jo0v2dWpejpALd/g0On3Kg8nGilSdoZZ/sfZPpof84oyXejBeGioKxdz53PawTHz
uCLTg9Pff2a9KPE/J/lPj8dl+TGpkJZnpHyzuwKwsH7Zs2+4hnt66cbR4Ikrnkcu
ihDUbQ0Jd56v3JrVIl1aAktD4NM0ueV0x8ANcZdh5QUYiwE/Qt62hyUC6iOgoBU2
nbInuIEhwNVzdxmmiuH4LtD2QSX5UE+D06HLcUSfusaW/maq4UIt+gBoTkP8sYc5
pKy34QR9gRqMz5x4JNQfM5v6GnyK5MX6M3dkyjxU/eVlqJk2QRUKsHbHC0Lg5SaA
Aj4SQyqthfhPfqYicnpVu2Qn6zH2IOovU6eyDs0jtQsxQBzvPOzBtTWPXJh2gigg
o74rGxkvB041l23TVHb7H5NVyZQGwTtKJ+0vOueXlfiAx7g7+A0i4Yev+EIfk+Gf
tR+/dEUUpanLItmHOxFAUuyQP+q/2ZegmhjiRSlHDtmrZ222LjJfiTwSK4wexvud
WgYeMexRSms+z8J05jkrW2UKrt+izcqncu1yRRk7Tifl5Fr8EAri18cbUfignZhX
JFeiVloQl7iKx0AysRBwbEH7AvvyTKtimqq6WMHNaSKB94cdbnVlJA93GUbpCyi9
Nx55KQc/K/UoUBtdYHGIxjAHDKmNLQqhXw0Vsz4cLTH7waVV0vNPMaXrJZajYNfQ
l1yj61lrseWbXm2K1lSAIYsuSa0ZjbyqJhjX3oMfmcVPPLCLufdonL0UZQ8lF3Q/
0aM6/w1hEqRJttSh/WlmQgyEGrAT9MbRlffHNSYsDa6xn6V9VRD8fwpWU+QO9hlF
yqDs0HWnAz+fWO1iyB+9g7WZYYM6shCquGCdsmS52nsMN6UTjRN0DhLzUdNrLw4t
j11rlxTgUXyPbdcekkrVnXG9mKmxJiFroRFowEv13ersTYfCq04duIjkqUMLJiSq
GVV+JpmxBijSIJgmTfbc5fmSIu5ELEROzRwLGhLMdBH9q5BFGZv2zUE3aXXW4VA1
7WSvwbRAlAdZVPsm1Gwc9GR7c+EePp43SnwP2mphiUWnnUtXs+YFIZkcyeTOxd6Q
KCcawEdZR6WXYyNuUYtgn4Gvg1cemLoAmnQmqBixzvUbxarYz2og665ZodTmulsS
7+WsE4gYDLSp3kZWtk479V+2vCPbz4NDQXpUp42EZjViVewA5hizC3mhbW2mL0NK
GnyeKMaYWDPMwPn9fpHlZIhpy01X9X6kwEBiXQ1HiZw/uvAF8NH3KM3CeGY4bmLa
w1LfO4QjGAf3RLBCNIWUSjn2ESsgv5IuftBPen9Tqcj5TlnFNovESS7jVp4XTzyy
ZJlE7LXGEwLPDf/mf9ke2OFnME0S4vdzCKQyKQWLqcC7rO4N35s3QGTgonsioQeU
yKooCYdobWIdXgPA3S2pe6dxsS1gZoJnh7G602s+ZQVRWBe3uJnIak3lKyKpuI2m
GYMJBoL2DvNwvPUoLKG7lNZIn57kkRN2jfy2FM8grp5gj8QQercmk7emfJ8suzeO
8LEHVKeZyRzQG6AqG1OGLCLOzAkJfUIpa+LLsV3tSJLV6qpZV9ZH0nqvvTgs/V0X
fqPr7lIX5jN3l6QeeEYiNgTQ9SawbdPoY8C3kqOOVC+lGRxg6thgU1qc2qAK0Pi2
KzGbG3DkKcoh0Tj+/U8dd7Lq4lZAMdiatCg80thZkNZphrTVYv1xO+2+XxzY9MI0
3yN6FoYksHtQScGnTrrLp8/mxz7rU91KZMLalrGuN3xoLNwkh68fzsm01m+yJYMx
gZU5xR/ycnGzEP0U9QZlhGYX6YckRsIgQ0JhfPC2zbtq2ncrlfrn7yOuVG/dwvcf
lWhDW0nmsxX9w2WHxKkov1TdcCZsR4vrCk8fDDEZIl7St2UE2HfMd8cnHKWDFiUI
ir6OSwZHW63CW9i14AZcx2OasMNvkkSGgOZZ3kDTgcU1sHQKJsmH/HpKxq5D0uUJ
UF8mfrwoYvanpjMsipyoDSYOm1043ar9X35TQnXKxpwwU1oygzVWYP5Yc5Dv+LAD
slc/eqFJPM4AQUAHtM80JHACITFh4tu4kofjfAQ/mRcvDVMxo+Db2BjJCOEiQr1j
lXNWRne18vuDk+E7AlzRdRjwmPeT3SfvfmUlCnudr5CH2rBXjq2n4yqftiU4DZlh
6cpP0UXPQmXbWKEhBn54YNLuLUnoNX4ck1NWnbaLB5mj8FwH0DQr+2WXPNRsUsAI
8BRJqvGg1TNzY7fWxOD20mvNdxYca4ltfZJ+mYsFyM/R72ocF4ASKZ4mY+JquqFc
hEQS6BzAbQX24wj27MUodxMz2UgQm1aVph9j4f2WAGBHstWWNl5/6b3yXY5qrejQ
iil2yI343GrXPz7Od/JnejdYyDLCNTQA+oiInVGJepW2pyL+mACwajBjdcpTNq5/
PyeUIegxMUEu0IaN1zQXqBHzQOH7c8fcyHLOWWHr3vb5G8dky+WYsOh+Vxq31afp
1vKq0HAWdguL7DcJfWEi3t1PzuZgDzJkKnJcyrrxqn/QTMoSOQf2j+9lVA2zrnT4
yLxhWKaE6VxISjfB32TLHYTkcw3LuTdsny0vwN3HMc51ntn9omTkNHCxF3WpqP2+
hfpRu+4XoAnXUq4BRV5QVXg5RWMaA6mEFbK1COGWJqSMGJUv7PwMc76bzCt0pDHh
jYS6AcGqaqtGLsXVjjccLursyTtd0BC4eA8x7a1BgZI0+U/lkAQfBBYIkqxzmo9O
WAq0HeQNySm2x+J9+OsKyX/YObxsKmfZfmEY/UFvR5JtAAomVtPa7JqzlwW0iRfJ
Kjn7XF9Ll3KR1gLhS/0IlhDMTYJdMxrYf0koyveodsP5Xta++xMwZJBKvW+DlOPS
OYZfapWNADrDPPX5GYzdqMDATrJ4GXamCNfUBlaL17TxW5dG+oawMt/isDKF4SUQ
9/2DidFnn5ytpfox2nf4q1m9M/fT1cyMgC7rdZufpAmzMBiGXDsSmhIgFpH8wYLG
UURQA1fetSMZXkyJsDGGZp/BLS9no71vwdhyB3lRyQMCC4qlYrhuftuRNDrcAguX
y8Y7dppB45u5CKv9T2Dvvmdn66NrHTgDX2SZcT9/3as/Srb1x9cKzAH0NRLedIxJ
L0aOcBBHhmJjY7Q9/+rOrB0tzMIKzqgU/ttDVRw9sCe/s7O+nUgxrSHlykGqXzW3
sj6MRg3Hf7r+u2I9iRees1PvuIUZm07UU0H67Wi7mlOdVlrjJDaF+FN+bYCz5s/1
ErF2oFFWBMZEBfqVm6/VBER8/sUFJ73YSqwO0qF9AvOFAm+12+MRIsjaKgDRVggg
kBxolQ6ADdRjmJeF+96Pdxs0kqL5DLO7k0HUuAwo5koIu4fNHyFm7R1hSRDGLCXu
xSQHNOMNp3ItCB+sJIWhxvicnAHMfufu/5HinZh4W3h7UZ6yYV4Toidht5AA3iHe
jiYt9NuGmxi3aBMa5MlPEP0+korpMP6l1+A+NlYJGqtH3x9zjylgXwigRbpM5RTo
0s2ttJhWihD4rouQSPv4RPeXKYpjwEbrl5aJdcw/xx8DoxOyX0b1JXl4FjbA/ZS6
fcl883bLYMz3o1nfDjo0JRbEyl4ZZnUarZGwiy6LtJCMdzLOcIzeAd7KertFwEnV
Ug7uWMgpSztJTwG94BwOaF4Td4tVionR0jVfNV/nNj4HfChxjI1/F/HhpOYzRrh6
lAlXTKEyNC8Haz8glgGoUkWRvSTw/XJDuLOlZpm5om2fz/lSJyJgKT4aF3T8vS/5
7LgNF5cW9LpJ6lCWl8hOM9C+rvOxSIinEL+w+KD/7nh7qGuadgNuBRbOhfY6oyv6
pFNqSdie75EXEg1DomCV3nNcEoRpKWmxXyNu4cGIKVA0tKFatxXinonSXUssUCQW
/AQSo2yesq1Wx+lnN8b5qIu13RqxGRJstu6ky7r94xelMgbNnziV+Tup9dVqzvHJ
Mq75QX5G4TZLae5afgnz3rqaGnMe3Es55jtEl6QQ6jySkWsF1ATH98y/ClovFxrW
lS/UzxJCg0TBXD/MD/4iR3VDK0MVxp2089c4wvBy2x0ceOX8bWfZ1RDOly9rqh2z
LPwRKM5ikAicKcc8KQ1njWYGI/84wUvcsZhYsKp3kE4xdd7QFO90hzjgpgbarE7S
sslKY78WYNPSX6Cleg00mCtg0L5GoqvuqtOkLwOd6CEQh4CfqRicJYUuqRO64EDl
uwoRVcDs5P8Rjv1PRTCaAWtLMd5GwYsQavMPqawCzR8YATG1ThvCmDHMPJgwbJQt
hT+tRHsHhgmN6Jj2HnETnrBsymEgURQPcoa0R+EEkEGeDYT1iaZH/0kY45HIVnYB
jy8w0yj95h6hR9EKSZSzWvEeAVNjaarO6kmw/HAWyxFNeIqyoKCEwzx9gBeydOhZ
cKKUtQMoonrej+e8Xat5VAMvkzZEsuQTuQlkS4HRvPyCzIqYJHc2MHVjQyPJSWLL
k9QcYZ3sOWFAoYKINNZwBNgKIem61MjpQ9UsylRlLefvUC2eCvP3N/hs1IE7z7gK
Bn3ljj85JCRi3PVgS48bsj9TRwbcJgQfFS79CnsYRv5XP/uTYTBrGWiQdtQ2GhbA
mAcVAlUAyijkM+bCS5xKcvMvlwA/7wT/BSTkxqwWFH8pynucDG9Y2cTGqcaPMSq/
D2BTbJb54FyCsSqRGFYsSSj8PBIgymLLtLIun6AiAZ+b2irEMn69768Hvpn1Kn/o
SALkpJiOvwfhXxETQCBGWogEgPQ23zopcIRpC3RPCjzSw3yHiQK6/6fhmtiJz3G3
z29y4Tq3iXm0oMWf0h59WtgmuKJ85allFL0oLHQ7kMXrfY3qQJual4/qYzvcnLI0
qahs/qlT/Qlh1dGK/QpUv7aUldjGivHCJni14rWammV3MaEB8+xPZSwfMG5rY33v
7dyFoirx0HxZ/bIVshcfV1dOjK+9Bz/ja7d55PDzTUKMrWrfTFX0Z67RuUucz17S
9rXUC++jAN+atW9/UXY2oCbzG/yFuwgGOu+FPNoq2n1OOxnsUbxQiPCCL0WIzWQh
RLH7K9xkjpap5M7Ysiy7mDNggTEy6+J7Y/lKoa/L6SEHcxNpe1ncXwy62S3aT730
eCIMzrc2O8ybSEUQNhFio4Yv38mTOnpxYfxASLdtnCujU5JAdoOutKRT2RaNKV83
3B+FW3Uk2TtR5CgruJeVIYpr/6u1KdujIy0dqzZqXOr0T/uD4WNO8zdVdWedvvot
o4NwJeGg/uowAxDXz2ea8EcKmwIJbQH/Wugc8d2xwJHsRYqkTxbd3QRlk+hQu1uZ
OTMt7MXaVU2y6HmGTCSaDj7ot/eWQa55rSKK1wcUm0ZlWKutVIq3oAsD+F0Ind4H
sg0Nu+1SGnWHqt1VioabcSgmVZM4yjVeuS/XiTCzQOEBkuRtybe2tzujBeKW9RJp
aWE2tbWV62fP5QhqJfH0ajaufQDJhYy21RRq4YaUsziyNgZmcsVprkVumbH/uqOr
NqeSyYemE42OLAdASTOI2KCeskMbTnDXCu1+1Qsg2y/1NThr9vpEgla51k8wwy4x
uZtmjbe+/xYtt1S+rcilaqPifcg3eysRHTvQsPsnSKfcmIuC8zEXR/CkuVShqTIp
lkmtoZSdSWJFiZgmqZ2scesmwLsohI01hprwxrhNzO/hCKxTGhHFDfUIvkkKCRrV
ywBeWHGd0dqZh5pU9rCfcplKiUiKBUvafSpWlGjUA6Y8s7bZWT9/IcuGcurAtmh/
WlWKCXPAvxIkCNF208oxFMOW83O6AoNYbdzYz/qNMoZpES9cPD7HkHKIyitQEwqT
/HpsrGo+vrZr9cKM1ZqBcF0V6mpufAnnfObLSSb4YLisUvYisGhOhGI5nNNNJll3
xESyLVO9h6BBxOZPeepa7Tu3cPgMPY4tq2nv9l3L0G+jDqmibQ3xAiCtFXAAP3z9
PBiQwLOGgoExP7ok9LU2fAwKoNmpIqBbPZQ9DeAyhtPqehEZYO9/hS+bysULsADL
7yY8z98j9BKnY0YFzx1wag8+4f9qYAUGpLKjq4y6M1KSM0dNngTN8qAepS5qUbYU
wUYNQjkNjM9/u5R6H0CHqIeTjDCbjjGUL7m4QcxbrAh99F8jA4/zcJEEa4Mic33o
0M4DcOt1Ghxj1/mkNbzLSyQ/0tDpbOk1+x5QTZtU2FHQnS/opcHDcZcv+aDo1tlT
fIjMy7aIhYXRg9PWv3K+fPVxpi3wTM+qnAs1PP2JALXTzJqwIvRKKts353No7jCI
tW2T+PtRBXRUCWeusc6kAdZO92JP2Y6NTvH3ACfaf5XGK5I+yN5xwswzUQNH9cxi
gWmQbgtde91Llb2WgosEoZ8+9zNiEKeeYUXbs5n+CX45tY+vVZ6gpBoQk4RR7mSu
PGjFW3ewYrA+l+bHJYZCMTb22zRLGZj4VwlwKyfPmycL1T9ShII8xlxhwj/QNmoe
MkwG3q4GHZqeJ8TSXwZewniEDlt4SRcVsg4r2DpxMhQKSOhDWzvF2broOWFrCOTc
oJkS79hcQBZUFz/BgH7xbKof51yf29/1Dj4+vj0aSddwtA5WxsfY2vN7qWR8IP4G
MZP+R+pexrrParjyEQFB6Y+RBeyJOvR/ULi0lympt+oWJjI/5eVid6+w1h1PXa15
b0B9UjwWaye2xO7ClL1J97yqB5aFU1j1tYFqiyIs88sYowyWFt/zffUD+hJvEyFb
EzhGyNv6AXtTaW1y/8jd8wdTUZINnqoyjmvAAQM42jBUP88ECPHAfvOlumk0vZ6B
J5DBrwQ80G10b6usa0kCcn8aMYK5UqF255MPgY41vhp2FCdlvpxEYr9gWJpUz4AK
FRW0VuGrELHbxhp2qb8IgWwlHPbcEpwJKWt7eLhdIjjH6HsGJRdQ7gKV6Yr9kEl+
u6s9ZfhaFyUYFT7Ik/9F5yOujIikFJD6H/JK01H42Eo=
`protect END_PROTECTED
