`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
52qPXAXD+G3bX0yKs/fI38jdQH9MTKU97QJcE8SpHMgpbi5lhHI0YI7aTh2Eexks
Iu0vbzr/dRykjCEpMNAk63JKU3msm0A449fQrbbrU1HXRprN6lBq3z+jm91l2ap1
vDuTFAiy67C/BdKby5GvXVl61xIdCtT9vfMiYRmUSwy/jFoPWIwIw0v2q2NeJi2q
GniLbLxpptI9DYkqUItf+OEHn7anIaYGoJ1Gn5BFCZg/qScREpbjxYlT92KmQqOH
1H1DZPt7wZ16gKQ1y7Y07N0vdh9mNACFJ2ZBTTkd7P8Xpp/vesEfi0JhQZauXofb
LpsE+d2NzoMUItKIPtTjDDl1QmLgxHBONJzTd3C756iADTkaUK045R+xzz6lmfxz
SJrO/a3w6iJzMtVyCw4vSSP9tA8q1gXUPIsEmMIlPn/SUaTc+YhN10InTWD8gEjH
JT5/+kwyZm2LgHg5SF2EQ66XqIYu08m2M7p+2l/L2zLg7KFDwfW6Y2JKUnZONOsH
eD1UiGhIYCLs5YJpkIbpPpzvU770N3uKWmDFbBC+xBAK1rWDkJJO5ln9+KgKomZZ
zDFnX5hyF+1+it9Ja06Kex5659rPA0ynUeAWZ2ZR4F5RQ4BUEpaj1vIduvm+seRk
1g7F2cxjaAuOwSyTGb8zWm7GfAfLOsV/grh93y2oAQX6yyDMBaMqcEtQfAu39seU
v8LdLxKNj08OMhUaQxngAdwqTHt/vtlJhn+eFqdAh82MwzKMSpud8w+AvGR6qGhU
bZ8777cAyTX52wJA0e4ormsRvvDJCFYdJq64UB3b5DtuSJmMUJdXvVdd0BylViyn
PhMc9fbTxwWPfrYmJxSl8qdH2/Yc3PtNF0FLi/wMusVIgcqBf3MTn1QwNWsUYPPE
C5SQgIo/SHJYEQBPN7BMEUpvfYPnSRzDNQCjwn6yf22Li52mue5MdppJirCMdtKT
5V3VBrGqJlm1RPiSzwMMksNoODssKYyKnIIoTcoIm5BLXzyP2kOTrldX6EDdLq5q
+5nG6qYfu7A9YApS069vN/eYh30XD4y6th4jKukx55JEkYp8auMZOO/I6jhbJxsC
tVHKNitRPFRkdsDXVuGUSE0auUqRm2+dQOGNlSut9Lxzs1ckj7YlYbcCXXImopdJ
cWfriFuNEHnX+m1NjFskyp4Rt3auZcvmLRyPznwxsEc71gl72KcttV0fnKzEKXi5
zqllYke9HjOr6bs3mspJzywNUuRLfLJy9xOCbx5oBgBCo/0FSjG6x1JJhcZ3LNT/
1pOYScCeJbdEGCcBA1YcC4K26dmJ0TjUkmsRSMWSym/GCaWUUV79BJr6wJuFx0GW
C5gprTgYGiyI/qxrC2guIDaATJoSMemyFw5EkiGS2woOQeCx+ZQmYjirW8sjynLY
XznydBA4dKMxfr3h65cp5S2P+p+l/9XrQxX4+oltlZtCZuW5sG6atIYvcJqVpSfa
IUBCZNIZNm6j8+EsL9q5+iXiXYUzozD24owbXMJceOUkZNDfvQOyrQ4N1+PsRFm6
T6dssS9/xMD/IfxwdFBVM+EMYSB/m+02MJ8gkmXzl0ygsw51fc9lD3jJicRvvyev
ywpzuhSvJUcAow/QVIw783QXZZpbgRXS0yvRzReOrfItQA34Qp5MZhe5ysYYGOHc
ZJlBBt1B1HzWvtdYYeRnHiV7L13yUx/cGnP6xjL7ADI30ysPGrae8N5f5GTCJS8s
bPn5TeJvlwK8xEhgRgDEp1ZH1G/2uBLJaO9Kvc95LdDtRg9FpKSfuHJGScjGrrQm
cXHqBz1p9McvStkWSn3zX+YGKTLSky0h/+7265BDir6HUXHMo8CYIgE4UrMMd6R2
PqWhttPFzr0SLO/JTs4jSeCmciB8mb+bbVYn4bMQ5EHY/P/w/fx49Jw3KOdq9KgW
9gHFcID3qf1Y+x0J5kngMOj8MJRBcg307Pt3zrxMWhOmXGz7Kud4k0Q2Lee7Fuv4
40QluOxpWwk6GjazxN/E28wjcQhBK/XfwIyLWNpAgEvFcniKKb5xLs2eAad+pRdN
mBfMFKiLS1FdWzKXknES+4F3813Y2TM13GboeVbqx4/wgVgjMnsCwInLXyaD3Nwi
h7ab2oxn0Opu3hZwhexZXNFqSIYavi5fU9N2Dyx4KOA6/49oIGyurdDIRt8Y/XDT
vd6UTAfJncrs8io3HdUjSAM3iDjiuD068k9TZarDOEcOJglFxmoJLTB/+KbFzZ9e
e8w0z2P7kllxeyWsRVGeMWewsg0AEn0XB3Vq8VEsPfLjZMoACYa4xZcBdEzjabAM
73LXOo4hFHoZ3tIb3pDMYG3Ln54tFcbfpLKgSzholytov0Bn+09l2gguwQCrLFRt
4c36eJTyKmoHc7wRVWkxB+7MSNjODpTssQRLsimf5MqChr9vlszxwu6YotGYj13h
lQ7OumG/ZzA15pwqTTe6sIq+cZb4ZRmJHA1VXbrYNcR5qyh0Dj8prp8J36Bc+Xjg
iJQ0Axzhy6MSTMmD24JMwIXCXCQTkFz3mLtWb6tWnIMd8IUoqlhZhD0c/1g2MIvT
CpNmoLuoj4QWBiSqO4OuKClF5vJBltNYaUYqg2RimKWcN4ECOpYOP1zTpztvvNdq
4wDVA6906s2+NJPiOCHQDto7ZitM4AtwAWpDB7Dvb4U1sVElQqebBcMpA2hXMgy6
ZATqNi4Yf0yx2Ex7PmeyVBoeqVGSR9q+zWQCvckmXTagHx+uAhvuem06pUUzPEAZ
zwxtYJ5uFI8E3/WwN6gVypcicPHxlzg3gRf1rROIdrNfRWYRohoXjA0OB4CyJ7vk
fWPVWDTthhw7wrcsStzcpHs7eGsG5uJ9fyfINTho3QF50p3g8p/81/j/3gp8fG8a
8mrmBttcRxoUXKnECMJhzICAnUsFjIWEzNXMEQ0/+2PHFzad6nhq7Eid5E5Bcvub
vLs0m7xiasrWVxd8M+/L9zz5DLtqMHQ7aXdDrrz8qTUIqEBlAqfo0DlZzKygTIPq
MOPNTfyCDqAbnR2rQ00MeTSokXZ30Rty4zvBC701eomLCPR5WLoRCLegFVoKYbhH
aFLnn3HaOEsWgogWaAgbQJt1ynfTdHCj04XghLaQTjCpsdy6eHmO/RjHTXFcAP1Q
MIYb7Axtbxga3KGkVbfR61q4DeDZndpdffKg2txvkRzHOq+fs1oN5GeSEEeevHcE
3laA/RfMr0bo6U1hlj9oGdOeQ+VVeg3W9m/D3TmK55qmVlqJQfAaj4nL+zViLO4y
dw+PmdYSAwt5HcQljqvydrKHJvOH4VH1R6qWGPZBwpS1+m7YVUmdarzQAbIM83jp
r52MW17xqUbwcxSc+0ahLL0XKpINYrOo1hallCzTBHR+s+T3uX2FTBjiAgMlndQI
F413eD4ZGuRq+IQnt6BYhgFCJcuPw8UZs0HQQdJgn3bnIFIOTDSa8mHFkBWJeOeq
3PWzw39wbaXfjw1fBAZsg13T5yOdI7FyKTextRlDBuPXYfcXS25phnNTGgwqOR+I
4PzLYA/LjJvtH1OIl98TsJKSn+kikPnc1REVe0knlA+9qRUyESZB6eE4yKy5yOtK
SDrzLcDD8ldXupVhwNdb52bvORWsdHbenO5fPujhd/q9x6OnaMbn17kAxNhroSqZ
t+HPuI3ByGALptWm+SaSP3s2dLIi0bKEdoWiYAkk5YFwZY0LYpwX/P2/fGg+gN9W
zIQFl80j38nF8P4k1yyaZEanUyRR5aVCuWBJqyWlR4T6pcjn2wTEcE36bj0A9qtK
GoGzx/Y9mWzUFwVBWfkB97V0E8/KwOJxZa0JIJ46gm0=
`protect END_PROTECTED
