`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ejLzuG2lxAODYL4++pNs7buQwo7QUuNP1ym5K/Fl54EYX3QwDUDFaahl96tXNlqh
Vgw7sXNN/IKwntGNDoFk3r598pKr3c29Gj1v+QJyRL1sts2qzuhRRxPAX1QifdWT
TM6db1Ih3xQw9L8qp7tGtCCE3Xi80zqNfMbMQfyEHLv+la9dhXoAoLk8wDrCPs8D
Zf4SmvZS5rj3p+xOBee4mITRroqRu62t2yjRm209ujVCLe881DLFS/7SI7maInhz
TfIz19ijlTmqcQZ/cJz0RYsBbsG9swYe4wFRWrHtn4AUZt5aHMYW/MQIXK215Q+N
VFyFnGLQMnNsvf+Glttb6UKrd50nECs0SCm5Ve7y/m8i1oTGMugz0GA/6dxQtMGK
f76CuRjWCvs0DXW5n5uHfzOpCYkbad7smxFj48kZWhcX0NS9Y47j98Gl2sIBQY5S
Hs+n71fxvL43Zead9v+sYgYxcHHHtRLb1Ta4TVQR7yEM7D70chQFfmT5oDsm8zqw
klfOYcrWL3KUnoYJi777ysCD7llfnwHocxu+2HBZiAMCoQvLYfiFyo9f/Gnwjz6g
oSY62059NnUWIz2kXHlJOAEI2C4VlY6FbCkrJ++VYkqXlMSIQKglvPh/Qola294C
hEGvNlit2djgxm3kTKfdgxVFP01EUUSUIXZW4KQHn6s/nr0+1Eo1Sdd7yMrkaSiP
qFyFuw1iWkht6W5iSy1T9wJRLnYVrmjOwUMVx/j9r3rgVgQXqDVkpPfWTT+iA4HX
Pr141zn0EVWATIMFVcmMZUOXgIKzM7k9ldwoKJWt2aKiUwQthMhbBgxEQy3XP2jP
qq5KrxijRYdXzQ0wJK49nNCYqrruBG9lb4mVWyp4MYk/J1dM7uveiu1wmR848oKO
5/25NvhcbGArmxCE/1yv3IHjsd1kcUKulrEzVca6LRRV7vEmLtNWc8lwJ3XEe5t6
YEX4SkTWYOT2eBAWqfbUBvt0WH2puRjEJf5CW03u6UZ2DTk8hRo8gcUFJpx7I3nc
0fH70zCT0Lib/oI6IagXdqPAqgTUrrxO8fwIMtj5CMA99oJs4A/SmMsq2wpPI7bM
x/j07o1JqxUmvcXO21zx//pEHfkMp2y0B63k/afhGiU8AingfU4Uz9EA75gTWoFP
F4hhnKEOktCesn8Y9JeAV9T+Nvbu66d6WUFPWdYZU6qAu9pTxJkUSwhXnHe9lauy
J2ETyIYBfr46CGgJ4jF1T3dP8oW6828RyAx/oddCEDReTQRCo3GSxnagVB+kcmdV
LAJQRNTwqDusux0wIORNGi0jfHSi8EUZKoSm33wi0jKfySfTAGUUtVHnrdcAzFoM
DsW7Y7WI5C2kIHXDxglmGwWk9upn+FV7wkoGjM9FTu0MKo+Vg83yFqfI6Pu7HcoP
KA9d3sv7wmLVDtee3faEt4Wlwq9xWgJKKdSCd6/faMcQXgkvOH/nD1KgvrbfKWbx
5rGapwbQnyth5WAPqGbtqpmEamRfzGkn4IOypbrZbGF3pD8SWp+W90aSdaffgiKB
S0QTqPkedCyhDuGc9AI++vbmr/in5mzyx7+onaUqnvCmf6iW0bpPDspa572jgfJE
hVsIVRLp8ktOY6wh/KBDul90AT9bBclFJHZV0/9wf3KdXFt0k7l6ZenurXVm7u4N
AhbsFKgTwxF19Z3ljoFpEUK41/+Log7e2wM3I9SfAbPsuxOxCfT5ejl4TSUvmfmy
8dL2bqnwGCRlKftUu3MqA1Il825zmZLk9rAf35BfjnwCtL/w9l8jCRwBn8Pf8wp+
pYUSUFkPq8qHqtMg8mPDiMUIXpDFdr+OPoHsSbc4Vp+edTavFmyJetBXcB5mWkwO
B4baB/qT+JNDzuDveCns8c0+rUl+d9NypbnnieuUVIATGMp9g+cKn0gApQLIVXyX
aOCHwCdqNcEQ7UctUwID9PjtlNOW9plc7sCy7xGeufxFk/bn7To/ZrR2rSyoxYi2
fO2bGUUPK9c1qwfRwro0mEjwEbyB96YzUJFu4/w4O8Q1BQghEc9441MCkFfwERf0
9x012nc3g4iSAONaXpt8GiHJKDl6lb8XAQxPXF9p4P0o34fdinab5blnPUTrBRcs
A25aD1zmAkeuLK6rNC8h26rdL4hy44M8xmD31Ij3c2y0d89/6ghAUL7hiiCryRNl
ocu9wF/wS332lQvR7FxIRNYVQeV9XkKiYgFSDC4rCEwYxAhTya9mox7E5M7zgPD/
u+Uqmcuuq7jYUNTqjFx4KcnE2hDSNbaCsz2OOKgohNDctotLWz/0ALBcBAYRMJsT
u/9EA2rxf7lo7eK1dO1lZPHnjOhdU4sxlz8KQ9UtMPl/VWmBgTlnaArWZgmd5Fbt
n7rV7pKwxbwLZd7Fjm9RB7t1Q4DfFDmixJDeM6ykirJLvMxRVccIOIYjTVhidgZL
cZJnor+5HzdS06gFyuxlM4mzMb9ytdS2kstU3feIpf62DatJ4WbXYdR8WtwoY3VD
ora12TSQYFuakLnDBaMkRWi9zjPaW8O8OwITxhh+n+VtgbLii6eDggu+yAQ7I+3A
zKBuIApw5P8eLLev7agIlMBKcdL+PFGhxCMt6F33JOysjHNgVKoJ8kG1kUuiAO9f
5vCdSHBOBVnipel7GM+OmSKna2Z+POHroyVjrTohRfgmZml70P7Av1QpbBvk75+O
RjnaKctbj37NfUXk475YMguGJgMByaH3adECwniJbnCEblYaXFFyIpzd7U2CRmMy
z8Ej3Q3XsTjZrmO+Tu2cggAFuwcNegTS8stUI+sPtySgvxwGS2yiX5VMA0wF4kR0
31/OPG7xJvTS2zOhrt/fo3Xj95AGkPyGdHGNqiqWVpYMufsoue1LeAukXiN54b3c
BtVCP0AG+QA3prqBtaWvg1aND01b/J1aDHadFOZ4K7DZ+atYquLk7L8CV2mwSVbF
33LOTdR6dRT3OeuPV0mECoVwQltRBXlNyFLIpMCDys3okqYoe6PhaYVsKJerk1i9
63kQG9DfVOV5UEtQKg1Afh03oQEei4gWK7kMQ42EsAAcDzrAQ8ttRtxWWr0sS8Uw
U4/oKMJGVys2ZVXYheaPWzR4fEHGK6FaZWPc3WQr7YNuJu2HVSQTCJK69icHRr/q
n9ohZc57MEU2Xx3lEQffY/XrKWBGU/4TCRq6VNdXMjL5tBGTBIiNSmjG+IZLOqoV
Ks8NUGyiCwG1kbNloJ221l6PW64xrHAiwesVEt2Xu5gzURKhPAX2+LJsDuiCRBL3
k7FThpaRA8ZzUzxJShp6bRriWjX6OeY+F4y1lOu/pswVAFRpe9pcfH+Ax9lVz5JC
wrmjicWJSoIK3bANmH6Zvvda+VpQRJopv14Kav++/OHZ3foyFU+1xdf+ZxasHHTp
dzmoTsE9PsymbAzfpPYKqbajm3/r13+BrFL1NvvYKRY4t2cHyDZgT44wYAuLm5Qj
Qo9GoBTDpucMclsl5Xz4IS0mDYi2Pkp136UTrUhIugcCblMM+LGeNfJXb6SL1Zj/
sUnP2+8Kaeo7xK5eC2huWADKiW4SA/ivx15qjgza8S2lPdVmTPR0UwaOIuzdPk7H
RFo1i7hn7VAfWBKDsio6e1isnJeUHwfdhaDTKPCMLqhrmdI2+jP7zX0cHu3CpjS+
mtCmxRWi2yNofGxnfyYd/0QTIu9o0psd2OaSU0/VsmEKCBhiWzKkNILQIaeApdH0
D0Vo2Mn77VfAE5b4T4SBYBDOFH+kQXcSCzzOKqZV96rw9FVe6MBQynIpDDtdNDRj
hdSrmWQRDD/zbF7EBzN6prYua5KDERy4kOKZGM1URkFb5f6lc4Ixytq4dEPEhj0F
LZt/vmOCx4rvMJIT10vf8lpCAeRyl70MOoFrSvaT9qAHcV8r6b7bVYJTxWKwfbc9
Uy2mEcn40tcQwqKs/wZ9TkzO1Lx0LQw4vNqyv9Wxrca6zLJvHCBxBITUSnzCa1o8
BA3YTHeON/4WT69OCzUe4XW3fNjzttea27Ng3E8BqU90TxgnZTgIAbHYFNhoM6Pj
iDZUT7Wzyo8z0jD3UDLFZ2zHJ9/1ajs1cE8Ksv8lyM9kV4grbaKPFVskNNIPaYcW
HJtPYfOLzN/XKRGlpiQ5uQ+s0APn+Npb+7dqSYIssyMZ4TJ64YywxrulVlvdOSTY
phNRkONuV5GfQqiSL44+BLkfP7ImsgO+EdCJMpw+Z59oWwzTfrQlsuHn+U9krx+s
c0bKW7ZgKCFWHGB5Si5fDXU5NubjJrsmSEncebgi9bM=
`protect END_PROTECTED
