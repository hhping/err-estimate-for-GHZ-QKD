`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gXIeJ/dKUZp1hYrfHuOpYp676gG0SGRH2S+elyLI8VoH3bx6fdTNFr/2iWVQq6cb
hPA8usad3te1WYGemvHj5LD0R3bjzLRurMe715AFw6c5mTdTK4VHKShxLgiXJiqz
oeMyuujUN1+FblqkuaeY/9mDSzw2c7ipAncdNf8iTyYOv9AvkGxtmIZaywsVLkAL
r+EZWjToJKt3et2M75RB/anmZeYSm9IhTzXgHy6zNzZ8V/nWRO7cIUK02Lst3euE
bzblRlUA8Mvgbn6QavF9+YrIJT2qNFctFQGiGSijMFc8pcLHpO+wppimUyTDUtiV
AJ/JtbDYu7yV0fik5UAbdqKN+NSgbBZ3JRyoEk8oB01hnkmflj5qV+vEQB8gbgV0
3pAUn/3Z6jsB6RoTf1mEEp9ZZaLeQyiA2l3nwM0oVbnZoFeOrzIRu6L/b5mT1492
Cybj+GmiVPkqK5QfNvU70fIsxifM3AuysH2ocIxq5d6RaegdfnLd6T9mhIdxxIIB
XFw0ZimZrns2ZxbVqiWUy8GvswZhAYZpKZ2Eyqd/FFiAJoFEbqOh0Ol7+Rd0mXLK
pfnCDZ23rWhlnfyGRyhe0YlP8F4aUU5s/CZq8ak6Ia1cOrE0yX+SHiNvCeLgtDmD
6DNWt7XjdrQnMC3Ii9+uhONFYFMbGdYL8JtdMybOv/jZdiU8kwCQiPqiJH+Brb8p
HC9a8wOLYWdp2JgjGQgJOsdstmn81+gvv1kmIyijP07Cuowo05v9kBpqMRAqfsin
eAxkRW3f4ut7WwRx8iA+d+kilUqPpYbo7rW9CQy5TXl4gC65HuvXgNPKDAXyJL0a
3bTYyr+pdNyv5gST0Cna0//BOJyKnnt9KrwIEd4tC0QnrimIz8408y0klYN2+x/C
yjsBle+7VOmVFfkf/qr1Co3nkLxfX3871G4dkgp0GsWRQQjmGkvSrtNpSkLJJqSl
42r6tINT3fQLD48PDEnaRx6mMNQ+/wT9CS+3bLHwHvw=
`protect END_PROTECTED
