`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m4XWGYVLaUns4lG9IyY6gjbSbL7AyiSPy/486vihxUzbSuP2d5YrGs21HkDVeE9N
hKzSW+1JWh7CHOJ7xMstHsz5iiIJPMeU2/2PPm3ZK9tiEcUNx7g1y0+dKR5eW7PD
2o54MRHVHDlH7ZhM/cdqBzx1NyxIx8ZXptVSq4l78EY/7E2+TqYEyMArk60JSXKQ
c0d8GZVsH9J12itNz+G0ztcgE93jCSXY9o0nWZe0v5b64WJ9jhAAqSe+tFEivqlA
YRuLJtp30dfkirh5+gidMe/oE7jixd8zyXrlGCiOp9GSk4Y2j+3tB+uLx04IpWUk
v5pzX+a5yfFkiVSESajjnhnXsYomiNlO2g0bL0CpaPOloKcbpeYRfsBSHRymOjEO
pS5wGYbJ50Xbt3/Wk9WcBW9Ys3/oCZAlL/oDMWeY1vo4s+2E4+l3D4Vyzb88zpbu
8UJW0at/LsK+fPX0Nxw5CLw43KvJoWGwBQ0gETsVAK97EvNp8dpfqHB1P7+v7Lv9
+jfJzslL5GKUCOLE0CzICIWvZ1GWCtyjpAERsv2a/nUjygBL+M90zCsQFcJSyxMo
`protect END_PROTECTED
