`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qppie/ckjVnk9Jk6wai97xhUiAUKIXZk9zIRexRukonBJgixRcSpL5wqp3SyJ1gI
eKprLTbkFO9jcYByG7eZf5Pdb6qJdAOWzi5fEoY6fsP0sKu1IQeMMIpuqEnx0tQq
IqhioaLiT8FImHlxtd7CS2GHKGOqUKazdUrE2IWXUTJGXQ3rmuCLCK2aNQp/mOSr
RUOXbP8bEc/SW7Xo+hBnSw0QJ2dsMa5rtaGBibRVhdNs/FofNdZ2PEYTTV+XP5AE
Aunv6GBTzrH/RWLlAemwydPVwsu/Nkp38VwUDw/ySpA3n+gHmelR2g6X8GbazbIL
+JsBmetV1XINPHxqBQKACDm7wZNirU7H0a+BWEk33DLHg9uaetOy3rRmfHfFg+UT
6RvREhPosRWoUDiunFDSrBS78S2YNJp9xcY8J2FfllXqorXNkGJ9Zh6c2Fliihu0
MErN6/VfjvgS0k3Wuymnpg==
`protect END_PROTECTED
