`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O7diftwrwnEfBKU3PCIiH7/FNyoryD5XRO/PYvo1ddFCCWcv9AHuvUNyOSg1yJjq
3ilhAdNlZaXvb8+DTnU8l9jamoGMOga6VuiPTT6y6S4NBqAyO0hQcku1RyWRihZl
6ZNxZ1pTHu9tLp8rR44uINOcsBorNdUZFrTjSOtMgJq8khbcC3vCmlCndxFEpLTv
iLSV1UXHHL5DghpuwW8uaekHfNnDE0RPmfe1tBxiNICZC6JitbfW/AHExjKw8rle
fnQui47xKFK+thgPAQhbOtgdJUPJ2N/7eBdYRblt7kle16BWjFaW/TaodYX4pEpP
cK7CaUIjVZmgyyYjw9WMm17ZQ+Igq/H5IIvvnNibVJ2Sbm/+nV7jdhCK/InOPnd8
lnvrrE7aFpk6hXuj32tm6lkBFgtG0bCWA7+egD8Fkenesc9Hhw+UM1mQmmpSiy/o
dfBC3+gd5ffMpal6yw3oN4U7zB2CY/5YZs76w+ykTe4ePNLYSRvqmPLkgiK2YDPt
UZ5ZQ74D4gwBUc0XVSKRwO2cwgyOm50O3IxkqbE/f9zbvOTaI+x+EFycUZI663uF
3aiXFXd7bxTGSfcivr0OYOMytF8zZSKTFyI99g8XjeubEg7CmGdxQZ8oZSaflbJw
O71u26WZay+OIAbQJNuEiLvbpvBRrjzywW9UUj9GTXW6mu7+L8wE0DJvYg2IdII6
cdO4eEs5cqP00vhiQfB2jD5qZJMCcKoiY9GbigPNdqI5QqQaj65u5+qf0fdC7JHD
E6uB3eik+95rXdEsWC0JbgeRmTFhkFH4KtH7ramXven6mFeaTIgseJnTQ6TUTewU
OqpVv47Kbh++qze8d1tiY+vpZBUp6bQw2agjcXr8qBZZgizcllPu769mr+Y0qI4P
etijYog5nrbpqyW7y6KUYGFJ+Lj2yiw5xVCshZp53hUbujY0t3VqPlHGcG6a1L5p
23MMybbBZBXbSNvrRC3G9AK7Zb5WwpJnn6Zzx2nJ7Q96fW4pytwbTMUGk1HH6BVg
64+A/0zCQ3YOCF9CXHhJlbOAtuucyqg2b+dvtyjW8jeqh+qX14ixFPz4oBMei7Cf
nUf3UPeqB+esiCMmpt6C1tG89eIz/nR9bp1MEixJOGYZh/Koo0SQDw1P7VO9mmCR
1KUe74gAlXhuqvoNeKPfQIwemR+iA1486YBk2Gx+UN6hvWDVAkXHowTXC8Q1/zuW
twugylQNsI2xvY2Jq6gV83qbulrslNzpAZn8yT62DUNrxcM42ZJ6cgmeSHt0p90X
LGynMB1N/Jasoc9l/rS9LA==
`protect END_PROTECTED
