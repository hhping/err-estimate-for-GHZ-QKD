`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I+qfHY/3GqOQBZ7uOJOjBDNFO7vK/BKjPM+DslQ5C/y0SeB4RFIV0YnzTKA8ULlm
89RvvEqSnD+P9W4S9YVyHHUwmzrBTdJ+wuLDEgbAmOdQ+aPD1x0bGGkpvcs9XSnm
+geVMqlig2RN+ERKwLtEw/WU0rVVDrDWP5i3qipNxoc3seCK39+9vwxg+6OHb5t6
6XyMkRoaOxTIJRX5MeoOmTbymA2vRqpTwKZig6m/MnS/rGNf/JEMeq/O1dzTzHE6
z0YVXCpb4M7xh95UF3UTszvtYaTDh0XpTEZQTCWqIoxzOejBkSwhrFl7EHYDS2NN
Jca9fdpkw7KBnb7XFGTWftpxYCqxrxRqaztEKZfnt3JjdO6OAR5+NwVkgNp0dKd5
PmbCkXl0Vi9PrCO4n31HFGhtIyLM0UooRx6CUm7LAhJ03axvDd61Y8ZnT9FBaOtA
66rNZePMK+b6mvy/fUOjntF7J8YvYhDmPxY2hq3FFYobTb/lT/PaXjrFN/18wIB7
xog0sB9KX0SfqeyiTNdRqMZ+0eDsyjWW7L4PwgNwqXnqYI/AoW848PJFCHOMrgXY
rcoOT69E62zID0ZfgIfH5OqehihPnKR5WzF1X/m/16wivP3kI05LilxVZ6iOiwnW
y9xfJEFSKvGQO/bSxoJGDQ6PljrybNvHdpSc8c9ICtmvV+1dy8U1iUqmL0DqHYJI
va4LixvYx3kvBkDYNHeBtZ7uK213cjKjP8RDCL/Od4O028hOwHCppuultKNhGBrT
ppykFDYKoaAgg7QkkgZeXKPELNDnfN6Q2cIz3iPPXwdIxREZd7LPb3LkKMWg3XiK
zgB6CGTAgLqn0HzOuFh9a3SInuaaeXPVXqiaDfTdu6HIRh5DVXgJn7WC02FxE3ee
GBXnMvVVFCgV7m9xVCdiGjQhlhfka73EVfKZTo4/xn4jZ0uI/AAsCaQx3E+HIgLI
xGX2Jr2QyeXR34LSXq4bOnp63/kVcs6cZydWpoFZlSc50EVwrehsHVbV9W1LyJoI
Wzm6HSQ0MjJd3Zv1Oq25SG/HADkIF8fqnQ2QTIKNOwd4ORMUcU6VJLUsuHjGldOr
birlZEOle9XskaAGPBbfZvB+IyFFeGdovVH1zzHCWDSy9Fus/unVhBveUatudBW1
pa8X2p7wCVqkjLw0dvlaUXjmjMvRK2WR/68redeuUCV9VIXbxdsuhdJxG0dxLVk2
rkT8mqydQMJVu/YW05tVqkbCon5a8N3cDvjTXuuP2SEp2ji18Rxcx8VBrnspv02B
ba2Lr4wDhZbd++d4ArtGQ/qv+1xOg0PXtveLyFCAV1Et7n79iiYlkVcsaNZwRCpn
yZiXC1wsOxfsu9LI5oVGcKTdRL/EEqN+uR7/f2hl39Ucpmgs+/8yywdF2OzUGC8K
S5X7crZGZftfHX0qbmOM928BC1qINW9rL2tSqDSRYYfb5YUhv5qPEZQrrbOyAMiw
Ge5At7VJwRS67c+KjOi/imWYrMedJSomHE+FofT/PytdyHAUaGeWYXLvB83Qv1Zl
8AvyBPEjfiyET10H6Gyk6QTIwq567WvXwmLiCNRzjWdKM4MCSymkFgXc++iR0Tv7
oL/lU173YYYbGe9wqIiaXTFan2H7aXCciyYQ+GZG3RX4aT10TJdOt5pVyaU6pvHz
xwFCftjBNaNGmQanX47QXGVldoZ8VKjj0z2btRJjcH8s/OUM0/lvQYnCV/gVZTLR
rsujbwLnPH3trhA3Umyj5FQTYn/gENJuRhqZ8G3taO+IMOad8EcFRRM8KZyVSqcC
poSS4wQncIfAEHasQdeARlAD+jCfBTGbY0DFhzCjpwnGQnQuGXOvwDOkGRf4UhN6
mckiT5JF9Ri5KVqE1+3fCiRPXAm5GnO7Zugc59Xaq0s7T8/l8xHGIqArW8g0HUhq
owyfA9upH3MXTepP45KSkf7RB3t79w1rBYxmAb3QEG77JROp4LB9NBTODM6uXUkU
EcDZQU/y1y3PthdDbLKJgk42vrUKqAHZxeaMU+o/V57C2GknxjKKHU1QBaESDjqF
gKvRHA0GIaVLNnuL47KdYm1r3iGUdylBEUzyZIB5mI/tFHPKcfXrywi/Ua3rgPwq
UT9QHjZDwe4qhNpT1YVO5Wz1uZBq2+JQ9ay+6+Z3UXwujYxux61JHDfkaMWLwLye
CCLo7CazKbIp5wQY1s/UqdsY1L1Pu3m3BxNNZaIzmELVD9JD0v2omM1kBdKN7+fR
Mhxf68bDgaObeXIjdl6QNyYVjea9nuPE4lO3JVqwSRDtesUEPMeQSc/asnL+wIbT
yF0Isxau5EsUbfzHAaKh/xtsRegvjkRjjMtNINI/tGd9X513lK9qU7UmMB2H978T
Y7dkodp8rUuA1EaoxkB0adkJrnjPS4xl9X+u8Luy08pZxwSy9uLi37NFYzr2EgOf
S0ea2xwjPPdsE9AVW9FySQUIURNdfeoF68wZ1qWDFHSabijZkvYv2oqHrjlEVcQA
N0Jwj1b+OFVLzb3kNQ9swQ==
`protect END_PROTECTED
