`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hONMWTivXw96BI3iugNLjOE/LFt7oLLniuWgYPDUCGYtyV8c2dL9QmuLD17d+ajT
S+CFz0A/cg3d7UryT38PV8cYThVDJ0gEUzBr2quERGYJ9MQ6BSnEpArgQmmqO3K6
rB221+ZW/gmsKs3xWbkON6v9cyhg+bpq3cF7yO6nsvWCymeXGV3llj0u5Oy3fPU0
1V/JESlMe8enYKpk9BwJ4YkRD9ACXUBw6Q2t+XR022bAvDRfASg7mObrXqCiUm09
utEdVU+Fdx81banE4uJd8bOYn/r5w2hFb31YRU0c3AkD9imo+ufZ673nEgTDjlB3
+iDAvZ1xQ/kT5LMZcZR2BXIQyvCOjPqeuU97vgEN1z38q3YNoa/8paTadAnBU1ty
`protect END_PROTECTED
