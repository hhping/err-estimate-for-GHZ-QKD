`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KBhSR5ZJFzbke0d/KQtcRq/aA8OfkNVuYQ8bQD3TtuSGw2eLeXxCkyKliatQ78H4
wulkw9wn2sYDKP4+8l/MORt/eyvDySu+NpCqSLVBn3ZBG+Rw51kSnJONk5WCLZAl
9XXyjVggnB1xamnfpxLuTqU4hSqVufSchqezH0/Lbfq/sSl8YeSKwE402ccOvSXm
TfqZo1q178nxesIh8Oj6aGidY03R6MOHzDpgfYfKTHGMJYDN3wKUKe+rBSbWL4Xr
oUGDU2QaXcYd/vqwuBZpkm8eCsVUZETgY9W3SE/M7mytCuzZd3jDK9xIDq0ZUaG2
GbkkKTtGjaKzS5OwE72WCjCoAo0CGl/45eUVnKpHM5eXS4gtIDYEVimjLlwcTuMd
staoWpHzrsjaIQUmG9wHjmyO6uFwuBjVXXnMCCGz+e3lgrV0Hw+UpFro9s1yMAHk
q2ezs4Qw80VPgBE+HZOTgwQg8Jc3D/O5s5vFy2dSBNiTj8Ksxw5tNH/Sl3mD9OSP
sDlw05WCsoawRMhzLfsSmcEWw2KHHSIFQ6Vk1AmVaqjE/Z90pvvVTzIqbABSaY68
WfECLEyyEihB27mTMMj65OaJLkn4KK3uV7a3xGg6/YOH+vAxT/Qp2AGjnsWELq9o
j70JcDRmcvVPX9xZ+RFe5nBjE+0jl1It8b5Rr1qzmcUYD6Zwqw4BmiiHGF4pQhai
w7w3cKOnkxbR7bmJVNyKLXY7KHP4oVnFX4HznXST44zgiNzyf3foY8RyeMUJBQoq
fOF7F9pYQEIS4gWt/3mRgvvPG1N2NDh5p5lKsbbSe3nD7c4QMHHwOdfKJIfg78RJ
Wo/H60iCQZ2OoiKBZPamjaOtb64HbQy4QFi+aOvi02+Bbf1f9EPwRiqnEWLSdd9C
0Nt72RnGYdbQqB5cPrRvlWS/T39ajAbwl2jBxP4zoPzSRjzSlmHaREK7fvOsErjk
1fNaod4QLBZGdBYhcMaJ+yyRtRPmrENKNHswv0Wky5dAwreoUUCdAb55WO02oboe
khhyKMm/BAVe3wqU//y1bTbUoa5/d29eBvSjubdNYQZYvCcJob5WBPVYbtpn5FfJ
woowbKX3Pmt+BaD5uCJkKmitl0G6RkQWZWMr04/GHJew9DRv0cqMwy8W57KhLfbs
yLWccTwM5XlEbEkApm3AsxD9IKovhBAgkK20w/OZAuw=
`protect END_PROTECTED
