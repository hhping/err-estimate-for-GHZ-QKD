`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MPl0NDBizIaE0nuMqilx7gqiTly2XRA4VU/QMHU46+ZXOX154t0RpSw/HdUwgWam
ENBiOw6XKeotpgLTYATWwvwDeMRgzWxurDCDMkOEf+R2ndKzahH+4w3Vv8TjjTlP
ySpH5sDtWk7cBRR5pKLR3wrrpuFTgdZtsKYXlpEdtaeUrTzgaKnni1tfBLFw2qED
uCR+UkOkZjYU89uoJ59tQSbZ9NrphL8M6USMVvrIUOwS3awy3cwx73NohzEHxNWp
Yvcyk3BcyeVx3t3Vq3b9PhGMYXZrDT8pZGYZ3Jmwelbg8fk8kUtru1jwPlhDzvcH
1lXeKauNGktpCqVVWQfkeiuyqfg+a6fgnNwnpW3jqopvKTXmTsJz+Ne7pkBMQrdv
MFV1ly12yxY//u1dgPqos5D6Cv6rkjQ5V193WvEoDURgMLKdmuY/0WTcZ6l+L9ws
m5KngO7u/5QYM4isEqeWKOVGSCFx5fy+MhQ6I0C8V8aiDzvsOoltzmabL1EqAF6P
nGMehRPodhDmNO+Xdp5tl81bkF8Z99QSUOFJhhQxdTwDi+u8tppQ69L7SB6UPPOy
A4jWMHQUOe+wbSx6Tp3xkTO5Fa0FC2baikVfGDrHrv1rcSOUMoWTLPQ7zM4JwhXH
Ja6q4sDeQdZPy5NzsTMqLz4EaflH3459InMlHjdNg8ozsg9WX5z3QJ+krHDOnzhW
csl4FH+NJHc/5+K4vZhFQv9QwzjD12URwEPaqX4bXonTCpSAoMeb+5/NyXepFUie
jSjvkt1wBbjHMVGidad/L0Nhr5iBbVHXzfVc/tnvfOcJHKZdXEzBxNuu3RuG6c17
A1hqb/CsMZjhTtMicse8zv/DeOen8hAvoBCJ0ZcdYkLmPObUgWlwIWbWxGfdX8Ia
tHA/CYTUb57YOwCwxnSX8rTrf4hNlKpQ8fqZNGR+IUWeEBn7zuLR1EeJkdePa/DH
Xrqjt6XsqHU1L2jUWVemfNXGhFYbx6sTWnV6sVroaYfqIofHx9cE1XQ4NdCkv5J1
0JAyxBZOkW9ChZKd7zUyI1dlFw2p0W2Hztx22Zil1AokZQMbL/OCbPhjpkkRh+KL
RBl+7iBUlXQfkM7LGdnk/nM/UGrc3ElVrVuxZyFYqeb/nKnZVWRY1IZWqfw6NH/1
WFsRQin/cHavz+4kPWNCuPbYXvy8IqitFwr5AWtB2hrGN6HJo53vVlRs3XZrgHPc
OrkPL4WxYiuztBRmpkw/1IvBVEs8A0b0Aoz+sVNAK+jy2eeGvsHabU/hlkoLSoLh
vBzPs5WdcfmNBRIgVzDnyhrAyImEFApdRCXWp3P9li0l9MymEKCeNwO6F+cqqRyC
uY3QVH3soblOhAQuNFfbq5+HxDzBeZOB4MmpiC5KCw0oWq3Xau29fgzuLjAClHrS
qQg4ZYatBMid7+AihOW3E0yewZVTmZbLxeT8I2Jcwgd//C+gfMN6UtBu0FCjR4Hq
Sv8w22K7iO5AFcby43MIvNEtiSvyFMFP7wI/y2SGpq/V2Pu9uUp9hIIdhESNPVz8
p+56ByBaoBU3UMjIqO/pGNhF3lZgInNbHlrtBZYklQMDkI3gTvyVrePimwFmEp2Y
aq3rXSt5kRblVRhireGKXogIUR3fWtY/ekXnIOCtpxwW1CtLyz/UXXJGQR1s+iEX
KdGPv26IQfgyW/jl9rdMZjeMtYlj7qI77mp6FMMFBqbtLThX0YFoputduCWA4+WZ
vSV6imtf2jSPc/20JFm0M0YX1KtPapi/uwvXtUjAFubdqYS1FNPTHCyIEbbeplkr
46UTqSl+v4AtK3coH4EPY/eeA3CvTahwDGYLJeCluRuDMEH0hvdBeNMYnjKQRyuG
rvIB1NT2NytXnkKG9zAVVlVSkecb5bf5nNkNtzO17T3jmQAsXM2/d2FRsOvX/QVS
FATzDhG1r6fNHKW+58xchgJeswVyvoM1Hej9xDFPs7Zp7LsvpQZQzsgWtm8dBsFM
vlywPXIWBB/lVpkT4NTJOuWN8vrNGl1JYA4RlxmqGYLd4t+IPyRxdvN13VnSb0JT
13ZUUn3cy5y9INMXa9Hqx7nr7kRPC5jmF3WRF67T85G9z4azZyJNOc09J4D6wu24
xMQt7f+dRfG94zmKs/oISyBNgDT6w61/a1PTJUYuGtr33pi7sJHNknUErztyfGD+
HTpsBxJJX5xD6QYeqgKc8+leK5DMofjktgzWCLp+XRXM2L5P4uMatcFiXXf5k06D
80TjPAjUghYuHRhUKwxmERk4+edHRl1E3seIC/fhFZDoeFAhn/UNzjkBb9O6tLM0
qPzwkrUUtcRhbzILaA6u1oDKwhJeC7mrRw7VHrN9iIqjySj1Xp47GdRwltDsOIfA
Llv39UnFTaKWQ5BtKXqbAziR8cEaQ+iY0NVU59DkCuUoIC7dwK2g5wCr2WXL471N
Ee/IjTQwwhNZ4vG10FlxTdvQktJyITVmXBLQoVDl8E5csubhhOO114BwCoM5h7MP
hl8tgUd5Q4DK0mjB/AU4ZEzFXLLb2Ng46OfudtLDnXDITQBO+liEPaIN+ehnZBH6
zUgiY7kLE326kRQwd95jhg0ufnsLlJo3jS+TH3NMZtBGKsQ3vrmF4OWL0zHFXqsR
6Dy8FofIltGqch44YIUOg8ZvCJffBKEgzmDhmI/GEQRTOiiAZrJuDPI0ilYmDeJB
wjjjt0Xi/8sQNqTv1DfHhts42teDpMfjaniXhOlQXJwskAUvainK2RfYSXhX7E8U
QGhZQHORX+mZOMOUAIpb693JjTnjDnGcMgWQ3puBTllBH55f79gOfoecrq07DsVP
DsSjPM6EgZ/G7ZlkXwVNdEyn6ZvgB72+LvrITA9ePQH/FXLKZEHpRSJQL+1612FE
2OaKAznYJlWVgVN33Mu0FP0VZosDZwxVR8gngRAC6g3T3Gf8Sn+dKxAxOqBV/I99
7ua5+LUS7y9m0koWiuza4yeCTOHy9GFdaI5AGDzdeFco8LU79VBlG2RNFB0jBW2p
yQDteAjj/ICWFvEuLQ5QShEpEmo6g1WP5PJ4hi8vS8JVGDEPnsqIh6wTYfN6uHIt
Jg7IW7T/f+Jpk8MXsZeE775vu2zgoqxaR0TxtnjCz/qIkgc0Vvw430lH/ldKwiEC
zZotTnDEfv3f+xtz3HCz8XZGQucTrOPu5fAusF2tc7vItJnQMdPqrBjsmIPr4YwX
WcHW9YyrDMCmLE/6Z2nhhlbip+VapUn3uMfl+oozhLRicK8ZJcvKFX54EdplUEu9
ToyNsVMXP4h8108TUv2ktXd3mGEQ8ulpuBzPH0910pv5fBv4hKAEF+7S7AecHRWQ
iiQ4GDPfvGWzKUENn6QaI84mjqKdn80ySiDuzgpGA4M+SLBe4mSCp4XeqsM2F3d3
yPllOLGUSQF3gjc68lkxTQ==
`protect END_PROTECTED
