`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZJDalPT1scYWrHcaWfkgVnqtE6GTCFwQkQSqHiesUwuzopOlQuAmha5wyHAghJYE
1Zn6yQCcAp2rRPGAOtjzKyLSXf/pYqCbFzkmz/1Z+ADf0jwfO1kAntCtOk58QsRm
NoEOR/Sed/ePDvk7kmb/gccPFoDjWuisNtsYRFNfekdmrD4BHJVBIRSQKpre4nok
ClyzutvihUeL+tj+7WaujCTJn675s3GJaHSHN1orFIBgZ3kxCu0ibNNJTh2LEYuo
P26iXNke/W6WB0ItD4IHbfjMv2lE2If9vsOZ5PAriql9zXGRc3pyhQYqLR0nkxuE
ruLA+3njAwfzhAQUMSIYSvTrK82PEYUV7j34M45YHrhnM46GrnbEpuGvqBmNk6t2
6rQZq7LrawpbRA2fIahWOhKPM+lg8P0xfAv+OHALOZeRkKSsaGh8ASCpn1ZcPNBZ
nw1pmPI9cVxiXGrPC426RS6+LfIA2AXKtPLw3gCJDW8ygHZiOtBlFDcMpJ/BtPhD
1r4oJN6cDNn1mu7IUf39Y4wFSGeYqA6kpPprFohqIpt8b2w+5YqUkVdyjKgt7smZ
s52eltG3U850z11H2OhsN/7GsOijsYn/G2FxR+1AkO1psgmmKipzF7rI8c+zAz3E
WGLWhB2XvFq3j5AIA2rPs+sLl+iUCZpwvSmAJSx8cPJMd81bBYutPQfbXI3YyBht
LZDI2tkF0HUQgfnEaWqgwi00df6jSNUIuo+ImfFiY/L5sqHDmBgrbOh0t8IJqblh
5i3kRszNDwWx0vMhQNsxUdzltHx6coNsIesKfSjjcdH9LJl1WDW9z+Ih9dNAJq3v
IgQrdYgaoZFhg5f/vwltH1u6bwTC6mUd+7FHcd8RugEklN5DKi25EKXSWiXNZ8tw
SuZZsppx6dC370uc584fX8dcJq6O96idaw9t5iLSUqgMMqu1EZ5ER+9mzWJsRhB8
8Rmmo638O1GLnfNhbvNONlvPf3TVmB6LL4Fr7lzz+4VDMVAlIdiSN+2wHiuJV3j+
DNxdUgPHQcNRf0SkxnsRDyw0suAcAj+trmjT5W/3j5pFk+45IEUdkfG0ObnP6yUT
FidXzSUIlFXW13aaogfqsClTcm3nGV2y2nC+AH3Lke/kdBVnlBHMW7r96Y+SurLQ
CbAt3ee2G4d20aen4RvGAaN67AKg2K8meA4SX5EK5OjML2KF/t0+ecwvh1Lwf1uH
upcovhVgxLEr63DUgXuyJInD1j2nbDfK1XLbHRm5HxZMWQ2jfY4x55hNhLr2Lwxh
`protect END_PROTECTED
