`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oCd+SezPEGPRdL32Csby44Rzijhr+qRR9ZgNikyUCy+GfMWuVgmdmR9j0f/CUJci
t/E44N7GX4dTjJk5syOOJjoty/ondPSLxGaTWL152ll2MA2tUSZ0PmoydI6ey5Zj
kTZKtsMajJGAnJN6F9g65IWsbqdEMHW7yWCvzwrDdJw3uCwGN1tZF9l3teJa8hSj
TMQOFVVl/ie3mh5hIKfDYW13QmRacmLjzdXist6xEm9lezRHVk+C7N+ga3WugocS
KcQ5GQ0xDbsJDkeXVRv+X+L25Q0jGlhAxqFOokrh2iGY7B0WrsLIjDYGop4/iIAa
AqfL/r0xLJc0/1uW7DvadWBZBh+hvO41E+eK9BtiJbS77UvD14Bw9ae1rfz2rfqS
5cY8m2y5AYsfNHyzCXLzm1aEmlVuz8C4ULqIqszLaBpPSMDBn1fmbraskwVqkGPj
8slMH6mOI6WB+aMcAgDAnA5ijiUmx8XScsQ7geZZb2dGHz+a/PuJyBQWTyC9Zqpu
Cqh9DaNkwTybmsddG7eoDMeFUpBaC3Qdnl1FR8arbl/Ace6TPUzujEPvz1bMC3y8
8p7BgrBpGwM9+qUs0T34Ql179wyz+4jNSibfLC163oVWj88k68zC3Qf5218+HQun
mcnvMmX1UpuItdwfdvLQ7vtdo28USDe5Fpw4MoQxsMSMbuS8S8/TXJKChFVovFYL
FKukpwG3phz7S6tt7sUOZLXBFzFGVzYX1gWqsmAgRi2dN2alnZIOaGRn8Ubm0apd
F6dnfx4Fo/FHi1dBbT+sT2xRUGFDJobJiH1dnQlT/3h+AzXP058xIyWnVj7g7RKF
iiwdoHj/KeGkjrPpUPFa0+Moig1j1/tiWNGiLuoA0ECZYmon+PhhLfRfSSD6RP5b
0jMpBKzvONRT9ElMiDbn68Y7MhpYweFEFEoF/EG34IsIeAGMX41VsLfhKRGaNrPj
4Cm/ROpqQFTx44gyZn2V8vuJSdrji2inQcVMFIuigkHF5fceaMPjMrNjGPE9NV4c
9oS6OEgxwUzPrtKaca9pFVPnUnInG8pNSTV3jlxiH6pKRkYat+46/ZTcs/xP0VOV
/mJI3N+6p/5niD/UnWUZZLhL9sOR0dxI7Os8qbOynT6wG+OikgyuNRGREoH8K5SD
q1yJtmcyn9qLVLDsJtSCucDm2IFhUlsmScISaAQ5sCZHS3rWVkCT7EtcZ/xXoRcJ
Nswb3/Kvw+cencf2mKmtB5qsYMWuoQ9b2ELcKqvdWBR4QBJZMLyJs397DUWdI6AE
WfoG7htjg0Ys8aJfOTnfrJaARChLcU7wBN3bz7/CSOpwxt0Q4pVvLf+SfPA4jPoL
3YL2W/lkMXPsqe/E9CSfJb/7OekhTPkG3BZ01DdYoPp9OzI/eEN4R3Q3m4KV4pvr
65gCAM1yAX9Gx8P/MQc6aucEpjykhazNQzKe7rFPVY0VXNVK1hx7OvCmtGhFh8Or
GZjl01nVBzjve/FIC7Jw1Y0U/Fn6GoEN54RJl4s2B3KWRuCFt/RLDKa9wspmj5gF
a1c+QagMWW+xl9yv337J9VkhYzIkSGT0r3Yc8197vjOK9bOzH2n9Nj7qnvPGJtdD
8+EB1mcygMkZXwMXhwnPa1cjCp5diPV4tro1OPXgim5pH+IAY8IG8898/pywYlBp
bvALgvY6MubhTAJ3AVBiGS9s1CH/62WsLLI+domBBZTdRuAcTp6eY2gN1xSMN7A2
CznYE9fACtNnsspkjI+JAbvvv5upmVYSGvMYKMLT1kOq3tXBR+ynfevWSCkbmegQ
9cfYLceRQdg5pJ2AI7/YaK0SXUPSpMqs46u/Lyzb+vdpmeUsaNEOSp8PpfbI5TGS
5Q/l/CdjGjd+kcOSm9fXMHv2K+3JXo1jw2H5YXurQo5aUJoeu5sQ4KiPkt5ZTdA9
M84toHkQxA09gKmUrdUpTeCTpk0TZiHzGHIs7LOmSutWzi/WwGJHYsKblRQVmao4
HdfmeSjH9fbOLO3remrrffgWvLUdnC9a/bnrA8DY1xcJzNRM0BrU8XWcK6rv1mYw
MuJ9z5EeorIgdJ6iLjFl2PA+AnneLQRdWQY6OW+IvXvQ7SuvQB6t5RpCzzDhyH7r
40cF5Y0XkdhVR+pj+9TLpkgH5penaneD5L4ZdBUROYd1nS+tatbBOzq0HncOhp6s
QeJDRJrkSMvTQIIhwU+o8uyWaFWt92eLzIeJDphyZSxmSlm5jkIMTP4OURyJjSzL
N/QarorToI4Gh7ZRN8VJwN/LzknInCc3+grlPBFGYX4JfT9hUxZbbO6WOK/qb6UO
jev6pbCzNcxQlG8ZyMtPaDW47yIBX/v3xSdoEWgza3bZ0hM4cLy+dvGoJ9+w32sU
pz0QcjQOLLE9n47ofiLRlDw5up3VfjwojuMVh6FU9S1ImS4mIM/nwvttQlS7SYKq
SgfXMr3HVXyGYLTv1OYlOZKSfg7QHi7DQaphNUAvxnzEzvr8R6b9QQkx41balogj
ZH3AVGvb5mBZeWdUjSdykpOehkdqQd4rsv+u9eu0Mh0pW6fTdzBBa/CFjkaQOje1
I9+W4QLiH2glW62ccYT1RicblN9C76IvMEJwfvFlteoW9lJI2722NTI5KxLDQgjU
RtxNBourlmxtRVMJH4JvBA1bpbMnut0ZsE142DBocALVwqAzW4MWhlISjqwGm76n
JDE4nDAjX508tq4Ri+kEg3OK/1OOtOqtbts3qhfUtCqotIYbDUs+8Wm1QPgQTxRP
`protect END_PROTECTED
