`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lYy8KguGRuuNhjIoeR8fWzU1CmfLK+GQoRMfd3RLtuy+lMvcSquy/hKrAFTD1LwP
wgGFt3nmK0C0fuiCxBL/UwUn2QXCFYTY3Z1RSeORIU9zt34A3aI7h9yR1zSp1t12
fvslwI2H5HjuSxICGxXLv/tEzDNM2u/SFYSiGMaQJ3fN4l2OMhU2raiDPJQSJads
qr3dXD1JOx5bEIVCco3doR8jTQXunb23bWUwyxNjkB6BFVJcsc8IrN9wTJCgImfb
Ld/Ny6ordbGmxO6vsQo13d2hHCxfQUPgwMJcibD/5XHLbM/dbfD/Eg3hJS8LXgBR
v41G70QGx27mWxY5fcuMbu0UI8Z4T/wWVPp+x7d5+lUPQTUQHkYKP6npQJDBQVgu
OLlOD8/X8qZp0LxyOWGanJePiKQgRhYphhciN6jEEEw3Kg4655Aq7p+GJ3zlPu+F
PYrW55TTmOh9zBKo90cnERTtkzDcmUS9hLrvGivjMgqGC6KRcXd++1yCA7N6iPQI
5AjMmSSr9p/Mo0jNi2+2QlHNGojJnBxyQ0pyea4QdL8s0+lrDPFSm5pEFSY3vOu+
H/Vs+BEXck4E3AD60d5XnQNm9Qjj5cXE5r00f4D0lwf9Nxq2CS/co9UvovEd7uRS
U/35WlLB1KZSng1LLqYcRXQVqrpclU3UAKY31Z/tRMk=
`protect END_PROTECTED
