`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TJ6Ej+BF4qGVh90khQH1u4tvK61h2xR85iX1dJzUp2UgoqklE104TldPS9SelesB
qmEY73OOb7Fl0Vp9JWEbZVcqWRkroTACVwatgjRIrO1MqwkBammMBVa9Q5EdYPun
rDCLCeAM+TYLxDS6nrR05jkpgEgUnXxilL2kOJ68sKRPqxQXy9xu3+hhtFVUtiLQ
MUZUMr1urqlckXpq5JatJmW+TmK0/McwwzXwFql3g3qKBw1f5tN/d17+OiSAF4iy
BRMwB9r6Quy8qyXtEgUxMu/MP7fybDfdjU70CiM/qcn1D0cv0CM50zyY1DiFEM8/
5ezkm9c60077TQmfNBwtq5hXjPid7Ple5p6sYeJj7KXOg+jAN6F3HBmtfPBz/gMM
TKzuJRnUIhMC8sTkRVU1KHC8bdrn6nOVxnZirGNIcwg12aahmpgc9542zCtSMygo
BnH9Wp9Ni8wVS07uArN9aC1GkLW/+DDpATYZKX/807zO9ZyZ92ms4BtiHnC67Ky8
h+SCmTjt0nzvtBMVbs4nCr8VdCG/F3bfAUnbi6qFrexPTFVWV/DtRL9oItVkhgn5
SfHWocG5B9d+riykQ59R6CKH17mTHka4feU4TI3H6lEMyMU8I8lAPLVWx5wsdfrn
sWnDGQbAQ1lQLppym7uB/derrrR5XvpJkRBMzkJE+lgw72a+bXZSLMsJKM0MPuCU
xRlwHiRCAn4J10D8yDcOsCsaM++mlpvTJjdzeKS7HnqY9yvgwhV19/bdO6kd3cjf
5zm8vjYUzTJU6XbGiNhj42pDq6r6yYGGmvOELmzDOd3l3CIOkIdR9XeG3ik0fINu
0oPc1r1QxdreK7IFzh6W0cOWCjtwaKG5hO8uTyILCZdozDRnGGIjd+bM2lHeWozU
izboKvFzyJYsK8i7h2DNBgRj9+dR0gXhtfaAMDnBGw58hArf3h1zu2R6os/nN5e8
nERVluykoUmuvUvQYExlQ+Kqexv+UnQ5kiv6zML6t8x0moR56KQ7BXh+P06XjNqo
tcf64daWrGG4m0cRKrTpZK2pVqRiis0aDrciSYhGD99IZrEGEAGeBPksL//VlRN/
kJQ5furRNq577JN0fv18pIwxgjZllxc0Gui9NCJdzj/0iyZggdxQy4VnOvaYc5Hy
H8IL+fPWHWrVx1KCuFxK1lzxreRVgbjm/BQVLScA4ZP526Q4ZFtjkrDYQuyzEgmL
uR0JnUbp5xQjZLQBGXkulITxrxlvndLvzj99Zelb6/SgddjE582aNeHTMHeHLH0m
BJN7gw1zNHQuWMd4gUmG5XJHiwvuBBmtfdxM21yUDdpysQSZhswNx3oVHrom03av
aQj56CFgOZEvn8IKKWrLMLJXT4wcHj5CDBEttChQol5Xvz+eYRqrqd1GeoYJKELK
n1kyoS29nvyMsJFgGUvvngww0Kl+vGxNZsifUDJMX4sS5E6nAVqYszY+++SYjNf9
xnrvIgZnnncHVDbgg69kdoWe5sCC9uC9v8O4dTCu3SCYdDvdxwNLCmWrnMoIxupB
`protect END_PROTECTED
