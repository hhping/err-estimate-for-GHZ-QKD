`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o8+TL5s4/+uLzcCJzwqpj+cHSb8fB9rkBrxvpZhnDjm0ygxy0yJTgzohKQVS5ByR
xVMAn/CmltZ8715evVUj2HQ1n01yrAQVIqrQgGQ/TZw5gwLqFrpMCm99DuwiXrM0
KPYtiAa0q86hTSABLUxRKpC1SdvWgUu4JPbcDhao+yWHP37puVXb80pudXDipFPA
SLUjlGVq0BsaVntv6tP7tlQ+TyoJ66ugbCilcBFYrlbUZgAMczxuw9/s+BmgTQSH
cFnsXNZOnEk5jduXIeGg+5M+t18trS/50Qvsjh3z8hLdSdeertkGE77kxivNV09h
QCHoTdqTWBL5GhiFNfyhOtIsCpN6CbWxvoInNxvEVDWJhUUh8CX8BJ6HAwddNbvt
AdAa4iJXijmmacqk6v4yChbmZ3f15jLnJS3ngS5dBsQ8mUCNMJSmOWrvuPh9LxIP
62QZXP4raNMMxVHQDHZaUAuHjUdif433iSpMYKSn3y5WenYSdNDvAWVfcnjPioHm
Epuyz+g75Zdf/yRX1tsOKqHU2D8m0T+8N4dpOZXBspoOIMyPhL0SmfXkQO2wZMeO
ODvLBtq6CzvNKGQOGyWDmVLgBsFZasojtqBmXB3VvoW7nVBwAtatNOcCZM3HfbFJ
FtilHfePqbt4utYNuvaq7sIYnXQprd2QVmk7Mntdm7Pnu7ZGhKNzCuYXym5EZ3Bb
vvDutClTmrQn0ZpaLGpnQkDDhdTRc1ZnkY+g7pz7ROwFMZ78XEg+w6s/ANnCKcs8
Tx1/SbnqWLjQHX0EiMEQWD3xk1IViC2WsMhsGQxAz+BWAT4B4dKTXmy1K9kIEhva
+WeYXiVbLUuTy7P2SqC5PGzaz4gNRQZqCKihWIgPmY8CcDV9H6fZdwmIdpthLH2U
AbJiGdL/Ymy+1BaJ0MmXGnebumfvGvQoWtbUVxz2ZRXrLZv0687OJHftQjCHfUO+
q1jYhTiRWZdsA6XUB5OUkzdGmW7/qMuHOKi7/Og6L6CdL1G3tDoYdk8HigOGZ5Jb
XAVHCQhxEiJVKD/9Dco1lZHhMgCaJ8lyqHGT8pBFaT414Bi1v1GmLRIndr4lzUnz
yfCCvESelzPioHOxy/Cuh/tpCJQHtoeRFBMPPzchY3yRU9BNOVIes48So4qGapI7
DUoA3t2rlZ66JllpyB+ojX+ZlRbGGa0JGee2zwRd0ocLTFm21dmEBvNqVPtgHEsO
O4LmkA+zvQP/YTqsL2OF9xB64w82U7EEMiyAdO7qF8MEzCj1QnjmJQDNdwprUNFz
6aoDmDG6OLwI3oCTC25WS2ioqIRjiA9Sd/XPtNP2tCxI7z/2UzqN8NKA0TlN5uGF
TDvQ2MJqKDPL7ZUiZVx1NK7Bw/TrGAjexRYvna8uE9izcDrPZKXv4KR4fymptFmq
e2QLmTM2a+H9g2CbH9q5XQZZWMH9dC95JU/uPtUjGAS7L5h4KNSwKmlCLW+/BHsh
tOtmHPhEYA17yVTuUdm0fNAnyxssZhVQfprf64FIWM/d7OX7ch0IGg9dQ5E1xLLN
QM2R4ybRRgQCZDXLfH9NC3bJ1D/FTBw8fVTs6eUqMyMofsplxB2XHIIn1T0AZzPo
pVbt2fW7M9U08m35FmNRaKT9siByQPWw9N3zhtsLtu3ZMyi5LmzUfwuO3DcR09Sq
ITJIFsDHVk/RsPbTyykeLBVqXXOlXhG5Vbi6f8xtbTfOhv39/5HTJzud28EoA6x6
XoboqcreoKETaZPLoCcsG2q+fF1oO+rSvlJk1viBBklWwRJXFcRreb9Kru3WslYH
Bu2TofPG3tXd7SDDvPXkAL8Flu95f7cZm6xMiWouG7l/z7atF/c7cwShyMPWhR+Q
WLcEi2jXsSJYUDLr1RskhinxLv5SSzm+S7HCNQNtIJkW931yfofDe9+KlCDd/pyS
Y4Y0UfZwj06IvlTW3Z/5AqNy3euPBqzUfuRzQeH+08n3mEPtb3PlAbfaCQLVg3aR
tEIyD13U2A8QD8MxePAPvwb4QdYEtkDwxq6Ejoylm20hyrv6pnhnNe2VJdONwEjT
Rl4nhb5pZ63T36dMDfJzL3K0yM4XJI/V/yhik9470kwN5qfHA8Lfp0mFo2YSFTsm
zM5vCbaVy1dxpMgZdB9zsKMvdiX6NTiIAEpPo0AT+pjQkeYLs8oivwk9kM/EzaCI
3rhPSfQ6l1Pf+XndMUNGsoiIgqvlRwSm2n/OmBwnQnpQOqKLMerTmaprMccXYkPZ
jwGAbGSXQI2FxK0PiM6prhxvtK4OT+UDBUyOaHBSUJad5Q2kdUz7bhr11UTlsN7f
6J8XvKgQxVdb/TnmxMDRxDtHT/nR8N4chpctEhUm+7XIShNDrSAyOnOp6mHT2E4H
ReRiovv3rvQoSi/30qal9krs5SfZkXrCQAUyY2YFETjj5G7e9RUVjG+eie1trFYc
Qr5All/TiQNYfh5DCqSpMKPPakS6ffPYEa6OWHaT5sQ0f4W92tmSsYdAq6QvnPyC
Dv0KiP+M+YC2xu4pyyzRvZonQqEkuG033sGXQH8dnkYvh37xw2p0FEkkPAZwDb82
auGKRC/4VwT1srvWYUV9unp0J6xU7Wb9fclrzrNQ30B39MT5Jy9sw01DRiO4bIB9
CUabFsVyktBkM5X0Fjx86l2RP6rCHIVKzeJxNWcYRXS/UV/08oDCqje3YCb6qvKO
U8RQAyFesLlG4CDrMjHfEgGyEG/wHcXhGAyUcTaYfN9BolzntdbS2N8bODjbz56V
UJb5vhbY0YawIfQelobO76x/PUHe0m76r61A6m+AJIZD6I7rD+R5GSyiZYiWXBXu
0BFIJ18y1XXpUVWLP8H973HJTr4o0pNdKOrecDoPO3dfs/n/fNSmMEWkqLRspMTm
g6MGPrgX2zE41lWVrVPgH2uvtZHYV46uPVJB9G1CCBrmyNTaEOIhtlh/822QPSai
hOl4nWpVf20VNRfR2vGMe+GvlHcGEteZ6dlasasVqmxi93nlsbU1+80czPLIfibo
ddqhKLzqxPVZjOWBw6nDwzhhfY1EwhEHDOCrU94sEyhF+yNQ0zyJqSy0kkW1nx1Y
IUvGSAAUcmOH5nxvZnXw1Lu8CmMMWFoqXZvfPva793cBdUc4gTu2xIQqJjTdKbEo
4Jotz7nCLE9SHoCdKtj+f2J2TmtQoeL7DEvwrxdGCzpIEZDeFpIBWOpBFkg7V0Wo
p9GMzFQ7umUecFMtQ3x3m5SpenJzeT5YMAviGykQmN0gVgl7nccibTgCMHvmhMSf
hLedN7wksVfBSTI2a2PMXM9SxlXQKCceVioZwjTpDlo04aKT5JC5tCSmaSWErGjK
++w28ZmGuIzSDRvgmlVY14SO/x39inmIgjHEFxfg6Wt3oybnuSoCRR1W7rA8XQTl
80NfLXv92aWjLSiMHH5t16IgJ6HgNDojawW4MxEp5bAULX55CUarggalD2DyUun4
x6ZQi9locWf/7ZqXvNUxyZwPQCW+sAWZrYMfUOlP82HwBw6Q10r13GA733rxwTG+
sDzhTxLX56G8PEdcDoWDzaIBtD4F9mltlEb4rqPBKAGngv0RGfwtogy+JZCZaYJj
wRHoBQA0XBidMmKRQbr1mCwYgPlqCEr+7otGkeum8DS1Bhagyh6t2SGrU/hcSUQb
5UmukwWW7qsOOxbqBIbxQbsB5IZb7C62vg3uyo8SwBH20mSY7sQ212SS0otV/1KC
cBDVKopEnuVaWU5FwrY3AWiVLzKX9iOzMBlhLj3ZeR8rU+11RqJTMY5ZpFQg7Uo+
3PlS7F0ZZf30lafVXt5/GMr27Z5pCfS2OltiGMJ1Tyhvi9wDOS5yPIe0sokB2jb9
T0VIO8/g5a7SDfM/hIA/o2aFQdKtCl6rfdSeWfmkfTy+PAnjDPDThrizEMtkL9zX
lXxDQsjkopAveWi0pQ4CpLaWl161JmO8jOtzljgqGnTQMfKKZ5yu/aKEIVSTICtc
82ajNhMSYeuUQ7688t7Aea+GT8Cy2g43nmLdQchYdsnZaP6ZK+b2mGOHIIM4RUUd
v2BkfIkq0g5asIuasitVlc4BWhDh22A/bIogLB8XuUUTBxUQlLy5Qe4erOgRyB4D
vqoSnJu9cQ90wDrD0wn188d0FsAS4+Z2jVWy4AOPYNYPtYLOJZuO8lAtb62fDrBk
go7OSwE3np4H+ODY7LnqnSpKhJzQPUU5RZVEc7hGSjNeBCa8Weklm5dfigcaJV/E
rkGoGG0HOs3Bo/04SQGzUi3MOhU2L+T/bFNM6/V0szTncAbbRZewiXiKCTpV1oVN
SJmgGMOWI51iGLhP0PFxnSRO6gGNTw/ak9F95ZVReN51Y/CFjeEDgOToG7YbNbGf
SdZEf3A43qip9Y+f8MR3xhrwxHiMKJb7ZGRP0Giq2c8uJHqtnsLC5AbssD56tQjF
vpqJ1vKK/I+hUKxBEWCVuLgyX9eX+vfy5zaBkiqZPTbFwS8QNuDUWqQL0s8r4wr/
0klsiOT7xdVWc7c51dPjCU78GIvk4xtrs2YAjWvq1cF71sH+C5XeZONAd0RLlWYs
vsblIvx+nPatbEn08E3bjEhH42MiefTokQqw9bvrCRaU6HPjcq1LKHz+hlnh5jzH
nVMOSf1IWi1UyQrHf4qmYDPkzvOAK+lWznqC9Q6UNl7615iHFXjV4DlNE/6AG9gU
GGO0GoxN9q8IOMOluDQxsihM+8zIB3jVTP61lcxIfrDBa4a1HCtGBLrNe9jkWhyJ
xGRdyRolR3Sw7dZ/1go9LbkHnbSz2seGNsmHnwxMM9E7x7M64AZiZWnoQHeUoZvJ
y/sLoU7svmY+jhlEKQHsDpBqQzZUbEsCr9DLT5mV48NLipWGkwg3ss9AyFY9fBAL
g8dsQ5d/7mqiP7Zjau5ZOEVteucuX0IaqX70ZUkaBIgK/KsM1/u28VwfAXnBphFm
/kfFZXRyp8bC2mUcCx0TtZQCU58WiAmY90LketI0531Ul0dnVD/5t/X8Wp+7775E
DmfO/oQBmh/DvHSVA2oxRBiCY8yHF4hmWBY6tJMz/3hUjCNY3eptUcIb+ZP1ok+z
7KMdySjxSmfM59KgB9CYHqjB+o72NVj0Pcyzk4GsZLTwGHgZsi+wLC918lEXpjgs
NYwTtgbMmGksdYrGj2R6AqZTHt7Mq9qsamk1sbjC9O2Z0eJr8Zd4bbvUp90U8cU5
F8/6Pq3+rFeGKH6eUhu6Pjy1wzi7FeFgbORVpa5E3tqhG2S/GVLwNSSNL/NHCL1q
A/+Uaow7LcldjzcOagp3JJTPiuOb+XSaoDcsVrNJTKrUMfH7VO2fP/Ve3uvcNUSN
Hg5h/qhPsszJ7Uzjv8VZOLgBoMgX4lt3M7moxt5+AHyk6jA9k1URyImh0OMCYf+X
KmsTMH7yIat9Dg6yOG+16T4JB1VHzhlg19sqU+aidtPyMf4WK6aKJtPouUX3xmUz
4UI0I5LjVSTwVF3HQCRnMphodgQVFjOO3LRmUcpVALIOkYM6AMrsgeb+ANBs7Kss
9TN9EnWS5ITO7o+zmx0bG6OvwP4yVfUiirAms+Sunojw7oMg8nji6Tqb8fXtFv5/
2H6wD344+m3mnkxQCnAukY8kcbu56GaVrIKgBtq7a/ZdAQN8aK7gDwbSsVd0VDGl
Po+hs1y1WgZn2q+q7Yyydl5nAB/Gtere4wFB/9VrmNakTGypUJl7Wo7/BFjhOATl
vHbwAnGBS37k0Z0zV56LcAg8dcTzw9JnSVU71GpDG7vS/AyTPKYO6lzqJA+URaPK
Umvlnti61mw0sScZR8ZWsmLH9Kv0C0IQgIX8+ZShfx5PMDbo3kX2CW7QAkQefpHU
ColD64+TNO6mBdLMktHjkuliWRwl3iVgTatqNf+V6GBO8kVcs41m/OnMKoTe17SK
FkvKDhrtYb90/T77xRdP4ksqzrt/yrOEh3BE4BnKysBZxT5hFtpm4utSgMBUQRJZ
ApPjbYlNupFP8jpsIGrAi4xqwaKVkT8ZcU0Pit3s82DXSMGPTO/UlBq7jdwRAceQ
fFmhYWo6SauuzTwCpCRFNWEgbx/WAB4lcpX7pLykccl728aFnwmGG0bJmEwteaOH
A4BJsl8jUExliBx7CHeCnw2xd5abCAG6cSFfJSMlJgywadoC2+8zP7rvdShVLQjK
pGxp3lJUpyGGS3M8WoxRzS5orQbV1BXGuLw8r8DC/UkSKWKkA8k+RmCxbT2B+Qti
D/M7ZylDeLhxGP6mYhT1Xr/70SOjN9447sWwYt0qQAcTF3HBfvKGfTYO+gVtbCYQ
xHsF84Af1IoauIAVlabAYakUSaUB20mZNvCm8EJ/0FzYRdxbRZA2J/9oBCNk30eC
n0+wkBmXce8mE0x87E73jrq5XXpG+kvgCDPIX0O2+fMawDR6TmMT6rjT6vhwGBYT
3OJlJxAsqdrZdy40IvuDt9boQEoxgDys+PCNrtNX+IVJUalgnTDCdY7YtUOgKpxD
pkbA9r93icfdH8DXDVAHkNPbsRtAWlWPeGDG9WmnV9rR5Cdue1EOYLtZAnK2kO5L
WMXV3xZO9bQm+Zy/ZRx8QM+g+MKzkchWmWImjmclFjjFRkbUuf6U/HNhvajQyKse
iYpoj33PulYjit9+D8giQD5V2qJ38grj/PSdi4uTr2lHPIUWefN9M1Qs1stOhjpa
8+dlgVQ2InTv6gd32bu9PY/I0aXNPKwDx3ZBgqtcjXUMu7USqI0pR6JDWM2y1hKh
1TKpyV6t0VwyvI/oaGaTl4/wNzEOj8UCwNzsLwamXSTwdLj3JGgRAoegjji1GvgU
ojRYP9lUJ5Y00L0Z6IzmwvZTwArIop7aaEPE4ye3U1LRHuLMFoxHColRcMU+k3W5
P7wcL3Schf3gXfRGdkaEe96v2ncstAyXUJUQqG6ONXMneACci0YC9V2QEtczSVIl
2KVzKV40QlsNVu9kOeXbY4rf1lDuvbrvinoWLXvvIb9fLW6yLbvG0C1Lt+8rSNLA
ZRi6N6B3jf1xftX/7A2GylyD1jpEjowo8KYCCnxIBpXaZgD2fkNoCXMiIvBJsmdU
ZtHlJw9YUon+rmKCz/tDCXk6e8hGRsvPSDe5fDsEipyOoD3skb6AhPgBIFmvypmu
psHew3HFdJWShTrEzdEQ5peQxPsbzoCCRQ/XR2I9NxCphL2bGJZcrnpegU5yiEge
bfkBWOWg46/cs3m3uZUe801Q4AICTAlxsvoBwz0ryk2oFsmuD7PBH+ULukIG+sGA
wSaVoiB/82oP9qPshmHPlFBolfb5wd1j2bifsmukiJ21Z9FMqzoh848ruMCyANX/
6sdH7vqmtrt9U1H+4zc0ORydN1zWhzNHMTpPvBTcY+vNfXjYSetCsnXrew1G0cvJ
F/gfmPtWa3zHjznxPyAnBBGitqrtPWNaRhcFBH+7fBPx701fSfOBFordZ6pbxqpH
v6dpaavIOgnmwoEhj+excUNQLMi58rtQrr7xXpwOMmh+OSdwNeGDfa2peHdIg41Y
2pa8B2gclkIGGLvi7LDKhShBCQq8iq34z/xH4VNHdF7a3UnE+69brScHK2iuKn/A
yuDucuuF0vdpD3zNRWOXM5agVcMwYjwjw4eV3onyeS1cKPFPlVZTxHZpV/ruxi+1
QgR0dlz17BF3Ug2jTFkwhr5qPiiwlkTptBW+SZphBrij8e0QvhaWzeO6azzx8Gh0
GciW8zEYFx6NidLYFLC6jkXM3FKF8CM/flnBvh4RNgAwadT+v5Ep4dl5sxvb3Bf9
Lsf9m7jde11agr0Q2nKFbMd6oKy0iLRPolJbUkNVBBWaJsK7YBtc6ztwlc/BM83t
O2EXv29QWIdSp8p+OWWANepa7oif5biAO9qdFLfkUlualIk10y7uE95wj/GsWW5h
NJUI4KoWiDeFTGS204kyZUPZyzdIfeB9ZmPtxik29IQ+d8olbHDolKPlE7BSL5Bp
TMNC0OppY9yLs2Vd8uceOoO4V6bu/KpYrDoCpbmicTv1Da7finrzjdsJLQbGRnwA
sqK2+/RJJ4ch+gp+iuBGGxSQzbgDorTLRzD88f365mnzQq4XBsAGHgimCXBQO85g
Y4/Zs4p2/Ihsm1nu5AcohZFflrjy1kgCqPGXe30OlGxvMYBSVzYfE4Vd01wIGTV1
8c2HDHi7nJQqVn3P46ifONxsDrxmbPsqc3p4Plh7micCvVe6538VxgKXRo3d6VN2
aKfKgwLywtfyE4wu99OFr8hz34NiYWI9r9Z/TqQMVCU34k5pdychSe38VgUrDDru
TvSpBXnkPkPvUWoJEc6Qzb2HQrIMojed02vngRB5ahWVHfuEuOBdHicse7m1bgwQ
Q1wqy6eWb3MUj74b1KJaLf82xiNuNQ7eW96ruXtLW26ww2NvpHbA8qkUeFY1MHW6
pOGF2rKq3GV0hHblp+n1OolieEMPUoZst/apEBmfM0oSAiHdIOzS6YQKWqvAn0Ql
0dKvyAsjsHAYvVoxZWh2erWZVaRCOeadUeqw7EGD1Bf2tpjT3mkFyJNNIExdKBGD
8/eq6sNlshdRUum4bSaIJUefwTNvLugPkYx7w25CvBol0FHLGvw/RogCyJ/ZUe1T
VdY054Z9f9rsDrNUOxFkRx7Px55xnIjo50yUdAmCF30zy6lQQ2emD8hk4NpaVmRG
z6axmIBteaHvh/eE2WR4Jun8BUrtl6hqYUzo3rl/IQf4B3jOMD6aJgpfaNJk9+0v
AfukU84WuMCcEwpdHxmcA8VOYQ4It7XtPWrEcFD3+TIihj4zHD7391h899KTHx1p
/6yvIcZLjZ9yKnOeu50bzpgpNUNv2fAcziVx2VG2rRa2PbqiNj4/pzqv24xUMhUy
10k5MR18QFBkM6yX9cLOrtbujaIbkavmxapVXaJ9WHfh9V1Gn9kncLfWS0SibJIT
YAFfTcuHCHuTjS3PU1EV/kujq4rHEyUP/SiHhMkhkttPrrnwkd3OWuBdq7sQWCF3
Lqt+2NHVFEGuMVgkjO5I6q5p1gor7gdiF/YnENX9alnorWvq/mSbz1lWUtY/5sh7
xmig3rUjLk9kHY/rLGFZ4r/l+YHfNIte2XU1+qG6ECScXfVj0g+6wmEbD2PtXrJO
4tg4+qvDivIxHV+MwDgEyFpBd5muBUYlOWNG9Yk6vSr9hEoIRqUgaT1bkSAoaRmb
MFi0+/bWNL/K5pTf6Zb2jQoBvB5bNto5lDhZoRScRHye94HyvHTXmYu7p/aoexFY
Cr0i4GFoT4J2RgMsX9hUL+okvDmdpYl4P/Tym73tKuxz3DHUgnJHYUSFUH4V12RH
mAsToQKWRytGkm+0c8tNJd6Ci8GHTQTDCCTZrZSaes3V9531Vizt1kgF2fpD0phI
yWiTZs3Cv1vGMhHkX74M2Hdnw1nVG79jImHcQnASFceUGB/VXM4zZ3DtpHKGx8hl
LdWbcTs0Q8+RjxSxB/+bQluaD9l4C71cO2t3WeiH6xVC+hmdLmhfho3uvoU6CToW
kztGeTb3GOHon8Uqc3UzsX9cPhGrta7HkG9YUmPNOmiWTym/opKZU0IPm+LYZC2U
B9Dv0/e0MhGstOviMCOZBf3uhC8YFQ78GZt90N8FS0pBW3c+qNEaYjhzf7wdLoMl
07hAl4wxzDJpeE13RwS1fltfIQSRFR564XqFEP8h5WCaD7egOjUB91JSNuZ9MdkL
HLaA/31Jkq1hq80cpqhvfkdN6yH1hWUwy8wpHsa5K7J1+qXXYHW/T4bnutLYTJBh
MenTBwFS55L4MTS6H6EEoCNPVb+HR0DQVVGI9kNMXpR7oDvePSkxo1NipqZ0UGGk
zP8IslcjiorNeDlw4N5NdesbE03pua5FREif4l90Y17MVxsspWbhzIYApPc77zPd
VHjARS0o8Omj8G3BW74R6tlakqvwZRb9DgA7TH0OWWjyO3SZltJOhO+3lWqTtwuL
HX4SdsTVI/Tu23FpVYM4zvEMnw95WFhG5wvVSPC8ua1A0wPM9A/DSZHHWZPk8Up6
Ah8iHM2hr9kNhJH7zjROI5YITVGAMd2Z5NuM1SgGLlQTzBaPKnPbtNkLe1drskbq
DbAp09mE2HHoWMJ+60HEk9z9fNQznCc2vRqUrzBBZ2r2IqmtriHPfGVDpr/dqm1d
Ov2ZnT3Zurvn7xjsnpqHc4Wfg6nl+O2OrmF+/leitdHix+EL41IzXJodTMssKICS
n0EjN7PBJue8pd87KG8A4mvbrGJuOLSVUyzmvgpVLagljAW9iHBdB9MWMDm/vR0v
aDQHfQ0VPdes33AONkp0W1NolqVVcjZbIYL3FoGnpWk6Hy8gqm/Hsbyq7dRmRWon
UID2RxOhJId7i2fHrKNhUPplj0ObN1npgLlEjC6CPf2xFKC7GO+p8gy0ZAP7YFKv
3/WEY5KTQGp2iDmErZfNLMJjvSV+O79BredWUlLtaiHtg+SqsKHLDrPkVx28cTSJ
L1Cq1W17m3j+Sn/19PR43mEK8CnrZzbQRb5rTHPNUUtsj1gQtcjhRSQQ5g4qUmdV
F2Yz35kld4A534GDgMtrcVlGHM9xyvgn3cjCek3fguZqa37ZKJogOZGT30PIQ0+C
I4D0mX/atnq3uxTL16kwxAvK9SL1U+acngA0b1qrxh8fGMGrlT+iLFRZM53kIuWz
vLDjojqWkCM5rIjL/yNms1b08dk6mcnoRjLz9pKOg4jHUiSV4Wz9eoiffm2apubq
t7/wP2myWz/Ih1+fmtM06Tm7y/xwy14ppTmZOIuQa8WmtQIuJsNxQwJW7x4Rm+oH
mn9BhhiO6RDwvCYX19FCREaD8NKuenRjPySGsNDAhZT50DzA5V1JG5Zoq8AChbUS
MBjhIzE4mDkBTeuvObjgNpNieE8DKNmA3oyrIIOrFg4HCapHOyU94pBGkkhR5CtO
+21BHpNyDMGtgm3L6hPtcGmBX4LWpv+44mfBihtcIMDUZ2FaXBFeMRDM6UhRmOoY
7XUlxK0K3/WiEQEx6IXoA3Sh9FLxj157ePmazRx8P4GDptE0oERx9kxKf1CBWRT9
DbD7N5CfVlfgDpm2VzwOGspNAcxe6OdrnPs+wTrWLYVtD13Mgth1OMfx/8nJdWrM
Lq5NmB8XZ0oIEW2INuWGNTKFdRaEe+irPArFuaki4N3esfM5bvYMPMtFZEyRovLN
rsv1z/A0BAp8O5gKHzE9mP1dD5ypvU5oGWjPcOoYuYL0BGMxMQRZarvD9xfoncGu
nc1V/uBwTkGdxTwPt/62VrmiYYYq4XjbAZIkyDw6T58ceQSicTyOAQc5pQYC+P+6
NTodgPE4K3bPBLQTrs/RpFaLmkkZDa3BYqBfIen6RwF+pu3GECKzHi+hbr8bFzw1
95MZi8rsGBk31xBw3xSz9XNRgjbI84J1+3yG9UnQWr9XimM3+6dSekZwqn0kcSG5
3MPyz9PRAZcIQIFBK6aW6A1ZjSsws37tzGpJ7K2oIeXeaimUIYYVU10lMzJPBEsR
J9TAKud073tuVML8pWi6geKbjVkKa8hiDpROTcQjIN8iLL7RqTcjBYF4emh+VSWz
zfljE4N8FwicxFIt6Zo3le2YODmrGUSxORxvTRD/OIEr5it8/q7hSYqnhumGmQdd
aAF0N1D4+Jjq2bRbR8UhRiLaCgwhms9PclUnqGwTDwAKfnpZPGCFdswb4+ZMboXi
lO41TwBkBi1cMOq7fUDb7cbKIMWXt4f/IQFLHt6TQMnHjhJKpdKmHSevJCA56BdW
PyNRkXA02Rfi2ErRuJzmC6Y52A1+UAYSQl//sWTwUzpo8IasalFSgE+NNUGlTk3H
ldznfcXEUsWG1knGUBTl09FKSuncNo3B8uXem+C95Ctp/0ITDo0GSssgWVHwVn4n
7v/TBidZBBBhQ5hx+fOoVobL3kRjwhl/5bo6W0aBNcMvmqT6I+QqUgn7iWXuZLnN
G6FE9Q8QUZzX6tMPNHty1leHeCaeXjOWnaqsFp83CEX6Vv/B2vLksv9KfqctWz3Q
gzJQPD22jR83XTR2jxttp4q40B3g2pBFre4I8/sjOuhAtp9g4CcbzrMaDersMr4G
Q5XQlnUXdhEtSsbPfm3BGCcX+QFkHURRrLWiN95j2CdC7YsVxif+VRH37flGrztu
r20ie3q4hTMqNZJnjfUwJpilIkCUb7tFkAXAZlKxPm6wgcseFpOOq/v2R/leIv1r
v2Twa3E3RrLJselrL8Hvs50SJ3R8nbcw3jEpWSKzJrXOZjEk7qEWWWSqeY2d4Iz3
vPRhK5UI31hueNrbZ1O96rg5v30EIqb0VRa+MvYrI2l02n16Ep84CdrUv7HIfLJ0
AxH/mipLqJJnySdGwHPYU7AJddR2BoBHVWl8RJc7rpWjPk4o48Q53iCoSGd//Tcw
bBXl5T/TC3RYhdPtz3Kozijvqvhi29Adfb2PrxAh50/LjEaMXJTw36uSWjwDH76v
0grsE/FoILX1feb8nTO8XYn6D0+C8gIe1pcYQWzWOpKQf11MBKbi/9tQhGFmv1JK
6E5rSuNdDTz1LLIL3fvLR55U5hkYIK13mcFk8OvDhEJqEMx9KzOQMelTy6HW9C6c
3vNWXaaAoaXxNDNZtjJSi9IW+J9cyyP6rNkjde2YoGcqFG6g2Qw6BQ6RKkH8ZWQX
pvmWIFz01bfNfZxGEzBRuZV/qNHdNslrm+1EeKZWzZEn6WXoKxCiEt2JOW93gTqX
bh+0F7nHZeX4wqX3Go2ZPWWcD5VnVPSs/eZBJfap3n8LfP3fYCCeka6pqjPzdUum
vLnXDZCWBtUvcnJmQz2T4cgrxTTU+vn/DxhgRTdiuv7ZdS4c8phNufNFCFPTzi6Y
QBC7gfQIZxmitUVjzgxWuSC6gJMQqIxdkpDuTZm1inF4BBY+RRJV2QHQpJl1OSjj
g5iVYMCnxhl/qlbUIsDL3RMzpX8FFFEPGRLtR28tUjSUMbw5dx/nSNRH52PWP9c1
ZEuB+AumpkmQCpjwT09whoYmdY22w0zZn6KgkCuFdWet7XEvFVYrXFiKxkuaiN7d
qBffSoFF9+jom7SF2FH3EAtrIHoBcRLHL5Uzso7+7rBmatc6C6nEJ2zQmW5eFcui
4CaeCfgJvpo30PPYAAB4gKGYR2dCn4YRYvRsQ4fflgWieOrUo13MYNDKVHU1z8xD
has1uWDgvmeK63AjTSeMjNkpFL5xw/HlcPokhOlGOSrOMUAg+LsVtMmlHhZ30zRE
aj+pOuRexi6y7emvFAYKsQccHO95XXXPIcH7iWScLLB3ticgqBhQddwIdBajrBEJ
pEjLtyUmoP1gt4DW89OlPSOzQDEgGmyYloG+S9nVLD95xoSXmbqx/tcLAFy5lejq
GoU5t0cFbS4/C6chc4Mj/vw5W2cb/OqlYRjpKXQzxBRlCMbZ1Lad+FF5hIa3VpoX
AJoSCMJHdGxLSVjLO/JiNYxOB54vB/TKsX3Vw0ldWfgHInM7VUnVoNHxERgN9SIv
BTzu3ra3vO9bOAlABFf3j8ha5p+X+MSjO+ryiQPDsM0+bde+aUXpOnjKGZZpLkfZ
fOXDuZgut585L3WUqvFGOiBIYy00liT6/7GvnKtNV40ERY2MXPIU41G0XYMZ5v3q
GjQEg4jrrqJnhXp6+yUWdzi7cAbaMaGvg3v1QgQWzJDIJJKHfjq5Bz346hFiIAQT
Ds/5+XnkX8MZgFZkDmxUSbw8SanMe8+hLnrEvKvUo6Kw2JTj0Cz2HkQ50Q1MSufo
xwsFYhr8sSN+JNzEBe8F3rWcFElBruRPWuZXRHzJg8oEUn8lQzgjol4G7nr/X/p3
1pQDR7+qmcaUWkMdMNUgD675db/zJKxoTS9/t2cWqqBqm7F51h1AaSSCNQ7d/8id
Gm/5g9bFpSYPXif9EljgDfLuRyJ6nhzjltyswFKsCgByUwQhjWdU53v3bMBFvT25
wNj68K5a4zvGXovoRgAHiLgx7jNzS/cQPyOgIA4XQ099rj/aiy98R3QO+ShWjGCk
VQoTqQtGC5xSaVm2I0d+grncFXAN2qMpPr8a9cxvfvEwrYsRSzNYxowC3JDtZ863
RZVaL4jFyC6IIx9cjcJ5rEWl5Bu9lsXXYFrXi64itmfrMEZq8K+Dbf1A69Ko9YIr
3wJtx2aYyW8uJ4xwUzyjYSPjL/4eZ0NTJDHN3NDwOYA3NdgUbWvPWOLc/gqMo+jZ
Hw2qVe4kfCg6pWVXuvgQstUdJ2IMZ+3sawRet07x/mzmm0hUwLC+JPes0jJWlctb
pf00wKvRDBETOcPczY0T7OlQYr4YyioLoWQY6sSsLLJ8M/Ordhu6Mgkez10NTDwa
8J/4JhNqv+4rjWIHV/Z7DqKjSBlhcJKGUeCWcFf5/Cywn+v9z5w1Yvv7Byxw5yTj
SX2LkJwA7mldXkcDmi66wQFblax3tG8xGOHRQfb2qene7j0vKYGWczaN6P75Iaec
QhIVSMy0zM6mhBjyC0xBvR4Aixwj/qYbdUsx6FKjt1xnZha/ERtBnS6Hd38H4vjV
13wz88G43YsvLWIK6uB1e+XVpcipCbjQmpk0nV3oXuyD8e7N8/KCLHys8biC3B8j
wrwsw9ICXnsNfuLE+0mxpGFVUOv6St/J1S4+La63WY3wMJv+KFubBq6SaoluEHE0
MtqPxBj5HLXIjK+hKsovT2hL65NIeSbb8ayO1NrFS8QJuggR4VqaxC8YPZV1qJ3b
JpdCg2uqvhQuNKGC22iC3hmXfM+WE5vgB13HVT13rmnTixTJkaeaDU/NRsbIW5bi
Eek0wl00VvD8TBNvI0PG9gmNETtscJtvDQKeBZwUTbb0hirPtUy4NeOZYpNo8kmi
uAEbiZz6K/BcZWe1sOYmrI2zByp9zVXgCBJ6KeBvdhcMpdzkYfNC71OaHH34qBRm
RuDV3umJnA49hiu5EMLzhqm2wN7OOD97xPY/Z8tj/9CyjOe5GhcsbnxdNFb3oP0c
r+T7foJw1fbYJvZGwM1dliIGz9FaA4xbbNepq3CyYm2ZzGwsK5nE4k3jSRyaDPDQ
ft2JVtvKgfR2LsR1FJaAzu1glPE8BjjPycAWj5lNeFAJ5DznYzF7FwidxuIDI0oV
5zd/j0Zf6bTq3cPCyjuAkKi+g5GnR6k7qFKdKstnPq1iyBj7Bpfwo3eVuGKqVxZi
u7GfJzyVu0pXVvVOE6vlCzcWdDiRQ3Fh5s6EFjp6tm4mHAW3bAtvrOKla1KSzeaP
7g3lA7+GV5H9JH8LErEtB+UAkYBIX8OQT+aPHDH9Y8LU24zm76z/Cqk8nJ3eeIRB
0BL1SNzTolLx6R0rMzaKo0CYAfxFMvV3xqhBoMtsqizYFjQ6HBaLsFJvQNztYET/
tzirjCLei6qwdDN8iPu07tfmOqUpNcaGsRaGFlKQ9P/PM6BrGLS86PZXpkGmRrGU
t9YSdmeADeaeXI9/o2zF0H2U1GGPkbSANrEH3DqSQ1IUqWN2pgYAGEE2HiarjoH0
ipVRYfUe3cVOvqIqzIFfhCnTsF4G+rwUdcJddlFYJPS4dbSWXC/FB5IoP63UdL9W
m+Hqmih3hMaScG4P31oZd9jIX0jX0pn1IjHd4ERPgsVL/BYMKZVPjRmxVFkoTVls
ZX1WEmFqJWtnSO/QykDbjM7m2WV52vH73CZtye0IAS1wbugNtjoTKmyakAh99SF8
onTau8bbeWV/NXTwWTWsxv/IaoaABM4gj51sQrYytCGR8g4ZQte5aYA8BZ6rT4WX
4nrK5Ay7mxYC7D7do3N/8UFqWtFzOdIcNMsVPIVJdWUkTtENdaQpshNyM97fq/uq
YfyXQElgQdDKR5viqSygm9PbUkWsO5HC9p70TNkoT71CSYl2+cVTcqGyAvkrABHU
YNAVLQ3vOuBer8FEm9tDvtfSg48zB2j0hotED4RdzOXAH35K5THPxjKQTTtjYj8t
V1w+Oz5+GITDJcXkuHef/hGsE9EH+lanIgRiniTPbjQ1IbBWTbcnh8OLpSe6PdVL
seqtYQ8UAC60d+31AZw1xQPF7Iwsn5hrle5yUyPi5N9WImrpFrajOcXlhOAOjcza
V+4FpFHdec3gcZH0y3YnU/AHhnIJKd6VPzQnZzn09DF8IEm1a6rg/QvhyffMN7dd
4xZbVZYYCFmTe7BjphqCpHhs0pTNvVnFN2c1y12eCioWJMINcFCwQ3XoruYbecgW
ur2Fgcpu0ehbpWAxmyyGx1BwBhcWB/gxhdEx/Kf0UU4K4nPxiFwR3HdugjppLLyi
HxeJSZKnDlgGv8l+wHF1ll9Ag2K+Dz2zkPAQuHagepges/vPSBya1LJajwlwXqt8
CfW1B0gZY8XHCtYUgFFkIufKQxBu2ZL0F0V+nwcixSKCL/kYIk+c1yIEU0rDf/L8
wHPK9RtyaHzX3PU52zkGQWmtOVean7wV0orE9eDkDtOsForkotH9xkpn6LFf7BJ5
+EQOorYw5jIW+QbaD/aa19Iz0N71LGOH9LeP7PG1ubajaI76h/sI6JrTC4v45wL8
p+w8zXaVU20Lo91i4eXh+/iZajtLcQiU8u+VN59fUwwVlvfROQwB4dNNG4WUQyjB
yQV0OuXV+WcUSZ88xueim0jV+w5gVTdngjGhDXojKEmSazE5woUcTfXt2MOOi41F
0nxA8Vqk75mvmCyEV6v+2Q==
`protect END_PROTECTED
