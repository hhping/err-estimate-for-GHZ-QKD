`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3VcGr8M0X6uoKC29BtQTdZYfIubGCc6URas90Igb8LazENMpm8mu21V1V79sv91z
U9G/YKJkibVg4T15UrEhsV9FTQ4zAJhDLfK0ZV+FPkA8t9FzsU0k4UisUGrgqISo
32y8H7LNkSTO2mk89wowNckZ6scnnsLx9ZqiDO83dG48Pl93qJaMyPiUdoVGNB11
xr5XG3FyYz8V6zuDOtJEx3KVUXyauFFsHCKKf4JAHuLjny+tjmibE9fZCmeyBsaX
INJRYHK3ApRk350f4Kz7cIenRP4VrvnS/c2+fwQd1VDJZbng3XY2qk0VhAtkPjgk
t2ZdpO8fS6RA+oQLpUazgGaL9EviX2Wfx5pob/GJXFt6txhOSokl33r26YsBwkY2
ksvYm1lHTSNDKG7pyKg+XWAawe1c3dQq9Ddm3lNr6BcbXPokHmSNp2/SB5pOOaag
NCufuKALouIBICxPhQXDog==
`protect END_PROTECTED
