`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SEKrBh9cD88+Z1gPXTwaABQnjmBbqMfuwvm+v/ILhTmykIaAdoXNdih82bC5WwFW
wIbRuVgX07rCAzqfjNBCaQqiNgFsvmCrc/BGQsO0qAZUq+pWPKlLq+/HPnGz1zU5
/Yi4hWor5+sIuKJHOEpYImEmZ7xALxgWsytfpu6IMIOWY781zzRGKiWabJQxAmT5
o5Rijlxe1aN2+0moxqUTvahDpJRw+dUpbari9GXpQLJJAgGmgZ+xepazsmSxP7r9
Adofq+MejL+ZfYySV3PfD3eN1Iftf8m0ZoNX0IzJpF+/DlV0QOstd4IFMKiJNvBU
2fEEoM4tab2fmL/PkTpYMO+CRJADi+mhe6hPUxgrUCTC8C/WEgW+v+jkrzkaAbCz
O3Oakpms9nrFe2RDFm5tt9NQTgkaQLz8xHgpbnu+RQ5blCWrsRd8JO66FFLXaPBp
BiV0KsPj6/y6PRcIpA8nlESOl4qmOmQfZspVDxWpIPvFczmBZr/gJR1InXoTzbV0
9Fw3qK/x6mMl7pXjw/7soFZESx3azTFHLrP/zOvz0gy7N4yvuDJmAzPwAoLUqT2+
zcDQtjVXapwzrc5WGGW1y01XiQ3Wwb6U/ib6bijh1RG4AW9aZCaBGn8dDvtl0jRP
D1bVrwWm0Gr+vovUMPtnYypTVR1KafkUfBl2V/jSUHwBPt3MUSto/nPE5LPNZNHb
41NUruNOU5uA5//bOOn6ZeL8zHFx95ij0CM946ipmIZD6mwPh18cL73Mk3n4uDT2
zVItdnF2YogOhfKIKAXEC74xQpxpO7IQj5kIax7CadpTs6j2aRhXfhVg2lEG/XrZ
+OlKMp+CR44EKdKfb0grVwWQHWkDpUXpzVlsuuM595k=
`protect END_PROTECTED
