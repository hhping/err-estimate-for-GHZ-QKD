`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wabWqaZnxZfkohz93vZ/yQzZ3WT1Uwy8aNanvojSfNNdiw1IXPvJ3pm7FDZOGdsu
va4y1fGYjR2xDM0rv3uwS895LydSRY03zyWmDCcrYnJeSO63ICSAprw4aA4doBMY
kdP5K3SRnicqm8ZF9vLzk+NSd/DdBOfpMczzu78P/kch1IRSYUUsSOEpUJiNqxGH
grh2N3BVm6ZznwznlQ8+lXUMkK1XB6MLD/Hxm/15CA8YpOAHXa/XZiIOdHNsqWxS
SjaRGqGsQPCBY4XTtqRhiueiucr9cFfJl82Xzl0ZWPGGBkK6gIh77/lcV04AKOIq
CdiL7bq+RpKxjMYk/wJ559fSQ7o/2XOkVpfwHXyvgt0fryJlIr4xtFrFFQklJUkQ
a2DxkT5i1X/86cvfOpr9qDmAwwVAOXZGQ4C6gij1oipf520L96f3p1U5s/CHRf40
bunusWlEMtX68gQ9VzumpS7wb+qXWVBGEVUaq9pFkefY+RFKqX+BLr+kMnM7Qx9+
scptOjU2QBx+3hkcFsnPZlp4yRjDeeNQwMuNxCvC6CbBXla1/XU6sqX321IRo6lF
uWZ21vIK7DTFjbw+3JbFgDWMkyVzSJMM5lfMVFNAVPA5r5Xn9SOKcNPiK0KiVl+w
yp91lfnwH0jEnSDaU4YgFxE/TBCJDRMCYPemaLWa18vfk/CNC08VRQPg53+xSmc0
rsRSYRYc+POEIEH2OuH6tOE9ip4X71r0CfK8j69QXFM+Qn6LQ1UIIgN/b0CbLij8
wq9V1Bydjl9fwIsX1Hbwkio7WI5OQtpRwG6UbNXV0AwFttKVEwEzhQShoZbe/MwW
uA0ZlX4gUacW8AwxR7Gqyf6iNozfMmFfDKbGxfM3QJ1zYu4AyVqLeLN2GDiMgisl
Y4+QjxpiefaltKlKcpsnFwckKZN7wmDPGZKDrEPqIIiOjlj4M9MHTeQOveptmq6x
/7ObSqHVGCZC/2NnwLebI4L+FC8Gre6cSzJEk4MycPD1CdJafWKHxUZoqnhHT8nN
PI8Phka/PUfs/7Yz1atbwtWXGPub9WH+Ouj0+eu5uxIDy28MyEi/0HxJnpsb9nKv
3Kl8Qj1H7MUQqBPb954Qwro2AhpcEndFacauUQ//qS3HSV0QCsIvENZhQBI4+qpb
AyUb8Rt5vVYM9Eo9tczwunNDZ6lInNwgFI2m5E918zb+kAgr1rjTJpA58v19dPt/
0EBQb5z/q15DCNYtVuhU7g==
`protect END_PROTECTED
