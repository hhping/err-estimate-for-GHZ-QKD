`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3RVQ8shxZ6YUHHYT1MjR7kJUaqN80+PHg42w83uLTmZwra81H6PvCiwiEk/qQfBX
yIIizhRCtmB4WNeCVooDZG3z59mCYp1gVIUIaELG3YXvbuj+YGGldSYNb+kXRY2S
QWKAD27cRucmmcYXhvssNp1epSgJQNehoM2nc2FSZfpNgIvrP4vCBrodBoEiLCXr
mqX9JQNYmHQBnOCvC5O6rrhtXl7NxXbl17gyN3s1rYsOfOHRqM8yYRhbPZzOmSB1
Mas75TNEAACHSvY9BV1/rQqh9IFhTBNRFHRbop3zG5YUZMDcBaqPQXm60fACd91b
b5otzuaTOkggbK/3KEdBJ/m99vFlVQE6M62YES3ZtHOdFqpmkSGk5Xt1d1yB5PIE
CgZcwFu/6Bxgx4w1stKkc+KIxbq+muqkLgDBkwupLE0EO3shaJrzO3EFiCYd8pug
axYdRRnseuTjzBaPi0Rjec581kIp6teNilDtEbj/+KrDmrdDQJV2ISc0Cfa8IP1G
kIxbGnf99jXNpt0ZKreIi9wdcIgGQTbtfj3acCJF3NCbJZXh1WgnpZU/vuxcvqH4
Op769Cx6nhpv0qSCfa+6T+06otTvfm0nFSr7Sw30W3uaysnjeD89joN5wiCV4ogm
kSpuLtdVqGM4N86puno9LOP3cJcdQyszHpbuTntWRHQF2F08Nmsux1UHhtsptIm1
q+Rga/2Wy+PcVue+9+zkYsqyjW5F0NEB2Ys1fA0ArO7crgQDDdhySRvDREvhR2OX
jDHxtJ/vUrOzWOdL9qUJ9tBDSry0Q6q+ROqfW8hfktc8rP4jWhBrEktmk3O/GSAN
iLvrl276y33VzGMv0MJbD6JwNjwTCY8DZLdZVfrasvZZ1s5Pah9SNGmbIqDx/Mdl
3Ec+zNyxAOO1fJwE7ODOLJUL3hY74OVW+9fuyrEzeAAk4sqYYrzhY+py03y+JBtO
VzCqe4jV9BiNDpB9sMxNRGfN1J4cS/jfvTWMnW1tnxriQv8+baQk5Cvd78sMxPNm
s4No3W8zJA2YpEJsbEsB/AOJ6STB2EFwYatewZQo7nmLP1nFVWJxx3baW9TMUPzq
zzJv1cXizioon67n540ITicOhYojeLmuy/nKdgO11wEwnUx07ioTVDAQzkHIeZYR
BR8XBp0CVN7MDLwOQDOHajK1VWNVqFIMmy3ZCxkDI/azwK29Cb71bQCUAon1ZqT4
B4B7I4WTCiGRFnJtNAAxqWMcjcIl9xSGV7/VP/OE5cwPGFQAhDFQMNQML3ddV6Cr
nC+11S8FcC0sjl6cSl2aTSgY5lJHgHqajTZjP+/QqKCylAKsDypK3oqcdP854o+Y
5aK42XRh2EcvQSw0MfIQvjHJI/+JQoM/nsd2DAuqdclC9u6wnNoHQBA+9iTilDHI
LFanu66jlWFeCuPnKDxW+wlxw4zVJeSSDznlCSUedErvtWt/6G7dcJ9AtX385J4S
`protect END_PROTECTED
