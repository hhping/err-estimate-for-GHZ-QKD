`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wjxmxo9aKIxsFyQtz6UWXvOFw9jldrT2z+H6pjGkZA96e8lgxkEO6B2OOfFSskUj
Ks/JJNvgGYf0k/vyVuUkjk/+gAUzI4FDLUcGnFXbgvidyKcfBwnBciYcBYf1/q7M
6HF39t2lRDgvSzqxkpUfvFgB2/mo6vNujW8qOEvdsqealT8a852aR+kuIga+gnIe
Fov8egUSfddRMZ3epJgAnL2Gp7nhGDc3VkBUjtFsoAlVScjbZdSmKbo+VgifpQIg
bKAV0IdOzniVCCqmEECdKJghFf0WMtn9PxuDQqaREkGR1Q6WtvUY90F0CIoWq+DU
PSiwAktRPFBgrc8H5VIX/iLL3nqQIXIXM1a8HLCSePqD27zlXmnl5Hxj7TPmNlUM
9st/hYyaVkb+JyBag6VyABTlTk9CeyXfpg7iSs2apLgg+bqhws4MHdJZEMsblkrX
fi3ekoT8LR6vWmIArSc98zXBAHOqw8IUV2Ip/yrTPs/Pj52XI/cYCdwwvzfVDwJQ
nTZh9Qb/v7OAh1Ng5M7q+KLjNLfXSgoTVLmuk8xVOlt7tMdsKszu3TBHhd8qsGHz
W1Z4AkIPEUO3jphkYtmcKgb/yva7ucDNM2KDfzLLNmtUpZsoGdig8jTa6mMd0RyV
XwiTsJQ87R4OfTH1ZeG1br9P9zb1sxjqXVTepc3cG8Uf3EhPacFfktCdmXrKDJYZ
ym5eUcMLV7kSZ93wslByjC9zinHQ2c0uFp/hm1ZqxIqA/YycIGzkM4DRgmKEZlqe
oE5AfwgkkRfgc+Y2voAHaQ9HznxLn8YHfuRs3So0YoVP6cf5dN51X0FutjTsK3rb
JKFkupIswnnfBX9I9BLBpQ2tCOw89GnuJ9COl4ODs6Oq3N/+ySfCxCst1xDuf+k4
MFmyz/EShF/MgzxFOZcRin6f7wfByJ8X7HLrGZY/YTpGSw6XOhg2hvJZMc3ymt6h
o54WUpSntd1/s/S0WQQICpUNS8VOsFjrP3qhM3OIaSVUN2vLkriFG6D82OBUTcqN
GnYgt9IpZqzSAc/7oQAe7L/wpWHMcDDc6TSmBD8BiZIBZskbB+Di7+6LNWb5rUcb
xqEMm+zM3angkzi3yQSxYP5pICs6RUx+vCxIidN4H88=
`protect END_PROTECTED
