`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hkkplh/+D76vmYNC3ntiBO/c2dKb2Tdxg/kU9OxS26DsgMBdG8XuOZR1MwBdTFef
BqWbVfmMMCDiCSiyAblfu76qm9bKtFs+Q+zbHmwFvc2rw8Kx2NGgjbgbMxIogqml
dTvrqRCE9UrMK0XbDkPkQ/EWQlbifVXEFgjQ9KmYGRiYeotWBPV/LmAFgTN/htB5
+jsw5UFprJgY+GqZ1BYje4fE9lyT2Ztaxw12YDKEyFLTrWBSoyXMxIvf20ZRIAFO
wPKEhlhkj7hSaeWfWZMG+PDgKSmOxShBUG2bDQNd/86OKwqy8jElbHaXS/ao1FJk
gNwA7np8grXbtyysDAsBf0RkkP8TTCq+vx+CD4X0iCX4cUPriOB/vXCuKHYMd3tq
AP0Iv6KgMePAmKZYr5Gau5W0+ND66ArCfdDqWrEBkbMPeVPlKbge1i3bB2vL8Hl/
oJrt1qz2dtdIijObNgB7I+DxjU2xPL0cAkYC2xIdGDrL4OpHUQvCcWj2Q0wK4t9V
0MdTFg7e73xNTuo3wNePNgQDATYOoqesTjBZrNtiEtH9WwoLD04OEtJC9by+s8yU
+zUeAsOK+6zE8VbgFrmjB6B0bnJIzGRoPyPNO1t3Fdj4OaUWei1LyFzqlYPNbFCl
/Vqo8Ari42aJ01hVBZsHx+1hErRe/M400L5FO+0DaPUwbSkJPxaevthVSGp2xhN7
p6KaLINe8aLOtIOzcBdJJdLPdjbGCKFn3tTb6nLl+mw7QN7E1BbSpVyt2gts3Q3v
aVIVQZvTNkUTJWPnbdSafg2VJaJIa9GhnEGmmYcWS5oZJhPL9x0hcIVIr9MAC9l9
0GiXv1bXrp99jyV2qr5tZzChi/KA7sbfHWYHqyIHxBtwPc4gTFSksX07NJx7ILte
mSSgq/DTK2lZ0xZp+v7CNX1O1oDSeY2L0g+jeXQkrezjgKep+dWoFeOA7UcxSzEf
nrhI0LNPQWyWQLDJzFNmEbGOKpRcuRNDbeDbo8ojqh1SrO9XUFSBL1NBLjiFlpei
tTgYh0dNYBu2qRPUR7RJvzkoxONs7//xv50CdBAdGFl8fDQBGskwg+uI61UOAToX
1xIVqMi9EyDSGv02cTgh84ozpCBgUAqp99M/LWtQ9LVEC9mpNp1UH5Kl9ns8EskK
6QGg4zheNDtuY4PbK9ZtzVJyjTqrLLglhWfF5NvLVAPPcgy09i2R5ArIkbjIIJJT
bsVaSqR9GSfjdjTtZo62+mCyF6S7964CV7nGJnM3Na7rTI4B9CPMw2FlWpZe2v7Y
e48B2pexeE0+RnqRG+Pv79onKsFpqdCQVsENqypc1H+z28OyMaSniBKwVEeerqOQ
maPfxDnFyolUDtqfXwyDefObyOq9TZMUUp43vRpsOA3wfBtkcENhmhEmavUq2KZz
ukuJzOOGo241DOtZRzskt+IETIJk65C3e97Wm4GYrpRZgsGgfXN1OGrwkwWtvbd9
dAM83d2LJn5CF5D2zOL5wNOzceP5h1L93aLihAaUBVYzvX7ie+9MnWpzCZNY6pKz
IlyxKP54gkG0CAiugp3Yn1JfUdDy1Su7sLqIRV8CKlQXDk/3Xe/MxUFvYVJdS3cd
`protect END_PROTECTED
