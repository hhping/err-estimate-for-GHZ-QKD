`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RUHtDlNy2j9q+8SlJWdkQOGgJsvxgsvV6vn+YaBn0RZ0o2n+YD5YYl//VUTlRZUQ
Prw0hc+VB23Fdi69gLf3pknqZxXcYgqYyxo42bij1rRTtl+PH3WND2geyR70TQne
20jIo6ajFl/i5Oqk2ZeVxNLb/Ik5oaVL2ScOdm+xS3D3qwdVYSGQVW7XRo9QEJ8T
qFdnuK6vqzeb16E5XP5qbfUcAkMqs67bv81gkCukVk2Y4UPkOjTEAeXcIAuNFn/z
uMHEhMXz50MIcb1LefEG6J9tICLBFC776KcehwAiw/9bq/JUxFOq8FaLq7b4AZnv
kMYHu+q/w76d3Z/e/FS9uYZYrACdppwHJSQ5Uh7QOTvwXRzjGOVCVomggJATD+0X
Ww9fvmzQE2velejgJlBHN+rcNGJbWAPQuJtCTZa+ffxy/xTagbqPAChGZCrd4hsq
sfmwOgJQbiI8uk6lqQVqWvgGjjp3yqoTK6Em9oPFX5iZAy22lP2TYJSCSP7jpPdz
NtwJ2VA0VOI5vNc8/x8H7lLAGIvMLNZaYvaJyVITZjvbuQa5ORgROvwBM2sdzuVt
`protect END_PROTECTED
