`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tX7QKcn2ss1HmsuaztpWepjlt8aIofpgFmoYNPzeFP7dU9MgCxpZIhaqIHOgAtwc
/1kvNF0Ow9RWp05xb5JRk7sJnrSA9VMDGeZkMXzzIoUmYh1d+04dVUK2xNngot+8
lXHh0K5g8142m+sZ2qv3NN6LI0WVGIo5879yRNdieiCJCaq+prTMchPpqA3mQkH/
TUXJFGGAnWYrBr1TAOJFbfKzYTwOf4Rrd6MvAy1EdNoRs5Vu8FaxD4m6vPE/Esew
UQxPuq1k+dba0MFHKSoWy4uZynWYAIr7oShr7z63HBSKur76Lel2aMTslbBU0kbo
sXC1j2YOQSNA+GZnNcsMiERGSEuzR2Erdavnq19GHUNglMpetSt7zJSV289F+H42
a2nVzb+ttTF44+tZsLK5MK8LgD736n07yAr/9wBo4KOqbHV9+4+8jkUJdnvxXdM8
aVUNQSKBC52V6H48bxpqzbhbFnSh9HJPmHlNBd+FyM9x6F5NEJiWXR68bO2pZps9
4wYRdm6Li8xbzm9VfDoIcf1whprh2YuH5cDRJnQdeB6b6JHA84YNLdGVLCs6B6Bp
1n0GABtS6aQjJcJ0iuONNlsQ4a3jxeNwHsFP+t4YPGNbv1dj9YSzABqyB6bKEdsL
YjMnK+y52WfQF4pdu64ADIfMlqbOT7yH1CDV+sMpJ7pPXzLGwbrRf2craA6YzaPS
5UOM2INJSQDanZzbBhx8sL+JbZTS1IQpKda7awIwl4bchkFEq2gn0XmSXFMnM2iI
LjUOmVbYmZ3qO905vEI7nOKWbmZYCxPRoy1JwrOuvbZLs2UIO2FwjbiWk2rM2n+e
JSLxeVfd+CaBXWpUjQfiiIP1QuDQojsbhz+KodMEufXHmspQv/wg7pXlXBZyEU6i
XUZBRLaSe6Z3ck4Vy3Bn+OE+NVU5MmraXsDaYt8p9nftqIti165EbbwPi6st8QpP
tp0dF0ezVwt1pS7IMHspX4bO0JSz0hrQeMiJFk4M61XshgJyghewgyp1z3kx+f9+
t+0P9hy3+LkuO/Bixb+Flh2R6ilSNYMpJdprYOcXPCJqlk8bOwHcLf5AnMBvr6aj
zr+j+2wZeDVliR5t3yBAgZcyB79KrdzeGM6fuK7IojIqp2toZ2hFQgplADZhNvov
UPXKT/3ya6MP22jgaduK3+sK9BQdL+V99+ySmBQ4eF7++Cmonj6mtNDVkbRL11az
dF5avZNDoS5nX9VfmyFk3FfjfFSgeQnpv1W6VMCaFTHUHT95yhbmivoFiJ9NVtVg
ykR+TmrIjSkbNtLgGINzU3YV08CqGhosYQXp74pcGxSCK1H9rhG0UN4JcXUn5A7f
XmpluvLQIM8vGOCNE9qlFspdRS3bqwtD/ZyoW2ETBexHMXPLHG167MjluxYUt4sq
2kDTRmr8p0ApZiClP/E4lShzNfapucWJlvZVNgVk1k2WEJqNFAYWP5r8GJz6wHFy
0BECFuuOk/I47iiG2p7GlZYIHT0Ep65oFq3j87v2V4GWtikiEmViXDqve8j2lpxx
0WxPKUb+076T+kTl4i8xjHqhlxZWKi3hZx4FyBxllDhdUUvv9uZbnPFVOI3rptPm
QsQaMahqk4DnpSGwiRRX/dHbyychx2sCOJzdVRSKIIF3Ww2Ve4xyI1crZqOcsfik
WrH840Ywwfvh5ss+UIW3RozfCS70PLlzgD2O9r6A2ruAJ/tmn6d21u4zlqJQthdt
36rijzDRRfH7pWQ0x3SlN94Kx9A0lN1Dk2mEsktVhGV+RB3w+kcJDIWwnpJ5GGPB
lL0Wiqh7n6fRew/UyBytQbQIlQwitGLu4PVN7DcQCyo2qa91BtA9WEc6gI7KG9bj
uYK/NrJ43wQnOMXpaoF1zUujB5ikXcxh1EGFN5E0hwbaPnW6DZZVMGlnLXl26SzY
eyhpbilEJYchQyL9/aggsA==
`protect END_PROTECTED
