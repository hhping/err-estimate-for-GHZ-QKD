`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JsQ7F3B4xGnS4DK5JAoiHeTJ5t3jdgdq8JnpTj7Ss3NHjaJDKSRFgcqg/G5sSSor
m6yalYAFnMcXDMefjDLNAs/aVQZaLA12Du6XCmgW+4BhxA8HijkDHc3beDox7gPv
nku7lDtMLlQpIC8jrzGzl3zAVQvbq8I6dvVXmu6GdZuF8U3xP0PXGVTvICpi/vw+
UpZGmk2MBuUU0AhZAkhYA30zmiTxuJc5iP0VDRKrP5AMyHUxJjxezDO/8CvzXg9f
vLrRHidH5sGq2E4DYRr1fFJoxUMB8KoC7xVSwaJ5kEBzsQ2N4yBy4gtX6AAiWmpc
GxkfIOfQqAmLXMaitYNRxKkbZa0teH4Ihe0in6U97EtQAk2tcGtgG89hsFBRTOWa
roQ9ko2yHBvl9yOf2UjLcqrYKcmC1TyswoxVuFbei3xwCFns9bY32fNSTqjmKji/
m2I/b/WUS145IUhQtLMzToIM02ADFRlXLd2sihTbuAHcxdTjNuVt+HuiX/qw+EBt
CzUX6pEQ3228P4cfUM62x2sTnVtkhsNJoxZnGqnvrhGi13bicbQ7Gm6ziFydCDiS
V62PbRoik9q+2J0S5LYtRqD5QOAlUNSNUtesgJ6VktoA46yZ0+alDHOXKX6zoxsc
mizyoxT2dvzh12fJwE38Yhe3Z/jF4urE92X3vWXgKI56qKJ1DW0ZUQ1D/mSxfIiH
K7LC0YpFJ8bCpl0COP9ehIYiQHGERIwkJhJUalG2E9+GpIlXSGio83x9V3bGUl7S
p0q5AFq307STrimVR+3Ze2eW3ZkrJWomt4SxKECunmGLImVRh789KfXPpPdXvHsM
+HNGE0CkgfECRq185tC9ApHOpWDDFGBPjw9n3NVR/FtYaYlaFSqpIxnCyoHBL0Bj
qEF8q29TAg2Tidk+w4SV2albe8j93h3PPvwKg5MR+b98QSTlm/evOMCA8pJvyT4m
eUG9Jrk4Cjuc1u04XMlDkgp1MWec/e73nAorpZcdMrxSWJP8xViEkZnOGYdroq4A
yl6tXn3PvsNvNkueOrHMnRVWcE/b6E1Aue+udvTIpOW88WOB1s8GCjFEF3kxO5n6
44V4Io+UbKyTJbMRSgBxipdGpGnHPIrsLAWQc1nrN8O1vZ4fCHEpwLbLZ4iZlVy7
CzQ2T4kRIpNAbpr6Kz5kbP5R6lQihOpb2MyIOCiit+HYC6OALBulFGT8q5NT6cYL
wXkoH4rYWcfgwYNHiIHNkL7tqlV1z2Tcxjnf7dhwOPu9ESBcxJdFWR1jwoCWZlUx
OBE5mfN0kC/+tPaABpOToRRMOQho/GGnNgtH5m1GxvGsE37Oa8ve7adup3KGLHNC
fluWdAgBvqm2TQqD2KMvx7hVZqwi3JQuwB1P9oSJ4MteYVNpDuohKmyzpLBhEDHb
kPryed6nY+Gm8iRfv0483tIF4pUZHtr0PWu3AY72d1OhNlL/u+2P+F2XC4X7Gmwl
BTvOs/KhbiH+/ZQxcciLN2RTEzLnFDmyq1T0E4KH5WXQUgXQWghPQa/BwIbbY8xK
z+WQj/joPWp51jJLCHPPqtB6uwTYtZ6JzYnqs0Q1KFS6dwxtPMULNphs412K0+Kd
K3G8kfxyhMLO7I6WLd0lp7Pyhgf2vP6dV/hcpl23MZiXohZtxAN3TkTY8UbS6Z1W
45TMFchq/zyIoOZRjV9GTpaut4LJ1HQGEFxoUsYIctdAfXSIMRIapvJP9RjvJ0YM
UistOZfPpEFnGvlvOLRBXJ3nLXRoclQcqSqj1sijQeJfhQ/pVlrcu8d79FsWYDo6
pIA/TStNiC4d30j1Qsrx0VvPCLFRDiShsN9AatPYg8PY/MZV/TqVFC0oKGNo3Rp6
/lzgpy2yDAOG09Y25NmeVMhiBlEUCgCCN3ArNbiIx56TYXDWvKYfE6KUAwnjpKnI
Pdmt+iB+kCG0ptimPFMBiqvymmxTw69w9776DZq+mM1vagEBW3JfOnSJMc9n3Gvc
clss18HssTczmK6PsyQ4LmD7JcyU33PeEzTfdZU9jryldO6kdWW7tYzm99iyuZ4C
BrqhfthAfXj1rTwR7ucBf2u5ACy+B6ZuEQOsd9FyTJVbrYvZYzsI1KN+LDTNSOit
7YmaXSAyvRgJdLWNGJzpzKoSR3URZAWQBGHeE3qFlvnzwTAjuxzI1X6AAVKuoQlx
hberAATDko2dUqbX4nYaWtgvBjaP2G1gTzAYzybIWE1Gvp48rEQR9yzyIWgpKbh9
2KW+4lUw8XZmo3VjYZxK0iX0CcM0Errq3Dj0JVj1WtHonOO7yjTFQ/eqx1MPDZqs
+UXhH2yZKvVD3/abGBFrgVfVrIJ9tIxU5I6iigM7hpe3/siJNVyNffL1QVVoUS4O
xCGD5Q4remHKYrFxTha3qUhUtIodf9sy7Itvh1R6vy65Fu9UK26ccNOWCUkm8JO9
Mqed8CIiVR04GGfC+smP3GDhHOsfZQOE2IzIu3lwAJAtH2/X2K5buSoEjwN2ndmY
c9mOwnt9ZvgDVIaL9JsiBh8pReync8ejrmyokvfKEDh1mtOOYC/9JTFxZqZr6H32
YHZhAgn1kimLkkE5im1Zsa9urkLRrsCO/7VD1QGIJ6MeBuy0wTit3QoLVYUyuDRm
OiUNPBwd9PK4G4HXT/mtM7ty4FY1yDQy4NwUfNGEK6BKFgcGxnOUsS84Yot7sIxb
53DiYqfBy2GE1lQan1l+NYeUIqRJYOD8P1XTJPt9mj02M2mDZ5nLtMTUEdoAPobc
UzG4BNoLuAPyv7h/1A7tH1y87LxM5JimEIQOZNu86yMSCYdVmThdQCSbadf39zZw
+2ZwyK8CbVM8fL1xtUJ1OiJrIp6jinP67GEhhANEwFHSOUgQ4KJxmkYzp/5MLzjB
mWR0DuHH+vAnDlwkh8SgwimooMC0OurWh/Ecffx+FE/zLni14gVPAR0cPn9uaMUf
skWTiuhKhklylUxUOHx/djQrTzKT6auDdu5+Me3aboI=
`protect END_PROTECTED
