`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PVN6F1vBF0BawyPF0poGsM4jm/F870ycmihtgoEQwg1RzLwE34Xtt+bMIQ+t2/NI
mRe16IQAyAO0W8EvMoj6H9tBcACEap3zbGVUJC4zOVVpv1FLt1v6HFgYbeNPLJmQ
g6zlEFljhGVxlXP7lnpA7KgqRivFGunuju3Q578j7yT0Yq1oKXcxgI0BMA9z8hqi
rjgy0kzZY24mbWHrXzVLZKETNQMkKR4/EcPSH13PpnQYg72uZIYpD6lyk9xwLELZ
tQq1UHsAF+f+qMNECb+hFjTzUPVfhk6LpZOSQaEzvZpWtqXEnHqCmb0NjJFEP+dK
8yYtuQoDHUQ2zDC9IGjDtLcqGDaDkT26CkYMRGjV56jRPaIbHFC9/0fYYZdprDwy
nMvrdg6Q/R0UHe2E3hTJ2PYw9FP1s8E+SeGebs6VW2zwBf2BlNWFxiBn4zkOlL1+
njP7v/+zOPgieSfYK44r1ykG93q2ioG2YaqbCHHlQr2YWa3fa8QnYd7YUnNbPwE0
ttyZFlmzqFKGukwhDNmulVd4/SPJ2loyVoWuiUz8dY+9QkroXM2Tn2vhqFnAQppj
JEkEfqyzA9YxSPxGYr7UqQw2G12kcvJBa/Y98v5pleJP3uoEpOIWofpRlEsJvhWx
saOdS4wjDaipQcYbKHZ5jhSFC0RlASwpGLDOoLPLFkqvxgKoi818qtYyNo5PJXrD
lh5nBOv3gxVUziUhKvf4R0aBHKWI+VfToFQce4Ogfgwdjf2FYvzFDFQhWBSrPY4d
ZVflKS5lLtFOSZNZV2wfo9GxLx5+H5xYmvheDL/HRM48AiuBNB7q2F94xDMBhvPT
tSZGgYKilFYOnyJ23bWPIHDm7KzzCfmcltKh20zw89g5yjvFypLHKpEV3dfLA76Q
X0YDcOG2si7z6K1vpG3yA+acF4sSwLM+Yip95lIUnCNQdHx8QbpZ5e5zM1ej2Kks
/r3gF9M2bBRTah0++wCHhTdtsvn5seIhl6jYWoR/gLsrE4IL1e3IAfgtv0+kFfSl
SfaLWKA6BkGDud6xtmH8oskrjXNLFgQgJAk3jP4sQmU7kMKQN7w9XtL1Ai2sp8HU
xirhSu+/wbY3ecqCSF7SjCYp99dW0fk0B4d+ymLL63SrI2LLY1qF4Q5zfE7HdOWr
pzZi0wbKG38vmQtvYy5SduAGIHqycO6MUfYUVzZbPpmIXPSXmjwqDoF0tUXP1AXV
leP1t/i3tceleZXQM5jJJukMKjfqq9wB7EF8B7uWXjHCJn0NsBrJhPq0hvNvSVrj
vNu9VamdIFjf5z9tRHJVtew9AdeW8Df3BPhjDurdqupcdMhMM6M2FvhQVwvVnBWK
qJTG16ilNEoK7ukftH2EGSVv/DmVW1VhbbOzT3FH7HPU6K8VZkJSEmlIZ4kJ3Zyl
fyJkCTTQGRXkEtjsSIQZzN8OJPt7XrQOw7Cf9/KYDBe1a/EzX4EY4rrucn0o/3fP
JrkNSEB2up8L7NQ2fNYbtHYKCFQ6dORZ5IxEBZnsu+9EZA/56Ml0FXa4NJdHtXBQ
609G99cZ4AtSxGS2w4dO+kQKBIDVUunOldqmkWNvzS8BfAYpzCmKVH65ODJltPfO
tjsYPlhJRvipzcXcYWDF5bqBtUJiiOWpISRVFJd9dx3bf+N2Cdkk5Ki68JU6OE9I
dfBZTbnD0HHHHoI9Sp1Y6OQDECtIlzlPd/xd9k4VcfQrOlfSJhFqSoOt861+e3HX
3YZ8T2b2GC/prRCiAXNoRyW0/xa6ZPePnm2wLVVewgdsoExgA9X1CNZxuVDlOeMn
NTWE+nk+CvifTNS8m6IBgoalpoWduz9QnOcmv5DwCt+Uo0upS0M6XQw/b/9+9BAZ
zx1PJJGj+mayidqTDkyslh5CGzIqthbTRGcjgLjDb06Rt6xrMD9bH+TsOjLpqznW
juJpfF2NV1IPtZQLCrX1tfa8WWc6nexwj5oieqQwcZFRDCs5xJMB92a4QprBqNW0
llsTt2xjWOhh1mZo+pQT55g4+go0ij350JWeVKQ0Vm0EIMZDfZIdPd3RkzR6qg0H
nErIfhnNTv++voDw559Lz/dP5yqk/Ji7ZMcF5OjZSmX6jwDuJTOShejwz/UI7ZNw
eKUAVO2qmE5UVL2SqZZ4jWE3PJnZScUCQwyvfh/KCRm/Mmv7YF8Ir1PiDdIIynpF
lndoKhsp7ntlJToJAnMLa/79rm7t50XDBiMuJoqVbAoSHQWmoaTfiUWcQ7S1uK8m
+hESH0pqM08/3AKa8GuAXX0I0X0BZDpz/NY0hB3+RQfUBkVAkR7abhPp0+OMwQff
SOV6reMOZNuqDUAlMKmhrxpwjVSZYwx5T6CZkZ74QdpfVTHAmNZk4WjX4m+OwAyw
DYyzYYoCKAaia7DEjmbL8Gc8Q0qfeb7kA/B8rXgFuISI9gexSt55m+9RTi8bjgdH
geaFJrG/pfECjXIHONtWZFsNusQJW5O26xRaGDqqKTSGQo1MaTcJ7W3gAuGmMpf8
Nl8Bk0CDzXpmZcrLwfJrfPyQASnO9OAW07OFYKkX6I6zkiuArg5yKpErXCQL7MxA
DYndj4JdDxbQUHOIvK0TxjbeF6FyZbsqPIx+RAdyEFzvccCdnshKKRh5a1aZU2dl
CwGS131dbETLnTxbrJxQhvepqdcrr8BCzCAtLDOSSOAcso2youp+fiTMS0OS2YUA
IcmjBNZcPsAe9VJ6TB38mxRUHg7k8y/u35CP7jdaeewya6437YBJxf58ggurEfMm
DcYPvDHA/vDYRKFBrd3X8yFYl/fK6s/MFajwkSy1EcrVfA2YdDcXVpUGOA4P7HWw
qezWvFpATJaJaU3E9GVJKw/3hZx4l5aUJfzBHm3zaWw2mnYaSHSdzhvDO/4pyMOF
geeAfHomnqjy9d8YNVYtOW6U6yO7X1jOVxpQJ3VZRepBH3sDKPGqvEkk4yKlcX1R
BCCUIJp/EPSQi981/EvnTeQEVPNl6lZ/v5jXqpu+Afk=
`protect END_PROTECTED
