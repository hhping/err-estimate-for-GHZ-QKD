`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nVcPrpePUJdf5QUCLaEK7Ml6V0IdmiP6q8nGGYVndZsVd1+LJX5vKXfL5kwfROZR
zgemnr6x3Gw7IMkqHZA+wjQY84JcmwN3cIKhOkI5DpnKjCNq/RjwjEZb60isZNxR
cwyEhcG1kQtkxujoN3CCtulytKfnIsmmfMR71PAE1IHqWszFKxqbcxaV9zkjR5ox
CIscGM78/XMVQ+B3bIBPD5MjbDk9P6L0TbFY0cGEt3vDDI3UHCIkI1sTNBFvpP52
Dfi4M2mMNhPP/5DvCeLHcu3cAeuR7Hc5pK+LO/K6bpikt1GylNB4KhWHhgy/SunX
9uZVkDPujEhntBoF+RXqyyWbb/2nmIa1T+JZCMdswVTC5DazW2V91aQidHE79Jtn
CffCpjjy3iq67eBDI9oYBv5uTXSJXQfwKlkfRLsKpDYJW2Szjilux5nJPi2KQ6ci
FGmvJzEn5iz0vAeneVyf1jCHS+EmP7qOioIQ2UEYi45dTzEBM0dn4ZHUXiXrmmeq
uz8C7Eocs9/WifZ1ijIr/ubzpf9b8gplYzILN+FFLzdg4+CfMggE7RVhJdh4C0+C
0xdAwdFI43EEfHAo59piOCjWfijcGBfdF+rB61lU9ByKwAz+iiSpuSCNr0oxF3Cc
rHQ5JY7bHYK2hK+7sgqavn4ib2wTlmgqPowatcD4oLn8jgx6uuqTFcOKyH4NFW5y
u5BtavSiGKWz9dcCInSaIGrjvKsqxkXpOjsmUJqroEl6qg0JVuqP00RMipQ9CXxG
kJgb/RjI7yfCvORrsc2q1tp8AFz0SJU9ZhNVmIPmBgXmECjAvsEzBUzGwEcPSMZh
V/MGA9b4nItgyFckQaccaaB8w1tzOM7FXCYPzCNqD2ESPHOSemefQG0o0pRYhkrk
+oUWKC/L52yYxaBV/Uq/WvC6p8S40NK+y+dS1a+yJuwuWY2/QZ3tSwlPFI382GER
4dU4RjcwnLh8xrvp8PhFUJOit+v8yTAxirualzU/OQHUWO/f/gtSHMotOrIBB/3Y
T9s9BzlvU0pGmifli4mUxx/CewMsZBodDB14hkHc6XrnkjkE3UxzI6fkUyZiFeW6
tevxET/aAEBX6THw5j6lPo3ekHI92Gtz+EwDFQbu9F+W/tWaX/A9bBgxCyRCDbUD
U0bw8+RstJFBIqoOohtl5+no8umMG3HBIToTxijC9fVs8Y6QlQCWP/fNjtdsKk1A
0Sii/S9l0cPQ+aNPxOTUiWrYA3CA6Y4lu14vYgFtvVY/YQH+gYlC2cPLeZhCFo7X
72tpN1h7+qjCP2xjZnGQRyFQXIawdx2+5EOJ3tnaPV1c9TtFBBN5X7J9bxfK38A6
F42qJmmcXbhBKuBtizEeA4qPd/X+T5pYVkcA2tHNfukcdFkb3pdmF1MS/BvI6BEZ
yd13QukDefg0Kn4p0qS43gztgwYs8W+TDPQSmsulwiPSBNYj5B4txQU+5pp6whg/
h5u7GfhZ4YhtBWaDqxI1Y6xf1RSc241kzjsrUXcYjGir/3TfyoCF1g1IIfbAsvSf
iyQSJTcr2+pnB7oUDC/ZZP52kK7x/kEccCnEp6Yja/B9z0yVapIZAz4hIvy3rnt7
zkR3tjBrCVyFOS2SCh9SkEwSOxBVWiU9hkJ76/e5soJZMHN+wzAdn5j7T74upn7J
/GPa+2IqBoED+hn27FqayQyoTjU2bTt68P5oHBg1DAiWqIU3L1z+jjNYtEWM9AZJ
Un3IZKhr8vfW7o3+lAZTdyudLT4EAuQWzLD6ZXuf3eafXx2KfI/qZ8Q+HOeusgjK
jPTkZHMIRSZO6HYpBc3IL1vGOniFOHGJ4WRCbTMNTaROWuIF14bwDah2IErjByqD
zH+OwM3FGg9LOy5sytyySX0tC3H7Huwkrm5ce09URB/pyWHzKAdeCV68WQio+V+E
2IBD6IGxMOnFBstXAwm12EglpPt6d/YhiRNWY2HVDn9pV2pVRvOozp7htXW0ZqP7
vXVKdPPmVtC6qa+Wcp6yWstmpzoxJt/+lKu96H+vxATWlr7u4Ql5TP/Y8v/LzDo2
9u6uLeNwulzrD3rPpRelKA50SKUgdGh0z+iiZjVg+GXI+42+zEHVRPjDvg4JZHhd
GSXClOiFyVAJwHylDl118aRahzxWI0QwNna+wr55yAfLhHIzEQU0i6hcfjz5UNmY
FSoaatMQwJT+Kf7BShdz4W1pCQq3688GC8qOa/JKJCo5ZlqEo2mvCaJQinbS9MOJ
aJ2zY7mg3AzlpxoZfbEh4JIjpXDkV4gLNYQrnptLTUJNbU26nGNXo8eWJByv28av
FuVIwecimjYbsyCH67NpvUprWmSn27wkIjY/IZ8V8k+r0iF4jZD2ygNi0vauout1
BQH0Cw19p3BHxA7XKWxe/INSppjMVSVHR2DhM4iCVHRut5182XaWE1/ZD7IhQCIM
2owL57LOzjZuLLBJeIwjWTXkI6LFPxYoVmf//BwuuDnyFHFv/Z/Jh8Z5Q1CiBpwI
hbrw/GH4QQXWg/P8sSTrveD7wRXOmdDQ02HMYd9jih1w9yAhEtYH+Qd4q7W1zrAi
u8TG8FcKxRtUKLD+R0DdPR62MqydCJ+N/6AzpRqvmpCuLHqiZVGSiDt5/m+VNEj7
wNbncvlYY3uhGAaegWYOPwgueHN0Kmhh3Ztyhi40W4wY4hWGgqCVF1HZlR0Rd2sH
xWwI5M1EAsS2nTRbM/LATi5Y6FVRl0CcyfQpFExV1HEbxbwCXK7MicJochOJQqx5
EIp63HKYwy7CotK5NVzPpjGYaWs7mdO+iWIzfgZtpqDcuTpDPCdoF0zVfTFufjy/
tVwQOywlDbU0/1o+lIqOBHdTDU7BXOv81hECEpq8ZSgOjX/HhUIWxrSrFnBm8f9K
2GuqD9dgKm8DpTJyqOXc6ixiZlLnorn+ohLyyzhVQjm9dGA2HvK+DZx6tS39WYyg
pVJOW3DTfVcuEKMqSw+DnpkgBpAiY8ECKJWKueF7eG1kbDGJsAHWjsZEvfjGiocG
w1aT0hKWMs/Sj6uiJFGlg1Ry9SFxl4qX8bXedRk1As6kCCmGlp8blVYkFGt8aXyp
kKQOycnXmiyJnWzouvipFVu7P3+giMmfW0CsAwCoWYGGHktR7YV3roonuvDB1koM
Iv5KLW2wG+TQfkpZUJXcXdCwa0SJOWrtLvVo5XHmknJ9M7YA6J/0vHnwV/Uz+nxz
3DxOvS83bIKgatKGMJ2bYlgNY0f0+2BtmTSJ6zNtBu+GoB+nI2dyLStxk4qJ6991
jHSBdHcAx3V0yArgKdER4aQ+rnYklvAOxAod4EkiG1ZCry6izzMxxzhYYuarvRYh
BOwQSUDK4udX81StKhFJjflNW6cp2IabFWvNzbCVChOWAyzY+A7/2+2W9AtLvlJX
6BVU83YivLPLAu2DXbDxNiCTNQLdyf7y1DWZVFLFTkPcJ3sVqIFdhOZc88I02tDq
X0ev+LAu7Xt20nzFkdWsbwcZiXVYimxOgfqA70yG4BRd7OUmCj5XfHV07IAxCDEF
KWkoIHQvLI8s7UfDLWVNN1KDsIVnAdOMVUiTb9oARmhBFopJNeMCnR0qaPnhNj7+
SYjFus8dyHxC0brQLmFAzuFlp5kGnNFjCbZHv/FNsdbuSEShstuUhbxR7N2gEolT
cbD2hnpwv5cl+0N5HMmLZo7LZ7GJ8vmOJhmHpyAnwUOPV+a+yTP9rlUll1nWe3b+
DZ5jXbGKnz/RAI8k0YFEOzzwslvftydkreSG4CtLrq/RrBWL3qKA9bCI7j+Vl50U
vf1TA1EymSAkkk3TP3jYlKn96uFHZEMW5g7K7md+WlxKUdfsRtFxZCdQ7MU9JuBg
7asj0Vo48CzHBO7lQ4Gdsu/TveeXD0Xyv9RUCiitcV080gcyBV8yPoouAmyMkbi8
KIpZPY+b2W2bop8GMW3/sVQhQwvHVEcW4A6WDPmCVkwU5dhC6F23SZKsSXhMabOD
4DZdplsNp6qOjEq3Oo57mxv+bovxpItuC1yiENhD8s/zfj62N2xD6KV5m6qYicLS
NVpLEeOPwn7X0v2ImQoesRU0LV4UssJcPA0fJzRy2UNxRHVVNZAe1evHkhx/r1HH
SZQL9/S6PkN1Sxo0WbF12jruOs4f/nkOlcLpkXTHUDmjr895DYbCsXsABtnV3jJP
wuNhlrzCYt46XHMvvelOqWEoN1yLtCG4nfm+dfPx8b7ibidY0hsVj3MzOm7gPcy1
7FHSGSxW070FL1XtovApH2o/ZyOvCDGApPtCbwHlrfpgloUZf0H1BhcqNDilM0Bu
yi3jVGgJ5oSmh89ve3cak85Us6tS2ebK0Uywg0qqujlh5ijWVKc5CC/N90+W7Q3W
K93SGfBgrPRHlCG+hS9ykcNOZmFfFuzAQiD7efH3+7Rg2gIXAv5/rAHOTAWeTSgf
kDDddGcr2KAxltx9QDzjwWwEdWJBT+IindXx0tbKFrhqZx4xtT/pG/X5x1X0nm9Q
J5XR8p6cD6FKSt+MEddUjjMhFQtGwc7zFnPVeDXRY9iz6IpLeZMhZZm2jTfKiU+Z
BsUvKdqsKhpt33bOS+ZTAV5hayd5MIprazL4QJfJKA0GQDb5orv5BwWd76ZT3jYt
cuN6UPaVVCXbxTGThOBmDm985ltpChsqMILlIxDAW8WWgMJPCajH3QNan/bazxqr
Gznv3/V79N+QZ9ha/KLF45NRmzE58S/WUNMNyD3CXcHwxOOtQ8e7lYn8CuMwARx3
lNAtUwguPEi0mSiEiggue8OprxmGr2dD0nKJQRQdZN03wFQzWw36xQN+ImFvdNgc
oQLq2hVkvL6EC78kdYJ2EO5VbNULB6YWXZgW+QXb8JiZhmCsL+kx+wm57h8G7AJ+
Jh8rm4TRZ/rNnj4IuNOc+fbtoj+ldGrEM0Enb3Y9CIRc2TkJqQG5N/2wcPTFAvjG
CDh9Sn3AhApPpHo82mox4D8/hTFbi1GtGiZ/VJFJ+6p2sVINv+xyLQRe9pSc/bNK
URaqEA+yPrzzjqaJvFN3WFbbdx6acvwnXoiidkBmIXTev03JfrlbVX6njbbj8aWl
c0IAcojBOpuvBEc6UgG8tDaIqwJuI+6OZ2rBi3PbQLcDnUykmD8NmPiQFYh7P0fi
H3jPybwhElNViv8ZUUWnLiT5x0KMsNXG4QahRW8r+Tu+QFvgf+FSAEZ9tXWNZXCL
edU4fVU17ggamdL3c42v2KdgkEGaqWc5V7loACP/iUzHjOM5ZOmQlfTJjsSwaM6n
aS4dc1ezL+afGTbD6YQ3N5kXo5I4lAovIHim7gi4/9QOud93YbmQmSGms4EesQxK
8WeSCBRz61mMJSVHt6FCD7z6x2Y3p+Mvk4ohz5pfedUx+v+aO84X/z5ILgNbl0Ne
I2dsGYLpLtz5UE/71YV+VMpQXXwo2SCdPmc3QZLPF23+HAleoLvlxuoLL0KMFebk
yrBxAlByK2G0bgSVZDDE4h1mUdFsz7YNunw5oh1inajMB0z0SmZxXcPVIZBH0Eba
1xlfKo7PEmmvAyEf60EsOfMEbtd4sThtUzyEL4j4nPBYzkhxkX0pq1CbICqJI5vU
upGZ279kwPoJP05icZje/r2eYU6pXEmRnroymByPEKZfItBYJAXkESZoUK1qoi8g
ACNHhLhoWjddiVCM7diDGnlrVOY3942JchNbfACjPKLOjvp7jxZNm10cdBF3E1UM
p5zV1s1GwrFVxEYPGMa3tTFJaWqboVMxDZHNEEnfneWdCY6jcOxakAaemwX6a04q
B2NHblvtdfkavsS6aMUCRfmJAw4LcOn64lxnCnux68khL+UJYcb5ML1wJhegj041
83wb3wlrB6g7rSB3hfiCkrxFarqLdg0mXkUQ6O5qZcoT2GFjU6ht1s7mRSsrRMDq
HAR1D/bySys1N7udNie2hHftXlmbMX4k4vrNfNHUwRCCzXuR6uoeFY0rtiuUGewu
tQEePFf72QPMrR5FRCsoc7/FlKVeEUnewBEgFG/1pxcuOS4WE77N1KGC6pzuFOAa
X+WQeqwVgYY/FSYQYU9cneWULvnv786w9wafn9jfe10ps0ErvlPNFdXo5Z37cfT5
RSNz+nfynrko+KcDomHh/44/ViFcFLqTMsdc/MKuMGbQ8P11/HGK/0pZvP+RskHW
TMaY5GC7Swfnkghl7uT4O8S1g9bDtlO6h4PK1NFXhcGCQmpNraPoLY1usRg/QBiE
NMXixV8QM1pp1vqi1EopikhldtE4psM18U4DHGjUQprM54OhtvKyMEvLEtQsHWBm
MO2LC25k7eAmT/OtrgM0DbsY+YEBFagrEwfGAjTWc9kDSt2kUPdiJNKia63n2uvq
witbGNDjgZ6UCXksvViZWZk5P7ubLpwSaAqn9nBVmByMcbNXdtxY9BMk424hFcnn
D2JwjMJTBpe6M+gCo0D6kEiARKzfLoUbHbYkF1RUniWiZCxxe4D0MkPGTyivS3GF
ICFARv0fH//Zo9Us2XPZROGYatCm9RpdkGb7kKwCX/B3aa7btboQEnNcynOU6dt7
IpgnXj8NYIginjH63FqaIEv2ffY3B0ndAOb4gFgdQioD/MLAiwfI+qQwmMwHbgTc
T/zLX6aa/IrkLvlMUYCmiqM3OybkwLLxHsuzAWS11z7/MgUYljsSyePOiyU1Ciml
kk83P5vJRI+NtP9N0mT7Jgk7oNnk1TVC9QFpOMhq7ARO1nIMisI6yg02+Jy+yI08
NLTI4MoGPJbb/+N15VMBdlmNsiHrP3zFKrgATixJHnEcyW4CJxUMRNPsR6n2Tm2a
ubMdfE75fFMlaRjvn/0gz+WCZxnE84KpH9He2Vz1mFMIdHIxdpTQHr8r1epd+s7G
ocZ0toIuZ1kaYBkCr9bcuOu/uNsS/xlo6r45l/WyfUKa5p3oIe/wM/Ejbwg4h2TA
PO3bRhNP0Vzx6RyYATAYobV9wBeertqzIdsgadFbnP2Yop9bDmE9aup1B7rs7q/1
KN3+DcuQ+1W8eMdv5BNC2aFEMRfKdavI3nvkVns05+ZQHFJdMQE3mhhvFiqYrxju
geEtdStiol7G5tpEhttOIZwM0J3wYjE/tIFXF9J2cRHcObZskp+Kp4docS0iYrdw
uM3bRvcWWcGom9SXl2TGUfyw9+lyHp5/V1rTNZ9cprR24c6p6dFxMqN9BMIqsjuH
KtkCcpvR1xGYUBLPgkaBOD66cM3UWWPWK9el6c6y61mvwErrkL+gxKhpVmjnzr5g
rCdlqgXRtG6juBtRPZ5BrE3YW48ieeeO0KihkByvYUwOwcYAefLw4kzqp/SaJySS
bG9uJYCGJdBuLj66nve++wcpT6YJqCbJJ62nBhGeLlSVbiaUnJACvJFnFfVbA3j+
+xiPfGpCFnVBMXBntvARGSr+toTRybcALlVeM6hgpknKJi/9ddvH2opmEXTW+6VL
vkKCOpUlv/iZR1QPlhXWi+XnwY6F3Dj1Far5JrQHBJHx5E2RwcMxdvZrP8flS0HC
JMpo079m1DB1y7LnUglesa8MhTDiy5VomsezGhlTLMq794E0ZPei0fIkaAGNDCzz
tlNlLMNCIUAY02fKBG3V1MaeTzhBh0zB4jA3cLr+sc9wkE9WmB47+2nk8WVTguLq
zuCAqq1Ow0mqU3WWaa//fVk8tI4EHZaouYQ5RkcP20p9TsTJfwiNMcCxVw9gO+a6
2Xd8LKcISnoTawkFq4KvUcCpm9oq4xtvt1t59yakUxiXMi0mm4XbXtBXnV2KZHOz
WIAX512zWEM74pm0YgCPzexQ/ADRxXOK9wptN3kYWkzNKJdWIo00GyMDcJduEPg1
HEX2eS7vAfNCanudKD1twheKAYUIvP1AR6q5guA6i/0XpbkDODAapMceFfeU114M
cldMegGq0UrqqY2lWjjWoWZhJHeeMNsCTXBeZcoGgnLr4oUu7aamcH7kOblceF9D
TlXs+VTDnmrvz5cG0hmkILT1YcUuH2j8ZDDfF0mZdq8YPxjMqMvABGaJSQORpBGc
j2f3VAHLsZtipsL4QTM/AV/0G4xJC6BAgH/PrPanTDld2XYUnbDIyGQZen4+HVfL
ee+/2Jc7Grpfc9tCYDRMaQBtbWV1Pk/WhANRRKgrxXQYzgBG4Fmayx6HiSNShUMR
EJ6DreRX+MWwg8Hk/lmSiPFdU3My/54xD7mQ1sFjs92F8mcTlfHroDBlCHRc4y1n
4nytaRx4berzITsn8zLJy5p3tK6r/3efMjVbLicmIcCa56SnTGcIUoz2Lw4tXHdL
6WraRRaVM8GKRD2w/Nf/RjN/SCCQGa76T9H/WBAaSkfeNRem8AtlqPpVXj5eR9lS
Oas6y4X2TjuSTQnEi3CHFulIJ346iuwr26tTRvPBNf/Lp4wKAU/NK9XlTG93DVi8
LEHKkkg8emDourZyLMTx5XPZoFbrKKccIRohQgQ4iqnvEKEqEihSlY/aA3LzLRmN
j1pxhvYnYqnHeqcE8A4IouPXOx4SvQCThsZnU+JAsNb4yE4y1G1d/tR0xwNgFsso
nKQgFDOFfMkiSsSiqkKoBNeIpBzKd88r3l8AshufmEFU0wm5/UNz0VPi2vymZnju
zJIjeNumHktbNKl4ZBDz7vLwbt1dRmL+RGxnQWJNKOA3GyFeNzTjtx2vKxEzcR4X
APex1YiHnATtq93Sz7edbAgxFYC2sGdN1LuaIDTV6cYZ2oLri1SxpXK+4uv/Nj0Q
6q9ycedAzFv1bzV6dQ+GtA5KOHdfJbYQJVZdIZsK5BA2K8pKBkCXaIoG+DfIhdMI
ixuUXCL+xYbRMfbwpah+ZU9byPNWAj6es++ILFiyyAstIPLVs/m77oj9ZsOf2JzA
ucnxHgyYzoQA8bH0/kx7s21o7vTEuRQsCFTnLreKzCf2ujBFxXQ5KrOuTS4Ijg7G
4z08fUVvpMnPLkXLGg88kSEH0GmcDjGV9NU5yUTRudD1AuGbxuXgvlHnwuqTkU1H
OyX1p0BThYFb00mC8SQx9BjESWvB+QRYweHck6j6DUKGUuxpR4qpElbNaywMRG10
5wNeparLcchwTorM7i2fuIpiB+znRbCN1Qo+Vqyqo+KkOYP5K/zBGUL5ZlRbtitj
1750303bigKYhN48zYNOFatj3MoOlzj5BeCUpNGEvqLhtv+LXadmYo8JjWs0U/XN
SVTHqmNjtEmlWzoTPV4r7Z7W655/sV5oXnWEWVeXxZkjx05Ni1gERZo4HagRI5tS
TzwFnOSCPqh2kg+UYqxAp5sbD5y6FFdyckGfDSqux8wQI4/hxhQruhZOa7DGwS6K
w2FcNLwyTjht04427cgZ/4TLisEaq2tRusjyvKQRwOJlzXOTy7pOkWK80tx4I+uB
8q8Ib1TyxDapMnzAOF+xOg/a5K1Dbqwr2TnWy/w3ueP11dTHrgcPhNqoJDbYEdRi
7yDRVqhnz6qXV6XINSO+E+yNceHAbhiS7mQ/v4u6NU+EVUwXXYKKJwyVG5Qa2DhN
TJrXOUfw2rG7adbtb56YwNTZOb11LDgrpCHD0+ixeBbb9UmYn+R3WtYZjLSuAQl2
pZEW5bqxmaXgo7OpDQizHR7KW8uEQXLimtI02/+JuekDnICrC4xgJTDSKfVQTuro
Ig2fqe2e/WONNr+xiz6iXbRG+xzfdq/y+omJqbi99Pmr9SzEHSuoTxqZsL6WS+bH
Q/jFOsx075/hcPBKymMfKMlLEjf5sNmC/vNKl2q+xtiH0cnQIC0SmjvyCvis2uZc
/U7WTOJh+aJ8bfkVcLSypjRCgN802ExFgQ86RCllO5G7xZBjZRO0TaPaYlaG8uUy
KaQvPrigx4CgZ/TPx98gbuU88iz/+92i607ulGLoltnyQuqZyJMIJxvpu5AiXSnD
iCsH210NUx6Es8MQNRPqY5zezN5FEh6LvN0yuLxhwiDV/mAQyPJt4zSsrmAoYuHc
bhqZ3GjUM/AqEEaKmpTVd1Liq1Hzluk9Ee25bIfhHwq19HbbM/RcldXuOaiXj5Pr
yr5sQwCARuqkXaRRdYlmhWRayWuNlw5KmJozJDRUA8Z+pj1ZSIQb7Ty6AAjGeNtL
D50W0XzejKnQiwX2QTWr74BqKViScMFrundmfC7ycAJZ+dXK5VlpXFIa1iz89Auf
BX8mCSOy9C9Lvr9DGHoxGjQjG9DPWse7NpYT2lC74IH7YshLvT5IP6h/Wh00MoB0
akf7HVMfGap1LylyjiMMUfnflGoue8pqppwqXklACBfxG4zHRKl1jyCJhcLITZGW
ElAcqhw5TZ1RwgRAJKmbnHB7kjbhCf9B5ui8T5oTW2JIxEsYpxtMKcq9n4b7+XN6
NmqivTu/kgjN33nlfZq4zgVdF4u8rfjNh4sp+mMQSN4/dVm9KOFxu+7saJc8qg4f
zzJpjYGYuksD9I74SnYYtU45D0ndREkYMGPRhOLddCeXDFaWxi3UUKWWbw3BmaPf
E+nchRvraXRa3gB7MIUBuO78RjzVcKGhG8P5+9RSdAjBkRSCTcP+3zeoqytKerjd
Ps+lH9yCaawaUHvyS0s36xdAy0YZObGcO1YwIzdQ3qjONYGNjluMRHmMUNOmZpzU
a9WhJO6Ss0NU2q0i3yNKqK7mMUdSLNTG6Afh5rSuilo99l0J56TXk3CmbBGhfrOr
HXkFoTurHL39xNvlWZXqUdvRWqI96BF+GzJe/r+rFhgIxjYoppOdpr0t980C3Dg/
gYtm/ow5KPQWh1qqOi8+dZUrqp1aCe+X+w4EHhy8ezGZ7drYh8qhXwRPWp2i+BFw
JvbnurJeSQU/zJ1g5CTnaZB2NpGKXNrLvD0HlAltbTVJzvV+fkDRq3KFBp5aNX4V
mamzjPuSmJC+RWuGkEw3GeC2LpCjI18ud+vhRsoDJI8Ic/SjOOfFKxbstKHd/hwp
Ko5S2BdE73h3LAXW84Zw4EIvCOq/kN4kiruOqD6NSL3td8mS5wMtrSX0y/zmVt02
ywvm2G870Qj3MGbjkdiY93u2Wd2+mWW20iSBrQm0rD21eCb+Bj85bIC6HPpSk3+6
mYJhPTlIWy6YedemCUy8oOwJPUfxOweU/QVpTRrKt+8c+/8BOY2p5ThraYBA6KXi
Seuql4iP34t3jE9kTi0Gw0C7vjuM0/CdrJBj6IfprF/uXKrcSf4Jq6+39L12pQE4
/BgjRDepdFx0MWT96/bRJW/GUbnasitkAbu+y4B9hetMgoWBhydAVsbsauWSRPIi
UTtl/xEuHvKglgEq3o0Q2lUWWiqcivFLIrU4oJuDTn7F8SXH8QmjpOjyr4rKt8kh
xBtLN8Ty09SKTIKEPQnV+xodEvLaoiBFwezHzoXIdzlnNgv5d9bv3j0+JWaP7IZa
0COXwNrm53U4glJg0pmQ38Ekkr+UmgnGSJ7Z3TD7gJVwG6Trx6qSSPqgMsmch4NK
uEoIsULiW878huIBOVvBFb7Q5CkWttACVKnVR9o32gGB+D6CfCDBMqlo1XsFXZsB
YYkj6XdIKy9JXbfSl3dP4ooRUwdqeNV6Goswj7ogaHas8Fvip6Il2Z8FLH1Ujcr4
B1XwkkcsWdWQn+/tQiR0+gN8k5BhJXHl9wKX9puKXoId1iRnDQQrFTOMjpjFMXqn
OffnPNdSrCO8V9dnTXhj7sL8D2ltXpcQxR2am7l0ncRn+A457O9huktt/LLV2vJg
r6kV5MDykusjOiGRYPZTIRzxZ76aTY79qciuGcCmOqyV1DlR43vzIW3IrWueElXq
i1rEfsjn8n0BGgf5nhWSUnMDMfpIy0AZ1wcTrjEiVBWV5J5pD/WGmgYQwYS4Yh9+
WV5w/Wc5LZHLqaUDhEzjY3IzyMWgXP5fpcXPN1oxYuKkw+GWbflO7JA7ow8dYn2N
oinDFI1YixDkgCRSi5WAKKZmfbgCg8BzoU7YEU9RiRZnnNmcwPAk+rLjH7IHv4Ge
jieQw806ERhWWfoK4GJNFpQlv2fSVQun2HoNuTFCJ8Js2q7wBXsdEMjFQW5jZZiT
1KXqR8jbjaSgwcPp8VOTKZDfpaFP/sAT28Av7c0dvTywnXn7gxD1aJ7OJIvAfCW7
A53spIGstGO+z3DumOd4sM9xeFnTTGYqgkrViiXbmckJE6r/bbLOSpxFXjVw8s2z
VO3oY01QZku+N646GFbol5Wy+ykJMoCcUAcn4OkVE/eaeX7V6XaScl2ftLrckAQq
OvncIGtZlN6DHyxFaapZ/vIw8+Hmajh9B02kHapDdnC1Puz591d7htYeP1q/GJJH
y+McyScBCXhkdT/afN468TPNp2bp9f08wRRrsiYEgYuVILdjLzTmgInAfJ2W1/m8
N5EGsYxku9dX4OdVL1gy/avY7JP419Gz3ke4cDphSmMpPo8rBMiLzmWEPjeLF953
SHMkwjyVdCwEu+sMRUA+FU9RtSq/sIFXSH5iOM1gFdwGhQzC0k1KJmgXIh+UPpNr
4IW1u++0/5twkK1FllS10rTACYhz7++TfqxLDaDRSxdytF4gUkuN03k5fkKo+tvW
mDAH3MaDiGNfeQ8TPxQnT9NLW12F04TvemaRJkh2gzqlX5qvaJmNIySjVHNVyc1G
X3bdciht2eitJovfhSwCM4T5ZIQhTIbnnOHolCUyQAWS3mq5C41p3WOTsf+5M31H
pM1Nr/t+KMnDJ8Lj7be+xMsZJ2dc8taA7iM8m9UaQ6ckgcdFtbr4dNokau8Tx44Q
EeUd4w3B1/1ahGI0G1OrBdFHrZ0mi5M3e19LG1OoDo2TuruX3t1J6msL3lf0ei6q
f07LrcOlfp+973xUReOER2S02v6rttu+HzyuY1/DwjyRtZohyK++v3NkCBPMyVix
rmypw9fuXgL6gPaBmANzcncoLCz7Tp9xZU97nh262OI13tfCB8+4k4RzZyW8MZ5L
q5+E7b/pXNf6k8jzjnAFua20LGi7EVSk2dEmS+0sY8+90qTiwAavJyPKH4NstjkR
DjeAMB6oyEZex4pSE+USw4vNAtv+o8lqVFF7BjqcfNvZmoiJ1szc0CuWyKm2XRNr
p0xfzWayQd2GLpuVW4vbv66FdK40JpZyFrZ9pjyfjs0CfosDzotMrUl/hsdw4lmY
qJ1BZlgHnexA0k2BqwdwcitlpJNHasfI52k6MLRkqf/nmf7Bwpqkw0ykKAGUXNT4
OHMuK6j6Ec4J4xcsealNT4YFL9TD4Z4iXWr2pX71/Pw/MwWTax1V1+XhFKAZ0QOq
ANynrrf1cRoBNrMIftfX1GaQyG/fkX71GlLzMjsSRd+xrVeHsthBjOrrBrv8DDii
PS6Du3YMyQvQLx9VKCvUSJWYqcF6yEMohAj2JNMb2RV4Y52QiAriYDxZ62xXaOX3
pzFNX/GnSv7j1p8o2leK5a0Ki0BL9vGKZbko9p4kxUVCAAQn4hOSnava0tLmrE1H
PPUk0sJ4bQl3Uv9DWRsCPEAxrwbtkGu1tEfS6gRt97js1WLIEXLXph/J6mw1gZyn
Qsu+Q0GyEiwdG8oRFpEjHXp5sQ98C2YRY5FvHom8MkyTxNov/OwPSsGUg8jrYBDv
o838cdmd5paToGoog5r6O4IFYbSVuCS+ZR0w5lN0qJ5DYkCUSXv1cw2AZGiSkFqY
rwSOmquYoBLpsIZOlo6sWpxrRPu6bTzwR1vh4F52TA3bzhDaxh4K5sOPyUU8//wF
xD2fEG+RN7OuhK8yK2HaUihQgAkz+98LClGrFMcaRVtbrECFr/jUDE8ufj/YC1g2
55ozt5NEBYkuEyPDwK/SJ2gWSN7Z53xyBX+0RkLCalu1hKupu568PkiTJ9wzis63
cQeL9hscwhomgikkB4dA8eqhILxuOkRuH/HwseCxkpraYN4fuECV1pnezoB0nGCy
xzPPt+KQ+8CZYQ4XL86YxhOBpXh3Q+6XAx6rjhwcqFLMX/2fqFBaGi4AuaK12aYV
i7ir+1FErO9zgJRamOop5BblNbl1UOAJyq11RnRn8Be2edWPFPSDciszFayvjmXm
PHrE4ZIXWn7ewkwOcqPR3RKP5rRcMcPIT1jnigdL2ssfugen9km3dJtLy361Bx2Y
Cqe5IuqWXtHCXZ0HlZE9XvWUW8fyVjdIaY3PzKEAazNJkIItIf+YwPLA7MMCIagg
CsawZbdl784GCPcr2AdeUlG02LUUcFreqvcBp2tKSeMZK1veysZLm4WnvP+5iyKh
udi9QO+jHWROMeOVJF3qcNoG5An4p3IihGzbRaaLyIO3BN4L6kyYITWQySSipuim
xvEtaF3BhNdCkuwfcJ77hRoAIduhAIhtxjrRFq/WQezpul2AjSnFnrdpI6F2YMiN
dVZXaUiPYdwec37h95hTe8xJCIcDoSSRNjCiTWhK4XbMQAzKufNDF8PnrE/p+/Ti
Pfrzgwf8dRNN1oYHEm9TgPPiBVJ3gKE4dh54uBRtbF/B7ErLkIsKSm1XRCq8EySu
K/gJz3j6wnYs8kMDhPURjE+66tmIg/+Vt71MERNLYsTjcBUNpPjari9SZih0fMbO
SNYT6EUgXWRBhDZ7vfiPCPjSHz5CB2e4I/ElNsH3IBwaz2zKpHT1u1q8VzMRU0fy
PZjm/Wfnd4y0HXEhl+djkW0rYjnSbitn5KhPaZTxXZ5zuVc8doawyS9p74lgGGwB
/tKa+TFH7y/DB0TqkpkC/+96wUBrZT6RSPRmEzYS50DDeK6497R90QC6Dx3qIPnl
W8eIQaI1lHj+e+qFp4D3rwcKLWFcKxj3bUCn8++URAOExiFEt6AW5Pgp7OsLiwxX
vcLX2CJO/4Me9ZuVEBAIvKVQv7/i26T8KrKHTIj9OJnttAeIy2I2h3QU80wltWil
D44wLE2avrCjhQvjV3yR0z7RwI99VYa5Enin8tP07gfTeheIS2vCxW2srB58ghLL
/RMwJvmZ7bspzafRTDBqRoxmYCDMs4u2tcg2WVePcIp+54IovTY5wCap+nR56r0v
MZeKCyJWFLykZ3ff0rvoyJGBgab1EFRbijj0IiiuE+inWQBF+UN8865A67Yzwz+6
SZ/h3lYmz1ugsfrBhV4Xa2q38RKoyLe79bjX3bZhRO7f3vrz6vbY5hSxb+xXAnNr
d9nj23r7zLSKounh8FIMsRvAigQrpXbu26LVApn6SjjT3dGpmyqO5lQNGvb5RMWE
cC98oNbVcqoe7K7BiBb51CabXToh20YS06bTDepqR797wpqbIz82V2PJ1LDJ7sba
OQDDE0RvqERzMWh0xynpmcskTmD1TLmkevgUyF9U+4Fm7LQIKsVggp5tlWuIqtYS
hvtILa7VdYW3GSrOu7w1isMKcJMu0ENgaOHXH4M1Kjlf09Xhc2sLWz2+y4tnLSFM
Xem1/HPVOXQEILurdFh/ccbWCkbSwA/JmSYogoDSzhkKKB8RDIBKZyDOXA2RUvPH
j2RnGjo6ZsK2ltJ3PyfWGLgOMovuYRFl1HvXrogXyEtHy+qQ4keS2zv9Ab+CWYoF
f8frFghDq4emrCj2X3TfEZzmdfLKVmsstAutuXjtKWk6u9f7yXfJjpp+3DV69Wjz
jRcf7z20+mcGdjvNnb+4cn5mVHCq73LydKS5az0+Mq/jitXyUymchKlOuoD94nX3
yk6JCerdQHrGQOu6sbUOaVs0kVHbs/PWbksCWjq1/4EgARc/EWDBbno4LpaaumUK
vUWKf+PVy8JqpgT0V/pFI7ZnhIDxgbBnpNLjmGyW5K34b7o4OB0LrhKpaVBqVP0Z
ms1Vx/703vChyRM21MEBQpZHrpCAdLeTK6IFU5H6bLrUlV0ojcV5rs2wQdVmeIaE
KpJAzLZP00CjPj6GM+6Rp9ZiyfRAMy76tCEUZIrISVKY+vijm4V+foFRz2ke8wLT
7bHCmi2d5un332HCBuplX7QRDKfP9FtHpNx75W03ABz5+zKwhAYm3Hvya4DPqveA
ZazET5CgCoIlA6ASo/ar5BUq5D7/w8D4YBd++JebQKf5uhmTumPfsmrf5f0dueAn
OiEjvt5nmP/043s64J1CNQrFUVE5kTjo+meF4uVb5GQjq4VKVVRIkbhhCehnvju5
dJXa2xf2z3lC3AchPQO6sigMVKMKiXp5t3S9/dPzysC+eNFCs8bJGUsZyOIOMGXB
0lUkzeuP1HxaF52UPfEWX+aaefvE8aObfhegYHtLyscN3plv1R6I/fcCtKHJIQnR
07nlCfQEFSiyK4rIlJN91mh7trWATID6QlVn4+y9w95Xfd2rV8d+HdPkfnAWpEV2
Yma+Uh1tGKCeNSf6s18jHanJB7aQrNtgOa9kfgDvJ+StO/2FTg/kaUch/C/Unruv
ns3aEc3bSG2tSzMUQzSb8W1qICIuW2KVYshy9TdBDzB6rRbiQIXQuPQHR2i7KytV
sN/nVOl6GVhiovN1NSUqW+/+vQmA5yrsHe/vZB8P2vfInUn1Hp8bwqL9LihsSFgf
8kRIh4IHMsWmz8B7hQbgTq8UL3S74cgi0RC2N0EfM31Ix1mTLgamz8tIFXSHCBg/
95p9+24WBHK/TeU6sU39sMtTFpTGr+dtOUMVx50ltuDVrX21y8IRecnfErGBzLBb
1vd8RU/BJ3X5YAeZRV0Ktc7PXgtCaIuq2DDH9/ta0anbd7uw+gOlxuthW8x21GcB
PkH3BvqnWsByZjh5vTUojOnzAE6hGflJY1VGsSTf0PzM2P0Q7gad9RT4+veWRY/T
vClRED4Ut9oN1mGVK40+r9XgkIDKT1UpVIXkaCEEH0aR8+DF7kx7TuzVgZ2R5JZi
62YZV3dTHYhRYWLjbLsFNqzhF6YdYf/5ZQRMT6gdDrNLLamWNQzt8NZRvzlbEhtc
o5eJ3IsSPyNyt5mVPGY02VYMtRVzi42aSiubtgd8XhZry27Fw+SUR6TQmHAy5bmx
B6jLnasv7Yr6d6emtjjj3QGsa81BMlOZx9ojoL4pAZbdiUuuouoax5mYgvfI/6pG
NPU3uRMihMVUE6y/l4TjS40uL6SjqhwQTAHF2mWXmGZmN7wh70+xWPR7/p3ZLcvv
uBVPLAr5zkmfriF+S021/fPeM56Gj+QnTssJMpyUOWFPEywuVvVrlxDa3llYnwXx
e/GmPd+P1IvWoRYSv4RXhy9j1RtKHmxdcSq296J8GuDxEv4QF6tQcuJFjgHveoLG
Yzb4LuRoP9CD7EVYVr73DYosF/yg40uZLVKxM3YtiS4hbgxrfNGuWuP++PYQNeXi
lvzWPrv7IcAkiov1dCvgG5sKD1TCOPwfA12cKkyCQdD13EvVMSKyNtEkaXGPGmpU
QA+BjHl+dnztQLKcraDrMe3hWHQKoaNyW2vaYbtESHpVRg00Xk4Hhg/lDcRM5bP2
lDBrhuwYtChd23UTskoEmEw2/k1/UE6gV/f5jcELAQkSguvV4h4jw1hQWStUHVyH
hqI3OzFdz/C8xHpfciZIKOzsT9d90Pdkz17hoaTOCw2H6cMR6tA/vT7HvRXM6mSr
l9l/1R7u+rVzOGo/L6C+C5W2h8TdCQRVCK3K1La3I5xw+GfFczq072DgIkeAxTeQ
yJjet8eznVu1GC4/P/Zcw1swhj524zCKmq9Hk8P4y8mhuVb8P6ftQvJ1gzkZ6FqN
hTppTrTBfYhZuG9EkUS97UUCV5KvLeZ2KbPmJjb4YiTdjuWcSO9uGotPsAdSS/Wq
C/Hbte5x1EqKDhqZ88+3huhjA01tWR1S6VjaanRCBgnUdZJy0tOxeGD8MgvO0R2j
atuZ/ZrLRsonAjts6uul4wh8YkUa5OvbZDhhJ45N8GMtTsZ+YryDuCDMNX0NUT4H
qlcjr+l+m9+qwpNXxu6tLfBeavBeFkI3/n8UsJU8dKv106hWDOA1c542RpdZLZTt
aombmM5XTNwddCwqTBEQ9+Fsdl8fYTzKGmInYN+z3M4H6QjmAP0EABnRbS9iSqoV
8UymvIOD2WAmUZbsDwfVrryCWSTRUbCee+HMABG7aWBfQ+Rkn9D2PeXhKriTyslL
JDnZlxAwtkGKQtw75kA8vAPpC8wmksLKTQ4wlfHc+OyG0MdvdgJOOR/ebadnCxer
Ym8sG0xra/VAb/90g6neygyTar+6iiWVmL5B6nvEhcwYjYDyB36C/gfJ+Zj3IsVw
GIQf7p9l83vEF/BNLq5u/Xxny+S93q+3+Ui9vS7IP9nQGxqNM5BstXNg00V643xm
dHChelqYnjPrd3FlbyWF/xRyK9sXiF+PZjz3Qn8hD0gwlITEyX8FPk/AfNM47qcM
WuutGIOu53jlgoLGCibXGFmWG4b7PNXdQCE9Cujy7EuxJUx59mnoGn3L8+eCFXt3
pbIfJPid1I6oWm/0NAzG4XnNY5kTuzv8I/V36JI51el7CnjIcmNQA05SXMkNlLVr
8ImhY+WMNT2JNmbV3ap5Sqjxy82UKcMOs0y2jxZMTWccHOueM6I7gIRj0wiFzL59
KzUSjival3ZyyeoiyE+GPmRMG7J0pKJHntL8hYYYEOz8laGys8Dt/tPoeX9/nLME
Vf6675h7/2zVw156gn5zoZcaOhBuvbDLKgIz0YF86XaNp+AFdyYwGG65xTghvsTc
fkDvo4EOY4ADSNwp1i9J6sQkKPI80zGTNO1M71/ZaG2NqQ6fjHtX+/IW06DofLsr
4ca8+XfpNB9IRdKlv5xleTBnDeph8K2GchRIlXOiRUeYwdq9U/Pxp28bCd3A8mSp
5rOEuTV27N6YieGIB3zeLVIXFFtO9ZkJ/jrUrnFrSxAGSKIIx8QHHVElLkJG5ikR
aBkREtdyxhhNjcZOgKN1BuvjY6LMiNLzlQ/E5X2xRbge4eVusD+LF8YGl8oZWIHL
pMH6f1U1CuMm1D9iqyVt2+5K9tC8XftOUJVnG7LbNNx47wIkxNJdHP+5tw3vlUhE
AY6pqCNFLONbEJ2HYmk3iqFp3tIiulwlNVf8s5mQDinMJ9d4oNrG1/TXqlxJDH3J
BcySVjF0EGWLDeiDXYnQ0yYacfBPE+GBsWNfXskMZO4AAZT1noW4u/O04VaA0PZp
o1MNrrclhBx49XACg/O8SJJLrkzKCBN3pqB77rFke/B3bfYQXyG0CSNegXWw66df
+OCbpTm7iYZPJbmZvTtVslg79CT1SlV8hPXPu3Ap5FhOO3sXFdRcsAawIZIMx7KZ
TtRUeY3SFDDZD7vPROADe4Ee7YZzS/xSpSGkssyUxMl5TIWsOjMa7LXpbUKBnyN6
7k7h79V+QZEUWsWLC3nasp4SDBIVmqH+szkdN15Q4DlRDRi6i7Oo410Hc92pbyRl
x+id+usccyOm1/nuiFDB2Fcaw5b6/h52bMAYeuJT2ekpm4VjDmupuJjQWKPsrb3r
/f4EZcRASAYpHBFHMzbAfPwe/lFKr10E4jXptm8DcUs7B0ojTwyVY0Q5M6Fg+fnM
a04akevsqCwY3kW8Mu97vmSRyVhnCHPhOLbFfUUUcw7KZ6lPRAHlEjlHaCXF/pWv
2jsP00//0PXjo8uYSebd8/qEqArtjVOtm7HSaQ4HvRRFGDGmLKt1gZUP6qTyfalw
Hn8yJT5Z4nK//4ukdv1Ukfs/OJe7LRMeiThQXnAN45hbCXVniS0wsTea5Mfr8PaW
/UfZJFZYNmxw35ASTKeJ8vAW8IuQ2hmZSLx3Rrj8iMaRqgvRa3KoPBVrzSs3GKVg
JiihW13RXR0z+H4G/lJ9LOglWHQ5+bv9/EJrroh5QZn/iCW/I1tqNdEmZdhQoUVg
a8Lu0lHrdpjEVl1vN9fEd0jEbyZaHK91AeKXDrchkYRTM4+FRrFkEYyCUWIJWQ9a
ZyaKjTt3Sp525eLbAf6ffOhdUqnsvSzu3QdMzGEzerbaXp/5Jj31y6aermFOFK2o
QK3vOEgK4qlLMe956csQ3EjypnmCofvyqxE6lXBiz8jvu+NctVu4QmonyeQ1449C
LtyMLt/Tv06wFCnl3En6mjiIF0zEu6vkqpUIpD6yKtD5/WUZT82vlqBHigWSbFef
G3Si1eA0qBZhJJVfCg+4CLMVZw7aPNO97nwsIrFu7jE9pVYlxoqnpaStWnu8kWsy
mHoJrmuAUOuLZi7AwvopuRuss7jLbmBt7o2LeD4nBfFtkxf/kEYjQbowbUFZ1dK8
opS0NDGQ9OEAE1U7trero1mD37tME2Xjgj5iDNVYT43hdKz+NPb+t0m2zj39kE/L
WX+bguTxJBeclmnBGL4LiaLlGKa8QEmrUjCpCYBTLJYQYLeQMraXBG8/XthQMnnr
bqhAmko7HlPSdIdmzhMuh2ad6MYQA2zCEpwgzBQDNPKXuu6LMCrH4ERbcytmrUb0
RjDwMsKK1+iR0f+4ozvwOrrtkSjYN7J/FCzdnef9+A1AzZgGzdnimZ5symvnTH2U
0+b1CiXDvOMJOy/1ozai46sSKUepkLJ2rGZ9LiHLTaOkZrBuUW5ADt29S1DAhFlk
ip6ZPuZWL7034rhtVU3zHmNM5kvDzJZjFZfeJ3t+hNOd0IbvUTe5iBe5tqUpIAoO
VdOxPJjwPIM3ES+WzO7bFOtUozgvcDoyNGncq4orqZQoDcU1qUFogxA1YOw22bOP
zRijEpAxjXqgwIvvPuR51jrxqN87YOhID1kPYneJiSzm3ZnezpMvMKSuzJzxVV7V
yqFlLRhqhAlK4rXgzaIqZkManDmW6vT2e9MlNixuDXp4XB93lGG27X6gMcY8bhEx
VG4UqOdo62rls4MJ+yRCpGP0hHGCGuIblEVnqjtdN/9RBT8oQio/kCguESpI6r3C
HtBHV4dp6+l2uhd8VJK773YujFmNe2qz+DRS+zLB7PgvPwrcDKp91e4UCMy4++xX
mk2/4drlajcGTyFbk+aZR9OuAKhz1X+HFVNdeUkOfayt9eFCP2zJB57BbM1NkbTf
j0l0KiO5VD8W/DeskiSa236R/Kndz/qERkRPxyvkWJvZNmBGbRiDOXlhQYBZvFk8
wDtGoUJWChLf4iU0gMNtkToMmr9Sa7HdcdHE4XoNRKpB6VD9NjA+qWzoGrN5Gi3J
+BSu2hxuAXeDQH4ZeFuwmYcxi8/mesFQjcE8cMolFNhohpBuTMA1Sjq7Eldpnz0c
feBPEkpba680mSQDWf5E7W1dMpU61o2osifgvORsHC/zsvVUn8ptqUhch4QXudjh
8W1+tUqD737euVEvWhlAPBkL31PgJ/iD9SnxW61OFqfAbQas0oieVlJz2lGSviI3
57q9n4f67fCcBEYxGq6Mq+YiMa7l4dV6vsMSPlDdZImcej65ge0gRUCL0tBLcXtu
OE4Quk3Elua9xJsEI7uNXJHg7qN2z6Vy0TVFrR7wtmNIJSw9ewO7TUjOQv0wQLun
Wn4//CrUVYZ7kz6NvUDyucNaUiSabUhzPhSNjS+vbngkb3q3DjKSNKhOmlUXkFYQ
cdy5xOZZG7UuB9RqJ8gUxmOC9REx39AJrmQNhJC7UP+b7qMlU/j3JEBvdum9EFe1
G7CDKXDbCtu8mHK1PAToA7qiVucl76/xkkPG/2nUvj6qRu8Xbdsvtb5cbvtCf9vA
cXR4kMjqnJwuI3ER07Pz62m+gu6dR9vE3mnYCLtYEkYHQzegFJMwpylcAPau7BYe
ORKwegTDQfCyYOmPn8PFQuOQpHInTKvY37qYz7KtA8A4TVC6AEcgveFoWGvO0f9v
PKImaXCoVWKaBXeJG0VPdQeAIzYmn+8AoOh1k2wNZF94DmFUu82MrfJKvXVK2kQD
4LY04Rx0Azp+Y/g1AT+1YkH/gkHOZjLfyM1ryUtd0oLRlw/Mj2nKhskpmhU1eWAE
vFtnsqhw1r4Dvfmgv+EJakav+W0rEGRO3l+dFn8GXe10HH0htUdRpIxYS5e++XSn
iM3U+4I/fAZc/Bu2KoSy0WCtHxbCvncfU46x7VEoeRMmQRWneTWTdE/mURYEbc1J
ZZHe9LtQZU2opcavbDIhpt6gxJSaqRd8PW5utV0kfrAfM5w1Z7Hhsp14BZ097KT7
9x28aPajPqzXHWNjUg2+6rmELMAJSa7rOtGXrOpkIRO6+xAx3LAhclYyWEYxuGeo
Wxjgg3kpUvufvCA/QOVWPaoIAqLjs8qUrEL08zV5jAZy/8wGTPzcryH77t7u2N08
erzNhwkDZMEzRptbjHpwxMQINeEgXEc3FFec61f9N8Hotk2xSDW0Ukhppy4twI88
1YwheRZ9cufJJGs4dfYdS06fqu9prYrU7N8VHnR6x1hHviEl1TA3aYKxQ66WZ0cf
m3Esl6JotYO2KnEerzeEBMEJrs8DO/lghN3WvdSLmtcS5YuRTLMAbarIqajLHFff
693q7xfGzaLlL/pM114+RXIdjNO2UDBPos7ubF0D7NJGnDIkfHCt2sT+PqbQ1tve
eWdDzmwMD2XgOPu0EyEcG0SlBil9jVCL5H7QFbqxs5raJcB4fGa8W/YD/RtzZbQ2
nK63XlQ7MRY5LBzeXW3/OO7zlsZcC8iVsbzr5YndvhswiU7QFuT89ehRqct03e8Q
mWuG0mJgo2YHp2fvQ0QFYKLwc75+uvfHHJVL0Yq8T/JI8319rOp8PFjRCsGcO8XX
kEexlq2hYkBhSeJ7FwXUHsapeY22pkuiPuXZ2FT535+I+Q3r67hE63gqBLMNtdPa
6zidoNaK2nqSyA2IH4gYE8+oXRHwfIqABvl3cx0/7IUidETxSKS5djixMGTa4T2D
AVMrQJS8FmNKkOKXa+NplPke4bjDHzv7gmfAxoqkQGkGp7x6+xgIO1LgWQAVlZDW
DlRkTJfHwP5rQg1l9/Wkgg6rHUpXhflQOhC7CxkAP7EEMQqAhNRM21ZjwU/+qSsh
wQlMnNWzUWok/vzP/sm4wcKPAYuBAAK2zmZbv7t2hkzVcLE49jPX73VjwLJSCOTK
gY01/F8fae59j/5qSFTkQhVIMRBciAHVXDq5ixPiJalTD1j33I4Iu7MxYwA8xoge
37qPWbKRZLzQSdYzN06i8B/Gs/JwDIhE2WhfD78DyS3bSDGHHOBDa66KcaxIZpVf
3VYjpJp7H7Ehb8e5ogwNzYFaSQGa7FwVGgwZKdbmHJjM60zgKMQ0h2m5gJWr6GNi
OkEGYL8IJ1voFpADsV/7UivYSkxEMMBjYqJ/2WhuCNqCoztul1iAbeapBTIiUY8t
MRQ89425ACtrpewn14uhIWNp0Ub1xR3U2PCj7yA+03aJ3vZxjOf44VGctIMjF8+p
7RMZmQfYFXOvP8B1h6F19nSHXxE5C+qP7+bNAhwV6IzabXE5lPc9W3exNqghxNgx
oS5RahegSyPPJWS59K8S2EzgtFC0nR5GTcRBeAemQm7McdXTq8yD4jglaHZsKj3p
qSU53pDm49UaARUJyU3nLLVaL/gXkI/VYj4XrX3AWPPEpAyEn9t17y1KenzS1eqB
wlIhrxJxQ8Oiesla+h5836tWNWkI04//jxvDoiV/8+y7cQ5KVHeiaGLKDGJ/OQC5
qn9TLxKiGrQUw8E6ScssIWYc/wD0jZHSjPGVZx8MEa6mLN3m21p45+v/jUoQsT2v
vwAy0wdRauuwPgTdSRO80VJs5nnHCgyMhW8JJ59/5Ea6suujQ//GjF4hIZuTSPJc
PiOp9dcGy3pRHusPK6gtLWiAWpAAO/9WeYRhYCbyvFyQ/FLu290JwRt78HkSUplv
tbFL6rpboN66+6f460RXZ46JXbB233ZKw8602QhCbYNwSvXm5PwyzXmyZzYNeTCN
VkxL3cHgKVWgxvjwwI87olkH9j6JQRxUeFEHQcQ6kTvmTS+VVxDHN3VQazi2cien
FSPCmT8EaY+EmYkhvt7IvWEDF2TNELKIHMJOMkRHt3Sq6GTl2wcGmvYMfnsrKemX
jHdLMMZiPMt9QLUlDrdZ+1nVNRl1EiUKshS0rh7HmigjF/628J9vYRXU1pjEuJml
gTwLrMk+ntLBc2h208ne6j032hLZDShRdl0dIFge6IZcCnwTPpQ89DR2wce7pChN
1teFpupPgb2f9syvtWZcGmca16UnPYOGWq2Z4JON9ZER1iIjL+6B87HRgz8sOw/2
nTZcZutbZiCLw5JT0qCHdOJ9SSKSIoWzPusdZi2sFS2IfO2jkBWgTXcfYSbvWMx2
aKkGbT/79azgDNlWUi7m40steyL5RejCCyTO9Rt9GS24qaxD1IHKa+RNq1H2hAaV
XgMZfWWmc6U5J8HvcBOOXkqNPESDX5nBkdaW3vwBDLFWTml2U2vsDOYYzp6jE9K/
+6YAbVxkq9jPHhccLxuHSZKWJ4v9h802D4KUYnZ2XMrYikW5J6DII0goqrmiNhDi
SfSdcVeOV6e5+X6iv+mCWgspPkH66xNYYk5Qm46FFgefQp46n22sozNyRRu55qGh
+0/3M6Yq5J4snqz7bNpuamf2w5OvYGWlOlMVPt40QRlMcSvqKoVNVZN+MQuwm2Od
be9QG8OXYxVxqcTpzNCAFcU3LxeDFD4ahVlD1x7SF/thI2lUNfJprNXSWwAu5r2P
aVDbBhzsxf1d1OID+ZEeATFYyAeJt4U2WBOnSVKo1j6AG/MOqlU2dLfwZxCA+y5T
lKCTZtJEzn3rK/ROFyHkD8hYM5kGU5fSguZJ2Rd6teA/5RJ731x4gi/Iv38xqSS1
LGsxKs6gK8LMDTUQ8MqbwIm+yGt0VqEdZNPsxVB9dpJL8rq/zd7Zq3j2XBu9uKE7
5xf/esCXl+SqGNuxHWHE55cowmx1Sp7FbGq6ah8ZXqsD2W4jvkxTAGXw+WP1BDSX
5Hfg5/B1UKfgRPU3KRV69qlkutHr0wGIxMRnVhxZoEkkbBgMeAUem2fZL388obwk
YsUa0GqurFpIMHCugkhWQRZV7JzV6RozDzSIQCfZN/A6rPr/DhZISdbbGnWc4tdH
4B9sYvtMTxCIKOvEmUNJtnMC71e16LzzDRJjc9suXyLv+iQR6q2/BfwHfrv4tgTy
ZjSwilmbfrbzPG476r+f0sHA/5Gm+Tri0fpTauqnIHoSUFwVY8AYMOHlL3BSlody
ISU3YYQw6CnM3EcXWP00OedG6pDMrY7zEd8G8tNYjFAZK20zjtYOdNpyN3chhSsW
lCUf/OuYKaER0ZV9FrsVZvGJ0hG4iguJAg4krymHsIV3MIRui5DHkX9uv6wBB+ZY
RmD00S9LzwlrFPmbkaezZmNh5oum/03Lfhzq/CjgnAnyn0ZZpjmJND9oynPgf5zB
KEjOWf6o32plx96iIRfzVp9iZyDBGC+mAc4D21lu511qiaHPHnx6CEF7xCUsW5n5
++bL//ylF1iGz4MlgV3wr+OMSzGJhaIlLuVfKdbsCsw2Jf2oQvlcVsu4edUeYfr3
pBzieS2cvCYlUCcDOrCnLgh+N8h3RkP0RavkN8NW4KxcelVak3twOxY/batvTG9g
N1RvwKw7a/NAxkduMIqyL+ftkmf+WvkTAm3ruOQmOyZ0KmGiaCnNx3wOAtbNJFeq
PrFkAGB3RKsMXaLG0mXikML7YOoTEagG7qGhUv3htx4FaSk+H6cbKIqUpzXwE0RB
mXlyGLPGP1S8/YpDgPla6DIH95ekuBGJgSqjLwLrKsSWqk3pJU6FQ6bP6TDqXJq8
a546XeT6vL8TOPYXDLlBHAM1BcHTbc3A1DePeZdI/wfsskQlEmBc3bRgbgXyO1zj
uTe1yAcnsiklrX/yXrWPEyABUmThCPpZfcOgnMnYethTIIMip+sutXtqNW4BW+Ec
Qx55GLHvhauCLh8/kxHBRtgecQOwLMvic2KkjkDLvNfGUalrJW15zxufS4nfsQYQ
6tKaRhsBIFbGQOIMS9AUNvchEWJmdyyaOTUlHBT/g6DUxFyLbGoGGX7dH1Ui+MSh
5jxxV/l1ziKJqiSnqvFCu/gR/Y2vAJ81z4jf51mqFLxs9GxsUtEPa0NX23mELhfU
TLJXAX9pO0v/8j2bZ7p8PiK8HtGsLMlUfZwblqVQSfu7Dkd936FYHZsMTAkS2lLd
W+6Oqlzk+WZmnatrdrsP3Ic6OF/fNBpG1FAi9mxazQ9+kejpv0Vg8lGjqHv7gEbu
BDwPmnb4DkceIdaMFLOUru2j8zqN8qkbzlp3X8n/u1HQeKKf0WnpN19g/0+oPOe0
vXe2i3NP0dhLcAy6qanlRiZXo0ijVWLV7W6qZkHq024cXN18oKH3L+9zFu4+JT8Z
LdADoFkgP4Le8O0Via+vhxtImDc2HIsIaJIBJWFyZf9zFbWtcD/64nbCkRBOq+SA
r4hZLw/Vmu68h/37dueWBMVnO86za+tCs7Zgq7h9mRPp2x5JPCEIzB8Rm+T7wixa
+vKmJ4y9BIV7KsnU3uOKLK2wrx3K3iBztqjYY0TLr9hALhx1CF9CC0IMJh9kgpON
SnlsDGmbee8PxBhMXFbijMAcJtdnwQPUBnIxYm8EEAMFIFkAIrUXOB+doM6QnwdA
zeC8vyCU8dQPTOIFKJvxDc/uvtP1+lTFIRe0Sq6Ax4DrzB1xgQnx0jHTbTnNAHA2
vy9uKz95qWk19Ug5PpfgsNYZvPBSePJ+RPqh2T3fkvO0UYUqA5IvCHXQMNY8Mmio
fOiScrTb8FDhV1cnBwigX8fIJ6rsSC5PfeduBqc0c4IJ/x5aa/U7orjo30EFyHad
YQ4qBWi9W1+5Ed/+7U/mZuLmNNzBmsezma3vXAh35zrLkN16sE+wmGzLdesNJ7QO
TBU/TTu1Zm3mBU8Za/OIwj0+L0Cylt25MlGNf6lRhc8Yrt+yYX22X/VHA68fCDly
ifDaBrMs1zMa7DCI9w8a8DgpvwJUKcTMQrrC24Ata+ehq5mWk1ta2Njt0NnOkSpk
8uktnUeoMane0s8iA3LAGlhKns8APstG9SnVtjnw5mBoXiTbEyB1nDx0b0QDSxsT
bEw/HQaj0JKvKhxQulYI81+gK8+/iZfLIpYUYx35uJoDNSuX94oOeTXtitktG4LQ
OxXUwlw7LcG1ezqCMB0FT9+Vd/cuJHja0pkCcxNXI+JR3DE6FigHwrvInutF4Goj
r2g6RIK38S2b/KG6vM4VwUjoXxFxbOk6QuM1RMZNM+0CPC9zpcsEf1X88q0hSea4
q0lQPSsILnF3uDevMFzR9cJ43Dudm3zBUgcp4Ohz0t81zpI00bwP8LcVMJOY2BVt
WMkeN/IRrDkMsteGSM8NEUImwP4HkcjdHuzYU64VV+bkHDFt+tw3xGh+Prr4B7V/
Mm9CBrrUgwybQBcPvejgtCpexN8tE5vB6Th8i8vAukorPTcZ9XVTHYR6SvCMaoIz
jv+pDeniD3Hl2CJyHByGvaP/Z/M3JSj5pgIwDMr0siZL/91qlI66AuursGorMx1R
fwTVLyUWXZR/QobQyhb9BoeDsp24LP2992e+HuVIJnB9HO41IA4Oh0wDfsNB/G4y
BsVAaIOJYQP6/9VZjpevzUxqLk1mIZpXSS1crzyRTa+MXmlg5JPhgFIHIj+ZOcOI
GSYGubTVMYVDUR3LzVpDSEuzh+WvSk773k9W0YvFLR+19cGc8OmCuiZx6J+i/5UJ
0lJIBoA62FD3HRxtgKCxuP9ucHqae0CY0N/dB38h1cTPMa6rQVoit5r6fKGeegjI
WxhllEe/ysEXsMpkJsBIQsQInl+2lRCxx11kFELTrR5cv2l5RK3BJif0RIV57jjc
vh5LRd5+GMqMH+QbKM88GqgFJ9vHpLCp2FCZLAiYgzuCKfMYoD/ulpF2thDgLZ30
GtY0awM0n7aKQS2GI7edCTxDE5n0sIiO8/a/zPstuUnSir7gh3sMSBv+sACm93oi
qj7DqW54Jc7qkM4kiuy4cBAMgrbMsH0yW1Fsrq9MPy/5su12TwYKP1r8OGkyDOqG
kmuSKtejsFdgOu3MpaFmNeXqin9WcxUDvTUG6Q4bZEmSrSIcp7BeuycQ1gTLPIxr
9KbGa6b/mYi1V39cFXxkafrDm3OgvRMe28FLrgEyrmXnjqwSr14I4auSpylEPm3Y
0/7Mc2p2GsA98Z62+BSzZRGyA7NNpTvL1ohL2ufM7wDYgva/FqQhIvGiR2f3qYm7
PDsysrrbn9dIGW442FsrB1dk5G2y6QS7frqBPWrjOagEBf85GPu8U0eajAPf6BHn
kaa/uNx9S1FL/VitrRh7di9ckMXaf0uiLSWt87liTGRZoznO7B7IJmj5IS1dXoew
HYXsPtoCQKZZ2kZc4P5H1rXURMPQHq0f20Egoet1yt5Ehf2eCnyMcVn57VYiuOl3
EVn5x2O7mG0yXqsIF5q+ZK2Q1ueixU0rjGnYST+CMVkHiYragoKHXliMMfxgyYqP
5PHkjjM++XAFcb5I0S0ol7GMqzhs9ENrDJM49b4WP4Yti8NvaXPLkpvej5K+mnMl
nmWfejyFI7xsIyXWp7iVpqhvTeSEMAdoO2ru+Lo00felZqaNfEkf1RL1BfLdF23C
8br6ufJzxCO/UrhejHJan8FdQAV7i3uyOBeVbA9SWTgz918y/blZtGhfds75ix17
VMTdu+4Md4KvTfYheXHKBTOdHe+9DC+CN1b0tR2ZtfCLEA5re1YYGu9AbuLXVUQ3
ILy9KHKJEMiIOzKkvgJOE89Lv+0TUkxB0lyH94RS/CriVOdxeiG5P8uj01IH/ZId
EdMNY5YzM+Q9J5lsLXWYe5aMBETbjOX0jv0xQaePUk8nivquQPPOuX68v0+w+E0K
9G9LiI02SjLbI9rr0su+ps/g+AjdTArCnVVQbqjp1eZnE7CEr4Pq3y0WTYfryHc1
YamkEiuXldtdYjQJfRZPi8O/0nUG6Iem8Znl1rK1N1UKJFXm4sOOXbuNZ2OFInJL
p1LndqmfuORy8KUkN/9r16nqBlk/D2E8duyAylukF3YcNnJ5J9TMd/IJCaATYE33
yAZw/Te8NA4SbhBtBbxut+fAKIJG4IkZ/QqO3lmac09MhO3ISdpN1Fcqr647PTEV
fLUgtoR9lxAIMMudssLTGMWwA7tIWP6hqiE/3YgcMAoeCeDSFriJB+/r9LyQnrtL
PRMCeXnvGsQl7JKq8BHQs55mGOAP6GTs7FzHxv2bPFDZkC/kCpJlMv7h6apeKTjR
FENtRZ35CYnLvBTJbsHDGkQVmdjukfSkOmV+gKjPaVpH9Gyrdf2JenUeHMmPqak6
1d+TsSN6d/pMkvPiJ8mhR/cO/sfYANdPfZKf0B1JE6p/VoDK2ECJuDupXHzafzhi
G7TZDSXtSz7gNtpk8BEuGs4vuTjY3Va1brovmztjj1Z00JebpP+7OfEgEayy7/7g
uh4s9yMBmCjKlMSE2w+1yx3JOonPRYzVSnqRpldeQ316WIuGo3lo45Iyw3sv+aiO
ShbqSvxEyFPf9SGUo7fJiB7HMHGFdBE85Fforl8/+zVLYKn3n6kfD9I8TxATuppt
hG8v1psNFhIOKb5dso697XdJYLfyGfHZQsdUbBedoCP28Vqf7Is1DDmCF2dEB2qO
p0yi8oiDhDGbvOkk8dW9/gyVHpsR7KY+Als2N2ES/BoaHS3S6EhlY0jrbeGACHon
IGcxDqXM5QeFPcn2pFQpaC2z3PzbrwuMMnHOVdd5c2SRP3Cbuv4304fTEXy8gJav
Jn852+WysLlyByL219tm2Rr8sObzjmxArwZLCM1TDNdJ2Khgp+elgBRSMjLkgzn8
zsp9c/gRWud/FQd7J+Xd8h0J8cHSncn63i1auxpQsp1hoxysYRwEg6Ee+7eAFXg8
UDo8UMgC/RVOlyv+BPl9LHuzC/7fG2gVvw9H4NWEB8wI0zyE249s5ysLaEJt4tU7
XdQlKc5u/2S07NDxRZ1UtglPzib7ltvRoUUkILK+XEfxhdlY0usuABnwmyVZAM/R
J5mYYwF46tMAJnv1MiUCmIvZK8HxyTppLEPtQKDR6eRYbmVXLLiYKX8kTGp1cQSH
4GZa/kLATIMthQCVHSHMyyoxhhvDJbOSQvntGG4yzA/lkHMiQ0kSYVmQ94EFsk14
RZT7Yj3OVHX9nDH1zaQNOIxp0j4ksBwipx4473xN4E/vJybmw8xZSro788KxdkRG
nPGraXiEybsM2Xl6IIWSnp8Hx8Fr1u13Dxaehq8zMNfMBqZUskaIcilSAN2E9/x3
e+Tm4KCGtpdOEFQqFVJ8QLFWm6QD8oaXGZW9IdYOSpze7OAgH5pgwFd5JQSO3NlR
a3E5DT0EGnkeqXsofPuZQaFdDPfWRtr8cabj0lDcXNHCDm0B167/H4ntt85edTgu
G5/x/mH9YyFwtbWIK9C4ojV8+NkFJmMlYcxYyP8lBdwkhhlyYho3jQU5pajO5H5e
41/SM4fIRDLtQ4NPdTRrtjwIwK8GlkLRSlGPWmhz4+usEhlIMUwuumbcEH2kjLL4
aB7CrJP/AfO/Iv97LLV7bMw8Ra1hY7891Jht9VGQ+O2W7BZYIN/7W3sAQiXtBngu
KxRKPxBw3nshwxxjOZFEd5RNPkLWZxV/PBvUHE8ta7CHvOX501N8zH6ZDAzwZQ2o
HByRQ19A1U8qOI7PVQrn913a6SQN8ABjX051CnNnHbqF6FLWeSrjj+DLU+jjMWV5
UrIDm5h7WpjlWZC6aTTs2kQ4fD1j/VGyYCcxdjvTqdD5fN8QdwoqF8v2S79+nzD7
ecYhTddJOUYE83JrXKYmMWPYXtLaqLOMYf/vI20QoaqeHbulAe0BZdrU2u/C1Oui
3j04akAuJI+D21Z1NJqH0u9ainGLwp1ab22yN0ftdT65jLewYBxuD/7l+mGwgekr
Eh8HZQnJ07yMXN/4uwn2G8zIVv0XdpNrKvj6ub911TQn5kd6nwz81LPtbbBUBG0K
tkDTIzn+M76doZ0L3Qxxe48xmFiigWDV15WcHQ5FIhDYpUj9pzUdgvBBtmwAdD1n
Svfr53HTi2N8QWBpMAdHxiYqWjHqp/yxAm6+jI1CX2GhlrO3iAYEvwGprSYepYpy
QqWVK9kJ2WnwZmOSDQYUGn8EzxgQh/pRWkT7Qi96pTPX4NK0eEEYOijmQvMFtsMQ
ZwDq9umDYyt4kt2NMi3SGbVCnVaqOQ5++j9TiFib/TocKH3WqzqTX3ZE0F0S2cCc
2gHsUkWIFVAw4PIGRf8uf+hJ1PUySuX/ZKzMljBYfWrno97jheh0Wg1rI8QFA+zB
+iTgkcWuOdOILBoBnJ1BOicJ0w7UcfxBeUixE9twcnUqamuih0AXr0lOuAfzUZ89
3Yeh2RTomDOxlHyu/QtJ2ZSOx3QpYCmx8bbXBdkYmw2WaRjuRVfeNsxlXS79xDHw
Kq1O1zYkkheRJ85TZuSthyCudsAmrdcHXHvJuzxQW/ci+2TbHQlPYTREyR3mTxlV
jwZq/ReXrehDO65ta0YEj+HZBWuzABcjHYmuxip7vFd7mD1eawFqVTMh0twKYT+o
Q7J7hun0DFuHerSS3kk2ovEdm4dULoaqOs9i1S+PBTpA7453fvSpXeCaeCfix2Gy
qtS3VobX0xek1h1vuq1IvneFXiJLattsbJhQZgm6B4NsbAwUFycLOAR+9AMblLj3
6hGZfHw0Z2x0jejEKwniDu/ej3WNlJV01CNpk8bR0+/o9YfJIV7XFny0SRmvBVyy
y96mNEqA/UKFUfDh1qd1p87JRKl9j77dBsZzK+MEx2wSj0PxghuEyfU6ndUl0p2e
/5du8Owj9G8ISseFd7th1UHeziRrjl1GsDKfEpmKMEPSiesxMiQq+8hW4eBnR+dz
fHYrFkygwlLML0QIbF7C9PTcyncXME3x/0wlJq+GWEzeXN2mAG6LaDpPQ8MSQ68Y
XJ3lub+h9ew1fT9DzOxYwNIg7MzLi6zZ7ebrh6IVogum8d+5PN4sz+Alkcd8NjPn
9ajR50E15ThnMkG0joRcZasljY/v5HkbSMNL1lCyzMxHX/VEbnsVD1WLg5vxYdyx
t3LTe/4jgwCQdddEHx8xb6mm/w8jhX3rHRgNuo40p2cRceJ0qD3lrHRKTG63RyM6
sxHLOppRNRD8ZEcFQ0Dsnrdn36d/vPTBMq8+WNc2Y9L18k1D/t4D7F1O29CJQ+o+
QyrAYyLcyIY2KnD0IaMoZy55VJagVvnOp+uilDsnoviY+nkqbLIrG+NdCuz+R4wR
Ac8SMJky5YpHBwjcScdJkmbqBR6VeFf52+nxGFzAiaNukbwxiILtfaRAqTLDRVi6
uOWZEcpaDF0H42vdYqFjdPTLa5dREnjbgEJe4R/hdTkSSm8/fI7tvnIwkHY5W/6i
s1nQncpTlZp9059IcjJQ/CxFPCKiPC1Yn7anNwc5UPywId23PU3M29ktbx3YmYAy
3/FYQTUx6dcr4y8J7I3hsPkdT/2M8efEf3XUEscz24hBhUjnp60/WCUJlEy31Y9B
60XO7BRoFU6laoSN81wt4+1+zZKIY5H1QLm1cd2f6B3EG9D/bwmvwS3RQSF7KYur
EMQWeDC8C/AF+s1D1qeIDmlO3C1DwGHKjHe/PBQoGAfrLQeWhdvdkNC9SUMtP6m6
d7tbWgW5QYIawYKOvxnmr6j3SZcwTbxdCJ6PYxwbcLzxfpf/nMoQUKqrTqxRsJ5Q
QZjJhfS0OKHGOTYfrUKyv+b50ALj8I5dexIwxxkO04FYKysV0Ru/BDOqRHo8/DyC
8C3AKBkpTWKr3j6pZBkumXXtwewlI5GYOxUfVkxeE96ShMXaQQ+oVjbe6H1rY+R5
5441gIwbYxa3B/pVA7G/EVCZuFhEpf8H1hU0lxbj1h41nV5AfrugOGQDdvXXLgG2
YqSrN7fkwbzKs4KbZ6GZL40mDKjiKXPghzvztyrp2tM4beGOIpAGhOMS0v1JeQPS
hdCTsJZNIIuj42jHRS84nbzMAu3NaZC19pqoaReYcGA55KUi0L/PKoYwntd9bmZu
VbJFu70SfKJhyde/4qP341Xs92DROIlBPqHIxysPMM8mBX3wKgcGIxh9jumK33F9
pQlnXg/+W+BaXyLaloMcb8fTlXDNlMYRk7jILrWRaYb3Ys/rgtzJNW2EBFWA96i8
XzwfQL6pyQdHyvnu95f73gH2bj3OQJDNuwj2mPk2wuPSjWuI9EjyJXCIbv/ZcD/O
dTl0gVn75g76FEcmbzxqGcT33o0yipoRYUkUbXgRd3AztX7RbAs7RqR4UyAi1xEK
huKUO1AzyXSqmf/SYgRare9/1MI+1a0olLqIw0OyY3gZT2/B+JuOrgr1Mo5zLCwf
449sL/ajpfKbHauPKrGA/C7sBZcl1L0Oqoiijq/u4MLefbf4UOjeVzgvual+O+1/
xdflIzGQ5K6RRt0VQ2nIVRGAiXifnjnVwRWysPC28DZziUIXFJhNTs+UEK/PHIos
IPNUEHuUhMf7F6rOc9J6Agizu7DAgvbSv8lmb9DaeBwzvOyH/KG2hYQefRn/D8z+
pBPyfd37rrVTJCdn7izBcwDRvk6S/agiIC2Hq0pJMVfRHKpAVHSetI2qU7q3CgNl
fB4ZxpwGw/7K2q0KZOOGzs5O5IA44R3RF4fPutYnOPRb/dLDXEI4PQGCRqq3REDz
+cadOZv+SB2wyzU87rOBmMvMrmTxhXE4wZcMSWc3A33BnEDTnupmjNwEdJzsvPCF
eN3ZmG7QgnYsBiekI0cA2DFWs/ssPDkWYnkgStav3S/F82dvMsTAmFjtEzeY2NCH
dnwgyUwycSD5uNobSRyuhyfd8kb5xMtjZxOZeIUglRNMOnr+b5hKrcYHM6i1yqxQ
ICInloPz19FBdzaWKAOIX+V8eN/S35Q0CB9r/bcK38JHNWfpVawut/2sqMHtgCy/
kVgo6GiynyUOH1Js2grFHTFKhdWhV2ddoMG6pXKZ0IzDdMWLokRoarUBIl5dOHIW
fG+RG+qvbWUCZKBST8QKvsRYhTy12FlHrBbvcCTHzHTLvCjX3hKlHY6593lp2tX1
7LSPBOOAT98C+qWUcyQlCR75UCKGoozAg8b98Arb66q8If4znZfVwLSUU8LoRfLo
ftq5XFQuck9viW7/G6cHrtBOd77PEF2lYGzRUYSBJFhRNSIIrR4L6IbJzSgEzIiL
5wfAoVop6QkdXJvvw/gYEe3HYYwAjzJO6GmcqPjWNOlMgCToGiuPwxste+fUPXEv
AbPp3kTvUZYmu2m2Xi2Ys7HrRSmfedXvAM3uQ2hkzFM1/E7dA83RGvlV6ek1VMVT
hvC4iGW4k9bfI+Du88XabhuGaU1rBlP/Z//ujy/WQcT0/EF6x4kINxFcvKHcroYX
KI9V5pEc9dgsRUNyZZhwiEsqYfGuNaWoUXFPtEo5u8loKA21BCJcKbUI8tQ6BABY
hDAfB+FjzKtwhcKjRt0Y2LDdpPBtVaVWDw6gA8MZhQYVBejublVjk+d9f9GI7e09
R3DpA7CAZ2+zaulBXi2e6HNEVSVCrrTtucXklyLJ0sGMZK38/T03NUoP/LK7AZAl
3TOUYSqqtmmzMseuJ8eH3RLjdOYnkAbC/7e17V24PRbTo7c83UANHalyO2ttEeE8
VONix6Q7pnVIYkaMcRgjL56iNDQkjoIlzeqHeowrmEQX+RV6zvoX0qhTXOHNzaj0
7Ipmd6GLGKY04eTocy+nnggWDXuOHMzsE/IQhlOPcnEsf6GVMvWczzTivbaoil7n
Cb0OLx1YtveGCd/m4xPpi6t1wU5NJJX/HAwyULtRd2sjArCYqNhClAsMYZdyLDrX
JBm6RkuSQ8KEMa1gcIfZ0E9hHATT8e+BuqCgplUa9oF9RxqSqrO7UqM0/+kJh2Zy
+98m/hrHk1w6cqCycZp2K/FYN0qwoos65TE18XpVXtcUerAzWLwkmLO2TqaaNLj9
ewnqurB86IZBjiHZYd3e4IyfVIbG2ulqGmCucZ4VS7Pc3cuI2VcMKc6yo08xXGum
siO6fqn0GKnDF5ukeg8Tfag8oXLqmrJJLV6BYwz4spBoTH+H2msDiNDTHzOFMwoT
oO4biyu9fqUBQzB2OaDpPz6l1zvK6rMYxmp7cH2Q/SQzToDqprI4qaYEG3arfk93
lXBawS4bTUlWIiBBK3BiWEKLh/5xhmqVaaTmg0b5EetOa8DCaTNMiVCmRpvxtnfE
SShJFNnhPuDNtwdBfw72H824h7BFJVmiR/wsAtXgSXBRNh/WCyPDdE0mFvUszASI
aHwWqLp2l01jMXzKn4qeedoB440AUsBxNwtW6gNRoJjSGjF6otXCjsrKjXQysdAe
ZTCdHhW8As/Dzerg4ZWOgU44JP9jGKGO3hsVHqLtDPZ0FqVgistM5yt2KcpoqRem
Hq+lenj27TC8SJGtjJx1RSIA+y9VGMtFHwmZbhOLwnO0gV3m54XZqCFgK7O4UBai
bhH7b0hRB7A8D2mH4ECgi+7G1LJFno2Son2w8jGXdKLFp8NwKJRbgE8EUmy96m+m
sXphKO0IKYV1eIycyY7XGqaklalY3EGbzC+hqpOT1uQsEdblPr1+Vu2dpe8Lmvzr
Gw9/bY3s8s52eH/F9ScmYDvHkC2s0g+O/z1G9xTNKeZfnhcQPR3DHe/Qd4N3Oefd
WzvmvprzrrQMybISqowoNmyxIFfc2hAw/zWNNxuC+Drch1Nu/55b/RwdPx/EVnlA
EWF8T/FvoZq9FXk7tQh6g7y/Rx5jZ9bTZG5Ct/XnMiLwiUHZcF6rBpXztLr6vuTT
ybR0Dq3KOEDOTVogOpACxqWYPHye+t9r3CLX5ub6BWY2O7gaxo4ciVRPfFqRgDkZ
bARzxn1jTZdFKUg81A+8SytnRL+J84YRH+cjZoJivSFyywaHcnTnd4/h54Vde0b6
VSAdbZZ4CoGdUmtylLbwRN6TJDTbCKla30B6QqvPe4m/l22sUbDssNVMhaa8VrB4
sn6OGMSYFu08hmGjN1GAsvwQ1FN9O+jEFtsKIX6h5LajxbZFl1/TGb4/VRCum0OF
fc27CqF+Pr7ZHyfgvLT2C+Pje7FLimUXua8wXczPeDkZJ14RCNnNArB/kXMHgeHQ
Xkze9BCRyNf/n1ySJlD9o1N3sEaByZdmj36tnHJYAy01k9N/gy/WQPty1PJp2XXj
8KrU+Ma/0R0fT388D6rW1q09PAW+FV4Kbiyd73uuyxBZiTi1wy6zL/EL38+dMlR/
vbvTxr31IcfdDgHjlnxxIxwZowwTw2beMA28PPGsCzdVeQ6WWfKZ3XXzvyqp+kVO
Prxgwwm/Cjho+cVy3Qv79ihuUNHoF1xX3QYFeMzpZrRa9tG9jIBuEvm6bT6YQaU1
l2oLD8XJiGeKuJ8R4pAlh6EXTghz2R/ig37DWcKfldk6PcwmcpcZGooJzcGdb25Y
ZtdRatw5CaAmE6ChbnIvxHVFUA/FcrOlYZDKhwQRPfxWpZYUkdvBTG5KhwqOerkX
6/vJnIDLQdn3jCk0B48fPvxZz0Aj/f0rpkFmKSOcpPOoFGPu6BcvOdF1pCictY62
jgfwUAf+KsqgFjf7hukjDWPK+SP1vb1pxr7SplColeZN9FN5OmgYL+tSoe1RU02u
54OMUyACgS2pyqM+Qh3bF4l8d6AfdAv70CxMoLMiVjSVte8J0wyPG1pUzzXDNWNv
jz6/s20Ft5wzqp9DWDwEPLbGco383i+paR+hwJpzrG+s0eGkKSzVV8nAJ80bsUVd
NXxTynj4c54Wy1tVMb3dD3KmA76w8VmV/5erarkm9tINtEThrZSpGSEKMnFePHOl
nZXezHAWmJdgjt5gqeN40eADg2deQSJxad7nrwzE50CIfkweTfo4u5SGtak+xI+C
9IQsfLPmUT6GQz88Wx5YCFtByMGgLnUVjf3hDkhzDPWkOv1QyNptwRV6AZD83fbd
QSqqNW5VRXPfQ6QPEyZsfjLhgMYE36rNWKmm3P1OqC2uLNj8LNmfTpiqFo6tkpHf
pAbtYTmDv6IHJN9PMl9MNbx9Ut4SgOCQp6RgY5s1LCS8JaOXRSqniBLoj9S2Ujky
CqqIgTZArbu6X+bg7U0xWRNpRasNPzhikv7PPv3OVbrwmnGAsmtjHQGlRiD7jV2e
I4YR7f7XrYLeSt1Phxw+8DkLXmiXh1yWjJ5IbcMZBGqfbhSVo6cTNJr+5fnyEIJh
XdIy4gif/Nvk4Qvk7WrE0esNZesgW21QqZ+q1KABs+JcUDt/9QZHbMnBILaeikwq
NKAIhPPtF886P1KraYXKmT16z+z5HE9Ag471wviqNvwUrHABNvfAvmyKNZMXf8n9
P3LtVFH9/dlrn7XzJahBZEzubDKwByiwbe8skHY/Umxn3HmSDZd2UMr8kpai9ed0
akgS9GBJAZzRXb66xCtVvDB6NADdstDJN+hV/ZXgEhcUaWZX+IlVMg21y0fl6LIQ
gukF5eA8xQAmovEZdYsV4J+Ub9nzMTNg8CR1GR8rTzToul1nliXZUn20mKsztizx
YzY7hpt5lAHvcE6FuaWp24NNNhPjHJp7N9bALfmhHF70ZXh/K7T//3G2WZdJyfyc
fD6S3MYjoxQTYE/GicqNKZkqJuHI3eAM9xPXG53Z30YUhCOxgYAGw/GWf07wBWDb
1ulFWUCLCuz24PFP+NWW+LfghrSD3+PnUjFovgY5EDXQBVUjbUJfCDiCpRUf7ndS
PZkkWLneLwW5ZVdRsxmjea5QRV5l789UDivpgrttbHSHrYXsE/vvDZdWqPoDqgYl
iI65A+s4rsYgWhQGHFLgoftDegVLuzdatQ6VTlmQU4CzFtS91l7n/KHUg21SR7Fi
/54X82YNDqScxJ5ReviWaV9ObjnORNveDFo9gC7oQjffucTZnj3D8w/1p0jeOJVB
fhrgNFDVj3hsMsOtMIVfIQu23+bgz1op28DppfTyjtE09ODcdyNKFWX9VBvKKeXx
HhduH9vp2F4rnbRhDMmGzcm3uLuBHgBp55dnpu1A9lI02OvbNaPjfV5Yznsq/XaZ
Dok/t/UhPrPA1pAZkWToH7mAkjs6JkWNBt9Jz57SLuiVvNMvOv91Y9Gd+YmVMfiu
QdtanWul6HN+XQAT6iU26Awpy9XqLvAFcUPOmi4R9j7vMmJ0oB7gamg4QmlMabLe
GPpJWceEGxzviGlSxudBPTU8uLg/pdU9fGY6m1yQ215mDV0ZKlJbJBCMr2iyp6qf
ETWc8s5ShQl6J02EyuetyEdnb8baowfpFxD1rPYb8lFoI4n+rFFrW/862vCrDtNu
vWWp+dmsJ4jwwYNtvKDAoZ31bEHdDwzDV8HXXOX+XtaefxeBItrz/4cb+fadmBbN
cY4kBCvO2XWb3GEwAcZN4f6f2GWKFHZ8g0jmVxsLrZe7W7mdX/DOSyLDy4yiirPC
xRtG1IB8ImFQKor4UleTF11A/Cx2nA93SblZRx+gYIi5VdCIyN3MLMRQv0QwaDdL
4RTVqVJJUe90Sgw8YMW/+MGLZClBQO0vK9VU7W1uiE5kEe8yALgXn/9uLgu7OE7A
UGSypyIlyon+FbH4C4lOVAOo12QFpcO9CcUvYyIzCC3nNobrTeO1V4PyE2AU2JC3
EEQL/gCnXYVp/T8973NrKKXG9yBTRpa0XiZ7HYfN1Tg5vFgvH52Agc1if8vaPbdR
N10m2oYaDgUUKTpiXPp5R4pnt1XHGmNZZzl+jXeQQGK1tYa+vWRvkefbgheVepe7
poPSfruGy8UAnCOHHxg8887lVQSWgd528j7xiXHB32zbcYruIyj+6XpJVyoYSOP2
+YIdfXQmL9Jqz7Z1NyM8Wk/tObPCuDp7bjndM1XhNCnYMer0OBa9GqVOMSYyW+Il
X7+i5z1pmkNCv1iTbZZ9sz9bNRo56fxAE+1ZhNP/sfK5n8HnNlWD+8+/Fjs596oV
jZAelD/hdlN8XaSyu686U582Br5mdnxrS5lP7oDGAiMviESyFPI2WCXlWZqSjf4R
rIpUrL+ax3VFgYyImYr2jS2ydzhBTOBuj2bRkgLiquK0uLlVx9iGXujTFkTSbed3
cFSJfoq9D73d6qi68u0AqYjRm1UXrCJZu/4yxmHbW7tBIaY+Fak9oT81POWLnFHW
eTmcw/YntDq/qNEZgHu2vO9SD4/CLrSA/HRwCFwhuVl2Bac/ZiLac0pw9uOQkMsC
H0eiCfhtIGLjS99GZrFlrZYfSjAdf8iHGdqhE8Aq5QOuc1rXzYd4xaEfwd7oCXED
yhlkC3bRpcHLM4AlSwQWUnGUBovFj6COSMg4/STbj9cII/HkC60jYPYeHE1SXIt3
5OKCax/XFmtVWBnQkUpBaSCLYBwCmbJwcUQ3Ff8lxK2ny74nyPYZQK9G1SCvi3cZ
AmslD/iuB6MV4/ZXYEnYerxFug5vBqC7L02ObFOugK3yvJce9JJEczYPRarDGfAt
E+GRXmkh+FhuEmU48KE+gUJGB6I49EWoTQQeQQPsX88cfKuWh3us2CfVdtMpNfyW
lu1xMODdy1BG8xl0+jEA645LEIvqDsaQbu5XsY7frwbfxwpvoiHkXeB1JYyJv0Ks
klg+bZfEa41y7+yBAjhn6kiZa0JE7cWzUsUo79A8PeFWJOroI7KjBOnOCNHXKcei
hx+Q2IUi7tszXwpCMkiu02jMXLnHSPKXO3Om+s+MZeh++FDsD7uooSjiDa1j5QaM
AYfNC4b4eDIWSp18bg19MBJBfs3a48BgZ3fNRA1VhtQiNa1FW4BToSTG1Ys6IhIR
mMvZpT47tnwJC6hLN3IGCxU9ZQNci95kxfR4iIZdPDqQFiLPUx4sLpHQmfXIZSGE
Vnl1q7QafpBUZYHkhvfERpsZLv+5u7F+1X3R0KJ7tkBf6r6fdaNgB7MSsEORv35+
uMota54W9JgPXWiMwtCCYXHyq2LMiCcRCGaga+0ICN8EGIGsLAXsf8a0xmW+dXZO
h88vG7xYIIecwHenCb7aWgE9yLhgM2EVcOXMA4ugg1dnubXUxJmAs77X9ynKNZnd
omC8CMltYvAYh7wMEvlzH2mMlhalBETTWF9FVzGKj9vPLZThwbwWDZdzI/p6rt+O
yI4/Sb8cOw1p/S3/bZ4GlLX0nEFaykYyjcyVmbDYz3gjVknEJIwGkVrTGeYfXyMg
1+tHWTGo4HNTMJHuRXi0m8PMH/sH0dpZMEKYjx2fjI/zUEG7T23UXPXKCdSaM4oM
2HnRbZO6ktdjIJ4u/1v+9Mo2vN9FX2iMr6FkqbMACPTkv/C+Mb8SGn6iNd2Hp/Ia
ZUB9Z7G4CKQ81Jcap/s+KK2oOlYWyHPlmnQOr0Ot6ppRyCB7HGk4wudrTHSvTuxi
77RrLzfaGX1O/j7Lm3gFLy/AIUW/90QoPfrI3WaYImOkToNqnGNKclm017PAaeWi
FWhnOc6o8CWOyxt6/RuXlLkkk7JDM9rHJXRV49wZ6aS3T49EJ8DB+vALnAqOYqah
qbhtGC5AfHDqptIPRkEaiT+L16Q8VktDTjtQ2b93NZ4ZhMdj5myba1PFwcOgR6jJ
36gIPIOY1YKNXOToXdGOhXW8d2a4XJd+8h5NdjznlXoVLbmbxftgMSpDOduMcxk+
JimwK5E5eF7maLjhVjm/66WhoY3RJlskyK06RJt80yoENR+14cP4/hN5N/Z74zwo
Tl4rjhVC5bdDWbWz+18BeffsMHC5t3IjnnQjMxOeIT49pLxCq9Ss9QfkOTG5yCTq
tGoSKIYPMkFKHITOahClQQ0wzOSAvHze3AJzdIRoQU19JZkch0hCPVU/ggbjUbjS
uqkXHM5Xhy4hY+xXe4j86FTYZjLJ5OqV8nIllZOvQL4bVWapoDn5fO9lcUWmL8C2
9+csW/vhHAN7Y00A+WATsRWXgdis6AaSJCWEdjpNidC9WzSzxFQZrHnD6c+qPp0k
M0PMq7rpLu3r9LsjtQjj85dMMgK3Y8k6f52zlhiwg9I3/nmTpx9suYMpacE+S+NS
WzpBKRTQhS+gagNVHgENLDW7A4fbXbYPM1IMVj6JVE8pDZJaO6yu3aeNEDbjyVX4
iZsu2YBjT4aYBiSQtythJbv1oqAbcJis683Dc880fCHCyeDBchWYncRHW9ooh7HG
QnWOHeYpOjQ8o7TpA9ZtbUTOE7e7vi8YigmTuEn8uJVnY2GARE+IFooNBpeR+vtu
dy6bBVeJQuwxL/7tEYkExsiFk5wCGirWoZnE3kOW4i4QA4stCJtH0gDnlsu4nW5P
M5uNI2HTeAJ9h0N8s+xaD5LwDvwgdbGOou3QPVSNDNs6AfT0gCeI4BCgttLdXert
VIwFqhPE7+2D6ZOmtmUNURd7MJZelqTtij9LIr3fUhGMDw3n5R8/Vul3MFEpLh+a
qhMUOr1tGviuvrQ+asBN5TJu+IkW3S6Wnr9HPb+4LOpymA12skAI3yWwQfE5w0XE
pgBZLbUog5qUR/7VJyoibjK+Culvm4S4DPr6IKJ4TAkvyJE6wEfm7PnoXKeHkIOG
tvhthv/ajtAruS9ec5DQSEE+yXAZz/poL2EblYvIEfC1pcyGBQ+HZzkWRHX8Ym3j
GYRmLwsvEnhqPE01pg5gkjJFJbLFwtuCBz0IEkW013wx++rvi5mv0UvfSt4p3LCC
dEl+FzlCYIdF6cuywthPX3BH8iC9YsTV3P8PghRDOtibxQ/LCaLJel0nZPTv+Epb
AjQjNH8SKwdoGwoZpmahvWih+vqnvYCOI1U2DZ8UF3eT0+fAiUoNxU7jezfkvBGO
vnM3DAKdBZR9bJGYmqXX/VcAgoQ6XPu/leamjE/4EXPu/r5KCX0M7BSSoogj7wMb
YoyHsNdwpoSx7f9PJ0GZKCAxbF2hVZqUPGJjwVRT8eAvtelMOcOe4mFa24wowt9b
lIGObx+WLx/P+rU6tQBniRpOSOLfZ5iJrSsVFtjsrJX0/IABpte3gX3mgcr6O69/
1PlpdwoQBDO4+2KDzi6ZCtahU2gTCEGfDkwu4UTYHBp6Iem7tdFQa9kjp/KO2wG/
4lDDp4pgft4XNQpIRmivtDg+6IT0X5vyzUuY2omWta5lvh4ceZvyFi3s/hdBTXnG
nijCI5IB9T7NdlAbbJe31Qq35MyxuZ/EYaKkD4J9kGLaAj75KXSt43y48O8DFW7L
usPJ8YT6dwq7caTNsKdCHkyxK/6F+xfpHhklQXhVYaAcCGOEp6P3nnshWGIUPeG+
bW7ZlHvwjzSYUy/B2CD+lEzZqDsJykStEd3DzCKNPOq7mtaK1KCe2o54TlHAOh9x
QDP+W/WTxwu9b3Qqs4wZt28BK+BhsrXqTCIIcdaqiE+8JEWBs6DakmvdYjA9en6L
vaQCCG2c6qHRbzfjSHkzO1HkZ3+MjkR/0/ZdbRGdZ25kWRczBKxixujwri+3hmA9
jQ4dBCO5dSni7B56iXv695eLBcSEBqbBgO1zxNMeM7SAYFTiaeceA9zhxnRstG+c
X2mXnq05d9l4p84nxcE2rDocpUHyIZ+2/io2gfbF/gZPl/EYGfHrsFAZ/KzAnWDe
ByHbwX8yOFU3Oir2S5APMcU70dpf00B/6igy1WSdmGqNwitm2vpxm9VonAlVTQj5
YqO76f2Qq4x6O1/8mIElrx0UVpL3WBUzRjNdwb+2pqrsi+UkQAJdjVXR192qlV8l
fjvd/9wOTis8akQiFOEAskzrngCPotLrVRnUGAr3X8qPdWTUeYbL0XvA0kq6sIwU
6qVldZjyiXbvlyWLEzkc3j/ap+PWViLQtBWgcVizUNBwftcEVEjTsxy5WNYT7RZx
xAV2+g5Fww+4+GEZrDvkcuzofCl3pOhkIXnfL3W/I32742Dcy3Cl4Bx7OaN+HPmv
4ambkyYGQLgS6Tq52BApzTm5WHrJzAxd5t/lUajtcCuNR/rUg5WE/ZEHsmiLxMLU
3iEi9aAgfmXfRNWOFwLUwr3/MMWufEDYBuKm1lXsNfX0LEVBue04AzYOK3Ndtwjc
8R2FFDJ+5128rWyzHdTneXSC5ix67Gtj9zkduGA7VSYAKK6DR/0aoeAbJFyxRJ4+
C8v6+KHzwpMmeMlf5pp61OM2mf7s9pY/WE4KY1jwFD4Sxb7DwENpxUSeeN/4pEzV
mCp5GeRE+WX0Vqpn+Y3NQB7xhP4kXJ6ju5ifb3XesB6/ZkSEmYkksgK15FE2v2ps
ppmKcuCpY76rMBZDNPC+Fa0LpWh2pgFLPYKPqYhIdeUGVnXCpjn3PZqgKSo6eiqo
TUD4tP5m4cn2oHWk9Iy3DXhBrZcfgZny9n1tzOjaTlrTZt9OmERcAUqaB4wwopmi
9IKMYraInN8PlYkqsPdHIMrCCwVKApG/wUibkUoSXVyzvez14+Qai7ZomME7QwZR
jfJv2b53GS8dlf7WJ8IMg62/19WqYA6XSl13culdbWhPxitthj9i5dQEtDR4kf9u
4B3DaMBJhKcOqMoHVqFl57Pmy4PkPuOZDTLynK60DcyagTMWaQvElcLhb7aiMz9o
syUS46rlPsQexo//S5ipcuWk87Lz5KxmEAWApGlN0PWvZ/OmLgPhoirGdnfTIYjB
zMUyRMBaItL0dD52lGGzW/zqnU+JLAjPcGgkqguFwZGFP4QZF9W7/yEtQnRazIV7
rBcU18PtUjZH74VfbETcIfyH2fd37SA79X94w7GlyGc0D6suYa6BNdWlRUyx4JZ5
Ju54tA/NmaGf3SwXMnjoSeZ9K+CtNdKJkwwEnSCM8qaimg4aTEqfv8uF1EVFv9vh
0ZRROghDFG4Zx2bonDza4dY+6oICipGHJ1HezLqPFTcz1ls1B/vWb8YVeeDyiup+
8KbJeCwN4HrZ6woRzRMneEi73bhREkuxpjHpKdYyYXyEwm4rb5qkM/tCylF2LW4B
04/kNpKmHz18pxIEjazjl5cYboAsXJLBuN3dnhmCJldeTqJ/I+Drt3hP06LOGXpX
2kBa8uCaFmzUT+9+M+A2wgULfwbhmqelyHlIVF5SmN0MLANDgFWnjSNTY4fNERxU
bwi0tT0L4SUKoWL0nhHEoLcsLo2EqF7SP6bNGOCc0movqTB44d0nXJqUuq/ktpo/
FVnDI221duv2GP1bdHDgg62fHuDmTpxYyXaRP6nwI8qFOGTCILQOi+EtDNh2fUaH
hoSIt8sT3K6gfJkDw6yiDI0bpArgCrt0xUPhW4Kb2lZ3YrgZj/LMY8QKCzfPIja1
nQST6nybBrLsuHMwhHKZEviWdf1HKa9edRokcufwhCCmT0YHFespC4rM8GJHkd+S
qnDsiUeK0WI74k2aMT54ZzGFDlgZ+2cCiun0H2Dpd8VV88RLvI1wt2qFRfjKHIFZ
U8H/hnWN45PjZTm9QeQi39PpNENft7ijzN5yirFOACqEG/irm33R3TRRZr+9qlEj
uV6sGolGjXOB20pR6no5XS9yaXffFgcNrHvMOxHPkytVFkuNlatQGkqI0+wKZx+F
ZAtCG/nDgCUhrbIrytG0ZZPx2WdgYETDmpPBpagTVnFC7wBtPDFq909MSRTlrS5H
zENn8GVPyDT1luKvOdBfDoCNKB+qrrr7s9yn1IOr5l8b9hwNUcorelHl35dAmijh
l1c4QT6vsBsKmFjJ9cUMgCsM1Khiz/RUv1QoQcYHpn5ZG3ReDvujTu6WQx/UqtHo
rpbMSgUXpvJjfyD836/XFwzTDeVvWlVtnqcpv+CupmAKloGv2+/yjDTaHUFDslNw
NguCzlIN+/q9gEUaw+jt6lf9f0o+zBpEzJggZ2nhHk9+UAAcjwzmpglDkwrbKat/
bpzhm30CStw4sfaFvgNFNFS1n3clsdZPl+TSNXwJClloLZGFXFIxI6FBxSNkYIc6
C7UixJWwWZFwLIz7lYjzdmDnQAbvQIgGt8bhaAJY69sM8yiaWXtqEqtpn1ePKZOw
/FsMIFjowPdkhs1ZdoCa8gqwFhByRrE6Dg2kBAxYnUw3Wbaa9vaQvw4JooZITDrh
apRMRemiIMd19Be9mT1T7iuLsdh+py1FSRHp1zU6XIGId6Nduemp0yyLVKyeYtfW
wWTRR9uwSIF47nGz5+3QJ532hDJsZNXR7YCLD1EL3vWureSQcGw1y+6DJ8LsCBn/
vMZa1vuBMuydNu/AC+oK/1Bm7Vbj8rJaoXsTgMxDNOmGWa2e1i5Xsx/r4ZZWh8oI
A/GY4qO1W3ZxCdnMaZFamzdfuckZ9tIuu2SYiV/HVmYkHbvL4PFx+iB4h+XBkA9/
5V/Hay7A0Orn/+5dWIzq0Tm+cYi3lDfEENYpngmI3LiumPq4n9Al5eu/Esb2BArK
IQJZtJ4cau7BEPPyTnZ9nvNMFWRN7nITeHG8wFXMICfPI2R2xceP/Af8cP8VtPKa
JdBy/NPTcT26hPnIcoyNSHat2jiglqs+3a7mfibSZmtfeCJov6MGAg36pHEQogq5
31dvYebzoZwD+867CjuzTE6ePEL4vuJy8ZL1uf1zLc+uYRA1S3rN9jobbCuuysIX
H8+9BrrWBvEaKRRvdEmaHTHaP3od32kb4XqJJ0HA0xwK3UDEfTBCSjuAFmq9R3K2
gdQpyKEn2wDMLjlUYnWuIrRDBpZdMpF9RPMeGl/EvhNfnRNId3tU4OToaDEX8vwW
kgNwBow++c486k0OkwtKkWogA6233tY9tbUC6xz2F/N/rtcHXS5v1zgEHWWylL6T
c27r63isoACjL4ff67CvMyNQKEcBhI9UYOEws07kQt5IcAZUfC4hOjQ5+dLaIkXe
Qw5Unz3PhFfX8jCUBXpUENVVAbNLmzjNvWhgFKc9yVG8fxMcwjU+rLmaHZXjeakc
W/PZTPQrm8G5pQ+Ji6b2n0Y409dTWiVaa3KYjgCVL91TL8rZU9Tv8OtzBAwcDzr6
8yI6o4S8/NAg0l6x19+42wfxKWDjSCyfnnJZ/WapC+sqfyHpxE99SyjQp6ne2lBK
8Hz5EIFOjG4/aS31zqPsSH3Q1xl/ccUHIp21mAVh+PyKm8dc2/FePK+JkQY3h5hs
Y++OveKjfV6SzDC7Y6OQKqVWp+5TRRtHm//PBEY2JW3NgJvDYkKnAZBP8A2tKgCn
IRw/oSqCerbSJ9InRPPensf6IjmX166Fkxc4qOdcrpVfVOAttionkZpdOoXobquq
MRe16ovlGOT/a6+UB1usEFfQtUzFEGvV9sKIeEscjQqdHydWIzR0aDl2YsacecUU
3u88/ihXyfMLoKfNYg+HzewiVafpLIA9NMG8OEGy3TVM7HLjMzkO2/Q4VlajQb8W
siGoRqmnJRuE/MyEFNmXbmQQsstqNLcBa9MQ4YBFz/VzZKsNxBpTwYY64Mu+hg1F
gjs+uUxLdL3YtvJ7F0ZX1wHIbeBXF1AYeYHmTwhxbxMz/fnHSQo4X3d9R6uze3W9
dnNhO5I9iFUNPLIKUFbXgddkwVJdwQN5BB+4ywmEqGaV5tEgetY8oqBq+koPL+7p
tzlaPBSdvRDJOGo4bMKUGq+3k7xGmmEhtFYn7TIqR32QcspqZAcZBf0pValc0XtB
yQOMLwFJgVl0gjI+2O5jg86U26Jx7NsBLaZCny1zFJXFu0K3U3y+nYttLeE4ffyE
4DlF1bpxm9GS96YsyRCmnoUCT80CPi3b/gpBfzjMu8lau3T6h/YDXlrbd5Q48Edt
QIKu6f8blyJCrqr9mXgQ2uTwsq9rAgiCcc1y2LM7ZatDtdlfllnBN7zAu5CT9CvI
GDCwepVYOpOXfO357StvMQRpz6QuW+9hwNIuXCdtkppbDZHK8GK5RRFhYT6pOGlK
FUnpFSrXAWg7i4OETh2oowG3gJxG06WbLulR9/Mt+RdRfyA8lxk/NXVkGSZBxT3F
Npx6Z0j0fKtIcPQLWkDwFh/2h28fcxj8cYr+4l/QPdIbezzxhKRMw+YYuXKX+6ls
pYTK2TeN1uougWyPNxQzIoJh0BEHGpnrjJXTa/Nk6VXRg0SvpuIMh3hN+TJsHG31
pAsX3FYwAxs9tM3PxQi+AKley2Rn0o8H+CEW7pI1Y0dDuQZ6F/bOIoknb46ubLmE
AmhGSv4kaDLYQmJXqZZxw/OgdfOXwiFPr2tzEnwIx2r8rwJ7NK1iTmW5DYSm/7Wg
pxWMyG+tIO+wkx6G6q1C7Sv2o47GlE++FETL0t13Ogu5eScBIdqMqXF4M9W4qK0A
O2BvXKbxwx9TBwmo79uqpLD5v+kGGBO0eJIJSPoiXB52szsKTtcE6cr+T8CMCw/N
TvL5gXpa8ZTI+c6GYGc/3FOlyY+E3rrsvr/N5OoOZ5uRWUjNIkh04jjeU7wNRAs+
IYzNM2rU6nBFAiJYdTwCX+VmroUPKp1RxAKsnEyyrTcsLGG8gkqUNja/nXSh8/59
mG7Dzrv2ax9FlkZ8NMeJ/Q3gnHnU2fx6DQPQFkpSC5Id0GhNYXF5MXOqLPXHFAM6
47VvP5YYc7hk8nhEsMGV0HK9EmLmCLlhlqL9dkCbKRU2nxylAs7CdaJWNySD5Czi
gb+POTiZyJYwzcFO8hXp7otBGk2+wF7ZFJqGG0Yb8bPm7sgvxFq8qMfQPU7erApk
98L1K+apfHvV8WZrxEVlawEqmJiH6M3I4HlHk3H6dv/ttyqIv8i+Q2eEsmzG4pF9
jOU9jhrxSFxiOteV70k06dPDlPPN9bstsXAb4PB7AI9sTtse7RLr44Z7FG0eG03l
z7DUrnuFK9llvgEYnfGAKct5di4EUb7SouL8VkCCGkREuUjGy32d5yZLIKVCsuvF
SxPRzefAOuck5g4Fg8UkIW0neAe/yAEAZvsPN+bcHD+5PFhP82v0KIfEl3WtcZnU
4XwysD5VhOzubF1Sw2QpZnXyTFDUsoQQk/pK4xl98T12jER9s8CegddnNGvJYjmj
lEitSbBGDLfDVvvCAFg0r70qSEzCGaD21cLHU2K1OQNz+0Z1snQrUI/fgLFFNp9u
Zi5IJbV3SLJsl53JODsdqF4oqo/BaWBKX6dNJlOgj49DEwIQA2hE+yaDgOEzvoke
iiNgi2iW+5/c/NidmngrZ9MEzBkZTKV65njiyWOvicfEB13MgoTFZP9BN/Zvsz6q
/ap1kdPjZk1demH8rUEjA3TZ0+k9LyqtmnYDlxUEPGh25qexVFzM7F1/bx9T7tAF
Stidy2+78xxaMnKAEC1aJlafjBCW5HZ10fjXZHET3U2AcmL9KT+YVGdhvGBtvwwn
K10ykJhgZoBKVuXmOt2+IBAnVhx7B/wbgXM7zfzwGlJbaY/IDaah1q6TYWbPfW5p
oI6ojZhRsr9KZFuz2ZOQ5O6AgY2e+jvbJiR3hiRPrNQf9Hyylo0lQbM/N8HhP+Cv
AEv0j09lrmdwgXj07qni9LAtlSah6IhulckJDRrdsmwKECbMK8y7RP8Xb2T1/R0N
KU3dUOyJ3BBb5cbptH94VkMsstuzC5ZGwDFycLzX6egfH4lepZOBMMzvF/Q0nGYH
IznwXJ8LTLaTjD0zQ0ylABLh6ItMtZHfBKdRdTiItwvG5dnD6zrYDH4wdE8Cmmx6
svF9cPOLccuZOdrzuuAin35vCyF4qj9wVyub1cSYkpyDGCv5uG0DdPI7AfYTfYPW
kOK2xjon1N64TdEQ2O2Gb6j6+8BKaZBTBgm5fYN/CODp3qUhSy6ZQwkfzBdf8jQl
jKJvlpHxGwn4Bgdf92EfmeBLcT/g6ImhNIpdtAVsYwqo/vq483pLhbrMLCZq1Lk5
KqJv3+6uVVYS/4/X86oIRVpbSFllBwgl97NYhJBKrXQ+Igx57IJVusFFBt8a27cY
6frGPEbr/eWy2SczxagzhoAYzofG4/52qBgOfcnaWFp5QFYU38qQVw0Z4XYPrFlF
2rgO8ctrx8aBV85FhkhOiQJhJIsU+eakq8vsBhdrG06nEK7e0zD06zg6BjKXoaul
nwpf8Yojox/SPpJ73VBBoJNKi5ZxWJZdn6e7QSEd8UoUHK1OuzRiXKYCv4eegjmF
r1zbq01F2GhCXBEhYWBut3KhrRphBJcVgJPw7SoUjfXHCtZMQ712HxF2njQ4zP/6
6n1zO3ARiS6PcCZuSeoEGV6/RmsLSkudwmy3TKWX+MjyPbM0a5hgyXfvfOMu+GLV
44ooSsCyWM9j4lhvT90ZYLqlaOaMiGIKZAmVJ814ImK8PGFVqrxiLLvEVeb4ymev
JwkntrqCafhv8MLbg1kVIQd+60OF4Dj8LCYVtSBR8KKFT3SYSTOSguEEJ9Qlr2Kg
gT7vknq3PuxVyFCI61wGXD9dgj9beGQ5NW71Nil+a+YYqdGW5+kc2UwdDiMYNLIB
MU4zRlvJdjJn+FtqdZX4j6/RdQmqbmCtjN0qsDacVWj6n6BW9R0R977Tg/5Dtci2
JoUdbIJaHCIyw4gLiYGOmxzCSeO1YusTev0hrFFo6TXOWVQwjG5Qs0F6Q2y9KyP7
oAohO62nc4Ig1ySL8n8TzlF/zKz5JOyv64QIjh2tAQYnIaa/T93pdxo6Vdw+z/AV
8VMPb11zwbAtL/vAQ5YCu9Wd/d0e5C2Q4VRoCR+o03iyBM9k+j325d4PqvcHsIwF
AADkRdSSuOsWnJd9w406/xHJeSvwPKEZkNRryq4SHK/7sNc/Ow7opCx4RyJiCZm+
Ljq1rG+Y5snXU0X5h4vnC+dOsDVcHucwdpqcS2mcpvWGAWOfkzB7PQ9zIKSD+RN8
WTgbhRQMbpNrvPvE0GBietyaP18l5E9sWaIgRUh1xkXzSsupxnIpO18khLAUeCzg
K15DjPe8PvvRggeVmjiIaqOk62S9KY6/pdHX56oAMbybyfB+XZtmTzmzbxTTgnxE
soRJWw0mocFFbi5oO0dbdpVD859MqO2LZ3/DfaHfXOeYUGgisZd/GvGFOC7l0M8g
L52RQ6yipXiW1NxEbfscQzPpQnl6F5eFXnK338XwJvbVQhUUqoBvyuRhagJc/PCV
rM8/tBWkzY53jkHNPz/vjUTDKI+flNCjxH6Kd5hFBtPKlUzmIdRnlxHd7W/HtnCd
MGKxdMha44WZUUE14qrjuHuhgdJRj0URnlrvt81Vq70uASUY0Q9zigywBKBxugLq
p1ngxndB75L/jnmS01mK2sk9hWOk0DnU8cLJA4pt6zvrwYGw2RBivl+dsYYVjV98
xTv8uU6GUMhOail4p/pYkU9MwYV9eeh/4RfpUnBlFYpDA86yoDq5C0IbLYe8VlOm
OCT2UeWc/rhuo+Vl27eGKpHgGti6kch3/e9pS9gltYHb+e6kTEIlHCsAg5JcpVDY
1PSgoD0yvVkyCICOaJPavgsPZ1WKHyxGGmwrIGw4pjkrv8uUd7+PbkmhaV1DixI/
8rgymebLO3zR38M+F6TDxL37UHizeE1KhK+XLgk5jSRvX99PZ80A7bcKoYC2zBbs
yVcodU3MMWr8FbuRUXlK4uR2H3Mx5JEROO+SkgUtTXKWFJZU4GvN+HeZHyjBoFht
fTogd6mybtoMECRi61hxsjTkDlMxUfUi1m/Oz1KlD7n3I+Ux9tdqL0GmY3wfEKrn
TNEim+4r57e6wXH48FH6hAVa744RQWefPrDcxfnTaYqOUzNRREUV0etIoweGfVq3
a7CZ5MwgGO0XKgkgRBzGAaT0l3bioQxv3lUsoiOe0j/vgqXTSkhjcV5EjaKkTtsG
BhwI4qyCd6OyvhJR0tDdigR7fkQ6A/Nb7kW68uoxWsQrkm4iOxaDyW6M65PxxnMI
eviEpYeGE/6+zA8mULh+aIXSrOfn1UzwD623Ep5pYI0wl7oiyBsiN36nV7ND6hlO
mnM20FTvJsgaNpuL4vqCxOJxMH4V8cQdBuqeN5gdGPOHEnrR/wbkMxd7nm7otuA4
LdchzZVVTCyq1i1ZDzI9ZrNsgUXjlVhIjiMpp9+MJmBCbUDbQEzLFXS29VWnS2N5
7ehmEKoMaPoPerMdLGmMsUZuMWphxliOIiixO9bEXOIxLG1OIoUIvNsGztoNMmwN
N1ZN4Dc7fZYFAf4ZXrfRVsCX5j2rStUNY81rwJZJiBo/6sR6zIQbVQJzWTpKd1r0
Ue/DqvFc5m3fQLv0xWYnm7GGwWO1bgLvW40oAq6sSrsIhyPEd23+80PY/0/qrEOT
o9YK+QsXMqD7/VxBRjs9theCUAXyzrvMtrSMHLov6/rHipOq0vuREf6OLb9Q7dW5
ljoNUl6L7KJj6M5lGupQdYdLwjT9c4arxE3Velkum3BMzewcQ28k9UlMhayKuS9H
Fw5hyfdKcbDqC5luPi0q+3bsfhOdyFvnpaB00XdR4jRgw7FkcY81HyURt5MdADDj
UhMqKW1dQ7qCtnwOrAlkIc9fJXlx3AFJl3h5Zm4trh3Bujz4wKDDkDwuFgI8+qXo
e4p8Cxn8M44mwK0zkcGBHH6llmDZpabV1sKHGtnDMRb8sQ5LVKxUPTLHn+CoDiao
ZjDunf8p9XtnRVT0Y70RnKStwTxnFLnS1vahszvCwg20S789T40saiJ+mDr2ND+1
HNlVn86gNWEFQewaPQE/bmP2uqFXjpxs+dVgPx6Xl1mBuuwlptGR8MYqM9ZUTzUf
6kx0kUHJAExYw+9A/tU4VkWYYkIB7lw/V2wYvsZXurhLmDWR+i1NQWIJhtv+S6SY
eqaNTVlHP7vqJbqEk5UK1o0n1Ca013pRNYPzbbAa2hQfbsENTMwK+U9LOaciTzij
R/qfWbzTzqolaK5yJaJp8302EE7DZbnLC47aGwgJUzf+bABYUbY1XW7G/3WGEoF9
MKxRJ+rkkzqoozUHNCxKKzApxVb+/9eQb/XLDFeeYeFeSbK7eb5VVfbETruKqRET
MubSEO8ZFRNrQRJPmqZ70Ebi5AgWSlrgtaLpvmX7eyfe7siSKKmDm+mubuffJrAy
BrnkPJIwOFbEQAJPb6G2DJ7hdLoBUrNNTFSEvUgq632EUpoIMNTNtuhrA15pkeCz
Z6qWf6lB82pFd14LoaP8PpFCBZYxdcGYAi3wTn0DyUUHzD0haebDpgOsRKE+twn5
5zhodkcq7QXfyvDdYpvCL+avOxBHQ6G4dSqKEqz02eIeBuwNXVsWd8AOzGinnlHh
ydxYQjlmI8WR8q+KQIodfT0Oi/0gSjD9zRa1qO3MOpiQqIxPQpaPncArx6VUhwPw
SSYDMfLvZX2I2witCHmSBSX576feXTLM9O2wnT5g01F88rSg7QRpwdAKmWTU8rOz
bWqhWpVr4bayN6DKudLm9ds9j8mGVwCNogggixYXlCoY8z6S5kcsGZFoAdd5I0+/
1t8FUtUHJh8x1zUv9wwwjLzCdltXCGRabmGH7mGPDU5HjIIYafiLWNkql33hP8Ra
YpATg2dJgmLRJGP8jzyB4pU5GCoGYjanXyjx43xt8UaRCK1MjaJi6sHFmmjwU/HP
9ZSoOwdNRJ4l+k5vtXhZoVLY1JnzcmQKYUHcuXIbyHlIocvZ/mJxZR+yLnQicjtp
xAQFJH/i/urxaNs3eOihAydEtnUOcMKtTICdokuSVgdFu9MUGgVlD6DZ87O//8Nn
NcaBO2W3c0lpR0HzAl9bc5yErKCvj6k827LJdqKzdNYUIxaogctEaUVfh/4/HlYN
+pIoCvPSZe2/O8DYlTj4c/lR1d5qzglcrJ3z/16mL+EC2LZbhMIfxOpj9ispPESK
PHoLb+rnsee/5SOeB87sY9ct43dPZ5bNyGrxCAMti868m0qQIKtEm7r6xLntCbqp
wp9Tm/nBn9QtU0zQU/d7EemjUcPj83xnWFndHP3pzDVf/+VpJny1SckZZqIVLqFj
CcdXnon8LSDPsXP4ihBKpGzQEPJs34SDMJVT8TTF3hLF6nkEU8qJrdXpyw66O36r
QWcteWI7lFM0FJHJka3ic9nTwzEPO/vXrRYeUEWSDwrW3BkF7QOqfYjhXtqQrqyK
nWf3o8r1pwara3LL2D32XYAB1K+Vm/kZQJdjnGZxXFJJ35mh2qge7yuP6EWy9Dkn
SnsITbNUEySXMXpcCk7U7RynvD2LBjhWxj4l8+AbT1nVUy20XtvhIalZtSd4op+M
IKsQx3v8cGlGU6DvE/0tSaOT34EbnNHc5RWl7rFfZ9qzg3QJkX7xN2lcevMYg75X
XST1JficsBpwq5Q9FiNWBCOhAJ2WCMFDdqvH/OmEFrWVoIlj58cOqC5AgNZEBmuI
RE97oqd1HDZZq7hXOlefoVLjuyi4a6/q8GYqn9SCMNaB5bZbFarL+eimstnyTWtH
3bdOGGdf1eKsnCsqkLs5QxM8frMjUxH/Bd5Ky7J/vA8UfXhYBK+x60SfLuLMj8r3
qEd1Tjv7GFjmNCbxK83ga4n5aBBluzRdqkvZYAAmfZz0fheb/5qHf2sB7Ckt3M+y
yKyd/DyFOoW6F+7KuqJbatWV7dR6i5yWT1dYUMSvBvLsFLf9IthvGAVZWex55xTG
0F0Voru4WFQfYgHN7kNVhEhrhXTAvQxRivzrFlbvLhHs9FX9VtBJLyV1GF/0qly7
xZc9/lS7STiz2yxAOg1eKBkJKm82bQVY3VVlh96yQ902z32Qnf4E/2UT0ypa3O3r
K8k+vWlxE8oquZiXSNzgVNbahanfYgqad7yuYVh7jLO4uHDb1V8w0AVZbkIOxNSJ
AsW8YTKD3CnTt+e5MXtaPaD9uTcBEyzyn5m9zQGpyBYbuDgmT3rSjJIXgF+Ohf7W
Fts80hoUz2jyb3GZFze+HRC806IHVsgjHE6ZdCsK4VJ4ILqTC+bWyVa/4UKGSKtC
8oG3oZWPpEbWZgo/AyO4wNw7rX4rWhE9WT5/WOCq4CpnJpqCOz+byRR/ZX2NBFBD
T4ZV4yvof02M4YX8WX6vKv505YIAvndrGiduYUMoJpnQJNZLayIU0g7dkc1LAjgx
l3LwCGbFyi+Nkx7xtT67expM1WPWjKsHKdz1Qsoj2P9wfhYClnqZPivT8gwbrtqv
nem+ssEE04elrpcFzIynvTzrju2v5gbfmi96G385gqjLiJCGVzciTIkj9yHidQTq
cDtJQ2vdK1alirwyHIFF+TRKxd5mZt2yA/gzErDoQW32qamnPx2ztXb7dBhjy9oE
C3cWQTIKvhtGAE4HwqcqyQnGVikZgMw0URSp07vakNdlzn+xjs7V4purb5RMamTM
Oe6Kp++s/asjz5YmMeyktfPNBygCF9F4iUvAEP7spiSGBIppi/4Y2rgXXwsqerMU
S//4/ssJD0OnL9VHWOa+/ja615BFlh4Yo/jMsi+ygdV0zrLRJrdtfgDgTuxG/GjF
j6/0YiUHwjRe0JJ/QYYd4nVkWY+UG4ev/P2mnNckIIime6hgldH30+qfd9QBTKiz
beEwfAGesWLwdrd/BH0T3mOQRw6UMLmX0XYYMS5Qmi6i5JEMfMGPIK0tP7CVJGCA
Fa8MoRfsePoIMtWWdcoUx0g0W56G+hhmA06+N1mhx+Th93zrCVIngZf/gkiAM1q1
rJ0fXPat+uWmtJ02xSOGsp+FDx7K1D2NYM4m9KsZx2M4+tB5Jxtm9cr6ucDd+aKB
UFpGBXJlSjo9K+tOpfGvVx+kD+cIhrvpRy31k+Etm0SI6khynDszO4mAS51WfEj7
P7dO3lzQdsDH2Ze44PeIb+YMvyyO8CnHX71RlVNp7PINQtpY+R/ke/ky/MKTKcWU
bTWQtMZq3+VTrVrtYOhCXyEJdCQ3XF79h4ccKru/weMp9IYnh0Xocd1hPwkvDMjH
feb3hPobajM7X6MgRME2suByRB4V64l8oHWrUQhLv4TDZ31vFRiRbZ5lP6q4xJhT
8F74LAyE9EJkaJ2tYZ4FABd87PU/MiKEmAQdWpNJZlDNkRF4TpVT6Rk/5WYYR5pZ
YR+Dn9p1H2Oq/nozgd7WxmYLByIm33xvouIJ2aIFtS1volQboh9zQXuHssCFsYfp
X7EZ8ctTjygEIIA/SCnnXhCcNxmO2xjuIuazx5Qb4Q+v2v+Ur/BKkcNGm5J/JcOy
SdKKVeDSMR/0xezt2/wXcE2EJ54KIbGPZBUhg29tNBgTZQEsyWEiMLukEAsVvKSO
1E+2AIlvqsdz1k+F0nBoA48KcwATXofzs5fnoqOOKaFHUhZLOyfBIFGXbEBr/GYH
JjLF6aImccXe/D8bim4fLOCMdz0p78uZ8Pp5SA8ty/mdVg8xwjS/iX0vLZBv/Kpp
gGFwz4PN4XY6dVpjXBugqb8BjxEN3WSTszADf/fvQZ5bM1NnLhnFQw32jjkydKJL
YeiBAmcXq2uNxYf4RfWUWLIO+0LbJzvJd7I4glNnewYzJXcV1WALPw4a9albMX4q
SCoAzsY/595yvhgzGqtVd4C1Y17CVxeF+O2r5aKjYOkzR1b0WXDzhj6AxSzsjF0D
y2NNzWhVClskDr2Bx/HZDIC1P5DXx1+ep/7brSMR6JZW5Mc9N2yN8wr49MTEalHP
y5S/mKclamEeCNwx6btS4x8Mwt6VCh2tb/1QL8RLlU0aho3vzpH8uExHq1mBiYIz
g0bm3dq3eIpPz2Gg9rTb7sY8GBLSGM37XNvq+4NEEdm7SNIREXmWuG5E78mHxS1e
fczg7kXG3M7q4FrI2VFrJVwnh3P3zDb4LDmx5lhyRq1sb6IQHPGtHSL4+t9Y890y
JaiCizm2i+AmgUjLhdeNUPf9V4HdmUQkP8rzd83kxUfaJ5IA4sGjpjIj1GC6hB6i
wPxksPhwyNEvJgSSQHT4iA0vGhfTSKZ0FV3eFQgchehWce5T8X1jTDK4zK3q8Ux4
BusHO9+CrXSOp4yjBbBWzMMuG7bg7KXkdnNc7UFlUqi6pUCOgzBNBsghQXi2mIL0
0RtUbr3b4n0ktv8kQeQF55EFH1M31jR68eh+HNUZl//m3+wIOgdJqHANdVRMO0Gy
T+nNYFsvnyiP3tOiFrbK7dPyEz1h1i8H++acsV6jAreM9ICZOZyZxLWJi407Imcs
YSN4Ut6ny1AR3QKZuvqrdGy02LU+6FZR8qpc7vpvljM3dwsCyJyA1lKkRaWO3+K4
07d+tmz7CqYAUNTAPbdpbO/jmU2LI/o5xaTFcFHWuCPpWorkjJtbCM87ryNGo8bv
vnozZ9WAZQnwmLLQdxiycLn4pc29Kf6H3l1ptcnCeqp7FfZr+Pw7WT1RiVW8GMkq
UD+S04f5PgJUUjZWbVCLF9idCKxHm4kbRxdEK7CsBs+FmLiclIGveBBuexTOl/8Y
2KLYo/vtfpezprBLFhHq+ffjTpj5my6vY6wV8YHlUe4vExInIwo9BXQYiM15N4KU
dZuWjwYmSlchm0EsZ35IhCBHvEzhtAk5PV89TzlNTx88Emz8h63ZCz9lh2ShO+S7
afxdCtcWz5GD6NN4aZEO3HJfSCDehXsC9C8c4Xu3MTSmNxQm56kfEKDA555gi37B
hUUWQeMPfwO41IwIl3R2jxXCx6Gq9/4QHIzZdYIn9X7Ivf8IBFu6gUO7SwGrUcaE
Aa8Lyy9/eV4S9SByeIAtxJqtG/a1bTJeeYQ3SpXCQNmBnYLjUYT8VCRyEdun0j3N
OFmSnVDRe76x+0EHC+xM7KiPGkYAh5sXwmoXCARNY/1zV7DapOypF0l18hKBqo/y
kxTOF1UR6WZBk2TQ0vsKqd19PL76KdNJ0vuuUB3p/TUseLgucdlzgY56Dp/+nHjC
4djs6ka+9SHLICY+4oSV1ymwB2YdA2VK/N7q66JzyrRt/PpHmUZjDZfRfCWV1FMT
GfZmWJP0X+vrBEckA8uOp1/mmEyDLzMtXLtq0wXa5vebbrgD7vyC6mojQFuu3rTS
yc+y7Qefoly9JWISt7aAZo1DBMAyBLAp7H+b2fvW7VdOMG4HlzsXCf4YBHSw802t
0X9lkbfIhz4MEgqgLVr9q21+q3uFBjjEJ73CbW1G0Gadg3XkMiCXtSCWVTd1jSnw
ACZ0zf4MEyCPssb41oiWzzmJBEUQ7zDnJReFIpi3u8+9itT+MW1d/L5CjG2U/+cO
runoKvWqJCkjyQdIzTSyF9UcYVGfMAhYUScnHo7dnN7x1VKZkt3jV8SbMB6XOv18
hkpvMzRwVVMTy0cAubn64Yt8FwpFtR6rqRhrsG/Lmxqm9BKqms11SRZz5lwvoFMi
Wrmw37+CobFGm56Gj2Vktsbs7aJar0ILqef7e6oCni7Qlu3X6bhsdkSLOu4nHhXu
b0Hr7Wqr3cihva4bFHV/EWKiGQF0uC0qbu8hZaPI7qf+SpntGhWLR22lX4eWDQGy
YaXoiXV+mufbQa7sxGkdu8H75sb/uAkBvbpTOsLxsow+7EeuP+Zv654pWO2Qsy9W
rGwBOQ+XjlPajjKkrXCLxdrfNWKcCZRjcdtGrUL9rvklGrAXhGxFig2F6dJmChTb
PHhWKT/wglsymdSGf8Jf1KJNgIQjCZpc73RRXX/Z2arscUpSmEUi/V3GptFrj+HS
YhEmbOyYRj0+mDNCCfOpI3fe7L+qpSDow1UAVNDtJ+bLZBg+/mIhCIbLmxGt9ub9
8dgLbhhV5AOag1/y71lcgtpfv6W1ltn9hv0fYqVwuWcVdEpmoocSJ7RmJcsGnLya
1KY/QzGvyW6VlR+YwfjNEMB9z3HGxAwvODjmmAkNhnY8r3s8xJgJsfniD/5KRoTS
+3od1J3pB9QfraEsjKGfnNon06w6RD2uw30oTiCuj90P2MkojNH6bSM6NZIvJUDL
`protect END_PROTECTED
