`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8dW9WhhPasl8LLrhzhuKD2/ur2blnAZ8s4jkjKvw/+WHwnjzHG5/o9db/wy1KW1u
T0hmAzqzJLW9DvgxaeNK5k4H5GZuKkAvnBCsXN/jlrQ0b1rHwJ9ptjIG4+crDpLz
4B69oPneGy1SNImnEoKm34tRoLrR3zsAwxfpXnGOM2nGUdNQgd4+vp0vYGMsOcuE
m4W5qK/MW1eXpT0p5u1v0+yP+Nnqro7spM+ysSyy9+uPFN6frYDrtevc/GPqF2kL
0xjvyUhzIgIaW7siwjhcJde6cZLRyl4gu8yKFY/AjIQYvRhAVwrrRHvyazd32J/D
OihAkqL8ZYK1hcsyMZkWS15rFPcmVJd0QchGJpIsahV3vad0nUSP6rA9/KbSq+ba
DtfSNXjt+riDiAcPUfK1Mg+GJuTXnbIXVux8kRmRT8RObu7p9RYhGdoVz5EXCNYt
qCUIJg4ow/F+9ZK/qam33w==
`protect END_PROTECTED
