`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eed97hHY4I0pBQC4mh+ag18Fl+hoUXU51TTifPDs4DoMXl9PNASpOrU3spPHWWVp
cJGEbsdFZCe9kDN14aH3PlqVCtUxigK5SK9L+H3SDdK7Rg/Azi13TTc/EQ3NUYoB
IXcLo3W2gx8tb2G4MRtwx7LLdlOAG22gmnvUuYf7tFcAfWAv8Gft2TaXqmE2M0KZ
on/1ZTFNwr8gogFKt4/C8xn8y7ocpuUHH90olYn5TgLq4B57E5szd/QmK4cdwuHJ
9UB7mpR3DcsSwfsU52ktbhEUSgMikED/YWSCGU6GmS1UpsrN/YkpfUciijwRS7vC
WzmJHMki0KeA1MF9xuhG+MjHLlSijOVMT7gHQwPKxwvk1C53uoqS3GpiUk3H3bT+
8U3otghTfSsoyBrn+T/JR9DkjLPk8Sg3UItkuMuF74CYGLrmp14U9QGQexuuKqIb
GvsSLYkTzua2xq6BWIdPdYW/jwYUcfIkf+eG5fc1ezdLlqAUqtJ0TxQPLbTIeFwW
Uy2LJB6UnqJWCMZnh1zy4IhKyYUU6QJT66YS2T5ifd3u0xLRytqKCJo79XT/F6Ip
M1Im1XubxFjP+qtGR9tivUjVR8+JzAkMnajmHYKwcEA/G6RUgbcyA6JFLVKY/VW8
qs+sBgvgHXoLGAJdha+lkektc4itUF8Uo7a760qUHHA165AyLR2XHaRkRoYCVdnZ
S/NHx9sx45H+h6PFDpD9e542rzVV66zIrUW8PdQyyHA=
`protect END_PROTECTED
