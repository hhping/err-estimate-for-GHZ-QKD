`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YFlKPd1NF0TAfHtHMLIq1jWV/30uheSl2K6zrVOdmBd3NiRrNjYWg/X714uF+/8l
FXj09AB5PSzdB9mq3sxX+3W2RG4XRjLyjUzl8/JGcq85OM00o6rCcWFcXA7xPwKu
rfzgb66Jlbo5Px8xsm+lh0/8tH5EKrOwp02RrRNMbn3jrTgns2BgTfkM5b2vI2Ym
Mk+VMqn3xj5uZdwmKeK9eJLXoPoHkVgoErEY8OX0VxOk5/OKSwiJb1gwj6py7Ig6
uw2FNPw7fXzkonYdswKdn09NyQgo0VvGniKKBJxzARAvaN9mRVufVou1ckm9vZUi
a1xG0TwM+HOq6DaWk6UCzIQYtjF3iOVWCHCwOMCKKOmcbPSY7B0wY4N40gDe6R9F
iZ3WfqJWj2wh8gE94A6X+ANihHzhhfDnMLr/iTNr4wDoH6q0CgUjd7DG/YPT52Vs
UwTm/kyh+ws3EEfRhwYzT3Ro76uLsRYBgiOxCR1eKPSgO2R1vEclhNcK/x9mZM87
y+jkVzwZqBVv696rH3aY1xpZKZzFXThe0N05tKw7ikh713NmEW+c51MblnjcPiHG
dahJstrJ9pk2mTnhZPM2YPCgYj7PRQLUbiby6D0W7u90Ebu9rGHFCsS0HCHVx05P
yAdzC+DeBNGU5jKfscKp+IZu/C7y90phTsXz59q4qUy99xrAsM4SrYxnCGj9aidY
UmHzj61ApkcnxX8DCyocy4Cf3BwnVJGzuVXXrPLMmWtq88fm7JVrp+oyanraWc9B
DZWIqhiIuk9jr1keM34ml98MsZUNPH1v3+tTWoFdxaaBvw3xM1ZREnuwTaSxsciQ
rhmMK+Y+PA7HfLq45T2+juxfNortU95AAqciYM3lYkayv0Snc5aBPSHg7hlRbpg0
`protect END_PROTECTED
