`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HverjTo7WJdZN0CEEVC8TI69pyRlGmxIzgqQIKznkjDJ/0PWFPHi73y9szWstUvR
NnYT7RVe7whqffg1JEm8XL4yEw3Mx05MRSCGdyObAuWCp99NKU5+FpRpQvOAfWJp
2JhkowWUk6hvzFfv7H/pfWnaFo54jozlqYzR1D50JCUx/zjIiAwcf6tmQgVraMt0
OJkR5bAABY2DovouXc12lcIqI4eVKuuMpuZBXvrZbLp7C2ga9tzDxGE1FyZVLvnv
vn9HGg04xStijempEcqYdEN1lAI83MR5h5iZbD2VrsczB7gBJCLc/KN0U8jsNW9X
9vWvTnGOReUsTFUm7x5nCOlA2OfXM36Qb7JO6ehkcyY=
`protect END_PROTECTED
