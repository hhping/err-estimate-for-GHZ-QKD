`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GtOoyY7SANC1hB4cvMDgQzuyNH+tF5cdLYs+RvSBPexv/VLJcElJFMGRa0+vo84w
SZljZG8v0qNbgsMyjBHYUuY8/whFzAzRn3YGefXB0nmD/j94PMBAOv2LzFo+6heD
U6F7M5IlhtB6WiXThpFLqHLWSz9t4k4WdRZ2w0+LkZifFmgbVir7l9LFXM/iD8PM
tghwrccsxhDDPijpyOoE/5OvJvvR1vin9nOrKnHInv9Qso/lDBBMGJ8gCh4UdnRQ
kWex2N0IuW0zowKdXYZ6iVYrwg1vBjHUBBiCl3zqTy12jOO8ekoKP96JT8pYYi5A
zfq3T5xItKLjCw2xBqepZf6UMtzDtxMPnyBxCi7bUAReWhoLIaaYdfOLoElqlv+z
fRfDNkblmaHb6FkvmXRyeW945fgWVJdy4WR6xbm2Zp6fMyLHJMyZDrqKyHCY+Z4I
HRPOR/sWrrIr56nuZ5Ni5xKFL4CCDpK4baXov0DcqFsx+9IvS8uhXu3r8YIXU8EL
`protect END_PROTECTED
