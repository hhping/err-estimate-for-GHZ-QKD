`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V3WvPBobaEo+FKUHc7fzn9wZIUvhaIPgVZVebKdg+s5T8tKAExFMoF1KvtlBc5kp
PikEGlbcEuZTxre0HNK7BToT2GSPWURhxk/KjTSdIQ5lastoiiV2WZBiGPtLqkIm
y2d1WFKdbRMauXAB1UEHBsHNIpnM4JrZ7ccivAlcDnX84UNiaMsz9mPO9xdRv3/f
AbX5Wy0fjCLRHgcS1Nq+ICWh1hpaBVAADVMUsrAGn19dEH/aKiG4JCm7g9CNNkoR
QUmKIeETrM6rEBs9m2vlzRerFFqMXAPBl4y5fCFSjjicvY5vzEx9L8MWAHMVuNui
buau9suPIA85TzTDLPJfELQF0rjvgsfJhZ7Efso45j8MNXMfIrrgMhkg5JGQndlC
bBYblSstHx5O9YWvBidEFZuAvhEugTYAECjhdnaNh9CDsg+JrZLS8qUw9YzV7f+K
d9znkIjosCO7FqyKzJguWv9+ZYMr5wan7ROZedryjpL+lO0P+ZZi92gnZoe/JqDr
7v+VehZbs6C+uwKetZXl21DLEzOWept1Ji6N/xsiBQWhjTvISJ6hf0Z3ggkCk5+K
EMckbsmeT5Ak3qi8O9639ZJEpvgrdSO0hp5kieF0l8qilhnhnDTxCN1ckStkcrhp
vZ5rLQpLPuyYBf4DNYE9zn3ObWAuEaXJvy/Qshy8La4=
`protect END_PROTECTED
