`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YpVIWjwq74wH3FRYFIBN+thqB2xY8ojGaOx1hq7JHEdG2VnkcBBc/hEHkt3vgzqp
JhdbjIMmsmv1E6ZJXRW0VF9ymvmN4737jBFKmTciRkPPF0hL3zDQ6rP5J747bqRh
J4t8ZzazAh5hj4F9FH/qGu9e32uqGVlTYI1Mdpk9OnhEPYUy2rQ9BF6Y8SKjLu9D
xOwbdT3hYAJ7khDLdnQ0r5+sVw21YU4Ceigk0xNZMm1upU3SFdgfckRbYkUK/UU/
ZCNMf1sNWLnV5EQ6Lk1pIwlvWctaPlk0hE++79n3v53ENJqdrkx4cWRNXIcqR0tt
ja0e+uMDeHXhVNc/GGU1ji5pJCR2IBco9eEI7uQvgCmIw/+MCNbQo+z2iS3fx+nF
Ud8ZWViMzOTqRkil2BJJ/dgluYI1+KM41h6E7oQTciVebvyanfbPnf1M4io9CsNr
lAgDUbXOeISVXg11ieQHsETaUkqBkqTGejm/OWwNeji0bPo0Vy+QSEvFVjXdfjwg
BJcdK+yPcvQJKK8NXD8e1KASUsfeChXTjVknuEGc4/i7v930ib4ExTrmyCpUFcKR
+RwDrXEI9PzMSdKhz7VkUWQltNxfnHsaKFtGi4QLCv290UYVdSVEMSXoqaj6RHXK
B5Rr8XOaZgabrwol9KPdebAogbnK6DXS9zdIMPqCTmAdS7cDPhYXmiMpgAyDmgjf
aF/f3RPcRQP1HxzSydnpc3fS+FD2IIfl15xJ8b9AifNSFHTqoSuI1XHNpdWmpYm6
rZVqKk5yBEZeZOn7Au0PstHCR/O97f+2N8pekZd1Opo66WjfcATTlCMl/FjLtIUJ
NkJ6BouXqIlRIbYGbcCLIIANOkEuY00ldhM/c8JbJiDKfJ1bYIqTQdcexgloD2F4
D9lXPryUWmzYXev7wYQkArcft1llD5UIM64oaAgdoYDlHh5ko87Ux1YureROcr+v
FQu8c55KTHxb5crSsB9jRDhAuGgt2d9pMRwLRLiievMPaVlC8L9RppWy66PUzaVs
W02MsNhzSfZk5WiCVBiXTSMhlqzhwfsjXh5V1E4xB/OAUO1JqN40e1dSS9o8JLKO
/SfaLbzBN1/35Oq0TQAWNOSH+s1ncTZW/znzU00QyHtE056plaJ76fNdHtdzUnGd
tx/phIRRWOiqBM7CSUgaWQXdsar3Yj+pq41+xoGPBVnbhl842OP5Q3sxux16NHru
uTE+Ehgorj0NVYiy4kR2s6jPKu/zY+mWj4ocr7r97bb++TikopC/2znAVoBYqon+
Exu+hA7n9+BDsuktxBeW1/k6VH21CVhN5/yn3P87ALJEC/S0XNUfq3QnsnAJio6j
ZLAfs4AixfA1qzT3MpLJJjydxQvf4ykZEIoVNRoA/9ENZJ0+74ZwRf0pA3CFz0S7
FEitibTW/Ojt56VOj4zpTTmb0CI40/Cl8EhGCp6n/FF5q8KcHM49Ob39yWY44uKR
Sg+Pp+AHQPtAz96rUVMNYGqPe5fe7/uRsa8F85/tQ6PutXVULC+GzRIg1wcLy/qj
9yXZahrpmP3UgHdmDOkPx3X6ZZ/iVEN21Y7mW/mRkFZGw6odjbVsjkajm1RYYfXL
zQalSKBCaK8RPkREwd50gAEU9eedBC7MT5xTVVDYxQO3mJgvN//LKKgxXiw/pdW9
g+tRBqKxTTuZR0pW9QuDah9atUP+X7lnGyYPphcckACutXNlffpxEbWA3MVCdqmm
WldFaR7QcHr44XKb7UY3eUf2s9rZItrJc8WDfVUth/c4kqX3w4axlzrENxNRSuNY
Va+HyqYHWnKky0RaPXjF1uRlucFJzLdiIjzFOreUA/et8rhxVShETvcRBvz8vHsG
VTdsXr3Nv+jn35Mg1Bahzq75+UrGo/2jPcB5QtNlnplIR2k4YG3igRR5/Nnw8YFN
mJTKmUmwxdKJ/gJB8szLb75seTbm9d+ggI2zXnXRJMQE4Rt8Pxqp7bei543RjSjj
sFi5rdVTfm+r1Blz2/F2L+mm2/T1xRes78Q4Hs/JOPOO3bVCAz/VHxo9Xkz4P17L
XjaGvM4KJZ0DR+0W7pfrJ3ZUFUcucb4wzQocnrEL20f5uTEdKaF2jGRZ8v0jVgrs
QG0jZ+y9/LMmxJUObL6iq7Z7XZrJqOztjoryWmsKNYitmoblj52M5T5f3b36f5pW
NT9//8JyBV6XaJEBlg2+PhDJnmm3Y49igMUdFdkbT7FMak6sCcfHDGznsny3meGj
sCtJEF6dHjBAYApV1u25xybLzvnXL/r5QLsxqIA35SaX3LQ0AUvGtPRGffwNOPJ2
iIeHqQ5sU3q1gn3EiU6ba/unjK7zpIVWZcozrU9iSaA8vsNHOsMbFlDrUUueOhYj
qymjnvQ52gXhJD+c7pgmQpEOBZYHMrS0zg7eMWrb3sPnDuQbiNZ5HtY14Z5AaEYQ
TxJ75AEIxvTXs8NFYcRJcWkvsC/Wsjm5ccLlJaJ5GB0DJoNuZdeJb0z59E5802ZF
djZDgid/a/Ju7TFnoHjTDx9XgDO8eZhnWSfy9O+/KZoZ1AwFKpBhoTbnrqB2/Mbj
Y4ahcsvLnSp58pbxIc8Ek3Hnr/cx/Pp37bQHPATSMIOpnNKEVlceD8XgBt1yJGVA
PvGFbIB/A22FCF14N45Gy3LUx7DTsq/UeMUcgTLb0+2/JQBK+rOasbJHrQ1cVgBd
VdACYO5ia4/7pXiukxj4JyY4tVYSgW9dP/5GXfogszclcwVYG589iivbVLDzoT/3
lJ93+CZ7Dqnwtyf+qZ95kIAazRGfvIh43B3GAzpsbj9gq4vY/6plpc97RVkGmoBX
1ikJa0UNVfLjLc10wbayVXXhfMnkAfrbU3fi3C2iO1gHD+04u4loh7+X1CeQR+Mr
irD542H0dWbDZ3h5A/phis4OhGXbSlvGUv6Ny/T70wKcxvl9YolocKElMcm74K+G
OKlpfxb5kY3vcD00tcF9N1OJNitYNZVR+GPiiGOKs1xkc/C9w6xZM80RwUlGtZiL
PcSS5YQtkCNaRiEAotKp7+YEZfc2FqS/YZfG1gzv96lEbVjp5mgZt+xQ4QIQBD4k
ZtgLSj4m0/hodS+rjwpam82Bzt5SujhUJRJg9tm+HXIMBx6BpmGuTr37VOnlqtvu
b4TFBSX9QRKMl5i7aEP2VWnLp+1/do+52kOo1exNd8a7wqJboPaL5T26LHWJcFQG
1esKrOl0G3YrHP98+zjUCVVQ+ExZPngvR8ubbR4YI2qG/OQaFvRU/+ba+wXZ4f9s
qvitg3Dmc3xm8Xv85zUsqvaiMA9djTM917VUZQv6gbqsyV8x4JinWXKNKp8L+1uM
71X8fpjXS+hqKoaj8Ctw2rnt/BhVL0cyzzIeQSIpV1ju7Jy46g1QR658+oTV9YeN
qGW5LNRVnco43vgpwHagsRt7KUKxI6s6bybkIlpnWcI=
`protect END_PROTECTED
