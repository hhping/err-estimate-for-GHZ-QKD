`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B88PpOQxL0wlMc48SvD5/jd25jGJ8H4EtEURns79f92xlJk+3a8+3QY3gri2yzHq
dfJ1/a3bw4RlBysQOdIE0S2ptrFptwxDWEPMKDjiU0ej+82/e5LU6np2XfwCFvqS
53QCcz6XDy+qo509p10V/KU2pRzO825PMJhjUeq4dYDqB+zJLsS1cG+y8c9wtIgl
4hOFI7cfBws7XHpSVEGK899ocvs6qmvcJ2jfwbLrNPV+r8RMMRHYueayrKmGQbf1
ziPwjEj+zGf/fThyEF2tYYw6H/P3pu13sP49oaCnxyHraXo5QiE5WibnLZ/kO1gz
59ZECkZx9nF2fsUnduUHLbSMKPKtF0Ix7iH6XwX3nFtIqIaR2DuCfYu9WyjicKXP
NHu0o8OD0bZnauJ9S+e0q35s5vtCkPfNHD1m7J15HI3QWfRu2jqp79oPjy6XDt5m
GZINBUi8Am2oAPSaw9AWshypyKsUM+M0m5aU/F3ac5vLHOdmPGBaSH2E3nOzUSyC
DIG+F7xaekhCwXIMLP4nOEvb8YXFMFh3KBaWqbDj92Is8ud6IV7TquXe3cGQ9cL/
vAxmoXs4imKMyF4KNgncdfafehCAN562qGbLMqOs0Xh0UnHHIcAb/68nfwPuPA7x
GR9AwA2CJ/b14+RPMgZ49IfWWXPD4Cym00HVTJgyZCKEhf7TCH6ieJYYDJw+LhMw
GT40XV0sSdod58HpdWCXf3XWHbevEddgkYrnVR1DvgMMR26BEfr5XISYoY2kUhdy
IXJSNMObzoKzgdW7Zi2GsA==
`protect END_PROTECTED
