`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iWceRPNa+lBlv7PSMngS7onbwnsq9zw+aEdJK4bz8hr0tiFyYWuGwo2q9oBojK1w
GgA/gn7s935sxlyv+jyg2dWQTJQ25a5uwX8lbaCp88sxuXGP6eIrzBxuVo1raY90
W79FbYkVY06BcYe2XcB7MlpvYvPkX1wB/h9poLG+8y0QtH1w3q6ohJTEqK1DgWvH
LEVeMYle4dDBI0cqI1eYgM4VmjDKqED8vLM8gpEQqUJHQM/lhxNhWLg0D+iukB5l
swTde37Aq2EaCeNP98aANOtDkPsCEFXQZs77SwEWRRU1ZQ1ra6daXTXi5k+Egeg9
q0ekU68bQm2rslNkRoo7je/EOKCOz1ZDCPk8nFcSwnGcIwfJ91c6oENj3ljx/akn
rVuGOrdw3cGBq7Pc5uaOG2e9CNRDMqmnoTVbkR9iF7LmdZoa4X+Yr1l0J7AiGmEV
bf0BHa7cQZffuCYSwTqnVWCqrIT1oRXCrrS/91/x12cuawRxhTOfTo8RROC/C1KZ
9Zld74Lt8znGOLA1pviSmhTYokMCEOON44I8zzYCHhLkw6sULGjF9uagCI9U8f3H
O3OtvS/6EUZaTL6o7MrUd7FdQfUjhrnpsYUccKbg3POLqCukNAYVoeSQz0EjUAVD
yc1V5W65vnSF70SLxmfGjDCiFjcThUcSdLV0L5WnuFxGzQyTcC1oz5IzoxGiH04y
2CotUNmkFp0rq+RTuLawPpynMBPOXogTY8jGeS1tyZQDRLCIm9ND8GiscsA/SNV8
4RMEdw+kAJuhJsEIj2sPskj6ngMb25mH8W4TfOpkfDTA8EGnm3coVrwhXS8TO5wI
9FQnAhTt/g3G1lK8m2W2aVv1GzGtn8DmUbsZzzuka65BGU+PL3FPfl8+Tfamw+/x
SsHRilDaBRxeFEcg2RgJmHsJuivd40GVR0e3at4nayjlJcHM7YxdercplT9dbVvi
Lmb34Z1LEUzKisDQv6tP3vlHvF3p/Po4vZQMuGh0ShkUeEz0t727vkvFcOMrhXCU
ob0rHJ538qNEujAX5w9RxLTIhcJZCQqLs42mQP4pKwcMe8oRSRrXN4TxhkQ3LXaR
Gi7fNhUuF0QOki3EMUe/aOhgUxcb1dFhs4LWnDlhIXX0AaeqnkcYc0pGOA/5mq1b
sItC0JmujeVYiCs5LeCSTcpLYwn9mGeKtsp8KagKrFFrs/J3ADJrQq1JXiRWY0nK
HhrVvWrnlJpaaxKYCCo+FwCpdt8aYTujO7i1vAUFt0NJZ52FJnoEdEeDv3sUE4Qn
bnrcbUh65ZDlz9NvidrWcIHsjOOB6LMSIjEBzkO0LsZRN5y++Px+B8Yq0ETFutP6
Vyc7hYPJQjw7Vpmr4WLpbtWSJyOXpa4967t9ip66dd/lDOIO1KKmbtSRlMdBT5Gn
RFiWIaAqMJ5GQvYNDqwrE00lM8VdKLHwlnyfzdwmj/K4MefWJnrITcsP6PH+zhKD
FigqOeZMxROLy2zIzletNq5TruSKmLHdagq1lctWOg/F7D+OyLo0JRfT95SIvlgp
840q6odkDpuPFLIOd0BJ7fNgJXWnoSQdmolC7KoZ/3uiRQervdPy6mcXH8T2XhZ9
fOUunQfK5RtXxkAOopaNZ1Yp2mwP7at/SP0S9r9aA9gmSjcYYrQLMxla6LMv/3q/
tLaFvGz26BRpy7nRYVEmQSmxV3gARK8z9sMkR5k6AnVRIk7kLCNPGFaxa7vp5wz1
B+3MdkLVs83FEJdyKPVXpci4ibSmVRCdvEfV+BUqXJjR+d1CD0WR1J39fCP8cCzz
`protect END_PROTECTED
