`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DYglonWPRfr27Q3dH0xeBjGN9ymHr33uic3WhwmLJusFedSWISQtipydGX3YZGQz
7Tqse8f0YLViKO182siW9zG/5p5OlQPE2sj8lejptQFhDO6m+PqjBBHmCO3dYL5o
t+htjP0555dBAsLAIV30TXA7IH6jx3//y+yqDxY2JgoCqmCVNCgcwfzxYPMTQxuj
oXU+c3TsRrFuF7PT8pdigpn0I23cQ/Bltlw/sUGYf55XxgPQzb867ohgE4PsFCxk
bVTh30rZjdA6jM+6DAIQs/FEjmXyeXEjJdymOj6zRojRoqSOx8yinki+HZMYye0Y
0juWzxiZzwQSjJQvWh7ksCaobRe62VKbVIcgsxRZ8GQT1HOcFAbYy7Vrj9wMrWnF
EbRrzLMRNRHWoQvzc+53HOF8tQF1cLwrvyVjaOadaFmJlNj8EIJoWp525iljhEOs
CDa+PG22I/1H64mdsEtuzr0ZB5+SzjZz+EdLFKJCy6LMgLDU/udJ4zc7Ciy7NpJ1
y5lvY57nJhM5xQxTFVzk5PqvqPDp4auX6uZO0S55N46udDB8TDzse4fC6kDCRyK3
OUux5rGsbjbQKkKkpqsxNPT0/OdZXeN8RSVWHEdcwbpXSZTcg98rV5xYif7VhmSc
4Hu2qTr634wRldwQJP/4rSIl8zqSEKoTexdFXL220k43F5naF9WKmWfLG0Eq26aT
Z20OhJoJtl3SXAUkC+rl5SGQjCBp8Ucyj2gPGkvHrgcSjsGpG2kx8yFrNTeXO8T9
xI4+EHuGxkjm9u7iHdBYzI1uf8p3fiTzYSnDjz1vJTJH7AqP48UrKsPnS6/KvuXi
ubzh79EnK2kdHAVcboZeknHHmnhtM0L88NokcEp6zPcnnRVFzONpRZKlyQK3kEAh
sYKdmxvoy30FjKXH4LjGx3D3xCWiKToo4wWMQEGjdSYcjlbHb0FcjkIQTEuk5fsF
005/nR8lkgTVcVve6ZmWIbHnbP+nWAhFty1sx1948/UxTvTFwCwAknPo8F+RRiwC
4XauyeOxN5HMf96BSN1vs3Ppgh8mQzUXPFtM5NJO+Nxn4akTMhErOMV3LwB52/WY
3ol0X+RLEUYeR+865mTa2brITm1v2aoiZS9K/ZM0gtgsJuU0OQNcpSRyL4t3HI2v
A0YcIh7WGjJafPlwwxBO659a1LDXtFWC8OrTfWYgNEE=
`protect END_PROTECTED
