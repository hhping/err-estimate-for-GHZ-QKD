`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/L1c8kIIF60Bk8/d0OwPgJ8yNctGOERILWPLeg1haetqhAeO5LMlqXwIibxyk2lu
gsp0VL3WVGmq0jDZKQFXHPAuoSH9MyhJAN1AzWvLDWNjp4fb+6pLK2kVk3zG1yJY
jViZiMiuqrctP3lAPKP4FWnpbsHjHBnrJVfGEuQQveYZ1CTPNqz7WJfKc4ca02fH
VrA+Bvh1PTLv52MToKH7lilodzKghgGzZuGHmguhbhU7gs3FRzteKKHZmxRbQReB
qK5uKSALwZLhukhQ4/taQfCGB4zPhOlaaIo8eCmrSLTuTcPXLXgbbaRG9LqP/S3y
99WGI+UqPHfqpYxwur/LaLXhgfwy0079wvji0fgbIAHk26dwdK4SyFPFBpgdzhdU
Vjv09KKRFFTiTEl782iPfcl2x4Qkxnbzx1MNKaEnRzzwFdEWEfMqCC2llMneVUwI
fLzdHti3e+6oY9Kxv3apHm9BuOQ6O0y/w1jCKjF/XlbfiCnQnFNu+VHmfk3HN3jv
`protect END_PROTECTED
