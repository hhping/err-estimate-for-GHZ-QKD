`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yl7Im5RJjS1VMRSjCpL8evKOSzKX32/PRI7EYO54x0iFJviZ7PEjb0khLkMfKQ1/
yCBabm8V0GhEFAOA3+hL6bREXxUUUjXjvHgnL4IepzgrRjcR2b5l6OuTZlopoeDO
4RNDwY18sMHUx8BbD8IjYYhmE0aCFPtsVziDXpVzOlJexNFGSnC6dB4Y5O9mK+av
6MGcXIQ6ggen6O6hpXo/kM4Lda+jT8OFYodwroz2vylpXoWzqsEBLNoSUAB+zIZz
uSK9dLWokoiRZdSQyWG/NUYdp6UbmyBnXBMos/n3eVGFkEi/YUZdS5EImhcQASOx
mKw50HImyc6HoTNRw1qMZFbgGbHG0a1BBx/iU1uaHCE6PDgB0Z+QFLK4jYqqCeQ7
2tMCtDY41pF07P8hPJlsUHINs3H1agKmHbLzjvA0gfL9edWE5Q/ElhestXoZ15dD
v2KmNeGTu9b5yRQPDYEOWLnjA6UJ8oEmpgM3hUiSuTCa1AA6DYuQ0FB1GTYYaTQO
AKgvxAGLfo5XeOlINTTtwKlJdBZ71n+/7PROqn23Fofg1hm6Fr3Bqjnc9c25/IZ5
w6/pEp6V4OvuOtSbB/RdNVn1WiQNtNO7LdYugdQnLjX1flCo6tN742BWd13TTh3G
BPP+qzbQnwk1A3LP3Xskr8qd8d7cdPbCfuYRHlgoSRi0GgpOG58ks0gIsEnC/Yau
0JfNqSA2r8gOmI0vkEhW2TMsJQ5++tjJWsffkUYZkOJ63GlrTYG5Qw/TeyR9wSKF
1YnwQUj66lZZGDMnDpAYUq3etZMVs24M0djDmXBoCkB34gEM7oTquJpHXzg8JJIv
yczXdnQlyhs/QWs4DdyzHEW6uF5m8a8ElEt/9iev1hnjw5A/GoFuVPmSf82LCXOe
imufoNMGLnqGdzT5fCyMDw==
`protect END_PROTECTED
