`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HLY0v5VRspiH5rqAeBgZm99PVyvL5OGztTnCgj5eB5h+M3XIDWehX/9gTm9iKJ3b
/Qxd3VzTWgB8diCP5OCyEPfZCBdGIv6c3cAbzJg/3pcgps3pLi7cO7WoBvmmOQrm
JwCpZs95ufk8W31GpORg0chFH46kzVUcrT6M5yTKmh7Jh2rtYPcaUlM7JKweutse
vMDUb5ovJRf5XQMs2DzWySpZilDmvJsP7VSix46B/R4Qt0N1WbiLHRwTCd9ZYtr2
PPstmdPwO8I1uLsTi3+oheDqoATb0yMI3tiDz09Mq/tMmKBs2mxSt5BxHaYAD6v9
c+u4a+UC+Q2THOUi9E4L14soXAqnNT4FwuxnFF0FJP324tqbfTWRWW/FZt7b9sn3
SIGv6ZuabxeTUOpwwqlcFa8MW0+uWXRteBmEFJRIb/f+wNhi56tkvnimVb8JAcGM
UaR5FVyLv7eIH2Y/QmVZaeV5DHDbaEAb4BXcr8OIulkhv52C+WZrRauRnXzEMGlZ
EnTJpRmr6p8h18fZIfDXY6QdBJFZldcIyqSJO6/4bIYAbhX+0D78b4PGIJfhdMYc
FIVMl9wyhpD1E+3zAZcf8aDVVZO2HaWaNryrUz8bNhOq8QRnvXw+zuYdBlcBB9Kc
qjo6E9ecqjYdhnNZOjVctZJN53tDJ9fJAJ+DWTKdOEQ=
`protect END_PROTECTED
