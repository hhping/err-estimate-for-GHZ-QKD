`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6u7eVc/HiRadlgShQtCBWbjG14AfuObFwAfv1iWGcCCl2hmj7ko2Zx/xLlrSXwmg
K5kZbXXopIAj0ctVcKR6tMxHLqr5pVNIFYC6sRQkifUGwQHd28B1qrya1qXFUv/o
2ty8tG9/NhEjn+dWButGWG2UddgDWB8sAczOcYDEffsUiGue33PlKxWzvZ/+SRMj
/yR6hIC1IkgzRML+5xz21CjexIfkTjPNwXTJHK9w6U4u8utmvxZ8TdzHbbnkrpVq
478oHyeRyyhS/2ol5ivcD24uP16Ef6WtGSuYbF0etpY4KVgRCJXmx71/yl9CqxS0
uzEEO5F+5B0wI8EeS4oykmLc43LankhtU8huyUcdkUGVX5MxcxZMvMK0OS0iJ6LN
PbIVEu2u14dc0plIA+VdXDFyuHFRHNfKuoKNeb2D/uxhQXPToYpUug+iKvO/J0+N
YExm1xYYgVc5O9Jx0mNi/bK3U7sjWE0z3r7IaVM4+c+ksqofB9YFUdD1RrwEcmlQ
c/nynK3JQ9BFMHmfc5xMTX6Vk5c7jgqzyy7mo91m5w/02R4qZjyd7X/ombv7atmZ
n/UinJX0kUZvJaE6Y0GQ9+2VpXGMZnmRVnAnwOuYG9U/LB7BpY2hTumD8Mh+RXbZ
T30VOPlAMIFxbp71jkUDdcAnm5Bs4cB2VzcTqREfaGeDP8LnSvba+UAtthwPTJ7D
vcQw23oEzRzCUOkaFIYkaLpK6HwQeeBAgmbvGm9AJS+7Is0viDBdHBqs9YckOETl
VIgIXvTLIGjAk4Wlxo0hcw==
`protect END_PROTECTED
