`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WJxYFpQIMiBTSJnHLCWK1h8ZFkTcc+avMJUG1UnppbB+E0f6HLk+T1u1E8UE52Bi
F/MNKACCuO2/B1NEpXlRtih56H2jBGDl7S0ydgB53xk0q4pcz066ylvseE1S8UNB
0o7ZUXj64flbtpQaA37IERIfvAT/xLC7Z5JviJnSzhX+rau9m10xzKmV+H7iopuo
90YDPXbEGZ14hjqA04hqNSKChGb/GOrTm9vcKDZT9B0bv3jtJNQDZHe4hSj5ZxRM
RXTydPpFhbsXZzT8/NMFNzMY7xHbQX63Qm9TTTNjIWs6ADlOYNpGVKeKPg+DAav4
OESvX4OJsKUP0W+UGKLQtbM40b7oc8YftUNu0u5G8YhMg8CiQYCxGoMx8p0kTHBq
99KFMy+QXV23v/do7iJ6rDo+7pDEKTed/P7ctkcL3JVoktd3ELXQLI8ftQQ9tAMX
Cqe7MFoV/8vXX6wcWInY6AB1wmmzX/e1sfftWB03/BKXho7U3TKT4xgkC+Wuyznu
FJqIdYZbmTFl2btyjrkN4RzOnEW86jvJalCZxTNBBGzsk4a8jQLjXL0xxP0HKUAH
o0RERjrREMR7hJJ4kGcqpIirtLfkeU7LG8oKYkg8wvUZGmYQgjWMBnAo2VRh+Zer
mSbDhRuvjNujNLbJHXWR7l13Ltl9bZhyEw5ST2FKIjkRWwN/sZyhY363xgBvOUht
u+wcgBtJWt8FM0JJ4gO8jR1/izaHeu/g6E8L0OqP/JWu9wrbBhZq/9JrOTObur0l
jd0NAjdhNDx0vxyGcLRJue1zYIfWni7m8vsOKkUhntEm68BXsb2PsuIBDWDh9/AZ
Z/eGGr729BIQyGZL/bfGYWuuxw1KACVUaO4i5rqtaExdAWxIeJ/gTGAOI161rTj9
2ClI4bcVXf4u7A5Ac75U/gDp+xweouOQoISFlQ9I3lupgjhid96huD5t1YcxgVgP
8SaB7ARBYBEP8s1I9g2+tWd8FVlrO39lT8lb62FzCfZ1Fs+peCNN2eE7izG1ADY7
SrFzq0HgFnudqrVZQKJOXzN8Iyce5e8tWE6Y8EZ/73b2SN+hk+7voxSWj6b5FNOU
WaRlz+brZr0CNUL5tORGbvOgSqiVDyuONDh2niS46475Bj8Pk7QDlSz/qtSgKujf
Ye8tPozTwk4yX/WsjBqf1ObHhY9xvXRPSTKu/9q5u5rEms1YSaKDEaLExiGcB7tK
H6s3jzd50JXGm0KAf9L32003/euU5A1YC46+qTflTQuRXxEIvNm6jRN3412Le2Cy
1VaU7HneUIA9FQYjMYFHZdX3/4eMEasIZ/7u7UqkCoJrCpUqLyfxGmwgCgswMDhc
T1hxs21S56jdiqBYf8+GUN2LzAtzcTQsXgCHG4cWPT+KQAr5vD7xXoB6p8kfOgwc
o0AIVoVpN8Iuao9x9ZjR9f4ibdSlUIDLoM3twGuOP1kQ/FLZKFkJq+2bgN8axdOB
QBZmdMMQ+j2TgUfpA61Ynb5hQZ6X9HXCtm2UQ/8kT8EdMM3dlkDdI5ZWCujNQ3LV
R9UILhjmbXY/l5lUBYhVItEDMDThVP7ukeA629sZeVw=
`protect END_PROTECTED
