`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7sc0CyNhXXkIi7AD0B8EfDcAe5hvcWUk01frROdjd3w+KGBCsQ8P2BpnvNSo1+V/
7je+j5NqmVhLLTQJWpwRtDt5md4YCPjTGVB8D4bcXBs4f5RgLcd686WTDktwmuXB
10wR9KvtdTUcGNEXEvWyI5DZl5NuGBoCxzjCMsq/G7+y8m8tMI7r4n2owMfURvHC
IDKy98gg4ilWfDcN9Rx/9ISlMmyWV9YqUp9StjV0jP/K9sgo/De7yO9d4sUdWC6b
p/v88mHUNu4JJ5WCi9m+D0svCUxJWWlnElejc8yhJ9Wl6ipKlMUZrIDJmiAo8uBc
k216ozOq5jdA2rY7Fr6GrRs4lZDiO3cXiFOljVxLBuKRYxA+dHr8P7hgGMOrb1kf
WGXlT1L+SafVWBTCWGUiyp1c6Pv+gO3sL86PmIUaqoPE/67vjG6rbsWtNdqhCszD
sZ3JGSBm1gxV0CAZ8mcq8hocO6Er5p7dJ/GJ25Q5tdWfQ/D3mfMo8H9tOD5vkotx
BAIP9iNtf6mJ4oIG/TtS+6uVCjfACSkRxPMUfhLCGgsvH7HxJ9v/zMUUQnGuHSok
8kQ3WYlYr1whBKIV2KB8x0Gya6G1k9Ed3HaEbl0dJwCFS/RP3/xcV87NCjkYCASt
yVq3xiGmSNiJUEmG0QNNtXHdnYSubxRstRM1PrjYjKoIUd8+Oxf8yQUItT4Owkim
4WmAQnBahc58UudMH6jFzARMRaiy7tjco1YIAVCknh5oC6Tw7aIL8GzPkQ+wHxVo
767lKKsDvk62bRyz3PGmG56GCUcgZkYqlHqWUBRzKy8vRxY8SkA4hyNChxqKon/L
gT/OVIj/hlunvOdrEhhnCyLRG3g7VvOJNhBGNmc9ypUYikADM6mAuRUrHl58lHjE
h4w/kgwr/nyj8oSeV02exVVci7C01JI+lz11W8LZtQC5OQ9qfop6dpPXQGn1/ZVE
ChNdFh+SO8K2rzWVmYEFWNzQF/Y2spnuMINXlKI1PLRNo537/qTNSxAMG21wthuN
tEi3VxMbQHTi+guYIzyH4o1knuqdc3FeKnOCGNb5lBvBIrg4ARVVGGs1dqY7NLCF
nZduVE7DamkZO3OgA3W+lPWZVZJg36ucP1ga8N09wyVfkTQFhYUoRl0ICMpEUUzw
8iKtaiYGKlHyrNmcBis80IWRpKiJ5T1JZYuBkY/h0D/EtshJ8hZuWAn8cDsrw7cW
+LTOUbnV5sM7zs3YCvxq2SNMg2MRs8BbME4VJPuSRv6klWHqj1/QxIxlCEj2xR6u
Rk1IUpGuwX3sVKDmFkh620+QtnSdnZf8eoxMrMS8YsXKyD/qTiR4Ceq6eUfbDcSi
wcibWSUmlASxNMMEXpnPbK0wPMy4mKyM2oTll0TaCSVnLWtrX9VmubEXtol4ig8b
/aPlaVUzc3ZRhoCBP/poUHUqAcpN5mzH34wT0U8I2os8zyWp5zrXxISh5QoVIf7G
M+d1zE47pKMTGTQ7pTsE9sJie51rjM+2oyMwOVQLh6GIiZ0QFkOFr6ED1ULrinvw
c44rPC89vTQquPhmy7wXdfxYlvPfgjsq386Yjuz78D4oo1yXgH9rqcApTy8eFkHU
88RXWEoL+zVp5eJHchnvGNBZIVPDy8bsV0XwBKEROc8mdWHpqs4hKBCdXN6tPMpL
J0zEQopMAJSQzSy/2lSnDjstOSfeEJaBJQpxAvyVP6Ih3YgIhO7Ez7+9/+JeeG9b
Qj6zo93ebRibR0E4w9EWeA0veh+liCQ5aCGygUpDNhynF7G4Iu7D+zkG0suCK0RZ
M7oCgHAbHt8QN0Nx5vSQmaFAl33yFLu16MylJ3ZP9dRYsMfnOSgcsWmueh1Ks5nj
OrChX3zBKvQexCMxYWJgHToP9E3fCThvGPnfbRsNZMZCSuyyfAXbgb6pbAiB/OQQ
Pnh5bpcCEjmq8iegr1XE1nBtHBC1rMnmRDF0ytV3qPV156IdZ9381HIdHFTuZdY5
c9aIEylBvP0y3PtY6SRiCzTSdsPW49ieeta1bIJfyiFOBI0lxPBoeB8NSIpnCQGq
Udg59+BF8+6CYJQK5AClZkt7C1+Cesu/vGRt0EiNojhK48/TV9P4mmOxTvnklKIv
5WL9ffwaYT5htwZjunNpp9dIchD7/mnLvLKkLmVNJvuwD+S3oAfsUaU6jic3Sm2W
PbGJMUONwRhqAADC63UocoIwgRJX191pR0H70aEMKgb69pYm7Cc0xG1+vj16QYaG
64msxWEdFmT/72AXUKuj0ILcpptfRziAUg6w/jhej6mfOpNyyaD4im5hD4D8Ki4r
muZ8rXjK7YGMyTvZRR3IBCxsRcOWjq60ThUpnyb72nUr8WQz8BuFNl4IY9+nfEtx
q0GSXdBqwzKzPFQAJPja3BINDT2DCovjSGbMI2E8lxvp3OnsYW7owo28VGjouM40
JGp3y9+CGDBJQd7gv1rMft0pdqUYnD9IhvoQgPhglpf5cptYO36llRtcJDMuXMk7
BSku7J3PsCXovNPWUuiQBASvmCtc0RyC0xljr0McRhmdPRPbdxUkHThIXVKoVyGa
n48G1PZRpOBPhEI6BjApeQ0V30tPGI3iPdmlXZ8br8Sw9PjoJaUxG++dFYEsPCL2
sLoIwfmHeCiHynsCzroDus/IO9ins54il1S8f2icxb/PjuNO/c8Wp6KGN+EOHsVW
3TDCN4hjtNVAQmF4pPF6VoZk+jx+QMLavofsBoCDgxpuMrLMrAlgoDGD4xRROMuy
X/V5O+aEUeIRrMO/XuP9Z4h23y3OS+fC0lC7EB17HDDjogPRnM+8kAnpepWFFjdS
ta5uLtLi+EqViJeYv+l5gNTka5SojTPg3VV0Q0UBXIo0J7ViYDnIBuB3GKLq/eR2
EJ1j2XIfJVkd5Pw+gXT/l4dtDPip9idL+pFhJk0fjAdNEeOiVKg3Nas5qKPSMTbS
6uUgSkuqAOHgSAy06iuODHaR3ik/nSukSDFODz1OtUQaP6MEpRITx5qYh5Yt/h+n
HTjtHbUnH4reNf1ZMGURsCTI3UAgdN9V78paiDfVJOy6PeOrv/DUdRRBLEWgdB1l
lvqI/qKzatV/zE9NG4v1VuQQ6OkHaYCjyaGcBrfRkjRgXNd/LzbHqUINqa9FWpwg
glupmriO3HvsnV7IUwFEnX7ccgFpuSMDP0AvVkfopXHqcpp1dr33aFwAlxU0rpA3
x7kTIjnAkqdHMpEBEN/YDRyMVaOxy2Xag3Mh3gG6ggeoWH6zaWlds9rRle3bqjs6
BD2107gWXO76KzQxvXL1y+IrDyP9B/LMCh244fREDiIIDA4dw3XpilWa8r374cTU
OQxbbytEG8mQmRdofwtCasl061uyGIAjJMO3GPvsIBQdoqFnURq9o9muhgxK8Fnt
7ZIF90RddnMw1LxPWZOnS0Gs6Nou38+WnqWmrg/RJNjnbPnwtwdf5jdPvhFmpd5B
XMEbxbgaCCgpCTlUh8qVyn79ja6gMepkjULPGSSfbqK/RBLAdnTdFITNYpcWxMp7
GvP1TB4z9pP1JIPGuemLF56nXX3pizS0rBNATbUv6VHtCbXBWQEt/LScrPTmn0tg
jruaiU7CBFtXl5wTCSfDUyeaWfEFm3dEvgq7/t2MJ3C881KqosVOhCS8K9+Vb5LM
7oyoy+g3AhCW3frFd1EgFcGEd3g4dKv2rXqNmXL0Q/nihx5I02UTRx4XQtpZvEQh
gA0AbnbhGumEsYK03JTPExiopWFbQRWqUNkiIMOFSQUJ32wFQJLGX0q7Zj3yCwmx
gm8EAa/kY4ceF9+y0jZoGgxdK7neEAEQMr9ddOA6XyrwtCrsxmavXMq40B/CLeat
4di8eYQfRdDkGZwFHH8nQ+Ghg4PKr6gvinW3lGwXgfuh8h8p95siDA6uOnLJ+wZp
j4tuRsC+fXAdRnYvExBYEp9VzwZL2AJIr4YLuoxBiBu52N1aQ8ua7MGShN/+q4JC
pZ+Prx4el6xnoI+72jZsSSCDQEQyB34bapCiNCs2k2PqwQ0IylYpIxMDP3TyVARx
f5IrcikQ+uULl1zgEwgkhOs9hxsR+G09yqs+r4tb7UZXSyWoLOL+MFcUQX8i+1CH
6w3XJ8xBp903xefRvYEjBRj7192sPt1ERIVAemPfTNrKqHD5d3DAXwUeCMTO/weN
A8gaPgrGQFddBEJmN0J1AFE+3qZLrtDMoT+zfO4V9eu3OTBHj5IjkRT4W76NDp6J
H/MupvpqVOPWBTMPEsD8SJnVxd2MjGodqtxVAYprIbWgo+JIS/2RPoPeCWw35f3s
jg6Z8/vln/MfUB1Pr1MtAcTwy9pJIGB2878LhdvSynSzLqJqC9V3uz66ByErLfrb
3OUsXlxGEq7PcYxe52oZd2HT4EteIJBEgZkZV48RMld/ylG3/oxz8XHdo8ICyxxX
3uRq0Jm6e9jBYtJHlnhv8ImWeXJOAXqIDXguoAdpXT1nLrMS2GN6SwHNoCeDk6OH
G75bMZT6ctPP4C6200nkJm3phNi2zFGIhXaqM3b0bknAcAQktEQEheGuwjveKjTF
dFTqw29fp3pKEGjY1Il7RqanKqg4YZtWrtuzh2MMCKPIQILlq+ZuCZypbd6GhcWB
4cZYUu+mqUiNGq/zR+I1uALDWyA/HuURV3A6CDcAzy2cFM8MGykeWXvkB1MyIh3r
TBetSLrLBS0sP1ClYqnD0iJjwTyIS30tZc+roIcTsFoEBbx5HgqsowHpJnE+NWJs
mnOJaSPYEbyzagkyEY1Ji3LizVe2DhkXxeRUhxMWfba9S27MMBY93sZwbsYeABeQ
6k/GGv4ZHs/tGYDywXbzNKG07wKyFPH8OZxBOI8/QVXswQUw11fsPmESuSnobx8n
ZA80UD2SeqQzDF+65W6y4FzRWwgntROQ9cKo8q3+a5om5+KF35NrLlxZWgiQNy13
FIzSUdavAKrpetmudqcfTlhIWQTXRSZGwrhfVUVmGguJhu4yEQM2X7/fqwT2XAbA
4V3YZh8ampOeur30CMCe+RDrvWwLD4BNkKCEOLDl1vhxMaVg1CORvpPCeQc+ZyjP
xt39SZApNN2vjGWunciwejNoTHNEvlMe62PUGGf3KJHqdPOtC13pkWKZ0pFrUAma
XVAo9MTBhHimY7X+nbTRCLaI/9g9T308KUOL53sAMQMvW3j9V2GuI8KgPqDER7yM
yP8tjB9Yqf8PcHVHfvFDe0zdy3dK6oA8OFPY71VdASQRWNKAyY/hE6KhxRNuvNe5
qem19WGKPoMz4PnpxSej6tub96X4m72DMEpvzf0p7rO7TPbFX2imsmEQkXp3LA6a
KVDM9NQbSoNUUW3dbRQEiKE/Ip40WM8fXwEbJQyDG36Ew7T3+dRd2fE636Zo+2Gp
gUwRToKrXKxLxwMVn/l9xYwxiS3+0JerZ13d5xA33pXs0zNexJvnlKCGJ9G2yCMq
IkM6Pbko2iuOv716iP0vGS6RObPwawys/LbFhew0LKY9iC765oMxwkndDUMtfMxE
WUb+bqhVxqA+vtvV+3bqCypy7lVs3UNTDTqVGC8Y5OFR4Zfqv98x++Ade/5zTXJ2
2paGYd9bVqUQ93LCiK+zRYD7CVfOB1T44hUhVixeNCe9ToOKFKFHQIT4xRo/DqPd
kcFb4Bo983w34W4e/QXmde9bVVoHQbziDI7TQe8pPyZWYxoQIzFstjTm3fE5qG/P
SCxMZWyBL4TH5ayziIvG6IB99MkrKzB6i5Y2lSe2OLvbkGCq5VrnUYBjOrpWYfot
WMCNXrNOdsciqgY7Vncm2A6/D+8ZPsrnq+3qEipcYeBn3sgrFctUa8/Ar/Mnq0IK
5LPdWwewWe0DSTTvhYRAuGoHGW3XoQ2RWpFQKS10MWciUqHA6W0408hVmPWWzQZW
KQ7Z03md/+GnkChQiaYmUBlB8PUenoVScmSfrFGA50cbaqnFl+qzCHRBdwELCipv
HcAO6Y1OQkcRAI++qRJaz51/GchqsxrZ4xZkU8K3GwlBNVsXcC9QE+bbodafaTXo
2ryqgZwpe2r3XqJJMqFj1mxmbtnccef/cRl64Riunwp/psSs+0+lTuwM9QxJa+BB
705FeD+A5NM1KikRCbCoGw==
`protect END_PROTECTED
