`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gaqs/cp2qNiuUxQj5RLfBie3eWWAZY9B9nWSvWUVopVk9sX9a3mAXLLiiECCuIz5
H9B1Xjo34HbrUWGzoxCqLr/EL/6htcsDitCGM7yCG63CeYcO+zMCObo1sGfh6llz
ayjMOxDrslyZQUTLJ/noVMZRQGja/b6OZXUwPVEjy5/yQTh6y1rhQynS1tdCcFBP
wA4TfE5OCEMDxv8z27O35fZnn+eXLEKRh/SkpP6sW2nmbPeoLsCStL46y8nEbkc1
mln9AJxPPi3hKlnLr6DAY3bD17qQv1WtjWA7JgNdw1mE6Z0DgoNz8TlvjRIeMQa+
/rLhnEp2Nm1tZlyScjx6IAQscyvQQWqsmY0Mec3jzlj+C65jQ6Jz10lZF93S6HOf
U6m06QxCOiiqTxnzNEJTs1WS0+43xS2TZaX0TdplTPomY/pNUez57iVuQRHEe7oz
lCoihvBMEjmTe6439LvZkB6Dje4VuuL0i4S+ARS5Iw4eGx7EKUr1cIPnjTcKd+CC
EH1Dx/ipruY0ne07j/XfPpc6yMXe38I4j+fkLggoNi2K7hxAIjM9no/KhyCUhJDz
1lmt51TQKlj3PWbmF2IEW5rKLJIh4EaCbM9ir2Mi0VvbB+grHDOgHykd2MQktc0N
X0Ma8LlLuv86FJvuxz0WD7ZZtqQNbPRQpGjFGkdz0nWgy7BXPVvCZgRG0CTJAJct
/SMt2zLBK6sXF0t4XPpQMFv8SWdM3yCmZabk8TmJ8CicyMu/GQfVFNxrKjq1zeUJ
gusX6Bn0pLJMODv7yOWjPoVAV0Kbr6TJtQOfhDp1XlOglma3zO30DiOH0WjGmaNZ
gddMNNS1XfQ81kf5KPk+RgIbvSPxqAwcCs7TBz4gkoQ2WDPYQl0CZ5AQx8wwM75F
TkdGvWZRSqz136bSD4nvrNk91OHwj/BIcJ9Sbg1/IMdAcB+ynNC13ea7x8gctucV
WESm9hHvrQeXejoqAywg/ixn1Kx1+nkRA3jXI6jbWsx0GkTLWZc55iUEC8tO1cdT
YGV5LCwc2QspVID30h6m8DDE/hU7n173eBkYg378VmJlfVW7mqpMDhbzhZbOGffA
3cZmGGVPmEdrUYYPr3uQmXsbEFlXSGGzK3m7bdXinUIHfYbasitwUM5lXVXoDl0B
pyvNc5oGRgrnqiQULvS3sQkJLQ3k07W5V1cmbYhe9c8U9WGUQvUsn9u+TQafDMHW
rZbcAP4Z1xJlk+2fL/zMR6F09BTD1tX9+oBE1IZQ6hDf0N2KK1FGmybEXCrl7qZ1
X9+9LCBdxYvUdQzyNBepBFC8jydIImsubO5mtXWVs9pgEFayRhdiCCYkk/R2WFXR
7LTqjfWhg1Sqoud22xJbLl55EqoCwAmfs2eg2LdHbqh7eGeFB0LS6EsX4/7UtoC5
rOdgVHIRkheZrI7OI19F3xZevCDvRl5ofSJBdcsHbPA4AxkPzJqKanzLX7iuRLV+
XCUvmDLahtXXHPNkBOHfOlNCXzcTjsYP9TVIgyCeo81SoQJl4+1tdE7WOXn/jAOj
TxhIwzUep31Qg9QQJsAJi4p1EjnqRAR79ZPdl/arz+jNG39Obw42xlKIpUuxPA+B
PcdCqVcvAi5jo0Xfu3GGxyPXOpdeWgKtaWns0wHsXSzGarrh+JQy0YwA7TnoH3j3
PeXWNRyUXXGL4Prr7WzsTE91AesAEbo+ftKT6J/BPrIIq8h1tO7Vxla+m5wfLmcz
u45d8iHmJm0WqGPH4QeFBBghIK12EJDZvI2OEPcnD2QLO6+SF2CUIBDvO2ozYV7h
bdC/gBn35v28R0z7Ixgv1aBxdjwGsG19UK9mO+9d6BJt8XPQEZ9ci/+5W4D+PZSL
dIydD18BuSzUPGE0RnsLCjAnhK05mAnL7b5gCrqx5ISz0ZMvxEQkzCSKQpuin2Xh
2Q5dYpWbJZCV2XzExYRGKa7GgG8fiBTPJj21sdoNXgX3bzulZVInDMZbeJRxWCtk
XOdlpV4NRcHTcoaY/7+fBgfJfX81+mx6RqeCjESgqtxFwFwEB0TiV0zQxS+b9avU
7hkGLfs5eaKpQPoixiNYyW9IClABy81AuqBHg1b75brOpL0kim+ZEtT4gsrRG5dB
s8WsiayCsAlX8zAhj7PJ0E2eE/QHXbzD4ywNqkTC7RVGg2iFcYpKu4SXWQ25PA7U
0d2BlUaA4vSXENCMzt/eevGn2LvfCLQ/g+HOW2iLmdNk7PmTyEbxSopcmOmqSnSq
FalSK/KUHFRHwxLAMTVL1r5C4SSaj68KdJhnO/2ztxq+1KhALX/j39tlXdnTzI6h
D5P+Wz3RGogckNS/dp9Dpvl/jdSb6GgeMLx1Vmf+jemAmc1um9YgnsIeq3biJhXZ
5qQ+pH5OrRTH0nY5zrgZ7Qm6LHHQIE68AumMMGgDKrA4MygNvrYEpKFK65f6vG7s
nQS0rfBdt9j1G1bZIbBjz7JBJY1meIiqdFltqvSSrdb0Mf1FeFIKfEQplG0WJOfh
ABm8y+6gERCDuX1Uk3KhPW6UOosP+fI8UJW+xarqlmkIifUxiML+Pxt1IztjTZQ2
hDpbVzZ/+dVvRa9E5fOBrbOBuGT8wL770hylRF9EZ2BNU6w8J2++1paM93NW4wnn
u67YtbnL4jAvGgTqIwFXmSgKonqo/OtMrA65pVOPh2Z8smReu3hpNUSfq44USo2N
a4FSHcRmHdkp90K6ZY/qMBO+8G8oiVkwr5B2Sekbmng5IBawkPmqrtHcBSYjuPcI
KipuO3ZOqV1sxc31eS28cEKPyhV2pOTP9YHuVVj0QpoJup5u67+vx6izYI6qFOQH
DHxlAs3/h3YCuNfiDZX7j/WlzFWRJsYu57ZU0dy4O2IVaUJNSU7bTxPTcDvWDqyR
WU/XMkchZJHMUaGBMltk6s1OsoWFUAh8ZprY9cTeXUljXIJ4uK1gAoQOMEZNcFAn
XQJUVZA1/PieIHJZc2/iw+3+8b9yT1rHVJaMa1PB1pO/C/Jt5MqdWZAOblPIu3NA
e9zN0XeDAtN9KWkC3IRkTaEX3DNQd9ezj7gy0zH6CAyni3IbRMydQ55s4LspsE6Q
9ESCV29NgHJTkdAHZaijvkakfv1TodsoSpK84IRoj8B/gVtKxcrOTui824Y/L5tL
JKsedSp/sk1fQoST7FmSFP2uRCXazhbBx95oIoD958SEiOvxIxSAjX+vv1EZqR5y
vi5YEWdeZQ51IgOKiFTGuIOWHLjcFrqeyrv4iiGzEqqHXFm6mxxPoaG43bFfrsC2
wf2ZDddnWa470HZQkFKcClWcT0bzjK9qzsT/Ee4zwyvFJupnaDAu0GxPzV7uPvMX
t3LWGBIljJXzvLBcFYJ+PRUawryEXzMbSDE0/rHHR/ncJZU6h55yW8ibT42PU2QN
GaXgAEMaNi1QMvJfMNYi4It48UHPQLXJJKJGXUJhPgCEQSelGRbr8JFzPJ0qXsfV
dbphyQwD1ueWoVzhm5Lv4E/3YIgtUTvr3FM8rVSKH6nC+6bD3ZTVYHg49YrnwcjD
1AvYZxhpmfa8lCD544GS790eBLcGrL0J4aa2YQmYQcTO/Cbdu+rDrLkmk7YjUM48
02j6G8PG8U5+nvqKaNFfcUOGUlw3Ipjqnh9cfEjAZOY0dWMg9iaEOrorrDRs5VJS
Rplf71W5vPdwcbU0z0Y1LPU6ktftMxTj5FAA/wsMG8LFZRVOpE+d/s2SN4dFXs+/
GFRogO8F3rGKFe8rFnmbsaBxkT9UqIEI2ncnSRez7kpDkzcbMs1XsOmP9Jru+06x
AzKx4k20rlye+DxUSquQrOANhqRtDywHnkIDavmovA0ZyglEJWi7eE9S/LLYvul0
W1PzCpzk5wWRiubKb5rlUtWWc1FsKuwGrZkZ6a/U/cb6cSpjF0CU2zasZQW+XYMJ
MZhNN653t/DCEUIBHofYxg==
`protect END_PROTECTED
