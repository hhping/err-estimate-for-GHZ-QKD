`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8mrdNLfBW10n6+UAZvp5gKF6xjyZ0AvoNO+6qKTrzvxpfGXvZ23MRG6kybIr4ZPr
wxhlNPWOqZS5buXTGurPGoM47/s/XD03QrDZRMsokTN6RBb4TtOiDhDrr80Ui9Pq
1Rr/qu6T0LdI8DC6AKQrcGJiKD0bEikRo+Oh6Z4AcISp1rAHs4ag82Y9+n12OIJp
n7uq1bCgeifTBozR4NDfBWgyJv6+eCsGFkV6nEEgG5YjEuGMZKy7rx42dswZkFRb
/fAzmKMltJnigtWis+ZnCWJMPRao9DQYU7pswsgdzRFnVpKah3krwtvfkhZ2uELB
APQN3Fio6XQNav5Iiq/WNPeMIkqBOD9AmjMRtTY2k5fwpNNyzBZtlokvo9wCVPYA
hrqwg7r/vIqhGBpsLi3KRx6+Yl38L/4iX4FuFg5Svc8lMHXd9raXsdiXA9vNN1xl
vg2RntQ14qoZ7qNwAe5DuwOdYS9AfiftA3cbaiCZXEs42SuYapd/xBfPy+vvIGYH
R9JCF5S+d6XxZeK0DDhiiTz9DNIBfdXJRLTInALLK+JHGWjLkuroA/xofMei5Mtt
ypW+nEVTjoNZTu9avxmR1ftWmxpfkVVci6YaGhnH/Xc/1/qA/h8jTQtdW7dtz7Cq
mGiC7CZ3uCv66IrzhucU1ArN0fhDuyQO5ft5UYsTZZxBNFMqIOMVEF/pOMPDYvc8
7i1/aUJ2tcnUqOo6O4PmWv/jD06czqT82YmJp2BLIYvMhFgJcDE+QVjzl1N03xOj
Sf4VqU4H5UHbX5xdhj8gdgEVoGXyDAkW9Tg1zdmtalYNUE4jicLTJc4/5k6iA0n5
JVu+Hz5LfZ2Sg3EqoY2dfkWlfNTSTNc8g/u8FQNMoo4C4RnM4h13JtLBCtmiHid9
EkvEcqrDM9GGxDjIc6kSq+Sv4s5W4B8yoA6bim15SSMAoyoWNKFWradttsR8huCz
lR7urxLlke6RFyA+n1XZlZDiF4vCzrZ3EplLAHSdfNnEBpRZuREFyS5fQv5jA3Pb
xt0wCN/RYAzk7f5l97PiwdqOD3k00YTChoufkMeebpyVD+zKKdyKeBEotMZd/cfA
q5ZZACglZwRLoOcnjrMCx1tuv/DMGuB+He2lWaJSlcVoh3NHBwZ8PI0Nqj0zo9I+
FDs5KcYGi3pDVlLnJFCr+ptpeZFPH5A7GcpqzaPax8TRYEWbOXcdXD1mWP+5M3TC
EBfLf19mxwa10GMPa04aXx0FPXdkVlOeQ57X7woDAlnekzZ9OWSVyZX8XY1Rj7r7
sxPbREOkEgPGtD61XFs/yBQA1c47aeuHs0d8mDh7h2J/AEG2FdWUAZsmshAh9a6B
JOL3oGW7Pk9hF7uPZSFTgV4QpaJrPcRExi32aUsAeLVvcIMfYPM9G/ZbC9FO0HK6
V/owMuduQA0pZn9LOG2MY6bJheXWevyyyrsPxfISSUPnCxLcK5Ymypbk4/Yx6egQ
Ov8+/ft75T69CHDj9GwBiw==
`protect END_PROTECTED
