`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b7GX3Coq0/SbLQw/5Zarm6ecPdjPRuqsAiTL3qDuAzpg1EUxNyifDzisohDB4G1O
+opK5R5tylJloTiQLlq7mM3i2cpd8aG1ma5BJMCaiJ5K2V4Tft3uCJthqcHN0wJD
C49nZ0gYWz4ftKKrkoHa1eXhQAaPbLf60o3CjjqAx26f25Sx7JnfkmVZise3vz9P
4aoARTPhiOa3R/mVG+wyHCKlsFmp3hoDEpBpPdJH3+Pvy/dLkjVGLRd8V7NceKx9
c/oq2TVQcaKoOleGtF9/i4UEVrzG7FfyiBpxjKTj1BcvMrI+UWX+/LctTicoMtxg
ZJvrsp2H8FCTWs9cbNK/xwLuvaSmmBqiYY3xeLwJoOLdjDIDidaYK56/xM1cksfi
4DD3p9unXorUW/Z4fArm7lH3+1udIi2nWqspFXstyPPngfklcxgrz5fI065wAiwD
pSZyAgNvuk7mel72ZqK+u2PpjbbSaCA0E86ztOQDB0cVB9ZMLd60zcks55xWSxnR
dz653obPQNE4XPYP+rzsF9EXfPjYdNi/56CpKmCu9RoiVVbSNY6daRnmdXRD4W4e
K/FTHSVmbXr6KPjktjvOjyOQSzMlYOH2G3mrCEtUO8doLwp0ZlGx5fBoUsLQu495
iXn6oWM+L6qflTq6UpQMUpewJ+uvAorjON9vp6ie3YqIv24K3HRJ2OwGriPCF0kf
yy6cuwdo62OQ+zlkvDoae8QybL7nfkypo/K3W8++plN3zu1goByizUb8synzNI+B
/mqCg/rAYj84QpvWQq+VgERFy0BPG4lS17wcbYPj7kSuWBKqT7zCcwGJNDGEILpc
To0GvuAR6V8/bY8NO8/CB1Bl/3mwmHJCR5QfOp4AzM6sKZfaqPfJHhvZOLvfqGVH
jDSuFUxUqWPQhGF8pq2SO5dp8ksyuzSL/83WFHDQBE62It80/wDgyUYG4avsHVFq
kSkRVsp6k+mGtnd0S5r0X8aBkssY+MBX0gjeHFAWtQMZql+PG5OQHosLP4reX4Dd
JQrpsaSU6oT4fdXaP62u6WpWeqGwvyk+EEwxJ04kzJDhYUFMIbdOjWSwnQBdyZEt
QFnMG5zKuVRNtgnLnxcSJdKqHTdz4IKI9VrUT+HoMfExaS8g9o6RnH3/bmUXbnu0
62aPlC5OO9Wc8S6P+p6Vpl5S4fzm3qazSrRtRBa6rZjgDD9SVo/CEMbXrTCjemji
qlKZicpDrqAr1MCVF1Zm97TrlGBRnVq4SFYFuneBW0rRo/Boy/N0GbRXH3Exfq7x
DH0FBZwa/1TC4qznPKpn6gzbMNbu/x03YO4+S4dJ+2i7s0abeTtmA6gqFazKvcxW
eMT4PO/6vj9eo4vSiY85j27OHEiTxaq9DkUKmcYnh8vo+23+Xcs3DSEOtaD/tkGA
YeKBZ5QuCesULD+piplwOPJJN8cv2CwHRp7a5HukTceOEQpUWmi+Sgp4B1j24n+X
5nNAKJw4/PYfEtfGuBioNEDZDv2rK7JZJUgCNdKSQXfk+CXcJRT5QSrGMDF4AhON
edRCgXfTShjBfRtbcMwZnirh9LzoGE59tyyoLFteJe/aCGZxpZ1iC5hghKjDfUMk
eRVe3OVJ/9bHYUW696xJoeF6doyshhwzCyIhZRiiY08joSARh5/aNWYbtcfvFTmW
TfN20ZfZk7gqPd7IF+pJTPigOqNXUBHWB1/fyf8xRfm4qSqoQ/1hIl8TczkF1u6X
LAlaIOfE6D1gnR3m8UPexDkkKcDopy9guUIbVTlzgGCWDcQHP3De8QNJbWoVYol6
mzxAnCZ+IUWmrirmmb9dA7fsJhXgXdFzEGhqn7OEmw3AWrYL6LgzQ4YR4np4hJxx
kgPTBzCZYjOKW9yhpHdFuS6ZbEVy3ROH8OzFOULIAEtIKthkpM20CfxvWZSGCGvE
+pAMzCIrF/u91X/yH7qKG5g/DH0osdTrBZ1eqdIn3VxINWaBtsutrGcbX37Abym6
xQ2WPOBBDTj9xxrtQe+d7XcyZgyTLAZM3Psz9aHJqC4nXEZ9DAYstYxO/G/YfeN2
UzHaZ7DM6SAXV7w25V/QtQzLPGvvhfQQ9vZvdBSM7rBrBeWR8mO4/GLA4SATnB/8
gnjOdW2aRIgrV+9YvByR46i7hZPNrhIi57jOMjYaMbSf6TPr83D21j3ovng86pke
N7n9R6wzyPO2cD31ua79HvBoR/NMPw8Qh49SCMa0BLqoiGEx770LqyYVoK/0EA7k
9js9NK+awxal2ibtrFl/GN8LAm3eWPSXusAs2PR4etXpxIGHST7Pd1Cmvd4S16Rr
Sdz1nUaI1tT2M5DFcyw5UiXu/1j4PmAmA+NtvBHggnMtIh5Z+eSoWA1pwhqYfi7U
X6GGtI6NROUSFLyiRj233S7hzEq+mpZZOj5sjQ34uTsS+YbcyeHCWSq/mHGl//ip
xFD49+of2Fe6/V5nfZWocNamOc4esqxZm6w9uywkOx16ExsM990pFG9mYu0TzrjI
WIe+dfpVlAs+Ttl+8dq/WsqBfoCmtvxq2lOa4JTU8IcMUtoBkt/V4jRyH92eCoCF
mpPhmOHuuML5Iy3ylimVMYDBAia5/qUBRdZVt0JHRB935iThgWo3NPKpaYASoDYp
BkBF/junofyzy+9piNKW3k3sq9st/k9HnXGfN+vOX8lILNvLlvct8bgMSj4S1CNA
Sv+hlg7MQU1p2itllbrEOVi7fn+0eJRSCKee0VByDiNpGiMDIq9ABK7lu0soV6Kp
mSf4hQL2EoPiDzs/72zaX/cGG2qqzupIs+SseoZP4RYsBjG4+emqYiWcmWeJOvOk
PdNXvknjNquy4pvVo9B4QmH6WTxbnLird457mtY03PNOyeIjvJ5VAGstPgJosoIC
oE3ipNw++jrqA0+74/4gF5CBdhQ8KUgG/LyBMkLIBF54A0hDAHLmIyRqcCKtNa7B
kqecZv3s/wFVqy39hD4yZjmEcwrHISGezMic8iR6U00qbMzck88pLzxiZaFUSBJs
HaZzQN5pF0Z6+FjVAh7ZUm1XFfVrQuEPGfBTfZ545EvVdslRTga9pgV0hLCkdjCn
FHOaTn/L/xjmgtsU5U59LqadrOK0CghtFFm1WIbadBGzEASW41NDvdOQyYgdQ5IS
QHgD48U31K+RO7XxC2Jo2BmreKAfmxRnvETx9UomKqMW+WNVWZkNi8o38ex8BtPU
X2NQzl3LfjrkG8Blar5Gee1QMpvvApSFZ4BX7TAft3SKcq7j7d/LOIfJZmXOu6ta
UBOPMcMt4NsriYTeEGpdMcsfYH9KmAoZFRjtFUW8y8CJDUEjRLA8qamO6HnSUZFR
i3vRROQdMRHXjPxahuOJZMIa6uwjLPDXnqmOBRiFx9oqLITre9eS4S9livxTxphb
Xl2U/hPppkAyth6MpfcJrR/4J0EFjvYzVxGLHwgJS2DtuROqcuvsJbk7Ofb2aA4E
t7FgEpbG9j5J8QntcLsRrkXprcRrjtHm7xGg1i3kuEdVARt0HijhJuQgL3s8qGjR
wDY3p+LxCin1zAcYPEe/r49azL7NbZW4zviANsme3LTcBpDyKVvNFBVXaH1Qo55E
vZ2SABaeBoKlwwlOGSU4STarLJOcxeGUZ8KO9y+TJnqxbvrD2MAc20nFLV4Qz+oJ
l3SwQDDYLSg4oZYMmvDp1Eytf1h+M2Yo6LfIJAMnt6s3UltUG9V7TI+dTh0N422k
48oq23rA0qHc5N/1OUapNBBMSJ4GqxxmtiQ3Ssm4TsXYyLUNOWrw8ekUiqhQVHZJ
Ecvc+jF5/RBwLdboQykXW5xbPoRRDS6Fx6FwTSvzQGtbEdrhBME1r66nr4/Jme38
uBCIWCjk+NF22q/6ENan50xcs/XhxrZwI9EDA4xM4kiRQkAgNPIMcQm4h8359XqJ
OxzLJolw/w9zrEQPvKh9PWkpGk7aSTRRUHI3R7ePsDKy/QgDKiufgtyQQiuTyYGo
U4Xh6lLAnt/A0NEiXObcIChmKD7CslU343I38++4tgky2BhH9JbZzrtQ6Y/Wb5hC
jwhcwujfeWyTa49+7VW/hyqOQQ6Z4yTfWlZYxH90MXb8NoEIn4H7s/boxU/VwsqQ
CsIShQmo3M5mSQ4c2sygujSI50In3+TRrDDuVo1waNmU9hJaoPznHOf/Hft9fRY2
KRXF0rW788u/KF5XIuxxJM/Bd0q/jktf2+5MUE8aosXsJQJssRGyMpYG9s/uT93I
CbyNddWlLWz5nhumVqDVqUoLcOivi+Q5dzjuHW3qWM1Cxf97+h6AI8tFtloYvwQd
CU2R8TSEgJTqwIlTT52NgDI4QiqNE+EizDYY+IIk5u/XrQy08qFnPV/cByUMe1oy
FutNKvzZcjwLB4aBL5MtoYXa9FSSefpiHw/m3L0NzR1dEbwYBDz6s43xFrAFvp+i
tRZ03yKXB8ll0//aPEfxWvrlbkgFwLnKVYcMojyruYw1UUnzr7L1WrnsCPDl8yXs
FZ0ouAl2Bc2bdZKbBcuqbWUT4Xiclq4Vn19muqifMoJT2jZq0SMv74yFcciBdakk
bBJD1UB4GOjxsjpGPdPkTjPfdZwlZ/7g//Mv4W0J2QQ6STSwhwzw4j0dcjiziImO
5fqgUURHx7nPjxaz5Pkth2nyRvjqiHpHCTn1tIDPI34ho7ysyQnF3oOpGYAqpPPJ
Q7SKwK/2oN9Wi/WSAdhgsAkG29HnAveOFlIRufYRqv+lY6eTz/82gvg0PcurI/qB
DVKZ63ePuj4jW/eLfwQDQ+39UuYBuLw7SsHWCnOCuFLE/pG/9xklMLNLPJPKbPLe
AwWeCUVFCpXU7bXykGjqgDSXGVDERRzLCFxMNsefi6jtPCSSMnVYoRFFkiHxAq/y
FIqKcxjHhJH146PHnqf1W6CO57efTPvj8mtz5OHKyJzuk5999qWneYlhtAUqQAQo
kjNEYJktYgWHyPuxrpTGyZeI2Ay0zxSu98oVktCbviyWp6MgQxrdc2Vdw966WrRh
lPRPYJCQag81OGQfh1RNGcbqkBY/nx7zUROJjpYY93443PkYazDRJJl8xnSwaFsk
sKSwOzmhymLw92p639y7zqXga862RGg2b9/zzNVUvEM+rgNzbAXgSXl8JAl3FZMY
dG+FKSUXv4lyUgUqAv7oxM/ED4lnnip2XODwUSSYn5sr02vZQNwz2WGLeaiKnBiX
MAOpczcpvjI2fCHTPCOqPT3eMQXu5mR18I4ZqzxIJgRUntf96CJx0PmfvHewWZ2N
YgOxCeyEJFe7BMdESk7Wiq+T9or183P6RAKhpD43FdGIVaGkVaBo9tAUADS4fyfN
G4eB/DMrhWR5RNW77Js6an336jTmkYBECt9cT1TjBpy9gnqCc70blbivyfazX7ws
N9P7Vt6UODWni+OlpctlXkze041NlHgqwcZdlFwwKDLU0G5CJ2A9yAqVU+BDdKlS
WSQ/4Z5ZTBS8gOZjVTJuHZWNQeQCFv83uiX3pZ1nVDtI9JVcAinRpVhkQV0aSfqR
DBhyYKS5wxP2j60ZYxpufslDgdwNcLfYep8RfwLj15EPVU/89gHJc/eht7ZRib3L
i+pmMEJE1aJ2hujtNVPgJHzJV6INDo9y0IUHIQXaCnY0rDn9QIwfQHvkgb1n4Zjw
zC01P/S49V3ERAIFLMMIPxPNRxaZDpfM12Xse+Fy9cKVugR9e4lsM91xpV6ICcbq
LB2PEQTXx/cJW3DF9vNgy+SzIALAYnjUA7w9yjYUCIznsi943tpv24RqHslhMQrs
udk8oqEbu/mPy6pEksq6H0zjmGW5ogJL05+NqJYbAMZHCoyWHdpVJh3GFVbz6Yni
gXTqiljqBePmDWRfZtEewICQiat7VsJaH6dUJMh5Dtj41aJVGKYs3wi5/fU11Vx1
nUajwEn8+R6bcVkr2C+yeuHM3J7gAH5P3N4ni0avxk7wNvAo7PN4XDGJtVqsPdhT
6DTgqN4JBHcenNLQ6iPMWvZtWwkmAdiHoG5CtwBpowhppajYAFbInzRNK/blsL9J
vZtpsXw0dQgjBLMzw3ySKjIe9vhvNstC3gSUc9S/SdJ8IczEKBY+2BKxOoKzk3mF
E/uAbbTtPk1F8vkGhf+sebUJCqaNnTyfmLVQizGI8nWWoReM6e73Z4RGinY9mn0G
KdLf5O7vRRhtJlitMUPInRk81844L7kksrTkoEKliTaZeQJHbsc8lMMiY0eGfC0m
HAcSqT5hobb4sQGQAm6yf+iJkzrBNTLQpLsT6etFZ17q/f3zBsLpt+G1urwhUbR+
IPtZm2HFgrGduiB/7C/YgAvjjYi+WWstsyXroGDE75/fbpOWOsH/kBvme4ck+XSV
b501Yi0KJFwHvJDvRuU0r09ypwOnFp9WVZeF4H5JXgKJyTLZ3tgTQOh4OKmfDnBf
ppnHFiNL6HBldl4ZeUyWRyFZJwoPtT+YxbyWGdsGXW04eac52dDkbd6+O6MOXW0A
4btwrm++3U6yl+BXnCUP0dFTBIu5swsb9KmEyky0/Ja8Qqgxcx76VlvMAv150nrQ
4M2DdlLCGQVac/BQmXAyu1hfZOja/tOFrHBBcpSdTzwG7HSuboYD7WRMjVt9oIR7
2A6zaUV2xZMSKLimk1WFcrh8bJvZiZgjrobyCyo+yelgKLBBaAi+N66xlisJTf+r
AcK+ZK5H1YJcxUqPEr2Tyz0n8DelY1yZXOzbzl6kTzFoJWd4kYbSm9fVHMAI7Kmw
RmjJHD5Fbw6WPPso1xxPf14SAiXnCCT5kJHY0Fcda5z4MrKbpeJeHzb2+UWBa6Ki
OAz/NQmgSecLWe3BQcQdns1OwVLniUGnzwKI2DHYWFPXS3tMV0rNoYrhV5EoztzT
Ggvjb7ex9ASLIcPOOpjFxXj4Wl8hSxQv2VyB/ijfsuP3tqiR8T7YO+xs0COROJoU
iMgGJqpuy19p8BzVBFYfhT8x2lPVyqwByHd2b/4Y/dihGtA/kkcxjUINuVjaFwvu
Z4CJ96+XhmRR5E+glcWlqHHKMUAlHeFD5Qc1Ua3JTYIZ0TvZ7oktPRufpi2erms3
e3oRngW/M+2LYbF/GVBBIXoEZiRAuSk+QeWXgxK63O1qo9tA0HYGHGOvddnOeYXJ
xOpQJ1i+CYTREVFXP0f+XICB3MmAZEvCp8uP/9s8xw5/w9OMRg92x3Xn/P9SAzNi
9JcKpxXvx9kGC01l/goPA8ODZNyb2GPC4C3wzDzosKAs3a0sMdFx0DhvRZ8o4b2g
IintRdpzt3JiAeqUx3MgXlA7zb1UCZcVTL7yhkxEpuQ4Xa8jBpaOqts1AcGZ6MDb
31HhwRcfDeJszQj7SNTS5Dt1OHLVSAd6jMoxwxFCUfT4cpeELnhZdRucQ/sbigQl
PtpLAO7mqmXnP1lgtZNYowq40aNRAXW7u+aN58yEojJN/e+gJBptI2o3Str0Yk3j
a9JRld3lUNhtn73/TVatjyc7C6KtJ6O7K4/J2ITDzeQaq64kfzVlbz6R/nPXKSXP
P/bVpT0GBQrKHcLW3xQDXvCKIUbecA8C6werjd5PGLv/uZ9tUMDGNCbtWmvBv5Qf
D4IsXPGEKtC7Cgu/AZGU2yBdZPpsEb/3W39dn4VXhD4R+ORCtLrDwYUXcF8t6m8U
wfnrMm3FSp7TfRO7pt5OWXlbu+mY63umCoyus67pvmpEtBcrXj0FAUI219uWtICp
ZPoAbc9+81ymZvs734GOy8jqa4adUZBk2GlFrVV0+FQ0oKAdQ3iZvBlsHxCB+BCy
C9gsRvaYCVpbBZJlWOIoH0oo/qMPGa+C0nU8/N/aJhY0d55aWx8ytyIvKlemP7zt
AOFUnBNMMa60DaF9g4DIXvMWGtVDPKiN1oPHfbJoAF6FovZfW3dSAxKfh1nVE43O
zN1x8I8IzLM4bqY31RXymASDzL84ArXCHNw+/9G+I3SwlV5jiHVqnUA7dILs5hYh
nxhrBWEVY5cBXEBd+WpYqjRm/jRhFmPOVANydP7Im+bAbOuvl/SB9AlE0hWfpFHT
TNr0LDOe23yITktEQF1q0ZqO4qfj2jEbQWdcMu1MRLL07grs5ZfBwGflnu3w/L3O
tVw2Xnvj4cKpeCVpX74ct42JKjUBeC7LvLcKZApFDWZds6dQss+GHo1wSbhiSmLU
0ryINLL0bhihfqqHt0tS5b4vsGHfAcv9Nhllwo43QbCJkY9jqSPxBBpJISmgZeJF
5hjqk4e344QgbU+4scpnLiT4Sss9yPoIkf+QhnFJnW/MMqQCJM2cmCd0rs8UPNso
cY4L1yPWA4OLFD9CYhVCOaWyhirjsJu4nOAKBGAqavgCUpth0XAI9STDkba/SMNX
w1JiYvyiHSY5v3/KEpXsixo6iFbWKgHSQCllt5QZdWDQwNa7rtr883GXpRyflE8P
zsjn3cgj3k1pMV/7gVbiiujuY2jM3BOP4C64TAP9mKsh40Ylp667I1acOZtxzty0
yzgz2OFEkI3Ct1FV9uyhBIUs14b1KIrP7E19+gL+LNUDb9ObejKwTH2YwNOpMclH
hnK7koRcmvz0B99KCOnbwiBXc8dBfVEYZQfyNkRGsS9LMF8E3DIuiHdwLjIw7SCR
y46rd+WrkwQKlCDQMTnynylhhPiu7fQyslUVoogxtwjTIJGzgPFQ9Vm2EBWT6JUl
2tQ3yTIXGbarZ/nXBDb+QpkKlUPuLNc5Rqr6vYAwkgFfrHaeRbGaSSUwiMXVeMzB
KM56D6pRH8ysXH/hFxITCIWNNfrb6BYj37Seq5tkQYduONfaUTRIvkDIbZx9OVmr
FH7EEW4cWQdue7q01LYPLazquo2SvXEStoYfVJNzHd8ehCukHBSlfvcibIr+/Zir
0lH02jqn5iDxiOP0LZcwzm/m0VHC4JMpthS8QBhxIhCuPlB88AnAA07WEuHFAkDh
PHiX6DJKWroQR3mQoo6LbZ6tmPeJ+SThseMcq1sEixuLhxgpyv1I9i54ZHQyO8P4
1xd4h+6+msSFwMXFK0Y9hrZrGgIh6W8EmdJhu7aFQWHKVTXip++Ksxw2Y9V+qmWT
ouKzkLXyBLFJP8iZD0vI8fJfujRU+TwDsjpwF2TcKjU1/Ki83DU88VNsCQi459+V
v8lFis/HASOQpV69sgreT5BXFmKgl9F9Ns7Mzs8nbMAo+GnAPZ3qJE5Konw4+oGE
SOF1gGjVCKxxfb4cIVU3Jv2MlkK4BstNIqsDvd+BOiecQurJ9sCAXfxANKMePbWB
QCW1rkLYMO3Vup8O98gpaNUrC8wnefKKp9myg0Yh0jtfBezMD8iGMTDzZ7uDvy4r
GdHGqWTvkIJjLIj7wHYeQRrJJeihyi30FoIE0MfpvVG0ajN+mvjeQKlOd34gfQBU
ay8k2VKe3/sWA/FoM+Hbx6KvpWQnaIsyhLlfiHa32yEU9lCsjyRoSrfGfSo+1yIJ
IBsjgidNRC/IKJCssqxHWWIk9nJJWAhPVbFvEQMRj8A8nRUZXFDE4ENhtVXmb6/i
dxOA+d2qtqJUeEA+DE2wRKNp6oitMu9kmBDmnHO/BTD7M+Y1sZH5yKoKPsy0FEnf
JgpIwREVJMv9agLEAWmhgXaAupSSMgVo+jjm7QB+SY1CQ41h3Qlr+Z5sQd8KQcMJ
Fswtp5hnI52oZxDCCfxA4sdBzvBXwdJQSC8GQI2xu5orA43+L1ywadZS33CUEPvY
S3TjzsypyPcDZ7rVND0ecHz1hkdURrcUndHt+HGmMWE+m5CgCt+Pih2Xc4yX/ZIC
7x5tRwh5gj8oFGVwMiIjabHIrVZEsFmlvlInmbNoCmsjb/SmUkqo/ccJO+IjQOFX
hUdUfDMxSSmpzoOmaiQJbG2CHgIWPS4dpGN/9NuPvOi2/MLD8qQXQqCQY+Y9XGjx
q/YmVuMC/RrzN++Ymu7LHXyttsorJiKeSbl/uj4Q3A/ObcycKEVVAXjxHQwXY7z0
ps56UgqNUPuj6PXbKGhtuzhWtCj/Rduvs2tm4CCwKr7Aau9Tb4fN7K1WrYWmgnWT
Py5olHtqxpRwD9dxRbbo5Dz2Cwb+h83FwQXCWGScjdYzaiHGYZPJ/yZgFSHnwzhf
RhTxMAMeUZ/n9ainfFCEOj6taV8tS0Y4vqdVqQvLvXbYpdN5zWAXE8xy1ZUYhmpu
Yti2pYHYRFLBgQMJr71Of3udmy6nG1IeDPE6n/UaY0pw26MWEar3dYU5+kSTgzbH
oKTvT6EtCXxxAhyGZDeF87VWdYoqgxg0sImBjrhjcGWrjKc6NF1RJTr15zl1T5iX
bXzRsDZtl4YORdr3DgJVGSRlgcjy98wmo8hKExtpy3h5VRBsHykLafkNUaFPvfwN
sWTZtqNHGeebnTHjTBjHaJcxks4y0Lvg9Meqrsqjba2K29AFYw+5nxmgnKrOG2id
cOBvjrNuwcRcBeqoxt0pPNc9Xb8bvsl69r4yGNPdx5WXG7QyWPXuhOUQ+v1ddGb2
et4YH8tVQCh1hwrWilIDzsPTT+Ga2QSSGdjA7jTY8PHRClDmwfTZXfaMv1iIA74B
HoBsoF1XSKyBEH85D2RAuPCETfmv34zBWMrBfmNsMRlOjsXKS+dB3n1bmis5QxZ9
uSdkAF6APrcaBmGVUCOvtbIjUPMmvSV71Uc184a6wRmx5CzGScxQvInnD2CYdptK
ZfzCGRftadj4cnZKXasAPCpBkvWAwC2gGDbA/bZsM6gN9GVg46xNTFtGKmSwaWjU
1aEMRzcAyVrU5awh1M9wYTG7qhQEcMMG7Bsc7yb9lqG1zDd47Jkoio5kmOQ2sQih
UpUQ9PVQizhgiy2uF/m1toDV9O9Y9iZ62clXII/6WqK4DCjRPaCXYr2Prpbr8NXQ
+dpD5vcBi/O+TGG0mNYmPxHI/NftJ2k6m8IYzCb6nxoLtvmFnuBMzweRDs/MXIW5
8DAqrZFq0YKD7xfu9v9XxX967EOuuTO9tnJ6wRE64FWjeypHJeV3gCj9v/Kl4tYi
LB+igHcCpFVmgWaND+vxWM8VjHx5PlTm2YRf8ZTEy005qshcDfWpXYWCzgmGsFI0
+wuYDkgHhVt1uFYp09TbqPZdxgUiWCH5czZWi24CrgydHeJLliRdDWm0RbfA+kQE
RiXUeX60AsCgXBZ3ihuO2UaT8j1l/jKZhYJgaB9kcr03rR8Qnr3zbd9caI3KHCTU
yLvuy0FooHWBLmnggItZYYa9VOQgZKklch4HjY02TAbW9YoyrWLziTmxW8O8AHEP
zjkWBQEx7do0Ks9w2VFK8SmoMeYXnb5PnK7YqW2K/iEsbcWg8/i4Ixl4USW3cjpS
8YWNB+OUJXTzIlHfICrJJdRyuzOmLK1pEvui63Ne4UUGXigiXPsOkzVOoN/6nrvK
JZyihDzBPCveByye0IiWxVMHYgcualKf/1MZxcgGRm94hOp7qP+CYYlycjPk/tGu
rUBEzUsyxzdGlfIOg6QXr7e4iF36XUFV0xtidQBuFU0GSUHic3XWcAOwRFLm0kaL
Wnf5vdHu/2hsZzig5oPusxf/GUHGaw96ImxTO837Ofs66qKAi08PbboKyi1wfHM9
1ZZ0dyqf245yw0Sn9v2ezJqJmqdwIeyKmqkFt60ipSVcQpzb4mlmqVmws+RhrElA
BRFS2hc4w39RmR19H7Mz6710UDcVAK2Dcg2/9lOkGzhPv4DEbIj9m0yxxKhkITJR
JxEcffEgKIRclKVQ4F5hH9jrr4nlznTwSwSgNSqghoGvqcT2vrOjBueGG/2HIQ7l
eF8ijM0XGh1pTraA7thVS0aAHnuGEmLWHFc5KJpvkU/VcfimUPDJgS8O2rdlJHLP
V8C0kkwF+/kyAQ0+mmuBAjJa9WzBjL9Kkml7K4ApGYg1KSqdQceZMl1oBC2Evf58
LxWo7ze7KWgh1oKl+5Q7E49U7EdRlxp9NY+K0u/Q7VYOWA94riA7GRgjUvPYUMY2
a1CmYnmy7pOMUp3NyhLqfgCwk+xdfzbSV06CtFg/cFE0SLY/0LKUnXRPHp7QJ/24
eYSzcmy7lhVWpJlnIpYUTS/ZdzOTWnpoBMFEMcgqIJ+x5Jsi4UxWkkQ+F/cFl2Pp
yQ5AtSpVt415yubI+m0aO0hbf+RNBMM43ICQiFXvuFfBnMeplB/cP0FbMSlxDpc2
aPR+dxOfK6qMnGhrlMMR3EPtl1masbwA31jLHk8biu9C00reQxBawoLNj09iKFFM
ENXgo4t14Lf295j75CEasI7UMYArwjyoGNJYC9HZd0W4AjuppfkscQL+pcrNQ/sU
9bo/h6V2uUX2vbVd0LW7A6J2n1YCBTjEWGUFTxpjQ2wc3WDIDMq0QZ+ekgYJNkLi
Lvg+Aye7d63VCPTMIvCCZd2QRlCuNzBW+6BizWJ/8oj8CcDN3V1hCh+pP+KZzF/U
pvBsSnU6MOD5e5RC5N14R7eoTZJDhuq9REIcwxs3iVb7KKAylynuf0cUC58UvFXe
TkR/mCKemyhd6EAJcX2UPEUnLyBCCnycY80yp5gp1OL8BFCF1kq/lfJDXhYsZYcu
fX3G2LmRNWMXaUNXMt2NaQuxtKqDF3Ye9Q33EVaOitv5XX45wTV8c2nfTjWVbs2X
3ED3FpFEsl2rH6EjGh90TwPLq7lJTjg+QLBKLZztqf96OcjyeQimGfWTGF+L6f94
YveUasMM8GUJe4dmP6Gnt+5s0UHbF5vCKDW65KIsldR7ZkOQaUddpkQlQHtZlygO
QPs0IXSDe4TKLbmKX4XOi0wP1qBE92mj+gjbjDvD7/oAFh7WbhMPnb3FgJSM4G2Z
iV1Ax35DOpja2x/dIjYoOxisx8qUo3Jhiv0M34IbFTznf64fLQdpRh/FB9oTaJca
45qwbWhnQS+aS0eL/j0Qpa9deP4R8+ocpNhDKsLvYX5+Rt/DwAY26AtJDkZHgxJv
mOCT3Q2rzKfkyU3BXTEeV5ETLG9DPpjmlGuilf7hOkQ93Zl20G64QUDNaN2pwYBc
ewIRrsInujmtwd8LS0aqwGMu9UjSxl9ek/TZev0NUuT0LtKLW/v1hx+LJEk7Tm5X
CwV9+0XDguLEelg3rhPPdvs1RV3N19LeVGD2fke9yiE=
`protect END_PROTECTED
