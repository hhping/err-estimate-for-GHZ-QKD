`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HGcBM681eUCyHKRfuN/m6t6TkI//veNB4D+1XImvOpWI7HcVQ7hQOvMGzQn6Q7SD
1XnZA+r+B+p6WMKkXyR+lyKdVIrD5PBOFNEIWpXzlEWkHu4LUeDi2Pk/iJcviy+p
Cpm54OGodTciFHAwGxTXZ7xwv3eKLXFuw1+0Xh14llohbt3d78Lj8NibezEGV9bL
XTLNh9r47fbEcXPubHKGjGhLKOUPaGTqGLdwWmzFBRnucNJUq5jxrc2JGh9wv8PV
E4k6lkrgqQGLAIlJEVZ4V+LhIOEIgFfCtFfNeH9whwbTeOvijUmuchHCgcyNYY56
8ddAFJ1MW/wz7SfNYAeccpDToLQtvmvgzXjvZD4tTr+y3R4gy0IhyhZJ5o/8DBfn
0XPDbaRUnPaqbj2n+xBICa+xRE+TO/2icQRjg/NvsjVB0Kj28srfC80OPVYc5u1A
WHyXqNVAZzBL3mOGZeWOa3LSAbc5iL0/X1iwieiie805mCbTdU7LInhoxSdBEqkf
fS3HpP2SH1yaVB9y54Oc6exRfYohq0wIuwtHd/Zf7CRSxUmMFBz+sP44zHRdYGZ8
+N0ztwzUFTlPyJeshFkHgonxmOEIj7rTYm9WXM4bxm+Af2j/lF6k6sRI0mJlaZFZ
JOmzicOVyc2+b/GPMzs0kSM0DR/Bq6jVaId5ZvMdIEEHVGXqFYr9qq0062lfulxw
z70u5EKDuwTvx6JmP1etGpoLT/JR0DolSpHBLzh5T5EH3Uu5tkfEnOdnGB9GRlJv
xcmRI1CJvopu9l2Z++qgYTICw9fg9SawQzF9apnB8qET+uHOnD7sAfy085UyAilI
JLDSkfjaqt/Q9RdGRWel+jGcJbDIjnbYSt6un2T66oGjwXl698iP7IT1t63SdGG+
bMJ0drTDCQbpy/2KtGBCU/kr/wdKSaMjxnZ76I0dnmFZSjZOqBKvEpyGT/cB6pjr
oGLXRxhC0Pj4sbNjuna7+9CiVUdRiCjFBX5Vjdq6bbkbdDR11IQpqgk232d4+RLd
S6exc6fnprYMnsgT6eeMiJAXq8WFvnFAsHvASQcyUZQjJf6odHaAoPO6yEG05hom
S4EcmAG+OTKsx9MNPQOgpEyLclL8oWFwbu528R5hdGWhP075rEJmoSS2za1JLCdw
c2hq4IWS07ogxtrx1fQhkEKcrg/5g52rv22tH8PXuA7cTGrP/2fKAdvCZLofEwOK
/p1EU0uCk3VF29Sc2AIeAnbdCgLpkittOwH7pFC0wT4daj58grzl4B4wHWCbv05o
`protect END_PROTECTED
