`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z/OXH85GCG/vRvFp9BJTDggO91KkbcFM+NIxJ/6LRvaqolQFRwr0PI8LYotLy7VL
xlcSj1TRO+tMLXSMyBbNY+YR0drjujao9QPblZMmm65EoYfAAHhfuplMtHZTz33h
e1vi77vFuNPEvzv/d73GKUQarqY6U4ff2bgiFkoP+aKgh0a6WIOyTUpRzs18gEx3
FNQdrBHUuHIo0IJ2FiuLEFviQjTl9zGrM+BujJ58si4BU+r2tpXo0DsmdSSTfslp
dPfQmzx+msiymzbCP4OiyMqbUL0WR/gEvimNe0MNRUX5ADOhPqZyhWmasutHS5RS
TdRrVPDSyfax41RvxKDX0VofOeJlt0clguZwEVaAGr6BfFZXZF8gKWW8+M0/NNF8
Y1eDUpUCGo7VJalUcOyTP8be6KzINYLJO2SKgjZbxsV6W2ny5aXHytRKmz9+duY5
unPbMij9I3tIwi2XKqvymgEGHFjd3sIkeEEYpQkhhMwzpmk4lPp+CBJA9il9hIG9
dvmVJG/dtbydTxIcA5nQhrTLWu+0Guwp99j1Qb47cZzHLD21mE8sHk7I0EZ1lBNH
nnANv71m4czWnVkwFlwdyenLPBw9mu8WzO6mrot/dtek3r1L0zVrYNy/L9A9JQUt
c66/Q8xV7U6EXaU5HhuDbSti3hzjJBR/Pw3o7SLjBXWupht0RE/UD0zwU9v3MJs0
15NdbftSeOlw4T2MTTmwLpJQeK6KgL+R4gTUynwALD9vIvBeEccdsssx62l/6HtB
7/sVuVlM35M+Il+qO3/a/XUMheDc59jBTWM3ARAbIssss8KkBdAPQaZwMvyUOIzd
r72JqU/b7fQfETXrllzoH3mxmrKReiaT9c8X/rMaF5jcRE5VkW/QvjD3Ws9cb84J
RLpcy10/6j8OpU9u0WuV5LjL+AIypBddVKJSCsRTtWZY7TUXBLYa56I6POdz2sZY
JQfkSrS8623KCjQWRi6qyR+unfU+VG8wUgNnfHOadUwKa0SgBVv9UdEpUQX2woqD
jCEBK3IzGIn91cNZNNYp/msaIG7XvHnppzTleyweiqg1evZxMGJe/sCX4DBlZB/y
egD8GzICULZCJRGCY1jZ48Y9oTD/Rc4QggNCkdTHvv0pwlj8mNqFTW5uYSGwanyX
3eGZz8Mk0Tm6NRIm2Q8EMnWMsWTpXl/dIgbxlOBVAFe+J5junHF5cD382pxhiFmI
QivxoYjZlXYhn0yMi0y7deJgyQFNWhOM4roNc8lmBWz2HGcV74Ze1ZdDoPCWHz2V
2VnXnfBHjxsoDVlpo8YoNhjGPAeUUPCO4XE/yxllgNajSWphhYvWlEGx1GNRwrZP
Ejfwre0jqtLHOZckVZrkBjCVqKeEI3WxJFaMg9vFZ02JRkRnovOG+KbD6JNQwVVY
/5ffjZVQZj+wZIUiqclxw0xzjzD7ydTgE6Kg0UFZs/2GTaQRZNujfuCsA0san7XW
MoYGiZU3UEHtsjWvu6iIWVCv+ak720W7GBCOknVwbp0djkEj9vZyxQS7PS4H1e6H
9xJlirCCfjzcGkcOkAoB9HbFVBpAj1Jfcce1vTvTROI62Aw2BXFd3vD4l2HEES34
h+0C4IUrXsAX5784n4wAibH8WA9l+T59csrKu9aglfCTjDBbTBxel3j1YCBMmGhn
WS9dDagWzsJ1JMrNb33bv8nA7xQqh3tdVSD1+f2Wm5LA7VOt83EI29cnJxXMeClY
vFmkosM9PtNr1gb4RRHAR1hSLNm0sBnW6qsr+16I1LtglNNCSkhfY2n7trDFQh2i
1O/o80otPDUWOKqajj0yAJZBsFmRxZNRR/stgOAVgK6X4tlCTR/nuPjc8j7xAS12
uh9rxbv2ybsK5zjMZk+QyujhID5//fKhG9PwcqftH0cQH6i7MAZu49DehtfQkON5
hI1qJoB9vqyDD4Bd7hf3e0AfTk3g+3umSnsExUnqu5JUvBQQUHxgPGHDgB1x/TRF
Y1gAVaes6FUBMa+D7lvcH8HKJtuSve7U2EWITqSf/VnbtzMS0kygf6+cI1Tyi0Mk
h2jllWjaq5PKgfEd29n+XOmyhTxy5K3OPDB/PVlzOOCQzu0aaRB/hm+b7juQPLmM
jGSntGbMw7O8JHlSoBVi9iEH6ntmDLdhWUx3C6xiMNnDbu/wdINjO3YW3ZIh0usQ
dKFCMfXkzsNUisJmdQvfawuAFLXKSjH5C3HcW/fs4W6IGmTQdttA7WZfgyZwm592
xgjKl+tS1L1V+r1/adds5YAByVkhKpY/OcByF7kD58+7z0MegRnFmLWU2TejJBEM
0vwpSsX6fYPmxU9F3Xze+6RWjpLS6GkuuEn4Wpuy0ZTnscmA0vA4SZi5JpRrcRDl
396qOCpfj0Yf5MMB/of5nIch1P7S1WIcSAvYbDkzvdZPr3AdC/9kPx8VTxkJ1CDE
cWyeTclR0zOO0TUXD3mDcr/EBEKZDSiSxOxH7UHk9EYlCVBQzlEpzlq67Yalumd6
D02IW7beJToBsg435hRhYoJFw7O/rWXWFMBNOfVSvGc+aPo7w3PNPGF96pCAxai1
guMX4cIAISUyk22QJzhdciGhE1XfEtVS3ZbDjC1QJ15XqL7XS6gb74BQ2cFCby8n
04jM0jLFHKib1D/ikslF6RucoqLddb4drg51jycuu7H7uJE4ZD0XP+fe+8WzMjAg
wMRKW5PUW+KLqQBDbpAvB0ZTSnePNk1DQr88Wr39Mh/bVROae5D1dXAabCM7Ae/Q
V/HaNDT8bWhh16LCkHTQ5SIwbPP3xw/8KQMgGZq3Hf1VmKhy1sUoi9KIbRXOtDOM
5UbFpr5xRcB7FnkpsjizlOOMOGRoL4M4EEIauQtMYudKqw/nKjRx9wDdROEVm1+k
xzwtwO21NtR6XK36dIsrf8hvAH7uwCYFLS239nD0n6DMxcQ27735h/eHDkTSA5Tz
eFXD0AMJMZjQoPaNXKAxUmVgvqZorLDJ+8wQ4s1UsERX6ly4h1b6fV4ibyUOiraL
sVAPW8hRUFGe5d14GciaVh3T5wDZfRXklkmAeUvfAjllk1Yv6v5/dEM2U9C6df5G
WOTV1acfntFBMan1JNNIFY5b2O+whiArZzFY5jawS+L5YIubGGfmUyVLbbnCpoIk
C6LyI8lD8x6oZDm02zRGD+VlCk5N2ilamEBApL2hfhV5b7e7Ea2NwEyt7txYaXvM
xv9oHaqR/8yYXIUAeCZjQuMNm1AEQpT0T44WgnTXYRes0cQ6ks9GyoQIygMsUOmH
RyZ9VxjWzBy2Bye033KQPEdp8Z8+/iCYnM46x1rizt4gGeK9VWFpmzrXK8VCKw5h
Knu6LesDyGCWHav1hbP8EbtUH4Z5F4igXZ3nptfcYCrsZXJhf6r1F1aQnlGbqTJW
aMafL2YGxWb9nb8Ap0QpnndtVpkOObjDzUpIvSGSKN5at7WqbtUQfZeEBJng572e
qs/kpAytBkEegaYGySCMKUq7X4EuMVigVzoCMOC8Wi+gTyKL/4GP/aUVS8rOc/Dl
VeFkp+f6M9BUQ5QzXGiqT/FDbtkC+aQVfB0tgE1uKIhI3jLGokVk+nm64V1kwU4n
3rjYAnBC3YzuwijmioTRZ2Ox1XbQ2wxBFna1AW7lcOl/u6yz7zlhFRKuTJGCc4tT
/ihCo8/FFTyl3ecJ3XjUIjd66HNQbjf/Ra59wesgyowdocRy/a+4i8MR1+P1zvSj
yqJmydD7f1jQIUmhKXA7SA6EexMT7Nd32HqoIqzi0eetoeWdwj5HCHnVBB1EJU7M
Dtrpwr2b1ZN7yaOE8NBVpI8PxLEhYMgdLycwLwApZkgJKjaVkoLEAZeeafaaO9DL
rL69QRt2Tt8dBSWYoWR3s5z5yfYE01dz/HHes8mFWueYY2KmwfuHr8MpuTgFwbn5
lHpRi93CsJ09252dsezSE47IM+KiJ3r8jtp42WCUTQ37oy+ISGXPoImTY1EC0INE
7Hi5vgdrY3e3GoLj0KQ3Iy/s8+16aq3GuCQ7AWqVYW7Ew8oaiyMha0q8YkmsZo7h
msA0B7Z0k1Fa/XiHyuViTg1nP9U/OF4a1NP7GiEG9xlC5YbFWeo1jQ9V7BhsZpTf
w9IlVBRaH8JTJjJN9MUxEyzVyZZbz7x8mDLFEbGtLojYtIh0xKpUpBKa3Y+zVDbS
+2I9G5zzjHT5x5P21BkYBpGsP2GRQc3GHEm6q1vkS9nAeFbvBuU3CM97zxifnUKi
n1TiNBRoYQyQx+jaidaPg88tEr84m9qX4gmMEJNuRCgG7SfQd1quTZ7LaUvftsXo
Z9d6kBL3Bf/M6UnxEkpwTntAG73qDJyd9RfJlK84xRyr1LL/1+kG6oZui0nUQkm6
aDdyyaDNsfG4GG5pMX+w24zLwFO71lYCqQpJ8dCZFV4PMnhih9CpyumWEQqqxmw0
ywvNxijpanOJshtaJ4Pf4sCsRB6LhqM8HRKNSsA07Y4=
`protect END_PROTECTED
