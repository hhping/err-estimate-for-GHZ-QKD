`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YKnRn9tmy0Z1G7lNs208Pqh5DQ4x6VWdJswWznKlG0CCBU7V9uRfi4Ae7fIFX9Rm
5c5U64c159YmGQMFAWamVJOqu3wn2GNV4SVHIeBGqddMhNUeci9Rk31Hw1PugDRn
u3wa+Fp/C991/sfOtn63s8W1f3D23d5KvhR7DoydhT6iA+77JNnnjTZ5H+hoHUhS
6tn5ar0auBNasqyUfouoHK9lLRsWds1Vf9rO9Elojj7qAUQ07TpseoqFpLyHGJx9
WpyUGWKr5tE6+QPB+3bFeU0dZxqcPc9w3xI/7kHxBQeG0/w/b4IQOybfp5neGW5s
Y2YA0177aCkJOu/K7zd0Se31bF4unOKgtcZ6t1xULirg9AvrPia/ICd8PanlNIXH
RTWGcRv8Hl512HLWFUqzM7BwQANr3z3MNbim+lmdyd7ZNlv38yHgEGrYci5+CpBl
VtVMrrhrJ8+Vakf2RLg/dNJjKagB5S0qaduZQ1LO9S7Ltjr1IS9vAJd9aWEPIisn
CzA8shGg9JiwQTYrqOXmN6jCpt8g6sifGQzF/5D3nYScTY9ZPHHnigp+9LG0SIAk
HLand6pmtyEr+sPAOYuYPA==
`protect END_PROTECTED
