`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gNDyvL1UnG5rfczW1r/hUxqn4ucZ/recFHLE9A8tZAKpGgZ5yDLRPtYvptu6GNuE
PdYck/67/RZMqUrQdcKL3/uVrj8UO7GkYj3Grn8OXHcv8052lUJAdX8OOOCbV7Xt
spB88WBT42ZJ96PEDzwsmUf0znCA5zgywblj3XjcMdRq/dLXfKTeOqAFkj/XbrgR
UO/rGJWzsm1+ThqNg9OC8HmQi0PUtiWwrrj1XL45j9pevGBpMkR1R9c40GrBlFNu
E2E2IhALVWiiXtbcVXsSm/Y/aVzcz+5uNzRwYD+p9DxVpY006l7TFAInLNxV2Xma
2HbijmkBHHhQxsaHT8P6MoW7dtEKCGByEkB4ziiTgU8GkTJbycQ1B+N5PAvEmvM5
BDrdlLSsUqDnHjznfYKJzfR7GRklk3+K3zUufwp5S1SdXG516JZzeOaJBBJTVkbl
YvsR75wFiD5O/tdvqQEa4gGHNTE4dX2zje4p5BUYPzEWnQd+sVPbMXHy7w0b4XCq
ACEhPPluV5oUIzruvYUmoUfyABQ3hM8BnrZiOAzQM2tMvk8gUotfjHlxZwXMt+FD
WrckcBY2LsezvOEBx9BWL7Y93xsdHCZevYeB0Cf3RhYsmyRfaCg2H1bnvIv+wAGz
`protect END_PROTECTED
