`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jgodkNUm702glcx5UfEf8myh+g4qmel0QRnOGooAHq3xOv7XhyG1cCF1G2+KHrfm
+GSMhi8IFhPkcfRjwnvlu1fPZ3TyHLTQD5W5UJniFFVCbXl7VV8tZsyjDTtllEXP
7f56KAmABWaC2pl+wJMMdaSGuUOGqb1S06W0dI79oNNaUAT3LVLzNw8pUMMhnlFr
TOmRvG9UDveeG5xQGJWxzYz1qE9s6y7y8YKaTDQaGCuVd/cf46l7pN2QGDVgqV2W
yE9kxmKapekWYD5VkV357X6KMF/ZCBuFH+FhugFXZ2KdZA6jzHL8FKtr1GPosSLu
GbNnwcU60ax9FV9b3pDb3NOBvBGpotwBhUOWWGFYjGQZqrNDpjD43c/qCGQAojWb
BbaFhWwxMN3HLk5960803GabNyiP9PBsH6yijdf6GHi8TItLtGbzRc9InnvVe2zc
xKeLjkKNYp85GgQcLMAcjyCQVt2ta755VoKzheiZufa65YoDViBPdidEgh8OSPXO
XFvfqBBlcB8P/sAOfWs/gi2K01BjP4PEcpbGRlgOJo+VFEBzZjPgjbwofZj7zpKo
bSIpCz22cTJlbbI5O4uqjoZS0SXFCHhYa/wuUhT61If2/E6eOm1T3bWaUgSM4OpV
nrudOZteBjl0ivW2mSgzl/DfX8EnvRZKDgxjk3gptElqxDdOcHSpjGE9VYTTNIH/
PO4j9WoPpmfStnk5f3bm+8pH/ttQKbLBwN544g4ycXDBFcyJ4JMcvrxGOakSVIzC
vB+K0vK6nL48j6eD9fziTBKoGlTsVKEdLwSUSr9yn3fbrqdFEzNI8pAsyvNTO+SZ
PReCqAAeb1LfsVVkHW7WC5+l+43+Z44XAz4L4nLQlXPnJBcGbWJL7o2i+hGVsrnl
pdqWRNuYM8Zfwi9VbUOshFBgvjuK+0aXelR4zIETxV8QbAobnUvAdYf5HnCULeCv
tpa8rluTI9rPw6eoREoAtJG+v9ne66n/3+pSzkeaPogYCWCeN1palJsDsAOli7gb
/UizAOjbB5glXU0d9ol+fni3+6ypjryx+buR8rqm2JGXXNFamKIhVUEPSB7z5PgU
gSdmJZK27uJw3sAUenhEDGdTbUuby35wp5oDGVJ8brrcy2c7BHeuB7S+yUTi4Pzv
8B3JAvhanApC3PgOgoFe0kwrJQsCLGMJQxrXxVQCfh5AwlGkirrhq6IDQzr38Ppd
eLGeb18K79eTZI4qgzVrXGZN0H5enI0rwWW7hlyua1YqsTEZvYATNmb3Jo2ARmW0
Nx28KWSStJtGh3G5Bjbh7MNOF8lmyO1IoV2KIW+ZXUDvsPvoVvcCbaNqpyfaH4Ov
jz3wKYrcv5AfTMRDcYs0ZGF92FtxN2HFH7xA8YsMzv/Ouorj1aKEsb6mrJc25eJn
nU+hfA9MIHTH7S55rccUAMAbzEM6rz7JI/yp6w4BUQ3Dc/CuthzLeVuSqZHb2Xzo
BwQU+UjP14z+iXdqccJsqwrr+I6U4QCXBBWIsnO14BPkT/3eZwl2nYb126Fgeaqq
mHxs1oKd+PwqdNY4RqTjvIySiFJSpJqNEBFf+QbbesoSjIwOmCk4C0itYXls/KFL
7lwAmA1004EXRWdVdxMGt3BG0k9/30PqDRNXzq1+idKFdxTC1u4BuVXaMDytYT42
Cmv/X/US5+/npgjV0FRRkh1dhAAmqk6d0oD3sH/vq4y/+62r0mktCqNSgbUSAPph
Hlkkrz7NzoNoNRpF5pyLohY6gcE0JPx2rVlQ0ovoUUerRFJ5qiZ2Xfmcv6G7VmfK
xgxs37jOQyuOIIXgm4skQdNEzxO0jwFsyBJ9f7Jw7YC28HkPY9s5e75k3wYRcwMx
wvIXVv0kzwXZOu9n3UotSXZC3vk5gQxketCmMFJ3oCP9baOiMyI0r98vY0qjWpiV
QW78J7T9ksn92usuG/X4I0rW4E2N1Q/re8rQx4liu0F8JxMtdjFgFI30rnpafKw/
I8dQI2xYJ0Wj3Xb3Gf9jRzSxOUQh0SHNDYG4wIx71E60jKAtsK+U/q32ivE+UnNF
jEb7NDdXHnoeHpMZ4K3BL+KDosWw2GjY/QGmcCUvcIAYm5C8NaR2+DTpeTclkMtM
JxpBgohoMWZijLSE41SvhyziqWUoqduzBqTAj1WQXx6RyjLBxLAWCe6m91CNkLKx
09x2MMmPdvHBb29wOcXzXWxyKQy95eEN/z3c1YyIoS/5f1YeX2Ws6hzZ5THFLROC
VptCyaDBwC3R5qtL95wLR3avkopU+gZLfVLYXwzibguy6nkbQhReJM92wywd3z5W
tHaFEXJ6Zqe2GWHnr990GoKNYuNk5hDoGiPFmzdDE2y1cu4/NcY2e/euzlgXzzuH
pUKLAPjz6/xk46YY6ok4umFp3lBMblG7H7bsKNN/31dUpA9jNrODw2opdm86y2XN
/lvsK8aRBx2iiPIVGGocMaiyupfct5e+YrxD/BDsKJ6nTnKa1bIc7BhON7GiDRwk
tuyfVh79Wyv+a5HesWQlb1SXvBIT/z89Grpr4RFZOGCFk3IYtpg+MSXYTUmsjrNR
1qSs5Wtzz5wHizdpG9z3dtI7ziEiDqRd3TU4V8hHDzuLhU+CioX/D92U8TCDXn6Y
5XfqH+QuPH5J383qhjMGULdylSKxgFFlKFzdPCOZDq6DBcDHy+bTiXIUx7re/ivp
gp7RUZ557+1bphw74EvhWcv4mCBpUcGVARbG9EM6SWSn5W4TIyJnejblZFn6cTPa
iSuivNEc2lwL22Y2bMsd3IpF28lceI/1PwGJVOWP+97Gq9c8u0KfKQwNrnG6ootk
HPKDLcObFJv394X3Z7R0oy0lUf1mAF/JF27yeSOftxBv0fAWaM41dfjaVmiEJh6i
W+kBR3UNAI1YezlqMBFm6yyveAECyrUcYbEh1FhQzjfIo+CM6NzY+kG4tfPZkdtO
5p8U578hNHWZwrs879dAw5tzqOgKS+Hb6t4bVsTEGWQqZUaVGZwzWeYtRjs7pCvZ
kuvcVx/4HcuWeMf0+vtfMECK1pNPdFLAi0d6yyfJTQparQ38iTml71ly6W/bmzxn
MyrmDmsuJDHMYjaH2aXuuRt0ujklQh2agvBY7Hy2IQLtNvx7fVOkkYIDA0fpt5fB
4AE9bVFbn/eJnDL3mvMVtGGtnwMip4QXvt4FaNWFPeJGoJ7WbDoqUE4/71UTyaZz
M+Qtk4vZgnb7edd3a16QOHMz3b/E7dIMIMx4a0TVd8P3Nuv9Nh/15pKZ5gsJUH0L
/gKRmiRgSQv/cz8TnjzvSg2/aTZWPJA1rXRHPTntmha/mq/JGYhvPxsnYiIiHMVF
XsR+fmy+7EEemGjlTElElqmZTBSoXoR6ZR0DzghdKuFKPRkjxA+yQB8ASO+D9GV2
KJO86W2Ca6OGbisKRNDdjDse5OdzkqaA423MlQpXR5OTQmRX8bS1CiEfbzZQdu5n
lGqWmYIrMZwrzry6cl5TqCjCssSMqt63JiD/w4myvEoeOHzY43qH5rQkZiI9Z7Z3
uFBsNyUj9ADmCjVgYIArLuN6CQ/93kxhc4B0XLSY1f5Rw28sL4BNXUg7BCKhTlV5
dZs/63qamvblnYJ9XgJMC5srqHqOwCqF+rR45WkT31STDLE1pTYtdon5j0lxXalZ
O1qswDrl35+T/GwnPiUBFMgbvGNHtqxhWmIIZW19UaDrZ6Ep7rqk61VtRkwvZBuB
PCIst7AytSXmkyQaMV19yOR0w5zwdEn2QL9ofpYbw8J0ZSPIlg0Mp7740u1Nu3Gj
voQYKTvQcsuA+vpRsBFkWHswpRYUZ8QuGjcKyJ+Q1vWXWpsZ+WSOz9eiFsVleiRU
AZ8d2MzQlr6982Vu4l18ZLTjzPixMMxczV/OLam9hbX6Y56Yek8lLrblXaSmTi/5
4JAdJ3t2Q4r/hhedp65E8FOaJQwXz6p6eTJyUdb77JUcmCqFz3f3e+6yZGJbP5MQ
i6uETbZSAugnsKvUWRmALkSy4IWpC34AmMucgBB+x20mVn5Sg2mlwF/2x4rITZX6
Juyh96qD1Eqat/94kwjYBBX2mHcxg2BBUGN6eqJiiwMk3HLP/3zqpfng+R/Vf5LY
bQiWtTy8QutZELxIqw4NA+vd0s2TdsmUSk+PjSMXvu3W3ex/vyHL5ySfiAudoDAJ
To7o4PjwPckV4EGe8ibVM6mPB2LJ8R5ki1ik9RH2260MGcWpkUP8Do/M5RTqERZv
3AcmnFK8lZGLMdgYFI5rgzD0S8FcPSApWg0+jvz+52D3cwD3htJnoqoMH3noo/SX
cw2nPVyfju8yem6BvGm1XoM42m5ZTPhUMFC2sq3iZgSt8ruwnNnwXjXokOPpnJdi
qXL3EYagIwl/5TJksgmF3wHp3J87VOEHOsyTqENtF0SvY4nUgbc2ygUrsBPj9/o5
LmLwYnfYq6Q5kaEeY+WENtX1IEPDkns8+u5p/+n4T4NQXROTeFonn38l2xBYyIst
u6zIUt8qy5W6uTz5k78KBi51kxLpLrREzDjMWn6hqj/84VHLKz61jBqF3uzu3n03
eStIB9q1SuRjUZqR9axMtQ==
`protect END_PROTECTED
