`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kGunVoH0+TSmeVULopY5hUbt6kt+MsR/1ytzY0SrtngS+r+U2bOyQ5Ac+C8arSe4
zYXrUD9c6VSrYLyN2u2DLBI/WlAjMvzCxC4njBOjQQ5BHC7cnVr5E0Mo+mKosy9s
PD8Umdm4QfpOX6T5qPfiQPvP+gBUFSRmZO8KFaiR9x9AXJHpW4wdzrrXLQDpEGsi
hfmuEe3s35C/mrMYNSE7p+83IFMOgjVjCOE5GCX+LOAND4FGge+UOGpi0lCpsxYV
V7jAId49oQWuTEYaJyg2SMiCSSEd33Le6kXtBbCQdhwGIO2FC+0MtYfzK1Cjje0f
BunnF3jQQRFekhrq2+fblY0/fATvoIXS7G+opKbpaAOuvDPfE2ZAHjx5Jz53n3or
FM7FrUQcKWcTh1jjAsGFKsIgXPaVGN+TogthRnuMdtZRO4IA11NyM64ItPP2yZTm
DTn3Rxmw7HfK1qy0e3PUm0FNTog8yFFV4IO0SptK3YUmAKpDLVJQbry5pV12F2sy
NEVOeDDZP1/VJrdGoOTqS2eqsnZV3nzFEmOpwMoHtE/Hl1MyfZ4ewDmnkpTMXHdG
ET7eYXO/YYa8eVPj4ymu3WMwSpD3QryptVhzO7FOz3IsTrG6lSItlyzauB3miCKj
IVsiDMKP9fnN/URAdmmvpGH1TX0POEKtqGzDzcC6DaxMVP61iANrut2dthNbbJw0
ApFN8Q2yMZMzwl3npMCC2DFP6Rxv1q8QSlxlaUnq3bq6HndhhydNX9wVY40TNrT5
adfadKuOKLe6p9QvLagAGaD5ZpwG7B7KsspKXpdXOgsfebpcrB5TfwufD7EUUYHw
sXRv1gNn/iWGnqP3eqM96NGe3WcaH9DaDD4pEsDVNpXn73i9HgZBDyyFuikk6zZ5
g16AVTcpxsnolwNy508u9ga0qjZvJd394EUpWqWps8yQ6+50Qv2j/f/d/tS1PJXu
y8v59gtwDLxHtbT4/nnO9g==
`protect END_PROTECTED
