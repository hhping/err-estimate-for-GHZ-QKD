`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+Ee/yCcTGmU7O0d3U5va85YfMxfEz2bIqqsXHXjZ1EavPxSEtLA67jZVhfYcPgjS
o6NsB2ha1+ofobwIQjSCFNdu5BRUfrKKinxj98DlxgpDpDqlRSFOQ4bmBvqCdI1n
XVHqdyYr7CzchwGzW0u1w2R5Sfxw9fS+gSlNvF1ihhtLrikVh3VEctXCw2i8kiwA
dwXiLppVcEuqhMj3ILxHfyofYMUjvG9kzQbYwTqmgpzDFFLZdBbnhtEZ7zqHdRc1
Un49P/wANkLOwB0wvMrGMx7AtwqHQBDxd9kTz8fmPn5eamHYWEmOXCIg1ox9PeJg
xF4DdhXiVTeTpM7Wx5THBuMvHLKqi3lcMqR14j6cFof3R2sz+C8/kJszE2+HE/cb
QbXZCQqeU5ybs8cDu+U5UuR1a7L7EHwVNanioEMlaciM+077qwSDmmZnrx/wJ070
ks1jsn9Xqfg/5oNIdKRkE2szSJd/a/XbJXDFzucCGjhV9WxUQILRKG28P4vl6p/q
QP7qqVztr9D/YBg74ymNOoJNB3V8BWt/HQ/0Q4r401iyPrEjHjNZPIgcWQb9cfmv
9hYCs2okyVx5Pr5grb0ewlumUAj8A1qPbGizN5GVI0p4Goi+evxpBJFTIcEJqFEM
wNnHtN7QJrZzWObLU+RFh6vPIriX+9bjbM6RFxRi2k2Y+K7ZuMrzMGlNboVdi8w0
4PKhYyH051/qYs1lxbyhuKFDs9M/sOwFKVodsHvzHLirNWkP6yNo074n+tlXcAtF
2gxHLoNdx9QWI1E9U7n5tSENVt0dWLHqqqsqchPLJukhDWKObxcli6f9KDr/DNB3
wVRGYHsk7kOAOng+H9QnhL4b8Uhp1SYJI2AwL4j8vqUlPFNVjPpyhELYVPs5qZXi
e0ubaVZ7Hysbal48l2kEflDOPN0v7hkjkX7g57PW+eLc+Cnf3ypJDfvDiy5wjijf
Sz3QmghtH8YPc3swdLY6cyTvFazjvunS5LUKwcEE9DzUJ1Vxbieic7iL+8qJsvTL
tUVa3vBtEK2slCC35560OQuA48GP8XJE+NFuZKAJENTxEMYmv/Acxyz5IQaCtTUI
aH69viCPfnG928hjg6pye8Gn4OAqe1oLwjTXXTHqC6N85AJikSWlSZgg+77Mfgbt
YjVyGwakY3+vqwmHgBj0ATsEXq+ycEd6Y8ifLhTL1jGdPxf693ioCMHppus4Bpph
7Ntu1x8T8Eh8RfbtxDx8XJITWf587GpeXCrDQo4oPSspKQQxhPneqErTIJCSv07C
TMWtxhEt7/DtOEzS7EWgFPEY1jlpX8ZpneISrq/JF/KYFtjUXRZMFmbclV/qYtTt
Yf8b54b0aIEi9huglKAoZhbCXUQHX35UkY/jrJJwOE5ap+EnnTWIjYnhtHKs3e7v
pDvrAKsry9bLMrgbCsjujTdFA2U3SFL1R6viw9yinsk=
`protect END_PROTECTED
