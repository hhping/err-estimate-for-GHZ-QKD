`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ldwoMyKv5iIVDCRNU/Mypd3MolmBDrKOU5ZaomawrGvt38c1IxbInjS9cEwV6xaS
YsrSX9/5XhoKpVhI9vmqYt5w+5OpfZtz+83+EjgpF80pTitCTs/dierzc3pqIui2
XAAoyE/Z/p802KcCEpGf96w6x0v9Bc1rVo15LbZVuP5HLiujpkFwqWc+gario6qY
B8ve661sDyZGV+PxbUoU5fSupKxr1CqouQzzxRyMe0CKe4ZFHQCPvcePiRhcTAXs
O2coT84cWpQ/er812WTsXniSwWb+N3YLrCX9g2QtJSAGhSuEYVqtmnmmUOYrYJXE
pdXsm+qmCD9toTbNcuqEP5ohUzk7V/vSbus0XhUuu4M8F17qaaXOUiaVoYJeTnZR
vFIAkcGwd4LbWS74dI3rQ6oJl/uHn5xkL/ln1FJQRrki9CRIXP7OHYmmCxETNzVk
hvZdAhjnM14de7K8jzmvqyeVYMCU26r4O7UgUBVUfskIyYne0VwIvVCS4qTCgzO5
TxIoOfIDH84gM5j6PEehr70XnwD1YOqFPu/7YTWJSsZGVu+wbdcLL3XzShQEwBjQ
8URP8oOGgfHE8ztfNjhxJhlAeABdYxNZgoJlgUZU76WpMEG9ge8zQzm4UyYESb6Z
SdJdVdcL98QvyAs5hc0ZiMGTwTYALGT4P1dQMPSrQ4IEE6WSDq5PUFQUILSndc+R
imdWa6XtHUjrBs+ESXK1/3vd2Y1ZXfKAED5bLMReiIZLkr3jV5frpEswE3+k/suC
7OuykFewG52EbbhqhcsnamXapkIXbs66Wt36L7P6OQiueDQDTBGd4m4G6H1nbvMF
d+bHxwCbfn12T7diEa3YHuh6Njq1w2nOKU/xWPRDw9/IBuCLSpmpG5Kj3YZIbe0F
vurNBJPpIJj+IHCYNlHkWJIQdfrV54H06B9QWFwoebw/Ns4qXB7FewLYt0hECxjl
0tezCZRVZBOXgOPcti+FR66G6YBESGTe3RGZoYhZh2a2nZBGm8A+9Eg+lDAXtFc6
/9dfKvYvbkAa43MqBRnVqnmnp8Mcf9rKpEMq+i+HFkjYkZcAmajUNz07sUVShsQp
Qmpd3nAl8ZJG3qJefWFQxyUIi8I2fhYqek9os7RHN/EFJXAGGQ4n9nhRmcXacSha
WN24fTkm7AJlIZE0d18vOMN4l9wIScnOmuKRJClZ+KUUc5+MxPwFuLgOxVrXgzfp
RPoNnTqTy90ToYESjcXkt5UNx8JlSrXrI8HXvTFF/L33ZVlE3aPBI/ZFg0qHG1De
y7jAUgv4RR65JA9ACD2u1k8H8kwamGpa4S8Q1PA0RH/ljza2btPmMtxATdqcxFTC
QO94O4NffU/f8mBVZOYGP2juIhyR/3ND2gswikSKQDcH+zD17sTR8iY82ecMW6Vr
BK7s8LIzTQn/d8Xl5Ai+EdWu2oHPv095B1pqdTEhODCL0dzlwOlmHWcn35wCNutN
5XcPHHqSiTOudrA1EsusukNM1jOvGv9cS0XiZoGJ1hJAIVyeqyoD/F+De90WygT9
/MqUzNcr/ZPL8IhMD60tjaeWUAGVXfBbJYcrMyXfuFswRMNfyIWN954UOsTDQM+w
5dfHbB5ddiqluWXL2yrt0Fpo/SapIWDPQ7txT52eVLDLnYGJtSnWSpG0RAdKhRKf
mZPPBNG+X6OO8fwO/FvYAf2DFhrRDCMndWDmUr/+B8Z9S2mKuK/Dk9E/h0K1JmTn
qfvTRgsZZ33Xxt5JPGof/umpuUKTs+SJbaaXSBKECz2agHmhZXiudhMrz0KfwBYq
fZodIYYxc+rDOqCBc2I+rS3+4HUuzwbtX3219Ds4h6bVALCWmAHSJnw1z69nHjK+
yIYB7m2HgNIqegr68T4Mq32hFHclUN1TQttuCEO5ZOq2t86sZsmq4Wfb/CUv9uct
YDCAGKWHwFO6Yg3kzJDVJQIwX3u/RIJ4K/2dsuEGrKhr/Rf6RfUnjbWIh27mpHDr
fV4DixujVNL55S2xYrn+1VOjrtc6sZwJ6ifMGRgiZ/sSzeqlsS7O/KwkexMdhjql
rtlIjlV7YfM18dP/Qhg8PdPO8jjT3W9Fniia28IIZ0Bn02p8cK7KFGNhTHC8ZQXQ
LkfrDhef86teKJtL8xGxLf/CC2JpSi5tWn9ASqfP+prrSlPEKJ0RYBdANfuYMOqL
xspCAMv3vvpn3K64RfZgsQ7++H9HH8qzb+Sbm36k/Vk4sug6dVDZ503zdznLnCNm
e8ceVcxpPFMdhN3tBeiRynPmtGUI9CT8Pb5cZ6sioSLWby5FDP1hdGVDefSfbDoW
oASr+LJysmUmD9tiOy+F2Q2R3Fhl47MjdfpgQ4qlfpzK6JVDCX79hWQVwuXrJOjb
j+w1Y7tXqZI9tqZlpNXndIH9+c8Hwf5XGtHoyMeicp4N1n7B4GRO4aGQGhuQrP8F
Mwm8P3qKVbtcrCdxZHac2gSsocsMjNetlQJaC9/IkHFWzwgloV5kvTza03MOaker
ievXjs7F+1Rnt6Wm1OOd6P21fQcVm8K17LUkkqD4uBg/3c++4ti/Ap9ZY3FoCnev
SxSxNTCaFH/YUQuuqEd/IBJrggG3R2krV/2VKvpJonZpW29D6Ys42P+uLiFcLDJC
pP2vNLOl0fmyoGKn8kjHu9qlZ2O5ApaYoxsgI5YNxg7wlIVYnAKEfUo7+cuuNdPd
O4wFRsRGVYaHcZh3FNkCT53oHfYRjPp/J/lVdv9rpjp3GeMQfpfl0ck+LWSocz34
xnpP02ZM3eqJeqo7xUEwLVLFg+vJnl/v8vXDdG2t5wbhQnCAUZqwblXQdDjdNcra
UKZUxEwBnBrQiCDkhmiD6Ux7+kCebvj4+ZiYpUlz/TtvMQeS4r0Ya992zyNjYZhF
voEeZ2VCuxsCLpGgm1wqgx1K3wbeIYgz9pd+wIIK/Af4dSX7XbBMM0tOITezwJia
SBv8rLMiHuiaB1zJqX+CF2DmH8O9TdntB3+BGjmHpnggQkBdQFCxB8xa58ulW88H
CPrLMNKtRHuCdJwDD4Hf7AXTastvDA589XRSTrt72B8lQLY8y3TMpNpMC4tB1+xL
XrWmydlk9q9O1cqDdzOclpqh2uOu/IyguKWhZ2JS2mE7c9w9O6VKqGBZ4O9JLW7A
Hq27UL1HcwBTM6wQFI42FGORi43AHHyJIFJxvglaGEzBcCLoRm9bT/3cJBTFdt5I
z15MtU09QZgkaSwBI1mph0ZF9hGw94wshwv2y+x154k8pRpYU01zXKkZwWtfjCJI
wNmXA3+LtyFOg855YoOsH98b+0r3PzRdy6kx1Yy8N16xp2NHU9sH5iyKIkasKKHc
jm1L6HxIkVd4YMb/NE6LYNkrisX2UOHbjIudbCLjqDdL0LIKmRytwln6yNDGxtSx
nf/U8nDdT198b8R8rclv50pxziGEAt9pDucnf2yVsxxL59kuhM1q1IRUxQ8kP6Ja
9WQoBFzypMrjUmbxqB6h1WvT3BzJDZOuY0hMN1CeiTol7cw6d4bm3LfV7vOIZ7Yt
hj1SFJ293+wYhz3m16555TLH996Tzokbu1bJn40SueWjgmnw8slZQJQNDgm/4BGw
1YwWsWUIQHR2YB4LMXxgc/JYfqVBfBXa1ePHrdzdFCt6lpHtswS8TVdxAukED6jH
YGHV+E0uz9cTCs+S6EzD6thPK7mDiNTqyFniKkwtww6t9j4AdPpnETLLjXP/F2B/
nP0VUxxi0qVI9yH/5Ch58/2actjVhuNjuudN/xHtfCF4q2DRXFfwfTpI3b1ikXKS
y98CUwfQK5S9P4r/Yrt2SCpTpsiUtBtg2xHVytStC85OTQvfDaqz1nFwQJ5nlqK/
JB+8Ue+/DqWxkEXjrSgoqxk0+T1nfOGbGSJ8AuUXPb71Bkd1qSSUjAEgGW4CZElm
thC3Xp4PDCFVGOQAPl+TJNfX5LieIyEJHJxKPp1elnLGrU8jeNEyEYX0KP20xqWR
xT4xYYQPGgzjlk8h0USmJ5F+25f/icXrRJVsPrgk+Gh3gd6jn7lLI8NNodEcGdvq
GrN3Zl24tqcVziPgIx/hglJW2icjArdAUFFLpLti4OhE9nCzaLPesTXy/CiZoHfs
xKlVnSoZRmbaMiMoQ9MTIsaIHChyRU5gwl9PpP/+Nh+rmSVU604KVVvSl1n7EqVE
p2giOY25P66VKykpy+LvtkWNrM9ZjHH9PHJjJmIa6oCo9I9BhriUopQMV4oQG+By
Dm/meQBHxlowE8bSxqfTHw4mP0NbekQISXY2nAfuzETjyuNCw51YN9XVTVRfdLzi
KgHVugvW3wj+JfQs52gd+kLv16WQ+OCgLvfwzbBZdEqRSJ12QCnrMQkRbQhNzIbw
wOhvuLJaBL3z7rnzdQGPiaY6pOLbXPScGwZ6jLw6gxIknuyOHW6HsIiyJvAClDSs
JMZoEAr7jcW99ie6Dr+bzfuxng01bCNtX9Nk1cBfTyg+Qey54SmdQgSH+Bj96TmE
voB/04rU0dhIeWILcCfg+vxOPcZeDaIObuzU+KmXXfMWi6cd9qMpoFai65Ss8edX
1nDxrV3R0VfPIq1CwAXyp1q7pdLKefm0cJqZC4pb2cHpD60bm9IeaWAE2R0+kmV6
5hChnqse5aCXPKO3uR+Nxb1YSkPcdfW5+sv7b41kksDyA1lfmhjjnXzQIZElGfwB
NsMkLrUrOCFB0lKpBsibTFIewHRQ6phOq18cwirtoLNbXNRm1llkYPBEYlZNk+eU
tg76hvl2Svboviem20VcXFFxk/jAZmH6cycCeGkhP/OmS3SJszKO6MoEkc2GPK2H
uX0s15ig4F29zD2+sHI7Szem6HpHkpkfRFY5LiLzUFSIfWzvDu3kB2oJo8f3XQ8W
oLxHh/ktoAGIJtYN32LcVWVWdHSrJI2kEDAp2BcqWBA/6ejcp6OkV2in18T+y7w8
luDifhrRnGVhLraFEBZa+mj22TsUDW+rN1bTQohHmxW9CKJgOZaSg7dTPESf6ycm
fA2kUf2RiUpFQqyadZg9kLvr5+iP8Eh+nkRYd1pCfhUtZWrYl0dVdkEzl7NkplOo
SmSZiEXVwefzA0mzjzs8jOIV905cnDYIKpc1PQ5gHcMVK0CcRzHZOdmymbZuw5d2
AB7n4SdKAy41Zy56oaTXZcZmehQf0/gcsfw7bEttkY68UZ1Q6ms1QeTRPH1fZKP2
OFw011m2aLPik10u6udsZD4j9J0/G0eW/pKSZBO2uVpQ0feGOmS4gbIar7/99jZ0
FGBlLa+gguf7DABQib0wJoOvKRlq7evQ+j840wAYuU/zTdOLCD2V1L44OIGbR0t4
btPEjlNI09fUc+HNeHA4zpjylktjGoR6WmYpz5cZGk+5t0/U/D1XOp8Y06jmwfby
khZAUpAZC1vK6yzv05rmetbTUII8doqcWipapU2YEnuP4FxHuGji6vczrvjf2Nsl
/bWiWPjx/d5RfdAcuQmoi2kTWliDZ1oIZmFZBsNJNGUvS0dZOboGUJlijZAm2oZY
KV7Lc1AT3hzpDpisLkMll1P7Q961Rn+Gi21sYlj7lYnwJxB1KCH//LS+A4vrikDK
WF24U9GjndcOIsthFPGAciKQuQJMdUc3AcxsbFh6JOCTLuKxycKOdtfR2ckbNqTc
zAUo5pHLFlsNWpx7DaNBy34exPViHkiB8W3QUudkzQRuTYf6FUGnowX9vn0OI3IM
5f4I0sWOY3s80aU3jiyLqTOf4L3faiGI07ZricxunofJNMYZIfNvbMOd1ni5aU6i
gf2qU0W5aWqILN264Lh6vEPNicoQRKNCOdoDItBtrxBaL+z5H+KDRIPAhmZfTpES
ttmaF4CiY9JN3OXPw6AQBwUNrZ8wvpF4oss6uBJvjvZeHqNNiu3GS97kHq44IDiD
uNPe+8UN/fSm1bCoNIVjyNrvTbi6eZojW2mQE5vZ1/J+yk4nhXt/83Jv1aUrLv3l
xmg/JSW/yBCK2zd4jb6ySbuUYJkkXIcXxGaVc2DYuiKwFJJhThYpcL2arLtbZFQL
ks/29HUPuCG8q8++4IIXasspjP+v5YPBM0Vri27+w16e9SX6piSWtHl93aFMJ+TM
mVVw3K1ou9EX3edGGCm6tdE+/Zb+ied6mVqYDTSi8Dywk9g2653PyNM3gZH0SlA8
xfwT0Pd90COJTfaNJhB7p03b7iL8AEH3r+VAJlncGuKaQVvjOQGig3BAFlryJ8BO
keZG4BKOe0K/ZXgcPvqXyHJdHy3nlS+qIznzSpzgdky4MtN3UrzttIghpCV40Amb
bb/qktmLpU8x+vxYNwl/HKartGe6mYipUyuFkd5AwsosBverKdL4ueYEhMvvJO0t
kSodQN3jtgSA+GwAhQunHgWHuj0NIGk/BU8eXfpmDBnCrFS19GB5d0p68XH1oMeY
N13qqpZAar7EMsLLewpzkAjRwMJ2nbeEpXGbvdiZ4Qs4Mvx4RRrSU1BBe3Q4rxN6
kwR3f5pXGe3VpH40A1q1S2J9BGpYVPVdBMnZL3zneExYeP434AR8Q2QUMuTm0Z25
pRhFpg1O9/zRxHjaFFeHdZhZlnRlmyHHNakCnn1dh67Ia2WA0722iChu6i4iCdF0
5Uv3Z0dnDkvesNEk/SlfkHkMIDBkAALfI2oZu8W/a1aHRL51FJxTLG7DhMBf2JcZ
+872/vUEK3ec6LjiYlIWgNjjWMRqHQpl/wc3nUxSYt1DwQDmrw7L49tteTGopTnz
j4WPPcs9rfKuarJu6NYWgqDnGeSBUNdzhTOhjQLHTuTocQl86CuNswwnDEpKI88y
58oZcNin0/OsHhJEzvEO/zD+Y4tz/tRaVH4ZVV2pgpdDfDAhqOLaNKtcDFnjeZmr
ycX85EBjTkjiEyZs6iDR5S0bz8G8dJxKUgcwxdk5T+PErGS+uWmZdgurNHsDyl4J
EYiEfwc+Q7/yPMm2ba1sj5/HNaVmcpCFyLQ81ZlNNGv5cPYoJIGMH309e4c2gyEr
3tit17PdS4wUaBlCA3zMDL/OVKDyJ4z5k5Ymol7BWLveOT3z8234D6ObWRtXrbfc
u3dZSsaQuO7Kw9H6aBtVWu7EvkTeJb/lHtAkipN4Onz1nuHcVHk2NkOWBJF4WADB
bbMdlbK0Kp6TuegejoNOw/3u+cWxEuCK1FA92d9tNZxdp1kzGATFjiNktYPoscIs
8mufQEarHeQ8sh1GAtazrviZaIkQSePbBg2Lp4YvGWY=
`protect END_PROTECTED
