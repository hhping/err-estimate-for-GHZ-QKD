`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fQWUYsmoAzznR1mcnjXa7YCtJeV3E7X7dPmkpDk/z2oDASR+ttVgJ1aGH2zt+84w
KbdE5ub0tDE1tJsEKeZZOAhDSPegwT8xmTM/k6w54rSefvCvEyGek3B7bqLBidgt
1TiuZ/CowjvsZ9HdFAvRfMd07EEIF7NOuXQ3DOE8ED3eqr3hHhLvYbGY6yI/xtcy
sBtOr47bR2XmXxub0xtI7W1wsEMvvSAjtKp4qicNLwqq3sbyLGh576ubUKsTP3l+
ljdwc3axKSvms8VoYEcfiJGMp+ll8N9KfGGPISASf9gIRCeZf8QXz7/rWcCEChWT
Q0m2ROwW0Bs7dyESdagNt3W2VJZaXC7rgujlrpsW0J2SUmlu3mXEjh9lrTasR5sh
MzUbvkbFypuJiR16GNXW1hhhF/qqtqPea9O4P7T59ozvrC4IPztHgx/IHZHA6Y4y
`protect END_PROTECTED
