`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hD4wGm8RQS3RCA2E1HZuEv7RpVwvOQWN/3U33pcMwXQRHzDrtjDxYgB1vT04Bufz
mPIIb3AaJXKEn6A9P/KEEneSc8UWp5I5Pa1BV792VwI8nuFAkNzZHUKZlBqJkDGs
BUsPiY7pwLdoxV8qjqUDsFXQqXf2fQo+gJEfYcxLGf/SORyCdunVlYlwDX+YdOS1
WCgcXG7EpNuleq7xBE/LRTG7GMYz/2MaO2PJjdYDU4ZEHnFQzgJdBkKeaHt6NxB4
xCiaSdVEfxN5y/fBaejCul2f5GcsXS7GjHR7euKURVWeZRJQYyWCRvmJDCEXEtyG
Y1zBEdDgzQwuHW8lx/vWQrvuJLzkVtu5zpH0P3fTBJ3Fh40LQsAo17/Sm30fbvis
AdICoNdpgtK1rSYS8qDXP/y2AsHskzoP68k8lwjKvdFouNn169+2EMXBEHjgBlMo
BVEMpz0c+sGxdvRufEMZwYJ4cuynF9k4/fGe2U7/DAYvwm3AUr+XCzJNcCnRQSnn
THPT/gRaCeCowCPjVm/1ifqg5s1M2eVFG3gy7e4HP/BS+YVXd9A6UCUDnPtaqn4I
Cu9VeivElVBGRP3AANrEgEwUHQoPmdIAurxDlGGuFbQm/st14dfNpjkxGM+yUqzN
a7urkAF6dDzH5cK5m18ulfdB5A3dRZSOjv8NjCLYdGXRZxv9k57xWZkvnaP0motT
hKHmz3TtuR+hZrllsDZUF88LB8LXAHC5LhMOQE+Px/OziW/GJIVRBD180Dz3LKoT
+Vyp8j//LR5BweoSIpUoiwOGJ52bMVu3m2ad9ifnPTRyuKSFyjBINgi+KZUw7GCN
bx5q5Cc7g74bItWO41dJgybgmxKbCWeqgYsIZPb/pXL8L95o2546aVdbGsfmL09Y
rIiUuaSgZYkOyvzo/dgX9qlqPEJ67SUCq2z3ktSM5YYXVjIFb4ekNaMuFD6rczz7
lWeyHAmTpb+rgFoxWPrIa+ERAb+Wf1dYLSbjCWIjOCwma9zTUqI2RdrQsmdyPdPh
Uk5z6Zf8wzaGzX6BW4zB9jBb5mT7a+su2PjXLuufrcbS78+mHlLgOH9tsnH8oFTm
nqOGvUOvrOLed+U2LHEwHJSFz2ahPgzG+ptnxNyp2fPEh8ti3aFanetYha6AIo1W
/UGfGbwfNCD0Aj8H3V5u4DtYqFi8JLHXBMwFT7TrEnGQcuRjVr5pJNrU1AOiyp78
q8HO0LYgy2KuVmk5EcGNyXO7mmmgrgq0eomImBUqf43s+3gVBZjeeEoGsX8YOVTu
cxJp91CNPBqwwpgdSsqeuLN4RYMJSYWq4FLEQ0BHnG9wV51UNJU8mAduWwtzABhK
MsLOnIapwfXB4ksbSOvxBzyTDGCUw5kvAy3dpHWRYOui33Jw9KsLCffJC34jGT9g
jT807zW2MQkjsAMWVEgVF2XLvX+kXJCrQLch5N2t9x7KpXt9i2RgXC385t9jczhB
RNTat4ky++JFMqvSAm4dmV/4iouERJhy01s4W2UeYrwWa1QAV9suHSkiRDYdCjPP
52/8wzlZzy73Ugyb+ftGkwi+G3UJtA+lQyJXJJWosX3Iw3lWTwl5NXyHSsNhjDuM
Hf/o+vSU5ZyowWYBivDP8n/PNhwQ0qkfHNblthfTOBs1DRgwnQ/W4hcuXiL/Z7JI
rswYU7dRxZ5WzcBSUH5PYbbDdVcRtQQnMsIFLyuHV3ladp+e6U5EI7nywh605kRD
S2I7aoTvodhLgKFYVk+nTDJYmUCez2AQwnI40a0d2VhKpsnqPufFGoRhej5fsqLm
`protect END_PROTECTED
