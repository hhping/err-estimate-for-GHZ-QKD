`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LUtEZg0nE6dI9n++2BWfMUGfS+bTYIF+67aoSry1AIXnKG3hxPXw/UQ4kcIruZrG
F/Ef+5Y5ELrK6F9B+gRiUSHcIK9d6pWzpposvG2vjVdjwDs96VKZ+jI/a/tym9Zs
Q65hHEyzimGYiiODH9cf8d2Y+bAPgw7ppuqFAnkB+ubNmAiWTgshwZ9Nl7wnuY+w
5kMm6/onYxqMFMBMQl3UQR2gjMVTYEXqcLGwnwfvf3J0b1ziZORrkrPbEO75FxSI
cYJHIsE08iXXU4WowGXXlhCNcyRuaxTZoaxRggf3Ng8/4Iz85IPsZZXIkITrWdBs
kLJjjX4aQ5nK3/0fWVPF7lKDsfXPcV4CqbchPjdpk8smd2wNdGq5pldU/jM8KYzk
QVF8Kuk5ndaPPU25Vo+RTMJ3i1phuUC+BEWB48FEo6LE16dEN3Awm+29tZ9uiAKY
Uw4txj9kTFu8o4lpsufMe5DHw4b8YrhG9zP5xrP7ITxU4mJt6JMxEEUpUQabtm7Q
JkrW66CZ1g/Y5LqI9eb2+7fW0Mk8nNcg0c4LpiaHyeTp8P0zrrm6+3iIshL66tU/
icNuTbyVt/wqPZ4e9a9gAUeVTuZQV3kkZE9f6BjJ8aSeAWNHVhiQ0fj1cq5lr7u/
pNDj71LUO+o9tLQlJxPDPuQ4uOx0XgPHvIOGBfuLdfxAN29ko9rBKmeadLs+D7W/
JWovyvza/7QJLhxHTLWzLIYS2dwr4piYdq0x0uY3YY2N2cF0quptMirsShoeM38v
FAucT8IgLCierH//Ol3Rs51upOFz+cIOf3E9j3LipmIlxyALSnx/ZU620qMXBQEG
EvpaA+9vI/KB3NkqA/aCbTDlskIAbWzxCZ0HYwzBE0uXJy6zAfgIEzo5VhnH3jLb
f0cYFX5xwkz8GL/3VFRn4x5Kj9MhjRziiQxVvkrh+krhWpgHqED19iL4KFizpEjd
xzX+BnBh1b2/9cpLHr9GtLwsoESGMLU/TyTXVc1dC5Ud9iaTMEXzy+wqXLQ7/UDC
fFtqSU7YiAcmH75NDqQT2GQBRGiyR7tQVJhAgycaAP413D1jBvj/O31LyuhEzBue
b3d2j+Z8Kqmplfvi/CTuDdX7hV81GsQogWTe6IFVShVeAAjIHKbbvDmjExXz/tlG
en8YRSh318K98MVfRKLq2/BlgYV2MhZaXNVuj0tlIe7e2qbojA1I/tziw39+84H2
+7iXs5bhqs+2UgCmrm1GO7BwKCcpsWSPIyJ9e+RxR9uMOiyVjkeWSlc3ZfKSI9M2
rmQjK4ZZD9TxT7lDf0YTsEDJ2kAs8OrOhj0ZnqoJ2QLbUku7omULYKvjBuOQOYDa
ddl5yKk6VspcGwNgIE19PdyvShGXFGbOmuaMkLTAtG2+jZjU5/NG8TmB5BShRmKG
APJWMTIy+glWjNUz177YMVB/gl6sGv4uHPCe+J8LmA3sCgU1gt5m6ayGzQOAsgmo
LoPQLq/je4xuEtK+d3sDlKedpbfb6qxiXrl5kgYW8c2h2Hl605D1ab8dkydZbX2a
ay2rnzM8668j5X5onmkuZg==
`protect END_PROTECTED
