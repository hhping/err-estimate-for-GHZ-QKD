`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qsqPKztL7QA+s4kRtEQGesUoqAaDCw9QDSwrCgMG3KILhSwusJCyyu2bLls+JxOs
OlVlvZYlgTkxHdxZ4unesrhYfYbk04fdS83ubL3dHks1eh0hDuDY/PHcVGVyHVsS
5r3XLQGDF1mL5YiE6p6j1X5ZZK+Xzhm5lE/jEIMk+UQA51qPc9XzJOd6LikRRQen
3QnHmU0x0PD6pKMvcn4z7c8qdshZ9ePKP9YZdyHXSL0CGBX9z6mFGV5f6dfI9AZY
8xDhrBWQ1VsKLAG3ZeO3/XCflWsJ4YBA5i8aLWLJ742YpAYFmA5ayVI1Z7ioh8xx
ypu9+56NbVLgFCDbt0b/tbhvBnFm2hgAyIIRjEl4aaXLVA21WdA2W9Dvfz8phaZM
SAwAEIuZdZqyj4OVYrTPKxS30pX09OJw2qgYvhosU38KZasCmyVcZ2LWqoALJGGG
cAbuAQjTAhvf1kl23mDfgfVAYQhivMs9v/q9j7Je/PHQq6PUZJ0/tYtzRqKRy15r
ZTHOtQta8UIJwWDFW7bpyDjF7vTqyc8YhZBg67hzQyWc6FnM+6+hSQ5UfBnhdO/h
WPm5qE/b5J8g5hlD4A1WSmDkln/LhuabT3RxEEBI3rptpeaNNARa/qgLtUryXOhN
67oM+yKb6rS97r03XJYCPNJUXiDFGgM26g9UNEHIJjE/wkXdu4P7GHSu7A5gl5/i
f0fDa/ZRHZYB8S3ZWlb94w0sHr5NsWcHcsoLGYwJgBh2mMtX23bEiHGp/OVlYUYg
lxwCmkS4m7Chr+LkbiDnbzoRE9d2GTTp0cB6DfELRmytu4OJ3MDSnDKaKWw2IbAx
WmOH3tmz0DVLAAmE+PNQ1Fl8nmm4WWA0L+V/+zNqyY18cmSZ9ASp9+PJ7eAjuM75
8u84pL3OaRLkKtyr0d0DNsjH0zNM6eNO4Vbqmh2j9elfp1Yj871qEKctIwG5ef3o
7GIHjp7onp3ecjpeg5zrvvYRylTxoQT6o121zalSJlfcsi/x8qwEhG6Bhn9c2lRV
5sMycExbB8AlTcE75iA7rmOE0y9Gg/QxDpXb9X4/B/GGT6ljU8CIb8OASv4yBnNn
/O955HLdKNEo6QzA3un07jPLIscI0BhM93F848fL/ZTuEiCynHBPKOsHVSnPWWai
bplSuwcM8Q0X25/f2w/+uy5zIVpuOzZMICErK0GYXk06pt0YZWmSot9JdjvQ9mLz
gaIW9+aIdGKcpZpydQ60Xosknxxo8wcswzJbAr6DTKE/jDpbKKyV1Vmn/o+shYKN
ET1v08zMj1AXxf76Ma4fxCRpRr0q4YEXEpS+8GHO0LhNM9UyJAoe7TJKmZvwVrpG
hkPbp+wl542bnPQg6KPMyzin3jeGK7efZmresTHQgmRDLb13GuIW0vmZHMkPm6Eh
kNqXhEK1TDKNfGZrnosD4zXL6hiPb7fHmjaLoX0R+CNYVvh12LbdRMS7eZp9pEpJ
r+PKq5bmhJsU7/RkpHZIVzXA0EE6dHJTFPPOtuIoSe2K4XN2kic7V6hhzXerW61R
UVNZ6PflnBbzdophvpLrxfhCfYQBr7Si2XikDCx05yl1kQaYsfZy873RYMA1f3mV
dgkvE2FE/MqZT514KsZ8Bxz7kSR3V8BAEIV9olxTtzOIFq5j1md/Tp2/18WV6YYm
yAyRSRhM9k+Rmiu2D56LPRQ0ycawOndCRZAxpQ/7qw4PYc2bDY2dCq4RABSqnB4K
kI6fd9DH5YyrWtrtOt3ZAQ4zhCyV0wdCOc8SE3HXz5SA5WB21ZdST+Z+toCzlruU
Rq7J6g5NJNVllRIH0qT3kfjRqInWbMikg0Q4IxyxTvtMGI0by/h9Lroc49jelkOn
Gtg21buMA/P5wiocjPnbp8+t0WFsPTbvcqgIsHwJvivkFEiMtBisLS/CLJWZIUTn
45CsVHU/gL85hgrK9+2Tbu1vp6rPfyUsn2tYH3J0fYg0L2z90C3BY1G+ofl3P6Qq
`protect END_PROTECTED
