`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jMPVSwN9/5+GURLUxyshLuRzkPR+rxYLUQN5wzfdKWEXbTAWqiRU8NXW8qEdXR6d
zo4EqPiVdSAtSUN6yJ5m9ahZr09/Xdtvrq0vqCehLX/1DFSCnd54+AL04DQDHqge
ce4pfkkdNcbHfUBvGRyAlC6mP9r/bS1gxhhKdPRT9FaIoUv/03zkqa+89ifFe1Ru
uuAVtJ7Vjupi2E57Ar9Sc3P8/K5DVbKdYhwY0C8EqTDJXQJ3KCVRDikhk++pGW3T
a+anov1qzH5S8cHT6dKjuWu+LRmdNEqwDRTqHx6r9wFJ+QqPKt5lbzRohmHiri4a
FoD9Akty89Q0bF0W2OTDu9z75P5IQG06d7gtA7k+oh9IRiaaW1CzFupv0LQN1674
w6ipuktoIDScQctyhphrEsMIrjNJcgLv+4QzsYZNI/G+uBu0ZN3BWqRkXMgVjDdO
ff8ku7TSbKfY4Nb/5RHmtYNd55W0hqgBOIuEzCdv3AIUXAr8EWc7cob5axhKoTSl
emeXZpxE0Evc1YsDd7GGyhV6tS/S64TBrQ3a4LkDi6tcKM2bsJeNs5ZWcyU+JX30
wH3pNXFhyMugEVsTi/tAGg/qWMY0CnRZNoP4Bl+i79MPf21a50lR0q4VOo2F9TqQ
/bMdJdcfXrOcPCzO+BHEmeqNzul4baNDQLVq+N2apuXgxIyGj8yZet2Y10mkb0U8
IEJec6FCGcF1WSA6K/nrtKVbctJzp+iDjjrEmHPIIcHYg1giIBWtzpLuiYCcCW9v
BfEs4AFsqj1AioccZwAAZCwRoSYHol4zwGX+MqkpPvO5+hlek434FxRv5+9fEcK1
kgJyWBwe0GU4l1EYhs0hDhz9+yuj8Slt5UtM43zHc3ccidVVyZ+FnBYxE1CMozpZ
hJi8FW1ac8vrdl2al5ZGy1BGHmxT6fPlAxrh3W3A/HYJlPrE9XB5o/V5A4ZxpDdq
BJbbafX5a5tFRO/QxDHYvglkFJrpYPNEyF/KdppYhxXR7dGfhUUCPJz4aCaqepxU
N2KQbhXN/gW0qQ10Tb1VkY4nb0WYswZ3+dqV9pmGKW3pAD6covAAoL+3qL7tWzqv
2PICLW1fI60fhdnwN10cc8ZLzmlR5fEaEHxUJI6+gh0zGmhR+jc+ZPRN/tQaTJnW
uf8hi3Ln7e7AcoLnAP3Q/WqoYztjqYsfMwN9PApJ+81MrwVFpW2qHEdiODDN0UHn
zeiMHzrIsf40yVnD10Eqpu+Hwu4WsJVAWhhSO/6dhJwFQNdstGh7qKrjun2AhzLm
CWEEBto7hnH81tbA8GAodVoe1R79pW8FpD2GdfmIkhY2cyeTqWMTtvdhBnpFukLa
mJ+0GgX+vZpqeRfRPBlgc1lmxR9O5eCVkIV2XPEFxdRtAlM8aGnL4J+lfaLssckg
VXwSFhhjZuXMuFD5qglHQxBPMRQFMkDFPLpS8J9liwDa6gztpph9lJjOX/Gx1gVO
tilsBZdRkj0B0aNypThHLIKNUK/22pUsvFLM0lMTSb3v9252Jz4EaT9vJ8JDAgH8
ci6DIq8C7+O++qD8rZ75rckRZWO1+7WCKiIR6QEbs0IHqqxoI22Ro1gBkx0Upmhq
aCC4TaN7rJp0NvsX9FiK2rfzsJqxRzW8JrhB+6XN887h6HGFickamfPXOKDeg3bZ
EDmild9keATz5klHNDtQxN96mnqXkw7hIC6dgUgTvmEhQp8uvLPNh7g4s5M+Nawz
XiAdhYlKPnFcIOcvxA+vBwMotqpM1U/x9vPaHKEKYpTWJPtkGc8ewrmq0leCj1t2
xOt8OagKcYlS9wFdv5ZVtBl6I+MoGMfYcLqYLc+m/ufy+XhsO42G9Pn4KVBfz7IJ
biDhgQLPfDWfQ9t8WVm9NFSMzels5B9pfTwLtP7Hjr1KxRxlbLIObDf60mpXFdV9
AYdHGzZOqLbuGit+qr9ZhtN1TJO8mDcEP4FnUADGH4EaEjxfAY3havx/9CnjaSs6
Ii0+rulQhCoaxyJsVwUiAluvGluRSLvPB+6aSIT/axFCmoK83cOHJFQqnkefR8CA
5cd33PnAws04/rQfACdPYSTjEAf/ErqYqPh9FhtcB8kJ8wu6PzLcYjPB1/1eUN95
p0j14C+dkexV8tY2heoyGQoGysuKZd1N0/a2swUa68fihJdws5QzW4FYM9qNXZP8
DH6rQOFkKxIaLp8n9cxWB1oKB8AlTi6ewvR4gBwcuuCBUIoDgqhnqkTzJkyo6R+L
yjL5jZBVoB61WgzElqUZFWyV3C70fui64ZUYNMT+lPoQdEMMgbRDMl89wWlclhMz
M+O+lU8RVUMUF/1CW+k9pD5EgtSNjU1mnJVTwq/QRGoLJYiTB1SjugA13lxucuRo
Z+gkVGTT7qGHNDVqVBrMpRbyOimwg6tYzN539k+kkptbcv1Uph0cGnNVerY2qa6t
DmmNewWAJDjFHhjUX1Src/zuFVu5Ne2ZBShnW+pWnaHTWMrO2J13Vznz2xSeH/iw
Vg2J0JQH4qUoyOr7NcY+5Agb5ymxdboobc9H2qzq3iQPW9n8TMIOWu0W6c8mPFcP
HWJ/TayGvAGViIWqVWNSGnHNZT54AxoiGc4Sq1302EV+w6eAUQTkLL4X8MZ3M3T+
bGAyO0P5TBl4D1/pW534nFytGHfhd/HVbgwwU0vRHkUnzbp5+VzD4xu0BTk24v15
MWnlVKIa8Glf8xlUE4PnZh0gkgmbozurJi5+c4EinojpJoektjSB/ilUdps4iw/U
bflsCFVP4lDPQAqaBazEn9K78JPvSQu+QW6zIVIlFvYz5+uEDrHxxc0lwHlrW735
ejkACNtr8cTYw3WIP+eLIgo6q2BF2dhVl8jFanVbgXS0x5a0OXsieb3EGf+GOnGm
5cpg9cjC2HsdF3A1ikHNU/3bV3DhlolskaMXqQ28getDYifhZ/saPE7JStBls//t
Dq1MPWWXOE3D8uhA47Mmryp5NdPox5zP86NTd4N8PM5Nz7kwNcWaDW0iJhDbLdR/
pm+/Xw53UWbDZu7E5lMXvJhb0oRHap7WYiP+AjtsOuwa66I0ulknZNJIhS16x41u
PUAcLL75I67U1K1wld4hhUzHGTnF8OpDjSM5L1cpXZz/HPUxDQNPbMHCJxRQmwQD
NMT/9ysNQsH18W9HTd5urWYchuGYUyOAJDPp9WnGMAdNlve88cET6mEhvTdSLEsp
3mUNhEgamd8XDU80fGA85OK1VwSCFOFwNU7UUCD/eVw6yD0ijDI+ojwNtFTnW5Lr
aqOUGLB+mohRfxX4coZiNDVJV5xjpyS1BmhmCucH47xAcZgkhkzdeN2GT0BMzAEQ
un05sR1p8b8vEmkBeY76ebH3OxHq3QLePJd9r0sc17TKp+OTtju6qcT9p1eDE73k
eYm5NglshEaG2xvvmHyUlr3RtjYoG4QVUu1UqV9RejtaEOCSQOvawVGWJ/V6YNfB
VNoDtA7hkJyE4792EDwtWdkV/77kFt68JhAwAamGn7K5JUck17xK5jllsUtvI4g6
iHM6CanUOklLDWr2sSk4tyuYkOs7UTBJIlX4KQ5M/CHd6GdDCm/UZxy7CaS7aOz2
nk/G1XXqbnUxeOS5oLHV+YUU3vecstSmHjnexcec+M56iUN2kpyT4pgrQbUjCxuB
Fh9qipEpImXSVQ4AZ/rCpD2PlLWjOv56oGtr30QL8KYXmwLJriWy0iklZuHFm3Bb
TWlWv2jIIoQqxwF0CQdEWN+GycfKlzf4Nq4PktlGyTEMEG/9RER/zz06qbSMIp4U
n+4e/xsIcjGox+ybJOSKQMnvQA8qe0AkXKQK+6zdF769yMl9qZMg5WbuvieYVl/L
GP/AkkJpQBrqsLQRGqvArPJDSY2+ci695xkoOPksm8fL7N7aEDidJhHk8h8p7odq
ZuURReRnbGnf8hCz+3m4SQ==
`protect END_PROTECTED
