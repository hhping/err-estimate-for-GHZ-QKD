`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mCeewUorYdQoFCRn0cFPM9QbtHORNuYp6PF7nPEWCgcbfUzKcfunBB0QCXoM8rzG
c3KMhGaFp7I+fQfzrmgVpt+cCHz1j4VdRxxO1lAU4LQf8ZHEmMKXba0l83Qg4NrL
U+LqWJ9tgCRLlNDMLYCKTh9irHNFcFpfk9LxyhpFAeuyrhVCfDkGasEuyES/MBeZ
nTTq5jvngHBEzw+etoUOfBvJ3gGQHJ+vpJ08NZAE1AY3iQRFNqf6PjxZhHUpfp8C
iq56UCWOG34G8j/JGD4/PRsY7DDcXfSaRU47NaQfRkka6pTstU+RPUJdhO+eo6Nb
v/ZXD+LJ4Ga9V4M2GlvZf4RrzLgqcDCplU+HD+h1vuWYXFp0r69q0i7R0Wy77HJS
+m7oYagqsxfGFQHJZHaJ+qq2wNQgsiXQ2j/mMxhTWVhvPOJosBlHd3OLgLhXqY3j
KvcgF/o+etSZz0GueyaUGBOXgkYEKIjpPyVefGnShWcuiuXzA7R5sFIU2UHve/E0
sU1zroePJBb5jfoxrvRGmHQmANSttysaLR/xAe+ZJ3lCSfj+XJNipOd+ZhKMuK1F
0XvQDR1NCdBHMDUoLKmveoBk8PPn9GpmLo7SvUvyrHWb5ZGl86szvq275oLFChHS
Bk6l/KxHAYNXVruYp+nJYWs0xcCkgc9Xk0iEN8LEa04fbQh1fUQ/sZJANrDS38mO
90yJM3oO9TObQ6VGTZazq3bvNerbxfjrZg2sWdyA0MbU1YWJ8FTlYljvtn9vG1XN
9bNnPFmOKqFuPuN51k8eO8ZEOM8g1XrEYW4RWVmZxg+tNioEzFkgRrgUYjebLV84
8WLOIjg0zbnTAkmAqT9U+IEE+53aH0YsjoSPZV27LP8jxCA2SxOUpcbkVThgfzEt
XZ9WDrhXHCGi4/PvHtZdJtS41GTaeRyhCsZ+6PflnVSgNQU9zeYpzRisq/5417Rw
wj9Atv8sdQ2aPiLAedb7fdMscMDvwDS6g0TogOBB8Z5BfF7OuOJ6LvoFaibuwPVo
Uh9h++te8wnHsIIRpEIDiKvSIWksJI7K5RE6VQVDwtIftKvJspW6oUeb/lPAOw5R
we9GVQDfKeiumSOWW7rBeuux9UnbgP//MmD0z1ag8aQ8tJbLm174pKccF3r7/5uE
kFiWq27D9pmbUoHjv0wAOTOKAXKsJA52dU1p5GO6NaosiiHkK48YpuuqQ5wYUO83
whNSRd6Y1Dbw+K4HSRbgjMHA11L4Qs7lDz3oLwU5jDQeFB3GvZ+iueU5kDNzvdRe
pSPWJeUy+EjwSRkTodvJSO4fr9KnnpvmYBRIvqSuIsu7+S1YHkAaDa2vVinejwl4
JJR6MCaTceaIfqEQNm3T8PQ08XIoYvZuSskocPtWBlKkanGBuJ22yDavHwKCASJX
lOMGoyxxzfOrPPQduKEpEztjEc+D2uRUCxPbBQH3odHh6s0xbP/K0aL8epGZ/MXt
ujS6VrEPVo6fox2NMX6RBoi3zOorHIndSj+4BpUTMQeSIgKwFaNYsrqOB9tG10me
z0cVmgetRVFcBK+as7PfxzAvn6AS9E8edlL+wn1vXYUjAYzrp+q7b1mJStsQMEm1
soTWuDX6QlrRSh/ggURotIVeWDMlWwn8lyPB/R5sJmq55+YWig2ME0T/VLOcbZ+w
DX8YJ97Xd3J+UM7copUwbhpD2ZHWAyQat5/xMyEwBnLfa1kx9GXv0kxxYHhd2n8F
RA5VVqie8LcYXsRt2/Snq+OgaZBtQ9EVVJBrPo/nQwlKHWd9LyRf7lfOzR7Ykr7X
SEO3MU8vFCzQ4NXXqA6/7Z8J+F+pl3+qULanUzPCRMVl+huZsFLEPt2BllHj8O/I
DT/5EQqAYPEbZlGcUDfhX/5iNzAusa2Rq2f/txD4/4LU+i+yZpL8abMMbVrQu/k6
Q+5Wtu8Zfq2QGJu/0ocK6zNK4bbR7LY1mXhEJayTrVGtguKS9IUS6EDpEop8QYy/
YYeMT1MOlhy54JU3GS1VlKJwyhgzYkVdZ/X9ZvqXWz3ZX6PCDHHTP0crME0ANB7x
o0Ss43caavO0Ck8NCO640RITkGI7vywgNY2Jl2y+ffA37Q1WtuiiRooElEItVvFj
+b3szipM3HcTGgDNAhgXOegiJ6o/Ce5LoRHhEcp4H0O9TE5eHo9v0kTxw+JxLtLE
uFZhaomlak3sZ90rUjr5Kg2Dh4+mq+2rtLZYQAuceMDro2JkCdG6hQSU6jYkvFYB
Te/5uJMGgkpusBsu2xD7ppF1bPAsC6JI6gPfLB3jNPAlJxgnGGaejtFv1eGa0IVA
iV3p5HDb7l8JRlf1DCOvtR3Olzpc01i7NnnrqcSgvD2m8iy5JrPKEydiARD/jqbV
9MEhFUxrZLEd4GOAXDGK67so7davPwgQmBd59F/bCO04iZp1dp42ALPBm1eUdEX4
5VQV503FtrZS71kDRbO44fq8krGw4K4WQFJzl1osqQeHZ0xG05LpuSHrt9TrVrav
SJ5UIziaLZZtnXgKHf9FCyxU5RYGahwz2+tJ65az9p4=
`protect END_PROTECTED
