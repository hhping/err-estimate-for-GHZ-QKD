`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tQh+xtE1Kq4bN2p+coxy5Ra1uQyknIoBdZeUuJm12jcNI+ec4XtEP/sQrgvB0wLN
DfZLgyJSx15JIE4Yn0Zp/SDVJk09s+yx0QiBF/WiRxNi/CRNUc/fcvBCXkyFZV7l
yV8XiGHFKsaHoE9EgOC4m7RKeQoJeWXU7qW+nJD34TDHfnoSwBP5UFFI3Po0pgH9
ygjnJV4suzDmkHR42JIS5Kjae0TcACA97poRZguvsnJB6xYj97ohiQJXkoOtgiWB
lKXBMpWIId1j1e3pR6xMOZqDSgGWJSoDGzcbfDd24+ewxeV+a7SrwOOvzdHgoUvZ
X0TjUXE7BBVB4Kpn0DZ/rsi1uh2ABmyCwxpHKWWd/BiWc4ua/VABbDo6Esjdgsan
18zR1wGgDnpBcVyIpa8oEAV6P2OLhq+bQhM4QOepCIXE3yNB/goQTjdxhwP9jbor
WTVDLr3mGIGkGjnok0X2CXkq78m1wK7IzG1mAH4UMkz7BUck6FXhSVKlSQk8/fRj
SXoYlj5NSmdDl5/MBDd1UVeb/B2sjjd9fsJZZRLBaytY318Ak5oQelYnGVe8SPhX
04LQV6SYJN9kWqSb8JyxliMPfTJzGLDQetg+nE4uyPd1Z+rSRoNlWDCn8Lu4bFMo
UFMiUDuhVuKWscC+x/AGe5mo1Wvp7Q3ccuGjjcIPtdlwUiZKR2chcE+340MLSyko
LPouUlea756Dnwq+P8d4fGRNN+Ny0txJc/CmWMrI3tBnpejoTs1+UGcPb3w6RP4t
bnLJqKAvPk8HYziyQaTo7JylVR/FqDmqHIaRjcN6RQo3y/UjMBI7UmJ9fWkx1vpl
dI26p0XKUPvgcGAwdw0TdhJi8YaIJOYSccre7gfgJQe6mOarc8yT+9xTOH/ksWQW
f++mjn7txGeFaPM/HVvrShZy+vh51S74QQAaK2F8KRJ4GpRvQ2B52FvoAVIhQy2d
IUStkS/zN5ixvVzGBD06m+YwDa0DjwdAT5amJI7cEsP3Mb3QEL+I4O3Eh4TB5s7s
R+EusuhejCVK4YKW/cp0fIaB/4OFfdWaHenaaSA+QdoybB1AhLeNtUf0X2LnCnYH
QPwN01I7zTGK0hp7UL+XQQJfMqWk1ntajntvrNt3w021Aav9j8zE9Q8pxD1ZBvU+
DBkPCmbEiRu+VBq2Az2sJlxsUBh91fFbuDZE4/9wkyKu4ztso41p6cmhDLCCdnrk
+x3NeoFIMNxHjU9Jm7hYzPM7zTfke1jYzthKFLaqVivlN4M2nDIXehVavA8o0uxw
XoIZtY1Se7eK33HQcYw5q1AM1Q230/ZbTw/mSG0yWpDGIRSJei42IF3XQdu6Qgb5
1x/HqwrUBCG9+fKQEqvmBKgCRlKf+0PTykjWsqa6HCVNjwq9Uz9KIRaHf4BIPdu0
I0CtgAWTH9B2LlgrivQIHv5695WXWeHdIiW1fKarSLlxTkcIvNGllvzcfm3IZj7H
lnvmmL1YGG4373/WoshcYvv689FbKpZfLviAlDehXpB3Ca3NwzwJ1ZNwNifF/cqF
dkdT9mEuj3W+Asttmo7/Cdzrlu/oxmGunRed8MlTYUDdW0/vc3I9rECcIAKrq9sA
CHQbbeTHj/hodTqHT8sTmsfgGQszZE1/4x7zJ33GGTMWhWtayAjngT2k3Bg/QKrm
9SVI5cUI++stcNiGeez+Zan+/ha+8w/hf4kQH/VWCSzAWXhgocubSgRkL0ncVD1x
j9TmVekU5X1uc1AecT02WRb6ipa5JYFqPS8LR4WsbSpjmiDCSkQwhhA6fHe9N/5M
8fLwdI24r6MrFyx16QaW1F3F97X4F9KRFfrcn4TDivVS0eHNa/EeZevqqXFeQB1v
c47oKT6b8jl7y360Sro7300gQ3/NIQGooTfp+MigqAuBzFONgjQ+mzh8YCl2nOmK
QLEBKbrsKS7kjX01USzPYYncPYWw8WSPYMDVYVstY+Y0xI+++6+QOB5IwbT5GCzA
i/dqGUdMbf4Ir2FJh2M/Skhqwzsjw8xLOPbYECd8erwBtBXnplTfw7ZFOAVSu8EU
fsezZb5bKHvMS/pkOKVmDAsjnZfAq3fk/QBKJR4mMT7lKLHBxtQyuOLza0FQaLbt
sLY/AecZbcp+2RnBAIuCdQzkXGJNiR/ThNNpFiGxq4ToGlLJqejXG30xsCSKXdwA
oS5AU1Aksci841RnTLtIWOfkcx4Z9YJHI0GgmtJhpn8tSBZY5NKl1R395gpWprSH
H+m87mMIRk8YcaaseLSxao6pj84vTL4wL7pTj3SGhUmF4IyHYFDkKaU3l4ZwQdJe
TDYj/fmqdySzZSHd5JjnxYN649JQFPW0xHmTDMbL0elJbwY6VWHnzTgF0DLkAtr8
Jk0Mn9oBqGuTVUzP8pLNr/XCyM1z0pgwEE05vUjpENYd/YRGIV3HB9bYc6sMqpTn
RbO4xzxjzyGBM36IoLBUfU1F5sOStoTpNOtaqiafIWVbAmFnn3CNQRqQPoiuOHrg
zyVCDwKl0Iy1FU3cs2DS9R/T3p0HnsEIoTYay4SNfgeLElSx6qX4vmV3Gt2FPtlu
UBoPzk3KSafbhLdDaBSOAD2GkUGPbDcX+hciWfR7PoJzGiBC2e1PJPB1Gaaqz+Wg
kHC6M4MbqnpeQUMR323EqfeqWc3Bqj48cvMQpDvBoTDCx+03pDc59dAxIIQH9Gsw
Tl9Np+VJ2v5QyxVo3FqGv1sNk4n0uQBEhCzicQuOb1ud2rrEhXHXrI+4S/6e+Bu3
2JsSlactemphxNXqSEvUGdm+V2OLASBHCvBdAqBZmdmXmYnJx5OFjWFZU27llVNJ
UQWqHIolesAzVKcVts1W2ujA8b7NpTI2Y86nJdCWEhFMGOLvBDgNZzDK/R4bZTN+
U13SjNDZt7o8YdHAxaawodL2fev093HyGxO4r4DvhoAZEXWhhpSpWBfQf69qFtYf
0Vf3ZX0iPSY9t2LoxC4R0u7oOZlVo2e9LnhUe6qYDlPIfIIvOgk30wuXOSqlwFT/
be+5bbEjr0qWpx6OjnUtsFuHFIKf37lHjdakS31SE19jDzWfluYX7o1foalgNUk7
h0jn1QTRefW9bVzLLvnRkjNvfKHHmgCoU9Hz6vZuS02BRULM1TvsU2kzt3XQElBJ
BUOW9jDjIF7FBBIfxJ713RAlMlFSOX64KX8i5qaHnTRQkN6XBUUGvbvr81pd3M/o
iqBNuixjrdjTkRZPd1Avav//mw2R3ViuSz30+EKbPwUm93Hx235fJoVhwELm1Gvh
mFq0Vui+djksx/RCCsJYuyieAVpP+GyG/z42AoJ0NB2JxOVXTB++Gmq7wZz7DpWf
K8dQ1ytmzZ9umgZaRn1NBkWGPx+fh8yJbLQ8rxs1iKUFv7FzKatt1cVdkyTdp7iU
kibyUtCBCaSHtUbmnrTvMbbFSIp3AIpNx66sd+GvV0ynU0C6+rXl1HLevWKeZ7MB
+LQza1gQLSkZheZ0UcsuH+Bqw0nMUu8wJiFSKs4afZ/J+TJdp6Ia+TIigahRKaME
gv4Cg0KrRtm9xAPYSCNcspzL/cBCMnbXQlvLNvsn583w7+1FIo8D+JdHfAnauHvp
EWMByq/Zq2lvvpDBjNR8k3NqVw3kr8KiTUy0t9Px+2EnY0EvCDMqHjLRsUEWIuhB
a1/nOyd+LO65iBRNPTqjQfNix6sPIXYSTPaRtfqaoCs71vkFuQv9VUyYjCQKxZsd
mFGJlto4qV08ft+CMMVY/8nLSskdPZUBdpfnSLWaX7Gyv9bQpJ+1iBblccRZ8IXP
dPOSv9VgaX3nvN0UGuCMvH4oTlilSQO1W5l3Mt39Dn2FmXOplwHm7l257VNEMGqX
VCY84kQb7Sat7ZOt0M6fwkSuyG9UsrwnBphb4zrn1un0k/gATcRZ9C06Rt0VKz5g
ESh/zQrofwj4qVAyLTIEVMXY8e8IJ3WtJPvhAvFyilCxoTDwPZs4LeIZ1XAKVT7v
Q/4eTbWUsZgIJTMVMZiVu5VH2Ta8zUzZSBNlXUp2LQv+VzB5NAM06SjUgvCXt+It
BH7LXhsEmsMs9T/r8oJYc/uOBpO2G2e4VKsZFnVdh7mVzMxJZ9fBGUzuv1HfsPnb
wnBXVFoNSfNR5uasSOFYg1+wlXre9UoBRVXICwXhpLu/ACzj4VspQmcQ7Rga+QGF
itjcKqURAtndHgkMBFIWuRz809hoUFxS0pHfhK0bSbh02C+EwI1BgwRpFzT944OI
tki8ez1wS6gf0DycwqrcL/Wuc3K1D+xfKESn/EXnGo+AIbvG1F920xQdovaiFZU/
qEvI/WoSfiag+sBa/5pXwPaccjYg+8YKrG/OSPj1aj48SnunHvV9e8OCjepUK2wJ
EnDgKvU40iQaEvbAWbFdQYZSVCMLrWcGtetk8RxfWakGJmcnaUGYxrCBGN6cCjkA
TNOky9QfRz+Y3RmU/O8Pk298obAgeCIQeWt9FKUMy3k3Uhcu5OYVdlDpA1wQHu31
zmEB0T+DKCtoibP5VAxMcGu+FMssWeR7l9KI6jdrjwTirytNTFPyUZVQm/Q8YPmY
O+H7JYXlGJzpDYI1GLZ8HsuFgdPmlVsekll8mUMcUrx8xGhcjc0hvy5FaU8nCOiU
Wt3BGK7Adnx9ErK14OCAN6ItTWck6YJgOnHsyqzpQpOcu0pRAEMSt7Jw3PqGU8+m
/PnEzsXbs9KO7rVuCGnFBVrl2FL+DCH4sWEFCHxZ60GA3xqHCkcSkRVpNVM1k6oX
6LRkcYw2Kb7RZst5XYCz93xG/5XhphqxBWEIqznLXYFsC4PpneqUjN2Qn15wGMup
ED+PZh7nAbTVP3hATkat0dzyJu0x2P+965B47fK7bFZ06g38Dehg+nhMerXskE1s
4MmzdiFe1Ux6AT9UAJZ/hbZYnt1u3ySxTCJlcYlNPtoxFLgDY3WA++OKiqX//vPx
TFXqDsNFnyCE1aj5o7XenAL8sozmndyVZpsetnE1AQxz7OAJtxlKgRWZKFrK2BwW
ug4Wv8YXmdwnQgWZ7/TArFZWakW0Pd9+I5FSQgs5fpRTAQhHP3xejIYY1buKrTI9
SZ3wMEBVG6qiSq2LwvkaEPGb/gPnQEN2BYpyCw9H/fX2RvDHMFN+Qi8zSLO/SCfy
ayRbVeRe4S0ClqSTgvv2PU6BJMHiLZUjFd9Xy1X3RBrYPG7GiU/nIfPTk5k7O/MZ
RhQVxlCDIsWh8DEEcp9PBytibRG9D2GI4xQrgPPxdpCLTnLHMawLoNOoFo8e6h7h
FCFq8OfTLnrs+mRrmmNULpU+X9U1Iwf3oZ2YE7Xycuz1Z5E8e5SCAw14+RSMyC+A
dZCYdUS3JsMkxdZ4QjTxXc4iH2+WJki6v9V5eTZ0f8OceGKRVHT/O5Mqe8TFU2pX
VfIA58xZa9qgzwYG705z3GCixpoIf1mG79YBCeNC/eiVzNMd9tPhPIL8AGo6waWx
jwrJjkip9LHQk/zKDgaTue9S6PVVyTXT0J5o/5CNGP9OMAK6CCuAAV2VBOPWEi7Z
a6ukd8tC+m89/tEZ9c4podWLAh5Lwi7luI70qvybp/Q6qqe5RB2ngcOUBKSlz/Xm
CDJ7BG6lrL8KQ2caDJVKiEl6YS5azUHMUmHTa+mKm6EbEAmRQgvmTDoSo6GxFrNA
faJ/m5qpYJJ/dcRxSXi7zQxeQmxNhr8x3EvVesjvau9HV/vXRyVn55EapPYh3Bdg
PLiyJbdfPsLzPzsOrQTbd5UjAHgyCZJ75SlNcTxWYWmcJEZcZg2UpV+i2EPYvpFR
Ye8AB+QSLNwgOLsqrKyPOV+i8n9ypgAT091u5ibgzXxE+KpVx3Miti/FRVCCQ+HI
xTXzWsaLiVkd021n0S0xFv9bumgLAORy4hVpVrb2uCqkJfTYwZQFuWEhM999G7Gn
Iui7Mr8UQr2H+QFpFESEK46sobFhoSZRBEap3IwTEglZdxIr6gO0Ccx5zRjf8fvR
B1AmTP01Ytoqr0GKQr5t5br/WvU+gu5i+4gw7KXownSGzXSxtihwZ4RhY4/d07FR
Ri1Kzw4ppyW9Uo84x8oEypi4wKvoKPoMkUocg8rDwG5TP+UM/icplc32VjHkrWo7
Bb+BZINFehgftBuWE+2h9wgEKjGNNT7uxz0hfYCMvotKgT4Iq1EysgFkzHqFQxzX
PRMWtLU+VKMsN0DP1pWOQDoqGuPaeE6etOjTfpabFX0z0x/8w3wlbL0peGTbOmD3
yPA/WVsSAPeFn9zbfTilGFU+l9j/2xiJXiwdweLJQeLYkdE5sFxX2FoJxsQxByMN
MpmtXD/JhWt2TCR1S0DFaggJ1I8b+WPBGyxp3+wG67PodbxLXaBjG9V04rNtN3am
cTM3g5nnut8KNkpwU8IUEm+CondqthgnDyBPGI/P1Y0Z6knrUZzjwhQNglJvbf8P
5457hSD54pFRlCAXPhPUG7iJ1uOI2pTymQZvX+VhnlHGbAvx/w8jgRZwUuk0paBc
8bwc+41NKCUGixHc4oxwxE+KfKsxWyqTk21yXSz/ojUdi64aIEng8YGEAxfeHms3
WmlWkpmDsFiJ5pNZZNNRvPuugp2KhRqsCF/K8SwuUc52dvxElpzwIUNk4GTudyoI
A8Z0DLmZ5VZ3tVQDLx3bigh5RCFwgZ3nJpgQTe/uTQdl6H334sH1wBcaC4O81dHD
TFJv0Mr7/JD/vyJNOo+0NMR7f8CLnrGmVz9KaKcPlHmal2/xTe4EUar0y/Rq4wcB
uZEePd+uoWIu4RSup2D7RMq3eNi/uajnzOb3u/TcS7slPxgYJfIiqCfvn/vYJWZr
7z5PI5dtpptWCn3klSPsmWnmwlpS7SDuMY8jd9c1sIH9vdZ94Xop+zYdX2c6OczY
g/5U6WlhbBjZyWd/7BH/NcomTl+74/D3UbbpQhzsesEzXtePpjEBeUeGItH3rwZT
2Vj7g4oBQygaGkxbYsCkbgSqO8CbqtaS/FTupgqN3dUnOCR6yTteEZbsp0MeTnM2
6s4Th8TjDP0B9yC/gpYp7F3Jfje89Nf3grLhdU8iGt8xKOOUVfKEmM+S0IU8O/f+
q0E5aEkpt4JRXlq51yzSY3zAeDqH/bgrivO242xRWQtZ0NrlA7weXQ/Eu8T/P8mA
Rj0Jn9tbhAYj+x/94LNXarlbGaUc9tWX0WKIMs/Oe7lDlgLxJ7Z3FaeQxcbYJgzB
anmYXMF8ydMdMJ5dq0FpwnUJDmxeKSZ2zLrNSlF7ruUTi0HEmjfDX8w16nZKVt8R
AaYqQ6l80dRLqP0guFOjiD7RgmyO5ZhGmJIi6ptwRTPRE3k9Ecy6tteOMRLrNlid
bnbonFQ6rtsSeGkYH0frus13MU4TNh9Yd3XkHfFpJOkd9I2aEPCWUx4ipMKjo76o
egLpjJ5osm0Is6Oy48uqgCNRBfyst/2dnho0/c1pkcL55fCcBKkelxoIpn1EszWU
yXOZ/h1nS0xQPPSo7SebGbpZFxwvMq6a2XoXVNCc/nhELQNY/68iZZXm9wxUVeFT
DXHqMm2uT9O1vAdE6RkgbCshNmKkz+khsXAVIWbSvvmnXXWcbRswujusL+p7VaP8
FivRVaRSPGVtwDS8ur+Zg07bFqC9nCjMTaWWJnrU9tMdM/SOHVnEM5aLs1uTHkFJ
FPhRULQ1n/iCFzVaZazJEnyveTZo4SHCorCYu8Rot9wcyh8t6mBmwmdzhM7Y0eus
MZQxbKkXVafZTLv1KyrPUKBOxF6ku0hIuZ0f9xrgwjEgVYJIbWJEq+uoGhDiYvZL
osrZIiWzCoT+yW9UYV+xGRamkKfd9T+3xWEfYSJ6/Axw3rVi5/F8CBc6rcOe/dGW
g+aSs+SRFZUQlknobUM8oc+VlpN3Kmrw7QuOZ02BXPkNVBNbdAWt09xdUgEOVc9W
WkRnCTs02GwcRrcXJrd+vDPqJmk2Gk8H/r4p0y5gNomfcn5aBB77K+SiXCFaoCCr
JwO1NWXD8z2zMSNzBgOv+i7/eDzNRbzy+Yh5kFd4c9UgS1ozFc6bK01v6PvYfL+s
I3+tLmou5g+V97fhC3Qe1cxRYME+AG0g9bF2bUzsxZ/C5Y2kTVYgoUyJOBBIHoLy
GvNxWSu4fzYTzLElCMsSCxThpFCl61qz8MYIaRS9D0DfkHIPaUhkrYHdJXhkEwRo
Cam3Z0it2PjhIGul6U15uzQvikyy3efaBH4jpMOjsmxbou+okeoi/d64QQ49T6//
m5w+r+AswWmPfLBYP8mihrVAf83vGtkIHuRNwlbzPsfiU7pkM2P0gVqfTBWZxbUd
XdSmhmdDFDX+TNNkq+uxEFDsMAShkLT2RKFJhQEmnt6PFhEv5DFJ9YucaT8Lwatx
1lq0xTt4Pri7qIGm384BLq+7L3v5MKU2/FZ0iYvddZ2Kjw5F/L8Z+7FVs4/lf+DJ
5jxw68lD5vXc1k4yTF3cJxxfW+ePpiTXIx+Bvc/5k+w+371SWe0OOUGdItPxGd4D
gXVvkkiyrHGaXmmUy9gq1Fg4Lvi6kDzh+C6jv7iZilQDoWMdVvgFnZXLXsa6y77d
Cxlu+Tl9Ilr3ClUFS2DYuTHxN+DKgX81w/FQB/V/jHQ8tdLmyhhy2ExKg3Lk8XEp
N+0Do7D9478JjcaZfEv1f3dZ+W3pRwcUqAi6eeXdbqGLlYZkWCXWRzkrGviiuxgB
8wadhBQBQC1qgoRy7wMuyXHQdZSoLuwo9yVTUW6iUczdSYO8XTvqT4UBY9UVtCMS
oFfvT9TaSM5efnKnMGcBacpDzpX6ksX6rrrVQW1QU19Qwqx3XJiTWBMkNweKuPH6
fVymLHfXTCHPY3jF+isnolK2WkihMBk03F53QCbU1i6cEP/LJHxPeII9zc+XANsZ
1F6vpaGmCeeh0mGXZ5K/lJ0zVkZHWG6GJYBaSb/l2vaJlWlLwPug2r1iArGasNha
nhbEAnGydFNWQ9FuOxaHymh85PqZsSYg95ROuVaiA3EndwSprqIYici7NRfVRaAW
Sy3BeV8d2a+GAvOGSkkGJ1u5mVQ57il3UT5CU7qfXSoWCO78l/9mvlPZI1BLuyVe
Qo58fozPFD5pg8FKyGzz/3auFdNGWSM5Azafus/lazMrCjOx6RgQt5qKU8DJfFkJ
/LyhIO4qyr+9jkTUxThZ27TFIfpy49noCgsceXImYWzlNQp7DZOL2bF541v6ihW2
QBaZeurteUbYtXVyHpVIqYPJD+cT8evOSEUqhrLJthzengKnDwcVrNxXG8+bzpb7
MKe+CmlGP6/nByMA2GYj3bMp9C026l69L0nyi/urUVX9Mw0+nS8Ouv5IZ6LmP3s4
yKkxYcU/TkV3ij5mbTt0m6hE6UvTNk8tu8TAw+bEHN5Rku5CR3qI8d48ADxZhjee
SYlg5s3NtBPmBt3JX/XoU7fAZ7L9+yU1/rzOOjXlQq35i9/OZGkJzAxyvg3kIp+1
VhtlN/pF144HqYcN2NmnEidZj8c29RUd8n+VYURChb7RBj+xQAkaYYiy8rSP2RgH
qL60pVBuiyRt++pTnC24jrWxKIJ5OrG5VjdIe8CI/4II3n8+vI+6bzfJIj0fWM8V
nHeLkjSXCbgzEP8/RmqiPsXv97zhoUNpqzbhx/qGVu2s53CFLc3clI5QHVNHNPNA
9wu5XGdwkHswQ5Sn7he1tGN/68mF8MlomePUg/9fpN6wuyAo3TMjKcQS+lAWdxy+
HRVZzsDtlW5VVvuQ/WA2H2qB24RdGyBYX1XFjeM9vCtCFT2V+VQZC7jh8jzcxiEN
pnjBmNieWa2R9jloRE7GabQvBhQOzyYJIv8oIXqSAn/a03cNJ1ZS7wjDPE/YsJA4
Qi1oD8YLOTg+abYYGpdXKKP0FBAZLpGqFKe3RflaR0ts0jTAMq1ASl6GdOeeUrIV
wIYYSE6vOyl7LkiL2xUUd+xbUjAXFOgUxCVIKj5Uf0PSDLcHxLSxkZ3EhXa/CxgR
3Si1QxJ6Bn1CM905U5P82IsgWfM0AOw1fVObDo/CIAZmmBAK+VTlzlGCMmqo0WpC
pAAeIvAfWKc1F5nmnsBvBZbulbz6Jn18oCCQpzCegWh40p9rQZd4KR85f5AI4dXE
jRxnQ3+Q6nOJrhcTrbloTrVwbGJ+9qb33gZG3beR/0F62TuyZSTAKiKXG7i2jgiO
axPG7lXY5E879CXz0kKwmWrl0skYEraqvNir34+32plZHaXJXRVcnpDfqBO7PzMi
22E8BkN65L1UhmZF+6MgeSxZJWSOLL+UP8xbmwhCenXXd2z09d0KM/EAmveyd3Ar
MBs0PlsZrigeeqjEuh6hlPOsSlbGXPzO+LfXmc1AJwd5F+4dr4N6Rk7Ov5fS3Lrp
hljBy/Fbv0G6njOHSf4Z+GWTL4uFOvfhrj/hDXZtIHeuDgSQ2lyZRmksFN2PkbRe
ESIMcXuFpJd/x5Y8yQp6pMxG1W8bbnQ78qHI1PcDeq1APFuI8UdAXkXOVPWDsHgi
tTjYXqXgiNEv23rVCKkU3nQ4FIun7e4x4ZXzAfGjE8y+193wDqmaa5agwtHWytFm
cby3TDAcYzuanlpFrpgxYDEPauBBJupqMFjdOg0Pk1KzpahQPR3ug5R9JP/ktEte
D/5B6mu+KrmQ5PTWGRkie7/fT+FTdn6iKgkmeYLQSaLJCNd3VCplVhdv7h2wmsNj
Sk9ecnmkYVFWKrsIHW79ismnBGZuNsQjhDZrR/JS63qCoudPKbLwv9LFz/FU0QOK
+ygnU6HwmEyiiGD1IY72oMPyY+NSYQN+ApG36TrrG5FFh3G+/H3oWdeIvshafLyj
p/quI4N1S2Y6TNjYwsqSkufio9Ot+QJH14xzOfh6wWIdntFdxxER8WVXIYaDzSRG
nC+JIkakUArso4nkGxkhwLkR8udEQBvPxfhAF1t4GNcA22CMU5vwDYOQz/+2RZ/X
/wrUl7zFMpPFr/DRSqcixUEPO/NSF5o3kqXoTlkeKL9LoqBAMO9Nh9+76geUEQBa
OpKp+2xSvaOtf6iCBoet2hY1w9CX0TTGwHY5TlgYup/rq70aAHge5sixiwyMsIux
Gjw41o08ZOuypNGAodZp9T4KLxuwAGXKFixJ1FfJQGQbbPyub9LcMoLWxr+b9w2m
HH+9Uve+k241yIC5OUDBxbpoVXWqop0hWDqTdowHlg7ejarCLSRFZFY7pAg5SOid
28YDZWwb2k/tz6cPvk0TmXoaE6b7o1bDhHEfzyLuotfsJWCub5oxakUNPRwpqkch
8RhejDRyCCIYgwODp6ghJ1gvUlSNcWF6OKZXhZEnNmTH01eppI9Q/DdRAMjd3rGW
iFMD9V1u8P395UcZYD2Ct1OCCxDyRmvCo0wzcThVuzOmIW8JLMDi361XYvbPHaVi
PX55eZ9291xnbmGweJg87Adq2hNpBSPpD8rRIl3kEjyKMQG+nLMAKc34GIFImEd2
tksdAufso/wVz1LLtKQOzs/LzNtTssN0O/vTThYfR+o0ShXmV3bCc1zgR+ixo7wA
Nv8vl0Ns2RhD0opA6dRH11+f0MVN43DNGJjjaenEWZRsqpQQS3Wrq2RPtDZRhdYS
WTvU2WoOVklhTxVO91baweiBTAXfq2szJnxFjC01Euk/BrfLCSd3Fsm3dTCBjyIe
pl92kn8ISx/rM8xdTxlwhn3uPhtNvZLLfxTZjjkJ/yCfgyqsuW/MJldlKsMKoC+M
OZRIY+Au75O6l0Oi4BTqWaEinKrxy4AL+04ajES2upYLmJYhKS1pcQUkApBFsBqG
X1fftIHSOXERGUv46ScmLGWhhLdfBDxmarcllCTjshLgpHpD5asncaPB+m90u+rJ
jkcITAJFQCE3xJ8JgsxUnmc7ZCotWRLQ7jb1y+fwhYYLUS4jwPfROG5TXAPciikE
Rw6M0YDU3BJ1ps2mzMkfGuwGOX6bkRyOvGfw12rOhMBpTRRJqppelQ9wAcrodR2I
ovrGGQF0sCnHqvx9KMzhd+VAi0ckVHU8FOA63gHbTncCFuv7ahz4iEJZOKJr3YBq
7H/5jtA6LRuKY0ca1NZaMGrhBoBVAuLypdyi5T6lqYz2fDSsV6Kr2rBluEFBbeHa
lHhriNoIFBAZGUsk6RpwQPH7PRhN2uY3g6SsGOTEj/J4LGYjuCw+FEjfi4wUgSRw
1NxzNryAxeHboE/q5KZSIb7iS9HI5XkBEip3R8Q235hYyYgTcwP6KK5MyH4cfxA0
YjPTit/dXM8XE10gB9ul5wfSIMA4uaInBTSu/EDOXhRl+PeiyMVnViZwWxzMYONk
YFw/3RKNxZ0U6JclhwuV37iaYBSAoN9smxHTZJh1sVPvG0VCmhp5FS6pb01A8f4X
NDoatntyh5kgjyoRHxokrlcBofXJ5q+JnQXnCG8PHYzl52qjPqSBqxKc4RfklqU+
2b0RzvhuZkY4Ke+OVM7IYx5BmQ2k7mC1RpVo09jQMaiuIVBNiFdo2cvEf/Pqzy1x
q6ryUL9PgD+vm94hZKOWKuNSq8jMfTmu+gzGrfGJbxhHo0sMlA9B4myduNqVjmVP
WXztUaK0/mLbxwcf5FuymNv39t+UJnvRXvK5eu3Cl/owyNsOfbCl1Uklxz7ijOlE
PVKoYxyhEwUZwGdXntR4fL2iJa+1QGb9n6/CbAwaufzXApWFmyiG2xFAbvQiz+Df
YhstGkI8D+IxUc31FawBzKU5+yTxuj90HbmvzLpAVgTGDU+nSE8XIPJz3GvPe0zp
imCMMPiVDfoeYgQxOBQDEdtUmOR8Svcz0VGqwIXJOgLWAhdFOVawe90ivQie7XxM
S35qdTeM3oGFMUwOiD9CKcfd0dnb7IaCjYbgkau1omH28o1coPzrj3UwKcLy7Ugk
XQfs6dpEuO1kKe4HEpqqjpRUWoHpB82iB6s/Y2l4dFvhf9u6yVnKCfpCiTdgwCOo
xAtm5+2VNde48+cpdvK1SfP1Y4nAJoBcCZy8AKt7t0u0odZO7YgVkWT3QdDbNQwJ
aiqeEYLqTosdLXxqFEHeSVyYOAJ8EhijMvcnpNt6moWYhY6cYa3EAd7s9Sh8Wvax
IN90i14il/YwjSw/nvIA8jH5tC9ZA7W4B0/0VAWU5G2aKRxR+fo4902E8Vf8c1Gv
kmjkzeO4eXu2ZAILCjlUJ4LFp+XLxGEYbPQ6q8q9E2PDN1wHwv8XuyW32z5lfn6n
XcydiNHoMnjtOOqHPnruJWXnG4BKVRbsRNH3gQaWS1baTCVSr1m8W3tFNoWwZdaI
v59mDMXcVdqrO8fJOrSAGwPF8icFCmdQE21uyBsrwgMh3M1w8Y40EsZb8trEN3bU
cuWevGO1uYiwdfiQnbsHDKKGxQ2vIsEvrQw0NxG1JFXyd4nlgkycAmCjnE39vQoR
LjgEFWr/zy5gyNYbUtQKpJu1CG0jCKNsEzufqaytSxt2L1Y6ReBWZdn++LRhJa+A
+vb99dWMdCK+EJuDdYiRkrECV2V7ZAcUfs/+I4q2rdRDsMcAANLvW+Uf9AP/jdKJ
wVfYwAbeF2Z3YFG3vnH27go3jci7XPHeLr2rWxJQ9HztK/QR6u6nW8g5nrGyowOF
cy5p88vCWPhhrGIDiTeRe5qsOmOGUpnmLIAsWRqAWm+3gRCRYSEyHLmIsKwZPpXd
zM3PasmMSB3hnXJyY11AAUc/trXlMdGVJW14ioRWH/eufahuwm2+qLJ84sUNKQ8n
sb09xhesDyTHyw/p5Q2HisyXN0N9YTTpxi38V02+hRHKG6lRRFwJ69Nejnb9odLj
9wbheRjLueWtoL8Nf0JKKa6aT356W6o+4SIK60Lw7QEZdvkLChNEysE1b4L/chaq
q5Wf6wbvOYxXR4w28xQAYeW9vYylDmpPuc8gx5gHN+4wfEvfSqQPdH2R9HtKB6gX
ZZnLbUvaiZ7JuKIt23syZIS/naCCxhDWm/VNMSoQAb2ct/lCm0j4mlm1Frzmmv4q
UDQ+lnWcz1GDz5S9IZSmkgP5fDcFRyWLj75/K57thOUfQeNvZRIBo/XAsAHSgsCD
2g3TiyrGu3NZi/XAzpNBk3Jydbfqhf1zroE/eEvnuQIPoijYxqG1tWeBl3W9A8Qn
xdqf/rOxgUBI9uP3pGgfS5Eb8A5YQEYJQJ0o/JolaN5nwCbqyMxXwEAarfwQ6ty/
Io/slYrHQKF0o8e9qKP8Qs+EbhInQylkHBDplYoc97+bE/SDbTkkDcgM0hfvcX9P
eyjUfbYDE3QdJzxc44x1KnXVyABc/OZxpSMEnF8nTFg7Wa//SBU455dAhaGJMXUd
rPfj/j1qqLgYo3kDdU3asCNHc/KG7KbPXOFsHEeZlM9cWfft8T3mIUdtlilPjVJo
VGSAR1sEo9mYYN+4+M27X5Mb/1Tk9Ts8b/GvNwf7zo5O1gEQ1dmEh73PTd/0cS14
h11BVFUUftRj+S8cgVk/uiI2+4Dt44g+Hl0fkycxrlUZZIIxdXK2ZVA9qxurOUJY
53hsXb/7JCh0I2Js4G2ovxBrMf/vZT+zslNK/QKYrfACnvXfbudmjQnvVZyJCIAm
0MtdItKP+n17odhT048Sqvsh04dygJEk+bliXoZjvm85Jnh/7Mc4idL3/Syqh9Qz
Pi//CXdVSRosv4Ic0MX0rPcmoDUQzTku2X6vB8mXJyz+DcMIGfdOZ3wtpg8ZDBif
EMgXSW8F2hTLrGHea057jYQAfzsBtNv8Mp6D4B4zdffi4rtkyRu76YcVpYFk/B/H
rExVukHkmu4UCGXTgCP9ei5pjZ8tuHS8d+vcbOAK76ktReqLHPtC/WzfviBA0B+w
eiN7N/bMfVz9BIUaLhuxvJie85bPwTQnp9C+BOz0QzuDVN3I/C/IT0TX3lhNZ38J
aNoKgymrPKvXvR9l0myA2y2hPxZm36D88mhQnxqqfsmQN41CxwT215AqPt+3A95E
bRqCWAlqFQ0ffvvuqodc2XsgJwOFrwhY5VV68c+KdGeh1BS3CC3kb47+s59gZR3Q
q5R6fkvY+2Eo5sthrx9BCxzbShG1fKOEjttW+llF/3IsHtLKxayc9y6R9aWKC7NT
8Tlz5XiIoteXT5Tc7Yku1VLEeJo0OuyFrqKh3qGb+plKQEcjl+3mO/rf2CDwDX1r
UiLYepeX1CcMdMNlvbGUGuTHfdLJqeEdsjOkmcLQXOfV8Lnmo8rR52CzGtEQWSnN
jZ39Xf/h4lKsO/cA03m1UH21JgWMYDl8eFGF/nBWrWApolSJaXAf8xmLKBh3G4t1
f/qTtgJTJpHKufa5VLsl8zPPXdoLkIJEB+X6jiNUCeXai93MKoNRe7xg2frT2qw2
6O3Jk7qaOg17cVB0jcMVoBMlwenFCj9B8mRM3YhTnji1yTYfxqebPibCKZT094qR
ZYpIHPAcme36ydlGIIsGvv2ePnhgcluntSn3wyPGS09vEN07dQ765dpU8F4yCats
SNFBiAg9EJoJ0Y/fwbQlN0t2P1FthYR2s0BzT8Fu514rNs7rYsuzTV7voerLu+ES
5vJSjqoirRpYhQauCuDladF1RUxl9BoFCtnsnGkqN5XPCoRHiFlRhV6T79mH37B/
UGKD49EbWaIuqYaXYN1VVhKvGNAgiVzz/QcKNE3l0cyDu60hvczKPCzVNsYtJNdW
PyEv3TSFihp/RJLHuoN4BiLj2oHDJo7pW4e5AZx9mtHYGTYnvrsCWuC4BceJ4JM8
VET/v8fyhzVTEn4njJXrDHfIR1CKdoOTJ+gRlX9rr2eP8/+B8XhkncFJ7/bUdsg4
Bq6B9uHeG5VrJyAMuUGpYGhRXqM99UdxtcImjc5f9IagCFth0KDj1Nzk+RGo0ajs
mPmApaQ4xnEwwhz4wJyRifehV+qhYOYQkYaa0T4mzDU8sPVQRiobOBA68Gopl8Z5
9VyynUPjXoK6m7PKpBPkjRWdhVMflQ4sLosqj0TjU81lRZuTG8/U159HE42ZZKjd
O2BBcudCcH13desgbC+UPjYO2SEhHQGiGvaewH4O9uH2okJJ/T0Jbd2uZ/aXoKYw
7zsNSOCiJm5Z3LOBgr3PgtPquG6ZO68lZhYxpLKBmdK9A7ysXBAjyOYK4hqNm6ZI
biYntkElS39r2Mdyp0WJxAwPc06XLYcn1fym5LUu0wrwQPPvWUtHqo/GA9LHm1ii
gHK5n/Z7KP/nbWqKvombxlJctX8enkGJhzLxcR3/GLtruAFshHE8GDsC9IVFrC3r
b+YGltXiqnlz1eGG/YlizwwhBLAwpIDxe4irwznsOr8iAyJDvYm3AUk3KJjUfkqF
PtCRygnoP6cwqZsPYFOHsXfhNoZcqdKB0zwQknD0336uSIj4GCjY4tElrAo7YX6+
c+hekoTSOl+bkTx3U+i58A4D7gJ2FLib5gyliLv1I53K+I6cJD+7cOUy+QKmSsTP
Ai6cCUQdv0O6KRKi2AqsdKvLejfEb4MnH3qkMOiv/BRYW+AboO4+gD/6XLzS4eGO
YAhtB5BzG046wdbUY+6jQIpKkCUmdnZo/Ev3xzK44cyu/cvo2OVPHSzyDI5OyQYL
m0bitCChCxc/Fcp+AAXoqyZ76GxuSD+BKgru60dKLUG0SODKEKOO+Lj/5JelJBZf
dZ5k2fRKRyafIbjkkwf8nLSXiXscPS7lgzP6HUBbdVVryMn4BqVz6pRkI3PcWJ9C
b64T5f/cnD6cmoZDSWsFZqD4j8DPwvuRtpD2WErw2m2r8iagXOCWxK5GcZQpQ3sr
33Kf2hkv41yKA6LJMPhPxkY61RA4l0+K8jR6CbNPRELOsV9q3At2wYsrKKFRjqRa
13i/hIg5AWmVChA8/lNBSyxsiP/QeGlC1uZQ+05D+SnXxfar3OAdApiKMmLq5SbA
odg7FoB7s2nUmMuPckwTqof6bULEY3LkJaZKzy2sAwnK4S+Vz9q8oItzpvwzS+NA
skO6fn9xuRUJuUa5RLvVcyCzboP/qNoLIKo/8CGnu5pUXExm1bXrStd+eFj4Kboo
y4s1I2OSKDGJmM/cd6Rx4+vRHYqZ83yqZW3Ho1V8D0hZtY2Z82GRp9NCutDhpsIp
ZoP3gsLNYxWmkbCSh/FBiP3ceKJRryr2R4hkpz1Byr/5Wuy/yO84FjjwKW5Ft0hB
OyPKbzA4SSZAi6vnkThl5L6/3dY1wqb/2yUE5gbzc7eMyQ5zSQHxltZ/1YVuvzte
1JIQaJB3D8QfZVQ9sgHfHQ/MQjmFwPcYkd74zpjO0g6mUsA6TAP+v2kKEKLDMYZS
EJtOHM0aKccDSrHSv8aX2TzUoFa4PJikAxmbQGti+dZfgzujM/2b9YCQF1H4IJdv
pEQ+M6vBLvsmoUbc/kPbcTlvDdvlf4+dLIUvDtsDSKC9PonwtdtDEjlXOKF8VVZm
bQ0aCEnVHr6VwCNMEs5n21nTxSQl2vAOdwKS13YC4H475qgs96F88GuivmEGsr/C
e6uRbJ4sPT/S7IK6uHF0Id4GIilunb0GH3a8bG2/d+qGPmXAgqBBZj5FU/lGY7It
NdwehejKKPyTDnA8kL+LmWoDyNWSNW/M9M7oFtfl0LKSDWwKaf1uRAQiN/VBisLl
JfqSr5aNMgk1UpGEAyLq0Nwp2ilI6YOdxsZ3t+tCzeSjE/h/5Z6L0feve2hXYWUX
kqeFy8jUxLI7fBlaPNN9rwsnAwqBFYulRe+t2h71SsBYNb8/HrVrDDPOsydIs5cE
7m8jV+8oTRwKHmpfqCzbxV6eHQIqLr4+Y94oC6KeS3N9uMEuhwyjlRDmVMGHuz3L
QK2PkiUj3LphKDiigvkdM7cKVTtslkoH/KGARBYKtTiISudvlFNo1iK91w1WnS1+
vpjMKrK9HQxEYJAeL1HcWQ2Khw3BpnmI81NIIo4g/3DosEU8MymxuN4ICQau4i0t
DNq8X0nzbG1Uia4PQIiNFGWWaUCAC7yCcK3pajJtdHxbK1MIYyCpZfYI0mAdy/Va
YJ/ROOTV9sOmbBpTVKiwnMhaHIeDTe0hMeRB9skor2kV+8PfC8PxuhM8poOT8DIB
EioQtajvKztkjSBuEC5mvxolegBqyl7Seqliyd8PdvCeRb1RmqlyQ0bmWXjPsPC1
hKgPy/Fe1CWXn9dU1V66rhbQPx3vra621fJamVjinyNE2Oehqxaxb1D6qAl1WD1A
b0BKXYEt7lePBgfTO3xyiRL+YhMKdnBO2eOSGl1i4NtPfV5zRz4b0/hOiav4Ooqb
9q/MH95dobi2Z3v45rlBQ6wCfr/oJXN2X98XrCcj8Vri+HEwGwtcAyisedOl7xQH
s+/hVs/pVGGfv3nmqMPWVa2xNtvG+K8ThATcuEYupds/TtcJIqbtTghVaDSclKrM
Sv/5bsgwyCXm2IjJqd/+b9SLo0hqzQ2joJkicanDr1drhOW/AAGeRMe4+rdePxGP
zfIkb7d1p/GN31ExfbQqtfeiNkNrwxH9XQG1Vfc0FX40ABXQqqpNW06maeyDHDkH
4LWtqXVgYvCgM7Ylh0H7D0tQzs/vP4mMiqsja5rZXnITjmq+RBZ5ylnbJ3e2cAo/
bISXWunwchUBj7WgEXQJLU0L2cY5s/3O2DSZXh20PsJEOgHeLmBf+f15b7NOG4N+
eMFcQxc1ZboEE8pPsdej/JkrtrX7nzS1UZ3hXbAH3O0IR+8STRAxumqj59sTak1R
rzrVnJKBETVMv+stGosH3gy1SsrW3F7+E2K5uxhjODBf2QVCtVUykd6C0pCdQSwq
jD/Rqj7gkEmxqOBUUhHPDXxq90cFOGyfiIVmEVxXfkNO8lHW9IOkn+W+DcZgkoEW
FKDu8L0JJWDk8tF/RS+KqFKnWboM8GIEuGVdB3eFqxG/lW8RNQTO6am48YuQ7hQY
41F/4OI8IbsGS4c6jwL84oXweiEM+Ppi6dTpLoIUkQB/jucm1feQ1sEDc8AlxnMv
QUAjBxwFImyv6hX2PmkjoSrmb1cV7+/d1G+a91WzNlqpy70PFQY4R28sgVRPv8wP
v12Qzr04K0oq/gPjH4vKwfdfcvqT2dPaA5QDbAni+FzYmt6piajWz5qeDfpS9d9L
f08j3K1fl0M7/KqSKnLdSKoBIFzJA4DEzAinni6LBVq+KLzpYZz++3cM2AC2exF+
2KWZQmeXK3EqN+WFkHzTgP9Edi1LxgKsW8uC/980gGAgtNg85Kgtcf38kTPO6TvR
vguKVS/iPyCB2175T1QXLxrkOmUCASvOB6i6EViUXqtbgih+TLyE1xM/LX2A7OAd
lCiNVwIJ5xRjFwfDDBNMIFqK4h9pI93SXnb/5QydcWGPopypxYixJCkJyNIFk7xC
EPCzyOL5FLz3CT8z76ckcXIjUEC3Ix/oS8HFirL1BV+ImXXjC6pZhRoBZ8JWqjb4
JLdX0kPtxjBhowQ17Rm7QQY2Zb4b32WH8btud8UUDCgCoxiA8ZrfpaDD6jIB5LlR
WmdAzhfKZysquMuosg/8V/M8k9+fuWFaHHNnYgddZteg9Mn/xSpRopW3ZtxONTH4
JY/5JA3npbrCyrrOVAsDpKmEYmLy9Pn5vDopyaXQebr73O/XnTJJYRV6Ad14sQ+c
k8BtZIWMxfOKHorxK+oqnnhvJuF/f/55NHo7vs9MxvA7cG//3I80iViqOFmcutkB
R9SOHPMJvOEItCCcaubDfJGNdQCSw5rdD17ZfG0Cgd/dL+6OaYma9M5/8ECzNw77
Di5eyndmFztxxHINWlbhfxvw5KRm3V80u4eEUW2eeCfmgzgpn0x1AZp/suAwTk9r
JVvBW2Q8F4/WySg/GHVfCx6Hbjn9d/shTkOW9kH3KfzBJzPDGNJi1kZjitLyuoee
1rD7U7bMAIg4L+eY3l8xPmGKNuC6GIGDVEQR4q9tu+xzdHCPkGggz4HYLIY0OD6y
3z9IalyyVlS4Hro1nR5MlOhdKgBDthJpXTMmUz3RrOaQhyijtLxmAMBiFPAA0ONM
KA3c7uwXpSqXxqWfDDmdAGzBtRasRpbjft3U55XMwZQ0ZCyX6nuNES0NnKWVbTb2
Zn+C12RMw5z82gyb2STV7dILN4p9YHGvGP/KkHB4nIw+Mx87cM083NFkrbij67ox
3yCKEOzLR3JnZ1xTYdB6hXiRIpWNFbXhMnJJ4FTW+yK0CveJxPf3KSF92WXcV6Jo
1poMUfbnI3EXBZjxfCSEexL+3rnbi1pEwsP2XlaPCtu5Z0iSumAu1vSRbY2TFCwC
vdqd/UP/igX75mV9d34/UDfU86uRr+GYYNs8We2euv8LdctewWANy7lINqNRWQED
6XZpGs4UX6w9e4fWG3BYk1MMhxx3cxeLitTPyXugt7BVAeXOvc10QKgDgj8dIcrd
CoN4cKaQfqNGk1RQqMq8U/bvGuqKzIuLoGlwGG5nCtW3W/oyCpOxt8tReCvXP7qL
p2eVYI/xCCZ4wGkYtMtkxVmV41ffusBPTa9HNKWE+1c9uWQwuI/MMt1VdQ9Pq40x
OmQsOK5RDX5M8FI+i8x0OqIew5fPuhXdYBiGSkDYPaGKcE6+BF2MGyS2HlcKr9FH
mBt9iErOaCgS7pGz4PVTdI6SXyt80hcqahjz43JYkOvOQcfjs+V1Ojq5uGU3fd46
8Y22NpbNonXqMS3WKKiB1q0dvoBXDRqhmbEEl0r8VlRJgzzXR6WbtOFUlbST+xfd
ZsN++tP8Ss5FVnvcFBj3yNMkYlwjCE2f7hGIKL+nfEL43t/3luxnzEnbT15OVNZE
qMHG4jwSgXRQsdaED6HNgLALj/VV3ahDzgioo5GtrPWjid/t+HA9ZIPrN92Xqse6
RzG0LoC5XNajszl1qGkCGZZed6XgEtNgFHXqFg3H5pd2ZVZuvkkVf2p8Z7D43wgn
WoiSODFU1KZ9F2KlfQpjZ00bSwuL5SuBzwLYBGlLNFPHjFpLfBF9mqVxK1DQZUWF
k5xKFno9Gpj5kNVtQTIj1NnqVio5ot1MdStayddfkdP44i1mIgieHdYpjt67foqF
fMz/VeYSUrXWK+S57nTZy8rCT/gAmciG6jzLcOz8UwFRXXylK5RTyPjUqaGk0WQu
t/wWsDwMwH0gQ0JwRdhJn7sPVKQIGyNSB9N688wr8rVW14tXydnLQhDH2oXbxcSK
C54mPvts6wk7Np4eE5ZkKP+lL5/s/DvBaftywQRIqHo8mzpJ4B3zfg8WBLpzat4p
gmUJCWiomYumpKSgG1dD2QNCgtBkSpmnUP9tZ2qIoX+TdCPNpMyRKMRfKERJYzMN
xqDSpZEtqppsao+sN8PkRiKu/xnDOmlkPLSmQ+8frJ1DkM0Ep19QSn3qKiEkicAQ
ru1l7E/mkaZ7wFflK5Nitljq/t3YEns7jXpTchykVySM2ExP9Y5N/yocZHOWadKD
GgJ+JNq//1c4h1LD/Ujx8breemykW6ob1cFSkkJ2ZIucA1nr1JwV5IAVy1EHHwz5
SamrnK1uuReITF12rC7swXQDVObRdstjJqRzHABjaAh3+iUeHoeOElYol6snyqdE
YgHsfcwjQaUS5jFzper7Lsq+t3ErK6n00mZz1MhHvkZ0s52kTK7D/muwjEOzHJeZ
Mdg/AJl8mnDmg9PK8et3nOdf+rzNdEDA7pBdMDMWOSJ1E2RCdkMqmuzRyaGdcA7e
doUiW98S1T0ReENrzXAneXvn6SGDak9fhPjFfP78EL7Cf0tbrPekJbdHKdTfX2E4
pB5NQAU+Y2sNvfkpEEBkJIGvT9tp4KBZncyCrp09AZ5wUWvxQ8nB0MF3kYpEBVD7
ir6U5Cpn+NIYwz2x5ZEaBagNQ1ATYYEEFmkABgvfxOFfwm0jHIAuAM1CrJeuPtcp
4ip7onEjZmQZ1c+RE6aWH67eJybZTbjvUpW+kQ+ot3tz/viM6K5vBt6ekUA8qApf
SYprOwqVUGmNGaOaaRvrb1KFmRiM1YiybKRSFufV7C7Doc0DCcSp2ODWZL/znxwU
nLA72u7Hup9rRv/FbrvpLSfbAnz61YOEWy+Z935X3Ydh1L2Bd0EXKsBTD32S9SUK
8nLuGOcbgPFcg6791TgXR/tNsRO02IHNctGOau5u4U68EpfkOT0SBICh0mZUAVhv
MoUbtNVWHNYEJpk9u0hjtKwxHL5VzauFDxKH6nVSV5YovzNJps27aFJQKcWjPdF2
3zGZ8FQUaNSIcbbjnAr1mKW7Th+yvKJNBnuPCnLuSaQvyBEGNUj7p8xv4wniH7fp
lNEH2uuu21AkLqmR8Q4y1/fjIC9A6bwGEXWsc2yg2NpnIMJCUoSpUy2GW2ckqRwV
vupMMogPcQeIgHRs5h43wxr6cQRaHLtQCgHpZSrEdJRuRcC6wJrGBt+i3BVgGvie
HXbp1u7fsbxnWNJ4sSHD95zJZ4ihYnp46QQpup3LtsLY5GpGH8Kem9thrGLXvv5S
peSPVjn/EcZGAFJLNSDLPlLLofWVbsp2CXus6xd5AvMRVw4QDpMOPSlEZ2zGoxbl
DH8k/0Gk6zvhwnQFeq3DO2GaTnUDPVdm7UD35nZrnfnhw1ea+PprX3SJfkiBwroI
WcTSB6T8ao9TA2DTm7EtAR+59qLqHtRhcaZ8riZVJvOBBFy5odcYZcofmgSY31mi
JpfHEWFWV0AP3s/b3jp+vzBIReVxjXZ0rhyaSgGqICFXZiagONXdQwyt5xpqSGfY
jmqZ00LvO4qvmUL0Avt7/dLOECYAX0nrzgy1RJjhBZabwfB10D5vZgmHX8gN7uLr
QoXKMEoDOZNBWT4E+uFXp6JSmAt9v0pUUXaX0wZvtz1In8BB+xMASU2bk3uCRroX
1e2hL+MLPYCwPveSCLBgJExp22Q9pi/do3ADovIZeejJv8pPCmOVnO8opNypu6/3
GONIbhhqYo2tkI2jpevkrvcKwNVmrBT4930LtIkuYHlJ9Bv+Z90kV2U7uDCdOBIP
2rtKEDWrZ/4yOMXdRCTFrO42fXIrBnkVgYGQexIsCBghBDZa7wcsuIjsL3JeWfxK
+/xEJl63YtylkLZUPpIRrVkqaBNfD6NcQgfnZ/svk8fcCwenrlcydDH78i88V9Oh
AT7/w2D6vwDVtGkQcT2srqw3qInSNo6d7pVnhh8F5vy27KGY8TFVh8uit54EZagi
XHtYKxbHRbWvbS3TE6O107F6ftRI3GEQbg2oCZ6G3VtXCyynGyZpKf1RUm+AxFj8
pqRuIOiPylMmK/bwMF3cBhV3+DXDwnhP8WhK5noUr18h4MNBH72am4gKDGH3hWov
R6UKZ9zG6hP4AV0qjM55JFMucv9Q4CvzTCn+DfE9wJILpeJIQCbc1dDlcmJ2dS3O
hBYsoFYCWzxhrm4vhj5DVhIeXyFijZ62fsQewqg5GHdwx93cfM3TjpEtERcFgmqB
Qdsd+mIbn+QI0L/oVh8nMCwnqh5HtLYuhirzDx8pZQcpeOm9C39n5NgatH7sK3+9
CHtPR4j71oTKsefosOitKsyHBBpjmwD3mzqUZbq2Vf2Yw8ZL9TZ4We9oWUhFZfmC
nqpvR5DWSA4IvKCa5DomkcrBJ3FmRz7cnuXZ+OYY/gYCJIUW+jIRT0uWy8vxRGd9
GVxaw6lMq5dPQMd3Mr9zjq74UTnvhg23t9IcBKx/BsdWtrKy15fKHjgOiHkgnvVj
C/K1XihQ9oLwK7lwRVvjXNiRSiygZDNNkTGDksyUmIvwN13ePoLEsSysi5P4n41X
yY93DVVxoltBkpf4QG2lRYDGVxs2sWrI0j0ef/AUCt4CvZ2MMlW/AVS9cnHya4ub
1S/czCGReaqV10jq4Ji36+M+9aaaaOYfcZ9gN432mQNi6G1Nl8aT973MNQaz5cH6
05E+sJXTO2kbXccyq59C76fXHiSwUVYNrLZeJ5i5870yQGGEjWZxrOTttFlXp5nf
z0K9T1Dd09zWBMo/HljOJlqBV1Owdw2c+ayJUJr65TkUeRqQc6Z6RBOUJi9h69hT
7cyNf3cwIBtRkMgJuU/WzX+jJYanco2Gcn42vxvTTOkEro1jwWQUxV67grJ4yXE4
iItdG6Fpvi8GUBSCopIToe9Y1o2BkZuY5Cc90MWfr/oMOHvK/FXXbf0cpePMNtwk
6XjZqbfYJuWFTyYoYdRpxn3vMt/pmaKGYHcCABADdHVUaBAJF4/aSRd56Ss740Vx
wyBiUPkViuTlSSsTUnN8Q9EZ9S6Kv5C2IJkXl06xGpB59Q/Em7cVuJsMO55xmU8v
eV/k+Us1qovOr7mP2lw3L8omkHEefDFsGrgjBBc6UvuAO5/Tw6MXB5hHpuEGl4M2
aRwc8BBehSzDGzS0vXa2ntmKluqg4s3dkHq/RJbfonFsb9fBgzMSHSWIUqkCOu/7
8AlVIUlwCsW6L5Pkon1m5CMz2PseYZCq1t//zjUnjpl1TRQ4PCo1sITkX81yWIRd
lkKjhMnMhT/bN82/6CcnULz2JxXs4GLnrTCN75q0i9K48ZQMnFjWCdx7Gh6pSN4c
HVAItZOnXWbCKLJtEh5CeancAuvYglBYUH/hDb7GlSPTXd5NFdf9q2wGnGSWK+kc
LRKXoo9NGyVfYhWT+qIxYalvqd9e8yA5ZPlk1pbhaQUxhSHEUZUXTupkPuTsd2hd
+iXmdxoSxvITMsygE1+TWANpXwYbH/XEkH7R9hTmSZxxcBMAnREF+zyhrwckwhZ4
LbAgCBFZdfEgCOQVelKC+QIjlkeCUbiNIIVlG4DsvlvucviatEYEdhiW5kryCVZw
A6ktdKJxCH2CNCuVKFV5JmR+4NBMJT68buMG0Df1Vp9ZuckOk2Vca+/nPeSKHHt1
ndy+zXPamHF5oMSrYWNpaISUH4Y9mv3CurQhb3KeIaJK3IG4gw6gTm0LRy7VYari
/PJWeUXkAlX20pZRlf0tTsLUpR4IIc9XIU5IGTC+aNaNriOpZxZRTaIUO/Qt9Ygj
J6i5JCUZbmvFuznqA4DpkXu5Y4YdmhUzD1TyqzNti8AYwYJLiCzi6F/UYb0MsDhp
ow80HIjagDfJfDst3d49sHu+kOoo4Z0RoUWXYLxF5CmLjdB8Urvcg5Dah008fykW
LoQ+tUl++2hj7DbNj6fLevi01xUva5+O9k13ETXgcybNHd8MqfHXFlrr1HvFRia5
v3TLWAb0fzPZkb29qGBoKdasI3ASyw9OisFAk8/S9vw1a/xMlO4WwrfcYu8g2Ag7
THlbwp0ObYI/P2LBMOILnsTB2XA7pQIAz4byWC9DcWOmxW0wmj5lQQiCPF+aHyk8
docQgUmJ3PO9usKJcVqSuxTQp9JDgfWXXwPbXc+MtMM5NOUjjRDRax+QCUbY6gw8
0MRbqfvXsC5IPiJ43soYmJaESXZQ4sqBSPC9asijl8RILWvPKY1yUiJL9ybkFzFy
qjwJWIXku5NGrCs1oC6atX8zdM+oePFWwiHLhl3aCUYoLEccz2OFJRK0exUw3K/k
K85GqkPJrgpmzlEyagtWOkJx0sBXpX0mydLzY97MZbl5uVi6Rjov0jpzW0zoKDYz
dHXVswacoCx3QQ0dot85F+V5ci3KTiWBhj/J/Lnc4I8bAbBGPdXMVtRCQQjVAk6S
vH6V4ljPR7Vy0PFN9YQ0bsWDVcrpl/7tZkH6tELg2ZAtLY2yql+hxi/aOVoEorVg
Hujv5ztEesH82OohwfHIZL48bPmpkReYMbpWkbnbuU6FYqB/86J6F1WQnl90iWI2
SbsraoXX22snrf4TfjwvAgtpNCfhztsixOh9zqTqzvCSph1maxJMSNxKmzF+pPD+
P3iNfgf4o5A+HqYdfe2Qasij9ciR68NL31ZE9rhCUV0oV2iusHkbkmEIxZkDkfae
xdbjQxlcDVqK5ZLE0ag0KzDyYY7q27ji/wP+NYjslsXm5RkEKxjQ7fIeTqfBKiCb
HjB7UZ84GesqV708IgWHhphHrArVJ1Jp9byqgAsEfjNKBQ8GlDPrQ171nzez384D
L0SlCsrahAR+LhEDkhYbZz1YtwqDHqNqOk/7RbY7EnJKwiufukzGf1NqbRTR1QLr
tFOyfv/NkqFaPkKY7sozNJjIkT495sryU4QGyP5lEYv3axOYKcq0ZR80frqfi/CQ
D5YkCy/e46JAMmo8VWqyj9qAChNnYi1l7lMd85CBeZssgqhCIf+kwEvugx496Q7W
veFjv/ZbGk8fvk/O54ilgQsds3bVsyC6w5QO4PICD43wRtpjdTwt7VkLlrB8G5X2
7+wEC3nVygdzqrYce0WcOp8EmXYwdn08fwiSLymr8C+XRTUAlanf7Ke8Dd6lbcef
F63Gmh7md5rPhe6Jz5zMGe2MJD/7NLExHU6IGmmPapTqwpT64r+ns+rFSgD0gvpV
n/LRykhhSR4RWZ3i9Nre4VU9JBfbJsvQSjnOeGmQLHq2iSUrtsxYkyZ7xb3pUU5R
nWBZhS+qXifF3Y+abEJna6Lg9gG9Czxfox8vG2QiV2d1K0fnjaNKs1aAZ2ROFHvU
pNXqkOMwsSB1YftqJPT1NICDV2hJEw9ANKU8JgkwS7PLlazwjr3blAmy16KqmurW
Yel3WWUhJR3Q1Oa6MV7UPGmjR04SPgOLK4KGnbcDYGXJI1HTB5KghUEN/bOA+7HP
jx0tB5wBbb2tRW6tIgdqUZgVoYBary+6PUFS2WIfPYabcUVQR9FwdThtE9yyJJOi
qFmlHqRtgwu1vK6SPKMBIQDI7Dgyi2tj0b1fway8LAd/87JZCyH0kRCaNWRFdDT3
Illma5OfNNk5nT2RAK7ocdcTY5wACceNZ6AT3g052lzQlrc5CS7N1bj721s9jila
JVK7cTEN+esxRpLbmvap8WqPnupOPCYorAmuABx9cFl2lbS1qFozHJtJXegGLWvM
YZQCCl93hZnudTAevicUAk86giKtg1DCFOQqG+x71r+dshEciVwozlpDeRaHq4fP
8tUZwgvHd9/PY/EXV04hHzD8BBTfgCXQGw6Gzj62apHGygEwAF0xHWGZsgRg+Hrd
Xl/9pSAAxPip9gjDo1ArEMAt6266n+Bu6YKk9vFTbnb3s+KsydBLIjhCjlLSSCiN
oYapjNk3Wn4a+rQMNyk8gM0SvTNr+Dw1YX9xEO8AuxZ3NvCyFnyGXXzuTN/3x5YW
Etrtp1Zek/uUiiI4C89cjmLdqYooPungbbqvnDBQQOuilfJEuWN4+UqP1Gryseaw
hPdSbX5aO9OzOvXlVrJqkmReMZ9q9mgAkUizw8VHHwgpiTZ7oYMstzw41q2UE4FZ
tKM3POrgYncaOEB81FtxlkQr0SGr7XZMgzRKG77uuB1RaHlUI6Ue2fUPAFx6EYea
YLb5OqGzJpqB+Hs6o1CLx38P76CxKs/JP+YqdQQqGN/Du8OfESAsnbZWQh0qGS+q
Qo41q6WR9NA5qIQoceFWoCgE2rFETOKkMK13SXUOlZQErdttsx00noWcyqR+k4db
Ws9tkUEYlnF7f+2UGkjZxu4DGJmBC49mAq5HRTNkOYQRpLnRZVm5nnS87K35lANE
lDoYzfxRrcblVSWWauaEaA0K50c1fu9HeuKUi7W75MHvFAx2E3RxWoXkI9KVlz7B
UrAqaI7K9Z/FlRcF7q8IMd7Q7fG+1WR96Q2hV1TaWjoSxP1zrNoE+C53K+rWfGZe
J97RUUoc0m3jbtcirQtXaR0/ytIVolzQg/vO5EO9dzbdW6yRMjB0Zq5+raxqArVQ
LvWkMxVb6JNjH+quo0dDbY+RMw9PY8e4qEsIE5d0ZGDhpkEueDt/AOnNOnidLxk9
C350NvZlmmDdveDjkLd1nu/vJXmjuKAp4wc/d0JWyr9F01yRfyq6tf9VqDAb1SOC
VmYVOphZobUycJDzgIpfDuUBDCvtK8WV+3JYbqM8m9O54oYkEEdU4a6E8WSk0EFM
fmZxNExqMN+j9bdn0n2hkVFVnQXsVZXKV7xNmWUvMDUOigGNIagdfWySmEjqs0IT
/Sg7Ea1+zl/OsTZC6KUdzWk6RhU/trVlMNL1UNz2kD5445eDnyBkYF9/Y05TzdzW
Y7rt3xmd96RPLiAnNGMh8qIs+1asKS9zpXs9kFGOaJBpSM+2DoAJZPm91EVgWhoj
d6Uc+yQ499k+0dFG9ehTQmgv+tnXSatzvN/dXeQbCTDef/l96VQgqy0ehNrp6hAH
0GPPCKxrg/rb2JvcgXEas/J5k+zinEtYavIAHFGbMnngA7rY4ShFLyTkZrBAVPj/
tV+8JLTcQpqau/emjlmUaRLzSTpFKGvEpGI8uBEQWN+QHQAc1IFq/XZh2w0NeVkt
axkZsGh/YMScBy+ny6JhqZXJmLYM2Ti6aYQ/WSePE9vdonzImeJSKmtyV4C5WFAu
DBhlH1FV2mbwGtLpCpKt/6WowiPy0HquCYKfm4cMvgF66oKEY0dcBvU5++eXFUMN
zJPganHxonts8R26rWUx4jMW3a6NsvfAfBCuSu6Ks6m/IjTlj3kj0YnAPBgMuhw4
4kKAexVF7I/aJcQ1Dh4oWrS3EmBYx7ay25N9Rs75f+QcWuiDsrswVOyypBFkOFbW
oFUdvNjcBt9lSoExcH1JgHICMhc/SmATyj8L56WIBaowYFN1pmLFCjfXoXGQqBqG
A/NGgLIdgHWR9DmLJMvlneE8bgrq6mI0Zl7TpkASKYYzwJyyfHC+AIHd3+mmxjcp
76rlmHgh1e+e8YLFeVkI3NWw8fLo4L0e/6qqn+Tr6pYi6bh5La7QeBQI7YonS64z
TnyPa7PG6mqr6oCNlbznNXf4EQ877t6VpVtZIUyDxr5Dw+3gtdA59MMj9QpBE0wd
XoXo+mAjG6WiN2BLAc7Ae/yPBp6JQSI7La/NZZhvtCgNKHK/5QverTehZpPO8tQW
iFodyuq0y1hXqhvKULyECKq3RxYHwEBAk0f8Y2GV2U6Z96e5QcXpWEHGKXLiB5aR
sgpMlXP60aUh/ibIy+BEhrozAQoFMex4ISHTdL8ZrLqG02vQmpRr2HsDTF7ha7ju
bc4zBODwaWd8DhaWRlqe1khF2biRwheHXqAgW43REAVB9s6cLkpoB4et7v/pI8Un
riB5NX1LF8WQsrXHfUeexbS6sq0Xs+r9WKuOsa5YbsUm6yGr4AT7xmo12caDhp3D
SRW8gsyBHRkn4uEGOPHhhAfXu99V6b9lg6BREgptz04Zme/PSifatu0YRyIpT2s/
ylN4NOynqgCNh7LiK7AvPAsyNVHS5NXY7yx8up4IVwznhUKaL4K87WrgnLKnWfh5
CjPWRLtbm1NweVSGyPZzggCqKVNofBA7fl9DRh6iDQ0U/LWOFJ5YQZWcnrNWNdOM
ETt/kO9GogSvpDRFGH9RD+Z2CJvToNBFlvZ0rtHjMzM5KGu7DM75M/O+4SEulOYH
TaUmavaEtdmXqKZSNxL93nCQbIFB+jjktyoWhDFz2k3hJvnxyN9wvZ6/ccioRlxy
/CmveOM8BQ+eTqmE4QbcxyiZJ35Lnox4KVm9oSWs/SzAdiifDHCofj1gN5+x7HaT
IvKYgtl7IM/5c2GN8W/j7AA/oNlfoNehbtj2LRiP/cVkUeFSOPbHJ/tLRBeFjYlE
VfjRvydDMXJfmhI4zKG3tmAt8ZMlNo4Qukqe8XFH7LhCALRYX1g4y7esxgrQEE8b
VXczeMGY453GjW0j5LPsM65clBHylI2MI9aR4AllkkpKHBahn/ZSa442Uuu2sCiS
FbUsqwZ+gUGq3WxjuLrS9zVz6bjchuRgz8ZOrd/sLGTagT419p2YdUeCtDsnLqOc
V6z8E/4J5ryMkFncS1KZVVX+0XuRqUVi8j8AIIbOucJM2f2LtWvCrfWgCofilmQH
jTt6POT+DFrLsTrGjtAOIactpRvbwbaNhDZba6Cz/UgpGsGYr9nc6EVrddkGCfTv
toFN0IC9IfRmjfZepC9/gnIlaKdlMptODJogxJsf7apCDtH+uKKFf2kSxUmJkJyi
8nQNNPEWutUcFQfcxs09+c9rmBfq6hLDNX2ilHcaqEkDNanaAIVbol8XO7ac39td
wMvUK+PJLnXdSDEhqF7EdiLbcNbDrfD0vvd6lQ7vkqT63RvxSZrqLH/k4fvNOGK5
24RFtd3ddRZtYlKfOU+Qo/JXwdmGUZtC/2ChHPW+3kd92/8kSP4SrufVfNXHfAv4
TZVmA8uWzBxBx90kaQ/1vxtPv6DkKexWWyBQwg03MtZ9Cj4NGSc5QGR3Tl9cDciu
TkgSxh7r3QiMuAEJ4OpqS5iO61tW5Mn2qcYsIKd//F8Nto2VqSAbqF1nZdyimnH9
Q+nuIHj+zEmxOxahrpIgAnayFE9iulpI7GKdwdWygcAPnXWHBC2IdnXhHhqqLrcC
O8o7h31NtnhQkwDRtfbstIiMrZGWLraWedfGnM6QkjUCMxKUhGHpSQ7HZHYkcUgv
TDYPS/ZlFWeJdg4FzuXXJakj310XX7T4GWrA3PBVVrJ7RKV+Io21L5LjvMDdfRiB
/O2UQyoTIeSGRynaV92ltq9imnsik7iGqtwpIaVDQIUIIgC7lrDEsB7oZJa5z2Kn
oj5Mc67FIYaSno5oiFMBDkyGpUhtwj/VAvX/VgptRJytTlEFRDaqPWi8kTO49VNA
ArRReOHFO8WSCU2MB4NbKD8xtinDCeVR8IR+34I39C4BGyRBV/CNCenyp1wqQfle
xzvLRPL7D6A0D2eGrhE3EMUumZ6ilyexz+iKCCwueE5doyXf0ldn/8oJ8dd5JqDU
5G1IgvXzt5Q/V7fvxd+BIcOUlRCe6iG1FWlitY4QNjQBDCJPN870CI8gaPQxa69+
cgGEs1ar7eXDYqQVrcjLcCy6sZKs2g8+4+Z8plonXVv7dv5lMjp23y9+fvwrr7jb
95pLRkvuTjpKJvSFMu+mOitRb1F58iSvgDkBNb8trebEFQkTOiLi+R6PVtQdifJp
BhF4aMg/IdA6J1o/66AQJPSe0vSeYI2lR4hD2RAomKw7PtNNr66q9IHH7nezrylL
8QWuxemNqVyZkT2Fc9qxdThr45BXsPxlagL0Q1oyNUFcHGo2uokXO5Iic+OerDg5
2D/ooAfeWdXbP6aDF/K4WZU48fppRoYAaQF0nBqHWH2v+B2pAfCYUrigiv91Xud7
bp0FvOB+5mtQnZQcYas2zxEkeUMwZqqSei0vemtqz/QneTJNl3WCosIp7hJ9jOcb
/du7wYT9zyWxUqFAoy5xwiRDiMQzGZhrHp+Igun9lzqxoSx5hjxoVCWwf0Em4X6c
WIDp//yQ3P60geoKO9kd63o7o+8rzBv+fykbuLmmWZFA8a7WVacHkRDOy+R9z7Ka
cypR+pLa5i7jBkgF6ZKABF4zREDgBN6XeN4sRm0nGIlrGM/iuuQZfP1S41QeFF6P
wPN2nwz6Ziwgp57+QHYM309S5ZPXIop4Qj7LMtThw/ohm2uy9+doopJmFFguSxdU
LZOl6rhxVkrs7sjvhaSti1aBbnviyvA3UUV0/dhMscid7+lDvTwlrCBeT4yYJAYb
lnxIyk9CJ5JUvSG6qCH4R7RrmMigFJYi91lY3Yh6he2wVU5FX4nOzOVY8o/EjX7m
7KQXQfFYIH4J2V4h2PBKteYD9ATiRKDk7oKnZ4Mktgeu0qicOuJChas5ZOFUzuaC
vbUCKKzsOT6b+DYwTv5eryQ09jsrDN3CL/3/6C7YCGo0mlrO1GwwR8jiyKbG4Oi8
7v7KyAEGZx9uCraUztdsbQaJgnqc7TnpfSa25EexeFP4RDjSj6bbhAaxj1eBCR3o
kPJjfilKBReyz0aztE9FB9yAC6tf3jakLBZC40A6dTWhkmyMBc8eZygJWuWDt3Fo
0iyYXlS0xlMqCngS4viH0YXch8WZj8cnqD/yFoMqWvRVo0jICqZxxFiy0/4GiuMM
jf8LzbDTs+rvckcqfSL9mJVbja7wsn0Eb5rly0LBPEg6PVTemZjnQ1qEB7N521MH
sCwGvqH3ZMzYUPQiyfAwA6PIyq2YpWGCxo3eFEbDV/nwqDG3X+cbNE3MIQACOdHW
n3libR3RRBHW0mxyydE969hb76UsR0ZfcuB6TlkeF0V6Oktjkf+4Q8PEAPqmrfqO
I5kau0mcG8lnAlq/mjNC1gT5TSt2MBD6svDntUHF+x4iLAufaTSMQWehVE/eAd0M
5pMUeSLRnYByr+4SEMx8vmy+I1tMxoqPLLk/NrbmUuhER7dFq7EZk1WDXagQGsW1
0DE2OKmAQIKCgcBdHDrtg6PdF6tw/dXnqetHszET6XjlQVUTtlqEY8LQhGXec251
tThQgos+I3sv53J1aPHDT8JDiXmZATUZ+61gk5z05sLMTSXMzEhRBEzRPuHfFs+2
9cCwF9A7i5UrQ72sXPaKN/1X1yPm0qlJK6GMBI1aQQo+B5oZrm6BpnGg4MS9kda1
cQ/qVttRUnisPV2DHf1P8zge8lUQv3IVMzDwKoRm3d/tWwMxpKbfQnwONOdlW1eO
EJ4a7jPrVTIAvrdpedTRuQzlpnTHIsCF0xAZgzZl2BBqQzdWsXTB2b8UlS2tpuae
UGW07Xas/sCqd49D1iSSZ5NWUCJ6kTdvDYrfYy3TGgh4YQYliLS275j9RRDvpHbO
y63MXl+oWU6axwpbrqoa3mSC6QXdN8f8TG/5jo4yQ80txzf99rLdsnxxaRI0Qh89
iHdGm+x2EfxA10jkG+H+Vi3ubppQI3kuIIsWWM7OuOCRMJhM/yQeNKYCJMM/n+Mc
MxOFtWsjyrAjPy0IC+PVvZPb1e91Vdp6R2vfdf4U6oOuxc0Jj1ixG+1QaYVoXyGI
B6R8L6CNJhErm4DKx3TEonlADxadjTOJa8WJN+d2Rx/bDo4bAC/7ixRdDZZFKif7
ovNSQKAPUmbA23ws7we0PTjbScDT9AO0xjukMitDiw4mCLb0Ro8KKojR3P/kFpBT
h79LsJduCzI15Wby+gbNm+waXY/yf8QgxW/zR1unODRVgVl16t0DCH+hnl8Xzxml
Z/x1PunIQoTA4T0vYaE/jV5zIZoOaTLsTuftCmoZbdBFTbDhkSy3ZuhF7DwWIOJX
L9bZkeA03g0JBIE7PMrQyB8zSDTr+yePpi/fuxkN7D/rzRoMivejgwiC35ZLP7vr
ivJud4lP8W+sUirjBcCz2fm28tXYUVMbJtABMV+8nw/LfjliEqyyiFQaxGy1OhH6
wKlcuysm6dDppqq+Vlwxvwew6fhKPdfK3MmDfmg2hroClivFH2ip5ai46inMgTJp
/khkiU9wom5ovps+KMJ2sD1+ZYPvyMEYAehg3z31OGWYobHeFS361l4m8nJvQ84C
wIu6GUZ08MT2mdy8iaFYxqQG9/q6EA4qUCNJO940rUDTT5MVNCDdogYzVvMvGcHB
rOdFAMtkKxZj9UmhAV7tuWvjOCTlQrsPJqLElyNIqhtUVv1j1O9bGIXr5m7C/oty
d2DulF8blLMFcOEVXck6PzW0YxxShEHHqt0FAH2OEapvEASsFvVbe6a5OD5XFjk6
h6SdEr5E8gR+bMjUFI6Wgj1OT00mMBHVqDtlhbr6shzbRX4I5OqU9t3CDg7wzt2H
FVmyZgxP6XcJmFhETLM4hiI8nJnmzj/n8Vn1+OH5HcVK5FXxUXBZ3IoZu3+A2Ds0
OP39vmp8u1lKBdsqR3Vk+GnLAiTsfFTQaxDQrs/nJhAGlnsrWPdrZhtejIRjIZN0
acl2Q64u9/AtRII7+frxXYIXYkMo4OE8f3UEhuhWH8uxlaMB4iyii1JwWKKmhy2i
+iQy9qRfWBCcNpMbJB6rd3yZLfjYlHJlInlP6gE+MBz7oVz4cMx9p6rXVRMQnZVT
z0lelBE9KbMs5insj2a6f2iUFfWrtFVZkTeJP3CHiU8p/KwhMIg5fLXHZPQD25gh
QgrJawcD8hGcWVZbziXfZKaP75llZ4kD0sa94V9hwXuLFO7mUF0LxjPHAGzvVvlY
9ybFWIPKNROJg3fXFsWmvuKM/mTk98ggFaqjXeQj+E7accq5PXMzXko/vd2/flIE
YkdpJPkVPmDLfCXgKemMBYUR3Mw24T4cQl3YQNdbE6xqUVv47VyU7u+/vLRRKcvD
Fey/fOPLyO+CSAZTmozQFzj/yXQX6fvUwMH+QjItuXudUdDAjE6h5A1IN6Q419M/
z2pf0QHY6yEbpwQHzREAk3oTfi5NIpYGiNXyZwiyB7yQeYE7wLSXntRA9kPhGukD
5wpWRlhPB68vALutdSyGcKDbCXSbYe5/7h4QchzG4DViGfiyrO6bqlhfl5flrHvI
ZMO9y2wgBub5T+CltV238IG/5eLqOnCMXDAHSiy9Ygpazq6RJxq+CvAUl3HAbD49
Y0RlfgRC9VuWv1XnyBBNLQ3UbFU2gBLK5z0dkPbpBIIGyoQs8qBByiIUuRRhJtGk
5SFyML2od8SK+Shfi61MM3OEDuA6joufxQZrJcKVllYT1Vx5jOfzTRJk78MZCAi6
KWTOhY0HinoHoDE6HYDkOtz7/6Gu/GiQL6bTDLW6jQK3GXnZNdK6b1QJPQ+VozO9
L9f79BM0Dd4JiRsZUHel51EJQpuaN1C9ONrSAGsTOj2ln78b+xNWnePCAJ3SD2ct
8tZEgupeTrSwKXtodxZDtkXo3JLIUAUk45ayVvIce2Vpm0IvzMJdNtR6DXxGsqS7
NK2euPC6hhz3bX9CYfq1rIDEU1/17ic+jQYmugvgZM+wa57SR2kalPhj4TzVq8I4
+fJQ/ljqRKtW1Q/aGvg2suMBNAMPmRIk8WLr4qFfxpTn+04qnSqgvyIQ25PuE7uc
bX9ueyah0h1jIoQ8+T4JQL6SME6T8orbpjUDVd5APsCBWIsVMmc5vnSzd1mvc6L1
HF10Hvjw2rCfVHyqbBTL4lhlcVeBRU2PVUIA9GeYQP9q0eOq0HofZBNiHpCgA69D
E/eVWBwz0jxce+W//v+zvqhYQt96axHVGZsZcGVLVPZ35fiHzAb3gsGrou7OYa8R
NhJryHrhd5pDdc00h0AD12taWWadj5ON5/mj66KQGVSp1n7rxWDAReq0whGtuUhM
J9Cw9ojL0By1vT5EV0vzth2FpdxXjUYV6tdqjVxdROsn0hTxEfPAaNpZxcx4YMSB
g/p4o37vmptp8R1M41dAd5Ly3ObJ5blph6KHnomA4mKpKxFg7KIABTtJWFiAoAOp
5cwW932wmwaXNmeXtmKhl2TQXHkdIkiGoWy1bv3JPdYzVxk01CsqVzHMRLbYKMaW
Bq2ihdlx0JR4gWBX884MIHXDdtBYLOIXHzjENPZZGMepWTUAarSqa3oGofgf1JIV
4XlMn/GWyUzhH598ozlO7Ez2DjE1rnxyi2VFPF/gpShJOXa7HMLzr++lmkE78UF2
A/VkAoycRj1bkrD488xoZVl1TBbAYZRQJcSuBL8cTblZ+J1P0bybJDvpytwBixsI
j9nIDRNVHNd/donsJSWtjuYGf/t02Usl+12eyIiTEPJjhnzRTWsiwMu/kIVT9fUW
b/PjaETHMAwW1TS+b7gfF4GKPpQC3U8gctV0O78iWgAXILFlRPn8iBr8My/NqMfV
9FKq0IdHJyS5N62tHnOYUjkszd9sZo608ls1n3JqP1y8E7fXLhDXKsnopanO1knC
bVDG301kxEsFRojK8hLq6bfsDvCUeSsxFq/XEzlTvAT1RcjjCx5lDERfelMlqUyc
74uXL0OBq/NOeoZciyrYkATGk5KwqzM5s030nfPtJZBszqPChWkltxYjeiFlhjFG
dgPfhIDimjj7fJlfwpQemfSxTS/3hJBaD+A2yWjDnnxihcS2U14resZVHIAW6pPP
aPjcBH4gvW3/XLxFBIO9U4i3cdLql5sXPhqCxzJcbWihgwEda/Hk/bZFx2pK8gO7
B0opd7CV4zufkDh58JhGzFxDDNArAuHaQl3bMJTbpRNfjEAQv1TVgrMKjXDhd56L
yvy+zpEKqNSApJmmEj7jyZv2supWAzAy5TAo4PHcRurAhO4GEvDlgal2nZn+G7Ks
yVmm5H8rm3kYtjq5jeZ1gyqkVQpSt9O7y9KRiMzbR9BwSLDNIE9uJUGlNYEuY5wc
JqUTWHVUb/pjspv+RadkmC4dPk6YUJfKge3Lii67qcdVFkFoBIm5dv9I/7Aq3vZo
43mSoSskbkWw6jrRG56ZNxGj2mg8V/Vam3TfMRv+iLZz37/NzVWYcfDAn3ehNM6m
iRe8n8Rs/tcL9AqQIN1BVCJwzXIKjkY/4ve/GJ4n8sXQUKzwgA7RnJKGQ4zTU2v9
2U9XC4jymHtFs+uSXnLJVrCA6H5i2HLgizoa/3LHhn+d/G3O3sU6vtMCH2d48rNb
cz2aGqYHfNQAKpSbyGszBgpx2e5Do74iDXHmcJySIsksMOwkuSwVuaRKgb/Zskgm
xlzPcSlC6LqtLgXgLrXvlLLOup6JtyaaLwAZ1STvUy6n9a9qEfQ1E8/v0EaIBNuy
wsmABnMSjwGUaRSHg5PiwTLs1sQs13slpKHXmEYpmyVk/pFf6DunDUaOGnxFxQmx
FdyPczmR8XLlQbmV2uua640i086oDBABHW75tADr/UG7Qj1sfrx7bx1tJPbFJmTB
kOxMP/F1WndFfhFluL1L9/5KvwLXxXX5jPzQszmpTjHpwRURUEnEPUev7jjM0l9v
6SufhJK1fReEelKtbmNBc/TMDtxN3zowBKPS1nm9nQ8l9YfttOTZhx6qSJP+4ajJ
92XBnc6AYzWihCE7t4FumfA5c0fgLjmDrDJqeC37J/Vgxz/xKK63pMhhrapVjgKb
vI3Ti/EtLTZn4VhjGdUVtCkAEm4fj0CvAZL0lF8wZVOD7Fyw7FJhkr0F/2643mXS
SncveOTMtS+eeFKwdQmKbXDGZfjAK+jHOgj8f2lRMOSAgksZcZiLivBJkm018yol
W0UXReV9vZmOkhGCxtU7DaB5Kqqu3Ptv9eGQvRL4G0U5qcUejU8oCo36GJKVPj3h
aJJbjdlCP7MIpB6UqjEBEFYVWUvpxwqkAiwCQ/kNCA+5Y8z3HmCBwDKc51rMK/5t
ypkW3UXDARG7FhJQvjoiDOBRIHNcEFP3swpPEjnJOaE/YXT+sLhzcdM4U2GbWu3d
jj/GxKrvOf0R9m+yiafuI3+IkbZOd0VisS9vg+3fV1NtihjTO8PhJVOVJoIfj9Ku
M7dhTRNb4kbe0eV7fZTs/CDtcYkceUICpLq0mwaswPVnnhwv76nXBBoOTAQt4E0q
XelHXij+Q0IWkAuRVgjs86jxMuSWTRikMxL5F++glqKuHgcQUJKnkCaaxuk52gGF
5tcjhtG3sw7w2lFzjI3jBImAWX/dJWmWk7n683KpLuIiognooJ+KYA7PnLzKngjY
mp8W/XECguXz3ZpS+wGLZ9WSUrPBNTfmh4pkI98kJWTS4hQzBfkcZgxliJJbtPJh
v6a/siUJwD5glNhzmiIKP7pYwUKN7J/Fb1/IADsD+cd5rD3IEDoAGATmRtb6GWcO
O2SB8RE6ONvzE2SePnDR/2KhD7yHfkMOqNMm5zvNHhb4VtYLpDVHpWvdeZkTZIeY
86futbKhF3TwhUeuS+VLswIl3txO+K2QInJVj1xOM83Hs7eBpgTqQQBKZswz0a6y
2L2QVjoyfLKJTUkraVj6rtZpOZVqtL6a0pwxd9sDbE6Jbe8SJzp0FeBbkhRDKXwn
V0QccDDcgJF0FA8pL2TsSdRQyQtwPlcRNElit+vkkDeurT+7KguELDE29OTzstpM
r6BHq/PQI5WLmQrLx0VXVSqA3ceI7m4QiCyGK6dOgPCKunqrbDAV3ttIjbpKCr7K
ryZ9LCM2SYLW/gUBfBSH1GElFModfYCuZxUhHNuQdSVuKDlnc7gOsrjy0cQ3zwru
bUjSQ6mOJWmgc5MA7ckCJrv7IlRbzukrtZK8uzuTCzukgzOK9q+4EBw9FmrKD7Bb
pDnGF9bNs5ZpBd1n6bs2+GwEj0L7UmgTFiGXWjyAdRUUHKJUxXbOTRsLoU5R45uZ
Pn1db5raA6p1SZdwpKDYZruF5JcY/jsTg1u2sayOEqRxcwjDifp+YHjF9dPAYdqk
WIsmSRn1mxRdal03PHszbAP452ydkGVYCbGuNt9izg/CpFcznaSpCIWK9d3vtvyt
otM43attgy5cMB8gQv/Q/42+W6L/dYOmcWs6yM0wxjmPgYyPed2AivwpNOnFTkjh
bSQ5oowQAEzf5XKzV1mpXHjkvTriOAgEQxD7FeKjaEk4L8ZUdiJAoWcOCHj9ThwD
o13ZBXT3qeSMc6OoRyz2LRJwho1PVhbZi3+C9eDjbXtk2DVBoLuqZe6RnZy0keKU
51UTJVhfxN+nnnWZjHL3uPzpDox6JiOGt39ZiAnFtTejpRu9A0G5VEO8zdz3NaIf
aCm6NrntH6zxBpxUyuoXvI64eFnt+Ro695u7IUJ6eq81FtwYK9rWKvwicem9hil+
oqsvy1ZwY9mkF2L+MCim6gl3xgH8OlnFvX5pNftQl96EX0EpvHriOqV8446AMS5p
iFJWLIEDvWXp+6v5sfZcYgrAdPDAHXDXHMrSgojIg6D6NYQCEIRnZp9E8Yq4POnL
ONMQly3zWvOORBYm3CfsWry2WVmHu13M9mY9q0B2TBiVNXY9Y7++xT46O41Y7q5b
5BUmYExNwZ2ZnhUNmW+6f2S0V87TEVvVXMo5G3JPoCqzRs733qJsvIAe13MPnEJX
Go9PRgnLcfBFIeDNlSwK0AZmvPtAl6buIkah7ST3SiLLoy4VNzWak+2f4HNBsuxl
n6cYsQlgUNa3tPpu0GuorvAU/FUzKkj5OGtuJ+5Utof8c+ssdJi8g/yMl98V9F7T
NaHWxb8eMCPV9dGDiYEiRjSEcZoWXK38NWUtZ1LrqZjWE1Nl8Pkw+gaNFa98vhi3
WoFyopFOMASIZjfnGt+I76im+XxAXAdtljBCADGQjaqOYRla34UAk0h+GDIhUdMY
yK6/+ADdhBEZKM3ikB/z9tkiqDGmD/K2xJiCi0tEyUEWPHJ2Uxd1+4w+5smmwqXQ
shPeTGr0aA+qlbiMA0CSg+S7odLhoDBh22ZyUoVWshOBpUCAUzzwe4jeEEUpFJ5G
wIFd35EQuREyP92UoDrIUe8pGqDX/MMWYwVOXSoEhhI+nB2dnUdbAQeejA+vfjfY
8shZfTj2tRULmV1AT43N+p51mNbr8f/sc6K97Jvmr6lAc2ix3RhTn6ho3X1+ahoE
VbtzJItTJe88+vjIDvoyd48+Yg6W98kBAxn4AZlcHIUGPN6NJl2P3aVNtnGgitwM
mhV3qk2ZVnzQncEuwMQN9F5nGpTahNSKpqua3w7sV+ATz42jLyHtURrsfdPqxs33
SO0Q87W1QpuYo+USMHVQ4xnOOWhNyt0EHeIQfbo2hVvxgeTSPAnPN041Q8hEYtmW
nc08QhYUvMGHk/B1heDim1ddaWoonOkFuCvY0EVKzKKy+lCLbrygn0Mj9oXPN7S2
IkdUbTlabImSLp3m15SxW6fyqE++JVPGR3IDTditAm+jqWZ5VHDN8iy1JJPE1C+1
wqPFk9ezDUVgWUqivnT6KlU5MNHP0jDpRQD29Z5yV3eWukW3X/JetRxHyITiO7y6
S1kAeA9Rt/qMtQWy6WPPVB7thtFE3z0d3FNJ9nHji5GQl2Wp8Su5BnL6bhg2OzXe
X/tJS45IGPdFwFbJz2a1+cj9xu8xZ1h9GUK7/lTEp/DAquvufsq2BqEBPJh3zhrt
lECsFGEr58q9/wqkn8uX4+PrS35qerB82Gvsu/RuyZp399AyUKCd+GEEZ+r+hKuh
ok+Jz/CiJmeqLmR064n/OiVV4sU937p1cf9+kKYbEDrZ2kTdFXSwh2J32gATr7l6
nBYjx0ayNXyGFdEFL9wSI6TZzpd6083UAc79nv64McZwXO8PQzvqEX+Q44xB5rZ0
OTQfGnQAa6W9V2+63UMejUb2n3P1KDfRGkdkuJSzi1sk+yJ6prUgSP226hsSwkDf
8O+JN34zo03ASdlDU7YlZCSPpVuYYWS7gjhfjGm3DP/SHDbpK0jNwyLMJkqW5F65
mwPufvt+cbmPi4tMK2cnv/PO1x0fHQpLnDSNoixxBXjduhabT7W10jdnNZduXvMF
zjPOcj/fCxd//YpaoXfGUOMCTv/SB7/lnXfVW4bS/pXzDEvmIZn7pp9oBSFrs60n
mVo5IjYa2cN4TgOlJqQgeXFZbNX/2Af8hudkLlhEpA5Osgc/WVpc/D3Rw+lZKEJn
xr6nmhInVUmvyMzfeEN4xUOH4R2oh8U1Qq0GdPOTcUmsjL5FnAu6I1USodin8R6h
XCj9RUV77J+UIemj3Qfqf1BOd66bhwTZ0G6hjuq8gLa4tYZwi26hUlonhx3GmMgk
OM6AVSl/mkILokmJ9cqZmFsNmGbbpXOpzcF1mQ/x7Pde6mlyyPZ9uWjrtQ2G0tDE
05KTikA9HoOHqnn/CHv+elF8JtnZyAOA7bUULbd9ry32JtklKYgRFbtyhZbAjP0w
69achLUCktxMhL4MbfJIYCrbQUnplr1Z36W826URGCUi6UF/MN60ld6OZ/LzmNNS
+LVxwbJG9nCCq80q+3Ou1WMYa/MGYDIelcCHBDMNpNvz4gpnvXm3pARMzh4qleln
9damzMl4I72iStkgm4lSzwthVgIQm+MxL53qD76vZJT4OT9U3rFhDzy3HTtXGbBg
H3vMmDxYJYsqXQ4OKVU247oSf45pM3QEQypCx2P3qBBILd9akZTFCMsrjZ7F5tBo
DgxLh3UCB0xfXKRxBBM5Q0Bx3pH7Mezy+pfF8nH0nvpSWHbddllo8+2fcoQXhEl3
41BGxfx9w1NOqXDat8rfv1oMoA1miJnWbqDjV5ZRnLUPnqChsX1COafngOrmIi+N
iJ8qOw2alidlWHxVIv+CITB/ixop/QfeasLRc5JVzfRZi0MuY4GDdyZrOqnM7KCK
XUBrXJ8CFUrA79Egf9A6YhMHdUpmKCVECSPfI/2uCHeNx1HzrVgKOfBoESH5V395
UJb5WrsPDKbku/Q6nJwxZCmrg5vKVKngbBvxLzVWEpB0hrpSl2HpGy/jt/ZsUr5t
pGQfL52Ogk5ZI+2ebOYd1QTnLBaYLs4ldbIwXSxJ4dPgj9e6gH15T8l39yZ5Pnk8
vCj7ZU/1Avbtfzef1gFQeCkWDvRLp3lHM3/HdEU4Yi6hHIXGKgugLElT2bCGPN7a
buJCWqM3JZveV3Ti/CwYGtl1vKLCLCIg7+gNcpt0r+VKFB1LN4atug2wkIMAgBse
xxPnm5sizVKeWi6dhQ+Ghn3PPB4X8AF3hajA2S68vS1domcVH0zKBSD9efWPHJDJ
VhVpfb6tLK1ONMU6a7aptAH7uUV2pC12LksNED7jGiVx9XZOhW0+d22h/ivZQc2i
asdk2Ru0HICBpYB+aTDyPMFWjadxEifuhfr9q/xsg7uST2WSeaEeXo615JfDk/+7
/EGuD8rZYsKa+o7TpCRWO1Xa76qro2QDTCX855Q0iOdxOMDGXAh3mhF/VyHU0Hfy
qUYBC/AbezCcF6pk4WbRgKlJ1+6vn1IvejWCOXCSQlfvWJGUaxUeMrDOSvHKG0YS
yHz4HEDn1lJs/Insd2NT4g+WxDsbQ/CJ0uqDo0zQtUXQia+DeVYZaNtMO9i+lw01
LisA1/sI7CcTo9YoI3p+4CVa7JuyUc+K1B3GQ8q/K8JHbLwJ0Jzfny5uRfc4L5Ff
PCk37X4o8X3u0yCGxP/xWuEmn9VZBH8icxe+nawAy13QvzI/v53qzKNDrNArs1ZN
9IY14G07LFvhmn3zuIG00hwFKU3/hiKNAWUEJdXDrHSyYOnD5DLyLxncjzclvNaK
oeIb4UWMDgBZ0WtuI332n4X4fr75Jwo235R0XPaIcldBHnZxSVowDphaJRIWWE1Z
6RrMCiVP14ZL+bkjEAcK2HZSD//1AF2w7aA7t044jXujXBmf1VlkvJK9BhzXeuL8
pNoh47fBmDbUGuYOL04woSpYYGXekyOd2FLTbbfE5U/pAKPNj0+EbTXfJTaGxtxu
8bn0C7Xva65qO0Uk1e8qxtB2HCyIoRzGA9o4yXnkp3j7Z/j1FU9bRu9cmkzFqCr1
fzmCuHqxL+jcquYlVbLxi7/FK5EVWlCq05PPkLjDZIntBSyvBA5Ky5S7GOIUg1Dm
VXW7aFtQDVlw7tWbq/SY4X/pzy5LJouqpBPNbl0aiytGWt/U4eFwQfcg9jrCB8+I
9TjwNb1Wx8M03aE2gs7muCW/NmrvGy9okdh0KTGUjUGM7t8lcuGKSILhPungI9DI
r8zm97kBA1DBgH22+rUGGbteHGgYvGDV1O/OreyFHgvFdD8sEhjJxkI6FsKl1Aqe
wd65XvtNu/UXbNk4m8kuJgPa4h3X8Wmyu/qdvIvCcW0KoPvwJ3DYEpjzPqYTGA+F
7bdHsSZJAbq9Q1ShWao44TNNukO3Dc0E0TKkAYqHI/hookGoI/LrqdbqUflmXChj
eQfpFeWCufpyBkd41XXBfbg9UCpNkGkrvSwW77K1qKu67WRkRsU1t+d9qSHxyVfT
OYFDOJUcaj9erpgJ5DGWNYX5Jj2RsMsibGD0SvB1R0vaBMyqbfpFS2D4l3uP7LPi
IyRa1romlp1CeJgamvh9Po6yCBZ/qeccNOz9Fd5ztZXULg5gIma1eN0lFEi+sTRh
RMJXK2Hrsst4tkbL6ja+06j+Q5eYxL2NQgwbNKfXskwHHYMABbhXvBoJDaG4QMoQ
YsaGGUXRu87J4irTa5cVRD9/HGD3QwdLxdnaTEHPXA0gpdKJja8I53RhVijEwjZG
h/ySa+tbSouk4WWn4RwIi0KFB47gl5W84Cs4jqlNijAM+nzfSEbXdJGpgCf72Zdy
cgRKyNk7Kw/N/NA5lMsfAZXI3WvIrnb/kjebV2Hofjenj3qrwlwNmpSEAPYuQR08
DGW8Y9HC5qfTUE+qytV2kzQL+fcASeHwXApwAHLYtUqldSB9hfEEK/yoAF3wkZIb
i1HCkKLN0vIlCMKGi0bRly/h9q39hRloZ6BHoxbh/Zuiubj1TJh/onFOzQyrClAM
S4AOT5oN60u9/phXuhM5RObJ+jZDtL7XNoF4B+3nDeBZodXMrvTDxwGwZGswKacT
DMOSEAoekauliDTrMxM3Kgl06BUKjVlHsRCUpnI1yJ44KzpZiwU6GHj3jIBkBAZ0
RXDOz7lIIdqJHpPmWEAMdhSItTuenovQRwODNugYqH1Y9jjJouoo2QMJ1NonftVz
7GAEtxkI/GMrlutpScu70nJV6bN1KVXz+HMpGWU0XG9YkVXV4ovcBBqJZx8Kl+FK
Kop1PX3pm4A4r43T8hmM8W8AKcZ1FHvhaV4k9URWsLQViuc3CTj6SR0MNlFkG4ir
5e0pr8FU2UYEg/ReV5bi8WPHiny8aEVR+A4QjaQnsf15bFxcZThIRSV95ebkkCX5
5uAwqpr2sVd4MVp6KKYE3suqvn+0s5ZPN1ThKK6UwN6hJlFZl8SUbCjrpIkdgkqp
NrlKo/JDKC7mDgcmWcCBtRKEeojATwjO6jnHuR/HTfzTeUSA+P3JySmnjR+6PfCA
arSwnbJ7/fSxphTilAFi7blJHsS466dvpWWuJfeih9g1nNuz1URpBwcsmq6gAJWJ
wwfhHttPeJDZn738eH2pIihWfKRdYkzCdxDPX+U0TWgXF99G8bWZGb8gM6krWUjc
7tJiLFX0s7Y5u6V0ath9CY6pSfVU2mvF+udeDBO/2y+FI5ZJ7U3AB6MrfdETOf9/
S4ajjs/9IGiSkGmeP1YN7damJogOqW7mQNwS9MiIPFn8mGCSFF6u5xV3/iyEY9mo
a7X+tlvtkNZ7ARtKqjYAsHmhbpcK6jFoDCx9b5o9ZUhX6fmXe7/C+R8g26L4rk1u
PdFZB0RXgczsq36cdQYcEuLePP+zATOBmXfL1yLvfhvzM58fz53LNBGmQVec0yDF
cAYv6hzj3HlitR1TiVw6JBvv0R7svA4qFg8CQbPOnszc5MjYJe2ggFJxvWWVrmYo
YRwvpPTmo810/japfppGILyMugEOBK4iCUCNKjuYBzgQpSe5ehAWBtGPWfLF8X/U
EbA9YEXtQDVaEt6k79nQ7I4J3ZvrgcE9SfBz9jVBuXd/L1XuFbweJVA9Pc6SYxft
7GXWdKYaEF7k7Kma2n00uw/J1Mam4e/uWecVthz3I0xLgSpjHnD/QwREvVAlOmw/
wF97HgQbvi6Mbfs5c8GYXAn9jc/PM+GAqDNfIvJbVXShG5Hepx5mkkuMvilb6RHV
+k5vDzbgjxEMnWhlzQVxjwPQCSV3Ji5Magt+AHi+WccHqOLgzpu+X5npQsDatQhD
FytJhjyQO6KutrjPwq/reXuP7eNavHTmB9yHN6ANMndf3SZEEu9uvz5sh86reLhE
14O8BMS8XWesYnBzdrkSi4h927J4coZB8RLwZkhChXb8LA3u6SMS5cPyf+cNgtVA
QXTMpO+LWi++HimMC7wDltW6advimDB+vDyl8AcCE0tAut5RGffj7MeV6lVVyj1Q
7a5Z5EwN3GxS/jCHPO0W6FTkyrTDSc3inQc5OYMBN6O2QRUkEYLxOw8SsFjxtSDe
jWQstRCRfgjH6kmqT3RbHq5FdjimjijeuO4OtgQQ2Kh6UFCYjUz9ACpvS+QkzIf4
SwoT6FxFjUsJVJ3AyXSsIACUfrHSPtkPraCMYg+eNULJu8N+T/tP9UUuVcMuzXYk
fGfbeA4FHfqbxoXNw/H7rSN+NCP5AQctcUgTJU91LU1qrQQdLFIArQoF/r8cfDzE
k4GB7Aai1KUbyfSFmtqwOu84lEio2bPiFw2L1KyfoIh6RNlwCuIdTydqEgs5pQ+5
BfDzFX9G6dIx9FGy0Sf2RMj6ps5HcTCBRgWq6ymj8reGuWP4E4I2F3e4WP1XaHMN
e4aE+Rs8+qoO2gYrAKsFfSXpma6dj+UmQ4uVdCrWuUjgKWtakt7w2jBJ+xFoHT6s
lHqyMa2IEY+VsN6spte2J0LKWlEPnYe+ivhQdr7d/8gYwC4bCcvo9Uhe53wCtJGg
JAFVPvigcR29GYYHgf8y/y6EN8jFLC5CAXDv5+5owlmTLn8dSzwvulS8VYtGClyJ
IfL9/JJSC4vA/5bwu7qxm6ojgjVh5VduOLQu3x+7t5r9hNTrjoDBaXuabS8MCaxR
/3e3BWH8I8JjsKMPbkV8GzEInLdErr6IUh56xTAHhtnkRz6OjeSoKkLIXNabnwpz
287Dhp95VJ4memMm9VF9XdR3ZAeC2kL7R7qlLSbR4vBv1q9dtm9+d9yVgKcYF58Z
3VSlxNubx0QjOjUFkza/o3A62XChsgR/Rv1mHIzfjMMv4J1Kw1lc26pSsEmiBcjg
z9EMERt8KKep3Rn7RPBb89BR7zJs/So3st3PBwJkW+vhoiXBs5POiwpZzWE2sJ4+
BapjdyFo6Q9vu1vc+PczMwV7ZVnhsvjOmRICnkI1HM7IfVsioeUQJdiaDsYAodQ3
4Axv0Ct8+OHUohlxm7qWcavoK9Z86iA9IpPuZSP3Ybjbj3mpOfUaUMDjozqClyw9
bpQhm7glwdXzf3hwgO4G+jycYJmcM6DeG5uyEv4MVN22+m5XMNiuDS3UeHQE6ez5
LgiNUURjLMUi8E89WBb3d/yU92JBa2NnczzDeRefwrZy94hb9uS5ZM/SJPKYkvqC
A3X8oE7ohNLZLuZAwcXNNCuLkXa3S9Cyp1meN6QX94O/GDEu52OMpBZ/c7fEdXMg
u1E8Kjx0j2uATaAMWOxepo71sDZtVTHvWbT7oCPGu1eq3m6rYGEyushTezJEWgRU
KbzujJdLfzUmyeILKm/Kwd1YJZySifkAvutzJR7rH0VP+1hXMu3kh5zyTjLLWF8C
QlI1TU5SzizIvYXAHm4IbcdftOoXmZTTgmeXewBwen3hwJHm61EtBDU9lPTkhJsa
hsldMcvNJwCCyxDlatSwDapiZ9eiEpRmcOjtRbNxDMbHaCNDbdeBONkRiF+J2sHY
vOFIXf6p/+IoIOfM9N5yidGyPhL6tMFJ5Ar52h/cA4TBuqi1coK/arcBc2msWddM
47PL37QLDmm0mMsA8baks9G5a3rGMYWUutbnqK47OsqWMCCKJ8dCVftCErJ4o0Na
w9zfzDuiOfEliQlCbux9RosNTF4zgOxv+/S4vx3vhvNgbStHjEoFfww4OWDZW+kY
1LP0o6qwAcXVbmezKXz1qWH7kqNaz5ujvMtHlB51s7cu4ZhF8uRQoeoa3zcX9I8R
3aEhceSAm1FXmGDVQSrufNHaOe5UTdYKJGtGh3p9AGDsGvNGK1Y34SVTEAPfec3z
TdicTHichKC/GBqH2tquAMVeaIrrKC6LhLpX7ZwIPf/UCj3JfQEcxyGY1Cij9OVz
cCr4yRX8eeXC2aoLCbiLXGcCw6eciiBwlZR3K6C/xbc5VR2re5lnU6tgypEVNWNy
B1RygZo6xec1l+aXGY109LvSZUQg0lh+HSmm2Kgs7stuTpFTKnLRaNmlT0Et6bPR
suAaDAlwxgXjqho7Li3vYGboxgd1atgq7hHpWA0UushbD57oscdeVRJZSa4DhnVa
x/p0If+jdSUqGoa34PLj7lBxuP66Hbn/LX17CZ2FsNMCRcR0dckPnP1LsbO2Ifst
BTvH9DGQ2ocSwVfu8S/68O8+olAUy2koGbYNgWIJiWDXcSPU2NiKCRg+fldx9Jsq
Bl6nWl1SGJkRn1W3SPwcCKXdN5gOM4eYrS3kNFHmhh7F6TArDFZ95e3EOd1iON0f
sbHsW/lowp7YDFozrDxGA3DYRibbgyOdeCm1TG2ts9p38ekuqeAoW/61s7qP5KMy
+N9i72IYgE15evGofFQGbDwFa6uWZYAPIawSD8ZmEI4yWJPI7eLC9hAOI3jwjiVY
T6g/5mQlGSw3deU5CAwqfugK66DNgMdP/Y+t/3QiVdjb6yM3F3XY5zUJEatx7kWj
YyLuFlgkOt+1sD2G12L0StyahnnFWV5h/wf0R7aipYYlxVRPxnUlwta03Ag1CLRP
pZQnjxM2giVERwkP3uh8TMOpyJHRhvYbngiWONdwDufHT0bQ0QtGwtadZxrtL7JJ
HRfChAwQMTfw4yvuv8fdApU2NvTLq/gAYb15ibh6S/o3I5LAFljYgjRTiaQy8Yuy
Sl9puVUSoG6NxSNlYbq62BS3lPeIzTDVNl2Ec0dfOvsEPwGKvm0CU9w6v17hUS+1
9OjooQZoy49KQX4aG5SECT5ObRAoVdV5R73eFN/FkSW9UGmahnCy6BQ5OXxdGwGv
RuOe+v5vf+Nlhte1ovr/PYQAoAxA3ovMcYcH7j/E5JegFUePAfW+ewNeiYiojiqH
A3aj5hrhJjMOIXsK0yohavdknZVwLVQo/7bD/t40mx8qEVV1yvRzGGih/KIUeE9+
cRZXObOrZ7UfFhzsCtJ124A+LJ3jZvyi4CI7bDcb1BOGzH4+2srGMuEy+WBOn5WN
LrUcqgBrrlryHmb2Shroe2IVEfMrX4POrM1SYZDkxaRC39UMSm4SQLzYTWrHrr/+
rreJZayW9/uchzQX3D9Vlm5epQl9cH/5EJyh+wBSJpWtU/cZDVPK7i/AFw/W1y5/
8fbbFRoMUl6tuI+/s+DBQ7zWOgVkXLX0U8I/VDwV/Lgb/L24uRFZCIc9JW2oMEVC
1O3MyFeDCBy4MDDvyfpxpKRHW9ZjcE4ev3x7pOZhY88Xmw+vADcqq5cVLu2oaXXl
WxkknlWnp98XudemDX6MAVwZ7NrkLfVV4hoVtBpajKj/iYXKTPzCQUvwH4HSX3+C
aeDPkI5GRchathQlBkR+FsQduKkp+i/gDNImNV5BepEsi3I2XO9YB6x6L4ufhBwK
scFDkq6T3oEzRwmmdbW7tWgMSVZq4GI89QFxyr7zgllgz4wVH8WBmZYyMycGBu2y
tRFWOQM8TyytUWttZ0AEN2MsmsaigUTTuPM3+EEgUVE9ZUBxNROqds3JKlJHgEtF
XZUVuyOWSfhJUPXTX3A2907IGZ+A5HkvjYnvFbT0a32KTLKEsFrDX8rrbQm3PwCv
eYg+RAxKM6Pch/X/2JA+kWQxAo33yhDVvm/IQxGGlutu/CYyCYf8g2GSk4xj5Qni
5qbf0Mv9x563CmXPIqAC4CeR93JQzAAPILgHQjtJumxV+VIEggGU7D/T/DZd8jqz
iEcacKhXQq/WVoFbA23QeV1ZRu24zAG4wpaiZ3hLEaTftWa2Lo1LGDVj80zMV+5i
bbwvOijGzzyvXfCB+S2Ez3SDcfoyUPBWAsHrTvLubODzKor91YZVPGHCw2hWH0sH
XGHI9t63NYxE7+kMz+TCKOmwTkJj+p9N2gibpex40AWGmoloocrwkIOykuNTcXPs
wNVjEZ3BAFu5TYIwwGV+lUeaPg2dR/TCJmlQHa0gx1Q7xXoxZBep6/b515d6RuR9
+jEgsn5PzqqzUCoyW+VmRHZgqdyvZoqd0VadSHPNya18dkhdRUxmMLeHWIUicluY
dkg03l3/omQk2O5xxhRhEwUU6YHg+Fmr+geL8hMSDE0Wfs+VpRtJv3UM+/k8vHRn
TZYpWdCn50ufd0JUwxh9NfEv34urxSwdQpsJ8+W0EvYJ9qfvO7kClp4syZA6d5Hc
kLmKlbtMTM7MXBVTYMltuvAyt+Z6T5Ibq5Esb/CCfHE7TTR/mM0NnUQPfcHm4EMp
oqs/DuDwEFdNiIvzQlzT8JGMggBrT7/N37H5Ct/1imr5+MiRwdx7WyMPa88KgyZC
DBqQNIBxUuQvUw3ifhchTRxJ7loS4mb6y/FIADQvb6XM+MgBo0V+t29bUlTItNC3
LOcpIr9BeBdp+rwIhoObTatKK2UHsHkdggXiN4M34FkGV+pQrPL0FKl6mIFim2Kk
ggy3oeK51uBvpOsBZaYU25LNg/InlGufmHYB14w2Her7S6s3aF5jXzD9uyg4+z3C
ZeB9EI48KHyDg2sFkeGyj2EsVPCXj+l553mwBe7E7tJl/Cg/3kEa6DckodtCnqgJ
fOyhQjjQDlnxXgC+pD8V5HPjRIGCba7dQIYGOg7zVhAqhPvWQalENITm7Y46KpfP
TEMgV0DwhYfGEKXj/kUZczfYyLkjNoDkOfhdfWQ5AuOydBbQeTUamLCkVhYo7EvT
dHFbXEZGg2r06I5kj09btrZqyvjTsco6qjNXBrQPMR6QTeZPRx6QEnPXGv83LHJw
p1UepYWXcB9ZCX3OUKpT47Mj4bNIDa2SxiA2QMo0pybm4ceH6TtnCiQTVZAtuzft
+ltgR1JOiiLt1mxa281rXwuSDW0tbdrFC3eIoUQllsfWSa6H1IOjs+I9WMpje+9G
Hr8ptDz/XzZMNs18RMjoENgcy2xWQL5eUtck2/KDvqaQXZp9g3smWTKNb7DDHxDG
1QvFFQVjyvqbgBLrHb3jWGNLjhZDS4JXEJy4FpY8DaLnB+ZoRLRfkHR/2PVeOxVd
zi8pFv5BFvEQbPuCgmCF7pg53KmzmoXWbaaR5HAwVfivgBbxPxYfYHQMx9tFEmCG
BOFO8EU2O3T/H++gG2tW+0qCfJph3vCYlnN8U/DqjQ1+QlTN2FqbLK5olrzLqdov
wFnLuRcWm7pUpzBi4gInImktGYfL7AYMctsJ3YcpMzRy2HtQ1kuHl0gePYguiX95
azbGyVkPUx3qW0UnY/txGMJ2NhFTcugOcdTAVlToLGp5AiCvUDyQNpqauMOzZ0+i
/a6Ke8W4WvX7lf6clgH4mlTwIx9v2Jp1Mmtkv7HvoLAWeKJ1J3DPgXVV5OMogY1T
MFCBulJUagJHtzeRfX6bkC+r6tnptsqhiOTo3Nil0H+CYmYrKJTWXmSiUoC//KNY
vYzjGsZtt/eqK+pWIrnEu7sFvwovkdXs76vf80AohEWE1j330UtRL86Qof1esEyW
Pg43mnCGVh0bwFWna57a6NT96TBcB6Xro/wTNjaz1s3EnxetKAe+LNW+N60L8p24
G6UcrPOSbu9bOIPQXT/NX6ZmmMwVpeurjDBBCcRm/oVECPFoxEY2lxH96SyLd2GK
817kI3wpuLajlhmIOiUqs5xwunmfHugEzS/C/4kyaHdxynDS9elt5K2TF312Ni/a
BQQun3dMpwnWXKsmN0mpBtrnJgn/AaTmON107eUycPiuNnl3xoLIIIPV2Rh6S/dY
xWxJHFap1K0lEJQKAcb0tsZrgEfSRSEqV/4XvtG1d0EVwzrKFpvAnpv2FDebEHrF
8fhystIkOhpd6ujY1ZpWgBm0jCdeeGyKLBIwHkzTvtRi8MpnUL5nkuoLMNdM8BuX
p+hC+HF+hWJWuKmoqywzTVwdLe/5ecPdEZo7iw+3tGkgc8CzmKFoWwkger8S9iaY
+FqfaNiReQvMldk6Qj/PsODkVloKx23xj8vrFq3CzPYY+y0CZ1DpLb3rzkvhUhcA
+GJjy44yBIC5P+JJvkRKWpdDgnpgEZ6XKXsWCfdn/YiLCeensBZt9Mck6C68/AFR
DQ5Lo6PXWUR95Qy+Hdsg+aFa8V6tRds0E9GHEJ3O4I3o0TlOU7pZyqMV6QnRToaA
3x7lzT9StBk/zZSn90K4JFwqtrvPBbVTEtSzXeGJ7VzWQYWyDDSu28Gp4ckenPGf
NRdIH64DhT+xw8oYp4wTbrc/D27qkfPa/wHZ7LF0PZgYOuuc/YaGjrLdZf+g0oni
fKbVnncEXcOM80G0xkXl57JlOHG22llNgaUe+U9e2kr/RAAQ1PaI997MO6i1VwSN
k0H+LDwYa4IPMjyS0KQ5rRJcbZMNAZxZLyWym+tJZnmzl1F1M6BhGrRPEdUG9oAS
fuL90sYS5rjB8ZsUV6gHOSdnTpuU2wqgwowOugMJgHHAE+jCbNw8Pz/6oh67Pf2w
w4TV81A86kAttOecLhtMocQOAwz9a5D6Y9XIkTv0XRPAl8+vdsHZPt/BlpBS5Mi+
AxvsJw8JVH7cmbtdUHz7U5IV8/m/1YhwVZ8GfZoxI4Ozpi1X2zwqx/W59/7Zhxz/
zMGLbcz+F77dDitXxw14qtb+TSdKWyTh2IrUm19ghiAoNwARbGY2KI5NwfGdgUEC
GaodPM3DxLa9k1FmXZ95qr/sJ03zfFp5NpmU3Idrv0MabeGB+OEkJReVQvEkG9HJ
CV8kV0H7oWplt9n6HOfChuUC91/fElZnJaAHQa1zKsJ8roHbql0t5HggTQSGHvC7
LWuLC0kQS44+cNQpCet0jAafVIc9e8eepJw4RdjAYJ6/i6OfKTixEPMYvLDzmrRg
HRLONAH7pmYFjoZHSIkY5fA0qYcsZ9MR1ufyHrwl0j828RrAt8UCbacXUutC++Wt
viuRuNHMYhoJW97npfMUWynBzAWv2MLbUj58aynWPsmuHUimoF6k3VDLKGsSAbJA
QYVXbRksJxEd9YyB6/D+XTBnfRbkdehjCENf8n5+Pr4pb+55+zT7kwByMZQLPD3Q
3WvSX0ITPPEaH08pxT5ypVjwou+GwBzfuTP9Nwwxe9H7XZGzu0PiG+vNtbkDtFn/
8ghGh2SGt5+074HbmbkiDjFmezPx03jr8JNq2tPJtHGO8TyOJjF4mQGo0m+bsdQI
F+t8cqBkFNqO3m9V+ofV0GC7WPnwiPrEDALh5pblddNn7ojIbYLXtzskZQ+cWaE2
FnILYvwQri6v0DtIjosVneedcNqrIzPx1Ygf4gpwZRQ10IzSMBdxTDs5N43Jtxdy
QR7XX91zQH6Wpih7a9bJWwz4BA/uxSd5Bnlz/ZVoZ4ibKtapiRFGCTPwIu/xRZpr
xImF9RjF7ATv2p5zQSTd/SE233hLv8tfNMordf/EEmM1P3esB3eE47oMuJf5ZKfT
gLpGXadVDoBJUSZLeT0Z1rhgMZeTA5alwlcq1Z5oNAeiUPRmlEc0kq4E1VYC7wyj
wLE1lD2L5l5PQ5L+z6TBy03vTnDxuop0BZTIThLCgZtHzDJsKYSm1qbOLEqplyVc
cPs5RZyYeguA83h8iqD6YnIEnzUHUkpG24IGbYIpgfhdHeeN3OzbdBA+Uy2xRjRn
aD/HASzvjYJcRoKA0Bs1V3+INZCwuKnpa2hlun6T902obpplSnFwKq4TSTFNeOPH
hRAUtMWu7bLIyphI3ZkLZncT0hCpTaqFHetpVOD/ns/yM+HaaUzNFqwzn2xn05YL
x3xBkkYCWlR5hxtApgIIXd9WxpQt8II8+EgixvVlS31/5qy/GeJK7yCdTkdUQu77
ic36X8lQEjTvngEHgv0xc6/NUtwxnwJ4zJ7zevUMQ/52ITjVssOcDTEBXI+FP+rj
qJIT1vgnrzABfvB/pMLcMzRdLlGalYbv5A3B542mhIzOu8RNG1IErFT2EUmY+azL
zOkpUmBW9CETFtEtiEUq0/35vNzB44lKtIqqExu3l9B96K0pix3W4N5f2RhrOgNS
EMGHROKqMelMKEjy/I0wG3C97r6uMcjSPKP+2/aL0VvY1zto1j/2nFG2Z6a5lNVD
DWmSlXnFxQprWqNcoxA7tdZNcHQlKX1UPCAldgNy9/M+PBhSTsB/03LTt8gklDdu
oNTnvQN6LaH9yr4EAENtSyn+sy73RSEYSBJKm6Iu/R6M9ElzNUdvc6A+kAVIG4X1
hIkujvqvbozYm4WCia8shhq2wwLlMj5KqItikxGuZHvcNikLX4nv91YUWFuHdxTf
et6JRwxlBRxKyJHA6nvBmw5B5d2WWPXS7IB1FvtFLo3j87rvuCB1XTz9cR/DkkRd
NeBmfFMoDoJMdlXjMWi5z+80TPZpwY1zWx05oGgfgLwYRnBreYb+KFznvX1BxL3J
D5y3pPD/0G0YdF5kDSUGFmYU7Gu8TQUMLeSIP/oaetQpDVbwtUg/r6GzcBouyASl
cvFmpzGnL2U4+MEJo7cuhPUKE+cszzqaSA8UbMc/BlyERAi+cxIXKmk/WVAgb6Rd
vvIRvTLxKVzoetEYDotJqePVS1zMc1fRPmHlKN+WS2q4iHeDQY4LpyMdEFdUhzuh
DMPpZPEq9hyMP1aPf/LMMwtGL13XKz/DFvi8evOp9x+kWfZnrak6ClRR/YMCawtv
zezVCzUgR4jyB6qcMmKnpQKZM16nyB9oLdUpMWOcyIU34dOfsSUcbOgcoZxlKUaj
Fv9q2mdDPBUNIF91hcDmotEfwYcSeKDZkdrSWYwexq5PxCHMJh3m+9L5kHmozWWk
gz9iMEOL0/Hd7R8VZJUB1QObexl51CPsuifHq0iDcr6V4IMMAfYQTa0N9PBIHCfU
OLON54WWcEp/G2SlmS1booy/pOW6VdY4zSYPCzcWetMIalpVelsPFLMqdAVxDDFm
7JJnn8s36FhyRfZw3LX3J1O4RvpXHIJHPZJwbvIb0mnn5KHyGN7OqmcLYmT55ZvI
CQtvXYGfylp/rNIPexvNEjcdenUQ5a9qccZHVZ4Rb2vfCGqWsLcsjY2f36IHZE8U
EZqZk9D+7DPg6CR3yV/p5Rw0NfEObTSK5h1CL39aR8+F6RTlRtGJ4Ha1bKxn22QV
RtU4YleecBV9HUbtJg9EHg6PHJkIrU3wS/pZkRR3iQ5fZxEfvA/LO6iXsSV8+VpW
GD70JMGyGkyK7w+rQe04M6G49bIWCB3X0bFY1NJufV/8zgD1lk6jOkB9UTVeOhCX
jkcOAu88qqXfFBxm+8L3cVfvPQMq4FtieT1ZBrEk5qkgriQqrcfWB7tg88S/887t
DfChEG2F+qpEliS5TKTkDiixmRdikxzCcz9ReWs4nfte8RtxyqhNCAapCQW0JqUZ
Ty/Lyx5dd+9nn5btVsewLtbUxUyK/P3ehaGqKWXnJorvbdv2QkICHmzK/0le6LLb
NN9Cjm7inSxyTaNkglwHAqsdtsQn/2j40z9Rau7gWXvD1HES7VpC7FQ+RmAADBDJ
/tyUZX4tspYZQdU8SQu9zsVtk80rc9kFqPbkUhxK7ETlsZNfyQ/9+y7z0b8dHkG/
TEIE33OLcbjx19KW29scmnfKiDKakfA3wclzL6R8zufV7TJMYiX2kDFkYsSweV+r
Ei/oQHLvFYAKYp71mWjL6v6sQiwkr9Aw9rkWOkVQ42Wcm6vEs1+cB0OW8eGveq2n
bRCCg6o5xAFR8mP+mDX6O2IjcNVJYugKIs8NZ9HzyR3ZyKMkKN0eFKII6HDa9czN
ZbQslZdBf9bsGTCWsP3JYFv0a0FkMkPIgQOkB7Q2AgoSQlvptVmI6wFxWEmfpOHe
Z84oQvn75RFWf/t3T64pJXaqgBXJimLZDo3nV3FwNJg98yMnIuRMqqrYth0QerPB
IfADf62cikp0Bdon875QWlqao2Z4P0Aypc78GW3/PAeEK8/Oqri0vOcF+nQdrl/b
4klEC95lO7239z0LsqhnEUsvTNBROF8HLlc+jnhyfr3THJfzMdASJai/OT9/CVlV
pwh+QUuOXzHuUaEEz8EMv9yquVYyZiaAVs08gTtZURqnEiM8rI4EQ0VS0o7RlrQJ
B8P35drx3y4NJ9tHFe4rF+IVUSvT4FZvC7zkV7hSRO55kcUNrGxuSOZKe4r/OM/5
PibZXAqWcile5/CQwWtxKFbfPZ+02sjQ0dJpwZSYW4oRIChAhGtnUVlg7HrRC1T2
iRKawQWwvy491as9R3WQERuuv6fVsAHdZT+TllUFUdvoYaiALms0XnH3ov1F0DVe
YFCbQPxm5trnvaxhY9m0iONTwokNQYhS0nYFDjk30aluv0mYFLA0gbzR32D3A4kz
iq2k6BASfEl1SyQxv0FLJ/uxoCTuqOgqOBKDce5gouVnlv9hs2HJ3xgI4cwC2tU9
F6eQ+/NQsNTyH8sbkUjgWFQMgWqMOe+C3vHdD9d6W1OMgXSvGZuSDGx+Bbm4cisp
R0ZfNxaMDXzI/cLEgy3m8gU/BetzevUEIVBHyJHZZTXKuOBjxUIhmzPURLkmdg26
+egMtJ7SYQ96ZRko36EPe4GIQDbr2PyT0tk36M0TZO6q4dV2z4ykQmE1xz+XFaVs
jGXDKTW/1tNosdXrnFstuMjskCahbxMB/IsBr/8K5itdbjyxVEPr9BSk8rUnh8Hh
kc+Ew6LtB9BQPYMiFbIuYefz11oeq6BwOE7nuyVhTu6Vvj/NzyXE/FZwPddSHBbX
b/5nN8vwmw8jAfrP3ybGf9BvhHfmgd8SKYd8qCjCsrMkooSmaNg1Wta8yAWVDgzO
FDj6EeDQMnFzko8f29b7HLqm8NJ2soZJdfZzQhE2QwRr0RBLU7O3mELKAjhN8dLI
8IL+7E/xDSsYgglKKi9fqpkk1jKN5E7nqgDQU2/wCQp26IdF6TAXd7C1jryIUYOX
JwRMckP73xwWEPhS4YfPwXwIB3Qeca2z9eUF6f4klE/nA7NTGWrTcCljtWFmKa60
Ejre7lrdaFO0KqSoTUbqqLkfV7OZjQ+I70WJdxixyC08gJoxdEFi5oYyjcAqqDoX
ZiRh1PerHjra+267swCa2UXhJQdnw3T6Si/la3pbl/Tj2OK3MUAlNlgIY0Ar62qm
xwnONeGL4Ai3Xt8spdll1w4nWEwQpBN9YNOc0chT0ZU3PEVxd6QoFUJ6lXVV8soR
2CLrRj/zmZl5Lu/gjCBd7kdx7RqDcR1uXRu+1g/HFMk/J/6gUejsmysKJemixbq1
0EvMM1JNbusPOZV34a0SVrRqbvumWOBHw5X5zOHOWb8MhgSVSHym+T2HuCbmpSKv
MyO56dVEBpyclL2VPXmPtgPIJsWq4o1IEoYa4BFJsd/VWIdzhr3e4d4GZUbyA4sX
umMctQevu9H7/zP4LS0xtK5JS8irbjXzQeCK7fjCo1KrTMO69XIqSe8dJi7VgTDl
5UxjPiR6QrD6aVmsmQ/VdqW99+sqA+K+f0bdMPrQB8//iN2gVG5S6CG/7REvo1eX
bLZdYrIc7FIhQfaEPlGrjS/udqaE3sp9XILoUrXTvSVZhNIbM5QX97oeCvZE5YYV
JSRJPMTYf0AKxzoNcjPUTj8pbEDe/NXEadRgr09VD4otBqR/y2P1eSsjGnWP+RLD
fGLIXWro7qH6ajSC/QWVD6+GlusKJeYXJtQuB1F+bipYCFV9V+VHLj8az3OwSCEr
DDuteieNREY6Jl72cP7U2zUMxXWxH/JJajY/zhzpB5slXvMimIkcVnfJb51bcMrF
fAP/q8udeASVUlUcmQFNUMtSiMJQllHneD53AdA4zOQyQ+PcgbCfJ7oXcbpGr/jI
68vri5ELwdDTZs6gW2XdDIMenak+Yua6kHVyqojIqNkBf2mW4oaUUuHWQOqtuohT
dbsO2hzrXVTP7bEhKT8XEIXDwl45h9BTKX+nGn4H/NSYf0cLbeoMIWZpQMBQHZ99
NAY9KBTdLF2RnZJTPdi2b+xvCO+lbVSeT6sFqZlLZMYiqdSRk9EuFbc393inN7VZ
2BqX08f2VICasEQmDKGYK8USWMIOjBLf/2I5WhPv0UpWAHJCnaZvJdsTjUwAl/oj
jgJ45PcTIkxGPuhswkjPAYG3XCHOKD0fcvxrc8hhsOral/YksXPozraBSPunGfqT
aphd9Ds0I8ZGruwIR5jwk+R3I8RGNhHfJaz3i3Gapzujwp/6PGgYsnxVJKCBNequ
8Ttim6CV7RTR3whH9jrfQIjbmflsMzmhPs9LWWV9cVxcgIAQzzm3Mhylq64VBRv0
9qUHo9gGD7KX5B8lHr2y15YYqTLu0wzAxYiONU+eCtU+f58rYZ/4bWnrX2RBOrGQ
Qd8A6HRxL/KgQ5JQ35/IecWqXNfAx+u2t0e4+ydtMzUgc+wg2pnz0lJLFYpZmGWP
Xr+QNRccAnfq57R4s2KD6ZyMfQpB7AIHILzI0KX0SqM6490IdqEGMR6CFl6ljlUQ
9x31umsoYt6oEIMO2ApI6N7hXTHKi3YTPbOPau2rrHEzivcERLNmgSZAbLzaKaNb
tN3z35l+qaBx0T97oWPpAbc6AT0HdDR3dT/AKQJDYKDwBc9vLcQG8DEswsLGy5oh
dQ9dQP8f7YokJBk4+gv/BHA5vik/yLzKDGZrDi5q/L7H3TPDwW26GA2765/FWl2m
31t6XIpNidafMChRoFezxOF5bBuG21JxY6heRfA5Pxow6YehbrjhJ/YBPKbuzjVw
YnF7GUGpG6Zr6+gVyrmhcOj8PThePwGGktBHPttaU2kiamYKbm3dp2agxU493q2Z
71MEnqjOtDQE6IVdPYwyQJatcDlGHNv5fGSCDtY9nAD1gOIaF5K4EFI57m1fxNvK
grVxam0P1benCtHwlwzL4VdhqNkjQCXpp3rQKfzg7y563o1e0m8KJeHmkzfqcMRx
8IYBeiRUeH9t8bG9CLoLGqJTU24ZZZDCN1rtzhAh2Dq0PB/LpJwTz6fvdelmydhO
mBcgC7JguNHwUGH/UZE+l/SSzIUv8RD3dM8b4YioRpCM8BlY4UDMhPRVQUNB26d6
uYP4qY/49PJN0PsXHlG+UDRuRHP5vKxDB7hbxhC3C2P01YuxDqwT8zrPSzVhMBfC
3b/qevivdCXIHZzxq58UiRGj+JH+NAO2ihKtY/UrKemnJeEGmTwRjdVBLkysRH7j
/Z3oc5w1tER7d0Ue/5Fdh8W2+1zY1/UnRdYO0E/s1+jBKsUqFevqIvf4cyhaCpxJ
XP13KnVVCxeAtTTxj8GxxmznbXjqlfhdue/aSuF5+6M1nb5ZCZXHo7ty3YQtwlAs
5SyUq4w/GtUK+AXrXX/Zr7nZWkBaFWPxlZmXU1Yf9+ycDfC/kcUIIU9JJthVhpnH
3DgmaRQJ8+kcNgAnFiyDt3Wh0+HLHCzf/JOCs5fBIitwgXMNDCJzFxnQ8DzYAmgo
nIqyLSBS2hEdIWfdnK/0I1GcmvTYwid5ptyFOcy+njq7lycLrhCjeI38jXfBpay4
LKX9hZlDAXOUaP+07tSVsDhUX+/BMHJcNlsX3kDAgJ3fnUr5LPhD5fq2y8opx8Se
Pf3e2oyiueEiLXciM6PKBcejYBMejxQ1BX6z/tOSqVuiLBttWi0iUec7mAvwrq/H
ulE1fcJs4W10tsjErt45seEqVAlW5QPIFPAPiPCQm9qjL1ZrRtlOYL2OJV2B+sYY
iJdWft4Tv4r1H3T+kvmZG0k3JxV0LGJuKYainvApW2FYoIwQDZ35+8aymh40PzUd
g4FdB4JhMNhRbcw1sHkx0Xs14f85RR9dXBv3olB15+wwKuMpYDbxNN/4NpVJT/zC
H6QXnUVnNP146pB17cX4lV6bh/uI1tQVOciWKMaIoaySmBpTw/wBRZqPxKfdKzaR
DcCUtUpKau3l6ROA7EpKNUUM5etPvQLQOs3OqUgxNlSgLsemcujIrLo9eUYQrqMv
SxDy+Fu3caYC2eX6ZK7xYyI/ETA+a13cC0dOp4zdK9AyjmscDTa752NLv/klVK0c
gsrRji/QBzv2DZjZ39uZaB+lkmVurgnGMr8735bju0haZjeLpkdLOrDfK50c73J5
ss0bisuFMLqAYQjhclkQNWblFoKf92saYYDvbTC3U4ewpN8xvzm85xJbO/wDtc1N
KAtSpFUxEOiGIPyrRnd0ImhYRNnjNkSoxNBV3PSiG6kZGMu8DSOdyq/MG3L1abOm
tCy035vHzQxee0pXazrctvlWm6SfYYsnQPhVzjFXTQ5UHAwVsGyaeILT9digWUpW
COLUuseb8nbHsTBYV4MylA==
`protect END_PROTECTED
