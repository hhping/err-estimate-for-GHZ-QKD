`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vZLnNYlsinheZvuLH1pPEvcJZH3sidPoIrDIdeG3kDxRCzuCgsE/4Au2ibgt/O9n
03OQy+tjwX4ZpCXkhuop+gqUMVyW6BYclJ4G/i1R67YbacKiD2atCZOqvaLm7ojE
ZxRXuMhG8gwXSbswHl/obhh9FGsn1jWTzcdYBdzi/R4UdGjH/IywkYoD3J3CKS++
rqaFLrYfiephL+gj6vNKLC1YKopgXYDkg39qdwYi3tm2XnmlMRegf/NuAi5MJcID
ea6G+Xs7+dwKCGDqjfu3y2G0SseW2Im/j5AcTl+ueAPrw1mERoT4mDE0u41f3qUX
hiW0iofNA4mMsAAmCmQ6eraTrklt0TupOgGl/uNxDtWdc+mLLYSwL3e/ywisVEQV
Rrgv2YdePr2Ar0QCV8+mxskOvBwKceREotDwLGuWlD61id1uLyG2E9EeMuLk0prR
cmwB8HMIoLJrDCd+DAJ482Kw0lLrDG4w0I/4YbCxO9vIkQQiJNGP8QyKgwVGO0LQ
2b6QiBajLZyKSXEvfvZghJV2op1IJAH9+0Re55Lk8YXIN7QUwj7LjETlIUhEweNq
3o0j5jdGputxs9nwsmvwnhjDqK3M+A9afmt+EPM52wKMnBr5j0wfxXgefb4pWkCk
QM1MuY7If45aPzxKO0zZIb3c/nKbVZgxrKDf7p87GP3jsECZ3W/iUGvCE63woT8K
LZfTcDQ87OuFcIBYxMgOVQx7QTWrvoItFDqESAtCC4yrpt4uM4JWWr1HN8mRtp3f
9319bITn7lOj7qRaCBY++4TAo8BAPKGNtpkpBpl0KYnLTSfoJdyIkISblNmTubTv
HVKEGT4LN22uaDA/ubIf8Ef279mz7yZfLU9HhGcM6Ycf/Eefl6CA4XOPu/A45HNa
aotHKPyw6oSFaNljmuS4IQzHgJfy89BFT9mlFIKrC3m+qr7CzyAE9VNOBVqD/3XF
YTGr2Xb8gt8G3zd0bW2uI39w0xEzS6CvaGIn6lSNmycPR89noslzGC8uwVmJMUXw
NHXVCp7vnxM/psO+RjG2+IG8mfzQuMB4g4VcFODfD8CeHhw28cbiLcvm5jow4/O2
vHtPH/BWb1e4GhnBkHzZoeMqveX/vLTt+kmtJOTsRGLtlC7/FdQkR14plVYJ7xFE
2tHzV+goHWtrk6M9u3VHACAOcimP+Hola/g0Or2i9KU6xplOU3pUpmJROHT1tDxq
+0GRx9aby7ggI2O3IYX4RfU3v9rzkWaI/0qaoujqMZlrpCjJsWgmD3HKWoqKi2kA
acQ47qMYzP3LhpwdeKE9i2HTnKoSdiHNMnwPVtbg9h7qsaaiqAfEEZ7NQ0jPl6z6
4lAKIW7hKoTOpn9SNhxI0+Uxcqv17DTOYdllPryXjPE6FrRxet+O/cH/Sw75P+MZ
D3SNmh8lNm3atX0zAaJv2BykPJ5t0LZwULtQrrW82SjFws93/3ebFBmJSuedjjcb
ma504U5jg2GHHLEkuNa/AxeOO8jNHemyGPPZPNREqjGR+ijTu7140XEUGFuOl6Gj
TStciJdRajQtVzzZVWCfG805IvYAqehZ5FXr2xA3I7JeIN8E5cA9V8Mo0+iRBvWd
bp8vkT9mESjm+TqsHHrNKJSi6FsBZp72bJ67umlOisKH9llbtYCCdcgvFmy5Ev3e
IjSDpaLHjBp2A9a75ci4z3L1eMXpQgVmxi28hHuAtukMpWRm2RWSd+N7TKcKrscP
+X32RKPnsEWMWhHLs+DB7wHoIkIoLzFwRtP15PokAspVHi8Hx5YQ5jiSMAzS/pEE
NuCz6VRE5K7AVhMbvhtfp00/NsUI/BDdptcHSuICLKdJ/iDLud7D4k5FXr/gLMq8
6h9PbqtwUxCQQbHigCbs7cukUAwnN+WMIZfRPyHgKniZ9m9T70IY4A7unqgVWPJD
nCY8bu/x+GjhpDFOf2oqyv0s2svzoXMIwj0uYzcavJCqLnDehNU/IG3K796pJG45
A7I+8QTpwXCNKg3qNg62wcwtcyzAkyDdi5WRwRcBx6PlwjXK1hEFRTC7wsjvqved
b3EShJ821CRmdmTsyBw7JbonjBDdC+A1HEghERXYufdN1Y+qNHTZUwCHRh/9xAFC
QNomth0jZa6ehNkM0ATh+nu6n0pUSN9quq/AlJiEk38wjwm2YdNCxpaEnt4B7gRd
ykogX6Uf29Z2sXA5VgUEbfddjYbstEWLXxRqw772qBRAcn7P86CQBa56xLhjRqQE
g82pQuEo34W1VMHSq8Q90J6B+YlIUSAqZUY/H338kYF60ZEchPSxdd9HZ+sKjaIt
+iTlXbV5GlDWt1QtL/SozYF7NmbG/U849ElDAnFKNOgnmmjjuYlaD2hzbKXvUE5P
wb/nDXNjWj9UD3OgFgfz7GHaK5mX01VXPgaFmsaa1xNDQtLl9j4a0g/NHuVjZt7v
uUoe9i1lgt90LaXobNJ+0BP4r89KOFngTzxx1xJ1Wt5HLQkg0LXprZ/3iIj5ybRF
jXQcQfRThgnpegp2QZUbn2Lyzy0rdLfwZs0GLIo8u+h8V+LTK3r5xsm1YsmHKjMR
R90Vsm5aRX3qCqFgtAMHm0u+JglvOvAesJ4VSBSdRNqIIpAXhLqsPUm7SapFbK1m
4dOQP5Z1RGs4OZXvyRAhLMu57ShrLk4wVRJE/BnkiTB7TdnsCb1KazhKOXHTJsVo
zyaZSMoS+NNGBZBah+ookzXe4f4Vo34yq6sB/4mtWWIgIGz2sR7eT2Npd0hGKdhu
Kklz0QFqeSJgbOygE6shpUweF4lcNzEuEqDQ0mDGR6Jc2FjLVnftuW6CpLTcaNX1
5jPZbxUCrhTfoOlykwTWS4j7ifKhv8qC5TIy/zqJcIJO917VtxLp0U9xJ8zLGTrz
s4qe4yqx3RU3mR3ejWZubswQIbO0vAZPezgqg37cPSxwzGt2H+ZlS2mRY0q81PUA
K14v5eZJORnc7pH9dmr+FcQKWYqNgpvw4TUzLRzj0BOq33t93LizG9wwbnjKjXhW
o1kM8LJPUckNC5edxqjLevOVUYzoM7/2aRBB+zn+Q+Ya6cQaHcTiv6oJjGG260oR
3Lq77eHXRlB572RsqHzMPXdh6ixMFveJ7kOgeIYcc54kiZ9mkyy2lJH++dywu60p
F0278AEcd9WraBuiW59nuYzjuhzjwyPao5poYNxEOb7A+7FCiGDP/Ue24S8ammq9
j6u68fHNhz4LE/2BK6DF9gG1k2cgyruLAPOiwJpiKwBvjMW7d2MfYPpopFRosV3R
K9d+fLRl0+rxAy3Q3j18iPUG2dXqOOr3NVYmNfB94i9ii3CMcWa1xUpvs0HT4fWB
fU/bzDKDvsGC0WPCINwCqv9bI0tOcPJ+13kEZ7V17iu9Ptoeaqaoq4h2vgo7vpjO
MiXaPd7Z7+gPzuexGdToW/uzTehZDLva9Z8ueFlazh58i+f/EdpLZ7Xa6yRahCcG
etIqPxWwVnaYNkUOpTNQJaQkC7qRtP0h7t6XGOM4j6BuC2M23rT0YTGUdnjhHXzO
X7UD+IwQ1GHNIFpE3AIWN+Pq8iQhnpw+Cvy8WE0A2PPjz3mftJoKz1bcpXnpqLrw
glML3/b7gjB7NIknIyWJ05SDswsY5SiGPNp0SHj/cZrdhfVs2vWPqURkdHbCTRQy
dBPxBKzt09CTun6tX1ErdfRl3Bzmjgjq3KgRMlkRNiiTcPJcQmwm/T5b8YSSsqEO
pAYP5Ryl8RXzFPFkoAqy5RcQNuwTUF1V92KsfMmzNmIs4InXMXriwVgzOjurCEgM
MbMFdOxSsUXJULNSdDBKWYMx7x3kR3You83UTlHSvp27CenqqOUKR5v3rTOwPPI+
gAUTDwZm5iUj6JT18ULTOSMJ5XCzJayYW67lnsHCGUwKTLzdVOucI+jhuCLDrMh8
GuB3gSX2VO14M28K4rPeLjfqwXEMpBZ+akiJa+/Vq4a9TKjEmHebsNk7zp1u9ACP
09kqaQZlYWKomZg37vxXRvv/vxOridEY7MLc8yyDWmh9jN1NSRNNuvrjDipuiZSb
RR+a2+fzgAEzMSq/BP7NxhYeS998XMDo3fd1jV514FW9g1kgzGq6/LanGZdM4QIS
no80JNW4g74Ep1mQpAd2sBP/weiP2HTZm5+Pnu6NyWWPJFyrr7josgDTXQgA0cUc
76LZA3Axcm7kWLEF9L0qzMyeglquevjHi/5Xn6/0F6xgiTLTAQC7PxCBRnWx9bV4
cNvT2PPkBp84UB4rqr8O5WOCt4VJcly1DgSBT0kcsxhsIM0mAGz8qjRxez4ABjRP
NojG77WfCFpMQZ79ZelEVMLcYngfrUY490bsPWktlYpRgbdKzhW+/b5YhX2c9l1H
88FzqHVwC6hdIei0CBc0Il2jv94rF91PQTBZZSSIt+/ZoOyR+Gy46yQdymXA9Udn
zcLo1WFTXzLXPTvTDCuDGKsuR9bUHIe90LxXHe5ZR2mF6OMZ5GIhFpu5iyKJg0gI
ACezpSGbp0LldeHUuuXVca5W073HKVVk28vCz/n7i9hs+g9nFxfzusYyoM/A5Zjl
IfSj16oQv2lOCP1jKvuWoSVFuGAt6CiobyKRWgRjP4GYNX4nZa5FEN5EILFPdG0Y
oJ0j1NcT2xUOB5Jeh9zJIXHD2E/pM9O6x6GmEhZhSyqe/fkgVYml+CgPjms+v9NL
Lgc3PBzQOjaaxYv1ov3TpnvCX07doNaJYwGt6QpxzQK0Uoz6RdQ0LTvW/Ai1PC/W
MAKkzlRDIFNU4hMEQM7nB6d9Yae4jKUi13rwnoj9a9akoKT5ZGAtb1kzZVLl65ci
sEG06NK3DpXjhCuHq9Mu2zhXcDzT7+ZPfxBemrPFN6vyZUjsWLTHM5g4ap/nkZ/5
O5pj8YFwno8orujchoZ4UokxoJKDnRmpWe0De94qrHHig3UyItlk198pzjJbZDf3
/MGJqVz1f4V2q/lJ28+2xEnSIpgwwvZEAkOHxP4wKBp93B2Sx1SkjPCzjR4ftcXY
+RUyfbNZS8+UBHtUDagIv5uNpyZmhko5Zjx/KJJ+uKDYAJQVoED8HEM4N+mNHeqI
FNu8u3vzSmU48P/LxrjIDFJhFvvGeMSq5B8VrnQKwWWKcxsI4jqYnxOH7477HDVp
3NJCmnhBa02sojoeKyL73REtZbggRYEnGAQ/gH9teKpHHgsb5Y6dX72oro3Zf/+p
9APPuC/l3Vs1tE377kX30pS5Kgr75Bn2gNU8MqNg7DM0S4gN7KPq7+ekoW29Sd58
pRnGuqSP+ADI51xUN/gXgfc7pKg7vAPhuPp+hHq6ISe0GRkmzjbqbYl9DSXIwAwC
dx//NEYnEoKAeduz2I8oekHSAxhmRUba8ShESkCUuyPAxBeZmTIKklXw7N4qWzG1
OAcCvUpH8ug883g+W5UtEjQd+fY2R6/MVw+qBtHp8hmybUSMG+h38QmwmTEXrjkd
d4qHAur7XAeqWLt34IJJEQfPqmbaa0uiU04d25Cn6LEBGhYJc30McaiAL1wwOySz
hfM3n1boI+ZxivuMSIY5QVjIlIoxB3dDtAidKAJIfiT9N8qe3OxAVLi5S1ipIqZU
ERpg//pFVGlAPd+101fhYlPd2tSI4LYvD6Kp+0BftyvFWVk/cIyHw6IGpTIR8QT5
`protect END_PROTECTED
