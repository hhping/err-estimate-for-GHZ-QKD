`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rq6qF8oIEv+tJTuSNYy08jOLKuKr/voyKybUWW6fUmt77H+AZmw3VXHYLQb3sHUd
bUANUyTNJ7ijtsyYyJpwVdcvmObSixJhsieMEXzHN3flPisHtS8K7AE+5A3jQ29k
USVf3GovKMiCpEOGC4BMERS/iiSM/Unct0iO8eW4bKJBTq5xx7pXadsH5kZiDCfu
m2rEIbKPILMCKjCCGYwN/avkkrYG4EUCDm8ouhYu+xC4B99wq/so2hV9w3PoDYiP
f0p5BbVYWGCWPqbp10S79H2JsvowxqxFRBqANC0dpSbszMJN4P1D1a6nApKq2lpW
KJbYMC8+gYB5hpNFm2Z9+Y3PRpMTqVX428dVVW2aC3F85bA21HSrygWeq8Qhi6Ys
zwuvKAXlggDfCcDwWUFOqEcDufaVzCG0LitiX/YcBYiyBu8H8068V78ya9rMYE2J
F2TPCV6MHX8TbxZWjKRGoTvVXC/hr348VsndK1RpFCgg7/EEMvTIxb9QuDXiIvC8
AejEKbjvYiGjH1eI1VOSPUO6JW+8gSL5TeTboD2qj1S0SquJ5UO6rnUWPbLSFPPa
EQzPsa9rzDjEBKIhfSt+9A68fzaQWQMnQjFzlxsSR2wZfr803aSsdJox4zZsFL+q
TH7uUCzEp7pt7puXOhcc2u5jhxpGw88VA4F8TwgU++04XFwW6Vn8Muwl7wzPPWJK
u73HB5vC01eNBOIyIMA5w8WAQfj9cfUfdtjAqk1Cpw0otEBEG0y0vud/w89uUELF
dYmrxF0l+ofdxJhB5Oey5lIxoMEVHq/miit4RNIdsnPc5cYkrVh2HbfPd7fUTEIc
gPVwqHS9BKgMf+FTBjfFxOhAIvAwCgMCauZ+bvwytUavxL4oTNT3WV5vaccIG29y
mR9WPr0gUGQJv+QL+QO5xMIC2qaBltn25B+buV015AcTSo2NA1Hn0eOqDL05re3j
AZNibuA3EpUip4U6m4nZUcGKqCX1JoQ+N1geHRSCdYdiLreQjFMdXroRFZqGR5QL
BnbNv/hGDp9mLOuqdvfG21LoLFRBoUvFZ5DuRbHV1+nJvNThQQbC+Gv30BQl3lG9
1Vt0RM6dSSmvBGGFmqfCXOauFhD7khm9RDWcqtM5zY4Bbn4yoB2hWeE9cVVn2HfQ
zyVYfo0tBROBjZhU5tM98nJKA0cFRC+BKgobmg8IhsukEReHfEdzkxL2XPbXVTTw
TJAqetuJ/FU9Dhbm1SqLXJMZWq4irV96t8nZrycHmgHGOBSsBMvIOLVs1PZXC+0O
XDoWAkIaWR+50syl0K5oDmvD/J1Mr1jSb+WXiQPH3981sbxmXQcEqs2Vg9dSUdfn
xIZGUceTIvUB9aj8nfvdpAipTKseI65tnOj8HxrJyVRIsu1DZJJR4F+M6jEIizDf
P3nvVB9yt2y/efELbtImwAK1eqfRC2CQ03CoFXITiurDpdUmmYpy/03YSkVKHdWa
BPZkAklX7CcNUAts5/qXZ9X1kDpCEa9Uv3cuCiz9rh8IPWdzxqKCGeH124nj420U
ATi7c8XaIilyjvxh3Q2DX/tSKHRpiFqIA/5mrpBm+i24BjiWykBF0BNjTXfmAN36
YePZA4LstloegIeBYKRf2ImumdvwfL6ohfrB+iXwaIDOti0ew9yLwloHoj7OiHIP
rUw28dYdL778nR4ZE/7Z5comTJqC4ll6p6EBmAWbKJ5O/EJBq0/mYRzY7tir6VbS
yVuwHKq+oEIyBeM8lWMYm7A52FiEI6/XGuxXGvxeA0axT4z0Q0C9tTmrRiH/LH0W
YFpTMquLQ52Gqc94quMJTl35AWNol3XE/fAxjipZUhRIclp8W+dkv3pcORIG/2WO
Tto8P6DdMaRLC8YtTApYFqjHpZFn+gd7qPC9iEOwZysD6Y0/MiGx2H2XFTxwi4Do
SZBdwjZoPdSAf4PPEq+LwMogUSmIYoBpJm9Tm/iZNvCZ4kb/78w4IAN0qF7O8da7
naUC3XwSH8m9kHXYkJY7U2QhuA0HsUs2bqmLFgicOatC2nEX3WaQvIVHKVApLSZo
kpyLRs/9ussgGbVx+r6GlfHm8uuhk4TOC8n+6VRfKFgbUJiTUAbzqopsjX3BJfdN
Adugdk+DeIkLoO6B+Ym7LYMON8okIFVVrHDezJILscjI6dBrGQRDl2QDrVlCk+4c
6ZfJjE4hmSyA+mXWLPdBSQ==
`protect END_PROTECTED
