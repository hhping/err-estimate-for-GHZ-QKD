`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0HX2sZ+9sq3rAgtejTzEmuEx9pXRh+vyDWoeWYJNtYJrjcCd7Q6m0KPJk1/FzCoT
kkIDTD2QRI+misv7+3OmhbWXBHgUCsLtSSbTcetL+i8SfQIThiXn79Tf/7nUjTaU
Mo5S7kzeD9ii/8bnrm+tMpHZinEQO259graeXGcYz9AdvTsC9RfJ9AOl2l5yQN6W
QjENqhlIhCgjpS6q0ZHOhIKHoOBFKzs+Xl50xll6YvPueCGnhA2/233JK1aDkfEg
Fok/PEM19vEDFfnp8a8wON/D1ciApOv2E/x8LY+QcuZDqUy1uMqW1ltddqMQxeRp
/5dHuemwt3AW3rC+lTXXFoCST7X7Y8PCXUjyrHv0D/QdKzpzf9ozNH9db38hguZk
h/CyHHPax479hDHKV6o0skaEHEZRW5QLaJDHteWo13NdsHm4fQIKEys9US4ihd/B
omNgqJS+cNhg+cd+nkO+kP93/lrDV3ycUXiL52VxCx6j5DcdmqufNCtLWOlxK7uD
pUsrFOGr5arvwkiVqWNuyXzCw2ZRHOJqJE2QvGJcXhi+uouMCcP1CecWc1qh2+K+
1uv1haMDtIQdVN8JcbmaKWgcuDr+1qdaEdds2EFP3YyYuK4yV0Xf5EZbZxFsJio1
LsIyijSC+0nO2trJwncrWBmN8oMxRZ9pdHOBQzvMWMA9SsdXYAdxBihPdch8gC9v
Z7iqSPmv5Vjvl0vajUwuVaS4eEg33x4ER6qnm3Y0qIzImVNdBca8HZMG2VpCUsoZ
RYi7HWoEq3B25Hy1uZc1vsAYXc5T6eEbcEAS+jPKRidXBR5a6Xt/8vo7rknf4gRw
AwTwXU1h1XyKPj4i0jzI8DYV5ysaRrL/JascjdoNDY/CFKeCMdCj6biHXnC2n7+W
+4aorV4lqv3ztiHmYCHvDQfAzuMJ9hcdBmJyUslPUu8=
`protect END_PROTECTED
