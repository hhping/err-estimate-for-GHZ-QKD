`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AT0rUXYSn35Mcr1LRHv16p+pKp7SbTiH4nHWWWq65wrWIm6CzctSE+ILmVpt8iPT
TE6sRmOxtJG9GhajjG0HKTkdEZAqd9oTIMVzLyRLnyPZUr/xG6sQPRFt+on6cYlY
JV1nFPYw5S7fC0vKqiy79jhO460M0Ex1UN8BTNJ5h7IBhgOiMe3qse3HVEe9FA4L
aSSwCeyyvhrchHNKjlZ+sNZw5oU098H4Jt/SCtCtw1w/rAWki2gnEUFrISP7f+GY
fdqUS2EOaQmeeRsKvky9tz4arbwmafzPF9uAdO2GCpO8bwi+RlFutXpl8uEztbtM
dy2AVWtCqvove6uFo9YQiGV3EzkU9NHrCv7g8fHbrh7K/59hOlt4J/X/AEiu1wW9
sK69nqkn5ugS1OjjfJHlPX8g2F1pbbSsVyMMKhh6Ozu30ZraKVK/cz/kLwp9PaSV
RSNDLCgz5XY6IIl0UzmmzEB1ZqDaA/JjROjF5DE5F5qp9tb7R6bdy9ZTNbf5U0ra
ziaGgHKreixOyRgp3aUhie+iBGfx1jiNLevrfmTNd4J6a3fVqGg3lldfdk1cO7Fy
VgKUpzt2wAyjz6gt2zbGvghhZZKex/dAftSGSEOPYsvF3t284RcSfr2kb5cbnnDY
V28EZq6zOhhRvgUzaY7A1d42xxF69iQz7XFUhJGQAI8=
`protect END_PROTECTED
