`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+i/FH/vzTE/KIbksCpmlWxifAHAKTgj/0RoJ2gCooo+iwky0vn+3Bkwnk8O0wdjw
lHkE5ci9vIDQ8DXE3+5sM2Dbkp8ae/p4BjwpaXJJAVoDv9aBWAUg4dcVKN33XhUN
WI6xjzMz/OkvFsgIE1A2fMnO+GYHaYQXx3gyNHtENv62gggHigdqVfbMHI0uIefy
r4ohVddq10pUeEov9u86WC/R9Oz3o0Op7UEZb72zEtBi+bsd+T1vQyI/ngwrIPhm
xmCVASBRQeyHEAl6iaCAqaLVGi5rc+khLbqIee62140JJmWu3usRVZH9IOTBLjEj
H4quu4AtM8DzqK6DWlzz3NbL+n6Km06XrqlJlPF8L+DNSiN3BRHOQrRKSNDSP54B
jtiliDMPRJyOQ1+a1rrXAqkF2sCgwbmGveliTjjeuBAw4/3K6HSdmg/A5i5x+Ztc
skxNYsbImxBez/mqlCQeuDV1cUyYGUh9n7YujYenjRH/31NyQObmf4BUEMDLO489
oP0pU88LWX66HYTrv4jUq2jaGxuuqOEg9xKBz7t89w/66KkWSx4Upd5j3TuEoMbg
6/G1MhkQNl4m0eTO/Yjhcpq9XKeG2kCPBW4LOXIv4KV3juTBcEIp+8lmUdfYmsES
UHsYGrATvI48eo9dskYT0n7DeIUsXH1r/qdY88CG5SR6o+De3CqmbweMaoJsN65v
UzJt0+RKx2Mw4oQAtzZHQxTJtqeFbRAgX8+prDZ78cEEqex6H/bixfMGe0rct8To
zLsRkLFmdfPgkh+DbJL7qkzPNMJxiy6MDz/uIGBdMWpken+v+WmigJck7AqHtOjw
x7xW1tLw9ZlZgv0wVfDQ44gw4WyrWAWY36/y8KNxZgTeXLjw/JYBwdfFxGmiyCgx
ueWopSKjp/Wvg+3Yawqadr93DoON3BaWpn/ItDI62mQ=
`protect END_PROTECTED
