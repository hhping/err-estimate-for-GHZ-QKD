`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wI9z2uCVl13HHHDquh8mVTc63v6Eoz3Ms5CMcW070skleWaRMZz5Y+dC3dVFvVFH
uemBHVKKvWaorT7kGC9andxbYSPB5QEjxB7EhZekSHN7bofXHhAhIj+VzOIhghxX
SDXP5NmtyFU1SkoN+xm6GIajU/XGenzSpDpUMgWc9DMhI5fJmEhDH6ZNCf6EKXNk
O8xcFTXntUBm8/JKVgKDX5Bp6sM8KuDF4xJ60NIFH3WoSezBpe4a/5szlX0uigAC
c5jKoKhjZdl/NwkwB8ZE/qmhe/4egav1WmpqaxXg46jMr1v93KFN8clZ7rVj81VB
kB8lAVZGpeCSJA8j3+jrtfUzcRZUYplzEXrTXc2Bky0bszqoNeSag91cTqm1wchQ
pPfPDZ6C7WXvLfJ+maRO77Legr/knWnxQ3FC48IhhBV78Hf1rmr62kZU+mm9RgOw
OVcHGle8mcrWZHPiU8dma7XFyNfnvy2CayM4+jg6KY9elE0Ej8GD980y/pt1DCbR
gxFZxkFIyefX99DoFXojKLHWwGFX9xkX/MVYJ7geR6w1vF3BxclyaPqqF5U1GSMe
F2DiQzVFUhVhdsXGmldQ2QsPt0YIpWocg8+AUVbT5H7kXT3+ecyk+UrezIBzAOzy
GUnRWBdRIvj0Ll5cECykveWXpPPnjJX6rchNKQKQE8MNl7XAFzAuTCLshe1r8Y56
fIWWINlu8L5hQPYCc/G2poWXIDptLICoTCZV4o7VV/1zM9x6xJoiyOLWbaR6DGsu
1ITLR7uvvAkJ4BkQvbrG4cL21DkkJAXNu2pVNeKMK6m+IvW++0N00faBdoPxuVvD
z3Bw8cmh3ExOh5k3KBzt7ZvBRyTV/b28b7ttiQKX+hbD2s6yNMq8ddsLViOVZ//6
u6ZAws+Gjx8YmrqI0lfyuuLdFq5mSTp+IFkLFWgXL/ezGVHf693zUCEdt45q1K3r
hdfMvL8KBsvf/0+6luPMRCEukop6fXCJR24S8/n5HO5RCYx27zn9vwAm+D03qeR/
ShiL6W5CItrj659iVHKTY7d4mbBrTQE1+Ebj72J+CaQ=
`protect END_PROTECTED
