`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XtTtFdRZaQR9xnDYsQ2yTY/QQ3v+MLnndoxBUye2jWm8qFT4OrFuMUK/h3dzSoKP
B+szeNBD6O3wj79SqSW/5rOiWLP1b5TlTpBnpAS8L97PDcE3tyiSmw/GnmTKsPOR
zYI5CsBfciSQIuG+ijqV1VFZxPJ8sI4sF6Q/QYy+IzW/tP8zFawn+tvmV9LFkQ//
7gneF6XreVeUjWnC7ZN9gjB6HkbRlPG6VUgyfhHGjyJKriy07CIWhOVGiuKUoipt
rwPfoGT60B7nlSkb8VqoYP7fHwxuJw1V0gSn7K4aSN5inoGOlxQXF/367+U0tIqK
rce7yM4yvTjZG5r3ZQLJFu1U9TJF8j8qvkwQ/GbYAkik9eLu5l/cOa/1LgkZU6sZ
MSSREBXZJU3UV+WuL56jqoqidLch9wIqyhtwgODA+t9181zm9g5mloOy0ejTitcn
DYKMTXSHHI23qV/hZVVdOUgignHMRtix/+cFwGejHPMSXaayvdGgAWHBDOjVlkDl
gXfR1lhe6lv4lCxExMhy7LvlmyZ175Dl36cVaAB0muh5WdU/mSOWQq1+3tqPz+pA
I1QV7QVGG8PVlxVpuy+72dWHbpVylPwzL5wcPEppMw3WL07aBZxckofXvNN2j+QR
NK77UlTXils7UaLaoeY8QkaIgRK3Um2n/2K7qPawFjEQ2bVRIYOGODQtovyM/UZR
a9vhU1vXOUfYiSicvLhI97PJKET+2/luxhapMLn2OIjPD/XLV0RXIJkmBz4Zs3Am
HdobjakO/B9bgkcrCEVCFv2+kXVlSFTOadh3IDiVWd3++RP/vL1ilkyd/KqGng1Z
0lYh55v3oorRmh16xK8hWMyLcEJCX3IQ/BOWnxmMaNJnRUgvUbO/KmbnLs7PJbL1
Vk9caJ9Rls4QFakDm+1iI3gjj50wsAeBQY7ReWrphHvIN6JT7OVxyVmcs4tKl5m/
OAdfNdV7I9RbxCZMeG+uJ0zydGenZ/mDCgxXGuT2510FDM68ghR//NM0tVMd8kAV
iUYK4Wa79+098T73Jk/5dHSt6TgRJ2xr7ia0RrDgfPCFM+54vsjXtpOOMSraAf/j
QnqNcDdg0ql6FxagTRstSD7CcbabMyYspLmntVQyTP9BjAeKi4V0d5VU5jlA3hhp
NgatjMbkLODhbx1uUw54yzG4AtfFxQn43YA8HDzCYcRobf48gSQlI4vPsxn42bmw
hUuNzC80DM4SqzAE01Qac+e06Bo9NGyC4T+yYifWdcftmUENDWKq0ZAvrwvM1cCB
LRwMIAUEmJhpPC4PBbSZAchki2ylzAY3nqwcfmRGJQYOlluVPCuLK46l4n9pFf9P
UvliH/WXdVby/Fw7a6TA3AhTyBarV91RFOBawrdm2gbiNlouKqWycGHsNJ29v13Y
T19KyLLiHMAj8nMWEIrj6WEXBDNEP7aICpvbeJaxL4xW+IGv4q0ljQlY45phZ7Ns
EwJDb2/2CWTJN916ZzuDNWxxYJ4YvZfjw7DGT1MIciqt6nz5e//M9ReLN0Dtll3n
KV/Am6yVj0b4T2zgS0I8g487KWStj+Bx1C5lOJgIb95c0N87W1gCO/MkH/GnZkNk
vpy6xs2Oqquwu2iSsXdhvFZTq+x/lJ/4t/UYqk4nysGdNeADx6/kzg4Z+o3PXOpB
My06enh832l+DMvxpVBJ8SHqibnNvo1y7OREikfUTtNY9FbMFlIMPricfP+aZXBk
5v/nzHc3M37N6HRLfe+K2Q==
`protect END_PROTECTED
