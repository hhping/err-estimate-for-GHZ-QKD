`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pw3ZB9I+Wnr+32tiujLv28oJ/v00SwYbHujfNidVPJXLAwTKp4wwJqNk7q7uYsWt
hf4e+28Je9LH85vIM4baO3pOBbW/6eIpU22O4xKwTOFeyd4HJZ2Z+/ScN/uCpQxi
pv0AoWVliVHd6SW922xZB1Gr1WN7Yj3ApFon+p3NTQSvxxKyHBwbbR71dk93MPIX
ppucwrerlrxVeS+pWoIcDWR7d+sK0Zd6i2vMkhkoZdbV+0s5NP56txkcViOxlDeh
8D5wqkaerIBAFlkEkkXZqkmmqwxkcLgZacy5+oX8tNkvGjr85vtZ6OCkAhmeJw3o
teq5U4Mk5J5ahM4MZ/CLAmrOcz+NUNq0ZwjJBIB5ylw1XfPNM1aX7jTA2DNOqezv
ZnFsq0OPMtqIRZLyadL4VIR3Ipc9pL0YNjXQ5gsVx7rNsIyE9n7yNGZ4ThtfDjS/
ZLlc1SsDzCvqXT5gmrU7nHI/1m7mRq2KlKL14+3qKuyXV3N/aqCZH0mrGihV+p9L
oqKTgiezqqyGx3W/eMUalrCw6G4PokgXp7VvxWYKeLro4Bc/9fIwjdFvLlNbvWOR
daFwMHiQKpbotulgsGzH2lLmJ0V5meq+QFiiG5QQtwfAg7ygIxEq8UAZiU7yEnPR
8jZ7lve/MEHIO4R52ywUTs9/gOJTxDyoKlRGhvUVEoaGHevGUUagge9AvmoO5fQG
uvosH6qL9nhH/XNbXhwWkne+9NQ1NsCi6pGPmhuMlw/wicw4xoNU13hLp3y5xI1E
TLvufBjrWdZDUTPLKlet4UM02LSplC21KIV1hOAAOVPcMDERZcn0H97k7iuN2fCG
VCgeuM0ff7OpIDzPfU9e1/Mk847wzs7nUYX8ZMMVKugBj/7WO/V+RWDT71Ga7Hr3
k2Qa70kbTtK72c8FZE42PgyzaVmnS4jgT/PQMQSW+YvJPFEVJQ1xIXfv5BkVVTgk
3fkWlC+82CAPFgaRVe05TGKU3H5NXEX6FBHL8CMx4Z5C9w+HQPxKFr1mVDCnpD9a
sGCbnvhQkIfg9mv9YS56AVvkt6pMcjSfLI7JqpPIgo53Nn2Qh+DzdtaMN84uamPC
sAQJy2CNnoy0jNciFmjJKWRKeaQtaa6JHUdFDx57tmtTRLjuQsM6PWeFbQ6I9984
kKkTt8UqW+FMBcuLj7GgRfgnyZllj/yC9+MKuxXQcyN8eO7JTdhIUfVJ1454jcGt
xUiYpz62chEX+wB9SWjLVJ5zRucDgrvjMAN6XUdXyRRCVi2RevKSv0SHQ49D2tgt
yVXsBEz3VhzNyFv0T1Nrau0m4+Fsi+GSpAITIEA19F7T3AGI0fQdOpX+9kuBDj26
X6wzxp+eiE9d+4BvwS8i9JA5uZctYrrdbpWmrRx7d9pBaQK4q+ZaKp2P21Bk361B
ItfAVhRqUhUeuhb3aql/fIByNB5TeZtx2I8kZeoe7XQFV8vGvB2HV7ESt/hfcs9a
H264Or0gnmBZH5VFRYWbn39rG/qZWeasuGTjvJd26/yBzkeGydtNXJc5hl4yuAPL
7hOV1SnONvmGQFAFYzbB0mmjlDgA6WqSAaekGRR08Ccv8LNkzWOWeh4LhxoTlDR2
b3prrmu5b8JmZAqOPAfFBLYcHuUdz++hsZo+kQT0bMVzmd+Tq+1Gi1UNykt8EA5s
Hxa1fKyPLHKeqBjV3iLoKbzz0LDDs+Kvox6qz/LktIqHHEuD4wJlettYVf4kQdvf
YSfYnW8qFbZXnTftI8xGQFZ3gIaTG/yy4mWAmixSXNeB1QyovnJbqc8LNhG/cQmF
eFZnJo66M9YnRIX4V97Xz6JeT432HBpF1B8j3ALEqd0iH8CdzRBf/NFMKKhfFO2i
3VHlQtVwZT2EPCb4GmL96yZX4VbGWt0hFmjhTezHEpYGr1cwtId0ruOBpQMqyZMG
OEnXir1mhXueSI7zcK4PguJe9G1GVzEMcfeefntOAJCEdj1fnZJuDu19yLcAN7iK
6VTwjeB4xVcXPEjbCfpy+mkz+RTlyTR2xngKjz++JM01Iagsj3wccIjQkmHP29K9
No2YNtoT9QfWQKOfsM1bMHJh+Uza34l4hQYUkW22k6mNWtYKpafYLXPBAQOVFQvA
4j6kvDSw0bGLPIO/UmlmEShd0H/BJb/bgrM3cMXmgpPMK1XRKwpPsqMnKHf8QHGz
GjyGN+jZV1NGfPDhVCmKr7bD3gJnGiQY6fTxU+xLB4aaNLSnrtqzyTE5GycqfS0k
/EPp4iUm/uga83twKEqmy6fM+WxCiUb0T/eFORDQ+5qVGBe/69VVL5ODkrcvWdln
yNm8DyDurJbMA4vAyCOKx0b/7o0o8PkCjrNvKY9N9Tw9UTMVoUevNjEkhZb5+tKO
Eyfw222C3+CzSq5YA93PSX6/+Hui4wCcUtVnclp4XCSDQMMqF8mIdPs+ulcvL2Qs
wPApZKR2i2gU9TUi4hq0gOsnJUC8Oz7qfEWGA3a2XlqCNiHUDCCfZH7xff1ZyIHT
`protect END_PROTECTED
