`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lG9PtrCK9CAw5RpwvkLucUoKxy3unPVEZBMhF110zcQIsrjTN1Vwrf10iguuxLrG
B2kB0CQup+JVHgYgidMPWmzGemc9pH4pyEt9plVCER6mwP4I0dLD2QbUBMkv+y/d
4FWtlkK+Lf6btu7VkcZYxmccE1dX+saObw0jnGeG23yeh+DXCbYveMILcAHIWn5w
oYelEYtVnOT8N16skWdFOQIhOxjMR0Xonm1a80TXu4qjPIashWib9wRZnIrEwzq1
xhHhxvOG0dhcl9lwz4ZmEIPbEKlWgOTtv9Mziu1llr7PlnrZ2k+KSBkuheW0Xy3s
Pk7tVs+xIjKZsVMGgZHBwF8dQ/DPNDhBaEBCyYd2RlT78uxaS2ti8vWObQg53Kj1
bgNKUJhralUgRfEH1fdKDaVxM7v/9lohQ2KwxTT4+emwVmO3te1Zc3lOFOXaCLAC
JigqmL0aMdWXCNjeyCKqBAia4acke9Fw4QxR698/A9yODyoqp1ImvAYPqZaIT4LS
LUJmGkXXXtarr0f0YOyNnWv0TYi5R+9zDqXPmVr3zMu0UASbm68yFPr0uExVfyGg
ooJG8Ty/elgBRI44DKbhLsh+1xGPCsJNtPtXyxN3qkoqwEmrLNy4tgP0SrInlmc9
NvBYfq71iA+9P0WDN0r2YAMDuYw1aXete4M9mylvGUZ9rmZzZjepcDOvTlb/R95y
K0HxLDMGc970F/41s/hlM5thEa2lH/SrKvQ4jb53zlM+1VkN83UPpZT6XknUDHvS
0LC/lm2ofMCQ2cV5bBK2DGcu/LDLSbl4VOavgWVt83s1DwsLAazJEypPYS41wSmq
fiZNzfalT/4GioH3y5yBwnccxz0vlkZ+qpVNoiunfOuMT4t9BG6x6t56ClWF+wzA
tCBlSeSptNKUNelLgOaxzxft0BV8rIMKFFIfE0NUZpbGKjAgwong7bntGttbUrI/
0cNuVSJoWd4JL7xspH244zk6moOYktPy1kwR/Lv2EUPCDqBU9tIeKkPIYjDLDBUb
Dveq5Hp+6PUN/NtxwpMjTA3pccBiXDjNhitCyWf6jf9eACnsnP8stiZGgRNNkj29
ePrGCr2B2Jb5/3kmNx9F6g6J4SJ9MwTe5uAj06UyhlOUNXZ3w+rcIATsWKECRGyk
wWKL8egDvl2qjw1sIfo9v4Pc068/z23AegRULe3rSU8csoPDgh30UAp0ykkGKkXm
kQgsbdsKhDvDcAFUot7DMH91dfLgWoBo37GTp6khqNfUTzwnu1ZteOqLWK8b9b3s
gMwOdD/0puP11LXEEdA+Yr3+7Y5EWYljXjq0/j5YBIH7Dubq/I4hg7Htlwm1vSoo
oI7M+2WhIQOs9W/J4Ghy0guu0i/sGcVN5zMkqFzD/Ep2eO5D5chBYxv4ZFrBmbGR
q/BPcMJ98qy48A4Ax6EeymRRhpjDKU7mQfdzpUZBfV2AThnI8eUB1HPt/KRF//C1
n7pZ4NAHn5ZEPw4HUfQT4WMAt41d5CY94Mrg6sEotud43Bl4dhhxlCj6MO4RbeAA
4bauaR0p53LGLyn/b7yLuYB+dpLGjdx3lzsdDLiEfA4/Lb+9XXAAJJl0lDraTpzg
Xk1TzbXmVpiFX8TrGf0c92W8n9LFNBimT5fJNsfLN1SkE3ruAPH4MovLKbNJGIPh
P7nL3PGTXGXC1ByqCaiKKlzON1dK+vGUPossSzZKdh/ud7fqLyAMp5O+LnIUifP4
fxc+C/q0xUYbcAeyC36rfNiZIt/EyYZTaKSuZvM2pt2akWi2amk/sYVjauxsEfcm
YY7+3Y8/In3xXbI3Urz7XbBOhrlOa9emAdyADMsvqv5wCwOy4xGlh4W6AxZ5zeUe
2IsRcguWgl3JGL8/K8kqvBVPIhwYuR2vBSm6f8B3+vox/DAhrf/VlJ5/9NHxWDvu
ORTArqjUe0h+dg+QmDmEY86xhZ1qODFO1BpnOOp6hTkP/VjmiYhh7niMOt1bUGtp
WrBbXdcE8jYHLwtgHE7RMdlo/74DqFr01rAprkXxa3AQqgiEIoG7ibA39ATD4yQe
QH24A/OnO5rjL60e8YByPOb8206ULkPf8LvwQwVs1v3epmZrQ9mhRWH4qaM0BYcj
`protect END_PROTECTED
