`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S/+8zDnwMCAb1lTSs14YcMoTP0gYtX7GqMo4uJ6oGxD9+Gooqm4JyKnMq2X7HAkK
2w8zjam2jl4quFiX4Uqae6rqaWaAlTKr0Y8EhMp46XTDuVQTAXKlWVrPILndsCdS
VfvCeyobtASUyt37m2rPdOC0fMf/JXtSCO7cuk/or4DeC512hfL03+WrL2Q18RYD
BN2AFNvfo7g90IsiZRRXltJbCtay18v84rquesu43JqsDrmjbu73DDBbTchmoDSV
jb3FMybnm/ld3xhCskR+6pjmdIx8BCu1iJ8yR4lDcKdr70fwmd+bDEwF7MDBsLzz
DTSDpuIDwSTNKHDHY+yy9IrhOJVCsnaEAvImrmF+YnTL8SBfV6Hj0Zv+lbbAjcEw
cNQSQFvYra4qRGqY0Y0i011hqyWXZa9GttEv8m0GGORFt/v2+Ldivarax9TvB6sB
3NG5U8xb1B8S/UhCuoG73d7QmqAAl3LQvWgQvGx4E5Fv1fRXD2VaW8xTNlKQNmV4
SUKLxrp+o0WpgUo2YrPt3z+7PK7/KDtOZ4Abe0DUbz/rIE75wSXADo3PZ3lH4Xvl
qtpovyHZ5I7FHFEZM8mZC2wjb41HBpu5XoDNDvAsKm3BiavSqn53vHcB1Z4/NJPM
9P+JVD5Luh9YsZan/cRQE8EsmLFMAP3YdrdY225iHU4pt1Y9/SALYEWG8TacmIFs
TtjDYnMv2adTvBkq8K4+MYCUBPD6d5nmBuEacQdRrB4=
`protect END_PROTECTED
