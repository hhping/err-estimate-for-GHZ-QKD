`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p04KQecnDiCFI9hY4i4L5e9jqmq/IKpTfryZ1P+0QcMECmiGHfQQCbxWTiTrkWEB
cpDtjRoJIIDvL9EkzjVmQT+X+zmOfhIkockoA+WasG++KEVA3O2IikHAiEMdFZoa
k+fy7o1meXPb6KGQv/jltS8KiFtd+jepYUZZwVpx6RYYvoPl4+2HGfmrz0C28WlU
cB1VfeNcCCZlkgwJbxHTJF9EvWH0yP2YBO9vDs2GT7b3h1QOdMUrqEEdXL8Hgu0D
DZRxRuADwSRcS0D9cPBVvvfCbBD8RPTzf8mmy3ls+gRhJEWNoRW1RtYzpg3MlFM7
lbFcEDgX3WRpWMo+8dCisQQk1uSNin2BR0lLaGJM4TxJ3c3hjjNwmgm32q4ZQyZh
uoWG6W652hjt5AzgM9TziGUJkDiuoj1v9StTsey3p+L8RohVU+0YoAf8T5JxI454
hxYcuyvDNIAbZcJEx8TdhvebKNO4j1lgXUCrRCdwYIVWejEdOCJZ1TqQLIbXiM53
Pqyvv6HOO8ykV4OYWXWFWPK3RMHAChcMfsdMpCRRXa5e/9EcLgtlbZOk0r5OyY9J
iHmeu3zm8Y/ZAGGv56RWie0kEXIUXoHDRLSsLfD1soYD+FSiTFi4yDqdxs1bR6+A
RTfXjwSNlSJE8Fw396qFUy14JMtuYoIHqLhBVwWn4z+Dm/3HI6uLd5/VBPey+nuL
oMETS98wOGYH8XydqIOnOmNekOd3rTXCuThob1B2Zlp+4JQ7zXn9fJdKmTgPxg9N
B3J9nSSu1bgkIpIcNUz/ugAVXfOdz0Q+W6gZl08QonRp8L8lLfme+AgUOTUue4rm
DucLzOOV1Ypg+PwqtQEOIguvu2KRf1R2QVya1+afw+aBOAo+ZUrS2vi1IrqRmhOn
ivBZaUSxF5HZfEfREACQyrVIrrXZVMGW++TF4HRh5lUQA6cYT/iT9dk6cXPbL4xG
V2p+P3A/0am9PeK5iVD8ftWpgDuUbsT2ph06QJ2QvDK5Nop4eAFHymmfeM4xAEnf
hnDlCzCfLlUkibmTZrGcvYmbPkU/v/DJzGbDkyg+VhVno4bkH8gUBjL4Edj4OZHZ
N5aJxmGvx03s7FqItnOyqpyJ6IyAMmIJKC8kN49mPt+3/h34psaPxJ5HwGV461Om
OwDEP5RWz2XQtXBXV3zguRIOULuYXtUFu3nTYLDfJHkjVRDVTLi6ibhKNK+CILEw
9cqxv/aaqaP8EbmS8k5EDZWROW28hjLV5ztnIdzKsowD6eA16sjab3aVPfH43k91
jprp6Xt2by6k9cnBpyI0FQbgMba5AWD/G3i6krkm72g2sgEbNuwZcvaTglYiFSkC
8zoW3zg8H5lTr+ALfKYdW7A0ASMg3UscOlGpP3uReqGFfGH3TD0WC1p7f1puN6cQ
D5kFV7sdrhKdF6/IsEfnlynFKLBS6JOxHcJco98GLG+6VdtktI8mc2tKX+TPyksr
uT2AIfkQFmSs0xD/ap5pvQ==
`protect END_PROTECTED
