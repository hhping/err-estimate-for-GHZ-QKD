`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j2NVHCf4fJw7ZbKn0Ss9rBeOh6xTY5Gv7EDYq4yMXVDJfoVMxrbTfFAZhBAAJM0S
vi34p5/nLH/JDEIE9+Ix1drQ31ADiMFfC9Rvlp5bqBAfXta/ZDszvzxE4bvOrVup
pICKQEESlAboYmaFaerTGBCTcRZelQAEUIlGSnQaIs6jAE+PnKpsAXAdtWw3k10M
Iubor2P3OqkibQXfenfWnFcJr753gLADgVRkoPTAGwGqv3/AT2p9hH8yrCvTm9Qd
E5UL4htvCCb8Z9990fi6hDdUocLwsUMQShK6PlfSGknAPi6qp0a8/883/020lyC4
/wgfmfml13H6BhmavPynf8DS9/0kOpgIJNSO5MS4n2zxda8ybAmHPmdf/TOGstl2
rnoRqFPqjCx4eedtJgkbMkGgNQetHDsilz4WzxpxXJ3G7WjvVeQF0Spa6lHx7nS1
m9EIVSC3oMwaKV8Wbc8n8MtMbvQvTJADA07712MjRl1ih7onTpPEw6tqDTSZkIX3
WO8Q9B2LIt9t0VnmYeedCY2o0WstH7+k8E7cSRsIlhlcOwgQWUCq/cBuPEx0CtiB
Uc9FDdPsxmxL0ZgKCC1ZIBfKu0EJJrAsmk/jwOYKqfwchuQvxInclQQSDzQY/dPX
CI0lD0x/bm0UyAacn1RlxJqZ8Cf5ujxC+hrZB2g9w8jw2qt3AEjLj5yijeEHMiUI
+3qJETVAy7d0mUGUR7VKBCwxb84BZjP8PBa0f08RMC+VuGynfqFJssMq0prZSzFa
yrVY/0WJGjH5+4kslNcZhulQFfNNZn+xEX75w0r0eFW3mJ8NNqwHJlAfw9tAPAvq
CgU43gcSNIA6aT/iw2EKqqOIm/UVEK0p8CnmwYQr6nuBAz8L8lD3fdCtF0Y6N4QC
DoMj0dNuab977ESLW++TIMDeDGXAvHmWvgBhCx3M5zUARQjtJtU5X+MA1tQuKoRo
2N+d1KbHZYLwEKz41x3WeTf2I2Ar4F65UvQ2awUNUQJlu0CNsQNo9xeoAnqaF3mb
XIMWE6MmFf2t7hxolX2kFHtWvsxnmZLiyljCLWdFJPu/9gYlONgXISSjEp+XdeAq
p82UlqPe4S76lj9xF9i6Xw7To7EvUuqdsS6Y/ZkFiJmmeVLNnpsmrTXGF0xc5EkL
Abo2+ETUJG++LlsdN+E7tKSTJPLfipRklZvn9763Ny7uYdsd0DcLqnDr4Q14VD3+
/KBOFN2aZn0Zcp6jKvE4l7qVPumM6EN2FbDAsFVVG0fX/GLCzXtUPIdQ5z2lbLGp
Ro1FiJcqFxsKQmvLYbS9scNKeKQydZSG+CsLRzL176oA6ohP04+dIauGpgSoXj0z
awOrj5yKEA1bJQFTBugq4oTWYqvaHe2ANhYKZwKQfOEBaJveYdbtAXdrqkJcDhZr
gplPanfzx+UUw3mfnT7ctq4XSxAWoopLuROmnrBO0+GCQVBq7kYBPAE2QFRJNlXV
pMcQDmNF4UtG3ciCI8rF5Gji/8kGSkVSD0GNati+lqgPnFXfxxJNjI2msG/S/TVW
5+Nf3Eqjl0LlvPJVjZQKT5LIjGlB6SWmdWID8T2GjEjJvQNEfwMYoSG1YJ/rppGc
GHyuZQj2/1Ch90lCm9NFJ+qfYZG4ReW4MOK2VJG6xu59rXz5hCW5QkyfZSmrhiqy
PfphQMe6B0STSHZGTKAzSO179GxAV345JkiY5W/KuoklAJH79NhYGRjZfnmzhqzF
LtXqDHFHBJYu/C6a1GCHhsyCEIvtNYYW1wB+vqF77G72XFsDnT4t/UmPYaPPzwp0
jAcktSJxX+hjMx3gdRgcOONLXYGZc5xix4xLYbz8Ed80zUz0ZkpppFnVZLuAMgOI
l0Rnlhn2cs7EI5hxE5okmbzmPAGpxLe2Tvrgq03GVEbzdPVb/tM6Ob4SfFqO8iH1
o6kfc8e3a+XWIuBCzZV6hYRBurEoZU9+jHP+pADC9rxgmHzw42SjFfzucMrnDq8t
aAa8lRZ/wfjlUIc9tRxK+LJrYL3x5X/19CirxTE/CPnW/xBzg9vOvPi2xCnAGWGm
Qoa5T6TRjXiMcZJ7Z4XVeahaEkB9WkvnrPADWJ98icpjwEKkYSFOptj+bZYd+KZH
g0EAVl//Ynd2vzbZhhW0m1pl8HtymInQVG7zIiWNnN1UJLSS5y7V6a4vb1sSIi2/
Vyl2Zee+N88UNwwEbcgGy73IzOpJ2TsDSkrGhH12l9llfv0szZkGnAB1jGF82OFO
DvmNAgfeUCR7XcY1OIg3GApm6qxpWa/S4K4HHAXamgGrF3ZXYj4q/TrrTN7UgrMY
8G5MuO/3iBlIpdXqZaNO8z8kR5/CHjR5p3fh3NWPWdkos9wv3VV+mqpyMGCmC6O0
7Ryf03JBjwTDIk9u6cpYHzAEH+0kBYNOcwPnjhD2I5COsJzJhLN9scKch6fGBpj2
dKuVLvYYqLaVPuG0lr89C/iokAO5ZakpJB8MSPSexERmuHGaZSUInWJfWOagwj/W
7YatjrgA+EGMDEU3PHs37AstdnVCAumatuec5kBhHnDm7ptKD4p2Z+HW4fre0VSv
UIzoxDjK4Wz+ckWaJwIO3CKnlpZchlsVvOpd27BG6CeC7ZdI1D0jti0cRDXHr2dm
5PV6dNr70Z84fkd3Cgv8qVQuNQiuPAYZSrNrjab+htAL0HzyQGLLDTa9pMR57Zhb
U/PCOfdlyp44tBGhVYBMO6h6LvrxcteuvFhFP0xyoYjPfOd+QUpd+yupFD1CWWBO
GtKNeDChYqVmrN6mtnwacl0qfQOFN4RuMY1c+VSPfCza2hZuBBSoiJQ+IioaP2FS
brE28RtXERxaikGkptgH9/M1PnAE9IrbjX9GqUAs3KM6QUOqKaAvqwd88H/rgcRT
cbzzbG11k76e4BphTJTX7/eqo6awm0mqlm/xe72a+Bq/EsPdTR6IWojgzpAzhHgp
PKfB9jI4yFOp069C66reqqVYZoiwxTje36KxNnDNAM+lZvOhRUMENVTYLo/7Plt+
wQSC+sIZl/LBLCNBOGIO9F1pikg6cbyFKUHwPij5hZ7KQMB2lGFZth4hAVTWTghx
CV07WIiXA4BLh22y8TPZf02IG9sOf5ZWgYJr4xfnJd8RjrB9qYA7sVTx7/GPOidw
tcFVpYDlj80/H+Na37Upu8UpJ4QErHiB2Aozncv8774HRJXLDcKwW5S+Maitd1R/
1pAD7zw+1bWaDBSmq+sGbzIl9RGvqoKRvKi1Z6vJB+PD2UvBea/vqHLg/TEY62P5
bnx1H/bT03QszF0wDF8eC9GKP4LDnwGp+yeqatBFmdcoIgvPaBuJLXgZNLVNY7+v
aw25E7u0LLwBmMcpI5eaMCA4ytGWujPyd4+sGlzxlNqv/iK1jxTHfeY0yEWAPSYp
`protect END_PROTECTED
