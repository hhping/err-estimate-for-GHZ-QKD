`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
483Jz5G0xVyhrQ2MaY/7QjXgNS4m7/rXszbWtCIXN9J4+iFT/9jDFFFgT8AT1YFg
MPr0XCohcUfYKeXi/MxrPl1Lc6OhIG/zVN5KqrpkIpbFLqsFenAevQKbO+LgnmgW
QTwyg+XkkOuQp3KrFKy9PS7B0kDROSuIa/XpzYAVo/J7nmE42CAwIluOdV1U0vIb
q9FNrZwSo/9fE3L085irSORTxtBhAiVYxJWWc6XRlMsBzSuddON8nknuw3BnLAAR
/TvsxglbJdJj/TIl8ItLWwdv53ca3VP+Fy48OGocvqOwnik3Fta7fhMVfcBUv6hp
85FKoc4O53+/QmTqlpFou37wDQbKUjSughHi9DqPhcPWhfoWplTiYWPk2HstCLHK
RHu3CsGOKdBYethNQcII15Ht5HjedHrANx7K3lu0iv1Pl+MLxgy6+ERhG/nRG7uX
TtARuOu/RFev05jon4YwRw2V6hKrEIVWWT0QSpIXQdPSKSdgGj6AHxG00n6x1yVu
W3JSQOSPBP94o3dOSxt6To1vFZ7ynTQJEH1sr5FaEGiFbi7+DElEOeGVvcvL9L18
rL3fmaJUmBNbOQ1yzcHO4D0GbXgGQqx+LUgLKz0SupjyIn7ZAOekWgmbXNQQAXmZ
DrGVAZxcajjk/2kBUa0qSd6QaSopfU89sWHQofok76zQ2i+aHV78LVNbsAU67BQ/
6xTILxbAc3niVvk43aPryJApB8VQVIXUMBoteT0Ya980Tqmd5HrL9nBkrr5PI7Qk
qxnNr3leyhcWAj9vsGKupyJGmMTF8ALa6/Fr3jnkmLEuOXDeH4Vq9JaDjTyPiy7c
OYmN/WIRdsG9K0OypIJnrzDTwpxOU2Y6F1Q/RjtBbdhJRES4VXdaufjc9i4oA9It
V5dRsycKFE69YnQ7Os459QtJkHE8DJlyFC8qtLw1/pU/n1G1dR9b8u8j+vT0pxzq
tep2o5DCbEgx6XmA+b24bVn9PokU62Jg7jkkur/XW+6YuQlglL6F1FtswDzUIEiE
S7ibWNNdT3VNqp5P2AwkKMjxcMKSyXbvbjmyK83jtTHlkB1geixU3tQ+TXPW4iUk
JK2IOmfWjufshHns2Ebs8dXAtrOPHhlbaMZ3+hlG7aT8xBa68XJwPjUWaxvFgRlE
UeJCuGHGuHe6GMxVBaRqrR9hVb0VkfvHQ5shKlU+VNUeB6xm1aTZ/p+pjK9SYYsq
WZIq0mS9Hnx4G3YCRB43r6rIm2df7+MhMSJSY9XeQTUY9lbQuCqz2P8xn/QrtYKx
+q6hPs8KPadbT7GMOiUSbgyHX0Pj8Y14ywEa8TeBZscCkrsSsQd3aP6WSl1CIuzh
sYzQNb0+0MIBMRJ23GMRoXRYjIFju+lgm4pnymdW5+Ed/iT3RW9Am/lX8nzvNc+c
AvwN576vidUAqVyVYPVYezHNQL+TVRSuTOypU8JnfKRgrv02Mv+/pPClctKS3lRE
ohOcL0MxBhCf7I+6kMJ3NJhNkwoa7bk/o4S/El1HPCtCzpGNlzHCN4AZPIof/OtA
DZiELDVYwN+dLNDzVVg5MSoH8doAklk8GL2krOoVSsc=
`protect END_PROTECTED
