// log2_fun.v

// Generated using ACDS version 14.1 186 at 2018.06.14.16:23:11

`timescale 1 ps / 1 ps
module log2_fun (
		input  wire [23:0] a,      //      a.a
		input  wire        areset, // areset.reset
		input  wire        clk,    //    clk.clk
		input  wire [0:0]  en,     //     en.en
		output wire [23:0] q       //      q.q
	);

	log2_fun_altera_fp_functions_141_dehmhdi fp_functions_0 (
		.clk    (clk),    //    clk.clk
		.areset (areset), // areset.reset
		.en     (en),     //     en.en
		.a      (a),      //      a.a
		.q      (q)       //      q.q
	);

endmodule
