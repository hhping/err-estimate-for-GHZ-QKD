`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uNkSmLD02/5v8ennQ4u6WzBnoq54+TzIL7mdwnUpb4hCU8+XMd6y/5dWrhi0oQEI
MZAfQaU+jrfO3fq8TEjgkt3PoMNFW0LC0KNqtEv/z8B4Ue7bpZ5OlUdw9Zhw9T8T
MCwqvrKlIi9F/jRaf27UfJthXiPLNmiRUGnouGDrfaACZJD49v8365/OTH2nL52D
lrSVzf8yazCgH8F9mmNaOMRTe1NjWHmkcdcg/j1Jr3t+aMdnBY0ZluBVclDSesFf
Sp7S6g3OqnJmzkbhuhgO5YHiGNkXVAfip2tkDvQZbX+/oSdwtoQg7pMljHI5pPfM
/8plCqt4XBDo38IJicyvNMOBaP4NwR7W8fBPiNGTFwhWuEAhWJjXsIwmH6clmxGI
k/qYg4+DCd7GpDLZF5Rkx9VWVPOVAnhOMwLXMwQg0bs46kK4FbEbdkUu+167a25v
tN98gTLQeD3w5/ehCSoCW9nm9uAQZli7FEbtLPR3jCbb2lZbNfc+kUWFV/AF6F97
`protect END_PROTECTED
