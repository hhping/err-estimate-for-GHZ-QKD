`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4EuYmwNxOHyQaEN+XFZbnpYLAOtgKA56Wc1tqDgsKedwURXlbS82IkFQu1HGHZGx
AA4ubqX8m68US2pXr0bJSOMSo8cga3H683V+JOB5VEt49HLd1Gx5Wz8fmdE26FpZ
G+O+qJIkXVjpcqCIMJpr45FuxlTvPMCXMILXjso91h5rp2IfbdvFUQCHMXEAB0yl
3L3da+XjtszIDcnMxqwiC2L/ZXPA3SnFcuE9aidH9elO0yyv2/YCEDkL1ytBpaNh
ndigZslxsmYXPHE+Rqx/4WAa8USVWdVO3jSoohGKHfuadPjCLI1uTrk0iEhMEAXV
h755jClizWPmFBvAkWwHjoLIc4x+FIYVVfVuJCxrRG6KNHqjX2bvg8box0fTL7nG
mBq0RelKbj9Sz76dqsq+kqJogPyR61VAgwuj/R3OMpThUj3JXPi9hRBuE7KA5ARL
sUBOnVI0n7+K3cnAMvziuVd1zbWqgCNqL1Msz6BKTF8UmV2ljqb/e3PGKZrz+QRz
YpGJXCd62di6Q9Vtk3CahF+1u423j2SubQAcChRxYhB0m2DP7xneXvTvdv13WddW
zJjz9imnmVBoFoe5TZJJfunBhUKQHTbZ2beelTK5r2ElzvqzMtDqbA9DEeVWlUoL
0Jb+t60tXfWg7yhwKEzZYSsx1aaRNAO8bL3Aput9XAwH76UfIFr/Gfm0BWX9+8av
Er2z5eTMn3rzFOmBPzG6YA==
`protect END_PROTECTED
