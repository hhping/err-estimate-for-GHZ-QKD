`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GHwWRdl+L6kgx9uV4INWCIDm8QbuoU8Mu0rq88MmlwoQVu0DirDeQVjdEzPFVIYj
s2Qpqg7nitpRtI8KezzaHVI7EUSGX55G0Uv7sZ0W09BF+2vMHvufxDciDUwtuWH8
ewz31qxXdNo2x42aNxJDrQ/SfswJ1+VfCwsL90nFJXaQGStuxk+4gESMDTRdlQ4M
KEnnnTTquxxHLUs+RDxJtr/Pi7YRsv00dWEs699rx0Scb3t/M5N8gpNqdNM7fEBS
LjrFPe5kfKUuPBUPfKEwAQfSZ3oDWHYgYWB8/hfSj+GMIEDAsXfATct5ixK7GTiM
tUbGCAP3SP/BPIRIyKiT2quh4i5Rl7GnetgDg39+kpJ9l0Fm6QA3QX0wbvxTbvNj
a2Xx8rwTSIKrKabCDMPIMTQ33uixcwCiwU25e/LV1sWAoZIge6wSbG68A3KJMGXn
Lc/6T7yZ2NhTN6UKZPqN9jfoTUNxedbSLPR38nZy9zoyflU1/FTl7TxCgWjcjUEx
99d3T2jzRxToXvHpAajZ7vywcMJyo/5N3oF/sheGHor4ue5zYBqC0PRc1lmAPdjH
55dGFVjUb8byidQbkZw4mGzLuf3BQBPoUKIHLXZVFb9WULjq2keqHVv04KM4N/Vm
gyt8/zGLQPRUFA6M9H/5jVX/0+KYWeX1nqh2PznBTh8Dw8TshD68JN4vWs671xTh
6jhZMoQGDnREkphYHnfT/XnUjfsP36/vCDww/stlwipLtJzV8514qz7DsnnPSmuY
qdqfEesmm7s8tvg8vuCU6VgcFyyzqX5VTsQth4PhCVevOwMDosKKSAUJW1wZRiux
5fC5IGbpfVeIUVOkuzZUYSnLUb0wUPqcWG7QurdiXyO7XS9ROaY747Ytg1HEEjg5
c9BPRr4ypdA6W1xqw19p29tRiP+JOZ7eLi8rcP3RivXWhdHm0dsXWAFSbWFjtPtf
259ONroyJwWCtpi4Zt1iLpfir1RKNzKPTFz8vMUj6GJPsDyfWXwOppcW/daL4pNy
G2ZOcJVBXnJhGeW0fYOIEueUayTGKGo6eLblp03zu86q/j6P5aZ/RqIHD88MFRle
DfyAwn5LwLfP9eoPMxKFE0J31um2ddxnBzS4X0VHrlI12T2Wrp0vDEAHWxp8q7ig
XWGKj4d2HirQg97mxmFJMlC830M8CNJBgd//ND+31BFPYJJ4CHtgNePjyxdp8xoA
1aIMMkFUKjseQ5R7fcaEH9yUWrz9HlXofqxMUvZbcikfWdynsIBW42o88cgR9e52
jeS9/ya20lyp559kw+o8Gora9AfrqQNQ+QnJL1pout8f4gWNiRq9xpOzAl4Xvoxp
IDzq4yscIXf6+hRqB9G55IVA5Za76zaEzEqCHbgRw1/dg7F7nVL95qfW9VA6O6g0
RA5O/YOKXHCknXvqrHmfr6im5WexHZDaWrHNMGr1AahgMhIyqH62h2hw9i6tDbS7
zq6L+yxnTg6NtCDW3Cnz1d7zOpYlDQExDPSRcMyf4XkDsdfZaKSI1QZZ1FSxNv94
UjHtOEZGjbOG0L9kkR/YjN9DqDqMfBJCJQJQGyTw1WBnqcfFFhLmBKKTWHtT/0Rp
DbrA9LuZIjyZjdSizuJ1G4UnO/CIWoN+b22e8uF0iPW09OUMpeqFZg9SELZPf1kf
gz34UltOV1PqHSJuDl9jjip4dmrUPFgnO4+RL56MzHiDQfRcV7+29tfkPWkFVVhM
eZ7LpGGTFQabG8eJqUmfeA16dWFpugxF1A3lpEonlYnjY5FMXzI1DLjJ9rDW8ZnZ
UdZ7XOQSfrTbCkB93F1epNjk2ZApLSueRp5gQ5589tZfa4pJCQQIO6QxPi15xgkr
/8lvpYcF+P6Zu1bSGvT7Ens9altkleKqJ4yrGSHP26kNPZUUP7qszsPAcQJFzrjo
0/yEjTAxUrCfzm+235H3PRCf4URtdCLUxWKJDoIN7PU=
`protect END_PROTECTED
