`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ntq1ACTpW1gGhj/+5PVxEIyjBXjvVFnfJf6uKx4WiuwKtLJEBaTKIwofcdJPL9Ds
PWmj1sdyUbjLyw1/gWh7/D0fPS1xmSXZv9uiFfJNnZhDe80A75pX+Qw3ToUUV13T
E/CD0GiWIPxspv3fW0CCdORLFkWMH195+biRYizKxRemrW3THLxgy0pFuC/FNreg
2ZvR0a42NrZ7m68SVGnPrFW4RVHCgqCeM8/t8lTwRE/mx0+XL2cRFZZyxVjMJWaW
oVQ+7Vp7cKJkfh2aFhfFo3YEVN8ZTjaqPvOOb+OnSiizdTzUMui6pWL+NC6RS/cF
JKwFBC3DAd394cpHFTvS3DSbCUoGmB9UGJpsNSTTu4DmIzcztOdgt2HxttWcfcrX
Zww88w7aXwHJDG7kH3K/Yt357Nc8SSh4yQHcH9rHBdVxiNHR+RtkaFCctv8siz5m
5PBfsEdSr8Ldgjq2ELJHPpd6DfSxcpjpkTFkebONnizCKQzfMY9CDgoUqND67Gmq
I5aauJTr0Liz4I0u/pEpAMO5BdQV46G5Cu/rdY004lfhG/K4p5kcXzcY3lBbwMqF
hgjhb5lY7/2WFpeByvqjLTdGZ0q9sM77Hy2C0DQ+DM72SOJ26Y6e4gXhL0/u5CWx
IJojy72ARtZxeXhp3nVwx0qgN37faMcj+QfurPY5LwAP2m+RENzTbkyBvrS/r5uB
5Bk3nQEV4cJk4Xdr1xSG7/7tOl3YEbtXUfRnRvo+4/xaz3y+OjS0JUrQ+of306QE
vNl0h/WL89o/l4bPOxS0ZICMjpwxqRAkWEwa/O9jR/xWCTI45MpQa5VaVpyoC3Bd
mGqWsIIhMMHGHCVIwuYcFRYTM7hcRUZFX7BGfUgrjiIxqnWWWydSobjEMmLa8Ocy
d+vPmoocn6PdCF3zI6VmVW+7hP0KXbOmMombmSucpGf5uVTjGSBdqdLKUQ2V9jiM
l70b+76rzqUBju90n69Br1vFoQliYUBWGoE9opxIHkXa0Rlm9dqZrd7wtI1P2HSk
wZyU6JOXmOZaZhen2lPddt8MU4iUeWWi9xlQZIDmCZKN/osAVOEhNoAsgw3FD33s
twxjFubAr/ftUAZos6K6sK314zAQX9//NbPvmQjN3g6Yxu8twRajL1DZEbnKJ89m
9GLC+UCv0NEMzJkcMnrIMQ5bSINZpQET23EJw1GH2rLyeDpJZQhZyqHx1tIgA0eh
Q0q4NkiYH/F1ne3HjU4wE70st0eqIG5OMk8WmyO2VS59/KMQe/f8xycw0+9fxrAi
6xJcL6yjag2dPL7MUDmKiWbRntB52WKUqG78k/8BIhzhSWvRPPrROSoNkzgxjz8k
8/ix+Yd/Z9+9DBjd5J20csbVMeWkoflqWSb5ICZNkmIx6qHGGwU87el8qDh+zrJj
hFfyT+kpy2HB0RBGKNeI4JLE1UVww2gTf2D/+JgcLV5+QZzZX8LAa7d+dh0BllyE
DYFVM321QakCU3Zw3aW+jkYoMD2MDLxhsZ5QS4CmYqGOvtuHH55PxMcYE/Du+O0w
sMGxJqUw9Wn0ML8Eyqi/gJvTFdxl/dNLHHqAf66xcIz37wSCm6Kjzh/M7YhPkNP0
6HWiUIEutiPph7/VzZE7luDaTOAsQuXmz8Vocrp03EI0BoritC1042p4x4U0T5aO
W3qfEM3joLveH+f4vDx24zC57mJmp1FAZ6MoTnSbDPg=
`protect END_PROTECTED
