`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vs2fRUZ5xGvR8JyThlDvv6bJO3t6TMmOWJZUrrheU9982+Hq8rNyWGjxdebTyJCu
Tdf8MN4O2fCzinXLDd/LXpvk2zbw4VctTLaRsOSJGRc7b9WzLEsGU4ETzQEyLZDn
rFMkNbB4mToROZQgNuf/t4NyBgPUOCY6K8Kzh4/Uw4slSLluk2XLsAVR2ZlAmaJU
nHbNKVhcbeOVMvbGQs1uq3D48NAqtobyQWbmgBnQ5UqrDGS/y/D05OO+6g0nqrsz
MiKqc4WwwsdEPHRzDxGrSUy2Sqisn1Yh3vowgcizKJGjANb6JaVs5Jtnc31azrtr
/SfTUD2PJK0UZPHX7Th4/8mqAf2Czdapy/mFsw/L7UweVqsj8hILGk73xmR3GbKf
EUD8PYdbI3dulvf3ynBHp797QheMxavn1JsAsctDZP//ASpXb42EPRHVGZl/qKaP
ZJzW4s5/sGKGAfEYowe7Cw==
`protect END_PROTECTED
