`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Xaej4ZEhOgBymMG3qLKgvLLW9NkQjU538ttzsNkoTHpI52Ekz5JsiLVaMN4mUKS
Ok4MEcQff6tzkux3gNPWXfUuvjzE6MZFeVbipokamdYUllS8jnDD1lU/c3lvPqyX
8mbnsi0ZJsb3xxo6KMK9zhscGAeuBdnPnaRG5BgqCADCOAnP50VCNPnu1uI2PS0B
Dg0Uil09TJ2BrkxePThqloK5EDQ/dCLXPbI/fJl625vqfW5Sran9DKj4fit532Gu
2lPasBDrykOfUhL/pYwphqj2/j5YmVGeNPy6qSGgX5vwZuyU6Mcs3rsnpA1MKrqA
eLrhGuaw2Bq2qv8lww+cgPAsgFfLWJ5ZXsRln3DIcIDFwAo4c52V5W+9XJkeHcY4
5OOz7lKfEmF1yNtuUOSMRA==
`protect END_PROTECTED
