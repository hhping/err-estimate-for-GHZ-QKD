`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L6RkK7km7VMc/Bn4eYMGDVAyyUUOyLB2Irr0d1CLvxzEFTbiE8Ld8q0DD9+8pklv
yPRN/uygnmwU5i3UcXm7QyURxsiYOmguv4H9NXYPomSM7QXx38/pNY0Cbsu+9BsO
9efMxxUxNXTgb9I4gCKKOl/KMA1cMmw27oErYO1ssjswfN0Bff7Y6gr24Fd2EBsb
+v+iHtOLjlM76W+UA1+0PYnTImqV1PopVKUZ+MvaaLCnP0q/lsx05sTl0KYS6CCQ
T9hAImX9ok79TFlR0Pvnc72J+G4ChtdRZs9zQkyXJTst/7BayeG5TlboCc94wXrV
yAl7y+IJsH5zS0PlUZFmEpgW8zTj5+zQV1zp5BUxq2+0p6WBGa2floMGNAwS+0Ed
HJpKxrGUmEFBOGyWwjQA+ifbj5C8qO3rOEJxs7fdEPOFfTjCc9Ipck0pWqJjajhI
ZUqNwdHqP/VhjKRss+a+AtD9el2ne9iUImEtHUEBcvHGamcojJuRVIJ0XCN/Y5fD
HDEmXtGSchPr8TWrVCW3tiR2l/FbH23cx6oyg+0iDc1RlJvT75KNXA+/ejFhmze5
4c4fFF8XQvcmIEdnLLny5iv3q7dYWSrMGYDc6Gkvp1LPXagnPrMtOud6VZFLzjD/
nCtQHEPOkR4DW9KoiNeExLO5UZwAehI4hrQ1AHSf6z88QlMeZJ3BHoSHHWUlWzTt
5Mhr5b5kBJYMdAXAKlddaXvznEKV02FW+MJ8/Ah15PLgHn11pKBDmyp7lSBdwlt7
1Em6picmG3OTIEKedHPv7Ee+xfuA7JcAKUBuBoHDoTxZpNleE90knGWB1dWVuoOa
Fm+qu46s6774I0TZ3LFlNxr1kDC8UpI5RuNfAht7qOzjJ6K0/s/n5RlQXCMwgd5N
aP6rgSa33HLiqo38p4K7/gSQ/81SEQFacYglfctBrm70zwM+8RC2YwKx1cmo9QEc
JgHSvWSocUxDd1OBOlgYeDXhWykfbvIIAt0uaRx9OfRZvjIkiyfKs4SxIGkXKhbg
FwEqrOa8tfOEdcL8c5EZS+DY6PVdvjwZsnMjMoQEt2m3l3yeCxaenIQLJ1GcbzLQ
PiScZioXIBqQo5vJs8dnBM3yzZhfL1/haSGnrUrgl0dbskn8ZGX+uPxZMJIAjXSk
xApWiXXtola7xV0l5SNH7ZrGFFNM3i1JEa/KsRkLyh7ysozzIPhPMkOiFrOZsjQy
knP9R6yPnAvfFFt9z2ETgNd8iT5fkf/8nuNe9wfxBUhFFrHaoH0UxHiCPMi7r/6i
N5/tlN0CxY3unFmnLJcxQqChHaEMYP+Zoak3UyV1FKRnO2sWVBCtWV45VX49tA54
wLPo2zN9tELr7uaaKsbnZv212mMJmF7clIZxxtWgOebOEYgzsdexPok0IOVM5Fsx
GbMQfAdS1emDkDJ5NsYGnQ==
`protect END_PROTECTED
