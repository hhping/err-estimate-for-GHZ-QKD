`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JkH4RnXPOgNVqKlyM4RkQpalNE97B0FNdgtfxkl7S5+a+RnrBpnft0r9Rn1e0kWu
uk9doy/KhTe7yYi0G0ZFv9jwm106Iv7dAHoJmNkYts3XkQ0vp0FBX4v1++DNTEeI
XLJ+28UNDAGutDywnbQ62wfzOvdpAYr0cMTsoZ/k3wYGyrmSN7qQzO4FF5zZ/F3u
PI9CXuYed9k3fS8blVK+4rIvgrsi2Q2Kny9xSF8d59B3cMU8Ew/h4vy1qJljGLwx
lXQmPcXOHIO/rowvfWKvu143R0czLXAfo8C2MVVYRBIFGHSfvbl4xkwJClAEquq2
q4BguP1y40jIc68UBFmBqlEDyWqKXu8roPp+TSbiZIlxInXiXb8MOuapZPWOE+34
qUFQ05TEF+0GF1DA03ORWx+va/qdzgmIGxmgTLZQqJRItvYTxMDePC4Z1jhDCaLv
MeYTX+3nKWrmeUeMrLHb6Xy8qbk3bKLzicHOa72I0mRPloW1uj3EnU9Wxh4ZG+zt
6u9F52uCbsgnfWk5YPzaaceZ6+AMKr9t1FDH21Q9UbqWyab1g666Dzv2elt5jAWY
lHBvbqhHb8/1MqtxaIHrfW6I6ZHefOHOFbylw2vzY1+72FVWqrI6vVyBRIwvBeJf
tVFgJnbuB7f0iMR9CGGxSaOsYXfPSeC0hcEKpCrT/D49GN6+sq/XslfbvZ7Ci0yH
3hB4pq4PmoYUx+dyXDldFZQf0FJXlHi4+JLEqpzFRZLGXsmh5cdPJ4M8Ac7gN6j2
P/RJRTE0RXzU8MHRe+xmxouZe+uMPH9kD+sWDLHleKbCcy7axk0MbPDmVqlbfBme
0ZFd6jJtCaGvCuRHQfQ7dXrJq5+yLMMv6+clEJloNafW2sn6sp2gVZ+Mm2jWKf4K
X8N6D/5wP7q3MLwKzZPS8G4iuwdbEc2S5hNCP8rCZ4R+AiHhuuRgl0FrTHxIVPP2
FPQQK6mpEj/e8ER+EJKivdG/PHRotMr2DrSnOkJaghzVknKbiyu/luBl6FI0IViZ
QtdJOoPMuESWlEA7MH8om3kOu3Qk4rsaUnXHXM5MEytjPcmULzkvzBcAJTBERpI7
B/pOQE0mnCEanGnx1WL5nMbd1/CX5sMe6ED9DsEXdu7h07Cf03Zk6CsjjP7NzYyG
7xhBBAAYD6eJ7S6GbKY/z52XroiMqwZTePqitomiYg8Idt+0JMpMdUrHZ6yhwlFA
cNgj756PxCDD/8mivbtco9a9iDFoGEFtaMD6USAupBHci/MOylFsCmTnd2iaWO78
gNTiK0+Wa0cF3zsWuO+BTZSX/JbUUVBjA8ekLngaRhbAoubpL6Rhwlyzi1kcVamv
nxTs3ftk9v/Lwn6RpA0MSnZBDgwoDl95SyJu1yg+XL74hlYr34EI2pSWp4rqa2Dy
ExyeIt1P1IJKQRX17bgHSrl7eoFbUgrbM44MRIJR+gA3RnMxpil4iGDazixduzWF
2L5lg9rFX0ogFJQ+7TmkUXkqB5rtT1NocOK1tygcbTZM//eV1/brF6gthMXeuAG+
i4fFs6KrWu106PwH30DBHWLceBrpeHQmf4KUbQC+o1S76mZSvrtYeNPzCwQxyVFm
LbkxQ2U4c7UTDnOJX0qNgcW3TiSEjJ7uvQo5WRTBCuE6AfhyJiKpsn/7eId1zQ1p
56JaFzSpDsiqGqp7w7LDCwwyrkbiRK5cqNF6fVYjTwIvzJRhil14soQKHvOjnvZb
kulzUMXmK/CviqYeUx6wsTRbKDnmF6hjfiwZjbpTPnLk8VQbOaiETSNLytwyHKmo
3+GiHUU+rW4em0EfQWlgffCDBo2JPvr4LTZ/Fsq8fjkzoxHvtzy/4AgSHfjFyM56
9ksLmodSNyVoWggKn4lfcg4MQ7Q0cp6rndRk5054pWqfA9akkr/lcJD+MZL3H6kg
mGdA8qq6XEV82jQcxvDOelJzaTIQGRVp62itFnqi9bdSBt6xh27k0MkAOkFo+QHI
waCOuheJmbIAQR6XKJAR6DNdL/I1ug9nV00KQrdCCgHQOwwjx+PSiD7n+7F0oigE
pwbk4cA3Lnvd5LnKsbbgL+Lrnz533z1QnbEPQv1TPj6c+YT9RserxsiAcP/aIEup
Vjctbygic9+nL8zhglemAJbLAXNXtquYS+ToE6EV6sdi0PcJ0NOEEbYFv6qSV9u2
`protect END_PROTECTED
