`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fA14coIRuOOgL1gNZ89iMis7SEuaKTkGcbOzYu4fb3wU1CGy1K4UYY3BV1AsADqh
VSmUynKFoRq98dY2Hlkb3e8LxvtqIfa0tbhiqLosHiLrdhpUwypS8XMPHvk0Ehmq
qPBchYivsys3EvdbGZmsOEyvI6Wglr8ZejfP6yiN8LmeNdC1u9O8+w24UKXdLOKL
2h6aD5BvMF0HeFPspUXB4Z1G+nPBJeWPzpj0EQVhZT92EMtpMUhQh9HWTBSo5hqw
5Xw1GemkARNJmCmHRQH6F/bOi82Ny1/aUOLD4J++Y8XVTXopnCaWVi5mgnvzXx6s
V6unZid4zXcFPcsIDEC7db5ctWCgcl9FdOa4uNYYwaGdP4q3v4WfOLSDdKcobGuN
+IgOan8mYdvHpoATTZ9Q3mJkB0OH9k34XuHA3z2+OWPYRO/D46aDAHYxL6U1MuUO
El0/shC9pMS9VJ04aHif1xz2Ygf/VrFoK373/7pBtuAvfXFbV4wP829nlN3+Upo1
wymRC0yUXK2X1IKpA75AsHkTd5ZvupVgautpV+wU9Ms7GkNSmekOQBPod4grQB2r
ybCs33P2gA9iYIHJKQKu4i3L4BLaV7JrLdLlAPk9PQzxsUOkJgDo1wWA6v6uRBRb
99IHMqvmgvs8XPSJRYwPHRsAVTZTJWz0SsDlcpbddH/dW5LWmxLL901hNjj5kfpT
EnlXxBv0rIe35DFh8HMOlyrdULEKOfeIR05DG8OIfX0ZE5tASahI788LhlTYIPW8
VsQQFkt9Qy7w4+nzAflawWd7N+YCUPKV6OwhAQg4/5ALXLZcFksvS9D8KoxCEzZL
XNaVtlwq1ba7QG9nciznefMEBZz2o9PkGioBGtu2VxEfTmHKE8Z9N8ZD/bLzlDG6
RNxl3Lu9QyJWbjuyQ0PbZrWqoWsMKQUWSdGIax0S/EvuzGbTurzAyfhp3uylDck4
UFuFE6CR4JoyNu5LCeH9EL22Wq6A9PrBsV+AOkEG3NjnUq3hjrbVVD+ABunF6f41
P3wP9M0o9ipPhfPDcgstoKgRwG/+X8k3mJ4N5We77ONIjbdTYOXWubFBudLy8pHh
uVFeyeEhueX2EXllLvOzdVdCF8kSgvF1OlXUJYsjKQtcrR/GB3XA7XeYubwIK6to
yl1jGBDyHGZ59F0RBvpERR7DAA6Y8yNilJ9WBSsUTi8T0hb0KjgH4zf/7cufbNOp
BWxbf1EKUua/mFnlJxqHKtco+rYtPD/6wLOlUL1bZO1CFO7B4IYM1I6WDdaA+Ks9
jf86D02At6zxIUOHiUYc35ccO1DqLzphCCRQBX5HzX5EzAeXoTqu2+2PjDIjRxBf
rdTdsLRT9KBHQlYvo6u+QjSeKqFImbytr8NtiKZmgohK7rk2uXn3/vRP/Er+i/Kn
zTPxLcPN1LxnHQDpeE0Nj3V4rHqhuseuWkqgRG/cXvm/VDlWlxPk+Ul+qVtrD9Pt
cPw5t3rhcGw/LauJTfBW0KphOTYJXGqlsK3FVMolk8VB0zQmo2BDV64G3tGiPIKi
9O4eLyhWZTxM0lR3j4kMv3rJT3bTGYzEZWKOLoBKAobaKxNtWL3K5+m8wYtFgYkE
shfHYqInoY+V9jvUjc7lA051I7DE2TK4x0CH3KWdtnhsU7onM2WyDEcvA2+bNPgJ
9nFygNMLY3oYpUnWPwd9bJvD3H0C8L78XggSiP4VvRHf+hAxwxSAwoCd5pe+8/XG
cEaG+GfuwhoZJSEgvt+w0ztjemCqCG6FXo0M/ZTl20K5Hrev3MPrQ4HGzzfnLNpr
44yNhqVhDjJ+O0ezh0F2yIP23Qh0gbDft3IKOu9MqgzLxSXkHM4kF7iBPBssODKQ
ZDcQeRs6e/GExBxEAb0aFL66Ye0kJyJ/E53ThyEO7y1BLYPYCF3HZDI79uF0YxPE
qubK5Z6XfX/BLkYMBxwvNcifCWCIZYjKI1zGxHv0rvjll3xJiD59FDOWnacGtvwO
8pjDNbrluG426lLBKKQtyEQEKTn68Vr7fiytUbxom9aaoXKponL4brWSx8rqjoMU
U7oZ/IWRsfwicV76ImKgOn+Kk69YxeOmy5HLxiyCQGl/ooGx1lOsoIDSVPM5aF6Z
ox4IP6LWw4LrjIGQ14gLadvoUGFnQQDKLqGWP9UcMA+sH9tQg381vBmuqrSpLBjO
2zWrXYgTnmQxhVaZ3Us/ZLFW9Sz1mOb+DTiZm7F3h6s/gn8V1SHl8n4VxcuJW+Iq
tWOYnM4ucy9XubUJQwTHYyYsC8hlJY60JEuyPTbzn3fLDDiH7jXfr0IKmhLtiHyH
VUmlbanBLMvtYMPP4+jfYhGT5ECpQ7tZWt51PASL5N744TD+zEJI+/8L267mUNgE
WiDxuXF+EI0t2P51KrGWXRRtVp/i19GZuHhZPLCs8AaXCC53pZgF0YHqIaj9ytSa
pigVLIT8qRNrv2EDgqLhI96Os/HwBbQySSDx7gI6ZCNNxrrysBahrOSgWG0FOBxm
mAf+kBF1T5mZamCKoWNsMz4Teo+oavk9l2GzYqVDKCU9ACFuvYAvCx95TcfY2KV+
eX1+H0W0tccJ7mXcrlNCPFSYhvI1LgLocSg5Dy5xEggUoniwFyyXuvGb5w78fN7G
7KIEAKnERvifkVuwWnzC269BT6qXT9YWpmpvK2GUbTv9O88xqtxH9LIlsHgIWCi4
tjkUL8dHbjHZ4tUHusLt0IAQcaitw1Vd06HRtJsFkcMrc5ZP+9aPVm7E99Si+AKg
aeMB2AqM3M/jr5Jpmyx78/dIegpQkLIj5C8pwIpGO5DCUO433MFq3rATyhbssyPP
7pKDmBnW/pIG3/dghcIssThJ5uPVMBnSEHwEpCyzpCr7fwXaMY938m0NAKp5p/W9
AtkfAjmYMWXWYr03JwHgpauM87H+yUxqqHiWs7xg6Hr7ufeLE78eFQK/kEGenOQZ
ScAdFIE9b5pxN0iAD17pH+IgOYXxe1/XnliWNFgAZ1z5ACbFDnm2nduhnf4wbJ91
YBxPzyunXMLH4id+/JXI8vhG47tBZO9isINqNqp5r8ayCwmXfoFNW3J4clfg/tzy
0Y2QVb/y8ZjEJxT3mukdO4QFqeDbrr2LYZF41ZOn6KgkA1JDuoEkk0MC19A2rGbj
DjVWgkY17ku0SFe5V65rTcr+OtttpycYirEXYwaZjlyvrk0l23IT+HStwkESoRp+
QPFZgA9sS6GgAQ1LabQgdJ8qLJD5aH4c0dZiroBky5q1j0Lym5/19p3e3JzEGjSI
sx8hAOJsZENdseF2nsrEnM5O1C+jxuyLlNOE2I3CB1Sy7FRnQkDGTeoiGRVkZlio
yXGMTBMk6ZIw1nc8NzVDKWXWaILPIaoW2nXvHw0grTjL3uV7wlJQA4uXML7JoWpY
JRpS0ql64YatZOW9T0hUGrjh2SilvFKhi8Ze+srOCvYzD+NQDEUrEJueBAQLulV0
crK546fV+tlEA5NO8fNhI4I2rKk+/m0nEdm2w5IL53NIfFHOvKP26ac0U9FxSHpo
IFygC9T90KTPj2nBGIaOU2rzTrrG/wml6HNG8UyRo/EDdYvUy+dkrAHNgec0o2QL
T5gFHlSEsqSOaFZaRZOXEOEGAIOHXXI/E6uzdlYYxil3K5qS618yb9Xk9olMJcfw
GYb6rvzKVCJSnGaIonGyUoHpJEDOpMSPGOlXszuU9gbOer72AogPLEbSiovPCHc4
wyRL6Ek6QKboIHPPAWSllPdzyuTaG0QqSl+2G7XqMI1JoepIf1nK7DYUrEOfohs6
9o5wiR0nbDPccDYzVipcgaQTkWQozGQ+Zml4/aqPP9f1gs2dUzG57o8GlRVr2lUe
o87cdH2i+X6ZBrocImb3Ffg1xEx0rAWZvAEC1ezL/cb+8cIV1hJADAUmAiK4xixW
x1LaCmYnwbm7ChhYU8xaK8R1u28fGSoCW37vGgTjMUofV1tGwZ6OPZuX0qbWUAkw
NgY1Hq5gda3FoAc72gpNzQm10s3uZwsU2nVK4InisLUlmaBCrxi1Wu0zx0yyL/dN
mA2/Bgb3AnQydJRt5Dm72EKsQgUfDr9CCPaKUQQEwjOakkqnyVqFcbvZ7I3BFKKc
XxR5CE/xML53lQeT7hcgU7oOtUjO+iWpjHt6kvHAeoOoAfpu1Hjd7KZ0amQQUMSc
wPdsQ87fo6QXqwinElkRclxYCV/zU66N8IVsfr9z3lraTRuQ9n8EaibPfHz9N3N0
FKHv/ECGcBCcYTX1WJbc1LNadJgl5TC6UxPMyEk2kBINLnPCz6/kf3F2nsZ50Yr3
HO/nCQOxQ1SoC9Z7hSbKxxWEZwIboB/Fauv2S659IQOKlXmgD63XKUMHH4FI12GS
HLsLEeYVhjz/Xhee3XAUov9cGlYVjahdCOzipeFtJghvCwiklSPObVbj6IqqXO7B
XKrVJtNlRBBU977mmFy71iMUgHRIQHjOSONL6J3OeZDpQQoVbxkWgviLZCSOLFiy
QoKeUPp+cX8ypFq7fTg4s0BjGEm7x7i75abhTTAowFF5+hB5YraolhAGuQbRlqFA
07xR+HM7cuLLyMpWjXg1/xpM5syW0qpSMRWgPtmCU8rQ+fEHRJfQe7yY4Zjl6bwf
QQkPgF9A7EnQw2WUI+3s68BYnT77lR/YZz8rGCpBPcdwN/Zqkdi7tl2usddV+cLl
vaPmtH+QcPC5Wn9CjT0p2hKBLtWeIIuhOraM9Fs6sMugS3MzV7XvPaGJFR1grrZs
/AuQvHUEclGMi4pYxLad3YqMET3LHztNY16M1p5Hpx0O8SFn7s+NHm3QT/IDZj2w
fSIAsOeT3MXjnPWJjrYcQrRRiXGq0t6PCZTqWcQBuf7kmEA+nzxo3R8+vcEz8q9w
VSUaKoXpHPuSPb7uqcm0EJA58Y+hFR/9atE8yQmGgKdTC79AOdruCW2vXWZZ80gk
uJ88K610JhnetAEWocAQFVi0byXUcdYS2r1/c7lZHCw1L73BknR2ODdnrN5Ds4FV
DQuoGAFQWTTYu5vMxMHS3bc3phEOzNk4H2fv+S+VdNp7h1kHNVi2i4u++Ed89P4o
w5f0OqYiWoJhRTlxfSdmohoASa3qx8qXt8VpyCjxneEsyndi1J0X6HzfoWdkoz6e
UN/RlkOb98oFko7UvM4kfberdxIvid58sy3ohCRYYbLFE3EjzF4uCYcgWpe/VLIk
WhTnAH0KPyplo6mLVDy7njrTuDLbdjh8FskttMx3xjuO7IkWg77sajzsSYa1mT4d
MWQHWf6jPjQe8RBvOFqwZyC2R7h9TC+aFC/oD43qVeIRgtI5PRYjTqrFYQ0SOrro
f+3GDLvb/Vj8aFtCD2D3bdYjD23VHJhE3RDnWpdaIb/ttdrmw+Egb6ItaSvLNiMx
15JGfMbCHbZvO7DKWGNQCeNmTSJDBySVYlqsc000wFiDk357E45861c0ZFCJOh+Z
`protect END_PROTECTED
