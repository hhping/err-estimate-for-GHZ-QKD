`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iZfnsFYfyH5cO2LTXTUw7oXYWJCD08JlcljxZU6diJ6fgelt5KKBnCVXMwHKwpfP
o40eG1kdr9O8NpA5eWBeF/vBF4QVUAdxjAuNLWo2DHhzM9KVTuXax/NoVKqe4m9+
tF4g+z+8hRorZr8TShY2KpuflYbMoOvTo8DgYTTiASitScN6VRX9vO+TqEmss5ov
fUZ2+/M1whunlnojV+VUZQzDr6aJj/DA33q6hKUA66ZTYh36MvJq2N4RfwUJdWJz
LYPScstvNofGccehpYJIBSy3TmOh0fr87o2SnC+y0EdHcIuxLAAXu5LrDa/xGbz6
hXlI44I1LDgYmzqwnA7MjsE7hROilS8PU46jqwc6Rsp/GjupZFu9p8NbdGwUzGlX
3ufgu+JL+B2mdo7zavbP8u/IMwnKqSFL1lKtjMxIYQYVDWvdozU8GblwcYca3Zdh
Qn8bcdO8RqOHIh1IwICryvxC7XrAB+rDpHsC/iTTsjbg57NCMPipDsP20B5/7BqM
h9qtPyIAmH0NSh3ukaCc/lQWRKZjZK/keP+bMzfuqRQlDYmA8wA87SsqM6/QnD0X
sZopYpNTt6ZB2k1Wf92S+zO+COMfiVkvG2Diczj0lVtk3ZGuT2C7ieUVUcDA2RdX
U4/muVNlmI9t+oc08tA5DuHe071gMkS9N7b64XEGz/N71LrQkP3KuhZDGSWcEDKv
dOrPbuRba1oWFS/siWcpbmMrZ9FuPZR+1PWCFSvrvxSc3xZNDL6emovXoLTtOCqS
vvBdM7vHX/UJOsibks2LMouSQT61MzdhDheS2Ini7fATyMEkeG0JS4pVqZPA3yrS
LNU0LDte4QS0thcw2QDve7LhZO2pL2P6L564yvVmi2Dof+f4AsyJfiNa7odwOQym
aPpQ3GHTmhbLzBgve4qioqc9wP+a1go6j87l8BpP2cGiyj74ksJtD3KMQM2Z//oa
efneAe5aAsvh0OHiQTD1vPEGmocZ8BEsLQFAFDLjxg8m27uFjeTH0Vjm6q6i4yFu
8jUWUGLSFLko084Yq9Br7oQrGph4982dCv90L07QLR+tgv60jkf3icGCKfIstBpO
rcY6pi6K4s1XwvxR2kNj1VBTUplo+DQwzIp69wm3Y18rXLM/fyu0DF76+7IoeGBN
pb8rvNo6OSUSiseSFa8qU8m3VShUw8Cfsn9xIHOtAJ1LnESkGgyIpJCmP0uZBnto
AfcwxWwJGeruelhJeK7mEVTwbBCugImgoCiQ/eijxYNGGJ8L0nCpk8fdQwAzWTfb
51664oKFGsBZgpSycONOw/zxLnCsfF0y5/29JCCYORBaHVVyjxYa8crHztckKzTV
xPz68K3vf+Lq/FroBIwkbw==
`protect END_PROTECTED
