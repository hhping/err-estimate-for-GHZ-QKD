`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C/UTtjg7WJhXYl3xqgYWpAeeE7l6J0fUK0t8nqxWJG9oiNY5aRTz2GxsUKRGtbXr
jmHgYS7toSX2m76qR4HXmW6FVzv3PzI0eB0+z0wt0L+4ZrM7VWvzuN6hJji3F1tj
5mfySSNUsalkS0VPUqtiMBaxpJvlHYuIyAPC8eCUXx8zQJ2f5Bo7Jn1u+2HrGBe2
Igbjwicuu67cHO0Goe1dNzpwWWWGQp2zdFnBL3bWyLzamjDIRmyuJG9xy7kVogLu
eV+GtGZr9n27Q+oSKousn8MPXsavHtwKExvc+pgbHzryjYG3hB76mKziVvbpKfqQ
WudrGa8KwDgHRjywj4yealBJtyPHCVvOs9pZ0SIZij5nmBbRjUtE8gH3G6PYpUA1
U5aQQqeRERH8iXlQ2ZofOo0XzdoOJBJdjHB5WOEvCmyONxmq/mZVTgDP10W2mCKu
3qEYvtzjLsiEXG61OgKA9Ohc10LNNXsiFU/OELE16nQPaGdI9anLqWkCSZltHSE2
TA+7S981iZ2PRaJj8y58yxRVHRleUYKs5FoZvzAdsn9UXM1E28qkQ1WJ60BR9oyp
l5fQ19xuXx8kuTtoZTTCT/u7KaTASL2aUwPJCNflILlIRI0RK+E53EoR9FDXzauv
kxd3ykOxqPqgJ9Gk3Yr5ImeYfHcW2ZJxI5vpuls7e7O5mSEioWHugbMbsqcGfsr1
z3cck2v91eDqjHvYKo+Uuq0ZjjmxSbYET1AbaZ87Deo=
`protect END_PROTECTED
