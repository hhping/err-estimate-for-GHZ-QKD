`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PJ6YvCstZ1qzQ8itKQXSm7EP0+c5lQsl1FdcBEF/1VU7cnB4r5mk99ss2Q6ZqdNF
RdfdW0ulLYodoNUNbR7qb3p5siqW9anFbXnZMo34eNrlpcL51gF9sTPknnQSHmxl
oRq3PLJct4CNE3P0xUkdR5Vb2B002eH3j8zg95IkeU4o5FF7TRzk2O82doZFDow5
oWpetbV2KreTRJHDNzr9mOwxc5Pu1k5968B5biJyNLkwHf8FGk4ap/ueymXq6yyp
86BW7/ZGjth3xYRnd1DEXqI5JiqHFrZRlhInAQeMGuyl2PRQnV09gRY1eqH2OP3r
O+gUpPlKAw8NQJM+07Xy3pdZdD25/oJC8RsNCncNuvKpZ7pwS7xT/D3RcQ6ybPOR
omhrkOidL8+Ml+JMjGyxy78+tbxETRgu5hMMILbY/x6MZyisMertA7VnpMOBdCnX
I6OxRWgvImyqpPEFyKrUWJSIuwiBJ2an9lC1bN3znYERSZGKWOQ4ef5bq0EkOlhB
WueU3HNw1ss7oBQ5VFAmz+uKcMEooV6kpKppLLMiNq2KpOE1W4EEf3aJa0ZRnil4
f0tn2umIU5Msy3gWC9Ak7GSC3zOhDHBm6EvvKuaEpR0aId2UnHodXAegDLuPu+J/
J6IfAOfZJEMphEat2bn+lG9uBd1wtK3LKIshT6vEQ1Yb8y4gSIr6q0j9griugvEF
IWOHyvqgNpRIer1uBcCG6ydXEvc0qpPSP80oKeI7+dZXX4cXylcNHS19iZxZIgz5
r5iRLAvyieGbdm40IHPlAgX5AWMwfImZ1lRY5UPw1ViLoMlb8wHlPuKSXD84Ixzt
xuJ+ZZjNstMvrulV4OxZUAn8k8meGo3qLkyMm5XK8/s=
`protect END_PROTECTED
