`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fh10jcVvDIRe1h1UibXqnPQSSYLTrR2D4zMu2HoetpXwJwfe+oGyKvErW7tQ6E3q
z07wTAqrSy+PbAjVGP+snp9qutLaqwIUa3TdMHuY72LD7LpLHKJUrnUW97+QzodD
1852ofeSuM5OoF8Zm9HQ2fEY5mW8HlASby83V9NCUYAqxWot9WIIL5joWxRxjgtB
ismlPll6PyPSQ30DZTa89Stz1OEOaKgthewEIfyaClIwTm3fmVzJcOx9ZjkKc2/Z
Gu1zGDFXSHA+CDthtalhHhwwPtpApU/qnHiTQdLrFv5dGYHcJpD8az3JW7Cx73iw
02+nOYgKJSeZ6hAEkHdKheJHUju/DpJXMODnoFxHgcXVFnUQLGd1GngSMoCBL6M9
4SyJ9CQw7UCgbDKdLoERAw==
`protect END_PROTECTED
