`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q27PGRw417P0GrzFon7kijEMr/s3VTbEZQjyuDuu6AsceJS+fHR0+4Zv0nL57qDk
6Kt8Pky96T6I6Dhu58Pk/VZl4eONtUJby3Ak6PasGLDBRNhXPHxaqsX19mg3QO5Y
4QLe/+uB02cspVkYvrYaoXqS1HoQ1BzWi/WhEPgQG+hCqlcUkhachEol6LEb5HPV
1TGIriXrfiUE9i6OwD32AH2afT1Rxo9Xpz2OBfYw0TUIGlJSXZ6C5FGn5RB1ihS0
JIvbnzw0dGUIXegxfyn9pg+/w2e7nPABv0/SLrezje4AmNsErm88QowKfSjFw3sA
g8wqd2UdFNT52jBVkQaM83p+dmmU5QvkANHHTWFPt3KJppuWcwBSbgHDcD3QFZ3E
VtHHtAPvxRT6K77n21jpgKUg3aLzB9Vqd25e2PFoG9Iy1/s7G591MB2U+fL+tiYi
vx2OwSfeKoGTjhXJ9QTGA/wTUojFh4w1+KvADnDxjcZW2c93/5RlWQNxjugUptez
tATm0HoToBv2NBOk8sPkxw5RRUCSnlhyR9WJyPK4xP3lmDMiCYKmgn6ys3S6UGaj
99mQr2dnUs8mX3cqu22oQE7JHHooSyNUEoDtEYOOvuoN4y4dmC65SdsgsGaqTBXW
HWrmz9KnXubu1hZfgLxxiSq7M5oMwSoUfi/pJvH/mLd++zME8ngdERlMqK65D2/2
udqou5WBaFgAHBT2XIGmWVQLDvg2aAuysKy1rDRJ5oDoYuOfnCWicIDum2Uhghoh
oFtIfcS2udUsoxK2TGNfVmSyMoXlkznxJWZASbavpJbq1IVuNL6LPZOsonNqQpYi
z+NOkljbOe4LLi0ty3ix4ocjWgTAxGFfeUeChitntZwwkzjEr/9Y5DQA93vH4esV
XgKiK0fGt2urHfKq8oYFLAH5vB0zfx6IIfL1EOonrWYMxpHjLA51/REZVJnhspiu
Q41XbKUk/2DSsm7y13W88njcEn3t5oHEgUGeiBHq9Pqv8UKXUeDCQmxgEungrgmy
LDrg8ZkJbKtN9DgR3aRJoTgLH9tYX2erR9Zs0IbdhirwZo59L+yo3uSTfPuQ/pUW
8No5oqts5NoK3LRphg3QWJ99IpBze6N6WYenljKU972XQZwYi3dE74+/r2/yAlFg
VanPtgmmDLAB8G3ghXzTiQhWvmxYkDK922l2sijYdrK7MFX2xthyVApMRRpK6miH
XCV4lBjq5V8AV0dENpf2E2kh5122/W3PXlYvvtuUkmO/lB93Y+MZyPBKCFms/fj3
Z0cCHdwIey4D8zimHrv9a26A7BeXlZ10azkOILsKWE9I0XFtP3WnjIqaT5HM4GzE
i8Rf+NH+hj3TqE/+aNligAb5qRVyzIWWppHfx+G3R0TuSc2zrgNKbkec7szpxFpV
URtkAZIctBmGbuIVy+r7BThKxlA1kcKxmDiaXchxiZROvKtwJUcYZZr2BwSMbG4k
h6RExqsAwRXfEaRO+KDsKIvRNFodhyh3NURWu7Rqx/GaztEIlfab/fUNmU50+W0b
u3s4+Ba15tHdA5xnARZ7z/lcDQhd6lVNEOt+8ZoS2aQu30S8mkmrcrUsLiYNcYVt
z6DZ0rubT8tIqVlSR0AagtVwD3nCWi1d2RFTah96m3M3zTBkDmwuvTf8h6oBdD6N
DEicGhQBjMiQq6V0rvx4q3MRejWttNmzk9h/kmJN75j2xAmk4Z7fapCYEb2LkSzH
XyOZNSrGPvXoC5yzSpo7YIucAv0E9DSuiW4OKqsl/r1eIyIyHcU9Bf3xuLT+1e3L
SVuu+5so7fK07/yHTRROtzd3sZSLjchiq+p9YssbiHtMyd+nEbdY81iNIFkhx9gr
GQXAUW5EsP6actmJWHbHr9FLZkPeqAouVZGvvHigbkVEBdgHBzgFRi64bhTtWD8F
MH6TbCkHTep2RRbjqqtXTF9GClHU9C+ZYacpAp+52Sxxg0WollWV1rNUuPyfIQfZ
OiIxmWBa+VbtJPCpCOg+fNmR+291BMyArlKN9dcE/uX13PAF/O+boTfjqPNlsxB8
A9YA3LGrPH2x2KtJcc2TS2ajkcLkIpHC3FOh5lsLdBIbP62h51J4j78TM5aCDjq1
4UHC6fnKsFraGugJlrXHBQw9vQSMif0p+Y5U0NU6x9JePFa+0CKZEXxAp117wW2L
7o+mxjdjy4UPzg/0JkcIco0dPLbi/UTv4yazLrDvOV1SIhJYVnm0qYUv735difiR
Ih7HavA2tzJtRCqWpSWCS/Tw6pAedPm4LlZPpa8ywAe5rcSxTNtQEZZzVSbTlh8d
17+LHWJoTsSdCebPYHJ7ESTRPPjdWfxX4dTrALbKLwmVMU5nDwHGqKYbgvIMp2jX
sqouJIkOdl1G5DR7AZ917SqtztQgjfUaeZpW2+1wFdnvRFToZxQYaa7oVFohPQdZ
8uR0Ii2PgRQ72pKT7VmnedzyCp32SsPqJRg880dy5b8Tm0RV4fjEON870Y6KP372
xn/ANLtRLj26xsW1+L5Z4ospayZz2EGx7uXeHqXkT6LneWVsxR4ilNVaZB1BEKd5
fzV54VMBW9mVq+yat2tgT9uYzl4l07l9M/hoCxFPesbmvX3T8LViHU3Yg/57azoO
OyTLlqFF+ddkZwgBnRlQKIvKV7uCO3k+/G8a2E/3tW5QlohohyFTC2rgozMZm1j0
/1i15Olpm7W0b5OBfwTLSafrkMqYTrqeQNn5fvoCPkA=
`protect END_PROTECTED
