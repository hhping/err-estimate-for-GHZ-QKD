`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6g6rqbkCDUMGYUox88GTZYNB+/SACjF7leSgZ3nVrYQg0PuR3pH5IO0tU50ThUJI
UvVD8W8u2dOdUG2eOHF8wgTdXRMzXUcm5Vt930qZ1JcrpJ8eH8LzF0nCGPbefbzk
jUfnhCdRX7Sxid0ijWTLsTq5ynj7m8ysGarOJOAkQE0Sofnh5v4vbO4MTcnNC6wC
/Nfe78Ls9hHJO5UTmHNAK3wUUzpw+io7EvFQGUnk1X5Qvz4+TRFf+f3bk0Ug/G8k
RThi0kwH4g/GJhWEmHvnE0nMpDs6NPfU+AM43sky8HalBFun1WFs/3XMCo3O71XP
l3FOsn211uXT1e9x02Gh4lSAicgam7kjsO9P1F/OsDWLq1+XnnZAjAZTo76E7gPT
omxDGK93nbn38kaNZmeKhMaxctvYN0FdECftrLq5V8RT5x9wP53O0Z4q8nwr4/VB
riqb4VubOkJ/Ha75rgzUApHfpLDuTvnPNLWG6NAmv9iVafuVAgIKq3YGOCpasXcG
JfrmpC/yqIf4azrSV8K+2Q==
`protect END_PROTECTED
