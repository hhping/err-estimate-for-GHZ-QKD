`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IFYDLjZyR33///t7NTX3pEz8enoEm2bY0GruoZ5+7BQv6OWAAAD9nctkdpun/40I
ALAFB43J1IMh4kPAG04pgDskKYLqQdyt4P5Y1jf8Mnq8GM2bw/D0OZLCUOQPELAj
/MFBJvwtW0j3JGJsISr6gA3NnF9nphlI1HM5t3qhOs74ZqVWw+L4cKEhnQhYDcdM
k4Wy8gzdyJstd8bSTzGRPAyBm7p6co+Bu5LwhEtKGobxygfp0+yKaeb5JiSJ9p0x
OrjjAh4I6iSM75K2lQe4FUTutxtLuh84HrmECMEaod7NTJMC1Nxgz3nvl47o/r/J
RqK9SqeO9QWc86EdVnTYjo3nX1rkC/zOwJY5g+3oRTMJjP4Z3JSmn3zfMqVGJWpV
kqGO2MR7Y0Pn981MGKM4ShZkiHU+EyrRm/3nM8wAMcxTGNWppI/bqgEkLo+ruTkm
aooXcaMmcygHgiO8ikEKuGonJdSYRkU5oh42en4kwn/dKU3b+uIa7Cm6uLIGuAdJ
xkNibJO+kWXPusblr3xA8WMiAr70Qlb5y6f7XUOE7fcDvYkEIRIbeGitu/NhVyt1
vHOUlAVai8wpz2DXehN/iqgtyH02EDQmTstelUQwPr+yyVpvPWWumopHi88yZT2k
Zzs7UM/bYZN2cwaPp2PInMxWCGbO7n5odfgFpBH6Z4ohtqwrjFlNnp1mVYei+LZ1
ZWKcKPmI7SQOi0UJVvUrqBtnGZfsPs9KbjTqfIUAVrw+jKBtVSEHTDxwtlHn7LRR
GkdYlIsXU6crMA1HWP1RtMGo+CdWFHnzqXuDI+qQSAxDfPEKavq7neMjElM1rYDz
GMX2Ysbn7bvp/hrGpGCcaaFgcWyJjlVZPjYdCJSv93qhy3rNoFj2XS8Lyhzfxzlq
akD9zR3FkYJwfQvdmmmgxSGrskNb82sTMXw9DiCK2HC5yPy4a7axt6kFjS719ltX
c+66+JLgohNMKH/crOIRyRmUndrSKfbtjJE/L6akQphjcBquH9lJHbJ3ZB/4Yo56
W0hgUGpgPGoCbntEoRcjUFBuDuqP/SXfVhZCHzOraUuxc9mTgKacw2iNxl35AhWG
6YrzoYKZMYL4KPym+sU0heQ6WmdS3X253DzPOvvs9ewF/rcAZLifMNz1uidLW2cU
FGyUqFiO2JcS5RxcA8JL62OFl9NVFpvf+Eh6eWo7Cr/hQ4TsVtl4UwZ4MeQm5gQW
wp3WXYQtXog827442BwtnQ6/ifd3FH2g2OboxuYCPwI1PibcKtoPzaT2uDyOkgb5
rng4eXZ6q/e9OuBIJS+pbyBWauF3PlPT2phwKh6GEAyzOXmFjKivTkFdSJHJG0oF
N+TN0uyXaW82jyUeWM1wBCEQ52TmMwjY6FwqV2GACP7vA2QGRhkie+atLF8Xjp/p
K4xbDc8XbzPySjcGCRMmyugD+8SuPBYk0J/uJqrxCv6UOIye80ciYEXHjSR3mE/q
ND7BELL8LlTYJn/FY+Nd36z/L+Kt9Z80ERcy35kCbah9C75qvtG0CQVD0gnZFyPC
82e+tN3lsREDlfWQj+R7kA6QOVZ0szFhYFWPNBmKuocV8+K59EbDUOxXM4U/IR7Y
lmP0fDepLP/il+jxm13+LqcDJJMhc2ZiOvf7zVKS/yZ87Kd7NN5+vSWcSXBzK3jc
ZXKLFB/c1XspZ4S7xsxRGCcZZ1PjHTWymg1TsLwYhdWjlbZhUw2ydUAf6DDgj4wi
wdO9Po+DwUOedXh/hhtpYWmme/vHIXqDorc/qsyb97NjYPuDf/0oNoLK2wlaH8V9
1LAp4z1GKFrRUNozXlAtKa2md1YPfOdCbMwXF2PUXvKXEtBAOZdf3dima7jnuubF
AKZomnCsxMscNH5G6Z34HA+GGcIh2NQSAThpKMVxdgGHFbnlLSTeNen/jE5ZZgda
NfHJpqiNC8LWixVFROQrh9inxEonTwiGbqEZklEAAFjny6/2U7VxzoGktzjZ4f08
kp0Frd0FOmdH1gvHk+y3M/Y38Q4BNQbhwLtqp1coGcfc75mQdUBwzK3gPcmXJVYM
pZaD/DgP/bnqg0PbwLH9rcd22s446qO/NV19EM8OmroHl/7krsiqOhHljTpPT/yc
d+hRGWfx+UTLoRzPC069NfYFZG8RXcbNZSPuUbJXkP5fMbljFFZ+X/jhD4Wgjeih
kIZlaJcnYaExHLBxRSPgOGyZWMbS3vzEdAoJUOPS7PCcaLApR5VZKd/djjnpP/9u
3xM7PfoPyVRRb1K4m52YEMJ527NJYoAypQDEeM5/GDCUduQ+K1i8oCnaOCg+w8YE
jHl5k7uQI8qztXR/qdHkQyOcnEDfxrqPsuntTuWrdJDpMAiYNM4xuArK7A8hHKWq
ZuHWSHHxJc6xL64C5PpXOVYBdV7nsxNx+bNsVQsybeS0E5Y0+5vpS767yhejjWNn
UuuXGMdpAr5ukV0o3MlVDm/7ysbwY/sGVZ63wB8Jfi38yk83u3UYG04aR2ZydGrV
ckHYolOIRDOb6cowH4ojaMTER08bTnmuOWLNIamzHYvGzEa5Jb5nR/hNpPgeCK6Q
1NneU/Pt1D2ec+MT/A1C66YYGFrVe0iYWw1vaRJz4hd7fuLwOr3c04ThHbXCbM0t
y5eMSwKdIxSYIucaXnEUsmcAuHRcW0hw6M3yeg//eU1AKHObjvwbhFlEW+mMUyxh
5wvrSNJlximHNiL9igzJpOGScsBlnh4hBb4Lqos9Kdw0rCH+CS/Tc129MpksQbIs
ikOh+UK35L79ozZI4TZX/XtMeLkK1nL6koj/7PllCvy2UKB5H34JF2ev5fSvip3i
cnvultcF3BJ0m+nLQdLjgtv2B/zGi6+2LYSBaEXgV2yCKwWHw68c8U40hJCVdWax
BtEo44xCf/uX9X4hyhPkTSA5o3glc0BmJiHwkQUZuO7OJVcO/rjMwgqksMfjr3DL
SI7dlzhucLF3Qa20r7d7lr3UrAb0oSCvv829zQy1HwEaadCEq42J747ZZeswelO5
ZGCbP2j7fC+NDfL1/yO6+xoMJylZnRsZugEAvHki8hDf9fiLM4Jqj5t244SQgZ4J
pZ0DYxcbaHEu/XkheOXDr/IEn1kfPOcW+Dap45V1hHk8yjIycX8cG9yGbgvNrOFR
ciYL5mf87QAriluwWTnLeutORa2899kyX6J2DK9RJG78ou9k3ZmtkFjW2XIAcTgw
howaKb88HSXWgb50diIejMK/vxPBo1oxr0KSZZ7BCJiXUbMigJcuKsaG/k7u0kZP
9LQMibPc4UWnKgYHmWMTMFw03ZDuWEvipAdB+NE1o55gbiUsfnnAlZquWQ2fEwDh
5e4vlLrpybJJS0hwvly5pJ1uDzqS8isMUwCfojbZ722XIqSlTnD47dtp2BKm3KnK
mPB49IMneC6VLqFEPdt5y44PzOILA9G9aI0VoubNPJvgUql7UYGEDcrhjvpJr+0O
bmNngvux1mFKIyHV1yMjn3dVhFWii9ULtvXdW/NtvMgav6NSBhCdQslJGSj9bzDt
f3ViaAzHYyNDRwqeoPcagGD5fOR4HoGAw0kGS038y93noqqazV3Fy7Gm8SEtLg2o
8sQ911tMEqwRXYKyYpc9+PIdKNCGpkA9rykp+zNDVGZ/r1u+UBUtn1L76cK8QLKY
A86/AwlfweUcPGF8tQUOrMEKQq1ftTRW6H4c0E9VAwpkTE/0HWYBcD3oFpD2CS2u
zcxhyAxn8jNt7zbo4Cf+W7itbQg2CgCnrruo6BvJFMd8eQGTbWP2wj6VYcuS06bm
PT2SsFzO34NpwHEBI7V2p3/dnqPg2Xeze+ujwLjW1yZsShNfytZ2OGltVTGtwfM+
TDsU18UD53hbRuBLKKwseiIUz/zWIgJZgjrSoKVnlYMLVddGguNvU5I1uAOozo8a
SwXScLSbCxCeS/1PmwU9dOUH3bFeMyOEu02btLfQFMI=
`protect END_PROTECTED
