`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E1NxTmZXJmcy0y5iAaFuvw7ytofNKayAw7MRCJ/b86q12bBpIyfIvT1aYBozQKcu
+NIEArepG6uXdHEL2Ov5fLcI06hIuegXWz/u11JDCBZGuSSmeL4RdNs+q8AxkiTh
X4KaJZs2cPUxJEiAZ8NAIfED2mZiCvvvyN8kgDHFsbhSjhcb8vUPaUVj1JVMKsNB
h7hf29VSo6krbOxIqxKW+P5sbm+b9Dz2duCwQXA4zyh9FGxdPgkaZnG9kYshDQls
htf6YuJS0z4xbpiNoFpJV66WZp9AwOqUMpkEJ6GfruoIEZe+rBsBpaZAYLyjKSGu
A4VJDUHJyj72q0m2p75nrsQqOvXpDX7ZmbxFOZ4Q5rJxhsiWgBITCWXmXpe8nUd8
qzh+nmtQAhci+f0+rcxvPgMMQ2g1AvVvfCFAqpd7kEq7ajBXph4TvGDcJspdawkJ
jFGcAUpQKmnCaOSher+CgupZwOQ2nhysjecUv9IgDLsVv+l7p5LYoJh6JiUKi1ql
jrZyGH1YP5EHnm4KIKmXoTLPxksobUm8r/CbQZxtQAk/3u+JgeibOL6dmSsqf+wv
55YvAEI9cJECm83V/LSwFCngIE0UlP8+sh3oV5uEs66DtCOCgKMbsbV0kIg7RNFp
7A8Fr9vjBgPE46DSvtEIDVtpij4u+3xNM2Jag6WOezatkoKmyHYqJBeSr9D3Lhfo
NpBuTQrzz6rGz3KqKTqHQWGvtIJ0RNRFKzfdepUMGqvVGh6m7DD2PvTAn7l+MjDZ
TqhSqG3NyvbReK1NvPk/Y9E00VmlCTbw6VTOHE/DEap0OaaKXbs7PO6EmFwz6eco
XZmbGGoZEHDsMuhZgvfaC14V1cbeDqz1fYnUj+pjGEp/ME0Q4MN/LaXn82n4uJ/k
eI5syB+O/BrBEDVd6bWtmJ9SKmFbJT/N/iRfMR7jBEDhQEi964qKqABaZ+y5rvLe
Q+I4WEHhF99fndkaE1BAIV2N0UJwjQudEYIkAr/hS0mSjeZ/xJkh/YSVZVO85GCH
kwCkTclQW0UadERioBNdpg==
`protect END_PROTECTED
