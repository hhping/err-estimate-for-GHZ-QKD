`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kYQtPOQseK6+Qk8WLlecon4Y8n2LhiUfguhNSIpUfwfzMQpYoNY8dzBOY5jL2uCl
n8GALeDGi5ryxTZOA5DpVULO7awDj2fNObUeKSyjQLly3IOwuAoYMTnQ1hsnHbn8
KOIweLJvtSzIOm9mL+59UMHIqRe5qtAJmRjPENcD8op1qzQnBIemdxbkCMFIPseP
xkStwTVTgnDs1PsxGRVi2AYD7NE/eoXPdGfbhq2bfx7YJOrojvxluz1KkaHlvbr9
MQyt/ow+rKHcCi0a7GtO1QsVdFZEVpzVrsLf0m8CqNPYw3nk91psFZ2uG/PMJgT5
83UDR+7I4z+QQYNpQZW9ncgGYz+7mN1NH8sQE0l8Ctw6bm4xu3Q+pFlX2iQVtSRn
JTUvtqAaYK0lE/ypJnCBmDOip4qEOVsLF3I841aNBu+NxFLOhhdyDpicAk/LuAQA
sScb4+O3f6ZbFJGMcBerFtRwTOY3MTVKcnmACyIC/MWsPL8NE0kjo26avgrnsmEP
sgZ/F4tfcfD6owI7TMHNH7qzZtQarPURafwMlcV8yDkz/nFE+rsdNjPFAG9nzZUv
Yq1xk/bgPa+RD3BjKyXUeSmi+BQYqI4l5O7KPPbcFbXmpI+e3X8YnewwVquDYVfh
3grBzBjlQ/iG81xfrSrzaPSs6X0NTjDOxaVJIU5HqbUi7j3JHA6dkruZPD7q/oLW
1PwO1oQFvvbwWJP/y22FDi94DvD8PtyloiGySEoOAAQ4hYsXK5cKdLldniuv01Yk
SJMLlBvFroisYoEpQzQLxMVZFNgqZH5cFY/2bJ2wHk59kD3knOHLL1TS7731R3nS
yiGdXzf8m8zTB2o40IXp/eCXXQHxMMW1ZJ+zz4tb8z8NO4gcNVaSZo7imMPOTJTe
LGRywIdepKeiv7ArEMw0KtSUe2gUCzl0YzsvuOzexDddlv0gIkkCNrLmlgNw3Vd5
kSw1PmNPEnGgvsebpnPkZKux8yBDiddwLQA2GS40cJ2jXKvgypKZRX7drFh3035H
HE+aQplmoTW1ph8g1TT8M5aTkkoCS0dzFTtyeevvgQ8pq2FeoAc7zK3wGbDDEoH/
mGz5VA6WeiG/puCVwrjygI/a/HtoGybeEPDdClaXUL1vnuwGSn0RaLKmOXzSDcnW
lOiuOINDbnWZjVYLngR5Q5gW9ugTVpdQAvscx4ZlJQoPWGXbwtf+paVZInWlqJsx
d0yS0Z0KkyTklEz/BEpjcqIi+E9vDEVi+9EbyvTMEQNUv8sosJtC0MPwSIeIjwkh
1yElRvBArXpK53oLJ0Ktbw==
`protect END_PROTECTED
