`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tc8ywgGSusiRFBLvbjXlOV/bpZbg9gKUYNnAQK9a2lbMIVCm6aMUSp4mYP7qOrWo
TqoxNjuBPMW3SCj6SgqWaOLsHkHLTuxi7x/WqYUAMsahmbvhViv9jOudRGPQ6qyW
28atjRnKT5wO5qg8fvoFFfzLfZArBDBxM6EF5dyDdjY/120gUPJPg2Zum//r8l9Y
Pe/IEdgGMKISuXWvGhuqXdVOO1BOEul3W/n3qQsY/LZ2hP85AxkNsltVnrqLi3dj
Uduum2LL0ALgZCGvad+FM4fZa+fBPzemchyEGDtOneTN8FusJu4C5660CQ+Qnr7K
cjmJChAO/mjoo9YoBNn48uRWVphnoMXESzI+fO6yneAJHrSxhaWCm844+8DDauJm
qhQ2ARbfy7i8qwoXlnLfzA==
`protect END_PROTECTED
