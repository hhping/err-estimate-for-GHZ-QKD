`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sr7IbCyaDTkfzOrz3E5LXlvCYN2CLQKDDzGyNqBm0mqhQO8lsljyeIVVkUmliDN9
U0YEJDTgD0vBBmFAYf8MCMU1B1Km9w2Z9eSHXRMjvEPRuLbnxZmmhfbTJiYaNE/C
lsxPBmuaqcSDfTfMrcE8JbGfliCjrhS31PVuMcamZfkvIQ8pjkRTSfmNR7CbOJOe
iH7P9lkKPZJ91Uh/YL4K7YhdzvbDp6iZHljn0eRamYVsxyFpEbC/Cif24C5/MWI8
X7Kdgid1P9n02ZMyI08TBiRXMIwCeitTz2FN7bundesGc7mg+IfSyfbQ1lpcYJNI
v2KbAOMaDl9stVeD3ge15lHpGxg7lKbXGA58T0DRYl5+NaqetDykK3kB2Jy3glKH
HA6NR9k6Kq4TwTMH5GRRTcSIf9PIRMtJ6KOL57m4N0h12JO1HAy4+/KIcfY67ydd
X05r0JkpYUnFvv4dSRIDzWXGrxv2lrC9ReMgbDAiRe/ygqqOuQtRVPhxYqK3PfwE
0sFb3OnW4n1g9PDP0aVGbIiFdA55RtvLPIJxb51zbch6KvLg4etDroQDIu6ouyFS
h6s/35feXtVd6iGqSFEiDMbcTiIWD1kxmJQ7kMB7B6bDfKA7CNZyJgjYuXXTbgs+
ZmiKw+84v61XvrX1Kkpkg4zoreCqJRWXrVoTE5iD6OLwxDcbav2OqQSOkgKHAHt+
QxXZBtJumh2aCihT3QClL7v4VGj0Q4U+L7+AQJnEV3VHLykeoyGVqf8YwFS0Umni
2AM31tBynjbA0pUWmt6imhy7u0hNTt8/PsrSx6ZgosY=
`protect END_PROTECTED
