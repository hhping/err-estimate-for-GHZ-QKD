`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XV51IsvXdvhgJnz8k4pTnoH7AV+XhLf7pT5TuuEsIrYDnjRgy8MyMZVrBPv7lDvF
JOHDOr+V8J1+ad9/TMJd6upxWx98Fcu4+/KCPRald/XrUEC5e+GEVRpO2cyNMD3K
mRwE6+cO+GEC/frxZFWTYYLBj3CTYm+1imYvwecNlTAzvkkOeawzsWsIm8kRwXQ5
EuR0UGaabiofUfGoI/gKzuke1kGp3tq8mjx5Z0Pc2MDAKnRr5UAQqQnmO8VEIHox
/Uxw1g3NuXabx97NMQDKOeOqxaUJU35AGg0tt/wr5GN4cf/70LnDmkRR6/teZZLa
g9tAKNBXf+hGhAMwUDpiWInFc9PxuFOYjwAiucsejmmn/fFgLwXepXTHZx7QzQ6L
Niri9wm9x6WEkbxxwvhJeeQV5v5mqW7ibqXwq/06jTpi1LxskhVUJQQZkximdAS9
AsBXPFsjGsZUJ8ur97acsk0qYWmN+dqooHj2g20R9Tgwle7oOu49IaDRxKLyX9j/
lbdQJFU4nPFp7AewgbyO5VgJcVVN7br/fHvXLTrQYUV3OJnFvT6AWgjfoA8wm6Mu
48kujlWD3yGEh3s0tcs/DPg26OzekpD0JDAd8ZxlOBl81EvIktMLMw4zMYfNzjFx
tIQd467iYt905sd/gfv7kw8I4zmh4y/nu2lSLMYBuUgjpaBZZgMad/6STCdGPXU1
q29A3i5V/3ta/vH0LOhdhFVw0m0K5TpyCXBZB6fFUoqjhX/UH9iI8AS3xGkbQJai
sPYHI0zAxIN2zGe81U5g0U6VZE4VJYGWJ4AzGNLsEIU=
`protect END_PROTECTED
