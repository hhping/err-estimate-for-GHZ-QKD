`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kdOweecHADXiRcO7vydDGL6MQtASjYIPhNPQpVcMeQWWvin8d4adRSsIcITHFv18
QWWMlq443yzcmWLOCyE26ynKZ/GT3tNUhooWUsg2WFBJty4bPKiqT33AF4tIcYvr
4fKCqmc6OWjO34rNyrOzLfDqQZ3qLoNSRrQnZL4aIZBE70WwJuUGVDZlPXAyy6HG
W8aGSj945fxpDkOabKAA+/ChQdVge/inhtzjFe9oOroktxD4lioaGA8Kwk1aoKHe
Z/1PMBaKwkovYcLYXBTPLRxEuCEL/V+R5xx5VM8++WzbtmCOn2FyP3kkWIbmmboo
Qd7VwH2eW6rK2E8z/+hSjPRBSmHYUhdaUoKmSX8/3FvmbYOcOYoDmw/bxOJQyRaV
qePyECHIOT2vcjLnwU4Mhdjnxa4QAhTy+aoTu4CELiRtNc7si69Spqjt5t5COely
CQqUrmaNLvfd+wx9Nw9IzP6tzxSJMrmjxO9fh92pKxHPAmaULFOAoBJmIYGjiMw/
JsO+Gjj9Lw7rLL6nfbui2w==
`protect END_PROTECTED
