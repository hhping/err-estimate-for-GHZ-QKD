`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5MFhuQs1qk1LesyPyyj9l0XGdOP71auzM7xq/S0KohQsoPlhlG7kQbri8yUXYr9O
2qvTwlOxli8HAadA+KFjLmKCgXnOoXrPFL9m6jLjveU/Ez0xzhnjHZR7mU+5LoWX
M+GIIVcvV5WAgxk6YDlf/2OnnaFD+DWVNeljOJ+yeqNS6Een7/v1JmzFUc+rjd4y
XbPRaQsnarOFEi135dUXO5d61Rnh+TGfVL+gZCFV9VkJqJgeQAPQ/6c88m8W6bHp
rdG7J0CEW0yPMfzxNYKK+anLcyQfPj+C5hkPEG2tdhQXcnEwXikTe3GaS2ESRQdA
f1Yhq9458gSs+MtYZj2aJ2zXQ9jIa/gFmOckCjZnJt6coluz6upLGQehmvjDi5pg
NPH+sMx10bl6H5Y8k0QYw1UVhW0sjQ28DYk2UHNDGvRhtsoKkkefjVQpe3kcNoor
rqJ+o6ZNSo+EWH5yhid2w31XMTrVOVDm3A/QYVlMLebCp2wd2m3LJ8e3j84Zi1MP
7GYsPoYw/zioqXC5UAXIv05vIbRZSxZn7zGyFjjMw2XN6zMWg7sFP0E7uJcJDbwX
JKQluCe5ObC/U7H71iog8ioP9uIrOTOMFEHZZJtS61W9AfmVc3LWt4hFbc+YeP85
/544+vYHTvqQzp43FNj6Nw5mamiT7Xn0s/WrtjqICzljcIVoKKyb3OvSAbDuT9ud
1/Vc78RMtRFbhWkdzx5SkUbRDfIfDiYCvSo2FLaQPQSmwpaWtPqFcyj3L1g5j2WQ
rPV+76+/w/RXOiHA2i/HPT2eyaMnP53qCi1oVjj/LjOxHtOoKSZ+R0LwWWWh0h2V
msniQP8oSkxXX+hrv1wuLvr+NnEpPyn2VBQY2WwZLq2Pf41QusiEJLeogsD+04Fm
IHgRdEVwsxfpTIrgTneci7SbMb1bOGV9OhxBirf51SgNm4m5BkzcPkG0Ql5pUMIT
UvHZeL1OBpOkNkt8NCpw3h1YGpbDFnE6jyqAZe7LWHjnttSJD4aLs5wv7fFhw8K0
FORwOtkf0mcpKW89oSlYjk9fcOFxuTN/UbgysdOPiAZPoP599HltW6FBDoKqRFXF
KgARcfhUx3Ua8hX90ARrETvY8HyK3sc2/jUOjSzDTzOnF2o1+IWlzkSB6lgZrvsZ
Do0ojU7klXXQob/PqJKm3eihW6RShVyQYF5p7S/a6weZgyCRYNYBrYtqlY1y5EMW
VuMAlzXEQhLacdR0tcWJkSt32va2ooarV1GhAWx8uTjdLN0bmkckIow+/LAl4Sjx
Db89ZNqO/kBZl4rFIMK8g9LJYsgsvD/xhZgFHSmAzPrrgJ8VUKDkERNDP4tFYQf1
O1vHGyKWgPihPkXnohGy9B5MaoICjKR1W215AvHOUz5i9M3Dl+iDsjsC8bP+mmVf
1DxBI7Wr1k1YJin1x5eQJdtbpIRCYx2tweWa0sNL3hoS5Id/gdnwsfvuwQW5w4yA
f+iNVeXdZjxa91LlKV3h3JHKB661Y5tIyd5xiVbcT5UXzvroPM4vyBmR4jRZ26lj
R3MwVLuT1LHCnLQLLBe3cxXm0U8eFhLG6/YfXsOgPnNS2PlZosj0NfzAkx2jnXU0
XkNHDSeuPBmKgZP9cFATlrBW/UpYp/Vo6ewWIMwqu3LlAfhdhv/WnjY66Lq7ZFA6
vlRHjDTWyRFLWuY/dtQO/5rKoqIrnotF2cig4lBDG5RXp5cgWCNw/04acPi+SNX2
XbV81j6UOwAPSrMbKO7fce4Do9uLSs8fCJqt6CDuNfnsm73txrvxot19gzK5t9iu
cknhUNzWqwr7uwr6m33j+Un6/U7nwWpt993oDF7ZPrk4LVMho/jX8uiayaAyQBSC
9gWjsfqBr5E621yhE960Hd071dA9mcRRBtDRK4+Dn3+su2vuDS9Qidi2e5iuNwe2
BzfHMEvS7wXT7qqcQm6J/CYOxo7ds4kzJoYfjUKhMdeKsugGUXCHlomYeh0HQeh3
aSF4gaTXrPPTm/2/K0LVjcP0TGIPk9vmX1AldJGHhmcm80TgAkJVP/aey0rA8KUQ
gJcsLIIhLOpuYurr0mSP9m3xmwKPZdCB4LsoMh0/khyFZf1xCDXAuCSuBWFCSkI3
BoqGk7ScadCLzKD1OcWPufnh6UKYafMH6ngJEkW0t5Y6jJ7KadLeVE8f0P/AkoL8
yI4HR8gZo+oQCrSLi2pPhXiTZriRzmJ/JvTyIoRRXbtdElBhJWCuIPsBg+skf4fR
Tkw8b3xh+gnm3c60eF7W7YHPreKpp85tXNVI0KTOIEUv97pqDgPbgFJPaxjA3WTJ
FX6x4uwdmYRAhGtKB69P66jbwLJhuQDaolIsD/Z7A8KAx9MQB4zaHiMCtSBfP5wN
a3Y8/qcYkSVCBlCV43Ft3Kflat76tcwphj3KQN4vWqqkoQVuzUmiqXvcanAMoVpk
M2JfrT76rU8W1/NjZxglou+zIjAMfGZ7gc68gw6G8vvtzjmPrpS++XPUPMUJpejH
sd6/Cww4p02EuUSl1o6aucXfw6UHBNyClLqKt9Jd4J9VtVZWnXCpol1f/UgNB9NZ
Z/g7+xJD83l3Aq5Ie+/cTbVTQNhmhZXai3qVKtkdskJySShXBYYD4FlxVwmVI4kV
25L2XGmJijfSCpK7mpiZlyPF0xj6TG8sI5D9C8hQTEFAUiD6LM65OuMbuJow+OgF
gsndH3TF14jytEZ98CSNX9fgWGTKYqEuZrFYfpcxbYyiRdVeOsBf1wlFeH+4RtJp
+8FyveZA1jKx4TQ7pqw5D2zZ9iREksotgG9wcUAsBe7BDYoRUhzUVQTynEqFXJgP
jiMklw8dloCCJFyU2SMXAwXvJIdXAlx3XkAlrIQUlhENUk1O8x6mFlah0RhyX9Zi
1E4GQ7WkKJxj4Cmnptedq108aenm8vLEbBSrRVcOH/TUotewJXBUsetStHxG2TE0
b/JmCRZegE5u+7r2pbdiAuRrjyylXxvBL6Cy8EgKkSqcvjYZmWYDmiERxs6IGCsD
WqLbnAakoc8gE9Jf58X+k50ga5HAym+bQwpeDBFsOR6EhKAtnltCott4Z7+Oz5Aw
yDTzCW5ARwy8sWtDdGM4KkTqCEzgHMKUIjATJyO9cq62GwDh0hBktiEvqG/ybG5A
0zKR0ZU47ULgjb4bQUe1ERMjMCbW8/XexBlvpTDq/bMAmewtqI1sMgR/Xwppe0X7
mBFHhVLkOx9CIxY979yOSd/0j7FWoOxATmR4gn+MwkQaWHJywdujfZWs9/6RFbZT
l2jE9Vvrpz8gHH7dn+X6qfq5c9SPeSt8YpeFaERVkHkTSVmgPWGUqSotu3aRtuLz
8n1yRcUJujJzJdNShCKjRvzBR/l8/DSySVafVJTfjNDgofaOzxa4wrs84A6+d5u3
xkptWmClKh02zywBdwjjFSIr9NJBr6yVvZV6K1tpRGgl/W6n2V8fJVecZ9Nd/C4j
10mww5xta26P6aa5zLoJmzKtvbwStKVlhIAFBwi2okrpJ3HGDLsbUZcp63s0vx2c
Cj57fb4u8BIzF9rUzRhh72YcwuqP9TBUGO4OOcJg9X2xBPlpyLqlxNI8+Avc0vJ/
WQZx1q1Rq9gXb74Sd65gnx6ztOhf561DgINgLqULNrw2x8znjvpm3wt8EgGL9H7D
/syZ1xgtak4dP7EDDt0d2QpGv4Ju0jVtlTiC9kfE9BRb5Ps7hk8bnXFlfTiUv37w
MMno4X7ZHD8AMlB0IMA+NAIGs8CpIIdiiDl4sqDtf6H0MbsLY8klRq2RPyZR7wI9
Srqi8ysQEeX6Gjwo9k1KUMIZl9gJZT05Ugq6w9650zL1MmssCLTfbyPz26E5ZWAC
6GUh7+NaU5KGEAfIH4d3QgxSkkaL8rkIfe7GVVtFygX7FJUZ8fD3xSiotJ8Hkze3
aN3B5+CLbQTCDt+0HEIh41v9MeLfuRqHNFZ+dmpHAxwoylyzMUj5Mdb2DLJ7tRGq
KytfAPf5rdtYQaySoVwihZoaEtf7jv1V3HFSR1TAC9uFY1J48gyiexdKOxO3t3lk
4FKY6nbOJtUnrYbcS6eh8TrY2c1er/3UNBf+HVqiu9wIzT/cP3ZFaG3XyrUURVy+
0Ue1HFHFIi6sBFJDjUUkTsaOglUKKntdErlC8sImnvbadj38buECbtaDCncuxaRO
s4sfvAgo4SYU91twucXTXHiBRa4x+/vSep3EPhdNKHAzX4NnQRxckLw2s3xMVGqw
L27pNjhgy0tV3XfLkUtlyoZfqafarqXOLCMaUosqOsvp5Cehvkr3lTqhci1xgzza
1NwiPVG2nELvaDY79R/XZkvevO+3qcLFvCGMQhj1YKSlSWbYkaEymM8TaAhY9ePG
qSH+2O2G4VNNyKkl0+IRF7oEK91xwkVdJkF0qm7QmsRdVDFo5Z1Fx/qstnwxNgT+
GpC8mELJwiYTx4bZt1faf0HPFXDcXxnOrW5sUq/xY0uyDjynjohUblVGpsuIehLZ
weBZVt+lQxK2Tw9c/5JbDWNksjjtE6lheDrv/shOmuzTYyetGKGvW6OUsqg5NGML
H3c6TLsiYyRe8M4xJVEG00Tk2ICuOOzJFZGG8EWViVSaSRRGhFgmzD5Zi5fxMPq5
mOKxced+pZvAfJaQce7KhVzNrWA0WP+LtaXLu4onWIPWITGJiTLuz6f34n5CI5ZX
RGufhdzwO01+fHTkJMQZmZBgzFghc9o9L8D/49dqxv5KE4YwuqdlitFy+XBr1Nzl
d/OcgUWJ3NfnfRKrsCR/Z2wG4gH37RzR4dFBn9Y8PyryXv3Z1wYdcE4bnPD8ZkHf
kEgPgMEPflB7yBJXGbW96CpqareEsjbT2Mp5E65r+ryOlYWLkEaDRtu2Vu8Xg4tB
1OGUyMoMLskOJRked0CAbpFL//5tlm1sH+eXiMMUJ4Jj6BsS5PzIX9s3FlKIXhF1
VZD9k7HH7rH8e0V1gN7ZH5+mcn6Ps/Jqy3PlqQf6hpqnr17qXF6oSchUTILizZ6N
g8Lx4wH7hGnS175StSbAChcVS+soPbB0G5rgEemcSbSdGsDszZeGyQkCxGXNzwrR
pgxs552PP+E05FnehWzYmH7wRBmmdMTo3w3DoLVWnnXtYxRDKpG8CRaEFAyUR4l1
Cu/HlgKrXdFOGhL7VznMMXnmXRAabWxcAmwnm7RcNbRgUaH/cW8VZM7rY4q27ta+
NlRnLJjejH2U44Dn4fHR59HwRDq+g1VHJxBDJWI5lmWfRnmbbYSkStGAKXTQte4u
dhnedS1wAac1WpS9IZCuQELOAc/bq/8ONVF18uvQo322Y4rfa/q60hzEzNXhs8H0
ePmb+zV8lx1rD4WGvy++2EdUTqLXCy8Y/YpSWDyg3LcYSE+hCDpetboJE2SfohVT
rOdkQ6tH26Ytbt7zD0NKtgJ7pcw0bIyWS0zzeC1ZcXgUMsP6PQaQp+ygkZPrvN1C
SFbs6BG2TmlovauiKYN4vf0hDDrW7qTwAMoq4dLCJZSBAfNQigiqikcXYgeU7InA
QRH0gaoAJuTqt7NMxvvTCYwHYoKojQ7NrYWCpbC2uDhw5a1LtgrDgfHSblOY6PjO
KrPkbQ5b2+DI8gWO3c9YWQIw5A1ukjWqXYURTQuWPVQsJry095qDs36iYgkjISsM
gnpJwZHv2SSxEeXtdW4QrikFgREdKO+O2EJKLS9SAYzZbg1Br2bvfxZgrasxTwT3
g2fkJLPmlGncogxoOoIDncXTseoZLaISlgS9ycmj0qjtScmQNeAy0iENMVGOrRli
DeCH/VBJe3O5K6I+yTxPTgHG2OSwEIvnWmZi6mJWMdS6lu+HkrHSPZ2nUyAm9V/y
EFlp4DwEQnUE6E7MWRIK+NgRajybzZ/BFFYqlD0WuHfOpjFX3VqtL/obK5J+90G8
lwpI9O7wHP7k+litN8vyCLyXBfmJDioE+0+S2NvmMDpqqLoaGI+QGg+K7i2E50Hn
leijtYMT80rIq387Qj6UXvms3muXRHh81a2AxIwbSLyI19+p7HdkImc/D0FTVidL
TzDoZPdFNKksfMw9OfdZL3+cF04nT8NXcwXhTheEiTHfaXgUdV0/u2rv0cwxa8GL
rEgvkvFLYe3uGfyLzcyrNu4gX6JjTSIYU4Gq2ZVix7n8zaeR0vWnur6fSQR1o6BU
tiQt49P/RyRlFtUkWGOb+Lin22l6HbRZpQPSAKznCsQbYQ77DSX7m/AE9rEb3utM
`protect END_PROTECTED
