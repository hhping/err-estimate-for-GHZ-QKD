`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8uYR7BQGZAU/ws1vKuzWL+Uus2508yy4igwQRui1WEZ/+shSfPGz++6TEyyssj/A
dZJ9w3rufwoM5wr4XWULbuL2qEC5XmfTt04QGAuiwUKKZMnCpQ4fgi5jOxfH5ItN
2nKikIE//ve88yPSf5WO59OXAoOTyXNpesEEVB+B+82qv5LZeUGh7CscqKVIPnSE
uHn5IQS0RysRfz1FZ8jgtVVP3XEepC1RAtOywQ0kp9Yd4nyg8U4JzgkHzSXnR1EI
UzXqeIIkvTVxChGPvvhMv0d5iH3LzQgbkr5Akr/IVh5PglWqxX5G+2Mhrc8PYBBD
yxdkfIotPQ5spHsURLNc7Ebw+oWd1ufcHzWCWlllUqmcpB+2T+CmLYDpC414ktnd
efGI2IG3GkU3Fr8MIXhTamJNPcHzkni4kPyxCAAhrQcvJtJLFlUj4oFHf2HL8JgA
pJrbHKZE2djjHnl4XcT2oEYq9hUpJoaP9sLMTjUO7qRsxzCbWk/hh0hR1vDK8x14
ICB/U817wTV/Xyv9qM+SSQJU+HrS6FhKI7/YK1DAKaw5VDzmcknHBc7lCgEKCy12
+9Xbo5/YpD3uH3zKpPQxkkjBIMI4yQ/q+16hlpj2QaIWH+0OVrK5orp3/9TSg8uy
Dxje2uMLPKt/d+aTrxPRMl/ELWUNJA5nXA3hjtdtX3aQjmls+jWyn7omHjoBFlIj
fnNi8hAyA2mxV2TE1BIpsC1GXafmBLIQJTvgSZdgccSzFEg+A5KeHr+OlTEaUfBd
yV00zQHHR44q+sBtfCnqfLzuVA1Av+EOWn8cBFhFroclV6GVmGWIIkoiwUI7mbvW
OEpysjk58XaAQbrQntLlCeI/oU1oWPw6MBoxZpBQ/HX2nkmIt1DvJii90kZ0gf6l
9jBcuCoonzqcgqK554l8bFf+50aoAlamMPhJvWlve6yrP4IgMuexo0wAH89JDIUU
bL+d7JIu+/Zn+DymsPtpzAHdMYwi074vgDbRznUBv1cyjewM8DLvH2PLmyPyrNxI
Zsx6FCOK7OlXfnmtdE1PXStKnTk4S6dZXmsyLdW9PnaQsMZiJfI2O9h9ucBQhnVX
cL4rCXswoPAq0BLlugSyZHkxnOLLg0PlybPuuDW8RRgGDnvU1VLz2nzKa+GgXTcb
+lkBXaeK0ai4n/jRpwO+ewj7CMptP05VXhJHzTfF5amBVsfBUbuz58EPlLRlQWAi
vNmWXZqY7LHPqgKheSD2VyiOhZfU+jVnc3bMxmJL2y13UMgljm2JDAGOnFN/cZEN
maMnJsxH5zuA8rlfemOxNQ5Sas5mzKHs9TrD1D/Ekzdu5KByfbz9+bxTvHhtuJTG
p4FQKlMFDg/vHOuSFxDj6UpgW/qYFPs4XA4ic/3xepyCfG5oVhRGaey/zYah1o37
2MJmaSc2tEAhxDqyLZFTjgsApZssSrKH47F57SnLyOPhI0Nq+i53K1TKWJAV0avY
41UN7zTnqgZXsKFwF5v+B7BjaSJHiAD/Pu1nOqNkPd1Kw/FfDM8I7QR0aF803dSk
bDGRqTYfGZMwnFyflAlkV2OPMXC5SHq7Y3yU1cVRlV+0JwBFMdKKE7ilmbhxlzEJ
B5BZmqTTKs3zA99IjMMIE50UiTg+iwjWry8hPGySEmxIWxsUMj/TCq+2bydMNo1U
y6sq7ghxqiQbsldlGNE+73uL7NhRvqeK7rRNvaM5GrssuF6h8Rqc3OSeqj1w92MT
pdEw5TlcdPGyYhWk7jkT4gcM6c5T9ATNzs4FA7Mt7HeQWAn5IQ8WjLXt3TZjQNBG
F5cZ61HzQjNdE4Dr8hq72Mlr0QRE+ZvQChbZsOrCz4Pxd068F5uIU3z9sh1LaMVl
l/R3T3Q4Wk3hhGVTl0phpWeik0PpyfWQe5wlgfaoMXiiyNBcpzjOheTzkqfPi8s/
ui0uta2ELri7CkNNBtww5P6HzDSullQkalZC2fy0lNgnufyxGkYYgUldPWVaM8BD
Ob8wgflKW6p7xy7LEPNrMYl9Bhn60micfVF1/AhkpzqbhqwpwzzKopCgBybQN/XS
3vlDQDr1Xwl/+q0GODguwtXGY70gSjDgsE2i7MAjpFGBP2zy8pq8JDf+1hLnYgQT
Enlb7/ou/cRb6zqKNfOeBB8jFcAbhIWzShNiYsi9v3hhNZtBXNBMKfbPw4nhN6cR
+sfdWY9UkwfuR9MtTTyG+5Jpmr3ytlY4DM1XHCIfan5AZ6C0Xrq6Fua8i6W6bwrO
s4V3Vr406VgtBXnd8XAPopusd0jQRGZv+oQ0JCAq4yrsFOPRAbkdM8GuM+NmfX8r
kpbAo4zvYin7wKM6IrVzn0EQ2pNYxMyvAvQB4DatTy8B4AB3J0//4N/6YptOyGZo
jfbawM4moDBDh/6ygGyEikKmIA9kbvGNIONh1Hm4iaeaXFP6sDSHLumqbBi0ELF6
VGV6GC0IjpbYh0DKdH2I9RvMk9943oUuFm3uTAWh4cM=
`protect END_PROTECTED
