`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KQOm3m1Y1wL/BSog2/2q7yY2FbtwENzhlFNlOEhw685YqjMzZXFS1+uSl90GJfe9
sSYKjgTtSMnPNCaN4rtSvnwColROD52UUrWjK2FngtEtlbJ37MsbHVEHg6fwcLoJ
CxSV7oXdoxVI7Ca/pX56eJpZjBcn4N+BgLODUuvvhB6QBQIY9BG3zqE1n4QgZBLa
jw85CLBWia0mirCRetAnFusD/mLiospQ6vSWXLJ/25TuH+8DypEFn0NNYEccPivY
JOePoN0FGiaAnT1JTIGXf2oAySR45XmrWCbmItYdGz2Cs7dRIzseILomRgVqkgPk
hM3pJmNBTAoJp3mLS33b97SCdIQXmd/fIhWTZ9aLtUDcTUnNm+rhorG3DSP7DTeW
Rcsukis0ohlOMsUu99xTnC79EOIDwKsoqMTi71qDD965Dbk1cfP24TDKLA1u57s/
VO7Ge1UbPTV5NuYbEHAolLi/Mf+i/HayLxOmQ8RQw3bW8ipPjQxmfFfSwv5fF6q8
UMXLQgIA4sdlDNqT9c79z9wdnnA4XJ0YWdv7edgaTP709uBZjYP4RbZ/w2nhWzjS
rS1lk0RsM1eSl4jAzf/rXWzYCXHS6IXk6NNd/gvT+FpFd8k7iY84vgsJCy01wH0u
rLBTJjx8LxrPSFg/RTATE8eG3mNMU35p5tBKAnJi9EzOqQD+hMZHSCk1NSWeYyYe
DpVPhYUt4axgY6HjfVrqY2h33via9j9xicCqClY3jW1yn7RPRoCeWpQgYfvyu57V
xmrUQMA4azNJbtnWMT31/2SHCeGLTUP3lXQjHI9ehtw7ozzSEs444+Tc3Ro+WVdM
QNjFNG5Zt2a9SnVXqFJZJmn3RnKgOSLA0Zpg+K7OkvstTQMWPZ2B9IRuaHN+8hP0
hUt+SmTc/AR/Iws4UgWs9nDidIaufmxGbOfk2q79HacLLrePsX+XQ/2TRyqPo4Sp
OCFFuXwoLEoIEQJ+pOABuLI3PUZhFO0Nta2jiJLKydIhVElkjU/Cb0jIhNExJxDV
Kbf/LQzpEoZ1R2BtA0nwyIZORl0WV3bI0nFHasZBcMJ6/qSwX9Rnjr9UE5GNuVWj
v46QrtFJO1h/ldUd7Dhnri2pF8FkzM0qIFmPemkfjJ8KgpCQb0NJQ70ZJNvxAN1Y
f/zedpLWZ96FhR6GUgIBw9tEy46hGjfzzyqqXCSc9vjCfdVw54xnLv8L+X7ASHpp
VCvzlG6jOlIeKdbvf9Jb8PC37k0OJ9pM8WLRNlic2UgdVeEymxSn5OQ7QbIPEU1E
oHpSVTkRRE0u2ZGMgcqARg==
`protect END_PROTECTED
