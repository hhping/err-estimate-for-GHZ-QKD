`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WVhNkiKs8J+pRLkNEOAy/FU2mt2RwYpBuIszk0VA2cL0vjo9nEZJ8AJZcfkWFBkH
ZiDk3sOijiljLaSyiGMz778mBkZMo+CIOpFWhxhzUU0zsqpHrd1BkVpPVaFYCg0I
e8Cj1LBKVSzedP3xzH+J7pxICFTdPDlT8dIIPo+EVxGY2BgsQpkZoJF7LVj+9BM6
D+1yu6OnChqVoRjkGnDtKOcgzHx+xjiKGk2NCM5c/oi8fq6oBJyus0IW3BHN8Uju
tdj9Ybrw9HiGnbllGfO1zECD/ZV3Ea8TsCsxpGwPv9xqAU9tBsVeMu9FAHRtn02a
xskYYP1Ep21RwHe5VvZxEZyctQQkKjDRPuKvyOuSHG3wF6nE1hRZMMtVUvV9S7Fn
fRQ1cjCDDZUR34ec9/0sT5zEecBowMdydrAOyxtOvRR7jqoRDX2DoA5nmaSnHkA+
`protect END_PROTECTED
