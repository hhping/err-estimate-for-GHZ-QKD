`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YpnhRpMOQPEBRBuWNthcvogkVLq+gsfYayS4wD3+pJTShOnaYuaQ20tIdGK1+Azg
6OTUUpAc7dwHFJVRkgmT78D/h89QKK47y9EIAMjE9pFML12eNADw+ypvq/dgbDdc
mjBuFKPHmhWvMIw11w30pPhiWRbRQdBIxuODUd8Ls+gDEbvqU086gBd0LTn4Fagc
NamaugwsFReYbVVzRQL41XeKyzEW+S6KUC1bOQU/gHAPfy0AkrB+aT17QR1CDASx
NrlCGeok0OPO6u26Wqgimcv69Rf/EvEfWSZhibCkyeNx8ia+oBaNTm0BbwJfMo/J
wFYq6Oao0iQDuiVflDPCzlK75EvknGoKyftI5N4QkGfrftd65JY9OkTRg7H2jpyJ
KA1kFq4NHarTO4316GjGhGH/2Z16Bbip87WDbw6Nekz41o2JPyGn2v5xphjug/AZ
XHenI0q+RtGBjYQQoe0BjK3fE4DADjm8iwR37qzAcQVDlT/B+pkJSDnwwFUSu0IL
fxhry9/KrW/7GvhmbNbERobbdHgBzJ7ROrK5BQOWKgvbo0KYU5uVjc4qUiPdoOSV
HB+rYQzvuNuMcjEIa7oWjBvKQKUKJtEHJGwBuapgGQ4oAGUUR9trEwsEUysRUys7
fnll2VARCl9FuiAW/Y13GNERIhSzr0c00V7eDZ91DGI=
`protect END_PROTECTED
