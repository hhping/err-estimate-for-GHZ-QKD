`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IFzWSsqG13qlWW+sHED8k7p/oKJpe9UZi1nf28dmxiVjuXl1xeS5DfKbiz4/gx0l
tSFwY5d0TDxVQGQWluAg0RYDqbgYDrt9RPZ9NMWV1uzgXA/LKa/zUujN8UUszV6R
GcueWmHAC1VcZ9SvkScPlBtDMrTUSODMxtEUKQqAq6aLtGAL5I3TSyDucUMHQYJy
Gplo5EWU+phNSmg5EOAaEDnIR6VDktnq3SYLWKp/8wr4qQlg6jTTpW9n8JQlWIGS
7K+kAnId7IvKBpqTd3a8OXb+m9G3iJXq2xtw8F7I5u98lYEqm1UubGiNKckJDyOb
62VlD9AbMBoivHds46pa90einjOktckKhESxIZFvTXxjsKYdP2ANq4jqNcsgxqPN
jWR+S4/2Lo7+oiR1Wcsn+WWzy+IBTrcYKBy7ps1q+NlxYd9TJr+ps0IyW6zyi+Xb
XGGLbgDk0k22eFJrIaLBLUgTXAmO6hWmY1ADsoCujdTHZQfMPhXC6ZHzuPPjpQzK
/Y+Bp/XOn53xVSIUkf9HlHNVYfBFksJ5Loew9k5wRXnsIpR5vpu3LV38s9TtgwBF
hjd3u9GDHb1jlyOTxLxBMQYMIlM+8eCBqQzgrZ7Kd9pfH+Qlvbg7H/MNYrCP1ZUs
pAk92BaBLzWIw6PFvTtUIbGDimE75VMzuu1vGzRwxU5imIvbRgtwg4Y8hb1S10T+
Utz1tGYSGHetsccbK3G/mXOTTl7e36xAJeOq+dnF9CMuQ9WEqBQNr3qizfiUc43+
IJVGQ6GbEbLeCN+gJjhu1WmIuY5LabYhkY2wS1peSF/eKXO77ixIjs7tkdbzO+xU
i/xsS7CxMvLqnG+z8ijE0Dm8hy8oZuHWAdev4XXea/GO+YLjbX05LFM6kow4Qr3y
HN/F6rcq4oxGcYz/V0I4HJeQz3zkjNrojnsLvHVKe2aIg51klTI1VBWcWIy6VLLJ
7MPt6aV7nJCuxqZgdN57DT9Rj09ZRfwHevp3eEWR7Bf8+EFsJ7/i3ybq5IOCkfQ7
`protect END_PROTECTED
