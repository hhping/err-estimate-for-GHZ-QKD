`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nK5yzkF6mJmAEn/UUNrP+TNShOF2WolecnBcSqQgolVj+xUlvGFMGgV9JWwTQC6O
fGHoYi0klbZwiTlFc0nx0UUNavmhGczrqXl5RaHRZ0T9V1vrZ358gEY7nQGTddsf
pevTJ+GVnNZFit14ALFfu92EYb18aU2q79d5sIOnsRsQQ5ezdSITQ9cDe5/1vUWl
l+UVR9S2Xm1A2g7VuZoGkekZNJXQAexjT6q079jUoi1f2d8RSh7VQZDPKmNU+jnz
4m0Uxq3ol8racKx3RJhuwCtRUxC0AM1AsdKf/7PtHcF57Dc6XbuJOA38aQzSYLd5
T6UiyeKe66FMdc4UKpCGbmMkVHbjA3eGUSsvZSGXaHNbYBbDVuVZFHBwGYQwxU7v
AQb7mFoxt2+jFo7zIX7nOQwQ2n0Vw7bOcTTs0L7wwQF/bZN0aOQpzZr6+Dm6Bu/h
OO1D3xG+WqBnjwQiMZu6jHhSPOTu0e6800erg78xEFBiC/aOaAIkF5ngsl0KkZ8D
5xCVSDHdu4dhRGvIV6AmNExDv0wfsKojZkQLPFSUfaTrdJ02ZQjgNErFvguCs768
OxnZgNnb2I1sx2WytuZYcIO+L1E8BGz6KwQDzEfMKU5uvHxqCjEoMgMMJZsJoQzd
Uu7oSmRmFXY+LY36iIIQNquWom+9OxCpyDs5RzhU0XOrDfehocwe6YFrYh9Ly/WQ
t3c/H/5sWQ7BJo04jehgNxwUg0Z0XFZjMIZ2b3oTun+jS3Ub15EnJ0aVMImbqIBO
DA16iqd2b7y2qgiIopWfRkQiW64uVP0sSVH8xy73MCI8pmt++s4juhvyq0bzAgWx
Sik9w2ImS9ejGTCASwSHaaQnCENnPnDenPJb61XPnupmPXuwtdvyZUJ38R7+hEtL
a2fTUkcwIB6/FrzVlWwMAkNB5+qE6zQwlB2XRk5ugwDf4jtqBVDbjMj/VhlH3MHa
Y5oR//ie9IrbL58reQqyfHdCod9AgtxYaZtclovaD2ZhTYoqIsC6/Yxb8OVMrPrk
P7FYZ81jC9QTkCSebaUYRoVlRrjSsyVPaR49/59o8nvvmILdh4Lpji3dIscLfEKA
yhYf+0sliMS6gqzZToxfA+dAHILQLJhDULeFK1zJRje+0FebgvS5nb/1qBSfQf5f
oLJ0OQvHrXO6xzC44HNh3S6rfZmPyyJn/E7EWyFasfuUAx5WJNEw8Fv0sk1JWHRZ
eQigpQaCNU4puAUH3nCRW6zhSF78szOVOOOwXZwtqBK+4NctJTCJvFZ0KmzyVaZJ
W/3yCqUIH5oKKJuK/73+IdlW7kRf3CDeEz5yuFMhPtknXssHx0TX0DileEAUzDz9
defsrVMybpocAMy/1aUuXxv4kyzWcUOpwfy0x6mwGCKh04s1FV9zHgZR1wyDUeFv
c8k8wPGDzrO5zS+gAlv829y7swmxvJQDGgKchJnSaM12m3nm56btGS0nhoV35tfR
UakQgh+Va+CBOxNGN9nbEeQcCixRwBuyyC4C2KWPCVENtqJch1pYJd1AvhI7e+6a
fraNNanv29PFgUSLBz1cIVka2KEzKb3JnwoMxiwI5cAUDLOiICa942NlnPO+U0UH
ZBNwwaWJ7uW9KwMjoc0DN+vy2nsjGz703z2OkqcEDZxNHRddHeLg9hQi+Yinq7qI
YZklY4gCkHAQss6Fja2+RdxUF300HkOM6igE/N779k76SNXrdzRnNf36VaIEVJ85
GcuwxOcY+KQ3vhQxPFBcsQjAe+rMLmwBGbbzMF2ErxG2BnwZO6yZOoR7k4uwdT4H
5t3IZXX0aGq7dDVV/CScCWXL+S1QpsMKpXkU+BTXhg+3pimQrRaPYfCZTWO8e81I
hgSMw0sqUGkWWf8Ah75/+NNpg3KwnQ7mbdVlbW5QGq8NPEmRawwtGDfa2Wu/a6E3
CTO2CLcF1s1ikzQaBb8RJeV6/qqNic378HRpkw4dXKeQo0WnNd1yhot5CoMQhc6O
F7f0uADxWDObnVGjy2Tks+TSE4YlPwRwfENxAbgs0WGlnXMP8oLcIeWVuENIyAAS
ke+DqEwRU6s8iL61umwqIjI2gAlUlV4CyQR5rZm+VcIoCEOx/x2T1sYupota6s3S
Nk0E86tb3uz3jriX+WznDar3/hhiv0+qlJqgiNLfYTCpx8Mx2h8col/oPk3rOmv8
NfuIjdCUQ+e/QVIQpaY18STrA5By4YlLuP01S+fG2cJzdN6ycparG9dtYZea++AH
JTEgcn6I1ix1E69VVdPAq02wUsRJShbMPFS/5yaAr3MbzlyGAWdMpOVv/Jp7dA/X
qTJNqylBVawdc2ZL8HmvF8gkEmSARaoqxU8MZ/t8RIvFTuhiPiUVY/Pyr1yt54QZ
hUcwybQU0wMuRqmRZluOuTlsrV6c2DC+5MMCPEb4a/KjsyzGNdUzxyz/j1J8nRTb
650l4MPG8VIhvXssVA10W2DHDiIoHxWhiD1+ZEkEtTB25Fabi61P+p/kKS9dqTPy
L1QjqldSF59pSE+DvxATEVPDtHg+OldnEpyp0WHo1Xv6yHhGpzf52P6MoweGMJ3f
iWmeNl/ki66flPg9zAsGQX9eLdGoOfG20P7M56r8IykgJnD1Jgp7AozD+W/pjeV9
pyNRkZfI3AW0GILJZQ18dCcJu22aYq8en2usWGeOnVkB09YtCHY8ZwTe5F9ATLJ7
+VEXwx/OELssy3rxkhBWx6q4FiPT4AQ3PYsZ5tXoirqhcQD4yOjJuzMZRwfXkDxG
bMwulcTFK1zDUjcuXMBax7gNXKaNbF1/90NUqC4lQ3GPUBFvKpSWYMrr9jXRLGxT
gh5B85/8G0NKWgc66soEL0jcFFYok/tH2Pfovi7VGoeYpf1dN7WCumOG9mHAARuI
Calw0YN46axi1WDaHXES8gSDA/5Wu6AxxegFNchNk1M6TG3r8GfWUaEHquyz1gO1
eFVyzIkMM1ZuTo3EiAwxfPdBKtqGQo5mmlYFkHQmhs5u/FSYWPoimT2jzJ+ry3e1
XJlZz3VQpqMRV761k2E08ut973CHIkHAFMIkdq1IL+fk1ogidWm2GUc8bdISsUfq
+RRwUeFQQKATXQxUdL45zXU4O1EOigM1wIKBTOcbZPtnJ0jGoXruD2WxutWRVnYP
6I63JiuWgX1XzMS0yDbgnDmXEuQungaLXYqgBtAFYmcKJkou+R2DAC5k2+9kQMgu
uDeO10mhTlA8IEuafazgPoQY5Bzx9Vl55Nq64GbwcGe6PJs6Xj8I6dUOKGWdydru
wccR200nmGmvzOPWrxjLVHN2tQkTtAuSyMgtwyYEC7rZMPkACZMFP6buVgZM//Gb
f2LqxvRf5+AWpRYNTvo2gK6algBY/vCNx+p9FHMve59VQEmGDWmG487Q26tFFG3y
RcIS91U4WeTVsTDsSDHnSqtHyTwVPPK4Jx0jqwfvxq2aozNMj/1UuJYZ3x9Wqb9n
qofIvHAKbZG/RpGySLagna/pCXgqIxbU7kix44H4QS6F0GaPzjwqB+hkDMzZmfYe
17XxSMhVTG5eSe2hcw/8wtTir3cuhrQYwf6DdnSa640W2ub38SPNqMQpVzjpCZJd
NDOxU7cDdYbuCFsQF2KBvpY49jj8aDYrMHn9/STQYJOm67++V9TdTg8sAxEQlOKz
gq0xSi6p1RElHsAIjH0RMumivrzX8kcGq6La8Hj2LFViR8QwkoMvoIDuuKAn3kRE
kFuRR15rhp5UIi3dPniOwrdWvigJEn+Jql40QXyuQkc3ikQIWK8/hIRotmEQ5e4E
31050UjcKxwGwOvjYngBDDq5tiGVQojTi3hJ7ul3r/TGe71YK75Rc8LSdBFR0aII
45pkrHhyHCg2sZhZOSgm98xV/ekUBsQXA2QJZxSyxkIBHcRItUJgk+ueenuoPbbX
6T6TA2QuKnIv5Q3ez0c2SOs5hUB6ZQiIoUCK0ZTyXbf5uimgjr9+h/HDqt8NAg85
R26K6T1G7C7jTjz98CkKw7Ys/TQEIxslAEJ8ICPSk+18p8/l61hzCwkuDh7aCRdU
j6BPtcWD3ArnDISWocqc7rN3tOp9F8Wnt6C2mPy8tJd1mngYr4VLDBLhx7zSPnYb
DLpuJP+FvW9QWkWeYasqFFPlj1N9+OjujzWPvgySW+0NKO3o0Ae9Nn8ZwgHsqYUf
jNSc7X4BqFmca1Lg9gZZJo1DHYv7eNv92k/sJWyt2UWykVg3KCZgQ5/LM9yGy/j0
sE6vo8Ncnry/2MQdyK7LKZlIdBMauZr9Uu9SIvTtNSXXgrT+gPRsi1AY7V1vOQLw
hkHevpK5ilq6tioZuzsY2mHKL79HQamqbMSLuZHav7VTY05ZQKlrzyqHDcPZzLn0
vEghSiEekWzvYrR3FFSOc8YYAoX8/Fhyi4JeeG0MkLlq3mZmcbR6QJ26kXBfBk6B
5gl2GgiHmkOH0vM3M0QZ86OCcHvTzay3Izm4+kYhB/gfwIqd4lXRmyoPvrQWA1LC
LYuMnF7TNOx9uWGdb4BxEuFSJqLEfkXMwyWViGEj23Qaa7wwiunhgYNHderCbzjV
WwG2SRme/HkiFiNiph6/dQ8MlOYvszDJRdDTUkG6MGK40+m0uL/dCMR5oAk8Shyi
iBKstXGPFVMwlVVnJGM5L0ROj4BjdlNmbvxK8A6jIT9wCgjIym/qcqCX0qYvFmH9
ihu+qCuW+qot2ddiQGd7wW5GZS6B82Q5pF+IwCTh48+2ACMxMbg3q5L/p9wnpDm+
ozqY/rfswprnfSAC6X8y/dZ75mahiP7fXOUhxgtISBmfRKdu5ftdxelfR2UgOAMl
GINrIpOIkAFEDJ1nowV21WLpJm/OIc+FC6jRyHLCRrZfUBJqytndR7fSFhSD+vzS
2fF8YfUA/dCzpqU1Vsn3fF26nlJU7f+5UxHSjRzQZ8qZEVW4STN7+ImvFaAyCuEF
5We21/ccOXJrInWZF4RViGKbxWnLDXfs2BZExETDBwC2+sI9ZQcs1YVS6aAB+7bM
0D+9VQlDp+Emq7rtrg+ROk0NxKdrhdzdYrfz3mz+c1o0YmQ1hc98j/XeWVwG2jcI
vHINIuJ6MYyGQglS4Of281P5DjdGXliiewwKoR35gRZP6ycHfM8hr/87e17fs3WX
S7s3tneIB5et4ATcfH2WBc9Akt1lwCMWFg88F1Ig4Gjh+1KuEIqNCm5fBqQgW0sX
uZQRxHJb+Th5xJrzc9Ie28w4NgUuHycjS1eI8JXy+vVynI+3515lWMpBh6kw3bAR
icR+2lZkHGmPaz89gaHoo51KwlYcMeV4MR/owJI27YidZOIOcKhvjlUXI0/L4aM/
olIieLWxDJYCoz82i/mTJsIHUqttrC8sJV077QH1Ual1c9B3PwC9o9gLdF+mHiyp
iYBvayRCfr/MnFSmXIPTRu9uUIgnP6b6oH2A+gmNzTVwRBITwh73yY1siHxOZcQu
aaWcnWPdu/a3/pstZO/+T9raJvw7nr35nbWhSG7HoKUW8AJxra5j+AWvAS778b+j
deEXu/0+fy06H9n4WqCTtlIAOGjMrM9IFPSzUEx9JSkDQxkGlrrfXNgT8Gdydb78
KMc/oR0qpytsoR/m5UVLg3gya6gT+QwUzLwjlxXSq7bWoS8cx+KvMcQkwuQHL5jP
hOsvEJ04m0NNAZ4gxDq6MFmbWSYheDb1CW+RvfUJ8PcVtpX9PbCAhxIbVs9EH3Aa
eHPldoZrkZIVb+GI9Cw4oRp0ss2Lo6TjMfc3lH07YLeczTYgSzcdgMkw/uAHnt5y
2UFbzuJidpktWYgDr0ZsCxO+bBCxA/KiQ4HhhcQ6nj3b3iESFIqXBCPx8WwzYWny
YVGKbk4mJ8fu43N6PaFjTDajjoUplHP7nr3aQgmcH7agrQkXFtwRRlvRhJnMxSA8
Xj7Ed2jDAYbZuGBLR2BeyGRuEMvoSfa/b2EiIER5o30=
`protect END_PROTECTED
