`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8YOvwCYk5ETbYRxSP29mL9hhJnlVLmp3fKps6QcnB6DMVT5mYi8bP82AaauJAhgW
PlC2G+x0ZPL5j2vMPlkdz+pZZUl2baV+4nkV6SlRIxDUcJqPKYvSygf+zL+f9AS+
85HO3gB6kmN5qzauVbrdvPy2Fy0Awd2mjizFtO36rwA02ajazwenv/r2zUZpP6AT
V/G18SVBSlE/sV36vhwB8+boky6wXiJ2bAUXJNJeclEOG8g4TADV4LFdtqExgHp/
rLuNW3g+ngF+4j56pXhiRWOR/DsgCE//Y4fH2hBXtspGNfzG9JI+nIIY9oqiA94+
WEiEH7LbqMwMl5JJGkipH//MuH/o08CSETJhgUefkfXbzmxHAeJoWE9RJN/CeFDQ
kKR+roVMiy+cwTbB9SJHIbrMfcEiPQE++fJQUCBv3DgW3I2cxj6HV1WjMDLxjB3N
LDOVVgZMWwBgztC3XAjbZ5YIt4jGAdfCEAY4q67Zz8lMI+Xdp5TOtF6j2xHADPig
hV/2UGDOtLC89wMVoiT4TZvVgJO+BSK3uUoAq2SLQIlq2Z3DactkUyMIe7y7Jyx4
Zl9EcSkY1gkPsT422yYqPuJoJS4rYoGBln9EuXZUgCrqpd/JWgW7iEVBrd/ex65B
On95vN1HPcmnUtpVSt4m7VkAdhJIuigOK6Kn5zW2WJM=
`protect END_PROTECTED
